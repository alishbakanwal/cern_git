// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:02:09 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Ak4Mu9eQzPsriSrE0PW1eVHB4U7mUajR1Xa43IjBEtA7+wOIDn/c7lu4QqBJQKrY
tGs2RDdklStCvLDozg+0n/86WXF929kN8qK4Mntjzwgpry3p4Yeybu0njjoRNgim
YtPF6W/vuTqGK9F/d/oVfC2gYdAlqmqFlSm30tXaYBs=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 15696)
13ZyWTFOqwJG6K8mTI68zh9lpvwneslpW+5ciTqEdoztUW/BdFcSGS8e+zsWE+ec
MX0gE5UntRlK3YnqWPVd8sc9PMxJRCEffoZ5nAXRTaTM9V2CRSHq/u0u+w9mANc7
Ccr4Cg35v72oGCZktIhT5g02dMd9UroFnujYvY0YTXBf9U5Q/3Ck/CAvozd73oEm
yEhQkWtuFZelLb2lba61kn5gF7W/Df3y5TZ76ieced/w25pzy30R8CWFa1auckOr
oFd1jQvqysJzGunr5rS5d1H1iDXztV7QOceZgC2nXdFH+RyzzjAC7NFl0Uk3w0hG
0fE66rUNOrTqKPtKn/RobDzn+DuTgbdm5RHhs0Xpv9TjehqDuyPnxuundWHoW3jO
p3RDIr1vdCe+GvOBuh+frv5WHxeIOTPZNwEf1BSSLdBih7Vd25sxSgBTPLiQ1gXZ
wFhT7QtIqADspe5uOMx20yY5nTLzsmHfRz6I9n938xWxKMjfSvnQ0DtCd1tfnw5v
gjHBwGwLHWxjipEssBAYl2lPYY0lljqie1OQTqVIvNQIzmMafTCVC6KOE+2SF65T
t1f/2e9viyMqcYKAqDRs3CVxDmRrWxdmVifA2dhtmt5OT+GMFiJ8/xOj6Z+nyH8Y
+lqFUa/EYdI4Dix2v8LaW7CEAAL2BbhgEz2BweVFothWf2NZQPyuJRzXYyM20PGU
7bt/7KayFNIWYBx7juJVHSH2fBK5HdEicZ9A8R4HDFyKtzKvMLUdDAeDBbwUXKi6
4J0dX09rIT42CmwTbe9gb2feKfODCo70B7PT0PxXIPXKLBXwT8wcOX9CsItrzebN
MGJT7yeugZvAp/oRWd5+Tw3QSO+Yvl0MBQh/z6G3W2KRK8YUlX3tYOPhVhZ2mXou
Co0Lc/Hs56xWDM215eIoSVJHWbuK+agUu7pjbs6KqheTXcM9pFmGeHKvlwCsV0cy
k3XQ50PERHpJwjlris48LJu4NWhT8t7n7K9HEE5VdPY6i5BWcJC64WFqexOq8H7C
6V+tBPEomd8HdBzQ/08lQtrh39iD0rTfh6Y3AXPGntdhcLNx2j8+dGu3a3v+xYQp
qDV2S0gUi5cibbLKRXbwj1yfnMOazQflTvWmCjoOGVx8AEqxhMCI9DQ+9IeaKrUG
WzztGD3Zh4QwytEIFeh0aSAHQOJoxvP+lF2EbFIdSsPJ6fdBVyEZyRa3BMX4sxWf
KQDoggZD7H+11Zv0pXnrs5+d4NokxKb6Z3zZTXK/GtT1YyVOkRPeOzPZ2m7r4DYZ
MVoeisBy6GlTa0s+Byg9+9+TMDFxDQEqSNNMgQjcfRaxC2BUaJtd5Thv2nwccrxP
zAVQ2AAT+W0o5y9FTm8W/05oMemNYP8ZORpIJMWY2dtrX/vpR+dgdN0WCWlUgkC7
4hfSFu9ulURnH8hKZLQXbuYqXUnB6/jUIDFxkZjGiLGxjwsG5tteSCrAQ9TR6Dp2
ClcnNkKNwm5RrLS8W5zCZyUahgZkGBELdRwrO2IiyNOv+1xmCReIwRkMcia/u8Hh
r4LX2K1Ob2SMM3q40q9fXoTz/gi+7y5jr69JDoHSFPqvhwT5g4hHWW5bZEDCcguC
as3JzaE4voTgO1+Zz1Omv37cKMxerTF7sd51dCrZDpBmTCY9j2nutNXp49is4LdU
4LCEvCL23cwQ8Ub9dbKwUvILbhxv9pSBAsQTt10fmK6yuTMUEC+z7cXwZEiUGTeo
ll8Y3zDPTvcN8Fz7HvSQTlNdgsFtee2jOPq25sDA4DxQsYEGEKOOJV5MYwLC2W+M
T4pZJnukNd7/lJ+oARVgby+8T+gOkY+c1ki62XLwqj4Q5Sk5PMWcjYlwvxhAdPQV
CAYDKK/tIg1OjWxGa4C24KUyZqMmXoEi40qbAcPYwmxgzkpSFARJyaHNBFiQVrtY
YDEhDGoZLeoiGNRDd+qzoFHXW8L+wL5GhNP0Bcyi8OFxjTAosqPc2AVvtG7v4Kje
hxa0g2v82X+DdyOEeDTXsD7aMjq6tZn8w+Vz8FQ5Qvv3A78/gAkGlQ3Bri5jNSoO
o4TansxvpIkcDfPidc81gH4UGrJeuK6WD/8TB3RnC7s7Ex7NmES+OvSRDnDvWaxO
uPc6YJdX9yZXktDcDeUWMnhdIkmHIRZVCqx6ol3PRX9DMQEz/FOe27MZiII/6GkC
k92aoH2hOBXdm5kZHMOoEmMRwxYp1XqbFHPdZL6GXsrBqF4NSY4qctMgy41rQhxV
drLc4Tyav/ZdIoVOdWoQzi+t11ARcd5Cvnm/TU+PPV/hELsbUy6PP70s6m7bnYmT
JLM60KdErTFpvjEdpBUBjAkP0ABElDYUH1trMXCJa8QRrH84Wk/T6Gm/A8F5J7Vu
LCW8AizToTMkrooxcGQefGbqkC+uHdUTS4I8+Q58Y3VpVLeecM0cUFpTDJPuhV7K
haocUMtYoVNwMAkoUj1Yd+Ym4CLJbWY/AUWv+LY6z6fEMK0t+rzLTKNJZY/S1zbw
JvEFYxOIV7CU8kKq9OHeXS5KOZvg9BLt4JIXQDFuivzm+N/grkn7DH+9bvoyZP+0
HBsREfujBjgmrqM6q8CWw/jVF/evkX/G7/YUaESscUedI1bxcHsNHh9+56hVDHh8
6OHGdbYLbAckRF9H7n3kFN1Cbb2fZuAIWLg/mNxO73WhjZVBWwdz66grnkmH4rIz
uf9l8L7MEoehBlJvWGaMGjiwVYvCDQ9m7NXy3W5GUMJz2KWHXCcsUDPjbgKOF2hZ
cmu3HKSY61LfO71YbZBXZkSm4QBczfKW5j9MhWHCkra6a8/6fxc7rM/+QnOGxak6
8btE5xCtijnb3wPnXltxZK83IzrhPleJBSpj3Jbe9jk8vXV5Fv5Ez0y47oz7IOdk
7s28NcPSW1++5hZLfJIKI2sAqTAqrq0Cko42WHPnshCpcG3XcFC/463m7JE8D9Zw
uHkUKr8uLhRq60hexYtOVq6lZq3VAyvK5Y1/bzkZpoRQEP1eoW0kCTp92cTMkT2C
Ap0J8tzgwLJUE7rEBBf5p0BSPip/qmd1U8y3Sx64T43FKmg0BcI22UZFzb3Gy4Od
6TGTVYBbxs0lcAPILSdCbeYLdTeRJbL7h1xAKwbG5ovHHkEAlFv1wrd3nSELJ114
7ndVv1GWZm8jQpc0XebIRPEGkR9RO+9sCA+3QyBM6Z5D3EkjSx2y3TLeIeq7jU5I
NzNTlWfTvRdwHjJrbGob4M7fLUuSlo4ujQwQSm+ZtFqPqTEtY3t29dSW7Bep8r0H
ySv1e/1CwTNQ411I5IEmOxydsr34HYvYrYa2klqlTz+FHhcETT8t1mTeYwHkIL7L
Tza/V8SAGmBEc+jTPaiemSn5vpbB8iHjsL88tj4YpSpTlwDojqkpb/bc+KbLkZAZ
zKGwFey9wjEGvxeYikCJRbT/oNlIR/CCJFjsrzC664UWdleUXwiEMjzEAb9ubEGc
CbRh918HbPwYpzAv8EVR4+2puZWUHA/Tv/jgcgzhmZv3h4JKFSBQDc/9Oi6AagAo
gix8wLv5Hb51IesvmjsCF0YfY22V5NL/qHxpgtJHi9ibUQTF4Bw1Vqw99wo4YmQN
XsQX7Li5i97Bx68pQ3AQOdX4UGAPNxHLdy4Jw1otUTu0NvRGKy72IkB8G9NOrQND
/nVagfiSGa//a1pI9KoY4VWjRfDuTcNvBnNFBMpy/qgw0y13ZFmlrGdwyd1HM7OA
vkgOUlPgxylpI/vCa9UQ1jsVMYTc1yuREsnxahLkIJo9ujL8NELnQSwVTU2j1HcK
lCUklbn6C8vTrHrdGDcpNTXoyduDjkC2VHAQ0qnYyrlJAfez4qn41JDWK3Q+KcsN
O+xWBt2OQGCY0BiLYXZS1jnFVuNymmZeTKhgUjUPdlxKBNw9vTHPMGsZBA/ut/fP
EMG7lG0CNNVHGXhrRrN8M3z+RU5wRg35eJ4ReAUfLE+O097eWSwzyJ4DlpcRCIr/
gR73wd2cjz7js6YQtHAAQFuqWfsrh7qKfwj4lDuiFZHVzz39SjSeHtvxtDEI4ewf
SvMcfQQeNY8Q7NyCzuuXiDddjcVu+TgIOpaR0ZSfLnR5E6RkycW/TcKrl3fV6QKK
G09gvJ/iWWv/fqbM800bnftylxfzxuj1X3WTBv4b/Jc3zAWzsshbEpUZbyW1NkrZ
qql+Sq8IMgbQS6yrCtnawFk2kAwUF2yDhsMpOvSBWRJ8gJl/IDayzOgjzf59jm1w
+ht/xqyVwwed3U6iued7u0ZsV8vIuYdIsM7UW5cCJRNa7fOJ/KW5RGAMGVfumoBb
MjiuB5LfiRJH56xfjg/TLK7oslxi9qJ+sPwnkea7iz/z0ARR8eZNnHXwjmN09adb
1wCSnKaWz6qs2elZ25GDQ9bdiDVvqW3qGzI5JXchKtTi5WtSN2nk7KfX+w5EhYYL
6sw0lMoF9w65RqMjNd0a2BKQ01VCOpCC+GSJikyBe09V47hN1vMOR2xSyiir7bmm
rdGIU4WD/PmoaMHHtM26t037ZAh5fWHLZhZXyw7rKCU/C+Lr7hp9a9anljqxtfx+
p6TX0O/z4rkzJlXREfforXWTeVbmZI3aZoP9EXwGI1CnBmWuwS6oL1LntTYX26W9
U3PNo8tyZySZXhOP9UjBTV7JY96sVNjZ7YSckNeTZgNM8SnD4J3ii2TZHf6ATrEP
YQrKnFVrN+UsLegAnc86xojnugCNU9R0AcN8NZIBJOVh57tmQVfA8k41KJYOORSe
bhIZrkM96fVuPDjYn6+SDAgE5P6oXaQjvKi2hs/WoszFjtEEc5jfG8BZ+YLqPX3E
p+POquJD1wRfMwZepvqaQYDz39dlFXnWwG31YjL7YeiqMftSyI/9JYsRArDfXy6r
FvNWLddljIhbjw2cozwvNyyZuUGNDRtYRUI46fmnMM+hwWT7dz6gq38We/PV9ZlJ
8IS2AaqrCe+uPwaXduZaz11rCi+wMZdhEdb0bSF4SP6bdl6PL7cOOPVvj5O0sRhf
KclesCXWg0H+ZIOexqui7RqXa2Lx02sUSkXh2E4Q2qZCbTeAGstYTsgmiziOV90H
wGK6iQrqy8gMHgGXh+ydkVUcXVw2gQq8uAq9kMdbD6SqoQIS0OcEuV6El7oK0IFV
oaqI1fPU49R89AdNWk+MLkfRHi0cLeaImwEfszMOo8XZ2ziqAD+5mEnqSpfUhVIx
IY4KR4RGPmjCuvjcKaVoHE6+6cGwxCIN56e1aYgv/rEBxQR16hnxn9ZFK4RARmU0
9tcj5ejWeVTYrIG/OaWCgifFHvA2x+CJfIUPuPSvqhnCzf0yIcNxX8QsTiFY3f+k
qO6S+aOoYt6MMZFUfEd0VUIA2Y4ttlADLqP6nr52nCwcfZ9S6+R9tbXZjAgor0Vj
TNSKTQG29meaJDvFxTvHjwYXpZr5yf6iZEYGl0lhurZkF8Mqe9+R4fc1OO4Z83og
LvIxHiZy9Gu4ZdEkkLj6XuyEY9pgy+qOMWu8nLhwF1NV0HotAI8i8jv2lx7SnCJc
Jsds7uYuynYZZlwkGl+5+3APATsMHBP2E5XI2ukbRzShUT4iZz/AP32KxmApFR92
7OOhNFiYcNZur+g7YD88sZqE1L18FkCjTVrlMwpuqga2aPX+wFjMQgB07D0Jf3FJ
nIBavmAA1+ZygEOo05cc1PiNE+hPjE/2uZyGe1Phi60B9lC1Hwg1rKwSrfVJx58j
Uhf0WHPoLLDpNjahdcrjh95zRFiMsSidsHigIIkEqzizmZ2563XKseHDcuQMYNWM
n3B3Wzd9C7CHTljpj59+e5TurSV8WRpevoORRXtwGJGoWg/hGhnCF92A0z25xUMs
qbrobiRMwHeqL38wXESUfWKsT5iuigkeIf0jjQf3IGPDP7gYLbOk+eP5ACimI79j
FVcNtzj1u7/4o7+wtP5IVvhdS4mbo6sqDELdB9ecKlcJqsfBtDRPdTOoGYRaHdmy
cXWTZVd6ZMi9exAjmqeW6YpYg2KCfpa1HmFrRJFkBor7jqm6WvK2ubkuV/0pVQkJ
umKUCmEbIV3IWjraKoKW9ojtoJym2Th+N5TDQeTgN1qhyFDCCO2nex/iwyzve0qu
aYcSOuK1wRO6crTdssM6wHb9eLVYs9bIAnzGsPeLEpglt2GesYwPMq4nSl5vtZrS
6rUjwdiY+J4JUmce691yUD2Bm2ai/vbpZ0BC5pRkiXQP/MelA+rJmLabG2XNFFBs
syzcnvOfRaWjAv2JSZ0Zd1GpkGFEjNztmu8vEoo/7jOVwhnSPsCvrLhcf+ikKt2c
l4pfqD5aIHltX40LFsyW1hr+sN6HEsMySiwcm3/X8xyMDcXdTOuUM5DRx0PmQYxi
TvdSoJ96WcJld6n3YuBOzX9vqbobib1L1LpedAsE8yaEKp8D3y9sJsmZ61cuuDWf
de7EAArb6O/rQ/WlJG4qq1lxWqR8z9ueYIlcxMQElSoYFGQZIWyJGR5CvmUqk6hv
bUZyAUpV8+faVejlmiHxOipXejny5C0gnt2ro36+HUOL1MiNwokUgAcXDpuWbTmo
20tUudbr1fL+QfC4FjzV+lGO3cpHO0JdaPrk4HSlFOkGR3oqj+LNHnjnGHB8Jgpu
H2fwWDrFr9/sYwpRmn/fB6IPZPKmgeHR3uFdyem5dfx2lRq6hJ4Q/n+1wZBe8ZOI
aS93eHHh98P+jtIbaIg+OszLo4cV01Mv2pa+jeMyGZMrtfuKLSmnGCVhkkw0+Bms
rhDEuMRtNqhyGeDi2UKq01JloYgL9w1nSlt2DekCuZ+V7WC88ySe5EdCvIXb8oYp
EJqdmPtb/bwDB86ZBe+tj84amFkX7aWNkpBnYv2Ac87B7iRfnDGdbowrw/qhDv84
U40AzTXkEH+WWbSdfcpb9Vuf/hthB+vldESih3JnFZTjOncNaH20iP+sDG6VN01q
Of2apTTg+isd6U4pzA++/P5j7Z6xKT3CckdeXt0H/mURsYO9aR/mEmym+9nQDYdV
cYrxg+l+Zg9eZEeCqYidPjmfEbdLBCWkW+OwKWDcnULkBCAiPFL9NVAmbjG7/RId
83ns99a+4QPY/huS5+eSuP3qCeqGUV4PRMDFClLzROaS/ApqVDic0eJVF+QjEG4R
3PEU3BWtuvhEcvMadCgZ0LBSKyMR3KVl5MSGRJY9urPQHc5l+02B6/9yRyTWWQss
d20cMK2U0jWPb7D0Y9zIaYEKzJzsa8SunuHaG2DF9SnByTqwY6xQ0zJXX5vO8Fsf
1fz4KsZicM3qgIh7/zY26CUtSoURkm3+BxbnPLfKzUPGg4Y/HfpfhuTtk7BZdCV2
VvQqIfMw3WaMPZS6OQrE498Jd5+bgLrNbt1pwY0BBUHEhWXzZ7hQQ7xcqpIqJuVp
9JDzAWl5jwpU5a3SIdiCFf8Et+NjF8dY5pP3w2ojFMYxVFSNJzTaMANQqZvG23xS
euDmqiuv94g3ByDW3ZQvqV2bmt0FrdTPsEMcVZbA29WBlxRJeYjUeUMM6HxgYJU+
/Jbx47ziWsXGnVuQ9Koo6DOsC4iaxaF+SwpwlxcEZuY9x3iRAVUDYweQIBhi+dHr
1acwi9GM59blWK1sux72q5WL2Mqxzk599zzEOj2gV/eH5dtYwA2SUl8P/cB9MioY
paeb8ax5CDXKeki0fuYgqFiODIbUuam+BjoaPVVGYeP+GpPznARCEhHWGaaWCugR
3EmMfxv6YcRuGP8CkBzrAbDeAGYSmWx+mH94hP9pUHiwYHvxB9pCmdtArdyu3H5n
saDcJ/q4qGddT9D6FgR/VVv4D8QVwPXBEXeagRb0CPjKt0jRNnqjIzX5kJZPDAsX
ln4DDURYmYZ/oPdxHn6gwgf/JC0JT/i2tJ6jWgasLn3PvQA0hkOf+jrvJLYoqg4M
3volrMRZpnFRBlu1HniofFABPh9KGJrQX+epVK2Ri5JifqdPVeLBjwaWPWITl7q7
rNVTFj1Tpa56c7zMTiYcp72khaGkeARoeqy5khfoaTBIIhBTZFjK+td7CB4i5qH3
N+hgo9n4CT7PvZUNk7tfNmGEfZlQdAxLabQYTNjE4in+1G7mft3so7Lnv33ez/1D
8QJDyYZWEYmP/p8xP5bGgb8igDTvEyF9GLQDetnrnvuQMk+Do2ChHRI9sa7a+TF4
CpBxg7AlDS3NrX1qj0KhVX6gsY2L8Q1HQz3QjOtQkBg2/8z+fAB/UBswaCRt5GTg
h+oSx7npkJZ8UiuMJ3JxuMdfWAOtXPdvCE/FbKL5vH9fkN0k+HaiADYVaLfvaUMv
+nRmeazEXZ1vR9dLJL/EBDIceQCXPPXaEKF6sac9EvQ/QkAtqlychMpiMaCcEz2D
0dfPRYY0QKaJEMFGwv2Igx4yIi8rvAyzdLxP+9QbxTGh+uAp8LmZI//leuA2Oc0J
fbD+AskIQlTeen2c2I7fTR8ut7qxkTydCdUPhqPZ/PGwbdU6/2TwJLh3usb+Xbhn
GtPlEy8dJmXoQt6TgS2C0VuB8ssNvbVIJz0pRONUxkQp11zrnglua2RHQRZhTjfv
0icRUme3gTgO9T/kG/Cy89TSnInEu7A2aZ0pbHGAxQJbwO1/cz3tW1s6AapVgtha
1KYC1aGvFludDdVEXoLA7eLpTLcsSZ/6HBjSDhT/BiaKuRQXilhYYvrK2mCxQ/c8
hpo41y0L3CGkfnIYi84fCw888k8sJkhXxM6b307Y1XaCcQmFois1we8bCeNQVJtO
Vb00mPhPTMDqe5jsQlKe2HnRcF4HGXmmw2XhzqZkGwi5WGEvdJMFN94RupyHwqf9
YnjIPmAZmL7ZHLmnveZvgzSkbySdU927zNTQVnt4wwlaKCT0KyBfpveksHmZIbHb
k9jMYcoti8cXSNC8kvDjuXogszhcFhBr5iCKLTsjGfAOPtk2OnRN/7EbJTn2CUHk
s7fL0t4KK1BO0yKU9Xg7gQaJ6vH9BcF4JwlaJ3FLjp8ZqVBKMWChTplK8Ho6egc9
fUIz3ykApsXU2B+uSuZvLw215f3hW6YutjattVvfp70VXfYk5AxRToBKK8Hb7s1M
7++0YaR65jXmxtLNqwubTMLWC+zisAkGvduPLPFJa247wzWuo76ibwXufeDVMz2+
DR8Ww12CMYU0q2w3r7v/IhQzSeDF7ooi9NmZV94mPbhqPzPJKwf2nkp7LYuOa2Ll
OQL1WvEQx5bTkIm1L2tApTSZteQCrIz9GvrfevV3r4W/cNgdSnhs8yUziEoDIiIb
K0yKQKupf/NA5K5D5isBYM/z8RegQAp+7at+WWPzGslyKcUP8DWyA9xlwHm4mWgy
tkfYkQtPStO74KN/MjB+rB2CHXG85m9l0Obif35Etu8XfNrGM6GHh9rtuWDozt18
SOqQIdShU8UpQvgZjdp/lElQ9Q3rYPc3OcIIDJ4UpZ6X57LwniX7sjrdvqBUIkL8
ZBo21sXZhN4svcW4dPB3Py3F7QrluP64U+7K9zFqKkcQCLytG487xQiS7TsA7wuQ
NgAQyiw7F8AjnUXBJlK86is3wNoFjUK15HWafx+fXgNVNxgGJDfygj3nCFyYQ2YK
n1KEmq9K7dTf3GmxK6LV1RgUIZ+99lp39wRYa7jWcy1q5LeLauMx760m3jIdfp1I
U4vVAsOTnOg2iTau2T6HTWE6LL2XC9HgReGIX8lMleLjqOS2A3iRyZg+PgciAZfy
PLmPYZmEVVlnglXgP8wBInBA4A+vxdURnE9E1EB5PtXGwkpJ5tPFqSwPdavAzbAs
p8gKW7Wlxk3jf1Rif91slWzY6YkSz8mmGP+aF9kwSGUmAPImMyAoqfzvaTJH/zul
akuqJzZJdL+75gs+WTt0ZIMzhv462R7f413bDLEsWvpsHHkjLsvt03l+qa3Hgsoc
/A+OGa7kF20GBWVJsHhJ2HF+ASbyXBt0daiqs/gPNjRFHKA18/kIgFZ3UXQqlcWf
Jdgu7Ai+ipiu/7fl+5zTolT5WlsicBjreG34R8bOGpS87QIC64uSBTdDmxJQm26I
PWYy4m2bfUG4i+ipsfBG5I6GaEATNFUxQjFfywCdfETjIdd6gjTEftt2um7yRsKf
4xu/YOQxH82GMNlIOhZR7CVfQV2EU9JsEOtraJ7YA8zNegtWE4Prp/jvh82VRHtD
jUfM5WK35u47psYKgyR9FrArUjRvOFoUyVHgg2MAI1AjnqKKBxpMWj55fd4Vhv/8
lHG7JpQ0Qg81voY4VjLGxnUkeVRPFskqno/1pZsn2HKS4PYRVgkmPvZkFbykYsBb
GnugzO8WoBCQNrZTOFJ9zX7DIRrLPuIyQvalLHvocP2LgUWOPUnUu+cwg3CrOt0u
hyJHrV/e9DL+ilixUOoIpCFJyG413GW9hM7ywlCDDrE82JWaXq35X+yEUnx3DHcE
uNYxDY/MqMIy58c4u1SgMpck4RqAQcPAXejJINyXIP6pmrtWk+0dR6HgWlsKf3yl
r0ZQZD6KjjTrYieK+f068/XBqFJ9zArRIlsFVuQsTweWzARq4J6MXgfR3h5mTITU
ghY3B+4CachjjYm8HtxUIAVyKzrfrk3YtSXQ3qdx6EGR5wH3z70eJbynP3/BmigY
p2snv987nzPOnA/1pZ2Yz2BiQCiZgpNA/eq0R7YLS24LJzk7/y9iNJu+YSvzMUVA
V5tUqXNZ2DTtJrkz6Ry8Xw8qggG4eFY2MegtOlW/Gi45Q1mOYTUW6UfuD1IVm/OR
3pQMYw1rW7SGPa/Wp0CVNOSTgGOHQBEvWCUqwLNVouMW5arzIbICT1rU1a27Exkl
+19I8mTP0GJaM52+2JG7RUmiCe7OANvLpmAt07Qe8uRgm2Rs40TQORjOJUGAdueW
NW4g4GB3NkoXMgWyWd+4C2YkH93zurG+omDNlY5GDe9XEi+50tW9sLqiLPzynm5W
sVTFZwQioWprKMYRq8aEPA2sRfg933cI91peZvOsYoIAX/EH11f27Q2GupbbvcIu
PWPrO3fF/LhJcVqManJ5Nlzz0+iwQDStfkGEi9WggSvXhuX7mb4ZsClFzdHn8Kc1
mxCTSH0w+9Vv7L7/cqQ/MvwMIhYlCSWRj7cYry5aptN2uBtg19XfNArsbpColfUT
POIz4T0Tmg/ZuycOjaNKoZAFC38whDCeFqIM9Nm1K6UXvPzGEvF9xcxedbJBAEHg
7vzXz566i7Lk3ykdxCvjjnPoWrnJD1sqmEQoquvQzXyKnlof9UnO3SNR44uDayev
q7nX9ru1GjrHnZmBHyGbc53m6+pQTt4FYv0LfdRr3EdX4QlQlem2LQAY3HNfQr8n
TT/OzwBjZjM7ed8gp/839lowUCDo5J1rNwCdNiq//baBAY0fkUHtzjlejGykwO5D
Wr02TFDY0YYMQQOH0a9b1kYfzZfG7DAVfXVBoyCaLtMj7nla/U6i5orq1YKrEx55
S5aqzf3C5Au0F0YVGpmuVwOHlbm2ErIzOMj0g2XM+AhwEkTq1Surtvv5TYOqkDnC
3jEpR8tmVkDrkS3e7w2YWPJNL7w07ZDtLge5I1UaU5iaSQ18QX4BFZgeYxTmdNve
6LE5TiiG3/uS4jpceLdUEJTqgnhlk5GZiFW4TktV9A8PheLQPjaBkDytrEWKVzf0
2aLcyubkcquvx0H7Jp9SG2MS8rM+d4klAgRsIU8Dwi+RQXIjfvxWhAPQfZJf6WxP
kiLjDqT84K7fmlBLjwOaea9IJUBfC3FJuSsTdiO2BO2kLNLmrw6P3TmONfFG0sjn
SXaD4nLV7bDiYFJVCkGzIH60tUlVOv5gRi1uCC7/rOmtQxECyiMjlmVHGIEKhDDE
3PISCl1QFN7SyaVZ8pDr5oJTXWanSFTD1w7OkLSTNQGfUBFGp9aPeita1lg2ZCBH
pJqD/O6KiOu1Df3OCeU7zVx3wLHmkUBm6PWDH7XlMKbNwzwMVDEz97eb/7klGh1x
fyWAIrmyhxSrhX0OEMGBklm1lsrJHeKStQ5yNfkdh2KVS3itviKleAOY4BjW6KZP
QcM3g8XfsQMmvadxDdH64s2I6IL1vMg8MmkLG4kUGXNZLufE39LAtsKh8UpZoDEx
dWr0BT7zxflY1goryQ6aaZDUjgaayVWv/gO4gtB39L4qk3ElpSu53X80v2NuJl5H
xvehP3MqLyeptzEKhN+Y+rjQkoqgXVM7NYGHk8pXeGmFDm6wL3Z3mbdrHjLtdKL1
8U9/qQk2rvN9T9F7pw8RqNxbTVH1i6pyCVgVP2BwQ7CPnVeUa3qH86AgGHz3bqzo
3Xy2bFGGcPKUqyTXkj3Qeicg+GskCISbw8ClALYsJ3qQ8Ejl4d3Frd5duSCUwT/O
UtNMj/VNR9DKJ6j/1H6zETJE3EyU2PBCVwS8huKB4ybWFGA+tNbx+dC4GxBr8njD
CJgONsEcJrz0CB5X3gRQDEHncmHIkgMpvl9hffbwcD6IoVZGKr2WZ/MlIuxUSa3E
AxgPLDa2TtFx6Tsupd0wFNZUh4xKhO4kUSoY/JMSIxM3wmLzB4OEuzzfyBlqyy+c
wlcb33CT6x/wn+LTO+y9W0IYG0DT2f33KMY9WMH21fJHYGard3QkYG+TXSKIAw2x
7IXzfdWoy6LDz2iLS+ISS8pV3Tq3arSdNnAALDWLxHSTJUVexSCK418+cZ/CI5yP
lRKC71plcU5KuAuq8/NQPDxhRYhuEIlNZyVyzhJ3XoRIOh2WHbfIUae9N8aeF+vM
MT0pIFx+pfyQ36rQv310PWibZBFKNR1mB6NMdA5SlJK4quCO40nN2prwmJkDUaH8
a6p8O898UczQ1wn7MiZqlTY/vP0XpPuDHrTZxkmPzamdnM6Lk3XBZkuTsqRX3dNA
NnJW3YsCShZEOCmN4yL5TNuVM2x4SJo4Zcn1gwv1R4ClqERi/OFJBt+6q3Hxgu5/
eBEB2rUlMtdMRhERCo5ODwZt9T2mdHxMXPoLvRumJeFvoNgI7BjNLxffICVjsyup
RDu6hOLDi9j0gOiQekeZbyll0wlcFmY3IUwN+SWlaeop85amxkWXZKjP/SWiyFQT
imOfSYoWOF5Xz+q+6urGKe6Z1h6rtv1ERVa6Jax1jL45r0ql/EkelR036BdVTJUd
Y1WWlVc7aU65QAH2Igy5yVnd9wZU3/DEo6RwX18m36Pn0UtOnEq8Gn8Boy684VDr
TyxFJk+Hc5wz2KOdnilM9yU/e0dGSpxtypQjmHt9EHTjNmULuzbj8H+DZnkrlGhN
Vaogl7BFV4jz6y23UhYHAJvITQzzsWFmG9tMQ/jLTU2Dfw6nyXkPkcizOxjDu9z/
bllgkfL9NNQHLVAv7yfN/Eojf4CWdyuZ0cEbnRJbdu1YlO69yStOTmVOxY/a0EG2
uF83vQ+7lWWQ8X9dVy2z/RQMZtmh2nG93OvVzwDhnkzURdFgvaw03xJ9qcgXwd3y
meOuhrM45s04u4eft5LMrLCFzPIRPoAMHrfVWa1KMM39/oWLygbZG4t4ocBByIj4
ARzOf3dcCyZsl1CanqP/XfhCacml0gdHbSKTZeMl7CcD+YVFhYsz/IJXZVv+KxV/
ROaUkT65FNQBj/FZHlRwOQWgXXnkVmSg1FTfu0Ftj+aXMMJUZLGvSMLHlwfJIT3f
0pwm/9WRbBnAvJsfrK7rOSpOt3CvuEF/xv/y9j1qa4nGVNoZTLQY6MfuHxS5oHBu
T0pWh8QrTDlzknPF66yne05GAxZLRyWUtWsSFtV2zDckIzoJ4E/+yrJNg/imt4lg
Ed47K7yLhCiV3ZiL1EPFwd0i4XKGmSAnU3a8eVDvf27NgzQzvWvqqJq/ndsHAuOF
oS/grkgiHTITnPFOrSd7y5j6Mmhek14SknyaZrwsjguOuSZH7/EKSsl1z6ZfrBfl
KSTWovqDDagoQssjPqw4OvFgN6SaUCa6KBcHbA2ccBAXen7ZK+1mdCgPeL4njkRV
eDkA8sufgamyNkNOiWsxfer6vFPJqHsw5mvcWrY5l+DDth1xsEmkKGvkwEGEFZim
vPZpfn0RNETZP/1SPcwEbgSHJvDlIYFag7nhwM/uolp3WMLmCMlBJdJMY7opw/62
YpXS/g02dEn3y6CIBgOoz3PI2yWMciWY9ZRbvtwtsmaLCPSTeBnUnt58FcndwqaP
siYTwe6CFNSsjUGcxU5HzHHnLeX9bo+fuao9AEl/gfKXTky2oc6RJV+9pIaonb7T
Qt0Whi2O7NfXRvp6DwvJCxBpIIVKBl5ta4joRNJCx+qwPy+Xbj0JQLXz2uwYWa0c
+ZwXPJD1k2HeF1TJqVaJ+EhW/s7sevg3Rn0RxJ9DgqRqjBbJUJDCwMk93u08TZDn
h7QXfnlXIjluo16bCWkVNx2ciLQ4IBDg85S2xpqgexSSZFec1/XYQmguK8mc7c4H
17f0+vvvmmtiGVwPYNEhCZz9Ic33JdWFVtA/nSwUe1NOB4iYa/9Q726JzM17upfN
3gYMiJXEz9TFEz3DWmt/j2+gYeFnZmeuKcQIKA9wV8pFO28YtZLeISNGLxEE/Ueq
VItoIHSQbY6GIlTzkT3j7f/Kg7UqW0IxizRnl8bBoPL+afyvvsWCwc8xCyboS2yM
+mEECV2iWg828eZHHa+PQipraaYLE3XnwmYS0Yeroc+zTtye8dndnH/1o8k1zewQ
5kJpPIbkKFzYGzb29gcMc1rG71xMv/a0ZG1KiA3AceBHNIRQ+E3nNiIKC0JrBcDL
DWO6JV9l8vVQl2qzavdfonDi021SWnkmnf8BnbtNNqemQQKh4itVWhg8o/nfXqXZ
mgmvHQcJkSqq+hmm3rwGq3iePBbofsBxt0JOgyCh2RbRQQJfZjUUDHLM8wNs5agE
p1q1njzWyOESL4QPsFQTJ1FOKmTBf1P6T6rVEzIpOKm1czyyiiFb4fCS+cWXjJjY
zrf0acEJiBddzbhDWuBhUeRI6qK9pDuMXNkv+rxua0v/aGkeoy8vv0peq5MIxmhw
DYvbMdOMtXNeIO8veVL4iZ541GAyF5p2vY55KuxhZItP2Xn5Qo3ilUr7qn1o7fyv
/Y2OSrxPpmHfH5ff9JQnOuV2nWmTOBCOoO0SY9QzoyqWEvrxQHTZqqnhWF24h7dr
ucO2IlFrgu5zoiw3Qc3X+XQ5LeRbLtD0J7ieEjjA/nPrCyjHlkwctxEsauTLWRnk
VvQIedUNCJyaHPV6rzt3O8fNy+RTTxxJoXDiVD3/EyDXv3Ye9wTFKxGmGwrqPurV
ky/v89zHwdV4E8VPorUUJSNdFK/oMGMSQ5F1POeh73FAZtNg+tc59o9GcMd3/gqS
ImGWR+gunW/rhbPJtgr4ejsmq57fusMMZXfFUirOWLuRd+kfrhN4uUJndqf+GFu8
aC2ckeqR2HBfqHoGySwbjoB+16l3u5+FbxRp5YZcxiKkE/eONPf6xhW15StUua/c
EKNypXsecp6iwKA9vnXahs2mBqqla/uFi3NJlPkVzyzhsHkTQYU1zb0OkTpuvFXE
eITpX0Tlr+vY5WHixMHxbtZVwOASU/MW7ykctSIXWmfyRiLY5s9FWfOup1bm2mHl
1Yp1t8NIHaxtyUN5hfbc+ZPDT1B3gKFxJuY0wzorJ9bQEZmneiL/yLQQR/3Icxjr
HSl3fpJ+9D+QBl9d5e5frQS9ZSRDYfLuw/z2Q6HvtSgHKUZApdkQm5I+t03CzGk4
GizceesAxy461oxfajA10BYCe70FebwUwm/6bIIWVAvVWAVX9LbvYwHszyVKjYC/
WJF4RnUrgdlxE0U1hGT3i7Yf6SLDUOrYjryiF33mwOFNF5+ZgNJkVn6pfa2Igpbc
NAVQZpuZPJe92p5dnkfBlcWX1iqSzyl6GJKOsJ1GaBf4r0H0PGlR5s81o3Ybze2f
httTlZLzDWtBa2XxARBxx87bxHiw7HWIBJFWyJJFiiFvLAv2E7W2f3ge6LjRkkJn
crJMMj4XMvMn/s7JEA+nAKTciyp4uf8Q5G5z/biv8rK1MZ5g6vB3VpWN6ZqzPNl3
kQW7WjTdnZPic14PSfKrFyGrqUUH9zS9xpHocEeqZfpeJI5Of0EpawCxEgRiBIjQ
l9l3HkvZrXBLsVLoqdRorRqHPjJKZIzwb8JhDxWQytJoD3kKMrhkj7BO3BMLkTIJ
eUARhrd/rncf1QWywRpCz5kP1//dXwPRkHHPLc05MiqRDJw8GJNgGh59D3edQPGJ
FvP9GnB1XNfcbbRlmVgSnyYxejtfYlSVWNOSBI50ADNevLFv+wbNBQNGbdTf+qxv
fWZFEQmkBTnJReRpVicpCFznLMJJJtB2fM1nQs7CH9gqBsWaSRDkf7dw1AAEuYrr
nnUbbD+tE6wG5s4s22SnJ0WJOgsmt++A4GpP+7IFGMXh0aG5Jn0GiMaGMTR8pz01
wXGgdQQqDfhehbHyk1isr/4y6JEgidOj+beV0bsT0AQdof6whrnUgdeimMDT9HIa
NDcZ40olFvw5XMW8+fupXY51x2lEzY7eRlx7zVEzOkmqwbPFV9qJwpxQ2IZNeIRg
kdAxAQKRf7RqIrZxCzwgDAMBDzq6VWrYo51+8GZJY16DNBMEC7hiBkKz4xNHVHnQ
rItTH4dPUWhhQPKCopzdE1nhkMHhbFv7T3l+aAx6+wx4pgJWRj5MqFokOJS6iujH
fYVAYaECzb4CIXVlicLvX7MxtZXTgdt4ergAN/gtrj+eFgW3nW2D98THj7JUFaZ1
C9NcyDb0R1ESJBOXHaj7WdSgKUihwr5VChoalVsbnRIogaUnDKlY1LPkfQ/v9nh9
+wxNe9/Zn0fbYmmvSKi0oV36t4YGJ1Xo7yQdxCetGwxHMG7agJlFgyhh1ps5ReFh
QyP2neAKyZoYfnryht/lP83r6Qb5jf9nmAy7eDdujnDdaQbXV8YyOBL17kaLu3wK
xerEJ4+Uq0VgKhxN15d//k1Vx6jq/Tpcw729tK7icVRw44g8PJ6LTzVlpOWuQrPl
vVV8//1vVf+eSlltKKuDl12G5WEMRXsqcpVON6QFl0SUbELFGR2H2te8B/MIGrKG
H2LRUKHsFL62WBekOPo35Zyo1BgBnUq/cmvP+HLOvryDJFfT6fi7YTBKWWk6ffMl
/zcYh2rz0du9304OR/AKPtmVV5N2eB69oFsecG1vCi7aRVP6fiahE2k23vAPvTvU
6DMMd5QCTfN1520ZvL+rK8F45udMVgdTtDhNyUzDmGMjFdDrHGv0JDutppLp6Er2
yhYxAlw1iUoImPXFm+AkY8Xd1Lh2p8WmbgN6c0qidMouXWOgteyAbDqHZSVYngSt
CG3dO8FZcxIF1XHevsqyEnW2pH8uSBuVehh4bQn07+NGSDDmjIzrJTIJdYkGotMB
yIH/XTSPmaD3oalBuJGx7IUhBW5uQiO5T/lvXLMJvuiJrGVeSVKwN1IK5bDascBL
8t5OTozK0ctNi1tqCr34NK6tKyj3MB3/UvOoexfJtcFz8v4xjGQY40pk1oh34fb4
AXLBK6nY3Roi0dfEqRB5SSdF7eV3eXZ+u+E3C2Ppj7qMRS4SjZJergc4pLx+fHsH
v0ObZQsFq1TiRiX/LvpH1XqLOuVzRceK40FzapLpdqG3mOPf/JwDGBZAyeR4VbdB
U5jnOsQvisCWbQ9V1kDxaO3jfd6r2oa5qFnn1kgMrM27pXB9oNdGJ4R2j1q79v7m
BasaYskqQ0lQlcXmcLVFwnFjBn4ta7A/kFtEGfLPamgEncJ4BdrFvGAaYxd5U9hU
tCauZeOqa9aj50ilHXK3gi3Tkb1XVvbuW2dyboDquTEoLzTbb1fFQIWIsinkPMyk
1yKSePJ0IXAFyXADXI1bpzFk3sc+sX/4vGRTIpcetaUPr0Pvm97yXCOj5Xs27kTY
ni6G1iza1496Du2aqzqonYrx5cbzxVpYKXZnq9k7d8gOzU2ZMbLBuBAsM4M29P65
6/GGeGPxU+SqN60eus2hE7LE9g8joPJvMnE4kGJK+AVUoYMe7ctsopvOYnDHPUdL
wZFUiBoNbUbxKWBae5lvdLTN0x16QByjy57tJtJM0xrbeCUNwITdrA4Ah2kCTHRp
jFXVwbV44b2YWWBCUHZ1QWcHlkQcdRKz6IVU3957wb1Zk+BKNhKWPn+Tmxb6fE46
39d0Ynn4If7w9HZ3k3DzFNf1Wbi8CCV1sFaaqx6W1CwNTOsJ1DMYW2j02C6L/+Cz
6VTyC0evyUf5w1NTUfENox22pc4AM+yRLDZUuUeLU/zodUJLwKhITn01MHpGhMyO
WxL1mgbbIxinTQAW3ZD1oa/XJ4HVWjdXNNV0jqMf/3g+q4fPc6O14iPJGMYYM5uU
FVc1Gkw/BjZsMV8tURD0r5lL713bnDQYPHWHt/Egk7NeDDKV+C0W6di66Wfjg6ou
SRWi7lHBZ27H30z1Axu9gxCYiYJkDNNNrvCmbql6mSlHRYsdQnzKOwIS+3m7RGax
GXyDSLOFmBJe5jIGel554ZJN8vN+dep19YMVPoCLQwvgUwE40ro0qquQ0neT9+T2
mW0zfNG6fUz3wJNqKQZpleyASQy0JW84t2e7ARooE3BF18uAktC2NnXz1h7O1SgG
5ouN7i0YF18tuLc7AYqsCI9E3vsXUFaKeCZID+cBhvEXU5zNSPfivr3/UEmJznm6
F2lamuiV0v5+7uscF+itmOgxcibtJfLwKFa3f+mBpUcNrMTYffPG7exALy5ghRw+
Hf0MYUIZSSjlGP6x6PAxF1WC4zgKg3AcDLdlmHbRcjxeTF5CglsKxE07Wt4E3Bbe
kj3vuRyQp2fajSkKAaNw6w0gWcK4yuw1kHveuRrfiA/EJnozMp4KhfaEwlyCBTLU
7LoxAGkh16CoQK5siUJi2vXKoxwRRRQtuSANS45CsrMn0V/8Ykve21QBS8KBhkeD
mzWXomFoYDNo+CgnutXP4atIXc7zxU0RBevaXJcowxRoMat0Kmx4bDnMOJFsGQa+
ttaAkW5VITut7GgaBeDurvPhaH9xMTbhmJkfdkXf2Jnp28GUxrOGmdxhd5FkpB19
G78gxsndpVlfTs5NPrFw2t7fkZQ68/WFtouTMtRE+WEL2tUgcEZlUvkECX19vdx6
UrM99SIs0iXEpKYC1Xr8LHA45Uw3HIkwGPKXbdxWWoSbFSf7yvwpuBkSRUUfyjB3
90g268oMfpagTu+7f0acgShszRlikdVonRjQzcZQqFbpz4Gs+v7iGOLkN4Jz9qQz
qXpFltZO2TM04p3mMIZWljrBeE7miR8M80FtB5KvLGTvgN3jQMew/8HomJ11flt0
DwJ1Bfsm7MyPUco55oY7dVqdWUD/TMubKGtt2H63UahsLTil5xw2rP+CTBB6YOfZ
jANO8U8j4/u/WbjKv7y1fR0Hto1Pdq4R4Lbe/16V5gVKfpWvpsMs1H+XEEFLvT7a
wbtulpylxw3Irqbs5gEJjI8W56weVqOGQITNTpXNe0chXJd0AKPvN3jwFHrjNYpo
bb8h/D4Nc2M69nHFm/5H2a9RskmChSvbVjx++2WqIxpLp1GnwfIMHhfqzI0nE/jp
n+gwnnpzV6TNW4gu2BLyDwaOw2rS1JIJ5gJEbTOjpXSHcOADrQlkV0d1Ec5i8mtO
KWxQHNnwaKTOWX5oDWYVNSUq+dADPq2nJgra45Sy9vWXpavvxCfMADPho18a6E0b
vZeHXt8t96nf1h+kiogUh585XEioSF8ntBHkPDVO681o00DZaJTCIDfmPYetHb+b
9i2zNEzGev1ePTKCEq3SCb3FhbmQWGn8/T2qpNfwyNsB43OdmyibBc0IkxUZGcQ/
l5D2KZWqKtBe1DIXsOC1cnR/CFHtNDNX1JfTNAjFQkkTteXQaf22CJxUZzlGY6i3
1YVvTMKNCbi2+nYWqVGTncrDhqfjARVJYF3n5K6/qg32szEgVqSLB0WuqJStczpl
bl5GJr9ahLt8weiC23B9RiF9v+bLGX7M3HT6/LL9kcvADc4ti1AzlvqF1J93c7PQ
JG4FaF4Mtf9KmYJ2QCdvmdRb8UL3cAaxP63HL0mrsyDd2F9TEPHFRu8qcetUb08O
zu6gTcxn681lzRGH6qVcmqcewuSlqkeSGRXsujEXmX9TZAabIWWz40BGI0eTZsxo
dPezCEnPtEtvnclkl0ELy7wNMafIgUagpy2FFfv8jfXDN8xym8rGbLZO7OP4R3fF
c67sq5wJIUXGZejuPmJc63f2inbRI+grY15ilfd11ES2Gu42vRqtqfjmVxoL837b
IntqPOoOQUF/+gu8k3uzouMZjKENBzKniXohhWSlP3dWjeIyflVk77P4LpE9T4eE
b2UzRZzIM8zyldzEoyMA31XRaaQ0z3B2GZaPn04kjZi0xmEw89eCWE49anIrRwqb
JVKXtvjokLdpI93mG97E3hQsSyFLyWtFlGwxo57xpsRyCvfavd7+VbhrEGuxJi9E
ImYfEburOz8qzAsAqfJiBwljP9+n05tAVIug42CbFRek6z9Wk6o9RuTtasan7nPX
UDjHpqI0oLWptprxWGmUVxg81DtmZuy5GcksUcoORqpqgQuFpcY/1FZFymJMrQXR
rEDtNvXfSObrPvvsrs47EIFXFYpbn7qrpVj4trRlLXxEZjFY8JH7bmDWFuW5YJ4O
99gup8edG0Vvz8yk9od8ewmw6yImjeJ5iLdDQ3wTZLVIrQFwAuYQDFbvqUGcmHj8
f4eda50zFUdU+D8+jlSTMwoCkRDOmVwnNZvDkb6hMoH6vXiSsOXqGjDVlG66k1J+
Z14pI0ylrXmO9zjZRdcP5HU+SxbF5aJiaSdZZsHLWOHjrE7zIM6exaig0jc6Mhxo
8uTMBB4DXHDOrN9ItDIP00xSYGM7bpEuRK4nbCYU7JsJ0hTI+VkdC8YPEn5hk9iS
vvURsFTnrXbWOVxEicY5mzgJoLPkGQE7bTcYqs9n1zvk8fwV5JTollDVOAb4RA0L
PdMT84irbm7NiZUoL8W3/QWTVeC9xEeIwezNOsT0Y2SDkFMl39TKvZJExj46xfx9
`pragma protect end_protected
