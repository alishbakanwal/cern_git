// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:02:17 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Jw6DQVpvDDgepSJ6b8a6SMlFu69ZxcnqaD9dO1mA3uN+o6f2IYnf+REDhHPOsz2I
Y05PlZvKI7AWTD34usIBQrdFi7rUoK0BEEPAna9V+R7cjA6HTzekeIjhu8vc6utm
uQb7diZNR1TtnCNJXQSwCeyQWPWj54ter9dsEPwtlSw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 28784)
BiQQHOfvRR6nu/b3Gr4aNoGdVXO8pRxVj15Y6lGozz6SLn9FkkwAVekjJQ29wRkN
nD6Te/5atWlHcXnQph/vSO/dkj9+DlS3D4ufHRco3AcZVpjxoYltNmbGbV+W3NoH
t4vaLyj5Y8YTYJgmjBIPESyp65gwY55LHRN3foQldCcVrlsCsSThS1IaWfIirQ0C
dvCqyUkrQtpVqQzRHlCInyWqFxkbAYENTSX9wsQWr5spDoIzOBA1j+z1Eyi2BbJS
6qB70Ids7reIMChAUOH7uOXi042Cwu8XDehMXhFG+/oKTRU8I6KV+3BZmBN4T00R
BlovONuOXN5fpmj255QYfR0cRi9MkTM9wctlUuZyno4rdk/dA1/f+27TtT9kiibE
7Hh8zfHBQ1YoZQxdUOu1ska1DpQnKTRjoeaoHZ33A4ZMKnZNjBUZUmx18ywNoxZP
LxXxJ9yE2lqOX9T8LH7dUzoUBjl0/swxBde+ZMU1WNYvHeqxYj1tZhdw03hgus7n
EQDDs16y0aFKw1/eXxMZlJdxF/KJPwlVSJHmnW/WW5/r20DKrseP3GxUNL44pFtj
IGxWk46JgwUcHyldHQN2Ob5U634xEtZwCt0sjv8QEYbK/VImxddSLNjV6riPYsAM
UhkQ/ci9YfVZI7LnCH+8VkJwxBBrqI7CON2tCMnPj/TKMLbnZoiOspCjesJnDpxQ
k6INxylEYEgtDu+7nJdZdWYK13o8gG+WVhm/hsq3ywvhQb3tCV3oQnpwCiSf0Kd2
g85S29T08/pqzOtWTP0Idvepuk8uKikf0Ztg+jI8aFpIHB6c9vI96C3NuAwYdmTi
YABpgRZ3gG0S/e23ptIHcyh/GGVK5Hl1zvzN266NXdgdhFM8NUshCfN+PueLxtgx
Bewen7Q7P+JbnhV5y0F3mVZTi3P/IhYrWiyEn6tSDvyUoVmM3BgiRZwtPlq13fwv
sBkwsDzTSRSR3kd9CMAPYgy3idGzcupzs1ek930mkOnmSucRbkPy1Hvgh94y6ixz
fDxw1RQ9HTYtV157Dc9jGA/1ORbxT5ECKxrankrCUSfQXKy3BNIJJDQR/SYvmL+5
Wwdur/l7rVActjXUjoNOHxzRNIC8sEchIeatWgnlgtLmclDBlOeXnYdsms0edmr/
8Ssv+UAEx5xzsmX2W7436hcwdK/JnquaBq4M4B74lTBsQ+xzJGqQbl4lTQubYdqD
Cr04ZGoNmSEQIiEbashtiSaR2V1hymywnrCheuV6EX5/mZjDjkj+OEtfrGWcJnqb
IpuDlKhNpkbxdxFd5QS/Qb/p2r5Em//wD/xRR8yRlL92cANMqbBO8nDIB/uqtXi8
MqpCgMOK/yn2XZeUDare0diUX9ICRvD8U0tweS2T6BwioDonLgCTPlWRSTZSN1VW
b/9IlcVKSbJgICwgStNG13qVcX8YajCAWUIM6j41J4o32zYZT5Pg+LFEekz4Cl4l
Qxqf060v3xFHtUOWTLgzyYBVCh9EyXtVLJn7h0f4UwwMsxh4yaTB64x3f83fRyhe
xiU1w6bArHXkmYUjgndj52TBKtGa2YESmLsTNnxJhVohywumHzXF4SGhxrgDYa6a
5wESgAvAKVstyjDkHGArBHaQ0qKavF6mQXgiuEz/m+W7T3eQCP98udWk2exz2vfD
Q+yhGiz4kBguLHWAsZLcZ0txkvPOzDJ619zwckJCHmQhjYUHyfz7gc2hwjRFS5qC
Ojd/0wJILjuoL47A3+5D8AZb6Ctq4G9w7IrjV2PDqJ6i8O7r3DI2/0js+nFZ7Zph
xDb3svQDu75PRr1PmvwZ0yAmeBPDikAOpGZyB3NHXOBMQ+LqSbVKNb80jE24jIAi
9jFdkukUl528GF227rxOKuQREfchfTrNYxFva2EoTKZiCeMNDWoSLBo0MdlUa0dR
roaX9erhjoIkdV3p+cb0ezmBeXPHJSWggNAtWyxOu/qTvgs/WEKDycWgnm/oAUxw
czG08ngAP8BF04vNXkSa9AMClQoEk76iG+QIajTI55wrC5769hj8+O2PvA7+mZ2O
+d8VDwq5GFEluXqJycrfTD6/aU/wwUDNnFpeGkc83HrgL7XlxyGenp6hbfQLwmYC
zj0gJQIw+JqBw6Psr9Gpae6Ef5mYfLXZYWhMZagFFBoTN5ghe77pI1LhvVHUMVUi
0gBjUf8DoEimu4isPmoz1kiPvTJ9+0VwMcdqOVlLX1fcvIMeWe/WvyitLkvHaF5n
2yQ8rEEkl/cl7jP15ccEcbIgTGkXe+5/oK0pw1T3eLrtjGRb/XPEnIJ9SiqPjF8Y
ZAQGb4pHPqt/ukELs5hFHm5ioCCVUIr9uxVlEffsb0hakg5+8C8vS+lkpISOOvpe
qvvVLjVH8aOM9OLU++WjWpruz0mUfKzOIB88eO8OVyBx9rBI/3Sz/mWrbj7QEvKO
wmv5DpGmF7JiA3ZIDqXaK8YHHRVYGdczA+NjHKnL0HI/zBPbb31CjWvxmDHzszZt
+zucqEImdd/PAuis4EWmQxL/VvYHmpCk5BzdXQsVPzkSUbBPACBimk9iOobjc8/O
lhYVlSNcJoVRN31gbA+UrpZwELKmxW6E8/5DHvUp3WmficOW7obbIfzEOSOVBoTu
voaupoPJug6yK2tvH/WF3liy3OZ6EGhbDJBWHPAObDMv0HO7FRxXyNopPeLnhRqy
kBL0lv+5550XC9wrhjzzNhisEKRPZMONGiP7RjvRVk6x6Oi1bOSyc8JCMG3+eCmf
p7i0OnIHp4fLK/OxlsAC77Kmkc8Zfd4ylNo+sWWO6EnW5jcTePR9q09RGNCYSdvB
fKYqc2pf5XuQWgiYVt0fsXQtFjJk8P7E0/mhYgDPEHf6tcJDQKtofskv8puocsuG
4wOKgHPd0d94AXD442oq5ZMAbAwMZG16RgRBGy/7p73qgAM3JYLFbjJ39dogRrtN
QI+UWzSosx/O5JTkMia7PxNYYlS/Kubj0u7y5TutjQZp7STu7VXZU0oeh+/8yaDM
AcK4nn2q/ZkqV5G3IR8TpSUTonzKvZY9MPbvM1dIgLi6wRUda2TwFDUxnhZ/8LKM
7ZeRyKMYUjTKDrOnUExEQ8vHNJOBDO790Dxqy8259OPNid4kqbfurwPROrnwy4Q3
u5274hCeJPBM9jS9mKIChz2oxCfm9oadA2hRK1oGfVPuldjK3Cx7qun/g8hTANzK
HSn3NYON4HM8KWUMIgYkOGlbSmGwSYpzcGve6k82tFtBFyP7SaJL28WrTFxaPiEO
mSh2yjtxb9yTNT7RcIcvoiToX66/kvp+uVCqPw7jHu4HYWeO2+aSt54CVzsdHDSB
MdpE5O+2J+EOLoxXqnKnlb8rl33RIf1PqnVo7IPukLvrbyU7Oz7PIvo7mCcqkbu4
zzKUEcsMK5eEig+yak2yMZlrLqgCpNfMC+A5Gd8D/VaBolyaXXdnYYZ/GsdgG+ms
/ajcRH7GvDZgi9xcwTf2Gm/E1dv0yANn98gg6bAkFM9ptC2f3JV8rydIrqdNOVFF
dMxA9JznQUwGEoSbSywsTEg4906aZq+jaibXucsee+S8Ljv/NntgUyH43dE0bxS0
eCok0iv0Z0gIzzzLpoAQLIGsJQovCbn97xptdhPPI5uVMrgZOPOvPnWZhIUP6x/i
xRUynjFy7bjxz29nStz9+T+GWPnCdFd7aMMKH15geaoYQ2iFOYGaUkycGo/Ydv8t
UiqYveG59qeKuBlSgqMO+tCjwrpzvYwCoNxlz1jBGzAIqBBtQkRF6Mh07N+4fxhc
zDYULbN1WG7+A++nIdqgwK4MOQnB2Zmo4HswxZUMHkgMZL418YKasw1ECPlevM9V
pv3bmuvXj8+wIFSFAZ/60255+92LPpIO3yM3ct0ULYJurLQv+ryFEAtFdI23hH78
VvJ0chb7CVhSG6hN7IKnULfTrT3Cqzz24dROI1gQjCAkYWoc/6N7QppqDsY+OWmo
pe+AuqzXaDgi72y5kwitAHWF+72wQ8IMiezNTruZ2RTY+0ktX/OrMtmjEpbR7HFW
xKpeOFhuxFZRYcUiPKa1Uqfdbbcx5YyPFQtNkSKqDTmpgxjnNjLqOjaYXm8lR5ov
SLc/qIx4qN1iAlQ2c6lYSOekTPViu4jJKxTq1mlJ2L6tetalW6FTqCVzkDJDl3Xq
tIQMFMbvYF7OONCcINMPQic550/HRxzNqBj+ejEi1NY1SoMvhGDXfK4roKAR/qAY
UqaMe/d3blDCXPMXvZI1ksZ1RQQHzorJW8GmgK9CdbN4hQlMTM5C8s/YC7WZmKur
L1Fa6i5D3UTBdCDoQ2GAf21z0ujQvKJLNR43IA202yDrsEHVSQM4jZNYgl36Jss2
z1GeAh2g/+b6M1A0/VKEkUlB58Fh4JeqZq2ncXM3qzi++BRgllxW8Dm39NJNDYaS
yVWvwmMXtOf5KoSuJKy0ck/V1tkO0HhqgEXW0qRxSX7bcRfcjs3EYmDYmJAIOTo3
a8yx7JPmMFLDTqArd5MaNMSSm7W+ECaj6RrXoc7GMcnPq37arzKCbHhdekTlPRzi
wBMfkgnMKX327xC2iENYJGTG+Y9KaWjOxKY7fRZxKC5S72kYbW7rtgbtigmb6W6h
v/XZ+QlxLWEl0eZEmhPjtAWIBqdMQORMqAKag7DTHu3FSBBhqVbBJ8ld3S6kU5Kg
db9qIk1aZOD3w0ZPyPwtxSaFoBa96M21zLdv/0vwHnOz4WOIMvAE+rRxXF+PTXqz
qhYl8gYs+JW5jhm0/66HurA/wD/0sRkpOOKBlGCxbaZkGfDYOtb9my1Pr/AEBifg
6yjTujWZ8AVvBlBkOt+SWtXI4kG+D1mpp8b6BF1fag7CwxwRUdcdf/P0GyGo7keQ
3THjw0N7px6m7E2XmibtB3aQwDoFxwDmpJcfhu2GCTuxnzV6mMC44DaUQvs7qA6v
3hQhtJ1IOzYWtp+4MyAUfuVn2Ln7fhTgG46a7ZJZLg6sipyWWUKfFRViVUjYpEhX
ZPr3KlsVaR6jSbSw7gzkjcifIGkpoTIOzXBhFbD79yTEEdEQpyN/hgOJsv9ADLfI
mpJmIL38zSiHJQDF+WxnjDpSFiF8U1pM7fqAkCozfPlfCC7Hu/SGF91MaHdWGV8q
qR+Gbu8rP/qSX9quY570ySYF0GrDobs29xxnk/MepWlDi7y1R+zMkYfgGYdIkVXR
7tI37ys+M16FS1yUvA50Hd0yljVx9KG2FPjn7MbclZoFPjdbbPxPMUpv85CZg4vk
RIr/iCd5HzHClmWi272QLoGSX91tz+9m8o41+MYZEjD5Nx50RjS+DNmyrJdDSjuD
VlZ2njKb9IbnMXzlTMXqPTqqn5Dmejy27nZvI54rwhKU4e8Ngvyqha/LNxQftvLE
fB7UeAiVrwUaWN+jpaYY/5pmmMzkszMPrh7Bu1qA6TTqMRwD9AgsUYhuRnoGdW+A
SG0J8+QrsD/HMouPJfmU4LEqHsloDrIAhG7ODH7huMJ2c8X6+t+/DuDXssMVWnou
8e4qbqz8spx+LnoITx2+Fb9RmmCZIvCAQydU1mWqY6hx3bjY7ogDSVFu2gb5HZpy
7zM8P/f5RNSbrHQdFWMlEDEVs8++yyLt1+dh77zuZk4qOK36RnXXsHKoVXnWX/dm
50SvAGCJwbWT8O3QLF1zrH6TbyJTqG9+yANN7v4epFaqYQJETL2cEgf5r4eN/Lui
uTrn1mBlZUMRG1bSsMEiayAFJmukVEiFnfmEGTOJc7F/parHHOyMd7GAZF4uoPKs
0WWmrCRdE1uaQP2Gdm1jVrymcN9eQ7BmcCRgOVTST8voI8/6wQ160J95q136z70b
GfNnbXgDz3F1Ppiwq14LOIuW3lIseeQiQ7EgC/htCeBE/LApLdAm7Hj5XZ0eV+XN
EXTB65JxFYIY8gKEuJ3TzZTnV8UoktzdWM+lPImWv1RC4YUEyVmqHvJns6N8hU2r
Tlkw/Mh5zPJ8kXApMNc6itL9KzKkevklySMdG4ZI4SXBCFkXubeaZuoLQpfSTlAz
FqzGrraZy9zWzlz/XkX2fBZ38vC8uiIHzN/DaslpmSuWr13fbAyW8YoFYZpkSipx
mAOoGrEhCIFOmjUhSPtVPA1xsGp4F9zaUtOaPAl0b7m1izI2y1NvE4N/IZtl7igA
6LBBc4MpX9LBK57+h2H5kykPcWUNNH7wxz/7eVSq7bpQHohqgzMEVsBESYuxsRFR
NuXTFf0DMtTBOfE1NwOI+AhAg1ZwB21vxGM/pHwu5LaJ4FzmMdjeL1rR2jJdP4Fk
xeWHraLOBM71LxGQIHyCbG4rYyTAoMSwsaBb7mDknt5pFV3QdcFMsDHDFvtY/zDg
TH0Kc2c7Ep2SfB5oJe7mwj4TOlm5TX/9q6dXw8mYGOgDvVPlobyn1l62dMVCpsO7
H7E/IsZM7CpsmZCyz3/PMBx+r/BuMMNfNxYdy8IvfV/d5Dw4+slqay305mtACkIC
Rn9VtrNcrxVXP0F2hIKkhHrStRqnBrINWNTQOtaJzH2bIt9RQgv0Lxpcz/y2zJpD
Lx6jbr/wu4LrQN/GqPiI2Rzn9S7z/X1R5fDWzsx+yN64ep8rqIwPIFMPPVHXNrlP
SxTfISQ5AaKiXeelnO2oOIAF3sQFUztb/zsoSCWUYkN9CuTgWwzK7gWAXC1uYY+v
mfak4jJ9cjCOSYsJj4L8DxfAsa/uhvlkAyUVZAVJEbu7DJyiJft4SJEczb5Yedt+
4iHBNrbBPC1XNgn8axXufgNh2vcxR/y1O938gQtW25EIol02QE4DQOWsEtaEZkHD
Un5rR1qtBqIxHGVd3qIalWfVM1VpIZdvHNMgh5dxM141DlGV8SANepRpbTaE3FLs
PGbGEYPwITABSv6EWAxWUb3xzm4F3eF7jLgM8ZRAhQU3zHx6lry+MPnBoT2+JilH
T10nzXauRqhZFY5wf0KUFtZxL+VMAIhdoCsb35Un7t4YeN8l7H5XYUv5ZNuONrOh
ilbqbE1ePYDLgbJQrC42leyx6m+1rILwyoHPYdNmo/WZiQ2SMimG7pvzqQ1DnCrX
4PlsNSLSfF40GghUlvUa3v7YPbfGxXR3yaMW+T3oqudydtKijQxBc9uwss4M6LOI
Aduh+sTb+Iw8jAp1Gs5hFU3mgRBjr+kPIsjPvGlcw219kYq5E+mrLw68TOZNu+te
tXPqWxf1tBfTZVeN/p+TkcCMUGefXbnEnnBcbleYh6gfAJnrXgtyhjb2ozlGHM7C
mtGq9ntdNVPC3s3c2KJUSMzM9/Ghd7+zanupPqXeNw0+s/aJTB211jbRmzzxFR4W
HuTuimP1CxKzuXbP/qY3Mojit/TvSCdkr6MzzmFoFp23LsAbVKsOjdJu6WSs6G7G
2PwCpHlxNaGCzQSrDIK3Yb8kHF6IN/RRVnkQUHwS69xujlju73xnBkmICpULgP6T
wWBVR8FkjkdMaljCZK6+AQZWPEfMwBQL2ClZgiCej2IK2Y9fyNMbVlAro95RqeSq
7wiS8kcw+o0OdpWWLvQPhoLtsJlf28H6G+GRenNR/+6TsPzf9joWHqcL4VpI0VCI
dTUW/2Je50c1kre3d1KSKhdv8fbFNLzyEcu1M1zF/I8gUevTKg8uRUn7ts3IkVPg
sTVVJ40k24w9iNmfHb4/7uSSt7MDPYRLRyGhp/L+FCuKfoNlZYdb/4xRJmleMKxc
VmdvCZbgSq8BeQbtAf9ruPc/PkSbts4JHZ3o4bjfmEsDPVnZKuGMzIUm0SZQcRdP
TOx3l1T5Zvlnsh/B7ZrFlOQwmWcDB6isjANnqchXxg30OCJGcJI9hl9QZf4D3Uxq
+pnce8uOMVzC6e/yYbHr1sV7l4hLbfaezNLOdq6j6/ksylKM5nhvXsH38TsGPyIh
oPRwok77L6Drb6UHUetlXnv5AFZOZqbtFB0ZSAtO0WYtlgFnv3Ni4wTo91YuJ2u4
CNhsS8u/z9L2XM0lICtBIAGJqlYutF4GAOud0XGuiaMb6QTvEzD5gp6lYa68UTBl
54jjBLyHilx54V+H9T1s+j6VRvd4xz0HcLFiGAswltsYlOk/rkU32gVktZOPL32m
NszXuR5mkh2qZFs+BoEFpkdEukA/rTat8SvEujaV4nIFw1TZjsdL+coDa1Q+Napq
bzSxK3yfVEjoxdnvk2kIjbzGNtcfQTgxvA2FlWlvS1NR2Obg4MJFl7tqpbzdwYsh
Ynn3o/PksBxGPXIUN9L/yUs3jM7byyQe518QzsBugFgUw6JIoz5e0UkHE7AgHR70
BnbUhkl/pgz6VGH69MlKX6JN6BhZd/+oYPJVyKawnru0ZpG5cpxrIklcddhm4ydS
YzaPWKEya3+zRs2fKZ2cWp/+tEFsMXO3h7H2bjMX6Y96dypp/EKDiK6XUGeti7eV
JIR7nGeJiluwQKVcZVg0g+Co85CT7Zjlv3bpW0tZEbrAY0YHxwJnn/8zdsrIwbcS
JewH8/MXzAK5EhsajUYLxStZOYLJNE6QM8VTXStsx+TKNPFpbwgjVp4VVvluiLja
B6lpAiQRKZPdkhfIlHOFypkT2Ue6SpdmKB4IwpB34mfdtIC1N6HUhRII8ovpi2XV
hkEmCdt1L7q3uNE1FQywo4wfRm453xIkw9i4JOPFsBtNexbFlLOBV87RQohgY95N
948GEDA1/vRlWO+4iKHYm7swV3lDAjZ+tvKxMqMRKIZBhc9qVlDZUhTP2TrCtTu6
ImpdzHcyRP2tkF75U0YSmyP2mhY7c2wlqZM51F7e7mSeunnWdCfJCh83vXrgYv6g
j/J4fJZ5Y+iYrjihGl2r0lc25E8yqDVTaDU7zrFXHVH0JGSB3v+OcVHYDXmkOg4s
M9F42B7G234WmQXUVMbvg6gjL5Crt3lymezmfg3d4GMK5K9J7YnUQmoXDzrRiEAi
BzSHSPqia+PWXDaRWB6hlfU+LSLUWS3zJGwWR7nvsuTuP41S2Q5RoiUQMdcao00E
DLxoejtye668h2Dz8y2CjhNrenj10OjrGklKNBcXj2Nr2y7UC/kRz2yWqLZzVDB1
2hv5Q/EiLAlYu1dJqn10+jBH8wgdgNWik0I29d2PG1KWeXovb0qnw1X+vyO8a4cS
fRPp3Ao1klmXiDm3S5KX0+iGTuCtbOaJ60c6Z5QPEw98b0iv/jLajqEsUDszCEGJ
abkqxH0DTrH3YRmi94Ro9u5ShlJJA8lCYbh9L/dZ9HNQaeIaeYaLYu9hj+eDE6Fp
VNW20RJCVvTWxEZl/U+bv1IODcqgfiCHqqiDGOwZ9zB6RaaQUoCy4WdQFE4iBTFG
xu1YXG8yLOOoISzV/DCPoSyJ2ixGuw5rUwR7MOZJ4jiMF9vCbgwUYcONX+F3fFuz
vfYt6q5nKpm1nMsE/F/xhU5iXTpryfYq6+Yi2bPS7uHmeqBYxpGeYzboQl4HlajC
J7YL0QQDM5WwZlhhML+RvhQDtQO0MHtozinTU5i3OzHdSi2dsW5mgD6wp7yNp97Y
9RQT4DH2uWLkcJYMJcBEiE45XcFi+czhCfzy8m4dqwR+zPpkvvOX0pROSZ9h9140
370tHUnzx304aTi2OIuSW8NwkK2laAk+zGmTg9NU9cwc1dwrwjfIlCwELIIvKMPO
1wuKuZwkMewtLEvNwm067d/1i/fpja8m0N9OwKLMeQwpgjb5wa8oCr2hdB26YvCg
4ESGo7iTRfglpRCbM7SGMjYioP2jguWRIWH+UpSQ0igOhUUcr4tJnISbLXJVM630
SLNccFCEFtxR4ojk3WpbhwHz4b5RfbF7OAjdJrdXVxZNLXQ9Tv8ma9yQG0qEc3zk
kNUY2bHsKAvYInXMwNtDxS84HvL8w7lBk37XTxcw7p9to62NXLjimqgIMokOPm2w
0SDou+KK5EPQdfXJHgJAZJt7PIz9BLSAW58b1euPlxpjeBRQcKyA/1Goh2mS/ss9
94KpTK7U97rcbXKtlg7xiFR+Tt5pHo0bZsfA8R/YxnJ8DdyV0Xe4Gtm/KC4l2gV6
KBiAZpBeFXKA46DSHx6Yyn0D1TefaPalb5ZpxvdkYRqiM7E08RWtU+LBzwCqC2HD
pY4km+JcYfk3wHnu2QaokEUZH5SGSuKJEcPeLyc3PzcXzTNaF/jHG5JHxmgcBpHJ
LcvhXp4Qw3RVyF8wMJ7lGFT1cmFqJsa2IPKZKSNKbStDSuqwbn7s1r5qeQ7K9Blx
G1B0s/qgrQbgx/5Oa8zktT+ZG5uHFM9oGwIUp0jmUNolWX1qClFuiFCIOWTN9Wo6
/dto23LVEPHlGYslDjfvEf+GjsUwLFAJ12ZtsH5y6vGRBYJ1Vg9DbTQmGOwN/xAs
g9VnvrJdUM7V+lgNFFr41XVeS+H+O2dteCGvxZWFsrY/xfdF1XItzxXKg1zdhuJW
qrN415k46BoiFUCcPncfGD7xCpsigUoQAp9d1RO1cFIaSHu/IMwaSWg0jacl4PmV
f0eCDpDJzIwbXjkDf/++4xS3wulXn5w8irpY7uComBKG3stVFDKnic5+azSLl/aV
MwmRzQTmJWM6nuFPHwTqMGBmpVkIplOnYCrj6MvLO5CHXEys9LnR2knejcI5P+Jt
CnMZzo035aFCN3a1VhssEGoE7OTMoeaGdFzBrDRrUO33yQhWHSGGjyMsenUA0qMg
MvUSCItp4VU/D4ipavMHPOk1WluEBbQHMoVCAMC3PyranN3/GNWiAeJD7AGTZOJt
QTdv/6sNpqp8eZs43myGROb4ob0dc4MtjsEfP6nl/S5aje9g+/5aWJ/G7BBrraqf
7v6POyIZtH+kDi8FR+AMhK+liXPfBc+BT0k++faqSxx0574ZwYKmMahUQydfBdVA
eyVu0Rp9xAHY5HmGuA5HT66vrmmIDV+BUqUXwqxzrXBrU239ou0Dm8YA9FOtT1jp
esLKsY9ukpjJi8/Z6YRGbLT0aCZYu2PKsAWr3ZNPEl6LNV/iNuAwlia7wO2IKSRY
lfT1GBQQ31KbunB7CtP1eoE/kCd3L8QDOKaLa8HpzFOjopg2J5EpPuQv+5D0SGxT
wp5LdjMpUmK8VIRTrjkNGbwt7d2/APBdg4gXRONLSY9aQmzQzkXvuakiUZ0Bw7s/
Wi4UEyDGfKx95cz0fhlU9bkK/POptMO0avRFL+VAjuDJIaG+LQzJWhCtFt7BBWVS
av12m90JLp36vgYCcsaHb+gLeT0eWemepgf2AqQ6C3dlCi+1vTb5NaCIAIahjlHI
+eROdYX1wgrZSzUuWbA28pJCrAW5tAu3VhnU/SCK372R4hmJSz6K24R59jSUITEb
3rMBYRqWOcoxw+C7PxTr+tYcT6JFFFO3Gu7pprw3fvhMN0kEGfpThHRiA8Of0cSb
wfUCMXj0CrcdSYde1PRzYAVxEkw9m8ahjJ9dunQEBsIkRJvBzdTjIKuVBSSHr53I
S0dPySnr6aILO0YBYC7uxrAhyL5kiZpyUxoZ4cfHzeGs5r7O5wxgVRPaBm35Eyga
wj3MjI+MtdzkuPs7oPoHJbyRHu3u2kandndDR5NmqIgw+b9BFoHe5sFC2QA/chDT
uzrzBMCWGlA6QJO9RlHl2HXgA+h5COqQna8PYLAbtlvRJSa8rPI7NxaM7o6jWjfP
ylRiXCu5LW0s7nfOdaNJG6FgqfD0IbgpZ+N930kcRXQuLtdQjjsTfSFjj1jNQaxJ
3rJrH+vOirn97ohOdkqfJCAgSJtyL+QXVYBLnMhN0NAXTk5GMlB3VtJ/ujaew+Ci
ds5cILFy3FqiCUaHpHEoymRwh+omXqtGpydQYg8jtnxQQh16QaDfzCvFAcUcuJG5
IM/XEj2CcVlhSpjCBw/wCLWZCR8J3ZgNNL/RY+3bymgMozVAy64st71J45TyXzpL
2zGGDTZ5RcOHNRbmqBeTqnBZ4TDLAt+D3USFuTu98270w1pw0EcVuBgYf0S5Shp2
6VRxaP39R2Z2rAOjuoCj6hi9rEGaD79ymwq97u6nQ13T0cF6Q9R+AvYcb3TUHNqN
uV5E0AP/WiMbEypm/JeVYVrgapjaZi9+PHNRowKdZaZV6VEsAblTB5VfH11dXK0U
z7kPbkuMdSvVqg90V1na5veo4o5PyUx2RHiW5I/jnMb4qWDcppT0y1hpRh8KQ+lI
vJbnOF6Wf/+stj73AMsvIue6hSGJvwNYqEAr28l+E0AoqPLQ4f/35t/CYaMHUwYE
/wVyOyCtrEUTePWQlKemHjBrZdYA77W4yeOoFJ+BWO7A1EIBO0NuCQwXGAffUF7z
hOEYm6ED8K+ZxDSey6tOcjF46e49iXj3arOtNefxLQtMEM46/HoQ9xy8Z6HqNNnZ
frZVg7OEqjOG2q0qfH4EchIyavYmTcn1TXdPuHzfTQJXGOzCGRU1iN9XgMluGrB1
5XNK3VusC8jwIKY3J2OKDN7kUXB7aNY2oN8lKZ+Q+0UKIGsBu+yk+GSZC01cXyM1
vfKUU8Mf3IdzrTKBTf+ABcGKRiICiqSC2k8cGTxbIqhtPfje+Wx7LOnjU+w9H2wl
wKeVrs/amKrR9ej+OVzoIRnPjIRBTrOyGGrX8tPFTJBoHyw3Wmgym6f6i69+fR8O
ZgBK/nYkN7fORi5DJ6kTGtx0RXlt+uUsKVO5e40UQMBPcVJvqm+iV92FxCZBdQBt
pv8z0EerQZ0FvkOMWTuXVj7vGk45Avk1Hnz8Bh65M6YF4Qdgt/MDmttSKfjEikIV
bXhY+jOEsU1SqtA7TsewRnhoNuEEiK4xaY42SuiY33cHFP4k5fPy7g+PzAPXkBvf
K5ln754TCf4K8Q+D2xPD41e2ULDi2anpgNIjZeCDlRVUcPhRGmaacLJ3MEEWyfVh
Y5XW6XoOEc9FxuRA6DcKoDQXfMtGhKMUDasxe/tZo/1CO9Klf+yeHbPK1JHa/iC2
h1dnB+EfSHrZSXr09/7oi2SCjLOw2JyWqZ1wZ1wDDRRAo4lsF0wkukryzx6UlzCJ
syJTDCYPnnf6B2slBNnRc0tRA6Bd2m1Fh9bMFFSjzjMcpjQFiv1BtLvRanI4FMTM
2ehoQ0r8PBgVhznkfxvd+1YullwFH9cTxbC0vqWTl2NXXsckoyWFgNKDHqk1srQa
HA9OLCnm0FgD0aQRP/WpzJyEehwWeCMQk8UG3sMI+ZsShudQ6BxAb6LOkX7gOVcQ
6E854LJb1hO8eq3AbojrLVM8ngp2ltZbrX4hk6CeSO7gyosZGxi4r3hmtOlcHpuN
Upy0akys8h1E2rSRJjV3d+iHsQGmS7xZPBFjbNvENDm1bKSYmIH0gIeHVFRJth/W
8evG2OEkaO+mYKergc5UGbGRq4rYXxtpAL00U5eqEibhnUVeNgYg9ptduo8xaHNb
7ZYiEfafi4pnSq7IVfSPI7YdTZKt7BzIOjFk8ay1JCoMy/I+JbcvwqwIFaQKcEuo
1xDCKKg5mxcG7WPGF2IOmye+8ylfAuBF6nTrkoNq9dbav1BGwPsx7r3D/v2RkC2C
CKqTQCOqaA7cy1VhV8VGWWOmC5csBI+ZQnvgBE8WEYVW9RVeEG7LpShPV9W61tPT
QEUERHkRje5x8tz7maVhBkABiHERp3K9yere5bD9Bdyy/NpfecRrpMa67tGXmnfV
jeFrmmUBnGmyJiVtNpPeV0Ued8H/eNPohJCKJGOtGdN5CPQ6TCGohWDgzhTw+9Ec
Z8ZXVYN0OOBBZiaekEWcROq0/ffEr4S0bSd0wrJq14Whb2TFtct+hgJpO2UC7k6M
54iOiTsl2lyGxd4OPr/sFKe/qzJXYdJc0MGvJX57gmh2sSGHQ2/6Jpo/lST05PyM
BRxqJkidW5j+4+0jPMh07dkLv09r1PKWJCuoETV7740BkJom6wesPCgQA0JHxUpI
OsHhZsgOqPeq0H8Sq8jDDMTO223VZTbPbn5dE4op11r6iMdiWheRJcxG0ZF03G+7
ydm104D+ZDTtEG3Jcg+1vFmXKu+YKbAKZ2M4pqOZLlpLcNP9Ra5bnsrZt8mwu9lI
jrTxRjvhjqjaDm723eqXch+0zPvJ1T58k49ywYECeHDGwWtyC0nmylCGgXqoAUJj
kSAR70hO7LrxwwoShqA8CK07BQ5m1bJ796m7juTqboTIuZCf2LedM7ufttnI39En
ZS3Gss51Hzk6SLKVaZ1WqNUrr0NZCethcuTiay68NSSFeJn4VLKu8J93/msGyAJe
D0UI0TmjiPzEqC+ZuOWr62RD84EDrTrH8ebXW7ZyUwuPvvH2HW0OdI9f6lA5XaWN
7+ExUMOy/4vRthIyUrV2G3BVBUxJar7goIkiGO9/ZCLQnQlBKM4bWwJ93ZPG9UW0
U9P1yryR30fSsTfly0gNRRVyKbidVtaQ0jeQnKSXM72pV2wUtG4J88+ZN2m9YgFf
PYRpd9bKFUU56pkDG5s2Gi1wSw6jpJiQj1RtOgJPyTRKem+a6F21r4aloV0nIwYH
tP2xAuCC3B6pXAaDrpxU8RJzk/oKJMbk3qjbB+zByC+HkiyNEq77q5KwhR5qipUS
sRzhKFRoxHQEvQDpkNOqh7rqHqkM/qCTXP7aMuN/rQjZAGr8uPj0MqL5bkoFoF8Y
I4tJvShKIIK3ZLCgosVFk3qR4Kj/71yojKEdRsCQJ8ogzFz9gm4TGfebhvdlkOhH
yTEvvws765yaj8ErTo0jwoamBeIsfRhkz92Q9NuTP1eiHNZndsocTwYSOTm5UoUq
zjWDc7oG8xVvlcKDwaDzVxk9eX1S5em7ZJ0KO9btUU43AkJad7O0QF39NlbPiK3q
0CG/C/QVvGKz9wTeGeXYMmmkx5R46K6sU15riv2mpf0ki5+Glid92l0EUXIaN+9x
vvnwcnaq/JIByC5S3E2Fwoy3iD9Ily1qqUDDDxgSyWxR3+cvtIkeHxjp8RKdxkaR
CSAq6Mx8QlIC1BkkEY2jdfKJFtvv7YHUyN4ntz+bKMs4iyerbWe7+jj0skGL2JU4
ZAt9Ez1VowCb9LFpllhfi4WUW8HICJm1ss/sVhBf6/9zk7xXR+Rn/gDDn5sRMcsf
2hdgdJClvWG5jGlBnLHOn9K9HGX1JIXnTU87ft5cdubCMIlPmSpPvjCYuXAlvBAT
evS9p3PNJLROmb4tflGV4Ps14SXqGumNSiwbjJuBMlV6RMVm9RRb9rkkTSXM/Jp1
ITG6v+E7KeGU8nhJ+5yS2ltoenZUYlyIkoxDeNBjHdBOUdOpeoqMdHT26dAttDMx
XmIFSff7ciCBYNBsVlSZduNjph9apufsBvt34LqMY0CWbuabuVUIcJWOuxBSAx1z
ChpAQ/YA6zQo6Y/1cdG3n650VXb6n/FDz+eRUTce2SLD+zVkLrbGTtn8dBgp8xyf
4juMjPJeCZCfPMZrPkMGZILiHa0Y6M2JCW8V9gBDQlI/AVmFwJHdIAZmW4EljAlo
6iLkNMZJqyJq3xhyS2aRzJoL/5hUNqXW3Rq6t+tC9OwHQ4WHVCtZvkfvDU22gkr3
igU5LmT9M5C8BqwvjwlqSug6sIUIHGnA/+TDPSDr4ZVxRncl5XPFR2gKNM4lECsl
/57j48Pl7CsTb/undyYzkUFJV2qctFg2hFEmKbF1KJuGGFcNZn30jAFUbnzVWxEl
7F5HKaX8/DRZmu6FRxxPfHgaVt+k3pgxi0Ot5QqmvR0PAmvgLJDlAG7GN7NvytXg
LMyWYOInGoGtVM/NmCSVzTlcY+tI6SaOmQMCmzNdnP45kfePSnuWXvt+8+Qkjut8
sznah6s61m/Wu2oDkQeiH8370Ydve7SRBYdRz7+1Wojwk2LrPd9qHn8d8nNL+lU6
F5xbnoP5uyALRrHszqAcdL7irR+0nrhZ3XA1hWPNxk6swnAzuKvvPgOQGTNmitdQ
XGtvxDWiZAEHjEuaZ8TlUtYvPm+jHiVP9IvPHK8DjuCyzjsYzd22j4xw/A+sQUP1
6fojuIdylJeIY2N3LZsH3xoi/7Gb5XZRfmavo9krxkNqsJbCuKTUxCw0At3LkwiP
bAbzrI2FTxRmKizFLIZ++Pmp95cVpXa/3AOJSMD3oTDGZlFmcmBhhfd6hx+WT06H
euEP8nCeDDkXOyDBKdMseeDONissHSbfV5Ci3GnUp2a+XParUTA6eNjg/xWj9KF9
hEVJpkqpAGRMrW/BEwMYcx5Lja75qCnty/hoSpQC24eEilHiBkbkiJib2HpNi0Ib
qrgznPdQxCtMC8cBFf3FUlUsAwLid9qXcpZyfvcEzsaJKh7Q1Fp8IMQkLgZeUGlF
YmlMSkGhGlz580DCbrDvOmKZLH4b+9NrpCfPa0sK6ls1t+Ecgi67htJ3Z5xaFCDH
1tYUicBXkAI1d/T7SztwFAw5+VfynSuJQXeg5Id1NbStvmBbgHkXbgVJv48mwRqU
j10eANg0sVmmO0/U7WpLx2BjgLPEHmnzXnWHMcWkWht10CdwgPufoesmezvAgRZm
c02Yhc2bBRlhD8JfmADf2ir6BpHPf3BWi9fL5VacgUaQpOdsilnwm9dAI4hhiFrB
PMA1ZbbFv5fKy6ZBWrltQzkXjDIh/99mQiBkMWPQYf0Kh33zJ4WiUyXFJvvZvygr
vEcGpJBGyRUBANooIUN02hWclYKsAAZSYn0pmHAa9JjvdpeYNA2VahFLfg2oeETU
HFN7aL/uWsCpnmfAwkhIvOMU2wAnk8eollvOsr3NS5MCJrIfaaFe+iGFWZEh9JRh
PCQt5xtTzW3jaheKOUwYJTZPYCuErcpENUwbSuXCCX0pvBqmIAY0VVc2qLeGdFPb
8t7Xj4+lT9DoIz0lx8awBnk2RytNvWNFT6OSsKpvobVttplp1ogVIrQ2Ic4bhh5P
kWlyvQLdayq8wxz8fV2IF26Lr79nL9GE77pYaRLIJlEo16BZOKTQtSeLXDR2qnTx
Tt4esJAbv0/yDxKoGNA/A24TOuT0FkSwnyXFffzMoVofWlmyP5EuGrPLO+n2G9Q3
81XRwFxZS6O6uPRn4qX6lJCzj/O3DwFxoojU0+IeihRpMQh//ItT71pBKAm59hqJ
jaAZudyAGiEjvwQZklKT3fWarQpkVQllEcnoGyIMF/LM14KOfU/xqWuuKG8d8qfa
LWxtX4LKiN2j7YDWofU8qmMsGkBI5AI6GTh/1NnhYsoBpFWLVs9MLfVf/AU4aRlu
A2tX//p8Y5+rast4pDwCbt0xazwJWy8R0SgkXzq1ZUSElSA3gQLOS9TNAAOwsN/7
SjLkMzRXYWy9FD3hek1LwkQ+csyaEWsxcImYHLlk0jrWOulx6qZvqYNqG2aO9rzA
UTxhueuhTUU5ko2KQak9AzTQJxbhqcTwVMeYbbSHuGthhib09vNWq3CyUDNKGPoA
d5GQzA91Ur7NB/YjrNPmUMmUCm6NkP9kt2LwfwY26QpqIKJC4YP8TrVTLSOaJuIB
qXIYh7TDdW7bPonGycH+6dzVWUzavf9f0d6FiVkkmvlWpFk8jS7DfEmL9+oQHrJL
ONRNgTpguIH57eczHVO67rL7azonIZVGpeRVHRb1xBXkm8+pZPaU8+iVaBodo90N
wo6OHouwfdCxTttwNQIjx4JJiIfQreFH2EAwC8Iem6uFenVX9VhzNUlalHPuV/bX
tca4e80ft4idYH3CwoqGhEZxYtpGzX/vLK07s2x1hvH4Bsn/EinTLv8/WVVcYdaP
kEItT8TuM1rlo1v4PfVnKP+SqDQSGgf6kQJncZDnEW2Vo2WwAz+0WrPXXBCnmMHY
DaDuIXDgE0JQN4zZWhwKsV8+fp7RFEH+KbcugkkziioFgPEjyr22AMHVUcEbchsx
dLRCUekLZcNc494Isc+btg6dVSu01TImcKx/oUEUBFapdq5RyzgjFKLbnZqew3mm
F54JW6Jv+TsApH2PJij8pYU8UOyrI61DTWdei9z0+57pEfjqVGAtWwCNYHHiMnXm
X/nSdWuY7jtn1XpLfXrqVOYtBR/A0sBXtiBu0j6sijtriZYJCUsvB46RqavjFOcp
Px2JsLx5xUpJOOSqS6DkssmP0Fm8uZX9pTJ/8DwLw9rhKYD5M3juE5Q3CsrhLS7I
xdxM+YNhJOuG0i/b3T+g684xhlF0eyP2438BZCRiiCS6YYD35G9wPJdNUrwJpJHZ
YP3qOvqAY/BFdwk4okVEylXJrN4kuHY+TYSQ3lGm+t0JnBQADnUMZpsbjmlxIlSU
8T/ECd3j/TjlRQjT/SmHv3fgaSqRDhxah3N+/hVKvg5F1wA5dkqELgsyYXiD1G77
P4iR97kv3hgD5wq9PQvBOyq3YyAyimX5gt9NtOK0Je6jSG7deh/cFBEENKIalmVB
RL0WFDR15FLq3KAQJYKL2nZu3Y7XwhpX6mj5zyqT9nS6tDHU4u5ioi4/nB1y7VmF
ABitZ0a2UkTYQlM5tvP0BulAZWz2XUjmrAwxB/QmU+Mdki0o2nIl/H5hWXdXOAxf
701RwQ1xOI77pftod5lK8m6SDd8ufOa6RGwPp0g4SJiI9zEYXY7axQXwVRBdJVNH
9hxVeF/pb05Rgq+RE8hpxowDe82XbwEixWJNFdcz1brK7d4oYOeHX5btexo57S3/
w91QKJh92Btx2V99ZymNVuJyt3Idhts+6mrLML6mZQEJP4LEgqPi3YfWSY4DTDfg
MlKyvk/6DOPTXRP4zKectG76VB3DzyQmDoE+HdTqys4UE86bQJ9YZlG2ob3NckGi
zuYcYymg2S57Ri6qt5ca/CispkGhdpYDgiIEpOTjf9njUKZoJeiaXvF+qsZdLcm0
ilWWUJgi5VeWPQjXSqfCfBUrVAz0LawCpL5DdDMoz0dGx2S9uO8dg8i3GR7XKvBn
EHpXTk98cewyDFumPTNwlPjjxfJN699ql9cOC8z5OQ5EvDRXG6sGa0TnPvutbJ85
yMCIEmmydpxYqa4w3n2M5Aw1d+Gkrk2HV1OFCfqePgPJLHYCCeQp2LJhbrhFHPoP
NtCP2VwTpez/qdVMQCVvRVWW6/eOgJDexQIREVXZWI+U4WflsEFHOkiUqq4iz3IK
EDSNe8OOrRiQQiLuPUd0Gs9UMXddm3nNVz2XAFp4gGalQIyt6rXik+Ab4R/Ifs7C
L+kcLoz980h/4oJT5FIyR9LfCD7Zp0+nJIwgoyBL1SObpanI7jzgcZMo5HzWQ5hI
Fn1E+jrH/SpgoSjCeeKd8ah8/lL5RxQI3bmDKGKOMyuCwLqhl7hH27tt7bnx0kQk
Z9nqyB30mDe4TUhpJshlRmOGmCJnoXdwKocQolJ/Rxc+83qPGZZwVP+DuVoNvmLJ
HmkwMMeSrBXqwh3SLPw9ykyxuMvbqg+7ulptYGbW9lFig0utPu2NgzdD1wP1b6PU
QBko4vlMAy8LWfwyfmuz6c8goF7DO7SNuA5xSoYanUznRjaIU3Ib0i5FJFF107WR
U70roEXcTVJIMl6U66Totf9Dj+FeXgoNB5JqVQk9A6J4ph6YhCOcXQXR1d5jqqJJ
i+FYDOQ+JTPUdz+RKUJCzK9VvE2i3Iy2VtfbViuaEo1W64hcfSF976g1n/GvROUf
W3JObSgeZoHRBW4Xrgffi2tKjQ2aS0gCSpHmeo3lzKj+XR7nPRL+1MgzZxNKtkI5
TTZLzbYQ2v3Lmo/vbwgWX53uBRB4DgLiIy4UB74cIbOlUSJpZgwMWLhLMkKUMlUc
18q9XsFjK3kA16LjQ6N7R858OuUJmkZlNw01us7Hy7yFReT4ij+s7MFDdvoNiIAI
MiROsfsNvNPUDwPwo1UzyjABpOXhYLJUTzxdEeElWQOeqSsaNkSvJke4yljQDdm2
g2+w9R2yt6YFMGwQlEl/hE7D+NVyopNQbF746aFe2v+QDifA7Of6mPVhO7iNYszu
pZSaiY1lAjTioHn4mQuKgGBixPr9q1hba4n0+AUUDdFdvCvbd3QczCKo2CR1R1qH
2LBebgT3EYs3ZbLRCxja0GF45rbSCoEXhl5VW5Awx4xkdQi5Qs7kKkPbqJHOHlBg
zpY+ar3UIGxEtN9rMvGZzOFyqVjEEXLkcWRZCQSuWvbVQQDtssdDOMZjRh6wra3q
ij3HwQ0NOiy5B6AMNMXNcfi6wctEmbl+gNXYG8bUNT7mICavrX0uHMXx3tSyiNfX
8ZWxIzqGnF15K6LBOkZ+tJlztghfWlFnUPN+n5JudJBHTrSeoEv5vX71JQlJKaS2
KaUrhAbK1nwXfoRekFTEVJ86M47l96Fx0XXid0MKiCJnatGqI6eSCxGxOyiFfa/L
R4KQVJXjRCJn+1Yk4biz+43GDSmH/avz9s3XlzvWz/gT/pFn3zl42rQMeF1dqTRw
7ieZ2SSX1wiopRP1Ly/Q9UPyLvivtTbDHS4Clovw9ofYBzrbchzKJvcXnkbT99zs
oqZZKIVPWxOSkOAJriLUmm27KXFZ4+sNVucZb+muR6bmciFm86+r5ExTEQyM26zp
FFTxa/TN7l8rIBDbfgvdfg8yAX8ph5ASWSC490s7OJ0m4nsNF4LZTQ4h0QmHQe4J
ANB2+uxPONqN05fN/5V8xTekctMjc8SQPA+RNcpdRAZoxHoG6pfsYqiNeb7JkcBL
LZzISpzfbsaj5DgsQVenYQJJHzXBMDoF3p4JWFVR85aLPFGGnbRfNfmmnasn8WHN
pw5tNQFEi7Q2L8L3/QlywwhVWztMV6481erMobfof5k8nWEaGmzomNB2dsd7G1kN
Gk1PZfv7J6DJgE0YE6U/aKhQ1v++tx5u6g0+kFoWbnTmkb1I6fDwjL5kNP0ADnvp
kMt0J5CkFHALOubO95b5PZ8K4+dIINZKmtU8Mki8nPIYa+XOeNAIDJq+b2wonH3q
q9bSgGBWjSQIelm/UWvyrXOPx96oFT1xWVQTISyXRgATyidc/O9mKXcmUj9LcHvC
Vbrchea8+kNQbdBr1ZKXWLt+e9FtsRfENFWL7RJShc4JsKv+FH4e9Igi47LWNrXk
ykJoStz7ewr1BTIOF+GMON7h85Cq+0b9dV3GZsddDt+SEqrOstaqtVfY+cnsSTis
xYLztQGf2uSuYt+bAaIuqpeIi9LmxHf6gAM8e8SH5Ry1+nqcATDcaFzF48VfleId
j/O4uvTRFENYMmChJiv84coc4P4yosKsm+HkntSbBMzZFC+w/kjT3i1vC43UyjFk
HvffRb/AcHidWsb25ab33ZE5UB1tB71+hw1UNyO6yHB1L7+4CmZYilqHKVWZecSA
HVwG7Fd335zxeULMhDDZ5i/51zUQd6La9zyNqH3RlpahtEiLTr7clcYkO32R+nyt
6/kX+z0sntMCii1MUDwBY5DK8roQng9Eekd23tnhL2haqIY4ry5r5ytQasEBoovL
KHozzEGINdl8wn7LvA3V69morIter6s1BfqTY85CXFWwf/Vsdzr/TlAt3Gn3V46o
2wV4LOwmZ7iVOEZbjZrqwXKzVpVEvodCwzP/4mPHA6MyyAVhGH9LvhpCMtqiFZi5
10FVRhr+LFidSx2/3IYY1JLOMQ96fOZpJCEyGGekIixnUkFbF0sdve7IN9A5HFy8
CnK5tGDbDpOhHPtTpiOTvEen3fZRCMS4svMW1f8OuCz+R33TMyWJellyXpxp36lB
f0IU5HVA+J2X/kFHoMfsSYu0H3ryVVLe49UYUm/Rj5V+DWUvy5m4BiPUp3VhhzNJ
oavnPAQDZAECWIDrLWAoVyPCjM8q12AJt+VhuA2iihAbxzFuYajHdXWH/WU6E7ow
5WSq+mjTefZPOFEE0GYAEhuGQq+EqKVQ8rGOHwSG3nEO33sJncu6QL+GHqyFUfPP
ZJrg/FtxiWldmyGReY9dk/Xa98cdYzXXi2/pRiEnMv+SPWVSea8426QjfVu+velP
c1bnWYuiOxe7hqvbwyAsndj5WlYTPTPt5CGH64FkX5Zyj19SiiPLBrC5pFAZFfKd
GtuHEaDKiXCQqVD30JJ0ow+c+ldfgmXkWaLQI0OoGuCzJsF6BMsb1vtWBuV6791F
ra/zMp4wjEbm+iFl9gSunHsIxiXSypOVpaQEi4e3+MAm6Hk8gWRTL8/rpWb4T5+e
/CKUmUX+/nIpymnkBVj8RQzcdOJoz+fPsxRGcnJtnPxHLmJ8Pmb+JxJ1fJ4SRROu
Ik7oRTtv7YMZgmfgmQOm4StITd9fW8uAjnCqiGIhS39XY95YW323NZKgGw4Y/s/j
26FalbOcDMZNJigmXlfnP6xUPZgRb7xGseVeC+cnTfijnzuc2LQFqkfuuEeX+8+M
qFQmWSOZSfVn4mX1JjUln7JS1ywGLk3Lo2FRRbtZHjkP0BWI1jhQs9U2eYia1D0F
tczx80msgWoGojf7NPKsCb4PHPVK8ONbPF22FNcmXstcallnLssSdp+T2wQER8h3
HxvyjWjshIO6MuayM+as+u1JiElXBf5+o7Bb3UbSgglDy76fXqbg1rWo3Jdrhwbz
NQAeabXgN3h9XBrv52LIrM+TdnV63r9CK1a6ED2y8Z4f9kw8tA0Ren1ftCJUB1sQ
e+VIYzUehQJZtX95F7IKkLCKBU3zVVgeLqnfJrCYR5oYqHkolRBMMGgdGhc/GzrM
lIeglwf2jHpIXnsIB2onRlxHUwFpga+fMNDTvUGQ/qvh5zQrrVl7hnLxG0LBU+a2
VTBvAjhrKbGzpAretxAA6FgpVOxhlek5GS9oFWwxdZUPGSKHciW+Pkf83r+RbG8g
g10CBULDx0sVmWA5h/4l6xISL9ups29jdA5K8xbExlrX0M7q8hnshWK+ntWK2rxQ
wV+fDUP+QiQP6FJOXaebJdZVPTVhrx7vBQVh9g1/U4FFfyc5I1imboFdWaujwTZl
J+FG4GkBH768PKbbvbhLaRYUhJYDWwmkZrhopb3eoqcuPSQHFEmW5zApw2I1Pugx
8+i7nhs6NZa7yDNBlekDfqamGtb2//NVR6kxaX6vSUo+2Awr3XEKHGZ1jPBvWwu3
8wbcGmpsLSSwvfkT76OrTk714EX2Im/tIljZVuPbKGwvlyEZFcqlitU7IYJdL62w
u+AqrQqBoRPSJ4AMDTbxRezrghAcMBWasZwiiwlVzN9fOeibjIulnDquwhfYWqVL
GOWctQiPXRql1iwHdbPzs8RI4S3r/wfczbULOqwkB0ZEyJlqq+B6ylQsTwQ5fq+w
J/LpJOC15oUMaL4vpiqY7coqdufkieTp8t58EzEhJqFsuKiWmQvES9zdXKrKf1eC
MgWq9ArSuZkE9gLT0/ufyGik+u3Q3QI6GVOkXIz46QrF1268xFcUIv/z6GTolP0B
HHXTiyHu3vRF36iCpsbfx4FZ4ftSC4TfxW3Yl28IowUHgOnY/DXifQ7UntIrKYdg
2GpiEkvPJV90qZ+/WYLSBgl8pf96upWgBB5/jFHVcJcDbss67/SMYwNDA5ei0Ky2
oJ6yx9wtAM5N23riuXhWJu+ogySVaAObylmjqbyp9SPIYsKSojjTA3HF0uQjHfLU
/pzTK6wrAUjkPaGlim98ezLmqwpge0JJAmgKFfQNERxdax25N3IKNd01Fjc0Bvf7
6A9nAr4tJ4io8zBsrZAPZcdquLwrbEN0+w7U2+GwIRq6QBKaxH+cj3zm9R+jtqCv
Q8vHs3qm8K8z/gmvJWW8fRmHGiwCRQ6txl3mb0oPkzFo/Wu7My6SU8eo7C6BRIan
Q2ffEEZfbmUmS3M1zitqvX+Cecod/I0OQVKTtt5OB5RwdozyBj9frRlXVGuRq/jf
kUEsuycr/FG1coPjnGu9Lq733JWsrIHCdaNWpgChpdiQD3yacAdUQDnJXKtNFTR0
Ca6sG/EbCfNaPHoQW3Oarq2KR3IbCrTwDlJ7/WNVKrOUN3qMrf7JJJjN7IBcRxHn
k5OGFBfETsbJI/Y74g8eGhPqhefpVx3v+CKZTKwazCTiTEc6rpRn2W9U5PSCVGNE
Ynz1YuKRX4yIUVdSL8CMsqDyH53KihCZZ/yWhCBeIo6BrLy/jl9cTlVqKh5KA+nC
8AXCik3ereNt8ZIPIcMqhauXkSorcerLd0kx+Vn0RicnLOdh3YC7BNLbNBcHj0wS
gzeq8Rcjw99CTmPkBnFDkA6YmeBiexMdOf5MXoPg/9zPhe9oGlnteJXgEQpcT55V
3Mo9HPftyr7rk85xqzoVbydCoTPhGi1f9FdwWILDZST6GMQJ8B8jD94vSIJH9fYH
Z3D3KZLzTqnBVhaWt2LjiLd3OX4R6CAdMiKlwpqO9w8rlgOgw6vhtdLavKF0MwFc
vj2uJCnH6lE445MR2Pa4Gv6na7AlUicK5/LsrP9cNzuC4ZpBhD+ZZjqJkgP9Igsl
JwEIxZzJcVn1DinMQnSD2DopGr9qBL9iBH5pPYMesOI1fGVN8coWTj+Gd+Ug9CWI
WeEm6HIEEiWnhLTUPhc4MZHOwhRqOdM+mCpNCYPrOaWxwWxCxziNfo0kB+5WiFBI
cqTmvSa7XIqDXKcnWqrUk2J94rW6NagAgoaoXoMQ1i4Yu2gkxJ0vMvQqrZoo+mPN
SRvP/KLy6wqgyAhCNyMVISZtjeRbMb7yAYKgXp6B5HZQsbFTyPP8V7XZHO9gngTN
03eEL9U2F+MuwSpnlZsqgyY7ND8OKxhLfhUn632xPnf1Y+R0WkLS8qUun2sIdtj1
I8q7KoWdLj0d+Mee+1+5dPwpg90m5KUStzKeUG4iiVBPdH+V6q3D8NCpQn70gm8Z
n22esNWoTXmULw2bL/0f/w8Qx1JzlQmAOl9xh4vsEVdsrRofl2jnN42cg3TerLWp
w2ppgU+FHC5ewicFUE23y7zfWqNUgQ2JtdnxSAQfnPD5hpGY9uIRGOctNXY0tAjC
WpT2/5CDYNW1dTdvNxp9xee0wkkqDOkW9JZpn8P0F9Ddv2VI+Wc74RELHrw712RD
8FX4dGGoB6PEx2cNRjvqT+3hnVa7H6h2chV9AgUua709IgkKO70fO5OCVVSbuHTv
ZBBFaRiQtpzpIhNf69yjU5VdSOx/A6/VIsDcraPPKjQLFSa5mKhMhbiFcbSbpMR+
U28t0ygbAqxbU4KcLLBXh0NFZUPw4SZP/0KbgdKc28stZAq174gh3KPYLyLPcdi7
lngO2Y8Q8iK9kl99eM1FMx4mPTkfmb91U8wnxiT9Dmbofg37/PQdtHJyBjWkVNIk
EjpJ6yPXsWJG/o/YMsiFwqeunJYH5GzOpaullxMdqcKjps1BeblwZYG+0mNkLPye
RTzmDtT/dTO27OZo5S4fueY8v/EOqBAWTR4upI7AGswEgyuUQ9nbQB3/QHYpo8Hi
tUPWP19qFy1TZc67VKYV1DH+YkX4szzaUYd8RgpOp4oA56txkWP+kshN6e0/DFIv
W0QJ8RhP/AkDJqEmT0LOxsTMuFjXDpN1xOLntXM0lkx+dhKRsS1iqDZPoznUufyQ
VRrYcQ32Eb4f+Giz+0PiKt3aVFa22hek2gmoTYS4C/8fwrmqWSY2ZwTOvDiIRILk
KAvmDqzUSkcjXNpBYCmNRWhHgA7QEDXFlpsDVbbkTwhnw33+u0AsP3h5uINq/2qW
//upvGaM2S6Ur5xb5L24OfdI4gJgsy+xbD1ZBCcIJBwt901e18MFM+4bt06qSkkD
9uP6zZMZKgR2ZNZHALIuBUOLe1yTlD2Smb4Pcp+ep52jMKAb8TjdJu3E/UIkvl0u
vRfvfd2oiNyWwcldylykqVGzmuOSW/ApqtGMR8Opm57I5IzSIG7EhvwFHC+dCWdz
T8k93v6jzRLtZiJzSltZbP3QtM+avsVst/hIPc8l3I/ytt0PwlJ5fy+2dSQaB+uE
0JyOTgQS/OE5FV32Rp5iK4hGr4Ttf+HzLKLcPFgYTK4WyYgF7XD2QdYD8hjY+8KW
umZwj67T4qxxnL5z2f33k5nY5f59opIiDU5q6Tb8PD+QjPL+RxK7JOgOo6C7bKAd
XsR6GvKFYUIMTBlf9K2cywNgNXvooWcMDRvZlvmTNCCR3fzqHWo28Tf/GvcHZNgy
I/Q9eCTTFkYpW0tMPYnvZSzaiHAHkXrfYsjzkGXLAATB/bSplYVbEZOEwdcrl64a
fpbq+RnxKs48kJRn2bPZxz6RC9oY5zBuSiACCOzVC+wjc4xJ/962Z93xiW/n8lol
lnr0HbZduTG90ihvZH2yiAUvb3dCenSTGkBb+ygyrqWCZu/79vj02kjPT8DgvLlz
/PHH9vrlLKcVDj3aCC+oskypktCkWHousVYcT0IhaSsgQ/6VKjOMgX2lp34KVJ/E
ZXMMCz1uJllsWJlTR3BLxQWY9KHIqIxzRczU78d6QzXz9iT1hZcqGoZHkbs9BN+R
uMEw92SsovLd7ryo68297rMEk2Ih/Fso93MD0xU/+5CTX7CSaa4n/9kSxEnhz57g
Jcw4VLujTAaXEM/rpnTRvZRXNpYJDXZpcifhNcLr00/06r1hIiRGgt6CajhrVj8u
hYADPAdvqIeA3fVVenr4p8vADV36dU8tFRmc4M81Cbj46gSSzeBgLVGI2EBsU91G
jCPcOf2QjJLaSD4pCRAMPa6lpDnb0t6Fi07DTJWhrhj0QCiv/HR3IjZ+5F38tbu7
bHeS/K6Fd4nabflqgzGGG/aue3iXwOV1cy/6gCmA1/o3tkPvFAVPw4k2Ls2Tisnx
LiZ47tV58kcVZULwafpYOBYoXox352q5RF8eJ16HFlRxIqz/6J0BwurNh9JNeHEL
hzrJjl4Rbu1UKGUzsu099cCn/oVszwts0SWHSVgMbino8/VvFUsTyPz54/Qql+Sr
GIcdyoTj8cJ8N/CvMnSteMPp6F62r6Ua6W21+P4DxVEDbfyZNyJll046qY5j4vzJ
EfMg/xDcsdIwkdnuU/VU4zBOwdavGisgO3JwaFRo6bz9iB65+37wHgWhv6UOycWJ
wzcvWZMQ+nsRhUipRIaKN0uU6vOjMbxQdkxj9kOFJqwrXjzHl9KWyM2yy6lSfLpJ
xPY/jPQBH/rttKwD5Va71vt+UG+rp4sFbs23TeFrFT/8YtYNo39ovygtGXmiwuek
PtjFgaMUH+Mo4uLKdEh2caDM2VTuAmefZgyB1dc71hU54KyJSZYjQcDZFqqddqKQ
SKn9qKPmO3Dgrk15YESQ5KK3I5pGiurpxqZzt+n4xVBmul5rrRTn8QTKlMygqIWf
XWLKGIRDoqbHVOYKHwD73tnIe8NS9+otpKDP45zTbOZUMzepKsGoWIny6X+j7rhw
FoHb60pmL+jkSsIPL3y32oSAuw/DBAL0P/0CBgj7unW2LOUJhKlAxV9sofx0ATAD
lzUIH1Kf9R3Q2F8lGw1f9sX2L0K/W2iSDXGmaBpc3RSpey7Qh2t7HrUjFwbi1NI6
4zHYg6R8pjggoPPv3w5jSWlTbvGFtdTGKOATMPHfdqpHOgnWnqQubAoIOgBC2uFB
B13/xUMDuJ9VpNsHsYL6MPpVnczKqZB0YjtnbC4/PamvlSMZaLy65xFL1Y6TKc/g
KGD+ZoldEf7/loXhKCaXk3QCAkVYosfXZQF8rzrJV/iKt4wafV+fa8fs8k3B8o9C
hIAot07nAsI4exMo+/PGPUEBN47yNp02fDIXddgd4BSBLMMr77/A2PWn7YLYDbsE
TVTkWADXNjat62hY+JuuyR2LoGM3gId3KhACJKKM7OHacM0pSEPSeX+G+ZOvc6l4
BOJta61Vmc3ZGqMRFNYvorXKS7NVDwZ/a3N4eDe90XcbbosGmI+tbW2prQn9X2AI
o9CK9oCWvRmvgUG8u3nqDIh6gOcVKAgawWTZIYWcl87upxIK5YXuXP5jwZ8OoM9c
7aktV4hF3/Xyz2RXzv8WkbPhDom+7a4epQ0MTePIu7EhvS1yp5CEmzhLgV1e006S
3opoYAwoyOSBXwWN+NNSulvae9cmDuicKq8DMDvIwAQ59O6e8g7tvyvMJ743lYnH
NXS59VsIvP/dZv2gYvV+1UOp3U3HLvcxVDpidNSou1YsF0PDjVsSDFCne1oLHjCI
+fToX99uYWB0Nc5gpn6xeRGcqOLOt7v8nF5Tfafo8M+Q4KuKKwjIdMETXfYCBZ66
aqdRqjnUobRd1VEeMtw27dPB3ESkSi0ai9JzVlGFMJVooNZT0o72N2AE7g/JzdWf
3XJVi70noI+sGmkJaOdzJpETjoG1xCXTSUocT4gCyJAWIscOYsyo0cSpfGEfNLLv
uA91uOhHzSfj1586f/wek2jaV/AZP39ha8uv9WYwFxHJKBtHiUoy5XCJXlIJl8Gc
eq2hYe+hf3dYVQKVpnJjl0Y+HYXmwY8F+LaSfh7hFm+8Txbx/IciAzw9LVZC+Xlf
5+7idqOVChPcRRK4zYqseOuj4Apj6xf8qtb1A+cnHWy0CVtEmRv6MCInQUxqLZbk
JCSUYaTN+F5MFdgY6F02TYAwLpxJuZkiG7ujGv5JIfb5JAecPaEh+elHbIcNc5h1
kmeceln6WmmHH7ThYq8eWZ91CaYf6+NYt1BJP1/nuRoLJh+OyXMDbpQEHB3wlCBb
9tQKLAlH+CF9gTTQhqmB8v3tm8VKkDVlcWjkbOvCGjuKoOiuGA/J/aGvPXjrR1Ij
Sqh/QfBgaTYsgwGP1PM57HLn9C/tjZoXNc0Ga09AyJwAJ9XevYLzjMrDEzLEGvFV
EWnBe4Q7LOo+3W6eMdWKXN1efuVI+KUgYviOxlETzM2JAoTjDDw0/QlKpcC94HpR
6HNeiwOMtc6hxJCa3PJ72L7G0iBDK+0/SAuLu8cYRWoOGlQBBT42hOdRXsPCFdeP
74ftShU9yTkSeeNrzUgt+cBWnbI5QQHqb5iNDuiDMyXWZRyZngjbluSSPiPbO8F4
2Ill0YUlP2SoLp/WAyx22sbIHDxGvJZSQfEkwKaEQZPvL3mPhgkhTTM8PkSPBadD
khm6vd2e5kC34/6UAl3T1K3bd77CWYQKtMr1C4NNLIqW1NV3Y1NLR3PJEYtc7mx6
BLtHeg8FAxkBgXGyOLb6AqFgapKjrgq3SlSAIi/rhu4TtMO5BUZPZNk/Jdf0WBgw
L/L3WblH9PrQp8JkHWIEg8ZnAws4xyHP17UABrrpC+tUCPQcMNUmKe1cHYxVDeoC
jYcE06YRAQ7PD7nDbymFxUVgqyqwctHczaThC+wyslZMoK+W2+hD4YFJ9LgqaEIB
/P5s5bYXCpE6vHDYlhODYtNV1psPJvYZ0k0QfjkNIthsBxAP7PGRLYwdsMxyep6E
8NdpOBg7fuug4HYvZ8E1Ag6ydQtf1x/IVvdbg8esIejQjV2678Sp+pB0vQz87oWy
pUZ7pFoJcKc4ll3jd2dAxkybumvDUKSx/ppr95p9bTksixt+qjFtRsAwh+x0Se3J
XVzNZGZaJoglL9HqcxyhlGAzXpBlJHUoGGAivw8hEov7Jo7I8LElUp1plulIQZUo
7awXrFoXL2DALv6y2tkPwTKvGjt3I4QV8yD7nHSbwld7f3V4JGFVNkxMUCpP5FHk
njrSUwaWYqihoQ138HL7a+GQ333BLRWWNOCuX6+5US+tYLl6co0kr8182eOsGFd6
1dkofS+66p7Pl05uN4kHjGo0mLtl4LgS8BMUUF6EicVynKHMfP3TofwAZMpU0ncc
AhGHfh+t3mo18h3ueKxksksCGwk7KMGrlRaO9+cwOgwOUasgF2BUAKG6AXH8hKvI
p8pV/6Ytt4C+EFl4k42EOnB2zkO+4l8g+l4UHqnRIoPjzhPhtooelXf8GUjtQeKz
R3pWvSH7ae1mmRvTyuG2OjrLuMfFENMNR8h/ICK7LoZEA3BYjeega7mGhdDTqVmD
UjjFy6w17emAYPbzpg9Jq1UURYxvlRv4eb5iV/zYQtnmJAgJ1J83zL+VI9QBe1O1
bkWMWxA2DKZMOVdFEVloEzt01PX9/ayNAQNwcDDqU6gRrdCbh3ae4msth8rQizL3
2UEoPv6pI2SvE24WByWMpQp1ke43FXAHEE/HWy9nCXWvUgdWJ4pWX+6WIQxdy5Wz
Pm3vY9G2lNHvJ3s6IU2oe9U44jK5seXO6IPdMT0yTvcFNvlN0r9nbXVtMA3XoIVU
yOAKHUkrIo/PZ+AmE160BRJTBoXKYM/nDqA/NbH6YyIUPw1WCHx50es4hrzgA4fo
kmBKrlllkFr7WYQqZie9P78rAwhzEhNw8vis9Y7y2jmLJ3h8eGjXTsjPK5ak2opO
Z5rNlGFQ858tOp9yUUwrwvkXMDVvTpZOBsBFE8CD46wTqvLgRE5th9WcdKW8iB9g
Xy68J5PzuhUeThV/+bFd5sjfLWS2HT+w9XhP+rbomsyAAxTewNBTdyFnCF+RtWsJ
d83dNmXov9sgmS1KJQOrP3cp0LdxHC7F1cW6bfZLiKjr+XPzQz9uu23mwc/HVfkm
fEBwsnrgQv4gBO/KCVrYsaB8f2LeX2zGsB83dz153Ecvco+waTluVmhGRS7hj6vJ
TGgOoYuVvBtUyz5qK0HfIOE7QPV9g3NwjhhziMhACJR01d6r7S/X4CEOE3MAbQVS
oKbn/U1lZbYEQ2s8Hfu3c1X84LxSTZ7H3t8/RV+4z4TW/DtEBS6Eo6HMOWhVEMNB
gptmFqGJRq2RMgkFMwtYJyZ2wHEyoIppCdSagKeFzk4eX1k/ZU8gQOqtrmXnRs56
7HJ9lpGwRq67A/TsD3NzcwWn1cXkJ6q5q+Cz4zRQhAJU05vrYk2c4QPJnG3vFfZ3
K8AJ+/oYDSE0bBNfH7ECEWbrBoivky/00i3O3++R+aftySE6aUdGHhj/7QYptkWP
dptGijs+T9XMkYguAfCfFoD5dBz6uDFm+7ufOPpZDcjOwljBFzNPxAhf9sIfaB57
L/g88LYEBFjrp68nda4Q8SScB1eBm7vHhCJJRIhZ2yUe2qziYb5ykLnisOz/wpgw
HKDXhlZrjaapphjxMqF27ySuGrTnOhCoC/7qrG/LKeRD01vEGV3KIt8e7M5w50wq
aai7Sxlz6zn9Dg0x8vM2XwxSNrDGHsKjQpqnQgv/Pi3WqvsrzpYESZMkT1IY8PwK
Tn0pSlC25GVhfW8ISFNlEmlUsT0A285hopuS1a8wTx+UrDyOFk/UucN5OVi+cR/N
3nYiM6gD90WF3LaRo4a0Rh5CP0CueoCDrcTqB4eHbGBZEH/svHENIfrdTA4z0G3U
DAXOi9M2TWjNPAlJLeMg+O5g7bQ+jN1+YgNUBP8MGRuPC2IX9lGzRcO5h99eEIjq
cmPy+gy8Qa/KuEhVyzZDf/y8PpvaOhpfo7eEVQSIpHrunVnaVzIZNNB9bFL7REjQ
z5kD9hoRciFzAm21IpJhcIn8chjCWwAtY3etV8O5aD520Y7q7RpkHrOabkmZgPin
gbav21JGIBSJniPwnG2EL7NyMbzG2KluWORta748E8ug0KtjSJk0M03O6VTyiqrl
Kv1w2fmyZNi/EsdhFGO7agI1xR8XY2PaFCY/xUSkSTul0Rbs/5Kw/mS12hPT4nu1
a1OeK2uHjA5YvYrboHUKglLcWvrP58JeFmEtYoipb6zwQnM70BvkHnWjFDqhqXBZ
wwlulL5yTwoT82WVmxI6rqVb6uAC9eciLl1ib19plNf97zsPzLd60+zvfE1qVoL2
QkrNGpoLAxjVuGLSdyT6gt3Y9xnixIBTd0ruKFMOPpp6ziFUddGJxT7bRzTkdeZW
P+nmeYFJYANywENwX7FpAR0/vXAaysPOHisgUdnRjMLcWeaoqMIwqNzhMZMSxWqW
nT1ISZ8OtMrMO48Mgl5bBWzWf1FcwaWbWkJ5NDtdVSlTa0fDJoT8VTQNT/2Fp6rn
5nFdjf9QKahq8kuzt0Bgx7uJS/dME/G0GSFxpf4u6qLx/2jcg8iSi9LAv+LLknHJ
eVDkfvcufFdMlVLtbnngMgfInLi06lADNsnNh+C5er3xEdym74NYHgMdtiP7UfLF
Mz/WiTAv4HEfnRZeUXnWozhAQcC+/P1p7THQGY+DB51ZMD83OJ8ZWAOzCOrhBtG6
BJEmWsWT7roKciZ+1HVxWz0g/6pEvzqg5BdqZNAa7iaPyRuasgSgLIAdb/LjpjEa
DH1IaQhgP90L4/Iw0gPjEV1YYarzWfZyGFfdXWgrTHt5IaLEFFB+rlretAo5t6hh
43Zc2akvpywTwbSd9R/x/aDE+jtOKxYSNaKuJQEMjzFtAUPUwJ7oXmPRzlCaqAT7
w7m+SjRHrFrSEi4S0ypcyL7DJhpbXHalRtWf8KR7cJRCAUjwZ5tPuBpx4Io/qJsq
1117m8N+mqdkbCFsv71Mlf0O7MQWA811x8EufE2Q+nIeITjkFd8G63mxbsbwcPFk
ebqhLnQ9uRTJs5nBGU/2FtV/l+s8HQzN38oJFqv6j2tQAfa6+a85nHcAkd1ITnpe
BMJP93bjtCXt+IY66I93dAQM7q0zui3nA9/WiA4V9PdkLB9xF8tAr8gYSBLi+FpA
gYHQ3S9v0eQ32VgwhnRjvKJiXVYokMYj6uL4G7JwgUCmRs+iOTG1AWdLGlMAbgC0
vaQPDY4D/UgilxnUtpcu12+910Y2fbWroYHIlieMAAQ1kqAjzIM4vICEZVqzjg9X
mmrvpaBT2gb00VaRyFWJ1gS852FAVVvaofgNg7wwgA24TC2bpz9KsaX2z2RDfhnU
SWuwkzK9DybP2fnNKFBvdcqiK4MQP71zVSXb2weK55UemPXuMgQCd6l4KjISFPyM
k8j/dQQNgNWU+y6tbVDjAdtWjsfG3R0VnIry4oAb7Ag8tMWYFS96NAlQmUfgo/y3
523nVy9Pmdit4KjJRC7CjJXbIwvlcS3iDlIxsxaE48nj6TZdBXI/reA5hdy5qwJw
C0U2+i1yuXeGM1QuIdMeIRBSAfi5ecn2I3/tvRsbT76rZ7Aj6AiOkiKca4LEl33k
7C9VnQsj+mhypnJjJ3xxKZtiS0xQFCZjwu/2gN+TSIy4Fi+hH1UjdF5UGLMbNp5h
r0xdzxSs/zJbt3hvGShmjB7LH6nwRMPcPYIcCNjEPvvBW4i8HtV9WMpngpygQ45h
D4ijuLNnd32p6+9qL9ZTSalEa1cneBlJMzoOFnThd6HcqtA/UtjlavsyDnQFIaYv
a7mKRexfKMkESnmEDLGJW0EmkH94PVx7QHlhhqtdpacyGlO7iJ0gSjAIL/pljF+P
d8RZ0wz4uMxpl2SXVckZLnbELdZzbFonA1akjip4kWUKa8NuTVGZEg/LHH2gceEa
zSU+GfGzG4vorNwzLvcRnHd+Oh1t9dc1eFYbuTSZGJ8oWzFm1NxXjrShEfkQA8zl
pSQ+K6BMw2MpEjfKFOUZHYQ7Us9zK/S0UNVDnDUOxJBmwd3CAjWTqVw3GnWB5tYf
0L9FXS7ed+8fPSO8nB3vOXsEkB4Zx1oRZBL6gw0F9p7nFXXmaVYdtsiFFcxQNEUc
3TSwdIE9IuQTdND+LMKUR8hXqdkzcUPGM2F85HlsUQxBYHCWlm8ZjZCyx1y+hzPr
U4c/6SflZtbYJqmCruE6s08Czp8WQCOtt20JK6zZH7X12QJcFE2E/vq3Xvp0Yzab
0p8P5/ERbhAXPU675Lwua/VIyCPtzef3DeuIymtVehCqGMbygOfzk7RI4uS+xGUl
y7I4Oy/mdFGoIm5a92ivKOh272fjZDXKxfD6gwuL890M/+TpTRUuF8I2PAWcyznt
LpRzWR6fEXgmGFEQH65VU9OOMXOnJnoVFLCnvtNHsF8xiISM3a+ryWwDxTh1WJGL
iwwvSJB1kCIBvU6sBPmU9u9Ceq5Wdz9eDsyuMHfKD/18mO4YRE6Yiml0REEaxfV0
14DESheebD6KLJ8wIkWbzUqXfSTKajZ+yNI7ZXzBAz3t2DGD3JzSW6k6AoNYFe+L
G1T23m480M3+uqvT1cJH3fJVA04jcxJEWB8S5CEeU5ibV1xUwCmlouui79OArI+V
4guw35ucmWGLzzr5hbMMKaq/FBrriy8VtGFv9dgofrnt43tWVKEfzwvmmuXagexh
lTfVdQ7ZuADdQPIhOLjoFYAlh+JQKgNCU1lz2+Nx/1w+jzXMlUg4ozKAhYhMS0/n
mRDxNR7JnEQp5zLQ0UHvtQTWg10M63Hcsq3RPlsrKWJc5iNqGf5ME/1aX/wPQaJ5
idNzOrBn0Ixl2FRVP2WBe0ebRTny6my41ZwJLCUZtp80fCB2LzbV+OSO1B1hVL0s
rJB172RDVaR3PQAnNRiuBhQdaqwGvf2qwB+f5IKe5KjKkigO3swgbPw1JhURNmm3
lkCYAuD28ibX5SVJo7x6NuIygk/9rzIyaXcJu9Fkq8tus+1lXDmEHHnOI2hy+1v1
ZmuN3u8swMfwfVRwi/LSbdawdf5RzNB1MY3zS9RRQVxSUt8s9j8zF8khVxnOQt6N
HDZMMedzJM3EofNkmPkRBb+22wpSxucU/KwHjcQmo8JaDq0osP2fqh7Pr78nu1jz
sD/U/Tt6PyE27P+FFcbqQ6dJozFwrI+0pVAkeQx6LJeEsrwvJArzLeSiC3MsT2So
VGEPnBqFW01GfhLa2zD/ViqzCzk/KSb6bp6MIL/UFH1BN6vpp/zJPG07EMiO+kEl
GCoLmHDc2TD4arfkpQxvETvprdU+RW4BSm5p5StTkSsBggHHF0XUVQKjasaNXn24
HZxyJY3vELBMaaEDBs7Zi4ipkadFxZbUra7652+XkYAoCyrOic0wr1zxdf0bpIe2
vzsyfKkVKkrCf0B1Z8HFsS2zUJPvPYK2MWqBvYNxaZ5Ry7UPT3s6PmkwYPO+Oq+J
Za1eA7sESkqG4u01h1UUUklgfxdeseFMYxWURzalfpQyOXXWKvXMmj3FiwX6GcBC
1u5EhCsRy7BSKXZxOs182X6rCTfETfYsKPS3/FZ/0RsbdixvlwG/u4NFORAuTj/x
zL9QoHWNQ/GRmaiDDT7HzUmESNHIb40aaE6AEZ+Hyz+Q4jZ1lkiEhND5hzu6yrww
8OnI7I133iC+qZpkxo439el9owKgT5UdgTAhIelB19920+0qEAdx2DxTlkoH7/HA
dEEcYl+jVVrifuqq/FDftJe7klnyuJUrOy4EmjLCm49CZvQUvkyuR0py21SFbMgo
0QYMF63kHf29+MN+Lncubyk8x8eCqBFdT/qflP+rkAh7BcFhBw+WiJbjpMnYY8+c
gQVSh5j1w8OM9XvaFBbOX/iuogPNNDRH8/4jxq58zDZw2k4HObozssTF4JLM2UWX
L63ZFA/nFtyGEQP2re9+7GAMhNp8rlZfzQA3EFNWmaiguwOFIGcni0xFa/aoaQ4U
RSrISKp+3zUe8yE0XZw9b+7kOoF7QoPw2Jm6r9oZud1kJYfj7TK29GUBZBcrXm7y
i+AQ7yWk+bQXHmam64nDy6qjx/Cis1wJJjQVJKR78MuEHHHJRL2ecCCCKoq7RLnd
K7a4LgDLbKJ5ZfN4ml3WMFDvdPlCLK21hY8nCzR6/Jvsfuu/pPeFAM0mHOCoR78e
yjB2z9Sc7rOGva132UlhoYBXkvZpQFgwaQOvfachLnvq14enn1pOk05ugrMW//bG
JsWKI1QL3ZFZzadIkmm63hIhzXFC9MbQSKZgz4zZaP1gHdsAMZYOapKoauFRIfCD
CUnFeACGpuWRxEX/lpAPODbPbAxhiMuKmYR7pIT+VzhJ2mSx8JvcTXCLmhbdmqKL
WhpklBg1VYzncuk5DH44/IcolXVDDIy6bIR+l7IhT8YokXOdK5quPUt9v3sT6+cX
JH/ermtSMXq1z4WYjxqpeQXEOjqW8rcccfPrAiiiCHQVfF6ttYQbTEkxu4zel8Mv
yIWNbriyZZuXizeguf2eXnk5BAv7+IH/4PW4Az4f2GbR5qjVPBcMpdnKWyulz+0k
aWIjnN5hvKdAtrTGexMNH59gdVRvV++5YHxh+3lPSWw3AyzW032l7lJPDEIlxFhE
543dRhw0NfXRYxEq+i46g/pY7yI0Az8bbJA04fCspk4VYhGRel/UCIAtHKtBXUww
fRjsvqHJ7IKWcKZbKRZPqo+yJGinUiQ/7LncxQ+bt1DXB0rrn2BoZcJXk87EO5VX
+0d6hKeDlkXE7ElKfa4L/xor28eGC0v+vpmy+OA3ymkRQH/W+z7TwmTGTm9bQQrC
ATG0gbF/5CAkWcl2nVgjOqYDEOkbkTGQ45zPlf7a0oWA7mmdE8KeKNO4+VOhFW/7
D+lne4dAcfNmmfwWv4PdCpz5D4f0htdbqdCm7SCM17SDix4qj8vbr4nbIfCMfpfr
zwujIlZVrO+yyZ1zX66fHw0RLcUDhBfcLhCBf1xmj2r/NF5L9F+sILCDDC/+rrdj
T9rsThqkozdROmVBOEvfbyH5SKYdhtZlaYUVyYqa8ameJv50Zne0zX9NJv7wRUCR
5QnySWOMUJtGxvvInZ+I3vVTI/SK4dRsz7PxqObdXMWRfM7wPEUav1qeUagg3N1s
vGCJQN4ORxLedw57H4zdAUM4f0+Q0qzue4wuwg2wAM59N//h6qsoBCxCE4D8gd4o
t7AaWirEJHOkUC9Z32dIhh3X7hB0V6djYcsN48B39Mq6rieQXeOGDW5aX5IrznY8
RFdIJmxButcmyJ3bn/cl2XIdQ5FcqAtVcb4Y3LRMKx0O5aauJCU0K1hL5DsGYaaR
INIy9Sqflo0w9h5musZgV6Ytk1M1EOFEXcQ1kmxOiC8EmlpXgOc0dJGIc1PeWYZo
HUkdfFJFcwiOYk/3MX4nquQry1bUcnwoYKG3MBeyl5Q2cX81WXzKFLl4ctO3cOUh
8W+oxECYKTv3Mohh3mJ751UMvzCf5ji1y5GYOsRIlxj9WL4wBHWRvckZbITeOuL6
WJotg8g3IZF45PqIR8vMI22XDE2lwPNQhhEWqIYhg4RED/nJFbcSOUxxdAtJdHUf
VM004DGXy9sAGBel1UovNb4TRGh50iVjuaLE0tCIsU7WVnypK+1sFi5nhM87UTS2
6BAPftqVjp/xdhDcbo7VeWGDMOD/K96iC+caV6ny/n15Q+0ierg0SY820RMyQDfN
+Pq4al1Kqi3vD291u1gbo8eOK9N89JQQu1bGYpFc62J9ut3ZzFYcNCDH3+MA9DEz
L1AebZdwgF8YIwuHNvcnN+B+W4OhuFIK+0qrAN3SI0EAqhuUD8QGTc1tctCQqfod
gDm3ZofFR7etuFlUUbOMzvtW8paWa3wzjGcyz64+fV4UomeKB/l5tCtvEMiWOCuQ
CW4AQCop4l1fumUAXKsAf5c3t5NcQcbYsMUw+VrdOYF2mkmaF2b320hurT0ufN6j
VB8qhQwGiC14C3s+p/GKpNLNAES5GnXDx5wlLuJyPl696wh6PU4Zy776T22DO8cZ
fGvWF8gnQI5tZJGMHMG8NOs9+GiSVWI+fu7TDaj73rikG1QZ++yMmRhf5uQbFyof
CqlxavhHhjLyOzVK3Iy/lne6EOHA3IMV7NgB4mcz4zP9sskakmY9+Gk0IvCC7Ube
+Ozpd2QxpP+e3y5agkmH2fvOoweL2Mx4j6CHyG4r1DgFvFVCuB/3Cr+PNH7RD+Qg
nAZKDJRlDGeEdk+u4a6r0t2kCTgnWrAmjCMVgdxgOKnyx9+QfNBpd9NPtg6ZfQfd
LfjQi32PhljZ8A3A6l80TTZKFYQ6NlmpTQaD9IgWw0jVyQy5GLJqqmItT2XFRGS2
jMvCFIn1hnKsTQjs0W+mgkeiSAzqqkmh8a9xzPXhzaaGdhRCC3OEaarYHX5pqhfM
BWOhRNKEBGk+iOTxj1nhhwEFw3firYeiLGr4YIkjywFtN+31wC8NcE54O7E8NC/r
PHRlwl5Le6zvrMGT3zbQ3IiNBHpkFnwC4iz9bypOXVFeFKACZdDk46Tgd0pk7H/P
/L2HVKCKIw19cRcKxRSL/qk5gRHLQCrWVoMYTV8NK1EKcyanE1mzxeZ11E9pV2YG
0+1ujrwHXNN39TTuv3corJ/S45a/pPBmGVT3mUh7cSNKJMlwIdXmFRVWZrysz4An
0/Pph0QcIrj+NxLcQydBOdERsgIv3fcazC7gBlIoh15C5k9YPLySqOrDMIBeFJ5r
RSF8bM9f53WnpykZVU8QTdL4htzXJJgIsgqyew7lHjmAFdkZBvWX+PDOeJNdrcD3
MVMa+x44fBYfG8BsTh8+KWV7hNnqgTQ+arV6hNMQPR9gpdKHizcSmXLJKSzs8E0L
yXTBoKzUKY8XuzGGWOzqcSxF/dYtBtvF/f8XW0SnSNK9BzcC95ucz80bLcmCzkc0
AyrVhIzJes20aATXUdlI1XRtVSX8gIY5NtXv06bJ5166aSVnzD2Z/0qVLswNo8nu
ss/C80KizGf3+j4VsFb8fo+hXlrQhpfjxBO7ljOfrzfWXJGPgawvcLmIpn6uWxHS
KY17douayjs5CVpUlIKRYFRvTdzNILoX1/OssxH8T5eKG4aDOt+K70JgVVoTnf4S
zStcDmSOiI+enDCI7h//BcO12+3woOlbOjExpdlmY3REhv6LQjYiRU2RjsBR3Av2
irWPbTbYe3VUNZGTYDrySksWQSUWzCeT9B9revZgPM77SPEcIbTqYEmW9qh7v+Wo
NUhVhOSGsUa3KD7NtIWksl77D9x+NjfoC7qeXCz6zwA=
`pragma protect end_protected
