// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:02:18 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
UrnHlQYEKr/+DQwNzw1EN9VJQJQKFnQu5eFZoK9UxLW03e+y2aXf/ntmuKnsWQ5V
f/MWb0HAUVctM+8S0nUMZA9sXKuPycWX7jT0obUgnOK3v4+Zt3Rpym3SPlu1bBnC
27DDOIKpHHcYf7T9utE8FkfKpVUpc3VzSf16shk+AH0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 12352)
mRz5XJstJHHDU2YXpFSuMoJfd8/BOL8geh5OhPpnxH8lAA86vJfjiBmPjUDMWDso
1PLiZKw8q7Wj/0gN7CbHhhSmrrA6V5GJwapn/rcCwn9UFoZvOYto8qrV9fJlJETO
T9tS3i/kcInPabIhAJPNeuaFK+o5QmaKtdyTkv63fsn/CuFSWFyzxQtZuD+GfzBg
gPCj5oi7RHr0DWCC7w/kCPyro+QIUp+SKpV093U2BAvdefeJyPYlzBQMlXAUDZZ+
Ej6MuE/5++nELJvIaiNZ/Yj/ivmVgOmb0YOvPwfdMJdMQkNF5NTSs84vAdpH6Ciq
1ZsCPLcE6lTSEEp2qhorS6xAsxOZrEyTEr8WwLKUs5lPdY4S6qFBGVZJQGek64Xq
+qwAU2f9J4j0aRwhEMz+n82dF0Q/jhwVZD10y6G+oE7bBj/7MUyH0EHbRUdYzqhH
YHko7Z88Mge90ult0zxPYk1ykdY0JdwmlfgZks/dwdZC2MZRIDdxJlRSSSspAcnN
BNASEyJlQCbZIH/JVX56sd6FzCqNK7IcQ4THoGe/hjRDtQwNJEIEMuiV5wk1iKpP
TW2BEcNwhV91Ioa6EIQdUM/D+OOgz9PE9zvWM/22PC1MzKLTJHFvQLsWt1Blq/zm
qo+Yr10Tpz7VyczsWn8WysHhyc51PDZYsiSbFfOsJf9GMqLRII+khe9RhGjvxe71
EvhjzI8oAwh5Q10k8XTvm3YGlIhm5jFuL4zM3JPbIjklTdMC93lcPOCM/nolN8ci
W3HOmaV5PNV1ky8gQ4DtWl+3+g2nuFVI0LoVtvG4NG+Z1kXtuOzRCtUqRRPZqwUA
x3BfjYlrdHGnHj1LVglmjxhtpiNMo68NMRIK7L5ga9O3fPouYdscnRyL5olij4Hn
cRBcj3T4jqWSbVzgEyfZwRQqP34kt98bkFhEqLQrvwm8yer7BXxyshPV3BoTRBJu
+yYc3stweiACJ03rnqCAN/1iQlOUOfu6QTsYpNIQZdR1j9bGVWx71o0cxYBSEGAs
OeEW7sz+u9pYKAXP5dny0UyjG/x0rcvDw4dQO3jo1NB9meMsCuxYifE4AwS7vhxD
8XindENGoG5NVHFqAoG/zp9PmYb3fC0bnYjv2RLEnqsKzC3si4wRDrsAl7HKpiVI
dxoXwl/2S+UORDsMZf7j618auyP9vKic3n5YWieg6fHlvqABUa08XgF4/hufEBmM
PwVugDQl9roBXiwH2jgb8oCTGoNkjLLickV8OEbyZHppMMGyqjKP8AwdZaCCDzIo
qSMpUr+RPw9Shi7FBZVc7dscu6ICQz8BtnI48AXflajaAS2Eobl1t8dn61YgY1Yz
69oJnuH5ludRTwDUKPYCb/PrhxgeBuq+JNXw4Xdq5MUvAhK20KtKdC8y1ZrnExqL
eCKk5cHZlVfziN1ZbE+ou6Yba8B3X5z2YJEGcWLIVlxT9Fv08VeC6e5d89d91M2l
8Ege0F6yGkx2l19O0iYpN5CAAskJhRAt4d+DIZqU92SMN2ttyKj3mWWnpZitwSWh
cRsq9UjJH1pSZdwXGheZlmE0NgP+WuzYqSXbsu28l5Yt+ARe8wmsEA6LIkEYFjA+
LKbuvYuRAxWIyE3sOcbqkJ0K1Wyv7rM00vNaThPcHWaGhK1B6OxSNoDCi+aWKXZy
+RBZkc2qDjNueGTWAnD/gKPDvxUZ++ab2tSZpfGE7d+4j4LDLejtpyJutBs1nIx3
2cUFEqw4Y9amcaj7MKo/9bRR04QbdlxUZ9EJ4HJqjLuShplCSy4vSpQdsNJnh2ve
Z2ZTDsgROoaToNPmYwdvK2LHeaOVEK7u+VA+9QJjKQQ82FgwqvU3f2np56ckNodu
5C7XrOXd+guAQjetsfBOL2fJ2eN03xqJq0OM52+2weq7s2RZSVkl7GFKGsQo/YZ2
5SB3/NQ4GzkMT0DwazIX1c7/LC7dMeQTwvUo7LKUf3rH5ZtkgYY0WN61ttZLigZv
sm1Z2k0gxkhG1+yCL+F74AfG+LQP1ADR5Z2XOxQO/7uFJottrqv2bOr0QBWSTZEb
uqbpbY6axZl+OhUz4lGujOojc/zzSUKN1iVposMxEwZ8gQb3kNUOeBTSPTfe++wH
PnZr8vsXCcvbucS9bwjnUuX7nhhzkNm4fUjN6CZUWqbQM8uL8Ux8M9RzBBWD2hKH
4qOap8JW8sVJn1KjPfecN4X8AmycmXmwJIs3IX6WV5+kTLQjwvAKvmnIBFt63vAQ
Cv2s3JMW73BUij0iBFNsS3P50NTwAauKviZpykGp2vRDvWxBaN09cQ1fuorANoDZ
LjKDitxPfXZxC0/OGxGEONKdnP+6yNn8uVxhNVrXMb5NHu116M3I+m0g0dmmA5tI
hhYh+8ke1uxk51l/YX+3U8fiierlPBRa0RT4n142YU8HGCUAI78lOgmCyL5CoCth
My7c512OheIsmbYaCSQrMeOrO/T60Xo1go0d7gCOIr+vBCAgzXLikQ3JsiEj3Bkn
pQVtAiq0tPfK2JRGbMjGHUxZ7VDfsrUO4Z+afeXCX3gs7eVDe3DhEtV9055MO0vj
PwPGgsi/GSJNSR/1VlZYn0dnUh/craZOsdZy2AtFs3LTguZ3C+FZtGdBQRsf8xLo
8QfBqCab3KbY6AIGmAEcWpEos1dcGg3warEVWIXpbxUurpnfM31EzPXX1571ZRsG
TmGwOtYXtfk2IIEQccJ6o4yrrEHJGb0kWBVf+ZTsJAtmBCh2T9oSzk9eMOoxRtKk
zICekz/O520mn/tiyYl9G2xP/6Dx/UD7xSs7O5xtthE/yv+vZ3Tia56gPbKSPG5S
Qi5QYDPUSRxyfplLB1xUPM5BMqd/CiSK0Y/Vw2rurE/OjVJy/HMxjanaugpRjf3f
BODFpxKM06MqR6kIpgIpPkQYHWJAyy65b4fZ/VuY6+pySg0+fQX4+k8Fnp1ACq+x
XABHHziadvB3lEIdr98yQz9H81TlYV2pHrWJt5q6GFkFflrsZO6EdTkUTv132ARL
7Ua0pe7bOgPK7Q8L77bBlHd/dfhxCV8/dmTCaTkl6YdJUB6ujjy5DZaK68prMd60
VyeCgRtGgwavt7Dav8Slxda2ppTSnn9gNxCD7riW8ZkFutISSw59VCe+LWQjz2HI
9O2uPhyDObiKTfG8W3TcT0nFoRmUmmAQuehEkBvzGsrxMpWfD3jAS90YC/JiOvno
CTvAgajR0ACmrceFmT2abwY9UNm04lxvwW0e4g3CDLpYWVv+gkxH7eFwJICtRv6H
ONUrpRfsL9dsvB5g5gcv/x/rAMzYp/uG/bEpCr4hJGm6zXM1BF1rB7uwAvqklicB
3LOuL/xfazDqfBEmkUit9eFDlyQIMPMjADN77J3CrpuVhEUH8vFG2VI5/kQ/DIw6
IOtCUYvFDx37DK1LdvW0ZUmq31NV5NTtaYYtXAa5rmgwVI70hn6sYdSQ3VoxXPZW
0ZujWPwefZfZpVnwTUWMTQKcFg7v7JzTYS4eu1z/vL+O+Bh6kfqXx2WWXcaeYuZ1
guaxk+FqhlPaJUr9DGPv43eKA7BonE6yTNX+Lx+CAc3vuQ0x4RYK1QHTKXG9fyVr
cDTmDZYBcpEduOnveVT6GdAHelmN0ihbANwwpis9KLidgRbgLaOXls2YFfWlKp59
7/XIUbzKlco/EUEdTiuN3jjr/qz+khJDqzdnFL5/4JtpzMMizbxPHFMvHP+ORtxZ
yoEHyohNAilwMrizJQ7ukLPtwn4Oyjhdo7QaHjoxf+PhyE1Kpf66Yg1Ly1qEkFNs
S3GHspbQ/bbLaKLK3IpkkS5li2/g5eNSFiGeJavCaFfPeZVdMf2lfLS9hhdJfhsN
LphuVqsK0uMOONUyk1ZlwqZ2ZnDqijINDVxdOElWnqhvJzXUN6yTG+Gg7OkjZzRq
zSoKxUMOiyqav/jnp6ptIpQNCEOq/e1O/q03rnXTz8NRFinDQQIarniQI/tLA1qD
ddk4r3rOZ4cXjuhsGXspMcfQyyj6Xy5nmmI6Y1zY9gh+rf1jPYaKdIis+FkSKV0r
EzDGMW0eVMQ+f8PpkjAeyNQ9xK91l5hQYGp3/CPy3ONdouYcEscmYkBwDBbmxrGR
24a29tGXe1J5s2TJQpeWDwM03f2jXx8QgCoXdx60qcVS7cAhl4OnNdauTuBIiWq2
SFcRwOuq47+MkaLt/kO4SzP0oRi9dQCDENDDURzyJ29XSzNisMDF/sGR7alcdgEE
KO9RvVCPJWVO5VST1ucuPSIJFffLS600gxzc91uqpkUGNQmqluh1ugW/MdiDER1q
bqLxFU1GDNUJdKn35uf0KdoyS4qOTwpIdYAUUnrIs+4X5VUEq9kPgoBWAlBkniCX
RdU26fXciNcRSUFWCnNfJpEIIDTXlSsPWecj/PpQj/TwcAdqDXOY9NWXZlqy2xoD
Xw/6M6jlAVoTGQdZKXDl1r+i6hezE452+oENzrqPGIQmNDgca+1g5BMMtjsURZGp
CRSH0g6XVSieN3A0TcpIauSZ3y1RRxLqX6vevav+msJGae/d/q18VmRZwlRBQalc
rNgIJEqyQ6uHZ6UvdiH052kQ4yXlMdZtm0xRh82m2nrnVL2M8t5PLwisHm9kXcaC
73Z8eYm54NdCxujHIYhj9oQzjYTdxSXKsxnzVXYxuGSI+FfSO63z5ECdlHkbUP1E
LWDQcLmY9Ms0SXwEWgjVGzWUQh5TE8Aiaslizt1JSrPlDbgl1BLARoIXjk9k4Bms
HxxZB6Qn09tTKNlmk65z9yWkVmPSKreQnkOIx/AF65XT+I+2alR3PUMoTF7TZ0Qc
VG+EsDnq4KawcW8KaiQ2AFXTGO57JYLLYxXO/XIdmVv0e56JZszCqZNOMBbaKqBX
4zuoxr09B429KXM3j4z13kuSAzetpDqz84lHkbw/lzmxiSKyVqNb+Puq6MHEXk23
Kr/GzZ/5rXxMzVnZlLHL8WPcrGIO8j/OQHQuyd0PD1NhwM+3eL++th+T4eOZFZAw
r658du9nD1T5eS8jeBwIXCrzZEGGIDAIt4yIdz+d91IfLIh/Yr9kHp+D+TEe0pVM
JpMni2qqcLCjYpsSK3uRPD+HTbCwj1zHj8jrMSMXgt5mSsZ7BJBY40enUcJEbsG8
iKhGcAgMVmurN3TYCM6FZaLO60A1TZXnd3bEvwhWjkomiz6RSaj+pKOvrlQRq3+I
fT58cdxo1ZlQoe7XBRagZ6KSg6RFAGhwKTK5dyVpVlsHxwBB9vamwmSOlithDsDu
N4pgQ0xjaLQPTUk8t39NIt+J/mL7O5Lc+Iu/7PY+pQYVLkVgEHJC9En4WI0XXOXF
SbB+UR5otXxhwcDYzOSmSNVnNn4Z2fe1D+puc3rlBPKmUpZHvG/hmBHawp9JTqpX
n1RdN+vVqxdd4xiIrTXQmau5Z0T+ISNax57sre9RD/PaZ0GPdOX1hC3p1lVGQBjx
Y7oPEAPIyZu++JbP33L9SsfLTj0/5bVOg2GuPO/36sIGuE/Apae0/GzULWq+zqw9
Mo65i2A7bmIfo+qAzIJyxVYElEoE/1bvIbdxZU3RIFKViXBS0pKcvRcGn21SrzBD
A6qxixkWgjOIQFqvvLqcZlJ8ca/5hKZKmwU43peUolcUogKdH5AJkQdyKk0S+QKS
3wsQ+fHIOGskK0rg7xsgsBmSLvnpApK54TiIgd/fhxjRUW+OHGV2w7Y2YssXoPOT
uPv3brEUUetUAOlWM82xHUSXpROFq2ZiyvrgwVN6yVT+8ia323zc0npG55ndaqGM
pEss2TaaHWAfCEyog1uujb9wmlZ2aJ2rfLxnRWyrgpZh5ygefMJbqcWXf8Y5adzz
AAmRP8rVqqNUwyhs+QVD8jxiWjvc4+JtelQ51EnAOhMjgk4z0LHYufJXPwW/YKi7
atHbONlemtITT9uS09HixjR1t1E1n7ka8+XxF4gjpC2bder5v1cEb9rCrEwVsue7
88n4BnDWiEE1vvDc796Z4EwUp56qqpKZCbL+FOLJVru3rI4ltxq+G9syxbrIDday
ywtddryRs4v9xAgxTOgCUpLYy9Nh6Nk+3cyzTZDIGhQrnfuPtYFsPI/HUQg/Ro3Y
PO6EoJXjnD7U3toBANLJgLj0UyH6bx0LtQLlcgxTHNlUibDfoQx0UgDtBCFEoSlY
arffe4hTW526pFnEcTGqmqZBaM+9zfeY5vG72ynAZ+6RTDUGvOHsH4soiLozwvzf
UUlTv+UyFQ5/61bu9XKFtUHn92Zvg0CzCr14LvYUxQXu80XIKHE5H0/akB/GRzY7
rQRocLYaHm6N9XbmyBhEdlVWgmlZBiuSb89Bbbnr7B7sDq7A5URMUedlEeE/KuMd
VW8p3ShR923KTsA2mOn3ZRRmrZxlnFR/lQVwBo6F3WII1DmyG9vAhV6HhnDr9jgD
KyWGRFCEjPBOz7WZlAoWCbqBHhEo6OYp9GDtJF6SRbqgNtQKzddR/zvOtyUPgwsg
dd7vPAln2qmvvJ7/LrulSVJ4cs1UMzZTloCtIdBp8g7JMK0tOJqZFHQ6Oyr+FN3s
Pt3bCt39taAsyEana54BLhqDd1CCLXzlDAQFFiI7KSp8wtv2nv+c5Z2yIbOuRCtz
FJQ9K4IZEzNFjPv/8t4LOUdN0UMDVZnjYll6c8Kw0dZJu8o99qKNAkbs3ss94igJ
Nb4d/CyZ2Q0lj2z/J9Bm1n+OXLLjCPN82P5bEZtqpefGQhmYIMS79A0N6PWsThJf
jH6Rgq9ktZ24o7plDINVnTVg0slWo++tSuPRN5HNFIgMg//sl19QLhkelcGF0KXu
F7NymBwSIaTSFRGnblXzOGiw7CoprJ+OcB5FOHIKByGM90rhXl9KwcVdSGYPx0cc
R+24n4OZku64zVqj4YxhkcIFH7f9AR4j/ElJPZD82UW1jqpHXUdQQTRhGEdahOGm
+wU8vB6PTvfDW2sKGegcQW4DaJm18/p/EruFcqqCrGxQzms+bQzHl80ckqCpmlaa
QMnkLbDbCKGpV5a22dCi+J49HY9l0EbH2UTuePeeDbAejWeruG5Bnk9SyR5j6kaK
JS2TEwhUvDjbY+bS86Yn9TzC7dOTOQaTYhfAKEPRbnGvxONABTP75b1F/K9W5Eo4
9y4VDTQ45WmOl+AvZH8IYXM0avva+15CG2CmJmGAjnZhFHQP+But7i8VFBvib73u
Vx4qHDdV1WWEx95pDuJTL5aJTj9Tx0TAeUKo32ZJV0AMFCCcSryljLjTtrupLXBp
y0reRjoQLWHG7Hqgb5PDoWQe4iAsHDjJrTSEZcHBBpMorE2VaZGlhTr2qx7RIR+S
wGmUFWzgLX2yXgGgf6aNG4cRPIstFtw+PiWCEpJzojskViex+4eEukBstGBJSdym
E5s/4BgaC63sdiP8Ty0xwrx88rDeDT8Qj4P1WeSY2GHOY2ElxdiilFk/9ENERtyA
zPk1B71mjUV9A0lgo5WceBGuFqf9R89asQV0q3RPk+VrSTh37+LyM7cMfVc7RsyD
MPgYWoVRq6zKn/jttdYa68wwjdXO7CDuKcd28Nkmy1vER5BrO57Hs6zm06fe7+c4
hxKvuLi+MOGYd08MoMRbygBfH45ijewI6WOJvF0zwYPpMhY4LJaw1IkUUoa8SgYG
k1P15cE9mfGm3EaDmrkVRQoy6P6zw3Re3mRuJuY7jY8b4LI6iVYP2ihTEKqVCyqB
R1iSeaDVSxVMOWK26JjuXfVK05384G8oO6SoxNB1MG1sX3a22tyrtdWGTvdw7dtb
E6845xh3AU3Tt9RY381c2cYJnmIwBCImUnzli3dnpSMWB7ncLv+AQaCGvBQMMTwd
So9JUza9eplvkoHbTN5f1Br112QuuRH7K1vFVLauRPzx2dHsfTOJGnrZs6mRmSyB
+G+zJrZ1ewJ3u2+R/AaUUDMRpolTIfqrxD3DHZy6JBlCdniUFSe3Knb6xKcWFD2w
Tg81ZlFre87DpdpN7g4ZOCoauhfGbjYy2oLZGjSQX5DaWQAmv1Xx+oLFaO9hvLp4
oV21A6dLCKBCMHgcSNfQM6DX+0Fal6yOvPKAR0V1tRFTEPZE+8KCpWGXkG2KDxNo
7Eg4xrKCiyvZM9UH1s07bFxD3JApVyY2QQKU470e6Ew8mnmk1QEXc1HpvK5AiWjK
HyDeqrcobmyMGIC3Ggx9iSM4O/i9G85tKFcZgSNEMDcM3biXaPosRzkmXPVTmOUV
czDjuRKM3w2nOvgoNXXoYmOaF2lBfaRkye7oTosgNEhy4Pl1YirT2rRdC+X0UOcl
EBG2EecaYjO3jCC4MDDEileMpcwk20ieh4O67j5YJRkRF8yOG31kL29344/SDblw
O9xtqX2waNARIDElSnvkJleNyGu34ToYQ2Gzqx243ksq0wNh2nb9522E8RDizwKA
VRlgmX2mPHA4+kUaJKJgZhpXzqZQGMntn+usqAE8AQ7POZL5GC3RoYK5J0Rx3XXh
+idQgXDx3dHzFrfLJaXFotYrpyKVJnQ/cEDbpys31uSurFoeut1yaJZaLoRAGwng
focRlXSLSxFTB+mRIRhdT4Ufn/q5gPQo58X6Fs/wXJPd2tXKg/6zJI4rXQ+Ujniw
GXjyNfQxw1s1YgypnjkUVaIABcI0H5xrtyjigArNaESsJDBLUlFs8hWWQJnz2b8X
B+LAGnPJUzyVj1yQmKYUFyJhwEYEnQ4/BOaPCJWe7+i9nUq7pJwWCizCDNQAHEJJ
KoGkr09PTF7EptFFYn5oZcrhGELuQ3DkcwJ/vqeowOCg28RpS4in8JT3vgpkvCyr
Ik1ZUt6pdoum4DlbGXqb4bz0WJNOiLyQsSUl8fX+mIva7ZkIcl6w4hfniC28NfDG
zy/ZCeSr8FoU+eaT0lMAbYK+lKKru+h6PVzGP/lA2KzkRKc4xUFGdn4hjHYfJuGV
g3XfL+ef7Qq+y1DTj2E/qg+bTVaqaDJjAC/mmJTAdkVWqqduUjS8z2iHaMNohnsZ
H/E2awbKc98uDMD5Bwlm6dI6LuIEnVAoQ4wQ0PnzqFpMDUqCuVo4jQLjrP3+waNC
RFIvi3Q+TKrY5139dEKbqUg2R+jJwNnzqQP06i49HV2qcDS8njuVrAoFtceAkhpm
u3PZ4z0uQA2v8pWLe2/JrsITj53RxchBELClBeHY/9crJ0BC4rGFymJNBprk93y2
Z48wsk935h7N10IKT5o1/PDp+VCMV3vtvtudfVW6i7Rt2l1lXxrCVczggmJOccZI
p/lgHVpMHlDCuoA381wIcTVOohaJkQwpChBtAh10TTG+kFZyqqrle3swur/I4Wd4
YQA/pTBf9MDku9FzjDV4+H18xvpFbHfBVlwoaKRsC7dPXHfWtkQD9chx3fWxrfC6
q1U2OZCuxj+gqQpl94woKBm9ddjiLbh6/qFiD9tkmYK6WoI16aiS1RUYP2hQhydU
lWRBZheR0vcJpquYL/H0j94Gkw5TljnSukwkFW/pGbsso4KQPA5ePWZgKL5PYatk
oP/dR+83DyQlCLeLkqR7oX5u51a/x6OQo5YW8c3Gp2MjMkcQDU1UnW+BUrzEfhvi
f8DOiJC7G7jQBeCNdEPIWE46cSFdFyClXqzbpXeWp2Z/AqZDPWZoqjl9BikyR8L3
v/dUGok91AR8slnNh+Y0N4r+GAyeNsjbP9JvAkic/B7oXk+t3daA1oG81N7HkO7T
CxegYh4mpNw3Sh6FK7ohWvpYQ7+chQmWFcoP7qWqX5ys6DIlWs2CrwcdiIMQFR6D
a5FrI711+wSUD6jVdHPOTB5jgkn/KxO5Pn0VtGH/c6IdSgakJeCsoLi2InMzrse4
yikor/LjrPo4EZik0LUOgkGOiuebveKCi3ExvDvsiuiqLg85XOHUo2loGo4CSXiJ
pmPu6OEtqVk9rYjLz90Zc0+vhnDYZ62Lmfzys8sxJsFuY5Z+jhEydlE2pFc0pDtU
9KVgdVVmEVLKcMTgUj8GFHa7JLus3tsNJXB/cCN5yxYhhsNjPIBZBi/UpP0MYnyM
bWcMDlHuMtAwUaRpDIBp+tmlx6QD5W40SqRgjVaNARcI5uZywXmccwyxT+JypYRM
185AYYZcPQUoaWny0fZksmuAhAilrE4JW1oppdMm800t2s8ZWyhefU2LPTw+Edad
1Q2xgNVoo/ou44AKRUw9Da8FIk8lEps8Nixa4PIRcRFjPhNvDzX6BXorU65O/9ua
vYfzA44EGHUcdw4iewGhkefoeBh3aBj3oEuimdi7ylMJMz3uApHIQDdhQwd1q5Ye
zLznYqAknv01cb9mVeuL8k7gPo80MQjfhiHIcyh+g9PZUiTKlTFxTKry+2Nik6ND
lIKGXj2X5Ja3Bo8Za7ZFgZrNJFXE46bZzUhHOiisMRjxSqFTf6bQYD6yJgDreYeK
GVcPpL6GTUTWdTzGIkN9i5t37GrUWEdG4u7Iz9/goo4W5QhDu+dQtHMVaI4nK82R
FvfqLhrXqmRf7nEOH8kG8WESRLsp2L9tcldzrY0xYikGrw71tFHV3B4+AFbQ13no
iYIeOHCc6Qfly9l8GRb5DAv236KjUOQ3a/DnzC2p4I75kbudlpn0iGQdgyUHJuwN
AZYNBweOyEP1QVs+UHYoKTwaZxWxcoywM0OsHE/T/liW4aAcvs7Zkic7Zvq1uYVx
awQ6s7thgIuvyg9mLOQwFkIAUD6UT0MvzY2zj4ekX3k2oji+iSQ8/njdk7WQJbRB
8ILe+/sYMGNQ1f8jJAV9ZDJo5RxLeYZNnzKOHkhEcTbXOFeQeYWg3+lXfyM2R7Ui
X6K7S4KMbr6DIAnwkQhqApj5X1J+lUying0r7IzjRshk+PNObzLHmUvigvjYFRA5
tkX5WPaPqklnzDVcgpsdPk8Ik58dZNF3VbnjtYo63DXCzgbPZCzVZvcW+pSAXM0x
hdzf28lyLkOFW9kXAX5gOTCB94tc3BtTK/dNvzpvbNcOwlb+maSnsRH0A6hMntht
wI2gtQdfGNvUbb0CGMXrxu/l5zzG8wR9nW+2ErqsqjOwuqH80R3LTPBpL+5H+W4j
KyNHn1Gz/f/rVtTqBaBAy5jQZcRtetfX7sjEjsw+2D+BnD8WLJ52Z816r40NTDDq
mJsg4S4ehpVT961Uqm32XilaoU+d2ykGG4zJrRzKDZsQF+pWfSTn+ifVe1XEN3pn
i5AqJ4+Vgh2tguPNT4fxv9kXth99f4GL6PcCikYF4eHZjYiH3LKpg+z56itINtMX
RZWkWXKnW4Mjyc6QeqSo2e9i0LZxIfG5H63umZsRvrcacUVdUa5wXGaygHAneqJh
6M4vvhReTLUmOYYttdZtpeKv1yn5JgGH8cYc1/MuRlceFYUKCO4Rtg6yZnvxTv9f
Llo/wUln35PNnh1hOXcgQQuSv/5+nr1gYBe48+/mxOCrjy4GJANHG5p9MER7Sab6
R6xL+k/fjlA4cy93pDgWFLXZZT8VjdvLya6Hu61EV5WWtJUWFB3ohuz2Rr/bp7F1
IAbx+VfT+YK/X8UPbGkq4/4G2Upk8rtZpSlfpYrHASnPazNtDM6b7ANBNwkJauTV
AmB/NBlRV4IoJbXIdexkfQE6iIdy6tQ1YGkoKpglvgXc/rDOlj6Rv8zRgtR2HU2j
aoz7MtUOlHCv1IZVJCKBu3HlBYC1wzb/Pv3XLzxmP0+jZfca/qi5d+IbNHAus/Ru
mTOCQBwpXpqyYEZ02gL0sMTYA+Ltgh0zWGBtzgEk884lFbEt5p3bfGiG0PEVBAju
rYj7+iFQSV2q4BlvndtLG2mHR86bULj+q191SVe27IITHU2mOHv3X9mNAM7U7scp
K21wsCnBcHYgu1u4yO2iGh+r0TiHGctOtCMlUgBcqBQHJYjmdJvgTETjmlrXU21q
b1HC06JWd3KbgKjTEsM9eyvqBdaqNDVfZvcQvWnna3wbPghjV+V2lHPtfzF3MYKf
RWJT0Na55Cn1zTmLLTRbjJ5fUVC5/JrCGxSH+yM81Eb0eCpwsZ5MlTawru58dlTw
OcbnmDNFQK056OIWldzdYsGIzYObRfoxd4Q79nWrD1h6LSCbPF1rmYHoOsk4t8aR
4Om+6yl8vAIAO0FHMK+TpL93iyoLxFYSMx5gdSxSe5VbUN4lFaoFJ6qmAB8PTen1
1rjag27yBzlAntBJEGnAZcWfUey0AI8dm71mpKAQm15L2SGpssJ04i53bBauThSq
qfs/45e52nBiOupdUfZuZX2GWrXlJFRIukYAEtUMZ0JzSdyYRl2gD9THVYh/BuCw
WBUEBZkmoisZrql7RvSEcmuMpGuQQJsG/K9SAoKKTeqRzEtj5Qj2giCkB/fgB5yw
XWCyuu6kmdZ3cWPkAejcsXI+1bbOMhjTxpLWxS+BUn+/UxOUj+mxqP9yJwfQpRir
EKtN1Czuc5KPW7FhwyCLl+TD7cYvkpJj/mevP+rIAu6Bm5dfmr1wkYHo8CyQMO8X
2AqkjmKyy0DpIwzWQRAMv5TSzbFwzECvizIc67H8l++8BcrA7Kg9/jcpBBTO8YRH
KSRrqfmqXZd5AmayNPMfbRPPs32PvGqdow0TXEl4eueF5XO4YdVmZ6owuIFworN7
ZZxx/D7KbSg5OAwMuNa3nNya6WkjBDJQ5kJkyO7Gkay9zzAbidufF7OwE/i7IWhF
b0pbuFFxtehw5/YUpK+5gZ3H89UECQ3S6gCRkoY/ekR9q32WMnPObBsX5pX4BKPu
lTc3DxFPYL10H0yTri4vSgqYl1sAiooOk+5Po3kaqpZyUeLRlPEUf3ZUK6CDaatG
Sx3Km1OvKpeYmFsinxaYndBuQ+HmEUlEpAi8twUsgcR/wIrHUWMGgXn0xNS0zYMv
C43+IclVZXfFElNEU6ytazVh6uPGnUEockbPl8Vu9Zso/C/0kPzG1RZHwX+CA4/b
b4gOYB23/4/X8sRtxmLX1NpCoSnguc5FP4javNSiafqveDIb4oOEQTv9NOAps+y8
tk6fEw/fw7HNnnsir7CirnquMUEF+XTbzUxztS6iLIZsV0Kgawe+xQ2jc5Pr5PC/
9cxQLMZbOolIZjvwFGfzQAHf04SiNG2jzD03nRBXa4F0XSSc2K+1ju6OERDxQLoX
qvbDU7lgw9qvybDZ+A1vhgW3TJANEqlUL7KXfIEcm3KGsA9bVE99UjDgKZYHOz8f
OG9C/2QMCez9Y3ysr0MRvIvkTrFOxzns6vyl5mHD8jb0CL+UjuhMJ5WTc9umGPjH
nfWN3jiQX5dwybWVjKLSaUYqna0Qc8xMrbz+7HpwFr+1rPBudmaU9oP7ZQNfKHU5
XyhdktrD7nBzbOrNXG+VUxkseMCJX/BhBVRizFgHAkxSyGGO0saotmcHFHg1gu8k
KtRhi7uwPph7MHsmy/TLvP/A0/oGqrV1WgOfftZULhkUdspBK1casEWg4k6X8A1G
4C3gnknJNtCubpd9qViTP/Rr2YBFiy19C3g9aJE0+dov21IlQ4gpQJElMTcg06kF
nrSzCFLjdgkwnhxUMR73j4UPVXVniygfB+582vbC2CrGt/cHM41UiXdHi/ugzgIa
2EBzAyUZ5pTJpqUWsVKfvEAXw3E2B32ds8Qse2EzU4OcrBXrfCBDNGf2KGQgNYGg
Pmhh9iuChTxU6DNUEN51FooLZ+8dIVVkZTxRIBzNYRieGyl4m7IWt/Wrw6hbG83D
g3+9EJuGLBx1VfgDWq9rib2Yn4n4m6PLNWsRuQgHfYQibsGXiVMEMk/FivjYyD75
AiS9Zb/5QEzAFiX+4bBvvSlDyGhOsHIBuAULyvubtfmxMJIsbY7zhRUf/MSJs3T8
3CHSputUVlUaYQcnw4u1fT9NLQH2X8qHvSqFiZzFzLc/7FI9wP6pKF+qE8AbvXrM
+cFc3VCllB2WyZHDj60UOGrA2t2FaPvI2p6TiqQ/CXqYw0rF7DGQgK7qI0dr7JE2
ixBThKgIbXu5dLAAsppZj/0z8mC5ZMHMACAWU3n5rPHbBKxTXEyar8dt+rdPLmvh
ElZRSzdZKtJygM5npMSVbDBDvjk+lTox9ZHE1PWqm0IhYZaDfyUA1cDMw/MYt/Dt
uW1NsGBDqM6muyqL16y2SFedLBZp3MPYlYBXTgvl6OwDd0le9Tx+ZCHaXCFAUMKc
lGWg4S+A3kpyjYToStG41dnq2rEGwC+ysv0DyQv2u7F0dg0seofD7SxUYCKbXJN0
BKZS3kFLhqlJ1C8tS33ir1cFy71YMY+STPCeV8O/Tmlz6WVf6OrXl/woaq7Dtq8F
4UhYygmVB/VCMmD8ZbTV8qoDsSxUvYqdD9gF3600G1WN9vcPrILQTYx8Mt8jvSZq
AhClKPDhZ4147Bht25kJqwGmmzmF665qCCQXGI6qFjklF1hCfXqiEwRPCwmeAa8h
t9o4w0D/mHtJnuO1Yl9o5zVhYT2y6eUYZiC0bkTet0/bEjH8dMllO+gmOpIF04k9
2rYlGj+ypKiQTVZidf6ZhuWD6Uv049BV69OL9bUSauaTEBeR9YIw6/CLn3Jh/lHt
mv1s+7otX4pAGvb+7R5xNFDsMOb/8Cd935IjvSNewqVsyPkBUEU6H6pFc/DkG+1C
gvUcvrJ8fMEpDv62YMS8NcsdzkbG9vcCJ3hZmd5QyhhidXCiSItKWlqDuoE3+2al
3Tdambzoi9NTGoYCb6QvxAU7WLdoA7RsKJLIu9lJy4AvGw0Z7nHFyQ7/B3D/iZzl
KOm2kmMbzGhczhBhK0AnlHxnV0FXlcliiqztMYuHtD5crHyeOawn3WELrKUhHKxh
/fjRO3s1fzpPIAw5WTqWw4Igvr1A3GfLHKeu8LCmOYh4HcMQe6zuz5ur9D3wEeyr
On2lLe3LBBrwzDPNjpy889+VFcGMM6ukOgwT7KRYpIjtGNY6g/ppCGcu4y8giMWl
8odrHN8wzOIbnx7owCj7c22LFCjwXB6+75HI4eHIzHkIftw2ed/6QASIF9nOm8aH
9/KoPS1zotlEObm20Wbmw0JNGe8cWzjEJfPU+kjs9D7o4QVxNdQajWPqWdrKgiCR
uHLkW38eEshfnUh67V5gEMfkMAQN9DepX+pDXaJP+vnX2pGrSQbmCFWo6lmFKvKT
Mxh8FHmMMhQOHs9xlsaNvuT96Rv/gV0UcQ/t2iIvF+OYqWB+23v9xu8NFT6vpDIf
hP5pYYmet9aZ0dxfORnjzogDaQFVi9rdw3xnozzC5Ou3aCaR2tA+CZIGaQaRg0aA
aSDPpDYDPNNSTCMZkmaLMossu3Do7Ub4fZlFVlNLB6fl/ia70Z1rB+8ErLZTA2BF
6TI6RCBDI1cBoV/F2uRj2+xxtIOtqRC8dzs3xP5COEpl8ds5Ne8zncb7UDqRbTVh
CQcQhOKjJpRuY/D4+a+40wIqrhCz4prn0z3we8gklljQU+5DJH9nNZVCP3QNLDZb
GAq8FbW/TxZuQ6jmwSRY/PkPCDzYLti76JaVoQMPg7F2GwndXnLLgaooqnIp9fXi
3Sdhxi1NveXg76zUktD7+aIGfFBHwsTRrAM4C25mJFrhpq9dEegS8bNquQQKdbwQ
Tf97HtpEXOvMaO9JpK/ydGsY/KsF9Hjg4+iPWiDYBGype7sZXFWlye3+fRVP+RB0
jDXYWI7ED/RUwwOA/lyQgT3AKciRcRnIg+8qdyPnQpvpTkxeBHZB5dIFFbazMjNk
+mPwJ/zyyEp8C1nCdlUe/LxxbXL7Ib6wRhRffXslINhC1dAjRpGGFgR1IsslMpVp
sH4FSYoY7QN/hL4eE9JR2dOBoJQCnVV0wzcwzwTK64oT7qSKW8vLxgHZFF4mc/fr
wL5K+njzRcOWzMGW8KzXU50TrtgEbExTho7gyu3JwbsOJmtrNoy8SFQo+p5aM1sE
s3/9DOjGuTkovZtlUEB8Zoq2BzGzIK+nc3MkuFUxCKtHgZI2qaxtgPkRZcvTAlng
orBLORtskjFSa1MScQI1rtGUaK9fLTmGyREakv+htPrxZIpqADgj2qK30MYy8OKG
M8i6cMNpvlgl/I3Hr9P6t+VnsN63mcfBjSXDklrSoSzMrvF++ahPNcQQqbKP8jvp
AVJABs6uwT0V0jPPOI2wosQ8NyS1G51ioKK7uAv6AozKnzq6osqcGJGqXPO+j9c5
Ncmp1oIRicQOMkg+gUI2pBZ52iLVoMr67tpz8HA9+jRDDmlx61cfpzaC9z/LatOS
dDzDQ/6hT94pG9zjsuOzYCDFLiBKkqURzIiU1nIq+sxQepxtYxqhpuLXpkgT9r7d
s+bfvJGEkILCRe76Ml8W0DsAPytG20ALIM+qaZGXFtUgI60bFWjcN5mh8oBVPip1
np2ZKCwbYJlrdNZbGSaSvqR82kii9Py+n1vgbsmXoEjfVz95uhgjnjSEEKEtfpfv
jLsntcNohXCB4MjrFqXlxaVcaHvUBiDJVReRN7peoTgdmRXfZYcMMaIVx5BBkr0U
qs3o0GhLbWysmF01MjAa5l7gbTLZ37AOJ94DceqVqPAPXltHrPJB/KAsPMY3pEOO
a83weAo67zJV/ekHW+1rFQ==
`pragma protect end_protected
