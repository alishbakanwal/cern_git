// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:02:11 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
TBm4CLcK6oSOCjmA+GuW4UG+I2niuXf94OEYH7P9idEOs1erBgZRV3a9CfKpdGEi
D4yRUzCCqDTZv5ZWUQXiQDIggOLb5cqDG58Di6lrxxvfsV/2B8riWQjfZQVDN7w2
tlAWw9USPh4XT7Sqwykimw3kNqBNxS7LLQlMenwbarg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11648)
Yv5E22YsnShtRJb/PuXvMkeE06pS+dY/6KZBndq6gN2PENfkBaCuT/icH3kU2Z0u
+u6c9ZUaQtBcxiAZ5YcYSNCIoXuOpmxH+Wa+v+2y6CG6nzv9zx85RNZthJlTU7nn
86nsGoFC2ML++OZ4tZMJNTYsmvXNjqvDNBIBxTqMjNA7wn9ChfPEMqPLWNLSfYeT
EckC3GJZe4hci4WLGabkkfgGBp52gsSkPqpyzeExtQZssqKbUk+JwhbBWBqAUu9u
JM45lPY0GO1Ibhgff6zHoC9apNBScEpViRJEb7EA7C75glYAou8OLnVp9m6B46t9
TCmg7OAygiiFRPTfN0kVHEFX27pqP16f7r23/T3ZmZpKKUr2QAqIs+XhMCKKZTp4
8t6PNaty41/6GLhInkikwHpVlgIO7+opzDRaP8mTwmZLzyEzzSbsKg2CGrF80DQq
n8Azy2zZNnitf9hgNzlIxRbnBMNrFv0/bqcVj1Y87vZiNfAffXQRvi4WXQSbaWqg
kcCVI8DkuDFXeR7LFqiXGuzxntgpLTs5slXPVTjoXYFeoB1xvWycGBrOLpQhWVO2
68MXjZTzRr6OK0Nd7C+lKL4/qBNdwJRmUZflzc7zmcuCXRys929LMcavNGW/bv00
gA0QacehNdkq106CcU9/a3yO37WxIPuT3krV1zotgzm3gA2DoKXkgW/dptQxLZmY
R+BusnKVyFeIS7om2u5pZhX0LC/LeoMqNBs7fH+ReoLjfS5so7/ii46hlTDz9wC/
TWf/utig66mprN/Sc52OVQ06Q8Rqg1g+FeuCRbzGCt3FUnQR+nMFtIs5tCAjpC1J
ShKpR6HfBtm3EQNv2zVC4B1Ej4koeoFof6dIvEXV2nsVl5ChilwwYJXielvjAvHr
2yDMF04HWSD0ZRvwBxBcs/k2cxdOj43TNU5DjMHyWMgdigzuLTBS5PbRLDvvEEtH
1OzKMbQNCnll8KBb5T3xz0sHdC+PnKkM2mryK0WUi9Asu8VKTGeXYyOaRvApmnH+
QRqHZPQJXu96yDYNNQFqRrKR8vySakL6VtrQrmrrgSXQNU8j1xVkqYJV5mUXrr5k
A1U2dHejnLge+apgzL9mBjiGq8H4wjUSZefgH4uTor4xEZRwk+S4zz+q3+XyNNuv
xTsZeeiarpJVHKdtRcntYxblatpMtyUKblZMk/WYYEafCT77LW/GIV0vAz0OO0lR
FfLD137Ns6ynGeVIvXXFjjh1Mhy+X9EkTdm8uHo8Qm4nBhGRskfqDeqR27wHOLh2
fS3WzLic/pTrL9CuLyyOF//NKksbX+uwRSMWlfyY/LO3tzXzFBgGJTmEOrP7bsN/
0IG1VJPj8Xj0NA+EkVHyy9HLIT+cWCqAW8YY7XYSnaz60Wzn2632c09ZU7LMRRuJ
M9QW6d5cNaqhsqIG66SFqendj5ZCBATnDLRZjcBbJVn7bVQqVweJbvIvt2egjpZW
W6xXBjzcde3zV4aLZ8Kkxn026FXBDBGUj2qgovLH2bKUpPX/EnLHhGqNhhE6jJ2k
5FvwiJKnrGfKmBvxTAF9Mq+I3g1XY29SUZXSD1u+CSbXbnvis/cIFD7FCnFjAinO
Lc3nou4KS96i7mJczgkmi1vPWWPglwwgiMhzDfNmazM9btK5to2JbOAYq+THG81L
ZVWrj1lYTjfd+IhjD0KH1VUi61i9DjAs+jyvenWeHdCHgnskmH0Wvfv2ocwscR8t
zxpDgRtr2TSNiOP5GMgzDkn6KkN8fpPV1sQ1j4K0cESfj6jxxK4SVsDcjJiIue/s
Lh41GZvuBm7gz8C06/aoCQ8oLRlzBpoWMfs2/W/RtkbR0PNeANCy4djU7wlzeE2Y
EoYy+6i8AXkbadsfA7vosp600t7GtopspMPagG+lhZyw9Bd4NPrlBYFrTFcG8k3g
5cx9pG4yuDfzuYiaFHBhvxg/YS7dhBEgEKC+BfosMEn/NfdNVRypdYrEv89Re2/V
eJF7rPZeANxyoPhYk5Xq3hW9UYEkNNtq6+5hhtDWmsABzoq3fG/yycWhX6m0bwSA
xH0HIwMCZI3rFvgHwsDMhMSfPVUAwnqmXJ0gntrT1f6BnL+nqnGQprm2uBR/3anQ
I/zd67Ok3urpNL9LVLn4tH5VPDeheTQMN87++G9v65MY779THTmy870SQWjjqo4v
SJ1RyTrcr8XJSq9KCXz/3oTnPbaHwpK5b8gK9tRCXVKs/vdxzbovEn6bkxS4xfV9
4BNN9zl27+BKnmlZcwjG3po1zSaDnm2Defi/G0beDiyhC9mh2KFT7csbH4ICCdac
pQqbAdUIpqXsLu0GvlwmG2Wa07sbl/38RdTENETnwpytGSSE6KSXnwWeOapd0+XG
sdcelGFAiooz423xtldQEzrVqdYXP2dcsqWhuR0vKWHONDxUSUbClx464zxh+gdy
xF3l5kkXyf2ZiudJIrAz19p5cBbIko0A7e5opod46SRT2ez/2C3yEyECTByajoPY
PfkDwNnduYxhd4Mys+/UEMa537dinD46iXU1QWKg583id0r/AUqd6McxS6EjtRw2
pwOylQFDKa+cGFPcDZp4kOBQTEIqeDcmqqae1V0E/E8FLO1AwW6VidMOot28opG8
zykP0NEUGOsFNKsHPpPwGCdBnI0P/jR+W6hcAFUbVcpMDg1dOR+6ZpcwmSXNxejv
8d1WJyfBGgPA4X4BTzy72/5QyfJfrEdWGutewicR7NNLQojoP6FuIUCsMBrze7r0
LruH4TSzEPIVMUjskCuRiYjG1/qXY1CTjQ1kgYkmXlssI0LE1jaDVN5GbLSXlA9A
XpeFBU1Don7OlzKgsViv8lpeqVd7cSMK+R71WUlqAfjpmanNXClxqNHdi34udiUx
GKI1HPcQO8KKl3JRua8avBcMS4Jfl3le73BF3gRaN/jaB6VDsReK6PAe+sMzoFEr
4Mx1zRsqnxgSKX51lxfnwjCZ+v8Hv4G3FBlgSF/YCrMQfnfiHWiJjLM+UMg9Eum9
85eBZnf0hiMXtIwOlJfv2mLR1SGggf4i3Wxpa972WoDbXABWhZ/VjltKAWHAKnzU
BY/FID8zXJtxJ2lMtkTcmW1KqGqK4kpfpB4oycWrlae3iUhgOB6hwPEjopY9Xk0T
Sdgr0LBTJpLzHw59SscAusMpv/YQrUEw6p3mzQN7z8M2bg6g1LhOZepKqcGwiJ2K
1ZpfCJOXIEGnY+aVsUpT+efXk/YuBAmBJ2Cvpyco5X4PbPM3NgXun7TUZN24tAMo
/keHWFBsgtOfrR8Vi525+sIv9Mf1mBfpb0O36BCxn94KkECnqauAz4Jrm0CVm6wO
ay34SZUy1yhFT08h3Sp9QsvR3DMWyojZhQEvD6IFaAm8CyC8+o4n5GxcUXmjBsjV
sKUewLXrwMuCndmyB6BW66BT0J7KAhVllw70E+r6O8PIbbrcAVRsfxykD3D07UkU
vWYE8oBW5Yu3fVlTzJ9vloTk3jYAynAmFWmNz1BmBU/B3refgCpTA32YmS/25olP
1JYJFdpC379D68IZYNQrWRCTFjCbm/Px/PkMo+EiNnG6+HxRv3EmhofNcTEsR2jO
b1k6aL9E1Nyy0qm4CjI48/LqEzJgEsWtrnzTEVGk89VmBOjpKWYF37SSmFX9agxk
RGrcaUBCfNiQ0Jx1FY++WviZ15SeWavaFj81qqScK1cqmhFpR6jzMBNZL4+Rmz/A
Ou8xl/xwQmKHPgJt+00r8iTq792IJM4WrG2MilErDSUWHvMefSzCFstwtBhD+8gC
DXXOB2aHZic3BuExQWeyCCFbe0+aivt/eeta/LZLEgSO5ccQn4T13qpHsGZAqDfJ
NPAPIHkD9N9ape2xvq2+/kkbV692zhod5/sHYsun9wc9zfZ77rQelmQAp/DrTXSE
9rVbWsGX9xhQK1QabL+JHGljCTxlqb7b8yCJ9jhlWRAI0czJ3oVLCiyAkWaGiVbh
onK6uGR1lgx/988yzx2Nou3xuSxbR8BoJMPps/U7VWrrz+hyS7K0q/I12O54iito
26g7/ZjTb40gz/qQ5y/IxVbjCOdCIzVatbSHQsXHY3hs4rxQFw2LQux8sOjows/6
AkE3/ABQn/n5KERASaccTmtUCUdffrV2jOVJS8ApiqSOdcE2wLX+SlbcXQUvGA3m
ocDyzvru/IV2AwmMeBaPxdp9pJ634PmyQ8U6Dmspxu/axr4u1JTu6FGW6H6rB6l4
2cDYOEmkhRG22z8QcXlsDUCnW0FVlFmgMuRntKVERLp5YSrbNd284ZU2atbUXcoW
ihZ5j5nF4DkZA16WcAkl79wk1R7IGcGD536O6R+niYPTUxeu26Vm0t8u4z5svJ+8
fCaTqJBBVDxI2aOe7TT3tc1jNWQcfEFFVv712B+AJNsIX2/3FVjh7Nh1INLNjmhf
Pko4rDBGbT/jRQ/y8/Zcw+7DfKkIeS2BWo6w7zo1U4HF6JFwQmLhNj7IfnYlsOPd
6xuvvDrgUavxGVTTOkafN+f8Clh34qJS/KNxju4E/tK6h74gsfGQnlXwunX+Jg+8
V+sCj5RLwXn9vRJccuMqkCfieOO2Q2aFaYTcmtSI9k4DsTqE1OspyHkT6AgVvjht
BLpywb5LeqRKlOi0esAJe7XitgKSC7iNJX5iKCIKT93LncmmE7w0jGB9MmBTvoE9
Y7t8G1MBOr83OuRMR0JqUAJheDCnWwU3XxtF+88jpVvLRPjiEHZahv62cIlVLuTc
QB661MXBQGDYcyhUBM+LZb9fpsm5PU9j9UDqXCNOMtX+AcY7vhrTGGiKUZBF8QDm
mtcimwgToq4Vq/lIwHO2JgT6X3muJ9rQQ/pcyI0p4EHGy9NOp9xa7Qu4n4f+CkhL
i/ijk8kTle+iLJ0BdRg6fOrwAL8dBMzPWaNM81RrrUz5ldV9sBwaZsZwrefTrWcZ
Yl8El11YYHMI8gqdxuNzQpItEpzYaibjesr3d+AfepujIstbZb5w3YEuX0DCq23O
YirVgOMyfXKBKjVTzxAz8y31pbN/BUDQnt+29Fomcr3C6GvYEMtfecl0hGuGMhx3
RxLdcldKbRLBlD4+goXaF5wWWPjblWejSZ4G0RMiBspCNVVBgm07wLGW7t8hO4IK
NonTiYDaE+XktHXjov93cYzr+2+4Fn14QvoIaz6hH1OWZvpNakfa/sMUwksUVfCX
lVaG8r8L60VdZGQOBs6YJQJWv4+ME4am96cdJetSHz34jXhWEQ6gKT8Uwe2uLNKZ
qXp7SmdneOEdPvDqUFqtu1G9XM3jitSaS1ozOxhGfIzEsdAHc/ALvAzNXlEE2Xny
hnJv336SVgAblKyA89UCoo1h0BWmKtTkVcFwm5/jDKJ7Sf8T0QEl9LNkPJkJ1e6T
won0poFYzXf579puLXTvdnYeCTzTN/bQU7e5HzvjT7FABUlmgMuad4PolChdLc2/
CANnueRdm9j1jA+bB0rXdcOPeS47wpA2uCoouA91+krrLGpxRu4sEbjlYQv+59wy
1IF5CjN0wzvN+r8JKb/pBlfT/RYR/h9ru8jyps148pyC3evREYAsLGGYGB6LyMiz
LFuUBixoSK5bqqWshBd1+uJ/Vpl+GgSFEm52UjpYgVmGMM12bImv7s5uTJUuiX0X
gVMuknqCM1MeKy1OdEF9dBN7kVYlIdYX7xOh5c8MCAGz/2sI1NqfJrGTiu8pHp4P
97QWVAMfjvHTXgznZpLfmbbxt5JuvdGkxfPyZmZYTsc3vuW1pRL6j4wXNeo+7FIL
D+BRO1+VQ5i1tucotiMJ0A9D0Kg4Fqy0canJEW8fbzguhSguPX6l3/BKlEkyCrHG
Ndy83sL1k/q8r+veuZQ1/Y+ib04bf+BfKQdFALZCafrGp0pcaiTF8wNs1x6AM3rN
KFp51bj2FBLDvPedlc3Vk0i66u0YqcvfN2Fy2OyDARgJ8d0vOUIkCyEutGBOqYAa
gib7lmIg3kxfgU5OLyw5lPJKStcrwJqZFhxC67XcjozAZwBNNoPzwjhfMeFzBfN7
UQcxsdmBM1m3vm1747Zs8RIJXH0CviXenbXRn+43o3xZ7f75q47CdzJyfn28s7OR
d882NRprNVvMLDiWZztfeC+jE1y4UGroIfBDeYcMBZYh+t/tPR5wNRQ6RX/8DdWZ
fi+zQUe4+cqUJW5/t5DKWCSKALN8yO4yT4TLVlFRUujAw6HeMTNJBy1e4qc8dZBq
BD+ROgjMmt4J5t+nNMrBtuYa3oaKSHWWoCbgKwAKNGRvql2VFJ+wZFtLrr+w3nUf
0WO05GVFG1EW8zfO2VKgwUVwxT76QQuZN/FnvG9lFqywUGs2VtBn5aG7+mF0dSmm
et97SQao4G1eFV0+bw4KnWPtlmNusbKpiAIeatY486ER4cXTfHMXezxsiqkmMERu
GTc1exH6WkpBRwF2nKD8g2NQRRRLhlLpXNrQvqy5hceWvWCuxWfHSl1CUFPzMrT4
UU2JchKeFzTj/7gqnxqxhSBtwsiFBIevca/RUpSmIavUusIdKoW0hzjaJr2aION+
PXWsg1d+Hg52pA4XfT9K5U2MXFI1xi+ERo0Hdg14l7TXo6gSxBpwq20NIEwsoWHm
F/gOmPI2CEkBIL89s5WaDLoaQFubSCr9zth0Wvbqrh5EYRVNktzwPoO9WAKVnXb/
lbcTHR1BBqVXxhwM1FKMu4NcFzANuCmlSJJMEg+r3GlDFSZTFa43gfdU8XTEHbKf
k+XVqfVk9WEBDD0dajnIyGA2FJgVBLIiVaKd8vhjqLAaMVmGFOGfZGBl7QyHRSgc
L0IiVwVMJYG8x7WlF+4xWg9EWwl8HJttr9yRWoEyK3zZqRjsFUW9XkWkuEnCSwVc
cn5wVAnLWFYnDNK8LoJmlSDGpH0by1wuiiX13IMRfRPRqrbqLdRGSYPA9tvaL4Nz
dDNHQ1JP/A2f0U7dMNYxXoVXiLCXsZWzpSrY3jaSKWVBV0BEuifCp0PFEs0NVIkb
eFSTgkVs8u/p5TE3maqx9DkTYhhM+/epi5Ia8p65sqGWynoclOfpLd89xm5ZdMoT
lRoyP46ld550bhDgZGLVnp9yJEQOyea8ZR8N2wvH9i/+31/SKLSWl0PNVrPPFoLb
F0iJr5dXjvI1Ir+ce4OTyPZPHsBXq6pFVF2/Hv54h18tBfK3GWZ8uLzjYrFB1qqa
KgMU219Q0afmPY0g8qx3XMVNm8lPOOjMdz4a8OHtmCx9QQ2UPS5S0K5MAETokGDX
0Ugbb54JTRlABLPxNv712mmBn/tHDLDo1kZObjROFIUkXI1Hnmnc3ZlAxXPY27mY
YEiRu0UOoqWCSQreHXi8l3pQ/wgflspj5NaMn65L4vgiUZ5yvwGvS8T/LVw7xA6A
esL4T2kb0VwqIifJdw5lbCtaqZXc9y4R0pwYOKA3KsxAkE4gnGXLofReO+prJqzD
yVFB2uzF33+yaAX5WxbWiPhREcjj79AB2DiXIF67nB2afXJE6gFST9K1HReeCeQU
iM3r4RaaCEpAU+N16Pw4jvcDvoatviWXB4mlpAsyAQhDIvD/G4V2gxUQhTNC4qdn
Ne5jobRT5lz4869yPHUS5VRQsFgFyUe4qMWcrqgw3x4ufYF0jDVGkKeLi7tPUvqo
xp9OBUSoNqay4gpo8K04VjH0KIRBBmG+/XLNp6Gkb9pLNjNwN/R+tGyaxWE1mG+h
m1/WmWkwZzonRKW+ydRJhXZIP5dWCnta3Quuj405YSRPPkdeIj9hHZ+ZqeFhzibn
SVZx6JK6kjqdO7aWkRQO+p0cnEsiGuhGh4C+z/Yv3Tm79KNVvaIBHaXxA9ChZCyv
AJXxujs8Dsf9zNv6QOSRG4QnBbJx4RRaO3e/6+L7mOzZ/QFP7AkWLC2xJA8tZxPu
PVpfEUMxK/fopuGUntFpoht6wNtO78/3FdqWeXg8cCI54hTOpQGVz4xKQshyXKgE
ej3gr7ve2VyLnO87CbRvrL7mLbhOFsfcBKeSMFxx+F0ipg1hwbEKw7XrsrfdVVu8
BQIaBiCY70zLYAsXJgwl40G2oVSnOBJbe64p7TBnvjagerqi9rQCW1tWO8RocTGR
151/5ky2qSF9Bn3mDTlfA1CtILuppukWF/gJ1CMkO1Pm9s7mKz8YIYZgHyQ1d1w4
8p2OsnXKp13/Ka7Hj0RaSOh71Ss8REggL8XCu4DjDeFjI4kfDNkeNF1wGk0IBt0t
BtXJF4E+HA5l/qTPRjcLY0SL41YYQpGL6bbl39N+NOM6AdLjbPGTViq13Vzf+FxH
KQCOvpU5svK2OH2IzRExRT95cnxt4/gSOnp0vjQzaHFf9VvikrsczeM0N8zvo8JS
6pUEYoErLWUmP/YXNv6fYP4480ABDuPpenlbddKuwTHRkygNx8kQxmofGlygQRpr
QpYgC5e5AqMULG2YrE11q+TyZj2U8cZ91iPHJxuuoXXbFJ+Q9vrmqaob82J6VFE+
bB/6O+Uw7iHe/iqh2aiQght9eDhOizUlyhw+oZr+1sYTwwZq6qZXyKMeChGnSzjI
ejhps2jFBU9tR9csOjv8+fJ7M/BFUf193WI78lyuxTMj8BarSMgeFMePmd1Uf0r0
puzpGAuCNzmqOZ0r9m/9meeVVfM77kQc44UDRum3PDNOKA5qlIFD7jIg4erlNJFO
E4e9IC9vkOZWmQtTGsRVEdT2P58+eksUF5AC9xKs3Ze6gcxLM/+hWujBldAeejTj
KBMo/qXb59/bUKoHL41EekYXCA6ayH8Ptm5Bjc5sbpfyayKqKQHFi04XBiErxgeQ
bMquC38i1PAZA8tz6BhP/PmOD1hWyymV4RTXJX9PGdvvKIdy3gTgno6PusBR+Dzg
MyPEyUW2nTxka7l+KZiwz1nCJXHuT8d4/mhWXq2loxNwQ7JqP7xNP/9joLZWe9B/
RdxFY4seglfMPeAqAJt5SPYPHQlUOEHVE6fSNHntYWbDk6mDWxY2A7tspulpbGW3
4eg4XL4jJCN2YExclPod4DSyFyn+xxCTTLaZ/m9pQeYqeVG7xhK15iQEQZ1Xx+hJ
EFAEuSLM4ILxchO29nSgpELUU3LTlWzyBELhQ99wf/ZgQglvTlTPaLAuwb8fuuCx
TPi3wNEtB+5GNvkQ6dUVPZv2+8HfNzAnOllTvAHUnq+bILsojwUnnpy5VCRNaHbw
mtF9pgjR2/7BParJ0s1XIzoMpfOfCeoUht9hjOMX8QNwM60EaTph1FHsvGzUMJfC
DSP1Wi6Jn7Y9gtaExI2VXEOYFskD9fI/x1y6uafs4NU/XoNyja28PdBM2csS1yYj
4ckO/XZYYPUxWZcSh8amuLRDv9LoWWDDnSuKxjhwohdsmTNfv4YoyJ6hvE/S1LSZ
rr9VUhWIP9ydZbylo6l73NhUCTEyu8M5MJ77qepcfP0rHfYFQB7gebF5v9+BWZnW
D4MC9vB4Y5ZFHxYbrZ8yjaEErtNaFw5P2G4KgC9vYkOns/xYUpXed/1C3sW6+rOP
QlU/ZWbKsHfbwxZxi86s1fu/A28wyDdRRMBd59izowTBUzOEgKZ9232QHiL1QASr
YnkThEMpCA0vP9YSJWIs/Y0MA5XDKeI+nAlnjvxj20y0+jM6GOoMtkeuQIueGwKj
vO5dFkg324nTMPYW3hPrnNAA1gkba98pDKF3IcvTNaIIOp77NyTm9tzyl4e1gVPY
qe/7OMjd7BVmyGdpXviPfnDbnXTfEjviqrRQhiR06KSswid8wmhMK5jxO/9HWeWw
ZRaiK43kqyHkYwXdbG3OPcnKXz/a/jvmfbvQ3uKW7bJZNrWSEggyaIBDUdPsP6aP
Sh9Vgo2Uw/J8HhItLNK1jmsvkUl3ieK5QGzR6yWzAPRi14kRrnsrmalLFg1NMfqU
6jShPMbm4GVfyeqoBNziEVuEzX9XCh9nkU6BLWf0facq4WZDOxeHu3SjbdTxG4t3
O2U9N0OwBJvzSvP8PsChwi3PTrm1LfVIS7raGeopFO0IB3qLoFru9jvgkFZ6wyxR
SXO4zPL24m5jgMuKuPliJSZkkh0T0bMlzdOJHnZZNNQeUMP+ItmOyYtXCk/1RNQA
U37MabAiOWJE92CAwZblb9JyLKid/JG7AtdAWs6nHJ0bsEVQGKY/ffbX8OeHtZYQ
IF48xFJMw1DIdF9f3HMy0XULKAjzTfusyr3nd/Ah3fi+YuwKq+Z4JNY4aMmHtOFf
CSX0It77fZAowsgRVikZndQxQdysrlwjiJ40hFSBDEiaqS8vbzYORtq0ncP3rI8S
nSdGdnuezbWe3vxubhjw62cYIXy2HioQ02DV7huA8/mV8iQr3qVXItzveOgadxeu
nurf76BZ94694ogfe62+6ayQm6Jjlc0lw1Fwwfh5+DkxVd49U7OJRMYeedyxYuLK
UBTVs6ui6+ixAL8p6XJIrIZcdM+3G/usm5ePUp+pJJtBts8Hto1f7rCtpjGfKK6B
Gbwg/Agd4iSYxK1LGV8GqKHdNTwjzmXzIIMoiLn14ivPwkK8z4E7sXnYtR/cUoFL
3XY/mzz2vGgLSkbUXPSSKF4X7f6jVvgij1NO0cLbbckynvzW07smUj2lPEuO+5tS
rvxPa6hHu7lXJKjZk1VPjLJmHa7sWXt63FXQVvsozpvTPL5SfD3eBxU4ktUI6Ewz
EhdualJp5xYdwAvnoUfRgaihQgcYKC4h15Z71aOjpk6VYWkDdGFFh6COk27CuLbY
uShgJ17PozNu5hkaJOdvB9cnfeFZL1NuH/9kPB42ONLvnyS895FVO3ujfLeS5uCP
7cEmoQlUCxnyfUhrXz5UYKX22DZQZMXgw8CVKytn3IH0OxkETD7MFMl0twkdsHeM
bqh4gQ+X8Dm5IUp/Lxf/OT2FaFpuVnGlcNK3KI+mGxmWEfNJ72Jdy8/cf0JH8Onp
KPNV2znnsPF1+ebdFP/NwNfpiU+o8crCxB94sNlOWVitmejWz+MKKpSVfxeWUOPW
Ybd12tVdHtEk5n8mzyv5smGj526ps4CVl+wWipCLZFdFIHFdjEQD0ip88oyIZ4sS
oPPLY2L9ltIO0rA0MOhgYqXBVSDg7CE1jPdXAfiYiHD+sofkm6ouCVTLaXPLWeb/
R/TH7FlUCT5HwTX79s7TKyAv1OE9i7FqU7ltsDo1pFE+EcJLP81Z066C4l2mz8dY
75KDjYzJKgZ9neDzrAxGqQEtNXpCcdqEGZS2t5e2ByOLj0gr2FxfX4TWqm86dnqG
gzIGCvqSjgpBHr4OYeDZlfU92c3esDPBTP2gHv2vqC/1KAQm3Ayyfj9SmY6WB1k+
pZ8dw6ecDeKKwo1icVcUAHxi2XyYBtViKh5uAhZbM3PB7siIPcdqF06/IhtFodm2
l2l9Q4+3RV792hTtpOdP9vVfueI1MzZY0zm/jxZwuI/MTld0Ezc0kTrlBg5DEa+m
WCytPO46r59bAHbYHCXSM+snQVHIojFil68SGltN8QPU2KWjBRTVYvPG7+HOb8fb
uLp53xTtqU9zryDB75y3JbEnuiGASAZRw4vMGlMLhOnI4AbPfOcMls+CSStL6ZUW
oD4jBeubOaSL/pHx8eMYjGjmRk4ip0mRQAQJYKylAm4+hFU7n5RlVFv/bpMYeteV
gvFcsG9WWoMTSQs0WLgierXeVKwHs0SIzcZZdE7iX/m9x5CAcHm7gsXQV8qq157D
CcbiQMIcqy1oOfYLSmuHDnCWDYnBllSjiptBEMLtygq+zC1I8aSHpsbvlVWr6a3V
OiEGTns++fOXRfnNJGO0yGHEJk3c7LOpze/o/c3B+cGFyEvqlecfwQn3InSx/UjW
DcOTlkr0YAEwacxoTBJW6ikMMOqXQdvW+cJx/4hVCU1iCVJ5Pb+EX8KueYFpArsY
RTUvzeIdgj+vYwxtBb/eTbQLA+93iaOsgbbsrAfk4koDE0n8+bK04MAyY8h7gant
5ptYnznl9obSNVVzyMzaAeGdx5Sq9vfOvOcgq2y+1gaZ6X35FU4B0kB3ZZST/WHg
iUI0xEV+AYm50utIcFpaLKFdfZSASsR+B3OQ0PMIRxQq4duGnmrC8qFAkLysl6OX
dEjIt+7eiZIXDKcOOu9akkmY2kRMc5HfsN2m4BrmAdAhLYre8J644d1iAWXUNcyL
zheQ/aoBT0ivlnhTbU4oejQjrqmytKqxkfSfDXMmL+3ZdMuafuXXFRnSBtSaeHvN
EQcXU8SfZ44UBWNDy5l9Wy5ipZeh3QtwTYnHDtk2OPS8N0+1VUr1XZR9cc4rckuT
bCATRuy3K/MrZSbzUpRRmz6QE2z9TQ19hfaEm0xB8wiRHcJJKu8zYdI7HwFZfBjv
T+f+Q55lawXzq4qq/BZE9SuHgE0p6hAGyPi5KGGeyhGASpIqHFf3LeJybGA8mXlQ
U75l1+v6XVoflgXFTv5eIGJRcqANXqfi9nlryVWUtZ39jGeVswfA0WT+tBgH0icC
scqKxxsfNATPXja0SXu3gQOAvtN5QbjXJqY/JcyVZAQj17iX7jJwXDTWkLYeJ1OG
OcVoPhEsWBwqzleRkVzI1Vly7VVKOar8xO1RmncLyB68yEXEObHRklLGjYUC4Swg
/7P1KAEOzs7vYCCgyJI2dKsIAPeIc3BwBao4A09ecr4Q8XCfAMkG/8MyNcHbi2Nr
VMxXxwXFC4RlTrxwMMlnZ56hOjXG809alW5dgUtbV4187ABHJRH8kQac1P3R5d+i
myaweB+Lw7V0kjj44SHWiqHNOsdvqmMTyia7VwYQDogh93Wv0IvYYO2OWlbmhVF9
dcSHvM/1LYT9KVCH+Y4DBNfKr3PP9lZNXAbdezwdVtJ/GKT6wX7ZcZmHYfse6oen
G0X3890RjbJY1y/sjvUhSvjV2xrMyTUCD8QM4kJgch/tAI73IfndJmk6wU5I4b65
UkyoMd430S9gndKyu6aOtIdB2pJ+lFNhY6cWlmY9q7Ev6mjVyazfp5SMPVcHEMT9
SGTzyPgLlz9tQXpo7bTtJX9kzM+5coIL4AedSDLiDjnZXKtlqDrPThK6mur/5fsj
1Ndlukyum8rX5lmGv5Kxf4q/V6VMwzuyKdc0bIRwbLv9JOAhAOHVo/q/OQp1fDJZ
qnZzhamvqI/Ghp1VZwXbdUEMZ2nJm3WYHlt9U2nXnhDTHVwvXIwe4yKvfhlPNM71
5nz75JOQQyS9vkwXApXKXGsd/li53Lc8GgbwYpc6mMN8EWQIDuV2etaUdahd3kdQ
fQzqhVlQd4CsGJOUcfk94+Of1VN2OnbI/hALVRSPZHAOeGI4vv20x2LBj3TSHSc+
KMWca/pYj8PELcytQ7g10k8PAQW7iKijuW83XXg5z4+Ch2EvNfJVmHLfs5oMq9Gz
ZIdYd7JAPTpdP8p6H7z+d0xB+fAX1DuFZB83rPH14+FA33h7QE2ziOtkvUtTnTbt
BM5tpNakowgIlvEbtKf2hEEgep0AuBjkPJyX5HJyys1CTLvZjBgFX4stiZyQIS1Z
isv7/4IdWeA2GWU49foLBpk+tIqX6Xf9RJ/LVNi5j953lGMhxQgzVaRr0DqGUaKJ
o72yTDvoGNZtiCjruhqCXaYF975jwYQUbfMr8d3wgzzy5VMIIpHnusyhYPjUObRY
0ySc5GJEWRDNQ7hYaufHheTSiO0S8jcM7DIBuzlB4AqR9UrOK9M+t7++42p7xysO
8yQPAbjbK1L5j0AFAymIkStr3CCG2zrvpHsLxEiiPsrexsQ51GZcX1eRFV2Uhaf3
s7zI1QQGk9uUmvWw9Ati+9+Iht7GMKPnBytrqa/P3/zpD+hRQ4XnRpo5vrRyaogb
COO+KK7lXghGa2Wf79G6zsy8ZnVvWK4+m+tKsDwzAByMRouj7jvl/Zv7kp5woVUf
2FRpp7RyoVk54PsYSytvaK4QY6G8Ev09EqBCVTM49TSXrJ3YIIDpvcq+IOZ28Wvm
t5oOvW1+UTZ10wWHDC7oxaw/GgLgMtS/TRBYCefmxCQC+jXpsDfFwZNFlPeoFcSB
xGDWZ1m0hcyXQHBI8Z08ZclIjkUPPWpjx0c8/nuJB0XDhDdalsVshsUXHVp7i9RF
hOX8m3dW3NG02kFbL3IZV7xS84QrDiMQynb44cWa1thsA0fjYqlwTFTEnM10kWKf
QR2e65Vl0GycQ50/8iT5eprmeIbdoyb6FfOkgcXTxE0diXHr3or91M4UVYF7EyDz
ROqxwSRl5kndsQ+oDfJd4TUxjy6KOy0LCWRByFgHOoeQkCKSlZQApXvvBnUcvDl7
6rOm7qAJuDOm7BsbyjhSF/niY7MWz50LeF/SvEvs2tj6rjmKmuBW0cUehnYbdV9H
YKq7efojxfVYC0pBoV30GMHpCRRT1Yw0RGLUgPrd3qKqOnPFodf93/kEbO0ywOnE
ZMqQE0Ebgz/yIJT1kizFv19JzwWuPr2XhKG24fHEW/RtmVgeI0ZR5wpAZk35aJf8
BM9sL4P72HWo4VxklrMX5BraTxTTP/rXpEQOURtWOpDj41nOCbPcFS+3/I7F3bBg
KWR96X3/OcleqX7VW+nTfdvs4pn5e2bTs11HYVFfNBjoNkuU7aqUqEn/LuiwJlqk
4GdlQUVJx6D2SHFSzQJmrb2z0oqTWTCfrsVfoorjhsCsvdPjZVgGlNN9l/GXz+19
9mkEFhtE58O2ZLa1lz3mlk9Mfi/TO6O13yZuBeaepGlA64YE7sZsQ7Pjdvc23Qp3
PhVEZPFCtz9jusclV6AGz5k5evoXpxLDzJn3PhocLPkUVtIPxRvwgf6cR5l261WR
Ys68CtHXhzWejbI+mLTjgO7A4xbWVxsLeHPDWZ4w2HKm5gkQ7JQAfckrzN0fiNON
C7maIB+wx/bj5n9YzuTm+RxNAo1S/0M9zNLkTvWoQQy/VgfboaNYRXOJBS9fM6GG
KNd5YZ9zOI632zEslL6QfeMTTB6AzEzZ35E8CJiAmlnXOPsELGOjm1sqVhoHJykx
ecOBWMOrrYUnXw0nEgukJstffl14ZLi8d07AlXFencFIem0fLMp7SQwRpL+LJRXE
qOkDIOSEbYKQwy61oXHF3YZ9NzCdAzwAivP5Q1k7Zxw81HjBa49u+rxxG8FG+Xxo
ZTmR/4h+a7RYuds/9BbXBlNqLih9o/Ftzb4/eoSfj7ZExKixBLEpPFfwu1ca5CkY
wMngQr4K+tTLS8ZjP0mIFEsRfwjne7c4LHSI976Ues7VuU/2Z4K8zHbENnXsrNp0
dZeR/rfIoTfKt1v5TMvqVNabKBK2jB5oytD5fBZ5LriJuz9aqiVbSHJaohpiWi/x
+kPpHo0Wqh7BHWCXjP0nsf1wS/VIQprealAWL8VDsBIdWJRc/KDs8ZJOd6IXU+Ng
CLMqgcxW6uVB5oQNJyOQtJDe3/bcgZapEUjqE/5n22pvTnAfuOmApGvpz2sGQADj
2CYb38AeagPuJ4kNo7+1jLvQ9IJEFPCsWD1XdfbL7FEE6X4jqK+ZjIrSFlpxnSns
F/u0vffAnAISf/6VXkHFiM0M+e+bOE7gxP4GrvDZsLACMQh08CNRTwk3ps91pTuS
WrpeymSoeJXOJz+QaF2Q+7YdH1DA3YzqYwFdu+e2cTA=
`pragma protect end_protected
