// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:02:11 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
L0eru2oDvRhO8uGFeOQl9eVVxXfiaPLAWjX9uxWEQMHry2KvW2OMIcHH1a+2eS7k
gX5spyZ0Zwhe8fTFpyvUbRR4CVsV90iY2ri13wPrV33iqrIlu/UNyGHpClQACmVl
/YawM10BNpDWynyaZA9GwjIFuj1ti1dRdqMIIgqcM70=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9840)
EQPRC7h3Q7ARBXKvx1zgK12xG80A6sizYpMabgwvuo0MvYB57DT7Bk5huoQ+2vIQ
ZE9YTSYZTkKRKyR+NN8WlWm5xk3aZW3xBJljW1ucv+h4vaHD3t+1QC1t1OxpxzZX
0BaTb+vrRDGhg/nIpm3ePdEnAVO5tBuB/UbNeIQ+UcmcGHWkxIHY4tRlZ9qcJc3Q
0qXdBytVxPYKH+Zkde8KLSqfid2qTDgcQo1et+XQKx8PUx0Fdyd31yKtdLZNeqxx
S8vdQjUvNzCeMqb1XDX7/pdF4kEra+QQlfuZfCeIBSx2mvkP8gqpq/+LPh/ywSWy
jZj74d68ItNYxblchgaFjTFEdZeLEn4CWgEOH3qqKy20ZoGZr8nXL5Rug2HtSnue
NmI92S5+X5cNZfgCATlbos4bS21GEmXUh0mQodxo0qF0hNV9ay6b3UTJL5fhEKZD
uZPcILxyyHp3g3GfdC5FWCZgvoIi452045u21v6lUjBSYjZ0J1fogM38qKZzGygk
SqejenEls67VeCcdUIOobKIHSas9Pmz3pWwV8oqp9XhHFnLhUrGL3eR/i5DCZ/M0
7bykejOjIzrcD5CERBSp28Ak330Gu6F9311loc1kQqu3pEcr4O9yb+pwsiRFsMOX
TIUYB30aGe6MnkTYMBooIAQxy8q1QC2PALc1/C6YLS8pe/W0y1P2dxny8nM3frRX
knr6Oe6YITpo9oTqPBKSnC4bu4/aEcdu4lgfZgj8Ev2+0Q7ZnZrvdYgrM1G4fpsF
YBcfKPEAFEdneGFuYlTioS25Z/Ba68ovff3GZZ+/j1KxRup3iuKojAIcllg0GAlY
pqJ6BgH/NKEYVoZ3H5y2ecxLT4nehcpOFB+oGiNYZk2bYsKyJtqBjWlootnQXpYX
ljr8oDusQMNvE5jt3+QLHPB9b1PAc5O8domvkpdudu4vcq3S5b6o4mlQMYrnjPF8
qzucaMJCuHXNzHWs3prV5uxW4cbikfT2rneU/A6Pco6iI0yOPePb6QvcvaigyGNI
ANZUBRo0ciUm8dXsQaFmrKaUqWxkRw4eUgaL2TExaQRtNTnxHK17UX+Ir73IGMrF
NmZfe4KrJDXDWU5la0v4y0ClsMvgTSC3eGGbeGnoQ4ilXWzuTO3bhoi99Js/QKsp
rtswfr2WvU33h4+PZDPh8pqDYByYqX95WKxVWRg7mu7t7RJYCUU8/K82Pmcv9xSM
joRaa3kQ7P7vhugzSXWN7nWGFCLMqgQFNDgf+qZ9aOXlsm78FQ2z0yZNvlwb/LYG
MzhmjchfSUw/5g9AU5GEN1d88jnLlTJYJYHG+1YM5lZWz1I/W24h38DpJmhW1HHg
sruNeS06O9n27qdKCIZ7xOFCcqACdLvDjAnuBiTocI2VLOFU8oR/44tfeBF4Yqgl
YW405r3vC9nqPnD1lOhWe1fOfcakiBfXPRUHRn0mt0u2XI7KDRB99NMCv/UCdrKk
/qYY77zh4ExoxNa2PXHSh7KIfDmivsydafhKqHzox0PiU5a7EsJNz+sZGjiVrzDl
+4hvKtfXqSQb8s8l+JArl6ftCZbgXZEIu8EwET+C8QlUB7sVBOO8GOqPB47wl7Yc
lzS1MKNCxpTfsEQ6q27chYYLl1ZDlY2OqtHdGsmwlN4Mwd2/BjQG35SrRuAIqR4u
UWCdEPeyEOVps3hEV+OuguFnQGg0GFjTvWSjD7EerHrEltjFjkOykyWwYsUfBGtK
tdYao/62saT4CJFoA5i4R2ZJdsDPl7imIWEeZVSBMZ3f7d51CksUnxQEGQ/Dxjmh
7gNQti0VtF2J5WzVf2FFCfmh1U+dRpcJWIEDPbYFDy5+KJpAoKTDvmxjKTEb489d
w4wPQ7ke57MlkSEzAEGZehfOVhQH0hV0FPfyKD05LNbz6woaVFGs48W9HZu46RY/
dJM89MDSrRgJzqLL3wQTsZKMWdCOB7LdIB7So/w2GipBZzk9yvDstbPbcvqw6R4r
H3P6cVVRpYn+1VBuAml4PxFscG5K8d31HGPsKhMxX1ArI6sccjMXbvpsEMdQivwK
FUhvaw7xRToXa5DZUSQbQhkOOLMXkLLOKRGrMl9HuhiWtN2RSLi5rYKQbvOELOe9
APUxMU6aUeyKAh3qSSp9IXLo/ziCSQX07SIflery029fA6ONXHlDM0VmTFXNp2J7
sEc8cqRCxCkoPYSg+X6So/s/DKKHIq4oiNB+4U/rdL49fRsrmT3AMeINHZv9ph+c
CWpS/YbqnJEPuK4FR9DSCrGIL9GqOsDBhMHGIPzRD6v7nAsflNLamKdUDRZ5wLCT
MC8c7J4Etkvlc1xUACLzWkMomBmOG/xk5Bjf9dlQlizxH89rOi7Frqp8sGmuU92B
GV4IhZR8yFMIgAhP4MVPMQoc+F0e6HDmlrjtObdveeAqRKVtZdf1gupzaDbwUbor
1n0p7POD1wa4Em7FWaMSpay+gt27H1xp/sRZMxmQlO0Lxd2ipUOIdxQa68XW8qoR
RxXYOhbh0ZudkK3pVRDeQ8/1mmO4x3jTFYc89wVYxVuHmp5I4jhWai+vnC74bgsj
HxORHD+7U47wxhtNQUoIA+8+Zhi8FIMuSF6rx31vgPdXBPC1BsQDRMrIX7CxSjLb
LRak4CLjLpYn+4zp6S92Yp038izmmaCRaGB384x/JdP2YmpWBKBSGg2fZxQLsBsW
KmRMQ/37Ogmxt55GDN3irG3NZqHn5FBH+lrCIXLSUWUsRKtb1YZFSYPsW+OV0Geo
xIBhBto/6cYTn/nvCnIvOlveKh+PWk3eWZFAMf8iLy9ak0Y5pFbcaICx0yM+3BNB
WNAbFg03npPwc59v6bX9Mct2pmSXOsUICHVm3evoZ6LPlHRNWLCAPNGwXfL6oG3b
MOP3FPkwbH0ReXcgnkdxd7RUC65VJNokeMzpsjtm5iCZougri0wExYx+wROJ8DGG
P/Tyhy4UlBOQwy0TUfgXgk3fhxdjEKmmciR7sAwL0+/v5xG9MAIrh7eOzp0P5uJR
Gm6A58TPPAqUqw3HttMo3N8uMUpZHHTaLyz0hMiys2+rEPeZXETLnimSJTwdMzwg
LhKbWoqLv72zoBuKOBS2Z0rHyPscKteuekGT7F5koAAmxM/kwgBVn5jlEZkbYXbO
DaRL4izxbNkmwpha2IlFWMEROIBdYHZzWjoMn0IsjZlW5aHneCwXnoqKK9lhDbKI
zK9X31Gs6yCzylBaPLc/QmRfFs1Um3o+lXNug6bjSiWa+2u6SYP73f/HwK8kuD31
CbXZjilbIArnjR4VU2GpJvIo72kijJKtn7NhefuGQF8zdf65yepnJ9AurB6p6IHD
Hwhtuic0lRa8LQt84nBjrEaDvk4Qj/QoOoAbdmzsuldn+A7sv4dVFevMOyur3OeA
2POx0ABKWS5mzGiWdw20B8+3XRPcEAvvO7usm19Gpw9U3HiPYWSKC2doMqp2bDI2
elApr9wVbLcY389UXsroxbWZ2UbutkoDhkzE2C1LNq0/Yh/yjpm+2M9/WGMr20X4
KLiumLlshb2aNVAa5A5UtzUHYTYonvEJZX56ebwHshx0bDcsRCQu7l4GIbhYPwfQ
M0TF9GH28T8ELeFJR6xL1zQK0mYRxvF/lDuhaA7C/eB7rNfs+uQKo5l2u2lJZc3U
ymctnXNq+pjvRfQuP0Hz2g7ZXEbGZTQTHQriTX384iBvEgjgw6wDFM5zDW8j/yaN
LiEj2H73zW0PWpa9cqL7sZajsFhAbJF04yj2Bl8xYLdMHpxOD7B323rWgtAQQCeE
oBgURDt+wFu2jdEHlDRe2yz+LI/LDETdbCkkSMjEM1ExcMHr27h9SbpEoPrT/2R6
Z0SnX4JSx2ajqbpdeDytHE6T60wy42WWQvwPPJH7GUQpRx2DSkTNSxBDetQBSqKR
TRvRG1AJ3xpTTp5oWufcHprForWo8U+s9hblCoB3HOBB7tmYVbCbCvM285JTUdAY
WjNtzDp1r7yFrp0O8qA/yIYVVi1cEvkicD0lO+bzsoiTZVC+Zvf9KXiwT9UPu6Wj
eD0FShfdPKnwj4ysj3x124A7nDFKTc9pycIJRQPJf96GTY+YOjXLRRnxpgvOaMRz
pWB9/VWK2bN1RPFp32E2EIeeDZkRmAKNVohelUpdqmbGtXgP2ve9rMViTq0AVSKM
jTzvoI2OhM80AngMl5nZyi67k0NfK0l7k5GKr9VdewlUkBV3cWsf6Al0+kwETvKH
5sI7cIDZWVaDUOEuRQa8sDOYkIn+2sYop5vBbRopPwrLZ59bI6tyqB6vmG4BnsDC
xD5i7JsON2vP7yMTCBgRHi7GCm9g8JM7dOmmIYPJD53UTF6YauwSygja0Cn2v6OR
Gku5LHPTHAsKUFpU2JAY6lCD7lNHp4MpPLe/S6rPhfP2yMjaeCN4A3vfcMGRPU91
yU7MtTgflOmRcbnn4XbDgK6mk7dspkY0e7jX3gxb1n/whkepLc3jObkW7lCkDsOQ
i/hgh3CaLQuNOF9CUD+v75Pkp0gR6XSKrkp/edFgWcMWXat2qYrDhE/zQukKiMWA
japFIb62gKuWbBIobuu/jxDTeusQ8DUHPFBwcnvILWP8gCvzesri5+kC3SPYyNZq
zuIin7r4LyBqujXkHrspfvLEjQuvlSsxd4i1e3I3PNqDSYmC0RAXHhlaYsQ5VZrV
91xmqeQZskfPJFYowXIUeLwd/Kat/8Y1W09GjvlyzwvYtwPGLXPsNKyszVkFYS+l
Rsp4UuL6ECCraRvchJxQyUg+Ph2NOolHXi9t0ITXqK211kGbGCk2KNxqTj5Q4IYe
NOGDydbNxLduIXjKF+tjq3N4WGcipTTj/yh//qpmWrrCKG14ogOE/2TDBbmOuv8b
dLLJ5h8P5+dSDijkLsX8yxve1pd6Jr8aV76A2bmmVgi1iPRRu37ohMzBIh/nYEwx
GRISWyw7bmYnsu1GNm2ZcwsNs2WThEbbD7AnYGApWR0WkBY0HJw9W6+G65GjboVK
R1h5fMcqxVMuhdGDTLQPl5fPTdNWCmKoY7kECTCMVirVD9sDNlNxL0q+wwjz739L
V2Leob1R6tT7RYFBIA2a/xx3efJb79BHEVcwxnJazxIg1YLAWh09y0devEL5duFa
5p5ni60e5ncMp+VXGGcPEyIX82E3eGj83lu04W8i4Xd4QfVUKMaYcbS68JssZB6j
rwsACyK/jhj+bmhCj7ZYhnEYuZczy6zAdnYURNR3TY2a5++f0aUkVc7Urg4xD7jA
aySMZh9AOybERb+x8EVb0lvpEyxsJhafZtXDjZ+odNkxDpbqU0Fa/ZChAJs/LuUQ
MSm9nU5iBdFjufxrUuQwewnGNq6b/iWQ7liBjJILSnqpk76kFJCTavQzpnGX3biw
lMHClpS6UW3zKyX+l6BukfKHHO5BSOaPMk5SyXnIAp+VVvfMVBgCnW/BzYpRhjZ1
7xLyeOkH7yr39B9IiBr93Fo5xaYHGkXjt8L3/yyCCHkVQnvgcZOkbuyp3DJ0gDM2
+DeBt5+faEuTQsXut/6gQzHMoZ8IhOLG2B0Zhpz89C8wXDVT2sKF4PrwhEipC80i
eO7EiByQ3evHJaGcAXGG6gc0gWP7yeXkrC7USHcyTe1/gRYi4CkUSgoRpex/EIkd
em1J6JuSTnTJWKYid8cWEFttRLWI/JUYWiWfCVDZFw8vBecc+d0xnTJf/T9yigwT
lEAAKV6EMP1FR1QRiW7J3LhAinbMtuKz1xV54Qn4vl86f3H87YfVVTdspbMMmOTx
YZ8ZZPHbC2ancPBDmtIvPPb0n1jYbIUin3fPqIXhX5GB6pOTpWu772ASwS8xfP9j
An8sxfHHNRAkavteFzFIxOALf8HyhLL9OqaGs3tuwN57eDHC+DbhTAbSIcPupnmo
7/w2EkVXsVfQQJd1PsFLXK/45kJ/wFgqZIZckYMaIGJ+P9hjtrZ+0KrjamOd9kfp
pMBSOpFt4Y9Y1qG7wH3wkSFtO8GA+0InC/E0TezOCTBXsfjAu9qEo2zhxdml7qO9
8wZPnl5tHo3Pl12+QiGVEG72Vh72W/P9Rki1FAzkM5/WX2RE4OcbMYd5Og0hEDqK
G0sZbQvl+qpbxNkuiRIHhZhQknMCXt5W9+lWOPuT7HOmYtM/6krWDv+tG/YVpYjZ
8CtV9Us8Q3iSGr7/svylJ+2u745R9clWUTIYwAVVy9XGQKdsGFdb4zvugqxar3qY
wCTV8oqV0QV9jHrQCo2oAYFc/vT4nRUrhO0LqoM3C43t7pL8VmRqQw4UZnsOx+Rf
eKU2CuCjFX4dxLnqAFyquDhcMIjWcXjWS9wj5IlzVV7dziy1Fp+l/s/XAnJnnkoQ
oYR3Uvn/62a5d9dHMd+iAnjSOJM2Sx5/EkFSrris81Hg3Uj1X4f0wg+BAeYIpeOz
78+qT987eqMUB+0mXIJlWYE7Hp3xAEEGHuLN+HK19WlmSp3kLlOt5wh4lPCq2lzr
875MkSPVVP9nX++JHIkLo3ANeGsuEwciauiIA4W36EZYJMY4pRIF+OZ5QdUEtTPK
wtXHv6OQ/8+AF7k1YqQt2s/fzyE0a3mh3cbDPJEBCnq0N4PJoooZgkUZykcb3rMV
INM1TGjXE3WKF/do4E206OQ3c/k821OfbRwbzfngE789DGKqJVxENCV4D8/ftvha
f+JdTKufSDmrdk1AYVqIiZxSbMCXUP6V+47lR5sZyRDiGONTnFNw1SV4gxiB6tvh
0G2xGhb9sPsOd7kZFcLsWo6iBEU3LhKGM85b90KS5xxUHvI0rUtcivTjj0JqQr6k
YZZ/Si+09ZDIqgFZvURaM6AWyhS3iA9RmvV3cDJjpbLPy5nOSFmEOuQUwGzU9+yj
8UitLhLe7uq3oESLTvCYJ/Mf3NEJiTt3iJmITh/fYKLn/t4wqIqWGKtAEl2VNRVu
ohHO97CO/P0dBBpxw8Rha36a6pjbTE3APGaVWbjxWl2dVJ1Ss54oHMGZVv9QC3lf
HtA+HzEtEm1RnyJmf5oIPMHfx0YGp+WYOdB3kIMTZuAjEy0DB9u5hhbLSm2oPWvV
54yGDM61WCsCU/3ZsUVeet2IQAOnV9sgsb4PLLSux8Y7PeudElrdekWNdyVwKQEn
ZzZMVG52+TXUaIVCRKRlFhjRFmTwz9b88O7/fn0WROXZRsXvvOMG51aqWOFQTdvf
KyuXHM4B/eYfPTQurNrOmrRra2q0iCff/re8SHcy8Y19Trv8JdMOYu6t6rnSEwWh
IuHz2RxXLs6SzOiLmYdI8qVDD/OcQyHGpzdh+fh+Lyvx+1cNXpcn6xax+EJQb+Hu
JJEUME3l1stcjrufAbiD0/wO59srfxQixxHYeZK3DKXaOuBYLzJOORNWTUVNtr6H
fnfr0wo7tZ/aKJiOXbWExMtQu4YHfeRg643CwoCLvO3KmMGJij5M+rTmMlArLhVs
gXVTWbHdJt6I3VK7uHEXaJicaZCwm/pmSGBMh3JVFEkT9s5Md+eZgR+w3ZPbNGuC
9x89x7yLqdB4zinrAy+qAYkfeDl/xVT1p8zc8p9Um/fg8ujiinYspsk8KQRw3Anf
9dif0DKDjNCpfvPq1XS/DK9Crjw37qve62FnCHetYA+on3+JcXWWMWlDuZvfNI66
9aZcs/4upVIfuW2GwZpLgIroq+5sdNOLXlUGOn02e+6t5L4+q/oL0D4PKAwuBUts
NpWs+19wayntztBwYlS9724qYqMtjnLuu498LASrlqtajjm5PncdO660sL4og7y/
+qVa1U6Eh3Tb6l7cNVejvipgB8pXscvKcjH7RW5Mv4pQHEORk9BYr0T/1aViciEY
k3dzL3qpu/w6E8VCwToQcNhHY5AfgadvbCJMWWXyDluxtAhz3bTpZGaFU9RKRZDy
YzqAu8TFcML3SbEaQcTW/ggUzwgEhERsbnBgWT/OKxUA9P8tmM5+IhxzYGma5S90
Ml9qEOZcmu5G9IpjZAEU8OtmYIVqhDFpmmRYJltHEkyZ1PDdm03NsUWDmiEjwi6W
jolqUdV1qLAwiCNywHn7HAiYcDVZ+GTCB6F7S4BKhtUKT/88EAn6QRpmdQ7vnnPD
EgEfGpIl9my6YCBNaka2pbAiEGXCXJaS0+XMa5/9aoUhSZw9vn/4HkVuVGIABYlZ
ZEaY6GkYOpNGbg47GciQP3qR3bxBkNAOvfMRTtSyXD7pIJJHUVdrtB08rK6iHVhq
ezrzUWmj8conusQAkTR734/RVZWJh6Zd26WP9Vj1BqGVTossjhXoJ8oVVrQF5rC3
yCBZYJNxUe/cR9aX6ElJiqVfJ70Dw/KUV0S97dO5k3vWbw+vcD+H3A/QMplpI9yO
fwajJnTKuz8FsSCdDGxVHJ4i5PqQxpvyGJEt2j/+0Hbt2VL7tRPg+9Z9fV6k1f1r
WWxmQVW61KUG6zoJPwtD6JNsW0Atvi9UXMLIETC2XGC2Y67DNqhw2qBdFAik69hV
es9VyGULcJQUiFge7JJN3SQNe0Mu+BXHDpaWyp1QyEXwGeXFLz2J2/Zm6hdyscWS
qqakuPPI0lSRjDVyzIS2Tcl6ZSPnD69fGKM++lbLSnWQGQDns7PvDv8My90kIkHu
r2lQ6QXlm/iZ4ocINCwOoO6e6bLK61zIb7CbWEMdbJQc1vFl2d2zy0Kpcsiy49bO
RSFGna6u7r/P1guOrqxlWq6AIB+B0cQECf4Z/d6PnSlAFuQ3MsF/xgaWeOAQzgdM
yV6uAblJ2CjR1qGHyaRRMmyZQF2x6dXwlTP4ILZLZOzAHlwa2elLaDRni6Z+KLbC
VB7WBgIkyL7PxjIapMizF9HSFve6JUP7sc3DQH4LB4MUM6u5gzmQh+OnuMC8t/O+
+MKO36AHbGCeRkwz1GU+ybXEbJ8c09uADhzLajwptxEzae2cf0PpC7AT+yfva4uw
0NhPUKPojx9WF/ZgPq2bGQkMWwrUFb0s7z8SqiqwtSsPKYUU3fAD5Cc4onhwpwRu
llSd1PDUZt0NZekIY1IFL34pSK756SCY0QlCCGq8hAbKBknLMBaJk5L583x9R8gN
PEJ+3qvFnHkyQXuT0ghFOogJKEgiWS+OlD3YHEbZgUmypDpNjo7jIrAUr9rjdgP9
IQmtJHlv0BW58z6lnA4gePcawOvDYlz69APMPuVC5q+553QI/JcSqSCSKU9PSQAS
3WdMI0jOWFPxGQiOgOT+eY2879skK8YiD/Ej+y/WppNbnMEn4RlD4mG+1wtf3HTQ
yqlg1wj1+mJ9hhhfoojthe6crBMqADCefSe66TKqqinWlX6kzoXRTWrdhBL9YwEn
dkjzV8BRv2+AY5bs1R6cDsuI3RWwEfPCeb+xhgijBGpVodKxGD++MTypOMkz3juo
9XIc5517hQXWY2suHCiy2fDpqnkeHkSbLvVkKxOfJGSCgPd/1VEZ6ivFR8xcF0Ku
x5TGk6tQPr5AzBD4KwYi81sfpJNoQG1daQcXtjg8qyjgbXJ0xDld9m2vLnNbCK8E
InD2y3/Qk54Hdx81wl+ftOkVh11F9hdx78MsCX0f8/nd3odteajNesZIIwvn6JLi
CWhBQcsZ4jUPdt24horGQOvtkLcOoQKZ/cm5pbpYzyOQ5EuBJ/bOa7sBdOzqiUn4
RCfSSGgacHAsq+ROePM8UZwEIH9iLHmTfVoDmPpaskETs9cWTIrU4cFS9BZoTPjm
j8FxQMe+lL75N/nHISxZJjsqaByrLnEteyl5mGnH3KGSmWXhgfAFZ05++7jXZcN9
IdYaRfX5zYN0OfQY7Za8lElRC8kFS9Hq60x4bkjXJ6IQe0Nky8qrdWtgGNQV8Lhz
MxiZjdsF3x+bIgJW8tDfUE9XObapHRWUDrUf25ifU0JYo3toLM4dEArHQSeHCzro
AClVAzNcUbHM1RymI3BGaOVkCk0XWvdROTXy+yQ47Cj2BBTSMKN2pESylm9WZ/O1
L//3n2h6XL4mSDOty3oUZUQicSEdkcfhEdvC0hLO1HG4lIgydQPX4JJwyoRDXtwC
WMtWJpVTQuVPD3sQ1XMYLPB53G/BAdzR3V68fu+3ycjcD0MFonYjK5lRcptWqnKo
AZVWvNDxzy2qhD21p0MIpmJtISQj01msSfYvw1CfcvKXEmr/vUrm0uz6daYi/fFl
9eDx3WZyaAnuTbHjoK2n+SQA/7jZ7r65dK/mvZyPloCVms6zemhAEDKg9DkUJmad
vE/sTkMU6JOLHPILL2MpuhdM0jbq47VlyK6fummN/gEWwrfggWHKVcVCRSbAuoYj
Pu4esoT/ZyvDgWYCq9r2bV/ipasZToYQItdEsUqo5bB+11i2h/DGzgKthtlga3Y2
8S3VB8f5N/LhmB7fwt9r3w4ZlzgtB9sCJA6AyMSXy/e4Ki5PHERJQvy9Ygnu6Uo3
h9qRnVswck9KpG/+BqaC54dAGsotrSBoECbRF/wNmR519aaIqjPR+r7/K3Q2G4t4
ueAhWuqZvxe83BFZ5O4GWPLnQHLs9q5BNWpPrvUxtZ4x3dE9lu/7Oe32PL8QrVij
rpk++vhLY3jKDIH4XZeyau+nJtZfbzJUGXZp5v3g1WHSc3Ezq4xE0vEJUasx1T/e
hYKOD6Bl/An/hR1sWrx2dWtn1TwNaoCVT29Jj4uV7Zs38Cy89Szdrq9d/HLoiE/r
crWrkntVkdnyb8HMUsZfDgjNJ17yujJzuKFGWd+Pt3/vTPYpd0n3wDPfrMVgGjB9
bBQarc1CnOE26ilyiCjmdj/LSO1EWcEkRktUR7pcB/uxBE1O9ETmcr52MOxo8E11
Ixa/WbiWSQfJeMiTK15Gp1ucRLG1LbdJepw7E9bgwnCdfFk+L6lEO1FvRHwjORGJ
Euod/fbJWnVtsXaHP/OBQi8yo+niC0Anm+kbSkVLuuHm44bf/GTt+w3mB37OWftx
SgRiPaLMH1USpy6g3i5eLxvhOCmurV3oR44julFNNScuOImFlthtVVpPA8NG69jE
aTIgNMa1dXQ20RrGs+hcFqVcBikd117aSglGRDpUHy8qREMlWVJPCdopqDq/4kLo
S/MPdYB1PrykftVDcFItImuU58YbkTP/Y7qa5CI4uFrc68AAHXoSsv8O8WescQ67
XoMhvPF3jw2N3py9Y3ZfrAVonfHjOYLldFuGAEerT+UUXsl+lN69BOeA5X81SK8g
ERMtePPXbMSrylqzsxAdRoo8f9WRwgFA2QIYmK793e0B42JsElr4KsmjPstNfVZJ
5mYpX98Q35khtiOv/hZyRvGExhFTWY+ju9Svus9FLrkk2RaFAh/pMTF4axO39Jb9
M/mvync9hS8XmZTIh2lXJ/btRViHg+aU8MbGVFKhM2dUzdm/qPG/4siPxJMOcjBw
Kw1s6OyE86YkSn3n8j6YBa0AnT0qB8mCBGULoL0djPmMp4z2vUuVvfmQCoJRJeJf
fyPEIW5iBzKZ6GWt/YHUOJyh+vLYE9OZBNhkgKKzNH4HG4tWdPs2U+CQ9jF9mnEl
/12yFK3lbX9QtxE55H+YrLumaa/sw88OVD/97enY4jb9TPBoeKu2Yp3Vu+Gtga3z
e99iwsLClUwdMfBQl9wIuLFYDP1Ohqtzu/3rTy7wv5z5uyogTS5AVu/7S1yGn5wH
YQAAFLCkqcuKY+rZjehbovU1Kokgqf6R9sx6r9az+2gQXqPXAMg0nUqsBrjjKkgC
WFrRGeE943dTDhy7fFxU0cHMO7SP2YZ6tyKUX3W1t+mQEUoFQXMn4C2cm2zrhKb/
LpFRCN7yGwp/PxJ1r5K0Z9wtmzoz7efjN44OV3Xuy3nPfU6Z+QXX6tzfFhL3pkfu
iX04H22hEGN9XPtiFo/qJ5ZUbKUGzqaFSI8e8n9zc52EuRGjH1g24+k3SNjWWFg0
Fybm4ANmkZkkL9HyvrBU/LvnDhGyFBeMSULRmMbHzka9xWrR+bHijlDgECw8GFbJ
ZnUF44HL9B8Wg4gLkpLX3dsT3iyuSd3c9XCEHzuDduDEvYtrYbgFolMZoG2tV0C0
DshGqZis9Q9WmceHg6L1EldmzSB1yLnN37TIfRCDgyd6Vgaag4qN4d+CUPVVgm9X
JTFdClqoTSHe9Aa66Rhop02S/R3OEGWhEdInhXWqpCFQh/+NcYKSNDzgxHhT6zHj
QytHboH2CDR7sTLpEasZA7S71V2yR+nJg2sBqrtUJVDXG9kEgZzTL63ynVG2DHo1
B9W/XZZYNtgx8ngBArAvt/+KcDO9RyWvg+hzDXE+Prni/lB8xpSQad8rhrGd8uLz
6EAH4YoI0j/BGyYgtEBkiVd/c0Yhmyyi0rBYOsqxvo1td27EQBt/iQG3BJmyOu4c
fjSXYwpVnRUCo80y6aGZaCN2sk25/3D9aaM0wztb0HC4sP5v+0xLO+23MIzZQwX3
N0GehN5l9VxmdLGrC6KBMO61rsdtwigZuoFRPYgf5dPd8vbi5HXKIbbOiqmVBAB+
hK9tP4EzfewGW+MmcFwaBNLRBNGwobM1DNy8rvu4bJDNQcKX57xP1gXrHEA9RQDK
wJzTQBgusRM5+B/Dz9ysg4zHmEj6Uf3hPXu3dLRxKsMEEl3meMCbIo8++JJ22jtd
gDRSz025MZKXSX1BICfbt2DdWCeVnuhGLXGjJXuDuBzwccDMq4MMeW4EP33QQCq4
j+dEShk7Owd+aGP81+NT1c6FoodBjReC4ecmjADC9B1aRNyGskg7TVvrOgJZO4fh
p+I560jkohIMfGwouga7f2i4PUjoUi+Moypcs5UqLBRR3E/DoBHxrYxZdY/juoDb
dbzG+bG4mzacpe90KTkiv7mqpwCLwpoCXi0uO5gXtaGf86FiZhoFS/7lYXEGhdwq
6Wnt/HR7Qn8KutDbupjFaSY+D+cgsmE4lEyHW4GrQg6EDUCmaCxsWkvZl1Y617NR
niFWvKdLcT+Phh9JquOKBQ0qS3HecGhQkIyS/EOPnVBBhTeF9pyOSGUtZ+/5O7N3
3zgJqE20qV3IUNl65hbBtMt8x1jAFdxGwuYU/9uNPiApzjtFkXX1NKojGynEPysY
t4NiS1ssJqmkdTkeoggyA5WMFQa9sDLGYYMkXjK+KKJIp2YadXkh/V7iW75Fn1dS
t41vVRdMvi0Z/XhTg2/kjDqzC2YO29VCzZ9mbwNK00WhIcJiN/Lr0UYQgEvUpgE6
`pragma protect end_protected
