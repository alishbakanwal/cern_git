// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:05:29 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Ynpcjk0wFqi/YEDuoX+uzLNE1JHdmxoWAJxjkkwanodUj1VctaTOzkbGaBAT89K0
ortGUKoMPzkOn1UQhzMcdMmsLy/5bdFwy1Fumb0uWN1wLUSBmxO9TBmrQYvBayW3
k81zYK4U6BdxAU7vCWIHe1xsk7MGHNd7QdXFxChpR90=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6352)
89l33k5JhqydpGIKTLhbtxfRxkK9kvnyMjJg56C4m7AiwsPb7WKRsrXjTDwWri95
N3jmyWKIEKezhS0fbjxQHD00NVNSmYKKmlHwAMH5H+4oyxYqvnd+EbXJrYV6SOpK
1VuiMpBIFpKymvCMakMVeqkX4LasnFAMx1fYsZ63EyNNbOV/KOLZmqTU/pypYqKB
3G4i5Up4PfgHeIslNa2MmkcxrOaH9SVGc5TbFmNWAfBtGROs8fgneiyAhmEH0zdS
xv3KQPy3NfcrNzHXJTGeNjW/mMppwPktXPD6+BnJ+9pW/fw+++5sKFiGxZMhubqX
GoTnBJHw6iVNowz4DAdZI/6QfCY35ACdh4iJ1G7NkmIYi8BytYNFr51jTJ1oLZwz
66mB8RIXR3/5NQYWmN7YDkT7VhrgiqZTZI30/qBSNAcfHAMWfAia6aW65nZEf2l4
DvAZB4sPpMtWwoL7fyZAVX9dmHTCF+uDxd9zKyhUlnijKE78V1VJWLAH6imwRRpf
WfVXqb7WxybN7sLlSoibsmo1g3N9BEyYgITZ+hpuISExyPBeob2ROivbJqdTOeKj
53a1D5/AYU1dKeQquEVVGMJ0VS73eMQYYpHdeli0OXdl3VZBgWxmrYeZr3JzvNSO
sHzXfCrEidXGOuqdtg/0+0u+7PwCT0xbuxE4sTk30zwkIzwoR2cGyCvAuvADvjM3
4LhhrsiZsdnCKcXFTSRZT2X8tZd+KjFF8iTr6+H83cGK6h2m6HIXRjx/lmDtc7AM
BAy4Gf3JHnUJHZw3BOrClbGi3tXBsrw3UlArWd8WtO90haeO45oQBBhul7ECldxs
1gTo70GR7BaIEmZnLjGefQEpEHjiS34FDEmEKap2BbUJhfurktiiIKuj+WK9MFHh
1Bg5JDZUjBKdneXEDv2dYPKTQ7hJUJgLLVA1JS1gxpmYzapEe4mLgVYatjQQ0+oj
GBzEmAjb/hjfuuyZD50AgqNZu7Z48oNQNa2IA/m2uppSBmGICPc3aRpRDcKeugKF
mLqyC4tfCKdRhaurBDMmrUKzhHiwd6JhB4juU1QQ6fi5wskeoSBU4JNSYcWOn8ug
/0Mibg3V8z+ykWrZxoP9cUZn0OEefL+bRD2GHdPr1VTxn6zfTEIpewgBfIOpVRSa
QeHIj/pGNVYcMjpkaThc42TSJDVMB3R5Vlv9oDnqBg50WnO488t96lmgKOUy5ZCJ
RvihpYWjWQi5I9qG3gaiJWqM3DOO5PWCOg7ws8o5Nzu4pHsy0/rfX/85AakD8OQ1
u/isTobklf5Gl326EQ04goGnlZIXVVzLoogs2uzmhqQS5LCuGJgmc0BSzcCMC0tE
EJqFAOFBqpsWthulXkaPWS8MU2MYNPf/+BSYbt0JK2gTTadt7mH9MayknUxG0kgS
RacVZYiCDwXogxvscLaLdP+Ag6QZxvmfj/81xZgDiR186adDKkuVqONkUXiRHeei
sy0CfZKXov4ZDDIfhcpkfSoQFmhVVChbPqvq8s5Ix0igcCS2dPH3E1aZKLGk0u5z
TYO96WSMZeigHo5cRjAUUyo8NIv0Fb2fs2aeIQAqdMtIuhGRnYhfrpXodinFLZlC
RnzjUNvm6wGZ4Prhg5Kq7UNAApMDA5zRvZhsHaMGJ9nDJGoLRqptlB9wcCQGljAV
dUTia0IM7/s2BFz94EvDUIb8YaVqXEp4qfT24GCCSeuSdcqd3y9rjP10QW45X3UG
MMuP0ZsEapLl3gA4zl0KUi5RBgkEgGa/pEjV5RgwQ3JG6p7n5GtGkzN1sXOvUuXA
NVlvG3gA2PfYmjfJlFsZzbYzG8devgK2FA36bD8Znbnv7UfGoAwgdrhFe0595YmG
HxA7/zhzOhu91ru8lV7CVXpudqFGcPQvShONQ6MVVfV2DqnXIoi7BDsdglqf3/SN
Xkub7ZdVdNVZBGOZNC7om7U8tBza7PMUjYL9HHw8WWFlKJrjfngrPv5sVf4/u8Rs
UAxdnf/Aozu4+/+KP3TWybAMXJ8D7wkABEFiibYKUHYibul/Z27DpxRVudEREpKP
ECd8eGyDSdOnOaWHgM93MxD175A1HQ0dTjLarVgnYLH5RSXNj6XUyxjH+FdiS4pf
nQcVToN8hB7ZH7Hrat9a28RalApSAFFE9SBi0Q4kgB4M3Tfgk8xjaiMsCouRaBOi
XyA9Mfz62XmLNBES0aLJE+n0/39Yw2xGTSMYeDO9aNJPRLKONijfntf4w+pNqHqZ
7mFu/fVn5f5PuSAx8g7HP/PVU+/mET1Vu4w5a9dqL9ULIEgyNHlVvTihb9dUmM2o
dBgU9vEa+Zsxk+t1gLxAQmFDVTRBstghTauM5t4i6EqXVFyRS15vidlikF2tKYeE
br7W5A6MuOt1vXNdMlr4ig0ovsOMryRJiYdZINNgyDajkpZzd8Mi+ZWntupovMiS
8WI5Nn56q1X9bxkU1HhG/UjLAo9Dedjtx3Ts4dlpZwaS9OZ2so06IpngyI/+OyE2
nwpR3hlaJK+P/akzVgrFSwpsshAuHtf3UxeBf/RORjkS592upVd1B/AD94/u12c2
6UVRM2Z/YS3OV3f6xg5AvMU7HUyhRtSrJxH+ovxj5hDy2G7wik2YoGjwxGefufaA
S2iEbkT695MakhkV2CbFyVXKY3HZBubVE7/pjfnigUFkFKx7hqg3Xwryp4rwTGq5
EKJ2VCXMTxzubtUl4s6cww9baA+Qc0n6P5Blr3PY6oKuuYx3EHgSttegWSqCj5+3
whM1LfV8z694scZaKTwTNTWN2BLfYFtKR42cLTxo/0hF65+72i9gHmvv9ge25+dL
gVJftvgtO621/fCCOhBLZYE3aPpmcjh5E6XHTydE+hp/bgO3rqY5/DRGVovghcEy
3JBJhYNqO27T+7CDpxFaWhvInfL9GYPDfQLBTw295u9RaYBArFEnfLqVM6jChLLQ
3z8PxIRdWfL5GN4Jr1tvt0uOteq6PxLK35kD9W9046v4f15vVTF6KbGr63efcN4R
26lLiYHIUSkleKXwE1Ysvze140tTapmB4oL9fzDDuQCror61Djd7HOLQd9JI0kUR
aNcNeVRsXC7g+wdCr0f/xkt8hDzEKuNC7J39+9PoaNunB1dfw4VxvSD5NvbTUUUH
3iCCkF512IxsXqD6sWEsGds59FjaHyY/3ZgJwJ4ArIMduk0rUEouLmSS+HXSXrYq
UpyAJwkTUt3uqku/kPTmHChdjqGd7adY3AM+DM1hWjN3Rv8LzPCKsQU4KM3rkUGo
sGUOO3pz6jo0GasjFEmDFqsTBxDQwWmMB0nNXRd5yQxUq0tA788ckBlR6NCblaqo
nRApfJFQV1HUrFvc3kp+RjkzKYdoT4CNT2Co9cpvP9QCx7mWCPZijLsAoRZOSrrt
vo09PWmD8B73b8cUpbTvbXwZs43TU3UPpiZWs/ahNcxa07l/tTpJW5RpGmfCChud
1cQytC2qWltvnSUNMrx/0M5IVBto3A6/VWBQlAqhVZVFG6ci3mV10FhwnGNoxUmE
xhA6QivEm4Zen5vK6/07D6EXCy9x6TG0H3srYG6hz6usZhGvwcD7w6bCODOpudRt
mlvN7pQe4R9F5It80WaFJYaBUoRyaYexe57HF1z3HeTxxUCsPfW7O7xd/cm9drZf
Pcq5WNFon4VfI7B3X6fYZHJTjuOdgOWci0TPIRYiHb+PMOj3NJeMzKcmRAeprEYI
KNupa+EbCS0TKnyt5qn35kOiIMac4uo69vu7acN+zOWX+CVRbtbKv/JlgLU1BXHi
SXNkYqHnH/nhYnYg+M+FoCBjOd9Azw3X2lvbl0ftJ362wucvG1rtwYJc7BPj6ZCs
lerNU3Yw4J4t75En9ZgtqDGwlRFOCcyehLIzdjC2+hRsZZnbu2A0rh8R+eJgSH+M
eTXlgCuavCFJvK7ZNn2+6d6gW9Ac2bjTkbfoCzCa8oQn/SdOU5pSkGlvaaMaswOZ
7Iij9OblZ9nWMU8qbW2DBh/LDQe8xnayJfJmC4rH2POKIMfPkQmpVqjIn1XZWaN9
H/wr1cDsV3zQ3jx3I2gDxRugGf1Z20u/zqWDaD9fvAy78Z9PDiFp39ALescE2Vic
W827E2fEb4rUW8L62iKDdh3/AIb/WNY9/QmVf+hp9rVi9+cAcpXU3KypCXuzGoqU
jHBvEMHaWg3Q5hj5zLRAqFo94xDCWXbV0vigXl8z/LtVJlr+qd1P8PYh7+kBBodN
28dFp5DgbalZ0lBXrR5XsqWCwIYfJ3qZjMFaY16yGiqbaHjZJScMMxxk8hGs+yhY
ZjQLlwI/N7AzbqaXMlUIU4SKFieMjCb43OCddiAQ1Otbj6JbvOAJfnB+L+t+UkHZ
1QFBvW0mJScMvE6IgmxwcySYqK7iJhpckoMdnXoKK4Ci4DRwZMs40vQso3V7OdWj
48DO7ywx0g4og/gnABjidgW/CLH1HUZuNJWD5VUi4AFS5bbZQ5OIMvc4AK9daOOh
WZt3jn2vdka7mWXH8Tsqm68nVaf4PErzrIKKpqupqNB3BCw3I19KcRucnM4hq/0A
FpotgdvneOEgxqa5vdCjUUQ+st2eO2eEmvbtchujJ0iuhONHBSQalN/knjJEM3x+
Us+PIeWyLmc4F0oIMlKJSE+wyHrAh+UtTDDH+78LlMrdB/o4AcE89UEcc2PeKiId
z7bj2qgHT825qRb97yvDHb7Z1N8vvUhAnqeA8so8WpYmf7Dfc2G85WTbBuc1NqUw
5JAI7qqAAgaEhy1LCoAwTm2/duY1QYLaKKLiN8AtfYPF9xufqU4fqygWbRWH7mHH
KW8R4anLKyoq7RY0LhvP6juiFvI6I67RSiYjv6aqJBaHpjsHZB6G1SCFQb+YkjRU
1wdBxY22nMg0D/U175tPViD4TeNe9XduMXZsLz233jsPcloJCpCTHVOmHNwUSRfV
utjtLoX+aA38Pv46rzUwV2HU9m5nZkKv+mztwq9l6IY2jyzNATgYmPrado9ioTyQ
7vRqP3xuss0uEtcA/a9cpp7efLnupt/dkKTg1Anjzs9o5GGOGqCaatQnb4OqoT+s
xPdwJwMaoHAfOrKIftYJRAJJVG6e6mAWnmE1k63+FxQF8CwFajg/v+W6iAq7Urzh
+ZvSFZJWZzkcDZR3V+s3y348mac0twPAuN6KjqdBd/NXPnMs2BjwlnWVZpqhmTUm
Z03b6tw+0C0UHZjorNZFuCh9iq7qL282tm77oGhXZzo8MKRa2x2tJQHEehqvoi70
JSxRPqLcYknwWnvlW9AGZ1v7Cjr3HSDABU3KYgB4WCpygr4Bqs64j9WKpBwTpNpE
iEr6kZGSIKk3cAkfup1StMGFtAz9w3zgXnONlgJNz2FZLuoPdvgShq1tHBtHYSyr
eBSlBrVEi7RFiWii+OHCTTf928XwJvCzpRcfTlzumJgq+K9qgOnCWC5MOcbJAift
s1YukJoJZlvzYU2vY47uNLGO2+Y6l+doALO3CzwsWwpHZWinvt/qpnRBTrupbLpo
UhcZjiq2qNlag04Aqr8sNnBo6t2IAxfeUPK1Pdem7og5jfJXdpGLGTMaT1STv4cG
EJuHrff63vDSUyDyXqLNy5eGXTDMqa08hhNh58XdRYm3an2aGDNrg/n4ivjE2Cr7
saQALI+HQpFJ/VXhDrOa/hbaH7xF8OvEoXoEO7uElBzSFxFPtNASP5vgzpK2uaXn
bBZy2Q+boi5csHm1fXxzF1omYyUWRNAZBFD6W0ALICzfRMnLqwjyyBTxXQfzL2mg
zP3eJoFCZDU7n9yEp7VWgqJ/9uD9SmjYOxIvYCBO5cOvzPU6i61aqQigzFjj0kwJ
3wo65HzQPHucGdMm8KaaJ+xicLHYZotYIASchWXP9PtN9nacN/sF0Vv4aqIokJqu
FfGG5plwq5vd4NsS4sMtTXWj2CKDtDNv9nnQQH5KYgs2e+qHjdeOqUXrvjoE6Z7c
h4XkEz+S6okOSL5b6ZZTHmYsAQGgvtgih3zdWmd+TetTQKk1eexJozLsNGta1znW
8mRzwZUSqZFG0nIZZB9TOl6WnNuY5unKXw3Yq3tQVXdesxhZhu0EEfyIcwUF1BGX
0WEQQ2WP7d+GwqnCkZouTBr9dAfDQkG7boN+QB4m8AM0j2LkDtNJvmRfyMYU/xtN
MtfZYX2jeMjsM4qLt1Kyc8X0dVNbrdwTocyL+k8+E9ICMrn8dZxhXDMc+UsM89zr
tdiX4UbhEDi1sMA2wiGpy4DaSderFMHTJrB1jomfkQ7OgjLFv1PW7hNiAMX3KhXC
t6zskDPo6i6EoP2g9yMRXTl5o+kIwHJ1BBIxPBEDW+YMQEuHsx7D21+IFoB7cQEH
dDLMqFmpj6kw5pfSEmrgLi3xm0pNt4EzW6nOHr7tKXQTAv0ioyUjrPa0332I7JvZ
XY4grmSfuURebhnljl1saQIINfS1hpj4TCeMfWYYvZrBILru1whCIlRsw+ox1t8x
65wYAc1nHiXYwXAGnrHLJfCmDY9umYVWYEKM1Yb9hSiF15Nh0dDXmedN4Tv7FZNd
fj6ZQNIxIYLiz+l9aL5cmWERDoWCDo6tmE3oeDYMuhOjK6Xem8BzJ9lpMhjfC8Am
hYuT0Rh+N0UdgQKqxGFCLofJ4af8tWIHpiCCH+fuUGZHsDByBVZR95BqZPdo9vSr
OmbRIKaOgIR96NWVE/7jwaXZ6kyf2r9vIvy5RZMieTv4gzaLGG/lc9QJK1VkuiBA
/Sq7Q5JZ8EN4+fvqzkh1CmBoHF9HuY7uDRqp0+cMeStP9zZib7IJV+BH63eZXW/y
W2us0m/C7Ixaeblh6RqxrIqxRQaLGcLptPJi4ooct9f5LE4fvaPAABTOKpR3jCYO
Y6+McH9n1rwujdrG2Ir/NgBvAKB3k8VNDtvJB2H7HBnminhMCM8DPgNM3MgzVo46
HNutx/vz8/z4LLwny6ZCfp/6yXvP396/fRdpVichSuSHKLwz/6XS7J/4YjzuW2Lm
FTsvQC5vnVq18BemZ+dLcGStGUT2YDZGwp50XFCLFgfTzMYJYG6BTr8gXSAe8sAY
SQY+hEvItRsx3/Dmnyn2Hv9PFFwADT1FXA/D2gvQ+xRQp5NxTe8WIx2cCCrxtM+D
+++CLP4zlNU7ZQyCbpdS0HWYJEHOwCDPvBRI0ZEw7/kI9XI/QxujCaQEqq/wX7Y3
ZWDsXirSex+3pqefKr04G7wuwAVzu16yJXcUCeYnsuzpRNtQntzzJd5DAJfTO9MQ
bqu4CS3uMBJYVxZ7LMqemOBfF8DA2TxE87rI9PYYjReT7UH6tedSFocZJ8GO7F9W
ZAKK9ZN1oaGnTh+Aj1WI+SiLU2KRuCfDOhstvDnKl3HlOD97jj8iz49z0irsgejv
Ti4MAo7klm5/zGe1uWMoc2HB2QpS2x4fpVqZ8YTomjzooMR8aDAal2N8x9M21n9h
e8L5PRYAXMb8ytEuz4vnox2jdEYZQjgBpmQjJXgXCF0/qmRgIkLpwFtiL0yrQwRk
AxCTgo4dLMUlPaPv3YtRN2GaUlgTy0KAU0HDSYRLSoEgHuzU439wJPF23wU+WX/+
wYT7rm+9W2DmQhY6Serz+FsfsNesbSGVwWYbu+0hlQeZW1x2RLQsDeJtFg5+QLX2
wNXBhJ9PIZwgZbEzIyJz63grH8/XWamoobQNZGOB5RBewAgS7NKOUO5R1T6P31xU
goakslxeQebvZUOipeul8dK4pFe+KeYrdqFIqCnJ4GO797r7Qz42DdoHw2zSbywg
6MujBm4Zv6njdgPmc1P03HTzN3UKd6Zbgw7QUufnst4JCK46OYsdBYcGGKHyl71H
odOJeg8lU7vvXNCcZCfhnFfpqqqnSqGJgXC/dM3m3jIGCDdn3zMscDPLPpnB9O9q
tOmf7OqhlfYtJtvZDhQeSVW4yAmfmcnXsffscW9dxDNzNZFe9MXjNu9oIjWmRAqK
dc5X4WP2RTfH6bvY8s7VeCH5e/MFpJYfpi6lICUuf1Z0RYvCQve2PsfX4OLPaFRE
OkA5zNMtVRlc3umaWEM6WfeJpJ3Ri4ccBfAFgr1UTdB8AvoamJq8fYL8nx1AZj3k
ZiT67hBToOGFH22pt2yXFEV1nYQErB3s6r/4+ndQluc8l7zldcLjIGLQJT23Jlaa
r9cr+Ew5qJ91AkcCCn0hHtEmU7MBCtRlMtdYwYjYUGPG4+hwW3VyxGG/isZc/kT7
gkqW7oyU2BcJMyZCLyX5NPd/20rUGh54/Vm5GxPPrgruqhrkQqMBY0Nim7h/DItI
dWrVY5RDJuZIzbmFW1nF8mAJsA1N12M6/D9vr40sxg4y9BVbWU8g1zYLIEsoYHhL
fBSQJOXtDEh51ZW87Gu82V5TjHBYjxUx49fpRpy++kFTcJJCVNctIYWlKcWoqXmo
ancw3rhob1qxqyy5YmQN8RiT2XCRF3a0/tVg7qSiM90f6zi8PK+/x3Wh9+Do1zuj
LWl5RfJTwKVbv0P8fujsfA==
`pragma protect end_protected
