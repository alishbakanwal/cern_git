// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 13:57:45 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
OfmqRkb71yBjvh5IOgQ3iiJdhTXvJ7r1SCRHvlkBfDFzu7x+Dj5uHxmWQXla9w9H
alxYkmZrfVRUvnMIlGq4Yiynkwh7pfvBcJ6S8gh4zp7HcjFToi0b4H8TCYkwUl+Q
OPVRVsEw4dfKU8zVD+0Wrk4deCYKpcZ20oEJxzmqPVk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 71104)
5zy8YpWtWbMgjlN7+9M7V9sXqC0fygs5XiCRlTP8jwVySDZyr2TnezzxJRsqcRf6
ZpS8pc5EBelmRGolraVh6Ggsa28J9rrZqND6nrp+NY2FVLyWoDvpkov3QN9qa9fi
D6XaQzMIOOHGBxs/zX8yp++UCuLzk2IQsOPfLdDhS3nhxy2wyt4+zUQpQKTadK50
WitMWdBi3wFPkBn2xM+vsSuNiL21YuN+RY93GIshIx6iqt5ST5Lyz/cFupw+BPf8
HQ8zkX1gSCZQmArCa8nbKrtFX+xwSSqQot7yq8BIAxG6k3qk8SDttuHiY1cV/q3A
gPzKNzgsf54ho3iWbNLYExPyppNWADtuAmzed82/nxmipG7r7csoibRNLyEv0iJt
+YJpn1YzyryDRcQs6i41pltyEUPlsv7TZ+PxMQFDC0L8VF8GA0Haxy0FriWsNaKg
1QnvurBt+You/1+qbKM4mQB1K4C/mgXeLNMpXv7J2TgKaWXSMEpkF0Jg/BD1RZyc
CGaBT/Z575GNA+EcOfw8TinxGbSDUNLrbO03GpXnfw5rFEuwwVM6dPD5UyNYhvCZ
UG2IpZS28jSsFcQ8Qq1pcY2HRZ4nbiaV7au9y88/150qetggTRnt0s0Y+eKV+vIP
owOQ1wEYsM+4KHa1pqZQVS8EZNuXvpV+HwhlSc4sBri+2tnhygIVS9oFTJ8SiTVL
OdXdGPfMsHaVepBGZ/gtLAMmhFXm3W1vtqmdgwJM7lXxoEanZZaUV6rgznW5u0vK
ZfktaZe2D0XcpVUR2kRUB+mtp/7/pNn6Tfbt5aJFid0Ijrn+TblnCqG7rsjozCJE
MyNRYBhTT5lsYD2X4cwjfDl+9a3+EdfeLgJ3no9UUxDWUfFNf4Aruo4opWg+LU/q
x02aPi7jubHraAodvVRpxMqIwzeSgSjAFoc2yL9GVU866WsYAd3mTH2mYQDEYTP1
mARylVwRr6l1O6j+8+ozBjOKuJ2YSMiF8Yp2GZ0t6rK6u+WZkBD/YIqNtgnk9H8k
2nSt9YxftrcVoPRv3UNsK38+YSjKhftOJLAP0sT31rDE6J1t6iBZFbveDwEjhQiZ
RQbyIChEg0/0eq13dkEos3ajFeuvE/ExRVtYKi2tvXcpnV6cSQO3HZo1W1SJkb6t
J6AMMpp+l0lrvu3H/oYaRuyIymyi+28igo/kWq4NLITte+vAEWcgi7EynS3dwHoG
RCGASu7EwLa2tCgIezzJZFzXbi+ASQlY/+h1dOEUjTG3JcEs824WhJx5IfKv/qo6
w/pDlGBCwC1AqleKVcC5P6L5WpiAoTz8mQxFReiyfY9+409oKSxupQD8QQ8ttZta
8xpKdmtiL7Dyczhk76LwO0eJGzbv62OUNPGUhUWQP65IlwxCrWDUQdz4yaAT+vl/
Q6A50ZpzojNd4pqDPe7DpZ9WPpJM4n2irL2ewjHE7SEiy/kmj0k1yazVGegWwehZ
rNf3EfAhf1KPCgET8Her+VGpKMdrZ36mNeSbIQkSmHsVHefUuoKx/TDkz6zbQH6M
CDFO2whAPQvoLTN63zs3JF1g3OBsmkurMe5b+UlooN5sy+Y00FRhJj6emgiJWKsG
hcA6yonOizbOu1+suixoxMSXLQqSWUy/YDQoafp1UqUqG3Ccq5qH5+QQxx3rN30/
x29kjpKxk22/JrgRJdH7eWuXZ51VMtqQZ6ub/8CY82X2xuqnHlmfoENNVRd6EJTR
r9PqM6vZTNTYN496sJlUMryGvCbCno6ISERs3PnYXTqHQRGEgjuFAePTxOlCXdVP
K3DxVvfO/s2UMah6q1EobCf4vq4zCI8IO1YieL0isgL2td2a2Segc+FKoc0Xxd96
HW0tBiviMnFMkjT11X70kB2LOKlzRPrPk4KFUkfyLjjUw+Miftc36McmS2cP2nvX
yZk5k7bM5QkAXAUHmP3Fbme5DgieyxuvBORex04K6SP9LMQD1UXWb5+cRVQw2DF0
055TLgatBv7CJKZ9P2sr2WbdJg2Pvkiw18mNYL5LwGcL9QI+yGUpEukCO63fUzoZ
dsdrpn4cF8LrArNMA5GUUYGudxDmQHF0S/Z9nWqdHMFPNAFsTB4e5Ge2wZHk/bUh
gF+yTVaHaKkkh2tpVMgo6jDCViK2XsUyYwEM+D14x/wX/khcptTLJrjHIFuF119o
gD1Qv/qGu4+WrgBNIrsDLsaiXNicfEYzFeC34VRKxJv6s4RN4xvxLN6s3PehbumB
fdJcnrJQ+DdXs7OQmt5+bdjwn7itV6vJAXAiclI7KEwrfE3wDXsJ1bYKJp7zgLR6
hA4Bs/730ucHBsbXv0Y3GQ0TjoFQcWN9FNYPzwHJsK4lwP3bJD66bK0qXaja94jR
oxdRGS9GH6WHSWw+cnJHgp23PJZIapd+zi+iw0owKj5deKbCR+D1gO+UI1kjZheg
qqz2FQxWS73q5mZjb/bCnq1mK8MPZVBpetlLt611ZZsSSrT+t8M8nKRWFRXep0kL
sr0takF1vypfjW+AjIvZyDVHoXE8dl/wkpSg819Ak/4bPrm4aWotLn40Z94FH7Ik
rYrzy34o/LhAygiBWcxx3a5BS7AaTYONHMDajDZOKAJE+VPLF0LZJnXQNIK+p9nK
G8ilMLyjijC495xjT80xFxSKv3j6rYCp1gC+v2PUdBMd/vbB6a574Evve263Y5EE
I2qcGJfIfFa3C9YiaAq+Pj27jCUzXe36XCj1j5E+Rbq5Cdx77AnLEraM21WaUVrH
Pl8chSYZdVS9o9cakzuVF6s+q3Yw5YtM8jliHbNDJOvAUU5KT2q8eiwcU/M7Kbuo
rr3u1Ic2OjuPj1xNiePK8P/6tbnIDFkDT969TAPskaou01jOoZ0tV91FDvAHQn47
NSYdDJbKS0hMnZRSxZL2pJxwJM3L1k00gpELfBRCe20MJ92RiQHP9a9K81xyrDa5
CmZGM/AMr/hBdGCcD9ZPQ3Xue5Au1Pi7jTS6d0IyCusd6q7CWk8tAU/9x2bJ84VV
00fIUEyQUFAwDGxJDNA3UckpTkfHzeBUGbHvJj/fo1e/NZU9NKPPjWmnIHKc5FbV
Sg9r0gxo+a1Ee08BQFFEDC8lTAlojvOw0HuWZO6Op1Pe5HiH+LXbAFnUVLbq/Hya
TxN5m/g6//16Jvi0lNugsx3EsrhIlQB7nHZRjM8w+AulU0600qSvYMkypyfmFDfp
3rXmqBdY2cA1FVYuBGHgcPYNkqJqyGRXvHb1ddQLvY3XMr9FGbGrbfy8ZJHUBPoj
FgjiZy8snoi3hHgJZxqvn0uJtYQ9UCEPMoAh40GdwDMdm0rW9syJ8sQGGGq7DDdz
3mk/iX2CCQ3BJgvtqt6t1YhqG/IsLCv29wlTNDwvm64lxDMw2TNUK6LWncG/d2/y
Cq/AgjK6ceBoJ70o1DKTUhk3bt8SSC9o/A5vpYIYHKE3qi/sh/5H3peD94CzneZT
oyJtk2mEJ5bYthLWbiameTTmpNI1abAjQdL5pMmOrBfasD1WKgQRgPft43EnIDN5
GdZ7HsIWKfBiGt1kZwfcHglFQOhIKzqU6keoVQbro2mqHj84DMwgltop3BieNJXy
X5VTrZc90Hj6innPDxT5nXISqZpiYP6489RIEOCNgLnBDYeyUeBq80h1LzbXVC0t
J1d6TTx2WwugxkORuWeLolxGhZyTPScS0l26PE5LTJl2E9V/EVKCk2c6cKQiPY/c
ITNjkf8D5xnJiyFN/quV24p6V7F94n7mJSN30ExieoVW6tYjO5jzCBb7kgwuX5pC
eajhgbTOMURpKoy4IM6SE6Gf//J0qUleR8C1JsPlII+hfI8ET1I6M+Hj/hBXq5ti
fpDDIhHQPkcxO5KRM2osZMJ23HMqRSTvYeCSfktf7P0ZmWznsriYUm6V7JcGSDhe
gEFWtUA9iknuE1pQJwld534JzlIX55ykmBwglmZltpRMAd8V7mY0VA9FL0YP/7R/
UdaIu+IKFFQM8EqdYJq9TLzZ1eTZhnZHIrry7euEJnSKGWo5Uy7PNQsWKpsbPrK4
6QV94tdVAzLgDNPLmjfvUKxh0LIfDYcRceI9MplF0X1FLnVpFshjkqIHUwnVrN6E
768A5yz9998uHM3R7DxVjCa4AcGJSCIIj9sftNmFF7Gr4St3LCOdZjgBO0keW/be
pQpAIs/4Zoj5iXrd2+iUSNRO0H04YCFVrSxAQo8l7A3MMYjIndCZnCm99exdZUOy
FbystJbcv6BkiQG2g4THloyKwwMnyDmxtjUC55IKq6tebjR5qoy8iSO5ih+vMpNG
1xy42eXxoFsnAGrre8U6DualewqmKIE4maeLF8rJpMi90VFcWzwuWEAgsrkYCMcW
Ax6gYzy5kJmbVW0BBHun7fuJYBmqtjzQP84Y1N3jicsZq8vvH6lokB3sy7JdXTWy
tKwe7XqX3L4P4WO04/adm+iOqca6MZajB0Usz6rwPrDxGQwcUSbLgxjwMJXFZEKp
ahLycQReOCU3+yRN/40CVWiV/mLzmhCQyLAokNsvocs2r/hti6ZDxK85DmkLOSSg
yddwUUfIr45bboBiIXysLzVOkoTudMDz7noxbjHGyGw1p1PKGBwdHCUVUNkK+LKH
sbFycd8WyMP9h6Hcbe/MujePoe/OkydOhVSGRm/cJzisPLPr1fNj+k+D2ZR0+iRU
0SXsS2VofSi6mSo92ZdUNLb963WBU+geKZSUEjTUNFq+sp6irnkdoJgiI+NtGkQO
qk1IEWcaDPJ84ZNitRo+m0CWl5R37jWsw+rf7J0nJIUVy49rvm3EDs1dWPVS4uk+
s3Jbm8TReT49G7PNcR+4GDKE7tvbvIkqZI4yIlvFSW3dNFIrfkW7Xj1TyUoERhg9
Uw/I42kqepywhht0qYM4+JqpZKP4bWmybmOaOkk5c1RjVzxPsMvazsSmTmGUDmEh
O/KoizVIwanzuE5nWPIFURE4DZ7ywGO/tOTyF/lwFIECixeYzHK9xilQY20zLDqt
bMBayA/v+U5KRa3UPtj5yasrY6LfGK9p1xWa/gEtb0NvRr24DUxe9ha6XHCGOONj
oQo/l2o41yihqD0O4tcQdQ1qsMEu8naGhaEy+3lfn12st+LVrYGRAkxrEbEiUHd7
bz7n4Vbr+rCTPr3LCEhZcMkZDJgeDen89j6NXpAD9J8khcc16DNl80so8NXljIhH
6sR5b0uw7DXH+DkFoTFjFk2DG9pNOY8SsQFtuHtPzn81dwaHhhA3JkxqPMqNcxV8
6NtWeQ/HAYxQw/wb1mRf8XqdESlKM+KISfF7oYlKB1XgDGYkKyQLZg2Eytu8Zgqc
yJs1WuoUvsCB/6H4k4hwHeErCgpNBRmjwct1ZSflRUdAYfeJLYRxgpj0wWcow0Sp
N/e0rxAUG3P+c9c8KSdFWn9B9ZXNxj0g26FTXd7NzGWdmvyf04BeuOYbeE0iWdMN
bBuNuQERGJ7uNxH0iDrcsrc8/hBTlU5dnGG01ieC5E4+viC45sc/qWLwovtu0n66
dLcfgKZ0AQw8mV3qrWk5C3pVx27NRDDyZX/TrNEyIYOFrVJpTqvEsULQEXDBc912
waxyrKt2bXra+jMSRIHmWPUAG6UCPk01HnV5QeqljWSuu5xN64aQaT7+u2Ico5ee
JXFHeINkW/GfOyZulArPkENEQWEm1yOxDUz1+VUJgEzhWB7bYnzO/VD/6kac/OYi
UTTySbaQni8A/blgqsI2joYyK/zRZ5XjnNOI6/oyYgveJXn9CXWAf+FcS2FmBxw8
lgd9v/mhPV7HEZp23YXJSkunfcOzXaxL9dg6MzTnATAFxH40BIzD27R0oDvYollm
QJ5m5BUvpDUDjHm+6GDZY+y7JI1td1krkW6aAVe4DbCA4k72rlds4gY/uzwuloZk
wewuzPmXLGbrSyHza7hd4cnH6QeVUfx+Lvmf2Ynu5dEPnu1Yle5EH6NqbhAMOvJN
+NINrCWxLKsQTFujfaw2DDYQPcleeYfhTH50DGd7ulcUmNAHIHm5dQ/iFD/n5I2W
zxcM1DGBX5vKliWSUIKkTBBThwo+wBe6v5hzQj0/EW3RYsQMppUBvbZYMOMaMK4X
YBeOX2I7wpo8zjmOKyr7HtI0lib4tUht6JkCXk8u3ZogwpjZfTgahQV+v0AtLdKZ
cGAnRH/lVhzuqq2FBtpIueT2dqq+CzeFdrN9kfzg0STsdO/mTf1BTSkgog8ZlcrV
8GJnkk/abuS/7KqhT5L2odwTgDYX13CGxLgPhZWHN4fz4TScNBk30w646PteVfMq
i3afWPM6mU2gi7bGFSalXYnW50x3GIB7B+FxyEOmehD3sJ0dEKBWgr+C6bQyKiog
Mw9/5SmK0CmJXtnllKRY34VZnVZ/cc8IonScM/0bqI9OxZM4aoNqjrNTpUtLL9lI
+oI5L5KxXEwl/+mErOWLOUDOp0w+k/BKhOUwoe6ebrgwGfD4RTJkNYo/GO+J1gen
iuETwkB5xL2pxh2NGowT7sqVlGgPAUeyf1HV97kphnOa5vIMC0lxx+7qGlolJP7J
X77Lq3JAnnNz3/Uk++zFxoG63Oar/+vp0FTnn+8CuFPjn/i9ZMEK6jc+0bhjRlot
RX00dekxZcp538mkPtrfEAprfyG5W28vu6PRBvHzVXoeYrBzpF1/ib87sqG7wpN7
fMVjutaMWgxK0wxAD5YgWZklBoRybHRQZqNC6/nkl59IFYxHyJrhgOcfiU9KFHkg
l1V2MPFg1mWxfHgMqOYpiT9by6wf5j1IW7K3u+0J/ZNVUKZtRsiDgP6UzGY/fv+S
6aFHUftHNb/c/sXo8+wpMQ5JsirBK6xqr4gWB2S/GHbeHx+b5g64TUAbjyaLgj4J
2X7byE3ywKXZskKu+eR+Kfa5x45xxmC8BKZm/UN3DFbyJgLeCe27dUduU1HT0Lpp
e1h1nXN7Wn7ekdNPmkGL11MzQftSlI13Y1Mowkrn/GWNXLEpzUXEOMfLsrIQiISC
gLtJGaDss7veynbxWgi0VnOvDvKyePyn331S5gMGiBilNz8V7ktl3FGeXoMSWuyo
NB724HUofGKL2O8rHaVBV2LGN5HP/p5CKSrYYeN5xck87Z5r+jRnXnom+L90+SmO
T/a9TzyxGtOFgMT2ZLQoRd+QjD87GzyeB86Au06MCxMjUkgBBnpVDTes2v6qvBSd
G2ycy7pe1yKeXQV+ur64bFCwHewN4oLkeg7l59uKCOC9Dl9ilUCHo7cGIao67ClT
1UtPIOvMaU5aGS/OWXrQ4ExwfK2j7k6XNZK+SOv5Ll8TaIJVGgAD51IuQjBTgz/d
dGMjOSroNH16wEGPdOLIiPvcatLA9J4KPPasc44nXz3mc/WXwuufrWTL3rrRu2Tb
PUPNIqmF79mkhptKQXTP1PHLIMahun/C+kaTBCi0vNXTSbwp2lbBq2h9m4IuEuD2
X0brhM4f/D6X9V6Wfvyx2nhE0KChOoYKxtVw1E9ktsN4KeYzh9EXkMi+EorHg6bt
71AWStdt9e4sEYKG62OGqslrhnclWVfLTv+FFW+WvkxyX08NURFn1lWtKVKxj4Tk
/s4SDEPEmsoszWgTMhoswt64honpnRQaLVVKERUC6zr8/KW7O8bxk4ADeeWJHJKA
P7gSCq2jUMiRBnLP9RQGT5T0iOQKh61PPMPnS/xvd8ddJmtvUE11RQlASx+7w2CF
qjac+ekQh369LRJXgMHMhZohqnJHx53TXeE8cgTRTI6dnwkl/KHtbHS+iWXnAwoY
/2dGu2uXMCKPkdKzQd3k+cp8sd+yE42SJcJgIX9NkLNWHrsnoRA8SIDwT3rFJSDe
PZlPmrC1kdLGBswrcVusHK2tHfHgQ0q7ry2QY24wYAj52TXrtOOFsS0n1KkVy2R8
LwuNXvc81fi1a4D0kW10sOQy66mMg+xSWrWZSTaq4cDkzmmUI5mPqS60rVLl+7G6
jOHFhlCpiu6y7vF1Dc4DnYRdFoF6luCv9jeXCSr5JCGFVi+mWDyDTVNpq3CGyDSt
yZxNCEw5KohFkiTZS5xs00aSd7IkebakdW6pGZ9TGCyS2qsmFZUtl9GRW+Cm8xqL
T1NFLQ84F0PrQR4PpZTq34oeq6A4kIYOnGVg2FNDW68JklrHALyLiTjcLWmN9ZjY
fBw2ns6/tLwJ8IxOF+dCJtTfiOYUanAshPOIbmOdCh5SY82V2qrFqZ8LfCedgrg+
vsy345He613MQmQjwMCxYlhWR1PbaQ1fMucSUeRLgUwIeGhYgvo2bef1huhR3nVX
WfbGKv51vp1Nxswi9HpxxHOHu5thDH2cxruq+SEY4lUKiZDV14+q1a5h1T7lStR3
cX+4FWKMc0jm/oAmN5sVXX10nWTplYC/OLN+OIs7Cyt7oL5FJ32DkOQ+HLN1m8/O
HTkxPGxTpA0Q78PfUkekgvK++rbkSzXh/TyEOZtwPHVSnzqyPJIju30zd4ba+PFa
IMDCFLIGuk+BgbLKotPH2MJ2XXp6UbPkP9ZsUi7VA9IkQJjxNGey0MeGjQ4mK/Y/
gE1PEjZfDjPrvKS/e7KcblC5giZ+eFWtg0XHW+85rZNbKHMPjOZbSNAamzZtZdRh
elE6sWLTnH6Xz3XgLxoSpAd5LooyogW3RNVODoAoHfT4+PR7oma7CLeBBt5gZmUf
ahRMg2hr7z6dCZDtXB3obwcXgejHhHyZAqz5FTeZaEilfOWr2SgluRM+wfHk8yOP
eSxTJPiUdYizBsMCnETFu9s12r1fmUqZc2tf5j2efcNxclZRDoLUkIOFsfwDdStV
Eh3Pp400J/Z2Z+bNizzIICXoVT8wi4wfUkDgMMkzLypnpnivbrsn4UKWdmK7Tru/
ELruvnGixvewybFx1KHl3rubD496PsZnE4BbyCyy9m3vRzqhb6rKmUuvost5zWL3
DW4mDs4BNRbl6pIWZrVhM/waSPM88s4yhKf+lknSxezkdUIgnL38rNJEZo9ljRnr
VyVt8sybdMZ/1mAaxnoMfiuMUi1IGtnv/H8tWLevqx879tnQZ8mzvcMIKsXDjpP9
u1GPD9TKImNyOqh6K3yPQM9drbRNouWZkaDZVkolDkHidp+41Eixj6X/wYqLa1LW
owzMQ4wNaPoYDqmYsPk5cXpBe12Ul0aO1WaWIE2a+/pl6uUw0BjzFRKuxnOSfq7B
vs+VfTv61JUFgKzjzwLPACcbx+Z4YTjewNP58E3ZEsMaz2EFYYNxjBBeg7gtBbNi
F2czKN8Dc/qFkXNd2S5rrJ9DdD4shrPh/Tng9vvAN4lbfxvI61snfcPiPG56c6eU
WX63+9Bpk/SV5nSQY2G8lvZsBKDPWJqfnTIyeknOG0okEAayOLhS9ogIJSY4CbyX
d4ZXCdBtIh3dbgCSUzArrIdcIyO6EDqRs2RrWf/L6H6lA1OctZR6cYgDuSOLrBWh
sksnwBSvuJv9KtBnjfFWN7AjajwbguaDOLqojoT3+zNYxqpyr4QYVclQZNCwU13q
RgJz6Q/p2yxwmLnO9WhaxhxOCZ4coOjiZsqFxjWiMFh9pSrZaUYX+lcyp67x3pji
s2zKd5HfT/9F4VJ1ShtDW04bmlyfiYtTpcLx5R2jZMw3dATFmVqsJgnh5E4nK7ZN
NO/FhpxgdNN4OiwlKPGcGo1VI80mx7yzVP4oDr4QuhwSTjHHvjzQ1/l/M+5KhUjP
RKH9GNxo9MgShUpi+CMCUNQKw6YsYoB2cdEq0ltoiYVuHRrMuqzm6ZqavxrFYjB/
4N1xwlBqX39/k8V9Loehe5rL/u7PG4hMbQePqHkFl8IqoOXXZGnZBjwzIa0WbOVA
bEhIpezX6NQ8k5qHCbWDFZb+hl49fZgwzfh5o3GhFeK1n38yaJfA8TZBvrYvxMxZ
4sXRR6eYCRkdYb4TrWmFcRM/Mwq0t3znpMs2KVmRuCbDqGHoEGiUAsRp64wYGxDa
ng7kbPNs9GdrEOrlvscaDgrhlEqQjqjYxEX8Jw/cx056v3coNifIvOozMeikL6L8
nF41v92Haz9ZZuWHWRx0MCRvDRXSjopm5x7rfS/C/A3ZO2vmGbpPWL8+wIRybtNC
PcY90xbTyPPkp6E5el1Porq9J+Yz0LtNP6v69gY7nylvQkpGT1s6l5QnGF6d++9j
caj32/RAJ+kU35MLksAjKAMlW+pG+6iNoFJ46kq0MWsRTbSqhMd7ShmwGS9bNOh2
qh62P0DnXUtze91maAwd/9uAF4j7/cBRy96B2s0qtwwXH4Qo+klFEtFGVp8f2wP5
NxcWIK+rBIWrZ36A/qXuGfR2xT7pG4fwglhPnEF//pKhT9A+2q2VyED5xAFTvUHM
hGL65Qml1aqCE4KMxX5TMDPCupLR2BtHHNjuT5YP8mF2TbY8j2C+QGO5PACIsncC
Z4hCwdNmzEwEctqHxZhwN7sE/B24CdV+n9I2pVpPOFAl3JQMStJBZ832ClSXlB8E
E6vncd4DkYknEu8wb85aftAFKQzYiL1dUTPFTU4Qt4oI8rO4OjsPmYMlnTu/sKNW
wRusniu5GqC6hCIGEHSCRQgvGcAzV2XH0yNLLlR0yA4bAXB2SHs8XSplsJtgQFG7
wzk0g5Hffdg0JxexH/KCfTnblWXN0KrT6MwOtiojIf7aFC0ChzICSycZt9b17HsR
C704DSYhIJEIc7JCNye08NbiCDA/L99GOAm7uTi31JjxpB/uRjV98kE+TyvluMeu
X6iYc3wl0qvGDdZ3nVatcxvhL48Q9Crs5cL30kT9dfr7OoL133WA52oK0tQN1zPn
BWhb3+D7aM61ZjEcVj065fvS8lxkWHMsn+C2VfG0UrBWA8+lvg+9m94WELR1r0eX
Owme786Tsxwp3Pe113aipSVUnGG4s6zfCOlO4DJ/Djkorc8uvJNmsWLgTazmZc7m
jmH/y7Z7JK6EGO8Y19YICc8oHvDsQIDZMX8iY1KE0Cx21vWaSS8ioTR2UwAxhMrF
PdgPUrCSYMoffRWQohg/g+eejzHy0w+Qy7VLaI4R2m+rsOTuCjm2CUrGHcWCrIm1
UWFE3SFbNN6tOV9qUSTZAO2YUHL1vSNkZDS+BOfZ/4SWPk5IU3JKMYXddJOjNr98
np3zWA0yOIAovqs9N9JpAtj41bBq3n4smt7m9SSutK6gzvh/H6QdfZ9F5hkA+WbE
VoAuP2+5s0Ow9vWe63q8o6TZ0FiH8LjbIyUNCAiVxN1TN1dhoQXyxXfJG+N8yiEG
Y5cnQfrxXI1OOyNxpHZm0l5UzyAMrTwiu0DOkdUHgIbBFvd3cFZSNTuKf6lcJXaS
P/g0We71I391W5sk4wnMXvLW7lS37nacGQf11Dr9SJVrMTvbfZvU8FTyTcUjSc+1
BBDuY81mMRF26zSwAJ+LueoT1xEHa9xm9/dlB/NcZX4JILWlXrOzWz2h8nruOL1R
LLqRKr3wlu/p1wH4Ew5XnDP8xIlDc6m7fLEViAVJzDSzFuX7mJdccScvfFTdH7dg
nKomLq8G9UKoLDabbCtr8lPzYnSfRne/CjRiTXiI086L+US4bEg5blwuj1oU4nT/
fdUhdzTe2zjdnVE+Xl2S8t0YysXs3+Z4drWi/t5YfWi4+iGJPt2uOHV/WEmsckv1
o/SV/htDbcPz1K2y+x6bWOGZSaVJ9wfs/ETl26v2WZXvfdyeHLoAafqA8SD6uava
N301K3bPlhMbGdu3BP0/9qtU11NBTa+BgMQjYIi67CDazjMuDf9y4bgKQgaevoVO
oJgfyiLrJUArmNPZ3sRBQlNIJH7veUUMwFpifBAYipidJcl3k5fEIuEbHSZED7nY
hmM4aXXpO22vSFhFgU2AYPP9UiwiBaK7GB4qyt1bWK2xq/T1wHGBu8BGwyn+WDCM
jSwN44fnqTgZuYTGBO4OBJCypVFyFhDBr6t9RXRQ7vWQh/OJBVNJngxfgNeYnoEs
kb5z/UGw9UE4b5U1CYGXLWI78xF2bQozrPz2o76Ow4xUJUwEDDMAHvX5Kg0hx5gw
mec1ODnera9l+6kjp+PktZXDXArRCsTyYg/8mRPexhSEZ+bfcHsUy84pwxS4LOYz
bJq7P0EZI87gY1YgS3yxMVkupCzOJHTutYGCdTUmnMi8PuTDyz6AeauNtJBwpYxw
GDul6b0a6gzZQPEsDcgdU30lY22jIExoKb8JlrO+sip1Fj6cAt3WYRqGbteyDKg7
UkPbCC7SQ2gbmCNZkNb9RkC7VFvcUdJtg/xmz+z0aGmxxGFjmFgXD6ci6P/GO405
G/npqej66SDTwPwcWXggvEtpFW4Wx9puTSUmMSQcnXsmEYGucm96zYgmOQQ/ovnl
LBW75wq53wbwnmYohoIcXd7I3j7E0HDYllhuEg/uOKmIFwKK+uCo2Z58sWjCmHfd
qOkgxx3DYYGo8WWy64FCBkgfcxGy3FfmkGPnZ2M4zIiZ+4eTwAh3Plewfx9AFG9R
RwC+dVOS1WbcBOmAng9yLTsu52i6q0sJV/XUs+C3wHWeDXWNdC7FYceOuOgrrDhE
H44muKHpKj5s4OY3nyOEPPkKiBhFs/pqKdJvyqmz20BGAMX4iFHw//H6EmoWAwKL
aB6EYT5Uro1u00o84Bi0CwqC/MvzHuBr4d/PJOyEmJqS9IUoO8BComDxEl9RJGMN
WTMLf/0xF/Sqq5aEpew9Uutjvo8L21hxFjfPqxR4fhRABqBBBonXdEpFBJlvidtd
tgmGc1Fyi03rs3HJqO0ZUPLLavXf6w4W/w/mnj0CKyc54yrmgAg2lA58FteQ7Jno
1hgs/7FaiSMLWTQNw0JXFiANWVLbrWJd22WWzmUTxVVbpqbntgOU9s9h5xd3UZIU
UAC+GcEn8GpdfXifzK0av0iqu1IWPDduT+xtSSOmP2MnPde1bxrU8IY5t26gUV2F
3gK+aIha8nLt1yCnWt/5FF92gmxW16ZxGf9NicM4Be2559JDqdZGnH06xmfZ56Os
6Tb7PQhUAhfcu6cFY4Wlzmq6WfTd5GNAWSIURZTquvYRiQ0iTtxfVSeDbEt3MzMz
KyPQu4P1Rg0QpzfbNlxuS71M1uXQbN6MKERtqfGrGUWvsgq13NBKxgA7WiUumqs6
YnoV7QupY0HP4HP/JxHqzmpMSP+9aNnJpFeuykX0KG2T8iOYcYdCP2CXXAnEwyWP
vv9TsDnNbnDwAhllnif63YXzt6s0ojybXJyJ+yJm+ryKzfodq2/JhTbmJgmPvcj/
mW0cooncbIpjFgr2NDnctg/d+McEBVYHxwvBB+uZ0Zjtd96yz5IzGp3If6Nc6Ksa
xD8fzSoZ/qCnMlluw9IWqklTCOz0A8jsdC5F4xtjubEhMCyzY/q1CpofvqzyXYYh
ANV4cgkWmkeu90DqVmpTAMoXrh+a7e2P721zak/lJ2Kg96yFoGXgdDHHkTlkJEvc
ObHICbmRHXltx3G2cscfItoQ2VuNOVZFV8SK7PumrPESIg68MzXNHfBDYfsijmaZ
2qcfVjrU4iw63ReyhWS+0THqztsmZq3T9eRBFtz1Lh+83cG/dRoFtbXKoqpWHfCq
FK2uOIg3/bQGcXYRUi6rT4lOFvK+1hOT3IOJkKOYWC3dIPV4lS0+W861T7Nm6oos
DsVoc7e6iD0wqE1vTWarlI7uy9ACUwhHfKM4Ecs2OWOLjMGM8GZIR/Hxv7Onp2iV
eYP6UsSc9ZJ2FS0ak7cqqe0GE6vgjYuUDQaTzEneV+w9fpUFiI3w35CFZikynto0
vmXetgZyQC20iOskxR8QmZXlMmJ0OuRrCJxaT3ihxtecNoqaX/WV064ESAZIKb3R
GKkNKTrKGTr7U5J1KYylR00HhJnDDoWjyynR1C/OduW/2357AJXml5pfatDW5+d4
I29ljtFeU7muKPnp7KeMal5NU2Bn73RIan6F2XlAYpjyFkmv0pxITtx0WDJDPjLL
tVaRAm0qpr0zWXZqaxS/6DgGgODil/50svqcf6FOgwh/9jeBTrMes74rWFpUDZr9
xLoYD0r0F749GZjy13ZWfZ4NWrK/i4WIGo1P1vtM/8M3hmpuAoyx+yZxTOlVw+sb
xW/r3LtbOQyIGy5TbtLH+yNFKBlhcRB7fFxZhLrsu+vsJYz3crU5c9ljmmdgUSh+
/f4v1OGyTK5Yi8dG2YCuSU2BVfpXnM2My+cCdQdFnJCLSRM4lnLLMeYQCLfNffK5
PFu7R1CSjdR+Gp6Wi19slCDmHE2YvcwMQRXa+ZIMKyi+kGBtx5VcjpMCwnrUqi5p
zfMdwXfQw+22QDJn6tMZ/N324ggqlJBWl5847ZFBtQuqC+9kf9SowUcyNh05K8tp
ECUYkJsVTZx/Nl/ycgTtnFVKmLZ7qRGztzLvTEka+ax8fx1dsMOrHZ0R6/BGDj8Y
eUqjcVuJGrt0YZJG8ZvHlrlprN+C8jhiXflCXYvpklL3StShjPaaaividzw8zKIL
ltMitImnFmSygoVj35rYH60nTyd2+FCxFdW1gCdM7ZFpP0WxvGcGOZvhyVHnRhEr
AAuH0z/qTV6gY068iw/amFZBzMmnudMITcdq4jzW1Ukz44ye9BDdP35NJjUHhDp/
Qn0J02lSGt9maf9eBnOdAxUMbLXve2GIN86vGK8b8SwKoULxo3KOuUHqbrMvcl27
cE24R51Klg1fjOIuEagIt2adBu196gMWFCgCC6MTKWO8+K4NeDZ8pQR3R9B3cozE
cYBoQ/ZqFCfjZzvd5NEe7aq/YHilDwD52p0fWYZ9WmsoxkLuQjd8HvTPKQxslS1G
vgg628R7L7gPu/BMS21nRXPlm28YU3Pz5HUJBzEGi6lVBI2vt9/LlXX8Yi7myMK7
yKukU83v4hvYCUsfe20/5hyExacT0hj18NZgYMEnZvAndNA/v2B5VFKEQWIAva9G
khMPKeJXFBtFIayNdLrYWrMwiqxJQePgh45IhnxtW28xwbbziQ+bY6oz7lQn2kXw
iWgVD0nJqTlk6jZWxKhI1SmWkmgGN/JzI20F2iu9GxntUuKhNVGOyl5ZfEz8muAD
eokbOvavQVTDxyf5siI6KOfVFzMbO4BFkAvu67Oh2MH15ZeqeBBeBwfNQhTp6OI5
ze/LAfnzq9XQYO7agYNrci676+l+fk4C426uO//d7+eZ2qSj4ngUrIMGKWbkEsk+
lhDbcAysyY6eSCpUNPQu03u3NOBbgrRlXeq1uVzM0v85Myt8u1be0QA5WDBsXlmR
B0Fcq5ivMySO2rAt01ZI3rTMe94xWuMlmrlVzjKte9T39mWyx32hI/ywrIbBLoQJ
OPiTd7e1xT5r293n8Qhy3Ehs2GcatoMb15UjPl1evTlBaK4rCKafThLSXQFEvE+0
8nhJe/UfUMmImakuTk18acOVIFxh8tyOHfPv0DTvC2C93VmcCBQsPyrM4FYnSI4N
oeradtWNWemSLIDtUk1Le7mU8a9fhbcE+TB2cPQ7UhtHhebGnx7sevHvOVSqEbXG
GKzKidPZzMThchynaxyT8Nt2HxsTLLTLimGFewnheFDN00Fk5nLnA+LWe5OT6URw
iBI2v5tlC0LTKDQyPmbh6PoZcCBSMyjhLMW2JWw1AuxDbLiynKNNGtOkbOux+OT0
XyEltcENLr2Fq0gYUEtrIJYSs8ktA122gF3H2hqUFu825/ltC4Cq3a8YkTkHOTOg
YqHYLE5pluRJbkkl9e0ksyl0r5jxoK8ZFGORIARjHtRC1wNa890IsZ4zPIOJt9h/
69oJp2JtK6UsK6irWAbV21YwgHq6Oq23XaXP3nREygO5PaDiQPT7eYs7b7V6oWJe
4jSrJETdJhdOyCZxM8Hcc8OHKolEwtmRyfMVIwcEKlG8x3yize1olH0R4ZhaQt0z
L6B7YpXyNqixO3uUfo+TGKRvm1pJemycd8UjFX4aHouC1Iy/nKn8OTUjwvkmhdQQ
Sbv0P9gLY6Cn6cD9SAvoYs+T6PkYyoG97W2hAPK+Yg3tuY99ynT7Rh2XfrxOwPWu
NmEzbsoZEKYd7/gN9HjpmRHjurDy4OntMmpso6RxLC7i76H3+eFS++gXlARavbhJ
HvviOZvbggKdSk2rFwu6xlvV5SVWR4R4Qr1CTDaWpBil2PbA75bl/XaJEMoFWkSh
+dD6NMidtLhOll/Elb2eh4N1AjGrjV+9upqYxQwliLDYgBFtZT4dnTVbHva/3qxY
V0TtXEPt4bFW/GkhrSnm8sJJGUKei7KoiDKjHBNdJTrgH+JkwbKWjDDr7QT+QK+r
ECfHKPGifhXpr6hugMx39TRxoOR/41cc1KlJGsbEZ0+bnBgnR82bfnXXTJjyO6rs
YLlcCHFk7yf0HJPKESVX5HCri6p6WGyg6fHxIKnK6jY0pO0VezfYfvFcM2cB48Nx
cPcnqcTK7u9ti/TCHXFjFL5n92mgPXJ8/xPBttgl7q/9SOdjVhSS6JZZ8NTNaEI8
GZ7wzanaiNm0qPMzBgEJGK5bkl8ddVOWbKmabLF5l7Wp6zubsbFkdRW4LoeuOd2T
1YSdHwkzqrBd2/3tFDaR3rINbaOT/s6je0aCsAKxV4qCJ3nXl2W0yRwrEmsfMwUR
83GJLENpaM4yrUrUoE1aM6YLl4NZlfiDXwhTj2jsrCBSAa9TI74hrr94aPbKWgW7
eaIZMLkv2rKVIGOQuDJy3MonUOEgbLlvdF2GgWa6Q39AU673gBASqI5ixSLNRzEY
WCA1EjcLD5+vVEB5kR8uf4Z9wKYQ8Bbqg2EFNkgX2vgq6tg0KJEv6RgJUDo6KnH/
u36BP+46H9278TcQ99sSHIDkClhAZsQtvSyOvrn1EBu7KTTOqCmIluGBTNBRSmEc
LLiAHdx9T7pXhE+Cp69bN89iZpTvttZZFB+3YjHQDENpMdXUC2DDFEJ4d8Hyrcdg
EYn8xLKozeh5EpPoCCdj74JER/LCx/wHdlGR/UqDXdxsipL7sXTCnD6ipPLDngiQ
VvOW+L7Wy+3qryD6lNypSK5A8fQvgM9dqb1CL+hSGtid1BxWxqfssMlsP1c0eB3K
RBbpN5YDdHjDWMecArdDiroVtfGDtNx5y5U8vhIiZbByYP/z005oKsAOcshxEt5m
ZrdYebKLajyIYz6zK0NsdQDKYHLAwSnKbpAPoeKI2Ty4VDfyUpAoxB+VJMFoi+s2
WrB4emq/PSwbmxpxW/TnvIvGPh0Kj4gzlkSvgQqRiy2sTsntAKUVyg9T0MRdZ6U/
GEycg07aGlFu6afBUFiyl9GkHGse3agdR868T7wC7K+AfXE9qFQqOU/3gzjjfL+C
DhC7vQlzgavRf6pRso69dMM0hDe6LLGN3AKd4ymnpbnFM9pqbiSDdLWG2hE1lR18
XMX7mOBdBc8bYHhqDUFTe1iW0a+UTkPbxf9VHg7DR3OPvH3KdPk7wLyrQI/jbwx7
WF4EUnvDtpfmuu2w51ZPeQ+1moVsYxmbCMtbHea6cfX1ks224vOexlvTuPr09WMD
8QEVArnwkr89IstFTWWRD9xu5iCDmlrp6oHj4s/9OqX/O2DmWisW6zsFGkE/Htnf
m0LvVhDCKlWHChnE2Dm7xBnaBTDN6wrSkhcqn6/RjZK9TPauDtoilOhoN53F2X7E
H/j3kCa8bZZCkXBUaleEdtiyOEMPl48OjEPT8JFN2rW4mPv4MkOdZRlCV/U8bYpH
xr/YiGAXL82zYRFm4VweVkuA4wY9LlGrekyXzJJtmYki6kDSUMMY+2MoY3PFxhCj
ACGSFmjwyDS+uOPustztpbyQzm/T/1zvqyQor8Q52+ixK5XbBTnpw8axOUAp6bH6
KG83mMy+cQd51twNM70rASjlNaApLoFkJsqyu/8elDoCKqz2oan95daheHHWR15W
B4iSpYpP3H9HG+R6gvAtFszaMD0ZZK+fmGdtuIl5isd797ElKCZwh00RCyPmlUps
jmfAboadaUA7cfI4HFAOeZ49ApSJzwXsbKrbTqtLPSPkEbZE0gvZk7Pk+og1E8dH
0Vo7eIsOqe4TDnYO4sNGmZaDB6CdzLzTGfuRQwhBkcBskNGhyyd62UoijXd+nxHh
0Q7O/CqSuEb9r4sZSH80GAAzy28AjVCLvo+Sbi0zLp38oBw/FCtscRHd+Q4+ESqv
FhTv/871rZ8RQYMzRF1o55fhHbqBvwmMSaW/ogVNT7UEVWTqbdfiRoiZNqaWUrgI
kcZOl7GqcGDn3GWF2vH0Cugzuny9Qk4v3rjCGDKHjzWftt01Nq6t9ve3qbGqXWOl
uw8G3fwO3fF/5IAZ9lbrUfOg82IlOt1VLxHoA8qBa0ThfOTFoYCM4WGttB5GTPyz
cxISb0DQGQ/8ZzyIlc95MGak3yCO9uvgS+ZKdyao1sqFHocM/i1vx28pSO+u9yXl
veLecS7kuHOhlauN4mj0VlLEhc+0yHk3uxHb3Z5XPPD/o4aWeQ9Onc4UsTOabIyX
qnVe72rL55YrBX6bT/qep9i9gkdvlvLMuTcLZDPr7EQrtdpKePBGHPqAhh5cVaSC
ZgU7xOINWzd6rEgM3b8D8jxEiBO9/fwg46OosABBeYbomcii+DG2AaQJj0DvWNTs
ywjDJ+5HDo5MAW4L7Oo2lGpPbBllOTvfUL/FYdH9lf0Fl7yizdYl2zUQfJ/2TxqS
9aQ/7rBSj63ssjZBCR0QNLSBC1CclVckc/PoaSiHg2C8tAY0qgjg2+YyuX2hZiRw
AGXLxUYCOK8YwsKWD6B+BDzkkg8KZns4gAEXFvrNL0jmcobRCW1dg5DPejw3Lpjl
f/1cGwXbgKzLbJVsKGY3aBk8nmMc7+foeQzZ1xUrf6xSuw8k+JWgSpd6OP44Dy1o
nidxz4iKSM/Jtg5Zf2PyC1dmWlD1L/XPfaTknBApTi3EAprS6YHZ/HKIZ+Ywu9w8
G1RuCKkfigR+G2Nr1nFlg97r4SQWU+jC/FsXOxYpEKLvEywyGolnwRcsGtK9kghu
0P+WoVJXhnESrlxKJtJx5RHuyBxmh0/1vRoPkb4opRpKREMZGA1g7+knHqc5WyVc
ULP4WhRLDKQMLIwg22YyxbshSGjY0+RyEtwsmbNGnNrvx8P9afpeVluNKLUyoZ/q
XVWMvs6Ce9FGNyRHUCsTfjdxCnl8GHJDkEqBZnzdaAYP9xsHqdrm9sXu5s5mbcGK
Nakr7WvOcZYevMFQAZYquUKK98GGeGbCQpTUDco6uuJ/ZXWa4x8/scQoavh3U/wB
tvSFfsJ3o+rzvlO3ghmHbjjeOklzyTTRJHHUwO1cGQ0Ll9mSpFroXVQ09md1KQp3
JnS9QodsG3H/PwoicLqcz1ppgKl8zij5V/JthavolPEf6cSouQKfwwUNEbWemccU
W+aQfTAIiRo3c5HCIXv9Wx+XXIN/Wo9EbsKBpFTxPzU9l4qhf+QWfoXGtG8hHT5Q
xaRiOiY20VUYM3AQCgFhcqVyVw8I5i0r5mah3UYJovX1zcTN2fAdWPoe8jTTLPqo
M/8N8kiFCkqOs6X2foCyRmQbRagS5688v/rY7qTdMhhh9XpCP0WP1EWtnzG2PBN+
8uugfT/cAgMpXeug3zNbY8dPM0/4IobKbhARvE52iw0EHB/07OTwxs7/0zk2SUj7
zmSeFqDpNCSBK7jTZ4HEX3ZL0//LbOERwLRU40JvfTYTxC5ThJfL0mHsVJO/fO89
mn/Kn0paM4hpt5LInXbK2AKRNuQ5q2gni0a+1Fr2DHvX7/tWwA3G7DfBEi70WADa
VYGkyb7LRvzhODHz6dfokwXM59O6WlXQzSkizMSBab07FV3VfWrFQLrqRAHHnw/Q
RsU1a7nZ3cE8gMlZj/Cs0ApeDDCjNVr2XbcuxhuT8jRank/j59VFwTQfOt6pGLpj
u1pu6oxGer7K9duifPrqlV3+V83RXwGwgugI1Uspr/d+mDqNBuKXxeqQCGQFKjxm
yiMI9abwbtCiByyqbLCS2byhHwGTM9+9MJgoiF5Y9xMKLKl5LNRY4XgcpRKMJwgA
JVylWH1kHM/B3fFL036S4r8qv99lltwqWuIIb8e5Af2jcwWabUZfl+s7i1NKUJYE
kziTVq0dumOhxcVzM4gMTfCivyQ0cMrhyfzE6SY7/YWNI7SCvhVijfpcrqHLhD6Z
gYcacfGPvYxup1iBa1UO6EQu0saSgWhqWktALf3fLNiTUOTMYks4NCJfEE87IVrg
B7BqQvZSMwbADlreeFlDZ/26GIUsbcbIlSKK1OOj2ewaTpY5AZqnrehn0zu3GPYV
qduMF0vxX2DnZQ+EUsFCerLoVSBQ2UsRkOgA/58mHtalS2TiOlUgW8DTQE92Mks/
Gq7FsLfSQucICgc/heYAg1FShXI7nSKyp61pFwXIyGofc4+ucND9ABnxWIJyt8DL
7ns0nPrm+CGBVp/zMqGhNRKHFAJGX6/j822Q50tnUnES5R4/+tfPUklAdVGuWEZ8
k8VGztOvMrNEMyDjK9cfPkuOP8Z9DjHztTIcldoYTGYELzG0ItIuobSFsa6ewnIH
aHwFWXkOk5nIYY7WLwy7Riia+c1asGJ56Q5WdCZBQbb7JRcezTqmcbwUTy6b4kWs
VeKkXVr7gjiGAIsv/DUyqFJAUAO6i24+cmqLBTaUHYBI6mbIAtnpGVhn+t6zHMUd
5r3WUOwsNQ6ONv8qujdsXLevZtzmnWYDDFMIzeecx2+EA4zQcvXV26Z2Us+wLIzK
nRDKb1huamyPazcPgX5738+WuCqi0hBbgEWiixUAnarMU/x85cq7GCEVaqlSg0m/
kk2stHE5IWZA2BZDbfukCGD0n6hgsQzXQoEK7HgqqBuMQzrmkno+9cl9fod0onWO
0ql9f+HYyATmiZ35UNtKuO9bD4y7aEb8fpKU1CFIrqspPnTv/GqdmLyg5OAaFjto
PiHFkd6L2j9uZYNZjmkz306J/OhY5GVcOUzO7nOHQhT57tWZFse1epEQcHKPUnOn
/8XhCQV9mhEuIeOwK4LJMMoUw1izGDKfvE56ULwjLb6Rb+WwhAuKuSIDulhd2kHo
5hIzOfhcQI1nGyKkozEvL1HYtFoi5faxY/BljLLP8NkgyH75rVP4PWH8bmnpe0DQ
kBshmcUSWJMKKu6ri0OdkrxoZP6L/dFj0gXm3ap+TGBUspzwU/djnMciLh3DoYGO
gIEYiJ4fiKCb072J0t4TDS4gODHQJZmVzb5L252ijsC/T61quFdLW3nD3d7csFhy
HCFHTHk5CRIzCpyQvsUb0X45W1cmfOIhMJhnBnTbZ9k0mHa7pv4RHVkzEdxfHR7P
VfpLK8HPVplqk0OcpXSH84rqWIH24xfLePS29XjCv0ZtE5VV7t3GXt2RNu4ja6w1
iLAE9KQl5wg8RlsMDMW6zKMlzcgLDb0ULcgxstPneYV+2eGfyaRb9YbpBXH9nbz0
4DzUk6oiOjKcCkU7EawDUd1bFE0kM5LBi1me+CD4BYFNsYCzoUzHUM6IYGQeEUZf
yIk31auHO6koHqIUr0SkDWAklws48Z75aNI/I1/k3sgweIbwU6ZSv+1XiR7aWge7
5JZsaOof1AyaW4n4oZugm5siBoPwFjZ21/6nks0e28PLU4PJkD/t6dnZYIi/uOD6
a0lbUPlt9nyO4EXQRoebTjbybEG4+t2mIc2X2O7AUrRUtgkUroaJ5IkadQYBofuR
6rmPMce3txAtl38NdekX+syWM3u5mG6wsKmcagNM1GqGaC7hc/5w7KxJmp2pZf77
dLJxFcatCYZqYgPn8fjKpaTor9boBPSR5lKPqSKjSJrcqtR4A+m3yNnkX2y+It35
6csYvP1p7eWvP0oU+WMcS2fHopDGdJm8Md9IQA1nekWUroPcJFj9gytrNs/6Y8vg
YSBjtWEAhHc+dwxLubx9yHK+0RZ5dM3PpMwNicgKS53HP15IJC3+/euHhfPUlRpY
TFfmstF3OAdUQcD+mez61+tNZUZCRita2wzMDHZH8YORHyqPNcDvUHlRjMCFMZZH
/Jv8YGRAPYcMqK2vrzbLRjNBW35oL5D0WmfJ8kTnxmuo5FoPqtzw+WU4EoS4Ul8U
PbVYrtisS1XIQ/zV0xSKylceDT6wlNomzeI1K9w/iRMlqxt1Vo8qo7PcQ6M5WxW1
zBKEl0wgoq9CCUTXsen7VGU141Yut6JRlHmVmMBSDw51gDN/hq/Pn8e5fBs9pq4T
Rm0u9LDn0W+pcum4u7MtvZNOYDFMsbTkl4eM9023ska/IjIbxmpnrBfJs77Dp9WO
YE1imo5wvVWReWTvzIgqn8zrtFRYEg175JDLDd69Z7aVS1uhmahzPquSAIFDAGCb
gyGE6vwPwPG1I3RqaDxniPI+O+hXv4da2P3xMtbk6peW9IskVzUrurASNKApuyAI
CXvZyDBOE9XI1+jSUDXjgaIgoB2WUKRbCS4OQajwRH5HjFs9gOjhi1MBudXMP2Ds
iVccm8NfMfQdjGFBJbzJTFlyPHdTBhGZzn9IijdqvvNfiijao3HHVjzPpw6xKdjJ
IhcrM5VrkXzJ7qp22mjXQ91sXrYmz2xjMfpZSyjI0cIUe8+yYJEDqqfAiVtDEn8D
u+DNkklzuV+J2m+d0puIGwrdO5fQ3Gi+ruKDQBGzZ3DIxyG8yePntvcGnjWRL01L
inGXmXW6y6vwvU3vwz1UW+JZ1/q4XIepwLUo0LuVhBFmuHhTvE0DtGcLQ+9v14Hm
1ynNWbjpGZoph+NM4w1Itv6GuDwVjuzOxopbOmSro13fY8Wrc9qBwOY2Q2pLNzXJ
r79EZm6eavuKahqEK2w/jVdbjexEglXtTN6p3Y1mmLId/m1Ldgy/3AZxJkkqujxv
aO+YZ2+v1JX3gYNwvW3mBGCr0JgAslSTE+BLm1+2XL1twUG+rS71GbbjWyRJOaXv
sJV0WFIPq/Qbl1vbNfRrT2ZUwQjRnzeX8feFowvmKuPxYr+kle2Byp3VFpoAu2mS
WLuiXKrFedqK5x83U4P4z1YMJbl8VaPW3MWFkfhPCEdwLC2x7ylT5880sPqJ3kzj
W20sAcht+SzL4YzRA5XCM+WoxjRVELlPWz6WbnPPdq1KpFTy654r6njWGbhJBUxX
3/C+bNI04GnGO16TjpslXioy9gC/JDmtLunW+U+ot8W5V3jLyiSq2edH/Q5IUE/y
ZZYkmgDrFXY/qzerxYHF3SLWPb4GazHhNQEtcNGWfVzw3Boso7uy+kfC/Moc61G+
krdiK5+x6f7JarpLeMclkm3Fntbf8DcnOgb/RDSkuH6zvdRGsWgRMhTVCVNcufEs
74MNCDInaTlHN/kvn/l2CLpAx5qAYnYlijrE3SGMY4LrxxlHsiEeW5tmjlJB/jdL
onCSlgHhuOTswXfhf4euqyEbjViJe0+Coi6qNJetfxCCtQh/IfBw61rfNFggO+ca
i3BAYdYWNcFavexOlTMNIocsMs85Frhe3JGQIE+UnuT5lHRQYCQ2Wz5vkiWe5T9h
VbF+lDZOeie+Z7Qloniwhvi9vNZUAgYebrn4PeZPq9mb4dGT3Aupe1BEodjFCnsi
iO1wRB31Ch3cJIC9p07WPqm2r74Oj+s5njgGLerYBj/4cHusz1TElBgY8krwU3y3
WfyxQNnn4kzGaLB+MWWXm0W/rV4Mj11AyQsXGxPGYGypCNUJdN7dX5xIb6r01O82
CsYbfZAGdC4oX2tpjkRRsGdPTZCkOVPOBP+4NjstSeJgaswq8aehdthoWEmzAdq5
HnPq86kphzjovorZopQJ1zyyErOdbV7srDgvrPa/HjYl31HEAtwMUceSu8Tyopyq
ZEBBtN7RXBpK7DRGD18yruzjNooY+Jiq1pU4tyMZmVTRsmL/2MNsV26HCGOSV2tY
UHTFgqH2ydXVAv7k1jfjOzVKcjx1IpzMogWQGLCHvfUupphEEGC68JhQtEUvElpO
AuW+/eQ7tjbWWIPHlkZSUPf0FtLQHYaR0Y5p16XFCRnrqq4pUJrTyEoc1Z8vKaYS
Ur7d/qeQ6GYm9wX55ebueg6hx/LReHliiCRJewYzvcoE5UlAYd4v3vG7kOGtTJeI
cWep/ZTEKp77OJER/9HWrEBP0e4O3IPq70G32NPsTmLLRFEElZtP2dB1YpAf2J0o
QB6IIGVDroiPkf1hmR1hjeEjrOPHfzN9knqPMlNhcfShEr29NzH8OzlDhflUsPgU
L3D63+70ivfEACIEkljyAIklXuGk33w1CltxpTcJVmjuUz0N4RejaVLlrr4tSQt/
O3ytjlR8FelfPdZKzJFkfrH7u7HpoWB1vUHapAvKMlLZvCwIjn58jHgbG+1JThzE
/R0Om5ii5kUkux1+/YqyFgOsMeMOCXMZ8O5DvYsCqWPPGv4dCOULn12N677zPomb
fEvmYKXk+OiI9pOA6UWoUeRfkXkiwqxFMStKiasFfuOvzWCYxHOhG40601Z+kJgi
3Z8EINSdsXELTsfc+WwmWGdEc8KvKO/xSWhNFlSUw5y8+Q2Pn/3bqzTEvLczsgTz
DDlOSnS3JYsgPidd0z67Jw1I0gzpgQ0uCIVM4p5Ic/9PbrbxBNkWB54CYx+4zvgA
bg3rlZcdexF1n0Zbp2AjCTlJQ0C0IfVjgidEbn6kzC9uh4t6etkB2Q0p3B2dXlZ2
4w0+FOOuMtGeFdDBqrA3eieMIdQrnTlP7aye0IwhYIeiRTNq4t92spNMGzk2yc+L
Qi5LCwCbiFGkaAThoWsJ4vDIqgVZw1VsycCCcULCALDHUbv9phLpss+9f7dEUMln
CWXR7IS94KGcilymZkT9t9F1iEUagVKXczL0FtQ0eBct5kEtAR0AVKFWZ+7DvmUn
2MWNdL13MMzT2+EpwwOqD8UF9Fwg2Wqs4GF9lXly+qRbXHyew/NsLR/R3X7QgPcr
SBYANuD7d5DMnyv5Wwow2eWbRQa+nmXDcHjJ+yU/pvJ4Tw0LOxeStekyKBDnyxqT
lJeAIwzH6jqtMuQhF70J3DFvXevmBP4bo2nkgLUO6E2UlNpDdbAgP0weLZUOUNwN
6qqaPQsRO5E5mFFOk0ZosgEG4zLjzbhpowXE7kBntLK7itRKsJkG0xU9PzcMtbtt
6Ph3D9TxGRNvNkrYslFLVxmc8QHHD8ms2A1hLrsLSJFjoN/FO91xpGDfcrrWQQtI
VsFExAe6ouArbV7csR4lEJNVn1TgWK89OZr2Ps97GzNcBs6j1YrhE45GvvMwpzr8
F7tjPJKLIsqJwIOenmIgTJfkl6fSbfNriOudHz2z8bnOzPhfblmaaq/NdtUaqkLp
iD2IrqYk4vznQJIM10NPb9xQh1sBLwaanLJgLEcNehWuWbuaUj+t0CJIJ8ZTiv/s
/4A5/wsFHvzZjhspB02ABR/hWqGRgyfs2ZuIHiL4CL0F3v5tqiqvM0rnSKqTOBOq
dqpW8TopqNsZSxc8mdDrmEKxpLhuVIJBsRst+CEfNNGhM0rr0vjxJhnHLqNb1EGk
stGzil3TQcPS6ROhVkgx25nbvRioVJ8ygqHDllvkBk58tTtgPXbGNNw3Ya1ePHwd
CWv/l5rFjOQutTKC8qSgDBsdhDhIoUyMZa+h03t7/EHKuptJI7iztYILQXnFpdI+
Eiy0V7UdrxgFHvr0vfaVsRdlxAL5qUWrjgXCBLdcyLDlbvM4pLqxqsVGkYqyl+2I
e6wy0W1tedVmB80HH/+X51tRBRYuDEWgbuL6UGbR8myud/pDENC+HFbFvqE4AK8m
j5DJDofXSflZxwbZD2F8nkNdGNn7fsyMuMC9XDwLyTebSOENSthcxxbulEN/6tso
9x63mF11/0Wd2pyMsja4+KEzYj64Ak+fk0qpzTHSJ+j+UqCw2MbTQN/Vp9cp6fHI
ao45spKtJ4IlOBzU2n9lZYwn+LYZDZMJM6OwvgZwoKalrTXmHPX3WMVh8KSearv1
/kt2trGqAP9ABR+ZCKjEgwJ93dA+dA+Yjm1bcYabIau2JO2FCEibs9d00hOWVNHu
roMflBtB/BNW/MeTQqNetEC8Cmh2rQgM6LShzhiWiR4Yw1S6xrdLOadEQsweiZJJ
3RgzqpvXISXQXJ2Tqknp2LfR4GY+18EibIhsYguZCKVL26RLE7J8B+m/QmU4HQSV
UBcqUFl4XCojnepgaTZUIHFYiGzv6rosIWzApaX8B4Wf984x7e68DYcuX3TeZEXD
jfpFZyQDO0jdMwxZE7XOjNCB9pqmEXSPzLjsjKJtOMEn0IhWxP+IykzAA7MKytkd
URZCKrLODjT0Ftf9R+EvXrXAWiq257kAclQccYkKKosOQFNCbCBrmlmkO2oK9nye
hcwNwe64tFQVUed/mKsM23okTaA/BQYPme68Rcb8zMmTJD6LE3pWnJhVJQyjZ9Is
roJ8zE1hv/QIS+2JRpUJ/I4aXntMDBTHfWC1/69tpCcxhtCtHFgHdlwhg/zSarGw
yL1pLcSCQ1jZirsVU/YHqOR2djNu0rpelzKSeEFvm8fA1xKrZrMCVvX6WRJcxndU
DDqgmBi1hNUJrF4c3pHSeaf2tmcKAFdF8+DiH6BH6+oP7a35HiJf/3QPsmDc8CZD
1hpM7l+0GAj1xu32p9xl2Hpl+lBp29KwJ5HlO3wwbVypybvsdT8NmW546MdhQ9hk
5U1PaBwBIcy7IKUCn1ki6ffqhu/9E0YTXHL2c5wtMn6JzbibGuAl0qtutG8FNK7a
316S3Bq+LIu6iaCmGsDHJgj2J09j0dBL5i2jqh7P4Kl9Su5iYaqK9jIfUCyDDBHz
iieSseTWK5uTDGflMXYrdm/DlztfDV/d0rsKM66fqJNOty9kWFhvhIT1ftpX44Cg
QBeQvU9oqnL3o2V1dp1XdBme+o0gbBX4DHBwUGnO+rR9IaG0FXpu7xfS9Nxc3+uT
8OSUYGd6XXnahBHU/C+D0CLciwA7Cluzfy1jUxioV1vPKMsBA5YXHc5BLwDmXRSV
jC2CUtO26syJ/IgK5YADxecUyZakRpk8QacLZVar4vv6ZdnTIsXhpSOsLvGlVgbw
lMAoeYL0wztYxop4iiKyMMJKBQL8ksdIqDiwzV2awS9ACBFDnHs2iaOSGulHiQHo
WbVrA60a0Z/B5EquN0Q+v2EPjt5HrpwppzF0TBRThJ64ypRpHy2u2QU15FR4kFBv
96FNeoz0DjXDPr9FOg9Ml7o9fjytVjWu1ZePe6t349U1AAMpeUdDWZ6pc9c3Lp/V
fFocSLpr6SfQ2Lcq64els/2EcqVBwTAquBhieQGdmkdpb79nqghGdjlpqnfxm1C7
Zsf+O3scCXyEQyKcntus/y4Krb/CDkmtP482Kznykl0BIVlxMYJ+zSoZwWmx+fe8
OuvLLkq+UllakWMWlBlkz7J+6WPXS1DVcpDkioERqe1fKhYk4blbQb71nLecwjst
1GzEKAyahnFm2IWm0leCOnxAE4HzQ6pJ+Wngv9MwlRBD0eE9c4fF5A6w4eBzxF6S
pcWhZ2dIBGcw5npXK4k5kXFIUJEEjo89voRrKBmV1a0OLjubxRFSs1/grxt1c6XN
ywXCC5jwBDjzucBHjLfPFFg49GT/n02g1TUisSg0LReTr0uWqJACYuRpGDzZGRGG
u5gue4tKJWWyAlhAAWq73jJrbKbBcHM1TxH/CdpOxJgvZHWSS+UwqIZ5ntJWypne
F6sXpWsl1IbmhW9m3O5HsUGr36PEqYestgNS21upSMsYJKJFlEI1SQFspiIQ8ZvX
2Vo7IumG9sg4e2/aGqhjMvRpiGoCqYtb76WDtlz8v0X3LsJBUc/IOtyouFiMOMgO
gVq/TxNrrq8l45Utz8rvKUbKEZnHhql0OutLwDe+2IgwweFsW36MNoNat5RJC9RW
Pcnjd1wldey9DHK88WPW4PIxvYFB+2ngc2hyMSjXTex7+K0oSnRDmQ7sboiBdTGp
jtGT75a85eaBXNHXDiOKju4TRFy95G89djFvhAqfL3LbydzPGmM6BPPfqPKIxrLG
JUZB7vfjejHM/25gKar/7WuYq1i4lv5ygStNdjZ8e4O7fMeHpg+8ZJKyaG13w0yt
Y3JZQDbVlvSddnC9dPP40pI44wXml6p028KyK/sRG8USdt/moQN7D5YrQm08C/wG
9fHXZpBd9nPIUradCD3IDAQ+0dr+UxmkbLk+NzxpPODl0MAv5SjOMGnUh9KEQXO1
p02lN+to/KGfgLjR48/CbX/ajBc20iC41S2TbUe8Jwe+FnOc6dH9O8N0zhAa1QPh
MJS6lytsHb/Eaicatf8pyWS/lWZab/FYEXM71CxtPDp8cf1MGJhf99E9LN9LY6t6
uFGSLqZ8J4g+oK6WmB7fAbGRQRfMsTcaYfskoNx8tfQOdWH2f6yJhRidSAlwvTrc
onpOI8jqnwi4MrKeOzFBkigzkZvYSwfhzseBkaeWVuSYsa4FdoZ4OfWv9S9/wVgS
pcobFsV94sGvGHCSd9E6Je6T1U3WbTnycpZtyvOx5rdBfdLtbomBxxDb8rhK+yIH
W0dOnFoefFKHZ+5iKimYv9U9I+RwVKtwBxK1HdhyWw9AdBMH4Dt36F+q7p3mx3k3
BIsAFpCrVQV31K/OhbXj9/TASlEdtsN1ShvQYUHJQO5hvXGQP8CpQ8yIEuyyq7Pg
5/HfanTT7QFQq9Y9rg8nBGy8SdurjTk7v9wVqGMfjHhTsx4/Ul9by1pUtvBGerTW
H5w50viAgJAiFZzplq5G0U0+N8qJC7nAWyYrxHPgXSjXBGPGu56xySoYjqHkZV9a
/oGQjI8u6p2pPLH87Fj8NYke6J+FW8qnKWd4//2Fons1KqA0bHbmGbw0j9zZhDFk
sOeMUD7+TT1oyUMznQyac28NiVdwAjBPRqQFswTohTOTwM2fgTJP/Gm2U0KSLzQZ
vguXvojKblkAHOphTDaBcptfecAUHWGtYLHnKTUvWuvfQwkvEI/uP6eYIOIS8GTT
2SYozQxk6PaO97uJu790hQYBNcoqv1P8r6Wf2ARJy9Q6llDLFFD1miCXJ2OOmdnF
9qiwBXQQe/rhNVnnMYqPECL6jY2l0B76tXFlSnsG0Tc4MEOSpoUENc/B1Mt9JXR4
z1Gs0GQTtxVh8gpBJ01cq9WxiCrmyvGBxum9/o91k6Ys1y2pm1qqRVQNLrMS7fAw
Pz4YY1r0mbj/s3CcYtaSt7Y3fGGk1GvHedhPiF9eX+TECikjBUFo79KMv42Y6qWi
FxCmfIFbiaS+4811ZdLE8e/2iE3mp8PqA9p4aTqRlQG90GRAoRyTS08j8gPCNTEX
yszoyGj4/Hw3V0+JuLJ0eyg7Kb3K4KhZi/4eDnZIBUl7Goppct4bXQYe0XCqc8sX
7T/Xi5z0B8IP1Tru3Qzi+Jz4gU2yqTfxjpFdE1yRLZE5B8RU054yOvWbLhM6JBRm
AAi04TERTeWuF9AlGzAEhPMd2bcWi+I62t4dL8p/ggiDeIePDaiys1WU8z7kg5nV
UOwxFgVAgyP1iW9SRttT4BB98MqkcCrDV3B2kGdOkzPpahB4AmIaLeVMvwdfawIl
DmUXaJoQLoWpId5Nlvj6ajkDHtp4tdhay8g75Po/Ek5H194giuMUVls7LKUHnz56
pNEUC+DQlyvf5aPYAX25IKbdEXZK7LACkZ/h/290JtuRHxudPbuA6A65zC3N6Bo/
7jesDgZnbdKIRb0Vir0scM2u7ZRTNSTs8XmgsfO8T1KrUB7bJDmSO90pNdfkbDnc
EGU1WJGHefCSORXTohMcLH1Ng6YyRj9o+xCmTA7sBT0M7+rpe/EpEBTehv5UVtWu
ICvgv/V67KHTejagot5q4QHut9GiUTXHLnuxVZcLiHTlRDt+FX9xnNDOEkupdmL6
UgZ1AD5oDJirC9ma38X5NtA7vY8ogUoPkzI53gFUtRFvUS9I+J644k/Ur83Ao7jy
Ul894YSK3V5CBc/M0hIL6+buRnGGwBfJ8CV7NZe19ZAuywEGGXgeDTvdRqWzTcCY
+R2c4AR1/LflWslPmwNdq0Le37yY/n0dD9Fjw/iD1iSb2FeGYhct/2joCSjbjchs
e1qZKddM66kYYh2rzWU/r2cgEIjT04XcqGarNvaQ4Ne7ZiNAQ/tdXrmx+iI1wJ2i
iTRF8bKReh038YiRuvXSQ0EfDfzgOXW1Lo5fpaHOFJdoFnqba+inWBfK0uoO/RAM
ttY8go5RqdVvcM0dw6CM/qZcCscvvrJMOshg9tDtZa6qWOCFeNY3uvKbRZpliJIG
QfGbAcIHvV9fhr0ud+TTxCp9xwUTWgAvgdns+OvqxAkb1l6tto/lc1fby5mJdt5z
yROL+BY94u6pb7c6bc6Wu6CvUgwnu/mzEd2bqKEiIOdpcPTb3sWI9EHgVEvUTYna
vn+EEZgmEYLWW+2BlKKK4QvVeSmEJbJOURBoHmY8S9FYPQNDvKS6y2EdSHjkwJkF
R7BDCFHJogqx4WlGQHGqi2MkmlB5wMc1Kbg6rFCV/m8znzfu1p7XoKwrvBi91oHw
yhTbYjApRy9BFH7tSWOp+dA4cFeDePYTRLeZSg3MoQhxbKTmVaBTUWmZ8vu6hPZz
tw2gf+l18SGx0j+XhDvkEVxj7gxwDaQ8FezjdbaM0xspk53ZQrwFNj1HbOO4LkTK
KaGZ06UT/G7+EFhkv0lKuqa1dh1Okm2ahskFoLi1e9AMQELTnT1HT6XwbmxnDiyL
cJyTiUihnzkF7vVPWZJFqOx5cxW45sGzr5rkG9dG9zdFCCr38CpH1RFSq+E9UnOz
rFe4StpFUIiqdxK9CtiRAfCF29smjBTPjlCofh3eqmmTEQGLaVoIRNjrHp97jdqd
UiCCZDDNCqLJzdeWF6Ea8hgnEOXREVQLUao/wWlsMk4qC4KBNB5vDOp3mbgN+jh1
x7gfjmKtO374kHQuXyGoReP195R1ywxdlDIG0lT7mTs8PksMPjiKCmmffU9irvl8
RfvactceJYxgSg9CxZgZyj7Lh/Mk1uunnPUbJWJYlbD0YRMCkWC0uI9koX469A2L
wVQh02pz/2FnHIwfgHzLn49Plt7Qzt056MAO+wTmc29JHcI8E8f4Vm0I6zfDjWQ2
JGRg0M0vLgnArq0UUd7ALrY3tIH1kx+g2L2Ok0swnmCKVWwcFCfJ30iFFAzrtByy
mtJgO5Djd9xtzAQaGrHbwCke/S/KM0lWmiV+X0KsE6WzsQJ5hgrMdfMWTjr5DcyR
IGuxSTIPCQSV8bHvl6ig+AsViqzelGZsdCpJz4ZtL7FSGNtwqep1SBShPns0soHO
VojXp3KJV3wwG84ZpaXUDQe4K/fq3KmsBcB/OjvjUJ8hRnK2hMLuA2eKRzpKcB0m
RkoBkr8NU8rNXVc7lK5WuOb86I4r9UwDhE4onzNeLPOmA6r+HU3bbqLOCv2Ym6UG
xJZH58MsZx8Jh6WoH4RSDKy15gY9NybVj4dvSfYcCDSEfj+z/GwczqW99MRZfJpg
uSAGot22bQkK2rmgavvwWGk0IpAUji5vtv2DRyrNLkIXHdlPNiD3ieuGJ4d2p9NO
8CpRVuwcz/+yyanuDoaZdLbY0JuJFx7MH231Nc9+RggV9tPekT4PkLn5OdLK5MJE
tyGAa4jzRqjHMqQVzA2xjffLTvy6SRMDkfYjYsUWJprC0elNmcr0ND1e+cmSgz5o
+bpxopcflydqfjml0QWu71+kNJMisIe4iGLiYPVhLPb8A99eg2YXFqsh1uan8rix
7JjH8zivigt8X8+buZosWdY5CbpCkqBTBwV6BfetUturMImzl95lHgh/dh8d/+9i
ldsw+jTGIpXHtBZNYOiLkhGCbnZBFHaXFbqwmzOBaYPt+v0OWP/ciXyNYE5AeXrZ
JYWPBS6QhjlJ7kF8oW3d+7cyLW8Vv1ZWCpVFBeMY6MOJ2wDosPXxozIFcWkWgjJa
1oVqa/BBRHZaMT8xWiV0Zwbc8OP7dAPgBdzny+Bz69xD7hUQ8i5LB9oALIvQcGXq
8CwFTF3VB03JVwYRZHAj6YEdhMxdZsp0z82Y0qdI3jAHpCgotfdTClqMTLuIjN8L
P/s6o66FnInV8I5mJbORhrzZhMmONVYDMPPYUAsFNfq5+HT0a/4KufkP8xskE+G8
RsX0dCBvT+P+cWkI9VdKUj/5ZITxAZlKY9Daarldiw+IKSaEvJ8gPSRTMZfSNY0z
v1cqUNaUUAuhbS+fHDLo/ZDT6+X3Dz5tw6RmWqijmK/Isjq0DZl/ciz5WFYYkfgL
yz2G1kCmz5EABqBbSY5v7CraL7Wl1t5gs3iLFNvyg866+3Q0oT2PTD0Go3xcGOER
UIib0Hzz/fhYKLnyEFEjbPh0npPeBDTLOxPq7So35Qgnj10IKd5HaiFl/kxjif7O
CTiGebnRfvdPwVqw2F7Bf+V/yN9QL3IAkXvdejtydOiSb16Wn06wYvR1VYwgefM4
rhcIH7PEjNJPahCS+X/8Q/SgFyBkZfNcZZtWDmaUIFGKM78g11ycZde3EbWgrpk4
S0yloE/i02Q8qboJU1GPPrSw9k7aioDX2v4HDv1JXU4CY4swVPlDnkfYB7sU1v8T
HmAEzfrEIBCp44KhKkU5XFvertoUH3QGx6p7nTu5tTXOVqPqmpxhDFb83yL5Db7Z
80iOv5JNA6NTRttsSOqtts2NGlqhMkajmFldOHdjO0JD3zoJ1lcUx2BaYpe9bRJ0
FfTPCqDAsq+arNLW8Hyrgn/FPTzNkvJovCne1ui5KBjLVW+IahbUuj78WftV5GV/
/xbPTcKIBEt0OoZhd1+vfONFPOys0oTtwjxXqZdf5+jlg8YVQZaWqnOSrZ8/ZtzK
KdtvoSrlFWpaVA/m7rS1Ht7fYXQ6ZCafQyHjPuBp2CxKsuzreBWO1YqUKmcverFQ
nk1yiZxKLLFpWPIdjaEdOQZW1e7/rHKe4lTOg8/dwasfiAWx3LU+Otc27HoYiZl0
Ltic2FHRFqlO0+Y2O+aCyh4OhNalGZiDXGn72eRCEsDGBdtZgXwBkEcDTj+pO1Qx
N0YKnashWEJRjIum17a3jQ8+RzFTisQKjNfx/+WOK+juhX9IGh9xTjtZ/eIsy4AS
R6nq/YEYFQUkpAjdeGl7aN4/bQuxOzt3j4UqeMmr1DX9mXnXO9auJk0sWWP5EDXd
82evKjQNhzkEROwptuWu5CKgOGOU9Zc/sDEeUasv3VJ93eA6DqvylC3TLLHnfIiI
sT+zLiPkmjgH/T/9u5bcvVNbF9BG6SgtDdCUyk5kI/gD2xbzmY2zE3u2zWYUbwCJ
9PXwrUFU1VhE0DIrYzK12xg1D2EetnmU8Hp4Mo61xSeeYPdZV9pDyoRo7MTLP2Hq
F4VupeKyNWBJnOIshCaJfGxXpXsrqcS41zCAnUxW8sToYpDLDauH1Zuztj4pBmO/
2ZDDMkA22cVChp7h9yY6j1RS7+vx7kAEfFfSiZv/lwE23j+wHVRTetlcOW1WjMNL
0v3c77+P/VHAMSJjGHQSZp5bkWiZACZkB4q4WAV8El+a61nSbL9BzU5jJdg59Aiv
WaC8zRQu8JQNosl+Trd7CAYGdMRnlk2QYgGOkFzTIskxgfVrKBjJ/znBfpyVGhmJ
A/mJG8jJ/uOmOhk6EmEWLzuUokH3nMYDsfqL8SX/WUAPHhxmoKKlPNDDf7/jZ8Cy
bPgXTv+gBzC68GlLDzNmzARYbpZgi1pD7aDwj4YBGBy3t8hWV/fVEwezbjr0kmZJ
M7XgfS5Ijit5NnSNqrzCE74WB5nc4pGTD2ZxhfQKL8pwKRf62vFOqggdsxO+4Zl3
rCf9bosjQycNo+/VvNQbYbm59h5JldEyR3ekUyTDHJ7gIRMY8rBDlAkvWnfPKfUC
ariq0/iWh/wS+tQLFDuOMJSY99Ncx2G/BYvv35LCrHJV+MolP5ZE+XopqstSGZhh
pA++M6D2M1e/tzkyq6uuOdASXvWoI5T8YhjH5V2WHgo8np7c/RQ3Q3TvHax5W+JU
UDeRjYt7cCMXkOskL4moEONr3oZZ+oicVPOg9/7tthWaOf43axUTg3pjuWUkdNE8
gB7fVnCwxir4W7p45TFs3WTR9WTVLL98JQf2oH7qP6FM8/5kScmVYr7wAtjcqC/t
o8ub+yRr8pE4P56Qlrn0L8pD7VyuhvOvDF09VDoowOvocBMA3gdjE27wcsBJUjV6
HS6upcBn03Z3jkCPZLzLM1FOr1xqx7EBr7iZzUrT4VlBK2VOg4X6vf1ejPiggA7E
3MWtEdBDgcKmiQcpx4ln98gTLl+mAtQCcogZKfkOmzv2ZJn2psZF076OFx53j4W3
9bpewGPbvx0ICPOTROTK1lVRVvSkUFxSdVKJRF7/qWop33lYVHcl6xtt/CvECbNT
5Vwa1s1DDwxOw5tpg3JPJ/sd/hdV979yRdfyRvqMj5SHboUk5Q/TguA+unHxVhYL
VK35IAiHgnEHJpoId90baPAI0K7DY7NkfxfJtlDbXbL3IzJ/7VG+Ot0xGSZX92Gz
WR8SnWlOmwlLG7ZtK5zzCq0pMN3f9sXDI8accnoVckZA3dwK9oAMmBa0dnaHLkhV
ecJBL5LUvUlRcy2j16pnnuqheC0Y/LM9C45xwDmNkNQTT4WFL6F0xhLW1EED8GTH
Lk2NHoqAmDAUf1/2MOqoAnIq7Ea23aFD52kV71aEC4R70KbsJ3Mkt0vUPwocBTOa
PSYBrIp31NFhc8ED/1L7w46WXKZsqLcqpaAdyxAPxLKcH8C0Fw7TJHTJvSSsKhgR
WJ98sEJ53Da62gJ1gOq0QKZV8mI+PhXjSR4C30V9LzQ5a8cssGkcMZVzRpAQ7M3n
SjsgoqgxGXwpXkkk5X2hQns0EQdD0a6V+xtX3Trwh0FxhxZnMRkXLw5XsEvY+BCh
HW9f1f2GOJvoEOMkznUq6xS/CN18iIS9fYH+GHOXZx8g7uR0cu7NcxDdFF1K+r7x
mL/v3LY3FlosLGNkXilqfS+0UZDe3eJcD9GbQWHluyEE42u8kG2KwOO+3hoZAqvX
WxveG0fg61XVq00SyLhYtw/b6yXWjIlz7fE3Ohjc7rCHqHUGF6NfEmC2ToUA+RM1
ITDhaxHbZmSLgAqRKF7H3ZuOt9DO9RENdXrObVsKv3PiosrZkAR1iLiZjcubqYVT
M1Wf6dByw3+GF2VNLU+wgJHRcZudrzXUYkHbqXnVymJ8CJ3HSrZpXfcNDOHkpHF3
S9RWElexnRXj3dWomdZnuB+Y4N++SD0SmH7LpJrAt1VyEidCYTsOoSfxht2aacZw
HghN+9hWn9wrC6o8obpiOqjfhtSXJDrHAZdbZs+NAYWpcBl3ALAgLYL0EkLPyu7P
UxUHCp+gH9ncmkALZgl44k5m1ZIiTFSwy2kbtIsAAV9QceyNyL+NmvmjvX078Lp7
hVhbufiqQQSWI1g/l5Qk7RgIxBw8uIVoYv/owc8q0XAZuyxZcgdc3602bvHnuI7v
rJBhAtFcLKU8jIWJezSU6yHZPS4X3XJhWDPj9PadbwMtQFjmIzGZhfhV31e/jLCP
YIpRM3gEqxTkXr9VinTXx9ll4ACJIIb7jOu24h/8A6uKx+HMEaOuY8wzIArPeenD
Nm3Qu+Jx8SHoOvpsd6Ff6pCf3/ba79/q9u1xxe6AtkwsN91ET1AIFOpGujRuA4RX
i0uVmLDgFZsrsBBKIE0H7tgH9S4DNsCmiz8FKTmnGaFQMTci0odtOe6jGAJvjlZN
B9AaWDjzARmucdgsUQ3KIqGcLGMcXSwE7JLF/txfKGFWTkwocP3jJD7/UV9dpumz
T6EKQbq7QykDPccg/dJjVDiI4HRC9+H25P5W5no1BZ9G+K4aau4OTVF0t/DTm/r0
Vd5Cu+wEq2hFQacOl6lhIslhzgGoXs/kVlEDdGMhe+SAkggyjRl7Ej9QEcAO31rz
qbcU4EtVAb0fybzmEUDkQuaL5JP1AW7QCn4yWSGv0mELUSU34YdLZRHVX8jXjjxn
V6axKyj1csKj6iX2VxR+x3YEiO9fo2YQa47BAPLE/K7ZSOnVXyKHS7rIpKmk1EgK
njLi1K+vCeZ8w7Ccy5RL21kjN2yJ+tV/Fv75gzyXuTfbSVEOnBJXzK/tzmW8wjie
wKbJd0y8jUnHNgxhcFJVAhkgkW5VQXgWW2Na3zEkFSr2yNJntBls3msVouyc4kxy
VO7T2B4BoYy5xs13XPXUG8SJs5J6rNmUOHAx+5va5OQ+0d9Hu85HnxXgEqFhyp5X
4njgoKss5oukQfrnSvpx9H6lSS/uKMSlhLXrYcweItJ4l4rIvpUac31wRc5iKumM
18Dl8Lnsv/ajE4HcgUsmyyh1Af07n2cV0xAUdelNvzTPsGtJ0kqFYtinBRfdxECg
9XivtPspPlquREsUvcUH4An0y4yA5oIF9G+/rKdWbsQo08Sujr9mK7ancxju2GwI
dzu83AymN8Fj0AZFuQZRqjT7g4Ndq8ISBbbB0WfTx/i4SuvzAgZ6SboXPifCqAZm
PaeqkHm2Z87pMOacVgarbgg1jln6R2ylCm/YkSphzl0GyiOW5e/OWYDzbZyEMSRl
p9zQFdK8xJyviTv/wczJksZrGsXUElm0CBaSnKk0KLxHtPbS1VCD2PxHLZz0XB7h
yP/lnVqoAoSe27bFV/IppkivmRUPsv1wQow3Yjv6TgNyGhmpGSkmXydN7nEfqtTm
qI2Fe0BtAoeIP9m/jS+2rhwkvS3Y65oZXtgontltU5lUVjn5Vsmf7et8ujJIXU9i
ET/cxWvfDM+J85qVy5+5efSKl2hZKOcfL5KN7bo5tOMX+LTsznRfDZJR2lFzLmLO
OxQLQkqPaLQKdyTDnEkQnrk1EZflrATXH3n0YX44sIi9rL//oGeAGK4dIuVs2yWK
JaGM/Cwfv9eRims8sqzx5A5QCLCdMweVLesFPUemhQpMf3FH6GCSRl0z9BCGa+hG
i05G82hwWhDrnh+NSmhUWxee/7WhWFHuapc0X4Ki1RpHjsN6FJQYvtAhXsGH6YmH
Axs1skSkFReJzgzT6T/jAb+MTlj6bQrZD0ZuUBZVL5XNEQsOccdjuS3dIXl9qg9e
nMAakuMKFYtpSIUEaEwcaKn8SOKWbUWaEaCdm2JWWPg7NqEg13OylSghD56Oj9Hr
Ib35xrweC7xu1Cka/ze4c2HNY+kX69QS834XM0eYZ4VoqFxPRhsy7gqr5Lx2f22g
q30psYFnfKbTxa/tBxyNs29a1D7PVleBrrLaW5E1HSi1nwmfI9a2haSHt0TrmnRJ
uXZPbaYBJtkF1tSg5BLe9WErUTf1EjZVKhq+zn7MQnuEwXbHeYX1vH7wAhXkKBAD
8qEAEZDYmmFU1DdTS0e7+V0eDdkx/HRJJSEKRdKpOQvTgJgboelcT+n87BsZa4lS
er3njpcnaDNgOssxxrx/NrqhvWP/5nk17i6zi8VheI+bko/qA87abqM3zu1zPpOL
u5A5n5yiPtd7FoKsX0isxwr4Pm3YIyz6oj+eaGLfsiPcmcOw5PugZoQl8r49f7FJ
W0PZW6Xw7rCA06W+ku49bVWjISRllNZaBMMYpv4NwrNiX6YDpaiovFbT0cwQKspR
OFkxYYJbFEp8uEksTV8HmuzfCegOT4b135QeGrLtb/ffj1S0US7ozYMGgkXb2ebJ
QesXVLWozkURyJoOBpr6rf0UlZtPN6kf1VieWoPAKLFAVkDhRsoKxPCjdbRd+HIO
TABMcUI4HBIr12BeqHY5coULkT4xxpATRcCkbX873YD/Re+08BWoaV2AlSbCbO2Z
5TtfYiZDuvNbUCODhnLsNapF4j6rPXPuS8wpdUZsnKgVM5Mr/TeQNQrH4T/T/I+u
Kd5WnrvVJ7dSNzujicjO+HXmsW/+vj3OMZixy2L0iGwwuLG8mtoal7GFCKIdD7cI
DbTlCLEwsDUNtQfALw5ZHfxdpKLbKFOeCPj8JkR9NCJmtVVW90pvs2sqpfXuZwBo
oR6qkzZi5B0M3A9f6kfZrNJXPyZfP1/gMDUp1jJwuXn4Wxtu+jAD38QVyHgkWU9X
kEzYMt1UyCL3FuhGiu360DoN/43fnvg2d84Ex7XGu3E/5FQp9c36U7BcsK7AmUdz
canG+wwuHHJy043x3lUrpyICN9xa7a9m2od0Yttqnrq9wE5uxdpCYm6LChwnsHDR
WDv2weFtzUFXxmrKEd9Pa9Qk9TCv9o5tcjGKo59+haHi/6HzxWg5RGP4+gHM9tI2
zuvwIeJXxf8CZnABw/oyOhQSGQ9tGlvLCTfssUg2Rdu6lzHks7B2kGzfQGmtsTHt
3nhe3ou+2rgs9TxvNNEv8liCDCWX8yFZopZBtaffkvhck1NBFee0YDk6CPUPunMN
fsKWu6/UwBL91AnClSccWL04ymAGGvNT16Llc2unyO7jh9a+lOxedl5JdNmmxr01
z0dhjaHCzKq+V1mg3/WzJOVLuYZUDi3LFCoIGcYTm4y2odf+StQylnXMwk8Wq/g2
aDEzW6ZAkNvi2/Oyc5mn6m9sRyAWC697DC/nKsJl6sJfugsGo8ocNgJF8AI6EtEw
PErNgK/4jvdlWKD7fJLgBFECfCAu3XOLIMXPkT2nB2eIl8vS0AeSL9Ek7+sqNdw2
RkRIb4/UPQ0bcOd1WdhaT2r+tEaMnQsDRejs++Wxcsii7CuMmV86Hrf+MSvNTJHk
n241rolFdAWTIOz/MOZWGMPbieKdrr/4bPoxPs4wEsGLB6VMj/CXbnjc0bjwAuBy
3zie5grFTF/+j2Baguj0Mp+QCYvqXAZPLhXeTzFebVEBXhsUtKlDn9GQzxIkjJcZ
0TbzD3BNUo/FXzT7vI1M7tylMyyVZqBB8BND88PleQbxqP+PVhCgYZc2letdgbVM
XtBp3JY8GsyTxzc8DAVFW9AJGqeXe4cjryMeHlqSLifwvW/PYoMhx39yqF+aYN7X
0aTrbNpVBPCpqqQhMHf61tYkbgUHzeP2JGm09JIOeAx9nxXC85Egpc1unZ7oEbtQ
48Y8aSAgfvX6sRKjAzn2qTLE4E2fajIg4MSuBY/HtWKiJzT0RS2nNZYn/WbCNERq
aBWeBGTVVCZmdHCtSX2CVcUcXrGZbBTUFp38fQJMRuFQIvv8fszN9w9QIwZpNyHr
RMJr4KUQk/wiWhRJAn23LQrWbNEQmf1L3gpBp1X7lC9VkSAnMdLBW6FhyeGIerd8
xZSptYckAtzSpnSRJTktGgk4Qm51v4ul9bc7Hl60n+NvNXz6UZgmrfUvBJX2Jr2+
tKmMjOFzKuFNcpvZo1QRDXv2JlTKnF6ES16Mbn2WOMDIsUrgktzHgAfHKAMk0kvR
dGc0LVjeG6zYR3TK/kOBWn5hUCNSyFOmm6NmA83stnfFZ0H+YkffNFuyDPQGPmH+
yJPIqWBGKHi5bkkpJbKli4J74smEDRzykPtCNRERvGw/hTM3w74xYDnUmLgZbtF0
ZcgtMBrlPIwDxALlPnBO3hdfqpCmwk+nuIMxG8PCcKN2rq8vzo6NfYJGagi+KLm2
ttp95HppO7is3/806lPRy/9fdDp0Qcfct8/suPYBInGoHMU/audtaa1hgqdZYip1
sGBBjRR/X+Uv9zqe6GRwtJitpl1HuLkMh1uKajJmS7gCEFjdX90YJwcXwH5L2+PD
hHjSwRi5zE8QFW1ICVnM+AJkIHpFEVJ3IyJWWVSnFl4RYw7XrgQdMwq4Y/lVC7Wr
XBaiFgwJQ7CNgBvR5aid8uw+hGUUE0Na8M6fkfh/S84IXhrrVIQCNaArD+5R1vgt
Jdx3bqg+KAoVccSpir343hv4u7F0N4sO6G02e0TctUDVvXJbjzNNDyZDvdT8FRri
tMHDpqPxA6LswncMHclxuizWXT0/uEX4U+VD3XQypnwl4JSSVRiwRYW03K0KQzj8
cl6j5Lr4QC+lt1ANrhaQTCbikiwxvOmbS2yfr8bQpbkDwkRQ3xkx1rxU/HLGd1XI
rRihsZOLjUe/+kti4oN0hf0yBqiWQGGXyf1lS1PGmW+UkzrhFctpT/RMvo0bGcLF
r4krN/qr/jivkXo6r+u7Attxiw6PX2Rzigrg5D5GMLkoMGd8otFlD1LuyDZGuwtL
9gowS2UfmrRXtUyWBb9oBWLkXKvZQvQTPyvqvn9lYiVxD8LMD2Z+pNa/Kv+D7J9s
F0Ubi59fiAymhPsZyeODTURYMCPXmfbbntkBGlERuKXBUuMvsQBTM5/Pa2K1LXfM
R5qzYs4JNim/wV4tQq33qNEAKm8VrRK2LW0k25aXLMxzQVep81mo6//0cGbV3oA/
MNaeb94eTCKtmjEE9eyF5C1Ly7yFVc8SQ+LBuuDRq3RtVqhFcVLdauhQlruxOy2I
NznuYChS14bwmm4qJ1WV0bBonJZAUTUNTMDkfmVTO3du/v+wJIx5b9c3Ujz7Gwj4
UcOWRQcec5ZGNPiDd2GQtrhF5DdO4m0MUkiS3EUGYwcixzdXTxPUBKU6QRGL+4BJ
Nc4goSLWwduVaxsKl47Y9ayXb1EOhYzmj45jmfbQpKwrIPON6tiSvhikVg22LBDk
FD3Je5WPC1rgMHCriOYdOhf+6KmwHV5WYWPA5c0T6bW45kX288dArJLIZR7DRdqS
ry+mDUX6NKKv2DEngDHZznonGYi9LOwfZK4byraL/AWbJHeM31a4TGsxAZiWIr4i
RK2hX0q/nj1MgT2lqqhhdfLDhhoecVLdQ7jHsgpLbG/UB63ge2qatAoJocStR2Pq
wwwfV7m5lP9hiQF33pl2T5f9Nwe6VhSSwi9uLAFcxRAy+XdA/vvZihxAGV7DqfuT
iagKBVZP6+h2+unDzGqn5rppJMUu6akivKlK30DwILO9uEpJ0qeCJWE7zodbX6n5
nkrV3W0VCYOSnnDMN6SrHVbF3JPu5aUZTp3wkPZgCnL2qqLgTVVov/dzA0TcpvcL
wjDzhwtaztdJC9XpQoxP8PrKPGlQwsCso5dYe2J19SSogEtm2a3CXWQ03U6wrjov
BBo3w7j4Uyu60ZhqhVhvd6IpNijHgN7Y5clQct26/nE8Gl3zNaOmGercZAfVzSDM
Oi4T5/AHcAEPN901n9oJ7Gbq136YLBC4Fu0J/h65H4qLPL9FUDqZ3Ml/V2B//32T
R2QFlanoE5Ui4pshn/A+M3WzH/b3WRqYJMD5C3S2pUao+sdgKvS9k2hmbwNpbUUP
dl25hosEheuK1IPD/WPuc1jkWnXy/6zaJr09ipcBxy8E4ruJjJUpx4VzA4oMDZ+r
0sP67HGFKcZyauNq5UxIsXCllzd6gkDAHeGXfmoJJ+pdvPs8L5JKW0gbbWaanC3j
we/BujWpoClBVLf4je59ysRq3uKrH4PeC+it2RERUda2POlG2nxQFWVuo9mBDITO
VCS6fcydwm7pWuqBO9NKYACShYShROTvVHiwkEyMvk9TWUStgK1MUcV0q3KLbAui
aaS7s5Fr8sJpCjfKKxBsPXZdgS2k3NkQTeSE7g2Js6SgOfU7jH9k74KSIGcYx1Fp
bFjjFjmvXrBUdF3xf8EkmjwpXL43LJr9rQupkkH/ORKVrH8UY/Fiv37r8qMxBnLB
A1DfGzr9IoJZ+OrVQsz2jlYeudJs5KvQWhbX3pB7XPSFWlOyEBN4cogEcskRUNx1
nCIvC2hQ8Z+D1KNZ6HCpcp1JIOMGzU+AeQW7+LeOfLSj3+pj4D5wvSigIbwdezto
R61JhHdhtgCDy46Gg/9UIyE2ef2/cX7bIpoxZUERRvH1/tsCVksixNETLxt3KqUE
OzX4Tyqv6wkTowCkAU7JT1a93vaL29nKm65kzPdEy8/4h/f9Go4VZHRghhoj25s9
w8s1ULfDMus8XM4T+oELTbXpLR5JU8tILEhwH3TDPSA2GNiBSa8E6s9y7ytXgfI8
mxx7XNyK/9CFQTTsstcRv6LQprtw1jCJtjyOdFfpC2FWbdbx3C9PAmAOss0Pp+B/
k4qP5KPCEE3ApKDu7xTHGlC3H2fHDQrQc6DUZqyxzsD+0sjKDxnd9k6AU8L+NRGH
odWJYY0xlQo0UmphMKFD6AUPXhS0cllrC+3Ep7WZRkUE2pzrBns/Dhff/78KYnJo
9UH78RlXz+1y2l9vXZlQz8KuJt5b5IhR7hSRC/wFoy6nbS81mbN2/CrpQzsIYTSQ
e/Jxyzq9vAtOJcjgbfvS6uJRFDGgWv7R+c4OwUmsS6BTsX6/XwEyak+UcvZnVxMo
RnHwLnOco+GxnLVBQTno4dUWncgfp0hnAK0DRmwDbTDDU9f/J6BkisVbOdzeqQFB
LDKIfx8WOHvjvaByTmTyFhL+Dez2DY+vG9yOg68i3iuFXr9xMOS0Ny58ZRieX9l8
xdDchAIpW2Pc1NSR7pD81Ci7wQUbNdy6JrezP0aq6aNsaicv3BF8cF/W77KmIt2x
O5M7/Rfz52fYg0flhzFac6YIfiJn1Q8kj75x0jMzSQWmgyAfx/D5niQ657nnrPuC
W8FGTUOp/tvxFanCP8QSH88LeyNp3DEcNE7TT3Ol6gRbqqfJ1wAUfV5rt/5cEjI3
TsXnHn9z9oyEVrCPlAPvW0z/9YSBH3lhyt974OAnRF4SFz8O5JGY5FvQ47vBqvJn
zY9pyqJh+u56r2juHeW6ZP9HgeGit8AAR+kYti87gDIbdLyAUmMi19MRy0fOWBi9
U0OzIOVSmHu0PHrT+BoDI6pjAIfKKgD4GhlTxGcGvvB9f0C4UW88Qn/v1IKeSLm8
t4OCAz5/vwBTlxfpcnAE5sMGErCUwxWwVQdz4EP4uInAQ8nDwwnZ+i++1wWZibDQ
N/I0Z+DwrU+GGH7w84brrehILG0m6Q/UC1gW+QDddCi/MVYThN266nqkD4Sv3LTA
L4wo3ZuFSRGhARvpbsud+vAvFzzmiBcjI6cnDBj+5GDqGnP2VZkM0GEClRGwg97O
M/MJFFdL9MuWrQPfxwIdL7cX5yVysWTqsMYlGmH4sLrY/OHuAKiGAwZy0VeC440m
lDRdVK5sFiBWDgFEhqF4rP1A9WgvUXVS+XQk7eRFW6Nq0d9KGBdYlglsOidn1+C+
PBEc89GnwCQ46SLsjhm4KJdyrGaof7DChAR5GnzzO8PytN47LGJXyrvRI2MRNgmr
Tugv6BdxICoO/jPICUjcvxe7NOskYxq9vxIQRawekgHBbwprt9X85sEikaJ/4NvT
w2wMgEBoi0XyLfOx0jpLSL5N6dWzYpHiFsan4Q3wX2RD6i8kejOXppIvvbmeDngG
n1t54QRP9/9aRiQemj5zOrLp5qDQPZqnPw/u68lSaDTCwex5qQoAHHPA4CJHWjkv
V8isZoKQCEZFxBc7+tIsGe+Wh1N38/wXWYiZrXWGfLv7c2sEHds+ZOnvOBhSl52/
U1k4huTQ9mCP/oHX7vO3nAaXky9on6LvVqLWzGofinCtOlStqhh3mafcZOUtWhdZ
ZUyQjvWRY76H/F1bTmFTIFfv/t7ObKrASrjcEe2YUOtUqHEPhY2ld11OnrdexhYS
5ZAoUt3zW4bVSbZOPr4mguLT/pcNwvlX0y7beGxFjjsX5jnfMrtizdf8cgeHiaNQ
sAfnvYeQi58XpoDLvmMJCkpZgYnfyQRbCOwPfGYF0Vt2qPmIq/G7GNBMO0Yb66NV
VtjY+ngIlEbVWoshojLZAWWCi3+VqGlhu0l7C1loOGSUu6MHPDAeJ0aoYtPIBSu8
HXHLViHMUffZK36C9eVS1J+uSxiFlx+9wo2ASi2hbymTnmLuq5psnYmR+TYiOHsc
+ztkO7CGb9GGwjPIB2q84lkXc/PWViWOVyIY8jdYK5BSARXhjfxus7+zNiiCTy7K
Y2zR2xx3BkluikeRdSTO6rMXgDNUOi1U/WFS5c5qvM3v0amxn2Nb3A5P9qDl+at3
sapzpehk4SsI7LfJZRodjKW3Oc0eWHmsCLZF0iws/ph31fifE/MAaqjAnEzoNcEw
ppfBJ2kh5/xD1urpPznEJ6buB0kJipLOqBpyFTAEDIdApwss0w+JKbiFZfteisNW
7exIGMSn6+oxsx8QlyT1gUTzdg6BtWrOB+z7Bxt1qobAjcAmIKzqX2b0w4Ldvfq7
5YbXRIfr5Rc9QaBKZOW2FmZGVrKMYF1NXJQlz423GBXSWJuAbh13pyW728ZrtuZO
9Npq1ZfOLBRVjg4cZa6tdfopgM1jPti8UY3+D2H7CopPbCm/8WZgYzpMBrNeoImT
pRnVCKOT+6yubGdbQc77w93eZ6M4/99xqd8riyFR5jV5PkxlUM+ssC63q2BCFuAK
ieefaI1C5Krb6Ww/V6tieioLAxDj63xjl4XcgTLSEDu5IDsVQIOMRwY56Bt0Vq0v
3JWZy83xcr7yylVgbjYxgcAozcPfwzU9gyUueYYzFBYfizVDMuRBLFrWwW6zvf4w
Ej13dXaDi8f1x1yfPBEyW1SnPSL2dSMHoN2BTbe8dkk5cb7upzCXfXqKp2d0Eaem
uk3yU1HvwHf0qXP1tVVU4CxNQ7kvHUUAoTZ3k1lXYiA/tISz82taQEkaVQB2lO6J
lUNWMJLdcgsB9Q3cDXfXLBC57v5EgMNyeYiYlK2Zj/QpuSAvTMHbzLlirdz+JHLb
LXH41uGq9QE9RfkRdJ/ZX+o1POYMGV4We57VvQum9InBg5NM8RGxXL+cSkhJTEHC
S/Cahd2pzYxTkNFkSrDGAUQB1O89CaQqbpnIUSCF5bz9CGwC1651PLK4UOFIxyBk
db4SvaHRoYHHPQR71jY5rwLuWnWxqswwf01OnbQB9edBqQJfZSaxyBmNMjVysdFc
50irh+i0wbKi+BlJgIaolucmr7duagehKRfyZ+hlmWXcnIY8DtoOrO0jz8+rw7h9
31+avw7O9eqUWJWzytTlslUXxm0pfU3VxQI6PzeC/fpW22mpubx36JeDeOrhJF3K
MCstJ08Ksn3b4kdcmnQNzUTbszoZpdw6l/ksAlqhK0LzZYk2PKB/U6v/93LA4y4r
g8zKFYMVzbDe9HdW9ohCE73VjtZMsiUuPcaVOVW9qQiu+eFKNfe6H0djrNNVZAZG
NNwzVRyl4KcmtmmyLU18AXykPBg+go6ixvcw1G32McFJWaAcH8O2jEbok1Yf/Vpw
nwyX8VSKARcZupRdtmYCcEL27PC/H78JpMPmevvcev62ycCj2BdL/8AuyDPqtG3H
9+FLYGV0lgcRlpszj3T3km9dJeNP7PUWyVTe/ulZZ75Vsl8d2lA73FZZyJW9Qqlm
UM9Zz4RhhRx7gsg5Qlj+duLwkVs8zNshdAxmDdsg78GIpRbLOJkhMP+M2x5lBbmW
CiojzPkFG6VLHnSsfIrbVsEdUDO39Mv2QlBw95FJP0/p87KSDtqgqvnJ6L2ZJ9h4
AfspslZjMzLQWLWq8NtKHolYgY8hPnKiMhsE7rMu4rByT9N8/tWGByHGcxkyc9Lm
1upgQxtRU4qH32MQMo6Id+dbzQC0uwz5tB0gkEP3pb0Fuv+2sH0XFaH537WmMSLh
cuRD/pUJr9wQtgkB4Q7ipL5sa+Bnt6SS45H4mUZEzV79+ShLTAHFF13Iq84J7bT8
YDav+XC9xxL/4Uw4wx4S71pWvRviOTaH7qytbryFGtEGSaB5xLwj/jMQBvJZ1A/w
wGgUQACAiFeaM/AYRtfOahs+80Dp+Ia6kHieOrNgB7jq2/+aA9cnozlv3UxpYe9J
Cka5O3eaUAq5HufF8gNdUZ6MNougNbdc2SAFFpjnq0U38eSUU7hsbJyAPn93F2uv
oRIcusIeHdi6LqpxuMPcENIPMlV67na/BB8ZOpWDzz9XQ+4xYsoWIijX1ki0tBW0
3bSLxbTd6Oe9JHjRa16Zvszs6DGJv+QFH8um2jq0V7449OJZuHeAc2NL5s6501jB
e8PazKI3K3MZlaJyrUYO/N31WMrOeDUdbNfOhbDwWEsxpFwu7ogISIlGC2RhbJ50
2ejy90z2uPrpnK5JYB0+GEKqua5lNajIJykpUBRJ/KuuZ3lbQtc7KVvvM0fsKXAA
6JrB9+id8V7KdSGueTUZ8c7Ezv/QWUnt0pm/FvqYK+sYX9Jz+Kqo8HBLBYTDnKeA
KYVLq/H3zg8DBGjQ9OQKFh5TMHTR2UuSU9o/cxN77ru9ZGmwHoS9g3yfNdn0Mqnr
dpi75DB1NsSxEAqo/cFsGInV3s51Wpu/U+T6LHJxAxv1V3DKlNMPWTEMMe5ZSK0O
gkNovFjGBl3O5aN/CiRP55QZf/wRnh+NP1wIi8AxMu8tg4xCY1fVaxRiactXCepK
Z8KnywZuB6QG2NjoZ9PlmFQWY6RCYJVeD13sqPOwkgV/M7GHoZB/UMBf+FfCVkmK
wmR0Jmt3atnFi+o8kVYoX8DgudXROOuQpYpJ4/dXOiE+dNsP9eoc5xdt85M+3lBJ
STcJNjU41rf1XbvYZvYSQ3ot/oKj53UMYRff/mP1M4d0m9X2beTop50zBrHOGFb9
4D3UFZv05sPjmObYjIz+mol5TrzJue0+839W+FS+UQ7UDMQwxoGOQBQrFRG8PzFb
4UHUPWW4KQ6x/41skhlv2Dcjov5o7lFa3328dmlwCrVYr5alW3RpV+rY935DnypZ
sSmsnj9SnwdseYUu937xopfy95PG7Hq1pAWZdCl8g6mc+A57cl1ODulr17+Usk+7
hiblVzMfJL7023ELS7bWZW3RQ7tu5bFw0mKMWvnHsM5ltPM7XRXrW+Yh9gnxpnRJ
tbuhSpblk4O+6jH3GKdfax4UFXA5lA2JpHb2ZY94r1Uqxg4deKdF1LqONBVdeQUN
98Hc7gwytWmSvqeZXRLBGam7vSDCflcEePQrVJKeP5kt7cwzxm53JK2BYZPZcv+q
3XwBXdz5n9a0Geeq1ntmcMrPyS1UxB8sonmHSCc6rGD0V9s19rhyYmCRSQyX7cN7
Fs7U9KCQPjglDMnL5hihbuXxFOxpBZRX/6QGpie9dPnd8MawkYP2eHv+MKi2f6nW
x18wAHWINaSOxNK2EqeVFfLGVk1LgiQvczD4lSHFoWu0CAmjltBwssADP1sPFTwZ
dmTfZqWhUJ+CsnyculYA2jbLp4+K9P8ssVh1vJvzXfmsqM11JSe6GbuNg77ZO69S
eXaYjsA++//EAaF5B0MPJsB+y5HQvjT8XBucw6maFmejg3xfg5GXPeQP3S7mTnpf
98OWutwKJXZebpchayNNAza6KYDPOvr6RLvcqjnZgDrtrRkjXAtly2bavwqFGN2L
FvvFAZKH4pGE6la3kUUM12J6DPWoFaHuC5+ctqEZsqsdQc0D+oKMG4CbcgG8i3t2
cpR/ELKR7xSqXtwoooUGAvZg+wQkffOg/p8asHru99nvVge8sPdS7+Hf7ENTLTZE
A3rn+vOt+5bVsx5AC23R7grib3dG3uo4eeLNFG9gjZSz2NrgD57YY2s5WRGLAuWn
dVgb61dr2gfClImvE3Wi0079HUhFqJ4HRjtb9rrzu+d29YjEpbadEdZxZpzTEHy1
7IkG39zGJrgTvbQo6G5jXd67SbWSNGPrKE00GgSbbjS+FQXzAtPSR0eyFOzi3nGF
pJafyJieX2MZTjT2Odp0Ch6kndUK+K14VNct88BSHpCx0WRfuKwbiDc3u8kplrgC
J5N3pgTyxef0r9X6u559OtHTlBmwljdyVQOVZ6Zgv9FANNekvGN75Bz1kDDjRl6O
SvxBSt1jhr5KiDG6qSAvB+LvAk1sFjo5Wg+6M4dyAWux2b28TQuZHsiW+/jrj2C9
nnU/8Jbn7VQjp20zlveYMpjzR5kwYjemNdWvznHrJshLbuay6VWecPvj7x6D9H4J
QNoiTBs+lBX1M7nv2xnHdVRqT3tBYSewkUixzF+0xCsF23M9tehBKb36+TuINJTP
U0HzO7UjeB/TdAwAthooRFm98hrtMnPYb38omkjsb4JH4nrjqvYCD+6nq5wTOada
+0gA/Ve9dppAw4zGv5mq/dNd/t0yiMzIsIHuQAiPpSY2LAop6yO7JEcTwgt55wwT
iRbODF8QwcZKQvOozgb+XLdG/Vm7O5N15qEr48PnJtzeBvthqwS7QlHZcx21sZsz
QnKlMdJ6u2bGAc08xMaS8Xw4wiZwnATg8Dn+vwKJvIzEPqa96GhXnKwikKm5b7Ez
ML6H2FfuTTZHbWm8kxolIl3dVXsrqdv5f217CE8D+pIhrNEHDQWe0U3FlDYFqlcw
lraOxSQ/KrTXw/mriceabIrRwTOlNfdb9DQxTazdmkBFkWMjSfuW+hH0EXWjo41z
NCYRpxDHLRd37eop1BiZpI7uqvaFnp06t+BCho7v9ZcmQlNY0vn2bVkLu1Q+ycsi
RkqsPy943mFb9IXHMkJUGPBsDZlw1zBkCjPFnAJF9i71oG0nWQQgDaAH/ksk+eqy
QnH9ZEUU7PFpDKHrcizUt0I8mCRi96jpN9oaDulwdqA/X390mVsR7W8QXfD66PGT
lNboZ0dSn+WCWcRvOWBg1X5yyXoZfwieficQI47sM8O2lyIZgEHrVK0JtqeDwEN9
53oVVarzo0XJhnznddh0jHi7GC2Ii4gOhkEYFzbMsQ3qdJhNCiue3hL4ksGsfQvu
e7dJ8N08PJOoV8JD3LGuDaun4nJIfAE2afMgzGXjhhElzQqB4nsJ5Ki0O/2pFqm0
jcL9SzscOm+Cf58stKtEdG3mBSggO/qt7C7YKE+wxG+2Uic+YSXEbdPVzhz9+RzL
eFDOcNDQYj4ftuWWco0IXW6Uxvrb4MPtnX1p5DEvixzTTGedls957G/X+3cbdBGe
kp+qETAocp2hXmWiuM/nhkqnSL8cRQQgUoQS+s0Bcy7ebxysTwXK6zzSqGcGLUmz
9PcM3eXOqik1TMvjuFFdYY59WAOrKmPflKNu+vER9FUvFtp6Kyemsgabx8gePcHX
87cScvR/TYqnR6VUyn66iPqB/andt2GrizHowExd1CsAUgLtJ+LeuqfuadCVVyWQ
iifIsJIZv8Yil2x/QJgkhF9ByVngeZXqdTUc9+jozYw2CIWzqUVcdOMaSwT1qVXn
KdswCo0qk4JsDOpbT2g10qo/DQQjde0RvgevgYCiOb56OhXPVCLeVc23M/v5tZH3
pPfMGHpXNYhWq6LM9ufwYmjQpiE9ldtKJ6597Nbsw8iHvP3WeiPkkVrk8JupqRwF
DRSmNpXIgHPKty8bjC61KB5RWKTn8jafNgRATH/67Q0SWrWJzzt+OKlHJg1brlEc
9bSdgL3RoZbujrAGoA3BojwFWTry/e88nA5iw2wCLEgTv6PE3BFF0lusZzJ+QWkP
mzseJ1PmLOps1nKoGOasfQzdAQ9mhalp1f/FXAXNA9uCEs91XAou4o7RqyXRgHke
eRQdJnajnMAsjuiJXPEUrHWgFOhHeDUsB1ZtYc/RGpqSsQIR2zTzEeJjs6eVMrE8
9ZFaEJ61k33I2nPjM26r0l9fvDBsS8sjaXCS+oReGl+ogJolMdaMXWbk/x3KEL1H
Q2EgE1AdOFUu08eTj9KMs6xDhtdSxqbjY4HwPi/bvFbwpU1lWgRMpVqf9NJM8Lme
GZ4zkpAUI7nQy6Er0tnWHLtp0RTFdo1jU/Hheijulkp96x6Zl6ijdgNzF3lHIWOE
X31+wkiHTnGYebXlZEHjFFp51e4yC0e2OGxENr3XO+kqms3N6PkPSdVXc5FxgUkj
aBgx55+y4lQp7XQvqCi+20f3DVvevHU7qqslgO18U2T8ClQA/3jIUDv//WH7qHNl
3TV9W1ewXfDk8d6EaqEqiXXVJ0wb+WE5dHxeNLtmRNPiMaRRBBm6KEqk7QnmmlR6
zAFGbsW9DOQKDJ5n5QGpmbmdd1ju10yVwfnrz2jYTkB1dYugmyFuiTbeO7l0tsRB
NnuVPJvyL0pxugW86ddLTVfnZstSJEzq34crbzBARsy0RovnjkFExyU5ovhatvN2
p/CHHRF3T7c/bH/rvN8b081FrQsZG8GYUSZoH7zjYNejVROHQORS6HwEG0uMFub6
PaI+cF9Gcf8Ss7EiIF0Q5X9FAZUuoT0b4X1I/+h85asW1T/PPg5i8P81OR1TAN35
QR0Uv+7ErOTjP99l7NIPMHHPLEVR8HN4usFScVrnGmUu0B3a0NLEoUQ/9kiYRLs+
mcPnD4+VlqMOvfQTr0QKFcWMAlSDXvFHV4jLbJaPndV/1ORngiHwVVvj0v2n/tX1
MzOC4HIp0gkxPQublqcU0Pkx/lvEVNY6nnNAbfvHjVb+dxmOo/ApfFPhXUqlkRnj
q1kZ41JCBDAR5pcskGOpm4KSpC+biFBDN5luRHrAc5hKOKjdo0RR+26H8cz184rY
MeeEtpFv2uwWwsBATePyOeiQ/MCeMzBsCwuMo/trzdryXXf5FEPCZt9RVzU5gAJe
NcN4DXAPOBJpY6ckVEccHO40G8vbBnqg9oG+DOTGmw+ebiaEjwdIKbC7wnfPxHVN
IYmCWzdcBcxEHzUMaqd0UegEpnfuyXSV8OA2IZmimnbIhl/bUWZUFymd5XofsExT
/L9eTFx7p8uZ/xqnNJxQYiNSIAXdwYLQnplenJbkp+LixaNa1JldXJtdgwnVFPFp
FHU+gNdIjUcWDq+T7Thn3tpNmDiSG7Vwtg/cuYTuEvwYFTfKGdR+tA2C/6/Pc/Z/
vSfD0DlUuXTvFkRwCdqL/zuKZz7emsZjttTxswaoFdqwXXFrpWUq5IuyZrPIrBtx
kZZWTMDAheKCJsw/DffKW+5PNSG+/JXSO0fiqQNzLvVn5ouVcn8EWDn9VpNo9X9c
9bTunm+nD9noTMtnwUUtuijsCFiJ6R6cAyOUJGhibHVdoHz+dKsEOgs1NH2+tpfC
8mqPhARRZMHlYfzwg9oaG6CIdA5h06m62oTG/NOjMeU1xgU2P/891qWmMSVHMD9K
kUJQLsMDMG1F2791t5DMrMvAZFgLbDT53nbo33EXACQJUhDUndWw7oRH7Q2a8H2Y
gbYOGrMUHrpJm1lXtlunejrINx8ktytJXArvPU9ChzDaF3fLL4fsCK+yUe79qgmh
vvh4p7WtUbaHcnSAR0Gmi+eOq0GNiTpoYKyV9rkWbtf+znpPqCv9fgdiuoe3FwTZ
bCpNqZBg8wkB/3e+0LmMJy/RwqyewpOghggif44M0TF/4SzxVD/bk0r3abm9eSX6
Uwk8EZyVlTt5K1f3EjZzMmVNm9SPj/1Lou1RAvdQ0d9jaK9OYdPM44Pdgl3ik7m5
xvAQyQprmsksa7egzZcfWJMvbAdU9ROMcuNY86znEEnaTkTHnXo+3RsTmyt1eoGC
ZqqcVN/s6DBr7pATCIa14JNYNsc8OLWmBniVQ0024Aqe6NvkghjVetVhrYIG+QLL
IEKvNyrkV8L3/6oR87WqZ5FKjwEt5QX2bB2AxQSod9MtJCx8l+2R3ud5bPu4L0Sh
I6H4asH3rkHBxMQbN8msaJI8K6MMOlkZoE+vv+DJLJDJ1wfhXqqfg5/1KrHntVZV
loEON8BhZz20iNh+XgtjVcYDF4l5XhHNGmGONAXeiZYrvJg6OayEwgbUGcXTnuez
NGugZyenQjilDgEM9FgdFyEal7DWWnxEHa1UzQX3FEIMfs5xewjMsLdmqi3WcVp8
d1+ESJSy72p5tmZ0e69FUcgSvtWneRUa1NBn7iWfcXQrRb9bnMmUpvYaWJCHFRt3
bgbsfcw4FKjOBRHvAl5560fzp7+mWnFcPx88hK5a1ilXcYv9z6xJOhqHgPlsN/Uz
O23OdNvYjjFN01XQuI2S5x5jXCmDWsF4yuNPCzlb2CHG5F3JlFboahtTwD+r4oTw
4naxkleBCbxroOvuzvE+wRDbJtQKquLPQ3Fj0qDfr59Nbc0l0kxbkpwt1HJvQvxB
rG6Y07yvfE7lvtjw911K6g8gJ1upzroGwsaZ9hd0VUDFBVyy954jT6NNZCXvROzK
UbEeN7AXVrS5nREIm0yhkFgpFxiePyUpM8PMXOGgb/vNVYwkh8yiNi4+A+hidDkf
eCBpSGrGmvAWbcGzDznuBtcuZ5ogYfpOvDu1XZmatOR3xmQw+WKEYIrhaCKO+ZUE
X33dBDYCx2jju2+OG0U/IBlh8+x0xiT9ynLRdfhc5bgKges18FXFRokWIBdECWWl
+LAiIPytMNhslSs0xNU+JljayKFlkWipOI4RO5LvdnH9NrrcLgBZEZFL18Jnc16h
oSoYlRnoLCdv6Ko5dHXYGId7dk+8/U7ksyemDnEjnuuVoY92GNZvZUOvmlm5XHMz
T4vvyFiQugNeryBunH0V75gPAWuf4/8ifw6mr7PwJfCjcgLiowoDwLAHJhsvN8KZ
QkdOfLbZR8c9/R783PnLLiGDqSTC3F6pMQJ+Tu2KkqTE8LVHf37/tEJJdarxZ9A8
ZZKKT+qn1pIquSaVkIl0g4iJyouCzI8B0Sl/IGgum4Ub3suTsUc3ZXYWStBln+yv
5m270RdWqpmUwzG6ozQHS6YyJXgzGvB6DPYv3hF58NlC9xPT57wFz+q/3/KmESNe
hodYqeeTR2hscKwj0oNviohhM2QiIIGaRkW5L4dRjKJ5MjHtgVtSv1qcfeunqN3p
i1QawS9y9k5jd0CPQTVxTMxL1aRS0l4Qz4atWhMYkf+Iv7d+hffjcIDamegEhrol
eQE/9p0a26rs3kKBqd1i6e/+hb1R3PJbnJTDE5lHbu9n64UkcD47bH9Y1r38RXnM
2QGPcAqsSvvGGPAvOnVXMvaR/Xpd/1mYD5PPyKPILcboITpG/Tw9sJ6r5F8L1VkB
oxw9koXeQo7dyNf/kHm56TGTs36ORgt02u9R36ns2iunwZR+mTeq+6igikq4xI8f
1LJtsjNYO+I5mt+ye5UznlKnyTTcKamXvd2jAG//Y4u9PUY+SNsrVrZRbTMRU6XG
MyQd2q4JlAT9lDahh4dHigTcj2WpvagxSj+JAD+TjS+lC5+HQeg5iqu1027WHxtU
sY41ghZlbbDsOqEkBhIog63DUHktldt3LyNltpTT+2zrl4X8rZSLkbQzsibw6MNA
SVg89tLVXM4IizPmK7VUOA3EEqSkBKIP9i4MA4did+NkQMIqiGBDQ98M2v8iTqR8
V+qj9k8GgRKLh1pHxJXNnvl3k5lSfp0G6YGQGU+S6CQTeJopfJo6ylfkEOPARjHF
fwikmY510B3GVLGZrFk3K5GnhudeikNTlBViqn81Klco3i7Yl35WMbLlpGK4/e9T
LF/JlP9UsHdak0j+mGEtxuFc3uokhIwDxjZQKvPd/yxV5ixBNvVcLyQMeIdp37fO
Dp0ynXNQkctfpKo23uTid9EU8ykvV8JWsu9ASaawZ/bqAqqe1p/7ESXXof0imM88
kSWX0Hs0uIlT2Hsz51zgwB29x16aVtYerCSejJ3vLULoNfpQSs8cPsZSn4tZg3Ic
anrW4VWIglMonuowJHF7qjbvOiuJv48OxJBRpuJ4WVeY3OVCiA2mFSFDrTakskYY
VQTDMAlHdbidxXQxewrEsEaEResz5ztCb0Uv66AcraXp7BzgQL4YD+qiixMynW42
XITKbOo4DWj9433z+T2bC9JfrvZvJ50jqc94w6E9v1nqxq4R/Ej5Gt85BlvSUx5K
T4cXefVKGTsDqI1GE+oIGsqD7EA6ssG6sZmDDuXph7GcV4/iPd3SM7Jbw6YhA8Ma
0of5yKkcyfQo7imtk9LZMD2+IJeOyaO8J5oX0SOkFabX4LMsDvzxL5QldI4uz2F8
+wyc6eT4N4foT7xX39sIFJY7oS/bSod9T6WY4nFDJwzMNywaFcsi1tFquWI8+9q5
ScQEgLHFxGlnq99eh8aYwqZns/dEXzN718hLaCBy950zYS5AwvApAj9qaC4DqyG6
cIu/rmqYuK8KCn/85ZoY5tIJmqGBQA+dPCZMHDZq3tfeAlM/g4OxkQFhUmth9KqR
fAppjuhWLQ7seLwzQ2i2GCr6wJVG0OGaqzmOkYncmj0KisUFJTy8oUfRMz5DLeIo
XliLfSkTVNUyy0h2dz1JaTbN62yg8xzKDU+Wvz+aOl5ysZ3d9wqdLjnyTnPu3ZBS
F6tplc5cdzOI7zgRnTkPbpSWYQRJIrRROf5hTD5bQd1MlHbhnQeJbHpAkZkVmizl
s/KuvfyTZk7+/C9CIS3OuLJBYbCyW/FgJs4ZYraMuOkcbmn+xHKXUlanhM6W3Rck
CIbckeURSip5/NExASunB6iDHxkaDQ16DQhnTvALL9Ft8PMDcVs2w8EqMGcZ8sI7
B94WN4LyN6IBmAfwPh515KvNAF5Q8t+moLJPWvZV/FdsrjvZTqHZqj4GH/n3phvI
oi1wq+/nOzWRvbORPaOc8K7BtmFNEauyHeiDHuvLJc2mW9aeRRVuccFD8/XGYAzH
Mg//whfMVxTrBZ16ULhGHCybTj7ofe26c+xH6YivrTTBTsERZDD1dMRn29Pqd7dw
1GgGbvTnlejnOg1jvnI1xhvMJOAFPLjh0aeSSQhKgOSHVLWKwZVJ2EQoBWRMDgX1
XFK8sv94EfkL92cf0PA0h5mf2iEu1/bkNfdM4yBDXLJszxLprpESRUClFYKW+Rhp
ww0/3aZ9p1bbSAjQuMhLY1HF/dP8KNgWTSWFlotiqiv0+4ZHv1g2whCLx/OMA10k
bAfYkWULoPPhjHogBqX4Yauu/4Pj0JCCmKIKjiK26A+Co9yyVHW9rYkPQRJSWKBd
kG6iG+Z+/34GWTkI3sAVHOBFAXR4p8vXySslcbP3TrrFRcR6Iar5KWPPm37EXy3F
CuggQMbbaL5htDUGujmB6/Wg6T8+0PiNXYuyh5wiHuVAm6HAB+an7FUsxRRq0B40
DqHi0k42t9WyIdAnouT1dQHrAXv45oIFDBA/LlkC1vobJC3kn3tlsmRwpHpHu55o
xnszGOsdbP1L7bhr9p3+uqK2AI5H6bH2UbAV+pgKtNS22nG7411cvZc/FYEnpRCZ
KNQc/ooaby5XVYt1tO8MU9Vfv6b9QbNVTgFRc4NN6dZXF24eLG28dd81t3vqLjHa
Zza9qjqsS/PXwvZnjsrgOEyToOBXai6Kx0acYwAdygkjeP/uSYfB1X6l3EUvE0J1
kt5WhT26xOBcvLWyNCJ/84nXwHwPLMvq1wtjp8AHnFDwaR7CmtlBRC+ZkRTNvZb4
YpoQAwm6OAXM3dZv2o5KKDGDk2HX35SELFKj/73LTGSayFvXEldDbYsLJS86CMPS
XpCA1aoCXzWJqP7aqqsLQ7w0mGh/I2Dp53ewJfIWaHhffGzCg8Hvp+CD91wemUre
VCKZG3FEX35Ii96SB3rhxEnnRVOc/WQeKG/qSuQ4ykO5dt7kl/EwGY6dLUDUPulS
IloOS5YywWzKI+2eP0uVfByGjXCdGb4JACWR2+h9XBPyYfDi7OF4II+cnZ7E9FKo
IQesrtF6wIPRUE+/CrEzeMC9i7n0UgbNTxdJMfcCVklBJMj/wuzBlWal677TtDXd
CYN9SWZ/bzqcQz3pWscfw17nWEnaCd04y7+g1T5lngGO5Qkzv08qBE+C6p2UrhvT
rbAeGZBHxRJthMaKGhV2y/J2vE8N7mW10g1u9sG8WD2pL4GSX3JEVyTJBQiE3kxJ
A4YbJ6aXY4SpGOU/f8LUq7NSr6vBDUR42YULQ7hsAkSHCZ8dgofN+3V4xnplvtt/
dcoeXsRFF91ZZLHi6SiWRCms4vim+iixVz8aQpTE43hvQy7+kVLRmv1FQP+wrXBm
ME8czBVjt1xf77oCBzZq+F4h5AaOFA0dUhdkSIHHYxye31Tf8QCAja0fZ+7urlTH
i4WfEGktpYNwpWnnv3/tb5Kg+dmuVvalZwTufQPCEGE+8HGuxRpAyeVANLHaiVh8
djqvyntjuykYzowYbeAWo5Cx81/C2CSyL03LlU4CanFVvDvF49ji66RcYNlAqiqC
izB0USCJblunipHeQ9Qeta3SGJ4WIQoDtw+iIZ0GxuOLfgl04FwWBvtlsz/MVduv
QdklKyajAFjPxKKfcN8B1UQEGPT9VukRl51X7meak2A54D3BjalL9R+4behZC7UA
ohrR1z1F57EAiWE2X9Ou+0yitgchtBC2dOiTM8K/78TcGPiRsGA1RdbzvmvGhkML
QbKE3SAOWOptsif8k4FMNmnvpZodIpn5yIEl37ti6KfBfxvcfrDvkJFKUq8AAPo4
rUhzdekiFOKJYcJ8S4AQJl2b6mGwCpCn3Xsr9SDFE/k2NED3jtHxNGitb8QtoPV8
6bQ0xNNTXmwxWvIZhT119gftkpgpZZv3AN9CnbRLfjG+Ya7Dcz89HBrHYZDMWHX9
+EXKox0hLbOXAjiE+32qJuLvSVXWqDzK9a+n8rn1teE4NFfvrpxXDZzorLMbydSL
aRgRwNtottrIwxFBOIgZAFTNtmmRwNGYgUiakCC5U3sRDb/eB3gQgwZT6qS0/tWg
i8PKyozM0GY2qAZWP6zafaqO8XiqY6ETiqdrwECKiT9OiZ5wFzaQFqrjlVdkflVf
Nq5Ex0Bd7CNItYVa35tFeLQ3hcgH3ttCkiFF/brTZvLtI90h6ZeCTTEPDcEsOM0k
gjALzLSh5U6X/J78594YNGIvpkyBPom9eqxrkhw451TRKlD2dLaMw4BF9bCmQKqN
OR1Trw7T19pL/ujv6Dt6KmEw6Ph2aM/KFP72yA/sb6MkygydLNHkBJOfRFoKNDXr
NDRkCZZHJnboyH3U6nc5PLZVqkoTX6bzcKWAWG6JxYn7s3O488eNprcdFHD7inOi
q2kHrP1uJmsnVeSdiz5+YmgIFxXCp7OdwG7vRj1lQ2AZG5ny2Ke5EGVIvpW1V28X
ZVIFRGGZXe/uOzBrnfwk2pguxxpysBEBXr2s3RpGFqrlKv77/pMR0MZsHutyJQfL
Pjk5ipeWKEsiWu2kcBXvltXNvQihCV2H87JrQQwHaWu77LE2lCVRydZF3ZQbhgI2
tcqEYz0mOivBVJ5xLjPG0i0i7fzt04aICY5TtAwhyaYAyx7RNeSkvw2epQyK3jZ9
FdDQfeZ9yy3lHmlEWQvfp4YABsbNcnlZcBAP7EJbMUR0K3zz4bIYGhX3+ISaVWjX
lzfrwt0b4GRwegp2/ZiPdi90jgFiXCN4kaWy1ASbcBemSFLpN4H7o/w9QjznJY/5
h4VOGOB7BI3m7JQYBmAn3pcM3oaraNBliIwUJZmZmsQvRUw+gmc+2wCHliao9mKT
y+UJvXx9HI8/E9YrKebiC5xZpaOsqOBV9kRY7L6xfTdeZCMwWAszZudOdpR65a2g
bRR4eCPvp9xU6RT3y2bQt90krSTsr0ZyFStMXp739mXwwUcAJhIVOk1nL+cgW5Jf
sa2ni9DFxzo93508jhtWT9UqwaAkqVFycpETPVb0xY59wzW6lAH1dZhHuJ3GHBmA
3DiDWE/qy97kPKkcunojRArcaWbBbYPaWn15FTQWNT7bjJ7C6NfrzjtyGAzlD5ln
0Vop17AtG8SLE2usTOgYdyrWEhEEWW2N1MxdzfbbV+7pdENWABeBoIhwg0KIHkYx
vC1dE0osAleOOcbX3DlFpaQLbbi2y8k9LQ4Vy3ohvzmgfutKu1MTTPsdjPipF4l3
o2rS43eco2Ig133NI0kepUxwBGMIVi1CvP/SamLnF36kCJx+oAd/klD6Tcvf0kLX
OaZmB1Ff5CSVDSXg6OoZ+kbLgQIKRaKBI63jMpE4Kb91x2Z/dDwFQbCKnPQOcrGX
R6dcQaVJ1hHtfnmOxx5DPqzko8WdvphyIPXN3DEzcH0zUXwF60IlYz3iCBECockK
p3PGEWAquo/wGZJcqukV17bK6X3GM/AJ0A2rLlq0T789y1QI94k+M1DoQSqJX32z
m8Q1bCdHxlZB5+tBjzBGowaVQAUaPWcVEgMHIN6MWUo5usVZYMItKGrwwYjWKe7E
TjN0I0OwRFhkbY0FazBzsHPxbhH4BIp33s10QrBnzCk1bIEjjWH1E2T+ePn2dQnd
+07dZZSPgIMYYAOlymOaX8Ps/YbtxXx2HB7ztzMWZvC8iEp3FiVTtWgZHceSV5yy
9O+j3iGA7z0Cqw5DhGPxkNyp4c0teZ/u1ZgiFOEyN6b572mJNU+/4W3tz8EBiORQ
sOHWagvKy+cIWW7ZvQdck02/Apj0Wr7z4m9Vy/8aY6E6ZEaQb2wsAKwpaOBP3ePY
saTLBkw/gi4sO6wmjqPabnAFWC7RUvIOf+JMrXoAbrPvYG/bXfMbIPz4qDpKwRfv
Fl/vc1eJV+hXqaGgUj0lxhRwpaYMdWdIVsODb8J4yuKqsgiXv8wqVlq7ontdQAgG
RIdVCUlHRre4g9uhdMKfH9K2yx+dj9Him+lxrxCvL4DZcvE2XLWEpAqneaZzmkrT
wv0gXnvytUnGSkDJVfYisnFrnTYXCDd+4wSzUTd8UsXqksMvmrXcePelnvecKGfO
GsxhZKSha5sAEQmMAMiGSFqRvzTBnTYNR9vR1eaOOsqreYHkXkQo0oNCoqPlb1+y
C6wAuGIV3hgOhSOkG2vmtAIqrWCkEBwVzT+XUNngp1KkXHZTTY5q2EOMW8R+gQqz
4p/wpn9f5Gpb5tIkduewyqtLP71oojZoxZsfljA94I753s45UyfPLXb82J3sX985
6AbJu7StDTZr0ISSttB2vUMfAH+lGj3rlUg7YkAoPzMIVu63xggD4jEQYuJKxlaZ
md/UWnxAF0ZJw3IEw5EVMB/nns5Muym2kJLAg2sJDIuSRAjbMECAY/8OXrRFtyrr
q7pBlvfEd4hjjoUu9pwwVbc8Dae6tooKWTfaHY0UjKtd34RaBcsTct3Cxj6+xpDh
ntIOrKTsO1wRI7LIzy2HFxsG7FfKxMD+KK22jYXkwIJX7mvXdJtZLH6XhIv89sk4
g+CHCwKJb22amfMh1GBlZMkL1y7Ecm9nyQs4a4hPAuLaCzlxlPaW08sHQlUtE/mi
qC4wtHxt5ZVN9LYn73LXGjaFDpDPzGRBALNfjCW7MKt16VtmxdRBIGKxdbmePcoI
UT/hh8jU8c6c4EKn3OV3tuzhXbfBAA0XtZvVMR9bZmSDAvl7sCiXDAj/zjLODLO3
mfJ+jUiuO8eGDxyW1mL0zQHEoglV+sFd6weZJUL9r5CNioxfIYraHwD2PwPvNcrh
eWMIUcOzhpu3Wa3FhPAYg3GbLZIyEL18VeaQoVwtaIraumYbA5YO7tsmG7QYiXxg
161IcPl+MijaHAHHRpX7Q0zHXDTuyER4vlvuHFej0gFdhXn60SsF3z8enEMzlXsV
ayNdLtFXdDGBUFCRJtPWfvK0M95wtFhrYTdVJJIzQRVlIPnCllcPZCi2bK4Wcu61
coqQ1OoIKnsX8dC+UYA80TXGsfJi1RQ0u1DwL2NjfsoMgD4uZdSoRzXV9X216WNh
OzELqfakRnfsGIzkoKmG3DMJ/YDmHJh8NfZUNy8/ZrulxNm+e+L6JcIubyEKyxLP
c39aa6crWetin+KHx3Zk32xYSXZgKPSpnzqT6V/3PNbv6uN70JBT3i4ZPONR9r60
NVcg44/ql0bxp7ojdqMPs3+zbEuJAIJaYMm7lJjFoeVoWlUaDfvzSpGR/xGqaU/v
BDc38BbFgjWwq/lejgQJiBFIWyitiDOjDC+OBUeqTYJ2yp2IWWAEyY1XthOaiuD5
lr46wV4a/GabH3YV/VzXmRVpwEctv2KAr3IdKXtCxDyvEmcqnwYVvThYGNssAH96
FMnj7TpaTY4Vkm1zInAN8AeS9b6xPOM1XKfi37WXxaxD8IUe0XnS1nDeK4oNb37s
pq3jAdngU2/tJt5+1cxElxX/uSQ8zfNUiVetvMudl+qQIFDJPdpH5lg4olGq8JxA
Zusy0xsdUMS6TtYhE6I8N0FU7BcSWAXCnjdWa5jXLo+UZhvCYSPLuydmLvANOhRp
H4Lm5s4UHZeriXommxPAdkNdVUbX93vcKC8AxDRkojLcSyDGNQVDA/xgap3NH0I8
H304IQlqsot07kfZuXvltyHsEldC01b8+h9sfXr8Sucn8N2BwZFPgRZ1gfK4h6nt
jxGuJ8FfeKzmB1ye+sbOg9iGPRXtHVZpNoKEJN2p9EyraBBEv9ClQYXpOWg7QaL/
HziPBxS9TC1JcZmyEMZxKFBIfLYp6JaR/DECqQ613S2KHqnf6HUFbR7BszM2P4Tx
Vi92X8jFtkc6S4fi2x/rWU7JcO+jdYqIcfO2boRsH9uq0OWqdbR2Lun5NW+njiQK
WLOmZzw2WgyBxfxrSy4OkrCk6gVk6fqDVEfxIlKpI7HrJlwFwdjdeCWe1YV258U2
tXFDOZW+c4jYu1txO1DPdtrosktwtul3CYn20rGFw825+818ouMu45x9S+dTA/x/
MH9V6VUMc4dCM3CGcIRMK6NCDXS/ckS4GE5KFpk8A1rBxMrrpILmrWeK6rQZUCbs
EggESlIaDtWFixxDThzjo7htFZ0HmOvcIg9zkhI03YXvA6w9ln5BgauSqx4LM3fQ
04PW0w0ZIW3hQPS8oihonC7yqFeUFfsGWiLD7LhreaBTejGoVkLwKTuIl2oKEnst
QEQR3EvsWF9JnU+DPF1l5prf9cUgEzNiFkQ/VYY4h1w/twPwiJ99awDMO+TZn1lw
VOlik/ANI58WneYJZKsCihPTv4WYMljw+XLFl53MJekBCRw+8XHRtbk19VvVGntR
i9fD7tQQABac/5rxiWKNIzgA8QSR+AgmfRaMlXDLNKK59FW22PTCttd3Sgq5Hy80
re+lTpOZ5iLnEC4kTlMq1fZoLOjC+q7W7qpY8tb8a1f0SnS2iKgs82Sv0TaFDfYb
KGQhqJsn6PizhcmyvYyAbi6tQffv8bIRPKls7KgjjQccM+jt54naKyFwEJZZwst/
cIItKjx9ej3hBMpscETQ4lT+ChmfZIYph0Del5uRvCiBDv93joH5KpzEuAlJOfmG
s9j1ZaxpAizRXwr7nMGjLCzs8ivu+4WJKbct3jnO7DrcjsmB2mR5QAvpvZMp1oqa
/8ue4S89FLmgivkSADFKC+h9CiUX4k6GjFXoOosQ31oqHtYjxTR11Q/BQlDwFk5m
jVuugCxfT9n+gAwtUPyJOUpw+6ODHiZb9f7Qiw/6KLyOZLCpWzEGkfFyV2SUJdz/
z8k26Q76wrRwIiWpA3eBDO4O/sHrnRd7fIrqAIx4AFR1d/MOC98JdgyM29f4TEAG
IyUGjK/8Ra2BgcB0uFpsf0fzT5Z1KrQj6kDsB5/HElaoCmTITQRD3ibFS+MORgDs
9Y1yYpYu5r0hheW97KxXcVLvXctnAirAljopgwAadFPPMPl/LnqDcJvVylibBh/d
DMEvU4azsI4OJqYRo8IfCtzdgoQxr6w42Rl34bDNUoFQU/3YEdCjm/5brxxmRPw+
J7RIFaqFK0nmJ4B2RvKZzLBJTtGzrtJC3Dk11IH5xeDcWLnMz36ew/W9KBZVJOZ/
Tji9A9TsT1+lUMpRxIBe6MSepBAv1FYtyEsN6e+XelcNhOkDZlXtTS46/NRMZGQv
W+PdGJnO0KaUAFxMjbiOSTt0CpPiGTwVdk8aXdMjwLdsvt4phTxgNsHRTcbdlNC+
YmuMGlm1P86rnPFAUTWYyLzMYTk6ZhznUWFwsCYM0408p4o/vnqtD1PzvjwS6PDE
TjOl/kwyt1+2JmrZk5PY1HdBtaMFgznjVgCMRh6wcAkvu9RkY8w10H5xMmn/Hgc8
vh6JsAIhMLxsZmYE0Ied90RITX9ZEVqK5mmXjsWlty6ypEdiiHn8ojGFRjw+gof9
L44R1xILF0dfXrH9ny0i25oTYrlpFG6q3sA+ZXQX8o2RSrw4hmUhqg1bpEkFyPV6
1wJscU2B1zF0Dno4S6EQyr9LZG9qvf8FGXApnIdZLT/Bp3jcU9DzXMnrFthdpAjY
2kVFwTVQFCGNhqlE2TdHBT15OzVEN8/AzImN7whA0tdGgEaeLlRdZimsRVfFFrXc
AgcxMf8yC6egPj18cSSAViZ1SMxcaC1xJuRidwGLmIsxML86mvV411DCV9207oFA
234fOKlt3XOAyaV5rZh1mCnC5/z0YAUWOB8zcQV7ViCEhHbl5J7lWAtq+qA8g9eb
nj1rczQHCVGSKrxcYUl+w14kbCK9OG5hown9yPbbQ4zf6Hchldlxda3nS9uTcMoF
m1Asd5u/SBj2bCA7ohkPMGZyC9jv0leWKcLgux2yG1clB/8Sr/gxnpunnB2Wd+at
X0aUHMmMXTs4iiUiX3ONkRAFh4dM7LefcZAkKVsjKprKlEt1kz6+nyRLqayDb7kN
WWDXlVMQcmleBCZofIXTiyKr5T1Jt9u36BxtvX4d/SoizOF2HCCpw/jxD2TtGY2y
COvUemyhlUpMPN1gw5ZGSzAUAyGfx+iaoy8gNKq9CRnH0hwqU1d8OwjCROMzzYa6
8Xc8zJVc6zXuecRhFWEcCxkgHFeH49JILrx5N/ickOlNItym1RtvMTjdO7wLO0Id
OKkW0mKL+HkuX6Kz4z1ImaiObhz2nkrFlXXN1yRWarIiBWyG9NV3ZEPKvQpGRl4j
+Rad44PEqUTOKOHzhXOnnEVBrojYn5yYWtT8BbOe85wpbMX4MdVzBnm4TNwaeG6I
oDf9aAf23t7FcScwH0tiQD5lAyY8Dl4CQS9aDL4BkpZlIhiadxFeJTLfYYW4wV8p
PbhvrAS+Wd2ntAM0tXI8Gz0X0bqR/8oj0kC3ivO3uhvbpZoNU1zUJLQIYEJ89s4Q
68RejpExuUk5NQ5c6dssTJSRnfHGMswf2oxx4VFLu4rFFFr/Fvlc78ORFc6rF+bg
16cEBFHGCoGIqShb4qC39uS3aD2qsiYzEehCY2zfeDKq9C7A4+bgLrZf0gsVWPKr
DMLuOXadHsQBlfva3kaV2tpJbyHba71V/MkHNO86q+DZfkORk2e8BCnsFKdK01s1
zGVn1Rp8XmDoeZ7WqachdKjnDnrjwFz2Gomi0KzYxWogCLUjdCF1JCSN6UJZm9G0
zOz9Ph0pXkaQzFM1spdqOjjCbkmBz0ZNroxrBAM9QQXX3a4memLzUw6gzQ04HdgH
+la/B2gmf82rFRYpjB8nXYYIXpMyC11Uh1IOzg/9NwDXdEism6buq4Ulp77UXtMm
R9gsbvnUXpj6DJIbQzI4EBLOnt7/binWVTwe+LQDo13ElcvANKpovIhp/5mWtCOZ
ULC/evtvCgx4lj+/VpUlFXcNnH623CqGuJ5SdO71gUDrrPaF+M0CvTKAFPZpfZqE
6FZD+IC9wmfdZwUkxm1jy6pxcl5cAtH+xLBGLtOoUIhw8YpTIKajszAtA48Sd/LZ
n1UNTU/zEPRv97RTVeW/We2HR01gTE0SWGqhBE8v74iQ4q4hXAcLC4Cg7rQaWetH
9+lsU9a2aqxhzgr2MhxorjAavwxIF5zH9TL9UQNckeOYL0/iAaHRX/SY+EvnmVPq
MKI5wmoK9MkFP+g/PWwMxEyFG/vtsuLKcwPK8cn2dS6HVP3mPWm1JowF/1Z355xU
1zpReciyk210UDPtn1/6kvv1pMuuHE3ekFLoyZcDQPdHwSUyDshE0/z5YChI8Tfm
YH2rwq8TgtV+wwB8uuKlHvd6IP+q38pK/hKnmL4Yh1jKNNfsJKo6oR+x8zmeGUC9
4Fv5vHQAECy0nn3DRAxYlBuZ6shGgPxASmb7AYbp7PmJtXaW0HZwJXQP8w+9fxeX
jzraQ/vBYnqp6NQY1nJbuArQ241nZwFRo8RbOUSL7Qbhjqvi3GTDt9RKVUONX6bH
IdSNDm4wbc5m+3VRToItWdU2flVjkf/TgrkBUeYj4O9RbD7h1/tRTSh2GOk1CQTo
5CuBjQ9AU54O5judcKc6M6oD5by1ar0sVYcPBEr+6iDjSOpne1X0Y8FDudJETln+
A0li//AzLmp+KOrHiN6cX/K1mENWh2ibTnB7BZx6HW7oG392FwhuuPKjRm5P45g9
vf5vm/N0CACgG2ZtXehKay5eMxVhqi/OCfJzu+OVbWjYKQPMxjJaZF9ZhsKgP4lT
jMrHIf8pibZuRE0//rucRKs94RHwbqO4tDE4kn0DXP/Y7n/gJ2b/RG3o2F9IzuLV
qiqy7+67VJUcqli0j3X2MsJ4bG5CPeG1r5AQuzAUL/ZcnWmLZnW6IPMG22O1PyRn
eAS89l4Vzb05A0gvSst/gvAl+Qd67TdCpZvdKajEn0yWIpYaAq9YNy1csj9zorig
bTpyhJjyW0VmhmYq7Y696t1V/WRbnIhB4Gg+kpJ1//fx1UZWHx1QGoRZjmu3qrc7
7769gIiBZw6NsVBSkeCh5TqLmD6BJsdulcTdTpKXcRDhUZ5AUC6f7e2hJSer96fg
yPBQWChMPUDVxhI19W9gm5SSV1BywQnq1s98zsZGOqtd486BS5O5426aCgjBJePr
PgizlL1RHufaC2WfaVlnqoVzlwNDckFnQgdWh4dTAwgLUUtySaPPlS68RzOEoZEx
6QdKC/giCszbyYJAJPv6dZmW5h+PW2iaPf0xUM804337PBPsMn9WSzK/ErSz8tJ9
LgQx2tozpcFr+4WqFwkmaT6a/cVgZwVhD5kRrPTcd+aXSn3TPurW2R+/J72nTo3m
V49xX3ftNHZ2zyyZ6on/laWuty2MsNyo+VqKVTzZ1T+omUuUir1boW+KVD0ROjTs
28eX3p7gdlVCK7Rp6YJeCKJVlD2j2AUobGWG6a7i0FPlBX8pzU1odkMN1XaquidW
BdOW9WLib9XdlsmFmpjDwVHeuJL6Pa9ajSc/pU4y3SOIJgUUUYLtads3AAGi4UA0
ELWd/9YvpRWUw3cYbDWz3yy5mU314Dy0w7NYRUwEDPr+8U6LEPGEMCIabXBxdq7K
P1PG/bq5HZ63B6osLYGVF++M2UiBsWxrfNIqhe2zPZcTOSPT3vsXs5+Ww37w8I77
PuHEzE86PcB2Kp0Y5LrYhZIjOgz+XTj9ncMbeDR+ola760IDBtmY0BB/9N7PmDg0
e7nFJUP6E5RfCG9pcW1zR0TYGEVI4DgHBwxSvLMSaL2UKzeUxEIXIrQApLcN4unK
jE2JkM5ZWp6u4XC8q+3Vw6W+Ys7zDmrgPVXQN8i/eV4BABwhAO5gD/LK8EV9gZz5
9Ghsu0XTxU29mfsAINjV3HbCeh9kSWcuRx+gxpAhGAAV6crzpTk26rfOnyxpOKbk
E24IDUpkN3ekReTF5V730CWu04l9ctevQ2QTIgHNb/gXpxkbC9QwjN6MgWm/8P2Y
SO3mztlU/izjZVLbhwn3LYHdiKofzdhA8Qhuv3brZnpLtZTeAGsfgdlb44DEDdVP
4ivjZdEgGLprcmtZJnJl9ugMCVnGLUfuUQNkF88LVvhElyo9A5WJiFhiv/rzTe0/
f6ISTT13eeqXAPX+JJpUVcRwywplFU/lnIZQuQyTNb4V9C77gJIvqdje/Xv/R7Fz
4/84Y9UdG0tdCFSHNzSzZ5+TYZOtKyDKNuzpaQWrHCAPk42GUBdsY8o8AFNTcHau
02RKlwubWa/BrUsmU2boMXXYDE3gEJvjWJ6zZcqmjAbFMc7AKLm+K3+COXwxzWeu
LoY65/MedXyufcYLkMrQmHRx5cEMDDWnd6/EEI6p04qbsSkY0RlF9zVyY6GKSpjx
wU8oODYRRyl0JK2hlrTK3OIOHWagEmVo4vADqQbNlRZAyAGmb0rHrfOXNzGu4y9m
2pnafBMfPjFYN/F7hIo3+h/EDzzJYzuOWl2OKXCbC+FCsyhXjD/eLcrQaewl5Fv+
FQGIqsk/+RJIsECaSiePrBHk8ztSrzzrNPCleJ68jKXb6GMPzXz8kLej7UgzK7Mo
U2pNeGuO7aSN1DH1TLNQnaCK8i1fg08LvRqO1zhf/QISKQhidvuD5rJJrLQKLYTN
OwkSuNrG4dzOBlpYatyuA2YGAVxWgxh8sYtVPq41uk4Kw7I2M7v6QgW1yfAJU+MW
60ZAUa5DJ0+LGNOB6/Wdn9Wen+IhHg7zYMyds+OtrUx9cI4n7XgK6i1ZzXrUJZQV
XH2G99zZK7z+wEZY0V+0gl9fE8gENyDEgmyyrHzBKEBXJutu7Ady7KIhJg77+7Yj
FXS0dOBpCLkLn02QXVSpf+MWdwEHvBmPhRTjKJQTDeomdhkT4qy5pj7zpYVfaS+M
+UV5lRQlsbGBtV+idkImL+vfFCn31sTNz9R56a4I67ux/JhYhi5ALcMMi0heiulQ
ZOHc0whSZwpoj4MNnH09qe5YMXNwr2ITruKI1R3ITXu75NT4BT2fLWfszk/Jsopv
8WaHpbP5U0neaeL8neGOStAnULa0ZPdoJ0zHHiyJDq3VBVYqHEhqoCg/FG/FgJss
bXcQvGlDxYGte1QDjLAGhIgOh2o4Je3Tjetn5LJVEXeh4R604J1AfOE4OXiEkAB8
KCUKRVHgLh+/2hyam0926NvBRGLJX0vIcD6eHrLOMx2l6/sU4u2tLvng89ZL2YdF
pO2AGiC+hww08/sAKnyUqY5H3Xexn6Y6+i+JP8ZXhBNF9N3pLCNvFaQ7cGNS1cnL
mqIdZlGYDBI+4sy1d9GMzLDwrMHXUosJXnqrxIfvaNga4yfuBUHKoG1fq7AP3VQR
a8JRmnG8DDFMOVILtv5VFzCUZqHXWvQ9tvf5TWhxuWogmCveCO2Nfd3//oIWv1ff
7MifQHY8oMjIuBIeKpYgjugBmS4FbWRaHiLnBiLaYDT4oMiP9tWxuAYCNllNMbf7
EB1Fe/61lAkQeadPzWsvr4PkzsO1J1nEtk1I1iumbqgfIaiyECzmb3cqp55V9/q0
VHFt/mLrrAQsDalYSwkuCEsIR/lg4RL7Ds+f65lQjKJ6s6L6vVgImhuQTBpCrbXj
Qi6LUtp9lI+qzpCHHc5alNJuFZzgW53fwN4epbvwW7JiFm89lFqvwFfZDwG5K1Qk
FFYI+QMlGNXVP+FRF1Q4i2a9CRj021R/2rRal74pSIxTl7E+nI9uj+p9+ubgxnqr
aNyNVngETfelZTyKwxGydj73Vl/Xa3+dLJhJUMfS0eXtJBl21y7ooWA7v01scXnt
37xCp3/s7vry8Yc2EK0yjREdCgPkwSTa2dMF7yGh2Er59BsFNEHi6nVtrymknygu
Royc5Jn00huzgRf+c1xWRoxbL1KaJe82fGEPl4YtEyXmpFJAMIcqIv6BRKpMfrUc
04RFaK4eSjNlhrs5HNXMBgn7b2BvM7BC/3MVihOR1tSU0cgWfEuvi7XF7Wy6FLnx
0SoB6tCgQRg5pqP/9SA2di4GQbP4evdzAn2yjBZBNHkNyUgggF3O+tpG/fQzQCf+
oFEJHEqUJCO5/HOlg60+vg7dL4wKnWijURK0sJcw0iLszARlswDVg77J8u4NTaUV
p1gjmkCTHMhYXBYieyhvQlOOIWkGlJpNHJtnjyfvA28Eacn+TuQaYG+asdNKlq6d
/qsivtKNN1H8EonG71v0ZeFhtW5LaKr80k/8GjxldcoJ6S8N8N0v1eF/vD6JTqTo
QDai/s+fpfeP0p4IGU0fvpuU0GT9c2af5v/oJN9+3kqCUcSZzt5ddqv+Rc7IHrzw
dD586NRvFneUDP9wOo2hjtzqgJMdQ43yWGl02tdVOchlP/NCRFUGvaO0ksi0J/b5
A+XCkDJxHNpoTJtJqiqp40cHbbeNnfF8NP5Ln04+CTqhqHvGouFCK9J/N8Jpxcod
tkDj1RVLkO/eDFMsTiYnxW0GckEVacHYMLnXJNEmfh87LlVskKtX9DHSxpJuYwxj
OgthRW1COWwWkhOEu0euyAeU2oZ6ih8jiqmsZdUQDz6Ancxy+XoCzDZCwnEY32n8
cCy+BJx3GgeB8CGKzuypCRsJHqBohW9rsPO6XhG7tuDYHjiq6YK4KjrGuWbLD9DY
S/RGfDfFxdjSNgVYKEwG+nnhvgANI28cgV30px0ogdflwiDWV3pqB1Wz0fcE+juu
0aIADqCscQ9A8+wPTeEfxCdSD99t9VxzTGCWZRblZzc6CeqEmWN5s0mF1i/PBgWO
36U3vkZ76Q63lU6q4WZfLK4E/A5dLRDo+awcQavjOplJ52tjvEWH8zgWgdOZmIun
mwGEzOmQKih/8Q2zUVUaFABsRhQS+YELMKNFIBwZamOCDF1v2JCYT8cnrJJVlbiw
63QlacflohvdW/DBhP7pXGke1I34QYxDA5h1eLaPhZuDhIHbrJ6iY74OLo0fU0ww
+Bwj/dyVS+JO+1qVXi/jlEd8jJ7h+ah1o7b8V4yE4x8zxykOvFDUpe5XE8LbVFWS
q5JJt3NcntBD81Og3oV6mzn/P7KVdfPXusZfOUhuD8xy4/Q7ZMH6zDNaymFEDDFM
48CKnTGW8PiBKSrI9SY2qx5wa304nm0A0RjlocL8TV160soJ65+4kA839YJIOnPX
YXIRNeOvo0mKsy9R8msr2ZLWtXPoxdSx/Vl/fxoYul5rU1+K8gl094Af3kgaJYu2
M/j+c/xcaarWoO/T99OP1SCBOK2MPrfCY/LOPUp2zlvjT7SUDWS8y1YMhpMsijWZ
ul2kOf9FN7rnLPcpk456tb1fdt4DelgQQ9h2kK0qeSoxumWMK8LitepfWUO1fyOv
fI0h/LCENj6HwWTILi8AzJdkuPMe6Ja3N/ns9R8Fe8MtzFxwrEQhXYbZZi/dND/h
gzCTQgwZie/PK3kP69QDB7tdZKrsg8d2Mg5q5r8SHRBOVfs/3sFEPYbL9Gl4t03+
ArbjKSIg6nOAMI6MBTW9+zgbewBDNeVrgXoZ9ZaTxnlQ3eIWBCSUrcMBpoTYbRvo
gVkvVWE8d+0bqzo1mh1YlrG54QdhEoCUTjWKJ3q4V550VQgXiXDCsVvIxGZD5D+u
vtzuaoUpCzRAFVyYQix1R4CWp5pNUlOdCK3h0p/bkOmwPovdimj7GV5f9iW3Yaau
zvcW+xgNM2EZRYjy4Qc7WnMAAjGzaYV9tBIroAs/SFPxqnwRqbPaG+6v3LWl1ekc
9X9YgKvysEJcreWI7uER75gA1gkLHrvVwHh+Wb2B6mcBNJjMEcFDOqryTr39tdkP
+hQewbQbQJHWPmsZlE/yBl6CDYEhH5ZpjYyCO6DQuz6xAwu3pSyej4wdpyXbu0Lc
y0THeRn90y+Jf+VEz963F2o8Q+sM1lJJb7JNVhCYqv1FV574sSO3nDykzZ43GllZ
Y3f0hs5HskLUmCM6AeUHWyTORJJ5Xe7u0t9ujTEyXXJg1K4a8vNkEdvTQ74FlME9
9SDqFMObZ6Gl4QCdFHp3VqaZwpfwNH21WqkmNUrM3y6qNxtVtIFJ2JzlQ6wNw6Ws
quMhrRLLGXePDDURTJG7ZqGIVjbJ4v7xZ2b3J7/ZQJzCk1L9zu8bDyuJgZLW9xNk
I+TnGcfiugs8m59jKqQEeaUKXpqaM68KWHzFsqbw/0FbAts5NIXHzVYDKv/ROCqQ
JMUD7KHHopyO5BgQPWTMhN3/+vKZP7kZ9YAjvpvyOw97iTXT2LDho7t3PO0FrTeK
YfsfI5m0y3y5E2e0Z4qSmezBMbZVLMLwl/UIYiJEvdTHTvVQ/5YbQSCXZy8vIA1Y
hhPUtV2AxuXFxiRYErW+cDmCHjH352HLPrviGsxugViykLr429Q+Lr6XOVp30Vac
fqfgjoBpe70nDRhSnyNcV6g4GL3rtRdSkRam2Z51NksSdUyobepLJ0Kl0iMMWyZD
8ly/Vyq7EBjqaEec5D98x4BIE2j0qMaTSleDJMwBlQcfgySCGt5KPybBNiowkO6y
1ujNEjIye4wEocZrHNtviCF99o8EMu5UPYKDda2/XLaJr1PhxIyJ9hGCv1uPO6E6
QrN30msATu7iKajhYO+nk+K6dCP74SiSVgle3GaqkfOHjMTHSdohtGRANmBYRf7r
kYO0PufMFfKhl1kONVzn+OqcJ5ITkSBxFhlmTa/u/nYkOffkvSlmoxpwvxlPOzUB
UQWH5eZSXaZ7DzB6SdNPvtUiNAlkehQu1sizb8A0q/68hx+TIzAVaJxGDZf0g9YL
QfBsVMcxIs3F7/DMccHwzug+OdCF3edunAzyIhcidOE6AVHho6S1eawwzhTZ+dJS
oNO0ku5IDwHfuZK7Z2f2NVMpoGbz1V5yFgMhSYu0E+gk08EVzdUk8FWDdWf5lWNn
nJqTiUT1UqihbAUJiS2ni7L1Qo4QVwR/MihcNkUe26GlcesE5Ypy9keANRMyuQ5E
eZ0VUwxwvdSJmVS1g03SRhN4+B793QKyyVZIP+sd9U+jYkyJybv5mg6t0T7t0mQR
vk5ouVVtP+HqteQcrC+ME3SUKsJ3xwuD6ikeUL+EpZVJocsDraKWR99Z8mhmPAzq
/oibR41kIKTmOoOJzhnQ1JCAHIegRZOV1yfzI7fxomV3E0fU6KFPhlC+Jh92PA4a
exLdM28Ab1WTK5g68WshPBRrSRVflMOBruqEPmmlLvmFEIhIT8c+7TT4S+uZbVkv
Q2MBulhYBOMHQ4e4k76xraanGlyGonarl6+diu/4WfMV53wqoSGStKHMthj1hjwG
UhPE3KQuSfSrjakBi+lxmL+0UYOa/fuT7JHztJ/LIWPHWiEVFf3bBLqcmHmqKWlz
OYj5qZLCwlH9S5ixCIe4TFB8dpHE1Phz0WfLUBOw3RjbJKRG+77eYELkK7yv/x6+
se4KMRIa6ztfnjhEdAG+qHIcQiSCWL0Hmu5MM/5DA3uqkG00eisesdyCZWCzITHt
b06u+s7SY+u7coYq7xaTxYl5rhkljIcxEuylhrQdD7f8sGF2sw5qlg2n741pZnqo
0Qq6aWOvtVOJOcduzbuulcBkT+0aSzLSU4aRiM/4PYv65Z9Qx/kaVgjZELwRiRsj
EsITxvkTEGZQcnkdsEfTL3+0V3pKV09rufNm/00px9QhWgRKvrbj2Qe4Ym/vJ1GX
5dwTPe2fGP8Oc8wffpk8i1ZdKlwisgz8zBiAw02jd17yvbTGl1C7NxAaMEixkReA
e/ouwmYieo0E4h65ElvzJrr5rQ97aDCAwKEg8A12TUQ2lQVebrblUjDgPKJYVTG/
LV0/hb/89Tx6vq5V1KWtwMJAQAppT9V2eE/sREqovc5KyHurUSECoDcH0Zb6a/fH
QSFTMp4wGHuygob2gBqHvI3ZK9l9OeFuGsRB7jXTcuegOwKTmr00H3Tql2GxC7AB
lJKe4xsleVwviz+iObN11HDxXvP2B0CkAnYGuXPaLtm+XDgR23ke6/MyA5IUGa8U
4Wn1gp9IFYpbKzPDRS/IU9HuIGcJ82nAD+G4fXw8zSME7AXdTNBleH9t2seLEGZk
c5mJNM8xmLudP/GiNAtj3mg8X5IZWZfI4QfE14BU75+mY0t4kTB9l4RHJ7e8GTkR
d4Gz2B2LZ/XpGBtmsIRQrPmeNy6p31d6xHlmA71R2YX+Fjfa0sQAUBWY/POCUU/E
r9uFd2ssjWnc5ACTJYxr6Lt5ee77+LHdJYgVc8PbXflFqznd2t4tZHv1+aWqH40o
k4dJH8/KNVdVxxxnac5X5Llq8XfxqtXAiYo89bVKQ/3mjjeGxPuA7xzWE+4tNCds
xkYWl5Q4eeUHu/gIIiVrHI8+XQvLwJ1L1GlfYsYz9gajKXffj7Ul3kyQOKInSz79
N8aD4cZGpOfSfdjMnbkOd42vmTbzjUpoVcy0u7wY7M5w3I376dNMwRryCTIoSPmE
2tuIo3QUFTu+HRXuBZmYzoZCrtdVCr3KiX0PaWRGAd12J21UXhJXH0n2+PEs20Aq
0Bw+8URFchR98QkU3/TTJNSeV60cvG4mDozImWlmYna4ttL8qkp8bWslcYpSKSGe
Nm1QIV4ofgHacoRhk0N7abnfvRZzZ0Yq+gCzzi4stECUirBALuzW+5bSWB0rTgIM
hpzJSCB81MAXFC/AiXS9gbTTLYselKx3Sx6xn77UTCmv2v0/gE4PWnXx9rWhSN7L
VvVEhldz8M8oQWz7wHaQQF5hlde/lEdDOoAgaq3fKHOhw98hCkT0DBxbepbX0/JO
s4ohv5HI6NEF0vZIVqtohkRgfTZxLtbjjurtKg9wr6sYm+oV47ryr5kCYnPxif37
xQurbWHLiz8NIk4zzVEhuQ3neOnrFIvNUZhbFJVLXnSNQmkA7sbFXqGQiiJyjE8x
XB7p+X9/Kad7r2U6Kg2JI45n0409+x6ju69yhzbTyG9JIHvcBDFjUrw6c/P0mrsr
SMXM5lVQwkdiSvKc1zfJ/Tm/6rH1FdcR8YrSi/qq1tDSD8IouT7/5GkwAgBwviYi
gOkWmdnnoJRzQ0dUk8or79FREULuwKhNQWCrsV+f7frD7NUSw2PdkqwCm/45gf0z
UEbO/cd2lUmol4e792CqOsgyVVwQc3lDfHEsVbgti1C4LaElGQg5V85/qmfF8gRd
5zFg321Ju/6xjqd3P0dFzF6mAkKTV+KTxd0tIDqki8X+RYsTOE/DdOCXuD9ipCJ3
PbiUn69WGRDPnpCRXWbiwG44CEQizMekSVyEP6oc4jgNHb6sT8sIyB3ucNHY4Zpz
0VcUgFwc+ModRqReh/FepxP/+AqeJ9dErfZZbiyNtMtVfrOrGPORNkgJas5OO8I8
BznJhTlUZnowLOF/1CJOjz2vz6mJq78+Cxqec2qX8gpTosEw/X+YIUTFUajNagOh
9DzKH4J4ILK2qs+Tx2fCrK09llJJQTtq+Z7TYHxenzul/vi+R5BHqvhTZIQIhuWG
zldHttAQov6xBd+FuLoUWB4g9RgUXAR7Wlk0W3ffESWjew0nmtJUA/FyYfT5g/nn
0uP2zq/sZlliLSlXZgYpvqYWYDwaZoQUvt2QGP/chwJ5habQTySPjgyzbeEH5aQ3
ACWS7TUQfwIFIiSLANm64tD4F3hXoRVDZw4rH2StmdwwmJVqBk8wIkNwc26lf/CV
/fw5SUKhf7f5RYSKLA1gPLgXhKVenB8sfr+5AYQN2wh424M5H8DLF3ylNg89q+fa
Yswi/9zCsU6phWt5IAPnZ61FGh7SzzxnZuUAIF9X4TZcdPekTxna967KWWzqtZkx
+ubUjactCevvEdpH7n1ZzEVaKv84k3KOUguT9gS2bIyOu55LuT7frseNn9JGn2XV
vPJ8Htmry926fKkZmnbosbNniorWpCI+juRvwh83Ydom7mPBL9EWqIryBC0pHqNR
OHhWoFHmTFMxK1GrtAe0RO+/63gI1HZ7TlOHC1KBdVkL/nqJdkyP7kn6LjIFwOrY
KOXIYfesnPQkHBMmbZPgoHAggyeBoL5/h+WlTV1l2nRKiRFrOr5L7YYMbeN4nkWS
tYSb9tweQXm7ktOZN9jKqyVNlZUd2GaE9QQ9Olyxsorq0ddq9UAFlbSnhtsWC09t
4LjY6JbYVdvulBsmOhjo3/Mx+NcGuvuusDiqJ4BPAI5IQM+sGGQMTK0+uMfs5kZO
h6rndjDLOQRGMyEYqLrTIyYmuu0iY5PpPjo14BQBDrh9dVB/bC0BFH3wGRI39i2w
zUz9zAUnAOE7UfIXHMav4lM64E8gKLB4L3N9k15EKvCwRFTXsyWCNOq1YIphly6r
Rojjy1tW/I900MQVNnb1PsOIOOE2jov9tfkrxsx8nmwcEic3NndePx0UCEiBSPy7
9LeQCiHEWLl9sVn2YHoGs7rlyIOKg/zubhrL8zVO0uMptBhNGX5hnQgqzoAmvhiZ
iFz6pZiSFByeydhRFCX5x7LUeUaq0QqTwd7w3SEp83kSPuYGL5CoTQSLFt7oec67
XKUQm9L0bnxAWlzbPur1SAEJSXPKB2TKwZD1tK0tuSWQJWxcsTML0fASSVxpkJtL
fUDJIFo7FWrm0Xs6axIPFFKJUvMEs8JKH202QNPAsnYGPoyedQOPvUtXHF277Yfs
kn9IlpcEvsJVM/zxE+1kgQ8DZ6u6ieWcn2Bu/oczvQihhi6WCmt0v83X1CWaaIaj
OVzUzAGQicJ1YuVq9BEwxPW1/nI//5yDSeMtJsULFgP5VgzsMI9ssoFGDr28NRI2
/RUMSCFjTOAO8xkFBscKwry0VbMVAOhsg/8S0cDn6zOvkcxH28+tKuC+eLq3qkQ/
EighNyxT/YmDah5RIAR4D0QxQ6M0w77vXtY4sXPA2KS9oSe3DeWXOGBchLNUuKjC
HyaCMJAd2ZbA7jeCCrUDCjN03blN9lq3mkgi+5HaubM1XFmK4MaWgh/3HvT5HZgq
BWbvRidH4DtQPhGsI8iqT7gYMyAaFMhR+LbQPuCtokKERWnw1+Ie3pFC9brcT2ec
1zH8D03ztKBl7K0M4AxB+wwelnLohOFaKztstLWJLPER4zA7OCVE5mB6eUPDgcyc
NTJhEoC4Z8rt4DPquVwdnWTrjTWw3pXspcNqTZmPpg77tuqPFemXO2kBK7JyH3VF
6okNcvIeB25H6O3l2L11azgq3jmVXAgFfV35MHJl1PLXJ+fGeLcu46/MDk0dF8Mx
cPuANWUqRsKNZoFhxQyP26GObjHgS5vwHFFkzcZdX6LAiFT4EA4w2aiD4lbLx5K/
uEfXfXPYBAfm6z7fTSr/G77Xe6v+sUWL8EcUNnN1Q3mI/5XdyVSSdEV1AW5Q4qwE
cvtC3Zq7Y79N+yQtGNJ200Lk+V8eWSJ8YIl9WGj93RHazIo9+UcmCRp/05t8rxVR
X2QZE6f1HZ8eLV5QvrvLuXW3UDAB0ZyEZWZbJKmP0dvceR0INPCdvVz+5ageFoPc
McijyzkkF9qDzrSaJvT6NpK7MNB5FSLeArXlP5XSvs2PLOL9Hn43WyRO6/S6T5fD
W9OokA5LvVrMUvJzpJPct1tYbJcCoqbRTAFACZqpOfgx/3YixvjBAS6zLHY7Nwab
ZD0Nz1fQR0zBBS4AIY1VGwrvIYSLWcJ8b0A7Mkl2qqvNaSehtjIYBguFzdkVyG+4
Hbydz2I/HOKuwSXOYfmUiZtiIoYmp0PSHV8QDlNYuTb7NIN/FKx9GbeS6ZOp+FmA
bDXeklwbHA95i63Q8aXafZYBnZmBEioNEcqCGeThyFeUUY9EQ3muUhR7Jvd6J8TW
5X0CU3Hu94YWmm0rxhsGaO7M3fcykHNkTXVsuvrVDsH5PAQqDBstAD8k0eGFMr6E
EYn6sCw/ycCPmbDNWFXOEyr/ICNckeCvyApHUx7ca1jTRgdWyDbWRZpKnWSj6mUc
o9sxM5rjDPhdmmtCWt7vrQhZVgENOK6i372TGA6KnB+oCkVY3PqPlAM/qb6VhYeM
HZW1KYrq306OFJhNDXNQbYe81zS1BA3BBFmED201mOUEDqkvVDcRHIqlJzqg4Daa
2nQfnrhMe2trdRNrD+CHqs2zxANzpGlCF7OaTcTClUBkfi0GMzFBXtCgS7xChHvp
IYk7q/8BqiBnG2VNGpFi91G7DTvsu0uobJNAi9N6SJ7ifPBqmv9J3oTeEv2ntoAo
b4yTQnNmEoy63TubJ9t4GrOu18pEAPy3Jr17c+IH71mApQ+8gu8El6b/oANkqP0H
H81bVkp+F6wG1O6zmD8//xihi1jsgbOp6S77oqmveKYOqQLt4Th9HjorFucA35qQ
PBc2lhdieqLbNRZnV/+3q6FiHyw1jt1XQaGIp1vnThVy8cMZqxmJIe+LZvjOFnQ9
5xMkPHdU87wKR3aRN/FiDHfS8rZIvmPoGmOD1W3aL/qkjXOvcE4lbkF/Y+OVybKi
OBg8dccOWcKU/kWleQ+/S+tm+y+LSURjFEVSekxKi4awHojc3kKUQVBhQ35RlFi+
YZRcXJfq8bmg+jMoIA1GYI1vTiQX317oJqmasf2QWFsssdq/wdbP+gCvyRO4/u+x
f7kP0xX3/zf+fAqbeK6V1t/pjVozpahuRB508jpdm9LAx6LS8y0Ha/vlY/wUqKk4
JNqfMH4WJKCs1RUm+1tpkgZHfuV4FZFpmBGwydAIHA4BoAmRYDCzFSn1nByEEdHh
iqrPuW1Yt5tbv1KI3zvfVD4St5o/oGAU9WaK+hTtuzfneHF0B8t1zPECUSn5R5Pe
Hwtmh/I76WFpxBKZ2lISddDNobyExRGt5SD7uMK9OyHh9INiAQ9th5mpMk6jkGN5
20x6YyiRJ71zrO5bNEJntcpLvwa/vIV6D3plee5sQCEBoRfxFNupgB2lEY0/8Rc7
dZwBj7hmb9mkqfJJ1rfyvdKDk0FIRBT/0jaedzRdQEIjdxCzF2pFkQtWadRP6X70
lLO527NmSuqtTF6/zSMMcMebT+swv4W8pz2YEsUL+5yZ0Ca5D92Sz/V9B6sWl9ob
YQQfJI4goCE80GN7PJr2CWWNUPT8hquPlKymA4/pdtdMSvbex0iLKainO4LJhm3i
KK280rHATG2aXunPAEkvxcFMj+cxlTyjhDpepA7KVYdRCzQeCLdROSemkiUpdd4O
bdL7sutFDbky1SDbqvgbUU3dS5xTUeuPJtLB6KICcJyYTE9D9TrWJ70J1I6A6l8d
zU3TilJLxFDBpSjlcTUdA2ULmKt2t8KF9bF04NxRIqLwG5YSYOk5J5vuXrUNwm9T
+PkBZINgfHtcA8bJQ/c77wGDhKpedftTwhmBl2Qx1PXv4aeGfM1HeYSaVoGS5y8W
14npK4NHwdENNc9PjUzOAaz+JrZhyrzToQCX44PcwDUBgTnQz2kb6GI8XMzT0pcJ
61+W1YF2yQoeizhCVpC3R4xkVPN0oYXvh216xLGn7Hleu3cVd34N9G6E/m7u4DTs
8EDpwyovsaX1ZBHa97E3F1zXI83ALLyAySZgOXd36Yn1AZ/PryFeP5vun0PqGv+Y
vUlKG9CffXNqReVCguslrwv2u3pyIr4XVpPr94Em6XwFVN60U1DKdg1QHjikJ6bT
+kDp167HP040PljXfL4G+9E8ZIsnMAtm0wG9Aoh4zujKVG+HAFowSfszLMZ4P9BV
/874u1Jp8QF1d4hX21S38+7kUahc1LcjyDjdiyj72p3FZ1KCo5ok9QA+WRpXgYr0
VxFyhFWCEN+jgXC+oCPpTyKP8Bc5OVBXvT/ThJEbihXqhe2PH6GP9IKephFHkFkJ
uL4zdAnqIxvv3rOml6mtV/r/o1FScSBNO1EklacKVHLVctIB4i/jJ8tz3LgjP6wf
zf5sEIgrzzGoK/xaMNcp64D7bIGUo2mufAjOtJ2LksmD5WHotmWl6FRbiazZspD9
/yqAqFDoToJPFlZbW4om0KQ4xoi7nyfHNNUMpUf990LEH3lFzM+tad7PgOBfOod8
X/MScxSZ8oZI3/d1VbwpkxCQnz293UzidEMpIsW6M7x8LntLk3ovFD6ZKn5v2W/s
747rXQIAHtJh5x7QlBE+v4H+7hjrUiAjLQDqyrbOy1SKW3yo3W6ewsOpTbnz5n8o
WZ8OeddsRxEeMZHwmQVbbVQFk2MTw5BD68EvhMGeALoqcNsSM/hyQndruAk6riqf
CP7Aq/iYUj+KdQsQDRxU7HV2+EF56e5L/mkj7UdH9oJ4XJl2bSynTkT9PIhTKr15
ynWQlUrsvWVUwGxKyWr+nZd5hoCWOC9pgwgkcc1vZs7NqAGTNDfhSb9B1Q20uF+m
lUmggXwhRL9ODtOP4ComLBQQkre63kKuF9W823JwfljfB9yO06NfAz5ib+Ue/jdL
FvhNULcptMrYiIlvlAat5OrovKbmvOTMTq6zgqynCnBLP3uVAsLhjXe8I3Gsy1Ja
iuLxh/CA5oY9QCMkiF8Bhv1O0bhXmFJq2BuOSRvZYOEiMZPHJ8sjBKK0qMeiagDm
zczWwm4ABWl7Vq0P4mGF3tP+V40wP57bJTlfPwz9kDLoJADw4GCHrvT0X6DDaZe+
yDLfNliNCVCd4PV4vtVDKST96JQdci4f3DrCWgL3uMvYWjK+KluxyKyVG24zy9sC
pGU/rdvu8KwkNw52VxEaBQzPmtA5yVR6DGrQL9fc/uOuf2JmAYVQjLOVUE0hpaLr
7RdcbzVd/lHhOR3pA4q45vovOpZBULbLnI5q7A8myXUiUOYR5ymXjBrLHdADUvg6
aCSypS9ERqHvlUTKEIP7+3fxBoUOt4sqfe3VCtdU0kwwkeS5nUphkRbkF3ZqmK0M
hsrXWZKnCbKvxHF5y35Tk5YnlYQxT1XMOHntJhetNeoPeW8WnQv7l73KDeS0x63k
zs43+sXpjlUDnwcumXp+oInvQd5GTXd6ECQBx6BypCehrVnVcHxyy/uY4BX5xzek
urxrb+Ys9dDD2TUO+5sWFslP9SampmkxC2Ws93nlOKWDMJ9YcLqnU6c8A7NFXkTc
ZAQRP1AwIvLV+35daNsWZwIwRuMZhAyO58qtZzCXDAH1wX9ilrntf0rdfkDtFdC4
XbGc90KhWm1DWBU28FCWqkh+LZFbnKT77G9lbaItC6unwGGaSu0SB0xapuxrnOPw
YK7iRIeAyAwtyKzxTEQgAVzGdIsQ7+lb9B8FEVPzWe2Jtb+3ZfRk/74tnj0yyEfB
PI7Ct0kTzTUEYeqCgdM8c1APjE36m4Cp4nOHr+Kwr5cTkc6pYRjDOgsOj3vFW7lW
PgGuX7tDDddoy7HJtHnJKBI+17WX3kSoLRSBkjwayRnZ2DbNrAxKm70ZoWo4eUVi
B1qaYTk0G6SQnjBrTtQnV7jAGSSn3dcymaGuTv0nLJPdxWFm1plpKjzoTcZwdgtD
EPZ6xj6dxkCp1rjWrJ+p0VyQet0lwsB4OtchQRb1FRCQkIKgJioUM4YqBvFE7tew
hN/eDQZj3WOVeNHvgiRUOMpYo+X2m+63YPPQ348zUN/7torn36+L3Xl6fZ0eidtx
Ud62wzwnCWlvGHsy95F88vjM2/9aHsSS+Da47oRoH3kXgCxMuW+dfaGNnUydueVx
joEmnVCYcwfE1kDoe5UFvyCTCNY4rFSm7HOCkvxB/ny83HFp/R9U5zR7vMDcb7qC
fGg4yyUCywaKNZjDGUl1DJzlx4gygx80pFXjhKDDv77Z+HKX0+FUxoLb3WKbSfkC
3k7acSootkZiEGyDdGHYWr559FWkaHd+kwpJpyKa7uh7paOb6oNx2biMNWIxQC1Z
xQq23GVDdg/rZ3hAejQlpmvYW6mpSP1i7V4SlnNxuzqusLD1DQD181ypYxFHHDJX
WsullR5hcvmNhzK1e9QzWvwQDJloEFyiiV879aPglcTTm6OcCurS/6pBjwaIa87/
zelFWHfQuRGypWoK3Jdc71byWgNpZLl/w0RO9ri7B8+lBy4QfCpp8tD0PmtbV324
CMbLO6a1fDpL1LUNErL3zejtK86woU3wsoF3hn9FpWmnRZKWdqJ2WwDJr1DGZA0R
Hqb0aAPGIG6WipvpHArK84Zra7/HSFhgFZYNTSNBv9mEUxu1o8H+zuy7/MEY76F5
UpNu9BvAMzGcuA5/ol6dZOXpT6Ouv27l5h2sRwRMIBiJe0Q/HcdIoSKQGndvWWQ+
whhBoN+uCigfwUw9RUFeIljQSO2oC12wlTXVXdIP9vrZhVTE6D/6z9+hNP5gBnnc
KVzwRaQ6EL/dh7Rfq3oUS4M0KHzvyh41P9jVzIs0TVVSoRV7KXcMBBj4EG2O6911
C9JxlLlKgxyXIds0yfrcuItJ0bchpW5GtcgqnhaeKycLiL4J3jJzOqeTG3zN0WCh
XQtxw09ymIpfaSf3FwOhiE1pEdvkqRt3aWmpLClq5eXn8FJNrRaKtBZpAU/lOMrW
v+T5jztuHJWeb2xYM4vDqojutb4zN5CPFH+/WzXl+QnLPGQhwdXob/uMi3gzBR/+
fTpPvez7arx5X29Me08A9SHwWx6VXu/bUne9E/db46HW86m/HUZNu/7RURIQCxHQ
bVYNsIpiVeGJD+GRgQgnb9JWaCw1PJG2cDIp4lzXLw+IUarjOBCAmrwKD/PD4ulI
oj5u9abIfOpOFmDrR4eFON9R1s1QstOx/Smwi+BEO+fipRhw4NLZJtCJc9SLNpIZ
MUpnj561ZRiI4e7ZqCHUGUtYQUg4OTTVANGiDbiyRkDjHSBlwAl0XdqO1amfjoHL
IDyxXlsgupXF7K7q+l6lpJwaFVglXx96qMzOfoAkz8cTERFgcuPww7+c/rx98F+C
S2I0Gj+8MqEThdwf4Z1TjugKVNZTXmgB6lFyK92ZnzDDrV6wD4CsIeYfaQOINgzM
lhQbEdxknDAYbht8GyUi/6p4Jw0TxR5ZF+7kTnsnoJr7C0Z2xPNruY0oAL88ZrvC
ScmN8k82OoGx1u/GgZG3HqPjAZ3bvuW7yrZXziNcKmLSC6cIHiRSoOOTZPIdmwzB
tycLW5cvxZh5sRw/dpIUnH8AGAozCAfD2h0T8mwYDdIg7gR74KVZSdav19MXMI+s
C8feUXZv2oWl0OTFW/gvoRd6OW3IX27OmSqkkW60cSRnfrOYr3mHiOOotOvzTp3a
YmxVb8ly0RCyqV5fpU1NpIDjJoqYig6nP6cgoITfR13C5rC1F11sJtkmwcq8rKaI
xnuYZTqbYHFBH/U7MyffoXHqjI4w6sSCROrr60x6CJtMQhNU9RzMoOWd8nXc7Re1
++HAetXoDXVaq4YCo90b6Cbo5vv6wY1AwGfUCYHZGhp2LQNj1db4zHA8ohAZHw76
Ep/U5DdlrM6HRTBdxIJgzZB8TfDNkkizvs1g5qeOdrogl8Mrg/AIQ4rtUqlUg84S
f/wNFxp9ie2bv3GqMPJnrmVN+Si1kUBD4j2HRKQEBxoejZNGHnHSpj1vTguJ7WYz
9UROJIruZGfl5UYeX3DjQyz7lFf6Lm75Du88x7FZYe2wLq5yCJhn4/nhJMZmWyKS
8VH7M+YTK3S6WFhF0avFGyK24N0MfFow1bPTmXpxSSTgZgdd1UfuFabf4VkdU3bV
jXi4YpRtw9D8EyV/FRpvKZLteTnXGsnA7k/5udJZET9lzJNpgevMoVRERe1og8dD
Ph0XBbxtSHb7TQiUsagI29qBcr8QnCTEz6t1nvzACrtVdb08otCToUObZrQhdLcH
bOYNKll/Fml6h1OgCfU5esvubfOkULLsGn9530haXwuzJm/K5JX7QCJ6MDDUb6N2
0UmVvijuxog4PoPZEEKdh1/2nNdceVyzT6yEfRP+EQSZGDhJsiL+5zWNMNAcG6WF
tRCkG5ElWxAYgTKY1+NIlJ2Fwxo+mAr5LSi12fggyahzh2nQnIIa51ioj27TMdAD
3Raf+ADlDzicyGflNKmXY8u8DKf8+jstPiCc1SKTZKo6r79IbmsNpoEYTI/E4x/a
zgbZTnb6QqSwW8BjWpeF3B3PTC/K5dQIlyfTeY/9PIWslZXWVGUDy84vOgWgGaCX
k4bXnKe4Mq1xeVSIypDI8vnNjm0xBhxbf7DPZOcnjjOslC6t1T6pTmjTUFnFNeLA
p9lGQq+cb1ejOU1MNjcTtn+YePMgVKZ00NUyNqMVkTxPbMNVN+XkFTRUvQE7XxG/
Zhoy7w1HzULHpnyM0PH5nDt69Ph0MvuccG3ybyJ0k3ngYIA8RXMQ3Nq91dmVc8M6
OeU2Skbi0ItR4pvih8Ljwaa3EPXznqvSEf2I7d5B2gZt8rbUGzl1G+QdN5f13GSo
gNwiwupabGlr1ZsOEjsaAAxbLXVafjhikPIdbU2LoUJjpMAO12NnnF+EZJ9oBu4S
g4vF+aMgzudcWVF9FmyqnGnA1JJRHs59IhMbJSt9+5L1Ol/EzkEwYNBrCveTD8WO
ZVMKs3s1AFjqHqsZ34eUeNbtjxwEfwDREye4w2/1dIZekLUtvhgu2UuK7NA/hjuL
5YSq0X2+5/Y+eIl8e828gzoC4eG6WH35UohbtkEcYg6gdWAA9djUDxijAjpK5li3
OQ9nqipuAwkOhCE375lcZNsIhUQoAgVsR71753LcFy6qngymgaJhpopW36N60USR
hw0J6a60gkhvlX9Z7md8hQbM7vNuUWbrwHKTzvLoUR4TWiKKZ1ZIzNWcfZa0FWUA
lon/lPKa7Bi3ri7G+eyhWbB5cwrepDv0etLEhNp5n+pSc90CbLyJ5/0PNYkNxn5E
53FF4ohRxgBKGwT4gcjedg1w79TbrC5anOnVjNoGb0+z24mi0OA8C/JxMeoFxvEx
WAs18OTlbOE61Kg6PeLAPQb197xDoNXK1sf5PPtbiChQ7CBHX2iGyte5DP+TkWob
a0Js9zFGwsKc9LKfC3PO6+j8NuxMlGeYKSq5rSnWsNadb8aYxKTey0twgzXAi7De
ZJ0B03uz/XfpfCGJPFA6UkPsFUczXnhywGa86DdWPSuvY1HeEEYSDDy3A+Tj/LQt
Jo7iEgK7yD2wpvHjX04qf6eiBZu7N7O+wSZxrAvYLHcb2bYqsSXuyoqyNIqsUejN
m8XAkGFBLae/WWOobQynng+H/nWh/wr3ZxVtVub6yaj8w0BsLq4ytsm73Lz1vl6d
PRIp3aOn5PxvnGulubueQdGckXEsAf4z9+55doMEtt0ZPpF1ekf5FbeA4XBX1TOf
Rs0qRxNnFbDhYTyY1wBxgy7Qmk8M1cOJVol8BjzZh+/j4ws8dJY/mU0RWe2NnJJG
C1m380E9JU09MsnznYLljIfiA6GNmYENgu9Ejw5O6RMb/fc2Uq5QaFzecE+WtVAf
Z8TK9hnxbmFXmz/VEDQT7Mg4DiAwsDfh4TA2UG76KPNLa97J6tJN/PG905q0GaAy
isovysoy3Q0TEOS77aLPUHAPjsdqACjPsVVdPGKH14x4lzU/5M3kczod7krGyiQq
jwxwGZZwC8rJXAETjxvG7MNzraSwpja662AEpFfgTlcVS6eiIU7oOchj1o0OZHEd
Zy/UZzJMeTY+cQkCp1j0DvO8foMmjG6gWTUwTt/C/TOMfooanYiYV/qPGJSVmDeQ
/s8b/lXGhMEiTj6wMJ0FWMQdBXhQxphCIser4OcORkPloFTvfA0tJ/gOq5S5kzzh
Sjujw3SX8387043zfv+DwWAz79P16r9lnEFar3gcWxzPr5mRzLX0lu1+/Fi8g/R/
xdavoxxMzMWUA6bIiLW8cXojYHg9rlQdNg0Qzv1HXb3zPswYK7trgzOaV6gHdDno
vsU8dIVwN+69/OLvj5/Fi53XHugnvUPZMNmXeQmSo4ntfFFZPlmEwrZ2Jpqqjmo9
eL6IXrtZr1tQMYkZ1WTgDHshve/FdlFrZKUXU0VB9EBHOHAU/extXKOzsdzOgsWx
idcBFnL+sKuc+VFKbBtQF9NlxKB9bz+pkdqp4MVMwqK0wZvAA15rz4dsAn7kDbH5
gyBTL/RlskfAQaNg+j2346JZJ4IjZmltrlEIdtj4I1nh6ba8hYPCvtoiAGr5Vrv7
RnTMtax0EsBeAiS75iLvukIPl3X7NKb2AkYRnzdUGTmGChzIE2ul8GVZPTdMz1Yx
R0fezdsOZQZ2kHFolOgkL985e8xb1skYC1RUjVwZTS6/RizLYaXYhi1izHhHZrQu
TwZbN5lN4483wBlwdvxtmMIItzVMNicVM4GDMapNpJ2Zh16bjlGADPThxDX7gYO/
JlDpVbK3Fn54menqGdHP8lRFppkWtmNrK1SZdm4g7vJJMQENOTJPN+Pa7Jb0226w
OF4XeT01fQCcDdXiHWvmGHQ+YuOtwGnm4HZ1XD3PyijX01QK/GCSdKIPE00jAHCM
KG0+kURvV6Je2yUduq6T6u9dFT1kkSd3tsSnKkTTwibnnzG/sY7gmVu4klakTKuP
by/orV1Bo4xoGs/uOnO/kzDwbsY49O2z1niQI8xux8KZYtclBsyFSeJ+gfL6xP4n
VUY8gfblDfFHSeQwR2Qc8qCRK8rHgkvrqb5Z64eAlqHMoLH0g/I9LWwxxFpzbroH
rA05XkKhNppNQSnSmQTgskkty2qWMUmJ6lGleWVhB/cU9imqhpyKeEzf83B2dfJH
EbgnHxoEDuHKfrAc9jVTRyzdFs6j6cRdZs2sQZ/vmSjPxPRKFbuQg2M9LQnR/jpi
lB1q7yivkAAP59SJew7RKNZypMQypJyZS91p8Pn2m7VUZFpFf0HQHCzzmfCTylhE
bE9zuSOAgseShrVBR349Zuq9OTsps7E8+2AJTB1A7WlPjCEbsv1rh4nQnHbc0Axz
Gy6IGF0ZgDERSX9z/5tPV7/YkgsUhx433NrMPuSZ1Doq6KaE31DITZxs/P2rWaLl
W3/bsl/gue52Qoxdxs8unkgA9Ctrw/eEAlxjm4BM1BiW5Xd60qpIvuajzhguqgl/
qnro2IKu1TGBbdhmTcyVpxZkEY9bfAKkG8d1d7ATDwI4B9zuCTxOxEkmwqHGWXD8
mf+tl9UbGiF4bbBWoOSAItWDCY8Vlz2tI3lv9/tpwZOl8zSxlbmtDRLjjfy/wxR6
bkv3CSYQLzDTCXk1qUTpIwFIOC31FqjbBYwZq5/J1ZmTTdOe0a6XDU+xt/VRN79N
AvYjVuIbTLFZItDc8lN6xm6dc9CJ+phn6vjplk87NTYebQM+ZGHS05ARlp12hJ1T
LYB4J3p19mybBZHEWoZJn64R8wL9nf+aKBFr/M/BejkIpHPz/KnJ8atYfCy7ELJb
M8Wh7ECPj/cBCHdCvRa8myjgDBohRy1zj88mvbulJiJ44FTWYS56fFPsnq70C2Yx
IHowtiIVEsHPu+sNwZHa9cpEmjrjFqmkaoDUwYMytsONidDQ36b/nPN3OiAaHG54
fbGxtuQTpBbmraT3qsK/U3hjRHp3Hf97tn3JstaDjz5V4YSa1c9bUqpNmFVnZu61
wJ7S3JXzXN46UeUzQvTjBTSEfEg4E8VI3K8thUzOQ2Yd8g4Vgruf2nu5W1/FidC6
aYTbmd7TtD7GSVFS0RFUJPYCocJq45DSSNL68QR+Y9UalN8mMNKjI8K/dh6ebbwP
qvuPGnCQ6mL90bm4y/cBg4Kwtonzhe2HTPmiNLNmw3WnvGIy1nuAISE+WbvTQoYg
Xb238lHxLt5+amz5NN4CnYumfNEmiSr3itZK9R5TVdzq7QOTUMm/xbIFaDTKD+98
rvpYhaFu+m5P7OBrHA2zHO+a2FPlf5WKWnZcI1V/7z/wXDW/ofhYAyxB1vIgGAz9
+f79Q17hFeXmhn6qGkrx9eDGqW941qao0NaK782Vkv2C2Iq5UElQ9DO/pluNbMG7
I9Hb3Q1dASlt9wqVQEJjj+lLvfKzgA8khwAq9zfhXEd3wdD/rQC/Bg92xDv+qMjG
k5665FuR6v4+fChm9i9lW0vcfIwg5Cvadl043rpXFUiIBZztTyB0ki0VJpFDpLtT
DxT/KcYDFW5QnuVPA6lhcWGC5AvxTxrwl0C+o6T8IpRW1c8rXJB2/RHXTdUFYE5J
fys+w9z0Ak8D2JwK5cSJdrfgaud6nmuRTK4dqKZojNF47iPd3WPf7rCBzANsisJ9
l1L67fiM2GV/pzmYvnT4/fDOIKLL23zuKqkU2qupeto9G0f5tw4Cu9nRefdUju/9
ldKhNWWv8khdjdVUqPQhdSNB2e5liXF/W0GrZX88aRd+kNB+NUKkPCVLCcXl1OIp
Q2I5k+BrZ3v/WAkZeW6oedysRas7n898eq/eBz0XROnz3hrTE66jfGRrBe5yEf7Z
Mv6WIADXwdXXHKcyOHIatRWhDi+gq+ovWvKS9ckhVqbK8md+/3pYSXUFWcbj/NPR
DBl3pFTGLvgINTkF9WmJbiPx2vqVhNKNWQ7ymr2EhJWLUuuQNDyfQT7+dnGW9/61
CfEJOltFXKYezRKoe/ks/hvI5XSDwqA/sqyLgJRpBkiUKUvPXrSBcW9JCl7IBXf3
B6/5jPRW9s4vKI16rcpVSOtBpxz/mAoHCT8Ya/dWr48aQfHw/ZJIlcPuWZ2VrtmN
0ELIWMweHtw4BoYGnyxS7XAy9CpQfbueNuhKmjkzeTF/lB6TudDe75sL27e5rbHC
dTw+gT3e4ijobw4GuynH5JiknMbdO3M+g6FhuSPObNiylBDHyyEr+XCOEXG/Sg/S
JtfRxF4/O3GaEyic9ZqUFJwLi5Ca1Ncpg4uFwWKCgb/ufEFKr1muzKWP/iy1zoeS
YCxYhGQUC1LefFpW03ixa0nDQOi7EOYLNXmd9fDzgHmZnvrge21yqF77Y6VrX6V0
lZBTPHSO5xYQccurk6cN7EhJjHw3u5FMrcPAyLh00SX3IJ/x7pVPiR6xn/x8LPdU
IcnFJ1XiTfy71kb7TOgjMdatb208tvou+LcGRqDFW9yr8fh85IGPlbrkGZSKnPXc
oqYz/4VM1XbC+H8jgbqHK7ct/uqsmyWEMPSW0J6QXiWbvP6uoY7PTqpF+b6gXvzD
znNCrqKtk5n3IH0MCwmW0nwBCREUVCgwZbcAKpM/GObV7WDZHNAVezj5pXURJdo1
xoHyylvifwFn9/xFl70gOhrS6phQMQfOmoz397UAi89z0hKR854+baYuquJOS5C9
g66XR3yMW+GnzMkTS0CZ0j+naXo05Y94Wv8U9a8lVzwRY57c2sN2AvBEtUlTxido
e1o+17KNgDn1qYlFxK9TJW40iC1maeWVWgDyMp7iMi7caFR72X3NBhY3+X2vApYq
a1aMs8qflk8q11Ujwp5w9ZuqL9mX+8M42uPb8/h5s+Plv5O8z131wqUMD6EBfjji
gAAMkDx/eqa029TQuk7MgXA15b/C+gepm907WZfQF5ec/pA4GF3NEW8q7mjplaZf
y7ZziHKqK35ODeJb5J9jnnLSliILVB5qFjXDEHKgRFBU0Ts7f0HXgODDZZhfY0P+
6WX1ccbY4oY4r2m3TuQ/vCmhoHgWXKCbG+bMkPwvK9cLMnKCuh0pP5Wf74ENnByY
01YN005yk+sKFgFVTnmmPKQ6WbuPfGM00U02uvzsI5kyNzX7WrU/sAy5dhFTTDTU
HcumjtVi/4dL+ucBTP2aEk0DvRdjXszukQUToX+/Xa4eSNWLk0NWrmdTghYZOTh8
N7r5Du9o94ZYlPzZCC8TBdOJFhvt6++E8WO02uPnWi3TPvdCkLF3mf1E9rq4f3Rc
S6LnaHfRdl9gJDOdt+fnI0J67Zbyykixj+hGseoofLVyugVk1846i2JfctgkC7tE
XLhgCQtvdKmk0WHEpaTl/3nN1XS0smlyqxfY22kxbsmwoXDTAIogBULVIKbSE0wB
O0Pi67oN8YFQoehe9K7otzkxYaYgjGCdaStnKjENA6O2tGXVedvEmMo4j9G18S0Q
G5/C98JScOZVyBTutBrlLpLnWAqwf+y9Wi51s4WGUBq40nrKB2KZz61t60gQdlPz
pTYFNhSNF5uSZh0ZKsyDlcXqTj9mZLc3AzUnsDzMaKTooRaLwL+qXYPUTBxNx1d3
nprSGMq5BS7jwqtsvZProYH/no4PpTIVRsSrbRGbXdPt/IyCWco1EzsZGHfiLnle
HYTJxKpl7EZ7Xepl6MO2NYu/vnDYSb75a1Nais6jDmx1+uHA8vNM1qK51aOlXY2a
BJCPMsVP3hnRpKth2ezJUS3//c3+GvXRcrqf4+A9z8196QdMxrZ/CUul8OsWEs6j
oFSoyqDAvGRlUK2weVoyOFN6wgsrPn82nTHMYc47HkMfSGAh/VcwNBU91/AL9tsS
jae06yie7IOXRMyo9xbrWPLh+j298kXNTkJ7vT6C7tZIVxbMQinkZ1w3KekBqlcl
FCkQEmUsKgxALWmBVm6Q26UfK1EmpRujKIq1ffZMgBHCx1kut+d7NKMd2woYTrj5
T7z0WFh8SqhoYZNws2kHch3M4ptfbosjsBwmeFj2I9sI1FX6ZcQYqorGsPe8e/f0
1VB78Kijlhg7vjNTkEzjFcDUNDrAIvI0OAmiuPeE0UWEV/OthhArChUjtWbBYQ+u
RUEnjkFB24AsoQ3SNJrevasokYEgzikDFGmrxs5jNg57o9CkllSyLNZrzesd3D+/
HO6/3IhLkX13zioE9DG9hS7IEs+ePwUC7HjtFfoa1jOeThVf9L+xGYqkZTQ6muUG
nRI9Jr1eDuGPTvE326Qd69Alb48BttnuH/Xdi1XyTlFPeyCPb7W+DfrqD9w/UFFO
dmcfJDrWx3XYZHlcpTreAzJbKt9XraZLo6frBAmtKzvHtuzEQVsKvwRJkryWqQfV
tb1URekzTFPI5KRIPbFv8mVTywQyYbR2wh3H89tJ2ZmzMnMzwx8PXB/qsFQZrtOf
UJMzTNVhqr3N3n8GhmMQOVH7GiEGCMCuqcZMzCw3M7lfg6aHpDUhy6g15R2sn728
uD0TstaoTpB8ZEL4tNaDymCqUO3LPG80XYN94eY0W1t2IIpK46gDU/DE3/Xueqqw
QiqIrNlaLIa21opbuE5f7MKu0stnltobR5dI6JeabXHFmkgb8Pg4WvCu3E/Z6bE0
mzE0mwwexvs//cp0i8H8EZddEQSbsSjZ7L7vBR9sRy9cwXSRRML64DGya6ApUmsz
GXMSFipzPwwyRRlBvSvz6tsVeXIDvQXQS/O9WgfWTxELtFQGJ86H+FEMqOxBV3O/
vV4S3H/IgTTjAdf6fDq6DaOqI2YJYrID2FpWPu/T9mMs+2pd134mdynTimqkPsJl
DTk9CledTBVJvFmyuPE5D2mCKRh6VTBllwlNujDFg1ZIh7N5ZSIjsLdAvm6lY9vL
SwvgJB85lb8zfX8RfAJHftbuHB1rzzM4mEPbZ5XIU2qB4NoXE/F3N9GuWsaPf+BH
L+99kHUz1ce4zxlvw3/J2Eylg22L+w9beDNxtXGbziC75TH0x0VrZVkmV9bilNjJ
QY2OYBxpXka4FK910FShqyHy7dmvnlQu17OT9NY1ML6o6Z2SgGfuS8AFXE4Acb30
S3w22wH7dpdxkdVbGBu4Eo6H1hkZzzwqCPB8i8FYbOg2MzB8oFdrk71NrUtd0DCL
fArn5lEClaMEPrnp4KCclA3fKMJhrwj3ZYwYZdAH1pfLRytv9tdsNVOFAs7c2eth
M/7hP9trK33VpWWkaGnkAlHctZAP1AAd78VUPnpexZBc/wnoIkEwZc8Z8N8F8ejV
uki98JWAReqft7rhE0cDHgQFsLqwIJz1GMRGc+PgctKNQEuNgM0cw9oUgeAH8gFi
btKuCIZ7HZRrLgQ6h8lOJzmmMzDu7MJc/Fq7WYbCtPb26Q15NcYETh4dINI2n8OD
gKZ0Ines8NN9rpchpesu/rcZe0Vdh4J5y5aXNtgTwoPNxuAsZuppjS5SwP+/qGox
uk5dIGAYCnEC7thSt4sgHyYls1lV/VWcanq88Iy8sqBHcCrQ56tzq90K+sWzPxev
3lxWKBpfa2lwvUaipxkdM1diGiw2Y1ecvpKZOptXP04bmwuuCECBqqWzOqQLR6vj
2lxiNqdMa6xfaw4Q3lPhFK8OxxxKy5tdaOtuqYpZZ5zxotTvE4gv4yFLlhscaqXL
GBg+KPy4w36ygtE0tQlvP0jk3s1gQBHKCdtFnagYO5FJILHGD63NE6uz00u8YOpC
mVEjDBYdym+jpdt1pr4POeHm1ffVaDfKs0JN0qDO6XfusOcm88zIcIReo/o/GFw8
EZXz+zXGxh+p9ZNpmhjAJa+M5RbIbA6WEUiaF4ZviUOR3k8LqxfJKJR5v9bNPDta
qzkAOqhgsV8get8KiR/5Yx9kOLcH/QF0rpTTpWixvy74Rd3u3hgntM8I0HujN3i5
Ozw9EYNRPM3nsfEgqDDTXQoC2rO4rIXKxpPZnFWYz0fXIRNF5U+DTVW/vnDlLRvZ
QZ/Xiz9qU7e/+pq1Eus8x3Rh1ePVDsYLvfaqF20+jORDw1RPF1ihE0d/yYp/ZCGN
hhAPbzdd8HMPTEsG98MbEXCbz6ujjnmlDy//vipiukm8WtKlcVUhnUQmfMuIutK9
TfJ0p7kciOSRsL0o1p/UseUWr5od2TsaHUMvbsmmS3mmrCI1UtRQWkJBwsNTN6Fy
eNO20AU8OgYFUPXw2L/E0uBsoTqguHC09RZGTp4OLZn87GZMkpB0Mo7BKZxS26TR
2eb4vlNSPb+to0tm/hO/Tt3OuLNw15Ae/TC+U4NZtU5U4WSr6JF/leZRFeOUxsBL
Nm5Vt5rR54IOk1J3Syvovml10eb4a8gnNK+dqrHPcnlENUdEvj6/hXNnvFJueG+w
8iKt1VU6aHk4oGSzX2nTn8KekwTWB66U5aOyCEnBrPNxSyAMIzjLZMLBJ2xlRPT9
LU0vdSOnvVj6OnpcUXHnCME0lm1WfO4CUK39QIe2f4eS9aAZt50hd6lmbgGpRp+i
Vow3EDf6tpqUWqjqssfUk0ciOaAe1/bq9i0MfP0G3yuJY9OWEVzUUYSclWW9NCPA
Q+l8f9kK8TbMh7F27UGU/uK8QQK5/Qcr8cvEvBFr209l6lb95AG7VIcAwdsALT1u
Y71EhqgY2Q7JYpjHpixHpGwNxYicak3WEV0swUX+rF6ygQ3KvWwezgolB0MPfHRy
JwUfAdiXoVdjR3d9cIEIjibBc39xfV6hjUM8wtkFB+olu0I4mr5/G4gwdeaukjaH
7XyLoFZVCKqMz7pY5V/oLNOLGRteLZ6JA5SMeUu6Ncsu2bp/qEOH01Qyr6jHcrJ7
qvFnHNPdZuNGwEgBaWjxl09qgRYsoC2hEvxdOYfzuuKROetXQRyQkeo3kfO8VROH
Pemc1N8YxKiScJECk75vikVbRVDijUG/73I3i5vWchepM2pXa6Jd3YoOKOzJQv56
O4hMJTCX9c4xrsemwzmcWNZfqW8CIzXsf1Ajq075vyvL3bDyttA4digsZ8Ak0qij
R9d7shVeIO0wN8pzOvXv8iSsmIxZ4qiDfKlX/GCxtIx8zmDgVP+gxI0AV47N6Dq8
WS9lAu8ypYlMB+7D2bM3bvNUfmlp/nttSoZB0vFeJqB6RTextU5XJW9h47XxvIw0
/hq4kaDdcnnsr0h9s3XLNJbbXr8/ZERF0DBbvDGZ5cWb4CLjpXX52tUYlFfBjNkF
F87Y6Y6NI1jn8Agic84MW+WIIJaVhIaqQp8R8SFC4+jLozJwUWxbCu9w+O5aHQKb
t3CKMTvynK2G3VXxJMnnxJ8bH5yVIf3lywaRM+8jbvUHXd9iEzmiYvE6lHwvH6LF
DJI46gi5T22QQyRijhH4p6AkcFa/BdBkob7uPoT47uMHqw3Bso7GDIX7cK8dZmL6
e50hMs7WXy6gtpd8IQor6q5/4rI08KNtlq0JHAt2dxoR1drb0Yv6p8wGZzHOnFxx
lS17ov8TGZ/MP7MDg03jFKz5Aptt/i7XDzSMltDpLBN1DwGAO0PeuwdRufDfwJRL
EpvJ0Ez2vJeIK2RcZc8t/WAem2a5AG+ZL6Fnc1+/doKc2sYZO2YD3Yin/TPbyKdc
t6ZN183tKT0q7ZmKpvLngEh0Xo2EaSOVthB1Dee5icgsCzLxv4LxxSMQHryKsacD
FacmMkzoqgSX6rxcLdlDPqKIEaSt6TeoAuShtD9U3FGsc16XzWYRXZXIXOlEKcHj
iS+1MC8+y0AoXejKqkXYU/BfRwV27eITloQhexRKSqhEU3u67pvNy6d1bxUvBU3F
WFJJzD8k7VjGrSTA4nQ26HozSEag3Dkk0kCS3YLYcFrRaLRi6LQOuTteC8yCHlrl
jwcm5k3VX2S52ZE1ezihE1RrdexxmiloIKWQ9W70l9Y34JYW16xp10k2sSe1oZuP
ncV3WNHZtQTjvVw2SuMMxIT1yYxImW9BiJj8U9iBTCnCI3D1wgQmOMmDhlwLV7za
CI8GcCeLNss3nZJcpVJHspm1L0RQ+yM9yf1RojlTuxDtvRNcMC2QE32wNdYBQFDG
Lphi0P/igC52gi9KrvLDLfp/Sa9au+EctGneXKKXfQUeP8dgL2YRk5ArFWTDwxWU
WERee4iAxweNtAuKn/mfLj40aflvTkjz0M+9iHfZ1Tov7AR3mFPJMOiGA1vI2qeQ
FyMg9ENBAgkxIIIJ4vxu8otqg52Z5q5CUpzPltiEPzHOsgc1Nq6WpwRMfbw2FpBI
+gGn2WCMqHT8bdejfVQbCNtfM1FAIBFKpZafNa8Z7KMy8zLTQ7dEYzsA+g2svTWl
qIw7IFik7aRDV+sP7qMH4tV0s/U8jPX39a7Z6YHiH7I/YZlEu5OI3cu7OHBNxuw8
FM9DsIQlwzeQRskWAUDSYiQiIJynrcg9xwlQ5P55Kt9YnFKYVVWeaLXUXLGTumem
Xb3AYF+NxwmAyGiQrHbfFyEVAnrwk/JEh8iTo5Oh6CXyDparkafflLZW7gIkhPKT
5TCfn57nXMMuG0709k19+oftazEkrNlelNd103QGyV+dPr7CnZATBae15Dw+bgyc
qpxu/e9bv5DkhZEHTfSwFgvvAu3M2VzwmBj4B15STOo8H57F1SGvsghaf/I/ugjd
9zOyLnW+D8fCxZgpxfceQpa8SGDauaaxnofkPdbjpwJFkdM+DiFiWS3Knw5Y56Vt
wwmdHGcx1faBOZnYbkBj1vM3d796rr2ZtaT6fzyjJc49kRBqJcMJIXA/se8UiwQN
ygNqt6yg+XBLccRItWW9abI/MMJsezOhUxkzaT1Nps1wYTs07WEuPa7Wt1fAf9Tn
OMmUK2uN2JZYRWB0gClNLsldRKROGJiofBg1+jDFouUTqe/81Hl2Gif55PL9c+CY
KSsGw3G21BiCnWNfU53tSWPP1XhwLoQSBrNMh1Jcv4D3q3pXHw3lfyztHRaS/GIp
wD2eTSF030YEx3/NTQfQrTVGyQmCI/mCivRTOAsO1QPsHkb1CQAxuTsLGNPU2qEj
xxi0wpO6gkAtha17ij/2ceI3yIXBovs2BmjnKIftzQA4IeA8BdzYa0MrWxYhNf2W
J+MnDfi/CYPPKe1TegLvduRBdv1OKYqTcYg8vCroXn5F+0Szw7OmuzSxfq+hDFFP
F/Vybl0vsYkQSMYZKSFqKtrbOBjs/2SoSKvIM7baAmffFZE8ajaHeoRwyEpw6SAG
ADGT2KUTOPPjgOVycyoQx8PCm2YPeItlYJNgVJ6IVk4vM0GJeHIiAEo6SUK++bJC
qU1yvZBQvMmnxAIUmumLZEjhntWWVoSiwvppnVDGTqqo5Qba/EBr0zjcT3z8LqyK
Gb0lKkTdZziuxMNSvqjezY0O67V/I6cv0ThVzthbTqdg1F0v0/LEJZLAWp0sumhR
0H7ygp/HlkURs8paYqXl5W0IWmwixTlYrPPG+jFDDDEX1Y4hL5e8DDfi1wUo4Jhl
nGoPhWQ3xq/51A0s5rjM1Gj5rVk/WJMQFW9n8Msn+SF6O29BgEFjMnowQ+icMqxI
jTSDKA9gIaAGEq3gWA3BEhbh23CmXgeG74LRK+YIS+pD6G2PT97F3dmIlTcE/EsO
lt+RJguWsOTrU7ns0QgbGVCugLQaUayHI5LRpMViHUp3hZlww+6IrelpdLiSFApX
A6KNEo4crKl9QBI9XZMoeirv7z3HI6cG3BGNLEIAs6ywGMH9QAtUo+QFJZCg7Z0U
HSmVrOE/wm3WMug9lplAMIdbkJesYQQZphlRDnK8G5T0W2nsrUUTHiHktELVMbNM
wWysSxjRws26kOMH7pHifTi0qnnI7InvxDS3CllXvvRNfgSlosTjWp0ctxEAKN7b
KYnHp3UrjZvylpBcAdi36IhQkwGVU1cNHGDe5lQ0A6FRYF/1tmNcv+iHGxv3M+mx
IwFxTIEkF12FE8a/qRvm4FgBIoXcBEEicX/cxsLcRBqCIzsajm1AIzbttdf+++MZ
EYe1aG9bcOUT3zw/R4+7rO6rQP4u2+MQLEwpClqyKtXO3sFLhfGsJnmFI2yTzBYL
ax/cIiuByCYOGOxfaFXsNqB1TvASmqMfZ5lzjXwLZ4Gu6eMKsKZc8FnfNoN9T5Wi
R/zOcru7XhN9sBxeAA/3tyn3m3JsLOdbYhl8nyThEGIdySzE3/wWXh13PJHTEyO8
6PuO0QFa3F8ECFmEh56Ebr68/SzPcwzRl6XB1ftQ5w5mxf5VKAvDSwSFQiSlPsTU
qCrBza0abkUaN+t2Up45IVT8hkn2+pHVLxk9tGXqRabFvZv5GIn3N9Ul5efuBOs0
LpBJooekyPOWX6cQC8Vv1lPqleUA0ohVZdGd83P5rJIl+uoy4BordlbdxJubjCE3
yl//ep1tgiRRAcS9CtOijZCOOXoRbKaQWQyYUSY9ZiSWgUf0xffb9+tohGjd08IW
1mXJT9GZoUFuU1vpD67NWTspfbfAUp4AZXJnCP/cRMm55hsVfKjVRBGFvlm9dtTK
KiJm1X/AAA9aF9xRGcL9MPLsf2YBSrsCOKW9BUz7S6v9mP0R23DUSOl3lmGIBdWO
0J3/JbZRu1ZqgRCd3LIpXcciWeSmg4f70uvxeYx12cpU8v9mM9KMobyT9D9RrS0j
3tGnsBRePgW6LtRZ0cqX6PPcTtiVYRqMW1HpLTZO48jnt67rLF4E7Gxx3BVP6Km/
X9TXIutrpdPqB68osyVHWi0yMmaypRnU/K6O2avn+TyHVbdUM+lJxQuriLWxtZlg
0cx6xugTCKZFqKsDbCNBx93UNQzXnAu1XiMBYUQfUeY0WB6M2lwxV4v6YOiLJ3U0
Avqf1Bs0YE4w7nQewjM60ZZYI0aMG11fko0Pn2NSGzpQWsS1IopurbEhxcFLDcak
3lKkAdZzvT/mUANf+OVW8PVa7v9REIoQ0phX01v7EYWHMSAyRZ3c3byY4swRyJmu
9k7ArSeM3W6mQ9/bud2XFv+ApjsbMMVtL9RizBseR01ngBnFv/WUPiVGTYA+0qC4
UErk8zNu2KIydv4aX1bdRJ4Y/lVvmY8TwVnSWjn7UvWzSz0izPp3Cux3TBTNC2Xh
LCWE/sibwvClZnW+OuUwe4ekkZyqaQazRknbZH9QMqVKrlEJ8sLq8dp2jb1mYZN+
W98WhSM7V+CHMJo6lPlt82pQ3Ixqq/b4H81t7N5d/r923ynQsSbmNXbDxBwb6M//
8GYZO6BWw4QupdZmHbfxwWL4Jvypkr19qs8HcZT3CwuymqbZ/+ZpPGWjV/iS5eTW
4BKv+PkAnNF6wPyd23h7H7wE/w2nXqnBZoliPwPHxt7zSqEuUm4NXKiJ1uTF6bTB
7wkY1/4sSRboQhIXJxoG/KKRH3ZRsJlW4u9cupPwEelu4v3KUSasS0wpAHMRSheU
fdB9u1XSRUmIvOwr2pYTgkZ+5nX7fq0zw5yAGuGlBZKCqiozQ8mPjT1CrlapK0KJ
WBsDTIJUPPlfr2W7ymc6F/XZQ9nxI1hB7sCydVet+BGcw78Ga51QXSDVHsjLmnd4
9N2L9Kuc8LuGC6ZiT/5uxs7AkxMa1xlQVcy5ciOs8en5hE3ybefSFgirqN4GPhrg
+xmC8F9kH8ngTxU8qmYtcJNMNsdp6Q4EJfi+AIYe50WvQTxtAcDjm2scqb36fC2o
NwItZ0ZfgGsmPDH2UUmOiw==
`pragma protect end_protected
