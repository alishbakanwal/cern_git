// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 14:01:23 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
r+Jiym12SlO7lmRPwmIbkcgLWHDzfw21Mv19HPuQ0nTSnJbZfK+ZoYGZysMgs+Uq
ljdp83e/x3sG+4I8PRIAkMXO00WVgG3q/DvnDa/SqfF+BiuaI+7IloFzjv08BtVq
WWGAciNry1RDhkUWlqqRcLuIfCKFS1H0NNCPOELxXZs=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 36528)
DlB9FwoicM0fJZKaCKrJbg0OEMrBnmUF0gvBQ14A8QfeRsKtcLpXun+ux/mfNfUr
NAeuQqh4rkBZu+PRQ+RtI847QtRqC9sfthNg+kUHIO0HlpKM0rudqT+t2O7MYF7K
2MKoLnvXxPf/bkYdzEo3zw30msgJ4B4VNlbt6JgbcXh6jUUy50POGXOsXyjv16pr
DARLBn499Q2ymHVLyVgcSjkG1LyyweMCKUDBp406yFXfgdNrizFh4KPrqb7XIPLq
np5ApF0qQlmxdXHE41/qIeM92eK9MxUzsg6aI5RzWX2syy0SC3SAW+hXFNQTzjKK
SrEhJ/0qRvDCyMROsiRtv+KvwG73drN+EvFPyGMDUZH4Hb5E2u+a5x42GnSPz7HF
D890kfLQBhKjFMpU+1gtJZODmcKibvNMOIEmLxKH9ne2T0h3z24avmTZEIcMHHP9
9fwz8Eom3rUHTR6aMXb+qhztp8oONUk9NuUnRwVDdAB12MgQIVbXSjJwc6blOMA1
sSmokykVESTYZsQdAtMEjzWX58R6PswSkijGEzxTPAs4g6lM3mTFZQM3lknXTNBI
TdioWyMCvt4ziaASil9DFG2yohlwFdsg9h4s08f6fDHD1vXUpEC6Ism5Q2tUQ+UK
MqRMxDvH9A6Wfn5FQZxvT4Ip362V7SfOvDYXBoAT9fhR/IrLVl8NSo6DlGO+i8In
Ekm20fzPu8ailkfneVlz2Otngf9AiGcgag0cirXfBPN59Y8wsobyNTQTnhp12NkU
tVdRY1Bz2vbU6xmNfhxizqtYlCFB8T8wcjy+p0/d2FNcxvE0atNEc+97EX+MCsUF
GoZXb/dRQHNUQS+FKXBDloYeWv4eQpVXKFGtKlDM3mQz8YWB/3exnXOiMHhG21cX
j1+7CZK5jz/uKZEJsnKyXo0ZaDGMg0Z++I8+zCAs39LQ3gDFQHu4dE0sUb3jsYnl
fEiu6zYA6YK1gi3EddL5PsORDthoql0B+J9X2hWZ3xapSYPjmuqqv6l/BHnikBiW
tnfRT4Y3XuZ/txJRsuU+mBbYC4vrTg5C09gQwFFLa79w3kZdDOVruV2hyuhZvK4f
41drCPxxllw4dqhUhUZQHW+E7iIKQDyv78GVRM1XR2uR3oCly2zWv2+LRryA8pzG
QU7GKQDek73uIkeHfy5gOFu9NbznlgU0qWwkCWaE5gixYp79UPzakAc/WhM8w3DB
IGEVV50TtMI+BXvE5cpLj9AFTBjXLIs+ALug//NF/b4ERBBgSXPue1dlVgogMOm6
KyJJsLtz6CM/gvN8/ZBkRRhojEc1K8e8G3/krAw6xfP55RvcKXhiQm65147p2OZJ
9rNb+5fE41Ejxk0Crnua/Cc+e8YYj/Gv4pQcdtNj05o+BaMkKOAW7UIHA867X3rU
5Q4RSv9XWnuoLYgPbVfq1GUpwhjGh5ZU+49KZVpOIYPCu8U+V8p2eRZn1La+vaPY
K6w3F1Wo/O4mW5xd4XVp9L6updFFUJcRMf3pjowYn4cKAzQ79zh6JREvPj9JcSqa
XvMG1gTWPPV8IA04J3WsY0gaXL2flvwSG+MzFh8fK50o1wQXEWb5tqIF+FmUhRF6
GQD9/tOz1Lvjrg+cFXl2G+2Fecg5PXFfY2BVGSG9eQfjyTPyfSPfbWP0DOIA9GK2
C9lvKwSynzh1NYNj/pw6AeRmMlJsutz5SoJK0lsqzPFCWHTGkklPfiaAccQV607O
1fc9EtNdhJM5UjWAtUiLo4LbFtd74zDjmTcqBSmjV2VPqDjCsigDym/DTNeaDyG4
E5YPho94+6mFywm9w91N5pA/t5fEpo37QtBS+0Bg3aUct76m5HNIhmayayzu0tSR
4rlvqaGMuY1zZ/UNGV9tfMqHStFvOxBQtG2rTR5AkX+1jM+3V3efRVZuD1R9N3RW
TVG7BplyEPcF5qICLQ4Zjcz0gad2yh2uqWQMY1trrwl2OYxkX9IPg9zm1uSMvAeY
TgyJtSj+ClZNBYcCvOov23Tf3klnnPn7YxAokJxx9QEjLjkIwtmMu6smzWUaLrOD
y7jvG047/1eH+xrgFE4yU9kXpLEc8PjdCExo4tQ6VcS3Gfgz3HZTPqERqfti8M8G
ECrjCiMIn21vUIRX2Y2s8mWgqOuRV7uktDbCjgZRxd95pxw5AkfUR5sVAui2Hc0a
rx3FNAj7G+OuaBtkVuEUvlkXzSidbouBNMmCm7W4fVNV+XT4NUMUGrsNt8pLMEN8
aBYm43wQP+X0KZ5ZHmF77dXyLV5QX3k8l/nJF/YNXJA+n9FPmYU6B9rUV7bHKMfe
uOLhafkYienQioxbub00VemEN/45+uDnfyVlq6gzO3w9U71n5RQNQ41aBpChQlQr
23Be7eRkX4aLOAuXhcGC/jD6NjBMPeRlzf5pWBvrCg56ecZhmJXxsq3brEnrYLg5
QujElvSAFH9FoWGwX8GyogZFNpdUNj+/jLdICov5qb3CZisAKNmuJAd+g1VZpOkP
m5AHX+ZVlAHcatLUkVA9u1L8gYTDMbUQGcIobdzOS8dxeRGwj8DrPd3ApkADtGsl
wX5T5Iyn1a4TWeTaUErCmSUd3V2MhoO53AhI2KahyyAP4IZqEeY6bI9pGkzuztO4
2uPrZgAnV7FTnzvV2zSq7qV3dx7txKiM3Wa4ecs5arxIVWxQ3zEOfsMlV2ccAavn
L/0qhbrw0wgVthrJRv7CIijl7BAwE/L0v14TZQRfvz3nODF+T3aYX+CM8OTEDfFf
EuC/B8OxoU2JdzmzJPa5L0lBAYpQuKXRySBTIGpMj5w3/dEilSFnkFdh4DMvNtPZ
h2UbH7X+XU1wBEISSsVASBeCFuJAT+Eg+Jnqj4+iSwRP684mhl9VaoYFAHisQHHD
ldFT/P8vwfLrQAS5JAA5seJY6lDxCd4VEDHaXiE9KxLClC4cU4PFMcuOvKRtNpXd
J3/dRlwtIa1HevysTl2mehZccw+dAqsadQwIyRRl9eT/Jb6qnPaMvX9+cMuAbEvy
yQY4LjEsW6LLTlFuhgpVGjI0dtdrDTVW5qVtL1BsRYcvd8v+HetumwWHMwfIgKPh
+GnES3lIucgVL/kh/usBeZBDTZra9sIYNag8ZH+IhJspS5d52D3CsBN+LBn1t4ac
Cu77mnSyxXHq1s3ZYO3kbC/mRUKpKc92ZtCBiniD1CEVwGh2dQCRnRbfgLjM/vvw
O9uObom5fLfVKHXDuTy6lknkQmLSd8o6CcL0w0jt/WenonJNYI7s31nC6NEm3tcp
SS9AeNkvW4OqBYQskfG0yXHqRhvSV/6yvgmC8bkt9784rLTrwQy5RnlWBDQnJq1J
t0LOIZv5jq+ji7Chs16pUxvJPOCQYP32i1vYGCd24oWFw3dEa5670UzaRNu2A29S
rJTTwLbzLvCQVDCf0aNMzRJ28PRgLZ9K/FqgMO9TMES2lpkAsxNji+PwrCwcZV0J
y6iMZxHKUKS5N4JVokUmW5+taSSzkUSy9fQ3bIb/aqvXZ2FFxq0AAcczOfS6q1aQ
+LbrAOUx4aSwg3jNb88pKK9t1fWlhnsnagTx+btibr/6s/62z4YL5+REdfZnaHIt
sqgnQdUuK0U9PFalBQ9M8WXeDErJYDF43m+t4FbSjwhM59AvAoMwUmiZmR4cGu5Z
OciHGnmJOaYRtXyphgATVPfOxWEZOof7NVYbNVQfRELpk/b6T/MFiZrQxOPhy8KD
cds+BKVP0AxWmiJ4KwYCF+PvfTcgFbeUMfAJw49O1LGfVK7setT5F7KSNrbVulVC
ZY29b7wXpfNipiwdDjldX68vf/ea8fv3mQ522j04bjwX/EuXuUH9H3C0V6xS3XrE
Yo++5Ku6dk427v0jgRc77TwKaV74wyKlLN2D71bw8ZbCKHLvtygH/nONzUxOZNDK
/Q/FWHtmik9JZEXEbUA+sGDdDfyxRmk2bUEgAnX9g4qfFaINjDoWAm5ZCQP0g9q+
0keOFIqV//gfIBXZWiG/Dj+0YBzNa/tYe81NkLXBMAIAgg5Rddpw1A5Gp605Wif7
8HM/BqJj1e0i5yTd6+zjwzXzermdrf/A0U8V70EoVNWS0fbwIrg3x6RUnPqm2d1H
zCjEctQn4hikaMmpy51quJuXm+9wfVPtv0sXMLid5g4xHgS5degwDgPoT1Rl3tN3
y42z2Oi9gfq/fCWpm2G3fOgy6hJGwmUvc3WgBn7plxK584aNLp3+lPvDkurDyFk5
8ldjiT5rIiWyNHKwuSQwNEjIs5Wuz6GEIczVePwoIODtQX80W04mN8kFuzusIGEP
BTl80AA6yZZkb3RoJ0WVGBDh7RPOUmvMc/H+klW2YLfIQXUDmx8G9RkElwrRxYpB
yFQ13Be3kLJAatU2UawasDF0h2qELF8VUAra89NyZCken2/zcrRhxGx/yB4W+/iv
4iHEfpH0YeFe0aNwTG9VMSxK8T+s+GiOu0qxu+ZssKvcd9Upb0KkYl+Krzyfmqpx
A/oRcVMZFrjFkmEyo2TGMR/sTCw2r/mchB059o/SfKzpGuYf/Xsc6F2rJmEFGgtQ
sekFbuNLARxY3TqONV2OD+2XFbnkhJZUIE9KDo3FwVeEckExwbUOyDYM61tXlQHp
afYBp4r9kfx7T5/QNDll1mBpg/VmJEGUKqoRQjulHmAX9IM5pkqdSJzPmjwoMMTS
qyATFjZRa5T8hlRixOlM7dkZctLb4GZTYZzJW5FczFqjI/wMlRMKoOBLknALx6at
Adm/KuCeKDVhlWR4qPyVcy1/aXIAxxW381aYNOypIMHAH4FuYczBbJgJ8Rrv2vyt
C7wqfuNcn9iAcDTeTKLVjEVJ5c5GZWbBfyz613omJIpsXJV7DmX3RBc0KX9Sz0hH
MnFn8vLvbBxRn9Dc89rhVezekChmp+drsu8ik/E2tAO2e0XJ24i2eur6uUcNpurr
SGLqXnL6GHCTnPQYflmLWtFceflw4ZNN85sIpJiJZGGlcxQ6Ea08947YeIR8V5gb
GpCiw0BKfzTYVg9zpux43uUE3nYLHERBayalBwZPBJB8x8B7C/hWHUqagc+zUGio
0fYfiSsyO9BQGNg2/sd1rcXubAeCmw2w29jf40Zbl6VLghLzEuXVVc3eXAGkvKRq
W12/65/iSTGSO8oaYtO1+pBxmwmkC99IBGXveFUuDrvh2jQ/f3nwNKEJctTtPfT0
06QhDANCshddcyHkcdpeTN8DHnA+U0qru9dXyYMacn3iIaU3eoh0xnvufvbHYH6L
8/2L7udMy3s8irL1eY/2dUnzrqBqzddu5wgLigefR6+bO6Y1yu5qfnOLvFAIZNvN
cqxKFm1plXfR6kqKna4bg02lGf6wzbq/OfTKZxqxHAdCRM8JUKesi8uxBDXXsKq3
fWsgezWX3JOuuLAo51hwwuqg7BsZvlllQVwEpZBkbjaLF7YftlvpM9W/bgbn56Ee
HDpLGS2ULp5nkJxN7NSuDUxgD7FUqEcUXbypezT5AANvTm9pZbwqmNoysXboZw1A
yrijfv2bX402/I/P08i86SohH8OEtto0aiVIadqDv98yxLCQJ2AyChYujx8QCVF5
K0VdgRSZCAS29jHJziI9FU0Sf8CI7/b3knBrhpoCrAE+PdZ4jvaQ2aqyVe1vgC/B
xEjXT3CzQ5pLLm7BQp+EHadKyMYIbmruwmaomGe/hvkdTfLqzj32vQuwORUG84Jl
4MKXtdNuLpguZSiS3MhBPKidi3vLSZ8JFN7vq0yrPC1ybBklC+7Im52Yhe5gez34
WKn2woLx667l2504k3fPotcpfyBXuDlDZ7bgF4/CHPQKdNJHmMyNZIYXO0DUg8c9
fAENoTtdH4oY1JBfuMmooBCxkfHHM/5gEO4KaSZ0bO2zKyQYIgEa5Z5Jwt8yFkIA
25olG3V182mlDLAKDSvAQ1U92OYtPd2GzWFHC22wPvJqOrExxgbsSwgq1vR1PCEM
lcrTy44D8vGirw3/uTAWRSB7qijtRoGmbvxramvsYSK1/xbBqDYAo/DxXEW0lyFR
LxIhNxFNs7ErQ6QQKH5snOeWoFCj/OFv66/HJTZptMXnbXu5CBawPmG3wTmBFWIG
9Wym0zg6mMUJSpu1kp7WNwEeLoAhAFRC8uJuixcOTNOrh6ajBeZGYMw583woPKms
ij2VmF0DoWsnkSkuUBNPaBX7CtWu3GkNbtHJT7lQBJIUyCsk1IIz2agqAZQbr75D
PDjGh7KHkxBd0lnFwxR0qY6KYEMRQKK/5QFYHaEFmlxmQbbf1536aKUUKdtj+2m5
jK/VL+IfFuuTZvHAKCzos57u2zsG2OVdJv+KokKHkWXKltBFRd/XwYCZX0riDtl+
JEenUtXcDtezBM6y9rmnU3NfCFkdc5NWsxhQO8VGxLvE+3rBQ1pZZuIr0YaRTDiK
LLplzzWU+8krDNT+YowhcgsgvRws+xwHsALAAU7oEtJJT08aLyapar8LseSEQOWW
Kn8EVtRzRC4/Q4UWVcJufitHgdN+UilpgbB630LjbxkvbywfnDMckv0JVsQ3oDCn
bF+rrDhcEopydy8OjQYo0k+aBqxdDGhaREMwByBJK+JaFD8nsKuCZJwqK5TJ8Tli
mlehzO0XZX4XZp00pMJZ+fBZmqnbM4+loWiPNVTB+0Xr/ktDRrEKCohDsziK4PFq
4VwqDSB4fbBS5FP3o82JHjqK7zIRQFvNkWdpdIyoOyLziXrdLq5f7xxVnkxubNbY
wXsSfMIAofVvqokxPh1JalU/3Go5fK1MzOXBA6Fn9LI55EhfylHrxmCf+KmbQNPg
/uwqaQ9vxc05iM9zA1bGc4CZ+Hl7dS7698xDUgUhdUxkSHNKAPzk9gqcrfetpZJA
7GAEj6ji/rlCwkO7mJ+CwrQagJTvkdw59RRN5BZn8mV2xZlWLj0FZOMY2Fl5ob5G
ZRCrUKMn4MdhMtW9WRFueVpvCD8dtQGzB04u+mAqXYR3ByfDcJWT2EVMWmgIFF6a
DQeOY5spmq6RtVjO9Ao3sczCiKEk1G5PZPz8CF171u8aTcKyucsipsjD0tW0HtrE
8kX0T6wAqCiDxFA3DZSJtr+jiHoPQ1OOxE1vYEIXKzSF3kgvfAIu/PHWyCFqH1Ug
7g92P2hfHPU0dEJJbLxj9rk/3GS4fRZK5H4/fB4fEOmMHLOSWHKnQ6/85EHdzFNC
1GP4Byb8qHuPkqXc/tE1gTN4sX3Zw/Jsuikkcu8TrOhBfOAdPqEZ/lD3OOHO8o4b
tn5yncZavMAAbXA0v+/JTJ3CyHQKxXdr9XfmlAQoWeVQT4btgBDQVd1iMpfXc7ml
+qUc/KlN7A0WVPtogITyrjc5R80xPYSKe6dkpfTiRDeAoTtGABWkZHsU5h1I5sGF
i9O5WnhOBfLP0wS73DAr75eegJT8fgsQN+lL0VIU3Xwf5xS77v99WDaqt4zKWpmL
6qdAQ5KdeqdYRrWf9OqnPwnyoBk02mqSHj4iIe7diFMQ6iPpLpy/DO1212ZVnyCE
N+tnPkiOI2Ys6zwfK0IQOgpy4G78ISRTwz5Ge10jC+AFPCiiDCnJ6waMA08j2LQz
MNbi2dqJ9tx9CCuuP8VW9xYRMbxSLRHjhhmHoLrgxhotQiBKwJUVfpUrn672LP4r
Ua5jdTOLRVe/idSlQXrPVdmXm1kMEN+xFS7VUkaxJC4sOYBNleSbG1oHR7WudLV2
7Wcylwk7R2P8JqeeQlRwV8sQAl6PM+0PHKe6vALRPoY84DcHrj6JEw+iQb8ay6EK
bbzEk8gawYWKdFmDkfhWIxbNfaNorKLqlc2fX58R+oEGEnxY1VVpyuxkYCwXhbVp
bLvHl8QmPkRuNRn5SVGlc+TWVBik1ouCRIOQ55j9xDumPCOt3V5PuVHpfKjpeHyK
sH3Z8ZBLvjWOhJW9MKsJVCfLyFgPylYt+9Uuw6ptkhzt02V7TXpIjjrynltxr7PK
FQELRGlIvaEIrq5FeEWWdOhAmMDissf/eUvbDTAamTmZGH67fk2POAq23jvgXzOo
LVMnv5qK74H8NLv2CfWlndDHesQhOOee35YWpztFcofQIz22OpcWGPXc7e7ePs5E
hutvQpsVDu6dod5GsgdUMUfYNL1pvPUhAfboOtR11dtrJZY9R6qPkoaGaT/fHMCC
r/M6tm71dUEhf4dJHg9ptNAs2QaT4fd5LDl5+xLU10hZFKsnNWFlcBu9IcfB8/vs
K74nLb2wwMRj2mERSn8AHfd3RpKrtVAZ6TLNBuz2wZEQFNOmhqj2w7mIfA3E29+S
khgT7uyzssJUHFx4rtgz2Hp6ygeOCdunZgk+pzE0luV+AHO2u2sFIA9H3yYpO++X
9x2DoOWehKro2FTsyGNgBI26Si7niDApnfM/4xZ/Sni1ruXK6o2+HpreD7AVkgdY
6KVYXqiWnfjIi6nv66zF8cUC/OVfS7dHHPSUKKoyMAB2z8sP9s8QQ9psJ+inqH8/
AAOUP7DjewNRYzc/nPtqAqPqI7Xlz84RcINQWV09ekdd1EzjEDeuc/fdeRZdL/tp
tKsdKFP/ULJEgFM3SVoX0zUKlxJeNeI9430lQcbIPMfpgALqip3vvrDk24EX0iVt
psjm+V7J0KpGAUUQDSPDEh8rEF61GGCz+fVGsnUJfMuEdDun1j531FZBBM7IodsU
vv8vbKBwNFDebg7s/bmNyccsDaEqO7AnzOSkkLWcQDMjvroSJtI+0QclkctcRT2k
I00DgU08WkODnvOpepenDwiwQTHPEwFEPuYHD4dhkXw3Xgl0ZIt0uI2B5H7n4Dpj
hH8mEQaqP08i3pcWwwXF615ztYxi3OuxW/CJC/Eof9VxAeoYJLFXlvf71BJoBGCy
IeMbeN+4jK4r3VjEzFY71ntNnBEcTylDsVDMij+I1Bzdo1MXP3fL3mLqMqzRb2mI
HblUKxMrP3DNP5ni9wN8g8vdovzC+/Q3Vs6aRf8jU5yfGRJeOXida1kPB0Vw00D4
ofiNwOo8Did+JT9bmFMlHephIde0/Tvv/bilbQlAe1rm/vRkwnuJx0LFhF8h8Km7
QXB4LLS36XUh6wBMyQshQ29XmsHcIlIV6n1caxIm/b+Uv75r+fhTUmt8Pku+iY9H
48t774V7iXNNz9pAgY4LP6GJ9Gzv8v2XvjjuNR4c5dO33CsAv+0SRsz+7yFYV4C2
CjycqtL8SUDtt7HInUboWJaYHxqZJl8Jh8Sw/youur3dQY9yfJyrcr8l2JygOVDW
7ca4Vu1Jn3UB0dqyQF1EWvXQZiAvWWHA5RRVus/cD+Dktc6ePRpje62aBEnSb4A0
I1W/oXBqQlHRG7GB7F0hCEUfI8wKEQRiRxaGTGRqMkyV5eMQpd0h5I2ZP02ZdwVW
u3EaDCYJ/4bpUhCJwJXfcRf+Qv+hqz84MUpamvSFtNTsw+wJjlFgcx3waTV5SYaP
rk+FgGzkmVLhW2sXHD/zbf4N1FZnR8m7KFQkzKyfJLPl3+NJmsxHM4RiXP+O1+ZU
yKXiLrmRAXI/gz5IfOdv5Y1V7zKhN0g9hOHsN1kTN7Uf2ZWHMQye1z4PBn6+fvBN
cs3z7eOh+TqKgQ7AGFAEPj8JZnSDhCp6fwISnBDuw4z+oi+awaKulgMNov3ritSX
A563dlcinqlxK58pPxT7KkTi/H5D7fGIHkov4sU4MN2VM1tCz+80XzoOBbXNQPs9
sXjoV0gjkXtRWrqAdTfEok7ff9x25Azn6c2E0EpsEWrB63OyLL2Oo9+bevTXxmGK
DIiiDkw2OovQgkHOdz6W6K86Gfrcyq/6YI+53lePYim8ithd6ad+eMvwAiiz7Sxf
TarHQBtliaMs1tKdTnHrYwT7OL+9waMEk4k4cgm8kqz7fTiPb+zCBWv+bvOQZhgp
vfbD1ZPe1GXAX583oni6LA/NOCY/uxhrwhZbYg4gbi3Ote7z4AbpQUYsAs0Y1bko
/7tGmd5HlCpF0TEL1D+Wx+mx3+JdJSkiIziB7OlFe0Ut7cdclZaPmhBYBfiWk43H
mTsXy/VfcsEProTWmLiI2kIMUNk6dHDUMlt3H9cVoLM0P4dpdbtK/UxixgEkbqR9
mCi/UMOxTrvdYGXewTX2Oa/m7XegTWKDnMEDoF/z8KbbswV19yB/p8IDi33Baaqr
ZX218ZOEnhaxlb500ERWxdAUtsbRUuclHco6ijrVGbrBG7xPFuNDFij+CBKNoLz3
QunGrV7wUrZEuZlVPpeK2kfDYDt1Hn/kgDgpbSqh3yIrI+g6ZNmbUA0SNYW4Ht6H
Z9JbOgjRxUiS8AWl9MBlpbibxIGTttwCr2ZryfuBXQvABS2sPgsg13c0PCwWq5pP
7P/A+F+o23RYSAbFTYFScnsPqVUMC1LYa2e8dlr6K4bA/8YsjgHKpNPMi6lDLY5G
HUUrslTzZJkv17opsgmyT25firGXt3pf0O7lU+4ifCDff7IGde0L6C9q9sK/A2gC
YzfEnMY8OrrXO/ni2cDa2Ht62zK+Z7vMANMd4KNnNBnhG1U9xtJo9JdEBi2Mb5LQ
wPmSGz8l4K5QoW4r62CQi4dts1KPE99u//0Aj84yrsvcqYR9td32OeAI0JuyGXJR
0RtXNZU3qSm5LhrF4wQoocti5z5WKkOhxcaB/9w8odFvizzHG3ubFnN2dLLNhGa1
kDyWuAe4864EMm0ksrsUjKDgfV5z7WMSADVZbf7uH98cE6fW26wnBovPOKjFgAOy
yy07+uP61Ynuw3nCOaymF8trTHqfKc7PC9fmGD212Yt3uN37gbTf8zTTHXtadxdr
I4Vpd8BddLt9msKVk3bfMEHrLkTQCceIJ/O7fixTd5ZYVqyhYRumtPBTxEfNwTkW
YUBaBuUJJRjOiED41h9ds+UN3XSDtJ9oHCoh9hPh3tx6u5BysppW9lQDLpLrVseY
Vunl2AunzMyewEKSq2bQ0/LHOlTGBeUkSmEOw1BYAVAKzAtM3NCGXZEQintAg4g/
VcgElvoNzJNT8QPI4l3I3dVzMsJVr26RK+wsaVGdZUqzJaUbJCIup9Rx2a1Yx0I/
pGxtWHLemp50p5KiBddb1wGHoPE/qlfPrFHFHQFKvRLZIGBhXW9pvvOfKKDM7Tn7
Ife5lNx0N+OYSej191uT9tP4whSvkfZxLOEELB2vEG8hD8tax6JyYPzkNVrRbL4r
ApbqNic42x0w1qe6EThRuijGdQajyxFbipbEU+3UtZ/sdr3FF6uD/2zOBr8cGgkW
g41NmU6vdrQZpFoUibBH8ikPrFpdIecLnVDvf/KZ+2m19o0Q5lMvBaEgsL6hdVol
F+RQC/PbwD7AS60ZecuBe66AuPcA0LrD8X2LICwQgRa7bGocK/KdwwFMXDxB6IsY
z/uIZYUjxDP63Er4WC6MCeH3SptkB+DZwSvYTDVvdUOhH0aNfP1EhF660kT4FeYL
AkQOvv7kcF/CMTrqDKiiBIY+K8fNM8I0SlDlL3K607rZOCXLBG3jxMBhV4DTN8n+
ExL6qX29tNzCHex9mmbmums2BqJ886dbaawX827zdEk1vD6zjN2vLubyHGVo2qMg
8D4PZ791Cq43fyfLHMq6EYfIls4jvR/yhrjVfkORPy1rlP/ocI601M8VbamAZqem
Zzlr9nBsh6yllBHOU+iaRWggY4sQi2u5Ya+/knDv5cUJUOoOEE4S84EuZ6SgkouG
UjHfI1AJ5w3YBI2Ks5aVbZuChXtytuCYhEE9CzmuHio0psC/5IK28juV92N5GoKF
Q0q/E78MP83XVQQCK390xCfRG3I0AhB9PZeuMm76oBfRrNKLl0jef4nIxclh7rWe
NgYAsmMiYhR0gRZz5+nJOOD98wNZ2vz5tmYbSPHPGo5qyrL2XA7c5kIDVHwMjFfV
LscN7aXAP73Ub07MLTo4DyVi2gx8sy8eD6mX02YIvsFsLzWJ0+z26ak8O4V2HuUk
p+OiVDkGYUqT0lfZ568/hp/xYwJOfmuGASfZcbqG3+d2GGJinjnlC5/21hAaJ9tJ
c43zdkjgqkL/WbYsVM2E3exObC9OkERsG1oOAb8XPqhlRjh987hi8500YQ5SMf3D
zvyxxgBXj/tXtuuX/Bogune/zx13FVhanAx/xZf457kF5FmUGu6h3/zRI0BTpGOK
jzh+n3IpoK1ak0ZW+qskvwTC/Wa6OKja25z8dtN8bvXzF0SVzfUxsQ/+ncOGpAOd
eDAgZVWF5MKHjq0tXUFCOHrd3hgwc7N4mRi4RkoMmjnUwc10DFyo8kHZuKm1umbg
6r8f+zbs1zpGPFfyPv8OfIgoYzCdb3Ca4flylYwKqXTx9KhYV6karDU+ZW2JKEVq
0jrwg5VcBel1VIg/Phyuwv27CnaSoa/J3WjVy0x0W+qBqbpnmmLNXWHS60KI27Wi
oO/M8qmNf1N8r9WqKr5LNFOCySBw6Pqmsp3sedBGNxg1DcWnbFH1AB9rPiG2BVaJ
R0HhxHFtcl7uxbnuXwdK8PmB/epiEh+ED/WnV8JXlblZ5/zfXFjzXXrm6KDV7Vg3
/VEWbsmrc4hE6WUqE5zV+FkiyEBDxdrsESeKKRuM4/u8zBVjoRZqo5MMkuG/FAkn
85msEUo/nLGwuBW6PwXtbkoUPsDC0HledgeVbOqxnnGd/zNDZ1n+MxwZP8YihCgX
h8g+Oj6Mceo8BD1LJSr4O97CzsGeLaJ8QK5dLgM9+vRw4fYE/3ve9ac8qI8muoPA
1DAJVK28z2X4vG5W07cjwK7Op/WvymgRnGZPMbnq78tlKDEJrDmr3qRV18RGGpm/
haYvc2nfWQ8azpMlm5tcTho8br+DucwRzOE81XjIxjoNA6Jh14PNX12gNRUw2Kwj
u+FKr64F7mEFWpHm+iTtPDsXr/yb4S21A5e2ztY0W9qYrSiqtmSZ7IdCTsG2Afd9
rZ039UUCcWnIvAVD8nP6+K+Z3/PBB7fp+d+QcL4Gy7xUYDAWw2/kHojvmZHFa7Me
xsV1y7s0s4Tt6n8VSid7TI1jG/pMix+r9S5xaNiUqMB5Z/xShI5egPtGUpSmwkr1
g5MnL0J+YNjYyvYhqwiow4YyBakICk2KA+khPFCuZlFI+jRWjYqPKT7jDDRNHUPk
LSBe63pn9u089rZFu2aFvWVw1fNGZ6jWprNs3w1H0TwD+JOEQwvuxrFm+9F39dbF
bvTzmuO2MxTcd8TgPBSZjUKGbKUpL3evr7XI7B5CySGXh1kCvSoCEQIzR1gaF3Dt
vdcka+VBjsBFBRUzHKxKMv3UW0uXb9jD7de0cRZ8LiYNJ2T1Mvk/fWEvwf6go0+s
hDqXwKeuI4uBPTybosINQBQvCO6o4Ik1yxMiCZdLn4i2CPdfJ7t+g7D3M9junk9J
CiCQIuhAb/gleCGixO391acBtKeqzK4Q0UOFwzyrgIYz7dPdv5gDqQaM6ovHuTch
MGUuShQLlkTzGRyVuRVgwzIYOksGUs3cOZ8ZROoPbYM2WJNXfEKuLFst6yIRWIGT
Wa+pU1UpeNHaQKy3oVIDyTz0cgnUK7KTQdpB/1iXf49CgD9xkmVm4GHkK+pxEZes
trQ9q9Swh+Z2Ino4/XsSSC2O+b++YkzPeuBmzctJ4Yf3DaX/jEAwYABYcwCxMoGT
+MpguA5PyV5z+HC0sP11OLo6RPLQQ1koLeFC7EIZiu8Q9RYj5kLWVz47MF1WOGxV
isiyBm/GJ2wdcge5jntiK2aqZr0hadR1RRTqLfIs4nb0qbJtIvwkxfcZWyXu5ebk
syGxrB6ne5TDNaFKqNo04tRB12Hy/oKciQLnQwPZcAOR23h5NT3Zoksjd1FleIpn
NBMRCK/8GhOk28CVeXwmyw+G6aiUOvU9TGWycqkClTRtRCV3pLHvZmUAxct52EF1
AYMcFt88CpupoHx2Jk4P0KqaAu+yrD/qP36RJl+wuC0vc5ucWk0EX5BW8jGu3kP1
Jjkp5k6QSAdOD3TfqXdnhkgSOXddECIqxPv8T+ZJHpGj3Q3p7UcUYqWFvsMZI3Bu
tk98Ku0lY6keFUvNRjjDgPbQFcqh2st8P32740iTY95i/hMLCcvvCU0VQjywG90E
VxwhFSQFeZXlWSqtgyXzA3REzZ9keqBNQ4HJ4bgiiRbt0Lwpw55ms+q4/aJ/f+3c
jxm6MY4xRJJ4LMjrYaIXxUJ+iOgU2QZhT9XPCe/9oswrtlniCYm7BAHbi2cnCVg9
epzcuSyVcgCDFybctAc5GWCD4S/dnNFR2H0y7OZ2Lg68uMETcUNhc2LZkhHf0eey
PXKVN0yDa7UUIhrOaQr4HRtIUjQA7WMJimhlGyz5T+a14/AO6O0wlBpLocSsQmme
R/T5Maw+BgGRFZZFwqiGLHv1U6AhZohoPS2FiAA2Wc5JegrcrHTZ9W/iJPcIHSA1
11u4cQGdOxiZoizHOafc0Y+W5lZK7DJv364qoMkgBiXheyOis+ke5pMMkOEtKtCw
dQ/7mkmfny9MqaTmbvvAyxsaQ73xt4Tgw6t9YLLqBKmPqSPCddDoVV/xl4nt6BXQ
0sVqTX50Du65nJBAK+M5gXNgZGQFbKmFGv6rIKdfw/Cd+d1ephf0K0Wg180Yr9M0
BoqUQwXuPKT2CZ7AfarxcTWitglsplKxT0mEzZba26UUOYX/vv2uQmykKg5N+h+u
PsLWGQlr+TT1azhIgSBCdKw5KS3ZI+4HiOCelJMgHVLuJqtRj+Wqb+Icj4+//4bw
dMzEyYa6x6M1yZ+FpqIeu1PffLZqqaYC75lels3EwI2lkiHzvvPxOID4hhuDCIV2
Fqv+zaPA8x/eeAlElpidobNDyy/hs+VDat7TfP4PUNoo7d75O2Vlkxp6DaIHtssN
3Ccmoh6DLVMxPLDWF7XwAc8bCdv/ZfM4XzBzgahqsC33LDCJukiKXm/cAuDujm/t
0s+hGwFKgvld+sRSz7upfABph1w+KC0LF0SsuwaUAv4VsKt2dvlbZze9ignWuK+t
7fbA6RgOuUc6VvKfIew41/eyllBYHe37PiWppuqYLkDPgOxK/5EC80N1SpmKBwgx
xgayo54VASL1B+SX68ly/XHLXRyg8i0c0UWH+Y1y/J00Lq/BLuEYhVRnkujmVr1F
C3eOmr63vnoYD5DF4efQiHN9SHKYh/XuAO/j2Y8xwM+gudSCe5qXBfEuLoEAxik/
YzEcgJoEqpnD4dIx8ZmvQwaJk66TRo+jMkXxcNn1ey13hS4VMEfkiXFpKqH8guOd
95n47V4Qm8XJe6VIF4F4d8nVj+Hv+tDRlrafKPX2fdyKnUswRuCe47/YKF2yFXA5
qqgqpEzqjro7qo985CnFujIS61fR8cODRWBWLbs9hsuBpcu7UTZjjavVzKQKxLYI
F5WOQU2GUG0CDP/+84ZJ78iamKoWLjDKNPLtAvw8VHe68AaMdXEi4btJ0BuqFtT0
aQoEqs0LbbEG3janOYqgLGIfi/o/6chFnA6Q30q+R2M9N+Y23jggUmyTTqFakqPV
KaFTVTeMFVt/wtNZSvLuZmkKF/g5U6x70V0sEE4EJv+e2VgrF2T741FXx8/EgAkC
CdOgJfwW1RWPiGe80rNSPKtwjibLVzBf3JmKgx9naiEVzP7fsqzbiBuPD1G3rjTC
5t0A18X+d7F0bONNkNHQkBMZNJZNbJrm0wFw9Jd0IM5Z5EE+Io8K7B+NXaeD/xKw
8aUX02XjkOprsvUHn/zpuNTLSYDGPWLqWNwNDr/xFEVLJzZSPGd+SKHqW+htOcGL
XJSwAZL7XJ7p7TJWbA5f/b2RD2qPEs0TUUGw8kL1aXoy457+w7kI1kHRtfuJrCMY
p+4QKfkIZtQu7fmODV2jExSB+50lLXEXhbqo0qy9kLrdw8VeE2BTkHVypkwAbdH2
OOLhVw5U+XCBlUcNIEwVmCKuNnjWEo1vY84svdxJwmJPa9r7RcP3mYKtpavcnFxk
GiOYlA/Q8UiT/q+Z1IkRDfyh8U/VWDCk9764P7HfdC+BizVps9WVjvu44IOYsK+2
gSBSTKQFEdZ/pE6ErYvDgl0/ZTJsAAsljARNwFkOqdnTWtPchdL0IFJDA07BjAAK
1BwTuZfhhK0EZEFZBlOQvvxFEzt03FGDZxSdTT6QnkhMmAOERNhgm0A5KLDxK+tU
7qdPfWz1O1x5n9yAGr6JsRzftJhPBLXJvKkXUltQn4btebeiTlDDF0x4zz4k0uKt
S+dTq6aWsWIFvQmNbIW7D4OW4AtrUhVxnOREd3wjdHMorDl1MKVXGgdLsJ2CfEDP
iI7hgQsvihOxsDE4IuOAKlRz9C1gPHchJcxuUJErW0qM8sYajRtGSNZlaiSpfo48
1J4DgPzH2TFon8iF7elVsNz2XzaJGdHbOezputHz6shyNuX8AXAheMbNuUxofK6J
WFVN7P+8JOYTdQR3aszwbOnfuEwpnNtGrIxHVJ6TXj/VYqAB8g4ohd7nodhphEAA
mDHgE40UElZGgFFz6JW3WJL/nIasb7QdF72nxJDac+PPgSIlLZnlCldrfPGHCkFR
lydSvgRmgzWEFpwNOel7Zr7sWzXiHvzJZspNmeKb30C9r60YRSNXmccmPsNeqGNt
tuf0yVTbQPY8iwjJD0N9T1JSI4s7ofKt5ZDB6GGj5dZxOy6tw295zJeAxPP91EZV
4fjSvoyQj9OIWOK6ot/6D7iVl85kt6Z8z/f4ABWDWpOHijYUGMJE+B+xdQj0FzSV
V5KnnH4iAVgv6iXvgtf1j7DDgz9COuYC5DlAuAGHReUdzeUpYyXlfaiaUVmZZze6
wIwZTvQb6zjCKsprQuWQ03wqeySQDCUdR3B6ailU7IdfKJf62utYwZeoHdm6Syzm
exNqUMdB68jp4oWp4USKGJEEwbfPfYpFLUjye/fNSNwgPJcIMvYnA4+bWpCWTr2a
zTQ2DdaT5CcXfsk9i4CxjQkOX+xoXvTWoKWetbbv8uLvRBc363Kr2PIwPPDBtmOw
fV8QuoAD8Vx6Yy/xmPFxaLn+YOTioCfHWGaRqm/RrxMsjflaCF+zAESETxMi1sPa
XofFcl0f4Z1Afj4vwShDdvIwztupKKNnAakRmLZESzpJMAqJs9cL4dvVnJCw3GrG
KDqgK17Ge7T5bsRvqQYVtGkUT7yXIR2UpGvViMYGdxV6Ox14aPcYkTHCHPuW1s2v
NoZISPEbEeO4M7leaevHQYsATmp4e37ZhPQTIoDV0GQmcBRQ3hhI+v/o9oMPrIci
l+E9t9i4v7QmTijvEmknOpTaqzxF7mnd8zhAmHOdx38vvd1NVE1pYNF5vEkL5zYF
TJoWt4PP6A1Cr2bDiXXdi0MQ/ubJ9bFfDVSn8CcX/kJ7BV8MjLPM/ZpS9eMklQC6
1V7Toubw/1uerQ4LpMf058oj2yevQ5xyvT9umsGy6EE5y47O/l8APlViF5sY1ubr
CSoTvy5+If+iA6cyOJ77YXMah9LTZP2I/K21aLuVFQvO8pNsARi99a8K/m/97T6W
YEHhAa74azMcQVbHF3P/SmWb9pssnH/jRDh7FDqcMs4ArY+YC9SP8Hkwm5uewx9u
tZuwpW9N0T/emo/cZmLvCYT/GFO0XrDCXXNoNhs+oMC9AGY4+VlyWuq3sqXh4K3P
+TBRQMpJen4k/iYEat0aGaCRLUjOvm7nxIKsgSHYq5Mu8T8GikVqGARKntiKlBtY
N+iRH28a07grFOkYtjZmD11K8D/rHPUduD9n7uJJVzQsXultxuUX+YIsGilSuesj
5DNagCXLGWj2PJltOAgpEeGF5/qpAh1GywcRU6VZkqRBRWoixcOfb9GBx6Qlrx3i
TL2496Czna+ktWL5Gn1QbnYgBf3hO08VpXwJ9UieELg2nmEeHZHwSLinpRDbZ8c7
IvziOnZlpFmtt+BEr8aCMkxxJ2v80Q56CpPc3mZ/Rs7c3mHbMtoSv1kThpc9ZAqB
rwzRVxZAXEbzvTaJg5lB8cPJxyssDFAoo8ewys7YVKeYxSie/QQ2Xu7rGJlLeeOI
HPK8AoePA6ndXx8qE6iOlwRZklsRidT0Qe/VnFLbpqxndmipz6wWjUQkWT4V9KIM
/nfqWBOD5+GJfoxnvQ/uZ02GTVy465b1w8wjJUIs8Jr4O9iuA/6T8zbe4dpV9nsZ
n7T7qjiGy8SdfLiKLTGQv1AT1Il+oO1yfSNcxpptoMXvZebTs5Vnt1qkZ3J1TzIG
qBAtexA09AKBBZ00OUT/oB43jzMiV7nqluKndmncPb+5cu03SFdPWhb9oJmCBciq
ceolA/oNb4Sh2Q0hOr6EqnQ7n1Nz9ig88qI5h6JxVEf2rKAqFOqaiNPOmLFoDG2L
PkyfbsdYh9057mzjdo4ASxCgIA9WYjMmZR7l+Fi0XVAzNVgIa97FY3FhdZAtvrck
utaNsinrLCQKFCNWuT6boKuoEFieBIy0Qysiq0hXCkgTuq+fPLOZMezFI0yl1kcX
vr3QGe/BNyNflN7as9mDQitdJW0+EZJKB00L+l9Cg+WeUMTTjM0A1qMPahsc+N5c
GHV5Y5C8OgYZADk5xguUdFQwumlPyZqWxxbW41ObJPwKhrf2tAduCI8N1ojtsEvC
uMOXTziD6+ur1FXQJ8p6RyQWUl+L9AxxLrHWCVH6hpZ3peWlgQZlTl/A2yhK8bBE
HyRU/IQWQ3m3LMUIomeQJFOqZfu/Yrp3mLrtcj8L2LXa018238pfUId+UtB9J3Nj
HNDrA5iJh/nBEsY31zW+dW5eIt/+8Ut7oCeov+cQFGJ4Zz0rvNoJtTG1PfPejZpo
xZKf+kSHepzb1rB5Uma9KX/fHLD2u/B2hSopZQkvGyakDfhOZklICJ91pLcTf4sK
y0j6/ioivkyREZWlBWCIF7BUJ6BaUcJzJHy7LITYqUTse4nCRjneMukjWO3WDfnr
gvKnTiojxv4rcl2o6yJqp5Yv8tNoeA78m6gXyOeicfdrFOwf+IXm0PJvsSFpt/Ob
/YwfYj3LuepVFTRJXqg7CaljFvKUnuK6SLYtDVk1BefvP/N24S4pqP201Z93RLaG
oiAMRdYKVVnP3JVSlIleRLSE3mxfW6WfaqVu1PSLxSRgN4Coe5vhLqI/ZfGx4RGx
g0fJJHmrUNDrZImOzyF5BreVeg+rBWaDax9Xb34FFrY4sPo+tK2B0nfZUDA/tzJA
F3NKmHypWeYdlSWJe0e7uidf7wYiaDGETEz2TBmvz+gb38mLHmM6Uv3PrNByvD8v
cQFWMJ529jYOwE+7h+eaaOYAV9smwoXs50Bz2tCccUVCtAYRJ5AQn+mz3C0Xht5K
Y0R2/cAtxgcT1s8q7+p/N3u/Wfy7S4QFLTd4JogH+xikxU5iKE2E2igqNgKv7jZB
S8bkHvWv+7JuMCvnTAE0bBU67i1TCjqgd733wrttKhOr77DJAs7PktPKrrZlaoDO
SwaVLDLv1RyDAikm2gF8Z7WRWoEUHWGJJx79YeJigK07jdMYJuW3EYG+rrr3HCwu
WcQkiQgfXOhOfIUN/P9eKVeWdv815t8hOhQzsV5Ri/dgMcWJgsCY1TtSm7xroVyC
6FrzisScIbsI0+z354R4u12jqYxaM1QutgF47NzDrPEE5rBw0GQ6sB5TwfnWMElJ
Ya/6PBog2FPXe1fdcd0LnFRfVDlIw+Eb1pTkO+eWI92Upx5FRttuF0OUbg4CiXyj
X/+Dx5vWZHdot3RjBltMVj9c7z1RayLm1AR41+ZJtc4LUnMWZTlvVVl0JjjBrM2D
f4TTO29avl1pAsAUGWjZsQ3lwbzM6SZJXj53eEY+cjvQsZR8bU+tB/GipLLfWt2y
8iNUQtNszvpfVdaA3vJpFALgGORfWNcXbKGEzQdAEmbq9X7vi5O+QhP4NbDHQ0fn
C6iDrTCWMvO8t8o1OvBUkhcALSEa41z1PdgkYJvfMUZMdgGupIn49KAbZHkZ9a8s
zuy4Jg+MfkCUr64Whbg8cPC99l5Z4XpT5B0FAyge3O9QvirSHj3SBTG81R67b7qi
cF8QeUxyhyw36ChVLLZY09cM4pgNp5nj7zl1HI7dgoxs8jjksjtYtEXucmvZXEcv
VSbthAAbJSXJuEj6fZh3yKtaB4lzvpwwn220Y+aNPKkg5gPvzKFzovmlGfiw+Z2K
vAMjaHDOdFRBgO7UfwoZ5t0ikGoMR5hgBtf+mBf7B6Cxp0/fF0o2aNXiKiLkfnJi
0kxvEKULL4VfZghqR8OfpbAxXvomdQFNzhBLuNWNNZ2BIqkLLHFZ7FaPHJqGwZW2
qYLyncigS62dPpkmrkFvTjcoBZbEr0UZjRV0Y/Qzqq1eYl2DJ2InDw7G0IkZ1udQ
n/uInNwQK7HDpl0uiRUPbtvXAXUWR0WZ8gvi9BR12ITbLodONHV5+YEfxxNjwZNj
OqOAyKffT6qkYakn4UiUwPF5WtgdvjJ0avunVUtIekz11Dr11wg9EsmggVOgDoZz
iumtdcVTz6iawZ77Z6/vUmpbrPb6BD7a6lTYt7mzdm+2wIFcs1ygboF34vX6iTkM
lxR2TC6DPzxSjWG+AnQFgpDmcWoQ868iZVofQMcDFj6P9EpMnEcQgs7R6Y1H78eP
QnPCvleU3xWF2C0KFr+sOu5owA1ZFLAi32869KAQEqqEIFYW3XTjZMtjIfP92zGz
NR8jpLLODJagGL578XjAAEegmPUGqefXd/4AYSr3Le5M+KiX5xNO/1nOJwwfpnsi
FupX6LqMf0JLOz2naCuHtpsS3i7fu1654h/p261f7KYT4VzRwg334PgFy9RoEfML
cP1xjaz2MTK+HTkgoVfxB0kDsRZzRTEOhicOm6Mp3pDUCHaIIx520Ipu03izW4G2
lZamPxr3atFPUX6z2NXLjFZm5fhXTB7FSL8HeS41QclUE6iVBCTxz263baK1juTo
EN95R9iR/udIexfepBFni350QMtXXNJbi7YkGk1E+q830Upe8fNXfStgs28tHV2Q
Q4cebi6nkQHzcsCOinWoB/nI3554AfxNKoPngT06CyPJGyIYcCRPvQNr1GmLyZXy
rkmZ4BvudSt0QsKDrhFnJBaCvdnOkBnW4HN6oHf6TKzYp1sYPYwx3BB5bfeOv/0b
brn8Ym5SS36fwDTPUqo20spLJ930sJna81wEQrq9NBvSTOpkGBKT5ZmY3MDc7yTe
ngLSFNw2dQDpU7RmGX23RMlkANeCR/BRpHQW5G1jGnZcO32lfp/9V7GShrqZCGJF
/9vJ22dQ0F64TQxfqi2dBcs28nM260zfTxSWlB5NWpKRy4Nz7KyyRNizGhN3IaS9
Bpz0R05Muh6Z4gW6IaFNJwxvJddif5qD4tervodSEPI4IZYZZJWbTi8mlyB4VDBz
JnA3k5iHeL1u7jyRO8JBqRYlMROd+dNyQdFUeChU7pNP1Z4m6zKIylPKLTEXnI9M
pqIJEq4g8eMY9udp0d/wZYJeUxPcKjS0cX//e0vohAd7x85mknyFjqACKkrijdVA
UyMtzvKOzqOIiXLaNCllFAjBCvMxYvV4sSOSpEgj0bS6zMXT/cEYUZUUDpOPTPPf
3IadkjXNzfHIj1inNgUaJ8le7vDdtPBIegcQCgFUfrduUpzEmY6WNA3sUis/vWAF
Ilunq+aZuJiFpXtSf49QRrdqnbHHLCNrGQa5z9N+sX0k0iM7NGzKD5SKch//Alkv
WN9cD+tNNJoDssVFBelG74uSY1vvwTt046B+N+f1h/BSFxB4WUjThNJbjNv4BXm2
3UjjpaEsDt+0dYkX24U/iy+3XiCC3Gi7cK6hinwaJrFvmQN/faS8aJtgTIrXyT7M
0BNsHIRD56CLFfLesQKOwEFAqeu4gQna7JNpkSpk+g/vWGDh0tU96wLJ+PCzk0I2
NmxZygegD9Xr+n9lsB+fo1ALE/7VzQdbH9QTGQzRiYToIIZM2YY1QqmWYnN/7FBt
+WvMHBWriGU9YWQl4qW35hEwk0CWbx40hJJ3mJTCPrJNHn/TFWeY8IT+9MnZcBXE
Wdbd/heM+3zkTZWYsxd62+aQunX8ChY19MKxTQJE6P5vN58uNL+sFZ+Emc1DG6Zl
rKp/xzZNRpSV4UDDLvBO7GrdfnMcz8yiYxqi0eg+4TNhh/NVnlhCYFqIOq5SMZga
er/ZfASw1nqKwdTTor8e4XB9uuL/A78injvfLSflkrGzJeNXMf6yDoLrhz1g8MJP
lU+O+Y3cww/DzPd2k4gRkfADcU1sDo2RMXwGpZKMFxfVHPk8hN4qJeucEbNwTEh1
cZmiaRmx7Wltezxg8cwLjwzXUwkgkPlshFYfbOJ2XkJ6Ur7/q6O0Yt+QQMbitkWI
sk47KwLijlg9tijBu2lhdsATGj5O94EOPOk5wIlfZrVdsaualOYNW/zaTifiG9p1
rzz3I2+uafFKiM81SFx79xmFXWX29TJ5ZmzQqXd/pZWCY7noQdfEZV5ZA6/gXvAJ
IjWT+l16aMp7jqBClG38LMKtTy5p/dW0iawAeUqG1oU+MdDMTR3J5V8qP73yC2Zq
i6PeGbRizllhbeo0ZaO+7myga3BCy6qbjyDS4U/Wco2jUUjlTzb6bQe9oUXqc40V
8bWDnAFM6RDE0OLpzOMIrAhTx29b0Y0pmgtTM2LJcTMeL1F6atiIh29NZAi3Y2Ew
bzmryZPWPHUXFbatq0ZycqDlZgLisghm5XYMWhfC1MgbF9l+c88iE71ESb4Cqmfy
/opdhOFe+dN7Mg1B1Yz854WEfnc4wMPIWg/72o5lODc96Yjo4TTITQBCbrMNi1EV
EMuH7C6hCJz/CmUO9e0By5uKq6VaiAMbadRAV3dh7XjPKTqLC67o65bRhsqUyKCG
0E7uu9lZpJwOLxDnwWzANqLSoMB7DqtJkLBS5DGB8jjF+3Kyckrqizz3xH4UR/sQ
/Gp4g3jyaSg9dfzDYv03wVHwgtx8D2FUKoDJxqcFnteLO262U1svicPTgMMMjAcj
aWLfywQ7lqa5hRUnBm626mWlE48H2woPaBgUqSyPRq3GsFCCEkoEcqKEQCSS70iz
fPUyMm1Z5HbgN6grei2wBi8FpI+uHzLHmHWyvNDblC6Sz94+MXQwui4YPJZFutd0
7wyBtUv2kZHKqq2zg3KZmkKO5OskyFUTaqL9kpEtFmJ44+697+IAcMPCDrhWpaPp
alSb2JWR+/L3RC6wgUPXXnIT31XgtijhYu2yZOhQ0JOEJtLMLZlfJiFMbaW5wX07
nG1knI0D6JkWVsiCazgNw7GLbYesIFZYCkkifQix3tyrEPbJIKG2JrBwnV9sR0Q6
DBDipcgc5yH7tgH//Ligmd/vQLE17qw6JzHwh+Gx92DfcySY5FSgk/JE/eWg7emg
LF+A/peiT8w/grFIE3dyfiwWibCnK6+p1SEqtsRFfsLUlCXet+gS1Jg7jVHec4av
0OJYhTvF6NQHAfk4LF7zqN6gfPptNCV3rAG5mjhz1wQa9A1w3nZfWPDzNiXSNRlx
7S4tCWwDcImc0JzWiirsKCG4tWeTD9NT635mhLlA3Y8VP4FsYXYwqpan+IEa6B+7
k6pnvWIQ8B4pitZAyAqy/wk3Ulb/Y3FfAqx+qxLcLc6PkQv4jbEONF+63KWM8rZC
nMduMO08Aw2l+2i2LqFKHwqPVPgoSzCQQW30Z06mUN+Hk4aAGPziL0yMIqUs4o7x
iZEMMqi1WLkIRObpejukRy6fqmHP17MjcFWo2vgCmFksxPYSQqA8lKbPnKoebC3k
DMDMBKWNZRZmuMS+6g6qsYh9jgBNV8C516rz5YEmUC/70wBIfvO1Yczb77/XL7XL
N2IxXDJtVcUNeRbGqdqZkreUMvz0XJEb8IsqCUFoJQ+mmQkEZX07y9ChZb0D+7Y4
msLmKsWt7TFpNTq1Uc9j6aNI40u+U5XR5vmH0ei5suW2CkHIoTL2cONwBsdtVwOJ
AVoxM+TIXWqOSinyCTPTQQYdADlyMjwJCLcDBKbt3+1m0A8xR4WMoNHvdNq4g1zL
sHJxg6PaS2T4WhtKrJiq4/lCFcK2JHBhcD33U7ZOvxzPPAfgygbpIIXfm14ETt7H
uBg3HmaobFjhHsWfH4m7JoY7sP4ZHNivsVNDhjUPemGZMd8k4/2Qpg6iP82dUId0
P9uHDN1IKUgqzkYLENdaO7vKQ1iCp6sRn9xf5DreS5SPNylJ7nzl03TPtmEsgD9M
yMDTh23kj7DQ/egM8DqJk/sZHBzFGFxkFklbmKCpXUuDsPjN/A/A6y6K1ilCSptE
qxUS43Ea2NvRLZCA5zuLcefyV9z5Vk+4AE0sYoCSLWDTUqNYv1nKVI9uOF7r9EFo
AGnkPSu2HtTvUW73W8Xyp/2vq69nY9NXgckZOgKX+YEgaGKtV7xeYBnd8lR+w1Lf
E6FGSYqfK4OqctEWlNLY1BgQ0wNIkES26QwpxuNfVZGm23t58PYmGeOvW/Y9Hg9q
T53f7qnjIU4mj4+e/YjTs3Wg8C5Kz6Lb+oAtbia5tX2nJZ2PPZtBfiHu6t4jNbNy
OE8TLH9gqDMFU3TpgIxhxNbzlqx6ry3Z1e0FflssdT832C8sY4ut1GzhmkkjZCj8
Te8czVtGPF7Auj+i4/cJrdpwuq5EF6x+LVqR3NJbIiVwk57I+UBE2fEm7RILSrMZ
UMY42je3S8uP/wRBGfhfUa+zLjmyxnByHSVSlg/5HxT49L0DjQECfQCPwTv/Zvhb
nE5OHBHygxpDpeNlZgE9uguVL/OLaOx0XAWSgznmqT5f75cXrM4iM5zbWQ3cM3YQ
nSHZcIWgbsAxbTlW77c8N7IneOyUzXXENnzO1+/KrszMpAXI37+MXTvpbSN1/SR8
8CrYUBXp2asRW5bff95ZfU0zdI9F+azcLNO6kjzeWKlrOjj9UnhxXqHZylXSXYAY
U4ZH90a8YWRSfQ1e7YWaEfqK+KCbHIen8i6GnDveYs3obi6FxfAoiMQK0Lh4W2Hm
RP87pRK7B3ChMZ2ki5q6U6+lNP9A1xQ11VGjsVDqaGTHe+lASJ00ZUV9c0wGI8Os
OUKN8ZhwHJX8XfjqNtuUpUWWkbJhAqGfUpno6N5GRCQFWIH1Vxx0L0qXJvtEEWCh
v2RShTwjT1atFpk/5tngf2zMxSdo9qIyBMeDYpCL4Jk7vcH1twv6lSN9Wdf45fGi
rXR5V5tqN8o0GIV8+/yd0WwsIWaPuqjCWdDPXTwi2hofEUZV03iz8Iv3x/Zc/iBp
AOcnsBy0Ctv10Q5m3MV4lpyzM48RfGtPPf8TR+rDwHPk/XC81GusCrBpEDmvksgT
6JSLXeDASd7UXV5j84iiFuNFS447AxZa+KwSCMuosNqSBynGbnSeOV5ruvEwjvnv
tlhOkEDe3G9QGAPQ97vkUZ1K1dUasvQGpF0xm2STrR7IcHpNl5opc28AOzfqB5e6
2UhSBx0RRMlpVawnobKyeIVSbsxaQtf4EZJFDBkgUMTvCGaMQFXbNfz2EwalMhgn
fYLh/LG3IwlsV9ldBnEHwfx+Q/ALnlnusr5Gp40Qy4X9+ttLbOcZusYkeA/k3PBt
ZMIG52xQ1guShIMFkjtREHG/0qXGXZLlIo5b90Oiter6o/ebAceE6LosET9XwM3d
PjfgjBqK4Ai731j+HkU5DekNphsMXT/nlH1SAi2aDJQKHf7RDiW3o5iPgJovlqGI
xuzK3UPSGzG/VWbTD6/TyRbuJMshFVznaCKNHzn62/kzBd9jHYh33TKqjKsoYG6h
r2TvyXlGKJj7+f3dfuYryWOiceu/K4eRlhSZiY+Jy//qqzNclyhP/785BuPh9xQy
mSNoUk5LRhiLWZhyi3uLlLgxta2c21+O4lvF8sSK3dDtZScxpdSK/xtFpWzveLgK
x4W5mwZ7sk5SWhGgSPyCUyju1wxTvCKGjz6pIM9qyt0WlGRN5SLkUnAqVvYasBV1
tp6cH2tw8zy+CJWCFYU8DLChlhcZXuao0RL8uq8ZwYRqEsH4w+MS4OI1JmCTMLOG
fUiVjAwOvZ0DVYRQXIJSlEc+VpbtwzP5urJAMUmutJ13uprghzaC5VMQMmwIXFXD
+akGaigbm6MvyYpvaDefQDLX3FM0lusclNRg9LmYkcocTAGjJb1MuCe/MZDeLE7f
Bm7/H80g0o3AL/zH3Zw6LmoPJ/WsoLpQKh2Bz8R1UorQX1T6HPm/W4BE8mjPOBNJ
QTACBrgwWWyoVw3glnUltII+tsLCy4dg89IlM2Y57OnmH3jfnseYK/q02o+IZTWA
qJxjB5BPjIrve1QcLunCTS+HCMIWVJPQZx3Z5iaFG7gNQvD/TmRUjnM1BeUcwong
HUIO2uujmfjCgaviHkYuRtFFg7MxccX0FVAFYDwjTKex6GuNie3xXuJqd/N0RGYP
+qP9hTonVVB3SsM5TYev03+F9dNuZFvKne04hpkYZz8qbLrpGHs6UaKxChwVMKx3
MyuiIMNG6TQPAY1QKV9cteJbr/WBFmb8ZDtEWqJ8eT0RWDEwshIwLOYEktag8cM2
Ft+9Mesl0wqcAR3yxiHh/8ARLJBuavOibA1PDOI8GfedTdSSxy8vZTZBdGTNPqoh
qsZd88FaknYd8OhCNAVVoKkqNR+8XjgXz2kkz+UNoy5q2FtdXjAEYC3p8VkiCkVV
2DZvvNRmjNaYVUWFHP3SXckQUHJM3UThEvt1pI3LIouKmZwypB6dsrbt31vngZ3/
eky+7z5qlTqXR8W1izb9hsqx5+JqB76EQm3lSNPvHUYENbYp1eg79jJoHHUySlBO
IRd+7uqeVHk0OxN3CJh95mqs3Si+w9KzQzU0H9hfLzQ6GL0UIoRErj0QJeneaMdk
amLgq4xUDvp06VZxiU4pG4NN0xBuA9bWkhuCr1sJO81GU0OuUJp1TngPI2klJ7Th
lUhtw0ZS36M9VnlYJQt0MOUkRC2lCaXWAJAxbDeCvewvoq/LRmCulUQB75VqCR4D
QSTO7xbZdw3dZEkucx96s3GZh/7yz5RPJaSoIx+3DQnb5Ky3MyGIOIA9xxUaQAPQ
9WBO/15j6qBMebM5QtTkiqMfPEqaArJ/SLb1vsKAYqsRY/Nnf9XPp1UuNBNfJxqN
Yn8JUFojyGh+nYzOEPBG5ewJUYxo6TRplxif+C59BFn5sp2x9fsRfa+7iPyKBzRv
l9vBteBNJvlSTbEb3f6vEfeZeMOEgTYur7FcKe0D2bjJNGs475csXhuNFYi+n5hV
jmpe3w934NGhEgkQs/NpZu1Z9LtSSuqOILEF8RjMTBU7778H2WW2GQFhq1yxqwNp
FzQhPq6Ekk3qYNNJ5whIt0k9gFJrNQ904lN5rU0BuaRjlzoTojq3+IrEiMZrtD1G
vxNywI0kQxt4Wc5u6+ucyOt6odX1xQyCueMPejVjHCaY2mwY/txsOlaSivpt5Wtk
j0TIwb5swm/BRYvtG1OhAuhsBux3igUlMLi65CuYcJWIxS3ac9MROFvrrIgcXHr/
fplTERkXtvRVOtj1xDqJ76gQ2wURYP+GO9zHPWCcBsGyN3PnAJIRwfmuc+M+T/r7
pRPQsG16M0UGqBkKRNBEIeIjhck770NsuvSewl0dYxu3O2a7upCY7H+q3KdoswKQ
DujjifoaCZhc3CBC7Bc2LvJvBi9o1yCoV97dtIr16iKYDXAyRhSrw6421d3LByF8
i35xgsi1TA65pOL6J1XHT9r+GfNHHFV87FM8U/J47tAIxxpyDLp40eFyQ+SLivVy
dtl8GS0uSqqO55HaldqYgEIEM6KkmDrDgtYbn+XfXPT6viLPlRTDATDY7zdANkj4
GeCCfbaLUO9lZF0PhSHB9PDcNHlhDr+yIyZhGH4XyphYZziEZBfy3JXkLY/OpHW6
3iiL6PJ9WPWUXAAputJTExe9ogq2sMUAJHzdvU5iXpRCQBbgnW4jmvrBJt4Uw+Kl
1bRKq5hNEm/dOIcETy/zkl0HKHSuQsPxGheufsayVK9hYNFYZ8r6gWgbSezU9ams
d1qZy/expb8JsyZbmf8lS0o44Vya13Wc9yW/R0CzM7yKTLciIil8g+0VJs/zXuU7
8U66TeXh7xD0SJ5bkhvP7FL+VG+lgakPCg7BSOU7AILLmFyVjqrhlEcUFOFNtn7t
lL+y2wrjE16qQJ8XS3iqF2CcOfm6FSZqe8G9WcWZ+/fUYNW1p3cND/DtauWYKWkS
A3NtOExB+tckcg7B1JeA0VPOuqw56RfX1+jPxRk6KJzZEQG1zLxFH8Q3dZQKDpfv
TwR6DR4KUBDQUJQbk05qxLdEYIW4C2bV0Q3PVumGdXxKeemAcBTDaD4lf7iL4RyD
QWutYWIRvtueka8SzA02k3HRVhmvAtkAppYxh587oRhJgTIfpy/AnGBXgeD7OiRv
K67y889hp06qSkoR+luVqqFjJmgHz76z28ATLTG7/4twimBNJbM9JUH+5f9ePTI2
yJWHtZy1VnYvIyMH4GefLm3ScN0yA4/465QXbWt5NRaQiTuhkNm2AhH4Qlr14Xmg
pm/8cMJ9pZc5YeHqdd8Y4pt7dW09Vra+ooZkCqzT0M4FjX2BnAi/faKtkfw4ABHv
+m9kOWrOV8ARMyF6Zr6E8RRwks4P+kSBbEDF5sEGRBQI9QtlTQq/uul1r++9DnUT
fvZu9El+RnIHLvL2XLrP0dP/lZzbTkALht6RJsv8a3uTQyvbyuN23B5qEc07Tyfi
ZZWBGpO6u0bx/Sweok5vBms8nnH17LWM0A/t4f4x4TCx5VuB756meYmq/NoXdWMh
tYoReYIcXfqSfZhELWzydxpGwSw/BE+0JS5Y+hs758VwURddsExF3tD0bA8Sns82
oFFR1faY8hMH/0+0KE5ckJhgDxweLGn38PaFeJvz/ITvAg7FgibZxZC52tqec/YA
SuHeCCriK1qgxYtbH9jMLtVwhcZjFsXudNCv+kwcYGGn18uiKLdh4zid5k3rdBc2
rQQRPrpjvxA2Qg5RhHvcc/hd37OrCDu6S7Fy3yeqy/gB1r0Yn4rWe29tJd7uAqP1
HyXLUjL3/EHMHYlXQEkPsm9iDDG9wCYIJEpbhq0iO1gRxaUMJ0IE+YMX7HpfXi1E
+5RiUY/mIBdwHv60T60KclPfK9lfeSXoUOMwZvtJ0adMhtB6Gt/2C7GcBF7Cg0AN
cwQzDwJa7FAITngC70i8Tx/3RFvjSWcqmPxSj1Qz0EOUEkOaTe0H8nm/YRqUqJPy
ruipvEW68cOSVLtc3ZFVLUZ8R81IgOAnSVzvjnQe64QQQVaiBqxotAwNMAmeKdvq
5eg8LM0GeXGS2ZkX3ZD8ZgelVTKxHBUcIDfSEBqwxZHlu15KZcSPMCiVgpVF4q33
ExIJk4+hCJ/+9qv9zero3hZIKpENGb89urBjCaWK0bmDCkZDZCEf/y5Cx87KA/1D
UdLy4o0xoBUNCQFxEpCgQINfabCQXQ1W2AmpV7RVlFCYRdz0CjIW8yWnA5W6Pvjf
HFWXSHddgjDVXsIApLKDQa+09J704zkswrtP5aQIeiXcKTl9BsBlvK8YGnasbhfE
7L24PO88V88zAR+94GIyyAeBP1G8va0+PaMKdEkuNr9f6916RsCH8tDNhUL3nlB9
y6nCTQpuN7wMCxHcscJMNMEESCt7qpxgEJQsERtp/bsKpSxmQIinP7siVtNreFNT
Kr7GaOFrBXSreNfUF8nI0HGFxnk4OtJX8xXD5acxF6gwH6L+FnAZ2BT1sRCYiHP5
0s2B9pXfFCGrVnSRdERuqzOto3LsXyQidulA/E4lTnqjQBo504bFfHz2rehPNtb0
sWF/RSK42rA0YXZ4X6TUSwZ/Ydw8Vvvstz5gT+YsF34ogpNOcDmq1QHdYxEFkST3
H6mW93mXOGcvDq3Dy6ZKsxJ/ewueAVjGwaX9OXve5lsB7bpcg7bzJMJjSt0fS35J
8UNJrcweyFKil9j9qeXPF7msVQK4LhVWS1lHVjQgPNhJX1fiIYzyvI4QXWFW9cYF
DmUp4aPvMfKorQhil/rjA4zeRkMQ57keaxg0sXd/E8yz25KPVjYFg1BbqLJkX5yF
W++vr6d7zQf7iSRJRQO3poIsG+8Epo8UX+CFyBH+QJmxnqtqmQQ4SX8qVU77wqTV
X9y7NY5RlSSvSirWds63+zEHxdskaWNXkrxUt1lugXwkbB03TD3b5oxGE2EEiH7d
yOM2i5pJjCoZm+Y8muRdEvK58BeD2lpnw+/JbbUzTCA6g/14emsnoFF5KlRSYyLC
gQ5b1/R7Y/ivbPPenPYeECJX4vpoovcaNqbAH8B4qbEI9nVE0x0gDUMFzH0fLD00
yZeYwtwCxljP/hnh0MadW5QNXIiKJpYVlqDhmqUz0nN5Py71giVUIjYV93QRDPzF
3wmlzBPy0qScDXLiCCdROnN/AuO3UqHuMvaN3UxD+tOT8Mi0eIF1qBMH1xquwYJo
R3QqKjhj8DlKQ9chwMizNLGT1JjwSXMjSL9ZbMudGbS2EkBjfMRXGbCnZv3z7v3+
d7+RQCieLEea2YQNZs/BKT+Zb8+hBwOQGS0XT8t32mVCZx5GYjqYQRd7UeWSvfmM
Gs9gRy6AZfZcgH+sE3F/Eo7M+j8IPv+Ixp7VwnqM/mu0rUPhhfwinb38ExlWj2OZ
q/c11t3wIY0g2HKJJm86cw5X9pbduvXoYHb6HGlNVLIzlQBcDbv8JSZsUUnLotQO
huk1LNlQYKTpnZijGOKN4ZaSiI5hzwoBqU2oSD34xD9PbPMpQpdThvzS4Bab8bBv
qMipix+b3WwVarGHfujtDmq4OFrsIk3PrNrf1c29PbKYa8hWz0PE5LleV8rTm36C
3XLTXXDqOZ0EjpXGrFRF1yrbgGp+/Ca1/0FaFG7tE4Cw33wWzNDVaCerC/k8DfM9
OjwBK8ac29r+6AzuSpu7S2E04VyrjsofmIOC4W3WfWZfXhF39EYTk30sh2ZwUEc5
zx0k3eCP6+2pQVrrx51ZPvWzBnEb+Owt90MTRCd5Db6VMGT8Q9D1bJuXQTEAtJU5
Ai3rnfCrT1Hd7TQRzCOFqXJKxhvZ0O/kveh0D2S9iCTQsHA7kh/YM5XhK6Ym9cbl
RbpArTYr1kD9Z8CUuSJZvZtHW5l7W9kEd+vdSxAMNtM5G/s3qbBUWsyYqilfYUgN
Op/0hVAw+YUW/m7fY7a31HlvSE3z3i1ERcOkzSXAm7dGFgc7iNyM6/gS4QlpnDri
lq6dnPAOeSWsVQEnNp2uGg8/XXsQ3C9a88vd8IhBqv5IZWJnVjnbL7d3C8ETqKWI
JInm/DKZKy53DHULIh5ADdrdGvaSiaMh6uGvuZg1J/JKTYmn3j+1iuuC9175yRJB
Qp3Lp/q5vm8cye1lfWtO/dN2vXOqeFDWZ38HPQDPjNj6c2Gx89ZWywoGirjeiVOY
lCZwBosCLyMinggEIESuBUCrEwdy1q0F5ay4iics3YH9xx5nZ3JTJAecRv1QWlUl
HpBjZ4gZEkUXq0gKytZOHC/rdet9SDyR/cK97GyxfH7eMVth9iVdF2XMrI3vqkwF
dauopeYKOAFAPb3Q0LJbCG+TrM4qk4VLoRbqMknVMNAP8rCiqkGAgC77LvwMsftV
VeI0y3ZR0n7CT1zqo0GWYTslCwuK9q1xaDDsq5xuugzD5PwEgjEM36Xx5D6W4BRM
V5/38y+RgGRT1zK5sh6K6W49ac59nBmEKxTM0tCn37ONcACFvl8LdRimKr7/gDhy
xkfxln1G7CQqoj4pHcTcK1WUFHTsOY0ELJlxTT5EwFzOigOfAJXQxsvraq/voKz7
JFX9IEQXBPvFqnzl887c+2yhWYmdAQoh3e4T+4AFxBwJKBMk7r2Tg8YqoTkqh5Ev
1zU6OqA3XpzQlA6SGRpToiGhAUWX2ZfjixyrTmZmU9CN473Np2DjOuuQzTmxFrN8
eEvRDRQckpjyR7CzicY94eVAboVp1yXFuOUzcDFWAogpXYI4SwzlRGy2la57kLkp
OdNx64Hka6bpBn+DHz3xCCuXBNF78ZMtr+gVo2AQIhHV7ZwdXFdjOTFYflgjpkGT
mLaiI91RusLbp206RD/W9+83scahMDyzDA0urTKw1zxfpYDnQ1/GFDn9y3h+ikQa
m6pvsM6OZrGY4XzdtGAdeWU2D1yL6HmiutYmsk8AiIIy0WhN7ADmdtE9FoVMOMdd
vIBs6Qi4Ki14GINMI+wsfnlJW5FhmasJxfgs74OZLPes0zD/dPKihxqHbM2j2eQ1
DTw5hzb6Z5BO/paehKnVrA7iagYxaT9ruWaTI71dc0DjC2l1Xd6v+kXMVH4iE6Me
u4yTUrAUcFvD+M/ipCkHWxgLuO+VpJjjt6SlYifnR+p4fhwnDZ6Fn/8OZ6cVOERy
ZHeqLsXZCO2lFkcKReyrk2ZHqE6mj9mh4mdmGrBljOVUNd7BOr/Uvvg9kqFC2Jsl
mxLaRuLLKY/FzcAUC0Zjv95zSHnHng7wWMs150gPxPSPm4Z6REaFgK9hAyM7NznH
y0nJrHjiumzdt313+EpbrLcUnWDcIAjOyQnnzVzolMg0YiLD3iBnyugaL+cyw/vm
TOQoeQysb8Xwm97iT9XNE/gq2JemeVVVtk8MK6TbiWyxaCJf8XXKV8mqlW6pu8eD
AzeHF5xJP9padkpEIOyZYuZzJBSPMzZyyk75DXJbfODjQxvFcSF+cJjJ+XLVwk3d
opTLAboSv8eSWXKzeb40Q/9Tc5E4GpfufaOKyEXrNvSDeaIomCqc2JG6qM/a/01R
BOXXeBHX4JXDHl67WbB22N5yr5dIwNP3cOnYoGYiIu8Kuq8HsZDUv0GhasJhmZoZ
zO25lJWuJvP+6ULaIhzulxSXC2ccJNaFuoG7IjcEwbFLZSrXFR/dPHhWlCShvsjm
bSlliQPyHSrxI8mlMY2DmKptUnL8eJtD4ddNdNzgBZdNZpZPkRU72ldSwrafnVj6
5+E6vESD5tr6LqRI2nOGqzcWJAgODxylwsbwWqty6EmI0q1Ypqb1cFFZuPoeDXZJ
9DK3LcY8kM1oz869DbBykFouO/uVHxBRTEyGhT1u0YMH8SnUbakcAyAFh3EsCgi+
inQCKtPeycWuB55uqKtD3nJAjk937L7l/36KSA0yNMJ7OeX6xsyFkblwpHh8zbA1
5b+p2nb7uCajo/doKTjocNLoOKXNJ4QaQ8hW1PFVWlMV78X5mitkVPRKgNORIs1B
ASx23la6FYGG/6u0v21ZiUUBBHM78uCxvmQ+8spgoYdreuwubCOkPP/joK9JW0UR
3Br1H0zB8jqMUNCeL4d5fUKvi/wGY9NbTvSgVBERhG3DKQSzgBk4UfgYheK3V053
5uYGISLVU2Jx62WFohS4BGyoKoRVmrTSvFAEyM8w883IyDlsHuwEYqAlPQtvAnP8
SOKSWIHooEOmunroBqpfP683HBEYXlup6ZUugJSOPFWCs34t7FKynRK0AoKnpNpW
GPtHZPwu429MgcpNBuPEg0hb5LOM9hmVIiSGpWEYcI5CuG/r8nv3PQYAvhPJHZyY
U5T1a5nqQRJpqkSqGHOM06FemCT+3Yv4oE02PSXZeNcZmhNe+mv048CVyZo9GtKP
Tr2qxPdF6aZ73fzabF4J8omKRL25zoFDWuJ2vASWvAYDPkwFH820YPYW3uDsMJep
pMeq1zzcdW0KmDpfNimPvUkE69+xB/V2A16roK0hyFZqXeqWRRVyxlMV4nH/Jc+L
Uih4rd7hsQCq7dgRL9lMWwF8hc0g8PX5te/VvngH8YlQhE/Mlgi4xg55FMTBB2UP
H/i3zAm3fiMqBdI/hNNN5Vax5DMEMzXoKjIWLH77YJHxnhWauSV4WuFLKhvvFOsK
WziP68hvAS+Atet+7avtANzyTLm2dMx1hwVzP7vkZsg56RkICuy2KOZrVz66WEhz
5qDJSsTQvmOWjaIm9vvNpJ1B2DFxRVoMNKLhceFKgmq8+ufjPnIK7ETzdDYWPiIK
LZsBZMHdRultJNZjK3J2GRcDkw/oAuKKiurKsPqv9D8X5uqDYj/R7Xv0Bq8CGaGO
VWQbjJOH7hdzljVUcdM9lpOJazzZCvdtfHuNGfKGhizeRVC6DeuzxxAZy+fK0fs4
zruLliYZDTDNTw+reUdf45ibdovlhwpvm6a3BaWnnj+H1sDbLd2Wd93q38iKo3XK
z21LmzTkQ9ALRnAouwOogl4vetWNsUPmQwy4oDolFPWuT8sY7BiTKIBt4UrpqkZF
4x66yGnexk6kL8PWZJv5ucx2EYbLFYCZYWHgGExbRqEUYA7KXiAzjftLnXHIJZbN
spvR8IgJad6sNUSQPjaOjhcDXej9Oy4NSUmYydzxxv9JPJAtf8oNVQXTdhWSUXf/
Nc4BfZ2mS5UwjC9c7x9xTd+VfZT4+YROn8+PZG0QEz4CFfcsSyQW8F7/glXWxhqo
+J9FXbPQEsY1LMu3WtjvOPpFHKwG29MM6i77gngRaHK8oJ/J5DcyI111FzSvOyZ+
qWcVR29tx+4V3rNQ/bXzS0hRfJ5Luj5oXqxN7yd29ksBNh3wG4KJbm0mCHb/S+6A
xXiOLXW7O7nnelj1Tx51u0faQht+oxkTC7kR8TyYNjv1Fgn0zUz5/4NH8xiIrbik
F2wrUfzgfrCibj8BpV5FckFv/YVQl7e6+KJAi0mwXY9+PZ1Z5E/DFpoKPGd45+B1
LzRv5xBtek5laaPwhu9HxHMbaMhScOnn9Yf4M0zPkbUugPjU2yK8tgxssOU0SSiE
ZGBDJRcuYXwww1zXtBrxO58a8hYRauqu2gVSQz47XBohmKnslrIbm9gzq5N6bFyY
ttPcN/WS/7wWy13P6sL157NO6csnEoM0Zb7hvO8Uqpr0aWTgt86yuUUff/vTonjI
28NZguyNYIZl7QjBX9f3ATJgRIL6MKJgyyXchFQnSADlK85VJWouLg1ipEWEqh3M
1HeetsYRa40IJajiv37el8SO0p7gRDDw4gbCfRaXYurJocG1UzaWgJARzw6q6Mb9
q5GdIbZ4APz0dyWQNDkRMt1vpXAORD3Ej1DTD/HufhNLnEmqq2Om3UuuVy3Q2Ww3
cwYyf3AqIne2W63jPGuBHqNEi5vFvjmBT+3FKHyD0eP6o63E6WS0QjgwMEOYQV5B
EZFp/LqJUASXMdOqq02YptWgtDwMnectqSePR9C28Lynf4D9Zcidi5SRJ77+YGfu
6Ukm6rzSv28VYpwBYZUHSYbRiSipeCsFDNJyoV5b22pNkxMPY8pEAkTvwJ1OghNu
KOrzXEjwnkQB2qP4OwPjBUa0fNBi35RcnPUfMRuYphQYoeqN6KKRbmCyfe7gAwyN
Wguy5tUfSb0f8d3+wKz/8IJUIwtRX3ZqRKJV9/L0gFiKhEcLkpc+vBDSYUt4jNtu
hJgJrHRSBKo3bKqFgl+qTUdccHNOCQ9DsdmJDHFFBn3zmOHO+adAJt7yQcQACkEW
Qgs+vIuA3oulXh+k5Y6bsF4nIzStx8UCue6SrYkS2nHKfuvnVfIgCYIEuywgwnCL
gth6yzNNpNvnHchpfPzEg2uGjGbhdcgWf0J7K7egaYgf6afIhrlixYB/Nr3+GEB0
Vv5wH04vh03GyC8DYLHSZp+AD3MGhmwi1R6l4n9y2NKbtEgZee/lIqL2EsQ2rpB1
KAUJheWXmQ0ola4M0kI1a8i3Bz0RgDvTY2grNIUBBiHtzRUalLLOvSz1nckzX2Vn
EOirTXs+fmn+Rw3wHwj7biIhgzp9BIyZEKYsE7Q979flJlwHbTLAqmpcraYUzHNq
eAWZHUGrUoqGoHWZLFr4ET1AUYbQy6ebWTN65C+IHhthN0XgTBQ3P9N7Z2EMXfgU
vAGIhNPSAHV3mLnnKUUSy++OtAYTuZVHaMVDerG1hNdMVYX4dQm5Kvf54JD9GWSx
3avGCdgvF27Trm2BLJ7aC2SxqS9AAo2Gy+JKQoy3vT3PSJAyVmwW6F+JbfsaQ9af
eDXImmX/K+aW2iS6UXp2soQF0qC6o/twmrV+DdIPN4S+8Sn9pp3dok0DH5145jlr
UmN9viN34MkgYfLO34vEQRg+B/DhpeynSFlNsCfFx/vYghndOPVXfnTwF2AFKJea
xbZAniryKh1BD7yB3g3hTACSLECdd65pchpkF9SfgEsBnW9fJGuTb6MmNfgWmlCr
h1gQnMdLdjOlXUdySUg8V3hM6bkBy/cAVk3agU38/Yrb+HeGuerkRhg2HnGl+lu0
8spuS3lqq3P/RMtuI8sMvV4AwSGur1Lot18ZemmY2nLjXlBnxiCxi8dTWnYkGPBt
RgA9Sj7kG5b7EIecOxfJDtr2RNaPLIAi8LTpyidiZEj8ceFktVe+SYdqRk63vsAv
E0FJ8lg1Da6bepV+bXOmuWu7q9jRRP5LGSERUlZUD7ejlr3jYZ8oqwqBbf6DWBn6
jAudQLk4jmQHSR5HwnB4sTExhk0IYPWPrgs6mn7YSVElWVXKDmVPX0MS+3GaDCKX
uY9qisWDNkaJ9rAwy5ygVCqSUsSHvfb78mHgjBxBBLy+WuSNS2cxV/R1NutawMGD
GL8tbaPoATx/+1FyZE/ay36S0t68iG4LLc3Wwsdb3S0t1AyeTrViD3T1504+M1En
Jq43oEbRBykUH90bPfNhaZRQkkP9J3OzK/qVfxjF6BQeikIk0c/2yBj9WJUMouc7
JBHV4+nRPC5L6W+OpmVJ1qo2aAUdQGGxSiSwMpufSktfxGnl2Dn4nCUH9Rz0n554
Hwaff2/r5eMVh5m1WAmyDMbRdSJh+NH/BHHoIymWVSU7oeFneu0okuNhkBSdVcFQ
NxWwxgemMxcZ7dQjA8yuqAAssn+dN/pNBSfOFKYwlGMvatn4oq6XpCiYEkInCuUI
qki8sa+j+xA/T54ohhAuuU/vTGNBLQ02ruftKqPOthmhj6Fqj1Dddr3CsIWDh+j6
AWytryEM82smU6Q2jdpRYjXp0ZbihIx8gljqQqYFDNt+IGbUHuAYpeGL9OKwbsO3
k9NyB0KkIIEsARx1wksuguFQRwXTPVxvLg2LmLJAXLYlMgE0v6CeoZMTUg0O4rCS
tOnuJnd1cVUpPDpb/kKDdLwx5RmjkkaTbNyMkkFSD+2xr68cXGrawtkk/ukwkq78
TwMG8Pmu8ZIVUyHuZ1y2mC0mfnKfBWMyoG28ymPNo8RTC3lj2AHlwC5ml6Ys6PgW
EdSRF2H1Fb0S/KESWjHWdnsrv633p1uIOIGQ8DBIJS+pd1hZhwe8l8FjIj/wDg4X
yt96UqQXZP9mpvJ5kTatQtp4sWbyleJeNGxVLlsMECqMXVnWai3FGEe5YsZ53ICt
9bpKYZ/8vqpcnvvDdTA8UFI/nKmNMV4VwYqARMEjl4+TnLVlNOm3n2Yxvt84Gy8u
ZubgLot4s2pSGg3IwMvVoz873EqRE+cTldunhHNHh4b3+8FgZKqVqANnzPTk3mM2
63adUATrWB9xY8+T2ZpOFaXygi8JuyJ48astsrqvsxsunxCkxFuXueG+4sejhBrh
ehKvQ/Gxyy+7ao6oVso+a7MswdHPUQNbTnwKdAK/4ALL5uRMBlLcnBQUuzwMcMtv
wBmhRN6urknrmOqdnjgkrDBHhNAgWT8fuFWvRA68s/ubn3VtvrlfTz18h9BaTArb
FHwi6D0FlCRQIelUGPLqcfpeBvH1toyDRirh13BEghYymRC2k7sOJ32QBKqtSGXM
7CrBjtqotqjujpA24Z4IENXElc92hqTUj0TZ7nSX+9vSGLL5Vogf0orWQMzGnLlI
h43SgiPQSpjnEmes8MdJ/HQ63HnQ3fsW+4LOnPhMa/cTL+0ufHFrdoEhQKLHCZra
m1ylCvSniC0A6FYsPaXS19Ko5Em2HVlEVCu6scqsz/8tVWSlOO3NK5yFGzkI7Qtm
YTmJ1FZIbB4uQmJbej446XWSEfdKhTDFPHdC4LawMeBXBjLe/pOaXksThnu0B7Ut
2NQhcOYetiuBt0KO35nu2QdvQrF6EF9A12429HJSmfD8kSc3elK6cblfPed/7X7N
6H5BrUOQjoT3ChYn7xOthpJcQtOOWp+tK0EStt81cDVlJcsjw1Jt/4x8wndbHa4N
S+wBHoPT7jH25ai7Klo3Rg2ZJJmSI4jRERffVnH9duLbScmaF4EpGNfoNb11e3K2
kyPuMxWJn0Q6V8zpx61ytzpYQJvkT5mKw/+7bAF5fY301P4vR2PpQ+WzUC3MeFyR
cvkWIZeNgdRoNomnvLLKdvHn/bhJ7t5J5QUVDhbVFzks5l6xMQLg4oFRPJ9A5TQX
K4UX3GOXALsDktybBKs4Hu3RhXocUDV7cOeoQEQO37Gb5V1d4MmxFMMVEu84qtaf
d5lhKolzb6vyGfPmwtTPp2mRKNsPQSAWO0G6wVAexpx+WnZ0nQUm9S5J1xAkszt1
SgLrrOq4fFlYk4Yks8L10H1l8TU2oQxR3zL+/YnhE/DM5qZwuZivIhvxGt8AG9nZ
t78DkiRJC8DpYaS7h3W11ytL11lIh8wjpwyz7ijyrF+Vq2ZPLe33QvAVkK55C2vJ
+YP3FfnDY48KRua2y6RWkWuoRTvsn0K4zgJjJNC6UrGO30EpgeWE/kwiwdWqSViI
poJzqLd+uMnNOSwhwtacx3R6SG9HUQL7d1hDvOemnPAKDryUCGHZtELDE82kMb8J
vIMcquklHBRfirTrOjANc8ULt/4P1M6a2VoHG3HVSK8St38/eEojzwYQqvftn8/V
FcnhnaUj0R6ww7JGV0MfXYqnb+Y78w0geNXCGfD02zKRem8Qbk7R39jhRalP3KRD
EMRcAtx2Dqnhikx+XzBWY3vksnGkU6FeW0cqdraIGaiZwmbdn5SopvKvINIvzlOJ
pGVWmDgSHIaOIgIUhKpJmnRirK8Xghu0Ffc+fezjC/iGz8oe99xW+vGQKqVuDTuo
hh7T7Wsn1kUBFpRCJ8Bu9d4QoUn9ys+OejdjCU80blA6UT7Eio0N6KG/VcHc0FGs
rVn9RsO46OlCmkDMUOBIYyjsr2NLGzBA/6EJtJkgYNhlnRWfOKvlATWXhJaEmd8X
R9zMz0NM0eUdGF9Ko9VO/5NkbreJBAjYOBfpPcCoRQVcaNNsU5SMhaAYzWD6TsB4
jLG7WXd+MlspfY2ygA4sGduhkJbxrfrQtJ+mlUKw+vty+20/KJzhPainic8Lqx7v
z9e+yf28kqxsQSMkbZnOZF12LW62Av0xwy/K4eWZZapZJP1dY973o2gGgAoraIRc
NJNO6ICXeplaW4IvD8aE3ErmH5ESWNohNg8VeYGcZRPQLudKiFC1WSi6TsWNYY3b
zPECxe0GZAfCE+NhQSe6Tux63rd7br5vRgIIwQpmFLDPUaLj/xq3iYrR+04SRr9t
2k6IT8c4GOX8c3HOqBozYJbpAsqHUeAeJ8N4pQpqGKLTTkdj6H4zwruMXDFnC8OK
c4nyIdoezCoQGPpC+tP9g4I/RrqEYRNWrtiesUMElNOdauEmrolmvCYV0NUEGz37
I32nse1/34Aghq0MICml7XCKclDwYQJoYOCIMfx2TGYJCU7yoNqR9dwLU6Td07wT
hOxj4pNWmDHtSVdOxmTz/zlx+2BPd+STM2okJ7R2zy/YqcWoKgCtVhAh/dlhwNXp
/G5b+4B/iSZkVFH5MvyN1/4Ztddt1AIp+rgElUbekn+c70YwdhKFWbMBUI+O2t4X
MKnq+gYaTh850XkbFdjvvyrWiXM1x0TPh47Zvc+yWXixaBk6KWYCHR6VRQ7bO3Z2
KpGhakBa+O46pMFYxvnKajeuoUb02fDUHzgG66S8VEuVVGZ/3Uq6fbsM+SlkQw19
/2J/5zAviebGFWmaXOUBnNc6KnipAci0UsZpUYd1tEwo9FPNeHuKoWkQJAOhTMXx
jcBJAwBJKIvONQk3vo7aOg8qFH3Ybz5pvD+nfTFU3u34V21nD3AEzVy3gLhGd6qI
yZmgXVE22nCHbwaw6HJB1Wiv+a3o6bSsrVvobj8Ls6D9tShnelHyFAbRcp73bEm9
o9/pSTyWTqR+kAKRRzx+rNcEzR74wjFcrCFHxAWNEIW2uYOoO93m663w2+jPaaR0
TtAVINix2cAn6T+xH/n8rYqk1xMlDbqVsJLE9H/4PRc7nLfXolwKnXh140jfQdrL
yN4i91Do4mgLSHojBv5VmcfT9PsqifOqgpm1zJtQI2+Sgwd9nRXKGFrvDbB6sBZG
uulHbZdz1GnicpxmYJUFDY7lvIYo1Qfhd7hRxKrmT2wXsCVka5HFUvhxax+v1mh7
Psmogs4/7QCX5lccWXLhB8n3w6jJKQ7MT8Z3jiCz/ZHNujsponcV9Lb17Rdlgp4g
ofN0w8kdlAxJyBpRcnDmxZYsyvoD1EpCjza5jY/PH4VOTUnjE80X2uU38+rh4i+C
X3g5ja+1GvxEmXHineJvPp3nbVnoFFdkDvdvyXzRoAcitgPM1tTmaPYUS7vdWr1h
q9jKQw/KiI4T8cUwGCd2MLhiXSNSjsq2b12UzdM+16wCLR2cCum9DjBjEKxm1I3C
fSmfeIpXdgDDHuEVfMScbr989jkIFoiYcKBGqHgrFWsY1VBSAGeef+WnaEzKcZFI
R5MQRaLJZXjSSMjgjMWMmqh8ZiYrR6AJI5+C4Bk4DK4FQXWZV/Z/dBNj0y/WTqrW
HU5Xeci/Xe5iMTSYbQa3l7UbQyji0r7C9+3j+z66GEjEcwZuJttch+Gzs0DRipj1
txyhyeZWl0PdHFobEP6LyYYdOjcAx28llJpu5Ycs/yXEkSaplxxqO/XeTp/9R/Zt
3BaCDLf0JvUig5E4zXSeH6D7Rz8u0xHp/TJlEbQv0waGaul6QVI7thoXAc0AN8Fv
gyR5qKYDWGZVGRracOoEnD++DaY9fcq/o5nG3S69MkIXg0VbU+M8bmThB/k5cVPJ
ag4XUAylQDguovMc+y6jEnQCMmURYdXYLbC75PN7V0ZHCuoP6Euw/GBYI4QnPy4f
/R1ibqWwhfySGxkABEFCMvEbzz28SdnmpFapf2D2NdgVxNKV5f3xcsp4PXSqGJ7V
A4GhFk6uOb0n+zDA5PhGHVwTktxl84qm3Wlc5be8Kqm3GGJitVoPk0Goxm1c1tHQ
714I0YNK26ItYc5iwzDkJt9a0y9pHElmUYFX/4EUVJedYDBjDsFbdJyirRCQQP0x
Q4Egv1MY0FumA4BMbbFGnkVIZR/emrtmkgwN/lbJWmzjgdtsMO0s4Z6CG3d3sS0B
lTikW0NyL1tOVIFKxXpx6QtMkqjWKOfRnK71e4OfM5BXRrElMMs2NtJv8C6N5V0Z
MOARL0Sw+dYNTJ/CveFxHGEags+wtesE6Du2y/yKgLYoRReJfbnZNKFlcEfS9cEX
FmIOhkc5JSBBT+C/ky9ry8Ec0nONmKrDeIPj2LRWOFM0LHPRuDvLcyUZwYnUqgA4
YVXEXXV54Uio95RtAl5H/OBdgjeiWk0JAUKIQvD+hngCuknsh8G9GEKyzDnA4uKp
iC190DH9YwTK7OLZslvAN6iAQH6R4Ri52Z1v+VlNJMgzWO5D0DSgU2ZNJ66yZYQ2
GWgCaYTX0W1FtMjgOWu73o9CAofTSo+kJqOl0Xbrs+4ITWvyHbX6DmvLVxCk7yDi
GVBw/OOeQzG1ElAR544hmn6Fh2aeCEaIc+866K5L0Wqz82soFm1uxA63UrWNyrSq
uQaPC7no4CPMDl6nbiHZtHuClUGQE2lzCTpGSnr2W57qHG8LAGvFz2R3IXbRyAKN
FMvgTYNjzEUyeY9EOVS22q+PY5MbcCLDvy84gnor4DkMVTrFQF8QHjif2GyCMaSX
Avl9OQ7vyHZbZ3PTFdF/Ro+X+FRdctV/hvxWrX6RinFcBk+e7Ycy9KfbU7LmFTS7
wwqQ+GpeWMjv7bXn5RT9DhfuZnyDLvs2oJBcW4iyu0NIz4ZtKOm6DuDRQL7Uu8FA
DQXNdXh5R9BZTnL0iVcn3q5pacUy1gisT6FiY0ToC9azaXzNo9/AiyI3pTNRRb+B
hiq3VVi9ktQ+cS2HAzso8zXjIzDkNWGhV5ixALT5jjrAKWgWZsDD4Fu/eGeTbAlz
ThFxMmH7oBQiOHmVvxcMXgCC4yHk9fmdfTxSqyDQ4T3Ao2Ijh7PP95ZS4EkM+ZzZ
COybB4VI8aQGQ/MwB8ciH3uqqMPC4ifEgul5IZLPRzrqHqXJIj47Fy7oEaW3yNye
WWh+L3vQng+JjQV4LNiZbv7GF/64QL7k1zHgEBP/uz1EsDVcrddQLUefGPZ/1X9Z
0dRqCZBOD72MZeNfvKbDU6NRrmxWMhx1oS0I0MOqpQqu9XNlB/gFaSgFnSSWEtW8
BXvDiBR7X1OTjyrUmCe3hTVIZ5/M8GVDkrwAddarrl29oqY51xOjujG+wY8UOK9H
kmiqkfxFQu822DB/MhntJGEzTCpJQ4L/0ddcUzyi99hE5h77xFbWUUHoYbEXq6f7
lsDTzYJs2jVyNU38jcU9o0f35h7diGq45LNCAWa4yHEmL3sm8KKL+pK5hmaSDIAp
EzMFNALBdOpbu+bhSiJQglSHDf67oz36nqs8a7DgBR0Bs84WQqf2TZGoJXkIp0ni
3Xsv1dSyqcpHaGRK54oQ3M1guNuBuDj6Jb3SzkbMPOp1LrIIgCBR6wIDliaRMpRR
z/doutrHZLqsY2feQ4GIqDUviQcoPzgp31JlpakuvH/WLbojsE3d+BisKCWDqEyr
vUJorfFOL+5wxNDXWYM+ASFGIa9eaY5N1AeRIKSti15zQEkbW1H8SQxD0PZEy9uq
HG/yrnpzcJzCrmK3EbCfKw7XYRJMCatnFxlsqz34UfWoNWMBv43PzXkZ6P/g+G6y
bb6nRaZSMKmaRMj36v5zVMq/DU1XrCDcar99W0LUoVCszxucsQPttQrAk+heLUFq
vxZpHC4C8AgkrJdyeng+I1oKDbKULJbnezy3UP8es3zaeudd6X93h5fjMNiFUesj
zwFaHFxt0Eqm6ZTYMIp/TjRigmP1Um3nyJCw54g8+weJgro7ZUo3eg0qgNeCEnWM
sj9I0gPTkXuXv8WMKRS6fLIHIq1RvlGHb9l8SW8zkRwRpOIJNkwaOZw/oTa96Xta
mLFzTA4jV6ZAcldfEzDQZVYRJX9tHXfyauY+v9ZXRqX/8Vm0KDBhTKWSir2dEjtg
9Xmjj/RY0+XUh9enNJhqx/Z7s5M7Oq3G5u4TiXezMCYfHoR/HfmHO2YqPG9xCVzi
Ll8gOWg4NwiUHeR2pl5XfE/TYSM17R/LZcVYeqAKRAc7gWF4sc/vBtwvs4vFRBiM
XfAaL9KenFtlemU2xT6KiPsdmhApJFX+grF/693XATukXioDQoe3HooFIAGqDNfe
o8tmqkVvUrYhOr43oHsmVeqwTiXQEk8NSOmdxEnzV8SYBHQOIbkKeQXsyoQkIphB
/Nigp7OFDVucfrOao8/4mf75qKHGCHfHYuqdM7WyzfX9LLwidA143PlYdkwK18SI
+evXFFMhrCKlB75kLz6Ppl2zW3hHIKHdA6kicYQFIj23+YeBdV1YYvM1oB+66nLZ
Nf1s74bRJYNiRNYMH8tEMRS6DG6EJaRkoLUKEjFai9aXn/gs8XNI2h14XHzVCJTV
JUXZOgqSfHkDWg8b0uTsxGdg70aYwXJMKZDz8+qNhy02cMAxzetOXrVOieUB3IU1
rZTb+UnBtONRJVd4piaz1VsO41liyhUlXMSQ1/IZSKG59WfQhzMMh9fkBZWRsu9/
XFVhemtnz8QtbrAdjqpACSTeLRaYuj9ES6pq2Ynz1/40DYK+DN1d32DhiIj5LX7x
RMR6uJ+w4mcb3EOHz23Bj81wfmNQURQPYha+jj2eJjCSJ72Yi1fYRE83LxaNYwzQ
m+oW2n4315ontsRGP6+A8IMa7taO45IACjNfjpURto4Zw31DFC4PuPwVZ2oGHmYB
aSEfW64eG/6iVBzXVzfT5Xy5S9HGPQ4sivcxwUwI/covJpkeb0kRkJA/ClDCNbeR
yR7FID2WA/A/Ar9YUa3t/ZZlixPyb7998Y8rEaolvrIgDMqIcsnBWg/fxv0BEOhO
6nzhlcrPNXOdibWp4+G/Jk31U8kSpDptAp1uDIQGo3rGLn2gTsrdzoBONW9424oR
lgU8tIML5fnDoxwNh4BKy0Sio0cDR8gwRZL8N5bPy986Z0jMGUmMPwwkXbjALpdX
bmHhzhPH/sloEFn9hZBE3rXRG2axLz9qN2UoJdRZiW11ivMNXoqNtbf10P3cJBkX
LMiltZW6OeUZufC4N9iJK6tqXIsY5q3yJLzmGMLn2gnAFB0q5yCdwu/MS6xpjmXf
0A/GOEjLzoqI7owN01NNRs9bxGcyaL4Zt54FPFXaKBbj3vzcvAqn0NZSbrGcxvDL
su3R+g0YcSSn5S2892yN+A+GMeYGKvOzHlBFQK/JT4mRpP1Ufk+y4Q77rfPiNXbA
9oOQjxABN6Uyp/Sn5+nE9nSfI6R9Dx667tkJrPfEGXogORUBhutVZbQaVNDDHG4o
pGyOht/EHeNHhBmC8SD7NctlH3l7cCE5/Qzmx2iqFTd4eAZ5k9sa9mRHX4B/btnK
/0+GVx55MEieby6Y6KXQsvPkty6Zt31ZPT+OxHfzzHB0KmUvzMplO64EFSRNGrJs
VqPAudkW1Tmx53u8LiIdrlPej5IT+Cdj0km+zRwc/BeL1rWPW1jDsJwsY0OK9YrN
58Xc/PVuDZ9zIFvM974MxQsy1r+H486ec/XAD9viQg3jjFv8rzY+NlzqHuPqlFjM
YvUxz9+vlVSxX++r0dh0/bc5K6LmcjUOJsL4z8DiAyy2Tl4azhmXVl0Tu9Pj/01N
0HIVqg0YLEj6Yy8ZaxR9/TIPI2vkEoek0ljtUYm0tTl7dejeQLPZymnl/KatDRTT
xoUTyKvFE8/yDg6bBSbJDi0XfyUckQw0HNGZ7dxlxlsdF6J4m5Wqe6ljZp8n7JS5
NCplCxT6kBxxX5ZjzFkGWw6gZBXwQvsELDzGJ9ftxxiP2r1eQFBdYv60NYZZ3soh
xRtwcctnL2TCJvumMyZ5EiP8WTh8PLe8Sm1PwlWqPgKVLEeT/GkIpRI23BQbXTtZ
gMEZKi6TJAa4yABWsvF/0Z7iPgSyVWPAa5kJyPvIU+BzpPqYfO3xJDMWwn188PzM
QnYJsGMJC4QU6CuHYn+aKQFqbM1QGc0l6ce+FMVPHa4rBIRlLMQgjVMDLDy7uQJh
2CDrTOC3huTOI58tH4zQ5/wLoh9CsslUZ7Wxu7orSE3zRoFPd2Yop4S8UuUzGr1/
Mh71CjSy01HN7UnSayoViHmv79e85mfXPcRizfD6Y/9zYPlQLCqSTmXnTisdzbrH
hjftMUtMiAFUGjU6/8eE7AxiRe11S1lAgyvWGNtzDZDTRp1wUdJPYIzEFWofWE0W
aSAIqEXNd1c5F58q3c+DmWwUg2qGNS0p3cCKwOVSlyHyzjsL87rRx2/Lm4zyeqVh
NiDmerNXZU2vlgYQkHipp+hLD01yi8e8bz45RMdBcD1nw8MYnubum1WPoYljMJq3
dR4oD/UkIZKOTOGGJjf2l3VNqnLDKXuKWPlUwVP5IJSSNgSJwZ09BxHUGkAacb5a
guRpieSmEsSRYC8dT3i8DRry6uOLo7eYXccsVSLEqzxu76wTqxHwnE9mqv21tHYZ
ihp7guNa16oJYqyCrVC5/HmIXJroSzKBE+croVR2faAZyb5TFAlvQzjygsm0vxnt
yQ6uIOqwyjvb9B1Z2v4yeCgf5FZrpWoH/h6py+wq4lHpuxoZePNOc5Uu7AtVfUOj
k9jcwHwvoYhs/RO8eeb0Yl2eYkABaIVTqjlaHCkALOWoCbvyT6IUVwnz6d2Hdgrw
GOwnQwUJLCEsKRgw4g4GfjRFOc22CzANwD5RQjkmqVGhn0sMXtyNzo3rwrM9wED7
jCB9H4jogJai9T1e+UFw2pG5RYTuwSnWB4WGKdT3K2Fxvq8G6CDO3fd4PztCkKVf
Sr3B5ibF0ZdqSwWwocQ+caNNAtZcQBRGiSEh6K4mT7UJTX527qyoPpt6GdGlIXgy
NcN0x5YBXGXc8SM3U0RaXvnMb7f53WoOyIHwILarUqNiiNh1QqLKg+n5Nrgb4c6m
kYy4z+6cWgTactLiZZ5qfUWNNdbCH/Q51WZsOEBrBpTfrCH8iAaEN+VYSJSwQa8M
soaZtCSNcP76pui2UuPm22n3OliLdFfXWpU+8r31FY1KId5cC1ti2FtUn+msny7K
tieatnXQxdRxxm+tM7KfRrA+q3ma0/z0go3ZIY5IihwXN2Fxx7HaaEU1undM9id0
tz3XoyBlQzI6wiDBxIOs6+HMJCNC8AXNcVvUxv8u3HUFNTT9sCmRL6nrUkBw0fSa
fYvU+lZZAWcCNOY+dD/8/sLkpt0paQ+7HZBMMzGsKCXoqdXWHm3TFz9x3Ja68Lhl
5KLlWhwm8UBhE7KMEfyRO5o6FhbKrtuiC+PS8gPVTb9oMwOCc872hLjQVe3X1438
HbiyZFAY/6ZWIeXs16qwX7kC+kOIu6Xwm4tAj9WSxOT5Z4d7oUrVf3qGjdVlmBlZ
ZdroHjY65wDssRmNh2MaRCjJdHM8N5gUur/B1fQvK++cXSVOPmxaS8MVmqKpxFws
eoHH+yTEtf1D7gU4//u3HLoLiEoMhqe49O/DTjQ1CsIAfRwqclNeuZ7wcZO4hlL8
OyrFXTC1Wbg7VNVVawCMlIWT/yNwciMA2a09LEQboj7IY/L2mRZrRvSPsy3+ZL8p
IDKh1bf1Rhp1j7C4w1EKHHQBtxjBYnxyzJ89qL0LlojVSrTl1Ntzc/yljg4tuteH
1DtgmYE8CQeAGEmTudu9Pe6IrCE+rnhDXd7pDySScYjhnGmF8ozh/E+EkDOLL5XD
ZQ38oHgp08qaYTB5VlQgyQrWqSA2IbhYjqS4g3VHnwvdkV04A3aRygdb6jbUcHNP
L/fkl0STdHKccog4BOKuAnM6BFkdVVusww6b9GIz1t0XYnpA81BTncraqWDi4BvS
EQ1ZiFSBkfKXlXeHphIENKQozmzkYI+o3PViAqJ6jmq9zXGv7Fz7lChNjGDA98f7
Hyd856ZZScY7BiOrXsWpTOHcmJWxSfvQ3tbnZpxjFkiAGFU8e8MOhhUJSDIlhweR
ru4nLqrev0UF1awRVq+ghddVLwhXl+dxNdvs0s55HQJLSrgho54/MgcAzxY3gGve
HfbLIyfRCIusvh52qFG0N9ONZp1Y9Xz7kKaJZ6YMYxPr7vR55jAwX8jlB7PVneKv
FMujIyQK1dSIe2kt9ji9YEH7jkky3BaVBh0x1b+LpjjT65d3GUEPpr6nwqr96xu3
H2xb9ladlYMeZXvAocrG3eyz3zYx+kCrvJ3YGBd5yY1t2odPbsrsBoJjlySSUdcw
A8URiRfUaSUFgO4d67zmYBa2IH4dW50il1c2c8andxv+RNHtsyS1cEhzZBSydgYS
jKEXJimsogPp9gidp1Od7wZFIdCMZxOFTPhLtLYFZHA6bZzvDm+aR9WKinPoCQCf
NI4UfD7dTIvAFBlRiV3ZItWKtkeocBeVwfaF1nNJgcyaOqX5HND7POYqz3ZSIs9T
nN3lDJSp2Y1g91N3oqnBtf9ra5Wvo4SiQZa/hZpiLF70AB1YW60weClzjDxacX6R
XutWHMSrOUWb/Ry1PhdBEBRaPKYVrpQLitmIzANopCMeh6leypjjw6OR8QK2DXTa
LtMV/Czhhx1PJFwnn02BQ2962QddnGliiKBf6uhTOwalBVuS51W5LI30gaDRKqPT
K7bB0nUzNk505RCnygwCoLabO/a91PAxaHPMKeAm77+CHwSe+IGq8mVqPbb/Y8Ht
ukVoyU9vhJ8zT6HK7VWzPRYZAGIm39iTde7rIzkiCvGzFNxTuCgfDRpZ7GZCSQYJ
z7mIbnPFnuskIReIkifFagN89xC1bvjU8NW/0Ivv3sVzyRlz06uRzitx1OCQtwoX
o2sqCFrlqNGCHY7lcYIzvVbe6h9+g7c5t3wu3y6FY4slZ7kU7qkrjcGt9Y5Jltx8
3R/6THVEu0bb0NfeRVLS1XUV0EhBWXT/biMr0P0SrJWbztbnQ1ALL4JRPxDpeyEA
TFqcMTx8CK/OsFR5ilGW1CkZcqOaCVIXefoZyRIDY1QYjKwaLGdzEiJ7pdsu5/NJ
CvqAB06YcjBXzilRwF33Q5cMptdAI+5EiGLlvxENtBEofYXSau67oKbQVgr8hncf
9DEcJs00pFZElrx5dMYXKmzau4LVru1nGKEQ+jktcztfuZxnqvHMl2hgrjGU2ZVV
3eBgpxefO5IIZyzP0auiiRPOTjPg8jOhsex10Xq0R79PUxaF/6GN89OKeoV5K1Pg
5wCDN1+KMW3m3Tr2umWkiMGuk+vfLTNDAu9vBBxGwUOwDVlvTr07xigCpugrhD6V
+6K0J2tAunF1k7wjf29ZPFFfkGTqE0sBOnUm8nZQlPImeBx56RDPWdGlUfLh2jZ1
Cmt+Mq74wSW1kgZ7nEnAOJQDH3hOyjW4D9q01ba3vfCbmHYqqxCDFmKPCGMT9DH7
Q1MXKw/OS+FW97KlK5HGo/v1ywVJ7dKLHmmVi4+lW5MgsCXHQaz7MBjLKr/aBuoY
zLw7+jow5JYIkZcnxeK+N4z9HLhIyMyiLspHIzKwdxRMVqh0Hv+9G3fbV5ayHcuf
HJ5XR6dNd6JvrFX44vsxwS9TV6YnAexxSyIqM2DJY0G5f4crZH0t7f33fwSXel8b
SkK1EYFQj1Wcj0W95M6krxQ43pTSp5lDCVlewi2gw3Ahaf99ZeevgN9OZ+TecfKu
V34qeg3RLSDuYp3GwxoNp/Xf3CTfWgOpx/tOqrV0qLprSrhme3P99vZhi1cQ+dG/
JwRID24pwEQOEneSHFMEw/zRDLbCHbqckbqCWGvwRSeQwyFOTaArKCHkjjb02Bd6
`pragma protect end_protected
