// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 14:01:33 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
nS5ct+xgBVVhkmkR6hIZfbajavrvMD1NQqxUtFvikup0Bv+jvzcDPrdBQ/yWsqph
1GzXRROUslaCOHCzwf/WaBDjQe7q35kB1hvi/KTCWj8H2bQIXJnpAeqXuOVCVM5h
DUJHqyaUd4u27R9uVCx8o+bLdJaY/Y5EASZkeE1c1ro=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7568)
8V7yKNmTTUrGeViLDp9zwhvA9K7jVqa2trDM9HY1+0pMS3QKZMxuGg9FqLTDwN1T
rnnovoN602I5hMFI1TrWJsXtJIvQlUMeQbaU0mHbNqVpp0OgUNQC0OvUhAisnbDm
lKJyzplkQBnT70XlkZT009zLAd8Cwk/EqPpsLg4l6shSICeSwBy0s1VY1IyUPsOZ
2CtiLcyJFgmmqbCTzQzRhv8RvTDcsd0a0buK8CbLfSplQ6cg3FiZFlIluKkNFX/R
s7CUQtBM0vh1HZejfnrnwggDPJi0CoM9b2xQ6ThCT43yJL7fnKAeufEO0qtQQ0pY
SByef0GMryJ2pZy44eCb9aEZZM70bB1kpny37trCQHStcghx2zHCRsf2srpd7P2e
tu+8QhxZoktFauKCRKqRpr6vYWpliEHs2GAm5qHfOJEVOkmJ3AX65BmG0WNRpSRB
CeTbLco57ai5HO7ho9/tJVr8MTerm2gmPAo5hE9PODAySLAzF9LG6ponC+d6FGMP
4oECg4SrdetzhFF6dpbJxv7KGZhvdOCwjsaaCt7otLT7wdgqaKhsHumuHKHe+xFF
c+Oms5XhW7SGqvqqGLwxbqDYayBn7cLExVxglFvHGAL9hrPqQSIPKKLPGy2KOIjn
fWRl4l8jxoYyPzDEWzvEZ20/A1aKHLWOJceSCspVQXAbL51kYW1dn1FqjLmVm+5Q
ZC7luoLXHSf8K4bscbxJckV2fsi9mWkfQ5HzIWmuWT2Bxogc+5Zr0oVOcRuxt/kH
wuYcA5JVPtLpHCRUHpyDq36JfsUfN64AO0+KJDO+C0ojutk6EeaVGp2UBKwUUl7m
dOjftYsGhD/TqRjy2nGiERPlzYTodX9P4YGS0O3vJPPgwDtFwfK8CO4Ls8NY2HyD
OtnlXm0f23KUiaEb3LH14+a1fVa3lX9MDvXj6d91z/ekMk+x5qgoPL9fbKD7nBA8
ZL9e1WPJsrDn4blZ4w+oMm/tOTQxuFMWLAeYbzmH9wAm6pGKBcrP/bnJt4bkAfDD
4mkDg5rWp+/rXlc6+VSc4oLdIlA9q94cAfgSUTnB+SzdXON+ov2blH6tMGLd1DAS
jK7zIDL3+aV7F1MCr1XHScA1oeais0O3/TKM54QIxt4OGMVl/j3JIGXueCW6YZ30
hHGxf8wHv5+Q6beBBjihQwBsIqftBQOW/c/1KLhOM3ZM2IE0rBRnV5s6WXO5U6Nu
YGOw0hSOYmw6kbCY+mxOTWjd44bithfFWLVLWPgP6ftAXQ/xeLrTVXEqTEQVPEPz
GLeUyTu00EBtJcoPxUgLHiUt1kEB28SX3iHeLKu3U2goknWjxN3aYWKeae2jQjzU
Zdij0+S//aseolwwq01Rg2tzlx5fBVMhCE8e93uQ1F/1tKRz686L+MLcoeydWnS4
xJd5YDLlFdEK28SZHEL/c3UkDGrpTbGxBPlP5wenRLu4FASAUIdS8y3rIEehks29
2mKm9LjnZEKwRDx9NTPASP1vXpBbmYBtS23Pm+JFhmB+wBvA6ay0kbYBQBHuEKLp
Y6M3Xc8ch6TWz6CL8XtvyOtGM7jICvAmJDRb+PYormU/le7TNCUpyV0FiaWwoh4H
5agdap+3VjAKzCwC8GxERxIsZQGFmz00Y6RzSQ0nVhNAkXVUTFONVw5yAEJXaVKB
nl4a1W7hLwffG0ibem0/NzwK8FNdhzk8RhFuZefvYAcgmCPCF0OGmYgA7NCG/QYf
ThDMv93BPDAYFo0H+KwK6f25ndb268QtTZaqNBhC7VZyTgURuCxuOJ8OYvAMBhOV
TqyVZMrrhcnZeBaLppmHP7RAYstsqBa+1xIWef1PUetohAVUnWC8QKoWvMkf/6Fd
DecfulskJ2/oVUV9ZrvlVDhpkxuLUOHiTtWnTuVvJGsQMNMjVp2ha+JRlQHvwi8V
3DAH/bw9zZt2lisRBZxj0c/IMbiKnuVLlIHttTmnoyXuK9pDUnYnDE7wp+DR+0B2
xmOMK/DwVQkZ1txg5CG6pdV6VqyvOuIApOU1+kpwuBhJqgo12m21J6T+0Pmp1vTl
DYrnwAoPUu1iS3qVsWO7jbVZhZxwKvZDqOw5znVM9+FAvyMmaUSVdThQm5O+Czif
FOu5puFxeSQ+8rQ56WlM0Z9OjHZWeZh54hJWWDcCn1EGpnDMsaHN3aYrcby+wsNn
5Hx/asGqJVtKlhp2OwMkOszcR4OFCipnRaxqZzWw485RnsplBhGwxnmqrMqNdmCQ
K1X7w5iQOD5w9Ss6G/O6ajI2LF1d9eg30ShhrWGG0Oat9UnVOoZQBBpSAzfizibc
zikA0FU8jkZIbqaP+FZ1qfUAcoT7ASF1RWk5+f5UmiL/sBBnM4xri0zIeY/LpZmU
p0OPxbmFouQU9hpfkIa4+0MO9V+7P7eJqLxZAK2aivjbjn1/M4NSMbMx4TYLmFsQ
rfC3O2zVv5Aawj/8cwh/oIxoT4vn7wRMU+eaD97F1nYZdcRi399t0dSrOZa7GSsp
65uZ4ia1a5HABZkuKUitE9sNBJhb8K9OLcE+r07bjts7gGyLILoPx15FOYjGHa5c
es3MDjAnjVHJzRo695fZItjUYk5uqFt2jVW9fsPjQ8HaDw7IfNYBdla1UvI7lQUu
qbkZXk9S/+ECvGq6MUrLf8NlSs8xb/KV88nZt2x+IQYw6swQ0haOON+AjFnTjvVp
IxQ13Oa61/yS4jC6E8D4DPf6VfcOVv5niS//WxZvJ/yc62RlgstcSY/U4KmkyM50
USaKXytdb2Uesc5j6d/ZgSX3agLo/mcLJ9y2rA8Nx56FKeYf+L/GN6Jcx7ZoqH95
pDUncKT/3G6PfesE0HGSCHnT5NnCgIvq512C0g258L2vL1fvNj97bpAzMum/K8/k
FmNRPRcH3+ZW9bHOAqSy8ZlJJdg0ERWb8QlaHTieApSdKmBy0lcOHZ4qYrB3r4sN
czu0Hi87qKWAu9vxp/NTP/ERLqk5Rx1Z9ekyj2diFkAEypPPKci5vvaHYwg7px1E
2/Mkiwr8DC8k1Z8Tmr63NPlN9N2PGSNnlzDsmb2S7H/GTmnBPFuAHreUcglp4XuZ
Bwxdp2pkJrAm1tsCdX0lrNWBygp6YWUTHirku/YntAvJgr4bfm1GE1qGQevLTZcs
Psgd980phHfERbWAXkMehTMOcwpCiueDaEGm8czkS/BG8AeLMFOgSKgMiNFUC/ep
YP1xZ7Rcx29NGIT2yU+wnoBPLgQMJ0PAHJPU6JHInoasyx62bVjyg2UUiZntXBuf
Ed4cc1iId4LVuCrE1WtcRjpL1JOyReNyMzWN0i1qzly9VO0OsH2+oGXw++nkhufS
hyYdHj2OgJe5im2uYuZdX+u6SA2a2LLwxiWcA5PNPTPml6/Ord57HkpUCLX4QTU/
qegvGMJBA+jiPaL3xSRa4HEIizQSIOGQY5x0Zn9HAvJKNFquiZrlvQEuYHZWNAqb
pNaSKDMR1dHMStVeH2lFSNfeI3aTZZFHWCplBzAXwpF7yjRkhRMWKMsYAeTP408X
v7KTsc7vQB/mYzlaeGRXq2sXeAnOJhw4PWhARdmszKbHi/c+lbNIPA9+NdsJXrZ+
tCDmjsna6BifKTLhKyyJ7rtZTnEgAmPq1TPpCZ/KG/2oj+zpz2mIW1+6styH2nr9
MXGcdDTFFG8GlXY1NgupYw4kO3yBzUDzF0ngtQc4t+txyzykfpyLkAoG4HD8ZXip
x0hqbV/PNy7KpZVsq35W8EFR6D1C3VrXNDpAC3D8qN7uQGzyOWyVQ/RGbudwdyKz
UjMJjnSR5b026g6m4+TNDRrII20EZY4nufL135767SEoqGkDwvVYCtKQomwdDkQr
HmYR2DGm1GFUkPF5AyRO72/JYsdVvHsh3ZqA38Onoyf2oYZizYKf5GFoS4vymnPH
AOevN3D5NR1aPhBisL1ugc4meYXFdMcEsGX4rPZ53hopJ13+RJe3yjW8RSRkVvmK
DQmu3al1MIXBKs3vnV/T9Ew42sy2UKTzGxXDQrdWyC9E0tUXP1yaw+CrVlPgqpy1
WUybnCoMWlhGMPzd9Y6I/DsSDZ36B6aBFAucpcu83EjZajj2BvgxXeOIk4Y04bPw
erHpil1Fda02Abh8xKt5BCG3kIOO9sbj7srSJc/ekF8nOpjUN1tzdNOiD056NrXq
M8aCnlTNb7S1m6XgOK50eDoBWT6uPayTA97grDfmEi6+Z+eJh64zSrICiAY+jplz
NgmB5aIHwqUm/GBQ34VDOIqemwHTJOoKbLLXqv8piiHlJX+i2eH/2cRn2Cf7YhEF
fj7baV14lyNpVKYZ5VOFUizDWVJ6xzU9QSCC2+8HbCpJJrfnB/XIVvI0XoefYl8J
r1C0jq6db2AFYS1ey4v9OlkWtKfyc09X5nWEDH+2IG0hsKBiKvV3Y3j0somwtMah
8caHRgCYiw9C/3bs/4Onuiuux7RKwdKnBWVZChIfitx0ygue1xRetSgY1mtNg8ll
Xtf/ETh1MEQ/h3hhb9TcAz3hAgpA5ZbpRuku0L5LXuGCfi2T+KTDDSfT+6nQvObA
VhF6/OBuxbNzhTY0Un6PCNudR7KQdGMXd65Bt3oPkvIGk43VeWYT3nhbXgtpTnBD
HiArjkSDBQPjh/GC7GwXJbpAo26y6/bL9zW+gCc/D4q+1dTAvCBXxfWDyZ8dUM5k
TM7faJLRdCjEbzJ6yYi+vDlIvPjjEU45C7MpgE2FkGh3yy4DW/UjnSN2/NUGg6FZ
rwb8u8W0PnNCsRXmgad9idk00Xwb/U7k+FIc9cWsSS7Wnq4DNlgbulEVIUb7zcWi
4iKu/kt5KGH3PV8edU9Amo90ukvBd09OM0cNrnzK2u6Sa7tcmJo4/cLLpfWTBJa1
hsY0PrBen2psnIdPrN/E9O0wwp9VoQlBsqmLRJOIiZd4v9ih8+iHksD5kzTrPiqh
oySbrrDtf4Cib9BVmZ24ybuiIdg4lANf/dud1sJ74OXAP5xeRF122y8I1UY54FoV
GiFXR7729ez8ehvKPmJUG40WddXPHFbJtNUUsyzZEqrPCN5x+JU2eAesmiIY0Gve
06l51NtxgmISkELJ8166SNEPy8Q9wHfwBX1UTGDn9mWjgFguktggCw0jAUJutn0a
uc4wayTiOCXkd09C15Dc2K67TwQbgv0ACOW4si8b8C5oMHJ5z6NvjHuX4u4q0lso
jtB0rU41uRoosEJrMYGr7EVrsDgqORBHerV9vNnuLXZ5dHa+wLzPn7D5yAFMkN+6
TviDcjdWB19jruIBBhir62we2JlOM8GFELPp0IlikNCl25CTSBKTopBn2YhTQGhP
I0UkAjQpr1mmOdua1KXg6r3/MRv7hv7FPFs82hTfu9zkWAXbJ7uecuAr19Oxs661
t6GvCDgTCxSBYYaVoHhmeOYELEwX83eSU/IvqGg7Y7wWdqCkI7RxPXHY9lA6oSQx
uGcKspACeMJalCKbF1w4qpydFf4L7S5vtBQ6vzyi3VZOCmFU/gcCH/rbhd0yyXSC
SBjmL6s+8D3kEttEfB2Sg4iAl3usAmb74CZv92aChRWPgWGXRCVKR0Ekvq9cvnhv
A6BRb2DLAwFyBeu9uxt7+1AdGM9TK3PBpL4UE4MBQVkGeDJyEr7p3Zu9pXyvdHYw
w5boeYo1Ahl0/Wb+FI6dXH/v7YFWfzHp/Pqg1BtRRXUFmlrYkAj8rYQCGeyjhC7x
ID6JxEezVZjpvIexSP+NCbipAqRuMrbVNd0kZAAjw0YvABPXGBvdDc8WpWt/tCmI
hetQaTaC0bYE+kkCuSZrEs8Ykiq8PjtG7C/w45/sFz1CFxKftyVtUyvGJsUVKx0G
MYDyczp+PgWIcwD5xvXRKFopD+63JnWNm/rJkzjYz9M9qenK+Tq0Rsh0bGFil8sD
KLeTE8N1eqRdswDx6ECEfUDdUjwD2F5C4aFqZ27jfwh0ccHgXkIkr7fh8hhNy7Ne
+xgmm+mDPBSU064QgxlybQb6uHms6tg7lfZiwpnWOnwtsQeIXIfLkurijMTg44p0
6yRvtu/tjLQQ28ZVBhFIdipJUEWbk2h58e75T+8BYnuXSpBSglyYJJOnzxA/ko3D
NuaIYeVLAnK7FUJyHw+nZSWJJ5Aa2xkoqnF8C1zoCCBjTmmcohERVFxTdxMtsQtP
yoRfbh14cuZMFPFaAYfEuDb8bq/KxO+ahtrrVbEIRpeX0N+1Z3sJLsQCVz/6aRcJ
wAbU0mr4pkSUgb6tFcNZ/MnPmz4Fekzd7JcfbDXkLLviw9khFLijAj+zSxeXETD7
nJH3EsxRBQXeXCzGiejDK5bZnFXVFL5ClPWEHMKaEsnJfmhubqqRcaVYahvEGH4c
31o/OtwwMLBorh1Tv2NbFKnoNmRLZOgmcpQt5srjKJ3fTirkgFVZzOGQlYiGpTkx
G+CRGHtAizji272dP1m6pvBjvhiRu5MFaFTc659ts5Q5WjnbK8mRYEdtRjogLThm
Ckfa2GPqkNx02c3ih8Mw/CKXomyK4LmVmTMJA1FCJ4Pwf5e+zd7Qhb0Z1lpX88Un
loc0YY5hLzWtMc2aT3RiMjyYZx/v3HFrNBYISAm6zaSjCYjjdvCJIkJuFH+3fsLi
qFcGViAPYdaPCmtO6IfRLd1JPdl1M17OUfG2+dTd6H1482RYtBkAGVGWYl6Achac
02oi39HUNZ27q7f8XH96fz272n1dMNFDGZ9bJkw7cr0gicmJm42YpD99jXL7/WB9
9PE+bZyqzLWlRf+6nTWoqTAIIErpuqSCsGVekPazCyeX63OOwedGAI40DLuE5FK/
/tWl4eD4GEekZMFGFwJTXKSFgTyr65urAb4jahKfhrkxSFschOn0KnVo+woP3bFT
QCN+7zLKg3H17/tShJKnT1P6LssVvkqxFzLcWq55stMACAQe2fHSk+BMwfmxlkUL
7xpnv+9FbqF0yc8Ttm6N97H5Ca20bZvAQcbSxmut+FnUKs4vwBvi2vr4PlAJ7LVG
+mOXyBfv88mJ+9YkTMyZSzD88NTPwFPhBEfm50e75pEaocHgboWuSn2jvq8X0Bnh
puTgKQSDeiR/LEgl7/euENkmKC4sfeRQpcipxlYqiMgM8H4+wgCgloz2DUg9TlkN
dAcrbC/E5z0YIp0kyVIW1xrx4pHgjxga7XuPxcfUQuyoCp6Ah7dBnigMs2EnJoWT
qRmBQ+TJ/xS/00o9dCt0Oo7GuFD5xJmCfa4fsbD7Op4Go7afFImZ8nN08tvYOd+3
16/VmyJCtWdzlAkw5uB4dSnYDxoQ7ZBT8ILlSnHrsYTXJITUfePfjo1AJXxgwFyM
KKXSV2dUCB/Lph1y/iP2TJ8OtdxcfYZYDJaRMktB9mHobabE3g+NMiTR0KggPxOQ
BBHqUgFlgg5lAQh55Yc+UYuU3gikCppWgskdhrCxCaPGXpOIj2JSfLhK3WAMSsZx
abtMCw2tq0nn2O4UkS5Aq4OWhqEY7TXRY0nwqWuSvcIfFrvERd29RsicLvqH9kWq
QP3C6vdZRs+iI8XC1lDpOfxYQEruWrEdsFepz77xiwDm5sznntJW4FofyyQGr9tW
pdGLVD3+jO2J/p9bO7H4sgXDD2/frKNuFFIKXORad0f+jPQ76CYdCoavC/LkYYBt
wcnlQpjc4jAS+sbNtwnoJ6lu/lCdRfoHZnn21L94b9PXvpzyPPXJOVF9Hkj30ycU
RpVt2kFRIfE+u/MggP5y1flC8eOVT5dLBLSPj8NrVE3rkiKPnINWjEOaxyJj7eFO
k5qGLPZrsXBQvjdVEqzLeIKv46QKliPS7qQO20k4t9/M9V0kZQ5jfUzR5h/7Ucku
r1DqVnl8USkEJxlZFMXMfxllY3s164+8HvFB1ZS3K21c9YH3WUML4Yv+gSoffwFO
RVs8FkTkW4N+qGPbmDert+h7c1bfRHxjbNKrfREVuYIpNWq70dH8kIfrygpc7+Rs
WT7UbZ7uvxvA+u8Sxb/ZUMNz2rZgvJpyqVrtAW5lIsxPu2Vkg5Aey/JYq7ZBHI2K
gSSJbp2twLWdQMYpOvVjjtEKTAXAiZXLOs4UlnTVEdVZVTxJxV/Qw5OvD16uQL1C
cUyJKyxSQ4t0zP9RiVNx2/PI4DHCmvGjHko52tbE5j7p2fjREOUIwnY+qbKgLBVS
1CWeyVSBDlzN5+RS9oIObubVj13xomLScIUxpql6oUNbKoxpb44NHHGrGBNlkS3B
K+I9mbtc/QNNdHMCeU9s+hAbzre1QNrcF/xUXarAIK1iALgLjVuDh6P4huWLt5pq
H2DgRb7LV64b1xyLnTURRt1zmieGk0q4tBna6LPRGLFQuWbtfE1H8/zFCHheWBzn
Wo5csAhxB9LM2AKwEf0ZXpd/ehx+Mo8Tmi4mWvfIPMJvQzcnFv1cd3WDAgq0EajZ
hkMEngkwfoFNDAfsbfCUb0sJ/y7NvXZ7YfXDdve7l9XJe/GAjkAahZthGLikLpwd
fCvkfD+gmi6AfugAz3Fv+xesF3oioZdI+3kICL57eKEF/2gfjE6oTjnQSHCI6trG
X/igNX8tOHIfkVxnO0N3M1tE7OHp7B2G+jJyL6OOVyU6VEK21ZQdWZVKb3AuW9cE
036EFIXxT70hyTktLY0bPLUnzDwXZpIYT6tErWPk4qQhjPoFP75uzUU/eniWpDZI
44b0neJVqKjNtZLg+o56/fNBCz9Pu/hEr3HLIqpWZmYDvo9m8G2Y9lrWRmg6yf0m
Y6y5paWefDI4skoDFSoRELPyEToxeQ4LA01e6FR9Eo3it4hIEBeEeRGDAP4pcrQU
lBb/yX6heagAg2YlEbRnlqSf6OsdoN/inKzuAKpzuDL1lSO82Ja3TKlpjX1mLUZT
Nk47WEx6M6GQbmy7Ho3wObdEz/9Jek5dwwGdQ9x3D0/4ZD05TBpUrJLC7pISbFRo
jYNt7+UfQL+II9Bg9napnEHQDRxAlYOcbkKxysNdmN5BkkV6mqK0iaR6dtwWXvQj
bldUZON+PfZJOdd2Pa6JvNkSZL2o5ZYRngjOf7X7Czu1m+CS5R4R2vdz+e6JYtze
VniAd7C342+9wQQ5V3mzTPT0ObQ0sCnpS/UAK/TZRruqijIGRGJsAG90djy671EM
nC1Os+IP5GdYHesDPr+ynQ3FXCjq49FB8T5Su8ZUi7SiwH7PMtkDBrDNIoSQHTQV
2lP3JbWeJgFYOmZn+tQhVjzXb4Oqt+90Ph++FencrJhVXHn9tFuK7ZXs3Kr4yRqo
J9ymADKXBjRmVi0/2pbRmvdhG/y7tkfElL1evqy0JzFNjXZvQ2v6tZ+46OKfICmU
S4skZFpqHFp2ZWqaNwwlHotuNzR4LGiJ67tNHtqvUHYe+2gsV4WbWE8bN/1S3EOa
x0uP06I5zSrTevKqdZL3Fs8Vdg1pwDbBugBwXwvRStjh9lk/ByNDofXJHinzfoYj
5ARM0R/L2YrmMS9NKQmPMZqOOwTxxEecgUWQ+yzifFHYQW9W+1Oo1K6m/yTHzgVo
UU0Hsj1Xk9hrewwlADMHQxG7uwgjhAe9sajwyu6XHm8vJQvxtK22JU0fJja1DP0L
sCtHO+d8OVYBScRAKW3NlhXqXm7FM96o6YejSCKJR4JbLp/CIKKRuDA0CoBCChzJ
jGLpmc4tQ3D/DWktrn/g1CeTeU9fRQHTrOeJmx4EeXkh5oHG8EmS7mfyi23w+lgM
aNo6vaLk15ZT40EFVtHF1elOiUkhVNJrjvnsXrA2XezHUlIVGAybiwxrNcpvt/DI
hh5RlC52y4jjAVAWyHUUDCbx/ewTlYa6pc+pR6pEO9tKInDXZdM5FTnz8wXsitZW
6ZeI0/JhcRBYej3DbuhUwZxhVXEzFZxhGeJzJkN8LZVqRYlhLiMFE0dI+Xa0DsTZ
N4nyxe/HuXLgqZi9ZdZB21zXbjNms38DfT8AwhbAKDfQ3H3gFp3ikWHIad8st+3k
UFr4/F87tKQM/oqcODS84vwII3bgnxaypW9WY1NASyExDYUkGwdvxtqW0tKc49HD
MIi3eraKjJIQkYZMJbWA3NYH4/xaWZRsUCHk7o5SQPpwtORtpjHJ/gLEwR4T4Hpu
8/3mGZ2sRPA+gRhPZmsHB/D/4xy79JTdF2433C5+nuQ=
`pragma protect end_protected
