// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:02:11 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
djEj2SCHRxsfdMsV2KNXIzYzZWTxuqd895PHqz7ZAKljac5LwH245qZcYecTN/Go
8Nhze9fyGi1/AcsfS6ynNfxbwcWr8f0sR7DvzIc7TLVPg+i12FCwtZ053VKamlCO
uIaisnBtuYJbh+kqnJoJxwAL1FI9WIKibgXkWHiYoh0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 10272)
BgXaolG+bk/Lo0ApFeOqi8decdqpscrt1wYwOiQsGzECyonFidz2M+gDahepaqDL
vFmhp0lKErFp7w7pbl93EUN1qRXSlcigJciOBattPditE1Hf2qbOX9lI07AodmQU
TrCXpMH9DbZKWRfRdOITP5m5se7kTo49y8fmFW7E6uf05rw7dLlqv8NM8vdc+rbV
e/bq75tK+BVWm2yNZ4uWbaCA1LdOZJLs1k33yxoo60T0CyEr09IV04p9t1ZTsn32
SdyMCYLcxlmcIwXI/hKl5ZAH5oxnr1Do6u9pJlgNO+29S70MQ2VTA7R34JhYYCs+
VqZamqwrmU9psYyWatj1cRnnYUAYS9LLyjFLKiPfEtfST4O8zF290O3OPXdycfOm
mPm+hCu0sorKNOQKcedvxclB6ddwtTXwP/f/R30dVfq4N/t8rVS36c8F7UB9FtGq
j5Emtbo9bNgcr91H+5UZ+Pumdx+t//l04aiZmnlwRdpcLmcGu31waFLMYWvizrVg
NfCmUhTGgc9GbDCKrmRYKMpLMrefbwFsGo+3rxnD+BwQBSm/SebBXzJVQWwRVEIt
AkYIC+2v84Dw+e2TsX/Qzvsw11JfDyeU8wjHPwZ/gtXTJglejrm6/FF2mJ8uPORR
rUEMAAnVMSAGTG86mi8GXJdY45558VwQbn+xNChHg6ITVHA1CGJBFbBVgvqvzS6a
enThbBmqnBgSvyPS11oF/nx9WDyoAW4NPfrP92il5lpGSfORYiYyB1VW9dySXD6q
/V8quk5EGCz1JJysdRZnIXqCr6qHjKgUkZcGSDdGJ2kWckNuKPH1pNqqLWjwEvz9
dFFz6wdkQbe6oANAjmKeXRFQQ0hcLoQJn/ejdrQo5mZX+zTtS/MV24aGoJnXGqdb
UAgUbxHw1pAb154W+mvO1jf/AeNd1l/jhbD5NwkIWlELApCHVL1uNHyOfUEbfJkr
K0PxUwskTFYv7ZI9STNfzysLEdOc80hQ8UUxDjBMmBvA2WuxnGfJRPzo6GbuMmQu
ffyQE9EPP58yjaOyazveeFXCpD2OvxW3dVc2IXw1by1Tl0ruJBrbekveBnlNo6jt
+wKloE1We/PGCYLIqHsPIlaFtZqkmB2HBePS2GdJ7uBBktqBzlcUOADPOgrEvBna
B4yl5SuN/iTTd7QJw0qfRK69D9/DGh4vkmKEkIzuga6gKR6aQq4WEQNZmZbOpW67
uRq9xFzvC+oD8d+9DPirXXJ1MdHHXAW6alh5We3bKJWMYC2493rMW+GEWO8BsM+A
C3PJ4qwVp31wFQCKfmgj7tBDVU55ajAg7NL5p3LQZGjgTpKsmx0oOJPNIAYXTgZD
65ku8GyDy8Mp8EdWng0jR5QBeiEpmeobpj2TBhAjSRR5WVE+RCjX+V5bIXZU27jW
d8pgxikqvgNxX40sk3MVvI5plh18O56XziIfUxNOjn9rGFGVItqbJ5CvZ2rlbk6J
bhT9MVjuOcInIaBCXlKWVVS0tCy5rDmIM7FNh8geKUiY21XQSouGGwgDouutghMG
dEEPUNptgWXacxH8AwiDe2ZJ1tvZUGi2142BPtKJ0FRrcAs3ehOXAS07FLZqc82b
4NjBESsDnW8rf9HOA7N+lkDFgSkbAHQjWZwPQWPE250gZBrjBAlkd39ygok36xDT
PVGG51lRlPH1eAFysmfO3mIpbIDBq9EWYz1t3oxw1y1VJZ9LtbdnvZdF12rF89VJ
Ho3fWPggwu6cex/C8JmC461+T02qyZY8yui6yHH0xMzMf/ppGkYhsPWsieiCZKBG
XGmnaWFgRLe0SWdE5ITITd3fubMO/grQGQ73vP2Lp0icclK4xA+9KQn47bCX+i4Y
xa6mqjG0PmQKIHbO3LVnTgaadgZT/J+gA2j694+cKpv4mqkrKldX1uvOFnDFJzAC
SqfEJN4L1laPGfwHVB/vLjOkhncmHFCxSjM/+ofqgfscXwlkyhEXGq6t7/xeeZ8v
+p2XDoINTIIoM0r+lbbEEOb5OGSNKOd++uDpVwUz9jNUpT5ASaKJTYXIqT2QbCk9
9dzdd1VesM9AJCfgzPQrSS7SCZaK2/zirOF5Lw2mksD0CrJYb5gjGXBkBAtL9nj0
M5ezmHSpkeI9XlaT+cCUo47RG8LLiZPJHR4UoT8ZQXli9no9xjxo5KJ31J9wuPSS
jS2e652AfZ21IZrMG4NfmTh8xJvc4xOoc35o94+Fj8LGU20y6HYd5bRdPo589JRF
KvICzsAS1lEh5qmkYO1GDJHTt77BljIQ8S44Gt0Wv4EV9csGEmmF0Nyl1w1YRgwY
uEQUXF7Da/DUBJvft6Cs09UMvYbY7hbZQ85rJ4PFjM4HClW+tNfWnDpvvf5upvEX
L8E7MnIhduVz8GtLY8FeySlf8Y2UEH99QZAF5sNXpUbMnW64V1Hb88ZVhNlZvQga
pFqV/LYGSkP3JBjsvauNhH0wkH0tyLg5filQs2yQqyBHvMcRUXhKhQ7HdL4S0ZPA
y/S1622sYeweUjOfbCRua7XWt2A9jw610NRNvqfkmBlDtfGhjxtzt/1zKv0d8Tcd
cDfDE8YN6GIn4FUO1RQwhx1cW5F4iVpqjpXJynNvjVzt04/WfFUHksW9Zh7FcaNI
Iy7p8gX7GB9q40kfxLpp01hqxZ9PufzVEeM2/Jx4+5DbBXQDdaUW+Tu+YmWluo/N
jdPk+gfjeqi3I5aVu9r3yL2X03R8d0iG8L753lZdzVEUbW6ECE/S4IVbD3T8jDqG
hMv5KCzniwhPXU0Bb7RZNbI/fvAsNOWMRo1D5z5lrAVMOTalndrsFMj71aLw/vqu
qJktLC/H+6S03XOutLHZt8g9GfsiYrRc9i/BeFVTNThBX6k2gWr2fSXCDIUnHM10
7vagBHVVY7nlu+Twh34uwhs8xvI1AJsOWjwjrbYashfGm+4+c61oRgAcfI/kVjrG
KCMP87WP9jl9L+GWmIqcFtWDSi8L66SkQ00PhuaLe5ihcEpV6HgVGywoo3lf57eB
LhtUWvUDePm69FiuADSqf2JSFu2OSLGR9szrRm+jOCL7X4+gyl8xphi16Jjj1TZX
cRlQO6rvw49rbuDzeQc+MPg/1JHlbSjYWQbhB9+Ih1lXADZV7U1P+UfW3UOdLOHW
Hn91jQgGExh7j/atOQyqKq1NRbUg8U4z9n7VWMR6yRu4gFtIosFAy2p4PHBBUwTq
QRgIuhT2HviaIjm9hr1Inw0KzvLawykTa+qs2MzumO/zDN8eSH55tXVtfVsnm3yZ
DHaMA0nglPpelj4dtiGPlHRU89aAakOXcEZj/PBv6yw4fh6128E3QCxPw0LmOO1M
MGA2Q0JvaTDHV2ktqSdIoGpUbvXy8GcekLLSOT5S4uKMm/JN5PMl37FW0wqAkl3V
9Dbb8shqojMwyBr0g38C765sM0HIV7ghwkrwpv0veC2oqEkspEeCrtoUDvkeEH/b
KupMcZMJYCWZhPD+S8ybzjP3Dd4ECJW3NVRGR9TmbAvWeVqqz684FR8snk1tB71m
3icpMhGmJwEHCNBpX6+dhGEj0oQz1lNTOcuIdrRUPgJvQl9f5LdUtnQHIWwNzZ5H
br1Mu78mz55bFYltfKJDZkMrhV8/dwfl8jib3xf5y1LJypt6k481KQ1pbu6oQAf1
gXzTgLed/k2BUZjFQFqYJzf10NgqdmBpMNEUlt78RcWwEemDR4pqdbqopbQSJW+z
OjRvMgncGro4EzlHUZ32gduypo/zLrWAUlaxd5EJK7rnzFT9RlFjClSmbLSZbqIX
eNPF2BA/cpvPKJ9UnnWFQpR723vjKJjHa/a1gRSTzvF9FpFT7aH4FuZaCmpvwf6I
rfOIIFsVGGrgepXk/x0Vwd4pCxkaLS29/N8aImlQ05a++V1JuItB2k1BX8fye4bf
d+2VEIvfsQmPPRG+J0Hwzqys3vopvuzvz49maYLSj/R85fW4viC+/wOxbRGWDQx2
MdhQJEu+paufFwEapKNVTfsrMNnoYINziA8aN8d95OHPRxBLpSJTI7oif1CUafG6
hVeYUcum/QM0ud7j/088oQimPE9a1cWVULHyeapFF7UAGoJwZxCAglUzzwoSFpd0
G66g+CDd8M+YrZ4zT+T1yApDzR5YS16hUWxtRHfM2gZ+bNHmAObCL+oTDsS2BluO
kiQrDZpDqfsrTXbZg8ylXSKXtYaZxvHGV5FaT78DWjN7FwEkaRI6FP7wYEAeaqIL
FRX1RnJN3MGr8ymjfBLq08BnqnVS5mzW3j84GXr38wLMoul1RLMdpt7OFAL3EJ17
zqBFKvFgZhETHQ21lYz7W3XBzIXcD3wZc6mk1pnkD/IYtOhOe+vjBAsTVh84ePWz
USJxd4JdBn6KMuCHXD8FMwA7fy9IVr14yLhFhsM7873YHsHxOyOgA9qr10+76jjD
xJe0qgABrHmpQ5B/jyiNGa69XkC9NRaBIzy0MyE0M7WABJapO5u0zpi5693bFs+T
y6hXK29ElgO0qOcK5wpB8pRw2cc5uMhvqkPuAdlYIHQZrRxZlDw0aor7T34hQZjk
z5jTduNHhLBSus/UZ/3qF2tLdOvtkwQMMU9hT3/sauJYBUpbd85hBWnvuQos0J7t
Fj7RSi94H5Qk4RHNVmf6HKSy8PD3vcpkaoB1MPvmYcPkCqSe/RpAM3ZkbxYDbKmS
Ch3WgdFyNPl5Ft8wbMYKi35sQHXEluyxbUwcWEGo2ypiVCNy/bXOuUYnxlZxH8Nr
PkInd6oOwK9fNspmvmu42j8L3MCgSJfejr1yfxIQPUULGtKo4Y9qBwm7A8Velug/
tjsMyYGA/XnFa3RvxdjcxBpDsMswL63Qgxy5J+EBnY3q5JJTfo3+cnItlsixH5qD
MSGTDdXt7j7AGBPyAJP+x+g6os5gfNUetie3cWBad42XfgcifDoqpmRPiHVOUUgg
rw8rYh8cTCe4XVhsDHZ1n7/ZxRxc8QR5Zh7g3awW0WAy3iJogR+7IL5+T43fpyYE
5d6gJC5H4DkDX57ncacPp2PqPPUE8i5aNlzU6MG/pAnpV5xdMngRlnXjNDAwd8XM
FSCCjIXKdwHd34+pNf1vIpLyLL75wH4aWOWGgd2D9SyKZsBxDYKogqL8SbAzTQJT
cSCUN6bt0NOJVxl3WClL6af/vjeP9PGQiKbfnKaAgFDaRs0QN6t2xEXD1VKlWxVZ
j1Qk1xSWGzGpuWTLdH57KLMdtDkCR8vCz6lp3ipns/Z/HjVkDF+ZqcdEXgUYIUW9
z/KZcZqKAD/dheojt3Y2wk17lKOEa4uz1jg0cG7nrRkbFQP2WalSYPPhhc5lPHT5
7h+dBYp5HiL+TupyZnjH6Ponlzyx2EyRGzkRWYXRoT88/AByxo9gi5zMod7Xjpda
fvtKvYf5moagtb6mnZrMbqQzhx9QJ27ieXxUINsgEaiNE+dFMMviedAIS87bLtP9
euF+QtqLIObJ/KOxT8R5Kwb4oiYbLlpQzL07GvyFRW9YgYaoQKlQ+cBufig5Jzvr
q/3YhsvRo2y3OPi09eJuTJaiWhBgniWCD1NlTz1h5AQiZRQSyJlWllQXMgmsKr1B
66iAlxnomoZOxORTIVoBTlz5y9pHNKJ1Q9MPbJOVV1b3Q99A0a1kSWBq39uicbpP
5/9XeKRauKK7KxSiav+Q2A9rBW/mDMG1alIIscUvCieMxHZneosCRHNGVfPCVgm9
YBrqzv4BoPJKz0HVQwkUsxkzMOjSHlb8o8DR0vscu876g5Xe1jwvOtF6FaN048n2
Ku3RTwVryBMKGeLz+viuu4eQur4EDLLNufG5fW2zrSTBZHe1Qm8LCzJ6owexcNuW
69pQr4WZx6GL6tnVk6xmcuAxNxt+8b1qEI11OW1M+ja2hTqLyrXBgYQ+TtC7JuQ7
gOuxp7TKnE1DkD/w/NMyc2RTg/7trKR/ULjmJz5O17lpJDifjpan0NRhs16irJPv
tD9oOn0XxDhXMmSgF7ylynCqjePwSjO0mZTyOKwxJvLbG1saUs+eox9mmTeVx7cE
SdmJcO0VvlLkZ3sOR2d7Q42+sNCwm2ucpsjyKrN8Y3DL+5BV/Tg2oE9nVIvKDcAT
yViEreRISmuZE9idVNDUby4lnmBNDQ0Q6h+vvcZRJZqLMOqg24RPGu3xN8avMJCw
FxDj7MZCke+Fe3aa+1SMFciNpcvgp0uHA6ywTCz3zQGPZNMaXPx64fiiG1+shxUT
7VLX4GcHvsGgMTs+LTpQ61+YpaGFeznGtszAzfI1Fvmq4aMHp1KOpURhUblQ15Lq
ruto8vvnKgeX0P5xlX9C6AGQt0X+t73LoYYsNais1+0WAOFtMSYYar38q2NeJuOk
0G9sZ71b2R04rtmHwVB03H4URoF7dmHuaDppiPgY2FwX4sZqIzw4CEVeULdOp6kw
QbZI8qeXdoYuEoMp0oED+X0QWzIaDMrfl7MGlz5SHEXZNClzkS3ZFIfN9nwIhL0x
KNZXSvB5XOatyZ2yOBAtCdvoA7DqZtDj4QPyFPCkQufZN2p2KxZgERhCdj9Fx+Dh
DdxWps/Nyik/hcnG3Vd0gRfvce0RSNVKReNh+G+5pk26/SKZN6ZCZZKHtQMhZw4b
y4ld3GjPrzyZL/W10nv4issrs0GejQE08TTQZmdOXxw9/ZYV6V1OicACg1QRVdJB
HNGhi+SJY7NqtD/rYfaCyd2osA6Rz/5j9p7mjlgwckkLtRa2iR1TWXc+62PsyGk8
pBqUmBAN6Kn0k6MoYeuzEpYYTeioBJe48AkGXTirnxfSaqTCqDnduLu3XMVqZrxn
9joV0VgMxHsPDYgbVBpNm7hCpSitA8kF5ICckQNRjnjSLyBFT86xI0rbjXGWiW2d
FZksXBbs15NagICLUpf245DSwrL9SVMscsUDHDhu5WOUZ9k5VRy2POD+nUSUAW9h
YhlM6DxSYLMUzzxUEBKkiNyl7mq6ScNb0Ft+WsBGiRbkaw5iZzif7db+ylF4Jlim
44iSlUefBe6ca6PQsjpgsmm+VQSqmHHh5hsFf88NiI3rEXXJeq1UKmx8EWU5d4BR
B7IMmWx7aVbL1Jqizmnc5JKFVNfmOBzdNqxElk+sml3yWxAcmHD9hbh4OxJdJKvk
SO1yScGylShzE+otY9Suf950R7UKqCnZOJ0ENi6S6dpsSrCl8C7HiPBk2PPYPcCD
9e5q8lBGCkoPbY+RCSI81TJJl+raDy8sXog9EdLcLPmuAQkPtQ6h/mXsOAfpcK8i
LViBOxC+q3FwCf3ax4ajunpFTEBPAoj6YmuiWRV0C1DSY8xRACUo0TLSaD7QwaZQ
3ROQjIu8uJn5sbizxihncYbPiXe+pQk+6VCPQqjAVutnOoe6BgwsrNhs0TC7cPDg
cavpuqrY6vmPxv5cl6lAt75/aZEWK69asko/5hcfV9+dvJCxYCXLAQ4Ye3uY2bMz
H7VbQPxeLzFaCJyIfiejcB8lpTKDrXGZzRogxfUtRBzMQeZw/lhIeoUApMSA37M3
J3sv6UOylAUwuvLDQJmVzQ3Xyluwc5CsT8f4v2zeeJrq68TzKgHdS+bUivc3OmQb
P9uhotM9KYHzVg8Loeydgmm6dW8e/NMcGBvPByejj3ANA542NBItbR5eHp1OX+mS
wmhUCjRVJymQdbELSahPjvrZDlm1Mm8k1z3BbBClMJ7lbrIyrlmUGIIWC9SFYuvn
kKIG4Chg7W9bS+Lpx1ZVz8WXTb5KC3CyWwBwAg8vMWw4mfsCv1Q9a8SRxPNEyZ+4
/5a/vNEp/2M3iMwAXbp8cNU0gsEt0pycMGalgKH/ktDzvApKvwOK770msxBHikbj
+vDaKoQVTYRkcxNIHJQRnErmdJ0LJTYOId51X9UGb223WJnoz4CCsswoOhoTgF1E
sO5k1KO/y8DZYcOoeD/l6qoZc6voilHEIDZJ7jorgzY4MlxNtMoq2HY0zN2d+6n5
YMlolTtUiEDy79sgv3cwMX5oCL9XZ7Jj/uhrsoQ5VpZSz48nPja9oHVYCaCKM0/s
/0v1Qf4taLrBgyp8T6kk/spC1wwo9EhIhwMs3GZ/uSnA1QgSrNm3GBhD5h3P+ANo
g2FB7vMii3qlvvD0L9HwBdSIRH3XdOdAPdjdtTrK1fzo99KhAbgwbhekFOJ0TUZc
BnlwB+jWCYy484wSLf2w6zGiEqsrANZjqzdmuf48hi4nJUr5uM9Fq+DQ1WRIkfJ3
i9/XpneIxYR6+J5F1ZNhEvwk3CJ8b2Od1oJJtLz+oYVeeqpFvyOjz4zC14nmRMwn
PWujghJZXhz6EDU6J7Dli3AcU4jIaHpWFrJfS11HRX50NYjYCOr3p6i/+Xnc9v9r
bDd3MQgnhvlLl0M74SpXJK31mxYAOoJjN58r7X5oesMMFHCqZnuw+qQ646TZ32Nb
7CCgAYDi/Mzl04C1RL6bcO0xmIiDmBuGOsiJKyL8SZn3ArAUUh2vqhs5e05VXskT
7OMIEAxoys1D5RRvDtnt8LDBHsEIXrskE9aQZUjuDE3LDBRz1kuDovu2gZkQkQU6
6Q9kCB7Iuvsqc+TEhdqvfkAuhH1shebwQjlpGr89Z23GeLsbrQLvcTdrHBl5keWm
RCZmWAQBAs6KoVNjPRxdGE1Q9l16EzMpSttxFWGoDjbPZVt8GBeWHZGqm2ulHM29
9Zukjq/SFeDnaFIq2aaKzpFdN6kOjR/qLr+oxRkbS5nHie3dvzgLZK8Ut0LTS+FK
DJ4LZPIm6iehqGa9V1QyieCsZL0H8edXRVheDl0/lV/Et9q3daqG5Ec7LsnhWVTo
s1/NHIqE4emUcALUFUPKYPA+ry1UKuB+ntW3MIa2BGzHLQeZxCWJM9gT+Azd3xYy
3/t9RyB3AlsKxPTp8rmHIAUrdJFzbheFNPqHcDPCj6kfmSPZmQH9hNWySsxZ0hk2
RfnGKXS/AVBIu4ldy81n43mHvm+k25ygyFVQRT9ljsX2HF1FvzXSfI+FiraFFi3n
0lYtk3O0T5sr1ZtozmzG0nJ+S2xyH6jDKOtFfE1Pxad3wLbO9ZnF4Kz82n1Z0OhU
w8Xli56LPsx5T9FzleVYHgZ8zqQjPivFJ8okQOGnQ/kxYhQoQVkAXC9iTNrXefoe
Nb+jqCMwm0CtVyAQRd+QDCpviZ1cAjXk+r2eNsG7C6+/FiEB+ATE1ysQXkY7TBO6
FyjbkRwdra4cEflW4+HbPyU5AFGJIWVyNy5c6i3XmO8JX36iXp2F8tS9kfQO1qAc
/QniGBc+khfeHpqytPHpRF/M7Dhbi9J3yR5Z7QfQ0FbdIglvDLA11xyTS7yQHdau
KMKjonWC5v2a1fhHDXTkvM18qmUP9hgEoMEgCmET0Lp0v3mWTnUy94PCKLm8aRAh
KrHsnfTqo9evAFiriJrgDL+RxwVx9T5Gq7r+ISY2HwQE7g2w+oimW5fbM99U2jLd
6z6mJHX2CmeqmnJzZ7XpFedsKCnU959xH9WdpaqvOxq72nNL9Ft3hxasUst7rtDK
ASxUA9oNyI7L2alLTRy6egZgAf9b2BRXIaknEQl1DneyS1kGexFQshNxOAcK91/t
nI+gXnuNuBo8scAHR9P7GQHpGpcA3Q79XoiTMWEpRT5e0Nm5HSOIVzH3ItspJhdL
xTfq9z6DaCQK7OGppeTIIA016Y3fd/dCm1wtWKPy3PxF8vSqG5S5Hh8/gnA8GVUP
W0hitFHumT8J62FcNtCZDhZxG4smz1t2kRdaz9Ap5axyHiTnqHNRGVtLbj3TTkhv
NjReb/PJQnIDH6sdq2d2aMGff7f6tEGG2RJL5KKs/I97HNHXfaDdkjp51nSqaJdk
rMCzMemJcql7KBroXWlyotWd+pAsfb1ZI8uS0aZQsdVk0QKXpw03so8bb37vtIJn
2Mc4MFcW8LRBwdv3FwCGjvyCIO4+hUsg+5IFkIUqIhUVsz0WDUDDu0vwtWjRau2Y
t3qyIgV1PZsrzc7YA3abNQq/nRfcMkINXpGhxkfy6CxE3y6aO78KCFcwQeb86B0U
c3crscv2xNpcQqq5vgt597tKURtKhePKqPYg0lDHbZVgehbVKDKs5fdu5wRdQnsp
GJPoT5JK+riL7sx8ZMW9cAWikXwcJ+s37+WCCpXbZLkxjMJO0eHgFUBol+SVQjuJ
ejnMPvsdGm4RZNGCbimlJEOfHpqNIs8CTpH8vwxfTJYrK3+YSeD/r/2HayRq6XXG
nNSHqrSeyO++NUW8iWgVPNEydpkQzDo1zbCjdGK3zrmsywnYjKKL0rbDWjys/6qY
YEivGrxdDn5mD14FiyvC0GsORcjKAciX1ujebI/fCo1k8lX1NU1HlLtEG7Yj+84y
jPa9ep0dDcX7tpYhp7ChjQ1hHkQwMFYXGG5PSZ8ZCYYClvFqlUk0EVbU8DYmESvR
eKBTWKU0Cw3K9JuhKl1lE6Pi+mzLbyxhSAY2Jm6dKEBD0Kt+EJWqZUybnvgYJAqf
7DDsLm+nGmsyWiEgzNBMLk6LvJ7an1ElMNN6ISzfN6RU1EcPi/JahP1XvjWL4BKW
HyQviml2IA5tIWGUaGDq2y2yui7wazYgl8FfUQgb6krHNE4497koO0uxBD5GeHA9
CZhe8Uc0v/PQ8guyuGw6OEMTsoYSCLRiYCoD8WIpYjxrpQ/8y2zSTpRvy28MbC8V
fmw/aAZUxaXPAdpBfDOOScd7UwF3L3KrskqZkwuGX9/e5H+fBLFBNzG0c58BOR5r
3RCTEwhqhcdKpJsqY1TbfGYqWwfU3GAGWBeb+2zXFuIGHRIwiHLs6LOnEcDSKlsO
bQgnOkLCMRO12WYNDDizY79pHr4PZCn0QZaASfXb4yCh3j+9gGCiQc1IBdkQ6s6t
2RB9sktAqNXRpDAllzchXwX+GZaQMyGZqHqZzQtN8QWAtX92AH07sjF9exs70Un7
i7vp7/D1fE+c0vGQdVPdpgvxPBvQSjqgOIu3vx8UEWCvxF8myoMlxDIf4IFC4cyk
xWxcHkIYSrUwlbo9H6CYMDFvFnxMGCWFvP6MNiYzg1bYD4vyqUUL+yUOq1BKIn/Z
ilpNGOZN4El/DrY69pXoyfzi5AK32cS8/HqMNktvMWDTRQswgb9AUD3yF4naKkzV
10+A72FkeZ3kJh6FzinaxnYd4WlVIyoSBBsImWLkDZukZ+uQZXgLPLC3O08Tk2xS
+xI/90Sz8EIn6bTtacRt9wGcMrzIsPbUg4Sk1j8qSfijr+NfvvIXGibhhETvfAtO
/j2sdL32oSdwDot71672IjekeMjKPDk0Vn9gYCVAKKqg+Le8COmqGU8PelKdeORE
/lh9tevqlrlHuM/VQvcpIhgSVrig7F3Hsh9eO150z/acHLEe9uCCLI4+W8p6SXtG
SaCNqGd3TD4aGKRkzO7/siljeulYPBbn3JshqAdeDb8X0mYYMI+72vb6/h8Sf8Jh
87CynW9L66g3Wpa+hl+i5W24+VvySeYmKkTx02ZRfgwKaPdQauamiKxodKek3ZYJ
1VFkBJMcogXmrvuNQ8uBmZJqanpHpmxF9xDUT0/4/YEyHff6oVX5myJ0a4f/NjbN
dUHV8al/HjZwlh3gLlbofHkE0uyFLMN3/E+zBrMZ8GhqMnQVZWB1CZAVCvcwYQGh
7NqkiVXyAtzpe+BRATZqTTwivtyu+OaxXVI1LYZP0umUU36k6+Oqpm+JVpACHZD2
wNyeG4jry4VmvIAP4488SsKZnnmqeicXscwH4rTg7d0ZpWAW2c3mGwBdFtsnfFiU
vSuqbyimgUdIWzmUPF/tG1JwyrEgRSRggEN75ju/0rRP5SpPq11nZuiNujRZjA7N
MNNMmG6CjJpIkN5r7P3VdV1k3LXhTgUcYYscLN/eC/oI4boYwdodRuVT/eMV9vIj
o4NgxDYEjRGK3keguzte9L2zgh624i8OVnmiofDt/5QINFhW0s2ukkC2XIpLeXt7
EVGccM9sO3UWCEehmI2b1O8sd5yEkAEvhf+RjWGr6B5y6WStT4KXwqCS5D7yECoD
pb7Kh+T+uwcRwxGTW1Vt216pOVqXddyLdPSCD8HHIWXjzzm8FjtV4T6R5Apo1ens
I6xm75Ihg5f8oO8Ot4Qo5y4LZGYHxg8R4niUJlMDXm8s5kRF91OS4Z9tIgRmtvtb
vd+kNdGnnG/KOcZVGTaSnawNQbfRIqcg2PKYZHsLOjEhJCtKCGxBKlZn0qS6YVJL
/VFLWTzMpy7D0AIkvVivN6ssuqCr6WIW9uNmOAPlV66QjbBS5Fdm8Jd4q9cHVpts
vGVf8/4hc69IwefaiWySo7Avhp+pg+CZwG74hypLKeiOBIVR4WWeO7S1btGtn+Hh
5z3aVSHRVolpDihduEPp+PbawXlDFHCXKEzEwqpg+UeJPuUIMbNFqXPoARS1HyYQ
5b6XV8YL6RaFBqNQChRJcj4O+fjan1GSdstIysfri4PW1y8xjjKUAw7nQYlIt1hE
aopaPW4i10iw3pkLJa1iIKgBeloYBHNgee4oLnidVAGmZyhRziDqUe4x3NQ8hOy6
T+1RGbM0yjeDsjHhNQSkxIwYxxHZFeIZZM0G6607s0KAZibP3e13zj2p4fbL5Taj
VQTftmPHHTXfV3+39zYxnOXpuf/5QpEjn/32j/qucehdRIO3jKk8YwD7/YJOaj+y
JjBFdrJXmA5r4qPXsosn0KBz0vTbQaEFcugGQ4UqCRXpGPhGWJKU5MwOxjkiAERd
gWl2VXF7FE2dnVPeulb7zKBvOwE+HET9iIsw1zaUtAVfEVngNf3NkH3TzODbxAur
CydXV5HIDISTeORcBReIjxlpIFQwSYLnacfguACQPBplhwriAodTGQeIxdymv59g
QfFZkPYzjZcDd9lGsqTjwlx/qKpyn3YIVHbnuKrGuJvgBsoxVkNH4TYNu1Ycd3NK
6Kfs6a4k1b641UjZ6+bS1RxswThEGRNXBzw7l7hzP3oYHGOuYZT8ZeM2D65scncQ
RfTBtmtgM/WPOEzN8YopoRNRQIVurjAGjulkz1BfxSRcW+nuo2NXFhIJU8NOT2mz
ag7VyIWesIdjdwA8cPbLqXub/pk6LscuqAIATqJnoPeBCgdVOozFVpV92x/Ti8vN
CVKLtulfY/WnQDLW31U9KZc1qJfzbc/MLA3xDTI9VkY/Z5zDV4Uc7sOMiKj3n5YF
ONsfGiaOFXZS6PaRN//ZDeGa7QDYBq9VgoaM8sx5zUpVQUg4nZqqScoEkT+SLByA
cixLl7Qsyhyaaf6UM8un1JTKV/1Ee8UdMAMB9OtsbmuWgiAjS+m/iWSTl2p5TXsQ
GVW1lj588yJXZRlNshtAHZNSr2+mI06QenoexLD9jfivF2NlMjJdqlHsvcoibZyk
tlkywW0OdVX2HN7aAatD+e9zhwhvXZdqcOItXvOiVmsuNl/kJvhQiuRPOezBLj94
s9QBYyDFKL9NGeahgYgnwyeM79w6rlXiHn6HQo3jvZEP/OFiZfeXthIiELU1zcN/
UQy7er2VJKiuWgW5kspIyl2GOOT5LshQ+sB5XR+nazpfrFDqDPh4l97k51gI8/4z
TB2D9x3yRf8BeyzQLcXya4b/m+k9iJShR0p9n30tWa+CapOJ95kRjOo31d+G6xJ0
6mcDm5Wig1NbKFjP0X+zSbaMC26GFOASpCy9b7aZks5PKxVVw8Nwnd+zpPg6C72g
EOHTL4LsmLFtxe16c7QhgjGEXCV8kVN9L/hopFv9d4wLcxbVyT/9udYW3tlDEgxV
`pragma protect end_protected
