// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:05:42 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Bkpl82RJ13H2hcCcJtCFs79GVggBTGTUSh/vM1RUXFoQzphfJma19N8Bxc2WFJjQ
c4ipxybVf5MW1P0ueignmUG/GVrJokEqau8qE84Lo7h6ZclGqYHfu1ZIAkFWDS8k
BEwkTUg1/+QHqc4pi+3dYKMiKP50qU92WseCYkyXCeA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 16992)
pJu5YkmXlcHcxGgVmNpr4WOsmDLsNZ8vTgZLTBBoBpMk7WhDtbNlrgNN+MBWLwdF
qK7GgjBpk0NG/fVv+jp7xC+5tXGb7HmULkizJ2miWDvQ8mZl/il1iwh8SzFeMfgi
hwAR0BFoF0WtulCiPinY0ZukRpZAa5zBBMpISuiYUY8V/pO8v6z+EnWORsVPubml
DobwIvhS/pegthkFYtnJb/aorzqXdWbHUmsKQmAD0RHczivatKU6BvvZvfxNZuPm
IwSq0FyJJE1RENyNlkGKXzsClX1m4VLL2WgXHCqndZfQ5RiKXj2obDL/LZphu7PP
7q500mT1aGESoQ9BVG/YrU7KG7mgZVa80SAxYX1+xJNfhKa35PbaUAxvu3qy8+YE
+1kp0FlZwqeiQHBuMGNClQFd061Ul/hL45AMvNfc5hkSdCw6h0hsG2libLZEaWaT
skEFh8dajGMZIBGrH8AQ8wXSp05vyjr1rwtAy/2eIJ0hZDG/wKayIcMescvaclzI
/EgpUPMaWV2MPdz4HcjtljuNHRY4qdo22wFiuJJ8Zz//JUaQ/FjQtvZSovzcXSrt
naZiOBjxBm041WBYjLxX91Mu86lxrDidyZYMjw4pEtaWJA7lbUsSuEmJ5ITAV4zE
bSg8JNkRnu1Jg/iUedbjaZYJ3naKsjU128UDoUxhE3S56EqVz72YPM0+TjjikC1J
SEpN7LF8JXhpjaXzDkS7o0iz90CARbizhtjEXLOAT8fuqeqgeWha+1k3I1UlWdmZ
gcndOUvFhHA5PbUOQONjbOgm3L9fniaY6J73GgEdHBW2FuX9n0i2f01TfZc2itBX
NxFb66ehjJZM9yNjpG4yDMb26FxMCK8PR34xL8sikORfffz39UYK9GSGO+eZXoHx
E7KE8wv229TFxly65rD9DZzrJJED8YagoZRwJV8DdOO7IDddoPWIAaowrlLmCpe4
4FZjKdvuu0RR/LQqvzz6QeBO4AzX/GohtkqGzmUNJJ6wD4bgr5BVdmjg3mzPcuzR
0WZ8RW1WKSZ5i1eFZcQoywVKtfTlmzm5ecJ2a/uwkjW5SWzB/aH7xI0BeaZ3tjCZ
qROfKDo4ymzUeK1qXwDhy/HVsxLp87GWlFuFzLgK/3mhmQV7l6PbaKHGwZEln7tN
SpDGfwNoPvc8hNQggB5OwVHsA/1DqX6URFrEpdnsCZ1XoPozMfbjmvv9eNpfUWH1
vugGXvbLIyFOrUJcte3nuOmQXTvXvpuYbi54aN4Z00nmPHUQzFOwmfMD6gizq/la
uKvXrqZX55tG/aSQLqk0xggkx+k1Gz9oGmFQC+sTLzcI9u1EkeCB8xncqEbZxqfN
iScJLGphzJ6sWtDdSIs2q1aeBF5yIJSXz7WLAKTUPUSLhpLxhw9ICvtY5YoVmR+U
5+xHL/ahCxbVwbFWYjH5yL84tzdkLT4eORNwBx6eS/eqx6+GBjXdjuwO0gAxwROk
ndM3eTWgmYu2Xj8SsdY0VJFGgucF3+pPgf2VJ3D7loZ5BrVDXaTsa3Q32fhGligm
goiiPtL4wIS/7zTFzujFq25FTaUQf0WGs/Z6exOptitRfWYrNIENEN2kIHWS7MqE
OwIV4N67ti0239fqWNWGK0eiuqNE2MjuTljnBTZ09KKVup7TtKCUqIsa3cSR9WkE
cn6uKLHqwz/3seOUEKxN1cB4Y/k/oVPXbWA/USE//qV1yA0hUVDBtCiUpdU7qEyl
Xxpr76sowoAgNHFLGu7fMn5DAI98WWcMTqHb/W2dMZH8hujKHrjEXZ3e12uIy3y+
pK4zBTr/XRT+zvCxeBEmw/p+J0dFVcWoIUGy7d+vfUiWhh4ElmkTg/waRd4KqzGq
8z1QXcrkSpjren8/nUv4cgLkvmntbPfDpAA6QvgVdAwf4f69QcHUAJzsprUHi/5G
xAFtngJPyEWrmPKLuVsrVX9ug4GNVTktwhwApL2NAVe15SNEcuuF2ATd5dUEWwv8
chJ8zVJgxiT8rIzYw8vvFNEPJUy4Iw6ziKeC8/Fy58ioTqtAFHjJ7B25vyGmBnE1
2zyjyqypM0nzsB4aKlPxs4eePWaIY9vnKoja8bMkfw5ZVCPTN4HbEpSkfmJ6YSy+
4gCYNMr66kyWMbO8VdXE9oRlMb24xhc+1cNSUEuHblzvgfuBAK6VHIMNRAWHJgg/
pMN+7rQreT35lLtJ0yksic9OLerkhlLwsKQ+8MdfUBfa5iBWncl0ljtjT7WInBV4
/kiYBYa79GDIA3pY5LFg1hnp8vEXT2S2kAoUsl91IqA4VybQQx+fotodkVLAwr4X
tPJL0TIlW7yAn9rVqfBFGZ9VXCbehwH2iuDVh2PL2TsfM0m2DbRYnfukn6WzzHQw
CNdwJQZ/pY1ogSybYG5KYb40uf1ytystPrTXC8HNYAHihx7AMnRIYOtN+uNX0ubk
8z0a7gtdfaSuOTeLMq5vOebjIMit5TUhNLN1nyYyRSIoL3lNYhRJF5/oJ54YV411
JSHO3q/WLPevXdKMv7FIxU4dM983f5XXNFcMASDqakBT1JouR74ec35Fk1fTq+U8
Fp3hG1L5yyxTu7ZkQe8ycfjrE4gNC2KqjKhFg/xNtq5UJJm4cD0z3xfM+EX6i15r
53EaDwT3TOFSs9k7w88cTGa47BdXL02TacsZTAOaUCfN2fEA+30WmuCTeRBkIgym
TN7yxoPiWFD+iwI+Dvuev5lUun+YvDsYHbDL42dc9pPrc8YZ3ODeABD9ZoilIeGC
JdilAaM17kPgJi8Y69uvRiIw4lOugdwFWPt5GzasvZIoAGqfWRZ9DMNfe+kV8R3c
XZl/55qD5Dd4odcsAqg00y9KR8PpFnhn1GMii+euvtt/rTEYw8KOhdCqzF0cE4tc
s2HMcyJjBFEzxk2X4S5dSxpYLsG34bZVfLV7UjxyWLKxEcPM9nbYONemUD2SBn1f
S6KDGzY762j4HwoJ3XKftpftTbPgPPAZEH/OFuYsAD4Dwr40D1oj2iqICKM6chHt
emq7nI8R128Dlz4vnjpBZ552mkoVzpSCAGV3lAWGClT6uLuWwuzOuudbrj6qJ7O6
M3Ja8FV8uqQ4Iey8jL2Ze7YkQDvAES/Jsj3zPmwqhrLWACTne055bgSFqg3ldnRC
sLZIPepkEUWseGHITu94yvLLWhCJe6fPgH7aVzRpvQKkP6HFQTt/mV04gXyvohe2
5U3SeC7ptOefZZuMtyfLZIAWOdntAUeCb4pl5n7+2bZnMbWlY3ZmGpsfI2fXV6il
7kPbjTvqV7oVdWAvvcfo37aIh4EvAN+E7X3xqSqsdLCWerYvSvGdgfV9h+Dd8Bnk
jUOH2DfX26wc8I5AsubV1ULJ79ac5IJB1X3Z4EIQ3lLmokL9gz9Rc4rOtHiLxfLC
k7Z5xVni9kWNNr7ZrzgHiUKd1glrFPd2hwdCeB66nHgwipzncZr8lLdyqNhY/2t0
aa3ibvU3P+6U59/Uw16dATFXIgLxyg1CO4lEnLULKUfbECNve9yYkqrc4jpLWjcS
3IOlUZGC8C4AQYEV7ehbM174NpIXIpGPVJ4Bzv+3iWMNg+VoGKsJfBQoWGI6y0M4
AN51M14kn//bs5Er1WiWrVEWrTQ2ULzdsXRkxTP/S2CqE5teUKmAv3yS1E6nE2Mz
ARD6x7kbDOtGySdkqvmPhVcDV+5/3gcDVj9D2KrSrqNNsy8LR7qYEX8WUmcD+5nk
VNF9BYof5hObIaVWqeA0Ejk2Pjhd7ZJQnCdO+Ig/RbI07w0tIwNLvzNpLOFOU+tA
HrjBSN34o5wr2UZjVSKCKHTwXikJ1VTJbfE2o7JqqXPwbh6ZYbMp5XPWLVZCO6Dh
9PHifJZV8915BX9coJE9tq1MzciRhncCqNxxXissLQhNTsUcZ24CyvuWG9sdCKbL
Bbz1EGtbBaWqHeOvpVaiDGc76R29ZJkYrre5H2RqCUPR6wnJEnw0isi07nxUuUSe
RHxamBUHxVa3W2hzqJoZUdluO3a7VbB7biTse7DprqkSVOMqoMVfuOZV0aGFlStI
826l5sjY1ufjLiA/ArGC5uuw0ULCs8H+9LX+6SAyDxnDOyQ4PTVY4vzHuCdjAbB5
7ETMO5YJfjtHKMXeediagls6MfOIy555KnynObEsPT1SVTrIsEsbHVhg8Twst9qQ
bddm+7UfDApKwC1KKfMUsCny0ZN6IfIG5HsrgyFU+sJnyfteBe+KN+YjrVSFeuM5
JAr4cMKbwrLmEtDHKvtAlcDnLS0voyKAfRGR0oXEEDyVJ+KUgrdgXGnynqLnxP5W
m8eJV+bpVq/rTpSxL8emBxBj9vjCwS3tedDDM5u6ZnICIiAEFVb6TV4M4Xro+aS0
UXGVZGUvlYJdUkxp3gbc1vFx9J5GBViU9twttkfi6khk6D1uNfFQMKz2uWP/x8C0
8nQ0I9M1rEGzP42uJl4beaiKy3sEcB81+yXBFDt8ru8RJ3/KWhUQxZs0Ttw87L/i
D54WbZYuJo+5lyH4tq8TfFKRjFpte9tsMyPmbXROqw143BoSsDVPrQR4JJvqqGrD
aySB9gDONa8PjpPgzKe0uMpfKfIw9Hs+orC8WnSsBMMfFxrsJ0HvfDHx+bBtSgJ1
p40wxpyM3XlSbcJEdUuI7en9sQr7medNbwydKO8rWxtSTjjIUT2CKZ+ofY2vc9Vv
llrmo+iUAEcyxodQsZxY0cgVn7lLE4h3gKryKkp58lJICpVgbcGw4z38uQwG6Cn5
PnJpq76u/thoAj99IDzKfDZnulVdg+cIGZaEo5YRwiB6DOpYuR9oAC/4iE8wt5fI
nsa/A4GuhTw7V1C4AYMTMJBtyYRmhxaTd5jSkQ5f4uIczJ+PAaQyfvudBZapLMGI
35860Q2Mdge8+G25VSki6hNKrHqS5UUg5P1vpVB/V9HXgmpTDvd2Wjn1a2KXR8TM
UsiBcGvnHiUEJQuRDPBPwu/QXgunx6DdxUgE0M+p9ZpN2Xj8ZrnJ9xBKEUt2RXCL
JrsB0giFiCYBeCZ/O5PoTcdIYzV7clESgybXWLlQWnc4FYcrHWy8QEEtso1inNrW
pmo/UCzUlqIMu990N+Cu5lamzQtnqrGXMcTtdT+NPeEGZ8aYkUGCd6IG4koaJMiK
cojRInp2r90Wf+oFEAyW0y0bklfrcaOQgYrbW6yXww7ZmBYsdN8KUPG82p6tvpMM
hcluuetwcnIL+Wd9pl2cs6bruYavH6J8+a0N0KC7zi8tVcpNG19MtFWoBrRHX0RI
ZSMViJnbmUPhqkCAOMuOoj6ni4gzBbxKq/+P8k7DH0qxks+lR4MtPNO6ueo9Mj2l
SDdjPzXeKBd3TK/v/NcXkUjA+1mssKRVMqiBkLmisE01SQbkdCLDnDSCX0tncRVM
sV2XODNkyKIeUipy8ugpN3UZmb5W9gzhF07SCssqCYR15gCYhpZ+uUPVSheBY46M
/NjCCMr/+hsjftaSweaTT0LRP9t4NoJxOvu/Ut+DCR7miPHPOzemNbQH8+C/dCsh
oDaNOdRc+WqUhO9I0ctFfOTcNGkZGNXdT5C067SMkdeORBpZPPKJZAhVLdwnCSW7
sLAmzNon/AIOSfAzSNQ3orYgTQN0fptmsniLq963JAFOa1e6QBxe9+I5m8Y4yWvf
mRV24znvsj3G4VeNGp982K1m6Js3j5PycMFiAGfkakQqtbL/dVRGsnGpnTkpkft0
itrJ6EHOJX8kY6qY4oUVD80QYALJLq/5iw5YkhmZB/+aBdzJDCBE/Uex+bWN1lzE
NxhQ5E52hagnot6RT31ZWuOuaT+1YQTxlifmKKg5ffu2SuqnzEnw8h6t0skbduiS
JaoiMaKqfyyRG6ACvb4OqB4ucOrwnvir+ounsbU5iTujneD/Rk67EoFdfwIgch0y
tUn+wQ5zAaVRc1q/vYWUpDtIUNwtTL0eJPmOwfY+rgNoRQ+lbdOqXE1BOYH/xS5T
jNBUF2NZ/WIcANpRw1iZweybUGib6uJmVD3e7u0tlMugGa9vF5I86N8s/2Q4oJgg
K75QXBIXujy+7YPxjhXgNBK8aNwNjeIGCGATwRfOQMghxei7325HhEbztD3q3dKK
Cgeo/gAQjacscqBxGdfi8MsgPA5JacvFST6FfTDXFwsPZZEJS/Rgoj8arksYCACT
YH/RKP5Nnt36v6S3Z2hmHbnKN1ujIisy5mhkQAOTO+jw88qjrWGHUhN093hX+OFx
ev+/1QmjP3E/P7G3q3glxrwwxM2tHzvJ4591UoujWLN7Xtja9xVB/TaSe2xEJtxp
QI/iiO2p5UCBqbJV3SmruCn9rpbUqU4vcALuS2ilcj4v9PRYuqOcB7OtvTft6S8y
mBXcCGgJKwefPNuX/2GBdbY5hq8f9jVNx4Uc0fJV++tXTPRrED+b3h0wbiCqWZ6r
CO88iJQZLqOzSE1CSI4O4AcKEaqwvS44QFNjIGkXHMCw+owX12tMcyCKfne8Dt3l
WgzLrLVndvgNILh70GyhPYEXZjFR2Lh/KkPcAF8ozycfo3830ng4eKtmUacDVfF2
NdUfQqYVmR/O/R3eLfwB1CkNcituj2bnOa5uTXmGQInZDJj7TQ7Qb1cVffN4iYCT
oYM+udWc0mkUmm7wDsp0bZybgKx4l9brFxzc/rqC9DSL3n5piViej7Yz9HOW8MNd
lfoFN9SD6JDolg9V+5SC7kKafkWUyrxKvUZB2Lekv1q+pt282ZpFknFUEpe8aek5
nzfba3YSnXGZSj8QZKhPp/a8AES1EPwvi65c8yHlzXeoIZtE5qct0WpbLHJ4yr1E
2pSoSrJYwmA+FdCNqfxSLwuk5lYQuYlwz0NtntmiGAtcb5yN2dO6+EYRwRHkokan
MNjG6ZoOMKfNT6W1mHVSuxWhAWugkKWthCXGZeoFGEoc2P4Ya2yBGv7IIEgK4fZ8
OXB0CbF0dDZl6XZ/xrG+AQgdv3YRIt+8KN1rdEG7M9bls2YxUVkw2aQjKovLNtLl
XreM1ZVeBMZuiWDz1azwX0foCMw59jqDPl1wgoTGX2zSWq/XddkgcoVSmh3HI1ax
cue3wPqVjhFi3joDWuuypVg73/4FlclHnkGlB5ww0phKGtEy4nCzjjIHaUwtfGAg
L476uWEcuCEuvGkT1b0S2zv/ATdS0VQ88x3uK3XiRPGJOqaYrYKANVQ7Z7kpHi2E
5qYqhvZEO3P2+Kmch+4UfJSAqDEEWGsleSIchs2aoKkTj7i4yDTmRRhTxRA+Qyym
ZXk2pT/V9U1f7KDNHLyY+mk0aAGBqqerttYjm+W5DXX3U7oTVQ6lFgpRnVh8z0Uw
SOcQKxJ4K8SCKsYV3pgCz7KBdg6+f8SqVZdPBPw0BnlSLqC3bYYOsZ6q67cITYv9
lqQxOXM3l1iyTLCF/9Vxu+EvuK9roCMsDiFiFcpapSrbCd9yAh2eBGN/utp9rrdm
iEuI5nO/H8Mnsg13n9Jr/P+54BZoz+fAQVhrMheCBFeWVKZvdD1SYv/+LMBxuwmn
ruvAn3vu0CR5lCKvOOKP9h2iZH7JK7FF+N18vGweimAgVdsDeVbcBTmFQ6zA0BQh
RyCbznJtmCGa9Qdk+tT7M/dKrB6An7UXphl2qTcCDTEVN3aXU1atXpo/WvzPnRdK
NFTah+/lnEL0M00QHnQ74hq0jhNQEV4IbZilZohDee0lBXvHkmTfDk/ze5VSWw06
Y6QiBOnpMdnYSZ56hSMIRCawt2OodemejWKiZysDdcq8fOgZSamfCZCc+qmAGFZM
xHwaf/5XLygDBTR5G6C5Ry88CT/jwlfTUVstke8Zb6d0hIuIrWeQNlpDinjkf/qx
CF/HSP975A2P//hRWt7oXZtRUrt1nr7QaEMXg8Px3qwtkbZs1+jCjv3CPLIsFIt7
9JbkJeNtk8uQ0hExZw4BvqkbzGaaIUYZpCn6EzX4+teZoHyRK8XJd6mqXfckZgUO
U95TIygsMgLd7RkesNqHt9KO0PrhI7PV58WSmEMTGrFsHVzFiLI9oOHfWVJOWlGk
HleWstBJ/KU0crmpprgLdUi+FPIdN1iX4NsngO0guRsuhYG5Kyyp/GNY/f+aEz0o
/Pe9nBYf+SdAnpsH5qS660xgx7f/wP7RyHZtZKvfDrmnzknI3DYD1EFWJN6NFjDt
sw4MpA2nxzPyLJYI6WmBDCUlxlbdqFltJTJGaIdJxS9wBFfAf/THWU5gsxXvQoBo
BMle5nGoK8B0e+X7UXKm7Hlbn4UQyov4raOlwJPMQgXKB/7u50mnHUdHB8+dLbE2
+pQCiBtanSj+J8AT0jcxWnKzkaqb1y+Ey622V61YoOy42KOdZHBSER9foAB2kWnR
/sH4iOe95p2KfUoyWraQAAy2+OjDL9tNfYvP4bYoRUJNKnpS6g3JoqJsrjmAp946
837mPtbjWAmKc54fUWI0ylF3cR1NKIBUvM3hBSfALu3o0RzynyOX2Ui/2t0mk/Cx
hznQ8Hd7tPF76boM/Wilhq+l3GetdF0m6SDVg97oWmeqcI/cM9d/RrZRKLYx6Aqy
7DgCT69IrRfaMAFjJjIEMaxeCZFZ3ZhmINdu1vvxhj4VBKyJfo6URgKT2dYJa/LN
zdWoWZZ0zYgySTFov+lVX4w/PpfSFaR+/RXA24v8uD+/SFoCKcDy6yT1tikN9LvW
//51djG3Pe2fBuuJIXANzj8tozWpLIaJF6bsDodP7aE1eZRBG3HOTNh1Lzn2+3wH
qXTsqRWeC7mUSE54qr9fSiJPRiHByLBYQPgN/II1Dp+jan70wVDVEhJVczrhRY0z
hz8x9fP1EwDR0zN1YA4nsGZ3ffMS6eF3PePZ1ez9DPfbb2pvEoUjI+eln3GnXGni
8CL/8S12LvCBYqELEWMR7S2pLrIKpEkIwoeHWAJL/Vuu+ynLhmO3xDsxfLJF+a6h
4KA2j3qf0O85hsCvy4slWKhTBCl8013G+OLZrcr3Kb6pxIyCyBD/S2rGsVc9W6eK
7+WBhq7YpGeJppbeLiXzbIDLM9yRR+f8QfH7jkVcU/SbcbeH9wLeL0fdu5VvPbiE
q0D+7wkekEy80nK+2L/uRNQY8I1zIU/o8sNsdgPnnBIBFTT/wbEalPqDaYV34cy8
0AFVrKAOc6zMLaSdPR+0pWhbqPIAuDwC0Qz3VTAgH0C60r4SeXYq6+aM7kDLVNwr
b7lCgKm4EeyG92S1CClRnxBkeO7VLkvt7rx9J/QzR6uqtHfRJFXZX+8iANmuD7hk
h7jqdTj2TQ950wbe4Pu3EUuiR0xigFgY6qP1KodP+I1j0KtXCFS8HJf+U6SYOTsb
lwtp9rFHHXsucnayUWiPPjAIAmPuzri+rHHW61xec9cbqM95cr5jonQcdnvr3Xh2
+BfXYdlVNO5nV7kjHNDbcRZbFbaR/bQGJBqZMt76u9xBNYNPnITCe578hS2SofwY
R5zxmo4YKCgcxRoA9p7BchpeUmJbMskr+guvbgJ5zeQpllbTXPUPyDcggrO5VWpI
YcanaUMHinBEWKORj6Uy4Lacidsb+Wqnb+U3QfQ7jpy6rFHX/soxmhhMF3FUNBEc
DYULJTpdkKtYH3HyJD+Fov0WWblRdA9gfVerks9t0RJ6M4gr3cLpMDd2tkJ1OgqU
L1F5muTdwPjb49lb0DnL8UghQKzF6qIVpYxDmCLZk8aQaBioE2kTCANjMALs42EK
B74lfQuVF4iSzm/ra920O3MmFHOty0qhrIp5HP7nKi7QC8mkhCX8/zMG5oxltYeD
NrM7brFP5QEoOQNmuzRbreIg/mkmhkALKGWZv4DwwNSP4U9zZLc6SzLVsMfeSEKH
2XgB5Qxa64NfeZaK+d2enaGXzne304EAhsVXRV+VaWQyp2ClAC7jWMJ7w+PnELaI
uJYv/+gf9SQM9VcHYZ2Of4AamOoa02x51hkCq9i4jift9K/ycovBWTV1Wf0+iZHH
wdvSfghGV8LsfpgFeEjpxkEHbnng0GX6Bo1idECSkzodr70TTJaLzkVgmf7qbyJm
F95N+c3Rr32MRm0yPDFRwqKX0xacY7jiGAW+0OTlB0XJAGR9FUi3mhx9MgUPPT7G
TY0FdVP/RikNMSl7sbRDm5PjhX/qpJ1+alebMa8aM8FXd8NDo4dISYoEpnjGdKeo
G2Krr9tmsjrnSPjl+Grx3DqTVdqRpkZIaMUfexvQrNbHZhc8gYVLrkgBAIhgHq3y
uj8C2Y8aaklnOpk2Dh9h+Qa3sAAfjv7SIJ0asdnE86rlr4UmYaQIg3EySI84nTcG
RaLz1n6o7kZOzGVm8ZkT7Cqf7349hpyhFlDqBDaZQz0JciByKTo4Phm74Fh9sbRP
QxjR8Jdy06k26IU1g0I+h1cQLZQUBKaFbJ/7AjgclA1772jdzbtuW/vjs6YAq3oh
sbLHtXThkKnkZkku4CnEd5reiM1Iv59sYkLysMl0ByGfJ9Zev2+9cpbkxx7LkJi/
JMXK5KgLBUvbRfDOi6rfdILOzUxBWP4JgvwC6CzH2P2WcX80KJ4ueGFqo6myrGFQ
YjqcEk3402O9t0l9oxa7gn7Kok3Sig2QVRKhgGmtHKAj0iOHCpsodeAY/VG0Lrcd
9Y8Dj9ndJs4o1kLZpBuL89IZnzaMO/an/W/671DDNHvNxGayUM7S2xQp/nri8PwH
e/a2KJCTvffhBgF5wClEarHBAHkqnqLru1CJkne/z8sqt81fDZORdleLvOwuzDn2
WAJUcKjBwnLNqEFbzgzxs2261hj5C7iYiWXenXOFi3z48blwxU1i6CqtfKjIFxo8
OiiQmTUwuTyTA5rTtzSBKVSzenxXOEoY2SoAvqSzFDycLL5hx53nzChJsIoGfMgP
0d6hOmlruawPeSOsGy0USdZAz9klDorcmW+J5pu9dC/wjd6XFlUkElyX84YHpNKQ
wuMCtBfYSkgocvvsfVnw/KVS0CePqFfBwF53gsYiY6Vq6ZJL/TWgAGN2LpCdfL4m
l6YrnWdeg2O18SDBwpFerNOJJ4SDTyUr8F0aJ3qdjBO1O/daYJoFfQEEJTYcqlMK
ryws/9mDZ9nZYz83Azt6/SDQaznZ3lQWd4g1ACa1AVmlTTnzxxpu3aQydTUuqUp8
7irWMS5TwCv2WP/nr1bllK1KBQiaS6AczNCXio9iSqeNy9gTbNGCfJ+yeuTG4SSm
qd0xG2h5M9Lwwc24dWIQodl0dL/TavaZ71ch1yQwauiD+ekCXURa0Xt2n1Yix/kJ
4SGyPjqQO/s5p/c2wF5mQyK3Rlc+QdM5/c5o77cfuUPuMcRvIEjIbUEjjFDvvGUB
dovw7rrPCjUFHzQ3OIopqNvK4eWUmcBPOwrh/4MteoE+GxCkzPesAD/J0BMZimh8
v+/cRvT6WlK+BJbcYtNN2XX3bu2xEUpmZ7PcBJkL2+e/Uf4q5Ce2ZC/9XAe5PF+g
+0NlkkLl5oxkbXXBQjfLXc9Pso+UTUtKkKh1MWP7XEsZX7mtBr59rOh1NSqpZsye
oZICKNzyZINAdjH1vrjiSo6dhm/q0qoObmgJEkeI9wwk5Y2Na+xDNr/ct1l0hO86
DWGmLUYfytlpsU1uXy5/vLMnpHypqiy3qUtCI5xQ5e55jnCR2RXdTt9DDFrpKgvW
Y8lBiUGxmkqbXzInHWRtau/2RsPCz6XOswMDHJlhr//PGBHxRYJflGWMEwgUwABB
YpaBvMwHtjc6KpWKF3nrD8QNu7TruGIyUvDyqJkXPYU6SauVpMJhZhOykzuODob8
YBqKJT/q7TyeJXhzxZBPtVLVlN+pvoZo9hTA8r2T6aIdmWrYkr8sa8yxpsOyDFuK
n+pccbJhZRpnvOqCyNLVXUUpR69YV9OtWQjisuLsShMKsDwNnPy/+ssLxYX+a4CO
AeUr6IBLfK+u1KX4P4rq8qbP5ECphE6/hM/PFjwQZangsiUcOgDKZtA03HyM5Jf+
QrR5ATzNKxRSyQP82mtQLpBlGXQXA5qFlEq+e9nCuDOP9I49rlF2m/As0yEMoiZR
ftpdVykPe1+ENaVUrReTDP7fwbhvx7sT0cKgVfoa/4roNUEXq6jAuEnrdj0Hyrdb
KTLhMDLVM0nVLl/HFt0yHE9nQpVq+xMJTOwXcY+hzS0Svh+vvme7+F+hlMr+BMbY
ORQL7tcUeiWWDBvPRv5OJu8DPoA1uzLMAXkqKtNF1M/RTgkkGqbdTCVexToFHkCB
8BmxlwGjFXEPWGyfuyOchShZl1lU/Aa2jTiNQ8V0WEinjkeTbR39dR5hSy0pbGsj
8scKDJSgHDzTTxVzAgH6Eh0cbajriqi+PZMWe+kXfy8IcLAKxJ2GA6MMsZwBxvVc
L5cEgLZ+cUO/GvlSlEt/+AEblem+oPPATNX1TV6t/P2C1C4jVELjtyKIhZDm/i4A
zqY0GUh4wD2HZ+4hgEP+kBo1P6MIvTYDyFVD29ff4HsHI2NTg7x80VJikp22IflC
/uuckEkq5ZgAce6OaBnvl/koE8k4+0Fz8meZdZwC3S3kDYmhThDfosuJaXdiJg6g
mF5ABfQx2X8vsueAO9ddlrIHcelVux81urQdEuiurQM7zjxX3onGL/YbMzu1gNht
41E1yB1uHvocBAK+Zqi15uB3WnNqI3jQkjGkNN9hGcSqwkAJ308flAxhPiWAa2ez
MnnI7uJx51hQm81AaofYR1QKSqBGIUw9AYL9ckOYmJuxWGLvdPZUu0pilCqgmjaN
/favMtMeTCzfShHZvxMxGwtY/uPg7VxazgpUtEWOVXGdBZ5TpfLGvoh5CLUVNlqG
sNG3xXxtdHeoKnMD/19Xs+hjU6SEg4ty3cNXAzjA/U8odEh2bDQFfpVAKverXbuJ
zzoG40e9k1hLEfS/xeO65XKTIDcc8Q4W3ONlX0o0Xg5Tcfg3v7g1mSZKe7Ht5HTn
SaQc9rZLC5zQXoCbE969aIqZLGUZVoAjjvdooGSimqDL0TTWZNAOftBdCfycyVk6
2ryPgJsaftejlc+6v70sewpcYawAsS2n94qbzfP6DQmIfuuOUKxUQ1L1VMi5/IeF
cH9Qe1RufxMg7zWE4hESYEIRxU6NlNsjRDt+Qhq3aQ5RUIut7IjM5ZWcBMXPQWxr
txFdaXrDNAv2i/fNypK3V9lT3f262UwrhBLMbHoAQvMt5Q3AjZTu2wfAqCeD06RS
BhweseQXRcq6W0gPe9jyK4Ai0XVStDc3BGGMJOj7YFlwR24qmIL20fGXaNTlRnTK
cd/1pjq1oWZhYKtE48+gO1x0ZEXHwrBALTt2pPvxPgFPGkknyP4TVwRhC3f5UkH7
6PEQuS4y7V4WPgRrS+r99jmVfaEkf3sPf8/EKq3B/S0tqAUKr0CarUcXqBij3wof
gXWoeXbXJf7HdGrSvFD+DuP076hPbYWRoUIPJCOXPi7E9aRkqtOYjw5a27NWpPys
2AIBbBZu4KKiiTZgB8wwXU4+O6MJ1FtDfv1X1B1YRgk9R0yH9uM2DqnIIzPe9RTV
4mnhn3GiFdizyLUxU/CzTBqef0dtdabcWJCQ0so1eWziRXuVkLxF0tUxoqv90g8Q
Vfxl/ptoJobu5QJnIu2t4UfnO42LnJbD92OL57po++t+uzALk2gQ0nwb8Vw9k0x1
dmvDQ4lEJHhIVD6LilOezdyqQvSE1pqj7rDcwgTsxr/P8i/dR7nc12+U9r2cnMQB
jd3H6MWC69SPi2daAzr5RXhNtxp9iGKVK7QvrAeGmODxTJ9W8deHwxvMkniaNP0Y
wL4Uzfff+aa9+fIZUIo4rH+vWqNrNZtfyIZHkJon01nky0Fl+ebQ4y0JdexGiLeQ
J+arGK1hjlQvu+YbhCKlWWWO0p47jv6jM/XfFjYAXZqtwUb65xiQUtfxF3aPhDau
2AZheeL8Qx7RMYR2OnAFKfvEybTUcVA7/nnu9lManYt0GSYCIMtbQomohuEw2OXu
Ji56Ta4gm53ywup5q3hKcTsPBBbVStEW2GZO6HpeYjNaMYRxszhNJSHCrmtPZNYk
8C0lf6EODN4ruuBRqd02upUvoURYVXbZkCHTjzKEcwFxwHn9+7qJDzn+GArnp7wH
L3KyK4zE/cI++R6U8JzYY0/sVsQqv6fDskiOC+S1XcYlVnctKHiDUi84iYKTMuFb
SYzXpkAdGD9vDe0S1FEILj9xJJ/Iu3BfAvwoKG9gYLbfQVS48hobXT/aogkZcM17
/PF5lUGd/O2t6f/O0uQbRtwvbg3Yw1BSpQOZ4k9p6Pmw2OwXi2gLwiGGVa7w2ico
oYmMOvb7vavXMpf6RNgPzpqJyXQOmMHGbF2FqXrWO9ncRmyBONwSmqH77QDak1hh
/geMEEtJIeU+o3gVBc65aZTBbQLyjEJ785A3HNBNQi29Zk0uFaq9gflu8tltiWJw
qrWe35cQ9srnai4LVJ/aRMAwsvp/n6rSUWmf4mvKqOo+PfkcJRxIg87AkHpXkdHv
lvfas/WI9BzWFCRKGlw+GmXtkQwmwX9n8rgP0m1FUxHsHG8Pnw5Z5ajDWSA4XfJg
FI/yQteNHxXaNNUGO8VHH/1QRsV8ZimC26qF/kAp8EWgxUbDjBv9uDzIzeavauHL
ggj8gJPEwJiTEiHqgQ9nuLYXRsQCjDU16/2uFcUd527a2SAiJWcl9doLTiiUX8Bz
0R/0GGgflglfwuO3amcYmBCBaa6hMVedL5FpQyoR8xX/T8Q5WhWIRCLvSfl3q4Im
ETaXzi8lue6KIUIVhVRuEQx8dva5TJKz8Kkue7+Q+4aZu3Gb+WsQ9N5lLPwbSMuY
q0mvSGrpvIVOa21WewPsuIwNvJxALV9yZWm6wy4N1u2XJ++cm653LJRCulv/fnlm
gUDBXXWBJVwatkIfj0ZRQAsUnh34g2SFfFWaSU7+r4nIX31DUsVymS+SJi5afvx1
Sv5s9BTktrdWsEkgsnYGQsvu0QBYlHUg2B5Yp35BF6tfFmYq1XQZkfXfkcgDYQHn
GfdCkkoxJ68Agokxaq31wLLI8lYzS6YxLUiLxXYPQTJznfSTxeZGeJlUAgdbC49B
Ky7B3L51BqibKqyQ/6IK9bETDcPXH9mIlQiPisQw31PCex2PN4AwP/qg2bNnO6tG
n1Vq24nm+4e8PVQSEA91UX43pgnGbLdt72iCQx5LevBFAbUAHjDPWQhzcIy2zj2E
2zsu+LuXELF1FplVYEc0cd1pQLyrdiMAq41zh58BWy+IMRRmWhQRi/IhntQZ6WPS
imLtABNbha2w2RrVIbH0Ua1sVoA5E+oy49kpH74zkBTZqAfJGZYEvc5GMBMFmAb1
wzzWXqnuaFpAoSNkSCPmlTheor9sRwRSyYB7DW1dtSCCnS8V17n3V7UW0jWG2eNl
sNjzhCq98jl5WzOXA1P9x/Fdea/Bu/TGa2UgleBXmNYYpybzMKDgYh1uY4SIxjKL
/GT6NuMXxxiLl18XWLNg3oqsvQATQsl7N6jwxQ/yvOZ3u5h1orveW3r+6PYOOvGg
8GPOHC7h5kihX5qFG8wedezLBB6vu5j/XDyKUXDgkOb6ypfZzOo0RUv2YHs43fzW
ry0vYHE4HN+bfgRniM2UZLWHnVKHIoupX96NPEBUlwzgsL2g/VD53LASCJf7Z8fX
9ga2aSV5TLzgIHlCIzYBKT4nYCqntumdZu97I8TcQ3HFbVxUqb/k8Z3pxv1CFd7R
Umtpgi4i6BSk+fIX6r9N0m3cx5oQXqyEFj3Sc9s/VcmSIU8R+TUPnVkJ6f9gu8i0
Sn8HotzjhhBuLlCdJA5H2FokKePv8euw+wdj+L0AzfUPa3Ape6Kvi0GGmQsECvTJ
MNPtQcGpwaHUUmrOJ1DHp7cr3+2HPVEc8G8sULYv9u6AzKkMxRIoCnnv5YzDnYpa
pCXK1/d3OyoeKqF7Iw8+sW0LvwlkSbM+7O01NjRxoCM3r+rLEgn9B8relw4JI/6h
kcxLgB9VOYa1ztKhsoeSgl1gDfiD+H62eg+McQu8yld9VeTYofPz2Vy0EHsqM5pg
rRPBfTRAQVKXOT0wAmTojVsVj8It7wi8jIMFAjrKaf0RX4WoM5Ise0PLbT5U/A4J
ZcsW0qd3j52oK1Tkg4m5HV4Ghj09PkP60srXlVYt4VIGbgl5ZaVIIXh4D7sf5CNd
DI+dBu9KpUN5Mo3TSy/N5bKHLc0yHLeoFJlg2e+TYc/u+3N1M2M4zvlwimOUyWA2
5B/cQeqN68G04WfJlqesUT1C7CFYhtI5YwtkzjTvcd2ESMSW4OJwb3wIWNmVqwk3
Q+Z+xaHkLLIUsHi4ec3HNYqekNOlIxsrcw4gAqgirZOOYSoUkGSWGZgqI5aqtkW0
ddvK4YiBdiEv610u0uWpR+PfPlXb6XMP9+8PlMcbT4Jtj2xVTLYWbiiBd5yS2nXN
3bZY8ZLg7a3V1y3wLUJEnefGUApssspMWcqKPnZiFO8SU5k0yGISJK5+1OjqtCcE
WiMfpUEjhLcFg9ha3JD7X68/vPezPY05/8GyDBr1HgYczWwxPr2T7g97ocxxtCyH
JSl0t3lbrLKXpKlPMq5vjvpBIiqf6aFtpbOMYnGdPD7MafEeTVCUV90BWm/31zK2
nZW9Z1VjpEKy6XK78MKnjiZr11GcILfdwtM6HRcWpFTu84cv1jT2uRgRA29ccD2D
m7jT7+TLwMbcf9UN42r/ePinixZ3aZGVhyTruSh0lWv61GXOlunC7UknfIy7v/KG
Ah/d+hC10nR8Ng60VkKabImnhSsFE5cIKZJdw+tj+uec95+PT8DH4aAkc8B1UXwi
LUrNb4dH+FEF+52XEVLrOEJk50YwewZypVyvrnCjIDGpFNmbezSBqPhDFWW29ydz
v/lxZ3BbveP5bCgi9L5yIMpmLvNgGpzwFKQPCk5q8gOA3+b83DA0MqGFyvAXCLx3
6nwNoe5oUZiYf55GEq0nuiO+Z6BolxK+YgZhgCOYMY3aFmihrHp9YGBroLlPKwzf
BgEMOZDGGa075QY8rr263WPq97hWjP6GKhRmL2p5vLMQIs4uZsFaT0Ma0Z0Nvebh
C9lvvixjgdegCmo6G6A+XkfhZK6u+78VLByjNPMrBeQ9MLVeiWTZC0E8wUKKRuwQ
fA8zgFEERrLZG8DIx+v4J4u+FLgKYO1QIyklv+3ynUYNaSdPm7IUamNBLg+GCFkz
y59LaRtQKPrlBvBx78xdiKDvo5hRPNBXwDNkNJqTt8EOnHjw0zLdcm2G5YvzN+45
snjPCm/6sisdpilwOODE029t0/ZUHogPkgIt2Byg57gM+ewCGPBJyYBguqb1R2dB
e2sMyJnQwm38k5O1p0w0wUiaWyr+novL6YEmPJJH/gh+dqxRV5vBi+XhX5fiB9N/
BxZQD9jrcY+4HEGNm4xQjGtlJupQ+tDAtWxsJ4uTat3gOVryMgbIE8cxRiFfwuWO
EGUs/2Wa8SqBYu6zivQsf75GlnN55RVJA8Y4VSRKlna0VPCZlN6bD5E9evNtxrNW
3M+jr6mYsBhwq//gvmRtLiE0o9yMe05gHDW+AhWUxhjw3rUYcHgcx4xGYH34AETU
5X2a3EQBecEi2+Cwc/66NNYmEFCwt972oYDJ6fI2O3gUMychBQETVBMgRn8g4iyE
dA4PcgGI8ScFGZxmFHzKYlUoD0IlGNqTtJwYRt6u/CiPE2iwNSxcU+1bRCuSsxUw
bHEcxd4jbPJzZkxpXZH0doAKyifTp4vYL7niCaohXYPBUwt6WxnfGDYwe0NXvkYi
1uAQY6+pRmQjD4E57TJJlNNrnOGPfNiEwmn2ygJLLhig/sXNEKJvTXUEizK3TcCS
XK1RNGflo9j3626igRGHQPaLLYsNtuLmGHleArcRr37rnTm6vxdpTHwlJsTP2sZq
vkHqkhzUeRn+M43B0QdhDAPH2twKmQhguxZZzhrB2B31H6WRe2CiCWkfV+P44ypR
/ZITbssIZb4wu6WQz8PdCbETuBbUZLh3CPXkZnVRBYOQ7fgvofKkyfSs4qjZvAw5
KHqQruCLqkNy2Bk1Hv0w+J7Oyglqcyc/jZnCNSC93tdzz87CE25zBqDh6VGSiwph
MqIETv/RYAZmSxPR0VU+7+WjME2eNFeZ3uRqICRYoW7iDpzXH/3KLUF6PZYR7m7d
r1k99L4zYPoWnLA2l8SIe+RbHJhjKfldixyCzUyl4Nvp+v9IVz8nz70LyruIDYOI
TLYgS8ipdt6KLShIGh1xyJL6AM0YGIp7Ye+1V5672yRjdisTNt0tIx8KbU/PA0PI
zQmU8klJ9GlnDtEb9cD2P2vKC/WiA08IfjY5s/siNiwqnda0uxMkidRoAEdI07u2
ipVsC+iw6is4L/RrhQFgggg1vmIIdQQRXNqOd2/94mBNTM0+1MU1Ke2I7wqzfZCb
SuUYgMFk5NYxJe9ptS0dfZQefUGVk+eCCRTKACU65jeSV960pdTUPtyjgzP85piS
s3ADF5JuWe57KFvHNzwC+TiE4BjXp+Ebte2nV2a1WLHiNUhDvhopMYLW8UbdyGEh
1Z6t3Xw+x2MEOHqfFlM6+0vge1Hk0zofMqJT7ebGgIs5bRItj11uQ8rcm3zS45h2
8S7t6t/Mw2phclvFqEyWN+idk/jEkt+uNCPkhqGxgQA0Sd0LCITLmL4j5zLmfltn
6XxeBfMJJbdRFAlyQxy+2iDNVJDMdGJDqf33V+mUTf5MqsRs5qDryXG9jaMHq3np
IPRePH41zAfXW3BZ/0LaHi9mxxZp08P0O+H07bcN2GPZvGxyWnQNtWTEhI2XRuJj
8XFlko3aGIJAHK813FUPlKaHoP+IjSTp1GPxy3gVHnMjazYBvdYl4QBk1G5IdF6z
2l2Yhdqs0wIxQKZg5Gxu/ZpP+XeoyMZ1g2fSTh0p5k9hdJLIYiaHkFV9DW3nTLb0
qZwqDrnUwNqvhfzb6h+QZjFu1oGZ3SF/tRjxVYNVqHn91mHUH+2Dl+iF31AmjwG6
Rm5+iGqBL0nZ2DmSn7wut2vvJzWEFFqMXF3//MGpHEdXq3kOsHYTgSJaoOz0GRib
QEc9oTuNiija7JgFuuRTpNeCyLyiPwuVXi1HFF/o3tIgwmmK8kv5Tdp01pUliwPD
EUQkzoRVdChyKmReA4IStjDi98goyaFJbv1TWvjyScAur0clumDGvFIZtSp5gZ9r
YEHkiEVLb7P8B51XFuxvcr5FqXrPpKXCd7RfjWWA25qnVf9uljy3plwfm8G3rg5E
ifayUnxAuXjf9/NbGiyLlQeFj33Sd5jL/n+8/uRqWfGs2W/m+03Fi/8gG8XhIt4f
qsvfhwZaRAlDrhromDQHJKySMG4yHqZX/4l5FDUZU/3IL7WbKfftUD8U44sX7TnT
T850xpHbrVfPVdb+IXvLh9mYtGuozdTOKfI/3Dn8i5CksiM2t8zvyRFqVFSFmgFo
0AifRyN3Y6kuvdfMyJwON4RF02VNOS6bUHYlP9/6UK9vG9iCL0kiY1ncj219I7ua
fgYt0VefyufbcbKn6OL9rBqisr/t+X3DUdAA+dRp1lLh7FL3GKjorzbff0nIEw7X
MGGc+ZA9uiAoLwi7Gyw72PXCXA3TvmoyLz5fZLCNrG6+DtO9Ox2QoLNhhWL8fm2X
5m/oKLlBxNLqSpI/vblHVhaf6B5wj7oss1SPCoS0JU/mbQpz0Kl2ZvDDNraumuW0
fwDz5e7tBiZNA7kXRyZ7bV81cR2OcUf+sv4rGcj/CEbAC3fOF4HY3ZJ6htirfmz8
LKSchXfrxNSqfFVxdEYro/8QXJFY37wGxXjvktjJPCVIbxfVxyyXF2ZOxfJnJBGN
7CH40qzsvWUItpn2dugExpUt4fWp2SPc44wCYtK1niq/cdRkDncB4TjEQ66ilkcK
ZT78KfhPZXaSvTwghdf6tPv3TtOJrJHIzrMRnZczON3/hAqG8wRWmzLEiSubZ5ed
lLN2qKn+rsGt+Kt65xnQCuT4yOwy6oGradZ/XnajZhZJMLAqcEKh7U2p1AhCvOVX
NrzkPuyXj774kcx9kYmiTVfy5jyjRy4p1S4ItDSEypRNVB1ajDp2ZYV/ZxIHNuEh
etfnjDmJyM2GrBgOjs4bq5HpbXKbDsweyqLi6B9vVbFBz6Mvh6EK+JCGnWKEULqz
VBttRpBPywvUVX/WOZku2B1D6bB4DVq9FwtStkbKloKJgimQVobn3mCK9/OYYDGV
CvE6PSBs1wyG5yZhp24Bfi/a3YXQQ+jjWVVAmWQE25wLvBhpWIe3GmA5oSIWQIU0
fFiZCCEtbic82zbdX1CX/HmY+HpvEo1ZNr+y4zbhWHrY+QxE578pPcIWGRZDvakQ
l83Bod702SXn2O7lVYkwaGDFGHFF5z0AK+ZLbtLcz7aNa+Fq3DnOuSnUdmGMIW7K
5gIg9kgp+fVcT4iy2EA+uV+JgAkHCtdbnigg5f7ok6Orcc4HnXg9w/IqYd/7j4aD
79uHdRn3nRNxtwDrnVWWxhZMqSrSHMrl7o714LriZ+STYlo1zKBab1hvaycpkqBP
YgM9L5u4Z4HKB2esk0H9E/06yhHL2Y0OxMF6XcAJwCVK/F/H4LXbAPdASI2J6Y0Q
EgTiJrov59e2tC6loRqYIzji0ooXanqf8F4z2OwA9IA44anatJN+tTwXW0Slk3sC
IrudrwYVT0EXSYRMyoDXHjS41tDbhK+t8MCrxGY3sXZRxnQJwbbuJOI7AJGhkZcq
bFiOTC2y8Q6Oy9zxLIA6kRT8YeJ+55aH0bcipqbzs6q+kXJOZkMffzs9XZeemUCz
cz8lQps16AoRPMoMg6J0wvE2Zp8GKGuTOhTcDsEmSX1N3egRF2H8ZLl8BXgF4Fmp
GF95Zc2cj/g1B4xLhzZAo4zSp3VISfxJatBNrtJQtWoaLNZQlXdYhR6RMXCFtuOu
vlANYC/bNd+cEdIuj7qndG4gtvTBiNdg/8FceAP4S9b49K6/P2DdTBZNT2av/HvE
m2/wDstGJk2m5WcbxcJZBhdhjwan91bofPTUDwQOklvLMfLDTk1LryFfBb6K4nac
VGrqeQhPgpm5S91pSzdgl3FfH/I8b76Q1JIO51ejw4Oz2SJMM9ZvP5TZsz3rIoKS
/AHDJKnGFIcoGxF+PByEu6cTyxdGhTHyUk3L9PhpzfHRqQq/ZkwFVtR6hzldK9we
xLPthT8ukAnWLhoQ0yMyWYEsZkxSnQi9H+x6knIMML52oNBXFX79Le5zZH2A5qPW
NPKZJKX0BEWd7CWgS5uc5tC7Qzp9RSfucmi77YRzY89Yfs/dBExYPIFtTfD1NMyM
mQmohAKyYhy0kaPAWr41ePcLS/LAgqvPN6aPiFoLy6wQOssXhJzLbKkW1X2HaGcL
CnEniQFEG+oU5HdzKuIrML3CJu3i/+cEgXo1Y1jCtayWAgu3ZSFtWwhJxhUU6j2I
Kj6+8HShXTEkNc/v3xG5OnTk1W/kb2jLgaB0ANsXqBm3XZKCFqz10UdnzdNHBQL7
sIgQSp1j7nC/+BcEAJso9Vd/cLgiDCotg6BFxtOCWBbxvB3gXG9rBX2uZ/wZQUUy
JNLH4W/hXWQMv++T/TKOqA4tOH45J3342GB6/A+vAYpsMBmbekvwjEONcdyfndEo
UwC49k63V3rDVFCR8PNs/MdC5CsN0cj7Xv2bvznhdF3N3J3Pn+ODB4DJfnZeHHeX
emVzAMxhmtgZrJO9+eSW7HU/Wb/P1ueOk1ZsyI7K1vTSjsPjcuDHhNNEx/pSAgw3
t8QWeOaA0wFRAMHtm2npEIJuJ8OWDESk0f5xRusCsgMmtltYA4bc3e16I83av8UT
JXLTsKCo3uF7anr+G0VuxxOZQjiPcKXdiyYJhid0XDCTY/zLUEG2Z3Bo0LAP1Lhi
i6eeW/fMIn78Iudcww/F3qxKZKhnz9KzBJcGkHbS6stFEOwIswr2iUN6DdbiB1OW
McbEAfnb2MA/S4JRFzPOrdDuEWkpTwmiuumQ2JIc5VLxHIE9tbTEpDCPmwcWNAxs
grHlpu8sF2vm8V4/yjoLh1b+Uk5VjHvH14P3kR7rBpd1Q4GUo16XnqeLNS9I/7sI
EjEC4Eomcxrnv2NxjjYRmlfhCrmbGiFnwMr5Kg5476kqPD6VGS8fupUcgppV3J2q
01L1ERjjBeAQryovqWGLoBKuansedqKKSZdeabVac02MWnJomz+pKig8efDg4nBw
YWQPq67JPv9D+Z64zYEM9N39nkTtBV5F/7rrcPEmql0G8/lNEJwHqr9xQuyhusHU
CEJovlPhAIhJWPrVcTQXmvwM+vt6EPXEnLT8ABUbN16JMdLGw9hGOJb5PpoCwEjq
BSS+ko5cVygX/LENQk19IvBDnN8hj6HqX88oNDwhhGh3+DUNH7X9lPbLT2Oh21BT
1ea+tqGwZQYqP5grUcqxlMWLsp9rS7r1G8puZmmudAT1NTLHJrJm9VIiQQu//xYF
g3FEAJcavtceDkKypGwcHDimsw/LQNK7Qd2pKxD2YtLpo1m+KOqsdE2w0ccYmMhs
CgERGiTEWifd/dDrtd31PLATtYiXHA7A80sm7eezLgtpyZRGDM1tw8horM8m2b1l
bjcfTx0SALesUtcXMezsa/3S6GQZ/lZBU8/Gl9L0/wW3PrrOmTu5A4V7RbqmUDxU
+/me3nmREaCFpaCED0BI19z36M+JuLshKS6I6JwLdFz33wU7CR027MFFcEbMv6wR
KVOM2NIpKjCeRX5BDSFdVwgQmm6n4kDosDyRII6PygHcUWCkKfeiNerVrZYXJUuK
`pragma protect end_protected
