// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:02:08 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
dnT2htiGwpYxsa7VNsmSRKNTqEjgKuKRdqUkcDe0sKyZWYTDTKc/QcRUNUuaXgFJ
WOBorQAcfrIvW7LQ3npKuP3Hth3bpamXCr410EymqCWUFsy+9RKfE2X1x8BaVMMW
UR0QnMa0lcT3MX0X533uNi+y3VrcN0fWg02Q7X1yM0g=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5600)
LJlNS3D9rJx+ovbIVlsSpeHqqHmZ2UDvTgGi5rUSYxyRI3Yf2A8Yv8sYjx1LCaHz
1E8FwTTHucAwPeqLXTeRFKyICTXo7XT1SDTP5hGZyn6d3gP32LJyFXWzzkxYtvmu
MbXJRJSggpgzIkpTGDWcNd2JwDT84WjOCF7aV9cSA05TUvuppcBvNJMTbTdhpLxT
ZRiS2p9pGyyhz+bk/CWPH1csPhu2T2ftEhgUIUsKj4GVJFHIVwHOFToCEqb2hbR4
BwqxDSGJbqrfgXSjnBbLjTNZAZl+KLvLKUh6d5MgZdZrifAAbWfzWuSErLrAB0D1
t/cXOVX1sQh3qTf629Syre/OTaIr/bO1eQcN9Dje/8yEaWm7X2rMt9GCNTDFDihw
fX1Tas2P586jrKiKfd2ueP+n5L84tLN5uJth9kvglhNkvjrWDbe/EVBO4o29GgDg
NijFvHTr+oWyUHzfBQ6mTloTbyd802xF4IAwlZ5A+khlXyJHM6G4/TLo20YKXGU2
mfN/7WEIj5t6GFMuZxkdxV9VGiEsCE2aHdslrHFEPAIsAH/G7kslo4DAkxLKMgXU
Q39n/YKd3sjzr1IydJifO8YWPftLLVR+I7FBoVgqgr+vZ7R58pUOEDperOHMAT70
Kgfr+la786N+6YTUxUyS7a15rF+Rk9WvNZ9fan3xDGlW6sEJRSKwaPoxRf6LtKbj
qisSpmpn4gZPrrmbgRpU53eeREd6u7QnUeN/jBzdA8IiyS3O34v/oaZTVr/ocAB+
+Hb543xakW+jqSuYTrSlH+wXGJGVifKYQwhvy8bdJ/MhnmHtoNFKaenT4YY9SwcG
DN2Ei3N82liadVdPMgYIcfugozR2APjXjfHL5KE+SZjACTn2H7j8mSRjzajhcAU8
5H4kNY0cR1tv0tY5ABaVMXilb7CjVANLAB6VoS56B+IMP+cGJeuDMbRjZr8tVLvo
ypE7d98Dyq8ugvrBGsIesDPKy6f65dYLtSqYLTqP4uhX1A9O27T2xZDbwdB3TPeu
txbIldxev3N5wQOG+F29DdUR3Wgpym7qq7ZjlQYSeuAe5CjyMl6Twt+bIpwuqCz7
u+zJwnWAxAWIdcsKCCHmbmwlCx7qb+TisnySm3YClNiYEV5Qre45275ItbXyc/uj
6ImuySNh3RB+H2jquwi6QHc/diGj1dVmvxcSb3l5kLyCA69tGKSPty6oSdME3Mzp
Ce083UKlG47YEsAo5bii43pJ93hL1OeH9EQvdW+4wSCRrwPnFuk7BHOpuld7W6IO
TL0CWSQKiUI9C6N197G0m8vAt6S+e3JId3z0r2883X11xKnAWCKp46LZnSZ0PfPM
yI4GSOlwU+yTZSp8if9yB5SkrqSGJ4GviACfvpSG5aQIcDpnX2SZCwRh4L0gg4X/
YXghPkPY0u+3LzKcu2u8vVynuEXc2MHt3XByFLd0tQ7N3CmnMDSsbKHuXi0YctcC
G/PcOSJcu4hu1ERDk/Sy9v7nR8Z9CKBM00hNpTpt6rCPZa3BXTtAVtGtVp3x+EX1
uaM7NcpF5cE5s/ok59zkSpt15y8682u6b7wCivmb4m6scZbkBlZay0ZEkLHrKHes
rwsZkcLFeqEBAV2XMXbF0KL/f4aUfZAvh2HBJgLAThopVaViPk1+L1soitu0WtKG
NvV9ksR9DEvP7a5MsGUCFBM9ueMtyq82PNZSXu5xw5C7h0mJxfdCcjcqKK5oTiZ2
cL+mqK/m9J+z+Z0xhX9w1fR2VSf0MqHsIkQeoM3wpAKkJNXUna0fkRt3krh/w6Xg
UkI+yuHdFgWXymwgVKe1E/j98fHVUgAeJ0PIvE1bRYZyfYhFIlA3eWE2mTlUrP0m
1wPypBshX+A4R23PhbcJaDszBaT5SE8FepT9lm24nMABYQZcqimnFhRVEHukZkc1
WF70LY2gHFMYrmr89Ne0mMX/L04dxV0T3yrlqIo65yLcMsK+GxNtMp70qy+zgRNZ
9hfWCjkQG6X1Ypq/cd8sRXMvhzkZvdR2NKeM0T69K4MZR0gfsYBKIoZBRKvZ344o
qutsAiYQzjWXtEUs2ECIF9f0FcQcvLguML2qT84ol3+OfkAyPKl1KjbxAzzahb9o
YV5WNq2k7+P2Sc7VqAnmMuLrmFBfU5dtKJuSWsBgmsukD1hPCNIGk/VXxLKgOhp7
pW2jYqC/FF7S5mBeqDXLsntq7+UfmThrSfw4ZvfZf3aojMvcO98qsfjkBDWenz4L
otnG0qFbn00+nwVAlGFCvZPKFaL5FebNV+Gm2Uf1mfrCbZnDh7q/Dr4Y9IzdOIgh
aFfX9Sz/Vy8seoeMMk7VyKkNQI8/qsZJSK+jERq74ietBTnydFN5axoXGQlkjLjB
JVW/m67wsCatHpKoCj9oQvno2qMQ32mBzEDdSGohG0Qc2wHG70ixBkZ1MnGsMpmv
u/uBlGozBUoZwFN5R6koAWCsmlyameYAIDMFgCOwLzPxmOtrGbi+BHBJ3Hx1ZijQ
03c5Mb+uMYQhp8/WPRJj5G8z7vAK3EEC5wADnwOaM1VcPjQ8TCa4WfWBujvPsWsp
8hn2DkYu34Ahmg9/opO3Ej/XdtUCwyZxAWTIP+IVU1eQRU6+uyWgVOozDZHcifZT
rFX+S5nEM5LqYZpIF9fns0cQapJhBS4Jd/7H6yJ+57bJyueS7mHj+lHNSkn7WNmH
JDkp+s+Hz/Hk1vgVwEn53zuEkjZECawgrXWSCN3YTXz5XlTEQ+xP5zArOTm9ihj5
RRTkmgsi+P+NK4STr/+p5XJqAXt5/VhWbVsGG6U7z6N7OB0ffIXTrD3cX+BmN/Lg
hzy2WvZr6hfQIC9Fm9xBdJmC6DudvehSTMR2Gtk7g6oVEGkpYWbJkmKI4IBc3xBn
mkreekTTUbKw2vWKq/AdWEDQAatFK2F2DEdGQRWBlkq/8CFzsEtC8MwUFtzzsr1l
DNVOhy8zimFbti5eULKKkr77KOkGrUDzHBQw2F/jAtgpO3saps9y1wlc6/zoQr+q
tp+LfeSYEvBcPCPzD6dlAlfIMn0+eK1cNUGJ+2OtlhJDWDYZHp4BPizlVQM3PE5+
rC3CPArpPHqMhiQpw9i650UIr5w6WEz9SHGhbWVpv21V4PqGgjGVvE1h25UOLIE4
6Sg3YfEe/KEDzJT2I65nbR0oVULBhcpt+51de8IKtGzW32HIrXsCB0mlr8WoNZQH
vzSBJjXn93QEb7AADyBHcW/yLfW66BnglI56URpOmHKD7VDqoU5BoIU8D+gPHqkY
JPOJkcFr8gEo3Ya23qX7WEbqPCo9EzHM0m9kiQw8Y4UpI2CYdK6HFpx+UcjMw2cK
XbAWd1ZQwnS6xKq/46I1tZMxCDnBptGqZsfUibysKEPciNCdmnI+QWq/oSyVvB8I
c/+FhBh/8n8LuwdFyT0JG5sgfTVhMVv1aA+oTuW1jWHZ89Q9ktKBwuNuCkW1dAjy
GC/raPJJgCgVt6DmmG4fKVmk651qry2M+aK+gi5SmwicC+nFPe6l5T19eiGvY5li
oayb7xKXSfxH/O3KpVdSSxBRduQvq3wLbWwFOE+erjCs4ogbccpxbBKKiPkvNZB4
gyoNFrWOpm1Xp2rAA6dZlXD2oeOq2NQAU8kYu6aLGiVKG+nroEvM2H/9MqEJI+50
NaH6dCOCuPMoKZiJ8ysdF9T2xCuNsL7afeZlCodiYPeFE5+uBhcMhaeq70TpMCAk
hO45R+uoEhW+9hy09XWlXRnvhliv/hHovnMjRnMo0M1wO5NT9ZpO/YptbGkzT1Xf
nBtHliwN0jEQxZY/fII5VVEGyaF+EWhL/CN+w6uMykhlsKdNyj8LCilS4GdFzICH
2ZpLbjYWFN2bK33HH656sIdrpqkXpXQAqMpHH7+jYf12KX6mESw3IpWGXWyKzAIA
qEqiteBNyUOZjZb5H7gW+7gdJTOaVvJQn6GAE/4QJmjyeS7JpGdKOtDRtcVhvcXN
KZmY+OKtAyK2ETvQ1AeNrteD3ye6Un5p6xbtBzZ5+KKnn/jjJpJFFAiCQ4agtAGp
RWi/tMPwXB02GYCssAGq31JMC+Hd7plt3MpsjDJoW292qHMF9fpw/USmAGL+5SvE
96xwki9Nsg4NKRyFt2MXT+HQiFNGyYjToHY6eM++7+Sn6vv/csU7RsfZFNHz+mRV
ffvXW/ukz8cqwvhPYiZnBAqU+p6JP7B75OgO5+hbK2x0uaAKWJvZexw3J6yB10GC
QZtyA9PYoxcyZgSWRoc5O26zqaX9xWhIIEyrTKr9abA85pefpFPZMsptqFpAG0mx
YiL4sWV8WgSQBQPWY4pikf23nhYdUKfuFKApWgGPmZ78iHCOYhM510WdEWgj1Oo4
4jqis8BtKjQgZc8efgMjYLF153u/UmxBH53RWVf4PgH4d4lxAdALlADuACglVFyu
x5iMhKm3w40a/XPORH1lKpwh2wPkwKheGs/KWCk7nIsZyve42ZVQ2SB/N6foxztm
5PWRGu/HYQKXL7AagxOYl+wLljsPewJ4MzTU5D67vIuk4VE5sGBBIEaLz1z6o9Xq
V19Pd5HBdapswagk6HuFfWtpuwZLf24PfhFe+PLantjg30LB2W43t2ILXTJ3LPLf
1TsfFbrpD0Lb8a+hUNg2AXUqo9f/jazHJQrGlVqyJq3jGgGeSmzwr9PgtSn+YZTw
ai9OEh8Hm6OCHoshaYxa3Xpc/25p4eJq8CxNHXl4iqIAQ+BX4rBIwXetP7JoreRM
fz3JH8GEZdtiQ7oAB5gBINaSvjdbv9GEP7DMOHejPzVQaQ4uQs1gmTE6FzqVaL3O
pmkAethZ25gsrq+hcgyAw7XlT3uG0UKyZkBMl92NcmP+lmPv0tX38sgO5mlagiXl
Ctxes0R0Av3Gpx2VFnd1+z1vcRSM5hm3rlZFe6JT+ZqFakPKWux/uu80IlJhxCMz
Nn30JjQDBY8l1X68FE5KkLKt0kuV7h2RiSm6W++zEccoHqqwWNTsUryTBh/i/Gm/
fByn4SvD6yjmChEcNbQenc36nP9LYwfW4OQ9ek1JITp9Be8hqiDBhtWoFckyldbZ
lLQuINqbBxjuT4xwqyltkSwrn2Gps/kXN05HxF90cdD2JgCVqjfmMIICyD7Spqkb
dCDwhjNAHTXD4NB1HQSSyzHoLSq3VxuNcf6eQeSRUoaGbGqJ+UbBRwopcDp8SblU
s7z5adVPrBjViAxq2Jb5Fm2Q3FvUqzJr/G+9j7gh+nJ+2Rx+EVUJGZ8b3MpSz9LV
1JpcEXfgEx1Wp1OQXP0yHtRzp/V5vI9NHTh7ARHrBFrTTtD7rFpmrUBKG+BOnkPf
PZmMBvrbr0ZdM+X553h+EYNC9mXKERlCoP1CaYXymB3747CE+1JVzsE+Zp0DaD94
u/GaN13z8y3Im+xQtsGbWjvH3GL6KO5TQ2b7XCASH8bctBG02QMB7xGwyLxhx64u
RWHRUho5UJJwhzci+/IjbtB6ir/qwfbrrtGVtECJ9+Ddi1V+fAHI+Dn7rXA342qG
VmqCfs83UCH1hb9qiDqq220L8p9iqxPs1Il+C7DOQtrVB6m/KSe8JqXtuMzPHPHM
EvVlcTIbywuFXLRseTrcWBXOoFRboX3QS6aFmVEsZaq0+Diw5CcXAdXBo64GrbVh
dFltjokcg4LExYYDS0uJXNUtkqxvaR2T6B1WhLaTULAqMBAhKl1XLD+DGJD4c31k
LbkvfwYxtrdJWBqwljSNDR4r9vPbw4fa6zkjnROUeeRD11TK/RJN31U/7KuSu/SK
hO5Qr5ApFpur72xwb9vdshKgV1+izGFgi/STVHreaLKqFHLisdmSXFRjRA0QNzxQ
OFCu0jt91ViL6W2UHgSRJjAkUhWPHFKJW1QyKdiPAzm2Wx9Hu6Gc4S+lHQrLMzLY
1rbPF4PQUwntcdrG1RqwPy2dzDvvncWS+hjQmMncAki99gHVxLCFyfyIvRS94Ldw
WvA2ufmU2eY4ZhE170tVOFzHkCLUa4AcWmCm2rDYWFEEelYEGKkzvXqb8oXYCKtR
3bawsJYLRTquM5IFBXV7/R65HBdgApXqX8AhSpiVsSq3FjH9AZPPVgwo+KXrLtTi
/RctQQ9JTZxgrJrCmqQWaogL2ifyuXyqbfwF8ttzHAbe6A3oZlA3n8V5TyF6cCg+
h8Au3pMA8cklW9c8ksrUZF0XVw8Z8m8VIhvf3ri4vWII4FKCHUZJaUeSTeh9GVzS
4Yujkt5a87/wPDKiRTdJMdbGbnFQ4pJhvlSFnU8jSoh6DKJqVaZNlbAmRJmYDOzD
QDyw2RIeIVxISamzpvwKub9BpvmuhKQ7P77FFYdDLJf3sNk+IaSGuYpZGBTOHb3Z
2wDB/tV388nICw0TyA808aUevxLOqGSYYL5Rw635gzQTO1kSNF1pFkJGl5ZLJ73K
2cFUEf9fkQz1lH0P5siZSh7yDVMRD7sZgpdqlntfoXYkWYanIC9/9aDwsQdF0WNP
thl7jdVzvquTY/eyUMWVqhFwx5WEr8EuX6d1X4S43+WJ9+gxTYZsCIrA6JY5FUo6
t6wPySHKKBG+yG0/XbtntDoUkTIAnGGd6ceohs4Oimc8w9+ebBav139YXbaX51oc
4eAOjU3HvlW8gGeWa2EDWaIKN6Jp/hDUr6I6bY5RS63mK3wqqb7zoJ7OE6QlL727
TAis1sV1+8pWpmkQ3LquulIt3XyzC3RS6IoAoN5MyQaUwyX+TQVGT9G1s+J0BcWr
JR48CW/jsbS87Uc0auurSRw6PYsZbAJ/H7P1m6WMTd2QrJqCUnPhC8pnWmbWW/Ej
dGHTY04okQGjd9meXvu4DN4VbQ7d15rmZaCXm1kUhLhbv0Lc9YqNYZXeOnuwkCT1
km0jYv5nO2oIKrRQ3T07oj9pLbxMcjUer4FuujNT1LNmKc1S6LtRLHcTUAZAr3oZ
kzbiqpMm+n/HSaxV+PfOmhMuzdDNd9El2qd0JZBRl75uD+A9BPycKSZjOMWy7xA1
IvFSxdJvDR1On8MdIV5+vEWBasjiZP6rWlOgCT4GuVOi1YOnfpddo2DuWnqQOdco
Hl3cQZ1jDAdG7+AQOPPWIRRLwY39hR+phNZZssXHabjP4GG4RYIKdQfroXWwzzoF
A4xYkilyStm3+ZQZSSm8H9tdb6sKJMPrdW3GikG305lXO+/6T/zANx/Wvr3iy/Sr
pdtq6iu/fuGE/Pv3o7l3nzHRF7svzwyo0vhO9R8xVVhcMpml4IwwXhaqiTytYYpw
v8tvfqYO2mbRxkORTHVR6fFPnGJ5Ki0t6SgAvkeZU8kuZtX17aqtScPBk7UFnKb/
DGJUaZItKxfIq6C+TRPd8ND2g74GM+WeUq9HZ/0SfCxs1zybYDs8dJVTXll6YnBD
L35KNXHbLKVGrYg3NeQthKCRNyUE4LNz3bBYbo/yg+biEDQ0FDNQaldUI5DNxBqq
oBcIhxAlqHJiA2fOEFhX2SDBB9UgWLnQsb0lgcc8OpM=
`pragma protect end_protected
