// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 14:01:38 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
N8QUD6m2rQ/wYxLRCyh6r8AIYWwTRu7Og0xXEy3jul3nMhh9E7zApfdiT/+F7UGw
z0K4S4WKZKqsfNauFE2f3MrwN6sscjZhAHmoxuh0vgv2iPxxR0JxLdqwrbqmVQvH
JdrMDmfvxGxyy36n75cCred2tjBUlC0Gz5nq7hCIZZA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 20992)
wmQVP9KrlmjImtX0TNXNU7YLEGKdcJwcpf9/pQr0ubHrhw9EFTRHr3kak8dMn5Cf
PTMeiVdVSy9Rb0H9qNuWtgrlMTwI6+vY8OoeRhb8tJoajNxI/9GlKMyrNiz2WzWD
fORtKOLtJQf1sIK+H04f9p5pwe5ZelvW3Dx3IMqb6tS0C9Uwd4hpO6EK7+z6Nhlo
Gs9Q0rr26JxI2s2op68BiktU1KKY/2oKUCnjcvy+6qj2VYqGw9+rEwWYyNiEdQqR
Rte83awg/54B1P8h9FsGoLBT0TILonp1sLOlI8Db58TOVEhI3buCj/OMgRs9NpPM
0znlhUXrxzzl5qyLJVj9VkBDyuVcIx22eDSqcW4sHvEZGMfiDM/3PMcHxexw0enQ
W3fRSIBYXmn7y2jGMefLgUeDShjyfUWA/QsW+sHMXvtZpqPf0W8ziOSbCNj+FJ/B
YLv7rzubFASFxIQ9tusI6YRh6+xGl0n8mgaz4RYM+cm1Lt1aKBEHftBqXvkuVADX
y2MZoFBCD/kVZJBbIihQIvAnuwLQGuOgCh3Ji620d3BwLP2hCsEjjH2cjTMsI6fZ
hz/j2L2N7be7PsDW6pYgJJHhllY+4SnqLRszt/l+zDVmUXyJeypum5x32cRxnHmN
pTNHqILGwhaEIvhYx4O9X3gAGd42TLPHi0pir1KaAzDXGyHrrpw9U0I2V3G5S9Jk
QWxggck1bZ5IC0PhT8ij1iEVhxrd0qqWMDiSQYjiEQ7E1/SJsr+BAH8nOWzhLAcG
a9fNZeHtfY+MEwrd7Tsv4zhKOEsTIU+AcwfVnZqcXtBEg+3WxjAvv8GNBLELP5R1
/5JgpsnGJxRKTpwl3XZELqtNHNK2yFaY6dQBcMOlcfnXSiU/bV05DlCNakHyfqjV
LaUj47jeT3kf3k3VR8wOd6fxwyQqkiFDCB27iyNoxMPzYcGqXuSHtF8vl2VGfJ9h
LWPqHoLUqtr6a7/oIirW5FW06bU7AXTZDgou7OgOYdRsi2JG0YmPPYAjYYBOUril
iVNqNQH0R1ZtMlvxfRd9wWTVW6H2rCxycP/IF99+mwHUvEW6AjBMgHsuWAbU58TV
xl7EwEdzHNK6dPQenwe51oX32vxFURDP1YJm06UrHztfmEFlsNz4Uqwj1axctVsp
YKi5/AQtqvU03LWwMBV2U/QUgqDUEKP2yiB5XiDdW93Vx+vjEq+DSB1B4ELe5q+v
XezjIjI97pFIQG3J+/YnUCtvuAH6g0rfICaE8c/uq+KlVmGqTM7ITRWORyU6KPHH
aUTs6bfxIXm/f59XJekjQGIOIVRa6sB1qayQKiL8VPhzPQRUiYuPgYMJRUYvX9Xf
UrpsFgtaoE72UIhQWAsgTjqJZtZq3Ktgr85kyYIDVh3eAuk3ULp2A5bgknuJvR2W
5VWEID4KdV0Uvf3eXv6s8Iap3JTHM0PrnX0v/RK5UoKvlH/383QIDO+zG31bgAxo
JlUdy92E9DnVKLIujW+BgxRKO+GNhiSRuYF8oLX3UyGeomMXeL4Kwfmfj2plUfkm
h06KIFxvV1lydvGVveVV6tl/Jk+S1bogZIySxHvo59mop+TzgfvFrdEQiZbm+Ql1
Sjkv88rJv/nx2aBxpC1a/v1RBnlzG9I41BSbjklB+IBltRtLCTV1mvhDb1yyqPl3
HWUVK1EFEkYtyzFhr9dNiHPCqkwaMbw+M9T4iWQdEGiVnvFUAF9THjYJJoLGHSMl
Ux9zag2f8wP0EAQNFMwJ11/ztNmG2OOJaWpWFVlBjW6vNr+b5guXCvSOGvup5GeE
AmL9jkqIfGRRGuQ50uf/UqlUFWUExSpoU49redhtTk6aLblpUp4Rdt1sTmKCk0r2
ObT7cFPiuglY6NyRoq7p1o67xCQ535eUsmW9jrq5RWcypryOBax26TL+hg/5xAWd
I2B8gdPVW7g+QBUkfJwXNKg5v8Sj+ZtAnfOlrvQ91ZYy5AdmQL99fJTcDZmgnCYx
6QNCYy9RWX+4sR4XRdU22z++XLxDNiJRCQ2BUou5jkH+k+/XnugeraN2eRaju2OB
ahgsccoEdlFThlvDCVKU1hwFByYDc1KP12ez1P8TVilUUrQRKOKh5mkGQ13ea9Q2
uvTGrjU7g9/EAK2vdPJKS3opBjSn+ixFom5TnldTESWSFeApTtlnp8XXqjZT5mht
Cjc77tKsjP+jcxC6weE25eF2p9dYXDKmR7V8x+dUepluabN1NAsimBuhN6C7Uk6S
jpP/0UaT/9vo3i0rincptyTjjRT6sdeRcPr9CfIJJBqfEFb3mGPYS7FSYuO1WJ45
RW5I0ejdGO111vvP9ouLAliUgg8tMF7csbp1unQTMhe+++JfFVgm0ips25ke/84k
VID1FL3ZYraWXc0p8TnPE3JgBIlL0F5LTgtqFiFoj3UfCt1TqsIdkAJP2MWirJXU
DAhYsE7Ga4InxiikfYxdTkQNEMYUx/wYNOn9qlUC1Ij3Yih1N+pWOaza2B7CCrX9
5bRTylHtwIOIMIXG2RjQKoldfj2DcbRJZzg46rgneYhjfrlEE5nDB13ng0yhqHYS
UeXEaIgqfdhfjtVhoGwRXomzUmxIIXJSOtxbl1d24lHwEJqlu20jHlMvZG4u34YE
5eUnNvSgwVfu7l+tURhIQSHkQKn9yk1E5BepzFsQgCjGHG6a1FSMedxb8tu5g1gD
TvcJ08yDiOs+SOopQ/R6JYZvYf5cERRddrCZFzcjS+X+IwDi8GSD5vMwLBQcfRwT
yimbEphAV5QJ79LfMzgtuUb9o/cD1N81ILpxUn1acAVUAuv6ZbsLbFT/o5UwGvCB
Su0D7eh7Zg0l8E+dVJSTN/9B2loPMnZ5V971yZ05hPb/POTG+tOpk4AM3qjFtczw
getskM7CWSD/akwOs5d0LYuG00Uw0hCuyIsp8NwWwh8nXuKot88MX/yRPQOWwPov
5TMDJ6fkCetjZZXOZqIkC0t63KSFeGgiGDLLtrWAaOKJkXNjPh60NeFAmck9euJs
O7VoN1y2m0Pom9/p6F4m0+thTIfY05quUi3KEdfL2z6KYvbt9wtD2S3lW0asJTZ4
14w9W/xl1wBazdF0ALTijOeSSJm65pI939fVbvyh1pW0RMygBpo3m5ZK+tt8+Us6
j5FEAcCu/nEA4i4TchXG5NES/fPYZEjN7sJIp+o9AqOhzNWFLpu/pxg9ePaeIB7A
fBsnU/mAlyYcLudNeN8aErTL8cpuMJRQCgQB1dYj8tpo+/qA0Dsc5cROKCyqD7IM
Np9AhvMV7VyR481PY2QAHLId0gnX/Tkq3Fxfl3lwax2w5+TfkaKvSeSX8R/wFO/M
cVw3o6kHYdzSnWP1KR5wW+qNlhbbkoXsq4zhxsUwUkZrq0ximLkBv2Q+X9cc+UhO
AyPlJcjKJHkkAnV05EZRR/kbJewMYHg0gV+n7MHMwglQUXGjGJlpfFf5JWPO7v03
U8edj27nBoJeK1HhkpYIivBM+3mR6xV50WOXZNkmgjGEC5Kqj37gyAJSZNNLxw4N
WsIC81FPBLXag9o6hb/5qImH3SyFtE1WOQ9JhFfcsRJPgxRix4LPXBx63jPBKQny
cJFds+F3rdv3LSSROABdT+o0tmseA5wJ6ueywe3hsFqmdRxxDpQqYI9q+fcUjtfR
inMVv4wSwh5WMtFdUb3IpNb5QkwRp/lVVhnqQQ78CqD2tXfu3sdWO/t8Eln0mQc0
wK1qs6lDAExSPbC95vhqK4FSUHiccpHyfQ33Hq0XAdw/n9L9zkxmz+dLDYP327dM
lWVwcKy1KYuzyDm+nVTs7zqVuqeD+V0NDxaCyCC21mMsAG4GFu6ao9chQ7ubTbIl
zwxpQ2G6fPcS8pTbmza4hXTBi03wG6Jj+fBjm3xGPOnqlKPm6ZQ7svLfceZf9xqe
aMiqsOjggKFeN+lhv9JqBmTI6gYmfos7U6Ua6vb09cePn3r+g21u1Rw0XyCAJZ+j
WaWySg2Ua6x4l9b8DAxKbCHayOUWpFyqcD4bqc4Q6Kr3sBaHju1eLrEII3VE59sf
RAqe9fIXjGuf0jzq85e6TxNDLpJTNX31x5WwdHMMzMTUwrR+bwAvYd2NP5g1EepE
pzzJzRd7jiTHo/hU7LOs85a4On7HeRG/4NG5byo3dAvVKzg/+UA+zAt9uef6q8/t
o/y0sakMvXzx8Gx4uDJEvVAWxYILxwbrh7jj7+n3ZLMprxrt5GLBmSG8Js3hHIaa
o4AiJmTXWGr8/vm95HwDd+RxwxAeCqF4uMyGh9rSnZd0j0Vb1PWT6RZe80xU7AZ9
8mcEeR0gZ3/jU0kasQG34ZnMp+UzXSN11td3EXRQ9N2UQeMiCO9WWj0HY6hpG8QF
9fv3PtzwFnceKlxCgTtxC55E0jIBFq5dUKX8VrkQD7n2vcylDmh89vjbD75ba6zt
1tbwPbYQapH6oOgiY8h1i7GXyuZAWxmY4CtFFs8DefjHTcQBDlH2BdOc9Qxzu1kd
1UJ+bt2o8GW8TdjMqvA8axNC2KPW7G/FMOP6+Apl9jFGthHqQiOxpqOmmx1oB9F8
5nTKFZibtDiIfAPPmy1hJtvoE3DWr9w/93PKz9dNvinTiiKQg7Jjw70xU3CqM/HZ
SbEhOMDNmT9iEWzU69UJzEVgabRIKTlnayyitjDxgocpIm4lC+9JkH5bHjnYzAnU
N6OyC0KtsF5C0f+6Vt0p0WNYs2BQ8hDC1+bC1GqDhIWqSfFtIASj0kIf4HcSEXRf
yY40ON5g9a0OJmkpCYk95IKwgWdXgKM9RvuzHP3lXDo17s73nC3YrcrPK7TPZzUj
oJqm2mLcW4qK/HO9IrFgWC6slPAbkD7Z75V7Q9lVGyZxHTKjip9CVuGZ9MoCJ9Ld
4RxpXE7uVs5PvSmO2mLQvYZYWTO4Y6hoTc7ZaYaa89u4vn1UB5IwFmzpNbXvdISc
d2EkGQawbmn0BewTNAauWphNhm6lpqEBmLir655rnMv3r/dPG4IdoObF4/yDiYhC
SsgLnT4DeRtN4DIAmhhAaDprmstDhf8gtkZB5WyVellpBgJOmUnxJhNm2jLyuwbl
5z7f9YbMtL3ZsMqwanuFNZWUfzd1csqtFm6ezmd6GN/ZTu+5cxy0l/UFYW+49Xi9
U+IsabL2bM3CWLtKQDVVZq2huJzzUmMwqx06wNLnrGlTLch7BXUHfHjcd9YLWKVl
liaAaymakhusdHWT3isTujqMm2vbFB698+fnjgf+2PTWkCD21JS5VI85xQYN1tyX
NRnbWDKCzftCaHuhp4i3cFJ3FRfVx5kYSq4wl3GGXBgdudedqhIm50UujC9yDPZC
x3Ig3pQWch93owXkeT637dBxQweef/o/zVxkD0vpShD1dT3TGGqXzA6/j66E6KL7
6I440N6uKm3yvbQjgVvJzMeM33WJMBj7L52nJ0lvrmXbrQKAeN+EUVOsfGFxDurX
MqEeyRts+z0osUqdn109nU+L0DTJUGNzfreuvHLopMtv9cSUfACF74uMAJ+ztOjw
gi+fTqk3fDnYoUfuc4DKlgD2t9ZE3bjz64cs9aYQ3mx1gAVenCv1pptTdu13lVqz
ednKCayp/KxUFtiNZZke9PbMEOS3/UvOaz7nw8KM5zDwXqfibWY1xagZOZiWrMoh
BwsWcF8XogsxKqH1i4Ab1io/K3wFeJYfOVjP0wnsGQFpdbBYVXx4lNZBxFC036UZ
FpLviEoQti5N2eUGBO6U7RrBrnp8LAovmCzz02kqQcQ9TH5ci0bJNmEOLM+x9TIt
7gL35G5sA0EXhyOWzW9MXKIrxQhFUm6P94YNEGtvshXwrDbanqB6WqrRMIRf/j5Q
qmDYe0Jw11oiJnryzxiX40kG/YyJwCbMxoor54CPVpSktHctDPXgiC65rTb0gE07
OFCaJwsVM4H9rZb+1ZopEGRuxTAi0VUH2dooBIuvqd9ve37HLCwbt77kLcZLcpyh
B2/p10D50ee66JUlLebPNsV9iA/9pSuPW4qIAG1Wa64ropUW8vp4NoBMkEQJaibx
xYQ9wncnOuFw3TwCrz0ZWJQrBCmJdTKQP/yxy2qC03MmLZpEj+/xKzDXUmvd4XUU
hjudO+uAlaj5OxpsayG8o6GTwKSv0c/Q+0uixs3lE7LmOJWpha2M6YQm9KoroZbY
QQlM9vOqamu8b7858HC14J8Vi6UlJqg3mhIqCypoaP5ycY+Et/eD/tWCRnutxMFn
s6Hswqt3pzJCH1LyjB6RxM8ySGbrtLhXHJ5Urb02NOxi4IJAMFZs2DvKRyxn/NY3
/SHrEBlG2lgtPMjaT7mpEgqw0XgugqWnnuI4m7xr1Hr7y2Byr6iQfnBX3ws3SViX
cOCrVKhpqJ8QFB+FuymrlGuoEmV9SrF+N79Vwrfobaq6E2RodzKp+RWQVfMd0a8v
bRW/us5kTEu3spTrr8zh3LaSkgx50GvlMYgedkGFisTQTJsSevl+D1OAqmI/6y19
Gt2PXpzksoWEVhTuajZMo+QaW5UMtLZdrMhmMto5wOdgllharRX9cUgeKLGfvHS0
unYHjsefVrHwv+RmwAVtQcxSzIqwO0iyXjpoC7itF8qoR260wNZR3+febrUYmpY6
MZl9PSLIzdbR9pZ/NeI/xsVTHp+j+kCFF75ZMHxdtnwHlfQiAU+oYNAJ4yietMKI
qqXnJNueIdkuoBqD5fBRQrRCAbXoFBvBxjekEXJIjjz5G+ahDm397sJvnSfyQ8x9
F3DT3gaLGaGJGwwUxf1LmiDJGwFcseV92D8NsOkxkkY3ef9xcwzg0M01icq1bZ7X
NU5cu5BhBwvXkblxhlW+QPnNmov21AlA331ZPN0imVIGqjrZA33LKPWoZOG6A6iM
wN+3Kv/xjUhcPi+aNYCRzEFfO3/JQtMZYW2pAdGNBcktuBQQd9jlPjP+jkHnJW2v
LjPeSBEo7pO3vIzcPI1szPZCLwlG0yMu/XzHXTKYCY0TDfczf5FIFXV9EWnnwx8Q
K7c+6InTd6UuBXSJOrkAy6LIG8mGezrbLkVdBeGUnFvoc5JPLMRtLJrnBidlZSBG
xksp14ppw3jYMmG0bQg/R9e07uya5qWyo4SLD2L5TfypRJ15XF2bmLBSyeFhfB9b
UmIQZr+sMH1/240D9YTTLSROHmC62ccwF/Rmtmp8zVawE3zeNzlJGZDxPG8xXt0C
Rd0YUmhNwQdnnsajC31Ld1kYAvNeZas9Phqk/xYd/cxqhK1arwuB4wvBzCQLKnq/
qcHbtT1KV0+RJ3Ni6VuMbEIh0vs9ZZHh2lzFdvTlv2EXbKU7KUtL2oW+6huRfsKk
7jw3y/ykv9bST16QH4Is/PTz4sOSFDrAVJE7ziBTwLGGqgSAf9b0ql88kCZZ9HJQ
fxMIIy4zQJasvXsmexFZYzYe573vB79zyAZd6m3oExNZGHm5zUnMqZGAuvOvJ7pg
R3kNYgxLggiB2wc2o0+n1wLAh2pV/yglmRZTCA6oefAOj/5OZR0wMSowvzNqmUVV
DJPjdBH3XjUPM+W/Bkhw4ziZu0WEpLnIQFmY6p5gXQdKU3q2ZTwRCX8sJ+i0uegk
K7Ly4Au3xYoGFZwH81mpGhvAbXegOjBhCJ0DAl52Mr7DEPiLbOB30LCpPk8EDe2B
pD3QaNcMRlS1iPzvayWFHrAcbm2E4rKd/G2CA5IEX1+naLmQYJ+Q0r/fPs8ORMII
bxed2h8wwk7dCOXfW5sOWfnBAGL1h31iUIR6c0UOZfDj1PbYDKmZCusm32yA5ZRc
zsfKL8wzDHSzxo7k1Bw+WhElHehOiuQADhIoJ4zAnXFKtE8K35tyxipUwv+zia8a
PDq1TNuXC27Jd9dNk1SnjafJAQKHtK3o72ezx4/sz6J/zV86NikfEGnUVbwSDqBp
E7j8Be5Hx2YmW5jW2sy6736zdZUFMbfYL1scvg/gxxyk7IgZCpYlUTQ9bZTUrSBX
L9MXfKjHjLCsTYIL8f8HNrVRwWRaKZ50Jf19mgrAI/iEx7uTIiDsK7tobJUEwelv
D8zxmi+FZPEfq1uSPnUuoE43JfkK+EDr+xuZ7/kSEzio4DD3RQCRzrrkqqOvBeUh
cSxzDAaplCuYd7HrGlLTpKdsHPzBR3TyRURyQ4MYUIzrSBTe7OWdv5lG9Qh8oJrw
sP/SM9mYGVKlcsXCMtVLw6Nokc+fRzvEHNzCiCmoPSRYIYP6jWd8aUIU8UQlUc9G
FU7bbJaPytLlAl7W9msNmphcRIsiX+FNl8fsOzCX/rTWMLc3cVWVGHPNM0k2Bead
0aD8qnGmDU9TEFVaROUsRzW4oI/rrGyXVxKupdOKHz0EK2H21Bavwm5OrRODEDkv
NGcLsiY2q4jRniTpylRy60JMJJjaxOXtDqiPR4zPgD0C5eUxSP8CJMcE1yrtaQkl
FnqfW2RMbcpI9cRwNz0Nw8IVbHBEPxY0224E/tjsztm09535kOAqt2ak8WmjOz4W
KtmGjzXqtlykjM4JyQebHYRl2iL1j8NfbK9Nt8lNuWX4iy/ImvEblpZf4EeewEhy
lUsdBAiv0xr456nUrISOeRKiZDHD8Axf62dEBHOHQOec/1BHRYehcro3cOqKM87I
I7vZGZBwIell4j9jTXbK7B6ufA1Q7HwUnU1uJrsBUveWCyj9oGmol/NNzxshY5op
cduQU3EpsxCtCQF8OJLimjLrNarG+fKzwNVjVHxApxO2H4TG/6otunnV3A6g+5fJ
yG0y881NhUIvxYiuHffQG5EdXhDSiiZk35pSajS2fU865r0RMzVLjIlBzmZKrHZb
O3KHT1qK7qHMOYuN5zi3g8fwKMOKbOeXopygYb2Z9HXst7PGFyl+DhuzguqslMrK
Qkd8VrrY3lUj4v1qjajoOQSqZT3uyjScqmGZPD0z2QtIToG331mt24536le5WYDZ
wjWiu5mGN4EyUIlRyQtY4YDRmDCexqQuq4R4ElR85Kht1tppEgU3st93Bc5SW83M
tyTRYXO4sGurOHkE/X2LKqlIYPqAZwaJogg09BKjfbhAeQjSxmnI2E3LOVdtytzd
T0cGwz0o99wn4o3RsGQlEi6soqv8+HlQi9aFxZs4K37GMLEAk3H2blcBKXfVH1UY
HMbPvwFldjvzNdzTxV9Mq9C/TPKhoPnQJ4lT0xVbkM7tc6gTCgSPgHFzNEg4wZSF
OXMyayn54NByKUJ+CAtkHghz9ArFS74V2aloyWOciWIGXYX1eK4tal0ll9TL9TSH
cAW4kO/xihfSyS2hWrakJJVhtZ4lu6Fd7XIxwnBB8lk1lq1wIaQv853I7XQ7KMi2
+obaISbp9a6MUeiMjWtWsmZqd+aLe4D2/+WIUYyTvW5lIlxCNJtsX2+rI/vGJaW6
YbZrUmMd2ktHye4zxpqFaJao5qtwuRGvxGWXyW+1T+JAXs8v1rugfccx5s753wa1
wyUBzGlJEXiKIQoRO4O/UQEbbsrDKAcO/z6Klb2CzM5bsWUikPspTK2PJbTn02wQ
iU9QcI7VEO9ttwpkBlAdWIeWvtVToVbqm82gJ2dUFXDiy2HRFiM46WuyNGSCq5Tq
BrhExkfd8bclOHUxszWKuI/fNgF19EbWke64DGRf7ellWKgrFaeps/vZaSw6+6Si
81xBqQZoO4zRStwCD5up9NKbKTMhDQ5WTLRlAFDVWc28aV0itSp+Cizkatmwfi3j
S6lUQXov43Vzu00fD9LyQDETlvyHaMb2N9VJ6nEI1X1Mj73YwIwKpHi52qK9I6ZT
6h1+EIfq9iRhe2QtbNdfIAHibekGVJ2ygddglyBcsp/MTs0iriXoyX+xNcIZH8iF
T6Rh06/nJJJHhhb9NfwR1uKoChaIcFkx5rS2n25MhY/FbZZvg1Ynxuf+NmxsSSVg
lw2EwfExhuIhwOR5zLTO8rFmewMTIPwbQU1CjaewiP2dJn/mefsig5ddS5m/LXlL
Nnnx2x8gWtxEgw7M5/jbJMi378+KHGKWqqtL/ZqGbB/hf0RgJl2uEXOvnFjK8FJo
GOVZOBMrbpVk8R4FgPHrzf/JFKSsbH4A7mdiDtFPnGDuWk1YBQuemzTBcvRfapc2
KTdqK9dRV3pcl9H2Lff4qXXs16G2dTJ3izEA40dyDBq7oBsdlmHb9867rPS36RJH
jj4bLjJPjmEr8xYRjZFVYOxirpnsk9QVcsqTBmA+qmvKL+9DGQ2jOvs78Snrv11L
aTtliwvd9WS3wcpAbLJw7noQI6ASvGg/zSTM+YTsrcp1Iv/vfWMgo8USajB4G/j0
uGkQKj+IvD2nuk8zuwvN0yhVNN89Zxe9emqnVgLX21oLx7bqPNC+ekn9YrK/Hx9r
mKal9mLd31PMIc8803KcvFnGb/uMWfSc7TtjPUIe9rymgpyDnDwUd3s6N+9Uetxb
wUClJxY0yueaAHz8tgFMaN/VnEuRcaZ4MqcmxYgz1zI1nNZTwyvryamZV5jE90BP
1cvF6Fi26U/CEGs6+l4wZBew+tGzIjao7nFIKOlf0FhtmaC9vSSvq2VJmxVQHQuE
NmqafudxKHG4lLEJsBWRE26hTwX4duOkRtqfCeCpZ85gHRhIneYwCdoq7OQMP9Xg
oUG9TQClIwmn6hpr+zg90eyZin0iCvcKnTlCMq4Taj/438vy4tLBoVsEaDtob8pU
ocx3SoL1zhGZszXE9k1SEti01pyWqKODulYPpEJaW7o27Uo93lWed4Qz33jz0l2C
nyqAGTxnyTdGdovS8dAl8xCYYPs+EAEePiG6qTtTcey5h/Mbo+nklvKr0EQpJ9IO
NZodVUo31F5RmKyGNzXxSD56pz4ch4EB5wDlsuj7YECgaLuarS7aUAeJb70utCrI
xE4yKhTQRf34X4CWSHrriQyHg8gwznoX0wE4OoL+Cj0BEPvc6XovNHMARWwHRALB
0g+OndyTUGaYWTJLKfKFONlo2WDb0Jdu1FDNnoJf064D+pr+FoS+kN14W/QcKr5W
H2Boq5JPDD93IgLUcSnRvEGw3q4jfqaXfuukjF6XnvqvSwLAb9+sLLDcmxjtunK5
9eshDqs8Sa7waQN1obvt4OXgryfyhuSPaAKmmZ7o0SsW3npZvuw6ajQ2cEqbV5Vd
41XWV29e/FxTlsvJMrSptiMjvjDfnxJtOcwRflObsmkTHQ1aeM4VrIP8YbUVQ1eY
mKHuOCVGQrTn/xSCO66x5gw/hcs7Jlxc6TrPcVlMW92VxbYC+fwvONyu3krhkYlh
CfGoMrT02ukDQ3HBnqOgQHK1taTmsRJmhgObtdfs9osADvLagwPsXuQGCdV4PngF
KUlZK0ojYb9XWWKnc5Uw8WAddt8JyZuv+N1iRqUGQba4XXy2tPR+MPE87g/y9GuY
2VT7sdjE71nk4grBXzk7dtTz+QNfJHfTX2RcDutQPvj5Y3Ad6hgIzZRrIB7VoSbJ
wY8beKJZ3TNCY+OVfhfmApDa50i7qMVXlgxfbmpCN9tSvCZnIkhTZlwyCCUTvqQU
U8oFwY6ib4KGC8e06av4Y9/7sx1bGUZ1wUWjH4Ezsd4KOnyw7uGUN6uvt/UV14yt
JEvRaupv46Q/1OYAZHE0xYbvDi5xJwGFs3pxbPzBCIdOkXqwURL6NkOW5zUbZ3Nb
pkCIEwQp2+UfjC/2YqMSc+15/khTPNmI2iz3kNkLsdIndzVKYJCd5Y4Hi8JQ8buN
Zb2e/qC0OBZejycC9JVISOaYyHu2ILvdlAD+ZL/Mdb07s28oeJtH0tWtugCGErTt
x3dXKIcH/BnTBm/aY6qx5d5mOKiwACmw4Llqtz8zTA9ZX80xdN+hjCupqxj8Bzp8
aNsGPG2Oev3VvAgt7XYZt7WjRqxjyff0L6dn2epm8xcWIDoV16xapyTLYNDMCFhN
Uf8c1XJQOTw914T8fXJosxIzcKWYNAA2aJrJUR6OpHpVYfADzYdwiG5s5v7qW6XR
+jjL61x9zhxJG13vPK3ebKOzLYVEfYJhKCsrYBKtOFg9FUP1dRnA6lP7u3sRs6zG
vSvd2k7Wstt8w2LA1ALVTb7XjccdR0t+SbtGJn7y/a+Mj0trqlTm43wjiGoxL/rr
6N/KdynuiPvxeEiEg8URcK29pJasBoBgGhsLsu7fi1HfuHQwL0QlNTutbRi++tEI
+HRWSIgpC4BUK/TNl3GjRaggNvYE8K51BuF0cikX0UQ44VyBvqzE2cweVvoVC0Ql
THecvjGWokZLPheNsiAx13oflV76LZosq1WFm2bcc2FpQj4AyakoBMP6g7PZu+Xy
N7jZ9NbaR8NMEFhxNLCc398sn80dVgDNBu4f9eArKEGZUYewg8PswKdvn25bsrRk
xfwaNUkVnkEjCl9TLF8ev4Ouam774E4vddtAFA8ieXKiKmtUXQ9TGVd7rQZlCtYx
miy6zR8i1m2kbp71HaLi1iOCubgihjrx4BWjhZhENj9FH21D2gJ9DXpzrGTlPQ7Y
MtGXHE2OofDMKFqSorpb69Ou8Y0zEmZyQOSeEceg1gF3vbKHd2uSgzo9yy9Pu55L
tMA2qxynG31lgbny21JL1Im//tAzsOIUhuYXMRuMtzLR1gGldQ70UlaBIfAg29Qn
8LmX25K6tm4d7JBP69c9ss4xR9c1BwyRvV9Z6YwwqA2q+UPWUsvtyuolLn4w3slC
6dE7rASp7ohjke43eVlW9+W8B/hWJ4Wc+du/4tVioQBSXMEbbunONpViMu5pI7rW
WfqzE3zWEiccP2/RcnR+Oda3qkImrHr9RyCLcJtd+rneqfkqWpBxTg2V4WnGsygL
rSUrK5hVnBXvviVAWjCEzDGrWvQhVIZ0TbyMQDDGn6wPd+ELSeRAeAiRKEBtf5N7
UGbtiTQ7lRdJawwneNryePutDlQ03EmIAWQ8AYUHMHEXymP58Y2pDq96D3xefOvu
MQE9C+k9guDhJbBRITQUGbdTWcvmiZu74nJgcd7LuI0350LohwipJS/Cv0CooNPv
QfboO6kEQXrmyLkPdr2C300LonsnH6NeBq6NorKrTqhrGs1I1hMDoIrQfO6+vt5i
FCfgVVPeMqJhTm/pk1V2wPUCwQoG/T5Q2xasthPpUfPABMDZdqSRuEm7w1eKcS0L
3iZv0F+NZ3GStLAZzsGh08+twBZGRg0U7I6ArxLHss7Z5Mqx8Jmvj5YefejgEDDd
5tcwdnnZ36ZPSdSLJRaD3DUHqBiIur8nBRf/viS376+L7lV/mThMRUmy/qljOHOP
4KF4Y1fsyCq2F7bfYQnFkqaGOwK6L+bheUGGMcqZaligZS9/K2Pkj8UzamSMHO24
Onx+RiKzZAwhHcO3zs0VXSdF8BDb0+pzuuEZZfEP8ljkWaMxItRSwkUpVF5MYNi+
lMzG9XXnzPDinPCXLUHkhGkNoqykDSXX0Vc35QYVqDbzkWmh2h0Xzey4YEUNAguO
2yb1pKsOjRrUXJkOG2RH+hao9vMS6gHm+1DcTwqHeMpiTf7DiCEEBa+saTcBVI0+
0FK/JpBX6tk8tOt/Z9ArZ2TQa64FZlrlxAAvJDMf8eZoCikQiV6unZr4PGUlgO87
Nqoi2cfJIOhKK3+mMvInAODcJrO6WIepQ9GjemvJ/lxzW6Sv1/CmJeOvPktN4UzY
cO3y8tI9rkA5rW/3hoe+UlLmuzO8Xe5YxJeK+ek9P78U5S7VECNjI38WowkMLphO
T4zpBXMIhpClqTxt46eGwFlKaWMQi+slKBWDcx3NWrSsnENfY0e+wpHCI7BNYRn0
yqN0rvuzi69IhdFjnr/ZkmFoE9SLod9NsbECJdW8aPN4LZkMYcnRrDfYyKeKRVLg
5+ktoaBYN+AEmHJmQqdA0gI4hOzAG98F/SOF2/ZFjmlVyeTEhCjT6VpvBMntds1O
x+60Unl3XDfo+u+wApvlSmmAKwNsWlQT38MmBrZhD2kWucuDo23BiLVgf6dxuoKZ
8bKv8vF2qx39LHFLJn3hE+/LUy2DdhW7xwtFpZmoNbL57xwYz6KRFwSeN0DaaKXU
oL0prvu0DM/RLBaBHljJ6lR3yi80zaVX+A+YPyhO5vEyzSb7a9rfr+uX6MGdZiDd
qBYs3N0ukdwyfs8AZSOn2LOw/pQ75ifV4GKTG1wZv2UdXyPEjMQpFTwAPeRfw9sL
ARDqCOkg1ld16yHQV+FYE9RHVXY2yFWYuOIj6ws2TKiDLPaKgXPJhspauegRGuHD
KDlEL/37d8xNZbweMHSQcexV5qO6ZbTjEQIoJFpRYPCAr7XgoYDohfIiFK8YUUuZ
ZuGuJBjbDcdpyPx3kWib5Up8JrlQdLrMrYLyY1dGpmCQmb9xpPcgqsXcVQS8dRRQ
CQXP3hGsOWzsbinfXYUBFad7ktnb+yCBDvsEf84NqSLFKziN+75Z1rjN+vXrDvmh
/cjNgYOBhkNZRW4fAhFamrmHkyWcdNm0DKzCYAXR+KedYP7KovLbUFk28wL2q3AV
TWf+Sl4/j4KC1zQUn85Eg8Xfme7Joi/6DZmmZjAWkLO4onKday2IqhmyjlP3njCo
sJXUwQLNdxiaIBiBitK5rVkvr6LPHeGVybvI/+/Hqj87hMVaK9uRWPjqvgdom781
jKSedYvjFQaVnpupIfaOiAyr1AF1gUbz52Mw4wIka1mp7Ec8D/8PyBkj43PjmwrR
WWFFOEutuAZY19kLH4eiTttz8zJYE55atefAWECm0bvy/TDHdLvvZUwzODv8ucc3
qXsnH2Rgs6IpPaXRbOdK6cYvUgMBEeI9YYZdSCdVrQ2FKUJS1msJgkk+1HiQQeF3
t+Hjr+aoVsHLmtAcbfz1Gtdw2YzbO7dgVOoyW8vF8YHuNHtOEmlBdXeURtWsoUMK
ztGto2G77SqmsyRzWIIP/qKxLY/HPe0n5wYTdG83HGV7tY0eFvnqjf5xsbhXCpjy
5S88KUePDatdKLJY2Me1vOIK5SFsZNpcdnEaaMwAeSL6VZnKgMXWxHPDCWUviR0D
pNO6EZxRxXCr8TdLhdf54IZWwxxAZuW1Cu2zO7b3Vp7EMv353hVocZz4q1tI8ZNe
1E6YiuFx77Je48k+EFuDES7dWppBTs8Hztn6B86x/wxKMpyk8AhuHyukb2mcX7/4
ebQJnSB/2LNmADmNHyCOG2FKublPYvdThlRx0fDEWuKn4oJO6aYPfGErZk10eo8C
2iI7eogHcI+HU0KJsJYOgezyTq1TBPR6ZYyD4TIhaPuAJeC3GBves5IvK2zmuzcF
Mcu5ZTjN6K44qerKIyCPsb2kHrAuee9nHFbKN9n7KDAbsVLtBQB6DvRYNPyyWS82
DddAaH8TLU4LuYkZQlh1122L9aNX2UVVdXtx3SguamoTjuWehOGMtBqgrmWuCm6o
xjmbQwchP5Q2Qom9OgAvJQughSC5MBJAOYSdIqasydfUDakMPEtkBO39AnCDCtjN
64J1vc4E+fSHTvEVS0rwBGicFy9TYPLYuZppjU79EqfH+zmh/WoS3E7hg/obWV81
vkOjUF7J0gV27pL1vTCYIKnPSM2ANSItl47S91i4LFY/bjbq+m510v1ePcnLheyO
ch9nabfFJicPM4NwjsGUG/POYVhsmqAQc+yV9M6F5QP9z0OG7Eex0d9aRtQPahsM
tAjuoKG8LWWF6jdL00lh9gQhNKKB9noACh7AQxVGU2ZOTBcPd8qV86J/GS1CuVoc
Vrti0G8juUjtwj6rL+ZGpIolZ0PIEcYUec3PYxLbHtKQE+IgSEIWuao0+IbDJtp0
+3opRafMqFmAK0wQT6wk9j9JcjMB3jjuK0vAHO9vqT92ctza5yjEdasFC4o7IyAU
r172ziypAQK+fE1UvVBbKmkPRf2hvtmZk6FNiuE4fjd+zz4jMI6t79cFG6y5HhR2
lNxt+U1cFzw+5bzUa+1jlRmzpooalDEQHChSXsxs8NQuz434bGfj3WZ7D6UooUlq
NLwKDnzBeHVmhl8dz/SHSuxtYsAwCJazBiU5aRXT+EH8ir5sQ+pYEqZL9ikEIkAI
ltwsEwlRB8COkzA+I9780iymR6l9SAAuPv3G6fND02p1/oyoxV4NsOB+l2SbKgFi
ZGOt7QdRSZjkTur51GNVW4O4z3e/3PLZxTSZkvjQAto0w3KGDE6EpKr7k37LKpI2
SA93sHPQXHOQGsLCMR1B4oExNWqSuxzrXRCujiiCaAGx4GHmK2oJ/eJsxVgjR0Jo
qjgayoJkKs4u9J7Xeloo18336x1Mumpt8Daj7z7ZYIgioFhILh/yFDXncV087qCp
haUxEv7ILoDje+Pav4ejzyfP72zlfrtV+3130PYNdHDZZ0bMyGSgDYNwBPWzBaIb
ETK4LTOkR/BshqwGNO+1JJvW8Ldsb0/rnCWJrMyL4qb4CY77NgBn7UmMQh6t1c1a
k3tF0YC491khHALQjD4zeYXMnja/IMEljePvp9Hgbo6wEgMtZsMxK3k7ZMVPqS1w
sNMWsTa9E5FiCnPwe4Hm1Lp0nZDnOUaEsLjPbmDbkT8SyOwxC+Zs1d/2D3Efn9Fq
ME0Nl1MLXGxR9kPCdoWcl0AfAoVjsfiIWRCBSxoUgLhrDCqx0NhAeHaTq2rta8VZ
yj25tSe2LLICEY683vSJ/M+y/0hUzvZgrBFO6zz3uFj65J2c3aWYEa6/WBRoNZ18
u18uW1LdOJ+H2OMoFc+nkR7C0t6tfBliHcS3whCbl4R1RXyZpdtdQcxo6L54xDlN
KjT3VXA41QQWPv2/ov5aFylXiytDw6h9kgBmZCtGfsA3e7hgHhcWjwlTGY2bR9nL
sNLC4UmjDFJXW/DuA61MxKx0xI3Ks+CPhEz2nkMjwZJz50aiE3qqB9MY1tN+r666
Hku+G1lUOdZWOeGNe2B0FUjG+381UkKig7rW/fyOHTL02w8vHBuLYXcS/otBtM5T
yTBsV3GkSOa/S43DiyuyY2FbJGO+EqJIc3OTURxAA7ZGDEEutFZCqnt244ZO1yvE
SJUp+8CdlsEPvcX1AoObUT1ELWbpcHDGSilIkqMuZ/b3TWPU8QDXCR7kAeZb0aA4
Pf7wuXU/y8JQTad2h5iWez1BU21OaaXmoYURL787f0uim2jf8RknskkSD1c6D9IE
PUCYxZ2aLu1D/6tcHo5S3cRTl0XLf5R4f/fa13ALYh0/ZUEQb6JaJz3gzVR/9Be0
y6czzwGyZOARchE5Y3lmwbejhsTFwERYY0Kx8S8pi5bGXvaiNcZ7+SbJ6s933+wt
Olvh7z21dmeb0rcwol+tmzjNVGmIQqHQlVSIXYZBAkWU6aJCooVS89kKp0ZwZqV/
cYYd5XUlABImqCWzaQysLs6haUMdYmu6agQmLmlmQIoS9u9PpxJ0mPno8vlCRNEJ
HuVlL+mFVT4RcJilF7mzhYTEKoH1AhD89tryhyJ6agN0xwyT73gj/MCaq6IdleNM
s2VzNibmQM8LK5LtKE6j8Yu9SkxZiEmar1mL1lS2/fuftRO2Fmx9hG5oycKf+cCW
mSUItwRfrCU8nKk0VQjYTKKVX/yk+MuQPH4ruHir/St1DSsOnwMPqtcXHZDk7SPF
dPFa/d+SPQdmFriQm82ysNETYxGkvnFn9bb/Vt/MY4Rf3gA9rpMhugGTU1xujIBP
xWNyTIQKIzRM39KukHooSropXaG886frzpziFx10uU8UDtJxKyUUK8sTjsIMmdOV
m35KK2VYUFGJc2AHom7jeE8ibCyOc3HemrP8WfE9tEhe0HJlU+C/FNy0y4gX7n/h
PAfcG/8i6OhDPVES0H4ifnkulkBYraLBAraeVfNbtKVage4O8uzZnXWtFegHxvKq
BcBUFZyLdKeo6xJxp+F5k83pEcIbXUdwYFjhhqCnjM96TudojHgBa3NHg0UL1VZ3
IEZcIKEv424JPD/WNAammPO3FNYLy83pJG2m+DpToa2RQ7+BkKzRIlt0eMmyMeI9
LBzAAwDIQrJ9nIGbasBVZLjxgNrP3kmENNiejRrVc5lyY6ObQNiZuEI8kxvkD+CP
330VRT2mYeaSfioqymNauDIMjwOqvgc+8DQdktBymMYMUEfkHYYSTdBJjBPD2CeI
6XHcuf48Rx3u1z5s1bEQHs9vehh2h4d9ao8YWv7XZpask1R0Pb+mvZEbrDB75/kW
jnS2mvniYGbcXJ5FX36QJwBAcidZsf+3E3YeZ60kJDFKY2IBu1Ly04FjQJt2yzVc
Y90cvt7Kj5k2M7BhnSz8xJ+67zC14wEOlNYI9qN8u26xgFRD8IYAKNbGQfwQfteL
95KmAtvm0TwZRdMhaSRAzPT0W8FEV75xGN6XhXkTUuh6m20Ci6cB+AGhK1EzzUYN
1OzeTNclcvlKaArIpbLHSU8RhK1lRb0t7JP4pSbwH8liHWpto8u1ppc65n2rtpdy
2hdK4OA3XdMvIhXtckPSN1yG/mcHfb41XmvW9Wu1+1Jw6WUS0gBrrH7DHTXxjNbU
Ao9E1E8+JvgcujC+WGkne82ywjBwZ/w9DFsAQNmJWNDAbX4MBIk9i5al3SBMS0iU
1fgBdELreBJiWeN63cE4Uz95uELSz3TjBRyz1XQktS/lx8xjgzEl5hSruBUo+14o
Rt2JQeNxkSehoqGQSX4LWJiRpJ6r0b1f3ZpJ06SAEYc4Eyw6/LNGd83fJL9rIJO4
3H4cbW/lDfFJjuRbyZYXZahGO/Ax+3Oqmse9UakcOLWSCtQ6ClHp48emqPN6P3qZ
IZdd/VGYIKN5+oLq4sBPPZfkALJKLE/OehNA5gJuk9MBn++8u0Bjb/v2Fds7aFF2
3znJQncnrqy5XSgMSndNtXcWLL/vKCYriXGVPa1sQUkTF5ijbGdFJn4J9Ljloi9f
424wwE3qZWq1sPcNRsUOYvaG+rTiBlRC5v9wFYWberaymECFkhXx8B2sttZlGaoY
78x2xrEyIMywHam5BkVd4S0/QOUahpqf0D1Nf2rGZ/Z/Di9Hse03KCJnxGi4vrL+
zWe1ZZlcOItrRYmarprTsYPwjUwYm9BjU8NHgkPoIkfxpjPw84GbcBM7Q+lq4ZHt
8GfNLzc/UKZaLvuwFkQaDjBr3gJDgK95RXzvbwapHSmJJf8oo/9mwnl8ovhw1Lx9
5VlAfX1fH9s7w7Qz3nQE9aa1xGBpwdkVdVkRdQlvAWhfZv3USU1bEfABC3h7xX/5
OLdSMpDOTAcrh4eeF51USPAFdgClbPDsmkTHxXkGAHwbIAelHukPeH8rdNfLAoV/
oyDJwuwURx3Acy5dN93Bf/H+tYQQt38csh8dkQmzDPM2M00M60duu8UOwKXE/K6E
VoKodXGn6bF1ZD+5hxPqinRX0yzyK2iuJ9MrmNcQ00KfgtXPxgRs4KVvntkmdkkD
8ZvUQ9OqASNaV4VgBN9TVj+RRmXNzS3IPyQnn2B1A+8qpH3CwM1xTl2adRNpfgV/
ofJhgmbiGFUCqVfKdHLHLiVdGDBvsoujyH/a3o8pU9aO9EtTMcJ0mfXCGth/+4Gk
hO2ilyGdxvnh4kqdHhxuFtLK6XBRW7ESpUJGF3aRevg1x4PfFgIi+BH7cQ9HVhWZ
jeemd1dzdPbQql473Cxp9/Nh0wNmhTma2+wzUoKFLno643bQvbXuhgaTL89RZz8b
DgyBt7rquxdbYnVijx79xZ7JsjawD6sOpFgF0fZh0Lslvlne71LJ5/mNYzXvcoKs
h6ux6DYFr9BUGPvNOMflGbbMegkhLDhueQjwVdjkX0u3Cdohn1aNgY2Cc39zysM4
WDR91/o2DTppujI2NBopLG99Prs21Wlr1Z9V3tKke0P6X8aVV21RCoLnf9qgcdoE
d2pZoUubyQxjJyWYNu00G/f/TEnEJ2DuKRoorWO5xjMM27u78I2DnCB0MbZY6ErN
M93Gn6hNHmhfUGsVzEF/UWJFLOYfCpxWQnDNtxRmcw77+HSBUamVMERxzddxWv5J
xTV0jUg92iBYYCJ3Q7jIysuRDvT3LyQLKpSBKwTL/a4INzCQRcDd/doTrT+hFwv4
H/oAOdSyQc1M84iOQrMb7PYbjZH5cffVRXe2khQ+0InaIvemvBV08ftB+nb6Wt7a
IBniBV2fJVuhQVUZbcvGezP5GIiQzY5dGRhVWYq5IFEalGE0ahTZ355Tjt4QHso5
EHcgDODkgA5X/Z391Hp8JV0hrU0m3oZ9hrgQG3F2WsriSke9P20hFyQKGxlh2wd5
pNu26pVyYb+HqhEDB/R+xscOgPFC4q0EV2tdiXAW7HgQWUl06fUfW6eX/YP12f1K
zOA1TXqhDdpmhlSD4hVr0hM5n6Q7nHsDvomsm+ERVeskajuMrG8mWL3E/ts3xqJk
k3Cq8qGElmFzj1XDsBh55+sTD0DOPuxzSot8Xzu/v67MI1q3hYoEfLmvQt1aPV8r
OvYc6fYm0DP1RHo49EQCAKac1qnDEWlD0mgwV83yBRvOR8jP3RRuKxuj4ic5KubN
vVRyKQGUAepKdgXdrTy4qZCwp7q3SFecRFbNEA/C3RbbW+NpbLr0Sx3g2D8TmV/N
ydebXzqxtSUCiYyp19SoDYEdi1NfXuVQVNW+ZNWE8tepKgmGvKO0H0qWHqCAqL2B
5F5KK667Qy+WWOxtFgS4b0IOjSG6SJRRAnhJ8NCiM85kyR0F66VJJIkRcE8xUnrc
hfMVDCJLOFOurCtuase89pbpAFxQZkjeGKL61wvw6y1mE3kFopzP0ALMLB9VRz+j
pdUohx6WZvEWZiNvOyphaWGRMtjWS5T1t8+Uzbf7VWX2BK/oAl95k6RX5nOh/I7g
L0Wc4XYeyFDOuAwIep2pp1QUWNkD8uH+pNWhNfqfB8UJ0ULNqyhucwIX/jIMXEvq
NUPzbfP+YrM8X7p5urD0b2Co6OaWYPjTb8Xp8jv0Z6mKHKPx8m0UAZ4cvMOzG+yP
at1a0K/9MBzJGfeBZQMeIpKvaiRa+OUGZbtq1mkFOWlEa5dWDkV/OPZOmJwccnzX
yzNf5lwO19V55n38IFOvtejThrAJD7cwatwlgRFpP4dtaomfHwf9yuWTCBkhHpUj
nbnGEU1LRHjohk2ppXq9NxuT0sMbRmM5EFKBspQlRsljrQ76wXNVK0enUrP2vw6y
CgkEemi3zz5KY105H7aUcYXA834QdaokJ5gSEHXdDeve9b2H0l4CwvHYF8VTSaa4
X0gp9ZfoqyUIYDLcZOf6FGuMplxH6gKPEGXfGOSACwN1qYoSXnciDpGRib4QU6hh
ZzLyn3sD7a+EfQZp4c3zU4cY09xJsln4ooHQVI28Dq0ANVNQh5iq8QjVqO9Yo7E5
A/kIqLZtvoa8oc7XpcpiK2biZ81xfkX0tz92MBGaGaLHZbjtwQdK8mPJB6nyDlpx
T5cwAseYMvV8WOVoMcPSySqKsoqDkPfzbYGor7oaLC9kiJbUjOYf3v78uuQYSABy
Y3jaqnBaxAt6ApaLqSgIh0VwSo12Opy6FfWfeZ2SgYj7sLw+JIWpaj3hJY9xtnYz
aI4yAyiBYqc4+Sf4MJ+P5Pw9kS13qsTm6WR4d+zSdEh3AfnpKk9aI/4LFzNRhfZd
lOVsuhI2qB1sslMmGYlmgcsen3AegJ2yhcUNchOvZpMRV0UUpz+XnRUyMGQw9osL
m10TyuEksjqApgQZgg/k3frraPF+92QL2VF5M3fUPvI9nWkeNhG3iUyeIpFIvtPz
/+BuV8SSI9OtCFVPmjW0m4TDwhxMNOQU+Sg7QXU4tNOqlOn1pTSbjoTheo3xtTnF
Zhb7qN3bGJcEi1WakvAA4vtrlOcZEovoz+3VtXWqssNycbZC5x58E+aKIfHJUEoZ
BmcqfbVxxLwJS7CVQpoBG8Iwx7gkJINvcc/Lvf4L6mRw0o/H9pbQODbSvfuzGD2a
kYqX3vupiblC27pkv4tClSOxgaIcJfqVILGHmznZVxwwjs6XzMmiEOTLzTalj29F
D5p5/b4l3tmCMqJjCtLjNWr2pUmv7bmOg241IWejv+l/rTiX2QyAW2mauqCJhyym
QBNIbn3m3oUTe/xu5UKGDJ9QsLDM3GWr/TKeJQPdIwv8EVIe01BAmw36vsl/IGqa
vQljJJcJiZ339OjHfwqnssT+52B8pFe32SPcIIgoxKSSctgt0tq0UHqaG9u/u5uU
2irgfrIbJ1KH/X0wJAz1ib5E+REjMOtP20jhs3AVFPyF4mwG+Z2M/BZsdv99EIiK
Fue3ac+HHWcj+F+/1hW2ZuQqRKIg2nUIoVpidvoPNTqg2UWwip54mMSID5UVoMRj
l6whh55/3cL8PHW9XvLcGAcqe6qCdf6F1echBDMqfL5RNUTIfObQJ686Qet8epKI
pNxxaBm29q8f1vFi1JN4vMdYCYdfiLWXqOWlgupK6Cxs5M9l2HY6WJqvQw7uhild
W7hsrarh8tkQKeMVGXtA1rXzJzgobE5Njp4pSEExp0rmk53UBvK/d4A3dEFoUCHF
YidX9el5RqKrzxwC/njx/e5oEHWmljf+f1J+GpSEqdaxUJOALRN/lwyZfAdevzVS
2D2tk692SAn+QCTToEdoEIkkF0QszWiJtqYP0znLUl/CE15nR2ydpcL53ujk/imN
8KDYxmh3nLam8g01c74+VIYZDFBo8xiBF7GuUdxTVZKx5KPhlSn447nn2aVl71Rs
SyJ3p7As1TlPJllAA4S1+6s9i4gK9enodZW5wHOre/3yiOtTjucY/FHVGNR2fdTo
Hnfl5tPZhXsf0qK3dOuQmqgckxP7SD6Qj4Hb54vxg8JkVh3oX1lcxgQuX8026pOc
lK8YvzzqjAidftCJD8rNnD9YF2JDH1SUZrYnVwLwlI3yxX8eRJPL32BaQMnRUfUt
weQ33v1Ao/By1s1EyFwLU1vFdXigHJLFy7yw0nZzFqIJKMJIqQvsN8x7mTTdFquA
YtW5oyohsysv0JS1Qx6ilIzC6r1BU91NX5M7NBVftn20146IVv3uDzswIPPBpj5B
3gDxgamwO52pMbKaycZZAw/8nRqTsK/kRFBY4+86c6KQ496XxBfOjwa8aEHYfnKZ
JWWtp15V0J1WQ2SeMrabdtghNfoVEJBcmG7NSravI0SLupzbOEvz+8UQ2zqAhun1
Ri2nIDTNO3tRBPvMJ23nm+wqmItDQsm5REoEuLfGXfsEKCc/68Jp8q3Lms/lGC+S
DkiwQE1O7jOehtGrzD/M1TReqo6zDSO7US7BfYhf1NoHijlF9QL2ZKSXAu1N7Ufj
AAYUyrp4nKzralOE3Yg08ZfL0NBYI4zNQFJH1VSPUiLygFUXa3gVJkwO1R24FqTW
kcTLqTmeZO/8kvV4xv8wROjwQvleogxv61S2mNy/ZFNwo/SIFJ9WKOhUFbaIZIe2
zaIRBr75QhI9Y3x5cfGUbsXFE8idwkSSrUnfdW2GOeEG/zQXLwXB0629iQ5XT0dI
el7Dxkw8M5yvY9eP3VCZWHlSSdQ6tke591J3p36v+QDgtnmEqw2ZB6ZqX/D9TRSt
2+BASc7YVBtwl3SJBa0rqcENW0wFBBMkQlJ1RT8//Ml5TgzGkDHd1yhWjFldst1g
/z02WPDaF96IQs33bomys9WXAhP+vntbfpG4s51y56+A89CkcIXmZNwPruw0x3al
9C/qFN8EQ7sPTLq8lmq01m5+uyPVw3QH/mqDLx2YeL0YQvOHGerjkE9zXod1CcQP
ggUZEZ+Mm2jBRbtqpzl69xzshFie0tSVr65IYlScxYyAKIpGhuI59BdQSTNRHgzP
8vrtwva7P/cxkISPBifg7n/EYADvEkuCAYv+SeHeLnitgDUGtAp92E0DiROwsz5e
I3atRdMAjKi4vXNtyXD8m/768PWkN4gXX1WmVMUjwyJfvb3hudtL2G6NRUlQkyyj
/JhlAonEQjQQZ9EmL1exmaFxxUkzzIfnSLHGpSICkFx2gfTrhuWNdEt//N7lnPD5
lKTaBHYizKRimfvJRTX2+qm9soAGNhahKZS85pLWt6BJxRMlbOXCcwF1gTgXyhOw
qb0vnYbqS1pTFA6tci6zZnwy9RTWg2sGLNwK6EKIORwjolPXV+m6Imk9/CMZGkgq
kE2M46PugInKFpeptPB+7kbk3NYV9tw1JRTGP/D7i6IaaIwfnyUFUAyWdJmSkHDv
APjAPQqp7rgcxbif88Vg8yQ70RQMoAL1SzQ28fLWe+OYoTJgaekOnk8GU/1mHJl1
na+fdAGYVq1ekWt+xtQvPifILi298v7JQYYiU5nSWOMGWONH0/H5pw+hZdVOlJRd
43wGppVBQ7fxwEKcX+JM1zGtk6tNHBCDQb+5JDw/MfUtwzagRMLB4GDkvttlwmPg
hSDdFtOimsXoSObJOSUn91FWZiuRHPPw/LjSaBpc1x2ENYQ8jbdnuHRKK3fCKYNg
KVqYPKHwYgZq4hPK8i0Stgv8SIJzoWvsl1ik5v/C5/gQ3GamBZ1rsaK1EgQB4BcB
yaSV73C2H10tJ2neExoofyYlpy2mIkBiZvHZ8DELE7XP6T9kC2sN10oeZbmp0oPA
wiWjUi1WwnouM3n9YrZZkFnoMyMcvv0LVi/vOTz1/D/URG5ulX9v1FfUKv/0TvPf
1uzoNc8UURxUogEgOIheqecKEkRr/r5n/v1d6qkI7ewLIy2ZFhlGbz8qNQtx2qaU
fXs/7qsYtGmdDeY+EMDxbse5bt9FYDaEzCSwFUwYMqjleUDljQz80++yG1zqiYE6
SKOUk4Wt/cjGPsP9nUdg2/WAlkIwjv4Bzk32V0aqlC2QB6C2BQKUNeHfXEEZDvKH
vot+nne1H6V88Tu8vhZFfKjGhFbTS1OMfw9y82CrMFmCoUfGdcEBA9V/Peg06sWm
BniB6iieCNHJyAi0RZnZTvgjN4jGNcUXuKQAiolWkBd223loWjuXtMC18ofp+rvp
huf6TyGWFtomU3Xt/fPgUkGof3sv6CCECVsJMOd6wuS7zASu41DrGRzGHVdx8T3P
VSvZXRKTl1yrrydbUYLnx2TH5O6ms44BNhwpYZY0OUiDH4aKc8s7iWcNXCBKaq+O
TPDigoyOWVsUmQAESyKbVv8A1TEac1eMGBBmlMXoq+Ft87PC6Ilhoii9rtitia89
pAzo6Xzew8aVg4B2B0NqmBhR6bhTnjtrHO2nbr6YVvwaKnRneTrspkqwVCvNs2MX
mtNf8qqMHGfySdPyxx6PO/H1zrYq2mCN7KB5iRg9oaO7Z2PmJIKHgKiPSqJzatcE
rkPyfL/U6qC+EwKe/JwnWCixM8tsSsj6xRa7zmQNKmIFcjx53Rc+9lIYH96bVZpC
wi7qZqaSEqJvhJFB9hOkw74VjkMaLu+VWPHW+pMZMTa310edd47UHaQ8aJWnZgGG
TrkjuHDebiciNwb+RBqA0teD/v22r9904VHYWkp+VLG3wuwsSbUP/pzh3O56KVh5
iPb42hu1EHvt4UWlVbGQA6Ru0kLaeB17IsA3aYwDBZlrD3Gin96MLMuP+UnW24ZI
QgfHB6eimpnVtaGdusIFBF6XkYx+irSWt1LaYRgld7t8Cncr81b6+VUoC6Zrxcj1
RtG3uvcN0kssK4fvXRSZbCxtP9lJ+kIQvFrKWT4ZoOPs4h6RM+bGOVdHOdzwF3FG
Lwe45zRuohlSxWJUv65d+rceIZgwp0JBXDsoD7cYr9+QxN4CekIlY9qi4cQFDEir
aOmEJa44jQI7lKjLiUI64YhZxnw448JIpLPD7HCu4BRV/0jR9rULuCaRQFYC4E2R
+G2z2xmuF0VReOtCJM0rPsQlGvFKU5M+r2QgBCb3rs/HHN104ApcTayo/7OAPmMg
ujvcwOrwTK2uyfe8rPa2kjkMtLoYmp+qRpwJewxi9gs0FURmIb5oQqqrWwkXOg8t
RnYAIQ5vACuX78+DXmyDMy+y1fPTojKjgSkrZSt4ay7RYtyTqVg9eI2o0i8o4ehz
FpCFlg6Aw3ti7MLJdzZ/jlpvvSZ5Ikq1Md9YRoqKfUnaKrEhe2s+UL6bJsti2Nbi
yykX/wbUfape/dQAHljHWZDtnRVbxoOdJ/68CiBNcWDUj0bFL0ne2daexf5DyoSs
1YEVIWkhh2diWWEeL2/a+d837Sgv+772wradL0Rs1c4DxOhDuudmLIdqkquWdCOW
f8s6iQgcCjcIV6rCP50Sc3WJvTRCJ/H9tOrkg48fWi9zbuwMyVG/vtV/MPGNY9fI
4+QbEc/+RBc9M6nevX5vyKlpIaFzXdzRC3JQSh7GO4jdM0LIE2kJ6TW8QIuM4rhd
9V16o8pTldy4oIQKYS7kJBD41F3jpDCbnQhFCqMsq6dyTyLZ1s8SiLu2wZqSwU4U
Wc6/HCfWtZ19GFLp0VjVBwAlkbQP97QqhUlFH2tS4lOQorkdM1y2tstSxU/vK0UD
keo5GkXpq735jzJZG4nJsXONqxCbCb6WBWukN/6Djm+SN/hMgj5WaW6DybPj9Vai
geVGHpluMfQIsCTmsUVwpLWSIOfHDXWyIn/skQpM082tkx25Xr8L2XA/Ss7X1ug4
vqv8pw9hy1Gj8nSX/Me3B+SjUbmpYON5nFYM26fAvOQ3UR00+EAWyheX83kVE+ow
nP0GY5qqRULHbIWdOYpmICaYjReluTOBNuKQ21nQW6q4A475I9gCaGOBWLESS829
EI99f7Xob+mJr3nNPUq27xLDfSBOxwiZjqz23Emgz8frsMYcu2ynltczzPquF7lv
6Q+Fs/pWyHxEdG1tMAvj57S3vkQZMK03JCF1B7YSY5lbcYpLMNQJ/CiuXPZoqLhN
y1KqEhRWbvO9tWK6UHjPQVMyhZV5dbMyVWQd74Qv04TzEk1oQIO8O5om05cEyilc
hmcozFjXaBEZyHsXc9v+RUxZ7r2k5MJqyRAFL1HbO8VY6VvnL93e2piwJBoDgtne
PEIWFwdepbUwNe0Vo+uP0nWyXAkjmX90eAjdHiSHtX6r3sRXX3DXc58bev510RrN
WxiRD8v3KdOC2ql5hGMUUY4prHiEBgZCwlMqyoklfZZkLH7YoqJyqM5Uf937Zgxc
NbKLbSvcZe9icsHL5D6xlM1NhSsD6us2/9VQt4KT5f8ehsr7O22B7OnUKb59RVXw
p9g14iDZBFD9Ww0peR5+4GwtEqR+TSHSH70sr1/vafRiTPlboV1CybWFXMVrb1uA
OhfN7Uxph3AfWbhDjlGfiojtLLGapnQwejDyLqidxEvHRbIIsTtRaaNBx2IepXbc
qKdHLgLQ6TCmFC7N/lFUzMJK9dpjAT/aswM4YIZzAisyOafc+2SMRwmwz7R/jR/B
fom14hqVru0sfXXHlD1ETgwcLGFUnoqqEgEd9/JoNlLg6SRwzGW4rEjj8Rlhd1FX
+wUq0p8K5rgA8TaQWTY5QyJSaFxxANWorI2lUooDz41NMKFUseDookw6S4OPnm2C
0S6Mj0CZJow/WCUi+5EMka2UQIlr09O84igzWrDhV39uNWU84tJbBvb5GPWQ1uDR
EASSm57LRv7oXwI051916GsrwxWFX8tw9fAQwR72yrt7zQCY2TeBOJaJxlzhHJOT
7ksTkM1dnt72IMHPC37IMs6w+A/5dVQvniEzBS8PtRTWJSEqeznEO29OPCr3x302
jdsghuE/1iwsqgGlufKYfee2JYJHHseF24+XSb88Zy27qgg1vxJFQVzCiWBvIhaY
JwcI1TGDqEIOs1kre2TR+zEx970X9qYvjU6Hje2Lnh3TrpkCyYbpC88W5wzfmGFe
5Yrkno0CPJAxK0nc8vfrAdHDbkxNWsnFIedaQxmTAxy/E06NzgWPZy77OnCEOv7u
IBWyrcAMwmJR7NhJew0fov8RytgwOwmZw1VP/ooZzoMFNs8zV2h58umUpMDA8AQC
jUJn3X4UprZPJLCNtgLBNBQmcCfuwdcz9cw+K4ZiLPoy7iPTtYRqJ0/gD7dQ9qIu
g0GQrQags43rLvmovc1KxvWpy7U/0S8AgjuUOirBC6zYRgbeAsg15M3dd8Ah9Pmx
xrT/2NQRvmV8L0e83qYpsXWFPlVuDzYsquCWx5ykbWLjYARzhyDiVuHtmJCQwyxh
3fTysITRWyyu3JCuuAa6iNmRIdt1uBYM17bp8edvAsiB8pBje0UB+CuGBOzYVxTm
wleq8eqidNFZD9QrK8QbMA==
`pragma protect end_protected
