// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:05:40 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
IxDw1m9ymrEoOVRfmfu3BIrzzcxC7cm19a5vTk/hEUcWX/4pSomzU+VD8Zfyk1r2
IrOaOf8Iw5XdaaGROcoYjKI/JD2Qzr3ZxeR73I/LdWlK8uM3qfhdYPvw6x/HbacG
eTvTC/TFymX2Uqp7uJB4g9ig8baR37br2IJqfwGyUCg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 14800)
Rh2ilwUWDTrQpaTfsjPDojDlEFzUTVyvPu5vXwp+FTQvGwX8XDXocu6QPUdj2+Lr
6SVKgdzJJYCkqKiEsQqHK2wzTAsn8ZJRytUAlEdAWnPCkegMxk8/AmYAeh6nKjcK
vGSYv/4iORP+D5d/a+KjadeuuomSj0wqt3bNuYTO/iXq5kRn4y45xmYowezPu7do
ESucnt3ZsKjggTP3x58jWhcWefFZTdzJ5SBUYk+4JyD08uD+WpJVPuDlj4VD0K8E
w3vScN2chKid00Z3SJbhTQEAwRLkGxSfWSRdvZNXjBsEsj0FcvxwP011GJNrBFqB
CiSkh2z0tN7gvLONk9znAydC8+zBNbcRyPGjaJlFN7ShVUO7lzsgHlf2XHKkydSN
n92/tXhWrO4YsY3CCsAcOgrpeHEwKCHZgop237amm0BNY/WKmCgSQFXC1dkzHecL
F0kJ+y10/I06xEXGeMZt/tfTxGBw0hIebqJpOUvwGuWCMjCKIf5O6h0FUseLSF3f
Z2+SS9FxEPbOiRh92pJzf30a6omoqbShiKfv82K+jZOMAInGoYEluYXbn6TrpUJ3
XRmjKBjWOrHcwqKSY2tGMzcxrXj18cZJOlIzkM+oJuVoIbLBAk6lOVehQ3sg8RCQ
gYNWGv3Aov/tMl7rcNCI00x/ASie1tvu7hcv+1TisrslsI8G7dtX1zFiBzddAX/y
x/rnNPEkihfffaC3938l946sKEp4itzzUbvFbQFxfLNCJkxRPHiA5dfX6/Q4rI/B
K4iYVvFjGluTTPDMa333Ik6sDhRAXlPdi8L2pI8FzMwonh/ucFwPYYB1oxgm1l8K
5ey676bAhQ/rBs5UpbZCZ2lxOr8v6DRvnowF3EHHmG+JgeCUkvyoMaH0V6NHam9k
IwHyDS5y93Uu9mBqr3w1PYQp5SG152i62Yg/ORXHQAl5zG3acuiv8MG2B7FqTpyy
mJ4gEv4aJXXyG3pZNYYcRCcOj35B1drGWEY6z9ct6Xs8aKRBEinQpbXsPiOb+jN9
GO5bePpPNAn/ezBsg8CcqNqKL43OJb3IGaZ399FzpdvLjzjKN0YgXpczJ4tTzA4w
MfDjiZZ4LlAdhOxsmyx3CrzVAZQiwHARvp6XM9JRK4hlUliulJUtDd8oFgBpKrfv
rj5+nqdoM/1Ppl4Wa2u7W/swh93f4saFUrrBVGDpplG1EAhUOKEK/iyg+kfKoNFd
O9X0X/VYFzgQxbSEDaOSJDBzhe7UR+MXc24T1cxPBoqvH9ehQak2n0GRM0GvVJU8
LkMQOaGxr3LnY1hVGvXhw/p5FAv0cwliJx4rmDpUuUz6Ei/ddOjRinBT/eswGv6F
7r+pdeTX7pkr6+Q3oxvGtPYe2XtKn4NSwtMNHZP76iyK56c2NtCyk3XV2I/TiSab
/A9IIeTZv05a/lv/HIpihjbn8n0hLkyd4/5MvjN8HpeeRMaT2/2xWovzBmpPCIxT
18IiwAJ4MMq1PSt4vH9ohhSNawnamKSsMIs4vrSCag4kOG7AXhXN2xkvKhVBTZDA
reK0enpH1zJfEzVsMXQmc0Pmo9vElvJvG1d/aPWIeYeituyDHW/6JTUsEOcgP+b2
F7W8kIzj8v0Dvt3tVsKz0l9uDfr9bsIVivmRG64zBOU9HXkvDCnvt5KN20zVfqpg
dBjnR8PrSjq4g0eJOIMy6m+80vnnCcWbv3ks8AZi8TjgyKY0Zh5mad940jkamut/
jWg2Zl0RunsMPMikLfYPhcuXQyxadxCsxBBjaLEEXLcxnasrR8EMqPCcUqoRsbjS
lk7hzQoP/MUEvfBD4Lgvjm5wAun9vwOIHmcoz/QrmRu5o6TCzfF/vcTu1754nSfp
0Bv0M/umtk5PXrr8hUg2Y9+yJe5nNU3jT25ZcISX8dhMcRtelB2B1Oo9VzS3rX0r
HSqsY+SsFmEwPUv0J76C0+vsePq1+pYFT9s+HY5fT2rFGJiH3Z2js9tHifZ6I+TY
qJO9VREGCTaMs2noL5FwOzDvDKRSx0LQ6ulhkS9PkQHb748SDRvIe0gX2gYrW3vD
nCxtGCqUOV5P7sfIDHr3T3IbEMy0mhP1fy1qbJb0pT04fyE+xd1+0/t90FPORxsu
XU/Ug6mlXtpK0k+e5fZG8XSE6hIzHl+N9YDaeOA6RmPZMnx6XJJLT+5P0c9j7kaq
WG0uEIANmoYM4d1Aotk3ns4pSH/39cJ0bI3eDxp6Mfdi4dv9x00/XPmIkM7/lW1f
LtHXtf0GBaptQbbdEOsXXnNiOKTs4oNxUikj1Rx/ZpdF0Pn1RtYh3IIvCW4wcMDp
gcZFhL96Vh3vKnqfVara5D1bRJuVOKE3NQrSN0EFTB6ESFULuRdmT4PCpVKipevQ
hjJEY5j2f0mGqc6TVFsfIj31K7t+I+bAH6VtkBJE+nTvfGOPHSnGaSQ6MxZp+GO/
Xfl2gXrVty9GGEAmz6kQj0V4YPG5Up/j4bGyeAlbS+6IXyeAXxRXZxon9D14kkoP
9De32ZZec+eyjxmNscNPbIQSvxl6X8G9ShI0bLMMLftArOF6NogwA5P6O4iZG4a2
G939EYuiGEXGzaOWYGpkB/jFpSpAYDqQUGXQZCQ0U8HQ0znkD1qGVXrUA1JGLb3b
XFeTIWG/p4witrdhVhvZWeVxWwPvqmRm3SM7kYYbvG9NDYVfVc+R0vQAylJ+k6px
eWe8vZ9TmWeKuChH5HuAavCgmXzvf7Cf7WxtQLZdXAR+mqqyyNdsmp2xmhOxXtzT
c1WdmJB6AyEut6ve1XgkahL9gvV/gZDpLHrQ8ivaTQk82OPTH1IkTxGMC6d1Krxq
T3XcPGLA0tfWaYrtL9hOkysyZrs9G6c1YZstGhWQHM2ghxPD/gEGd3lKXbOHBJzO
4kAKnTlaeF2tIdxzDeUfIKKVEj63XGR3dG6HDFQJc1p3VkOPx31S4mKr/+2ypjI8
+Ri8F8c2PY9hhuJ4/1+WH1sm3Sr7JT+KZYOagvyMedG5ZvyLZTHz8f+dCQLS1FsA
G/A2DRx6+BQVd2/7wx9TaXB0HdmptPZlZoIepjWvch66LyDRgdH2yKTQ0JXL+LTA
IngffGfEmZmwQzUZ0us2Ibl2i0jLnYZoVIAUFlqm3rsAYZVkS5uSxAAhWpY50NJP
6jwl+oqyKtaEP/+3nTOqilLw0QeuYaTVZCmJdS/7tesGAnRXK0SAePb+bYhAhtrX
93XZZtcSryL3ulmD6uvPJuWPw8U6D7GJTqZKn+uxIc6MKfU4aVphyJP6t4kJrrbo
rfA7vYwACq4mKnnnSPyUbzjyGy67ox8ZgxIjVLlEiQoZA5wxg7uTwBOUObihweCT
wibRStTOzV8waebuEH3RFex32N4a+Z4fFqFClIElTinYJ3YeuSAr3HGXlSTv7awO
/297yVQTHzhvMbWzbU3VrhjBqQmEQCAeYOvd7LJAn71gfw8mz2GINOzdyFVREv3Q
06NtrevfBVmpwkX2XIOBaRv4N1tzhcUS9K4PQhMc/h1pvD/+kvCJntvj70Vxm+AN
spjKLj+mdj8QZFq90PX/KppWhhMBv3RDYQbMaVupJKwdZ4EAOAVTtL+rC7eSVQV/
waJiJ1iocK8htGshe5GmnkIWWWJG6jxZt2FNunhFK5aWQTW7HeEbgyPHrxLL/dN0
FIgWAj2dYqmFWirOXlBvTyrzU3OUhXyXcakGIVhp+JTRKYvNAn/GzeadIQoX45nN
P1+OEHuFnxL2oOanVqM4r5UezpkPxpd4p4l7V4RY/4xjsx3/l6jAOXNc1Ub9Tw69
wRLRpGA1OFl7h0ZbZAcYiyCjA9431fGZ9DrfVxhTxMunn/7lxVpm6SbMgwaRgoAV
zph3JQWXl4EfPUbCBngKM+7wmI0IwHdqZdrKrZtNIBkfW3ZdnaEjIXdTTYaFRt8d
xta4YUagSUA0ztFDpV7aRrZiidU71n2xWi3XlTb01XmCsPSX9xFL2FkOHNIOCg3A
QwhrYdIfxOKa38dJo+nuZHuJZDMLl6W8eJO8tzltpibrS0DSHS90oxt3vfhOnQY+
O+E64aqxdY5Zn1i2j01ZbkERTd+pJXSmzYeP7IV29eWwlr9MEcvbUF5rCXM1eJ93
fLCu4cZgVOA7I+wlrfqCbDw+7GwwqLzFJVUUUuTzfy2xARWwsf1q6/C/135mwE6h
lFQX3MZFgy21uqP748I8xyV509swRn3056dH7DTIEyWxKNVmCGUHsPFdhlTRX4hk
vQE9exABu1+8ETEOH2qY5r6MA4db5k3OfoznutCHxnGz2P+n3B7OrMbSGJWSw8ss
4ay/oJ288RepKhvcrKnie9SvIazxon0FSmv9NwrJdelmwPE4gE21Holo9KSxThS0
jgyzsm+yf0n4ximm+G9iGtEThJv8uDN0P7QVrt5qOqfUDg10u9F0aUu+7k7GEDOR
aeKrc4Ap93J+9FfRn+NcV/iV1gx6FFNuZEcXnH53wRv1b2jyyA3CgWql3HGnWdJH
iHm/O6AGD08+zm21XF3kukxkoEtOwjomzJrxgnPqpPRBicuiQ+MGFaEcUNNN6DWo
sdjbk7ZUXcjsVYLJL/TwjS8jPo3FHbSR44X/MAK8sC0iKbcsat/q5daFVy1UEbfU
htoDQ5RucisuDOGH21G2QklJZMR3qMDnRQ741sFA28PffQKruWOjh1qaRUBhryng
EvBfxnMAVkMRbrv9gMgjag4bNaA/ztPNavjIYaGhy3Li0b2hFG06mOG3PMY3w9L/
4teJkZla/Bvxk4VlH2EsOx8DlNJ5NrVZkIIdjfYfyxyklLk62q/roftPatu+OA2n
13qsFcBoAKPRQCNLD+0NTEFELMdHjG5ACsIDQ4uoeWYrLBEcY6x8+0Noar0jdSFc
fdEPCUSeAoOKgFCcyi//0indRNiHNP3gx1Hfk90drPDf4GwzcK8JJgcMuhJmOk/5
YItPpk6QcOLXAugs8PVgH7VvOVCcSyHw7qlxE0zZfmtRy4dLYGFuRXZzuYKxdKBO
dKKyY+OqB95A0TOj13QMY7iEcajnzl1K1XHDoJlPVah9b0Bu8zCtT9rV7YWHtWra
0TtrccGOMvnAc/5N2VmEkBiTWNPTUmMKYeFMGNzN4ooIpipPgMVWyT2ciCSDTHMZ
n8wdCuQk5JXP8uUZymeFQTt2mYfvWQgN4eKqs+MhDUAuMYoR69GNqnnK8wmX3zED
1kTKe+eIBEX2Q31tJwF4CtA7DDyl4gvFwdHB/ySb8ahRx0/vZJyxG1NeSuaegLBW
gFPt/92GGrSZsI+fzj6mXh7pW2BKCZTmwvAv1ulYjCMXSKnC3/k1jELMRxlj2pxa
Sjglw6smeMRi8zpODRMZcDvH2coIAhOEZK45NrdmGbrvMZwGGiIysPXo2244/r6c
5CF7F6PVAtOP8DswX4pIWUUR5ch1ANB6SPFUZThdINpmsbocrMgDcSaxluBdCbzE
C9Vx/C/oRTfnIKXllN3pHcvM1tKIFpDqiEnW/97RRV5byK7/8ga6/40NfXPAYvdm
8qqa1uYpZBQAsHb8eIAETV1LU3avc6GwVh6+9MMMrDxSCtp6U9FnwfkLGC38jL/s
fR5H2rNFbosKNve398/LjIpa8OEnK4tKYwwDZa8QVw5J+2dxhZqfiEY0R/YoCoiq
cMswGDoIZvbfpAXYHmjripCYlR8VETH5eddFYwkIhAfqxln457lzLnSx+aNbXSKx
sVGALCGk2CDlcH+C9hKFy9W+U/wLNqkCIx4jFKPH5/MIASY3rA2EKQpg2c0Firbn
8KnpYpVU5Ae9LHc+Y06pBprkazvJXQry0i/EYwcL7Hc9fj1wyU0FxlPJkQCSMtQz
eEGZ31x2ygv3+Sk4Fm7n4PpGbGaGsxj3WcHudbWNQg2GQDR3R5xFZhKoBNoETi8n
dmKlUFgnMb7Geead7ODDq77uWGxUFhh9Su+QiY29pCEtwjnoOBP6vhDZT9pIPtn0
m8gX4dqd8xnosdN16b1bBgds87eyQqcandeyxB7gftZIKttPB/epfEQjtqsWeOoB
BSZon4RvUVoHdOyl1JZsp6Nz2VUo/zTWgA4frf7rWeGzysRA3qtnSsuBNimCad1T
IxGCv3R0aUDlo7LOsGv6Nk65a/K/St26roHB0dLRQfI90ZU74/esmLz3NXWgygpf
T5iEhPLaPsQUiUaOz85SU7vGtkFKD0KLQKHMuDeRTiQWLnWwdL06kZ33JtAZ7X9b
hiT2b/Ed6tF+FeFUMYS0e0udKPjayxXvCXPVQtz6enJZxcYWHumEn8lGYw8/MiqQ
D3N5aXO7Kydt9IJsvP3fW1XshrKK9hPGMwNO8t2/KxjhEie3XbtStEp/tZesi7KR
Qtc2wLgE0ONcqgoCQcEYRVr0WiCc4kOWJeN2q8rj3+mJ7YAqBI2BwKU7IX6Fj6Tr
zHkm+JXr25B24iCmktOcR64Ae9Y1miUAomROiW19sQ+f8We9m8MRP4jXqUOXYke0
FypNTfHaN2mNQyVGh12Nc0SNsmj2PQQHaL3tBa7jJuw5zrUQf1x9Z64mzg4fZEa9
/rm1GNoPnOsXZO0Wc8P9kRqIbpaftSMpfe2A7wX+khaSBFalZ0XfQlUitR6oDncd
Ot4JP6LSFwg4Vj5jcgsZ571BVQHT6XGjqbyWU3e7AYFZNjusFnde61XFDkTT6YC+
dX0d/MuLmePJawhgmCLm2uwwdgRQXHyj4cEFrgzqOzCmHiuPIn9ySCyqqH2+hniY
SwQHmtdtT8KCv4SriHR4HV8X52To1bEY3mJhtPmOnx3oJtyEAicX8Ta73lACfoIt
7GlYwyJkV9jofk7AMt/6me05pkDBA/YCS+6Y/J0MH3swj6VlBNgqX47Vf7CqkLuG
qcpCq8DY5C8L/mlnjUt1+f/bX70SgngM948U83GhbIhnmoFI6vWMGs8rqwzHE1E1
s6NeqIdcU0fNhipIwjxM5/cWmN5pSu6xTcqtA7//MVdF3fUk4NCJTobA47ch4Ooz
baIxhiHwHtW+aveIGDygg1PKHKQkIvOY7ECvbV8g6DduaZH9Pe4t7zRK+g3AGEW/
J57TSxWtBrhRcdqgV/ALTsGcbponLInyytvFUA0gGRGVv9/b7v41aXTbD1yilJj/
MwBbEXLU0/G7imcfvoCnsMF+Vj3U6jXhuQT5aZKst8kKstfn+9b4vbFKEbA/RPGR
TBC1bSAYi6Lca9o0XjECkeLI6WHEAhPrLBAeC1MLOcWANMP2A5GcTJdPE8MuDUrp
WrHGo9yjJem2zasPziovzYpS1Lwi6/kwUyYgd9KkbSiFFjbhS3XnzfGGEfiEjCRh
9Jh74ba1lFPBdwyo1BrrzgsSKbrwRDFBbcGJF+PKIS5j6t6EUdG/AmUAtPwVR0vG
tLayc6nOvZegJ+vBM4o3Z859Ki7q9GbyHXKPJcZ7kIgm5J50ac+OEhIr8Ls+ASWy
1QSfekc5HmtgSGDeR+xp0rlKuiT5DyX5BQ1OtmrHXTxTG6/u5yI3ttCLQUusrcnM
G+gXnaPslR2FAkvqmggNOsNlVFsv8BrlB5zggsFerSP0ypI9CE63jwQDb0n/33pU
3SnMHu78rAiutJCQcyFFiPxt4keyUVks+XxRaxt2WMUOahEYWvMTtYq3+XIfSTnl
g8y1jnhhrA3rZiCHXn0X8vbbwT0xlO5zHByG+R5gxFzlVNN/zg517MDu8qcolnoT
ynQqNWeftvd8KymGrVvzK1C8wHYpdy8zo+OlR2xdbGTaWz6gD8A8TncIk7iPlEzu
oLToXzDtx0ynkP+9EMcvp1fourpoPz9l8V2yP+iDftGTIEG9oil6n/oeweum3/d3
3xjjARdxOfWVdV/lGQG0DLzl5FrMxoQMPUupOCPreCeGGE+1EBNPZQ7dH75m+jx4
cMUx3fWCiH3gGdgRU8o6x51F/06Hh/DJPLJVJUt9ajEjuOPxU4kCwwXWh8yelsWz
loqPaLd6HsVQJb8eYQLPs0ONSjio8efVg1bD5QkuRW5/FBrLtyBOup3ynktE7D8E
sKw5IWgWy5AA9pryMiI/j7wJzQ7GbXq9oWgJZd9E/Ehv3EWxe/4JTLMOpYhDjuwd
0TVFFZ6ujLMcrTU80cQ9Q96zb7Hw6xIO5ovCdb0qkdLSHkqkJnyNr5sJndWyVDOu
l4k8niiEhkrklr7A2Ouc2BLDRazNzpXdJXzHp1juW4m6KNpF5p16jKT4CD5ACqHP
zskZwVhCjSWREpO0t2hzfFuchuCTM+DOwHEpO8ftvp7mS7mW6HHKU2YH74kE6+wb
XG1uaNID14AnGmS8vkwTISKX+bagqVblT/qNpGHE25KuQTV0PKdot57FG37FjlD1
3Vob7f51frlcYYv3Q/nEJFp1CxMv1WcnVDpNv07dTkaAq9eqPC29WnhCLTFNCUa5
16B5FVdSPNVTyAq1xXZQ/IAlG6LGPGToycqMNiE/4EmMzUiKD5U/ga51MZ05gMfK
A7iQ8V+n+4poZeWDnMOvNhhk0znzlIp/XQuJoyF/WxZPobwzHtfMgyIaDN8i3URn
uHenXgUGMz49/bhL1NSOn92iqoH6d0QQKAEGljIRCP1BkgNtq6gPPlripz8Fjfad
P1OafO914iBl1+pKUQljNsP0R6KGFm2+Dsg+3te+IqBydlj4VzlJGP9eRETMB12h
a92ls6/1VywE6whw67F0/n6jaHCp5SDkxikICfECWz3j/d4C7gPxBphN5JlqWyqr
gf0Qk+AaeA0HTTbxpE4mJJ6XAXhprxSF8/QhMJyGnJBVPG4yQjaNx/iqSQP59q9t
AGgwkbVhzr29QyFAi3k18P9llhcWGOx3y8HUoKt0mFX5sD1OBjSrjT09O8g7EPdk
b6RUnrMZZdsgBCt76x3V8PO6lCeT1s1pqjeUQS9gp60XrOrcBJ/UpWliIGFfW/P8
R9XtG7jSZ3CCPBBe9fSUWoxvCLGR0nPFKxIMvNq/cbNO7JpvtIlsFuCDY2ybngfV
Q4CzvzNCFVXEStyA/aVlmx/iD95ZrXC07mvDZQtHcopkT2KKUVqHMjAsA1a7QvLx
wgOwhVPkWqvafizaeZLBLz9F98VWtyUfUPIRbEiTsifr12EneHvANmB0yUaxNtOp
2fv+w7qsTl8Zn4rVPOJpy7IGepTO249+wL4Lf7key5cCG9M3DLsg2uiw2B3pkI5Y
HpPuGxUNi06fDJn+SIUJtiv36PneFVG0zPFufWkCdDVi0Lod/17EVlD1z2xuKgkO
5yGQBDVF3lyr3llKGCkDC2A/g/Ye2QZdhpERuo+24ttRmTxTCmtPEsnWDK5OvvuD
VU0QklFmZwa22tXC6WNeg0ivLyuB8tqzYUtgYbcvhv5utD1YZfE/4n50y+fQFA3T
rlR/Hx7+v7Nc8DWoXxL06JDVOUHAJKfdCxQ68IbK7pb3GMDOlRfl8yP089KtcBJ1
TRyo3JUp5chReTuRAvXj1ZcF+gr0H9Zq8OBNzFikV5PXDX1lpSPJgSsgUmbmSZT4
C810kV5pQO4UZrVOEowY+3nrdhgpBFxndXJ21UJHZ+9dc3JkyM1+xelea7izMrY9
nq1A1eqDby3kJyyOm/xv6l5k/eqIdXfCZWnOOGVfc7eU7LNkGwoiqHR337Wt0Ogq
Gpnjv4kxw0W80172Y/YUVsTLa/l1V/T8ihArBKKCIu8VWpe+Gva2qMiqR0rncdGF
P4ENJceNEeBZGxLRwgKqyCmWgzWHvyD7X9ctYbmeL2EQpV8yRcm5n2ZrhbO9o/mu
CZT6cdwmGhk7wMuOWfjTWLtni7OZhv1VYqgH5KbusVpXBgv2QaVqMqBc8qTO+g7J
1G/7kP9cX1lRTgZdCrwrYivX1HelUZjg/0RWcDgkaGol6Saib0l9lkNba6nykiGx
eLUAK5W/xj5rdAaF00trSB3LXpD2QJ+l524WN5mFvRYH1LeoRpA9FxU8/Eoeib6V
6V/Oo7XElZ4jzLYL89TcG/8P7lLXfwJ8I0cSpkS8oHdL+RucAcsQhXUT1gb6uDaO
DFW4+z1zDqIWYvrnm/PK2B3kGFTAN10vz3+15GbjPSfxiIoWdrnqJ0jAvWP7h+0p
+FMZL/3rsGx4e8GmiY4ZIXUP07BMl2EtaEVnDhBZBt0Su2cb92Ih3Vv7qYqdKjn/
2uApS6SIt50RPyEAlLFCBOp6V9hZuohaKuwGr8lDpLzYVyE4ZLcj0eu2oCAgJYLy
UH30ME3L4wLxWF8+gPNe/rrQghZh6JImHHpV87A5fQFAo+HbooD/5qUIom/3Yijz
5jTUipv5ybVFCjw4MA6a1mia3t4huLh0GuKG0vD1ge1R5urawXZa8N4y7GJRYno/
jg5mOxZuEgCpzyqdmRmZTUExnI7oXr6hj/pcExICtco/XSnGjc4KUb69fqGMmDMm
TjFYWqVJpzUAkY/gboGYEs/raIAuYTjdIs31XbCIeoD+7NR1pyIkXgQXOrtjA60I
ym0RBdUhY3OnSrAKJAlWAXSJk39BvsgkQzTB4JX42d31SqAMrDVkfF7Riw6CZnfO
caZa6sTikvP0koD+EWA2igzbDdnOXsWYTCJgmdtWXD71KJtSZjP0723jhjxO3ogC
xCMWrABia5/6o7BDyGeJgtyY8OvV5ZgfKWA07YA2BhUiP2861N+9BWHudZgqOOBN
M43EBfXbhQjV6/HeMX7dv8hXULNRs/+qFztyZMIWGPq28Jbe/HR848YyvYNz7ZQx
bjGNx1Z8Ewi+e/NtLiaoETw8UN4R9UFk3DUQJOWcKwdxty8nVV8CesRBzDO/I8nq
lHXC/29a0vbjg4Q7aVxi/IBExEXbgbuR5Dy9FJ1ocsDBKoPR968MysphHTtHPva9
AzchKkK+vewo+11IaHB5V8pCk4EUsx+aU28BG1lHTmLtQKbXzcBqySzIlYDZhu70
th8wYUxSeb/QBYxt6MidZIrm2g4m7wd6ELf59bybAlHdSNa2zmsP5r7r8WGZOi08
tLdmU+ezhfBrWcr5U55iuvaK/HsRZs0QaEsoo2tR8b6tBXoFwrCJBk23Rz6MJ+7E
5/sNZCgZVU7C0p0eHO9okv4SW0u+VHFtuJVTJqGTxz8oGmvLgM+0E6DiGyb8Tvxv
wY0c3muYkBtvU3lCPZfs+sWDrm5GJTqoEKlD9WLFH9h7oKthex31WUF9OGGioPiq
FxhefALw8RXczmHVZ5tiiAQJoXUOlfMOz+6oq9/KPqW09ZzHW2Q9bZgCH2L6se4T
Q3vs286bk69tq987+dvjMEg/ObkRrYLenuUU/zWa7eBO/DSbXVsUliC3BFgtcKW+
hmS4UsuDwZFJXw6zx3NusxdCFcK8hUcWFxJxi9yKzJS+gSf+r+1+nouwVlb2MnFD
N2SpenUnwBRI9ieMpN8ihhF5ZYd2tCTcsJddqJYZZTcRXnP2jLfb7+VCpfkW4ETJ
aLe2KofuSr8MVhbpTalBT2lnqoXSBohGs+iUAyUNCzSPOjTPbmOPJALfNAGX8M7H
LskBpVfQMEB+pyjGvzYqWZ78xvwfB/Qk81yKSae4splOpC5vay59lHZkBZ4WRnab
F6PLTlevYAGpZNf7D32LQoc4LSqne568NzyW3vubym+bHCaJzOHOlVF1Nz1W8c37
ql39XYe3jfnNoqxxBgq8oDsGglVLHMmln+NgA4NF6MW62nMx5SsVQyXbNl9r64eV
v3Hdjk2Nr4VqW4ucUSS4+rmykaOPlDYwlzFYrJPWpubL4iLUxMWnmXhFfTIScPsa
W1dj8I/iyptgb3uPAc0EU6fzzMiW1qCeI/bLeCvwlP9ujQYWCQqpiJCF7dtC/LhL
s1+qsKlnua+0mzI2nK3ignr+36SqiHZMagguxGPhxTEYzSn4evWA25w7o7Rf/gTE
K68+AyW0kDXcZFarZMpDH81lU0PZRRX1NFnWrbW5l/RvugTX9kVvDUWyFuCliiR4
zwotlHmtaxBLSmH7k23DCnTtxVQXHzJQkEM/pnDERYje/aytSqZifposG4VY67C+
zaPbkSJ+hew9XzQ6wfkhx4LglxIzbL13T65GMDh971rNO2sZUqOxP2bsAo5I0mYp
v2qOf9gxM9tv3UcUKZQuxNlK2TEFb3tlVO73sgdGZvrUp5rKQVlRdUP+v+hvxQJQ
kV7pxIQbaR0WJONvxsUotWq3zT9kyLvG9WxG5/kL6tcSf7VWmWzJUTUiwLSh0xta
f3YXfwacRwxbREIIj/hnA1xETPbyQyzS3BiYJ4XGdq7kvfsG2O3I3Cmf2/UQqS9b
NFYBXhO0zlSczvkP3+WrtR6DfVfXkmYDpqY+qek8S3CFd/chTJMysjMz9eazQQOI
vQmqvtPGjfd7ULe2EWZewi/cP9s1+t3/JfkCk/HiHHdnu45lqvFyn6tVWHRtU3wM
KQ5WZGrKOLo923hyoqlFrCzd/tfg4vcH9sk86dYFmmPrubvbiBFaCKy/r22GgbWZ
PLesCinQt2kD3uEYIaZV21cNqIefkuWGh8ZQsIaYPb1XEzOQ7NS6R9cv/tTGfQ/R
w9Z/ic6OyrZ9dbLUwcGE1ruxKJ113pQX9HOOpaE7Fyp4vSgnFf/GISN53YyYJ842
bQyJE5Fkx3KS125mdH2X/2KvTItZLIXptu3H11IXTZTboENb1ugHrTWYxD7LFob7
e8weGXyL7+eFh85Swu6ymVpkMSVM4U07/eECT7viTHaqlK1iBMxTJ1eQ5LCcYK9O
OPHmA38KH8YhMuqMhq17IVW0SRQB7gaCO0c0ZG2FFPHaPJ/XfmET0yUbulwTkGb9
RfcpEYZfHoIJYwjwdmkeWpENu2FQOG49xVUomc27aPGpLQ1xFlEmqZ8l6W04wgDb
woqKcGzGUlQhs7j50Hlp1OS9AceI8t0YiCxqcg336cgB7HULTOlHnyR5YIFfTVCv
Ibl69LpLqlNvYnQIRYsUdBO+aP+L53cgvGK7z3O6r/KI5yXC/eFFIqpFrcWEnBDN
W1iDRd4ncfYYQ+njr1FjPwShNiXrN5XIvKWINyIBoniOdMMr/acoBHN7D+4BK3Xn
yPwzC8b9hRyDUyZ457fQenAVe9QkPzNQUNvXHWsymm0hv6AbrUEOCMVd9Zyru6eJ
y12E71uhu+X1/WgRIcl9sjiP6lJUT80opVRADnWu1gY7CDk4xeSgdZ66EEcFFRMl
iUcq6HYuXruCdLbfDEVuFDVBdoVqgRpCkArAeSORBDCMq7jC8Bv0yiEuds82h9/C
q2Fjc11wEdmLhXnUUNxppfzaCssZpxpPIXpJJjdhESME2A5555SlrLD1+2xCpYco
k84CXpY7fIl/7rjjqYX8MCugYqPbvovy8Lo+962j6uCGApXpEjOLnQ0N5n/uIw12
Uz3owiIrvCKt/jFCTjHvoELalUb7ZiTUgLsLvVTqwpQlKK/VIvUPqzqrHFgBscsQ
Gh+fmQrjFVjsLZmpNaoNztghkIUw8DMQwvyMMRKUtw5u+5x0bG0JL9oJFq5lqN6M
6hxSyMa7Wd45q7/A5d4ud6Jn/NYQkYpjCsnfQPYXYsrz87093Bq4RItKuyl5sgcm
migkrN0tvspykqW41rqXk3DVQi+/QBKO+sAtKy1aExil6GTnfbZXTHVN9KVZeZ2Z
OZmCBXD0FtpwBbq+4yt2Qm4niGE5u+YprW+koAaYqU+gUudDgCLNbNo7CaDvLaab
nQSeiGqrDIYpO2MuM+WR9QIqW1pDOLoeRG9WByfobujKJYCntqau5UAQ2x5AqbGK
vmISzgzOdZyF8Xnn47AiSzNTfsDiPbpaYtAC90aACbeLysXP2lMF3V8m4dxBq1w0
xXekNA3F2gK7wGjkR6LZSmQcftzcjvf6/63xpnc4am3xIpA0oYb74DcBB1jsa28q
IWLXzszCMj78KFgoOK/q5/DWbGfHnbkOSgiaixGzqw/au4YRnjqNwgHVzLCiOwsi
M/Jvn9m9O/DJ+2W0pce7cKrSu+MyhwlGwvZ3mP9PbU6KM0TGdAbDTQpZEo1GxIb2
SnZ2D0L64f9OxYhNNCRtalglJemvlhdAibl9i7Ur4lrgj6ETdfepXv3/C0hu0H7s
suU5bYeWhYWsY+QxKSx3IwLkahIgItHU7QP41sRM+eB6eukeEm6k0iajXskNik+z
kubZkRY7Oyg4m9JG6i6RsrAexYlg1zvlmSAohl0nAiVpeZqg9aeLGcfB4vhYJISd
ywnJn5j0cOT2NH05/Nx2+eIdqIt6mv7lElYlHqfuE4aHkJ7aHpcMTlceem1zJS8A
CfVjiEhNWcvizvfBAL0b5ck1FaWp7vLNbf9Gksq3IAcJUTouxcZ+bvikJ0T890e3
UvWDwidwJ/bCDurifW014rhy7jAubqxgUT4/yKGuqUcwK2VuULf68SjGhgiG0uj6
7AGEXGBJ1bfsuZrbmO38DLe/S50e4PUyFavE/RJm/1bl4uDHdzzdm6/H0lgB316G
8VM9RFtXvUho6EsqGWYrXi/aedr2IbwPnnVt6FkmH9pkEjeKqITbnyjd3XXxF9tF
qiy8Zc+5g525W9SiDY6673/OZGvUGNQdS6RqOmc5zm+a2LUFErq8cE9OtcBNTf6f
zztPFcVijYVlF/1gkDr5uasMTw1RYZfGXZ368s7eMoOIH1SHBOS2UAB6JrDGdQ1g
YecIr8Ty9CRCy+28vgOdPpuDIGHx+JO3G0HSuhJHCiMVDsk7rOJux/7BDE73FOdI
Cak2YFaxvZM+sjHXaY+a4nD6g2pe5NqO7adZdUEcap4v2R3OP8SofaFcGHbcZBuy
fcwLXxfVz7Nw2fc4t7xoumTwhStBmzfOXOmN2Dt4uhNNX7Dnnu0lfW6YEIjh0qhL
ybuEHv0KVZiQQpfWmNlvenIAgvAGdnIhR8nc3mjIMXrQXqAKoT46MmPOfRhMiNTy
pzeEzsAq6pIKkVNryoSMNNT/p0/qB+gEQzY1N6l4PKNoyM+RbbZu8Nme0PxLSYGX
pSYbI+wzbUreeWRyP2CYFuKG6mLgybHEAd+6UflZHS7PEmBJz+t/tCr4JaP3Y72V
XaF0TbHQpBKaWbbsJ/RiBzJG0yE9muyAQniqIFS3yLlTl6qYCW7zhFGiDsNBA3k/
dLQy+zCKQPsK8TxUbHXvvoqQKh64O+2k4PZNy3jA39MS3iDBVkenczoPXfcsHNel
FKhIic6RW+7QjCfUBZSoTsQ/RUIrl0G+YJtQwl+rGow+0f9WQV/F1+EVhOlSGDnQ
Axdejon3nH7fs6m6tn8FzWOIe5MpQxNTEfJKWMog8GGGdKalYc0ttHmL9BvQ2xA/
JNNrQM/y46ptj4aUhMJCbITFWInQq8yP+kFMACAsOU6AtE2emt9UAyPitAV4LysJ
mQ1G6bxr1vCKQzXCb5yE9CSiVkrvRiD2oW9KcODNw+9JL5NPXbqJbKLlb/vHmiqP
EUsRJw9xowCWMs8QPi1xHWXCW8SDao87FKkBLYBi5zY/90ekXt8SN7bsZkOsVbCd
m4PnKG3BkOQw2H3HnS9mjUtCBgcLkghsPAPp/igEZDGmuMS+mj9+UbvH37FePugG
qDpTYjoYevk8+amEfvqpNG5ySZ+ywJp1J6ew/V4EaPHvFwFrr2Bz/SCdD+hsxAwN
gFCOtSxUM9D6efficELnAQho4WOAnYpTfhJYjExo0jqcPHImfoupHBrWzb0QLxDe
EVHuxucmr042mZ0vNFFRjyGoa3Pu5MEb+y7QGKtX8HvJsmfp6c8Qo7BAsYQnShDX
9jq/gyrvZ35J3PcCDnbw71LL6qvn297YzJ2abeGxYwC/tXvkY85x6xqmaaBhTdRV
FjbocIaOMOqemgVdbdT4y+QjLwzupYMabNcbMQcaAyVvMYlMNQ9pZQIB6ogBAEAz
vkDRo6LCSJfUuLu6Nq6CfnWYLqPrG5SBFqWucvwKgBStJZbPIg8T4GfE1z+5nNNt
FUUyX4ErLHeJm//owSRnp4YucOTBDb8a+pYXCN7AxXIcQmA3bI34QfSDGDDCYaQR
yl/5AtHn0NC5puCZ4BoOQGC8pcYUDcCmSxvX5MFPAQHjk0EBqdaAq9H6smUd+At7
lxrmu23rUN677x5Z5H0plGERoFAr2KvjXowGl6Cv10cmhQa6v9+vfNYbMfyv/2gS
3IiZtjbdj5q42snpzrX7IlTkGOYvHBLpLw4UVGpVSZgYheAS1YvZx40y8jQ/Lpr8
fxt9QsgLvT4/gEJSbvRGe0LqVqXNuAxM3iYtTz/03/hMgMFrwL0G0UqAW+OHq+T8
NfuaCoCBzAkkM7X4AvUVWTo3Lke1cCnlTC5bOoong0CunSvqE7cagsngWmNxc7+B
bC36x7ubh5YaFoNPdCma/ffQkN97MUibuHl6+CY+//BRUJ8qMxkSumDfDKMhrzUP
JasRKr1AgywU3m9IRy7Wkj385dzzlCMRKf/ZSdg7I3gwTZSddO1R6D20AccHmORF
gzLHNkyeVl/aRrCoY0fgc2NJtNggyg/3HcFKRieerWzm2rFw5BYPM8AXRjjIFqfa
OoVNRD4I1T8SczE6vZcuAmcOesxkB8tpmrq3YMlaNAjS3xTsySWkcqOF/kLnfiy6
kVtHRL23tq4+l7SIkcpru4WcFGLQbCN8RVaehzhEbFTj5UKljpVFjGWSu8y1r3q5
A54TZ3lV+AvwOh+/iQGvA6vK/5mQ7a5ncHQzHQRyotfeyl5MAem1BLNjx7zEKSox
Du9FTwMRJGJAJXwE5rBoKwUueXK9I4nMPKyjxKddrzebOlaSDdOGXJc2MA2uEF5m
hbk5UVCN7bhNOIZzRN5qtL53bUrldz+coGF3RLp+/GKPbrFNMhuiovY8zEpPJXZc
mg+rm3O51e8nFmgnTL3ISKOe5VxR3ON/jroZpzMqgVMF+v7+socTeGxcV4nyZD1F
mupVpsqOr/jVPC6VD7WKtQmvXaVe5xvt7/YhnLNCy1mWVTi9wKG6btHsx4FvY00c
BpFog4SNpNH5NELCcASb3GMq+zgIj8xzbFx+NZR1b6nn9I/RT03kEjP9QdRRU0Nh
DSQpwUivrOCjsd5T2iyXXzy64ykSVIkXAhef+qCrXRyW6aSsgXyZBZ9gIRd9Np0Q
NhIKzuVBZDBn9KxLeou5U8iyz66mQt9fRybrmm24bftb6IAV8byJ/iGZe37X9j0W
JLV0LOypldnC8ms3t24Z8C82ftDZqEWAESFHCu0952ECXMBbqefxaUs0PA5qUkFG
gw3JIl5k60B3bRK+DyAXSKgnl8Tf5WgtfiOg3S7u9V0IIwDEXENAPyeAzzO/82u5
do0DNYClVgQLcTuFDg58r6Cx1jfZiZ1m2O5AVPpkX6BvpiZa4ZbvVUXEb0to7uDt
oOLCOgLbQRTVU+CigbTVDy7VQ9CO/99K0WyehppDWQcqOwtXzdKsl4dNa48RPP5m
LoR5EyBSTA08QUCsYnaBNyTmAIx7iy+cgZYgeD0KNoUQIf5rCFWzrAFR/RLk37ZW
+koS3yy9xMfbRZ3uL6IuWLIGMrgzaz0azP0YTNkdc9YarqLPqpl/9GvL5Jxmh9Cz
GQKz9eoRu0vVDw3ABSCo7OAabrlb1hLXBuPhLOw6tcaElKSGTM6Y3DSCPE5DQlH/
KX3GvjOB9gpxGDg84/UasQ9ZdKFeH1NQfudkVAsyUAguSt0kWQxxhZkMKivz6Niy
uSZ5jVRWUbHxtYkDWQG9QqLeS/aDXeyQu3NasQrHCBVZucDKKY4Ued2Z8lfHaz/w
kDvsIPvax8MSzXE3IF4f6Q+LeEQmv7tj3baCr5XfwyvTcMya1Ti8QGWYyL4HeMHu
P03Ihe5f1hs47nyRND64PdbKXTmI7R2x35J1EMZcSrH1bTZndh0Gyr+FktkxmTA9
acyEAZmwdl4IWapr3AzPxUY4Gh9ZPVLNpP29cUvPJiDTgfmxNyz1xb52Lqm6U01T
shvLBqz5Tw0mNZwHo3D+NlQEcv85T3sesEbzpKwcoUYWXkikHKViY25LNqj0QBhT
IcoQsg5VXRTSqIkhtRhSEhSAaE07tcTLc/a9GXAP4FKS2TV/NkvoPKPKDbdK2UIq
Fwva7zwUxTff+jOqNqfMqQUTvyZ78fiUs/cd0HPtPl7pqIDSOc7Qb8qg+DsBi6YP
3ShhRMm2y+aDWJ9iV87iYBK23BHW6OhwIgdfPdk+/BU7QemcawQ3DNPM16aYHbkj
ghOZ7lNROKViP/RWSQdIXe+dFgA950FaBlJ+MWAnSIGNamdDfvBrzw2yZvUskmY5
ix3c9mfNrt75s1J9rwQfwXgvElBXz6qYPNJEL6uegX3i7rWSSyu6qS6atE6EyILF
JsQMglTebZ+nACqroCnp1yW4M95lwlQJrmd41GghYk4llfvIjuragcBTWaOYfNry
Ou/51y1tiDjBZR8JHQ9p9kbj/yg3CMZIwqzNXfgh8iLRbeoxzypff/02hxx2KEu9
WtIA4gST+7Hvkgxt1odiNCaaMczx/jzG10HWxgXjOif6oNMawljFEcm6iwZ/uKma
VVNs9iqsfnB5lUYZJfhOH+7al0gmsg8jveyCGVe8rLbXDRw5rFNypiE6cjo5MBpH
6YiEVMUIUX9WCukzL7Yq4U4DPsjqV4AWPIf5q6uOlsfQ1Ht+gBpf+eqquyAkrD7q
o6Mpd3ISgqoWTLb5jM9BlVpYrZsACPLpusWOV+FWq9ZOsGoISsATLcduDravJvaR
kfujbRF87kUAlREOoRj6oxcTWjNC8oQwsf+0hIaQ9esL/huWwTDjnwRe8kn0pqxn
y6pp+fjX99LfJhVSIiZq9hgnJKALyctqLQrhnljnlSWOiQWzuJ37YfvbzzF74+53
d/y9GEy5ttyoLysDNcvhAl/jZiV4Ux05BJemEOphhFcqVsRAJp344HD6fujdQQdS
UGT6gR9aTuOp1C57L4/RQW0ICNNKAmfjzCspX1WN00o37TQARO/j0pJHTzF1ZN6R
60/AbEbwZqy6KPp/FmMS4l9sLuCTIIUF1Xao7sS50dHEENWtKjesY52grwWP12a/
W7Rbw3Se4Ew9dYhJ85XLRzmS8uOsJCKbMXoQ8QIiPVTfvje95m2qsEa5sK0Mg8dt
GSR0Me9LelATaRZCalx2GuzTaMLZb+v+6cjw4530q2nvpIYRKDFHHRnHIul7V9BO
Xd/N8cGsbcEUROKWStHX+9AGevnZuaZxEPuU79DWdmRVQZOTDEw2DV9es4lg0K4z
1FMAxNbk9SE3UqHe6KOhXbu02d2R+5FxL7hucSIdMaDnYR+TQcYMPrl4sHF85WYi
53CdbpxFSfXOYcLlgzp6kNXa65epk7ByliWal9EuS9yVIs2ndfT1agu4G+1p8fS+
CNHC4S8F4fWzX4KgayI1QAEn8Qcq0EyGRY7gg2zTspP3EcpciI6blTY4PEetmTMU
hz1jdUgjH75GX6G8+AEENI6KFGsGOKBaxrF0R4mmWbIdCCtlL29YuboPbjtfqdiG
/HsrebCUTjBse57paqPGDLQfpwhN/xP1uW3il8IBUjbkvkSrKCH3W8rO5tA5tXvf
SSKM+GGLGYItffHa+Y4Ufu706AvYIfrZVchZ8qfksEcmvePk8RbnBZzT6r8gyw2m
aAaqiHkUg95c37a9RY16FBNUIaMnpT5wf9AUde18LIoBn7bTpr/i9fED4tyaLOgB
EMCPSVumbJSB9WTA1kIhGhPO1iMskKTxYv8Uq0hh+lo2TlX0C3pkmUj+atZMCJS/
wxt1NhmOZfg94hLcfepTjBYzFXGOarseLHtq9InYkciUVu5CuWMurHcoWIztScOS
ICyorynZFAvYNg7rhAQTLQ==
`pragma protect end_protected
