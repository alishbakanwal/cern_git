// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:05:36 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
CWQ59lzuccRGQu6kNnJGL7qtnq0kjho8I/UpWL4RlxBdBKksi9OuiCWTc3pONnXe
jzIFQR3KQapBeHuXfXSws2c6bNqsLc2ZFzzJnO09ODzMEDiz9bLnPSHJK+ygO9ym
x78OG0aRtACFEPb8mCjLbnBqsDPpYGcWBQ8lvSQGffQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 13584)
uRot9jP6flkrLkWezmw/kPwnAH/ike6y8KkHkR+sMd39e1I+sKpkBEtCfTVWY/q6
9uWf2ykF5JfArkyoowW2CO3wdJbBqAUkJNuPsC+owHyyYKBNiwM4I9F6hQsabVQ4
pO49kzpSS8HKK1MKvSzJ04WOzJqOZiRp43dSJp+nvDZLUSwQKEzPL+fxzssIltiv
4uf67LX1QfaknuYOfmrjDQZr5FOjKAKojKY2AZXPf46W5Rn2W6XQqAF+OCFqXfd1
YP+id6z+KpEgHsnCWdTzj9ggmixv/LhF3mmb4uSnchla7V/ZO7oG7T0zkPbuEQRH
fIX5EfaqRfrwQnMt4SILHZnZxrdbsG3vgCR7cKWepfR8voovIayTcCgbUt1hS2u8
31uQEsi+buIE8aSdVlSgDfgwIn3zUbY/uiarlSC2EoKUj8ju2TRaA9QAyqMZy3xL
tmvJnhFhZvaCvZtntxRk1iWB19x9/ZAZrgx8TIQ3d+qc9EPpNAmBVx2wvBbb/H9F
F4VaL7u9c7l/HealAa+QuwOGhM9nmXGWI0zVW9O5M0fjzG4XLQa4MpfQUyluXEiE
EZOUvgnB5J0hPJjBeyG2q4JXoWTL2LQNJ8wCwJlxW0LcHEzAM8/X+rdFhcqbJrk8
GuhAtd+sq5IlinM5ueTgWdolORGHtGSF6sYF7+jGy4/GzkyklHBg1yjAV/kmMMfw
UAzzQqaB/QlB7Lcl6FCNihHXpLtadN5HN+1W192p7/FKbvOzhXKz/hihSed5nQ5J
d/sqlN3rqPzlLHm/YqO82B5kHvkZRGO+hgKKHdAxy9q0ld+SS3jSrKuzomSFsVPk
Nnu+cO2VtsReaUON4ewpeXhdQ00/qKOOe0HaMwaRd/BwiFAiw//WTNurqSaZaqwA
tTo5HTZ44sLmdmdpQ8EjIJKTYDP6SD9XaNjyj+W48P7pxOX71yscaMUsuy9OQ0Gg
PbLiZnOSX/D0JVuboO/AqaaPyxdIAVe5G1kdyPIlg6JSr09AFvZugpno29zNbsNg
QS6SG658zLOEezewu2hGikojqG3YrwnE689Pqdg7m6g542Z+W+p/cl+bOd5INRYW
J4hD0BmVuUXLjL15nENa7C8wMfc2j9tgCc4sRAGHezxg0MdnxDggFKEajv2oFJyG
XiprYzUgvrpfJNdfm6T+r4F12fuOuyv4m8RJ3nJXVAd3PNFSfaGXxj/MYfac7O2p
f6Gu0KQbCDEb5tPQT4d+s/1K/53MV08SM3+K3VDZ7gIyeKgW7dah1LvWy46iOW+w
2ltFsYp8T26PBzBte0T6WVVdJRuF/4xgLJy3pQEv8P0FHz7QxcBrckvf3/xBZN4F
f4Hqq5lvYgsHPa4Gufu5tpfbzbI59SuND9Vo8bEs9P/5l2xGKubzmf7idGwLCLwn
gMK2YtMpeTOyrY11fmDf6h3Hs8g0KRyN8oqIUs369wZebb9/7BV0GdPYeY84yfIw
7SqUGRsl/7Vg7/aV+IvXyp6xGlLzEcGR4EUIcVCHWvYh9AAiywuXCj2np9HFJRYP
jP52KSGBfd/WcvGu/dCxumBePqwRyZijg2TGsjZWPc3x7f1kGiQmGViwQX34wnOu
tVW+BT5Z9zbAMM7xpYnqUA0t/eQ5/EVotbTzzl0jg3UZzyuwttbRRrryL1mhYvRH
HzevqM5FPkIYNez0UwROVeZd20Ofd6RWcEK37Rv8GcuUwGpSH3zBGv5CGP8CiHLW
vMq2Axhfocx76LPxuM/9qOf3oYMxqa8Ea7zo1lthBrQLa/ETTR1HhPC56v7M2+JX
WYYd22wSL/sN4wxjRMdjn1WBr85vHUMDkB0i4wwtmE3RBbkFpVyDzorpUK6yrR2D
ByNmwgEwxph7s9GSRgfJj9LDppG/D5CU3GOL3vQoIICm1smzJNpSbktxlLiMANMB
9IY3yXpyfMhQ9R295f/lHvWu58mujt2plInMnmmgdO7jiBD84v8hwnFsCBpKYv+Y
LOulFFHN5EKkYoUDqC+chFHHPxfUJi2bBppS3eVrotZOXTeB4UN/JizJwo8xpy5E
zNqTxofjgbZ8MXqsp/svrcWsdJeBs2po8c+PefoQag5bdkFyz3fV/RgegYb0Opwl
ilmMfLEyMsuhpnAHn+EU59q9ddB8JKEbAxvcShCrXaUE0hdPibNQcUlEvVRc33BC
ZCNqLs0N6PoHjIxqsriQf49EziT9l2KzTCG6f45u2cGx66cJnu6Mm380U5IGtjXP
d+In0vqK5X1JmZDGSkSSwVTQFeamwWyFW45RbYiywRURea2onsH3V0KVRoaErH8q
qAp42lhOV5613bMHYW6L6oy3nDk/ulUj3fNobZzOlAKcW34eTF4fjOol86x+vPLP
HMJWQvhWFYyFYU+wFMcySo0PKerON6PcNLE/3jF/AIQ0fLLtk7jxkl73HcTChqrK
N9hCtMxry0tX44JEUPDYnpgzoi1YzRZXZckoJH2pKNlh4+HXVdqnff2nUoaSF1TR
fjSb160W4YXlYVsgFYls51URQy6Z4VINnbU4f+4gsGhZE7dZYAC0nWpsT1l9mFI9
FXbWENjr5cuHXT93KQncMMYE43Jurine7y1rplO0Zr981ZuE8JabyMO6V66ZyvF4
DtwSc3sHJkgoCAOQ0UUEVfDD6ZOaV6DCTiAesYt/SbTmLLa3o6sxBlCK3iVWQd1V
1TNW2a/8CL4CHFfMx13qf95rVgk71M03dqwpSVRrQ3WfdAWsEeHWapc1Sxw6vbWH
9jcXCzH4A4CMTiutJ83sMyVEeZd5Hf0KDuwJJAnc40jro2ZnK91JWqiWWAP9M/aK
CSV1MvsmnGLblakFqSaTLZoI4eBPNqIwz3ZjViCfd0yyBaGqu77+V5PFPOz0rD0+
EprGcB0eMBw58+8nG5sIIb2m55XJ8Co1KoSV8FxnRBBicVAexcsgVFeitGqmj5Tv
xu14iRRMFfP9iymrSovuWcm+2xANVQKtmIsPqA/tHmjR//Xcrp/1LGMR/Y0F936F
jhDX8UaFqp3099G6gX/9E4Ozp79dojc86EBEtv/pKZ4UQxBFpCGRkDAgolWwDohG
rEnn4YWi39kD4N5f9LO0eNXLNFMVbaCGI0j9ZE+sgvqpPypTFECA8XpMEKkv9RNV
pEDegj3LEvcvn7gP+XVKe1uk/JRW3A3fMlpxPaJdmlN3A6EMJciNaZUAXKg00o1q
zYfhCr/2v3gummDCrMGvXqrp/nhmZ2YZOr5EbcZMleuAPG4PpTjtyiXYlPzTCwQp
2sS6BNCNRb/OgstpWiV/481k5l2kRZY6nCuwRIff3qw5HZB1z71mCV1DGlxBJcH0
cTxIX2nYUCLgi+GkVzpgDseKH2CqdJrMYQ5rdMxbiNZc1Z+Kcn8Z5FXpS6GHzXbX
I/hZMlE56lBlUcuiX2L/cOVoVii/lyiByXBmyF47C8Sf5+S/34kbrCFz7+L/sfrW
uzoJ0CYi1pDcF9Hs82X5bMIEWi6paFqYzUZXmnrK6SMUbWlmdf2/2ykAfJDbWuHW
RMDYpE4A/RlnqDvc3O/MQKnbSEYx3d7z4nj6NtlEaj2GtmuBZ6+uYqOEnU9t7bLs
pij2qCiidKiIhWhh2CxuKel6ahP5J/Dpbhazmx7W9X+MBg+kNMXb+ZEK7saNIB1z
HqMyFA9ZhGxfTBUxx3Uvu1/HcvF1U4zHUBue5OdztGmCg0I31g6ZaC0AP7E4m8Gy
IpsWVN5Jw5lwQmH/ZmjKu0Au1ua/KQ6OB0ATcUCKWVaDSdBciDkgdHO5hbEBmIyb
QNvZzGabcOrEeXoTCi5aO0d1HF49/osD0vmfnCnfwa7iBtzvE7FH1IQ15CZoOQqF
YTdZSnuE5rpcbrRkBW05iUwHth6OXozougcXGmTzdBoYsn4CeXlHD4Lk1LEJjuqu
vT112NQRIFAF5fmAEq8MLfhni6jLJ3+2jIE5HowGpCZUBaN6lgAtZAFNcOADNnn+
wUuro1PBkh93azxu1JWxguuAOH9AtU8ukyzzxFPTIOYQFS0YyPMSMhmQkLKAU/h7
MswpDaASWSXeq6v0a5Da5GLzkGdepMqJR9NzC3XogqZN9KFKuxHQL6NZZi0WZoa2
Ml5OPVuwauAa2Ndp2Z23enbF4MGCCHY3Bn2TNx2tRdSbWILd1wMRqHnN0zXhL3Ij
svyBrcchzyaekohGGrh9ERkd7mwy/WK560LedWzxxuRHV7fd9332AP+Lw0+fQXtS
NtbwcExJg1YdcRR5CFheKN6q33szVPrPOuSO90fDPla/UKQsu8y08SZD8U4/ZYw+
EPdRJNkWJ24ERhOz4KlV3RMkDFJ1DLiopkiY9qFQoW2QZIKhH2TyXE7SS3b/D/bX
98pkYdvG4DcaEpqSNZUgiMzUQ+rAtf+eGBjRfNUVbbOjP2jhnJNuZx/EbleHVpA3
PJOMnIbO1EnvelbeUw0yqFY9l9iats8AAubjkUf0XCWPRMmUEEk4zDDCcOJMQNUu
7Y1XzfT4HuyjNgCWfWIiZWAylhXMeLIodJOw9bMWX6aEfXI8KrbbmZCgulbUk2uz
Cyl9nSuapaW83CmtgAluYZH9vPJD+X3i5/T7pA13cYLcvhabW5W4sbi6r7+beISf
xS14wyqymmY9ipKN1dXLgQrT7ykBabDXmUpoAqimY5GzMrrnOC0BGta77bhWMFU0
P1F7jiBKBs2JyHKkNSNmJaa4IO7XN50e9gTKpnvG1qcTSNzR1YD61S7us+YaSIKn
z7icS/5o78f1o/8RM8y5LeihrN9mFgjSNPLcSpCua+JvtiHV43jpTFr/zgmpsWRJ
vaO4MTAcrsOfTfrrmnXxwBmbO1B9LUhXgPCjXz8N8RRaHEKk0aB0ZOGuxRTUz2Eg
B/LyTx06MXKzkIC4h6XXR5RlKAhv8tepwEPjzWTRTYREaUCBVagtIyT/f3M88e/8
ekrj7BBvGG/3MF2TWKP68WSOMl7wbDLWnOS2zKD60A8szM03CjdVSUbXuHVzWXHU
SOtGRBjmIeldbZgug7oFRzo9jBEs0TCD7T1OR0+JajeiceBi+aLpX8XAyfPyaq/7
Oh6U4xcflcaZVJ2UFCjCE4Z4iJxxd4SEy93/HiDasOcf4yWKvDAPekqRHZ1oogIw
Y3AeeyltKB82M3MVEUCDsHoEdjyoPbB/uI73vqwx+uj0MLiaBX8T+SDF78ePA34z
qQAA55C1rxfYs8KKbke15eJ/D3O/igxvFGSjnY32AbKbZC4z4MXJ8P3ejlvLVV2b
3II90JV9ohB/219on4DD+1h/EY/YEFl56joSQ19YTGu241ZVHp5YBZk51l0YJJoY
8vld7X2kqLndTGonGJ0jcooT7koKinUvhwXO7NmnPQhK4SAWCUoSOpceW3fN8oyj
gHefbD19a6NO8E3Dt2yZOxuGEa13lg/rhnRaMfrOGGtojuRxKlJE8KmAYJQFkk4C
Wm9MBaMpmeHFej2n2TyXpIhi+Cd9io0pfZtE2B3RRYmuXDB0cbjXY6G/mxtzqVez
DMAxRusG2VNnLUijQ6q6bsBXsWw5e9+KptmbBCdP1PetwLmhQMRsF6myWY4FPmog
e6+NKnuzzCTitJrVIo1HL+jDtgVqtXXuNO4FXWeDTj+eVI7nEaKc6e7zD5CBOn0k
3dcMQACuMJColsU6GaZ2Tth3a+rDVbjLOxkiljRRSld0BL0P9JTgvdUbaIssmdXZ
Wv2679Ak2m00D6v9RDL6foSfL7+QpUuHxUDp8EHUMwrBiFP+N5+CHU997NCSNe4z
stZH+eKGV4oKoUQ4Cwf4T01gUaM9KUokm8jBocW5D55gIq+7lAhP8ib4npssghXn
81t8URyBkg0ERldHj2DDpv3KyHIAFsHG92PZErTcxZYO1YoDLP/DaIgUwYPW/BFD
ZB51vXybWolkenwhiAmUIMHfMV0RPolYwpj3mhjdnSaHc6HTlBqvm1k3aOY4FJ1k
zmJzavxVP8rQMEhGYawSDveWEwKjMdn5oL45baliQPWLIzkQPdcdI5vfERitGdNw
RgPdbCO7OwQOJllHS20z/HbU27n2hPSFjhccsVhzY6/wkx6+q5Qe+l65G7t6i4v8
b62JNGRaCnkVuBFa+xWLdwzSXhSv3BBxFg1mbhd50+ON8eIgTeifWjPRjVDpNHmh
5TkN/zgbdH8ZDa90sDDqx7OIgCXGJD89hGyw0EnW9ejrYv9htANbfiyw9FN2uaio
XGLXXChVxF3mWd7HPqx7ZSImAE5qemTsvr76H5oE30jOV7Qm8tRvoWvv48mNtj7g
r/RKMZJ3Ltyeg2kZw9qT1xwBk7lR274JwjIvjusY3GQeBhEt9+IYvzXhrb52mhK+
b9yI57tIiPSJMaYZ41awcMn/nCP3UGNhKkBDULuTE868H5VdrFhGB8WgyMerhzI9
OMf7oA0Q+/s86MLVPG565gNWaTPJZySbBKHWYIDjpDzyjH2ghdpXbj6PkGFDZZe7
iBN3+aq9kh4C7hNgG67hX1EKqvtG1TKmnEIoPpSJXrRxuluIlkw9SP5PH2t6Q824
8TlvpP9svckvatkIlAVbixU1+nsW5/FOa12+rNH/y4oqf4gsJLITZIw6pcVBl1CP
A533EpZ6FjzmdTyp5tjaLOPiy0btvFm8aMZzAUlNHtraMaO22ApudkkuFDvwpRn1
kyNVZcv1Rx+yjNE/v/XjbtmoYp9N74p6gvaudOdAKKFt9tyTSC3KIj3lRn7Igb0M
1AmZZ4g2u7u12YJzQtzoA7KGjanDuDaI0WK8Rgbw8fu8UYkyy/mjAG3Psx+KYCt0
NWO65hV5BAM6g2OFZe9RfHNLmAe4VZjG8KUXmlD3s7a4+TzUcDc291gJpDQJFgHZ
gDDVYc+QUIgm1GG6GPx2yLkEbNwEiTKeJKogOHNKuufPhumkuqAcPLti8keMv0uZ
zORv4fv3WPBa6uJgho8yWYOgiPVSEJKl6deTJ3ZozVuZNqDGIgTZ0CwlzUui/IhA
ALktNsiWYuvlWSQyxi6MM25KIonxVXl3Cyzc76hDMqTZtd5EKC0c1fwnERAYZSuc
6g/dNMxg+OCehg4P19hWTW/e2H0Onq/Z9mhbH/gs6EmEjA4CMOUw+VSK7gVZZX6o
66MUshkMXOsEsq+ShiHdKk+1H8TI85AllKZdzT3rhqwOwGBTFakCRHz9komm2HFy
DFFpPjSj+UycoDCn9K1aoBF4pXHXzEyIhIu++gmLNxN6uYkiO5oaR9kHAmNUf3xr
NsfoylellrCEdFdAa7vIIVE+V4XhmgrkvFo84YI6JyHGSD4PxAAToJ/zCyC3xB1m
bwwgSo8oQuHug3zSxKgMQbsateEOHzrImsxr2jdTJnVqeg3y2sZr2jMRTl3wQ4ja
erWxJgnqZlLM+k5KiNZQAgXo//NUU6Y0Z7NGtcgvBrYq++BYX7fEaZVr9q9no5Rf
ZiHv4LGdazGjNa79VBKO768L/WDNDRTcYHXcbHKydHWxu8FK8EHbtj52zC6mqAmB
VBUcdUvDX1kcesM0crzfwEcqmTWz6q8QsIdwxin8o9lWYXhWLlnSYcEN5E7plS2J
BACN5xSnvyOop93EieRORGFbJJ1L6ZdhM/ThVaRNwtSmiv5Y7GQzEX7mUJQ/+bJG
PHRcyg0KY64pZAKIueq1LEpofyi2WzJVePYURS+wuflQo2AD3OvisNWU4oIHGg62
KkbRaVHT4zhZZD3jre/Cf98PmcSbXTNJMzbpHyk1migTwq9MD9cce4556PNCHDiL
RnJQPR0qHFlb7MnRmwwZ/+I4rzRTjkHx3rJ8+uFu3+2wj9tkIoQyt1W76xVi4lD+
bDHIXTLNWvRHNNXsb42ZKJe1ApR7szEDIWsYpJH93U3C2KE0Mbr5AAtjOcl+4xB3
ZaG25tVIsv8PEY+UQOwx0f7A9o8s+/MM2Of8gFlM5NqD8Isbypt6Z+UqKlXYJl/z
d9FYhWPMr6PvAdz+QKZLiKX0I4/qnjhHR/MoJoPHQNVama4zkYBmpTnhTv/SJJaa
kHaxJjPp5xYKT7/D25oCxvDBMQeZwWRgeFwXt4ADotzEsaCk4aBbOOFG79A5hVUB
ZQ6ZIl602N5zZiWMC/FtUbdsXadMdWn2brg4qN9dBbmGWXmjbXPE40W+Ei/z0zMV
q4MpX4P4fQPruGrJiBfJH7uqCmLhNHJjySRne7bRhgUNwVrcimNYSYdyrhInqNmz
sEoWXZrx4ofdG4MOUZ8l80gRheWfF7Ui1Sx4dxWX+QYYPAPRJCJ6Tfn4m3fru2qt
13OoG+AEG5izFhGh/cff5hPwknI+Qpi58jTfBR09xxJbcJRDlTMuPx5vSQM4+6SN
zNLuxSQMakrdiP19nKpO5W8PSxujuGijS5HFBQl7cAdJB/HhlHsciSckphtZcc5+
IvcIPCAQ6rx0pXYeoV20Mvm7FfsHzlv7Zmdn2VsirRVtoKTpSC7IJcFggWgAzLCO
l046l6meBuG69jLjtgXAuwJMBAmhJG1FtUAWnPjrit+UEnZeRGxB7ev+oCxvxgQh
YRkybcdVdD1BRPIKTHLIKEIfrMeu5fRfOwG6sZks9XKz5zzZ39pQ34+FSyXRerUC
Ll6FyhR6nO7kQ29oKWY/8srs5tzWqVON9Acoq+i6O0T8cYFg2C4gE3HZwZ9Saowh
6mVxPCXqNePkuKIgf5TQA4tqW+9232AGCitUsE98ooR3cqF9uQRrKFo6K9WkQ54N
VZ+u+x53G2EjrJoRCy8fTkIC1UtbKXpU7v7noPShWvvlpwauu4PCG+fjB7JbZKho
S25dt1+owyWesvd2Vrka+530lM7fPBopHsKS1juHw7tg4QcD74mYK8AKvCc13ZY4
RbOJ0M1sWNNyW6rl//TRGZBFHUrxF7B3jHBPa4pAJmUHnAYxnme0fKZnNqFxeNJB
yl/YiGw3LYb46kSNow7jMzesA++/BfcyNrQKQi66zNT3pNIPznCc3taB4XQzHOYb
C2sVCrCcgSww76arGc51m3lPusj3W1W3kos6Ekw4476J2zdnpMbcYiCmr+0QPxMD
tzNBeigq7Cl3IbXxsT6eGHGzITLyOPGf3M2oecjcwbfYm99xfdPi7vnVpRzBjUK5
qhSVxtcCvFOrxVd+J79ngZgy/X4h3pnxGwb7o4ndgrKBJ6nQl/G1R0+G2eKsgP9i
6E8sA1EsF68FcQqMsIERd/4EELEvpV8Z58kH5hIRs1mX85OYd5Fy/q/vgFlrT9Gk
u9F7KqBqF+4tdX31/R1C1Daa7ToUDYhjrRKXdEU0DpbZXOqVC7RmINFFGA2vLt8r
l/Mh8d6tVCR+UtCYjir2HowjxiVo9ot/FW+Obq733MeNN+NE2UbRKabqAMH88hrH
bwfANAujRw2cZ9CRpwce+ouUm2P1dGMHItvqFn20tu7XdGT40m4QqaXZeu0WdEnZ
+Bcix6UQuvGIGCWlYD4ONwdEU3j8TYu9eYoQ4hIMNIAS9CzJG2uKDo0f4Z9FFBhp
UhgRvTkC8Gs0O5u6ECHFhz/NfG/N9DZ1F2/HXdRL1wBlk0Yd6lAIcKCys7lkZ4AR
l5O3Xkalt05VVGQ8PTqOMI+eSabGou0/o6ISiCjXIrLvueN4D/fTxGR6TT5AktWM
UJGaTDhHzghXD727DiSbKyRi2pY0rpvAFm5E43KOy+B2o7YGXu3m3sTDpTIe+Sxy
+uib5eK1tbY+jW2Sui5jqrJUlt4Ap0sDAd/KiUBm5NsYZhiIFY/zfc13hfSyStEw
FfHagcEYvh05a9xTWfGIQjs/1zxPWDBdKa5SzFu+5vk13z3OgMtLxo9lqLupb88A
zzQy5Kxc7jxikQTZWPt4FlcS8emoT0RJY4LuscwxysDtImOiyge3Tqiri6jVDvGI
OWppJ24U0QJTtNtBec0OW217rT2hsVOLqwPtjRcnTNwYk/78NSbLRTYAErDJfliV
utgh+GZ8W22luDw3YWYB07jZfB0hg8XbvlMSc7JosGcDZMgl6Q8VBXuygptt/phL
lQC/3EJOiFe1t4AHmj6Xk35uXndIVnHmo4fIEj8CbNy884/1WMSJ3IDf7ET/hKia
B16AAg09ujR7IxoZOeFdR82V2vc8O6hppf/qt1+kUPq0KrqyJIQI6VX/B8zhuKt+
w3AaCfPMLdNDbb4na6Qd2FJv6dXhyntx8XnWFJUnvlAy5EATFwGWCwvPhGpsgyjt
Iseo134w1PUmgArcGH7Fs4F1Jek7UML4EIDSI5f4drvVHr5S9yrTRS69asiOLHvp
yR45mdtGerfRPiQg4KfepmtT8TwKUSDQ4MgnhHNWJrVOC4DKUYYgI5Q5/Ku98on6
krhdlqzLe2dCshm904P9CNzM5bTtmsSOjbSWtdjiyPxj9uIETnQoOppoLK/Dh188
wf0WGsdaVCewA89Q6g8KlUmR9RcC3+73lJuOTJiEcJ8c0BAre5+6EJhNu7p0HAKR
TySRMXzFw28L1aIoRkAGZBbK1N4QdkG5e3DBfyy19OWvt0hXWURmvgryMK2tns0G
q5cXUzayma9kTu9L7dQ/+Bz9X3RSQW9aR048GBfmnFw4AdpQP6OETxhxHg71hjgl
A4WCUeh51MNdvT+BLCfldpyK+nEFFaRpjCBwThs2FeyvqYYHcjR9Ark7+k8hNhM/
uHl0tN/KlitfZjcRPtWrDCJDMAw+MNKfI8rdsStwm3MYuHxmq6BORDOcXkUgZNWO
60tYpYyEucBqq59myj60tGY2ps8JzuNRm/g8MihOn8P7eFD5c7cXDIyUx0+uTaCo
sLT3OTo008yx+YtCo0oh2jBEwYBEuBNFoO20tC9I9cQry64PcSy4jXaVpah/gJWN
AzDh4UavKlyxvaBsGoGuiYYWcGtudyVvbuVLIRlBTMjTPItn2h5r2LVra7LtgxmN
wxR2jWSynSkxQfN9oQyrwgh4xLGiRmcst0xjy5jOOfJiIzrVyzpl+OwHIuIcPqPP
79mPpULtXu3BGwpNbTXXIejFJh0jYo7i6HRRA5J6z/k67ihiuKxJgrCeQrf9xRSi
DTRWKQvHZpby2e+bZjuAT8RKetc5Io6m5MeSHWwZqo2c025FXaCoEInQK1lAkvxH
/nldeR48sdQPR9MX3D0pooYKctxRdZcCdkRkkfuLoobST8bZBn2ils2fdOxvDjnC
hKtheQLleEC0R6ShyQRbOT5KbjoKe9lRI0AJx7SHGgOr9hTaYQelumCrWLe7xcfX
pg8rY4xYx0flenS5bEMuaRIvbC7isNaHcsXKy4ZEQsz9rqCVfr0Q+htLGD/lIfPN
wHVx45cPXce3OKX/xIMpcwRzMtDVzWPtv2u5LK17BropDW0UdRp14elaoF37lcGT
/tTGBReIvtIq1u8+/1141winWfRDRwlXM1A0d/Ix3hIWM+rlkNcAEhp0rtYvnU/m
dgP6GFaSYjj4Iwcy0hyqO9TizGEooU2LvGUl5vev4fqET+6a3ziDsMBgZiFIy0u7
iX1JuSZ7sL7g/otIHI3FQG/3ovDUa5t97o5fMyf+uk645c8DYVbQsTDIeZuDiVJ0
itxcbBhnf0hCv0xVVhzAHDu2wxJ55slaSWgMXz7MyGdUt/ioSAAc23VXkbZJyT6s
GNkYY75EjEsWVF9+LrgmNj9EDOSnWCUMpGehGMADkngJ799F1Sc55ffJg8l6HXDv
D+E0I00je8vBZsPy2XzBmaCbmoMWLgjXHbuEs5yb42Verv71OkFd/HLKe/Z9RdYg
SeZs2ZsvikATGZFl+UVZdN29P7dx9cICt8t5YWetnbZJqMtNnMYemknDazMTnvo+
czV7nAuHVcnCBh/Wj5E2mPSEi3vYXJ/hgA2IcK0S+QUXRNafybZeeGjFvIbAjs8L
nFRDGUf2fJNGiWfi06uiA+RKCAbf+TpRVE4kPELFzSfVvG+tWVQJXUoD9hHriV7+
JCUGoaF+RCc57/+A9IrNpMkUL77niQj3K8brJnO0gJyEHSug5EYeMUyB7H8on/fR
uP/sUc7JXwtELtLZSKmj57DV2P/lQV0Jtfc4P6eu+CO8jasq+Hqq1UaTASVOAAoJ
7Djb8u+6w08hTI8LACs9uvK1saIjej/9yTHSTs6+KZbz2lxtNrslPenrxQKgaoww
jV9zbuh8O0bRzFx3KsR4P24eDpmeJ2OQ2z9ot+Qw0snq8K/hkNqMYL/TEe72kzCR
QtXGpSnkiiZP3Czm590g8toIcXSyCDSoYVr3Bre4fQ4P2oLCWkdEwVgCmsP+k8kp
LUNi4rVqsrlS8xbfaHTZxnvr8FzkLF0CA+Gh+j7WFG1z5L0r8PMt02vi+sbBrBte
pXazd3j17+pdKUqMPODpQCXmodfFjDCbkN/Gj8BUrX5r1i9Y+Rdjfk8ipXtele2C
BzvrqGV2XPcROv3czvo/1Opa+zf33M7DFQNATwQ88DBByv1rNlwK5/YrI1ZWPZG7
7B37j5AOP6OzVBSa5AzbsotHPnHVvg6EHZYlhXqivClncpIWl/bhTfveRWI67I7I
IEurHF2Uk6BRm5hqpKXhVj7Ru69a2FVG+JNUE380pcsbXrZO0V4FWJ2BYGvn5OtM
PQKrOuQGUaR854GRZHJflwlOocEfDbntYmIrmLFhMDReg1AojJ7hP9rZr6gnAhbY
HRCjo5tOzrxSVscm/pmLzNo9hp2iL8b+k65bKGBCULOcaYkzrPGA19MpZgyCQbc5
S+qBEPulUqnO4uQxNEzaXUTvoj55iydwTW8SSkKI9QJaurciEoGluLpYzulYlgYs
Xho3FrUANXHkg5IKjJ4fnkjJakkb1JkfEc/m0HKKvW4jT4tELSCy1dcJUlabvS0K
DAZlyio49JNhuMYYbwDWI0CKBekP4GvO5P6MYlCE1MD22yLvcuNXWeVR6znZ6NbC
FqRB+N5jx+g9DWqt2YvMUvGiBqhQkBWffdmVlI70fHRgcd4TAvL+Xzzfc4vcI3Hm
UMimeVCvhCx+IFJGxG1+hjd6GE1fj6IRNqXFlaQ3HDIWCPUEaXHyECRRCSM9ddtJ
YGHtuIfn5mDBrwg+XNnMV3ttTjMn114LQ4MFp0wK3qtRc83nYoq7d8j6OV+Mi+u+
o3xD2UdprW49Xl9i8OHFqNtKy04RUTmGYEQdepDtWnWVNctp3eHHGZRQFHREMi3h
+72q/slFm+MQ/6XHMXNvPpNeDRzL64bg2t7Xl6Dad55AmaBvyPe8O/XgJdew538I
AeqqayIskqmaWTMCmMErtep3cfCbZEaWrIk7pmiIfzMJ5Y0+Ws1G2apbCFQ7XMCD
k/mhmBdgosYWHk26ENrm+Xfl9FA/Diy6aawJgRNumgRAhVYphGqlHpdlIf0Jh0vJ
PZkxz4F7UXdHUlNkXxQbqcdlhGGEpYQRRq+BuRhribKb+cpbVuhkApBY6XlzYdA4
xuE1HkVuP28mZsSljyn/6S8ffQXQkd4KKeod+TiMTPgbUdJkxz8NRlxngAuYkKVd
DzfLX7qQ3H1sN9GhKKEuYCQAqqFVwb0FE+UjPdOGqGPyPF5kJadkL47o3i3Ucu/a
rMddYb69MRtwYU8QJHClx47/cBi1VZ76mS8X+sbNaU7sKSNJRvLSllUzvvhR7pBL
L10+4cCL9FgF33Vv37E5PteqfAy9eIzr3n3qJenAk+5bhGr9EnqZH0Q/oxI91llj
raKITAC4Z8p20ggEzsn2sbmhjv81hIl4jM1XQZy1O4tjso6rr7xPKL8dYBvyGqZo
CyX4FTWm05uvk8tTCwgxJbex6fxGrMKGnU1srKII9yUGsqOEBHa+yNpqxUcrawA8
fvTcNYMmGFJ+FgwkHRPWvbOebJspyqG9XOUw7PM7Lad4avsHtO99KIMrh1XZZcPB
s9bxDcwdQSqTP/yTGuOXAXKXjvQa8pIlpjY+9IO65XspOJHad7Vye59M+/N7EzoL
uszD2RhIMP0nxte8NKxjf3on8mMEzcGrqomIhRcbgVqHypvTpQ7U3pfs1cuE/CZI
HvyheVbAf/FOuItnMja8pBcKk4/n7kjIevE93NC6wrqdAqk0Y3ECi/Pwt8B59Oot
EFhWt1lxpuUGR/AWe/kTJZLcyOT6SU30HebcSqdMdr3TZw9WNG6jk/W5Qn/vXDjH
dAM97SQYtPwxEdFT5Q9fLh1ekRF+6Xar8Y5Rpx3JYx0HdLROQJYwjFjqLYHXxYDZ
9i4rRGVLSBMufacbmjtrgQav+WAHHw9Q91lAEHplHBUwz/LHWIwrLOjZB+9iFGdm
QqhZyqyutaYQly+Ym7eI7ySmhhnNadeKVUWOgja7rBRPsD5euMTlilXytAiuXNdy
Y7D2raHWJefMKQsNZPIbXnj9o97blLRx/MUS2V6Ll0D6OVz1E9isazcNtT7a269P
8UOFFJNWWwXxNVocPPS3mYWHi3Il3wIRLC8ziotVqoUsoB8bfBbMAoVnor0Gb5c9
yTwiVD5WC2QxD70Fi5RKtJsW0KdnHhphDYZIxH/aiyMY2c5Jvp4xGLQIm4ZRiOgC
quU7TbTtN7tMbBjNQdudITPOvpLak364Y9NJkn9KVGNwQZCgbp5mk3eMZ032mAXc
OEnHg//1qaorrGe/HeFLBkZt8UF7p/yXaY8wcczNuri/bcupHhMoBgS43J4JlppQ
91MjRnrWuxWDgXDWdnDIyUjgNT2+cPiA2DtHPlg0IVJlRiKzAAi9vRyDrjGXs/cU
XObaLSz1hOoof5phC4worC8jF+sgZypBTErnAkAZra6oFm1VQExHAfPfOpVSu207
QRDiw5jJhmmNr/4RSTlDUCKeQVznddTh7z/Y7QA8IG3zThhN3Zq+J7I9tVoBWwSx
+BFZywESa97UyJKiaY5if+BtpTbINycGEgKcR0HvewLS+JBTn1D2du0J0Kxculb/
IWHAbTN3nSlmupqJSdSOKk+kTd4aD4byzVDO27/csg1sZgKlWzCzj8gORaDhxFNk
hxLfq+vDoTYx+xPNCTMo5giFpHpUvMcBF2UoxVaseXI2MR5Juuw35cVamAt65hLU
0eZ163BvLRPrKWEYWd0Nc7BEw2PnfTMZSqtUFm/PI/ziWivkas+UFo/CnAnaCwWn
lO4TWZJDYS1G1X4iJ3aNm+qoSxY5mV+GpkJGiNDyuSId7OCJOu1sXNOsCrETuR8Q
eAsAkiUhJF+2AQ0gpQ2MRY+FVabhCo5G5Ubz6x9A6or41qYg+hcuvKt0fESCipWK
WnT9JTTV0KVR4F/7teqJoZrJCyeNxaOVdSMLbZiqaFCTKkDgdNFpQJcChMC/OtLA
gPKAhZMl+QgNDd94Y9kY69kv5OpSebt19xkG7IWU9Vu6Z0rH8v1akfFuo2iefohW
mW56+EaV90Zm5JI6DNpOrdpVyTQoQ/lQGOJTZ2WHN2HD2Z6xzYZoDLwkiKcGTS6J
Fo4KmI3CCc2DkfzmA3Bf+0sFMVMVX/T0kOdckARgWXrvU//CreT4suci/gadSqOC
71PiTEfYv+NoYftcS3eBrXPr4baJqO7POTadTgMV9I8nDPeGc+PET2Dv71AWUGcn
wTMUJs5YK3rVlLWROua5IbTFIbxmJQ3i8CxCKn9BCtYzM7H5xvAjYxxBosMshYxc
rUrtlJN7EHfWWVnauzp4Y5U6VGFFRtzBWSVf7nzSHK93YxFq1PnY46KgrK7bFFnk
LPtVKxgzRZabvT3hrYmhDr0h5AGCm57pR/zrjPT8yRC9kfzeAINf6b3PP/sYi5kZ
xC35qTQj1lumGakifz8Fjt38k3ghRA2EN3RFeZTSSCK4PfhzkRhgx8S4WVv0WX4Q
3XaBN030UT2rFFoM/5CcGzT6HGqa9Lk1s+/UGsUWjbBnUNDKG89WCIrcpssfCW4P
0mD1Z1RRsraM9ciij1Mh+RosGgWyKjcqGlrUjzetNSfR/CseVnjWwiOVdPgefM9P
y+jZD2wpTiV0gjbeiwgiA3lJZHwImJL+pv4mGQJrr9R73V7rweOW67cN3F7YJS/7
AnBq34v+l3cTyyJhQVdfYJv8aKzduP3++R3pgT/+5fRE/ZSu7EF340sJdfSLwPwO
zpLaEFgMwHzs7P63YN54Xq81jkOvc6e1DLsEmYi+vwGEu0kwsXP+hZiArBJmRoFw
JnN5uQDehPPMA68lR8Jl8rUVTGXZGX8pW7/CIwNabEDLhaS3SNwgzMhkKIf6c6c9
bZDsZwAoGZ1nDMxJBWk2aWHZ7nAcBWwv6Rt9v3jN1jaugHw9B2KTIO+Nrp2Jvt2v
OXD3X9LPqauDlCH8G2uoyw1aJxKpfT/DRRshfRpWl/F26bYZaKz27NgbvnjWc6CD
X1YejRy1ORMOY06kAdTyt9kVliZm9pd6n5K83q+BZuRagJyFuHi9RscdqbFSaj6O
uuiAoEgIGnxR+PxisxJzQ3TX8gkK2YwbyYpl/1yC38+PFO5x3hj/LJVqd49WB811
KLHF/gfnk8ZzErxb2rNz6ajzOAmy7nIbuV+FNA8oVjq+dSEl2w4gFUY7ehgfFEy0
qxfFsPPV2fe6+ptGKl0FaEqs1xzpSCTMboO/OQi/L6W/SCDjyrolWEqooe5KICJd
rs0MeQiVEPqGuoEAnH6+9w9zwRY8w7uwCsF9l1rLYzmVaL8/U2HW2WT01ucq0A65
rQF0HMlr8voqzIegNY4Xa98lXybpxXLwxBi0jZZQbYNkpHGOUzqVJHFsMbFpOsZS
iozi6KSH2jSABvHqcoPpxgTjvGLHLFRA9Sa5EuahYRNRktrkBXtvUNOFFtCtMC4y
xv7JPHQw8gz+XE+Lsg8hM55N5U2YF53CV7TL14ReoOwB88JfMHS+JYM4KkTDxVGs
r74GUQpUXBa08LDynQa1Wa7mC+xl8/MaKPUCHnU4aRep3trgWW7dznrcG4bt/SzM
4equmW2hfTe0Y8w9o7E7/r9qvwpN7//DUpBOsnZubEr2mU00XoPTWVUh3dXukSGN
DkALyfPjHfggTnlyUcDE2+WQNypNCjNqXxDGnPu8IF3fOpzetuo7qEdpSglAE5b3
gL/mVoqavXYVkRACM+FQa7jFOWh+3r4SDKkDtDq2yDSMmaxigS4cyYJdzpcyfNN+
nnbpssB0MBRj0WuNUMl4tPOij8QeAa5OdTWObOYMjsJ2Xx8UaZIzT7DWD81yr/8C
CmS2HjUfLDQwkKGP1WYuAsm/Yb4FZQFEhCBIkIl4vXVujy21tWXHtJHt2w9CygdT
brNkwSCX23of7WEMhwnV6Kj0qRGqv52mWz1gUW0O/dE1WqrfkCO9dl96IfhiMN34
er8aw/m8pUn+or6zYQH+THNsBmVVav2IXICvWcgXYjbgaw+B9FErYejc2qsMcFGq
GRd2IxJc9u4X7Mn3lvwwpMAdSSB7nIJuprwVVKX9he5pU9T9cKexk5h2Blit8Bm+
svJS+lYJ3Zy264BXdudSUIJ4XPiNL9jhIClGOoh0Q3+YY2VJMbt7LlN/f0QnQS0L
GV/Ccq6cRLUurAD5ldoawyQsw95LYf13VJ/l5fdwPrwSeeFBtqT8Qm9tf6GuLwmG
61P9ghOhVFyU5ZtHSan5/NcYZ4xrORiYx8S+vQf973I/ZebQVwUxr2G/HSObHZcw
cXVQR88A/jCViHAdft7wgB/HoiJXs6f+xwmRyHKrN3T26+R4cVMQs5WT3tE4GHhu
47ID5ACOZtUgVoUouoi1Nzt2gNAbYHwJhKvBTXgJaD80bgDa2VXsORake8SH9HE4
SDiq7BrAnnitiKaYzAxzp3dRYq66WH+/ro2OnzfCw5yLA92G5DW3CpDE2UdWCZcs
WKQ+j0LtXsgOY+fK/brlA8TIw6NBn+6PwW/KJ8zPwznMLeRoD4PulKpIXdP0f/nc
2VNO2wB6t6y2RShVhZS7QVGPWBEfIUvizvC4VqkshPX6Qh0uHx0G8ZC5+geFfovI
JKn2nBc23hbtfev+dyKBZidY48mPFDqBe+WGkOT78mht+WvEPlSZ5fzg82i9s+RN
pPsb6LrA6jeSAHV766TEbuxz89tTGNl3iEO92ny6zmHXKo0gxW1uVH6VHa9V4MTJ
6s3pJYAq/aHfuIzFGc+M1vFRidtOM/yag7uiVQ549JGeHIAySxtVKUWqjiSka7Ra
8monf2WKo3YuB9F1IzWlkmALIZ6jUKex4Xh5LhVgIpGdNt+m5IcZB8jy9fMC2Mcr
`pragma protect end_protected
