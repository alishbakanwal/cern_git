// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:05:38 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
MOg25mqkmM3vId90aNHi6UJJ0FYh9juwewOyulpcdzWJKBnVy3zsFLwlHyAgyMpm
m1jfxnGZAHFmiGMHCQKK8pSqGnUsIkrdcyv5TKaiIFaqrN9T1S7oRogBHlvqWszD
TEtXH7KrAgki9jA7OWuWDJ+CjS+LdGv29FuvrePW6ks=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 43696)
U0keFKiJ8e8kl0Yqz3IBHbucMrpd47LneAZwq5RCE8vOsceF+VU7C0dCv0DERWRT
Vx8RgiPqUEsEZastMnu30VVNRS1Oqui+mRxnxB/oKfp67IC+GQFT0TF7hwUXiFJA
bde7LdWwNKIww6EyYZEvtZwfqlIlfIqpsE/qjU0/RcEQvs62a/qumSHdkL0zXgDD
2DOYS/Y0p2N+7JbNBt1vJFYNwXERl9E9orX23ZmZajKogXOKxjh8oKtteYHMa2Qj
F3rOv/FYiKYzSfMuqCOCyK0wYL2IZrn13laQs5t1ItIrXnqy4GN46x+ceyQf/2LI
xyZRg1fZLh38+U9Phok6qG4gLqW8IYhlmi8MpHD4R7WW6JdOvDxYN7xnKyy7OfJ8
cwKOCMXEa7ieGsfuJ0tUjz2M5gzznBvBy1M3raXkkDGnwaOT0p7fpSEO5nu6L0ld
8NW4glsAVgUayYaMPJ8ndICpbqvaLInYj541VqvLbIs+HNtivPaj7BD72kVRatps
83Pzw7Z9MYHlUOeLU2DKbrXY18WPVzGaxFQOIgjnHsTxciAQgJp3esHPBJ3n6jLH
nSfQ67yXuO2UfPbcFTZiCWgxOjkHYP92+ME/k3Aim9IBL6fkh9pUBOW7RLt80Jcf
EZN1lFMWVKt+v9L+7D/9nRYJFwNHJ3yyJUgMHbqf9ZBIjrbroFvkpmBycqhlgoYz
fijvA0yLxpSE3zKe29OV8srUVGe2re7AkU1R2ZkGEm2Gr08sV+RhbiTmQJRvteIh
dXM8Vd49sTorJdLX12Sqf2mf+FP5CvXQqZdwllGapNGZXNXGrYSVC6q4smGK28MF
L3a3EFir3hdKdHqZd/So0876slLkANicWLRa/GHbgpi85oaqDYSS8ELM7lQQUhDo
UJs+r0JcCU8gIoW2Ow8f5V+7CbSQeFgB4XE84he1MvJ4+Acx7WQzZQSRtl280pxj
+vLNIAv0ZgLavlKJOHJnn/1EM9m0OALhsP2ixbGvGUTdsQtA61IEwgognskNxkW5
hDdQnQip9vSuDFQ5W2u0In7UzuLfsg1EmaUDNeqwyGxov1lfVXrFrY24+lRLJpjx
oFlrODg1C8kcdh0n/43Gc/vP0pODXobX2B8vBJrh1oGV074eAZ6pUX06zq4xyl9t
IF1wr7MFMD4wpLIkQ9sIFU/kqiF9YAf4UhbQB1eHJbttV3PPwFa4HP1gfDj+f7d0
NHUouJllxs8zK6YiVySUqg3h3kQ14G8cpCQvpP9S7aKLPHi80xdMvja56d/3KbSk
WTKcB8Zxi2x5R4m7msnKg8E+kctpQVijSqgLIoaE/nURGd2/lZXsQpOlMepMEtGq
lV0k9FcMJgu2u9ZzXAaWCRGiJwomwy/sXi31lK5bFVo0vNNBQgs2CG4zSvqSajyS
d4eQOVe7tAtYoDOYP2qfFTR/bxcM9njpDf2Om7iyZJL3OI3gZ4+MMA9ZeIz7G3yb
xkkqsvhml2pDWSET83wdouMN7tLuTC4e2mw09zYGcUZeLEETEgvzyXxrdTVsThwG
NqgK4KEWJj7B9VePkmdIrJn/286ajouCwfsc3MnUJPQ8xDj0eHNIfkplDKa4Z/dl
X+miwarqWkAAgQ3G1qv2LXTEs7uOh0q2USUt6DiURJfOiqHaVFnnK1OkQj9JBpc9
Lcm9E3t5pyrcxIT3elPUtJafqzBmhjDscWhFyK2y2FD8bWRDkaSqcg7iAscRBSYk
sfKQVmY9Zq2nJaEyZHxFapxJRUCgdcSAo6SNlZ180jBjTutJTGQHypr5HKB0jdTf
U0kb2sUiC5JWn1oHyyc5x3bD11zXo8ytxK7BdtigV7MlY4vmB+57B22eHWZdSu25
pzVnElfyiI2GaRO+SE3rN6nrK7Bf/V07muJ1Z6TWRuW+puU5onVF2EwY2CA6RALv
kvvFYElUQaaL2BKeeQWXteCIAl5JvZKgubEolSJAxilO+XYTBtce+tXMbvvd3gnt
tRwv+P7V+NejVNwHX+jgIzMdxwrqytT9VK0An/RM0p5ycWsJHjn8cKoRJzk1cIQR
2BkuaNk3XTjp+LB7uegYS2mVGN2mwA4UjhquUJ8ZZaHrqufUl6FYP3rKoqLuqAsx
vJKjGfjY0IpDJpOgHWqwBFsoFXfENmgDVOYmR6nf4odODwDWFxpBrBJC1AIaZdAz
ZNo170Pc5k9Wo+2VxQtC5M7/nPXynmNlPVg79TaiZBZlX/jK9ZAxSPRGN/fyXg6D
Vjz7PzevaIUsEz911Vdu6hjiyL/GOhelCc4kyHpFwGxKSLwgVHG9lqzIpkSxzgSK
ehKU1p2C9j9tQCzl6ppukWGWo0pioWVPUh+e63RPHMIxnjVOwFFuW6A5y0QhHvWX
SKh4o7zMbm4gOEF2+1666CLOPzYWlTK+j3IQEjBYWOFSE76gVn6dElmlXH+G+J0i
R4bkWTbsFtqn6JZyt8y6Jh/6SrmN8PJJfhXolbt1Qa8ZsRrOFmLyvDUNPKk51ZYl
JGH4MrotTHNIxDIn2VOmSNFHNOWnsUhOX2ah+mrN4K9Z3TNUvy4d3pKLNJe5X0R+
T/FEf1MdXFek6/4MjO5KI5OHz083WS4je6/WyD7DvIIClzRCkOtlQiH4JNEekg23
kjMoBGSjJpKirsO8trk2Dn21NYSGFFctydeypyHMu/r0scYmMlIJbbtROOhYgLIb
REgRtuRvcVCW087ucM6cnwLfROT2PqxOdHVcO8FcgWVal/UqXkOm6pUuY2X120OJ
U7/gR2zF4sk2XRyoTFx6tfsDw5ejoaFYJOLHjLKAQnWfLoOXUJtfvzjNrR2slH2X
6NH1B53u8u2xox/xGHWPchz+I80rDCSyGIxWq57zg2YIAH+k/XOCe3FYCo7zsTQe
6PdvhyxpaleUNHInUC4L4J3dBalP/17d1Q9fAItOuCH9zS2DJENZiT/U7wtvhOVF
ciashCrryjdbt2He2s+v8XNSp6dMQbXwCmGdpeqMLC7f5rDBLxYh54RM49TwDBp4
S5tfkrB7LQuCrMvZ+g20R6KKOAjhY2c3h0JedN4bBbkqZCR5hlIAtc45JsJV3fvY
QifMH1z9X+MbktRV5Kn9HUmdu27pJ6nztMHa/xREuT2Yj6J9O+J12E1xJrNNItoG
CYhL/GDjI57n0i155EgpVOWEYDv/px0qTHZTRWCAY0PBPg0uXVVKvIf1BavXIX31
/au7h2suS2QlR3K5v5za3XMltm+iPZDyNG2SCKI5ZqyFimSZWQP1N9JHtEC1ZYv+
yIRXZScgRPvS04ZegxIVKWRUfpvQvbn0BzdjS/LjM9DRzEKCUAS34QFvru8aFjTS
vQjDa+YcMdmGZyRsxVFE9WronWwK0RH2f3zXhhN+N42aLOfvCvPkElhIaiw4ZYRw
a7qWXIm/Fv8WUH8/+w05DEa1YTim6fUHiMv+641N+YK9fEzzjB7J5XYRu6uxJWjy
75QALf0Ug/cwA2qvaPd8gGM7LDoOIhbxLdxErG3F3BHrr5fJcsqV90TsWznRifTW
IOaHfhNvjN+1VS5Zh2Gu7XaJAvfprnl7kSxlll9IAd/dnp2ZuGbT84b8RIatKifB
woq+3mjaDWBR0zdZR8FN09XiO7C0APz7sUqEe5bjbhwPfIRShYrZc4IYwgIrr8pf
CN+kE6DEXC3WBK28KSOF46ncpGyZv/ta0jqMNgqpf+KZ3gyu1ffOuRp9Z+J96QRq
ePwgftfa20MbRZAEZALnEGGOT4MIIDPk6PfGFj3LeC4ewIq5U1QxIvZMSDpgUxXJ
0pKe01kRTgJgDtS+PzbzJtOEwRzp+xJm7/pCZif2FXmjs9np8Y0WQGU/K8FcdDyH
KyOEexTzrvVxsG0adOohorXHhnS3vatvJQUyB17oEN88jGiP9WrTM1D/s4xiCEh0
sdhly2RLK7bBqUN7fhEkB4cv0Ttbuts1zJN6V05iq8dlZx+ccDJ0MVi2/36ojA4a
P8/SVdzC+JtGZNQ/g7+YFO9XX1WKX2yx2Ed5YOHs/ZiXBSIaXg4cWM+kfhZIwVM1
A2h+X3vmvQbQyOo0CrHVlyfDQLMhKdzfQqud2Di5CKBmMl5XsmyY4x5197/wq+19
qIES9scwwFzJYZT6XV/1fp+dHR4F/AwDLXh4Za7HIfup5Zio3NPFsGtksySvOEd6
4l2UJ5jSmFyLZoso3/IYuUE9P1pc9LEaEpXnm0IbxzAqmdjNZvrlDqH9kSmLRbgC
FZF4K5tFr6UXTSM4Qd8hG4jqVcN5dtse7PTzoVUBDg1NDA/ndWBj+jNDQg651OJq
xUwJ9/riscmgmHUi1/9Q/etArt2bSoaE+vtg5aMAoOKe7Ubt7Ep7oD4i5WQji3c5
aN3maA4Hi09FtLTqH6ktkz9OeByY0zLRaD2t8tfwP0uwtEbVW0XDmxkNzCx4Yzof
1+PzWJKKYUBkdZmYqEQ6SjxigkafjrH3fOCRtuOidKytb+aL36+/7pGvx4GjyPCp
Q9yJOT/AzLBaqfKVEHpkv5DWyenxEOb7fGZOyidzLkPajLga3SkpjyHFhIdTl8tL
4JxlS32ZCgKcbJESZr9LoFnexqcPrpzyjadrzixJOwxLRXblJ3FalI4bxK414Q/d
Yy+la0TG86KVGtSb/Y4MrMxqY/PKCMKeXwVxcwvnN9BhXQiCkTB5XKagwB+x8M/E
VhKhgqFxt3xOnzTI5n8t6kLEq4tnhz1Cvfw/X3lUvWouLSlxqwqFXeYJlINRG2u2
1YprhTCXajsZcoJmwBAzMbI8BTWOcDV+8L3XbcIizpbpVM7xswBFO9qdCWrwA4CY
sGGLqQOQnMwOdcOXs8s5qnw6YtN5PHUmeMqCdMXxAWNZkeq++q568MX29kQOK+fU
ti4095dlqS8iH1XeidTZiMvWlD2mC52eGLiYk9uDF3S5QBOUfUDl023FuuiLF3xX
zb/TWqKs6pNcftTJbrAAZ31FczeIGZRi01rcdc3ETV/wtaB5VtsSayukib87mGCe
UBW+tCLZIBFdxzyKWp5JKuoaKupsHQFDaSC0f8yo/R++wR0wuESKWUi7D0aWdCDL
1+mCsBH3JazwcWiIuiH7UkkiyEQ3b1pCx4ExVYspOODeBShO7yk4FfqlT4DlynKD
5Mlq6fqRiuNA923j43ihxbFMGeFaHnJLe4o1BpgKvBALbz5vAoOYV+mzkn7+IChZ
3oA1ayUD+wmk0+UQdOJRynbXNiGt9WPBZMmG/bmhUc/O+nXcKQLzN/Gd31MbEM4X
VePQueZO+9p2a+8vlL7yHZAAt9WwdkZMvAH+KLWbPn1fVacLpNQFZ3hddnJF9513
eErl5S3H26f2gr+VP/pzWBeqfFc95xwdo2V6XLDyoNlDDN5OaR7knqv2yi4QCxlK
Rm6lXyzTiIgjSFwNpTnnPaUxt4up4HQLS5jzFCAUdl+CEUZkryvu4fUU/Q9ucJtU
KPMfH08L7TT1WiF+WSf7G3iyNFElM3zetLaQRsYgg91ElTFxW9Brvp1uRqp+efSX
VcMfrICJ0wfDptBbc3hhSffXRnQGiIPqfVUbCr8esRjwJ6L2Ngis9HFpujgJk0n5
9AyCu5YEc8PKL9r4dB0tSP2mF6U1x4xsCCZ6ZWDEnLNDf9x+5E/6OdRVqYifBHQ9
LrFEcvCeoVCtDog9MKE3KJ+9Wwp//c1bwM8d+aoKM+wi8VgaZ+TCR8O7qHi653uN
2CpNqDGPV55lYWLzaeOsO3xxUagFtSQKPV0bxFtmSgJK5ycYaR4GYLkjrJ1MuGm6
KOG5Wem5JkjB2bSQdajuXAVSrn0ED/JxyTZG3se8yDtG6t4Y0TXCs/pru9OOhBd7
OMo7BNZqPc9Jfj0sy75q/D5c7qYa+Ocf1Fq0cOBh5tXoVnliu4q64ZOkvZojUkoJ
Y0S9yCGqD9YvCg06nXiYYiHfgYwuuK0vm5R7L+YmDXZBBo+ywVmRQeBTTAycOr28
1iCaquIdYAeuaQmhWFi2k2gLIeOxliciGrWNMfl39VJwlvygVbRQ/esdlh+nbkD8
PU2M6YUql1jRmt+QZCMN48/El8N3+wQL7PJALUd8bIrg7JuDSO9sQsmnhvU6sXBK
x3+wahGBhq92z+uZqzGdQIOhHhyXEYc7jHGuIbGQVDUH00VLPo1tBZVEkyH0DUcN
0pVNiim2WQvd9luhhu6zzGQ/mfYUkjO0CqvBgzGZb/VqDyZ7k6T1tdjLGt5QHcFh
ixwPtLlYP2dxxOnKnM1AjmNurdtxUIDYpDr1Wq0bngbK/rrZmbaU7dGafiX/iEJb
16oNx4CJSuPNBQadtq8AdVj3jfUoYgxFprygx+C3n/ObKg4dwtb3Qa3CR0Vh5IW8
c1ZOHJ8RMk84cLI6+aqvh6G+RLTTnbh7h9V7jojblFAYwz4MGWJ4YnXnfttp2fZG
sPVqIVi8p2Cm7lvi48yiRaNGPTqdXMFZY0Ptcxvffgi6QJW8zQZI27KDxpdZRc2C
Po1KEYly407zkYubReEOIikKLJn1s8RBs9wn8Fqae0yc0dleOLPOvKjrahSiC4A6
stbAp9QBfgwZ+DS+b50FmygJ1abV15Z1gEiXYtavetVsnCb9mOG4SBswCVI3eQk6
+V0BllICNyM4VxEdbMcC/k7T4ixW3jPCfK8ahhsSBFdt+c7bJt2fZBYbzvqYlilQ
8Ck1VBIac/AtVkO7L/vWzbRfd/E2+K7fcRRjDKhqAYL0zuWharvKT37s8sYzNFbK
vA3Rqzpot+iRRhVlAYKkSqLedwYQcuRuDsPrXth0st1OZdgTxGtcwIVVoT8Lq0j8
X1n2ujbftLF29IHjVOw/0t5/JoLpHv3LysK35w1PFIu9Yrj2E4t0QtbOSIUo5rH2
KA+gp3zK8XeY94rUPWuaklnkqOFhOQJOVhld+5voaUSurz/MjkYRKpNtLQeUrGrN
NcYqDBWBIEBHbee0Oy0VSrhFI+7l3J/5NeU7vUBQr9LRNJpZsTWi/GpCPc2DdSPW
p0JX+k/3u92UG0V3LRoZYYDUNXdMk3FiF0AiaAUkAbO/WcSYXaeoVCqUBYh6HDI/
elcUokhMWQs7iEahKXZguSjGpzNCb02/P7riqKBMqjVucVEAV+rtOmH2S3Fwn/sT
6CU7stnxt7JRGKvzA/18T1wR1MedVrFwGczr63/DZ5dlD9g0OmEmgJT9k4bjQdps
ZwdcJZsx7cm1iY1mxvI1WVtL0zyKV/wivdVu5InxVpfXzUiKtc4MV6YQIXkA/LK4
w5CsvSOJEX/aWTRtjWs+fadAh3vfYmC0A+5w6cinQoLr0TPuDxnMbXvk45AmeOLs
4bCTrJ9hUQ6rZQ4tNVpFACMJHo7FdAtkmf4CQiNuElYKWZGWpz0hLuiLn6Rmaz5g
qAD4KYsiLcRQ61GTZELt20Lp/zQVeAAbhm/fV8RAZ6VB//0tjDxCzGSDYmPOZGa0
krua2S0BC4jD+qDsEXaFQKEgWRqZ/+RiINm69lQYKeYG17JdfZ5/lABj0kThmYn0
48aLkyUu0XcI7k8aVJUjP4y+pn7I8JvnOJtqkepbQAed2zZBPrXLYVuVYFAxX2CN
P/vrniMB9o8ljJzocWTll0L+GxK5Q831Xf9XpsfyqO9ZXINWx6bZpqh1SQrJIRK4
D00oKmt6LsNCuUUHMmCV7CUrYhGNLtT0oqlBwjrY7h9rgaox8N/vp0v4tDYURDR0
hQIxbtvpb+hWzRhFTYX1u5z0yNOhzwrdJvswRLesJmlRE7DPHaQVTrtnchFx3SBL
P5/3qMwf5ZEU26lAsc9rjX4jcBYn7mkjkOY/tJAeKlXthrxB9dS4hQK+b2ylcbds
gw+ZjL69q475bjRGQjEYsRPhiHktuasEnIRAanrFinPz8eXuSyNhKf04oweS9cc7
Vdx/uT++NMFmKM5bCRV33ppXeAis0EO9sgSkcUUp8g8Ql9nX8FtHjiaqz0rmn81B
n+/pvT3IUpcz4LigYS/9cKZExzNnn9MIyGTyBrSjTTyPvQ/e3yns06mDBC8ICUnr
uIHsxeQMr+0KP8dPqV0W+VzCs+4ZnxNj7+tilzBflVjDOQkbaVxqYi1Hrzg8Zv73
qaYFuePXt8MHIpw9sNMfiyZ1sYuoDLczado1nmKWwIZ8vsZgRyRzTCOm06vqN6xN
Mwz49h4cARS6G3yI5/0yEsySL/cykGphNxST20YuM9Jlt3BJllGmRSqp+ArL93gc
BlGPh1ZQzR+EF8P0b18zVr2sBy1MKMnYdRKHLOv8Hfi+pp/rPoky3iW2hew7HkYG
SSzneo1qSNUX+WFn/WLO3YHKclTJv0C3yOWCRKZBkKe4B+sLAeGslHjE4o46hxdv
ZICBx/HZ10WNXQSuZzZqRT1clLUBKPEZKawY0oM7soZAGVgiH/QREymmpyqs2VPx
+2IzJC42i+/2CezICjHI/UVx7wL4m6xAhTyyE7u59zJ2snIBxcW8KvY/9SWiItyf
7YbVA4TlZzQ4cMr5dqwDfe8V0dFjrH/rpYU9TfGsWQzQa3SEjbQ6yGH6gigsGX5n
RVIA7io7zO/Y05NetSX5j8eUtbMykucyxjVOtAZvBwEHN45vkQEN33iJ8d68Jc4B
Me1+kSEO5K8BNvIHsQZtwlTFPn6KWWQO3YHzFBXdjae+bYvjEFoktU2FlA5p52jA
mL2066nCgHZsphE0KPauSQEAFrVaRaxtzsMk44At3Hkn4dC5MwynhGgAbTIFXs/w
ftbVRWgHnzzk6jPShUI0xBpwda/82SgsgHmfwKAU1utfuhxPbYtde+eD3y9lekzd
/PJ8WGj2wXqE8lE5b8QVubfkIub37KViT13f3ojqdDVPJyeHV5B4wKKtYe9HZVnb
EzkPWdoEm6r9j7gIM1Pu/WnF4YQcLLbdOx8BAI2NfZCiLfmi7OUYzodjaPZW1PSH
q3tiFREuySGQECeXrzMXDCLN1m3SSPuoUtByjEHxgwWqqfyLWLcXgaE8kS19LoWN
a/0grwe+lSqhvoVVXuiMLTJoXDxbiuQ6ka/qnP2o9oxOUUcb70Ltc9137szpmxY5
Y3kpnT53jrNhW3Q623PlHWyt0RcfCh2UsDJ1YE88VM4dK1DdPU1Qhyzv3MIMfTwK
oL5T5hBs8YgsFOnE1OMCodPpSxGMqQrXB03JXMCBsHvEevgpDHtHT93CAQji+10G
THIgkR5wgwX2UboIBk9873oH9ZKDg/43SnyxP3+PXa0Gboe5C5K9Ls3SORUpUkLT
QdzPGi4+wtLAfnFJbRNQhUDwD+hQ35Hb/7alivhFo1u2fqrDTFw3RyViIbPlIg7v
rGLTHSn6vhyUGC89tktzynujM0ibyVBRZZblQEJRLvHKcoxkfx8vt/euWNUyEohp
hOaFKp6+vVsvmJu+B4TJHGBJPYfsUo26mMKL/NfrWhcFXnRPY60fPbRjha5/oPGk
YqPoFh82HDiBQl/3gaNLj5NI33LMg9As6tU9EXxz0K3kU6likuR+VDTmiGD3dW8v
OLjBZQC9T8fMrhmf8tkdJYi8BZW5OU0lyOjy1k+TRPFniOzHRSv69AJF/DX/B/Xb
2xiIna1LO0x2DJNYP3tLh4bhXw4AjeDhleg7A+R2quHaIkcMYsxFcO83/Zu02kus
P5xPPzhN27gtuvhjcM+GEx5LXgkiUSwy6oQNuCqPccbpMPR2F7oTAjeL99X0hUQc
JT9iW0joCAkAj0c75Rp+MDT8FBOHVEFhd52XypYtfHtxdtY/psj/dQ2PPaYFiQ5a
WxXyg7dFMCdCsA25NitUArkAoBNhhVdomv+MxzSVSRP+7K7LzwsayxpaHoI7tFcB
j/mYWH/14lKOAWvdqwL+P/XYE793MgYceufO8qEu16oxM3Emx0RIieZVHdHAbRPJ
wLyig1GHeAPaNSadfsecuOzPhVAsG8E2PMm6vW9CYIxDMVtECEupRgChwxvYGPKP
vEcHeu6TeeLw0yO0Rlelpco5Z1qD4MZ+sdj0rWz2EpA2JWCSc7lyOY5Rh5GnIqoV
F6r+fakpq9nI80eLrnXGQteomoG93lYtXxJHWjXhEXirAt9AUyPiyMffSq1iWYt4
c7yY3762lm5XyPXDoMlz9tPI3vg/uE8tWQM5H5lHZNKr9Un/u1fJp4w7Nsvg1WKt
2Xr9BJ51a7mFpgI5Kq7zFE1wd1hrh9aEYHHnnKcSoOPFRvF8JeaEI4Cc1b4gpzAt
fH6ddQEkkqSKpu1KocZiIZelCL4cjOCVtEPwBq4hVWtFkLWSYC0CBFbFMOzFpuJ1
s6IlSLy2gBz5xkylUeXOumbSkU1fdYQnHq+yPwNLLOYtD1GlYkZDa2nBMs8vPlJk
K12RU/Ik5t5DcVSljQANXHzhnuM930KputIUjPHcaFfOR3OvGtfK3RCoqNbDhwOl
bz2joL87qAHcTJsikJiLsUNlixlhq23cjMSWT49BMTUPa1iaFfyxX/XRMFSlsrFs
s3yONSNn4+KAgP9prSWrQbEAwiaqs7OOvZ5DsgMpetnE9VGevO3IrDqNeLTsNYBw
gE5PVfr4fcSR5K0tLEProS0aazNZfWr3hc7YHVKtYjGwQREFgfMjEKt0WBRnLfJe
vzbFt8eqcp2Qwx/QotRaY9YOKQJdKduq6v3jdepac9zYrwn29c5LOEO8Hu89C+/F
85cRImc/lxdji6Vjc9Nfb0QUs/XK21ZFWw6AX0vRbztqGxX4VKTGOXpRAM6LLNob
js7T8l99ZriK6716JreogPSUfkK6/n6TvGLgCsMcGhIVylrK3U9zmyUU3fAIyLtM
mBrrlSp5gTIyKgzRLsj0Xvoo5apJfCmzXqFCCvjAiR+YjOJ+RPQMyRt3RUbFt7aS
HGNYyCtn+C7VD8y6bo8hmyfl6dP0pwTbGCJ5tEsotNOeAnqqVA5+o8gcqDeLwaME
E6QD0BtWGZYNIzxgpRDnRoE+8mBXyKVvhVsQYEdkzkwWswBTtgekvovStcwDftJE
vX3rM4BmNjA/kr7MCDDoPDH8RoGSFxWCb5T6BNf6L0zwYtE9GZ3PfIloDs7T7WT+
1kL6IQ3guO/VgwMpG4+naA7ie3QjJb8b561qg5SC4Jd0KEWYiPH9CZ9ucKrBQp0L
mMvoIDPlfDLwoeR5edm5xO0Xv6TIt6mpvf9a8Yh87YI29Yq6T9R54SChuk3nerYG
j+/LWvBt+mi1+MUVICJdDWC+IUCo9J9/aDlacBie8qrTXWvupSVbyohf80zGvqBP
W/MnVTOqlJrZlh+XmOTc71v2L8QukHjHpeU6pV2STKKl/qKT22F5lXEgKQ2rH1LX
oRsF1pMfIAdUN/9z68ybhl3Je23t/YlSFHTjia4XjpKwkBEPDJFH62+RELzEQNJQ
q9D9owPAktsvIYGw9rd9U/Mz36HGvFk7qY3GimwwbLgvaWcKbbw7Te0tvx7hN10d
8j9YhIDAlNDP9tRJskvAkbZXLqCpkXPmfXxBOg3m/zaGabZQ9AFJgNZzk9dAUKrb
Tvp22ILFtUKghRxD9BpQ9MFgw13ahqJcnC7XzxP+rPaiqdrmp7LJAs9SOnBBvEbo
Osg2CQwv0bMllIhxe85eAWuqZ8ByTenfO3b+v5q3MPq+AZlA6niBPJvSJ0XfWbRR
+xH2kXSRkxop2Ahb2UQKqs9w4BWZ6so9sSoY/I19zvRoUdviYGVskGmH/3boBfDi
VKAqAlB+/B0FESFFsSd9CKhz7ts4cuzZvvdMvKWTpf2PQvMZy9FNzolntsGX9V5f
BQxQuWoojsOx0Zw1EWoNOXpvUxblDSd5HZOa2GFUknNF1vyWNQo2RxmYy7cBJKWB
GEjb1Z2wLoYlHNTh/kZHDeGsL0bQ6OljHxBGFNPa/q5KA/jYa5vh+k1DM9XO7MfI
7404EtXPwIxUsIw4ErWmgt3VhJTYi1mSa9rths62Na/JEMsESma1UPvOtNAPmGks
0sZ55hN9rgz5gioHqbKu+zqicH6BSXppsw8XJKQi5tXwRaQ3jUjvX9IIZzPtKflI
/nbr2i6+DpjXHUfdRgSK6wwLFd1+EMS+Zp5ey1zYDhYsXs0+9gDlHpSu7n5NAV0W
QEElFeD3BYMcHQAhf9tHZkkyLVHxKoaFvNXaSACFziD877e4Kw6gFFye6XKpqNU1
CcY8S6Y6/PJFjx0eFb8AZBnMR2CdFBBxweC/U+mRV4rk/fsyk5vE6BmXvJ2fTr8z
hnW/mNwxxXwB0LAQw9kSRoD0c/yFKiDr85rSkuxKKmgP8YvXszbPQlK7tyZDkYsp
twcUcbora9gVWuUMx4rKbzj10IxM/eWu652/tEXELczEkd+LY2BXodTvhT8BERVI
9qBFeWM8BAN49oWullQ2igB46ImJSJXXJmLXMtbiReR/k7T/tysEOmb3qum1zNqW
usUBIJQnUwfp5tm6W6Qxq61zWVeCsinboP215T+VtLBqGtvJEN8aZkAmAM3V0xLE
CYCBtZUHym05uZOeg/SEYVplLaxNL5OuDHEyMftxsuySkqIHxmu14+ObONYSYV67
qwU2RwJc0a0CzrAgx96KXHy4I9QaKocrtqc7JEanQjkwOFsjc68Cikg/Et90dte4
ETabtqIgrfgI0XkQpz1ml6xSC8hCI7EDX/sQ79bEW+eIIuvrJ/jozGc6NfbJ0+PX
yPwNLSbBPdzkaM8T1VEoYwLovgX9wOb4RVfAMvi99lIxMy7I2L/5L5Vwk+Ta+/71
tf+nkpdFgRiejFj2u/qw4xluHE1pXdx+y/03pmAOr+fkq+acYy43S6ff7LPJDYgZ
SZN2UkCVaVKcdH1v1M9qEAh/zHVNhq4GJ6b1mR2RKZlhzYZWeHVU/i4sCnRvOolw
Kl8h6tgugWRDXkyhoSxehle25g4Z6MQPil52vXvNBIFPD3DnwlTjhCXVIvbX1ViA
s8dljVlXjHqh13M4tV3aU/RdJTqBdOOIfXe1RCmnjOtDmyzVJUaG93skqTOhviLZ
vOQDhyoEVPiPO8i27zHEIip3X1VNHYM+zmM93RBzbgkpMgEXMsqJfPO1+Fb4eoC9
aWdeVKm4Y2lPErsFhtAUo4HvWdXfsweDhDRCNHqs9roAQn5y9ul1tOx8zcPQmqy/
Jo8OcrE9D4YYAtYpt/wI18f++Ctqiei9R9hsN8v/3O4nl4efjcN2Ew+dPjaqocPP
fjMrSVpVARCDZ19ukSoE2CL5rOPErV4esNm4DHWXSDLLyvF7L8Fo3A/I9V6gtjtq
Kml22/0J9t+sE1hpJX2d0aoWwBQdZ7lvhMjHbD/a0iVXw8/d2pC1cvvpgtXksNGz
y87GsngAwUTO50Od3jEkrN1mKP8xICQ7IbKNNNEVAOCRvKS1Pw49iIomLqwvQ/Qf
UWo3hbW4DDTOXfgbcKLScyReXHokSt7vB++MUGwMYaHFYaituF1lWqsQGRPj7soy
zKHmUMdZzkxvDHxdUFX/7tlTljjfXpGel3IFwSMXR2RWlVQBH0hN0lLzY4BHYyuF
TdHMdEo322kdAm5pzLU+tzteB9yyIrtbQqsdDdfw7e6N66R/yidzOFKsnQGVUs1y
pyRizpcDohQD2LMHaOeF//R1w8mch+/nPc4ueeb7boeepgnG37mBuXHebpchfhmb
DlsE0g7mNFeHI4SjF697wzIoSK4oablFEdnEctBifovZ3XPZlWTpSqGis2GL74pw
AHFi6quCpfzgizxtMYkiraE7yNEi+xk4zl0qK5plqOCWx+1C3owtSJQRiyN/m9Yg
RFwtoc1D7WZaexRUgRYxJJv9xV3EfPR8WGZGpdq++/ija2BMLn3y2VxEcobRCUr0
x+/VsXQTAtMxYYy+W2/uBH9uRRJv0pebt5OUbzXhDfSLqXMZb1h//l3J0ieM4A6U
AGtUSyJNIy7LzaaUyiqs+iFv23ugI5IZwujLW3u1gnz/AKzDCTt6AKs3JnGTZN/P
hYKfJ4Irjr/sOeof4W7sfzLeuGgqOmPzR+8a49EC97yrIapsLl0Dr2lKShuH+gdf
HVUkf5DUBA0rsBsg1OgDcgHEgKcrXzQUd+GfyMqE1hFJfhHmJgn79WE3oEQgTLPu
L6yeqe49HbLopM4BROt6BJT+WsCxHwIBq3BmDcpKST0uZeA37iIcz9JQAkJJbXOD
5hJCxVg9c7AwGL7+KUJUGf+epNU8NjlBelLYJchxyKDzz1mG/d+fN74bDzqCJV8v
FTNo/WrO06yAcG1Zfg4e7LhM8lmPU7fLOl+VjVhmU9sTIIEvUFm42KLxF6NvLREA
DYm65QGxddPeiqBwkC4iqcfE30voJl0C5ZsH3V6XJ8T5yY/qTfv6EyZXFZrjDnPC
oOCurUjBw5wBa7orTCis9a5ZoMOBSJdgXVNrksjI41oQAocyYDCJLs1Rc6DqvU3q
8Q3wRIGN4ZM4iJgT8MXMr3bmsrrZ2KIUTW30b6QJ/T24kNIxI24CqmNfwPLPAX73
WwSEQXonPxKC7e44YCFfVDMhWeKq858M/9YN0ZBgAa2djr4x7H7O+WjxTMJAJd9I
AE3IUR5A2sZewOokn38XGiGgJ0PnqdFKkBbFm3H5BzfEZxXTHwKQ8neNr7Z96ZPV
uFnSAMAlJD53nF3wmSzzkazIvp2rLVTs9Egu3I5uFo8+EgPmaoeApZOqR3i6zNzk
CrKWDrIKA5Yvn9C+7h0IJBBoQeeTLUNnbp348d7ca1k0u+z6dXmebhljr6x0Ia85
mgwYbffsP3i7+b2nMaCt4D+jtjiyouN/qJwuKd+iQXXMQk57sviVKQT2plZ8sYf2
ncAcTckWJR/aYPbMcHGG83RkN/OmkAmzC1WrUpkGIaput7rPdz7a0+NLH7Vt7LIF
7njUyzSuOhcufJ4WQMyRIQD02Bx8nBVKnFl7K6cW+7/q2vKettm1W5Qxpusvt7Xq
RYpquEgHWJfl4V0OoSQ5VzaJgRucLsTYMUrCKHUaZa5P6tJwnXoMYSpCjvL2mCBv
xMkTlfKOc8OLqzjMMSJeq0izbJAiwKEfmRwcFDuLOrPjamfPsgJUJMqHr9XtULi5
iRfh0KIWBkWocTPemjIMB1y6YNeQFv62/1Nutl+Prg8WT4yOJzshdnugfSsmpHOU
QBlgayw29rqr+ViSbaskS4HmqQpNzg+41ovMYYsE95BaTbeE1ApjYjwniA0+/ojT
J4UjRwcF8LiIFWSMnddGAdkayTXz4gbNjthUMpbI02KbPq17pYtKkNaOYebAomQQ
/yB3KgIUOiEHPCjy0aLB8dtUdx9teM96vd5LfICc5uin5/cyDfRHJoao52w3PXQQ
P3LVOIp8IZbVRYlvJwdgDSs2AMkM90vnrwe9N9xfDtj3NpsGNAJ1GKM3+N17fwWg
79/Ul1RqeS6BwNVi4FU3rdkvygYnU+7PO15Y84Y7CdK158u13bjI8nuZ9gxVwdUT
EoT8uFXBxp30S0NG9vMohhenAtKjt5/Kox7s0wC+cfbv2RB+QiiiUaX2+I29MwZc
GFmSTbGBcxUmI0XL8t484tHNFpDmnFUoousAkL2cWBDM/9LXOwFFwHXlSShAFv7C
/bwLYlKVpvb2OvczUOR3Ko4+9KaOgTIB2CdChLUCf96vCdBGPK401RiJr29VJSIK
fwf+Kmi8SOCHyLgrskP9QgvAUmIOI2fEO9kJ1rxA3X/BwdRgrSiEDC3jvOQh5veI
gLnvWuY/usuUBz/WreTFkj05eUV5z+ZFI8Me1A5L2IgwmCKjafWWOwz700rqITRt
0sZpuXlul5YVgbU3Q6jTrCfMfeoX04NUfo+4iPbtL0egi7PhSh/Er0stTej4ij+H
dwqaIbtrfwJfQkZXMIbydsZKbz+a23dioeeKQuNJLqy1FCJ7qGeFizQaFLoqEp/S
5Ji23zVbBpohaSZfC3rOoo6EAlJsz55MHsUcy/NBjawC1jqOgPi3475l5z8nwGPI
2/qsyOvZz45N2P3451/x/0jgZv7/L+TXvINW8ApwTnSOtoZpNf585+OQ1wMsR9FD
OKL0vFB+V6Ul8RlPhEK/7nqd9IhOSAQ5nZmV9f+KsjEOiLgXuK/3NundsRkv3X52
CDslOzI0ewcplp33CKZN1wS0g4ZX2DugaJpU2XnNqGhCDnFK+ShC717wIHiGG9P1
7K34AVQURRUrzap6g7ON2sovmdDmXw4beOYdaojqeUHEJ77gEiCONA3zwVt6yta+
Z1xj60ZLb2hApaqEatmknCIIebzinwjKGrNSMLwp9yypyCYZXGqotdm9dIUIZeib
C+CtED5LIHL5Rw726UcZ/iyxAucvbhSBPojv6+GiDiOzYHCHOeuA97qbT/Gwnvfs
h3sTY6oox9vS//0ra0F+esHYLNcNntpHjFtQ/dkyawyNNEWyMIwMYzy32iNTHAxX
mHS2aOff2sUN1ll3nCXHOXKSnEUrb/utdY5lGQyYrIBTaYxZZPzbrPeC2zr5fuqr
hvOcP6aiGkkURy1R9vfrYJHbEXmfV3zattxDrIh8c85ub108CtcWqzI1dDMvVkBB
gnJDTlnpV1OC+PGmyDdJ6FXuueIOAYPwNWQe2rnWQapZ4VJbGAmu85JuZOg6bLoL
xxqYpyMygHkWW98sAPurr+XdUTx9eheUUVSWPzxtzLtutpR6Mi1ADwrrLZOANVGT
7Kne8+ympcnylt8NgvfPWP7+B73a7fKRVYKa/EGDb9aEszg0B7OGa6hFriFCwLnt
zNBfjcGrKLnhrn8Ey3hEC+Rv9UelgXiUMTvaLR5WoiDLOZeus5m6zqh6hNG5jef/
Yqei60xcs66DghzyEpE0a2m1mhZXvLd6F7bQtfXs87h+tDejXSnRWHJmUH5GyOz5
vScT4iVR1usTcA6b5q0tLp5D8AcNdzZlTQXylwHoloxykbmhQHW4J5vgDZzLX3+y
fKg2s4nLONu6U5qKmvZvGvhO5/mbcgT2bOKssS2LCCotpkzSGENnHHpBwda3Ewlf
5kwGqs1vIYJUB6fz65fs1uXCiIyBD321hdwgwC0wbPPjfF9OOAEt/QV7Do0JcgjV
Ruvt6EMZoy5IoJw9FjjjwmqqPdP+WLQh7l9bOXP/y/Snxl3YYh/zMwwpARZguNNA
Ir6g+Hu+ervWGiQVifpIgnp+SWzVnab66/iN8UolAt2W5hmu/xukXGkmI8DKJMZf
lNJKYhISXdVfHMI0vUdO1Sus1siOwSziQoz6U7JYQoyZ81GGVq3+bdR9kMwV19E0
wtsg1VFDbxV8IPc2kQ1OQEMVbGxl68knEwuhvi3O8OCCuhAKmxiZqHVKdfgeMPLb
6m65cOiVGj7uA5DBo2bewxFe7EmrmrNLxJzjr1Ob/oJxK7vkbakuHw10eL5rJSzT
jh3f+jZUWGvkXCMpzxAQgXM5vwr2DvLpbgOo6M/99FmzE0tPYSyhXw/X7eKZpE2Y
EjQqEELJI71sFWCwE2cqBKIN63scijZ/WuvGWgdKXuP8uEOJRdHOiLbJFgTNbpbN
GUbhzLcD0KPr8Ttn6CBR1qr8eOjCI0950me0RXWdOICeTnT+oNqM1T+V2cJBMQb9
78ruOzVbSbr2lzURW4s7xCDQuIt0t9wHIwjihRkWAHEgUxrDGBdHjKlJGK+MBtt5
AkMARtWhaM1KQkx4gAd/h9lHH9JQC92pbti1IDzJ6RRgklusST/7pFPovhq4s0k8
LRXXVrPhPsypc+qO35NU/lZw+it861A7dOBIZzAxFZGjsKLEoU/zLT0dOR2liJ8r
xpC+fkwkTwtLKegPTrYWh+ZChp/2cQWuE9hg/CO57IEmqKdmw1ypb3e6uIZXkcec
bAN2WXacq4gPJrAmIBpeXLDSTJhGgPs6EQ4TuIpfMoelwKPWIYFGDSGyP0wxttu9
83J9hc4FPjGjaz3OnplqGQ1OKrLgpH3VFr76NqMGo0NiIwTxvD5VNDxg97IpzoEi
rJzGWtc+Z5gUMbFDgabSDlkPlGLr6OgKF8JTFnMQBiJujjnRYep5+qBQSc5MuqUi
W9RQ82ICzbx42CnxyjovopbiyZwVXv+iyE1KsFE+9EYO1J3ILseOd3Gk3IWe9AKE
QyLGNYTnUJEjR98GfoGarzOT2rnRp4bODnbZ1DyIcig06+nHZUDnc46UiTu8z187
XMVyfb3D4KnTa4NPEEX+oH5vQAlVOqmyN+eFnzkTKZs8vMpXSRd6WBV1NS2kD84h
jEuI8NP0vcA2AbbC+9bf0fAFeAL5bN+sCV0sz/9bK1NiF5zWOTHlnlBUmckhv7g3
rVTzD/i2W1lF15xCCkKucinoED6tdrNXXhyHhyS1tnbMH+S4T/IUriWZ1botfvJa
wsHdYtgY9q7JgEnCLe7F/a3760inZaFZ7R3rf7O+WW2XNPvyXqCRxR7+y+Dn93x6
54qKRc8eRyBA0HcgVecgYHY2UBJ1+92BNmn67Pzss/nY1kxD5k+gx77cwnq/Y+VL
5U1rKNFVHAA5Azb9nC09MZwipS67ZRTNEEnhz5ZGafhkx8nzM8DkI+/GteyFmS2b
IsGGIswY9DcJBcSYAPrXQJ0BlStGXOKYf3jQVoZcirH6pGEXBJyWjCDU93av0C2F
NRW8yUd4YvMi5z4zsEqkk46NpOn3HWEkqKVa7rk7wOpr5YKjquP1DrjZ6//5A92T
9MQ6uwWaBkHgUsAsvf0FcjT3Rp2CnJmtS2Oul6FvbJjnz0TIizbJeoMGHIFFZeuz
SPN6buhpLvKvgzcW7cWLcCkTwNo4H3eZ1dvoMtWmF+uIthBzuBHk/8tatdp80cCh
RsEbvnsRys0RZzT4IqtxzXPwTRwlqcFw7mFAf3bDXPre6ByyGlF8DESmBr3cqJJQ
1TT5XUQ0+2hsepG4nxUFG/BLojsFOjEkRujpIFQ4nLPfVJxQ0cbRfu7eXrVKDSN+
XKQ4pQfVcSJNVqueFccQprt+cIBRNjDBh/VJeJa2dKVR1+X10N7/dbDRFnfrnLxh
nhpZs1cU0+RreUMdxyP/hc7MSgQ3KJhbC8I8JUf8sC2lG7pCTORb+3p/yLIfKNg4
FXmu+BDs+xXY82ZfutZNiZbQv2ofv87CsgDZuINJ3rLgWnQD5eAdS+Bqm2J6iXpK
lswPdkIdL0oRlZiQHL5aaeDbUzC+Sp5CGBAhtI86yrfqiNjmlwCqeSI9J/pi/4FM
UYhyeTr4gcvZoxpZWbFqIGmkJoHePk69yDUYKA++8qNB53K31T4W7vUXWvvjGULP
ZkDykF+TUKeJ0Iy+n4+rG8g6cirS8C8azcxK++38BNQc/zWdyPNqF7yfDng2mLcA
Ju0aT5kyXGPXSazVIjxUxNS+Ul0TE76tDzoOJNHo78jUvX1zJwA2s4FsXRrsR0Jz
OPtevM896UK4cjpf4echXb70UvfUeEUHemGvvtEcy9Jy6xU7yDItCIPta717iQPL
nXNcvrkqXRl7ftjGydb5X0Edagm8Yrks3azujD0VGGxnQUyGpVoVuf0/3tfrUY4E
pBVks6yy2bTVOe2D2jRZNesBfPsBafh588CzNkJjFWc81bW0xcoD5oLngJs69rBF
Lg0uO502330t6AR+WqJHVQOBhdjvUSySUlzV7cckOeoargCISvT+kc6XPTrvwI6j
uHSKXez1NYC6CGIZNOftcv8T+p4ZtXsKe+eFpNya7hyUrGoVDRvIqbFOYlSCBM0n
knOMj3hfRef/9KdAsdxWktyWRHOV++8FVdN+6tK+CddP+eNbaCKSm8NIYC8U3ZUc
r0ppm5jhjcc6kI4aEyZrLhjblhR8HvUJfZo+WzED9+v6VjM4c60YBTk0f4Qzu5FU
BHjLyv2ncjkTb7PhUnPbhna/T0vOLp+WcWwI5Z0ElZiHP8ONoWCBVrXKC+iQRxu5
PVOiojNO57gW7AwOWx1I5t9AxVGsW6hOd98mFV9X8FIi7JwWn953OpaeU8GvQ8dj
5ZqKb/vr4QwpHQ6zhQ892IqkDx5hjDsGLAX00K7O7OzUN7PHKecUMJvK8Uerr9TN
wdg3nAqTXMEHa+SMn13LiAfym7HnAs7GOla57a5Vnz0b85CrhkOj5k8o2IKGTJsy
HD2sgH/aHsVfKtfWzwc+LSO7CGbVUoSMFPuTdDqNwW5ixSGmOlDMPSws1GGdPycr
PwQ3Aa7TkAtIFhhp7kE5LCUJ2f3+WONOaru4iRcncoEq9ZS4sh/GA0llC1rNp221
RCjCIkhGULIq6hyO83NVpA/AWhZrJYGoGc0V3gQj9c+x+kOo9wBDR8QfsgDEwYdP
g7UQ+T86xY5TPTixUrF88EC37Uc5jQbblGckWg9LsEZmnt8ktCkknRb/1OK/B+gK
zTAUGZp2ivp3ubcnUI8NKBbpBDdBeTb1O7QDBFSAC/GZ7uq/9KMaxuBTaK5fnqlz
cFtpv+SRin9OICDafiTqmK+FxflQTW0cER7elpqJOka2PjGpjYiWi/qyEvVW8Cc6
4DtDQ/ZclPYPxYfw199FdstanFHCVNOjAuD2sszdRShW8oHwtILIYZHumvGCcsTv
FhDJ6BHeDFvG9owR8Y0o1+2IOt4PxVvKiVX4J9m90ZtcVVMctYZ8XyzPPfPmUqHO
Nd2EbUjoKkLXyNCyyjXxRu5CCHOnGAJnCGyUhD2vrwt7o8nBqaHnGnGT58nsqoCM
0x9kYYvLJT+G/K1KB5gFemJVbJQd1MgrP6xH1dMzyLZs9YSIeXAyIm+CgTGZepCV
YdxKonuA6oyJx01PdPvOBCkrHHN1LZfc7DXFfHUhzzHRZIW2arTHujnKV35XTqED
vIlylVvOAvE7wq3tYufWQGgbCZncHYklU0874ZAPdNOlRUBKMAT78UHQQjPFM04n
NXyENV3imfQ/inoPOJohD21YdQ4kWL1v8cj9Lg397lxucYdQopjf14rOq0Tg7O8H
HkDENy0ujND1OqSynKkwkSDrT0LvtxdLBFKE3tVfA560dUpZ+FEqvWnkx65SvQdo
KUky0SSlItI4DDV2nG3maACUwWX1EOdhjkpWlTB9J81TznSdd8dsfpb1zq6IwotI
ogj48Y8bTPZlGYQbYDm+4JQbLMz6DlhOHkSPFpS/NHQOqFt6CBr1FH6FZaT7b+LN
k5Iozg73sX+nArT4Ms0LEHLIb15Hotka61M5rGKSIo2p+oIVh4gM5d8hMCDRlVRd
F6y12/tPEzVGTDkgMDNUirzdD6cz/s0CXoy2uegsj9dzYfkIrDF5QBEXQzuUS3Rq
Cujbbb1Yk1UV+6rt8LoCsfquXwtMMXVPz9N21LUIwMWZDmxdSCdQOSdZgzNyLpk+
BBHXMTilDL+jCL6Ar6nj74MeUgnC5w4EvVL0vEyH1hMRaAZDCJpTmwRBVOMg7Les
RltEWUPCZYvRLCqU5/4+V0mvmcL2Rgwh2bP+/9TzSTbxQKGVY42Ba6lkvwQy6KZJ
pcOwLTvsjCm8I58vg76IX+aQbQ9PizYNSSWy6JeBOVfrEj2pBVkFiShaI/TknrXh
xu+BWRJkvT6upVPx121h9F6baiBnr0YfhaR2MzRchvMSX59vUj30bDohYVTDVq4j
AHIny6EkM7sBlvmRwmXugdEB4iGS7rPytS2ersWGQKWiKa1n9/TOBQNR+PVVbScS
LC91Pphdl6dGjoV3m1+xZEcKCrIOTaA/ry1Zwx2ASk6LIJpCABXxzqoZSrY59r/G
X4O8GMYPbQ/AkQehPgDF/bjA1CT4Mi/jWbzhM4qXs/9UAbqJHrWi4X/GLZv3ah06
ViVDQr8AAR61HG8Rv3ruY0I4boYrX6rJI4gUR5BpFgl9BqNWfvpYZUuX75f4ctRl
O94G6O2xLkSqjhYl5HlPJizEV3qqiwd2JKCp0HnnODm94sqkS5A2nGEujziKzl/Q
Hd9gb+RhMBMJwuK7+WCAGYcvuI0MRg1Qe8AlAMiBLQJp/b9AB7JYgZL6Y8I1LwMi
O5NUc2NDvOkhJWSMbjBV/xvmSTT22cmWZP1Cj3s+pbkCSanXfgzgxJXmMn/dKy5c
J3Zdd0MJ15e4Ft4zdocfktG3NXW4WeFgni/9NO/OKg3E62tYziFvG83vfhFKxYJ4
TQEuLbOru08oQ13wlM2vXVI3PnSAE77kIFyEqzM75nL2ZlHrG2tkZeYDeYs08xVK
FlScYYqH8aJJWnMEbLzhmeLfhGd2V37VMrM8R8LOJ5fVkF15emRSX56mfab3Te0V
k/AgcFWgOLWXYWSJJLDcQoOvXWztg96aylU3/nsHaHhhpQ6joPwuS8IukV1NUw0z
8xCrXTwUNGu+CdpObIkga1mwplluul3rxrOgeX80gjLW2IhkrfWbfyvYvLu0psg6
KfzH7LNRa4xfhLqqj4yw7S9Z4hqrLBKJTH8oeB3GhgE2aEaX4micor/rlIHfHjB3
BvYxys/DzfU1tcMbPinnWIY1pRBjAQh+OQaUEYJi5EksEjLbZ0tZsXRce9lZ4/Ji
9cXP0TQq8sisCpuXm8F1+Ufn5Utobv1Ccs2dszkUl8k4AqyWtE9drYSaU4bRCpkC
IX4KhzlXxpOmrCKWArBpzPfzV5I5E2PkJLNKuTAxklqtINZcICHj8A7kCNScrDiH
aIbJhLkaGnmNArFoqkiiK30a8+0xFtCfnVAmcQCMiP2jrm6vuh153s9keyiR6Wb0
LY54EzBEHFz8bEqW9M8C1jv4dZD1i4zIF3F/Yxivx8nUl7sxHZZj17J3OAvYyUmA
n8jr+RWfVRRJHH/maaxFOjMlGIZVBXxW7K1EE6wTeBw9nMAZSP/Bf3JXS7rj31Bn
D5R4hCb17zmOWyQ3gtJDia9LiLqBdHRRFS1Qk6L1TKnjKGz7RFxye71ZO5LC6lAq
mhn/rmnlpbRSyqBj2HtDYt8IssTlWhiV72dX8FxuekdQd6MDAvngnR/NZ3QvqxS/
W1LbXSb3G3ECVtnN1k0JG03e4umzKtX4/czbsgVHU9yj5NdWoUG4ok1fWb4Nb4O+
1q0iuwYCMIMjd/ZDVJGcLYqQJIJuVU17eDw56iJX13k5zhOKv/VmhCzUaESxm5EJ
muzQQU5i3+kpz4m6x9hITBBYjx1/muUZd829OJLI0aE3LsG9O6sEh+iZ65P3sVwF
4wISZf6wAbo7kQAOdyUilWwvQBt2xX5UFbH8ZkpAnM/7Ohoud89ORogDMSTyHxth
cHne1NHrtJEqwEZggkMF9w+iuLgvxLsPCdYFXN74G6VJkKC4EKt+ApIRdI7iMM63
dDsZFnvuTHMXdyd6nWOX3a2Y+SRR2pZU/8yFTUIB/cf516KPv1wNUG/lwm7wbozw
3G5iVlPBEUxmw82Y/qp02r7IiKFX+jQeLT43/hNp6zhckKMDTnQ2SVlmoPLUdZTG
eWB1Pkr6dsQRNR6LnFrfR50PeqbB1eUYCgKgD4MY7ZNr3NVRFDPQhmjU0DluHxZc
pK23f0XvgzelKPhZ8o6bmFLxww9HCfkduP+qhx6kYynaTA9/PUCa+rCwV4URQ1po
/Vk1DLah1fJq34IcQfSDROyTxubBpFAUDqy7eqsmgHV4wAy6uYfDYV+URqjRojpB
fqh/4N82xV9cICmOhRsBj90C/JbrLrrCjF24icDtMgqKz0beZiir9vH7/ZaYTlCY
+y3pyn8NYSGDFM3dNxLstODoQH17PIYAOVAgBm5oKUyGb91kW/vrRZ1mOhDwKt5c
ZhSv2EGVVLtM+FNchEjAMggY4eIdW2W5qQK46DEFVUx1mavUWuP9rw2hb4VikP74
qR1UZtdlM4/peQiEc38OUbpkzhf+zWwbmSsSm1cEPg/hwMa5AZGptzebyAjJWL/C
2K5g1eW2rrYaLt3w+HB3x9Ca4a250QNfWbCBqbdMmXx1ZM5jaW4AlPC99Y3oPMqy
Yr/kXBUVpgQd/WcaR3NcM/y4tTDn4q0+1yoK+4iROYIw1wOzpACdGmpuuoPF6e7B
T/zADkJ6Am3c4E2ceQpae83rUWYYM65ArBoUMhgXaUfNoRZWuKUnT8JwuVC9iTeB
lu8MYP6FBRaQDbebBDec8+V8IGdgwl5okDtzwbbdTgc8bAuk+HdDp4oNF4m5+9iq
cfig7J+VUfw4ebV2clp42UsJ9HsdGrJ1yIGD+RIB0ew0+9YNGbXIshDI3SZ72fz+
DsDgCtq9j6LvwEIN45OvAgLeaSh1uRZu/gyujnHbQL7r7+SjLrUQ5z4NNkX6UGBo
0MtBpgc8p4l6W4M7iN+u+3uZvSdLvNcLb+MCaroNjsbfrW6V1WjM3oAFhyZrjyV5
h6fFgUHJu9BU1YohZi6Lhpa6/RFtS3spRyjMQX/n6D0vWZayC7wq4gdZLOmj07sk
pqhfTwyVcgU+L+2qs62dJia4nreoKvtFtU24QEaGzUTZItzIt7jzM3I/9fd8D/SO
iWZ8cF8RYGoumZxWimLrHsEc9HHPkiakD1I1Zjv/6oB138gjxAsJpLiIH4eAHsAh
7yMXT1t+4A83rD+AHN+TQYkDAUHLc45QjTIRREyvagYaJ8qZ8QI5zGYTV8OMsgHC
nT1o+Do6mZswyByMFgNvgC0zYMOW2bZsFTeVSi/3fSMcvwTBoLEt1K9o2nyJftbB
NvaOP4xljudYV2mrlFj3gb8mOd2fyqaU01iEibZ4oNyEOBZXrkpYHs0IvRt/q69Z
cMT5c+ms3yK9+bC4qZkyvpiwdTtoCToxpGQRz59ZOJkty50EyBXgZJjr9jPY6UP/
WgjvuZhZYINVT6S5+BN9Sm5YJ24D6BQ5wfcMc7mV3VFONsTHqptlwihjuIsMiyHx
I530RwzPpkzqzqmjwh+q9hOud+uHL+MaXVotz1pJT0esuTWuuNpdJiOc+uQEpQr+
2r92Pa7kjzwx2FzuX5KdXvZBlst/TCFJGYPY1njE/UjfkGwEd8i1ge0K6hZaaOpG
7oH+ReLosdPGPmZLHuozfQmTr3gU17Yp+F7L9YZ8J+GZfRqWqJ4HGocCHtUrmqyA
7/GqnPDdxICs7oboQFnVHqWmnBqv45hlDs4kJRaoy26UDWGqfTZOsc/P4Hwl73Zm
X/TenClZWETV0bzGUNfwiuk/oh5HVnzJqjHxAurEo1VJJ8GLK98IyEuY8nXcCYnj
sQvMngzhtre8IngwxpetRVZvWgwWsp2+FaNVl0TDqG9rapLIxRdMDURC3sKdb4KM
9HF5onxyY3XLfDUEfy6uWH1lsJA8wNm5ZXlB7sAil+/7+CwRqoJ5Xoj/H8nvGMnG
u8muOOcSYawQL6BhZ55IRbo4zTs0ScbnDx6TSlzXGn2oTFlq3ZYzFLjdJV9EE3Nc
cRMrRkEAGuQydYCtmtq/arildHvBHJ0NsU53Pnjf8XIOwJhJFlbthcsqbmM3oLpq
4ysCFaOUyf78iBrJCOmVH2n3d4x/K9Hefh3SXNFlJaFSElUl/vFKVDBjUW/ABPFg
kuZRG3eI0ZX0RzLS7mmlebqC+H03qMLzqhWp9ohI6fq7BAMiil26tOy8cev/zjki
IaK9MkCFqp4lHibUnN+xiyhZqUw/2mORToC9ll2imYLF73MD3lCAuX9l9KAZWWFD
7hMAemX/dIiCm644I2MT6zFJJWrTyByCuaywZf4c3Cu/eVwmb8ZcKfsG/NLabWGr
rk/NmkmUe+CNTC+2/0qKDdOTyRpmBR0RCd5MpwqgH3/0WG7U9tn1VtxTRlF52xo6
qrxyA0uaCEiZjhi6p6vtQgqMmUZXLTYks11wyNuVHSQS1vZI/A9HTWKcctiWMGRI
mO7dW8SGIOd5PJoTUy7JMKESp9/Q9ACmSj/OjgpLEkAMAr5q3UYhVx1eRMg28UeU
N5vbMak/4Zve4uFRQBaSuYUxMO3Lw6nTOCRfK6jZKf86UNbXGfDp3+Pp4Blo6enG
VlKfzLxN0jEsASU3xSJwT5CtJHzUcFSBOl3fddkxKAC0RYv+xpC85hgnll9oL4MT
mB5ks4Haz+ViyEESRXfru05dkGHVj2ciYnh1OnPoMS+WJLGKJGhPb4uvkAWB4SFn
1LfvY7o6r3X55W32RjhZ6qZerK432HZQFV6y6ySRkjq3YNWCFgFIKBf0693/WzYW
XG3J4e0/iNWnnV+kb/zJ2XKyJl+565O3mvJw0JmgXWgeFY1x27MV7d/hNp3yWQZ6
G9ZAe8eQKeWNrPl1yLorsOr3hxdwgminiOr7O0ChdaKrbdfa4k1ZpK/aFry4XZNm
SGjodghWqCYmVJ8E2/2oTxuKqsKeGN4/CAtvocpSZkWRTfBCPyTO3bZt5fe7vjrQ
AuHsg/obLkkVydN9qPh2/5G6oiJPz5pD/bgm2XFRwUuomzL4JnXSpO6DfB1l9KuU
fmmo9p+VuLtgHJyTS9LUfv/HqIvTpg/zvhJ4sV0SjsfFEZ/Q7GEIEv6TueZWLosl
7+GPHS56V4FdTG7XQv5Ta9nfXEsQM1i6OQRI6c0S80RpDBeekrRuwjkR58vCXYJa
eOCV/OBVI81ZXiF+HFLN+TmlVZPkO69wteVB1c7XwJJYgZ7SPqUR5CPO2sgIWqp9
nnbnCbGlxCZVFmURLgjSDloz74qMqjYBHXcmvau/sPMnOahpb41pOIKQ6xzl1f/h
3U/5UoBCofB056bjm16MqjKKmmoujlcd1AgGlpS92M6YmFfetsBaI11FdDviN1CO
thZKfHsAfv8dMK9aHj8u6H6WlhGUXQg92DFDVAmo0/ybYTLx1SF/eH/EaJvf3iJn
VSdZoufR3eTtemq1ltCHvnPZWMJoIFHuKhn8i2Z+16L1ZlNQTJ9qTz+hml2girAi
H/JafFHNw9az9+3APsA7SIhZFMKHVkyvXpxa5gNAqzQitGwVbIBxaSn143kMh3AW
Os3A1ZT2jTNgTNW+tfjuK82APfazcvxHsYOPTUa5Us6AXxfmJvRT1fr5BDt/L+fN
7zy/zx9m7m8STVh/Kc8o+jPgjTpU/GA7WOqcGEN5UlVxD1ZBYSZsuYGgScBqy0QY
awkogHFWmPEZZepBEtBHNhtptDb+ZfpS6Vze12n4utWCxBoTqLbwCAqHHu+8DoKq
m9Zot5zNRX9useA0+7cSDplck7us5nDaBCeCE1mk+ktOivTLUIp/HUJaBguPWNJD
kZntfcYgQrUyTCKoALQfIS3sqAOTtg1q74U6NQ8BawmHg+xCqIB6PsMp8bSMh6gs
Q1699Jp3mScm1d6aI7F7GZ7euvzyWd0TMD9eeKt5+YPTy14VRbvugOvpxXOWmFzY
73mApAVkonWZP9Z+fOJ9t0p3X6DOiXgZBWFzka6OPbQB3GGQR6ahK7YBbmQku0/H
Ev1QGrm5IAFMUL7Q3rK0OvUhDH/JVqFF4UZ+Fjd2rDgBBefzoVZDpPRRdBtXA87O
FGaGMpDFhsQwrURTNfNGiabCI6WYjBtssfNqKEqDPLhthdasGvLHwFQhbaSt0qcm
T5cMyOI8FeFHr8J551z/JafmX0SvC5Sy6GxTeMGUIThOVLiPpdZE1Ik3Ib9MmPnG
vZcq4jHCDs+e2p3wdBEy/wxbHlDcxeVNNMlD0cdStBcucg0r1nVaq2lABL+pgRfs
rb/SPJO1b1ZVp39hxDEqD91eHIq3E35mkeeWovS8EkQqfDrponB3v7IjG1igQ2WO
INC5cOfGwwCgGPQQh+EW07NOjIe0MBKBqR36vSPbA4CQx8sCylFt4FtnloTnHGfM
P+On9rAUbCwgFPzhSYUlzK/y02nmKQw4k6AqJpXUZWN/Rs2QfhzrXHsfqjEDby67
wo0PVVQQujtD+nnXmPnd8FGuwp7VOdYV0awqGyor+Q6a/bMp61NoHCddS591IkW/
gncJV4YgxqfHnfRCMaGt0DRrS12Dp5jtt0dUKLKa9kuRGnBwpZivB7H6Na7r1gCp
8LNqJUCk+eUalSAZZ5ZATfVwaB8Lq7ieGVlmvU6TDc6UXfV4c981yhsnutx5H+GF
qyndQJkix9k8Y+3xsmYu2jJaFpPFR6nY2A6I2+AhTAojmjrHXXyCNRTKIwZEvpFn
PfKCveeU30VKY6p17JoVML1YpzMIo3pefpw8XoCcPMNOxDvB49rA1kzikT+2NRfZ
9r3sj9rzku1hY19Gr4foHd29whBIGRcJbjeGH7E95oCf6kekX5aq/y5jgTAajMPU
GiZej73lho1uGJRjRgjK470JTdQoU6my5z+mE5ZL+W62R1v5FZiOjwBPNngNc7cT
QrTWzXEdYs8Iektfz9/DfbhU89/fF54Sg15NX2NUTPCXFWXtXagE7SZasj5b9qvi
o1J/vQ80ZCRsL+LT56gqs4UFjSUL9Ia0c12p+E2bRfZQufUg4+XBVJu7v7rduUCT
A19H1U+VVl1zRLuGla81M/8shiJ/gpo7Vzsmn8ndm7qC37MZVzVaC2ko3xj93F5g
bW9osXAUFaF01PSznSnVt7lI32YkW0i5JiHsXUaysmo8gRc0Fv9kKQsW0ernvKCj
9cY10MhpfsLDOQm/QcQid7kx3t8vbmrMFgIO4nDGIWscrIgFNYtQ2Eg9rd4vHJZE
3aJIoaOVOjPj20OSo6Z3oQs4VVeok0TwcHoWkNeMcckHjJkktmOl8XmeQkPEHAUG
EHzSykGGZaqw72Zf4dUqhTj9vdX0tbVgvZ9cOvSqKG2riUB8AmfhfQUxH0ES4SAS
fiZuNhctj+ij+PWWawapjAv9Fh0CITeIgGiVlKYRzIDc0Ne9HfQS1LyhfqevcB7s
Kom/dfsgRGadeb83GPZl0evuxKaajxmGTJAh8E6u4UOPMNxMqkgylSLaogRQUUqF
/g9lsTJZ3BBeHUeByUjlrbn66tVieLr4hMLSd0fZYlMfBIjzxckInJUf+LVLJGK+
g37vBfU0QAenfDOLilSQ7dfWte9IDrwKVimuR+8qwW5PI2mst6ke3BBgkctsfPSx
/fdlxh3opgtvbZq+2KFh9+I3peg9mZUGCs97MqPTN6pZ9VO9l6FMxF96/OA/XcYN
1ez/bJwZhbBzAjucdZ0a1khNUjm8CYPwjWYUqnw3CFPuoRKmY1ifyuUQCtb1eYMv
PZ8/NgYsKk4aSd80ZDqMqcjwHnEfuMXeVskZ8GNnLfNaaS2lB76uMgExKImqFS0V
Rnf1TTgGjyfZ3NjkwfSDE+r+G775UesoQCRO8LlbDLcXlVtwCq80OXALFXOUP04I
UMpuXZNYya45rCVKP/O30up1zoW80FH4Oxz/Ql4VAy9mDF5kXChPk27p2n1Qjbop
IELUA2DQBc9frpEimZDVNkLoYTLrIqEmAGcjtmJpZMZb6KO2NVVeaQ2pHzhfr8PN
9xUQmoFsF89KMBRcBfUTUpC+Is7665d7Xd7B0wSfZE4MQSnBB0zks2GB3hHem1Ms
gUityLCw70G/7B0nd0rQJNjYv+0raWCb7KOS4yThwve8T5Gcyz7FJV+yxDew744W
XegVgzYHbYUW28+LwLujYy39n2nX50u4hxkvxiKMQ43gjkfsVL7gcKGR7NecZcLm
i/7IO9YlW/2MCge9HVpOa7MOEo1w8zGPDGY8XDxbaKqEOzV6jn6MLvwEBbYFM5Sg
YjNhazvuRgktetDx0vycUW32zEYK3oZDFwvliqy60APVV7xcDOYEJKT0KNHKL0xU
FYN2AtHD2Iswbtm0X/5BrIdEBpZx0wG+7zsxr9dgvWH1xWuvKY/A/CKyaOg8YnDP
8E4HR75AIJqj3v3+GweOQ738xeJ/uNPSEbErKcrflhIB+rp8OGwY+pYVOmRvfvTz
ou0Xog4pooS1s5fZbHc7m4ZD/b4fhC5ui5U3uqqdV3cDXRu3NOtDQInTZ08fwMfh
Jug+FKDeBtvoz8O3Itig3pGrTzNKoAgWcjT389G7Y2e3Y7RBapJyjsIs7R4asqi4
RPoli9/bfImZoPCM8lAp5+SgT9KcLqbsiti3VkWVBAlIzMusdwum19MoQvMkOmcJ
b7SpFpi0C1YWX/OD8SNX6h55g5Tbc9rhn+j184I/Jj0psAdp1jNYaAIjUD27mt07
9Lrm4/WctZjAQ+x6xRtOkUFSC0MPtHjpFGx8BN1GVpAxcKvH2qe+zHSX427MA2TG
z/nJIDR+CNDAgL9MdbeI81Wl2c6FCf7Hd/+W1y3EQJ/8YSh76uBCmaYIX0Ao/mE/
3Oq4hWwgRx3CdH+Bs84gKjcY1xkb6JuwIUWaz1nGfcT3XpsbwitCQJVKLwRnUMfy
pFSlFg/glmEb3Ql2n7DdzXvGOrGsChAKLhgPJonbmxO9SRMRn8GPze7WVsKZgrp5
9ESkxT6uZFyhvrlr5Bu7Ru7KdjSlS2uksw5+dBbdHEuQZib2ApwNGG+vuVOvSCS5
FpzOFRg17CUlHUvmdYHA0nrh9tnZ7w4EYtUx0+B9UC0VnNmcISYobgimEOE0jB54
Ssd7/Bz8UJm5BmqIdWRtYEvL9NGdgnDlL/A2nzk7jddP/8EC5Dsf0tEqsScOnE+i
RH3XogzFmMCp8Ez9SsZzcZsOhA11HySNbxHCkUT5xu9IKNNlsoroLp7nIcy1jcqZ
2C/tNOu04/9EUkzDrOP3nMlCRbHiewWG938Z1Cy7PIBd73F31X2QXjriVxEnBI18
ylfX/siHmmrwstVCVkZczH8aewqyqwBsssYOvoZqJ2N/QA7sANIPqZD+sMUZ/t/F
ls0WW9YgKlfRVSCC4RORbiYe28zDSRRZDjJCA76kltMtbCvc3NatoAETtI+cQuKt
tI6pu/B4UGdFDbj0Y5VUA5kY7AlHgc1ONJ+R2PxsKbHvsMWuNI414b0EY9mUMu89
yqyau0Acjv1//hgTW+qI4lAPIMpBHcp7DtXO328fOLZPlJsPJysh9ZLK2LiFxbJV
A8yr8CbNnxDnGoRynpsLS8VAFZbsqJf+BidLiUcfjaIn3bNQuQQdAVq8gVKc2Erq
ODGn+3plhUsSC032mYa/9yEfiwvIwmI1tEYRsIkM5rwD9TsQ7o2OrtG8iCncA36i
pQQAuDn6L3fTUyyXD9IKycuCtu1/Cq+FgM0Na5ut/yTIv67bnfnLiYeytNSa7E/Z
M9Wb/f6XH3ZLPjzbFkWmOdnM3DljoRBE9JQ86z9ra4N6jLe1l7mTS7ToBHe6Duif
hd5KmKwyZ0CtvgHGjGDZtk8iYg9MVeD08YuXozuQ8Wc75R189slnyHgg3hdM8HHC
JZT0rqh4oPtayHjOZZvlaQ5TTrGGBgjYUYeo5ujoUblC60qrKu/mu+xSzTLbtDxD
tCV8hEHUiS5Qj+Mu0qj5Biq9HZTLtd6VCFUCJ1WLd/J4BXJ7Bhr+fPeNJElvcodi
0vtPF4N7ZA6FQNkWQSfjeVmzvvj73IhcFBNNQbpSoAd7NjTYlgJr0OKVRFhf32Al
hTT2j6KQNCjNHthjhHdDLwNg6FRd11uINCZcLipCze9jvZpe/rWG9TGmWpb9sr6W
jvEtXPGczPl4+yWRrqlSKzo2SGVdQMCyhf6mO5d1MU40CA1m+eCqNkmVuLQ0b5WU
I+sedEJUGwYxP427w6v639DkutXsrIL9pr2BQMjoBVmb8ayK1PHg6PjeTh+F7Pmp
tHHpNx7+qzEs6XmSDzQtRnNlTiOzFRzmSVDbyefxsq1BlMFFoN8kgVVpbn8JtdlD
wV6Tu3V54oViIsJGnApH1EihUlCN1MTIkNeIfMYC620d2FgW37rgTzZfJwSyAAyT
UtGRzKqoylZgC/dSDXucBU5F//TBIZptypRwh6maXK7ckG6iclrJtbRiaZFRMe2s
n3FD6R5BlPZAUdNKicvNqQhN3hH8wHnwp6KQHHS7B/FenbEdbW6xJPRm4AinhVc5
6MqEJenQPj+Wj/YQ8EvEwHy1cf25xpZ4G6u2nqncJoKDJ6IEqfVhPrV4mOkIMOBQ
mdhBjR89/hlaQ7cYUzyOHPrrKQzQd37QP2GeKz6vJyZYIBPkYSA1ADpQteXmwTQc
B9lGY4fKlfQtxdzhfPTWYiQiacvhS/WypY9WGCUVRVNEdMHqYZoiYIMOaT2cdxE/
bt/jmIxe6twGI/A6cWD256wOehqkdnoGB4XXlmTNC0C6EHin719RqsNIN/codSYs
1+O4Y17BkIoq/RbV3aHBJ+C8ytio6+8Pz5tm850vQ08ih6ST4LZrGuySIiW0wiJ5
6YkYgk315lDXxmJ0cTFG5qro00jaxUKl1oRCa32qtNWi5OLvwsIw3gl5G1Ic0QX1
nRaKl1KgA+aKv30SvcPzaOW94BAN7V86ObYcUgVbymoYMjEVzZO+SZHjXgwh4poP
phTRrP9MzYdwIM9bHS0t7zv0oI7HagBTUtOrh0JqgTnJN3iuBDSZAdts5aCBte5O
Co2WVh/de3i74onO1kmmzgm0/hop9AYf4PNEcrg/II6d8MdSIBUXdfb9betu/1M2
WWUo8tGh1kMJIc+2VfR61G2MnyViMw7wtezAM7YinFZQ8GJ7Nhl36vedeobH3RDZ
5hlbSHvIAOZBHcJ6lrNNX5gZ2Lp+OkBXkDpEVndZuV+MJNxgXBnvZH/ognuKmM5z
nike/7ngEFEUdxnlTc5Wlgt9spI5tJGGHjSTWymzrJAMOu96KrrPwatv3RsySxO7
JYWpa4a1kUGI8sYFkayNs5dlWKV9Eib29zU7aAB/KL/RERB4zw8q0R9+Tz1qxn75
/zGfXMlMawxmopJ0G5/qJLAKhfvt/MFoTkBoDnjNiQQ4cy5ioQF6sY2GWgHJGqjf
ztOPWpZ/ww8tkCKG78BJurWesQraRYInUi596bGGVV9kV7YL0F4K6QRumWEpNAW9
UwYERYgHTGyps6dA6tzI0b/5PUtq+1ocEJn0704Ca4Gmgt2+Si7Ep6qy1i7Sp4EB
QV4xn5m1ur3wThR30+7PWF3G3c8HUIvbaqFjoYPi05l1wqGUp+ZXCzR3QmzIGozg
dBwxlGMm8yJMZFIO1+BllbivS0uuS8VawyL0rIFEMT55hYBbf+Ga9Dvc/jYFlLhB
A3/URRlzwTvB12KekwQJm/Dr0CZODCW97snb7WlBlYY/zGP2ylIG2nQ9AqnhvkTe
Z24Ya7x6cc0dLbyLqZHD9dBd35aFzF+jgg8/LZYLtApLRXw3/8GhpbGcK+OjrlSU
ebXlhFHMcWjYumdaS2d6N6vAWylK5ihc90vnHvDtMc6tyMil9kyjxTK9vSCQRxem
bCaA7QO8bfVGwSsA7CSwBmUsuZEzwVDVRmjnap/QJdzOC7ghpg0axxfLLSfNXiCW
1kDPQ13N7Ykgz79Cf60RqIgts562rj2+ubGRjACEB5u1yrO8ttlxmloigREr352l
1pVs+FItGjdMuLgrvH8w2jcIbVaLM9uLNPfRLVObWs250qdoYfoOEHsLA+QgQFK+
s/M7RG7WJKUjgBLDqQVwYALtUTDbkBvczmrmwN7xHIN3lmAyFRDNIXLLYmNQU+VF
n3W14y2AEr/jY9v6xPmtqyWViyZnxQdNA5uYfEHVlIkGDqmNPCZnPaLppYtcaf9a
mYceLJySAJb2voE6GPMn9I2DE9E1YwOAXooais0moWfUZblChHlbU9wpdSaI+ZXG
dBN+P15djiKMjuaJ/vO+jBISk22jvTxKnNoOxOUCmeXpV6CY8uEnxtArYV6eQGmC
Loly8me0ZPKPS58EQ8/Q7uOcjkImsjHt4t+ymnU8WswSqui+glwUsyrARK+FQi09
PWuL26n1hbPrnyhtm1Qp8LBDADFfrE7s+Cn0h3w+rAPLrVYPeUifAS282mVLRYM7
2qZpRomUK1g2bEz6YM8v6vC8BPN/j7lDIvxUj4DLyZBHO6gxbivltCwWraspTjIc
BhTPrmROEtIF6NMZskcfchiZWiaY/+kSqGgfB8tVgSAmDpe3srxS3lee3qzU1Wz3
RABqXIFE6sU3MCywQQAmyvZjif08hrEP7ug8Uu9SfodzkY6lpHdshHPH6mLyQVdk
N9oAS9kqIqUto3PJfqoUwwuShI3md3kJiz5r6Q0QJS6J8vp/GTpcAseJ45K9Mkog
6IKyStP319/aJbv/ZWLlCjAkaBOwrwJM2rGJi3V4ZikN0fgCIR8EF+zCGuyVLnLb
oppqABwsdfxleR73WY9JvCGurB4lSypCjOWSct+ITOOmRSTbgidfba7BX9AHXX89
wT1UicBeNbZZBwzSKH4aio9mn28/VHirbDZeurvuMUmQ/vUuocwpJclPnEuYQm4o
lZ7S8vGUkX8/rTi163baK4xx1Bzw/BU2h6hDYD7NWKot9WU+BQrbN15pnQa2NLdc
9dRfZjADPBBqGPOplIeCkfqmNVl79Ki5OlG0QONtnPQWKN6ohLuvYzDd1m8m3Rys
kCNYxRRNq+y5EQ6NUU3i1OOpZ31VB4GT7cUpti5yLIUsWhxpJ3Mahed/4K0cUje3
7C1OYMBpBt04maBUjLOZw9vSHmiyFKfaqgsRyMHwnxZ6IEIkKnnMh2uio+laKwoK
Shnat20AU6wGzPJYTzLoWqxDeE1MAf8NNE+Rh6r1Yt1zJXHb/KyX3V9UI8s6SRh1
99GZAZ4Ho5X2Gw1nwppLkJXuQObLduQLSU1ekdkxms95puCkEH93/vK9F8IdjZUS
9o48erZTE6WRFz2EePlMs2nZCJAry/4L/t6dtIc79bFainGE2TV3ppVAu/moCNAx
NBKK+OSOrb/kdHq4Cx03Y2DjRRbjZLcxu6behEiwyVB2hc8seNQf/94T44LA2sYc
pOoR8q/z+4H4SGgS66+HyUtBAoJmbBg5yYw2we04kPINa6fP7nwy/j/X14XXEXTX
MlJLp8S8V7mUTJFlBtPwWAdNmjmRsl99iWbpskWq1X++kjh9PuloWQgnhvpq4r0v
KGBCxmO0l0jJi66cvxiPhV2v0IFFEz3MvJbq0cetxsibmtx2lY4c2lk5IiMraDrx
Ha6VBvm35OmgpTVh4hmNkvrHmBRA/Dz27Nd2ndRV+/r0JMvIzGcCWYDPuFweZogD
Xi63dDjVXwKaz7MrQNM47fve3QTv46oiwFIDbm+rqKXCXUupFhQKNIFEgLJE6gGJ
SdMchL+5P438cekQy4HW2YP9M1JeM+R5gIziNsoI2CXhZ3JcVXxCRdQQoUZ/hRuO
pIhJVoxBMYizKGFDz9fp9uIoZgb8WoryFewqbyno1JvhUoOAYvZ2UABC2sIV3exy
AEs4rcnXjA0o+1G0E3N4FLllzscdEak2A9HpSUASTbB//g912PEVqYK9PUTGcH4g
jon5i8kFhhIVmUO3S2bIcaEAKhZ5zPOLWWPEznDChzPfroL08o0AzgjWRAzUHuPP
b09diaN+dXSfzIcad+Fe2a5rbtUbw/HDe8Y21rbF5MzCQ4+IQXxUDAPN4VkBYvdZ
ITyhzOcEabMDSR/0sW2eixNTrNeM7YBWfaXvoT/hEz+VNLuWsuZ+/AUfRYWC5ngW
wgxO0l7quTgDdl/eRDXnhzlyLkRHmbuJYAmNsi/+dE7e/vs7Gp2Bsv2s5JragYVh
rh7/X4jPc+pIXf1qSd9Pa5YovW3E+StlGmAM0DKsjU3HYfkuuJd+bhPaQP6NV9wT
3l1YHaFBzXKuDnmduadW0kqMGKSW9jqC/L4+oGn6JwgfdBlf++7L5eA5+EY10hhA
QbrwEg0LL2hhfcekMixfBy/JLSDB22Re2TemxuymUGd/MOHUDGT27P1JbrcVx37P
BABW8lHZSgOsBrNHv53o7PZAFt/8DbAryDqShY/souHQDMIaK0PFsBqLBQD8I06U
IveDBDFhWpP/iCuU9CNHCvfT3DuuU/VeIUm3wQnvsR1IWShVSEbL+guKJhaJ8DKp
u5G/J2PG7AwVF2bi6u7Q5ddUPoYd3d1eETsDdBzWGImxjyv02P7bRWRTyteMoYaz
yXZGoONBW/JPl1/FnuTpoLM+e7iasZSHWgxcVbNB8kWhiluww2qZEfgAfHlYMjxD
NaExhkSnHC44RJ6cbQ+KvfuIZ8+gjW0Dkes8h0uvAvX45E2vfLXAg6vzJyGgTLFM
Gm8X6rT2K35z+asPoPUzv44E3k7CKxmBXl4efghPuB0PkFOACMQqpWB+775+2RRE
ceVQYOgGKPJOfq9KfmvXDgORdT63tAQVHa/sdvejljZW95i5Wv5bDDF3lC9c99J3
fxbTiCdsoVpc5B1TcF7SflNsm6nfKD7RA7aYXvyT8o1off4ZuIHJ/H+BareeB1uf
wGs5SA9buyye14uWzz5GRqr07stDCdJrSkyOEA1zXMjLIBBGEBBrZA7dgsMwlmMD
yqjdA3y9HJ6Mc/Xm7Ve1d2xcppwjXCYyP5cYd/S9ET4NiLG9M09hmy+dxxM781Tm
4p+Gsjm0uG3KLvZsrX7+14JQw7DSrNdKyLXgOxZAKRi7zRjCKtHalh2i8iPw6xjO
yQ3DMWcVv/B1nl+Xv++s/ATTS+ltB305Ontf7GQ0SfaYVxAepJMRAnJt58Ir/BuN
JDsd1YRE3YQxrqpUawhCgH9aZyGchVS3Yh4jphfRgfmiPCzsC9+zbdcEdJw9Ywnc
iUFaTkf7M5QhoiXC4rGtdjzReLTySsMSMjH/TyKELrMIsiBijjWvlEAHMgDg2nOi
NRC71pnUasgyJqxSsDlBL7FtNZq9u6WM8Ipg3q11eStniw/dyR5wiyxu2HDWmQRo
3PEIYmeEp4Q9JkSqfu0pOZJo24hS42tifxPlcK9vgZqbKtXpwYzaL84clT4zcJVG
IErQuq4rWSkhiQxo6wxwia09wliBCBlWV1X7WDnocgOuJI685FuWN/aLSaa4dFlu
UnQMgEhZ577jmDlPHFrzr4puqOOoFB7vnHslFRW4NOCBLNwzf37Xly25r0mf2eB6
wi+P85aIl6Fjl65v75cVYTMkpdJ+7Lv3cuFjXdy8SE652MTvSe7a2Lc+vZiWonGQ
NxK28BzUHM+B792WHluKHuW4KpyxnrdQt57rHrvBLDs5drGOY6wLYIdrvCxKySi3
KFe35uaz5rY8+oxZI1IVELQu//gHXhyrqz7aS/N3bl0i063+D581N3ZX6laC1gj2
boz/B5eLQRng+bJA5wdpb2RHHsX4gs46r3uJ3P8v8ckLVgNR+7si1WpEp8P/SEz0
bsR8vVzzL9SU9+oipepkxjtM5hh7z/qZYmZEf4+rg/3Yjf9BEd/5jHo9+MZJgYmU
AhD4tk9gKk/tA8oS3jY9foYyyINyOdJi9O38zPcrQIa3Tk1zb56KtZgmnMWYb0kv
3dDHEdHnZ73SDXPPi09hd6n6f+DZbbdPgZgunqUyCq3Gsi8TOwSbe4xAfvdY1Khn
PEVzezkj0DHzpsBu07OdKbdN6jwt1IZu89LmVcRG6ELhWTdvRB2OE2MsRHdSHbp4
xM4yaqBjgiQaa+8pem9KuQAFB9JBmE3C5eRnLsDwYJj7vxOnSQEmSJaHMRai7Yuj
sQWgQeZ+K+N58bg2gdO60G1BsjGO/n3HiYUuT3Sw/qc0tQrsCNcob+NOYlGihjXK
PGK7yxQtY5Wje3c6zlmkwOsmIMgubiwMcbvRB+pJMyRTpCKNLWuYzvTAnba9nLod
L85+8KW21AojkYCoEaglj78p+zg3skNYRdpKrZPNuyWNT+LIWHHyv57mwQwIylJc
auVfNHO4WF4utqxtl3PPT3g7vp334BvUevDxrXbzRKcgd4rDqPCVuJ0LglsICTmz
7W2oqQ7Sgclu7G53IuASFqOAmVim73c6KwntnId18vOhE4Y7NHIZiCmcWc7/Vtlg
VNERvVItq+IkQpPyUa8YxLCGIupTAk9UViPsjjvH+sg992/d+WgUGbAfu3WDUZ8D
ri/mq7TTK9u5yQ2ARhsyO6e/Ir2wvfyKD7iG8ujqXAN0WaVHHCSVZlQfQVkAas6I
pfv9NjhfC7S3cMg13p9+KqKRo/ldi9KpaNgF4Xc4qsxKAYEwheJ6eSN/CoW1RL7Y
RHH/lERRkS2Gauz8AgBeVAF26FgkgS9Z1RaFKEQVCccoEiI2cQGPDnjMPyusI1UU
n0oCXFttK0qfjsYFIgA7BZiFgxwJBBsViRD9dCRx13TBQ9+N88z32XMRX/6679Sp
B/cW2ofywQTfVUt4895+XZnhpNWCBSO9OJNEKVWSQv3Vhs6eppv2ch+2jHllyVsU
Y0D/Z1FhEYxbvsi0yQglhXQPPtMuwux9ZMMezsg2e6MHtHsopO33wQf+BFPwfp8t
zQ53oPj7tWnlk4aUHrLavPSP6HaUVA7B+0887mIDpWz/EcTKTJe300uOVbBEWpsi
MN+wV7pn+bLtSTwexPbEfIOV8wtK40rmN8BIRCG4s3zR42iKBEmCw4aKSUBGVlqM
kFUyu/kNPXt0UifnG3YG/i6WUwTg1L8p1SsLnvX3ZcupaNI4ojd6e2dr4YXUU2EU
vitrGuyKVJ+b4KGYa+qOim1DiMcz+AU4jGSROJ2lVSbdW9tDKn2u5o3RkA+z8FPz
jdXglypUPWOaHuJwFBtvwcj5DRFS61X4VHbD7NJH1DSH+MaraJJzjEwaA3WkEI6a
BXU4DTdSzEUPhuWC774dFFEgmt1Y1mOb5JuxHhO4L9jmdQz510c0/eV5HeawhNGY
JNFZUDfWVgy7m+LphuNexwD5LlwbQFrTCNtCgKTC8wYDUbYc8kTVRlxT/uhi41gL
cQ/aXf80gX228p2ODXjsoeS49a2lNOEWZq/arWQMmOBDBaLlq9i8N8LIvA+bTtsi
kbFwgRbAzUsJhoMwsrRjvM/a4VxSjWPr8WQM0YYAA/qmqQ/CwOZOnUoGaDoj8FCU
RPtcfYOq9X0DVb8m/g8bYIf6+4JXFYPYaZtHruwf8VfSuwiqhEln+k+SFZhJRw44
X6wsRZKs7x65KNzNH0OUV66zxI8d2anhoRLrANz75fbx5yl1vzTqTb3KJ9uaS1QD
Ibm5eHUXY31HFEtD8tDECbFCS72hG6kWt4XSq1fslv8u8A5IocYBfgFji4oz6ToV
aMGOFpeAiFCS/0aHg7N27gW9a+l4oIV7Oc9B4G0ktjP4yX/XwGsqJb0crQlXJS8k
70X7EVdBFvj+zh4CB2qXc55L4xZJPJno1iusUOzySTwpTo4lohWpqd9qFM85NlAN
dxOyB71RjaA0bFSb2Yyt0EdYeNAWJSo3CzxT0you5xRxCdkWkshI6haJz1sGXRdj
sGo2CR1un4porhK2cf8pNPPJ4PMBUYvq5/UDbon4nSjLsUXqXokvKaTeRrcziJoB
aQ/DQ41VuiXoBPthLMxUQKMV93NWztcM+qPCWQvXJhi8iVZt7T/lL4DOBgFKRWl3
QlNKjAfWIPXe/tn1U6+vvoVjSHR+dLFKhMbuIbeRWn0q1++SAF4VgUWt+qBQo7o/
XbKj5QO3sUD8iJuwsykXKpuVCaJP97nnKIMKjTXQYX7bYrt1DCxVGs0b5egdkp/d
HJW/iNMbreX51kyFXWNsskRt9zOJGBkRjdI6HnJjZ3QWsXh2QUTKYEzR4sXsGrLj
DX+CpHxiR4EjLQo9ZtcvUiZrJjHuO17wncH0PzrHDla7laYcur507w4YK1stBQGc
OFZ81ZptaGq338q6iGO40gvNJfhkTX6bnUtFri8qeMbEEwJJNLxrRZPw5agEeK2i
KasIuGBYSrg6Ph5N00nP2GUYFasgx8ovQk3nNocwju3Hh5AvevhrXl/6ybip7VPQ
VWo/3eODk356X2R2Y/ZoPgvKI4N9oRXawTYdd7aVoQZ00DAZ1VUcyVPdMvUHiu3k
pg59WwnEu7aTyP7NKVoAwul6ws5DqK099ok9aL6s/gLFSQ30+P2lm0PjIeNB1aB6
wt/oF8OqcgemogIb4HSAH1XjZYIsAU4q1T+sg2Nng5zuf08++UkJ+mwi7OOdvCsc
kokikNrFUjgrE/n75P9MS1RyRRfuQGpUsSOkABfhJGYUCJg00bLRyaQ5BjIDqrsr
80kVR8gfXYCa6bUauajs/V0M8KrxJmGaDU0woC6oqdVXFVlzeS01eoNcRy/UMP+q
EmLb/bNRft//zLmjkSAVJMWwJkyS1PPOpFZtb53P/Er3MPPpc3N1yGzM7rN7hULS
whjpRcbf8V5QUCG5W2Ah0ce2AlcHhwZDA6WoccFIgUDoS6tcRu6PeR5/cuCaUVjV
O3Lx7PJvbeb7pdhv4ShafcBU3T+y53vh3uJdLb091P0YWMDjUC7MtJrj7iubfiIY
ggsFd0gKI8AzZDfI0e+iUBhyGWFv2dt2N1GPNaMbipM6RxC4UrLrrWjz3OqevAwi
Ebfq+Q4tpGqzgIk4jeovJ2oHpvbuW2TxTXH+on1X/HW1sUqhGa8xnCS/x8+K2Y9q
IH47AxSlb5qf2c9Bue7y6oFywMS0/MYU9b5m89Ex97QV4vbHvJFE9X31Bu6hlPHG
6G9b2h1SWC/Z4HRl6ZFOUHiQdGySqUsDVMIw9+2TZ7jWUmdhyE4kwWBVH+naEDSL
4CGLELWlnVvnpTMe1Cgc5Y+/z6eIMrcPHq8QbnHxRm2BXjnB/LBsaXTK5lz7Gjkm
mV405qxM1P7AG3F9RZ/JGHKJ2aeVWN34LGus73Q9Oo35oA+UnyaQBzLvm4QWzwfO
8M1MqWgMSzqkBVmmS3SCV0jMorZRFk8PdNwt/iN3n2gmkFZxk1gcDlxlEYDwyXPj
Ohgs31mGORRGE0o6qQOYnCWlU2XYHHuHw43qTOIGY1QKk0BaQKHDr+AmBu07Ilh/
gi4j/6kbg78vYlFRcZxK9SsbAPy5T8KNKbWXzoszzjE9AeF/d/NMTl8Lf7sLFOAT
bt+2KvuYyLeBIG4V945yXS0EHYnhLE6QeRbo5TruCZT6VosOfVoIcauOEAMWt9yt
KS5snnqvr35y3yLpQGIDnQTwQIhTkZ8OzjP3AQ5DBvPaKexOCAzUqDzzGXSVFLRw
46M2KhybVFgjhb6+ZBfvRB32+nE7Cgf4IMY1C4bwY7fxNVYwnGOqgVH5HPlBrXfL
RKtbd+F19fXjQ9MqBA3HEqFj84zV+G2S2mAYdgx1OqXaCh0YD9JexgnRNfiNimXu
EweInn3/9iOETTrSZAjYguVHKI/XKEiVBw2MJZMT5A88cA7rDP5Xla9mqAzkXRIF
6l7uJiD6xQDne3InZaRdmhm6bZvrKmy71RH2xMEBUQwiFCalCCJ0YWpRG+R8llin
R120jZWjmyKKSbzPctJkGYgz1Y3P/w9iFN/BwByklYtU3R0POoQUPq/2Vyfnbm2g
wUh3nsBwJPEqqdcvTrI/k/T2tT/ab8q4vnMP0VafBiX8sD/bvStttYmY23UNNK/E
4CwvY9Q9rKuuGwgnVUoQyQhYvfkwp2UgYRj1XjTUIdM+8Y9NGh1Ez+HFal6I/pNq
7iPItvgp9fbujlZ3bXP0k70IOwpdFyL31W2HS4kFBv5EJWsjmqTzWpqlIFl1YJ/O
iLkK9+y8hCgW5xydUswHZ/Bn94s3jThsk2KA1uENV7hKGSRW5A+A8Bz8GiwmR7yX
R+SQ75en2Z8f9XERUBUGkc9OXWDGw5gG07+mQFdJCI+1JQ/cg06W7mh+6BmxGWk+
FKg+RcaNCUbPk6wjrpQ2CYPQ0Cav5ABhc7Fx95wp9CsMjGdW9M43QF1K3Vjy4B3f
31cK/OPaj8rBXTZ/2GD0W7EzrdIc59j6pAB8x2jMyKLQCZOOxTy3prUPiEADNE3S
vcTRoMFit4EugfSrKjYgSdn8A3BlV9+7JdBBG8Fk0ZxAGcYchitj3Vc/vefc0z7L
uICUSE+kAVfo8iwmXTd6WkSeB5rd8xFgvPQ/qdzmrrH9inVZOttwtET28PDu/uY9
xYpMGB8v7eQ2wQxCxD3hv9k6XjUnsKBvixxzFkehjLCmZP+fXSBEDAuV0jNcarLb
Kz3P2x/gbvsCTkz0HJhk33IYtR4FoMl+dA8ZXHSvsJu2fE1PDDpJD/We66PxbGha
XFxJvZklXqnFaKps6pGGWiYJ3rqkM3IU6AlVULbNqr7XsRrwlIpthtsmjaLgDpfj
8vvk9C16BkgNoCj8I7lZVLakUn/2ULsJbEJMGXxDLFLymvheJMAYS87sjz4mN9Vy
eloGKtomdruPxOeySkiB8xy9yYnWPytSNTyPs3gZSCZlL6ORneOkslBiYWHPmS9p
Vpu3QOzGkp9VT0GMUmkrEC3gm/e/U5i4mBXKWxubPe/FAbOZXuBtr1PAT9ZFuqnK
DVUoshqAfhqourBhocf1KxsyuhV9ZaMhQrDTkUitfI3BYo0CF8WlLI13TSwrzJu8
JnN/o/YNOvJ2QhwpiWN0GUvOJ6hsSz3tDZ4o24/ciMax1rGSeTd26BaswV/ghHSW
sdwC+u6U/v3/8D7jsQluCXTIajG2BO8POA38FRwyG+A4IxpTFpT3HBAIvsZ+GqzZ
40DTruwimZYwnCbrCtRXomxUavLXfhnJptNgTWgJqk42SlVIASvvQMkZLMmMRh6v
ZZsD6YCWah6wuoXk+sHcW9hcadG4/l1UOugNy/IwmsHCKQ4fVivwUP//e5cyqNyq
lUz/rVTvVjb/q1Y8piVjqFFIj4wuIhOcFFpUPyhivTxIZPcI88FTfTZ9mQwS5N1H
pJ/TAkm6H8dNe0i8Tux2LFm9CwL9CflP7dAbrnV+qbHmJkfJc+n7LgUy4M/lIMfv
R9s59RB34khz8UJ543yhlmvBZR7a+JrOlnUTDyqlvvcIo/75x1OUIEAKOv4ggCp3
GM6KcAxmF4zsSUAIY+26rslWdKytSIxwfn48txBo+q9Gozvr8dDvXhG5VnyRYopo
I1lQpWAg0zt+X87YvJ9Q+KA3LetbpWRSbwZ5FU5dppMsOL8EVytnbYj6pjW8/fJ/
hhf2EzNVuagRylwi3dyoT2IPW1ifGP3SzzdtNWBxBzE0XnVUqApF6mHVamOYCnrq
heMfQAVMwkmDiQICQ7det0xtuG+ZPWiDV6V0sCJuaH6cD2G8XiCmdqamnt14txDO
uMZWwWzmFsh7XhMZAFSVcuvfpQPDIpZptQ9H6fPlYeAIGr405REn/B6c9pesbL88
vWcwFXETiYPJFdCAiiE1bTozoJBss/N8m4rF9ItdyeUAx7Oebi1H7JU7u+xhNkiw
6mAVFqSN8nmGKWXAkRo/Kcug3e13tvBndwSyFfUIOAyeNrxRVgR5Z4NC7HkZ1It+
YNyK3uUCwi4gY5VxU3rGs64GvlP9JCfC7z7Iohd8nyXI9iucmuHPi7Fi7bZ0S4vZ
+K22C4x9c9dbbxSDmDF8pl/yvhXvCxEOb0D2ET5Jr9VKQrcGA1TwnpDd7wMHdtOG
X2fVI8yAiDlIKjWNInv4QXS0viOuGkpgA+UJgpU9leMoA9WfcM7VhH4wbSAVvpgj
gWFv7pFCJ6Is2IowuOqDQJ+KPCE/WwtVgAFld1y9iO5Wwybuy2o0J0J5tl59G4XA
VuY8TxxkEDStvaFDA7GsoLWBh8sZih8qPLh6MHX6cBYtGsxglfelpBaWaYtBT8xD
wFrpcId2uIB5+e78V9XiL5+K/NgtXX1j/KJSvInouJwxA1zqh2KC1SX4EW6RRbQN
Lf2UtW8Rr0ZbIdDL73kZoLCHi0s8OKH6FMHMXp0KYtBtp8c59wrl7QXZ5NmMH7lJ
HZFDWc57PUO1H+hOftuvIlK1QX6qOrApHdWJyRzlrXq2E17lmwQdWmXtJQBxFdlQ
TvMbOgTC57J8pvuA28YEk5nOZm8RGe8gAwOiH52Oo9eCtdTfRN7TOOqo+n5OZ3lI
OdgJ+9ES1BBmYlNbbyxwp1DPBsti1Pb7H1JTmZ8oh//z1C9PruejRg2/Z41XcOCq
eWBQu0sazbf9uncnwl80I0G55aRnOtG1ykmaIknAWIuxydMXCY4sLZc/cYm56KGa
k+Z3Pud2Vn5kZ9OvKGWqco5Hjh0aW/m3yiWq/bAL0ILrD97WTOA9YZ77EZ82Abw9
oxEeWfnpt5jP2pk8sYX8kYrvfI3GKieiqgN9ffAcKmi1PPI7SA/+CkOAilWc8xLu
hcM39UuVv1BTbGppSOgJHuPBBQLEos1hYcqQ9/rpqXf1K20eNS4n3la/0y94z/cw
Ta0zb0PanxqHWexnKZYkZsarvq13kbperkxmNUrmahK2HJT2PpoWCdquvH2XnmuP
otjYjv6dlbxhAI8g4oUN8sO8DVQusfAFLNOvnX2bG38OCxOL5okLHJrVBnv5YRJ4
LRdWiVDiuJzYnbjZxooWR54sJViZXs5VlN5m0a8ic0b6lM97sitLsNJWcM/v8uT0
gBNpSgcXzqgsYI3JCMBDkMMhaSk/Iw7jmyMwx2eNmSRc5+n6B/SYD6mhffCbHYpY
c4D183sdaajNnlevEOtCtBUNm3tVCd8d4E+ctPSl/PDLbs/gSg8wSQ/USnIJ7XfN
R5Dojqd9ImqdI5Nb4dESh4EWMNUWTnJFs5bZ12+TtKTOyfxlkr44UdwzgoR78wBl
JwV4kA+BZWtpQFZyZRBZZkScYWAwbdDUoI2eHrhAAJZ2xhxaB7QBqPK2Y+SPGqqF
Xn2QCYPpvB76cRKkjeMPOCh/7Nqd0N3BmAMliQ/0LDDpcj0Xk5kl1bYYvA7m4/Wx
Qh7TPmfj1a3dByqtm1fUnkqZqUl2lt/xkYHhTTZU+gesCd4gXivCbdHezabhk69K
Pc/sJaAUMEB57AYZgs31KmRPqwYkz3krah6Llx9A10tLi/TrSzqe6iV+1lUph4aT
PmC2rofbrvGonMWrxuWY9rp+3UzterPxP9uujrO+WWXDBFJ1rQrjLES2RYO77ysP
vxcM1GdbkYmKEzWI+RW0nncn54a3v6jRivtwiCMeiZHKM4W0cswIdHcDCZLmpW1U
zGrVhaBk7N8I2PFDyspT/vRHU8bgc12ta5oJl/hibXp4teZl19UvAt4i8AVOvQ2d
/fVDIv7rsGocFhnRcmWa107FrLwhNIyocB/axERX6+3afPJqokWAmkR+2yTMPQtN
pp+lGW+T0NGvHuspZXoTFgJxw04mwtGT51GZZpyH1nGgvzwwZuDK8mEz15OmRdhO
obPT2H7hZV+R2sLxJYzQGa/ZcMu2APDGY0kAbE0cHWavjwFK8XsyWyD7b7D96HlD
gFmZQAj/HjIARM0WHhfRgX4bMrfyxZqDf/9mvZLJiUsN7BBWqdbA6B3Ixlb1USsg
qKg0PS1SQDDl/CLzvn+v3mGMe3SlOSbCSxURYwWdoTUz2gQvN1pNwRW/vxpJ3Lj3
g1rLUnyBv3DuRee06Z9YZ0QzoS8wuWioqhwPkjFkVLT2zs6XkQz8ivEm2W9l4gBY
eZk3R67YEnvscfJ4qR1AHWACghVTuohyh1mJVhb1QDUQnWHhIKWCo1Ef91if2eXo
xcunxjYECpFhuh0rlPpd1Roob12OAjqcaXXw+dsh8SY8e8p6/Gm2qMW/evzjK5br
f4MbpNOGf8jr1qmi6g0Q6sDJoBubSc+RU5DtdAshhmH7aJ/YnIguCGyhgyNTCtOh
MF1xQwzHJhgt3zlVx7rNpgvQLp3uYUIPwqkFUCs6Ds8edf44JifgamMyiK6uwAt0
DLQ9hce//SqAaZ8SbmBpcQDOGWOnZLWy4omYGhCAeC12WYv0CDdsTsHaW0YR4gye
GQnn39ygf9UthoofkjtfINvKa60PWe/IT5eukuDTQERGOOdsaZ2LpEWauM2mQWut
CKrTG+tAJj+iO83l00LVYlmD6eVIe7cVnyhfNFnMNWB26U8RG1+wBwpSjEanL96A
czReXSudw+PVU/L1TfPCUZWUULR9iq9MFTNgN9aIGwgH0Gkbwf+hwoOU4a6lX0o+
ItLPqcUjjc/mh6cfQfMSDL3AniGp7/JGJeyXVBnMLWgAACPy3yL1jF438YfM4R5L
1RcOwXOEdt13PizCMPwL8WF38KyWy5UlWOkvNTZRaQdgL/SIcxGfeFu1n4EzCNRl
oeT+I29aNW/D/xclyoQkw+J4F9zGYmd7iEj6xdsafTFa/vriA+Hg8mq7dMO8P/3i
Q0cCW9zEJxZ2+hvuskBvEk7eOmRiXZcvVkvPhdvLUpjuErHjEdaoopZqB3FXQOKw
dnoerOdpkYtp49wCP9UVX9obmTd+pkgvD6wUeGyOJoAeZ4o40TvB4TvYWw/nbifS
Ssc33RgHoPqb4uTetnYkY/kBCY9LIHV4DH+UP6JPY9Lmwx8U+yE3yUR90QrTytG8
roCKDyjUw6dNx+rMgRqItwcnpRpeIaKb5p4Q+RwiVnxOk6tygV6KNXxO72HrmvNe
9dyeel6jTmMnlBOKUSMDc6RJRUppBPlZuHEXeEEu0B0QelnkUKlqei6uM1Q3ueIW
i5LKPmFDxvKvHGwQQbwv3v0SIwYB8a50cNIdl9exS+3Ez4BN7OspNpCKgK6mJTa+
D6zz9V2hoQOjqH9L2hGIJPS9uRcU8ZkD8dVcO7n0XG2GMUb16bQqNLl1FFf267t/
/EgU+ifqtcft7y3QPC+l3JJ1OCdMp5PO+vtAt6DGPTa92sruQtXDz57cNKkIDJrd
i/+UMP812mJsN7g4y4AdbnQAO3Xrj0/hAnI8Tk21+EJzXDyXAo2xdox85qfVhgL2
i84OmtoV3I5xORCXDZQTn2chsagZAaVaB64vsFsOBcY/2OInGuVGOHZ0GGhMKHxc
KwTmywZ3/o9+tCTCvrN4yyCg9op/Gc/Mep0qbWA0XZV1ti2QBTbKU+hX1ab4msF5
N7W5OXzVDYfjsbVQryG0Ot6G7bO4333bfx/GgeuNLvGurLFbUm8KlBC9Kt4d+IzU
guKWUbZADVJTF6eJsDDD7ETAWPQmFQ6Emw5z7Y27oWYdDMXqj1j4HaT9dh5Rj3bs
0v/qg7hhX+jkUJCMA2qKoj6ekiE0oDRvfZ4Cf8N5Q+UP03Vl/BTDgHPS1U8nH3Fs
YGR7M43e8Nq57/egqp5BwL/ZewAuSPC8ql5DBw3Y8Q8x44Ah7CDefejg0894+Eu0
cuio9h+2rMYp6RL55zYyj4vPpdPV8duSyC5PWgyuSvniO0UGu7/ReZdNP9rjpgxh
Fs0rN9kyF0kEhB4pi2q4AIg1RyrgVf4TB/a2seeeO3aLyLdSQykMPldHPFPhJzDD
wJwgjCAW1nCGPo6+Z13zpRSTtm2owgHuLpE4FlF4GREZPGMBbCcRw/yJ9gAjJeTr
S1TaSzOGj5DY9Gzn/81SNTqrabaWki8Zac1Ob0jSOQc0JpT9lkARBY/NxalJUENs
JgK7Y8ekOywSHINtRmGwA5TYp0u7Oj0czph2EyNcPzEGS4GmQkJ//J29maL5Brml
Te/vn5NB66zschp+29+M3uoJfajAFKmQ7tlNV6bM2L9poBY+7jSBrGt0x/4mt5wa
GRIUq8Z/GblL4w5Y550vS8fYXBSWlXjf7mVRWLFhBv79D0seJkTTasK+yo5+g7d3
rw6urTbshSS5+JyQZbZ4xGM9pOvTQg94GUs9Gyonn9JIuM6J94iqqE4l4/pKZzVI
kTwXXf7DWuWPhk2cTt/Md5ELNlR3nGZWOO5/rwHjhbvfGX8S0NjF1Xr8+dLH1cTK
G+/r7BvkiQgHNdlV2is9Q1lGkzFL+EvcuPyo9unqNf+AUggvlr/Kvmt7FJSfp4kQ
g9BodDAxotMyr6QpUMAcA6b/FZ5MWdWeBsrysbHe+H128wPELofdBXY3fV64N8IE
evWLPRao27YQ68IVB/GEvQg6Z22TZ5Or7IUaqpDlTDcA+fEQpqSvy9rJYVwLjwP9
OlImh91CDE6bfJDuofkBHTNE43PAxAuxLvpt4C/HnOcQ5Bm8oOojyxlcyuDFFpyM
6sv4cewh5eL31SwukoMXhubPOBE0aIPf7FnJ1cUunu9M8Mty4D6k3kEINiRo1yil
ne38ZsUZK4FPKeJhsKUUgqfv252jl5v4SB06PKlfeBnsPvkbLHDGJQPvzElsr4qe
RVSWoN+rSgSkimDj1RV7sVwMNYY/Hy+v3Wx0IudP4Np9pc2/TX0nOKPRNn9koSYk
Y+6KNN7jRuejbE/goZ8NuUbBPuvJcWxwWqEbqYsYGTXmDXsO1KAQ1V4yHn4GQZbz
ycPiuyeDCh8hGnQO1M2le1ihLsPE39rr+PSvE5N5nlw2JrM0dAgDYZxugThWdg90
+PNKapxxhSH5zJ0YuByrHVfD5nuUTASjp2Jn69IDkUFbuTvaBkuvw1jH8vQDKrXt
doDocfk1V6//+l+P8vOn8QVDTaL7jZxHpAj7t+w+wKEZD6FTF2S5c/eMYp/fWKfH
QuiaDLSDvJtUPJ4GF0ZjK5MuoRZqLgVNQvmb0CK28sxWw31XSXHoFz5+HPvMyiFG
0808GEyIAb9lEMRW3GHKtFMQLV4RxrXKY556N4udKG7OrW4ozG1mHKm8KzhZsomi
kp23lXepJNzTO8awh/KEKjW/i41h/7g0KuhZDKkP30zLEM+N2L0B86uOKkG3qRWQ
6khQNdKU4POw/H/KoDCyB69N50EaXiTa5ZLIWGQ/u5Oq7qh3HzWTdd1/w+v2AXdA
mNPTKnk1nbjY1sl8HyX2xktylw+jrEDqEj26wrrfRGjl1QQ6SKXutrZzItSDRj3G
I1owdHpzP8xPBsdNhRkCGrHmqgHrpdqZe8Xgsox9hWcSFpZjBfwAW0MsdEkDFqbW
49t93gaA5bGzeRVA+RcN9iVG0terCK5D9XFKgqWZ8FwFS6ovWw1DMzEqgy9PB7Bj
6XuL4gL0t/d8h6eKTXFcf++fmCK+IwNEBFgN8wfIyENELBgXUm6B3fXu1tT3f82g
qUgmJeNqfAs9UBY8u5HtmTGVAi1MBqmDM4Pk3tpecjRb226RiO1Rvo36Q5YUnsX2
aYrv+K1b9br2eO9TtR580nXSPgi5VKjyysIMJ1leAlZvL/uP55htuPdWzUh7oQC0
sySyXi2Gtx896nxz5wcAdqII+AQgIZ/7tAags/QkMf0Bokp/gsz/amHd18/PLgdL
f9GnyPTWziymItxqtmdcEqFT2Xgvmt+gW61ZTWOmC2CbDtnItHXpY7RixfDKit48
H56G4ZbFlVedUIVbRCQFyIUcORXSM+ZLYWG2swzTkHhKDYPKxxYbh0AGrr0FPORh
1+9GE6EAsVI/g4gADPpttKVNcCSRzJQ8Ppj8vvQ1/TR0ECQyLnTUex3uJRlEMfVa
dtvqeU3bvQ/AoZyJqll/mr6IF5IgN6+27o76uNYJhVO7x2pbr0wyRxdmMDv9A6W5
p1ajahPZuTJkMkSLrI7HwVOlkpDWQ++UMk5zrvZh3bkZAWkyOG3lShzViS6TbptX
QEFiAzZub24s7y52PTEU9d1nLS9c9bVrQsMpnruxzKSywpc3mQQVUH0nbTN/bDJU
bEjEAOlLoKNNXv7XoRUGn57MQCGpSzpuTEGC8CjTti/X12tMA0EKaeM2/vCZqHDW
P7sjwJ2Pfal3a+MndeGz6Kvh+hPbhk0hNsGSaZyW161iD1JtoFUawLcgXEZYGCQr
GQCQ03irKHLLOiVNg2CzBXqFIzyInz+73IHgAlEwZhEIJRn+iF9Yb0FqBbXu1zk3
qUNBM/PHwbeW5FGzaThAhXSvbT+EInSDLkHsHmrdXG2xwF2g0nzoGINHJJIGOShM
tX/eNlpC4d53NrsjVdGa8ZX1XRLnvgvV5p1HIFeqj8izgZXHjMHjJyZyBx9eqAPi
b9B8tGqZemiwo0zrIt9gz7JiY54b6MWNHbbA2PtQYCn4xdVY2AZ+rPRQFkeo3R2p
9nzdZahfpc4VunszG3bAr6a+2y7nfe21igJDXZ6t9c/lGSYuJmCh524ch7YKeioB
EOwfoD9FaHbwuZxL1x/eD6n85E5ZT7pNFZ1hd5qInWj1gt7Cjgp7YSxhfxXciOLV
ixKUu3P5C99UbTk0yKUWumkBpfGzYBpB5Ata/QEYaVlqoaas9BjLtqLPR8GpIfSO
+S3A+T/jO/DzVqEeMUHdTf/nL+iu8kxBCyqu40rHgbuwe3flwmDKqZv8U6OTu/w2
9Na+6eUcKlFwG4KMpxyQlwm3wwVvhtDP1onQE/GyWIAorKCX1Z8T6mruT0tjn6VZ
+3NO1Ik2XE4LZi3SWwBF9/cE2JTL1WyRPbrHcU5syJfeJPWIFlnRNfBlvWsw7IOh
X43FZH+ECHS/vcWSs6UnopzP6fmcze/h1vpn28l9gY4IzgRsnVV9YsHtfdnvtbNE
1i8AEMHh9VUT0YBPM7AkIWhzXLGLeHBYIPUbxkDW/oeb4JKhCQKO/Zab1WcNER1+
VQjKiwOGM0Xf6+Zx9NeYLa46RPCHO/1wm1aO6On0HdGqkKzNtPOrbxfFaRfCqIIm
YmOyOiAy0l1zzgll95MomfhW5iQLWMLtXdO2IkdgWKAXNxOmFSrE0mBI7CSx3ayn
gwHe1XWQ7IXpHXyAlB91j/SCwFB6XMGo5m/dkrGbj8P6KX0FdPhqlxx07ygZ7w5G
kss37GVY5LZskGUgNCBio4YYngf4qKqO/BwvGxQREACWjYIogber8fJq9o2eUs8R
KQrKSNfeE4nu/Urok0+xBygggyPCTb8Xm+JsL/dBXhfM/PWG5SxvkSjS9zymUDxQ
IziE9kxCE31E9hLdjpdzlPche+YhTE1qQpiPMmRgtPCxqVQEcH4rhoj5hbyitpIR
5cLvQni5/DEwEks8jlvLPBn3Dv4NDlDD8jNZgs+Ozh+WeFb7jvGs1wpFkLCJ5g9P
pPrePyRDJwsPN3IIOpa5BO8jij2dNfQkqdXcOwCpJbOnoWY1icCBkyYlDNZ8w/JO
div9rH0ZCKGj/LalD6s9ExAJwuiEQ1t9NlbGmOA9lPUUrh0d615vq1rpNhOG3MDm
0D5BnhkL6toyQau25Nfbe+ucSRMLDryFcVGDWoFN4NXdIvuugS26s46G+QeU7CYQ
YoeyAgCBtFDAdOldwUJqBGDIGIzUzeDN4i4Tj+3qC2rG0gsWLFrWAdrxGSvkgNW/
y1AyRL+CvrC8QgMsGxmuMrs3Kw6fCrlxPWf5z01P0hP9mKiZ0QPRyxb00pY+tMzN
2ZAR533bybunMUQvvZv3z3GAOqoJR5dQqy6SU9/in3y5Dm8s73rS8oR2fEjJBO8t
HgUD2GRVVsfLohbw8D32PsgotToJBVSmKCRDzRBX/6IYcGTCbF/wtsI7K77qJ1jv
C/jEZz9JH8vWwa1d0ZqSJWu2SOd3Ky0VC9g1/2ov1zyB7M9V4LYCaFMobLYeJMXW
fQ6OJT25ckMsGQTftG0GUCTwJYbuCr0q7QRYpcS2OAWQ9E7dZWbB4RcXGXH3NCtJ
RcGk2hUqYy1XzwM44Ps6J4c1/UaYWZf28KAvBhuahA3zAX76rf+YxnGVX21gSQle
e6hfYGWWbQHkesLc25XTHFKONsDF9xj6j1g3Fz+SVaNpoyScYrnWOB82TR+6nfPv
GME/IVI/NXxH7XD//bKZCebr5LwvzB1G9snAGyt5iix706PoVMObddXq+sMGVkIv
OEMm2Bg6brSGL2SJgB7+KBaD0TLNLZOf7hLYjrlmr2jJJUlvMRsuHQTeh+ftBcEV
I0elX9eI8tOwxKurhMLvWScOOIANA+E0soPAKoZRDAmSXFIq1avWGbG21ag0Sytz
1rfYns02udt/pFR/6mVVIwZ1JZgtmDZhBzwysaX8NV9n04qkJlR5yMOaoMzeaeMG
h1sANCyr395WGrfgln9VDnjA33sGaOjd372wQV4Vs67AhX9nV45mMI0gP9SKjwR/
L3GdJ/DNP26csKYFZEh2ZoCtc5ZcOEKJ+BEDfP4wkG+Rkv+g0qpIgbBoxJeTMMAt
KrTxXPO8RREMQ2THYx1iXycuxEKJB5zqQ24oKmbiG/yvtYqYJI0vdihb0akEE54F
YjUrsNESJmI7tPgdkBT7i1HECG6MhbkWJOZWr1n09UawAYWhjw0dklYwT5fF9VyS
n9L2cSTgtZqFIh6wo+vx16scqbdNw7lHi6LiVDK4uRQw+RyDx/5nPeCGLinEsq4Q
VsZAMv9Nbc8w7ZxFCswK+UOxJJBecRHQycuCDXaIpxSLq5FF+26F56S6QBs5a0Nx
u7fenxAzSwZ1wasCwRg3PwsdclyEQr62WsLn1lkjanLqZ9Enx0siPoQCZBuygfz3
85BmT5IYGLXcmeVqgItfKsLQGOHdNGtcmVf0m3olKGcc7QuUxnayFkbXhVzsafgB
pQPymkXlb2hUGuHCD/ADJUKPQ88veK695AutdRLRup/k7YeTYwyOCOfZ0qivVxp/
Y0MOptwUGV93Put5RByGhj3sQxN0eK5aUK0oTG59Zkorvk/rSFD/tct0UwEaUpyo
zVtWpDaJP+p/a7Cp3AkXJE6mPV4RXyRqsqIYQxSNLNWs1xMwcCjMy7AlgzP3mI9b
aKSxJMnkQx7qYv60U8pNQi4DweGHLSDcE3K10KdC3B7Bs66bSLeLfhvOV8fZs3E3
/w/AZ+p9kfLLU4uV6zduzJBHTegLmBC1KVnt6ncA7WfPugq4EnDa0ySbASnjDUnM
upgvBWZEYTycQYFGUAY1R3gkQGVlef5bhdlEbmBAOLKiNICqs1ZBzpsGej9aSxJS
gZ4LGFumpKY927TASRn/4FD5JjmtH/HUdLYU1ZLUyKFnZ1AYKNUpiIGl2mlxzxzh
7Ilnun5LvFYL5w0j7WRU2ho/xVYi6kw793Nv/o6vrHPpaTmlvJbeAOEF06Pt+XVt
o9ZlV1cwPnoIu+DzN/oJZ9bhA7iMpg4Aw2ZVJqMb4YFEbNaZ5lCFmKOY9a/t/T5z
UrMRLo4vpsVqtBZdPmkN4ioKp8PuOQIbMEgRnzUHE8cWg+IoTviVabW1j+m0Eope
TCRQDHBv9PpgHkqDs2zs8GpsynFqLuhlAzhDKT8R1SSnyjGoGLPYmfYIh8SrpQMq
UCWYvCg5B7UtkgBuGKrA1ZZh02p6c+KRCIHDBlS/MQpj2A/vkw3V84I7c1BtK0va
n2vd3bJOebMvvOcbNRIpuwpBXo57ryvOHqdr5kpEg2VHVrYbEY19w+R8koH8PEA+
UumWrIAVNmT6SPna9s4vMpGqFXFiPT0NTSuigfPyRcBwr3LWFP0ig6UAAOi94v72
SXKNZSoexn3q6fkQElHtVgmcVoPO5QNBVCLJdCpfZspueajiArCXKgTlhyaFca+Q
3NJn2aH+AyiC9tSeqRMjyl0FdJdENFqta/X/whiUCNwmS1cDqtyVMzodj2p8YzBd
rHoqQx/7P61txUr6hG/D6RGQwEbgnd+VOc1oqbH7S10xZOe4DzYDJYIiQF5jSPz4
d4bvtKLve5/9t9AYtFngO3lBUG//fRSObXUwWLYL8L4KExvePSm8xhSb0maSZH4P
riBgy5kk0N8dRErjYfUSElLFyo+eoi0kqBWJvQIk3b2XjISIPkuUgRV2grHBy9k/
JffAEFfC4uW2HGyQ5JAP77qk1iRVjgL1pZJeAKnLaoaPhWu3gT6LpAci12JSaGlo
rBnun1jJpFIGZoSM+X8bJT/hcPJG93pYEGfLsxGZn6UkE6/j7BGjglF32QrB3YGk
CR8rTX6A83bfTc4j9Qv9LWtvQE19il5iN96PG4PLsY0N7CnsSnegGjrpShuN4TsT
C7JsC5rVJvIXlL7iGuB5xYnkgDnpK8lxs/JOKjnLwxOO0XBeh20vNCo67f0VYp+k
hZ4cNz4bjYZLxErjseAswGhbYAKgJem1K02vUVANK4ZYCsYAiLCxcOgedEyCa7j2
AzomV2ysidYbkNb4WBtRqMDuxjRVFKMIm982ijJOLHnj1Nz56WKMBqZrhFuKKNCI
p7TGcW9PQx03pURz/deBsj8Qy57J6bdkwPN+hNlOIHV0VMf+0iTN+HrPIWIahE9D
w+2PebyaLNPeE3rnpriaCQVoSnZsZPOKpx30STtyN4Rf3NP+pukMIr4fzFNISJ5h
bVbtLQ6vzbZDtv3PSTDvijSEygxXqZzWm7NJ03wtzGmAsVASI/MAkGVq20hiDvLA
DSMlRt4o4QZmBDafiAvBgFZuv+7fkDJ6DeAwVLRuQr5UNygHuCeb/D4+6qw8+GG/
u9VGc841L7kxeci1ExMpYCmnqAIo5UQt3jg1gqI0LfkIXEoo2khBhqu5yOaYfdBT
UdEHd0UxgLolaFyrwPe1PxzDtv4iyEDFW9e5uYAB1gQa79JSKol1UYJGM0QTg/js
2deXn1ug6tsZ5BSA+pOCePo7rF2SEnZDxBku/dQ/Uj974ste2jPgobLJX3JqaSCq
d723PfeB94FcA1gKin2QbmXR3ayXXx9R1If96srCCiapx1IGrrl4jgyT40WILol5
amZ0R/Bqq6T2SAajsMzvJdmBThiKRm3SjGQ6+S9aAaMlyiJIEkPhhdTq5InDUYAg
Fd5egyw0aLOy/xTLfKmjl6May2ez+Mtd5Ryy2R2hW1M1R/bPF6t4kIOJWohB/KdG
o1f3bf/Ihl1o1bUbGZW3RWylGj1/Ah4ssjiLMZ25okVogPa0tw8/ygF+MH8CXYj3
nAo4dDU1WGxo2Cjc/SNTntNXv+PfiAXn0+uMYlzgd1g9J1+mUp++UajmyThHjpjA
xs8Xii9z6Zhd2zRl+5GwFmu7W1rKHQggZZtUYOkH7qBOUROEOo+ECgPDr0F0Vxvm
XFqggqZ/jrub/oJT77GKT8nNfOC2QXYbqzi2XWSp4hF02xc2YbyE87ollG6KSKso
Lati9dygiVzQSJyCN6hg7J32Pn8H0281hcVrcnQK/4YLHd+vZ/E9N3FtVF+Vv/uQ
14FHTOxhrQNzDYuxQAyLFeLu2Mp8PGb4tMgqMuDDT0CrifMsQFCArVM4X9J2v0Hx
Tnz0wCAkxdLBNRYaA4quxo29zCrMMrUqS2t79/DVsGlKMNCtJldoyIDGIGb6BqxA
3RLrcYaA9Cd/uuARz5BE6DXKRugNDoHGTrVD4pV9AApcvbvWq3OQLXGAEM5+9udn
zSRaUFEdbMOEbdRbO+O+3ug+Xg3kWPj8yrr8QhOw2s0z7YEGQR2nV2GqzwRnNm6J
deeqrpSQ8AbXtl3we3aFsH7kOevH2SkgMLhBOPb/1OeqneJzSALO3+7qoXic27xU
Co84pNOYJvubvcNIBGuJWCYzQPWW7yzqmQV0fXxSgXnvAkqpshMZDhFLoP0E09cS
8TPVQmiKXvWCC7koG/alA/a26fVv+mvH4LhAcBJKPoXtg6Gff4fki8ht2HpUf0B3
tmsbhiH1mVruI+6yV+ULuDyZ/MBdxZCX4u//oTi5nqodU5LRxRV0ht80jGe99xg1
mRHglT97JHXM0Ae2Ld4Kps+ACVB+amEIzc4ZdENaJyaT1UPVEzd+PtHvq4azfstc
OzEMZMRO2zXtwVf/kl9+FX5prhihDJqtEljDUiJYhMnZ0NAFMiynOnWj+VGz2TUE
o+Cf2U68WsrUY60g+nskUPmweAUW2n9fTrmGpGlvn6QVzq7PxkMtUyV88FrwydxW
C0U33N1IqaOEd5zQ1vyIPtISbhaYydd4zHuV1qMS1h+to/o38iJTf5XiV+yhJsBd
qxqrwZ4JmANlwQ0EH63xbZyllIYg01wMSAMIRt5yc3H6wosO3PtgLIAevZWeEUcL
F3RYrwd3Gpxr1YIDNPVlNHxURkyhSbjpLrgv8qj5VvhKllBOZuD0A3wjOuYG/VQZ
1RbwuFpsGbM8TizTZP6AEA/jpl+4ejBYadIOLBV+a++NK8Pm8c5BfEHX7Y/r0zrT
7/A/A0ZpAkAeUmAGK90MtLAdf6T7xWWKh68/GA3maOab7foZx4huN3+S7MwNjqQ1
MtTyyhuslUeXpgLjU/2EgOH6MEP8sQqitYwj/hCpmFJ/1H6u16IMF8M+86dHpFqG
9yosRmSZu/VxHaLFi4aT0mMYSi1oleRrgG3b+3YDekwFS3RFi3e0ZFFlUrphIxWu
NMvwrbQYz/iJYbMXJhJrH9+e7DrOKudrW7kn+JjTeqfNDRvk8fI+68wLHNibVYdU
IzYnPxO99dWvxUHTRziJxd0468Bem2wQSzdQr2hTfJdLI3GdJPK3RRZxAMOk1OVK
U8bi0TCgCoFRnN47sxjz4gDBoAWLpohar/V4Hq40XSDuyaWVf7FfZh0SwuJBDJVe
N1LjF3itzes3yNkOlx24AwHwrB/OaLwIFpIbpuNxWgS9dSnDSYrnBLpca8OFcfcb
pnkj2brBjTz43Mihv2gVmp3+9FpzMBFtfSv43lHPfYzwxubkETUCq3WPmCaiHjH5
nkyl1r1INqctpPnv2EVgt+LCMYrKMLqlBS3gGzxX04sOj1pJ2jVcHTxxTIsqphB7
teIfyblAn8FGecLCW2ZmEpwnQUgGWr0hrLHh55Br5ZX4LAcDyvk9ogG2Vs953XN5
qE7PVqIOzmH7lVoqurHFqeBwIvDU6gnEKyK8kOpSpLUjMmc81OSD7TkyE1A5raXp
mw3NOU1/GKXP6kyTqd6jSLdeJbevtC3v0n60rnkmCnwFnxLQ5Xi8qvtNPoiDYcqz
nxSMbh6bPDe8CnqMC/1SPkJMvTTmPwGce4PawkSg8Wd3He/LQMNjqI0STeWhccxc
Sm7b3VmE3yXXrlnOyeTLV2g4YXlm6+Er9iGC+2tdt7m4Q8qx++hNQ6QJTjVrsqWv
QvFgAhO8dIQ22I2IQVXD4yz2CxEspwN+F+muRpBMrCZcCnIGiF6UjIJ54Tce3x9E
drCxDqDrGDk1j2Y0AT3LEaoOLfn0Zarx+wBG+7RwwMUvFYvDj57dNqL7fdDLG72L
UUkxaxv+q4Z8CNgycs7no3c+nqZoM1egRcpRjJOdnduz5sB5iHVdr0GuG/jZGK3t
8jWTdi0q3QBZGeM68RtXfd+oElsQaAaLLlCuTxRw31kjH1nRRLmAsVQ0zvPo2E/h
uV3qdJ4tB79pkzTaUgxgIEaRzO0VPyv0ycG9PqoMVUQ3sraXgHzQfdgUa8Swz0o0
EDT1TWfZz4+3HhLLbCvdPXZm7GCtK8D0n1ob39P/Ydyd9DsEQwpUL4LMSuHwgP2B
0UsMy+lL1ywraex6Gzs551uNwdMLCLuh8o6GkxQTvp04aR6w5j0QU8HLt8aOtZqU
WKm5wBlsvAWF1tfywl0IUFv4lnqsDKriX54o5zq4k5oIOUJzWLIjtarYyjmP2pEZ
aBGU9NJY6U1LbWutjFSnL7gZPJNIhX4a7upCwK0NqFZkY+cpeoBYRclU0j2YK1ru
3XdpNMODdNm3V4z6ttIAC+dLHgytOya7uP1QS4DYEBXv8mmEs5eVXwqCWHsN7A9O
wN0gAR8p4qirxqyHNWW10h3ubum4Wg+OonY3jUL3CUYaC9RlRgwLi5E6uHwXKqR5
FE2C158ywXXjG90emEkbWneHmRKG6xp8Wt5Xz//ZyGVMI5zC0nlQSBp8O2qeANxh
dxoObKQgFi58Gqq/Nc5Jty66D/PMFarGyhYENoi+pprDgEMS5Fdg7Ek/xGLrrXOL
gm4mBgfpoojlhm7mDrpC/hQMdF9ieeu0YH6/Oeb3C6dhlrao6yMGXiD9nS6Gc9yZ
A3Z5sU0yXo72ET/QKHUTXSDF8Zc5Wa+Xdn6O4w8tfvYqW9JpryMQgVaJkSERlxyT
BIge5/eJTI2e6j9CwA6QyCogDt9PHXyWh3Ps/nomgo2LzXHSUYr51LRwnxq5IMPf
GmBYzFpeyZ5+9NI5UhcomRjuOm0uoXn1KRV0Do19Laa0ZL+rxdCLuoHbTdqYxtHi
kBm+uFO/w3lbdk8uHe4SaZ9doYRceI/wEKn5qP/N6ipcnAaUUlttnrvE5jcDZIs5
0rE6lj71M4u+o8hWNxMWL6Hm2sCDn1kmHc3/nVuRV9h10aujS8sgP4NArBICSC9+
9PUp1WU3onYIgVTdDZmntcW6vF5EYsrE+fMYqBv25m3MpW/pSzINO4RY9AcF2qrJ
aQ3kq6BXRUY7a2ae8eHkB6WOYms2M34R+JEnBEn0cPdfob3oQ3bORR100xF/bUDh
MJSPQrIg2MD+a9gdZtc2e2/v7f3OzVc7kZurWkkjVKIcxBZ7LkwzX/2OY8qzL18v
vdJAaeYiOa77lKfC/O/6yk471gwBc2TuklDUBSruIlMOUbdunzSn433f7T99VnEH
iqVwdRx2q0pCrmGgFiBgM95eKf/u2Uy7iliZvv8Fc9WApAP4jFVMm4t9VKTIaxWh
FmwjKeqDMi+r4qCYWiGKzRJ/ZLV3f/QJvkoUnI33MYxjettLKZ10VSgvpQGua5zm
OGzdhfYLgkNY1pKetHcCrhfRoQCIRv5xOeG5CJzbh14sOda2bqU7598UjPK+nZkl
lJUHjMwBoe1CDruXud/iEThgVGIKmYUOJIMqM8Ow2BqLopaOwjNkaLn5BAHD6Q1H
3TetCZMcenPoResVvg6VdTxbFt2VhlxfsRHNuRPiMk9il5gC9imJ2p/jSHX0RTIZ
+HQSfIhhdYKMzUMIwkJ6sV4jMyQ/IfNpNVv+ufXVSgG0sOaNDjGbSrFyhF35oMjo
9+OCwueNw2Af7u9g3MduvowoBcHA0XviAil+s7UIbP1eqeCrcyHjgfy9us3Z1oTP
KNCd8yxpQEp730RDjkWx6vRZaTuqmJUjGYJa5mPZsp5KDqtVdtEsbH5hid18Iqit
rnk66E29GpMUjLZ/179O5A==
`pragma protect end_protected
