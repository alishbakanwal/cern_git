// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:02:15 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
mobGcMWr87QHcL9ZRAby3+TQVa04ulirzvh9KqmIj6BpUwoYyxh5s3zHqWa9n4vF
jfqLVpzlDjjwMW13ZsmKlcM+z9lSHM5FWvINYwMHpblHm60lmROC4UaJ/FVkn3rC
4oAYBX3FsxQxkkU08NHdhE0E55WidgfSwIgCSLzmy4k=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 324336)
458557C+MXnpyqT0phq3c9s1iUiVtm1Pq/IAGzDz21R7lJxaBvNu40cNBFfuwf0Z
7d6BBwwpACCzYkIQH7FC4PyuAS5KafnDxbweywQ5YJpp5naBWbwYut//jf3HesNQ
dBb5yw7Vm82WxQd2mBYVwrxyg3A2vsIsYkuxlXyWzxU7iNHHhfyPq/BEeHkONRnM
evdrca2s7cHM2vjmJIwGQR3DatE9dtIjKu0wZVwF6UwAZbMo/IHLi2Nu9cSt/X8W
EJUNMXZGUXlXtES6dpfvOnIl4DVpema+47G64oc9EmqT7H1I/7ckA1GE8fW0Pf7z
jXc0pq3RYC0GxjxZAndIdxqM9feP4FP8a7WxuI1sB/wrO9UB19NGIbKES0xrdZXH
E1tB2aSbnZpobWxHMBXu10vfbMT0QMYrMdsMs28afyL4z1+c6I/JdTPjmlgUpvCB
9E2W38RuqjQ+qk3uB30Dz/i4qUcahAww9SU+DHxQLczZBfC1yJsSB5DA0u14Um9C
FxXuuHo8T10z+Zz/XtERQtPASa+lQI1cY8HRAyeEeievk1zzw8cotPYZaSH+uBM6
PJQ7QmUHshA7tUNQUbjbYZZuSnKi5GCoX4iLAocrQ6L4IPkwv4J4AghQlMG6Nz6c
3ILgSEM6uH4kf6W8ImAoO/i3pBFcwAc5zhA3OT0rwrmFcZ1Vr5f67EwcpIg/IXIm
fgm+1j5SOB6QrTfxYovhW4rUAX+CPnQcinloo4Xj9lLb/CSQTKWOKcW1PN87vzAj
s5j15U6tVQD4YhZ10MM2I7/durVCkqEYfvI7jhYXmU3wvQ6lg9dpTppTMkufrvVw
FN6OdfughcJ4VsVrUIZvG63M/Sez6nf2iON/gEcxuowGtB+GXpcwgoR9qwZ840CJ
JyUH+9NoR5iNSq7+JNCTYKd07qaN3vyPd2hmNipl9G0TDdfs9XYlrSwYSqgme91l
kEmsJWcIcc9UB+11rUtegdHTh1BnUw136/BfECzFm/4Cpjh/MuZSWvgfjtmsxefb
JWgU7HcvXz8G0Qzbr0Z2U6Goa7wTiG/HXmoD2TISRaVK4Snr4ERNocFo2q6oaZVR
cH8ck5jx1HwBzMKlr1qpmyZifi+ALGLv0ksG29ZSdwnoV3OhjKoisEPDe3l771u1
v+ikuOcbomj1EusODbp+pPTlY2tXAbNWW857zCY6RrWOK0c2B18qQcEnhhUR0Yg8
HNXEN5P7UBN03q7MCBFaKwE9Bv5XGu2kgX/zaxRcQ430utsOY4QFehqB3ZyWM2zc
gKSKkrNpn4GhJ5p9583H7dB96cNXQTEGLsVklorJ8RNqrlbPHgNMdXGkEmeZyp5x
livfhcKvKHA2zwSbCwpHTZJhN5u/S4X3+PO3sGGcd0jV2OhoibLnHJOEgYioJ6hK
eBlEs/GKoSFQ0OFzot4sAGaMX1Tp6X0zGOXvl2yIwifCfo4sQrqwLXmjrkeKjnXT
hmpYSfuNac4dOFPIvGLChKSyy/GCCcbjpdsTTtD5lhwCMzEY72R402OQF1jWSvAi
68v0Ax2WEmezpJF/ZDvdOS0HKTMt5uVrPFWtjcGvyASyhlEx3K8Fs/+RbBFUjJcU
a6EUih4UXGtZFToVa+oTVEiykWsuWz5mQHy4pO1s2pe07eon/5Ty/Aqcylip3iVd
rYXclykhpL30eqZJBbnnwmCTBQBVTGHgJpUpDhBu9e51F2d5tC4d+ttGMbxAozNK
2rLonTaRR+ZuF8flbPYMTgsFSBXRe5HOWBKdNjmmmEH54p04nM/jRFmUPMq+Dl2x
O2m2uuZr+HCg5kCE7oSWy3S31iHSqYg2FqYKDzcT4Lkw31s3GNhibqLyUzUU60Rb
9VcTN0Ac15WfBtVpBB05JCibh2LPp6rlGuOAvkeROY4M4oOmXrWMKnhi6Ai4ZhS4
sj0BjuOSIpLY0iIZJ/2Xw9n26e7MAEocREjK6PdCbQC/kbqdbrT6TngVDuiHQGPW
86LYJNorVSviSVJAIHCKKAFgpfNkWAgxW4UOrIIO1inCL4CfWJzrL2U3NFS0rHME
vcHv9Y9gWoJIY5sPYcRx7CNx67SD+a8m95lBYacgwYzzf5Adaf0CwmL2T7KeCM29
NVwp/nGXMr9Dwf9phHP8+BhhbE5TtV/xyPpdn7kzh++rmR32y6RGZ9nNvKPLzN4D
dXj3mTPm3UufMgxafFLUsLJSrKfr1zudUw9V/L/Rg4MPvCKABRgkoAQIIaYe32Wx
qBzrXEzN22pJzORzoGmZRa0DclKHipVHHkqk/sezaYz5oXIosFMXSDdYosTG/zCY
8VqqnoyqGbNiYnFukeXF8x+lr4i39fMSGvPUL5zKvZr6Whe+m1hBLBbJjX57gBD4
mjSN08b/0tRhoOev4ZvS89Lp4A8T0OIkf6sYj1huTvIVHJ28TJny0LNT2EKR5Y0O
RdG8z05pRUpNUMSeHxg254RtA5UlYp7kuihdTvaM8PGFxi2nAe2ds/GqF+48YRNh
yjAcVTVAiwIr3MUHg7/kncbHyFkoyvmtpzsHPNSDLNjTrKIoTDObRzuRUabBGk9C
6QDohZAQkaumTI/FVOw4QWDj3TlVMCTmeEJdlSM/nq+j84PIaiUrWqYxeUsMUxAB
kGu19Su16mmUK6JhDsimgmdv9Qt1kQ9MYuIAUN1oyocu+YX9ufqAKv/tkgobs32u
WbyRaRRfYc7p8WoU9gwB7wW5xokPx6jGKZUBocVH8K8PFp7GUt/iyduwvFejFZAv
8JRYVX1tfwX+FIQl/pD5SmnT+o+zoLy/TGOZUmlf7JJi2nzfaGYotpV0l1KiBA29
BWZ7ZtxqeUU1rbTQpBPvypRHTYe4acwKkaDLxvsWT+R0VgqrFMftL5oixxO6gqju
eFY5wlh6AtEsipSRrL1spMzXitKhxza5CCfcPK41C492v8Ng/lzsHiaw8jSNoBXJ
uDfZEtmwTytU5rergDWuRNlAeoaFOlTwtWpn4B1SU+AJXLz9r+f0V2BQ/OC1zQXP
4vjsYPMgVf4RGFseKdaP5jBYRPHeC7ABL8HX9jOziMc1YLliN4kUicqb7dLN695o
SsfdANIhdEgbLO0BZz6qHDfrpmY66O4tZWIMtAsXQnHhTPfPzaRVY0WObdNL7EL8
Lntvn4boSUgsgln6lSzy8rPYU7FlHWzd4bz38e4m5fgJeN0MRHhJkEcQMvRZ7Fi5
1twux2m5Tdg0NfJ28P0s14OKfS762W54MbBkDtVlxzpL7qn0doignN+Jd1x/mb2s
WhtHgCkg1m9N7QQJxAK4jQXJ9OKpFNfM6fkKZOWkYZw3IeDa5nKoaMdbUazNmyer
TUBHjv0EzTIGot5y66s6Hrgnk3Pq13V1b1exNwAOUXDu2yipQNINAL/WJnNa4WP4
n8cjgw0RzGJfkSXgu2Z1Sox4rXLhIYR94MvT4gDj856U391KktXtjJdMEv8LRoip
jjITCuQP03fetenY0UScjNhMd9v/s1nETsEtSr6OCmTUzYuDX8MT1UvYtX5158Je
ni90iFg6COewfWF1Lm4FnEM/tXtl57gi3/v2RcVbxUjPbf0Em29d+beR1Mg6rXgP
2Ah3EBHWidvA/JTxtOdVReq4bi9y9o5vLLpdHY5O7HbQlhxwRDvE/KLj9sN/fdd7
zTODmwwYt5JKUz90QaFp6gai1RpUkDEusp1kV5Ds/m4BdV60VXLooNdLYfk9x+FJ
OYxFulynt54LnHYJ7zliNNmzlE1k1bHjNDjjwUtn1oUvCdUwcWsJN90RdVL2p+hG
N1OK0FDA+b441S7BM+vgOz24aIyaV7hfldEqXYEttc43WsP7pDfWgyALOo2KtqIf
GOSPLf+Dw57+O7JmHEJI5/ogvpzczjCp7cDPrI56jxkqjmGYfarmngYHbGKSng38
I6lGODu6XokxEzRheTjdUF8UvuJClBiPZvdNLPPK7M2qWS2cO09wqnDefHhHmuNR
vsow5jcy4q74KfldNCOf/owA8dtFqt6fut6bLFS9vloWBzCZsPevxhREHYv18zkg
8azMQctnOS0d1kqdlZzNRJs4BaudE6uHeaKeobzbcb09NbaRDUYrIlTmMQCDAqZs
VmY7CtLwA4P5FzF7qX/XtMPIVFifLP1o7DudAjqLihED5FagMKtNXlnDSuEAWHF6
AMEQsI7e4CtZTJjkdM3XshG17n1Z/aebA1M6ND0y+HSQfj2XOFxaaQFThaL36HiN
xYQHmEjOyNISJOeSwE+Jw4Sx20HgB7ZaAwf6sRBpuESed6GuvQsaTixoMDf6DLe8
7UCDhn0ncetP9PfjD5hWXiZihkWLDN0quj2h8f1jxIXzWSad+BoMx5Uut/pQwonh
+aUw0Z743hZNFUNlckvjLZm3jzDiZGFL7NdW5tTS+a1c7tvkdBWTRLkq2y46YTi3
aY656h9JxJNMBr7HkISdAGnm8wMDhJlE/z/IEHxP8M8kJ8N61KrEhGDQRW6j473V
BuUqD+hvomOYs3nygWF8DvXUR6qudlrR2Qqbw09CFVNGWyqWgvrAqe5HY1F917lS
laqiV0SvR5mcEq65qdGwWsqnkUZly/XZ/+C/gH0415xVFVsg1bm3D7uXaqVw2S9j
GI1qJdN4r4ImUoAZ2M11WkEfKS23WKO3J3EcK5W/eZ5Hph9pj5svHsr7jFEFZoZ2
ZQT9y2cmY1IUPrLMOfiviT6tJP4uDld0W6ybBTXout1gwwYkJhI6vhn3756qDHXy
W40zpFLh3fbBn7PetQx4mD8VeL+QuZXJIHiSdNrTpCGIfOZPCTqd+CA0+ug2BOj9
l8z0EJFlkm6t+R/jx6VswUYgOAPHIdNGvxTV2Oiwv6sLraMJsj+O8VyDscWxa/8G
tJ2WDBBlKoZAiXeFAlcuhsKRt8JD3+oWd4EDv4qehnXPfGn968W8QsDyTouqpmgC
L+VkTZHm4fgviuovlQa68Cle1Ht5PROH0DWG6StmWRI+YFHuExz+N9D3ufCMNcN6
4YC9dCdIVxbfhtZ+64ybZgQfibkTnDxOwFA6qiZnZ9hFrPBPvp7h8YW4Ajzz8U7p
CzHhWIrOt05XtAp98oG6/J17NZBwuuv15+jLm4G5LmASH+HyThRGVlzo1sqfXrhf
ybOEodtFivi8mp/jUxYij7/E7muB3nknL9C/79HfK8G0wfgLuhXidJkj/7S78UZX
+6igmiIvQ0THaIY4Me72/OfrrjDyy77OwtSQYvejSBjapY0RFX5hI8lsCIIJIL97
KICaDiEBeX/D7QYOUkYdjfehwivSDrxJ3jldzBuKimujbJejeIiIyaaorUp1y13T
95wMu6+r/354UkBtFbqg1bLmxHpi3ISlafigRHCiNMSFPZY8irOXBb3XJvlBqGTd
npXgnazjNaHKi2KR7fzJOZnHtpb60i0fP9tne5CETAobcWGrKf0/du7crJr0Vnlf
LZDUu7zmj0ePFXbtnsNN/jjGzt0Fc4oZgP1UTiz6COIwjDjvr0pAtLEIreMfgz9q
m6z+D2ecahS4JM6+SEK+LpMEhd3/1xq+25HXaDoh/AAuyoagkR9Q77ijTlYflFG0
ES4pApct1N39z8QE1SiKpQXcuTlUhWZDGKWlvt6Mdot76npYQ7ZMuWeGP6ZyfPwc
Gr9jmOrPiPNAycCYnVNcE+GH4pbNo+uCisEO9ga7YDLiTJXumGP0FN5UXGkk75xF
r4OzLqcIDabQ8PtATKAYIavJO7Rt4migMJIcsjpDo+ge/14vBNyjQxgoJF08BpMi
awVZqiU5kDr+zPcumpedDmCmNz8ZGkn0tf1843SKa4NnZLSJrjJQ68TGLYXowJ3A
56tR1afADx8BTwNc/nbaa3ep7GzWX7jHzcxewrWpkVTDrOtqZ8UVlTT1NidQIYO2
zsJeDIOKYiiRKdclYpMzkMp3lEvHNysjhKrE357FAI5khWZnzkfPVQKphjFtlbjk
6r1qKQhmeR8fXHTuSgosjqMc2d+6jK5heqyD9T3hVIgHvNVHVdaQB3Nv5HVHgrfd
e9Ig2/BsayyPDzfgEO3cer26P2+4uz7Ucbmrn8HyiwVfogvzP0ylFUQ2qzPH0zRz
Ul7W85utR+e0ai2BPhwQB6VwBapfXimFkMw3qFj4E7s0qWzpqJJ+kMkKAhRJ6dot
gnyyM39FumXNK87w9sAWUQV/Grl6SL2uWwPZ3hO5TUR2Nz0T+xZDEbq4XOGlKtLX
T8pGJMaLIcyDrTnjawvVXmcjjzbnFpUyP0jrJ6kdhveuBSMPamKUOLdvpTb9YIrx
XFBYHGPoVtcT5BTzZNUlysvC0dmUUuHDz4EpJSJVerdAqwMKLqDjoWNBGTFmTo7F
FG23t+2kl+RcFwrSaP4jn7XxwsvW5sL0Nua/xkeJZwhKo9dwbOM05o62EhEpBLV+
JbKQIKc5c6vnt5sRtIXM49T8tBfwjSjBplubEnqKrOV9O5rdPLPVgbQCSXKTM4g2
ptbT3Fi1G7F+iyzs2L6G/SuT/72YTg3dEK3zFOIPKV0T8vs59FB341NelcbTCHR3
dxn58Itv+FMWEg+/XT3jgpPWmp4WicUOQJ6MD9ZKsJH8XESxIM7lcz/IRYUXl0Mn
O9TqN0QQbX/0T+2cAZ4zjthiwHXBaP7/LrILrD3K+//DAB/DphXPJSBXrlx5UeNS
IjTApTKF5UUxyAj/bBQZG+XLdQSvJ9uQzIGBivp87CYGE27b+t3O3NHEeQ0lVNgc
I+hTROZFeDCZPWCkFmp7nprQ8ybc0WDnJhxR9GGl9fcdk5RCW7Wi2H+MDEHjWDKT
3epnmyjMqWd3VwS9AwewZ196Q4ZXvQLsPbJL+4DhkD/sFZUP6LsmNMsfW2Q3FH3H
gWtAP1saiqtfDyw9zpN2oewGaPEBaSsjVhjB4gVGOLxZ/Bmibb2Qtt8yqXEuzZj+
Y3ebb7oWAIYTcdaY8UR5n3BI3/X4Ne9A+7wTYLLXTmWdpruvXgRGw5zfC8YSIDAY
0dLe6s4WI+ti7hXMX1cK9dMBNf4GwcaVX2fxR74nv0OcwF9uujtU6tIJqNKGWY9I
XK3sM2zO6HJ/xjINZ3m3Qhd2W6xwobghToq0n8GZ5L21P2nEO0McNzyCiqp3yJls
M7bGJ8TR0tJJgQfr19xtoszg536n56EusZ3H0WZbLtTXkqFf/xloKOwUIcmCAj1m
6I2//JXK/nmEkQzkcGTmdPbz/NtfDgp99y1BJndjtpBnJzew3uiN4Lj95tQX5kO5
mItqq6h0y7wuLXl14LDwwXub/jsvReGvs/K8B7VoLWNxD2JiOtUIrdy+rwgutk/3
gtHaA3U/H9km2yaqkVofi34VTgcjRTLfKHlIJ6UnWbBYs6mLIbtDiNLQI+dRyLsL
zRdkds3LuAGgjzkjwIPl6dCcg8ilUzNZ0Z6Lwu9zpFS7SxhuL+TrPC82brS+Sm/3
6jfSyF90al5dhrLK376VEdF4GusPL/VBKGZtN4Js30UDHYEO6d7aJLIGRFZY2BQq
uJ2JZPTocn3FzqgmM/ZQPo9rrKNC8ap6h7f7LBAbqHEIeKH5EtRnp2h5f6ELeKht
eWuj+oRqOFeEMXB1Y9vNgPhnwd6RxPXU+/wPMwa+R3fNqqhdoPbeoKxywyZAQ/SP
ylKLoxvxkGu7So1cJy7dSekWqFsr/MqAp8AOI7Pzb+SN1DfXmFQFAC2B3Kvr42Ul
5wUOMNgX0RkluR0vBqYh49BncIdlYmY/m8Sd1GIANGUiKaxj7HFk04hoeedg5h/K
tUjc+0xOkWrwBFa/GAMUQIkFMuOpmszZ6UuKsMh1EykHcroY2d2qshwa90CuuTRM
9mduNzYTES/iZ+4/ISJvuduArF68akUWonCIFd4Xh2Pwsu6XZ3ANFUTNLTyL4ZP/
JETQ93X1l907aUef+UQVcMbT8kG0ylhmDJUjHLlOYSSR+JTKbqc1N6WYm+y1cmz0
YnP3kw+7U0lFFiyoNbEVduq1tDc7fIo5ew8Hpxbr3tPbbs7OMvp28AP927m3JFff
t3GHTcY5hdznqK1OWBaz/VoQ7SUpBp3QkIZ2eJc3V5F4tMLpTfu6EwIMV1oMLifv
JcLdZd8QCiCsEUYhmJ/u8gBMyf1PANONJtV4r5W4hYsk7u2LGhQLFuWHBiKIYXHH
zELVT3D1wNKpw/OvzCS1xUnZgmoApIDgK8URT8CrlX/MCT2jujyWWofxJt2FKy4D
pJowAnDJam/6sQJfROUjdQeUMeKog3IzPP5zy3NzytImtDsR3ukz7yOWbZQEbjLS
LkETdo00ZbpQG+NX67n0JMbEO1PX1HUdIQadyNJLhDzEMx4y9pVYy+h7nXmBxSsx
RMK1tkx/mWHIY5iVvhcjyBqZuR6dTqY+SufXfYCMfqxyfJCgMM+h7v7cLV5Zw7Z3
FqK454wdaJo4dZVatg866umS9c0krFjeN5CH9CJCGV2rDp0oaxt8lvbOfbURlCeR
174b50x3Bu/sc6exYbtFaFDH7TQrmqgEE1OsL1sOcLUvLdxoien/XjJGIGUSjZWt
G+Cca4/GtvR1DbgwIORPaEzjVofNfAac6SZcLBtrDygwNpiglUEgi9zuFB9X4UD5
ylNiSs6pIsEOVzlRejO02Xw5AKu5qA23fXMYPABFVHz7tWjZ5uwRy5O1aHGzybfC
d0/hVtb6diNsbRh8UDIGGRgIgUI1BGOjd5thSYFY+Oyw1u4MGbOT5o+Hu8B5K1gg
BZRqL2CylTvACcYePbm/cuuzj2vGLJspfIP/K8jtc+phxtOgzk5gv4MW3sVX1gPI
t2xhuXchc1GcPLGctyUqv8KpCAF9vrYA/dy7OD9e37GDxxeKuKsJgr5wNX8vD9z6
J4G8d3oG+jeAde0qSkVu7GQx5l6BabWp2TSqitEfmmv9KeBRKtYDKXln3MJHM1Cb
qI2H3slicLv1VWa4yWSfZyPDFkzj4o7EVxnjsQoMG9XHD7Y/UoLAuZl49mI4zaUy
4rVMLiFVyvIpfZreT/Gt9NJ1B9G8Qt94u0o2TPxD5rAo7PqIepGRQsJt4w1zp7Od
n99B0hLr0C2z8XWcyYTk/ZuKWM6RNIax3qBStDzp4RKLCO3SxyxnV40+45/Trw6u
emQZYSBa5YgnihvYXtM4lkLifbj4eQRHPM3na7FWzlD8BbX+Ze/LJ9JfKdAsxXOv
cHUfGjGrKEZOldfU6Sg8Pe9JsDUUUbdOXJZugQaMKwy9ICCpXbv4+69Y8IwrXXS4
wbZOE9J0mhipehngHJ/9UFHLnth4teEDudA4oKlzyXo4tNBpQusU3Yg2ESsxRRK+
d4HA2skPO0jwLxSKy0BMpx5xSWX10CH9JFLihNb/OYbGTi443bDINhmdZ2oyJNaI
IR07C6rxMrI/uFOToVVCXeQ/ripEa4Xp3XPDm/A+WkoJyDQxRACJQ+UPX9sJOJ6a
KrI9aBQbEdgknUp07kx3I5mNqk1tfo8XZTz6ffaj6b1ZvJcetHa85Wit4CGDjswu
AAQ1R60A3LlT216MXyy++jpw5ezM+KLarbpDtSM2C7mQRgeqYz2T0NMtfllvaI10
KcWJiB2XVtJuoAp6CS19amw8RPlvoHXHrmOyPSpp3mUXuQh60diew4FCuowIQCOU
MLFO0Z1/cfyBWYdX52VeOXfYZcOME4b7oCYTuhvGzQOaGKPzElLbVuges3j/h1M1
/hgDcKCO+/QIUTPdLMGyTpYna7eSd0kwU5L7ZzsU7IG8qQC2Na4pwflki2Div7Kw
varqj5p281WNsrzXAXlRVOLd71U5wnZKuE59Xe9vmAaWmNrGwSbLrX6LAlGMAnqZ
W38xXZlpDc0UKzdL0Hi+zyz8S0Ie6gtopPNZvgJq+G68YOcNPsgOWI4KjfzglRil
xYjZsr8TmWHGt9hfMolq0plTU7lCeIn2Iun5UNLpqDen25movfBBTFSYLA+ZXhAX
cF7UzyEK3l8Hg6n0dHt+Qba1PXQ9LZNVFUJwATSss9dqGDVSg2PPDNi9NkKv44jF
6JMOkoiHQpnyIVd6wgt6i0qHeSdnnVDrGKb5okbOrNjc0cIYs8nmOoCrlDXyJyxE
urWBeAXYWaJeQP+/cFhfTi/qVSH2V9l70ofpwo6b/MAcYiFm9chrcN0q8dHDy8/S
gsaTVumfEcgFP2tdgiy6lwiZzywHlxrnOVoaQbx85DJnawfFfHgzVl2UWKnw2mOP
GJqu75VdKFCKJDLGpI4AkKXEge1nBEt6zQ33gyuQOuZWuI/uBNn1SVU3mdin1KVK
NnvgXQSskM9gxQpm6bTQoOGb0JczStZXlzfud1Ra3q9Q5Y5NLf6yLy/h7KAsoqE4
LIoMv04w/eWky81LDz1H2aBN+AL6CUcDQv6OWiSzlfOMvhLhu8IMjgtaAegQihGY
IEiQoiQ/vPLrZyfxohQS83bqn0gagHETsFgwHuf1OpnlNMoIiyvef1Okxd47WneN
9l8uapVuJJUIGzT432MHKk6T9bVpy3Q3WbJngnoK4XuAuVRfOURNiI1uJbITYIPG
/G2g3/U+4USGdXomC+rJiZpYvRNUbcDbsKmwbBns2OVmV++hdJN1K/txaqJ1HzKP
eciyo9YesaPZ2emRX7Go73pFOQOmS7/w4ZYuQSR5tJppO+ipmiE8P08Jn1GYhorc
1H1kCw3g6DkFwpyGoUZRJHX4xyKDsOgCVY5ZEwoGVIIEtBIzenH9+Dx4zJEOjMpB
yWa1UkldCV2mmvx2HQB+dx6PLwlaf70PJfXe1OfWrno5TqF6iKsv4AiTBp4XJznE
q/g5Zi497fXvs4c4s+lVwsQ9WvrfShDCwEV/ZiPhn3LlTM68ziLvpZEQw4/0EeYs
GCaNXIFjA14P4dxbz0Mjkxov+vSbVbHk9ICCByn50paXSXzezQCOUp0Z0k8fMYg9
sYnGhK5NYCPCohpYU9N/xhmD1wcudiFmrN73vKZRhy06o9hOT6jusjBRm+CrZOjU
0KZ/4lVpHEngH5WwYjLtbTzbp9sOS7HZyOwnCViVD0Sax7jtYDUX/vzbCssmNvBU
EI/QEIaoilPxprsdqr+opTan1ahI0b86tYm5RYWIXEmRMHIUaQd4sr2lm3uGJlYQ
1ECkjFlP37nbcLd/smEeGdeEuhnC1+eu5uIopdPfRTHJCN7Hrgq0tUKvz/Gfpjzl
Sa2Lym3n5CiBapK8NfJCCI9Ua5gXPx+jvz4RWXen2Mt6wf0Gm8jhSF5WQ8kYcLLy
pol9u2MNzAKo+tg4VOw43AyzXCOungxCR/K0p2Ju7ZTovZeEak8r3G8v9ZKlU4CV
P7KMVReFfZsAMdsEcreGLvQGFa+WwzQOgfPhfsdSstICN57XTzvi7Ubk1piGSIqH
ISW/qGclxz4wlCx2YjvKk8jevB1i4MCa4FKjwzY3WwzqFoB3sm/vPK8PXUrb4ArJ
Tyq1Hi76hGD5FEteuoqE2/YBLMbTVDrUKSoktnKF8TYQ3w/Q6y2Imz7IOISa9TlI
N0nvd90E/XkhEElgMNoQ2V1HVx6PYPqgvUmX6ixj4A5dn7lXAEf1+FnfmZZlVCMe
W+pG7kG9f2avjYL2GmicOocqBvK+rHVoqLv7it260U4Z87dZNjYcGwN39IJhfS6G
FXqFR8m9tf1dox3bWtokWJTKSMoj46mw/sKAFLSj2dX0jFWCSDboJk8eH2Wnj8vR
n4+vPqM5NlOucSdh1JOy6qjngpGay7QH+cktCmMz1vGeJTOOzaoti9w4cvuATfnz
gFioL0Wr77llZoteeGxaG+84XxYyo15thX1rKzoARvTr0lSL2+ljzn43+Ve/UcDK
3jiQapgyFJNRjRvwgwRqc9v4gEL1fHM5K0XyoQo7T+Ju0TP83nhhak/O3ZAzKk7P
4KXoTcmDhwPbhwm606umrnKlsRsiEGuJTjpdtb8KF9wP70pbknI6MGUGsc75Tv7j
YzpJFOnkzuqNRhdNpZz+WS3M/jfOaqsmcIYbxRov7avuhm2i9R/hKmGpwemel7e0
CLoKxqtr67GqUOVqzoJEVE8vyJ7a2c6xZoEAKGhhf+xWJqZIZH+D0Za+Yx2g01fn
irY0IOh8YBbttfy/waEbRQ/7u0cX2FNXj2B5oR7f/+XVYhXwOopp8gPQajh49Yro
qxBKVHywwYgPdsTxQbNlWfyUpbsSM+XjfLBLwNtC+L60nYJe0kUnmCG9I8lSyppP
UyuYeoTgxTpZlnzrMoJ8ixfNkFVqIVSbBW/a45FSJhSsbOH0nsWPXsKv1V6I+6gm
+9SKQe9a7jpKKJC4llgOoCzB3MOWHFj7Si54E7H27KeggTPrBisSLvuVKGmmCnbU
DF1WYiNJDqDSUUu3FWuOgTCO9TnnVLweCGvHz4FN8kie7deMa5MTQ/qLkwKi0oJB
/9emtPoLxhDbveLqOa8EDVQVhRTH1lbkPXWvE+8PuNuNDtVy6lDYXSZt7HLqEiot
2Wc+NglXDRl63QbH/087bIvogAAA3YRmiWwToRcrnFL5Bsg24zvHliJ65hYQETq0
DORRpjrdPwgCZxugZTF2Ornz5DsiFmmmUoqr8sEQY9cP7KTvZzaJwW8Guz89heLd
UjFOIfhvj1Eocw/pb+yXcH4dJ6IdQ3c57B8UsfIYe0IZblNQ97yXABugRjwkybpD
WWXpSXBeiqzBje4FibEyY+734jKIvC2WEvHDtJpJbrReY/gwG9ZyZVlcBTS5TMKU
dX6nYWevkCgeRmHFqx8Y8oQzP/7Uk6BmK2hHWAo62wEfS21nqjAZTuRRcQDravdE
cL+yVk2QmBlLOHY6QAa4pg0pxCHk3Blw2J6RhKbKg3HYcZenvsW0MxDIxgZMvpwj
ozEiByO/iylhurb34kdC6Lfkrc3I4xarkCNOxg/zyXWALYU9h5IFjpsanuFcIzYo
UA+9dX6lU0bwGu2F2+TiYjlaGNan2KCD7qE8Tv95ioP6/Y8BbsX+jaIQu+0qXQCI
CafCDDzECynV5YqxjN1OV/jd2G1cdHuJoR+CeFYnT5e5IPjPfGALWPHqHYYvMz1+
d6GbwVBbY4sfGQ04sY3YVv/HCbOUpYed5En8L1rQmkC/Rf/IL/UyhE/q5+YOJ+Ys
C6JDGz1cEvourgk6Iit0jP1HZ+DAu0S1MX/7UAkHs0oMT58XDu/pap8VuFdSeI4y
dWskuLraO9Z3eY05qIsnQ8Bw/NC+gfTxUodT6VTHuVUV7hR5TwgFgTahfnPQZs5H
zfw0wMYIU6vK4z4GweEOybo4JOjJEHtLzwAscma7Z6YinJMEuTJ3ir40u05/6i6g
ybjaUdhp34Hw1U04BsRN6Dv1mZOQGWO0Gu2J8ksGFYzqCcIj6VOjh2CVOZuJM9gB
ZI1ExVtiONViK4fJZBhSuDrWWNbZgfQXVmXs/tHdHCEyxoYPf4bnbx7uGYX0Q2MP
7hpqUQ+N0F4u9U0Vf9dXpDMaYzxwSRFc01oNxScw9HSNv3x8gl5h3yY3hCeQ3ZS0
mXxaJaWwCptX/vpStv6IQAcSI8DCVA2A69crrFAUeirvry9QXr7K93j2S13y5MsW
d+a6S8JCRvhGFFSzYZK8RA3Yw5M4/A1szLKRXCAsGqZIibLpVlzjIKsaZ05xP8WV
kkAfaa2Ch3a/mENUnwEtU07pVBEUff1vJc12EJT/eNpe6Hb8IGIg6NXQjNxeeNZQ
Km1acHZi0hdpG/Ax3QxhXQB1Mh2W3imCXymjQyxv+RUETTkenEcUt+ru74VMsQx+
LvDJV80T+2whHOIHxrZ6yP1cvi59a2QuAuV9H+0N0VXBsCTObpwGiHwVXF0y0wSN
p/5pR1j+iCXZKBc551siWAJPD8E6eUH3z4QMeHARGXtR5x1LOclsyJ+abEhxOSeI
JbiDkPYAr/sUoi8ZHedAYoxIfA/BQL1Bj0oIs4djaJbilqKRtHn1HcmHlVIuWTyW
TzZTXXospzCN1MtEkJ5z4GfPq8cMEPvEFVqJOXkpWs+9MIRLDZUaV9IxgMj+8p0t
5Fq6Mh/myOXWDuWblUpREesGyZwCLfNyHaWLasxYutsiZSBiJ5G/9erEWARyKiy7
V6aV7/b4jy3XtoSnxYZN++6I3PPYMSAZCR9GpRlxy8I7RVDXRTf47WaiYIDYUJbK
3m5UqRxU6zBmPYlyw1AOkWA47aRDJ4+crxo1A421bzIYmPn92h1ePh5NxPjaZwfj
FdB1tkQXm3aneyoi41zRBqUQ5ivbbZpYsrbuUl18GkW0otjyy7Lf4J23B+zoTyPB
qgjwJnyx0nmtqybRtPq2dAXK0PuMYfBCWOvHEnGSvcpfKIQjEV1SDCU5iJTNSOrk
Gptjnf+8D/X8D+s0m7wKDZB+kaqtbcDVHIIEfiA1L9vGhCWlBrkfyttwMEJUxhy7
4vc1Td9+ih0IhCFPsAMpUb/btWElSKVzu7LS6xEo+6GRkCU2qTlXkV3rew2A9EiX
nB1pwGok4B76IKaH2g9EKsoAbwtP4eHtOrONCHSHSsk5c1OkJRRrW0xrOHJyTS0l
ZknYyihEe5hNGKMp2PsHhxhswGotHE3yTfB8VfUu+nl20tZq/AJgAJby0fU72NdC
pI89oHe7jx9avENU6TRcjMvafji+/hJk6ktC3MSWHHuBLFXTfw1iHBdY/NFyBAMc
tmMu4Y3FlMxoZtsMfeMPoWYDhRVKYGaXboghVBuA7gpb/yt26IY2kxHxKJjaCbXo
v81SxfFTmPnKzijmJMBAiN7bZKeQWT6LJQTagRQpq9lIdK+hA4pKH5utTb8X83nd
03mvgk3GuFVWN6+nS+0TFXWza+gZNhAArBo5Jt/AC2kCj5e2ztTvXWWSDQCkwxjz
9fjr/0tvPvejCSC6DOUP5SD/29B9GSAnxt3LZjUvgcUpjgNGdqs4XLv2vxrXV/0p
nVSlYxpIiZlbLhVZ/qYak8cyvdZ8bS0JRliTUXupb4nCTUKSERUWWvJYXJO2nYD7
4esH1uhRAisdUXWIzuRPj8Ed7o6+YLcJVe91pndDvowm6TPfit+3RwTuPqBfNMUc
cQk1p3xKwYhaf6ovgdrH69721MTHXjRlaTSws9IkCjZ/g1SuSgRCHoNf16UdA1+g
lqdiqSP80l7gfhpeYZAvpAJI0FtrhACWJhYQrV/vvqV228w2iF4KJwvTs/dAS52o
Xu213R7Rz8zP0ZdlCROyb7DgogguqIcVYBEvkGFSbHyqWHUhIm15wswQpVajchK3
OBYN1bNnVsme8UmPGJFxmsE2UbW85Zv88f70QLFdXyP8wMh6jTrUKp7yIR9ikRRD
marLWFpCwXd2OUOdw4PWCGs9oKuPzqeuxS1GE3doCOfzUJscavFc7H1w8SB82Z8N
EcQim6aruTOoihC9sLgVhPGbs4DuUhNdJMGnoxQEu74B4zVKJ9USrKzgWhj+hUq/
josncA/kQ+wE+bAIprcO8VLfxOpNwilEDW8YJmLu5B3OAtPOZOfhdA1nRzfXHQ0b
F241fTJRxc9xvgLvHXG1eR5MiE6qiK0k1prREL8E/O2Yl6h6JTh1ltTXX6JbvQkS
N+DuxorbANfYvkVNaPf+fGnWZCATY5ydRjoxxong/62YsBJT0NtnzNowtkurGMjt
0GxxLeiwdOVOmfLgSeBL8cnRfc4pkQm9eANBe8kUPw4QiEOdGF/MmKV226OyJkzw
qraZieXK+0R/PFZutjVL8XFmqDx2VKhOcHUNJrO/NLSDgvnd7N068LUqhT5ahf/H
xKmOYBQgu0085C7hQKeLYaV68GISDBYUr9HHEkdoUH9xEPGSq8oxOp1sT5NOdJmN
8kco8x+KoQZCX1VYkx+4whhX6g14YheD7mGLqocIskgX+miQDHSQyPLfKZWtGuF0
Ld8jRiyMezgnQdxGph4qO1XHlJ4w4WqDyM5Q8Y1izOGGLcbUddSvs+xJOLRgmQLH
1Ozbm0wiSIGRcbgt8i57gNRUophWu3sVuj6T2a0ItwJ2g6KVL404mqpETb2lkdQJ
G8Pd2AliteX2eEWxYHpCPf8cTauyk4DMlz+e7cNHPfiMh7zhUeoI3fUAq1vvaCjp
g671I+oGN13r0YOtwOdxUGVJp4wA7IaAHwAbpWszsUMTQdwqFewuwXdhXvwm4uOT
gzgU7Et9LzwQR7OoqCN7usVkrIwvDd58BcunFqNe4v72gBBcPgYxQNEiRPB8Fqe5
biB5ZGeBiCfpTUmUs+KBsl4tiJhiHPVZSIbZdpGV1wNdzPXxY9MfIzCeabGTXbYh
pXkZnPvPKGWTF7I/Yh+ENM5KAkCMq6r54pNh7tC0qDYrd5/3NUY4SYZZqCRK6q4D
xeljfbrC0DsEYOFv0T5U+kNjM5RiWOQWqPJi7smIeTEeDbk8xqLM9ywcQL3DvR6b
U+NVFPaL775jjCQGLOOWOb7MIc+tA1OqvWQE1ZGV0iU66izPELO5nAG4mZVaDlSQ
3aoAzpsJVtTgjauNns4WfjI4CIP1X4pEdIa0bGO9GQbhXsmj8GLq6NBHCpCfqswA
4opnbzKkwQUV5u8gtfoGm9MybMNxFB096jXvO1iVW+PqCN/L9NbX4OAjrYiQ9KKg
ROaIUcucdTiuf2vQ//e52E9OtbZk/p4cgIbLt7CA9rXqoUScUY2mtQxCqFTfMP3q
1evKNkBEKxGp0ABnpNKj6oS0Gro34PIlNYLlqYm5jbY4BBR9AqPU2jRRcdD27ljT
wlz2kG2yZNUIAf+lSe7KKnXstykWDS0ONgg/QB0aLuDXT5DJz1m5fHlKJKsl7EEB
9qy3aFLlVU1Z0Qw1l2NciYgl1SS40s1LBaL3HgzZubwrc0TeyB4nYFRwS5ODdfHh
qCpSGfjifQ4iUcKg+oW7eL9QHZvljM1lQS8TWIDGYgHGwcpxhpNtPBBbSXQiX0xW
2So/nPY8FDeUn5DSpHAhnO82qxVWfHUw002ki45tDg96bGpTpUzL7fjvXx23HWCw
bemFeNKlquIi1cJcYbk5apd7SkgTIZ69rESGbhPM2xXlwAhpyHlbREjK1yamEpa9
NY+4lS1WlpRu2Q7kPcQD/1oLfu549AEyh5HPRjS31aQgEXACICrr6SEXkgFLobgV
qrRSgXC+F13bLYTczWFSIwlOz8kY+TX9+74DrFKFXUtiTwHW8+vswhHhw+pjvKNV
kJCS2+cbFDu9B924X9vbrvK693tGJ3TKYX9QkwNe2sdcPmW+dr2OSuaPclPEFQbT
Tt5KJSWXTlk0UT5WaVxNvyobBOOHueh0267y07ktyhOS0au7Kj4P2RVmJBIgYsYI
DupvQPU/ePSjf+IG3VPGE3ehsYSEB3wty8nSF9pQHsG3dDAk8rTrgi2aKTz2Brso
ngFcdrEEAzalQWdVYNX1R37PCYiGvSHR4nQWzn4X/KCshbDfk3P2E7QpHyaF8agI
SGc6d5WGznQA5rhE1P5CArUMg/Ya/5fmiz6dLkKYBufxYReC+777yM+uObQyL0bn
x/zCK//+jc4bRQvUwvp4iRXM2B4/Ya/p9uqOuuNf2lBg3Ft53ZLJLIM2emkLdDJF
pk5FqhLPzoJ02MxsGw3RLdDKXuO1fk1jCtkb5zmtgH7cO1uEyTeg6JPrfZM5h1sl
w0B5E0uBn9/VxPGfz/+lByJVvPpctdLWLtTNgfOUfmxXjCMeeN2Z66PepEL4KEfg
GCx769LbCERPcJTTHmyJDsU68328Ugy+5izjkZT+L5vDQrQW62WQTYVHGFgVdwyi
rBT1VdKjZBspkWxEukp8BjL5B8tzSrdTsBl46al61Kr/ppiSMpYkav1FuJj3LRoi
8I0QcSW0vbEfmop9rYxu5lPBSavFlWK02TAjHof8PRjV+l4xO3nFAURCVx+tj28b
kLbGGoqZ27yVWEbbmZ5Ml8iYF9oVUBw5WAUI3H3Fy5n5Nz/oA1bWBWwUdN5gXXIF
rm2d7MMbbenhTObZTvOsqPBdkgKB4eEqGHNKcwX1ojV6SvWzHqgMue/cCjP0Pvr2
9omehJ9HyJiNU/8yidwO7Eg4HqdcFNEIXt+DVGDkZ4cJJXpB4x2A7lJpDiOo/JdG
jkvZGp2Ypq+ZGKt9OCmG3yF238t8U2S+yKXZH/sYZ1spBZu0ICLC8DGKhRg7VM3R
v6rgA5povISLAJLBgX4DbVW31BJVdPZFQclBD3FCOyRYlSpg6gdiVr1ux86nGNt8
xdTtYCalbdNKstS4XpmK4dGXkqkaoYhQgyFAhoSI3m9rRgMiIuRAeN/kwCood2UP
e0CMeAJ0usJBCswIU9ZbWjE7KMOV5QX9JrCAFfHUwk8zB/fxy7jm0zAKpot7pQyR
0aFmLR+WV480C5PWVaGOQyfc5oD2ConjbvwR/O/JVBCAoiYCly/2jYgMcI8biT5R
UJhNfaQddAhoyrm1bRBITNmuDCc/VtxIsRTTfq9xmLYm2EVa8bHTi4Mio56ZX/qF
fIdcpNu7T/59hNoNdaO1BhXVRgot6R5xXe+aV2DLBBGL1OqcAHMDBtEogjeR71wn
F4cW2KmX1QD1yxMVqjIUDyotptsVddKTGYfMT9kEadEBQXj53693S5XGTBdkPkCd
tUNJAT95MsSaQTGnK1B39hcLVhSZYFfb2s9z+RqRPlPv7/k3B8Py6Wx/Jq3fBHqZ
167nzUTFF3D/p6DVJsqR5ie/SWlHM4G9mLVL9WomPhpFD0rSDxBr+dnFi0il23k0
ycwKrhoh6rhvuPm2qKRznA2TcLabcUlTbZ4c6ryRoNmQqQONWWjPM5B2ydOPbtWg
uvvb6sitzv+w2lqPwpdpD5hKeURFiCuh4xfr2vAPdDx1jNlKfxlvQLdK6kapSL4n
DD8sBEs+eF7bqm0PKQIfpqbMt4LMDd6WmESS26WB+waFnN4+pAOcN56MkuaUTB+j
VwhXKhT7wDG4qzjyBTdU2qn8DVJG5/8vgLcBclK4CGtbqivUmCCucZGasheKr8Eh
YoPvJUs9Rt9fT7Xrw6y35OYmTl5OlwceTopkxbKtM02OdHvKmWojwAQllkmYKM8p
ooUCHKyth/GwTbJMTQZsGX8PZqIQY/fPJZDNE5zgxdDLe/QWMrovtDiMqVmbbyU7
mg3D1CxsULZugXhEMfioXYJ4SHDNrhdzfD6SXDK4+OLUimqVuAKHblky/gFrCxk0
DsEJO0H8xssRuv/2Y5Lvx9FVjcIMaTWkfTdRiIG1r1k8wOnsd080liAQjw7jB1DQ
OwFsLMjcW6QWyxhMjCmbDRBKMVMtWCXO2FQQEZQ+nFzLJsWnAwqaG66BzCjA511/
z5SStkE2BPV1lCi05KAe5VjMxg/MAANBWW0t2MLnRZZTSrPijEzXlLcyuDe+oXWB
dQduKqwrSNZuv+/Qolf6GvgWvdZot+74vMcv7XwKoZT9N/e289JW2uTsCGLW6DEC
GZbzgq3mNhA/m3bXaScKVVXe+13RBh3gY9TTOyljew7ZjrKQ5A2HVoH9h+0WmLI8
vjYSEv60iFdAj515AryJdK4PTYIIwCdWs7uoLyy8bvRjNp5XWr7SJTI3EFDZsaAX
2WMcv223cSB8/Sl3i7pvNdSwL2aAKWEuKid8w7ETo42LXPnAvGV2+97sfqenPYi6
f0HLyM6lQ0qOL635Sl+0Unne+hl21zA/+HBE3rtxoEdDceJ1/cMGz3UY3NON8Yc5
kaJh7MgipkPMEeZXMOVYDNQHjeh0h0fqebReVLA0meRCumU3x9KUK/8nS/GjSvU2
ods4HEGHxDUInQfMkLfVAku1mW3PdYWFWolr/xmpveQDUQfbMkHrt0TEffNHA6xy
TIOw7xyt/ldx7G5byMEYQRFoqB7VFyz0Gj+K0oDhYf6ZjgBh3AdgX8OVc2G27Sfo
/INeaDa8E5mlETciHbvsGdWmv7wRMyqVoayxMGlE5xNiOF+tuOluJ+sft3vh4xNe
BYfHhPAVaWJUC4J8S0wV8CFyNb8CRSUrez/1F6Qm5mBn+2f9iLV8vhYHQiMEFNh1
xwPubhTRNG4HCPfVI5c6nQ76fW5VC0cWRsttf+Df6YNZUBMnJRwNyigmnbHGJHrI
vUcyvh85Gd6l7wA18WKY8WeVI78FtXv8rOzWDoJQPkvfpPWtxLtgEqZsun9E4eMI
xAx8Rf/0U727Yj5t+zc49l6aO8im7/Xj33rQ1crPg10WPXMh0VNOYctraWjvuOEP
bJ/5OKgNGLmfsiByLk4FMcCYROsmvNX4XGy4EqT9V38pTSgYiP1pFDrHQ6y3TXMd
CIV/Ft+lEhB2EF7T6b0iTTYN8CkPmH4CjiIXPywEQ/RaX4UL0723CZl8vuXwjjOW
v01woajGDVqT42ly7x9C+KaVIx9p7gz3tuLZWL4NwfGImVjZbD4hR+5UQobtI9f8
emVh2JwnSBjbV9r0I0L9wAy8vmTKuvaem1Zqeog6FIy8/irmJfQ6d5sLSMYm7g/2
NuExuuoRdH0wwc2hssAepUp+z8G1exnXR3Zv/aidaEJI6ZkdK3EWNMuQ+Kpo1UKy
nGI0Ip0xcmB1HLZ7KZmGdmfNI2tInDozDT983Z0jSGUfEYgAhO51JZtpg0dDdDPM
KvfiM84sSNQk3+dXFl2oKXv7hsHH913SOHwrGOFNtopmdeweGNu5oeL9q3M9hvvi
cnUSiXonVPy/Jf0OEM1089J3cD53QzpKc2xD1OIRyPVA7x7RUo7txXCWxaCykzcZ
/aLjVzruJQg7c7Soq9FxsCXfL6b3t4T3SXIJWy1Ak0/7q+4Tad+CAb2KRnJqsfnG
4ttd8YOQlTDvJiqRrLZ+MV28zu+xokgyU4Mf3yEOtzzkiQOdP9GPz9oUoyVr8uH9
V4gxGMW73EnLK1GovwZTpRTQTU6fMtoFghtaxKBN35U9LlJtgdiCY3rjX5L+UqgQ
ruRqLCwJc2c6dFAzqK83ZS8ygOKIXd1cZBXmvW741gCe7WsyEwWdO5mPzehUSISG
ZID/QqXgJf9fl8oPp0Ft+wLuIhUhXUYzXq7/B/qpThzW37zj0ESz1tDsmHQ8VNcp
9A2iqA1WRqnTIi7b6sMoT2d4pm2r2pLdfdzYDCdhIqvvEhAdOLOny8M/vTkUcF/r
CWkchlnXHbscNBGfAHicjWHv+nO7I8T8DeUElAgghkKAdlNfEnl4+aeoYeeNJEb2
enFY6PTPJa4sjCe+aC0wzRAPXCw0y/ku+wNJvpESvzhnsAAtAkUb1fYYSzb2nUoV
6aBdC/PdCB/j4GdlfNTCL7URd1YgPAJPr/rrQhR+DYMzsb34bS8TNWFOMYwYTKYK
nEsVagKEbXrukUZs8Up5qjct1LOZofD/l1J++uPV0YY/QrkQ6KiEVqtI84ZhOY1Q
iLIzHP6+ynpMiERYUbaEjIkZAyb6t9Oj431LPbYjphHE83ZAECdcf3/RoDN663SJ
hanGYJUNVukr9kehfyhku3nEhZnDQIcjlLZm5SGPq9rInnU4g9unIXeWRPpj9u4J
TpWmJV51WhmAFue+VQdOfZC6guFDhN289DSbf+EJpMp7x+IvBsSawi+YqKiMzS+b
VqJ0NsP18OW4b3/zKPHw2PA2Evg7Wa7HXKDHX3V1pqNFqAoVlpUpTxO6zLDwLDmP
wCyHNGZBlJ4Vuh8xLS4wAJEpUSFBsx4ZKgVx6lalGl47NsFFBn+b+BZCNRMAhhcx
ZjLE5oXsO6JZDzDZTLe9ZeiQxcQglq0gDhyDQUcx9gD4Cx/zmiyuT6/msUTXAjdv
MacG30W2eXR8GM9aBr8DU2OXt0SDxmhMwpGLStVnWhmF7uWl/bvjB2IKqCbyoQOA
Z529ghu+t3YeQf2RF5ndFY9r2fsADu8D+KTT9rhnGWvmYADz7f9c3+RLY8ssSYFu
WDtK0n0cUJz2qKb4g60J+kCJClq76F198q1GCRNBuboMXn/P7eAMeE7kOuL8yTEQ
WZ4ckD4CX/BIlHd0TojfkeiEMRr5kUXjGBEuVFawjfx43LCCpzWMoqN56DQrqzPg
9s3HWs3vWmJEA0jGkTCpUD1L6aowMcVE+RFmjrnZI8Gudg6XHaxbejAe9BHsZel6
DEe9XlDwpmCcxIwKwZfDqPlqYu+KfRjG+IOfZajI4p9vGGjUHqcHwIkrLJ9lq1TB
RCZe3OlvSzWAMR2UU9sB8I0dD+QNh+lp/PYCiJAD8KHmYIXdr43h1oTC1exkZyBs
bTSV95fp8jokzRS4+UTbOUY06dv9+i92uGRKpBKfxX0DWEOaxW2JihxTWuttQrsz
8zQRrDgwGsbjaBMe9zCHtfzTMPbA/J/HJoqaqO8P76qluF4LU5s5tZ21PAIDZqJ3
U54GqlOR8YL8IwmZbFHEJZShINOMAm3G1MgWRf7SmTErnDFnOn4kqFPxXN6EGhTa
To0hf2JOt6ZzwPVJNsF//94vpd9bR/uauUgGrKhiQoByFBJxBjkyKXxVEn5Ue1j9
WNfXaJlFxV4nMxiFbAsFEXN6wMUKus9ogacGzKkEccLMPlkodOocfn/Vf1TgA9/T
P5cKgbS0BbKGGnPUoM8vc4nUzSKkHQFuFNXggonBzT8fdaOpJIpm/fyVqjZV3/tf
djPygL7vIGcuzWbCfqQoEJp5aIDOSBjj9LmkkSa6ePq9lS+/LBo8EN5BI0b2yvH5
00nOhCltrUSMwhk0Gcg4vORUY1K5QnLgPBd7/zN1MvppOI0qbAWx9xuDMHZNAaC5
Ycd4NVgiSAhTcnS7zqupfUl791jQs8vBnEJmu6Wl7FaOKShh6zn/ZetyuYQtei0C
LE6Fyvh50LmfjHU2yH8+V0cftIQhfFmvtgsyd8cVA0zENTleGF1XsrxQrxUVdi46
jO1e/s8vUY8zhcIlK97TIhUYuAmGKYztnHWnUL48Mj257/wlXOPgo6EWcgNt33GB
9WzPK+dEt/Q41zIqaNkTe9JxOcMmSuzgxmT/dqWjn8rjGQ0zhpIafpkC3GGPFhva
sRmsYqbTXDBseA9ZZ1seqX+KfEGoSK6/4NLkWat0LN2+CO3pX1YERJuabWEfD+rP
8XcTswF6L7EbyWdAPG9aJuaRDihx68ylNXleN/QX79gQtiTDu91Qcgk5O18RSxAs
Jz0somWNZHiCveYl8AarZieyppAV1RQKdCCn8xdIpj2nSXQfAjft/VvZKLUWmgox
2dfONVataeTn2dJmH+P7C7rRTkyYl1Rpx7zV2MengEeOlwt4RbKDQ6hoa7m9Uylb
yeKkqdqTRTdBVqUCe2wlrEjhVZX/2RgSurxUsqKu7bPW8z6I31BaKP5e6S5A8m8V
heZ44+q+hEwy3+D8inaFB1e7WFPMqA7rDWLeBvFl9r3WN5T6yLJ1evn50+HDX7WT
1lgShDO/TjI1L7/8ux5pfuCq0jDIhxXKltE2qiCeW13vltdMpe54x5RVt2Rd2ARc
QYPwpumdPPWF25AQquH4zGKWLDv0lhv+oddE7eOyV8HouFBRNP2XK/JhSH0rwEg/
IQyQGHQoWyUD5qRhNUMFLwI7Rq18XgpmgWXARQ5ctKNKnXHCZwLki0AIr0nQTHjr
PuUxqYdi352JGwHQkU00H2Gx16cJxHWgQyKd0ARJSh4Cq4qRMhL2j9mk6/KGzqLE
Ees+gqjOWNJ7JIq9Joa2ij1J5o0VjwCWSMSpH/wo+4+lpYqHKZ9V6MhzKt3azk33
xNwu943ehLYQFXs4i+jOWwBWVv818+/eae2wcr1DFXkr15jwovpiiOKJ8Y1DMznL
tEbK7K+ZUuiBUgcdJheLN1OlkWN9/RN4uDxAry5ekgkjVRx+yNzUaeiqwAhRb0U3
TKDeNUMsehpgGHdgtkj6e8HnYzvWMSl4uHLU49F+r/Qy4Lv5DJ5KsLzDOAEXx3/w
iFWn6ycJGLQ3GT99HRjLAljJYcpZqmUi/gASbOtbNp+naL0P9GCUPz54trWFSLmE
JjZEfYhp3v9h86bFIKtTEIZYtm04DvrE6Bu3vGXowytTxX9ssbC9MuNIFxOORpqI
9VEH+D/c8TqX3jvGPg88uAorK5M1W5WpbfeROuAiCYTnSf7De1xELJaNeXKMXPB+
qvEclgWRXsIEP0w7uZc6a2e+ccvRE/HkAs+xvQYKXbkLk1laeVvT9r7RDTw5U81X
VZqXZ10i3EhUXADbbhq4/aV92G+ump4T1JxCoD0nC9mMy6B1GE4NLyZYly8rScSp
xGlXnUHE8N3MdgFF2/IAPT1PG8YCoQmNZZ0BEhjtXeKUYA3P/dtJXuFfCFLEGHnb
BpCZz6zWX50TQWHi+j9j1j2aeFfTlQ/pMqE1uYd8rpsgUHYUmV9jCrPfwaCq6RAz
KDMQjcI4l4cGm+sxcjDLIyUpnVBmEdjhoNQ+67W7oNG66XuOIKMUC1V/y3qY5+8A
glyJVpU5vrqM1r+BtIchX/KYt8lqwiNGhVkYnh5S0nS1qjZ+vxQi1LPykwiiDGXb
A7PoC+91xj0mKbpwlNJeoCZBWHoGgb1ZJ477cAZcNNy1MRF3gsTWaIm7+1y1Fb9Z
rsCsSLRxVrd/vumPjTrpBz7RGsqv7KdJRQtML0nQ6HEbixUPmRuT5YpLZRZTgnTb
QCS2vV1APJS/dbeKYIBQ7NV3uf7EeJ7o5vBWkT3FOpvdtyxm3qwQa9DOUOl9Cnkh
LA96ImO8H508VQT0XxIi6qc7CN31Ixs8VpfzdyJPP9JdOO+jrsBZHKgwQFGBHoPM
v2kBx3V4f/pfsUCspT6AWx/T3lRPsSCeQOs+2CcYxTI5pkGMDpJV9VMYhnlRwCDM
E2FA+rCasEqVHkWmYAJoqPI0nbWgVtaNvyQ8ZAB+JN2H4zqNlZGaRBkpEgByqTLw
lPrhnVM+nYQo77XiNu9L3phtSt1AU8D832ViPV2eiN65VLTYTtdqMrNEDatQ3tpz
zaqQwvxWnV4HZp7VSBc7nVAzRhWzUZ7i5hc8aaDjc/A0oSCqpferTy7FTZueVFzC
aG818nGo96jxLSD6vzH8BUmSRGB0x3bJlQwqkr5gATLR7oUftT89cxVGPbCWz/MB
u60ZWYzJVurUt57mJtnWdPhcAOsdaL53pT2SHvdyo5HV82yftzOwR1hD7QoKbV9Q
Ed7AqYg3Rkbh8H6GAao/D4ufKwa1G7gpeuBMdhUYKpRRxR9Ar2UMkCNvUtgENXIY
iTM/ZCyXH+1PoUUoxq/BCwO72mgRupMsLuSNYUCYNH7M7zxj3twoJ2Z+ZovVLTYX
jH7f6Pn6z7DjdEnPbHmIWGY0xESO4eODy5N38FqW+xPmq02WKe6VZ0t3i98gNqOT
PKectzUDC46T8cLDJxo0xk9JxqBgQiSgg6cWAsOHtpQBQIVORbYb0DjGss6HloLK
06d5xBBcHzAWPSwUxUXzhiGa0zHo+4NKWMV47WZP4Y5h0QsQN+YVL9afbs5IFyMw
am952sllNqZGCMHefKG+6xo8zRm52n5yejY/dHpQWgFCD1uLFF0FSNmH+4nkzuE3
2szKpFG8h5Lc0V6JcVVIv9LY1i2+mKJ4qWYaUFzmDqHiJzGlDfHIz20NPw7IsMJS
nnQZeJ70OvHNGSmC21Cj7yceec9gnuOPw5WJ5ePQbrAIMhMqDzvPMGZthi/EZMW3
njWV4Uyh7EUFghoL0KyZW9nz8D3rvejKUe2xIQD/VctkCVF2fuet3gSD/UgYL5/4
FabGFNE5oUjq7MTo57NQ1d09i8/7IPmLFwOD7XUcPui2xCMHgmpfE0fenw5G0xgH
6h7nuNwGUpeCp26QHULlVtt6NfwmCqw0qI9xsR8/8TJxAR9C94kJfiqko37L60uA
zRkudzqYIHtv1pzhpnlKPYwHBZ5BUBBfxDcI3SG8ff3w8iENDOXmj+3ZVg1AYiBW
bHzKrWsAkJLUixYdkpDTr7ai+CwNVpovcMYxdtSLzPOTahfoJGc+lShDHTFyqsVT
nWLtMn7Jg3Zu0M/g8L+d2oItz4iEiHVUi+lVqURlLoLHMKfqqedpS3i/Pzqhi8XI
lDHkP+xbFOHWYu36K2kiy10/2ljWNVezYSqJdk50TJrXboD/UXBbqyt5D0weEE4x
QnDHPnfjcvTGucwa7J3HfxUh2G5hnbYSohvSsnSEUL1lbvvPL3HvXoZAjBxZ6cGP
a4UPacMfoPCWYrKglEBqXAdvVKaGDU/f2GRL3TckCovGu4j2LxKNZ4DQuBawcyXl
n5v2SUjCuD6ABmOETlCtN38uJP3H2jN/dWJRakeK7+DZXv/WKcIzYBIGN+VC4Bm8
aEWZ8mlWDdworVq2bJLIVcIQUbFkDybwaxbn5olMGrXUy0LHCCPK2X92jGlQB6AI
VAvjynIC9rU7+G3Sfkkg6Oc3VrjZIjBIV24q+1OW8hSK5Gdq4HJrTqyxfRSbM35M
IbWYBJj0Mo3UeYV1KODXXEKcBYuNtNJYQl2gq6PR7VLmyFEdVttabJdiFw3Hq0IH
Us6UW3aviPWtGBVcE7+EA53UAikTW43+/aiAyDRD7G89UIXdRfDBQjtlKUAr2IB3
3irHxf9kMkofsOeUCeyHTJyOE9QUzSJRFGVaM+6m41S2Jc7Twl/wY2bBqit0IqYu
vNqGkBfiJ6xYhkB844q1lE34E4bpXl/+O6wp1oxZ/05V+8Jpq2C+P2BI6SfIJL5J
4uOyyEdTpERzw+T0EWBMGYkOMG8Yxkbsq+bHFv3q50CtKT3GbPZTe/Im6bwSZIDg
fyaatolNemCwU/xcgLGbKkvr2re3ZYdSSIivx9SSS612k9SD+UIb+NWrA1UMvpxg
7EXZScVhBwzx/r5WcwYTYpTMI2e0tGNRYtHfQwfmPPiJjBNMNeONBnBMHSXj32U1
z0BXfUqfr6io5Xy2bBgOHUdevfQMIqGS5lPFCUODIzO0fWgN+FS1/t6NCy2OrnBh
22KPoPwhYFGPByPLMIIVirfyPwE3CpwBpjT7iYzMw8G7JwH2JcUjvebqmP1SUDfu
b+NeJPkNxgX+09hL+2KPx8tmo+cauptNPwEwBvUPW3L/mGTLI6BnvrfAw6Ih9aFb
lcn7S9hkd3XmDyTjDgkJPDaDUtDmKbvnR6ibkXC6+hTlrM1tS/STv878V0MipL9T
UwXmhX40ak6aCzeKO8iwMjzTQIK9NQC9tt7l3pYu05rG0Z2lsemwRyQKOFppwEPE
wLXMdNlv/SlWo75iFQcwGHTq1EwV9C9qF8lBhR+2GLcEYwxDSN/laTKPVTE4oME4
C/TUzQWKKAfjsUJUNHDpL0eeDgVFw0gj1AHM17XFI4T7c2eM9K2UpmqGjDr3vj+q
icPn2E0HQbfzW4ZtmJK7wuQONfE59S+QksEftBJoK448gMKtvUbSgxIep5jMMnnm
G14ZChsTXJv4+kqH27TBHUSGRjTIVV28puc2OAbghxD/fRC5NCb20Z5SAqiafZW2
XyEINaO5Pim3fNtGCvPHs2fkVV8n/k3/cAwpPQ53BdVzEN97PFcwJzjNvZV+P4A7
M4KEdms984zN+y2nHPTACN69KLeTDHC8+bJ7C6H1xTqWAAynce02eryiU4T7h7cn
42MhYyv93HRZG/9RM4PYY7yfNs2Jnd1PmFxVuIdY+3xHWMFKvkSSxWGKR6xoLJlY
bTs79z/1e/jKdgUEbzzOJ8GXMp/tYDmJCIc50rPZ6THkHyDHg47dBifweJ3cMbiK
kXFhgb/1jQ3BbeoXWcNZ5M1O9gY3lQeWXSLXpT2dROXjAex/+zcH4xRhPgQi/aRs
5cBi3x+1hxW71OgRtDslIel8tlkNOzO0rW0NWnQG4BY3oH9g0et8pvbt33a/ghn2
Kz+oTg2XELTsTrMMkZDcilF+g1mvFBBaUSa5DEMzIrkki7gI85bIj9jtYP2BvWv4
KfqnPMX5rSeBmO52Qy/PtgtllXrYYUEGtK2vxrXsL/gUskBPzcF6JV7ziICxhMIx
8by3MjB1l62C8gS29ZHh9YaGBhB3g7X/BwsiEJz43XdodgrNKLLjSjXr3ccQgAoL
t78tM/cXwwvu2zYphD0bLrv4CMD5ULJVZ8OwbajsolEDfoWflLYtaV7pgyQB3dUt
B6xHX85frEcYEk2Zcu+zRK3wdG3GsqL8rlxFkNFcXKYb3ZsJRnZtfIq6tn3oowVT
ii6oABiTncCdA7VQst3wtw3NAhdvWgo9rL0Rdok+mHweuUFGaPa0TBTtXICv3As7
72cJoBU3y+ZfdB1PFhEXU/1Xh5e/UmAe55XmLID3PblMMoWrjP0swtri5Fu1FQym
xvUDYB8GGtpwW9LPAUeh344cHUoYqB4a7OhfwTw1Rsx7JuHhwA01tLXlio9HbKBD
RjwcmuN2n94OWUK35CO1+EaR2ryfJENmKdkX8rSNuJiBFci9LmR/5KCJa0vCsBnE
gJv4MOLm+x/WNtYJJe5+qtvOReKNawWwfaazkyEruX7WcEqFzoXLdcgDTHLZtAV1
1778ptSdDdtVtusW15S/ZlRA2Ws2ePD2zThTCOsnwAmXKROvU9kQhvVj+F+YlxnQ
Ys7ggkYif4YuYybPr4dY804AwDeYzlT8uN5AqVFfRyWSqxjFrx7DuMqMXVfw4il9
zrG8AHFXfXqoCRtjS5hTgYQpjYZgnfM/LHbCor4i8qDTGxsWApV+aCRb6AuC9CbM
gi/gMsQHc2Ij0JDuIaLIQXq91ArF9PN+HPA+wXTqE5PFDoi/A30/SE5iDjDgvLPW
F3F82zsBa/5GFwgA1CZlLBw66Pmp8tkcjtUpNbz+jVM/5V+uWY8MxPJQ39V1TQbL
4owG9BgGOneA7s4lcAPfnbcGbhUa74HKTW+1I03NvwKIcnUupdIY1cbsPOp8wkyT
FvCa9evEcah7cZwP7ZiC734qvL85niEO+koWhPh6CLLAc4zYl/zxzDytWYI6xhY9
dEXuacEhDnKNKGY1PjS0j2diQIv8xMozn9/7f0duwHXZ0zHkWmgJeNF3+h5Drl6k
oQczVefQd4UAigiZwxe2XVpFzOmoQkteFdNlnTgMANrj/XTMO/9NwODzwwRoJQfq
dzaHYRh2CBtsQTijjUS3m5/6m9sVO7kc721LKY6gUDqSn1OsXaqtNROYw8y3FCct
BHCYcug8Gta928pVP91uadonq4uKzBCh0eedCob3FAIPcvb+ZYk2UcD+9GguyQxX
A34SqG4O4TrI7h5S3LjbHxcG2suvZpm/SZ9zwPMGPJsZZFL2vS98+gzjjUP+H+7i
tupxSDNIHgYfQ+PURMqyttbUMIbRrFwFo6oCEAbPNnCjg3SNjBRaMES5cRJjw5eq
wPO/pEkLJk9d9XLOQk8ZZUu0/5fY7WrpWmvLouW7/PUufYPA5DqZQUOMc63i68wA
7+PaNJmoCEZxpW9kCbL07V7LVAGA1kBVqJnYrmAX6Oi3RozgF2LGsSu1gM0Cuta8
LqzJjTuuqzGaQZBenRPpvMCOsIEtQAgwxMeVjvd+bCFR8TGxMOqSHwm54Q2jMHsR
nwIr10hC2vWRXTf6mCnYSrN5DQo4Gzuj4b1VsispAyk/PF12CGleTFUDmWRwOlxp
TWWO1vWW8fte4oHXIG24+c61lEwO13y+ws9yYkaW/ZlZnY1DlaHjwjyC98rink0n
58TRU8dKjhr6DgDjBHq0nkc6gEclRCcuMyuhLmTNBCFH3jvC2yD9Bi4HBLdcTlRc
EX1xEFZ7XA7dWFHrwsGW5jXJF7HL/6UIhu60ahm4vmyT/zze2bwA6BggRLU1xFJN
d329itJOZncfsW1xXc9QI9X/jNnnxRb+6XSdq55QXM8B9mtmnE8oS08nhR8Qpy59
sE6XEXfhja8UtjnGQ9OcinetYw0qpOIi6S9SP7uK6os8fkFCD8dUq+1+87/KKMQ4
321JTzFl0MDuwvNWVNNPp9s06BIbbYUAtoeTVWPeCrHD8Os0jhXFzfIBFBfTgkzC
+Q2UlIIl6hqWYXZZqG7xh+Q2DIKfMtk3/wzfVGiNb2aF0H0yzvHtxXc37btS4Syx
YWu2Rrd41DzWFWJuymrcluiF8LZfedsnKqw3mJ5rfh41JNENzaigRNRduts6jM1x
r7W8Mys49rZzXXe6K69rC4kR5BiCqtoZDP/RjPu5wdzpjWTzkFNf7/RF+jzPTtLu
Fuvaf/FqInzuCzuG2ookBaO9KnD2pQAJlaPPG1JDYqb3lLZffjMFLBYgQBuWdBdn
NXmHk/q3IWM6dGPaDP3VfTsftNTFjktvoaFNAmSyskbN0PFV64VWp/9v3oKx5etr
FeZ9Phz3Wuz4ZZ/u/y8QKN+l4IccXE7aM9ifRuMJyxCfXKMc6axBnjJ7MaWOl1rz
Xlhdsmt/ATVkDIRbB1837ReSYPhifL38PTCwtrEmb1l2fuQZSb34++SPDU56e9H1
SmPSgIxaIEWrBHQppGcvMDOK9slw82kPMA1ir3CUie2Vc3HNnM7u+vQOXgNo2CTb
VHhml19NqqdTkzEr7/Dd6NTZRnZgm74DOHpocaW/TfXEmurjHAMvuQHQ0ujZp7O8
KCLzLW2/pqgV6nSW0LRf2jPTUoiNtc7vxZKdPNoF4HGYIw9jzR+650nkhbYVUzEx
j7k8v0LTDCAByEkYe7UW4ORt67DdxB1/1vhzUcu50bQ0ZzDe+1C2VX2juNeIeNAd
tiNC/QVmyeKY7u8liFWCqfPV754xA4PXus7W7cnUlv/u+MxaIju7VF0rMaVFi8dO
wXLFyFo++5fgvoSST8zBHTPVtc7Nr9YCqR3vtJV8szB2B2kYqDl5fGrgZ+xknpG8
Iw3HkM7AdwGNNLCdxX5aV5NB4lRWasPPElyVb/zeFKDi+Kp+lEQ6c1KSmVT6TFEf
C0dI9ps8/MUXGTZVRpvk+HF9RBo11aAXXuysJMH5dMr8VW9fRVFqNQR4mtp0fTup
l/XJaQg74geDQZnNSBSfRy6SI2V58EAJ+/IJBEsn9nN05NG8r6K+x+cXLxFMGGLB
dpb+HdgJICeKHOmpZMMl3zeLTiP92RyRvklSHq5CmoJeT10tcJy8CJvMJDb44Xqb
ypMzBHcaFNqbtdszu3hxXNMYDK4koqZ7hdLtfXnXhezoMeo00coU0B30kUokZbId
ajpAm5UgGhencq0bxRljDzDTb6njdtUCl3LwS547VYG9iqSLgn5K26Fr8F4N1/nn
ez+S0YVHRpnGMYE3bXj0e6n/vk9aPQIoNMXy+VNJpz2KxVFBqKRQKvDk8LSOzrZ5
fraQVhmfRnKTsgScF8jxK+HQbX1N/i3jz50Qi4B+HLKgdxzWiKBpgYCYG9uTkOtF
Shz2V3SI55by+fHPl0v5v2vv8cXgIl1TdhS+pHOuFR44A9xRgpqBXnBcfiQnr6v5
8Is51ned44h0OZZ6ZjogF1USOj83qnHM3RpDWfPWAXW1vYD2oiMWkUKVjo1TKtO0
qCat8jSva1+gJFmRVYcskmqLSGYH232rj/Q+ke3P4zhtth3nAW5QvV0w2gtBdQ15
XmslOz3Ar8aOl9x+4QnDDO3hu+ngeNL4FHgYgwwlVbAIFL2PccQsIhle0NmU4ex5
dGTumqpQipX/m8+Og9gqXLSRaws3O85OqPVVlqiGt5E+JYoSPlE0iq3pAPkyWnUv
OVBlUwauWp25O7PmmAzF47W1WoAYCzgX5IAQ2GYUFYxPDW02DRbxxzOqu37z+8JG
9DigbO5OkTUcbhB0bV6r5n2A+WLIMxQaML0KTrkBKA8BtXKkRTyarggnWcOeBY1Q
tGxxDqBbizmWf+l4jIteDyqKhG6/LrgdlMkTXeYW59ISwemI2w2cMSkfwGemXm1u
dmZNtC0LiEvw7ipj7rovQZMxMl+GAtWopVDHvdGmJCA3r2mwoUlK+pH3QvxhVWWK
6qcVHHVzslE4iUrYwTJE8Lg2OGKWdbbDc0gVeRYYXORh26U973Ud+T17AtZ0I0Dy
2bOWt0lKBZQgiv1ouNNffukTmKYeq9HbkBrxUnQRFatXzwdQO2sOOfXQPPeLOQAI
Ogx4vOk60qarxvch72tvOoeM0ROckBDEagSlT4JSBk41oHIe4tBtSh0ogBNG37lI
saQbu1X6BxQTZTLgWB4bMXhWpOn5DFGXTsfGdQFbhbXQBEMA1ct3nKI5Yq19I1e9
3Fat8tlMKvl1aiGZMR2R7+/RZVviGlnbexC5epQ67LxFeOwRefCuYUfJ5kIH92mi
PUeuh1viQDDci2hGlR60+zzvSsZ7PkTYpGddbnFeczkDyfQ1Yw0HFZWUO4u4YrwB
cP12qO4uPX3OW7Y3NoKW+7QNzktTzCHo8bZ5lZrBvyp0ywK09yQJl1I3n9My8S8r
TPuFaMKH2qxCRA82PMzFdmVOOXtY8i6IzBBJmPLndtha05ZhlztPCFU3IoDBEvr8
En4AABf/Jou/4w0ldD93bKbLTdtoWIN/Bq0cQHGeDJFdTHksFcYCs4wk0Su13OCa
gSoYpMgB6PCqYAY4G0OrLhkO5QGWdrSG7OjSBbiBNQmcLOJwrFG2M2i/PWwM5foC
6t2UgBHcP2SUXCfTIB8MS8U6HpO5Mtz4Jc22qtYPYrG/j1+8NDNdPWWQ81o/9tDm
o/egxkuw4Kq5wkjBnwObt3c7G2Kf9Xapnu4XFIevmsAXuguETJkGFErMuw67dSWa
oEd1mAekZ5QyFIgUT127Aj+QqBfqFI3l9u+KPRRiyTnfrWfl61tOzEmpNcjx6Wvp
QAFdR6zWs01VGiFLHj/6oGOfLhb3cPspncfYRQjAe3Gc42MY//S8PFYeRQaE8vjW
O8c16KwMjYx2Poa0OC0S0JYV5SFTtb3GPcJVfe5jKroIb5dgSBQPZGPrj+Z13RwL
YExJ0tqXYzDCZdwPpgCTzJafH6o2e1flQIbFaByyivLGTdjNSvVBOliBn+YVq8wi
KIlnJeGjBZEQNa8bbuMn8ltB4gicY6Cm63ofvGxcPySwwe0pja8Ngqi1JQpVuh6D
xOF78W+rq6yQtJgWhzNq99ZhJrX7SrZjuA4YE6rbBJ2psXUhqVJIedUdzlKHcy9S
bpusVek3ekpm8apJV96xX8XYuUr6QAcsrhT0B1xsCRqQn4r35zy7oqKDXQMFYaah
MQ3Qt9XMWNy/Gvgmw8Ng6JgDD5Nt3u9UvJy2IPHF0AyMbXVIqXk2d4LVO2UNsaOi
dL0g4xM3tjgwtx76P9Huyu0wkuOQ9MCHqHNYRWXOtyfdTIvmqhkCRHh+v9uf9SIV
K1vYlTLq0ra20TKL34Gq0tmdV4VQM4I7oZWaWnfvtgAxqVdWOEUmjH3p0kvXvtaj
C0oMTsDbY7ROMrICED1YFtgRpTiAH3IADspWH2AuDCpv0cwqpp+jxfXKT25edWwm
4seYY8QrluDfIQkVh7r98MUsSV2wlAz5m608/e/tPoMrrCA7QsdUV2w8hPNnXfNW
B7eGpJ8OCuDQbE3bBl6lhtbCxDbAS7p2K0SCORUhkQr//zkgBI5VyJAZp7Ff2NX4
lU6McMfh6BSFpXTz2lYmIYwqShQPRWY6ec8+oEb+MmLJZrDCzP6qxu0lFIS0WQX1
bIVxw8Qe37aRNOXZZHoLW5uJbNslmvHJAVmKQpMhlkQ4ZLNJJpxoXypIN1IodFPd
ucjE9gySr9d8x7TyRiKj2672+lDc+YXvYqroxGcFSkPhYGdyvg+dRLVayLW7ouBM
d+xIQrC2rINjaVOTxfs/ACat24P6gsqlFBxuiNXP6h6ZC9ifxPPXhmSzSWOuHr9I
JgTsMAjKNVqQg3uqhRYNJPSI9bxShJAm5BBEGm9ze/awF7xlbuCs7wjftpfWSyrn
rkLRA0VrsR9amJ/0YjE9wn3AiSqf3+8t+Lhb8Wea51+HVgljRPwvVdcZoH9chVAD
AtJz9FDGhiv/AWPLkKfrLkBBWr2k+/qMUrTiyZyF6T0xeFGHOoZyf9UzoBonurH6
mGi27Q14d+arcToCzVT1B6/I62td+cqbAK9PCLbTnlETlg8lEaMy15xSQHeGXqFc
D26v6258tieSMZAQ4qLtrDiz7bue1h3tV2ufVrc6+roaOSXDCeuZogcHSvJ8SVLO
u+iGaC0XwJOh3xaxuMQXP0Icgd4RelKM2tOy7/D0/GTNuBSPFWM00RP9NZYUZxWn
09SJ4QFG7VnfrkshW5IwgR/SzJHFBswmReD3WF+hm0l6nYiRWN4SunCl0t3IiY9R
3hfhVPwmws5MU8E9G/b4i5WCwH3iJsIT8t2iPXCmrnDDs4R1svc7E7GzokByujoy
iHZ0TwdKRx+l2O66dmNbOALynx/+7RO5L214LqebqDrCZSOIjExxn129gb/mk/o+
x8dzMWY3UFsZJxu31bWMD0I5jvcQy2PKSzoeMl9LhMMCl3LaItsZm7i4cEDZfNcz
CTDw1XECJy/fCpjqvq//eaYTfqGtaIx0SDbScmnf7e98Fx6J1UGES7TIf+oLv8Yc
EdVEwA/oFJqyXxh9/ZRtFICVjBKNLcED60wk/vvbKXOf5KesHSzKyg8y6ykdq1FU
iBtlRFetzdYkFZ37gL8vzGHzle9dRWVu9tETu9vbf9q7FA4V1iknRVikb5wEsvxC
beU8/g76mTsuFBnSn1LXgLB6C19LOJQsq04WnpDFA+VrUlF/RLuXO40U9WbKLu5A
KvhUnDv5N62EAQzQvXFSLEP7Zy2K/8IYhhVikZbHkA+yQ8yUlqS+fmn2kDBDdHdJ
hn7LM2CB3BIMRAgNh0JUZUOLBBpG3fZGvvNCs00MyQsQq4yQuSE8X1YT+Ivp54xj
Nns02fLSnBQJoN+MamZV5xrdVdRrxCp9L/FTDA9EZzEhRGMZ528Juq2xe9sqp/e+
ujfTGhT1Il5tMCBYdENv2Axxt0WjH7jQRh4FBFpPUwB6vWzhdpfUp8E2Cij67vUf
avORtRbN840NxKmRbIcis3baG6GohqruJo5r9uxbEL+MQvFrmToHvIZ/qryl51/o
act62/+D0BsXhO5WIlpYRLZpDqF5PTG4Bg9ZnjXw7UzfH/tXGg/4YdjKO28gXq06
JB1QO4cTdE4En1Uc+sxcG9h2V6rx9Bxc9M0ReiFljwzWnTXrloqd7ZVdRmaNPKS2
gtI+e7z4NBxR81DmzAz/4ZWVIOiIKF6cFASKYA9XBD+XIf//ZiittXP47z5DsbWL
+AlWSzCPlMIu6bQn0ytsf/pplD4YnTWaPPFZ8rxmohiO5P7O1mQ9Srfk6bP1mYVK
BWnuXqB8J3Xbnj1UVCjJkWhYGx0wdykghIvUlCKhPt2bZ98X/Rj+Fojyu5zzQt88
QyycsL5nEda1UZS2f3NmHAQEj26W+5PH1AcR/slO3c9nLVQFTCzKtkFz9Zc5Xgkr
OopFFTaiJ3/QKHygS9EA6C0a6Zr648vul2TrssXsONxox/os9CYvOnKcFZ06UU/o
Hzye6wi3b0vfZwymVkNvGAfOrPQp7T6Nd5NqynGQcUupfvYfSnF/SOG0/7+vaREu
fJnJxDKpEknicV0dhzZ2F0Pcq63e36QVnnLGKacJJIFaoQ5IGhZX/MsF4Fn9n7in
zywtQozKGOpPLq/8HQkmJKiYV8JB0uWuruTBqi10qSOqfPMHax6zX/xYOg5MeVYQ
NXdWcA3qlbmqwOpyv5x2t5vdq4HxgjehJIGsn6t87bNQ9MsHwf9FElc8ZMKHT0eQ
yOtuW8HeZGgFXRmhy3Kazal7RngfVQdC/piUBBtwpJoGX0tyhF7Q39UPySn6KcLy
/Doo1if+RZounjH2nsA9MRF8hz0+HdSAdbMSkxzyzfILyh7E8mQJfymJ9PhLjREB
ROVrEnjxf3+3f5U9afks67XlLpvSbdddg3K6mICUGjxB4ca4+e8UWDVj8GwFLTy0
QnTO5en/o1hjB+asIk+G7TYaXNVf/8hG7JVQAJye4XLLEM9FOSuOUbs4PqP4nK4i
xVJFxvjjdLl9rXu+KGUSM2XBbkmKT9V2uwMhuTr/YicC6K9NQTSDVpxUvL2S3gp7
cNr0uxLjg87e/nA/7EX8t74+sz1jYCNbcp8L50K2wxPfPBaRDTGqMIs0GULXmz6k
jfJDagSx49lmuTKukzkDdx8XqIKjDvze2IHLa3stKGLy0pUfa43D8Onf7id7K4iK
nsPPrUQpgo2ryEziOAhNcpuNdZhmW52Se8nZKZMgayWO/qPwTdqv4mOjU8Oz9rkD
1VV6w79JacubZ7I1AN92hwhGYEpKCNytnBgDvsvvIy79kmkvr9KRqtlBdT0ryzj+
jaCeURVPlc03Lfuqf494pO1YUxYh4w7GT7yZ0wh5VJG8Lirqidw9TReYawDehUN+
RQ9/MXU2AvZDa5Pc+T1gXfI3nvl2EBCnR5XGFyok2uCKS0GMo3rR5Mzz+d36BY4w
Vd0EBc3Odh1p2oxGMoSdZdprmwVTmotfIFQdy8y48zDJMywPKruaPM8UiOYbOdjE
lOJDG3leYaQcbTvu+VnzfcBXyzIP04vzDMJ0ROv5oizjr6cQ9rlYZ/226Dot0hp5
0O5J+a12UshKhsij7gtPSan/BJMthnIUIzKKCCZGaMXOUDRUHCLAw+ym0xwkSpVG
3YBZ6bdiESQNzmNYJJaqEwHFqjl1kjZzVxo7hv9GFLqUqBaTnJ8ALMP+mRf/Qaeb
p+1MGPiKQz/TTGitQpg1SKF2xM2gkGcdhMGiiH0AiVjRm4EGmSmZf/ySRlFVJLoN
/bqhY9ubS0rjA4jXYpp81naJGpQb15ZXX9mlvVHr7Y0hft369KLGeRC+uXFdc+O0
40F+skKw5dUo+GMqGfvyWlYCPzLyZudNmjbqU0EC7yVsQsG7/iQF5GsNiWzsDW2u
zZDY1ITM5YMr6ulb0kzklmn/2jTFQdo36Gc8m0mG9RL8lblEPDAoJrIm7WqzYKsb
jl1r0vvN6sNY3z2GVI75rpaN9qKb6JlJyBF3+w4FuukG0g16a2CuU58dJ3QgYIVe
OkG/HvnOi70MXBbHk8ywBhoAHilEKt+pWWJ+iIMNolqikF2Vl8dIF8y/nwUsRzV1
TfvqdepbXo+lNmUI9RUM/ScJR5DBTucxNqWRxVUfn5i83yReEesKfZHbhICfgX84
K4AGIp1ksajSIkYx8sc/jw+f/6YJUd+s4HMU7R+bfKNbMJfIA20LsFoT30RjTukk
fet0w0saQsVB9XqXNf6aq3COoKzLWm8W8S8gL9GBodvB6hUstHhFuC6suhjwE8/U
9VTxZqZkFYlp14o9OfI+owqJQWBkrv+j8R07r954PDMl96IE7pPH12mRbUhS1FjH
Tx1VUwftdCL2cUkI7dU9rNy84lLkjKvGjeQhJHeGIQ+Lo1/7M4ZrKzaDSx946GPJ
qKSrzD6TdXUceU/+UoE08x0HgPUEU1Q3TIMXp0eqhaWyjdQUwsdD0sT1pQowIuV2
hOW2An35Vo19YRVEn4G/prKNZJ3MK1aBh9l2OG2L5Q+/3DwQ/Qmt3Jbt4dONW7Oi
A8q4AqBOAnFQGp917wnXPrm1dOcZ/zgwxl15+HvXIs9Yz2n2Yho9Xjrz5MZiONtG
ElLM5AU+/28X67xQgcj3GhiGWr1tfuMiBS+G5G75PrVZIUM+Bw2zmbtYlTptyyg8
RHGizzGo9COi6HVQEgWF6cS7sXsZ17vt5A/lrBdZbVnc8WROnOCwmiGdFBQyhqVh
/yOjULc15ghE6efWhrhC85HKYjALV7Lnr8QpcX/dbpPMWwMf37SBCbmltWOpGkuh
7u/pcvLq7aetNh76A39lTYc9xATu/MmfE+d/0+5D3s/3cWhB2V3O7NljLDF2YM3z
Hf/O37drTFJ3lG1MhwCiJSpVhDSeEV+dtOhXP+2j3pT2RIxX7raJnAlitmILW732
2j1N2x3KIklJrSanacA3HTl8zboPOiV8Y6WdaA+ORzcsleVnmjgnailKz6unRbqj
2SHiOW7x4UGXmL4377kDOL1nILyeHU/RCaYVW1P3+S9tnBqLCQr2oE9Yx38yHs/l
J8zwCBzrUp6rrcIyLaUjG9jlkcbuABzT5deVaYuxdgj1P4J0EMyVpBZDZh35x5ZB
QZQP38q7bdcjzdKU+45acGf0G/3k99HOLe052iiQ4V34bII6yD82IkMFA9VManEQ
BgGpLhZn/3s9EE2IaiPrwl/ICk+EXzr1vc3BQkUamkGQBDf2SNKT84xnHzf0JrKG
Q7HhDAL2e53Oavxvi9pKmS5OKudRXXp6IR4cmhQaCLgmBRfrj9JRJgV4bnoLRKtk
1ZX6l7C+/URUkUUMC3VG+3ofcMbp7AyGdRODWgjYuhdm+2XWVdlr+/uBxq/6jO18
KEGK2UIyKhQfnQcDKCatnWMXJz9eqPrhgY9Scyj23DVQenMq7ybooMrzxCYR3XC/
1GbpJjrjkOAwvD8I14ZuyUFGFVTmpQbdCmQ0IT5329hvyKElg+GakRI48D1Anx35
oEGBejPCHekb7hMk81UTvfKbDpmmHRzieKBOT/qFYDFjcT8XLN5zIPMAkkVMXPhk
5rgWZBfsuS2dg36WxhYsKMurgVb/uMRwXHT6EdWMxJIyuKpzoRclgYECr+DpdInf
ODWKXqn/z0Ubzrp3kVA188k8rTGO7DHkaUfFJJBPl3HEuUAeodRg+ej7Xmeq/yeH
kzBC80Nfg5YvZhe2J7cyq+NJI/8rVn4p6ufh9NYKHWkN6mKPLNvFZUyvvANxc136
vi8HC5Rxc9ZWat3ycyonwnvCy/asgKrRVA3f9o0k4VEL/tDwzz8ynEvpCa+ZmIB9
xFLfOKFzkpTriPJQa45PuieKOK7O90LRZF/IFAhyVDBIkojY4KORs68azuT/7gjU
HteUKjdDJe0XOhlhI3Ry5j0oZH+d6l+zJefOnvMZhoN/zyIYNrx+Dc7En+XtObjL
LMJA6nEuwZkWX7ifYAObKkil+t0OctqLxjFIyH/eNM52WrI4y7BCJ+e/B9zwZxes
ketlFMqDz/R1bM0bEPi8bPiw1YiGblfcgmGfHqHt/gvJtxBZ1HpjjHFvfs4ujLQT
Fji3g6HhFgiGPNsIo+KoqquTNWsxYoV9+5DPKWy2MRIER+fCOQ8CEe1B9hnCMsUA
X7Dyz74OkZdozJ/+7Waj5IGgHNrT0s6suySAyeDN9pHAWs+UCYZzj8+qgrkQenHg
+QE7fa1ojb1fNZGNMlP3Il6hF9yTAuMx0f3PSI63ugWWnVZhfIXxGQCy0bwAnCiQ
lspxdqcFtME/zQ/eUNrTRkLx8HsP38bgRPzv2MxuIz4XG8wro+WxkY/Ri6bmcEiI
p2Q/t+wJHJbuGl2ZffQfIwWkniI/NnJvK8iw2VsSAzcAsv9mXxYtcH9JQMoBPE2U
K5LMlniq+8duq+WbCFBC+IP64ewQUKjC6xYdKI+oNZfR9AqtaMNojY6LvlqUpF4v
8gPgHQ8QsDsNpMU4SUYPLQ3g1+KrsC56dPwGfadxVVQaJTbkZixQp0QxBPYhEKYq
TwAujapB2tVyymTAW2xNFTXD6fw8BUyLlXFehbdx4i7UdGSgbHRBIolWSUwuKA6S
ilzzTmknuhgitGAveIVFH8/jffM74Nc18nqYaR7AnU3kvuiVTI5qVRuUDRLU5XJc
W927U2VvfWO2/20lZBhkqnUdS7WdySH0d7V7NrDDpqWT3cO2j5TplnMnkUvR6tJW
O3iSmO62ajYba+r5UtwaK6XTc6a5/9044BjSJVANJJP9ccWPp+S7aAC4UHNg148t
BQyEdT4hcQAYgYEk5Pf17G2BE1QkL+7DNfGwFsXAVb2dsN5Q4TArAVejHgPfUrCY
u+HuVDuUcoZYLHaQt9LJ8UGJ44MsBGUH2TjB3qzoJLe0U+hPj8O394bPVD7hEgnr
/wVr7o/sU5LtqelSWxhVQGLbif4vubERHcVWOoXUBP8/mVvQi2nHfq6PnZvxlPZ9
81nOjaQdBUwn53WbqeUsIciDbpXV5GjC7OFmvwRtoYrNwHu09mGiC+nevcpEN+06
HTn39BcRHrpAXXemgjZus3fMQ1CMXlJrpkb/g2cE6t3Z8RHfztETWeIdB+coK8gZ
pr2WPT8J3U3kpDfN9ECF4Yz1NDkfkOVTj6f2smIa8ft0B0SzKzbXshh1Y8XdtTmb
Bpms9BN6lxOv3gs197zdVyQ/ivjNZkz+JZyIhLHNWwxk5i1wrfdk+rHzAJV7nhk3
LPBIqKi0rDy7UNntyKYR/MRTMi9Vpn1vnon2wS0kHvaHO/DcwDUakjuTHLyqPeq6
pOqij6GYVAk+fjfmYRcVW2C9lgXjWnD8KY5Cr+fRjm1jVtpt8NrBePbxICIkQVu6
Zc66bdO2+/tqtjns+cF4kuRI9Qfz0/uGPNL5mxllaXJOwYZ9jKTh8FXQBpHNWfqX
4c1byRi0pkAOTl5BfPk3Qq9zlzilpJHPbIgQsxQzkAUdzOYtaGz0bqIm2W0UvFEb
fuFKLDyKaFREjyhyTHqYw1NW8e80kKMnqJVYXCOMpnYUM9W+mG35zXr5BEZD/B4v
mLxuTYSLLza1m6Kf/Wof140rFG8Gnp7wqhEnjiIgqEkwVqBhhn1H4gatmpJiwwJO
bg5K7oO+BAv/QLSiBdEFGcOt9HnsqVxpQZyBWUeNrJ6uy5UWVkse996KgNVVF/0P
H2V2b2jkwUKnI0jfGfcHgSt/AaSh8TxjVdYAN82xgsXbbx5F+fCykAKnhOCF+o88
V2Q0Vbj7rmi/n9GSoCl8qsSUuWzKMjDs9JaoFwFWxHKUUVlQ+cQFSDLM3zKkEvcW
oWGDMAax84wbOU1BSdD9NnolJmGN1IEOVatJAi65L7uqTJaYL18+abTIqCo/DcXv
8wDPICO/+3u4sf2qG+flxZpKPPFarPBd/SQ/SGryTgKUKaRDlaXgmUz2ELjaR/Xl
vUB+Qo3hqPsN30xag3tey/g2IGDdO/ZLWFp2E0z+sbFQsT/DtL5oAdOE8rllDn3k
SrJMY1I/CU6RW0Knzy88Xu2Ibly60PDEFFpKDsNd1bwxM3PlghiGgpMd2mBoYZkF
e0q4Una5zAfinyF3FzIzQORABXXXS6p/n6dqhSAbAMgPOWoPs4hNGIeT6yjigTFC
XGuFX3zjYgBg1ZdlFAsRIYPvSZmfD+J70c7yPLWr7Id/vB/6IvW4yzrjsn9mNqQ5
dfsKiebj+LTz6sEXz+Ok0cAc+UvCU35bNjwUnNno/9hv6nsjvchLNg7v+OVnE5AV
NU6Q6sysZkm/nWN8tRfYQH8oWBtUj4w4baJO3j6g91eqqARXz1YKZcbtOW003Rx3
bh9lQZXT96AV5HUui2JdJSjxODiXvsASpMMZevB9Hs4MneSOqOo96WvMOJ4uqvcs
dcd85+EbXdxGpkFo7nW8hycaaZZBnc+gPv6tjaH2lVbno10ciYAdc0sX7dtn5ENh
x0thGErOjoYI0g4NNiE8wFzBhsdg42lN57oQJkZRt7Z63BiNx0DQUbKMndOL4dPC
XKOEoWaDxXol8M0VXQSexfNDC9M/vp9LLt4aKq1EiK9EzR5tJ9Q1CzqgAA8fC+EC
B6GfXutgcqFv/DlwbNBn21PSPpxn+qt+T1L2fcPMGHPuQRwUvbz3bgDLethgfRG4
G56DN7Cogrnki6PIl6QcnqcgvG6tvkfIwz7VIH5qt8MTOfq8YeFzstsxAR1Vp8av
1yjnC0jIAy2IuRgDspdP6u/dhV32FVHfBsL3YgOqQ9idRTZ8GgJjfTTc48nhjt4g
RkA2A99CkMvGRnMolcigaz1E/qc6hvQnk0uLQyBqhVPosfsqxYeD0D+MK1c6FFbX
5SHlnj1/W/EefUk6QkJbZ5tpZp992MjGe7JUwJgYOmjAiJ9CHxgluKUpYlva5axY
lSevENQVlaDDFyWlu8sdhCvtxH4sCywDo2E9fs5f0chAhp1OGOLZkErjX7iEUFRq
UzJLsDV4XN/I0mIa87TLWZ++cvkRGppRfkMqxkcnz/ulqizFz7KNeN0lV08fdOBH
ywapcS0sU17+8lhtKiF01a6ld6nGt9N9RJ/Gmworl/aKhSBUsjTQzuwlK6TiAhln
0q3DUcFxN+mX+2FJPYyyjv6b4hsdmCKDayg07RMC1QeYUJctsKrqW9m+/jpBYPED
dLgyQWJyC08ueIde08LmOUu7kxUKYBknQw9x3CS5r8CQO/w2qv5oO3jjcY1nPA9S
CFnd9SGR2WjhGR+bWUnRtEEop9m98tV1DrevKPhTqp970oV4y6JdKdx/bSHSqREx
fcFo+YytDuCwX2q0+pvQhNBQTpYF4rNcwPuntgpzSqBICaXj2jLS08eZWzxRh2XD
92F/G4h/2WKSE9TfVT+h9cNcyNsFKpDCWdBt5QTzAH9xn5C/B+U1Wqm8//ohXKUF
EXHP6jZv0z3MD3PnplQtpNKn8P9J7RtOFSCx/kdlGPkby2oqH7//QWo1HvMPlQja
A4JcaBrEfQhZ8stqHE4EjSnTWEtqk12cJNp9Luc67sQ9r3uZViEX61AJeUt/5HWJ
m3LNfYy/Klw7oVl6HOgn14bUB1QZno9DMnHTrPn3AgCcODmzIm/2mvttgIDq7Q1C
oVs4vkbZ75TFdE4sbAYEWZwwMsougQP30trwC/U0DdiapHJ5S2TdgDpVo21DJlzK
rMWR6D6D9xDRe1txpSXDhvPHOqmLcqsxEl+XPHsHWQhTWZQM2CHBNpW2VM4eSgxF
H82st9iXDm+iACOTzi6f8rJv35Xu8KwMNOWtHC/zGon50akUprQ9juvRT4tUfZYh
LzZrD6yUuPSJ+/6OkUuXGH8cbUHXBcY1rNauOQtkVmaSEvzJKXueJ6WVPcaOflwf
idMtwtS0cRsc/6eGjT6d0BB3HullKHXHSbErza30KR+ggpTe7t8Wbs05i1HJi2QB
b6rT9LaDgykvhZeR6k7gLEAO/iW4wrj8G9SRDiG1NFsc+gf0TXpyMYqO8ljXTmfc
qrb18Pp552AMZ0sWgIkyj7oBKlN6MjiplE/O1lbJ1T4ec0xrHDl9frVyBfpH6MOK
VQ7nS2s5pSTG9dskVJOGAQqMD9Yqyd8YpiO4WEGlNbicxs5zR+u1cMeCdei6VOvf
4GUjpMpeJ+C/x/bYkxF3YyUTULZy8ils5zRapW6EkKqQrcrazIsPPtD8IFgItca/
MBPfyczdKf3MlSHOE0jzNfSmNL3zZuzItILjpwaKfe9RzGENjk2vzw700Z0jpg6y
BdS5LQqpgsra/0q5tlOtZ8yWufoZ7Z2Bjmp84LSOpUCvhehTAG2ayo7CqXDncv0b
S9mp8vFzuoJ76l1bo8sLa8fue2du9Fu03szR7kk6YyLquF/l/X6sahIa3jktgkaC
AjxcQiyuDEV3fQK8FMWGg0hEsdpZTqgNXRikgxqHjVrTZ1E6r+sACMhVlKZgpYo0
P3EJiU2Ctgt9677wL//J28HB398X5GF/Ymn7TE9LZTQC2mCdDWeQdon910QrYXKR
m61HLlz5rD+xYX5jAb5RYjTMwRWgQnf/0JB/tNWbdEqXUESA1eKsuDMlv2hZX3Pk
gmQBHaVtksIU9i0SSevkBHLFKF7FIOYCK6u78Mql9mfD58ER0wUGrFD2K+3+LVRP
Yq58RPd4G6lYz1iWwDuyU2wXHtLGERRdSK7rFaS/t87gBl/RjsKI7rQcsK/q7CW9
0XwPzg7B5o3+YXEwryn7jWR2SX/Fy0nCZCsoDo1JlwNPYU4zVO5C/DyHFC09qI41
dbqEHLyTp2SxH4yh2IG8503jem/xMPQbF2YSGg1WiaPC0+OtInBnd+TiDDoY18YF
VElj85CM4mFLJsyZD1wsA6ONa4GR6q5xfyigNIvMhBHDgRXUqB2PMe5Gcv3/Clvl
rDL/aBqjj7m4d2zRQnJjmBQMOt3WGdLil6+06dnWDstcqc6gzwCzvYLlI2uMPPmA
ynmgCFT4Y2VDnMovto5LRhAGEjd5h/MesDscr4q540FoOGw8eT5hi3peymDyuSpU
rK4K4j2dDDRR1uhUoujdzo2msolgYwKgy6RFbVg89KJ39aKjQHdLhwYre6Eu3ZMh
8US1+cFSmT93vkKDl/jrBbgKMEskjGrmL2b36qG2+SYatLFd1tI1yufLBXfCG5xX
8kVasI5Rk4QhHGBzN7BcgbXbhM13NzcOVLrindOHC2xqIvI6zXonrTAJj4xiKHgo
X6mOpykiNVTYdCPg0ZP6Ch3PdNKVOQbcBalspNXdWWjtRl+e4aEElfvyp9fiQGr3
PC3EUj8BoDS3mM0so2KxMHNjmVY/3OAZhbkDaoTUd2JUW71MgnHRx+Qnw76fE6rD
C72y4E/DkamHPGF0vl/x30+HIYP7bZVQN9Q8lfHoRfWWzGkT8Qgi438h1aW7TZRc
Vgx354QHa7ZQXAENdZnYSxGAG8igrDBn/c7RmISvfow5tPpQkZgpLOkbDRytT07Y
NCYDUsKvAycAMqEgy3LGioe5Wuq7ebyEtIEFuIKWKB7mv0uNNejfgjgkPjdgySZH
kSHf0AhZ/gX0WMawwNynrNNnN2lwMepJ4576dIsUzSVOd6pourCYmH9hJOQrckXx
s3HGWAu0T5/KygtXXHvX/opbfgXwUe2glg0BxcqIvLLjdJWLm8Sm/25SYAurXFBY
wlEIR0Nd8oztV0SNoLKK0SNFCV0QzxOYibm+k/vVhkSvaTeoEnvJnbrVx03Xa+9T
+He4CNbYjQ+lmoo1hDWq7bMXa4wG7HFNFWkrUh6fc5JOPhxoj3SyleUzDbdzk4qK
MhSPtwfM2NEpfBcyMzqmX2vetzVrxT0RX0QC/9qOEbS9D6CmiweHlCPWFu4VyoZl
Ywp3wMuhyi7foC2ncF5dm1rtJZYjoBIU8VNtIpuXHxc9zr0zWOmxIqiYFTU7GeHf
MQE4k4/u0ct1xDATDgkdub+f/BDKDNV3bIZxf4PnKdx8xr1A1sXdWLKHl1VEdx1i
R2x36Zn9ERJV4UxfxJ9T5CD40cjAoB52EV2kJTC0C9cm0MvyCb78kmg/qCx0PP/+
JdLD/0/R9IL/JVMdxLg9Ul6s+V9ZZXizJHp73ns7mLKRwc2E+rzUY+Iv50wiRJOO
+yR6ihby0CqagKwhezreIHqGnPZq9ZlWHrjxSrvV4ioMzXBzrD7KN12oaOMTLiHg
IEIFVKqeRvktdKHzI852Dt4g3helYqFmx4aXSxYC7ZkfacLWSQOSisOf0wa8ZnB7
ItHsiI6CnB7Mb+rjzi1NDzmxQ/YjidgF7K/JtSJ0swEc0CQAPmPwyiabsJ8SaOgK
kNvO1uTf2FWqR7vp0Vs8C46cbIe4vKg3ndG1EgW26z84WbXcPMn/26+HcqRY/5kp
sL9lgRGI+WDQmSBbf6abXZSYeBaidFAELhHF5DdUpqby0MSCL+iUDjJGkFthhUBf
f6l/W8cgisl0RBNNUW6pkcdDZLivfsj2eJRt7hPur6vR19MMVX9TCdejBapK4fZb
WC870So3Rn/2x3k//KCvvEOTBumztHB7hzzw31QwM919UD4xeFyO8jo7LySihZTQ
ciJLAK1UU7Icl8kSM6o82Hn3ieJHoN7rBoZjzVZo16L7AKkWMmmQFIthf7MVqGm0
RAPtBKUyLNPhon27B3nSna2SknByhA5BU3QZU6Bav6rGJQGUhWP946yaMsJmXArD
ZKQVnDOKZZepu8C4ueeXCk52hQg8/e1U+hDNKEBtrvS3TMa9/ZaqBu5G2UnUS/bd
fbLM1w+aDSwK3CU5xiPquAcLmxqDD1kH81Ylgzqu9e84X6w/iwY6krdaHJK9IV1D
LsVZyq6pCWSMb5g/Gcguc3sygi+Te5+LlhsbDNLsHrA5f+OIBLPYAML6l72oMVPT
GLPmxcjXrSU4ygS5KK4wNHUpAh/HiVVwJOXOFTHjH6UCAdUa7h4hx3Q0xSh/+chE
5wktVV3KjMy+Vfz7Dafy14aAqogbfihGIosMuDofV6VAvT/AmwyPhXEqJJ0EOgpG
ZD2SRFl4VkXmD/4JT+ABNf+fl6rJGc6DmYjK9SoEsb3b8CKEvL8esMb4tqmZnVvU
Igh+OXMysUIv0gmG4FxkqjMvVcreSO0LmMqlVSJDxsC9NiK5DG/mBU8kfeo9CDYN
AcxiB4fhc7eB1M7xvuJncO6q9SK40hkzuLrX13+6DZer5T7uhQe9N8qwr2eUmk/a
muIn1sqUc/GPl9138yLKeLL3nsGvjo7f6u94cXpFzTnGujihTjQ32388ApHaCkwD
qaBbKmRKmyDd7+DvISamxSb+iHjwMKIkxvh9PIhnkkXvI+pDuo0NLDEO4oYA3uUw
c8efsGsFCdKciGmoHkclXqMIMjeTtzjjEjYN4r+yjB7hNyIpb+F2oAlZ9NXX6TWT
xi9k/o+kE2l/iti4uWt/O5MQJTnfSA903xD8rEL8SEvQmyfeL2L198lmqMInxkn1
sqLKQjtW6QC6wZjQ9gM0KBSllk8a5rqFxP/81KuZPGhIx3tEqcytayHrwzmpfOMu
/xonIswpsHtGRARw9we8VVpeDZaF1u6g4le+9UytAnCL6pu5aYq9NmBrTJN21Qn7
tfDVaapdH5dU7yAqP0rTXl9yamZTFWfiWyMK/ZALvxoV/7o9XMAp759lEStSYpqS
E6r4VfaIJNS/63gxppADO8d7l2IZ9DoJE3YOcBq9H7lym4pmk4yY11f6yXr646ZJ
jqj0B2yF0Hp218/6tkJcmltCO7soYqai4spfNeRQkS0ysncQRhOKQodpgq9pCHb0
8eAn6Bhf4qYT3HiEPnWaBUpw0nhmnzqA6+4FxntR6l7gK4hpLgVreg6pB1LNHUQa
/I+RE3hTbc9yg8xfj5q0F7J3BueiIc/6hhKOSDKz2WjbosoH9uYBjYGWDQenRq7U
5Z7sflMKZz1IgDiNwLLT9AxzoaUzZd8I/fVcinYIid0hLpxTPofVXdQ4TBTUkpbn
71o9qHwiThX6rslSxTgPDY72p3tmZqhn+fz1Aw70ujzpP7CGlkVQ77OGWs3PO8CS
CTNy4gBB1VD/h+ckdfpsgtGTkQiPSZQ0qZncz46qknqNjgWdis3z6JpWViL8qd3w
KAMKsvY/pnhTi3ftawwHxLvdYyi8l/MVob+LY1Blki9leMZlFTPTQHUVlarU0YYQ
wf3cQO6HTg6P0r0/fDFkPdZg7JPvh+5MsPL5wIcG5uaBtSAT04AmNjOgRQxrTZLG
BtiiL5kv6UdWTR2WzLPnNc5idpGIDcu/qhJhRuiNsR8mkqAm0MdoVh0HUmMt+2rq
k3E0EPZywU5k69hCPcE4sXfLcT3Detkn9Su8upQ5zBib8QmMPisAcAv2gjVJRMcf
YN8x+XKIpTTxwNM4oSfCH1Glp/2D5z7l9kZ+jsdC6Wj1qWi0AvVtM0oc8yq/eaAQ
cV6n8pqsu8lElFO6HQne9lL5sqkI8Pfxhdf5miXozdJhJE6aJzWHBrt/VU402g0g
AbzjoV4r4DGJZjZs2GiP4p5eCCny3J5M7GcruVHDd06b2MOlf4murTm6sOaeaD+y
ZV7858NCkw5ShJkzfd4l60cLRIxVtZRoRtXvvRx6urfkJ9cL6RvRCo91UY9aLiNg
tirCU1qOLMxDgJcbu2H4zLPpLmS5TgqM1R2661CnIel6IaLIKVIBVBHCmjST1vrn
QUqhE4ohc3LbCav8flI6MKBUOvVu7uae58dY35UZ4Q3sF1hGpp5F9dVZpMKNaIAL
UQLxLGQIR1abehzT7j5RKo7TT4mP6OksDwr23Xov4JM6gN9TNzPfqf6E4GJwTns9
nl0LAol8LDo/D91Gu5fgbDo9MbSUUM2ScKIhJsShKywUXnarv9jEQVJ2wmERkGQS
kYtH1OwZk+QHMAFSFjGSOl1n1T2PvTjxRK2qBr7EKTzu05L7j09Ij4pwnYkG8LZX
QCaXdXOe2cMxWc7z6aBpVyDNqdywuBjwQ06Qk3bKltPBqj5h7XItOPVnw8ysh1Z1
pk5RcYUXEn9n4LXpuqaY3SC8MbKyURQWchYFriRooC5rjtjWwzdCWN6fpshIatdl
8qFX5rlh+ZKQlo9MJLtl/9v5z4mefqbvvWaBoBlGG9Q2b0lLbOjwohg4sy+D4tMC
NhbMvnU/mJGQs4fIjyi4l8X/rtEPX66fgrIA/uU8eOjr7uK5KDzx+iE3s0+1ypSZ
4wn+NwAJQAl6REkMD3nve11EwMcJ5OXCeTYcjH90wNS+MhDQL0nMN+dbpbQ7fCA/
clxk1neDvgDeAOxJiu9t2TC2pYoJd457zboola/gC2XHWYmZqV8nOKt41j8nvpKF
TmljqPn+QGxYy+/ZgQTlyxNov6VqDDIZVNotZg/KRwBMDRcdOXk5Bw3F+SIhuNvN
irci81wCWKt0CNAJV+c0QB5syOzH8wgFAHBt4pXO6W1N3RdeJE1tFHobpW7eeYAp
uD/nPybOBGKOMu+ewUv8uht1YajmsLj3xX20x3EElPmDz3x49AijAUlMJY77pXLE
i8zw90HXkRw237rwRpolhKRRYcun+ZyR74JI6Nt8vY5XvY+yjRWoickqeGiAODoK
dZQo+7FSN+X/21kFfCqzyOWHjLGuHsUEcZoKHFDqFW+4y5Ln4n3CSzj1ZeJO8cTu
weMgWdH83g44EbMwetWe59WQVd9nxbBLry46q+CUZOAiFrkxLRgQw4tzkVOUVrTG
g+MMYWxQhvktS25BEC/9jULfscKfr7uB98Ca92JVdMXCmrGzIntJR89+f+e/Hihb
wdigDg0aAEsPvZZRuV61QHc6EhE3w74LdXIIcA+90Rre6U453hz2YZEYNuLzIG5C
5kor4rJVNeiJliQIkTN7mf90XjTnGCmmR4ogS4LWqf2J2BfRG+nUqoEGULIpNo+Z
T/VzwtL4QzIrep4RcpwJV055zUIGCSApDTKhzw69hANnFBgQPNklg6TJvJVjluWv
JyYZAlq+FLJ24i7SCkAhI+RvIhT2ydFv6Uh7RUFNk2JtW6W5+ceQc0cbJ46SUryT
RXvgdISoTKa/jCh0dlplX29tkOqof5dQU68sdH2+L1OVfg54l5sz+sGAszBrrFaV
TqJHpHsIF0Si4C2be1/fepQqiD6F/Sosuv5vd82z52WdRV5shIG9u2CyDJJYoSCA
YPvJNeQwJ/L42kRUdD7RNlr1q0fNiRKb9daxdZvXKpTfH4pCYSfu/jVk2MJlI5Nt
nbIq5jVJGTPCnYxMnc5DY2wDnvxajfXuKhOIpaTpsH2gwCg/W5tGP+pPQyw68Dos
y7iygWcOfBmELClzlpn0NiKOLJ3jSY8oXEupEbRQeARh2S2DwUTW/ED/M6u4rHl3
80xylfLIbzwVxDiMIXXCcb4xcPQwrAk5j1Z1SVRD+fxsoe04NxR8uGqWy1GnwoEB
BX1n7KG/6FRb2wTNBFdDVWTTuAwp7aFaWehYw22gBFLRRp8+Ak7OvcrrAmWuZT5q
KrvDjEgQ9NDgpZiscIcYDH7Dy4JDjRrK0v6o6LqZgwsTXDgUdPvmbYaIUKE1BLVu
yx/6eU0foIwfBQQEhoDyo8V6epNkDDHBdKAZ69WeDre5jrAJXaJYOS4iMF1U/1Ar
Ewx1hlfDCMG5UCrzl/1RZaxDMI3Ix8FVArlUA2DWe99n1vkfDQh5ulz91xuPd3dv
lfvVVdYXaT9fX9vQnljElSJPj+B1dY+5zgIdnJQrGqojEwp19i9/+miN89wbIHr6
cl7WuE2I5XsrE2vEydJIBUWgLfnqheWGuyjUVsI0Cjbf1R5t1nPyD/VKAXN9AobY
RCdbepEZddA1EoHKD09ftlQ0/vQbzHQVEJQgYooy/C27G6aRZ4CY8A+aoxdkTvuw
XvB264OAywscF8bak2HFYj6b0ODh5/QbpHyworMHFiGtexMeKa9V3LFTrH6dyfQD
5/jOOGgQspP376Bws7OyU8t4Xg8sTcuBL1rXHhe5/pqfqNnLtWXBOnxYNmEpLCNI
Kdd+iLYaEuZ6fmqgUkG84KrHwy7jNyUBlGl66MIwv8oMbAMrE6hcTfjI5FlC57z8
Lpu2mzpAJlQ51IGORN0SR98KjgIVS6uMqfs1KfY32vcQxcJaKOzkELYq10gl7udj
0bY4YaKPPgbbfQO9Igw7o8eRo0WHMuh9JgQ2rKaHI30l84H3QlVF5b+StGP6Oy0W
QyehSjLO8vMqqTT/F25qbh6LNp5Y4KivW3oyaEuIfLUkqJjQvRUBuKNRAWl9pdIa
CCCW2j5I6neOBaSIFlbjxRxFd3yxDvrtux0uW+lTxFYF7NDnt7P1V11W7JK2E5c7
S4OBesO3to4r7ZxyS8XDkA50ckaYeP5m5P+fG979s5Ol+78hb/suIqbKAeX6liZo
nnLD+r2auhU2lWRZP/HO2HMeCD5a6ve2G9gEm72IxNyrydQxITDdp1rityO3BWIy
e7UE5ccdyJQ34SdCnwJe9ZLaUtdJTCdVvtZqJH68tfkEoaoG8Dtr+0N0diNHOnXF
axslSr9qdIpka4+A0tl64oXCIAF7rfIqhB7kUXzdrUOl5UbH58FpLIVNv1uPC9B9
TzEuCmz1E3HerGkE0kgdCywuG4nGJIsYSLZNIDfSWvUFagffFPPrMNtlL0l8Ok+q
bY496UZ7REzcTBOIL2d4cowT/9vpeIrk3ISSmmwi11c4mMhUMd7zuYuRoMIaeu2i
vHHHOYXJ6DFbEYgTKSSVjM9wtCVWVfnzNImA7GO0X6SAwBrO6a84ODi/+y5Jd0qC
9Q8enZcUMQLYb02d6GzmYzedwlDZ5LeDoMnDPmqa6zh0D6l7WGJVrrMte1qWLDrl
915Ocbl+2qsLgLpESq69RU1E5IaWkOM5OS4vTtyBrEV4jnr94N7o6rL2d4WiunSS
TtM5R3MBsp2XaairWNs4da5mL8OwqoAPxIzuR/+LHSSom9CdoS6Aikl+gzlWToHz
X1egPLT4IsRIUVixSHPTywoGFbRnM7xLNalBIXtFGDcARi6fMIsUIbPCrye2x72X
lv3kyEx69cfgHKaPkECqEZUVl+vF638A5U+d7ktIhETSjpcZwtKd7yzKGeGaj/AV
YZe0i+u9AlNeYLkfCl8sWU+05YzysFA7SdplOHwrKINhr/zFlummmBw2H2OXViZ3
XBkp6RaicFfplaqVhCRenRiqXPoinoZBWhG1daIJEuuUeCGHlj91RNfhKP9JISZ+
20IT0KfYdjSecYJOuh+P7Ds6JpkIqhZiFOJ7lRkYdwGka6yR6AS7gkZRvHCmLvj0
CZDj5OrsXkBEiqpimNFn+CLDy2KKeJr3RjNfFRUUaB78P2bznvTgAHuw5kTdLZFB
vjY6i8uBZVlEof4lVbucd89fbJwKU+AIOp0cnf4Td9JaF8MpaYOrEwmZnl6FtaLK
rHpBrw76lYaOeJtZ4c6xjh169/9d1Rt7Yy7LYW5adCVv6KrMYRXHS+WN+avWLN9+
MH6obxBTcRwkl+ZtEEiPLr1DdHisFcdh0+BaB578NSJNdXwN+GM7mxtIfccD/7+n
PEP8n1QtQqZf9fUgxIR862AH+BkSAGa+hsdfiJaL4Ju5yeUxaGZj5R31zsQRZQIK
KyDjBF9hrM3YIITgr3XRsQCLi/m879h37BOoALns4kCfSrcw2pbYqEPMF/7fw9rN
D8cEx0qAO0PvyGOksRflH0z0jw//+IJN6TJu3S7XxjR5xWz6mwtWCC7gsc2BCNmB
7swJVvfmerzJla3Q8Ot9rjMmpdjeta7F8stlsj8iZHR+SmfPIIUUh9tRb2eqpBWw
9ntxEtNcINuse3KuquEgTtI+3BEl5NBBTi+Uq7me5GWPgj/b7x05H5qCO4v1WS/4
Epg2CKWxUIGNzzVgHLa45g9keWPi750NjdjFBxEEjJa7NDFw1TWtb0laWfXKFW3t
yZMyvlUPajvnJzL8z3BZFCep214+ZG4S3lMYORVShYH24mfZpk+CTL5Jp+J4uiJU
43KCqTonQSL7I8sCUASIx1KyMoyxxBEiS5Ykkg8RYh6tQ6UGywtRWrqRZZwzMAlj
4gf8B8ftwQzidYMmbPOUQnlEoh9PYjkwwV5AeH3f1Uz3V7ppqxN22/jS41GjAX7+
UYtTAsnk3kfNUDzWvWHKtJ7ctWgHTED8vi+dVIk4tIovY5EObN5UcYunyKe4N7vE
f4GF7FsC6mdQQ5D4/tveczE1pT0oK4kUTMGu4LtD2uiF4LDzAv5w/tL3J6yofd9e
u42Kyw+Lt/XUXpO9vSd6dXwg6zvyk04PRy/8fwoERkfDrD3TiyaL0R4Xovxp0NFd
00QXHhdvGZ5FHA0fdpc8Tu9BD96jaGXqhhV5R5/TrNVT/9N0188iuKHlW4cqNC6K
ta5zkcbNX5o+A+eB30sr46tvSAmSsnmkkrZeB6b5poW8y0ycLkU0NgbbVW+lvH5T
+ed2qsoYe0YFIyLwT+ESF8Jfwz/mLOCqev7Bf6FJxBFeFwVSKMP7vYC4oGSWlRo5
4+nIJyFjAO2Hiuc1I/WXrVFsHy2ROGK8N24sBJ9OTodCwTWuSvBXL/ZlEq+35uTv
aE4S0nBbOC3wS/9IZnMMkLcQFY1+GisSGawJwFlCrHhaSD4tmocl20RgvOMiPtv0
rCSkI09UUYdpHHcWEKJQgsaG/hElQD6kH4GMN17u8DEo4Or0+4usKB7HkTRi2CRm
6RqpsKDhZr6LVYO1K2iUA8iUJJuott19ZHEFbWb2/3tU+mQt5dWqIBZwYBmzAPb0
dVYkDPO8Dw/CcHHZomZC5VCMA5Vptp9moHgg1CkR5v1OxlxgqTEvQwmnowhHPWB4
YWDK75GlWNcLML1HY1TdCKS99C3vF34BUmZyLXdHm2uJ0c0qeFi8HHWkXB5wHiBb
s0Get86fsSWWM/YTrfaOvuBmfPLhD5QPaNMq3OZx/7DHcCa8qZIxtsOvwT/yCA++
r7PhNq85AWlod7beGWQpZJopCK1aWeXLtEqK1MUePDLd526daseonRJvfiZ8uJnh
IsTipbBa2W5ouPklebBsHlKRNKqDOlPYwPbpxNXPeqtaZ08+WmegyFja2J473b5e
7YVZvxZnNGIbr0Ew6xQyY1M3Q1vj1xC5VD8alN8Hmzf1WQWqKbRHVZIBQPWH14Gp
NfKSE7z++tfnwmy+DeJn55qQQmxUU43Y0ncaKM0PM97VdYZ+gnQv4VqdEFcsh6D4
/fPKrmY2jGxH6U9PKF1+jg+zQpSrmh9NwO+ch8tuOgKT5hPiwqiS7XeQV7nJe2Jn
GngqwxWcHd1HpMkYlkjUXb+15g9UfCpeqA1Xjf6GPlVSx+ZRIsUBwb9eeHpq1dIx
dHhkefthhA8QXPmFRjS2MYtyebJjUv1zLFc9up/i6cWFUKMKHbE3gAbs/2DqVH5p
8XbZ6rzpjfRK3D2wKgao7MkvaJnFeXjp8/mB4lJ9oUqs/ymDBtpo1Os3qDvzSl2i
UGmaoC2578kD+TDQpRVxqoNHgz7TJf5ppZdoxVX82dQ6TtDvytrzGq8+U0wFlKZ3
FioF+5en27JskwqM4aJR/O98b5BgtapE4RpoyXD0AjxksPyvtDXGr4hgZwST2bQo
BbsU6j6HKsWMXdCwTxB5q06rIKaed5Ekm/0TE7AFeUyZmwOW6D/KN7nnRlwFOOUb
b6GCC03GXwVUr9f3OZ90+K4rYlMtPYqyLcubOvQwPTbXX2sOgHJAYB2m3LaBq9nN
STr86LBHDeOiCxpC8rw7VAREMeUXPPJSVzWasxCej8/3CExUci8wzeePYiHG7rzJ
JOIWN6Xnd5SrOAuaC8JQ/dVzhh8ince3RQ5Tlwd9Sl40q/GTPLP012PC2WlXUSJA
aBsa5FYKAWE4Nou4m+ohCRxf/hYq05FXnkyEdE2AxsEWN5ZeopGhfbDIfTuqefKY
piLMCVnf10iMTxz1qJCU/LwpBWPyAoGD24YeDjGyu6geePTt2s7KitD5FBC25NOd
5I5vnHHfcysjuvOSkWQYHOLfzuFoJTXDMKicwhZg03iUhMg7jpfXqGnitfU5ymlo
e15AF6lXrunMbzkCCtTsxLgQCEwdG5r1qYr1R0LR1FQ9nGq4adv603OUMyRsghdh
y+BBawoJc058U/PnVAyJDnuqpISYGQHTYqDqDKBlxleufWTB60Zu5den/40jzv77
kukcH0dWvysEaRmaRylLkKGSuq5KjMqsSWelHEKqX/fX6e4W7o2Cdjm1HAMBCUs2
wyYL32TZ1Avp9W34NtO27MBrZFARH1kwz4kxrmmWoklneT9HKXHffR/REvwXzrTu
fGiqoBelDXyLLavjI2WyKil6rS1L5HgnnEU2yMRJYI7sSg16b5Bc8BNOBIP9ckKi
kliQjGaS8Dv5GV9s8YQzUl65n/4JCAbxfWpbqzWtTqDPFRznzjipvPYlojg950CH
bojDl2VWlFGAJ+Z9lcmuYN8o4sn4T0VobZRDTWuCq5xBziBeKx41mITq5nFIqZqz
NO3shI+mWNrPYuLammYOUF3QIMGweazPQymuFzRYJWvUG6qJCbsXd+PIVNQYRm3M
t28PfuwlC4Rv65UwAw6xufhziurPgWghu/4XdtZaF2E4A3AEOZiiRO9NOUtVY+WT
v4a4wFiCiFRxFexlD8Fpnk0DGJRHJTd7x77mZA/RaaeTQmQYbSIB224+ZOtW7HXv
V+8d9RYtbo8DQDNWb/HAcUZXZZkpo88vlRQuY6YvvylnOG+YBYyZKRmmixAbSAzh
IlVwMe4BCLSMiQ09H2sI4RuWksZqRIqHln0mz6uBUll2xVKU7+7Z4Ro0zJJrBeGn
2mGxl5gn82Z5HnMol9BVujakEttw0xAMfuAq96wrMQykun26gXbFaTi3WwezBQv4
nsiUqnPTbXpt/hRmmWxeGGTtylMK8WkEcpn8NSwKH45izcg9iu7qHcqUM5qJ8htt
yVpIlWnS+/MCIv1MAS8vxt/Q8QpodhyPAuHS+fR1JxnLTwPyUcPmTBBoy+IpHnDt
p3t4zCMqO7GqEcCTBjhFj4WzlpXYp4mCcoAGajfZY2U0swQsG4rAifT4LJnFi1Gw
2u2Y84lzzGDuLeitiFFC3nNSRJm4B6a5XmgvN7B3mJ0yjWNqhSXXRR5g6fPzn8Pp
+Mvicyd4iY7fRc0C3ipbE6ZSImyUiX45wvn49ZpLadfcDH6wY086woD53duvjRIo
ggXyzPwEIrK0IDRY3ElGUGQwyqwQCBsllVY+Ljd7zfvuV8YJdLPUVFbi1EE5BAuH
9hQqa0+rC03RJPR+ebARoTS9IbyxfJlL2ISndhl3brY0D9/5GhEk1d/8itwJOOru
l7FtkAgy+qOU3d9EJGXdpr220ldKjqG97OvUEgzuODwa/MCpzy7TzAbKojPmltpT
V+CBBYz7Fba2plP2S+4vDLJlFmoLA0WIiBWWYUw7x4yBIOS5uIJJXxXKyIi9TPKb
oMvzJc+zSN36D2FRF01+mnCoR96zvGhUwelbLoCJbVYV5De3/X5s12lyHQWLndx4
U8Mwv7jmTrdM9PewlXHKCrJoezrL4f0MDgKoXxmXQte6zfv0vkCMqqUIEvdKdRyj
WnnfgvW71yI0xhDyZlcvUvJMwU7i0Dx/4XhcHzzq/qfTyt/V3kqQScWnnmf2zIRW
7BKLB3YoEd1YNJeQxwUvk957QGSjZPeSifYjWN38X9esr5jK9ur0L6U3raSVyFgH
ZzxcElfzgdBGO0IAqBtWjBAqx4vbhhLy19rmPhd13fLup0LUsmtMoij6MDrHi0Ot
nhSTXaxeq+zfIbfqxeM39k1J1cHfePBY2I0SNZZ4clf4/dykLCGTVrKn2/yU1lD2
4SjWiO0RpvIMCevLix0cPPTGf0QtmYy7YCdccR05/gLmyyp/r5z5WADJQzK8qyCU
GI8KmBc/wC+CIG5MioVYTX6Tew3tHVsk2XnOTWiuIIp0kGnv9arVg+MdLIi4eLB4
UEIEGfEb90gn5zdq1+HaHATk1rEjngQF19QUjsctaF6h3r7yYAk1AQLLl4QAwnxD
BmcnAiXUKFLr1lGEEjPmaJqEYpUYbbsNdoH7suRxAXr/7XEnpWEjhnsmv/WH88dT
bYIizUzRQ2E+tXmTXMJ71P3UDAk+JgxFYBwBdoXSwibilWf4qLGZMNWE5Ps0f5+q
13R4238f0BFfdCPeDssxDZnsstTGObV+ugopwo0CU5zIilODBvFBDKKNgZEo7l9s
qZ39Sfwf/vSxkzzyT08esWV2zGQkJPSh1QYTfjA3xKauEZhcGXQY9fjzMlzITl++
fw8T+8dxAQav3dVbivOlxnfWreHueLPZscjvNFJTSV9h2nALWUed0xnXoTMqWGkU
Er7uZl7294kmFegUY2wdapC5VtszT5AyaArXVOQH61fv7yPvJvn0itLoSS40e8LH
tkMB+UK0ttWnD5wYQVCR9faumD9fMHdV2GMmnN8JjE9LQUO+ey0pK/WaCAah5RUL
9wTiY25X/y0Uu8++08AsiyOfXHvF405tESyQW1XFzW7VNOdRCJffftQIleH4bVc2
UQsRbaA3Mqktao3FJM2r2VCJhjlfeIsPIvU3lNhvK5NyPHa1NS6q8rJWjB263D+w
SAbc1WqckUUUHsYGvjWm7cdB1SpVHzLxlUT47R279szK6VCuZh5uabpzsXt3ENNh
bECYy7y7TUFt6Zr1annShTIK0iNE2ws1nuW3yY8RrDMC1KEaCxI1PkpNg9v2vT2O
o92RTu2qdAjhL7O5e/yD6EPR1fV0MKyf2IOXEm3mYuugALNcU0zNAxac6hJ0FXAF
gkZWSAJN/OlYV4EFCHYsGqnq9estTtvTyHKbnGXh2RAiOxXO9TcetrPX2mQ0OA7b
rffBUf2jO6Aps/4ZjNZfYOe/I/c0rw8R2btY0cEyeL8oFsGzj26rTB/LM6M12EFX
YSjTvKjFx3uvaB+26+K0owxKlTkiJc92dYLL1SlTtomwyKaFwQABMjJimNynQ9dE
gtCMFBSlXdvFGPVFK6YmWbwxN+5yveSiejEvfzNDgpJGv4vGcy5KvhYBLKteokm4
cTsas4VyD3rPnIJdKlHO1xtJw3DFgWhVTSHZaKsAjZkbLmvAFGwddsnmlNC1+P3H
M+dLpH6Z8ZTIYE1TsVrfUEl5Tb8+C7ztGfB4CcS4pTDzhgDm+B9dKMKiS7NeJWe5
psSZQnLmJbzMtTXubUgzN2SiV2TU/pXP2j6skfhgNCL2FY5NaubsVMCtyARhinFp
k4BxIVghuyTth2oW4TOkGtR3QyLVrvazBL+gXnLH800B9+6QEuRxkiBwrIpBa/uk
b926zVFA0+R1Hf8hkcrRMgcZxv+GN32k20jzBiw30A4TvweDIkYYrIC4yUIioRWv
cFKCE0Af8t1W1Dbgwlaccx8wRPEyifVdnBZaGLCpULvEK0LvMrVZaPfWRmjw8BW5
Na2WlRflEBG+OZy3ycjYr+U2Mv65LqC3gOyhNoCFO6hy7/U1sOK+wKJmAQ8dMdcE
57MTvC/Q+4Si9B+NpfMlyyRZmC7LEZVbqdTWVJDemE2Pw3s9ZtvbD2VWa4jhcX7o
lZKPHOXIFru/Y+MKB76ueWe7/DidGetBknh+pkqevFb7htu7tIlsJlUgUN5337c2
5w9HXEU02SloXyIX2KYnoD9Lh4fimxYXKp/ZkD1muNfiMCm28VEdvjp1a+Uewudz
a+UkoFf40KUHIScboBKXYhRxUslmifNmrdtfAFDb+zMFzXBXHQhdnH/dCxgaXirL
005lKFq6MPIRkerS67xGbXCfDdtHGc+zo6Q+3glxM1L0VOOEUEi2bOlMmCWyv3T9
j4O3B45Ysk6MSiP01XKJAI9tK0D2cz7CE8hKvs4Y6dGOvIYzFyvkaG3XPNK3aad3
MthZ/HsqCfL70ZcclLJlG62Bei8CrRbocH2XqgvpRZuBAOMAyYeiiADC/FSrgOJZ
DXRV4dFv9x+kBj7OamfL1I5fvMvs9UGOYBq3EZIaVRC5diuqVW9ucfsy8gNGU0BX
2UzenSb47oLtzJdbI+dEnPQC3K9An3zutB/URxqggb+0dqpKmYXmasA4P1Ra0zga
En9yMBZHQ8WyvDCWL3sBn3ZK3DMpubVf3+7VoDvTItk9vRJVgM1OK+uz6UpWxkRL
6CZf4COEWd8GRVyuJMrWcyEHYgwGr7k8nih26nbii2q+SaOzGkmhoeKmlcMvyA9/
wVjPJHBdjrIBj6zCGWTAOwDgCTUSnFvqm7R8EsLEqz9tSX/CR8F6tNxOBZxDSjUn
jDLdPr5VEZgy1Yahr808GBuBO0fDYscrF0N95CtEvz4Tz1S5CTt6x8wrxXrBm8+e
CsFT67vFjr3g9P2s0GJ/fdBhhrHt5NEk06WAHPYxrxN08cm4BcoKlEC8+7P7fNHB
JVEuL0/7YKvrF2vcnK1YUAflJoBoAYBkKDUTtvV8lS4f+WKNYBJ2NO0zUwacOd5c
1M22jjFhZrpfSVMxzIvKRE/EKOdM2ty9F9xs0DirOQhl1E4Fne2swKwI07QsbzVv
6FSYxIxq3xmQSe9a0NYDqU63rgXN95szggYhb9lVRktljFnIijD7XWnV1FyunQz0
HyahShwU38Mk4biol1hR0JUpk/7jTZDpJfAVd1YROzNcIFTab+Ao8+U3ygEhMg6F
fU+7hI9/01g8uVBhJqhYkWaB3uWskEW6KThctpTpjqO5KpTjsFveeGULdlImKkLv
cHbWjDeMcy8owql4Fwv8XX7oVShMsVwydB7XaVMPVXCyicYLeDRo92IFMIEmRhtG
GN/0HEQrZou3cOBOynkCk5FekyCuGKMi6xTU5VmIt9bV3kZ9YkO2YdlzMBXlZKp/
SmGGSaCks5bDsx+SiKamHZo/p1T83fwlRD52RTKj7YNb++VoZDpjrdCht1KOjl2w
2fiSzW+SA0cGMRLFWAJauahu7rXxk10owq0vFUj6ECStl/s2WYuLW2mZePMv0Oxa
C/ZuNxrQ4vDIPkbNQl9YfCDFLfFz9O47mFTQgjW8MOSZtPztqZhl+iWMzg7/4THe
iNvSfBse5IeCVG5sCK9u6nQ7D1wjnz4Yrvq0NmV68XFjZlVeDKRBYpcOO5Stzm22
NiH8z+1aKyt6kegLxImT4VIheOMGLjsnIzGE4odmWEYdlO4OVl7bMy56TF5VNVL0
dqBWylesoQNg6OlXO9zPV4zyJuDj5N5xsE11g7Jm2wZqtuwz5jvfuK/EIlHZSzFn
9i/CouR7dLvMBXdk1G1/3WOgjpx9q19Zy2Sp3W6hYTTBSoIMpNKtElfwnW5ouO5w
vM3NABcH6axbqxbpD7fDymAgLCewzPgCMMYNCgFN3oA6U9tRhdxbAQvq7olEPOKd
Ds5HgqmhBjvWAtMxZZjWDf6R68HNO9aPXqwJK9NaQfD1bszTwznBXj88mYJC6YZ4
1gsadqy/OvLxrTI5R83Em7boVo1xFazw4LAEhzKZLx360PLKKYu5HM8+Fjm0FsGz
2eu/mbIbYsuvfMj4FcgnE8PZEtDf2UHn/itaZ/0LfagAgH+bqCQeBErbPglbz4oF
YQYZC+53eRhUpPVPJPna6WJjsnElVDm9wtIS6uOQSuPj/chpk9PiQUSadbx3nJ2M
CwrY4nf22luRVHiGB+MT2p4iC0DIji0df7ZJU85iagtb0WileBvdcBkM62c4dk4l
wxg2fZB1Ao/tnTcEl9TieG/awxXob8pgiOAlhzDK/1/Pfz+a4B/Ow0BA9NZyNBho
WASQR+ZL/ROAjdqn63mSEJ7hIdi7IV0q7JeDK+ZwybVYeaPEnW4wHAt7x26Zbh7E
fOJTigskW0at/OddPY2AMxCd3609FP7XQlyM+o4BHqm3k4VcX6hXCyz/cxmLGeyA
ANu5fYbyuxLmPy+srLtQeAbqglBGa3bh/sIEa4/m+7JUzMo05Uo6EwRFG+1oFEvH
9h1QX5QHGlk+jm/bcSwGaYMkT4pXb23KyIeoGhwKyQ3LSZ+Cxp3W23fF883ZoxG+
2HUxSZqETpFZrxQqHeY6kiJbo2/h4mtHRtwdDbKlkSOKlI1tIhE1Eme7mUfmEuBH
DQ165q+cYFzIx+mLBXG8R0jGoXachNi5UvLhaHCO8/Hu+JI1ZIsm32ySiqIyKKcS
TgsYkGp9UeFJO5oKcrZyhoXoBTQIGc1pPU7/msR29GsUs3drb4Ac7Dbs5SMrPbk0
eesU0fCcZlBY2Cb0czZVNPCd8PD2lIzbF/Eetpqg3vm7/beZtDltMCLvGUSg0PSf
BsEo0QpPhVGU8BQhduIATbwLF/ocVYKe8SlSLllBv83OJCAH+Fsc7Vd/7alHaoYU
9xXLlzqgYgKPuSj6ZjJFy30sgl4pi0tDn8koTO2GJ5m1yYZ1LdSS5EYOMLlh1wXI
hgC3K+Dv07Tx/dSGfg8YKqgXr77gkiE3VjMCBkTMdK57yYweiIjFtpy/CAnTqiuK
qUfQdRes0RVQ5DcoAczsD+KlKKqAXDMisHsu+iDJ+HtSuo9UVke7y/IulksxSeMw
OJsJGKDWgqRSqP/ElKWYGIm9X4lIoVu6ZHNHgaiT5CiWBwdOCr2gBNVlXQRodso9
9FwkqWRdqP2AvNFPGlT+0ebfxDfuOonU98bS/558lvyqwwxRU9elQsogeenc0UaI
fChr0c6/FDkrTTKXS3pSxSX062Cnl8OnapyjyUFWYna81opvy+W/zo7ZkSJhR/3a
JY3OPQcdpKvvpB8H1DqPnZ+xLU8CARkO4kJ1AOjln+NeqtkvFOSUbnazLHnwtVZJ
UhjXTe/xTxEKzf0yvO0K7g7A/53AzUUhjonBZaFy+daDAtv5W4TS60UQNwSw9hXt
EMYzrqeFAaG66S+Mrm6vz/+xSMQ+FfdM4reE2UPCThlD3RSAOO6yHu+SDTiCmKW5
yEAJAOKM5GzAIdb/x0ybKW4WOR9kq1uHjKhkyl/fetuXLOpjXwm6TM1+qmvNILyt
pHHz3g+tIQH62cYYZxUpQUARz6eC9/0BP0U42F3LBDcYk7jLcjUeAvh91xnr3Kj3
K5fySmIMgBz5flU72vr4VYuBVE6vYNG0RfOeFlo5mEp5En+AmqWRLlv65WHNWZXG
OnOf//AHIfPflL4zzYMmvb6FKN+vwrlgm+0h9cLO0sPHSVADpXba6AKCspKrUbYX
Tq4WRqH+U1xeRoMLGykLJOvhdCJQBvam14vF2PGOgnuVKVWxxJ/drF+biONQ063U
7Mv1+R26J0ir5F6+LLyJXHLMW4kVSrLFdhmhkCv2No1kKjI766WcOIVPoBiJk/lU
y/TgU00AZ8NmAAchb58br3pc+f7s7EzE/qe/FTBHWRYpW+rG0UZa9S42DSFg50DT
G8byKmoBZiYrAurH8b8GJamE2UrQzAXr+XgkANLxP4e2Gl+/YUcfppIqfCNaGudt
SAUyBfD+4jOI5mA58KPkzRYxAGj9dJF65eKmOxw1JZjADyfNQfw+XNM6LpmQEDIh
dl4WDLGOtwsqSOOn3Z1NTWOfbM6x54cneko10zpHxedJZEIROp3G6GfwtXQ3nGbV
9acC9fKFEpuP/pDl1fFh+8oEbP55Wp88Vv7HrnYN62dpzBbemHtRX1tblwNg80SH
CAb2KpnX6uW+giZwiXeCKYZgNk9PpBpIOFgqS4vzl9oAlFId5JKp6QhDtj6gBKDj
SSxJnUJu0u+NMl9bi9d8W/GNopIZXtsNHJibo+mL+tH8z8qnjjUWW5kdgszCxNeE
YCwasYZVNIj68pfV25Cz5qSg1T63+ZbFQN3zUU52Y01apJI6ykS2txWA3u5W7Tfy
hjV2FPBatUqi/iFeg7uKfGcRx9jsHHvRRDRqMIIJ/tFisQW4b6x/nBWuGcATXiFf
WS26c8/jVwj/P4lHlBxBHV38KVb8n85tABnFg2q3Wplr9V5otu6TmrlPhrVvYRjf
PiSnThtI/ntN96qe5N8qqqmiFkoAWyiUKdqLNpjNatNt1xwOvSnVYiyWy8ImPYes
6t5KcolJAmzOGt/DzCncCIBZKVM4gYXWkYPlHjIcy8x9HeyEabRbL66gsA/1tugk
C3N3M9OOkK6kQGjJYLiyjyleNjdZo6yEIF3zukW7QAA5M18EKowImMHQO3xjikwm
/i3WWurtRS3DepTKy+82Oj0MGlcufagi4h9mD3PEX48jP+o1uMvcsmQq6sMR1zBF
VF4QvRBg+6ZsVYD9UP+7oWsJweTFXBE38HbNbaZy2uKvEXJ2HicnAS07Yl/zwPRC
51RoSrVFhLs2+klSX5DoS6SjYskbGObRX9qoiboglM9Y7NxC4tE91XgBrJ23/PDs
TSb6ykMyVRE2HtWGzeNcX802+L3FUlbZq1cBF/ruPexZD1iVdS0sc74VMm60534T
fVB+gUdWcim2LLBPlMfwp+6LHanBjSWRVTqKKOsswcfFS7U3j3HyF9tdszAvprFQ
9QxWyVIYrhzyzSpBFyiutr8b/2vT48dDNb7sUA9onaUly6zoqKjTWCKy6RujAGI0
SXBUZ7TI22pGMxg7ryC9T0arIHfe8zpafI+kQN7p3irXHRkwvgWZ+z4uTzUB18zp
k99fYTZ10icEte2bmYi3pGVXp4p64GzibhSpO4t+RNZjd5IN1TuT/UWEgz0ueF7m
a4eGmwx3cu/WAsIJf4XTnYLc6cF4LD5Drbh4lEnBcuXuLPsvO2S1lXlgtK3n1d9s
6XMJCUTxYOK6OYPt5H/rHRf7Aoivl8S7AnadNT9ZyDyuNzkl5aGRD38W72pZFLHP
LyNJcs9so3932lLCP+EG7PlIHN/Hj7M0exbfUq6TYZ/94liTI9CpD4w85s7hDbgU
qgDH1A3ha4nRT0kBFgYOii0ZrPOAi4rK4/kBV0vuu9oQwUKsBsfCXkWHPC7TSFhN
RyWK8uJI6QkMoJeBnLYsH3j2f7F2TDMj10yoObX43kdxovRXsQoT1VWQujvaL4L8
W/A1TNNAQX2SuTQesE0rqzGZO9p3OZjbCCPO3V/fkVHGRrPl3ggWbW0nWk5YVmLP
THgsgYPRbR8p93WQDARdDdwIlMBPbdu4VcnQj1/PrKGyfiVSn7W0ETQtEjuwAUaQ
xeFZ0v1CaG6DCcpwa86OY6aWGwvsIgam4kHg86AddOkYJTBmhjNhtuFYX3CCXhVr
HQRdP/gyeQfDJE5EVsc9643wsTT9XM5JBSAb7S+yPMiM/Qy6Np9UIgCMZR2nxsW8
uTJfcBLmzEoQbGc3kZhsbY/7glBY+PjnxY15wyAkihHnlsY59G1xtnC7hZoxQw5L
RMC7ceHzgB0OAF5Xbr8V0Edv5i766uAgY/s8swH96bAYjvYU+qP8OQH/JOyRVPi9
iZHxyh/MNAbOzpjUFhnB+oEn7Iz3rbDsiJ2uuBJ8iN+GNZ86tBD+yBzZjh9Ye+wm
T8sMQf5Wlij7H2rFWcxQ4EHt0MwE6GCNfKnPK54B7sbJDv1seOr9tzblyM7Mf8U7
/3vHYCKswlKSsZc8DLyMamJyjbEJALPv3bM80Rm/YLJMZGjXBW9T6BO7ADFG22UC
adSuHN1bsEcPMj+mO2WF1Y9fO8uQVHI6aQcBWnMq0u4yn7NLIvc9cmhtpZUdale9
pYP92sy6t24m3nzk8WB/TggAmaRx8cEAJNpFrl505oFw6MNic3m08ZRXnZpK5IWr
L+9+8xNPal8IDausulBGst772wYfLNep7y8K9VlYhYgqu4cLWRFG9txlUB+Si1EL
LhjSDBRzBy2QiRiAOtEnF0qeIen08oGms/UoccKmf6nKsOflJhGWHngFVJejuMf+
GVWIIGLnIxNAb6td9fryVsDHpGbM2B/N4k75pF+SqZvm2CadzTnwY8iQiresa/ho
jgIpw8lHRFlDdncuqCmap6SrYL7kEbbZA2+gC/rlouEx/GOpA4ZIVXyzr08xn3Ec
AyUeLfuaZDlLhltImd37TMA2MYQyAy5aAN5FbSQjTgk0hnxyZXqE3uFi+xRqD4XG
2cFABDgDnqx6Ljkr1KUrrpylFRiE6G/dksH4ORJvuu1tATevpHozeCqgRaRI/0M7
vbaK3FQf2k+14s+1oiYo+A6pN/xF8wDfS82NQgJDyWtgjehTPYMixMy+n8QO76t3
SbN7bIDelkPakKBuUItmIFm/pzuOXO2IIPuECNbP7oljQbVunjA1+7fWgB03SGEt
V2l1jWo7tSYcEsLwdD21GDnH7469niEG2OAH8uDToF0V0qOGNfsMOxteHXR1LP8D
Q2z9vn+G9Hvt1n8kRBnDSYDL4G8V35/5DoYi4Ywu1KBCnBRBeVz1GALLy1UPNE10
sAKbfvRd/1xWPjxWykSSKItoqSwNumCbbRI22//A5MdAe4MSs+TgRT2csElEBiED
p+FGQIimT2VYj0mB+VTK/VZB0+igFNVR1XwyZaXN/kEMW/QMW6sVlHqlw0jSK1wW
ZKvKw2oE/2OSn1ftBidybYxrPIWP1vh+4fvDq6xyjza8SbO5AmMObtXWgArdkvyo
UvDf+Uu9vDdYyMy4s6IZQiAcXoL7rE4OYAhEVo5NCfZyc2A0hi0WmvuQ4JdTNTic
16bSV7MiCR7O/2MSWLFb1acSediBUk9uLBH0axjpfMMkx6gyRVUg9HTw84KrgHpz
iikzyHrpJRBzD+MoTNVWZMo0S7uvt4gA+RPef66cVQ8Jjnwxjerdp3jVydUk40Gn
ixJiuwSISPeMuw2kQkCLqS0T10SqVrxGtMnK6p3qrhroCyXavh4wVk29RnwH7lz7
5YnXHCSkA4LYkLqoXxr9O+M5b9Yd5wves72cC4C/tZSIcdIohnPjkMBM2kZBi6Nm
NjH7bcOFlZnsFwPUacXzKQ0CNizbAjSnUNkB+XJZXTSadLvCu4ImXxo8qFl8WqkT
j+vzQMJYzsVbY9S5P4QEYyNoDtizogTUa6m7/ABNcaSKO81VjnJ2IIT0SRcGi1aY
4PH+PPOvvP0wcR91+zsapuiL1j8IzOMp/CpBABM05FU550BqDZhgY5/fj82KxKAn
U90oJpqahrEOftehHIwX7EvwoVnl3/pEyWhI23CdGlrnFauwDsjg19hdN4CuZwYR
xfQBlb3j/WPw4Q4gVk2ADy6ke3kEoEdj6HenOjwotbgUMgAdY2X+OF3cwwCTtbxa
7jAN/Z7F8PGBLiLKboTwOtFc/pVhuAtrplgPiPz1yoOjTUKW+RbTynrGqfbziVeh
20HIQA6gwUHXW8ofnTOr/Nj5Cf+etp494vhYzqPdtpKMtID770l62u4LMV7nLTpd
Tdyqj1HvIAN+kgMyDVu1ynqXjDpKzmT0jAW4QBfH7Tm4PlyBm2NoQKqI+AuSZp6I
V82H/YjZnB/x+EkaEnslclIIZhVYsIwzMnQJL6kwtXyc0WcIsSrpB9wImk6Orxiq
PAhQrghSRU2FcTczoiwOaX1Vcs32QxYtldGfeg1WKwqzjsYHQC6ojNBYrUQ6nG1e
fc+KPCQOKIC9oAo1D4GrU0S0m4C1XCqkccR2cLjAW3Pzj3Pzo7giHLd2Osmzk1Hk
6oDg5NEk/laKL5kj8nK5fhDP5VY0CyO+CyqtbIVqfeLeCCmi/AXhzfZSoZpoVATc
qNgLHv3pkVmCZXYeTqxuI3XVFv1tA0pY41QixYSvM8M7UIx2YF+2GMzv37QBnOGN
axoN/QD9cb6k0SxO0PCgo8anvOZfKS6qZKwt140xYFin9n5KOL6xKUyxjDEzX890
GvykLnRrGhYa1r7PTR3V7fGQ2PbvNBmaBjQjLyEKZMATtJ9Mlf+ZZ9rKT6AQzqK4
FZQKgJF1Y8LQsou9SadhmhBbnIDWDHh6h380iBllUQ7C2whe2mXZEY2i0aSG3Qst
QU/5bVhHNPZDfnSaRz1j6Ac40WksYFDEUAxWL61ZHWpY8LFDu1gH0d1nf7BJNzt3
dNzzZsSWxwCQVAn2pDcbpggPwenI9WQDJPdWPgwjdZYGfe7jwShnmI6nYdJ8MNjE
046SS7Tmp3zXHYqAdo6amqV9j483MhaSIGxGbu0ACyDoFzkY5VxWSfqM7kbXi3Y8
PaIXBdCyuFThcx+LaqAOCZBGBe7fb75a2Bl2j9tr1+r2BLSw7Zh2PGLKn6TfMC9Q
yxxwFoXN/IDnNxRYnEVyJLtNmKP3yc/gAHv+Zak+z3Q6qQ6TxZTUjvdoPJRYwWsc
S6pQYEvqCaejaZLlzX7leFNCUMZewo6YwDn1bmCsMI3G/iELCm8CmSyRg3BTLouy
XXBtIKt7+EaC967VNU7dAuANsVKth4bJtjwKbLbdMYulSub3Jl0/9socA/NoP7bG
kihqUwf34DcvmxQVncT2iLD4lcsZbWN1tUTJl4FxyqyBm/Raps1v3/d15fpb0CJY
SAhijWDLkbNpMzBLZ+IHjBl2NFa250onci1T46rY7KAbMxBrB+BGtEV98l7HcK/T
YSwTcVXBsjc3XfleABG/89rSNlgnGf8ujAoj1waMpTtYbh0kUz5Ok87F79zS02JB
/Q5Aj5z9maMo06qrlu5RsOfOeifa2JOraGnX9FZODqF9nzDuI/Rca1jFj0yg1dqm
jRAG6CxHX1scvwBuZcC8iYhFgr6RUy3PKgUYzaktRPit5ar8DQ0G4kJprJ0c85mn
SlGXLuu8RyLbWEZCOxo9D+eKcw2UAkLqnpCY3FtM6lbjXS28t5Qin99URuf+55VP
rBzT5ifxjdbNTbX8b5Hjg+2D+We4K5S2+08hOKLEGls7axI2+5Y+Zq97GkGnfiiO
QHXcUSaGPyvmGt503KSxm4gZb+imXQTu15aIVL/XfGCU4GWTCVhUG22LD8qcYuAU
1JEkAYCk7IDWmjPQkndFSFcL2iCQhr5TchPU7afyOZictA80L8zsGZlfTZCKnp/j
gZkTIbXVjIXGIl3UosMO3qv5+24Aq9/KD/SnqzkbswWB/xCLyBqiHHFT68YxxOU9
QoA7xP+cg0sheMy/uTOsSrhFitjDXe+dmFWaqnmuQ9zwkGu6Ou6+co6cQzDUgyND
BH6bJGBz+kU/0F4aJgrvKsX60PqGgo2xH1We8EkMLrBSODgJye0mXWUGtVMOevQY
OWVXhonRvatF5JPvHLh+c4bTNaE17tvJTRNtY0E6KOlQXrQUnPmZ63xcNAt26ZrD
ex5h3fLAmIE5uz9acCyEgnl/UcE9Rd1yEw5+FKb1oQ+mIFuVzQ/pUgpaP4dHLkcT
9ez5s78fW1kcvbBXQIg6AXKWT6RG9bUhx7HKyijvcTg5FSz5VQzO1WYjChOeGCr8
KnLyUh4V8B4DUCkfWPrKHnvLVj9flNt+ofdSaccJTYSqCtociKhNjwzQBNfLap8J
e5L+UqvDCqkKOAjVC82iF16Mn7P13K1faYwlMIK+eBGbkO03Fd/kjGfyGVRQz8U+
ernnLa5g++P9TG6cEHR75jgT5ao4GSBH6z5OfMj4BZmCGL7PYy/Aroh/p++IZANy
KAQt244mfc4CxWeuNqsTHbNj2EKMCFpvoVVa4Yt7UGRQuxyUr+TP/XHCZiV/GVK7
HrJsDbYcCUAwk/BZzVjDuE/h/eWixsHL7Or3tki7fEScHT9HGTR/WNt26pXgEuOm
K6vNI1MozWz+ngo9LcFsEgnOEAS4JK5tDCmTOv1xH1V1PoeO9T04eNcHUqVUK2HD
IDTmvCtepyU1IcTACJLGOSErKhXX+bcKYcCJO0gfKkrASaBz+VcbqPMJGzNRrBF9
FQJdMPE60m41RnSRteYMMQEhGxZCN6NhO6toNQn/DoNIZIf2Ud08Rh+RbqifVCJr
U1JVEdHm0nXYRlisSED9eSdE9VbgxrSb8eoexxrJFVJluHcyaKgSCO4qqUGQLpd0
EwW8HR7be87D1bmJE14uYMKDpVOt/n9z8eodITMSyNxP4R6bkj17yli6sm2G9ouJ
6RAxN46SfsMw+eik9C0mRV3r2dvo0qXU5jjur1Pw2hNrZoGcDLA4tEv+Wy4yabEr
R+7QKKWECPLoEsRxP6aVynyryaS6M2gvx64OjJOce15aZytyusBUGbajZnqhw+rP
OynsNc/c/JRC4YQBFJ8TAcIk95l9E2jjqSoFuL0AD5QvJKrlZ1IPGOvmAuDQEC7/
Bz+zzZmmF5ozK8Nh0HzhsiMAmFaoohkKfk09zFjbHDjkMNTzl/hIUlcUixgcEmDA
jHfy+cZfaFG/q57yJs48a5s8SFts4v3wIa3Mi+igNZiXs0WMVT+RIaE8oKBS07kQ
Q17eE0RRJdEFezzOpPcTi+LP1nbYgRFm/lT0v7JH9HmlS7aP+8GH7XreHNcgUKPQ
teiXa7o7UTZf+HcWqpp1BzG3wEQKeUhHYXDCNIqzM4nCkUZt77BYhUI1yvg46XMy
MWIhmiDOZI3iMQLUAclpYFT8blwViTGcU3B3yppu/1xukn31wXIBn/UlpMpgBhKL
fFz/0s/RauDxckt1xWolA/ZIV+HorW/gxiEUbSVoDbdHpPYNyeL4doU38t5bDGnr
gWD4mKvyAk45EDdynTEWs1LUTglTB/dN9b971hySIgLTZQ+BVtcDqFAAYxdNIq1s
s+GmadiihjJ9J+o0CUB4zsniUMK3ZHlZIlEr3z5LY6rQXz0xh4teUa0CQwFMMztO
v9JyXURMx6rBa3jo9FUcN5jBvDjr9edAv5DW9Ypun6/05g4lQLcBGS6425eOfupa
zL6rNlYpKjn+h0Avrq94rFpS7PL1s9TY/DwseN6PtnWwhe2JhyhEpmyeqWbWDrwY
YuumWYuqwVI8J79HH7sXAgdtE6SbzJgUOevo6sM978S+ZrfXwhCcmYiC2aIYsAat
iSDKz4Y63/o78li4r+rQwQjptwiSvefY9YivqXuMKE1+/N+ImSaVHrSM90WP2FMS
0mNKf6L0eIzHuGlGfzvIATnCadPizVnyqHLo1I/0ASdddKfjdHopsAtiS048xpAX
SOygxBu6BcacDM/aKv0XQScKMihtL+PC1cqY1KIU/FLct2plX8vbJweGqR75/O3t
fTblgJFqjXgfPmnx22YzzrWLGUKnmw6PeN5/8rPd82Nkh7zYoGbJrir1piCKN1FQ
vAn7upYtcsyZEYoJFkYkxYwFpJB66WFZngJ/4hbMKASZL/Na3aCqUE1ZjgmXuUVa
BlItX8XnHx46kA/1FU86h/DclEy8V7+MSB5DtYjF2zDE+kbrMum7qZ5uvpF72iC1
FHwujQZ6mXL/i06notCXR5P8FJ3LTKHJ1OJSdYH7MNeiSc2ZI8olkM1mrpA1cQwj
VonnxSC9YoxsxUOMYR+KMdgP3c2x/DEX59Zur5KE5xyNoFlh7BsDokcQ7ANnzg+E
GL/Bg0Co0eGkk/MtCMrDL+cfVl5liLNsDxwsn21Ls07w4A2sasvjm0N+kEBPKnUG
hm72zHeSJFv3Vn8/L3lT5euqNcDMCD1E0evqzWK9ZWmzcqzt5uq8hnWaQAXMPo9K
Zmd/Fpl2cPkGz3VHYkizOiNZCBCgNjaN3PxzDDrS2P1K3IV3wZqFl4zB/WsSfrwk
NwcaSAAAOcxuaIbGqzUNn2Vt5TmFf/uUk6071354bWcVyGxGYVWuuBrWIrfXF53c
kwDgBxyFgf1JIiBXW/4biPmw3qO+Nxe2smG2EGIN3AX3460oZmAJvqrSlqj2aDW4
NjA38tGM+IT4nlpw+amAjuy2diwjYDcaji4NRlndI9UMfgKTgNErd8kdTScWDtSB
ZuTGpKNIExyVlQg+dWmAE4mgAOdE5mxi02pZytGy9kF2NFUIWjfOdc///qVnsDoV
TPlafolZfhzOnwf/tI16SoSS++PGrM7rB18meyt21UpxS/j/OeXWEkW/RRrCTeWV
76eGNhRxeHe48oAM/XJo2puxXHAaPbnseLovxYDiHXxCziqd8w3bWdShGLCC8SJM
WRJDtapUETxaNluA8iE+r+02MSG1BN0BjbFRrwu0+e1085R9D45YvtZ0D2g0zmZr
ypSwj23bYTLLKG9Dthg/0szVXmC0/4SHCyei1Ht0qcbpREc5yDJQxUDSfO1wAF05
YeUfvRjrD5iBVorG20gR1ROyIQ2vnihrn98HlfpRK3kaveCRZ/PdVIU60Z93FndD
D6VRpSQG3IpYJc06xX6HE0dBjMa2S5yT8FZvuClh7a2m5jbV2XCXCO+nBma3j+yZ
GpHHi0ucmcnOloGt9eC62nsEMex/dZgJuseMPLGCi+/dFmxrGecOLms6gaNDEAW8
lKS6J9iY34xdF3T0MPquByWDl69nNyAU4D6/nEX1TUNA+sykovge3exC9Cp+s7C7
PjUB+t6e7a0iwxfM/xYFpeWfKXgHOOu6t5hut2zzlK+cFtnwD0lsfbIF4N7k/jS3
MlOTgm/F/IYZE+w32RgQBmJjASpQm2VddslbK1c6tmho2DKQf6+ulr03WPZ9IOjD
cQ5qhUEnsN1Dw8nOoGUUCU8sJZnPZyavXr+BJw/Feh3HfELqrFLvMsdSDoLAeiGJ
6EIqb1SBa8+4/ZTCXuih5IszrQujnnLO7JYVMgPoQCE9MjQ4BoaCaMg0SgL8Unhq
BCBdDosFyDpFPYYyso3O5iu6WP9echNNa1lSUx94mA9n+3PLX7z6ni+Rc0YtmW8u
BgpaGcOlb4xE600hik4PgpgRytr9Im4l4+e4SRLcjzu0wTDQUB/BAly53ZXGCZ7D
wxsSfAHqvVucHt3C5hUYAMnZ3OPJ1r+7S/Dv9ooBClLIuBAzJP8njSggIUXJube6
lfrFXd+x2ciGbR6f2wVH/aSEHftAQpJL3RRNR7gvd0lshhWfbpqbhTlhN3yItywM
UFMZQ5rRzdxpyM6ybbbP7XNE1seE/VG5YDhgBSb5Uo3NUuxQYVHz/NVtmzI1l6kb
QMpHnfB2C73pvGiA1eQrKaALpYVP7cLO/cZsB4ZKKlxKti44yZd10Y8sppvtDUIM
OlnGltbbNFQWwYwql227W4JqxPNHQT6kS6UzFNkAbO11Tfx6bwPrZd7uuWewLhLH
76ucs/bVy+9KZJQEoeYFejGI9T46bw2fPgQxGmCbwjZRp/s0Bb2naGcRU1ncCD1S
7hclAFqrLyodBpMsQ34RWdOrTk2icvAY8T7tRKNQ1GnJI4M+Jl8ewoxdHDMTjEwz
7PCfobW47aTkAJ6rP3+7pfXkGVBVZ43klxH+zZP7jz7e8/ACAo4jfQLgpiE4WFnJ
ci/ykDoOfEVly6cshBwmBCZWHp8XdYq9RkwsD9I4cvpqWvlSKKKiGG3y57b84UhY
U/bDwrKOcxXX1pD4HGSeD3NvQe9S77pE7kCjiuz232gRNg/5soSxWaoXerRboeRj
c4SebRPO9nX/4HAEFSBM7bJCHNWySFtrSJhEhKMIanZ/ApCtthyhAtLLHz/sUffm
bFRBALSwm3TVjehsab4JYdMl8ZTdOlYUbIxSHW6GRJryEr7R3aJNNb3m/sxMhIJF
D57UH8DMTNgsVQ+jhMkrG/O3M9ovz0qk8/r6OEAA0tU/6XeeaUsV3yOJSpvjvB1B
bYMW11Mivzts1O6s/2wrSB5rzENWe56ga6GmWYuR6PIH2Av+cCf5/BkHWw+wDire
fD4m18DN1Gahb/MCxLhmUcfoh5/0+YeQzo9Zc7JvUmxcSJcA28UvvTEdcj6XsU8U
YScZHMwKPirIRlHEqPy5sHrCCDhK9/F+dWBq0UoNpg2My4/6MeX189DsO/r2Ovqy
0o1kPrQdBQ00tL8GEaa9u5bowZg+cs1WuKELKUmR9yjLeNPABLBB/pmaH2wKA9og
/AJFPf3Xuggvf4I5xIlVnuOcNpEQhiVjs97I+8trRzDlcb/uvvoCLXUHK+Jn/hpB
kwENeecLf+bkZmRkue7zcbElxwVDoAsqh5sQg8HrBC7gPl4dSTPnNJo1LEfEgh9+
dKD0KaeysSx2GPHsa/EEyBSc5UIDO4gGzDLbvCsu9UcfhYYZXbaD7oG1IG1S47mI
Y0n8uuTfSFxiz0Y/0NnEzbQ9pJZLWbg3+82bxdgaYhPUyK+oBy0c4beruvVTNLKc
oyLRBTxdJMltD7ruxmy/7YA6b/Y4YjrkdL0lzWA+nozdc95a90WnhZEXNOhri2Wa
9DqI9wsmvJfgKzf7XLgD5GmLtkcoJjjVwyUYxnjZQJZkvH5nocMgHY90/XuvDfCf
NNSiDr+07Dyi7FWzFa9YPg2FSNluDbmmuUzWqucM7LZ5jiOC7q1UXatpxmDFPRpm
RsqBRI0foP3B5NHpitYCapbWLM9eEpCvHtGTGTsBmH2bWO806KvDy/lSjznW1UfG
8aPzk3BLW7ws2HsP6Q2qq6OWavVRWPdSvgfV7FCBHzgfYMbdnnURo9UwqimBGPpU
wKrBFv5J8avfxoFCps05YbQCO3bqVOZMhazh+ARenmyChBrUuRELts6WGFD4+ib7
rFEp1lqz6hgXLR78yYkXx8eZb711e+cBrhX2TovJVzP2tfGK3ocXGGREXjbjrvAD
AUkULCO3XVRREVEDVjmH19hyihuXuftJD7ITCDUT/eEWKC4bxitW3ykk1iuunzAI
BqeJ7c9BrRZ7foywnfkRnkhma9VeTFi7V9C3svNqRvQ/bXs/URVmOe0rck5chm+b
4FoeASLGS9XcdrVw1dkKyCH4Mkr5Gn5/xkjUuAJ9et56tVLDipiK+fqa46OkCj4f
UJwXW6jQWseSYxmrgZeUaXTb2DWt0LnkzbPEtNAHHKXHjWy0k8HeV2NtzFMCkBMv
UHrRyNrjQ5ZKSjKsMxCDfV/FSWLeK2Say4k85i4UMQBiENyxiCKrKKY97trs1OPa
loZV16JXyfbtsJJaEK6zhQ6K23LKzW2ndisSe7p827ZnKoqop1aYxJCn6lo3sCw5
ePGZuyZHwUpr+XIwevtjqoNMKQduj+ZjVuXm3nUutYYXARPEvv2syvG7L9oKcQ8L
P04w6hZUwjtkKKENS6FAqrH1EYNH202Jubl4QHBUQWn3hlVqyhI8iGSEcBC1D+8v
uKNwWqJkXVPt2vyEhCk9YqGHMR0XqU6J5/VTTrFyJhya1cKiBZ97vswn0PAMXvYN
u1tHRaW4xEX1ixz549kK8KtHdbm5eq9cXcOdvNGNmcqH8uLxLqHoHybIoEZb9N0B
9ZoWmnCFtvqrWUi1cMK0kIbaaove3GC1YFRr9DbCTXwNgx3/OQwMpn9jOGI/IxF5
7KU7UEgWxDO4Z9P3iXyKskn6mU6qPWsZdgRgBClKWCapP5fRIOiE68EZYTQjUfpy
RRy4WcT/ntfL5RKchLhPMa30iustOS9PXTajq1avUxJAx6MAidsPpeH0SdHwYVah
GnipsD/vwyXKSkAw0JFt2/DotoIFLV6QOnPJm/3inD9jo6c142+wTJf51rLp6QOf
61bePx9fvZf3vT6rTPvI5Wq5uQG0r2xQhv2HIZrUMT+dWvwYMaahcLQXe/kReAM7
abeoTsnMFrgB1vBLbvlfbagIZ8WozTHZVvGbgxU5dUQU6TyniQZElVzRLh7uQ5wF
tSlIP2vBzdEg7UAlU7gAAH8yWsBY0RhM+fVKv4F7RbIRXQM62gkJC9nNWZ/5RJgQ
sRjZmoBhJSc8Uvtii1q1q3FmPGseZuustN3Mu0eQrHzU6PjSCOf0xN+I6N+ktZ8M
18VU6TGtDMfTeGvQShW1UWYYa21d6qDlOeD4uEC85/usJvpA7RlIvV2kAVJFsKXE
vPQ6AjjcUqtjjM9Uvsl9VhGgIf1KWxxy2XRVQpRhKze2s9t/MsfeQopSJg4VoYkV
J61yVFNW0f5myvM9zNnMrR/LGhroXpN2ZEWrS7pfk467749S4/vbM/HS1/n59WMO
azjlyqEQWLaJdcF2lXTvbpwBlAfCNfC3z3n5r1MjxF5PlyDXimTfHeIBQJxaKNdG
FZ9EdKhH2tzgz8LMsEijtyVjI1EYU4Mb+Vyy+tqQBc505OX6aRcmy2wBFd/bg18X
B3Ojbo2sMZJNx/uEE0Ex8RRw0ABk0+7prmoObuFP0pxR3E5Zhbc/5gCBxICgA6eG
fhXl/amPZGEmoyHaiP8C8tjoHnyxg9LcGZuoAwcWX7dp8uzOZk1JylGjggYMNZ3q
v4Bi4yv/G3LRzySaLaUataOXDZqeDL0nUOvq28GqVlO4nw6dnAIk2DoBQU4Bv4u/
9/8KhNJPy9T1iZ5Aab6LydETq0FIJ7nLjICQrc7vmbEB9iszwe7zG2akx+XMPOCF
DuqkJaRau+9LX0G3gpHWJnn0wXqsJv0h7sqV3eTD8Vm08nQRgYeO7dpCkZtpvYTQ
sxqKCMEwxQPBhuefHmY61Gruu0rqfhLz+9tNA5+3ghGehESqK6uxORetRmwDuuyc
Z/0rgx50rnRGF6C31bo8gJ2G/RUHYh96XSy3W9qP/NDv0MQna/rFXjHSzLmlf4J7
r4TKi97DJmgbJ/9KpNy7czlj5TSaKYHGcfkDLB1pm8vVMF7PqxEAai9J7TINCXei
+Bi7D4/yGx3CeJEAHYd3a6uwEen7SCitmkI9LwL8LO+kzHcIrEWn3we/TNY93KiG
+/QYOla8XEEnNFNQSwBcJzzSdMGddfycYrFStSx+QBg4wYVG9VEUqrpu4e4oeld5
Jr1bWGx1WXVc3N9k/xhWyDBtCwLSoG7YE81yWXuVm4aM0INuNbNeeDA1d5BLXvBH
sGaBQB1+dyto7OhlAYsZaCgsIcDvbKpLWzzCA8ekgFINqQ8RGCSodsXZHY1OUy/k
XqtIc6B4rfGRnNuAfUq6vBKkcitln5pZ3H6lzMmAA7+Pow/AQfaECeD4k8loAAs2
Q2np6Hm6j6JUSnrPAonf1szZ9O3u2aiVOtqgC0qjIVBZGIfIkWjd3Xd15XaS8LYH
fKxvbaYOwcrL/zKB0zsojRPwww+tXNo8TH7j+2ZLGVE6sIp4QuGbwjnyEz9XSWht
s1RSVLHymMrUUto2JBDMRm2kDO31FxU2aLlDI1Smsq2S+Qt5natYJbikfmh8TWim
hWeZ7tysiolzdNK+/+L5P4hkJZP2kMV5SAeRtcVvnKhqfIJZL042s20kpr/9TsS3
xIiJsBE1z4GzmS28NzFcUx+tb9j230IZkW0S/NOp1Fj0WFlH5zVSHOZkHpCTDykw
hL1t4vl4W7s19B6MsyWzQlyHTMumt3YOxDooR7fV/DsM8S+ma1JoH9qQ9JYUB3mm
BcDJesEwl51xykRyRbPk0KW9oYQarH1tYumvDg+vjFBlzf+pHQXYzUDjGoPEFnt2
N9ixVtOKUfVlvT6z+A+LUr5xyHcTHSvYIflvjWToguGuad9ajwZfe2YHSWnvVWGv
RmAeiEZ8g6BiM2wadazs/XCh4lpfsOG1I4+6I5vc/aN0hhPQq5L+yYgFo+/vdKy9
gjlk+gE+i+cm9WRvvrLLAdhDRm7YFDbeIi+56oBVxiitS8LmRK6tJQ3BYeQinugO
lNbb4OwPj7g5POEBir8cT8CalN1LA0n3f12vitN2SFSkkDwFYX+w0bRCpaIOdHZT
3fERxskRLyI6Tdi1047849ikVa9Gz/EAuy0PRMWZL4d8MrzrflQOyfCrnz03Ss0o
kblOXcdpzHN0EKyIBV0YE4rP3UY8qAZ+WnYbhBicu3QiGUZNrjWNjB7XPBnGBMEG
kMWxjv/TXPs07hDxsyy7yWVsbESOmteNvFLkjDQ9yKdVxVdTyDVzruK093+NIl95
mf4cH5/pVY6K+Uy9E6sTJDO2TU8dssS6h2YQMwFsuuXhyq9BJ99FTnjOdffdWzxf
R+SxTOnBSwt+Mzwx853+LE4DoNCsIr5NufaIKchzjfHNRwUO9JoHiyavkrFJ1A2q
40AhPOkIEwR4X38NfTlNOuUyvRjWNDvezbCb2FhEzdfregVggIpIxy0cvlQdKDeL
hOobVQLcAAbY4TZNKyC8oz7vY0GO9PR4D+jLRUngqgl+4EuxTrbzFpS/kdSP00m/
woS2aJJLLXmB0OGwO2a0a8OFvGa+fSfRZnAsE25kA6DURmnuhE7BseMKmuK0Cev2
fNRT8RRqv2bCKZKE4WckkFj/7as+0AfUKCAUd9Pex9L2Af/gVuuaoLadj5d73U/w
kJqGPtL/m26XoN4Z+0To0cAQ3JN6MOecTYUx9/JeF1VMZyovVR4SztyQDf7lJVXt
1tQEZN0q43NWX2iUxNRCmhcbEMN5D6upepXRrogToqX+ADU7AcesrMBmruJFezNo
E/Huxau6Tc/vxWNgf9ppOwVLfNhw7MswuLyjKq0YGWiQIdQiYizEPVmFvhf1oQiM
y7YhnQDiOcUYbyLP4gO6LGJ3sgAhsJhIqxSqY1CBip6Aslr1gl+J045/Ri6wrd8O
ol6S26rXU9TBAns2r/9X9mXlni83HBk1zcgbDUfkySD7miG8H2LNQEGnESm2ujP4
STaEQniyZSPt/0oIsStRnucwyj3rEAXE9YHlUCPpLPLfpNus6a9FRYMLfciuVid8
qZ5jdQhxTVbGwvud40nT9tkt1PvhwHdoJddbaZLOjJNLncQ7zrcnm7XcTDu+oZcm
PAE37Ro5y3nSD2uM8dh0/wRFW+2Qal2WGaLKzNb7u5uaLNoKsKY1eCK0tqIvMwo7
zj8rpS13mIq15E8ab/YfVpPBC81xWE6sZPsvvNPISA/hHchpuUAUN2kvvIuD0Qmn
VdOE80MeE+ApRt7Z2kmiSQU4egk0RJdfdeuvRJGdL986lrovyPhxUAOCZRDRK0iR
97f/AYSW6oIV68T3OulKJcVIJs494uG8QGcSflXNcjYwoTexZ0enfeytm4r6C6Fm
RvE9kVfR5KYeVTv+tJm81qJyaXMwgEl7l+/O+NlbiO9XuHqKDSD+hKBX2ig99Ct6
Gg6jTlJA+LXZ/+E6zMzjWbsSesBtgjSXU+CeDpLuzilFHEAmmq8Mt01rWmhSxjwi
Cv0GtvLuHoXjgXn0PFOlow0WH8l1KIP6lrCA/4U/IJq87xMQXRJfdzdToIbVwfcl
QVZcTnSwPgpvRH5Ng+ft7ahVEruWqbufPfJG6YWn3ysz00coseLeXm13sxx0/DKW
6zNBhsROO54WtrbUwfwXRVEr5I8YmMkoxJ7E7g+45dlPdRj1J6XbMX9ZiZfP2PaC
QjNNr9Z2xqwInRY0r1176Xp7hsk+K2JcmEavG++irQ8IaSHJvkUhFSqZq180W1K2
Yg2PrNASQzOr91KJ8oxeN566rHDblhq+Vu3oIjye15f1+2crJDnH7CATLqc5gNXm
9Qwb+5ZMym90dXPgQFrVRtKbOCkTqXJTEMzVXGq5ldZx+NRss9dTaUB795fHUKrM
2jXML7RcBam7Ztb5jgcaw/JD6/YQDKJ+dyqVYHnLMy+C20wGp7YIin88RyYGjiEl
Jsgot47+RM5Z4T02ho7WaarzgMiQ0MQryFci84qwMdWALkKEGueAV/Ocz0j22QG/
Qk+muf84nxh7Kc6std5Ns7GmlljCScdmFg73zZ2cCXQlQLv8XEK0vz+EVV2RrxbJ
bJSdHaVII4YiKKOb7MFH7d1gIM6qeFex2CBPUC+wXEHtya1iNeidTp2PmY16DQ+a
+tYEG1XYp/Cjq3ElfN4ZqEZM6+5nVyeFa+KeIm0Ix2fAyZ2JD6ejed/CEOetQLBy
cjEbF+V4aCtZM+WWV5GGDAwjk2xI/15Y2oZfb14IuVR0qt7Zo+oTxy4rjbUmWspN
lb9Dns2Bj/cjv9uzV+Ox0bUkxJmkIh2muPtAB/YGNJne3Q5NLg4GYZxxh0ZsVHxp
+D2u1GGJA5kn89O7jMs0YFYOt5K3FaKabVDL8/jCRR2hPF16Iohbh320706JEPa8
BwB1tflARk7spHKrUxSRrYRr4Pyy9cksMJSe4Mqr5x5bTG8MOKz1nsgl/IO+DinY
Dbs6ne8NprkSg//Q88hSgvWhbO5E6sze8ITOlEEm7CgtzBv+pwFKt4n5S0sjuGJb
wRoVbROQBW98zkqcvXVOcJNJkXEapGncd7Y6VgUpDSXf0H8LVgVRwKissS5uT94A
OMmytqEOwAbdQcBIIBZawQdaMb88Bbgx7jvRMJL8TZMhe1fW0kK34O9x43wRqvoz
6v382JzOgmiE5ir71Hd1da2puhDMpQhNz6hw5e5wOCuv/sZ7pzJ/tmtty4lP4rW6
8MpjOWKBRDOp9ygZHO4MkgnDX53QMerz4lRYaEtwhy7su30XUNplWbWvv+cCh6U7
p371i+GTTWsa79AalxTrc0o4d19zL6fN/2ofNYV7HJ5yGHVfc3Afyqg4wU4Rva+5
lPPIgUSFsGgbkbgnrcTgA/cV0AqD5nxN3bOlF0Ie+oUg2tzXtryEVb/VgcPTtSVn
m8IiJADYJXCrrzPRwJ64Xvxfkx6b4fiWYopkujpcsMSAgFISF7Bt6BRv3GIY4yZx
VY2HenwGft7qrNsBIBKreSrjONxYW2zVVT7fFO39AyLP+TitJa3Yd9sA5SunsQeE
PqWpJqD//0lPjio1St7Ap3FimMmpo66E3G3AAjAym5BtEk07PFJem6+6BHu3DpOZ
eNpQxrr7EAZS26EjGXgccLg3gUvKmdHEU9XOfGBWDOhikeLiljHQkR2HDTXKntUv
kwMYwJ0eyrKIz0WNJ9JoglVbart3MUeZlKqI2pMrMfsZEDLi7SKSHlARDLMaZqbG
/LUTjKvRByXyhjwwUCul2qmjgGrtADrnVdA4hIs82JPHSX/V/Ww/F3J4cg58BZXO
8+Tg0mUC/M4ase4UKATpjUaDyKrjm2u0QU0TAIdvSblO8kqibIYsgfMQCHNagLXo
SJL5GgY2h7InKDSzG1w/zFmiQ6WAAyPqMdl286YaWIoCeUv05D3N60o+c0X4w0Rp
6MhnujenyBiNo0DllQHZI//SBCds0QYmXyZxXebsij6RHkA/3uAczkGSsCyEHMvw
n9HZna1gk4cfOW3K4YKlAWc+VEnIkMoFmg+c/wrWexc8qt+PCX/gmE4VfRocJIIp
/+fkJm1zvR0v8kfewIzu/coGFgGT8VBo0vvhCCKjdbQY1ya6gNuLkrBQRWPRkLRj
PTDit2BclOiAGO+drEq2FFIejr5oSvCiT9niHltXZXgSu+qFe5xVhk1OFHjTbHZD
xOLyikHIbk7NR8YtW8m7fs/ySiFXwK+GSjHh3cGIe4uSmpuGG3bbrRLZDsVCyx9G
+2TkF0ZyukcnxZAp4ZK6z68NfcuJ/Ofkt3N6F9KzpRkJ4pebZLynOrCI1qytbVPp
u0YVbAjjMoWgrAKLCPegeFLUIDrL81iLRX//z/4iHFPb80Ad1rmIVICbWa7Bd58p
11910cqbYfAezfCnhkXldAEzeC/LzEAR0fAvmw5vqQbGWLR+KK4UTcIXldQntvq7
5v49eP+C1TQ+TcV2BV7w0IKgtf8kgaod+2I7KL2PKIIKEijdCzk/lPpR7OgGMbaM
RMQKP8kOCkIq+XBVA0fK+tTxXDHhxXoeML47uSvtDxeP0/jn6JRgpZooSu97dwIX
B0aoRWsqdpDJ+BFjueGg3z3gdX4BC1DIIkf/H5pDmvK6vy8/wYO6F4ztYJZeDOcy
5Ay04JwPjgel6MR+uEAP2bDK+88ufcCuM1WC7X1/iUYwkR8SBRdO53dlgTR+n6qD
iTY4dU0hPuuDKW9wYN1/gw/w6u3Tk27EVVKM0L7i4azLrDXvGXe4lmE2ss9CH0eS
9YiJOGa+YMtl5e1eK4ZPE7sX9qL6NQYJnBxwWfGhV9oRwyoWCtWP8ACPC66KdMq9
UJlYIosRvtACe4XSoGl90X7LoAvjrrgKdTQ/psdiOX8C90tJZmsoVAl2upUkGqVB
QiJoEB/3LycsS7ir32A603mXxmlZO/gWtX1uRHiFjSKzcw1gjIl3YhxihzVz95oP
SWHk1sq5rY09BVNs1TNCcdgaboiDjCC4LjfE31Kfdwbnfg7hH/3lFKHp/jNRUZ6r
3SEULzoPM68+yYjYrhFIZtzxgYfLSZABOj2Ti5g4aYXqCS4q3eJe5umzhQKba221
qP4kXqTi1F7obkN3+2SlXC/RKznvCQgo0VKHPkeZFpGcVbgWZBNURk0w2KfEYF0j
oxpGWrdDe9TCbLhAQEJbfHOWP9VlcAPLyoTrCh7ZSFVgdUvV9TQLyRcLPz1wN3Mh
4ZAvymmptl2PR3j1wWuT7zn24HIceqpMp8UAXTrmi9oh+nzrVqNmQZut1XZobPeB
rp519O6Tg78vW055yPiRFHjn79pP9/XWh5buAXUNVSP2Ij0jd0mRMT0NznunbbSv
7OFeiNJ7bEMAcOtMo9P7Hv7gJw5wuvUR95PdPB1bin7vmjhH1nGDSEpy/LSdJ7tu
MvZRKS/6tNp0I1CE4plq7FgbIrac2/2jTwv6pp0qNPYvUnfxnURRF/9T4zYD6syQ
oQQFMX3BpMyo/56c9AiYgUTCQU0D3om1opbBJ9mqt8mZIlchijb3s8BZh7xRD2Cl
fwdGLuD7hFb1V+FqIg5iX+uRwm17Y3jt4Zv7BQzX0uLYsNNnA7rIk7yb5qsVLRAU
vXi7nze/t98QqL5h+b2ph9Yv6fTgDCHC0uO+ZycCasSasaHFIsnwr4W/5P/qxxsQ
nuDyG8SDkzMfsbGz7kZTU9kUCJ1XiGWA0vIkaA3NkMAblwn5zd2LhYA4UpAQ+P4+
Rt1Ma1f9ZqyWpDBa/99hETq3Sse4w7VCP0sLXh6pZwKocGtc/j0LstpTAh16/UrT
KvFKihUGs05HHZJ8YdjpWoHxC2ssDhUXUiIU9hyAZoZ8ZCURxZIl/yy67+r2T6ZM
f4h+fspu2mLM30AJnn2GuCoIKD1lUXAdr6NZwAlNMy87wbLkW9n8q0rcA/kQfmAo
+lXZe9kMYWClsgXpOxnAyXTD63N+DHDM/YO26+a9trtgG4tyez2pFdmmUzpq2TNZ
DbU3DxtMt4CHGWxiaPK+GFi6/xSrRsbZc7pLqrgBhr07iTtX2vrbBktnuZix9PfM
7UyZydFqKy0s2Z5ZvLny2DPOY7hXqOVAKOu/EC1/CcigHbOeapdYseLprXzykhXd
pk4BWR+jLbGEr/LFeuo+rp0gZFI5oIkbSSMsRTqw/lKKRtFVPkGKW3ERPNLRfScW
oDwlvK8SJMa65oatGrMPn07758mYHYkNrgsnD8QnIdL/uJqu84HjSXkZcnMwCxHn
sN2aBMWdyeDTpwWEwtTR9W6KOgtN1ZufyQszcMB3nvvPMTV0/sI5PWKFssrRwWFe
2JKMxnvkWOdAye63byASdwNWeYzGP1MJ/wIu9n3zXPeLXlcH7Qd6kwaVfy9BiedQ
trhpzq8+6LImvM9AvcCM4MMERH8bhYEDmsR19+Hu66IPiGumP3RSsJBKJAfFC9fy
G3dpMFhUtjorbnZH2UwdUcLLSnIJxRJ8FA76NozseINoZ2muT0ujcj1DHRa1N7bJ
j2KLbq3elVjb8seIzuzELzV0jWrvKyA3ItiV7b6zu1FpLpU7M4bDRH/gdmc7GeiF
FfVqVF533YhrUPasRgXfekNLoYmPJfSoNqNg/GOb4Yf2wEKB7Duu9jmpnsTTpPaE
13dPinxG5aXYEvEETBFcU007WcGq2kLOQA+ezs7iVw3TRFff1ExTsPNTPPtIqffh
TkOOk8rk7SlfeF1WSSNmMRE/hAh3xCJkVCIwZMIBl+Jb0BYFtsS4ENU5q2bZ/ozr
UPYouOWrH2JHkZ1QlCli8VKoPH1LG44GzvlWiCXXn/RMMBrtB1o3K1a64+dsNuuL
4JkRpEBT63qYjhkM3BcRbMcbYGFgbx/JirfDz9E4OZU2hwY0GhloYhi+tSxJRTEY
li+2PiTihxJ+S4wDwal+XdP90MahQrLpjMNnJXMlfu58MkIgVeYL9Ai/f/IChTNt
zfEuey5F1SqmKwUHOg1nZan7WjTM6r5Vqh1u4cO87DFrUPjDQcxZoCuANqywANvi
49f7AIu0UKoHwRnqqt2SeIPBVBU9q8MNO20tfqeDT9qEWowbTROR9u9BX3+mhqsX
uAq4o99isw+CHhXjnxpWgOJihUBkVaH1CtxG/QIBGv9llRDMgZMHO2sxDHqG4sJv
Mlwt/fNF9L4SBzA90FqL5bpun3mJc+iTrnXOdMuzPTZW/I2SabfS1PPE+uyx2PxR
wfAXKt/tFzB8CG4wEYJEYXcOl3TxCB8roUSAgM1ufiQCqYp7DQaYucdrvh+q1zxu
oe1rd7a/aGiaTpx0ZCwqnsAcfxHidoEg6XnZEH0hCD2bvj+HSgPVq92G572+K6Mi
tadTBbQH64mJ/NDYxMHTCyTZSnl6dWUPc89OlmW3B7PKXQ5rQ/Mc/UZnZTq0ypcu
VBPx0BQjBye9SHemv6t03HgSNZPATUzxkygIjdEf8nDIr96ur1HsDzGIzlAKQys8
bUoDGyerpJSEjXzK9qMKNVeOIv5CQfrHRa74uztD+J8rndUam7xWx946NtUQTqie
+8c9ujDVohYC1CDceW0WUG4AomLqBddRF09r01lh/c0SCN6MpGtHfreD5d3si3lM
rSu1mo1cam173gOgwIV127fMqVWU5owH2yEADAhGnZYop4CU0TgzcztNPlq57/U1
HFCDkLnH+kMbgCPuPfJzJ9nd2ojOCrI5gLEOL+n19su/yo8+nLlxwqp4rX90jXru
BTa6Hyihk15xNrniuPKahUKfoxMZJ2BKO9N3E8qL7b4a9IFJ/KYnH+RIjhE+fOMy
ncTHt3iu5/QKFHdMKdREjaO29/owp2SC7em4IPre6ZmNJYCHna0Tha6VXWXCqnOh
TNTV59/WhALxbWN9XC1aI67NVudrnGQnewddRUcn4EOMZRdWVJuIeLVBoNpYbudY
oAKi9AYq1MMyKR/L3WYJKF49s/VKwrvhC/hbxHwN5fN55mWuevhL84AUiapga0sa
CU1dXGgqvf3xA0bxSNxt5Sjx3XxPezIxUsI8ppyWFnZeHa46CWrCDUm5fBH1qPNz
+92Ta/oqF26kD1wxDS5CayUZ+7/zaAIv3MrIxfvljHRKIw6MT5gdDlj7pcYYkKR2
BEV8BFmaWIf+sZfbfG8R84M1AcZKsM0NDuy88TmnBkdLTxia0tFs89uQI0D3BNrH
tvgWPFjwQBgpfOXXjlZgASr+UbwHwtwFD0Ou+3tRM8U5hPOOIquXmjYUag/z5pDX
4RgBXwNocbwtbNo3CQv0YJjnJ3b6uIN31YiQ/8kgionEE3CpWky2E5ziXO8ehJvz
SQ+jfK0mH+fr0lmoQz2fmtZrvcvg1QDqkzitLuMZLEdzYVuNa6LQZXulcQDJ2aTy
IogwLYU//Teg6SjAh4gPKoqzDP5O/dd2s2mbjE6inSfLOAipDuIESmqiSPmJC3LT
1j53c9+BrDiVNRA9lCVNtHH8aGD5PBvRdYeAVzog850lu943WtTd3hFvUXlFSsrx
YXPfuNKM9ep8kXua5ahZmyGU4sDK8Arb5yYjGhB5Vgy//79HI+R8T25J4GN9jEdy
bLjlQAJnlCel6ZmNbBtk7kVZ7uuYFsDma74fSM3LowSZSFmdwV8iXY6vVuUWY17p
iJhkiRFu6bmSL7ivQCXdqCQ2UPIEfW2UZY/UHn0bGZor/3uHM8+nRrJRU4i7GMRe
nx0zBR4MtAL6noT4raJ/NqJ6SV1hUzDCY+8KpGP7FYF0kC48FEeLusynb+A85nOx
RfBLywrNrUFWWRqYfRe4AEp3peytGadhmtm9FckMtkLK5hfhd4PbBgTp8F4D+2M0
+mlXA7Ao14XcBx4Mb2BfKJBC32C78zXcKAovKW6HBsawm6ua59rEUZ8IZ35My0T9
FaG5zruPphKIqMejbVK1T+1yAUsmiIfLFdngyxhFW2JJ0tHGB78b1WBvZn4ngHYR
2Nd4XFGiXJXjJ7CDve2lU9MlGGcP5+RVjlPVldXSpzFs/yo4F8cxcfY714feLHyo
ww8SU6mQ4EHR/TeGJsq2Gc8fyzZVMkpKoI6Gf9u3fRoDaLBLtq+8A/oRpEiyiSCe
vs0Lt7CBIT3MhE3bqMPyzJ3r/Thrs/zvmaGFqks2Swq1pGi5LMgBX2RRQN93RsNZ
iEIXCWOnLY4WrZVG7fk64rQZMsrt7eqyYSkrzgWviviTUmFFcTGAmEVnWidQ48I9
IDRLn6VOdJftiyokzTPNWjltZ+oYI7AktHBYyD/+h/xPKKJa4sz11ndIwOm0ggbg
dYPWXY+qtsRfdG6IRIblft7RT6nDCJF0v8Yxtb1QmfgdHePNJO1/Eo64c8qHqGqg
/NPq5/IRh2bywSzYeZifn0G+B06wxQikB2Pu3B9pPeeUN8KVwX0PZ1GL8NhH0Pqy
RBnfNEdvkj8HtxxZzYdh9QaCIZq3V5yknJe44Pr344IdSwbeqxr5EJ7wehqLukLX
lX0d6u/KEXtIqmiQmaGSw0yfA96T9UIdRBMo+aaVM33UtDKv21ZGghm0Hp8TwjUp
cq25pA+Sbk0kh7ipmQkc4wshNP4wEXcSrCxKu5TXXU+vVisw1af47ftPNF3Xe81O
oTliALb6MmcVgVf+OprGUGjjCPp5mPP7xLWYrBLGOm8ts3AcnPbtzes6yzlO+KDq
kBsSAl6pnP/UCrZPh6bWVrKbRiajdMTZ/B6Y9VnTZ9OZvE6c5S/g5bAG1NPFprUf
HGlMEtgWuOJXMXkvmutY/kW9ooQ9qVCX8/cW+MgLguCH14OuWheSUFzcusufL7Aa
qS9oyQQYfAj0Qss/AU3q7FGZh0XrPepjHWaG7gEg1rPBuCEpPSh5nVcsThcv6IDg
mTaAkbff4SX8f/g6U5AIqn5eAcjO2M6DgYbcTtFrV/zkQN3RAo7u3ZvLn5JAUDBb
hIhIsUoeVdnGqjlzxqI+TgH9MYdr9ASFr3b3P0ZaUxCrj/ePSLimu5YNXuNxHKYR
NnL+IfR5jl9e5vs1P2qvXrO0Crm0kZ/udVMu95EVLFqRw4zH55Ht0W9OlJQBU9he
pr7dcr5ALHPuOTTIm+XBF1xtfyDCwrvYHsTrW3yO0LlQC1pa2imxGupm4zRpffJ9
Zif0anPu/DrD/dBEnnlYVsC0kPOc9+9a4fk9uFJc7jitO1ShGg9Tn/1iJpIu4YLo
Qgvmkdy1d1LTfn8JckNLcjKJplkCd7aF+S6Bs9KmqgrHsDwvxO4zfQ9dRyHCQf/J
elhl1YOAk06MQGDGVsBM+LnqKOyWfRWTmOFd3uttDHTLpd6q6KAdwKrzo9obGmRY
YUfv2zyfre/IoCHZzzXO4QPVdhKrs4Uj7kGOlhqO1ocU6/rbAYwy1ITeLLcPYv4N
MtCZ9KFdvfvefM+kBncO0SQt9pop1ahAetFDatUMnnMXFS/pC1NrvPVkiM/c/ok8
w4aIG0+V+fQss3f4ZPZkYO03OXTTwMEhFkXl28XRWRt1NMNJPifKkFXjeYaJdGYi
K5e0GLyR1v3aSN93zGe5a5Y3WMNVa5DqA9MFOVVw7y4k/Iu+YBO+MZX8pZWblhs+
DJTxLYeYa2bDlA7IFCSu8uNicAK7RhODVtF/Episdd+f2XnwuLpaWyWZPrQLmwNx
HI4FeLsEdyo/xtkfa4BngdqR4MHgHVdaESxSXinr6XG12X24gzhusxikbGODW05F
n7fQmn/4sXCqPn6lgGEnEj3jUYgiJy4acVKUhR3H5wWrtkzeiBXHIncvgDXSKLsv
pPpzFdWFl3R7NqP9khJKN+xAU44mpjCKtayb4uzXdCkbT/MNPPhr8haBMKt5f3li
HqRZcu+VlNrQvR5GcQIwJm7eojhN52kXSfQ+QcQI0KXJjdsirzBokI5Iq4l+Xpu4
Hk6dwa4NDU7XistDYASQYDq+Cq9Gho577rIuNBPYogViZ5+owrdVdlHC4lUVsF9K
3uc8ZFc5YfROn95MtgrhClLQLMEfP7l197rDxOAS0jnnNaFekBFamIQssSq1V2aW
VhhmxSmbS3EDMvZfclIuaW8Zg3tF89VbEW5wI9HcGX9a5U/k87WpoddBLi5mn2hC
N8XnBl0GxsfVLuwLGKWvMjukk6AwwcfsrJvllT0OZrix4P7bhRqtmStNZCflu4Nv
CtkJ71mmCNEkcu3+W5wV+8+XkEm8nHgIgG79eohlWHU7CouTPbRcovPmCk9rwTb6
fKqGp4zZP3MwGP4y2ayM4o8zcGWO2iqLkIxOaD4CSV+/NI/o/LjL9xAj4FMj0yUJ
LIh41qL5A5MHRg6PE/GMg6IZ2w1Y4Lm7uqXfGxg2m44R4KpXpufgMMLKi72fZ+FO
52hCPDcvhC3n+8k4Tr0WXvSzP9R8ahWencJDpnHJdXX5Ndl1lYnAMj09+PrvyrL5
eAfBJUdFq0du0hpXhtyP3vi+GlJH6UaJ8Pa+GhSOmqi7HVDKqBTI1+QkNQeKOZ1e
2OO9QtOhG2CypCph5o6W7Z1ZeZnB0OxaIA6oI5QlvqUmJgeZ6ukWyy28kldHYclX
R096DAId8W/O9mnxGBbhPT6hTmru8PgTnljWcHupNCYn80Hq42SoWyUeCxzfNoLZ
PqbimDrqD6Gwg/Uzih7ZW4+mqdFSymwFauKGMSR610jmHD8wX3G8O9zYWpXo2NEB
cbSeXhMkTsvBdYe062Z+yhCmmw9yGgxuf67t8qTDK/Y8F5F7+KNOC9nmJmg6FIIH
9KKgaVqcl7GfMaVZXTmR+uZPuSlccynX2r80puW+geuN4vf1UNH89dizVXVuEv6Z
V2QbPy1JCh039+SKYwBSTnQi6RKxst6vQJp/zNoAb5mj82W/JHjbBkE8rH4HZe0i
lv0yrOA09pNk9laxONspm/2WkoidsDC75d/Ps9+UsdBt00lclowSkW/JGaZz7KbW
OdteGNba+gtUJHS2pyuciU0woUuAOGlXBp7eSq13ye4SSwefviwn/p6RqRsPHZTZ
a9NTwg1gcSa/aB4PrbKocGHBBhAP90TYIjDLxHQAEWab0Ak+gczijlRw09Hq3zfU
dDuKPFIZV9mX0O9CrSrlLl3hrOVch4pTVOGhXJiOlWZd7n2D8W8EtqvrDHVwLQPC
HCK/HuCrcfmpcQUlgopGrrKj9z3gSoB/0AarwmJLgKTr5b+fGrbGC4jqOKZ52bTK
7bDgEWpVYwJ0mN8n9oOvFB12Jl+ZUviDKQQyq37W8yFjULNCjJdtAId2/6ZEpDUl
6BnBs0KdqI5QkweR7wCwiTJeJ3kz8Z561R2B3YD8JrLNdEltPMEHJ/eOL968/xC6
3zPkyrxckRMalt1A8NL5Ck1gP1SOAsNZV3/dRyb8lKUOUZTuFZ+sa4jA9mY6tzfj
6DCtJ7SB4ewwxlfpyhXn/Jdvm9xbNggntY7iSO9NsAHlrNUat0ppakhb7QmFSbP6
+1YYOlYWwskIs4tBkFMuOhqOVb+p8fMVBO98+ngZAHX4HTeeG0J4fyxs8UZBU/Ii
Jqg07fUTPTIDMVW1/lTNnW8fmx/yNwTltPw98wYaI567z2EMOjhQyuSu6AvUWLnF
XTW7bo21D4EZo4pQGptVtT/g7gFIj5ez0K2MoA+eIGogGgGvUXIkpNVR21GNDrgp
oJaBPrAHvsLEoFnGePDrxl1mlpxxQhPu6pI8/ltwJcszBwHTk4kZ/G19adumzzm4
zMpZzoIgjRESxN7EnqL3yPfhRRoynySQtxfGr5YK+7BI3uu299mFtQoMh19Cf3Qh
m4FO3ddiIEq0hdZg5WbxwJPr4Ii8LGwGRlxu4udnwTAmowqVATYuVqVx9IhmvDh4
VkwWZfP3NRtY6CxqtRqQEKrO/g1dTxxpjJcotBmDfP/nGK58o2gUthQFbUTk4Ngi
Ao8YJlurHt19KD1PEl5BLg1XC9/UqCSEuOuAHxbS05+wc0ACmgGHREocIKKpUJmC
2gUHT5w9HsWcVy7zG36wIQwL4X3VNBCMYfT9FizO55b7byCv7FdKflhzz5i4UvG3
oZx/BUDZfE67FO6ySJVxTu66FXJDaZ68W030jdE3DeVoGVqqiJdjAzekLzWZWW3i
ES1u0AFIaeKNApZyUCSgvnj7oRBmJxwmcVFZWJLYh8vnuhcs8VjMo5vQkgYE3Ypo
IIYNTF9Y/gFCl2Gsv64CR7TWreMZkdhT7GeyE1bA2smGZjdwdyFqItAHzHNxuYVT
WNs38uOvEbiSBFVGvb2BzKPxjfOMkIb5G7TuUSI1HCxbOEPG2RGgWmgssvG7z0EF
YATPvJ+5ZQVIZH0zVJam0HXTapptEqXy/8NlbJ/jq+9TNFbgZViXFnUUK3LoDD1w
f1d0DQyIT0SVAYWOAvPj6T3bcAljOmQ4+gA0xQjSztjaqj68aBBhfbZgfh5Wl0YR
qrG7wWeOTD6E2aIYh3N0aXYArdYbqq950YxG3I2qxYrexhpcoPSPi29iY8cz94U5
xMMw7lVx37IbKPq6Upm3h3VAL55geO8lz87WDikA4onO4i9FMtkKpcMBW0duokWc
0oehWc97bC0ibp6h7dZRVWnjl9sWJMaPLJQWmugxkQ8aN+cb7me9p7H88wNLqTAk
lbG/5FgKNGReg4seIUoCd0USTEDYztTXXZDfhERX+/Lms4LEhNBVRXAC7aCi/qT5
3n2Q0hxVodD+LiETqpACVHd16ZDnGJHkmDRF7DFZXIHb/5C5fVI6LeI+72aLKO2P
z11xu+4KHgjxKWCxiKpcO8qiM2iMEW7TS3m7QFZWxt4JWr00MGFNcPVdiN4NfaDc
iHsk+FitVmeZJLm7cWeUYIspiTfMa1nJxYSwDTOI2LP8EArxt/gIi9sxkpok27Xp
lETX0TzNb82nNaZFr3Jr/RYLX4511MOJDSuMmHM8PxDrQa389KB5UsghlO2dj4CD
C9dM5I72bXdR9jRXBAXrAqr9yN6zIFSMnxu4X531QBWyqzO8xPnzKbu425NcBiV9
xTmdqv3oo9wmiPH6QbSddSb0rsmXhGKExg3pKWonalbBXkkcTM4S4w2qTnsWGPhe
H+84mYgYGySbJY7KxQhssz3htnC+TphQq0bzDUKbvDp4nIt+1FKoNHGy83+khJXF
Z8YY3IxREGmIFx46urnYSM4M2EK3r4RXdwMt08r7cCIsplf2z7JDyqCYBe6eurTc
vQtf71/uZbxZfQNiP6LOpJm74v5Hj7M9thu6HocNxttZrwfPGbxw+/bCRLNkkokr
dqYIozpIItskVGnFIjSp/+fPnmTucd007ERgUtIcQHfT26dsNzD0V4Vg/5ihKY0d
0tF5Zzn97hpmXITDr8QD+OX0nIPJcJJ5dnCx3arC1MSXkTM21b4lpcwWoDSWIx+E
0TBzrDJJDEgnvuvex24lz7f7Jl1wmw9g12rFdKQe36xrJyhauvgh/kI2os4mpmaT
/2WVkIo0/b51PgQuYQwcb92xRVoIUV6x1HL9O6JECwXjs51nIXP2JbCsmW1dliV1
3qQ69duofe/HeveuXiSYuBU6Q242BIP0C7d6pvHvlpDDRZ0WVULpd3iVjrYJN9+E
2CYNoaO6bJfmo7F0Ny1E4j+bOVKmjFGynZW7I8tMzUGbusY7ILMowfCox61Qp7pz
465Vn1GKxF5fVmrO/1POiV+SADs0pXl90JXbJBeqXwL78Maj3IU22k4GqyePu0Mz
14K++GZM0ecvAzkWu5lD0evi2yv3uFX+3a6QzGkOHsQwrIC0w1kygbqRGMe/0x1L
pZfmvCX1A8l+2nRwHwEZ85KpFK2WI2GdI4RirQ4WdTkohkjFgRNMyL29u/iRhpAo
2DsUd3zL1XyG4tcUTRHNMLBnzWV1cZYuB/YB4aCFUgu89leWcSbftytg5Ayy9ysd
42hyYmPg7wtQebDlwU2eelVJfF1/NJAR+feBj6s1u398gSWdlv4qzkyoz0c6aOhZ
v1bH1V2PCzgZlM4TIP+sw975W+NfrxgqDVyurCCacMtBjYnIy1GzmBgx37ZozdvM
2QnYpZwpPLjsIxATC+Nqd1mcuZTZ0WlRHRGRFfPxxgiK22fmAAWIJgojfplLPL7E
K88NO7Vi1BAK+fxPRnA5jyLxDwRtKSdAxa8NUCJULSoPOZvsZ6TBo0MLURFFsZ+0
tZRIc9j+sUOulzucSNE8C1sDFocmrMjQ1QbjFFHJyFYxOCw9c8ur2tOkbB56BHZU
Cvo9BIo8uROIDsFccyL5hTqPWgYSdTjFdZcrm1G5BMvG8xZ8yol5s1qut9KPkhM4
5iasVtHOnOW+KapBsIAxbSQeLLP4AuUl4KaeUkA2uGDtnmdMVaMlWkbHL6nyq17c
9DizmeLCPX0LmBLNZiz1KEKF7zAZqX+XNFpUKO+CuVWD58POSs6TfP7rwUqpQKoU
pC3l3qXYsU01+as+0rupL3tIT7CTD4kFaCV2LoBdaJWznd7FqzRsYXHRsL5v+se6
Ar8d3z/7oNXCxXbCNHHWunJQ7Qiz6X0x+y4bY6WfSLaUPxkUuoK39PRPCzUEw8jm
p8i1hlomHaMaG8zFXCIgmZ7TxjUwB09icOEGYFmpe302P2HUPw/q4/3kX4yMGZu4
lpsoohyIVrRwBuz4sPHhcU9r4mmcgDfFodZxb7qVbnRTh1s+zSL+YE5Er/ZtmFKv
5HPl58OPBoWIof/jrhhdXDBdcTa5AJKBLem5hKdfM/gL012i/O1CiQja4yEj3XcF
Mty8GH7XTE50d50WojnTqVaD16D2qmSpY/g+NM8W30Nd+2ed1D5qr1THCkSeUUVZ
34+hmG4grG8QbS6uqtTTlJzD9uwlVCkKmzOPLlzHvf7tbFssvQNQkF37x0+DTyLT
gaBQyzOyFXn9RYLxo1K2b7JCuLfp/gA/6SSwcbBplb17OajCr6/ZQjjccPD+Lc13
2hfF0jIF6t3cjKNGvp+mZ348Qx+DvYymhmzmhQuY/UUrEgGGPWWPno1HTkz1wYIP
uU36RhUf9Jjn/oSSWo+TXk2c2CuJ+l4VUbP8gnLWk3spJ4S3OGCykTjH7hsZ3uFp
XZLQAXPDMWhwdktnlR3lbG2XoDJzQ3yXHx6wFe1k0GabcXcv02oFYrNUXGcif56z
WwKbxhhpAZfjUB9xpGvc9PBDYWrPbtg/pJRAOslcU6Rg3NbBsNMEZ3CS4hERt6Xd
wgDvIhdmyymXKWmMJziXlyIOR8sMq3HN6rDYnpHXCrQRQ/iMFmhyiPZJKuAqgJ9b
ZwM7obl6g37tJyIQEe4RWXQiWgWx/vytAapgjm+mJj6dBGpFefLFwir1RF03665e
hEYBRZoVIllqlGrCQYacxAXxowSNMEnJ8qjk8ZNFik/nPWT4gXZL6oDW8p0K0JTU
eFBKzjkhdHpgZRh/262xJ5ANZmlVSVR7Wy51f1NLERxbk2wbfjQzWNoNFG5v9LQH
DgVQL2OQpV8iQvCXnY3rPyXoofOYog/zG0ZPSU9mAS8OrtwPKM0CKmUnNCqOo64i
VMgLyWXYQ+Gi+w0TOwqaSgxLgZMR4UBGiXdHHIg3f1JC6o4x+C9E5aF2gW8wNtXN
ndnAbOXRadhIL85PSjJ+fiGsqRKhjdsuTQtNp90tMNZyt7/41MZKLBmmkTf618wD
nD05tVHOqOhHwQ91f4vHlfXbTbvcMIJoa9WsjwmuYqZcldGazjDCGSF/WOLiaPa9
tSwQtgm1jb/ekRt+/B2i5P4o/FXGEed+DTC+qWXAouqTJjCVnqUix3R+FFuRRAjy
hBCBkKVghLz2wHe0fLq20EWVsscHH0gszhk7EneyZuY3+ArfBrLbqoQqP0WSs29m
HfibNGeowiJLxXU3n2qIIFOGH1xURizkA60rNCZMZR9Q39D44S2yIAXrXcqBWGfN
78t5WmcHa3cjaGWV0qWVW33rtfKF3sr5llItctHvoB4FMa0g1a1HdnjR6/u9ZDos
fBxPe2uq0z6XTxUuQKRCrO2G9cagrhHcXA+tPMf9nB7YtIY9BMHNZST0XbOPZ2+B
wnOZe4346A+lA7s6vYVPLSA9u1UfP7/gidh81CU58lPkR3mL0MwNRwM85Jb1Pzg8
KM3Hs+ogCiJPOFh8lPLWWo6y9z4GQpr1i4IxaSM+h338ITFo8D7nk0zoy05tx2qF
YvRqyid+Q1yX3TmYYuKzp408jgD5Sp/HpxgE6wxQ9a4vBUSZ211c1Qz3CwGNGBdx
wkphSuBk7xSvkxuS7iv2ZwY1uHmAA0TsWUtLR24oQy9RPHFuKdLFqA09CzJr7Zkm
X31tP/wxsbs+gb7Xvtq52/2o4186qBAkMIVk0KxNH6eYMK7zzkM9OcecYnEA1u+0
SztBqnyibzaeyOe30LFgcFbi+FqAktPhTXPRztVLwysLOLkuKOvN6pcJwHO7bk76
vIOayXrTFjfpQz9aDkcdVsSoqznOpfFmEiOAokXofbJ2Cx+9q8xR6TH5l/HwTa0V
HKTeof9/oViA8XogU/WFWGA4VnhTFYtygoXhwLYZWr9+o8Q+swGg2V1RlxqcXrPj
agrP6SdLCTMagLvyiuDJeytWCqapphc/B9URXuyhqNbYPXYR4jDfc6/1GBy7AErz
1WdMarDbp0ctt1r2EewiBDw3ULHKGWOUTQJwle+KQC3E744GMtx66bnRg3+UJqLu
xRg/6Hhw16l8gv0eA2MtuoLbcO94mJsZlHj6SZ/AEmTZBsVMPzUMvv3SmiQFpEOe
GpsjF5H2G57lqixtGfGHsgxlfEekCwEWGc/PZTFN4yUbIslCuTvbbceqT9xg1Z0O
0e6Ji/oseJmzBS1vBCd3u3pXKMnZOmGQzBfT9m5S5aC5Lgalk9S27ia2B+uI8FKR
6iHGoBRgB5tmBSg0RlN2Ok3x/ekVCEiBHaAwffmF6qCP2B9rzoD17ci30r27UMtl
sDQtqCSG/0mRFqAKmDSMAfPZxjeBTe1fd0/Hk8yHR+uEycyVwfGUj9Hq/yna1ekQ
Kry8zZCFSDlDyFsLmERoXXZyQsxIbd88YZNVpb1rSvsasYigKvMZ5Zti3JZK5B8Q
2Q4WwkAvNi3OAasr4WGBrN+qw/wNQp0vwfeNxqup7mKWLFDG1SPgSmgqrIVpXCji
kzn183eRZdiijUcNyvTwBxf/SQaMtFYAXAIT2p9515ZNkx0oi4JbM6S6t2vZ/GxK
ZvurKTWrKsyOi88sKXR100e33PZoTKlAB4LZ3nu8b19oKBfrsR/UZsDV1wcV/LNv
aljmmINanoZoxsJ4HPGQW0q2yMN+WE0Qjk1keUCI4AxUPu24C0+iAbDOoPZmONhh
QzaJpEQdEscAuwu2OnyRQBxNd4EYKLAoPUhQ2r6KuZeVMIA5jHEKg8cLpA1DXTsn
fOJouzTK4ZphQlz2if4MANV2y+Ydr+foJpq/CNcVcwDR1R6OjHA8AZbxAybAzWgA
NVDMtOuloDwcRrYvKeZ09+j5MBAcJMMJzeiXjNw81gMGnBZsaKm0aTKsKts/EzrG
Z29cLSOZwpvbbYiky7k4oroD5dzTn4T/gqeNm446o6HoCPHkZQaBk7SQ1MPcXujc
8uaiWov7IYTUeY6aQAWNl6xwOg4607Gb5In8OwzqtZPXS6U/rSpqlqCsin/y8kP1
ml+6sJJ7osYTgrns8j3Yr0FxAoXDfj0LNOQ7Yr+k/roA5oIkii0Knul+rdnhSI94
Hvzo0+FPPgY2MhtixBZLSY9jE277sOh4S1kgLX9ZLGzTane95ZnMpuwstVHiVbHr
pp7A+v3e3HdRNCI6Xb5jMEJrxzZhw94ORAbYFr76HlvNQNHjzJv6gdTdQFtz9FRm
o9mPhQNB1TSTOmVpypwfEtBl909JZ+9VTNxcOQJ72xzL+NiE75XkojMjYSJ4gJIP
l7m/Ftx5S01wno5KeSECLEhZ7l1K3yLNwxbL+xL3x1W/96QBOOkQCeLRB5pgOLgm
AimLGhzqKrpZ/HoaoQx1Yztti+dXkwcSd9WTqrg89KvMneXhbgaAKsS3ZVYi+obw
+Bjfio/ZFfzEE6zc9cs3LszF3N9LuMbaBbhKUGEWHAAVxV61DV7YxnZwvgWpofpu
GQ3USQOMs+M5RwY6UkQY43gljFNDno+aOkjjYLfe5CWuMX5OFwyL5T8BXRC3L2fX
r14H2gHBynHAzAg7D+iQtx25mxyh9y/j3jH7ZJhE7QwP4yKF2Pe/f0y4cm5A6H+K
v4RqabvUFPPi4vfVqRrf0M91LX+0QiJyxqw8Y4nG3kHqr4G0nRT7PmMdKI2FqVXz
nDaJSqUPDyDAR9mUqxlg3UsyzcXA02a3QWVjIYUTr5gNWSiyamdycZQgO5mrviRW
g85EYqf8Fb6XCQn7oRGL/w13yLG0yNTivc5X24CFEyycxWT2U3zw7zxyLv4Y5ETV
QusRRciioPOUk0a0TSfpCPReI4vvdzcyB5oaex/mOP5WT8TqWDQloF/1FsxaPAQk
u+dujOD7zn4uRVU5jpUV6roXX54Wa7EvfPF1ws1FV/tQN1QQyCXOrJEE7UyW7DwF
lMEEa/XfjK+XPFbQtJKhZEjiVPPelFTLnUFymj5rvtW/sYCqWpPhEbd6BbGGtVJs
dq1QHX7+AGB/fTlrsd4QTrs6J7j3aSNF1CEMmMQc5amGm9Yt/gqON7LqloIwXayg
MzkasKhKK5i+mwUCGch3TjzTNShP6Ch72XvVIsECOVLcceUgfLUC7hHPMg+A8kjZ
ciCqRL69i77PCttwDTPErZvCE/eyo83bI8IuD+26nS2WKwoAV9MT9bRU4pjK+TmD
OPgGr2cMGUTOxo2XWkaduj5Zo21Dex3gaPnSTmO4OQJArf7qQLnl09p936PKKcSN
8VJ0Bs7BrnBULeVCzow227oaZLvBiRfwFjjML7Ye3wSup+Vtcw9OukjUIP1vEo4s
GGK4ZOG0owwfR9+78Vbl62VTPI5VljwblUyj94XSKM6nQA9FNMLu9NBt6CCyvFwD
cb7Ck/pYRLZ5iVI5o9AQPkeJjMR0dbi53jPQ1LgmkqlHjmx4pO8h99WIEqT00aXT
KcvKHbpu1inahtnyW46IrX9Ne+XIaytKQUTeP1VW7UH62Ohomx/QWuOIUcdvjSh+
uvAF2kdaPVz4U5hbqC34muvg45bh89PwbaEXKfiTW9/L+DAdJPBlzWsR9mKc3F7y
OOIqLOzDuGHiEUQiaRo3arC7BGRJ0SRY5qZ3mpCUukrqcMR0Imxmk0QC0ov7STht
Uj/SgBPc5FJN3TZkK320FygePytt7NGAQNB9AW55UqITCg6HuUjlayrOmclmFOpB
sLV8leBCrDBiORSD1+CahCjiVSglouUF39Ixf9p28Bv2F/oBKsaU/qrWgKzg6Kxe
x8LppzAu87SZmp0yokzracq6o2luUkehmjBaulDpxXJKI9dZKk0bdI1saUrDbsuo
LOqRHdkwA78wBY36w77f6mwwDxRuTP89ydvi/2SRctu+7ceZW8xFbUR9eV7FAygH
KEel4ZM4u9ZfZpKxia/IOyKt+U8soTXACvBUUiecdVq9gvwDBamWJjB8eQwcreCW
efXp+xaXyh63doubjn4eggNLY3lIHomZYaWi+rEwzUQ30v7VcPWXmOSNToQt53Er
YtPdET0LhE+M3EZtRQ9AJ8bcUuVr8TPi3XpdREpJDGgHHCWQmCbu1CiNZEUOfZXW
6pOe/8uWNETVS2R/FF4UUBns5mfYyT4LZnyD2JE2QQKJTMBDtgmUbSV9yGDAE3lZ
7pCWl0d6xhQD8JxEwCQG7NJY8NMIy2e7F+344d3rWBsmxFRwIMSsE5FnYHzU8qht
awQ7D3UFN8pC01ih1H5XyrCM9aQngnki6eETUzHOADmCFbzSIQQIF7ZQu4xzM6qc
3KwVZx6oAQk7SEED/wnEO8JbpfBwdcr/gtrKt5zdArr5xBxDIDUFuLhsXuCyHQ/o
eZegm1Vywo5MsW0WNRmalnQNDkzQpNIocAchL78CcaOb6o8o2ocv+1/Rd/nwBDwY
WPNW/Y2F7RqF+Prw4XzGvPWah2Cp1bjLWGZMcsxYUiwSbAK3NN2lnlg1L/nVQWah
LUpqIRAkPWyJMegW2OnGamNKhpSNqe0u7knhLrvwkCH9B3+ciL6tLpUta6FjSQ88
Rd0o4nY528cFp7v3tQ3u2kDKQhG/Gro9Fl0qyLUKGunK3TMqFKvUKzjqT7fiaHV1
VrsXjLm6qoS3oH1XPFrNCzRIv1cjvbiZreReKOLOM1rVHAiOcwrmIjTytahIZILm
cQsyIu5daBbZQ1yfwnCdhONQuRpkZ+OH4ZEjJnisuxMqMGbMUu4KIxvBunkRQ5l5
cTFWj/z4GFmU3tRMXC9Tb1GprPf9Sm920bdHHt89t0buzQQWa1M/fPrqbLchodtC
ik7V+ARP7QJnnu6+jgsGQWprHZqf8KSCGHUKvTHGQ7PeLvWPYCPwb9Uj9C+rWXwn
QjcK46FFXFp+EIVxZfozRS+MGfb/Gj45XR1PWgla9qw0mVvKbGYNr63DJxAOscHw
nP8zTbis+yQ+SCcgrl4TEYICX7PkwHYytdJDLwSuhn3GeD8chlmhODXf6kDWXwFp
rwmUlLdj7FGvUQ6OsQ6a4cKS3RrotE/7i/jj0dCHrIYEEgURYN6Za1HI0cmo72S7
D/pBfpgIsO9nzaxm0rStg4n3BQLu6apUc+uc1ci5+J4ouAFuDwoFCgvzHmW1aOT3
39pb7oCOkYOEo6DAJB0frMxOQKlcywFxp8tXJG83UUyf12yzsEDovCsS7zNypgc1
rMy344zAFkZ3GD/QGbOCG+SebsKjM9bbYTo3IwocX/uH1gYZidJyIReeKtDjzjyQ
0MndnARVf+urBLejVZTj7r5MxZrtzmxJzUHs80DnVu7PH0qSb786K4SQQjboIwj2
48A2izp9ElZ2u92XHheK6XkeIFYIPjjXGkgA4bP88/+pzfRUCB/B0/FVv1VCyNP2
YHasxFdRmaXBpyEa3uuXSekKr9+N52CJDIPq3ApH39iyBpyn0iY8qgm2h4HPo6mO
nX4A02urhqUdPFgI+20ITVFDi+D/RsX0uawEoW2woOorPNWI1QdvRZLrcE9NWREG
j04REfTAzUqiu6RosKPcqsFkxJ75J93yXfHNeONYUux+n31Kg6qYJcKAcIlmgeeb
sJefdoCU02E+8K1rZBazhcqM/ZTFchYPILqjZnuT+/0AuZKMYaqwS7J3zNVDMTmO
E9XEGRO6DjrIP9Zh3s7LKxtHedsBmr+cCsnJF+FfJfrplrv5ETL1QYfQ1NZ7dfUz
ILRoVbBbsoobqnO+4zG1/zB52oDqm53VQhkdBCrpSFyU7sX4C+Y/KfCbzilRLAZi
yHXeeEqxOSjNpKzu+XHZlOcuDoSB6yG6BeDA7p8snXN0iqkDBJkU1T1zboj+SuQr
+v6p0mRTLAUsq0D4JIHNPHizZVECwfdWvHlAwchrlxVlf3owEA8jikj5hQk0Tlwy
FSGyFPvW7+g9OZs4HnlvSlXBAsJ41wLqVpVHotJ2rJtDoEtjEhx0W4bBESLAMbOR
jxqVytumZsG1ut8xqRQN8768xry2iB4vTs4RtbUFl5EnNXznxIxC6cahS/36TAJW
d3TAq1cc2e6NWWDITmQE5sduA4GK9JtR2RFEaNfbnptBO4Q0QuYd4UXyTajMqg4f
d9SMiILMlJVahgYLcjFDWnATbR6YjSS7yvTDdk5AgXNgs4s7vlppR0gkoFnBUp6h
epIqAekiS2k8kFu7lWQjFdy23U0xiIwKcqSNa+BKO/FXwYdRvmMXE6CHgdYXIH+f
bmprKMDJdwopfO5mDq+HJA82cpaCL+zeEhzsEqF/UQHyaahEtU3dyQwl/Pwpfipg
9OaKtKQ9r0Vt1jbDYCNgnde1aekaOwGm2zBh4CkkEfozzCBn6lNDkt7n5KVpm7by
QS4dw0w/QYAFaFQdR6uKXUdJO+TXgBZsG3R/BcGYTxjISxRALi9aa09gym8/d4Kk
DBHo5UiWyi+1h8yJPsmlxxUBZ55oiTodRzprcl2yPSYpK6jlW+vHjVHGpaRXk4pu
/RO9C1eoIXNm2y5u81S7kNKLGzJGS3QW7taM3zMiMeLjeJJVo6K+hm5dSoa6Lmay
r7N1ZzS2pTs0+V60fo3dtGgegdJC6X3xnAe9IQ5n1SFYXwCIPwnKOioYWYN7SxHS
VyqIJ868MMeU2/mRuKx3e8NChx9UJgwIQwyYoJQ/MVNCLb5bY5XYM5nBW31cXSq6
WXtUYHaCiSkVcPac18iuLsbsaK0FL3QgvvjMhVhF/nsfk74OLbYDG/V7zhir/PJl
sSY9DLCo5NPLLuK/EWvF4eoixSTTSJWeMQu2wEhHkYk1b6477F/SLdzLt8Mh5tnZ
SNEVUzOg9bn88usTR4cGIfwPO2zdp0e/hHJc6wMr6vyBiAsePkjHScefsj0hpGH6
MHE2CLcfthHnH3q6CalN6qMMhN2wmFcWybMNXVqDonL4QWXPtL8cPXME3DUuYONu
f1g6BhPG7O0QoYLAZL8uq9Ks0HIcIfScqDaGU3EbYUJSf45aHo2m1g0j+T3axasv
ycZTo9jM6B3X/EsqCUrfcHz80b+HBTifwwNP1n8CPAs4I5O7G5XT+W/2ah1u8q6f
Cn84SsJ0//mVmJMszOrAU6RTIdNFedMFL2SCR1M0pcciw0cPTp0XBTKH38xbiXkg
Y+ZUAhP4/a9h2ZT6JbWtTxLIoz3ikBQrzF24NsZTe3/L0K8AuwoopHQgOnEj2yWU
1pNIpY1EXicWYtmcus39CwWwb3x3L99WPrbndXK5g1y6QOxwPLJq/ChvjNnzZPWA
Ftf/eWfc2ika1se9QdBIN7gCMk7WkHnC6s2BhheovFtF+dPxkqEIVH8mfucWog6x
CnSaz8BmJvQGr0tVlvBMdZmg/uPZAzc//UcApS8ikaF38YyrY/y10uMhSLRQSr0/
5byvvuIxgffULiI9I0NMAeVaxY2Iw4p92+HdwFMdhJrcyXnjiQ7aIiLF77lPRN+F
4PUftllbvvj/1FO1lFcErsaQuWqPkexKu6OcfRxmTHfBliZnd3Qvx9NPqQ+6fgUK
8MrX1NRE39jbVNGBhDHuRl9K4ToNpqm05HVK2M3EhEs0gyd6duCkc4WsJMWLBG71
mKRUDSWIBPi/04WspWeNYnqlCsEAHJhviPyGI0UI7eaeSUUeAZ2lm4u2EJx0ewRo
HMDuxGydtdjf7CgV4e3emx5+9XTaWxNbfFZ7ipsmISg+B1wHE5+PXt3qXOd66jiO
WPSpDG5EEhpaZTR/AEe3xIRJT39qL3YwZy+wj2lJfK7qhuY4yymFx07hlW1WrVtD
ZsoJZ8syE7YtEIezgWmLP4vcyjlpQGoRkjy+IYVFi7Up/CcBeL0L//oqsdgJT60S
VUhgTPLeStgbYTtBpKiQXtKMNIoNV9EEGlPI0D9BjlOySnSAOLiDqH5gJbSE7G0L
mc9B2LdTRgdyER5xC0iugmzBdcVTiY2AAQgdNGwHn8PTHKFVChmLqismsXFDI5Ko
QHsZ98jiNtV6NGFKnHWIH8EgUGFgdD7/sQpgXSAdyDC+b+jhaoUKHYCkUbZbS/f3
Jl4NHWxo4VHdGgU98uaK//Ohpi8MSGvly/ByV23md8UAPrIcZti5aeYZp5T43m1y
MnE+U4kYUngU7FJY92ZITsAFPwfAdJqRJ2xCc4afaOEGl2LLwWYD3H3Rbiqlz2du
gt/+ZbZIfWvvQ99MpFaOM2ckz8dm2Se1pFK5+V82S5zuvwncPocB+uzZnLI6una6
N0Yrp9WcxQl5heN6ts326OrEUyY0bPssMa/pUbT/UBhBTC4MgLMcqrbB8F/13zZ1
nEKmb2L4UcJZm6MDB2ut1e9usGNDQkHv2Fci5JtDGFjb/r84OISegWcH/L8drlCz
tLB9GYuNaUKayYLyrUdIM5VZ5nmn9Ki6V0LDBSlD+e7JQgdS3jyIAxTi2ode+OCe
fodaEou4lSpU9XRdX7q+huYtJ+ciuTES5IeDHJMNBJEklvhkp/JE7EdEBqd9DLny
QkW9SGXaEnX/7DIs9y2xRpPjpbrG4J9jxLaL04+sIPxz+UvhmUexO0y4DcHFBJgR
aOZvq14JFcmSHWCGh0sSoPO/igof13wS9LLjEcfF+PS9drvhy5zMDGOCXBG0cUgT
Z2eYr8zs45f8P/OhAwmHKdKB7nxxMbRaGBP4JoL6ZDf+40HUm9V51HyY50G2WMiP
UyFq71wmlSnHO5U08iFHT8cex3yQhAi8IsOa339Lzt8sqAO0uGNBgjQzyOTzjmQ0
+/lZeamJPAHoxWD3jcLQ6udj2j0w76Pg2VvMzzJa+5pP7ZcliNo3fcebq/Yu72LG
vaVTNteX4jTqgE76QwEPTsV3qdlAq+z1+iDQFjuvUkDB8T4yLCYshmVmvB+oTQS7
2ZDJQ3S3wRXmRDJMBg2pvT/wYIIs0RPOh82Vi5/EcJM3FaHYsNAL49cx+JutTkgH
QfkzeHcan5V0DyP31pau0VQ/2znEV+SIhYRZY26U05flXS+a8uWI7O6r6795DjJi
s4tNLHnRfsb+qZBTaKMdtWKI6kqwC12qS4d+eXF6pDFcYthvS5shd7GIMJMccP7x
WpiHCIpqG0L0yEo0kmiXnwdIwxf9aR7AxOWwD9Pl9huctgdLqgPpe+GJ5TvLxNEW
PPViMgvwgyrkUZO+EQ81zJ5SX9yc1eByeWUXAy0n3PPSzNpt35POvaLStjmRkHUM
Wp3RfR93DLofTjgMwYpsp9BbUuyiN1hpi0q7XOnYLWf+vyfQrlca974bsyBWaolC
Jpdqspw95lsBxCWXVg3HxgvRJuvO5ROzB9xFrE6f1E7N01IbZ2OK+Nd0Go5PYwok
e6qdc4Hxfv+ua4vMztp0K9mnQNw1JoNRtpO3B+4bFvF5DBD8aoOBQDKPAJ40N4sB
Ba0Nzyi72BXUsbDTwKH+Z/IC+L+wsXGp2U/y/2IgwdM6POJcTbbjUjTqd+h6iZcI
tCD65SC/yhlXQTh1WRg5eLGQB9lACxtba0EHFyFXFxZORlVaGo6IqWvN+MEzKI6/
UrIcHyX5bbYgHjgPdwW8t5enZ18oObfK3ValmgtBx4xupyhTT9sm5L0MznHAJJK7
c4HeuFAgr6o14+0pXB/fbhvmBE1kC3BcFqLZF4RxW3NABrhpNL4CCmxhQE2Ll3bq
109WIx8hWFa7ez8+0HfL188OrTIAvU/NCi67j/ZeunBOKkgVTkZWOpYZTB2gsiFS
gl3YaGjn3DNnQ8txJivnXikJ5V8QmVjWtCSJ0euLeQizLvf74uaKv9vrj+oeIoyZ
QdDa6AFxYl5wDfwPTUu0BtD7j10K7fs7QY0/JjqmTNkVxa3prTh9nncfokkjeKmq
v5wlmbVPAuORLdm2HvDHh3P3+6HCzYFfXmDwRB8/A2QoyEG1W1D/8yk2SeWARE++
RGBU0R54EJp9h87w9kC/bt79/UKSeGn/oGEw+aP3VI+cXiAK9uzPtgTUVTQdVD/b
MMfj6Jncps82iYkvvMjkX6I8BJZyFJkB7e6i56gByPR8ko5doweYj/MUiRpURv1S
kCugXg6Qv5Xya7l1XdF1aHZG0r8zE0/mrllU+IZYsFpnkPD1GFD/cIjvtZIRbtAy
KljH8RsW7p2IB65aN3pCSaL8A9BswntyJ2SmHbgyDh7xlWFkm+eWA4G/tyII9SPR
QEDfKCC6AW+rDs/hLJFEGVjX89AV9TwoAbrsKuYyqnOndzKa7sF/kvmBJd8gzBeF
WKyFoxvKxd02wsMr43XSH2L66iDaQpR/Kxx0jGFz2V1oSoj+mc8/19rtBXpEGDnb
aO9jXyqqSrNnl6P8bcEFoQbiJb9jV6zIXtxhMUAxFx2/RIT5Y12uu1pNZRJo8Iy4
Svp57/w25cEvLzwvUxMOp//96+9NL2NTINVBUQILE2C/XzH+Csd+aiCZaZdMtWl1
tlThU3wxLaJ2E+nf4TXxH2p8l7gO9VyWCt+6sNHOqpoPStlyd87PVZf9gxGUmw61
VNfSkrtRsNWA7sNrOl96nzQBXjviYfxE+l1bibtfHffU+8xyc/LURWGkltA3fpxE
3IKwyFQvGvkvlW34GHYl1c5IN2R2jRJ3AjvgRBUTIiB5/Dd+OsCnoL/n8v3wxddX
A2QgjRfr9Q8+UxnY5YgECipMufa8f8VYNBvPAGsGhGu4tFfsYDw6vc9taFwV27K7
QN/iqr/T/s8etBdhvAZ2+WyZ5PrSf3es6Wlc4hEXIZtjkusdmMBybxP/muSM+8Rq
5fZIy/YrLhzGu5qFwLKK5cIGpdd1gl0aUhY9x9jTDGb/kg7SKVnFLzj0oI8AwQEY
bSfAC3EMMzkGnbHx+kpvw+QKJ/qMGdgIhRK6qBdnTv4joSsyMHHbdIkuNDzjXYgD
jTRQvdeFZ8gvUXAGKJLF+Lh99YcFpr8NyyPhw/WFXpBb/jlBTChVguOqyEZPkjok
pvyLLb4PjVLDgMiZ0y4rJZFb3ihGTglw3dWgvN2YHfNPH/ybG3SuNJ6YFcLqqvGh
h7aXW1H6DpwQZdwO/RhiptCYbJYLv1oQVtZNq+lvQKmXE/4o9hD6eBpljZV9GmHi
+dratsqPnT8xkMwlCzdrCkONzTtyEPHNr7irh3fXSdFfsKglMCPSWPGYLCe7e2ZF
IJQquRSk8OKpCvENPJzOfGZQs+vKikdySeZ0kn/jW2qb7NJMin8zhy5Y6zfHSCYT
tWw0LAr7KKJcFbPbPS8znK5bVxbmRCd367rt7Uxg2X96zrAY4wuUu+TOR7qxXkKK
YPnMWjg5WbwvFTZGTUQmni78M0h6b6XEo2clGpgO+1Eow9fgoq0BedqstmZBs6JX
FSJMHSrsr39kiUKTkrM9Yq6hY0dXp66RiZP02nis/mcPbZh5pV3wCwWJlcsy2FiG
zcgV4cBZQlVo2si6mJhbTPA4Z/drF3rMmYMVoBdoa+Q5oI3NAly5kgPwvDpCrvnH
u3TuNR/rmVOFVhgaJ9SqRpfG6cH/dntZGIxDf839x8Gmqj2w68Hud6c2xaKej5Zj
z+TnlVVu1n/jY33cODzCNR3hPJVqBf+dRhKzb7MDK1BvPVsSZityMM7dI350ea5y
cz9g7sK4pGWtMYBvUtQO1LfnLwxiGmynLO4AnQdPk/cK1QEFYYhwAyL7Sr81ckNt
cjrty2+9yKd/l3riB5TDioVQ/9vrFOa9ay8KTiKX1fRbeHWB85rXOEdYEN0N3gWL
2ZkuVztaxpczKSLlOqR5rAhp4Paw6KMuXkWm/LNQyBfzma07gmJoFsBh/dBtPAei
hQruCBk2K63mLKjJz8rQ4GwX5YaAj5eg0cc/Lq4xasH3/5fCG63oCUsBgK2ge+Tc
foPC0Fq+skAve2j5TA6Yvmkw9qh2IXEgeIQp81+JxJpHXZUN+2ddn/I2LLHmJfoj
edmP3j5nYT1CkZrE2z1Mwdj7T8WF/o28GFPBNYR8h979ZZ023ZvSKXYs4hoKIaF2
u02R3XnBwp/IP3BlgihRGvJKMyspkMT5uqrRp5rTVRbSMqKRRJvPU9bmun4VXowx
ea1mN0dljo5lp92tfVllCpNJbDNuovNFuFPTk0zTLVMWgJrGNhO3G1eEqbc+/A4y
e8fAdVUf67g9/oMB1YaaCWZycOtW81RAOD0IHJDQwJfUvzZryoOzPdld9A+GuhzX
mzzgtFeYeWbOXq0nrzPTIZfYqKI7K6C0K2WQQJvMq7F1xZkvIjznE7pNMotpISzg
SBvJxRKHzUUbhOfq1xb/DFeSmA4A9RXcyClYgVzcl74FYJijNToFcc0Pr9YkhfHT
NL5zC010rs9a+cHfn41ZhoU+4OStb2QbfirkJkPNjMtUwKFe8CXXCCwpJr6EPRkj
AIDJOe2QDxafAydRwfjDlj3un+BDbGE0x6JM+FARcS0/zQwCyn3JTEG3XlpBu2OX
CQVl+l271o/RWHGCDGASzljbh5lCc5GEZMevILNMqOsylKcpOo1GB1LPADnRn3O8
6ngb14/zVxdfYfm+0oGYjotnEfZc7Vd0q6I+uADIcG/zzdg06GpOrOUJqZMs8b2e
PrMK/d1kP7YGJhy/FudmspJvU17GV93M3bQ99KoCyR/v2jZbJ9UzsMLmxt8Bd/xJ
NKCQXxHSh0vO00olSg+QJFORQABvVw0r7PQbybjlByjUBMSxjJh1sVl94bqQpjwP
2SL35Md/937/+LojxTgO1nsP0TCKlSClMJXrhc9MVCmWBmzeqiknAL6sTRgoOuUd
sC3pEfB6s9/R/XZNzNVDX9E4amPy19ej6ibIk67XsYm2FfeBPuLZLmpjhO2bxmAj
ZhtLdhDJco2VES7tvglJsSf5HbPCZCWA9YsiInULQNVhBzL/NaW22207aB/Qz5bC
Z6dnSiU7pjjHFr2VLjQSwVRNbAHoYTsS+LxKDLdqC/3YcakIhjgl3zaNfUspFJlP
L5Ic4dBk7MJx+gSMNJ1E0v9OOlB+7CfhlQznXzu1N03GiaB9fKilYSWD5o5W4rRq
mLvUz6Uk7iwMH6uS/TPqYlBhkLJb41o6OBfrhaB+BZYmLfqSlAquqdEp8lkJplVr
YnrBUgaTLMh7JE2qV1PRqTS/xeHPJF9PYXDQg1/E9WjLH4JtFv2PkZQ8PvNLaTJk
gaC7QBuhAbaVkzEb8ud8uWbbRfX8PSX7I0k81/TBt6QCJN2q9oIZHKgflPQpQpVt
3Hu7enjp30nW6Fk7EetV3hZEYwdpSKjuV8N1MazbUnom1WI2Qvm/abDD5245ifmc
8qV3cvkNILybj0NCf4Ahf7U4FuTsIuentJEjs6gn1DzJybTfmO0C0UzsfUiCsVK4
Rsgkanx44G3IhvdLzK1bdZJnjjFnNKAgA7dfAAj8RIKvDiVWQBUPtHmdZoSpR4k/
fZX+cZVugrbxbhH9oUvWa7e/HRUac+yxd7Jcm4ptqYCybqh1dsj/4eQbj4lmMHXf
lHxj+mg1PHzn1CNw+AW04vBaAuxRSfDXG9y0MB/PaYOpGfZBVH9zjFQUyYcFrJWI
C/iL9yCZ89l27HQP67Kqz9LzdSwNp25GKm17g1Cutpm9aIN5Tnftrev7ypa2UQ0V
3VPfCDQdr+pRcyuvhYLoAhLi8BdEkj+f/HMhDd9Ud1jjJP0HlbynxTIzSNGVuW6f
XEddJvG5FerjIX+mL7S9Ynjh2Nx3y0ND1cZY5o7CfQIQt3KgJ8I4hYOhchBMd3nc
Cb3DiPrNLsZa1IJY/LxwEGxQ8HPvIw55+qzkAclV0B5fh6+HGQ29uZw9EI60KtJL
Z6b27A0SFwijgJz5viM9Rh0pjjNw5K5WCnjBN3jqexm1uodX0a2PgcgTbSuMa/WL
ruHLbWzcNqw+opNIKfkC3IeMzkBhxtAaR8WVsFzPt0PSNbrBFN1QE9eEgMEw/CfN
6WsBzWIpxhu+ToyyFxTAwiXYexvaGEWsMZQFRWrG25MP5O6ggnxEIKdaBWjBZNw7
QGCUSRa5U9nzN4jEixR3y3b2s6H/ah39SMEVfJy68OMe09taLhmPTWrcwWeaBe9+
Tj9bID5wYwGyme/Zylmr4450uMb2PL+FRdkrZ16NTtdDGSvQe1ywGgWnOSWSB/iI
Z5nQ4KlL4IfOMr+XRHUpcQF0W6T0idU6y/i/q8I4FFjfrm4vVi2os1SEpOuEa/Qy
pvYHtnKAiaGtUCPyYQONkdLQsBtoM7Rtuw7w6Q1GGENxqbmhbIkCAEycEIIdxAaB
4TUVmJB6Kd/9qxeum70rPt7T3zQUSP0mcUHrLs4NG+PsIPaJx1TB16KMVk3HNMZe
VSbyCbL7FANVzngw2NCVSneFPtcAbY1l6PSNdQ9QNpyZNPZWTz0PZP2bSvYv4/J9
yEs4aASsF90VIDqbf0zAaEqvk/2oPsW6NSTCcBjweXi6v1/omOk1metrmr1thDCG
qxxLdbJ6hcsGff5xYXA02NnHPalTM4VNIaScwoRMfCsOxdAHW2k+XZRvgH6Zy39U
+2EewI/B7fjR63bkL/zN2ca0QMm6ASBYD6pmIBp9Egl4cPXHPzkRZB3g1NmQiUmG
E8WUYsgGce++JS4RyJnlQRavH06q9ihNhohS0KJq2pE8Jk45gqcbrF6KV45ZzVl1
BoCH1v4B73BjyZSZVSDZCmV5Q5A4Tw3TwuyeukBiI6RP5h88ft3YdQL6BVcjK43B
BHbKOE8AoZGthae/mWEHk9SUuqI4h/+dkuL0AXD7G8aOQ+2SGjDvtsYTLp9X8kwj
yNoeDL7yZ/PPSeCRsS/bpMZNuWM0Qh8jRuCsjW9MkOY1ldJYyhxQoMcsgqSf3mLS
44TNUSPKfA8YIiXooelhbylvG7FG/vwn0q+tGPaG2yYXGjKm+Wqb6MMHTFwGlxja
i5EnyGBOdFRmaMZYZVrYZTRJnN0CkVG5qP1QEVPP7fYb3A4p2zeYsHnH9+DMqEW0
f+pPA19DH9HDA6aG+93SsFo5lekRpnI1v2SP/dP7YMJIwDSeLtNWjHHls2YIotVC
6ndOqWJFUsP8h1b6HwJXHa1hUg/O3kqRe2T+BtIGGLw+SBDDRwNoK1NCPj9MrgFg
IKXvjUsUKwxDuyZae67vMf97J7tYGOVxHH1jc7IgqJks4tF30rVilAANfk9MRNK8
X32Pa5NWkvPfep+zZjDfSfHLU+vHrsOK4W0mYSJfaiEYs7kL8FZbGQMqVNGzZ0gS
Lp4FTE5iLZf0AuzB1bAavYCSKXy6EY1XIGj5B1q62JHJR6HAdaJeGeXKmjCFH4/V
4839diwFOsHPgNSFIopqhUo+gLpEjA3sxAmpaAnBxEYbOKMoke2SBtRssu34eqVq
PM3qvoJ95X8Bz3nllHA3sLr4TvcyEoiQ3sOxycNT1e7YtGcF1aPdjLe+AmhhOY9u
D33LCL3vSvUiJBJfpXPcg2lfRZnbBrfSwlSkjvB+oZfeq942+3gZM0EedsFsUD6n
PXxKK8CBX2Iv0eDf5ScSgLDv8nJdEHf4NgLbNGdet2h6UVofSlQLs84f1fD8Qn70
V/ubuAuU5HxY00N9ls1p3Pk36URiGnUgZpRXajnygAm6YnIVf/1LVjFTYGdLG1NX
ztVGl1ZqqwIX3+GaofxmLcrCH2gX6cVGNLgOzYyZx02WvNxt9gqdnuUmMfFAtIUY
hyvJhgFEkX8b6vsEg8cSAJxJAFPhc4rEwSHAHNzZKWrANFk1l+1PtrdLXs4KptFF
ZLEEqjKfieS4M/mBgeluDS2tT/LIPHeJMHimzxolze0n9VouIRT7GdjCQOXNZLQt
x7BZAfgvxF8IG5CbWGHSy7QXoLgadvDx20+MIDpu8Eym7BDt2vNi/hjCTJiDROhU
TaKkt4dUqlk4q120PJ2RZ51e+I3vNXvKOzHJWkSr3P3k4vLC9VnyBw7qdKLWH1vm
rbQaiJu6roz00gb1AkNoQxJIKgdghtkHBdmApyjV2JH73OR6ivEgvPAIRVCeka5d
WBuuLlqnJYVcEQMcODayllGoO1p6a3Yttla8htbfP6xO6S3BHrQKxNvQ3SvB3fiJ
4pLyU04VX1v06yPOC2Zbwyqn8+IJnUcI/lcPTtphR5VT5MxvmV9jEdYfU1oApkKA
E1taZW8YWD2Ndii08erF6dxiT/EyoW4+ulxk5BjkzohBS3XLUdyIFwzbt1eQksDE
7dcIMSNu2uHK/GRHKrkat6WbJu0rOcR+B1Azea8Sj57srdEtrmZdKHU3MPRjoFiJ
CdYIwv6gGZVq6u2bN6Tq0Vlp0744eY8U1ItOe+efz0BeqSXhnG12YpWVtIjAXpx6
ct0nyEDn8bdjz77e/Ylm+IzRJ21bHnTjGzXPalnXHQzsGnmf6VmOEjfR6HOX+FRA
6N91j7KmqBTyPt1o8BWWZxIL5mT45Zd4qpfOYiwZC7e68aQ32cqYmRULVyDPgDf2
jk9RzSJYlCzkUp4utuOwP4QaiLY2/1YqjuTJrBb7RP1LZ2X8DtMbXwLZ+iFYU4qy
tLp0LxF8HKVyrkxDhGjJesb+dQxaqccrtj69Q16YmR0YdavvqiYx8CXXgczOtA9s
KBhfpqZFoXvD0IfTs8T4yL6Mr0/nUjN+K5fCdHUi+gohu6ksYzCwf7b8jkrSjw2C
vuRkyKuxM646gBH1VZsPzUDamlEFvRhzfnyzRmSASxQZVHG8SZFcRk+TuhV7XsQb
stal54URecUfm8HG1X/PE7TCydsRgd6zbOuxf3tbeXH0m5whBCi1XvdJpFSjYR59
+3jd64388QmFZoXFWopzEUzm0htRQHizeuaTM/g4HTMm2v5MaefM4ekt1uhb5CJq
6YZdsnZeivetBsoUML2RSarbFxkYewm2uiH8xWuGwDKkqg7sDON9Own0Xqcn5u7r
td7KW3oZ6K/Fg1E7wkz+KUxUlzpF29Jb+rfua9tAbi0fN6G9dNa3k8+V5sZTBu7C
kk6QuTATKIu5wUKOiT9GWkD4B0KgFmo+tyTuHMHnah+8EjaB4/+QJykNSMM5S5Zi
FI0ikqNmGJl6+t99L9aZpzoTCiOqRE04pxYGGBQ4KV/OFInabevTOGIsUUqaXYjN
qV6fwktGr3YvyFD06p7QFXz+PSTuXXaMEqUuMO42sfqiy4wqW8OG2Xe6nDv3IgPQ
+55a5OVefBkGBl9FIfMag+kzJ+0tCDyZXu8hRwfwktjtjpyK/IsivOfdDS+2ikFf
UJy4O+HGZu6uGptKBJIwCjIVkLHnW8aqY0YR9UKOjbG9S4m+7WGpltfzh71bI/Rl
UPKV8nzQM16QW1QgrT95FTJvif1nBBjxCmxMmajDqyNHF2CZz6vgxdL7KUsWrcAJ
T+XWLqfGoSHeiVM5uy+Hte7UuuygwnXSpcK1YMQqxRVnNJ8QY/Kr8oiQTRqjKpST
JxbQ8NF1UAlFXJqAnuwJXvHZKJSPTFTq5ISzMUrxDKgVQErS57XjJQOFBJiiymhB
V4CtzXkEDTu8sGUlGlnwPAN/CZRTCIrtRPH2W2oKi+8p6yrFBDWUPu+Llb8K0rEg
4pEP80XnX+Zq6OO5CSCSzOqapnQgot4m4r2rUJTWcq73qaEavK2/7RpS9/mFyNVS
Xo9u2RcgwEpf0xxlaTCKbev2kFi4cwNlMq/xCuUvUQT5bi6r233SsNiwdTw5Z/2J
PV/LXj2kdCECmXieO9m1DpvXUGEMmQiSkv0w1KG9FrhvZq/KpQnfgeCUk0aLxZqU
pIj88bFbSp9aCh4oDSNlEVPqckG3BX/cDnIM0D9iR2QYMm45p9daNfcanPZ1Xpn7
bEAPm/ilHvWnRoBwo+UXxougc3Ae0qNinzZfp/VgtnR59yzayAodizmh8Wox+uiH
v4FQgBs1cV/l65lhdIzJxg99gIPkS3WcrrXT/EetFXvI+DdlZ6eKk+mJ35C60n0X
f0pzg0Wr6+Z93eyxUQzxK1OBresBIJMdpRJ6/nXXAAYFZwPOoaOl3e50CGlpxiV3
NU8GjkHsea3Qem+iWOCFD2BXJiJGHOJhsDeCZcoaJj02LN+lqKw/b6s3zonteDBf
BRPRQruoYaNFAY4z8X2lgBFPxRBaJ58/nTlWICc+tZAMsm+02l61oVHSg17IxaHe
kVYUNES99gi4YFaQkY0sSaZegyzh+vXHqHEd01Vy5PvIFmVFPj5hTTscmoUvFA4a
0CfQLDQtDIzy5V6Dx33fjaedILE5M6BP5mkCEBv0Earb+bgFwWhRyzpGcXD2MWHM
S5ZihHIcp1DJSQLlEc8S4c5rLUMElYR5MzDoR19OCAi9v/2tfIP/nAV0RvU3kjOn
2tOgXOR/6Yf8HzGs3f6QBy8E7F+ydVv9hjw/FXs3beUc5hhxuydVyHOtvFLrRhKZ
itjT/Q6fc78107Z23TMC9DMJkZGeBsMUOmKEE2+4GLPjj+v/cWkU+Zz3W86lrMUu
b+EHOJQeEVPWIL3CUgU65R8KUMiOa8ahJ1KV/W/Vwt0WwPrC+oUZOGvvBeTJhG3H
un5UcI0wRTy3gQfhyoHxcRJ548lvU3kqSaWm+O6oEU7hgRW/ESxzoBzO8fcBUaCs
Quvn24vcRm1fJJGA95mcrMjq4Kw1eDYkbL4rXYu1pI5WFOkE4NtZfNv7Bg3t823J
zqhlYK0J9ATY+5c7ZwfLirKJQJqn1SLTcyfOXH08ySP0pip+Y1dLygQknGdxJ/bF
ceY1qSTxDWAcAwOzvKtO52FYnAkgt5uKJ29VZQn6CHp4M8+ArHDB5YSqNWpI6ZGU
pJ37fgh8sXjXlS9FxrB6rJ3I/3wpfyLfZH5rlX+xQRAcqpvHkJ7A+ynus60tUgw+
ngd35PnV8x4pHvwzx3SsI7X67PSvYsJbdZ0WiUixU2mpF/fx9HCtC+Xc6h5jymHS
S/8zI+XdAyGuR+MOGzzChliog4CYdvKC6NBA2goHkc6v2zPtgJz7GBTscrBvTzGr
cWqviettLdXVb6LhbevLFGVldMhHpYGSIrIKWpiwVbJy0VM4dBiKCwC8gfPTJVqj
h/b0zNPpVY43PGFA+/MSl9aCeOdDHS/Tj3zAWVMraCFCzlwbz8Uuod/cojIsUj1X
7Y0LsQNeVASKdbj+o8E38lCIlpdMJk6U3+oOQuLU6/CQIEJ+j2snSrtywADSg3db
NcAmF1lrUZsB6UyJFpGGJf+XBkmRwdS3sF6eDOAy+9KQxGX+LWumO5dgWjRLiR81
wIQtVGCQ/KWr8X+QoiDFSbATA/L/uNi7YQp2m5ZzW1cN8oThsq4Hqprz3anHvSNL
qFIwQwZ7q4EiMD7ZZfR1vilZxox71Sbade4MvD93ZTqiFz69oDNT/u/y/rSj3HAg
PqR0R1o4W9DjhUGzX1YzXwKTk7qIwYR8UhVO9eXATlPCEWRL4ApdfLyDNRDJtKZp
1b8OIWrySS2k+2hrxbz0rNb5uY24upSXefs+nGEBK3wGij00YG4yERo/tlKfLRtL
xzdyOIILHQaKVyGawTW6MfvkAE/iH/1ruE7r0RHMaJpjim+o+5pmMeOtSODwJCNG
zk8xdIwj482saR9U4Ia9BF+1XZSvLOZdQaFNnfyIHBFFM+ANuXJKIXOK1KvHWs+O
92R4i3zKvuV0eqZhXEV16XFbn5o53jgkWeailC4BbKCA4kKjsX0YPaDvw2LdEsWt
UXS5N9I9CjsW8k6xAnY7e6zOFCMHT/cwEJc4MpR9UNAIrxGroZFttQoalQbW5QU0
n7PGRTfpSQDg1GMF2dGRkM7PeW2HhbF6ZX80y1odHPMo/MbICyp/GKHJ9Pmoyz46
/BBTJQyHV/+BLl2I0/ODozHZ/+CIRUVwJRJGAEQl3fzk99DdTyBHzUVvCS4NVe3j
HqLTUhYcLLAg0nNcBv9M11vDVIOYW2Hvt6Q8z9yTicxK1xrjeIid8ey2oQ0nxDBl
+v7XgI29JtlO30eo6K+iaGf3RLgrOF5xbsHYTrDErHnfB2UCRyDoklpnXMwzbEGz
ZwNGulwkO9VkMA24vhEwLcBRZDsam8knEeoUz9f/sgR/sQCJOU/6zvalnyCN1pgs
nXXjSVXdl6LeDpvMiG91J/PWgGQIUfCydNiRqzeoR8F2fK+/cVkF7B8AkD60454a
SfkHJusW3tqWDhxDcmuTLesEK6E5XwhtY2+nxrsk7oZ3S0jQu/jyDHIrAiqBWJjq
oF4lyC+T4oxgtZ3hI262OquN/vQIIYHupNz1OAoUB6/PltZvi9HDX1tNJymgBS3f
vNjZlSk/k6hNsggd5UZA4/yND4x1sUonBZr5P4nu0t6N9vAhpCG4hkoUdgbpA+oQ
a/EhkYYEsE/8BSw+nPymL2M2j9m8TqkYPd9WVvzFCzhGE2KY2AexItYNvhyq1FT4
EBZvJGPFLf37HdsT/IMuCDsh1iumKpMHo5TbH4iBW2jKJObgAAJ4bmOEotfwfklF
IvDfspO4J3vfTqoCPF2od64uFw09Djy7kDeUkEdte5vIA1fko01MiXEvx2HoVo5d
fwf1vngTIp6a3WkBtsVqz0j6cvrXtgpTMbT9eDHOl3Vo7G7H2zpAB8bI4Bka6LmJ
uU0m/zQ9XtiSd4PBotIx0lp/oSHA+9OsEPy1Z1hPQWmBSFCxhIWIrPn4rSKqlFbf
NSddfoYBEkOf/G9coZx2yYa2f5GyQ6pn1p4O4t5SbY8/MGSI/I24hh1sX2f1wR/4
St/VyTMjOoO2DYAy3OgwSWqDJEgveLVhckF285j94xnr7sewNILCNCaZL6yJh2V6
UIj4Il49phagrgNDNtY4mwVklf90k5I3cNmZ85gS/qt2fP37bmsFR3pWVfLjEdQb
MVxwujZh8IT+u8O8cJ1uHuZlDALuQzdqS+4pIVWDrAe0jdQ0P2uoJRRR4/J3XXoy
/aP7BaN71mIvlOqWGRRx+NkmyLcWQ+dpDuKZw6jXbeH3g9372YyDSYrOK90ZGGdd
fi2JJWTRpG0EuuwHBiXbLmVzs/N3/qDtmk4Mh62TVLjbAJQK6NBQd36KNVKXWJCi
8qre81h83pyxHqL8W5OgiULRdg6drPwLwuPHCdl2voHFqrtsXW97p937tO2ZHGar
WswVy7a4ymSz/8N1GqBIwf8giSPVprbwnNPopBsVDNeZwnW2di2CsUT6tUq/EMaG
wHPV8HqkKqAa9TA4fpSbPUKBXKu3Qliak6OiF0CMs3UgVQ3lv+hqeve1AWijgKRj
QfTQFVTtDWF6i+LRPx5qMY+khHXw6/IjszZq7rEwHTCVMHNQwgsY567tukO7tf+t
+3hdc+vzEYB5yWWHdaLTRAd3RbH0D6Ox64K2JANsBuFVJeM4ktZl4nxJZhoBi/g6
JbNd4+GBx53ZJFUlC+Be7u22TKTpJNrQXi1Jz0bHHeW5Iq6if9OMqalZBh6NhfIY
hgZ70gRfUCURJtyXZp4rAxr/kUeu6lwrb5N/BV2wWx+g9LViYSaMoWgTVjIIufgP
RGDBEoxz92ySUktv7wAOopwD7oSAJQpdPowCNUetsd36tvrebudltBQz68OWZf92
7w83vvfL9lobDaxpDv57oAE/LA4x0/MzAvwAqlOwdkrV5csrfL1VPJ4ap/xlFkni
o1eZFavaItwV/8Vet66n8IOrWHVjTYtxF/qnEEXYFssYVedTD15/VjTpgaQRMgDY
PZfPxOJtHc7w9Ys5lCzcVaNOpaQ8E9zLvwtNPR5dsyTFd2qp/nGfiazEYCMOSxU/
np+SmCHoebiYbPxtG6bQdbGOcT0YLdKn1jTi4D+pAO8fhy6W1y6C4n+p7SJOngx6
bZLRsvliy/RZnRi3APO4cNSHKZZFsB15vYocgC24S66I0q/rIFi7cWTKx08FgxA0
DjbzsV6RihRm4ZfeLpzv3y2LAppxmMAcrIMdhrSga4axWv0ldlTbyeoWeYHc6M7A
uxTYmnc/6ivKOelsxHKzNvm5QeXNL+xqmPoSLZZd/3BJxODC+MAbsxqAzWR4UfzW
DjdzaKNkKUpELBKcmBFqdS9GxZGisqFceOA8CBlufpvbjeNNhyEKLQB+srEY04uz
1S1qPBcYoSHfUGz8EOaaGw3hyjIXuFaF8mohqvdEmnxEnkv1aOzdUBnl0Kq45sMj
xedvrgX0S8CEWV49ncNFXQsPJMb3GeOLBZ1DYw3esEtizTt+gX1e9q5vFK+Sw0x/
mh78/p/LxXZwHOljQ3zXefC5TrFL8pE8GgSDHN5G3Ta9fUtMVvy0qwe7URXCwz45
d3kkY7t7YYUwug3hgqB4aMx28lkOow3wcbnynKHRcxjX574wy2kcFSYo+0RQ6LI+
NGorl25m3EZf28S/tovzuaaPzAj1Uy794r4WfrvQi8u2xVd+MuLuf+dd5gNvQg87
wdRf2MEK7RA8KAA6eGhVZM1Ae2clZWJDt+T4pt5hFSG9VF8cNgVLiKiYw5vHuZJP
sXCAnkTIh9L3H3wtFv0pe99K0sJfm9jCq9tOKdfSttLp8KrT9jRCTc69hpoEEiRw
NBV+B3uCLCoED/5ZBMesLEQkd+DM4S72qRtimmVzkOJkRKFTrsIp26MM1AhL+843
v0Ii5xpfVH7gq/eqiC132QASdqkc/Bc/b/XX8DfEKWlWx2iuCe4yx1nALBh8YL3U
YTvryetISGrpWcOxgNMTdkGotRdSbBKTiSU+YZRg3pdUStbMst47X1ZqVAC5JUQ0
8GdES8f/uXaohxP9HrZ+yzn1J+6TY/Q7Ietxyk9zIDkPIrW2Dl/8BHlDW86+4O9T
C+iIqH1YX5htOHwbn+BIFb9NCTojfHgp0dBlVH/2DltNtHTJ/0z3tu/82O+AIFtI
d18ZBMvjHOLlXkbTVmHcelrueyxFpEffmdS99VRw7BQIasI3fTBvfD8kqmxvOgfa
kQ2u7AU/Ql8q4M67usi2WVarNzR9n17ATibVmdxDIlqZly9u5NQi7M0cIwtEXfAn
OB5ZkKQAERJiDiyBAH9N6Vv4gnr1f+I+LLeneeil0T0Y13q7SAUNMnSKkN9RqoZ7
P4sZt4W1OuinjfPgCnWRlpkEWU3ol9V6y/oYbb/+3eA0+cpDRljvxmbSLXSVcSNY
T7rimaPW8mkS7xhZ1sq+lRk4eLlasf4mCJHRCOJXrVeZcFdveuYdyqOgh4eP+Dta
rXW7lRiHjstaGO+1HEFRTYBaC/J0gYCYjfXe8PPVavZwZ7r2+09+HaJhdKDa0EyI
OdJO+bG4D7/ODgxUEQUrtRQ+hWZqYLZNAn4YVGIyNVv4YSnRGPxY0vaP3ta+vlRF
iWJ6EKwimrqYJG2pbxpCeznrNhNg+duSE1Onryfn2JVomuCcjkkCOy/Rdvq+XjxW
1g4GffWX1iSxXKvmgMPTM4aaPR/w/toyYcEZAdQs5O2d77aSCAcSQX0SNF/bwla7
c0obm9tNYxKNbwYOrYj6IE+x89JeI/5bQ/97cBJ0KhHh1iHWVG5dyBXt/uLL6WZ5
2IefbOVo6gRKIdutU4GJRULim4ChoeX47R3HJm0MwFtOMhaKYSx9c6pcaEoPqAAF
zRkK6g9E6JHFP54eVXSNB8Y7RXJaqaWXAkkBpW2TGosMaQc2bBIZR2yZzi/zEm3x
vruX0zOVU9WERId+kWeyNoa44BaiwlsaJQ32rk5qf7JTk4/n0z/Vyaw1KlPNZQrS
ES10uXMpgyaqr3C35eQlxyAZapakyRrZIxHueO636ARu9JGKQLjnmdhO3Xnbv5iV
NqUnNmcvGQm3+K4j5UXOGjwZIVhulEgYPRlinXeBsxXcGLpTUPAMTyaM4DlRPJ0L
DBOemK2UTgO6cVFnCtHP7Wbid5tV+oa2zphqw3BIrGEPcrjRzRPCumV2y0E8W3gQ
ybRRpA+o03D2u6gTD18pwFMvM/sjwNXsgy2hqbQQBRja+t2SdvzwUsyDCpOi30Xx
MAL7t8fExFy1i5w6PwyehLrNKqj70FUfboqgeJn3eNjDvWWYR2TE2rBR2MBfcgqk
YsHrKwO0V4MZRnBbpvM/V53y6OFJ32CeXHR1es32IqaObN4Q/SeffmJEl0N6uX7G
PnyZZJm0DfFROqSqcDoHmkbefFFMZjONQC8G5l++r3ut59vfFkbcaB+5RCjPPONL
W9Se1e6BZvXm56Y0BR4pDC5LA9IO9WCfh3v4gBdS7GhboUck65OJNwZ09bKrL74h
4pFwr05X8AW+FDLD/mDUb1zh1q78OnfQC+gJkazSJIH8uarCXcqXEyo9M6h24R5w
lvRXxyfk78Kg4wEp9Kkv5/hx0WFN4z0iLpIHlkMdgFz4y/HG2v6qOYmQYGW3Y+3t
VCiANwI5TkJmXdYiA9xe75vzph6JhBNC6ZQBv5DsDlpGZ0pHs5V1U76z7v65SKp4
j5DCqpaO3Le9OOpUnPrP7/TrgjtuV2R703twC8z0dQlZBK95hQ3mGpeXMRPbrFxR
z0wKpmVArCPYR2gHhFBc8Zq72ayb9/+pDUtdQam2ofnKoN67G4efzbb2m4ek9HZw
q68pUea+r0tT2CyAToavknPhGeOhI0LajZDrVVBBM9+gcML6rlk6C7r51LVTYx46
WIkY3gyxqXE/Glv08ZuA+maJ/BHHuIH5dC7NijUuYDwZrAHDCn9imyLRoANSgjUy
vqNPTGFdxKcLhGkE14xbX4W9oJBLQlhDpH7uKcz12QCUBa56eCrJmKWbcBLhfXXh
CN0EXnE1113iU8j7ZRhFe0/V1EfcBDz3xKTx9hjacPdWMIlE0VL8vJ738yiB5a1e
X/q5ttd8KVBXxNBqFrcvNSYF4UT0m0+JoTh1HhJ8YnI5xVGo+YOne5UCbX+HCaGv
hOuDm8WJ7i365izmJDv+tc4pro2QipTa8c0rVWf73xXJZoPbbWSwnUVI4x8z4roF
u1Pk+I/HSMFScKF82kfVQyXFdCncyD89ePMdSDAnuS9tGeq2msjTtapwesFYgXI2
Vo7qN7/HhF6rsZ0HiF9dTOiikmM8XX6AyBnJoVWEqkcU+ZLUHZDxmDg9mpmcld13
pNDxLKGtygwaXFDtwTACT5EZNnO/yplWxhS/Ya/neYHVR34cyfIhi9wwQvpNSIbf
ro4faXKea97yTt16OAWT3AR/Ny5EOxYHfLd6rYHf8Jzm5aTM0DSiYyqjPOmDwhSe
bkd8ij4VWUQI6Fwo1S8TC99UocXNbQT4nPzPdtMUvJ8Wwf5Qv7BgIxCQL2hsDnUK
W9jUROI/2N9lXcs0sOAsflBQtU7vniNvEeIt9iXx9a4w38Zw5ecr6tkfQKgRWwwz
udm3PgEuWS601Al0BZxRDAwlj5gVgZvxPyk3PSpn56QunTFA4KHGnAs3lv8IAgdP
26w+/uOrwfzyXL79TRvn2iPvY+O/UTo8kMs9yRW2d7oLRA0Snact2KbQCnGq3Pjv
A171+yuxw2FueuKMSRMwn4ymz9vW+QZWH/ymqZLkGVnaU6M5Hy9BxS0oLhSj8Shu
DUJPELEq5wbdgCovKA+Z6ltDX2wigTYKItXgGxu0ld8Wr6/x+7DqScJTWf7HBPYZ
1muWKaezHA9p/cHH7Kc1usVGaEsH9ZgzzPz65AtQMEoMuhFR318H/9ZNBeLuBG0G
PYYJRqklQJf6jtza/NdlmI9oOBGRNhy5beEd0B+uNXlfyuKuluuNaPJkOWJLdWFj
SyMj3Zw4096lrlwFn9Hrb0EaFpOFSF5Laj3vA92YF+OQ8JdrBTcxOHnmMJh4Vvj+
7uD7JPsYul5nFJFMskTlMO9MGmbgD2Ev6MF7gmvRvrObCtW4476vNWYF8TcjRQEN
meSkBTKtKBrVNkmuUrRyKbpV+xY3flqHI+IramGHorLKdF0ntRua0HzmTcJYOqsw
Wknyw61dUbkMPot+MHeLo5k3+XMwOtiOgc1V42CFF27OUDnbJtuLrmLVdQpAzYcb
EPFiSDdZl87hdiZf0LHv6ZrzTingfZ0nYbfd9yN6LFGEjnFRD1f6dRWb0XeA/IBP
z2FXhjV6XiRKou7FJkGAGwacJAVe+pcf4ufAaRcXOGCFEglbk2Q9uu4wfQDnuQR+
TGrkDVXIOmkBVzy3CWSxniBKJ/KSVdR4+YAyo5jbrKumzus65TdZGI848Zr50sz4
YFcCeNCLYmrefFkcoHlBnxYpB5lzlUoH8+IyELaLo5r9Z9b+okXG09mlDjwZkjkv
gN15YGwfgaqdGY9VKK7loX0T5qTklyQzcrqbRTo3qgFrF3mI6F1xnZyhPa0wKA73
vaWrX/UDPdDbNxrCdirbAc51VZqLJtTBDb3RRIZYJmND/lmr8T4OJ+wBbdjOPEHe
rXB4+8YKIPegXzPWMJgBvN7ItvGQRZfyAyxvNaQn30/erPSS8IQw4HexCHSQSTk0
5qlEQwu/1J0DbRiaiMiD2D+i4OHGaYpN3kHuQ94yCfX0J7CXtkWgHppT+3Bstbuc
N2crsSUirasLxiV76vhVWAYM+KCuE0fXpY7ykSX/FPV0RgY+8KJGVzUAH6LN5EAb
4+10jlw5YYjmG1GUh9ifWft/wMvxZKpN0nw+zP76Ofr/H3zEHDuqGoQzwyZgIWQe
6JP823T8RYQF7S4y2QbFLabWgJb9jU1t1M/tqYb0luIR4+R1ufmt/J74hKmPOs9z
TEzQNvo99UEoiEVx5SvNKqVnCcEWJylYpHEXsx6+N9UfLuhl4HLsSXrdal/XrPzX
1ajNwO+hYdqDhEH/q0hix9EDQQ0Y5qjWmm1NTFzPdRyy1deRrIT/6PZPuJeWp/Tw
96I/8UEcE2W/X4vil3VSAs1t03/1WP9GhpHtXAsMB7wn+9Wu2jX8p9B8Lu2wbjr4
5hJwIOf/CxorVTHl2d8iW9gYhnSduVoWdQi8TJwxSYKbhdSCbYKGqy1s/fD3N8dL
LTJoYHcghVEjazYkQz32aKer4ilgCjWccQkFyqhwtmsjfShpNEjIFKqkXG4dA83S
5wsZDkHvmJAA6FB0/iXJI447J8g5IDolXWLw4mghVBS8EvAD5k/TEkzC6Cp7kaDA
XQQgZjs/6mJ3JT3t15rKR0vbM2Mg0BgAyJ/m2gzNSQnB9MEIbRiYOjS6wf29NZi9
6giZyrBTdJX4SCy8k2KXQxmu9TJ/UKgFsJj7X219VCGGs7HshKknHv62n0tu2sNV
/zkClsqFImZ9i234DC+PsWr91UXYE/ttwLHu+QIXn5H7dYiytWCB/941OIDtGlZs
AtTt9dc/GBmcNpEkq3cX50zn3kD30j+4JQr69po0uUEgR24fWIvZN4hBej3X8GET
cL/KcyUBcsHJW6ZyuVH5AoOMykT5SMRV0TAw5PifABu35jYOebezM6mXlgTALZse
5XPd3ks9j6eFTrcw4D2eMgDS425h/tw3D4RjEpDYXFXBj6vBNlS6kOZP4kBVnlky
boFQvwMn3SkMRyllpPC1Ypc0K3s9WT1fq8CNVKUfgZjt8cPMhfQ+0OU1cZkOQKA7
I78qOMXM5ADH2hNjgMuS6UfKNgLD8drzP17s4dPFVAxLJoBU2TgcjJYJkhb46rii
N7sTcEA8ZRnhyixqduO/tckC+kmzpyRBCg9TEDok1hJHWETaiu3rFYyd4EpX8Cxg
yrEgc2P7HxYXAhq6WngEE88oJNU+NPkgRKWZFKQgSwW3AJFSZ9LVg0JKPX8kn4UL
KvRlQEzgzd8XlR8ljtn7eYAkV3ySwulEDj4k/ZcfNh0+X+rTiOKmXp18JZW6+Jsj
N1UwdMfthopdGSxHKsOzpxC02vKWGqsQWttizeCHPo4y/KUzdG+7j9xlw5tIyYFa
RkJNF/i8UQim2HMWHlsYZbuL2/k2Ilg2UZiSkdvfrxuNFNWO0233TwHL3jcfmTj6
XXTp0+c0HZDKMI6y+keV+Q9wMcCq90qX1rYHbtYBVdAlTVFmz6c5KOLm+SHJ45GT
5Vk7v7oQdfKDZLxFH5G+z+sC8NDlne6QSVXjjf6pVL9e2WRn+cpM+HkzHroVoCej
4s3rMO8wN9JTldZEzCKG/LLrD2/ILg7/YS6ozZTUPFkfOW+ejFCFftXEtwuTzYa3
dSUicik05pc6GSWHSaw8Kjvl31oQj8k9jlSaF2ZSwTXW5Wngd4f/77cV066YmRZL
EJVPzrLsVGPDPBWdGjjp9c+hbS92kmQZqnRA7VZ7XFtQmY9O4VQcqnrVPNTodyi9
2XKjfay7QdUyauBkrS1cz2VUWTapnM7QKX+YPDapbY8WCPhroTQRHieBP2U+IXap
ArI8xbyIzlmsxToMs0XHGeHQRmIDTu2IZHeAFwJ4LoyT5FB9HPa5lDdjnATX6B7p
JWGdVZGoGd6KBe9LE90OxpLypgtTTSHQTTPkz0WTrOG6qMse0jCNPJ2GIiVzDP3W
upgzCEX4csiJQOgY2+gvbykkgzB3Y9F3/HQSVytHcV5ddrAPHmKZkVwNwvW5mwIt
Gdtp5IWmHhvRUDtkzuItneuRp9ldedfIREHeyMhbjdsAhbo3irQXSOaERZKlAW2W
jRBWQVgo9QXidZoE5GE24bA6CnbGYjhYRlKbR22c5FyCB0C0H2OKk0aZA+83j/lC
vyackVTuN1A6FnugIToByWSendZFad5Py8jh73vQ5UoulbAy9gjw4Fx9fLvHHqfs
nVlmrh6qGfcot+K3sC9ftrlSUlU+6OU5ioQCYtfkQlBOCigFs5rAkvSZxKVuQJSt
IMSMkwUylGbBdou1NV4+8/OafdjKzcULKsIG5J71kjhBMNHg8t8600ivPQQbqkJN
meZY4XJxZa019j6GaryLQTM0eofVLweCu8pPlM8v+vzLislwF4pqO8YcUcNeRVyX
YiI6UTqvH1nRycn1MUuy+5xn62iuIS+avDbz5hNqA79eC9vwWNGTh3omAtteRo+9
AajvVmpLgSk9oNTYNf35Eew/dE6M1XHw5kk3RF8pCD4wRKBpK1jov+j/C6PofP5g
EtO5TbPVvOTVu7JGdl2lZUk3c+BEMj++z0jJXO/13ikKwQYzaIX5PdhxgJtcP3Gy
nic0u/ckzsYxa85StmTOY2rP3QP3XYyq8yn+eAHpPpP8wDuCDSu+GbeKHgep/hsO
/i6YDZlTMu2O+g+5yZwvzGNsUu5cVuiJS4605rLzIl26l4y+umZj9nomZwH5jjFD
fl/7icZvMm1ZofIcT8qHg8LtDqtmJhQzU9zDSRpunx1PhZ2OpSM2kjZJaNIR62xw
k+55/voCQRTs+sZ/Lgpn+vrz6qiPQoUhhBr+Q/asFLyIaADNXNjYKteRA0eGgvyS
/yZKgEDk3sfX6DyvBxiTih4GTDJKvwAH+SYF88m2UcX4LpL2Jh9AgIcE7nOU3sOZ
r4g1DC9C9jgtDg9iYgOjTKwLlSc3uD6UMMZh0rvs1567bRdoNaVGhxEhLBs3ml3M
mstcom6zToX/qPBLbk4S2n9M++RfypcZ+RYe+aHB8VYdgqrErjuBuGrmPo9Kdp+U
vW/eFAxCOv79lT8O+eJl/wu5TcuWcg6nhXWprD1YEBpSGtW3FS/KybFxC3fLK0Up
Aqz9yGPRRfcf4wSt0XLjPM+Fd16MlzzmI8hqXZ4mC9PA/tpseGsRf38xZLpl6xD0
Y99r2gubcZiqwqmNYm44ein4dGNUwsCNYDwWc979IJLqJ9cUKtjuaY/2gv5IGapK
JdZe9liphjFJcmrVkFZcVGtU/x8IQ2fHWeMwUgY7XGL6iT2d6zYM8D/RuxQzfydo
T0f7C0cmeKAmVhL7lem7V4TYogbNEj3MtN6gJCBshaKv14c+qV/LURCI4D9Sz7lI
1IISYW8rTQnkr2YpjKEtyfyEX4zedvNGbuqdfKFwqN8wNtHRmVoa5Y3dH0y5Vn2F
SS1pNtIiftEBbzVArARAw8fFTNp6R5VCx4auRHKZtDQ+KIvF11iy+cHZA8H8MO7V
fRhwdSxIJQf3zEzldcbcu0b6YvAGqsy6tTrXG+b6ACY2vzsVH+ggdlSFUvbh3wmU
Pg975MpYT8psvS6LJK3HWVqxLGWrOqPsbs0vtiMTKnuEsAE0+4ZobmJtgF1102gA
ebwolM8kpPsZI/Imxd7KI9b9H7hjMj9SqbtcjAqU2uIeZH5+OA6PeIsdTNEWRXFj
qHHSGtjQ0ua3nra1H7U2BOvC/ZxZ/1ptKKPfkkc5PCzfhQsEcYhyk9Pma9thf/Z7
PMH15h00N/kWQu1C53hMzL1xUooWmS/hjuBxyCs7q9dfzhvD0qqvrd4hg2h9naQN
Kn2E+q2nzqU8kbDcPDMijzBw8G9TNDzAfiJKFEFDjDRyjMCwML2xfXOLSMUL5WW2
XC+uSe1wcVrtC8fZAbG0VZqQKHVd8HiiyqVTg4DH6kI1lQLWfYNZ0tp3n/7yirTG
lt42SbBUopaej4d337LVk2WPhvGAQ7HpN5vn6QGrElLPrTj5C2GCK29bM8C7KPY9
kiMg3UW4osyvJs5Fkl3cXaFqHTh2kLrbD0FTIBFF8dy00igAkbEhmE+lb9nTi6Gl
zkxJVyAra9szcg2xrKPxNHtBxsnQqztrKoIM9UngQ5hpajeiDnljYJDsni+C2jv1
GUCaUFGjOmt7wfWooeDhl026xJs0358iplwcoUsdXhU66PANQjR3Xa5H+zeIFRqQ
IouCUWfTBFSHzoRY1rrS0zvO1ra1eRWXzbJ0vZARhs9c0DJZNQQmBEfLOOBbqUZ9
m5ziLKnsZvwJNz7pUIobSY++VagcssYYXQpvVbXAwaG2kuZiNBKOqN/sm5etXgRw
OoCoYTOzVYNzb8PR846ncstnZHwt0J+losLSfTQ3D536dA64OSHHV+j5qW1PWQut
Z2Nkk+txZ75KrUrsS1XpjZ5ClVprQdsvlXvIunkyRnVuuX27nMflfRUlaGq973It
L+TJqg05UCx5mjkWn099B7epsfvAPsLCTaU6NA2T6qeoQxScSeZMBCvCsqf6r7ri
KMsdOud0bhgqG51UeBtE71gpUXk+Zs8gq2mEEsethIwrpwrDZKMqVlHIOPB7eaYp
jTxhBNheMixGVJAA2LwvgEENksBgo72Z38QQTRIBCt+hWF23WPlGckhNIl1t//b/
DLGL9IZeE2xUPkL1URDnykPySBmsl05a7ZvwedHNxA6m1TylPcJJ5fX1QNM83nSC
D1NXEG6wOLUCmpACYgS32fF4JLDnUA2jLFJxrsueiMCS8nUEQa7u/+A64JO8COh1
eK1zO1n21r4IgfYBkjBHaoIkayQEXIb9tvIYjWJv8HPCB+lPJKpXoyZGCR24dmxr
3RyouiADQEeJwIUA/frUv8SOq7hQhGcZlnCxszmRfvvx1/7iQu/ig0yT9nTRNozL
J3YDNcaNwhKmDby2y44hTbSaHld09QWXBJmHxclnYsBG2fwWjZdrXSjldE/t1AHU
2z9OZ7neCHMr01ikn/x7a4u9UmgUgO2+P/Xo9uPA9PbcSe2Hs4QRpyoOpGUY6hhr
rzXdIFSkNM59srBGt0x6946NNozqFRPvY0/52H9oXr9sme8McBMD6au9t8JTeVrc
hO1jy3GnMGWr5E7VVrhnV0ZhQpusPCfkcerE+Bnll9icZIopeU7/w/3SPqj9cPem
UXhy7J6w4jMf65krQ+g7Nsl00LUhulgVj9o5ViFhq3+Lm9/yH7UhMqWsTxcOahkM
Er/p939C4cjTTa4Labcek3tVmNdf40h2F9q8kLJ/qKw/OGPSAAKOUW1DB9MKYrVE
HbeoOddsWJIhYO4NocnR8s9ul0WDXI32ngzCjRdZeTrI8/MErf6UiAASRPFvJt5n
OXd8v2xdNYwpI4UBoobBJRWUKC+l01JEVnrMUtz83GzACYyIBY2vQFOQebUL00dr
PEFRCluA2UtuvdYtSG6szSP3CmY9mBffvLEOS31bHuTYeqNrpNlZFdbpMYr6de1L
npYw28BepdFiz/JSGvDCQPrxphOshBdO3FKtkxF2rPIZt8zOLU37RAQX/gaDBH5a
xy6eQqPlcTdjtNMP+pPdvsXOkgcfhFcz+lVUOgYoM2dlyAb4D7R+O5gV+GokbBJ7
mGwdHlrCbk+NHgb5OflHKM5s2FDWzFwA/fdnR5Hz6ZlWNJ5Sril/5E7YPmzfyega
Bp13LwgXm+u4YjJuSeWzNyC0PZw49woeVK4DPXZkFGTqwKW3opnPrhj8Odno2WAz
yfR6lFSROu7PcjK8N0+TcTRVUiv9aXClPR9OgKvEymw0KrzQE9rvCWcylVs1USHn
wABJDmImsDyr1S/3HuSGZjc3VTLtAk0DioKYr169jjZUN1j+zaOJv7DlF6TsG5BB
UF7jeWQ0qSnU+kQLtf79Fba3yRmpJBxzxIw1qJJeHzLtnX3o3ar+eLxEhs9omkld
lZI0E4e14NhQuMYmNxzolURnH6HaOGGM7EZkzAU2yUgvQiuIgCzlMTlLFKE0XCBo
GwVJaoyL3xdtYnwtzkl5ba3ewboJH9/4AVp/bHMBFZ4r6zFddJ8WN5ZIgwivl5y4
AtBCQEugQlSzMTsMDIqAHZ7duk9TJwBuJjg8v4ENaKGUQ06FdIQZlGikMrEVZ509
ubYa3vFyQHJxyajPwBlX5gMHHMgmzT6O+IM9B9l+crdpJuGuk/4ThJObpUZBptV9
If2ltjuY1izNyQM2vOWy2P5uvuje580tR3GZ9yZMpsQp9gMtTv3QhYII1GCQP0zA
e1O33A1Tk1q+w2BykMIDy+64cUqYAG0zJN2b5aj6tyrmWttaFgwmVQV/+ERcl0Z6
RtwKA8Nd9W+Ua13EVM+IOBlTYfhlvDmSbF0Fq7GPISswpkixAPx9LQ2hdL8Sb/UZ
n+DlTgNo3EKUimN172HLCnFSRfAoqKKAhASqR2TFbQN410xWxrE4+kOLNPS1MVAS
M7H9RKZWyL87y58zFnlddhbn+8b9WVhJuuqepSCE/M78ZDLiD1B7MOCC8zYp/7/I
xnJ9Jm79UoTNWJHktGtjj4iKT15xnU0jQGOanY9eA4Ykgs6UWYdr51Mg7uPIdyRn
lZFfWYKiYCcDkAD7xbO65k2NbV2S8++0k/uAcYYt9N9FejRqbziXn7JHrG9HIhuv
7+YPjYTqDYo6xD0kBM0XwVCh9GES9r7zBwjsSSMs2slfeQPQv8w1St8S8lXVhUcD
Hs/2HQ1fGQ9J1JX6td1Hz07gCua2BEEHgscnUTkT4jB026/q3yH+IphLo6Rhgmg/
OqRnc51EIytld5iTGbLitUVPQaIG6ch3IFtsXHuTQ3KKou5Q3h1F/UC4nVBuvuMD
MLK6BaOJqSEoLLThhMTtKkIjfyLlXnPxUu2Pp/tb42RVboa26UJRGonWNOlP3/AG
kj+v6pSxh61n1NpXbrUiybTW5iJLv/giz5g9guSn6M1Ydw6HgbRIO84WPHCFuA2g
cZUxeqlvQjjO3RRkyBowhSStdyiWS/Pedi6u/q1oUlaUyai3J5yPcw7JpFIz/xni
8RrNaarbFxRz7wDsCPuAI4AnCG3HjBhH3nrnHSi9m+f+zj/UxWs9BDC61m3Ad28Q
e/tBW9iUzcO3uzq/0W6LQsntN1ffLVwqSEhNuZ4WJ6jyCzIv3c2zat6XeLmZXOQJ
TXxyF9aL3rdcxZWoq14IeFTWctOnkr104yTaLqRCgs8p/kgQbstgGZyCnPdvlH4X
hw8SmbycUKbMF3653MJC0Rraq5+jA3F2VkFa0+Fo1Ixxm+DHMYXjNktOINrzeap2
vAyCDQlTHknJYoGNPpIMgga3y3cryS7RC9OOK/AN/Ce4ODEICwf5unM8qoNK5T2m
0JIEg5tXmsX8J31THyUj/faKhkT1sKs0j9N7a4SlL+VFc/i6EfeMFIHVzFvtJR1a
OQRBCneoV7tf7K9J8qpILNHJLLLtsjqGih2Sl9XL2JXXGKJt5acj80SAvx38nnO7
cbnbwjxQtD4tkCUifiwbH16LHY3bSKQTipau/RJgyepIZGI+F4IsqTZPooy9VS9c
572RpHCbi6yDxWMTK7WZPBJEmpKH8eRjWfNLhln/O7C8QD8sbgvzn35pa+L1IBo0
2wtisB6SA7E5N7yibHSJWX5GXAAAxw4FDcjGdglHu9RKEt7SwwImVGDz+POSghpz
JQycKpltMDTqhBbTccVqU6AlfLQ4pmQLrSmOu9WTQUyYN0JLVQNlcIqf6U7pP8Xc
zvWY2fJXmQ7naiDjcClk3w/T9y4teGo8immpm7fpuCMvtVga+f7Cv8xqcgiROmeE
wUxlHJMEyHcf/5/TiSldj0Nu/3re0gNZ9zyjSSS0s81LrKWEXDjvyLSdDoj/TYkn
UIYDXGMrIfBepyDDXhpknKRbjW1Lhgv6NoYZDCv9N8OKBzXAV2R+3KGGm+FdTV5i
IfvcIo8Nkip4aT0K8h+x+j1mYKZAalSm/OnvgZMzQ1FRmVmtMZI/VlEV6oaKWbnm
vdA+/+x/ON7nvfbxAok2Fh69Q9CWVXtoVHULE2ZbYn12/K2/fLGqOfovGEGazuE8
oieaFbUxqtRF5yRBUMR6Vlo1D4ORbpkAUYyomIWzL+7vvFKKSkj7q3epIndXObuL
vKr9Z4g4DT6OPcSCA7bWzM+JmPui/3mekOaMuQX6d93bSHHX+YYiOYnU0kgleXQV
AHkPXsVe/HoGc069An0vMTYUG7msNmU6cUsIQam+RuZeEUpTjf6f8ljwjnr8FQL9
YO2B8YLyGGPt1lb4svYAQ8S6NFrHtgMNpDFB8gQGmowrQ2x0E3dvycCselmebxHX
gDQf3jkF8A7CO8DbtiRH9Kfy6Y68llInCXVUOmEXaLj4eXa8E8a6DIEE+5erRcZD
Ya7hLV83mZ4R5qSyON6zCizvifHbk/5Kkmsy+My7hCm3lULQMqPRw5tM3yBtaUuF
iXf7wSjs+371Ps9PtP1vEjkGzvusa5EsvJl2kLp+HDtccJW6W4AoCBvwVbniBIYo
GFx0WKpZfrWrbGD25/x2GJnakEBvzLYYr9zLHUo/xxBS0bd6csxgCNrDFGj9kJH+
/jEEIoRJ632LcHRHv5EwEutH9qZmPgiP5Fe68AoZZJAMEKOso5tr9uReE6zt62SL
/f6EWMCSmOJR/53SPUyPbUtjycAsAqCcKxiaHqZ9NFWm0OCa957NsOJUdXDoN7xW
DEMrwADTmhkjh/SXRo3fstYqiXNzfxqOh4IoteSJbbtvV71EyKDuLLXi4fvndsdE
g2f0ik4WYcGFYqMdVkHrMs90YUTToSzg94SYE41zzioVHNowtjqzYIvvsFDS2dWC
aOfmWg0sHTwLVeL0vqWoed2UCK5FJihdFDrZPyuzk5dDGxcNpin7q4tP05uVZkCD
6kwq5/LS11p7uyHqNo3Dg4DQKptaAJbv7OIz1upF8wBz/jICyke8LMRny5bGT2vh
1C9pHCZMA5+PSuy4YGBVaIOP3KEAL+abgVD6l2HdImZGcvs9mB2b3f78OlgRu1aQ
bMHJGVc8FiJinLjkRRJUoaSJuQ52feD3VtA3WiVdHyj/Foi8wSKDBUXm8Vd8YUOV
wslrK52ngZuLfnaE0tF+BZEF1GmlQfJabErjpJTStIxONYK7RbAqeGBNq1TOA6+O
jre8Hxnqlo1iSb9V3CBDU0WYL59YB2IYz5jzdHG0P3I9l2cvaRwuJspN5rmymt3J
ozD84yiEk7PfrMBNphF5P8UqmTG8FFtYU+xIwML6LeEk4L9PF+HcbXHAWR6+Lo/0
RiboD7N2lzExpSkPbpzaaAVG5df+oxgQn2hmAZIVAVxpK7hGhTVABTL0+zK7/OT1
6hu3K6iUen8BuoylVYEVWZE2eOkiuJvxskDUKwkdsipLmapoXgCaIlMbPXYzvuwM
yWD1zV4qC6Izpc/rY0jQOX1xvJ/9h3QOKpX6j47/R7DRcQhzckeDstvNusDCCTWP
8qlFxJGX0r6C+WUiEpWXo7Bth7QZh8CaT8szM3KRiPPIkNs81wibgczHE/ihjaTO
CFOcw7MhkqFT740pZfd+GCGsvaowz3SFwSd6SYMSoxse17Tx4YUFqIN+2rQy9iZM
Rbbj90GTnVAz24FjYd0gwkFa6ZuPridHTg0hHC0Ik2b9iOgeJzYLhtTRaHfUR9QA
G22Fli8vuiXvo8Tt5lh25b/vJwH7nIcAsbWCU3v2qsMKnjCX6xjRMGhXVrZorIMT
4yRVI6kzia+vGekNHzTs3QIZ4DFHqcUQd0Z6sfofIUBMrqtdVI8e0w1ZOXcxnqwE
EYIuPbSqzeB2FoS8Lnq1qtw3Zl14QvtnfamZna3sczRLVWq6S9AaW/xIuTms410T
wYzVDeB37tn+O8n5LPL+7GULwWBituBS/5J3ayo8q/wGNrJT0tcFQyF7yYheGXdV
PeXFhL+UB2ISD84Z8kh+6tetyjYyRovW8dGVyOU5qWeudD0Q48KOw5H1niEoFL1S
A2e+wn5Mz3Ct07djwGcAQWKP3oehHg4ZZLunQShuozvGMYtFhhAeYJnF2SEny6hm
074LsXwrqoynbogC/+uBkGbM3qJbDsBHlwahdssAE8OljyXNeV3SI9du9JMY4jJQ
TJhcSOBJn7BISbYHQm8uVF3DbtkOhxL2d9kmPjPTAqcGgiW6XSeqYFQKn9Rb8Qmd
PUY2Ta25SR9YhbyyjvzYnFIRjjnpLY97Mf1Dv1jzPP/LtmHks5zeKLNxwoAA6jcq
fZzmtrwgUfrGVYtHXu78Q6kKYMJOKYs/8Nbv15RGYL+nnu0zqHlic4pQ0OMlwlFG
JNh4+I5Ggt/K69Le9+vb4C6GCkpsufVDXtO5n7wSQJpl6qn7fblXHM7fLJcgLhA1
A+k/PNM6YEKCtrfqgFnyzbY6qWPvZGIlmHezpl5wVbSShPVj42zkpqZTB2fq5+CO
LuXCfwRNR9p5BR+PIb5myZe2nWtJJ3xJvRgxGHDsG3l9r1rkVhuW9T242ZK0Zx7d
90mKqjWAObfvFWf67DBS3ztdB1asy4rzW/5VyYwYT2pjhRdDatRULgcU0irIXreK
yCkIQBNnRjjWqugFovz3eUsxlRiUG12uEi0ZRy+tE9n9cl4XsKXPZHC1VH4IfgqJ
b7OrhQZyOgFDrapPZIHGD1qtSxcjk2X/BTsUtbuFku+EC16yz4mtK2D6sGyLXW5I
0l4lgn76Q1JLpP5O9Qhk/VEcPyvYmPYFzVlZzFy8P4Pfvxo6G8138J7LaNmHI3DX
L+7dA6hK8s+w6v7gE4cFKz1ugCci0GKV83qPdBmn1T5juMQBLyDdMktjid4olghj
dur2CUBR+hnIoBkihPjvpNyp9ap+rAW9AOGqk4cE82bCxP4lBrotJgwEOZibNi9S
YzveGklLS4Z5KvUaB7bs35YRBPW5y9ixtpK7HIRyi86L+3tQ4rKtTjoq7FQEKAQc
aFXjGgCb9wjTe4s3eFJEgVfaeS37DVMFVDP1O9meeeQqHcDnUEyNzer7IMEIJ9t1
SEcxGjjSYl+riUBWQfbVVelXxemQdx1u9F2iv9tkqifJWINep8ZkE/mXOJZi9TnH
z77qW5fyeS5uFcequb0Po+pZ/ORd4X/zI3KvoNIP7nS62ii27pJUkpCmSwWRHR4H
r7e/odr0oe4pmdZPfUtkUVG9mgn0gGqRGo/iOLj+HNN6k+y1mQD8m+C2T6fB5y7O
B73terMkvpstEAYuhK0pVOUN5ksnfAskNqKup6Xc7D4FPPnFRhygudo0NA4FEJGt
PJHEuWwZuxTc0xoUOzC0lJdhqi2gp2fUa/lLVLqQRWr+LJt6dHO52PZfiqNPBHgY
+GhsZwdkfhnvXFEKkVwZFDCGtZVmi4ceW5EOJwu4IVu9Q1W2BIKVICoUqeZoYBXK
Rde8TZAciNNVbuNew5kcwlWlltr887vMsIWZPWjIg5enrToFrdU5MkIV9PvQ1QKr
4oASV7IvfOmAzsoYMxLcHOcgcKo1vVWTRxsdSdInnw0T5OiysPBuEyhgwL6sjwRC
2VtOxL/OOxblR6KNixJb2RDuMR6niU9y2L2oO/GllPxtpLUwua6+gW3re2USWQ1K
MdHUOl4DF/+KZzXRe8zQmQXyg0an3awGAPPmT7DJbTzEiMKySBy5kyjuNfy7cqSq
Kg8NPKN2WomBrV/UGIvfVbZB5kN0/tfTuIi7UEVGqheed+CBj1MWvKiCl3/vQa3X
TofXlV3+Y801oJc4ps9wkuOottRcye/ywNxL/jnF4e4iELdqtAYQJZ+hllRzhNjT
ptJbyYCPm8IyRlCO7Fz+GUZlOWBiSvOgWfLEIM1oFejxDEfhToxALmOOKe4g3kPT
fKwmbCB7oe+z3Ja/396W8BrMyBZx6XOTmm5t1WvGKewtoqI55GIvhpwcojxVCM4R
bX49qWXLfTH4V8bVCZ8lSRq/7yIiADUW4gHNX3MCrWZ/kDBcyz8ISxMaVE8qzZ8+
1x5gRvd9HuFPXea+ODNAnhksa9W342y7jU+Wk4fw4ZKLj6SfTxmYIo4UZZeA4mXj
I2WjeEDOKNE4kdD/4/jkaJhuVNeZjUTIoydUvPkJSM/WpbsK+9uej0Kj6KBGliop
xo8FBG/9KP2magSGFryCiuST5ofJq94CWPfJ8/YQ3e7/4DFh9OEhz2QEgYoA9YCT
w4rDA38b9OxuAZKzPuVJRDMoEuIF7wLB1OP2ShZB03RFpF2aywLNjkmrvgt77XVi
XPY3nV5TfT1ZzeD8GDREw08u6xA8AXEuYg+V4NPnAYkMN232Hbks0t+IIrYPn2jN
8Xny0mKiHO7Q88SFL6vpAoWb6DeHLXpCrRd0AL689fgJ++5O4xo0ptRAxedSkyHy
WBYYNXrrFZKkMW/fh6WGZ7CWlWOFdaotK+XALRtok9+ZNGfOfyPY+k5udmjPSB2t
YKkt/GONHt4gmNrUO29xgkpzeStNge1mnhz+1t6aLwoPUHy5TeLFkm/QMuP49DOY
SmDanI9oogTfrcbnw3rhORWjDWhL16lC4OE66fVzB+bqnFosiZtYjbNjMX20Ntmu
MPnLSvIXzgH3PFVSDbg5GHbOYQAI2Lm8FaTwU1aqUuETG7jD8G3EHW9POCVIy0gz
AO38gTUbvI0uI8QCVSojji4+r8omEDEP+1oAgC/JMb559hRXdmWJJfIhNj2fCPyI
X+XCf+olVBC7Ra968oN6625oDyR4rUuUW3xHKi4bj+bTTG/1DhzU00qDb7MqTrIb
fE8ZwSO3V5vGSd0R2GLt2wsuWFy5c3dpkZPWP0/09mVojdXcVBbeXuaLo8uNDHku
h8ViqEQsvAhQFEDdpN3Q9dlngV+uCkY8IGIT/LsUzbo32XXkIV9GOej5YGn/3u8H
sjJhs6CMACPg2futzYJYxcPq1WKl4sjStBHfzOv2lZ4Tuqeaun23U4AsVKKbTEom
RTwvarnPA96DsNBg2hzZYgVL5Ma34UcSbu2d6n/LLAmbnaGv0VAr6sObF1Z8i8v9
Z9l/NkORQNNnzSiG7ICWxln8PGudYPi1Zi1auFPOSbBR7WUd73J/HffatmXZ0zJ5
6PLPbRqoWQoEFH5ndBW562hvV3cwRibgbuM7xc2fRCTNjSzvA3Cm0k7hwZdA/mzz
LBkVYdaWG52qhgsAJTg8cw7HtJIoyTuV8h6yAr7PIDpVxZn+eux2dz5pArqA1/vF
AgIDHCNbVp+v3sOek1GPPYHkDSEHgHNmXt3+b/KqrCTXprkGT8x/haWL+Ycvrqor
wUThRexUvxjGWHhZZUafjUgSIC6xUuL28tWjmXPfECJHBh9SfT1vvdlLaB4gtmSx
bTCzbof4U9SzLsZzahEd0j/OjPxJE9RXJP8IeI6hsICS5WrClFn2VnHJdVYLBcdN
hBRD+T4RJItmwAlSN87f7kQOkAehvGQTgSptArYrzPGZv2WfVoPaWMyPdbv+wi6t
9llg/IAC1iQ7BuZt679Q4zimmfq7P2lDBx9u9p+69JMUVxnYMsoABMDaiGBrenFK
t0BVUYrw74eddFaRgXO2Qp4foQ2BWojzjDtSWyzJoQS48rEzNUvlBAGwIMLRhCI9
iDVYEcfCKgGMvZn2VoXwldKo357x4WxuDKkpENNfc0ywDM4PDZ8K/9EUduPfvpN5
N++ZbWeaGilKBkjdzJYRGXK2Acw7LsSCPU6afBTEDg8U/YFUmJnz3pd4SM0NHLNI
hrd2W02UX7ZneKESAt0GPtz94CAt7U+UIEFWOc0Q9PR759wQsuqeb2NJFmdShcd1
wZUnKrYbXbMdK7bhA/HKi0cPbilXxyLL41p9FS26zARMYGSbZmi+pG0cd5yokRyG
MT/tagrnOOz1RKhERjZwAyxjJhnw7Y5KQmr3VpFO4wtGJstbCQhvu6XD/MICQDOZ
EA5r37jIK3Oppj0B9wuW3RwU8dZeDu1isx5L4zR/EBFUN4tqVCeQtP5ER40F/93Y
lgZR7m/TfHhi5gvHKMAndXQ/VwKqa2ih825sU+LlUIS2MDzRavY+h25+ZgPNdiw/
c6caSsNuyDIBl7eKnkL9ULQ3A41qGVTcsG1xUXg5PxWCCCqELZgyiptjSK2JHnTF
9CsnTFpX1lvIUmZYNG2YwkyXoUATkBvOyPsAK95urWJqF0ZNNXSfgK/6Q916DGUf
HuQeRngiOdnNipIk4QfVRfRjeq/V1Uc8b4xRT5s+5m8JrLLzNoQzyEojJewga+md
ie/o+j2bCEM+ABTu1WBQMIcoMqmt1wYSNMBqn3iGlytkRfWYFTBkkaphZkqwM6Cj
bN6K4O9qwePoS7QpR8ylg8hnLV8encsqpPwf06nYpgzgPXGREj9r60vqGGorT6xi
xNC1zD5Rp6rh8vvWP685HjKVcP6QYPvKLz5oQZl6Lq70EkFzhpWI5WuxKTUxYio4
n6MSPP2AALDd9mgjosCswKX0Mk8JFXfSMNXs26c18QAAQk6ry/otad7hWgKfAYYx
MtcnO7yalTe+XaWzNa/XnO5+mM86HPw2+1GGRvg6jUsc1VJOXtSfsaeXIYDf5O6f
nxOFALtZS8oEA5OuMq+cw0GpKlRBSGSIlWdMfPa43bzt3lBv/zwNKGKdDmYVW9cp
hr9zOlI4eXDGbGJr8MRBpXr+hYccHSS+uqZfCIyE5CM3krVpVZ60WtMHM+FOK7DA
BQ7glwZsJklbzPsgasJi/tuKIe3V0bOgcHo+72qZ4hpwBZogj45FGdOHPqbb3Etd
U5RUaYoDaFSiVsxz7TrVjbrrIRLmZ/tLRbHSmQ7vXFGvC7KsRvNRUTKhxmqai367
JVbKaEbv/sZ43IXkMyCHG0kSaqV5OcRGwCBNODuVl6nvgr0n1a0ElaHUwv93+zgz
7IlpKofgv46RacA4AVDWttYGSylnRk0Tx3Rpd7B+PvgEynGctetRSTnSwL/RKShD
D1vE2sbwaariv3hve5NrTuNdzQOlSHjsMs/bYgvayD+Yw+Ccx4WeQo1nqyyDCI7g
wNxMlRVVLMYqqhEWpaj0+P6T68TiPpp4xGXBt16SC8zznheOO8AroGERIINHdmPI
C5UveOVCJs/AL/iIvWtJ9f5XxlzytEi0nQrriXjnqDlpVeRbJw4zQj52lH1jT/8W
MDnbqoPXD1fHMJsr6NMdLAtJ+prObmr8zziFYuM60DoB6QO7LFBtxPZvKkFKOOqD
nHRR5YNTuuExKAMpFZFtRv8T6mgk/Je52pXrfvixYXzwO2McrUxmPg3YRC0NohkR
p8Y3kb0CyhuwSIV7PzS0l+zYes2jPLqtbfmbpzGLG8kDuTNVB0RxbUMeIW2P69Yi
UZ3tpWMysQkQIS6ORdahkBVnjQg5BcM+ccmH/K6ymwOC2UE67mDnDMSsHQbGxsiW
cZvZitMdmyNJAhvjzJgHhDVVjp6MZaP28VdDvqyjTMqXrzmh8Kytp2CqbK0RE8kX
vm7Br8NC08Gt8Z2d83MLCiV0WwBSAcBhWHwM3gITjlWgeUPAAtwVdRsIb1VS7PKT
2IfOMnrCBlyRt4s8/7CZFTMEofxkeFz8BpfUbIyeoD8rsED7E9LiEIlnESOux+zV
6OBeoP0MQbAIsTjLNRuPneE1Sxgk/DM+wO1hjl1hCfRfVacFR6FX1FjMOcqMFaSE
5SrPYONn0yDBdcR3Pdhw1cRVEPLIywsm41A1kUxS6zMTLzIFbM5XzLuPL8RHG53+
+4vHV4EfEBR7gRCFH3EgMq/1wm24DLnMOo2IYVQwQacmmBStynkFJuXKlYCkxTf5
8+nEsO0g8v3qJsKOP7VM+al/TND4OCMaN/rBWD+F2qJLCqUusfib9GEoPeSzF9zg
0ibCKPASR0qJAOn/HFdqgG2drmagJvqvBgu5RIiq4iSsUBO6P1arABufF07JQb0Y
4Pk9QsTfOkbzWiUceRLm5qZPRu7AQTL8L6H9zj28IIKRTmqSLl8Hl9GW2H/LcjTZ
1+PsA5Mm46azC/ssmH5WpIYliqs9w6zXDBKvb7/W/hvs/Gh3RVhHLcMrTvchsSRs
IjoWceg+Hl4waOmnVz3et+wss4IQD6XZh+HaYK1knU+srJ6Z0fYxjwOmvKTZjtPk
GTNIl/dcxF3FShP23ecgrGrtPFAlEx5/7Zojq5cyuqsPWuGFswhpKHJXwiO+MXES
pKCFF4kSjCh+yz+y+Wp4aBUgS2aqX34C7sZRdxu20XSQVZ852HvSWso88j8gymCc
GnCAATJGGNizskkzuAURujnCtbkt9i94zDxO5iDq13Wq24eRVPhiBA0R+xKIfWeA
RXm0U2QR7MumAOSNdOZdb7R3w34lYiMspIJb4zI5jKM1+t+MMs67Z6ngI3ZNhVPr
QIxFFVV2x1bC8FhvNU9Hs4Tox24xp5sa8lHENK9bRQN1K6hVbrMp8VF70DcDNQt1
UcRa9ys2D9J3uzUu7yEEoiXXcknP7/4+p85RfWM1wjacJUt0tfvYzXAspTIO9yeL
z85gmZ1hA6frRvV1YBOzauFHIJFDrkkZnwwSsvgNRato7mFM7vGue9TxdSO9Xgwh
h1/uGSReYNEKhnJq16GN5AqrAmL2tcFWr5Kn90jlrC/c/yHISJChMN00vwS3+BYv
OHr42466hIgEWo+rthHZYAAWJtI2W5mElOetjW1JLtf0uVEINZQm4LQNYhVJm2I6
uKVgq+KUgH5SKckp9uacR+wS/x7mgop+ginAvL8QmGULuWzp5s1NV1dOauz0F+D8
SiJ2huZkD8zcOOmbPoVMFNdlUpouR9CVVmmLny29/8V4IrDFFyg8ns2/vViW2xEI
TczBSWewM96HFY9dio7+MHiS+NP1STkaQzofJxbi/rLQltj5/Bk/4R7BZJ2CBwJy
0lrexxSK3XkF99L0dVotcEPFNjAh4QVFG29xhF54Wyy9M4VIHLKW36vzf0NQH38V
j7XJnSfwKchbmz/ymI89slAeykuqqtc6SAMg06neE+Uun/EbmpAhFOlyEztB6HNQ
Xf7uD2S5KYGOns2SRhQQHy76OP6ohXixGiuHwoJCas/ejf8FTfAzWxW4wy+vX4vS
Ay8hfS1+wF2xqLFF+lIOlwS6I4Mqo76D/u13LO33D8ZSferYKOSgIfWdpUH7paqj
MOLTdL7ggkqW3GU3VPFwAHH5ECzwlbVeCV03mTmLey6DKLErlQj2l229UDPN+H1v
ffzDsDBWv7voif+SY1CahvzE9Y5e1qkHrugBc7TVhdxR0mtbaGvIgdII5AHph2ol
7So626TwVqRpUNnLpanLWttNqUXWN30LyLYDTOYbr7iQE1lg5cpHd5cedblrhtVO
CbiAPWqTsEcICuSfNpVYQnu1H8w0uS2tike81utygodEYjDAO3UDJqV/ISaA+ZvA
YS8FbrIzff/sx2pKDX9Phid7QqAXPiAP2WJi9I0soZI7Hmis01WKTnohgjJB8T7g
JLhBXpxdVqxQ1xPEdWrdhcfArLFSq6gh/YhwejmhdwrWRdG1mTCr6MPTmiWAaAwu
GyuCeczNfhl5Gh8/G/+LSUcITj5FF2AtJV8MeqDPu/z4xqhQXDFKxbCgktUS9ITD
0J+lpKJtSjhHM0iltg/7erZKXHwAdlooaCD+4AkvRo4VRVppMC6v4iaI03MEh914
W74xVu/4f3KLiZfHsaJl0lgQlH9AMvn9jzyb+JiMmRijd6YLE/gIho7kgdzqle6z
KgliTZOL165w9W3ZWfELfsU7iaDorJyAA0kZK0Ncb/HAjUOMEVlaCoJgYsgsDiGV
xeY92EX66RpjwbKt1EscN6Af7AHYInR1RveRMX6Y0NjUgyslZZ8U3xJ6ggp3XzRh
S7eldAnMkoPtELT5i3UFZx4ZYmpJyvlMP0CcpMmHbPyQUKnndQzVDz1PAWeAKTZr
CBMWowbiPxeniNNT9rnpp0p8LJTj0sZ89/1emCsmvxPftf9AwgK8I4i9KofhiX5/
+XBC+Da77ixlyIuaWJhgm7PwQPUuaMwjgMC1tjc1Sn/lCmB/GZNVn7c9pGX/MeBv
ZILk99tFDCq7uUEPWZKO2I+DxGvrJy/6iNuHEgsqaQ0uJxnJVqRQ47ywRxZjZxDS
obe3bSqb93MHSqq2y/J17+NYAuJdOoeBOtcge0FJN3c53QdZAAQnZWPShJhWTfCM
+ow2iAJ/el2WBFqAxq3Hyl5qKmFGx71EJ0/CRYWXRFEO9dEjtaZjAEEfl7uC+5de
rPitodxL4br+Or6dVzstRouK4ctTyw21ItXXNrIVl15+YVCxzjXm5suY4CLpfLj+
9CgrYOFq24pSu1oCDiKRB7nOEV9wRzVBpASzj9/y5DIUUbxjU8M8W2MlhRYa0+QE
lSXnJhQTuU5rET/upCDD6BB146THCO2Z+ZK/mJzMEak8vYX3bl52DNf++zY3hvsl
atMhnSbaAc6/pMgsnlyywAY2k38kReS1VNKY0X7dgKQc9mjYzr6VRZ9rU7624LvD
YU3GbF+q4ZhxrV8SsAxFFBI0SOdtcTkSOOhzI9myJaFmnj6jLewJRutC0Xji8Spw
Pm8mtuRC3JCQ/EKj5WkAykUroJc6E0+knBM/fNCNRKf6ZyaFum9mBWiGnJmAHpuR
1AuQi5CQIyVPutQuZVmnccltL3gWTuOfCsvDHm3mmkOZbOZubNb5+ENhUyrcps/w
Q3DTWhQXWrm44vnMIO4P9VifSKlFthAUSzKYiP6LfvpFEUGdRVn5RswxVjUmYUb7
W4a5oI3wYZqLbVV1PWlHEhM3Caq+BKLTnTzBoiT2oT2Mpgv5dvDbdJ8Sh42iIHLD
/lqPzKcEctQpH2Y3aIqaoO3VqmF1rkUR7wRWxdpN2OZu50y9uazdJbPoI2VTEbai
+LqPVkGncjw3aw/o+zluqz++qpGP3R9auypSST1G3ZuSqYxggz6HaGZaFNQL6Jx0
Zc9Zq2czSlb1SWJsrxQo9AbiSWOF+K4Qvl8/KkqO22aqZw/DxB7wodZr9icB3FI8
OuAMgCb02uWgL6dcHupVo4nV1SpB4enmDGbyxUInxF+HV4QF47AM+ma+2w4JKqsd
NeDWu1ieD2tjByKmBUNmWCIfY4BWvbX1a68MVbsKztOUFuBLbfGg7fBqiP6vkjVe
A4w/qdoc0us8ImRuuV8flcNPmFXr9hodkRHwiQAOJPYizWMbB8ZDT9cq8VXgOV7Q
9scKOs+lgudz/L0uUSRJ83vNDAkudp58yBKdQVg4wDP2ryU9oQqZeIs2pon0R9iI
mMsNRNzmBp3XoFWTzOelFR3sfISGjk8v3+pv8mYjcd9d7av4pnppeDjqOBYVGup7
B/COv3/d6vHp+Lj0gO8u9c348G4/bYC4ZKwchoX0DFLn+uZEb/VVbEmIy9DofqtD
KzFq0RfgKmofUE2uIKW9OYDZ9cKmd1pvGfbTKVrYzRH5LLzRoX3Wm4m3+q7+98vg
/srK8CalWX0rXsnIZEtqRaG2x2C9NbykQXBuamZj7h/NYirB0YtPfzdkDlBpdTaz
WvTk7phgSBVfD11z+dFP31yLVv0FAs0Kg++YFyawVTbMAEoZdt+FDaOG2iy7/6MV
i0PgxyydMhpT+MBln3dGhA/5twH0NmI5MGWInbG/RaDb6pIagldGBzPs+fMV5ONW
oLccko7izB9s4nV59mXwk6uzy/+I0kBkax4INeXUEDHoDc74HgG9kvMxbNSwt1l5
YCM5HiyNb/Xax4eTw8+SC/muiWyFM/6BVNnrXzzGUHItWUM5OwXjrenJKJymNxmh
okNcBOkBGaafzZevE5FQVPd+2gAMYzBfYkxiQbxQ4gtzByse0f0LMBuImRwXVDo3
gm9a5LjcgnCc248+5M11B0CtFn4/ApK91vIPfSvQscLp3nclkuG/nuCyZJd/j7fR
Bk91oU7SH38aqrW/Ji0+SYGIcCjp5laptnGfCYCmCp8bkdM0ZEg92sPZv2WGjxaJ
Gith7EtUVcg9VZChUdqD9amocr0tr5c38KGV2NJ9BlhlKcTOvs/aLn9dUcSuhkWa
2OhYZ2j0kAptmUO77LEtNvZNpIQOFU6wmQBhyrvU8wzmPTqH6O4UfbILKZ1EX+6E
Tjf0gs52DT1uxdixXK4eOXFDfDA9biaXy/RTw37gqHmIiqzE1fu8adPhDSehIeB0
JnBGn4totAtgtUIJ1kYqmPGeJHlgA9yDkYRrG/K2aSBfgky327+TeeSoXfqVCt3g
IJdNZV96mKJTGsBUWtPLpb6l9/jobKDjIephFHtvknpRtKFtRvSGRDfWYhAYhvVg
wYcDPPrWztLhbtSeKx9+CYB+sMLLMiM4HyBzxQdu7WgnizB9AWV6mCFVGRHyqX0N
72oY9UmsekRwHMCFu1n1cgZreX0BnOWG1yLiucCqontzXqYIrq5oKCDdkVxb/zOM
OCQbo77zgPZgy+NVwAAnExnxHJf+TNoEk+O3WJg6Gju4jBsRFrXRInBwLxexnbfD
ZJ89xtPVcmcPjZrpaFOO4Ue19auKAgusq1PXh4BnZlRhl/USU3pnajTwL2EEEnGu
EWg+73fw3H8KHfJCpA6rQn30WdDGI5HzQlD1EmLaYN8IpFBtPwQJUd22lOJeJ87X
KCsI/6z0zNvwbXJnLvGeYHgCiRqvFEyf+H2p8vsOlnLvHFh+jVKQg7fix3fWJSmj
C+x6PsPsDXnkYiJzBAQr28/f9Xdr1v77VJ2BzufbEg6W1vC2TkbmNTgpNn0ixNhP
315jjW/KmhZxtvho8hcqIYb5j9UosOnfR4m+4782KA9D3BU0uszeTvZIeWtkji8t
dLtQpMvgCz/R15hLcPqLeZLfkJrf25F0Xsn6um2wRuC4R35fxfNQQQx7CC9M2nwr
sNqWWYDJSeT6YRSELwitwCBXzsBvQd5WsIEUG2kNQQwkIEk1WLc8aEdhB3QNOVbx
igRYMxi65MFmteOU24rKAQzZf6ejhUXcNddM6dU64B3DoFYU4rtr6ju6xT8JQWTv
w8gR0pLbCVPmz/qD9uWWpdK6biAsWR4LiK9PWEqzDfewonxiT9lh2ZRDfZ76JyxC
c0Zvva9Ayqou/kklJyPNzcOuDEZBXAsmLl1KM2CfaVCOksO8bH559KuDCoXQppdy
n2bb0/D78431lwEG0LCmVLS8tBVeKyqL91n/jvEX83WeuIV8qR9/UCvao8GYpFLm
RIQNd2+qLgnBob5CKGkyfrOFhvPGRhz212Hm932fId1sK4tLF9wmvpbPA8IwdRZz
jLJVhGkgdETDAb6jw0RhbsxCfP0SDSX8z2xIoDwd0DlRV5GYVP1j3KWSJjLl1UMC
9g1ol2og7mun+MOCAGXfPskluV2fuDO7XQWr+uV7yMXbE1oThrjezn5P2AvJYzMm
da1TgWqQQ3FRKORnxRKMFdTYWxx3qCH6txtPkKRBWMk+CJTJAezoAeDBMySVyi4c
2MnILRKxlhFPAEU1AAQi/BsfJPhWrqYEHZD/g7hVMJiJUU8sTuT7atj2zt36Hu61
q5FN0r8nPZal0/gvonRwxbZwIEgp5GS3IZsH9GGmuPqeAJ2vp3VZbO6Xx6N3VTu7
OImboBXHdUmGfYMFnzOUspz1BBl1EMi12hxCmd3Gr7h2N8rLSaRIurOpoqjMH3QE
o7dMT1JaUSDtBWhSd3oixlEjUme0Swh8oKHXLjrBc0Jg4M6Pvgkx/eHbc39cF6SB
Q0PRXnzQgM8eG2i8PcxoIQCni+6TwE0q0NEltHUqrA+6VKR0APavKAkoUhcpTKo8
kWRneM6A+osWRa4noICikKtdvR5Wj7jXgIEa6nsjTEiDDUa9t8GA02PJ0+LCWu4s
2XSMZJWF6hMRAUhvtaoyCTopd5w1GTkeLR1TlKDOt0BGAD1s2XH9oryYAPmEhCZW
3yeHx9UfR/R+xlsC5aRHGUWdVPlkDM1Nla5LEIgcquB8QkgPE4OwVutAhz151DXB
8IhdES28XZkC3prHPk3IQ2SaOeu0JTSszlB+VUdRKEKn8SXzeAa3WjQtbqQnFKuN
CraDIyA02bM+ej8KL2VjmsLWFSlN5ASJZKrbBjN2TwjEXWbrQ3YA6w03iONtnkUn
72EElyPz9iRcoXZEzdqm7gGEdE9YF/3csWpymRgWvKvesKghj3q5wjpKDOOj3RoP
/hV0oWl/6n/BU/E243rHwvcF6WgUfOgkTkzt/bHDszZHYkpYWo/Xdqa7jik2naoJ
PE7SF/ySMGL8fUCCrHF6pZp3P4wflTwr+XLmNvti6iYs7gA6eZyxoE8QmqBk2VEK
MFXFOQwRAkZbvd4L/RY9qJi9FovsP+ZcLsluGg6V3r36lzQgDPdIxcboaebmkOCb
lePGEsATjBoTOwD2ov5CwJyci9rIHLSpPn2OEJCIsa38w+fTEN1xLYcDkcuD5n4q
viMKn28zHSZurYNCiNdAwkL6kLqr95FsNXLBvxBN3fg9wJUC4fan+NYkNOCzeg2T
EwmA8sFpVo6dVka1+WvZbBEhNCLXKVUXUKrljvKryPcbSpWxmJ4a2Bs6DOQNt4lM
qlA3FL/1G35JCllGVKaWj5mTAhiDZNpn7FniOMov2mDf+UyNDCTiKyCySGKRsKcC
kT0lINO+ojSFObOce2XoryALmLhaF2dPB52k5jN6LWwfDcK9FYPByWJCGi2sPbVN
a2eo/23we9R38TD9szMi0806D9YFREUqIhPVqvFN8M/cE9R+PAgWeuPj0+Ybb+G+
DNGoNOJ+aVND7zbRak16KAtwvo3/FBO1nvgp/BrVVMMu+CldkKHeixXI6+M1vlWd
tp/wNSFkfvJEECuF8mQXc3x1QWiEeWSAyrkMi4z2AHLy1642TKo/pfPWKZS62Z4Y
piukgvfRSZubDMEzzOKn3ad0FiuDeQr0cRcXWkb5dlemO354l83fpErgOC1GIi9A
o1CH2pm4eCXbpTbKjEhJgoy36ihzWAsbzQOaZcwzccg1IHdbf19s1BgQYDTxHL3m
JJeGeeG3WaiIYCP9D+kUq8wYuc7vZ751b6gfkqGgpWLEbWxQhaLek9QZXBiUL2QP
JOkjsLjkn50PWX8DWgnabK/eBS1+jmRT3keecB/tJ0V6M26qShfxa62jrGJsBGdH
TPDYYbmjpRJ/9DRsYt/my0Z9A0xNj2BgehrjRJcTiey5qw4SKptPAICxRPIPxRy0
jD81OV0Pjn+Udw9DPd1LvWx28Qxe1VOKDkAY2MwzRIftGyv5iVTEqYoTE1jzV/SQ
Ewl6rFHwHeWsVZokLd1IcCWt3aivFS4UsVNDmzMy5iY69D8ZzVpM2lk4BE7iianH
aOXQ6gGUuUQaGxUkzFZBNyc+IZ7FJ59YLiGuNXZy69j8aPc4RWKVRDYEF2w4Y9AD
JvOA2jtFyyS+0epHkMnUsokcIfokY0dUnmBw4XDFE7K3J7kkBfEMXR+vysh/N4T4
arED1Dff24CjGFOp5OweeUd7//gEbzzhh5R7/44O2A5imrms3ptqUtlrdXsjvQEu
V8G8mfAto7oqqsTHrya4J3GnwNFmQ1yfBJHJQQM6YSdokkRkkf12sC72hxF7a6hY
vdw76XihtdhU467vuipJ9TqUUvqgIA8fU4y7RL1fZN10IWjkSO2FsBxUbqhGfOJA
pjmBk+3zRhZECicDgRnSqMnjwrCfZfVPBx2F78MSChxl87iB/5yQlprxpYDq0tCQ
w6R3s0WWLYm9EwwlosHv9cO3mUPTc0uVsDqw+RXx8GSFBVtJfSCiieSO7HVh+sI2
jrqrpAxHJpU35rwSJjCwGdNWN9bT4yvFKxyYbaq6vA3VOgpQPjK0TRn4p2vc2Jac
jlikc8o78OmaEkaF6+DFioco8OkE7VYZW0HXf0yzf93r1Vu056J04yVpB89blmDO
HijNiWahX01hXcPPmd6MCwz80S2a/TMqwnxDUbcc1qUyFH5RnA0zoCHCJTSiq9Hn
tizNlvtgKnZwtTOTDrTY+sR8KTxdADDE9hWlG+Ipg0ExcNs02/j4XrHGSPaP9kzd
iuTt5FE/trV2ItMeQfedaPIb7DlMDlUCgQEFOnF2PdEphEaXE0aApLpEAmlxKnwc
y10qE2/okPMjUENsW4UMgczm0voSzaLXL/lXQrKfG0+tSOwZpLZvxySy1xZZ1hvJ
cPa5sRDQojGJsAGIO8k4xtQks0/tK5WmNMvY9rSyQm728kd//1o/S3yyVG+s7+sl
8G1RXLVntsiB9rK2hMKSDatUaOEH6uyfhuRGIXEKfua39Vp0fXKJrebc1mkex/Ty
M+fjOyRPoUX/wDz/haGAS9jlf5J/bP+S78/dUz6VxOoRA5wMTPv21r7uJhV5uIIP
IY9j/1xY8tQ14y8ZwPS990N3YL2eva8GPi+Seqpk2npsyCNhIgW1kB5+RQ38O5bQ
mQfzSnhHruLRHX13StvBoebOu0ocVvZXVESQGYkNP1XyiUbhKvxqRovZjDsvMYUA
D1JqMLfImxyJdiR3MUa6SoxLYh1u1YV0vpqg1buRQjqP7aGypPgG+3pwhJ12DlG7
hORSwRlMTLkxOmcuFyyHkmCBaILsRVc3xbdzOoNW6EMtvX+lmkCDKbTc4ljuOeub
22A7GWir0OVT99H31RfVPk2Kiw1K40UZOctx7D8uNkdYtqE4kTzbi3ZCz5A+GTpA
R6t8m2AJLthaCI9fg59ifFDmFpn53R2xOSeE/CIFVMro7yxfCH89fxhwRrzYiU7P
a9CzMLiS8bGGyjaGHNyU30kP3/oosF/9dAbYKZ9hdkEz0Ju+DGUDyqGAyWkIJjr1
yvydQPFFvGo4AtvuUu3FHarTgLCGlSea6yr7FZrnGfK0XQMD+RWc5CyL8YEPcYvX
fOPAuObA/7f7RDj1ByeHB2wDhCq2l2iLQ+YOrjcW3kK4BxYTJs29HOpFxSs2/n7h
M88Ff66iu8sBF6V1Q+aHOfPCG0O+Fj/Ed/aCqp988kKeaWbHEssMdGzsbd+Zo3qE
pFasRlZiKw9ilSWLbgXOUWzOKQSWHrzhMTE9zLPD+E2IJdFod+VJNz44iBwquvg1
RTfd+K1n/nCQJnYDWULoRM/6ZNW48TnEOfooTF5lYYxksFwMWM5IQ1ZHQoi8x6Vb
HKBwnQN6mABwp7h9CKFI80pvelsEWqIHGvAXNW0NfCkFhNJPf4wZg24AYRDZZkZ5
C+GnAOkERggnWP+sxUX0bw/u17FWyE84zw6tqCWlq/R3BsgpTkRMaNhkKbv4IoLj
e6qz/IVXrcwD9decKza3jyNoBy5XFaKX4hF3h3oLX2kW41RBpmA5oXL/EwED685R
rPrsyqSe+h70jc0fvA23drB+IUhjP3I9ArnRBoIs0nk1bwUVo+3Ftwff6JInlPTg
XAz0rL1nPMwNB6BKYcW6z44f5bO8vt7Otki1b2/h5wcPm0exdqr2WfUgIO76gZyX
55ZYKzmp1Qd0bEmvoqC9d8wMmIHS2KNJgWZ95cAhHVPYg+v0zv6b3GEXxGr7bcAW
eqqUMBUY1Jb4OrDdG4aDyEP8d1/izPosc+eSwDUgcJ4oeObmqabFFZMDyyOvzAYL
/daY8uA+Dxb+og6+vlGarAThPCvJt5TDoI7a8zYqPTc8TWvlyCZ9q0x3IN+ZwBq0
8j14H9wesbcXhWbnnRdbrgitQU0uGIzj1PoHWWgZpDj8HWUE/62VBMoRV0GmM+/9
NWFk7uHg84WMRgmMS6MxvEQlLj0pj1EuugJLMTrzWVAUMvjX7aLu8TQBY4GoA4yC
EU+wuVxCyWOWToN/Tjfst9WEAnCVbiO6PR1dPQA1GKrcGNSEYuUoMqWfuzZWewK+
cate5/ax2ADAaMPaYjLFiTwCvC34eoiHr9+q3HBAW1UkbpDuET12Sp0UDQF9f4Pn
uUv8x8r4R2qP6O/wcgF9IgkPUUVzmxTre7x0kEgNoy8xUH0FnDxvIUt1xb+tue77
i8pQ326IaSi4wZ9AsK1FaspQJjxNyp1eIOhez6uVRNa8sDrfT02AmNvkbS90unUa
hdIBrn9qZTBvDxBgNrBSvhBmBRBEDKDhYTBUTtE/2KA0HZ3QdoUQ5oJmsiMOrcKe
b0GugDx8qvucEF/9yGeaRQfbfjyBaERWTCOxqovNnuMzo6yUr8Z76L55iH92Mh70
ee6rw7pjxUSJ/Ky3ON1V4bC9qtJjrdWGMWN9Vh2ggh2IDhazUnouBUXW/AdmuHY5
hX6MjFsbYS7p4hqq/Z9EpTIR6VYXVD7lcc9orHoNhglI7Cgwq8zIfovcpDONXfzK
wFQTT1nqVoBUkfhMJZJDVDFF6eFIhcAp9MESpyb1362BlqpNmix0At04ELLe3qvf
GEGn4lVqgddqMvApzFunI8vJZzBjFiHfhBPKHW6EKblgmm6BidesxYKGzJSC9pQN
J4cdUBOxMCGp2ziXAlQVVn9Vxwev7vjS1+x/DI7C4jtgb/h+jaEaTW6FBOdiUfqu
acHiypvfJP1o+9xW9X0Yy7G+WMtcrJhAeTfK10qjmnBShOBZjliyM3jzh8ZAgUSm
jX4stzgPOhu1OKzrzZTB0YnZUQkwei6APyNypi2F0NPcDVRI3uo0SSf2hyUYKI0R
61yxQfTXj2f46g3v3hx8ISmOOwapgLHOvo+OesawivcBMootAyPXcuCiK0KYiqoF
f+i9QZC79HI/Dp4cq5uaaNSTAwux+1NK+rFgb01azMooCy1TRKy45DR9s+EfV2ug
4vrbkxMiPw9zFu1yqmk/kHwOQTPfC1N5zhfajM/mvjnP7vnp2fETGCkKtbuisq3/
/YvQtBlMrLmSLVa/FjbGygXIl3acjTZfT3eMhChoC9jPYcpWQELAGHxRm6Vk29O1
AfRaRNPaV5kHzbJMBYYBHLoJGaWaIdUuP/1pRMtWWEqVDR6dPi/KQoGt+41uMprN
ohYcMKXQMs5ZG9yY4eppZXfVTvl0gL4VNeXBJLXdnQwtF5Gv7zYNATD8PktZzBVf
Xgb5RMn7H/ypEqnJ3di6khBYI56DbyC5yK8gVYqZCbmGMDvM5iiGGDLcbzFq3dkM
wbSi5lITjaNNe/MnzjE8ROU6HA97LW5IMmYS0s7QplBvEjS0sCJ1JBKHpdYr3Yxj
zVb8SFm0X9zL2qzsIJ+YpsM1CmTRqF17wvyc8iGi4W45GvVOJIXj4+1aHv9mLqo3
+LcEXvLm4j7OuSdCvaasvDxKVh1Y3i2+1CQEwSiHmh/paoEf5lGXf2HUB7/fkPxQ
Iz6OSSnLzodW5Jupt4IUeRIo/D7YEgsU8y6kAAxADL3zivI4oaQy5C0UbIJdyYoW
Hflm+1oWgH2lW/QLgLs+FJApxumEmIwl8IBYlcEYNBnlq7aMeHNL99utj0y0ODBy
udm/MpKw3AOW5AC7nIzhHkW/ixBSwzRB9VWVBxyu1oJ0/o9Zt6fGHMdC4s+Vk4Y9
3ptQJINGVHTegYWUdW38lsxpDevwy+eAoy1XabJuMso2DmIq5VI7id3cQCYnHvD7
WZmdKoC6JBk96viIY9/csbqfXTCsV6mu2UqTNOX0v3iURt14v2wuMTh0dNDZQlhq
otPcnrcL3yge/4GIt6uaMmtHO98mnwVJej5pnqCFDsBRsJTNJGqzi0eaHqmee3+N
8bT6GgsoNlULnUpjhr6iUg7Cm5KJc7h9zcMmmjdWb1aXHTJJ0Mp3uSS89iRWZH84
tVnNf5Z3AMJ2jRTEx/H2EOalsWVqiYpZOQa0lf+VQY1oghOATSTab3H+jc9oPeVf
EIHlqLt9LZOkaFjNQmISef96gQMjjBsHAohNwUmHjTIwu1ikD8cCcI+eXlgjp3wc
D/FKpl0GfRNsCgJAuPqIZIfUN4BK4ZnG96jmpQUjKyU9CE7H6UhJGf92WuKGUhdb
HE3eGWm/LjbEAllAHFps7cKwE8ZXKURNsf2/jYbFCHYObqWpcu4XX/5U3ylHbjL8
Z0KKL456J/hM9JMzGAujXT/bPYNaq3gx8Nc7jOyUEtUMf6Jz9AA/bxmWSJoDd3gW
DlNhKFs7rUXSP4OV9y/hR38v8R2s0j8kTCaCJW1Qf/zxOW4nJ9nfPede8hfyvbNq
f78neb9iBiYqIMns4hppg6r8UwbNJjw7U0EfgKv+XoKuqwbkV84VjVXvslQajxPV
YKN4Bzx4d1rVFpliCptqp+mJnAHpVVx5fh2mTBK+eV9/WHjYe/Cit9yo3EhvbXws
3Xmp9sCgtjIb7dOw2OV1UpTiLBGCjY+/LObI+ICVzYF/bVSi3e5s01k7SkMNlnTs
oKNYgrEKtvpmqGxbd5zy0bK1xluc332AnViJE0wPb93NgXJURqo9NpLkH0QyjTl2
3yZHopmNYRn1WKGeQtef6Q2PB00mWWTOLbxBCgYdWnWhzFk11t/7GmxIH/j1boiG
J33OZX/NTUnmyyLWys1t0rmzKkv7VsaAhyIVNa+BuQvSM6k9t7njGchI3pxA5Owf
Vp9t+FoHIyuDw36tcM9YDIHEeGgCSdZFi9FMcZ2bQE8NXe6dIf+oUMSbJJrwWbO6
rA9z0Eik2Bl/km07d0BeZEOCxVl/o3R2S1CzWOIOSN7B7pGuZoTfGtcc1Tt7YYub
QaksX7+q0lrTMYKWBNXcLu2OVsU1ug0U94Of2sm78Vjy8zvN9WR3YwqrsyvN72tc
X1tueZPjV5dE8xbwGm1Uta9POyoFyPTv82URdmO4v8vdQMwbTJBgGyfEVVMQkEpW
RKxJpuDMOiDejOpgUQhfCdOrbxVfZn+caW7NctCZmLWP6vPBpHhjdyHB2ykBx/xg
EAcPaKP02SYet8c33pxPuDAywFJ0xjfJC+dmPSNR1fFB4czAX3UFaaPnyWlPQExH
bXSUS9vy+7gy4jdBfiKuO+pAtF3BH6LIu1xD6cjDjrtiOKunizxazRJXj75SSczd
ZPKGdpJvqhGfFj3V8vttdI69mzEFG8hi+lwn2QUL0KexY7YaxZ4Ji43x6XjtlkrO
/LSmWGCa9i5D0HrnMNtVWl0ioyNIAgO0dW/t4ubdE/uNYJX1vuZi37AJg07TchvG
SNlmmzyipW4DR4B/Bkz1XdvcYW87AmKH0VYfXDzJkWNGOVFvTezttUhZVwsXqH34
rldmJbOXDRx6HsyNpwyQbiW0sQlbA37lFYYu4elnKkMetphJ2+X9W8sn5cdA0EqK
VgVQj2XdWOcRwds0IoQLvT1RFX7vpAj5gHWyXQu2RpvYPEm4Jah8jOYaSfop85RG
CUn5QtH+6BTTr2Zy+64UgGeJ6Qo7dX1Ayaw9w3mIfcRO+sy7mshH6niPTMuNOF/T
B09lG7ro92TBF9wlAM4JbbVaSxXyf6bVKs2wEvnCc2HoBF2L7QlnI1teatNiUsV0
yEvPWqmAuVhzdGh5vBtJB2+BlLd0veBIJSn64zxMATqIpLxv8J+EZgQwdY4l8IUU
qp6XqUEOhKtPVpqoRvMqzLz+wCXp2qg9YQtijLkpxeZ5TLCpBoQGwLk2wyiPYWJM
52lPE9lRTeCT0kL9m1PkCI5eGDb0oV3POHlrDcxSQtIDuOwJUmSjLqGDjIrofXUs
IZ/xPHTwDVcuQgDVBWcahLPQZxGqR7qSdCbeok3aoPLx+vEzRdxCs+lGteWwC93+
ZaffLSQ7fldSOH1NgETawxeP6Z4t2nmj0Fs0+SA6kPuJETKIoq8iSl1HH0ygCZ31
vuP3Ox+0rdGfwdggH9qTNE+WO/tEIdpzHYO3F5fYbMlNRps42dE29H7SqiYVFbmW
zVFHNBMTpHH25ftn8n4CJLzqi2Wo95llu5YmDELO/QCpuPT8TyzV5I0Sfiik3O9c
TuHWE6sYkzPK2aBl9x1JL9oH4Z3VnQaim7HoDoXQjbys2KE1+4lwm52Ex8O/wF7K
XMLt04At2EHxslJHrG2cpKi/sW/5doVttRMFT4c3iLPOQA1gbSF4keTsNSFMP+CH
y886WiO7JLz9V+3CMxHmAH+V9qHonWBfdjyMURdGAdV1aCa2ALuVZG1xSmCqJCr9
Rft7bRCLs9d9RlElqpY9+Ebnd1Bmvbg6nDWJw+2VMVHHMMgQkT9slwYKVxr3vIDX
+n3v6CaORMBuXZdbpRCI+3CEdNSj9ByyP+Hk+mMi4C3yICs/Vr4VMfj4TVoBJ6jf
j6TCk08F85YB5qX+66seNTBysThSmJSwYj4kgIFAYBp+pgXZsYqHOJmXH5pFipHY
sH5uGplHnWYwozxy/ouPJkVpOrKa/C0B2a8DvMcwiH7Kjs2F2n6eRJeIhn2jnY7S
gnCJS7b+F6f1d7ssCC5gKb8TBT3IQc6Pp3G6si93Okoq89e90pXcVCXopLlUSoOI
HicIiq4naGMmihEQICNSCCuJVgl6Zcd37ZArrvsB6xOjalINrq/KvjZVvJlC2HR8
6Wi/AX0YO3QxoGpO0hF1Je1i6BA0mNlTuwpCR3sHhWX5EVamqO+8W5KwJpimukhD
cJRIWtNPNDxD8mFnHZRTNMl7St6t8y6WhMGtEYWIlTMLFrKg8jPeu1qJ1zyjBGKy
w/OJSFuAJd7EYBgqHiy9wxtbqjNZ94jk3YagbTbFztAqMHTizQO7W/jCX5sEdwnt
FbKVU2Uw6RoA3Us0kWZFY0SABK2E491I1RZD03qHym3jzcODIuC4NIeK60eEYc55
rCR053iowugo2riUR/JsG96Unw3xxEEWluWQE1l96Zn6MPJAgL2a8ZHmgand+iUY
8YkawEZzrRIwp/cjjSUy04ACrKakAtONEhiaUZJKuOmQwQcpVEn/+gNXNMRkZBA2
gc+R4dDgGrvJ0roShDpflO9LhcEdFxWDo9R2RIGImCxL1LAFIwB+CdmyPXcDyCJT
zZx9YOXWMqPePXyWG9ihIRiUQPuId4gCG+JUxxMxOJkmqvzZtBIMwtDTJXn8FOrN
RF6Azs0oqvYIXM5R8kwKnLFPN76e0aRghjthJb8KVQ59nlj8Bvo4nyPffdhzR888
ifTc9DbIq508+YeS69dhKBB05lyhqb/txD/cgKnOdE7SapvD7a5gFO6DL9v6IS4C
HsEXssZnuRa1RyJ/Xo0Zb3Ts8K3Mrx8nPYDomP7d3PKYh9gQAzIOZZcLsDVVHgKf
I58rJzfwESjXUtt3b6oLOPxfLows3rhMC3e+Far2FukvofgouyY242D5mdpjioSJ
fIEHRzByOC6XSWBle0SXvLro1EH9PnC2H0xM0WV7ce8WqogaYvHqDj13+5e20Q8V
I8P3O7QXafqjaPv7+j+aGN0zRChmVVt+cPNBrPsgaI+W/jpBUKVtc2c5c4WUp+4R
XACmG+GVinzINVfPf2aufg2JC6On57fIMS7QbbK3P0g4IVCbhs4P0FxQcAQF0N3w
tL47SmMugpjxvREZ81Kh3siBYKqEjAJ0b6QOPyhpHXc5fEMxuRcyxYxr6sCC3+tI
/tIfm9QFP6KoaxZuqQHVnF/8/M5qYivxFPcm5lHHyd484L8YJwHJ/nWqea//HESe
m5bh6PvFx+hzZ+9DZj5Vj0OGs6uLp62SxV2FlpFIvEr2+IZ5fadoxBdRpN+tNZEx
7SBoaw2fB5SH4fKHiaLwRJEZUcOA7+0NNBCV2CNUmKCxQDn1pfU7RRx74uuwmNmD
ePN9X/8m1vsMZepzmd7xXTEQ0cp4ybPlGvo6wCy4cb4MQoySBVck52nJGt2XoU98
BLbSYjmnzd4u/ayu3FuGkro6rcwadXg3sVEypcZa91MvHZrfMBy8t7XKMFvonDBR
qAwB9XCDtQuuLgUxlmq531cBntGB7rAcBZkNCP0f4bBP7r7o4QGJydQfMFhNpyyC
TibqkPG5Cp5mU3v9edumXTTrmlW4G28a2c2AmigVgPsGeAabxx4DnuLCSpACr8Fu
SuTtjIEBakkKLG8H6/FZiAvSzVSYABJ2GQ/zZ5Ko6naTSTMINVczbK0rJSm3edQ8
fkTeQSSgNTNzaYuLZmWmdsJRhRgPCN6Lhi+TZk7TjXbh1sHTqI2n8gI2wc03GSIm
UrwRmyt27RhsjoyXiSOG7fcCYsAM8mFjqULcuSPJUywDi7uwNodEs4yWu729ITZ0
AFY/rUuHXNAKE+lqYdLwHZdGRR2a+7EtVv8B7s9sng6FNc5TPuxjgbCsWJMnRtqF
Kmg38YPIm8g8tYmZLBJTxnMlRFQ4MurFzcn6GXacbxSlTWXMAqFSrYBoHPg0tJ9o
gP9/bZ+ahYvzacYhFJ37uUI1Lh3gR06dYtM7UevObUTAr8WWtPaeJjZtDtbs4Mbx
k+siYenQSz3b2AA5lT1S2vJZUNpeg5tUTN1bF8j6nb/jUGZLlbosqw0nfu3pdXUM
RUvDRHXi5K6SzVjg6OGW/v8ICVV1l4+xOlfnuX2o3akLUt8bkkkXpFKKywv9tbCd
Wc3X5FNw04/eJqK/2BlvI3+0Pfdu4Xx0AOviwrIK5U4+pHhZi7T9jlNlUgzhzTxL
rge8CTGcsjBWNzPOGFOikR6ym3zi+8rHdhWUrXOyB+ktRtSSrxdHWJ67Z8tyFNdl
hYc6M8/7B39ThRsFDktPbWj0GGkJ/sDNUMGHp6dqfMGR/7XzZ8e2FmcB5N4s96R5
uzWvHk/p8nslbr4zOWEh4670wpTIF6+mPIJ4DqLBpwjeKpZaVVAixPLWx8wHH3VZ
NpPlEltFDm8TD66ka5TXdrL1TJIo7q7TKAnzbqKa3zJSora8rt1e0CCII4sgCUYd
L0pajmcGpKE2sJ9i/rkt9G4u57Ujx33KrqOTpg38Z6krX7poMYTu0ibIlzHkT+hQ
OKpxvPxHtcjNGhpC9uISlExVrVIQs0B2YEYgGZTBWSbkCAfm341Y19LMJwkqWsI/
7F9bfs+4o6+8byNXbHRfNJz1+HQ/XH9SyKoie7w7GWq77Moz4XI5fPJaoZ6t078J
hfb/LKdAn6kezjTtVw+xxlwHT1DVzLMLbuKlGqH6zZcPhLQiBMeKnHVt7eGCvwY7
YPW3DNmhISkRUUR3/8p6fBtyhsBdAZjqFC+sMdoZ9+9J5J8d/6hurKUCkgvQ4uY+
w68q0N7Iho+ffJKl/YDBTZVehn49d+BTu4QQIf24diHsE4kGf9LqGeMkOggutNUy
z++xekgxlijVimbJK3ghRIR+246CULGPoFAHgkSYhqxqQ9J1tzW166W4Hk4cmwDi
Bc0HomWyPim9A7HSAlpnXs3IPrR+XzaBV50N8Ipk2m1BYUae31Bf0+4lZ7OzCTLh
HKB4OBMLcF0IY8e4lPv7NxI18t1TihqhjPnI5Fu7+WVxi8lDVl3DPIlV/hjyIDJH
zpTPFc3qS01RGzUasejU0X7RNQNkHouA0INzK3mNpm3u6XhsMdbs/YftZclZnDdv
6Y+2h8Q4LDzAmFb6ZqhTwYoB9BEtmolRuLY2rFMGDtlnbJELIDDrlV87bXyl0NJA
s+1v9hlpFFe9iR456wsDKuTL1zjBigz0ozvcerdXVDEwizsmGHwx1V2yWzG+PRfi
PhsQY2GaCW5RR9oOzvmNHUcsCvaiEJmu8Q//zWl7XOzDOKH8K0IyRuY0UXCtZKy1
GLtXIdF54lgT6OVm898urx5sNHtq37xdLb3wuazQhgo3Te+w4L/QGuQjLrKESK41
2HygOGuesXLj9Ihwrc8n7JddBIRupsbDr1vsJXvMqhAFGT5ytaQoYILj0uNwtCwU
JEgly5YhFD9k00kmAE/MG6Td35DZVP67LV1+nZ9XyRMCI7a7oQWsmRSB/gIHyt2K
hHwRCGUX6/zDgc3Eb2F+lS4tcHxw+2AHv22aukOcG4cqe9Nha1qLs6/0/M/4Ckpx
UHkFetpR+/QHQHRm7vKsITM99pllIBq+viLekir7m7Dgx7ck0HD6tKPWXGyPs98n
sohNytHtFjYRSClGhgJ97QEac7AaY7OZCLZURxT9NX6sk0NEK1f+JCepeBwHqs/i
DbDAIQDuIl+J8Oy5YMnNUeHOF5cZVtn1Fmg+mdC1oLqTCJOfiBlAvVJ5Op+6ubwl
JiuTbQogVDM7CoOtvT4F4wTE6G5v7WHdV9BFG+2szqYMPzPjUITroWq92SmzbvPd
v9VFBF06AKZ9e8/N6fq8GXU6IPKosO3l5XMh7ERkDRSyg5WwwIhnynzoA2M0yDS+
rBrwpb2ct8b8JJyNvCMOAoq0IgsQPoQ20L4XI7NM8GYng2tKM7jnrO/JzWZ5fgAX
o50+enuvMhoets/ZnScIrl6jWKIi/gwc4wi6S5gYoAam/wpVlJtiiA3dVR5+CGuR
/4RwGFqW4RGRu0lMzEj0p+ZW5uRc69ykGNryij2umTcHsgAEkr7AijQluWAVAIPL
tVHdmBGip6inL1vSMsFbuiiaxh5OJ5jrCCS0GvysjCn5srj74RBj6ICs4v1D4dND
wEDtphCv6KkiIuUjKvFAdgTYN2G2vx0FcNwlDT+N0SO112ZzpAMMNKHEjanvkQN+
wa5u6Kbl4xvsNzs2sduEkZDqHGVi67g5tNGcs1tkO8+Ozkt/Z1QMIsukuAuuF51t
VdHWGJ1mHUWRHwIc/2yh9XVaBId9Odcz+ulTMFFSdN19SwItpUpaExAt2FMwThFq
agfgOzqXtSmiNb3wcIy8lU7Olfsjb69XGjpACnMuvzC6IZBWmzfvoRNGy8257lva
M/NPJuTo1Rj5eQjN9xnJxHcJKUhCPtdOz1lwh2UY6XEbkUh5T6OJMkpxOzIK3THW
pK1ixhLMD7a+via43gQznsyCkuAc1A72+VSY4byihX/DXUBiFrK2+/cpJmQSsibX
FPqs7a3zTaDDuijT0VtAQ5lE1zh87D4zBDdlJBzGHPVZ68hCzwwjsV4w0SiEtE2R
8o9mX80ASiSMTyd9OjeA0Y2WvC3C99dt8ZEE42Jm8ehB41M62hu1QOYcmu/wK33P
noRb2LfC7P+osafebuklpFkmUmzWgzWacepxrIt7h3i0fdCOiS+6yrluEXCrdrHq
ryQeoGqyiDJC69L0vE3ovG4lLHOsuwB0HN7Qecvd7vcopaKp7A5YCYECvcbcVo9Z
rhXM8X58X63Zi4czwowAnBJmyyfSTGVfnQwzWrTXB6/CPAGoZsSbzXc9a0P7YLHa
Rr8eVvtm27w3MvuWc2dAdyWNWBSb8lafabvDefx3qqBnb2WWs2qsceY1D/lQrz1o
TNXJ83ivlYBCI36IUcWeGjxNEadnS+RNMIhOUXRpiB4yQVs5qDtSunN2UOXRpStb
sEo1V+sByjXyGciJjsSDMT/5sYUm38yh5rJ0gKM1WNXmX14iL2dM7E0tbBAzZztI
vRPEOaZ6XBaSu9vuzdsKwND1VIRmOrwjDrbgPCfMQUFpNEqBx35Pgp1JBQU2fc/N
uW6s91P/r2kVo/1zhXceTtY/a/J/+hJS/YiP2gGHZAgbli7wdNdodeAeC90PihHx
3j8DTGnYHv5Mb2TjwJEfaFj9DVl/SET/omloBlMFfqUybR3F3uhPpHKdtGTYD3zT
H0jmNxeQS5FrrCu6krssBM+NDegIqkL7yD0YOkeZzeLzhW42Ct8nBZdx44r5Fmzo
Itex3++G/mfI02Xn6Ckop9KOeIiDLzBjBx8JGrZUGIQ4aIlP4FOhN4md1E+LZYqt
YIM99qGaZtxc7/DUISgUpMueg7kqtVV+9l05ijAr0dGeJf+xlQcVj5Aqw/9e5eAZ
kYN6eSk5uwWBnJ0zfP2JlR3mNx2PRpznguz/4uY3VN8LYrT3GNM5wqcgFU3Atzpi
ruHV8C3ecJv+2+p8Ee8zYT124a4iPs3dYIutK3IQbvCLZhBf5YmhK0+4VyahJ46a
NpJ+l0n6wX5x/G25EWynmju3+KK4/GHX7jMokJjHSHzjR9FihZZWuIw/+kDWs6C4
PUfMbga8jEptza2C1uo5RR6RUCTPdlP0YQCZH1XUgmQ+qvlT4xGgazPUegKiKQaV
RoZAZBXyZ4KOnoQ++kEDowJeoGFVVte9zL6RynenPYYhRTA1QQaAlqZWAJ9+6CmR
W+kOpIjf3i72M4pxDSGH8nGnivFzGCvAH2boyQz6D18dM4c9xw2/YuYkeMmMawFI
dxPtNwtAusiRIFW2hVzC8btSuYDCKomDn3B6lIlyHZXfr4OxlAMgMzwmS29QQ/fJ
JotJFC1M3oGSDoIPGcDp5QjSGaqKPLHR1oX5UDuqPSHWytfWBu4hU2/LdppNU5uO
iXC66HuuBKyT0a+h1Vcrn0yv9x1zsjkoTLj9GTSv7tC/z06Gdo5w1ukWjl9UcZEW
dzTznpDDZahsm1Nk9lsfQ0GUWw5+DsamIhSMlrmMSh9PbFMoG3/YyC+xuV88U8VD
TvVw3xqp/0scuwmu6UWZ6jUEcTHT071RQEJnE/+/J/y8nfd8Zh3uN9ZjmbPRNRaG
/FZla59NbZQY1+QzoktWTeuNGye9PAl9hugGp2AVwx1g07XzSYTQGEejHcCMkBtw
MR/ZJxcH6NBMg7t65J/aA/bTsfYmPJgNudGKJXX0tfJp/cNrTSUA4EpQLKfc7BlY
zPcVEtyVxC+WsEhutHskZwLpY7lKsfSA/T+jqW+T9mX5p68MKE/uT+9q9HnOADWA
wY4ZW8nTbF/HNEGTIxr8Yj7kAzcc6VbeFCal+r/sctHvch032igxdd56JGSuoLim
DY5iDpVF3I58P6IYEg636RQ+ALEXdq/BI9YGIMs0oj1CCvuRoad4gyy3s3G+Va39
/N/x9xBk7LPYGpsOJEK1IDwG2lHpVBdxxNh9Rbcj10LSXsB0gJ/ai6eXK61s388w
KeJ24ntQBf4zLX3IDN/HGqB/GJYWyaNr0IKLo4hay3rH/JQWmOEZSEZvTIZeH6v1
25qT0TJCjaBJ5X6sJzpqAqgRVoLpDtAew46GMR6ghdcTfJMbUJfhj/W2frs9rMAa
pLL8ULrHjLi+0yPVcCopRrL53wgqzKrwkGRxKcbJxM3qwuMerotxZzJvqx1YOp3S
lMFxzgVKK4BCMBuaOSRgKgHiuZm0ncZzDmXfI/NB4hArwQCjEWrEZAhGaK9vLhOC
37/p7RmWh+1SHzway66yOuEIxnvF8hik6Da3VvGfWCJEcDtRB2FOGRAx/Xk6OY5w
UUvGk8TX5zeFSqc6O4rYRSMXRv48cNUU8MRXU3OKk1sX44KYRChI8UVc8tZrFQdP
/d1jfi8WOPlcG4PRMO3+3t1cvpFd43yWx/8mYHZZbyfh4AHjO53wy2YfaEeCRKh5
pINTLanCN/Z2YCkGwUjlj7+4un/UxrzoZU1CydW5yncu1ggcx7eq2RBLRWytoa8E
gSXmQ9ny2aFDSnCw1CPVk369uEbT2v8IDUGJTVvfPPxo8rWy9OX8cpQ+LwF99NTS
dHR/ZyoHs3vHnXPJuxGm/iUn/tEPYoVdY41O3/65FqyLJWI13EJfq1T4M5QdZqQN
A6xySwrXBaZKDSFh3/DJxw2lKoc1wcG6j8qEo36SnS3z7KFTKOlsY5Odd/Nkn4ht
UY71MjkDykD0/+lbxWdHDimykZ40fsCmlGx8iYMQJN0oiGFLm8Lv7ax/3re7DAHK
M4tcuYuyWSqon4bS05jLnlAk+pUi7qbvV2uNaCAuoKGrPc/hYvZMWxDJw53GgJKi
3yp1UyU9Ardo34/NPGr/T9r6505hy7lvIZVhSwnigOIngcz3iH20Qzbzjl4r2+Jk
TerOMEcWDji/RcYtSi2w3dSV8uaYaXjRQ/T7bKYTO1PCmFiyUvCQYSZzst0nrXnO
WX9f8ApZCUWJHGrT+k+3pMit4skA8SWO2+Wovvns0q6MH/KY6k9gnVuckTXFaJMK
vVsKapAXS4znL2UutcmYA6Z46IPLHJ/VVgK8giNjR7ht7XWNQAvNJD82QACGlpdB
vdFHZeIzGSFJy1xJjua8fOsHIHW95196hWx1sKvPwLs/2tbAEvOa1VX2OsKerM6z
5rn0jAzv1Z5xJ1k5MmPwpTazfCnJQFYPPQGWiPv9+LPS4GeZx5qmO67vOT3KipK7
75HRgTE1k+28h4n/V1ZCe99gKoJNZ+Yj3Pf5hhl3+uEXtnKjcVJb9qVRXI1iiUnP
kxkicR8gO87ko9u1MoHWph3SVX2pETjPvAzRnW3PHeotb3vXmogIL0mcaDEQvVAP
PE2SbI+Cgoyu6J0xkpWwaGl1I8qsdmcNFQT3lWmR1X8lYfkLbBZHZmfujEz+sNNu
yexb2YzBht6dXoz2687aSLUX2U4Dq5iUMjTzpDRnYxB/KuP7GKFbfoNfFRBYB7js
8QgdY/9t+HBdmUzurpx/iDyYxAm56j8NItdscj0gs5T4jgnFst+B8fMAjzM1cczS
2PebpbgPIaBv7FHe3JJRSYs7Fw5AgUabtmWNhkPuV5ezlN/vhiHl7wSNt72tMmM6
ZyRRCxzQ62kwQYH/va8Q3qLJf+1SEbEUOD714lvCAivcIq+W7bUOe9Wf7eQb7FrL
3+P5iG2BPBvEcPfDcs7rWSq3URnUaDIXXy0H+sYEmG00CCM6RXsPJlRPM9RGIrV0
Dxfj+84/oN9lVjbH23pBvC52zIjevBtgdrlP37cY+fvzrvMdJ3zyEyBTESfBQacM
bh3XQ3+HXdcRsTCSh6XhlNUdhRTtEvATRgUw5iQbgx7v3Su+TAlEhvWtC3NqbRNx
bTyqDiNBVCDPsc0ABnrpCTrUt2Nl/sdJWXN6ijHx5LARAiZXWfZHrjN78fGd6U/T
IKR9nsX4D2QCWhePo2uWGQV6FeHb6ZsmjoS+pO2/OKsjBX4TrzS2RIPNURbYNv2b
1jJrgV16/j2dYAUDuOPNHH5yTdohUmpjucUTAckRTti6uKfFMWxhw9Xm5gk+FUY+
8pGSiQmSkpnEWSHZatelnbfKjoSjqhgcaDEmU9rHlUZMu63atN1Edo2XbEuzmwvc
WN6XVbHJDiBdNRZmrqZEpSY7dhhF16IUCqWnEJHrX3E4cIzegGpNLc3qvSxJY+Kb
LeMM6MwJNThZc6Py57HLeCoTzLw7DJjPSVcVL4oN0xd6e2yP9MgTVBgfw7pV9q16
QqKUr8Fgk9n4n+4zq9bbaGOLgqhvs1M35BXvxc0P+VTTfqXSpWEYLI71MXMk9Ksn
+o9EPSlq2KTI4IIhZyHXeTMv1eShWCzeg491Lryp6c2akklVt7ZEDL0NBeLsK8C9
D8rH42kSGKjT8q6ybL0Onwc/zGj7+aPME9A+gbDc0/l56eu9FBa9Xuz9C5FpjVfh
SfuPad9J4Ap6E8PzU56k8nteA6iz4VPsqZ9tQ4U5fPjrIwpJzp09uZN1MFFMoAGG
tvBF/UbxpRxxIKJ6uSVOI8eNd648ta6LZHy08OqKiuvqcZw74u1uF/8D5uh4Z30O
SXvIqvgnfNLV3Dktwav9Ld/tPNrMqvSrxUkKRD9tcQnr1jT9Y9oTbao/r5dF8lSB
kVs9E3K/vBUOV3Ql9NZe/XiWJOsGAVReRYAXNp5+FFBMBGBb2Z+DaXAaM4wG0Z7L
d3NRppu21hlhcNVXK+ztY9c1kQQw1l5LGsz8Sm0N5zdB8oTvaKeAq/ojTAAGbct9
/eqzv2VKfmOs93H88xOuSMnfC1Zi2xEIgDUecbQ1rcItJW2D+/znzMl3bXrLAsZS
7br6axlgyNFnGg20fPTaP+H0e0NdQL/C9b/B86bK9dlCgWS6jSUxVqwn1TBCjROV
uOXcDN+NrmOHbqzwO6QiYuHJ8q4XEzGwjKe4vFYaw/Lq3Y6/keSAhPjz4fUTjv0J
ZXnMzuHf8ujvEIZS3UM/IuHUlPipekRGC8KZQvO4IXESCtlXnMPGKsvyWFV31PFV
UUbdpsDmFwC5z7lCRzYvnCM+kk5EDlREgy7vP8S+xLdlwDvix4PYrTI0MLUK3rdj
vxN5XQUOjYWUiLtsmMcL9jjC6K2GPGrwvKpMuHnI3CAmmenfD3rWSmRTR1rb3gbP
67Xxkw+VF220poVphqubt5bxfTulPGrFVeEt6URY53HYGn4P1qCqt5n8aIYVh9Vr
Vy15iNAh6vPoQEu11wHhma0U9X9GxTjtzebmAO/YOkVip2HgKD8WnjzD4xvCCs7d
FFFv7klEgYeCHWVAxuZVs6E/tFIUj6Qp+s24vHzBFIsaHsEgfI+IwHOAJpbBc8u/
WBP4qD9z+WvLLQA879OZpos7NP/q10KJUHMOFYgFklSPI3eLaRs8krqGaQ9o5G5u
cg7l8qGBmCfXFOA4e4z/57KY9m05UL1TBOAC6lxqvVMxGzVrX+Mx/4l12BH7ihsh
FhtGP/1YMpQ6M/EOA1esxCoot/nPrGw9DQkZc+Cg0Y/v3DDu2LVCaOI7oRXqc3yf
du5+OPZn6kNN8kqO/AKN9/cH+P7bv4mjTkMwCashbypVw9Y13nnp3MWX6m1KHBGq
UcuBBlH53ubGrlJXjaINJoqfe6ESbvwILrq8kFpL10hS4I3xqCjYv2oqwwByfIeo
pCni/UllQsRg6UQPea5k0QDV3KNP8uq1Wv830JamUJkyRJuDiJa9BBfUAFgTOo9c
sSriVs5b7oN+QTnpFcHYnR8Sees0F6b3SPBQH4wMbJWXphg8XuGnamT3LubGXKSI
aAjH2/B9gtrvEiVg5S459pRb77mt187iE4hBg8qd1iU4SSGrCjlJ3JJla1z3dlck
TpB8i81w41awl1lIDse73Ix0TzFG7zlycSvsEkQ0tjc7BuMGKvnnlnW2TCThYz1H
+tqzR3OnL5fQve9VrLPKgTTSJjTJafHAAORIAhcPpzABPXJf7rLhGFk10ySzFgLD
rbvrTyefWKixCeYYac1oRCKHKyXy26IKJFim8K18vr1hjwaycn3oJGB2ZbWsA7D3
TkOqjLrANhC8fp5GR/NBIpprTozmf1RlmQkKdZXJqoEJgznd2a4BMp9YTcFXIdo+
OyYm4PHX3yQTWdp5vxU/HtVyKk8NqfX+zl3ilhp5b+V/qDlXojmejmO6ScsBBHNh
UXuwP7eBN7bOKzQAxTkKNJ8psTgU3qykSWZn401zkDyrtaesZoVntJ0ZSRRJz2Hq
nbHb8VYlKLnoFTHxWFkgIsC+Owy48j5BoHLgXYAKrjW1PBekck4+PYo84XawgYUP
staWtcPyQXm8seeU1XcBYs7gCFgrAcGiABxrLTTRcRQ9y93/UpFJYbzI/vq9gVNA
iF5iu/SiDVtbvcYasg70crTWqNJ0i/hlPVg1h4l36MczBSha+u9JjdngFstucQyG
fdDkjY9Fl4OCyUm2LB9PSbidd3iG0FYJVG1jiLg1OA+9VDwYDcC2lW9Hiu2fc/dw
x8no7HBL2idglKbKE7WtRdhpi/m4gCZ7yVsAeRJb9L9zSunj5F7Bh9aO7xULyqTA
dxrKZhVObvTPPku4ZyyXxRmEmisMXM5yCzF/qdFst/pBXuqy93gaoTvyZt4L7CY/
005BPAJjDMDoiiHxpc2zDokjyl0VuBmfYKVHNZDm7255pxSZR8JKH1igEpRcpgCo
gTK2hNW24QwoH/0lZL203n0eevzUTihwh0l6C/IE+H4zSA6baZQQ9L6V994HWulr
ygEVscMvtC8gWkkHZlImapvFQlCT/wviu+jaIzUPp7ZoKeY3DWkvhiPWJttXOiAZ
LLWBIHtWP8YuxmepdIXMQIxkb96okZbIrOjRl/bmzPy6p68ErShV3UN5JjgS8DKH
WmR8vPMrZnAyxxTXkUAKrMXfs2fXJfuW6xTidSQFZUysQKHx+xyTUV2p+hzFlLKA
0o0iAphpHwlKigTU/wn1NbMZ1VM+QErLssUSPD/IwtdR6svAGbI3srB5mYTjLIC6
HKnHoc+f1vcMs4lrZEMRlhWb6qE757Sr607xryx7viQnLi7Z3tQUxAuSyK3ea82S
6m2RPIgVtXkD1Bi6EUhF3sfSG6myv6Nok185rXJDRKewroG58eTbDnTBps8eFcqF
K3hEdKDx2QHE0/3WF4+TwhO71ZOMZK25cGWZHvbYoLPMBwA32tsIi77fV5sESlov
OM7UCQn4oD/YfTLhE47MQNcOUsij1xDStbxIU+DF5aydbEvAMcbiAGgZqvb9ikYG
P5MCpffYqWAaw16PlGXZ2PcKrI8YTMP7KVLpZoyFhirmXAC5NiDd7rL6O1TLJBBZ
RnL4031l1to8SbMapG2QDRiBJqXGtk049BUrEOQs5LQ2n+IwUkumye+JbkC0ZSZd
HK3hLrRyBkwusJHaV1mSt3aFcm06AQjNNamymeOQAcw+5n0Z85Z1Nnk9eQcPXRyt
/89z2UsCiJB9mmNN+HMpeRwIA/MlDMg5VhxtAPaN3pfyMwGwO7J0vGdf6HRi+mEp
oFWAj7d5LU5j3FcO029rTykE9CMEQDwmsNiWBR13B49xugnUIOgJIt5Veb2aShJR
T7pVbqCisXe6lAb3zVNv2xyoG/KEihKxWKsFD42sw2nxg5cGy6LrDGBhACpRPntu
Y48p2M0ImOOca0WMRo8aaTPcuzYNOIyHtVxoOZy0nXm7xKq5hZA6b2dtPhcYIXQu
K9140uGJNgGu38L14+cEnweVvrRWZnjDsfS4g5IpxLPvQjMa+gDq8+oeZgIB98WI
YMwFZEEYBHznoGmE1YQtUVIeJPhgJIMLPwJ5rcL8ligCn1XL2HAY74zLE/BMrkH/
MojrxJzELm5URlMDohqrKQA98kc8YUBElJZpyAv4Kan6X29cck/jzHPoHXl+pGJv
93ohsfMkGJBfB/CtL5ggtrnM2D4/8HzY8tPCUic0pQ4C6Gq2R6ashy82psJuChij
m+RTwP12ked/3uDIW+HQGM8OxYotX1Drd5E/Zf4X2E3lEQqUE/8BsGfvLILpKSW5
xy3rY6qSr2y9GiTE5q5u24rYu3HvsMAY0Now2zGdjH08D80D/CJNph9PI49Hr0dI
wrMOPM8SvLMYTA/Mb92QrjpK15eGKM+kKglxjoHB/X0rs8MSSLKrbB7THwQIlP9r
bDFp1txCWoTWKJyA4oTokNiBv/PZOskdorpvW24zf5xFk5M1SdKRtU8fCPASVnHc
QRrQpkFxy5scHuf8WZkeAAhrjCZGjG/+p0wdO9XMOesWPnZ1gbMqp0J4hHzqCAr8
lm3p3Ty6fQi/OWaUyYKWcGfGldI575JS3kD8CUXm+ALWgO964T5HBq9+Kf9QOwg5
PG2YVtzJjBsiH4ub0rqSiQyJpURiA6kD1kGZ0Qm4LyWu93Y3cEFxM2eSiUMub4F6
f6mP+qbqvqfHEuVz68xzzGvTGXRK8ujEvy3LeaP5uwBzFeNvtRXsH1wmVz+IveNX
Xv06QYYaIv7xYN1EaVICMk372Wns8xML1b+D37FZmLG6GstbaypdMYuy101vozpX
mjj38I94X+FyaUF+5gzR3LM0fjRPs6Q0Un4EtH/mTZFYJP56WwobIRmU+1SQS0Zp
aW57Ns+Jq39J8wo+66b8kBKEADn+Ygf2clr9SuAMhpddCyqJqa+7eeGD7/6RrWPh
hCoIiUtcfu9AcWpkhQjfPB8Pe5jVB1KXvivX7QZyo4O7sFVGpBoTa934z4DdT1Gg
0Fj+u9CYzA7wzXWKJqAOiuOgHa4YcWz2fKR4oZBFkS0otqdfkCIQUCwwOww/qNhZ
/Df9wJhQqXTbswoQuST7xg7/eWE3TveC2Odhs6dfGHJ7x1MvdtmC7HVGbtooMCU8
4YYJlF0iJMYcDlKlUhYASCpySXTYsQjN9I+QJgVl8UQraZ0/YaneWYe9jrPbvE5W
BaJHtMINA+is+M7o/m6Grh9hMu4A2nNUrXKdYDEYaUx1mFx5qIYYaJSUxaxAvtXn
MfvHRiShB2UMiJTorlsmpyPzskHpZewE+XstHkS6+qsrkidf4vYRymQbjJO41VCn
OqInwY602GKz1gJ1qT6R46idZ1QyOg69yV9T8MIQC9u0acelBB6jrJxaoFSyMfGn
+wUjOe1ijC3q3nMhCcYw7CcLmilAlkm7mlWfruzBElQDekOKmsW+W+o10xmqaAX0
sjwYWupv96y6tBOWrEGjCYv43qL2T1QgmBqboygDjW3e6xUwuN5wrNER5bZcfvcC
xNiGmcqMbaSHm5KwRLVUaVpMs4pC9X42ldSeDsbYMyvC/CGl06SWUVMpYNnXguTn
b2VJKXQbHQLcBgrIeA7n0pUm9WeYP6IC6JODolJ9nHabksFiBYW6AJxor2zOeqSv
VGiMJWSdF4nzENrZbS9W+Tk6L5ASHxRZfv+Bn3jOUiSEsFWS3KRlNNg+TehCjOMm
SFSd0eiuSrnmmVmIxvxmSLEkGdxwm/Ne5AENmPcnCsedxdpQ5taBoDkPNg+HKmq8
Ga8DZBloU4YqohNJ3fkemTLlJDqnRHe30uhh9lCfmyhbK5t/H+aRyNoGn/p5z6TG
bmwj2QgjmwKRmUZIyuGK1QmTme8wylkZSRQRKcaum79Gg9OkNNQtU6+IncSedXId
zJIZIemBCXIh98Sj43Tybizphsg0OCy11Q6e6slxtpU0jA4SMtUImeuhn/B2ucyz
1e8blj+NiGjURcdwlGUb7DvLWfK2y7reYBEkS9Q9GHw/kWhedMc0vBu7ZO2ZvlRP
BOn80pR9W91zgbagaCIYOSQ1bhsV8c64JsPtwhpPCVeb5R90PROFIQHsl7CfGjFn
JF0ay7KUC5pbknTWWZ9GvRZyZaX6kFgsELdArse+g87xnexKIG5fL6CGpzoxVQve
0Yfvv6iTe9PBYIg4siueuv8PbQJjI5Vbudbh+cxifHjyXHlbluJRLCVzSWxDZLHn
NqkjJSLJYNH26X+2AdNyAH6BuaDboqcSbk/5AEcib10EbW+suXrCNfLx7qAGJLiF
RBieSALUzJlavkhRtjxsIN/q+F2GwGIluAbOuxCTs4OAmr2wVv6Y0/f4lqiFZ2aH
cMwD0LtX/RYBc2O5ncUcexR4YWV7KPcVbLulcuCnKDHWxjD4u5fp5EobnryoCp0b
GipVmFKyyEWcYnzT4kynEZ3L16kV8QI+AnT02E0Ru3kCUU6QeYk20cvYJIPKOJQi
z+5KFsB1rN3RHOf9tFoncEduNvsCt8dZs2TV/pPtVsYQSy+kBtZQkIVEoSIGMrFy
E/SAOoWPTqlDgIbisA3RydMWIo6GcWR+J5lUsS9or5JeiQuKxjLTc3hLPe7ySf9d
LXkR3KBG7MRXCSJlAnw/xBcS61Ws9LgSw23p0k/QCwaPsJBXFsggssojejB2M4Hb
G+D3DkUF+NN++U2IGxiKBgGMGBbJRcfmM2BsDHZFlXkkpptcym2ExT7DVlvaQXHU
m3w2CIBXF7JoLcwVOUX9C1c5AoEsNEWKXwQhE3sUrfxt0+Rgmn3YmWUItjkLzACj
3EfMBSgy85CR6pHP0rEqkF3S1unRzn7huZOjBHrQkQ33VklopN5XMg6MFD+WEtYf
YunDJUAVa9fu8LRJNzGpxZ3k+Oj+OfTh0bRvfGOo/r66YT84otqje2U/8r8cugIp
I2dNPTCLDZ/R1Q2h9fsOwtIMo4tGWHioPB15jgiPC0uBLPe7/ly4xxEJ2mk3BF6r
oECjcHUK/tiIRUw1thMq6BxmgGrfPdwQ5isIxoTW5UFZgucBtHjQlI3Pe6gCox6Y
k3+8OrbBiOwS865ZaOTRasjQdvSGzdVqq3qg46HXSz4fsbna7cOurK+hLLBDvNjy
2rA26aJS20B2LQPqSqlnjwkagehQPUICemCFh7l+NaWGITnUNXu6lpHaHeY1/AyB
I8UrBP6oc9r6mPz7CL5abilKuHxtLwwC/qXbXzk5ucbmPlKrg/Iw9i2i1u7unVRD
ys2mc1tkw7cnmJGexLibEu7JGZyl4Ee5RUcRwE5x03+KRWhhL0dWrVtMkEiDwLbW
aIEm95LTqEi6Gyyrj2j4rVuUu/0W0KVvYeyzWmvqNDdoQIa9z1OMVXr0taFPHhRL
QHM8cCS1Gq2xZubE/Zk6uIcCz5DFy2Lbz4e+2L1pYgqkkf5kewNa9l+ZULQg0b6O
HBlVeGcm9/AGasQiE6CPbda/yrzzCuVueiubXjwjqrBu9R9vBQeyX/gzhpR2D0my
YG8/PbWcudRc9m/POSipsE9S+zc+6IvfwmFJdpsblA8LTs+3eBpSc7owV1rndbJn
u2zkqx8XE9vDYj+y7JAlSskWtwONKtnRhWMW8XTXMLlH/kzaqcccYt32j74cs0Yl
k8/H/Y03j8T8wskYlBUrNiYBXYsP9TW8HiFKGIZv/tPhKFgElMZ88kbrNJwkXrpf
06wVnb+3a8JciuMeHQ9aQdbQWR/e6SSV1fTFy5AfOjUtS6bcHyl11cFc7McRrHqR
Z/MAHLJD1SXZizWisLMe0G01an8nKPmTI6wYlf4J0kAyzxtL0bCKniRyCrhVLxPD
QOCBbHyiomlTClPyCL/XlJtOkd+5CMWggpRPmzX+t5YWkk3LarAWabp0qUOlm+m0
WPjQCJfHSPuHOzs3SZvc0DfYJNiMTaLOcTd5UG+zRsDaTR9LLT3A6pSqvm55qC7A
A0qSHVcMgT2KMLop5eNyMfXza1cBEdM4NvVtg6mYZyhyrneO/Q3HaMzyfwHJWZvZ
6sXxZFn2jgPQS7Vzbejs9Zv69hqA0eh6QOGsc+AULwnPK8bEMPp7Byu4B6GyfS2h
mQPIQ9Xg6eLycn42K/F4UQminpcpC3N1EaaBRQSW4oV9MoacqjujcPi6S9O2JGvb
KRppqsq19glg5doWBGXTiY+7nv2gbZbWuU3Ohfj1NRNECz3RTl1wyu47WHXljdiQ
RRdaD9xFXKtHF1Pkq1J3WmCV35XnAZv0ZjCsh4eRlw2YatCVGf9wX98gOYEqKyfy
4U4gGhInn/MkeWRFjgC6EJ/79M2G2ct6Hb4Fk68wRWa3FrEz//kzE/Qfdq78R9O5
fGE1S0V+iRYvGY8SMUhpB9tCXUZ1m+El10cfP8OtrDOyCbLbCjETdmW3dVXWpsro
5mBaFSDvE3e+zXgQ3MbgMKWQguCfBDRbKCLqnpW8rTiBZ8Q20zTN/zqAQ7haQCRk
pc43Pm0CclKD3accq1KlF+ccVL13dTOUipEHC10MD7FFA3+UIjMnj4X3xTKz6L8p
Tm3nzuzIH8BYEpcQ0laJzuv6F9UxtsqG2w2nnbIniBiRzQvBKnJLy1Rvs/EFqGpX
ufgXwNN2sduny/WPQpm3/v+Wep9sD6OxaDY3H47oOLR6sZLc+Bj8Do4J/cxZvDrQ
S9b968A7Mk7nGwv0bKhoGMesG2kmgc6Ppu8cebUFgmI/Rjv2rnpgtjEmb7u8I1nk
faDk3ZrN96Wr0t1eAZH84De1RSOWMi/u9AUqF+47uJdZ7e4IwUGirAuNMSqHA61i
Fhn98VuKu8quD6hbrp1ci8ZLmFaQDvqLafOQ+s4ebT9IYbF1MSJwlxmYbh1bMlQ1
EOTWAxD8rv8j3DLUHXss5Q4C7+sqAVLVG9YgYanSrr0FSE94dXFG+qZPu3aJzqzk
jfvo7gUC7TBZYqIDulZwzjaKSN0xwkwC7Wvr/xUtg0PD0OZerNLkWa2MUlEbQAul
27d69zLVHO7DLWoS1EC+jKy4ac7Kj9pTnymWneQq74hXndmsK13TRsXLMJXLTydp
Q1i76aANb81HwPnbvNT00vA1cbAWo5Fmw1NmDz1pZtiVQEsFjRtIfaDB7G6pr2aR
MzF8J5RpX4WuB6gssHFYR/QHCQ2lneFgPbTXQBdDjNQGDvn9WY0tGaL+WiABcA2G
GqZe5wOEuJoYKh7EtamtQDCVrqZ/n2KmEEtDcBRf2WW3lRmJTsy+fa3//q2f1jOg
NaAuYG5Inn/k+8NPGHuugF8WAtJOeXMB8qjrwBpIjr3nw2tMEAYJ8sFfRSrKAUFx
q3wsKogi4m/LWSEG1KvfABAkqCdqBknZZwoqRWuXrGz/Fv809qXZmSIw+ZouAPkZ
HewURpQHMgbegGJxqiPM2sq2RCinIItU5nnwzsQUNsfTZLv83Eau5PvTamJ1OlR8
yy4xPS5X4GeanihDulSWhbMIrCUvBtX9t2yW4FKsGpSZVwF5K1CDT0GFYbapWxRi
9A05yKxex0ALOWcWVsmv3H+3iXS5DJygBF5vDW6pLwlyvHHvzQbjEyRDF8QT1ToC
CcIBvc6jV461M8Skj+6daIOgsZ2Qgb5xNV1OFv0zkI8OjoK1OwfefNZkOI4kW5co
IoA7oQqChFLONmBuRjTCFJk42V/gBElh0pRyz8qllz+gpTJVMSPJpPTk1AW0iYz6
H/iCp7lsSFwLKj+k8nSnbyQiU8iOKNDhu7/H2JGJeip17G3SWxT5vAKMHveEGaP0
TpWVG1gwku6SC9BpEvub0erLjjw5Twvchu4Bw/BusKcvNFp7DsxfQlp+5CRwmHVy
cj43ZNIL4mMOVW1ii+DMoWwpCDsvHjs6wV9ap/c93zI2k7r652h1fqrLivfZrory
Qe1f9Iv809zC2/ZGM0ihSPNcmrWPPIcXEUl5xbAt0tR8jXN4fZ7bxIfJcrzQZD+h
a51HKVkS4O434w2VM48lur5WbPQ3XXvupp1Tcg4fJPC0u5I72fr9yjOUOvdBUJil
1B1fIFeW4BIfH0qnx6N5PD8qVhv/1lTTqKVZGCzjTmO1xy8V6P8ZbgZVh6aTsKBf
tAJEEUkkwDE+FLxXq9Fh1+I2VzvTd9V+T0bJ96qnMgnjOCGdc0Abv00uThTnAsq/
rx6M3VwKAuRHfCAMnQdQDJdCZ+L9wFMh87X6tyQp450bsyCwPZeIJAXvAjmjOWGm
YIcQfp4c7Y5di0MX34M/5GN82cZpHnsFliBKGIFQ1U92bIGsnKKBmzb/I4ZZCm8C
nGYA11A27dUR1r0xaFbAMIegGOWqwlfxWeDaGkVgO7vgxkhN5dNRdEgRrRIhh2YJ
Fs/75t9Ub2rblI9fBaUbLHLrdtIPljHC0iRgXcfpCIu+sAUoxxyPcofvm8Zk1Eij
NKwOCfolQHr3asVBc7jhjHYiIgqo0aB2HCBbk2u3LNgPFAp/o3MgYdocUBVw3un4
Mahvc1CuSAwJC/l4FCUsG+RkAOZZJUGA6TRna9j6ELNLLWbMu8jg4biAyQlFqVK5
jnkai3LyoAomH+AsB+AiiRkZ3O+AhELYEiY+0sq/0ilSi+F5JXockw64QrPYh4hx
U0gAZPzd2p02I6ZcfY3t7F1y8sK4LiqLoq7y0vrH2P+w+iMW3WOIQbMQwBrz1RQh
RZKSGaiwhWMRc9sPuBOShBmBTLa0Og7pWFWaokhJkmTy18dyuBfAXLPWti7zNKQo
ge/UqqbSq/EPfoMSIf5HiapYyyPnA4BEbEyG7V1pFzu41FEpUwrHMtwu+K4tRfDY
jyS+t+Q99xjaHVNpYP/sEQ0Xnou80D4bmPfwrBprxdmzkuQRm4CiFC64zV4uUSly
XTdaR5a0jzjfYjMuBhlfP6+ghKH0uOL2XkRhqmcLFYEPOO/qhHIocUCJpzyMn/fk
FhZGuftefef5j5KVfpc5p7Gic/Bm0TRdL3LBMX5P+IgXJEME2CMTErSSZqP4hxZ3
uV38i8PaheY6W3GoRXHr056rVITO/NrQ3lRUHn5P6DSw81M+jOD+t3LMv0oEi0P3
NCI6Z/w8h6o2zToOZbXj73uVqZLX7Uuu+BtJIFxCodqcRjI09XI99J031n2gA2bp
ly92VDzakHOTH2NgImLuNxYbInmdxFFs0xJhFBk4THWWdJErlh7r+gwSBoRlpNTO
CNJtQDbvnV7HCYXaeobEbDwvldxWBt+ZbVDtIJkgJnBcremInX9VtnK08qsHEfKG
zevXJMUO88PPCUefVOunhHEGw3kf7kdPPdMKu5TrBCqESIs6iQtjOHNaRf42Ekou
T0qVuKKd5RJWVqy2NgjAMxBJU6fCZSyNQFi7toPY1xTzmTuIHG5RsQUfsLdNm/u/
yOIeghQmzSySKJmfa83hCZsey9L93emu9NIYYme6MB7wnQTAABAw8gANYbyFPt+X
Y0XLXJbHWxNPLyvTBAUMPfzAei92tQYpJsgBJqKgksmFcPlo67Qpp3BGt5but1V9
Xe2JcvwhHpgvQhyjFzYLHw3tXVmuLnuZod3N4I87wlPgc1a28sfiETZYPimzpy3w
69NBBORZutesxkDcK3qSvInCqCPgjXCzAU2ufBib/hCn6TrJWuJs47xVRhACziad
alcZVH1uo4Zahfl/BSzEzQ30tqhUQEU79HE2klZ+++kYZ/qyDP6YeeyJlkT+UasS
FocsX/J0WsCz/vUqNTQ7psKBn1HY6irYAatwXrUssyiYHlR9SzrUiYoYr1qT6C6b
941sUNzmVR9vUO7MK2dyY6eZs+Dk5x7T0EOVMS6Xw2i0oS5Z8Ptv4M51g+IZUHGx
+yCTeGcblTTV2nMLkYo2vFn17lADM7qO6iR/vvz+eWau4DxEmpG8hmhhgWrwOrTo
3buP7UoF2ZT35flp7J/5qRuZHGef1763gVq24/Ok2ub9V+ja/ai3ZGcumpxhFOQ7
rUv0XQSiK3inwz0VdgOHcaLyiikMDxF0GheF4OIovG4VHfzoO5mh84km2Gl9W6hd
ZdH/JpGzylRu32OUxE8xoQZiqRC5OacQwr+KwyuGzLh+dSDhh9YlU3ZDX+yotBCV
/pg9gp9VFKMKdK9g6++v2NWGRSw0lxyQfEVPQ3L12qkI+Ovi/ZMinMRCQHLucNW4
z+/FTc5/Mrm3Wb5bjyqPd9D6yLgLDhvN983FD31uiW9Upe1Ln6d+bIm3XzNwXJIb
SBqA/h90d3WuxBYSGzKY26cc5/MqXwHASxB47i8utRryOcUBcTJivzJWW/8Nj9GW
yI16avDRux9ZHYf7V/W+ke5hdKjsrEuEAwQSQzXcp6c7b5seNR6m8A5UIBmTvG58
mVuJoi+YL07rA7l1fCp06giO9IYEjAmGugMnkUToxTtVDmEMAU4VzfK1ri7YF38w
2Xjk/9P/BjrbENLa7mJ0xGTvHxVS9yArJfHjM50puAk9qDesxXVrwvZAVXI/j5vD
kgoe1A0qBsWtq9aKK7D1u3GUvFBMOHTAv7OZIWkA2HD6FuVH/ol3SjW/mhInThsg
gYjw8m1pBWYxduMBuPPLabPRk0sFgOyNypbQPOXDduAmysUgAoxqkVI21vb9HRbS
U3nbOFHO5el3uKHEH++rhvS6tza01kiu5b6H8kURMa+EhK+4JHXyWh9Od2JokX8A
UemuRpyh84Zme7NTpjm5M0Q4TCYto3asi37DAkmZOUjWCjNcD9qaKJpuXP4rk7Zv
t+C6w+Ss49j/uNCFw7HNxs6hKZvuBHhKvM/RHuA/KgXKoveRLlz8eMfhVR2Mu5yt
VjccozC9+UMFLM4gu3I46OJsH5/q11KmfrmCHcKIktzMCqv8c4dUCBaEcaq+fBb8
Y6QqVp6wkEwIlMFK0Y7R43PXMzO6NiAqYT1ylkqOUxPPxkAIfJj8bEGtXpBZHWJB
l0NJ/N8+vY1Wfrd1uRcjHk44CIHyfqjgODaDy3PB3BAx8ly51/Pm/RtkgRTXuSLO
DEL+bDhBybr5KOj6toUiz2oYRo4xxyTPWeibonyycAxhka2GijBLVMFFAbxKV2jk
JeoD+sXitX8mNjVqrZcHFpzRHbYCRM+BQ0ruQ5B/Vd3ehqKm9i+z2YfiKpF6rkxN
O29z1/gUKXUGS+gbTbwcMB0bQ9+SM8r3M89x9B8fvgLVjDHXwPc8NMPBm0bgzFVS
5n3lnjYMnE0Kr6wQEqPC7SPgCzL1hZUksTqlWv4f2XYH21mTo64Wtt8llg2mAFQk
e4g7rNlrnycBbbf1JhSp2RHsQ1d3FSw36Vm/jOAE72LETsQjWQVLczDn8Jl4XAxs
CgssfeZL6dNV4hl2+8zQXGsNej42AH8p2VYMj5dZZlNivkLaN22EpgoEDFHCKp4B
5KDXJcHUpcEOTf53TTe6a6eu5zHz/dbkg9RqoFQSSnEq6AQkMBcvPhaBFZTMa1uE
wsestxZE+onh+wTGkTENp9sk2Smw8JinCw5HKLSL8DHFEQJzo28OnYelA3Jtlnb6
MSz0DkTWfamyN9E786v5ruEbdnwAIX9hwph5HVS7T7Os/2prPcYnHPvluMkPsnu8
OPScaSldB0wL7Xjv4+kzwzBQHhbsi4RC/vHVQk+b+2xBJK21mDu2BeOkWRvBsx/K
s2kbYRsXgvl1Tek4L0PJXlc2J7d7iR//cStQMnTR/cRLloyCVn74KCtp7Wm8qJlx
Cr77Y+pbJ1moz8FX61RRNfzmJhHKwggVgIvCQslybQFPoERMQZ2pUv6wKqpE9kJN
BQHz8PB+mcKBPyoVNxoaI9BK7ehofh1HLfRs/pJABE0D+S7Hmgi+SIAMrBqpW/Ud
f5oiqHq98XuozgGPt8NQMbEkkzRvysU4V1U5NoUxYx7Ei1F5N7PDAiammPDtPiop
vbTm9vb6aUrxdOyBmzyb+Gq0CdpOCqy8ZMZahNI2KTgWA4+BVc5vj86M/QzWfD0f
3UQNh1GoxSlA4cMnuO9n5XBcp9gqYTBwtzl3ufT1rh2HpGYAccIcL10yzXPd/CTO
E0VzqzNiJUDKeuxNy7SqbmmvXLSGBWBVdgQNsbLb4AQ65H/deNqfRysxaYtRVTga
+dAXl4NiDwodjx+yCJZHJRliC5bPA6JAcgp6mQK2NQfsKkXUDekV0atZwIP363qd
nvjLtPYpp+S3opzAPVY0CkYRddoxzWKGVWOdEJuBGBGPP6fzEzbU+UxUBWQJEVkc
L2QaLcv1ruJeXRtoyaO/6MxtclR1jo8VbSYLW1QynQGHTkzykqdD2dFgNF366niG
IvK+hSYdXh1vpJIGgsnE7ANNHQYQHK5t9z5oAp9bfJe3BeGK6ecFUW+WqmpOs/Ub
rjM0+xXaooQWQgdc0VRsH5DT79/YwXw0yt91s3yK8T1eeNKgzPTMLjVlJ1/4ZGlv
GxR5dazPtdkWhMydqiVdPKG+BBVgjQEO1Uk0sF58ESLkB8MscAfGDzrVfZni5th5
AVIs6qy9m2p90DUu9HzzsrC/hBRa+DsehVbBAIjMfcmFceAHRWiptG9+F5ZFPttk
Ona3kpORxQLPi5XDuEkgnR2G27Fv21S8GBpA+ms0cv4EMnbLVPFvCMZ1t1QCIv82
noVTE4BJz347b+c4+vs4KCHPd85XueWd2Wx1nsbQTQFdM8JDaa/XYzdOnu7c2I2J
BVhiy15XkbtI2PLf5kserzewpWiNowM+Qx+1/GbIY7Yn+z3MCy0p0tbv9IIYI9ja
hjBPXq5zYOSZHkv9TfOlI/jeeP1DKbEnXirDoaukoYm84+JWopAo5mykM+vsXPgm
S3lsDrJAf1v0OK/v+itwWaR7iTrA22UXrYULom2TFKnLoE4xClRxS1mZ9xOnKATa
hIurPl8VerpBq1CGzdfS/CevxaZ27ZnK7qxMvrtec4j0VOPSXFLfrB1qw3xHhnxA
P+VbrJMbbN2Wc+ZjKbumhonjIXRqiEK79wo31s77qJ9K9GG6CdsiwTkPilpvfmfB
RT6fNYymmWlzf6RKinfwVjPgRIcMbDNZYukYrPBSsmy1Gu658HyhTJfrgIky7kq/
0Fw4gyA+hAWMqkTru3ghVCy7wJq74cJITZqlPG3ZW6dw3hp4UIIAfpZ3FtE5rrdI
5yrfqy4XaTiQWGqX0MmglTi8dXdTu8pdj9qm4RyNHZeuthPCkTQdTttuyPzTCvRK
wNZf/GgAbdt1NytmNZ28H3XdTxMtMqyNPKCrqGYH8knAeuGTIb7XNcHT9JKez3NU
4OTIBHbU5oMck2qcSCrPCf9jX7yK6dvj7YxX5Yv2ZQLAaERHFepRoEfPDbiPfneP
J7354TgLaRraCdxTaAxFXigxH3hauwtbD8c+2Z2Px5jXwUC99m3dmJ5oFIGUto6A
hvW/2V0MEpzhUOH5eKR9N9D5+4PkIS9ehRkQtqY6cuI9Q0KSnQPc4Jnqt45bZ6SG
N60Vt3QCveOCyqrV/JCtCXfGKfCvUTGmpEYf23kPftUF7jm0TK4c2MeFmKIDktvi
kP9+mOCfK21UzdwoLsSaRW5HsPfKWdlEpo2b9R2W77MEDu+RRKB8g9yzIeVd/EpG
Dj/Q2CfC8V7dB4jxy9uFSYkvbBJHEMRKUr+F6k0gEMj4DTwtYPop7Grw2PzypeTl
JbXyb44+ChALbD0KQSm87wwBYWJRncC8kd0+9aFwIsmRHUTWDy/fcagKK5aa9Mr5
vw4+6S+X9sBkS43pHKUgJGBYc4PLeDVqHCHNmiz9zqmpCTnNdg+WZjJkX+yt2Y4b
/kT2VeSVLSao1SLpDkB9VvpkuQmBHRvOwC+29wsVvSo9XtVWIzmqEE6dFbicRZ0g
ZJo97TW4zxr74EGnb9vPdsA3MCfQy5EfXebiIz9wcW+MPb+cYuGwKfcgNkAyYqlM
4Gm9IIEns0M5x0FWyOfuvES2dhH9b/KuzMHnW5ePgW9fw6Zg0JpR9WSlf+mWg6mM
arrW3Yx24wGMC4+70E6C4DAaALCjsQecr+ZqeWzXVKQRjs5EOIMH9tYPirOCSuDD
NihNBdaaNxWOGkhbtIUOcMfF59lC4MyZD8v+OZW3DdUaR3ZvlwByOLg+87ZI53Zg
Jw+kNzGKYSub8LvNnNU4WZeM0gv7CSSeHEOZS4kw285lTNsqyg0nxFlU2lrCcJa7
ebKSItKhiIbRAfUCircvk5nV9m4/G326QMuWKyqPp1P77SjM4RQIhM9lguT4b+z/
E4u12sIpfC6uSq/qTQ5ZGMzbvntjXzxss0qBsNhuDWPygu1UsWxDrO2WYhjwPGRU
j5aRxKU9sIDkW9byw4cOyxQf72NhGXE7SUvpr8Hwp2kTBoRRQDBoUQa/03TOJ3hk
WTt2uaJ6TCFDHgnfp0Rc9ikhOYkIweciq+xyqUk+i5kXSnTf4B+vDbX54UwP1InC
el56yiz9KzTUnt7klIx7gYydRkViYceMMk61nUWzdt5wjR8sFKq7TZjhO5sGsiE+
Xo190rjktg0tnNCf0JZgcMgezIIAWBlrDZLETE9Yl3vXlPkh1QJS5lGhsfUYrv0M
dGBFiHhwLX8VQSSEilLq9au67xNBn4dH+auj9WCaDXnbGUIoyZh9HAESC2+/cQIO
F0iMEuw6LiDTZTkyzngZtGmHINXHAndGiP3kmYJ45ek+pbNENjBkk/oygO0A/1pn
zsv3xWinCtJkut78DH9QSdYgLLR5Jv4SQBJx+ptB6rNqSO2Q8SZ2DNkHW7dGzAss
caJd02pH4sGorGU0af1/jSDC1/jjSYn02Ib9lK+yiN3YbLi8ExhMAkQYlfTCKGkg
0zCBet78zrdMNKd334eLCpSy5FwpRYeLyoBZLtvn4bjjumehpXyIcScSW9lAv/XH
qVPNydEyJZWgYMTy7Y4GA9H97p2cGIOPANfu+GJ3pPYJ1CJtChwAAVIJ+fvAdX6g
Q0BzSXAsDctFCYeifJMuO5BRSqSJbiWnwwUI57F41s0BGKyWaPcOyxKM2bFkc/Cv
vbQ4iti7oR83XOmWakApylnaNbrkOMWUmmJv85Nb/Z/NSlOfGxx07iHHh3QdTXJK
kibBA4BReWE8mr4ArK/jzETSUHnf5vjqa1Q/xqSVU0QeougnEPv+O+r8Z0/gyjth
fkyH5+XcbCzQgUHu7zn9ZGMMJ4AqfZ5BLVDcHDAew1+LD1FdAeG5begaYfiU1Nmv
gcl7/csMVs+wXBsJ+O6Kicagvjp92xURk+VtahxLd/hBH371OMXLI1D5f+JmuyMw
YeiXb9I1NASnJgb1enTzIg8poYuAAPEz1mtsFekFuB9eUncN7XuoiAiOF6UK6Lxl
2NFt121OYYYlS1q+9pzWpLrXlhfmt0fw6hRQJYXBnEmO5EKntpyQyd8ajON5zImA
fbm65qSDwvs/n/KR/GWxzNRvM5TldMP5U0MgXF2p0ZeuDlMJa7nZUJDbYS96gFz7
D5ATRGeOcIEkeODWECNmWhXQPvMGTgUkAbFfbOp5UBdHE1AHsl0A2B++hRQvJsBN
VJ0mRehMiYcDp/lfZgO3tU4aPBBpevS0e0vSeK2gHVxxA7KkvME8lEaFQkcsc+Ol
C3uYUVTQteox4vYhj40FN9cAv12PG5Lq65BazqZBmE0fVUlOx7rSnTrbGx/ERHa7
zp4UTQrG/1iwDgPGbyDqVA0PlIFyYUfDy+p8ECK36AoQmHUCFCChj1NmK04FFiS8
PZcRObc7WReAmSOYDvNbL57mpMj+5PPtxk74eF/ZNX6AOdnmZ2DNFUdpEXzorqzV
fN4jcYa25cREHoVX6bzQncSx1AlSxw+MPM8tXFrIx4c71P/KB7Pw1POygetywvQn
e9atOUI5plLNnJ4WI1aVq31o7aRVktB5UIggnuoKLcPP2wcMWdRRHid4ORkS7tUH
uMOn2zaO3SKR0BkNxPJjtY6FibbOIrvr4YFN7BBeD2LKog6GPu19Gf0GM99Cryff
wmG9mkuPRT9WrkjahBg+6HaFpdsrec8bhVCMFLsDvymxE8otNACa8dS4g0p9yKQP
UoajFW0rIs6vmrgA0ADItvCChjl7B1duXwYfZcNdT4fBVTgu5BzdjdsqfbNLuDrj
kZ9eaehUq7H0Cg6nhDhUxrTSTQy2XEcE15reUM7az5OQvWf4a+TKTfv0wq3sW7GR
Bq7rHzBzSuNGExrII5PWjZTIHZF8b9Teebp37QYpQeZhHB40QuVOtcSTSetrc9M+
PmcYF/rhP4JzaVqd8Jtn8LsdCj/DJgaRXfKVi91GTXhdK4rLpdyzxQktwrJ7dK0P
yipokxndeOYvuba+TI7m7yBdMS0ApGhV2/UTOuwfp7RdRn+ybOktwohN4QyP0ol2
6aeHv47isyiH1deOxXayxl/ketz0QmHvMjeBZLIYSO6M4bPDTs+Kn0UZQ+rnNRkG
Dpl5wjgfflfgDAFsAinnlYRfVmSVLyDn1XfXMMVSedcV8MNrrw1Ont7tOSTktqB9
n88RV8dHILeV1vVkS7n6dkx5+CFuasXqhgrqxGYR+HgRY/ryrUovuXt/VryZrVGo
xn96SArohvW9++ydh0PYyHCJXikJ7Uu6fEfp3wBn8uvmAGRuznWmIxvzSzX0AEIa
HaHUHoNNpePh1FdNJnCUSDCbWuFdIKxekODJyvzBsq1HQXW2bLCPPXHgBrARNIjF
N9UAlhu57+K824D0vVnUybDVUB3x2tbgqPiz+w6ezztjpW7Nk78LdrHU+P4kIToj
qkQDpxoSb60yf3s7w7K3ftx+CmBhe8GKoQVTtQkePdX4nFHL6lXrFgjGx/TEc+GU
dYWyh38Iy/x0lJkBnUbSz1fyIk1bqRxJSPRsDFHzirAULnDmwJlIdT/oVY/MR2R/
NHJOU3YFFmHIcSp2aasr6cY4l4itelYJVhSsZYCnxFYkAc5bZwgt6miIfKM/xwGD
VhN+Axz+/rWGvy1CdG3AqGA0gbxK+QvsoJ2gM6uphdzALT/kegDIhW+UIncQRjNg
QeiSbBTBn6j34h3bHaq+NhGCBzel6aoICcT+2SuphkEOGtktIPosgab0xS+uzH2W
fG6UulSgXt9eO/JmIIdnLhqhi3j40idi5goD4ZNp5SncoostLKotL4flciRjInaE
K2p6o/BgkU5f2RTNLPtTbKwWzE9l6rFhE30gfJ87VoswQvOZNBsfIHbw/klp45Ue
SAr4x+wpXY84/i3SpntK2ZNqVS7FZ3O1XwM0lwK36t5CZoHi7xTXckCKZla3zq2h
pI1M9/MjTZm3kCeOygkq3Tex8LzBY+FYT8YM4HtlNrbIrts52bQ4slmmhWj6jQlw
A189Llh6OhrFcUfcuVIFkzWKAyhnYQ4aIpqhxSIwoWL+J4qjIwtSbqK8T0Kh6v1N
D/UJ642bo8uFBuXwlxA1j7qaJq+cqhYH5D2EZDop5XBcRRycxr8xFxM7WqgKQ2vL
ZAJe3JMBReklbifJQIAARkCcSLYPtULFw0RwqsTt3ddrZ8UBI7pktXNxYf5c/DlL
f/RVlkwkpca4ENBPNRolDBlMoFuwPm8WDfBfTK9+s/N46o9sx1Y9mZMw8dHpSWM/
ThL6Aej+MlzOSY5ftoLiXg0diFhbxTbP68ulZfWy/rbEE8e9CKuWkvo5GtFK/7iM
Swl/DNJYNnNA3gKhkrFf0ODFtt8QlrixApblLgUdvs1P1YXh/fXB1kSvrea06sqe
BoAE1p6xZSB5dVHBlVUA2ITyYoAjVxqBqIfQAwQ4I4KKP8frHlTzP6J+RSa9hMNn
QbxiShBGipDflUTe26I6L/QAUx+bcvpgKmftqmhEk3d8TYlfTZQnueX1eijPoAEQ
Ouw0zGwI/MdTPQpSTaCbIvuaDKLeMTRkn5nqv/pF9ZybFTZKd0ZgeGfLTVLw61wP
XRXiPdUoD1m0WImYzkXWZkiqZnqPv6Ul2frflcSN8LiJVYL1osmeepxT81ouWz8y
GVH0PRtMXxVvCPXR7dDslX+951+lCJ0okkg1U03hcwD/R5cMuqBFnC02b3TuZCLg
awzi23thzVTaUzCTuhh3NmdhyPZBwNJ1pONFgYUgzi7FOKkBwTelaPD5Jz6xZ7KW
dOsIX6bAFpRPRuBWumhxG07ZJaSJ/Ja6IAdgwoMmhZHnULSvUivnDo6WqIfjck4e
wnQivGcV1wtfKqyD9PMYlD2+Fa3URrLNluziCRTmPKWVC0sADBqd7pJB1Ehbr8wR
Vn4en7S9hrSXae8tgu0AVA7JTe0Vll1qn61XX5WjJLxhlUL1Ck4Xpz7IKceRjsNU
fpttWNlQKk04SyR/sAQOeCZQHhYyVLbVbxrbYRPzRtAEeJ6OhS77EZFrnB+SWlYs
UF1c+fee7nF4b2+5C6UkqC2nv7xeTWBEkkZ3Tmy608wb3bj4W4kR235Ja2N5VJzg
vNyD7D37kqt4AETL66ff2sw7UFHonQtjatizYdEbdCuyNWGwTTF7z1xYM5jAJJfK
kznOe8jjWfT9pScpvP3ovmMDY+baKWeOa/JxJULMizhUXTDhwDIDhRH0xwZh3dwF
2hnsk7iDoce/EnAzMjL7XUWASTbtTnlgDTiuuguyZaaZA0lV/KR7nu9xqtCM9/Wr
NN5FmJ6cwSaUwOv+oj9LlqTy7C9HCzjBPVMWJa/NdZ2bceI3w1A5UATDzKB0+bve
Iq1/WKsXZMgTINyaa+9GgfvVOPPSdkdwW5WJ8/AlcGFUo/bzRFY5OnIRDZ3kn5P4
9kChJfolSA+vtZF6xPTDicWcwgeVXEVl4EH7e1Bhb0VjCmhmfYmE5o6OkRV7BXzp
Xd+nUcBKwHYfsFhoF5hAeNTh52W1jkawU++vBliqHaZ3i59mXJBD8iKOgwrcWZ6Q
8Bt6q1sxqjDp9Y4V3v/0CJiiCYSdnqQSsZz60nXkZczVXpPc/szQHjaXcbJJNahx
Ki0WLMU5Xbzpus3ut6rPz0vqAVrQ+Z5xDUwPAgJyE+5ajmlxlDP01ULsUUFA8ELz
TWhLjVdzVYQI7jthNqSk0nkcRi6O/ClPcqqH9eFqp54VOAo/Vq/LveA3/aSLI5Us
Ncp8JCqktqUfFlA+eyHTQPq53lgfoTqd1x6D9j5FRtY38WLWta0AVYl7g9Zz5E5T
9XBl/3WUET77m/NgLy6mgAO9GKxhSKMM6AczHXL9HdnrIgmo9pjVLSdt/Pt/RCX0
hOeYjimIFYPl/ZSTOXoEeIgZzPLKRUyLYotsC720N3ZObAZ7VByhH0DU9YILp1zL
fd5ohNGU0XtXsVn20cWZw9k4h1weZpqydCyCDHafD20uiyh/JS0ZlXL0w9VlTJEr
+T4Jj9LVzvfs9FSfrFJLjqXNU/OeHGlnnntmGvg5w5Yoo0S3w/POlUqupp0h2beC
RKXkW43pkXX+y59OU+oUyjBzhULGArr8Q0m4arOaxjUuiudfCYXeuyAwRylY0adu
Xcf6oqeIZwutrLb9CE5FNKrtVPsVRmVVeggb+uhBE+f+Zf29E6mKcKh+5iqicyC2
4JLBywT0IuHpw7SKyE4sK7dggOgywwefOFSPSi8V+QauQeqbnP/yhGAuOKU0IG+7
NempAMTvFNycBlZ8oEbpakZBHq0wCD2DbyOSB4jKqtu9udtTRicgGsWhac9qalMV
E4OnFOIv/JhZyoIOK7qo7pYM8m4mkvX7B6nqILOxudgIG/7iHej9wf7/4Lx0quNw
b4n+4qIzePBkZRpfnufg/FNvvek4jArDWvXYSbvWcXVPvZwofidLUN9dZgTvM3eu
UNtObkdKTsmNwCS0j6+K3Rff8aV6bBuCIwa84HQZ6nEgD3Cm2IZtNz0nv8+Vtueo
Lh5uwwnzf3wepFADQ7iN0Xx2RsDEyGI1Y302FjqoqN+mV8g82W/b4g0JDpCT+SA8
em4K75NC9PUhOjM61gF2dOG+KCEKRHXPYtoK/E69pXAvS4QZAWmwnKrxOseAPsSL
jqWA8CN/n2mKgoWGS3iUqZQnG0M17ztFmqX7Fuak7W/cUEfCW+nKT6qXhVLWZgbE
MzvMP4vsywyU7Tqx2Yx+CG5aX3fCdbxNBbUY4HFduqKLc5+5G3FYTYCN5/lNlU6X
2Ctlsv3SGJ5Mia1tLa+Sjyx5NIEGz+JA/X7EmBgoqIjCS51eqx7EUh3qGQvSUUBX
vYLbMz+tuFnTGJrTo4M1k3kAuNPcxZSBAfZa979WWykv1d2+vxkYFqnCRo2x8juO
9cXJXhRJ++WolMG3tMAd6rLqzUy9AZ5O0ntkU69ieDxxYUqoASZ6H92YII77RZVd
Dzm7pPFWmRUhltmzJJbT9CNfyDoPkxdtIoYH283LROQf+eCXiBo+NnInevU75oTy
iW/IRdMFSzrIPC2tVd+4ifz9lb6xeSZMVjCYIv71N4pqZrXSW0h1AmAxKngPoFzo
Y7lFr5YtVSOBaSzZmM6nGrFglhprN9RFT9FfRb+bkyciRi8XphGQN+LpmcEfHfe8
UfUftjZGeuMYXaUxjsBPC9+evlaLlK8WWXIObzzwkhUant9qC7c0S4GQcliAC8Fq
fn3L1w70A9nCL9aq4RJK7n+XA8KCHZwUmPAamO3apK140J2bBvrCpvs/sbnM4hMC
p7763KOLXDoX7qAv4MX+G+VyW+KgBbtNA8FA0aEyFJgNG0ndrwR3u9eOrNpnXn6p
0LCQlaNQmBDTt2ebhDSdKD/Of32HhJbxrRcW6XUtiUabWLO7SUWv/y0LHQrSMSS4
6cbaA3NIvY/l8tBkl2pU0Ybp68XT0/fueTSJ3fTxAZPqfFeqQiIN4caGauEANkme
QIhN3E4H2BJuuyaG2LReWLJYCH2afFOUmpJfrKO4RhnWSRumadm7II+xi4AY0jTr
sHYiRhtoAu5LZ7QIBqWivc447H4l5Sf5c9GSZD+BsqQB22gNCUFgwD//JmsZHMWc
DEiwBcVm1UaB8OoeYr/c1i6ua09cZW4naJfMSkOWrgsYsnY14uCj8Mx6qIPOqt7F
0HclPF9rpSboJivOlnyW9k5GucRfQA5sxQ2ORC/ehsI2jbpF6T2DiPAcOmjsGuGX
Q1LJ3VviHCUF6vx4SL2o4F/YgtWLrtOxDOsPwKyjLtc4F3w7xPTTeCr4yZYZqIFs
N9So2eL4dWNEqSEFJqYWcDMDepB6Y+dscVSKMQlpmby2WWbLBwChPvsbul4cgL/L
5A5DTAAA/yenYYSCRpV1XtuQgV4tRCw+UcYSdtsyjScJoOHE2o4wFx5bwS1QrWLG
KVjSkXTMnLBZ19V4AgJM/R2c3MgMcfBp/U15G5o71WBgQsYpIPXL9X1OJkWZjdLB
+aWGRkkJySAwLbt+CC0fkc0E2H4vfd0mlSldkglXZdWLL03fGPKd78qy0nI4NDfj
d4kZKcdp1pRmZ9QJl2xnU7bm8FXuvPzVYySZ8jviu73PW0z6wpfk+UzrO5R+0Qa4
sBrv05byc51kwwKwPLGxflbLoB4/Wrj1JK1+MHn8RoMAImLx2jH78QmBZ+xo5dcy
2LRIlKj3BpOnsDkKKSkeOnOayj58SsqIjtFzJP8BjO6sw/MYJTzTGKOfcbhDqPyk
n+o7BBSv5C9pC7UFHg1pRCYvUSOrvH+MktqtJQjQFZz1u5zMD2tju1GUS4NeVUlV
1Psxcn1tw0PdEBRDsyKDjFkB4zaYBBmFZMGJ/+SjnQNe6r6clReaHTCyKDtG9vuP
ij+R3sjdzvcss3L34dJizuNIfC/ZjDjlirqWLcSMWCy+TnddylRxi+Mg4QMkhd+Y
kZStkhdVIAPUufMUrtQQ4N3io1peWBbYtjnGoTsZbatcUFcJHaT969Xug+EqfFEu
l/cbgeWUVTsxUbyKvYosPueSBcGOeBJrEAht6fxf9oQrgz4FGvAhfUAC8r23fxar
70Qgyga9yjCKQl3hk2/DXNTZMbUl5wlpki/4+z9bsSLiX5wXHGbYmH5dv2PvY4qd
Z1Asr47oLqbzAh/Cu2FDROegBLaoLnSh/JACrYyq7NZb/qyIFXEln8UBBSIuHU9Z
QHJbLVXJ67AzcJZSY3dErshSsIpJTOUniBVnVFCpojq5GCsmEQtMo1AVIDNEDUfa
Wbzaql4OAL5S4hS1kGNavzZo8sx7j+2lm2oYLNjsSPfMmpnghxS7W2SDgW92A6Un
b2bb4m26XSgFr3ZaX0HpXUZi31ksze6MwPXp4293GqGLbVmpi98eNZvfqRJ/CCSZ
pdo6HYwaP9KAbvj4SizogYg3JV0u9yfp/RA9OPRx7I9tU+/Zfa2wrSoOP9g0Hf5k
blUi007BvNb5AajXqtsPe/FZl+6xQe7AqVH2LHCPsD3NTdpHVpdrOFrqZH5RyQEi
ehx88qQVZu4CJyATGFMsnuRPjOTShUbHNKq3SWXByrZmOKpMWZoJMCcD9QoVriCJ
WuM2UxK4qFEIISiE/7bHu2vETgyQzGAU9pqVhMxGrUR8TPtW1Amorqd1zfpLXXEm
9I86QVNMtyuiYcLOFFPmsx61qT6NmVARju3srWMlSQXvPNhEUsQhzhmWigLmn0w+
d4pcyC9J2PkhC4ihbSWmVPC/AMsFvDq3FZw8Sdd9Dc16sh6QO3JL/iMl7+ArBufB
zNUAjreG14vxojrLYJYDeGjUQaLhSwwGnFOn1PWD1x3Qiwr+0RD70NJ6M4YDnJNs
XcX2z+o5kOgZazu2ujL9xub8bdzyWU6NayC07z3byiFr2T0ud673/PZ8bPN8Nwlx
6+6PjUSgJWBo2JZPRA/ONldvYh23z9O1p1H98T9OU2Hrt3UvgLgjEEY6jJXFV02g
fmQJCiDNs6lKHBcgjeyZH1V4YkU4zqsrq+EO/0M3OidrDZcJ6qJ5FDdEWhRwzEHG
etfuRCFjOdmTMHcnjF5Pu3SKF9Qcbq7j0Qx1JtgKMyOhSJGzXAFDDwVZpNefxmY+
MU3tms+DW660SQ4JEhQDq8mukXgATvPPC+64vpBk0BBMlgxsUX0WI7Y1ENM/wEw6
ZCM5ee/cs8TdzFxG0Ia9ve988QujLmdqZN3re30F9VIv/OO7krv+SI1vT1eCHci3
+sucqpAoEOIQ632HnOCkNZmgTwI8YUQ/Q+iO8kz/eXX2AJvI2VvYZFdaMAKKl9hN
IVmkWmhJnoQm0XVu8N9aMolWkIZPkRCvBrzboHT4OZSA6smo0HWHvuQLrc1j4xhT
9fq+2GArosM8zGo1dITmTNlK2Ugc2E+xV02NS6nPHiYrxanY1Jd0S56Sf+tXn+QI
Q1OQ69qeXSumZXOPNOgOJRHgxEOPfxhs6ahs53vrL3yW+dxB+svVdN7W9FbzkHMv
iiuZfQRpRlp2eBgSlAP4wx+hd9ySsmoNgbIHz4Vt29Ve6U41q30J41Y292CBnUX5
xgDbSPsAfJhNHZm2E/4AsymyMHJjIbt+27sGgw0uMRen4mF+DPgi1EKLRwlp9uj2
XnyrijNNdYxNF4oz6/J6dTJgu+Vm6m+a09oGbgOv6IanPlWKCyjJpk1JtPoPSdXS
C7ZVJc6529m+jlsqmJYRmOAI/qHYhBrNcbQlRQtKUvWI0IzS9PtwVKEIkZ+E0AkY
OrEbKa9cLm7djEZfjyMiUqyqtNlomaFaV9N13pOp3wbWKod8tXYaqI/+q50cdqyD
ljWflRZq+S4YsK2BgiVfuyXkLC6+WWUCNMX7eyyCA12lSiQu7U53mJyFckZAnAbR
5NrUdLJ9v5dWnwocdWUTyOH/ZduAFNAgIEbBIsWBSuAGHu4UmwgTpax47uOlkZ1N
gYtilclXa2KJMkHm9/0pABrK//yRRMXqHeAJtlOPC3PGRatSb5hEHzG1VKOk3hbz
lrLPKhfs6XcThsd7PMmHdS9QKYN8PirQ9kZWF+U+jjrPBUVM7g6kkTvDHgN/gWoP
5vIrr1Zd1xTx+c902wRO3Ff8UxWddUQehWMkrfQJRTLclT7j/2UovX7LhEnmQ1eS
4ZtNilHrYyzP+9VKzq4cIncYZ0pp17TjE7valRPzrvkOpeNy/ZQkJIJXjLYx3mSG
0mtRtIINRTcAFbh5BaXn2JwK2WFZ1zPn1jVEFC+6vdFn9dN9Lo5gbQwHWy5i5VuY
nLukA67y3keTZDaLEdr6tlhAPfTnY+By9uR9D0gmT138/fCaJV/S8jOP8jgvLfnA
s2P+YhTyy/9smPoskmklm5V6Z9y0DvPpBuzaS0j0XlY6Amv1mo565dq78YQ8CgOk
atF+6UsULudikiksFpXBct0qcuxqav8KwR56nLiY8nPLH1SipPRjofdbt/TBitW4
snnF270rRocXLMQJefZy57dd6wKUfAxo8hTFULCzwLEpOSIoHHX5KiWbzV0RuxPE
2FwQhUoNsif2AQLE3mBxx55Yqg0LHiWbW5CbAi+UQ/d82gHkfLNBdTpGrHE6MIMa
GNyhyx89ubH+VhfOUJ7bI8twt7XNSn8PXPldj6KMTr9kKh4zovQxJwoGFlNMnASA
K4vY2coguW21qS15LEZql8xHlqaAA7UbcTMgCsfXwVkp4dRf9ozrK8q2+mJ0kQyU
sGI4WBSfDVFhMduVoJPcI462JrBrevFWXwPVT050LksoC4gUMJo78VRtqTMfoxZA
tqC8uAGbsO07GHs4/h5zRNtiCsSMdTvNitel2Q5IhUhvgVhvtf+S79xRCSdEOO2v
4GyaFA39g0p9R7BXsyvfePxbTQX+G9A/FEOOa8Mc8zwuxjBSUe0+IdUKPLB8kwV0
erZm3qXJBw1R4Rxfdc/LP73GJ04ZzR0CIhSNP0m1WKD0R/abbXoXClxmsnBIPPCy
alpln8F5KejucDFz50gDJklwuYkELwNzVaud5BGzTrF0UElqJM4gmJm27cUJDB5p
Gk9akX0ZPst9lsEVzk4fdR7jwD/Qw8Zx/0DbhzHve/8MZ0cVmZ1ukbl/7f/HVZzM
5OmAMvIhvV5FWb8aGQ6+e46BT7WHDfgjPSzlZi4QOrdSyECVhwvzujFH3gpvd50L
hTCJOvl0RtWToz/A9JkUIsDYKnh3i+0pIkAHxAsfasCGVZ2yZFf2gifL+FW3XuSS
1R3iRdsaF8zW37Z+JOfM1MQKQ9T3Tm+P10T8caFsbA0h0xAPsa1lllPKeqV1A1go
Vk3eQQg59jDpNi/fxsy6HDsKtdTyRHAUS5TfucCRwFl2Ca4pE2xN8pUcG+BJGGve
EBwGARi7+OU0nQKXCfI0OeCTSWW4FZZ00/NAUN6YRroW7fJKLDlV59nih01NaubT
JzqgKDSeqHsnY6QvLfHJR0M5Bxq+vM53QrrgYT4YNS+tSQjvzUuwzLciUWFW4HgV
3rw3yPZvU0dvHtjQJrnYgz6zwo86VyAy97cgxQ3kpK8ngvYB2+bUanHVuNfmPuRt
Bm9yAdch7kSVOoT9XuGMx4Qgtbz7z1RFpXH/0D3oCK6XuesfYJQXOnN6Xw1f2D7t
ZGu2UjroD2jV76cL+AYoCyJx/UmVMl37xSgnI3RN0Qx04tNKNTqOuf+gQydjsJrG
77GuUnK3UoptwblbVZF9L/WEk7sx8hPga2Qmci4GQY2uWT1IgUxLMPbDaGKDK7AN
5MEz2SpG1conGM32zOxgqi+y+fvsTgLdStXstqtxWLVa2rD1Tokt05FwBaDT8ZQr
fVCeu3EFaJJL0nuhihriv1n1T8S3Qujigf5ELE1/TI8h5I/5+aZMsGp0LSP8gVps
xO2VUDPiTXqJEwpZZVK3X/ycAr1TemoQgDVTzXCpYbj9ZozKlYtABUXxUGFpi6c/
UTGOr/BJfHQuETlJ4chflCkTScCoshwQG0uiH8G4eWJvuS0Qot+aSmKiJnfmgatq
v8hUDkR69iFOGYb37t40DhclVJzsOkMcsOb9ckeYctogM4O1uQklEh4kqPxG8FDh
9UXNhQXbH7jOQeWOsQiMq45/YbLI2cv3P4YXmRgKhupDGCvSy45XAtyTyfbW/kF/
/Z04PZdYR3kXAD13+VaQtstgUMjN6Dk6kvUKq8kTR3YuZtvH1/51sx6pwdwCjcGx
H5GKHPcbrr+HW49MY2ZNZ4F4X80zpEznQ2pJyW8sGLNcpqcV5DTxAuSekOtTlBzT
YkOE6+XWvq0r5PdQai7kVIEgbIoZG22Xot7nzVNQScl7H/fHyvGmYQWGsLYTvXmr
SgKMnmV7QPDt9f2pDZ8VgCRhwgVr3d/E2baNNuZgW4XjHbtZfqo4sTRJn/Eayz4N
l5+1raUNCG599lxiAu+Akmn+UIb2dkdHA8ejYFPFYbUk83JGES1Ra2rmS8JhMi6j
CY9BeFsR9Zh5SFP+ggeoIk8VXv9WCxf2Lgxav8D2L7I28IhkVPKG3fOrxG4ip8mM
IOSgYvs4/FA6p2qgeohvMy9/P5k4IC37sviQYAgauRanmC0up1YRradP9TWUeipw
LIaz5dM9LWAoFLTgkNCmibd9Cn227gnL2GMEjFlxLmxU/9N1aYMv2P3hAXjQwxgK
P155DzttOFZ3ERnEpwAGZ+HnRtOpegIpgAeUIrBr9ouCX+UQaTaspRf7Jy3gbzIl
R3HNBZkaEiBzKZq0ZhpXABzGKuBMdsLpnfSUiA+MQZWWg1ty08an/q8sxBi5bfw0
DPuQ9fqNUmmHGdkgJ95oYUjUAXjI+E1n5wfDR0ZR5mE2s2/algQ9h9sStvZTsEZW
gy4k9AoI/xwZ9RFuXrV0/X5A1yOGSU0/LC3RZwvtFouVYQzesuzQdKR5NaSVjuio
Uuzq9GQaUqTMBDcIV4U6x11fAYDg0WcHaRPgBzW4Owl7LNqTgEFg0tCpSRdNp4ZI
x3pOOOIPqRufD33ewDqbhBAPwD1/h/HVCp6XT6qx6TwNEaE2CMfBHK23QCK6bMSg
JTCCQB9kzBK7y9ZycFFlxkdMejBkF4feUOaFaPXIYiUWNnL2kAFYvaigv2frGXYz
DmZGjSP9Z4OJI5cCqxvpvBNw9AawhQrmOdyN5kkI4ahq4vjVlY9W9ystlqP00OXu
m5AoT2AnDM3C4ED0IWMVSgYQ9xnYBd/TAypFBc6YZGwkYk1eH5xypEM2CHXoICij
SDFMI7RRfJ8fWTDwHVnDmFoE7vKE5D2ZSGOJQS2P90oARE7yC+bY11AyfmlOtfYL
Uo0S2LCvgY4AofyYnPu6w9KXcXKqjoJ1mNUPGHmUfOEXadplc/x0e6BpzQdcQLCX
UhbPaWgm15YEEnOtkVGCK5itCjv1NL8xD7tXUjEv3ZKm0zNrhM3bnq1a+nR4fqNi
XQWUUtohLyFSeXtGnFU+O//ner8LnqHE0nk3MJBIvK/XFftuu3OcICESo0u6nZLC
VDbDuFPI6pF2R8EavB+7jgl6HwcCS5eaVn5YjDy8Dwn1CDUN65npimIdrrD+9nfX
mBWjn1LqWKn4a8NfXpPtr6+j759wG0vm8MPsC2FoR0Bvi5WlHmEETucGIeIzPIZd
FD+bXvmYFw0j/SKDegxI3sM/ckpLTo/wSzABPhDZbdmBrzxHA9mfJk/1QDSOYT+I
REqB6YzHz9yqvOS2wW30U2ON4cVlh/VcP2isALCQLxY+SfLvIRHmkj3nQ/otF+oZ
lb2qsN5KEyOmp+JnjZrFtTAfCiV/qcagJuNcMymotRNfVAF6LqyhBWybYnD1S82b
STnI9rFZsrWpcm52Qf2l5uPKNBHVzGuXvZvwXCPYRrbh5nuXPxSRpI5ARAB3AxIV
I8VyI7QYzrN3IMx3bahL0CTG8INBTf8iyrUmrAJ+YuRgwT2cfu1F9HSjbRhJKmL3
QwudELnjTbS2iniI2DxmN5z0dByzHt9vbfCpNSS3Tk7B9i0YkFAEGKTdNGauKIpm
rqaJvh+XIfLpICDMLtwwQYHayG1wpj9HnSTbZQQ8WEYmxBeTeorQHluDa/NWrOgU
G7cw7NjVx7WBxZrYZIF7iqPBo0oqVYmLmMjusUhL9DdaVPiDwuUgB8qeYxW4flco
c4VZkafxlFbvYRM6ZP2VonypH5ac+xCANy6aAoeC+JfWQTj3GuphyTSKJAW83gb6
K69aP0FodgYMerQLfv7/p07na4ILyeuW9GmPXNYCWmjMjh9rKnvXl3cwnXhqOZVk
pWrtU2sJt09A4PYLQSBrxM93QX2R1Omq10h6IpDCwnfpDhmwZeU++iTx8Li6I5rq
hWncflN6HuPHVZOQkQ7MAhJmeskKyJP9Pwi8WWHHyOq8DBaFQ+iCHs8UDqlDVYtT
GPLkJT4vMmQM+0XhxEJY31lhXI86T+6XSZ6VFah6zhZNnw8BYr1hDRpwzgyD/Mhi
NOB4DR3S1YKSjW7vjH6sYg2uUMskzSoRaiA2jyNZoJbxuIfTgg9ua9uHZ0NJdLcB
zPFJ32XO4GjFDKtZl09ZVvlSrkYPAzu+ioW4TDDRpuCqsT1gXIn4+F9Q+SOhuzaa
9CkEf7oyE0AYlH4DNiMqFRdoyeUINrcVqWc8rHnNdl0M9nD2SS59mqbQ1rXgHCII
0dUb8OWwMcy5Sox4z6o58L/kywbsdpwwUmSVu2fu7B4Z1A+KyTKdf+Xarkb52XHH
04TyjmMUPp20CAzmO1RikT8HtM4zW7Pj57equ6tf+M6UNwBIvaPm2LxMyMdTvu+b
Kx7oCWrlGepZSu/ENlm+u0x5uySTIoharMUYAhiopSuv/gzPfYKTDjYcmbviThMU
hdPbH6kIqQkOEcI77uj67z7+S2qDjIfXRWA1Y1Tm5GiMtGZ8qv1FXe/93o3NMIO3
WK9yhE3sRBzt66pwSNzztlOdknP3ye/FKmMCOeSGJg3u+yM13hLQ6KqBh8nGB1sN
Jxz4670lDZg0Bm9lkWuvU5sGRmf2lFvOopvySvJ9gA85LJaOw+DWyMr8Av9khl01
xF+BwfcydKbrZwj2oGQutErFP9NO0fpihXpniE87w38R2eLQt2KmJ2+wtvy3U6hf
25CuflARAKWyvu9ZbobPIcv673WVkdjfWIk5Jhp6B7rGJ7GvAU5b0KP3hLPaMmZT
g672BXch6LFde7Wm4mU4qSR+ukyWu5ZHMgeW2t+j+JfoyLdhvF7YLxrjVhUpdv5l
r1RtGLCsqrw8emI8ImO4cQn626LnQYi2ae6EIOXVT0HmCNWUfth1ITCzZT+5y5yJ
g1/e8K4BZ0gcazm6Tp0yf4EmZJfGjnFybvC6ScCgUXJBpzJ1Tw+sLhOyuSFGwOkZ
S+/z/5YOUgSyoYWMhTQsEs2lNCkG8QLIPbqu1X1tijwzGMy/Y3Hobv5pGj5kH6C4
pasY8ImS5fni0Op/TTfMWH2pp7KKv/G0iQ2dAr+gxs5RC8CzeOSAF4lbJ93vAYxA
xUuqzy9IJ35BbRUyZPfW0kn4NwKt21q2b8AQuUEPu2uiUlGoDCL8wUNx4s6WfeDb
ucAUNZ7VuwtskoHYoJ6XISuE3JOvOuGzexTxw1WYLdqt4/pvOhoksVhYcBERMYm6
ovNww+hTi6UaCnZKOBTKtguEA9HS9lBa1jmjD8PlFTfNmX5W/6M5cvVo8jKAqwCg
MdJAPNGLJo5OfvyZDTf9JO3GgyruJT2K84LLk1258009YubcJyR+C/pnx548kIec
h3ZpQp9xEN+8y5PVeXkgTQ8kOvp6q1JBN62nsQVdPjRtmt19qV7KNqgUnSWZd9UT
gSXnyWX/jE3ka7JO6biDwOa2GLc31N8bUqBAvWC4CoaZWoXR3H0bDBo42eAvUtLT
TpJI1M3P/sFG3ZBjcc0t5bXiCH/xOPWfqlqrtuwk7v2wyR2t6oIAQ/zV8gb0FEgJ
QDiADwlsHwydoJhBC5lAD8pbDeVZlBABObU2LDnlalOJYY2bM8taHck7t7nLUMDN
ezmUCWGNpai+ozk5tkzthGEn5cFpLvRlXh2TjHtqYcx4jN8Rv4vKSVwzflc3Mmjh
55Uis2uAHGjmrTshf4bliJ8u5bnB6eqMXEbevZyZrLroDtIojZ2UjGHlNi0b+Urq
A+ZXcAtxclJkfqdhn0Ly5DxzNMAcSJGyxWQ39vauf+97Zea63cBrJcKje7fX+ocP
YG0hYGitgDQrP1DUQk/Jk4rJ/ZR+AQnMHBWmRJLiOJkkq41f635iuouCgHRhuhCS
1Yefh7sevy5AWxGiXneDjTO13eQxIr4F2a2qp3vIofqH3a2hfeOylFE26L4vLQ00
9jSTZAQLZSQIrDtxX0P9CJXLAuI24GwcF0NUXski2SUHwl9SdQ+nLM9hCB2+cjxo
gqa1I9EhvOYNfr1N+gvy7/lvBlrEy24g+D2yhN3Cd4Jkygt218arUszImA7KlQca
n3xQJ4c/3phtWMkGJAjX3Mo7tmdqvpaPzAH5ApJCsdROLD1wYOA/70ahr77sU6x1
GJ5SspVn4zVob5y0fNKMHJb81u7y8Xm4GaKFlT0qCrar27RPc3akqpkE2hQbFe0p
dKdKUIc2iDe42bSdHkLx36h1x1xdDUCpX+5y0FUKXGXolxZ33QGd8ZTMA14faDar
0SUI2uxh6S9A2gnCSWDq7EGK+pvf9oZcZo6Gt+6rCXI96mmD/N+UOrIZ5wfNTjAt
5bRHAYkNAZDbKTQabvXFvdi6kmN6dP06B4zQLN62al3mYZ0v41SezUp3Rs26oPDw
Iy6J1T9uEZYfu3KTg7JwI5Vg/oJu5nNEDFdgv4aE4WFZKB0tqutWkr8Q8TQrEmwa
OHaZ2pe20SSGdLAJGG/csVQg76kWPoXYhijdZo4Bx+sKTY+4pHSOtSW5/xsXX6n7
ziJSQdq1cmelHk7jgX5dhEq3i3PfpwYKCfcZ3o/6mYJKahLIp12g4dy8yvbWYdQr
OYAyycaggBUgD73l6bRCj0BEUiVa5YnuV1OAM83k+VembWGzE3Sus6qNTSrz9Go5
1OITj5uivxjvj4CSXe0BndQQDugnd33+gq8QgkYNr5kDoSjf5SVwQuq8GGbK78pO
d/F7ye9Stg6DquZZRREGcw+5mqGgByyBXhQZ5eq6rthur2e5xLuESwBBR/2sLRTS
lTon5XckRAEVf1j6krMpoLr8obVt0W/kyTn+RgI8Vo8mVx4gmD6cJfbRRUgDeI6p
rXI8T2f0Oz0lIGYQP6ziGKtgc7tMWEGySTGjE54tdbFZrdOiJ9vtujtKKajejuZF
jSgTxKGSe14/gzYzh+1AHFirjUzAx1tM6sBHtEN9o0dMlWHbpWlUVSkKoR9n7jTl
7R121piy/J2euebrZ3649oj7T4DEsEImGCosGkoz+Ub74mcNeMlza8pYH71oPNj3
gNIcxoOyRpFr3cX2Bi/Ee+k0psgX0E50Wv7vB5N4oNL+FUlfEA9O1zrGPTUAz8r9
dipI8qABBOGjjqoo5oPtt1SPd6r1yeVyfa8tjjWQbNgUcYUggIkibkC/hXEwD9Tt
nUYcxQnv8sQy/4+e/LYsc24HJdmrNCyY39+2Av9AgmoWs4pOFysezj7ERqpb1X2U
rPmNJ+Ug92ydgK76PnU13C6mXNpBJNVZJ/xIcImt9KQR+PlGoFmJCFHG16qViVIw
luw+VP3FKWHt5/f85lrXuU4wKkY7/tflqw4Ya9eX+an1qOm3mm3Zi5OPm6J/xvP4
a3BkNq8T53qXpAV9+Hn2Z1PWf2MYbFkk7rvMS3jKTVXdeDZM6k0jXMhCp80ZgVpt
VEDBMQDxD05sc8PCImgifisbIDMMU2XnD+3YeEvtD+mfFNcZmJObZZr9M28+7LYE
E6O28S7klGejBOQ/0eR/p30Dq6BtkAwJ/vRGWF3np6pamItxe3VCmVIw2qSvN5Gz
IlVPbdeX75lWWLvOwlKyt64MUrnG4cuDbcBpD9FdzePSk2KQ/fj48hkhFBqz4REF
fmRCNTg4thW+5C+O1vcPaCbvcD2hTlndh3zlTDLRr3b68rjJuZwERvARow4BPTkc
doBSkkQ0AqDiZimb9kiT+3AMhvV1o+TaJooKfwHAjTPNeiLi+60e1MLE5mERgRBf
YO1Vb+1Dkkaa2UfjmGvvCuoSjP/+uWyDe9zRAnjUTlHYlHe5AcUthtFn28FkJPzm
duthO+MSFdECIeg2SucKe0Etabi22G2xPrynnRvd4SH4kt5OUR/td8iNNzAX8oJO
RL4ynwOF3lmLOfaosP7mLIOlZH/2wl4IrAf+zcT9b6MS8N1IrtOBC6fZaifHVpSQ
iv/+7Z5id2Rm/eAMXai5jhw/VV0BrCyGuqA0W4GeSwbZpkVK2UG/l/9fy/SlILXR
ae1xYJsYq+QqUqiU2cUPD+CMgs+al9wJPCobtCxxbBoa5xEZBS0tkA2JFeM/OGnS
5+SExXQBFvarOxHHUwfMNDDqV6uk7vaWI+42iNq4n5lYYWnC9o7/wLTAcx1pq/x0
GNYaBisCRPGr+1eLCnfJYycyO7vNfuxOhcMZ0y30TAMjM1NVMU2Tl74Ls+ra9f2o
K8Vozhtd9Vtriuj+Wf5uG6sH6KLEu8RP3oCCKVT5uFvVsmVmGlFZVyksAbjbKoNB
WtmqKbUNINIF1AwuEGWvFOAE5Aj5vyoldEhJeHorfmLN116ey/tl6dvbr2z5tmdd
uM0Eorv4ppJd+FbDevBHJl3IJM+dum7wD7e4kOwqZvhkMfPM4bKjpEXNy8eoNDzX
fZHLg72o+ku708vQ/YEWWmXdtyQ4uCaInEQxnmGETj2G9hM/bKSbmu5iaObJnQu6
FP4iFDTV6zhFDapELRKSoNpJcy4424fXTpJTenYya20lEyvNEpYTxxP2NJtXIwUp
iq2i4saDD+EjJCSsiMLahgMh+OgNNHBJGq2RUvkZG7Qapyt8oNASpaVqJbuIxixg
H1s9kcP84ip5YA1Q2D2sFo8e9JLEPgMSzBCtXB/c8voT5Q5WHNDS+p9tx5Xt98tw
1jvNJbU4/TgVasE9hnXxdnQU+8xQG2Qyv6aoZvubR1JGXWL7ZIid4cSCyKeRjbHl
eIGZQOqLMIH9bPZg9RWr61gOYpAyvE+D7v1gU6KkndpPZVHc/uOeINZSp5E9fqiu
ZO29hi51I2uVL6nlpQZzYEfLMWav9UT3MJcZSH7u9crYG7zj95GQU6vkaFZxHL4p
K5KXiH1lefpKlxNmMvD+9C4uKvKVVjLI4AoSclrmIr5M5lI2o6u8LeErg5N8xp0I
vI8biaKm7lP+bnZjjoes8LetvZ2dD+JZf1kgObCU/FsIJPu0MMF63s/BixNuOAal
DMhnYhDCSeeKyrODLbYymshMyay4jZCal/J44avDQ3zeP1FEjdrS4v76y+MSsYde
/LXk9T9kltFWjxntV+fTWeDsKlj9cxMKfBLEsj8FB1GcsqsiuJ6Bhwuya6doy9Mu
5wyWMMwO8ALZmeVjd6nD4Nr/u3bnpQUkJN10jplVd9t2ZCVDUPnzyqUclQml7bnX
dg5A5lTQi24YWHe+Os0tgr5HqU3qE3xXLSxtVeGzKQAlv/o64XUE/4J+H6JRnkq2
yMWq4nsIKNDBZvIeN1kJ91XHNe8ZgSUxW3LSi6Rz6thUNg/37WlAsZdpGZKsnEM/
lLEP9ZShMMe6MflmzeeDtoKM4VSTUCo90iClPeWHKTF0mPcuxeUpWwrZupeEx7aW
koTPmj9RM338kIBwzqyKu11GK7ETgNJk5ND3eU/EQOb+sw01Y4eCWZXzj4FTScYL
BkKtNzTxgCP+WCOJxC4PiMAQXDatG4KXBGTo1JWTEsbg2OuszholajMDeosHMrJo
ymPPCCKBZjyXri/i8RA9ypk5cu/g72OBtdVJxtANinb1nuD7nCI8075gBUhDKrgr
a7ZpVeCoDoQuu0aZW9sFTrCiRH6qHfsDDEi3FOSN/MYcy1H8pB5s0ylPRxVK1DdY
jbR/RvvIG2ymnD3iOw+5KlXkVXgmB1qC1zBGVW7uuZBu7zHKjSiPmXCO3CyfntTB
DXWStn+b7vUdY/0JXhG8pZiqIIkDDaVSBOq8BQuemqzdeDnEEEoQFYtEUc665rx3
+rSCqeslyhjffpkFfm5CTrY0BdhJiUaya0D1ryMgn0y+I7Y3sHfeNX90Kqyp5VX8
e79CwljIOhYEaEB41/hHNFvKJg50P5JxCsjdC/AOwgdt8HU0yoJDFc7JSz8YMOWl
QPW8G+cOiZUeq+8jO37LP04K1lXh2z6X/QC1RzeYYU0av4vfcOerBpUb4vaYt0Ta
xEe6zCJMfPCJOfZHDRJDLpParKfQDxdomXnVGLtC6tZQhPoZikklP/1dg/a1xPxd
NPOk2v+mClC0JmC1Xt/5ROCm3jW5kxBD4KC9Nucr4vyMUE+x3MyWgFVF20IS0SpL
LrVewCDW2PVsgtmZoT5z58vAMsqflbr/ugUPEAMrtZIGtPWpeHLHemFvqNBa+eVm
l0EEXDPn9VoFsgIbgllV3SqWO0i6vgJKyum7pZREQZyVjMg2KG1g9ltIaVg1OqiO
KFt2uZROSF4AHQWdqm3w6MbLlq8VGtr0ARUpBa5lAqsAAcyDd/OmqFUynXsVNO/C
M+EgUz52Y46hFJLtltj+IXvRMNV220kd9zes5ks+RWyPwccetF/rgl0+E8N7ZK4W
v9eZ+HIUBHLFA4zy7P8BIkNaRgh61CTNv5D59FUwO9yBZo3NWTuvYmvLjeCouGxM
B3sqiAQW50+mifXEuBUDJ6SRTexSYFDF13kc4eyVbj1UUMTVv9swOKuMFB1IQzxk
kFlaRuEphbmg7V/gZPvqNttUs4QFpptKlAdBsMy/AiCHCrb9s5yMu6XZlOgSw/ZL
qs/wfDNbRHKQLzsYzdTlt+eApafBX+cXxwqeqj3moYZ3f7Pro+HN/8mcYHIZEZM6
KzQ2d6tsUMC16Qg/qwkafcNYNYrPSjvZsbHTdIiBQdvqN45Z5J69YKeMkgKsgLz+
RrpCI7jhoxW4iLY/rMwRC+Yt/AiGe3DSiN7Ida3AW2qPp36N3Ddm0RHJA6MQihUl
mrGE1yhZTfu068HUxVa2xtVVM/p+OM+BWb3gHzFvhlJFotdJhGu8XaXMAY5R5Gqa
tcPgf2Dyk5GR9rtTYwodmrxxQHLiQ+30mOJLPu6fRCm7gy5+GEgwmOtWqTKUgXFk
6HWQdjK0pt1FKoy8UuMqVjh8LARbTHj6PmUujlskFgQtCs+fWEM7Fb3wg9tqp11Y
ZxTAE3+Pfpa4chtugfczMSlIYwxSotzjTUDGyu73wc2ElPll2MZvk99lSEgVBpgk
pA5UwYUu7qnHYOG+pY9T8HA+MZPLxUioUT2T+GVAww4myk84PG4IkVAcSvPin+XY
6VeBO4PhHxW+Vsmc0TZpt8DPtloimpNKZO5RkpTgcK8x7CeMg/ObSLSh7L5dDdKS
7kn5hDvusmbC87xEu2OnrMTPE6pVh2PUXzzbp77aNdOGdYRF50wA2uv0v524RgDv
n7tyw0zwzRKohjoXF7xWtjsHJDXj5VwJgGpjX0IopQGeJBaX+NFJtY14g2d/VYKt
XZfBfghoTsjTUR0R/MxcHfvXtuw7Fjark9iBog2mCK9KFDzxFDqwykOu6H66g7mO
KYkqdqrE3y9N6eqRhtRsdHFds/4lJZb01YVacEvPrkxiKufPzHuB8BEB51G4Gj5r
8CuYI1bAu5TWqmhxsl9klzkfUErPS0OELE3BW1q4EDXi7bx+xkJCZGy7ZI0Oeq1H
HLCIza3Ul+WKAL//D2NjCUHBdK6AcNvNVjJz72gJqtUZtz8lqBKnZE++JZ9ePH14
FWh2w972+l0f85bgQIAD3VBGN8/YbdnOtOKhIUneTZwlPhMW5QKBRUE+cU1pQsPF
4YTUIyzL6uXBdGHczz5b9t1yN89N1trEWxPLy14LQWbBMi+qYYqZ5xXb0zWyxTNN
ZqhBFaKQq3s9b+pFmCmYnbVLiavq1JaBoDO30L68IB27Et0IRq0errgfhhkFq7dv
/cJlnkWFZAe5iQKRxkTosUdggUUrShikkClmixUz75syZdbghGNoMt1JOwY7AR52
CcqW1KJBgTh4XTaYBJR4ENivOCKYrJ+1zkP2MshVSm5AYW47NONVzB/wYqFKPPA/
yvesMRUW6y9rQaKqVKASaBB/XcdkeFlUwkLc3X1LmYfqJvbEQKY7UE5bKBTgte8F
pIU7usxzA0CfZvGN2AELZcnxtGq8GA7hVVnKxGfmEwDQmzqSQT8BCDw17h+DgP+/
1JysToCo6sosOTYV5UZhP6B0pCEUxlbCutRgAJC0v94romPHSde/j2x1LnbEN8Qn
D7M296L2dbMPNgO1QaDxaYbb6J5mgl+Eh70Wcmbw3lccN7BqXIOPSvc5BKf7/Q7t
7GlU44i9g8PBMnrtciEjL+rZQgKDNv5DhEaU4lwUArc1OFJ9n6qFHSQwWbhzPJKi
Xk8OjiyfOr7x5ZO0hq7GpcSTHfFQ4kgpqp6IcxTkEopNjhggOKfnNT8NApY//q1c
lKXLL+t4fmMZJOR3bsJKNchbIoFbmOlqSNaEg07xsneQiKUuHbo3OQaTkExhtm48
g1IHCwWyfuWRClbGsF+i7J0n4W+obbH9aMa/g4hmIS+Ro3ISDPFmxUdnRlRXuS3B
K2ym/bGsWOJUrw3MQ9sMGhADaWoLU7ugzXv8Y/212h+N9ArxzSdMhHLKWteQvSLC
ustAc8lgNh1e+VQehcwAoapbuQzJJu3TxKjkqGuhUzsNrdv117X+ivfDiAV9S4/F
4tXGKkTujs7pgbbOspZEk1Ed987le/SuEulT7qH0cBW67FJAaQUisTiSJ8gNMLxR
nEqf73Cegy9X6KomRYgf8QhUDn/O6v4f5H7mENId0Mxyaw7zUXnjxjdGYIxul36+
GITLSM/XHrCLF0U5NtiIzpkY5Oz3HEZt8UgVNMmmFAdI58glDZW0T8Yfxltvohm4
Jc0owdCfwfvvUdkXpUQ/zoSDVZleSLeYKc84SLZOMSi44MVydoQcEDOD5cFA4TB7
H/Ozii+0AITUjtLCK9bTE3qBy5/UmJF+8kiy+5OYDH3hF4ScKT1RL43xFKmc5LFf
hPYPKkDH331x2dDBnfy6upFsu65gKQFmdls9j9tR1LBxdBCckQwyEGUpxPRqB4oJ
RW84r4ys2s+NlpMVo3OBj5N+c6clwrGo+OqMc6dVQwwrxkobbtyOxHd4S5eW0yHj
4TPAtRm82SBKceMSvBfDwl917U3Fy3XM27Gn4MumPw+WtVNlUGJkxWCk8aF7xviS
RWKGhQuMRa38WhGmNvm/G8RedIKb0PAz0+EGIJZPK4HI42kQJIz7y4HawMWeFYKd
V5aBdHigecKLiV6Sww1czDbtRTFeufnbkcMQJFwHL7SR+9InElzivGHHpax5oc1D
KFVdy9wkHqrWEYX1v0Kjtqc9Q+lQsUKzhaA8cCcUEpc/eREA7DGO48RXrPYpgvp7
0x8c87X+yks0JRz9v7gHFInQ+70ns2zz86/mEQ8aa4jNOLMyCG17b31NvRKSEEM9
pzh3wU/GuxK/KN/KI5OkblxF5Swnd16+GUEVzpFnN4BcJ5aaNvaRfIcPBANrmHoF
TI+FMWwlAtRQ2rl58KR4TmwBZ6Nswdr46KBDblww8uZJb9bDG1lH4FjZ85kGHjKw
M1JzrvyU/EYl1QWj51a9kgqQZlTccsRmWcOzO+jL+NFGqjyi2VzDuTcV976jdwhj
2aIyLfQFRGph5jGg7SXkUhmuQA/5dbzUwkXNZNvwm216kOvsvyOfb/2vkpFObiwx
noXCzLamg7Q8HOeIFdUmAZRmwls32Nf3NrAWjSVUuQBSrkwR++mL1BTMLkWETT58
ii2WX75HpS9x4wGhE3zEqY/z6vklVRj/uU5KjHeJVn6P73SuAoS0pEZvWW/XCA93
rO4HZAIDubjf4XcKeFUPqbtwmWvzoDt5cUpCVz+NvC/18IuE0ub8f7lArBNRlwTt
WWFiR8lGzTX6pwAIwkKXKtEKZgAB8wHk3bBSdL0Ki9pxwYUeFXOdkL8NLP3AluUW
k8/yAVMCEp6AjmztjBCJnFctrFOCbVBp2y2b9RANsTwD758tjRiF0lzh4qym8Fx7
cykBFsRXIObbn5bR5sCDnKwbQYcQayCwFLj7EDZaUAgkZvA5RwF2O5FuA9DQHJ8r
k+29mSRtLtsXbsFaVy/GDgQ7MSXn8VPqS9Zd03PBujgnOedVjEEnVwwIOGsRex3Y
VeM7nM9QgZqFz4CWt4q9eq1N5/6A904SV1EQMGsgIskYQzfS25U7hvBUv6jhCDmK
19yv7e5aTiSzymgzbncXpkXrdx+F5OoJT9D6G3MimfPlhTBQeAyzesMNTk6z6pTi
A8SvjYmcfl5yhHMbQ4Xm8oDOwtpypobnGOXx6qKpHdjtnbfxF3MJK33hy+G3z1pa
EFlLIICsUCSLYE1MT+5toN0ds2SP4phKjfSW36Krk/5sOaFIUF/Px1u3yEHURGuf
eFsI/wViRw0MXBFBocJ5aWiDDXWsSVJ4y5DiIXSgeu5AioWhugdYh2+P0fHcSjmb
GqVqQibCr4q8VdtW14DeutSMvUFoJlK3l3ihhuZFz74DxZil9+VBIm9ITgMcRCem
usDoC2UskomkV7qYGx7VhPkBe3qPEBIxKT4nIf8vcHLnaGEJOgusgVNlNiYz3hOT
HRv1b+xFsIYcmwPOhwER7UqZaBaS7DCftOrKxBcbfrNgyVU4sl26iDAhR/ATrgkq
OATardSIghJRgerh5+9TTKFdxinbQfhTfdHaHih+9dHUeJFbDctWZrm++kqAFPT2
RZF1nhHUVsYMT/b83//Kys1mVPCi0IZXWkwUBcykONAJ5VzP5Qm7hBYUFuMQwrQA
aWRjLgSxp8O2JIei5ALUg/ek1nq6ns1iSwQnoa52TcDbqgb+j0OLxg4yISd2U7Um
bLsiyVPrG8LZxlisaB5pIP9wK27iY1nW1MX0c2mSiy5in8AHweqMUu7GYgVZcNod
tbCh0GoKHHGzNciQqs4QfFvwl+fXo15p5LlqlfXpWRtp2ERsZMxurzhU4bYeYNIZ
r+veN5NoIwsbJd6toweZX26AbxwqSePrLB8xHcJvIXcfIanXaI5DgJLCZESGs9q0
CE53ZWY8cb3Sp5ZFa4q5U8krzG0s70J1BI5wB9NExksXya9MkQB8/+0YknibMvA7
+hgZbYjyeI+7E+oHrFxP3kDjuMxatHEQoNR4/fi921myD0xCeU/ns1tKWOfUv82D
1t/xH9pB/drzFPfyzDUoIiPQwaigqBY9mDfxNHGcMZj1C3HMBfjZT3Z/wRrbhuwp
dTuVwg2UQRzxWsBLiuUHADobnFa6rEsJN88wTxVzC3LXP3gRNek/rdyxNJSvydL7
vtgAq+2j180wNtpEig8MnB6iq9jtgteYFCb6q/+I1tYy+Q8uimmZ2Pc7NlMD+bwG
osRy7A9jRZErAaswlqm1q/QrV70WHk1JXSGywYuQ0PbUAe4TnvS8e9sKvk89gGUw
Lsrl08OfFeRU07qdBoYj9SgHr+i5a/r5pWVT4jOq7kUXYuhO1yiz1OWku/vwM2qP
XCl0Jc895SiSCI7DpQ0Cv+fWRCk53nw+xUdh5QRxRsSUREUI4Oc3XNS8nTrJuiMg
XgzorS/ZKuyeLEd+7dxQS80kRFUoAP7I+3eETYFmurieasxkBrPaCbC+Alx5//PP
hNA4P8L8kxNlrIOmtXBlWRI5JCItXbB/RPo8BqHJOVsI1xnoAxRWuaxiFbc7LYRg
gDAsFMKyoLcp6We0CJIir5j/eTbWibysvSjr6D67t0++gc1MvKKykN2EYgQ7N8p6
5FYlHqawZ0yVjA6N8JnPZOnpGyyYrrFX5uIrR0JFFkxosm41a9j09k3IrWulDGB9
5UCfmBhghOSvnwlwk4UXMuz4b/GNvNn8B6KwVR0dWRBPx1zCJGQAS8HYc/OqqviJ
57Hk439BFRcQUNrZWLiwEGOPD9zLh0Uqsi9JXWU9f2JM3rxWNl8v88KIz+Hht+mo
UWsKdH1MaWo/mQpN24h96GdPduYNKlZPWW/39pQd6NTfOd4f95ZSDc4awPpRWrts
URr35R7wwOjjFzqUe75TmrfKoPk0/oqTqj/nI1XSKFPVvgK33h0O7qhTIqcILB9u
ScF1UikHrCsx4hiVrc93s4PKgbkDSpKH5ymJN3zd7FRSgLBsR5Y9Srt3fTYT42QH
7vLF5a3xHkzrP6sw60zENPhKddKcYp3YuxQZytM1RmpybW+BDjC/4lMpDjuZ6oJ/
Ee2carw4XSaiYoe+pDW6pcwdM5jrIVduHeGq6KM/Ct2i/cyQQ3GMn1OxFmoS+/8J
zw5Kg+5k28pq089eD1U6aZqmTX2Bz5enogSvThfE3irv2S+I/Y5xkNhuCdriv5zY
E79KwDYEM9s4HXobn7o8So2i0YHm80obYKUvR+j16u9aw9sLdXxnWGfARCKDBFS4
LVTPf4ukwSuXTcpflD5Yg63r/1fG1sK1EU0dwIQqfXIf/+u+wi4j5xpzmz1YUMFm
1SrtJc5DIYj8BEHNzcCGdb1P1260ZjbkxarX9O3fTcpf4a5UcxBxEhV/YgBW1UM6
ByMhMANfOs4kmgoxudJ/LO/sfKz7g6ZF5t21NNLhU/SNogHSX7QaEWUIwW2Anb67
GPVnd6hQ3gKXLiJGlH657fmj9qaOfqSoGfWYFsLbzXNdcTqS8ESQ7t1f2z/CnHLc
laNi/bH8sYDIuy3+Am6nOUC8ne4tDGTi6+Slx1M4M09ExC+zeh4KcCCGRVdH21HV
kf8kAzugI80GYKZXxl8gDF1OOZfJ6SVtrpjsuHjaP7Sk+JxjD1hMe2SuhNGl0Pk/
p5fv5RDbLeDviyAHiBhcYWnqlyqzvSOtClG4Rc+gBvXvZKRy9L4rsPkylGwZUHn5
StnhzbaXRQctZUN2XuxWwV4grlIoLuxuwKszKhGuaoNzXItuGpw/WV6tfZlu/y1b
2ZV0l1/SMnjJaFO/wLAOd5tzkOqrXuOc5Eqmd+8bMbcxvMCUMblkIS4ghZapLjbK
jyluAiuQ81NYSBsURBtqfBi0gE5LHTVrsvhmirsBs/9wp8VTkuM53hSdgiG8tSZC
1BbSdCcouLVrZRsqWyUM4WUD7lvVm6co4nE9VBTDG/XDYWRQWCoWSWXffh5y4F+G
v+mKhgxf+s/nflr8E64H6Bdoh6qvTLjaKG8aRKkPnBe2UjmL6MV8c6gIUQP0Kvty
bWEBJW3TYGKQeUF1hF+ph/D4nMZ3D0yoS0mpMLXmbTlNbP4DVojciJOXgzHcW9Yc
fnSegERlwJd1A8ePMos1fVf1dNUVg95L0dGPEMwETXTkkpYkWU/DbFyD9JHcg7Uh
7MtX28StLMzhsz4sVHmpGfUJE4Rip4TnRvoffSIn79Jq3EJiS/4gfuXqky2vgTI8
QgBeDEn1WCZde5e7S2/WvjsNTnSFZGMc0mxsSjkllwa93XJs/50UgES5XMmECdf1
4bgMzuFsUFDSPfX1FpCPz1InC9ARVDl91ApegkOSKYESuq7tlsWmE6g3DfGQ9GEj
/fLV2w0mPx7jyMmYm7AcxD7O8Ft5NkAJywGmy/80dVrtZV8e+y4ByXZxbeEaLDKd
cZIqB+BLrVDEL6wpZtSCgp9SdB6oLEe7TPhIzlCny3t737dsaZRVXQnFeJLAbE/t
PzVoeIOnLgDiAj3P1lsie1brnCunsx8eFVBCM/mDrWkvGaDKr89pc4bY/5mAwdjd
vkphu9f+kfhpx+cn5ZtVNYvzQUJO3hMPul3QmcGlRL1/XOJO8g1sLWbcyZNO3sZ2
/NyhKKb86fdCkzu/X/BpNRb3yiLjtzFQJ8emG5OFWRuKWgWJKRbji8jZi074hXyK
HlX6QuHZBD9r8b6kpvk7mAXQw15yYr8hRh1ful2mr8xMS59wJw7oHXbByzsrgVmw
gTgOCyM+rUu4A4RFJ6f8OgkCHT+6u06BVOqRE7dpOimAE09IokTWQ3UjoraDgG14
iSKNpRFEdhuQ1OLiPbVrGPQBLHrPZUgJ9IPgpNd8ulHRdqyRk7s1ZbhMjKuyLuyv
oyo/RrsZR2F+OolOxSGrpXAMexOB0sEALKgkRpmeCXHw2PVX+Tj7xMXqlW5ilzpu
fLPD7EXH38DCJnP869LSEz1OV2Hw51222C6S+qcIaUCDy7jJvkSPN1FkCu/8NXfF
UXEpgkcc8+892VDfTyEuVIfXTvlBNVNFMlo0OmLaY+AfIy19PYOnLRIt6zUJxIWt
+raSkfB5XbNr6RqHQ1Zhp/ipWQj0lyaVIUMP5dYxqELi7smC1HD+8SO3VUIUkdj7
rtMAZI4xsFd6JJWR5chGO6ZkCsq9hJGxBM6P1vTKxQoJWiRWQXRu/ZE+NoAhgygP
q28sa3U+LxNU5YBVJITZHfATWdwbPBEu5dYlhJgoBS/KzmITEyyaWyrVdFZRJHfB
SmuzykjxIW8hYJyZZxUMAEzgGvkvVIIaZ1Mc6moc5MAyWuyG6BwqZxFCyhan0A/y
0g63YrKH9B5W0DBu9yLXLhVRtDK3Qp4Rek+863coeMa9cdU4iDrwdcRCd0OA/5P8
5Zs1ft9z1T7SvFZqHrb29RjbJqwSth9QLFfJpWvXJ4F+uY9KkVKXZ8xdQZsLeP1I
LMb2T0aLHrIGPzt4kES/KLAZMwJE2qViSaLWM5tYis3qlXSnvBwvvjlsWGf4mSEz
DWUwHF7uveJLFIJCaS9nTb/mOefboL3lxs5TmmNXyOXIgullKdqYpTwjRyfJsFJv
uKTso645aPHFP6HIbdK1EoS/n/ps8FY3xWxbizj9LS+roxUdo11GVvt6zy6dfIcu
ebKmLkH/WOprromB89qlhMWdRpDhPn2x/PMDIK0aGgHKMTDJo63A7feViIrUliw1
XTj5jk3W+/lA7/GNaVpiEUfTTlke4ZzLhRRawo/N1GY++S6Sz/Jx75W2oq1rWkih
nVJv3AIeDWSPqXT8qgkKdR8vmoGEO4EunPfpUnEMv2qcLrGEewndP/O78+45l6CT
1EypLmL+UQ9XxYxAszbkOUiyTvBL4yPMFQO3owB8ee9oqmBpyl3Eo023bqeO5A7/
ubzY9tIFlXcNX5gQP7xlZ90omIknpI6lI6/46lG0Stjev8OMvmBTxLAG8INtg27b
anzJdNWCkRkJ869B5eDkiJgTYHXELHjULuvjPkvbO+PzWVeLz5LgPK+N1gsYcerh
OqciIHtJg6hfmTUT1gy59c1lQPgQvJHDkRa8coUCjooSJlbTOrntoyntSMJRA8sN
zHek2bvg9DzZCoLYz784uQ+dt+aFxwJVkubATW9FJ4ZzUv/MvxCyPa95K9gKluZK
rtut3TXKtzC9EdAcmV2365iH7FMamBwMYM4UTdljg5nC/J1JOPF+nah6NVTyDEM0
qX+iASQUbvGL2wFOEpScD75fZad4RT1K92EpEjb46duwaEkT8G24fBKmB4I3ry8n
fQ4zrWYGueXLuR+45YXZlsq5u5yGK7mEULySJoALux3aCluGASGDN7PwCjsMzvp0
QX9OcLqbaJVp2RQH1GLBcH99bdIYXpbFWcmUQ2LdUPTtHK2QXmhWR7jyzs+kx/l5
RANeuJZkW6QMjdRfPHxLNaf5DgYkQ2v4o2mEqiXyvkis0L9UaiHV8X/FgaJV/OXh
/Xjvr2LvW3HW/ue/+PnsxV4tXPloa1d9y0nSntu0TcHxr1cvc6IGEMrVHDwAhXpJ
zRLW5JD7YVpuh0bw5/1ijR8c7Fe8jXDedSbnOe92tuxr54GKM95BuIC2peTbdXOE
z+1DsA9bFZFL+SFqn0DnDQnW/42NK5rWtb2qGt0Sbd1AZdxBdxddr18FL0qp08g9
JYxLOtlKN+Z4SjyJoLpA4jsiJebGXt5RpEjlvz8XiFcuWHDeQv9mGbB7/k+iO3XH
A4T7FkXRDU8VpSB1jyNmZEqojbA2QSlFZbSQutFiZhkKSNI8S2xWS6f46Q757wjH
w9AYS/SP8ct37rLFeTkC9O6RJNXGjCPNuM4r+F3CQvz+FfZRfxN7P9oDqGpQu9gQ
cJbPUJpjoCFFjwTsUYcVmGmdBfP4lKGKoVuTiSa0FKm4HWXTY1sKk9HFwUWKVSV7
CPc3ubGHRtX1QQ6ha24CEe4RpyMgCi/t2UNOFjU5M+NK625PGjUVSNsuBkrtf1OR
5Sl4b+T/mi0MwDvGU0tuAUOYrDKn/RSRbeqc2HEERagVAiMObFL+IMC6OczVc/v6
OKS0dL1HX3kU0M4lfY71LYHihTMcuII/tubfIwUTxvxzMJfIbFnLWEcs2uvwIyo5
3f1T6JueYklXu7OkExwChzOj4usCebXXIg7owVQgK9HZYDQORd5pWE7/AB6CX+Q5
pzBah833aHiFq4Fm0YjVrn3BzRcBvDbUfPpUmsi9G8p5HKIXb2RGhgc7Xaj+FxfD
dFY3B0u3POROTx8DedaKtiJ4KSk84q4e0emvfjlmqfYrN9ZsEW9+DxqACBnqbrr1
AyDtImCIKM4hAE2/LfxU182umc3jHJgBqHQd8nhad1EhT77BdKYD8cIKHJy/u/VV
CT2clRmz5dM6pADO+IsJvAjRsY2TlCCR2o7f3gq+ur3HYa7aFND+uuSGzTaCFBm9
cXvU1fW2eEwNV85s1NQtkmtU9QgBN1AF77TnlYygVigfQFXfvT3Fna3x/UAjRqhW
nIvqkAbO5DNpMS0wQ596tltom3Im1XB5DUXi8w0QbLkOZR5HQSGl91j1B/qN/JR5
ixR/aJ8UnXjlEGMsdXG7SZTWnzgk79dmCEBGACw86EEoKVE+ayBG7cHxdLZgRUU4
HtM9UAkvbVhyNiWVXOjHBWxCGuF6eNMKHVfBqn+uKaau8tk3IgpR9GMixEjz94s3
+/uaqLuP/ot46f8cKBBtcfOxat5CTnxFsIXYBy3fUQhzssidDYAXgDw1gmed46hp
9U2AwiX+rl1Pl4Mc5qjh65AvC3vrO2hkZnqhItUHSz588Ejhu5S6Kw1mNuxvHRxf
5hJnCBJDtMohZuU7DkQlzij71InyRyuO+LD+6xMCIXb5NmKfS1aTcjZT9jSGxxd9
8N7/xuozVwS0VeLtf1Nwc2W1xdErqILyhM0TvMDm4GHO2rLS8EcYHWzl6HJzRwut
sCm2gWoUiskaJNLtk+RDhe7RqrYCPAvh2d6rM96pp65T4VbHTKYugICleHgMcwNw
OnTedLTW7XAiTloRn4TNBOwBbNZCAlDuhIjdW4QTsPXKKRjpRGGHljX1FOfA9wE+
/P2BL6bQgs1NYZG9RttrOR7kIfZFgVIXHzVamW3pham/GfWgIrDlG4O201YBdhIi
0tGkYkqCyGGzLMrFjhuCeB368c/YzZXqkcYGOv93mcWPrXJ/TandDQipDFysI5Cu
yXTuudHrv+Mtwi1Ot9kfnmlwAYKkTVubaR2+Wgsru8/KkwK3NKbRLPCsYhESFinR
W2QMrncY+YA49lFqAA3zPeOnp/EZIDG5LdwG+FL68zAuV1eql2HYWd250gjIVth7
TGrkkYSNLLD0GycsaCcTnasgFW8Ki/Oqwn8vn0d7p63T9b0i+ZmOny1pDluGuic0
TFujwCTgaM3XUhbVJ/Y/ETd4QqxIBEnp7CQvR7L/BEHtKkgPIi5BjePH1XDjP21P
BNVPeLrre2Pfiekm4QwBCgpq1A99r29qvF/xnAOdRe3KsciOCHtpd/0RKXyWKeOl
UxfTM/WYv63CEgB+fCgLdt9AwbRSDYBtl0aPDwVSFf5AEUn9dsw1uZ+nTZozMO8y
WpagWrOZPiBL/8RLkAfoXEEIUBcB6AXTHPc53QDwcb4lqBzoonMeMEeCe/E7Xbt/
4gY8fitujzDWIeySungLhMXAZGuNj2mJFX6Tk+Qg3+03FYFtUF3j1dzvJz1InBIJ
TloI05dcGhz3pHOpTPxKjKtkQl+KO9ouRHH3KYA5+drT5ZuY/G43Il2gy6wyLdw0
qUVJ0v4uGGgDKf/cHiHXTaNkOdrEOYMzxAXIPNUasvloTRjw8rGT4XQOGTPzodNK
Sx3UObNEa3MtPRK2NO1/Ze3mGkpxGerhUYjM4ah+SJEUdU1HfoTdGcRELA49EW3e
hCJg5wqvJz+xaWEX4q7RXuYNJz9K/Y1lnwb3UPrsfIYRf7d9yxx4KB9sDtToyF/V
JUF5Rt8k5mkho516muvKHTrCO/htUyoOdFB+ycUDKuiJIKFpYPoF1G7ipfey1Iqy
KcxKKVmHTJpIpZKsgl3JCx/Ea6VrN5jcAm8uDms+u1lFAl9ALVIl9HVxJYXmQD+4
KD9zEWgDYWPpfHImxLgWLcycvhuRPrkzh4c4hj+RsjIjO51zk6FD9mywu31gysZk
cmGn6LjlZO6hVN5ojmmHGSL0eq7TUJ+rw42Gc5cOL9QMV9eoVI0lz98xaXQ2+G4S
6bbhsa104J9LYDC0RCwnYQFknJdyWbQI1xeA5M5vF47wxEszsTnhHUKcV21THUkT
Ph2pOGwaIOrVrvf46kPm2Ffmy/3mX6M8X9xGR+C0h6CY3QDFS5qMbhxbpEIo0TiT
YcaXXBi6yhckshuQTWilk6CFC+D3LMgV4rXhh/u0a4Beu3jbhF909cm02qkjuNBt
TUeeQNwE2dO5Bf0S4tv00mNRpItjWWahFQ75VdUKeItfTsRXTI689R5SEmgjBuId
NsuRi7mpGfhZrOHDamUhmv2aapoRNDtR/pXFq3KZOvdPyk6r3yPPzqzPSUSnNnk+
r6D2N3k0wd8wvpOsTrS5n08agGYp0xeQIU7adPvPVJvcWgV/xiqPWhw/PX+aXW1j
fHELKi0XlTkeEsbuIJ1i5949AbfqZWmM0FKCkaLrZJat+l6vAt6GzJ5mvqIduSZq
vh3YZ7sAPIRSEdzwIh6vVrumaqxAY04Vksrpx+3d54d2gqdcs1A/RZhl8As1ztfc
54F/iZ5f0skQA5mgJdSCWM0FWExsGGYOYmblilc0J6azG783vCxCAjvZO9BpAWpA
pYKpBpU6nPgv7ot3pitOFDZ20uzHDoYn1wjlZFGr3TkaAcEH2qrP0Liv/dEydb8O
MA1p15+G0nClPWamP3V/SKtZMd4CB09AvEpsMgwG6giSLPpRxKggu78tPdlBLEa4
01ojr8YzMIZ8mdApVYB2c/1f2mMrGwYLZC3NXlHamjHPp4pHnpAniEmAneYTQTaX
E9SZWnXsUotQIduqj6hYdGFAPQSgsgADV3mG7+rfjj1Ipni724gOtfNHc+nLq3Gw
fJaI1iU7nyR5H1OTHwrHFJ/LzDIpckT3ZqEnsBdGACwcnlDnsN/0THgg8hS0p/i9
PluTeajIxmpJ6ggaT3mtdJFQIX//bsl2vWgDW9zNYqQ1YjLNwxLzzjAIAZxLSVMi
BGLl/j1rlCg1qf4leM2ZCpKq6aTuEXNqkiuW2ZKTxV72sGosYA5m3115PEZGUxee
DD+FVJKCyggyn2idTdrtAzObdxlCsdrtuYDGVaNK2l0iAtJ79++kkKe5tPXIBWSS
t6hsQvnqTCwfAX04tcHlu6+HJd05BkexzdaYlR3CNcLgCbi9MXvqKVgoNT1Fenmi
F1seSsdq3Clz8pGCvpvK/dorhGRqXq9QUzN7KTVCy+7Tdz1gKlGZp8Ul6T/Vh+ht
zmQYDbSQm1JwCq3uVB3yPDIio0BMuv2VnqgotGFmhVd9VMu6Vvd78T8VGZb2UPRK
gQ19KTK50AGcYP9PzuC7NIKRj7SUbA1a6jLpbVRcz7YsvOnLRJ0dIMGW3ciBX2vF
xKKS+XPrY3LmWcnEZWnmFovZA3qKCmZ9iWMHPT4r74tzVn/2U72VF59H5DroDfLz
AJZC8WnzHZzBu21weROCKZVlWR7ExI6Q397RB4Ls2ovQryK3Ie6cBa+aHxYVwT0z
dpSTHqOqEvW3YA9r3P5sKN3ZuOw0IPF+zBaWekGOH7WLYzW8H5lvGA53kCe4J+8h
SiMnmVa/oXxW5o+WhjU3OETQTGaCfe1GIy51gE3taicPHGBO0fg2hjbNXh65e3nC
vQduVoENXymFZHdI4b4huSC6aOFpzLfT/3jrEat7vyWXT7Fzjl09ss1Qe1ZnYPgi
/jhp23NgQEmnZxPHJPubaLqRk8H7BSmYJAVe8xN9WtOzVTSY9wmlNj4VjzzWQHxt
19dC3hhAT2IV2eNelqxcM7i8sgxyJczsaF503eb1FMxNuKxh5EBkza05WMK3py/q
IdKffAxZkKk5G7WCaRoUXvvLfJ88aJdI5x6kZxTTeQZSYfK0kfJVExet0P7LC2Yl
nl8JFvTostV7t1V+LDqAlgN/LC7gT3xInRsCbVMBNo8uJeZKP0DTBidrzj5u37T9
PzjMDJP+frvsdb3fAEPiIMyeqET7lFerEDeC7RqScf/bDZ3CSwm98zlFULSW8swi
FCAkNKkdu1jZTmZjOrXlIWfbgWAYAoTxZkuz1qKuNIWl8SO/A0XcCE46on1z6uQj
aIVhjoNSkptQ+B1WrycpkYgQBR8GmraUTieTwhYLRlvAyJOZPuRaQj8kgKenLH6Y
uz0m2wdn8QFOf6YWuU/Ev0kKeRSSbrKpq6sI5KEt5GeaEKPqX03OunYqiQmAEmTH
fvcLkxv4OqQJSbMnLwCHhXWmgvcOqcUIS1HFWSNXDyZ6ffWHKlXCG1Rbc1fJEBxd
GfuOO738v+SbDbc7QX31e3JBSeOazvOY9eaD5enGd1pEna33f7V6hdJaMdZxfzL8
7MdxjxlRnogIQdgIKt3ArL5ubg63B4DZkpRv1gXacB+TkUltkBw94aHqN9eqMix/
OvAVV1UXJqAc/Ls5TPSLYfufWbheAOpunaFioMID+uy2QmmzSYwLssG2v6jrlILh
p9sQEPQEoppNBSiWGFklyjC+eyNJ0LRb1OjaloqNOAoBf7Ky2vSqLOozMqvOK7qp
4+zGT7mmzBhmdBRsVPL5ZtWksqXh2o1kd14/MpI83H5L9UWRnEYpLTw/6p+T8z/F
WGsb1LA+6BG0hzHfL3yrAHqwpGBYOW65FS1dViy+p9vfVLl9J9C3Otg7/eCuvAJD
BNX6jpGJwvaHH2NKkCjkhuUzHk6NL6G1r2ajyL5CCE3y6S7hGaE+6Z8wbgQyUJcc
TK+NwUgECjO5sNFzmyOA1tuKw+7Ip8XAeIaINPIM2nwEjLMmQ8er5CojPq6kU2lu
t2goKVlPkkLkwJQVmbWvIgsLBOx+B9djBsm74pLRXXqXUVFFbXVc5920FHpYTd7d
mT6DBdLC08z/CcKM8+w02mHO7CW6Ty9yXd08z11A9Zz415QCIcsz5jeh+AQ5vn6s
HHzqYYRwsht59o9HA5nKG/ZUWetrVwQaqcN7hRB+9c1ygvuxzJ3MdL/vXkTGxfUC
jPzqk3SisqRpdL4sapgRmpFtR5u/G4gFNp6YN+Jw6g6fSKG5BMmvF0NTPB5Kgk2C
I+xmEReTZgWKwQ2wISMCm8+0Uk+9RkT1GwKqe7b5ALqCNEt9wymBbQc/d7+PvS8r
hYwKMKsVWs34lgU5Hya5zT6ResdezwLlmIUuful4EgfCCgUbPWHUf0N3mG/xSKti
xDpl6mcJER6DEYxCLw0wtK4JE5230O73vwIhEyxOI0QOsEHDF6QLCTIV4cMvQQqw
P6xuUICPDYm0HAFtLEIpMMBCOKpa/GD7yFigCt/sB6znhELrgXD1+vYrQv5Bt631
rvcDte1QhJmzdqSqZqf6DlWSQSyFk65mXakydbCDWzlmgKnzy6nQYyjf6D9oARSu
uvbQqwdjTuiOwft8ahYUedosNtdB0SmtJegCuFOtePsAaR7+vc8J9B4eAVkW9HTc
ioWTn2+vbNNqQWmPisgGQsMN+Y8g2MsPKwCK+/DCWiaoSAehUCU/Zt/FE7/ApIPN
dKNf6PUDYsla7CCT/dJrSa0MIGtp+45RxYNmfRNtjRnm5Ml2JwujONlJ4W2P1xcc
9Ujtzp70jeO8jlFkFrztCHoowFn75pYW7BYYHjTuuA7DEZf35jjh4BMOHPUBWjDR
7jpCZbu+sLiZ8SaKKL5Ab8xBUBZDj2MbgXWqxN5avgbGPhAipd+YmiytOzEu7Vnc
VOeuqlP8hdQGgnpAznr1QQ6gW4gScu8bDZ4gXOOozuS/lPajMqm3/Ge0gAhaA3WA
ThQ4iDVCcLjs7TjsSyx/8sD72xn02ilzJUORQ7agsLwSfwrEmqX8nfaJNCj6cvz6
iBHsWNHtalmg1JCkvaJ86KB3/od2zgaTMXBsXIu7U4Uykn4Jurtgw9+dnL6BNZS4
Cnse/7b6F1TyIy03YdeJ2GsynDPnKnrENlzoXP4zTTSF4y/HmYLaBOJzDKeTZ3JR
KpqwK2L4UxyEjd9HdNeutr/Bl+JbTY2nrKEOVEh6Hxnqsa6JWHK1ARYJKuTlEIQn
RSPSwVqqDwfZVxMF+jLIE7zsptv5osGES/rs9IunyNUQ5/tW+9+Bf2cJFWKTppAE
XBimXm2zzqg51K4lwmBtAg7oC0zxGVpf5SRxRkt7Q06i4hN4oamqSq6994mRjcDp
Qeg4dSJatfCdjpIJhTogipfIH0qarzRssQN5VtXqSiZtoLc3oxDP4YBLXyzZXG+m
Xg1lclhtyP2DS8feYW2CUJ0alda+sIWQRcylT8yDx39YzXXHByyBaqp8PQfzHr7Y
db3gCmo7PF9lviPAAmmlhHBjdHbTxZnL8hjndausTo+OKn+9fSQeC5C5OyYUCo2O
DCTNGaTaeqd8mg/2wjwj/4Pwg2GPNbJgfQKYM80YWYlsKuBViovoxXZPTfNDTJsx
rB4pfnZBCgnOop+sxG3IRbyE6tuJA/Hgyr7MdCMfJUXgBBXeOfqRHYLBHKcUtLt0
JI+6DcnCVt/cjY0BUdTIneWTmR/c0GkBdWpk1Erq+C5v17mwvsGLq7yajV8B7egq
onxpM50wdZttjKJqkRx9kcFTT1zFxVrk7GqvxCK33bDM/O433yESOnzn9KjRRGPJ
jyxC7OXfb5cosnodP7v6zV18Ko0JBUDVSssgA5ycPDI2mPn82zWOQajdwXqfndxV
BRkxuO0H6WIb64V9jTb9fkL/cULuUoj7wx25LlkCpKzX4YPTnLk7avg5w44SXc1q
7KE6gC63S0tDCT4LeiS44xB6xxehfHgMmYoQY8k3Vc9K0GtvRqKq6uJMLZ7vrd3k
96ZH5S9GSp2Qt5fgDT81yccyFMwvubmjRiKumGPuqfuW8VrSKyx2p4ch9kDVoD86
LIrNmfS7j4rsM/lGpyUFv/tzpxxRozpC8jy/9WRrQ+ZPemf/oPJnHunS5Rxhb1DJ
E/nM1G4d7RkgTIbhOCrOfc8I6QP6kVV+In1hRjA8pOwcYSua//BVU/tkQr3jU36z
Q6f5MgOkPrzaE1TySkNHk0FWqtSyOV0Fx6iVAXc+DVYqVd4wfaJtdlHiGDHYHWQT
poLyTnGQjrrC4nWBLjkkEPc6MVcL7Fw2jT++SLLHRAswFXVhVnmYLzqYsHs0GPKP
17MomNVP0G8/qDnN2tcV1iSGEJiAAFSQFN5E+usBrO/3JTGqlHrMjeRzbd7ODWDg
8x9Ht9SoAQny44IveI6Y+qDyS5xPsRi0D1c7crqSqx/yr+EiaW5l+6ByudJNJY15
e8IdeMEZx/u+d22ubApnshKKUtazk/Shx+k3dh7jTEX7wZex8eAlgk3xbqjxGdjw
vfttL1b71CmpYNpv4yV9vsB4znr7Kh+LZl/O+YOIigc1w6k5HMzSX9k/b1DvucwX
S6ZYEyyifGkKV+gy63PN+CRKBnEYNEdIZH4ZnfvKylOqlB2icuSuGNtxE58yr+Rg
Mz2SGszYQxnZlZRwwHn9ZsgO4tDuPf62BR5LaY1UzcJ6/715Uulwsc8n6XZChwCv
//P8VCeHWSc2WuO4Zsw/luVzEYVVF+pgL0ArNhTNfX29vwKpop6qbsUPkKUSgKPV
XwUf6EkHD+rgvZq1jOuUDHERZFcIguGBDrXFT+RGnvQ0myKE49P7CQTYF66udMSR
IpVDf7Sn70T/M3sZPmQL/6orFSRXWX9416j/ka8avQyF17IQp4Rvv14r4LPdnunv
moERU0yxMpdeT5+nocu8APqVljfq1QfIX6MlVJ1IT5SB4gfs8rUsKPv9WIwUQDIB
0iJWlHbN4h7ya+S/O/2w4kGQTtrwjRNGPfSZv++4tej+cbgNXGza26eD81t9R7En
WWTTHPyxqnKLj6KrXjgiL/BEFOiC4NDlo+anzNZVkU753K0ixlq5xeB2qHh1Icyx
8XXUVb0TfJpBG8AVfAAyDGe1zEyqZ2tMdBq3TjqooCd9a/+rkcZ4W8a+xLi3mJAj
ss3Mzk5XVHCZkHKn2OiX2ebJFGT4kvbFFPyLpWsMSrxHRGQXFa0su1daYsDVUACs
GOJTYfPF0WzskvOgV9l6LYQYJjnuPYHKoCKuRun5QRaZhfiNKv3SUm/ETX6gL/wV
/j83m0E/7FpCiym+aWizV3hwQx0sn5qDdJtmpWsJl8XWDASrvywxx9Ny0uGGl9o9
FLx3ia+8OU4Asof7e/kgQBG4SQoTMYhfF7JjOv/s+dkXyBKiAGjSXUyuY3DUIcqC
J4TFb0Cwv5Q03pvjlHDw2BkYioWB/2uAiH0gwA0Iue5+HArXNpH4cdPueWq91vY5
xQpVN245DB2AaXue2Q5k5JrpA3Gx0bdZSVrF1UnN68dVS9xmZTt70A59UBgwu/TV
Yw/nw5FRkyz7t/yjR86ggUrtHwzMp5z5orcOiFwkfTiyDjVCVMBye8+J8FbLhSsB
oaUBHHd2Fphamx00JyACneISUZ29nSovCDG2mnLqNjkB0SU/nMH4+dGytABrbthc
JYr8Cpsdi0p+hxp8LKkJwozFf7AaWxp4/O5Ew9abDC6X6/uM74cEYlLirCJlXKUT
0BxBFRB4LQ6USYlE5ApkSHgFI981sAodl6a8t12QUYEiGTgA+2jkzz1/ZsNKWMw7
st1ERmgFVtXUy7SX6tNqsWSlLLNMH6FCBgmBbUa+/mkGz6DRHHfREkl5ouTMhomK
aLf0wnM9D81QvvKfi1RcaRTl4zGQQRVCZijRe5B0/Ew/1FW180xDDxn3NB+qr15B
aWAVlIg9guq+en8QTjll7EDQvneOnbxUFZ/UsVbc07/xFyr6QmRvFXcqzFvvK+UI
I69yNnNQep5kBRPrpunDplk0jqqAqKDSXdoOW7h1ndIQOJn3/3hcLqcajgXg11bN
s9UVS5O9Bvc6F/tQ6w4C0uwj0ecgbZjTItScPlpCjvAGGTrozoISjVYDLLePiHlU
liLh0s/RD/iR7YenKoCaW4HtQujfxA5CCzcTr6y4HKOH347HFmwXkyc9fCWY9mXR
0iE4LRqVkfRkO8/ZxkFKvDuZMLNXZ9LtfiXU1qwMJfjEOxg/q/xED7NuM+SSfHon
r0LY/utRS6TBDyP5LfaZE9EFFaK5jHP25TMNY1aVOnPHhInnOw4sqv/s/+vBowTC
4aZMSPApWNrgsGHnp2/AmCspWPDRVVz832gkLJ5kHkgF2A+YyR0DFOyseSR7umYy
3DILkmPfk7rBj7JsGZBbCIYu9GEc/dUg1IxIXeyidKhz8SytYgzrovllTa/KXdvN
ijbCQnbVmGCKdr8IwXVWwy90KZjPEiGYjYHfa5PFRqvS7ftrv6Zn2VAU2AtiXkdC
wXPefdTm7Aw92FgVIqc6iYACLXM+h3H21OTjOLLMGzGzs0CZjKcRDMiEwgpR2i/7
TkArA9BOoQnyQrXuFoF7LBo+n6lq61oS5xUJMNTBWCJTLahBhCUiCiOdzP8kVndP
sqLaQQX2bk6AGhWnhjOGpFbUV9hRivLyCIUSSpj9ZOgHKVxWcqlrB8LEuTn7iLPU
jqmpQu3yaGEdY9NYGZfzqHH8a2idbrO+TdelH2P/29BIehDR7u+A2XATINF3D19C
9ZU/ycdYSvnWJIPVpHTvxii6koSmYBMS690LnjcAbVdyOcnUU19V0ONV4ys7qzYa
liXlZgFbQQXmgJBYsFDzQfUcDttdgAbACDD2wQYDUdhs9b0llghzdcClZRPIMTUw
e3UIt9KcclHlwH3EoCcPFd7It+pE9zJPa06OVRQ3Lyiq8ZLFtDeQ5c2hBXriidVF
Vtt3iiYrkENKUU/Zy2kji3uPb1Ljj6QQNxHNBCDSstiFKOeteZUP2BmHkDemy/WO
3FgqIE8Rg7pXNeB8qedHFtHYrNeulbzw4WfwrDshVKt8ajlBJwCt6cgRwaJDqsBh
I/GR+5KwL3Dgi6jgSwxis/ds884f+8mgf44sfCApiO4CXa3ScNAgDYRO8BphmOZu
xIf0uvHXVyvWX6HF7XivDeTGMgiBQ4J9hWwUDVzSccWgtO1hHs5cMsUBEHc/qAbX
gGsws7EocebUsTu8WLNDSYaLLaBD7iKwkz8NsagTVg7rns9dL2Ef7jf9qTLVOvh8
g3nUZjGQQ89FLsdwgmoeNLp+qqJKIHswWc3gf0cu92GYrX+1SGrrWroQ7XoQgQZu
CHXgDJavlpdIJygUjdJO6oahWIWLNRP1GTC7KmLZrpvxjbCcYdjushQ+g1Qg983f
VukTwEFoS5+PpGpJLQMrk08KPJd7WbCD3rCYxCY0hzdTbQ6sKLVGpwhZCqISOAEG
Z0592sxDZwAy+AiLEK53W5vpn74hpv+7yW8RYJGXBfbSlzDVyy+GbNhweQO2s+xo
j0gaDUUmcIvLYSF8qdLoD/8UM+Y+BMROFvB5EqlWbPU+sWYsOfVqc1uTEMYSRzNf
lVLA9LFbIE86CnrOsAG4pdbXL7DU+C1+0mzcAHJLZeUwIp03SfIs23+ELi6dtBKD
60LDEeizv+78csIkJUWAbvNFRKpImzJEQBaKsTaSzwNDa6Vr/UQazxqHumZDQLnY
/hNK2onFkoTgYLz1u2DOKlhDiy0IfhYiWYBZ/uFgyKxKIywW2wUhHdhuBsSVtoPz
Jmea79R1BT9cugA0u/BCUh8AP+G3E/+7ZNTzK/kdkXN9AtZDUnCcKZgahqbElwwl
/O84M1a8nUzN0ZMt63vGH90k2M4YtW+93teWoTFWxm1Y0pOuAHtAJMjmZ5CKa5bf
AK6/gZA9IjsMS7A821X6je+B63t4Nko5lO07mxCzk0ouARY6YnHLhfhLDVW0S0+6
fYgDNqMPKjWUrdm/f8zYQl/1mocYlb49pcw5iN/mK6K4DllAxWGpB5ZCzQCP4YCG
LUmRnCmpq+wkIJhRK91PRWjH/9k0ySG8qPOn/KBrpIalfKpDXEyv7QYSw0vEHWti
Qc6tpblni/Jkp6p4FxjAdx8KgJPZSImYJYSKMXENHAKqWffWPbcF69RDeabx2tF5
cKZNJmTFcWEou+nKJZu2jRLn3/nbD9x1FNiAtHf0FHxtmmB68J+zrUu4+dYbfGyh
XrbHjBOwykpVuPVb2w1FJ+4+PpbpTIIpKbXkppbhjr49A8bgRvAXeSR0uxB8AOPf
2vpaNSb8yBoIFxEefQdS0JKrt3JgQd5oOZx5gdOURiPRxLvjsy8P0p+fMAcRZVtG
YfHKjDKGgLooVIEYx4nuiJl9PF1XfHs/YCsr1WOqdMQ9gfw/CdoCyWSQUDOPNLzm
f+jKgidmOUkYb8fYruqHhg+LOZFyLJ71XS2nTsZYPpSZACBvdAgUVhJJBLdvCVDH
7d99c2I18X8WGzpfxva980huWkhPEBL4PTkp3QpOgiI8CRTmWmHYNVdCO6sd62zC
Pd/gMzPP+KQW1XnmrRgp4U1J2P+0e3i/qmTvmnLqVgd00AjKb+0GM2vOh9xRHDoi
6mIjNXRm/Mg2dq5mqja+tDhOn5JW01iKX4kFTZz+mcXchp0HOaZpCjMHL7/oz5O8
nf27JyJyDUYLsxDt6dBH+h/sX2VAjzlHUduZKXZiMd8FVjZGBtH9/COB2o84xx6A
15JPAZiSx9lRDCA/XmQkeSnjCP7ww3+z6HTUA/rjnwvWem5egwY+PpCHLefHsUG7
+kuQZIdbbky6qnBx9UZ6n+uTBrwGk9X4M6PmDnvDx0yv5exfl7X0yOyjSSTgX/ta
pIbD41wpAcQ7LNBZ7BFQADUPdMRWug2u15bS6WtcpYpS4VAJKymzqFcsSBq2cUbv
Q++iwtvitFKlbJj0x75zmSRE4nQB81fmxVmX3dQLfVP+7EV0hiLUrICec7HuPWqG
CJnmrUO6EJ0moXB3X8SeF2/REJ/fRtmqaquagxJbwMFB1AJdRF3wpjbu2ZiKKaOp
KX+pQ7XlDTETs4BCYPIEIfNbTlyLkE7kaJ7ZHxHePCH/xPnuTqKtxtFka8F2+3fX
pHUlJTlDCH9LuLxxzHEb82BoGIOeysZ8tL1QpmdhlOhI235fOkswkKFbxWq2/ro4
sHSGNbMjG4SAxOEmZ9QjMZloYiPz3rq0e2qSN6deO7yltlJhohDHCFKdAAld1JF8
IoMBq8FwAx3/87FlRiNq4ckTpmJNV5HL3Ebfx/WzZiI6NEqdI4WhGUj6Gky5K8lw
+0Bs4RjM/oaUtaMhgfUlxMXfXA5LUiCptOqM5tB/s3XZdK+UcJzph4G1a581coRY
GsF8a7E7lOfVR5fKisFYLrC/eDREJc7FXFv22zGuU/m6jB4+hDanwaEXOygeWQIv
x5ZwgAUF/ZqnUNGpE8PMzPhZVdeuo5NY01DlkDHtt8j02tzGtegcVtfqgQimcAg7
AfCbcvj1mAqnYZNZGNSGPyvF0YPuSYp7ShvRknel2BXQXx5BxElfBpkleuyuFnYQ
mCMfOd0roiv7Ih++gnyrj4Ozaco9xKnTh9yqG34BmG3LzFwtJK0DAoNJLEldiRT5
17Y7MsqocZOzyS/DAjfYu9S7Yoxw4Gi3r2NAVr3HwpmUZMpMgXUH07ZNk8ffPvUM
0zzl5mwfMRS8/dz6h3OQQ27QVF34RY2B37eCNIQd1ukJY/7+BLYorJ+VaYRn53rp
SA4pWQZzfiu3iU5HzTRYN0hBIAFWDpP8aJ5fJ+eJKKFUP4fIG1NNbVKCh47GoStn
guIFiwqAK+YMdVcsQZLPJGHzFhkyvZnrs08/YVtIXHTytVcm6+VLDjxsja1UMkDh
o8pSL80wFLytshazPzuN0sNXyKhSFiSNR9BjpH4DPcHREm66oaDdnXgKwsWCOvgU
Ma6yj1O3icoXhKK7AIbDG8XRw2XuXJ8fSywZmJRPD3yN0f9/TdGf91zrt9R2ZwmS
feIuu5qAuThwarYfaX1FGfNV8EbMm9A1BQuirGnC4f6bB8mX4O8j/xUkdEVSKFqD
2mWUzOfqQ3ZLObcTB04z6zkkI8vjAsvrX4FF8cec7ebV7y+kktjnHu3pZsWF2Wrv
AkcgydIiNL/JstSyGddzYkEIiIyqv5QETXJaZIL9As4LoHQ38CKYarkcGyh9MmEK
gPdcChJyToGu3/49WmlzY3Hkn/R36C7gVDqMB6OpehKIb7kRny7b+7fHZRCZwWyg
I9q+WndGL6abkbfaFH0HsRW6lwZ+j07VHpesTGA8ZRjNQpJolkP1iiZTRQqzMtCo
upFfjDS0eiutuYIE5FLb9s7O8a/AUtFFkP3/uQ0KOaPHPV/mc4cxgQKlM2MtyUVg
lh7ruLt5ytACn+ooluMHNWmvThwCHUf4FQYm/uUszc6U/LY3piRnsnnbggfi6cW6
Z8zAMgW8aRYV2oPuFxZWgduB1lU6UqRLlBwBoOlzP6mnFIthmrX2bmavd2OZ3jYo
SO5XkDIq3LvyL3AAt8Ru7noBHMkvRUH2ksGw+MYmLxVQZhAplER4ul4UOAOAaqiW
BpoXTMKONXO5xwkredU8o1uIP7CkEso0Brt7hOieg1jF1vYVUiq8rWzCHXOAI256
6S2BDCD+sWM0l8EoDbAb/6ydqeNcDpg1QNus20ISjlXREdi5+kpsIOb5etIiwScJ
AfdC1FAkPEXp5GCLimcEkQIpDI0t1sJK+N8zsJK2FHYmEa0Dn8gzcDS1N1uY5tqU
8MfHilSdkMkil+ksp5q0qnMz7TQgurkZAs6OctzNCGcMmex8RaWUR6UeBnnh5pkt
KZE8jgU/t5GDvrvk/VbKOGlQNpksMHcltPTDxMyxGef2epcq5jvBW6HwiA2v8wjf
RMVH1XvzUgq6+aZ/Dhh3ebZ4XPvyXAmpzUpUN3Sio4ntJnxkEdimhX6ci90ER5pK
uq4uUDyrKMaaKEVuMW1aCn0HLdZdGSI/fBGNnDR0jiPlLYYEN9iVOiujYrHLf88Y
1J95iZL3PCgvFDRNLXzBc5qNdAVLf/8ODLf9Z6/dgXuAmqarK5l3YY5WbN+aThCG
J2GhnkURl+LQROi36yWAprFJOm9azfJZE2U633/pEYJB7ZyPc7dHAPoJNDpnzmy+
2r359tSHrb2x947puJ+kAm47d05iYhnYftJf9ljOu5miWdZbDkUJIupYHMUj+mne
go4Hzemv4DukZuy05nDnPpGAofPBuNPfeIwR32r+tTeffjxC7AWfOhhGEpWXHYP7
NAYT7SbZm24tlhHN1Llg44uVJoqdEcH6Lm2TvlmfDQNTgkf5Uir+svcw1oM7UCot
rZU5t3qPLT/K5Wj5HEXx63T4tj3/PmJZBOOqRXw2s1+P3UYrMxXl3Y3GBKe65jwK
QhykBBgHWpioIp9OUkjBQYHHAHn3SxnIPSF676pJ95WR7KFjt/p1XxIzBf+owNtS
u1Aw8xaJoZajX0/BPGjnzsus7F+1EOqh5SdsL9DZJ/h6saB+Uwz+ZoKDtCUOg0AL
2NCRwDj5kfM7TQ3mllx1oWTQURPGJ/PM+d7Fd4q1dR8ONx54I+ouuUu0Z/r05FEq
B25xNauFiCHKhpGeYxNsrgiZKWN8IGxfPxt9A00D8DtykTzW3WdON0Acb+KKCULZ
CbA6hZbVBZTVrKGw0JEy0MXGzoO7gquKUyHlUL5E9Cc44zvKK4cH0L5yodYlgEOg
dO93856BLyxAZQ3BoWxiu7HaaxLy1EmPcKrBxvxUaVEJP2gAblVwpkMwpdb1DV0a
3/jg6tgQM0gx/yVPKAaV/UlNaNgzorn59no7jU5dx+iPWHpjiNlW7nGev4ym5JcU
bQgFQdESlTO/cxMJIabsUWMhULY9JrXdS93t0v07ZGDGGsnyP+wFEm/EqjAm5ZCP
Ha1r7/wK8Ps1XSmmrPa/oEJnoFqIOIk133PVcgmPa4xIkKVWDVAgTKYia48J+mkd
E/OgR2LKaq444X8Tne5zqdDUpgfL6H60UnaDfj0buyJRLsz66VyGcK/rk+++kCnC
byVo00M3EPoGBm7MOjB3Wp1ReoNk2qkKPNXIh2lliz7bbZvtJiJYe6GMk0Ec8MMX
dDvRPePQ3rPxrxrjHApmeU0Rdf+nl+2LOhxnOu7lBte9bbLA08ZmXFgNaGMdd+ZW
g/3v4MPpknBnTYc8IO1Zn8uprYzk/fxHH6tCm0Z038RAsiq5N0znKZ6NqLVRdkP/
AQkOT5RGVNqpHqQxQoB/h+M5j2VSYguhUDGdaugywoaKuSpG28DWAWfdLfmhsI35
U4pUR4Ezl4VcKtM3b7mjw6LLDyS9UsvbCw9/UIaCKSUXyr91nZCtPnW5tvK3Xh4a
FIJokTcUjvzIkmVgs4S/TnXUu99Tug4L4Qx49A36JlW8oqbSlQFC1Ja5CvPfT897
rXJIYOk1fokFupyhxlqmYyyUMzR8y6b+aP41Sfq6gdFxwZBHCKRPC4n7l25Xb81A
xQD/vIo+epoIuSSlBOBVQasJ6BCKTLoYVNd75O1dIZayW7fUwUlsm80h6LbiSvgE
auzIGXZfLH2BXTP2gd8pYtatzLkmoRNFme9OPBi3hCQUDHq9SdtvJTs5WCgVfcE+
aiX222CFTbi5rpODCSC/EH56pfDGlqwoQKOfH8OHOiO5VdTyJ4vmSsIOy5jACgnf
4Mc1f7ELD4DCtxV9GV9OA1ulxnDfEDKGG7MYdD0+XKKHyferuAGC0cr1z+Yw9Njp
UbTPQ0WciX3VTO1T9XbDHspt140aFNmiXK7mfiuRUZg2QAHwANwhHmamPOWHdbu7
pgFNhuPT63bZkF4VQMUZlhtC9LY1ApyHXy+q4PvgVYGq7A59Q5Mz0EQdgV5WkH7J
Cw/AgGp/UR4RngJYYMPoheQIcu/CPUvCfv9+/W5OXeEfZRHAA4c1xuGLOkELognP
Awqvr+bE09Kj6YOq4eOdLl1N7JtgVyeQ4okNGSj35iIwVGuFFvURAQtDD/aM+ghU
AjVRZzvlseV3VgS4J2G8Br4eccYQc3Jj2rzpPu8uCRpl90bXfWOLg6VZOhWnkP7f
lxtqoG91XU40H6d1DS+b4ii9VfG2kbq4uMmoYeKO4+qd/jlG9ASFkJdXFQXNNuz4
wp9roiKgNdq6ww2d4AOpkVKTjh1rO4eMwx0cQ9vqOkUQlVWFTZzwdCadLRObUunN
fc8nuTXbglatG/aq7WML8tzL3O7JMmrUgdkZ1ixWU4vzWB4GYNtUDslp4dim1Wkw
revaIusYi0eWoJWonqBifoLxnIn0yES0hI+FjLFjS3YGH1j7OHp1vvZXayONFB8e
scmLUunjsQ/vWKEo1qUnR28XUtCZ0loDaEHg4j/20ArLeamseiF1+TctZrKmyY5w
qzmfGGDZ1wcl4iEZBddahWzHL7fcvWOzFfIDcGeqcaw19hunnQsdxe7XRpxEc8m9
HfUjrvWFPNf2oQvp1IJbgOL8fw0Vwcewqrn5m5K7h8AvzO7uXgCo0npGF9dIBDCl
+v3wNdS2U46yuSRYy8pogCOMr2mQvY8RG+SZSfvBc+ziTx2f3YyldKtAVsRC9ANA
9KsmTdaOG9LK/9qjbd0vdOu459Mk2LSftg0nlcjRi9R0xZI+0YoQCs0UcHXO0vNX
vkyGn4QCFVPSgPuxI9u6v6MfUWAffhrkbzL3i/ig9hKrSk4nLXraaf8CffkZYpRn
TEgwDom5BVnwttmQn5tD5iAhMoSdnV7mCYUhPB+GunaF/fHfy/E6Z14D/7QrJlaC
jBW2AHn/UNuPPdkSbPu3lBqys+/L4I4bYdbNTs0u6VnBqnoqnlAylCyL835z8CDB
bhUow3P8hXviYfX3It/2hT2rpKhniNJrrzFSz4+JU9M9o//g9J3uWPXiq/j+bKdz
zO94Qbgm5aM5dDzsfmE4aHiPM5nPtoa82PSKR7mkIYnvSHUei7Cy72VrqpK0NtmH
7ntRM4p9RSBZWtZ8PjDKAZKu2qy8/5zusL4ddCp5HhkCJ26fY8IGRwsTUVwKYiHM
SZIXMiOy7dg8+YvFqlRXszHDAiWHMauWVtvGNblhtCjNrawjSJTc9bQZFk4dumLN
HuYNqocPtnVQJWPAQbdwn0x8HnvhMxFfyMbUbtpkwu2l11r2v5qs6xGI5lzsJs2h
lV0Mbr4HV23kwh5Zr/40aBeqJch0x3PyuR4rLXRGgm/Wjpg/bSP9SPJr527kmScf
o9454Wh2EsVvXLYOMKI9VZLUi13sCz8qdAQ1RkgME0QXtOZuyRNkpadK5N6xp/gc
l3jWRmNFOH8/ODBhzZLYcJwO8VsqebrTuTVZEmHJUOUlv3tkdvn48l/Ks9kBWcrs
t24MZ/M7klywzl3JkQSmDqCdKbrz7qTvL/1+DOP8lAlnh2+fy4NTuDEt9JcEoaNK
zjrJLfJ9P3DCbrNGK1J1S8O9sm/f0BCIcMWnc5HABfj33uaJHb49HlqLSSLbPee2
iEy464tOMLxUhyae1u88kib6g5MLyL4LZo1p93u/w3nLw4NuglQxryougXQtRr3V
5g9yH3vUWujY83w0pKbukstn/ghBLxswYxQ2CGl9lL+OLrYood76i55fkUX2PM4a
lVQNm15iXLeJLVZVPiUWbny42E2hlCcWWbUk4WirU2gQP9ynIc7D2FBE6W/0y1l+
7+fW4sisca55QsMMq5e+nNhBEmigixXfLDOEc06/ebMuO7MWHFQUStesvgkLS1Vw
cJ679vPC58UhZttW2iD6ROtKPU+p7kMFgsinai0FsUyPu0mQrYpzoUFHLTbCzj5x
bLDKg1VGsyqQTxS1gyE4cJUu9bakag8pKf0Pk08aEfdM7hni9pjFEj6J/YuZnGRh
ZoVPHJvE8go02SshOCFnMMFKjoJXGc/BQTiB4O51rMePS72G5UL+3uvxnJXHNXml
3ArsaTzpmrqB45ekdzhloZluHx9fKgZFzWHB5BCKdba9rwV7qAOU5jEmYXe9A6rb
gBh84AxGv4AH2d/dqRYjZZDm3U+5lSGGsZQSMsagPr88iIXLA9scTdcIJGutm1u6
R2CE5cpbIgXpwqcg5v6uQ9wzoAbqFq/G0GC1TOG77fOIAwRSy/Tk9pjODm7JmDiY
2F8IzTNgMqhJsnTDCmfVWEDD3gArJwf0+6JciG01aoKOaLYAgTVfKeMzuy0D7JWh
qDwjx4XQ2LTsusKyUcq6W4ExZnhk8iFic2b3cwL4zRWqnxR+/D4CRTmOjwMsLPTh
aZSCIUO10g3oJ8c97a1CGMAnFYpD1hzxvvmZN4KE+CZsmYczqhyzjsKNjPCcLFlV
lnMyn+iVNAAPN0MSntVI9Rbrh1lKLVxisIA88Z87GKHw70vm4E1UlSBRYw6ryhYY
NTS2+uGPG6CdhThY09vW+SjTObfY9HRI3RLQj2iPq/rBX+MEqReglEnn3XgF/bQB
P2HPOCp8/QVG38C7uarKKZHO+y+ZDcChsjqWeTEAaKR1G/gZwA7iHYoFIQc+24HV
H4awqf/d8Ydg2N0k7xEUURZmBIIsO2LOOmVKS996txV5C8mryh4TkQG4cIbNJqJS
hZVFA7v8K3G618Xbsv+/mRVdbwAFRw284umnguYGp+Qs95u5vwNSG/44NfFeOpSR
md2NxKmeAezAlhddLoCv9GG27xcb3Ai6zxwmZP/OSTdYYT1Utl7sCxoHgqNzt4gp
Pljw7JqXbd7qsQJ0s5XpzwJD0t1iDYgQ+C7wjYC9RK1w4iK76sYlqgr1aU8gKQDM
4VzDveNX3PRnwsM/QXj2sKZcS4cX3INnCa0Ggp2B/00dRozoA/jO8YQIh2CxRBDy
mCntxutgWgnWp4aEgheDNNxTbc9f02kU61sSoH8kNFiLn5M1y+ymXJCBhmHkDK7g
8Yhb2M8sz8YvALKyeSoVKrHQebLy2/UD7AzpPYnbsSM0SFAb1kg3ZQU7vhC7pUVL
wwKPNFTlWegGxCbyBh6VmBrIP9p8i+dL48iTD3Auxw30xua0TiS1JhFb3TQFDG3g
D6FRZYNhpFeEuiqyroLYeLJQNCIfnvQ1cI5QQgfqg3hlKBNjJf9ToJSnjFZpgl8L
LY0fZd1eXxFKJIUZvoAIHxRs8zTwAyP0w/QFoLt4yTFPOX/CJNpYbEuQ3PstEG6x
dWcEpo/jPerh+oqXvvVUNsPkxU5kEoVoiM9jGJ/XX47OW3p/qOX7dslwXEzPUr4l
DlqJcCE5J7K76s92Vsyr3Cca/tmjlUsXFwbc/8YYTbCskwAJVnTMhdDo6PJVMHd/
YmoNhuoVPk3YgglDNtSjp+n/usnX6jnhU1C8/LT+O+OOmecs1OlbrABpaeaTuj06
3zbB5SqQtNWp9zDQf9ua55WZLFWI20oBoyIjdske586tseMaMo/1luGLc0GaewYl
oKScD/GrxNOjghLunBowWEqzJMfh2q4ObhwnSiOKTIiqd6pmDKdtlM9XxghjU4WK
UwEjxqJxWLmzBXWs1OARaC4JJdmQjx29KoOHs6gs6CmzfBvnSkhQDhyB5qkTW11L
FB9s7Mz1dgVBECxFO8oactYGwCpluX1UCSW3hk4UDPKzor8YOeO5eHRBnp4PlqL1
r3JGPPc1h83VSPMXf091pfpbw51Ge65wc2y1pNfbYyBJceZBf6q2LffXFQwizk3u
pxAZsrL6cGW/COLnQ+OTV1SSjuPaXi7C82bMPVCW0PTCd6QjYnFVjEbLyDSlJ6s0
EHxluS4MyMbElwoNSjwZHBg6uRJzlc83FE7NiXNWP/QIIv1LxDoBBA2frH4R8yPK
pIfPZNGzIFfRwL5szO8/oOz7YlZRm2y4xMBPTxCt8jjek3wCEpjYPxfzmGmjCcFB
ecWZBYTOVtHyHMhC3wucq5F55JLE8fcQsuUnr/qZgLwKNSnn+i3PAp4oSqCeGD3D
jt+9hmAxPB5wkogFOK88GykXjwB1CyV24phBOcPqUZatgqoIaxUD5XEbfxV3fm0U
HKt32eBJV9RX9lvYB7QWuiQIbV5xobdaSGXK6+b9tEeB95+rTyzwWijQGj2370GJ
Ug3rZBJepME1d9BpmOgK9z4NlDCau0L3ejwQXK15lMoT8OEYRr8jhoRcOuoDCdh5
hAV7WySLCpyYCz3V5Vm4R1uClgu27DZn6eXXj9USG2G4AyfdkGrw2yJxIlIt6zDr
NuNDiphiw9wq2iF5hAX7bSmbz+VnG73zj63gkXFxJ7HBExBdaGHa5b1j7DhRCKHn
1qI8e2RqQPUvp1a5f7ZGH64ZH/o1hUoB3sBa6XnHnN2uzd9sFScirN4J9TGsO3m4
OGoCkCmOJKOAR081WSlsPACEiRVuN7B9D9EQYCqcY6pH5yAE7tNJdgzNscCrHUe+
DSa9yg2pf6axwhXPsFXUMFilGn0EH8yrQAHYOwiMPMTCsfBsSrgy22OV7dHJ6pQV
3VN/W+MN5ygjugPPE/tY4F9UbNepmEpeBZdYw7UxwTea8buz+vCgN3pk7Nqod+LO
YKlSp4nIUEpBKdNddU1RC1TKEGLbkS3Hs29IEJZ6CBjLOduE5Mn+4MYJlcVtZDtw
lUHFyeCNpGC/JNxt9iByZySuo3rHrV34RgE3L7dIYJRvqupWw1y5Qo6mqK15th4X
3imL5tNj1IhXbp/EbwgxHh3EI1vWXEnDESP56mT1t3dAeuPlz1iq7L2wQBYdsHc8
Vy5YxLTaMIXR9iVfzSgHgvJpTTGlMhIkokI834pYBvF2/WyrXGjSnxs7Llpa/L4s
4Oi9IsFDEejoAPXdwXbIJjh3jeqQVPgYXsgSrqk+Bf5Qj0KPj9Jh15Wc5m8Phxe4
ct8ldiq/Zw2dn++T0vrwoy0pM0AIVi4RWjMZS484D5JVYGpmoKs8saZyg8Jy/e/P
3WlPKEDwvDa2drCORP9WcRmJD36nurJYOdNVeDrqXDa9PhJvpN/fEshlF9qd0CBw
MOO4nD0Icvi1gb9EUQeZtNHeGNZMWuOfz/sqN0AcunbUp2CP9Vc1bTUDpXrQok39
9j9fzDkhH89GVvSpKh0SPjE02VZ3MVk/vqMgeejoMNnxGNv7e1B/fPS4MvvnlGQg
u5ANa6EiE+vjCXbNCu+p2Kh5qn2aYOyuLMcuhDTdvisu9fybUaVLIIk64UIRklu4
9S5XioVtZDWMVQHEGEeGRFjq46MuBmuHogLlz6T/vXbhwbBztfcux+FGd3vQqnuD
Fp2ytU3cRTd4XKqlARg/F4H4ajVkbggcXaAltYR1M4y8oi7wqMfyvbr3d84eH9NE
KHSr+2h6GOTVKiZ7XlMKbWVQQ7+hPMoPSTKPqNNsOKiCTqQ8B8Fwv7NioP+nQwLP
uCOTMfhqGVJCL9gHbsOqwAk0L/Ejnays1SSDdQCI0N5JSWKHjckGhGzkaV64OGhe
FoLHTzTzWzi0mAVD1/NWHqo++GTIMQzSC4+dK9NRFTKumlIaAqTEEebP9i2ir80x
UiRXn09FHd0AWhRT5FyZnVm651/y7VQ6H3YQSIv9Anoe82yX+dfT+hlUFaltRt1n
sxIisszQPITqBKCeGLMOLVXSFMrwJnmuROv8FoUXNruhbOsZSI8dr/IxIqN/Yafb
tUT8qHVao7YZfnZotNn0T/wtwpAlPHz/EIhlvjBOcY/VQzsZNC1jI2cId62l1wY8
JmApDu2DVV9HjkqiBkvdREJVZtglU9yXe/Xb/66wldhZj+ehIYazpKSHpSOy3Eit
802A9bf71abRE6bLetJ0XSmYbF624QLsMrIL8un8EyTVmXubI+StvSVDmiKsBScx
/gRCjNlJ18pF3l02JnrTHG4Zjrt9PylvkkUywHMjzLGPqcvWiVxum9+iqpztsQ09
b9A6gqBJ6UeKEAK58xNZ2bilDSi39Ys8sFv8eIju1aJHnbc5IH+Ihyp7U6uXdf07
mpwCJH8nxWcJ59QtVf/iToBtE8XRvxmrqiDiVRAM3uMbzBA5ibjadGaLls9uAN9D
3AdrdIw4NVkQWmXRoUPdxnGR/qsu85elkRaoQ1+7gYgG2IX1LTC2UR0q6wHfyLRv
BQVAAmWvoXKXPwfAFWgZ5IRfhl1305UhFs7FGZ3bPKnb8S7AEhZCNF8DEPSktK26
WsBV5gNfU2aoSjDmlZQ/0Fdmyet72i+KU4sYQYyiTqZlITRO8PJglQc1lAhgaTap
dv8Mlz47oCHU4fyYfbpLEct4pvEo//BFL9ZCunTX+jl9JE2E6U7v6BUgr+pAiX3D
Z5TGQLN4ntzi/6RYQ/yRM/bAZeW9RYVjo0Q/pFPMslWdkbYDUU4GuAz8m5KZdZho
5kiHvWoDtTi1y3k2qQtICvRoVXUIIUzN8Oihx/e+Opykq114wPwSlwjkL0kT+Txr
8SDEQABoJO9MxHqzNyQgiBCEJMhAHjyMw8W1/K7z97Yk/Ah9BBaxadifo8GXHMe8
U05Tr7q5gC5qYjh+nzBokv8uMVRNbgebTFiFAbGLi+VXHlyfLxzucu/9JaDRQ07t
jIdhj8iyjnIawPNo/m7KkUq5raFbaeONyX+488rsJUiC0awCpkgavSuIifmgmATk
PIMj7vmT1Di106uZOdTE1bsAgUTFLjHp1nbpedbj93d3aJByjkojIaZZpfvx6TBT
nsa3bdwW3c5js3lu8TgHGqlW3S2brBzs8I1o/7yI1Vv0d7IjqljuSNyUaKz6vfRD
pTrHtjJh1CajvchKqUqIozy1CBWusxodLESykbO70Hia8ouadtiBk/XqVOx905NG
AAYPuUmBfDAGHrr24d/9wYy43/Bk1F0YzpWh1sBDVmQsL+JKcW+nEaAEcJffSjKu
KRCUtT5Y7cg+SDSjXUVJO+3JTqeYdzwfc1I4OUv4eKc6amsNJglvyzLM30dbs/Fl
cF6NsFHh8YsDU2CcXOVnbhruH3UDI7nh72OFz1cNcZFH4WXT8kzKjqMZa2eba56I
2AwKXcueGxdNvYRU6Nfe7MAoL7mUWk4tvIawvuKkVeIDViBLCroEHiARYUuMiijK
a99jEiG62QVNu3xs1qTMrA3WgnuT7nydQANbGHlOS0Mq8VThpVGL8vIyDOZU45Ef
rsPRVDIZUprFwXCPBdc+uAwof/4tNMcIIlT4JESvGYWDmGI9SVDiDOHRazFfmfcP
TGobKlzLvjM86FWRmOBQfHiHyygSB/Va7Kt6oQGXFL8dWRNDy4JK/6ne5kODSlXC
Kf0FvP6SL5EaCf85NBkufO2IWDmBiaN2qoNgVymvhRFGEbHQkG9O3furNKyOOESm
cpkT2vOeAQyNBUU/4a0EMcmrE0bhGPmWrf94Ny/sB44SU5n+ZEiLqEEMaJKfwOGj
kjZpRtF0dS2OeAtMb0Drm6Hpf8bNvSl29OMFInOHfUygZ+YfupxORNi7iuauQK5O
i17uHkSO3B0EBtlxYQSuXcx0FXButsKdxAfvGEcY8hOSflndDHSEXvws6GOVxUKS
hiBmldPUH67V207CanM4RhGwn8YhcMpguz4NXPuPTcEyo8HOjEnvFxeMZd8gKjg0
NfpzNu7DlviEaMpcXt5sJUaTKG9tU/1sTLv4Pzwe6ZDrmVW9byUQWkBmjTUqyNrn
iPN9cOHkrGT7v0iGNr6HZDHEB/YG/kIuO/LRIrvOxIgr6sA/SSigChP+c7YHpi1L
pbSsdxckfLkESMU+dw/weu7E8fISN8b4S4h9j+8mlhhq7zUODsLv6xr7x7CusUbb
59wEbKT+ezwy9ujnUH8bojAQ8O/kzKnCeC8vVG/LVooVPFe6AxNqor1okEZ8NGxH
0qvxLF/Ip/XxTIK2tSAgvu9r52wXdnxckk86qauljDFq4XDb66VRFR8eqQj/oGzO
zOXD7t/yY2hBfnatBesIf0Lku4CvQACZ/RFDbwOmb/9h3c4tM0pofGn2+cVTjyUp
kFbVrxx4bAamrzfIeIdRxWLYySRe+hfZSqAujOWeAnKMLq4BCXS35tcjmiZqAY8X
2WkFuzEHAd7MkDiC5cvcYeM8Z0OqlZCmDVxM8r8VG6wTYba6ErG9q+3+3dvVSlkf
gNuvCaOx7t+ys213HtCUDerj0qjPeHjmHLUAgcHPP9lhb03iR7fWPwu03L3od9cE
Q23O6OasQa/vn7NasdDg1X9yZ/mi53qmyk/3kY+uvQWsUTodnUC2gGJCBUyvxvKU
WS0LjLTfe2A57UQRx+7krapklcBHziuZUK5XnH9EmdeW6NgYdjJAa1PYk8kADmJF
QSWyXPq1TC1TA1Fn8wxN0eRWcmn5/jy/Sw9vb1+JAIv5lbGwTQBgv/geJIgAliZJ
5vvmNmg49DC/W7RA4PC4rSPGWXItfkyZiFoHswFkob9Y/KfBHWIvJX+SuTnVrg/Z
AR2QHc73nUjdHcrYedqzQc5pG4mX2xVviEBbD3niEYU2VEe63YyCxbV9iNz+El82
kiVbtWCrTgdrmkzIXGaRvOpvwSnyUGZyjKNld1ICg5g5g5BPe9KrFpLY2H4k6bNc
xIjR1nHQQOkou+AwtG/QYbKTzVU1oRrvOPFmw3N6e578Cjik3gVYXn/NzkG8MOyV
gZDsYpB7yI/+94ciXwDszZ1UkyQ8SQcjmuqLt3uHG3/xoaXYcOPhkWKn2qcmejpS
iAoPXNUTAfqNRl4QSt3Hz8jAt8WDVnueFXnOZg/2TQDI3CT48tziMVLXff4VIuVZ
9BbTwZv8SdOMnv8n1ffeKwVosAoSEdZ/F77sShmwPeskJOVmgW4lNp8rLmKxNgkC
AU1TWEhfdcKRdmRymPf1zNrze8iJquUaBJIYpEuscns5BkYwG9D5bdfEbKH9enMs
rifJCti7wVVIiMTjmY99Z1q6xEvnRYhxLg2DdzSZIGRc30/v2Rcxo2vdg3pfMU7W
vQA58KXk2DPIXxDM8qGb4gKR5FyYK0MZvf1ZJDJpO1kQ/7sj4eYvX6m9gLs/ORdf
p0+i40leO8K3PTeZHCxKMB0WXHhD80RFqRY/xPHAOl1t76GFhKcV4bDND/aVh4IM
biieXeKLlhUwRyhqV25vUqMLTFt3CJPsQ6/UnPSBKSe+9NWUWdmE17ol1DDDEenT
FG+w504pHFUlyvcpBHT7Kn60BtT68d41laP9/4PrxfP71lYUobmHlGFQa3DTAz/y
hbiGSYjnU9+HPtSuopYh/nhkm9YgNjJ3ijUVJ4e38mhStGRO09Ra/uPsiDQoOnqS
rfXkvSiLlcgTvyPqh0C0BthkMAg55TGvCFIvT5xkqwrMGbszov4kpkTSwxplz23l
OYaqnZXwGXu/t76aE+2taZStcVLfbGoK0qMzM8NvykCmbrk9sMRLVtzvBdCvjkbs
10T8t8j477XIyeB8P6CHcqrm6MWWnWMji8L91TahNz9lvkGuDtpXZidz4mFEBfMB
+EeWwAZtcksurGjS3hgVI5sGgzFhynNQyQiCnc+WZ2toEoG/sv80afUxT7nqjvbj
AIZpkNqZsbHemio7WDH/x40TIbMjfWeYEqYvZzFGyjtdRcah02y+wzAU4XqG2q7D
x6dwVox6rxFZE3GEC0oK0XjKXD9eq0huPbq4SCd1q7kRx7FWNRpt+PALwptH1GWd
DAhy6uuhHYyC/D0siRxLkvuqninE9R9qh1zKafR60UFwIpQ3zu6WQS0NCtiuL3Pu
VHIXyCzAmD5wNgvBpPf0m3YeLKZO1E2iplgvqFfK9qhZuxPnCgWQ7SOtwgoKmVR3
Pp9p1CHgHB3fMi+H/ha6tnrDpyCTuck9bbF+AxbxT/a3y+Owyf+rIb2AoK1kM64G
gJPKtdhU9hY10yH2t+m4OAbGbYktXaJk8m7L7KhU5Yr/h6KceF4mMmK5In0L84xI
Tgh//06iOUy+x3CXngvlfKP87mwgr/C21ZWmE8ltjzJTuUs7GOiXZ0UxmP1P2JDX
QbzoEiia5fpvRQt0g2xUeL38n3lJSy3jgAFqJxHBOjhzbYyYlK8zCPwSUZYKYZLZ
lHr6Wi6VLVu3nVFYFZVpMoAq2DjnS0ByBOO9uKtfPVVEmxOKkgTfZGQHPJKcSYUg
K7pkdmgEVl/ujHymm0bUGx5RlSepOCscosmUmt/s7vcNG14qz5ezCScaB8zGSWN5
UiQs2Fxgf+yTxqugITiHF6Xt4s1k1mV67WW0cF1N8taclxVF0sGbu5ScBpCHd7U7
mJRycO6z2ilW/FdeUVsSttC/OWwr2HJg6LL/9yZzmx1bq5M9m2du+IcOp6sr0UEI
6lmq6wLO8rkh+80YwEnBRG1bEHzZ94pw42Xtg5Js66Y71Oc5yGUtb5UDx4ZTgNC7
JovCyITHGOD8p6A9JzI0XkcjjxjkH8j8HNdH/UxsseU9lHBnrSq4CK8ZSX1DzJ8I
XmusJJUH5objEe25Kj4evgKve7DXZ5ifYJOPieuxLjCYFplhX/t7gzf0cxDfRDpf
TK7aHpJ5HDOUG7t7hu8wb22y0TEeiPFvJ1RcfgMJeTUVhHLAzrar0uSR0tBFQxdB
eUFfPQ1cX9xQosjWXg+IgVyTDR3edZzQTAgnAXV/w1eCNvFxp6YVxKBRwYNMsVCR
Ejf1qyvR9z8OBU5Op0tt44FNeR/zzo5e8o4kjUXa8StI0Ks0dslylDVhvJ/wBt/R
irpNLr8F4VSPbMfcVxyN0/V1FrWNI+rb3bgD6wu4CobpbaKbhLH0Ls5ccDd/O+Y4
s/Oc3f9I+faj2HO8DBaYhwZZC08PRVs8GMSbICgaYlblvd6GLQ9XXc0+WKyhiYg6
h7hMafM2DZey9i0LK+UWPpdEhowsL8D0NQ3m2956UXiJesHMiDzLB945VixkXooI
FPDayWQyrOGVML6cfqidqW7f8w8qvVCqpeSGrpi2gU9tZegM/wATfWxoAh962Qgx
Jcwr2Gq90sejlMQOLBEeiS5JJz3PN6xyiZ0dveu3YJwEOPXjxZ/orzwsFJ4slOVa
T/fe9BvMrPUaOfR5bz7tgzflMY5M9TM2B6XrL7N57eoYG2p6mM5CUcaOpcvGwws2
wxLWjNnPnyFVxS3xqGCmiP77BZjln+0skfd9nkK1GMuyZns+YhiqgrFvc8DfKdis
Gzn4Zwx2cuStUEASL8iC14egFH+SGL2sH6CMu+iDajl+50G73GxYkKNVz/rSfN+y
h90CO/IkVT61+IwqlgMPwhrB2G04U34HtOK+30VOWwpzebuC9RKXJJjfFmIkGyDk
5GQUGkQVK9VeqxP/msk83Jf6RQiSDfNyRZ6ETRiarmQa1Kax4iHqgD2+HvXac+ev
nLJFdr4GHGq4rU6WD0coy58EhEPIMsVOZWALWim2+P0WD2Acs3hemKgqyP0uhBD5
9RZwQbS8PRYfYvG1yIwlE+3xaJJ53bZjeEVlzzj42uwynk6v2HUsbtLO4ke4ygTG
XY45zU+ZQ+qNKazrGo9SyVIazIKCLIfHZRSOhKtJ3gBg5a5ATpeo8Evc/RPnlG/G
/obCzwiG2aajud2AL8SUVGE6VPrzWtmPw8dbDeSOOtKs/ZVgajCCtgVXzMFswl3W
Z8VgCQ0Rkfg7uKRFK79PmglzmCdL1iNK3MbuSNDu3/4c8DJyQAARSfCyYA9RBJpx
r3Vx4DG+KYEiFjm+7jOrZYg6AIzosmV7a+mkYDq9IMAkVYGiTQa3n54dB5fM4xHI
fFu9QVWG2uOyzUG3cpinAFFfM4NdwfCsrr9i6nCCraV6cMmnFBP476S0pPout1fh
6KWqayJLB4umvkw+ZOX0xyOceDM5c7dezgSpBS7QS1tMcL82GHLPz4jmU9VQdUSp
vTe4sZ2qqFo8FbwSxKhZU+CgIfYXxoXBXlpTqIWTGmKa7AeyVuUzvZPt/rZZB8Hk
05JeyHfw0YMUffAZNKskyt22ldbzcU4g68atF3hmenzhcFTZmizPCDuELj0vMrcb
oFBHED5a1AR8L0HTTKDnGRbDWc/jRF3YtFAFwa4Rb/FjI1MVkD0au08GBcB95OVH
XhVSgJEEHOLWSBFjvQzC5AFd/0IpUzjg+8Pqsp0t18PZyOXD0h1YXDFa5Bf0VEyX
u4wSEldcQlnl1eHoKN0HfyZIb3EZTxodjlGT2jiVJivk06PY1PVlrGr3Vz7cosfT
ALEsk5J4T84BPrGkaBp6ZH+yfRTfHGvixkm5pVfboNTH2m0aQQQKNxsdzXGaRyzF
AqnN3TG98SRdb2TBgGPDUa3C69m7r97EYMFwksbUQa9GO4a/QLLd2hlyybQ3IROz
ynlN+5vcRtJ+IMLKcfjDrlA1NgaoYcRzX6wDyQkCvR01Y/ZkQd+Ya2c8naHmS9Ds
ZRl24d1G2ATU0p9IxG770/WYdJ4ANqH80KBtgkjqVuiYxWfxenKrfXRocHXBamsY
q7TlgTw7qlSSz3OcqWuWizMQKWLZK7mqh9HMyV35zjH8iFIHyPnUTQUt0gByczYU
Ffj+9yKtEhm8QbUNp42d7fo2WVQvKT5wNHUQzHV9ofRneaaewJNWl9uhV3ghTa0d
k941LZFefeSWp623VbPTqKKPs29qazqAceyAxAI3cEo9unbXqc9z+HkgOoEuCsYd
NG2N3KbXfqz4Ynp4QpTRSUXF4q0KcQvTyKLlplYopcX8g3AkRo4pPjvLJ9t4+RBE
AsOd/qAsAECITKuOQv2nQD9X7gI9oPs1o9awkHZYw/mby4S3AjsPk+TCg5sbCdC9
pspdov7NkbBQFBI2vNu5FRgjPP7zlaIbtRQLifdoEoaFzHNcZ8CjMWDDBOhI6bMj
XhVHLOwzXFEXV5rTjYvPbvxiTe0izouGHSO7vwznEI7lKv5s4oVyWuKDbyU4X/Q1
VirrZCmpAch9kl3bfeZa7zm78ZtbPiB0XeHUWbTL5OgocDLLKzvh/u1TElTEMg+q
jEB2Xr7OcKplPnGUopMjI+0V0T09Z8AsuHycXmAERg1x2mQeBcqHnoqn9+jMA+DY
BJ2gVzaOT8in7h9X6cMSw6cemCGg/dBYek0rRF7Ty0dV4WI7Mda7XRQKFo3veZw0
Jllg8xNLUeX8aQGlGU364JY/5NZuQfR/cf/eUKljWiy01yUzxPtCw065TlED2Zwu
m8wjx2EWHqh4r9n/1yIR5QlRVOJJHNJ1q79KS7gcmZmxTBfwy5GVcp1ykdz/lFFH
Y6HgozpNz+/i7z/l0Z8+06j2MhOkRpLruANBuoxc9AZK5lFN0iuvU6QfYgyYukUs
jqZldsXagUPxSueMI+D/B7s9aJrEWd4/TBtgmIfYxCN2yl9rlNv0rVt0fCOFcbKX
sH7LgK8as/XXQ/KjlqW2//6ZFQ7jGM2bYKGiXJT+PpHk1IFBTjkbdGymi/OzYPS5
1Y9VPrg4nfzTfMbm4U0u7utI505jqYZdEWwY+bN+5vujACHOfNLLWJ38Xx31s9Dv
ZDzegR4YpVXrnCCPGi9htylhoMGKHe0Ko4vIEWO7S8FZo1hTEz20wEmfKClapXIE
ltzlWC7dXFmdccAuWnQin4IKGMXKGp6SS1ZENhtOg8YBmBat4pE+yRV0bMDuZYNy
I30//b0tiZs7C61AbKlADpNvWb71YkjBeaML40PLyGjQU3sq79RcYsAcVErq9KPP
kA40prupybwhAzvHlzKNMB9r1a/KpI6AskKIrwNtvez4B395JbhLJAlZv7xXkSzN
BdhL08wITqTT4KBggJ87oHjOs0B/FXFMO0HXNZW0ZwHanHsCCGVgk2uXXD7Qsv6B
aGh7sa98HQDCuKDtX17WcuooyHQYx+JKHFrkaky9w1S8C4RgFGoN1K3+7tef4FAG
lqnsmeiepObFE5HCyb0+/rEy2epjE4Oho6jSoQGWNXvAJXKKdFvIgn+lJZiJMav6
zOBQ/1IcaRjbYZuQNt/JlIqpbhdrJIoI+rqlp9QPFtoW4mBEJ27zWGr3DoYE2+sZ
B47fMxVjSAY8rT2gu39ztAtBKhnKv5gIxxwFJk1WPWK4bw1CT8mQEoUnZZq0xjjo
sMBlhVhGdNjy+J6Q2g4XkJu/4gcsuFhk32hX7eLa9X5JXx9aEkGOm8m3bIc2HcMD
+ld83qxrNSWwjhX1En3kcM9Mh3pHZtpa7uyVMqn5CRT4Fael5NctgbqKvc1RaAf+
UukH3b6RYBy2SvDoKvHGzI4oZ2cRq2idc3iBsMba2G5bTTNrRQuFFYHknugVKf5y
GyfosWFR2Prd2xLToGfG4STB4rK+ZAXrF48pMJegFYkHtvtK1r5MVmRjufUznEeQ
c/3YK7zT1bKQDyM/DNGZ34ko9NxYltWGGL0RC7EXZkAIXYHFcO3/lmMMsePuYbW1
QQvHsKoplGW47RSFmplv6SUo92Kr/lziFoyURenCdyNHmgYsyjQ3SPMat9RoPvKc
0hRib3POuUlMra1g3zfNVG8zQriKYvic0sfJdI7vNTuAbhg20GKrra87aAj4WnOd
FhQp5/VCGXWF0jR+r9yAvTbO78ZkuWDf1GxtucT59axqTOXN2WKMMNoiBSZoxfTR
qIZY6DRPSPH7xVSra6IxoUUXmD/AVwCXlYothulx6S6As0Z7TOcaBtlCZwXl3jk/
aBneSrfuAUQmp4bt4Zy+Qz+beHzsGAAJb67F/KXN7HeHJJtQEOdGB+LfaZsRXI13
ph6V3/HFLmfDbyobvlF/p1HIHxWsN9WqR4JJkV1RXCEmjv/OhFWtcI0oL0QlNzzY
HT8FfpezeO+oT3tVswrpASuwduGmVf5S5tGIDDKXhCOVmVXtppyuOxLNUza2sNGF
4O9YC8bexqN5yEh8Hrpl4E/nv4MmqNfoRED4OJeXBRBT/slgtM3rv+BR4A+wqEy8
QcriVjD/hLRfT4tfGuzFHzROzbdZuqe2YWNQQnAAu8NihVpz2M6yVzSDueN8vtP6
T4wwz1KLgQrND3Dvzbe9SbwAGwqiJrDbkRpX91ttEti6UAKvzK6EyRR+CM7QkPno
0xsQCiUbz2j3AYXVOrGNbL1HEeYWjqfI14iZi6DkipbH7U0ahbLKMTh+B0Dv6Ybk
zQ/3EmygFcMniZwlynpLlFTGIYm7t/de5U0SU5I7u2YREPkr9plE33kEHr6IXX95
MJ785PsdWaWS58wt+dHeDx2k8JCjexQkob/wr43tsjsh1+l4KJUSyAIE/xOybGeH
/AHlb1ildSqFIahKstMJ7oRVUao+kJafccEwHM6xxM7BZC2uiiP7UpyuXU6IHFv5
z+0EbOfzXO1jY+dygFo+x6UX91Ncfs28dThjRlsqnYkdQX65imj2lKZKZVwiXonh
4sFe3iBFkBaMCRtTtbLz/9bMoK+YumbFX5fJoDH1hmGZWSyRtKjvZ2kxk6Wfh+b+
s8FVaPQB5UToC/DjHv5de7uSEJMqs9Bp3PEXTUAB22nYOohySV2dD/GtDmZNRWsa
0J5MO0xRoM6Q39x+88zNF2aS6nGvCglVfsy5Kty/vLpypuu3xCFP+JQi8bkpbj3T
bbuYdHd6YdynNk0WwwfKT5EFEfepcBd/i6+Ecl3C5nIfIDZGtPc0I4XemlvLKpPM
+2Q8nrAbzh8Id3VelQiuozEY5AB22erXPxUE+DrxcTfH+nbf/uwEK+A86TR75ZvL
gK1/JWC1b56t+bhO/oXt8DUv5YqoQ+ErV0mdJ+nyJ78dPSj5QVGMdtKkCd0cdAbG
fTbryeTjGY1T8jLNqRkF7XZOZheclOIZdjEtTN3qC/LSEJT0ofesTk8/oKO63F1p
W6MnxNZETU7h3BKMAYzGTmBmrw1HZHkiyEtPJZLf7wQAfPVlNpuX+4P0dCzN0n8S
C/oq6lYrUuU7pJP9gF3bhl3FO2f8J3PLfeqndc6aeDJ5P5vspxtntRluE/+BpEID
cy3f1cZ2odoLTLAl9v4fbKZGv+EKVX3C1k/X1gTmPP8bkfO0j5NUloIa0pvkb5jd
lh0MNHMcWiz78xn3kPC150Iw/HiGhAMn7uTHlnXvfGNJ2yu52shSRoHqS99F806n
t1NrEbpMw9ocuZoKje/x5AJ2PAAFi3cnm/2Z8VFqwGJnpyjwkrS5MEI8k6AK5ghd
DJ2n/Qw9acvkge+hoZ8orGOVcjWfjBiVwcmnikzdqKabqFyh6DY+xx4QxAOXltHt
pVF7N37j8yLhQLhrPRhsdg/1SeFFjRmKyZ+SUolP4x4upfZfXZeenuJOBe/Xw2LY
B87Aqpj2MZ+N6VkGsImVl2W9MSdtPbAfv7o9MXnZkW+WYUCSyD1fBvXNx0UY5jFn
Bh/P3+Lkl1InebUv3Fsm3kX0ZxcQvnKj1qSBl7/Ax0BJDZ+A1KHcyeXCamv7FbHx
qF1zF4FX27ZG1N6MPtuARUrGXnX34z14cXQQH9gbdAOQyDv3ARjb+cGB8D3rY5zm
hbE+Xvt4mNgWB4mHZKN3zjhgERhh8wYcQeE9b21yMpygayXmZWJX+53iHHoHeJBq
G463pb/dqg95pYWQ9IN1rJoRsUjP0RrB8A3CcuqMzjST+TRsQ2Z6pQxXqeFBqbbO
lxOJAhP8aGxWWVEFfsDzvvfWXB7SDlZ/MGHHFLfEeffOAP3GVTlyILwfwHIa8y4N
kw4IkEVyBUZCoqlaRBd/BxbLHZ6MkwOh1xcDNaVEJ+GIy7k3U2S5XMKKKRnjTIFr
STL+dNzqf7HVo7bphy2qTreOqSCVYco48qSzHXSScyOF+KUDbX+Kc7loSFFlZSzP
hsmeEI1UG7Qjl4kvP1WEEjMMMr2ggRdhDTDwmDZGp2RwenrTRD7QJWI/oEgk22M4
VTy5w8Xzd6hZnpiSxCYrTLYFbi9BroX9YWOaSestxyORdRiTf1MUD9+hmoTGg+8h
euuGv3M70LfcMfisWyLMPffo2L0/Ib4077nC1WIHlJrFmcdQVCaDKq7HkiYfcNtR
Y3GctjDbyEnofVpGPdySIiiY7H/RdWIirsxA34QlBACeykVN7uGY+tkgOlAj8kGB
rl5s8mp/3arzJVIj8zvKrjAagom7VcV/5l3Toi3RKQZKFEOyvZ5h3CxVlK27zp8a
L3289gE/SMmacGGLh6MqXbS3qNZ0MsMgsnVVnW+AINp+TvAQCngbXh2JyQJR0N+O
NtPbr/cwRuXQtr5N+jC1k72TUqvc9XdxcMkigwy8glxo/GaeB9rJoUWmjCkKeYvu
Z/AoFxF5ic8aHF70ozMJs05EL+8+3go+8Z9lHKGbfg8p+XbS5pUl+CUDE6m3HugG
HqzcTMe2OEHUF/vo1Lgagzdnwtk8GgiQNPn3xiKjFAZeSEKH88cLGmFwWvpguFye
hAhbWYSJpYn5rwv3gEnK/JMGgH5JGagoh+TyQBdWayaeWymzHqeUVmhMU8YZjh5m
ygxUnUOlma6am6BQ/ozaJC8CyI+KIiJ9cUQ8nlxad+KD5Sn6sLyP8X27H/Gx1mpc
HkzRXzaGsLsij2ANniEyYsEvlt3WggP3ICIOg4BzyrKJ8Pj3lugAF19QBJbOPlC3
3uM7/rlnydHfqIQvo5tWB9WL5d9Vm1d6J6pTpHJL1gz155MjD9BwDwh7tlTzKBvu
4KH8iDgZmXTPo2yaaKEgJhbQ64QX0TYKSKJVbANoX4OYcN0OaYoZfkUsO/xLWvIs
H0kHg9hwSarqmy0w9CpaeEEc23v6CTeM3jGfFGH+S3V6VK7KcGVAIE2Djp1hSSqA
bAem2VtiKoceCGpR0dq6qXdh7OsYd9O3dJ063J/KlGWIdULgZJ4rZu2C8AZfDn3i
4xgOYCI2iIt5OXPchFEKTsRphV6vr8aj/6/V6umVPalU/nqz3fto/mY9r6HIPprj
5PYvDziaIRPZ0kKvDqvIFc4zcW9pL+gATGpKOLXg0iyeuFyR10KBkbEMYL1GWT62
sYXLYU1Rh5WFAfQRyaOFWJu5WF/CUrw2mddOLc7hk13kT5ixGkCl1b7+vgZcuxcs
bur8lCc9OZNxQ2azmZ4IjIvOIpLN5e4s5JLnVwisT8S9fBH6Da4Gv7zWzBo/lndH
mJKMNJbUQi6VC8v2rXvQupb29lruSKl482T2WGq2OYbewzuToFaWGvkcLzdx6ZiW
ujIkuD6WSaPayKBcPDM6lCLD0q9jvuWm6KhY+ntcxOpT50V7TJCcTSaf0MfuTAef
XIvx+heuCNNrvMBcsb54XZILHN3Pt94AVn2gwn1uqoWHlU1H6mvkQ96qL3SW37uM
jxWMRQI15K2k5CKdeVK7svgAb3/Ks8s4vKpTYUS6dhuLDm/yO2lbQnEeDRoVs7EQ
/EBknWokKfLjzCWW5/yD9XYOMrQNHjgZbKJOv/Anf6GeIsuGv4jlalCpFb/93rrL
zUFOTg6EweDgU7tus6CkBERim22x8QcMPQgWduBn+E2M4yd4gNhlE9iwiBwrj4jk
y81BaRH0qk/uaJbGwxYxPesylx1tWUFaKVvJP4YNyDXcq4E6qcY/lGcWiL2BWS+x
Lv6XfszWhz+Mq7EoQ5gG/fu1yj7pwjCifZvC9J9DLDleE0aKM+wRmzpJTWvwJyO7
ysTw/hyWDB+2j8dYJeJkdOzl5WlbOHRT5ZVWo/HHdMRCIApJY9/+EcgeVtwjWpvN
ZcZiFhIJwTPnU7XTMLrwQyPtdfbnTybrpE1hWL419Ft0OKf1Vgs1EjvB1+LGQEOj
o7D6iEXpGRKv9Jkzis02AIqGs8yLXrlU2Bmq+edYUNFAe05PBupOYKEvE+FKtnrZ
dnCTFo2BaOyLXWHloBCkbxQu1rgICbDklrGXXcRBjIdJf3rdRwGZ1okhvRc7zB7O
gU2RaER6rVu2KezQoXXDKpZcZv4GDlJxRakEqtHYYGC0IhHEIWejUyXjLnvgoboC
7SpgNXyt5b5hin4JKr/fWYSelDMxGNXuXT3tzwVzpC0KaIwZwbHPItaQt4S/cfmG
qYucB3l2g1GKYxaY4RkUHR53NLBp44gjCLUtDeqbl53dkE1U3RFq4IF9+R9WuAqh
ZsCGExuPKjPuVBPA6a9zab/K0ySWEOp3F3JakQ4MRejIixFACkKWUIGDVRSPjouF
6IKPxoXlyDEgXBYLprMwkYlwImWPgg5Wnl6+88zwbb9loTk3B1YbhErg7ekCoQOl
t3zBh9zLdNR4+ZYPAK2HUFEiCtmStPCO354uycVYwIO8BrNPnWuikNjworFOCfw5
BhGrRqS11QLw2QpTdWcYDPTzjkYJNjFrxKe8rTOe0lm03Ct/00ZXpH86rnMX+EhY
JiVfmnIBcah2SpDmwrMRODxW9bqQ8kqgqbbbAnwF2DqEuXfeeqPRjekUa2wmua5x
NRDEgxO9p3cpQW0YRapwNaaVqFDJoI/TiDgpAST9P22/p7VLWFPFOrKds6cSn6KH
8InUqanpoMZ2vjR4WAFEOfVOX0BVmQJqBY70zjnG9+51AEEdpavDKjTRWO2ObSHy
vV3HOFebPpUrCM5w+OmK2HoRWb7b+aF8Um3IcWOEW1QtBILj3xJT6vUB0etDmLm0
bzBU91dT15joDq1KQcLaHt3p/LY5h/I95/GTufdPeX4zN1pbntQbUHBwPa/mQwoJ
2mIL31Ym9tCLJbOfngqOKdcBtO/Zgw8n8faw1PNdjs6YI7tYgv9lZb3OVdzaDumQ
8HTYSE1ty3Y7pleLiIDlMAv1lVPvkcS5i5rh/NtMBFw4eeCjnPjQ+frVA94hUhs7
sQd/EMWNJszyAcaRLmV/nBOH6eCoVaaavDzbsUpG5S4Nr4xd65afT0xoUSvQCnon
Dnc4VT2Nq+19H+/4JzbpNxwnwdXEuFmxkrkcid8vjULHBK+wW6sWiqZG1cGRgeqN
JNE8sxJF3NrCO8l4er+Jxgzm4i9PRJVgmD2Z/TJc3aYNJ5Yd5Y0cp/vf80WJ22/S
SS63DXIvw23pnYr8cMllq9UHob9/SVlftLh+3zLBzyUkzPnjOezY+zuyovktBUqa
gylEuGqWSsH41SldxsIVkHv1xhvlv0bkdseQo/luiASemrxlBgpWDk81ZTKKwgs6
dWDhXwr2IgncVkjMCEEbDp4ccVe0rNV5gDbU0/t3Or+T54X6WHx7ptaI6yip77lv
hkEVCBqAnTxSaI56ZohVCICY5xWU3cCKZJxLNb4FptA0SyKijn3DrwHQn2CXGjO0
n01NWPxOiOobge3IH11BPuG8ZC6wsaWArV8Tzm7RkC7O0dELNlQC2IW1NXwCzQiX
MX2/r/C9dun+yP+XU+i2Y1PVuwg9V2Y7sHXMBB1MTksliIIjpvoOCJkt7TgD/xeR
alK0FB51VyEP/xpFXEfq16XGbJtONlUmgK+DcYDwMV0s7Wo/fUyw3BhZeU5EcBmJ
b7KVucl1dEIhFNgYvSgSH67bOcQoxDBBqfBKd8kV9rmxZC/dQRxHuFSwxJVNl7OK
83fJNGhZ785A51qtyFvE3+xtGR1wL5Yjpsh+e5Y2hqarSXHnl7E1UNOq/DnQKPqR
JpFTShYLFwoF30d1I3M4ln20z/VICeFCklq4QqIBT9mAJp+y9mignDzkrKvjbKV5
NN9QX0ic8V+tzmomnokpWvWPokmb25e6Itjbid75U5hnsIuGUIdxgIiyJym8MMuX
RKsfYvYAE2uslifC5udrmm8j+FDq9qs6JqopVOhN8IYyxpPOtd5m7/Yz3tAXLaom
gK5w+GC/MOc7VqFUqILzU3EXvXNsc3NdXmEc1ycN29lBhODPqM+yU6sPSC4gUwFs
J1CA8DCAa1O/KEyB9AG55fYEQycZPdWCIherty38H6z4aExukoNWo/kP1zhrCoCA
9KbbZhhcm9PvNWZNh/yCZJDb5sbbspOC8QSXIWDQPcNgLnaHxfEEWjFebxFD87pK
Ve8pqBIEM7R9+gVPiuMFhqoqCxNIe/4rqZ2P3ympk5jWQCtp10GdMOySfKUIPc//
bvOnSOSpOMyF82D7RvoSEsSmO0juEOrlyeBETDeZoMRXYf6lAs0JwJaMr8CYvUKO
X6i1tfHxN5Oqhl+kpAX71njK+Xkyzg4WXF9OUR1+G6HddS2wpLbjhsYZylDGbdS9
WMVb+lKQ031mWoMrloiitdQEdl9M0BCeqhXURyZFbsNdgjxze2IgyWrFB037O0rP
adDYC91NV85Rmzc2thdmiyQ6nc7Xo4tGuWqTnhczDtrPXg9+M2ocWVDofwuMefqT
Y3++lq64vPe2Cd+K7p0uRIN8rw2+H8E9fF5uHtny5/ARXazOQv+R94OuGlWcgtYp
D2NmeIXg39SHE0Y9oYRaj8c0OFwpCbbPAee7KRz/XB5fog8LH92sCC7f2fuUKcc3
FWOA1/o3zwFYAXFWmingwa5u4Vzxm3mtwTlhMJNrFzJ/i22C8SXaJ7yxUNYG8C07
yy2N3ZPd0k+pc2E66vaoHqJL7mDD8iNhLtV2yU0Cy6VXgiAIv0MDiZFvw/kHsgtt
bGVsn6ONNJ61hCrWc2whIWD3/tQ4Y3uIT2mi2hq+RXgdXMANxSxmdTT0nwg1ZTys
NlxaDXriTuO+yelZFOzpDPGB0chFkIrYhc13h1TTg/Rhb7ndhQWj1hdsHp6vxeV4
rdf365HRXhYFUt50s8y49pBYf247+yAhVVMDMpmxmtQB9rEbNewALpMvRL1Sueza
zYUmtBZdcy6KZRsrCMmz8Fv4+tO9NwRimuO89fEMT1KBxyKlmSo9evjEZj1uy0mv
7cITqiGNrIZXZ75+NCjixKh5OG6IPCfS5TFJyH+uSUS+MFbx9NcNgFUy3iTyQaTB
P1/L7VroPeL6tqPQ4vr9GfKSHokW4SEBCabCVfXzkDphdqLRsHnp9Cf6H0118vnx
Qu7SBV0VWs3F2wPsGIaSLULxqMjvQK6kxDCVS9DXFSM/oNTeRRqST+JNgtV8hig8
01ZeDNWC+XgtaoyMYCouEcpt/Co4R3XmogG97+LM1mWLZbVnGA0YPqzSK8MoC9Cr
ZpoH3ONT5mnscpa4peBA4/XJlvggGgn4eCECLcIHnUId6uMvb2x98L0kLeeofhX+
ckyIrOl5IZPVgLxue9p6TP+zOyH6t3kPQEt/mLdDVJh7g3yuWpNsQcHEZWw+l6dw
s3iaobRbia0vNCpY19r49dF9Q3pCCEVEhdPTwBIKJzqPOTJNnVKHjSQaSf6a0uXV
vK4H9aX5EAWbHAUSZFfQWGw/GFT3dPTMKGH/qGuLaGsFMm//Wb45p392/pEowgm0
9o6Zv9bgq8mw9Dyaji8iaq5zNj0H1l77+NKSFjUOUlqijH9qAWwFCa1ksIl1f0Uz
ClfZerDc7V2670hp8lxRl/6odrksEK2vLW/pUy1JInpPkUJZ0RUuMRqdpoTdI1E6
lt7bdnxmoppNaPWRJeTaB9B4z/NyoEQe7pjbbi6f4vmbEb9u7WANr6OxE3uHftq8
XqJoiPX8I+oZqh66P5PkMorqZhsYIDKyrrCjwpfAdhelsRcxKoWB0ohDRyo1KZLu
48c/KdF+6YVDZwdoCudOKYGdAsmvR5129/lPaytb/XGsJcBE9ljoPQTieuFO/W+O
uMaqavYPrfM/pZBkda+JJQ52/7f+g/UeZqHh/u98CVN0r8On1Vp4SXkAEraeOKnw
sOoWKI5Ir6Lo7tS9WGNXk3mgTNJ0YcUfkS+ZR+II2uYHhfsHG7dAxY+e1PD8SM5t
VMuT8KSl/eIdlFgiZ7v3Vb/0vtBwEz+oeGHUWHJKQY5SdkBlqKhEhzsujzOXvnsu
Kjt9sJSCa2OZSsmQHpKBvVAbWSUvnaZbKNQVRQ9XYAHwiWKP+2RpNy4za8xTpcK8
05sbfywe5wqntS0v8cIP1fs2Ikl4+9hpoD8Xz+3kDpIdYxBri/KQFj68uZ8yVhHj
NyLZnNMsTwFLZBNKLT9bBLAzWrvGgz6kOt45XWnbJercamW9nkpJBasZSryZWISH
tKtINquY+Ib1wxAOSMZU4YfksX0pRymnPi3efts94xw15xyJcPlMUFJkuUt6YAXK
jEk2InSpZeegPm2kCa7ASmCdU2veG4FGScTQv/IhFTSCAr5WEKWXG9DEN2ko4V33
baXa9qym3YzUrwxEbxZkiFuM1fWVWdfB1y7WL6SOnhSSate4zAD3d3m5aEIJOOZo
rYxasB9u04PSfNz0F4vr4amp9gUq3SZQbbPN5W7NpdDjbzETbsyno+qsKD414S+I
pZ2uGc7mgpXgn/Ft+uYy7hJqQlCAIGZkAQ0PAyWdHYZx7uezW+b8U8mno88+Ult1
8+SYrT/7kBySBCHiKubueNFbckwgZBuo4mlSFwLh2Ag8ku1uJU0yKEKLk8IqMiN6
7jVm+LNRQf26ngF+MYByf52WC+gHazKrBqfv8y9qW3rTfW3VTIXFZXbG4TRcvfGl
XRLnij1b47BVHOW+68omsJrtUrVYJXmMUkIoEQGmkjX+6ZS+VCFUr9Z9dlj2pwtA
6BNvFIgHrJCIT/83GdfdHvzuTgbL1nbbLuiebFWtsgw9ZydmtTcvMJnvqKa29PYD
d3yuqfjkNouMl5pj6zweJO8Qpv/fjOgw10KOh9ICkAjH2Gwvn7CuFoWg5njWvOdU
ocZ3SLmKil5tzSEJ/P93uRJztec6dvOe6OjrnTZjVzMBtcG4xoQPYb7IF8eeaXDe
tn7WENAQ5y/R887cddhgCXD5GmrG8oeJnmRaspUmdWVpFY2tkjfZ1ImH+12eykRg
C5yfv4TijDSsYpqCBjFV4ZXb0zd4BiJrYhjYM3JlggXo6VxBaF7HUUEZ4QLSLAvC
meYCBTRLChjtqxEZYmufqF3pB1eS+GqD3FAuHWeinh1eQ/3KrPQF0kr9PbJBQ/oM
XQOAACx5K00atuKqeaZgqZEjzZhhkIeGRGLKED76PQQlz3MqRJEKGxAD8VMJ2SmW
V6fJKsLbGSAkbY3j+BVdB+BhqHNWkEXLb7yrHGXFo7d/ZLfBcqr4TPSHvCwIRXRx
Dk36SuVtc2mYtbzxgupQEXeeP4Sc1ieqHnJT6N/HodwuU8xYp27qSjiR7eUJ4fxJ
/6m48uH4vm4VbMqL3vh8utAEOxp2I6fily89uldkkKWCH0HM2ri5SWf+o+hm+fsR
+UEUp4fTVK7954m/nms/6RGk4OrJ0fmkfl9NGni29KVq7SKfK1QTiB4rj6J+Tax1
iM/DvPDbo09QpvlTv4F+jAuu20TeP/RKK4z5uEx4kkdsZlSMVoaNkHwYINvFNI9d
6r2bGcyrEX7sATL643dJKr6OkC7qr9i7jhEcbJRSfiBWKY+br61dAVmPvAgizs9d
wZI2PhcEQ3vWsRcbTdXlZDpPkd3yDP1K9Tlv+j9XASXzqCtmACsgwxmIZjXzD+/c
PYzICHqdk1FgFiMU9fCe3WmVmVzt5pVd2+QPn1JB0lUyeMdRh+yYtQPRZSxv6xzz
tH9kpAkXokj2xWLb54Jwys4YAJK3ma7oQ7ijCqeIfqz6G47wXFMKJCP+so2k3cWn
nj24jVcofBVxoK44XU4znAdN0cPMX95gM3tX2MhwIOysPLZdEsMFLVPhmwIKFWTd
i3vdDAMFg5YFC/Qsp9k57fyHYRdnKvObo7NvnJzDDNOYeMb8h0qB2fi8lmXsvQDE
ie1VepAxCj//NY6DH0DtWX6kG7L24BFoCCbK+BVaHuNV9UfkfCz3WEoNfxomcqbt
LSA96vLcovH+0oUAQDAs/RbSWgpD6oZOTn5BwJVegChJQbDL0UurNvjq4ukBnaGF
c2Pw0jIxtmVblnw3oYzMdzvDbfXKoz9hvDjRAYOkqbxuTth0iuiMmgxeAZ3xOy9J
VP5VwRLLwNNZTuy82gXPUYVa6P0JB0Kzq2oGxcraitROxM27uGa925jnSPL/40Ob
Dmwe9BIsjm13fdh6Mx0Hx5LILHdfNLUfgpCCQmvwP/3MH4iau+qcYqhNMX5kli5v
Pvv5ofQKTsLiLSrwdXTWRoD/6OaHncNfOemfFR/uB2exgbO9Cg1UOSezZbotML+S
DtK0lqq6Y5WHkrXPqFQ/f/JWvAGuGofMk92At8ZfKdnBAUg/3L4xURAErKNFeNrW
X+ix6gmqRUSgguKS6Bikn9CCuif3C5w/f9/wgjtyBNAkVlo3TqLELJzS7ae/tTq5
moh9H2Txvft0VtwXbnbIwD2xy9hi5r29luul6hogw+VYtokIUEgD9Y48MDkiq/cl
LOKwFn9gkAO5BkiinzT5XPu7PzwFiEejQjtLNVvvBr/Q8SQajLrAlWfrvgQqSv9t
n4pHvRWPDr5Vfw10sMPGIK2ESBK4TwH7wDtkDhUdwN9PKvxEDv8AL3IJCMRKuV1d
dsdiV4Kdd1QVe+2kAZHnwSpsiFS1XKyil6E2dDfN3XNPtcG9R5vJlvODauN9wbwY
qot6zwQbpQuXvl3EEtidQMvBKRAZFOSCdYmvkcM0Cr5SF1h51jKC4Qu+DRopzdf3
75579w6+VhcJi8BXvsJGl4OKgQuUaJltUImz4YLR5JHiwieV0TfUoy0+n+axtTaD
iCyXWDjHKOTIrqKd/j7vjEun39Op2hBcT/wWyqvanF1Rkd6y9IIOk+niAPwMDztM
VbN7+m5MHdLHATtA1eV5qdkUMFzqObvM2NCTKKbaMLLKIP3HMvi26IKFhISY9qDh
N/DchdJbNcMQDMDgV5bczQUfH8vhpieOZCmI4ZDe92WxKwgqq6iMo0hITrps9aup
dQLhpcMz7ZL4hQuyejlw3Eyy87DP3SO7jOtORgtJ+iY7kikQXsdhtVwKVZXOSAkx
yecZtDndjz3sRX3/Zo/UwvuRphXwWYjaBqUylOT0luXyMUn4ELYzNmmlpQ9YQEwk
IX/posX3cMuOf3L+vRM1otM48KVVbynE5t+aNsJf3M4Gx+qtEAoqOzwSo1Wa8/Mb
ezcdvUT80xqNUNrynsUrSM7W9qaUkHgAdgGmWIn0DgN1ZFkvGRXuz/c0In06EOUA
o0D8GJmo1Tz9HxwcO+mAvbH0Nsw4FvA9RJEoAVTANYPitoNJMg+PSA+E7EQWbmX2
4ueBLtbN4+DJakmiAaxcvvGl6XcJuoikeNfeAl9vViORhJSaTtzVG3IfDzJtqzbT
cQYQCbjpEnyz0WckadI8tKo334lg6rYy/cf8/n8AghejpRXOYpsDqe8UZLZlJMZ0
iC7ENJLktg2q13168ixJTZdeu/EuxUM8cAUbgGPKbOS8Qwz2UJuX+25AdYMuxOkr
ovYs93JO69DXDMEjSOCUH2q9ZLtPyMTRXmNvRJoe5KF3+oYoHayXZ88Jvhp5gYcy
+VeUVr6/kgCUuNuGdxTo5i8v7Miq3SJ2gwTUlaTnguTJbxRb0cA3pxFeb2AQqSUJ
ReDfmntPd0XBdoA/0x7Cdj19Ub4Lz4vkdpFsGq/B6ig4QifVksTh3J4SHfLjd0Nz
jEFJboVwR6Q4LBFyEuyN5YxaV9tdvdnNcuOmUnGtCgz6zv9Eg/qcvNRGKkHUczCO
r9oKh8kpEWfcnILIJirf4WqCEnFIdy7nmm0iEbqE4X9LXzI9KChDfO6pWQqxnSu5
3VfOkkrBjxL8QYxeDwr1q//stx4TvdKIlJsLe4nm37FbxOAvizCTKV7NiHT+Shks
E9SdPAlKxNYJlZ5YkxfLrlMAM7C8pPsQK/ZNciwAhba0F/hs5hR9RY/cJ1Ma8X/R
Ip2JDAVRfZsCohEeBTd80XsGPPyQBa49MFmJgXQUiijpIl+oFPKi3t993HkpQes1
nQEQcf4TJtucqVdHyQxznTX7WTSiDFhAM+cveszBtXxNeyi9+n3YSpsIm8fWUk1Y
3yzYWz3TFm3JkiPV1dIV3DTpJOV7A01g28H1dSvlitzwK8exTE4YJm/VUzsu64x+
SUVazVjJGegG+iQVT6E9Zu5snEbVYqGVbpeyHqncZMoXLnH2nnnlH4RVn4qJNqHK
LAGs9XKdRGL/9awZOMbFJIDOhBCy8lgguHHOBVSGc6DTGTMWF8AK1lWwySMBkkTL
g5ieRhNWERjs6cbwwJ1K6o6SbroksMrCchuGCLqk0WujeB1PeACsqL4bfwFP1kSW
568JhpYN6V/8Sc1gVxwL5Luh6O+oSyIua4snM340SmloN75Ifwh551JlQUVqdgeq
UrrB9oGXtTCvAcL10HQ597fuLmi2iTYPgs4CB0U43iRQua1FXxlwCLOvgEhoZr7K
WnyCuBRQfv6XJnuWuNwBXzGzSbm1dPJ0OW3ZlX2C26dA8mwYrWExQ3uIQZAW0e6v
f4eGYMYnGU9ZswELaCWyJ0TKZ3k8uaWPs+XW1l5ZR9vEc4wjLtXWTS+h8FRVW+ry
shjgEIkPyJ5lMW6vl1zkRvw9nGWjtWhSb3/6CaVMbhhG3/Mm/IDzHuH0fj2rkpkL
fN/fj9S+NrgAKubENAYOYSM509Lj676zySuOvfGWgdD5wD5LajZQ8IGXpVhlqpt1
tiIHHlaeNOUFAtqXVtp8Ohn/6UUPVkGsfJhkb7MTS/RjNqiWb+K9hgyWAJY1jjlF
oJX6mZkEuBhxL05vnrda9x7hEnizpkeVSJVvTWuUdWNdt+yjTxivVi/uSPG8yuLH
ydyd413/LTUMiqPSmQZFZPwANaqAHBdVamuA3flnot3OIO7LghcASs3XAYHKVyZF
/TqjUA+QbkFs4cxfUqEChCFERgkTFm+zr4XHznwYrYjhoDKt+mCTC1cREkes1XPA
LuyddEy/4o7OoFFypFVT1Q95TZ5v9dB4W/kDGSzI4V5SpQCxXVUokpMQQR3RK8+v
PcfCfkYu/4AbKSbCi5bqjq9HpG3BpW8058DG/eJ5+P+UZbxY0MXFnrFJs+AuVHs1
yAza/Y4iJTeXmv+4c3sYYZ3YXYGKbmmgd2LzuSb5yncTLDgG3O7SzAC7BhUuupg2
2JHNouClGoGki52d5uwNxnxFdiKVOTPI4c2JFHKMb4M6q95a/wlLhAcSVbpiKyc/
hawHVrGLGyRC4ee7xdnBcAzce8H0NZndJuabEti2+quNyqLWf/kiQtOrHyGaqBme
LEssV635VtTMpFd0BqBl4KguctHieVan/TkEellXLFnSlarjMatoMFnAf5vz/Nmt
VnezKy5+oAcUlcYpp8CmbuX0+r2MdzWo70Z5OLRs/DN60peoqhLPf0pGoedeu+bC
aYEfUDih5gEf+DYjxgUUrZrSgEJ3Y1VgW+g77R/d1Dcq1ALes0vY0ann7eXd7Fm3
3C+aYHvbgbngPO6jrnM5qvCE4ta0tKkI8QE/XkFQsldAgWOjhaBcYhkFmdddLW9r
1dLcT8i/4/OlzeyKNFO8wAeqa2zWm6ghEWNmLrn/0Yefp2VNIOgHUUF6fYNR4qex
uXl/jGnOF0xYr7QShoKLGZTKSgdbjz1m65BsjD+8vLL1i3Zr8JCe+KKpkqDaRcOX
qrM8eeL37lHEEWQzSqRWvUtPHbgU3rR2dCOKXWWaLgqOOaHWRgz+oQAo9xssr9Jm
dpK+H4qFwxnJEcs+7rQrB2iRA5GFCJcDNQPxTGnPXbR/dwEjz0LQqtyH+YWzopxV
okxrn+wsmMIhjuTZ46fE4g7AlpZrnlHCAslbvqquvGAPJKaYuyoQsSKhXeg6eN7E
TEy9zaXkx44SMV0qKaJbQtgtGzgMRjwEPkr+XHdxx1zlVZlTXCoVlWugq/ctfK+o
rf4mPLOXIrVU2a6BzK9M5+n5DdIpMn/dMS5ytI6u00HJ81BhO42MjYZzH8Ixl0UU
4cxWyUrUbOv5zScKkZ2i7C1pqiV5cHbn1abOyw3Kbk0OlX1K8q/GGoXPQsoHVUGC
cOR2ERdit2UIq+v1z74UP9JiMlsJUUCi0tJiGesY3nUZeC4UamySBAUvcf2DU8Ix
YSqPUpM9wRSb7H78sd/5JK1QAl2jNJ1OQxB9/VDWxJdRBYdyJDHajG8KbZnULzwJ
2OYrwGNCfZujRv6Dp8qo/74SVeSaVAxxNprAbnhdYXflN6rdv0FGlLN3PWt50l6f
08ANhOCyxGWN7JQ2M7LBV1H75szfepr5ZeXRIpaFl7utffQmdRefz+3SVHTQn/xT
KrBX9GuZuKJk4M3kwtyndQHXCNuEIq+PEFlFWTZQKoBa7hlJnkvDWP6sNHrrHZBo
ogUK0IE1iDOTXy7T3AfvOlREzX7Z0CjuK0Sn4xJA5vH2h8KbxlkZKmSuEHtxxSUs
k9oPKm0CUnZTcMA5tXlfrlpJedsgm5RKhOS6tGTzkC8p0qBgF6NtoUQboh6JkVQc
mkZzWB2ALRTs3McHyQyUfkcri+x3i8vKZyjHyIhdeSeVnR2iWNmBSG0LdVMBl0lV
NxU3wkz4Aiq+e4nb/zciPWM4AWcqwj9xKGE7tOK4tXd5rgLSl1ZBjDFc2NxN6hlP
0ZRuMbh3IkpBbKQqfo3dlAY0Nt8vtTmuYiLSl6KifA8bXGP+E3oAOmDAV6bx9AAf
qXjapUemGH0u1bAi9JvZGBpa94ZTYfEg7zZq/SOaJlRsOVUKdQGKLEOpasxHk+Dd
iS7tQufy856aWHjWHre0NhYdVoP/heGsR4WeYMfQui7fZ4uqt7jwv7z2qj9zkquY
KFPdBg/Gk9+ct51nr0L7iLOXfc5GtrzsWAXXp0B058hirgdbMxZrx9vifo7sfo+y
01sIHzs/ZwThWqdHfJSIhEDGTdrzDJwbHvTP7QEfoOTjXwMbAOvPmvk0wu60t4J2
QApjYLXszhbnajpH7wxqqUKo8SYFamj/R0RCszp898Iju1VAMeuWFSIEq7FJx6S/
IjfERVXF1w0kDEyfKIb4XD5Et2EA3OYwjHlrcAESzt1ik6jVp0c76Yc+R2HRG6p8
hhI/RAiAcBA4b+x2hDl3JkEVeY5utIRh85+RQIYJjLTveV/shJhXCx+pmfxGPbNo
t6HEp4oSM8uS7Z1zE5+iFY7MYqctLUIKq/2S2jgPeOnu54nV82W4olHo3yA3sAh1
XlTo+3Px64pfJ+yUIRQrdhUTPnsBUvTW3xvk9woXBzjv7RJ/LMaYd2J8QkZjj7Ec
2qdF0oFb6PZhbk8UtP2McFpopUGd7EDYNrGaZsA/if/uGOV2GSJ3k+a5V+yFn5VB
QOtxGW6iSKX45bELt3AKtiKI85ODfD+PwQytZcR14ZxvqrejpHolBZ5GlGWNbdKk
niZe6+vdV5LRcd4Kw0zaI0GfUPaXHokxYQD/d3LZprp5TTgmOWMy4iT2cdaInLDB
iPE9bVxsmBZL0xmaj4bKx6KfQW/3BFlRl4oq/NOV+jKcYWFp8EB0hjkMuJxXaCD2
anJdRExEnPRPgDThzh76G0KuizM4J1/SjsHmStgnKWhE6EGD2CMbfmPgxI95IFk8
8KabPtWtmFfqVhjmnkp1iLkqahGAM+IhywoIKA7Gj0RERdEwMnp7nF2wCFTEbLRH
cQKVRe2DoPRI0dH/9ZKjzVxaSPdYO4a7aHyP4ep83dVdh89QZzuHd078XywkA3mU
dagCaat39fm0gL2r+YMBgOt8MuEMQk+sPVGs9RuIGnPcfI74jpsFGWuhrxP6o0Tn
TtIFkoF0fySFWUaCstIg/DmmLpRRA2lqRX4I5ithnDtb4yV/tzNY+S3R4X6Ap+QI
grNbdACIJdqqB+bWKJdj7bNNjYMw2h3qHPc9RSeaKvl2Eaqz/hAAF+8BCBFqD8Q/
w/SeyHGsy8FdMQ4geuHOQYvmzXZhYsahIF3cbsUsd4E2I9R2MovwgWExYO2zwu+N
arkj3mtxfs1zevZsL8edykRjs5BeBOBEij9zaeVwYAFhT5uF0z6rmTeZCe7BIKg7
zuUKCbb1GnUO3FvFGD4vSPZ+7T9KPGnnSMYLlrNUeRYTEl7VO7Yvy7tU4dJJZCeC
RRX68uVXoZEZsc5BzNB3qbTbW8E0JWqXWaKjmFdvixapAw++oePnJSnxU/8HrBDg
et1rMWBuC/S8gGU9D4bn/SHThtdoSsZzS+FLqJJMP4sljFRAYRmx7XTSoqy8ZRAU
L0XFoljoBpwY4d9T1BVzjYxsrCPN50J7JOk+gOc6piXHOv388zgXrxTHqQM99w4f
H9gmS31UXJdYcRN3Uk5PFRcy/h70P8c8TAcja5+/FcIq0l2CnbcsBiV5ytEIkjaw
ktPC95k1CXvL6tRPhOdtWjcJibA0bv7DwDfVxJEsfZIPNlR3oh4S6oo9ZsbFB351
3gWXtYfFRP4Xh5e4hbT/NprUfDtJ6+Vq2TUK6usrEwm31pUsvmBVf7d2yZVWFK8/
Vi0UViTZ6i0qyV0kp6ggw0xri8Hb+fQbVBZ/BnEdmPDSN8ByPETUzMN+HPoeIjgL
q0730Y3IE6b4SaY8vzQcNrXlpkt//vyWaOEyfG3qBXK4EsAa/EER2mc0Vky+vwus
NHSt668dOVPXOzvHSNaT6cCgs6+izWCegYUdi0lteEQWK3RGkCqfaJOsywbEtW46
PxPxdQayCDgd/U5ST6r8Q9dZ8pZTHeU1g/U3TfBsG4/VlHA6XNc703q8ZvO7QFeE
crXU4cplOk2vpd23EnUCzo6b8Nq9XIBuG/0P12xsAvR+PZsadMXp4u0uSpCFgucV
FAIUkoa87OIzjHAIudXdxyucfREbqD7cWsR8qug0ePgbw2FM8cu6OynArkQ8y6zM
ksclrIc+5bctC5fEGPJDKDnW3veizJSsanxYhY5uNsgG6mGTvMBlFonlI+XNXzDf
FHEsKudeINJMqkQbHry194vpiXlHASft0rDnyJ/7hPWLa4BHELVZo43h5deA7z9U
0n8afIlKF/gEzReuWotyxJtCwRv48B0cHv8SSLqORLuk6SjASZZWnIiW2Hyxi9x7
A8KhPW8prQ0f8T9aAL7hkH97dVPtdveRDd31tkjcBfJ6b/FFPxzpGsAvkVe2P11Z
1I2NbdCR/+LL83dujQH+6IUQAxmqz0gRmcHayY2TZAhZx1lAB1xh7VPteNyRksBU
22YJ+nlzt6yz1ToY31pxypAXNyJ9TKA82jwidUucuw16CcJJ0YXJPqrRCcmTUtfP
GmV3iM0m1e20mWvaBMAo0SsTJzAzrC5+zLo6Ok584WL/iHlICpXsuNCtIWOZn1i/
1D48NN1XTPvWEvellhfi05wO7FFAojCWgGDzWdAvhaXGvni3EYALMRlnwOlC2tgj
3mLMeEUlHIvd9bE1x2GLJVjPzgfhdfXKxf3a417sFWvLgVGnVjOi05+24+zudIFd
23lN5gvgv0iktfeChAo8xGIcNj4qRZ8oj5xlDuV2P0lRzPJiIp3nX2l1Yt2lysC5
5mlYekUHNgWugHSNwqH3wxFCGtLI5zNBNh01zmJ6auWzc9NhIAn4lmryKz/eXEK7
Kw1S+Xo+OW4dxhNgd73gRrzcccl8FMUkKJUv2XZONnZtWN1sq4GlQQxluSZwAYwl
Px6mc9WxzhVRHFG9qp0fceqyQiqvLgqCg5oAG3I3hNtHMTrgK3EoZmH1A1jbwgrb
JhQxfGuVy1E2kXLSvf9xgGtzxJtHnwQDru+9gzexmWZgDYWXFd/bve2RG5NEI3sd
bsSWM9BAPbNOIW08nOgWMsmdFtoFNf38GXCHLFqrWItKoqI1WvsGKz/wtAb5wf5m
w3lZOUosqvdHxUGl3lGNmbmyOB4A49q7KYUayd1p0BaldGBB6IS/7UsRVgspvHkx
XVR/mBIrm6aZaTClTgtn0QiD/4dyHOQtGNWQRB2H6FPnLiuJxO5fSlmF5LM2NjYE
o630ehRK/Rg+i7tOjNE1JwLc6qAfQni5e9BCsV/x20PEhlgC+96UPWNNEMptLLAh
7CGEoH0Gs7AVtdR+ikIIoSqt8f16MZxtq22nOk8Ig/JPE456tuXklv7wHXG+P5b/
u5um39VBYE2DwO4JC53YA4n9fMRG0Wnc474se3c/gS3Ap2Esn9eIP2PECfTA25IL
PVCmpYAssNWFw4au69zYWYfDQfnzbHGCUjPBw8404NAugH1plIKQEvA8DWzP31+z
Drz6F4Vrx5IE8S4raTeEL6wRNIFdHyj6PVYXGNmY0awdizaP3uETN9dzr9MCi1Vu
pZKW79pJEEQNoCXSxqcXQLHtlmfuxUMIIQjOqRQE0CvTTIL28EZfdGPc2OqpcEyB
CEvf8JWpk55/NnogiW8KBmkKr04HPqvNma0ArSPupo7XYe4gx+SGPKtpXBtOJjgR
mHQsh8wLccCidjhlTSVFi2GDIou80GMY5yCwMSsMfWOEkKKvGhA9jbewlbhWNOXe
mb7fKrhHYbn5ooAGf5w8cDplOC2gG7QzTIAq8atlrKUyxQ3U6koly911fvmRKZ4j
UkvDHUBBL6Vch1ov9bQ3qivt0Z06fHVV+SYzR70Hb33eFHNBOFY9hGIFzbt3wmW6
JCLdMl+tQruFPBb3n9tclaHoy4xF+DFA+4c2441Sr+bvv484Q2z5522lsIVUX5BC
8kZZIVmIVknWC6kV5lFjTXRKxH+ypEe68hgyEBAOWkKbWwjqwIu8Hb+DVt/zoQRb
uJjY1pUnkvpm0vQY3wyqpel2fTgsCpCUVS/qannbyF4lqZYw1tgTL4Peo5plfct4
LvbMOZ3zv8dnR9SnyYU0uOlx7bCDZ2EezuwZIbvQzYZiqSnuG1marRBc+2ZQ12c7
YEo8Vo0A3Fa0fJJNqjdXi7XpJuWtbsK6PA3vKQUHH3vQgeczWUZ3nFepM26b6NxW
wvAlP/jaYD0N7KvVoWSDadxB6MCf/1FUlJfzBupuxXJ+ZdZasP72XDLoWJrc9kfw
fbE/d7iK/BSnjyutcodb+5rFb5/LXxzjp6HcbVJeFHjtsXtwgCGPfnnP2CpFj/QL
0aln89EwRGm9FFa1SW3ZC47kPY36feKfXPQ2C0oMUrYkZ4WgXwZc6An6HlbbelIe
1VIk5323QHXjcg5O1butKoW0TX7eby7BElFwcr6pGvRyI+opIxLmxER72ImvPWCv
BrEJq8JMwGbkMPr9yFlpRQ3vLnYkNDMoGCrst5LDW6XtlYwh4cKvwqw+Iix9k5IE
Yax25IHypPkt6yxVWFaa5B6hrKtYwGj1Zcb0kGr10ZadlH6SVUGrX01WVN4PI8LN
iW3KiA9zXc3vvAJbzsF5tBwvdSH3CyIAro5wyottr9gDSzHpYkbTbr8z5i0S+4Za
MyX+xgSDOc9qr8fiqQvqm16RbAlBq+1Qw2CjaU1wn4+l0N9iIgYKL9ijNNtlp9F1
z0UDE1xdfDUe0gFEaO/jAksMaISv6YHqC4fQ0dl2f/qb+6vt8SpmQyLCnYCAM56j
y03SMB4NfUDpz9SJNxmQl3YXVvLLblDvOhQY94PVxFzMiD5R4a7gmgafUieTDhQ5
uUaJixYCfsA3DMAfGY6j0DqnGInwWvkAdu+mj2kW2IcwScAjYmzEC1JPNX01xGoj
73efYSOpHk9pMamfMkQG0R7gZK7c3/StuYg0EXjiPtk1FBU+MAXH5U/IQN32zCY+
4Qaif+tOV88Zd1K/s/htV1YUYLvEXDPHzbnuMJ6qnHze35BJYJLuF1+SCoeFbBb5
61sJ2elcqUaK3SZl/kOQ0ioJAXvQxF021ubyNW3bl5e1wl6VjdVkKr/sgESwOW+F
8B+m+Mc1OaH0+hPIq6RQzy7ah9hP3A8tpwAVxS33seg7fjmFG/izdjey8YiNmKoA
5Q+82eXEg5Darn0BbKsOJK1v67dfNogbo8pC73Kmlu/ZHmxotSH2h1/aYHBB7Cz5
iS61RmMUJxcoRGyYYi1zy81I7DqMLayL4vVcsN2zcYwVppD/CtvhmzIHglxY8zFr
fJw9zIMVVnAMoTWIDNUz3FAplFmDBzv0MgZOAqdrVpaz+EtToQ/z6MqtFWkwDVAt
6mH4rSh832p8fNKqP0pW8k8uKVN0Sw2PKhRAZDix1eY7K5Sk4Dt4HR+UC3QEwNws
YR0sRcKZEPn91+MqAhoHVsNG9NGoLNHqhzTBzDnn4Vi+rPynlaI9q94Cbpud0gxD
8xZBPxDFD57vzomVEe7c62lSvIgnh6kgLUfA4N88ZtYEOrrNiI/6JD4tyw/ldLTl
XvADQaiLalTNbHltdnPfev9Ixs+jyp7WjzeqYLlzXR/0BqW6kgli8rvGlxjW7wAR
npATb9VPVU7Fzo+pMUs7HtzoFXKSEWCyRCHTUeEhyEUKB3GwRFix8HNMx4eBGGgr
CziMUnU1JMPkAkP4Y+ZaKTF8XJZM7mjGMBuvoUhrpSvaqJYTXsrbsY31zgre+ukG
wAispg+kZsWL1a5+1QzUdd6hLx3Rtqh89W6k3un+85xO8B/Y43eq22Qcd7YsOZPD
HpUleq/HtiAooayNBkyOSAGZbW7T28s8p+jNpqnHfMDB+lx/vi0EZBwj+ptgfdbB
FLpLipIO+qOa3HSpjDM4JH5jUllUm0DE7Bb2eYXF7y/cevTcXj/mX1TR83CXZ06u
Ho2jqM+HOBgbZ/RJfVxr+h8HS1lcQvwOVKKQRDgL2O0nZtsKVpMchdtmnM8i+VPf
ez/3WBIFAVvvppWTJdVzxaSAyfwkUx5A1k599fGLvr2OPr5sEVm1NORXKIiVCxrZ
kaKg48KokBs0bAUHjvRLIrqiP7KJAyaRXdJLwnWnsJh64Yg7KDdow5E+mcw8MxzX
Xalxlgr4+NTEpbJVP7XZbdQfzCxwMWJtAcHCuWRT4fiOvQaD0vsnwuUtlxxhb2sw
T3rXG3FVdq/QgXO7c+b2d5JNiM+pZEf3UJiSCC8L9MuS4mANU3SKHuRsGh+C34Mo
vaGV3WbhxrXAWX6DCVeolg9b5n8oolZYNInDEvGCiio+C4TAvlxmFkHJPy97vkhF
SHdxgzLUovIJ54PtDFQ+Fs73+BEc0LHGeNaj+ZFpLAp/l9A6sovsIkKB7YRdyNqW
5AuL7KoW/A6EtVWbxSwyCbpH4PPC3VCkgH7T++4GAWFX+NjS5ftD8YfHNZPlWkd4
CrOzTLMrAmOa5GCdinYKwM9KySIM3CLixWl2Lq7hz98DBS7GsmXlHgknR0UvGis3
ddfUerLhuKjnIQLSslr01V5zs5iTI/FiB5751GjI8OD2SPhckny3ktIVpr1v70CI
JvKzavpG8aRX1GllPcRZeiEwPOMiR0TeaMxL0QbKBYhB4YrJqfLyesoyYYIw9UmA
BLnOYPDIbK6E50lyeFWSlo0nSAzLskqzWUYOFm54WYMxsShCVuu0jfkc7i+uufTz
cgOcFQ7jqcnoBKT2phUuMIS17omCjkO88WSxlFAse4YIRfQB851QGnqIoMl+BipH
L5xSfCVotPuuEKBUydy9gudKv0PpoyGceslGo7Z4uKITDE/O+TVqbZe4FfeS5j+0
7Hfomsb5meF1AfKseJKGNaS7cETbF7qI6z52lr6vWS9wm3/R8PLtwQTvLMAr57N/
C87Wh/8ZUIi5itZaqhAnbKJ0iGuYirf7OPrpHQXqPFCZ4QC1KPChMFdYKGeddVxa
P+Ic7j0aAtyg50ISYiQC3eWdDcFNVfehiLw3RxCUNTdWhwwiDnNsVZoL4V/xqmHf
qU10YRm8gA0to27KGbhoDsKFxOGZH2l4M/z8EB2zK2xz7a8jLArLHnlA/70dtvX3
tnn/UDqCp56w4jKpBuXZLG2m808nzJ4biIBBpJNKK5hNvKEGwJs4lrohjUMSs6A+
JEb9m8/gEH6clHNBdoWr/UPDitxy7UFHB1ZHtewikxoZXTLK3zo3d0B+rR7p7rsr
nJQM//1vkYZimDtofS1zh7CtInjGCgyhTOHP31eTvICLvAISSYdSKL40ZolLWMjM
UKuDZfjs5pCvLD2wfv7aG5mARfJk6nCe18MxC/5Tafx+tTgnJAKmoB8ymv6eWOZI
i1JgD0fXeh7X73RJM/MWka43T6v61y6Hy4pu7phow+URtODmoZbyAincFb9Y6Ueu
XZNtNTUU0NjBPX6o2556yxFC3bkrSFULGxBR6Dl+UrG8d2/TOd6acRinnkjOSvip
o4SdZ804BucXjjGgK3+Jmj8ld+xTkMj3oTmqLLIQ4BcZKk+Qrkg868L4LFrnWVmM
Rqj4gfjXiafpwnYr77z0pI+SiZnoJzVrmW78998984a9E3tZCPHTX7ohZFDXIZrR
XNEnUyqQxahVyKIgHKFh5phyusbB9hIZ/BksS5ts762bfzt4EcqdbqZgJl7dmqL2
Fu0b3ZiyV/FKBWNiGbEWEOUIWeGZYgKxYCWZtb86n7MRggmudV43FrS9YKsxOPaQ
FeP7cu5agOAYc2dUpi6C2oVQgC8piHJa8VRfRyqogf+sL9ddFcdw7VHitaQstWsY
+rRxA7VIr/O5TuNJdYbUTwe3kPDl+lfxlRMbc18aO9e0EKjMbkfATReQGRq15ehz
p8jY37uJwSy+RmNBBTYs5Hem/nZ/gasBHhGn250HL/CyWhe9zmOOPX6R3jjLNtFV
BTwqK8ECOghznwg7W+eAUI/GjZsHD7GpLuctrrNK4tC7FFzivzWgoyW8jB/cM2Kk
8jCqtjYnATspqdiX+7QZs8VLIhiDRKw/oit0uDx9fybEgvNZXyzkaZxAfVvynH6N
q1NxXMxqI4mYqc0uZlKZsrpwubsckdnkP3tnIaYOGS7JZkO90SToPGD5knSAJ/Rl
xqB4SY3kRUnlKLnnJI5+xp5XsNS+Q5Z/2ZHCD423LjnI2Xs8JmaQromeLX6DBtOX
EVV0qzWckvWUMZWm/iQ6du7cVc2iLHseYAbNlhq8rlryVy0zqIS5anmO1Rj1E8iR
3UxQKeLAM9kLc8YPFk5Z/5lDqz2gJsVSae3NvPtyrUIGwfosE08AaysQSl9p7xxm
NeONVR+/Q7oYJIhVVXZ66+iT8vHGbLuuMnAX7S46c3D+Iv3EB8iXkzFK/kOIJ+l4
8//h1lSSniSlD6Z4Q5O0SY4oyp6FE/Lu2r7xtKDAvq1P+d7LCzyeLQHphQDKYPpz
171CUnozKTpjfN+Jm7e1hBXF/oZBX+LOWvtty0AJHhHSpsMEp8krEwBUubFBuiGI
qtxrvjuSLiLd5NNkmm0optGLnCz+hHh10wxJH0TcT+wvuQlAjDgewnEtBc7jTaPU
xPakx2vzMn6jxbrqNHU8JrtT1mr8KFgsJSgpuSQAOYvNlrcxoDerErpomWwAQBc2
Gr+rhA+rjy2HZk5urpYdr1+SngA12aqdwPy2XSHs5y1sN8NBQ58Wt0BifVdsGhIm
smVv02bSKUeztgm+qaETgOotdsSWs4gnSCaq7msgwD5nANhOWmLUzChX4aWWuoPb
zHuAg8WKAXN3O5BZ3SUGtb7JUdh10BqgIzgHv8jQgFEJHgQXfGLSeN3vdTVyuqcJ
XznWNbWt4rzKaOKeqp57ij/aO1Pu5Hy0O5J9P6M5Kr1oUBRKBIACkjI/GGhRiGN+
9LE5AgYfNOm2H4DCOjT2UpSobMptZ8Unm3U1+2x7kP7jOF/hFbkcsq15bNVt0QFc
AS28ZgzOLdJ9NEjpoyg0JYsnqG6iDBdfn7YhBX+nwZ4Wvs8R2jZqyRxPw+ycsYgK
FIkcs2ZfYlT6zhlaWgHjitBQfYCfWTyTBsmeU4khddvqu7QCExoP5edHFjhtIgnK
0sESL043Yp2Kp1OcHzemFZbMRm4jyW5LBFJNSydIGwhXuJOuwSoazBgTW2IQeaq/
nIDbWPRsDkJLS81CrcLIkN3N/KW3AunGe19IJJjrR18hulaTSsGWUQHHMbcYKtQe
6L7SRjkOr0+K88Hw7yeGcwbjCjQAXi2Klbt7SG5ee1VCGN9EP/jGjLKEc1HLLcgg
JDg8kDrI7HakYTXWEgKVTG0o+uv1AB3I0JrrnLJ87I7l2Hh5prxRttK6oE0l1Mce
3vpiyKBMRPVXD2ZSk5Ts667Pa328dX2wG7+sMd5wUJy7ldzjTLID+n54km11SWtT
EzASGhRSliD38vDu9+gmTmSTN7uYhDutoW8yIOXUZX8h9tZ7/6FCo73yvF2FITuh
9X95xuS0x686maGIXWyLtQ0qvVKiZp6bP/TtXGn0nOZemdSwoFs0oDMzYjgcszbB
DtTtnyno31ZA2RF03oE5VHWkedgZ3hYxbxFqOxp9QpTLWjuHAKLG9GtZKVEb/DYH
h2ERPDUPUhkM9lqoFhf/uwRQRkrrRXeSsgElptO0GUmsHFiu+QypconDvitmR1rV
pyyhHeltfETXNnfhn+Wbylw81xAz9QYJU7+pyR8/wdmii4Grib4cvQEfAWOC9g4l
5qh2LpcH6Auvf9kxRswti1Ph0c6+pUqJ0++GlUciY29Gl/b/J4ykXQAZhwFrERbu
TWwAbiOyUcHAsJGIQltP4FnN+Pu92vjpUi/s+IlmzCjy9e6wnoxDuyjP5YTYyoOt
bE8p6quk2Eme51pDrLpPVSoJLo2REqlRAVmdqzjn8oWeMUpq/BwHTaDfDgXA0Bbz
1DLuFbT0jmS4b6SmUYjkoN5egEWXf5CILTqAeQappr/bNGtGiv6wInslGInbnjUW
HvZM1pgVzlMep5+qLEEyJIuhRPtSizvT1gW5+ePjErzsg7dfVCry9H5A+jcoozfP
No2L7Uvc2Gew0XkWlaGqDyV4umgvt/bXLJ3SmlnA+XfNYLqD1Gmmi9mvapaMHr2Z
ocwe6ZR32Oyi/VHcsQikrFMy6p4IuSAOQC6bvlvaFn13TKVb8SSK9LL51NU5SZuO
1PGucdqvC/Q7wY18IElW9qRbNj9STh+X1rDq/yR4+4Nu+30r7+riy21Ms6BaBVAc
gtvHakWXkxk215UKVwjpg8tTaOhXUwYxk2yp3voWJGozd50rKCbLZB+LDCY5Nz2d
mC2+66LSOtBAG2MIr1YgAylZiDSj68eXCyjwK2iHijJHChyDk8pLrIvjf7oCf95S
sALNgKxPKGt5j5fEDIEvIggkRrJ9wdjXGJkF/HVX5Lm6WVxIY3MUZb+Gbyk8pozk
KyiPw9A0EnIcZwu/3Kg+KQpbKxok/L8A9jl8ivj+hW0tlAq4wyTP/OR0s7rn/5S/
oOgG5wHccCnL5iE07XAUQhOO6gHjb8B3b30CZev7NMEPj2C0QoKzUo+6/DeNAVqV
dDNCD2Vxsf9harH3qM6UlTMz1DQr0lYHRqqqa8puu9FTLJ5IrN6hk+1kwPZ48P3d
0IPDbJ9O7zMwwP7POfzthMf+pWRNUe35FCU/Dk1LQ/npNUBPuk2957mDxcdx7TDn
tH6NoH9OAnVsecAMAS/lIgOcgz+ghrqWnfnpNSXIe66FO7EJKSRzNLukHGsMpZnY
oX/8FtL3PGXib+oYg2AoE7MJERmy2yQ9HxaPfudTzJniQvkVLlEAIdQ+OU2b3JAU
8eD2cITqXFON6ihov4F22u6I9OW4W6p808SOWpj+2rozp3KiVrVn2XazpKisodTp
q9mx+Yyhx+q085lrw7lRbEHG/6n6yl8YNF/7Q/M8ObdmsrrsKVM+uwXtkgIk/qHW
r0H3TFK7ZYxzES0LxBbJKZ1knb4xSmyPiZrNXJ3CHjmIxmVwN8btTJX/CSkgNS+I
PSiYg9/bX7xShUD7u/T65bdMi7fbQtmJvVJMX5xh1aCGC8T3fKlqDm/JSCLOIPFv
q4dQY16NtnBxMSA2mN56PiFWlun5HsANvQ3LZtgpQF90yUQJtJkGvSjAmMokCPIi
LjxX0e5gbEX3jDp0DDCps6l6AW/AKnwOStivXnh05NJeK24DlQfVqcSjUBgBinSV
y9Ris19QaG+5O535EP6LKk2oDYsio4QwE/SkeBOeE7yDtWyMqQgzor+SWKQW+FVW
4rU3myYjZePFU1bG7RY8x8HnHV/9SYF31uPP25RLM3Jyb6UqwBoMya8a4EEZl3IE
KeeIJrO7jZWf7Aoyyqwid2jYcwYRTPbTABYiT7zhL4ew4ne5oHFrM8L2mJVMi7qE
6DPj2bTgvM5QUzv8ecAW9h9C/O5sJrUPvahig/vsDIkxtfq1sewvcbAaWcUpkONG
SEtoE1HPZ7ET3YOVXQ/5gZrVbla3N9dHOzAtFCzZAT7vJP0icyDs2KUjzE6aeNIY
R+rc7vyjfeh8S3Lt2n/i62QqhgALPgfxxFGzgrScR3Aoxnn/NEPuJLm5NMNBejNU
ja/v8FUarcCBzT8zvGN24+HyeVTsgJd46sqbXg2/IkTpQ+GgOwCCzD02un8qnf+j
sPlFxkt/tLXujJxxSWbUeIwjOwdPULVJ1O5n4YK9S0jrvgzjBNJLnkzMRYK83hxe
qO56gXRPw5yR2ciDSCxJdt0PooESmLF4gXwtxWsQQnf0UbyGks1PdQG1xMO0j5kc
Mfz3AWkgplvVXUg4wED1d34RuaVHrN09MCnPq1akVBzW5pAWevqzmp62LB497Uqd
nCSncj5oazCPIlhyadXfZmVl+/Yd4BchD/Bu9xLcY1A1okjjLFLnm/Wi8eOVYaY6
i0JO2X+6swH3wC8UncNGEUH03rDenj+4hpLMpaPk8L1DYJFzvDRnp6h4MS53Nlr0
avX915HBuT9tJinfVd+v1kgcimAtdAEqbBOajl68MbgvwffUOZ5mSr7P2o6oGoRC
/DqSum4xOXAoXxj/lzMdhYCrJKhnm6Yy5lqBMBaptZmc6A2vbo06isO5CcEf8BDh
rB9Uzx9YQW2psRmZOiSr3N5vmrX8EAbSfxhzMeTIBWUITWOz5saEmQomBKTftmzU
Mmtr+JlbD9NSQDPRT9V5XCBYiK59kJ/8kwYe6pYDDn+wYZLQv8RzuGkENCcJUMoG
ONXY+zg3fg4F3FsD5pmVYqcG2QmwtaUgKV2BWItOMxytP7N1Qfvkg2/X2s4r56r7
3f9G2Or8kqbeOVn8ZjuW5KbdH+nlvwKKK8RKwbBjDmS9nZFCxTbe35T3Z/C4+7fK
pn/mlSz9ec3au2U2R9BWk2TE8XLP3QgZUbNkemn/oc6VyQwFmx/zO2AIaxPRrlJS
SgiNkCbu1YkybW+VfxQezAcNTC1o/Oq458pA5Hn20DuUeFzzDrsLLJCKAdHhnzhf
7iNSjuHgjPUfNd/DotbfD5SUdPt6zcEkFj5NVygAbnCJ+Y/HV/yiYWu8VZR95T0O
eee7sJrZ2dCsdPzfhRCfiR/1CBCjyEyFIxPW1OGCq7IuwTC4bYelQlV4xnmvIUFz
sbf7zWXeHZ1qfZf74oFUnfMfrcLKGLpBh1GIbcEzlntNEhbKcBpczyBBHzS1sSlY
WLm715rFoxSBceb/fxOEqxoWUwY2f8k3yz/8oXN+jYpEMbLoynKnYUU9AVISBGoU
qCa/TdZu8WkbcupVRUNgnXz49HNyQhfSrhF9CwGsoUJhI9Z6qQtunom+0J482/ZO
VVNMD9PrQbgJqrNhLKk8nlRBAi+XgDUgRXzJnan84ikO4KqphcEi+NNjBYhOgLls
/mZ217jXItZOOdWho6ygjDoOzg7p6sG8sqYMqTmS7R89vmnBomyX3jK1M4mu8hoY
JC7EaThQZHCEaWOGKlXbp326NBeAQ2HTKr7oMAvjyL//dYen8JBOx+DDN1GbEoVb
cI1VDqYF5kBzbJlU6blKrPoEnZA4uRVcFX7TKuCftuAj5Hy0uyYQ4IxeguTYc8st
5Zof4/0s3t36V2z5q3ZJysdLIMPxZjg6YCfvWu3DI4C6wopowAXWLovV4dRcAH/f
Y6Wxhs7hnExTpQoEjf7bdXCa7V/0bkuNG8GdKZfaT9jO+s3EVRxpty9qRMyC+qjv
P7UZs4UGPoJ7QuHEzSju8q23pUVGf8n9O4Elqy8jdjQcVyOtYtOwpUl4g6XPSUUP
LWTWKYZgx7Azw4PK1g+l3hqLJNuJSr8DAl5yvnBbXLig/607QBLqYYiVdNIFM/lJ
jmT4myVD77JL6cKPfK85TwDS09eH7KDleWufRjL6HDk2OWstST+G4VBrAuWMg/kC
QJXdNlh5FWgh4paVV6wxob21D7R6gdAzKJxa0Fhm95MP8JLmvvxq1LzUQBZf3gVk
1zFK30YiFH5butQT39h90kKmgf+eHMCEAAjBPWiPEWZ5EzisN2fmPQJhaqx4mMJ1
bSSzNZHtyZdXqqvOHKWuGwWxIs//f1OqVrojMrCXg7NT0nwnuA2S10Ku3Y5EUHGp
dXOQSIWTmCEQeQefEtb+cxZWJ+lavur3Ts1qGFUl0MBBW8edL/VSWghAbMA/jL2+
mBmorHFMKPOsosSCCfpTuMEwvZyHda9zaGJFb9oEamItpbM95SRwqyqW9lFlf5xF
OFteFf6LlDxkWIA4HXwjGeE6WUzaFVmlSs9OgKJUVqgq2N/vTJ/mFIq6DulpNsgh
NYOUwQlaCyZZi612tomaaJWFBJ0iHP54qIsm9/kCnVJIEUd0hasyN/4C6acNtQQu
8XS3o/hbu3gqzk5FZAXCTFukTrptyGOpKADtwiTf6Bp5ShmkIXf06zVH37JR4l7n
mLl/4vbYnAzOzETNBQRS64mIrUAY89MdQBZbcUdc0bI/gs6zjNMwwWDOFicI82v3
hAlJE4NRhEpVJcjF7lAxfx4MgwK5Ad94kCs2zikjjS1Sh8DEGNZRMrba79qjsojB
hbRnHVD4csdJjsgcRsst4Cmhfcqxal/ulWDjimZkyX9fKOf6MAQNfcxV0RM9pYNI
PLChg/X/Z+TwrlLCFe47pi7iv9yx2G92U2ZJOuBJ9xLloCESU6swgthL3CPpqiWz
9nJ+lZwoJOZN230JJJ/zL9Dgp0vP3n6nGhO3Qr9wF+u9C/zVoQQ+B/BnNZmwl2Z4
l1vJ48hwLzZN08EzH5p45fJbXuQhuTu0xTQhe6y5H3VxoDUcYFlzOWzduyNen54U
Kwp+nFk/51Kv1PvmVGDKt610Yu2qra0/LEMMgCt5TLKMREOzQ2uiQ/tF+jxSG4xi
t+QqTGwKuI3gqKconVyvxl9Nke9u43+WPGiH2oKWAJxw4zHDwQ47GVnc0Smxo2KR
AduGBQ4iuHIT4nefw7WZgYUH/4imouYKc2gq+J1wGjzqPcms7GFsC1hb8PNKXYTJ
j7CWeIlKk5G2BjWHSR9OZkZOpQc8zwp6M5FVbyMSDrqHibcP2IXAAHhOE4o8Phh1
4FPoeBoDCculXQ6q5Dna9l9Ok1fSO+3PKSVfjnLsLCbGGrIAtBnRMG3VfaPZuL0l
azuZmNzMnWBJ7ngNsE9NP7V7bmc+lg0woUUvmdV2Za/BZuOAgoB76Mjq8MqZbKI8
MojoFcPbr3sqWyG2KgjZZUgCJHc1YpM2yMdXb4+2J7b7iJKPj093P37Q0ukcYvku
2n6iyk1/FfNtn+2qdbDg/BktbHA+/HY6MOm6l+lmcDru34dqI1MGdwYssy0r5oTX
92cBCya3XkzJa/y8Lk6TXQg1/GdPIX4gWRR8k/TbgRG/94m2qDlGOnWh1KpAJPJl
5CunNS2zgZXZj6MxDC1TjkDulear/LimwJ2S53ls3balFhghuI8onRZKoK3MMcnD
PQYAnZmjRgeYPObrK+ZUo0P6/nXBM/vMQ1lYhuarIVe6QEpTjGai/7ciZMkavJGU
+Vw8e8w4icf/L2BqM1Vx3f0jjw2X13MBNVeN7+mki7kaQdyHci0e4pcmF47uPdS/
pBY3nwAv7NlgacqfpDd3rmzGN/GzOR+YYW8M9CIxFxeiAhrXPIspz0hzHfkuTQkM
S1P8LZ13yuNPndPIQ8jwaKrPJrWRpLzMksT1HFKHjgJOS3NYlUDcElBiMBZsCamk
mX/GUMtp0yqEiKBT8j9sBdsGq/2DQSACUNWQLeS5ARw61R4G3uIRdCn1Wk3LVQa1
o6hTjNwFJMNcu1Tj0yTHrMS7yhZu/RjNywsefscypnHhgrt12F0N+ZowdgYOp31+
GKcUbhe7FY7gZFxK8Wc0dCDeGLdklmO4UYDbT14sMed33SQxqIwORYPR4E5RcWky
XkhYbmSqkQOPTa2z+FFBycH2J/aDoD52Wb5u4oWHvd3PcThBFb6gFNtOGmnPzxvo
Zqa4PCCm1qPrwFcDZsuvOP9h5Ed2z9qHD8BmNQGYy6A4lN0PPhbvLoYkFCCmvEDK
dBaZGZUlSzrRDGFQOh5q7jZAF/w900tg3GWfWTeLmp7XDWMvN42vkq9IdU1ImYzW
njwqtIh3uIbLBwDoH1j4tVNqcXCkAWTIfC6zZa18c7UrlUt9i5+AXNIzrTgdcYCb
QkLbiV91m3Swm0sp+Q/duvr+o1RXnvvzGnmLbakogi21ebvDJy7xDSpvHW7Rit/W
UzDW7ppu5M83Ll3iq06EFHI1+mYdXJSaLQ+0zeK3L5aHRdm7M8OUdJSaT/QLjYnB
Wx3IPfORGeOLed1UlQNrOjQS4BBemvRKUUfry0d+1OlocaiBAtNsNP96dSHDMSjG
ZEsA+Q124ZnNeB5wkymUu+2RCkH0bRav7y17MBxYYpGpQ3cJwqmvNI9hwWIwl0qB
3KsGi1O6r8F49frJ479ggZrwRY49Dh4KtgQxUidLIllPdUL5kt+6dn0Zaah13Uif
tXhkl54VCSK1GmVj0MQBRULzzd27OwgTFZKcDXFX8vGNZqIOAa8vMRxwh5To+7aA
xi8aLzG487oxKY+sglI3nq94nhJTwC/hSZb94lMP5BVtamObMrNRoAqwi45CFLeE
K+WmscAFxgiwwBzBW4abHkGM1LZrrOJ1yKhujQYCrspcdHfLGydaDLWkxz49hQzr
R1VJ0AhrHeA6ZEp4QvPVpeVH5RY29kr2CcyYECMC9ccY0l6adKgolToakeBPDRZS
wYhYVR5atlxbboUSMdbfus/HCeXGSf1XWpxmOGf/Qz+uqopt9ZDh+JRL0GOxmphl
r2biIdg3ce6GKqRXlNxsmsXyu6CmXi9DrnhEG/qo5i0GgDvhroPa8taJ+d4PR3Gg
ognYSW5Op81NrfvCj2gpDPVVFn46zRzg0J94WpF7GlS/K+RRhhxkgS/RbchAB3mu
THklOCb2dlvdEsHGCwPwbCraqtPVmDZi02S2I3Wl88i1ODkM6Ji9DyXBfECk3/dp
25+KeEi7mp8yLcjEeUdBkZkfy8bjlhHH4A+6ntNbZbOKXwMJaMrnRytfH9iETebM
WCHqINWZkaHJPUjnc9cAjr17Lp0EeaTAkNBwr5VWUsPODbqYuTAFE4wffQQfz86U
BQRsVmqploIKJTQDQ2lmw1A8BbyolX29ljXGAtBJ+TIf1tUB6eYkyP16eWW6BvPZ
nmi7mSUqV6do9nUx1CoUiaCLn/gU8Vim63xa599K3HORQKviM0njZXxsd9SOx6Pb
Sirl/RfC/z7QQk/3HLPx64DdjGFjvpZRMWMWWXbHTnjW5uA1YaPeXbVAfI19AWhX
//6wN5bxdBVzyT7lslU/bU3Y6T/91JFWZ356MYy4d/NC13H5eqNrlszrYWmgAPMA
zA7Oq8B+tmnnpr2lCxrqrAfkQ73ynQnNm3ePfOJ2OlmafvD/gPfWnfWvYzlCnz7H
+gEnDIDBdVmeKvoTs9B3uixFFjLmi+Q3QtAoY5n6wzJXaJmchuQ4UBds6oksm3K1
0lNWgz/lMriDH6zGAQPqFhNPrDeOSlyD53BJiMrCNTAPKfh1UaraIMVLoDSS9DhM
A95061WLg3NmhmllMltoFOiNC4jWNek93h3b56ESzdDLdeVfH7qYbVwfaFPh4oIP
WXyp6D0ZGwRnHs/ptdKCeeiWa0YdJK8gbh6fLXT3ua8m4yu1el9r2WQcy5THgGgc
3ydNRo7CGJ7cC1iHc4Til6iFG9aBpwMG8yVDXIOtMN7xuM9hjK48I99/H2Gd6TDC
lssDny5jNB5YP58tnv6t3DJqwe/cEfjaxOjdoGACh/r1ZKgucVunL8T7mcbLkL6Q
L039grciabRcTx3DBSKt6tc+7VDg3bxXTPh5IM52p87L6uJQb/pB5Km4pyG5p3JH
SdltyFJzAS4FBHBTKLswl+Q6PzOpqXXqHP2YxpgWpqWXuLVxyVo83w5VKoLu1mmi
bbYWdump90yomBp3pM9xbaL9X4uwQWu59H8+0XM6+NGf2tIjvMhA06UGmbJa87ts
rI6oLhqa0CUGIo1B0ef+cOW2haKPVNMr6eNOmh+r+uOi5kMOvHd42vBkkTbxIfh+
ySwmHYqUCh/FMv9BJSYGv0KFE6fZFMBJ8hQG7P2QL2sZJ2F/q1bvTmOvvOHFLHT4
iF9xkviIHwzJPzIfUz7eJvxS+ia0qwaOBPFv0vkK8EGuF+Lb9PrY88HQqNG0R3Dm
y+Su0fFffbKBfEdAgFrYhV6QBFJb3/Pgd5JMk72EZm7pjz8nUyUFL946Nt4FRgoC
VF0cuRSiwQsuPAmHRqkWza1EfMScEb4/Si1Giv8DmpBw/3BMR9nhe1M5ZnW8MI9X
wPBcJp2yiZqKB4y2bA6NrAoc2fdm1uVn6/qHn/UWYUKBBpmNmFcygKO6IFRlNnp5
bKxE3moMCO3gm5GxPc0Uh1TX9WD2Lqqq6fbRiY0gHNtoAN5Bot0RLcUXXqJ0G+kR
go6O5y5jM85cYsEvLBIi8jLGKyOgxp4EBkApspPJF6GVNqxecHIVeYDG6mTsWEt+
r5Znks1wL36PR+Vlb/0TvreFPBQNQW/yOSl0eAvs8eRr/RmMFvaizXnPzrvsBHbV
5Yb2Gqw/GWsYIhccBc7D5lvGRCUlYnuBjydsjxwtOpF5BNmM3xd6XV4WSSR2h5ss
26Ovw9zJ//vji4xfWBonVTiIDKxWL56h/iUMxlV95gU2/fRq7woyGse5ZpUNqVCw
7jTPI61YYM6UOYwQwL4GzzN6N2K2uGChArsCc9LHUib3poTY5I4Z1dQ+Pxy06diW
H3M6cpbG6xMf8eLohKtRrlDgZVLhUP0/IZV9otX0j7b+mjNa9mV+s9UzkH93qijo
xho4WcUJIALbazmpbFZVUHX/2VDtgPl7BuuCHX9mEOSFotS+QlcMNd9Qhij2bD/J
LHndIxu+zQv4n7UyWCwGtEBT82w9NajdL2Fr6APCfURHCOvdiWP8vw9GZs0ZTttb
mU8agFG9+jRkihdk81dLLflTpYTZzqAW0HKSlYj1cip7aBSaDRdRkZjyd6BIJumx
KuWa7/Zg0pAWgjALdHfY3hBFIcU/OJFDK1PfhkP0odJW/O33pDtL3KAYZD8WLhHb
YNd2pfsWc9e1l7tRENd/MOMqdBQqMCbw4tJGTXOhF8e54dSfIvtHbVWcvM8zqRsH
s+JeZ6Jt7dOmxHyz/DhcRzRo0hHMT5k9T7dKJJxi7HmeIrx6qQIczwzTVcmmQBqF
6zTxh5avYbjq7kuc7ApTzG2LMgStVn3mGoHXpPKiM6vOqhZL9bKivW98wk11TMqm
HQAdpz81pxBOHzXIz7Cb+eRAJFolZZq6EcF/NOvSzAiSiu/y13in0riPjAtXdIQ4
FaGqZNpZczHn0knV1pjhyz4W2OIL/SdTGfJhQ8fKsla9Yw9EtG7CK5CqkOaC2Y5A
uWYsjIiLS6DguDZ3fuyv2vAt7wlpbpLsq6lz7anCyk+h5WE2AjivGVWDUjX1zVQh
pZuUo+LQqxK2yur8OoCTVq347+j2sFqWkBUFlyOevue/lztUsSGom47Y0yUwCPhG
rtzcsj5MvXC7FHTIIpHAde5AVtxdO2UfiZHmj+/B3/P2bYTnquWoBn1GpCitkX0e
pAS1UxdS7UFgfj2KJAKnvZ0VLURgTwMMpNKSwoGqtZ41wNzRXX6ZqKgUeBJRzwpb
1jxgxUcRCzYdJ/RS2W/bUfAAvr/pJerYbFatLyvC19Z9dLLQ4vTRBediurbbGMue
pGhE9ZSBAEQ1QwNfRV0WzYa8oaWh/fGZnQdBmDhawXKnA1KtGvdExD35eBLwOHA+
0rWT6fmSEqRj5qSlyUQSryQ7evBwnBxBN2nTBQTUkKQrdKY/V1Htq4GsJHaXqolN
+tD5g1hmSxpwMFI1FDii7fN3ZwKjM3EwPO6uOfnwM8CuuOMkeZFgKHVyVQrX1y+U
KArSh7zTxe37b1z+pqZABbtl+nqiXuSgtOtz47G7mWTCaWCEA0Glx6nEyM/H8rYH
iyzo/sLumlG/edkJgLpzAifIVfl/mvJ+rPGZEjb8KYCk9gz0Yzd2b3deChRpQbiz
mIiylqCVB3t6hMnMKldvodEGrZSdBW3J5k07iJbBEFnjzSeOtP32adWV0w6dkmm5
si3y2kPQFdsD0yRtnu88BbnNcIYsxrZFVkCnrc+9WSK/S+cbOhXEF1Qwb5Dy9pcb
vkrIV6EXCnTusi97CRXW3E+4jsJhOrYQiy7N9eaKiXN/oG47HhFbCth8EeO2/iKF
AbObiFHzH+Ko1CQcgZ2OB3cWS+kwb3gP/SXn71T2kJnG21WHAVOj3TrVJBZ6Weg8
4MWawibMT5+yRsq0IHBD04PM4+YwA/QtYZegLQTwHrjRKiaObD+bfz3wN/IVtwtO
fjxAR63zwmbWPAboTZrUhBnsvl6FAY/HECQM8h2oAQjjh31kvTahdzouEi8nMuVC
BViLLnmniwVlrxBpCNJHWt6QnJn7sWGBzCl2lUApI2eKqUz7yiSPjsmwDJvwCoCu
kHoXLmlEWFhPA5+rl75xU2fkPlSuYeM2QdZl64u8NAHctS/yi3+NJSGH2Zp4M8gt
VGWCmOEq3Lp03n0RjuAYE07DxzGmSw6J/eo+GiTzV+yFLsVph/G6Rq/vVKRD5QTK
F+fXmB0NqQGSIcA4hnIXinQWI+GybHStpf7yd2Pibv14HFB6Bgx7RuoFh1TzSq9E
v26grNdFelptflfs6NzrY2UvNih00wIW2JzHTHBJFYRXVpNjYixHNjQ1t4lRzfpl
nFIDHGWbX7XdGmk8B5b2nRlSK8g2GBh6spCovc/D3eDwaeK0vl1caAp0Dw+9BMuJ
pxYtslrSKBzlM/XeTjQ9foMRIzWkNmdvoNoKMKA4uHgQE84i2ARypMSsxPP+Ywrb
5Q2Mm1DPn36Id8QG9cXyedgqacAwEpcCxQGlQhOftgdviWCKc4k4RSWdL5mzav2o
8VXtbbz0kBkhDs2LXpmO3mSA73ojl1owdn50OYSKhDE4cwvypU073xmiMHuBy1h6
SiMCz9snmTLXidDcoGlV4LqzL4t7c7YKNR5hEWBqH53nAXGk5GShh5F+pbyx4ROK
iinXZEz0iszWqid8yYhVmUSlu9x5E5R02o8g/q6oJZTGU3cltoisBM7ccmUKyeoY
QFUzBCRdM942/9vFvgXG7jdnkD0J0XrDKxy2RZXvwdk0/c09z4ShT/ijjOjmxLyI
T5/xp5uBv4ckicDY/B6DRqnSt0B6uveV9ogbMdH8ARotoTRMLEO2NO91IBjaF1wH
goinub6WABv+PRnGhdF95/XNeKcT0nszEMBxiM3UsmZJwB0AdE9bYFecdQYpm03Z
8I7hxI7eY1V+RBwfv8X3Mt49r7UcEQHQj/5NT4+kzTJuwg9u6KfS5UqnqB++TTsh
fSOHIb0k51VBgnjRroRur/Sx8L/Z/R4Asjz9uxCKOsbdP9bTp/K2LPWbXqOYOg4j
Htb4pLhgXqOgoJvgxCHQz2aYkRMwd2I6NqJJDuvBaSDxlFBiQem3EOhGsGj8WXzJ
piy7aJ0a7r/wcw43ofmib6wMFp7DTD1CB5JcHAnt+o/2sTW8DanpMXmXTWNEcM+v
7Ti1DjZMMy9vlro79kA4uk8S3fRM7wpSMXoWVztglN4AFx63OTRTYzRLcHTlvxBh
V4otUvuyvQooat22kOd6+s/YT50o/ZajOTFER6bBhHZVxxaaxPgthOkmbSV80x6l
BTTg2wVimvQi6CTCFnlGH/htx5XjvqeKRr5Nwd/JqQIjqplZLW08xC38YPQ4N94P
msIyqeXTf+KzHDiIpyRLwZL0oidYXKs52EQ4BGv2IM64jwLezkNX6wTzXU+6OWE6
U9RBpVaGNp7+0E4Nvk/oFnIyZhLUeRd8j17z0bjk+6g9RK2Z9n25dJBFFEU8cmM4
HSiDZgYqQvKTjMIbNeAVKfTL9nZm427HntQ2Y6dlYWsjGlWwo8AvqhWLC8NXddyk
xM89WVLkY4qUzl9JxgT0CfVI3t98BW5Yo0AGI48keMAIQYcO72NGqhuMchKHLK+b
0U3NHkeFcUO2nhE1kVT/bZJkjql0n5ew8uKNlAz3DwQYDVUNl3zlvC37FSaW3Eso
LvsA8OAPWXrVzTm3K3tmGGpA8nWgyQg3llACtoPS/U0FCfZ6qwxzMeQvxkXjLXye
aTxLOlhavDmOikgnW8I0ej3+vrf4ak4oWKhuMlX10ErqXtyWX0HBm2LnERS5/5my
gOfwUKwuSM8uu5JFPvf+znl+8q7LYOkmRtv88Zu0Pq9DGNHJ5uOkYqT771iCdn0a
EzwnXN5CrmVHgZlzzlNoN5gvU4g7aFtYJD2ZLS9TlFL1P1tiqC/U7ON5jzUJRip8
tM4Y8Zi0EgLpmWkTKe0pZtsCmeesSZn9ir8/7rU40ZMIVgiIenYNlAxrClT2L3NH
O+i/Pny2TSuMGiX1gGQpNO0jy/MtODt/mRK/vE4BiS7/bBFGFRAXQ4YA+sqcqBgI
slR7C2TCfD5SE7Eq1MyutSlq7WALPo5H3G+DUnxgk/RXG3PER4TsfN+KPc37a4Ou
wV7UYRt7lnlfJXT2N4QCYdGXcKPkOf4e+kwHjSzLlR2tXmlt0uMskMnGZJ++cg2m
hLVwx5ZlA80nt2DTRK2pGZZhK6XKYALZ5/o0qu64TgsPhjexTHZ3UNUgf5t/YeIJ
zC6MabuuhJZG71OP9FvpI6Ov4pDLMCdl2Qc4cvJLEq8NyO3D3QP48rCR3OMyvthn
C9ibF2qfPCEu0sHAzy4shPMcDCPMcW8mA3eH4280UwGRfT4VvRyzMuK8Hg3uc/6b
yIDVbHx2MEiASowvqGTtJK/OjENxbX4gcQbtwxqm24yPWguZ1QRZFJCHqH9XblCU
y1rXVBoJ+9OR1t1dWe8dIZeAXNSJRT7KXxDhygDk0DYKfNSnV+J60ePRYgmct0LY
LldNuF8JiucHIZCdGR13kjYj3lxCQ67J07Tcb1Zc3mlnYRfRqNm2hQTYrT25oZe1
LobBh5o0VAmq0Qk2DFxyhfJnxkWJOyTLyq7BFJ2jibdfEZvkZdzqukIRttvsibOv
sQ/5v2TCtzbb4GZaV78j5nT7VtQHiGVEWMHW82f0HqUFh/ed5yinCwmjGQeoiyX4
Jjle9VQwlN9dWyyUo1vk+lgUYNzrHGeFlinZ1VtmzKB0hNbfJuG/BxGwLaj4EuZW
/TKir7viUweWMKtU+ID7psml1XhHTqpMTewGlpathiAnmoKKsTnl8lg6S+xFZp5N
RlocE08klmkeaG8ei1nkvajESIBlyvtfn5OZWgAT/Bv7bl2T6IreH326d0qYAv55
w8zj2IRHwLrE3hG3XT6sUnewDnZavjTHzNik9fVtgBf/YPZiRZ9EGhoa0u84Sudz
pEj10wJ7ERJpYtVLqIX+0A9Zvl55nHB/2HPLcEZxJurgQLcC1fz/XbtdT5se2eGA
cyX0ULRSNrhq5NDLDDKaVHiEJMUjjjpC/aQvOTJuiZEXzaOuwu9Meu+yyS51XXU+
GryhmCseYnyFiTBoVI3RrbcU4M3SH6/x4rXnOVmuY6wUM9ypiwJP6ok5ZEeaDOaS
TydBz4TrnN4YjL88niA0R3GHfZNvdyMrBhVZl2wYO7EjKYbDrP+uByU4FZknj5fz
YkAg8nMIUfBaUhswb7SbCNi3jo830mck+AYAtiQ/c+uAzq/MZAy9R8Q/t1+8wAIw
gpSCmwaPm+kZ1gNYOSVdCM43q8gLJJPdYq5sPXW5GnnGAlV8+ZmFJIypOQk2FHCG
sSPJg4Ru0wq4G3gK5EG3kF6A1SOGwXAz7tVdwITn/EvaAGRrLGtFRJTChTzsEXmN
B3R/fiHarN8TfU98wnSbJjE+H4dg8fJ7E37rXCVFKxgI1ZjjcmtusSZa/8StjgKH
3nbvULRYRv5k1oDXE+fn99TmnTzEfR50N6gLB4mlXeD62Aw01rxwmdyib9rdFSpn
ZX58rdbOFoWWE7MUubZ++F/plpOh/RMyKnUVy+JpfNxpoEBREh0XyDtaoktgddjD
Gjo7nqsT7GX8yh/cPFJzPSXaBhNlvmu96SRQ8/R7j8jxabTCZHBdDBdbOKzBjla1
29+FxqQ2iWP86K4/jGdAHtSvdKoZeyzYGqO8ssppK8U+LqDNLNtCoCsYz7vQRVae
1nlhOOBgpJIbHe3kup/OrN3Hxpk+5VP0JtSadHlqOijxpUqk37tqE3/VgD1Avqmu
udxL02cJFt/ZBtYS/uG4h/okAPbFW/3GBnfQtF/LylOuOOsVd9hwlCwj0xxdAnq+
ozNXPIQFXKsLXvS1Ddhz/ELgTcWlUo+zRthhYiv80M/uC/iVUNdRwzPj39Lw8B2g
/YUoIcm+aaopOjObxQb46XWt3i9NW+hxjFMFWcIIpdpH2dH2DUpdmRQCTgg6pmHk
ko2RyfvtosfurfddBjygY2XyiSUh0S9cevP2OPSSEH/skZfWJ0fdvIiwOIoB6Cpn
NOzOsNhBlhYXZ9HciPAzk9eRYElxrLgSonRyPE+kTKlKMOZBix8MG5vDmKL9krFi
aBKQC79z1jRbn5xH1tGUHoEmsoGRM/mSpeRQ9hD0BZ0FA4bcDsA+MWdEtgu65cJq
863oH65P/UqCU6uzCmENMtl+Fjvo3eM/NCwormgnM8ZXkrBPmJSErkUUwMu6UyGg
JpDTDjGweKGnZQZo1I3HMu5sOlrDWVuLy8JaKjMsY7AV3xE2wSFTYKhuKQ9JvprJ
A9RcwhQKA+fCtIyjrg3JHLLdetPO63uAuSJ6mMSFPK6yi5Sdl0mVexvapnYWLpjO
En+clo+KluSh/FM/rvBxfiGOEDA3aWTFDPUH9vjRzFPlLCZxspuqirz4FulGgVwl
An7nxN3uUoSHdLjCC1KrrWM9w39Wjdql6jpb3VAQFOgbRX+hJg1GWUFRuLty33+R
DCYBIPAt6egDYvvWEWu1ePjfl6tu5DEpZybQvNNz3FGkYmCNxTGTGPko2kghaPXb
LN7lwomkC+xx/a//28cQ2euKm0qAow5BgTy8qUJv7uT/PRdkGC/0SOtRlFQJb9kx
/01mFE0Ysw/cHgUVpgH3dAWO+lF0lhCLxVTd1XNIgwUCnyAdh4BpfEt8mjSAi0y4
rrEk6MBrHOEJfiF6NFonaxTXKVZTwJfEtmQaGcy7FjQWMOVTcah8HjRvF2SCi3h9
ckstPnC/ySZ1uw2RN7h5kaUuCWUlCfuuBMx7YVq0gJsdVu8wcY4jEKgYlmFjBEQ2
lBeTsPUWjjkjFZc8V56Zmjf50wGRJJYOdDN+ueFkAfXwEaAcs3NjeGVxr9sFKZbl
nEd+OoizlH7VAp7aB5DTggDzTzjJSKWoBrh3GaONsChbMZMMDDO4sKFN24XOMjUF
KXbxRsMo8SlaCdJgVbYL5u7mdPrmGmsNf//rjbJofaV9ATLB05K9zhc93C5cvxPz
lrnCNgTreh78s9ENlRdUfwNVU9ksewzq1PuuUg+C62t4iJItmsG2ygJs4zvOaPaY
CNLXoLQ+CvCusuPhrR/sP4e9lFcxSJjBIvD/srnCoj1DJfDlQv1DWzY0yc2Mc6Vo
06iBfeTWiIWKEBtP1l3QEnGQy/MP8IYTemi9VVzRHuuNnW/n921nkq0y0LpKXIo6
N7J8gTgqOO3HkHkf6P30JtBEbKlIwBO14LCsaUUOb28pQHcm+YxyFTrGffL1Oaha
/R2XbSR8zndnv/DYs/LwU9w9VcriKGTKPLxZ1KRiqnyKWtahs7Q4oLHde+dACcKq
YDity0queJCVi4cKY9JszcrBQjpMrH17hrDJHHg84JMj5RZzc48lCpK2lfY73aMk
cUBTshwE8cTDYPYQkEUpg340Z/ZNpkwQ4uM+YNKHwCt/HvzVAY4SZDXjjSlQIcqy
3+P0zPGwzsr0LkiKR8IC0gL8nylRgltuWtlULgOOvTrRzXAtmcK5fjgGi5RmpRfH
C+jfyA42eX8YggcMz9le3KxCithRteoO0Jk/MGKEFHxBnSX3tHN+IfZ0AfA/hf+w
J1iSY6yUK9l1FHMr+QIzIJfQJmk/+iN13FcQMfLaUpGvWsZodBmlmNP7SXMJElzf
gx/v4yw4kCQUXVOLgjp1UeUtb88AVBWhm3iZqcRScjvs6y1x34rLhwha5ZU4Ay8N
Yp77lCBGfiofpWd0sfMXfc/CNLDUTLqy13AVfAn0P3reov+SnuGBAteujeY+C7pm
uql8X7KQzHL5/5oGHSKiFOKCdKPx0dbxGo2ohKJ6pIJfE7IDR2b0wU11leLNpeLW
qyjRQPcmYTc2Bo2giBWgsz00OE63XYsV7+FS9RyFL/XjCrnfOgvZVGoPwPGb49I6
YTkEN7EjE7wPn+k/WoEPBR0RJUnSlEKlINwxVNH20dQImp+KJ1KMOZqiMson17S2
VJ4KjAdITPEm2V8nc1IDJwLiVT8BwHoGOMaEPiCkXtOFjVG/hGeYGVrnVGToEzSY
UiSeyC0H5upKhMJTQ20tjzhGWIQhNh1ZLHCavI0r5J0aW5aWfi27NocC03KMQozH
sfsiYz4lWrRQUhYnAMoXP/bwFRhvNJBzefHkiYObx3CNmlT5fnEgNteNGXeUzjKy
2AnSd1RCLMfA0e9HP5qRbo+1MIh1ixJJFT7xuV1M4Un8vf/kvYnVTWdfjaKjA19K
zirbbwjOV+pp5krvYNO/snVM/O5iCmdgXD5jyn4abJG25oTPck2USfpLZ7xMSuRR
ygLoV7HLZOP5J5FqmAlAhKbX4/FENiJCQoWX+VoxyK7xpJtudVKl6Ux8yh9HLXxv
EE5RSAJbsKypsxtOvAcVVMD31WjU84mt714zseWX6affkusP3KJiZtDnzPuDJjzf
V5hylqAbAqLkZxd1dAx0fUAEwmJPES/dTHkuz3W/rdTHz63V009ddITIvvsALwjc
VMRHqt6QHiXzfBDY2dRbrlMlhKtzrUI4w0dqDRcSxqX1MRmnRpMfs0v7uZWflDSr
xoHwz2zg56C5py8fc2GyarD1B2ENwsQRV4Iel99N48KLD+i9bGs5+3jz+cYLlbHK
BAj3a5HimF/C9CxjzcmF04I3iUA6Qx6d7Jhlzh8pWZx0H5314njwmm/kqwYZ7pfV
iQxWNGzpuec3fHdeYbKq1TpgHa2iqhPAQOfRn12MGy/9W3/VFmrck1lLEIwyqf8v
6vowpIl+fuxJtPmPqn1koOa/OGIww82+vgztxl9890IAyJhq/sJpBKAMLZhs0PFP
PwYv4NqoiNHL28r0Hb4DBWtDvez6XExHPEo5lMcxbl6NoJE2T4aJBndLd0i2OJR3
JfZ4CrDU8H5GZ9CCDpZC9Gg+AJ4eb0VfajGeOfOASNYzUPyv8LDE4Hy51kh8TnY+
D50GOTgQJZ+Lj8svx4o76etM6kBSN4fqimd7QAqJl5VcSlOIE679xFfo3lj2BhH3
hyang7vVUP7rgm/GQTcrBergUaFO85Cc9l6Ao0kU/KfCcMqqpMctS3SYpoNgt9D5
0EKy2WQFZhPbZEzfdTofs+LDqSCGGv6KEUBSAb9Yf01sx0TVf38F/lOXZMvCFVba
zeKMwjcRwNBnW0b0bXzKFzjuZuxVLmGO+L/DNCv2WGR20080dKyM+lYSq6ysw3jo
x8quQNsWgg8QvOxN1ej6+Vgm1/83D5TJiOGpbL3yY9kUtRe+uNiZvqFfg4VInKKs
elTL5IoUN3kHbZPdS2wf7DWHsLJc70+0EVIm5R/lHiGBPhZXgy9HHTmL84xUeO0a
o4WFN1EGF9BZTd3iSLJpD6eOG0ZP19xnYB20kNIy+1bQ+3kyhmPCE2DQA+LSczHT
dnOfzY4WzkI7BlWuIE5RIf2IlhHCHuqVxzHcO5aqUVW6ANLX6Z3hVOyWjuZfDixQ
+mkitYThuBlMpfcN/puyTON6LLmtLI3jn+1CiRuDECR0H5doyRQtw+Coo+qwUw7f
HBecvUAVgYaa7H8cDqgoMtdJ9k2McYdf0YdI7R+T90m4v3jU9AJC5qpgrX2DFnRw
uov65SwZ5soazgXVaznWuMj0USmOZ18LQLL5zeteujE0cyY3nKukA+La0ahXIgkv
Fdfuo/YmKds9o/0v6Dp5iYUinQb/j3yBGCq3Ucax8DdkKEIAG0jgzpJ2zrwhxkCy
e67x8GcimZuRz/tyhkOP6JD7fCk59BnaCTZgZq8edzSwSg76k+osNOI1s3XORWbl
fdt2gD49AH2ihd6cyq9UaQXNHu3NOsE1YQc4gyiYRtUnCWIk4lIALuWdc/Si92Id
L6Svc4kLWT9z20fIGb9NfXc7Q1RmesJsyM9k4bcbL/Sq4qX834ZWQYGqt5jOSd8H
DuQQV0V1yArLRv748sYu0uP7X5jk7lq/eFA/uVKQdnLxiLL0bxBe9XemWDJH8nrW
Dq+V0nl4pzdxZZACNGICtQf8mWWghkzsOBQyEhiYo64AyYYe4DIyUq0HMyHYm4/e
EJqYMy9M3WDNPk8RICs+meGtKowFyDm2So4WPhRQcG5/sBK556V3Tj1G2AKrVGC8
Uus1KzTHgeY6FA23n/2H92abGPKzOfJ4h1obeSj9/Km1YpR3kdw1iqL6vyjZBGE8
pmSKTM1kQJ46gzQ7Cy4Qhcm0VCi4w1wHl3eSbBlEYc3yfFRtjjj/dnkf6bfC/NJE
OEY7UQlnSQsf50uE2Ggq+f0CN7HmRkEnxTBe9zbv6rWVD3ig7SxLZVdpLTbG4/tF
ht2eJPniG90gqXdxjIyr7VByBgJ+RlKhx1BCXevfNfZXqYL78KBreMWAR9240CAL
R9kEnVQLdI17E8ruJ7/oY/15JO0s+3M4A3iRY4WinNXmTQXw0m1yhY2w0gptudCr
QcaGSgNUN2E2NJBgVwlaW8wtmjTQL1RhPwt6/xu+Dkmyq2tS2XvAAh61ObfyUWXx
WhP+R40mpTA5BaU2E9HuG8iW8c4ghqvy19nzHdsZOK9Sz39eWBfOilbYzbSZ/RME
v4x/BbySiz+t0gQv6pw/Cai+foF/X/9LXXSgKR3YiMT5s6f8eD6oELJoc2JkACMn
HdCUN0rRb/8EPQvqiAJ91rFOla07o0Doec6TiR2eBn1E8YuyU9fQj3HdWIttPodr
ivAk1NRormJm9AQgvW3euiVQuIR8SvaUdjeqQqukt0T7Rjan49Wh/OsPiSArPRJH
N/L8lHWN1OznP1HsK1CinPYS8CHh5VXKq7M90+JLLIXcmxCCXlpHD5VKq0wT05Xz
6q9qdjBiLRLsT5HH3W3st+WB3BFBVIB+pi4ZjxIM3sU8K00s5HvJqP3o5mlW6Qbs
wddOuW/b3VGWXcFrWuboHFkYWASr+XH4ReH96axa0ZBBZcQPufOjvsMglUTHF+U6
/c4pEeuis1S3BmkF8YDeyc/Eh94tw9w3ij2UrX/jICwd9Glna4uEZNp5uHpaqk4o
VkMtRf0TwPrl1Mksm5EUOjc0VkaWha+z+Dwgg9eUSr+QF/CboYyKe7mdsrHY2T6k
ebtEz1NFW1mWEgIRpRdNIrzXqRCXFQESW+ks6D2Fhuu6vUnFMtIVX/8ADfezzbJd
R2m5arK7GAHv6NvbFUD6p1lWlvwjwHMh/h8KT2+XMOWHCoJ7jU/cj2hrR1J81QvT
m6d3R//nOe4TBUV/sDdL2dLtrm8Y6se2K816QI4AnLQBbg8Ku7EQeO6o5E/ONFXR
QrnFq8sTjb4WHgPh7Qeido73EgDihEDP+HhsjHxQ+3/V+TSsR20bUqyvW+1dav71
We9V6bQk6hjjzrdegsGIbrsWYNzTvZUTHxETl/7LAmAJUB6A/+xK+3Umy4rYXQKU
ZgVTL30r3IDabXt9Gwy4/yVEaQ+wE29oJgqzyvnxcbHgS77FEHit9pRh0EaKjdko
xdtJqlsk6aYk3joEYIs/gYYUFOANOPKq4F++CJ9UeNiPAVoCRYuI6mdesdvtFGxt
UyukAeaLikDEkp7Tz+9qPKRE1i8yWj8aAMIojZl2JC/1zKdFLxai22g/hPUNbOzt
ng1UTBLmD3njlVgftHxa4q1fE3Nxw2m6LQqavp/tJMD5UpaWsEvRI8JHlWpKaxUi
0mqS362vodAH4UCvEpU7cHvAj3o9kqTQ17plDu8AYR64cHDItCs9IhNfouNUIjdx
FXc25O6XiuDqB/XOuvlWXPkZLu0FeundmmYgjYXq5xFTyiSW314N7ioEFCzJRxce
s/EJO9xtPmYWWZz6ju7HIpU6BT3vUwanwW1G+3mQkLhqPsZCGuCF48/ZHDls7MO0
nqgwuaQXL3QVz1MzU4xfdQ2jbUgcO+b5bR/AkgR0ddoelO2Ak8B1VbCBCvJKFE0B
+9Fgq+wOhbZeSru9GzXc3owDoCivxJh2a8liqJW6qKknjB1+N2UX389Px2+p6A33
E6lavCXJRgpCC1MxUFkWDw+teq8sZaNt9ZsdI/Vgs3+8xjsOSlbmfVUBZDeKSl5K
O3INRTOr1Eq3glG3CM/QQclP41ydnYJgyjeLCbG10+OqKSjV8GHsDzVytctefTuZ
EJwfQDixcBtQAk7v5EwJqPujCwD1MRJW9J1seFAZpgvQat46HSzr3J+/kjLZi/MF
m92gJt/I0CC9rM+WDbr/EwEnGHAuNMiUsQ5OPv0XN4qO7T0YdiEGUFWxjVSR74/a
0mJYeH2cseYetOky6/gQgdWfPuWWsB3Bd4MGfqWP/KMUYQmftUEn/bncKpFel99A
sIxaHdNgkXUed4fEPsZIzPvg7n82dOiWevMpVZLhjOFVHG3vxiFuHhAGPACXWwo/
wbiKNLTqGNsKUCZ05mHgFf9rdN8NuWpc2TCIcQn6ulsWlBm4ufzcMmhj03XkaZrh
uqx+9Q5WZ9WrwUdhbZ64dkRNChat756eIFJQpn8pC2kV/Fb2I9mxzGLIJqtdtKjs
EZ8XUIJe/qO2+zjxEvB40dSW+y8cTbJhGSZCIt/Dxl54GTBOP9kuW5d65hz4v1Se
G4wLHYaBrvEeT1Q0xvUM1Y0aV0maEaJuYorVNdQv8w3iBVYtmhnqbvlZ9ge2KVe3
X4wth9iKWFTXF5tINDtNQycF+trMmfnAmwfoGXDkTcvVlzn7spubgKw0mjddCwD5
pxKnIICza5RLEo5mDRj7SKnl9MZ8CBeIdJi35F82Yvg1IVE6NmjT+CoCXJmCPAKv
JWtEYYeklBC4G24JJe6KVBF9s4Msa3IbLb1BZPm7nygd0ZXPannSPEjhZvK2XHr/
e2CImdsJkrrjhvVp3l1RrDTdS3k5glqSs/ZQJTxRb5Cgb5J1IiCSAIt6B0gwQ6uH
9Ozmgf2P6JeduD291p0EMWPA/pPKtNoLTRTNyDxFTJBuK4hEW1Kj7Oqo8ehpK+g+
KFVHNTuhtXgNP6p+jswxRb6hPMum3F49A2ytOq6SpHg7Cw9yiAUihON6EGdU+jWq
RFkssYxi9D1mW27S8CeWDI295tXQdixkeIUXzlCfR1IwkHgDIHNP5LnjLddVmSyl
7zGExXtpnYzjSX6/2ZWphKiaSTK5uJhoA+egvy1Mpf8RMGkGNET9LaCzBWxrvzGf
QsqxFgi/HAX7nWFK/Kh66plJggt9i/ZhQvFmgbjyg0dclKNLykv7xUM1C2E05TFn
yRl31vC4lrZzU/AuTGlstGgImezFyCNXySGXzpan3+pZz+8VpMtDZ6n5fQJWSSLH
xLOp4J/0MKOSUJOeA4vqJdgUo+0BkEndX49TeonvC2DYNpzya/BxhK5ClSkJvH87
UbIRvUQc/oO7mWrwzHN98H5ltohAojNL8OIyaDoCzYhu3m5v3RwpxJmWQ2zWtq8v
xSQY1pK05wWk6xjBsrCO4OAwGqd75F8WuNL1Fe8WJAQfgMMYInkNYd0HtFSSbExz
ImI5zJyUWdoNUm5tU9Hd8+/D9oOe8XFBks6weaz5noAH5mesZHl7pRYK5gxqpBSE
BUDcMqcfeIC9LnQGm2dUjLkzeCAzX0EHUz28PApXV7jzmsvNzr/Yj6Plg0r+XmNy
igh/HSw8K2vU6lu3eXLQ+D19UFA0I42QL29VFO88t8YqwXNACCr9L3mqyXvHh3RW
p7Uk0/r19BMhU2lfTti+/G+p6ItRwHcAricvX57t7hDOQ2+4v7M/6JTIrYc4fgm+
6WzXRLY89xja/QpnN+RCyr+FgqYgyYxNgJhkwaK6UbAvK0mJM+dADV3D/KNpD0zQ
X+fQjatCLN5gW+xzmXijryIeSA8seKOz/q7Ljw/9ILjjGebjaQvWO5WyVtr3D8pW
ywTtM9M8mmbMoCESusOrOI2Zt7rlg6HUw5MheczjnnjYO9k969p/3t16xKq1KOIL
aN9+790kBc+SGOcOuBrm76/1gQy/k5SB1bOi3+HHSFWIUt2TePUqP9+uhiUsfmjT
+FX3GIR4nbMwfHFjZml86v7m0c9Z3K65K3TKPfSQ2QIZwLMTOr9j/gGHSGpmpB64
WAI786NlRy9tRbURykg4TDPfFb8vhba8unheHbnWZq8VcPaQivdCzz2xVqTQKVYd
bJ21gcbjhHHnPPMpxOCfpZBePnnONUEw3CMZnGoi5ln3WgS+9U9dGP5ObAbUjjk0
am3lvvPn3lwmXsOSOQnHBYL6ceU1tqqyC/SnrB0sa7moySd3QkBfbxXLs6vHhfYw
V+D2x6/gvMdFMJGmTYB1HjkZR4khHAIlSbDqnfAee4Ovi2EmfLI1P2HDeavvcvaQ
2GLKsT6tzI47dGgbNaaTc8bIQQ2A2aQcr1vQ2dz+mShrKzJenC8j7qg+X19ygRJ0
MbJSonL+txeMqQZ7PMOKONyMkwOmwK71niwUi2Fb+5fLMHIRgeRnbYEaOLhWTEIe
gv53/nSpxo98xhUtV5lJSY0qTQhJoZ67HiFCm2H082iLx0GamFubypbx33OxsfE5
lOai/SAjmZMSMdx7FGSxCR8zLlHd4kPFYuZJBAIw3FayP8hNQM6+Vk8T39w2lQKa
Dv5GUuZMbc4Wx185WSWE/5kHiw9HIpmr9GUPZK4BBjXaQzrQEBWTzsqluWILFKOp
fN3d335Z05MgqHXX00bLeC8ycJBCpA74A3MkonxsxWtr2HiNGb9RyFQ3Myd8TBGU
Egm9+zME67Gsq5u+H3EmwEZ7R7+tXBF9fZ7CsFveWq3wA3bVpS1p91kxLsGWM9PX
5N7Qb56PJX7/KR50K7MKdTpMk9SV5jKyb0x5bCf1jdQ4qcO1p0rpw88ejPO0PJsC
Vc3TBoQDdjuJ37WjGmRQJGfkjtMHLFK2SR6fWoTRUHz4WxP+xqAaSBRjz44tB4dm
GB45q55R/jMR1ku+upl9SwN0Onr0uDYByxaq0PwMB47IDZ7HAYVxzn1oMK084/sh
U6VXWmf0G/W6Oif1awgWu9WxMvXBtuK8OFWdmelW57REfMouV2AnHiA6fmTEp6x9
t0ZcfOwX4ALd7Pd8oxR5Iqw1sC0yNk/8cMM2q3zKOiOF3ofz268O5lOW/2VuscPz
C6N5rfBETOs2rn03fjKSEBOyLLvX0THFoBUtV3ZDq7SrfueVwtzAhIS7z+7Hjo2+
AWkSoPiju7uoIeBp1aSWY/N82oQcARRM3qey3nyX/3iioOSiaS5Syv9P0HCrmPm3
ON/AhgMf8cE59Ygi563EFqyrP35C9uaq+yzlQ3pn9UMI3t0ryODFaQ8kntWa1/ew
/E6j35LbFoTGszLci+oDnZLy4K0wH5ZsgTKQRaBqaI8lff2lLyE8wTfX8/cSIY2a
dH7mj+/fqFzJkftVKIkvhkRfzB7TQozEHe7/JgUOJv3xWE4a8YI1pQBaQ+bGnH33
R7VKfISiT+7SA4Njj1ZI5aSAvEEchIzyDVpzRkxpbEk8BD4R4q6cbPQwkuqQIASy
ewZ8nMGp9glywyhQ5wabe6yBzETrDA2qOa6ir2Y6ejq3oupyqfRUZIMQqfzSy7AX
cz8dIwmxRm1z1UVCjbB6Zc/A5IbFxeUmmLN9mXPC9H9nZ6P9aBLP1Hqre7ZmbAQH
MhtvYjJlM49PNzx3jAphTLDZn/sbeFIhfKH8Ohn++b230+KA6/at8p3e85Ct/4SE
al19wahZd9nWLEYwsbSeWKIwPdy6Pv6N/dd9MFWIW44MjkqLwdwmmcxN1ZxCkphc
+2SZE+3zKY4shP7EMCBAxvj/ELGeiTmMgBmPWeIrOEGlGVXkeV+e5Kdz+v5uYgLj
EwfxjXu/EfBd940p5B08n3QqocIIG9zbtZIRmg9b+OgbwHiKXzjUVeeFmQwx3H78
wbmnSf6i81SlSAYYKZW9PP/+7rt9d5sXL0qXG5s1EsW6GT4E+rz171Rf/rFgtToY
fOF8Q6qjjLCFzGRCFPQvvP4GmMf0HcBgHTeiaQsNRvi/KrblizJXScN2QwgS6mtd
Cki9gFYIfdhBAYSx83N71cqnlhdtm5KmU3/XjlyE68GFJkuAZrVuw4TJlNCnoq1l
P/LkPVOpZfymhCkigzoDA2oQIfJyJu5tgI5hoa1AJ9tWPZ8AIV+VsCfQDmTTD1lx
5RwOuTaoUqD6t0GgsQLi+lPhx5LNIUFodeBAt11wC0XxBMT3cIhbWkC63tRVdTZ5
L5ef0+q0AJQpzsSJeS4+/tJ0ToBF8TfJ8TSXGvvv0+rc9XkX0eEShgC7Yjg/KJWE
fzWFQ2cyVUu7Mjl7S2BUPkabuTEIVtg+niNbk1ylzyHt7N1Z1xcPX+RfUZNQlTYZ
FehGPjB+VKhjtd+j8ZJrDQXyuKQaucC42SPT47pFRcNnTlLpKYRa1m2Pfvrk/mPm
HS+zX0x88E2aKItxkMZwsJjNXBqcHig7HaD944GRCSOullttG707mD5AOyFpqkcN
YZEsqCawvF2jJR6BZFQ8mQdYMPOeQLxVof3hdPvbsn9nw6nNJQmCGUPb2Y1cU1Cv
06DMcxGTPFmBZqb1/0dIHgCe/jmXzTgglEwCCDqEoxlfy5/xvzTPP+IwZQBuv+06
LzofE2YuwzlhBArROuiEpsf+u6XaXlQwNwAgSnJrzFU769nJDDgUiCeUwBgFlrcd
pARXmjnI1UCHFIOzJwQJToC+fsnm7VzxE4egJwyf1zWjefJFFk7AoM6re0NYySvp
QZSnkrb8j0LR0724xUr96zBGtIn8aeLK54xvbixRINIKmfOsQYGQWMR59s2BZwSE
5lTFGdiZUJSf2w5EFkaUwqwsut3SapHyIDRDoU0P4ZbcSkjfYD1d6DC8l89qZtmH
cpV8gBLrHLxoxNnRzxnKEJgHsHkGRFsZz8gUXpxnKQ1rl7tYvHobsETOpCgQlBtw
azn4YDvvPWF8qkAM+wl6EcW5I7CK0Q3UzvrvyVzKPZR0wUtAmSJv4L4eudzSoZ3d
lLDSiU3vn3a4m0hELQ0jn/o3Yef49Gsag/5k5vTnPhRuD9TrPrDWz5wdVvcPPA1g
VM9hI6NtT1oyXR9sTg+1i3OUxLTSf0WtZm/e9vbifJ9P8dZ1b1yjcoeaW5NFsHjD
mepxCS0O4vkK0I1QEH5D5GxNbWSRH0h30gVy6LRUTZejm76QXl2+20cjLndnkeoa
GEgYsjKnp6XBWw2tyY6ZminQ/L5K+DeyrE6N9AX1EoVcAbVHES8JZNUsWPp2fF/3
a0yL+1cv4JF+bxFeH7B6bMrzOHId5aD03kwhZuKXbUcPcyMse5v8x1gd7Dj66Jpl
H4SbjaeAaXFVg6qtEWpTZihvYtEsT3QUutMIxvZif7GMQixGgfcbfv8ilZ/w+ypu
Dml0iaCQkDCMbqTB/5YhN9Wg8vdZB3c+wo1GPwLvkuQe0o049XSyitNL72dRaENN
yObuSQL+4Z574ILGoRDrgTo6LI9rlKfh7YT7B9oIANFqtkwvtlZ+BmW0WRyQg2nx
BMw45R2zwAvne8YDGWKcWRNK1BjhBSvx9X0GkQbv7dAeUDdhDOkCbKZJRKxdARaQ
X8THM8PXFnbz6sACH1gqnlbgKYLMarG4y8WMsbDyPLS9UrzULUCrcewXcV7tZx2j
healffbEDLXh6GazCYrK1R9LbjP0S3SORafztBI6rGGwATu60Ctb9vCaQSUeelFI
rtlq+8IEn/q9AGnKpmRJ6GrJClvNzEfl8+NYJ86DMuqXeq9yZIH2X6tdHocykmAZ
5Zz5RYCxzp+DUfaH7bdzXBp4hU8Kh/WJyjU3c935OcpaFPyBgNiq6SZt7lcw/aFj
EufVmz6tyfWym1Hpjd0qN9BJm0Gzm7z4cXX4qQ1el29PkqK9+1e6HBzW0lu0TWyE
LOAVbBoy4cNKdeW2Xm1cXRmsd217Y5lgv6kV/+Hp9f0sprvHvaL9ce6JvdYFXCjV
V5yKqQKtuGiv8c8rDkoHMvCSeX1R4G+6nz4nzCH4fVxcxV4gpTFGe3RKJ4xcMcLF
0YBcIPfdc9pZLrMwYtr3IkHXg3h/x5YgWgTfeRM41atSi8VFEsk2Ds/WB9e+s1tF
p8E/Ct1foKs55ZlYcbTjzt9DImkIzhu+sUeJyN02MQJH3kknU1rnRqDutPScOfPF
SUA6qQzu0kK1vch7sLn3/d3/k6sk39aIjTdJ7/oIirAitKB3FwFQEofBvo+8X4ya
RZu3yjxFlFn6wbdT4GRO8+rWtnvqq33RtHr4WNAZIyMdK9nKK50slEEoU+zruwv5
F5FQg2uwSOb7plEmy5IlLaVc8C1HLiVS8zI5LzMtgN3LPcv5gpqSvvRj1x6c7c2U
ANGVfTdoKRZcIB5zGCz0Kt+D+nc0ekETg+65RyxMzaLVPGoHMycrS9TIDmQbJrr6
G49KPmbZRCtFakHQN6bxn9/wezsf33brdqGc+i54ZAtfTBusyX6VtxAZeG28LGMe
wSFRiA6xSaG4CJVndEpZt4YqZgprdT3/UJKz0Cy/N4mjTcgsvCRC/2FCju6wHu1j
z5el3FDkTpJlW7pbReD+h51P3PpjIiNJsR6ytPU74GUU/53THLermnLMHstI0XX6
9fLs25nZUOCvmQ3GWxPC1McmLuo7znioXjn5bElVwv8FPY9UwoZzKLnchT598kzY
HlC18thiTvO6vE8Cgtg45TNdMmUbRDxhc0mQrt5xCtzkSwquC+vJrYfNZ8tSQBgi
TrFjATg7Xcq5ArpW+7/rlnKiJS1E+BGZVi+jBMMCPN9dM+6AJ6Pxiiyd0xmKVu32
xQEH4BcVmFq9aFVUzfYlXeXAPWyPj79suHtpc3ESG3nNw7T8Uv327FiROwo4a9pu
IAtu5Wef7DeRU96r+pqBc4WcQHcQ+mv0sZxL0K6/byU7R4vdhn3hqWfZ2mu2sawR
A9IOkwFv3xZH0Pk5b7XGCBGyEcf0wbYmv2xuqbQwUVtaOdjS230t9zTWdFhpQ2wI
wXL5lWOuHy0sy0Na/Z4yKXuR3LVFjqoe00MMdKSP4D3APae7Y4TAr+jOeYIDMMG7
TN4MfAihkc0GI2+CxV5w4s861o+E7u2r3nCHCIlcWqVVxUdtsZ3I1T5KN+BGjBvD
WGSaQR+qExwR9Eq2HOXYNkw5IHNmzpbeELRCkCwuUjjZ+aCEeV1bATec0pnR8t1Q
PHyzwu2w54TjUOsKw5pa7lpNItK9/BLyDPFsdGlCcUQrSRvq1ELBnnsjNgHDTq8a
tmqi0SMfK1zzeTOkqTzumAiYSnF+Z8SQgYjuuup1J8m8wSTxTpVv3vDoVXHiov9v
GSFfLQo81mpy0SwO9evTrNhGDat+zIEbKT3LRhMJqvMLSWc/bIdF40IyE9dKBJtk
AbQJPrJTFK8FYbXpUUfjjWn5gbRugOK0f4XdNSQUFfPhP+RU49aVbmxEHGhoY4g1
fnuvtIUS9XYb/EDc9Gbml8IECbSfihu136+xqiOWYqWWGM3S24pu/hlCkWzbVuJ9
L6RSWV/x8nmaQtWewyp+3bo0iKeCClxqnWDfVE2qSOPYwmuxTCIDNvfM9nACMmEd
PV4J1LuRMiJlKegXtlCk0r41x77gYvTZhny1lvTCISBacsi0esi8jFXP4GkkD0W7
tHfj56eU1fAcgJ9yyPH/sK9Jah7zeNG3kCEOS+SwT2LNeuSJw1tFMJmKO+BHBxdq
uzCNuIEiEkYiQnoWUrSqMoIT5ETxUThE9/pvBfdc0Cmw7cVaalqnGfZzQGJrHaxx
0MK7r17A/cqdEDzCR+6+Bdco+4s8bLIOsEhhP+F30ekGTlXipS1dzUNjR/UxkSEK
awqCh0dwn803wYsvmJp99QSpy13SMIcqGRUURUf34lZiOscym4Mod34H4826CEJe
yoWFjVx/Kgy+hx6mnwLxKxD1B7LKl2MpjG11K1xgNeM3Q4aGKwg8XY+n6Gw10FBs
kV7inWKGq/Tj0dmno2QZ/oUN4qESDN99NWWymSgeQhfi+HIHPcFizVrE/HHYSWAu
XC8o/MPnNCOY9vDqt2TCLFHRJfywoZu1cgYNw02oMavdvtG0K7ZpoTwkWR5OrFQb
2moe6QrYBfmLtOPh+GwhTat/LaqdxRxUXj2EJ4jVyYA5oSiBOKmWljDcoPQDLsWo
7pHaVLTuQkVNdMm53Mv80Avj81CmhFDtogCeoRFIpnP+i0NIflGDQm7W7ojP2DTs
BNWz6oLasghLEvB+217jSzvnQmrsDfqXsdzsyI0B8vhIa+s+GOwQQqg9XakTud2B
HlCNhs9l+PaA0utWtVzkFqUC+3Lr7Q3wkqD38/DW10KKVgVscyjj0R3yDk/c61gu
e3qSM/WlPeN9fzdYE3MJ/LMzrvG/SmCI4o4AOFdmbWZbLxeP45JmjJNZvO73fkwQ
277WoPARjA0sjutQehygJIabRYPz9MoSqpJxrNbLWEdAMLhG6yoxUcsdL+KucuYd
AiFgmIPGGvDb/VNj4/rtNKSpft0FI0B2VJiUit7iYWEg19bwmdrMjqhoxwArAgnC
wYu/GcFnjSi60ERVgW5bq/iO3wNAjczlS6lEW73RkAxUKnLUgRvCRdeQudyJvN/a
10htagx8nWj6MLcEbKyPZLV4U1LfJSpmPy6kNyQwuKE9kZ9PRbMZWqZ/GbAhcXCh
HOwFGtLQ1P07mChi9kgN++FP16dNN7B0WY/q+eDABKhP5/Ul5/EJOBk5slDvD9WB
v5yfhj6C+OxbV9AummQjF001HjulZ0Urlh6zfKQWkamB5Zb6hS2WFy99JMOQkO9l
B1Io1Ec6CIPNPrhJGQzs3rKB5899J6VvG94lfm2kV/QRFzwmB7D97D+u7HfOm+ah
on+vlXqsmXlhfABwJ1uEr5+qZtVunJ5MOewOpDRdm12uNYj+EwQSDk1JyafZNQbO
KG3HAJ2+o/sbsF+qfrNqNwClSmrQLAxAudRMnZUCREcB+LEl02yMnnr//jFxPvNv
SuaaaraaGj6xrvNwswVDS6dVgQqsQOStw57UZp9jZCR6oP/qtWrUm5/UdXMp3bc3
9HJwFKdWKizv0rcKN4nBL9ArvuWWkay/qq90yQjhnAKktRhHzv6lO9FTaVm7QX9Z
gnZ/gFFlvu5PLv3YcDRlFOp6oK3kWqaQhUpr9LwrsgWB+/TJ0Hf/1Z5ZbbRydjTa
JmxZ0LScdzjqW+h+HaMs92F+WmEe7Rchw3YV/IrMgQJxdBB1j0scGGZxgcAtdqZQ
CnlvBPuWTJRipckuyz3fpCrJDa8EZ3IzlzoR/dCIhyFz2HTddZPkVrHsu8VWyQk+
BEDyOtro6LBU/Q9cirqQwbqOaV1mQp6fWCv3VPEywWGhd0u768S9IniSNE6jvyYg
gpZQHtDUQUNIPYdiuQFwLiW19TMtgNI4XxJNrNxBV0of5PsnMwx9ULktjpScQM5A
a5Xk7YTTqJzuYSpUUlVlLrkof2X7zaTEd/7Nre1L6Vc6Kz5RxpuNFoH/gihBZl1J
1LB1WRt3cpl6fNGG7YqAd7HjpwT8X06ZPt/2Z4m6cDOnEcaMn+pojBBHz6/0rwcm
kAaFvuP4tEdM2GD6AKtX6kUouRhInNto0JTGwd9npjtl4M/TtApO1oqPXI1OOp+9
hJwk+IFgpdSjyjiwhTJE1sWGmDgD0qm3NLHdG6Wg8NGDedpKhZbiX72NAczD/VC3
wX8z2W/NuBvRiPOv1KUYS6uivlkc9gx8ZB9KQrtdNXcT41vxjqLS/X3zPsyhMaX6
KZDE/jFdcG3BjLFuF92otZyaxhNmlRYozH+u0j+gIGPE99ds6jSlSfW+b2+gHbr/
mVta2DQNSb+cChG7R8xeJjkQots0e74CVLs6yJVojagFqFRF/pcgEo/qx/3oPmHN
gR2zEEKgbT5zaFmi9BQMciYCnc5E5HdeybO2FtLJ1NYKh03ASODK1qfIIJw9rDF2
WDXluQ3r7USIPc9Z8GZu2xGe/fdwXj+so8xE0iS9vaVpXDSpXPcNzpsIHkd2ZFl4
2A4/2njWlN2WKgV35dWZtZK6WLI4TRU+BbfWdog61ak0ScvAJDh5Jd6PFqQ7JHR3
poqQI0XTRb2DC/oC2J7M7XO6KXlQaaXfIUqm24cplTqLM4TBzw3hg20oHkfqqitR
MjQXukTs7+Zy2PJLqoTPrSuCaGnYADHb5UeaCgqqTU+1omOvJH/YbrnmdC8+IsLY
Kg9cqPQINFR+NZj72z1cRkbRptajFE2KNaJf1CtimXfSiYanOR+GzTpCsoH8frLA
0GdNWrq/oPfBq6FBLzh0ru0RupcXv6LC1ugHgmeV+JpvcfoXg05nx7G7eeTfIbCY
p0bexzfAcGJycIKaIal48vy6dY7NnCxcktv9Xj6aJkZpYJK5uR5dD0fzYLs9p1x0
8WF4DfD8U/NP5bsi9vMHx38CNmccwx78sdhykNKVxxE/2yOFQhEiC/iJYC3Ut2KG
NaBnCC/Q0Qh/zlSCl8PNOuoLCn6ZjPQYd5V+0iFA7rmvbaH2S5SzoaW2c+NofiCq
/gmQETY1KUzHLLvRF/UFnRNvlQ/xHyd5UfbfxxUfS2A79XhhOQA3CJZ+FZ3oX27V
cyfctDyeb2ttggcP9+yLcGAn0VIgXSOAjvzbqenH2Mhwzf16M2MkWARi0bYIS2Uw
LyN714F5ldfqTlNiMY9ukx0zfvyv5KcM8utVbX7tcQ2pXn066aRuQ6AWfZTFndL7
0el4dWgN40u+7vyj3y7gIUIjVPoRMySXfrV8XYtcVKfmZhsa8cdgPMWOTd5xLVd/
KqG8W4Scfuj+uis+Qh4u+7LEgKNeiPGg4ffxLAD//XBWN+4fBPvqZgJB4rs74GZR
OLdNeBOttMX5sKrjhrf2asK4y/XlcIfT1ANSqk6/t9T1MjnnRaST6fNvIe8sX+Vs
NtOp2+reit/TXoDV8+9fYI9nHWD7OdmxsUyte9X94eWFACYeBTQxXTy8Wl54NcFO
UND8KpPsaFYqz4gMDMIUg5fMV4AlVY9u1kk4SGVb95kUlZZrqqFcESNXDVfi88Nr
Qd66BBM8g4n4LqCXIqy4iiHdbfhzBwnrTSeYnzMzell1YkDo7K9G6dPmtJIuf2Sb
m65tZzNK917KWqx3tOFW3PojsBzj8BU7eZc3kGvxVb/ELECxWPR+LTByF/WHnS0f
UIRj++5+7I3P6XNVKn2iMaSIumYcxhx9rtj4NgTHHLdnEosI/yssXm2gpKawLL9k
RvqaPoCqgIGtkXrGo9SmuX+XgGIHsu6BncLVnnC8B50bRJ1I0l46RmaqBmiNZA2P
bxCnx6QaquAUtg1qMz6KqQoY4r8XxjqgB6xizwNT4uYRCYhfv5tbmuD728qXdPba
2YP0rbvhdFWJr80URRDQTs7PmZKnq20I7shXxKhQY8THgNiRhKNhjADZ5zBAz7HJ
+h7+re0kq4GOjcxiPoZ8D5BVI3Vz8vKlU0mdrDZH8Ecf48sbgYAtWYW6aqa6nXmB
Lr3iO0dUmdtZI2huBCxpnVG83BvQbeBwj53PaDZqX97NloQZ4ARCJq+kQGvPrX0Y
tlWwD9GmnGm29ad7se5REldIiK9i2yOwq/rJiaqO5M5mcAdEA+ql3h6YTr/fOuoO
Wo/x2LysA3pdpBDc9SW+f7hZD/fhTcSFr3z73jHKwrnMn3PzfWK74BOfQLG8B4kG
dYvrCfJvgTMlT4N175SOSrp+LpFWHjRl4ec77JmeEBkDd+7GUiM5bqxDJJz5XKiK
oIHWU+VscwtfOqA2hoXtPaOQpMia5/3XsCE1TI/Qg4iLSOqSdV52g2/syqU+Azk7
2FXUsQ43SRq7Trk5kGsKm4DKbMIe2D0d3wd5jiiaRZyd+hIw3dvZdREpZ56tyiJb
M6HYY4lu807LRz9yk8QpjfL03IoRhCBlYUGfsdW5/Xf2Bi9KeSRLYeICNx8MogpP
JDICwZCg4u/JOIGHDUQw7Ks3bGZS+KqO85spuT3h57/g87FTeHFZjDwOInM4ZFKM
zxv5YWnzqrpBRRKKSNLn8FQ3eqdYOLsRaa+0nNeoRZYoLPuYuS9HYGFV43b75X9b
Tr2DS8HRp6c444C9h2eDkVNDfUSllu8Ri5QRKyoXnOXNBYdTX+guL4YDZuFSHKjr
jMP8Afx+LuaWfAYESRl8uF9mGR/ZgkWZZ2eGhJJnwFQH6++USLwtUf2Hhg71Gt+n
hQlqZldrMDcdZJi/bfJTP/xhY3dHuR8PyXdo6MouHyIia6Ds7MD5e/G7hMAjXFmU
9KGzrQO6lV5/1VanAiFpFqTAHF7YbDdCdSe2KRhLkqciNTzLHLFo4rf7PV54lR0o
ma+hI++AW7w9Vme0QO36iECZp5WSfqkoW/9LmlU/yfdHh08nQgqo5U8DsgMZBbzq
pIWA4I3h9a6TraES6pg/1+Z9318O50OQ+sWsqSn+wFB1yKK6TPULKCXwDZBU9ymZ
uDmoUEEKsk9zRQi8lP4iIJecAB9zjB3qbRIOV7HUINLksEBg+UHTMu4/xOVqOb6e
kSVQ6kwHs1aei1EAVaWy/TzQ+cJHx+BZpMbpyoO8vKzjmCCYoL628rMure+YhdBR
P2ZW92HJWYgePiKNcxoV07n9BXzbf4coR+DBowWV+EQHHzdu3XiImRf5l3PLt1i2
cFMSSaQm4DQTFomh3uGH/S6QhHs1YWaaMdtT1qCXRGWJiG7c60H7aKukJLgopc7Z
3MLfmZzVu41mlDe8mXmozARYbcCt8bKTAnBLsXMtYtRSLmyx2Lnawdq3JUaxAheK
sABVrhZSfJgBq9EAtXTA0hifl0aVlNui3Ojaa70vZwn9jIcpvFBCdNGHndEJTqU8
JwSzsuTBkUE3ivqx8gAqQmWbLhM9AIDiIJBF5AjXGkTvhi6hGPbGD0mM+DnkCu0G
CKjp/glBJGu59QjLy9mU54YfNqwSyXs0bBuWd/mIUQ1lV4k4FEKJiOpKOomjIdEz
Ip7B77IK5ZsRZWUXBeMZRrvF6Sn1tLDeI0H4ahDdhMQpdAr6IxKGrytbYNFOacsC
jLH56fTXNWYrAYQkQO5LTMoJZf9dPQjvqLRKpNnigYQLyBKImkGrg43NA2mR7BQJ
vA9olU4B3gY31Y6B3XZBpH1Es7/3XQhmCavM5TbJS5/MQKEOkkD0pXHwltglnpPq
owVQ6WTxoFnQQL1Oc4hGqohcEQs1unv+w2jPYL9fPog0yloGk1wn7NoUi5l64lqf
xY5x9pD1svyz/A4CrVnpDzm9gPy2HA4hZLe1RBMXtTNg8peCWcEhKsLiAmwOlL/K
VV8qWzNCVXYzwmiNvrjLwYAkG9jIXSfnYVL3stYyLwxUmANIu1O7FDfHqzA754+B
9YS2gtyw72yNe3UULQAm+zHMLrjgwiardj340lLWElwp4ez81mSZxNxdM55tNVYl
B7l9hMA47J1EvFsFPlpb0tprtZUcGpO6z+tGQCFOtw8ZCqjJYp6p4zoHqn2pnJUM
jcfigPdMRQPP/fbHdDuIS67cJok9tT/TXeg/NkgWJ2j4V0bTgDC24gcUJT3pZ/6h
FgJCEt0Qnw5lG4CKBrybHpRjSxXK1BcR7UT1B6/ZZCvto4ezXEYanxAyFMAv91Yh
/u+xR39L8f4nhxnpely5joLmsiwDgYP+CItiaXrxEdt1+LilcDLyEsfDKYQjGAJi
7unHoB4QrbRe7ADMyOgJkdCsOakKBQMaNuR5VFYo3qr0U8c9l0xdsWK/C6ERk/ND
AxkYOqrrcy/OfWYvA4T+XEMaMPk3mNMHgN3CRPILSVBEiDYuD/yMo/cpAdkqaUmG
9D+o2TKkSXMNQ81eyQpdGQlTNtRQYRidJEFYe4WO6bwViZuZwt5tHCg8Wi7XJAbR
swIwXtpLBdzNw26AZHwwUiCcrvmOEd9QDQCbFJShuRviUXwnWg+MnyvAm301ZLuL
dF9N7lHjU2C7Y6hMy+9MWrxfuTP1w7rmjOZ7k6FM2/nmpon/jS5UXR84H8ASSqn8
cHA8g/nosQ33a1j77lU6PKCqhrciyB1wsT6R1AwMGeIO85H7xT0Xrvl0Xx1TtNS8
6s14JdHsMbuB3YbNXj6pFvTo2l4/2WGW+eA99mTzC8ppAgAcY0H9DmXbTE0av/Hb
PXGtIgQMeQMlMMjJq1BMkDgHyVQ28hFtRyOXAb7Eib9GpcfsSM26QSPRyVqclXsf
P9qhv83VTVvRb+GYUD5CfKmD9BdUFKntIIzhZqfkHlobPLxAum6t2VARzjiwW+HS
XGC3SGxLcnD+Y+40Ti0wlamlvoxXb8jAc9Rn3YEEST5ah1Xwwx9Xk2LUiKWvGwkX
Rn/EDbMiUZLluWUno2O/o7RxPoQ66RaJ99nqJ126o6tpkiM/icxGT0jwkpOUKPF5
8bz0rLRSIwHKvJOtvEzQiCasnPDGrS4fT3S3kw8u1BZRIGPZelIf8vvMTSJh4jZa
u7EvYxkl1c9bwN609deVa9MRhujiE6NwTPTl7UdnJdbvCuoUO9tjQs9FeLgO/xYL
is7XOOltzyzAE9IDpVJu3ExhAbTgynHAy9BUgVByeae5H8qiuF6cBbepd/qklV2v
RqRz90hXtm/bVmpH86IkY+ytjSS97biLPBpjY1wWKlDhyN/2VEoKcqmaaMm7hVB3
WhIGd5yTlXqLURlfP/96npi5NLFXV9CuicIuzxHhkwqOexeRb1AgGo8krOwKZjTM
bCIFsVGa32cmFOS7VwDz2DHHcrW9mt57+uoTT/+ww/gOLRduZSVq/HlIS+GOvQ8w
ukEv86bsjhu9tZc/XriRd+TNCJ7Q9BbH24BNo2OfbvY/WRXJYHjl1/KlcO6MktrO
XQIy5+167TrR2RO55K1Twbbqza4mfjtPjkopOw7odUGegk+KOn/rHiH5kXT9Una9
TGh+NJSgzBdyLAQ750RYwrzhB2aL4CPkOA6aAj3SE+xwj8+nxOBc9P22oRLiwJxl
p3HKRx5Rtm/DtzY5Rdj4aYmGNtEUKsO2nHfFcGtLa1wWfOYzR+wytdhWbccVmxad
oHgfKf0IffVp4Q87uxRUivgeWORLnq23lCcC2eKfK12QuKleZqDBWW8T8FqYlQ/y
9ew0M3QdzrcnCqX081v0pDAkt8JQ3xK/zvFPJ8KMvozPt5lyC2wW++V1qlGZfSFi
4bic6xDeDkIcAUFnOOXR6HjOiB/RaJ7C2EkglrjZJkHAGA7+fq7+poM4bw5kH0Al
RzyjRaw6rVSr14OI6uDYZmIowwC4x3qUhdAI/nfF0oLubu17wGZOogx23Y44NqVM
/uIcR7Dg+CgLn7O8jvzHHNxbllBP8HMPneMTVxuwibAklcaoI+9rS8RO62/ewgnn
kAvi1G35BH+CvyZr+t5oDH8/1QRySevByN6I+UnlQED5GDcxm7eecktQjX7pwLOX
W2WzhrdhRUaxvx1WYOL96l2vTNfsHLv34zM+cjO9fLB/eUP0kUtZcJV/CLKZadeq
kjzdE32fix46wJAehBGNVeYpYEd/uHohuHDaT3F1yW0YFMNlG3sKNTKvVDBMGLRC
YMVcETopJYWR63sA3FygWayKa2TkeuxsUf/Na+2LRmhqY/1RsTEXaVzwEnozKXAa
JZpgBwCZA4BOF0JCKC9mIcerIprRo0ZIuD0XiUcdf8BMietTymT84W04iAkHrT8e
L+gghWLdHepY0Zcb/EDMNjgTCX+NnBGaAhlAvR7viylw26xXVzLxO+HXkPX2Kmod
Xsd42QgT61M+s5swUKqAz1vBEEoPmik5T5zJLYx1lZXFmVHGHh3EQ5pimI/9EdZG
mR5g6XXr5nIAvjI1DkRXaPfyLtGgLnXcG/QOtic/It8VNYQ03mE5r5ntIOVPrdEt
S0bpr0qNY27qTwyUoEUtBVcjy7Ctfs6mUESHEmm/fpYRp4873dxLgX8dGi1+6Umb
tz9wp1V6T8IHYYdKklEa40c2xQ0LbTb7wx+/EtR7jQOq/DTGpQhQHnS07QyeR9ai
J5hkr9kRpoPsWjp47lAquDsqflYOGXj7ZDfPo1gYdKcTLQG5yboBDn99CT2Y0bou
93l3mlil8mxoTNeb0GVnAL29CQfHl8IxQ3g+an4kd29VegTq/jBb6o3+J217/xi6
ZzEMMO6BDUdtFJ7wiU4KLGAaclR+LswZXtTVWdNv7CWjkHO1qHxbCadx9RHX17ar
dt10GP+QdvYR/nbd09O2lnTV0HsimjBsvCDrxiOZ9bDz4RmMmnceeEVC5ZD4t8Nb
6QOW/0vkNkZhUyPXsoELHgXulCtcSFNO31Iv9Hf7bCYNGSuTVY2i1gqNwxfYKSmb
ILuz5uW51woDfV/2RPHG/eO09ieRfs6bT/NcjV7Hq6aJ5Nez4rhwXtRzmz0rsuIJ
ybSFoZ9ct6cBk/9dxXS5JHKgg4qo4GI0eEfqkRW+MOYtQSnwJEg7BntZTARmYR5k
efXf/2I6puyM2UYaci4ENPToGw+RQq9DE7gLHrJsG26p1OtP5kAT1IHMeW+px3a3
Y5EuRXb9ORascgFj6uM4ws+sm/rQW+/+t26k3QkTGTI6HzsR73pQclrCrVb7eKHv
LWBVhAvbQNRdk3NzKR8WOBSdRBRXiwzGnk/h3tvm1oC3LNftY2fQ5ieTnd1RQV5s
bYrWgn2bpL+A3+5n4t4lyFgjVswBooX8DFRS4dwr0Z77BcjZyrdjHK0nhXsDSkdS
3OAmUi03nOlpj2/4RtdnVsFXr38a7nPPlkJBR266/wJDxpuvlnb6z4KxQr2gC816
e8Awr4dXDYVMC1y3a6mJLhIquwh0W/KZ52Om6QkaCXww/A1EbpuT3EHfxdHM5chp
A68URsRKecF+xFqig8HqFgEJhPIidt1Ah2tTUmcHdp9qLIqU+xxEcqfzPDnrqXW7
wn9+xetG//W6ycKqw4EY/N12bsx44TzUeMuiPwF+q3tmuA/QRenpH/er+uEgTUBv
DXBtYo63wjqZGHB8SIQ2111oJfRoRywuyQEmHvNiD4QnTLCbHYQek8lw+FXItZ5p
KE7vvbYytjJz+EEvFWYdmu2raKemBRmij6fF1V4Nds9Pet+QfRdN21kHyU5g+nYT
HrkeD6nZbe6qq+BssVSEFhxyKIEqxcsXP03aKyDDG/szJyilwjHBBtKS3NXlIPcF
7qmvfZld73EwPfttqO6WFwathOrizgqemAvTFUPlmdu0oK4MJqW81J8+6oqG56wo
4buiXfvk5VRB2ZPCLTYGTqI3VE8z5Nh2ouwChEBdOkiin3rRGowKkEwlOu0oohxT
G+7Sp8KW0QS0p25/dOkusIKfA8QO5AfZciaGGy4+MsGMYMWB7Z/KbXZUYlYzBZGk
Ib8dgoYRYzajdn1NY9T2vFH1YBhiP5L3pidEtj2xyP8drbfwIQV+8gyOVn7iJWMH
Mak1Mz8Gr2fVGfEkFnKr38zEEgX6Ulh/5lNe09pwsYArTU3gleGoT43wYgYIg0nB
OQpR6hM0Z4y1rKZHtakEfFkCyOdk9gjoAoO3AxKqBFXEZYm85Z4xDx0Jw8ncEhnc
mWCVfsHF0oiIASnNGOkt5LVOW1MrE77nip9glKReKvA+epiAfRDfz1MB3Fn7pm9j
3vA4cnUXBBctTlHcTzSqb4odLFKf890YVAQnaDF/6zkmiKkjPfp+kOvHCCEcB2Ff
EdPlI9FjygAk5JZBMrKV8Yi9VX7IJgPf0w4BaUqEA/05ZJas2Q5ua9MnpVBpOb+w
X7ww2tSdjl+DLfYCZ81K8gVWvrspgYTKUSVsqb3ZFqdvEpX4pQuiU4Rc2Sfo+rco
pIScgwVhctQSy0TaIfAIBNjTPp2XhPlZmHI7B4uDkYt71qWzaSdBwSebqmuf/wuW
zrpAErH1AWcdA5LPB+xJvdHpAD/Gr9hFkMpaoZ9XXIcuS3+iQONV4Vxu7s/5N8g9
jRDx2F7kssU61X+JO/uQFxE+7j31bzvPAMkoD8naYXsRueNnAFg3iQ38pzr1wOhY
QsgNCz833YjlSbJPJicgpEnSTty0gsJKuAJ3htb/7zWuhSyiL/PqcdMC3QKRCaVS
cHqYq4rbe6lsxyjKWdh8+wDfIele204jl7gRDDlcp5jFZd9hEV7/227JA7kzvJQM
ApOGXkQ7RQdYb4e/fCLN6uTCWP/RZh+hCSaASzUT+DGk5sU/doeLxomwulj+XM03
/AkPDHcyAG3Zwcg20RFuFmOKEKTEALLahKm315mra41sPd02OTxLIpxO7QNpX2I9
WV7vbRxwMWe3h3nQ8WfsFo5ryBm/dsdxnaKUx38+cJ7/My3mdb5cy0e8KdgrKMuZ
AnBxKFayJbPU11EKmZkoKk7h58gwe/dSNSiyNyTLIv0T0IJh9iBB5g1k3xfYnb8t
fZDa0zKcWjE1FqAa5jfnnBvJFSD57gOMFDACxMmHxE15nE1HqhAPDiUA9tiBWWY0
NLwIVr1IgcK/b671kXkP9lHMwZsC1W0Rqtz6mHXU70EI3rBQp42ZdJbqTLH+Oii/
WPLNuHs5oV553/zRvztYfUiWEObGoB3NbIiMkRY9/cF0OCRGDnsX9M1CtRYxc1eX
jGJykZqYCB2jL4LjHcUP62imyC67YNVDJ0ZrAFL8WNE2RlJjj0o5c2J8e+pS542I
voFEFyO46ixoi0g/MOc7GnQGTpWAfudrDfxwTPWtu7F3LqsNB/EbNzllKVafn2LO
+OpOg0kQAa784jm257To4iEQVIPIR1Rxs8rSGErKhC3xUnrPZ0pki0CmQMX00A3y
FM/VFNdxsD8V3ekQDPyfe4Sl8SpqX4WQwpAZm32XzFKfYMf1+LzfO92nRtv0qz8m
cbdZaSPHA99w0DeMoWZgmuH/ZxcbTXPtzrKnjCNwfHli7fP1jFWzjHOif18/T+gW
56b5O2fK1VC0AVz7seL5eSDpbneaEUWIQes2MQa+WBDHaCfJ5Hi/pHzdTNm9BEAz
XiroO/oNMqYG8mjTZ1jcaOrUMu/X3rTgOV4EKVwqCYdvV5Bu4CYvKVzNQfTDBmyk
wsh4dstFiNjFETRNeARdxm7wJKwp0zeD8Zkk2uwe6xrl9m5aUwBVAOa14DUaBfVW
M5x56y7sUx+PTKMcj9a9s1iCWH89oEUclpdQKy8tHvfkQuGH7a01SwjEauM6T8tW
joGctlHkNxqBYy+gDQdNI74UbOXaeym1/JhKCu64kaMvwB1dHgdhbG5gVjr1GPSv
5QUiCtmSQirOOUD0lUB+Wu0v1AzsJflYN/gzb5c68toTsLbCS8Z+KEaW5UezqXm6
po8QEThjCDqjNkRSHjBiTKf9Ctgt1BOf0ovL1ll7Z29WE71SixSb2nkd+IBLUyU7
o8Px34X5UgBCsoUMhLCRQ4PSERkCtutOZHiOHKqUIbPhHi6Mx2h4dQVX5hnal5xl
BeDoeakW3c+EqOU/nm+46vt7YKor9CzXdbQkAKyvf2yqqCdqIZYxmadr/KxJy2e8
n+SofETLT+4Y4KCqbrVJS87LJf2ubt199oO7aSlbVQ+mFbY1QdmVFFY5tTfzpw13
Yg/LC1fa/hU+9r34cyJICwPugAUaAIQolNh4tvxpWWHwNZdAfgaAk3zovNbugWVs
WUPCUFNLJPdNynvuid/8+GR8HSCGuuz6StAT9gYQNyF3/1NiECQxXqtjJ4A8WPtl
hgX7mLzs1Lz82f/oMftLHGds8HLAXCVCytGVjmzmQdjRG7qIzRVbPzYghovKAvig
mWmwFcGdw2OhGXEo6oQlkg2qAyjfDczyAomPmSr+xmjbw4xVinpjoKuYibgx04ym
9cq2Q6w2mxfbKFaZK4aI3eL/0qNlBBlNevtSgqcctlIo98I3Avs7+yCc9hfKh9Dt
NGQ3s4v5h0cmKY3pluB3rIFwObM9Z+Uf/zJfI5LKmX6CPm8dBIQeKVLbDKXgz/IZ
RYLUEktQj0LiBaVt8TCR6RGO8kgnIm5+W+2WXpZW11dHYj4Q2mgkjg7vM/zL5u8E
/an2HosMQFOiO2zPZuUWNY3zHC37Y99IjFnIQF6l+DsdXG4PNc9mOmqDEEerRIaP
B+CYtQxUYQI6bA8Usi82ZYKxPDk1MlLuabQeHE4sU+Zf6AYdlLjuOIo27DQq6L3m
Jz/VOkEFr6yTWX8izu7XoZeECCmbjBGwCTLH/2+fWpOjYJECDgrTzIXwoVJx/TTi
Z+HQcEZ4icQLirRkUP7dN9ormPHD9FjZ3ZaR6QQI+XibwJhoVzyhYMC+2/PPnnoF
jPy/CL5xYlB12wLAenWNiga9qU8vmjbU8TWL894+q1PgS8JyzIsjWwJl6c6uA4AN
OIHoTS3WJszg0kVjtQus1cn1tSY5XnNc4pUX1YN2dPQdi/xTzUc6SnDdLCJhxfwE
DriYBN/YxlbWafr96jgnKJCYR5SIpxE+p1PJxQmtlf0cx6L6LpANu1yRRxwPeTjU
WRiG4TlgmWBxFfRjnICqkJuBB88uj6wXUZTOvtYBN9RoAhCn/edhuGU1KsSnCz/O
+sHQc60tMosoxJrNSBrjs+Y/Bu7pcTz35+IJDx6TkKQlOcVSMqqaTxQm9NGBRtOu
k2XStLshob2qI/EO5D+XdNLAXgN8LjH579Z2x7/6PycvverfZWdTnOWKLMMt0jVX
cT8tGrpIFf/O5litwokyILZSGxzcNgiyXbCQTT0056vTxd1YZZwIllgmFW75htkG
ATXRNdClDpWElYMSDhIRrFQXLDc63MvOSZH1jxhwGPKkjC9VU8jP9Cdxi/x3zHAI
9Vo1T1BzmuQyRs9etYU7IVSOoCGHx/yq9iX6ARo32X955KljyMk6jZPDhoFKRcTX
YkXXkOJ53gzjgbVmUjh1oIbnU5sddDkMifpzSWndc3joawm17Z+ofGyDvNlMMKmE
6P1WvycXF3sHe00P84d94QrcekTDIaYMgUSS2LpDdXUEODbCo30VadLYP/5LRmeY
5Naf8CFFdbF/oW9MOWbvMXNXEhzdzRP/Ve8O3upeqgPz+2ZXOFCwEj8azN5jwqnV
Eq4mwGADimT4MkDsDM3cmGhE8hrLXcDcqntwhWSYq1H5piHpq6m1gwIeXsqCMNQY
eRmmV0UjSdFX8oLfXyr5WxL78rymXoLkEBZ2Hw+hDQ+gouAfBl1HMXvlKkvg5idd
trI0V/4Q22aROq3XCdyvRn95nQIdARQdKUhmVv6R6iQCsRj7MryN7G2apD2FomGX
nLUM5GEvg/NX+QPSJeUNqTHqDXHqfWcH/99gmOcqU3hicR5B8TUhJ+LtgAAdIec6
7QrTRX6/2UjLr0Hfa4mYWfyDK47O9aLalkn0H9aXUcuAWbm5FGL6wTa1RZQW/o+T
whCkuLUdm4/57RV3rmectXtDDgB8JiD/FUrnvoFi4MMDo1a5uAyEm9TzL6WpJKOw
EYozZn1leR8ethIXEWCp5aEH07FL1MhNeYEhogqONrvl8Y1IGP80yaaXOGasRsB+
thUGi/K1UeYFLqg+swZQgmY0mXyGJVlg1m27UbCzY8meWpQ8PqdK1ng4v9jYcZx2
ocGKxPVAaFGF/uewyJmIMUwuqz367osBsmM6RhpOrgk6BOTn1l/xftpUVjEcAwOP
o5aqB/gAPnQhcrP/WuNMlc1MWftgS0a5AZ3sZA5DM4rgjFfKDmiXB8WIM1R8JGrj
iEPJaoCJxTbpI7/2bKYz+Qf2SQMPDDnFwogZKOdEXaea1RZ4Z9dxrcptJXcDcT7I
CJvbaJO3JuGzwW+X3ZVqoyeulbSrwQSRFVq0/6BmoGFjkP6hXlZzJAU/16c5pldF
LIH+iJDgfJm6R0zfa9zXy+pbiCGqJGGsN3W7cUjaiz/Z4Gr4bv6ssLsupLvebqjZ
p1HeXe9nPyR7L5RX0V9khuCSLLwyWt5+8+UmLlEqkgePVV4nqvUD5dtprdnmiv7I
waTwLdzkvHZB+lqlsa8QskUC8noObTTr95VTL1mpZcOHtPfvyJRI8mvwq2Qq6VOW
rFVnjEEyQZvsmtmpFSo+Qb6JpJ/INX9XReq59IpKCOwm3rdu0JvHuj5RNrFVSI+5
xw49pcDxkmSVi01n3gMXj12IJuWbaXhgBUltdm2WAaSyUqKmqU3woFK14Cf08INy
biu6CQWN4HD4wIDbPEMgIKOaUAkCwAt+zjmXWVEBlak122uHKmLL2/Qw/y4gG0CJ
gukNufsmJfsqtvHGMCLiqepqzjNzfvoZ/3YlAScIL65p2/gKqf2nkHcVvCsJVZTs
pwMZPwo74qpCZmehUbK+Cz9oi21Gz4zMlMpB7DAhXhaU/SKDUA/bC0XkiddNLYTl
IqVaDJsx6H4XQkLSBUP8D30ZVi9vHsMoE58NJf7GRxFFxosami7aGamEQwiVwEeg
eAIuH+HYQ8t41chaVR/b0jWp3/Tg27EO5dAL1e0v8vMoRhYi5MfZEY+PrzlAr51K
0ZT7Vx/TgvnoI50qrVAzGIEjK5nqcWRgLOfMAqUzTOpGS5QSz/sOLH2Faw79Sizy
dRrnx0Jp1fuTU4x2c9RX8qZVlVRrLW1dhj5g0daMSGvqM0u7KLcoujnIeDdE8BLo
FZBjFZ8U5KT8mEZ8tdPs+WW8vU1rMWfhkN7IrC0iZTqG5vji286Tmm1RXBUZnG0H
tZ1t2CvByi4YCsBU2G6dvgvMdl4Jt729tsQOcfvOqLa1AhY4bac5ruuBA2W5GA8N
WrkDXEvHQYNeuTj7mKw4YN2PPGab4XGmHF3Npeh85k1mcz+4+/8nmW/svG992NBL
p1qGzK2EiR+c3Bt8CZrn9dCi23UjcW29iuNHXYqmtYns5ItlUdJmhhmQDv40tuhB
E6Dfr50HGLYw0RSyLBZ/bKz+bB5O+d2BL8TUfwuYf82QS03ZVq4reMf7Xz7ATtkd
855hNj6iOTzwWG03Hx+yI9QF45+azJmeSxOJ083146wq0sPOPyuV9Jsqdc29iOek
h8Hy1Dtl1FSk6Zq8nJq6yDcHogrTxmQuWoohnTHg2nJDvnAfLTV6rfTjk/3hEv4j
+9Mvy+bNpzVw2ncIo071xKpjVnQhgnJYdNqyNB4ZZXSIFOgeelARySa/9zDScy51
jQoXd80r1v9RIUzSHgD+DkfBL+8uj4vzW5WUGpNkQfXeI628zt+Ah0G+0o2dfAxw
YsHFGnWRYdAJKqoi89SRzI/V2858DJ2hKGSU4cmqrlYY4X0tyJ0OdbDupWKgRZnR
9KorPspkKtQUrAJwEOnWoCY4oTmXm7+qSIbQAvrm5Q5G0bjgiBqLU+ISgPxKC/fs
Xw2Txwp/L09uYC8JnvdnahkfF5fpPCD7g7QMxKELsGhLjZFJHXL3wHGF9gVRCUzW
EQ2zZNR7kscq5+ngpzOGG0s6O6ebnV7JhsRAAnCp7vQ1BCBmYG5LdaV5fDS7osEP
ZxBSGwnBjF3Z7pGKgBUnYg3jfA1qfxO1qcmOcG5xhvV+tltcICHGFH0FajhXEuAP
PAbUh9SeChWVXiu1ByOEcLGTlcO/OgSHHBvS8xiJarIAgZoUj8uNex3esP7cTjh6
RJGkdB9QfVJEpZ2d1wkJyg0KcfrodiB6yRRjKno6t48OUeAisI4ZkunX5sK9u+HJ
zcFQmDN+CF8nTuVWK0VTagKQEaZ/GceOWPiR748zY1wzGblxd0MkwPvAqFieisRJ
xO9/est+qwmaf4eKeini8A/uZgbyI2DDRGnevJYlU+RORWOULLGStUMku3nbvbiV
hz8xav6iLFljn1mgKpExRQW6BNKEXRFHhJdxf7AxeIYUsS87Vup/M5w5oNRYHQ3Z
XqhmsQzDhVS9wJkqSIjd8oOo1lC/UVyDNeylzIfH9MyHRA8RSuMx0fw9ujN05OVd
/fRE6MrgfTE5mv3sa7DUD9geTwZrjzQox089qrEaL+MLbbodMei+qNgwZiss7+Lm
sVRVRKnoclUjzh4bTMewsUVq+3EPYwocAlXvJueJysp6g3t4pgdmhWqv1+bWo7Aw
fEY92UJdDKcUZQzOuNJSLpcNOapxu2QuEOGIrkGe7/q2A4h8bMTaZxa4jfDXSTR/
p8dX0/buOMnbse1YRxsmJL328ykeJZQA0MePwSAI/KDGKr540NKCuTE9eaVC4/f3
ggiD0Cg5BHN9i3sk7wsuIeVz3lE0ke3DawuRtbzpo97TCMhu5ZQbuBZxdHS7IJ5L
YFMIm6h6FdnfEU6EXWjVdRr3t0ir80hJUYFarV8F1GDoxdKlfh1ycij38aiAoDmE
rj6yZ2CcdvrT1WMmaYA5Ca4Mfc+RW6PIvlwRUItRGmp7+iOyG2mazzOwWCAZMIr9
N3mH3mQRGVJ2gZvLy2nN+41mJ0bsyZPdIYp5hNio4O/Dw42fYbdshWQRyCA2z0U+
JuLhe2NSKPZSdrYX89KHDTwvviFPE/Eq2OWpFYYpyPWKCVSwzbe7400mbERK6dh2
SdDCVlFv/0kpzj+T46Wq690wATTClKoyfqe2ZUNOAOsGMar/ujRX4EwhrnqLN1FG
ztrVuVtx/1DibiH391Q8odoBpRmv0CPwi5feGK/+DJEMJobpYeJ7Z/0EziGDiPH/
0yGLGKeZmZADtDtIWcTd8oliJ1WwZZ8d3IALcigFNvEaS8JPMcMzp6NvyckHwisf
+1QRxpRupW4EAsT5cagjffLfBS1majkf6qwgtnM1/ePNlOgKaxYoSyt4+coGz7Ar
W4Fd6paEIc1iFAwpD3bmFKDY2HoxDpBmZ9nD7K7HA1hPoYdRixPZoozKlxY3+Wx5
RRWp1yV0kqygBKNQZzL8eiEqEaTZpt1xFOHsFNCgI3MtY5amOvbLc9JTQJQeqANI
gg2UScrpETa119QbnZ2OefBVkgrZh5OFT0tjzunUbdQ4knyUoHRrXYaYdgy24/i6
bOt0Q6/Mi359PODoMLEw2BqucS7Aa/MTxD15T+G3mMPXsntnndKmVU4i3lZeUbiv
YkMv5BRtmepaVvV7FZxEBIaha80cQ4e2HuUgu05YV1RPwJlez0F+tTEesKQ+hmnD
mhZnEEOpxKKlpW8KYtYr+969vA7S9rilwPlYNxkoJepghXSYp6HOKcRktbK5/dHK
ldKauQxbVVGuCcgx3B1e9OAUrxT9MNO1WytxAYOI9ucsBELlRKcRtRINw/4ZmBs5
VSwfEsmy15tjgt30ly6wK8ZJWp2ze3m++Lw6bEhffLL8ylj9ru5Ft+u4+uXkkAdY
0wsjIJmhoJ+Pa6EpfNR2gTByVztXUkyBFFkA9Mmpulxs8m7gY6anQ7BfRYhZNgwA
xa8enbqykzh3b6ojh/XYtKoTuluBGTHVenqoB2BUzg2TFRRRr5heqqaE/sMwYwEm
Lg3lHqmBSsKR2GTXcTDUwhowvTrYXXJeWgqLKELH5yaCoOA2SCUCHsYplka8uJ30
mankPAaJ4gubjPEGHdiEqfeKhMQAyTVot63+2DGbSmZwmFyF6C3Yuu5VPnzkHIvI
Z+p6CFEf6A0dw8Rf3WfJlEyOI7x+jmH44YWeKRgBoBUlmyI0Fbnk1+1AXhfXVmcf
6ADpbalsnCNobjOX85oHurOt7/Styn07dksmHQrOc/mwzPy7bKSUrhH5FR2WLncf
AopDQnV8e8MkZnTbUeG3r6uNsCQLgu05g7+Id2gPZUTdtGlzcaU5ZT/wGNT/iT2v
miQiz1XyD7NEZoIpeLRzD6XGjswPg+hRkTU+zPgX2mHq4+L+CtakayNRMKlLT4M4
1dRvx5gxClO7dnM+XU0s0e7+t+E7IMmxkI8I4N/lda+WzqDcVNFrute8Ebqcv+Ug
c33wxQOwAkklJKjUDH3gFTg7XTMSBFkc9RNI2fSwMobVko44Zg3cpOlENFNZsuzL
R7zpp4sxL+wOkIArR8VxYnZVmuWecKYuX8lHjk3/2RxLb4jsye1F7fcZzDyjGL+D
r3ERfmq0RAKSq2IMsJCB8QaDFX6sikyhjfbwGIAUt7MnTXVuL7TRQrazoPi1l2qY
Ex4I1Kd/SB0ZIKinYZ1XZAmBgpoySk5R/wKfmn1Sx8GcayfDj7VJDL5hJ/GgmtzU
QmClewGv48jBR8XXKGbTEiVTiZSzWHf3jpuMXxvjzd9xGb+zy7AT3swX9hBA5FeL
DCLeIJiJXfMcWX8DR6PeMFxcUekdrpaalvX3V7XKa8o1lb4kPaRydg5HoLB3Ppix
q+6tCJ1qp1UiMVFO6dhCp6ZNhgB6xZSKVuRgVODFDjb6OeScoeoinY3dZlbPcQcN
9HeeAQCfVBcio0ptgF7XKFp6zzK00Yyqch0/8gBlBiHVwLlVArgEITKN4tNOM9mR
f7u4VH1gQ6VRf/OqXzSWiQwN6kSL8LPWSOxp7AAHXIDdHWf8UZ1I3Ydac9S73lQf
Sr1OeLI5CmKeILSMKmV3q6GubK+aqQE0sP6BqsWlKdaA8XuiNGAxO0smz91/0ShO
/CYYMGA73WGVXnHJjyqB+UowlGtEmcPd+VHJsGjPBdgAPFzsls1NJhOgrRXkENDm
O5KyzMtO460oCzpMGFz3iJ9NCN/+H9hXpgCShHr0B+vSJXeRTiP0PpH3wBhym3Ve
z+xEEOuUuu/iejx9g04jU9nBHqwogRoimXhl+vr0eOwd2qSVaKWYiskOu9XjgdcG
bUSoCNIwg13/nHrCxRB2dKg/RdJAkU6ffzhRGlXZcVF1Yqrage8bzg1v3zUYbXzM
MMQ2dkWGWDwS1GvGRwM38vZblVtsqvu0dM6L8b3i/qdFyXMT+hbFUh/MxS4U60JW
MM8aFu56DTWnZjvUZ1QAEGEdGZnptTKovmko+Joh5ud1nZjYhJpLZkKIPX/DOZJ7
/KgtSmzy71vifEw3ayRiPq7OmmtPZoJtBc2xaWdXfTHiduWZ/Nr7aBiH1EeQUp9I
tDJ3zKrv6xMLapas+qkF4XkwwoP9atVXbKQ96ii3igSEU8wTYE4BEGHxrwlGyuHX
G5EIWre/TZ8nrGrJyr83Vv0gLSm/h7q/C/aW4no1hR+CNcJJOryPFGfs/wg2IMRm
Ep3JeEP/qYAd852uK1av/1d/lUOVy2Rmi9QB30zeLnofETsCimNWshz12JyVZKvP
1UnIyckSfTwDw46bfxM2N3p3lO7pzHQfUi8toyI7+U0Wq9T/zJR9XDwHoZHXzEGv
nFj2DZzzVFv1sGHf9/fXTqOmafTeDEPv1igu5l4ylT4OUL4RlIHvneWB9BZ+yVw6
udtdD7ZaEz62EnO83LXJ/0mplf1fLe7DTALjbZjgGvqX/PKTiH2oO/SmG0bLt8dM
q3L1ZUuY7o7HoIR43FWL245MXvDmhg6TVnbdu5vbUBByCovPdiAGDjaXzvMPisdc
ZhlxHfSkTpzFHlou3Lv78xgh+Xgdl+cnmr9ihSBMv3k87ikbHiaKQoNzH91bI0IP
OTN8WixYZ2OPEiQ0KtATFlWNL4CX+38rUuxsVmWekRppniX2FLjwxrJhAseA6e7T
dC5Z9w3sfZJOx4gtBaNFWExT8Y/7v4+ZK+sxGVWEFsrg8jx/revcz/bp7d0WINCJ
Ef6RcDYHpJpn3RVYEjL8Xjk9aMGA3KHoEr7Qo2kUNGwHeAHN8CuGdSrOWe8CAVb1
Y4xlo85D0iOI4QQdBL/FNKcrymaNQyztqQANxJuCKD3dITtLg+HtjL1YyTgZHFFl
5PWOC5+nR15vum1aL22slDznkngePbi94iV4okLUaC+wHsKr7bWhGKy5euGgKdkX
peng4/kUOvwhzq8VKFekV0hqgcAHcXtYjG/3mU7W3u2NrotSQGLmaPg5LntyT34T
NQpaRJOPSAU6PU6LglC7ICeBh/+M0d7m+wbykIv7ajrHl5hkEYb/B7EqVrl0+WA7
yseFkOTot26UPj/y4vZzIYBw81XN6V8uipOqKQ2QV9w2ah3P7iDSftv/Vm4Bg737
x6qpm0GSih43GLSGWPo3R/QpeGnMCfqPxzumh1nmBHojyC3QuIrdx6MzzXsDoGNY
6Vfot7oaMDuslUnMBpu2s9unT1uWZFzN7mzLQX7Bv11wPyhdUTBacJuk4zlenyqQ
3B6o4p2YR+VavW1i1kcOmutVOM9UEEMF+YWHqazKcZ/CLdaCjDxFcDdz3hEMZsP6
j4EDqhw7lm1Cio9GnIB5CuxcrynzuWPQGZKcmqyh2fnBEoLLTuPem0tswfOnTiBQ
vJhKW5ukv8FoylnF6X/bm9MrXE+oRNnEAyr1gxCMbnUfQf/YwzQ424Hk45IcP5yl
a+ml6GFtsg8vBxDlZj7GDP7WONIL9i0zB7FX5mKXvL5jMRjV20MCXXMRq8OFoNEy
u8zKwT2FTe9XAnb1Dtqa+M0hQqJsqhGQq9zcA5ewnOEy/r3bRqEJ3eSMLPp5QU+l
4/ULzVcpaDBqQ/jlfMzuZ5rdcYEaYO6XuQ1PHY5z81LSq8j4NEEcHMbezQDqPxZ+
qaFVMU3vG4Sji2W7PIBZ+XxA8k6Pn6OpWBtICeppIDETbIan/o62D9mhlF6KkJbf
q6hhaAG0HerIpE26t+mylOHgrsET3FVNiIylKn6DM3c3Df9u0Fa7OZUj6CXeHYVg
sZfRaiD2SNT4YzqpUrdaoFpjq1oU8LUpoRdQbKlp3EDpIDcq2SgvaiFA5q6lyITq
6R83iZuiRZy6rbJDRSH7yJpi0yi0WMhVElg9HcK3xUM3uQGcCSrg63wIZpZDLUDw
P0t5Weqg+qscxohtlC6xBsDj4k85RgDtRa/d5m5c6JKfW2J/X5+8fYsYqWK7Ag37
ddU3NGB3px3fvF0rh9JD9RXEoFFvOGdmLmtorxo0cg8q3i4t20dOtl4eNRc8HcwL
8xZbaPBmpGnNk9cpPHaYklRCfbOWhNXkxrMM+DzxTqKFNbqLOgTiXzsCzAY+DMew
t+4fA7seNkh2acM6/Hk1XgZSivfqK1dzussZVEpMYI8KtSCJ45GH6PIrME7euNVn
kqDMeuZ5Ef2bVqUq8VXk04bzLIwAHJtyRPor13YMWFj5UK33izKm2XtSLZFtTs+O
xdziyu+Oq0zpL/Ln47cPuyM46DUPe9oW1MdVarVtOh3cjhMEMsiH9ov0mtBmUQ3q
zH/ChnLPFpbFfNL78c9mr1QyjZfHTjWfPZlw4rHYVFuFe+iUG2WxtinltZrwGW5a
ebDZnbV7Q+yWNZ6PA45yQJAi5OUQJKv2D8WsRm8R7RAbMFy9irlt5FYnvxZa/W2Z
bkkiIUM9wPE/bVxjTAMOx6wvnjzMLBFJZraqzsa2/oh3hPMrlQEc6CbDP20NeMbV
2AhbwqHmOePyBh45pPYDQQCm8+rCzrT6/JkOv6bqGhFLwKbny9VvOzeBFsSDcvzh
jF2v3/9Dzae21esogEky3JmMVMqV7XZ370xbjs3Gb1EAMRr8/DczaHNNeqNb1pqd
mywXmzTMrFblhPBXwCFl4gZmemye3Y5FCXaUXCA9KFMdfp8Lto/aPV/YtgfTwVGH
netWX+47DD+tu5XWJdGzotGWz/6p5Y+0OGIJ6ViiBTe9BgmuLowWmfZBH86/ffIo
eHI66201HfK/I9Q53IsyNyyhU52+m7Q8Po3P7kjxsH0q2QEe28J9Yn5ggjBpkZ5Y
D1MQpL1EfzEfxueCfTYh6Kexeuwg/UcYzQF0TtOhzeCpxSBXI85IR+AaU5/+EYec
w0TgQuMZDzliDDaR1aqjusfvBzbYgbJIqh8CAEXEdP/7+QKmAyUuhMjUrGh8UL9E
HsSgIHjtOXd8YqJ5HtcsPLNZeRn771SwXmHiFJRU7vPRilp8gDgNlauV4cbIxF/4
PYjeX1H7QSHB8KAHKxEJwcIL6nkshsrOU/X5zafQgklYWp2derTCm1MAXqUFTW00
qPctMyd3qOhLOaJcyDbBOGx6QDcW0+xY7AZPyQYXwjQDWAXsPuYA6Q9BK9eVkfcM
dSzMYvivWcjkMVrl6aq4E9h/sPRa9Nm8IO3RgbDR0yXorE3g54snI/l1skgnqcxI
N7ack3/y5ywijCm+MfNogXoToeAe/MTEhckvufQqxv60e3cRom2scrQkt+bVBIi7
jnUl/URljY6l3wu9y6HTHMIl3FUhat9HuwVUHFU1J7P9HZb5/QZXdfjGQ6vZ07hp
hRiUy21B1eNYpneWGFp+aWjPI+UkPvJny0+5TDYGpvD1UlMB1cNRlNjNaTwAv6cB
V/LbpPtlXbQRr1/GYvtNiO7ZoBeQLX4XVU0ibICAIigRZBLwTRCu0J3A/KuTD5uM
fGBY2lmdoeg6mtUnB24CuDz8RaajJ/vw/QkhGy0JMVgfgUmCjrbJEEcitcGVLRLS
gvk98jJZQM/i2fiZ93foZLnaFA4BqBowasOelEdgmVBExJM5MMzkNwbSuDB+uDif
OLHlIh2oL43AiOkH6keAwobV3oxELqI79rdK4bCfLthauTnMgzg0pOhjVMHXoNac
kI+J63QWxPw5JMpOTZDo/S3JQhHCqEMjzxb50fU8oWhE+M4NWX5huPsx9ith9e5b
RI4AVgBaShU22gJWOmoySvABsnL/ow5gQ0cWNMAcpF1XORbU0RgvoH2eDIp/WObB
gjjsvcFCnq3/v0ZASGuw9aU3AFo0BsH9p4lS4MKeyqVSvNuphCe2aWAR+Fo4b+NT
NYXkPYKqUqTIBTXn+PJeW1Ie4CTeVRxRsrY+SsRvIvUk+WoKEJcY29PSUNCC/wxy
3rW6xJOlFfTXUq//9oB0dR0d8rSeY8wY0Bu8+Cs9Ecarq48GzPcwYYx9D3P9grsQ
KNtF94WIVML+nZWzjDDj8VGvjCbecctwZA7bB5Lh3qwdeGwn1U71CM/T7OVdIyyP
TEJpvRgfM2Gme4T0wQAirbEu7VWh4/DdGVgJ5SyPDPdgOHrCFSbu1V7feReGVOIB
m82hswrMOUBFq+LiHVbvHAgu6cwRI0WF3yikdFiWMzv30amFB+nty+M52CUisrcg
UNDf+2DxgX6KmfUHWTuhnVmb+oodBioHaz2HI/f8B/+LuEBHXFrTW9Wcz+lYX13T
ANnofHpjG/w6ZCEP6jJtof1VBOmdhTKleyLH22MWIzLjCQbI3IH1cALWDQmaBaKT
y7XQX4xM+chy1w48CrmCFoa4M+Ta4fMwhHEMSVcX9roFn1QgbUGULxFlil+wyojx
0xMPHxNlD2bmRY5KVBIorIGjJij4xsZNcHeFyeYZq8IdTnIK0C1Ehx5J0Rm71KBa
BiErNc1GlZ5iieWAhVDHBrFJrliaLafE+mRb1xJSPrpqWy1LbMG/TtdQOyzygRfD
KD4QeUvIZ5nv85nQsugcNGMYyeadeAVmf61vDB7G9k81pS+FLmESBU4BzDq712E/
B3+ecrt4hnlKrYx+SOMigpMbJYmx5s912h/8t2NVlgAySa/le8jvOglMmd5dUvOJ
c4645yq2/OKn4SlrLS9qlVdDbM/ZToMDoFgAEdfRoCGEEMUej3BkWAlmcycmfPhX
fdm14kvqkJcfzWy8GqE/hpxZ/HoK9EbNdrZ8sPOkq/SDdk43K5CRDE1yAMZZfyX4
C/Cutb5S2t+i4J+rHFI1pjRQdi8GkVusWvPDhGcJFqChSmtaRrQSvwZz93CyIkY0
hxgi1XaQIFTbTWrkWJYxwdm/S/rwn3zcQKhisZVf8GOPbT6H5Z+GoXPwYBquDHxp
a0auvFOdXtz1JASCNhXElMDPZon1adrDdE3M+OqqtgmqQPQYziRa5Z9fljs5fedu
noOFbUyFI8YfIrRkpra9dCoNKTjYskW1O1ZeE7BCIr9WPv7LWEpU9KJ3hTFiopVV
DkwzFBwpVh8pXSeYYLHtynkRyxsD5Ct7lS7viS4LM2lgy9lL7+TlttEOngjnMbii
O4TfOmt9RTycdOSbmT/vt6sJxNztZTJhF1RD4KRRaxKUqyQOkz5Bix9rlugYOi9Y
NZSz6Ets97d/mqqfU0LIpLhStrWPaRk/KEI0knXOE3T/sRq8wnu8XotEdNs6o6Sy
4ruFCaPjtiJsS/ChxyZYETnx4CXbZWemZz7ReG8qAXfQy3TRJvXCArY7HtAlKCv+
L8B178n/a27VhnSG+nYsrnb0MEd1I0B/v9ENQy2Q7t7KITvu59ztnqRPIXsExurv
OUIdC5gndyfOxguqYrsJeNP6yHwGwOhJHjmEPlXEopKeURxvxJJj3vlgOcm2+TQC
ek02N5uaTdjiyZBjto1EIRIIpioG7qMFN2ggzB+vGHSnH8/VcctsXMTEJkYQjh1P
S6C8cHI3xxOmu08BlkoESoKg8oaDntvkgqKPxtHIwUomlzi5XiEFEQS+V7hyIuTr
O/eo0q3knZce+x11pJn0YcoIz0omSnGzsf6ZpaWTRYD64rbo8A332f3zq8ZgFPeD
hDnZ8AkcZxLFA1xSRnt6AJ8oxuaovTWZWGD7I0KOWI/W6a52FjojvkkAq3kM9+q9
O6QGjeFG9GmasDQGP26FQP0/Lp/xoakHAjjxogEwYfkE/3aL2Tfmgc1F1e/Mn4WV
EFzd1FD45hZd9vQa9FV2GYnTnvxgy6bw3Z1sYPz4zxnzJ51TbM8GaueupFyUifzQ
y/+X2sROvwes31EMzYYkfWGZG4DH9l6b4ptVUCqkzH2T5ua+Gc9/6XM+nBCbSjLI
yT45dnuqdLGvsth/p7UEnZbYaQwqayPqxfN80kvvA7phsQmCf6RDCXDcX71wVcC9
DKNgzmLOjKB42RPLXp6naQtm+L5g7jmyfb2/CkJXE8yQrWHVa0957cWiFsYWniE0
sj0j0FVycHUN/uo4jREIICA2SYHy9cfjaTpaWOSoKkg4J7sIyH3LoETdm7A8moxe
UnlAzokbj8fWOgYTq64dA1ndYKZ21C3qr4bvO7cqiRfToRhdIhqqJLC10r209Lax
wz4yJIUOu4nVLWD5uPU2q5SL/D+6x6yLRm9jEAmqqfslK18t5GFuhZTjGRb6imBh
+qlgYLJ2fCZoC2DdDJAibOA7U97Gvs7la394462hHEuQm4ZS3VxTzDgIIQPxwZ9r
3fPvSsRIwlgY3Tf1R8NFMt4I1CCjK4b+zqu3R8UEtzxStjEc5hMdG4sVe89C3Naq
YPe67VTyRs5iWRiLrFGum8v2GBjQZTu4xcGwYN8HDtKbwPvQmafwwesHBmKKcDGd
0mImbdDJI/VIfh6JnmdWapSIBeUhwu5O8WGFGOL82ixMCZQ6u8xzVlZKP28W9YRA
KWGZDk5iiSwgVnqcgm9mNwxcjPF28QTocjkmPEdfJTvg0/ChmyPwRNJomtrumq56
Ky3rrPtgAdVM52FiDpeLEy1xrraeDdt1ap9Jeb0Ud4OVCNpZy6to1iyOnftQGaVK
eczZaMD9oNzsGoWZeUpWLgOK/fT8CpHwEZQkBYpRJjBjLS6264b5lkOnpiheP0TM
hg38UVzdxkSbs8aum/A3E7a/KHPOmkWnJHLXYI6RmoGztSXyaUuTQR3lBCxnj8QC
OQKLMmBATcE//2HMKwf7dbxxmAZ7ItiRcHWYYHxpIezDrV7pXmn8h+tXCl3gwD4l
kG4ZKMucNLQPtUsYLXO1s+1jOImHmiaJvNv1+/Ojidu8gWL7Ccrr0ydSy0VHVpx6
XFa+79Jjc90XIPlxN8n7HknrAp0SXJW/GU8pw6Qhh+FbNWJwRfiZf6w1N+njtRjW
IrQwLvOuswjeFWKFzJDoOp9UQ5pbqW8hx/KmhRk240Wey6uaAI9K5wPHXcOYXkIL
Nxec3UbK9DAZ3gnXJZFC3X0n6xAFwSUvycDPNZh6ZyNGsQbbwsaEOtbDAP0ROkEF
1f6I5YxhnOOVk060XiyWtHm6umx04EL9+RIhRFokdKtR6GJ5jxpHy9fZIaY1eU2K
XR+FJv5R7fWBrmPzePkeXoGBwxHBtsrJFHrg4kqIPCy9CKTjMpv7T+H/04x77e20
nrGWbQAgusNZanK781cTWfzEDyI1/f6avw+0mLwtwseOtWcx2tjoiWq/6E+1jFtc
BJ1xWDrabHNw6w43zbsXL3ENFYP9RFFbx7fHYsF7YkIUjYiIKbGkbkkF2B14wtYE
YW09j78THmIl+CsOiUpmuI7UYlJ0BovEYFh/oDolz0tUzpBkZcAgZU/yb8eSFoy6
d//LgN9FUAidQY7uv8x+9cogEfdIoKr8oT6EqiaGnGsxmVTw4Q2zae5DCWdYRBrv
Oe+IZG3jB+Vb7+A54G0cYj45KVf2Eg8tf9Lh47lyK9bfhAN+p3hOfWKhGvjGyz+V
QctanlwIAXO6SJ8Zb8co9eghBnWS8gqpKGvOTX/qCk3NgeVjijWQlzUdoZoE3qS0
geLqGTawUZ5xhi8btUya3oLMvCC/dcMUOdgfd5IDIumKfxufMhumPhrKYYKWNqS7
ulrLFsIjsLJ1RZNwlggOJca6M7nJ3s9iuI9miAnjxCw0kTiJfkmW6dp/f7E3bVpZ
ZGDO9y9ILDIFEjt2j/1q005VAZlv+NgQeCcglSP2Mb1LD9+fzkjwuxnQ2oE4niyu
zBBB0iFMRZkfraxhHGpe6k4FfSZbIwkB6ilfjGNaYGiL2ajIgft4ay5etZYfJnwD
zFcVBxmL8FrCxIFRxuqlgx6A2WzIS8jmdbsDP8xPNQ2oUbWx3iw3DqJt0C7mVZMr
UhZ0myA8c0Wmn2t66aOWRKjGlvVMCA/J3UNgR5IY3Fm1hd65AHLUgZhHz5r2cMx5
lUWdrUJzQkBdw+Rlv32JjKKFcH7iLzNmSvxUKibQ+vcO0bwHzNyWFGtGGb4yFn5X
Jo4r3gy4Gc58mzl3UqN3PipsEPdKJMURnFsRyT9Vfv277opk5MPpopSKLdSU7nv7
snh5J6ShDtXKFaovOtXyaeY85UJFwFwNf03XhB0gw9aO1AqiV33E4LmWg4KaPquc
1I6OBwg7zDQmtePvvzsgSMXhK1Rxj/OaZ4Pb8U+qT2wOXo3t03uV8OJxZCmXBEZG
xfFUwGgyLywg197ca2iJjyDl0CHRdI58NXFYlmWKbAVyaA+AQs/jQ5fxXEsACT7+
0T3hdLytLbXKUXrQPFFXOD/jH4OQh+nepm+WKUfOruy2u6fsHkS1Cg4BKJFSuQsX
9i1kmSEchh+dRq6dDtjUPOmXvhltYCGYxtg3UY9JXs+vuMRoxZ4/qu71MReqASxy
jVofxWIL2Q1GpN/hAhpTo+wmQ3HJhzyQSS8pP8qBWKnt6MbsL6V8m5eLFeUnU9kM
cx5MMAJUJ6Vk7O3UZZMfukvZiEB+mCqr5cX0Ci3w7R1JFNmd5CsDQCnZJAajaieS
RjZg2WP27zvWEDovq517YZ/PyusAwHHAb8fdc7M5MpQqdwuA4DS04wRdPZAUj6c9
prA2upHm9vpOLk3uWWuviqBY+LPY58U+T8x6XmM6U2njaKIRww/VMx6QJS/8rxdm
h6Z+KADCz2riXyiqYaZdn14w+MEQwftsrdLuPRGacab91gtKKsbYCUkYq1+4kdHC
bvb8yLjp2SAC2m9yTDWSTtsDkKgw0w4km7P2MD1ToATuIBQImM/AKpWQzx4hC9Dk
OhaSOmGFmxxkLkPXWKP5ceqR/5IVYpBp0Vpyi3cR2gKELRkoFzI3oR77yj5Ur42D
Xcjr7W3oqXNzrsIzuI2yAMRa+cT+hnr2SN+c2cTamInbxF50fIjidMVKDXJ5+oR+
mey/6wGubchyIj1+YwU8j1oH6WjyKhNMY6SzzY5mzdvSibdkI5KF7EGRQPpDoAXi
wF7/YhNnvFeP8LKk7NUbhYEBof+4dRCPcsJGNN/MgE2VaGeRpgXg/Uz+TvyDvlY/
b3L3eN8vqEp+6afe0kCE84WrFv8YPZn2l43/mIRR3DgtX8bxcKYAG5XlyImJDUSM
OFv1qD0VRfbMJCN7JkNfuK8T1+CqCZlaOAz/K9elHG565Z/K/Qgxi8hBp4R1NTZi
6AGGzPbDvscAEwzc4tXCXjCX+0lZdVbyZBRLZ6tjh2uBvWNIj5ZdrQnoLd4v309A
xcnAwBTAZ4xukvrIU2B8nTb40NX69P5Y7CbNST2KtmswHFBbJMrHRLGi7Xw0U42X
drC9rJFDVqXB9IqQaHVrIchxWTq9VCVkjIg+DK6rPU3ESpr3tyi1xrI5twb+FISw
1s/xipINMVx8UjG87k9acGrm79vZiXDtd12yCpfTcFq44RQH556fhaNTdheqUsXm
jLsl4T5RDSLE5JVQpIPTfiWCci9QwFX3BrZ0yqX/3CN3W6cJXoZHAYuTCXxuoPV5
k+eUziqczmGO0bOcppTR2/DgAgG74TsKzKiM/IkEkKvPYYWHeGmK/M0NP5MO8amr
9qpzDbOaouAdGV0GcxIQr9nNLAa1fgGwHEeZo6DW/sO7tHXy+KAeu0Z+WK5SFX2C
BITx9CIGqXscmuIhP4M4UWoJhXh3wNP5R9BoyF3ribU2KC+ZV2UwjXEghB3Dhzlq
WmQO3JghPOeaM7ZcXYGPVBn5eNxOuKWCiXnaF5am7VRioOjPTFnNEXVG0eokKYiX
x5jF8so2Q0OgJPSLOt4bxMhQ/lPyZp7YWN7/KLLfskBpEKdGTqjLcw1clsJXion1
bEXFV9BFM/yydc9gU7vdBAYiTHcuKrwyHnIhsKwt1ioFzmuAU3EsBrQ4SLauSs8W
SxrLq/Z1zkCETQWHWIird+1iRmb47Vel4xeNOMboEfzlpd9wWLfEh+aFIqrX8/VE
t6inNZGtEbPif0ZgB8MPXzHPyZORrFyijfcrZIt56E+5bc/e5NHbqfCvQw785ORl
aAkt5n8MinIyyQG/29dpleawQRsHPl0wARpHk+3LajT0+NMmxYbU1XD+YYMNumAm
2R1rqkHG/hestU+HCUrmTe0g5LfbK7Cjrhxub7sKeHCLhjsm5bnv2GqBHnvgTeRT
II7Jnq/ZwhuRRpYfwa8E95FIeqUNoDn0WSml/bXuUoCe1hX42N19tvddlf1LTIil
ZbBQ+9/OUeOt2GgNL145EDdPTc3Ex0y4Z21QNAaq7uZMwo27SKQtVITRV86KdAYO
XN5EQo8r9ZqSIc7IfpEeVjqBfbUsY2sbAcdLTn6ROvU5CPGq/3tUh+hKhLlfhjHx
FZcBvJtxD4SNdNmH72CiaXRAoCmLvOXyz5s/irl3siwDsgL9/QJenUB/BV4chyfH
8EHZvHseGiyEPp6ATOycuZuihibzgATWi+TROY8P/cvqhaCo+yYAQrlzelHKc8zf
1VgGQma4wM7FKXmNZErLCn+52+P/4z8UHqVRPt6JsYDi+d4d3U3829DqOCW0LMXU
ARnKPpTRTZCfbU5PANDjYHvLv6sZpxPLXzukHTNbGx56zPRZaCv6fKxD4VXMN87M
jBCTqtfXZlbz6jyblSLkelrCiS/ZK24vSKt8y3FOXiev0tCeuU47GYaiG9gypeLO
KMkqgdHwPRC7pWNunjQIEj1y5UZWLM/1mHNJUxRtrKuiioead8tDscR1TooSzh1x
lIAs3NeePtwZb7odCwjKYu+qJxktzm5JUcJSqC2fVlShIcgpaHuf3TUNCWWP8MgM
8F58aOpW7sYnQwOBYSLX4B35XgcCuxQdpuebpRuQ33i/cHV1hhAwVCtoTYYluaR8
r6Kv8fxCbsp6syzQzWMW9hYz9Ro/6M0gB7Zc3pzGxyEJEWNJzIVn7nC9Om2Fk5fW
nnZxLbYvSpcg/7jIaTsZqDFJRjiBWRf1OYDge5TtUax8Azu5c7X8ZWc4lry+frHh
+a99MUe3yFG8kdMUeGz9whibNtpFLkCQO0CCIfQ5YfjHApmAI//VUbyqRfm194Lw
zp0Tk2qfSkaejuFZgMQTOB+PKSOlzGVRdD7yXY3ZQpHpD9/LNQYIANuTHCXYxkRe
sOgdwEX1agoHybjG8MBsaeH8OyCewraZoo37/uiqf8uEeNfehwFnzdnbvGQM7Hqz
uSzxzxTr58+V8LOJNBiJeL/HYsNbDMbrxHyjetyZMBw1FXtjvPwIrQA0bqGRBUTn
w/zO/2aOnILiUOQ1YRfpY8sGTkQklvBTZKyTQJsRcyi/rkx2JfT+rufo7BGeX3VM
QRLT4O8z6pMewjV55jxz0m9MOr5ViRO+bDFSxGfKZWoltdVsoPrYXJBG6JeH30hN
ggRnPK+d4daDmY5hZVfA0UqHK+NBbhMpJ5uRjmHPhiYvMNUUHQTj8GQEYNhtlOsZ
GV4E4YoISXKY1UbX+WygEW2hPUX+k/nNhULCzX/jeo/WVwDjGtUj4r7C+Eqmgc6g
4dpbUygCvdHp1U3RxyYyO2YVEegeFyEfZkjGlZZ6uIR/IA7QUEyeN6ACfwGPpJXl
14Zk+bS6r4Rdzd3kVQ+mJqNVZK4aArFuQRuIPVOd0P4sfYqQoR3O8TQeeUynbgRX
DiF4cBJVURvMA1NfY3Xbr/Zkh054xM5oKng0LhwV7AfocKMLeSWMqCEgJ2bnr3e6
XyMW5o0fswU+v0Fv4J4mi36p2oYsQM68AKI85jRF5dg1Kp8jOz0PCjLPzKnU3/sb
BHzAh2JEmP0W7RAKnzrfMKLQ3LBBBWlFdVNy+wfJqlzcXl8+lwlSflWZyNofQAsg
g1KjaLoU+eUJaYGvAxh9QVJXbuYVq7vRWRuECNvDLRehkVGzO08nCu1r6aZ94j8C
tz0yiKO39i9xE7YWTGoIC/TjLUvB4CPPg13yAv9oTRPyKUW1dASCxeSmjJt+dnWn
IN/CQyJViDxdaqdVvc7sOE/RF6PtwWsf5baFigQju7k2OjYN0ARUZ5pbypG66NWu
Xt62iBhveMcNUSEvnAuCdm2pcHO9WPh9ewy/QHucZ2UGOFDYKEEPI4QkwVMlFKmf
IQFtZ1QyM1xtrTXPLHjPl4kJiJhodkpkwkrwt0k9WMsP1AoVL8bAvbr1fIc1nAD4
GGGrGmfZZNhMX0y2TvfDwHgZsV5po7UYGmucUVaW1i0k60R/A7TLUC83v/Sk4J4p
tLG78Y7+NHxgaj3w0mGQvMlYWw3333UrEgaZPJl+7ObMbHU/uTsZzwK0xMbfVHHf
2UcQLvyzd8YQv7c2gv9eF26s+VdjBvqSRJ1kprZdmlsC6Y2hKLEZu4qLPbhNq2Dk
XAzh36pp2wx6PsH3wryydG/2Gcq1FqD9gHzzEZfUPod2Y7P5cxIHDeKjaaEmO0/Q
lgesSbSLF2ugJBvVVHfkD2oTDIXUHwmMKofxT5HoDPPAjmnSQF+UolTVDq2do/0P
QuG+SdH4nl0yr23PG4oMvzqJxrbMsry18g96Shma60AcwxEzcDfXRHBAHXOMX/eP
KL4kbBt5nimoJB36wKClfgMB1RExd9lylRs6XsV2UZZccUIr8dCSW5woF6LAW8Bj
9LCMHFfbZdTdRoQPr2mX/RmbBjCGCxwpMvcPfV6GEtikb2wWl4oT3yUBrvpGKgxB
5/qs88WnC0RQ9nJzYAXqn7IiQdjOkWlGb6IJRmaqlmQIHb12jkwi8t8j9SO77Syb
r1alj2sRt2Dc5vaZkXZWZBnWrEEHqMG3NyiVkreQYb4eZqa3ku7P9BXxjHJy+eiV
PvDEkhmIQgoKMgLsZqyQfm65AvixLsyaCz/U8bTMdNkb/xjFBYNRzVfCcOIPTGZP
JSUWiboQkix53JPoWiu25RtoZR9mi54sofRT2p0Yyfi2bhuYOG67k2daJMFfjZYJ
RUTRWitGDtyWA7Z+q3Rl22K4QKilhAfpW16I8tOxmQXMlrVAb3HUx8yaLN5+HBsh
Obz/xEopYM7lP2/NlVf5Gz0FFU68UoIUu45E7L1Z4tg8cJ+SA7PJFx1HpQJ8gQLw
Jlm0SaEnza2lvcr0AMo1KfdDHnc+LRnATM5R5szT/VL+nPHnOBaWXzBPLSmYglKI
YLk2ausDjLABQcnd7uvVE04ch8Xhhz/xr/kBHQBlzvFwIvv2iHDnUzIlAA23EsZv
/G9ycxkg61IwGVeLG2A28rnRKb0WhDCHwaVIlOgY7owB90Ycsxn5+tiuuLLONWAi
K3F5Mc/pn7xJD0A4XMhp3zR/NGd5ikKJn6CT/Tdubz5RcgZrBUxyv4sYe+Ajdxb9
7A7u1PY0/GYWrjePcjPMU44DQYoyKyowE40G1X1KLCvHDrVlDFt2tLSnUzSTfpSQ
jFzIzkB7nrGq5D0AkzILgajXYdehovlAV8BePRaZtHtlS8E5TwqiIJvxTQ2wPy1r
ZzC+idblcpzepKuYH1laiWEqwb8MZxMZa/73F14pbSLEj6rjYgjjixAAgPDHdyyE
PFuTg7mMO8JtcdJCHmIKQtc7kMbVfOajJ27tQ6/gS6sRR706HTO+JzNL6rFtMrEw
mWl4JeRJZYJSKWm5urnLgehb0gJUN0iVDPGpknyorRl4GWbVnn5mylgdQF6DzjDh
f0/Jqfz54AZY39Gh/JKQyHWW1JV7SYBkfgqY55XYli6oEOMgIRqmHLb+SPEJGuRw
XVzRNDKpjvO5I5iTFoDtabcLWRj8XAUHwd5ewt9VkmgP+Yf6jeURfdzGPV1DRDTk
L69qb8k6iLKRw7x4dF7HaD84yke8B/1s6UQskk5OHuHOIz6SwKsg0Sy0wuOlelff
pCJTeFDIKpcQ2UU6aGEwXFPhEf1hNZRiHhAK2hwpJ+WSG2NedoJS9y6dVUS2ZadH
3ssK1JmdvlvZGDbT3N90a/ktICY5Q1hl+KpxLjv41E3PBIIDInDd4mrwZhGTBL8j
yRLflNT3ATrt7XXE7yQ8aPb4y4legIuRuWSPeEZfKUFT7bukDPV7D7XFtBefux+v
4v+KqajuST9aCMrEusG3qu5GfO6Mh49MHgoTqYiLrm/kluoMcyreKEdxHINeTQJ3
//zl6owpOOQBpy4iY8XbVZbI7zny7ZdIqkxreEMuk5HP7P6VB0n6l3bd5Y8PdJ1Y
zYHUtMgsrSRAn5+HHigXH6viFucZR1xYyUPANRtTzw271bJA1nT7005cR+ZySv2C
sIWBZvBwBieJK1itjajcZ5yn5h47W5x3yEZPHB7egTz0OPHLoeNRYnCqTzVH4AX1
L3w4qaCN7AQMIMfhg37tcjq85XtClO4fmqvYGCs+kS+rsh5EOPk2W5gh3988Ono/
ddJK0B86XW+D80yOE3h4vPBHiBQZg11zNmBTSMOZ7JtMFqQQShP6s2Fjv7+yohbc
IGeoq6nlm2JJVbBYFMx5RO1WvkM0MLByp0pbkfuzoLceMf17fEHxrFNPUIfDUAzP
BnUFgX1+z9cWgs0a0R+kBDK1Hfx1rz3IqInqQxkTZadOeL3uKlqxcTXhJZmrvStH
+MOPH8bhRBUQ4pndAJfrx6qyjlEWlxMGxrbOK54k9rqHRJ4u+mU1N8cpbc6yJLiI
8445GqTmKnrFL4cAYQYl1ehkZAMtEZBTthhZLjxEeL9l79Hb1e3FMEJEIRmbq6ln
lnU0/j5Um2gTHS7ZDK3DGynn7wA3RdBxBLJ+bkdmLEemRfFeF3CfaB1d6DfVd9pl
/Hgey2EeK79MG+r3P2dPaluYJ7P6r3fC2avvRmi14u1uKpWr3exvq+OQ6o1bnD0Z
i6gT6DGlNBD8vLR+HYvIinHbee+X9VX6NeSkWTlDlswRPqLLAVubrKqIGeyPajFd
b7OV9Ycu5xcz0lomKGGwlQ7b1kaBmu4rcgf9Hde3W7ZfVb4dioGvtRzq6VZS88um
tv0qbb27rPGdE2x8jYn3lqUSWJqfCz0G8W4tC5XwKxW3RbSYL7yrQaAW4TjVGsKA
MHBXbM6+Cf++4PIr6woOzpf7wfa8L/ciCGXYA/U5l9DYDA4d+ajs4O4m5BwBZ6H2
fbFsW7EMEmF58g3il15i3uhOIGwaH6+dhy96EN/EgtYf/uxz5YrrqgBetaJvFxnQ
9RmxeOJUJX/tOn0EXQW/f3eLRiK4JHlWbl2mHmYTg+bXITvzuzkw+STsZ1wr8/HA
9B9+qvub0IS1oNrdHjHnz9oJKQTsplChasDd6u45n5Tlr9Do1btDcpwUy3ZrFFKp
Cq824Tzw21BnsWeteK3kwnBWrrX1FqNb9u1htAuObzTgzqlV2kL93NPlk28KOyQR
cuwd1Bs3tbUSwBjsI3h1t8t2dTdUotR0DFE+meNz6U0bx9cfjabMlqhaTW+5fUUn
ya6quckvXqyYpt4OXDYc9mAsEYtX5/Ozdt2qibkII7sxaDKVMp9Huzzlb07b5bI8
Mq+/9BersMn1AtLbrjQFmc2QMzVTxANWiqPg0xxu64Ra2QnX8TsvRta2YANoQ7ee
xfLCuvKwV/HlmKd8KOtsed01H+G+MnRLUSoisGLLXu7NscggEQqD+SNblvlZReuh
b+Y/go3bw8D32QWsbi/Xo3rmsYsRlSNK91/H35P3E070x+A+jVF+cECl08ko/9pl
yBgWzTuhIzLsJwcnsOiRKQNTpqhhE9wWT31VTajOoIXGZA8WnBZ9MqDYoqjQ4wrb
IIMcSn9JOPXU5+Co8WXmw7Pzx2d1pA/43GCfAYaU+FvCzkNnFi6jqgx2vsIuEsGF
9KfsgirWQhiToIq9AN+55WFO32ejTuJMDjJZ46oCwHDivFCkjWQrCetTAgCbcMbU
HyijovFLnFZ6xeTB2hbA3kjWsDoN1xQJcKCe7EKOSpUi3GkuKidYNDNEbpMFDUpj
Qe0pft7KA7WcxtIivBGoz2txg+MmukwydTkYv7G+c7uq86bTDBvYQZp91QojS2Qq
jdNI6mKKCddmito3Tz53ZzyZVcWw99AvOsOK5o5jC9smjJ5gK2vfzNNlevcHr5ZK
GYF8qYrK73g6xTdvRlo2MTNz42plLX9M3ITgMs003Kl3SIrbHbKnHIswRgtZ2OsG
rX2OImZJ2eXXI3kQyrTBtGjqYD1uHxVMOXsrlQhkuKawIQvvrTQtsh0/+3SOKw5/
pFeH1xmWZDxWdyu+7UHhYom+dLwCRy/oGm+h4vGZuNtxeCCbecMVgojkJBlyqcTP
ML2bw7IFvzcs5xydHuCqX/dmmpHZCTzqcVZsJzVAEBGEAoEFUcGmKY9rz+nebipN
0J8ADHflmI0Mhoss6jTsbHaDmxRGmU4fiPpfvo7MEwRoVnLV9OAyWtXRwrp1Ewpl
k4o/lvpHMsoNj7TtLkwgrFkr840+vFr2VyXB1ewdBTpjAgcMwgP4EzquVOQ4qPPz
1oYUWsjONc07Lo/LSdPtSMzp03M/jYRcfv/TwkVLKCDgkVnICOGBh+Uw6wnfCqNc
dJW+HBLKbYjJWAF9EHhqzcZMFn3MLbiCZt0Ea7k1GqOnuuY2/3DbNnPtyfeQRKe1
Z5MpTxMdGd48ghEb9ju6QR8Q1EIZ0Ayamt6jrtxzWBf6WR4NI6S0yLozInkMM42u
nGHLgNW0PWPh3va18Ipf/ZmUXzH06+vbLwlbXeAWXH3J2tEBC6PhlxFICBzscvHN
gvtpjUiW7RRnJYK/aUOmLYNZzitqNhu2fu9ykNDourWJdhDrBsqvjyUQyLVkbgJ0
mpUQhQ6khUHyOXvf996Cw8PvlQ5Hclb/9PvhyPj2HJjyKv6QAruZhf2AKeuFIVtS
elZi86fEXowX/Ey6RzzQc/OPV+32fhM2sVL0TPzWjkfb0dBmWHEscpcBAKC63AD+
bYNzEAZrRrh0M6hOlFaxlPmKi33Ywyebb5W1L2VKf5Spmn3e05sw35852A6idWWc
xi07PA2YMd94xRGNYstxxs6G5eKc5DKhDAruMsnLYF1EpLAl7A9tgkaO8zuafHdl
2TirB4EKWLOb5RsiETmGnxZzIJspM4ppI7U0jiJJO7rxW2qxZ8AyQEetiztf0SxY
CMDe1R7TGV7JtlgIziRNC6+4AvyHfZNEsxil7e13UZkxbNNuEnm4wfVWGY944+gJ
kZ4F8RvtTp3pFe3v3tNtX4/I7EiJuQMl1FSrT/PncR40Dcm75P3XziUnXWfdRMcN
UX3LXWhjzLyyKSCoEq49V1lSltOuNISrNsL+UXl4QrX0wQypdoSYiLi8RalGF4Hi
goqyirjAY8phF3SsJJYBsKb/pZkTIbCe+ru423paBwqqmz6f8veIuTVPLBUuPnO8
jPE8zFqKw+DxOf2KDmvnnm9RQEISIotSkv0bE7CqJn0hA0GypYqOsjinJfWJ8DpX
UGNeD8qSY9CEu5/IMFPLAimiZwfgDCyKB9glaJ4Qj06QTqxVQf8//avUaCkFBzy9
UcEN/+RMhVFHrSpiQ/me0lM8ZjUXaSYvMmgrnCrolvIl1v2ehtTa43/OMkvfgVDO
k9LTo01q4sxMQDLchlBd5tPiS6q5gARZmL5VhcbaLo38iflM79eVMCDDN8OVgOH0
eqrSckXj4Hy6G00qCMx4t5shg2mXX6iBpQ2EW5b1SY4JElYr5YowJc/tDSC74e0/
wZvXvUnrCUPHDYENjnVPJiiX9CnZ8l1c6YK3pHJYeq4F+uOF4QGzhVUgnR3f7Pyy
CQxUPNpVnc3fZmS98UjIv6aUwLxyoIiWqBIV0UNyQvzVgfuObfqZgV4Sj7GqKYPb
okz483Q9dqNQYsqvorvpWO8QuflY+bhF1MKButL+vcEURjBMxkU4PRMSUK9T7j2N
ymUaTr7wiTCSuMbvW0MohQw3j7iHlbCx6SnisB+fgKsl8SHxZQtSUgGeUpIb0TmA
Hz0mCIDS6jDvqPO/lH10O/Z01ZlAf95oIv/ZSsMd8y962UWH1knr0BUipfYhx5YK
dmKLzvdzeGQI+K+TCGefOZf5Ii1XMFzWJFUXo0B0AzkLlPnNzHJegQwgdsFOL04y
QEGOyvJ6S7CygMBgPEtS0sgouqRSq5sSwX62n8hggphF5mooNfnPqgWzxZA9RKzA
Cx7A8LHqiwG6VVNc1oaa6BLsJdtzHJSAJ61VeCqRAeCDJ97/J2Z+5/lklMKiKwUU
ajh1PSYyylJUWGszPUCptrMqWpUasU5jTvlr00fqBN9Pfj5V0ksdeCRUl3K15Wd5
dYq9fBPaCh5JUHfxQ1pxLAXF4j/VtvHekTjAlJr9OVnHYzE4Czxq+pBviLPbOmYY
xdRxu04b6C9uGoyzTTK/Jq08p/ExM7+7e3zvaXLb7CXWD1M30pZtbNzy6pP8YG3F
oiT7F+cYWyrDfuDijxfZOdCESgBeB6vd6fV4WzCyHU595EPr8GWcmSSqTMNMLK8O
+tid7cl5I4nS+0UhyC2aXlY9d7ms1+rYrZ8SmbZC/UZBtL3DEaIjQvvfXuWz8Jl8
MKZBhQIT0UGRWmBiHQtyQ2jRIlTOVbCBAczz6xG7smHWwmePGKXAUAi3Tt8N45cu
tjnxEFVmc5r4yt0uW8oR1qJ5Ow19P2ZpSupn2FQsrVmw2tFpe+T24USA8TvMaTiI
wbbSDesSkybfqOK1U/cy0N+Po2Iv2Vrv8kjeYMvJdm6DWKv1i9bS/hrTT/5RMDSH
LNmyESB+mZUjL7Rs2EIboMefGyrCOyM0LTy01KDkTB78x7PL07GlHOBQYELaHqIP
FmycUSTo8TNoUcyiZFu0rR5T3YuGA+Q+YS1+L3Z+IdSjUJt0cEykKwKHTPC+iFKZ
MkN1/e7tqo6AChWaRcfa9T68dLEKX0AqVpgoDSwmG6duxt7yf7A3sGKA1sbul+OM
98CAvtT4TjSFjvcdDdZadHvNYM5y/1OVsdLziSH4TllgBepmsaNzMeze2rpjy/oI
yuKhFDg005rwvzcmIAKUwy7HgC6MhgIa28NpJeW8Pz1NK+DRYALLtqc0QPuA+p8Y
nyQvICG6mr4N9MaNMoy80AbW4Vo9H3agimlZ9InlW1FWHBeNAGOuhHNt1LIAGgFi
ZNv2MlTIksliBYcJZLzdn6gXr/s/IWNpy/IiLads0uPJy17smdPZf1K8vkaNMD9Q
QBZIMYTUAv8velWG3S2g61vWPWOJOeJDPTGnh34sJxYbYM6Ctu2EiNXmPXXbFkTV
i3mS82xCYvXCibRXBInTNzpL0xENok/vqMm93OB2+pj9tdNMwP6wA6iRxO37JLN6
pwxKU+IlWNC6USRPL7U4qG67tZjoTvscWwRxhoQEtg+iVvwQYoy/knopoeconaLV
lSCVZSNb9dUoRdwunp7n1sTkgh9N1NI+3578NyRcRFDmXuLfgzIkZKmnjOQ8smY0
nyw7s5unnUWL/JI6JbikzUSG8xuM8HaWAk1JCH4rpar1DrkpNEbK4a5DJHaPpc++
m24rcsAY0iXEHMrDsCLhrBtvD8E9PVTFiYLmRG41vFdpgD6XB+bQxRAJUSEfNO8P
lGMaP88vxh7x8QIdurjhth+BjXvNoxb8F+Sqx+urvbWvzz3H4zmBD1GXhwctVES+
6jRQNM7fUIaJPT2IDL98x7PzJ4Olaq04dEGja98epKxtfwe7/vB3WS3Tv5UjF+68
I1rF9D54tUhF/DKnCZ8eRPgVAZncDsKTzrh7PAtPkCr+jEzuk0b4n4zA/1MqmtNd
ObX95yCq9i+Mv8oZF5/6MLUIuPRKBGBIBB6hdO3UrvLafmadpjDRbkIUcS5FjrCd
EW9VJgo4Lfgin23J30ttx7btPVKgEOcwwmVI42DdcovSJ3hFcD3wWJXl8ieFNeoX
gBdQA6l5lKKBGC7LnCmNm4WJbvOdENe4OXSFIpu1ljjnw5hwKHnJmiqamZUvZdI0
riRd9ulo+u3c2GxA1hYlN9tXLpAN4WZOgKqNt3/PM2B9XtlNgG5/1fDmJY62MECo
IYamypLyo8luav9kfUUwBnYIXuru5OS0YltbG4vq0OP9AA5oKAVeD4oziDOK2HjX
5itLYJ8bf+V0/dg5NvJrbBRfKiBbYcwLPVJbtnsICgGncT/kd8qArtM9+ka9HxGe
sjXNBvQIWqOKGBBzSbiMnGI6eKVkYUOkUDbdsi2rFZiJNfmhMii3rwUlDbgUcgcA
qOuSXZ+8FH9wjzryVLyDX/kFSDUdScIaIJb8WiqKfM34LB0ldtK9zLMFf6Nb8yLq
rIMZWpij8Vvdhb1SR1FQ+cE6a4ylsUva9oOB4vLqHDu8udN2Qo8fbLR2l7z8sMc8
d9kkm4cBDTKWrMOKSjqoENMZ3DJBYFZqCAdYLqRFQ/gl1PZiex8zmOX841WXXiOf
SA6zD3of9rWT4oIPUXaI1y06R+xzlivRKmLeKOM6neC49m7/sdutlClok/89Ss85
CyIcWZzhbcTjkfznWEojHCzY/D1w1uArNi5nHLkiJhwJUqrGgfp0PR7i9yT66e5y
SQrien6kjXDu0BwPgvo+O+kSrObmvVwe8gERPUWtXtJ4SpzVezaUTRa1xGVQz+PA
dyZuwsFdae6Gfa0r3f8V1t2GyIcmzweC+m+gQ93HFuW8klbqv9FnNLNotcnmjWge
mogk1aYAHXCOw58axa88QGdxymaUoHcZuCk//295VxNhOOhT4DwKpi6RjWaVlkCd
n/rmdSDbEjc3g692Lcz6Q+d7Uql5ca7sWDwfmuI2dJPgtcwMpaVwtave7GyovMiz
PVP3RehVhzv9bh+uc0ySh6jjh+iZ17QPVvTctRVosoQkO0t289FFzTHRNYOeU8kB
y3WCkr8rA3ACWvAFhzD5jj+J9PiZ40qIm86MDjJtgP7CZv0yYu32jXwbsI2Gnw/k
8EPwYS4EI1N/brbJUuFy4ZGNFpvn861UbSM6JUJOLZd8zThv7j6v12O6Zba3OvL/
4ocxTrYMiSJvGNzPlBhT3yPQ7YbTr+++PTQJ/hKDOyTrXR5Dh8qMoVo9To8u6bjZ
x2EGBb2C9IUsYO5WdtQB9ah4ERRzV5/AqUKDSWYW9L6TZK+4+WZlJnQl633X/v7t
z4NToM9ApOK7Lo9ZMDZ4p2oN+vDB2PwDgUqkjjAqusmw5PiFjjGn4nNde01xVA0f
1NiPipVIwDR0B/lWYtEKmTr7yvNIlMYwRJCur+mEYLSBSdJKKbojluiI2UvAzhqV
/EscGMjoZDxz+ncZVOtkzV9PJtrCzwfZ/Acb38qkEfNKoTX3rXh0gQjF6gzNlMFs
7njHG5IoR1cSH4gwytiGeTp6a6OsXJsqulYfvBRZHKq9rSzculwWVx1DFSfVRYY0
twb8ZAUk7F0ZKjNrYBekr93Soya+3i74RLCxzoBNOe5WNYwK4SxXdL4q0ZHMCbgA
nVYQYsrE0k6dWlbSfr9mn95YaTHZLSj+Iv1V+t4uu1CjcC1b0pFBZ4uZBwWeyVSz
GSJJLC+fdwVIelADfJjynp9ZoHIE8tKCn57uAdB1kC6roj31vhkB+s25rDUS7KOK
T7uO+v4Np6IDsuRvDxU5QlYd0GAe1gJpMnqZ3qCDCESnWpCMsK9j1VV4gmXgzRdd
+DfBdl98oqO6+gxWG32Cnwv73cgR9rn3ztmeYWTd995Cj76afIcF6dy/ZQ6qoKUk
NVy9GP6GoXjgDHYk1EjFGOJRROVG9YHQ4mYEkBdc6lwHJK5eAxJjNueFog6HDKLI
JGFjTWtmOqq3QAWbSky9oPCV3sa+r/z7GoY4y8SP9kNR8e0lTtcn60HR985Am+OP
gO2YTXt/1dXT0pRxpovbd2l32Qzk3m5qVeVvkizsiImolX8SAFjfbNclWrp9VJC/
7qvDd35KaL78i40boN/921sIkESpWSrFE8ZeTvt5Z5/HF09VpWFk7nnfhG5/uKCF
E4PAQLhX/tvOSMdO+Zz7ZFpAmElqle2jZhQ+CjfjLovN3/+wdU24VmIuoL/Mt5Sl
SL0HN8DFUJGOCqnyPb22rj+dKcL0bBMDTCvdvrkSdH0C5z7chHOd6RgR8itTBmw6
MZi7h7GJPfNHojBG5Bkt3geLKNS3jPWKaZCQB2CaMVizhOCPUdDZZv1OclJOGq7A
LoerHuVKWJwopmfTn+isaqJOiOI/5qPJssiTf3SSza7H8No39LzIzud8x0reZZBD
XKo5zY1xcdYD7JieB4pNUyK6XyIaYpTV5moTi/cQVddtDpewvF0ab/bKKmkkdYNS
nlwzW7sXiX4AYdGy0APewJV+wL5lumUGNUgCdSuUgdjV5rtfReQgt1Q3x9mPTfs/
5ZujZ4/gGsUFFwqXjtwTMYVowpXK8zaQpn0viHrR0FghY/ju25pWXtS1TzmeGELy
MNUb67Dz3XxIxjtc5J87Z/a5ZshgHBjP9DoGpe1s2ZW/VrMTHbLbS4yupvCUiHAo
yJJGV/j5zBhOopJ0XQMVZSNuzXmsweNnl/w/dilcEPF0KdOg4hd493wG/pqU/nT3
E6vm913kHzycN0ZUzGTu8iFpYWiXaFskoylA2M8zWzxt4Ei66jhBJ6u1a7QRvD0p
voFHma6A2Q0xof7QW1ULUuOIIEhdyGH1UW6+mGucIuYucKidPilYJ+bYvHmn5oX+
gTybFTos9fEvtLdpJl+Zkx1SpUjeV0+PnowKtN891isDCXBh1/A4aNXie+4dAApI
4PSNksRyLGqQu/ZM+Dcf+cEq+8EPEJQs1G9F54OhB8gwx3c9UUnKQNMg/vj5ddoB
MPm5msLjHETLsEeiKneOlRxkBpcZnab4MeEw0XSFLVXBv5raLiFCKOfSqAcNmEWx
mvWMMEbpBkhi0n/BbZVYqKtnu0Tt228zjtJ2DLHpzbXEpaUrzkOuucuexN+4lNbE
mPtiQGoZTUDGgbhoeU8D2ruWiH3lBni2uaKBujF3EFtoADtqwCpVfWZb+nzCN0ME
8BWNDOTlvNhzskTOp4k6tmeuvRQHjjO+S4agIbUrGXiQkeowY2+QQjQxE8g5Mwza
EDqEAfZtFGCfHz1X5hKXk/dY686r3OuurnjGKHZBVXrH3a1I8O5ZA8KBSeePEUDA
e58Rv6cY9abSTqPgLEqcNtaQqZ2kg1t35Thk6rRfXjDqa8ZvaINeo06IjPloi9Rk
e9g2Yb9zVXcdYsHHjsX3MMZGVK45D3IsS/h9BzMryYeyr5KNZtfG3/aEDKRFuxTa
RsY65u6Ufmoc/d33cBD4Mvnxl4QEazocnuDXyC3eFSjntpnITXd9bvpoDNMXk/c9
5aJPghwtCA6hMbUyoGsoaHek2v9mcJyEp24SxyO0eK7G3U1y8Ghq6z/12JyCwuiO
3hFCGdiGNT+DED6uxJQ0qvNJkddP9UOxjHeOgOODPlxWtbnzyG0RztT+r1uyNpey
e3lB9LFxGtLqNxbJuxB8rfOr2wyMqrSap1VB5YPSa6NfzuNGPdJJ7gFLVUsqxJLa
bjeufqR7XlMgg4DbmdyCG3D8I4w56htH1+fqLc19URFYx3r6ZJ8DRinNYckDdEZ+
ZTrR1mHbKJ3HKDpzi8TlQtfNR7m2mQUmA23G/l1NFJ2ZZ2DtdhOGVat3zgP1a5Xv
QXa84k3aC23OJDT6+ivAWIHr09bMeSRhnwYVNnr+oqaG/eC+q7s+9h7VucIiVB5N
L3lK42W3w9imvdSICm+532qmnMTz++0x1NwNLAQyoDVe2cFKQzGkByqCXE7juXo/
nx8+ic2VQ8MFWcWc8nq9ph7h7797U6Y2bazG0At97ElW3VH0JDeZL4Gc2H/38cEe
B5whP0lk90DXS/FAr8AUpwGsLURZ+O4M1EC/gmjY7YAbbXZceRGlkZ/Sg9HJhpMr
maRTDmKe9/lhqlFFqZGOVJdWesalJ1gnUL2C5oePsd+NVqeqUykku3oT6bBg4Qav
1QmjK2AIhHeoK71qTOWrTHx5nmpumRM9WWgCfzSo4BTdFtEhdkDzAbV6uA1ynxiS
iH8fvhxi0CupUKCa9qjEqibzi0O2kzIckr5YxcqbjD6c0SoXxLof+LIEpXttVMta
LUs/CufZLHQG5e2EWIGLbfgnhll4bMwpFxm8b9ZiAy1lkck0+f3p/RbRUsZ/AM99
5Vf150cWgssvTDPnHPIuRXrXRGpNsMRx8j9T8GnrpmuPti4ZLcYlMYUo0QfN4F9t
DQIs/tKeqtU0buvQJzIhgt80dQ/vfwvGOtTAs7S30dLKVjpnamDCmRislsWZbjOg
8oSVpZQeh5NBl1ZYPzt5Z2pyNILwEj6ZfaevBP/5sxfJtlBdi6yv/5lPIphLV378
Aj0ouqgGHKTYY9y6I3pa5n0YxjAO8HPd3P9oe/dbfirEEx6KnyLfzgLAQMjmwMZi
WVVFa64x4YC+Fe49R0wCby1vZQJcz+x5qWNnFBhOjzeedLq9r23y5EC1SMiKLgD1
4Cl/sLvgQv3IZ2Vu/bIfsAyT1KsF6LqEjPv4WSI5g7hNF5OF117Ku0nEDHBHnLk6
vJwV1csoZCAc4hZors1TuIthJ9xIA69Ln1QcXREGBPHZHPkvEij3P8n/P3eo9Cb+
bbO08gs78nIkMW2bbyqWvLjocXt/oy3lwDYrFzTk9raYIN6gZzsFfGosEFvcDbEF
JvvWjAvIkPWoA222m3zASainG3aUcvDlGB8CcnzZ8//s4sweu2o6uitu2AgC+6AT
pzHpaZX5zWXV8QXm5A4mb+2nhHdcS9NIupsjawJxlOgiA4jeiqL3jFEMKom8mgOQ
xodI71hW2aW6M9qUOuxOJ5Dpl2ylBDat6kBOPi3VpOBRtK54UWGrbyR55q6eUkoz
qLeiTObZaTcyVvV74no3khpqh6eW/d/HWpvhdsIVynr9vP81VBaFMr1ocJD0CY/a
QT+H6OeP0iwsoKCg5+qmhKXYvk2myyDjcwX4B+74rDBF+DnnOkj8mfwACNlgRr4F
AcFbX4jWUSEoy5yHkZAkJPa1/DMoIkzKbKJX2zycULEmT7zXxCUNLP+hN2DiAdOr
rNxrwjsq609PQ8SYAXNqmrewk+8i+HKTpw/oGgBdApLReXnUZrP+M/rTGX8gBXF+
iq4Bpcip1FXxe+aOryw02AU8VChYXDJNhl6r/q1z+Ups1aWwjdBR82ZXV2TKhdV3
eONfSUub7nEhFEPxllRby1L4Vt/PRlcwMF+Tzvit4YhTAAHg8l8/Lcs/TlJ5N9mY
i7+zKUUm7A1tvjMuhdoJetpPFZIVKFSBw1Rk1wE+zMnhq4hsJd0rkgaq0UPBQA3V
uXZeJCsqwbO3NvLzNBi4GRtaDPeEIpiMaOIdnrrtPC+M2W9WDSjlDdSRBXrvLO/N
5ykeuSjlbY6/MI5zGzlw5aLPGK95Y93neQ/z5HOUdlSCOiR0PwGEPTcNFl+0jM7E
b6QpHPt2GwkND3VqprTAu2dAJ71KkjedHUgjO5+usVL+DTy1Gw4AxwStb99F19ri
VkMKnOMs0NaEazGxejSaSYBTPmPzfft8kFNB4nOBN3pIJiVjEJeEXaGFVrUPfZEh
Js2F/8cGZgJAzjexO5+7WodsbGZtT15jSL+tr2cqOSSBxwD2jB9gtBHrAooXHWpm
mfa4GEzB41pW7pEH//sKxeuQyz7pnU9oqt2PLMBCgSD8X6kGi0exsu12cAVJAqU0
6aya/19KbiTmTPSHBkOrdUcKV6VsWNzrJcMa5oOrEuZDQgbhHX4pb817cpsuF2aC
UFFuravXoRh2JZRHgmc4Rpj5VDU6R+9YIOI4ssopzlXWZXbiJ/PeoxUdUy2FWnhQ
m61j8j1dVzI0+0XJmNJ1frBmFsbWJqSLrnDUEW56Ubr/TBjKIw7xWW4NrbZLFff2
XOHo/+nLe5oDn/rbCrojak12iX5LfUI/0hqgzw1JN8Kg8Ztjhgv+kfs7lPe6DH0t
Uv067f/xkTxSKKCXFUnMVvAbx/4syIK8yieNyYRbqDhEEs/sCf0S65yofbP4BUtL
NZbp2uslLzEnNOcXir+G6fZVb/AUU1PMtnyOPFiQteWyIDco49PAhGQFINOdYSbP
qAfMzl5h6dE3c7n1Hu1eSgA4V1XJfYleQ2dfeiitYAGweaS5H1RBRStfO2iFlTdj
VXR5+9q8TozxKg9mdKA2rmzthd93g/vx0QXMxI3QvsI+3EECstavOcOKk5e8xAgB
we5/lYLB/Ur7go1tYQQr/AXSUahKllLBXBR6KPCFEej3r5uefzMEMIxAFbzy3B9b
sa9KYun4Ibi+5BajaDIpZNVdJB9uBtgEISoY5jv9OmivShnnD3Jop1hl2gLs5GNe
fx1Nw6uiNPXDRBpR9rGGuOYYBUXbSJljGGN5vDRRE3kog4Qg4i7sHK9NR6PaLzdR
33PhzlLcTMJlcUC1gt4ti6MkAjqZ3PPqjKAeSobYZjbwF5JW0myHRmSWiMKvRHrU
8Muy20jD+gYFb4Glqt3vehW1zWBBUcA38epat4xOpZsLaE4n+16cckDDO2Ehgafg
l9wui6JDo72svFRQNW5CVl8TUhnDmkWSwJWq/pv8YoBGEEO3KOT8yHQ/S/o3DS9h
fjZmaYcEVwlDOFzWwyw8Vl1hE8BAKAbSuqSym5W6cuCV2/aDe3wBxErTduZ4DCDz
3kvSQDPCAIfR2sMZktrcJoFm48NgFmkfm9quR99bRxm2Aiuo+WiB/nOJj26PIpJO
Pd/NDXKIz+xO/OOoUjptcH3mTIZKdTnERQxp4HHPHbtiJc4Hh0/G69C4WIIEumLw
X+5jyowAbI0+2NPmZmvkT5SLgoz57vZKk+DY4cMxkZcAYeZgfC6S5l22rnNXmizf
292bLGX9D7Yc7LI2pW4hNWaGbDqTlkcFo4TlVi8f1u5a4AaiB1KuLSgUrRZCuYYW
VQh9A1EwSDH1fkorm6r4RmUbLsdbt60A16oZ9veu8R/QzaCbMl7YfRbuvhAGtCgU
iM+fmWmuqwcuwABPWgKGLSOMBMbGr99rfxX2IBX449uCd/qbkVA9BOCQlt1sV+v7
ibiNP5qnFjqc/OWVCcNhIpgztyC27slXhvOvclexcKjmEn24Fz6upVYwltMfrjZ/
lztlAkRUVJqxVAEuXYgB+mki04YnFpScKURDZeZP/axgp/P3164e88kpNxYaW2Iz
ELqF4Baxrnq/K5YFq9JJh8FXbyIdEmO8k461QQBup5WFK/GoDtoVuQckGVOcFWyX
7N94kJ921qvoz/uQptolMohun6+R3/D5g8URTsOwqfs2DWAMJDCOi69sJXMVG3Hi
Y3fXYgpQnK+fZg27g7o9UK/kpdx42TCS7nv2wDf5HaBI3QaUCqKHlxMRk7i88Pc7
gNlv7ILYeKLJLXiFbGL61ya5F7NgEy2mwdCTHJKL4dSu6Z8w6ns4KHmInrynlzsl
tonlgi1Azve464rNXuVA4iGRXHXuZxsUdUCYUCDlDXm8vWAz7V7k8Sb/9k6+Z7H7
fWxpVqyv1iizFVqI1/tbdki+VqxsnGxdlM8z5/zPa1YkHkss1oyT6fDXXIeiuWwl
DDLC/03+JxpcHRrcOg7lumjV0Jb1hJDABJncvDpr8UxFAZiUE+8Cl1voDMmRHHqk
kiTKcPqElLDj0JUH78AzbEQDeG8hEj5yre69IxP5dxmXnjc4j3IoS1zERohZq7W7
n6jE/1X9npNq/u/pgbkjeuMgfZ/gf5yknJlfOJzX7VlpCbxLzCb8Xf3tvwBwsQGR
mpWDrJCOsvPujhdkqLp4RnmqGd9SRAGgbjhpc50JYYpd7JcfhEW+n88zsUjj22dc
AUWgc2KhuNogVABhqN2DWrIIQtRgW7awSjh207wmrjfgHLe10uTZqMZO8Po/EYp8
jW0LgvamTzoOLF0VpZqvO22Fba4ZO7+UtzCJpWqAE0f9lk7Bid0qHrzJPR3p4KO1
a0opiSB90VGpCXOJ3k2zVxwrXkBxGqlkFEo+TC5M4FY6NN1/9xcjrBYkVg2b/sCK
Y6nUTutWxIuxNxHeNnf02CmNpdAHSRWUOjfgP3y068vFiIQ1WubPAHmry3MkcaWE
mPN+LYN7SiPFMsMWgChzTimDTSE9vnKM+4mRLuucQVR61PM6EIEeTnZHUDOrpLEN
IfOI4ILsbPa0NLEYreu8VMVTpkAM9cBet0oJaULh+N8F5D0eBa4k6BjZlgNWkwiP
PO8zZmf9gk2Yqj6BYVdaYdZzDsjjw9jUROCU5jDsbrUmYE63nOcPLRSpZ3v7Pnx8
fC08ePNIaigb8yY49fS7tTEsC5c9qWKKFXYxEgd8j9NpBVKDnixXL1MZVvt3l8vx
2YC2Zln6Snm+818U4RQ/ltlq7rcbBtq+qPwmypdexkoiK0PEyG/kLtIvQSUsA7pp
OQvs994h/NCZdFItFJ+voi4MCKHS5gPDbi8SIIcbMWZzILICHcfcd5C8yXS86hhq
I1E5l7tHENWuJMOqrry79Gd6OfF/dUUQPaXKtaF/+EXGMCBQ9/oM5iDr6JMVINme
QbkSF8w9gOnqvOPKr0zREfwb4S/EDvtY3LfDSti/jyvNEhr3UcJR+t0Wg2IdciPL
pNuoUYhjjUikiHfC8cAoagqSeeUSYkHwrigG1/6nXpYQmk+3hrig5+BfSVe3bUXk
tV7+PTsim5cHTPvGX4r5cmASApnsovVoIR6qWdy+npObhOuVSjo09BwalICT7z3c
MwZ5tPrApYqA7eC+nqrNZjO2nggEEF9ivxuJsR4k6ZpoL0iMWppidpXWg3xQkozZ
iE8q9jGb+TtD2bbLMxs4ueA/h9zJ5XIFQnyjd9JcCFrqNzdj0yQuEjNcSnA2VTwI
enBBvJO/FxHwH1qB3urykkNsCnFZRImeeUpN4syZKD2CIItG8lceRrHk+mQvtozL
uDcBh7MeiU2Tm5Fsgw4OAPLbzC2Qt5xh18ogD+q0sBmcZqpO9UbZ+aTNCY78KYZL
VgSmIm7nL8YHPLNttB2N9Lw0sC0AKzYa7iuO13TRlr8XPbLrIVOjOWzEqOrEtZ56
wn9grcvbYrX6hf41iZ+oyhJbo6J6YgR8OocMnYyqOUfPFG+hPBw2SSwKW+gUTk1g
1GMqgHWjH7hDh4nmHHdQ8tSk7wZawbdRYzXXkEVC62Y6XIqfO22RsXoaYPOxEO5F
yjjbZws77JxNRNRTB7ISZOVhf8wR5Syio5e8X6+oMcI+A8YK/MGwTc9KaeAho5En
TNgb8HZSAbtb1LGOzujd6wq6p+KmnoDVQA67Pd5/2eczgRCcsvUqkNme8zuei8Kp
52x/E0QoHsAZTs6p41ag98WDTdPYBiyCEk5Cr385hitmgnDRgp0Miwb8aPokq0rq
YDZvIyO91dMPldMNRVRY5qFthm7GEwLxADd3J2ug/4khpXhtHGdDTHTSlVfrz+2J
klZHdPNEYoe4Ftl0CnQkivLc39T9+soFzjMs2nI02Ihl1ZS38iKI8IlVagjET4nv
qdt0lB71gscZLc6Y64lo48ciLCZaKM2jG3mNcDKsNl38wNEcEQsIj1zBa5+QYnSj
t/sXSl30bAwBVil5C6KJEXG09WKU8EbiDV2VtJOSJnwTsqvC4ouNeyYthI8l6tsP
n5NaErRG/BkzZ0s3PrmAP0NfpfCkvas6ER4RFXdibprU2c3uP2TJn4GXCnk0WFb9
3C62+n0VpAuIQ8QZ+5vnI+9nqHqhlT5flhPKd14idFTij0d1XYsflZ3pPO/+khxd
YOtfnHdRUwJHthR2/pXzZKAdF4VEulv0bAJQgG5bUVGYE9mzzKOmk9JvrZzlDGoP
YoE2zhDkhjygglP9pg3UWLdQ6RHl712XMe0KeF6G/l90F/FiGnD7UPCn59zrswms
uuwblTKhLzlaAlA53GI2fIqo/BbTJoM8XS70GiPys/EZ6ls2RyjQNykiCTlOexVc
pKOf99J94EQzdxY8r40OpF3BoacT57kZLdztLOoaYCD8qWTDFruc6o0kX4l0Ix6l
x1dBLPpt1CTuCBZi7EmxBK3n7otPTNNK+dsmWUM5xyS3y80zKh8PZ2kU/3LTTpUg
+DBq8kKaVXQZTscyxIQCCM8WBIc9sSkAPkHsOWDdasGbuXDOvzygwDCH6x9mOSfh
3NVVEw6QSZoF6UVcWlCD805GvvKQ7hZGzsiJMxZ7365ew0Kxa1s0UGXHywxttFAn
2v57PUABfZOKdZXsRnJodr6ZxuBsfE6cjr6V7tU1a5c+T5N9u0WwwWY0lO/ZW9hm
3Oo7HnDJYe77bQwLik31PKKrTxdvSD0spcA2e7pQKLOTiOmIg1UIE8Sb7hnzT+ID
nqLuRx/QwO1QY3b66df9eCfgS8xTFLe5ci18M9T1znpHqHG4LdOB+9FDS0Rdl0k3
6vN/u19apAOA0xP5LeCOvM5vk2Wu9cbnghVA5Y+v/lPE38v9HXxhaMG3Nb3RPAnh
hKe+59sGvpfFutTUNg6BP8J73VeDwSBfxrcvgGvC0MpnET0cnDnn3ftTc8kE+KcM
n7iz9KJ8iN+xPb7ioFXFk+h0sjRKtp6s6P5JwtoeCljuZOWpRFU3iywtrYlbsMYr
DOAEOpnJrxUt1RxuyC1OihD6bntiOfxB5LNbKHBF2IsdB2ghHmIHO5ZNAqxbjsmz
lEAPqy/PvRI/SBWfUoP3DThFazKGcICNAjmX87BD67tq7GN0+a35hXnkVq0xf+UZ
8ZIVV+LZa5ISTX8HW2GNnyxqhMd1QpMCfUxp8MOYiJB6soxPhaJKYGtLTzTGge+6
Z+jXWq6Iy253pvvh9bmUTU9pZ2394Ms0ACCqaHyRD3+iz1blzlgtz0Dpnuq+k5TI
9C6Qva6g4+6z/46pWgHqtCTpuoxihM5UwEgpjngRs6dmyKLYjwMt8gJWjixAwvNB
Thr+ZS0djFYXFBILqOdrynPr4Kx492y+Mrvpy3kYUOHObSb2flCVwKANxK+olILP
tHjB83VXQR4s0jAR9jB7ggSyB6GPd1ZIU3XfRlUiFo2/scH21X7UEXMRXNeI9CE+
/qLqkEXCH5eBV7x02pi06Cs4Amr9E3pvYy2TDlD1Xl4o0e6ToUgwx/+ac15vrfzi
AdIu6GI8zXA5fk9nuaCjgRA6RJZFV9Y5YbzXNWnPWqbJMfxR/JbRGpgGXyFEEqs9
o7FGcULNrONvefqGOrg0aSn0XLNai+qZxwvPt1LBXNlWLkU4A0F6WbeuPDqE6CLP
d+9Uxzh4p6Pku47GystX1UrRFGaDWKeTJJwThR+lUH3lw+JzKjrkXcLSH1Qtog+S
EoPpk6HJkG1z06sILIXCQuP3R+kUelIl5VnG/MMpH1S+qkbWR4/kHmiuS09QMs+W
iWpFNq0lf5LOZycPNtFiS3/2Ign1xMfZRfp8vFekjjAxJ2/EUSZCZCNFxrkBEOm9
XNVKwIKIfwDymaeAmXKPoz+RsusODp60wcX6P0sdL64u16VI+bL2NxPwL9LWL0X7
1A0IOJEwMeSa4PdtvMLJlvMTfpTGWg50fXKgdZvDXImr2d/VhW2Qf5E2rYh+Izre
2DdQ63sVbK0f6nOOt6Dnbf1h81cDc4QKM4L0gwiZ8yodJOumhfB4ahIKkzLVa1vU
/UzeMIwKm0gDoaMs2DguOOOpqmX9CbgwOdpCSLXl4cm7Pvny0NnRv1vFgbfgFxqC
RShJWVuvwKckQleCq9+i0T5mhOXkdzPqhe2qBUC3j/l6HfKcvvi3G2Q2pIetsoy7
XKHy6PrK2xRDr4nrE4HU0dNhOa0ovznRqp1qpl9v5NIO8j9unY4y1f0KYIka2kWZ
YnIQ+bxHg/gw0KdZR6Cql3FiqSSn2PWfkq/X0nAvWYpktYZfa8icWi7czAsy23Eh
IaEla0O/lQai2QNDD4UV5sJH622UMrhoQPzctR3dTk+iy/yK7eLZJXZuekGo/n9u
whdRBoZRhnQtAWs7arFMKTQyu3EPFfbBc52z0Dw0pHpTHw6ldSL/ZXf1DgtXHP7t
IvSvo4LisC2jhWXEKhGpzMgXskGDJTBTcAkUwRtIcNU4ZykShEkUmHkQliV/z4v9
ocofkNzhEi+FVefu1bovbqzl/iUMK/wuttgSgKF5pYnm6M6O+Zb/b65/hW5Vjik7
mEQIf6PY9OQ8mxrQlihsvz2W8D6wckl0Cb/v3niQ4lkwLwLIhkJ+6Df5wtIEN/mW
4rZGUefYQGvD/M6fdMYAsPNiWPj37aEklN4SiaLGztVc4mEUO+QMn4PcEBvl5DP4
LKtcU1zxb1pDXkElIfGHdK/5Qrtsx1hkzMP90ehJBCuiTPNL9US0EhksojTiHkU/
F5F8HrJhGEzReIuB0LpoTRmYCznVXS80OXw//jQXMSfbQ/54cE7nbd0UQLNTzqA3
0LfJYxTjvGvzRHKX5HH/7o6PSmjSLxyX7VTXL5fmZTC8SwXxmDzdO/vnUfkkhnWm
oHoSDToy6lSYzFwxo+cQvJrMsZnwnj1VixS0C5uFoESaX4Ivi5TBnojhQGPNPMIL
x4X+4g+UeMzsSpAI05m9oovCyB2cfYAcPEkcGEyFpLdEQjMeph1CWtkfoHU4ei8f
+RX7f5AnT7Zaq1hvyHLOy+phDHUvkRMsh8CCPlmTSDtN8Stmleio691jA+HcX3h5
FuHrf5LLvlGnpJjMqd5j0rSpYD4P1RtKYoO6aKvqPtAhAcGnr5it+809CFT7jJ8/
eVVOYEs88ovrWiDrNduOWWfXzpif1bQr7sLBgsThLcc7XhAlaM4juYr1F+z/+4SJ
NZ6f4aG0arW0flGfswybJ0MJ0h62zlmq80/+iwDpwpoo207cspD6WbFIS4hN6hlR
x5RUhiqepOY7i8ft4RvoHQyTakYtspQqjxMz8y7Mzbehp56Z+EfC4mIX4Muj/LNo
bad8//o/8owDQFa2C8TUiOgl+qIZaBzro32iA6kEPY6nDDbVEBXpIzht46pSBplB
P9GwZPXpN6eWSIlTpLQExA0lo9i62OqLiNQYDh0x3xrTJFnTkGwPjM2wNY2ml1a9
PFOtSro32mwiNs7Qzbv01Aq8klBqk4ZoU9xNHdQt3DgIA3vgEZqCSOhtjICFSXlm
m2L7hsOebS0JpKE1JsgAkuX92JK7zZ9sH7pldyrMFuav+jgtogLPatJkk/CVY8U7
fckAr2xrYHvEOxkVtiL4I8OZDyFGEsa5ufMC4yVccmPxQ3Nqc5qIQgkWUPRl22bZ
5QHIwY59MP3mSRHwwSW/xbn5KBx65bDj2uOrqYB7XEl1HgM8eH149ZuPGfD4h6uO
6UksQzgnrupogBeA2+Q2vdW97y7wTjMSFCx43XZ/j6w+9JEnIxgJtkhNuD6Z84hb
r7gzwDbm/kP8oxd2AkikWeH75jY8hJybVUqDCGNOWElzjWhnQC+V2NnVUYTgQpH3
MY/gAxPA69xQG7SgAGEIWVmAx1A/2jBxXz7Ly4GK4lb7cSeerglae/LpLuSTcmx7
XyI2qEQWLmF3bNw2wNnf+hq57bYq2/bym1lswJBKdDNc+FVLVS321hMn7YkAiweX
t+qyGokrIUS8lQMa+QLpA6nD3jI/mRxBsi89hRCOTsc8ifSnjnfBWpdZfaTmxij8
UTAGgwbE+xQ5ADuT/w15+VqNnluyw0XPX1CEvBdmQ3icHuKB35+g/XGujLUK8GNe
GncrZ7mkk7aKvYFyLHSmDnCujUkZ/pzvM/fPgV2wjGmc2P/ayadu3FvChVhy/8th
xJUhIqm7OMeq3dWckAT4/rQTu/JOTJLg8TBWpSCrJHd36y8qcSnQ2teQZaVxpIuF
DoZ4lI7JSmW0y3pM59CcMFSUDE5KoUnuSLhW0WTl0Zivz/2eqXUnEZdUBoCimKS2
FGXpCcI1ampmKYzLkFjTJvAsnu7SMyJooEi7pfxanuy1i/4JiKmf2kFNpEDEW/eX
OwsD+lJt28RHLr8PXrPBeehgVdzZu0vAIX031ooc7ze1zweLdpB8OgMjYFaxhaWk
SG34FP0wrRFKkmTRT9W2TzP0QVTWK8ROnJ83UyBC33pI78AQ7z+/j1yNvEPm8wT5
J0M8YHDi68wbKeCk9h+LBWEetP5kOHEiLBWEBvuUeYKKE83/sQSTln5OjeJyFUHk
ceQshLmAQ+PUkEAjCdI6HKNxLHHRWPaig1hEQafDie75wj9k80hVnXEVCoroJk/c
ySnJdh3S4dVf9tzLzKKXocoUBb6hCz08dowDdR6rjnpmhAE72TI0yZWuHAcjxTXA
Jss/836QgD5z6h9wze/Uq71whuSVj2dwSYPK8HVPyislIXOUK/bw5BG6ZihMIXl+
X6MiJ5BKhVhAiPWrOLRWF6K021ZFettSH9VeSTC0nddRfXIsxqBNvPLkpOAKAvgC
aDpWm/l34lkMsvlN2uB97Pqyp1EiUcasLLSknT5eiGD6Aec2RTaVCMApgxzDBJbS
zl/TqKL9tZS0ZEeHhRn/9uxURKJqKL9tbPviKiMpiRikkJxt2OTenzjcBWX8mPM/
iF+wyUL579Pw14kPd1yxcZKWRCi7FIocepCZF+NiYKl/s6hL1Y9LOHmqPLMY/Win
5WV0C+tJ6+5m7RZdsDOH7VsjPACZtpyoIlHW7wuO9NUbQosVvEEUa/ApqnvdUhJV
UO0p7Up3vTYTDPUg2hf7TtzzCkBXW8NOjUjtYYIQdNoKkUXYmxi001LWIFQJ6B6l
JBp6MyliCppdkqvoBSIuaspXx8O5RVUGd8vl31A2NrEzGKIRpuVlbSd1cOZYcGHd
qsVLCnyvUe85/5Ft+aJJ7GTOcVUQ7hcGtdXjbPwEuJdz6+x+E0WWnwhtCjN608uk
v1y4ihW9TDGZLJfIKigUbHNB8cQ91vRop2eLM/pHpSFVjBDxe/z5iHMqdgXxJKHh
5RYMcMm1vYDgWVMlrqr10thH2eVfVws8tUFCJBiMzAiD/mwd8ZJQVQaJaMtDclOH
ockmmUtlFFz6hwsqgl+9w/QxbV7GcbKRVEhl+vExq1JKwEnC9ELVbHCG37faiX+T
D4b8Tid+OumcDk2dW8bI/nWPzO8wd0t386+p9zN4k3ft8OPyIWRBLCWYSXicqNVL
3YxzNKGqThMUMdTXbUzl85/kCv1uvfdqg7k5hIX5xq4dMk94UskSNU0GCuuZoxXz
x0H87u7mhJxdr3mEIKpwc+LxtoKAyu50nvl4d5BoRIbRJJlWhM7QTq76lla/WkgK
J5rz9tPMh9mmwJGD7wjcg3BwGQr0HZ8dwZtrd9ozThdSfc7dvIkpKejDGqPe6vxs
yymZnrnKMAXO3XwhwHa+PMAbwSttDZN6bfDFPnmW4mmiZoZpBe2YB6DnVcSwIYtM
TtBKGTenuacOdtdYmgqLDZHogOqp7avmAHppjD693qpI3lGFPFx7a6CgHUBwidVK
vW8q4HdwmHdNkbhfdJJnmmNpAcPdHjF/f8b3gsetVkHHhZdkeZ/xIlRyLNh1OW2t
qmx2g1c72oWlJFpAKIkz9ZdFS4/mBnT0Kpm0q80cYBx5YyB+F++y6RFhvuCmxqdz
Ug10OpcSIqsxT9o9+VDrUI5qdGnqlmJZSZoTvPKKB3fPwcZ/VfpCCHcpfQTLY6fJ
hzY6+YlrgtO4P63wgA/zAfdnOhf8XgtTHOuIRp3W4JmkOKocuqc/K47txiyWNfFE
HIHnoQhSJbCDLXZRLw4u14lNmjZNhodipzK8vpI2zEIaFWvi1rwJL+US1McSwJMd
ndif/pFkb8sb9IPuSnXEVzgkpHxsMHOUaO22LjOMuRJ68dhqGcM6yjrYXsLQQ1Nl
VOt/INTIvh0IX8HoSi8jFYPAJFJg1DF3jNAUhOs5wwCgc5GNDGMxF2QRcGiOBGCw
cXv84n6+36i0BsrK6yuppBnZTQ1Kum6aqcVMUtmjDHyMFO/k1k6/Cx8IMSJOo8ZS
6I9EAINO3uEWNEZY4mTSy0oGUQFeq4BE48j1ocam0NLq+Y3fC126hkdZ3K+zC1FT
9lu/tCNzt4+Ad20McK6qqRLbX2WDNgKODBo+3lkZCrHvq1+MjpYzvGfU+tAJzAnU
0yT7WprIwRAZzb06Jj1nhmvycSVJurYhLQ3cLPShCvYwg9owZIjBPLtL3DMEbJmN
r6AdI9LfA6Cy8XE4e0UH8kVNgNsrMjG4KCY/OKReH4ZWd0ifqoJbaZzIGxlPdxjF
bnAeN6GGgomFsHj5N/nEhFoLdujsuxrdWob6Tc0rYnY/oqemHhToqGIezlMIIIbz
dLHsk9kGhoULTG4TnqS9zG65+MzPMAFuG6GgopmXO4fK36Pi3/x9tYl1SuXScZE4
AQz0JXuAiCF8hIsEur5aIu7ajJ2YD2A8nzs3ijijnB1pFt+U4LMHA8PRUNsSKNTU
0e2/fBS6GDQr9rlLvoLj7Xt5SBiwzu6rNGgRrPLm1JpEvYAbDUFzD7UF7Ds4BJ/Y
/JnqY+GDPLM0ydLc7zihyxdMsQjjvBfK2xGoyo57K6WosZPd+SJ08O9qF5AJZcIl
X5scJfca6Fi670X4qf+2Pws2zD03xxqAQS1pqr/rfTlMKLKNbarc0wB6FgWVLqo1
KPodpwd8RfIiWU3YXrj5A4Y2knSZ5WJE2hzCMAfDS3jvmXGs5lDl9LND1mNNEVmZ
Qw5hR6t8jAtQlKEP87wTYMG58x+6GX90Qkk+OuC3gsuOfwzGPFzlayksp1pQFcbV
76w0gW4UDjewsApImM4fHUiRP9gsQP8GSI1ctzi9JW9uAr6MDB0QLEPI8ekDQ5YC
SBytbLhdzhUsgGyW1BEcsex9zbs4Bl4Cumh/weuGISbcC1lUfmctkyrwhkDdMIy/
KJ3rYhlS8uqWpbDjaQ4QAOmsQoeRKNZfl39C0OBNgd2N4Qkuw3zr+/I8ZAAhUGzR
5DFH7diSwCWtSlJlrwe4zqsOXmbPAMpTvEQil2fWOpSJ1ob8MS+q+T4n8Xh7SHGq
NGcL1nnRMzvEAlAbh1Bk1PPubk5fL1av4R7+u0igyhNum2IMJ51SKtMgJ79EU95D
y0QHCOxPGm9Wk+ZLu2HQc4ukNtSCZJ1HFFN7ioXuoh7y4D29o5hJ7TbtpIWeFSE5
orTECfdYPLFFyKKyG+Z8oMGHatPC93IdBmHv9g3FfnhgIhqh6kIW1bzPiGm+UgDF
cpaFvmo/XlXQF6swP7HyytcWwXjg9JS6Rl+GKTwXENyDqXaueO5i0LD7j9ICFQCI
kXtSX/W4I95t1Ak/UNPwaZrxEqnnARyHZkZpWw+TaTZuIZ8beaKri0YtanvgRhF4
NTcuZA3J5wMuZ+DlPExIYcjtXvtyiHv9kfCTIUrT5aKeVRF3O+UEPdVCJjb8BOPZ
SZfmdyrMplBB872jK04npeRz/uWFJTvzP77/TRgl0yCsGLlxL7GayStkt4ug0RB4
LUu6nVEMWe6P+JZMXN8t/RJz/BuNIC9erOYHdnAnTA9nbW6huFQWwi3vJMpaZz+Q
v9ZBRJ1NpmKs9fUxXZqdWK9qVbcp+x6d3Eqb3mJQM1eoiB5pBFFs6CU8m2jB2b/z
WeGRaQnG8G7v+byRi9m3IYlbNMgF7JcnMoGwTaBAsLV2GFnlZrexLmpDEgTWbUxJ
Qc5Fa3x56hfqZjboe2r1tfOV4QfnhdIOluuGDZe9kJDmvSLMLx9vao271iO71Xfi
lVPdbvosPuE4dDGJN+m8+6Zf2O3LAYMSMf8rB50JmfXvTAof9WXIqZ1DKRxYhnYx
0Z4UIsPX3MmDNYposQLMBkvI4nJJR5c9pYO8LXNPuHH/dUGUh0SO7oOQHGOl61HZ
lTry/AjR8RZqTAhpiXT0/GMlbsydhhO5FWr2OQCgqaABHK7+McwufX7UMlBMwgEo
KgCDs5+jSB4f/0H7Pm6o5bCedJJbXHmDpNdRVwte1X6vyal5hNnbbN9DEfBezHGK
UG6WK36jO71xlLdb3JR9Fl6Jk84vQBKd+H/GbqirC4BBLIxrMfH1nA1T/WVKeTgE
4JXP4tWoQCnEbIzgvO9FzJ6YGMMgHuZDmRm5o6p6ghEau/T3sh7wt8LWDHRMNTWY
z32wMOyCupGJZ905XJFbmIqcqg1fELqSEBsHESpIumWfWbCP2B4O/pFPWbb+tUOq
pIXn0NjAVqsmhcNK38QyHHOsSbrOOEWcl5Ke8KxUrrucnw/5/FbEI8Rqw/4GAHT7
nvHPrX4Dnzc2VZY2psnNhhnoR8iEa3FtfbO8XnPu6HJhQe+tvKyL4qXWEd7C2HHx
xJuA0qQTjygsU2Zmyaz3HJm/dZac54brqVK2iM5WzCjWtkAin2YnmODsH1VJFfrU
teixxfwzyOUu9ITZXkuerUeHeLmssl7x1NcsTO5cRTmxuHUdlzncZb1GGWKdr1do
z/ApAqvv6BiveWZD5lzfIbItaPbHH9NvtbcFfC2I7xdzGWYo1p7fBiVvaOAHE0La
QNssuFO4R2CZN6PPKzyPCWIJ1WoXLaqBBuYRJu/hevH3//pKcfUWu/37d1GDOAe6
B03nftLfBERSZluk0zZU5lxMowqPwUoA+TXbCTNEGZlCg11U8+z1YZ3P5DfTpxEw
s6HUMY2CBKXJICIKNp2s91bXWktBLjGJga5fykEm2tc37sXKmTpQLO29ktxgTFtq
mILc59etnNCyesgZEWbrzVgpFCEpOwL7CUSEXyMCkHbpwh+PQ4GoV7cX4bDe2Ktc
5Xukwq48UPfRwO/XkpmQPNvdzcEOr4Td84vESNu/aT9KGFYnG7082xoS3tChNGgq
7RcA7ikeb5pBhvTAJ5D7OgQEn5ocrxcChXNcZFgYOBQQSKGMFFfQe3SU4IglzSl0
krnBE/sDXKWaFI2NPfyAimGKiQ5wolR6dFzidNq98mMD4GYXWy6cyafsjItwu/ZG
lDbltrv4PjUzx8m2OfUQWmO8OowZ4KNk1Ca+GW0x7tghNKvIz+JV97oN9CPu5a6p
d+CkRNgwziNOxRaz9XcQu5DiwTshvYZlxJa6lBLpvD9UW7GDSeIp7uJdiqXyLApG
yNZws74STpIMmo26Z9gMkN+U4S1O8NhRShBmh7AwOkO3zmWdraxITtjNm7SuxkLl
z3SsPQ5fr29eaG3qFtgK1iuJUVeHSK+Ct83t0ve6hCUIFaN20g2s/LwHv5d6un59
DbluTGBWveYukKvI9bbpR2+xaYMjmxGucIra+bRLn1mD32Si2XVHprD+z5IGp4PV
km9Fm0Bj/3Z5R2JkL1I/QlGE5/iPSwGnxRZIeL7/qlz2czoX9SHYlXhIqYWMCwex
OKQjfKj98mlPD5F/BuPcUPMDKt7kjQfDOAwLtUdE7vi3Yoh/Ukl/ufnECZxTGXjt
9SSiMEu/og+wpntu7nrsuUaGkkFKQlHwghziayY5sozrDuTRgo+dYfZFTkktb614
obExRq3FdJTFNRMt96zhhGILKwz9vkfMtrxPyTxfi+6eiQcy12GYkzk5XNhi8vdx
OAKcTtZiRGonO8U4bCRtgc4HSw0nHt3tWkTfpCmGpyQbDr8QHxs/N17iIbRDqyzt
j4ZETc4VqAETQ4iEHD5eGEePPj4tsqWc7siKbAlaGjwwYJa6KAd7cRP9j2wav+me
XrHVz4u25unI3Ofy34xc29wrpEqYUPrQ+f6+Eo2ZMrON+3qeQdTqk4hl1JwGbBJR
/aTKghTy0JO6hk8Eqa8aKXXe+qtV8Si5Wxal0aOfSCzljR1C3EBxOnTB5eOSZuPB
YH7q/ir7Goet1/k8ro5XhuvVwOoM7ICKumAZcvtX4Zeoy9gCt5j85bQ3CksSZQHx
g35xoIY/LTYudX2tkqqq4txVAWSH7KGiGSnuGKDEyFBIUZtfeUY7fWizkj/lzz8a
6QqXb3ZwsDnh4oP5aj6iYooWdJPA09hx7riexTPEkc2CK5lOLHewK2BFsKe+oQ9g
gDjuavyKZ2rAl+oZUDwZryO/tSDFblqrMSm1+M4Sswp3qDIK7+UyeU5BAdMTtvQB
9DXceJtJMGU3jWJF1mEKO/bLC5RXjArcoq4WOMFi1VJdECXL+KIo3GsHztgIKyOK
HXnzmS8rxHkEX6SM8aVlm0bDJJBBa1pY4jTtZiBbxJDaux2vsr+NfPCT4Lx8KC7d
giBVT3Cn4QxNv5P0u0bWp0ZGbO3pbpSW62HyfuEc1g5rEEz7cebYeeQVJwf7Ahil
GE5XomE5hi7/CxJWcKtXiu3aoDqH6yNdhOta7qm6e1V/kD9VTlXOwcG6h/cAIyCj
qRDyvaALsvYc5kqq9Ona+b+xZXs2x61HDchf7LFKyE/mas6no7O04Mad7KuNWn2B
/4d3rrFpzz8wF8ZTvXmlN6e8L9Tt5BXp4KB6Zp/bZNsPZqujs/f0B3aqQp9/JbsC
R5kP7CNoTKcwbZTznCqHqJ2DQm6q+ZGSXc9UkndDRPq2DwU/fHZFpJAdM3W7zoaP
M05cpXlOUWtRoABrzr70pWZDlADoUjppRoBZZiWBDJrHjt94aTSofDDDLC63iAwe
oWGYc5Jk16XqYrsB2dc0nrC+z6Q5EzPzC+5EryMiEmap52K0fv4LwHYZPo6EvSfI
GPIN9gZIhJWJbORNdcAnUBj8hDmY9nZXaIi5p1daVMVYJPLTAsrjSAx7P6rcZVYd
XVsck6dWn93FO0OVBhjy6cac6YSxmEkQn5rPQsANuHF9lGkH6VeMrdJmdisjTjaa
+z4Xj2jngScgR9B6ni9nVXUYZxtjttT9cKuVfZNJz1kHouPiD2HDrbCxbtdCHODh
Ox3+GngsAp0bpTP7k0/61CvQYDnP1HkWrGauCkWqc9NZiIYoGRGR6kcqu5KaNpdH
ec7++M7j8cmQSoAURk0GkjjdbpI+mCnLLgYN3WBVaEHBuTYcSFJVN7y5EJnY8jyp
H2hgTkLJY1zPk8OSeZmn4T+rjX5RXjNL0RhTDIw0V7Fzr/fWNVwvhoyd66EVwUeU
yeTI/0N+2EnNdl5JZChVEi1bnV19Uyit3vJM2uwMxPn3DAf5c4wYx+lGINacE3HM
ychm4eFwTOGacqxNFwNkYaagcpHh2wZBTz+5psU56UEBhsrpBtS9A5nRAHLRX6mu
NfZd9h7W8e1I+Ru6XEpAFFP/JaJVVH6m9hntwj+fuvhkDDMbH4H/1xk0srr1S5fo
YVlGA5OXdehZ9iTZ/IMlzAhxD9/L0rkVNa4n+bN4VlYD4PXSzl76XMFjXvfqkc6d
mFqoAv+kkF2xmclxkGrrnORZxhDIT552r9vlffDos8MstmbVHhHC1elZCxNvxXk/
h1Ri3JKZHnGoYv8AFIkRqx7Op1/KwvWg+kalPcfacwv/DVGSBj+a6P1U3ak+fCbY
v6yGcs3i3GYmmLqgY5g8jmkEtArv9eeOCMqFrKpd5G97gx6fKcuhQPCqQ3JjNzMt
ggFpqKpQQnujRythGJsMGPXaj9LLt/y4Xee+ZrSfX2OIsJ/OqSzhDttBcYtHzJnc
O/Ej6SN51Fnxg2/PuPxhYvOaSP9Kup7pb8yp+XFZLwiXmkny787SMz542EqN4/wy
Q+KTky33FoAPVCHrE5YGPDLjt7p/XezajUlpdmsJz++ctOwQUJVRDpBXOtjJvAz/
7aaqbatZ5K6kH1jY3SugnhYmhxrVTHO7krOmVu+bsuoyYGn2l+L50DjESYPziFrt
76sqW8mmtGo47EHXn2UUxR+y4q78c5mi0PpC0rA0+ifBrtmf2Esa8X8nmLMmXQQ/
V5CM42k43TyFZ0GMnrIP6gunDFOgCSAO8Win4YsYNL2pEeQeQnV3OoNFekHhEVOv
+/gPvxQHjEe/Y46m2LOjDD5TZNrezEE5+T0+zIukAAu5ZbQNwyuNdWvnohlQe/UX
fd+rdcTtFWUNMPGmJABTCcVmhq9gv9wCg56AYq1d1qLuOrsHey6UbXHRzu3WyIk0
P/XDbLkEnjOfOdm1WmIWMu3Q4XlKmSvGLyjwd5tH0tgqH1DrizpDxkrLvQeQN143
lSGiqAGFLFNM4AtijeCSxENO8Fcj+DgjhL81aA3tKQ2gzhfTPMW8L8xbWDgdRGVe
dR/9wdona8JOY1ly119siiNY+sP/lpKt79xcBeWQUN2o5c4vEKPDIZc1ABG81zeS
4G4ZfTU/bmtPu6T4rF3ekWPjFKYqpsIHwOEp2JmhBqQIbBdPubcty7WdnGcG4C6N
u2HXJkPpgEwCCAmAes2lo6JH0eayDSBtnX+mre5NAxBfmCXtLajQ+6ry1zNssNrs
2kmWYatrR7oBcugxlQb0KbS7CqkS3kbGibnj2MHKkDNPVDWko2YceVLXyoQOlEDu
/GDGL5ZyLZC9Jwc5pzceD8xhiRdKUi2UetcNFMC6zAzb6n3Z5+h2FOEvHxrgteQs
hjgqITHsEKaMZmCghPFEdPmNsIqQ/ZCx3yG/VEhyUo01LAzNOC0xBFVwM3fexjKb
eHveZn40aTyoUDlhoLVDJhMkQvn7e2jovgBlaCgdqXtXGazJji5uHpoCSv72hju/
2xJGcGPHtM0Ws4E+zibUP0fZyYEkJG1CAxXEUhiMXAq9OR55d114+4XBX8+re9bD
dtiMFdsq06sssnYAZ3XCEUUOTGRVd4UIroIaETD975GjzR0EO4opBCWemhaSH52f
mXtDdZpi6xhJFVSX76hKJ+OPKSLtm+26VkGFZyd0DUy2j4rwVeEizcv3a4qrdR8z
9SYc5+NBiUBK/0CBS7fz4oE6x6VDUDaDd/a3olwZDWgikYIKIdWOZEaz3h4Vs51L
+OTt42DF0nMJTXohbjoKxcD103DKCuccXcJ2/OAqDkrlSOSrCWNLZY1O3ckxCd9t
RJFBo1yRvaefzIuaIf2RgS7EGNwKNnGlOYeeCfOITedRUZYV5WKK5sMr+kkz0e/J
C6DugZ0W+P1Yrtra/ULcR757i4zdiknHiYloE1sJvQvrlpWobIJcsMeA8sQ3Oo4W
mqvzcFRKTt4Kl1PGa7/n1/xb11mzAwTVZmnSfb9XbwId3VHGJGrypnj+2KZ6APW1
U+tYfu/p8V6zrUSdPB0VfkhqQMJpB9cbdcKX+I9a2d2h3YA3n15oxOtv7gE5tY3x
pbh6ZMWRtVwlvDbZOEC3OdWl4qBjCzh8Pb68XuLVerfWONpCCXtSDIUpnh3C6Bsj
mtjXHgg3e5UrcK/gqzh4yFDB7BXl0m24HyuoMRg1j9L/xRlSwVymy1HGeJG3u/vm
g4sH17puYk6EZgEbaQ28Ds9uQDvQa+zSvaY9dvXgbBtfDMDBq0Xc6hNFAkn0kOMO
186O/I3GYkEXzePiB+KJ/fO0g3P2V58t27WZwFl+HZJlXtVIOSdTGCI9MPBufOos
CZH5qia076uB95u6+sOOaQLL+fOGl1+30W1MCFLMPW+aVeQbOot2v03It7pLj5uh
FvrQFN/g4sYAGCVVt+Nx4YKw5UgrRFaijHttW0Vpk7Vj/N/Pco5kDL1lwWJgUBq1
Qxjr+lM92p3sA+z/A3/zktbIlYxJTQWr8lmLq4JMhjXv6JdRkVE17x84PX565it2
yHpepoXLCA8kd9g6/t4EalLOmVJD/wuU+7L0tnZjG+9IE7BwwgQx2pq/BYK631p2
V75gscjB45MdBkPo4RRlPgi6N3r611sa8/EkN/uOghhRxnaccU3S//vgbwYcLwXo
MTW6Mw7AoKFYB3yi6CvY21MV8ov/MeeJJFz1+0w8erGy+KI19h7BzcVBeFQfm54K
lA19ZTklACVPjLvgrBE/Y7cVAEC8fifmirtjP7VIfzYtmOvNJIozncH2ex9hQWdh
VEhFe22JU7Sl92WKMyBl5Nggt5w5wlujnm3f1ml8xFcHGndREvjTf8jMME5M3GYL
z19zsTNQgow+99oxmsHSN8Gn1XvpoixRcXPud+UrTYGdEuZTOwLmkv7tYBqnR+yO
g0IxZ8IcSaz7CGtQEf27ImM3LURQnkNAT0uprHTXhG/B/yAAyDj2M5FI6cphOZrF
dcts1hZ5f+5ab3en/SrahZWOqLQfphlL646vUl4zb4L07lL6mf20dRGwqQdmpPi3
iZh6VVNMbK1h8Y9tGK0eaY5Hawq+DXZ9hlfqMbnrAELIfxYZJg73KC/J78y5J2LR
OUjSbfLksKn+tFak/8/ZMq9O+QBCTIqVum6bG9Hbx2oAnONvMBZPv5+e880uki0f
vlK88UjH1BV44upNZfO3lsrkA1uHrV2fmDCP821CzymVafmvbuWa0zEQMpd5Yrwa
jADuK/RBtUEbjJouhodL6oIrKlpUaWznk6WQqj4ouTrxFMdV/+KAFdGneMV8Oy2q
9OPgCnDRealdJH8m6MIK2FojNzHkTebsAhklkzBblmREJ71f2MG9sOce5jHCu4Y1
SOJIoqDZBnsg8eoqNlzU95NhkLmuShgNcgX+xTNp+HR06Wh8LkS1N2Z69ESULcmw
RGhnCJtlVwuuYg/p+aMgMvAS9ytjng5DUH4rblDaF0tgqUx53grIubZtIUYHO6rb
+0iAEmb7pnGK9L2h1PpfDyvQBKn2xYpAyWv9iRn0SaNskxVC+jpE2MfSRH6MRvbm
xDSDz4mOshLKwpyTjAb2UY34cmvaUUbdNNCg71qYYihVNGPVytW77cNzugzrgkr5
9ceYn5lY3UMuvWkXPc7da4NVPKZSjcgOkkLVO8Cx6X/79zL6/6oSnepzvn2jL2wA
ipXSFGP6frhiyGNyqF+4GkF9KWU7LPtehnHjU6L7tmgJO0G6uH1F3F0aw8c592SR
g+WWHiz5mzNzg5yidtWGYDEMjigSVJKgmcZlwi6h+RGxwscy+lWAJGo0lO7zIm0g
+OxztcdAYV2i1bnICwg9ATj3ueG6uElys67oG2XSCoSVmisx1U7iy4gDseD+oP7g
bcHsXpsHSEAqKTACzPml8e8M407C8+a55ihkULSCSJfR3sNwu6imAYO2GEHx+HgQ
uCt0yYWRGQ7d+96xbLEm7rwtbK9FnVklLs0aXtEoCovVAppHGWT98ftJ7fupXQEA
ShZG+DZ1GnTjujYhbZB//mJhMc2z4PkyNUQ9rZQsizhT2YzEBwIe3Mb3G6L+4+4W
troE4VGcFR+R0LGzRRMShe5E3/AVYvX83BPmdTUodnFVIkiWY3ffHEVv//l3NhaI
+mmYcFAW6KL/hewjV5pMktYpz8KAhY/MvOBXAzv9TXUhmM3bGK+dvNJkTyKl+9Y5
Aud8f71cXsBLQns7W1cXGLBegtswbBKrR2HNHt0ZxVdgVL6wEI+11xw+Brr6StaQ
FQAgIjoZj1wXqJFxepMPxffPMYxyrNWmFTt82aan8ulRjXUw2u+teuvxhd6p0xHr
O0F/piriwvUe3OE6Po+NMCznRdGa1fYyZ0uI02GG20/pgUNV+4gmz4uVZ+KFxU4I
Mw73BK3TLaO3qQLvxxb+9/WyjQO0gWbYTmj31e+w95a+pTZ0WwhLDD3iwhJGmsz/
zXWVxMzAwZondmBapEIg8LEKv+oCFUYtk05zMGbdfLx/3gNqi2GU8awF0xjPOv4A
ynVzOvunVLbqqalPIe/77tcJmFOAP2DsSZ8ZXYzBlqUSAwbbMvIJ2VOgb2MwF0cN
h/vlTmSMDbAItm4KenT9x/GXRMLBBbpYrr7dZ1Q3Me/AbCFK+UJHu/ivFQIW17D7
3/upZHvziuwMMK4psm+DodokQREqJB5niFv5gBuK69phm/5CBY4mgLI6RfZbnFOD
lGr7lN9Sn1G69GDmZD0JM6jhf0EKjF/XQ876hAmfp+OU2AB2e6v3+BoM1oPZD/Gj
lscmFs/7oaKs+7np/BBdGAN9b3CuA7uVb3eiP6u+qRGw93ZFz7yiqBQp+sufnx2+
u9DecZwIrGc69dbcqZXeyUOUS93XGq0eAWFbD+RUkj1ZjEW2vD00sVrQi3EetOfm
LTflfr2Cklf8Z3ymRbA/monqEzEbOatxLkclz1gj1Gf56dKWKIR6/2YUpIA+/yjx
XmUieBCqZXxQbuwnHomMhMAQ5Vaiz+/vcbI4eYfFybkdoO8wQycJtnVjAozKMuQD
zAEeUX+yFzPu+B23VtBFCdcF7o+zVmn4YJkbYGTD+RwcoqcnWuVcLh2RRSGalDnv
yfIFLlX/QWqZeRd4581AFgAiLuKzN7hnkSbhIMwdMITgG1n+2aoIez22Gd9VWW7W
6mhF+LMzIqj+PCx/CCRW38vCEMbWV8k5K0UlNsLHMXQrwSONfX3V9m7pBrCULkCk
NL2CwvcssXInGbBMHKQD1dNVt3imUd/qWNCOIYt1zTe1UGK0cUyt6i+XqMiy3SgX
0c2TFds9fVN9NK1tztwew5JwnCDL5RZuDYbmOcVjbM6AeLhsO/deg4grVyYistM2
jglj37F6utxe44KrPqg4D04ztOsY+34Ii6PCU09VkF9gqzvn80gtyvdQMXaT4hyl
73cYHg/fwJRf9wzgPBcnW0hNzlIhQuqljqIsIEQldk9sBD5IYXlrsDH9bEaffobD
asuJJBYCK4Cu4lwwF3U/CvckUEl46BOwru2epnR+cv0jAQ3blCKKQ8kd3H0JxD+d
SxxW3U51oZ3Yv0s5qy73IoIiKL1dMEjhUBJp95lbXcza569VcOyiP29RrtsZr2V2
VU3J+Zh8Ge7v4fHxnq2rsSAHTe9wOPJPQaWMVhHz/RviwozxqogZnnuCvHBRuLyw
q7t52UoUOr5FO95AoPKn8xIqLR2DV/MZvInTxWNlUIz/U+udR3nAMxuLfm+pc9z2
6IpLPezg792SzKEYGdMrEXvOo4p7TtOTWFq1ot43XNh3f043/I1MDBuCKRtwEEoE
n8jTEnRHTcqghgw9xmOSpAGE/fA4DUvt2JipgWLXnxEd0kyaY3q9z5HhySGi53mY
qfSn/ItholLUDcrfyzckImHi0nCwgWc8gO59Sn02aUMVJdzEb5S8ZBTiDE3fmS2X
5FsBH/JxXE/qbf2unJCkLrOjeCgdTv6GZLwoXjuQkV3TY4o8LqpNXO0S9mq8mYU1
6CTKA9sMW3WAVBWZ3mTh9JKheYI44BRTiLNmkoZAspaRZJY8Mq7w/XvPy2qhzpLt
oWt88UBZSB/MvXA0dI2vkanz5LBXzIKNuyFQ7TVJMJSh9j1j1ZciK+Axli97dSnj
FhtCjAxDZl8UlNNz/hBy/3y0RyMShEFH9SNtGDhg/5nrTVXexvEWqD4QkHAIHX9G
c4+MzHgyyqd76G02S0O9rkm6FpNhO9DInlsLhqnEW2qAZ91w45ivffX7AAItUyAV
rX/AndXFSMEtclEKXYhZJB82Vud6uH8NTpP4Efu5twC0CMF7CKLFa3q/v+cFi93g
CJbHSvNhRmgX5ZmEBgbnVIsVoCI5kf++W+hZyc7XzBGZ4pm5kh7zKLXl1tUcuf7R
oR4bp7ChWiWt18d/pHnv+J5jpqJFvOVP1e/wXHH0DYlPKyuZJxQ5nYCscIHFVDcO
wCZW31Dy9iYmXLOd9S/JY/9UNkUgeEpsSmah35DOZVRWQJ4OcFxzXTBXA4dkCJpD
uHNf37QlN59GOgaSIgMiITP9W10QfJI68I12SxLrCeTLGnRyvoYSusTwEBohTE2c
IHhmcd81qjsLbGxGAVjyQVij7sSDUwqih0wsghVBJPGeFdlbQPQhxgVau0+pVEEA
W8zcbscjS+c2VzN3axiCoXTGtu6Cpp2jbZo9p533RZUHnLVh2T5pWrxP85HW1hbz
wSq0Sud7epU67yFeGKGyUVrDRn6XPToBbKWBCP4i4QmSGdb4/nTgfhx+gn3/tC33
KP+eVhLzHZJ9Bo1lnhgCTNprFh2L6gMbKIVViK/uCdVynN7Ur6mxDVlqBvlBUZT0
MlpZ4pG8xYFV+ibgGIwuJb/nOXAlKvlRwBwUqlGdjEF0ixtJk/8cL2Nu6L0FmOGl
cxvnqXHDiQGwkbewRP1ibuuKyBcxJfzJHbkqkYxct8Jekwa0pHi62ZgIP6uvC9Tz
N0Lhvec/WDpcIOJGar3Kv+TuVVhcJojoWOF6/2oVp+PxBy1mMOS6+b+Qf4qFQjNz
4FqRwoQoIZdp4Na9gac0pPhOdR6ZgWMGx7yFM7rcTMJ9Ly+8iGSbf93wwdFRSROh
7r9Uvnls3daPG6ugWadCzqfn85htW1tJVdhWnbrp1JUWCASeB2Rjr0uFRJ0a+zyx
3VdIPi8lF1xJmDDuNzV9UArf8YzJQNxmbgvWUrBfOJu2EVscRAhayKSUOeTQ3rxt
/LCR2gXgrPsdgW3Mi2alntA48mjBc28YhIJwUlNU5e4adz4/HkHlkxi5rznSrRjN
atkZ3sLYEKlKN/xVCvVlzxvWd+YWFH7MAzEy+h6xCzhEOq1v1c918Wbq8coU3SSC
q7BrB70/xBYQaJIMt4MWO09rpKLsn45wMZJhIzZSNKcEQu2N3pbeEnOR9+5dYni3
NezYAGHeIXbtbbsP4uavzUquf4D0RblSrDlqXL7idb3PpGi1eqMusFZHokYGu1LX
rye81m0pBMivz6CgJq9HXQ2a5h/IQmx9lsD5flOPXMCCH8NCOKPcaIOQnGK1LU5D
jiABADzDCyN5rgytTH1uhQ5oIdgo1yudPiJP0pJoQm3M7SzSwnvTOcBZN00rt4Yw
9Tgh+MNCz9QDjcvs+ehop9PCy689pv6DN1zFmFfrqwOyrbAghCGZ0YtKnevIXnwY
PWbgB3QhKN9qCnpPYcDTFsI8hPW7K/rskAFmI+rHV1VeHZVjoa3DNihX3dq8MNbv
NtVUUBPCPu60IB5c4IORfRUfbWI7Xa8d9j8mHvK7zTe4iqLy6Up1SPNw9aEm5uMy
wBtRAWFGl5h8QwsfA3T8JoZGPLVddx8NTI4FaiHWpDQplMHhS0PxDR4sdrSpU2TO
5WecK4eoeeqlE+nS3PaJGlGH0g4tnESabuRy+T4xtgUSIn5HMAdeG2cXtA2qctz6
CzzZzW29sb82OvQDExR9bwTly9FwaZSpfanTHtayMK2MUXazwdzhD4P36veyfmyE
Ftz2Q3KKdONIcQTsygkFWNGL9WiyYwzOAnHWpwjhNeqij8os9c5IvzHgB4bQWYb1
uplWlVMboSohohmsrY1XEXFh+VjiFce+3GG89hqXgxg0Tj887ODd6ZLEASXRQ4aH
q/PBq/EN+tltZNyq5vRyjqRXm6C9p2PRvmqf1Un22mw5tfv9iZh1OBAG15tI9WRv
8ve+Ht4+x6+dHt6v4vystsuYiC/uBgLjOk0jEE5NHLWcnuvJwKdvSC4oWxNlz+/i
dL7qo87e55qukgbPGvU17rKeVErbVie4HHfxkNj7FDd2PUQ8gOiU3+kDbkAmVebP
YPZQPvZX+ciX1c7uyx1jC6lZJDU5gpFpCqChn/VtwXOyIRi+cdvuhNTdAZryLlAN
sQ7OiZlLamOuWv8YNAjo0drVrEAX1POUm1tWN9Lx3LEZcoEcFGpImHGZ9y4PXv+M
/AqX7dqr64nnaLUMi0oXtZLTD5QxmgHXzj24PYN8Ijle9J01jO1notp84wM6rxWk
Vl1ClUBemSJvHEucRaR2Hnz4eisg4Oowbwxdtubc5vbfghWSsKr6dXj/vqclxLcH
/cx/B/3ZklWYfWQwxgcWD9EFTRwomJi7snYFkxDvymYVUdIAMwyw3BE3YfRU9nb8
ox75v2+tZo1lfSqzN8e+W9RMOR291hkJp5lb+IxmF/BXvLFK8DjQsXod7HAOh5ny
agnfPWfMqmzINVza6Iyb/1aO/KReh1TIrC/kcrDOJwrbt9pEzgdHrceTs5/nOICp
cgXEQNOyP5DBHkg969hDnN519P/2GlClBxgQ30Z4SkQA9VJbwOKqe6956JOSIuGA
sZd6bFZgeCMpctPGm6rGUj41ry5zRXoZp3WxtJqTtbz12xISNsjVZwfmfXlOPvT4
hfExSc245II19Bv/fwk6rNT9xsmU7stD4wvuZD3xBUqGz75lO5Qr1g1qfWUtH7ZF
jzSD96OZ/reQdWxsHvRVFHFkXxAyVF0hojoYrQhCXX9l9elcsehOeZ5KcF06Gq7i
zdCYOkd2gmAC6HAIElkMYvJpzImxF4kDaguZkM/XzvjwTkNNVoF5KIhMf51Iapn5
NXDfVCxavRAHuFiaDB5Vic/D2OTRvgP3Rn7MjHPgkMvzGw+wK4kGx9LA6Yz26PGt
kEY8z2Dzg/FXC91rg3WQHLc9z4fwNnE3uPH8BLsmRSMq7aDpIGdT7faxp7lvCuYf
x5oR/zN03MLE1okL14GCTrZpa2mTUGDzrsEkS5rYZkytT1nvwv1CZtDHkxCUcZXc
svde67Ak+4PlGYF/IMTiAZifG37QVmKj55iUYqc7dacfYvO/6nmN/ResU8Nw5IUx
o2JWHooQtm7FSzrXcP7VQwtMcPIZ/RtC5OgonddsUbMfYF/ZvKMNayA0dLEMpqMi
4bOD6ha4l/yDaAG0n3uXuWMJwy/SLF6UrEscS6To0D1FP/eNxPYTVed0m6chttPi
l+nC8q8LlGs43aYvTO84EI7jpflWESL6gw+AAKw9hpjxO6uOX24R7qaLZlL0pxjP
S//boen32OJw97JVnSLvd/g2jPHkQwdcq+EGSQePdOF/5I50Yv6E5oAZGT41xMiC
aH3RONMEuMJyS4d+cLqHHcTEYrNqqDI3OrKmLLigb6FrqMoEvEOFNI2R8gWDuemF
jMEr9vMQnmfHPGoNu5VVj7ew7Y32YHN1iy5ZEcp996OSjkra26cF7SAv0F0pBE38
Gxgtgy8XOh0jgLWEdD51ONwU866DrVGoVSQW9ZUsEwbuyZtp6g83BwB2qYINp3lH
Q+ZCsIjXxD3W7KvHU7cDQULE5do1gks7XWGgTSWhwxtuZNT8FvfrrY8KDDd519Nd
hLFecXGYIjOlW7+iaAOeYkncSeGiSd5wFsY1NUt1WK9Dq9xtLicfHbKTH5HC4yjy
DRGK9+MOgsGvozmZAnmnPftu2G6BEBYvxBgLMMVvfLoo+uYATPqX9p3bf1hafdmx
g47PUmBEl4s/dOUl4ANYY/ddB0IBBKs6bvvs4shGTbDWqMA/XqstNjAgHb16xY6V
OVxrdVlDWJnZOA44xjIQIWAHeq/SOnYFKhbUC98OZz0AkMXLdYQT+PXALNZsDGYn
dwNcagcc1zRxNMwWfir345LEzF6yWydBLyMO3zR0wrOa1pqaU2f/XnwQkVLrA0+w
V4RhvuiE+hF/UEDF6Tptgv2xDS0OF13DRpf8geaRJwk4e514L08iP1Vs1zML9EGr
Pn4IX9szOS1BUB+/4cJI6r4Qk7fqIfH7H61l98eFmI1AwLM2ENNdHlsBrzRHb9kj
XL3WR8zBf67G8Qsq5f3Bexobz50/RlDna7uQK5n/FKIFLOmjsurYikaU9ObQk+Bk
G5Btv33h+Tj6iS3pPtfwnTtHubgk0kopxZytWSiCemw/coELB/sPOsNfXdwCNSCo
/Y4dGaNsZyaREDjqaqTBUqqc5aZNoaia88BzOagsaQ04mbZ+8sBwRQRNTy6EKI1f
k4/l1rjp9CaSW41J1BPSZNKAEC+fGDyySfucTf8bX2/080geABXtk/qMXMnrvI+P
lFzbXUSRHYhgOQjUPSGxd0y3cUkwHUCvHw3YbSJuEKi7azzvDSyIJSOUbFz+VpWO
rmDLTYuihd9/pncnePZhyoEN4HjXGlW2PWEKPNQ/7tzosxqI8+qqyMf2mSeb+r8O
jAo9TDiSn+Shca7JVL2yqAbIr2g2auJx07Z6jcTJG17Zbh5uETdgrtQnwssDINje
pXPoBmehi5/+j4+7gAUk7mvBRNaztOLYxWsA+OX5kig7lMkk1bO9lOkhYwAWZeNW
aCQ9UWSKpRmIRvbpnB7FwiyFLeS9QdgmSvBs3KIyoE5x7+TS8s81O64p8PB93lv6
ufH52y9NZYoHHV2ErlRYx8W2mwFxOHcsTEMOVVSeTwL1pF4y6h1A7Nu3eGjcms6M
u/Pz+vjDon2QUADE1fXblvGv91IVt5IzGor5n03lEH9Z1WESqB+J/kJ/c0ZiHunN
CiRVpJzLaSrwle95UAMEwmePl5ABWcWSJSIX0XCpeekFhPho2trrdO4XKCe3eCgq
DzYgPNsGdDA92IiUmdp8ktAICT6hF46exoiPw/5RHD2beqRN+kBmOBws2YvZYSht
Lss72OzjRujPExqp+Iq/4KMf+h7UWrZTMSRzY9GvULNroJauVyy6ym0qYc1VwC3i
kVJWo0o7MwyMFvjFNxUI/GecjO0/CVApUhGidTVe36Q5XCHdGreS/+0x7Ai+q9rx
HPG6ajY4oBVOQyyk1LPwn4oLWbYsEu2HUat+2P24eaq0JzChkUnSvnAmZRyZYa9r
xxXZ1hQo9TpiIJ7FSCXugIJ/CkFJnRyCdU/sffZJ/BwnwXcg1XTXE020v74l9aRz
FzhC5QN9aJpJ46fkAeuCJCPrQ19sWj73himbkQV8UBLvy3RcwdsNFg3C9Z5AoisR
+zCm++TTl005w7P6FNaRINbyYN+YIbtG2IeyGPIg8fcWPT/U0mOBV77F3zOl7zKw
drHsf0oCzRaUeMbk19DcxZBGG0Z1SpX3qUdJeuN5/WV761WaX9XOMq2T9K43kuOH
/+2+Hxd5GUlKYzWUU33nY6bS8KKeW1O+HZ4yseVmY2KJRSpmrNHTPxCWiE6zC0qu
THHV4kQJGvafvkDZ/zW1YVPYx5+f8n4Txf3s59dXh4ECsmN/c48hxl4DbP4uNMr+
ZUeY4H4Rr5w/1v6Hl94HLtlS7VaqLDY+ye0yuoL9+ZUdfdtDA54B8tUqE/z/qWbh
p1TnwsEgRvyJgM824p/GCiSssuDSX1NZZWpfTEdvE77FwszHbHSdOLnpVP/S7len
OhFGplAmAXmpQPrvZamd3LFHBYnrVwCN5ZKJ6/74dCwDWwuJ+qXRrXjkizcs1QMZ
VxdRSqfL+s6ZVF1VyxyCR+IAARmy4TuoTXaYXfSIQlSNDXLPYKmiNvCXvZ0DeSPE
oXxJEG3LKDAZVj3pKU+EFOvP9K7y/eSsghdsPjCZFTDHg+wZxP05b39VnL4CRnXJ
XcLw096FXWk+eq59r0OvW6G8RzhKDm6XuoWi0MINDt/uNpLXvjjDTN4exU9dC3oM
xyM+uh3FT294e8yR6yWO+TV2UsaGrYBPNRf3rwDuQzYoCSm8M7W1FKv7U+fJxPfI
X8gMg82LeNvkq7StDZFqQJ/gcBEYxLQZX+hr2Yypbw47AKNN8+d1OkydWkvOmnvY
2DAWYAb+Vf8FrH+6mx7oP/+6jBIJYNF6rkkZGGSFcqD7qJi+wC/xR1M7XQqEJql2
64b2DYYD8ujjhf419A8tsJLZOTBi+HFWoy8gK9s0xcG3+cOc3NycrkeJdvHeVhjW
oqSjnICrqFsduBVrRLCxQL+9VYhVEgdWD3zU/qo+2gYBzvfWXvgD3dVzXEjqz0Fn
luaCCQzcaJQDu3pFHzQmtpznCBQ6a50fP74IbtYjd9pG7AQcxMCcaPnldRoTYTPc
xyFwhAb94EGnQoAOLc4lxb68vivtI44I6oVhr5+Aa5bLx7VKyVMM2odLHClIuO4L
GIOpry1HVsNN/FvRz8LkYenBfH+P0hhWMX+p1wTdkwWxVNxvdmIFHJ96cdktCwc0
uGYo/sihCbj+a5H+OwuASsX1fllXnlqhh2fl2RqYg48sqDgZUrZlmMdOweJOGySz
9XTAirE6K19sElMf1a9pDwYEq7V+Zd+lcF4vvKha3kZhSzoNNPvGeJrrhqwGkmN1
NTv1mZwa1Adld/h0ZTP61zCr3lOD1ehB83m7V0iiaHCx7kswJ3kNKSxQhUgCAeQi
s+S1xZ9KpHgGBTqsmRm6R/0D9QsogPLqVDLD6TVHd73QDssGfWGjpEsTGJFihjla
vVGkq/rVHRoi2a+fzDad2IPojl5PTmaQPwfu4lrSERs8cxBxxvaw8go/FQjcS91L
skXaVy/wpbHHAol+JHeZg4klEO5m5OMn/EtxjsUe5Li0TwPLAgvmGQLKgEjpOMKZ
0HkyHpT51Wox4GHbnxTVG3HmZw/25zKwqDP0rFR1IUGjN5ht7b5rEk4zMlg/TPDl
yugqtnUn9Bb5i94Iw3XZoWyMmLuaG3XlwnMnBHT2wY5RYWFgdR4/icTPy5NFNCI2
yam2BKVT3png+dsrXcdZTPD81x26Nlj6xQBoh9YzREmPC+bDZFxVNsvv8bMlj8aZ
cbbq+mvLL58ywIKtmMC9C0Usyi5yhaCQydRYO2ABM9eYfHVX2Iunc0Fh1kVvXcZf
7P2l4h3RDl3AZMT6zJPLBkzZc3ZNUejBjr1W8na3RMhlt9GHPsXsf1K29E5lu1K1
l2CFKPUifcYpnQ8KQgOke8Sx/xfXQb5ep7nrIfvd54w9sj3V+CAUyI8nTWI8ZTnw
7Vmrhpdwi+TBnunbcqCj3pmD2E1hSOxL1+TDtcT85y75b1jlpP85Kj/Z/MmeZeZ1
d6ZETlwGiSLX97kXgThlcKtEbAr5dEPAJw97R9RoUkuVIc8mhQ6yiQgS9xqYL0xH
dLr0u7fYwXJ0Lj+lUqDe8IrTMcjcD2wZGqFIweRwUFX40xg3A7drkcd3PHNgDwNu
W1Rwo0LxDcZNpGKq0kFM02MN0kjpNGpekafkWnlXDAn4vx89Ys0JPgoOuZp7K4DC
/zfCYikmNP07miaNpDYno+tA2CfHaZeD6XuL6wj0BtDW4r2GCcjkgM7JCx9OcMKT
9KJrxOHXN7daJ5MHBvIhPXRZhxMZ0AbvkfCCEiTIYggrHg7JCpEY9Qjw5V1DBDeN
nvgBoNSqCq4oXM/3WNZm0JaZbctf1mIZRe5sDSTk+1MlOoE6OzBAgGsyBop2p5sC
jXDEMxRwxMTBVwW4mZeguooxPpqA65qP77YDAJEWiisObdt1k2WI/5IYcuhOvcu6
NtfzeVRfIY9r6OuYU33EJaW3Nsy1Y6Z04iRkERcTaqCPb5iZjMymlmAKP8owQyMY
iKGsBHfFLUoL0bg27S6AdrcR9XvjNjf1udQTfciVJDCVLGjuzFJz//HEzZHXon9g
QPQMfrV7+/wYccqE9/FMWI6lcduZxDGfGIcB9dmlMXvOeg+VXztOvPZoiVgH7p6S
nMxsuq6aaX1SOKwuHkixviCD1PyGhYDvnU74D5WxqHcthBfkrxC8ti16yYJ5ftd/
COKSyyL/kaG++GDwIeNNTRIplbBjYjWk02k7mp2kfkvFznLc0CsusFQKUa+m8/r0
MwoO9Gr70B3CzPnjru73ISlZ7mh3acU1sSOMVBE9TGL7o16hLxpTUJ8r2aiQO/ID
I3SDBwzuec5WomSdUZUMYwXhNepv9q2V7tW6twUUmSXkWnsRlZQlf5p8pRrBkD+s
AbBaVgmxr/cCmt8D4mnpFvR13RAXPgQmb/KJwJnzZ/sO9l79itLkmD+a6CJu8BjF
RbeuEbgzOJtzjCJQT1ptXpNxLbXnu6GewcghaqXHa5wqNX+jT67HU9JV8Z3eYJ7F
zcMkY8gtP5vnZSGcewQn52hk/cvCpy/TJdD4SeLHVzzZTRJRrVhM+tGCGkf8Fr2a
hOQxx+e4wpPAKuBGADZziVEu7AvHlWvpYRBNeTq1AYXNPeDu7cn0bFx2qf49YRVM
pMIYSQeZPSnTt+CEZfJQYOHDUFIm40S0fd6hBLapq2I4EM54XKbF1BUT1ztgNBe7
KqN3Q4aVia4EHFDTMkdYMxoK2QCpZssZQF+XfEox1RjoNKH14y5xUZPLreD67iPe
Fd2kwSTZ/U4ni/5qL/5Btmxrz8J9LO8bnOorBLg7NHeJdeZNHM6i+whyzXBnH6ze
2vk8wM72vsJgwE8QCvTeLV1Sjn59/y7dK3KcUD7kLl2DKfMVHrRNZHg3jyF8WuTt
6qo+HdcwaF758VGRd3j3I0SwLEUEAI2B8CziVQUqnZcuvbYiF5tciiAXBM5+XeY1
HD2ziF/sSdbVSHMv7osmBsLyBuWCSZs+bQFlT42JZhCa9ii3GDucxeDDBPDVlbSr
DnzGkshtOnZ6rVIhSTO5RIPJbm1+WYbq0rsNeRTIkcNKOmK7mSkw8fzPKzEsbgfr
2vtvDp9/Iv4e84OsBaHwhFeaAEUgobm2Wf2v3EM6FEbTrGFw3l31Q2gZWCZVLb1i
NFYc5V2bXn1Yb2cAISR4P8eNq6Xt90t5cx1AJqw6VbrFnhx55PNZNUS+nxQeqBIK
Seq2uDKM4IPPjeGnG6A0O2JtAUJORMu9eZ5PlAmjYz10B70Tz9jgt3GgNQZU7r17
zgjY3L5/Ngjqil8ahuoVlSn47cGTSWcOppFWYrLsAeE+WdwWC73cMyvpN6kDDmPP
jtOXZmZXHHa/VDKhxA2RDM/YK19Cj/EBmLf6gvKoVkVviD9tF2yWDUrltV2JqNb8
9fifJrLAoYm4azn/ROK4wVVp1oJgpNOpvP20yRUNpcVNzfuvSnP5wvrkSHKyePpm
U3md6UeCyEx4IxSRD8FFkHKd20WFcyZ3KjRuDk/tw2wM9XVIFOK5TMLjNyaHT/D3
2HuWWQ7jNafoaV0Y23QiiiRmIMntviU3pB7NAyStU5qTeA48HLlNAw620hyX5C5B
U/NsdXS5T61dsuX722+gwWHa9xzVn1iIoDQvQnLAi/lPKwGogvr7hTuWUtO0L+NX
njzogzmSNWWzGUWqKVXXOZUtbT74Jw0y866IWUeD7IeXdN38CgNifII0JbKCqnTj
isHQCIc+dYSHydpreJK+v8H6f3pQvJYTz8OQanuq2VCtKeYQuNcLIJBSTxkpafiQ
epuJ5uIUG/cik2QflJe2+8OnYKXTIuaeylBXYi2teBzwRByRshRCZqhQdxsTD3oO
Hhu/DzXWlbg8+y6e9OdXyYpBTQ463XMrO1kIzgTA4pc+xryMkZseI+zOKDFHt/Mf
PBofsW5ogyS8DXZo+c/nHQ5ZTX3OKl8YTTnnRl9LaxPIR6FbNcLy0fQ8tsPpqbGO
Pjx1oiCU+WUatIVHdCxYbs5Ld2M1Wt0o0kNfqTDR/DWg9mZ/Hzzr5pXLh5XSe+Id
ynoasedz9bCr36FBJ51wQS6YacvfVFKFAxmLFcNPBr04uE5Lfxt9aIvx1ampzfZQ
zOPt+B7Za6GYjEOTB6zX4EABWV14T19FkVqypTe4NoyfPF5IfbD41ojt3bQyDuL3
chydEuc2iGX1PaWH6WAjI0th/Qb/i6DE0aEeND9u62VhTw7Vv6wtrP1hBnWK2z1k
cumrOzVUK6SwFPoI6r/bErbMV9cKoIvQZXRd7tgr9kg90yq3cPVb6/CxEhivNfi0
85AMfjqEWB3vXP5AD2dqMU+HcQV0urse+I9PkSqdG/XJsqG3zRe5VyYY/gtbQjpP
UknAz/y12R3F27v0/yM58PzX7IcBK/ypyINE3DYIcuBCvAUNjNQxq8aiAijxcRO6
RVeUhHXkwSOj/YO6FDJ0i+hNwpq9z3Vh03Zfuu8MyY04Usta+Fw27lr85bHf/QSq
j1QkYrt93Yz9hjjmH/kUSgwb6KfKA0ZPNmJAOgix/7duQdmiecy5s6eqipEA+QWj
h/ZT9qZ8wer97oAFDs0QyonmjAQp0lLF6QVnZ9mH69sW4JFoAnkMRW2CuXyMWVLT
Pa2xm7zXMOolLxYWRI4c6d1Ns7zqg6FU2KQAQ37MikAzMZZ6az1OHGSv3dZjVtYN
zwE8TvG0pbZAqyWkUeHibPnnQs34z7TUbkWA3N5o4GfafTTkenoVDHGqo6A9TDzp
GlYl2XEaBkXYU8OKoFxh5CabTQVnGHQB6AWeTI5hc9nyHYrmVIWUvy1vEYucOu8s
naVLzsZhs3jWpeDt3Zk5BTgpAUiD29BDAFEnWOakC6Aam2NNKTzAXPoRUxsKEV1l
6RLXfFqDJCvPYbMf8eRYdiYKmJO1j7IMqDk0ifnWvWlONL8z3dJtegJ/Nb+9cWd3
+aUMFptu0NHPTfto6MzuPAh9oDLXgHoO/FOQgqYQzmqBU6BjLG4WIzu2kCDP2/aB
rM6iiDfOUyx2HDMCe1CMi2MHqMfI7+e+oQmpj05Mq9tqpIRsQJN6fidZbqMleIia
+9HpemiBKCzrZ8C1CfAQcqCAOufAr0g+97PfZUVsUT6eLGnNX6gUwXVDFWNkjA7H
J0UuV+DGoqQD3yeoO5ibqe9voAzdftsWRqpbtqKN5IRu90PPHoAA2zC0V3+iJ3+L
b0r7d52ijZL4APsXf8GS6ErfXhLFeZ9L+YzK0osArOE+TQyHkGltEwrw+tGRRaY8
uxyhhHYmU49JruubQGkg0HA446yuBxf/4XmvpGSjjUqkFu2TtjlrZXSSCXO/HQGI
GQQodiNbXrrzeymjRYBAGyOKh8L8zSmBikWjUzCQ07v0pK4eIrJs6d5kFRyrgIBP
QKzjgTl+SoHer+SRj+sv5dlET6qtxkgAmWMZ0G+FqRbbEFDwt37h+yHq5jAOJ8/b
9HMi85aoIzo2muLvbHZ8sgtZBYc9a9LvAStxLAOcEnVCJTyeZVnTM5b95/+FtIIU
MUxgZJm8niXuupPKgZgCiXa/7kXJ3gYVDL+pz3DJR51gOVeG3r/7EFEzjiaj56wO
7hn4Pt0KGx4FKU+DFNF8DmhcbrF7kE8Vn1jHOUt0KVmvKSNNX0BDDWz9WSWzG7B3
v0SzMm4ahpnKxUNxPsggiSTqhlNqOj8s0u5d6p6fH3ozHxk4b3+G+VLyksknYPf4
jZ+uKthbsVfczSV7airLSHZLYh5BsDR5M8LiRuh/hdG1vLPotGKG72NYANg1um9O
drZL7HadzO0/Eo6DBfK2o/2K2EOz4yS1PVcO2xBkwlZmm2+NzbjSR2j0zQKpLLLc
5gKUz3hbfJ1y3oYmUirGq7LjccKSlp2k6Z61N/90D/VF2lgDUIcK6G7fCJFb+b+Y
zrasJSs7bNaQ5O1gaSXorIxoZs+/3xIX9f/vHRd+IydUG91GkvSWFI5Rg3P5hDpg
cbp0ykFndfrTmGZ27QqpBq/tyo658nLodiCVWm3oiDFTl62sUeVe6kLjdBTgRxNA
6ijQ0KaBHzCSLCWSr+qvvAR4qWALqdCrPZByq2BdbtXsYOpgr6W94MK3lKjR/8bb
h4wcXGdgkI812V/v/GgOQEjZBtP6mPKzmeEjlWGhsjWVM/lZTZnrkgeyEmJYBAtE
WkVo+5jd+Du0NBL2kEKuXUyDgUU6fiipt/EfqnQlQnFqodkXr/S12ho4OL0FFPf0
E2oxMGYDTcqS4/4umZex94PnykEaCeYWq0nNcIQKQFMaDVFrnldDbsv0jKH6K9KB
rPziNs6TkaQHozQtZN4Z/OI47S3iDfbalBSvFm+mzRyC8lGTbi4jxKAsua7iKd5q
woXq5Oivld3f5lBdrek22lBekf4fCAdBQzfg9PkzOL1KU3Mq7wxHXVnEPvMiCPud
GhCZm92Rixj/kNQP9ds2L8958tNNGdcfx6CueVJD8HyRThl2JqhGJQ3Z3gcNVlyZ
H2ebqoEsGkItInANf4LLibp7vJRWET3PmMFwVSgKwr7mtUXt4ThzEun+WIUpbY0p
o0qZX44XNw1E4htaUd96c06vCgJwLeG3BiAJhD3hPxv9Ko2UhFdKKInS6Yq0+OBS
5okM1lRwFVqtCNtg32OdbJ7Tga6IlBUQuPMskxmbbnfKtazRC4oDhVZ3g9ID9Uu1
g7tQ+EKNGsyUIyioKRuO0WPrsG5MCHRdjcAKbUI3Kj3ZPdotutdPxmh3QNwCuhct
YJ0VyssYACXDhzBm+L7AZgehI81DvqSbVGefAEtdaM0vDRd5ubl5/ENvTQA5+5l7
G2pqUsQHXqMgUFhdP18dzEjZVxFhhEaVzPMkj+On1Eagx7aC6CF/hl7rUWJGkr/h
4PC1qmaklvVnsUezY++HR7j9OQ1PHupw7lheq97Pbtn98FTWkDrTDu+BrMF43o5w
YskXOiQx1JZhI1nhMTdWd7Wg0ZV4DRx5o6s7GAk/yEea8ALyJ2XjWRd/EkTiKIoh
86y6WCTHoyFVcyyphqrQudg/bspZC9RQc5fmlYYQ1sithc17vw+j6Fu2398IY0OF
W2uYTcYeAwKwFaKQX4nxxkCGmV3IzPOZWWD3ZAmJX5eEqtT3qglAn3xDRXuFq2/2
8ocFNzJ67fMvjHjPJ42RVveGCbHBh20uZTI0vnvOh4s+diqbg5MaPfjtxL7IOctj
amOjgZ4TDDU9O5XWtsNqvfQUcoyuFOcrjTLd5i8td4dKMVZbi67tDtIY7/FJ1ZmE
45rKX44uetcaO3tOUw7J7HGUCwzi7h79HhG2IjMZOJmZvgwGF7/8luLf7UC5bmfA
69Q+qHeVXrdBdi1pccx/6FxaBi+zzZm0kCr4MMJ46dcTGjz9LJlKcuujGxN7gPE1
gomlbomFzBt3hKaE3Uihedj+33+YKups/ZOY5y70BXtZWzCZHq370gIsoh5w3gPH
3lCN8PPyNa/fBwmerhGT1za4U4fmbYG9YxlzpI2KhoFBs4HaJWYhO/WlQ6CaDSbf
VQVKvTYZsSQ/enV/6znaYjrZgJjb7XV6CUcEbVIqnT+2kMOck7qLKYoY5mYuW04X
7p81cBtEQDNRekkuIWg50PCbrDqzsdoTOi9/nsNreCbqxE9wFNSgMWZau/VLIMgD
WPWTANqg66lmcPCPiP+xWeK8F85vzNL7gDi9E48cuv2svan0+GTDgcy25qQaMou7
3NzY0yigiS6aOA/4p5FgJWUMkm8RwCHOiMHdxoPcpfBqKoqDGfAwpvMDrQxvcXbm
6261qX0/tno4HTGaRgTQiNUY3BtuHmBVoCK6u0TLixJnUsgx9bRYkfxc0neTThnN
Vb9i8FiqtSR6PG+6k+h1eKbMRgQlB4OjVAXNKcT38zzudiRYYVM9pGuX6aAygPIV
qpjLA/cVaOHxfM88t947iYRgnWoC/8AW01QTDpniKTMYY38Pjvj9MP8DRNfsGk3W
drbYZPyd9QiR420BIKEAWXby6G6CHMikKfQ2JX5YLjs9MjA5HYjwzqw8+sdbkmMI
jw4acwgoyNjH3+MRe23lglZOudPDjxsygvqGBEQUaO6BKfol64JpSwmMVxjQiSdY
FOJ0bGKEh0OfONs5uFTwgFPuqpKamxU4L8pWvH1q2k/G4AAdq9qLdKBHqKSW55Rt
JnQN4D6Vq6VK78SVsPNalFQMw6In85XR7sy6rRC6aSRCiziYHQDE8CAvVlb4WaNa
eeqWsLHhzVPd5b0IJcHfwvSdGyTduKAMO7S7QUymnpyL7t7tegSHhK1w0U6NtUh9
0tR5jReSsVqZXZWGoT2qZz5O3yabJP0d9MF4qvtps9i5h04LqrHli5TC9Zo5BcaZ
ZoGA7q966FPS99wjogOHzY/mkeKhDmt2B5JlGwlZdz7+pH930Rm9xUhKNlNGxUrx
/aQPI5mKovES2idHMOi1/0Uj3wWMCxJ4/vXSq2ciFDyvc8PL4en62CbZuukjWSgl
WcyT9+oo3CPF1bU6O1cfq7JVi7FzWq7NLBLW209y4YTDsRZJYuRC5vJioKBHI+SR
tlq/4UDyDZta/fjj8CwJiNCyqKCPDwDOKfBTGYRadw/zU9g+/TyHhd6y6A6RUoA9
PYRNLc0fzy9lVZFiVjjJvRrbFnpJzYdVTaLO9lnslhMSNNI7JZI1b+OZgS8L8Ck+
NxtnZJP1+O9KnRZMowVCfQFiEAXecjvyK1sSBHLr+eMOIcRDSak3nSRHp15+e9qm
vOiMfrKtx1ndNlNcCfMK+vunbIkcvFjL44DpebnV0oSUkjNizeY1TQ070lEPwHR6
tTndtyMFUS+wJD+wAk4EevP5LI6foR/ci6FbXmms+sF+vwC4u5hf9b7KrAcUggmY
ADOK1XlQzaFLh3odhQbnvCdgPk9BX1O7fAfAfpsWX/fA/uff0z0p6tx1p17VVnyi
pBivvBekfrrVFtnCpPxvl3U0B4z543erkqO5ke7JWFYckEDxs78vLUDhN43gPbLg
z+0DrAr18nBkcKkn6IW5IqDPUvf51MhfA4Mys9XAk+r+dKCO5QkX+Z9RmS1Y5AwU
tJJh4VPRneD9eYpJQx+Ld6sRGPVqKZB2GTD1Y3yh3rvFA7q49X4oHJo712N6oRR0
Kqw+eUQveEhVSV5rIJISUTNOIUmWUhv9LtnohNd/RGklWQONnO04kKC9Dd74L/m+
/WufGVUcy8xXEl4PBSGg/qbi7uAEMWx0cMcysOLz+QvnttlaLvHVFSmrWVZ7gw1K
oe0SG9fGVoWALskbeohTfhycEmlgAbplYk9Ge+j5cNbBoycEr6MZVsXGiJAs0suQ
P7oibn1+/DPI+X5xpQhxtlPi25KBb+SPy7tED3mdNP0Bv/WU12XFCzNxWYw1RZEw
+7rmqrTO/5R1WvVWmPB11oo0com3MQ7LZLpgY0irIHtRpSogpgf3Br+OEshlmnlO
X1VdJT5ZtbNcVULGsUihLK3L4pRXng/QHDUk0+QcW16S58ANpHm2YXx8tD2ECqVF
Xkn6fjBUIGk5+DZS0N/oTBQuRODeEpS7/txlnX7t0eeAwjJbrFSlz54fuJ2xsmul
l4HnIuf99dC8jOeMzQgnfnj4GrRAr9UOQKhfWwSTAtH6Lzrp16WYaxbCfbS9VUBv
o1zJvUbLhgNXMgto5OEbLOmnhWrkClUUMl+M9vfuJkh6627/n92R065UQYZX8yzb
tB3qooY2W93Vuvo7IJvoRQOxAirSF5drHoMerl90QFO6+3aOixDjTfU1p/P55VvI
IZ5wgCCoG2y7h9CTV70dvGM0JZmk3o77z25elpI2aUpG5BKxiJ/EbxRantKfKlz1
BXxYc7IeLjEPPAP5dnFEb/wT8YUvIYCiUZoRCUoL+jK5O9F6ukerYF3lzkX0SZhz
Oq0Tr1/L6AXNb9GBvAbGAKzSsjd5AN42Gi2+BHjCno5i55Q8kZTUI0mCFLLND//t
Sy6LbUmjMobucApQfIlvOfd0549EJXSsL6Ng7RWvUvDN6Vxzcq1uVX6XFDpY3JP9
nwTwOCKY9UoxeOZFVsbROkdXAlFvkZ7xfOH/iy2REqPi7kkWdWRMedmQMyTCNU2t
FcPG1W5U5teP9g5EXbiXRq1Rs+kixgKp14v0hOpyFWFuBABk84EXStAjWqHRFAqm
FUJ9fM6a6X5P88kQBN54ASb3XVhI1tl248sJw333SGsl/GAzYcbNp3Ru22dq3244
Sno6lgp4BNaHk0joiKjyjwyBY9RXIeENJh2suTYuqF2UGy4JAsMVPWrjDpKYhoxn
ieNmZJ0S4K36Mo8juleZnS/79Kdw0Ra57+3xZOu2Mv/Fq+WvLZXbuuelsTcO46jP
ZKEMdFxkDCbsVKu5UrcvZuk0ExbGV7BYdQPOGUQqSJnSJkmSSNPpcuhVW5LA+0eh
hjz5hkgvcbTvieZ19UqRw1PUSP/FLo8BSWIyn1PO+2KlauEU98baEgxhWYLnuFiq
FSfW5uHMsKM0B4NmI0YdZsgUq8lxFBUnFI6GQ8ol8WO35zBQ0b66TxUzGNbcA2aM
i0OZABnSpXhuBSWcjgeDvKt38gV96aMQpGaLT84s143/mm33RgIOdPcB6aLRngKv
JluVqnZAKZdeB2g7KS8VSiYJHnqFASymHf7Rque2qOcQj3ZcEdi5o/3KxJzuMzKJ
k5xZRSZBVaBxEeAwcs2jXrdXbO7ip2QE6g3gcyXaWZKuoVzqeiHdDr6d1rfAlElU
STidW2LlTdFWqruzcidM6CKVTsHSNLQ0E+/6j1jJ5BgzOngYZWG+h1nC6XgNTA0V
4L6n7fxH4WIq3dSSB32dJNStdgplWA10mtK1IY42RJ+kQyPWa2MfMPgAVZKmi+sY
IVVfD2dSKjnSCu2v0QPpcoKPsZEbrslcD9Gkg6/v4CML9bVVSPZaE6OxuZiZCbTE
NAH4wwtnkfw4VPOkUiXWkwFEqX0LYTcnf3QTWqMtW8++6d5Ys4J4vz6b7clFUHzW
Ur7T1jgPHRbY/H2Ag1A1TpOLeaD7G0QuFffbNNR6V0Ybaw0l4nvAgkjafrOghgQA
ZifP7N0yalOx2Rvf0J1bqW3ebhtiz2+6g+AXRWMXFyxvVfElq0+dKNyeYrYYLEeQ
7ek2CVykDncbekg8El4BvZiCEwsoIYD6RvE3XNHbc3byXQ67GgvlgXsZdfujhO7y
S5cr50JQaTSdGnto8YJORJjnv9rHD7yyxUj/9EwgLx57/aOes1vnjyqFqbZex5LK
NULNBuVCu56zcU0nN85RzHg/mL49ASk5eijcCZWyzuAChWp70owtvmti1nWH881k
1p2Gv6ke4/vNJ5lLiLWJ6S2XGNvP5Nj4mTmJXdk5BrDMaaC5JXgRknIR4txJKOAs
Y89foVIVyCvLohuust5subNmSSlUgobilxiXWVLcFLfNcKsafr49rakK3hSjy6a/
aaH0SNd8OkXbSHM285ec1MLaMHMkqkL3NlsOvpCrCLtOrCCAEc7BSyXzyxwVD8AZ
9P4sV6mHc8i/uWTFNziK7Q/hwGdsAY4+3FYJaGtv6FJeoR2GrHc293TDxVcZAC4u
yzA79TOb36ppRLulhYu989TgAMZxvvhWcwdWrkNMHuUll587A9LvMFKUWMYqp1vx
92qSDMykjZ2RXnmXzAxd8bslhifLM5YqwR4xxYEJKiQfXJzPuW4rqKE66UIpgqGn
t7oTSb8dD0Kbx5HlSYYxMMth9SIZu/Sl3ZFJ7wPogwIzGAhpugb2npJMEP7KgnlF
LpVirKo4564mSZYBrz4Nu8m7k05mhS1bAJVxMI38h9q9UqM49cyPnqlxQRwrzUVO
lShCsErPJvuHOpiCFKYAYC8buSY8Dp7lf6rt/IBK066m5UxUvYyfPpFi6s8ARo6+
nhOUlDZZVPz0TTVXWNIDPd1PnRKk9y1OtwDaqQimk9qRKBs8vo0buEtvX8GC6XT7
qoA1kLdjNXTwZ7uFbm+rxmGAqSd2Wi3tV4gPrGLaXejK7Cd1i2YqmND1Kd0u9bbf
kqNv/Q+IUxYHusR8om+/HHC7zoyxTkRy1/0V6MtvyJUOonO081cUIx4vOO5rbIoC
s6j7KfxwgjTsD/08UtPiBJ9oP3vaP79+75h0wUHY2qpX1YwvssrSqGzO9UmVb07a
VaAC+ycW51n+IG7qMe5lHCkljPYHFgyc0sLt+gIfaShDucPS3FG5LAQN0SsQAF9V
C2z36aUeN854hvKydho0iWcUMQhIg/JDydhPkm4/gwzq32+hOHaq/h4bJAHgaKoS
XJKyPfKoQC3U0nrGUO3XEgSbSQgtHcowYixMYJqN/bB9KbUCvn8YteiXUL+WFWUT
vuYEdUurYbFUEoBwOza4J3QpXZ5mgqIBV0Qh+OK3T3tIMmPaWqN4f5+8kGtwm8QP
bmf3UpZMArAMWAtsk/57ndJsPJYwWd0qPJCX9IsMYILWcZneeb/qfq/YOeP/WPUY
P91eO2n/I6oPt0aMX//b3531hMDWXV2ayJJXpOXGB8m/4VdDdlx1LO/tLLqqg7TZ
/Up7NdGfWN/S+3dAZgsg0Ohd69DwnojpbasuJAc52TmTLj+Ei7l+9wiQLFzAz5sT
iSZ6IZSCxHNe1QNe7buE7QBd3hagC0WOG+D8CByM0ef5wg2tXW/W4VeMH7W3vq6g
XiZuR70SYKUWDBADoR306lZGvbP+jwgkyfogikV5PkTJTXXXyeIYKoI1uDe3pqgm
B9ZUcknWO+pEul48TAr587OydsC+/31+pm4/mBXYpg9Su6QLtO+Yzrom0C4B11U7
xouEISKmmlWrqdWYXYqNoc8srKXz+jFW0OVmAplzYEHqUkk3LPDXQu2vOgPGL6++
ztI4PVJrOSrMqZPbhOh1x/9KESYC/trB1qdcvym9kY6ZBSyeFl2Rh50IhQo9R+B5
HA9oagHHRM+jL5ezn4WZppOEA0xJwTM0bVW7D9+sI1+5lfUQtydXkq7fc0ChU0ZA
rDFoJAVTGzyrt8TOElEaNM9q47eQteIYpF6h3ed5P3Sd++cEz62dCHE64nTes5Hk
YVQNADvznwRonuy8k5gHTns8yRght5FTVbKtVCl0WPT3IItUBrNd5pUlHOhZi6qH
1/ZmMeP5UPMnVYBMK5XpIiSyJMF+fA4qR2KbfEO83lR+aaY0v4Fs1ZDqXBDwbZ65
7ADjy2jYixYxXH3OsEfTdnmmriqVo8jO2eTYL1YRMS+kM3IWMmiaFz/ZdZ6IB0yM
Yydt2hWHvO4pyiwnpivvhtSbk2saAUy+E7SL6xqepJYjtoYTfgq3+Y3AjBIDlJ7M
oX9zHPPuSVnMnYSXmZbZu2Sl3swKMNYQ1bXD3mdZ9W+KQJletPN096Qjut9IGcHy
Ysr5xDna4lK7U7t7V/i90p7gv4QvPcsvMODtO/R5doY+XeCf7++tErLFtrrvcz3O
D75QW43K9IBXMTLiKK/iwihPbe3NdQbB+LHAmy4BAJFiqqOLiQJ1c8qLAPyMjFqR
id5MQMnHv9XaaFcta9Qht7zny8bb3+30zsHpEgUz+ViD1ryxwZY+Ima2sLnYabrE
hoAHHYVA3cxdPWN6fYkbRRRNoDF7oMVqCRp+ggd2sj9gLIqBDBLNrwn63NeBvUV7
Z6EiTukDZDBBfcstf4mNqFzWLdSBSftQ6TT6J3asTb9VboCMoVn8e91AvR00NHqd
cEuq91yS3BNJBJe3/VqCPMl/Wp69DKEamWtx574ir75VFBIovKOeG9Wi9vd/kHMG
iGpbCTZrPA086VJxuwyX1i179MDVIPuTHxPE3bBB0ANMgv0mn5uHsjQ2eUxvvm4U
4dY72q4nLRkORqSVLrALZvTkI7hiL2Gta07rpnUbvKySEqA2F1AoQrx07CF1Iiq0
eJF4W4BMh15A3vLOZGlBSrdXx4sWB/1dpurTU9V5IEOkKem55PYoKFBFsUfvxYCN
CUUw0s1582D8+EOI1wz7DavrDwmd/bGLk5xRdI/x5rHcZd5rNcsfJ1F/tw1ayjvL
s4EV635kSmq6obC8EmNklyeEUfJlrIg0UpptMzRhlU3EiACa1EFRQTLu2nmkETio
ZC+4JXm1p3364AhNCe+5A7AFbqqANpPcOa7x2qUUirwsL4wbZY3DZDjoPZ4VhSRo
npbxWa07b0xdha+gVeEt+Ck6zQ5SWTdgOHNNTuaNlksz9fuVgE3U8WJkck2CfcX/
BC7Ji6WaSo5dA4JOJkdp12zycHzdvsTZlSJ+wI3hl/tQRUYczlsEQ3U2TvIRu7Oj
6Ernvn7mzanPPT5hsvPoKebE5H8Tc/2KeOIvMuOVL/IHUEdV0bVnzULNOS49HUW4
ngIKxLVx8UiFQ7wzHyTMByBcdLS2PSxTd0kluhxSYzemXpdGG1zZNg4blEXBITAA
sJbYH+xXysBIv+4R4/RYOopbKUl+h8y2Fu/SYJR24AgfiHH1EgaMeM3ey6pS1lt8
RErx/11AXHDO3oWgyMqidFqKQ/n2lzpfnxFeWEBCfxg0Ty/dHTUWoM7iCWZX7XVo
7/0beZG0aepyqWDggLB6u/bYqt6cFaF9jjm3BKihs5qIisUEbbpLRZXrmGRpzyrV
sEjoHPOZqrkoeQ/h9lyaj+eMfjkeduNfl2qLbI+VjGg2dfii152SHwGQk1AyT5Wn
S3AppLzTJHYqOJGpzNFxh5MVLglXYsmk8cl6KmaX2zaHbsuGfQiR0JdRGuOtPZ4J
5cgR4/L9yyf1qiulu1xfvBdniHd1T8Hiqe96ey6+Wdu0EluCzIZc3rezkP/g8WMw
AVNzRWQ9IV6sw7HCgwaLffYkexJv2zxp3EGI1oO5VwKCE1R5A/a+17Bb1vRs1m62
NH0W2KY6YaZPF2biFUQsFZqyWvka/nmx/CGGlVXH74dbtBdIy5YcVmhkucrf9ZJ2
nu2ONNpFzX7HeJdCh7y6AlrqIucjuq8LBJ+KKoRRh3468UKqPD1PzeuuRdglGlvD
i3m0jbyHtDeo3advlSRW056SZhmHjaUdJ7zAiIaKnybgnWgInkj9N4X9Z6WgnQgC
RZaEg+2dIyIl9n+MdM9zAUbQapd0UNcIL5B7ODMmIp+0YzOMg8DkmUGSILJjpOQW
jyXBJm5XmLEOleRnDbn28n2xDYab4R/d+LMR9LEkF3j9fNiswsHrttfWXuT+GfTa
vn5DV0CJE0N//xSoqxJowTgQ3b+UQ1bWd6hQXJcizIKtI6KcOpKRM8lI11HmhFrq
XLOabS25TNENKeKn1MpGARbNcqBN04d5wFT/ZrHul1piEq/fKpmzxOtL31Uwd8Gw
As7DtX6crUnH9zeCYvq1F+AbIQ5EkvJ0AXplNzRf8/J9yjuZmYPNDo8233w36kTS
ZigSCZE0SpUxGOmYm0vCtNomJJZiTm+lUr7juMhCbPyWx0RpHSpAqgxd0dMsqWkz
YrD++HUzHphtPxIKCuZAHUStXz7X9mnQ2j0SwQ1+CPPIhaZn4lFzIcHJytg/q+tq
67XpGeYgvO1Ov2+5bwLWhv2VKMxDz/AnC2A/3b/ptJdUCRjHNG2c9GbcGDi5KIXn
bz1MHUuBThPc0ZrfEKqG6artiSXAvk2aps3zdxtFdjnlQ2yVEfcyHFg1Wr7B0/Dy
tSR16hCn3yXwPTyx/VUPzv/ARXfNgBbsl8MVjsafrbTsMPpMOA/Ze1m/GSMBIAJt
Np30GNyWsPkjaPIqjhBQpp86HgicPngokJ5SJOzCHg36DysrhnC25elXHyR+Gwqd
ekogL0Ebb2nI2FcBIEi1b+2MBZATJkdTEw2MdunjCQ+o9nkV/Z7lCSQTZvkSpe91
gwWSwQXmLBTLl+GLANGtjEMSXO+uGYatK2ntzN1EAtSWlfXZb2LnQ3DOxhKoXI3J
1YXQ74BVMgDX5t5bOp3lyPHpaqmyAssVqngvrE8Ofui9JsMdcvos80k5Nwh++fWl
Tmd/iErOiBT08+f8JOb+RYUHpNE5WCz1g1R/rjYT7Y1Fh52hsISKfBRnGb0L3WbG
vUQFmMxZsZRKybbJDrx6Fpr0lzrsX3H9eI6rB7/8n4ags9My9eaRYhn2phXd82m4
nUCFuba35AcGgnjh1D5EHQ3Xj8MbfjITujv/LYEmWK57Orq/Jm3/T3qmAj9g+PJ1
SWF/GTp7FAuWSQt0X2vHQ4ryeBYxLjHdftS96szHl5fbL1Hw0fDYz6dSsmAKqx5J
7/NF9SRBFcGlRv/LPKWxGqR0+Mdn+GmYffimQYIQyRKpznYEk/T16EmpmUMiWtPX
NvsJ8MH8Bm8Z4dL3xcKN9os15/r+Lc0iwK0fnwoNJxctI+xqCWDTtmvuBDzV+f+i
S+TIIWVIKLZrdBBCkikdHeNCco3DE7GhDntcEW5pnKMbpQ11n9ZqzQWVfrZWF7UJ
9aLNx0gLqey+fSPfQ6puRa8Kzvng3XqMuP+6aUg0MnDvep3XrfwKVwjUp5oWNqzl
59xx3MTC+yHCqkW+jg5zg544t7x+cqxNznVmMtfM7+Nyvg4959uPltG0/gRBi0rd
qWfmxkP/ajQrPv/dATOD/vOwSHGSUhZzgr96WlSCk+ejPy9hGT49xVGsJmZv3f1R
sJnmXKYK8hEeGZYVVQyq8GczC7osdD5CQzEaJp7t1xhu1eei7iTR16VyOcL0OTGc
W7g1BQUC0rWxWzbfVmmIsWOaAmaoIHlIC5jXnLIM5k5uQ44y1iBzUyEf7BvpSUa3
1OObk6/a+L9aE8HF2OoaOR84UYPdp89qn9OmYcFfPw31I2mjFk8Ygl8KMIt/D43y
gNTLyX4rdc6M5MKm2UiVprqGqhc86YR2J10K37qRSV693UWbT6ALIHj87elOQVbD
KNeOHpnddwPrOm4X4aI15CDfqz4xLHno7DsnTvHtfR3gPr7478GTNhd39ncG9qMQ
e2mOA4r/tMeT/B6g62x2Mz55LuuiaWF0jh6pZzjAnt1VCkEAvCqPnlZkl0D7AC5L
N+pg/i6OOJga7KNurg1Si8R2NczbSKioUiQtbVLIs9CqJT4pZpX3d2GFcQ+aN2v6
6fycvX6QrzDWScJx2NvU5L+AtWcdT2clWOgPzw9G2kizf5z8skWTXiycUWnp2heg
A9ss/uSyyoaJCw5Ot87L4xo6IcMbb+YvoYLKEqDBlek40KkAt5nL6T0mZwOOWnNS
zMnKrAbgnFGAdYTtpxVP4i5ICt9FVoQ+69d4JWb7Ty+DQxA1w706w48vzjT84Mjj
FCw2o9zufyzD1LLERAjLYM6dSBxE9phKKM9fLVO9E37V/ivAzcXbOiEcFd6/jddD
+DdlCBSI7FmTS2cdF/5dDHxkgnHSV8hSGkwFptf/xS9Gk2JvyTRVKh4nv9FyzaSA
q7YsOe/7S5labAJYhUcj8vA+/iWid+jq48zTWctEaRWbUoGxpU4oT2PtSQR9Uefj
U322GSxLEfKY90h94OtOLXA3sLgfhIf9s/KdQB+vic/MG5Q/toT0Bym9E1gka3OR
YzEz89mTC+7eTi4B8oyC658lZ06NCG/v5RgP1dUUYf3FriCHxgsdhXQXjls/BUVy
s+ak//He3p2s76KmoDmHD0EYXNbTdopo+vOadP7l1Nqk8UC9Bfx+ag3GNeTGD+Tr
cOubtQcXBV6CHU0pwPKyBCNqw7Iebe4mb2EfHou8btk1YCiENjCxRoTBR73QV+Hb
Y+LM/iB3nGN7u8oQ60M4VK0T8ae0reUcU+0loPG8C4d3N7u1vX7II3zPmUiMDZ3U
t+HJ3zfzWIhXa5MBEf9y3TmVBQtDaTddj2nANGHUaAdvt9pXvUSCPOa1oP44rYAJ
OdNN7bw5H2J+Q0CzlLAhPK0ekYUHW/EfLGhlB2Bf4Vld3OYopWQQMRIR5BhSIV1x
y5LNxRI8JAXkZv4G7oaHmz6WjVgFDzFIzJClX2TkYeH+CLUD60XpHNIYp2uqRgO/
bnJ2sB6K4+0yGCbLiKz99YXpyd+fqYOBNF6UfDkO0iSzPXqAeFwkZs6ClE4CbhuU
rzfeHi5hY/gN22vkvFj7SLhVl7Y9/ICDZNKGwOyG3z1n7La8purrtdsTg0nvfNhk
AESav6wecRblhIpdt/9+oYvcRQLugS7mFywvICRvSfrZC3x3cUdnyvDD+Tmdkhua
PG8n0ErBYQYWWj5iXmVNlyeOmPFPxc28hxoOxdhfQD3LZL8in3+gLFGMJMoYh6KL
ymDSX081QPc9kcz3EbwFz0yV8lLD+6zPBrTuqSdqNNdO3lUr6HpitLi6PkfnU8yR
ZQQ5ZDhPwkyQ+d2+2+bwceRY1U0LwSWrAN6JVQug65P1sYlv+htScI4n7mpU0Tc+
nktd1NvF/0DDOcytjQIRuysAov2y/45aiLWZLsKaAATIMnBu3d1+SOR1oL+/xxGb
3O0PMQxF7JVKSAyuii83amqG0RFVc4QpwkslhGSTLzVtpxVs3vDvf9RuFZphgsr4
hSU5vBnAUW0FJbZPg7epmq3x9LHENPNwHQg28ez0MrV4azwE1/lwB01zJfUDy5FT
y4SoSN1ApL5y3sL1FDGENLDktsX6nUnc/VuWulBgmAgvk+DYmT8xzQrUh/5vnJ1b
i9IJaBw6DSfhOQoeXWLCYczaxfP01KkonIU6UtsP43ShqemLSPPiv1/SWk322IAo
zRmVfYVAPrnTjZmUoMUxRaPYO2ktlblpZ92d9tSP4iktQ94qKFolfWbMFiALEhKx
pyAIMEbbFyIj0cDsOVe5MBvsDRhKqyckgcyeq+EwW/SpJ5QKqprtpQGCd1UUPB6Y
XrtgPq1f2urW6OZcZpRZ9t9XILVmUZbMvDW2fMQW9Qt3QLS4VoBu2rVreSJnuRIf
ceiwEsTLNGX2BlJriTFCLESuhwrVutqX/BL0LTyEA4QZYvi4HznR1sUDEXXSXIQj
+6iq2AfiicCl17RkWvAdQMD3aJQ6QJvy1Pmy7nMi3XxQAy+5QarrgVuogihv7L5C
6sJ9BIbTDheifXpfgrXwODHOq34z+deC0eryCOsLGNjyc8jpmZ1ZRlmXhwPnr/ja
QzQojUTsAxOaunue4+N0ZhKMw/sekzZiCoNt3YybOVB/8o8OFPhAbsvs+6pRw1dA
WpZchk0Zh5vb/RcjLMJ/TJdU8AnV7QsKTDrkrVFhR4U+yzQTB+3Mx1m0qKyAZXes
ulzW09YY2diZhd0yFzt9BAM8Tljzwlv5HJXrJFzJxnCPWb37Xjp2kJeX/X+s7LuF
6tkZ5TQcMQkxbEz0uSU4XZ+XE9w9GxUGHpXD5WDmGejf85qHsgS5NQwBAFCPqTe/
7K5Pb114gQuzjJHUaIYo07vuCaivUYTQwjFycDuK31tRa072sW7cIboGJE2riKKV
eAzZF6UiThOStmVFqTqI9yH3xK3qSDZ/6vHCMwZGP4VBjd2Kju9Z3UHedc2gDRRl
RJcuKP2uWvxsAFbjhYXviBi1xYKuX8+ADRwZFj4k9kTu+czsS9p6l2my9Xog8+Sl
gxftdXSDl6KyjAWwXeLPLHuH3nUu6BFMc+bsiV83AzTqQW90kqvUJhKq3klv2ALn
i1HD3iJMlnJOsNIEmQ5ZWZBwyPN8/kBHb97yg7+pbJ92Yy11WPuAE8MMRk045e/C
OrF1zZOsTYLQvkdxXxIRlP///UYaQsYTaZ2BvIPbnYiqePmT27IrvgYYc5e/Bi8r
P+aXjV1ZOk0gkwmptQh2Z6J/6W7jgNrdo8//YPZ66lCJYoHo4k0zsairVaxvfXzs
IrN/AhpsjxEnDlLG13SPn7tAXTf+rJLHaHF6ymkjSMT9m8m2rOJfV2tQYyO3hDM2
mcyQgCEWoxn5yF2A3eWks4PBDY/loPYtuztm3+SrM1pdYepuCHJq51ZZ1uEWPcmq
S2EjxpknurLrIAh5/65OSlY5ZKG7m5+QSOS2VlgCuL3eb2de5zeGexBi22/wCE1L
+iRNGuE5aGTmemiGtl9T8+PWrcTwILaM3YJktKDLfGD+P44k6DnhkW7O9HWLt4q1
YyI4iC47+hW7xMjBHV0Oo5bKlGHwMrBl0JysHUEAjIqXqqyW5VYEtpsa2ZR8q7JT
mORRCk11ijwHE7X5Wczk/lGMuXHz1D7AdVY6xwjwLEIL7rp8R8ErM7BSJB1tTDnR
eLdNR7GMs6Zh2Si+WQNw5TDLVREH2byRG5CXUem1VTpVowsjGdeQGD8QsjILyZeX
3Dr9C+EpSwnDWMCGXhyQNV645l3iH0nxUpCnaUZqbX+idcEkcT4CD4ipx7RjErhS
lMBhXtbm+accDhzG+cFKTxqbGFtIWUGB2dP5JyNCY05ZL2Y2kmidMOa8mfTau5og
No2cCOALqYEXvljGPrYBVFe4V68z5urZnA35yEAkU6C+tBCCA2/g11pp738Y8DVX
IwXakYwVet88eh9C0LTZmKIWuDey9mdE1nWXXA8IMTWwo/yVd+JYB66Im8NJJpvw
QAI2EgzlTpZmzsrTkbwQi+BJD2riyVrHHeLt8RSptJr9X1Ywhh/KEqM6QWB8VyuR
jj0wyDNrodCWRgoixVn6+K5f2OAfmlf5hAO5It/iAhjtt1jhhbV1fPekOe806jBx
9UMYy6gTwLldEhtzruLnlu6An793KgNag9t7xxuDXs3FpFxbUmvByS2EtFfJG26O
d8lPxdqtpEDTWnwtnPzVvCyIF3jD0TXpMHWEZGzdONcv+JJg6szueyc/tLPoZywG
coUyA66D5Y3ifSaMSUMGawIvuxRnebal66wTXqRuhviQ7IVPqPkMFQEm6Un/3M4P
qCQapeXR9CmE7g6gFYpvRJDzfOuXD2TVXS4IhxR5q7kBDG07Kan1Yicq7sH4STvf
NvUqN5gjf71xhnXeTgGH5HICABeWF5JhqW3lyD4SQQ/qMcT3tSgT9a+1BdWH3r6T
lbkSEBgmNhg6oJxdYBiu7MRSHesRkeXZXmq6/8opw+o0LMbOCJhKPDW+y4cxCkUR
6vOqL4628HqxKkjPYjuuWYfgmDzNOwIcLLI75+H+pIxQcdm2L3t0fKCI0MKEOUyF
XGTpkz67A8bZh6iQgWYY0ChjpWJX2pw07nj1RurQCLiKFcfVheP1ixoxLx5+w+2F
aZVJmcoJ1CVWiCoOUvJt1Ji/pC1Ef+h6c2ZSi7PRhrksjvnrJ2XaiZATm3O4Hu0K
W5oLj1wMRO+QsKS7WNhn24dntmh+QW+2etoKzwSc0pxH8+aCIaC8+2B2G9UBmzTd
MWdffWFBgaERty6s3pfonkncSyrbA5bRla26MIxYov4UNu6RXUZqx31tIdn6y/M5
hUPbBRXi2G1zy8GPsd4385NS0RyHvfan8AbQTMJdaUxP3uYV05tbf/gETXKSXnZp
97FnvBo6V+kLPVt3KBVZR/dgIrgk/WY9Pq+AVtYZs+wSfr+tIo66dCWWj7gvoWlo
AJIppookb0HfU9qWKzW9tyzovvqLiFOHkY8ZdmzfWd0a8NZMOcSz8ZnK4LghqyZ9
n8D8YqMOSH3W/JjIDezYWf0j+4pH/YFqLZr/NsMoQPwNh2VweRstsInDhhNUCOyd
uymRi2KZJVYuyPgc3wqKfe6nbHahYM8dxpcJSWM3RLhlUVALovmYhIuFl8ehLFxj
RXy3IXRMbiJ2zs4pzeE4QQhx1VMIWf+dQmSWF/xbvU5DMf6r7/mSPg/YzBfwN2oK
lxQIfvR129G+zTzTVN2PRrx3LgfAIOzW6zqIKEoffnuVXCSvtlBB9ukV1oP70frt
InCxsKzvmYThHVRMqhaMqs2U+rWbIfqf2Pfi5oaii/rO1uYh1c8wcRvGpJsJvYLX
pTMwDwYQeTgSrpR+oI0qMIO5O0CV6eY4RAKFQX1KuS8iItF2RrmLpi7l4hz6UZva
d8xOFV0iAn7ILE01mQGq7e0vvZItzhxE1s5uLSDfir3mRaW1pLBM9SxFPG7lBrSP
PF+qh9TUUEihaE5w1xmIz4X+BmBpmSARJjKiHlyEnBh8xZy1RrePN1ioCe3H4SjX
KwG8mYfgVJDfEN/kxnS7dO3lTg1gJSLBb5WF0aCc/Qte0rgzf9y2WIC15lr8b1t2
ChcWmouM5LhhqiEArHt1KNTN+ghr2XKOQdgkGHeJMFGvvUzs9hj+3D6n9lVZsiCF
XIn0D2UZ7eJ7ISDwzeYy+ONUUFHeqQ6ugg3/9vTkaK7iR+Q3OZp7kjqc0gD7bHhq
pnBiSp8IgHz7aUl/qyXtSCN+fjkqQtm5yHWnJBsi0FjM9NLeWEKBNdUNvRiGLRVQ
qJPi4VYlz4Vaa7N6PniAD1q4gXEOLxlkeuWAA/zfiG3o9MUhPjAW6cLuy8M32mRP
3yslpYeS98JtYq0I3ke/IMg5/2c5QDlGCh65G5gyP633fGWI/3MHHeQi3EXsSHXc
Sd8xRhpn2+2CauPbSv7Ex2Bam/F+IOtK+IuEWN8lPiNawDsWb/FMupbvCb8ZyCzu
m4c/EXeDHbtf/xWc1t+tt/q2bQlpof/iHWvtDxvN9pgQ5g08HVIsyIVxTp+d0rPA
diBxAnhEg56u3gVePtiPujIrilALIrsXWJmo7L5qweYsCu+rr8sz1okLGKmFklIz
96QDqz8rBw7Xy/o9hmqsQZjPK6+J0QsK917iaw4MJ8rkhAQDpC9ZHELB0qUZFRUi
PSuK4HUCBALkb8B1CVTuxRd4Eunbruc0FMrCT+eMWb6NtSdFDFD/gcXPbjN5RVmh
T4lEEnRqYEhwiwR2pZug1AIlDRZkKbDpZfLA1utWXqmWkbvbejodwVOzU2eigGtd
HTyt91HcdRTNO72D94mTareGklrcH+T7WNgHrYzwFYWA7v1wvprAoSL4PlSt5La0
DFOrhYA6+ZmjSgPo3c9O6tYyAX6/UTWqZQqXU6usLAqn5FZsdkoSxo7BmEFfnXmJ
djxlAP4qr/+oqCKzl2Hu5YuUaarF1c1GWyWWiOZVZCLjwOaEkmMTR0LSSraDkVuY
pvOtk7tT1QnAEstTeViHz9A7Fv9QZz9e8SWI0DRPDz+J/8g9fpLLnr+yqzwYXZwl
uJVFMVrvn73wZ1FDcXvuO9kAFzvUQggOpM/871uPntBVzN9dQRwUtO1taKZDPCg2
3n61n9epDB29vvZlnOoR5kF5ykyjsZOfC6vYjLq1fkDkqCy8bWnEna42lhrNjen0
sfKqf7RePXEo4+F/3TTfPGFVS5IVfQv/9qCsretMrI9Yhh0r5gCwjajtn7c+0wtK
WTqhMdnRZa/ArB2FiASFk0MDG7AitiV+Mvc3WtyoV3WZIltlUXz3hh53tzGL16vS
oBH/CAZM3PO0+PTp1+ULTSqHCn84CgARsQmLURobUPQOxHjZvSOmkI4qhzDYQfj7
h9FAtvb9CkVbwP6lhcAIItfOV/7+KWj/iYx6Q+PpQ/FQP9Z+O7klW+uGD9aprYE0
AoVyklrndCG+XsMhzsQcI2CixEqzlyONmJvk0EW8pqFqopxecXDRPwEzYpb8qzzv
Kmfz7qAqoGrHfjJj+qQ5xB6LanDAbLnGpFbtH2WxsW3frFz2nBazxSMyWHSmkpkN
yigJHBvjpn5m/lR/92OCEjXrMeOfeS7al4PSga7ffH5EkfgVF04QUMB+MWSHwwUT
ifi9G72yui9bKNcJ2kAT5JtKHMIo+MJegAzQWHyb4WfRj0plMtsHXAzZvPQm8bKN
5NessV9OnttZmXFl2owZ6uCJVyPFIXEpxKhecigvX5JQLdnhx9+45H2hQr3Hf5X5
i7xwlKD5uA315u76cgGMg7oy6baPcasiwk+0t8CWaEWQi55+iD3C0YpimTPitr3+
SMlnHpphW2ikJ/F05O5II3s6fEWMS1NehxVFkycb+x1gMyeSguGvhpGOJUdSL9O0
/fIBv/wHxS/YZU+dbiA+JqumtjEC9ymXQmIke5MPufR+EMhzZ3WHyFXZxeV+Flx2
xryu37GqAs2ABjGJa3LMhbfGUXrrZkTPBhir0NrwvIoJoQxG2eyFCsyRhJ32qno0
ho0OMubu2GS1UhA+pzmKU2ZMVz6YJdlHAdZiGHREvgJmCpAO/QhuXNOXjPzHV6fr
AV6+yBI515tBLzYVmRqqfFaCekkb8RvtDtIMBge/KcUZ7/MJ+PCNwpF84tvowwjA
qdMrKVdT3veV8d4MlUZSzzXVsCg1t8JzdVl0sDaZaX5zyletQ6Rizbrz3j2DUy7L
7JWFNHb7WHOYW9RuDCxwDJB+53xyWkC66El+0u2WJJv2ytvUGOOcpFeCDEEGelkt
3Tiy7bAIDxCQhZOOVN3oUrhWCxMCD1aZlaQToLUARYUEPnTIBTogsQ7879wLPjs/
HXW3rUOL2KRvWHZOWQO3w17HP9WC5yDcUt7v40X/4QuARYtCE0dL4ln0zrFkynm7
MKhNfhlggtQz8ycFk6T2fWYYf05MZ8M0iiKFebtKxEnzr1sWTyAOxY9PtduyEtVS
kkHsqljiVfohrjtL+qWMvurY5Z2R5zuam9S/5IrfXcyeJFeLm6qPTd6uuLq59txZ
MEF3LJ098wbFqorJBaMNXNBS/zPwWD13LXU0OGc8tbGscmEJno18NZAIm3Yw8yDi
wf9UrKAUk37k1InIfd3uXEeNT8rVvF3wvyRVY7/WnHulYo6NNhtgOHCbvSiIdU0/
AZnWH/uV1lfgHsrWNTlsPfzNjLR9BtHKTE9vXFbrQdr3T8QRIqZlcb8CLs82Vge6
nVTw/Egl+rDPrF9uJN+qu3qvcvvXkox3lifdeYpE/ImfnBtYkxduVPrF/tYu96Ts
VJmp8wh9rlANSG2cEFe2JqyjzqrxMJ4PLv8qN9c2uwfSduUmPOhS6VJUl3KAdmwL
Ehv9f0KHW6RWaaGc3WigDKIaJRgqRABkAYfWs6AQLDJBQp+qtqElxVIUB56Nf4iC
d6zFP1/Ht3+wfyURktrblc4mEKpwlqMKO/p68DqLWZRwRx2U84leg87KUvg6tXAm
AvuYxApNZGQULeAvdJiuGMaQabikQ3cdlLBCWodtqPCwRB1LBuujrDHiFY/gaajn
OcDemsrd2uq6DTXyqj4GBTqEg4BdU1Rk8H3FjDIkzxyFjMTCe+6lth52fSirowgA
1HVDpHA9uzydu57oMRNBzIc/fXYPQ5RDNOwQdk2TuzV7uHFrCM0++G5iXHc0T6UO
a7dx7w3kTPTgK6pIlcd3HgtbQoPx47ZE5zg2tfBqluhCKjZqZKMJmDfUxJRDINrg
rTn+z3ayz3lNFCmKMBJygMOkIfVoouLokkgwHTYs+xQKC7ba34xCjO1ycsq3xv6A
IS54Tqz9FnuqPYBZJo2mhzjZJMTayCfFKkHgla0osa+0jFstpKQf9fgqJYVYWTBD
d3LhKtVx3Emp+hA8AKFChnH21GbiWK/Jumwcsmh3GErv2wFUxkG5+b1FjPYIHo3i
Zg4ijOb3PqkPNONkxbo7mob3TxqKqwRglk/hhmm+X+1s7uxLBhu6IWyqcqoBJggw
FaEGKjlMGz1CdKj4sRTRrq+u84rqfMotd35BfKoUjuTgYEwyoBoV/Mdhv4hXcuE2
yCL9ttkUFlEEHVYKOQ8/7qymEy+CH3kocoL6TIkrP5fsBuglYRd/P3UxqVoJKRwJ
V762c+cPCKT000mQ5urtRfdVnD3wt28QIkN7NYSWOwHQgmgRUFYViZoJ5DkrherG
UbmgVJDRd3F9QLNBMcmzEgZ0Fhn5xU+W5/XonBeeQyEyC5Rx3GYKfsxAeDLalMfK
E0vE/r7rzzY0nO8ILA1Tu8w6lc+YesUbQDJhZfMeTmR8+cQB90MIY/Tvd4nYBvTF
SwaAfRBxTO0AcbsF2Qq89mO15gvpLZgW3ReXHueJ7KXvLcJ0enyyGDH6H2Td3aKw
gob+/3bzJ/EfK5QBKQt9nBOLhc0uER/GpYHkFJhP8rpxkFvX0j/bNNJlBYPQ03ac
0Nd6IfwY9ict25sFhEt1inNd46vxyhdVDoHpQqcAGY2U9jPYLqzMN5d8f02gznv5
kefm1S7DBDISE0n1pGr3T1fWDxWH8Mqxrg/IebPf918iA24TtjlKM8cb+v2uCpfj
VCimjMiEmlinAvTZs/czi3TjvRoEMNxK408eOIvhC89Px5N9KWWmmPJZChhOigpx
bXsrxLSpiWlTNO+2ghZ3rrqkOr+uydJfuRbOoUpd+wgMrvaZgdtdsWBtrs2escF2
+fBYjNouVLfkwm95Jrbp6Dj9bHu4Ob/eXJlXfF0O5/AJrHkge7BOf9n0SZxQFvk6
HFgNziXPwKCMXBbslwL74seAwBg0gTzr/GQM1JMjRhbxGILb92qtvafgA4ZaupNs
CfU8Gi8lt7vVcvZNnMxcwCRlSuijZqN/S8bdj4qygXjfO+J2K1/H1h0gpgwTG/sh
MQbbARmNWyd/89akeaJgKAab1YaXPkrzWAboiY0Y5snbun5tS9iXTU4rtmoHf5vb
ihaqQ4vztKRxuLpeAub0RDP9iOogkH9dxQD7qFVH85y+kVeMH7ZkeW5fVf1VtK11
P6RmeAyKf7NqCKyU3IH/wI2bCcQLeCyDxLUWyZLswjd+ld72vY75a4RkCPCLlS/a
abFkA7uUU4su7YDMqjghCd9n/oQySpyZenR9bY8NDFh2XaDLBz8MJpQvByXDxC+V
kAh08h7XpkSsIQrzXDk9mYrcDT32tUMmOzQDVvTwuHRMKaRTFuh74CUSb5CeoL4n
jo4IZfM39Dzx/7S/GNfoew67Gq0tz9dMyXlJ74rJHcyEc6TrJUC2Bj30aJS2DwDK
0mC8VKxwV8mt2tb3VxfLvCAA9YDTAFxHYew0eiz0hS7aVfxMDTlyDd1nwZCmcD8z
0vlFJ1mWN/eMMpWXwXieiqaJkDNKCX9u+IWLq6gyBFFmrWgazQ3Oxs1UJSx0SJWw
xrhw8saWNuvv2jraB+2AefPev8iYT8yGvizN7n86lzWTg/x3xxYm9m1kOUAPzsMX
V0gecWtIdiBFLKXEJHqNss8VgwhEqfTX5Myw6ES3f1NTAYGfeeD9brwa96vVPHQJ
hRRu+KW/6aNrC9roxI24LsaXzpJh+bggiBpjotqAI9UbM+fGPFQ4NDl7gacCKrb2
JJJF+jtJCtQSBK/1mDPw5AkCP8wiSJRdkSrj2CJMohtMbZOeaYL6+l4dYna7r2WI
CRPHkHVQmU+D4867wkbv9i5Dm1Q34rdmx/zoiUp0mL+NvVC+ZSJpeeyz8PvdepCi
n7bGUtGck6cAFFeB3nShsRqelSPsZzU1DrzfMLCo79MrexrpwupDBQzNcJK1BmUu
vc2jC0883EGsvfD0ZQWM298ngSzsYyw5c3C+fFt95X6X/V5Tl++mIsXiuQTGvqZJ
2HMUgn6bJv7+8cxF1rv+fWCeRsa4O4QbeoGjTJuFxyx57YFGvEi7Exx9NI4bHS+q
7tkAE1LKDzV/KI2XEmFIQxMlZ6J8mgIYg5gNlEy0mFCyzvDJ6U1rXM+VpLWfpD4h
oVlHl4WarvwBHqCbHU2sJV2o42ON/EQTbnXRvlzzlmbJVT2s6hwgfQK4KRbi2aSy
tAJKjDdRgj6dUjPMq/YLtZIcvsro459RXV/tAuAyEe0MKlydHdxyqpuHSESQxMp/
yv6OQcq8tla31zhNITXUKTEo/IggW5R5VThNIwCwEJ6UOtVKfjpg8XnA4HrdO3C+
9b1STfox2HratLBQzDp70OLn+GftAGaYpSJcYvUTb/rfWiLP95TWA2jlog/gHUyt
2zOftGseYT54AFt6QXg/73PYMoup91YVnLqhqTZy7yR6V80wu6OI5/7JYHB97Zaf
LDlwPEVe5ndMmo2pgeoHMYEN0gIf647fGm2TCD5gaE+ZNtt/vcou8rAl4+buOc8Z
5QeReNksIXC43no/an4Ot/FtGRAyZWiF6Eduu7WxlS/VYHbGX4AE+k7yD3SC7r++
0n6WAS9Qw/X24URHs17tIjxgb3RzObREV7OdhJvSohistfxh7phZH8vYcs5HnLzb
XNt4SCfYuoOyuPgkSXWqlJPn0SIhd1hwyqj3AXI9QVdDSRiwMHh8PNIJFgzUAXex
MMW5b6TU7HZLr2BvtYT6Sh3uJ4XzxG2Ta4cXBnrU8eZI3QFOPeeYvUEQPzcm5BkL
pi50VKJvHvDoapmzKLcuY8eOZOG+U1F61jZ+1HHQ/aiJl+HshjQ8JCZYJo9fplka
rSe76pfusv/UBe92OVFAHo7LO+op9MhNU+9QnML7qxpoFbCwL2wl+WmGhrM+OeoA
FngE8/IIYQqBBsaamHG3ssHzVIL1zOKh55pcgzamMyb1B1rRTpA0Tfxa53vdHWjx
p70HWJCMWZvFS7NiVlCsUTYgIeJvGuAwKXiw4MEpiwL+ug5lrgrZ6bFuR8wzYNDl
QouaXlzEuKX/lORw1gBlaiPMKKZuQ1Qj3NM3tYq70RosEzDh2vTU3rbDEbcqvaXz
Q8UriSqfi1znQoOkmD46b+YUUa/YLFRNbOM/UocYSQSdF59ttjn6+i0/Xn3ghGj4
2Ity77Dlyp/4PIS+vYlr9rPk/eg/EUPLd5cjVbWggtxsP304NOxeW9h8OJGryqHX
I1QFZz32e68+ARIsA+ElriZl1nuXZ+YCE0KdjvXwBCIrdYtoboGliOCXeMiZZc0/
gRd27A9okmAJhJuDLNIr6A03Fq1zQAhcEiwxkUlJSjv3hdGfBw6WG0++odv+1NMn
jKYOyOK70YaADfrqoU24EiVYPGBRJlMrrY6o2nBoBifG+gkj4/j5zXlQgPzQcLfs
sOckKQinzBIdXS0/oee9xSP6EcuvZD2qm5yYjtBW7EPoVja2gYO4AF6v4qEsQAgq
ITCZL0VwuRhtOiAf0ykyxbHTGTjIdyvCG3r3tmhROczeWuxOvU7637zvanjgaBg6
tdQETB163ACQVciq7bwN8aKKm8RnzHedcnM10DHs4N9FwAzAwDpSgSgllzS7PLJ7
lb5RpvVMLDLrK/tWU0r7nOSbPBZcR2ABvWNkHA2p5LFTE537f4RowJPimRP8TJsw
uKL5J0yHyGZv/b151Ukp66P0av7VVLqAKmQo8ZVTwzNrsaSQfHk8eBLA1wLjSqsd
LawrsjpGfz82x/8THPOMsbjlP5ggHlbShz5tF7JKcE1mo/Yzoh/YMw91TmFEGWLg
VwhiwHmDDyJhhRrZnXjGF521L5qkFyE8b34yZ7lgnSDOdiFLPNdvbrEoNx4T4BBA
JR6NVS4umszAnUTMKJKC+w/Gt9JWULagDeoXSnjzDEuX3HLn13cm+ctdINaCYBg5
vuylzXE4AbndEYLqyc9aZLX8SqiFVzWrALbsJuxPm3sGuZ6Nu8iRoMYSSX+5j4ar
JRWJvPxWXhFso5npmiV4fzWGv7SWf9L6lEd7V00rJkTPk/rTg0wfXXD4fJFcCo/C
NL0fPnbuRARArXeWEPWuiEgpnheNH5dBiRIz4qcnsn2zawh+SOfqkffwYiW4zoTK
erPYePAbudRHlq0A1suKN676R7M6s9LZG+wa8nG5mbhGP0mZcjpSEkWnxllGPF3m
1s8gj9Il6T1i510IiprCYs0T9uPVP0oJtKd8IPe55YCsSS3qgyQa8kKzpZVUaOoj
l2ILfnbtH9h5eKL946YAjyx1RcPF+Zf3z++YS+ZrU5QrjaHIQbP+0N3ArvFSWBa4
XS/+YmEN7L3gXx01d8LpBSLZVkRwjg9/JG3WURu72hrcOIzjf8zkuR6yulYJEJHX
gsNpwa2T0R4tBz6RoOcc7q4HZpXMdrnnj2RFUHyuxCJlBj4kVVuvHXkEMzzJDvQ1
9vKj9p6e0kBQ7VPtoA1PDMK/LodhZeO4sAo9xfGts2jDXIypmokXSfMfwGDxsNz0
oi7jafOyOQRvFuykGG2Yxn+CcgHMQ2+XXmQJ55NRWFD9hmAkX+G6qGSF+wt9P3Xc
UUCTqDGXTn6VBVaNsTbicwjpnIOGq35zTjXeBSQQh2gvBoSNPg6yN52XmmthFVsE
0+u+rmHmtRwRzUcdOe7DLRa6kku9wmPgqYwUZxDHdDi8SY08gJM32XXy0DRjHKQX
07mTB6NvSxfoKKdgqUfj6wvBx4nZ/Wi6Y/B7Jg30UWDR8xWXyEfq+ZqmKgW9g4H9
rUf2dhJCXHo9KMxuN9iebO21jxjsBwOC9N32/eFDNepRyF9WHQG3r/mtix92flLN
hkO3Ol9de/jTa/MacQvFZhHloBJVVjcAXF85+abaNpuOtmcvDInigx96wGv4pEZD
xMbn1VI+fjE0kWwa44DqZ3I3w1IqJvMBWMzxPiesZAEN2dvpcepObI/EwoIU5HBo
OdTJxHl1gOO2YPU1MuivOLVcdtPBp4NLI48bgn9rj8K98DTuJyojX/dL/CZqbKwd
1iqYgNZoOVskMT7p1zaBZdbJrQGfwwTzgG2s8slcvbDx2/DKZnDh09iu0lPlFO7m
C2PIi6JDE6eJpwdv0XaYLgJ9/PdqYLcfr9QJFQVxxqxSvVFcfSnn8SHqvOGwUky8
t/Q1qYJWMGwQt42PZNakffimxPNldWckDojWeWVmoKiQW28JAiuhBJBBwrjlNDLY
g0BR12b3lQ/Eo4elllU1nRA9wH5+dCOB39u/gv7ZKOnjaz3Zb8e6AyRvYdwlIus0
267TIXRr5R8Vj/gqkLRKGSzQXaZDbb2R399DlnEwR4vKNJ2dfR4feOu//lSqvT/r
T2WqZ/Ta3O1jfpppmrr0Q+XHRKqvCkJy3AzM70PmZjBg5zoJUpIt3NK0mb6txABY
c59/2F3z/0Yfvyhr9/CnN+g1ITOStgyXBbdpC/dq56xcWhU5xdaEfz2g40QqoaZ7
SyJUeGBtp1FGYz15UAOUWOgWEi0hYCxztIoGHxJf1eMe4ssGCAoQv1EK9U+WIwLb
LgBatq7sGDAclqKLeZTN2HVJS4Sa43lCBoGw/UNTWaLcYIm/GP4ALL3wfEfGVwzH
6umgFqFUx/OosdLsTtI7xA4TsYfKR4T01p9I9LHCDKLUus05FY9kGGDJSjunnTvr
Qqs0zf5csJMeN89RW4M6GrcBDG1FGXZW1oFv0nyC5PAThXzzXa/vELmjvmbOv2bv
GYaR2YWk9R32M05Kg9orf2KIqjSloupe5TXBKxLS6lo1BmajrOp6le1mPOkhMoCZ
ZJaMUcRiqsq4l97mFZCfn7SXHGnwWf+3BSVYomOFRGcii0vEWLL9XTwQeT5NFQXi
yohWrpBtm5zZTDtK2xHg4lVirk2oSqsCxh+kai8vWYFJgh/q1OvJrk0dkZ60kweW
GdwgTe88gb2WCAq3rLOxsU6IxXQT/NjvwBUjUT55fSTef5vT02KLJ0nE5Z1ycIqJ
OM3u+QRY3hVNCvgQX8V9goynU6KZPcFeyFFlrdp8kx8ChGtPVBmvLbaa8aXsRUbs
IRvRmCDspRafY07cZfn0keli6JMb0J5j1h259/axT1m66zFOlacmNP2LCmLHUWlk
bW3mzKUIGo3BLWGUT8QbjPirnlnMQvLFRqKUO8UmdvbNOeCcBqZzrASmGyP2v5ks
uiOWwiKeIiD/Yh5sWN5+vBIL35ducb4unynQyex78LJ6qqxrpIyEPmuUS/psI8UK
du4Jcy8kkDW8HbdZxrEOrwdOe2FuZkW7Vh0KjskAu+B8xwSdc1CrIccrgdiTtYtE
1hJfVB2rorVkz09c8qZ4iKXme4JoXnLSRhH68BB3XsyZNyaHHEz0vbLKMLEnbqV0
bwdyFuaPoOnPCRKOMuOyJIc4uE/GO7nAex9ukyMLE8LD/1uHCzV8Rw9Iy59pEcoq
O8l3JaUG3lS5SQIKtrXol45d5VqoL2jIJ9Md3h7fZjZNu5XNAkaGbNJ368qfAc6L
XwAbLQrgB1l1IHNBFiYjOMaff60qJC14g8+1dkvhsjEokVV16wHaIwHpkv8PLR+l
evF2GvjqhWJIfqLfSuWZhIl2R9yMDIR0/8Q4VTUaKIGev6oXRMxVZzuWn9ytLXxo
Bw2QLwxHoHchGEJB23BH9lar+MRB0BNRxZuae92hLpJJ9oRT8bMKe1aIYZC8aJqF
qTTwZuWe9J2DHQ10gsQG5WYdtrygejG5Ugos5d8rUx9VSdGqwsspZ01LSL37V8OT
AgMxjHSLcqm526OTiU2ARKUhMW4C52IBwAvP7Vgo8t8c5CtoSkbwCs827UOPXpAo
rH7+Y25PKAlq5ZEBIoxJvUEpXjUwktctNpTOkrC86iXiJYdw0f23TLt0yJgiftSh
oFw2ocMQuJZyAL/0uRdjb76z2VSQK1Q2a6vWgGYIt2W92Bo6aeKP0unwPMZYORGN
qaaH/IJoQiKt6NofU5iuyoXbhgq/5ah9XivliTXJZsJA6xRdjMH0rE4W4Vhc/8rF
NBwTora9rASYtk6uNwedscT0SBOIjrepZOgVncM6CnUMLvZtkeGtAv8TdZeXlIvY
Ql3laMWrLb5mvOG+LWwtG8FSJwn2/MP5fXnHKFtm4q3lHLLiDAAZIuwmOV3WhHsy
2U/fn9yhAeI2ecMOJYiE58F1NX7T7vQGkgMGzLP4ETjXV81RxxCd1sCIQEQWQmCH
WqHtKA2q5FjZQUO/a4ClW5eAfajbS1ohKTQ5sB6WBFRuBMRWfGcCY3wbM6DdB5dk
ndizqfPCGO02HprDTK1JlztZWk+UMMWr7ikwJ7FTBXvFztU+TK1F3WWrh5h73EKW
ypF2rHR6NcP6N2wRsBfmKi7q/FHfg2OYk7v9Ubao9FiTbjusJTTaavr7JzpAXWRX
C0flJudZRzfSwNhoGXzYA28eYgt01QLkc1Q1H1EQiRRoxiPddPkE4nW8AvxM+hbv
RVcaLHy4x8BbpNC15By29vtnKuvro63ydzKBVf77/g/rLsUjXsV4NDSNe3pOz2SC
G/NNX42WyvO2nrJAkIHvsEw9p4XBHdirEOFaEg2Nxs0RozXubNm7DXHPYuQre/La
orUybHsKzBFQ4h+us6rCXrqWzYh0CFBpyzTh2yg4m3jS0aQZx4+xWMeEgpxFUQSS
HnaWABs0JZodhdu8ni/hQyz7t/dDPDaD4dtGbrqzOqSzH1HlZFNwuPbD/RQjXp31
euiBiXDX1XJ+QjscIj3zfU5l1lB4aQ74Iwn4/haldIE6L23VFgDBDtsiBhODQD88
dsLq8t2jpm9msAS5CEjzHnA/2mecXv5Z88Y4xwhM3ltIzdCd6vvCixp/4DSCVihM
NFcuz2z9kQb5A1m7kHPf1AWtq0yphfblWXwm/gX+m7I3f3pCkEEbtKbeIdh1Hudx
E86GxqyjVEQXQZ4SmvmrZQuUWaJn4psAebkFTDn0PK9GPWgWsG3x4cKdr1N7p6zu
ltJB1UXiil7qg9tG1dJ6ePIitNbmQ6ksIhnZHmig76c2TCp4L3GJzIbj+C8QDyam
YWNSb7VOiAY1FHmOf4gaxN9iY3wTOTahJ3tStJmSHNR9i5WIOTEkNYaDrC11gFgb
U4BWZw6kew2KLaNbvCW6tV/KA+1GYhz/eEJAcGO3GqkaevWgL3fukWcbTH/AnPoW
OIQHVUQ1/4Pa4tmGOeSCTTAK6fb+ajVa6CBhzQHczdxUJxytOBU9jcp4amaltqNo
bnUxmXJYW4D8eq5Tfv/Kxb2bIfXJSJqe50L/ul6DlpMgBX3V971NDuTw/kg6ytEX
dSDi4MEXWfyYWEiIUPBfxNfKlhJOjwVdPjOj42vpQHSECN+OCPk7Giph7nA05MLY
QZga4XHjkd9etQxPThy9m/ef4VSRbplCRboo2iQDf6UPoVPOpgVGP6+6C1Rk66AW
4BgeIwEGcKWBL1SUZmmL0LJ65TeiLDHzzX5AtvX2b2fbJudulqKOGlDOupnE6ceQ
OZmuPR3fWmsglkbQTTz0LBCGhi0bhIZvrZQP6UW0wIFUoZtGKqjriGRm1uP63ub1
jb3sFQH7713XTvqf3Up9oOjRhdt3X/ZjjcmdNHF9ZcXQTBwTryVhN67rt4EveaRT
6sjlSUryK0K/Q9VwQRu9M6ELI1l5WLC78jmzz5PdOIcl4AUQvnWL007wlbPHKFEZ
5ot8VlAQX0nHNah7v0ilyZIDEL/MR1Z5DsOu8/+wXOgJ9cfy0honQoUV9RyMT83L
m58mDbeMsuZwHPu5sOrQp1wIFz/PRTcrg/uSFa8k4CoYYuHKYc5lVcHpeMXvwhXx
PNgpsbZbc2hC88VMcITOioklqCDxLB/HC68dfYOgahLArrWfB3Xli41km2ZbtYhS
R1h9XAu67XnDNYYNdFBC2pyP4ig2Aa3YNf7BPwJgrHNmBWIqbPeKAnmvKmPsMFiR
DEhLWaquLf7pnKsg1qmRcQRGtdp15BCXlj5q+uOo/tcm/6jujWDnUHzQCVDnbqNg
ViMFybi/yXfXu6TOlV45oOGKFk2db14Py+weyczmlskny7jwhvQIkqKv8L6RIYOs
0Auf5exb/XjUb2NsmSL4ZtFKyITXi9N4/KhdfIptKJ6iJ+c9yxE0RjHC2Fk8uty7
VyLOvNV6DY+hRDmmt1i7II+W8DtZ3iTOl4RG3ofj4WjGM8dnynDWfn2/5Jx4PdpM
rWt2eVBWU+AEjaKApveboL/L3y2kHF1KbI5Hfju8hCp1w3iIQyitJISDincYZSs7
z/NEhMWzmgny92/aMkEg1hzk4zxfCAmQGGoJ+OjH89mxYBDnStDvXXOsFsWaW8Ey
+YJJ/E1WcGXim4WTkHsuZ92YLnn2NTHa3hzx3zKNbK5zcWXTcLJwO2Npbx7L827C
6BymdX8nA5NHqifnGaXXOlBy+2Gs8v+bdVX/X9TonQWdbg+g/2QEheSmcXylIAzF
83Jilod6ROP8mlZjb+5/jLuQ56SSr6464X7AA9kIOSR+U0IGV4sQMl407YSaWJWo
ZbFSFOj0S9gQ0bSNEjESd3SvyHAS323UwJQy6HYAix8OL8/RCKAaDt2eFojUubz8
n9rzURDmP9+7HZN3Hh0HMMCBANTLdhHOXP6EYrmfxb9MIO11liWdhVmsZDS+OJW9
iNZO48PAEEuFYyDR0Q0X0aWjtajTBW78bL5EU/xtcymXC69gF+1g2OWpbcN8tI0C
tX/eUupq3Gr5d2Y/5mw5YAEPczfetzydE971nYY/qodTakStdTfy2pGH0umCoQE+
c+vG6KbKF2FCq0E9Jtelet09s07Glj9cwfdMz+SNqF/KyHj4dgfBf5gJiLMtiObS
trI28U8SQ29Of/ztXdzDyEet0p0n9dw+5L/zB1Qfz1p+NG5bFIwRWkoYDIFJytvC
sP+LZAtfhDlxWFzwMfFxSkvgJOQleUq8aXmH3WYX/N6rFFPX8MtKSOkz6KFG4kyo
be3JrRD4J9NGo0sqquARbfpHrbWfuRMx5/RUC+KRouhkIskUcLdrcMu4/brw8gNw
/7r9N9byyJiIKQ6k+6Iphws0I9VeBYJK7OluKGvyjIzd/h9o7K9LcBR9HzoOHxoc
SItWRs9FUJevwsh0gHtCAFeDp5KMMrOWyiA7FRVJR0DL/UChnA8NN8Xyt+9TlWXL
gLXkOcQ7ON/jpwkoIYBfre8e/tcIN02xwmhSaoal9tu6sEw1xgYGrPieQaOLuFBv
qHK59yTP9BpTbMO+1VA3zbkgR80xxBVdl5fFsapEdigHx0I6uc3PrwBtBizu9HX6
FIHhOxMDKw2U3XWGGlf1yVXdfj1td32Bhwasi7ZaLSbD/QE3N9Lw3fQGI5pw1MrV
vai6zs3taCjCsTQZwmfxR4SBBHzuM/VhnqoiZ1tIXwm/lfInOEPiJf5/2tXC5rQH
HEAwKtpxfJGWsiaBK/Jc1uBV1W1a4jXU9P6X6QhpM42MMJolGMlSISzONrrZ4ZJM
nV8nXpPPQnDLeF7BuvqYcgFQirR/Q3Lwu4W+8ssxjvG7+S0XgOJhH7mB3Mybus01
UsG6qoFsXIAzHk0Owbo9ouOsuxWOL/sKsXjXE3UqVxPS41mevxVzdPUrQrTDTjsB
R1B5I8qa1jp1Mj/U4R6MNegzNNfFjkJ+3utjPYev/dsmsxjiDZ36PyM68/q0naMg
2LTwIvwsZEyHZEfRXGYhKV5qrI3yNRWT95GKcn4yAg3IQtPGzdrz4Sl4ehqLux0y
4Ozig1D+UQ4bJ6/6I7LEdsYyk8oE2MjLCTw28cdezLC4yxzP5weActpIkw6dQ4ej
+ttYqZRPQV5BPfgSKjR6IEE203sviMwFDe4ioNj5W3EBZTzBtDruvptbygpY8zgA
FZ1swutUliSbSHpMvsMbEUzZNuwjq6vvRg04XpFqIKbmfyi4VCEG/jwSd9zhBnV7
f7o3BXQeKFhMGRT5QM2sH2fRxCDMfi8dufCWvX6/aKJW2P6Y2o/6rXO1zTOEXL+m
HtVK9ZFWpyw1fvtlqJC+rjJpOr9eLDzSVvlbTitok+Qq7gX8GfSxWWc48Br1uyNE
BU+/MrTzRCdrPzB8mbhXG5HUE2AsIka8hoaSLnGovTfVVjCW17oYvW9yWROzDwdQ
tiJGYqQt0FFEY6XetDHdt/qsBZ+ENoP0ll0Hqj5kqvfwGoEG1pwuxTGHyhv7VuoF
jab2jI+D0EQvcb4kB8GgR38EElOFhdY+gjs4YM6nBKoAw/b6GuFJYpfGhisbVKB0
mdmTMK1TnL5FRbmvHHtatR1l63+73DPSOj32pCCKQtuEF3g1j+wC+iq46u2Qq2s9
mjtlT35x9Ta3oevIzal+/MNTpfb3jXdsxnZoNxIKsyunZP7dg5LmP4qXvqbhaIbs
qMba1jW/RVGFG/ZXglafm+mKNX7/BrFl/BcCG6t8zFzaqRxPxCIOY7tL5u2uePZ0
3pzJ5OLzahzAEtv/LzQBlZn/3/oGlqDhQy3Z1KbDbZj99oitzO3jnfMN22bTUzkA
zBo26/bKCkCrDXAOAKdbwWegpLWFUn4d+63Z8gsTcwhjO5Tvnj8zYCi9YY/LD8DA
z4RxkRJzTyQe21g60z9vmCGw5eCT43ujp7BgSd1xdPfDhLWTEwD0Hflw8C98NOPx
nMUyZOpSV3r0AgCGyLQqVVl6UmPLleznPHOSkGmYuGKKI3Cp4l2J0v1powEsP1o5
o+EY7yfNAX3bSa9ydI8u5tzAwjMTuJpCdiPp70USyrFPTgVl4FAq7+6oGQc9p04b
Wl+hsoPN6/H4TBoVBn1KOTZZ1yI2Hrj5AXVN25cBMMAWrkydevsaKPPWxAe79XbG
+zlkjYJjSQv6Jt/7Vri84JeFyYwfxD73jWHZz3usk2X4RPzuMaNQJ88XDN/UHKfH
x0493PEP3BkQ6gnaVdOVnviAkI1BHosSE0b2DKBG3qepa1L1QXygI0z8ozv6XoqF
iiDI1sVp3sZc1DuIcQNhzyh5xo54AKcDZmnIf0H0usel+Obb0KS8uOm0qz4tTcnj
Y65QRdJ8R2yknmmdXk8ZkzZ3C5+wqwIeQKw5WIeT3YsfDOq0GdrSqPRPHlnKZ8Rs
L8bVS6ZB32btk1/talr+ZL46Uwouyclbtq782276RmV03rEdl0y4pTqlXDnfH7KF
6IOXq4B8wbkTa4eZG7rLV1OYkFX825xs0Wp95d2YNgWEmerowKRT9QeWnvuF3jl3
Y1qmNCPbNv1mmpW27OLnqed0JE1xOxUwhoK6rILs8lh+U9FApRndXeNtNmyt+pC4
L5SWGApMInKFuF6eCtYL9ci2WD1eAoKzec2cyXBz0nox6zWXPhpvdcqylqePRsnB
z8Ud2famWnO1jUBmbxur9d5RA0ZZLyAFXpfOxR6sSfxCAT3rLL8pnUoMyr/9DWqj
wDmmKlsYZ9OvBGbMjhh/Rn+W25qbU+tK0havWU20eXLSsiCNAPdY9sX/VbCUk9KP
bGN5azROUIDdUnARjm/sGqwPSgqq9cpZ3f/okRT7moJtrYFi/D7LseTKCAsUcBo6
RrlfpKsy5Q1p0gpo+UJ5Pb0zd8i6ZSISleIWtC4LYhSmJtHEW+fk7WvmLeVMWseW
0i8lS4FFOzVPEG1clw7RdT7FuCz8migpVGdJO9iAZojzPVhFxZFdcZeifTP/OhiB
adeNAjz2da1/OuVfdT97bKjjx9qwXISdeDWLvowqiDTwadqf7d5jYxkHPUX3NGeb
ullvy0u9h7jn59QdjbO4cP2SfjYOfOCbQDjTkKqTD9lwkFC65vKDkogQAKrd6WRU
CTEoLa1jnqYiVHdFO7Q5df5JgIfVNCnGHqz0UhjC+JLZdGIz/cCaLxxtaM3sNm2T
ozDFLAx9lBXOW4TNMrxhIfCOBedOaUSDI8z8/rmaj80gAu07gZSnoOvqNbYNGnwc
swIJLfj9L2xVzzNd5uu/vxSt/oDHznoHFer6HvkKMXcAxZoi+okgvJ4UDRfv3WL5
Do3ZvGiaoWGU4SJzF3JsCzSLBwOe7CTJmxZsqmO6SYDsnLcKq3B4XuJdYqM2X85I
kZrx0O9bVLA9U+16YNyokmhXcjC1mMzSq2EbdpiCOmDplv8tNxM0E3BGeQQFdJww
l5L5flraCbARC1gBEZupIKfSE/m7Ybf9GW9yRLVnfhyjLrCzOYWEy9ySWqDl0eo1
b+mAN/MdnaJKCw+mjrNqxEW8JnY288806c3S79Y37F2kWwf98sOEET8DF7+caRZX
C5++wX6axQg8ni8c7lbgT/ntydLYwzlmHx5WwhZf4LOEbLoxmyE715c3sjmGy4DD
r3LppbLjbhMMN/3IIQynX/91RCVpr/qitzlwXLSE1HgsFuQ7yreZFyW7rV1Oj9Xb
p4hA3AjRFueBjO+imZCDOp8wOl6wlp/PnMogk6MalWVbg1zIvTCkR15koUEVOkgk
9rQSnarHyTzOLa27Ysez2W1plU5x835QDa9YT+IuV717mvg8/nGrLn4QR1t0aUV3
FOtcVUZoXsuq8ZL/5alhU+PjWbXLOpwKqLQl5rF2mBnfprj+lyDZ0JUPdfeB9d/N
rFPipY1leWTvwgG/BgxAIsx5jzBE1x2HGa9W4WtvOHDnlvJTZuQcSlgm6XhHJ4ip
2t2tDnJIaRyb8r0tUzUAfdU5vxddPkbuUFYwHVbotQXXZ2by4CMwAy8OBVSHSng1
6oche/bhEBR+P8yzM/3KtIoS7nKHSQFF5rD2k9RR0b4EaJGja+VRq24hF57jdhqS
Yu2k5zqjXdyGddhRVnCOIhkVKpnAckzvcg+8tiGF9sUqnbomFahGozc5s8/q55wp
KTToEZ057SA1LSqDRks805uo4xw0TzeDaajmk2SyxbTvpdwKYHDWK65IZ3ZesL/v
FWzI2IYzdmq72ojL9ZigpLF3NxpeuuIllholZBLu8nPnRRd7dr7KrclLQ+M0otMI
56gex8xMlZUT22ROcKVuyG8k03zJIKTAb+StPLJCelZgJhzHRrp3eV+BezIwnRz4
LzKXwxjFXmq/Rh/v/o9nDqzSFZSme+btExYtYvbdY6R7jJKjVZ8cnMsRGTq+d/ub
+AxIHejojGuhf/GR4SRw5V5uAbv1WQT/LhaRkh2trqQp50N6Q+bGw28EkZf0jIbu
JkwcfAh/9dzqd2c+jXm9aHoJkgBo+olAJ43EYRpFPlhMsY5u7zZgtyf9IecLodCp
wTDhjSVqA48UKTsS+gw4XE7VMn3TramZq3n08hWug5t/aT8YvLiUrLvvSTmRKmVb
N9LKj/6Els2XKuH14VIyPdS6YgMOdfQMDhxq035ilyOr4Q9fJoiA3bIimhVvkpFU
aEV5OvDf/TNCNMqR+AVzo6BrnK2wlUXplwVxEOB1UkOeTpjGGWjlJUzWZk8mOhjt
3hLWCxLHUp3gLVEFod9BcMiLJLth3Iuf75JslohZpNqi+S0r+70f8rb4IZmmbR/f
UmJpZgnaqoVCWeFKP/V9x68pmMdlaQR3u86AhdpWW+Ou+SL7Ij+214L9gfnX97av
OnVS63ZEIdHfn1J81GBnuXDog8l6gMjoFiL4C9dcZWutPkScjrR96TGDKmnhRvvb
a8ENc3VANHi59rwzIGeb7n3saWtxwdvoYmNDzs7XKwn7ml68zK4aFDjskAHI3FJN
QHyBWbr0AfT/77OzkdE9P2GPeGBZxwSeYMKj2PgtsYW7PYrD65zelcKIiFMS7HM4
UMpWlNjb/nQ6XaXqyZLLJvol/l+xVPUwbkVQcIAGEnKiPmAXqCaxzkkzcFo8NnvZ
akTxox+uVZEZl3c26bHLO60crLwdcuroPZRaM8OOpLd3UBpwXuYQT1PGRJspvkaw
AcGRcmyZs4KpJQAqNR4xCbxaDdfhxKPaq3Ed72EWX7D9Am6pJKaj9+vOqVzMSktf
NWP6i70RQj29Onq4XWGtHxoHfFecotsf2N0sryHNf0uICij4gSC9M/fp7MAYJI9u
VNkfabFLJEQr3QOkhbVN4NAPq8aFTFSvgwuSgbWZcmLLT7Baxe/tkaSnsMafcxSJ
aXrTl5bL9iJ6Pv4EuWvWlSL0Ra4sqfyuWcqeByRBVK1nAglcMRElWzmzuQZyR9cA
mkz+J4LsD4tIV2UElKIsxuQBEnz2bQp6fmkPUlVhuLHIZ3ZtYUcd/t3YBs3GLkly
90LrQdC2PGtetJ9R46wGfxbdOA4M/GuX3iObN4orHn2RudfGULMsm9atAz+bB2RP
jOJGeUv9ArRrdUZ21hnU0LR7YmVutgcMl7UHARaiJ9+TbskIf3MB7StZPjCGV6IR
qGgi32ZFV4bCX/1Sm6i//ACE88iByfC7w7IlM7QjzQixBYTozae8zGwGC0H7Iv2X
qdp0TxJZqFaJRdmX1MCO4Z1vE7mORgmN7DiKTUraNRprTGAKBLaauenY+ye10Y3y
KIpcGt0R/WHVvAVaRWAYs+osS5bUwwP9jFe5wI6y41DXk4plA2TDUkOkgNFtjWkx
lNyoOwmbM1rmLs/fw9KfTqPpa+uzPstRH4XsplIi08mWj9oBIo5uWAKHhK0QzUi5
X8aTOqpAbXlA9mem0IU5Voa59kWjBjEsO7XrkJBCZ5piwSXGdmhP8YUBf4rqLfUg
zBfKENYhpnnWp49+5w2Dk7whbRPFqQfSBWXhgpfbEOaqI9JFHZoipPctRb0cUeUL
D3nueVVcxFsNA+5GnN5JQw+DwYhVmjn8l+S/wdRkl0zyGoUwCllsa/U9XrgKVhG5
+IBUspy1g+y677C0TV9aqujNCZd3DMzy4wqTG8NSB/NsR5z1F6WVwshV7+Cd3aQV
3S9KvfDkxvX7S+TB/e201+ZGSjQO/B/Wepwl7pn635MJaV8Ddd/jMcBVU4KVtWgk
3X7hdI32IAieWUIfl9N6IRyItcahjmEJVlk0DSuQkLYL5CqgC/z0KJ2inZ+w98u4
9FUE9ZLxON6lQZUGzuz9ceVvBr5YqFNRP4V9LrRJCaCd6vGWxICgT+6xYEScFvzo
/ssCKWpaxcWSiwU7slHEnA6+Vc1ftiizBDBsClawR6wLww9NZNCBNglddhP6bzzc
m6gR6jm2i768z0EJ5wXC97U9NIVh6Wty/BDi39n9pc7WzLK8BxPLBALkI+jRo4xe
O39xUPa1sgGYggsjUMmZYDoffo0kDeZAgeJl8H0n8IG+16cqr31HhyEiRwcptQTb
lMpDz/OQHBerzDKkg5q/0CEMulIC91sx3bZ9fQNoeQ1iVcly7iISmy8dCUnIS7wZ
LUDbs7R7kYQnQa+WCwFEkhKQKXsTfF2otyv3mGx99Lqzjf3gmMW8DWTbUXKOpepp
U8xdx0nbNkGGCDUTe8r6dhG34jR0eYm6pb84b3kv+BMyxWvqnbJseCArfIItQ/Kv
dS+ipmIw9WkIgAo0CyFruzHzzkyED6wCKZUs6vjncebWUwlJqxupPClLB4sxAp92
Lci+YXUxgKlFbfw9kJObd6swZfsqhDE3VzLNg5ayPh5dUHovFCiKlyrFKSqGCx3Y
/9nAYpixOT89u3fpgOnIqrfMn2KXL25BDEjxOzneVaq5VECXDcVkKkQHP09KY3Je
YCM8bGkVE2zDUMG+aWig+aoRw5YMbmXLr7Hh8l/Q7/WtV4kclCvSZ3cyYBUg/pXY
1/S5vw7TqH7sansOYHzvGyrkfQeNhh/OGAI7vpKheQbeh4RozidHy1JpuHnSsJvY
Kdfy1Y4xupNvF61OLvjONcI+fe1L0znSGyf/X8gVOxGibNNopCWrp1OSFdyKlscX
I2TdrOvArojK9bVjONUKv7+G/SN9H/AAkYlew0+p9lVAIMJSKTJ5UYzQayaEcJb2
W4WdwEI+HP6yg0OeUm7YWLhiTX7WL7LFAleBPR1wHTwBQ0oBuleWLZ7c451DpQMN
N5fzDEREONvChwdrF1BS+DEiLbT+y83tw+XnvZkjEwAz+f/0/MJE5QMh31f31oQR
aueJBVKTKuLvlZqjjX8GOcb6SvoDf7IIhI0Ny6fQVQUywp7bLIrgs8jHNQ7s3zsZ
Vk1wEQUTRF/b5XbTN11qqwGYnl1Fs9IeilfUsm/0WrLYZ/qOFW3KSiTY/cWtlPqV
WGNX93z3XRKGVi8vHLMlOblMkk+t4qLf268uhwpR0qmede3lCaW9ebd1aHFm6Xup
BsPJEg4+y4kwbf9OmASYD2j+sq3b6DREXfGnMGJSJN9AKWSwrcQnNdIdGgt+Rap/
CGxT56FYestsPNVmI98diJ6Op6loxQ/mMt2X+hr2fAwv+pssdstlhKcfKazR5Qx1
XWw9cth2Epyi64eP9krsuBiJZOxIQQuZl45ld3WS5r9YjFJhyVxR8LZvsLmN2agH
44lcOgfqERsAOAjjD5BAXSX1swGQdA3BUgkJJXg2VY1uyGsCPU2lg5ViTHXCSFT2
jvZhZivN40aF/T1zXXUpJOPo3BfRgFAmmZ7remJqj9u3u9EGP9sviU9IBFOxPyYH
9dfEefat7FSWR8YBprWFdh/7l46VsTlh3Nm/JcBQcD9CA7Aaa/IQ5yXe7hXMciBm
fApnAT/iepl9DntDzzNRIhncL8pHMnp3M4q5/SjO5lrJ8gNJe4tgjhVmKhHlgJLh
btRwd8e0P/ufOqbUl3X7/I5gjBI+rqX6lZLjzA4/glWNYpMz6XrNJbXf070ePNDd
ivgE5eSBRUVXE+SOl/xMGvPAOo2MgcLuPIUDeLLG5UunLYFdZivWIviXWHbMv+E6
Rqbs6vV7vo3yL4tafmKGCr8lIZWO8buU2HCQ9w37Zm+HIdfFE6PfgFxj4WslqY3J
W+WrnZL5WFQqUo1Ny1wsT5SGXQuh/ZQR+hwKOQuGiahi89ntd6K1UUk1FIKRDmzy
0N5agNXYjnZ87qkcYGi+IyFbNwHAlyukynM7lyeHSRfIULs9lcr77KYqk6QmgdS1
ktsz3K7P4rW0+WSucTKF9qDtZVLhF58TqbLdnvxtKNgGOcPRnUAWQ/tgh8MhcvIL
nFOVFESt3u5Ajcux3vhEZfKycEQ7GkASxRim2YR1AqUKhkNM5qVN60AZlbZzg5N6
i2Av3R/TkA/wSgt1jII1XEVqk2RqG/h2XxDI2MOgzLQl9vs6EwgTbKbRaMFvkRcs
LohXgx7JTlOCAeA6b4LDvOueNCuvl1p2QDxiXzcaDZIFdgKLXQYLLhQtZNk9g+Dm
su9n9WXXsnEN8LfpgxkHVg7qnb4Jx2KzXabFu2Mg7CtheR+4fn8SngxH6TRShE5l
bQSSMuyoh6IqIsIoG2JnBnm1VfjhMaERvCDa+yTKyJLnyzFzAYMvQt6ouA4Tt6ox
bGJNZd0aHmmLMMkXh23ZeLB4hCtVk351osHJ0coOFg+tOLKdMvyyUomtafIyvIwA
n0mXESyyZVs4NaMnD4Y9J16sWeqPMxhES7kqABGDpcxEOhsjq4k/VAQUf+FT7Uyk
80ZZBeY+nF+QIhcyOwKNmoAz+Ffa7/KLztM/s8BdxIvlDitNAGYkLupSvYb7nivc
d6rRAxKCH6lhGKXoiN7j394xJnHKcxlJiOQkKIM7DBt6vUBR5bU30/kUFva0tnhq
fle0vg4bHgV/gnKAQ9j5Ucxc+YqLtTjNUhMnBZ2pczOp41COpM1hm3bk4/KtFLm1
XJnP/B6npcdyx9C3E9SJr0LNVwidoxkv9fwKGhnLDHnyczT7qDjcduNwQ0yEyBgA
co5WGboRJsBWemLKvxn0n0vy+ZO5CstSuGGUWfAAsDJ7BwJtSuMzCR8UTPwtYS/8
PQx2pycdfbdE6YiGPo4SYJpXTMeMlNEATd/vPycVaRvtQ7dRP7QQGXFSgJ9/dtGf
Oame3AiMcbD1NYGIsEgAJBLljCfzqj2CCaU7fJ7TrXR72NOBizfwPMV6f+aXt6H8
HpiYacplyCZj7Hw/6VCEzzTqFnowqkO3P3Ig7v9q3HBYoOjiU2nFbUXH6TfdIEnl
p7zs5xZK9n5jG0DEL2Zgpm/lNVaCg/D1bdCcgAVN76FGmtGH5BSgB2h9ZBg6Bdfi
FVeE1d45vLHpkSe+/z2J8mqiSTRLUJBkHkgYR5kG5XyBLdwku/oqGl2yYjmLii44
VshyGd8nmf1OS29sCmIctmu7sBc9vFTrXq6Xs3WefafMmjgtVixEP+9AQyJb5B6f
RXReK9IbziqFD0n/egEbcvOp8zVqdZHaWD1bvknAifOYbkkvGqKRVQjtZoUE/GZd
fqmfctlaLY/9MWBSg6FJqhY5fvw7IEP38u0X31YGrMg1iRFps2sme11+vJTTyLW0
PEgfC2u3vFXOe/rweWeSxtgHEoLpDRA/XdTTPl4CkM2+5S3KFg8UBowVIIMwP93n
Q7ENVB262qNcAvV7sTcS9o3DUM9QIiBbblfqup1cMRnz/wqCmO/TysCEYiiG0G37
Rt+zviP5gqISrCTrR18b+CqTOyAC5W/15U2NGIhqZ1PLkiRnJ4fmP8ERMU13Vg7i
f8jGCVwrfI/nx9dxmP3wLyWqn4o8wAF+09QqjvSBXGLr7Z3pKjIgqT3Pdpflqjlu
cL8cYulMOTvUDABWg0byt65MAE4sJoeftrrQdo5fOr2lRWcBS9ZGZXsYNFhyAEov
0NS/fybjNq9DnNIkRXcG2nxMAB0IOlsOfxgIGxcsNq6R44+Lp7RwH/14kBVCA/0+
Os2UAttuYHCacdHhdfhZq5U++INkrbZhL1lvVStXVnTpG7jHGOO1fEwnTIixNFI4
rftLZK9mNSywKE3KYPj01cDbsEIpQNr/aFTIl3o2ts+ny8ecSbSMLVS72EUta7w9
SNdaxU5ejDlbwUzkv1DxaAM5GZlGfO1ImkDF6FKGrqYuTbj4ivaviXNjYLBrmxid
lfXyfeROT1M7yc2vd3FrVp641Ighu6ee63nIUiH6vuEYwahu6xEWeLNngxC2f2N7
SFSaWCUFmPz5jjkbnxy9K2O3sLeJ7UeDl6m27/B5angvIMDdXVEQvckhBYQqLZOS
P1vApPyn0Dc66wkeDRGOAAWcYNwHLQrhg1qkNHtCNCP9+eo2CYQDz3JPvXcr/n3f
lEL6wOeAdjwbpsZkkNfdSIkIhOMYI1cdpCaq7FA+rP0s36DOW5C9B42k2FwSsVrV
GjEoQfqmtz1RpLDFwrqxN+8n/uQMVKvATZ8JDe41eoH+FGPiWlP5G2uJnoPxbf/E
S1RYSQsrbqzhmJ+q+jBd0XCYdqWe1cvITE6qiGuS/1mOe8ioG5NDUhsRa67cZqzR
ZwUTKvq7dCWl6MpLvaHDnTFZNrFQoUCP5soGdRlx77oXmi4It4oafajaK+cJEyIu
oLriiVQreghcyrSzLF3p3NlX8aM4CsXe0+vEez2HLzOzQymmKkS9AQULWqk+Xl42
3yy8tRwokGU5EoufCDAiPdPtYshkxL1WiDpKupgGWSLuyVSSBkoe+6kK66go6x21
TxgH754Mti7IB2KaNikj4YyPWrLHQl1llVGBFfXIcQQMOfWtVyH3pZmBNKU1f/vx
uGBZCwrkyrx1Xc4ObPOBU1pAe31ibCeBSig2MZRLS2s6F2IaOtQDPROYkIlXnTd2
y+S/xd78VH1ilRAeQC1uAr1G66Eh6EV0F2gOsi8hvGF56t/HczURHrQJX/6XqJ+a
91jvHoA6dVcsQKiMpQwJ/2SZN2NG+Hos25l2TBUy/0nhBu2esJaRVyhKkyZpVzAU
wFor42xc8FNzSnwLhDtF5+ctQIhPslzEZciej/tKh2S/0Jnr4/KBoK7mFeNOUix+
4WowQF1ZHq2v4IDVq+inzWfckn0fD8hIvg0PRle0okL123+SpnpeiCp18i7nagE6
RPYUOMjSfhVPvNvqwmIuC5ggboUtvFjFlopEeiRmp7MbP4R8tUhp0KFAFLKzf3zv
Lmus6YDbhePTMpbstrnHsNt4YOrBcyE+6lJyLjNdkFqRsq1/1z6TWRaiDad6NZaY
I10b5h1C+0J+vPQ/zqGqwMMS+6mVJzX9x1LmmBMI9zspqvkzB1FNnwNN1Dz1PO4u
r8nyasc1VdSrud6v4QPwJ83/D/W+Fuy3pnb2JmntGpVtSWGa+dKipy2dL8nciS6h
19HQmwreKPnO4SLrGsBdZbbNVxbZD3JeyA8Sbh2bWGfmAsYlDa1w1wabtsZSfWeU
Iolx8JzCrE9U9Ro8Fx7BXz37IDSiFKda77Kp5O/j0+J9tWtumWQvN22sMkfPW3dS
xw8KUcUjw9fu7Pn+ZuD9/vjGjiLE763OnN9pIsYWR2qEVY0JPr8OrsaYIhMZiqG6
NVScSnyCBZt1xf6XYfwzjxh5IlQZetvPwOmru23fvtef1OQpPkTqQ3iuwKlzAax0
s+teWnSNfFqWuzUuAHIPGdNHpT9KgD7P1BrGjEtjn0frQKBITz9G1GxHCDBwtY4J
EZT6FZKSQd4cGmw7kvqj/B9y6mP2K6wLo3pt6OiHddoykDWiATKeLl578kuYDpRT
H2Wh/DvtKUPIVVaSD5zf3cHk08sB8CH3mSScg4rT59SDxgc/CDdNbpFAFTPOHj5v
0r7hyF+LkqepVdhLOkY4xV+8LNiJ8eGJbBESl95H8RGAVojo++t+SoJ/3BDb8Y5K
jiw/QnK3FnEo9nJpqPiSOEg9g6QruVk4yoo7LA7TIfHiThpdlEML88AWkOJcEodV
7HcFoaDg+f43DNudWzZOj0QF2Qc41j0w0KYNBLVIn/OG4LoPdpEqKSc9fIVI1mGf
7VUQhmhehl0tYOGzQNlU0WhqoD/fUUb6NH5AW1FNUy1CxeYf7ES1Wf/z0swubnfs
rOn6p9KzgfrzAxRl7/KNRsG7kt0cOW57TRuUVzopYO+cWlvRNpJoFxLXPMUlKaps
OHIZSjSOGanwikjYj1xBjN0hSKXkbFEF1YJOct1xm9S2LU5E3WYc+oa14f8T4LyA
a49dJwRbRVAQhwZ8ZpdsTt1UOpNae/xlNM5X6925Emu0vRHHr2Ev+l2arr7gA6Xo
LJGy+mIYGXwz0/xY9EZWCwyi0JpY5iqXZgHvTnGO049SHonZMEdtyH4U1TKRH3I7
AP2XgMi+zx4WWo/nFhoiSJaftzqOhpvPkocZAxoAaroPZCtwcbj4mqqdtN7HCwcE
8JtVIzR5j5qeZTes3TCx3405FQlIVuS0RAVXPbTAjLnfCPh42qpkWUXMxj/5Vu7y
hlXEhF5UtpgR3vphUAnHhu4yjo5BA4vy/UJM1i3Ti+kOSmHrAqgB9xCWEu/UWDZT
skH5pQJ7E5hgiXmLVuPlkzimEfY9d00gWoaGTTZNFvXnpMdi+CQvbL+SCwyV6FIG
0mq4scQViw3Qgu2iuLx8TjwXrdjv0NuLdtYUxA7XMrcAbCKYfp2qayeYc4PoueWM
WuOllUrej8aHVkXfvX3FXSlOq8RHqKAcXd1AQsVGWA1POvFiqn1R/epqiWjrqnQ+
8np0nZuI7FgxIMOPCYEpDAr8H1K98nj1tuGDzoSfL3bhKyDRiDuj6xaXeR1hU906
PrVHwH3d1/2mQhKJQ/MaNNKfTJoe4gBBOqbR2bFWvWEaQ5JzZAFhyQfpEknhgd8y
0bCtfD9jluS3pVWhjDWph+Fm3N9AydbspkGVtorpegHsld3+j2Goo32hpO3cIBmJ
JWqPWwpyW5PnmaDpGTfo9WqkL0LcWKGSB291BB8aWW76w9TC9NNAXXCS8RtlFOTh
xcd7YULI7ZtbGJAdkSfoPib9YenjYu3QeVdnuM8ezjRWkVHWC9UCKGjJ2njU4rIf
oqkumdb1hzX7lH8OLOmMRSye9uvuQduKNX12jzCpKRHUCT3svekPPc/SZkTZiNZK
7/xWnNCQOLJhH5hzwckKGUea5gjcYDFRpfBLQ+TGcw8j/Rck7NyaKnJc/ktXc3KM
n0Ow9UG8br17rgrQL99iAWZyVVR5578ihQpRNVnzKI/DRYmaqvjeGgnSYQ4gIWUR
SLr1zHcAbUUAdZMJh4kQtGdcnE5KrXLzZwdvdESa2clXLqG+QI9s4U0OPlfVMd7k
z2c8Y9BnU2ZqZ8M+flajTkgT4AEhaBJCBa73u7oj5xIDP6KFzmepDHDrakT7ACWh
GSI3XIEIG0TBhnyfWn8TxRMQS87FO62xDJm4AhAwvgXB0VNRMMQqt/WnQvXA8Xdd
RWctvFz3jilD3kqp5s62BrIA3c3tr/b6HWdwkCk/UpSJPw/5OQkHdZybiAT/dVN1
99iIMvwG9/a0VEvQZuNY/jLi94iO78FXIeDJSzwJfdKl9VrncWKW4f7s0t3K86N7
FGIRSTag395oxMQ3fXS2VVE2218ZNttbDqpXcB66PwP7DPd+Bga9OauSZTkE2QP0
kAmPKJ0kML/5RJz+CR7IH3ltKloi0KJgwUsUzpj5LIzHcIcmf4j16jtldU51vXKt
U9GZRgopK9p8EkbhVpe57M6wSUMvZDNvdqLBbRti+Kt+atzMP26oT+ju839Qt23R
wjEpsazHGT1sLJNVI+iWtrGDeSS2PNs/rvWCeNIlzdiD/+8hGXNE8GEYdQ0w5X//
DS2E+wmlxbDRJ1OQcrIOp1hzQy++g20QSp1OKMnRDQ4A7I898GUuJgd1G7X2Uzx/
jnOdKwl3i5PY809O0Xr1rNRZ5I7+KwAAIWVzxtCFedK7hPagYs+Rq91O/Azvl0dP
C+HOSHGwRmJ/mb7sjewdxPzGUjNDTE1H/q/siH/MV+TF0vZ+bcf4/5IRBciPiG0Q
qWScqYWLs40aJd/RPsz3s7ZqMkr3D1dqc6OJaIw3EX0kUnCltq/p5LVDb3ElNQdV
ZkrvLA3jRiHQdghOV88CMWFOhhfBVmGadHaEMnegCgw35lQfsMe3VscPcBNzXQow
hG49zECtnuoaAZ1ERPxo7I1UuglBjto2CSHd8rKuttDYi5Bubn5XT3y3bshjgTxX
QnoFnonbx3yKfk57T/wbO5+HE1QauJk3bC+pIV++EcjNJaMBec7n8pVnpsAZdzC0
FUifdxyo6h59drVkkvFJnqApaxIFLIXLLwNo3bGfIhZMB//JuuztVAba7B2lrezq
sRXoHtQdza8d9OMN0IHDWtn6ay2aO3mVNW51nRmimO9z3Wu5/RTMDXjKjWCnxJD3
IEjOCy9uEASsqtHLiWdeYBWWro6bijZMQD3anCtkDGmNcEMdDNqKZoUjJ2Ewpt/J
8nsXizRMIlYy4QmRYH2CReu1ckXNbXrczg2mhY3sedb4YpxUi+ryzBJNTopRbvJc
GHPxf33baMQVVFUvb2dKLLjMUalSwXbFl1gydbynTKjCa0OYRwKbfR0IAC5frtrY
garGAM9yzzsWfLGboC51k8IKxW/dDwXDOMxsyCw3xpI29Q7H++Wigotq8eLp6875
usRYrNkR1N7Z23qDBL0cfr4KBCLDXPjtqXDoLGtmG8zJRzeiZWxqLWZS2dbmQkmR
lpcJszWYSF30NxHXPsUYRZBpkNZiAaf48Gy/XwAapxrIjTJJIws9utjglr25kT+Q
tPJ7WNJ4WBWe4Bu5kPIpms6CMdwBZzPhA9W12b0sFn4ZU5FFYia3jotgfDTUVWwU
cslYnPSSqH9pAZWzjivbpj3jKEf5L2tL6JM+RG5kKIZ5NKZbx4sCRpiYfBqCxGBX
fnnhdahPYdghV2CK/LAfxDPNeDMm+uTKrLxhvrc2PmxJt8kTPDb+S3oCHjjEwfub
OWQycRPzViz0PnZWJLiBvFo2sRvn/68ecUqWORDVgtas1KK0lidqK8JqARuVdcl3
nYnx3R9V7kPEgdUIucRRdalJh4sax/DSEHDIdd91SLy1aNPtNsjoBnGncD2ux2bF
KitcWXMtXBMcZL8X0dSzaeE+ztqa3inKzzeBnRwzY7DmIOQU4Z79eFgBrhc21Og7
6I2tGJVsGxpbCNc1b8KCLew61OiXkhjLz2YUhl+y2zWslZDT5mzoKeb97jbje5r6
oPKfM/fPbJdyKvf1pdWyfTwgBhRgmwYBWiTIfZVzc8uIlOSVKvC1wEvY/EbfqM+C
Q1a1330MhNLQ2pGeJn/4bt63xDVn0WGr4LgwBFYgDCCcSs3qUi4qw0Zujf7KBV5y
k7pUz5N5VR1hcPqMIiR6tgRr9RxW8930uiyHF8iWehnPAVaQvkIwDCrV5IeGIVxa
4Ea/7q7EJn5553DcT0xe5+kOAOE3McmZPHKuxrw5mpWIvzIrRw63T+Bb5Ol2V/0x
ZLa5PPXqZse43uvn2taX+DT6X1QoTXTmT8udlzULxM3e2rGUA6etW6eMn4znQs3v
JWj3+gIHEig7x9HY/iMd3I2dGIU6qKRw4Z7J+YSeTl8OIzdbRXMnoJvG74wqNNww
kJ51FvPsK3xcfoJLjMWH630/DLQFbHAxhYy0t/PHA0DjGZO5w7feGLz/2faHY+JA
ptZYwn+qglCNPR95XXCGVH5mz2VjKjjOl/mvzycvSwF2t0vDrlPuN6YGXNGouM0T
+oVF6ajLPA7atBGzF4Cw4NmW3GQpyyxMXlHJKqlsbY8VBEStVAMUhxZUaGzIirdE
JA6swQ1n9ehdMdw2Ec6P0aREaAmM6c6kYb/q9WERJMQa5LfO/pqSkVcd9YIUxcy6
4AU3IvhiicvvsMxnGqGzDdjsGvTQ6cX0ngFPjLAi/B2sUlkvFcTMcjgEqW+/NAd6
O9m8/1Cs/xCS4zz47ezkpKPZDy/QIax+LKsQeGz9TzfzgyOy225r/k9QeLo27GPk
tQgQQ8JRdGcPXhq88gXiwRJF55HsbWZ8vKeAc50zztnDKEijvzd0EFERTDguzDn3
7VlBxDqgJDNHu1emwkOhdTzztYMYUec02bRQX6HqRxWRRqvneBw6P45sJNE+z4SL
fMawI9mC7YgoDJTQosi+vxf9KTE6B64Vu1Py1OMC3Uud5ksnQ2f3rfWjVm7lfbxT
0deW+Su+57+Dzdi2jdot0t5koNnSZH6/JhPsA29dXnHFk0avR6psBPNT8N3Jn4Nh
kuxLDOUjwv1cXz90ohfBYReca5ATN/rsZyX+ZYJFy/iwExUfQH3PAprKgsPBRSol
A9yRRLT3gLx/5oOFQ8WBvJESVx5/1F9TqCwk2HssBbs9LQf6iR9FEEQhqUY9rkF5
M+7yrVpPIpTOM865ebnwx7mxGriHIGjzBn9XHKtYMbvmT1pMT2r3qmGOwHmSwTV0
d53B551lxolF6XwxH50CfXmuDWzEIdqF40ePO3gOPhv8x3MsEpbc78rNDWpUCbKK
EQ3DoSqpOKAcfVV1pj349iHdpWmd8OJ89YuMMZuiIPa8ywfCkOahyVIgoz+jaGoQ
3QuLDGZ/AFkRitAgALf+6K7VIDMwhtCxgkicSsFJyPTqjfkUYRRSNrGUygzCJOdq
i5JG6VPmugXGTSUDVlhYk+cnQxoPcaQwssstOumwUd/TaEkOYqAGq4gnNSBHJ+jh
awCTntGuQYW7XAF/BeWOg77d5vrVo5BRwlEs8y409RFSSs0FGYGHDrCUUh3sgya3
zJLSoNV9Uzdzr1XboJt3tPXu1GQcyDv6RUxYgx6BWPvLAm81EZjkzUbbJpg7CGAN
8ZHxZuFWVo/+w/3jr4okdKXp60H3oyJTfHY8X5Oc74sNad0IB3oua/VZlyAsChDy
KlvEYMzS+mGhTZ4YECTS3dq6GvnEqbhsXZgoIZS0r8MwuWk8R1zb+AdCLglhA1JQ
qKsssfuuFc1Q56bxrn1B1fnaGl9hhIX05t8FjjhJ/12XzNWrOwderBEPPKx5QpR/
7ERQ1fTJ8ngDVnMDEYmEEO9ZCIC+O0TY0s09dinHwXvFyK7hMY1vQdNUQvE+KErU
k/AD1YuBM/vYRDyqHU0zzSNtXkkEZ54PJdbD5S4PtXHpjl1X4kuIqCK/TpWRObWQ
uVF8SFXneNqFxTBb2saUjasfnKfL4Z2h7KOyvnx8OvUiPn3NbHQ2DrrpWpMBfnxJ
sSjofgNGnll4JNKkJuBjMvma09PpfuyLZITBehCKB0m0r1BJd7HtDHYzteIKPWK/
agbvPm1C4bTdSZXNVif7mFQu2VfyaS3F4nZ8ARYYXHQ85KUbHKu8A7xQ1Q6J9UBg
uCa+tGk6SoW4y7nb8e6dOzOM/2VSk7n1ivKQ/V7mX3Tm+4xwAusJOto/I+XygZRD
1I1DiZ//wJKTUhSwJF92JFxB2oiVxSf3RLkcR+rz2ONzXo7Y0n25YeTmwCWgRAmH
fPcEi/EmDcqsgjah/QK1MdUDJNqzxXbMmDH6Ak1wBXwAcVf4F/2F8BbLHoYwzAVb
3ZZyvn6W5uEgZwhm9tSzS2R6rM5QQ6S2WH9F3Pfv4b965x920Hx6OkQJ1YhviWNf
qR98WE7YyqEoz2BiBlnGQDfdZ6GQDGrNNNW9dyuHzmvDUBmB72qBNoydKaVOxe3f
Lb67/i4KQ3qBxPJ+X3MMGwq2kHL6z1Ev7zVkqGE52mRHZp3S+Yz+jGZbvsHLobHG
WeImWstoVU8lfRuo970ntRerLfySqu8qL+AxKDYCLFHY03m6oR+z6b+JnpoiKpl8
dSIOx/k8c1E/Mq3+jdiYHMflV+DMf9gAdonudvb9gqKa/Cano2FsmW1Apc5eFral
/bvL8TtWZNkqYTdaz27+dq3c0xOjmSB7qwdu/rjXqh5iQtPYNXndyWdArWahp1VW
czNqLbFcLbsLuRtPBxkvsM0WHlNhtJJNdLHVAzzCIERzHD0lzchlmXv/T7gmPVJo
MtvS88LCR8Z1aVsifDnTxKfKalpAPeHN3s396JRSvBUQEuuaM+VF46gqXJwO4qAP
p7xzD2E1CqEh5XVXMkttLw6SpoEodSQqqixmY4NID5VeLutlXvB0J9fajGcsYGRW
2hz9p7R8Bd5POTweHTcnFF5VaqDzWEI8mEtWIFarxCRovUosmutRCK7Sz9DSJ7mY
yyIymuVAbAXx5yEZmpOYrJw4cmrdxsCx7EcM3OjskSALK477vfQ8QPy7ZuwdhQpe
EJyem+zSbXvcjgqci5RdcaUEfuOHMPvaxptGdQ/rfhR0ofTkUaDIyi5NDgYG45qU
DuEHvHCMlxxIhbhjf9K3gj5H57QA0FAOlxH4xckzXkFuwWU6cwIGvBN7Ohb4ZNCa
x8HSNVvMR9bFVKmtCkxfREflPgvpXjz1ej5fBVQq/zARyYD7Mt+qWqEaJHMwwkmg
LAh9Z7gtQkQusFWg45n0nZKQzy7oF8mrOGHvs++5iPU+X7gc+9nMG+j7MJCHBztY
xyS4jUZwdBKsl7jEj2Cph/UvYcLTLfAFIaZ5BswfvVMeJaBJis4ZT1BNFA+V5Wnb
sXdqgVCYnyIIlUhTXh4ARk+r7p5pYR7R3Pi3SP5zK1D7/IXKfwaNv6bllB3p2lY4
bhXYwerXepGgWjdRUBS2c9K6Nk7RKx1yuNdeDjtSqzNiOb76+Z/b10Eh0be91J/M
mDW5qBt5oKZOWe6LMVoXH2eqei2ft3oFXRqtaNGaxUpstFJ7HTNivmK/ydFnwwHf
Kr9d9YN0zeZgn+vRDdetNof/suQWCTuIEIShVyQLvT0zPXHZ+5uTB04wyp7SWT9D
cCun+oYlGsvLFB4VqCLPq86qHjtPxkRacmDOTl4Uvyayw2nnpEVvfzOrjM5OHfQw
FUr38h8nxHosVdcugGwWONbpj8RWhJDv1KlYNDXxd7E7f008u4CxZBF/Ar8+HIaH
vX8fCTRgE0JfuyXQpY5gDQ+vZRn4fVc8hxXX0pnt6mXKaBv0yQNzPHV+lOSHPP+k
0JAPowVuRd1uXW1wrTORp3lJCU94KrN8Sria1xSm0KVQgrJgiAVbcdvg6m61vkBO
llgeXLu5DiRfN8dfZ90sCm5EOOgjpXQdrXu1OR4q7E6TVC5Rocd+LY4RlKveBkPU
Yts/GQQaomGH7+2G0KlB+99nVKEaKNlV90+Bor2QFK2dYCHYBgM4Y7yrRUE2VJbJ
KLsG2e1qWQ3E48Sy2MoZ/2wF57qTLYRih62oXW3otAdu8E665xgJq/hELOC+BYtq
nrM2mOXJ03KN8Wdkb/wKLthW696emBHjTW2UUhBIGYJo42vzWJGOP3VGGo3ysnL6
gLHz6ipl23IP6dBCtWzO2j/P5dXKeo90EvTZPbzyE5wJIIlFG9oHgOo13TJKobm0
NsHdsna1wWGU1idzM4mErsburUhf9nfJCHjagiP39vLEOAH1Cm8buiQcozOJXGFM
BCXtEBHaW6+kGnjR7G1b+9C7afkKeQIWDhiTxsg0X1m34YkIpLVbQzUc29QJvB8L
fQje5VLskb05BCN8MiRmOL4CTt+z9fNsDIM/tBTfi0FvHb1xRaKEEE3CFH/rbupC
j3/kK8xgVuYWxGF3z0M1y2NqtWu1X+KAcIUvLPRW7qmhTEH6Gq3tTHMT1VG+60y8
O4vmmhOgiH343bdTAj1JoLR99mA9eRQKShN6AjdNJNmgDLv4oN2V9Qa2Ulgpzkq2
VXL9aPcIrRi+9o+MQqQYhc+VefkB4NUx+2XA0M2PgizO7e/N8qey/BkZNEYdkzTB
tL9HoiS325+s+VeaLB6H07OCdizVNmQK0z+wf2ulP+RHQdsj5QCYWQ0sMyuqmUv9
6X4F/gc8A8G5SB2Z8wBed8/k7HbiEr5h1vF04LC63M/3PZ55aq2X6DyeCjO5InD6
FOhR8NG+tltNb3B/KpftubybCcsw2OWVSOfKYIrHy6TF0NZJhhmRihXO8wYT9kAp
SnoGWRRVCNbaVBK9dRCfWASu4z90EYReEHl3nPQcaldygAT62Gf54GiRjvIJrHos
R6O/x31FGTqUuksTpvscT0+R2bTzrxNkT7Xw2UIgQwtM7Bv9QTz16iLIE/ZFzaiT
imlCm3/isc2IMpKidu16bjQFpKE12TYWid6rgjs+zhGj77XX173kNArPz/tXwQ0N
904QSlo1esocdk9r206Oo4dXKLm4fBYlyLXjL6NnNBsEtC1wo6r1qQUYD6OBbFBJ
H4tCMGFY2VbPs9Cr5Jsl9DokXIJgdrLf5SVuI5AaIknctdlvP/P2rZOr2L0maeBr
jQ82Z8CVNFajAqDmEHh1yiiAcfJ+vYsQWrSnLDUJBMOgALICvWbiVZ80Ay8vdIs7
ZDdIVBe1jl/rybCjGo8rD+FT7+Mr9U8K5b7hJmTdULGJBlCs0+mSaGaeq0vASouF
ysje+wHVHOiRWd8dkNNW4wVHkTcUJNEL/99IhXzJyNzA3L6yBVLgZmOKx9r7nYcz
xQZ4hrM7loBU1BVza5uEWo5vRdC/PVMH14JCF/T+KYH/vKuERNpirp/4U9/+20j4
7Z0mGgvX6x8fQynbUVJfh9niDj9IyW5sRoAdkz+Dd9LjN4lldjqi3G9tfaMpYKmx
Nz5JKPo1A1D58O4I/4Bzb/llanMcIPKV5zZydwyennLxCXEGbp7s/oYCyfJbJhnt
S7fchBwH+12ClfcOdDAxO0UupyfT/TFUkyBIqtT71jRB68DqPxnhOAXBOEjlrTb0
lac5Mz6bpnixxrJvBw63YAzOaTMsi4CUM/8cksamWZJwfxzdHMHbdsa7H8EoJzaB
SXTjNzpPRy4jeO/bqOUmOnMT6z37DQBMQEqF+Uc1OsnvFoY5CtKPpVtV6iDH+58q
uGJs94yntAPkAoanr4RsISoDbz0jUxoyhUS68znGZO+HSuohyMnZAayYLc9H4Ulr
xLWW71Oa2LV30wtTgNb0dLQpCILpeX2TsPAUyF0/O06MHDdM4fTTrn9cBVEHtopa
Nr9BsuiKTbUlKm99gR1xFginNSascaswj3J0cDQcQ8gdYvp9x8enESj7vrZI3UQF
Y9LYsF7kEXIO+qUd+s/o7GgSlLOgeZp9nu3LrbGy4k24El0N7R2H5kwj+v85vLpG
RukOdyRL0/MJr8YHtNxL0FfSskMg9klJ4D9GWN+o94RpsBfzjQzK/DNsHmwPHQ1+
/doWWWRbuNTahuReK1O3WxqY762PwNuS2lZeMY9T9aOw/Cnb5i67BcwwpEp7msCc
HnfTJAIU6K9SdSwKcpU7ZnavdCqslncq8i2hMVl96ajqKqI/7lL4+tZDl0LIcukx
eZc3Wo12em/FMbsmvL/4KVnpMrZ2JI+3bWuZgvsFAH7pI9rwrmzwqvacthZv0u9S
e0aQ99BpdoIFgRaVKvl7eP7kZRw3/xCbEPVFhAH5Oz9kC+WWieA0i1kAYNeAmKcM
gp8TsfOKg5x7do16JA6DcsC+08azY1PChfLsytd7jSPGuT9V5SYTv5nAc1qkfH8d
TB5j6S6t1Mi3+PyUF5ZqfVV+K34J+bspiyVpU/lS2bLody10FnfWL0Puat13tO8P
KaXKeZEouD7wJTaXMmBWj3cuaXH7KPye1pOqOsidpzes+aBcynEV0MRKHg88nspB
5IvFQL+UbVAYmoJuhg4ZmfaGqBpF2KyEN6CNpNycLYT7Cre5vsZcQIARohxZSz/b
RshvKeRaCa8pfGb5x0j5b3GCSZLoNTFwLFJ/m+ozCwofSRdf1s75UFx2c81u/QkT
DLjq5WWUnCSDeOANFi9m1L1bQO9farERTCCFpC3DFy7nXekaW5LgAuWKqJnIDHrW
dwMoWlB2Xj/nLweWuDHtwNcuwq12cbqMSXwzRGD/fytGttv6579vj46uD9dRJnJd
waQqJ+1jggWKjfA5Pm56A8xUKaaQYoqE+1wDzTQtB3EJeHYahdRzOMNWp7bxXEj3
5fhiYHEpNjhUtU541QBvkyY4JtfwpsR9daOq9WrwTKlCfuVzfQJbWdOSJkYiPT32
XYOGv7rc+qvt+YdbfVhE1gVsyMHDQklTZPK7paWn1V5al5i4cZPQwbDnytWJNlrL
uMxUaH3ZB4YWOoMPduEe/OGt3c7Jw34QAGyl64UezyTMUsNtZK/4MhXkHftOUgPv
x2fCLCgE9D4HGmdN0aYSKaX/tLyVA0T6iJ8d7IVk1umIe2uxOUp4Tk+e1+mVUFx8
NTxcSFf1lb3u6ivfI2XrVJP5fJb8ntYJzjM5hDiX56ivN8W82wJeKDbG7A24oL35
UpBeYorlSs700cJDhj0pyG6G84FTkgzdYVBKsMX4qMMhS1yox6kMR+9FTmM6os8O
oo4bSKuE0vzZ4AYleULr7TtyYVfDrS3Riw+OPjRBCAPFnZi8/B2VDxpFR+Fbcn61
7uOBEP6oJAn28R3s1f261ZADyBIzsXCE6AxMESwkvrChn6e9LuIxl2qixJELlW2n
XulA5CMQ9UjIw9qUCfhJlzo6+ps7mWC3apFYJyfqxiUmXxMxU10mTHvoy7dx24JK
k27x3ZibOehwiOerfMBFjICCK5IH53rF0Pnz0mhqJwUCFDCQYqPGluzi3osciIrp
3GxL4ckxD+WTFQkDRKk1S6WQ9B5IaWA1x2CAi96S3D8IsrfQZVEmvdzrR+isWXMp
FCOba3doJdH3oLvGGt/ulixtxV/I6VTh/R7pRZod00h34xErQ/Ih5HOLuKAaZVVe
NT/941gD4MCP+N2MxpQwq7LParPZzKqQqlqaKJHgmUXmyr0yvfUCdEFi4rA1TKKA
lMruUP4k77eHqkha8ZdFEmxwArQtaIj0NLOS+kbz2wux8+EiSE5zQ6Wnh0qMQFBu
GdC7Vlwq0/eaHLrxgRzVXqDUaulwFV6eFchTDyreyjphNEEi5H+ss6nyRixuLOpk
KbesJ5uZmk82Lc1bOY9xi3qWhYxX7f6nHhTAtJO82CalAcQ82qk5/yn0XAXBGJmM
9ycnA+vVfWE2nvnurXMjcOcEQQ9qi5Q/4AJhrizhDPDBPZovfUnWOzOTAExUBeGh
MoyIgAnVJB81/TMZAk/fgAdLNZTIoQceKfKlFlk7IZ9/5u/oH0xG0oTXitMapL0B
pB9lnbhUqzFEAxZnSM5WpWHVZR8WT3JQ7ScOAmeB2akCEVVa1V+GBk5JnATDtCp+
EnzbQZLAdc/1hypfO5/xXn2gTWJzCwWjNm7S60U1ZErkI8ywQNC2OJAlUUYvkMsW
RQoxDTE66sA+Q5AiTtfoN6J8EpRzF4EFKofr2wSTWAWYbFNumrB8VyBA2uBoRGG0
moQk+rhqO2hq6YA6VF4j4lpc4V5UcM864TD9ETjwvthw8uoOI8OG7W/QqPIxgKYJ
QdqeH5R44pVqtHPndCokuOCnZ99umGBLqxAtqj161pb8MVMGgHveu2EX8z6mBins
n/vaJIOf9ySR6YbPBGcuoCJ1zZXlySj4/2s0lAW4451Yng64DWZuKSfDrsKjqH/u
cIDKmPBMGWz+Mz0dRIGYWrSabOCwM0fFYNxkHHtc4b6IoTAnvqEg+bHWsY2Dr2i1
R9fArW847N3JV0YfrEGvwi8p3yguWKJBna2kr+v0k4tD+NN0fZrk0ZLKjSCTTVdP
FvyakdhkhIpxTZYx03I6Zla9DS5buvIsXPwhEa9hax0kIYvqHWOESrrpPfvBoIHs
DSOdWxMYKeXS5g7S1937Yw4+JKcmAwhfbjTVRp6w5DYsPKs3wtYc8CDf8bz/cDks
lDKj2aqXI4PnNQNKVGUBoE8CdgxqWcNNuXVsbogon4EtNpdZQXqoSW2oo8gp3MWN
+sVajTHvm3FHHkb7Bno4avPEEqRAL2+djKLnrtIZnQiub/4319d6MUi1L41hj24n
7yhbl5Ls9w/o0NKVWHbxxORaa97ylYdGQXJmWW7bglsVKa5dWlJi7cddMHQ5etKM
sQwmTksrzJ52/d0uOQt0awtqkxeFzHkUuvG4SQnYS72m08uLgXUFAW83G66yxhtW
HzXbWeQtBUWqVOR4jNXICshnw+ihWNHuuEBvyNcP9NJ7alMqRiD5TOEa9oK9sh7v
vKqg4k5JkboEHQ0675OuFHyHvA414NO3tQ9Y5TeyNglzv0TEDXkjDpngq25C3Ppx
1fRnG/OCqJjN66nFJXo+Pwq+1iNH6pi5op+7php0IdJU8A4YVY2VU9YuAqNe/vzg
HijD0H90jLcAjYoOZl01t0hhri4baSAmpJZkOz2P2XP33k1Pp0FoWaW0HkQASEPj
PsXUf4ugotGgyDEIP/fp7JInADwuRpdbMlfdk4A52/PmhJA3rgbF11Bdg96YBqN5
CqZEbBVPHgBa04qGFsVfhTauDP2Ylm9KeHet4LF02Mo5y0/We9nAfTnSEn2ny342
j+wUAJxZwP7KLMty2jG1deLo68KihWL+Y0etf6wgI0LyIFyLWbRjxxJgsFeZHTDW
KPOljFQw+fccik9va6tKfjWE+kHFzCejpzJ5DCT06BpgXP3nBC8OapkqIO7pBKeV
KyFOp5Y/r1j0In8UQrLFd74iAq6k+PbmSa28X618AcxaK75LJkFQTkcbZBUNcuTx
w7Bz0V21VG7pnrBZ8Xu0SkvYGfxXoNvLR9aixXbXOtB4qw+ExbSEELgHuWlRgTqt
4QMyF0zFOK3GKaY2kMjXITv+gwf/FdKaWuwhHvUzoNS9VseayfUFQcKDJ/iN5zDG
kx6XrBNncNPPFgTqwALxoajEbTn9OfeofEjrJouyha3/2MCKjthjHzeI0nPnE/8p
F2Q3vGpe8ofI777nsKlmp3QfET488YO5yOoyl9g2Q927Ble3srx0as40RPpUNnyy
JoxG//zPrv51+QZtZ1qU8wkgcSD+MCQz27sHLwTTPA+Qi7ljzDSwHg/BydwyRKcZ
zpXQB5pF13llNIeMS5MWGuq4bd/OffZQqz7GatrhlTwP/EQ1V76tk809HMiSDBh4
CzE0aRAm1ZdXrg7xidSUcrnCJvxQHBK0YWiUsv0dIVEkusjBmy0p84kfO0K9fBYp
hYNt/3Nzqg88KJq3VEXUhc4k+EE/IjdChJ9eh8fpB70p3LTAv0Mq9RTTMyXIVFrZ
4wI9NLKO4W5r90IyuJvjEjKQqvAqsMLSbKCe/VXHEqw1xW7m4/2J7VAWbZ6IcLsF
G1dGvVg4JlO89WsGtjKkB8RpVRuNDce5C/TjFvRQMfPTSqFqpk2Q7x4elg4xTyMr
9hlgPChFUFWksuiyTE2/zaH3LRoVOKmP3lDgAft2KBQ1Y/v9le4qfYm+xb7wxKy7
FmfCTQQyFrK+oDGXGp0LwRjzrDsxzOj+ctEFuY6z6QDxavN8OtrNuYTVm/egrdgQ
FoMHg1r7rizOxt0IKYlBSUSzpLbALcG1AwbkiWfmbkmNH6tVnqemWQms4D+yDnWV
FJ9rWMB5b0i8py2bDJRMcIre0HHijeJIrJj4MMvF1Fqmh4SWbhEWbWMzx9Tm+Efd
ibySaKWBjZRLyW2TDDk/l+TE06S16qX8hw4j0PO776mjEgPnxo/YtmEghIbqKynl
wa9RBRVafK6N4cY+u984GFHD9r+JzjdY5gZZWKlktaZTprfQuGLAOy76Erbmir/p
cWGPwzkkYJRf/AxfYy0VPWzD2k59NzC5Xph+IUe7EUNSy8hkvWDJsYRcju/Me6JD
T20Lac6FH6VrUJ3UHe72HAFNWAiwo9heCuDcrsRvhM90cpCThsEILysKziRo/F9t
CD+2pJKvXp1E7m3jZ3qP2altwJV94fH7LzrpWeNs/KwAEDkzQ/VsVY3jlYK1QJQl
wzH49iOuaYtFxQf/PROR85EhnL8VcPcy26I+iGj+eEnsNoFspqK3YPPeTLLXtQfd
zRd6TW9WbACY9iP4BmsxLWSInwYefwPpMsTfJj2APyuLcr73CdT0wTMo9p6U9P4B
LLqx1Eu2G++2Ca+tke2Ag0ZPBdeS1apSsfWFmzN65hlbYt4Hj2aYrV+ZyBPRa5nj
c7JGQrLCm8BS3WOTxPUjphSoGqssdgaelOdDMfa2alK1yXvrp1rN2JnYC6wu+wP0
Zsd1Fy36E+nX6TAnaYsXnU8oW8IWNtxy/FI6ao5F1Jfu0iiF5mi6/E2gd+7wV46a
g1nh2okjIi9BD+IMr38bIkJAmjGBnBeuahBvaiE7J9lf7WWwYLuSJukrS6Mj9h2v
2dTlgdcSciOuBNzWZHq0nbYFZNaQJLS/eVO3yoKZnvwm6Bn9onsoEsd6DzR1em8c
rPoElqS8tOPP+rsYrWpA+G94RFKD36/MujMU5SXqcOFedpQ6XQsy31HfmvwZena/
CgodArSoMRU/wu/FdYUXP+chwpgf7XC/bLzUpZer0H5pMiCuHKVHvqiTNbhBwgmk
cHvfGX94tSm+44iw5EMWbI8YIMsnMrlrwOU5HB8zPZND23hLIUHWDd+x38szdr0a
3FT9I/j52vEE63BPzpqd6cczNGBM+wK+m8B4pJtCnrC7eZdFAOcMVdtzOF5O5fRT
aopea/Ljv5rH47k0ul4VYsuYqQohUfmx3iOG6WJvki8xynM8btCpzQxlyxUAI2zc
23sgKZQ6JVRwuwuN2c30I5JGX9BwEXd7QOuH9AGEPPT/KJ/eX3/vvx3tmW6sWx/i
0qfwBDeXeq7l30YVJNXkmcPpNVc9PhN+mR0eOVkMaxjl/4iHnEmlr99R5nqq39qn
/RvkFT/qcZ0HfLg6b3wiVunu3rw0lU7UBrM5G3RBD4xdIVoZYrmabx3OLKvH+izP
cBMAp4+mc00OeE8YW7R+KRk/JXJ3V9tIIut0NP3U2sBXGifZV6om5ZpWQNq9qast
FQ5zh/x143zLg5SM6YGdiy78+Aif3vnuZU9fqu3e2jrRokROTqTuLO2yKxfCAaRG
XTg3/tQOxrJt+RAXvIOwNVM3DyQ1dvyuOVzW9LlI6By2MzXMfR7saxn2jWkoEYaG
Equwgt/CLgECUmrE/gJ5Taz1I4v1K0LJSKRBJebgRcXG4VjPiFrFxkHRXDRHHt0i
gk1kUCdi2Rd3nVBLMTQfH7C4qRsH81168/VRTMHldDILM1d9qoVuEKUMwvb+j4+a
vnw4HikCbPMFqG3c69jTZ/9MzEC5brWbhUQ0vaO6PZd8ZSGoidwNg2ToqNnUtZac
/3WVy908fG+/RLgNAf+MwPKDBA5ERq9Fb1mnN9RKj4inqB3bmvd+sS1YKQ6WpjgY
H78ZoceocAQOlcw6fum6jCySiywiSkYb9L44m9ULUZrwduTGBw08TWOOASWvaRWI
jSD5SI+IIKc+X3c3GUe5aYyasV0Igqtb9sSgAr970WjE9KO363tT0xO9FYPIXzoY
4alVuRHhpUVOJ7k078ND7Ji3nzk0PcXm2khKNoyWs/Wl1u/9PEHK6VlpST9SKeOb
IvcZLidxbfw61DPr66LL1Y/+uGRlVVgbrjqI21c6cc2odmHrAR5ozVFiesR+dl4c
EdMojeajQdKe7Z+ztEhPw0k0QH02ZNB/kbC8lD10nUju0RlLi3+/9axqP9NBBUZg
i0cM6ez2IBUkC0T1r1tpnVo1l9SK9InXiplqmjoDTdC1RAuPdppoUtlWs8rJblGy
AP5sCnYFHGV4qhIYCUVkDreKugoRdA4Jg+aqUzpetPkGDWJCdvOlkZ/Ho9XiK8wS
ymXipsicY3RWbM2zidvwTphn5zHt4x0RGOMpNQ4uL1sbfw1eO35BdhkHt+ZOA5Te
q35SJBreGC+QJc0bVI8tj0dD5belzG5jEoeywYt1/o8j36JFdd6KuyLsfE3hs8AI
YiwQpcLXNy0SNdLz3p+KNRNIXtz+O8v/Vyweom4joUaCTbJPEfiKb+XSQLJz2Cih
ABAp3sypl7lmyTIO4Lrh923nax1r2PSgbF4i/ivaAaDz3zuvL2belAwfxcD8O29D
tIVKaC/msPG8fxLgvnCpG7lnaI5pN8iBQdKrwzXHki0axE95FtmswhLt2OaaiI5W
XeJpOZYFj5PbU6GAjaDs6rJxYL2GUFYMOaDw0rwqKxiDeaJI/sIyaB821D0p42ds
9JMgw9GtbD0RPLtWRN9N959aV809xhXj711KzSIMHGFymbzAZZ2jDzOue/rjxftu
VFKEz6OZPd8XBql1NXIMzFYpR04SHVzanKtQ9DTQ1QEMzuOwREZjHT843hz4Ll0e
kUSIJ67kjEZh9cOOfUTXaTQOaw1r22Mv0qzekp5PUC1lxNMCuUtZms1qq1qscKn7
n25EHMqsXRT27RWYnDVBKnUMvx4izasIcvf+9fRd/Sc9MZ4dRuXaIBJBA0YKy0y2
zI/BUbyZkMlVscfThQTbrc46U5ZzHp5cxd02NYljZ+PMHBwdhW0ANt0nZDmCWYo2
qmsJ+VO8R4hqfRMW2uzv3QbVutGCirlSn9j1iuwfaAtm3Iayb/8HdtodZ0Y30uF/
YOyXam34WTeIuvJ0OYyUPrx4Sd7c0RoPIgAvGB1Fj07alcr1XkGnxIr/RTrMDRif
fBMvWZG8a8abhlT0mbVXxdU/zLeuZpNbrgX9aWiAqKxQ/nxIQQ/BkTDhkfj2Vecp
7Zd4vquHkVXpFjIAUKYorJg4IeprRBMlq92i9380sfgKEBA+qsWFaP/hMbkEWYo9
1aSnEq8BI2LM0Lny5LH/Oi0D2KlrmQjJeNFXhQpBgCkZFzOOu9cTcrVgM3jZMlLy
VDYww6t/C5tZYAOnMSxSP33+RCzAimXhI+RmYHvekVbpqoJJ74rnYhmNGQLhBaH2
wLhLSMoflGxi9MSGiLKSvT9SHXmt0LbcwTdX9hx+n+7WB4rwjAi0RxRk32FHsWrn
wx3jtTh9wI8kKI2A41pAo/dfM1EORbigsQ+XZI7sI+o/IuqHb/n7JjQWPJVk/iyL
L+Unr11ACdSxbM0XinQQWCp19eD3ozgicH9PcajGRjI5P1u1Xyi7oAspDaYwZkm7
DmPQPejVYM6s6ekSqsswQPXj1duCtecQUKBxHpYbVrXMZDSh9vUSMKuDunwUSkRR
PcsHsK5IUIkabRAVlr7dkZnSdRzk00FKPi+WsmzJI3FpQxobbubgHhUbmCwkOjoH
T2iObxTe4ZO0s3AbXHR4ob8tvoC2Q9dCqBRj0nVIBcDKKuhgmZkwLTrs/UsHZqAH
e0gn6+ASEbgq7RE0qnUjPWSTxnVw9yCoqC0DKzbiRRYccfzyWwcAJIB5A+ndlyl5
L3dcnso+KhO3JDZMtPTVpgdFNFDNu5lN4atImJhJfT+MU2kf+2nAFWAgjBiaiJ4/
YbnqATbwZccNHgNOoQGktd7Tl3hfU+RdKkMnDe+Y0zi8/tCi1aBkT1nMKwGawm98
Bxo1/IXwSbYmUy/3POTM6Th0Zk8lUkciJqBdhxAlAfsyNXERE4WoUleEfXP4WhMu
5VJfeNICul3W2Tc4OOHwEzHVo0c0jxSo+Xu1qPdgDrw35AseuLUXAUluw4MrJ7fq
AevAhmBUWepjbszLKm0dxqnb5UCZG95dINFr5mDmk9viLnHN8bSKysBmGpwAIoeE
0tKEDbNs2wLzkXXhgN/a5YfA3VP/uSsiWlGlLPUo6Z/5raiqxuRyYUoiTQL+MukG
EqJd3VVhTlsvCA3+HsnDYP0AwW8t5g0Iywejk+lNUyu9hqhGn+XfAkWYG8tMwsPz
0EdVqzd10RgClnxoa3eaU4skn5xETWhzbMUd5xAVKKO98Kfyo8k0JnmrPRP4X8dh
18WECWQ+VVAygRL0Unmp6Bels1SUWqZu5hTar+sQRbWBP6TmHFsbm+rdXY9gOF8x
/bZ2gkae/CyZN88tf33jqye5xltnLGitpCXLfSBFmownGnAsQEyfaiQcGinDWq11
8ObfaF60s8QqsZVCOC2DPwaiDegDkiPjuKMVy11K4BEjpxcdUO7blzEiIM3zJ2Ba
oTjk0LnBKgPUx+juU0E3LTlmwjLz5rrp8LCM3kXRQ2/se9ZBkL0wjdD+Wp1O61ao
WUD0WWxpUGRqOgCtapsKPiAWWlSnT6QrT2QkmXgnD06ifPL9hl4dR1RXtb3riCkA
7zI3hA0TBQYqkD9hhjPDm4MM8sULOQyOMzueYNE2N5skuyWkjwhiHWeZi+5K+n57
+3M4CLiWfNAUncycLhCvB8yIjmLROzvrutZ9qk/tZPVrFoL7tEpfwrfh8Ooydjrg
YwX/P/6C6t2u+mcWH20bEY3hl3LYlO7IBT+5ecw1MNyhpP9amOVeftVlHKXQPnLz
7WSTQu9hdGIu5x0h3cSnF+UsuMtQJ9VGDVVPGVMFEtyQtDYjn4NKtq7zumqRe7by
SnTeNwVbHQZCaXd1jI9OLnTHdPxly+ahGN8nunxIQmSHcrem6VQyvf/hoa6dV019
Dbc7ZQnERqVMQ8yAVO53Uvlo61e47OfPo54oucDTTWe7N7EXctR3HmTNwWehNOtJ
a6DvoUl3t64O49rlZz7mg+dRcer+XSI6OR4CtK54K6AXgYqwxIvm/meUJ21kAqAe
jVWNnTiMho9X1jeGXVkN7wukcU29AaKqpevE7OWxq/bLOY3L/m2WMCafBUBvUBjk
Oz8+5bApCcda/Jx22FOg+9o/FjV6aPIb6X/x0N2IAIwB6lQ2AUvnKKbuGq3qylw7
1Ch9NyXBSLQRbOJDK6EH7e/kRZATRjufIYk9gHBdmwTfRQVM3iz57CAFoI+icESF
n8XDYHQ3QCiN9NyOd/ifIvOJ7Yd3ZnMROz6dxoIQ9+UlB1aY7mBCYs+q2U/slgrJ
Oz4Gf9j0Alws5c8EFvXAYwAhfPoR5nByQeXf+s1SPhSolZelPakh4qw1BYHoV2AG
pzgqBZprnnVF2lZSOSblXezb2Sjfo9Jkwhahkoef/zFEEoGDbhmLOALRArb5fa+1
EW4Lzj39DOzK3LppedZT5UyP2E6pYbL6UJWUvyQChVphnoTifpglA9dO9/fTKO+v
bpF4MUxUWcEmrnIG8vLimWkWGkYWsIu1cE9PPIjIYGByOb9oBIMtNHccFExyIZYo
vZ0F61Tw7PW0sPSZKRQHqMYUus6q4Lqz8havieBpJ7LWSEKGAEDEf160couP1uyf
AB85ouro2f6WH+lqLQ3u3GcJNrSQ4Fg1dljA10xltnj26UfbmIltoIMrF+s7VRin
+Va3sJC2RhgQ5uf/tmigyuDwGY5tT3kgyI1hsUv2RyzUT/K78LDvFqYa0JGKD+U4
pKHhnLPhtsOLCK40LFqSizUngzkJ8LQqeOt7fgHMqiVDjXW7IKZ9Xvz2Z1r/Cbo8
noGTjaH0PL51zvv9mGHZ2KXhRk+AlKjR3nedwDi+cU2xNClFc+aYW/QwsIX+K5rO
RG6exyIIyLURwe7Pah4B0/bOyDnRrQZ1hbQHBU4kCBiohWijca+3IIrSg/eEadE6
apFU6ZIFFuPl76sGtHsn33p4HqmrpTCQwepKpWD2i24FHCoNCHKVfnt7En+2z2rU
Yao8BC88zxiCoTWx0kXIhOJquDH11bM/uhrub6lQx5NUj02vBbl+gKopRutoR+nV
p3ua9VFgYBsLwQKAMHv+rR3VbO52p0zYeBJMpuaXWVPsvkRU2nQgk/q5ssa89Val
1f8iYy3fcSVPe3kXb1lrqEn2UuYTHg6RII+Dl0VKdBmqqhtFAWos5P0SbWjNFt3K
YEdw8KGZp6prsLo0p4KV9nvTId2ENudstsMLMoCUGXgpisNxu8taHwsvmUZMUoxp
BmJS2IOPW12VVkXl2eulQjmvyZamrvP1LBqnEaZc/i8CrGNqbkhRh1M7ShQ80lLp
odB9/PpilHSuHjGaY0pg9sJbXNQrtkXngKq9KYF5qKkjp2edLLXlRxGwvsM0ruO2
Ib5h0YR/73eSI07Uwhe0X5/wF7MX7xyBrYOh3HqYkyyBRzmoL/PpHZtznyot06/n
xt5BgjVqEanNayusvadsSSw0OONX1vzR9K8agJ/5UifMMNP/J5+b8sEgHUgdORxs
QiKdGu0iOIbVh5iRERifM9+zu7KiLcX3nIGJfDRW5AfLGnMZtDFW9bQt3HmnupWn
Sk8+lGI7zqMJJ7Ix97N65+3WzQZuK6TRYFbun9NPPPz/ZOZeutKz256DlzyD/wXv
80Ddnck85ggToHRnIEdXeMK2qI0V2HFUz5kexhpHk6LBOzUm2HKsqtLQsXXGRcyw
sJal0uIyWC+wA/0+/3qtHATU1NYgjWbpnubP599or1jguXZSp25ypV35kQVh60kf
Xc7O7mB1/xx5Nr1ZrdPti81aPsBmOhHix336Zgt5EgAQj3HuOo3X6An25WitXSQN
rH/g3t1luF9AransLkLRFEX5eyvlmmwpH2bCb0T4xN0Q+QQD915xmihtMG5/kQTX
OQF4OWH6RWKtxWEvQpw4uolQKMfhKviye0zF50vTVqbbixSAELItV+qoxwKD+uWg
1T3pc8Of4tBAQRwD+JIjlrdltR9Omx7ENBDA+5R8JPuunYDOubnM1K0PUuIgF7cS
cgj++pPRLTrRbxVo6XjB9XInFb3QSZX/RoOndMIiVvMT+LxrZ/JLVldG1NpFk1RM
tyE2w2NvjMEDC5qmfXNCPjoGHMlQ7t3QnKL08Xqchn1IWUJJLAiZlIH7bT/RwLXS
dWbMk4UV1db8LLPjLWe7TDqac1TbiUR/qICnBXZdybnHO46uab49047gfZy7fR6V
wMLzpczMOmvVJF79lwaQHxIwtjCKdWXEx7hqj9bWoZRcE9VYMrcAtcA5/FaZnEMO
duKhdg+Y+LWBCaHHJfrtMgvYCkTl3Ols5ZEkOih4ck8hB1uMbALcpgqmYOQ/Xj36
/dTu64bZB05xSe/YglNe9E/pNhJ1crwPw9L4/qUxyGMNwNplnLhf9h1MgnnhgWeb
OVmB2r+wkmimOUlbVqdZ9S4fK9/jsp+YILCm/bP8zsXIcoFBUbp+zo7Wi59F1Pa4
dgmz6kehqRgKne8LRxGHferogl2epLSuJVhUfxHexfUSttn436GNV1NUlO4gvxXs
gI66dthrNl3oGKs2YsvVPADFXSFJDRLEf1i4ZHu369I2qC/xjhDw3wd+Nt/4+lFG
3LgoK7eTgOHQOb449/S+XpgBDdvCfwE54iKOV1wJteqOWFUDSpmotV8oYqTPsfzh
3TAeNJcu04JbG2Qhf9qp1uY8IH3gGIyqQxFNu2lke+JBWzx8pV3YlcQ8Mcxd0Esz
K1G+LpKLRGTLjoReIWbGbmLYP8sre/RVVUkwk2w5bMgjyRgtoe8CaM7a5dfFI9XE
dcLvQe7aj0xpBokNPdOjVq2YaOWOQFnyumqWn+isyswrEUDrNBEBjOWJEE1yRB6+
nIoFYOtHPgg0NP0yg8YVQ+a2/A9ClpNyXc7qxdwdfoLIohmA7moJLgpc064mEU3T
BwhCeRge5rPP86gIn6OT0KW07KbYzmcL6Ovys3EzpsBo9gYJ8Ch+/VWqJuhHF0mF
zHVygTEyiSmyEcjLy8APqyvIujL6lchnZSBXBjodjz/ODFsPCooJS8oN15tdSX43
UnefqpUs2d7tjmrAPK0+R+tnG6Y1P/+lnjcY6Pfiv7EWbf1Lto2IqdYnBOdqOVXY
ETGYrr0ElidDdq74BdXQTDHS26Yc9EimyBXQ5UOqBhuU37D37rkkb3DsY/Pe9g1M
EkaK4j0dCLUn8sdzZSHEr/hAj82mLo9DisHYXgTwXkFAWD2FxBK18goE2kxfB/1s
IE7ip5md8F79tHV4/1PjDHGvTV+MNMElgPzvKtvxb16bGQkMmWULL5wOOZsjc3Fw
PlbS4YFSqz+o+lGDjy1bJ4325poUoA8mZJNaaaJRyp6u3xl700Z90EdLz0eFBaCo
r8nimZHvFzX9VTQ98yKgs0iIL4LctEOUh1baHPqkkDdh0Y7p9X9yJZjPWNWgCol6
rzdimt4E3WQNFJJ9YYASdVtQJXOA0g+XVmd0JvHE12XfDSz+jNpuV1KRhoJdEveT
9Qx56k2EZrLGc/Cv4UfmlhnBd5nvMRWuxeUrohg0s4xa+wCIJtImynXR/fgJxG49
PZa0qkkVEBWHLevEmdZ5q1cqXCqmJL8pEcnyF1urO7JlYczVR5UbW3jtG07aZvrK
zTMdAEMkoyTZYbpnH44AAz8vMaDS4AVOdGbXYWJwfS+mTl4Fu9ndIZ2EbaNbHs08
fbFF/0sTbdOgobDFRGzuoOgPPNHBSTEARppFwoRlZ20UNHho58EsITOjiHRLRFDx
eXsF8yO+ixH19HEbke4aDWcOx6lnsabIXOfu152KcAoUCN1hLWZiMLhYHnLykrCD
v92krKQSRKjxTEu3WcYivAGRW/qmA57jp2Hk+j05Yer0d/uudrO/pAgCeG7HTWQX
REGJl85maOGhMF3V2t3Y/N4a5wT4EgDH34LjQn32mHBevG73aOQHzTrORODtwCBH
JP2bIuljh7NhohAuFjcjbrsz/CFXeJeidXzPZBYhWW2AU7w/66g8QkXvBNPxhhbD
GilnRXrM3zb9ABeFZXvZocbXQwmKUQw1pe3PaN/Uon7NFNyF1LiS7xrPExofDwRH
v5Jvc2SYOQr8fM0I2YZcfKhgEWxA2a6l5VIiN4PFfzwoScXsHDDg2kEtgxYqInCq
+DiUQZ7klCq3M22/InP3MlwErN5GXlGSely/85zgq9J5Khv0fr3mB/40dQYBoYlO
eVKqRtHrptDS6gEgMocvcNJuziFvH+SdJjsRtXRkzdxPcQ1V4GLv1S33VgM+ecTO
v+sqwMUBGG0ou6njDNboHIPq6ikJTGGn+SihCaFUq/432cE4sF7R5kVracsxbS2F
Lco1TDggn4OXvm3FCuGnjmKB1VBI5gRHv1nLfG2defbTXtbegPCmaW7NjJ7tcUQb
tO3WnY5jF0TuYChBsFJ2uQTmLnQp7wTsnY7Vr5MQMWoRxr/e/DjAnxndwBGF7yOU
ZIbOlou1FZYLYW8p9K4htLyh2VsHlxWL9XtZMquk5Rr+c6xUAHzTAEum2t7fnPsS
29wbTLm73ZhWkt2dnG2iSmMv0AAiqyqPm4GrXEqSkxeFUKV99n+IXE0kDHzQjc3W
bfVywRg80aCeMsMGAQcAsyrsvKN9MMSUf7bNn3P8kF1ar14qir26AoTgdJhtiekD
MkVPqYEX7Bf6jXNIr2l4rrT03+MZ646jwcAMWF/JoCOWEM4dwlnVv8G0iekNTYBf
MLwz9NXgAvwJ3/Z8EdaLDF9fyUr2QV4oTntJh70Gt+ZmTvL+OLkhkiDR+RSI2zyq
kqj2D/vbxV06CpLS+jhzgmWZGxbCZkYBFAdLMNUVr92/CtMXrO0QAlBbnXNp77Cw
d2pfUBvYQ+9YqTRSH8SqJt6rSRMNmFeReYfcbfZXNGnPdCgCNrK2ag874GUbMtr8
LKSAvzLxJcpZ6bT0dXt90pTzOU1mqTcgyGhf4IPbYZUKpTzp0XVyGJhyuuGNy/KO
PzulSxf7oVwADggCl8Wv29V7hzQoSa7aDQ/8VJpEbisqX10LS5bKyMSxnibozvJA
sdIMyCEY7uzhXp6gTSJ0coTdrF8YjqxriehY2Q3wArsCXnuBIvAIsFiFc/oMdR/G
AY99N9z6954Hz6WfynX29TR+ztlJe5OQghMQ0eKDCa9gL/O1CWCRd2gKkBao1toZ
4kS5MebqZmVl60UJXiAk68ikoQUh7VrCCanBKoSXNrJjzfLiE/GPFXgsudghiNPT
6moaKp5dlYXtFUb7fDTivjlEHrn8dtoY/PD1cBrE4H2CXB2J1YckvFJH+r6q1wQg
MD5Qjalb6A44Ef8tR05ft6kLQAbH7LUV9CdWpBSNq/jZ1Lku07ZXRG2VuRYrrwZ/
OPLNNgSmMsi0C73+aJA5VH/I8j9bJDV+4TWFCYuDDgV4LYnhollsIZsi0kQKfBZx
NjNB1YTMWs0+k+2+mQ0ehcu5TJkaM6c6vxwFUAMqzNSEddkIdIQelf4/C8BF5SfE
PvxzVDBAF1Fal+M6MCC0Kcbo5WVsJF7/E5qCWLBI6IuH0u0YkAwMhl0z8667qtbq
ia5wWa5mQJtGBlwwSuKMzOthnlm8T4U5FlIp1e3pP1KJjz73EzUruEM63i5Rdi2u
U/kahjOmr/J2oo+DWRspIUCvJhxYyaTfZ75e5n+s3Hm/wN8oeNNjKspxXPzn3ATG
sAr/Ed92J/t4szZNGTxo5VfVDHqgFME3Bg6pbyouawrcicqIb4aYFPirBNQsE0vW
H16uYgFSTnJyGF4Xy/KlBiRXqZzzYXF0yF2YFOatAVZa+INvZ7ORkxKhkp5wpXzv
jKKu2HAICJpQ6ADDwdzQKj01IxRDLQ926g84kggjYvfhav5rA9CIhwRXQwdaPsfj
EvekeH0tCUYxxFk0DY1toroGbSWJ8Jby33eE/CHsf0mLs25fVFkN4lmR4OUEzvFA
90xxeBHuyeGD0MLxVkGs/qLa0T8sJn170mQmTWkOsh++sm82thmeMWH0IWBgfS1X
XRwr3U4Bg8ECa9zIcflnIm35zxswuo3aPpJNVEwqbG/keM5ucZxrhWflum2zs3nh
0zCen7nFqoxagS+i1BvkEJ9PipeV9axDVhGrKwO3JR/zyoZzd3rjiCMF5yU0b0Vp
msruItfQ5/eoE2QGmvweYfuKLmKYOSLgB3OD4aVjYc5iOVxnEeqwpRXWZ7te8WuO
qfipTdfkaA5GSAH6so97oFAYFbOIzZtTW4c+8w31IeqI0zLng4m9lgUsieVYnah8
fQl+Pun22nad8Z4biXZ3C8EKPrL9SNAtBuYhvyUHh/vqpKmKRoOuVJt1UTXcdXJ5
Rc+7m3vij5ws7iPi0W21uqQDiMI7YUR/bnl2WWx2FguqZ+Tmqgl0omWeWRt67VSd
n+STDqWfX6HtACxa9eeWF5cZU0LIjf2EHGeMVgKsqTKsW2kyfoQ3GLVFmZK58Cve
XLlzxq30+RWnQ4AYQtP/HF+X8nBXhcel02on12E5M4mMLzkGYsI9KWCn063cD1QY
0jVBef25WLDSO6RWJOvp/HIEHz5uZOQSo7O+9sMvzr1MkgLrpKyGqrR0JYJUTMfx
2L+8KK0t7OsuHVlcNA2opoPeCkHlOn9whdmYT+aLQVwRerxpGeT9LKGYGXfABra3
KmR0XgftVXyB44FIY382MMFfjRyAOr5GspM3+FImVxyZwc3eq+GHXopSK9Sdk8vc
KdtAPlvnUWuMxKBSDGJ5eTJWf0RoYrQw8SAgrSPyHl7d9e+nSRo0DX6dcQNcSxJX
XIXAsaLbKObVUk+nyRB/rrwCXACCEcv3k9RU5z6hZpcdawqrzd8YRLHff+UorYHV
DFBshUhSykcgGg6diJ6nBuIDV556eu/0AjnpsYGKOKbcNWumNHpLYDLg/dhhQ2DM
fwlDbeaU5+h+nr6TQM14uaI/Y+Dtu4zvVXhlNqVN++MA7WWMKv4QtSFfFB5vd+VE
4DJTQr5ssSGCIrd1yVLdHz/dtVaosCOc7CugyMUf0DkNFLtb1bSnxjqPlGRyK3kB
rJSy2fB3YrYN5dWJCf7Q52029OQMiNbWvSyGAw/9PuYAonFXlIDedZQm6YkgR4Wl
Mc1qCJeX7aFE2JCcaY4XBoUmFfHt3oLAMeymjOCf8iXNyewjPhgPpUpHW41oCQ6w
8Pmhb7vSosBEDJyaJQ65pk4z4jMUIqkrZ+klGDOuORaOKk8YwRNR3E9iAhYAW7iX
/endjZByfQAhmH3k0IgeFJAiyHgowN93QOb5SnkTCOCnLsyQJRrKMUfvU/l1bIw3
dXiHzoTX8hGxJaQ0U2s3gZkw+Mz2pZ4QioeJPjIk9MrTUNov6OjEQ4OixB8etNyg
taFx+1lCnSZ9TUFS4M44JXaX0Gvls05GuUGlXq3FpJMT3fDIBUNIkm8Nc/Tkdcsq
YBGan8sqSwZwqO0ZM3ZR0AlaHpvFBMlOub0OpRAxozX3arskJzGGPHmO4UHZYme9
2buk85ei1hgV2lk60r0LGV3JPYgcGRY4MlipxY3vzzVJCq2RijTSaszlHUqSR8EG
e8f4xQAQxmLp/7ZYdWY8azDh9Z5uqzTxvrfgl26BpdNX3CmX16C6eE3DB2kj2RTN
Aa5ICtsU84sl6P/T8CARVweC9rETGY8DXD5gjD+tMzv/Dx2Fv4S1ghjL3TJwYI0s
snrg7yEwAg842mECBTdnBn6+KObxuxoiSEspw1Res2cxyCe0gKNMhpCSwa7KTHiG
eUqvUWKlummneCiNmWL16pAHlMtb5nKja+WtqaCzYnfU32ZDc9QfAn88mGTx+UPb
A2ng4z3TGac1A0H1r3aDvo3Exo3vkdU/n/rTg/7rySYAh5BORGA9pekUiNFVfBlq
yMOFee4wR2fIPo8HXBTT1who6dCKNiwgTLjET5SS+IzQciESJxWBxKvia2V0NkxD
iELFIaIazeJkopfHfwoSy2BbVF3pFOuN3SK0vOY1twD0mLzt3ZuL0B1dSzrkuUO/
FF/1Z36eHyfBtghWgLuB8oARyOHYl2QGEcZIQQNwWnA/vkwuHLLNXrcAkABNNfa1
PobRR1l3qx3hChL/EOJB/E6A0/tH1Q/CVSPBzAskx2M7SWGGWQgRHnmhmzXdVocw
fPSNpR8CSn7JUVgIocEwtnzUdG0mQGzgRx1h3oa5WaoqE172L8Sd9HBl6QE2DRDc
WlMQcz9s63W5z8t5kpReHLAV5inZY6/ItJEPQKlqcHEK4+wNzy12AhfQK87NpOGf
5N/YJAsLLY5WTwcq9rSSQAlPwYAcN7NLAfWSLv3JNT1tOIkf/UyiNN71idJgT01C
eC5YtN+nfXGiTqdGyHkox/QIOCNymoXt7N+2S21h6aRifyWarJlVkRuD4BHhrf/+
ZBycoCtOlgRCEQBlgcrUHHpsSfGiSHdfv4ASdh/zObEwx0MYXAazlznurGqR+ZLj
/vJIu8jRK+ye4TnKzOkBISsQ0eiXQnv7Bij9pM4PSPllcBCZc76CS5owjTTHY0Bp
fOzi5CsgagPwr5NKW8kTZ0NawcH7/zbAIRmcZ9uhIgxplzGrji53fCMRm3G7sAyK
JnSbdFyEfyDfoDpj9m8FVrWJojUgiSwpTNGjhLVkEumOvSRkHwCF7lB4kATzdWIO
VtSYHYyytD1MyPxK0I6LcrwwR2nxyywT0Z7nXJXyEkdzA0DaXeQ2DEhI4KbusA41
eMOEeewHn2upWQ6ywLlhfSzrCAwmGPj8ClSSzOZtr9wAamf9VXj6OdEZPiqUb25M
LSvVmwiaoOB+5rkk4+eCxru8yBKAHiF8k3rsN4fwXjOX8PVOg198aqeNrWn3U4D1
QPKrW5GpM5fCIEDsSjjB6vHhRtOp20ZJvBb7UXrJ8bGNJIWhVbEl5h4e5OY8Nhph
/AZYL9TgHvFoup1OieNo2KLXbBK3tjOQl5RPgXQNN7LoTcyemcx0jIBbgMyA5rZU
XhbTDghb7Noul5Y0S4lxCTAx4DOqdos5PW/l15lGohZduh9EvyynV08Ge8WGuKqC
I0S2Xqi6aBiJ95i3zalQHLA603a+Rak9YSLynljtDfLuIIm3+9YOybEb82SBpW1g
2tih56Zg3bMsAQ5rlXcxALy/eQ+RmpQL/HlQlNwCAoNxnv86dgCP9q0gSjSRBiFm
Tk8u9DLupj6rWVZiGistDHftORaK8VTDxgaBnTJzghfuZZweEasxzKB9V63GH1TM
0Jb//NYU48B7fZBZ3bk32GlONXmpdVGP3hPu2Aq31F5RzyREBI23lBSeL8rCr6H7
lNtjSp63qqDSS9bNNLj7o4/iYkoi+jUiaYssCbgH6lHZC9ZhEPEFkDKvW05dKcD0
qQjKCTbzOE2xvyrbawDgifesYl/NCTiC4mqui8czMl/HZpeh6ICJbrIewrNe4AGv
gG12U657tozeI0mCOwvMVYzwWJ41oYki9tVkqNNfL10bmmwQ7DG+eWH1UOdk3Nnz
ofP2nDKU0mYyKIG3egqIYQ7NGqtxDC50VOsz9ExqNfLsJc/jlqvLvBfX/1PSF59k
Ja8+E9QikSvBj+v5PmuXy+0Vo5Aq/mM6LA518Ql9T8eTJyvcWKkb0iDV3CSlDLRM
2/IWXIy/y5RZOTbkMVxAb+XlhsBU00T97exwvmQszbBA+R+VUqd+0j++o+62duln
CMlj2SrGCtnlPkNEPg2g+NKAIN6HaA2Lfl4BnSaOWJZdcVy2xpiuEpFJwlbuckP/
0HOz2oXKNwEAOEAkPgIVYNFjXB8MTA0ZbRLfBM61HXw9MDCf45WwGUUvTuABVrux
ORuwp/MfYCGgORURqO60mtcst+JbImz/DPMzAEUyFr+NlJowQuB+JoKLkDIb5E7R
TrgzdR5jfPF57XaSpMmYWO97o6RMB1YKct5081+Kc2IMvgBDThIlzjN82wNSJSPt
iWSlzAlE60wPdpWhJzynEQ3wrFJXQBqqeFQQaf87sEvJA/xexOptrR6qjHwK9WFx
YtZCAzlEYX0DN7XFuREIm6Ui28kz9zdtYsp8M0Z4lV8HADA63RsQermy0B86HAEJ
hOmpWDfdUgM4aL8rkVQI5usE+26mLq6GOxn5yMp8iMoZ+q5+VMS8JUAKy7ysfXQg
s27yq6fgIaCsEgBIPl7QCYlRBWWk1EuA3tMrnYMdJB3Fdal87ZG9xvje9Q4kbjth
apHNsd54Q6KvC+aCi8NiIRfw/HNzgzmVWvIXiHw4kkmuZ1DDhZ44/kffGjaZfLA8
S49AqVEofIYY5GaYCjhfDwQ16kVVMVtx0xSgbxBAjvbmxRToNPDplFhaFKkWZ6xM
49FITSFa0LFNtxaz4VtzSl5Vz233foyxhSyhJq34zBrewuS9DXUZE0VPJ5v4mat4
Ga9nNOSPsgQYu4lwjqVqt24/FPwWQ9We1XRsY61lbAlESgxSQs4YgdCxN/ivwgzM
sQ25rk3Hs+2/SndkXxzTXtR/D4j+CDZsejPQgdG0c6zzY9dlzVdNrfQ6kgJbR9kv
skI8IHLKBr3a/nBbi9NLmE4682bhiXOEDMSSd2IVIVlFOIY6uCwaaM4+9u9r4Vyz
VPuazrzowOXi+iKgp1h5lTXAojw3piXal/wZNeS8rNpxuFmusUHommjtwzQ0gg/H
vXSIp7VfcGZmPnDbZx8Wgr/VAtIBxIUNizBLI/jAko+KTfFruXV/eLZiTV3KecMc
BK6ct7+8whvVGypKpWzqzNZ+eh7wjCwfWfEq8EeCoRfkQYQ45Xg/LMaabTtfYQqM
MVPMAQhXl+f4KrT3giC+D9K1HUnovnZrSlnqXDKhMUGUmg9/stvD35JukMJ7b2BB
SQiE06wst4IaUakkMzaxc4MMREw3KYVvaBsk2KesCauxgURVDxRS5Zv+GWV852c5
rD6n28a7fuPSxsGbRDKU0QvaGjT3xP8D9lrBpWXFT2vJMB53LHdsvEtowsSRHq5U
lRjfNOk9MRTHxWa73okVvQjFubYa4UKCCJN6SDu0VxNR3UxXmpCn12ZSWcwoaef0
yaDcU5id8AeGIcQVUd7d5MvaFC6lJKW25qlbZJtgyEwL1J3eX3Iee4+sg5troU80
rqKxnngmH99S5KH6Iq33j9X/yt7fR9am9JP4JaVcEZ3YIt1f3RqudXSkB+Fcu2zv
MSpci4sLIPLdyraWc+y0JwzJqr0WFvob1zrVyxTsla7Nj9nssZDOW8m67dO+TsC4
gJceNtdUSt0R5hqUBZRIm6bpPuCFeRD+a8a1c1jGZMXr8mT807sYqGtXJsUvK9tI
X6C3KdvqUzczLuMz+lCJHyfu+rOguJ/YTT4mUaGgtzXtxbS8Rbz/cuz9qxfjoq0v
+/DpvJ8GAj6RVn6RE1VWwD1urubEITj9/7xpQHhXpJG/8ezZOVkjQEle9oD2qd80
77Vt63WnwfGjbUlaAc8Sgl/ZzYBdbSRPp7CkPPGm/C9jerWYiSCX2vlqVW5Rkl0f
Sh1c7Q2UxFBwVStTJecVWxFnBxVUO1YAwE2IVLzrCKKOfCtxvhuBuIi3Vcok3bBO
b89Hdbakpxi2qAdq9PuKjLWueVZ4FbvFmkovFOR6atupFWJQjDbR5dvWFqvOqRpd
SkvUF0XuwOPgdD6nLEtVJVqN/m660TklX9sHOvU9zYytXsQjdvnPTwOlmNfVhOaR
f1mx6e+ssNNGWyY0zlaARpp9YvZ/AMgaZd2inCAXtl6N365xqJVW1KZQl699WbvP
pdjwMD27EVhOVx4TY78WIhBeUA0azzkKGkR1a/h7CbvfqFQhE5WlXQU+FyRwLBTA
Ar9aeiXsy9s5+Y7O0SclRol4KQWvbmDbIsTIguBmD+ji/l/OsZMNmxV/arPCVrPD
`pragma protect end_protected
