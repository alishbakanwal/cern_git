// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:45 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
kx56C4egvFeiMHhMWNrgwJG9gmi6P8l4GsBDRSPt6SyaKG0YbN7sZIa6nB31YC0l
En+uPQ542UsQTrZnMsXPNe/ByXtXMZKK16KwVCaE41jiciybpHmTpvIhoSIxTBKG
gNMZG/JKHQ0OreMYIG+8G1FgdT/UcuX/bPeX9R+m+W0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 18320)
JKFc41hpHriFcsTTa9cUW/UIhQkP0i4VXqL2V/o9b5vwMVTCZjNh8kl9N1/tbGfU
IUXas/Ag8GO9BS8qfIwDaKE2oQyOlHfA7WRvXoo4J9d9gsZOus23bkENKpcNjXPX
ysB2vrHPGZ8KzvrZ58964uTeDAAqPnDDkIickY5iLzJOroWGQtNQknLMSvL4o5HL
BHIWJvlUcWcMfs+vc+C8rzEfy5kjZb0Ca9srA2VRYU/AyjFpQmbb7o3KuaM6FFDd
84BKPkgSJDchlPzck/XCkgiP87om2pyG9qmBw5a5aAk4IprscPIXboefij0utTKM
ZUuskxxSs0svZEWNUWOcvjCM/JlYE8YJD4FYiRyUog7cJHkmUtXtz+gupx32fcVL
qwiqJYXJhjSvTdjiQ56i6DdhYX3Rsiu2gKq/k85ZnAATJOwfej/MFEorc/bp6Qfg
ETS/rUqd0xvW5v+CnHHz6EsCmVov39EmVDhxvwojg58AH5KXsaZ8amSKWoHh9NEn
Hm0S9kO/1lSRdTHsneAEQLLzqkVYmOuntj//+k3P07uPAPNlT0xBSsjqI48TF4qB
FroDyjTBoTrtYvahUXBh8lj0DDDAFJ+KcHcNLlij73d6Vynz42XciFWd4NcsCSN4
JxmIvxFh6MdnYXrq+e1YbXWhw043MEjN+8fQRuZodMzYUXPT89K9Wusqt7U4waKz
1clfU20xSIDjn5MxWmauHDxnpVwtpyqAQ0mirh5cwI60vSzY346ygQ5Nl4ZMjC9V
GTi1xb71US+bnPaYajwsqq4RbAJ2WfKuHShj2AY3VfIFaOA0eP4QKSebVJ1Sx7RI
z/ulX0bnAwVyc5fX/52S1cAQJ77tjtMWGQLxL4P4eFL4E0PbvIXvnb8jwD9MBMEr
6kQ62qLYHH7KwYskpjYL1nBnzsPI1pTrA4+ztr4NjFlVZ9u7IbrT6FmdApSRVBBY
gngR+TgqN59qpZRg+qIgOB8mfzzZdDIDeFPtYCkSDHPmEgW7Gduh5atcHK9B5voo
8VZigrEJI6vrou03gmsheP4g/RlQIIa1wJLc9dziuD4NQIMty/MILlIo7Bcmc7ON
kor8/Bt8M80Eo7lFAzaUKLAXJyIx/RFM1y9AM4Ltl3lKPp+VPfYaruYOSYwz31Kc
WCmBieOjjeQikjcrykmAYVrYIYH4e/QFQBTMGI9TTGxxrfBRxO9dnxPOXpQ4Wvd4
3mSPV8gzJa/O5MQucvlHMkJNYClj1APQ72MJ7OsxbuaOLOi04PmKTmsHwzALG361
k2JzNMCBuKwszdrzVAyE9q1nh5bqClDtfGE1CB9HZbN8B9yDWNHyFXMBG2NnxL3P
6sge0kT4Jabnut0lYiKeybL9RvIcQXdRoyFgYvdS+LkCyKxidVDdszrXvrSH8mUJ
Q4h41bxIDE84oMd8PinlqjNcRUxiXKQ90vOrpeJKRT6o1NuXbD6R1ahtV2qRJ+aK
DvWedGPtDhfC6SS9Eln/B+XlPFYQbp4AcounoyUl7VZ8/b6IwD1EROtQCAKD8LW2
RqVV4x54N0hVt67aPh5BMj4jVSLa1vfD++7HBw11AOL8VTOYHQPJOuIC8JNAYsdb
KrZazVDNgKv60kl5UhwhsGpAOMJrA/9KGUKkCZ8T53vsBTnlKg/68JTnUBZy3Qkl
4eOrfORVBZvx20b7vGfgQz8FwHS9vh1SAUt9SxOm1nfC9q0oCZP1w2LsIxjqtt6v
Ekz3p5yv823EFt63HO0s8o4iKaKhqR9/WuIya6V+f7qrZ6bEYfSZpk7IGuUJmjN+
OqoA/qYzRU5Xak7rSdGAWWrFqSPt5z8MflnCsj+9Uswhz9m3FdLK2116jbfkEvmE
m1tclIJsHjl7bDmC/gP7wnRsHnqFENYpEbleDS4QBzrNZjG8hcmLYOMGwIaJVvLh
FP2P1Qg66FnKOP7tlI+wuui5bEd1DYXCuJcitBT+kLzE+RBRLFKNdXO6sHBYorlD
zqwAhxBJTfvwpbn++9CvIa6QHniC4SHqhaKlSI1oMWyR/xUne17ssTJAxS30Itiw
y3+8ma6984MDSbd3AKnfE3+Wbn+EysjPN2s9PL9HQkD7DlfOJM10lzfVL2T46TLl
IVvdTH8U/VRc0Uz+cR6+ulDqAFY4sBYoH4bfn46sDXqKnosUzD0+zssVdnuW/wWc
INy9gFp3GLX4Rz+/ztwp3xAxatGvZsZYsaFCeZ6jBkTWmS9oJt4+nmfsdkf+fR6m
rd+knEuQr1pW5IaGb/M7pU9XJgnCgbwEbpkiToausYr1/ehdFwQvXcabBOSUoSm0
WrRwnJyMJC5hbF2S0m2X49LZGe6DU8c3b3jia5Q+idzWkzk+5fDpdfldDLqzuBLJ
GWRZVbPC0mJ5oyRnVtZEa7TS5KVxEcfqAfpn8TxrWVFY4l1+BFIpARdJn/NV3ak6
u4lfDZZdA/fAo39q34FBQMaHFcPpV4FQePV51SQv2hgaC/9L2PZdqU9az/ZX6/dS
ODBZH7TF3IXRPtcjtcJiwYdjgEybvIjiaTASL5/ZFKGhAKlK8IV6Ag8V6wSHwmyq
FCYEmittR1tykqQ3QOHzohiHjj6d/YMzj0AIUZ3qZMyDgI6kZnC4mgyMFWwlWrAa
kKWg4MxZ7aKIfAjRr/pYv014914DS3BMYSbSIDfQEIGjjHb87+7+GPpZ2+JiDcPg
KQKAB/kqkRBkuFbRSf43r52FB1E1rOAR6Vs3DAz2oOjGp+74NUoPhkTtVlI/qCGE
zl+pyWusG3X4Grh468eyOkyfY9fyURgYYOLX9y5+n36Z4C6GUM1U9PDYrXH9Z7cQ
evelR4DWKhWrHg6CoSNLMVzSENC9EA23BS/3AeY4U7Uq9v/h7paz76ItwysPPgpl
cjfiC8HKSMy+YSlk2xuiWXcORb1+x9MUKFAy1ek4f+zA79/24lH2z8bBhMKjeb49
IS94PwR2bL6N7RB9ZD6WS06Op3k12anwAzjzPeWheUP7E6+utq6UHj+kMNkxi745
X+gwFpcUeTqvFrgukrHhAd30/pTl0fTGIZ2vhpRXQEKRqAVwCJcFck3cNYCnGYgz
/w8zuYP1WIystj5dlMdtXRl+8fjc5WgvrtjgojuRDfAq+nrQP/LqwPadRTYIrtII
kgS1XPQqFZOQi4sDzgmxzyfYiELXwiKliwjx4/NiC8kPsHWX6hhbD30oGoETZ/pD
kJupX8r+xfl2oWLL//duW2pV/IPm7G4Hb0nqjNqVbiCWj3KI5CDbCOLlDViA3ZRj
pfKcVLlF93+MdOC7EzjGdAaVM4kTHMaTBXw+qNbo1ncMgqGsn+Rpn3cUeB1NOKQa
FeNl5NmTdscS+L9eI24r4Qy48knMl6eC9eEeqOvIIIiL75In/N9vEWZPtr65/G48
USeFsbOnNVCxKDUzmhM4IP3oDnk1qTQPJvC/rbIikdrvnkUTomK9GAMJy58RQ78z
EeK3UV2unEDPwLfu1mMPWPwEqFbd/g0lzxtXUYQ11X60s9h7ESmH6/setcEKAYjr
iRxmookqCfpCJb0m33/0ufGoQAHHMjSqqSWUoVozSIUguGD1w5Sdy3F+d2KrlPX1
vb3NMDXEdekmsnAXzLMSPW9qBIbgDDaLZbH1SAeu02veGnFA0LpUyqtwTLHgbiHK
AC4mAV+9PwvB077oGCkClDOlk5jsbUhwOiTYbAIlNXaiBp8G5WGQ1rT18M08sf3e
GrnsAt50pavbcIgCmdX9XRQeyPJZdt5LIX39LMUKwr2RyW939UBQbRk8EJxcjIq/
Po2gj5xbRMQeU3eY+9zIdmQg5jq2HagTgt6/JWPGX9dtqHOYqAlgSrhRiy5a0OOl
mG556I30161iOF+0aN+5Nq6qn0CTAmNuvLpoxEBBLp+Q3a9mMGJRPee7xe29dQ2V
IupayBtqLSzxssFXjlMwjhqJ1l/KCBjkFmonmETciAigxUYG1QvRmFGpGntJr3FG
xY9XQx78fy2LFrqDOS122xxvnemBD5Krb6SPihz+Ln2uSApbqvsi0EduPQOPwtAD
H9mLJbEPUJ48s87byYHydxd6xsxtiI/WUGwLkYHoahaymCJAd8YgjzsLjI4bHbLs
Hhk3Ze10BYau6YRsvGr9u7Qe45FMyq01+0OEQx2IVIfDIC8/Ev7OMuvbaOzmGvHh
Uqmlpr+3fI9njYFh2fe7NNnipDZp63+rl4CqYkSxrNPWNBtGkhfYK5D79xP2mvEL
o6QUo2TztqleASq2OOBzF4po4+0Dr8O45RYIOJz+A5q6VKAi9uH6zdQoGxKpOl3I
c9C1QcQIXgqCuUdQQmpHWaA7WGOtaapoNd8UAWLv5PFTkdBGQb9C8ybH/g7Qz62i
3iS1YEAPqggAoP164ixZ77/gekY7v0oR9CKvQapUF8KFO9FTyb4SACvpf16zX3uN
u5FZC4KoRyoEdmal811XQ7nXEZH4FAnrjOFMBlUd0U+wd3ZsFcjd//VZUfoI7MF1
mgZfArX+Yaf0g1Fo0wYBR4uPWiFG9ljmUuP/sflbwx3GSToPnjCDxFhmX8bbnxLM
kTr6A1kzGqtkQPZWJeoKpAQ4JWK5Rpr+J6O2U5hru0gjqjDgGZ5QVFE/JY4V1jHw
oK/8VH6+rr6VfjM5s6akDZcSN2fh9J6qZ0Yz372vaPCCoMB1TEY2KtCMpIy9bMCO
8mfklflOvYeDEvPxXtfTkGACKrH3id5Ve763/6nlnoLzUqEUV7u9OnzTen50dIys
c+gKfZLo8Yo6ugbLIAWvTmqzuPMpMFG6evAlDimC5/p47Z/q4l6q2QOlxu0OsE6s
GMtNbNTVS5V9Ocf6lpXDEGApfW4sY3c03VaSnjqDW1jdOXT28YvZJ82CjbCnPPIf
INvwj5+ioS2RKrxpinV2drfIwToFk77lmmQxTgLK8nDCG6/VCs5YOvZSj9AFkzaa
b/6aAVLXrRsCy3lE96vT9Z0VEURAgyYBkQCIPaV2/md2R6JSwQtJ907Z7ZqX5jyo
KlTgeFQZHdd+eJEniH6kfDgR1Vf0HekgxvMPICX3lO9VS826yx95uLzSqj1jMxYL
KtGxGhT6SY2mlaZhVpGM/FmI6oMPC9eqzd4jtXwkKFLBODAWpC78F1FJ/zQrT/Kl
S+OvCTdq5R9LZjWQQyqTf5Y4GMF3X3uPyNAs8u78AsNxf1mYNm+0ypZG6ftF2G5L
SG4Q0tm1NcGXIf40dkqiQdyToDC7FwoBXC4JZaeCGlFD8sPh0ajvdkV8TtJdhrO2
Xrmz7e7f4GkghRnmxjlqlDZ43oIto0zcus5ZqZgd4pA5Y4UPvP91kDOt/WyXvlcC
w8Rs61Z+sWFwi/ju92ZwQaRhpovsnb2zaVzh1eqIcVETvPQnTiNa5vLKYaTEh10Z
TxbWUs12i+V1x3c7yOMF+w73/8dLkPdxRa9GJ3vwxaWc7mseyypyIUZ3gb2VrKU4
ikz1RFG4jiMQFBB1jTEM7IZf6p/r1A1jNaP8Iq6XrEhzslEwIC45l2sFutGNPWZr
itxzbJURi1jo5v0LQzDp7bayiGgfsksLGKAEigBlgj8AjqqtiFnODhEqTBBhnjAe
s/+robCMO0yeu1zhA3u0WM9aHsc32WAA2287dXzqatJu4DkqbSqk0pWI5pY3Ic+A
8eSfWxYQQTYu7FNqevVzqztqT6v/XiQIJDuV6Y21h4MIGSN7EwJeIXvkJLunlfAS
rN9Q01nurwFFdTe7lSd8AGAXWUtxbjuC/vWkOI5PTSh91mfpSdgwECCETgBUY4h9
OIIDq1d6OvMhR7WOmKHao0nH00EYAnVvN3eMwHRFsi/XEYdlID99Bur0HwQ4fxDb
9rIL1I0M7djfhdsi4PXqI4hVB0QO5HoHRw3ZX0Jvq0IfpMtdfjPMQNeEjAJ5Mkx7
MpXSfGja12QctgSbmM78YKuOVtirMaQT7sHMGyT+Xwh9IRRZyc5NJUW9Eo16a30p
QV+lnHAF7UatEDWmsokuVUdXJKoSxhcM0WqPK6rIFr9yztEXp8niHvccAhJFQw57
G5YCFr1RN2jdIyhZbI1ldKwFkFoehjpjh1CiWBip3aKUuVZMU9As7zRktcwIiTS3
sjDK8v/k38R92BBR6rV+Bu20AonqNZW5D9EGgbS8JTbkcrIlf/y0iMKoYqxCDNTh
ukuw/c5/1k+zFSvWlHXJvW3MeVEjkwClWrNZqcJ4sD6T+olKMLSwH9jgIEWxQfMS
RkCI6LJKprb/3YrBaT/ovOlqOKf+GcrLjcYAg03zmTJpqIaM7mE5KDepaiZqhvLB
wKiKMrP9D5NDWpe4WO5WmUOb/MVyOqKb/rifQNl8YlW3f6QAdNhlMekWtq65IPT8
/M473D5IlXiRFr6pYERiDqk4NviA6P7iY5DU3hHePwnkau8EJIPeAqEXtK/bgXnq
oDsxfPeLem0xjXF0xmoJ978EqhTEoqsfcLeGA66AbA1yLNpCXn+yqwgn1Lva6nfT
HAbyRwzHrZt2rC3LmkPUPicN5mk7GPorAM3b/cUD1Cmm5d2ctjqjXn4VaLjUFuQL
TFMqqcbXnas4+25kSypaWYrbK9xnzhfQaUjHWmbANPu4xGWBvQ5DPm4wcm5K6TzJ
SYIkHilcbyWKdtz9zGmliAFzxHUR0cTVJkCKJewaqZDQnnPsCknfqti6DcvYueXC
2CaPar86pQCkaE2w4VMf4H6UUiC5cLWq2g3ZY7G7yan9IjiIImczgNYGtgGiLCqr
RNnmrBpvKTW58W5SsyuD1H6m9K6BjTthie93wPrHraQnc5D25hY03ejlEk4t1gZa
bVMQvGm6VFu3NMrpfXx9QKXFYOX4cJ8RlVUL6yjc+J0K5X1VI2LvOpWjCwH9wumY
AMIDtZV0CZhBEvbh7CWM9BQHxsp0GdZXYaG4aQR/jTt2t3PCgmXgPlsOpy4UsQJX
gND5EUW+5BMs6zaVwM7zccJe99KdTF5e+QNdvqetlN43qbOFUTh5B6nGubGxtrYz
b/iZYlq3lDhXzcoNYn7J+7f+HRkqbP9NpIGwb8NPpJlFoy0MdtObxloKK+rn3rEV
mDwNjsWFt8BnyA6jUdD3I2hDwhBlD8fXcU2YHlUReuCRhpF+Zg2hLUz0Ba/R8IOP
msUuNV0gXFxJa2cwTbl46bXG1DRvT7HOFyyk21xv4L4EdLtFZ08aIxP/eSCLBlOu
tYmpjuisgSVCf1S+/Hi1Qg74ons9+0v5/CJg8HV1wTolKKbhF5uJwmpprme44URY
dGEBIIEA672Jg1rxhiIvO5OzfRpfvPAFtsU9GE4uUsDwzuapqxcv9tWbYrore051
gq4d7eAw6yxQQ0xd/RClE0Emv0Z5Q8yjmKRZwZ2nac2KuzlA5/OW6VWV4szO2+ha
VJfAGuilgdz7rSVaNsF7tIHL/Iyv+LMVz3SA/B43xzAZEBGTnJQUWt28YF90oxds
83i4g2qRC5AQg/aSogKOGWDCUwuum+UX9YcL2woaU3MAaF887xhhJvftN4MuPIEZ
CpRLX6Q34N1yffGDFpMzMMTlFtl2R70sJrZomzrNjVo93A+XhHEScLOzJOvigTDo
rPWy7NEZwVFrq4oMFtEr75bGC82MS+4/q4iwO5eaMZRuTV1Hgak1LTFEohvnq27t
jX0n9T5e8hiPPeUThvtuyHK1GAaxCZPxR7hZvPrL1kln99KlXj3UXpwoljbeEY30
FNgOuVW/DntZKbFgnrs4TAm0mYPZeD6NVjEmueW0F9yinnIYx9ex4fLiodNGyllo
frHSakLustqbQFpPTqrcJxS4NOQFUlSJmeFxD8990DSkFJilzODu57eV7s5BgKtK
UG6qP5QYAitv0+eSXS+QJdByF6MmhxLg/WE6/4mRqfYTMAPqIlvnt8eH560QKsWb
iPSkUvTPgL8Sdcp3pgYe52Gs60VSQaVedIaf+XURFdnJFxcTKOYUsgOEjvkLRW6N
vkVsZY55mripeqYNp24jW6rB2XmS06oWuXgJJRFqdWTTCETrtmA77yxt1RWmgePn
9TDW0lUoaTtc6msjcyciGT5KwCuWOmM/CeLGLOr3I9lzrLXCRW48AV62kCyRj+SZ
4PrrKRnB9bjliFBDS+ofHetfhgIOYwSSq/4Ud6wu+9mKhWsL1co7B3O/Cihf26kN
fZzrSYh2vZx9SFypLIFKZZB4P1mnkdXqfMkJFeNi7ezH2E0sFQwj8kV+cXvifJ8I
khqwH/wZ2OKmiCPc2McVJxpnnQ8F+lGKZ4AGs0EK6C6rdiXo1JHfDScxs/+FezwZ
t/r6J8xRZ+bgwe2txsC70MlN3VzfJLI8WeJOTPO2WhxS+q3slkkdtZb4znnx+Lia
0e/d+YlD29TCoQtsyxgYb2junHZ/ThBQJAXVr6d8z59iYfrhZg6qeX7OIxFF4fbN
CdeThm5Z1yG7mU+3fUQP+by0Kly/q5aCWYaKZt1KpD/sR2UPWf0vFE2GB9ZdJe8t
eff33B7X35sFoNCftr8t/xoOYOyg9WpwNSFj/pSbrqo6MC6yTzVvQWg2TRwKFmH6
4RGzVWSx8Fa6Z04cJGOsY52FklAoSYOOOoCXQMrt0etFzvFbTP5372RBFlfp0iC2
ifsmRC7XoLgYuhJZh4evtz7//8pe/Fxyi4q+lEBdjPa9OAnQHrkLL5n07Um2f5Yb
cxVkvQx7KGBrutRPR2dKDOX2XYzEgkVt/uhoFD90MSvT8ZooxVUA6+HGinwxrh2w
70djR42uVoXd2xKCdc6+ISHAHiv3zo//gsjgP0buMh7ZrgL58ctn/R6jE9IvYrn2
38D1ELG06rpz21EAu4/UiFDO7QhUTCLJfmIg4Bk6HHGcTWg8jobjy37l6KEVHQ+k
v0YO/CLcTEMMHzeckUqVfPMDRKFAcLtKhowWveUuoxaMomd/tPzqkUA/vHS2chm2
d+HE8pIIZBlYYFsWU42E27RHgghOP3NljRDk5KOI0CTr9qW9OlXTf//UCUV91Xer
UFDzQDTV1Ap9TYHNHEp3ItGxDpy31z35cSM0g7WAY2MisZx1/IRB7ZsscD0qnxHP
hrdPHpWYwvVHO51SguDbylt7ShHrBRWqgOPiVphThq4VZnljl0gt0djUr1DKDHNL
rKexyThGdToQ2kmdWWC/v3233ZAxqPp+YphZtHYL3e6xict+f2KYQlRqIiqs4t2c
jHq5QBAJfKfwa5eS70+sjL1usQIqP4bnCBXwVSHFMZTUZa9xAxgMCUk+1Y5UvS0R
Gtr6xsRlas96oDct9DqukZKSB8xAYlNm/Jf7NSnxZ8dBRSZGAQjW3hAOdjAMY8jO
voHJsgK/lUjeuvwifL08F0nVL8d/u9asLdEj+3OO1UoFu+37B1CtpOWk1ALVKPq4
naRcSGe6NGYZimoUUXRSQZYPM4aNjaT1oXmm6dv6lNhUBbZe0cgkMoj7MYYRdvfb
B4xcV33iE7sa1fI1nB0EXjkKvTTR/EOAF/b54w7u331+T/uxVmJIOb2ooumbQUMl
zzGqeXvtmEtq/Fi9VCoIH4NKFs58l7lwekp9evQ+kOCg7tGSA8mY3YqfltQV+Dpc
6wt1ydOWxlBufBwQFVfbxzTWY6FoqTYk6t3uwcBKP5LLSUL4dUPvAZV9g7j80YNZ
ITiBmrTgaEAZvvE6mDFiv8I8RgZ+/bdkdx5xADaRK2DzEkb3ZcKeFxjRWBY3kCG2
h0N5LYiy1GWBGXCHgxtEmAjCvBbJ29yqYfEBWH+xmjiHTzEmODDRfBH5Ok251sTs
1SYG6BlCNxfbKPJqvpTWWhPlEZxuZIXVF97sIwXJU7/MwiLkTVKEJlv1Uo5hVPaS
M7he9hEf8BUqkfYwPmLHunV5zz4Swgyf4kxL3ON7Vii5Rt7P+++pWNkbRBq97KOc
lit9FOKFofKNIMUIld1YYHyq1+euISulPVqM4A0WZD3Hxtv04jBzL1uJ2ySlq6ss
5ytrKWe8DEWbR71B3DoJo82VUlDGY80HHMfXZSZZOSWOCUGLv8Xi1B48AFGCuwNr
olp8NfQX/Bxoi+I7zEfSqJJeGuSCiPqgUTlqruYsMigHVpKntK4n9FTuxt46smJP
yP2CJA+RzQkxLTPDh7bftSsFVU4YMbYRAS4S1qCZaeLeqJpn8RQ5UB1OSEfnJ6Iz
kbhpucOgC3+YUb4PNgckHBjpwcaJC8OMsnPtYiypZFlow18rbJLjrsYRc4mwzpq6
w2iKue337n91gBEtYvaKME2xXn67i7aOETFjkqc4WM9jpoa35JzbqrBcu474Obnc
LcoImSkL7pkAsUOZALhHUYfSBgbanq9gkFgF51ixj83jEK9Nme83Txgdb9mCz8DX
4nKWJKLm7zMBNdFhMKBoPspZjlmpoIo//rViN/98HdP3S2eV4eVyKdf+CBgPPrtJ
6QpHZh5mVNFO4nZHw3HZZ13joarz9BcP0sQj6i2R1yEbsmpSLq05wtCdSFrdD0E8
XNQm+hCzS78ytEEnFZkU71bAHR/Tf9gDZY058hZkxyDR8jTR8P/KHEaWF7dhQECv
NO+UyubNcPVyJBr5S+Hl5tlcZmcJq+k8MUubQGcSpFsIF2A5Zj8eU5CtKBtg67wX
p9onLlI4Ixpj3QrNX8oOvhETt9dy+MfzdDhBawPAAzt9MjkgsBky8KfjrbXPIYJc
WviqSMDzedjg4X1e6ohfdSfqg+hXRpCygfPaPxBoRmLVcUpRPcvbmWOi9oIjOgtm
i3gCgvgnhLXquFY9BrensQMfNBtsX/gC3VDeXcQoqcvGwa9SzqGiheFDnoHRZCln
2+yw70RNcfBp3y8v+fCZYKp62LJC/4cQEppBzVee7VWJUdLVbd9noMdbSlht4E4B
UQ52OJ//Ta4TVVeaqeLPBu54aHM1j24QRtk3wFPlFZZ6HBMs38ZMY6T8iNbkMllW
1fnOukz90pdXiofZFPzABnEuIrjW/iH9JX2ZZQZ/QoYzm+mCFW1cvzwieOg2AGxD
yNXckpMEVSAMmPMjCI9uRQlSczVNqyCRRo88Of4WAJqF47koiT5jwNMPiV0C5o6M
QWmze3gx/UZ48d+YmzNIb5biRvuGk/ilr2mxxvk5/t9A8Gx88O31+bnu2ED3i/37
H3snKVt3riq6C9M6MFXjkRr/mdGE/smJ06sipxlvoaFCjxzg+yzAeYfip5liDylA
v+oKk/mpEU3eS7liRRM20iBZhbhc4lXzSTtS+6ek7qniqw2Ah5G4wPv+QdKznwln
+U/6kpbMR7cUFSF6CJB4JyijOSHEH7QCXyxfyEeH5/newFMXjvu9b32vm6KVVv7p
EaBjTc1+aUvZBoDUldEFoPQNTLEo+B9USGpGEgmGoe/93ZseQdyTl0Zo1D8OmH4c
xAWkl1vDtFzD1b0gzDusbFDdl8h01l5WGetctWdd/WYMtsjCEQeyLhh5TIQufEC+
L2yjRTKP4t9rbhrxE3TWNRMk262hrvSCV3KzY67kIRPz3bo2Mr8l2kaFa2PYCfGD
wTwAnHhEuP2C7roXL+zvfBnZ7IOFQ6EFmrW0TNAdOzok2laJKZa0dgmddYxJBttQ
J/3p8mSqzpu9YA2m2nlUh6D1zL1Ape+PtPNsQIX7ABVCRWv148Iqjd7FPYY2lKie
zMnc9NLpk5tD2CPukW3XrH6bJqdlsLLYF40VKLwgk9KvHeh3xNMZ+9XNsZXSS3wz
32SaBg9KjNpdCKC8jB8Q37/WL/v44yqvA3J4dla4j8gmsqoGCqSLq+hp7OJGY5J0
+S1X9erhPxy4QJLnWWlp7EkcWkaIfkcgul2bnfyKK0SeZwGjQ+nS4lzaFOYaC7iw
DvLmAWt4DgCRlPSXWChlFhMbvc4fR/8WzXX6Ik0tDcdF6+BAUI+jWAaQ7wsNnwNs
sSfzJbvOA3UyNgvAFrwdAhl2vTNVgvihJUREz62FqP2pk9JHZlVsdIioMFNbvjOi
3NOclpVY2cEG20RbAhbcvpNkOYR3oBWhEx3mPQe3i4V9LhtF71D2zjHSTSL54BLb
SuUinH1T8qY++5+22ZLVLioiXBnjgH2ksJ8rRFzKOrwQabo6v+yX6nI6vxOnviVO
9lmZMBzi0/OJLGcLBLFrIw98BG1zyf1IKz6E4AWBJ2LwGh3QFIBtz6Pfu3m4saN7
+bUvQbAQiuJS7JMqOjckddiJvFzg82vFAeN4R42DNUZkdC5sVM/NLv1rQG+RM7Xm
Cfz/5aRgpSPHIZFFphtCUWRhbZ2F/mUdnaVw9Z2c+o2GECHh3W5tjUJ1qb/42CWK
75smEQ8W+fLusC8gO+wObyVkcdP/e82eCE0zaq2KVUO78oYooexCgB0ylb8/aZla
fLi/BNbYRqr7SQMUC2CcCrzbAj2sux+PVL2uAksp1gI+G4diomp8ge6Rjtnb4YOc
X3GrcoYYuHKZm+gaLg7BFNVI7VsVKDg8qA/OJCvsjWMSn43+xHJWA9FUnJ8B8A5M
eH8ipQzpvk/3z0xLsOIE2UtaN4iF1bEwjeLAwQbXFN7LRfeJeLSIpdU9dxGjLZb+
Aw/XHDN5IawiVh2b6uZ2MR/JAnxZ9x4BkWhUPzW6DyBNtc1Lt1o/39O4dXSwxHK5
0M6H1KKF26yclkhPqaCzBdoCi2S+AH2df0Smiw5zFezyVUAp01RFuV3DIR7JSYF+
v8uJhFILLTH9DAq2C42Xn0BNqY+hmpl5mRlQ3UIk6d1NpUQCrdX2hyw5EAe3ToeX
VDSGSnxqKOHno/cq8DhvEC1cEmUnOUzU6KkW7pEYNBqZwTUyk8q0BOTsXKBJBQ2G
9swo+t14OSH0uHQGH2mgg2G0fVV6VptcjMvNon5icHZT4jE5AJo765HljMtmKyyC
z+536yXCikFuq47z8ZLK6QYpZzqt0PSkI+FVt24oyABVDHBFT6OAjvuhk1TetyW/
36a3SqxWFonPGAqCbyC6IgPa3hYgkn7rBzGuL8jvTfGV9dpidGnk8ZEUokmW/ALm
dyoG5SzApnTXfI6kLJSiO6oJSus/oPNf6HlS8byM/5ZociJyu+GRx7h2ZhzzG7y5
JH8+5jSQfQ0AjSb3oMV6eWpwu5EoMbkI8BuhxBt/W2d+UcpX0fhlISKGXx2U72Bd
vXQLwSuniuenkGAdqgNA0ehuh+I5OWIZC+W+XxnxjweYXReagQRbSEGi/aTs7Xer
/5/azrfhERjZ0ADZLyog5b8VZ/GiXIt1mepERHTvQNNKA+Y5SYyL0ZVv6yvJbTAQ
Wbv0746O2cBBew4LOCfTNDUi9IgsBkZMdIpnoTAgPHV/I2CplOaMR2s1I4WWWdtZ
WgbSQVypZcx3HtCAvNL3dMMU54CLgeYDdYBoTdS1lcHmca4aAxDIJFlQwNtIVWS7
4oOMxlpTXM1auf76nPUOPM277C6jAqdWj5ehQMAe7ML3I1CGltqdaAEIR4s8nymv
POHQ/DxS6u2Gskx1iiR3UbfnYMEDK006djwPlHEhshfiuNUz7Vm23CVghlk7C/lH
bc36ZItRMBRNN8hZWl5PEXL+Fn1j3MhJNBEAGkjMjmXf4ECYbZIE14kZegY55M/k
/pWcmPLUDHM4dTRButCiJcZyENJ6qOEx5/Jncu2OBMWILlrozEijDI6Ulse0aoci
E/ByN9IVnNXCuJjMaga08ZWo/YGyFV1Iz46bdjRrq58v9Y+cnizyrs3xubT/dnNb
ydIQfqn11SU9RSI7weqrpl5sohXKUS4m0a0X5+BRQYfXnzbzPrsFntcmXbAqhbsa
baMOCHsLo35yhhxEPNwJDe3OJm2hKjvJ7lWwY77Cw03wDBM9+thLosf48tqzpt9g
/2e7PfDBxnBEpoFACAR8s+4x4QFCoMOA5oxq0x33JPA9kP9tBR6H9dMXMHniR/2t
VRZ/ud9ydv+4X3L6y0JslTYxb6q82k3OP3s1CcAxH4lMHfHcP8lFPqELRvc6a3MH
1jpOXFQW1NFMI+Ik9SYUxyuU6C2pZgqoSjojdYFXBLKTuHVc4vJaw1+ll0OhJ2Bx
WasBKFMy25AMIF7qWdlKYe1sXGVWq4swcqm9w+zKrnVqHit1mJYQlUsdwq6KjnGS
rup0wq76mHKA43oCIAAl0EH2L6+hN7GOXE+8uKd170FRBjaV3y/My5z076fnOOBb
ohvoY8i7+t2EER8bhnOtlz9opqu9g6NhQ2M9a289Olyf5jNmvxeXgTaYH6GYXIKP
Bd77ATUJBcLPyG1hSxFZBrdLD8t93c5N9g1HlGVz4NPv7DZ+pR10mPCstMXSl4TR
L2cADpudZEo82rYFLp/73Pr8SjhvWmhHlqnUQVCPSKH2rd6DTmBdF55TEQ9Ueh/q
YSJRveZ+u4wY8Si7Ik9rBooZKHqlAr9dLU6Y5ENpRJ4ChZyE/VKMemPpO04UyBJx
05Yn/36DWr63lgJ13dnso6NbOsPuaHuobUaFutBztqcnS1ri9+8q8vmY5B1jV3MH
8AxiMw+HIUwGVt4+Gvz108ZTzA0qr3dQ9LcR/O9wh4dLnl004dk8AX38eIrDJL+b
j7JEXjsqwfCA7jr6lKjt9JSjKnToPkLXy8cW6SmP244nTV0VmIdmmZPbyFWaclTt
Ce68Y9byup6kQbwPBi91iLjYCKsECesV5iLtifw1ZLGL0gy+qTpCuhqzszSk/w6W
1YccnIrqau9guiwR1jZ17zWHTUN6dckTultcceWVCs/7gQZWB/3PHEnfBZP2TGhX
Bi9uXDH7RWCF7WEuDscQ90AHVTGduq5PFqhDLOSpIkEsiyJ13t0oxaf5v/+BPFBC
VZ0/wh7jSoyJsBYWzRILm8jQSTfT2UDlANYTD3D4CC9qJe2vCnX3JTm7ZPV4j29l
wMj6AX4rmrHihVlXjNKcXlMI0nuepbjjEgEZJ6yz8uC2ITkBv0YVaUWmC5BLnH62
lu8lwlJm1+Jj+kI9tyi20BkXzZHPcqv3ZJUFwwh+Qxak7Iqmfp/9r5oVi0xw8pOM
9WObpgJP+3Gc3ixpr23HQrs7Zc+rYVkx1lczdm2P+EVz9hr807S3Jys0FqPv2avZ
7S2WI8C8Dn+TgWiycd5a/3wP/Q1hoP++JdHEoBp/f9fJ2gBs9GzOyYVD5JPFN0Df
nAesh5WgMmDW9jvw3scFblNkgXUQj3BrODIfcZxqWjPBeUHTaDqNuxCH8NTzcIdh
eU9WnwgSofHpsI85v2xOfHorPyj5pb5g+ULCabozYbp2knGWlJZgZfAC7q4QBRey
1EsiOplynV+ZhlSmbbBuk/RDS/F1oXpGFrWRZGghPiaZ7Mi5piU7/7sih8ujsJXQ
TUHj2wgAzmUkySOViMud3t6hZgXaolVsdt0LLhuBprNePs0etyWvRBtdelnoXEOC
hEGI7jPC+AiIhtJ5R3ugdzYphIPLBrqGGHOHCwFHRVNMdqoIzD22909iw3ubn0oS
rVKSpC3vlnWOKyS7h+cLJAafKn5yWPzGIG0jVsMqEaBAdv69frCdv/kBFGvm8wYj
hrwhFf/h3b1+Pu+VCBjJxdQMRR22vnX0ammp7eTnnIuFkFNPaNTdj2d0zivet3dI
lE3/EknDVSPyUyx3QpZ8uoyZa9Uq01FIUicI/0plwfwol3Zlso5f3NsrsXQFmzMI
v4Hd/2DgOUK4XFgx355wDyP8rtjPh885028CxMkCyRurAiZ67WQBUzpEu8Z5NeuJ
G8cR3Dv/66Jv2kAlx+wdWIvSeORDF+7S/ET7QZHHSoPc22HQqOnbHSDaDvIJbAfU
xSEYQk6FgUipKWW2iBeSSLy6Hs19MWFiOzbHPzc1MaFGIoqAaLv0yhKk3j8Nzg+1
p2Y4scwZ3fxqigM+/eE/pU1WM3vrbMkNsO/GJkHPyQskVpfKOVg2lkX27eICbpS5
8ergnhyVq3u/vPFrB+QoxlZAC/xvI5SRljEh7bT5fak2BrWzneQTZco86/3Bd0uq
Ts03yD4ZIHnuk18X/PD+pPbYHWChEnE5whfu2prw6z2dTiWJ3Vyt0fR5mOSl/kG9
0z+0cHKYznAhLCAYzHwOYpXwyG3LofZwPOHEMkcmmU4g8evrgXs+EpR/CVZTQMaS
rQHif/Q0SGInxegzHVXvcAnzbEGUzMuo3A+zPjrRlql0GnC5pIyzthEZLxu6H0uV
XjdISkhQn0/PtOH6xVC1TTFIcly2DiOYciQVxu/2r0e4lSogsWeBqhnklmkmk5Ff
wYOJobEgRxOMrmIhxhLe5dGrlhUTvQEbe6NRWuvZNdBFlr/nVvTHEBIKwPYFh3UR
kzodgM3NI8iBqxGSxfPIb1WUiqXmzMVNyV6XKS9eaL6esNcZBm4NgCr3GqDgmWbL
1BG9GEyFUoXzK+H71wxzSDQIalSE9HaQc1NSpKaLp+uWf6/GkDrtwc+EoIlFSy0f
JN+qByEI8J8bSY0vujhtjOq9Vk/MN0r4Ju3q6bbnrtFwUc7Hq0gDvozp13ObBhbA
gvPZ4Fzh44wQWfFK5OHaIANixZbybKH2mXChewL4ebGdQJTaWlnWZ0eb8OyBt6jV
Y7AZbc42wiHnERsxw4SCzYG2uhUEUIBgEcEzQJzSDY7Og9ZlGpHH95VLteapEFqU
VY9afFK4CmimlMCSlNNEu5j2t3hX5RXfjJ65VKRj6Yo8+AvBictqIKna+/Xv0hZQ
7BWW/y03HWsku16GysYFrU49JMyZbq1TiTBnYzbnvvP1sLjLpP8whqf06hv8ferw
AHW9qGnwRAQeLwYOSkIo77e+AXMsikNQvHEttArkcrqRJNFlp0wUkjdQOQA6AAy5
JEohj0lq5CUeuAICPlMmEC9OSGeXG8J2yUQTR2hRYDbsqroIy9SyDIz5LZPpu+z7
VwydBmnZn1lZCbYIT71SBooGWPJFgnyN7MoEcyQ1e+Mw9DlLljVWaHvvRyJfNn2q
fOQVpKzgUqUjjInoLgkGXixL0dy5odch9TPHFrW0LgafrYbJ2Hsxc2n4xn/8qGtu
ephI7ql+cb+LYDMpOdEhMRFH+lhENiKhSIyBB6ej1QXTUExcpk1YmVpMagWG+2aI
XpU7o86FFf5YNz6Qgz6nAHPsXY6cIZgO6rlByPCZEXvodkNP6a63Nr05+IyKXCNG
E1NNMYb5p9MHkAfuWhp2dN22ACP7ZDYVEi9vT2fjZ9ypV3/pt97j9qjaX3SqezHf
mWlvciOB5zM6TFtPa2JPS1W+OlkBFfd+v1AD3rGS1WDv0o6hZMSWP6fZwmDuKPqF
JtB+YoEizlUptovBm20ScBhk7Q3A0U4kdnltP9YN9j3KxaUOo5vzlP07EYXw8cWr
X370mVQycWygwWP+JdauCtWQmcRNCSw3XM48As3XtiFnSbR7cNvakoXG+zA01gaU
z/p3sGLLJqJq3TwtLTvLWXTMHyHg9fWKfw+mhWjLDxiujSjH/7yMyV4VDvYaq2r5
4rtuEc+ZnBCHse32nJCEMnopuo8pt3+XOK8ZMKF+s41Hvz5h+MELWmiP0fCLE0yR
1S8Ej9etF+/i9hzmZBJC2BQZd8wk6TW1Z2VF/NjPmkZuISYzyoEUwRJyuuq8mGC3
QmQrF8yNpelx8WbCcz+lhbp2UAl2d3PmK68USt9SwsZbWKui8C1Uo92UiaAJmbFZ
v28U6PMdqgPa+2IhLCrITqDLMF8vEEgtDy4Rm2C1+5O8B09WTnaEXXLe5CpK2liH
j83041+19QH/pKImYieGMNWWxuhpzWrq8dESDyN4F1y+d1ahV4p4sm6puz4HO3rm
csR3O1YMV1VdjrDYccb7hBz/y2pyul+ANO0ItiGOA8dsdNj8vaSGEbsfaP0uG++9
1EtJOwZexFE0z4P6QMmGdSwREM9KzTVScw3mHPOf8h78op9FkManRbKVr3B/sgxp
r8SbHc4OgwDhxVHc7j+fN4O7E9pUOh1mVny7zoMgxRF6NyrwPknah1y8vR7VaZK+
FsNQJ8SwOHo5Oee9WdC1iYigLmgeKDi/YsYVXBBdJ0jaIXyEVfixUO6yoxUwPj+M
L42ogZASjTJ1r4fNKSzE0P2g5q8bCnF1ZaTsQ0ftKns1AJ15B6IMcF97nPecyniE
59QZwiJi9t2FA1HwS/wBoWhpYxSWTm6zY61z7X1EdKhqZNFSiI2+ek20MQtBvpTe
7F/Tzt7Lw2iRhRiToLuXO++/JbVwbbQjiml0vNSu5a5XiZCnK5z2fQ4fH5+VEv/B
ouwiGqhPTT7sEyyMI3bJwTLr7j+JdZBMj3j6BS1elJGuoUGlDTxiHIi2w1Agde7x
s5+tPIyVNFIRWlUcEB/Jz7mx/PKIRRvTTNKd+ubpKrgXItfUZExEHCRcylu1mXbr
/W6Z1QXzWJd44jtZS/VGFcvvQzt30speKlZ1mCESLW44mhm0/7BOdW04mcxtMQvc
1It5nsUCzfAyIAA0PKikvDGMnoPI+NZsSnDjXJpJTsVG+5Cx4MxxUVOZxtbCvmVj
9+Juw/zhV5kuDh1pCvAxm8s6/MxSmBXeWO/59cfNHhO5iKSXIYgtv/lLa10HHQ+n
kIcGQonATHvhYacX7L5WE7fhNkVe2GAen0HQosCrGpf5sGPEBzhy7nXoM+pr6sTZ
z+OiRCZ6H4gx5NsMeVzcrR2C/s1qhnzsKhVyHw90+6y/N1nH9AGitOaumGRF42K9
QMyKLgj5DmTFCj+F9hhAei5X2VG7+fAMQZVXWhMVxwP8YwZSlvCz1GspJ+Y/Zd1s
VEGF6Acwr4GaZYsIT8/mH5gwENZ8wCUVLEdWGBW/xGMb0+y6By/T9HzLUn+3SwIe
mn0DasMmBQ42rF7L0Vg7u3TtJSgfQrtFILQdRZllvghNIXpfGfTZXj3qRNrm22i5
uWqusMmD6nBTqC9UHM+Rnmhyk3IlH+/LO5JUMC2HOyk8dR/hgF5UoaaMECv+eMti
6VhlQdo7xRd0IoVZtPAfs6QEkEonUEcef9UtCfwq7ASuu0JDecnp20lxIxhuP2wS
eYl6nYtD0MP6cvndMdeR8sOjDEQJUtVnFsXNrQHdI23RxMWuRFMGkQyWcPiBSJu5
nokaMiF/lsD4F4/uRu/76jNbV5AFEl1vSrVVFeUtydd5DAS026NspKNPbEkqjbA0
s/W+LW1mZXLXjczwb5izZDqfDt4/3AUb/oyEC+HXso6tjaw6u9/x+nAaJ3iV/uXk
PiD6zB2ybCA+ZCH3zUf6/ia8k7tf+r0hIxgXMqfgSQAHOvFORhAbXTl8XtaWKojx
6egBx4v7sBHczguC9yljZNBc06QvQkrvLVTT4em3BZoOES6v27GeAS9TJN1M5kkI
P6PGK9YLnULUvCjpElgQ4xuSZz1kS1ZfLd1dlmOndO3lppFOyofvbpKNLg/FI7mS
yMlspan9NzodyfuD7rwSvKb9CeyNCVwJFkU0lEOTBRlKtRkbn+ZFjuJiZ3fMKvLd
wz0SYJlUizti+1wYxVvCOCxSdyc5nymvBzK37oYr2DEUCiZGak1f9SiXed9l9JoI
eGWME/jfOfEi1lG1qiO1iriH0gUKw3XsP4RuYu62jUZy3bgPS9MuKHE6DaPQ3qEm
OWBgKdmJz9AjwuRLYYa+pO+sjcBVw3eYoOcvU+ORu+3pgR73i5MhNU9YDBZARRVJ
h281+/H0NNK8URiRkMZofAZBs+2sR4tl/4uqHM+wfvKROIjivxkwAVjGbvtYXho7
w6JPN/lMiDB0Dlyyk8T/DjeaG0zQxngLOvqGg5gVTe5bMsx5WflECjAKljqK5iVw
lgg4eTlDTBr0Y1FBFUUr07fHSogR8Vkv+QWxb9hdDZIkvW89yK/lGCWnqOuusWt+
2xAjzh0z387a7ehU39Xh9+Sr8sNPX5IJW7x80KW4OBPfAef1G3ECTMZLzLk63ppl
ADVmRx9efeC7QDBFiS35vIErZ9zE+p/5kZTi6JheaBn/g2HV7XhI6Z2NAQVKZpa+
oNnG24l82ZbdUC/GKTYlWUsls4oL2fllORnwGXuTNQrBWIeW70pDp6C3wwuhRdf4
0+nfpj18GJvEO6Y3GTXda/T4p8IUpVhAsm2nltwbqHPXRkXER/0IH2g+weUvX4n+
08F31tG3OXoqf92bAlFHFOC2E8tz2eFOThETwMw8FybrdOivGAG0XwWbYuHA220N
L8c5dWDHhIjYNeEMBCr3MSAzVHBRWbAax9AWb9p4Z88UzE4mOu2ReCEXFHMZJsVI
OcrjpeK6162rtJBbQ/obsQTsMfO5CvOqJTHIaJszG5KuZ40ghxnXkNm7Qu6mgbXK
IZccHNVj+B1/uEhux6CjoIljZK0Lw/1AMLcyNyhYpvTzFG8NOuBasi38iYGXa+Zd
2neHjDMlrmmtgOLG3ktkloP3h4kIn8yAf/y3BZLcTL3cErsR3Ip9yo33B7xsymy2
31EP8P95LjTBEuSRsgb+4oC+LppGOakwbdCANXNwkp/ypueaFI6lalocJ/OwHCuu
dvP3P8AfNjgGYXUslFqi6NtKkafyjwNfysJmQW6KW+03LqPygNxXEqJhtSAqOWFP
jAuxg364q6slffYjQ4FVWFkoqkD1E8+luIMxU/zp5TYQb7j7sBn/1kyXafmt1R+i
4o0ognstK5E6vgB6vmVXkY5XdIm3grVeVCLjTRdALmmuaWOKY7a4ggivj3AAfarI
rE+oAGUcyyFUc4DKAbgIwo9malrYIWuUJe74zcZmTViR/Vun72kOHdszB6Kq/dBq
My8e5VzwhHykpz/1SbkhLpWG8z35apLVzOVeST66UGimQOwCLhOlqU+YAJqVvW8I
dC35iTr3sr0+ZPWzLUDV9tOTCs9hgsiEbabP+/C7+dIlVn3V/cLRJTGYMmgExhfh
Sg/RsZD7a7U0271jU8s9RhyEi98LX2Q8fr1eQojtlCiAZ958NmaB3sxdeM2ZCEC9
hcUSj/UsBv5gxdKqop63924dupwx5Rk3JmaK3TJa0pNL8c5cHy4EwPxfyJ683Uzv
WjFYQ6aoVAM7lZ9RKmHUvP3HBXVrKYTwPmWMR7zVFgtm4JXniAUiQ0eXxWLXs92k
HpOdpNMYJswQge6rqUj0iceux40qfIrfjlLOdbJ9N4tdE/zM+k/82MmRXoOJDP4o
WqPwcBsHK2y1iLv6PBtPMueM1vbVBacQBXgiGRW27o7t81bMQPj1pjj2KxEBoG14
ekoaX/4MXp44wOwat8wagmIhN0Rm25CJ2H4Al/IY1O6O9fqM7CXjH6+1OqnZuWmX
cpAd4yq/FAmAYGL1TqUF6+vtI90T7ipWHdgO8CVXQFF4Mek3LHVTxnG+flre81vO
wRw2hpfj/hnQ9vuh8UTbKxSxw4Mtc+sj1pTNU5ujztDtoCg9UfZFEXcssI0lAENP
BzzrXYnG5qJflXet3qsRaI6Fn7H8832T2TI4Qz1Q4MeT2WTWHxzXN0I0HhvA3P/x
vkTmNeqYtbrH40RIHqsIZJKpheiKHQiaIIAO/o9dvkbpwbEW3xv8gsn4AAsywGVg
U6MBKtYzr+T/jpLJwdnhMVNTDcuEVDxtrcg/ENFNDHzfIwWVA41dB3bVZXlAAt9N
oVZ4Hhmhrw2x8LaHoocM2cer+WmmhusW6XYBr8/XXiDihom19b9MUCaSXNsmQ0I2
Cl9BFnw3RcNYXO22AxZRLELq0g9A1iH85oNvsW2/UmOQZiyQp5c23b7DCdEeQic6
buqu6ieG9idXoPBgM6Zm9GWmUKG7yMDuluR+mOXq9Cq3Dv3QVwgkSu9Bw5XOJcj3
bKewhKaXUvCQthXLodQx5aDnT+1/BLzHpiMTtF8S7fSkpqEakIkDl5KbVm4bUN3K
0uuq/EL3oKZFkSQ7Dg2S0T3JOXcjt+prW9Z/KQYCe7WfkbnXrdO7XwUrQ9sGrwN3
eGIHT+pSoLUEcNnA/E0CuwpKXz0s1fIEF25rmhbOadEYfw89CS/VAy5qUar2oWgx
ZDaWngrfIXdBO0RsPQdOWVffVRMRGgmoPRdVrJia/Y0eH2pk7cV/dRaQwoQXMIda
MLuzEzruvUSm/u+zYMQBw2F3LmDgtmYIoZnvvSdFZSdPZDZ/wI0efWTaRKideKL1
wzwq73p5rElyiAWbVnHHoV7pI7zpZbsIRCzrz+7AIA+OMF+y5kRXbwhAWE2ff9td
fDzM7T6NMq9uoCjO1T/FFhiHwi678JX7AetqfjT/zP99UTK8Xdk0JJ+PNpBxVs6r
hbSVvGBZ2OWlzP2xjj1jAxlSdFG3VrlWmVwMB60g3/RrdAJGX2tbOqmQLHeFdx9s
kYc1E9n/1S9HhqTa38v6Pv5RawOnlmX8sbxNpi6pSQ6J1X2jdT+8kzBKqSPPPA1+
af6DHeguT7A3yeUJ8p39tYztRH3JF9NG0e22REsSw9f99+dcYV29hloGvOB/tOOJ
DEbuLEmJ7+la8eo8+y9j7YhGGigCvwTuLY2Zp1m/yEvgB2mR2bTcRWU0tVc8JnSo
DxvaiR1507tdExA7uOVttDR1V1R3EAXN0XFB1iphDlcT961BcmLDfBnpcAIJavKn
j+ewiOjhQPh09kRXZ9SGdZac1i/EAKMCkS53KYqIYlbhppoJJCEX/OtXrSzHM6aY
cXcSITxcrdBs4XalRArCSYl43SF6F0QpUpF3kZVKCyvlrObTHGmUCMVFoq4IepKG
p8WeVS/6UAwdYaTV6GKB4E0pOgjk+Q8A5sOB/du1tasVMQWQ5/7H/kr7/8x52Nrt
A0rUX0tZ8BTPXgMbCo6WzZMrLORLMdvcOCjoKq3f6dAJlalbORIoX+qq12I1uccC
bc3rhi5lyYogHWTBRtL2BhBa+tfin3mx3qNgEb0kW+W1hDcgy6mAdXT86Wlhv3hw
Uej3yl9XxfyozDb9TYwLzWCaNlcpOjbYmmKqG72X0/meSJr1fK+o805BK7O7R0i0
b0x/cU9KfDG4jVxEVCDqWWy7LZYl5tK3IOXshxad4ILQMN2cBrPM5O8FeeWaV3ei
/eiDRyMJ2sHonFmQMmR2RkFtNkRRXUWn9WWPM0UlS0gn26dy/8rGl/s8a9skcGUn
NX4iqDMpE13pzQ5Ci7ui97cl8YG8MNVcPkzDKr+lbgCti9N6AlhyHRVE+VZ/rT2v
OwMO0QqfyBfTwuQtBDnBIuNLWUuHmHOgVHORq1rgDcxuEHx5iiyVwmWe+t7GNAIb
aA8qUY/UvCp6F8R2xPSC7fDYuYUxWZQP1dB8znY8xH9uYOBITtkT8vMx7e+5izif
OS4k3d0FnxHKaCu9KEeSKJ8glY/GWHlqrepv3Q+jEdhex40gXZIPXI7nYIdVXnt/
0gytQJYhMOOMjrrOFvYfiiygnhimDimK+wQPS4kRYnG3Iy/XGC0TV0GzFa3aab5+
1TBRejFTT1EstsTUx/bcRv1ss0/WC8zeM9TitMqbpKS+iPpBswWCcp89I8uK5/b8
CbOgbFd3+ZGKxeYd0U9GT3Ho8Xfwine8oppMSdgVOFUxThRvzku2Aa3vX6KCwva0
bOAbn2gBFB9QuvpPEMXoDIZWkqO0377PwKEFOZPNXyXUcAtR2zsh2V86M8eopF3k
pdcT1M9h17Yq3NZvFPwymwZ3k83GT5pyq9k7Bss0oQk7ALqU9PyC/8vNcFON2Kpb
3JL5/4wxQ+jaQ70AEbGO77xRjYclXIdcFOunYKAm/8xN3naUG1Ypa0fBUl9syNq4
xJyj6fqxQ+2LzLgyrbnIafgt8LMLfPFFLYqsFglA/1hj64qeCxVDkH18M2XOkDOg
TXGQl1jn8/AkVezlY3MknzHRxwF+v5Tn4oC0om7S3aXAejKeqDvLojvA2scItJAv
uRU6muNqHA+LvTJ9zWnbffubD8ATXhmGRts0/57On0M+NGVEqgEmo82zuok9IxcI
uArS0CSKzLSwTBGe7VXLrI2dZyWKxKLpykOil0dRUU6C5yO+4z0YkuC+W4dWWDi7
RlRdfdVWBOoo66NVPZMj1OOich2GpIJ+7/SaHyiD+FUekuY8ax8I7HuUrWLnqOQY
8uuyfq5gtqarOortjPQnUhb+jnjvGYuKj3ZQ9WnpASDCHjpTuALqAmnLXrH/X+Wm
E994SiQ+fdpCUS2I435csCtmbIgpPsT9i9CmwizAiVy44Pb5W/m1A9IjPUHlxdph
x9DMixRCjFaloX80TxJPamVif782lCn4xcc+VmfLowy9RhHBVwR/KLbddDxBspue
jRsUJimDNEwtTjNqr8V1vkN6cb073rZYyMYWreuFI6L1dmbcgzedaHkcmBQZ258i
gpgjqCWdMwmxe08azvZnXS2M4UBdtqI9zMiKSLu6wEoJMOtTXjf5UM+T8SYXKsPo
uWaAZ2bV+iUgp3icVZW3HYPAENi0qlOw8khQFxPI2hsAFTSM2pAdH2uLDU2vXgzF
ntjoAsFydGX4ZmFHlYjFK7pOdRXPAhj3PcTS1V4LTusQLABBfScgRoutDiCIGbCi
pwWqJbrspbcTu0jcqoPKtINcxWunf3e+0WggsWLY2szwaDpIT2UlfXxV/3/Kz4I3
CqHDz1cokh4TuF7hQ4UVqhbEFRnhTjevGSzhV9ntGeM=
`pragma protect end_protected
