// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:02:09 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Hcha5xaOTLyyC1wHuZ7Z6Tn8+OTTRHXZNa/arDrFdG3UIgKVxflOD9arOhFg+Wn4
rhf7TIlfeSwaSdgi22BCx9cDjiLAs5upb1buznHxS7ykTUg3oCvab2OIPNw8zmih
CdybP9DPOGyeyusuAMEuwBSdcdf4sYwZTo0dOpvB1wY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8416)
dyDKtocdPV8VP9Oj+5BehUQnhNSc3bcBFJcUeGWjCDhNZt85KsX/oI+6emQIu3Bh
pTkUGUUpbCys7AmU28pZ0TnhWb1UGG84RVMFDPwbEtLQoC5js7Zhd58nST63//f+
xe+rIo6KcHs5sHLvkbJnmC+N/JhFEgKBEzMACbRMDUM4cq13kYxk0eLREkVfFkAq
smD5XGMmMmhyIcFJ4BfxzbgSTRK95wMn1CPCWBFuewB8kOI830Xw388rtXlufHot
h0W8cdZUz8mnGzo3tg2yNdL1A4QBI/4r80Z33pIw/4peZnlbyiSbEbL3DXKujflY
SZueq0MsOx1371RcIfK4ImqtCFEUonHZdQqKi/8k8NgKflX5rplcdYGWR4/J6qye
AA9m2eRw07ZbWNkg1D1cAuJtGOCMIdqQOSmRC17Yzh8Lz4qCu2XHF58+BlO+yXoI
R/JL32jV3bNuVWJkMMLRcstQdLSR/uvp6lb71+aCf+3p/y2l/bSVH5jrY1WcACBk
USKcqTofihrHieZHtOjheK+ki1JMevg78QIhuZYggua6N55sd7xW4UdzlUe+NKdk
il8qnQulso8BDGQHVFaI0QHmhMedvmp6w4awDNtXazKhXvDxjgokU1HIUnXFEfUS
mGwdHWKe3BxvfR08jRaGhKFXreuyCTsWTYZ5GLHm//TvXWLMpZkbRxcJ6AZwfCj8
JT6c1gmJ0CFlRdxIz3QMvvDtQNmZgyJt59UN/TO6Q5NypsiFI0seA7fO3Lrx+F3j
JC5yQ6YJT0PIgF+UCWrlPYPJNLWK9zeH1SQq759ixY3yMJpqwedE5avqUn1+7Rtk
4x+/kYr67W1i0KyRtlBUj4gohzZS4LpJVbr3/xKXG0hukXqyfDkn2jKuh3YX2QL3
fxqQbd8Hn0KMXIWJHKlMne+riW5gNvhFUWrScYHep+SlZgFvDIw3fYkTTipkkULU
CuFDUMruk89Zlw1Hq2E1cmUZkTCKug2DYs3q5puqn8knX/uSZAUQ5EMxTndWOWJm
Qw7JrOEKs9UJ0Vdsg/LcHpLSief52DrGWaWIFOaR+onYgQhhq8AjYNJLlm0mgBxd
78dBwuwwb7umTs4/b3n8qVW//kQrlnPm/hSlK+ec3KYTrStzBUUZrmgqrMN1xFVB
68kCOUfcwNlKlK/iWULQ6BLhnFgt3gv4ly8abh0fuAafkb7xZJ52xfqj2pNdzpYl
aCajfLCrhLQEtFjulwnkLg4HcvXoc1tdnUPq7OpjKXllXzyV7eN6xF5BXN6gN8pT
c+hy/j3Zp698mj+g+qnh1LnVgJzn0t1JAy2gH5YL0UGhKIkIAzPgV3rBrj3P4VMi
gIiXzDo5rUgKFwooArrSlf5RC2ZXKUlfV64EdUxdIJYX6CQgG2gf1KnOlw2U3BoO
0jaVKYq02H5aj/b7K6U2eqTPRS5n69QGU3ZqTb/Zz3+X1aTDgS0qh0n+z/1CrniU
xyzf793glonhb4hMuIqE18bl5Xzg3c7d9rIBTpVTkDVwZHWpkoy9trtJo43nE8M0
/8AO7QhgKtkk7I83kJ04c/nhFy6T4wSrf6NDgbTMK9keC2lwbEqOCii1xKI9HDqH
GP3FsAoM0Rw4zqTCvrv5OPWUPyaGSc4Qd3oBvDaAWCjBSxd9AfNejaAgEwUDm1/y
HH4jSK3L97/JpJu/xuDRBqdz92NWg3TjZl3hkKElu82nYE9413+y1sAiujh89cJH
J0E3Q6ojx0CMOdcivHw6czixzjO3bT5osKqSg2+DUY7tceX/jwzS2AjaKgYQVzto
e1KX4Zj6fstO+/p0Q7HPysMnTxvrIsKxHyYLDh2IefMxR4Fmf9PtcoG1Wag4GHZM
2XtKy+qyAWXYOSbrZ5neXkphJzR4SirAAc8Pte9TPIAPxAy9NC5Tm6hTdTWLfupt
1OYiKOgVcDEse0R3rJVlE/Ffvs5A5JW/Tpp2gKobYDQTN9FLqYPjiK9r+wWsa7vX
2inzndRh9p6A56R8rP/yrmB+yAJzbdLb3XambAteWtaTnOhW2a0MQNtEpf1ZzcjP
IpmH3mAy1XA7fvJeyWPYh07PHTlF/tvmNgbgR1uNbwbypiMri3P60wR5z98w8+jL
kpzcOpymZi8S3RIwDaqveqb71IQApFRNXo4114w2O1JL92CE8TOLkhVS2kIWN78y
ghnijiPlB1znQpyMT4Kphy/8ynSiNXz4RrUtcxHHyEWH+wCB7EfTT48h6ixzxVjU
Y6AteDneRW5qP+awEOk6zf9U+lCVCKTK2mYjw9HVFuBTepN7MPUxLznhmsPVAVyD
oXDkGsG1I9pBFRh3vfioMtY+bIqamlkCLDNvBDzYJWjLGv+zUasAjryngy91lWb4
F2EMtzRpToYs59ScFuakUnPPFOtk6NaLjmJ+CvKdHvS2E+o10um4+ILqjlJ+pcF9
cDHPa2Su1JN4Zl05eszGM5xmBSZAv7L5MMtv1pk16v5rCEwEbYXAUXA1/241lRlQ
uN7PAHPB2AcnrVaE7sTZRJcm1QyvJl2dWFkkn9THS6YTDmJKiasMZXP8fR/Iofii
g9tVizYGCCsO8IAAE25/sSsh3IZ5O4CovqZDB2bBULJdw9gcTXxO7I464GYrVi4B
wxfVUvvWsg/BdKZ07RIRdYzXRHvXKUcoVmCPhCabGIXI7DmyzcXWgV6up0zf37xc
TBrYRNPktvNuyGoaHW39Sys6aMbkGe+ihzzn5reM6gQWqwjdmtJc6S2TIEATbAgR
lNpLYwYOosuMEMtFBz2gK9bOFNSBhFQ+8Eev0hYx1/OqjG5/Fod306qH5zZk5wPx
0XyknZi+mV9h7OFj0R31SsSwye0xTphQiAeAiCOfGDaNrVXqEyKGj/V14+C5gU8m
oAef96m3FihrUslz7jTqGNEXjFRpWuzbm0s2l+XE+Tbt+DqQ2YTJYprxX/0SmuCF
QVaGwYlTlOhf5im8ExURi+rWfR0VPpQqwxLQrYuOxLdkyTdiqTmo1XlNAbOlgFMY
xqGZ/exhiNLWmXEVDhIbR1A3o8HpbhdUbkgKeWP6bLazX+6q2S4jFKodjF8EY0Ed
/ubVsjREfDG7ol1tideKdCB4GL5v0TKkIIPhUZbgpPFtFp5kVGKqWVkiQXvIotRH
AQCOd6AMkYTG5cQ++J/myKCLp1yCzp7nzNDg8Y6u8NJYjGF1qKcy9S4ObEjpLoGo
xUMoTKt3HHToVpObTBdOFkMz53VxwMUl5ASfarud/myOlvALUT2odLaAJEkkfxyQ
Md39J0Zam6OVjs8p46E6YwWsFe4tun4wgwPo3/McvIB7gC9xc5W7Ibwcv4wdci5D
954b07n88AB0ehrVHIlPTYlKw57agfgapdmxOhsNGrQc8hw4hSratQmMcvq6Njyv
hfdflxriRpSN5wrDqZ4lB9gJjeQBXWoguE82UcFvrIxW/bUrA191Wxsv6YysjtG+
+RoMWCU0yHDJCRqgqYHmztGru4+WLuKhXNWXWxef1XASHhT1cxIim7mI+bMvS6SQ
NQWYxi6I82wZoR2aCjRvAsxpfyfMMFnIIkK7HDZtJyNkj7G5oP03HqfBA9TehjFq
PcXHm1sR/j8ZXs8T32FPQ+v70nauxDToKTUprC5PNw9OVQYR6O4MfGnXDHkFUXwF
IXbXLhR9Zay9G3qjR0uDVJKY+xXoXcescFVOFc4pYI+La1PYMm1zGsIVzFI3r2dP
zW6I6cFC+aXkwb1kqHtNg0R6QEAgvDp5BY5fbJSSes9THEkZEbuc8xPjRyWKsChb
KN1YtYmpasqXgaus8L4U2PmdKMkQsNQZ4eFI5FWZ1tzloIGlgqEbMQov7x+E6rTU
k1UA0pKOCXA3doA+g/t87N0piSzzYUd4MiPLMn7h4FQmz+as4eT/gTjMPV9yeYm3
thHHovJM0cPs+4M8P8WarVxPKIVInoaAzcC0/IapgaGaK6bBKub3RQugtM8A45xj
+toXcwyQ1VVh8UWbkinS6nOr4nP2Al3GmhUuseAqh8KWzXQItoIi6Raqn7COGsmO
j9adktY8DFxmZsP3R51qaFgrpZEIt8fQQak4XFyU29gGLuU3nkO3G+EBjuwJv6Zi
ya1f5DQZ1usJcok+xe7ACDnOO6EDPHs7mOex6RrIeGWN2ud+DHf4vzFKw5eUT7C3
Vx+10Gp/wFAgWoypnuCpZ3DIqNWQUW/e3OzeURvcJIqaDYrx2Vu7Uj0ZuYkqGZBe
RKKx6Xmj/vnVTKxu1q1E7tbBbw2EjYQTn51iFTv3wwnq2GVgYuzB1b+eN0+hkdbm
2hoRW9j8T8cSYOe4xHTiIyDgCPRz+FYLvbg6Xs3NpUXpM5mICkGTt7veEcviw0ZX
Alwr39wVIIoDMaoD9QgAWwTQtJotENMMWQ8eOVOWgibnVRPqp8r6rrJCjk+4Nf8E
oUw7Qu/kIuCysS0gxrsSHi3aCTsJupoDcBRzhwBH1Q7V3HyTd+gdp8zQQwLgU0Ic
ikilJA5QvfBKg94DQdM0kueB3LUO9a8TWgXpZC4R2BFD6gcAubdwcW28PD0r67G5
7KlxNVueRVv1XIXRCka1nHhyF6bbBU3+hS4M8++UpT223t3zbLsjitY5l8iM5Jxy
qnbZmm8efe+h0vrm74ohUheLTDA3Gx3yqzAYVhD2B8Uw2AU0avNmh0/piCATPav0
pwmGbNUNTB5DfX+t6eqH3oBdLwpeYM7pBhhetP3PaotVHpg3brFpEVhASmWd9fTJ
V1nqV4mTlWHP+JkU2Bj19Pvj2FoEWm3a7rgfyl0CD2ZzOimPnaUDaGRnQoNQJaFm
YQPJmVM0zxITK9dM1YAecTI+PalZ3CFvj1v/3ehnHOEUZfOwO34PKcd++CYsTydI
dvVJ6DBOdRwHjeQRCMi5IPSlhUmS7xwkzDwBV7aGUungY9v9wNqVqVXSCQpeC6SJ
I2Z6bMT3H3sLkCCRjaR2GolwklTRaqif4cdUhYoLUMQ6RiyWFD6wGrqUNSPjMCSV
x8SrZdpAbggXS9cX7aZJe2AhPB5lAHlIQebkAgoVtUG0/lksrZfdnvFBPkd/4CFW
Fl9Yl0sgv1llEpcLg+gnjO+LXkISQ1A1mEUrGE6bIhwakRMTXocd3fWt96Usp7jr
j5+C5cCxvsSYxiUxyQoZTlZKJ/GiYnboYFwJOcf2O751uDzF983xEF8k5ut94+Qt
1y6AbrU9n99itljsM/hTxegYblZ9KgLTC694b3TTJDA5NvOIGSmaWzHfjo8u2Zts
/H75xpBIeU0F4Jb7g5iPz7qKbOenvXkrVp8xP3ahzUIzyYeHaS0Cftvwp/gznVWW
KYT9E0RP4ayuFOrLfFWfEpkLocgqaij93rt51xZxtJ+R/6w5+SF6Q46PWw/jzgxD
y7lmDcX+3tn8K1YZlTFJKv1DG93kv2IzNxOQDclxszmpfIAChUAUNAN1xeqUvMG4
syP/3jl7CAwvtdfM3HZptJuVwBGpjBMUygQuhTJArIz9aqkLStn73u2MtC7V7eqP
ajXG/wsWMZuSliv5H4G4IoRlhlrzRueLstXhjyyoUtKIKl1NRu7ATia9Pf0AOFFn
JuXj1boPNikucV6rkYfTxWTUu5Edoq50/NyNr8891NlQqwutcv4Oe+bm8aui+zq/
kUKEm8EjkGJO436WOW0yOZDxQmmK48m1We4FItxG5IPqtnoREman6yHyMW4f340I
St7RHmufAtzCm3VL69j1pOble6iD5oGNPdy+Ni7ymFWQM3I5s4LGGr/q/wnFz9nZ
LfQGzDlm/qZ8Ou/Mk77U+CmdXDaA1DiiYHybfW1nf9jcxrBiQr8EwV04RTHr06vD
ozfWGcIMlL6EQ0e+hXIJ0ZIokG3oxaP/atAceNlRL6AGz3Oz6fIp5EsM6X2C+67x
VItqrXl3JpTpQgCoINU9P1nbZQtfpHTvE75IUZrSBeKe9iUVCoKi6o09mZosWgOf
q/+2jcZOmQVQ1SY22CGZhqeHHJJPD36D/2ySYIrE62RZ9uLLcnrjqE75d0Vr3rCT
i3epqGia6NILXMvfy3IrYJHoeqReE60SZVz+fX/0ATuu8nbjqKw7lWPZv3OB+5gS
VfaurfaMC7a8b44gJd5iM+zR/yjWoLhKneCD34TNi2qDPqA3efNofUPrpuy9AThf
89oN9Xbp4MaIOS/8LOLutoz/SXDHjYlMaYoyoQy+1V7rKyHvgSFeRLh1IPkDw64F
3M4AJXkK00Wbf0VJTt2pIv/pBX4L67TJ+N3CTDjapcEnZPJ68MfnCEskKnXewYTL
96rv1i3PV+MDgsUKnixmkL/xFCVySZesyf5FBP4A+j4T50qLc2Nfcp6pLWiORYkf
neQpl4iEdW/sCjWNIIf7FEoPDAvKTMVY6AesL0ghiKPffOBaTY+h/iH9cJzgXZf9
lT7skmnQaYZ6vdMtoD2ao/gmgJdF3GLFg25I7Ui0BiitUTf7vV9ThtJW7UlL7dCB
gmB4WkUfUB22sI7VYGEMvkd+upc3/SmR3EC73nXX+dfeboUETjs2PiTQW1MqKSax
FHtmsi2rAdLEYMZYJF9M7eT8INZhxFXkh7oMtQogDQzaJGt/kQyjPj28I01snjdf
BX5ycmx/tGnsbGjscumbAEG1xwsYWf5WdEon6Rzf36rVji+I4aZd/LDHdOOGzJBk
Drsav/M+h4JOguK+DRgPpX9q8C1GR2Ukp0d9lMtiM/NyzLyRhQOfKuFZoTjJjvZ4
VWrObxhvvPJd69f/YoqWutnC/jUbCV9dH95Vul2h7QWx6+wEVSaI9IyNJ56f+LVw
we6d+f8YEwI6Ulx5mMBhjF0s/bxdyxVU0cd3pPFR5QM+mJ822yw1YutuYTruDELp
+KC76AJcQeVdBQ1DgwuAq4b7AHZjTU9CVNZhCoteZ/isIImxY3u+1NN4SbwlUonU
Dg/QmCDUa+fP5nroaFdJ8uTFOnBozy0uQGU+RJe2pNTuijmEJGfF3dwVI6TVyKXz
FEhX6WZywDX6rwFQe80QNPzWkeeM6OhDzdzE8dR16JVyeXJTtBfvIuO7E+z3Rjxl
jkPzDs6UOOT4q5LiKmqdHJBn6s/5hs+9Pkl4bcuw7rcRr6LgZmzcpkb7RtMQr927
JBWXUJI6OXLTXwo8SQQv5uparvI2iP/0KRRXfmeQLEc4SzjZCVdPYeQn0jE5T3YK
nou2jU2IKi8jdKY44OIhGqeJwWKFjmADwU5j+Cq0VkT+HQy1InAR8G4W6v93HD8d
0S6cuDvULceTqneiY9SHbLyP/dHZXPGXi37206K4orqsRXtt06DVsd+jWYHYpTIw
1wb5qYDQAAKJv8VSu8UYN2YLIl+ofeXuEhQy1dsJlxO71uYP0N8G4xFITAHTJwrj
MXuFKsc5CxG1AmUSnJD8hNVAH7rGFkEs9bniTVyzB5c6rRuUckPyUWOfFTiU2UlW
Sbe7Covsn/mnaHDyo2uqBssH8pgnSZOjN91VdM7McfP33rkKu18IRIqeWVVPKPZZ
Hgz7TIzU+2siFAqjpqBSS4/F75D+Ezh1YRVgo++w0Y5OxnJI8YOxnc9ZYkkCUy7c
xdSX0YOgZEOKDfPohBeAG5RHoGQlBy/LRd9DSj1Zwwy3Dt1McVxGfww2yUJ2IOvz
1MkFE01hYjHUjtw+s95bwnKvgAdawRcc79w4tmVqhi1tQ3qRjj8TeBNry3QBQAtt
VhoMM45XEDaf+WF6f+Qsa1P65cw6IqYhCrt3dQoHCyKzz3DxWDB5ptNP57lBbPX3
gGapfN9aJFdHoWD+rUiZeyJg2KVbWR0cm12XrrXhSHnBmGHO/ODcmQ3e6ZTiw0Ng
6XNXpV0FqNtWzLMbGVRw9a6Kppohmv29FP5OXQuPGBCy+K0KW31sf95OUZzvzrXS
FV4yyRTPHmY4MryzCY0FZl0/hv9/tjEG93cQ64kApW+/OhcahFYoL1IEYi3H7cb2
D+TzNL49al5jdn/KEEuwJQ9KxfzjxsxCxd+ADwQVsCeL4h6bRkbhJssgZpFYz/aJ
Z1RzVGCyEG+oWLbtrZ/K7vBHfefAgKvCGzIgVEN5h4BUviQHwWnafII1lknri59G
c1bqhF8jBsGlA/VDEgAqoq3yVP0n6aLBUpqiDShQYsE9xvZQPT4j3kt/dkWeo6wb
y//MAoJQkgvLnrQCBPLT+hkbdZvtmVuGiW/uVBMWnk/3W8wvWbkbv4LGH2WuVFSl
tOn7aJDi0SQkNKnyPwZfaAacbcCPIvIYGSGh3dwGX/doW/iS4XVwhDEtoUHPlz2A
Svc/Ez6I86rtk2q3nbd/KZ7SLe7UHM9cGB1Gth/gg4GEpcE9xo+K0VujKVYS4QzU
BGibKfc0qa26/J30ZH84PCR9j8moLM4NO80uYDDS/CTU14zvNUxHGd4QLb/gxUnH
S8GKLPumwin0iTBQ0RQTI5uA8lvrO7wt9SoDCszKMh71eZKy5z7Ba3a+FjGqAqyj
p/8kakEBHznZ4PRsuu16ayOJECwa9ydiUdkcx/YYWmC0HQC9lFvEI3YRhNDGvkCe
cyN/nL9hcD41/9NEpCJPsaZ8ztwUP7l/DXKC9g8K6unC+u1cp4Hjbo9PCURC5U6S
mW1hUufcHV+ZBJp4vj6jQj7EcA1ayQ5p4VqzhH+QjjlhyvQda/Uw49IJ0AQFl9fo
OwAn8T5zwF6SOyA/2z5/rvtjQfg+1WijXTQqmG3kWs8/mlRL8TYi86ZlLo5jgURC
gU/nVJXrGlnI+RjbtkjPz67/MXldBSC/3AkRyksa83kdVHgXaKBl/LF2BQ1hgQ8J
SrQfenAhzNAg1+HqYjjofIBw35EXgaSWrMPQ/aMY8TvXPHAu6HUekLMhRJwbmoU3
cK1fX1xKI69N1B6Af8cOwPXTbjgJ8sp+PD36qOy8omSfWyv8Ren1yfnV0NjsmhL6
vThVwDeev+7o0T94PntCvnH0Np0xNzS/PhqHoyfbZ8W5LX3+lN1LRk4hJhHgg4MT
1LUP4rm3skZrBDNC8cWEtEL2MGv2dRGZBOluRgOQWrAd3AEav+e6skDO1PPyeulw
+lkth6ik4ph0XutYaXSCtBud7fC0mioNzWP6juSEBURQdXo3Y+0LkbiN5xv+FZxo
WE2Ng9LZkHLqZVXqVFtYW3wj/WgHtwZSpYUnp3kXS2kT/dOGjf6kZwhKTcqKpFLn
RbBeFguFPnwCD0iwYx9Fz+oMAncj5xqqUG8JDPRSVOofZtgDEadb63h6VDJAOn7J
Iw/2ZO35wv1yQ5zJzXK/SHSqboBo7xwVpVgRn6BDvjvQRVz/CXUdH1okXDT074sy
MTjiiYcOFQ+bGuFsPOvXNBIvSP+82djmQDggSxB/91XN4ppejKhVBSXVk5k6gflK
e6+PE1Ctl7XBXFBcUyPCgMhLgCuF9HC4HTIo2PFWLLEbmFhureKb4ZzjnS7k2Fr5
1IyaR1eb0Nkd4hU8NgMli9NVFCexKMiulpapzuc+ZsjfK/bTQjDtorNt1n5uMbtr
L8ngq1DkXYzkYfLdhsQk9MkMHUZyVwTStyx4s3wnOm18Sdvbpsdv6sLuWFW+hDZY
xDuDAqyotSO6y9BfUo5ex/Iivq03UFWe+Q68kN6AXtkeDFfa0GHtO6fkvi/9S4lS
x+YKA9gp4WlO92FINynHBodNGLGxMAQcRDCHiUoApvL6k1RhtK8rHU33cbWsqsb5
8vR3u1v3n7NvXjS0G4k2c5YZma6kRoT3LdesHtIzszFMTcoyipEiGhrUZMfSE0GC
bK6UCXDhHf09ofIj8Jv7XNqq3pR5O3edl0tyx4p6XUA+81QuFANzrPb5MOWVZw3j
wIp4Cv8KQWCdDy3dNrAKY/Zqgc45zNihWZQdzBRSOrfOr7h3cQHJmYmMgt2NWI2F
ShUwhvtch2NzsNsC2syPVGIPiBqQU2BxPxOiuuyZbPLsElimn3hTnzU24bL2+7Ka
Ra2nwYwJUi8hHoFI/BCxInf4QAfENlC0KAVjCQSfEu2zsAxvbBNyPIO4/Xf62q55
KKtwDsZWYkZH1Bcc87HrgEmssTHYgFPtulyZXjiW060TLngCSjgAjdCvl7ieQint
ZOkF+dFmTCiLDDZ7TZwi0Sq9hQtLr2zL8it7r5oAEKq2Ck+zKTeb5DRC30ilZDtS
K7eFvrZkfeeDKuv+/HogCOc/fL6Yv5leqlB/JhOPDAFM/EhVYt1wbgO+0Q2E2//8
mD7t2CtLIvpxDMful85GKOKQvUayJGo/gXh4CLCPuSf2ssU/NHFDXUhtvHDzGTez
QrLSAxRYcoWF0ZtX1lLHIzpp1DVo7KNMhgHymzYNwyn8AgQqfQoV1LJrMDLkH+tV
CQh7T6RSWb3h+FrfM2aYT5z+TLdyCsxKvIqAAtHAMTqNF2zL8l6BgpzM2pHJWlHs
RbUhJeX//6t7nxs3xm9Pg2qXvOLmZBkt8ki9t7zw2Gy4TBurv1IWupU0+ZKbrwB8
sZajQGDzfmIntMkPNIP20w9/Mio8/ysX96SK9w4Blc5oOBbDOjaxlfjnog/OGG5o
m18ebjG+BaEx0xKCKqbhPYv8LFfBjqxLzpyoe/LLjvq3aBVs3+IJlS3C5TpiwNS0
ooWAJXObTKgetgosA+khcyBZQ+oRw9NqflqlGCWa3xKB5SQPnGMSZJPi/XMTud/S
qE/52Hhg3q0OLkY4OBNMRdVlf/DxDCoU3blHo69b/93KJnv+XuhM8hrr2SDyg8lm
PCFbMY328/mnnvKaCpKSGMd0sx3x6dCU+aGfk15G4jJZ2va/Nb5v62IeSq/LftN+
FEDRkeeCYjFkGExQWbZd0ox9dlvtqTvP7RSPyAs+0kPdXZIDGyLym0Qc9vpiBvpH
4oNJDsMoAO7ZRHLlQV0Ch8JW7z+cjsRQQMjAh1XWn+P1LgvBonyYhisCAp/fyCzd
U6ndOO1+KSdzfqPzMxUDNhiw+XxUEzX0TMTtBk+T0T6RB7cm9TpBth94mUPSv2GV
9gzuj1DxeYQY+KxXj3C5S8z+DZZlQq5qfdX+LfonPUWJwuhu3IIAv6Bz8C2Zs/98
TzHl0UjZJZqS7qqN9gSN0QGmP5JeKmuVWdItlZ00B5QScr3wev36JQElRSklnsB7
o722fPbPOzEcoxRMWHjAwJci/0wjLihH0LtvxRygcmt5l6yR754ycH8L31B5sg4U
ZD+LYzxYgDeE6GRAquN0fVVTXabeNoDPtE4DQ2Mfxb4/o6PMLmsEUXVg6JEtXV2h
DcSQq9h9BF3q2s0wpCB+fQ==
`pragma protect end_protected
