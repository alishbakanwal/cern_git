// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:02:16 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
HppGaZKhvjCTvDz7bCgLtWqWl3CeitkINE5woN+Jec3uzZ7YEM3QaFL1NUWURVlN
RdEkk9/gCZHzu6R/u+H1g4UTkzHUsHLawihemg4NUVWVVo43i0guY2k7hM31z0q/
0y8/S+0YpMo/k8zYaY4bdp5y7dga2QGcWanl6dpD3xU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 25888)
kFf9LyTn5StcWhcK+2RchNHbJxqkRqaK4O5Y77+qdtAbki/JK+la+HxxPfFseQ6v
kcNfKkno6dUXMlg98QzGlwVuEhs/G1Rq0LZdxTERH472yt9eucfN8zioSPg2BRfd
tuEptREmVgGG+N0q5U+tBU3wIW4zfwGIOezA20nx2awVAm5qg8R3ZowPigang6t6
7PZ9D+W/AH/HIJGgj26kvN2J/STWofeOJGHvjK7OgnqCv/At2Q90upTNwnvd8+Lx
ag/qOEZZ4IXqWC4wsMgAD1gqAsMSnmr556DYn7g+qDzmL2T1t4FjXktrXL2hRSRA
VJoYzwEOYPA0bTnmpbFueCVgZvRyo/QnQxgqcKB8v4BWQRBeD++M/1CKiTIHJGuF
XNhc/ar45I15rZzpwSCAiV/YVp9UXBAS/CYkyDb0d8q5LkP27/bDW4SccoB3hAnq
XZde3ZVkqNGbJDWD0KIANWvId1XW+5BjZQOwfF17spva68ARo9JukmX+LqcvaXlL
JuE/9YtwZNAt38NS4DS6VDfT3B71xmw0cppX6iy5aMVZk/1jVWB7Q4rrXUcw9Ssk
LmKTBUECuLMoBEz3Uwy5FZRWClnbHDHZv+hmdTMGF6Qi+Muki/aTcJItTf2F9Y6y
QLKeJ7GCYdSmzUzu4gR25vXk5rOcl3FQxum0oMaNEhNKnm3Fn0WCuZ4PlCDTp01X
UN2FWPsR2BuHkUgnPPIr9GjusJkH9PMdELmQ2IKf2FnBdRTb7gJ3QdivTvURo1NY
TuYcsr/hBsgPQDpabpONWXGgXQfcamFhBk5Knxnvrx/5iP7+ggIlXgPYQpQtNbBF
hO7cgDf+jrTLm3V3tQ1FYfS+OTYYCh0rLnGEi5cHQSRzzjCkrAudbklMZNgrUT83
RybAuCukB0gBOfne8KNSdMRzIqV25Sg0E7kij5DYG9ZdDHS+iLFuVTomSThKR+bZ
fHN45L6IwowjUF2tmbUhXtwCuP9p34Sp2/zapDmyntzXIBJX1N8H2z/KzG5G0SZ6
a15vFUUvSNCxg7YGngvY07vv+C3T4LYjbZQs8fn9D1+pES9dmrI3vmTGp9CXbP1k
JomKo7bxHdQlOHtCMmTfRxoNQ33+GSZwu7sGUGpPdLgYQgOmEL4+GEG4TUyquGRd
eaCeZWsCc8BQAJeMe3jSgisUH6G7L691aY7L0ANuyabXkmiSbYxRDSql66ndZ3hS
jkHTK8TvmbkE2Foq8Zhf6Pt+wq0WMC/o22fya6xfIRavWE5U5eRCzQ2/bHnqWEog
eEKK1ylBBkOnlRuEKgV53XPp8asT0yu0ONWjt2AoRtfPlfl+/sWU1LQt/pQVQxUF
LGxlcMRlq5sxbTr0J/7s4CBhmGoKwNbc8YwPZuOjaNjoF490hOXDSh0+Y4CMTGm3
zHkH50+fVONOiwWVdNFnutcYO2YQsRX9aXkCboOyfxA1qobPq/M7PXolK/BXjB2H
SLlqpgjQpQqLCd4X8hX3DDuOij1hCKp2zqi33c4P2UVAsfvtwbAFrkuU8KAMoFd2
Qlcm3zRwWeL/hZFb9fJ3fYPvSRYxPHxb2/kM0M7wnstYMr6yiVQDpjlf8L74E0+u
Nz/T0cKC90z2pbBVrdXK0SeUvGxYNIZcEMDv+UcYT7qsu+/dyFEGFjpW/by+byGe
1IVu0pWrF8bR68khB0FZk4twMnO1HMOwjHh2l/L5Bf7kzwv75oc2R/9oMJl9SSuX
78HNDZTiYzaJg5AcauFWk0rYTJjpUVN2GA5GnxRQB0E7d7i7szxrSB9B9K5nwwUj
5vCssBgZdVydnc3Vm0l98NXbx/sl2z4a9TnGJQfHEFNTnpBYLn4vymuWVIun7+yf
fzTc/OmyeV59VVE8IXJmVhW+26aBE/u/Dl+VBcKX+WCTDZMWHpe6NrLcqf3QiLj1
TbFcdklrm0BLocOt8hblsgvm4Fmkr35xSMYHwXngSlLpg9C4MpTa8+Zu1oVRqbNx
tL6Kc8STOhzQaMX+i0lRzseWi6XRz2NLyt1xmNFxMuXzC7rsaZumGQiCpEPwYMlj
TvajrGvoa3yJD9xYj/w0QnRE8q4Q4A3zZh4HcRmJ0f8ALE0t/+7fBqMlkeBoeK4k
dAPFILTVqG4rDQiT83j3s07aEXjakc9EMCR85ZNvIG0IDNYw8YaUICx4FnFM0K4M
nyBRPIcKLU9kzAqPtFeeIkDp6Ly15BGJx0v7aeZeRr3ok7s2qNNLj0AQNCYYEUAl
4azmlNRZDxxRzXY7WoX7aOewXWM7Kq7HWoJEpOCVNqWzYvM46FdRyFoVjPu/Srlt
YveHXXJ6C0zPRoKk6Uj914V+Oa9vQuDytQk7cjWsald+IK2sHmAOBrRfpWvlC9Vj
rxrtYkiGURhzTOcWQ4OkwYWYhmKjLJludrJbwDYXWSOl/782mlufRYGc0IUrwoXG
s8+YmwbvcrHJ/kzkYsPwf4cM1MTCqnpfma0FwIX6SZ/Z0zLaLSGmFMcI6uSAxv0X
JQl0Iq+CmPCqn3AIhjnNpbyW8uU0mjwRQDcqyem9enB/bAGqFjLlWjPM3jH34OVF
WZfEt97Ooe6nb1CEAwbiBZ4SULAf017yaBha/dT0v18ylphiGcxjnsLzVTmDnxw1
s30P1Re6S81GrZgBbKBtIPF1jNxtvshW5mueAcEUPlinX5azZn2CfArHYNj3jJnE
uKgw8zL1oLaMvrb8F3/Kn4En60kEGj0GhIuGIPOdZgu8NQTF/cac6dN8FnLn4C2d
r6EsmS8BzCh7j8vTs8kn8KZyvcnW3WTU/77bWtPiL6wI75jBFLLhkLKed1RRj7gd
rA9Y5lP89s2cLa4vb/ikJFcfr6HIuJlDxoNCq2IPYF17ZkADitTdp2i47JY1eAi4
82LsAQej4IgVcEV4qkboRBqbXGoR2mkRJTS4lmyMQXPuc1MxaOfjeIoUHrBWiEHw
6U8qGVaWLBDz71YBsBMyx2IWA0mfXEmCeVTG6BvbmsJStCuE6GLJdRr8yoo3iRGV
lTO67Ib3kJllT9Eo5K8Llpo98FMjq0Kd45FG30UEiq+v1OiP330gC3mL3dFinvXW
+LgeAjDet+1DU08EUNFUjAiJ6ekIRmLxLt305QGHxaY8YxM7pxW8O6yaIAA/51bg
Bxs0loDFzEBQ/v0fkkM+bD070xwHtGOghLm+0VXqjh37dBfmjIdfdLjbAAttycJQ
S2x5QXGxj7EZ1Bh8ZnlChVwEwhJ6lSsD694IwKByiqky/m/Zzp0mzHgwzPvvEsG3
aAzuhUaM0B4YYb3EigdE2W+BZwKhZUYlnFEjRZ+A7YT8b0YtShjAdWKvUSPTRO7u
718QcJC42nZkDd2Bw+8H26ZrqEddY+kSXnChQrg1081pn4o/7NcoH4/7B6RMCqSy
KkL2NSOzSGiLnRWLYoL6zrVfLGK4SwgC6KKgKTaLlD7SP4ctRSFRiGY+jqqcd9Cd
nzbJmz34xKv66YP9wKE3lydSoBmQm2br0bKBcu8cYURkdOOr5aGVFPJF0XvyaqW6
r8YFeoZCECsZiTmf2uoT1+z/3jZCKlXCGhnHrs2ePQF3dXkwIfP2ZDqqMTpNr0pX
t4/dUKhSiTdanBNeTjoYpOt+9VOr7SMmf0AH02UHEClIsD3N2II39oDn54abqRPx
8vtuFZk9PpaSz5mLi9h/9IqcMy20TwXlukiDcVmXzaxcojXdJ1ipUuRaG6si2FiD
nTpcg712g8EmftlTDqQrwtC3a7egky7Y2+zAgimCx+/d9z9Xyw5Uq7TUOsEl51Bt
v+lipmx8+XWDLMHaYgtMawkmSdN/xg/kvTlbTznsLi5f6JH4z330dLpvnReOYfXn
j6NIMFrLcR4Km4XvSiiBbepq9dyTk+mMsH66xI9mfgUQ822oeNrl0xT7UClJ55Yl
CIY5jdc5KYR2ST7O+jo+tACcBjoXCMYZoX7rif7/oAziObhLe1w6xsGJBvvmdzF0
joakNOsD+tp/tu6SDab1J5SNmrWFj/lUbjDp6oTrnMq9C9lvYQhqWD3FRapPVP14
LYoIanga/kYMFWHNb7TqWU96C7KPPjLlinyvC7u+oX8wShedmAqULv6WrI7MbCd6
mMKn++hmndFjIBC4oUQapV0+zdYu9AopnMwET1ubgxM96vH18F95vZCD+FTBPWzy
S3N4Qa1a23rsQ5JC1+m1PShMKY2vUyrQpgWZrmkfqRzJFX3wLwnfock6SrMIq+Hl
/YYyHHhmvaIOg5+7OT0ISBdyqIAyuH3IHRD1B+lIG/zT0iS/4n8nG9+9VivLhE80
suGDg/xJdeR8QTVc34MmlsntkrIEYs/6XwAS/jzEI7WAUk9w8ez/nVZpL7OzCIP3
LXp3WG9Mo/g0EwF412YyqlxoRTOrtRM25NGdFA5oKPP2Rx/goMZfIDkHbRgoRaZD
/awmW1XuDRHdELDqDWU5aSQWwN7vx4gFECfS/F3ojJSDYc4p62oomqmoaAk0W66X
i2CMXieabQs8LXQ8Ro3pQZ1X+nT3x+/3CASoZqftQFyugGXpO0Q5/6Ojq+Ychm4h
me38iksu+jluKNauqEMQ+3m7xKzS2yILeGmKs/m/R0MTg/9mzWCVX67QQFV8PxQO
gDz8CP3TdbkeLSWoBfFfkXiyDwccdcUFyT59jCL4hQ2r2nDKlznNKXFjJtE05nCR
sfO53jqYUyhis4bkO1iK/O9CmeX4pICjM9dkch9gqDeAHS+tiuh9REDBpJVtVpSf
PaOMJ37tv3g1a0uqG8gxsbb9KTl31yQYwWLFTUSZaCFtMnpHiXOSuvu6X32eZ1nv
7GTM2khc7kdkQBZBazCvI4QXPhf7ruDBEjPGzcJOjaMPY1jvQ3wMVBdEdnsNONVT
dz9mLA+1bxx26wWXChSOkHm9JTZeJGkMOc4NpfwuzwZ8BVrAtKweTUusUEWAjmmj
9kz1PrjMldum0/l3s74U7lxrfs/1RiGNsR5q7tDMJGiQQaUK66IvrG+qS30RHxqM
xAaP/6LC4354YUqnzwdngetRDbLn6H4Db/xIpOoenecHYl8wpmDuqTB/5j13PrFj
V+h0xFEN2gDkfXDWUChg/XkFsWUjT1NcrY8MM8rj4HZeBq6NIdSxEbnrm9mhbNua
Z6IGya6IPe5mdCBP2JLdtYnm7qDz2UUES30OVwElHQkBQxOM9Natz6+MB27lSGnP
M7eWJP+21VpRyDQ14dF3Ox5W0IHhrJMKZsLOXrcbHdqI/IfpguNGO3KKoS77TfHT
KaHIUIMOLQMSLFi/Dl4ElDZctBf0r21O2lS5ThfgzdLIstbPROiS1lmE9Bidbe/Q
1AS1mSNwaK6ywfJILFZL/ijkgrV8Rybxd9F0wHDQQlat8pko2w2bwsGH8JrOvWav
vzccaarBWoEvyhrfR0hJe2DISqUd5MaZl+/gsMaFHHWfL+qhxedCIdLYWcV+IfHp
JUwh/acPTgqbl1CyRwlkVR1nMIY5iUn6GleTZVA/yKinvj4Het/VSp1jYtIaas7K
HZtA1QFGBKAg++k2DZLUnWFVtrjGbK/15GCDoGjzuXVvQim5smvXBTVqYyYbLnbF
A96O6nwHX21kDSXUQTYYiIcpcR68CGHdgpVPCo6YorcUtnNxBDyoEhK3diPeCVwb
FB6TfAw2inSX9Lu90oqWh/ghJ45TfqgBincglr8l3gWPyZXRQdIgOgZd8IpKv5wW
kyaE09VJPPhkkxGY4/QTypsA6jj7JybdAeMm6uwV46fmfMEdXbQpjtqhEzyFUlna
fpR2hLYmC1sF1iPrtffqNcSagG4vag9za3U1WoWwHlsTvzjuryNgzGBehb5hks90
dpMeYKKuy3rS4VSJBroPHbyG5TYHQU8hRamNjzgjNofl//C3uQrGH7h5jGBs/fdy
wfbeL0PVzy8wE/CYHtKpWl6ZPT7FkovqpW5cEGKNxzUdhy4s2P7c2dcHf+Guadlx
n8eeRTFVP/wk+feqQX50i3S4yH7uJVb1NTfbZ4eciTzVDYhZwUinFKJLtXtD3wTi
oZP9M0BQlfatI5GkyneO6m3IYtUkHMLueGd9X1I7TAYRaQs5c+bnbzMcfhHhJdSc
HHxqvKeXvdmtqgSBuiqv3c6fdvnX19cxVVmInJvne3SB7k0PMK+D8YQpGwpoKkwl
idRI6EY44ytWv4Qf53QpZsBro5cGm3wgfNt1ozQ1XfR+L7u4G1ntB7LQ3EeK/7JP
m//o6m2FlgFJE7+oR0yxZgBJv2ZF1Zy3vWGEZo64tHRettLklv0pdn2GOMuS8g6Y
ilevw8HcxrpAtfdZvx4vdceaRJYKw+OthBUV6h8tBO4Jgn/+d4LWlJDZIOcCNwfB
JHdjDzuQGRk78Ywk08dkiqjO/7K8L2A/GDS5rsUj/KW0unTNGA9OzQLvHw8UyE11
eCBupgCzMiBcjb0mlqTT6Pd7ANuDLSYZLdy/yl8m7uqLLhw0shKAUQRS52fRU+3R
N557P1JGYTLmSQOToanCQHVxlU1NRLp5nq0XkI9K4L9Ra57r42oJrwH5DWGfxUbu
aitRROLaM8aUt7bOCYSHEo35DIR3KGXLFSa2v+K4AJILfqY16XKlK1ImnVGutrKC
c0Cp4/JYECQ4uj5HBXfqgr1qAT0dbant1p7XD4/5/HKFb8zyDbMoxL/6hKuXrs06
7oxeoL9KB6ui7ddfbbbJ4cyBtT4xNQsKrYKRAOK0CFthIN81DaYULM6IZUmGRMtP
D6kaIyn7/DBRAfoVB4Y9VXkH2dRnLUCXtF/pSasYDA6iqP64w49DCG6zRkCEdt8z
iHUbX3pVCt1j2JxmfgHXotBEMXwE3r8vBOuTuvGvICxyjMSpMkhNTnPsFp/rMUIa
hebUiWgIJNtk22Wowh93rf3u5EOt3SF9i3pkY54iMA3ISbhgF16xW0I0AYM0imr7
G6Fv4SGCG0r61BC78haUinGgNjkd131UZJ/JdqSpne0exxGjDOkxxGpfuvH17SA0
42azzt2fDqLg9q+aHlccFY1FnvEgW+4fsTJtp3hTcOsGLG1n3X9QfoECAPhQtD+3
A5IvNg/291sWZPoj5DT8K4JHPxSLV1skoYM1DUpOfRAn/8a4ceo4gMnxy232q2hX
ubN05Y/dTp1ZfJfGd+qGNElT/P8s+RK+44pJmFAnXxCinNavZBvIMt6i15XDIfzE
r+MZCV/Y4nyPu0NIQoW3zHX3Ti5m8h5bs2HIM88s0n5gIsbI4FGE4futysTzpQal
l47B6b/DqrOqMqQ/jdPAgZ4EyxqaTDZVsEmfLrJdl+L7yCfw5+G2oJzbQx5FMrRT
G0bajlFZjOIhgGD1fyu/l7WlqrkJEAEFMpdD27JqC1iPBr/4eHRPMymlPoO4X1Y8
b6lxPl68LKX1Tz8BHtREZsDV5Lxb7TkOjW7XEgeuie1rke3c75oD/bLQHCj7Yan6
VyySGV44irU/DRpvUXKjbTDgneo9J0FyyeuQhxLhnNqbXA3EFD5dir7HuT2UxQNi
GGkGDmaO3E2epiIf0DkRH5UoE9kQrlSpv/sRY1anHfUWDSlve9itpaxiXVZOxroh
3EzVYysdVaB3cpXQn66ZyrVS+G9+ZGkBRqElfy42Bw3SHPXBqt0YjTO2Y+SBb5ej
rNDiYq81s+4c8h0lfXIh5hA32tpZnEanUHzfmT4623Q79acg+tyii1v3FnuluaZx
9bhGtsyVT+8+txcKG7Z6FMPMB7zIgERY356V8Uelx0zHjooOKAujgTFn6kgA2Re4
QC4WbrGmSE6W0Ur+LGFfP4pSjdm7JM9C4DcgxsbfSp0Ye2OSRg3syIk5mZbCvZlL
D7w4YQOyMvCl3+24yWdqo85+QQbVGRA/yFUjGFrA4AmsXJoQhZ7cn3gKq7V2k1o9
7DEy9hKQU891EPiDAJ7qZ7MuPNblQoQT2lz5fhLeT5CqpLOIYZHhX+6RqrgirLEW
Z4XfMV0eIon5uTlcpi25InFjdbZStG0kKicKCIODbEcEBXscH7qalAEsth/O3GJP
1skLRg/QGhycFlmRB3cUfdasrFFSxWWS9VHkaAwle6XO/lLLaDO310moUNjM6xGq
hWb0jYdvWvn+m+O10mxU9w28ebtzuZ/mpwfLuBtNR0nSp1oUegosQv1mdWXi7Gbw
wCwLAPC+Ssa33LcTI4Jn3ips2s5vV2cSOc/6E0oHbAZ3w2UPKrau1nAQXHSO0J6F
7jfUDnd+L/WXIxraNeRomOhkMGKUCiZBU2Wy+JZCQ3gSggW6OYgaPUF6Rom+d2xE
wvsNQ8xtgF1AFFjkLsza92Xb8oTCS4PIXU2XJGqFaGcyiVHwyz/ovoe9riAwnpbO
1SPo1M5Jt1GLRFmOKdwkm3o762q8OzkVwq+1a3kz1OopAHlSIMVqW9yfkEKX0KcV
st3dj3cyiVa0XovlrhLts9Iq2hdlUOmq/0tkUXPVUelV1xubMNotcwlTUGXCIKfd
F9U34kL1ac/KtxI30SWmWX3doBdVcUIKKE48Cmk4n7IzsSwo8CfsUGE6ccKe9r0K
alxwXnz1uwIzWJkLyqVj7fkgrZmj9oUIWHpPSDeP8bX7ilCBmIdNLgx6XW9IBujx
m73Vk5++KYgfcNYrl/KWcBKcjIuPFjHlOtutqZC1M7mIIxpX51EjV2xx6b81b03i
Rv9KuZKSBWmRE/J+qBRnWHXjvUXLHYP4p8dxoQlQb3zk6fAiHBUPTHOYfND3hobS
nIhVOatSH+ah+pNiXKsgKtBXY/4WyPqDY0Fx94TJWsbReH7DMM1Jr2Mxnqhe1DFk
BxzMl5aQZVwSNa+FIgkgXIMdHH4KYUZWG/Nxqff1RjMkrqBlKWCBahApP8qyzGSF
GPnyrdwgQJ/5aW8IwqHH1URePrHQ2QRB5La7Y3qby7fTADTDrFpDduHI3IG8fBUJ
qvgdZSUyio/fmucL9H+c9NfRUJbSMWKwmJ1cE+9zp23VMhYOelm5D50lOEN7yrLO
Puhb71bZMox0eDOcpuf8CFlYwsO4Ge5kiIAmUKlnJ5AM7wSUV1ZXyh6cVBIV2xGH
url2GXc9PeGDBkwK+FB9XNVJUxq37wPcqON3wNC3qTwK/ayzclCV6JlAlGgQ9aZK
zKKDjaUws5B4bd7VmtfhbVhINy+VpTW+qvd0zCJx+bjBsXht+p0mfYrrcffpJ8II
NOjU5+AraVFG0RkxNKWmFZcLCDF4M8kj5qRku7hUsN9LcHLT56CnweJSXSArzREB
lPk8UvJamAtPojkz+juBvwBU9eXA7xSdNC+O/tkCfjvaPESA7HuTSA/COauqgxn9
AoVhNpviWikBrMOkde+XIEMn4MmGx6wY3rZ2q6e+sK++2Nl/O61BlNyNlnY94jCL
qho6dkcyhMLUjNQnHdDPwf/2+WZTJx+691ij/HJ9Zpw3PP8//qYbxhXFE0UTTfZ7
j97cMbR6bxbXsSLVNc/Gcyxk47Em9HBtAWDrww8bcBgqiV3xId1uPQ/MH4653mBj
6edHfOaeLwgQazDKvrL8lyndS0uZzOAxCAGCxMOpSkC4+9PwYOWNS3Ix6bA5PS3R
SXznjRAa6jCWIWOwtQytgtz4asXlD3qNLe5qmxBG16rd//t4jbm/NMUg/RLvm6oa
oEUs774lnqluOuq/Xpd76mzvRIoAjuoJFqDTRQZF+cunNqGzCDe0VYJR0WYZZP/+
TMv1mUPd3w0bB9mV2TusjVVTedj6fdp7/I1596SAQ5YujPWSm/Pnq1LYcfRE88oG
7qpId9Ub+jkiCQgNYm1/bwLeEn+1UvZX1ujfmCSlgSi8ziDCWEOGglaYPc1+00uE
y0WJyGaCBxMGWYcdovLFgjRTLACRSkV175SCqMcf+xkYrYzL3SyOQju5pC99Z7tx
cyKrT0aEU20QK+csanGJIugaQngaaqqQI/bgmfiZ/oFNGjh2A2/4ABOGMttRNoC9
9aONfsGzmGSkEtlheetlX3nde654we2It2Edhq55fGD9LG5ejk2jsMgI5QoEZ2YB
II0IDkF5gfywkPNlaluG7eguGcuvQR6W+wgaqFu/cWQ8+jwqindPfvwTIHOPqA6B
xn1iklLOA30+asrLHf6a3gjTr2u117J0ZV+4/MiOOj9Zcjrf1BBG/XyJrg8pgU6k
NB/CrOQyOwdIYeyjkRWrzVXodMl9mjmBP/00PyV+3iUxSacijWUthYoMAcRXmGjg
faFAcj0Ur4iMnCLxyju2FHbWkxQa2SaCaQJWEOYacYhrfaA6/HOT3+FSpdw4Eel5
SEhQEYLX9XAxV8VZwPgV84Li2DokAHaggrfXryONM/AhtGMzcbc9IYvJVj4jlaMq
arwUhcRSTil7Xl3giz+CwYWJx/KTEd1PUBeLMb22ldcu6BtTm5zdIIOfPrNfybf8
s3jlqd5B1SnUi68J8HkTG8jIjDlHkbmRWgfGagZbEC2dpu1VeOOkFSyOUB/6bK85
F1z43pA9t6f28N0mh5hO4BAW4Bw356Jd7GcHjwvuaHu/Sxr4nBAfMtR5DpSpFB05
xuvbfdbHwJuwOHehyMRMJ4OrFDYe89BBCZLLbo4+Of0/y9KFqKl1xVwwrqlfHT8t
cE0W7OtT32XEhiTcZrgV0P29apubaEV+JtBdvet4g9bEAyu12vaBwpG2OcWAvk8I
mA/PfIDZlfk2TQ42rGNgXnYZgjvZw7h4TM/H/ThewF/J2naHr74pkfNHzyngPWBU
mZmsLq9cbRyMrDp3jrdJkYaydp6wmep4M4ByxXATfuYWeeUpxIU06AWG826l7GEu
e/vOzhPGSNjjKsCPSVkICdzbDfSMpyosyIlSP1KqTDF2JUiAEkpfj4m1MAWJk6GR
ZPX9dqRqRvDeeZbPKcAL9kRwpaks522xOHDOlfWUGplJavROivLamYPHFxoWbss6
1OvBGvSwwgiTkHPDRynGjh63RcHOr9vEKHkC02AjNpKC4K2IjoAvvoj4oClV28up
k84HJ9/B29a85hQd9z25Yo5dfAlgiuSGvn9l3h+9KR8sJr0Gm1zjRvqFDWTXy7jA
yy6lfzrNOBwkFlV5bEELvz4p1wg+7IWCy0u3XVxCae5IAMsVsN/0iFFbeOlV5MON
mbsi6e+SNYsmVko2Y1+eA7yU2oSh9JeZaE+YT2i8u3z0ROWuhoZmEA8EAX7Y7rcb
wjEOTpKQh3SQmw06sI9+q67IhgOPXYCVKlsW+15x2ZUWzHWzkWL+YILpmwaCX2Ei
AvJOlNB90fS7lzqnaEzQjyZueZBKZLawgi2Qviy9t/lXI+ZUi5leTnpWYwqmB06W
Xi1p9fMAWDcV+4Dq0zg2RogCjQ00ZRewp6hXBs61wTBI2nQwIzHMW4iUhdhsINUp
TrI5yrW86hJjnNF+soPoO7t4DlZHPK1mT9+AA+kRVgAMsUI18+ZQCt2zcYAJ+1ub
szhMwHaew0nKunaTVQCO5bA5GUBvZbzbWf1XrUp+Ffqixu0dHtAhE3dbJALg0S8W
0fmqOX+h3bm+9iXax9KU2/sZevyfN+p/kl+kWk3ils9CNmGDlhbOf5WGm3ByNMlZ
gpQ0dtQ75VrV0fVYetOMYs8XKVmJb7SDrSL4l2fZyHlWsATnky9nF/1FVU88tkBB
NYw/ymUJh13UydvDFPKfOr9/KGS4sOFYIsRTUKatYTCnslmk/xLSQ6w8dTpQKzuP
w3hJ9znlg5rj7gFGaiXAvLgXMGqdnlBAkd39qrxkc2wht4bLlVO9L2JSw39EgHKW
DZ/pdRFBD9++Ak9qisJTx4Aj7auzZ0IlBxQFMQQI5zTk1NjPXq2D8ibX3eKmItkf
nSzLPZT82MZgY2rKwKESmkoIDGVkng7gGK0ZowIUyK36nDY6iVj7hb6ntjaW0wAQ
CUanQVN8f38NvTUAAVWqZkLBYGOYqqhigEIFj+0fJchPp/GwptAL5plcO9e+cYTc
tDJpnGp4sP76CLfbeHIDlZ9S9jV5N8HBkOk/Rt2x8+zUvB1WqG+HeUFKyc65jzEI
3zJT3PQJEEsJ3y43XVbWfG0Ztn2Rbev/r+uHW/ooKvs38D5dBdcpQJ9MWEN2DwFI
gIxEkOKOVN+0CzZv4JaLVh12qmPP4CXO7be7+Ljt/AErE/6Ay6SEz3wDSbhi578p
y74Y6/EBRRpj+8qx+xR+/DJNlS5R9C+kw83pZmIMdYqvQccEs+guZjf0ctWzGofV
1UUAS7S5TUguZjxb/HVrRCWGG0KJ1haBP2tliwZJbZMVhu5yAJyksErM523IYYW+
gcwBYlyoMoU1MCnatFlvszisVO5rIJ/QTWrO61mfs0iENDb+K/PigdY0Y0m4oK8V
Xm0DsZSXAT/JjRI8gGiBKkBV4P3avP2fP5/GCwbWlkzkgodQmYwqPrxIy8YedfDs
K5fWcJC04177vJkVBuOB6iuBmiOc51wQyuBQZ+Y2qkbozrpBlYEluI47W0Vkx3Gi
gw6/YcPoq5iqduEnFJB5E4nJ6F6yPkSTKvzn7uMIEdsdnOiCabmYQZUnCDmPM4tR
d5U33FCNRKYQ3MI6VQgyuqTxedempbDPMnLYF/IUCHOzpQBHzwN8+tFo9G+GhT8V
eAJDB2szEMBaB2/S1+WJQJ93NIwJol47wK7egc0F3xkCzT7rFThUzVawn+v9r3P/
goxbaTxaTUFiUZwIEIFwkJNpTg9e/q+g2ftMJWRCPq+rUlftFVyNDnHNNlwOSm1Y
9I56Wlxk1sPRMb0/Wk9y84iv2CTEAnzlcVc93tsM3Sm0nwIvfUgQWMCeOCbdM11a
8Axmv+cS2j5aDaB1V1c4k68YUReORuJn4mnp98ZsjRWNP7/XHph2PP6nTs58edGK
uN5j4PuyKj4xgpjGwR/DxxjJtlvHIZggGGg8iC5vYlDUbe7IGqKzeNsRsUqvtRuG
kvtnukRj5eUmPY1JzhFpT9a0jImuClrh+Q9guTrTfbQxoUbJ/2lQuGmkMc4OkLw7
ft3SnNmNgYY0s/KmVMPrPQCd0Hl0+Tn2dLrGjmgY/Pecis7wQC7HGaYd16dzUXdy
sQJZgWEyDR213TYDKzfoVIPK+zzlUdVg7X+/7/DGhAPeKCsXkzwAZk2Qfd0q4aBH
7KffmSbhDaRaN+n8UCcmAUs+9QGbjKmXXq7tuY+D/0bZnl0WyE212HIDdihAvLKt
nL+3HTHV9yYWO63dh5ghek2+4mhbx4AHWI9DyIDRhCSkWAvIYOh5PILrirEVhk36
VqXYYbpqDYc6SbBpS9DyuxeoZliKypl6K20P7Ba2oT4t79IwMiT4Qe2MqBtsGFD0
LdtNJRZm6gyO0aTxAnDfS1ujlEyg+XhDAbOtpNq2DBLH8SagSzezADf/YbRWb811
qqfngap1DTf7Ft7PYJu7GH7oYeJt1zHNHZ/cd3nqK+rq0wSoqGUhNMR/47tH6TP5
7aCKTIgAwCNLqkOF47FpycTFyikuHb2ZejYn7Rw0U+OjxTYo8+eQyGCM8quuNtFL
Vd7FozOnmol+KfTpUkc04oSFICnc7msJa3fLwBr39hUCDv/h/IjC7/NK0SC3RFoa
vc6FP+w96yYjpJF7eJS/GW3Xc3Azxak1qv+lJOdZApTRvzte4WZeP9aJMXQjVDSz
UzfUtwdrHaonvt/RbDsNFbbtOcMR8XZ3ejLKBVToshqImK03TDmziYQ2NQtW4BPN
tkzguTghmn5PzENtE7Rs0LEbpdxXkIe3JHhWcB3kGPZGoEwQg/bN//Zkmoly76vH
dMPBWnnRttICxvddJxxaI//9fBpXetp/Ag/doBp4huVGxszhbK+7b7hjHOVT53hZ
nfraYT7+yMPP6JMFL77Q9voIJxTOO+68s22cn8+AKWuOzxL1evsDjNaFxO+eba7M
UfDGc2crae94TfWEB/TlJqR8Qbjnn1F3fdG9YJnE7NWkDiCax8FqRYFAe6BpzG8m
OyZY5jKBJ76XjAmWB7C2lzVJPraMFOykqGEp0urCPqpfq803PB45mLYiKRYUt5Kn
eZdELSjXluzG71rbq6+NKwefuMXGBss9gOohQ1US6RAHHCjT4LukehWcG++DYlFs
67ruMmXSf2ABaVuv/Ccj+BhiHU5zpp7mUPFNyf2I/A+qDv/Nu7m/QdpTrE/LQ2PI
D4UX5CDYdte8dbKbvg7f4NUdn8ljx6MAI5FKe3ip87adHADgNHtbkLuGs4AB7MVD
aP3+MGJK3/iB1wP/OJmGUFRn3j1QjffpA+dIlBxiqFww5kTYj+Yyr7U1g7OMtoMI
oso8AZJTGZ66emKlj/2fMICPUgJoE8iM7ze3SCgeq95r9npgVqN9wsxuFAz4Bslc
B1Bw0haXGMpkl3KTf7feBlhEYS8ZJ4mrbH3KmMNMaromRCtEMqIvuP9UQ0KkH4iE
JPoyBYf4PuWW+baST3vXCIEP9fnjJe020SU0Y758v650pqZy0t7Id2xZknaeMrbY
Gyer4qMiSLmVfZK4bhiuD2VRzsUiPNdlfD1an1zhnDJ37b/krJCjQghxv6Gcrh+N
s8tANAy/Lm4pgcKh37wdqkJszG0NiA3AQHeOI0nI0GNcOYkzVpPLJ0YXbKows+hI
4JONh43E/SHeIiWNsF/I8Y7HIQsE5DJQi4FvJgAT+JTQOwjb6/Ki6Lq8XJ4TSz54
AoF6oT3QrdwkpyheAVpEqUuGI6Vfsvsloe3QuWbExg2iV1L9e5v5caw0JjbKdZbl
/ArXlps8YIRTNwvCtPE5gXaYcX1HAy7eQIRpHmhC3ZNTMiMKUJu0RIVN1fy9Xapk
Vlh44acpWiUjCRhy72I+Ai7vfIfdH+FZwv1E+dXx2KLA5+o8qZeuyIpD59f0Ejjg
vw4/ZarAOYV6K7FEJZeEb3ptfgPw1sgh8WwiEjEums+7jvICSI7XZbuNEq/SzgjY
Rw2GSim65ncgcD5xj4nfzIko0C0+VgugI3Mn1ojTETAOHj+QNib4PYzGxWo5WrFs
DQhZZHqAwwWUHJkGy5Vkzh/f/wO/6w+KFhPU5JI/z/E+F/qTUZp0mBFiOoGPpLpP
i1VR7AKf9LjWFcMLrSpFIt0S4fAutsofGC3/+PUljX2fOQBy+ierHh3JPEDVtif5
j8tid2FwxuDtOgUtmbqSOHaO/5zGbp+N8FPQEZfqRuWLWJ5SR9fXWzW62PP6YLb7
7d/OT4iRgXseSq5PawwKVLalHzSKNXfRykmRwk1H95nC0Ks4IlFCAVPEEpHnHEqG
PSe7Zv+MtmaeOOLT+lZqTv57pEP5yzo/tuK802OIV+W+WgNNdWLXGmD/L7A4Uz2p
7prJlgzP0TsY6KpsFRBYz7JY9Ps/1d/GrHW87btSKpRQR+LviGnvk3jJOnoSDWnu
DbqnjlUIgNby85okBdKnLYJMuvD59bo0DJ6ExSn1vDAobDPkGVkHj36UZgzfXqLq
r8okgxSrQUxQuDhDBEiAzxyfaxlaIAITckKP3ncFZ2voiMPHjE0YmDhDk52epJQd
0Npw8bgkw/SJj9KeJT3KOjsyLI0G+c7p/ENra4eLUmrfUi23UYROpRFr+DMPjqPK
YzML2RrbOdBOykFgg+RZ+VFv9aaRysi4CCRncTwldnRx4gIyXEMZlIpNw7KIUOpX
wcWayCMCtwDfVtK0t/azs4I9iKtW05RTF5Th6DMkWGC5fHJgfx7bqP+DQff51okH
noA0teeJFI289wklbKHu38ASBYajGUl9n6TbQGcJaHkNZRpX3nJ9bYtYxIKCdDkh
yc8e0YSk8MvGg3QvxWP58oUUT8GDDvSPhdDinLvx9/pOHK40wG05SvPBu4oYm5UP
h1pbPupzReObbDNbY6+iG2/MMo4MT99U439arGA+OULYwmbCiY3CSpKJWlE30hcz
Zx/gMn1oTIpxa9oYHeIUkhAxLKxUWG7GmIN7oUu3/4PbDKb3bJpuFVaIre4A5DVE
fuLyILpv2z3/po4W8HDTYBLm0qwAfIXgg78ZU5IYCSYMM4ocRwZbzHwyyMs/pHZB
X+heq6W5+wfgxiqChGx+t7MwI0OboEuG+pj2QWWkr4iKc9ONXfDCS85Le9R9Rlh/
1rFQSax6LisrdNuUpUFetuKP4al5PlX5Bjs8ihGAa7wdWWp5t0Uot8llaFmfA9aq
drHhR4gMviwDTZ5PEAveqxW7D+iJnbyMquj726uDKORYJNmn9oaD1Y7vRDp2H3Ej
ZornivcB1U5u0JMROnFcJzJqkf1StIV98VuVIVLhPiICIwzJDuFcbCoQGSwRNgnD
adJRpG2oUkOGyMsgGrBrs101s1y1vvV/JUe1R7zJhXiHjEZTeeroHhVoCiPcIA1N
c6jY6M2C/B0O3AtbQltShoxa97y5lrRD2qNc+YdXavupgRjzKGPtNaPuGvZ/vlsZ
r9LPe+cdXgVEViZ4DIG+rMx3Hua0fEUTUXKJf3lKna12uMI/HYYjCjiXkkSFVhTQ
EUWgsdoLuLTI1bsS08B08dSip/Tko70CqcyaW6E9vC6Boi6x8DGnCLQuB31tOt1N
J/WTd2ky2xZrrMAdjTCDsnEka8YKw+nHZU634MxszAoxj3m1+P9D8jDDpasVwIWa
3wr21XDElybo3x12rGbXSw68KAGZbWXYY9kecInv27w/ehukrUT6oojf2j35Q+on
PSPNaMY+XeYGtipjaPU1jXpBAckltaX/iIkuMef8qwFBLbCe9qtm7G5sUviF9/Tp
DtNdu5OIaBWZXQuqWe54vf+a4fxBEuVqGVA5GXJYiDnbRYE4Vhfnq6eqHWYg4huN
6aZAq/UVCfNn0uF+e6Cr4UP9fx7iPzep4Rf3N5FXnSGIcSU69o3xHz2SrEbTV//w
bUbCxPZ1F9P2O6Oi/JjAaWvuJv9tMH5RXNYRD919S/Xwu1P03eOo7MgIb86BxBfr
+qzo59zq46chhT3wpPrsq74vHC138oG7pUxf5Xo9WuDVTCvTzu8iSlsPxeFu5D5A
nY/dVghnX6mmH/yseiaG7AICPbcS6Oh8LX/iToMwFaxtiPkaZ8AZMo67uJlGpcLP
rdlqXSYjNOpOtqC9WLYyD/9Rq/HS/Nrs1IAODsN7xju3msnZHN7Z/MGMFuPv+BnS
NVd1z2NIMoMsTy/ZXWP5mjKXnIE+Z5eCwen3NkYRT6rhazWx/SLfOw2/fsNGgYZO
wihcUDYukfYKIfs/9eThiyvTRneJZIrg0SPLaYwRIpu2bO/n/zKbOmanzxZy5KL+
TBGL8/n9O4wZbdkLeovYVUHrdiZy+m0L/DzTxoYKtNKDEABy3o40H+/0y0GrvH/Q
+C3AwvAwOweFTkT00sfFPaF8Z3iy4bvcKW9COZ1aDPlgxFKvYZFSZcIQafc7RuDk
rmjtPz+MkMSy/LVBAlXkqR3nFskMUPHvGSAnpZGnddvLs0gOBg81yGQLOaKLlavV
JA6Rw7FP2dnzI172kcnkHRQoy85jCj6AIlkNI5bDlkFkyHG1ce/jNFtJf7zXauxh
GQp+tIe+UmSxGvukoqx2XvlFnhpcB3u6XELvyf1P76PMFuBn7aav76BRUAPvRlmv
GfjkpJcewszdqSAiUF0/ADQujEwGvc5AYWiLaGWUY7Aa5QYViRC0XzAU308vDq8H
9909/g01I5Rl7xuyMNBNin/PuhauVGbAGYaDbh5Ztf4h5cgRXM1mtdC2oPes7jkr
46RaE1EF2ZfLHu98FEhHony7ZuK9SAFDiNDNu4Mn3Ndi7UMOCIS+EBTzOSCN6lVC
/84ij5eOHS5QQwS0lk1Q0jzReQBA5w6zwwEQAEyqpESD/5kTpipn7mxIJYaTH4XJ
Q82Yo4GyNSOKM5cuazuTjlqOwi+RPks07mOAzGVlZaI139cmckw4eX1qAq6TOaAi
mISjJNUYw9ovUqVJV8wsSky/L060gfhqzHb6rhfywa4hia87pEDjlL7R/Bdm0xUr
gPLpyqiGQcT4upyTU3z+1BDuMEgSF8D8jaVHm7aBUtLbNCa8MEWFsrHRi57vZ7dN
QS9mlZ8VynnpD5bGtOyojW7qBXfIwy8wwrN9tsmmB1GBtR+pXM3skUUmrUE+L0Kn
IJuhCVCIIUK8hD9WgTo41BtQZ/jvdAD7dEKHdEKlYEifjmuWaLzz2qX0cHzL4+qX
d/9kylM2jIOnAEpq2Ogu2nYy1AWh7gooQ20biHjoEl3P9LdUJxKIW6VvFfNpO9PQ
clD54r4GZoBwjUWk0Ot8gG7YZYXvUHelIQVL7bWOnesiqfm6ZtzT0upXf16rqb4b
L1Z0NO7lwQbwLDd9agML2SL1IHrS8vR0DxQip0aR5d2G8A+J/VuT3cBqbGQADsqU
TigN25It5Z9RmKwpRhAa6zEQty3MU3RiGEEujlg3wb0csZpcj8b/FngJNRjJO3bM
PuWZfWgDLKoFEPqeepgXrd3dMxkOXd4F4DBxCH6stRUrOlxdjVFWu5VvtEqNL4JF
/hRZ6X0RddiBWpSMkDJXOXaYpb+pUov9JTDDJgT397Ubo0pkB/STuAgDcXXAi26A
ytv3aAJdP3LTkLVAb9PkHdXOcfl0YaPrjA02MTGoBvM4rOs01owhwcyyfRfHdR/C
n2E3BZZvh2e9G0ShHuRbjUffw3A4dtAtYpAbSKra2TBhvMaURDpFwUbPuruOrMgH
zqrun7FUTL+ldwWX9kHnw/lmpV1VaoJPNp6zX+xP11Q93z3JTRTuZuJiYjeKHIQQ
KLaSrTkdWaUGVmy5cVW8QKA2eLx07qNj8W2mlb2hix1Hse2EPEsT4lz04Jqx870k
oy1En13MIdkO7o0D6j/iJCwZjztOPvPYgWmVzYzoTGKHdeww3hBQyg7TMcgCTKHb
UOfPz07CD4cDEDg1eGSyRQk6/ick+Qv3tW4QmMN0VP7nz71ZZiDvu6ARvcTch5Nl
K0yj2wj6Gv6exzPN158f6XuMidScY3Io+DJsHpvccGGHUCwPIGh/O4DqpXFQ1Ze5
Vxrz9Q8oQWGDaMc+dGSkIOJ4FFMDez8XcjsE00nScNwinhViGST8mHP2eS0uVv5R
kHtSieQo3Qy8zQ6zXRT+Pkbl/dt9IZ6mjpou8aMW+Z2KnsDfsd6X3DLZ40/bErEY
+tBRH4Nt/rfP7tntrPlnwIiLB7f0oWi43katpIJ1iwwZYUvnLualurW+J+7PSbOj
aL1MBs1oDk4H+8rcdgJEYKpZLOxG20O9ly1WbxdSozno/N3TNC8wGFa6A3B7No2Y
QlNgagHQ3WoUjSdv72m77/vr5VPTNQ0+pc5ZAmkN8/vmpBJvg3H4hQWsofy0e9hh
veuNr1sNqgptZXEpdoCPe64gLTVFMqMNWdxPjf1A2aY3rimcUPy4qfJqftf7jVxt
nNXjN0j5GGMhOzvaGtwXcNCFnptoHn20FpS+jteguNjIoeWIEzub30zarexYVLD0
103a1iEVaM8FTpgbJwP5A+lF9Y0jlpVKotePJXxYY6OLT/MkhkNQvrL3/6ev4bsh
URy4qWp7o17OJCgjCuFcm4flJrY5Ur/za3hA1d5a/PNyBFvws4ejjlvke7+NnY/O
OmgikUeIDu8Tfj1Z5jv4FQHPYpGPRJXPVgZyhYiJGekl89GvcUbxy2AsbrOxattV
hHX29ZDTSfbGVKdY4IyW3FifGfmSzzsjUBTO3pT3QN6BodUw+lnTIzqYDHolBK/d
4/IABHpnWBydMmZ26bKm1/5no7e4sPbbpCz/3BVY5f+xz5fVzoPKFGAqP22FOp15
ECCZLzhHqQjh3d+s5COi/Ctjsw5tbJtIoRWqoq8KwvkvG3worEbziVtm4jHGBmzF
Daa4SwuU81voGt+YZnFYfeAkbWIPyYhLwaQ2ES4KgqKMQfn5MVPSKdfXRB4ZmEej
KMRKK7V19X2ZrBxead1bPTkJ57otlc+JwIDpRjhz3e3h25QhDHvC8eVO/OihIWaP
Qraq0COkN0VpuD1P+aURnkIjtegEyieYli6lrbh79kt8Sr5vajL6qslhwwRnlxiJ
2LjJWHwgyWBSgmWfInfv6EfRaWE9O3eKV6UbbMj9ytNfNimYRByjwtmHliF9cZs2
e/CZzUY/VFF3Df+SpjAFErtwNPUlnswxOs+MLM0yY2ij9JatqIiyxiGTNoZhlkN3
QftkZ7v01+2B1VCICbC5V+uCywmm63JlbNO+rwVVT7TWEU5fLuN7KmKXzjdrEVbh
fZ7k8sC4LYsoWNMmOX+Gl9M1HFl/gVb3QQjh89YC1rmFrcX/+yiWq8vlJ9GwcRAP
KwtMKjXLLB8CPKnByH41LYZghOATtM0VQCpFcA2r/yaU77as9wxeTa9+tjk8/lmt
tU9voyL9/llyS7N93nc0nHqNQ6jngGBS8eCeEYvGdk2lnznMSvR2doxzVmim/cSj
Hjv/5CmxAVlxBQVGby01ONExPij3BPMbjKCGta1/fegBjFlSBz4/8fi2qDRaX8+m
T6oyVHbARveSQVAMf09FKBliQiqXVtIfqjV/l8ENn9cpVtu3+/Nmp9Q5wSvB//tV
NjtnRM8/MFr7OloB7Jk2/6lIxyiJ0+6qPMh8fDR4wfSLmq0EKJqYGXUxZw3kopSe
bmfBvKQEFOaj6DMrspYW/Zyf8FLdqCgbf76ipeNnL4HIojnK5e9udjvANW5oC9hn
rujlLnIpNfgSqf37ElOX7B+Hoc7j/MlNa8Ndx2BYH1i9h2u97/BDZKwSmmkNRtac
egpWRIo5WKc7i7mf+C5xJ1z1IUWHvZqJZvNV7sGENu8TvgpB1hS0oRTisKSDINvK
zKurc3Jf779S7oYFB0LZCw30/GjaGwF8bKLtZ9FCzromvyLK+CyHTIF6BGpgrRKr
PiE/rhCEHYFIImB7f+Dk9jym3jyMxubQ8n3xGmNAH1id7vWPKdAIdmTVa4YIuobA
skBGtQkFtMUSUB+bSOYw5es3f6CyQ3shHPM/ty0FWvDLaIDQ4zb9D8oR1p0SEpnN
HJorgRCSs3uwILerH0xVl+R2QA1/XgJv1NPc4tNv/ZqAZEgifja4mVPsL4ZplAbH
OilpVnJoE6a/TRd0D/O7lfNWKHssu06iljzTn2zzbaJEpGMfjtChPITZUGE6+GY2
0gtKNgRXWhTbGpgMge1nzavpTpRyzHfCKY5PUCZQGFgVyWAJr1CCqsRSIvwBLXFM
LuYd4eVRC5rBYr6UNViMA5/ER9mw1hHgO2VV7nF/zoUmRT0JVCfPSAugZWhRLnuL
4L7hWhuPbzp9IKb7YrnXwCB2ttLr/wQEH1LNwwcEG6ZQb/fzh3YPdbgO2FTHffRp
Z6nXbSUtfF7bCrfaH651oOqRxTf01bRE+4/TE9RJOGwDa3+AzaL+rq8qGaEOcSdV
Il8+qkH+iohFQNqaAYV2/x3GgViVh1hYPqSjXr8xWF/l5hfwWC8wEn6JAa1crMxN
kauJVIj/qO3LjQvf4QaUqD3OL2PlxpnER9m2oqiLi6oOGT31KUsIcehP7yooJ1VL
LHtBJBUYvXFbWiwireb7BcWYmSvqwlFGYCTtkYSvw8w/wEel8lSeoBtBjdHHixaF
L8lQXdwAGdZ2ZFJZwlygghNFDFL8/lJ1UUn1YGhgsT2ICN28USvhjA6TQSiDAI/N
my59KjGYsLzgigSO3PT2jT4Im7nBkeKwx+ig6QoGEvaTN9lVfzQiIh6D449CPK3J
Ik/JPq70Qqi3icim4qjGWDEvusGIcwPpCPtJDQr+N9kzlzKZcTc5gKiG7S18DxYG
syx0PIvQTWvLlxWUCG2EmqVWIz3VWVP1blcOOVJ7zVcmVTnI2SRyLTQ9RmPRX064
atH0b8X2ESa4byQzSFh3zRSH2Z7mireVnl+3NQya+1rN2v8L+bZsWwfg2rWyjLSM
TU6GiTyeV9mS/UQ9uGs43SROLPTs2qRZHciILi2JNRwd9uUbrHGPn2tTd0b68IuZ
rxCIgAM9Ph0LkdmoPSnNprNiXOacYT/xP5y49EZSdM3SNoEFYNV8KGoEa9hhDbGO
IuKQrEGAG3jHLSepla0DuZOe//WLij6jwuV43wIoOH3EeX5yUuuXArqbKq3v+405
GUiYT1DD9iSvEmS6JIYfCz7Bx9stVV3T7iMUWkTQrKm6yDfzXFEYKETm+47/rkFq
aOVUGVS77h2Uod+V4iqC0EHZJtJSSXrhpD5Ud+IUiTUO+S/4D6TMvlus2r6Nau6u
M0O5/dUJ6+9NEHTehqmMqv+8iRNRntdqnOrbC/sEhqylWmpVYArMq0TzsADaoayA
tBnRtVi3FoWcSFTZIR0FKIyavIFAuO5/3iEHS3q4J6CoapCEnyGZoIo5ezknhlhB
3h/ImmEtcAxjolxkSDGaCJhTTOOq8t1PsfzkaWw3zdGOLgAU6NPTKXqfkqO2cHHM
RISy586k2OhK1bkGf6FvcSvKQnDKy/8TBZdKt+OUTkmj45g7Ys/esLtOtduukI0v
jjzSyCF4eU9bvas9SnkVZxqaruTqlUT1YXfJv/a0oH7jlLqm/ZBNgB5NcWpZxEpd
XZ8OVEc+zobXnuLKOcLNiyohGHkiTUv951RY94dDnmbLiG258o6R/U5odywFhwNR
USCB7fVUfcQGi9h3O3uY4X7cNDsRYVAhUEY7kJsahDZy+JSu/4oBqbBgVW0Nlczi
NXiEwXIRUfIi29sl24urydq/qGGirEmlYgte0ZGNG/3gmCqMWCkMc3SsLCrawSxA
hOmGeXc5fGvVfs6JJtb38LYCJajL+f61pVfBZacrz2m4wFYb/cVJFFPr5EQiMFxH
DGmvZCicOi4stF7RIUflEsAE2k6gSsFdv9O7zLV15wmmNioVWj7aO52vJsoq22pa
5ooXrxFG+erNPTeJqw7Fbhqy6Fnz7rlmiFFU9g00d6H+FoXTmzRLveFDZ5xQjy6R
E/E04IcwaG7tLRoGNFHuQa2fqVhWXLIjvtOyak4jMHh6ZUqlnOwNcN67aMtymBDX
/XY9BOLrxe8a9TdK7xYOIiSmt9twZW6/KjdUpFSGW1Ggj35wWjsvauh3WA+22hVq
D1BtQjj0oEzSZuXNWHTNMwhtVY0gSOnEpBTJCqkGXwUWKQDqhaP2w6FTBphi80Tz
iTRxfwQDPL7Gq2Qm1NHpt0S41ZMs9CVkYCbJEvgoM3GwB9IDIUDBq4CmMwPgZRsA
EjnjI/RI4LMa8J60f5ma+1gG4Vc0DvsoRKXnqBQsT5vhFOgo/ErWKVR+t+1piFQa
irGmVZ3GYmallewRosRIuHiy9rguj3YanipP2ZO4zljqSI69wXAxkWUSx+nBP5ie
DNb8m3TVhxETRMwI6aqw0c6LJLZY6AwDFkXmAoLMw5ejyh8hZhX64jB+pZudbO0s
YD4N0av4b1VDd+U7q/dOYR+usdDQOT2Zf6J0osPxE4u7fq7Ne8t1ovQq72pQl4Mn
viHlfrRJ2zDDGxChKnq763T/bGrfXBYPpqIE9cj+eCMdrG9lG4SMA/i3c8jrOysD
mSdjjo9XbKvZpH64thubrL8lijHgzpRmgIZeIScEtPewdT6+XQT8u9C36+KCR7PX
FVFwHk8rq0D4vLBhBv+SA8joVpokLzREGtffIzj7orPj0ltNXc6/qrnml7yPZok0
dSKx/LxRkGDo2WHrSK3bJ8xMX+UQy7Grb68t4v8VhP6ia3UJ3xR8BPoPepXi0bAg
emi+l/hcGRLXKMoHCKKOXIXEQm2ZVyv3JdIuBmOCqGbC8aAoQiS/LJ9YBDVtWw1V
5C2r5P4vcYALvjWc/fYNz42pOvGBRaF5YO5ucKyt7GA6QJlN/c2si1NrK+9w6Ioa
eJIi6F3v0jWqRIns/J7taFyMFqSVz0YrOJzjhfcVtqF0QbQLqbFmB856Kpj5Hr0G
1oGWa5kLBpqcLUNlz2uuKcVAy/vZIgdrGO1erRm22xlYskZt/rlWKdJWGtIr9gIa
k9iW6YxFt0Ghsw3XYofRtY1MW2YpwT9NoGXYGpw1kyczP8MCkwDw89QseW8ECXn9
RedMIKTHLPoA3EJRejO0+UIiVaeeq2Lof2K0BsKSLdor4gv9WFLQCBE056Z4vDRc
k33Z3K4pdFDEz00rhni+v0uOVJs0PpWycCHmMFdORHOASW9ExlcLg1D7SSL0XLC/
9Lv/3SxSG6w+sF0jEK7H/k0SV7oU1Ng6rzRv/JH9x42H9Bwo+bXQyLNvWPWM/IZT
wyXeEVsqA/4fxB2gsyXknp4XbBeB4sqsRea7GdIzTqZshqOJiYki7bHlgvb7yf6O
1KBK1wmE4Hhtq1xNFUlgV5SU54ZWGdEdOmDH+WLz4zsNOxiEQ0W0Wa014Tz2f2hN
rXqR0zNNHsM+9j1tfW0UGMepQz+hDBUcxsBPakhilj3czFLmhE+NVsqCuSCwJGMh
JMTHIrdyHQli1JnTfVsey316tdj/YtW6gJuETRc7J1g/OBNOY2tSx5CNGj0u0NQt
nlXWtGdiKTtq9v1zzYvDx6sjR8I6Bogv2PYPhbR2etb+MlxHaGUgT1wSAO4Go/p/
YcQWH03lwNBAO2rtYzVZBNWlUbh5x4yejB0+NfpGvcKC4e9SLRzuO3DjbbT/0Duq
lYqm/mwJUZ3r3QT5QsRtud8tOkCY/E4DWNzeLTKcklMTdw+mZ4vNMFP0dqsWWQYG
JCqMN35ZHuaH8rhHayUbsbPBOLHup6jIGabD+9F0ooeZ6ab+ocyNTyOs3oVZ25VE
yr+vo4/lkhgeb6zTIfUt182yNnMTL07m5Yp9SfAk/cLeyIbXrVMNwnMvJVkTyeTE
DF9sLStG2cPkgsFqEmcrcWklcNaDq6znoqJoijIfXuW+mdg88VSviFn2Rkhw3LyG
BmsufjkbBGPW4BMeX3ozeoiIJCwBK+ZcP/sT8h170grUz63T4St+HQUJoHLbXtFN
MKKqkqRc7pOWMR8EGvHL4PmHx5+0dAV1KxYG/xb+mh6fB3xD/ojiPzYgrtHxLSQo
Bcr7T02H+8xLQzbp7JCo2OpkhBieg8DPkYAj+ZOI7ZNZybWoOKdKwyukchUzXSFJ
31BTeR9CoQdc8lgvMlWdYBpYXiNTZgJUaqOdCQz9H0rKUfqwbgv2zeBAO/yDtrNZ
8xdNStkBM5/g+LxV9HF/3tyMyh74Haqr8gLKHkI72zDmD2vHa1DhobdoAkP9LPYT
8YtrGt6Q079I9W5FRu5MbvwPDRIngg0FaP4C2/SithZst5ilUSSiEaiIfHIgocC/
liBqtF+DB8Hdpf8xnSAs2NzcHlmPSA/EDu0/Op2o0/AsRRA5hxvJ/Fp0hMllmu0s
I9yzTO5/rR1U2mWaB/Y8Ohyepr9d51ssqEdCXagQb75jfwU/aFYtDJBa2aaGJ9A2
+WG67APnTauDGBwtnZj9yLEuQQtS2/NYQoBcLckVyNeNoe3C/wnapkVIDH9wD67V
LeDm7kLYX1GR3qchOdaZ+XNpk7NvUXihuEx/E98OcGlTRRd478ycvh71oJq3mUiM
6LKiTOpcJoIj+qoW7IwKP10bAk6YW98i8og/gb/vkxGq/fwimf9fDLpEEPNb9wMt
ZYIf9n/OQJfrLYQcSsgZcTtrKXgmMedgY18kBLsH1lFOFLwfEkz23VHkwhgRvHA0
6CmHhXt0oeeB0gaiop0w7FGD5qS6exkTQAqzSxL6rfxvdO3wwazOBT1aNwOO3x7d
xpD1EskdOARzPKs5J59aPHuOgsyDyjhKGRwrtkc/pW0IjOFcaoQGovDSsHr0Luep
8CBXFYgfS74/n2vHd0fKiwrfhKnunI6W7eO1z+RI9oJUhrK+k5O/2xIjWFV4GYqf
IFp4D/5KBkF7ZC8sDx6PZr99JR94gTlkTa1Iy2ows7cByZGAcPMUSe9El3mtt82P
PZtfmsW7Pj+SzvD4hlnuamx3UAZHUGW7EMBr4Eyxaqs7lS3WK394/6wpsHvVwH7O
jAJrdA9WPQ7SXcK/Lewb5QzB4DUK4OidBxlCdiUdhE1w7a1xXXr8Y0t3ZhpbPdXH
DGf8lYtX5ImZTiAK0k7qWSZtIO0x22f0PGSr3joRN8Yt1PTXypFITawSyNNUp45Z
/tQ8+BFsUfqHWFmP0THWuPYfakrFYqlqtJUmaIP5VF6EDt1HV83L8unn3iYGlp0T
Hjchx8uPweeFF+gvqxIwRhFGnLaIm982Kz1I/L0jShcO4rTRONrIo4rjuPFgMAH3
hvPGPZa7ln80mIz8bF+Y5ScXVPg8c6efVKuwrQ0h4mqjTrb5TmVuiWij6sD4gdD+
V7CsyoNHa9X3epdRzsM81/OsGVtdxHPs0cK9pONJQAZJV3kqBr/9+TMlQINPV3C7
ZJIl9iXNmF7ertyyonYQbxaQWLJW+1njJCgVW6u7fOrI20h7gOge/6E178QCDsAy
6OLSzuZBKo4wAJhRFJNYDPgS4nnOU+u0j3iwxUYTfSPRZ+3QEAS+n5t1WmREN3D7
0lttuIxRmOcTYVHKoOBsKYXT3XYnOlYzsz8kgECUMWEaqgpwO9NNJxlhGwdyo2YR
RAwFfl4OLcl47OVylq+U7JRzpygXFv8q064ZAwQPZ6oVffBJht+JLApi6OM44yvG
NN6uES3VfRaO3u0sEaFSpaXVknqKSCttZBjcJEEkYi8WVmUkSCSSm3ebPyWpWZPS
a/siTF9OxraLq+9B32KdDf8Cg7UYbsw1DAMQOyiwnczm3Oo6NuTgp0VmlUgiSfXa
fLIQTpIzOrMg3dUK91MMFYLrHTARp2sspw0a5Qv6cV4qdKAAddKpoPjda+9sDJWE
cyNcqlxLyprauG2jfcz5svSi23e8f+0r4ADounrc+3b0RFx3MHNYGRTvWeH+Y1c2
6nj5YILUxVjGFBjBSxYAfecqWM3fpoXY+Xey61UYYfXDPOxpppRRdKeUwgGZK3ps
htiuFTjU5cVf75TXgeKo8ouGDeGlTpB9gBlXU87mzWNpaVCZkchKGt/Fh2FJxYfs
W10/IUlbvFRYdsoffxJ8QfjpY5ECGp28o6moBaV9mwB0OliiI3jJ2S7jCBg5mZE8
R6zmKSmg4vUHLBBeOhNtok2SkIawvETc2nXD6qfhfdTIXquVCUjrS/26SOxpriO8
Tzi+bKbA274BMNXpd0B3jSJ2Gd9WuuG3idAGefuNTc0kR7+v8r/qZPq4IcL+RqFX
zfPdVwO0ZjCMsTitB6juZoFLuqKxz5q19EOhpLzP8gMj2FXfXY+QEquGPjqcjakZ
2f6ghE8LyCI2kD18uL++k3NO+q0BwX7ZLTwBTAIrVZUiTVF6GLz4ZdIiFEqvdooE
dROvdsc07R95scXc/QQYXuwk5a2HS+1bGhlKMcRtr3R2CMM22lUqkIjxpXsIYVpA
POzDmyFaEeIzqPbhkPPU8q8Urfb81taiYfMMOib4XINiVH1edJZywjcozTY1ga6j
ykjecKvRkLF9Pl7j/RQVNTJeBBMgSJIzG5fbB2IswM922WxR+uIbM5wzcPYsEfUv
5xAL8q0BuVVUchqVFggZ9NCFNhJhnPx5AR2mpflQ5Jm76SWKo4hQlWifi8ZzRAjJ
E/S+G8bqnRI3PUFrGz/VV7rvKsy54DAUQTdhQUWRt2D80E8IJwIfeljRH5bAy69F
5NqB4vmJMr3qffy22O5gqDFzzF7ACpXBcjWryHrJ7aDZEomhQEzlcGzZXw86GADy
FcvcZMYRkcK6wOosTCzX9FbG+ZQYipH+Lyv2Mfz0bh2evuSfRcyqJGl1C3ZCFYWo
gPXsQtF59LjplrBKZTHIW5CFIPh1Pnku5O3D9r5ZjmvMQdBqH7UMCMIdB3fSzix9
p1azoncMQCIDIejnE+QcOqTz2ZebdOhFiybUqRxQa0k9ltWu+UgJcvi2u8pc7cds
1eVKsORzs4Lcg6fj1EzIix/5SQKi8HhU1ZvgW+chHfGHA+rxxwjMEglvMHGn5Ful
InuLtj7Uvcxy3yT/Rc3CWeg4OEEY4vU0Qtp7yjLJWB6otSrnICsVA0bPUxClQ4/0
vtld8j5i1fleK6u2AG1SvbKjMWUl2kZuMaQRqn+zqw2f6UKGqZO7w3GHi8TXXhuR
UJFHdrFUriIWzOfJVgWJCokie5JEktRJobcURPj/GCWIePsshRslbV4KcSlIJr1u
UX/yyJKQZn5aINPdZQOuOCUmKhZ61uoR4qGacIs8BGmFvhYUVm3OTIUVQhZUfMaH
QY62zeH/VNejOjgRmxf4JnLvXhx3gLXv/jb2vkvFHILylKxJ3Y/c0rB32M8vbeqo
izwNCx2wv6pp0Dy6EY5G31FFnCkK+Ykm6WJaJX3LI0AQ+hUkA+4rf4u2AlzXen/f
cFGLiDugBRneMQVf0Ymb/V/WaQCDdR+92b5jyDlgjlAfhETn12nDJbwA7tCiKhMw
xseJE5vVVSM6Lgg6w89RnXoqUEhO0tJJHuyvsdZA/5KD2lOXLLWBzT04vjw5JM9K
c/i7aZqVuyvZ8aGDdwDxAPa0EGif+55C9xTG1LWZnlSyGSL5116M0RTCOcV3S8+k
1qO3AI586oKIRG3nHWVEnbsSFKMY5u2egPfvUacZwUQ4AXpLRuQVvOUu+KHC1Hkk
HXD06lfEqNOLIaqQaR8LO+BB0AIyfFD3I8c1Apkczz5XG08WLFRPLBxMzWKEL5mY
S3wZ77+2c9Mpu6wae8wcqO+0civxzXFFIZujmpofdaPoNkgyX5NT+A/76A+Mjj9o
2exn42vIi4MxqVEO8tjfVnM4QK+qAyFnN6bYOmpeU6nq/nwR1S17OHzQZX7gpk6m
RIWfR75f9VaDm20JLJ2tr1DNCBO88IMBftkhYijxN7YXeaB8zRUEm6Nj1lthSU1T
RgG9sfc6PrMbsPcGSfofeEzUyQzelGTIAeB7gYFp5RcYzcBF+pBkDez8AGgPIr/d
qltkutmjQ2UJ6kKElO6bd5jt63Cq071sRLetqsLTNVNfbBUTgHgSxbX0pbcEwyTv
QWdBns2r9ljcee8oscHq4v3C1SIPd02Xn56G2nFk2BTVvsopscszD5yUSCUfF42q
y38Uv3cTivk7StgABgF5EnmsZPCvFNxLu93TfXacuI1w0uAslVsaRN21FdmQg6NL
dAafH09Kp0uzKOenZRK31vEU78q+6UfnI1f1suQzTbKYqJ1z4a00NgCNRvFMnsq4
pRinDOSZjILLPLIlIf1bV6wINDq0P3sm8lccGUEMJk2/leMy14+NB6l/t/4XZaMR
hXtx+8ZS+ofJGbgYVuma0nP8hkURcBVVxPtHm+7g0u7Xls/18xhYPzqGNAj/LcTW
qx9CoVqrxpzzqvFP9xXN+ORuKA6QOMoxaMMT3CuACtsxjpY1ePXXk6BKojx88Ydh
9CI//gXeh5U1WLpkzf9Ph7/BNmd8kCfupsSECL0xLpePOdcrUaT9/bPS2iUVVQnn
iWVTD89Qut9PQKNoxIpiKIyJOMtu1PZ8VmMXmRJBFaUVehULHHLNjyNoh+jwkwoY
PCUWSyRJxNbXiBtgNJmgLrj+VbGl09RnmUuyRs11b0SnR9Mjjhhz0TvdjnU9sxdh
jF4/a3fPUHTWnpC+sPDiJ1Pl7WC4kXYd+ZZTCpkvKSQFmqOKiiQSWFYdTnfiIAqs
79b2PK2YfBcux3LR6DqIWaWDIa8g7kwRcRm8FObRYSlIBfxq7K2mkQJ+CX3zOVsh
5VH0676mdHZcnN5Wqk6vYo3KjubNdCiRp+ujrvIHQYOlXcbJUZ2txtXhfdojmrDt
X4xwltXNH309RxtU7r+YfqS2WZTkaOC3pGcD3cBRbwUJL6byJZjrgYp2S9S+vZu4
xe3waOxFoCwmrPzCig4Wzr5OvkEjy1KvrNKIz5E6XgKWom1/yoA6Llzucs3DChBb
m+T/kNdwFElaxT79ky2ZCQhEX785SVGu+4l7BWQvNBlUvw0zLkkLFLn4jdc91fWx
JnuukgLWwwYBp5K3nIJjF3nL+eWOBgFUlldGLXYq9voz1J31PZu0xcEPKcFvlPvX
J25b3hvGtlG+p198+XLXmxsofp32AY1lyVrgRAIJOgZg3mxSz09/7esPZ5wk5JM1
rWdI7CsVta2Vj+XAmP8BSkDMW+KZHhJ47MUd0mLegLTnCYIiOUIaA4aylCZHAUwj
uKS210qbXitx3VQ2ocittRdmIGbw40CB1FJFoHGf3MjmlpQNt+DjSEHnVkQBQ1fM
USKyMFdpwGceVruhPc2qqVhBnjMX+y4Ok9H/t252MDSlL30XcfMQQTHV/4jIRkX+
90eTiXgbS840+XMSR7htlM1splL0XMmbt78G4p1t7lU5c+1jd6EWI60LdhSKpb4T
YXD8ztgE6opEUHnEMikPYwa8PXPsYx9HhOdx833YtGcdHYQnXjac/2KbjMcn61S+
uj9Rp7Aw6nZvTmKFukWmJCY62PB3Ng267k440yfniE3lT6DljhiGKZPsHfIBBnQS
R1/dfWZ8luAiEum0/U44TtSk/n6xDvpmEQYSL2smIWntBi06OjlxlDHYfJGbPmNO
dx7vHlsyaoa4ZjqY+CbeAYe5IiVsncwr4AGt8mkxoiAW1aqnPfFqKwba4XhXq/X3
t0KjqM96LW7mk1p5U3Jtr8S3pJv+b+T3657QPT1p3nMUANyCNk0Eay7HCZndKkBl
wAxUcfzdeN2w9RiVDQ2oVRhosAcLMnv3eeGYkO0WpkZW/pb7x1JORVAtlCuOLfnv
BIjgzSNg1a0xAVUSdSB0E2v/YwjjiHS/KXU9G/wRO2CiYlEZ9oLlEsUsp1Dm5hM5
Q8bWzKopxWgpssx+efsW8H5+Bq+3271UIZu0VkAFZzmoY/fkfub4vzJYnZ8JytgX
qiN8puzkZeO7PQC2HSCnK/vAcoNgzNHKPJ8v3nYUDBYyLH0OYPQP0jHLztmi4pbo
Eu2vD00J1BCxP0mtSGzV4Njt7xCebe5MbSVNsCvnA6UHNSs1k2DEWyusLZKywtQ1
chGqRgVk3sPRd3Axs2I0DlnvE3l5zhYWIiW2f6poLgd+a76JQvNUAQCNJ/vM0mD/
MGMiD7AICZbi7oymBnPh9I0STAHz7v9cshkuRPAnUzKfGeNqgHuXleOIwNKnkmPf
xh1NPokC5xU2scvs6YNHBOr+uW/nXV4ZceMSMnSeHKLAqGsuDquWn0CDuBL7cPhp
O5oNN2WVSEflQwTGkPTffTiHB2MR8aCIPsfcb41VvUB7yVZCQsYRU1UFASWbVwqj
X8pIZcbjOUGsu3z/h59YaEvNjNe3Gi4CiIYttxPw6aINsXlKEmzXmnPgjEXarsN/
3iwldzzFCT1g+KVP5KRxby7Y+cxvGfd5FgHr2hZmcSTbb3U1nKw1mRyM9CluMgZ5
wAk0IACnxCdMvBRMJPRQU1nlxIhvOBVdP+tk09CWoNSGRWlhbXz/TbDKNpwdU5Tg
yBa32LitJorQj/Zsm8a4XeMKKSN7tCEgfng9zQSQk8dunre0D2PWFMD+/YZUev5D
bf4Mkk4b2uqyf0q5NbvE2wAz3n7cUoflWiYNT+cqK/n20+kCqEdGGpmjBtBhU/G7
vHzqhTceVE792FGQxSvfxCkCGEKKrgVPkp7gw/4IZjhbBCrFcjWzUURcl/wi4MqO
WBq0yBex5ihc+o0Q/xZzB0oh/BFnP7ZI5GhLfxOSAqSCXEJhIEbemifeNwnUUOSx
qbvfl/IJmUmlfkkrgVFIoE7InM2WrqGEVDxeUInGxj/7fyGr7K65GMMp2OxzWfG1
zz7oDIC0ZhHMzoTUWTxlSPKpM8bgPE2ecqktUDTADsquHSyQzOafXlmh0lOKAPzs
ooVVFY0oLd05V6BW6gTb8YNDQDQPIA92do/4t0dx5zeDtELdPSzJjAQ377vXYH5u
KI0Wys7AIbaSth0OD5i4dt9IdDT89MGepTwxACFBv1886+hhrbPEimsTwyDKYg4T
s8hOlTYmg18hG1bJ39oGzy+4AlgMyNVTVaU+u5kYz2AVhKifLt2g0UOn1rsHuC5I
HV1s2PsyDmwLDvi5d3uXFOvk6GYKzRwyb04Z+3X9iL427qRFzL58B7gE0FCeSkpu
oyPvK+hk4Fi+nZioQ7fe4F8gB1iD69W9DADm0+23EG0NakunLVdYjz1ASIDdAXCz
CiHcKUKc4De531A/MnyxFjyvNfzwFP7SGeG+OjieCQGu/I2RmGf0l7osP6oaNSr/
ldR8fGiLbBDWvQTr7kClEolyhAVqFvjQ7uiata3l4MY6la500HjoGipf3jcoI60t
onkhS23B/8b72ETSXlS4OWvW4rW2NXdUF+e4hlRArj0Lk2AnYtnP0H+0cLbj2hE7
KKHbSW60vcUvLak+MZLC9JwA63d1LtsQ3ajlTSSIJq3DzWcJzLVOoJDGwHtTbNg2
FSARdAXaShxxwubJgu1T6/qUhJjBSRDbKzWwmBHBzBNwvwAnFOzmM86RIGQgjqym
uGefVyH48E89FbXd1rqBs/KHHqlzlA0mrF84tZkL6JwCQqWxWltK+G8aJLGFIaAE
vUgQctJNutoR7OlRt2Fi9ozZQuc/GQV5t1GZCWJV9HogFrByfIo7KQnY0HZy+E1y
uZ6pNM8IxO1W5jDfIIhctSLTkr4QKgWVfyPrmDJf6mvEELTineylYwU2c7sG0xgR
3ch0HATO5kMPeE1SXFEhW9BjlJs6ug1R+96hAdTV68TRpk3mEOGvA2s4Be0qmuKZ
XNkWqufHbcnK7dlwm9qsLpuczRKxq8qc/nDWhp/LVDGkDj9DsaIw7uWT190rpV0C
SpRX42ik4Hw/gKfOFmGxhqc5NPKS/HIOWqJ8aOBnNyu5W/s2skyJXKZl4s0gLEuu
v7PFWm0pnEQjQWByQ37iMHC+WH6qyXxjE6ANLdu7KAlYV7aXH2P7jRwLV7qVHMMU
R5q8mpq0s1rd8uwKSkhLYKhe9DP3aTzT75Abstl6k2ZH9yx5mPaP8xTd+wwKU4Ra
SZxeV6CHV7LSD2Io4/i4fMvvgK8hRK8COCpetZPBaHRMw1JcHYSUnUTICc/VlFQX
l7+eOf/K8uf2/iJ4mXGJuFNZkMNSom99mwH1LAU2MUz3Dmv+2YXClUiM2P+44LlM
T9mxN0e+jyDdQ4BeavnrICLD8p1LG4wYIJyMEYogcg+9rS4PqYQ63qqJNemLjuPP
IO24IyJGmJqchxDK9wB6ktw/arH41jQhnERLCFdM8E+ai5Nycik2hwyzr/Vn9dle
nKZoo7SUpmcHyptgk0V3Voet/3PXSCC2woYTXDyut43GJ0JojXgguV9ul74rVlIg
DrN4hk0kfe7IPm3gjoFzG+kUp7XHTiyEOlta47Sr7sspLUaI7q8aV8hY4QJspUVA
LDuVDnwgSf2LZra4eXBixR4TOgTKvcNxgsX0cQ7bA7njrZWipwKp9CCZTcu/oKI1
hW4no4un/LQ7TsqRlQ/gcBLOCIk1QXQfrN93ZcFbrZzNl203ogpDWDofc8q/GMAY
xLVXCiO+PUnvoeQKqOvFq7fxvGsQs16jo5NpZOYs1ZruT5K6dfjmRHlL+ph5srdz
CQD5BLWjKbK0vgUSJTqDwDKRfJ9WIRaBkce0DaNAxXxekyuHE9D70Y25PRoK34Iv
tOSUOKA7aMI8ip1Ti5gHqvRDKJP3bNbztUOwZJ3OthjvQcCYTSUM2ZLfF39nzXKW
l/bweVJyvcoylS5a/xgUVHImE1/wYLrrKZfat1m6EPrhI94EdR6lV7jPNARm5yP/
dtRSLbz/8WDBUwBEXzrA1YmBfv84LwnoYFczywk3jctviUeJdoSdsEm86jS/RUPH
EuLfo+6+8NGvMYEBdDsE1zxNncBJmLcoTnimARh/IQyC8J+9igtzeSssBa3zNUI1
S+43EXS+r/dQiAD0Qc/H2tJJcc1iP0+oipEsHkQ/thDXb709YUgoYu2e1Kca1j0f
HK3NgJn3ij9AtoNAf8gmGQ384lTgZ9MHfszivDP2jFESD6DW7QAQY5i5nQ5sMpNR
M1OQ/9TUSAW4veUje8mJrcT1wI0kSU/93wk815N2V0pdkT/WpSwMHshOiHRxUrnN
EY6eanMXOZEVf/dbtcnb9EraDscMVVI587Tfuh8IHq2/dHIvgcW73BXePRhiK5NN
NIDdu0nDRfhv1D2cfI1uPSnGPrXRbgtbz3R6wcncLDqCKZLf/Wr5A/EByNGqHlSO
0iTzCgmCyXEynd1MfEv3lCKHcQhC504JlBdU1WCRZ5S7MCzMns5q8SFKAQYk8uK+
GziPNeL0sqKBRBCToye4fhymo4RLi/adbaLtr/aS4P9DirjCZv5OucSNRY4UvNWq
5FaV1eAG8M50joCOm4L1kFy5U/tuN2fcM7TtcPhdgEAMKaXZQoR0HZRI4kc1WjUv
OHcFpCvBfdUtgxMoe02e0R9D4HfhIBzGj2n9qDMobK12yMF20zThpK0s2k+5In+7
V75/UA6mlc7iGfcKKzlswNfq7CaZEKlWu5KsrY+ACszoswyIGz+SbmlRQBlCFOJ9
BgPBx8jTWiOq0fi4E8oh5TPXpqkleKnCN4lxFu/fEqccVpm7oKw5em0DU9ch2dKi
l6UYjhhUAYthg/xmszZoNxt3tiKW/IGBbRIE1Wbh9Jg8mCyo/Mt8DE+elYKCTonG
/gyddaepuK3q5ZuK09sF7/dFy+KJaRMRAbc5ajK8zTYiYjTCp7VXVrQgKEIj8a/Q
39Vw2IkViNQRTacr/04qtQ==
`pragma protect end_protected
