// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 14:01:31 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
EpeSpqYo+OlHfnuYoJ/Ogr67/30NKE+So8zucV/W0q/M3EI61TEFird0Y0CSNKgL
76V55fPPCY5wxfJQ9R804f642ELsb0reweanepjhhDUKQNx/cZTkOvKk2QoLwinJ
zIlIp9fbniRu24hRkyUFT0GSmjW6Ali/KrLhLOkA90I=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7232)
agYXuKPxHXoIbv/PALcD4FkZoW7esXUxbPpZe70XjlyLL3Ylq2aCrPUDK2pMPqPM
v2936T50HSpeWUvlmSm0sKe0S2MVJvJgX7Vg6UOB7D8zybKJj0+1Tv/Lg5N5P2+V
LayHxSDtxlYLcDuQfWnE6ax4uN1fkQepWyPI+llhlgveB7v26MLp6VKRxTbduIr4
ZiBIu2wwHnt7WnakQz6aMcaL49gD0RZZ2spKj1x16/Q3b/oUFlQRUpX8r8nJ9hSp
cEjvzehklPB4F0kJzitXmXbyhjbXIVrr+JVZSqUWnJpg3T5sMr+cI/j86aBsk9rr
TaoIxTW0kx9Q5KXRrQrNffvWLIqmpImX0KTrBPLm4W4S9bfVsX7fp3QYAc8QhGVr
G5lTnfcIouoHq2msPYAg2d7MTxXv3QtQdcFIrUEG4m481LEhAHDbkRM4TnWLF9Yg
vVwUemWRsyrrMN+y41d17B3x85VsZQ4tK+eJpOihQOFbqTNCDjtRgUbHicbviLxP
5R58nC3w/DY+r7joDYtiDNjlIqYMpGJwyE8qOK06rCsaSyFJIdjkgU5LfdkYrFNb
WPiIvQkfkg+5hmkihRQom4XLQckuJUF3RJlF1cX5AxKrcO5xThGP3FdUuuf+Slj6
0HJa9gOSh+5R/7fWIrmc3fMT+XQSCCG1+PtrhPwX5BZHWfuZC5b4xsdji9J4GXeM
+PDaA1o5bNSbHXeRzawgcxPOFm3IkZ06oBa2m5qu3ViXR7Q/2kR/WPWYiu8Q+uK8
6t+vZO7CH6DHp5FOyuQc1E2UUdSu+B3rYHuMUe/7Z5M/rHGqh21jvF0Mq84k9UDS
awSd9KfO4GzqsOx5oPRtM0ntpR9oVVRR0O1Szh7hGke7rKoscazugrYt+GSp/96p
P+iSHhEwuRms8AW1kUbqSF/GkPQlCIJBhj+BN0ZfOxkJXvO2yvhlWdBAVD50yXko
uTPB7kspU6PQE0P68jqWhwNExOAApngeob9Ss4g+LKC2tHRNHAGVCue+V/fhGYag
5iqVdnRKD/UX/xHd5XNS8sSHgBh61/dkmBiTnUGUDGm9pJabUYXnrKGovpG0cLr+
2zBX8Zq5QFxwv3YEnZxBbDhpkgfVeFt5WZdstC6qBWqXpu+POFKMoNh1zH9ulDJM
dla+p4jRBQJYrlYc7SuafpI74KvpOvCG0BUNLA384WJufQtFo7nR+OVIh/ecBcKS
W5lID+MDV+gQ2OsoaiQ/6fjNi4JB5+sHuYmSpgE0+1J53w28uEmMxsvU8QzOJBDq
Gp1lrUiOTCEKd8tMb0WWkKZmywYYiBtBsdVnR16NzXA+Qjygt8adCGHWuib9W35y
hyZPUWaj8XhuKWcxd2f9QETXEtmsUf0ZJ6GH0oYIFJUFpmodZgQorcyVQ/JdmBIp
FdZnZgsyAZH7vgZiGL49DtL3ZWk6DDL49N1av6mFCvR1cifRaB2COwLMReW77plJ
/X1BkuA/0a7ypmsY7xTH/f+mknVbvgc8aJrFi4lyaknJDjOsf+YVu/J/XLpk86VE
XWebYlyKoAf9+8oEMTKtzjSlyMIuCsAFHzbEsIl3xjXG3yx0dB8jVp8BTi6Tt3M4
u04nd7LkyH0pYCmgsyoVqBcxZ9kPk0TfLXONFOyUMX5MkyFmtq6YhyL9bopGQrsb
YDsFtb7SzTLgZ96WJ4Rc9r55zFRgevVRrCd2ZpwSE22cLQ0JvtT65CVw6sYGxxn6
G662w1fYXMMz4tRt/UbllPOwrO1OwQeTApl1wrhRa3cL/KHTMJsmzxh2pABHIRTP
Yt68p2AtQB4THq1VPc9e/jQ7orObGxhQN4Pm66NymOX9IpSyWf2fbKo4g2JrYUpM
7DNUciNePxMQktefjJb/X9JFp/iM62sC6bUB5niWIb1hbg47XKiXKX18FSh1TpKs
MOVD8nXfYAXYOx5YhsYe9LpPEOrHO4404qQH+iKwXxpXghQKXlwn+6SbXkmTk+SQ
jJAmRTKNQop0rENEOx6eoed3dIRChbaNRAZV9Tc+kBBzIUbgGb28/e9bMpvdyCkv
ACfHBaQ4UA1nVIejWH9DDe746A9xx3pj++mmylqbJzkq00R3ImHrcrYa3RPAxUpM
RAolvT8tGzFr3k1lkT59vfr8fvJYdlGNn3H5l8aCKI6bePSx0paoKt5hdrOFyU0t
f84G79M/vSXvorPQtsv5t9GcRVXheqFjeZGHLByMCgszsAovKOeSkyHbn9PjJYQx
O5OmMuENqwQlZPtf6Yc8LBwgxt3idl/Qco/2wOjdgbjTaAOn9bwev7xDQuWg57mK
BZL4KAAUo61Wo3fo51JfWGuT6vNJvSR4uskyUhXMIyH1UcsJBu/n7lbwBnN+ScIB
fWuT6spdDkkzSk8d0rOByv1Qu4dPFTXI3Iq8jDr+vslC2fXeAW9rPlJWtAQ06EBx
pPrmGN1hDXRgy2m31Jg26K8kXldUOogwLFzegd1HWyok5jDlf+VP0pxMmSgJryfm
0hE/m+mOKc5l6j4ukYQrnSGpALIge993rbMKKx+Ukb4d409hmgtkKYGpcXuWpENY
x5Ague6Sqg4IZ2Yno/UV3SNOZnwJzx1+0rpNCi41i4PVtJoe4JYnquc8NZCXm3ZH
sgW8qkbwtrBX+sZLcnkk8hLqxyXZJQKPQkzQaLXC3haePM4EfyIm3BQZrqygPq0L
X+kHkdA4KEGvf6v5CKGAl4sNCgmisMD4xdwHJ/08cXA6Vrb2Pz+LvtWlhWCMw1s/
//dHpX/T2I/lCm7JxC/RsbCOktOjxx7G+xQU83UWB1IYEkP993CMqiC03mCj+f0e
XW12IIxTYyt9Fp0MjCCso+wTD9OPzZ4gckl2MhZs1SHyUAz7VItuPO1pEljMSe+a
S4hDHB5Hx6IE75sfF83Dg7ElSTNLPIDUTWfacgq1wr7xpBS/ee/O603HODhA+1yR
VM6aZBozAyhE4rloT0F4NzgtRBVxSGSriPp+95M7op83NJTn/hqrQgbcgbh1Kpyn
4PXaDAUQfMnEIbZDsoeWgMYJ4opTr+KHSgzQfe0bap9KNlQOjaJ5DfsmpjbeZXlf
5/H5rxLUSua37ZZjapF5oxWquiwx+s8PrRbxZqCoRiDj9u+6Dt+1t56IG7hjgWXp
SxENG/cgu9FQV+2+nyWM+jGd6qyeQTCs/QAUwuOxoRqS4ca+/AjqdX4tckFmKJOv
ONMuckLygDMj6ph7tt74tcLNAKvP5+O+CCeCVE8DNJqdJohd2T7S6NNJMeDJGFDr
fzY9kW7YsFopLmhcM3T9jKv93A6bu4zySPxVQyieQ4A0pAG8rWeSgXh2/HD3YaHI
K8fPLKdK4aQvmDta1DP/fWcNw2wXzTJtZ2KkV67CD8+/WCv4SQ4zjQt+ikT3jCdC
+qXrpDfXk4vtye5CTXng8nC1j8534LIJ9Vru5KNO5TtDI7ogqFSnLidtGpJtSKTc
Xpf+2oebsh0y3IP0IFQBlzn8FD81RXqIE7RsHySLBSLvTAzWbxMi7TbmjI5GAg1r
RAdU0PT5zQVzIcyXyzkj/V2MKa4lqV7AIPVTJPV1fozRVtjTmHp2rOk9aZleP8ue
1USOFqig9IIahUMWnlIf0l0DsakZgGoLnYfN7ao029Kmffz0DHVeDQaUSVayEQgM
7eDttPGZaYXRMeupnkz6g5jYlk02E3K+R5VWhnMWSTwuxFEKbnyJdhjaZ2mBuN8/
tislPQlJDxl0xdXbtCTrZgzoEp20euZuRObvLpZieul5nUu4Qa2pyshngdohroHb
ujnWsVkTRAL5PwuZwX32gxlQskeLtwyy7ZVHVdEGr8sNehEi7jVu7tGDkftHZesH
SZLUSyRP7JKN+Yf2fXvBGAy5yTYOES+QYBdLuoLpVloZH1CC4XOQpbwabo1ZMN8d
YId4VcnFLEYWeb1MLMRaIRBlnk5yPSzboTTi4j/17WI1VB61A6jL+FOCgHdpU8Ph
E44MB5fhRbzJPH87zj7RxQmUnNHL5HLcHQsUCYaA0diRXvhwudILbOrMU742M6Cd
WCtSnJ51zP0W0QSkzxYcjerWBvejx5FlLDnXRVk4jD4KtYbEcjUCf8OTUjNIrbMu
2Y4TvAh/DulqsrckmUaZxZxJbQPzdw3ZLCB4ExqgjX5WHTgK0duszHnfgVDzVvLY
XLlvz3Ue1cGYTMw8sIp0O8bEaxJfDhNTyo9Dl2DXHFEnrvZCNekkUQvUNoxgMjaI
MOT5xwAbcJ9cqz0RvaGZl9CDl3kZ8ZqP/PK+dMga9lTBljhXX707pP+EkXTHWOCS
2uj2IaXouTwBiP3VA+k+AiZe4wG8FiTtInlwddp+ieuTZo22ncf1gK/H+dnmw3MY
3GodMglpAoIHKOCC2nC2XgJGePrQEeg8j5M2YMWMMw5HWdDm0DwW1+vy3IqF28s1
1jRafOKLrgoFFy/D7gllnt+WpKuW6NkfveUGK5GFyD+P85KmWh8wXv9jzXICvZKZ
Cv++dRymZZALJ2SvHhHvCKpkxpk+X4OrMUszitH+dp/UDflfK3sTP5fZX8rCwXzE
lBZoiHhlZdumE+dw5bpuEuZzDX3lNWF7fIBXfRadApG7mCv2zdbR08HkQMYHQVbi
MjUhkJwY8r5U1tDVe6ueSXg3os/CpGYpq2HT267l0JrSrhWBr+VmG15+CQU5/zfl
O7OgReMhsxQsic+lhU92RTB8ziU3BRNGRlMqJoTgkMxMpnSLTdZzC50hY2Hi8u3s
ivx3ZVSxQuAsa7pxMYmMeSN0pxE0AwQwLb3/sbOXpfkWzoPQI7UXExYHeO4SBFqH
kkkqCatA60YQWojBB00M7OWEN0I9UqiSDmCNFE0NUKiUdzEqHntPrFhhFRI45ysE
a11Lbor7tRnhJdjKw4QQwazzF4ikNxh/2FhateA1pYVRCtJ5Gm0sViplPb4PXDZo
woaO7DLPltmSYgrmJ4OtS4nq0e2VVzYO6M9UM2Ei1wiuyOVB3BQEkEQPk7916bwx
1OqvOs1Tj7uDvskFaXYms7jHseNkVaJBmlTiYHxS+HpsaV4KzOBrPIJ9eDqG/v9m
zhO0CY80TSWvO8VTo5pql34aK+Gp5qWtKhPVlN7HQdSW2Q2SJAKeBnCLXyEdqM4o
Ws4rGQiMTJBvuz9ANuTaJrXlBzLoFlZKYjh/BEsOTVxZpDVJQAAZXt9Z4x73Rvfb
xAzAyinE/nlVXGpmUWVslT/RNO1m88YyUPZNOUBYWA9NhpvTR9NvpJOFEuoVM9DQ
//ZCrfS4qa0lPDtzC8gqWdSHiKoL9e+myepcwYq/vnXGn6VkjHM2JvC574hzWk/0
ZgMpNewpzZghAEka1IHb8hAuMP7TaQ5q/9FeTFPtxduBr1/CSEvSoJQydGwbPQOg
0yUsOP/MZ6bVNFcebpdDKDgPuNVoQWNb2K4JCn0/ElyIxmFfkpXGsVmjJgce2oz/
XcD4GzuHRUcHDq6TVa3RbDOwAqlwtbyxvdpCzgay9UwofCfQ630BVYilPQBaV/CX
raBCHBvgeYl80uhvPFBT+GNU+zdgWVgFpr7NhPgVDQHuhteyRTh+dFPJY0Lc3dXH
BYjIfm8RyxGCLmAPpL+as/lT8PKTZsv1hHrhOEEDrerKYEKHSO9BHKV+9uYR4bRx
mFOOFxSo6ec5K+sA/1s4mxdtFJcQXhlx36lHaHzgg6eIgWWpd9fxN59CLq/7XYu7
Xa7mnV/apvKXJpS499MG9569KnGVW0RifCh9iMPb0q8OE0Mato20BE0VXsKfYk1O
TzZtPCVwMyR5coWNAQuCapUWOma2P10x48sruLTKKKSIFQ8Ohhq+2eQOh3YOJ6BD
Rn+k9Np/nrE7/Vk9NzmGDe1x9vI38/wBaj9LfFaLsgmlz5Ycu7sMvgcPJFDQjHz/
7e5C4mx9vOuQ104vd8Tp0QJLnXHC86yKuEuYbOBdyQ33mDDXx5YIOLwmvyPMsKal
ZRVrir15ZMamz9/lGC7tlBRu9RIBz03F1lBVmIOKrsSGLjVlTz+Ss5PGOIxNm5VT
XWJkKrFDKUzHoKXyOea5TFflJ4d8Av6pwUktw+grEtgWtxNsNoZCmxfZElM3wBKm
tRzqfAenQOdB6rJ3Gc8dLCmFrgLfPd15j4dS1XNgbZpJrW9PKlkq7GnfbYA/axGK
5PdxigDXzrhzG+yKW9Bp93MeDPz24c8ENgC/vMyUoCZ1sL7AbwL/99wYxUY0KiA/
pTy+MaLigPDAJFW+kIcfaimY4Vnc0B7AcNivkkJCxU8+tBLoMV5T8Ki5PzX3iduu
/d7w52hFS/DVfzskYgnqIHHTDOV87J35J+3umSeA0+6DhEwgbO/KsojzLmvg3tgn
MjuURBNXkBpH1pxjbFXMPeW84FDbEm3+rFB7/UoXPQue9NX/Ymn91vgNo2XYgSCT
gteMvxxNcYyCxfNQKa7PQa1w2VxZ3IwA8sYGTgLWTX8WLL//lNv1x8GQNulxV6ZX
QqeXNs27u8mlGKj+n5agrtswCzPR//HGkNKsrGb+7grEjSg7UHCqGmPmLY615L2I
GDaPakq4TT5Og8sdDOKWgfdFhdjSLzDCFacTqwZtwLQMbOZAhaRbqiXwxtHuwcGm
2O+JrgRXqxaisDGhuD6Axik/FJ7NuLuxhy1BAGlA7/KLJH/OVnsI2bIL2/u8jNAd
2PbDK7Uw5FAEhNEHBglfoM4s/sFes3GTUFTxvk8ohTeo4AtEFDkkG7pxRqUqxoB/
/SE6eYOdoysvuB1vYn1RpemMMI+WZFNORKhJZr/5mFQVN2IJ7HfBzyzND37rCgWd
pR8XKBO1owRp98U/kQlEMR5IBfq+boA7At6mmXKPE9Mw12rGlIgCsCRG0nAGFfvd
9G/EjREoLOrehrEIDXqrYcTg5+cyT7CW8nfsYX2s7z129xFnaqe6XxBVZyp6EHKQ
2JYeH024Y6hyRgL9GoUFf87WKKU11TF2N26zrvI6Z7IFs3eyIgpNWMPYk/Tf1Dam
noxpUDV7ZHja7Peqwvg23g2egIcsaAGiyMl+o3qYPaz76fOfv5bxxt8iXKlkzqLr
NV5mThvtiAUrUCxAF4m7e+hxR/GF4MebxFgf/TWNHfZPjgt3CYOpnrXXQfp93oKu
KH36IjCnPFB13cDBOjk4xqwSIJKmh/4Gm05gSGZovOhulTE+671+37Kkj+WlisVC
KJ3ss0XQNVSdYrKUxieeUAGlwwb2SqWa9oAIph/ySch4HlEo9JVYgzTb7PQL34KN
CKyU06yq8R0qlWdXYtEbvkMKtI/Ilqwcl6kyhZWBsZ3L6zKG3htDOSyGsOUeuBms
OcgCdJEI0hZRi9NuVmW1xGhDUEO+W084b4YLhsmROK9WHS7AIJiBr513yBcw1sxa
g2mlu1u6hsLCfvjZzjZ/cGlYhcoIkpvuCCAzUbPwYYAvzY23ySclKhkMXSkoUM49
XvZ2Qfd8PbFdGSLunjDC9spY7QOfI8rCVDBmedueDtFsZ5qj/s/LReLofZs1cyic
utHhhxip+1t00sPeNNqxVdudKFzR5m6D+pWRxvSBgSBfue0SKfmctRoxhxqdNX06
c3g496M7p2X1fYUxAzBOG1xuvECXEiZWTxVl8R70Ox6f7AV+hf9RoMf1dhr5vLU/
zhajoThHbhGjEx5TSlJIO3fehxGFNvRRa58sM/F5xo7qtEzNmOq7n3xnjZsWEJ2y
EBmuUIsCDgwhKujhXGOO9SRBUN2h9x3fms4/2g/Ww6rmnokInXklEr9Ps343Dtmc
CY22GbS2MQ8SuJC7dlvifUaH9keSzX08RH00QIfgk0dgL1856MdoVfaO2ZnjIghy
QZZL1gN8kwm7pW4KEqJ2C3V5WojPppw+YicJCA+29+g4pgRzQl7zgwijwzQjFy+Q
phfdqSb2R2KTGcPeAt32oBTly8pv312PR7ZblUedX2wvS/eZIz+Eddr8Wyr6l0of
Q0siUBx+/x+3BFsjUh0NGIUzXU/JatussW9xnNUU8ch8F1alQ71kUF+Kd9mXAdfj
jfCarn3qPTXuIacXVvPTdfhrW0vKR91xv61iKmJc5Bp9CZeow5fkL4OdZb4lvgs4
rXFvdUlM+yfgBrtdWjn/YGLqt5HXI71RsUJjp2iSPAmYzdLvTgiZGoc+LN3c/RP4
RFoYOiHaUFG606QRmtZIZmeqGfqKgPEtSvGSTujUlyxt6+GRzQ0TcuwinM0LtAdC
KWEcaRxVUcGbQvk7qdvmpeOKw92m7kNw+mBN9iBVL1LC/oFztt5+nKduUs8t1s/M
ix7lb27hgiBPiSdlvZfvq7keYcQCOihb9qkJA+DPaFADBKX+itlO1LB3mi5syq6B
UeoFJAN2gpfLRrrX3BdkCNZc3NWkRep0ad57dImC6YS2ZRDmR06LYLis8pbJdT64
5+ifH/Qy8bFf/4IpUrwrwfw3lTDaB3NsPr0m4Ag9iLyUWwEPagM/gZv7oHwrP0Ul
RN1MOqunPGVoGFlzTBTYSChhVnRyCwUrxhs/ekRPDycbnmUjRwHevoK4J9I/OExO
Y4bBleScLgV03EdSBAsOn2MMfenS2au1KgHc69F9psa9w+8lxGeW4xk+Ik+xqNBU
Xag4F5oHyqHXfwtRxtOGTrgZP0c9DCZrpNVILkwhXQeiG74RqcHhUavidb1wq4UA
BymzBJFExCKWr7XNhQAyNbw5cheiPewjsoc7nkgWuWCZR4IOX2kSwObjW5Vw8SPo
pQ+re+y9KmQOnpSp075Bo5//1PtHjk+fKn68Q99GcYmRTUStCpdDjdNduRbsxFeN
pwmnQqKV9843+yZp3r15rWpB/aZMMzrS9sjepUGhWGHC5Gjrxl72AEe4uFKddQV6
UN32dEQzGCEjfX4TyQtqDfOGBxDzMMfgFsEWqXlynsBpDzzkpUmu0WYf6sXQbJWv
tVXAnZAa078JJX6mhBTS7zjobA+EKZjrwhlMzCYj3WE9CHA7FOe5TpxAsDmpcr6/
UX7UnovOcHjlXofG7Svw3RiKTVJGVbaG0MxtZYp4nDBtr1uGK9sEc2TQ7EXjYxq/
FD3MsP31aerH2NubjE0Tzht8VWgRcXE5FWtwrBJRoAKUkIFwGWnYXvJ3vm/xIPUF
TuJxTbQWu2m1IM3tqXOmsEETf0hQ1Zs/JMR4jvFFtrP8Ie0zOkPdWI9PGc2GJEU3
AthGpAblFjT1eghdZ4NMhZ1HtJLS40n2aW2cRl2TImXKTyVq3x2u2ym22wYvaPaD
9zp7+bO1r898ZZj2nsB6vb//Fhf/ae6K5qpbf94Q//1eqEhjFFX6NhHRqn3eRFZR
fHfgD0jUmn2nFEG+EI1vk3IirQrsfch5FWgQF29votD50iIxJg70aer29hkILaC5
zq2ctvTknKLn3/qRcOw8pnfWYRDFi7ZJndhR62O+8QyOfMQ6IdSyFenPXvUWZTXm
EyaHW8OzX847CzPBjYWbQz47JO5vsOMwo95aitkxcE6aL9AHUuw0dwxxtHBqV/c4
GGLiLA38nF0FL4BLYlHe93PIKu25iVb4KNxAyD1oIROt2GaODUOwNi6vsz6pjF/A
Z+JqT5QQsfricHCGWb2gGiVCxUXjl7Ig253UQxZqX9b4T3FSh/iHCSn8OA2kv5V7
UiQcA/td450iG4xSLAIx4Nbyx3VuZDl0VmXF1wI4gXo=
`pragma protect end_protected
