// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:02:15 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
H/VD1u9oJme50YXl2QbPSU4IQJEMKSF34iXNon+abQrGZrC630awVntD90BjGA1C
KrJ1flqKMBOtgIXAZ810TlgHTDH8cfdCHMViiyX78DI+e/wJDJBYt3phMus1GZTy
+PP3M3l5yOpX1JRlBkVmWwDYCzfzxZacxoH4SEoJelI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5424)
9JzfmmLv30QeTkR/+AJAx1SYWe93QaOnYOqk4Mq+SOASGyAz50hDkckZU/180ndp
mt6wCj/MM8zK4c8p4Q2Z0WDbK6oNFBVfDsswbRDbpS+KuPsdZ0oDPFsx6rSiH4zH
Bs4V5vDH6F1Y/a9H2IFaswpzGjC5et1QdSbquCtb6b1sY71FjFKZyxfymAC+hXr6
VNyuJrQ2n4OqlVJwthSKFQYBH4bJfQnxYnxJ1E4ZDWThcodTXcusIpvD6pObzYX+
M4ZfGpaxEAFesF0kvE0R4T43+tmR/kGsG9x3f6OmuChMtOJ/cDS/zl/n4cRVoPTi
nu4b0qleviE28ofuGR6ETJ9TqtjzP4ixJUR+VQ2qzKsYm03SkYxRhm1pTqy+T8Db
WQGNLme188Wlm051OLOJuxz7ygz/GOYPqV0ih2QGCK4Way5vHyQqFrCeXIe2YYLA
zRa9DkZ4aQcXM+TdS4wYBP7U5Z+2O/Bma30CMX61aCwiD39MSoS88u2WMMCcTViH
R9ynnWJ7PivgVp5CcICWCP0uA2AH4QvxpchVjbqOBtuIMHNaWy9h9KEBN2+sVAVh
HEPjrwrBTia/k9ms6Bc48WV9JeO35g7Rhu+OzB/PMnIZ0hyc49fHfhhx3n5bLrIa
PPVHquV9vUaH57W7BArPAmofnPN2yw3Hi0RuFeDfAG1NBVesSspzRKiuHW0fxUWe
ODVXapfTjuQFdjrg8cptbd2mv9w4xXAitIHRYE6cbW6vGthE/YhWmjHKmXc0SYqX
9/jCMPnw2PEA1rd3Ui5RMQ1suGtAkzbIjIPc6cSqwM3Rw61j+anWGqWsMIa7cB91
9muh26BjR3QGaIC/2mZisskHaddkS3puaXPG9zbFK3tKfmYZP1Az2jZJxDkW76Uu
wrQ4TQ+ztv1WFUbFI3U4BCQuvmbVAKhCLPw7oEcj694hlpX5lFEdN/spKo95mUTy
hhDrIB5qOOUEKbwKZDPd6yFlSa9xooIPv+n+xNA3xKC7tK2VfjjAuu4QVDUGKKWM
O1cGa5UgZsjECQTgK5vmAAVMVD80GOs+FpCkK1IrJYN8Q/8mHPfp92vxreNIqUix
aI/9I4XnZY4zCFpxkdDqJtTrEsBCIDszr7IJ2sXpjr3QuFFIAomHXxc4cUTfhk+W
fa61hUqjEJ1kSUrscvqFvrOnRVg6QPO2KqaK3jCstammNlNs0gtiG+17TylZKelr
2349dNjRH7m8Of9ruvOPddb2dxJ5Ih1wx6VNDInLibTeFV3VW81H1wnVfGjgMdoD
UTPbTJB8AUfbjvZxvCPlTxVb0ZROwFuiGUaoD1Bh85HxJoxSa0t+u/SCecX4AwJj
0wDUVKz+44riWkxeuhVxHCSA6szbLOyQOPli554cOJD6MfQTT+oQ9vFf46AZruie
AchJ2iP0JRy16BGyGxaAchzqqm8BfxHD7ZqwwMBL6/8T2H20KeDbeRs9poUA8gbU
TJMPLz76c82aK06PXOLdswGI6cXj0n5aYEHNf1Dua0JXPlCsw83+FChU4g0jhFmO
VcjXEX+xrKJoFV+gtFQtrM8fNVe4zwvsdEHeK8wEnrS2+pmGjaZU0BDcdzWAxgGl
nN2R65aHgatgM/cvL4sOvWzaqTf27vmB1U6eQAgIS3jG9yLvbfvNeP0cxLgdQ30g
5WpPkpKs35iNw1JnPUARTtS3hrQrShj33zT344/FqUKL6twPyJ8AsBawEb6lIlFl
1yKJHatEzYWITY9p6kCJ2hEPKYhvnwfCcXPQUPpVcHRk7fn7lvDU+t9kkXwZ48LM
OI+UDL0GmpNjf03E2CVKWOwsrYhSG+SnhGNtuGRFmN8kuNri7OOmUXQguEuBlgfL
fTxImHjHmLTQhAIPpY3F7hQ2EJXStQxrBS4Nm2SezMaPUgfE5BOgJQUZIom8wFyZ
hobVI++foKlmQwQRGAr5ehBpNgxtnj5mKjKOvZ126fsL8xlbtV/tyirsOGle86UB
jRw3FcNDuAPirU0yBEWmMCFY90oOvGzvZskasu4WL2xzUSOSv8I4nSzSYYFJtxNw
vuMgB6ZImNpmVGi7TRzdSnRpJpYMLBVdMqsdU7ubKBXNqQpo8JDTViwtD9Le2UPl
93BQknRy1WWZOGr418cHuWL3VoxegZpWGKePZB/CVmcJpx9+P4iBcN+HH1MzhWHo
N09bSPHuKVCFu+Kbr2HiSCFTw+w2WYg4SrutNLk04WImnrwiyBrC19ST2LVYtssr
dNDpClzKqu3HYG0Pk622O563XVsFGrhZSxF1k1KkuIgFk8QZ92IYAlPepAeu2GsQ
fnUxvEC68+e7vocF6D+bhM5qCOjyAg2f5itbACGDPAqfXhcMJRRxw/jzOa/UKzCb
N8KHveLfuUejqjJxEYOdM3v3mbLyLd99NMnLHaE1XP5eYzArdY/Iz6bZBkjiV6dY
R2wEK6sSyTwNo3DkPyprmIqozGPpBtmqubG1LD/eGgkoZ1tjznzX8Usz5rpiqMj5
k+utHfcTf2icSbjU4chzNxEQjLz/QD5P9sxiJhP4W9JWFD4chHn6C5fCg10yttmH
gbiIz9BM66utWWJx+FdbVeQpYSOzv9WCOvfB/nzSn31q6/hwkOqol1fbW2gEP447
OJIdytiALz1eiLzjIYFcSg8vF6mqlndaUDEDsxOEJfu4lMk/64YNK3HtI1oediQx
n+ls812abWIJPxIVd+0NJ1O1SJK4+SS8bSuGbR5qgIkc4uOiBuEuUCoe/qdh1gh5
t3xJfNgSYAjOh0PBQS97x4C6IP7OI2X9d0byvuLHxg0Tlzy3qKxE6BFXYTFDfrn3
xRw1FAH90Sw623cYNwEK78/dqijh6gWdfSVwaV2JTpOBXp4Mc/uQaW2tEBNVrTZg
1pd5zb6mZ1Ly1fOT4hQ7Iyxg6iTB7lWcKCrwz34RK6OVe/LhSumzU4v+Gwkb6ext
cB8A8C6DBTPUr8WbzzggwO7CxwXhrq2bJS7jBYHstr/yyyO7OLnUmg7oIhbImfZE
RsZ0T5VOObd7uELubdhzyvZYOiHBr3OLeYGCD/jo4ZvGEkX25kg2x9NusYTSAI9Y
yh/kbk0h+9NTH63goB38INwPSLYr0ma+PyLhasaSQuIce19CfExHUwopIvp+cQw/
HuIFWbORL09KzaTNA571jhVarKBYArKc2QYzaqebfydVw84u0rXz8x4Q1aRAxJNh
fWPXZsguTsSBQAKqIghvNssQzvC5SNoIIAS5AHjqPBymLr6wLRe4ajwqi8nzPRkj
6deio65W8JhgsNmmZyiT1g7ksjG3WOeJc2iHSdCoNgF3C/6Gmd05FtjsohTHa0tJ
lTWSR1OCWhNsatTWvLLxD5L0yxZP/0zySJ1dJKZcOzTP+ncTb6g1oS8GbS56Krv5
a5z7Dc76PDhrXk6LBki8R0Som0IkJ1rMj+tFhHGPGva12eiP8KeOP3U4Go+bp9zP
bFr04kS5K4DCLQ2HtEuZfRA6Q+0SYp8SNnUumb+Nmm+GFW3TOSkxs9RqfPet7Nm3
DAmxc6Z9gOPBH5CyGz+nxhQe4w1h2dX10Nqm/Njt6oGa/rEXBeOpDMnnF1CLFZXL
vYiC5W57p2gSLCJGU0ZBnWltyaPYbiF6tLClkxu2lD3CF/2YudUd1hsVwyG2qccj
gCPMC/SWPvoY7DSrXJ2MROq2ob/CzXdaV3PnUmxOaUmDprgq7kpO0B+IhIwlFtdy
5TgQ2807XRr/1kfFC2ie1FInqzbQIo6SYE9/C9ObQ5SRbNykT6yytPXRO4wAowGB
Amhd2o0khlQdgWnijfBAu5juq/CmBgdloQ30FYn82GQK3vW9ool0jXziHXOzqS/6
QCF7T5wvYVjHmoov8clMLI1w5Y1dvmLnGjGwAJP3GPpZYbsmSl0PiJCiXlMSlkap
+NavDXFAvVo4jR46x9OHIponVpnRs8mCE+FZGxVCLK6LFjVzUd/5jb2FGi486N2p
pxiGfYx72gVNNy7RWOYUb2t6pM3734C1mA/ejtczfeUYlBTQnWYMtjp+eTbCzyZs
wRtHq0Hz24jXJtdj7EfJEkxVUv3iL7kxKuHFFF59a3183ESlHiap8a3TqXAdvkSG
Jrz/Pqst5pbegu8eQuK/+bthtU/Ans5PJHPByCRUFOHOOfixZUsUAln4FTSYkxeT
bTJL/9g777uFV26RyW9XseYp5DCc4ZRVnsz5LRbNElQUDny+gevUou82La8KqLH4
fBgZbMR7JxkAtwzD0Bz8R2JAc+jXFkiyjq5/zvmPsRi9eyk+BmyptdxKQ0H1Sqg0
RBMUH1rsjrQHcE2RHf6V4iQe+MKQbARXPKC+t+yqw69uQuCQ75nmlHVyOSjPafJz
5TCyBoWmfbSilCUpCFjpXgT6RWPwkdC9UTKJ7wMAvU/7jIOw0K1JYDxGswr3r4qe
VvRcf8lJC/v5+oNL6VgzvT/yZkzkdtkHrCilqQ/Wi0qS7lLD8qURrGKPMax0oxMd
tk1jAewsWwXtGOAgIk0InVMOVCkjgjiTH8mY1KmLlg7PRwWVmat53WDhuiMO/uOb
sxAa42otxQLCvYfDkKLGza4RTTS0sqk8Rqdy6FOnDq/vYe3mpIviSKID5aQ6N4MP
qb3NwSCktvHGrgDHMQoin3gk39A3DTMnGhfeFk2IK/1kd2NJMm+NdA7W0BnL8dU4
gyCZNGizSeYlRSSKrax86qztHqV1HxzGADRqrrDpdZvdWRmMfLIzq4/EPGr6RmM1
l5aQlOpfVzSKv4Gg6zc1detkTI9RllVVDFKYFGzA8ao0zE4TjfzsY+qsspuzFMN2
/uwNBXKoIX1DxXVHC63Fos5BC0ZR6tZbIaiYrDdLVAnScfqJ3GyVJM3K83gSgGu4
vkwxjg7vX8Wv+3dyz1bHdp9mLNtj7rTCve5dFjhW/ArgyUixwL6nMXOoefE5mr14
mnwrfwn2UiaEH231orAKZNpMpM3kYOOjPzUNIy5TsYeCHK46vMzZYBfQsYz4N/gP
K48VV9+wTUfRQP5t1N37pJie6Ldc3ldv94B/y8+Ckt4vz1ytXq/+oaur43Y6uQLz
5DUy+wKRHJWGGBK5t9rz1TKFOsTbiXx/BgXDzvuR7sBPp0kIZKqdBNjifamrnoQG
LijIfDA48rcOODJoTNR5e6XIbA33MoUNmgJTYH6RudMkbHKhRiydM/lfBfemGaai
+AxW5nRjOZOhNeZUO6fMzupQLjM+4/zNvrp7jrbxNbK71JuxsnUWHahLvODiVxQl
D3ky7Mc19Y6xi/ld4LgLCNW7CY+ConMll3NazGrBzh4+u2NVCqi16RWFamB14db7
3pWkde6yOiqa23XzuHXAXEqRcPrc+a2zHIRx8PmPB3cLu/PZd5hwPiROZB6CY0zA
ILa63tio+s5BWSE3LcTzrHxW9uQOmETVF9vmeWuBBu72vDPKnR9fcNirPD+OScP8
alIz4HUjL8wKxgA6m4C3zEyQHqaSJs7EfZqiN/znPsQOpt2FSjYWPRWp5rph3+6X
libNd9CSzy56ktQMZWPWgiqjtUx9kAU/w7Hn0tu1pk1V5cm76xBqGraY4kcQo1RN
T5AAG8MqN5VBOoTc+TjuR9vtcyfu/4P85E+Ng4Hbz6DMdUwak/1MsK/RiOL5mDYV
WgQR1LCcydV5UeKa8VCK/j4bXv8kpjnZx/v2N7VLYDJZHGzs0m3chqXmiBsNOjmz
AG0R0yOxTBmwBwlMEXk3qCc6+R8V5rTHLIjVya58EQsBlAlX9r/spjGSqD8RE6tg
uBXG2TgYVekZWRBCpwLCmPztbFdXy/fDhR0Cu74WYQD8pHjPiR98oZKB0RDzT8xA
KIUyxOiIumL5Kx5tixbTKh8+vra4gfPBOsYCQCWe/22gEs5oH6oevbVenDCT/wfV
tH4L/25Dz04fmvGXb1t5INmCIIBrVFRj1LGtOqu/MgXOAj7EpcrJ7Ft6oSxbFfmC
3VeAV2licKJsSqIu3HhpT59cDMod+DbSBuxqvoAcRfhsyjX76iv/ELwl+b8XMR3a
Z9AHs6UkGH6V+9+oCPnVZMBI81cfvjI+mLEJflcIyazfCNYoni0gRJY6H/mj8Zgu
5c66dcvTGPpLj/i8Q1//YR62X5T7TgfQFHZE89dMPngg2sU7wKiYwY+/tzm89dFF
6Pfwq1yWjpxQMmYtFh/LMQz/lxxJsYeWA8meUYy359/KHQh6xDdEt9dfRqwE5QyU
F/q/aIWSdYKei4jq0lYKYh9Z7VAsksiqygApUQ7dtiQmt4ti5eZfZ/Y9pl5/wUni
KURwiMFy8PrpMFc2UQHkfAl26D9XUFmMWh8E7L7zd3XboMODhJB4Pm5q144ftsvS
VGARoIxp5XOXmaCapmrw0KTZihhtHoUGVkpoO6Fkmo19ze2sfzGOYkHkIn4IqN5L
C7lzKWJHUjGEiQ9WeycEv8k34GjCE+bs3fxxkNx9J1mxvnMXade98COfP84A7f4i
l4c5Ac/i/VTmI95Sz8/acQOTTH66YDal5/dlAC6sQ+YnJb2cghfOYnISrjKOEYn+
HWOfK7WaakV9EkGtnWyKD3SZT7c0TqyiyBtL6HtqBots1NCuXZRLafp5am6iqmW0
n/VC5Ot8tHoIXj/yFyEwm7yZloabj/uy2wXcDWNq7eFuKL1NeqVCQr0UOdngzLnR
RLLH3rJG5WthsqdriSV/oX3Pe2K71OQRh3D0mbOyjnBcWUFnO7u8TiyQISI56tZn
NDOlVeobfSsNWBl7sI5zDnBBatdfpapfyBhAtlcU7VpICMs4V0vNWaBRNF2UDeY4
/1TaNbLXv1r2xl2x0VfncW+/5O/05RtDhiIG4gKj6VV5+aKwUVKokDda5XIe5eWK
zQPozcC9MbaWmagxWZBYDwecvrggJz2JDVoNI4BTxKZf6CKsRrSlcjW0aFjL3j+L
JHI7EcPBhGaqujOF0h7bshAkhd7RIEBo2Jk4jE5sWTyZYXoT7VLbmsGJcKKxSj0X
nZUe1AuEqB25hz3kchzuZFEoRsX8jeHjJvK7sYo/xDdp7k361A59fa4OHjk7dnOl
7PYGl1CDRQ3ae2dZtg9Sa97dZ8OS4oYjN1CVjj00YheHTz+0bXvvOIElX4J9h7m7
VKJTvffVRREhs76dd0EY09W66t5J18q6YHqHmJ/vTi3wh5DpyREcaxr3bLG3ilUh
YwDjKpe5YY3auybR9EwTp9KzZ/Ltahlql+2u5SgJ/wStCEnXQ6Gr0Dd0x84H4bL7
`pragma protect end_protected
