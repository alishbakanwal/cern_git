// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 13:57:49 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
nCr+sBSQ4BqjO5lqPwT82ybQO/u8IbVD48mUqvDJuT1w6P5x6j4kcGYZcnmclHVv
z0A80pI7/M8JF+7mOhU612blq5g6Eta2cAWVL7D0W6sBw6MVV5qA/yh7q0G5ReQG
Fy9Wpt8xn8kzBHvluCf1Va0HLYLamGRrXO0Vbyd/MtU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 10272)
KE9N6EfEuLSwO4hZNDMcyOo8oxQGpWRW+kb6BhNJrXJfyFJQTt+LYtXbG2MZIKlG
2UD8pfLUIkxhQWwj0utp8uqKqiSsYbrjS+faDP86NWgv8FYoHx5YNQq3lkkpiSrm
aKMc5+WzRoVvfrrRSwxHWnFKn9MnmmK1NN0Hc3A4P8WV5yUASXzY9PKwOExYtrKf
Ds4tz/7VmCsUd/P0xCB6K1u6Lr6BRqRZXY+8SwPLIm518oTX1uN3ZonxDhvO/l1A
otMdOYteGsDUf0HSDNNJcPgQg1zdYBQNgF6FAgfmVILcXUMdUw0Wpr0AvU+5F5dZ
FLSRp1S2buFDVZtR3stfmcIFPVKb46y2fR1rkl68Hg1UAVUwkAnKedg5zka0d/9s
Q4ddcYsZkiCEiARcQkQ5yEHzQyFh7HHH4ujv7rYJ8GJpIPiMwAX2gIF8azTC3COg
8Y7ASTRS4YfLO3YYfqH45dRhBt8hY7jIYMRqkVI0pxZ2jz2P7/YYqk0EBPDrAsDU
CmorYYgFTpyZG1fNQSdChCyLwtr/kQuO1B6WCQHctZ5KW7DQUQ+U16WgdBOmV6Ea
0VF1sguUNh/KRFSHq02sgYz9Zs5vHrG5TmNCW3TDsruDSbNyC7cpum0slKF0luw/
6len6b0O/Knf7bN4vy0FODnU7eWe9NXX1K/saBNh3A1Et1VaqrbWgWbPu6LbqHDU
pVdIpb3bzRn2OAIMo0fah3SXPjA1oqLfX3jlyIHpOTn4UmE74ddEWbv7woh5tV/F
mdmuj1sNiZlUrLD/8iHXbkJu3nepzihaJrkX7Pyr2pQGVSlkyXpcGHm1Gf2J1zV7
sYkfP49vpCZ7c2uFEnELumqtqGh9A9EaXAcbRPbE9btC5IqW2YbRuAcp27Nnt5xS
q4CBTm2o4mrlKqkGHrdP1AfDXcZXgNjuFDwFOp5/cZ8I/+zFK3lLkY2rmncGrE6D
+9jWK/fz0dFmQMArSWDv713PHZRV691pdnCy1jgD3TDapn/mzpaDZiy6XUTg1vWg
W0OlRvDr4UiYksK2skLvRj17scGbuRGbbzvE1veS3CH9khOavh4zCqrtyW+CqyiL
39DqZWpozEm0mkp7KFZAErU7TN3lev6oJ4o706bEPtq9NOBsgwr4dg083TGH3Tz+
nR1an980lAanYRAIsgQquYFWo3qAVcinPIirBs28vIY4gDOtLlrHbckJtyO0WipT
PnEVyAk3qtaFQ8qMUfJyqzzAFJ2vxLOuc9s/36w3nbBM/pGW+oyjtCqPhLEfGarJ
qOYjTu0vXr8jdZHzl2CB9jKfmnpcG9SvIrtrebEbkcRphhyO77zvxzw8HiAbTBGl
z8oBwzI27HOuV/b8QlTprlcsi2Gzba9pyP/bFgal6baeHfCTITjSB5jPHELhGuZq
C0he6KLFvgyn6Ef8f1aVkG4npHhClLt+12c354IlswSYvZw6A9+nhj9jRhca/EbM
wFA+W1s/owwWposQ64IbawMdzeoYnidlK3KZj5rBiEZgTdVOyA4LOX/hA2I2KMIe
SN01lfXkWxDjXEAZKf5qrCGJSzgopZ002jRXyRI9/aBDgujY0YwVD3ev53hIJtDt
hovPytFPd4Hvd/53Icz6DISRvOg0sn/K4hk5qttMBePKy/b4daud18uHz/u6Pk/f
L1vt94EQGPx8whco23mtrMvO4ESKiApao1dSFd2vQcONwLO/e9gU9Pp6rbpucz+8
QrisgSqPiCvwpWH9vTFSSt4d1GtoTAl6LpUkC/g1v/vAzWT0z7nnFuexAUaiYmud
YPtV7Uz8YPLLrDbmLMQeUe3iqkkhQINTgDL6moqNC06k5IHR5i8w4pNyRmf20GRn
Ngoihu0J4mDrGT82wr4/tVZ3yE4vFaqsKWv5vwEOnArVIKo67JGAt3/0lax7mfre
IJmSBs0sz83oTki3ObU1GMTBZ4tKjzLMlsAkvVqZ1zhPPt2J4rjaRroVx/zpBCet
uVd8giIUUzc+cV1eny3Il73kD/s6oOkCQFTWBuR8/olI35T/5JG/GnTQvyZHNWl0
DfBPiP9cBTQ0nwJuasWzcK49HAaS4JK+AfbCJ7nFmeCUaqAtIxARo6uiHgQmeDOX
K8gnOmmaQswKshBOkRCEAOq8el8ikB+M+4WZY6MpnhlrAGuYrYeyzetV5UARIpn/
LdwP9V82wp1nhuK5rs2TTwZSJo9v8B0Tb/HGBYM/wSLyK3A+h+FSHJw2vxvQpado
3ZkVdcohIOcG2Qzlw0PablO0BLWJjzSlfA2k+7RZY/hhD8Bwq+3VcPIUNoQWHO6N
lqzIF31Q+vt/Vp7N3+FOENhFngJ1+0uuA3IsewFqIwhw8E+AyuvcA5LLhnEpqdeX
XDQnOMvE02v1OhsRlQbVL2aCza7AoRCYmEWQEmxTNEi705BM+WOwMZRY9w75FuwN
dm6eun6LzSXkEnA7lmOz1cAtoGK/weCfVJoG9cjr+AaDzl1BvBqxa34Tk4uLaD/O
iWY1gyE4lnFEbL03QrqhF6XTQ9uOwxepislnUh/ucNWJdmP/9ANBocbv6rnBxWuv
89gKCwlQDBDTqmi2l//lbs1SXACQ59xAr21K4iSUSvfbLbg5ef5PAiIH8sgZpmho
Jyl0oDEGvD4WPhxK07q9jgbgIoOP4829R2bJPdixp5hc7t+qHXFj8OZOxaQ7ptWf
i1956k5/CejQHFXyrR0xZeAH3wrq1UPd/tfvxinwevmGPxkWRkXvx+byBXTUD+VX
YF3a6qR4uNOUzcCoCMW8UNAsmCMdA79lKLENUceuXlp9P/S+cKE1J/TcE3r2+y3v
UC0kB7yEvD15+bY2ddJYk/TN13VzgUU5pKlwjZo43DqglyiBXs9U36PFm3dX44FP
+KrP5lQJMGePSc3tVUgK4V1to6lSkctGaEG9qE3DI0qXqEpLUMWdEWM9KgCJGwAN
zVXUq4b1DE5Qv4xABy764yxIXAUkQ16leijYhk1qWkXI+6W3gYz39tRUyw3Opgf3
otOmUShTQA8Z2k4oHxS1XH0fNd8SLQyoCvOY3bib7H/YT10N9ShfNquehV1XczOh
hwqSrpta6b3x5+Op4eZx1hHwG6/ldal+UbPcFANn0gI2S3E0B15bRbKSFrTK+EjX
4Uzf4tkrdIouTq14ANpPnm5atIxHgLcx6ZAqdi4dvkBeuaS04vPcTY1lyjM15+Gn
2ar45OZbu83IZW04OQMJAzrYwm1lH4HYAtKOopo064P0X+pSTE8UUFCJtREqkBoK
oqC1KTXpGPdZVWt0V9bGNoLarQ1j0Qdzep4bvQTS6HS//FMAQXmNM6fqUXAFE+db
Gt43Evk+q9bjcufZJhBDDIInIM4zfJJi5rvw46WmcdCeiWll0YMl9cWxGSSTeeMC
b0cja8sRpd4QIz5LWlgPBar5svfBNnF6YEGJVsko/AsQl32qTT+pFXBVmcUig+Xk
qxZ73DRJt6qCeg4v/X9J1QRETqAKSkX4HvT7cF+P/Kye4L8SOC5D6lCBL7qF8Y9X
pa08htJwo3PNNSZPxZB0TNc6jDszaB7XtNJ3WlHGD7DItFTwr1B68MaMWtkBITZT
AZoIe8zMj8fkReaTW6QEKCh+ryKaWuFFytoqNjpaHLxjIt1d2OUPHbX5Zw1TUsGA
GUdUwt0fLaxkXagA81zAf8Q/zAtditZNP+ts8Hq8RAqFhuMInijPTzU2+CHzs8yc
vC14lU4EeJ9QnMWPeUCeF/DAf/HCMvJr6zY0XyhPIg5tiI9sB/dZ65dxIqJzDU69
rNiD6mbYKtDJn4HJfK66+xI5ZxMLToje3axbPOBYJXUb5DdZZQrVqRY7uvy5YcCi
TAjrVguW/H6Ygb+j8GbSn/rZjFafmQILJ7wSIvWjpLsSOAYS0F2w4i8ODAmk2ZR6
RjziIzRuxNPfIw0hBwnu3ZSnJQF3tXWXz1qO7Sy4owsYyFI/RlS5v96CEw3tZVkt
0E4hrU9jMxNo78U7+mrY3juREo+EWQ+Z86vBAWliaO2lpcRwnj2udzOh1JrPnt1O
mEvXN7jDeKRByK7RwNV0Kv83UAr9gFVC8lNN2yFkLxnushfRxdBmrypTspp+Fb5O
5uRpb8+/8ANP650CQwk6FV/RsfBT3XEDvltcDjorjkAUbfMzts6WiIbbIi8xDIj/
5DpXodrLvNUdHpEMsXjUPVPLISe9xFkOUWnV9ogDd7WRDfPA1MpbfroOLrv4wSWp
MDDuiCCCVtrQrw0WcGMbjYE1zyjddAg3ee7+2DjcYx0ttDtUljLSpD3FPdQBGnME
oXVkuasVrkT/8H84ufK4I/BNbOOpvf9Q58uqwC6Qhw7ONpgYD/ouHo0NqGc0JXSI
mnqPckwHPug2b+ifjuBiinLnT39rd8fsG6aSwxDVGt6nczn1OwZjkZUjzGYRGa8i
ERFRB2BXjRLoKt5/aZFR6r/Yn3VgZs4NKsFUSAY25RCrSVGuYU6Tg+ekz7yGIEIf
45HUJtLef32XrhFqN3F0aWJS9GJdMwNPPlypQw+Zz9uGJhhjcdGJOpXgs/Et3ymU
Z+eF6FsNZ3/xaMgejA/woOrVIEtRcJ5BFiHBzEVf9QsY4+Jzw8DzoYZQfoJ3hqy1
IhdnRNChALcxyhOhxeCbsw1UpFLlSwQUs1Z1GJY0OQkw22rSZaNY2N+nWpMco//O
PsU+XdhvOBjplWtdfuzIJh3Z41R7HEGT+s+0t67D2+EdaNofsNbvWPX6zjeSO7EF
Pc52SF5CrEUq3QyaDxzpsN+i1qAto9DBVKLb75EvHZa3RtKHTG1VRUCl8f+vdh8r
0HY1VA9mdpZcVaXjrAiealMKYB6g9g7mzgI0kaFIUSKvlbuyg6JopYALd3b22DKs
HZmnAd4PEinf9v137LAirjKYhCXrt8NemiaYf789e25pOMyH1n/WsDfOwjLzTvvP
GApFvWxhPLZDC/NgCviqzXkWqxBz1ZG700PVJIaMjFBJCd1gJZSJLsrqhTz0GeDE
YB6j/SvDvUslVPn9L4JBdin3+UBH08XiWJq4x67QPMXMkDhEhiZ+e305Z3lTJnzA
poROHCZ/R7thOyE5jM4ZBSgMY4DJqUdJryPrA96k5nwLW1IToCuOngy94vm7C9Ly
ptehM8TNkmzukyMF3o2hYSGhYf/nGqDwJNWGtq4JXqhZo+JRP+r1djLoka2OHku0
Bj1nonzNFqGLTK4N4MgBXCWvc685xxBpFdk41vrijuvPx4HD0TESFnC8tf/7N2jv
/JUjnUx50TfPF+qvFvaMEXUtJWkVpwp2G9po2yXVHw/ndIm4z773w3wXFYUtta4+
WmLVGSnXjxxIKLadkOMCDDGTM1r4yDhp23c43I95i5Az9uvjUhnIT6d/TFw/45Ql
D/PzWygNM97qG6DgD7pSyITOmH/iLgwo7FDTF0l6uGolLc/EZ4rEddHa5JF//zfn
KHGL8L3FsXWi6R+tQ9Pf5oCVGDSNBListV8QkTHDniAndlpM5kiMlme/U+LVzFDe
tjO/wZW0zOwEOQ6+pfELJ/xt27y7w7a6SaGq9jvtbdHMwSHbuK5Q3WRWbyjIhgYV
9Pw7MWEJlcTFAzs6ho5UB/fACpydNgY3Hz0Blj6z/u16GkhiQ7Kw4Az/zLXEUY5L
wGnxFd3Brt5gGcoaybbCx73XMMlP4c54RtTr+FlIKICK/9+yqIDZlMh6yqFFgnyQ
JPVh/Nnl5gOwyO3RPA7WKyuzMWtzhLn32Kz0Fiu7fLAa9J1hKI+OnWzIL9Aj67c1
rPiHur8pBcERZNgb4g3CiHanQXP7uJN2oI0X14vt9q49VPBb50zr2I4NqZKn5v6W
ct6i0C+bKiyU/TG5Wu6qS5ZLDEmvHagxifAQ9VnAPt7lYbnEHYoE6YDQ5+w7gb2X
y4Ok+MA1VWtg+lVq6Wfie05uyCapMEhJdvCSq3EOyzypFGTB+jLNPJaAfPOgVlhv
lF8XMW/erxyW6pkBAN5S8hfx54HHEgO/tB3nzJKH63o2F85dC50N+7K9k7FvClnD
97FiEislPlKAFcWo6odrlVGsY4LczdJEjd31DoZIltx5J0NmyEZyP5cvLTuStYLo
5qZfoVC+vk2vmnzzXxuTSH63sKrsaov4BTHG+cXLdH6O7BPsOLJ3uE+d/iJlr0mv
RFG3sgfZ5Mw8lagCgGkQhB7dCyZcz1bSLTqutZ3eG2AzRfr/tyObeIXbDPXn6LDB
3oXZ0Eny+IriVv3rYmIYVEO89wSTSbx9kMYfHhsS4AtSgiAkgg/C7Hwq1b3xAwig
KVIk7CsHcy6KpYgH4+UQlD2vAg+Xz4QHahfM5e5iyOlLGZ+qujd6cetpQLq0GFMu
Ml6FCj/2JWPL7vVqiqDrs7QO2G7kABiRj1eiLdGP+jD1cDm/Kz7UCoIH6YUse65m
9Yh+3D1HY+bC2lE7forrNzXPa996xxTZ6Jglzvi9cRVxw9Zuj2lwFv5KWmm/TK+z
WPMHI2Uz7a7BVIRpUW0NJPeJbA9SUs0jSdV6t82H17JiPFgOWbNL/X0CCJxzfnSA
u4fYEG3Ay+rF0ceu3HBIVZ8Gexmg295sHzVN7RcjSstLFDyBJqEkGfP5yzDFn9TY
3YKMxoVVj4peAJm7NR6Hq4+nXxrWgdKC0FMeR2w4kgTCXeR1qHvhi5xDCBsNb6xu
OvVK3y5a3UeQ/IIXlkKEi839ujna8bUk0yruPig5aUWO/nABR62KgBcT/R6IIFs6
A2m+/RYuMZuVvwt5DtpwO7bIcdSoAK3HPlTe0r5p7wYYUggqxP7WXe/rTcU0awo7
BgMoeHLiHzIcSdSHp6//Z4CTmv1bijQ+2fycj2FosBhkdeQhOFZGh910QVkHI+YF
BRvbUBiGhlOiuY3tIX/69eMB7xDzgpthkhvDmML28hvoSyGoL42iPnPVpcFRg0qs
vGPGquS3RkfmD6T3UqVDNBkhPZk9gr4gindzQxuEYplc43AU5HZm8Tit7A99VY7k
ISlXQMZmvb8H0fSWeB/7x1U79QeBe6iyIOinCN4WlxB5+02IGNN2gZqVGZiJxhfU
BeVrErk+4CMeFksJWAXlQ6txQkL+/TXBmeegID01Zv4HSTdwFr5liKtXYG88RtmO
OS+Lf3CM8l2vWVZfQN1ug6NnGupEhpballZSQBXFlbgksUJY2EAq9uJtfqoi2dmH
GvvBLBncUapFd1BBQVTBe7gvYTT4dKX9z2p1B2nKdrSdLrURgHQkclT3dWmCPM3J
I0zfM59AtAneeK0tkMO0CibxaundDtdcxFSvKN0g8VFaFzl6s6SZxQU1poRNYhmT
a7gqlIIpDHIbIp9hqOU1tL75ghSdnJpL+YnCTm4qo9WQN7a7rojZBVgOiPYjNpd3
sI0zKQl1WqBCMbeNKVLLLvhCMEmUWbbaaF6TOsvA2yBiIJr1t+mTBeM5Zzo0CcTw
gYV3+eiTp4Cp0uUdLOHiCrjxNhSR3kRMGu8hLC8OVWKKtSDiNQsGdNN0WJIfbKJG
N+p6Do87SIBCsj7u+KJoob4sMHgBeJoytm33NlBTz5mx0lKcmDCSQ1gx6u4JeeCK
N+s24cugVNhO7FUiMv4Ocuig6oALZL4yaV1SrEgcKWgC9944j2mruY4sbaCKBhcV
GoK5shyg4xiJuaEiga/riZGR6dy6Yd3gCeljjO5OvwPN+2JBYaxaf8eIG/G31ZXr
jNqa9LiSVumLcLmCheJ+sWI9uvDWoO0KhPI1tjbc1mHDa/1zKdJfS8V3diNLRo6+
IAXh5YEZd+vpj4GOef9yIRC+hL9XqP9bpqBmAvkUcthQ4XbAKzh6ajXO35wxZcHW
xxj+5tJ/g6sZ9EKQ+Ks3WRPnKWGbph3TFaP//uENiKeM4pxhnV2iID2dcCIULQF9
b35X+tTO+OvUu/Fx9Fm2TVeseCH7O5rTTy7OwoJCn+V48jyHa0haA4bLoPW+qX8n
VwFMseEl2jPwqo12jiDMP5KInrH9U3CTBp55XrQBHRAdI+Dd9nNHYHvtfOZrkocG
9qPAAk1Fs9pjLhOzdBXTceS/924Quj4uUxHxFAHAwcGePj1Gkmje9xDciG3rSmtT
4Ujteefr933SufBN0rwlMi4x2e9JZQsZCcbv3NDAX2GjHNG/0nq6AqgpUsoKFZVa
zpX+rLtswzZ16rU/dnPQHee0pN4uASJSbcHT9lTDeP4f8nfLIIukaE+440oJYS2c
6Og/EJHDjNgUk0Xz/awz7LVbNcrWgGC7c8rG9kWXII+4JZ64SEWraMBPN6DKVO42
JQDSpguUYZ8x1XauIp965kuFLcx/OPU40MLIINWVs+R7B+6HnPpCMMiZKsI3ksRH
odRRae3XjpuSxZg5rrKaYbsLYE7/8HbsPCCRy256Ls0LCXhGJ1EExEkVW8NV1xB0
Xbj9DsWHYi3L8ut2gjwiiIL5WOa8clIGIRkP6eWc0HbswG2TXOBldIMV2APQCXUl
czv6nERAi1MlItxKVryBpXn4IZS8dJFLW/p51/+QFuCDj2u9ggTviBEnui8WzetW
AbRZqJfPViGFK+DFc+/+jmqhiukWedw1kxDfHL/T+BOtZvTLoGkMuu2TTT1aDl2L
bfB6mpzYdY8GLO6dtDf5/q6B16+pF8SZKXr9a1dotX2VkHmHeiyyNIDfHMfgsdZw
KQmZUdJHy+xdIx+rNsEANfj1aygNrjyFgnCSZ0hMxHPppXLy/nyw7fYJTcOsA3/K
kO5JJ/HobgIv4ynH7TDctjkq/p37iDzA7s+/BT0gZdVTp5iVE2okcdRTp1F9KdrI
+fReQz4EvmG5XujZCnVRwjJPRvhQIWm7pWh8JmWvr7TvmDqDyw7DVAXcKc2TYZyJ
SD+gJAXFRCsKXDUL27LhniEauopoQIKnBpbjoAl0w3jzQzXiIdQwjfZVcUban5VJ
zgZEm1MpyTAv6veuEu9f90HxcYVekx53IcTyLkGh0sQUIwRn5UrsJevyn8JdFiHw
SRGOMl2d4/UFr5Ez1hxz9KB3Lmyvpz9f5v8RmNDt4I/WSHWUMbjr+raDYB/IPd50
69K3LptSCNCO0FyJXsSUrzWa62E/r3l2NTF6VXGuC/cBkDc3JVLpVzOoFDsuGOt/
r64vTef3EkRL/1bFLcYuwERlLzrkVKm+LhCJl2INSpdXFRCGdljSBLVBkCYxCdNn
sdYmUV+hZvAboCI2B80JtFiUcjG3yqco2muQVsWm/RA9kYD9ZquRLNHw/4pGMWDn
hSBuA/Xr8pOpcN7JvN4o0l7BTDsjAsEc5+j1pKXcZNzdnGGnVyjDJ5ciFwxSGlzW
ZLK/6ruBYZyF19CtE05zrHkJ9VRNsI6qtngZg/bRvj4WTpVKFAxOOvBDYmWNukqR
bNh3lFmXkqSnEvLbx1C2On7ebZUIZDqJGSJ6Yl4eAtwUvrMILSA4hhbTovgqHvu4
VqkGDWaDrCIUdJwv58bbQEE9ZnAi17WCGN/hlveGFS1lfFeuKY1XxZbuvl0y8nh/
8EUmBFbzVBKa2YcBZ9LL+FyRI1mW9mKnDkQcpoh/1uoracOR9IevfWV3UhIWBvI/
fZ6CEKNImgcRYtvrQBuc+3ynAUyXTvW4K3qqD8MFMQvvvxWHxtEqOLMP4OCT135E
hNaVxhXkFBvNQc64/fInle1Sp48hKokRiDIZoBZo9TV4/FOkwLkV4dwcaH1+vwxW
8DAr3WHformek+42W6LzEDztrIYKM6jqVl7VM0Se73aPv0yvDPZ6MGOdz6O0Y7GT
LfOrreGe2xmfrU1gNXAdNA/CPtoX+4PA5ITiHGZPnWiiJBtg0z1K7VVvVdGokvFP
Q/LFC8sck2WNyX9o4KFukGSswWDfm4b1d//ojP2QUEYECJDkZ9lIgRJmkM73bQmP
Sfxcu6guILkIL2oJ3bPimxRuDfAaKhMiSyXj9pd3IxqLJjQzesOwz27NCXFaLxkF
XhSdDk90hEc775pPy9Dif3v5y2N8AxPBjo/jWMGzvlgVCnoJoDaZb3zDWXZmlmcG
3MxfQZy76+YWbkL8WiqN/cdzDmQnPtkej1KnMWuJoF69tSAc8lPN420x7RLaOZOl
/mGMo7dboyJvky2HN9akX5OJ4D5XM8r1w3sam/gKuxtpm0lGaveeTlzziqeaqaXQ
VNigXkowRh1ssVnwLbm20EcuSZ0xkr4ewk2DdZp3s6GVpAxZ+oc72NTKw2ALE1YC
J5PHTsri0T8OqLy+CB+2iLKBKN5IkcMYp4dhk6fe8+NH041r+l57rBK9gjt2lrVr
iYCniASVc8/jnNtAkJSC7EnjKsBzDabeV9afVZ3p+ssZ/Y0CbKUC/jcJ9x7UAOm7
I4WrgLMbrbEnfPzkVj3NFauviY4pD2Z56sk/YfwmQP8MQLkJhoaSO0HLcg5atWeS
tJx2ECn51DpXXLxTaMIuIdOyRfUcmPei4tuM7rkaVdGACWs7n7G0nqv649WYdHTp
tsAh/qC/fSFIzaMGysP2PHI9vwRuNKyn5WUmMOH1uhWgaTR705qvfEPmTZ5cp3gw
WWe3INTBnLpdAr+XQdsq6q+80+3EQW0Gs9/AyKJr+7/cXGtLot2fE8xEZcFaHWh+
Omr2GQzAg1WI85E6EvF7n5YXqIYuBDd8R3BJZ1rUcnMKFr6MkUVZl6gDiWpwSiz3
Eprs2t7be0uITvbwlyTc8E35jFL+O3iVzQ3Fq7D3FPnLRY4sPAjeJrJTIsSASJd1
qrHZBHaVgrjMKjSZsGHI3ZpFuN0sCdcbg1tJx5mzXvU2/n6CCVc4Ik3vBB6CtrZE
wsScMoPCLyraOfTrKKguitbxaBRB7wIcBqWoTOUJ4E+dGHi7hRYi01LyrQnoDiV1
dFXxP3i7fW4GcTsscYKDSgy07epr6NN9wr3BpWLCVT07ytHVwKMqcwEW3clueBEz
WvZhyGQhVwb9/yVA/vMeJ445HKBIaQlmN+XXndjKNOKTu/vcz5iZbD+JspGM4aSh
IOiqjFIqXDK7HoLg699swOFDUWeLKNEHz1+8m8kQDoi6Iry77PqV8BDa5uNQ/xRV
pFzk/4WpZg1ebcC+V2HaFEfBPv2aphatcvc68npIAHhiXdcUX8jgqyPBfylnuT9Q
wLvdhpj3wxxzKknQPGjVbXfot0Xwe+WBM6KspXD7Odl9Lm9Su3ZFTjn8ZwfAP00o
0wZl4B7teOmQ3whTUWQ4hqQeeuUUOXUKsN9OfYsHzAQeKisMD7d2cXDC//iPbNGn
YsSD1wFRE2IlHFozDWT9APBrDqN/niDvXUFxQWxs9xTg8FAQFS4CciuA2vXoDr1i
VsNasBAB7owGL4XBGx5tUrd8EBukmqCshEuSke5fbfFTxzhiHVGQuOjg3dnvDR5l
UUpsvaXYt3p3Zuu95KZpyXQ4jdMVkSzhNmZLkQLs7cZvjCTUFfWNq/CUMncEhqpk
JoVqBDJl9tnpUxYS4W8sPuidvJVJIyaGfcYqk0uURktXTEstnKb/wn+ZNzCjb74W
dF+cftGM3wrWx/J0HMlJ1VhpkA67W70YQg85888wIzMb3AqFpH9NoghJC+h6jBk3
iAQXM1Uwy7xWd4j2buj43q5oTk/GA+cTwLzBbQXHp4ZOuHGeBiwtgwCv+jPaWP3v
F19LHbzzVio6KWbCYJEigM0lfdqyL5zv+w0YKkWhexVzwzgUMHhM/rcU17UOwrkd
lRCwJVbWuYUyPTTxucme9wVHMNWRic6LP6ibTWhiLhcq5cZxL6aKSMkf0JmYRCx9
FcxUpHivgIz9jd3NIc5CWFjbwQjpZVzLkrdSAhXKhNVLjL/RK5mqCNzLWitjWyWv
rE7sY+G4Izvo68lcEn6kKldYcW6dEtAiCuQlFU9+wFW/QBJ0AL2ZynTEDk1hMnqK
R5g/43NQz04x4JytH0roUTj2oLJLvhvHfXDmJyvhYtqyr9J61Ng34Cs2u12UIoFZ
OxcTz8mVsSrNcZda/t79Z4j7jdQovxcGrK5TIw98+2Je6BCgIMT3ZN7IKt2i7jPS
Wg5aoCVTtPlPKyAARhYacgc0EbBbhs0zPNbe06RJN8FgdxUDsDkeExmZtIHWYyW0
wmj5x9MbcLOxYV5Byi8RWNVh1OCGi69Vv7+ZxnS1qpK3JZs8eSqVLBMP3bEbvpkn
naeQmS5V0jLTn+gFz1oONeRQAbAYF8gUljq3Cl3nM2rVe9kwGBYbhfJI8MSjUreh
+VCkBlecYJXiu9UbV9iZBpEjvIzTwk12l5Eh5pSJsrNfIzIAn1VvDa1bbhnzgxs9
6FKrPERV0e7+zRSYN9URysXvaXW9Vn4H+bWC/f9cXLWZpUhsQcbO5TYJpbUwduNs
X8JA1hChAG30AsO+1lRIQzB0sE7ko0AwEpTG61Ov/L58WjKxe9bTlkJeIf4HDJ2G
vyKNBrtBIV585ndHWil4DzX9pE2q2X2poF/J8xP45S2NF6/vcEpbkzo+2uiYSHy/
COd6UaJVH0Gq32/UUTx8KFhUyVXIK5kBvQDz9umNZsMa0lt0TZ7MEqIBmPRGUbIA
JxdVI2UyAuo6Yruk+9iUu00evZ2bo5SKrSnX2ezr+3iKOexofREN97gSutU55dfR
eHfFwd6YYM6ZcyYkUnbsiKk2zWYYuHr3ihsO7BIsNNqyQMvRfcZvAarTtjWIsA2D
s48Kh4nCxrUPPNUnN7D1P377h7EUYJv6d7od6NUXiQ7vvKHVOv4ZSB/FC8WmnJ/K
EIp62HKTWtEdDE80WrI2lSKzChZoXXC0c39okIdtizPYP11pMBgGUKxuFWqJ73nQ
dUha6o8xOeLs5mQxTyYs3eWQps8wkiZnpMwUshwDYuvovIIN+hGxk+2VQtBTFiX0
vK4CaOTMoXgkGvihd0eMrWTWmSlMBQmXsO3igVbDK3xLrxm+8Ku9at2ZppWu9uTS
ArWfnhbgZcRruhoeB+TUm0kmFGPYnU9OOGI0ULTY5WnobO9rONTVe0WqsypQNAJU
I79jKaOfrPpF0wGv/D/Mo6JZS1z6c+mQk4FJE78ar4sY/u0IF2xpA69xTG7YJ2J0
TrigpDQIVtpWGBJ0KUv8FIZiC2Kq6e54MMJ9+0Jw2TyV/NOyu1jvISALbKRL0NTW
OPvzQd/npMNfYt03AJsEsv0IoUBE76bIMaFdT+CqcAFqC7wh02XKTlMy3JcmLrYk
usp1xxZhVe+AY0CTN2OFgtZ8u20wq09JFHzvAOqWc5oG9a3edfs2LJdQnQLR5/ZN
BPPaplOp5Z3zbDUzpirUfTu3hkq08wfkFjZpF7vdHNDzUyr7eyb0BvgBqn+LmebJ
vmtMHXAGRDWW2zd/nkq+YjbTjYh1ilByClzBi+QJeocLyDBKJZheEeh4VOhCU4ym
KWlz6rVum3DXtdqgwjf2jYG/4yVOiJyCFWwT73TgdV5kez2A+yJMQl2h07YVzmvZ
V3a9iUDts0yZYBSUp2CnZIIKhNKvgJiPpKv6QKM4rR36I5Z2kYhw3Q9RfMZiuQ9u
kZFXL4o52EppuzO003mrP/tERBcYd9gZh/s80OkjI20ZTGdtZnW0KikhGysLKSoJ
4q2/EF4K7+Wbxo7j8ipjGgZUfhWR470oBAKO6LO2DSmAt58V46Th5ETSBxd7ufvo
IV4VeGoEWs1RmbpCe/IDF6I48uB4Uvnp4CqK/+W9ubXVJ2GIQcD3VQCih5UB0NAD
gipYn1yzpzEN0P7Avm46Pk+OpMelxbpbEHDEBpZTm/yB+GjXkmXGRUAd0sEGFN4S
`pragma protect end_protected
