// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 13:57:53 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
U85v9gsDtJ31/Oj5J90+u6ERKlFV5RpMmXNisq9cYjXzWK8aUizCeWn02uqRfpc7
V7IoYkNfC90iYmWzctLtvc867MCU26htWv0aVPDVJGuRQ0sra0EWA3aSSjtsB12s
aOU5fd9g83YzQzK10fRRQKLyO5S1adeCWaMKdxp5yoc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5424)
NgjmXtbgjqCM/jDpSx8gkmRhbkPWegO5UP/uInW77xGqlAt0V1AUtylreJOUP/GV
7etwy14yg4lwXIGTDSxowmm9AwiAQyKiJd0+ZLiakrwQWBbMcFc9IkQw3gsFIVsa
NzK+p/7VO/G6aNEboWyIP7XYga/bumBDFlttfNKvxN8x10MAQkyLEpdlkTo4L+ps
1mogJhoNUhzlSSXpZyBf42locbsQG4e0/TwU/QgLWGeI1YoRI7RGWYrzHIZZ/0s/
S4idXCGCRb2ogpwE488+vv1WGT96C2Z4nvKuf3sDODKRE1gDFSDqzBuQ9ydyl8sd
7YyiGockqJFRjPePCJaLSK3atFw8hI0qEK55YBLwMPZ5zSuMW/swJIcdOtPUB6zV
rWN6/aF/i71WiC6DR9zlNuU8YLb8YYroZCPUwmx3BFustMz+D34dBcr/xS7z7CB6
3JD1TBQbaMOTzwvQecvVHwiRU1k8zQU3eDc4tpmu10U7vcpUp06+al1xLRe2Uwg0
aaqBzL/3UhlI9xeePmYh/fxpXSnEKfKEjHIG7ZXcMISclenamnB0K9Vjr8wan2m7
mdSRiBOvutVKDNdWEa0uSSzuODmMBGTwuk/H2PEV3zqC5JiROSVZwSSjgJ9y3GC4
CdRtmxmTc8nxpH4MNXqVc3cQh33MMY9vIYjCvfezmoqvDv62mhOTxgGsgBY5LqD4
CV+LPlVrugcqkw5lqR91D/P2lEei09fUO9+BkLZWOWpYvtm2zM2J3pykUt+ynyfg
MaXy9/7TGSZO2cQ2EeEkQwLwgKSE1RfLb8OhQb1LlUF0z/lH46qocdfYsL35mAYJ
vkzgbUincS4LW2wM8lMcsxkSNBq5MFN/kFKgN04ma1hy4c546NzPgp2ZEfzOWVyp
+we/UUK/Z1QRRoCNUx+9lkERQihbS6xhp090sd8d3Nal12ZRu7KPE8nF44XCtAbV
k8vZABH/vHUwWovTTqW0ksRSTFMv1uO/hBrkh06O1G0fBoNkC3pMUOgnWOgrjU+G
tALAX+cTAaKM2ANUcENgwhW5J9V+cf104d7dQYqUebl9292T9RTToOZiKZt+h7Io
QkRIHQAnF6B8gQ8LYgwHHuLZNjdONTcApX5cO7nzyUe56l3xT/Ro7exLRp6JHzgn
Im/kcHMDZDLu4R+ryUI98Yt/1bvzDaUgk+gcWtQ9Wxfk5iFNTw92D7/nff/8nwuY
qbuPWAhxh7TxKzrtoRhezWUiARqSL9vIiPYygYIUOAE5LSLe/XjFe4OKxgyidlJl
aFUMssrglQyTjrJDQJaPGxSyiYF6YGhv5y0NEeYskjnMI1QZsbjGFoJZEIkzRlgb
l7eaGk01Q3EO7BhQAEfuTXlQa4/tCCZ0cjsYFlI2pCMjIZHfNFooKLfbHSUCpFQB
GoWD9rOmeNJrSdI/zgwGp6rWFGL4UGKNl/K5sMcX9LOpFRUmSohzEmeyDZdDfntt
/SRzZrnaD85gmNONWnLYfJGYkI53wbgU4g2tKFu7lftrCnPfydwZK3kBNRROWEwa
7n6zzMaJx8LNl47cZbCXl1riKPVifuBhVFpwCwjhDd2p97L4mtAHmLJCzPrGP/ZF
E5i99zwe/5L0yXCr9hw+o0cbBEy9CRq50fCtKqVR6/y8AAhR7Wetm7eX+beECUUW
o6CSdQm/hzWcg4/JxrRx+pPpWsonMQWfI2iJ7si6h+5Gk2mNJWPQKaTXr6Sn4k9V
VOhxdXZ7M27frgFvuV3shr4hA/pTBFzeYgGUWvAHHL49BlbtzJhJfJbEQXx445ek
DbL7AyzaZeDEi3ZYbSBT8fqigzoyLl6Kum6/sEMJMRrbjZaRh2runNP2Zji1xOS7
JEgMGFQChhU2IrG2upA8+wiNkGk3dmfoiKKeiG/AGIBMJu16oRTLzPG8gVymgmii
USTl8sWtv0kSRBdJCwbypbFSzk11VW3r/g/B1jo9IzBUZKpeYNjUp+NBuDqUR8eY
hHm3W/sqKDPXBouMDpAjq4QT+ZTILvJtVBYAwIx6qEQgSgA7COOSL1PTnwmYxox5
Q2LT2dhXWuso6h7sMQgpMUBvlidHJVTNVnEDwDDmRZtbngnNlgL7bmN4xvQWbdfE
XwGUxIuxXn4ea6R2yCpWW9xCreVqNOeu0fPyw91yMmRGgHfQSA5M1oqUDopfg+nU
D2iIBQaIygcYLeFK9O35hX7P8DacUsPXeCFAg4CxjHZ7R2UrPaUXwYz1qqhf00TC
Q3ayjz1cChzlXz3feIrMeF+u3oCEoUQvVo3CGIUZYPKs4fMiKPJ83yU1XwXJqgMx
K7L1EMV9vayhesJM26Xa6trec/WNwZViUrVxBSbiAW0VxTZgbRI2HOl3UntOTR+G
2V6jyiKWiQsOKvrWSmol58IqZTRADJ9PmhnrhGqSEntGYNwkn1Sk2flNSEBlfB8+
I5PaoWsh+RMEkNCgMwQGQ0Chh31VwCr9ZB4+BFgcFsGI/Yj+903ojZ1nqpZvqM0X
fxNyeyQqqjaCWiVkZzYK7HeOnqE+DF0GOpGc5pjTOYirekYEL2NekE/N0bEkmt4/
GyPkAkbqTEJzzNtBDfit2a1N8JWlVOpMWcwpmW8znlxfuwVgFQUlSpkCdDJXoLnw
GL8IMU7O2AW1UQqg0uj+Q9Y++acv6omF4xQaM+aEq8XHhdo0NydyPCdyLBdhXAvH
/7lxuUqLCP2W7fDTgNxWLrEoSeHO0E6FSSv0fW8Wjzd5uxbTFTgCHqDGTkpcl69x
Wru0sGqOSBzNOUyDq4stceyvYExbAPn88+3BIJDkoYoGKRsiatURS2T/aMBS16dF
FYUgV6jQWJNhYiSdk4iStbaAX29iP96Afr8u5AeafKacKMAqgw3dWfPblkEX2SZo
2Jiujd/YCOmGzPgmjfPVZHV3A3ppyqxanK3Xc01nzTQ6ahIyvBYhIuuAGSIg3AlX
zh0khxGaCbA5lLCOd5I62bY6gOggvFnvFkzLWJztsFS6MUlwj7TXyoNM0GE88tOj
yFgni4d1IFM8jkV/UDaBTbRXUzkY08xoNLeeiVeKSLjCIRVS3wK4oxhpLLerr7mI
RipwfkhEigd8h6ZXD5pO/S3mlfGVe4N7th4amiOl9BduHHwCkOM7j5hLF+DjpxE8
rY8/Her2tPFgoCxSQxp2mEdS3vHlLm6yeU+gnPfhkkfw/wloiaPQl5mkhm0xSZ1j
GW8lrEbrKX24Y28yOkhdecrngg7xnkA4x2J/Fp6tjT4BgWUYidelor6P6L4FS8C7
hS8/4qU8HjVAfmJ3athg7pJW3xyGT7Yeuj+DDeL7/8v8IkbtCbhC6FQieYLoZaUU
PCdd8S+jJiQwisP3VxLjHwrSRsQaZjMMJu1t3fmFmrHPbvmyuuwX3SKWtPnaHlOf
jeWK/vLqADnORqEqSDi3+KF9O9gaW8qH9dYqARRGfOBlvz9aX6Oo/SDjRnnudHCU
ciiLahxbWks/V5c/9VGhuoGYra/2OWMB5yeyJV9DZN4FVXx1hgZV42WXcHBSESK5
pc8M64mPgffVWWjftQwxwdW2bUe5sdweqAJLm0apaOenoU6L6GjxIJeveBkZKxAv
aHOOnYjMl4YSMhHn05NaYjt8mjVt88QlBdiO6LLcR1ys1C3vs92g3zCUf1Hq2ci9
Gk70hi6U6bbcxsxRqc5hRMe2PeSBLuuRrjYKAQe/v9fb37e3XzoN8/Aa4OaFgrNR
848ust5O9gWbfy1xfvXkl20FYkVnRVzl4G30PCYR0gVxQa98oTtoxrR3ADSMFiD6
Lxeuqf1u8IoXrCcyESeNZt8kfiPfETc4eWOepAxQVYRWQPl2Suad8zNd6RV3Iq+J
MgwvtTb5Iip2OxQFEFABRtPYXNn8wx3rpW6Jwv9qt9g/ygST63ZJiItjhoaFaOyY
qbb8fRmNkN1PDuX9lNMeNAeRnJoIc5w+gn1OdIvVOAEfgRZJxYeiphO8mcSHBLiv
dsseTEUUT0+gyq5rFjDBK1huriimuV56LF6YNyHS2iHQ0exacZt+j/6vV85CFQkD
FwMUMPl/9SBDUNk7IhBFnNgSywbexg0Tdfkq5gmHyCSBuI1CgjSSuSBNkRNPKrfb
qAJ2BMPjDjpcW72FbAinJYa2hrc+08ZaTc3XzR3NIMUd4RcBX9sqC2dBra/Rwmze
WLyfRTITXdw32wjCH5HbqNjDSEDu/5oV4pfKkHNxO+Eg+jcNZsENM5orH5GAnZs5
rU7zo/tReLH8T6UanttbRrM2Xrw458kLayIy03TBhU7Ah2riyVo1zwi0rkfd/nqu
clx0hzFPYj2XZ8vl5sbrKMLnXJL4cAPuVv2Zi/gcN47qdQNlUsZP7HdPSLc1dOqb
KgnEoOFgOU/47fHcr7DUM+6EJW3L8b6x4b0pKD55LcRW4O7lpufIjXkRbPE4XEdi
4dwPGyLbYkAMpjduvcATN3X8ry+6vG8mERiY8bG0MSjmXBErffnXmBTbvkau9VDK
9p/JtihqrkE/tcH+w3KZr7ylF/srAL+gdrY6te/blXZVCczj+gyatSZDcKexdgXK
zrcS1VSaRD1dte6AQHoVJM4dJ4Mk7nKnTzp4dvfiMCdqEHa/PVqGEdzozjaVgp7b
grSX6p9idDIK5R2WiUiA/g3lxGwJpJPiNcivh1zi0QWB+VJqXjrLSYW61QxkNNR0
xtnbdkeNyZ/uJWWl3t+gWvQf9zAQ95wSbYoOC2yXDRlMiKgtp09nGCmZyOCtN1gc
JpHPEIaPR7ht5w01JnxuKNPfSvhsyqZrdTdUIQ4kMtpECSC2YkuIyTt9n5bqusjV
aQeN7fbAI5ghvz6V6b9jE3NbxPYG6ECv0ddzFUYy0WoEuxTMGVXgBc/2Sl8mpLlW
us9MHvd0e563RBHkFDHvxWzbHmVsAdNtoUPPcLQDVI81pAQfrLmDFpc5nR3skmDL
NJtkx9MwshsLrO275qEphpls43OzJp8Zt5sMndW6K0IH5mG0OkBIbV3wL5hbbOUn
7HUwSTphddezjCWlww6O/dD1BwfWKj+lz6a5bVgneptJr5CJDE1x3UFaTTaw+OQu
5qqdbsbEM9XSLSOWaC/AP/54e87pmHDMRcickeqB6Gq03pNnCAcD8Yb3xlq6PkI4
kK0Y0a2lf/VaH9DD4TifVZXgJv8REkvDCebTi2T+ehYY/EPn5WCu7sTkZUMWUZiR
Jqt1HNeHH41AiMI2xah2CA79sU0x/wdyE6TzNwUEnHon//rb44vD32guHJSi3iC8
IfyvgT0fqLjyHR2UHNKiPILLgqzvxpbpT61mQ0p0oI5NfO4tTCqEnfb2c9yE4aB3
T4UN2oH3MH3v1cwdUS0Sxmg1NgCzuDCHsoNd9HYKZEWNzvaqjGZIfeWcZtFy0sEo
EhOp7gGq0C7qX39QnHoWzTA0tTSahekvigHg7QAosJpZXfi0Inbv6cYp10r4Me2C
HXlAhgKJPczOMAu8HgsVvXeZtDHJ6HCstj9mUAnX3/GjcKjhf8csMZan/I2hrux2
bgkSU+F87rGsK/6NhlJ5BUf1IOocMsTHFTtH3lPGI3twxD/NsEUxIRb8o6M9/nWB
VCpXzlX0X+4IEqoLT9v9hXigzU6nRBACwFo6Ey21ED3qgyIhJUNreDh7cF8jLFUt
hKO7kvLgSAy7V0hvl87A7mpmshXEoormVdvZDgJdeWZHLhUYD/eFca6wChOEXsvN
DFrfQY/vw9O3xCj10vORehA8OMX6QKdSWne8SpOGfm9aObXcHU/P67arHHONMLYu
Ao1b/IrDyBDRzylNthvxGLLZi+dvkQUIq99IGXjlj0+zUABwD59x0dLTuEwE34rI
KAP/DzMSHA3KNTG5d+45kMFYTprp60NihM0yHRt6E/plmjPWRggRmbDsdWKT8wVT
tAWJEeWfzBl9CuLp/3oBooaG5dJP9xElpnT8VfF2Aa1F69Y+myiVCmZg3DVCOhNU
Id3qT2G1Mt2Nh033VORBs74adl3XFS5RxhqhqdZzLVjsJ10wBh2iQwtzMX+xp//W
xlFyL+A93S+KmdMJzksERy2zMzYam1LV0NfIwg3XgtHYl2H4fmpP2hCayj3nDO5i
lCgoc6HgNQFBrMXR/RbJ1q9QUy5ivlcwoxjw1nlietNMwXuVCsYKrrX5wNgAadz0
PKKlD6d7V0SRdn7KhCYnw26Gb4udXCWs3PkjmJ+Hd6jRQ8kFjUFz4VW8o0BVViAg
XgmbGVpg0GGu72alPHSUHGLZ5Rm7zLr5IWygUIFYhs1oKCerCUbMOOyevc4kY1i5
fxylo47o8etY/pc7IcSSFnlnrxjjZG5JjqomXQCNAxREiqC4kepY9rhmNQwCivDK
0iIjxI8EtsFgJd0Y0XZTLVAMBItwDO72Wf/tNGA2qRyG5qFKaKiCOrIdEZ3e5LUH
pEfIvlBMziWXkSKZqSADKIb55rBmga1Y02HXshmjk9l/wS5E0vy16VxLnYw/8AUA
JRLjGYd5h16VHKV8DePlJFhBz391UxQHZhs8K4n7UamxrRMq/G72NFhq9fI6eJEJ
9SCodiF8Yh1U3eV0heEGlUNoBR6QFk4p+nr1qzo3dL0kbhyLkSIyzctjTALplx+u
wJcIeS4RYXCOxxkgmtjAByMUgjEPROW+ggYmxJ/j8tLvjR8Zcn8541DRonD873vq
wpFwkYzaAnVUq9saxj11H4QKrZ1HrjREav1rdiEMyzlSkc3YFKiQSpgYCAWf4Gy7
rSUV8M+VNb+fp+YYZ8HGGoqo21BvaowhY/C+qN6UUItButdFHuoeCo1g7FLhfhel
oaUXKwNJ9123RCsm42DVLi93zHCcmXRKyIE4sjdnGwX+fHQ4OrxW/Gj8N8bIGfo4
YYtrEGa83xUFRn8h9zka+/BBFQLjvWduW1WL2JehNBCDTW/DeUNwwjwWLa7RXPES
u5cPO9GsIXVph/e+mb1Rd+TWiUwj5j+UkTD5cQn6B7lhswjyV1N0EN3p8RIYObKn
tEKtNexB+0lj33jQWrVfBgrVv4PfO04jO/nWyz8samQMd0DRxD8iOQpyhEjJU4UN
obqJI2bMqgGOZmQWDyVwcVbZChcJhtcyNGR1dy88K4XMvXRsjubBq5/etx0OT8jh
EDFG9/LqgSwSRjVlJHsZBTig0/bR99E154iacRcn7Yz1j1l9Z33QULbevHsJv1ou
PedDyozEKHfI9wqRd7HagScqOzsNDnYNRn07ltCowggpEAqwU1ltvD+Lq8kXXZKm
`pragma protect end_protected
