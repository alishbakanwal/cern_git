// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:05:44 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
hIvm+iKsf65Z8WRk2chYESYjVKJSmmomHYkCNYts9MbtyqcLB9AhAEvRSkqlD2pq
mddwJNNeBX5J/zashqFNjHL/eSx3K68xX0s7tVIitosMPsMBTkmp3hCCJVbZoWiD
nzxpFsIreq2lyUWnq8Vl1Z8grzc4ws0iWl9pHmSYoFo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6416)
PnXpT9FJRJvhO/zBVmbzMcXat5zG9tUxDXDiH2GQnpuW/1A9Hd3hMFVgofwTIojB
1ld8NmBDIgLYXXx5/zzmdGFJIhV6EmWkLE8F+OUMJyBd1robt7tJ8NQCxhfhTxxA
/CO/kUvsQLg87BzZwP2CdI6tTbZ7eexP1jaiA5K4Wz97LWtgtIC6t0+AZ3xtT+AU
Hq+UQGtlqudwG+85piOVOIwDXACzoDw5h+CX/o8omfiXKf2IakeRVHphROk0hZ+v
n+GlmKLBvfRuJTvPxcnLjj+vc4irJOJWNDVLT8nuh8iG8XVLpzrZfZ/7hk+fe+xK
BKYVvHBWCheVFmgbIsqBOXcVvWa7lOD/l2mc0xJ3fOMRfQxFko3/EYhi5ZMIcAfY
CSkhsqkJ1SJFCbB/0pNA2CA7Q4dDOVkks/VKgTNJ+6gNpG2iY7+I0S9N/yzc586c
/aDBEAx7tJLOD+R62d9/JAzsNenan+bW6V/5HgbqR0+lJ0Ci3hOLe1t0uLiBw9T2
Cxj/hghF0tXEYooh8D9uZcVLi6ReE+Uixlu6VlueCaR0FM+Cu7vj8iONqYEj1Aqo
piPNeD+EqdsES2WTBUVvHHxk4/5WRUN4q2yclEsomV5xMAVyEg7F8P1AoRIRj0F/
PTv/OIlvdfdfhporL0lUA5tQC7+BGh6AWRZHw4ZGHsTXcU5CMrdycAAhECWHq3YN
xlT88I0aeMIswfYVmLbWvSbxSCQ0p/OC8kXw5Uma+OdG70ytAczL8miXl6OrYFFA
NZjMYf94qe3QjJwHP+TpClLmZYHix8CJ9wQQ8R0UF5HKfTeLCbnPxKX5v1PDhEdW
ftWaahrXXLa9szwP/sk3w8UkEKN8QM+o9AejNrlZKLDEGDq/YH/u2CQEW3jwxwKy
4GU5QieryjnQY1AltV9Mpl8koHesj3fRLVcf+Mc22mULkRUl/UungPlH2dO/Sskp
NLbIEsnXNRf35wPIbtG8OOyVzvv+1Whn6NqoRKeaEDgfAcbiNbNKTn9ryjZ9F/u/
raa/dpyjJkK/bUGFlsHGQdMVDUEYHJjj5UV5Nkl2/mhnpCeVcQeZwoESKIJegbFK
IKCnW4KMkzCLJyiK7WEv+Us8G6ixzcCGzQlK7v2aUCcPb5gUvVsCNRaqQi6hhXNg
l6RMAmfAxLXmSouNtA1U7CgADszfLf24TkDJXf0mmkI4YWlqgxUj+jKFUbRgB2Uk
f2UAYdzdgYEnWxi7opj4soDqMh5pZI3SbP4E1DsS81naaLdbI7w/N1FgTtAxeM4q
xmvJ7VP5EDn2Rmp2DJpxEnpx8Cns7bdrIAQ7P83cyofNrnBq516FgQg4w6puS6SS
lPFwPtolPdsBbbx1URP189ppcNLdjrTf8+fwNU5KYNccN8XLttaAQd0clMvxsxpR
8q7IvRQpeh5bB+Hme8rH8LlrmeZXnm5c7GBGoLMFkzrr4kwRVpCLsrf5bnUE+f9I
0HLWpmTRlfJq+sPeNQ03Zjkyu2+6I1IFjrqEZ61qDQGN39xgvj1k30weHFKibRbY
Vv/86k7DTZjWvZP4aIUKqeH8GTxCNH4sfgdgDeUU//oB1ZErhsBU0LYFfGWjwGax
B8TLbCfbjzKzIT8rOdWQcz+z51ju1s14iJmt0Bnn516DFyHHH568Uo67N1/X3Lwl
37B9KgLNsfeKdmKNqWIjGuy+ZU97XSxeUsiT3gHgMRB5VUuex0+TPqcnyktkxen8
HuvQV7BsPRc9L8/o2UcMwAIQGWI3KSsL27BQOECWjaVqd0b+Mv0MeUTPVxv/9EKW
IFMffVB67mUnSQWporVrTk7sKhw+OlemnAMiY3vDYQAkXd3u/BOFvc1MQL0WxEIm
/z8eNfioxHLCBvNKUxzaxW5aEnGbwv5QlrZMGa7hoq3iS5qck1AmqBm/FnfcOfn7
WEWczLbAxRTwqv5x+i79GR8Se34q5nQS3/jPDfJ74dLvYiH220EyJQ03iS56V9Zx
nQ9OIzdzQq/UBFrlOs8wEsajJA+W+iQRhBfPMHRF68Ci+05Ais4r3CFSQs1VkjwK
ZsaiAyTgzH86u8rHFzJMFh0GnaudXOfB2Kci9B5ywx4CDIIYV0m7e+dBPgWdUjpN
kqUn6us3VfMX0aHVVG6TFgda9UPCZM3VRARkIg7ORo00Mg0Ql8ZmnTYkAic5fCcm
AtnJrdhuxIZ/g4cI1+TwSfQEmIDksrfr776dy0wAtk0XQ23lBfLeXlFHEemU0Zej
29UkcO5HmFMm5cSTwHo/fE9pvM3RSiFgwbwAZz/hVjcmhA+gz1BNnOsi0sIBCGnP
a9oRUIThD1nleuq0p98CjdS25D4QVxCvTHVGRE9ykUx6VCxAk/qC2t9hr50GFDgi
pove70IO+Ka9NhxiP5PY3jaBpZ6VJnIk0AedC5dEFzF+12D5AewqG9yp74hE/AqH
0fM9hmeHlefeWjJAkUXjQgIne0qbRQMqsRapwm7aM+ctRvHIR6yZHFRU73F2PoL8
tclKQRy6fFZE/RF2xFxf0YouXMeLPnwipqzheFeid02klSdpxB/Ai439QYfKmwvV
pd8ERvjUXdYOahFx/RJuGi1tVACvPVQdgGbMBnELiq6PryGS8n1gUBfI3XLBryPd
BqBKHEUSwWx9txwelMEZOBOeTq3guoKvIEddTaCa3akWI5GW4ifD0uqOMUwF4kRO
nSLCS36c/uiJcPAMtvlTYcul1TLc7vnuNTDtRQxUeqjT3DMYVkAxa+y/5WYqb3gz
pHwIszM8JGnL9HfQ983x7qi6l3SnuI4lBUWAfGGIjOag/SZrQaGsh3kAxPmKF3Xv
tJhR+7YPg9XHyD42XXZm0FHMPWEw195YEeZjU4tAmY6DgrucVe1Lk1cDcglJ9+e1
JluikNzE08VNAmUcsnS++yXfYwN9xWA7k9Y43Jy4OdaqIwJTw/BbIWgHt8twIAV2
86Oc3V41Gbd/d9hzO/DsvE7d4gFC5Dxsd0u1hWM5xr+nIdYX6XpwSicVeydMPIC5
3uAS8paL6U122REAzAggSBXuPfZsXbvsvfaZ95DRqblF+yf5Bi/DUac0SS1+qKga
D2C/ekDf9B4isrn9Dqx/E1EZa0Tor5y/35VE4pz4cIzMqbr3BkP9nryIzef76wbx
VJfydnSHpUuBebU/Ds3mF6b1ppr2Bc6LdsQhGEvsujLgRSotqBevkI+jtJ4MHTb4
lHddDM8osY3YHok8Yul5LVaN7tozO4uBZ91lk3vGNoy4zd/UkumQDqyp5azOZW1W
TWQcQ0khA7taJu+D+KKghkbGUhhjf56YWlkiA3LGLMporGbmSaBf1Nnk+i1bcJIw
J2/C2U9zNwh9zmi3xIEwvI2qq/mDp2nV1+0Q5s0bYm2DNzfDOgblPAzXauNN/ood
VA5CyFBOheUZuzXFTDq7su/CSPfs2vWgsjUCNancR+kX6x4f7Ea59ujTaNJFYmwM
xZjkgmvxI9hd/Km7WvWm0g8ab6HPvfTTQYTeULei8twsvGWW+0dFUu5SzA16zb5K
tKr9UQ4C8+SoZduyvDaysvB6YUnHkxZrWwwVvh+kz9a1rQy3Cm/qrOecy93nvrWp
kB/8Jhq+lhp4cp+73BbwslJBm4EIBgaYvUB+cLS8h0bUy6O+rzk0mktztYh+V4P5
rYgf1fOZ5vQjEzb77t0CLXQqNQdfKPct6A1defEaCX0OtL817RONNA6BUNoDn23m
HBNgBDkcTz/Yw7ed471/IJh24RW3HAA3VcAaH4psWwhoODrIMSXIHa/Cyt8v8d/W
oMZ9q7y82n2qyQsrJnYp8+wZDpkSUO/AnDCpQasX3eGvVpuySdarLeyQBVrrfu78
nfVqO/r/WwhRrFTvRIuvZgdyhxCBfar/HBYarrvt5MSXHgoihJXaKWZbpjBQLemj
zUfNe+6t3Ht/irf0wNOcblEsbJo0iysninHUgZ5bGXtytBihU6AUDymn22fkUC4j
Ya+jzfjC2is2CTlJyW2oOwhGwxWFK5jXPz3ldvGkq10cZmTfVfQw6eecnvXiS3rK
WTgW7yfaQXrdDJeqPmhD4CM07oAJA9fk8T+SHTJDGcx2jOpHALbZ5ze1Vdy08xCH
Vx9qeSGfa+FySANg9q4nMyCndi1dgxCklI0B02ZEogBynCDA8JO00KqqHAQ6SkkF
rHmB364kWAtuGSD3sJvg+kBJYoyAHCLt81fWfapDW9mFrTunpLPJt7bcLJLHahfc
/bUGYwc6qF2NeAaAvnMFqHJ+yJ42XU3mSC3cZxcij9XTR0ZyV/Mk6JM+rT9O1ljg
3IQGYV2inkMXZUvbkqyInhzroGCBa2BlTC/cLth6Pvp1/FJWxBJZlynj6wqYvb6x
TT4B2BVhMnIwzDTyHMJyhfy72jpxxRuB3+pB8SfUs8n4CZGAx5AgRGoPGj400mfi
VRrA3YTIqNtY/GF33zMaFpYNHkcsLaTM1KP2XVTN4+hgZZULcTX6aSgk3O2cRm28
0cMlp7b+8AN8d/dPlWX2476ILFjH/y6kRUk6BQLu4xwmEWJ08/yNbGRx7TaCIpVR
A3inA97Op+fbdwbD6kV48kBrPZrLTCiCg7XuCTDY0lLHUQtmRISdIBEWwlrE7UEv
6eUgg/4TWWkjwgHrQvNhYgh8k1gyKQXjBAPf/Ia3h+f+LQTt96BVopOgUXZpeXw0
5B3pv+X2X1bjHjNYfApTYl2iSZ4cwQbusgbdNqOhyvcogv0XwL1/d+svovgyh5kf
COXgzBO6pKm9+W0Zn+ThUhVeOnFGrurfuPABxz4Hsc/quNfZC6SLXz/6oQCrMrwz
tf1XS59WIvJxIX1HF6H0HKDf4Gw9QzuN/2780JmTkNl+RZZqHjrAymn5vpX/B2eF
ojHcxcfe9KxQWOsVFo4Dry7MwsFk/4J0E3rexXWFE3GalTrH3k5pQEoRxP7Xq+FG
11W0GSpHNPr5QsyEbj6BiD+tgPq4Nk7XcRiVxnI7cbFZaGGbvi0xUjxh5+ZVujmP
BSYiaGw+kUaUjP4VgOMNapTJcuQXUdJUeekpAr6FFKYyM8Jypd7f2jPwErbZHfhp
EMMTwpbyGG9U25Xjt0cjB8lxZJPY33+ekhAoFMFyTLub22cQMxRNGdCGoI4Kqf1i
D7DxLe1xcBtGpu5dFOuErogvRCtrysjoimiU3GeoS51mXyJL3CdLYppNVMJQBO/n
Tb7RiKVtgf1dWutY0HOZVJ8RfP3fIy/3TOsVnrpXmWSy/k1KvLwjmdUuhF5r/Ggt
DhdqHJM3s+6we3fDtDkDbY5n6U8ea7W1B/UEqVt/PG/o7kyM+Ie1p+blCXx1KsR5
HPDAxDt4kCuRq1qIelAU102McRO6bxj1qSN2zYHxHzVLPyWJ+nhhnhEDSLvJNEeo
yGN6P+rW1qdrX2Qfbl0aGoAEM6F0NmLVKWdyLjwqEv6dhbr6eVptXJJdbk80O2Tf
fQphYFJLxpnEGd60jzyiifR6l3Ni1cXKb9/6orqzVbbqf2mueDgzE1aVhOPGEpky
eOTnGxg7t0CTeH8FkGm1OO8AIP3R/hob1CrcKsQxm2zjM9shJeJU29aKgi6d+3N/
3hOG0lx5+YGvEL2ohqYS4j4GT0VokU/M1k9t+XQB3N+Wi9uqXrF3KwNbXYQyFskI
aTGVyuuFaA6afTtKotfZlgWLMWLhvwMuz0vAoEnckKsK+QGDBspspktCNuCYvvR5
6o0rNSOeAHwifrH9Q8VXMGyuEoA01SSll6sFi1MK35eJzbvMuwEqAHoizQm/Km9j
5YXElR2IlcIzs28ri56Ukcr4dBod5bijWgebTi/OhkoFVyHoAbpoANLUh9Kxs8CT
tqf7u9QXUeM2j/KlAyFprW1rwsLthnx9bVk3Yl6Io6rnFXcGjyFthm83sZGJ3kDb
PqB1T88jL+JNV8XxgGYdEsBJpxHa5l6F1v22Q63o8Agdwshh6FGbRSEwGOz+GYhz
YFLmU7EY7PZq95lLdCgFeluRrdxfAxyvn9CJEAoqIrvvE2pLNkdXFeHlseCyZuPE
5eUrvX7M60cyVfAulFeVuYn+3opsM6QfzYNXg3IKFLh1N35fLDui3xnY8t2tDUUU
LEkCwwEc0Ym/N0sDLQN3cCa2SNJouWnzVIUQNrf2xWvGMAJqlrnANYxnnJiaZnHB
leWDzhrbQqmqVd1rllfdC8T4+GEK57tn1wEyIcWt87rnz51FlWZDMRs1TkbbVA/E
dHW5mwAsWzzAyFu4G7qiM43jnq9CZw40AIreR2B0kSYsH5Gl18UoKK/ymPxNLROL
CxIk6frzldufsNhEhgwFRfYPhh1WmjLz9nClpnDROEiAZtFekd0o7ttWqAbNWtq5
vLKJX2XeDI/bbCex2WRMrhHIBK7Hu5PqdISwxnGxCZbWHYbobrnalF1gnKQzQTYY
j4iBKeTSy9sT9ByXw36CnYIQ5LvWLL8LX3q/cxQb5nlVYhd8zUxB0UexktoRbStK
7EnNfyn3MB9K0OYURpGtT2BjxnJ8xP8vT6f9h/8mCNy18am3yt78iuSeorh1uY94
WTqxUTQ70SvnhaLrw1Kbp2nAhJzyILteIUAXIbbT2V7QTKxqQB2QDRBsPOqPbwyw
clinHBhNX8DjNduCGLogkRd5DCjdGMZJzKNg6GqiEEKfk5qksEZat+FYwaFZT2Iy
zaN68p8NfcmzgdSj5jnDgVnZ052e31mDq6L02BcZckKAPdBfaE0U5PcEgY9ZQyLx
Xx/OStVwdS1IkWleu1kO02PlJsDGdOvn01wyH4+KvSwt+q4jC9XVYVWY5uZPrb28
/pHjDWimv8WLfK6SXg8+Pe2NYfVLGOjToapunUL5iMYhYjsQ90VzxaTKty0Z82X6
zW2nfG5+057zGb5UYIfjUkDdl5Yj0sSOmAlA8uAJfhMNM7wnP2fxlopK1ul6njfb
LbCYAQ3tuSzGZPzZmpcujUzO4Z0RsCwHiRMZ7yt46u1YdG6Xs22Isx7t9ljLbSPy
0vRMUoaEGteQqWBtXl2wTJ6TIZvF+qMuboOpMEwYbcfXpst6LgR5rSuOu3hyX+KA
El/5w1hhiSp0SydU+A2P/ym2oZ+7E36NvBXmtvyp3jLSXXi/43pYGi34XGuPtdrm
+BZ8MCv3RNDaslciLggJApvEhkjBE4Tjslm9Htz7KQqGWwXNkCLXmUrUMMqKmAvL
mB+Y0z9Hr1mML9e+zWqExF6TNWlkax/E9FMDobHUje+IovP/pmpVYBC1udNkyH4m
gj5ByRB+n8thd7u8bfhQftVaEEEJZxnNGoTJ4DN3ZThzlpft7h356e+CT8r04gMB
W1qkpA1WcoUrGzQBU3XcblO9lI+B/qaLrZMc3J3okefCQa/3L72douDyV0e8qLAm
tceD91lK0iW53QUF74a5uGXXx0rUIgbZV+XZ187KlmYTQUpyBOMa9iSGmGLGxCMm
/2UHgudOosSITwY3ErswMY4iLnNPNB2/uc9d5OsiZgTYTodkk3Hx9iW6OjFo/xKF
OICSj+dcM4Dbs32tRF1y8U3wdiZ50CLh1vQTWipN8zt5FnLU/8uoaBuKSIErekgq
3M7QWEEGB5RkD4ol3mNsCS3VvOrQX+fOvwHVAMz8hws7IslfPOh1hkmhh2qT7pGN
kPjPdqYcdnGxdX9VBbMyyRY+5JMa61abl+MAQwI4ycHpMwHW3pa44OL0D8cMmr8A
Bj0ZPa6AoPlF4bK08LosgQ71tOLeyk2jA+dCGhrBynp/iIIjD9VY3tUld/Ma3YVX
/z30dtYEAWIBKnhRG5zyJvSCZOvMMI6BxTTnvPUjW7lcERT0tz8XkeQL1HLyXrno
vc/mufHCsJ+d9x3SGg/ieyY0JifBROrTzoogt4f5VRztgf5sg9HK+MwDaaOCvCvy
4WeZ1FaGHXySnd98ItnyFdPJQD/Ww7QGlA+9Vpp75uxopxr0fd+9Ik4LLGoCQF8K
Gk3tHVHxIrhOmlH25F4nj3wVyKbimUVcL98+J0Vy/jvliEEmouqpXPFrgWX5PGf9
6PMgVmESlWuMvofhHTtmOCv2p3GzIOtsW04hXauhgVq5P7zNO+H0S0MVYHUa4inp
urhQM2qWTBPa4OlqnLAChcV4Ff9RCZ4HeKZw6enshLSZxmGT7wcgEam+T2+uF42v
6iAcSSQdg65dPqHC/fxGusEkAzWtH1CJP+iWBPrt9oHN5dX1am1mlsMm/61HRREC
efqbLr24TJox01VkJgVkeQvNeMI/6fBAxlg49HAdLcFgyK36pADZ2IXrWtMTrOHq
Z61CIEl6hg2IlPPs1mpNf7iJ2c0JyHLdH58Uuv8rR9VqMckI91M9wNq8KTNmJuk7
RLtzfey3I/7uqpTqDNqkj3ZctcUmRTx3q3U/fdIFMju8ow7isXt72W0GKPTgYjMm
tUe1I1wvrOeC3qsDuqN5myPuXxTuLzr9GHI/tet+9LjEeMPN8tL77dr6nv3Wr1Io
AwYfooZVLzBFLWpn7HDLr0JRYq2/dXsBZ7QKXiSuJTCKr619BAPYGVL4sianXOG4
s2Xmf2ux29lrqa58+OS3bC3Xh/KaQRTfnvt+hnKS4oI=
`pragma protect end_protected
