// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:05:32 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
QAOa/Piiuq6Wl3S9F811Pt3OzgGbF2XxyNjCIbf8TXVjjciuf7iINJCLgl9MMyfI
Yr8WUFqzmfURSRg/PWn0o9YvwpwYUqgd8XPuVdOZreDCs9YXaUzoBWhcvS3hhLxt
VRlYxY/zr8U50jItOemoGT4NyeDjWocX+Mi9SVbakw4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 46192)
eRGqm5NRYrXlk83bXrVVEM37tYUi7rbjpwuSTDMwz5eOq5ZeBSVwTj5nQujulG5h
C8DbLBmPyoHRB23Xi/Q3USlZyyUZx9DmoVPjFm64hL5ycnG9BtbkDKrktLAfamZz
iJM3XC/yuYYR1n4sjRaMHEwEzy84dpMGUq1o5dJYAj5XObQ3XwrfxTGH7nxLQ+07
orHVMNR0Ohxfm+zif/Y4my3agOpz5C3mTdxhMQWI4TFHe/+E4tm+NCa/derX47EV
sZCyQSzb8hvhxgpFwhzHLbjdxM1PZgLw6DLC7AXPdoYIvyjH6aOeQtGqsdwScxY+
LCZEQXFkA5sLsl/uvpblSrqza0OxK8zKR0Yac1stiSreEVv6gN0jt/jsSfcxEMp5
pEI4kjwuiKQ+Ag3fXZPKJ4H8lK7T69Broe7GSkPM4TQ2wh1oO5REpwFezfy0e8c5
0AIpOeFu44cWy2VNATUdfLU4f8y7ZqbFh4XXWkGIl+p9Q+DMqbQgNYOZ6zgAwTzn
7r8dcho3o2RZhI169/aB6/vCpxHFIQ3HB0At694r6GOQDzZZpfcTBzFTbnZT7eUR
R9S8V4rbKN1yo/M1vot1+T3is7ddEAYxG6T2B9VA2xJq65fETdbQbV0z6p3EjyOm
KJknkhrOVfofQfB5VlLOld4+5sTrYcfC//NfWeE6x78EFlXdMKokj6/9/Wr32VrH
8jEwix3LqBKidBs4YApJbqBDkamFkk1MP7QOebsqDF8Xp8bv/thEwMmFlGJ+g068
7V1pYQR2zr1VY/uxiaMAAfgM0VzRZyTlizMeYGF+lw0J6ezhQKO41yqNR9Xys56a
QtxQwNVfzldTStjFN9LUYvid31HLVqMvozABNG+O779L4UcAQul8JoruvF7zn4FV
79KBJYEdtqK7Sej5zZgRWmFHlcjblGza9KkPSmQRtMX/cHAbyH+UGztPuWM59Umt
YQ4gw4vgm90z8yMMsxeBef5Kv8Dz/9JSJoSB9LVFf8HAtiVAjuWadrZmSMSLo7It
cu0cFjDX1QJqB3MyxLAAkTRGbEJukba1sBvo1Cw1JKaMSH3KLBKiIMjm/pgRM3qS
lFvrUuG2A9mLlDSsgxbRs8ao1QKsqNGAFWMla+NjbQ3DzUm6zHAWOeyf0mZMEpLZ
Qn82RQ7ML6cFgEEACFjgLh+4Iub/qdCzmaTn9yATeTOXwIwI3CbtrVEyVKOOk/Z9
WMaruBcPFaA32AuHLQo2OGkSTg8tpsl18YX0YGJ/+rpHa0qj9xc+FWRyLzNvZNb4
32NrNYmdTIceBfD+4Lw2H/WVELT2kl2F+DcwJme9vO1xlYXg0DI1ThdkyR88uduD
VCXl3NA058CneE0jQo/X7Leyh24CXwYnqb4/oOWJuxHb5D4N745eWrZPAwsklF0X
YUzn2J3wnoBlOCY+ZtqHEEWCCv0T7E1B5QM5zO/hfM0KLUgIerF0muk2hSaEHy7g
7+EzoGj3VZp6IdC8to1MUqsnzdu9xZH1GHlaK6HX0cRvxfbN2gcfPhha3ysKp0yL
93WfG6CiF8Bp3sBgBmEItAf/Vcg/6I8tFA627DCj1nWuuDEcxxH59O14MOpmCxZc
/XuJ1SYu9yP6cbkGyAeR5BeyJhALdlqsf8a/ZRsMrqPxHfoAMKnDOVXN1ebjLs8x
9luwvY8i58UT3r78BYQ3+m0H/yXh32fublGtKpwisKxKyPm3+PnA44QeHE5eoTpa
PZ9Jmc3HuO1sq6M/8ie0jpDIQb+XQEnBYKRITx/IhfL4t8ckT+NhOLJvep9i33ez
tqVq/Tz9yXXaCVBnJb39et41iIHrNvALaJHJkhnz/SWxMoHpcl6O/QHLBDRUQwuj
001EXIhW3ZEEPcYP289m/SRduIxcvLodvsXNyMNnl+4xqS3sHDK+pWB5QXhNvn7k
p0VdDq/Or+rgarpZy9WRSxhRSTIAml/Xddjs+OjGmHGo3Gks5sO8vXZhxDKFhucu
nCXuePjck/q/KJwPCQb5PQJxEDef64KMEcnSPDvUkHhz9AxayWxpbPQsnnYc7aGR
OE4L9fiXSnV6St5TUl2Ww0Ed3Ox5QZpyses5NCVydPUPZOLGvP/2c3tVJZ/MkNUS
iv/k9k1QoT8yHpT5VaUyulzcwRZc4wZiMLyqwf45dkw6SA49w+SErSa/E9BNYBxN
rKHwJWg6bifkyoSsZtBHflImWuxAHxc41SGuCrOnzmHr6HyRT9dc5zvIIn2Hth+d
bk9eixbdcIQ1LDvpOxJY6Ey44FH1UtpsumuOjmGLhDMbhxKR2O/pYolxZ4d8BtJQ
a2JJVdt1lziFxuoSt+OvDPxLCLVlxIuaMY/vaqWn9d2TL8GaIdA5kjHX/+Mqw7cs
M1WbiyllpYE0AgmAqWdgan1QWBNfWvu6B1LWlrzWqXpfSp1DanldkzlIHd6IRKYW
w1lWGcAvBOkO1sGfnYmzXyP5s3+3DmqdpzC9Z4I0tqH0/yyKcY1NPIBkfWGnA3Pp
/w+rmF1FXELjW1XlgL0s6yea2MGctb9ZhJrHIyzp9DQdEGSynNi8Dl0O/ojx0jWj
mnqYmwsc3LPVC3Yn3npbRa+cUTP/37Jyntnc8N0q0umAE8907CV2xJfHIr/QfdPn
7yK5Z2fOiJLu3oyHHB4v5di8Qac3ny+77iATvXzCQ9RQq//77YbyXmRpQ7EEInv0
Om7Js/03fgLrUViPr1o1RSWFw+h8TubRjrpz7/eaBCsbogI5py5JEx7UusqQf3za
DSp5sYURO5iuknmAzaEgM8kRtHKkfgwiJu//3hhrNWyhEYZnNH2vNy3U4hh3MGFj
PK9zQhA6IBuRuWPVNN74wSk1y1RPJo69wlJcBdajhj/iMgqw933yIKh9YCsIHzzS
WxaJQAchE5g408GfMxgWYMN1l2bG+s1A2x2xDWJ3VY8n6U66uzQiZIvK1LQPpsXB
KERg5z9RrL8Zay7KiAFTMwNE0so9RBAk4AGam9c7q/I584vk67lN86m+8bupY30z
pSOG38B5j3jGL7CDaViEhkgHDBOIOn2gCN6OdzpetqKe0Bxpia9yE8vz+xWQ8bdN
i+/u0sD4kNPEuvh7vXcOuWtJd7EI7O1qdM7LBmniu+yVq9VphMpX6YioiLMCO0SD
juBryAm693IHKFJBp5KcHvmR/yyEpKSk+Ia9PV+E659zkYiFQw2DrHoFwYzLXRHg
h+DfpcEucTPcJMnuRldkfJeX94G8iziCpWRoQTJw2TH2l7HepblGCBxIvzXIleZ0
gdJhR9FLFiVTGacF1XD4/dFAbbb40IT666A8KO11U86gWQ1+exQL2LkK5VyrT1j3
g5nisrOTHrlQhqN+PsIRceY0IbNPF2zOv6sv/46zaDiYRdAF4hiyfIr/FiMXWQgp
2VzZfB4qx+dHox5Hgc94hmHH3VyIuMwRfoiTqi5NKz9PSLRmTUr5evZMn6nHsiL6
vbK5IYjruaorMEHrsa9IWlnEvgYLoOAEFTkC2rxpJoVdcDidDYGoSXo33QWLnbKM
gOWCE4BVO7jlcn5E4xabEtlN6Rfsytks57+yEJ6UQKPjsA6PlkJeQWBprmCjX8Hv
dZJmsEpkZPCmy+1TR35IUmh1JKF3vaU0jVkfM4B3+kN0VHehp0BEhlLIfYSH3G7f
HEAGiMi2w9QuYd4w0vc4UlN/lZzRQoGdJWxmEHc26/DuqMmdm+eb2peAUxC2NLvi
snNNOPX3JGTiI0jnHUcUXutyjpfzlRK4/fKaFUP08y1WqAQbD+aI6IV61OoK5Pt/
jKlP5leUem2RyRAGwWUoKCGOi9V6jAUktcnLGgRLapD8lyzMP2D3XSp/jXtdQvJA
UVZ9pfNuigHR+UCo/PYvhjWHJjWlJpxdaZQVRCuQXqcPILQaUmFW1wTU+WUs8Vkt
xormpCk+rAeEPGFFmdTp9NOqH1vqHvehfX8i8YSUMGLmTmVlXcO6un+nVrKTb1yA
GRefRwKlCpbbKls7XaxDpafR+uCl12iq7yjLGb0+XEILltrh+g/CNBLYtiWAaYM8
pyTKaByLSrlQzYk9C1LS0SMn+GoXPS/cJk2vjGqZo0GwuMM0Akasdf8wtUGjh6tF
nmmKLQQOayaa4+wOwx6ZZRwbpgeLYPstw2QLz9iyd3lafIZ6xhonMkQORVV5S7JX
jbIpUCF496v0uY10XCYxlX7uZU7qbKPzbzRrc5Ch0S/Z37d3nRNPOt1KAwoqzd7s
TklVmrM+hDwE6Wd3z/RWNN6bIy+n6vqaj/vHh5RH7Go7h9QdtnZuaFrJQxqzKe+p
jpJQg8tmr0YkyfRikzGUHA9deu0Prd60cHH0aIWJEjOYgLCShANzwYeXt29aYjJQ
6HUBbi80fUjWULQDek7CqSxBIZrveJ0B2myYpYLeySUU9GtS9cSAgcag/UlR5SRg
R5tK7D9QVZ7bniulrI7dgDoU7BkNoKcPZuoy4t8C/FPLA7BXNNc48eFpbYi3M/Ks
8w9ncs8ulZIPUJlto/lJHu0fWX6hRsxjbepI0056sLPYgacMxVUgpvvemA7BY1e7
GcIBgjDpdNZlVdhPOML0qfLye4KpUjN8BiOVHUP1xf8obxG9gvk3buRlA96CQ2Bl
KSbu2ogkRdH/DdRWqUC5gWxydK0B3+GDR37qN6iVMYo3DFAU0iXJTTkIAQNUdt8d
yWUct88SYwxbGHLmZ4+42brSNVl2qQB8Hzuy3+3ym82B6WlvOZUgKC0c+o3cDQwA
JfM9sjjBbdv3DuFYXQR8uPoJ1cQkvmqXFG5aLD+GuekRX+nBoon8syYuz7RWwueV
8WjpP+1ps5nxXq6NOWMVsf3nxXY3SYhJmYiUMxHKSBW5rhibCusblPn/i0YhBnJT
0uNpdDUn5KwBYQPoG517TUbloi4jfdPc4S6vvHS/YBvZWk/iogBeD/XIgTm4Gefu
mAxVH2Wy2D4pz7aS8RbmpDz8M9AXLatyCq/ASDpk6at5NneZAlnt614Z1n+OFM9o
7FRSEEe9O4TwQ4FzMaTpMniDK9rfs5SrvongLG5vCNYhVZB6tELVD6C+OsL2WdJT
UPvV1kkiPmwMHfkufJnrd0N4GHoc5pBaihCNxChfH2OM/2JfN0f/vrYbafq2X1Me
TjjaYqJNcyPI/TRDV0yMcHLObJUOJgCNXMIN48Wb4RjtKyq0wfzbiHNR0Rua72pa
KNlFuFsGPMg/49L86OWj2w28wOFqTwdQqntJZqs2kP02v9Cd6at9hV41ELplR0D3
b8U8xavCXR2zlwKsb45gQQGhQLVbjETUzf6AoNNwMMIW65Hrb5WiGsGbghwbm9Qj
JosOC3pQpUy70L53Nq6DIMBb9eXMCu/pA/U5Ui5GDiGlD/pXym9TbnYQ+w7cQNlN
6L1VO+t94+dNrPN0dqWSZpvvhVztnCUjY41rq1fO9Vqv8oQbcVRlowTfOl8BTofp
vb99itIQb7xcnaS+1F/TwGTOlgrgPMkS1TIVceQWa4oTwD1TjTsQ4ogHJlrIUMYS
XCz7GABsrQW4sc4COAojxM+oPXsqpXzuWhMu3FH/BA2IYyrVIBbywEGrluNHHboh
hDBXtrnR17L2Fwb65wO5s/k8zkN9EWsWPXBEAA10oAaSpEfhhLp1ZwbLbnTEHGdU
KC6W8TGHsWCXcIt5ZWLPTm0H+tp0acPhcBTCCp9YodMFRYKcbkdmiyEBhUExR1Qq
dowK82Gh8x4zCgLGYy6eitahRzranc4spPzcW6wdZL8pSrFaayxQqZyXDC4mTBIG
deujxfIl6y3+gvxosYLytV7nEBGgkxKztPU70c2QB+XZxR/9+WPExBXijnG0h1CR
+LV1yOzi2n/ka8EEGX12/9OMSFEahMMsM0rYVIbwZLvkTuT0jnsw/RIz/ViUr7D1
2q7CryFMnC3t6ERUHD8QtDvU+v4epP+bsJetJyb+KSfWy9gNrpRug3WouzsCnHBp
TE6ImAZwMEdmanF8WzWhbmBFxKAD3jE+0TTXZ/SDDbkPvbnvMA1rr+FOca/6JsQR
/nB4NrIJWNtmgh3VLbxnLAzqasIiwmO5wpytBJ0ngcYz5d+g2Wsu8ebpiSHhmJiO
EQQgvkx7ogeTLDfPKfGra6dIdV8ERaQ1YZxImQZ7PKuRYtvyi4ytVy/Swaj0SBr+
sZBsv2/ZNhuW1kF1iQvTHaupGJ82ZGKrPOnXOHbrStXeRVLLw+1oby+eKv07lIf2
7p9skyjaybuT+ewE2z6FL+/tpLcl+vdBx56QTTHQzB9BjpSa8N5uDNwGQYoCGjER
GjrlvQ0O6b0vgXTJw15oADSEUZFOSCk0mFAdJlr/VBr4QtpVxe3FdTYPNLWSLemc
6oHjDXWM2dJOF67P002StXgbaHTOTNUKzxmtPuT6RcmwRCdj+3wTApPT62pUsauY
5axo69Fj3zYNvXdV5UQIzUonzUWVh8ZFTtri2CUP+8+BfryoxrmcZLCWxi3HUyC4
PSV9zWHLBG8UAfQAPgMIQqtZbXgSkV6PcL2T2ZG5hatJfwMwJPHE8pAtpn5YEszF
l2dV1kgv+QF1Pj9ARQG71UbbTLtfvHfs3aOeFfLqHdAFSPL2xFWpmNFaL3sQF4vO
MccrKILJahsydJvBrg1T/h88C1M6oIHZMeaSwim9kSAaVay6GUJQtFwLZcIXRTpd
15RlJIfnk6XM4BBCp/vqQgFzobS8SLSY9HVDlCKL92WGl9KtamoRP/7ySecR6Ss2
4w2JRxdHvHSTXbCgAt/eXXjv2S6B/73IgwVJbc+DUauzyDjNJ/wj/zMb7kMsE5IN
n41HP7B2BbdJpq9Gn6PYOUjuvkiQ0G8bTaj4yuZKBjPJ2+20JK9xyi/6bIkuLUlN
IYsARprF/HXUeMUHL88m14u7XYfXVozQ18VwWvcS+yN/s7borS4iE0i45wnnh+jv
qh7DmyJXhi3vbF1IFqIbDVbJUuKEHcFjL8UB5aRETp3FIp4m5frt+lVgfWEQIzrh
ibMXldl66TCz1jjFO/XTsYkKOlPl+670xKJNUfBkxarCVyA2v4VB+jCiioevi3oQ
zuBhKK9MLdgGLT8Pqzxkh2/xIIfCO0mXDlzVRvFhULML2Qt3WsTF3mMCGPRZdGCI
ozNn86H98BF+ME4nCQJ98uERfsBlAl4VFKJAu+zaKwvi8OQ5yzW2nhj2iiscBppO
teVQU7Mg8VtxphOqGgKK1c8DN2Qgv5Tcx61aCwqP3iSZUaT6dta++t0+rYuK11ZJ
jTOxe6RA1pMB4HMnnrcDEBgnUTw/zdkiobzaI6bLWo+bp06tYnWKxkMOkRo/5mmv
9u+Mpf4NaHe5oKXLbXuR59KzIcC516gzoDPS/9qoqLe6Z1cQ82IajIFIEtuXEjd+
ksSWn/0kjEixNxAJGLF3kLcRgKLRhcGInkfXLFcj7CY7QPlO2r0EwBUCBqQaROi4
a8f258wBKZZyRuAAq+/6VHZu0eYBO3298WAs/7i+YFZhIqUYABq2QdJZfvj1gwmm
URe8Dd3aoaXvjV4IJxkwFiFLXHqcNBfIpW9OpPzLtqjwFndfodHUbQz1du+dhu7Q
LzBfipnNKRieILN1ErgNYRXr25W+LGB9Vu+O4MKtO9lLy3x4hvnH8UuzJEii3oi2
scewBy+e+GB4bhTAl7oKzngde0szsAIU9Pyg1Qp5SBlMP2ZMETXLXun6FQ9B58eK
iqO32l/SWNKXzhqE86FUx6bcoEPzul1oiosZQTtAPWwHngJMdWePbWPcVarzi4hS
iYiCQarRQd+jNMwv7wgIPrr7yN+jL+NY9gnLoe1LM0ALlg7/qM0FejhXwkJeHGvI
PNaF9JkmW7Z1oFm9QltLZqXSZbHmuTIf2DYjULF7dAMw0ScMNv6I4HpUjanpY7Kz
VjpqZZP3neErrubfwfe9JbvUk45HyPfkRzpNDCRIYsnIwLwYSKgJumNgvCzQ7Iay
TqC/3FZsNGVAO9OS0uHQyGOKmQ+bespbZHe4BqZVapV8KBsG+6T12YhuklzPKE91
Yz4Iz9lkzCYNgQTR/DtGYrmQ/RaYTVXTW9JqHLwjd4d4nsbM5JbSrXtDw0HG2tcW
k764NYQcvOKVOUNaM+qPmFT6TwP+QpdsmDyxojyolzMOPlpxgyJ0YkF2c/g0MS5n
ORTDYkFpR/8mceSM8dIOSvf4KfpsOAGSLC1qpQhV+5V9VWG26k018tSRtAHGetTV
4jaCojsCRy8sJziD23UO1UMACD2R9oxdcgXlQrtpKCdSbt+sEkO+wkS98icP04E3
MhYJhanZ2RPom3Xf5cN/lEyN55oAWoYLMDAC5s76ng8dpARK1nsRH9akySHJjaAA
IRSlYVq73jicI8SfY3PEGkhqjqI4O53jmLoOrINb3fGLJNlqRwoIPSpZa4rGFQPM
2UWAd43CkhnHgsv4oTp4ZNXpN4407ppVPgYe9jxxcArOGMPWlpA1m8tBfXFhwNzc
XkRkNU2Qz+VBm6FzmdhAhYVnKFyuMWN1GFk7tUcDnT+53sYK6RiSnxuSl/PkZu6E
saMnCpAux0CvZA/DXE907cDl3uniowzlPAxG3wbfqwviJ1PP+z6GnZeViiLHnbWz
prK5PFid4a1j8eul56VDFGFIC03+1ylmDwkn9yYFNDrHgJq4lZPiatLxnz+Dh6C0
7utRui2pvKQB0DwYQzYpnNNn8jTz1494Peb9hvwvQgOfo6zGEeYLALtRUamF9M8/
AxUyAOiE/pbIyzNdSJ1K/DR8iYfkcIXP5JeUhyjTH9NU4nXZnjK/YIfHxun96/h1
Ug6FyDhUCn1ZXCJ0sTYgHDA0sC+HSquq5w6PBw3HNDt9jUXUH9zZlVdBkWswGAFZ
ECVvHUGOs5myl1UT96n92OKa54hx+Cv0LEkPBT82A1v6ttFDCjae48YMWyuEDPkX
pvfzurydTzYgO3uu3+hMAmau64nB7/4Lv2iVUbiuaCBlpNsLMZY4JKKO+ZCoBw8G
RPLmQlA+3nfsj4UszKbY+kN/2q5Kt7ZrAIKdbL93OebrXaBRc0qEzrxCu2ZsEnNR
2SB1JSmcaEVLy1SUlqBw9UYmN8V3cYjoAUIz1v9HHQNEJYO/AZUTfK3dn6tv9ico
5RY1sMpKJ52fNavVNILeUMa7owM4WsERa2XMlE9CRiZakszraiEOfXcKjljQENcS
UnnYmW9bOWyrAf6F456+/75ai5No7mMpYMwcsh2aKdIrV+xcL4Mw4ZuSwHvWF7Ac
RDzi9m3oo6epuNa/ocdob+LURSbD3jFqcLB3ZSxkuQUKZxd8TdD3LOCCw5/6lxoR
VC+PetAxGLiykd7ivj7kwcFjTrwRFh9hJ+awn0x06nbLMjaVNz2L4BtNK53u4H87
qgrAtr0+oeoZ+4XMOszPVz7Su0w/DYjR+pveHan8iB9G6UQOMxtkC4XQZejvq11A
zvFp64RXrXMtz9/CpqKz8Wb8OeDb12LF0hZW+cTxoumi04XErDIb2uFombaE8mv1
JLg1TvdsYRZIY69CBzs2GE7vqSzxXLNTlmd5ZUFS7OFhkgrUQRmB96S1Ru5F4iC3
8GYCN0CrrFn7p+E/4PiS4ggP92/oiekO3mD4YVOxXBYGZMd3zifAT7v68V4zzJ9Q
bTS3jdmUFh1zW1O2lCz7oWzFfqtjtndDqIIy+3OiNiD/yj15Oe60/WTYamk2f2hW
gGvoCy0my9VtQMD70OpP50koOMPm+17Qv8r3rJdpTHYkNqcR7wj47ihIz5Nh9PAD
3FWSMtTAjeNZuUlE/KWVTWLXCqrppikfzjw29i10SiXD5QFvWJnJIvm035Gvnfks
CbIBXI8ncH/F1Y9se5eU5EwhfNi3z/ML7/HsjzqmxLAlyTYnw+5oBpmlwbvHR1HX
wvsA74R463Kyf1e7kQ59iXuUNe/9/j7HUoQUUJByDCrTgFKkYtxv3lbinJanCNyt
M1pVI5CyD9Bkz2rRdYTc7W8veM1fOzUKXpu0srn7kmczJcoG3GfWETmLlaujtS26
SRRmyOd7W1dNO0wYUxTUDGGhk3KeAFAJKuF45tldWHoKiF5lteC8znULra/E9XxC
vx3i8NicihkGRD7GktAvIrJmErirn/5sCNDArD4Qlsr/a/j7+xufw6qkvjssL8bX
hogz0TatsVKkhWAnLUmvKWG8JpzZ5i120K6uOvEy2iXq9TIUatPggqtpOMqRxEIo
/Kei61wNleEmfAU1JM1O5+wkw9pPwdbnD7v0AbXDgRqJHNrrGl1zmvBwmD0gcCOB
Y9PIbublOUpK/iHeluaUYY7eJpRtEcaclznnzBpsi6uT6hWQJsMscw3ewYnikfEF
fMu6fH+BpXWvEhRc8dzDtYUwEVX7iEge+T8RXbksPRBVQW2s+Y2pHLP2GohGLrls
c6DJpZ8N0Rym2RMqRLuyySGoV4oma5sU6f9NJIwn+jFrDwgdVXwyf1YPSb8qkBOr
4g2tb+oetKxJk8o8sDs68gF5m0lwYdopbiWrlm38LSmf2rqHkgv+aM9jYJv3ANH8
zq68qSb9QJ2nUbJsQduVdu46W7IFBtAPG2+w3SZ+7gY7sc1+QkaEv/djtQoDZmjr
9L++IICuEUXqVe4f0Jc3ZZru/G2EpZQvt9O531lOjtXP77SS8oNM97jHXHCd1dna
HJZE1NgMiiUjIu8GXM3+hxgLEzoxp/moJvPsWbm/rghXdAnWp3lCaIbAdOIyoFBL
IylY7uH7qSLHLC3EFK6A1aBLh/pQpqmZkaps0Q9y6sDBL9dTzxAbpuJkQEi5vmfS
j9I2iYsrxG6rpuqbMhQe5gX054H8pZPBeCi1EW9NgK/cnCqAOugHI96OPeu4sBXN
c1mF7EEc5d5QPATkY/evcWnAmtyeMixwGTs/+xEwVsMZRWnQnKuScOddrNiGU66r
TB29h+8SOh8XrvoSCrmDqoSPT3emtnNMinpDEDQ82NUGq8TIkVxMwQ1Bp08hj3oa
ngGeSsrIB4PBhyBWRkUEUwfvyEIsv74SauX5FVJwuAynHmx7msciv6DbNovxS3YH
/UMFov2e9/ohTr3mXrWFidyBBQlblaaOh4/rukoIZvGWH1NNd5pZZC5z7N0KjC+o
1rsAUYZHZhm8Thtan4/T0DFTaWxdwIpWR6c+8gDF6td4UpjbIMvsmfvlj0+uS1NF
6bRgGI5vn8m4BTh/Nbvq9lz9HJ7knHTnitmzAkWKUylF1J6iunWzom6Bm+Rdh0DQ
hZeORZjU+sR48N9xjdDQWNaSpOQJIrdCWv5kcqG81MXxdJstNFN5AbgP1ba4N7mG
XtvXeScFECijyu/jd0ZQcGsIG1n5rHzABfdelaguwcdRPSZBjtasvYS6/+gGgrzH
cwrdQnru0CJTrc9tMymNjRFpMCZEIyi6GZBxdGUla/DB8m7ijtqoK6BNKxDZsTsB
r4pbjHNx66toqbhDrnZBF4CaCUQnEwZsZatIsOEAsotlH5a2lF6Pr3dxa+o2dbJZ
hJVGG0kyLtFC+bLVn4OF5FJIuSnWCd78aXo10TLZUWZqJo3I4zwYuwBkVBDIc3Vm
9zIhylPMlzAjIEhDLUeJ4fbmyJ8/Nt8ir1gyVjZ+UFVUS6ojiH3ch5ku90OqLlcb
YmFcJYuVFh83t3Wk2e2knfgdxO9qBxyyQH4ZtAaYRkvl8BWLTqxplE3xol/Wr907
0TgknqPkFxmlTFO9Lkz1+6Xjq920TfhgQ9L+2JPdunr12PR9KfiuQzlWt/8Bv28c
vHPkOGqwGNdpeKnBNKl0pxzLn4AdHoACq6fKxz5Xrx+eyR95IBPcP+V9I26v+IqP
X1Yp46NXCNdKksptdmCoiphkvqscRL/LUnuhzr0fr6hudARhpKwwg7A0/7mLjFx9
uHaAUdIK7cjqbpPNYac/Z7mqOHmTMlDdHQSlNwp15wFebYMvWtEzQrQfSbHL6SU4
o5SzbjZt79QAm7b6tUdcZ/sxIlxjVNV7GyLGTKhhnwY/A4uLZxtTSH/mIIB0REoh
jbT+z9syPXhaqfAeea/vJsLoBSAnWRIAZwj339+H3EjxQ5wfpqq/MkK+QwAQuYzB
VVIP+eTWJwEt1CRHgiapPzP1qvcn5I2SD+9SWfi2GemIPijHs6iiY3H/+rdgGzTE
MypZloqJh1KReTlOF7yRiQ8AX3KBnOlQrQFkqvlXOeEzPuzff4kvaQ/FIgfdAIYR
rA7dBxt9XyuBasdhkO5wFdbM56IUoIgtRxAJ1jXoQgeIlR4Yf2MjlU7d3O/CKOIx
KKIEZw/RyR09z6SmD6XEbSu7vYCM0CrF5k8IjZ6ZO8cZfTDrpq7olP5m3A2uOwUL
UZ/Ae84rtzjR4P1LumNjOfgIQy81PaSb3GLo7lpmKpkkRzQYmjJ4+SGwdMIO6vgR
oAnNAVACBgCg10sPJa0LYgeFGuDW1yIfR2EyUVfwP8OKBAQIFDdkeftaSTYdUBpD
a6XC2QFVUgIYvbP2hQZsdCwN7ysxQn24C/ZqShWHYUbbGzngFa3hqcg5L14ZfLDm
/XdoItdNXWBqI6NNP2SjW3AUco5W05kK7T/MC41VeN0m4wRQupbUPK5w76xoj7An
b1n1v2z78UCuGyKmO20iXs/wF+tnoGX5t79BwvQwHR8KBzXE++lEIEgY0ZIEo8To
YSaKPZvksZvj5Fvuf+d3P2AQLgp2XaF2hx5HOGmLnFAEsTF7sMyweDsN8DWeYOBZ
UEo63h4p8xvz+onF0GbMTi4jlbMBAcVD7daUWhouu3A3K6tNFP+Laqx5Y6rjJdt9
9JK+jZibshRGCSypV8UysbCbfbTDAu3o8AQEguyIaqJrIoK7jijWIw4M/BYk956o
812tqgQRIbjNrGqADZiMMMObETltFnz9tbIMfDiGHi//AnoA21sFvWREOR7WYNm6
Rliu3ecla1wFb702ByYq9DcwU18f0Xzpw7NNBsFNnpPiPI5mOq6F3A70bLSmWShi
MXcBB20LfGdzLkOnvwC7V8EPrF5fswsJJ6sO8rUDfabFD9PIo7udfSSx5BwR8NRr
pQ+DdqSs3GZsikh6+KgdmZuH5n2b87+Vl7sQMgE7R2tECnYkntyK3aCUgakY2XI5
K84RF2saFU8YNSD8q4sesfhMEZ+d4UkiHw72qOMmR4Te5FrKpX57McTIRCXYm17X
qB44RISrWG3HM9dDAh27hYgiCKt6Twu96VdMTcge3ygSDJ2XyepvQk/DRe5lfNMV
0YALYQ/ao4DEQxmzGH3GFu+MIldw9p31rFzpg18mLUhBDcT4492RzGr2rJC5OEsm
VHzggFZ2CDuUha/NmhvyhA0C6L0U1SMVvGqVuXEJn21Doz3v+riCl/7nQGp2bGok
MspylKh6u3M1kpuCBsDjdlZvvtJl8gFOYK95Pb3LBBLJu18RD4nuB5vIfmO6qGTH
PEF8yHfJa0DGmGyp2XI8MVshN68n7sNtM9Du44j+71MDQnFM8WdHO4RC68Z4m5ST
MA18VbEyhoMTg9SDqOSBa9vbI4Hmup9l10ObGsi55B/bI1AaR6iNcroRplOIQ+vj
7Ma0q3B7uhXEyMgpM9cskRjVIpIqcW9PfPPqKHkhUfVBbCCCfU+xD2FDpHhQi4vF
BdLs9Ubn9O9pYqQ6KdrJq4sedRym8/LOwhtAYKsPe68LaWaatvnMD+JxyJmN4/aJ
tn93E+uWx7zRY5uAk8m3LQ8ji4najkKPKh6FW/5A906Pa0eO4GCVGTlaeTs7eBic
eqg2Xx3p+YPt6FiqiYslXC6gb1UTUcklBAzDw6D05okYVR0eoJ4x3KyUIo/emAPb
vrPqHzEKNQjdkeM4jAtis2smebsC6r1760aMtbyzQzjsSi7KcCCL8GPN2UecvV6i
TCcswMueTopHhO5xHrVYO5mCCHF27dhNWad3qjal/eKkyzAhoNTrcxLYO7SANCqo
gvjMLfELP6duL7qEobRx1MEo0Cd4T7Bh1YJbxCoLtDQ+7kAPruw/42XvQrGGV4Og
898I4U1MN3eudw/Sul94quHarb0/Nu/NwiYWt1/ZxyZLqUEDlrfKdMIBtSZOkJDg
sYsQy40+M0r9lTRVUbOrkeo5iW3zZXEmrEwhDD1H1yE7gBUPA4iOyv912Dl0okT1
eOvM7degT21CzJIBMrkcKkDRi6bLIpqDgqN9UmzsmOlaJvqV0TZeI2s7DtQ7Wm1i
GWt723OoMFAQmi0IDzo+oRgPSxvKm5pHTAes49xojydOIHuaMAEOh4+FUoRNiogv
mQmbn4te4MP7oqgVjFVzi0FVQfiTciGwYJ146oaqVyI5epDnptqPUoE66Ldk9y2Q
ZJj27CZuqJ8r/v5Z0+S7c6hm20mdD9mLqE56EoPkbS9x6Ucr1ZCntWQTRuqfFVDG
DKyg0FY7xTrc3rg6Zn61w+fGyq3+IormZRajF1c+eJm7pxwGBbJOxl1kRsROoVd8
zkZIAw/+0PEy87n6lbusbXyT9KPJHOFLFsoNHFgAa5N0kWAMiZtdEM8iEWoBme2k
rT6+4/xH6+10LCWxn0azTV6jAsyiCg/OpMxwiPWfFyhXMe/C4rXC5dm+sgMu7gs7
R+WeTKsghJGKvI9F6GDkysOLxY0yPnneWj19C5nC6DJrkmGb2FvBCecV2jz6w5aT
iKfvu0M9uTvxMEZzksY/vr8MN2Ct+Y2OPjuiRyl536pXFLbCwthi57cfmLbBvam3
U7MJqVD31vxPnNHqaHTFr2tCr3UqIyiMzneX8CrIWWjjPblX9PKehDsf3GtX2hZ9
RG8tSoZjz8/nLguo9PwAK31DRPF+BjbUf5X6oiHkgZYgEGn4Qm1bsZjhcTJObITt
Y00g79MJGX3FK93aM71f1lz9/DiaX9G9oGPOdvmyKxpTxrg4BJJHo/U0rmiNfzdo
dmTS6wG2mfXuANaxTF4YctKbjyJp+T53gBf1W17YcstTeNIrEjNjhTEVXocTUQx7
AwbZv0XLWqe9qR67Twoki7zvcfM7avGh8X1n4UZKebIl8lAj0II5VYO6zhSeCQm9
3HByC8Yrqt/j3gEm+AkyvToNKrMRHSMW965BlaxxQYERTgW45zZkWef7apG412sa
8cd4Wwn5KzHMZq09gW7u/SID63mI6SeCOrsQjey2m0fuVgFjooqKzck2d/uXhAO2
kbAkxX6mocTw1ZmK+v9QKrf1VUyrlSMtNcoICAtkwozxkKCSPv8sh25tsAtE/lY8
EAPyJ1mcTzP87NnekCEX1MoKzuTevBMYRrBmcSj3NZ2araWPkj1DClY/Moika869
NZkSE1+1Z4Y73bFpte4udcS+OJzrAZz8TwXEwPz38lchw5FzcsuEvIf6cMUZUDgh
E896dOKuUEEPzK3fk93RxC4Bsq2g2RZzPM1o5eGl3fAxfg/LjupNlmC5M71gMb3P
Ch0b04YfecNJV5+tZpxxKUnR9NETqqraSjO8ku6XWCpDSvICJ5P3teybumxdVCR/
2MC2DPynIMItcjMGQTA2o1NDoYfoiAFx+OAKSA+hPrCEAOjTdT8XVJHRxC0MQSGX
5f319RxuU+GHoofL101KLUpCm+/f6QEsXNk/dPzbcGldzVmvwCqZhFxrE04nR6wF
LBPdEARVtMo8nDU7fhaNl5CAjlricwishoXE9Tz2e+flKDOyHfwX3PbpVFLA/jLu
pGiNrLfrDj9DqYSoGVV0g/tYl3v5qga+dEB2fQJM6w2898Ylha9fDu7ldR55jWrv
oIrDSrFURFy3JiHr8H/XIFS/aZ+Z0+Y8HNmRzwLC+qRtJZ9hxhXkseZvboNw6YL7
g24Lklv3P9wCjx1fqFYhP2YtGXPcqcIJv8G9P9som/bJomcaPNTCO/1HZD94XPwo
jU14fqas5sWNRTihVoqNIZNJlYlmXMXU3LD+SukuzdUppAsWo4Pjx//xug3k0Y6/
r9ib7HK7onbXbqDH1rRz+QDr4Y3Zsi6Fo8aXd6pWxFZ7jdVXoqMUfLVVs2nfGZwk
ZR7MEqyzHZdUo8gzRwagmwiKb2zN3i+ybJJLLf1K0aYIhyL15yvJUE01BnMODxlZ
IlCGlnzSb9K/lpuyfwvo55B3r/tOzQ+owo4cJKSRBiUNI8mNpSTg1b3a82Xc1Njf
1DDnaOm5HPxiX9YDm60AgMXPUh5qkUBWUog/C5dtW+/O2Z1c9NwqvPiFMJJnFPWk
1Me9pkGHLf1Tfdpxk9xdX4e1f7S5DjzyvzuppuZykHwyk/5a/D30w0CR3QHj5HDr
+9LKNSf8cdQmg9EM4MXr7kFDHZE6KaPQ5HS+HaKILqvYUqEpYSUGJmhuIvndqSzS
vRhbhYDn6PvheVLBUik/7+dCjZOrz2rU65ovpFR5OZ8zl+ZNE2uSOUW6Fv1P6yV2
IRfLE0eMDht+Xhuoil5G3tAOtUqgYa3zKgSxoVYocx2sc/R36OMAbfX3muoDR1zK
c+iyKF+cXj37mJyzpjIiAg7NTVsN3yxBa/a55UUZ6u7mcR45lDSpn0ZZjOfBcmnk
WHODamXRQkD1BLGmKsrgDy7PL9Ipui9QTWfAA3kjswSIKFQ0p3rw9DlMLzzZODcS
peQXP30vYZIonCadXCqcZK/RDJ66fERsQ2LnIFF6YRAovYD2PvTVPsE51oeo6/9p
w+axRjAnLhfRnAobEKt4ULecFt4WG0Pwgj1b8DtoQrNcTju40PFrnS8hQKbN9F6V
PxI8AzECArh/SF00iSdTRNmN/eYDQZfjiPIwRzxpi0wpujK9UDfPEK9RL+Oi7J/l
bBCFwscknWc60+lP837F1bZ0MG9jVrnbGNbeCjhPqa38GVUdBDxE+QjTRlzPwRWF
VS6U/IXrFmK05TlVgYbRUXaOYxOT0FGgnwU0F81j1n13lhyb41kfAB/2ywzcBU3J
Z+wZZDVseeKaEOrRAjUBzjVMmH5sBwDG/YHVg+WwzLbJviYK7EIIBmBcUVKECkSl
8wG9ZEwYfTP3ACEiZYqBCVNiehtWavSw9ryKgIx8fAQq4SaTlcky00fhfjMJOyag
NLQ2Izfx+P/p2IGuVJ7vA5Eh7UQWB1jyDkA/172bCTrk5k9zO4ISsIr4Wcr+b3fI
nV/I9Xe9o9VL3oo8kv0lFcY3Z29y00sHjnxjxNbkv0j2bzW+lLYlOknEStn+S+vN
TseZcB+C8YqWtLycwVLB9oFK+Pi3g3ZARRmeoZEXCOTNGpXlmpA3u050e1pTYDOl
UUh2xQa/5QmiB4EjIE0YNS+iXOCEau1oSrMV9tfqEo6gTf+gN1BpTHOMcZDgwjQW
eOOxYADySHQQENJ2Zf9BnR2ZOTKmYv0HaoCRhXFU5VGpWYztpTsIgESnjSWTX+ki
fl2XIYXeIuNGYh0i5KHIj50C5ixKh3sZC8bSImbGruXEwn/WwNR1vAoGsq1knopJ
cPyhTCmnlkWnYHeYHOuytocqkbNXqVH3ceIxWhL2PTxjfxonVLGKLGmMalFALKSS
WMcma8KRrMBqjaJa4A6SCaid7DFlxbG+pcwr2eiovnLC1DgmqKiVCG5ghH8Xu/DN
3yJ2VBMXWI+KdB+MhNL+cMC/Txqm1hQgVa0bAqOyq8q5o6G3YJEs5vrwyOFe2RnQ
UcjLZZPz9a/S2+ixDT0D+P3KOivCSTkyhGV0qYClU0ZH5k0Su52dtJfyHvlwR6RM
P7Zs1ut/osFVpXtQDeOx+QUDmC433IW54o/gBp1qaSa+WKNBR0i/K1nqwiIRomSH
lO9PrDWthKKHGvecQKI71tOlLcj5RHdi9knzlffJW8ZeaWR2q2IBTMFlPxIjNvBy
9g9S86UXR34qWXuMCoS5BO40ghcnLwWG3KjKaRK4oKXFXmOejHjWXftGf4eSEM3l
XqdIQ7GSPdgUJ5TuFncwPSM/jF9hYfErINiaCmduPeNA75wGP7r8r7lDTionVtuO
b5CwkF2H8mKClQ5WOMW3pmGyvf2Hu85tKKORyCTQXS+xYCNWa6C5Y7Kfw4z9+gQV
2N3bn46WjMyKb2j6ETmjfX2jQ9Zg/E+4apx8NWvtcxfSKKsAfQXkIS0/QtLD3uYl
44/NThdlDPCZ++FF1hwFDLgc+4TRlWPWQkU1UgvyiL2ilMFni6ga3vOv4PyZ9EYI
kfuqzrSsp0nQEJ7YLcThPCjsHR8CnT4SYxwXKNiKvWpU0P6y6FpConwsaUopRwuD
qQI/OS900ONNqsdTR5siUObsWd6fMDb4CY7xO98vDfQO8UhndiTKAMFmzMVtFwme
LdO8wUjH0Q3XEadkDxL+gFAJuAYG6+PfJ1RTTu2JW79iGBPoCvipfJ3sHmQDnFHH
+hfSpKEGvhELPQZuJcYoXqxt7TIKldU4sfH9NERk//HdOa765/oPtTq1gzsNDaKM
rxItvOGGONeLx6B0/fKHn6E4TJl0pqdQoYGmNLqrNKaGpubE3NIQhg1HUaKOrjtp
T61kehUOUxgT9NexYCCFXGSm6T7xC1UUwb3LxBiqtj24wO9TlvVNMjVosCeaYunw
iIAbbJcNZzP98PjWNh7xnbYvE6f9ELebWSqPIh3kVsdDgQVOLnwX4XIupEW8xaaU
xJjdOms9irwx3azAu0dDFHRH+kiErlCiAOXgjK8Od1zI9zjdyb3MKSGxlrcs8Tup
f+7DApxGIKMVLOu6v0KpGiT8gZ0tTeh28X68GYgrODJ252szV1mCTdW50xB/LDN7
9e4SXo9op/cr8XxNaIT0De6KGbpJkt0qVOnxfHOwecWsnZO1oY61YTQFTFLHJmGc
p5mDOSqpfw/K2wM2zpASXJ/zt3F+MTekwzuOQABjPDx7450vtNfK1PNIaNwQIgxH
zThw89otmicfe8TlKv4tOFNL/I+7mahrOI7gvve9YaEIXjvpkXC3vMK8Hb2F7F6j
huWnanhIxufOpnY9GAmfBdHtZCRBWVy/BjhiByGJTQlSyyNM7fJgcuDPiNo0ljLA
CWTqCA4p7zpgDarvQOy3a/LAkyRQoj81Ym1tGKBnG4TQHMJ5QgX8WRCtW4twzdBe
92tGBssWAbdcnwKz7+z7H2yRB4ssMIAFHPjGVja4EryDSYaHeJ3taD/Mls/nNh8l
h0cGxwcLkKvgBCzHoM6Zyrv/OmCN/0b981y25RyCnBzff7Kw5k2A/+xQrd3C437s
l0zDkNcxeCHNXCqwsu1fku3LXOSA/5RGQ0T3VDcIfrSLDlKnH1EhrhwjQXkwhbqJ
B9zV/QKEh6zAJxTR0jJIKZQOeRlbzl7UUDCkbD5Ew9mFONjt8lOpr3reP/N5ju+p
jZgIECRug7jW5iBzFzXfCYzFX4pbsydCnmpIR8LBeMw2wfXM9GKfAEN2BJJe+fQE
lNJs6I1+yTbWXBFlFDeBFE1BA4gGGFYd5jhsZwjBImGRcEBUDhhllVNKD/LOcqX3
OiG4KKHKXBjgsV3pxjSo4R49CJ8h2Uhyiqnp4APPgf9V9Q/6cwEfyBPoiL2XMEq/
JsvjKgkqNy88YQeEXLuu1crKrZVYIkqUqPp9cXiVFC55h9kULnSlb7xaDkjyENlD
R/FzEjd3c6kA42n6gD4WX1e+FZ0SDJ17a3QwQTeBvkfgKUUBQVHeaeyO3k0+s2u8
KM0syR+Rl9t53DoPRwzTkNTq6sSlnYVT2gLtTgbvUpHcpPsKU2GGXLgaAFot7rrP
TTSLLXRjnvdxcH9BaUYG8BKY+ahcrZ9rwK/cvU4L+rZJIO4iS0jZ2MtMNcf3TxvF
gRLhDbfu1dSfQtkpoPhXBELMv4d2GkCSHvoUe5mS/1dcL9vSh77Hz5BQ4xX1In/1
8P8OTDIy/RFDSCHX595Ye3iSB7O7QPcFwM/9R+i6AA0wTNX3W5aU/iWFOJznUvd5
vWUeoGcY0ieUYgW+evl5jtfPgz9mc8WsZX/mHsYGZX+DdumMGZfyHZPBABxwhE9d
VSk6KP15+Tg3agXAHNbSCm5X4NKr8K5U5NSd+rke9M8UtSXNH4OzTt86+V+G781y
+2vT40pIvCtrWQza3GvawWTfeZIVKkdPSu0WLaRy0DEf+XL25KYg9Jjztnafci5H
jZP27OLpF1Y5nxQiSW7dOfbGS2y2kqWIEVm7rM2XS9nJSCtqtJAvaR6V/cuzrcei
b67ne8gVreLVJbctjR266l0lNA+nAo/ghW+Uc6KxnN0sWOtkvYTf/QiMEf0T9EvK
OFuteyF8ERJ1ZcQlhIAF8dV9dib+eNTnoLhTL0gzmHrPAnivhhew3KPJ95DU3XrI
cInqAbiYvAXhEqSLKep+O1f3Uvy1wKP0HFOVoOpRPtydf5zZzSuylaePzoMfUJty
gW0nvrYLCYIRh0RWa0TuNLe4yIXiCWud83jeStwCPVoN4FQquEpPYe6Xnv5ar6wD
0RdlTufvttyHaSxBehX8H2jpeA//g5u0vUQOgm7lpgNyeZd3Am6iPoFFVqa5JTYv
iUIa4Df9EhR05LvvZjXKtkz2VS8dF5Y1T2Y/o2WCGOJs22TFaNAXNQxxdfBupL6Q
TZ4OvAYnd2p9nP77Qt91MwdkHNiWB+x1IhYjuOyBZdTnKfhQHZZ7kCkpVdjilC1+
yRAgLeSePX7sC/JItH6h9rpJPq0sQqSbezA1cWlj5gVUv02ntbOuaAqmCcBhqroN
M9LsStTGZazgWxA94GK8ME+9uNfUh7phs+grzrn2sDijK9vh7BVoP7nnFajnHo3+
dOgfbR7JI95I0s5N9ia3lgz1AwBUhz0mS9ULelak15JHZizmY1NbIf6TBCM0Co1E
rrf2Jqtg28EjeIeEYXmXDjbExN7YzdiwORGOYLdkI8o8J709/C9h/mR48qJw2MEQ
a2ma5EfhNahcTPRyzaJVupXrUq3v0E5mjNzG/GEA3V5Dqa/zmUyJohVNxLRf3zT9
fdEa1SkRC8Lx76ni6YAA8UATgN6VV/PbJ0MPkk46lJSLQIA7ZzZWlQIX7KseFTtn
4aIOdyF1sqar06VzfimMYTpO8RU9G7aDfjmhruaL7MGqkCwPZYqauFCT/i5ZSTXh
rJSTSsp/KMS33qmwZlX85PxeqxmMqq/Myt+IXd1ZYCxoCwmwcoH5vu4oMj9d+4n0
SgqRgQPt0v73juYjrGSLcgiNFxUUjNENFBfwlWVcg8veUs12dFOfoFnptpm6afOE
aKzMGd1D6Aq5IcKKIXOPqI3ViaHM84GDffBFO00Y8BH1yimOo4qX/TAOJpymvjFB
jM3/H8nBs/CKtXZUX762bGymTBNbnxILf/y8Yv1gYIXryyzW4H8pVkZSCF6K3oMq
w5AC15on8AiPJriPL7DRwC5I4il2JYjmEj46g6ilPqk3GBYidb9TqfHAuFx3FxRA
1JROOgH36/LMMg07IcD22XdUVdxIfDsG/kn5A2Nmb5dA6vVOOkN29ZgX0qzU4h92
9gL5hNFbvFb3+X7jkUbO8HtsjWtT81p6r0c3m/gUp2djj+/4itJ7bYhAcRgf0eSQ
w3hi06vvLNHrsXuebsysIGzhgfn4CJeSXbhi1q/llIpX0sGONl5+XST+1T+9Wmgw
g2KMhpDxMxLpWEtmdi8tJBZ1JC5i1WrLiMjPRW4ZQOWAZz+KxlQH9gzEnHKH2IfB
gg/lbHH/gzme66yRLuDV0eJ/XlLWrSIup1erioNxwVxsEaJlynM744bEvBlfRECX
pLh0ZZNdDkbGJB48JY6Ja7S3WyhuRaCEX2Nwm3e/1mC7Te7Cdghmo+ijogmSMFK8
FyIuVdP7+xVl8nPIZb7LSh4O98qzZRjfV5YUNY2C391bUKKUbQeDJpUOQjOPuKNp
vSuz8snCQaMmy8/zr/PK7ajZZvFx133wdhe7IfhBSOO3Tq/BBfS+1rM7pqMHBZC1
Kc/JEOO3eleaWwTXIrSaqUDnPI2bd+zb9QBy+Azy4eKQ35jmh1BLFAUgnxKwMZL0
50ZqFtEys1u8fsYv9f38ZYzXX/QQ56tkfzn+uQSzeHhq1Qq9SYOgFEj/sTh56UY8
JjyfmQBdJ0K74ZGsP9HuvjaGWmGij7E16xSRvPCK8hi36ByGaw9fgwz4EANcdQpT
lm6aNQeROfx7hyrN1j93xrJBn9oubhK5HrdK0jjb2iE4aI8xICLi0xBfVBY5Z0kH
/ErQyqMQL0H9SQ70498+ilZId8nHzXMleG4JjKI7U5V23pWk1cDccpA9TaJ4VkY/
Omz1a8cnopjRuYlMjS3zGpPkqFl/rNwmPnuMmts87aiMJ6gr9BESRERFZ3oEHysL
paDtG60f5is3QjoFxuh2Nq+OnDO5tBQqjPN4MNVA5kbNJxu8mV5Ws4L9ZhVEbsNh
oeX3qHxWV5NiOOAhOuZipU98xKPeOSVCf4FMfVFyv0mrhY7kW1jw7/GG19zOUS3r
RMbazxw8wdBehtWEpyEk2VXneqmZtuioIOyxM6C1XGth2LJHigBiK9L75XRhDAeN
iu9XZg9m9wJ3XSrGdno6fnaSlj5K2NkrJMff/NVxDtdGPoLDCeWaHcofunhT0rMj
jqWwR4tn6PM3XIJ42ZdNH1aJXCIA/tpPK2NJMo+5CKdBY10KZAlSIVYbaFfaJIC0
tYrZm9E36uFjh/OB3HaxMEL57zsQVrQFYzPWgQx33oWo0vJi36jethSXEx1iUwKU
rkGxnzT2E/LJqaf7Vr68DwvE0jv5rR7IzLmoDGU9Db45Y8J9p09N8VBH+PAGlM8Q
GqVcY1lgfwHS5JS6tjsUaQbQug1E0G4PCXgsAcGbkEpVGuyHOn8pgY5+o7MSzKHX
7DUIagHK1m4zDNuQX+vXs0Qkhft5+AhVhNoKnC+/oC8ijX5/ew24QkTQxGYzMjWn
NiizddZ1COvBhJ7hESvIbqkbBThPQSa+CT2tuihpqnKd6WQJG9Kg0vKy4K3aNiHT
iWcNRk+mQ40xbDZo6Pt34SHJGIoTWZ9FCvrty8aV+fMZPSsd06pNLLG4rdr40VAY
s+3GL08SNQMGpee2c6buQqv7R6Xgu5rcFBz9pBD6qM1zaS+Fps/8ToxU6HHo+Obd
feL6UseWs/nge1Tux/qFUYZcXyfNKi2uXx7gfg4H+5XYhp4xIU/pM68ggfW4/JPY
x2q11jVKv6u0Yof95YNBUZ3cY78vw0tQ2fvtBl94FqpePzHuSW4Aibx7zPI7ypMs
pStSZs+s61cmhQ3G/dfDYlz8bbGHlDwH1/tRE9OCqEqNX2i3NmeRomH5czBSxgTb
2if5P+fPd/1T9BqJL5Js3rqXjFt/m6uuFkMSGH+M79GTDc+o3MeaI/doGtxctj7Y
A8dUYftJrWK6KfLxjkYH8MezF/kbKkIbc0u4qJxY4m41RHbW2r2JjSP7Mq8XfEbv
+28syMrz1T7Re9SnCEdOtMCgSU/y+ZCc9b9RbmY1S+q/4fAiOtyonNSW+2bQgD5/
cFUokUJYExx7PcgJMXmzQeJx1mbFlevXdxfw3b3P3hIWb9Qd3gVqICNpdIazKjgN
v/DQ75XUC410TmXjIxRy3Oq8c9V7JL8YhQRPbOOKiO/7FxhP/Z3vZkTNBome0dnT
imr79C/LD91tyClyDw+dkStaw8Go1q86MOwuru9lbjh0h1PVZXZ1o7Lnhvw5W11/
TnUFkUVfZbnJP9euYPRUA8MmUcBg6Qf5KhHRHtpW9CaeCI25k/xAziElGq6GBk25
E/P57YFJA/SBoVDe+ZAXn3H373SWQn8eVcWi5ZD505I4rD9268h1f9F+u1Wo4rQ5
dvg50ht9MW85p11we9qTjWuNsYtLyv/zb9RHKMTwnR92XQUNtiKeaP2d62dpU0zB
k3Zy8YEN7FE4zfZoX3UTlt1rkT0atYLJJpSh2sq4Mi4adlHfoeAiB4JQET/7Vv1O
3NI3igup37JEpl6roSnxt6/mJ1I4AWV32zLCnFgA4yVWVbuVdZC7DXpoYAt2JEqE
cLyOyi5QR5Tw98D7qBDWqCSz5McIELWN+53HpD4K1JP+WC7LMfvvEZHQ2qL5cwE0
8k0jyOf5KCBUVuF/A733wotw2u7t2O6HChphwXZ/4co+tcFnJqrAEwNN+pWi4CkA
rtB8PIvhRs4V9TtWSiuPuXnVQbuo+ds1C31kjcf4Dl7JEbOgn4aEaBWHLAnvFFIj
WJHFo0EeA2kaD55v4ifqTiBwhJkZOl4D9hsoQbwPYGF4reocTRl4IjuyMA5p2zVx
pqVAxJuxGTIJRVLMjpuK8tvsISvehrMHfs0oc9Ae6OXYFESCUCl1k8qQ/7Wyl5XG
QqFR/35ORbYNYHDkedaxRIKhy199+1E29cBRLf2U428LufZUwiYsF/3DIMHVMLsU
4Fk7g9W/nRgzDiXCkaA5tWZHQhpvGipkgjmKQm6efRJIO5eh5SYy8GrJR8miMJCY
ynO5MJPiIifL7hCdyAXV14lPsG+XZlp23+Yhti5PkPbY+mstQ+c/Y5iMS3DdbscL
yDJALjq/x1ADzBlOoOe3aN+EXWRKsquqHAnIeQDa9OLbOHXOJdyZaHwUogPHLqlL
5aAd3ljC95sv0xz5tV/U84R7boAtRSUujYNdAXYqePZV3TWI7fW4PpK2zmpwuDBg
JDGeu9nXCicCkj6N8/94ypVaopKE2d1Ed6w6qC92fyv9z8Nunu2eMTGtDqiY092d
Hq0ZwFmkNroC7ZXu+0/4tBsZTZJ+vOkhouWym0ndaTaU5Al/tWQmOhY8zvWHVAu9
wqb4jf2tMc2wMlBG/jU+5d6t6OQHfMNK2U20jRcTjGKQJr+fUbCZ4bEI4sjsC551
DytZvOfYgkCPkzymLm0qmNhHe97hFUe5/YM6i/6s+IHa6nMqDBCl5mHW42iUigDo
KAE+mr0BRGYTRZcwK35ee16D6HgQ4NYKNvD3xTlIkNK7qqXCwHsj4k5vRZUoXfJi
8KGtDbDIFKc4/y/Yp0ViiT0ZL1QuiPHaDZ5RBtGLLvOUW666bOiYMFe4b2EXRQh/
uceAWiBMWWZuzZV5Fx5/LAozpcITbR2XLWETzGD7BqgfRy+Bvv+/d1OtvXn8xsP7
cCs/Rx6ZuL7bd29wfGxTFNxkq3rfm+56nPhs/jL+Y3G5NC2tmTKhvRNuOphOpuKi
ryZN1LpWAUcvEpfpTiK9f5fAkgtwEZIAEzmg3sWVA5Kzkxa64q08i6ig3pnvLr1/
gpylPyjLyvX1JSIvvFaT4eL+f9UZCy6aQLjCKbYC6HaE397x0HBZ+HcNHVi/nOWD
pM3Bn7XUMT9GXRpS+8xCsW94a6/cI3EhBKUT5/1kNYjs2iUFhReUly72Q4NdGMFZ
r+o4c4IL1qH0tsNe8kQOhOqqeUQEs7Qx96SN84MZQIu/v3Qozfg0+udDBRILrOgv
/YGYuQVfoy3JICq468JX06w8kzayEyJIgnbiJe2pLBMZsrxG1fCS6FENGXzQgZfj
DDhqGQ6CGhRDirSh9waXvxdDTv7/S0Xwq/yRGUufZpBSM6+XQsUirv0G0lELqmHS
onPumJI+Vh6Nr+9jSr+faec8mLfAMk25FeiP9SUopJJYnyRQn8FiG60AolYSstyG
XZLjn9V5H11SqRs/wpNSnaSxm+bYJNn6/n7QO8JWw6qNlieGrW4agXn01hsqqRTs
6siqFfZR42ZSXv3YP+fbEIHwXBkSa1xmq7Dj7wElwjA5yhPEbjcQw7BOZQvL5yFG
YqhZ04IErhiFJqjz7hBdoG7AaI4fztrpIb9TZKdz2N8DtBJzaPyKxOBWnLIGWuHP
mPKvUFDItLtkyQVde8CfGUc3DqeJHJafNsRg+EbWwloTpPh4v6ZAcds5qY/G7MsJ
hfkKOVJvwnZRdqABVHirqQeJbUfVoJ2Ef89cJpryt8Zq3t7V9E9gYDg9KMRvwo7D
QE9ou8tVrng41ZWw4bpC3CaqxVl7qWN+QS1eKee3YMcq3lnwb/SVts4lVyMG6NMO
tIzSc7Frte0uvky/ce5k2K1Suqel2AXzGhCWUkUJx12Ekdssn5Q5ZL0Nyjs3bsqg
ZdygEtm30F5+t0puq107b9mK81JncVxcWRTgZiA0PVY56XU9YIW4LOTPwBDVMIAO
QDJWfy2cc5vSULebMYBMOFSYeaOk9f6an1GiLKZvnOu+WZA59VIYTcoYhWv7OV1n
bNB5YPyb2P7ksvDu6nTosz53b2L//SqkbBzFwg9PgUKfIhQAbHRLCvL/ODRmZ4jP
To4Gf30PwzkInvDkciKkby5S6GECUIdXiiptX4xCCT46G3WAlKO/U/fchZSxGzCO
btz8klY1H3f+z3nvj8rwW6dUX4w3YroYFTz3yQER4ygA8n3wBrmI2B7jljTHIKz5
c2waGB25LNDvbhfCsdqlBN7EPrtuJAPuGun+KV5IscphCMqkdz8zsJ94/JiD/onH
j2w9Pk/eDFtCzxGLSeQvPffbqI/jGTAfLwAzepoPtK7n4am8PHpZLRjAMYSRCFCM
Ye05Y3VHHrI8hZmkulnAH/OOwqsC8YmkDzVRot5p8ssAHLch/EQ1HEI4mNIzpeF1
nxJWMpTRxVeF9ql5O1N9ckxFGuil4PftJg+69sw03XAqfq/gSxSntZHa6Sb73PAG
ARKQY+4gAWbYWeKP5lynxc85rXNu6v6TcxUR3QGJv54h8ca9VzwPhmtuSC5xuK9o
kB3C55l+Z8e41c5IxebtmAGdF6qVcyuZ4iZJy2jeJPcf8VvGwlJAwDvWzjHpKnd/
QL85ganVefMpn7D8wX8aofiUB+qEYCR1B7RidLVdaFAgT6MLeBqdz/GB6qVNZr4q
6C6V87o06cucCuzjA5jJsxAuIn17Ve6mN81sl7jM1CxIbcfHzW5fq5OW1fEiu5X/
mSYJnxRj3FAlO1DNcxxBaN6MHgfOHYE07vKvnc0ET2KlRPhl7ljFR0/mlhmX47mz
ghEwjdYgY4cc0GkiyBAOK1s+7j5Jc8jR0YKJH+nbp5deP53Ghqrb9w1TTHLghHSw
HyEFIH0FcWJ62J/qmWjKWV3VcLGRNId197npFKDOXQLSw+fNxdFct/Ij5iiPOBET
ltEon6kHvLsLhOrZURkaMnSmGYp7nKR3TNjsk0uPUXnz1ZUrBa3vaChyxZ1IyTcE
3wjPRt3q09KcU2zhVkihVZ7WZune5rMJ914UIFqHqfUeXJRPKSbdK/GFYHRpGSAy
+jAt9RQR0iPCroT2J14sG76einJZrdBm21xRpsoG3z3+jB7LQTp7uKcvK8V6DqK/
6upmn1adIOn3SEDSHEryi4+5+jBXfdE4G92CQlDglzGeDn0RZMumEy5NWatlnwIY
HoOsTK4j5W6BEMPfGmAqnTpIfUHKLEUu1kkzkQx6zXO7J5WUM1tQkQeogDxInKsM
ARB+4b16lym9UQjnXror7IVVjY7dTP2UPaIp5wZ82xFecoC6hhXyqw5v5amevq0d
VNHxcXhSJpJwZsH2rkt6BwmMmctwMHwfGFLk24JyuaEuCZVAtzvAZJJhYePW5TfD
pNUZOz0jWsAkNDf15JKdgwBr3Flcbe00s12bywjD4csfgnlTRxEiHFcBv6JgLOZI
CTot4EB45SmgYK6mws2TcrvK/UAcIfWjRw21BvSnAADRRCgAh8vQfb8sHkPOepwm
jBeSGmOrzwiVv6cNKukcWLff4hitxwpRiFizI9MFIJibOp9WdyMObXGlleLj59WV
qomE8PnhN5NVG8JGFBkpETdo/CQM0SyY4OnZhP/PqnuG1ijiIrRIebUSn0HvwG9g
N7tdhdWi8yjMkJa7nEtRYUB7WMMV6jEHOWx0tOe/R1Vg/Ew686Arn6RwVqPZi2td
aYmCCSEEgqTEeZlddpcDdieBI1L90CHbj4Dx5vwmdMy9nv7cesdwIDWG9+tVm7AF
9mk0j8ptpu2csZRudDPlI/1KeIEGuEGpYGpdCLYXTTmVsOwrnQQOm++/YtTc75FE
gBjYUeoMcPTC1YiXg3UDhbyvAobqKtdMZ2Vgdwpato4dI4TlwYkT4esw1K4UfajG
RbuoTV/XQfv7gn9RKtc7fDktRpInG7xlWZRhPtItUWnVs6/FgGRxiibYhOFbER1Z
hvQrl3pXSiG0HVURoUa6gdyvjZ9vIgiLgu12K8wtrEOxhMOQWajSY8yiR5ybuT75
0Cll5j2lKnDXjjlFd/Cs/DJuFyACjiYItQ2khOK3rvYaYK1X9c8N3LG7hnxf/xLZ
S5g1A0dk4Qob3JKo9ygQZ6w6j9vuJ528n15/nRwj6lHkL3YAcZ4J/UjM+slARIZ1
/QIi5n94k6Jok4NePxJD9I/JbHPm5+aKcingHbqsJ1wynfBCgYW6oeR1bUjVX6oG
Ot1zo139oPlOfPb8enw0mcZZ9tBc0ef7/GIzdM4Q4ZGiDstIS300Ia+eu3IPAiXv
PVH+sEBaKYQRGzxG6Lm8VPe/g9RSCDLurriMNVPfBeVN7U0GNvliFsC8svArPN+v
a+y9c4v2SaClscUxwUeSE60pWUln83vVjwonritke2VQMErt+JRzgtzclP0/eRcf
Az3EXiczNIkCBwvkcRiZVX8s7+m4XskwFE6ILYJUa3TwWXlKPSO98GMDJ0OvHNn2
2O9uX0hgG2baQcIrx7mHdutv6QpBC7Csnr7PTArtTzz+LUtEPNIJrcf96WmjNZGt
ATzrdKFeBje8sc+M90VIzWqTGy+QRws5iEklrk1JExhosjkv55+6m5k8FjDVXU38
V4vFUR/4iBCJgT4K74kvo4On7ihU8imeX7DThW+19bUMSP+B7H4KrCQsP67Xc/KD
l5um4I57Drw0u51C89dpfR/IN2kfvt606vX/chNVO9rXpfgoVvWQfo+XDOXYlQHu
vXjSfFabOt71rOIWiz1Ees70PhjD/qLsU8vf+K7aY/iSjO+KLeJcthlWOSO/uBxE
KorP+CNCEc/j2iAp6auPpThqOj5CS4WPLWVq2VU1XIeLIFrOeqfLsj1Crq2Vl8y1
UbCniIeP3xJm+XUIHtNLn3bfGuMXOoyhe6pBF2Qr9ngQfnshHyTqDkmO/l3iEBVM
YpX/Ko6OywCz2FSe0Ptiw1/b4R81NleMJ7GLYxquN564WDxlML9OF1SkHdeJH/co
xVqoI17fXMZJExIcmLoAS869nDlWPG/JiOKK1T98vGRDFEAq66J1OnKlbuLTzSja
ZjCQiGHaHKbaSf+G2IXAAweNdQZW+PflzBmJRRvZ+B3nah5p3JBJpyUGH3T4eI6p
9ZffMvg/N9Ccu/W6EcmJOYVFhzGQFC9mPNm7g/lfYIfwGOIPaTgVQbl1INda7nnu
Orjz8sSjL5eZAeKEGa5shXM9jeQVxj0f8/jEnbs2TNL6ycf9ksCHpHP3ZRInldyL
8Xs/Iit1+PHR0jlNJrGeefCd3ORAqw4noOYfQWwspD+Kg/8/UM3FiHdweMER0/Rw
XE0U+76wpIpBBrdZQPTo7KA1sMwOBDKtfP/5NIN+6j0PVt7/eGHcNPb7R0ZXpnkC
5fDBJv9M3cFoPlI8y9LhvtSGsaTW+tOMyvAvHzLrA/3X+N3P45B4glT8w6CSRCTv
wTPvEsl/UuMoDK5X/2ltRIQhGsCtDlwViux/ZFdxcLXykRkEioBBy+kmZeS/sAND
4q8QIGvPKP/20l7uOxN9l7ZG6LBmimOvQ9mxJaMg6UE5cHVX3ueEkj0FHcf6TzWW
wTzFQiYFWTPBK0VNTr5hQ0QEfG5AL3E8N3TCcLGLNYcn8TCGh4K9FGec5dl8hUEc
ld2CNPHWKBSWnKyCZM7rxfY/9smJEkwKQpyXt5a6lMnkl5XWkQZakOJxmg5e385h
rNYk0SuOTi11ffQoPwDh82/XmJ/zlUzUWA1dFhDfQo0Qa7TnvZRCw0z3316nM9/Q
PwEsa0sC+REZ/rdL2iRw8WI3s+SVt5xjazG4QQ78uh7lyikx/EaIaxpDLW/M1RhH
8Yf/G8uCc2sQ0TXAA4Yvj45mOlgN+/N/3NxgeI9h6ANIe9FBoDG3WzhokPLz3kpk
Q1n3pAy/scxGepiYwLvKDqmg157+h9MaHNFXlfynEUytcKalg+R5AXkih6E4R5um
/69hY9XEG7dfMOFpCy2lL61g2o6u+T9Np8EyueDaISkurb39eoTkl76W4lsFlF6q
NFgSFEg/9J87HlE7EVaCVx9sWCoHpHze59r9lj/H6QAPnqeOxo/KOzlUMVkSqXA4
PTbsa3O1Q07Wm8Z/kJiJYoKAQ/cqnEN2b+RWlwmVKFSiJW/BipSFCgp9WDc/Lc6K
6faW0grym7MeT8b4RPPawTKzUfx1l0ywRkibHiykwPK45RS4XR8xsvhHX38VsP7F
4UQfDAM/MK3OUs9DDuYDCKDE/qy/HQHnwiQa3gYwwGsuSNh+yEPH/fz4xkZokeg3
BtBRF3+rY6uMS3dYbH/+ffKyj5xz3jPEZZT86UoI/yj0xbQ7RK6Z4uNjU8JGlTcm
Z793Ewm2x55hK2U4aMsmb+afrYYfnhHji6FtpTpaFAMQl9HVIAskkFqS7v6fyzUr
Jh9TXVuasWvZ1isK74Kvj2+EN4UQohehNQXy6nQXIbJc1v52JVZwERzpummjW+Sa
w+9Zh1ZKL5yglkifLV+Gh9PPlyXGBwLLQlosC5VbJ8bke2RGiwN3VUpewB9Hwe39
OZ/iT9t/pJTI0fdlt45AfRelmMBr1NDq6u6EdTqpjdJKohWIPo+TaaucG48mk7Fv
wOAoPmMEKH52Q9VOzo83z4zya11ePNu3LXDRr4zzWdvAXEdZmSkJxyRqiC/PGOC+
PRz2cNbXToPSq4ALqB7r8vduG09APQPifDIykFBzm7AHnJLVxNdWuK9rGmgLXNKz
8gj1zE1eRK+l74xNfi85EbFQScblQb90o0x+s3RRa9k2BeyO+4dwg+HKziKyjEv3
px6cHuNnmzBcQv6p4IrYjAte3Fhw8FF144vge11o7cJxPQlnBsLM2FpMqWsxWE58
cKQ0tYYta0al6fr8UuaIGONgjJzimB2RX5T4JX5ZU1p+CY814LK7Br1EqqfpYRYR
6aHIwZfzp8mLvM4p1HWZrha8+94jvClHkNDkHLD7NDqX8d9S2OUqip8SM6Pcvzv0
OAYC9pLWumweWDNVpo2JWiYJh4SQz2MM6vNrqrr8+E2DRS0GfSldyYxnf9i21YDu
FbgL0wsLB21vBO1fyL0XICV/tVMUumRUQ2Grirn82c0oos94PffK8E1GE+4h0iha
ml8Q3X2ZNMyO+2+6a4uwRU2l9uzHdW9/t+yzCuSI7qdrmZoO/yCKyuOJOcjOHElh
rXZU+hqnZ7cWgjWCxXjX6QxaA8PzTpQLGNmcQYAPDCv/u44QreJHylohYcZbPcFD
UHJ1qrJQ52DftVcHXTUpQDPomWvuPOKepr6cfku22dAvf7d9kD9Oh/QAwN1/sn5L
jH3K+FgfKRuxdwBn8+rIqMf6bAY7rIyfXGPBLh+WjLU2bZ+qdgUCEidhveylkdFu
NVwa1wFj50aU2AVvw6LugYBaYxNUc4LT4gsXrekDYGg+Nz8oh/r98hfqqc1pXu57
o1HK9qoXelO2fWnc/2Gs7LtiAl2icwdvQIRBnA7PMTUClMMTdrnqKiCeZWPlkZUt
4o+B2Gy76dA+eEvSUH6Hrhi3Ro4zcPkoY/UBoYBd4aeawYRszRKZViHuR8TZl9Oy
m8O9H2N5TOfzRxEXi1NeiP/BvdMTzGaeAV9TVDpfezJAciFMNbIG6zuGegssu4Dt
JJjLdmB6O+OnOQxgC/hG0WJ/qT/i3iHSN7IBP2we4YTrM5fxVa1MgRL+qkvFQQWl
uXUGs4IbOaBQKEeIfZCokAJFoSTRVyb4Zwm4ofA9LLzODYX5OpXzCsuYs8blyJoR
zrux7FeHM/qDx5kY4y0ryfYjG0KtPUp9i301HoRnP6pCtXFJF/nNTg2bw3ypFAC0
pNFE01IGBp1O4hA7GCyDCTGtXTRLx/wHN+gyoaw03UpDTUX6uaGZD/fm4f+eBl5O
fFYereTpympBor6AiZfie5mWBt4yX+0vB/TK668mv6uFPrmyED6Z87anW5nrB3cv
5G+POp+jb1jRozzfTrJaMu5e6Y8iplIhMsr8sxt0N92uw+1aN3ZCZSufN99YpFyk
DnJxkPsVovxbCAHH6CzMNqyWofq+oxfA5LVif+ITnnclnB9c0mPZCncVI2bmBuUa
cEoS9PhnnmP1vmnpfTZcynDoW50ZJ+Zt70fs4fxbnDTnQnOaSJS6+CTbqr0cLZW9
PPbp+JTMy8ZjhFMxUD0wcRI5k1Um5dqj/ejnvgGURQhQEKjrCTArIp/akWCEpFML
CMGA0l3Du7WWBQJQjRknzJNPpr915EC/4jJCkJA+bOD9P/oBF+LUx/xsV5EnAEO8
1Z9NI1709+KEUPPgrlNOE9Dz5vTv7SEzyhw5lpZmIIqYV46Ub+cQp69Hs7zEKCwG
tjQXF9SNgbZfX54q0mO3X56xb3vC7cQS853pdeXxDUvEtASzr2HC6vQt3Xy2SYQq
+terGmdbPr92FbIJpVyC5fKAXjF+WdzqDtRbx0miz5c3ViZHg0Qf8H8hoNnR93gC
fRWXKvwYuMlJxvhKUB3bpSuJWz/FK7EYZQK9WnQoIXV2yeaUw2AY+R2MZVu9wSwL
DRwU1UddWF+ZZE26kxvJEXLet/Z799zTWiH6/P0O1JAWCcCGraun5Vvht8OKw/ub
+bYCZZ5UYtbqJogX5MGG/o7NCJ8t5L2ltazPJHk8Yt3ZrPZrJNYd9xLufG3j9T5V
O8OWdLeu5bc+Jpx/JFCvAVnW/nCIh2KVLB6nrQXKBpUD37jDW6oGhav42XFwZp38
F2VgZTLvR6U9CcYqtbONZ0BbLGaX/Vko3Yf511V1GEVm0Yb7anntrK9JPJ+oDrFW
pGtz8mkhwIYG7nT+MjHqckiMsevkZGVro4oA4KPAuGPVbCP3p+BoEOGSTD7Tw00o
nCb4y1/lKcrQTVTPZHDne68YgC77jrFb0xKuIybqv7vJ9Tx4f4ubqN9G6ot+Cw0b
4KH2mLwph4HN8UiMTUSlT4+UzqwKKJUci6qWVmQ2eH06/OgXQB/VjEjUQ87Awv+A
Gn7uc1yiwTWW8TdAJz1EhqzP9YbP4WwvoNgk5+45CHzrAUuYmDE+mqs2iL1N91uB
QHkbRJAEhVcMKCjZ3W2fPYA7tiV3mNPEdOfVRkT6vz6us8HynSoGsNoAqVPVxXGC
GFWgTE1tiqgYIFykgXQB+FtT2pTz0fOfS6bYSzmICBJLIToSQxENEuQXVxucSgg7
wimDXMZ7uk3pDHE8r3/HbmBVNqKqo25NG7KGCVss9JsLR1+9MOTj1UlaxBPld3D/
oIAtoWRVZk3My4ec7kdkef1DBu5haITerFgz46kkjIm10x6K1RQDnLO1GTuXMIGY
fjFcZrqv06Es7Y4UtA6taComzJkO1zxXs03co+2dhd3xbu3y1W2km6AMvY0frCSJ
FICpIlCUVHn+PCglPUwV7IgIZakhZP1rQ8mdnipeiZXmWdq8jutTe11VQyrVdabH
If3hoBICIZ0dPZDeLydmNJzc9T0RtdD1sgVd492lsf8gmdg2DsGjW+AV25FO0OB5
MidJEBIs7VZ6bBeW0gT0ZkbRRHRx3b1j/zZJQg03EPW2Dcxjxh4v6MAqSMvYx1ed
QRtM9T1zV+aGinfloQWjYRqhfPQOLEUER6wzgu1WTE/3N5rJ0UUz/kd5n9oWiiuQ
U9pBRb2BVlBPz3skAIWWjPqjhQ382s+CuzoAXVVLtS2UjtZklkqSAXSjjFgZZ3/p
LSqH4/NkEuZOq+z0TLwzzPCDlTIP/0q2HYIxzKi8acS02ezc6G+DNK89NAAtio3B
9Nrywt8B9mB1tzdQlJ2Mfq7Pa7ECknSHWKVy2VYwh+kpkDq8E4Eq92grU+d7vk6d
JSAtugQtg78xSVFmEtRBIibTi7eaSmTahZNTJbrRdngXVmXN5eeXDAdY0m/Q54In
xEgUE3N/zb4ftEpjXsVVSWooWLBzM1Mfy+1w8osYhK432ntGkQqrPbdRiq3lqA4v
uBVmNeQdDlyh6NPj9PoNw6IYkqFQ0wUyqTR4hHz+VzZX0Pq/fHq1bN/y5C6hLFVq
8zxZ2OotyE3unqcjMCvm2HMlJN93vOxMnq6bfQ+UAu1ncenZcKbeTM+LwpvEOolE
hYKDhj3YWnjUq0IFQE6yxCElUmRrfZZLzpwlGeOMx353BHudNfnOBLhtJc031gIY
+rC4Q/jx6VLMhJ5zzSv96FdQCEoK0AW5vGH6sA2PPJ6HlHyviM+ecfTvkeCfw/MI
ACZaMmOhD5wsGBt0EPfV5XogoKMQr98/7b8H5VY0NBKAeN/GpkSStgpovrh69Y0e
J22Xzr5aVF1+ybTfnSFNc7ZHI4zHteD5I8t9ESXlEI5eCjDQSviun71eeX+1/DUN
Gt+OOHFeE3GIOtscvWozk7nEDbMb9RYqNSmLS1Xtc/tMGZar2qoHsC6QLPVJULf5
385cdVKHL3DMC+nvzJ8iEYXfsmYUQGtlWDda+x9ISRqu72yz5X2kKb8H+8siUUM2
Cu0K4ijUAAz9JIrjhfTh3JLmHXLzXX7fVlUmhyG7A9Qs/5nx4QG1sk1HkOkWp0DG
yO7M3TiQJ5p/Si7RfgOyPqrebddbWZ+I6fs3XTNAzsIQZsPT4Idr3MsTDk9/DCge
o9S7QNYiQQrjD0Q90WBrIBsycjWvDdYY6rkIvg5zy7b1EQpeF8P2XYQNg/+sLMEU
9zTWBy7/oFNcjfGMtBujHtFxwx7oXkwR6Hxdv9vX+KfQL6tV0T6BG/oMuteIzKUv
BEWOgAUTxpPs516T0tigHsS0lmURXlo1LyQgBpKCh/nIyokliFOnpudKCz8WgeNb
3s+zWGjw9sV637bAgm7fwvf4pv2p7ESAqBh7E5JRjCJHqACWvSuHscFNMMfdB9jD
4rzw3AmGwPOpjhr6zITpS4J33Xq0wQLtvA+hdljKtTJfVQuR0ym6uFRgCQglYnac
J/o8ieFNaLYoHJ+QRKnkJLn/bdazPoSTRG5jtVeqgUSxIxISMmNBaVVC1+1mDiJ7
w4pkzNEV0FxpaTCdPB/bPhxUmL55cId1jp7krLYqpvPR1TQq/lcnI1+qVN9VfsDS
Xp6zlXWMnqcD/BAQ/6apmGekdDDqRjz8PU26jLQqWEA8NPP0B11bffQ9DWR2nacv
BOeut3MGTb/U8OSNqVSSNqj94gztbSygq6jL2FHx4nqP4ZVUsuRjOk7kHCV0l6GZ
92BMAQaIlTNjSAbZKrhLCw8Ds5Qp/gNFMb/jYVnm1w40Xw1Pufu0fAeXgbBUxrC6
XuvM4Yrfr7JE4x63xzmYxk7UJTSPhH861+EVcjV/QLDqPstzwIUEciLJzmKADoGF
j0xtueah/e/ZQkChBn3+EJDHqpZGBisk/GN/fPx1MILrDYYMfmlPt7B7ahwX0eE3
pu4YseIJWN0gBaUdIOHFYw02t8oEs7uqt/Yo5XFf3P2g4lXbhszwXPEkCcEXz1nf
pahIvJCw7m+1QcIoeqY+WpWX5KMVUrn3vggUldWrq2ZtETW6NZAyblkmaZc2S3Rv
rvLjN3rGMIX8pLoD1yHwE3JFrhJISyckywcV1dwi/x4Drbcb3cwQYTey4RIU+OeV
8fLdBEeKQ5tlwtnMj5BUHxi29ZXzBtxjJ4vKsWvsxZ8kE3miv0/tHaKu1wO85DWA
4eYvM1HgJ7YsM9iyGtSlsExlx0d0x/SeKwbBZ1VaC9zyzR1g5tSWELncfStW6Fxn
lUcRi5bwD5IcfhxUYEXdHHkkhvMfJvJEKIDa8mu57enz1hsqdJTUCsAjdlTlQHLh
qwPWZQQPkxPYJHPwArVkKyPB8yeZ80Lae8vlw2kk7lRLB4Q6DF15FIaeI/xhnYx9
fj42R8455LiR2v8LWxRrFAuGSS38Fep6jUxShZ+tcGEquZMYVrS9jnZ4/9wajGpi
RNazxlu65P37jUfVDYQiSjrbtFZSfl3t2OtDTDXHX81eFxy5oZQbYXLBVgmyPhMa
yykWBRpXfiIAafQ8deHmkpggL6cGAKU/Rt18zsUC2eka/TUs8ZtUMA6tF7dEWp7R
Rq0BQHiSk2FWNoC81jwZo6ovAiXHUiWmE9lMu1mYrfrrXbdJBP/RgINI7v50T5ac
WYBUEo9zmmZauA+JdMOnz92xJ8Nf2GjSehS1/gJM5VE4/R06SQpBYLzCV1rjYcHb
amRj3I/Mwc+i8YJmTgx/gUpq9UN42QWdll2g0JrrB/RsHWFML2qZXytjKw8uev67
CYYP9vCg0P1WsB6Qlp8GKeD80WeRNJkUaGIVrNBPW9p3xhV+5nbiMf2JFp/e6dGv
sFvH0GmQiWhhzXrhBVsJloTcr2+SXdJJqaV5ucTZb98Wwm4nD7xBTj9ufY1TxXt3
49h2knyV3nU3TN4TaL9ej7wBtjt49WRkgVDH015X/rQwEE3V0C2SRV6YYmzfvzhQ
CRRowgDx++IdkLHI27ZpKLcVgjgXC7cVHzBeuUWi4RIEm62tyDwnBrI5xJIPsg6J
pXvVsYSNunqBrWQkmiYkh128iQM/JR+ulzbvokawCb6vrCMhVVTrugLJuM2r4D/F
/slZC4TtxG0C7WiJzInmbitSEGecbgyuzJeca+m5LCmXP5GJM3lE4tXIuTTkU2kC
aYxctcztGrpTOO8Rtk+f4x1/lP78ymraq8epEo6iUl+y077SZdqhXnzxg8OFGCXi
z3NrqDzpvNotpGAzbBYI7J4DJUEMsqCoV1sHbOQaaIVzKypW4xwUIkGdqyKo+FPB
1x8kHfR31SDT1YkYBxaXe1k8xMA8pG5225hnPMYvD6BjjvwZsip28ZA1xe89enhK
si8SYzEMlBAe5ILCp0XEZPQQ95js2HAB5nBxiM5dzmEF+pKXErTgKhicJ88ZSm2P
MyBSlMqzjcaOn77xw06TpELxMnC7Sc8ckajKxpzlfFaJ7u0FCJGdIkTlZhzZDgYx
FHUHLxHAUIr2mss4mW7gDAYIft2fhKKJ4dJ3DKo7xwXgn/MTRRY66zXFqsvyegcH
jFtZABCIaWFRUnv7jgWswgKyCGoIVvExHEO7XSTDdBqbuPBa3mbveUk0r6HD4KWO
REkcNM3P6jPrIHO2YAxbao3svb53mASsuE3CRqKAGNOdQRBaJIYwkkv3wHs+S6aZ
3ctO1H4sT1PiWBTU8JwAarLNT73n0fwlAVoAQivJ6fNSpr7T4zOn6SFMU6xLQxPC
nVywPKw5/yk7l741PyvCO6uWPJaRTJDDq1iEUVQUqJGsfKQdsuKhIVZrKZq9+Urq
7Oz4TrbOBAd5swXLtTwwbnoo64VCQHWqaANUbUgN+xmcY9I/iRvHdRvzH6phr2IW
nTs4xol8bbibowgYfrOwdVB23Gg4OCHIJppdu4/hutAA0weDn9Txm24oMjYjvptL
UN7veQU8gfLdr3OH0AWFLJ1uPfX6bK9mSraMYSvNhKCZLuexHM2Z6JqGm0QL3/nE
B1lH3xMyz6qeG+kpoFGANcLmbBUCc47UvtgQnA8gKr9CsHvPBWIPuueI17OXFqrc
kIY4HYXk48puG81D8rFr4lJOxESnDlxk68OiA5/+vU+IyC63QWDUxZCbwwWUuZzZ
xSo5MMnOFol2J/AAuj2/rGS3SKlAkUf76PEB/a+K70FJGkr3lNxD/Z8dXbW2ADf2
7dSDWuNahZGe1RjhJ4RpfC0EwJV8Vp9rlLWfttmwV1t2DLqbF4b6i+PHsIrlKgOZ
yx5bllfOQRtrBfpEC62vhOk+cWMMEMvh7I+avgn+rDzbYKGdn8FE62zWvRlZ4gc5
hoLrAQ2sxxqD5uqMqwU0H0Ca+m1R1fd8WLz0aoQXB0pW+o4I+eZGIVebv2b+Xvvk
iNsF+NUKdeRJnZVZDZiCp/i/cUYW3Ht2co7bABCF/yERCYmkHeDTfpoHhPEr3JOU
iIB+xmWp0vPVbwb7T1OFrdjawyPFlKUXJ6AT2c84UZfEvG9CeMv5qalxI9/QCxg2
q2Otb/NHt5ngP2/PdKAaLtPpv+zBqrvrzlpfSnnqwm2z6GZJChTRTgLjD5i6ETrs
RM0T1rVAxBujgjwAT+QFqVdC9MBNLMuz9qdh2uaexZSSerBvvHNsz1WXJYXYwDbp
0umJa3wzvG6Aa5v7JJr1zBtqR7WDe4TikwSa1pmUz5041MHTPBMliEiwZbncnjNx
2vgWtDNCSeZ6lsnqzql29jOgdEzBtpA5DH1mF75H7ChX7/uzaBCqTpy0MsE+K3rm
osaYKVLvxZp3LL3UQcanF/vVxeQ8f4jxuhH912Xyt5Wp7PtZfyoxl68KwuAiY7TD
gxPM1r7weiWyLxFASWrdzGpVhFIpT+Vi35FXXKpjYfwtbwPaRMyl3cU0052BVOZV
2dSy56eBOxMAnOus/bBLyUVm7Wo6wFTrZycqWAviZqld+6ZdZrEiw24cnwf7LPOV
IxUidMM8HrFNVLn9psxGhbsbb4VFCywx/9pR6yyjfskAY3ER2PZ95OOYGyeR3foi
WOqGZIUj5JibNeKxyrkdlnwgSiThwaj+6yLaqPnfBbFDA2SxLuUyFyCpta309tKe
WfjCzsRknZaHbr9PUqVGduNiGYO6ZpXjeKNdZs2qAT7/PthLj/sqgwxDQEegSatU
nLyF3So0YG4K1AJ6IwE2BjtcTs+5za8jE1Fjdwo4lpQg9Hmaz70T93/CVZSPxkAl
Y//fc6tKdRZRRMSYfbnGorGoq5oOYaPe1o4SNH3sfR0h5gA5SMusJ0Ji7EzEjRXQ
Fx2+jIddhqiofVCUxzG/NggqdrSuC8QttHQ1f/mx1lKE0xkRI55/qWY7o04ZhgMF
i+yhSzSRHdypz7+xhGRdVTJVMC3rn53SlnetgeGJlL3bPJz/6A1zojuJ//AxbnIR
EC6yn1zrQ2MwIoFJFFlzv7D7ZXAv+aRrvkcXEm0yCnH/+SqqDXaQBS0Fwspau8v4
WGVmaaY8KdcTbsuzn2dNEw4W1OKfCbFUuC8bh4KPZg9Uh+lI7nFXhYN8U5BYrDDB
kvtcXPTHVZaE0lJdKHghyLZ6pfcRyhdGy6tGjpyLnBOm0MMiQuTu5LavlhSzTp6+
o5KCaB80eDdvcEg7GmtWNmHJIvWIz5tBu7dSpIVpslpOYktRfhpr2fbjtkJpXRSQ
4Yr+PlC4id93AWPHTZmsqckJ7HPRUfIGOwZH6wnsHRFKxHp2GEcKt7iES4PdX3c3
xlIkjNPz8jyMC460JuPNVrg+Js+SQuIH7+zwFAp8Cri6wIJUA1bBFRveZ25RMwOc
aI8wEGVbLYFisZtgswaqmOIRVITJbHvUxw6hW1eXHnTCpcD6u5uOIP5O9jvXNAzH
vGEM4EGJauroBzbihdk2aQFDmefyK4nKp90I52aNfBGdcmTTOgb1tsQpEMx6MlSV
aZdQ8PNNDRFIxOGFnEyrmVFqqkfGVuYurNGjRF7sbAqRSadPx+TElKmISExikCkc
F30rYHO9rpyDMDHsEhNLaBgft2zDIF2X1jwaAP2cT32fOrBz9EicE7GGADhZaaWZ
GLJBiiyLFpkX73qfZ30wTNnoEgrat2PefHgneM4CXOo+Cm1VI3UdmwYT4Nc6jLpq
feSTeCoXWnMyJCKap6Nt83rLqqOMC0NJ3Cexu05Fyl95Lgv+/99qi1jfBGJU4+Rh
84yux2TK3L3J1WkbepwW/m7CHq5K490KFc7dCQJSpJREwRWUsekw/bQWNIkaHaI2
s9EU8LrKjo5rWrlNOJb3iPlNcIQ1cRawuUNQMqIqK07ofi4eThzNpcRcWbto8Gyy
XxAu6x32rLQg/7X9NW8fL5T4m2wIbqpnc6ayJZdeTLU/HCYp82vRM2WXV7sYYRmV
evO+gNaOIFk4MuKs52OsR1m2XoDvtVgpJvQFSUTOK87Xkrti8k2Yhdg/ZfU1+kUd
CkR9/SA0bVgpTRIljP7uZAZ/Om/s2GRno3k9yqEs9fB/0oSEr1wEV2ix2xH4NiPg
Hw0tmlOLxIAlucuE1qe8AGPeS8DrUU27B9gyezQ2XULb2O271nrci8bFYCRoozX+
kSGhk/Eb55lbdbCLdeDpeFp/79GtVjlbj8E9Hd6CRkBb2KY4K2+dNp1Wdj+Atlsi
nTCssgs56jHLhotFFN+rf74Z0/a6a2mFHyYU9Adc4mqtJmlLNcXwR2SOgT3m/BMZ
FZqsM63LceLbq5QSfUTPqX7+sWx8w+cQ938OqXh/lAeQMKs5rYxU+OmjOQEnxsce
VQ7xBcRe9sg15oRMhiKlBi8vLZrh07VOWCFxHXBP316fONB2CeH5RM9s8mFiqB/K
qsOOY4jT2DQ1LgTm9ii0y+ZIWHUyMkmQzNkJW33KhyDATA8pBGC0V0BZElTbG3jV
Db0cPepzaQRuIidqwH8Q/hx7DZULpVeTfBvIp3lS+K5os4vD5bQ+5xqGgYjkIFSe
BCB2c8yrFCSElbOUj0D5HxlAMytY1JZMsNbv8E/PTiaUsE2/Rh62x1ljagVz69E2
wCTaTRvr62h46L+5idRZYbEhMpkkUOhU718ILPfa2px8FH9+eZqPWNAHtThGG3Jk
6t5ow/uj4rWlCgbomr6Fun0LQsD5BOChRiRcxY1SU+AHvfLgRHPnqdwV/GjwrGEH
NPI1QGE/+qR47wBqahH7gDQeNMiFp7DR3IJ8Rmdhod5L5hyipdPdYEjK6MXXHECp
UpgzYilmnzDAuuO51/5j+KoxUXWaNbo/ziHO0zPUsg+Xx+CYI2WWXTJrsT/cZMkN
EELZacI70Q3SdQwTierST64OtQsKFogyRxtbti2rbckbkvxtvPsmgqK9eOIfkNKN
BkTMr2+o+/rC6Y/j2/P/5MslxhBz3natYTqyZ7HV1FHsMzvivu1pYw+UMTFveDec
9Lx0yfDYx1QLBnLj3I12OJGZ19b/zFYHj94XfUa6hLojkMO/aUPLnRwyVjj3yxiv
2j1L3O/5fKXVp5qcCeww3xI+ZT7ystSZBe1ljnlOE72cKKTgyo4EJAnNIX7K/iCY
p4yq6ZLWosC9mruasjuvpfTNZXwXEtiHNZ1dEgMFFEwkPKC1RKWhL1X5dUMwH6uB
lBWCGnks++owOBxOtJs5XowhFj7CBI/pREAJ4bUWN0EnchMLy6+l5swzT1PYQ/l5
gM1GGHPGRc+MyOOes/eyK9DBJFlr4eQF0PcrcVxW1sTnCsD71Jgmgg3qcfkZhxPs
Rv8at9j2wDBmZ+MVimP9k5NoEy56GKjnqh6OksDn6yGEurZnYUze9OmKYClGvQtC
CRA5D1rxX7tYXbAAZARBxBZd5tyQ5rjQq070t2kf5ui9aMdx84SSf51tXEK2+xrz
YVnpCLlwWs5vofueNYZJN9x/qjWoxTsBZ7s3m+CkTse2nKzkaavNP79TbLGSY+kn
9uo8h+7zGGLwrk/JmMZjjHVUOPfToPdD7WLGkixTD82vfvSnrxmURt201vNz9MeM
8Dkg79nBuDtqA62cfFsQLPhTyQoFLxhGRd7iEfUKWsm13ZEStRTok0aW5ONmRp1w
XGU15eAEO7b8EFlf+56Uo6hOIeq5reirX9Z+Q0PTKBwH3XEJjW0HSnF+qrz15FPj
5gkZ/atxhZt0sqfY4R5FCedDsN7PU924e1eghmV23uKNqGG4NRPAnwLMabFXlrq2
FpruBrH5c1th5bCvTY46cSBlojJ9q1WJk9y7xkt3W4y4Q+/bWrwL6XtZLAZrDMyn
s76FS4y7FRAVTL/HuqFZECFEJ/5JmJgzg8bCOVhiQcCX6C3IiyEk+dt2RnaftRA3
2FovAW+Ohvk+1V1Fm5Po6Y/GyOKYJP4jMVlste7sd7NIWy/AdZqBiLVhNpwFg9HM
z2FA2g7je7aLT3uxbj9YDHaxRiJI3P8QGBVamZbV1K4UlegsilqTpTGXkYHI0Zsf
iuer6nO+BaQ9pBB1umN/sShYk1e3NWvBkGFHedXAwNLcCBPfHX/gLgMdxEWxeN3h
fiFyyxr7I0GvVSpnEIr0xG8V1kIBx8ST5grCeb1CDvAA6NJuToouqZn0GMa+sT2b
9Qbt1dV0dT/qsCPvUOI1dYfJVG9qu97eUD7ZE57FBTxTo4+k5avunBJKtyoxvmgt
BdrdCkx5KnZyjZOHG8myNfag0fa7L+aZEH3obFFQHumQBq7hbB2GmEg+9DOs5kqE
beUFIWuVpWClVApnB77VchCyn33UsBiaFkQJSgedDV7DytulxW/sWKUPbHnav+6V
m8yd+gONv7lJIgGX6EjtwdTNjHK9oroiMzIKB7EjoqvZVYZcj+en7Ou0r8GZA5K1
H6jCeB50a4DkvEMnCWNjC71hRNrrL9MH1YqLwxWqEKxIX3myHvQwxXycV7459W8w
MaBR5urPdN2HgwFCfGCTEfrMnKwYWdJbIdKhZUDIzMngoPS42c+94tyU+psHkZr7
c+rzt5tvdI9j8LPG+9Br/LHUeWOP+pBHZY/t8AYr1CsUaj3zVUARVSrU80ov7NRh
QARXcacmV+QFhEyVIQ6Ye9tkmZ7z9uWmhD9xGIKD9WHHVrsXTHUYUGToWly8rhzf
/ao+iEmfBA/ZkO+R2O5R70mIaOdM9vTpVQzRdlR+LrGPyjUh/xmcYS4sHKlGzUVl
A/lseiBxID63+i4BqIMcqsaDHUUm4L1GINp4yeLZpR5MPLVPzgok8wcoyQO3ovog
BYR+Jqng5fxnYd5yduPmE2gUwN+y2nhKwEl3+LiUvmQdKWVruAjImhsCwDHFt4+i
tybOGv9BftTC/evoypxz05SVWoW+xUQmIx2k8Hoy8Z31nKeCfFwC794pW/2ll01l
LfklJvwE5Of+bWh2/icG6AUCpPUAcZTfMV2cRy2OHT7UUm+RuybX7On8qcvfVbwT
UjhYZoLgsAiKb/WBEq51Kk+Pnry4fv4YdwYfsBbxWK8HXEzWKsh0v9j0Ootnc/2s
+yex5ruzoUaw99P9FLvX5vfu1zZlwWJiPzqbZRCjw6yIE8JLVIyJv646+GqxjbcB
kowzVwnkXgNShTf8JFwF1o9v5/33w6E4MIvrY67Iu3UJT4x+9TLbVi0WXHR/BKQO
8pQn10xcYEMry4KZW/UoeVxHNJhf45qPFuj6PKmM8cs1ZVQmuJcNX6UGcfmFuUGa
qZJAPctZIWn2uWQcRh+ODO/MU1+iIOTTniKdi2fSD95RlckisJCePq9gvlrTrUBe
LDevnkVF81SQ71d4ejIgwRzz3O4sw1ZJ7PkfdOd6ApUxznlsoSp5zNcgRKv73y9F
Kkal7s9strez8FyxYRN4hBYgh3JWAHS8MSRHKNHKxOn+azdvqHvhnluhyb9SWxVG
TKsW6w9HaJhe39HkVnCDg4cKDfQSbJGfYKQ23zRdAtjtwDOe0ilb/MDIJKEZB35M
NkPNxuPlvHoJveRO2Ke4wpLBKnS/jChOCkIp+1+vA0JbeK6cjdIxm6SxMarj0x7J
rr1jkS4w4dWTFmwHxF71taW9hjbiGeVEYk/ZPTR+UcNI1kwlSCIKSp29Qzj+00Kz
q6nHDQCjJlO476ZChR2FSCOAMXOv2qmSsprIdN/mvIj1FALEoksXSB1vIION/1Bq
dfMR7xhM9keI0MxEq392Rx8Kac+GA0tuqxvu0+xRRTnMerPN9Pg8FaADCE77Cfs4
p55TyPJMD9/S4JFXkpEnyPlLDGRLGn4N4IiiL2EUbxe4D4Irem6BVWQJU7+XK7+y
C9JLBxbT+JkpN+0X7t4qqscAqMLW9ckGg2n/e6spE0T7xz0taGGCDibE1bwVtSJh
wHIksl95B2036IGXkwGbMWDOfGXtejlH5MTS+ebYnGLJc/QQxQI5/VeBmSd/a1r/
8i/qok4BRM1w9vaAmhAbF6D2LGKh9w+XKaNkvEcWHssO/Xc//b3usATs+QuH8Y6f
bjmW0z8R7eCndgo8uM6uf6Wx77qHq8PlkrRpXR5MK6HELWOD1rWJBgmhtOfTFKH3
5worTbUeSOerHXVxNdXZuS7/5Go7rHNX5jrW8dox+rbZSA1u4ablbcXXlcSaEmwt
jj1Y/ro4GjqTDgRG7A881CmYWLojIxQbrn//csnoi/UEwixptL4q1GtZ+mwE7brx
X4HpA1Qokb86KQEP9wB2f3VFBlSqxI6bLgBNEAdZCWcYvDAQYczCIcFNo8Z+kEyA
lat1QhID8tpY9nhM9j3d5jx4+xne6oiWq8ovZey6l0U+ixi99ifXD38onENjuAam
aTM6r+hlp7b8/eZ5r5uB16Z+rYuseErtB0eZWxlKoyKbUd98rNaxDEfZEFv7tb39
6pEsbDP9PZYXd/fDHWytrYV/ylrimy+N8UOupKnO3/8QVz7RmT/U4D6M9kiy8sVO
SLcyOpjaHTBxBa0UWlTMPLKV2e6r1NAfOyack7iL2sSd0Ch0lW9DU6OSHRGTIKwG
ERr6rz1tY2G+0IfPF8YsAaEeMEFFmm/w12sKvbD0KuIozZNaYVUxLn57clyWsEqS
6UgIiMG3EJ32K+JafHAR1i5GAvHRhtODuo7Y3BnvsdA3OTWy+ScJhN1uqCpBtQLX
iOW/YHj/D1G3kcLrdhKc0PfK1ytDfUsTUb0b+kpVnUzsafPZtlBdmeBXtV9aZzV4
cgpoa/vASr5/W/21iDONjVQZJHqE2H+05UvYfaiFvX8rQw4lPHiRhX5IwjcI4I+M
ik560kBjah4m0+CIBVa5jC0TDGN0zglkFVP8X0Y7B/s7FCD/yS6BGa6+9NZJvKf4
qHl46GEY7YLG4XesnwaBeeyCXvAGYJO7nOLBUVCYweAOaN6YNWRmZ57TnNw9xMlv
1n5RDjweT4iDDXg9IM5qRN9Pi3fWE8r9hyNzfyLByTQPK+MUKjJ0SQeE14OM94L+
Wht4NH02SDIQD1jK0egsIr9JN+D02g0Io5UaHo+jdfFcujj8kQuqwI+6ELmlOHxJ
TAzyGjI0FpPU+bcXVzTjVl8uhyEq73arg+s4aH9YgpSB3WYoGTS1YLSr6MwWx/KB
3ALBD74Nawzpbr14csUhcWWCeP2k7QoGXivs969QgYO7NIPliaauLNkhwx//g4ze
QX1IoRtZ6PqXpwkZnViQfv5tJNe3TsYdIoQw9RK8LRwsTG2NVI89oPtdcxGKkOXK
VuXV8H2PPb3qsALDTPnaguX/5ekWZ0taInpP0soR2LXBcztw6odzVN4nZ4lCZC4C
0miTn9aQOiMMUXTpWPSkPvdhH1fjFDvsMz5hMxvmpshwRCILDq8aeJtYzDIFX4oo
HBCHfE8dHpsqKkjwWrI+iDOPChs7sVvUtA5VK0Yo2ro+miBUrGbHqWGZ+8suPu+M
priQOqTbehTqkQaZ585BRkOfx64xdZ+/hjCviuaIugzQK1nMmBzZFHo2LhqBS8cp
BE64xKVHRXfxQxCOjBwsdfFJGuOfD2+M2d93OsDOwSZkANT9dNxTIg2Mh1efHGij
wELpfPfKm6OCV7Ntjpd90idfw7DZOMfd1uubX80/9nhEy4yumxMx8MuuCus0r7Nr
22P6rsHym1yVdPZeMK/NaWZSnX4dxEkt5kHjhXgdheGHvzPJMY5cUwBcLjShlUkM
TAY2/KZlwceoKM5yEC1boZz/ZPr55YfDUrAG3pvFsao93ppxO8GFeyLw6yYWHZuE
CBjMea6GLqn67jzCwTwDJDp0gvvRvLpujJavE90rMbFQOX1qRuUdThfMae5SV0Cy
a0TgpBjCOqrC39Vl1OVI4SEW6lqUgkvnhmO5JFmVsVza1l/d/mTEMraButNfqWrs
W5ktbwCorgqJO1gpLib9Sq7FTnFEfs3fE1OqbWL5qaJ1xBjSoF+v9qgehNUtUfAX
1Dgax3anfq3EH2zhUgu7VOJXv6sCU7osTNfdjOLMLELdt04m6yJCjdLMcnIK646j
/UaZfGHCyt1gmKUxfpe3zbk+JT52PyrY3+bOH+3CQWDyLHWo+l3SugAUyJeKp6FH
JZRh+lB0D+hlq81oGGvm2aymhDe3Rky33aeOgnT+8KwakpnWk4WA315mVl2A61WS
I1J8lQe/i3qzqHzsr+6pP+OZ8Abg0HQvsJ2GITreIVoV4dh+7PQICBccjaIS3X6/
FCGYh1c+xOaxn7qMib+AT5s3hBblPp+lzRM0rJWsf8jUmQLA1DUtubFSTtYKhb0B
T0BMr2RwSj3yozy9cQFkxW6V8XV4oubNDEii0oYfRYJq+18RZPU1hIFYEZ9NGNGV
rZCdj8TRqdGpbyeB7D4Jz/cw333NfsvA7EfiECpwz8mxXJSCFNB0w1tTcH6+SAsw
Q5NQrOrjLuQOktwueHpJApqEkZ0PwIecC2gwZ0JfqQY7Jrig5k/hbOwANvp3rTbP
Nnl09RLYGct5UTTjM7OXxRxx1U6tQt0wB6DWKQ5CPgrLKF0k7htsZipedLXlCkmH
dIZhSPQSmhvgI+ychQV8Sxj04gCfK2qT28lMIE/AXUSXQXMDy0nX8Yf7r7TwPfsE
7Xdzq3StavcDlwUUjXBZE+wTFmJPoYEQDcivVmSdfSR4+PyCG7rpQVV+1K0njcCu
ZMKh7lLy5WhpikGSqqQIAmJZHkm0mDdnzBkBdgWeW8JK7gdum7xNtyqgnTIru172
RJXEw0Q3lNa30Dokpz/KYJQwvXO8ZCY6QM74DAGQD8dhC9TkO1z+OjA6KG9mFxzh
y1/su0VNkXgt/QMbxbtloODHHDpkEBkXaRSebHb/kI6mAMNaUd4+oUtwMdpyxbMy
F9fhUAa4vXhbtoNEZKuPKMAmz+1N+HAY3/58VND5b9luIpTNL7B7cL0VwLES9Cm3
VxG3Bvy/eUYFRZtGXCN/e3YsnfUjFheFaSES5/c9AyZ7eRR+lWF1A785EVhiu8MQ
Ut+NJd3xxPDb4ohBYmn4g1yH+i9Ef2ZfTtidgvscj1Us97QIriQoJy6cGvRYVBCv
kOp6oJ+TZTe+aA/3TVl7OWmdcPp3lT16Whe8kK2Lcsw2noTkvuxOXyqtFiU9C46m
zK2joojB0w+W/L+Fi4r+GYIzX7pbETK7r+JAZAMCkS81TjAFch84fSrmKVSZT2Bn
alLmU1FK7jtorObvsz84DOAaIGLVX4Q/fpnBUJ2G6lt61NIQZMSdN7DYZ1y08LL/
VtwWqlg4+Yqb9grkcxxlYbJLXiUViKobf9wBX5t/K/eqozcMwNTwF7fE9IShL+0F
VroFltz+JO9QgBWksyrFrPoSiakNAoN7e8UNZgM6sJBSpM2a2bTTEMMevw1Hf5xY
rDxPZ46nx0x0kzVvJc56K7O5N408bu/K8fO6+nkDcxofNl70UHsMr/SnTBloQhy9
2AUlGl9YuRdy47gij3gLJYAsLLScYvj7rdvi+mD2dPnAdXIKEKNEGzf4YZ0hEDQA
fmAjyMWgK9hYSSjGZQ7QEkyqYr8haTR5WH91aWzByy3/FHJmrjAGkybTPfSc5bes
gkEluYs1A4qbmKhkEMxX6OIclJ5iGR9JualVoQHHyKgNYoHs3fBTiDLYWA3wIwh4
rgJlKvj7zvuUgixj1nc6uqrsoNNVlSawEhVsJhV8Bi81LLIaSr+japu6BuIx3I2u
eHxYRJWehCRY144vgH2zB2iEEGS5YNZ1R8X80Z8jjCtut4ff3Pw9L4FZNLacIjQy
HdqAu2QCKtTevEImZ/i/RGGGFUjsADbzO6rn3VOfjfDjO8WYIgolZcXgReJPCSF5
/irFTX6bMnotvEQuT9pu1Z2daCtk9Dmak9rhI6ZC9p/aGduMO4ksxbu9ZJ/ay53j
kyZgSkMsqW0swl7f7g02xy1DiW0B7n2eU8LqXKWam7lj3hTC8A+EmunrNlk7FXdj
Jra9MsKW0WJORkzHI6+e/94JW1uLXi0+3xLslPYJZMCZiWfHh13LBiu+pO4gE5RW
nZtUYDQxsuVUQiiUgvGFYwsjE7+RMXzA5DrO2eKFnG2guRogJUrANuWCrgmTh8vI
oI0k1idJkRrkEIu/kP0n7N8b+i0J5ruVBD3F8pTB3QZw+GoioecjcYAx4UBy9ep5
Zg05oDREnAK0rw2nX2ItJzoKYao0sraEy/6AKcTXxJI6EKOyngnwveAAoEPBZfz/
29UPxJXqD7M3tHuvdelB6kBpaCo4dbZYiiq9zgPPpjVkb809CKdn94TftADr/reI
3ntixYL81XIyWXAV2sGSUfLHQPJiZQtC240ML/IeqoDFcfquap3HaIObSC0vo7fg
vG1qeEjiVbzaCQLJc0ianRZ1Vk05nyJqJYXekMkpKvmVjw2GYdommKuHbxYo+RvE
G3Iwx0awbTpfjvFZqJMGf2KaEt6ygrBSTNsnTh8Waj9B4tzxh+48iDdXho3t1gBy
mYfLyRaKoSua4uPzWnDQ/gM+F50M7/htyheceBO7TvY1EwbLerAQAA1ds0yJdKWC
G21Hefh7FErUfS3nGwHlA4GWR1qXuEoX84BkCJ82KFnlDobCGgQqfHMxsRL2+gxe
VboAFj5yK+1Ddumq2WHOA24lS3cMuRyY+oIvw8OzwDEXQX10bv+rxQM3ufUEkphO
lZCSbWd0R5dowUkwUKpgDZe1RygrOZPXiqLLbExo0igFhJbNIB3aIh+yMufJAvxJ
gWWkKt2qqkWH+Vn0QXOecj9H08zvPDNPdG3cIQu/kd7NDAqLDxKxyyvAbTsgKwo0
dKSdGMJw1DlgKKjbtzXsTLDJnZFd8XEluj3eIy4vLGAdRdM5qpWFkVpA9gflrcUN
UHcTWXFcaE2S0OYxm9qmfLqiXhzi17vEkPR4NTvpJlvuulSGzxIrZx9WFYRjBfF3
Jx4oXXy3SBw+WQ/mhSMRrVGahqBBh40VtRfAUkEeT3wxPo9DBmxuhHok5aShKfc7
Bq/PAqP8XtAlxTbSnybsASgodLhg8v5qVNDbWEvIJR2DpAV4ZsqGqYgIb3LDvUqH
sBld8+ZV3c3Rpt4gBJ5yVmVgsiskDMSlaZN+74wvDlWMuEMxA5VAYwmxsubCdcs+
Oa/knDmJBtciOop5EAbwtXclnaF3ysNNKPhvuYkLSNAbsBrIIKW0SnnM2Kk35thv
D/JTBXfkWirUq34ujszSjb+8xRHjZFQOtAFuVYjZDr0DmVUVrRYjGLsWYfVIzyPl
4chXV9WibU01Hn8yeupgyCH0q3wx2Lf6poAkiCu1uOEMh6IULcoQpjiWrP19eXtt
T2khoqN8KatzIo33yMSO1YdOH1k+qQTrJMkhW1ty3DRmQ5bHGBpKqUjP3z5FgSKb
r31K8mqYaAUNkOAh6TcPN921aLue/a9iq+0DiqtEpKsXJNKRe6U+mOOEMYw9/K6d
bHYQZSwPgeCdVgCTlkrqCjFkvefDPohQE8100lrTRTmMpBHs8Je7g34M/MDqhP5v
AAoTNEPOhrNfj1qHHpoTNnEhZaJE8ERXNnuA/PppGEaA+yrMTGr2NG++WWFFphnr
h9+tqh1ERRQGnc4Z9JO5VfYw9Hll73QZ7LUzJNnSrL9lJ+fW+zi7No4oanLEshTF
PV4Akes5uIP3aGgfUHMIuKNaO8shWzZALS2iPKBFV6UCPJdS/yIl8MRDMESnu+oe
AkXBDG7YrNizE3Fq/hLMFGkYtGhSm4ltNjxqTWQEKnm616imrAuXH3qwrbNsEhnA
YBrgDSqKUktVyn2q3cwI49GnSJPO5q4gFa0Qzby1Gp+Sj9Bj0RxE+nNLKvg+P4Il
XsCYu3wWTomDAPtyiGIKD4oi50r6eviM8VPXUlHGltOLu0L58GvKJpW23aE0X8Iz
XhG8KPORGiuVYj75jfnajkvfnNPdq0I22yf+jNPQ59yI+RM3DPRAwEga7W2O9bFv
OwrwkRWCbSf8BZg3kz8JzL7jou1UGw//SanVxBrITzbMf9rxnIx3eDeTs7ZmhpCr
SgCyCwcCwklHGLoUin9Zg9a++Tsxjwjp0lG2FD+9mBPs7VI0vQi5KoJktr61/Nz3
FlSb2rSwEQFFdl/h4iU52Th9/RwT7EivABboKpRMdXk+Fr6oADkeoFNliqy6llMh
Txdxz6fMtNs4QZ+Bph6pt1yaV0W4lJRyCQ9hGoSpEss/4Cmr7cSMpguYP/ypXLvg
anL8YOWnzANTWPTDCVUR82G6QjUbvBq7NLbxNAM9Vo/JZJms3xVpSXbWx6mnB4rm
XBrpQKUxPnRbcuFC7Jg7f+RSzdamY8IWPUXFmSKUe6N0LVxoIPUcd5oj/5pNfM78
/h0mRKAFyEYmnahNW1HHvP96gqnZ0sy+kPMzFeOXHI35Mlyat+6h4eMyqVgrhxWB
ezg6hyJ5UQuWZijLejso/FTUW4igZwzHpf1tpdc6CCV9CypFzJpU4lEUVREwPBLJ
vvHMTc/06QdrZ3Qv4inWzvK1ztWYQ+W6CovJpta8lSDpm/bWKzUTM2T1VmsYgmjR
+ABnZZ26vZSfl7M9zhwCk29U27vmGgXqBLU1FIIwPYXZJjpgsPmHDn5LHGIGoa5n
w9r2qlc6QBdeYYKc1KNx69BQoxGu/w7+CKeqqVGRc0t6vBfw7pOtnBQHMHAxNP/f
q8ljeBMZfRv+S31Y/zvZyffablFK8ufFWU76oRFkIw0ZAVLvD4D23flNRQAZN7Kg
qurNyNbUnbvv1saYrCzEAYWj1XMSvVYTn0Nq7mjEALgyliEThy4yhhtNeEWL/e9e
CNcxdIFfpsKl4/zDe33yjj8lai2E89cNPWs8n4t8M+OLGauK1FlNpEr2m+yLePQa
Th071WE3/Q0pYG2H4YWsz7R9G8p+jEi8WpDMVO9SK3uCu0Ik9lnIb3c6nmAPaOyU
QOHDnsMt7Xpm2QbZdJrMzb8hB4ChoKJPjdIFutVlfRjKG3vmXhY1dnBvPte4twJx
SC6hnnjWmmjRSEwdE4ZgxwH/AFIM3VUrKdJ+Q45VV3SXjhNSAwYSbsKqR7uKqowJ
I+EpTT0BHq5Zadb169JSNFSBj9s7lhZ5ppkngHwwNf8cXGXBZPnF4FTBD/IVcDdV
fPB6CEq+o5uYmlADekhMGJPhWzZsNLVuurmhfQTnWkAKrUQhEFZiSIZtbEbWfeCl
uIQl2J050DHgBHkduj8kuGxKErsg7IzABLSsdUcDaFmoA0uKk55lGrQembVPMVbY
5XuC5XhdGsiEkgE2b7Bd2x2ewS9xJqi3H3sRuIjljebk1STCSbFj09YyrYfclOdl
76e8ERUm3zI6NdHyjjMd927qEZYNZIHsRCbpJnCRccDM/neR/4rNLjXZF8VqQLRm
dEjNVsQjuvDRg9ogI+7UmnV+byx0sxeveBELKRMXExMhV7nujkTAUPiZWhpI5ac9
k5ovj6ttZKo7vDIv1gvYzxHEKVQvDmiqWx2FQ94IaTyG71OdNcHo1F/6P0XfZICd
KGE4sFd7AfNbLbbVMMo6PTDJ1qJW6slf8KHIRjS2dSj4bXdoPmy/11FZfgr2K7eg
l2GmNVJm6Tm3tarefuAX2zEk79inUJP1/gh3cSCdOcgXmE7NyjuCfoOgjzRInqCH
CMSsag/hZ60H1vQkCG8+K762zirQeoobFxT28Erqv7sq+eTK6qmd0rmEez3PRWg+
sOV5/jD35J83Z5j5Mz+JgCKxhX+gRLKztslFKMtCVqhtRTiev3cGK7yKESJHuL2x
vfdD1w49onu4zo4mb09Loib68TiOvL6KWVwW0OcX1gNDHwbfzN3OsYKxWOt8x7x8
z3rCoeBPLiYr97g2ztBnCTGrY1ZEOqFnbXZkvof6GEzBNKKTBqi8o4AeqYqKjXF7
wkHa6SZ+bT/3Ncz3FpwgOybgZIiyoXPchyMi67CMs9aYC95cd5D1DKrdvH9Ohd2V
kuiS7tBR3bp33oeNqLLzOkCq6h3AM4E+sb3UiFS39ASgaYDfky8iKRzVWbszKYP+
8zB9syw2lTgkH7ccKjVupk4V4tjKIta3gvJW2CCk+pNzqmTkFoPjJuPYbwpdXYCw
zhkdldJFJ6pk7DhbPwkXHU2sF/ecWYuXpGGE4k585N4yvzWNgH/DQvt5ISEPHr21
HHCWX7SuKJO5krlwwh7xQHcgqS8hBjsgZuwr9+CPFEUgW8PgiNMY7CGncibEbTXC
9cu/9/hy2WxQMfzAS9ZVKMuooUmgzYLnI/Q2Q9rC0/rg1vEM222WFtR9egXoeNuf
WtbMoZMtJsUvc5++Mhpf5r2q06DmVk+XIVtFOzSOqjcnhaGVmjqSAOzIWXb7ihdG
gXsOOQAsndJITHQeve65KJqFMJDpmMJPytjKTLYavLYV90p0zE81/WhebQ3W14g5
g8Pl4Z59WqqTaS1fimmXIA7cQ3Fz51hM/7GS6zKruX2jeTLWHqCeznPOFC+6uNaQ
ryvLs/VFTWRVc4MHtZT58BQg0z/C5DfiU668KjHY8QDrMW70ljDcjB24PbTJP31P
JqmQ+QjDROcJ+ycVkWArX748qt7/qUnZHpMcpJv0OVcE0o3jD0IvejUCRNc460DJ
unZt5Q4tQZiAd4MV7Wa1OtBdTEu1kYaVF5+rhTwoQkyPQHfpkeT4tkka+/Ecpdyj
OBpBnsycdeH/2JHZ//umD9/k6YHfPgfXHpJuCvkpP1d1QIT9o655JM5nC/Sr7RHn
WGuE65U+B22dVQeDIkDyrf3/O/v5D/3agYxLdb46XcX2tUbwDiSTktcP6X7jBjI0
5OX8tjXrQHeTxQz1dKPQRyt4SSChA6vurfSmboNtBGKD28ybUWn1vWDeM+GIrrs+
xbK6yJK5BJb2OAkmK5OVPXmmx6DOykUvxHkyiKYB240SrWpDagjf1RRlH3O1VHru
Nv0Jc/X+ZhNZOUQqJmkb31yKohKkI2Gk6p0rDkIXsh4coJ7I78cPa74yODh1AJqw
WnGa5s/4lxBWI2fq+Q9Wg2P6p/s0nBq0Z5HqpsbBxQP6UqN1ciE58/Kbu8Ks2tHi
1DmjfLzs9apkUKMyXl2r3eSst7XHC8iD6S37VER4p9/8GAq8DezHFNURhpgFDa+H
YnMxwQalUHh+UwHizu2CMx63Aj7RSBtS7d/aLqlGFt+oup3G6PDwtw9WGUeEtXao
/aMd+nvGZOF1G9OmheO/OYKjT8ONlT8BdObDuo+uSUNJ8mDz56jJXhREdA9KYfsf
y8pDXCCHTx1GqbwNB3eJfdUXGFVu6rhG9+Gamf5Vz3YMhAcrZVyLHyuJKxkJ61wZ
cdrBmir7qHUzTYnF3OaeOq/1HbxxvPBnkuyJS2LuWyioXWb6/1EapiQkbDw5UzQo
YuS55Ow56e9hz2Q/xpgwqptmmPeCmGaHPbJG+gxjsxLQ/H/Ejww2e1UIqixPh2xl
20HQq8KkclL5qYyFKsPab1S2TW8mnUZSmX3HSAc3gAPxjOJIDjWIjIDD/JQ+KId3
R7iVA3G0gD5Fx7gup0Gz5u8Op1OQQfcBg65/7Ki1VuEwHEk2i+lj+EUUCk7q2WbJ
dzxc5DXEdwihA/oGlSW+4yzY9j0sb5+bZS8wU1HhC2m3d4gdGDUUjlgR31igeTvw
ZB9wObhNjsG1RsWMm3RheijUSXWrv8bUKNU/MibMVSB0G70Muf09cIiraaz9uKzX
vDbANihZ340BYFDVlzh7dsMgYMsSvlMqproRTShTTGxEGTHzuPwzreDC8cyLtITA
zGzhj6Pq8B1QVn/RiKj6/d7O9yhYwG6eFsv31toKwJAFJWSZsC+ijvmKZQW9kcuM
SwfBK+W/WOd+d906s44lnOj72Yz+lFYibi3vNEKi17OFh3xO32MLZhSbodXvtS/e
NGYVIqjqifu9/e2BzwYtRh88ya/p6CmPH6RvyoXHhYnMVlNhGGAiAh4TJZn0SlqY
gj1Cya6bAPv/z5gmp7D16N9k8gCyYTSaT2GWhhmtlHWtJYuwfrlnnyFjPXQBgYr2
bdtfYzMn836LFJrQxuaHr3nZ6rF3zdg1tJxe3i/dfihguA/SUEdE7RHfulwdEQGE
+xh8Lym/KAe8E7FAOsjcAk04zuDShKNoDUttus6DFM1P/AN9WoM+DvKHSFFNK38L
szxzUspfNDTSrxEqZFIQx91lmF+OqS7hCy5I7GDSPmvhIsUYjZeR3lMmoLDAkFIY
x2VyY3gWQIma8tFx2VJMqgqbcBA/t5k+4aFx3yhQq7XHGrD/peVryqEck/iP3hh1
y8rG+m2ndwnL0DAkftp6DcE0LwwfjWwl8iDA/Ovs3uvkFG7e1oK0dkDBX+47CZQY
GeZB0PzBuGiNOUKui6jXlJa8MaZiP0W9nYPEtiB29wieP/ZZXivxCxwk4XozgfZc
mP4zLpoVOTQRCOhmKIebsM8EHv6GGBu0E37mrUDXHtb/eTwpDH2tc1r+fdshEEz6
HJdG2h+I+jOptqm7D10ccBZvozgjl067GHjhbmEua6o9TeecHtC8e26w/wKaBYW6
DGsdLcYoHeKI8J2N4TZLmjvtkLKUmUD+utOo6CcAw65YGxb0Ha6/8+HSGsJPXq5i
0LcRsX3eeneSYNifdrA+A7DFRxJ5L400Mz2jku0zehHZpbEazpSWe91LThe6nWrG
pJR/lOVfLTI1RNy0sxqruLvpEKXMAvvo5J3yRcFlqwPlp0Bw6Ut9BwD48+L5RJML
Zc62IhK17+aRFts97yGUoDyyb8m5wI4Myn4PPxBQyu99EhlwOhxZxh3CvTqMCtpk
qtwSBU9MMhehEVMmoDMxl2UqNgoXOcsBK1MCb1Y/uzSX4IFnAgJh5zzVCoNl04Nl
hds0W9r01t7jyp0tzdnMqxuoZoCfCtk9WOcY6TjwyPRgVTujT21Th3w7nXWHMjWq
dIdOenRNWHSQHn51ToboDojoD6Rty0UHW8Qa/F1ee232LsVQBqnFd2ke2cLo2TSU
er/FSXxC+TWW0hQIZTrKYqzFuH3gNk0jxDDpVHEupXsSUVUZc/QtTFQuuMN+ekHI
r1i7ZKkBM/RtP1pqGKBC+rSDyTPVEm3SVP+bobNm6wFk/5tIaeKg6VkfUu4ppVi9
l2nTUexBIcM1EWS9VwTIq7gwWbTTFMrsKo9borAXwz714xWMIEAcAaQyIQEiMA0h
rfLKYAgffqdQDCwASBlL9wFNhFB72AxhNkN/itlmVKnKDW590GRCrQKB4mX5o9Id
VUtQKONEMwUL2HnHlaJUXaxaCp5SuP7h+M1jvkFLP26rwGTCXjmxi5i/a+GRWq8j
fFT6sxD6KxLg2QahUdlBIwKk1QDZPg6T69CFQY1tJOjgbsW1xX+52Px0HHmbSnA9
jmFuDHJV3lnVW22cDvZ314lWVgghstjl4aZpjWMnbAE38dXA1znTwJecLa4O340H
t1T80suQVOuiiOzc8Ibz7p9TwWYqXiP7IQgRj51kyKLOvJxKL4cZjeC5rFk8dZCd
sh1Ao5vofY8BYms8UX7tvqyyyz3JnEjmJDdyK6rHlcbzhr7Mxj6uk3OfkLsG7V5y
ddGgLlbl74D9jQ+Rx2DxAZbEyx5nb/ZQL1hWOwOTFqdnzLVB8HWGMXUzyBIdel4R
BdKJuLiez9zgqgDa8r1x8pmYXgNqVDBCimonqlRND84a0RTUyK7/4kieC7Tp8WSp
Jr+L/g5Bd/IlUyPPP95eLTIMubpwabsNQkR6g8dYNcIpHAJH90aGo/XbsYYi9Pgn
OtZ0RYQU11Q/raODax+4H9Ce2DFO4RLzB+nCQ/ew0pDl593Uawek3xwuqsqentV3
bJZtOKwTdA6PQe1N7UhZV1Sq4L0cdS0p2CS745lRZufRvzAwQ1z14EaI5G5FgYJ4
RtwHAzhn0EPsdsuOzenXHa86QVz/POS7W46tge2GOfdFntYDJCC6L4SKePpypp30
trQfblRvx0KX1FhrsXN8mYa7asgrQQLQpaW8SWuHuH+wz75uwr/c9YXIX5+CF7E3
UcDGRfPCExfhH1ZFgWvHZ7Q5C/VyLQuAudScJv1/du5xaqMtcLxbQA8PmMG8V/2V
THkkOJ3vYWO/EUwuYB1mFPgK2LRC+oBsMxEdSA7eFSl652fW69HNi9hHWGpcihfQ
4ChEhUgZ/PEbDuBROrM2JulLcKScey4GAxhnEEbvIpLQ3W4fLZ+bz/VVRpXCkRry
CCjtrYuGN08s2aDCGkMVQxcCWOUcNK4j1kqtbt/Typlnk2LxwyNGjwbljJ5pe4p4
nMtSi8T7wGFqjXg+6Nf4sXQAaJfSFAs95J4OZGGKnymw8yTK29m004bk3VIY+glN
LjoR2R9ZPhEKr+8ckiIFrzCFYeoFJxeCaEd/nm3pNaITxSGSRc9tBa+y5SxoJKNr
kro2SLhefV5NsNw1KylMUzrtiGTZUt0BMrf/hjhMdNeVjLPat3yMc1N+ptNJfO2E
JZtlYnfXsiP82h88gHxUvyKnLDmFzt/CEa++c7gJMk1Uak+v3GBvl22ifpjSxLQF
3X/zt5452SIzTq9zHYufSzId5u67BIfWdJsfhgIO7cNOxn6Ps3KUEJpahHm3dNAt
ApqoMHAJxD7UdrzW7kkronfxX41n6keYghC1zkmMN5X2SwKt3ssU9zbClBkJuw4e
4nQaWykJYWf3gYGVjIwG8USesd6lDeN9Xslqj9+iznpX4M548N/lqGmIpSmu9Ye2
JRL3e61nWeKaJ7AyIWmPhlfez7CB3gHfDRyMA1F2RRsJ4z3IW4Rcp6fGJ8fJXnAk
asBF1ZcV/7fvLDa8hp7DBb6LONSGieX+++SbwdiSTvAztPqEreCbgBfrfvVJ3Bgb
CHVKiEj/55o6X/sL+5FBVnR+A5rz2JITww6ujeeq/c4tNEeOQPJ3c4st1hhmwMsi
FHm7YpUiKYIC+ozq+VWM6nokOQqJnxacBDrA6SAldajRFp3U+0vASt+i93jZ2Qgy
DL27E+ttPb2Ea6L7MWjOX/dvyIq3wXROUJvB3vMpLoQfAoiJALGBQLrjnWj15wjp
qzAI/IHvqG3Yj02AEtr3iJmYAe8UtQUjheUJ/1e1TOIAC6R9mQl2uz4O7C3yK94x
7KQOXNyxe0v+8kFsHXayMkVuabXfX14YCFbk116L8hA35BlbBHEvZoRIrAkt0iPe
sZni2kXYWfGZCqefkERwmKhowxjV2pqWQA9XZSHLVbItIJYZwq25A/dDHd3m2lTk
sv9qXNSttj7AjltGAIYRXWwv8VZHRrE5DxsXh8oBbyCQcoC+M11yj5iHvpnX67SX
XapuFigCYtYAyU79XDRkwAygQCXRCfxvyDP2fWjqwf9VYfeWy4qnD0GOQHaNhzEI
Lq3Irhift4mw2M7EMJK97HuxRJZ8cIPNcvTOIA96plTBBfizeb14jW3RRLBHyNgp
0TodkkDE6Nxpk+hMka81+sR4y8bjqYKbosBCBnujSQkpVQ4CT+umBdZoLs6NJ/ts
V1614ZAspWsw6aHYOfRp04aPr1ePhMu9EFwW2l0iK5GCS/h0AVHcjptKQInta4EF
+ohGOKV3xSMHWDTleUnpoWhACUuFo2vFqN39UsCszWgkGS/5VW6osPhhD/7X8bPz
BU+Onlt1oqNI3CGro2OAKnr0cpvOVkvHYXbSkJlV92pP4zeArTKzit0pC4dqgXLw
NnksAim2G72Tdq19fo1gNmjdfwqBbNv36bs6VzUtzYLTHUV7zh5mMxD7YYgyPb6b
LcbHuimMeLyE7Tqwq9lZhQzsTJe5f4Ik29239XmhpUkIX227x9rs7jgG0HHOSaXL
siWTLI3Xfkz6iL+0vsT8aM1gOR5rhuyd3p0sQxXRGC897RJHTBGI3e8IGek6mLHx
uL2hjTCKJJ82ttmfOwAVqUIgX68RvMzqT0iWLCBJo1Mz9rnApR5hrkaDspjKD8y0
j7rm/1fEQ1/c/DyON/quQU4EfgDp4NjaH18/r5VvqmRedNEFv/gKL8uHUFcBP+nK
JK/6+GMOuH6zLB7TWCamqZ6vwfkJLJkbinqmapdH62OkScb7RtaUM8zJ3ohSdHqq
PgX6V8YhhVFwInBj2rOgtpcCwfJlXnbipguyAwF7AfvoEhgC3gS5ocg+0cqXDNvP
oqdizZJP9iYVo239JrQtqT9DlrPPDME3VqedwFoNvOxEuOtva5R/YVBHKN37X+cc
8hRLwaVK3F1mmi2POOkOkTiYSEdUCqE7UEdLNPuCfPjSFz4C1Qu0yZ0VH7kyPyEo
j4hsqgFpVundKQ8ffmIre5y0OMxJUAXjgAPYVub7uchmsoXKd7EzijYv593Of4zi
no39Ui/ToDY+VdkaX6tITF9Ypt/ZFi1c3rE09NNmxOVK9FaLucRL5ImoSQHgTxxp
MMs9HAtW0rLGqijFpDQERFJBfmd3QE5s/+UzWoOd7MvTU34voA81L9F80aV1VTH6
sDmBzvP0LYYLdd5uxkcDrLBuFl382SgzyOW+rCvwptiGfuE7z5rdiJzgb0rvvjdN
aBbjJNBnv4rKlaxxF2zV7R8dH050DnaJeqkc+uQbZY/bcU8gB6YXPBi0LhxSi1zE
YMEGZQj+n+ndNog1il52id4+3MUE+67fAUtQywA1DUg3PNMZfLNJaYolyyCVD1TZ
UdejSBkOmUlCbeC7qxdGrmqMmqe4qLlNmpSkOeKHeToR50x/OI5HllSLHQItqkVg
6M11eqjGSjDbcy6fT2xRMmyMI1E5YrO7M9pXhR4JmFWfSD3xAUux3m+zXUQnYXeN
S8tIopKG8pB7QLGxn4GgkpBeI6ED/qKXh3kW2npFAm6S7idGWd4gEKK4GuLi07g6
ak2vyLJvhjzIauQ9S8VDKGLTCAtudXiXgbs8TnP+ytKVZ12Xw9fA4QCOw+Hs5VsV
6uW1RsdNZ59Xoy5zdKbem/sBRF3iDjEdphVCh6Vp8AMARWOPGa4E6eVaeXGW/M81
X9Lx3LcxLL7ICKh5Hzw/S+8tgrv+WEMnolqw/p6z/Fc6ppLbiZ2bpw7LNW8wlBJU
7WXzHzUjcdFCYU0p1Svir22eMdENyOz5HjcaSTQ4FArQ2yFGY/M2r5C+aPFd5bxE
0HUDd42cQ1iTAbYc6qb3C4AfkG/ykVmHVF+nTu7ammTzRTXENrJr4r06I8Yo5Iyq
yDX0E13/BO70OGt/aUPJwWS77m1Bc2juL05HA8kwNoifyaS0f3gWEHktCsPcgVo2
7o7hV0YXKAcwJ/U3h8SnV7trg/3eWNbdfRDnVh2s+R/xfcvZw5oEisKe0v7XcsQG
BrRD17yf9xwkZJiQL0FpLaaGHIVif6v2AnIzCuunH05EAKfT9xqivjD4M2JG8Dcw
dMC88Ads/AEVW4vWnoq2YkanRQVW29wWEZcO9rrx3y8NfvLYa0cOF8Di51P3kDgX
4GdM+rI4rhJiI+nHN5xrivRgTfnaFscXigbthPfMCurpN+8hflG4zXKOnWsgnivp
0oY4zRL4NqAt910K2INtUgZp6sjp9tehYUBRzE2zD5nik90xKftTqmwsD/iBSkya
AheOuIiEosv0Ql2OFuHnHatEICKWqMBWVyedj2Qg1RGSMuYDOEISmeWB5hRZertR
jGAvj/mkcCajZTwiy5avxcIVo0AJLvPhREtilvqceM3Iqj0+gfsAAB9uWpkdNrBz
LKsepvXbdwo3lOSIRlFOxR6ZqNVvjc4ew1fZ1RbNQSWdbcvDE43c0PvMKupULriB
swAhd7X09oBVK7v/x5mtgsiZEp0NOHpahex6L9yLvAs3XG7JHbMRGAPG1kGlOsbL
8IhHBdOlO8DQbMXQvxdXu+Sctd2CjUAhHTaWzNJ+/0O9NwJpBP5Lqz0Q18fF7C3p
ZviPyvmQmDC62jd/mIu1P+TkNRK9YRHINj9kjh3iiLKUR1h4bPy4qlo1NTtpGPjW
SbNKtkcsm+WHYbek02hgaRa/nS9ZVlc/U/15Q2fm5oz55GU2SzlNhIDQAgL9qGOC
df39pgGx730or9hkMgJz4eY/gBKjfvESvS5FSF0RXuvaQZ4bakStXB9uYKPx6cNw
HnMZy6D8Yqq8ItscnMGK+3sWnCO2V6p6WiWmmSS9W/vq6zNldy5+JDiEwVKxoCMS
JxP1kThCkisPICRSyUEpj1Y0MAKJZYMER50B+ZBUDCcUj2+rhlSfheCrHhCzaDM+
4Zj24vX+i72YmrICmR9gM7BGPZFKykpkkzja2S9UClMI2heXT4WZFqD2Jz6VQqGN
HKJjN8gwvNFCaWimhp7GSTs46IVWhZeK9BeQcR1RymxfK3Xi+l2RnIuEyQq62AgX
tXLzorixyK0EzX4v2HUj+P7iSaGbEvJNZB+fxbvhBDMOCTiZRbfJGoKSYvAKun+i
Ck6MKr65rSq6gZ7mODvqnSFs9efWUjVH9FSApeMoOlJqNgtqfEF0H5e79Ac9rcHb
QyfH3O/IuRdrX64q+KeyVZRIT8CG6b8Dyz/H10kLxrfZ1qS4HF2L9hDSa5NPPBDY
0T+6FfX0SbUlhcx51dR4fxldtDHRcAdozzYR4uxNbiotcPiKnp9lyEOrXFOS1w6P
XgYLHki26wnNNADKd1ouQPivv0Eb8eCnShv02MKCwZ6A54+xNDYNtEJ904TfYq+Z
lKYMCrAPdmD823QF5BrvzlUW9HSP2fzuzLn36Eo40MKGHoijt1ryR7Qi2xqGjjqW
spFGjYAhiFd1NkfXnDZp8kPECz84w4HChTNXe3cICtYFW3cax41IjMyHo7OYRo8Y
qTm2VaP01o54r1MQxOUc3D8QM/RpX3TGP24faFvBrl1YIMsDs4rSsA3HGT7SKV4P
AoR+QE7Nh0TRN73UMumDK0nccqh3y/U6hzdQD2M89kKjN5DuHxkANpsAHsLng8F3
NO1zWrcuFaHTaq2nY7qknCJ1Jy+93SKCY8SepjFYefYCsjs/MY+fduzkifL6xzSx
1uiFRlEEFOfSMqiMkRSSUVFf9BWTIwXvoo53jztOOk32nLIkkyZaPY3k7ujlAtnB
rnbQ+s3Bc0fAAJ42jxl9Jdvmj9yR3F3f4FGKfTSDNMY5Za0DOwdtk+X3r0+NoB0g
V+CPG0YpA0lohWv3VAt6RO/lohOi/NhBbZWaWimg9uPeAcB2Z2XX6nqMv8uBywSY
yTwPiIkof1KA4I8+Xg78xfXdvsfisSBQ+w4EhA+LRzOTkrWebXXecmhyjLG2hb1A
EOulIbnnIKUwpOnlTxi7z3HILXMbamuIRLeskLOUI6q7VwCQjXmfrtHgZzvLT+9u
06VCWiMo4ryTHYZMYEScjYQ6DH4/MCmksyohlRvkSsuhbqP4MvyDooaCe305v4pr
KQ14R/okPzq+3a9x8IGv02zQSUTYHmews5GTxeMsge8m9i9PvN21a09vrcWInPZK
YUUQcvA5jLr87ofFBaa17XNlY3kbAGm9JTJXZ0XcIVCrrdsYsXlpju6BxHh4jE9Y
Z2Lc44DbB2FxzA9L+4/SMHTjXC7ePc3q2HMM8PZOIRdnnZlZdiXSFHwlnxvhWI4y
hM9R0kCikvfy0r90lHfPhWrMWw3BxAQcPbm9+DLR5gajlQ/LeqpXGxM6tP9RuhQK
W1kPu/1+7fGoCTPHqPMLPeBVHRlU4MDM7vXbIa+SbJ0RznvGCGaReSeQ3EmVeNOH
O8Lfqid26vPUjdRq3LfzotXRmrSCuBVS7CGj/WJXJaR4EP8j8zEF02e8/SG3egQa
Xyt3W+y4f5CloNO0tavQ0ACzj1ABEnFOokXcLlpznm5EHGYr2e9rkAJaWKA6F9ef
ngScfis0yR5yZALVtiCBLEImzPcJOXUOeKYb89Cmyx7VAnRquymWvYkcOlt3I8R0
Nxa12V+xctkxjFJD4Xo/Fx8r0/cw2H9gySRi4MqkYzj+eRW9MUzqY8Qlrr6rupy9
HxtlEmEv5qjAGosjQXNsU5nVAtYtVPlsodOgG2aqcmLrl1V1ePGK4wybQU0ciIOF
46riTjEz3/bpn29UJ2v3qw==
`pragma protect end_protected
