// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 14:01:40 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
bN0RwllSgTX9MHiatJoIzEvyMmH4Tf49nm/Zcf1HkENhDz3KwURZ1aHwpmA0FbG1
jpzVfzNvxClMuw7mVDJjABPVyOGJYnG6C69sJulr3DR8NXfdzOysw0HsUnjjIC6B
FY05VG62QQHIlbEsrhurX9prE+SFjPWeV2cwHj7wmXM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7920)
cV4bX0AQOhMTviXtFMPuxdlOHjTWHkhuVMaNRCUKkgbI9NkFjUJdQGyPrfn8AyXB
xzYgi87JWL3l5DnuZXehNx/VW9M2HAKbEhzAocqhangEwQjC2vPF1bxPSLIHy9Id
CzMziC3vnDi/KCVlzPFwTh1CCBkyvvAGorrZcwpM9G/e6q4cVO/nM7rJrCQuS9kr
XyQ7ZtywWTRAJFpfelG1wauD/X9JDRe+pTKmhpKTrPixaE2ry+OQDx3D16okZEK3
O/AMcfc7aojAV32EesMhj90pH/vx7551yucv+JBgQtoDVp2X/Dp6xgbBiFQ7qrUs
wjH0JvAx+YD4U4b6ZLG7X0Ko2KSs5NUKd0Dn1tgv4juDRG48m5NH58uVWJ09Ozkk
eEO4oObpByfKzNxRgfnxMm2ibwbvSh+TKkXBwr9/23Y414NbmAxRBaFZrdIzDjUc
cxfmhSPraRAU3t12z1cXets4SNsqNQUBMRnoI8WioPVWGukZYzyHBTGLrp8I6tvf
BHbv0U6frKaHQKxc+lIPmQAJiytjs1tzJTzYVQ6zwx8r1PHVuJ88o8gmKb/KxCXm
Jd7T6LK0iUysp4searNcIdfueX2wIWYiui4QbbHYZ6bEZO0KS2xed2BDWxuabXvI
rcG9owrqKUOmqKZmS8AnZHpfCF/Gcq9yuuuDBVlZ7aS950K3CpkxydXNEp/k8uv4
F3L8x2GUENK06rryKD1AkAGGe5nXe9ARtWR4jJlEXzl/VfjMIOcsFF1OxyxEmZio
fJBKaJ9oGf37nYIReCQ2p/BSRF9L3OA/Qmmx6PaZXMOuzn8+zTDEWFO/rLqldnQL
hferThFDvQuCVcSYLIV80EyZPQAZ21SmsyotDC9WJgGIE4SVeI8l/PQnlqfYbu7d
c/dNyTvXKrksCr4j8knTXTUBY61mEtKZ10twdzodv7vCCtc7XI501v3JSaj6cPsE
BeuTL9/nYQLfEoS6L1XKfkxbSRs6y3ifpwVGD8MHd1fWcrqNyAFMTyqDgKQ2bEGW
BEBQhKkS9aPlFxjDOupX4zeHvUlCFUmIIMyoSIR+FngGbNWFBjxeosuACAPWv0FE
taRuN9VUm4DEnKnkgvYg72l09Ss6KxwyIsh7dPXOA78dffY5UPLCEZ8oMNUJc/Nc
4xWLYkAFHK4vYM3WyMtHEAcr5bhgmf0wQZbohirgtDO7kD7fWCAMXkBMkXNHdFDq
sjDAOy5zNQPECUExUuQnMRrI55FEw2aNa+/FbNAGwBMagL/TMwA28QlRPlvo35PA
qFRRVU6fsEdETqz71nyk/8zHzz4NrY4hxCcrPsHyyyQS5PjGqwjL0t/9TBN+IcLY
E0lQOz8/twKKlAac9wKOBZrNEeE8nYEQ6nfVoyKFkeApAy37lXe5edtePIrb9yT2
AO7EsBOU6m6FcXhLkU+ManYA0aw7CDm1x0rIfAtAaianmagQjlZEbZ78l+mb2JtZ
k/LvapAIIa36bquoDu/3CleKWSgyNTHt3fjzYV6QUt3FJShdHp+SF3oh7SZB7TbJ
BfSIu5W/F+3d/PyJC0BiRw8F4fEpLBa7NSpggmiDrS+7mTaxxwsKawKDwqKobzyr
IzjuYBym9fPZmv2eUx8BSj3xR9j0N+vj0KY0Iu3cjrSkqSxlIF4LbNMLjrHjf0io
/FkK5BIp63wKS9CcN3V70qQ5QnNCxhd4OwQdtK3RI0Rd4/v84Ymig2i0rpiYVDqV
oUG92VjqYatkdFMDgduggq57Ah6+PV6Og2bAPVW4t3lhqLoW++oiq/S3CY0VfWUy
PLL25C3lhqEWVA4q0zelstXVC/SB1eYgJnaDNsA+mkonngmbFMbptMO6WQ7LjEZp
t7OEkhPe9RFmbjnDHGEw2Jw/0HQP5Y7ZCJWMKQ8aVWyGaFa4EQ97C2E17luB/qIk
dWILuqNl9h7/ici/efw3bdO1Y60MuHnVHLelt2uHnrgROP4NcVda3BhMTbKOY1ZB
EgtzP5SYYQCBUlYAoT3BbsIiUXetzFVMRtlAako4iZ8M9KovS/ZYG6v3PxNcBnjI
Zg4HNAYU3USWqkR+5JpSwjLBLA5pl0iaQno/OpwWFxPIY5jDEKOSwuokx2zOk0IK
WM+tvNkLeCUMLPsEUuyfsj4Eryqa175aYlIG6k8I6zRDFzkBOmvlIXDSmLwIDvZJ
qcWBFLS5MtL3AQIhECmqHhkTs4iJrByYqTHy2TP+ytZNdiWXGknjOm0okUZu4Acs
UnFBGoM51dWqk7Dl4PNKb3dVk6NZDZj9IsvjzR9s1u93d1L2fDnR4O2GL771PwHf
o5k2EISSXL8eaz7mKm1nFPkuIcIT1S4N1hFpOlzyVV1PRmO2lbN28MWvzavq8na9
nhzJCc6cpyeQo5AItq/yI8SSTWqYYACKK0+49TN8VnwAZ734tlqTv/4mFvOFfSAy
igN5vE0q+fifvef6345on7HsGxOUwGznOoIzD5/CWxROcFWNJQ8vpLnMzkb34Rer
Sgt2G7UpXfrUUm6u1MpwtIzPQ1DSLf4ptDBt7d/A2tbC6wagmJ9pJ7y+GKoCv84U
3uv0XuDstDlN/p7jPEjvDcLfqabuQ7PytVGK3pEY0HlPiGB11c14jcxa7qFbobq+
Z4zDAlzAKfAbXrH59TIrgP36te5VzQ1B0RSP8UQf6pEFEbvMMF6XYy5dQtTgmoLe
29K9kWwy2pTl9kwchd+DcilbtwAXSuLyRfp7bE0uPPo5FGOeO8L2de9dJYco+lGi
r6UVykkwttDfOzcL+lNd4DwRDxxcSr98DpW5klxebi7fzRfxPPXbvUKSdsparcMA
WOFVAiKFKF2sMQLWy8CclSpqtXLUpmyYexkRPmetVHbRButHmEgAM/IijJWfbkhv
7Aw+thn1kGbmDFkqH9c872gEdpdwwiOMr+zcd6LZeDupuUsN1Z9Cg9OyMuPxDi9G
aDQVQ7C5TASX2xv/u66s70VatxMQBJFfxbFNZiE+mvk8WBQ5kgQ7Fn9bGHYO2Gib
X+rg24gmkGZ90TD8IEg9FFVvrqIX0790xmXLPlEdp9EFsi8CwuTuinC8whHnfh/E
/lSSxSM+l3ASH/CS/se3ZPa8dbVMKOe5572JNSBzDPENkjJBC2NC/QowXdNgeljk
ezYmlGx1HR3uPG3JFf6dbdlfFTrKcERi9jzhHT+yTYQkybt/SwnoEw/9TA7HwLC0
7BXHigH2sKw6AbSVGP0lwtGfRssFowScrk15hdJpXPKSzUKpsOZKY2zH/gUNBrtB
OSPntFS72Put6I0uq7YeGwU7N9jUFbXnJ5ZUBqyeF+apv4lVIYxl11g0WkoxgDMm
c9occfmpzFO6zgMqR50ZR2CIM2BXK8a1t7OM4Zj5gSIIa1/ac27pbJXXbJE5UfCK
CkVLgnfMNR/pLfgTQBsHKSnkix5Ejotv2+f3+8ciYtKFs3zM5SfDHmuIpu/wzgyM
BNPe6Curh9pWa35JLFe5UgN6tejwiZYv7zMIinjexi3fbIHy2l4R+1U9A8HaqS8F
evZNPMusy0LL4fQJYSuudJI0mkJ5SzkZIlA9NCjFwlr7Wks3zqVUYuxaQ0H2gfit
1nTzTH4ez35vJK2ERcrv7y5SGsZIZVcJotbJLo5Fkef1UCWnSaUzvQx3ep78B0Ah
k5KYLY8wYT3DxXac8jjC7gNgsg5uBhUg3WLSxKLc2ZcK6HNQilgnk3cYwHs7CV17
iLtdX63/UV2ZiBurDZKj02fkjLDoIbasSfW4G5bhrXfK52Hg5BfHCRpoGBWrckG9
cf7qWemb4dao21x8GUy3e4zblaiDrBrBO1Mn4z/eXL6aEPwkyCFRaqAJU1Gl4vWx
GnoewDHCg7tibT/Q1UQZjHTYb3tpvQNOx+lmfJqn5DMAB8ZU10KgFa2D+DC4dLeD
3c/VBOZWJp4mwCk/x6iCb8f5z3RDNhKzpYx1G0iFV28fKxeFH8XYYuLjzpmcu4tM
df+ZiDKhMMLIehXGlTo6byYF1ZE1FP6G3r2b+2j0t/VyFqFJkxxoq4NOX0Dxc/BB
ECsVEkkdUaS0Ssowne+6jo+yDlbg1OackCtsS66+tP6r+xzbRCNpp5WAYvmQzfqv
gDKIQRit2oMcXlh94Z63Ki3V+p282bIWRgvNkuAyUNvtLaZ+Bilm3R7vAyDXZKFe
UjMNeGpOOVujTgcDkXWyT5/ylqwTRdc/cMj3GmL+WNTIXBhxeFGDcC3QluasZ99A
tjbXborZN+6jkUWPNes7Yo/9Tn2z4J96DFw5pqe6jA0xU+Hli4eWKu/zP/DpRJdN
83BBWHWDEn4HbIrLAi/fhLoY6gMMA7HCGfwWLfrE1ZdxgzkzVQRqTp+Wr8+FrGZa
2dSRlFFtlStOmK2awl/0lSXzv+vm4NEkE/BpEDZn3zgQN141xeYWRvKB3Ln9WGWv
b7gmfngsQnDPVtlJVgyme18971mVeT1T09g3L/OCMMbXny7zGcRbngeiazm0JEaq
FBN+Ii8KkVNxpwNyuDv8Y0bnaH61cTqMc0V3J0UCmNLZoQJ7TVI6hKbUf3A1jCj8
rN7gBU8auEMnMaApmYDSd19hcUXpQKgHxMJOi5JQllQG4nJpDpNeWVq/WSxcVTzU
QDN5CjlWPajifotR9lLqt4vf0NqoPqAEHIaVso9pebn6y2oxCHd5xYN/BEEiHBGH
ocH0H545/P35Upv3GKq1MPF+XuMwr+YXoq+d9GgWTdUdqzf5M4NeYxv3JHpOU1Kj
SmgaieytL1i+5omS5HysRUYiHBv/u4WdtqH3UBmHWBxeWq43+2hLRo9oPOt6ikwx
mQh+IS7x3J7+JcnR7xBYl/zuEEKX/JrMK9K5tI1XTFJSYOK32E8xU4gZ5CnWiFQi
rZ4BejWEn8T9NczLdLwdESRuFPNvJesl3XwIT/YKwrIAiQmXZNISSa9Ws1sO7RCb
1X0e4QZcSpfACpg2TUu9K99/B4oexXWTqpWA0bCgXIZ3X6fuTM6QSdc3qu1Jwl4s
GIFBa8AcihgbUhEJOcStqzCgkC05Fvs4jme/T5LZ+pt7dOH635ayq+x5nX/Dk0wT
LBolfWRBh0wjpf+4dUA1oDhtU32Bml27fhKzYyt58mpMZoHUHqJ1iqG2t4upYXTe
nvO7fX06Sxh2F+I+rXjloTnYgOFg3xl9p3H2WkhWgQsGNzOv1yxT12AJ6p/dVxmg
NzfUYV2D+3YDiW2YNlX+m47fnQ4OVDWYkBhpYpPRXpgdDmCJ+/WbrVkQN1mK7Sdr
pQMSBLzMzOhrTcVy9wdZJgLKn0qoKRSLZWP26HaW0qx8q3Af6Iaongx+/9GnVUq8
L5yWhkmzY6oUY9dVuQlaWoDFFxPVdlB+jmKiHnOGYPmC2fqZ0WknYLw4/JOc33Bb
aAKDJxVawHmQtR4WFYhqHg1oCsnwAypUSjXCcsSdAM/oVN+rzJvJNu89icj9F0+b
7pXrBR47SC+NkSm18oBz7l6Xb8abOqtcs3TqdP2i4/4X/hPhfUUr+jtbQwqul9vw
w8tV8gLnZPADQoHKT1zTtrbLGpJux1CP3s5u/yRYeYOojOo7u2AvtcIcJEWlxz1S
2C0X9X4bE1j9hKc3cnM+9BJln5r4cLh0MyJlOgaIC7N22Lbv4bpq3UlibtJnYg8o
zGTOyHsdSfyOLZqVD45SQvvxytl6Q8iaTmD2SSVOLl5yL/vSPV/LtFfRZnyj7ZRJ
VSkgfT56hrjV4KPKuweh3zpCrtO3+xcNKWkiogpBYFJhYqQmWcwGpHjEhLeTJD4A
LKcLgkuUhPgmk8Pp8o92wsyD9HzutM2LK+VkHAYal7gedv3oUzqKnW3MAs5dyFC9
ZCB+aFnfwJXvhMfz/HTVKDEfn2Qx6uFytU/C6+bg3/WEYYbRE5Qpy9IO7Zlcy/nM
/TfU87j/8YcQACkADEbkN8/Yyx6IbqYwEspZW7Pvm8pcDyYnyKFp+7Wmwgcy6omh
mNaVQGMtEI5muk+YOlHVS+JkEvNu4LIky3U7fjqbHfmO+GyATa79W7blZ6uZJ8E3
vv0p3xWpENbuJUkztWEQ8PGrVh/icYa4KUx+j4q29oTbvyTnCiXUDQEheZKiQpFe
7GvtZd8WrGm0k1n6ZUYjoEnMDby08i16B15YqMoIklZdqYRbsJVuG2FaPHYB64Nr
TEWm2YT+S1N0ndESY7dFII1IfiwId1J1xQ7pKliTDh8HK0F5kl2zTsIbhS6nwXWX
iHh2rOXAP5et23UpsD6/mGi+/RvoaYQwy7Mn3JT5Z2Tw29HGxRAkqGowChmgwl36
Tna9TcmVy8LOwbaAyyUjTd5P3qAf47AGGT5SXmBCMhmwENlPe1mywCEMG5lWiZow
mvVE1VnCfP2Uvf/D8oiY/2AYLjC0qqwoFp3ls4ps41R5u3XbVvDz/WVnKGDiLKn2
Dkc1yr/9BhFtbZ0VPpeq20QM1c/i8B9/uoFPQkVDOwOTPDooabMMlCfEAo73hrdE
rIjZXbQnFp8UZeBkGn6ofYR97kL03T5X2yljnoZN4sGZPMO6KIjMZqAcPh72Rmb1
y81r7/7Pytu0Q5+HN2c2azhg1AOl56dcqxfhPvk65pFQYJge4OmWlIu1W7LIeClY
uBCwUCABbqo758+TPpfMw+QQM/FpTvf/rQm0W1C1XUqPZUBB00JXKstSC8AP+MPH
cDOKDjcidU+9LLyXM4ZIU3DZHjRMDnKajeV/dO+e6YeZH94S41gnBXTuzpAyK04B
Ve7a5V2aGfujAc//VD1EJoqWvrZCFZaS6cJTPzegseaFtu/KaDWVQ7+TQmfFbBSN
mTnVqzGpgOqTffgizd0oghixTRyT+k9c+lt1d7Ezw7W+SB8OGwPnFdn2D8VaSHHM
cryILO0wlFmAzuLdTBaQUoxXIz1kdUZq8ROF7DrpKLqv3zVy+bY70zYMbG8odQqY
yFnyvefMDeNVTlXqEab4QbhnyGXqf7+LIRZKZTv5Dn2fcRicGxAl0fOLHbz0V2+l
zn/JBs2533uO+LyFd9HqLtvmudVcV4QU1rw1CIjypeoFnsCo5HGf6U79kzXOmStV
Ev6U2XioptTHl4N8rFMr0jBColi4+stBKINhE2ydpLSQN/HWCIHGQIWdEp8UiJMN
+KXEnGK0S43+WG0OK7AwvExG6o+ufPUd6/d6DFHWt1uSMRKiAI+s8QyAGhSOxmrB
3jBN0+8OqvzzOy7D/j4H+iskc8WkyjAgx26MHnce0OAXIiZ/+Z2Idx5jfknE7cqO
jEc1jDBgtuaHuFaSV3nd7kkVp0TBuaE5O+gt/SIdXTlXgYXup+eV1luoHpPo/pAD
4b6s7tz92fe88Ifva3/M2539WfYv6sSyTV7u0e7C238fK3bR0t/tXM1wOGjburfn
+ZKlmg3XmHiqsBDZw3J1izocFOInPqGUSr+zYqzzXi+Z8kOgecLXmeuRlzYFurcj
xYz2Vv+SwFtw/eTALv3XgLVsKKtQdDrZBLVfprOxidmk2pvJIXAD6souF3HyJlJY
DgVtPIrDWcwkhHBRVIANSQ0o7G46VZwsF9Vb+fyHO3XEUMjfnHw97U0X05tO/KaX
FJ/tWhsHo9UY4wRl4GrO3LDdH57bJzSN3H8UKuNAcbK4N+9WzfSh8evZvENiyZuw
7zFEA17a3kzNwBXz/rTpyUJfn+Bcgt1Sneg746O/zxFb1GMjrK+LFIwwZqv6oT52
zpaNMePc/d3zxog0f5k+PA0FC5yNRsKDUhU6woHJccSzwrwfCvYdtm5eKXca6m3z
dfgi0OKblqkuTcmmTE3VveIF/rn/gJtN7SaI3zEpW1hReJVSK4ucu6QY6mKVCb7Z
hGioMWrbtZEIbcW7j49B9vql42O4VtYYkiHTLo+RQ1q1lmmNayQwcFTPpaZV6FPu
lL4FQbw1tKSz3ZWyLImDtpvbNsqEFbSGsYjL1kR+TlMpXK+/2n42YwFnQSliBofL
mTGJmNn+T8B8tCwThCpyk7QebpcEa/ciE8EgFXMWLn0sPKqxMMiOJLuEqu189AH5
ehCdpRFBcchXoJkzwg22ULuSlBzgYkBant5J/A1vyYlzVkxPum/by2T48VPp//6d
6ZvudvHOqH3KFmGVfN1nmXKx/lHHX5EaQOHYRaex5YCkPoRBz6aKCs8wzHsOIIjL
Qv0vh9sS6gnCZ2XD3HfOSANzFtbQnXV95nfoqLMAmbVzEae/S8I8CiUqhKQowtiC
Ao4gqcZXvzkugqiJmLgCsAtYBxDOFHVz0/qO0VaAT7wOWXrATGw3aFdiBeLD2eW/
xyrg8P826MmsszIq+ZsTFxhpV06p3j1zESBQjO6wYb0WJUrDbORHQHCKyKBJhNl/
VMfN9zjXzLZhBBdxqFfd3VuZLuELJelvfyHfnP/CHrSZoZOyzArA17C8qu6DkwAY
3ysexoboZmKj9EZoHvfeuUKpQYXf2tNx1/PnWDEQB1F9BPWzm7geN0yCV20RYh9J
Sz7HB992yOBnNSBssNW5huDnBoWugmM1thVOj3khj0sMcMHEULS+0xJwOQAlFO++
x7qLiUlqOjdeKAydY2Xpkw+uHbiD5iREYFNVEc8aVqfZuqGQpk8umtGh8BGwAGez
1rn294rq8FDx58iMTnQU9+irOgHjY05huCiRnc5Mj8FJS3WS07eXiwfBfbYCTPW9
x82TjAc21P7o3vZ28kVkNUZtTSr2ZbKKTa+MZH+QPXqwxDuhtbDmkrchtXm7Qunf
imXomogqIs6BflqHMAGAk8MEri/nIxMXF0RpuBsY2uA34ujPserl52M5cYq0TOot
0yS5CtZYPDe3fohS4nNWOHxzXV+myTdTICZLb+703vCcAbFnzQh6n+SOMBdCTlG1
/njDYs6OU3SRlkBptaipdUL4IwXD7bNw13YyfKdkYh+jUmMdHHdWWNeqCJTisP3F
3ncwfSjg6difbN8uzeeqD8nwYz3trMSixh365oyxQQ6dmq8jMURhcWEeq66OaIw/
dgRdHyuRwiwyopK9cG7dlCIxtsI8Rz2zQI33RPmP33wqBHRoB5J1uLqS03ArYFzY
soAoKSNzKEu6gZy8ZI9pZvV9C2NYFkPq0Z2ERYgoSDehQNYiBoUZyJzv76z2RmLm
f+svgOinfWsWWdbJXzwGt69FKUw9C8L593wlzGRJnxjrF6XZPGbPbg53cVOm3yN0
BKX0b4Sdcpx6dMNCfVxcOCnzbImQk9m809Hx2I+mot5T7aizIZVabMO3f2WYKhwI
ffY06XibrKoPqgp1m1gIFhMTFXvGLjYlnuPVM35/9Mey89WLD0wJQ0oHt9OUJYyA
CLJMtqugclvGW7UxT3jGpFmvkgxhBcarvW4wqIXMMlb1K6MKG9pErNQrDcgifSay
R5cWp6eC9gahzAuJFgEIkWH+EQPkX4kSYw5TaQ8D7jh3a4UTgtZjssjJ3v1TZ3AK
Zd1s78UaILS4n4Yndapsud60G3tvuFxkF++L0zj5P3rHfXFXCVqsaDQvT81nayYU
V7fXbPS4KzyQCdyJglDW428PYTQk2raL+p93iLCyAR45brm5ycfzCB2P4kMgKgTr
M6hlCM876+6tn2YxiiMOlRWHKdx6mUBvvHRQ2pOn6HgsO3TsA9ft4ORZB7Rynn60
mYNzD226t9b0rp9r2FZH3l52uWzf5l11ir30Ur8z7A5r8/YogfG388p0GojxhkCL
Fuo/fOaQ+LXrKc/xQ/qIhHXBkeVu+eGQlNu5C2lrEqTQJDu0DpVIqpklh2z7BIpM
eURmpFU7PlYA/T3qBbkwjBBaeREHB3wg0O9TzqbCE+E2JKRjjgV87rkXi3NZHEDb
jIgpfFIKCleVkWhSCfl+DIEZZWpkVBm33wI7fPCBKFb9YY/363f105lKtaZ4nV/P
7nxk0YfVIg79Sl4lkzwUzVEek3RQLesI6F6uQAnJj3Ojm68+BCoOrR57vNukbHFE
ftncPak6+y5Pq3PMFX8B94PHkfYHnQ9gIz9p7Wz4+wKV89chjYR1rpEqvHq+wqAt
0oLrVE/R9Ldqt7yb8yjdTSxlMzdf/lQA5ookFwD57kx5JR7QISkc1W+gHjFVJMDF
oZ7z9eY0aMOkEcSd/0XHLrEWZ1Bo3VVMqJ8DcNLUiofFUSJD8JsgclmL8endiNGE
qA9ZRhGaqqVlCxg/5Y0y+rjiuZQ0bHYsC8OvwCKAVjG90ptg1byp5tKaGHtfqRpW
D6WpAD5iCBOpthMcG9+vFgyt8QwVYW8rhPNbx8yDWlcHxHVM+f68d98SmqHlIdBq
liJsG1mfFxri0WY0zfqFpCa4nAUI9ikerbWSuHAcq5OWBIAFUL0FlI1Tz+6UnWs1
RCpoSVobQQt2HbZNezohTGN0EdciDNuKZVhy1/QtB7Pqla/nThBlzlWSTkAYiwPL
s61mGG2FDzUvdlkV7Qv00k5ZkegDpgKl+ADJCwhqJDPSBwA73uanOSb6idcKIMe4
pd5zQ6QOhXVLmz3ovBxrhsgjUnKDnIIx9ljP3EZ6rSeZtmJXsdcW1P91vp5YkQgy
3Aqn/ZkFQcoilhny1soAssViH5PeCWVIuT8zBj6rFeDJX7txGemmUFHD0xr+npcM
`pragma protect end_protected
