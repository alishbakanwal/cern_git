// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:02:10 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Kkh4dfHsXDK09VuuQ9Thp5WaGZvZbC6OicgrN4JW+cjFK28rrGWOyY8DZ19+MJ6d
9t95S9PQoPvRYhgNmpNWXNapreGZmUnTZ+mSI6OPgZFRqogx6UNr/9PGSvTga9HB
OvNmGD/EJzbUhpczqlfW4VlFjfcn/MnQzgw7lAwKMLo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 28224)
DQswYnnr5Db7Vnv6BVvMwAIDlCMQxk1uFpFydAKdNXVxXNttaWY5zUzfAW2pPPDk
PGehZPm/qQap4AduvVKmWYJFrX2E8UtMrON4HKEObTeR8hfXOdpiwffOxiaoosR8
TSd45HgNE/knaPNWcvGKhYow+p4t6RDZGsgNz1y9TVL2n64ETagPd9X+RqKfclQ/
BbXJwSdrhxuxnMx+Nh19DRpRQyeLiQIQihKohzd14pf85kQCTZzHMeRScmkdUQYG
KsTMltIUgeDeqXxBV7JaZPC3XZZkhT4MVir7UmJkb2cw5n38j03uAJ5XLEDhDHHX
h3JzAdJfsjh7e9SqEcbjArmQHFZmvpUvb5ZS5+RrOQIUfKXlBTo0i8eXU9cuWo4q
OmyDQCpPYjU+Ndbt3GUpkGb2V6ZWbkd8VRLL9iwWk0zRKZrB/GtWqp3NW/x6onMK
MuFXv98wmDynKozxdrnYp706gN/PzgCaGnKiaBvxgrq6iyhKIb/AQCLidj3cgRnM
y2h09g5LwNPTJfD78t0pMDQAjnX+SxvDEOJFfuYGELPyv7tur06spunKmmYTyMYt
VHq1dMKPYeaz3M5m4eIivbmMTrA3UrENwTgKMRbdvi8rCQ8lrbwj81a+OJ59hkbS
/5l5LBsaDsVGRFTBM5Yl/H6ceKOBprop1qbKzt3ZPpnFoYPakeKIlY8RTpmmUGCr
tbmJjvdpqXLyBzdU+w0g6BfBxbxMwKk/W2CO8e6zzfe0Ra/6iwtLSRTKvvlevrNC
ARk5IjzizYJ1/eMRpnXe47eYPPHxSRP7C9y7MFmOAu/yyrIcj9VQbEbHEDo/AHEI
VI7h6TOSpFsdwtpnsDH11KDAnjN+dU+RRDpH9HNoldGiVQUwR2rrBhrLn0HmKTVB
2m58oW9LWjrdz633arrU961TqoXU7mQKmjqi/+ruaMWy+BncaJ4m6tkv1rZv0Kew
ybJ4b6Rqpt04fR9EnGbXRo0snQ13g5yvVeLABCHVXdcCHVQrwFjMvuSAdN+e16j6
trUWm276D5+hLd3m20B45lDZOUS5gD/wHDpCcbLZsW3Uy0llEyQJD3cfT2rAQEll
D25zzw0fTFyG5TE2TUIayi2TnIJotuL54we331LjDudTS7SMLpv8+w6KCMduUJXy
RLkQAaMVq+5XvwY+ELEwu2/cpeq0qO4aEMP/e/UJKNm0ix2FsH9aBbwDvWTpz294
+DWSRCzMSPxzeJ1vazfLRoxxWnzF18X4BO4ZSGFEe2rHikI9JgUiirviZBNmU2Aj
Wo5YImYd3SiupfnjneHMst9sIF1vqDCO32xTy3J45TBFzHi9iNjg5/B/kzdYxLRg
8dBCmNsV0wCEr7bnmvbbEf6xnRdH5oC/fLekAYsRdTty2PLynLEaPKGVvQMufiKj
mq0aveZuXMdkjB6PSkhsmHUGBY3AnoN8sKT5YTMb62J5gBicV/8CZVOhCvi8tbeS
pXQ0kLZD07egrcdlG5iNfD+XS7vNQpft/Z3TmwgVZslC30uzNgASM/7mTB4yr5as
UzZ9979r3cLOtHeM3F+Q5DnJLJ872sOJgj2Uen1yOIe1Fjf/LNEZLb845aAqYeEd
FGvTzGpGB2AlBRfKfc2UuW+oIo7zXp86YDjg/9xjZb1BabFI2LrXwPa7Tc6znkeg
bMDeV6spUFWu0CX+WwDzsXp63ceB6SRle4E46JfainFPseImAHRg4FS9QCp7RmDm
vE1lWFuP9gsuGZ9H3hQASV9gd0XwkADy64YI5os34OrZKxKXLfLJi46Cz//yg02y
NJO5a3+R2FnBlnFuenP0K0QkpgBrApi9V9gOacfiOUuuCsrpbyePSBPzbHJ1FTCD
zCGRZXUg1akW/PABVGKK4OFXjsZ+fGt5DCr/y8mBQyFk+fYKMQKHD3tqwPaJi8rC
NDpfgvRnF8wjiYLDNXkD97bmpxYHTjnPz7fkULVgcwBypiETXPAau7G1JIJKd3cG
lr80jQC/mJoqtOt/LVmOOgT+PhdW158HQlYzuBOEUQ2zvxnrmsLDXenwo0ccoO3b
q4h9Us+x97m5fjEqkljU5KjhuwGRk4uFwJa4EiyGOImfWDQO+6Gtgn4FpjCvi5kT
qdgPWKPm50qI5DQWCc2Oy0XjjZiwqAHohkrgc1MDMd8BAEXNSQuSY4ILvzdPO90U
vYl8buRPuUiY/L+4fyoHJKkRrv3UJgKDXYtXlPJYiISq1z0ft9bSWz2mTm2cOWRx
rS8cTGpK693MLc/ROA5fjurOqemzxy76AVv+oAVy5BkgbhLYK6yRgBZPzAjUGztz
2b6iYOD9yI0sFiDdGaSBTb8QpU91dLLO0H5omNcSm4XcAYKl8brOYwfiYrJaoM3a
JThCX3mEwO1hdcE5ZJ9l1pETyTP2Y2BzMnvXKz2s+CBeiOfZ6a5XnPJbjaMc9UhD
EWGNtm/709LKoAa66ovmPUqYBDdMnDI6r3NIE+S0fhPjpBdQDsALwm7CNpnQu8lx
zExZJ8pP2vHssnmyA4YrcTUfnuCMK6CE7G5ozFMvZUnrgXeYK9QaECRlqVAuijO8
1PoC2ocIoxSUPaiPD/XB1g0D72Pr3GUIXyEtNh7pTJ0GGFH3r4QkVW+Xi6OI7YfZ
nTUux8yAHycSMabYGSXWCgn+bkKZ/30Qfj3JPvFFYRaE1ppidTv6EWX9YScIKkF3
DW47mKMhgpFy10I5SVpI8KXpyk+WDOMh4xhujvmg+vnY4dkCzfviZb/ciiQWVqfs
GzRmS96HVpmz4UoBlNX5f/IzZJvKkqoTTTNUWmux1iR4QzIa7d8gFSlSzcqgECMR
0ckRpPYGoPcssXDApdpw/16eD+IliSwPk4bSVyPtrShbiFmfl1tnl6qIxSj6WEaM
7hLFdfurxtcv2onGy9eY4gVYdhKa/bLINLojX1JAFaBwQ4VFSvu9Pnc6dxJFHPrC
TijkX3LrWjVHpWXQyEu7ei8Y9XtjtADjFpd3AJgzJN8zeJCA1omDqwxJiuzpeQ0Z
hfBa5bbnApDypbvyouGiKp1d39z3LLohdDessg/v5Y5qAEg57pmuNIex076xjOqJ
hdEUteg0yRbHPIK1VNLe74YE0JUVeRmPMZ8mUAigXw7aeAnbwZNW4C1C75XwGvO5
adFESf48PGWCfX2Vdxog+ofXxoeWuZFzamcGampcuA1BLA6r27UQD5ApQ9KNOKJ6
uZRWqzQwHVIs8JOICCqIRRwZmBTNTS/Qr6/9hzN0e33KMH8BL/wO6uH2dVhoFMf1
ZcJKLfhLpr3KQ1I8i9mYNCcLgQH2uogTyg+KErTf3jol6MHmB1SSrPm0w7l9ve1B
zvK9AC3+FIEBi99WNBDuqDqwhJvqD9bTw+9qVVJbkppydL8xc0TvGVCM/dYYEFx6
FYGbsdpFwuUl1TeMl3GQTiCcy9dra3nH7+bqbW6Y6XCcFLym12wLjo/75Kazx988
Ys4IId8KSrQ59IUxCQY2dHLiOAc9+B19+yTMNf8y9CEkpSq/4LMyq9vMH/uz9grR
+pGhf0pjIXqzzR6xKYcYDAN7JbwtaDHxntkMrHDTCCD/PNLcmNx7FdMfrQUl8KIs
IYJ4XgHQ2L0+gD78gjHjSxmZh+sbNr/ca+REfXs4YpiAKwovwSlxvRvvf1IiSaBG
UCz6f4TjgqbKEy6/DAhPfSxE2ja1Q7iB8ZBTbXEoNfQ3cWFywz8/Wx+Pwn2PFaA2
hKhG5JSf2w42Iw5UkhJ9oYpSRzVOBxfRuipBLrVcGwF9XddjhG5ydUriwWB7qMuJ
2j2ZKESngCB04TcyMOB6quHhw3G6ZQDMyfQ1Vgr1TMhG8Pb06MfCrzrv7LDNkPNX
ggHhrZB3S196kWixgDcae8t+2Y0QpTtH85qHrPGDtplHp2y0jR2oXCfD+rhWv2VX
kMqQO3lwpARgMGIrLxBj3t5Zxowy77tP9Fb0u8X4c97RMsh+JnATSlYggkKWMw71
lm2vll9egWwIFXlUKoqsxdgIB0wI+OgOiVNA6mUDrT90RL1dbqZPByqeiSYF8/Zt
F7Yg6jXTsgTS9+0wrecs7nxVepz++4C6/NsqLvz+3QKSNhF2IH7xyZW0ZID6c2WI
ZYchtcu0U/qnQaxzd+BcdPLADAX0FYofT1ZGJX3fpfBhQsPx+aeH52We+XmCF1IL
A+L3TeIWkNXvZEp1AKtrb0+5lSQfHpr4wtUNphBNcZUPyHUOzM5s35oim9+yj2b9
OIUFZ5fw4werrTfAa3VXTyBReLrqQtBneio3+anDDJRfMSgJfuenfHyoB0mbxR4V
zZHv39XyCMyJ+TYk53FtUyUBGM9r/l2YkkAciCSNR2//xSNVTM+rFhMKR/mzmPyn
eOK1+7IUfOWk/vQJoB8E8UL08YC/rdqG4MklluMV6xYehpM43Uos/COPaOWXwUzU
MOrjESASvxIbaEO/mV83vJ8CH0vexLebTCmc4gC9ktmPYzzyqHAFu4nHiV2PG9ZF
V+LDzZOLQB9R0JMyZaEzbF3h2WeL2/uLaCwuAzdZ6y+za2/SX3m7WARseK/Eqxhk
vHvgEFefATxiDhe7Ppo5SIpi/zWAqvGWjFUTfUL6yNYO6Hwj4301RJ6HKvvpbKh7
Y/GkdvjWj76hZVHjsx4JTjrekoMRmSR6qDlzDZ5Ppl1K/4WMcAYLPTaNWU0u4fct
F7xoLkB03qsKiTYG0Nj++Ym44I89bSNP/5ItEgYbnzBP4beDJeev9mr3raWxdZXQ
N0ZSGQxfNNDFCWqrO/whzqfCLuvXSFjbhn+T2NAVZTtudWzyey8jT2921DYNrzFr
TXu6Yph28pcA0MQszAY7IXTjie6q1jmKCWzFlW5UHulTWagpP0GclBDWOk+yUQX8
yYUH4i4Chiq89diVts5lSVg0aJ31w1EGCvMQsnikauxt0N6dGOLPvxAXBZsUPR/s
UTu//QnWYOvlM/BVpnlkOFZ55I7Ny2Xcynx8tdCAoXd5avfcM95BuKvCm2HZNvfE
Eg9RW5vjhpSrVJZeXEvC9YrPTnzJ70yTh2KipZ/A+0ambzmmDCpzwAQAgfW/+sPf
bwejHd9yB2cx/YSQIaqxrQvJ8msDUFpZf4A7w529LNrAOLn+TxTm4VPVE0HwwCo1
Osp/l7/ofC9mE52Qsm4o4cya6RukdrAeEwfeeLZpAVEfPARbhjNjPvOdO+CNbLZJ
nmuPm2K82ZGQS+pFM2aThyCwYAH87MDqx6BDro8levMM0Uie90hp5phXa9BrkQe5
E7peiBvOKuSP0rybXmnDRtRIYUhcoXN3Taajj3AX3je/IyOKGOh+2PSNdQgP6tgn
mLF/2xaOy1Po4P5DNu3gJYd/7J6mAUSripCtuwP7kCburnRrCxasuTkH6/IkM1KL
63ACX+gN6SQv+w0q5TMrObhV0d4rHF1kG7/L4mb9oylwplhpp5QepooN2OWP9Prr
40NOZvJzj66sixKvuE68eIuWTTKEO+FweKw5oHQ9Zt5KL9FmKGslcxmMmjKg+zdg
RqbDDsKmjWJZs0Gf27yNzZ8V9UMQtuZ+b7+rqddiBY9BVWetb0cRtqcLY/6vebsQ
meZzTYsFhxt8tjRZC6pfM2la+4ONzretJopKMvQoGF0CYs58GFKBZnmNaxILlQA4
AD+03VQxFHt7lMozrHNGi8UnCWmZ68OhMQcXvdY/3TtrVcDM2N+IDJMw4p0dPRoz
ahnfoPNwt/62BGu1yyRAMnAuhRKCn2eg7tGTrDAkmEFfRRh0s0n0Qh7zmbZlSo9Q
0y57KxH27V3qcA8b0ArOdHnXsudhVu40BHk0HdwFPSi/AyCRSP79IVKAWwU/cJ8q
Xu+81rfu6PC3Sf+f+xLi0yTQaV/ViDAofnsk42MtrCUV237qSfgAg9pm9VBYqu8B
x9c0LGf5wbxacoxfyvaPtOflE83JDyeIoxeBUR5uBndC3b3Vgm6Cbwerf426YNbR
30g99jCx3kXSDjES7q/sxLFMWd6kAdM/vZRDBes7nske9sHWBoLQh/s9m/D1YYu8
UD4xPLKilOXWLIDUN9S9lJjJ5PnJKP4Xl29OfhTfW+VHJQqAa4SrFd2qsID6UFGU
OSyXRQdTkQAvV/I/IovR2SsH+Pccu8c4dBvz3UZ/u4yEZ51Q0T7TNYrqVosCQjX2
EpQWlkZ/RrWrTPEfRubTFM5Yyj0KHyroRgd6aU5NTxiFRfZSeLVEaHumMsaomHF1
rMjZkdYb6rs6hDkVpq0JlfVyrb0jCYQYeZh3umYHnSDNQWGOvIsVYJpYtwxYqjpv
LBe806eIeyD0zBH8PrBM+fD8xRaFQOInOa6Swg1RadwKo5oVZ8HnA95MgrVVJDTh
pdgmKsgQyTZwSbKahpwfSBY22DGZUvKcnuXefAUuAiyg7zESpsLOT2iPk9CZgb0N
GP/wU97SKydds4Ea1v7zYCUXhMxLuDc47vvGrsO7q0d/cGCB7j/px7nHt0as1zF1
6jTv2//QAN7nBR6FBH9g1SYg1ihnF7e6b4jQm9zJZ8bivwyqGsJAu5PqffWaVTLi
2YdL6D1Z/LstTueVZ4SIQLJ85UMZD4yxWFqxVoknUceYrUlqR5fPEJwPbGpy5ZO4
K4twl1NBW++ryLrBIZUiJPKqxEZKKK660q+RccVfJRUrmD54uOVzyfuPFbEN951k
vMIroKyUYCiXg1HOMNydNCZvDjkO7vej66EP0Z6hw5uPm6maLcesQz9WPkpi5mWx
kNW0LeUH34I5ehdc6dIOzefK1uJFYvTd39IYuhsGOZp/uEapmaKiC1gjlor//quO
rgEhurnEacnE2wUkMK1AYxqA+fVZzv9CQ6MqTqfiw9xPyf6FcP9EKNXk713+QilT
AfBUbHJzoz+4M/oe9AW6TU5YMjx6Wc9OTGD5VPJVO2UCJQyM4Xs9UXbzGmqpXVde
T68lOTn8CSLHWkx/kHaDbecq5zNhz+WqKlE65UztrpuW2mFou9o4PqMfjzPO2H05
UyJu9Ro3kyuxZCSvFmfaEhYV2BgVgjYyBqSv0TKcMksLEd6LMHFIcClqFVpdtTm1
0gTkJ+og0whpzLBJhqdFwbT+xo/irFC1AeUmdyvILUaS2hYM9YaQQBGN+MxKzEzJ
fRuQ+AdDvU1h4k+aDOr97fJ3WGIaS+hc8EDNkoinS/AEh9SVU1WWB/jUwjpWENMo
JEo2cqpFz4kruWao+eslMN0EKxZmnTqGZJP1bmyR3VgaKLYuvjTydYZPMU9ssDx1
AayTVVi52sCkZoJDomxC6Of2O3k3Q95kLDhXjq8+O5pEp23N5seOHGo5rz23KSMg
ehPlOJMU2E63PZKdulzFy9wQm47p8aGHcJ9rIQsdFY7/ObhpMO9Vk8iLNawHsuvE
dEtjDYVVKYvfyOpZl2uIphNVhegexrQ+G+IjL81x6ROvA+H4ZnkKzOVaaK+3gFiC
diT5TADKryqlFdQdI/J+4a+SJ4h7is0lZL7DhesAc/ou1jIpWffhwsarNE/Z7OrO
uUjcPRYaoF0+yZqAMZaDZyiBy/83TUCP0XGz0v44tcieC/JPz6DMyUD5fsJZQxlf
BnK03pOcWiCzgzbeQHS6RvBLerrXkwnG5fVExEFI/XZ/nLiM6bCVQfxS3lIpu7xm
i0+VOKaT8yULz+lAMvMhatm6VndWGZuX6bupybyGTL/LuVs1Q4882t+M105qBetk
6l6yyE/XQgOq4vydsAX7I0e2houT8dsN18etoOlB90yaBg3BCGKDv1zPa3aCnyM0
6flNesBDvV1LPXwQtJ7KZ2AKLBuRcg15gAVVWhQBz9pPVRRIfh7AqpYfY+vQfL3K
XUYVbm1+qSz6uz+UJlbT5D3rEKdi2hX34Tha5bWF65fSNBh6YLkjx/7YSl87ggsr
bCxeeMWp3TXZ7J78MNF0Yji8Yys6O3ZfttR7aDv7w5/XmW+GFFIOoKOpFZL4b5lD
VFsNBrvHvDquXkblTW/i33TZy6xhoEosjB70ulvpr97OtmPifzyuYCzpr5++iRmg
if9DHRCYQzvJkOb39wi4rokxocfhwW3k/OR0jAq231yR0ev1DOQpHPq5zl5ib0kq
y2Fqjj8u4NPtO5vKuODnXNcHiFPzJ/nSpMqfRMy3TsX9UszcomtxWaKFoKTcX2aC
w+9u4BfqbIMGRdrch3gsI+QoSBwlVbXAsh1aN3zH4lISRfkkfUQu6J8w4F5rqK2E
WBusXR6o/R9K1OvMz+pHNVgsCX04Aw2rEtTSjj6cLOJDTeS8doojQNcZ5H/It0ie
uidm3DSTrrpjP/v+0YSqSkXPa55zcS8CRRUn4sLP9h8WXObPSnPZGyB517PPZreR
GMRcIg25JZeX1T4n/1dYsgdzXPUcNnHC6VbIJTw0kQe1teEefNqUXiSG9kKY6n4R
SBZJ47xA0NNrnk4PldrArCdt7qf3JP8Dvzyu/kUzPNF6uSKLSxpejcX/KNMRNkOH
F9mXlysbSlRvfwF6bcn7y4Elph1r2pD4DJt1g9fJcNRBT0bagniOePVDKqj4+Tm/
3QpeWNe9UZ/UvGGEpp4IRMhvqVRYkaNuxT84ktH+nyx6uNqHXXoIuGSH3uIYlGHp
R+jSLiZb4JyQmM1nJdyns3DtV8019OJKdiJN2E8qj1O26LXHffEVvSLLZRaRIXQh
ednZyUGp8lVbyg0qq5ZN6y9sH7Vj7JNT9velpD74PN5WjlG0Fwg4+iXnupYRwfRZ
7eBx+j1UTThy9TAAivwiagOGzlQ3vu4K8+ap2MzWCDIauHInz98b1T0FxUtMSkoD
I8v+niFzD2Q3es7CAQ8GrrcKqzK9j0yBx9jIkR+lat82oLXnFJDS6wkvSikKNdnJ
AoLGABN631vOP34ahnqzAin753ZDLq1yF2Te1OlgAxiWxDMgmmTJmuYynwKKZUje
fuchR8xJW6Fn57hlA7c9/ns7fS+h5Okhy83dJvm5WQ2cDNxCvorfTsI+UzmjWCRs
sRAsTCGSFfHvzhKzBDHYlf3zxqrbDQnrzKace6XTIffat8z9lQgSO/HHwSjcYk0s
Ow4/AY+QnNali43mNW2HETLYVJfEVgs4kMiMWHkXlkaXSl4IxjMuDBrOVo3wOYK9
Q2V4ArnFXfrccgBTUV36ws0L+Vrr6rPnkosJg7OuasbrfLPOZ2jtqjdcYakIKrKp
8uuuxctOJorMRpifcNL3pjkNvA+MqXSdXPHT7X+Jnr7P5fQimpM2Fo6vhkYAi96H
dG+3rKXTbQRmOPxXLcvYaJBHTAD+O0qVZuSKKxLShLb/g1pltdLMtqCvHr0/lPJ1
bvjKKXEPU+1GPDLxJCrRYXrqBr5+W/v1ZBLKDOg9rH7sOuAAGrpvk/BlW+vApj5R
8VWXogNKeMFZ65oqOBB8IuHxC0VYLyH0SiOyh2gMnxwO3e6C2nV01uC06p5uNCyG
dNKI/3DeyyploFV7o8p8GOlJk7Nf5S9Dnpo5bG9nNiKylQwkJsY4jaxaPcGLHWlZ
xKztoEoB824W8YuwqWHZoc0OX7jmun8tYP/fn/ShEnlu2EAWc8v+t77nqWIHOQES
xl7KdLmjPgx5dEBjcyY5RDc9Ry6L64HPxbS2GojYyJIQjPIteF8VBSN4JImFlolP
b1ftHfYeAjrCkdFiXGV1sMu/GTBI29tqWW6r37R1Ef1PWwwKH9aQShnn7lR/G+WZ
VF5wxrHKqJ7CU++vwVMar/XCxIJKvjGYIR8BieUn2eXOSOZyfT5uO+QzmxfsiF6W
k0l1sL65Oup5rxTffX6xb8tehMKWrL9l8j1Du+QWOWNM4WlbsuZucdPZK8U6KjwU
CbRW4Ns9xxueDtXtZr+mAaCRs17LYMRUYUJfMnFiGZLYopi+ergZZ+mZ1yhlO4hj
VWbcsyp1vVm6s+7OD0Q+rAWtV4i4SPsxo8GFu2Hdg+ywoBZw27r+QTyBFTRHTM5B
RCFNU4nTc86nhxBvp232hO7hYvmp6dlLK7Jh/R7xoegcYeT1UedbHh/UVaZjhol1
ySkfxIZy2A7EVyIktpjKydB0bfZOG7rMqw8Fibx8b4a1WS6/xgu7WmjALKoI4Ia+
PxazsurOsFqNj7MbH0/gvvHpRwVxgZ4FRBSeId0vIe5gpsN6S2Zj6ddS472llqIr
6i3aXQ7xOjpcrkqeSHIq7Le5s2JXyaK8BnilpNiCtw2hUJAnm3UFMLb/kRYfFbkW
gMl7HMD8UXe4DRQBH7C72wWCugMuxMtSuNBmJf8WlffM7X4RlO4PD1OHIPWj3hYX
upea2l5jfThHoJQoMM0VIZhPovWCntucYuQ+YPY9QaDIRTwB7Mf08RIzuRxRkvSX
KFGEugkAC24h7UyyoENkplS4FHY1+JKdRCrKeRLkMvWvOD89j0P2XVRUM67ASr+x
wwMI82Y9Dafoa/pzPnM5VdE93wEbLzZmzPisoAFuZjpx4H3EKGqfEci5Xx6jJPc7
IJbekbUie7DHy1/RYQu4YXqUo2+i1QQW0gNi4BR3fcZbam6AMJ/RrqoxgCSDwlhR
1/x5jdFQD3Kk7OrQmjyZqOSbzq9nUGtLS/EbTCR9WW+J/nepG3QhavEfIBxLz8sy
b50MUjMFLwyFW6vH30Hf+wh1TV00/DeeqyG5VbJrK8FsCuZrZX7ylYZqK/bh1/Zu
8ZQxMylaxGO/dMAVxt1lS3bFLflFZg8B4jX9rJskugWUnoXQP89U+MjByrTArl8y
MCSStKDjyWN1MbEsGwes9TNBOx/bdX1IzxtgtaOWkksBw8QSc8QUq8DEET/jIAi1
GycAZX/TJuFFSWAwD+lFZ0wDfBIfoppD8L7ZKiv3rt8H4zF1jDi/a8duKmqPpA5E
aKAlPlgSz0D+4h7COF4ObU74zMGLKKu5lDfvxc4K8RUD29fskpvHfyD2HlyxKj0R
D0XWOQsXh4x10m5X+Zc5YpbgljimDGS8i35i03qWrKLTSehvyW+Ot5LLchq4GLmd
dEd90vli8jxEX5aXBEDicdmAbUjfGJGC752lI/YvlkEVwbXFFuyOrTZ/AeLFroPr
dOLTMUk7T/Ce+nhjaHPLDwAhiwLh/QxIFSpDatlfnlc5P3k5PZ0igvNkFqsU2HoB
KbDBsqCNoFNUisbq8TWphQfoWGS/a7OAfw5UTIDciE/jN+cplMspwyzWPEcf2h3N
8gb9FUCsMTnOtKIvirQqHGY+WWd5dx8qYwH4DAR6xZOf/fpDsb3J6hz3BcxKoc53
eajJiI1f7OAMBdA4ZzFyybzXWkSiqvAjYZYXaE/ZXAESVISZEiF5WGlTb7FqQrKL
F3ccJpxUndDziIfxEOun6LNSipM04pDR+/aJXVqyvOAvnGnP6UjuIvzL7KSbKp2r
Kel/3QO5GRDwTQDHIiYP/lI8uQ4M4kriMDmxVMthsBN6qvq2iV9y2ziOhynkSghn
zPr0SKMJ265YmkMP4Z9Gs8QFpwj02mlrSXKDpXyfZIRuTirfcr3/g1tGrfzh310I
MhqVAxuDNxDBcvdjIquird91Vu8NqLLAoc0RY6MhS7nfVqKWtwZZkyn8lBHB/gSL
35eZW16S8BQR5Z/kk3Cm7FHcUfIWScILwVUmIgHER1k+ioHXDWWiTMtr+NeOKHGv
Ynrqk/zkvg4H1Jd6PaiLYNLG4dXJDDUMv5nwt0sCqCTk6g401zNrKRuuW6i1Lw6C
tTypkEGCUl57IyuHjmhPqXcjnlGlR7mtNklyFa8FJ761xsP666iosfP68MMsTEPK
EqCS1BL+Lfdo5pqcPK0J4fVkjShVyzRggkQjG9rNusbPs8lEVs4PeHGAPBVyCtMh
cf7xKviUr0tIXJivvpwlI7nczFnVP//fw4y5FuvHaJvy7lOXN1rcS14yAJWNAM/w
qzS8m7QzqB9zlyijT9h9gYs3TuY98FwJHKbY5atUdp2F7PWFG6zG/RIRDvcWUiNd
U0kHj/qBxniBovsSC9fgp7ZF6Ifsw29OkR5rxhiM2yrOv5yesE70kqOHfBMhqX6v
NnWotD4TEEli6dfscdgvNLzPwXPAjnHryeE8WXItwpgxQctMHHANbDijsQV9umsE
hGTm57gpAGc/K3mY+bfldppYLbPwHwglXbo3jNgdXOIZk/lam2L4TRJ5J7lF/fnM
wus3jY2CxGnXAQPSlPjMoctBmxihMlAeG9tdH945hOImW5eFlMBEI10VhxwLaV23
Ji+25NJ1r68hjmbQJRMMxCh48QNXXTQM2Cr9zN1cxWqlHNnEB7Fkliyu1vmLWxKh
AlIxciUAih6pnkJjC2HSq8UhxqgkJrCR2kabR2He8wMqweE+dfWcH4E2hjXMWRfu
vsP0Uu3JF+WfbMmR9L1e59J94eSotgdI6RaFnw7n2je+wVTMKgarC/jM9YS6E2Jc
MEuJ+bTUT1RO9sRWAHIGSjAhd69IXPhGoCsbYnTaBIHM7PLUSYEDYz6Iyg4ZzGyJ
BhG71RoUZok+D/F4LU/WsuQO3GR2r/O4t57Ax8Ym+vFY1vOE8OZU7Nkjb94+FmOH
41P68z8Q7y3sBSmPnAWQHcPP4EfytVsCrm4PFi5avf108Bv3iAGMjKCiQZP7afuy
LpxXqSAgVS4yM2aVxm7JATYiNKL7hROD74V8n+oKsDltPdIrO4vp3wY3N7wd+om1
doNsMmUURH5D0idDXTrZiMRPjaH9F1UZTVAcO0BsNMP85tjJUoI6x47ZGDXMRGKs
vLbwcvo78jf5bmdNlRn6PHOXjFS4tDeA7z4E2WStzn1nYjxjpmPt0Ur2dtOrfQqY
4FomCIPjDCsufseETPfY+axAOczFpcoNPDTDUPiZhuvYag8ByP91rCuVfBwLj8TD
HEvWwqEZi4erDroZQ+Y7l/uSkZ0ACSUsQRgxtIuCjWPSqMSKZlN7u6VflqMVO8kP
RJCRvYon7FAiEAmbHFHGseUYPxTLMd+g2ZgEtze76gNFc8PwYue5HY8rMd5PoVYR
iv9AxXk6Gc6Sz5hIJDNlt57A0eDRtjt7Q52SYNYwmmX1jvSwRSCP8Ivj84yzZsRL
cZxuPsRTy6wd03ddKUzlE7WWwecYdqVIZ0w1hibvkPUOVtxDNbmiyi06oVWQKx80
1+evsOpqpKH5T4g31qpEIwyNt3XCSZnug1j6HXL+5XUr6IODLKOglB71ohWOHI6p
zN0xMc1UBv9vAeWZo+rSWBWATqC7TYG/aBLPsaXMYt7ywP6EhYAGrUQK0lb1oHQ/
EU8wuVrFwEvadCrS+tSoR7fsa/AOOVukjv0sQzDT8eUDU69DQQE3FwzOGt3MCMBi
ryZYz8DTohrjcBNK0lSgOOWnv5mtxUfIe1sJbz1zw05WgH7ouC/b7FDRKeqJZSpx
aX+bns9E0moqeXVL8fWdFymL9oJyq/9FExHIM05g46qlj65RVQQVLew7e8Yl33/K
mvwl6N4yeY3Au0Qmh6YzYjsaqTaaNKA2AgO8klMluXtV8D2WOnaBpLqgtTGOT9TV
zwXqOgg5BVreYyiw+zDc0XJO3KGKmAuGRkse+Jt4CJEunwx/8JSBJAWPKJe4rHub
F6KBftXNKydq+VkWTiPX9DNVKdSLbMhaAQnXDSv11GVoXP/jvhAZB+O272aqzguy
+B0M6O/u5VxeXL8VtQqyTaK5+tS/Q3opThiswdIGde9eLAE/LEd6YQnAerRpflr3
FYM9L+geLJrz6JpnRM434KCFEuG7ZbwNcmloUx9vpF0MIwOO+jdZCCXfF0r4c4K6
PXBFqA2seU5QFihCImRZukNW2U9amYZGdEqayn0fX4Zp9H79xBEwohGAwuadrFmB
o5z011p+ng85mp5zlSMCPMuyCPFyfoRc7/68qws4RWDXRs2SWW2I8w7RrZMxBHXV
KcAfAI7uDTBO2CCtiF5tsIXKIqBPtPLSNEL3JM9sc1xCko8ikPXc7dy9u+PjsC4S
1kQoGg+lD83bmyfhvdv9pJZ/0BIh9QAGOvHBYVjKMjSYPRSnAyybVYlinHbpxgRn
WnmKBRXiBdpUdX1/0WPwQr4qqLG4Rq2phauvuKgAC5KXSylCBUD8UyoBAgyCBjPs
7SVPr9kWTlUl7qk32h7zAVOLG/rhNgubkxT7b4tXUnJYLvib/c+scVTgsnq2iUr1
WuOJ6QTcn6lYCkEqWOn4dp0e0y/w0Ki9MQHyt4W/NjwLbCvYIxtLtjKlatF5CIzd
CR5S3c3xrOem3D/VnWf3jEvmv+BwON3NlmA97rOQh26w/tH+/u95boavsDcYvR69
san5oDkRyyZQ8fHqu9g7Ui3+oLSfXNTx4ifQzx2Z1w+ySpenbnnRzJAPDvPKzndM
NnQFW0L/uLIotK5oTv+oZxcvKtpx4vELeeqTy1i26+EwZ+32zVszdPXq21q1PtmZ
DhywpUT7h+rKWucjrMb1vlrI/B0UU+TDdU6v9u9e0FhzO3hsf+ZOPwZpAtpcemOd
6cVP1YStk7+4gmZtYIyy0n3t0hLEp4BuOmGvVx0DgCcwst2krqfriA9sPQTMPLDh
SapIWpEaW2muO92owkq3Whawj1OJ7maII6iKlx2Z3QhTmQNzZUz8npGfWjRShfeI
b62Xmoqa35+3LKSQlnDYZBTiEo5VTEjUzmWHvyCSZjYJ4Js9Iaj64z4Od3BLWsqk
OxQtYJvB6ddIKSAdhpAJnXQbtvakWWxC6yxDgIOn7y0UoDN39If/dIVLyjC08JJm
46XJyj4ODpE0iNSWSwbgiLRrDeGuV91wFZws5soG8Y1CzJeZgkt6/qO8bjO/qyHB
72HOJK6JeIqR72/OK8gyeHYPpWCkRfX+aqD22k0HOIgsOwZQcslLfZK48uwp7pvs
5KxU1pHIPZrL+r8jPd5L1K3HxITbYajgyiZprqQ+Fv4IiX6fYT/E5YpKw66w2n7V
pQzlZHlO5MfPO/wtA0JoVcOTjU2j7iE6saeCTgMPB583hv82UoW1ObgW3d+GH/AC
VMr5vqAZgMl2pu5A3718Gz2eG6Kc0fwvoJ1l4pa+FeIYTY3j5nM6iyntFrO4dI/P
nwUnD2h0FK1Ob2GEKYdfVIjpDJOu7cEYDqVqfZdBapkPgz2Af4aBDOhr1z7Vz3Fb
xI3PC9n+BoGhlEzJqqRsSqKz0AyyApR+gHx1vz7kFdYuc6KozKzZ1m/UstQ5syta
4RosfDc0AefrunSIcrFleIHRRn0nuUj4Ah87o+nS0fEwgmAuPQHGw4/BOBLfCM73
9SP0jkF4W0WfXIGZQi8gTMjLaRnn62XM0lV1A9+R3UEjpwKxnAAIjI3jJh3sVAiR
ImMzbyhvu5Xp5WipM9W4t0U29shZCqHUepPQLPXCvgdY/vOf7zw6p1M0T3I22nkf
R7QpNmgNqqC6d7s9HsejOHoaseeCeXZq3wjiuknTVyUS2cXoIr1qkxEFCNGnb7/C
UnswjtVsO2/+newVdpTiIfr/T7yilLM+sdtrAkfops5YWZa8tQeK420hYUFdB86u
CVaGLHD544nW7KQ+HHKdhUysWkm2LxYjVVIU7+GaXiYa3zqVRyJlEg7Mt2L2TJjE
pSAwy7nyU+sabR+cw1RpQpMuNTR8KtbNKFldSvNnCVkgl366jTDwb6OMCzaUg/WV
DBPv2ZOWGPnjl+5U7ovbrle7AiNX18l5eAsP0Q1qyJOc/kRAUzreO8pbsuFD71Dk
eJw8WIvp+1wrBafHozV/TnahavWTLEi3luBCu6BaIwj9aINd0CbmkT3C/T15+qYH
7hlMzyrTofd5zGq0IRp5sojTsthmXe3yASTcah9pXANQaB6vkOWIEAZhjMPStjTl
eY0WD40a3Jp2gAAJhrxjcn2Yoe1etySt7s5b+grwSsM9VfSswtawG/aSYG2sn0YB
XO5ZqIp54PHK/yDnuUJDGsw4SgDSO20ARSgg2joklBl01m4gv7CIgltao5BPj52B
e6KSZBEPyLLM+d0EEn00LQz73pExDSSflrAtUe0dd262T9ZG7teUdMQpuUxey0Bk
Y39Jxx+Fxm+U2CBn0bkV702Q9KUIN5HYGIhuwephKANYeuvEXTueQwGEdPScHJc8
qXPzn2vmSXmCyHChtrG6ueox+kLmjrdZcfQy/Zw5UtOF7MPqlLhzT06yC8Q2ALWZ
J8b6GRENxcIpwohgptEvsWz5xUbYGypChWjRUxHB0dAlWsfxCuZXFg/uy3udA4ZD
hrFxKFEf6VvAjKluo+MzPUM+JW50oEtNJiK63rL81TeJrJP16YrOPnmKb1da8UYN
WCm8ydPIyVJMfLJZ5zjfAZdO6zDpAUP9t30DGfl+Q7Ag3cZwpWYoIRyX87mdNQ3I
qX31cvk0I0KypEF1f6/rFazSTOQ3j5D8H1Ve2WoyFHRy77yFzzh3/Hyslo/taSa4
1lgH/PThEp9T+Sc9tP+vl0+i1oIt00R4inY5lqpHM18VMzKBfNFNLKTMuntje+Lc
EK3PqsFt/BY9egh69C2Wk0ESV3ph0JDcbd0AJJA2Y3tN7lx7PyCNwFCamyIMFdCI
VEUObG5XYk+QGtJa1RgyPKkxsV9c5EPzIJu28Dumztbarhu543lsrLw/7smFJ7Mt
wbRaj7ajsLa+K1lG75AGgShd/M/6bGXb8QvzfthhV9QLSx7e+UxXoDvaLOX7vzCq
I46W2kkdkC/tHpS+THNKb+eOs7FQghDbjLEpOMVboGh5pNKSw2lWn8jm+VnWK7wJ
6/Foj+Ep4ZtuWL0S2eEUx6hwgS1zo+97Y/j+1MEY6MgAeYOhnphkLoNbD9UA04jx
tukdDTV9jl+1TaaUmN0wMOHGI9819IgwDj65k1pstoZuipa84dcVA26IVuOgqIcn
GIR6WZrgFFzmPMgVpM5B16kO2rdnC9s5+WLLfmuRpkS5LMqiQpEgq0DIRxsNkPcu
2M4qVZRmuZagsSHz7+pcJTdmjhHkwGW6rGsgxiGBwMcbJcOaTjZarCPRtmNupmLu
22diIVH4Apzllg0yvHDNRPhZGByYRIs1y1qwvzySOEhtlQGEfFgT7CqT1y0x69fh
M45fd3UCtHbyTtGWuuQO94eS2+xZkxATNXOpBSd0642cifG6reVVGlTt4hlfTCP7
aECVGEX8c5sbR2K3olkTFurwrncJf42m5GXuYnRBIaY0rasdQFbPeGPVphUs0rvA
DZU1clCzVCzArw4Lj38NRGXqans1M0oSwGrJI0cEyY7hSK06ktW2+0b6na0eDfoD
It8HVuFSaD4I+pMIM6E0OSt6q6ydyuUA+HPsmonkB5b3lV99DZq9Fw1tVSYuku3B
jNKrrwRLgYy90ol9hyvFoG28bffJcdEdeZVLKSKYllpbPgYLKmrhEEAcluiKS+ox
Vzx8EXUmWCghLwE10JRrnrwPsOxH5Ga7L8dPAL6IQ5EwGfimUtENLfXt2LgZvJ/f
QlbU17N8CccqlOUcWxGTW7wbBXhkzgVHGQF7tD5qJNQjIgZeKJhMhXfxW3UeZxYj
0O49OCjRDvFZjNUMtLAdEGUczSNH+6rVLVmMN/xn8Vb7Jc9HxCKb3ya3lv//kM1C
kQz6keH4JtQd1XV6YABRAarbvr8Jt1xDM2p933xKhPlha3j8bb4WygBHsMfK+oEe
aM3ScSg5no3rNUektbtOVTDYrGL3KUDIlU2KWI57uWIwxHNLseBz+d3/bo6xJUgA
zN234KMPQ+m6k4d6wScdOko2bEdayOCPblDIVtUyHw9CynDPEPAc25tnSZ9btwIz
L0lq+9tGgxlH2Hqx5fZnfIsJMyKkYtnSji2P5mofRkgV8uXRC4cwEo3BlRJIIqwR
yPg3FOMOIgxTXofY1wN4su7fvpfTzam86VTL12DSLqlqZVePd9S73bFaSMy+x7RQ
l+cglbsNFljJ67boh/mCh2rCqllDnMBGkx8Hu8BV4bNIqxMVgGbl2g67vigzJeIj
QDPuEIr9Yg+d4dQDSDB83KKQr5V6jseJLlgMYGoxPKl0QT90gSKMYkwyw2ec2yyI
EYQrfQg9xYtVoZfCwvY4cREL3QgaFq3ZtMPkGPCdsSUypsC/MhA1R84dI5A4+Ni8
Nanxo6C5XvR+zrz/Ajvr7kUFz1dJ1XzRzuSvb2HhOoiHoUi7CRNe5UpdtfORoLVE
81kOS5VEsN0HFE8+cP7wQxV3zZJ/gVavvPmjI6gan4J6j1CbXCAa7of/VO9ZqH8a
qxFZ5VnLLGzCGbwl+bTYFe5Jq/70q9CBsWDGHuXJVDlFCN90ahGQKvwFcBKaQN2V
QFw4giAzGlX9vTDeEz9UHvz0SlYy2ukPi7kPI9nPjbQuatwZMDLqC+/xDXaIMPP0
WCknjmJlBA+P9ZyRo89lXhGokBZzTF0b25AyS8PMx+X7/B5Hc8Dy7F7MahJX1PG8
9vYDtcORpPl+rn1bXRgC6pxWgQoAOInGwdtHiC2mBoQlPUyMRQsiaixKMKCPR4IS
nOy23BMgJmcFZuC6PxPSz20gIDXcTabzGdDEWEdlNr23SoZTkC5pPLsD/0ZVy6Dv
xPX7zu//ZVoK/ISg6ocysSiklXXVHQZTwXrvwqZd97eAjGNUVaviBp9CDCM8DqhT
bvcVYNkfCwdq54nNQ7ZXq17EgHaV9EL2LDDgXJAmEucu5mYxR3Z8j4LxJ2HSfaUG
ZlSxaJLcqNDkRpupPLClWvw8wkOlf6RxeiDyEkkolns2pYvJqoKBTYADEfGJEDQi
eJrUekSTbZjLsUoTIf9OEH1+GAQw7aiS2fKAIU+qFH93d1FCH1GtDg2hgFl6+RFy
bu/MWKN+xbe0R5oJwvhApKs90Xg0oHvqXWOh5mrZFuOEQOIIOnVfTUYj9ORuFsYq
MwuA15sM9ycTonN9KeXtpkTCkc6dkOfCwIHTgIdkFEAC48B/eF+2lzwP56Ku17Tv
lAYg9N+r/hlm92AieBZi53X8nRM1kJRRL2AnZ0id5EcfwfNv0gBkTNQaF94HcWNg
f+YUtrSSDOuVg6nXmQF9ehbQaM76KxgcDqh7Zy/w7h183IbtUP7UdwPNg+0oh2HW
2f6D0S3lNYYfcTEyW4Fl07rsFOntyC6HUDLi1D/bmVoKktNk/TV1hqo+RYG3yRit
Oyc78RWMDMcqnJeXIvernxO1FJcwRzGBAiQAI1DB4GTKwRRpBnz53xlcDiT7UfiA
ygrvXdqdXNrxRbrhUTOB9rJa4vdjtK6V/jipBRZgVcf+R07+RNpcMjOh65lcLVND
Nb4NpBxJaiBxrAcODlHIQjsa6eetJpbjO4uzDpgNDUp9auMYj+kUbWe8IC3J4DfP
fPm8ba2BwAhM5vdQmXpDFBLYjuhDR3bjl5Di+i2O3rdGPkfNCGrSxp21AN1tdgLK
fbqj/dm7FfuhCvslXMsNdPtGCVQqU3ElsiUFJo/ZMEJKjTgXXt7titk93vf5RRI0
+iiv1mtaTDDKfxSNaBaTKG7wl9yJvkaIIhfaZLeIN9r7ZYoixkZiERTF34/JraGs
j9MYJUtxEWwXdxsEu/W/eV9G9VeQ58XPO4T5GAWrZMh6n5XOavh2b8rztpMrLBpz
CubVxCnhVlrDDk0D1ttKm+GjF2akWJyHA4TN78/BdWYPuGtuDiYPk264GsGSDj52
FY7R++/J8nV5gh3KVqrMeiO0gWujoGMXR3Gr6+o/ET+N3/epC4+nHpCv92XIc8Vf
YmbevBcDQYWBbrP9jM17ijEnJOuLLEGXZF46v83wl/tTwlp26hYqF9iU1yxeMnxz
HLm9ojn1IAfkBILRXIQIdL2HToPdqUuOT0XUp4F0uzTQ4ga9Rmamq1gq2HyGJd71
gLmRZ2ehNbb3vFYDXw6eFBd5zKJ+GYWYXbjdSdWVtxeAduHbQAyIWlmCP7v8iS3t
V+4IeLX1E6iV9bvWOERAXXMd6xnPJVwDvc26Q1s/m0IlfUuy6UKnC+Ju/isI/pBW
L4OWnzzWNX6RFA59FqdYbvgy1/6ZDWWc7UQG+8b7EJomHUiFz9859G47NT7Q+wgZ
CBiJMNkNwwiAKzqyHDpA13RgrAXkfQCTMCHcL4Vu9HqC21UkfatPbQMJ5HxQT1HL
1e0jgwlvqlE7p3Y81XlrVlNOZxxBJLicGThfgHIVPknLXhF9GrmtqRKGJEPVaDgT
mWJoDS0MUYbmkMmxsKSUj1oYlKuNjA3fUZ9P2OGuX7Gda97V6BrTEhE3Ksp8DmSt
CkBuuVzk0gnoRVsjtYhiA7S9ndKG67w2skKuzgfdZbMmIE3helinngyUESlCEB4b
uyAsyPxF1UU88xcFQlaSBN24wlOj0BdDaDFh7G3OF77TzS6x9BgfKRq9Fe9B6R8w
odk+JEoJ9ooB8n8D3aZh5mPCwjoKwtrZ2DaVFgvaAVudczOWU7Qa7b8zft9Stp8t
58WIIT4B7svGiY7G/Qr2uP7M42OqcU9O74oPTUjMWN6lncX3wHdNWBpTYSyEUpwu
Vk5n3OPsoGBluYhilPZjBv8wUidEHjIrKF6IN2mJJ2NmnwmoJfgw+I1VnrkXZEgT
aHF5KosQurNcqeSfvTkdptahPhF7xYUqbD+02ZSXCWBzaaFIkond+Zpx5F6RaAjE
qZHAlaHUSlrKaaPOKG6GttdLXjmK3z2ko4zEkH6j8iujxL4hiKy5gesXiL5CfJe8
40s7yFhndGZzTgKVr2nx3SROm6fNJeSf11CHK3YJXRQ4M6y3dpls8+OVxkmfijJg
syVoY7eEriEFx1y4e4khYWtzFxLIfyr1swcY3yiL8dQBwH4NuxTMU9XOIPTGLU51
8U/klTHivJY27Qdvd/vNmBB6GDAXWo9jKDYrWMrAndmECbWgV2N6xGtlV5CGnb48
LMEX0OGhD3smdquB4H2yt9AlO7FhRPyY19fOUny2X7yT1V3dAVHtn1GDhtODn/nE
A7h2dbb2McgqZiAw5Rk87W2SpnZy7U4+EbOldZnbBKXo2TsiTR9H860HdcH/Etm+
/aYsYV5VEvSnFNLoOV1Ok1xmYekDV5xHTaQBDAEfwNPyIX8FK88198sMbPNLjz8O
qp4doJn3rBSGk4g9G664enuM0ISznDAA9wyR3OUEx2JUH4gatjO+vo1+52Cam1Ao
HCRJmHs9IwF3CP0A4NZpbGiwGP/FOjSVci4Y8ADwfF6GkY7tRgORSt36n4n/x9Tm
0tN0DU1GEGZwZEA+HNvW2yuGXK7oVe9aEtC5l1McCDDqrceX9RmQVB7gW9Qr6UUG
9KIpB0EsL7YFFq84HyrIBr/ryQoh9TarGnASMoEKbnKkxvyOcEWIUHyynxwrl0Su
YuCsu8jqkVEIlVERCBViy3oAufCjDddUqWvJ5/LiO0jLjXkiRr2wdDW3SpoSdIcx
VFpK5Akk/9swDTMnRRjhJZ+PeB16Hq/TN3Frs4nyb+5jLJ4cA2qie+5KTgzJTCh9
nV2zqMws965Yi0GgZQbOvZeioa4o3gVO1I8NPH0273hK8SPiUJbxIvlo/2Y7JV/F
cc86tljRjAEP2ofsr6SbcrmOntSqZO/0AFiVFKpSWGMOxqAwEitNu7/lFM5sG6Rp
9D2fHHt7GTMXkUvtqGe6HSosgvb+MAsNIpIJdyKjreCWrFjMJthdV9qe5inXMrIk
1wtVdkdI9pGK74ccbD8t7ZGEbcgcC4jNBTO+sfYA27eqKamz6vQB/j7+r2ciLlGD
Sr5tWJ+lo0AaS2UX0xOoNAFTgp5rZ7XkVcvR2nh+NKcJ29MOsl0MQOlf6AGGn6nP
3Po9JTUKfrI8dI6fd1TMBw0n15Lu/Chdm2czByc1Sf+n878XIRWoapoyvvVxJZS4
1mOr3lQDPxA0YqztyYFciQpmCVBvs8IkI6oTNGZ+qmR5rodJT62I8tleplR3IQ/O
4RYD5JrNCtYJoezch2micvzfmtkfUjCVl7iegJCVdz4Q3RK23k2+PKfiL+wsDpIm
0rFS5Vw42urAHyM5GGQenUJQ6VrSBS1Yi8LY0h369VJtgNEm48jSycpNcUOh4oM2
FwmG9/gmPV7hVpDm7SrdGgfhz7Xio1Hh3kFI4O7TgGyQggVMTaY/Kts1+VZ+S14t
6V5W7Ubr4RntXboJXWpDiUFJ5q2bSmXRnBtO+XjVv05oGvbOS8Q9kJMdivgsJEyO
w8BOmnU214g6fjiSd85K+MHe/9Y8rFEGojhiil9Agsb+kK20Zkqs5Lna79B2is6d
lszYgK9xopIaV9/ztAShMX8T91SVZduVTYdkQKewebNFGq4AvzZXKV4Y4Wni0NhY
2Yg2qyZefrZ/SraeInXiI4KF0HkrvndlAzowB0OoL/SgndMYkkTaZGzH4zM00p/2
ajLkPiq/7lbTp6oLhNjORn9dLNMNp/3ng+zcLrseU7NK4mxLfPfaVFw4uCVZWAVT
KEe+qHFkg1laqIW2q9LZOSvLWoPq85pI/SNC9UCU+7I2SwcL3+hBRwCqXLW3lf5P
kFmi6YG4HmCTcZJMH0hXGrt4tf57CdGiloCm5MTvWf2X6f8Zj+g0YJau95s4A6RD
jXiNJXY3HGA+NTlBLErPSdF7R3qATO5qrM/ZiDnhmAnRAwZdd1nWabo/FhKUTzbK
NopCU8grTjdWuLYq0PGnOCr1ziRajS4MnUDFizwtf8SC2KANxCR/IDw+v6c0zUbp
rVPc2wmsCDbWdDLPhU1taBQflvcaj86P5eY140rZJtV4t9QLmXvMOBc2Eh6wfdHT
dv/IliyBrWediQXuuhCFnUwIhlPI/kjpEeTnWtm5QAzw5Nu1bqnT6zH9eF2SiMQq
KySNNkZQOnYWTFVCYfQocxj+uuIC29EwGq0UNkgzUMI/QOAkgaHGqVhUzAJPq+4J
RIjKXQx19spQoernR8Toe803F+YN0zF8ugfnijRZ8JPWw+pjJYIMK7h4h+CiHCdz
57PZU0W6gsmU9yY5LZhmouV+4bAXylFdjqQsMpJldRuZ2Cxl1SIup/uRDfYSyOlO
A9X9/8oAQlpa71p/pIHpZ4oTfBkv5+2AOA9e8B+PXBNswtvLfjd1D4Yb/v4vtynZ
vH1vMpTh/hYHtqP9hY3eqJIsjZLhM2HAaDqXA/Wk4UUplJrk50eG6/wCvSKlDn5x
hGO4aqz7yvNSb/td4NjDNgrahDdWpxJn/wA0S4SI4wmlRFycafz5UgJS1QOsu1Z3
Y8UTXQFdaA6OWj3seU6wOrp6ApB78Pbn+9Byjq1/2Etb2uFdTns/DiKNiMH/veh8
+1woyhs7ZbcDSrXBoM3CoraV+Td2N7AaEFvz5PlzgqWmI3KHHqmThPG5uACU0uTs
Jgpz71DcRgbqOu5zRx8yzSbb3eeWrhMv79TRlh57ZFkKoqz1Spj/k1lO3/3EJGXw
lW0D4zlpFbYwkT1939BCizkgZ292UCH/EJ9kUhDb6u23jXwmy1xI8IrPKI1lqtCt
Q7k9NDslqQTMltzQXbeSAsDrUXCLlkRAN3ur0U/B6w4rp0Sh5LlyVdcMj6b1AKNK
zXB4rS+eGUv9WkDWqLlgcbcn05kO6PQ3nAI/mqLm3bD+rIeVDVxfALlgOXeMVSJp
G2LOwxwMJfsh7P2QrRZkStyJk0bhkFKKuhV6IGbuWA706U+gYAuomjoXImfl7lK2
PU+96H11SFE9wTnOzORN+NcJ3W1S59n/zDND5+rrOsdmcrKgqlL/i133z/fkfJFY
obil4kCRBatqdFv3oh+OsZS4BCWE/KuAD4Xq1je8O005E3mRfVS+mZ1XEVGtVDpX
dwWot9ENA7CuEZTOZo5zoTre2uTlO8Z8ucNi0LmJu7Y0xWQFVSzBLvvAhXUl09Te
7mdRwcn4v1M0gH3YYoRJOR8sgCHnM7LdRBwkUQuVueKS5cVeyZm8kVHSZAE/+h8x
706lMR/X9H1L9rFXL7Jgnd6avIrz6+zc2/lmELmFBpQBvbR98CrCxlF2FNOp7zh3
y8qYgfY/vau/6mOFIYaeAmeWIagfbNDfgQ9D2h1SoqosyIHgJQ5eGw659T+xBP88
hLWa2Vc3sqLJtPumk+HFFamoi8SxHddbGUOSdJnv/MRl0Ox78uqWsthOJ/Yu2YON
5qoWNqtd6Uqh7lGr2FKj44lxgSsPwAuMZ6/iNPERuocn5ee5G11hLpVplRB/nIVl
zOFKV30VdIOx5rKJiHR59gvLh6Di1wX1mMUdXkIRaIg8VvqpFqy5/2oCpeP2X/oZ
SPuLjiB5Ys/XtW+bLDWSeGsurSdiKRp8Mkh66zqZTLuv8Q72E38ag5M0J2xT165Z
nZDyuSrP/3ls1Hi9x0JLzeRH4X7dMsBvav/duvgimq6okjzQD28+PR5D4YNUx9v6
qyyptX/1AwqnFfgS1PNlE9PwvHut7NAZHMxUdIzgQHlp32TDXl+YG9f0D5dch44O
bbPxJe5eJYKiJ+kQO55f6nq/HE9sXXtQ5jn4N2/PXj7PjbC349Zhm/RPF8oEetZY
8LThXlXvo4cLm+xZ3Sy3h2DBnaZ5XgeXTNRRy9GbUthwcvRNURAHW5/+zWL+/a79
CiG6ktDoepCDSKYsZAc1H0sBTlipemTmonUDviCT2Duera6atoSQ4gop2LQtt9VB
UK4KIATl620SzdPE6yaa77B8CL5ih1qHlw4fY+ngVFABQYy7QHv4bIHA/XIaSQdC
ZYgmygV+F+NlGNG4oyRgrDikTW6Qv9btGR2nc6BKTvw/QfzDaabA6QR3/DJbGHI8
9H+1GQiDb7XA2JbA+W4W9Z1FiC6xbmkMUC7UyjZw2K7zid9GJtsMwj8fUnY6FrQK
TTdhOwZdmQSGrbZs8IQNXyiGpHLjEA4UyCyXnxCS8LgXPPvZTl2rbPEx9QQOZdnr
JnnBU/1wmzGY1j/OqRWw6ZOEEDWsCQgsaWQUhWbMuoXVffZ0oI10ji60Av1NC8Lq
woDu4QiaBNFpf+mCSc3zXa4YB4c+WNaCaHePo2rk468eKDVwar0sELrHyfzR1wUf
kh6KQyqrZXGHIdLsHpb0xOiVozlbsOr0vOqBFS/EgI8nHRf0qNj4k3JupNSm488J
WOYGVPaKFBs5aE8uVJ0HsztdZYbjRo3/OItudCjLDkIFsOfZ343IY9nBdx0+4RCY
uYv1U/+EA0jzic+sAodsayau0o3dYgmeiNYqDgz+JtrCcnyZj815OrP+1/aoOXdJ
qOXwDGF8kO+u9J4TNTr2B2rMfMYdbOYVihn1rKRdmO7TzlT03OBOrOtVfpTwLXXS
OU3HEnzH+2MosSD6V7n29UelJ3OA7Or4odIjof0fC32b7gw/me4h1xnRDAnUbqbF
L1Xy0hqYMn+Ym7KLkKtDLJ05N657QII2CppsfN8JfuBUmrDSzY0g1U24GV3LZ3Hr
gSMkUlwkRgX9diZ2TXHlPELTzTjEyXQjhrCWj2r8vXH2mQ64wF+sOMD03bwFBEtn
vJlmCKq0uHDD8GCZ7RlNWMk8Wh/rVPBepIyjSI7xw54PGpJL6iodnZActyjP27ym
t7OBd18yqQzdrYDUEubbhFcmuFCV3AImJNWYgfPf/HuCzmdjMecO5JemPyG+WgwG
4W36WhQfBds4N5+BrWMJBBEHR5J47FVwosZJ/ZolhUY5yFEQx5VZubMRLKty+V2d
3gryjNKs/4x/oCOxVi3q9dsA+mz4cwDzppDkdohmI25/xUjkLxyGTRsu2EqvI8XG
uFW9R2xjyHfOtZH+2o8MvnonB0LbAJ+ecFTx8rSPkotZIeYKgGk1o5UikQgPE0IS
GomhXsB1r+oY49j21E48cqS3b6FJ4aMr2+RwgdqonHv7msxZ1AhdG2r2W5PZVnm3
sGXLmo0FRJdkQZJNG5TJq78MX41yHc2ArsmqzLYxzbrsaabul+ZsNcPC0paYtUzV
xwPSNA+n89hofmOeRh8BgSrichH/cn66Rhs4yrsrtjI9kK2dztixxWYbBuDwNboo
mr2l5HqkqmKBVfdqx8685jmS3egK74hiiKLjtAy691S2gocphhtfgeYMiVDv9xDM
Chxm8CoH8txpG6ikKqoCFOfATBJA37Luyi4QPznXfPaOs7RdHCsZQKFfMAYUAdhS
n+BmFqPoaSLrj2GyHlCQnyy2sz6ogCxaEn4tpljNNB73+MnNz85JANi8POHI10Fq
Ge4o4cNGdm7Lngow8uj00VU/MpXcaKctOA3Ic8ngSSD6g4tiyEZiHBkKsUZV6QxG
wGPBSszSgIcQFAJNvKfranyeX1cPBkeJe7CgxndZx9QqKCCI0bSt/rAJAYHZrFu3
+M5p7ZmJYAyN/i8Jddkb0UV0Zg1bhbgTq7HMzIaWXHiEuDChmM4AiIQjBckdTRlO
XH8Fnvmn9zKTpawr0fdjxU5B8NpgZ4VgZ7PRmYVD1OcOLcSqMSGOzGN72O16U8kL
FnIaIifbDklJ3RkKgB8Gbty/y5zTc2EYf1YKVLgvOI9EBXAu8Oi22RtsVo7AFcYD
xSS2+1r5820wgtKmrHhav4Fsn2HRMJm3bZqm5PkbasSI6yv9bIba5AKrnP0J4jSh
Iwi8YomkaDm7zYeAfd7DI7D7txGZVoqyzMmk5Zb1Ja65H3tL24bDy+2kJtmCsvgb
vPmeG1jni16NhRQM9jd6pdV5Tl3tOb+zScQODVBr03XSiqfcg7KzAlz95xrEr5dh
YjH8Z6yw+F3YoKqo4OHcfE0qs2XvN2l/jOkVSNRU1mgbh78dCETXbMKr466vbrmx
E0u/kydl6wq9Q8GZ8ztPWm17JugeRT3Wbi6mqnOVCKYxoWxdl7P4rMFx1z75QTt8
wpaLhtZWNLolp7osqS6WYn6Y3IH2n3JGruDYZEjTC+PKQo16nLJ+xvX39FsPME3U
ZVmIXQ8DuEHWS2Gqs4HLlrPHiQ+P4FtB/uNPhnLwq1Zvo7pZikOJqyaft1r74cie
tDk/tLNTzrQMSYQUwHC0y/Dmbjh0Bu24u7gNqF0fzY8RPST1kVM+m6yv9SFlMZQU
M10wg4rHY2TFW8p9Fww3cVYLO8SXxOygPvpNkwuRDBw9EW2YPdgIE3VSTHaNvQIQ
ld6AJBEfbQNAFh6Poh/uwldgWxTRhN9BaDir7xa5OUGV2IA3spUWxg/uCrO2heqw
c2ablMh9Skz7T5SQ4cPp1v0AlQVt1wkjQ14i77xE/lYvTrHVqHJCfFTGHKGK3NC7
dKC/FqLvBA0eghKq7CztU5qazkVUe78tFrnus7TXj53U5Altaoo+BEP+nRWBrHr5
WM5JyE1hWeB5tWl5ik+9NBknaMUzaHUey1ZWaKg2eknA346ic+VeEEpD4HrnjnCA
a1XJXMZd0BmnRQh77DHu71/l22HHLVvlr5TIzLoUiPNdazFxkd94gClMJSioU9fG
lm7wbpsZ6gZqfU23vOiRnx4kcvR7W06agT1wq7RZMfm4mehg5MHZMCGUjgrraaSS
4kmBnvOOOm0NvRfaco+yD46mnfKKJ6AHno5HByowgO576fbkAs1YQ8J9k8y1OOtj
QFjslwRADFEI6PIA9/xP9bDPUjUH4mGvT2neL1teMZAZQQ/dZ0FEkWOAfhH2Qg3S
TvZk0fG++66+GEHM6B5YJUyz1sHidTOvfJpI9uZSjAcNRIsGzuJmQ22oYPxoaeBD
BOhQeP9tnmTwUJegLm+yblyQjVxnzoo4/CBeHGjVgd1VeV9WvEHfGqNJY0yJuhll
b0UcZPdbD80kPRoXJ40/tpI5qCFBd2d/gfllIdpkZPctdwfULZ6QAW0DsVeDrmS+
Of2GgIW0KMwx/Seqss/Yj0F6CCwIpdDbngPOJ72Bci0jumEOWQuD80jDZ8GU3Jm3
PoVrXBm7B5WcAdPVTrO0zXvM8E5jukCpEB7PKew8757PpLk3w2asgYDJ/JBSQ5WY
bZfIL/yZ+/6TuiGIO2Mdg0/IbBJx37rY7ouEuCgqMLr57yD1oH1U8zG7+zMrBSIG
d9fP8Skd04BjscgSGOkhG9lK1xD1xm8Dniwqtmk4KJRuM0XgpwAkL8AqxfDAxWum
efXtZLIak9L32nbSO86Iz8WFReiwVwBtSsTEuHXkhUVhzV90wZAo948ZGDGQsyaD
NzUH7t+ud6nhcUrCxWjl7cyVwSPOybgXuPijCc4LCzvCx7BZ4CSx8lxdoX1z7urG
KpbDoEBPVqvIs2bb9iO8iHxie2YwaerJKU+FcGDGZMSD8ydboEs6gq5RyR0iHcac
1rR2SFkqrfyzVeOLzYsga505zT3v+RsZTaXywPXaJImKy9U9pDCTA9tny5xDpnpX
o46gAGpGkeWurHlHJml130SLRwVwTF+3lACjKr+z7I2G3lA29VNf0d7OZWMWjpvN
yMeQZq50vUUPoHwPeNQgPL8qPoCJCKufnrPIz+AdiO5B4oEKbl+9jBzwat4KXBLA
m42V0+5xJT/fhmf2OCkDBDaltPSkH+nmq4e2vtu4fiulD2AgXWZAbZsgjQ3jm+r7
hOycHJZ6DmjhQ2gRlvXJ7oN5qMVJJYEZEtI1Kv1GuPJncKJUULVPDqpYi92HocMY
9xtgMUrJmLjQz+NaabIX4oYXUw2S6+Zr+fEudculULoq8UBrkLBIYv5neQvJhBMP
X9Zd+04FN+MHFkE1wWWAnMx8xEpVPyYkZlQ/t7/c2rijtWcx6Sjabqt1BXkVmm4V
zsNNdH/nYR/wlIwNL554s9JGFEoG1KSr+su4+i25yiDkX+nMmJxxJxqzTgnGfFcm
tsodjReaOE8y3n6USUI6z35BVUMVpNWAdfHuGPzUTckftajiukPysUEj75ZQZXyY
dEtqnh0ppJkbc6peuE9EC7irBJS57COhnKZE/iZblxgyOhcsyWTIwV+0FV2so4cx
lpl/XMocIBqu+VqGV9yCkv/Emvrr2SlRkKv78hmyeRkz69t2CE0yyVq9HIpLzNGB
eyjF6Vcq/+U+PY4qcK7cCxsFF1UheTltpFRWh9q0R1cy/6Q9q3x7maQDiXGjQHBq
OPlN0oxg6L70ch1ibEbaQis7pLuvwGiYkRlpEYe7Wo5AfelT8/FZK4YNvxP2Bx5u
VIitH4g2crN9ymScPerb2MJwiuqAR/IaTnLLSk950uhAKMpGgBTqUCc52wLGJ0JW
hdfL9uLjoweWSF1hKzcSNqMxD6Tc3+SeX5lqz6vW/uejNKrtxZjELGhyK5IABc30
urB/YqevmdxRjC2GvSQHPnl9lRZBvsYRwBQ5PctQN3DWmja4YW9MmaGcn/le35BL
6FCb1e8+4zlJNoSVQJgLyc382sjam2suEIaqjxi3auhEaTI5rkDGoy9SBrxcks5L
6oN5LqJHqaoYYaGX6y81LaEiJwkZKXX2oEukjHjqVFB2cG0/InBHVu3Wh2jFwJge
JAq6OtpyHbA/gSkfkI11j7BrivNcAkcYY3yRUtP3uCPkghgfLk10UTbI9/LMqYCo
PFKXBkdeJGBSLlUEH4UUgycIHr3cHw0bXF5pV/bfWUSpxQonRLKuBsfXnI4j5vgQ
kwHE7bZn5Oe22snRIOLJtswoweDqPBQTo0iZ4QPDEsW9cULdHhfqivtMICBBpguo
dq+anlyKBnqnNruk69zhLrxkODYElklRBBUvLOwfdbbKh0iQNeIu801zxR80ysOu
+Y/cS8cZyKn+UYcTCx0R/8JgZXBVaRXRAJF3K0RlrGkoa7jPurQ22g+wA+Hw+2wt
NwD1tylbMp5GFECKwZ+ERlPu76hDJ+kN8IsQ+eXk1f8EecQuVuf5LmONXbWgQFms
042RrelCfvPQpRwyBhAAEzEWn3SQT5TPUzVpLPnyDCvR3tAjCFA3773HStDOH6vI
3/ofk3einZHxGbd+sTv79/qMnax1Sf2ivjF11UA89iSKi1pi8nrklSusbmcP5j4G
YMmO7YmcTgE2eKsZNah28a9TqXlQ+2qMExpCfjdRyuYXcW901oX+ev+U5cCBAPc7
hHyP1Bjf2lO+pd60Ve9AV/JxJkyhsBPQzokYvc3ybvoevWFtkDqzbor462JheA/6
LBQ0ikr+tKuySnXgPkS8kBG/GyzFNxL+G96Q+mOGez6IaJw0ZG4FlWdXaLpHVMeN
dCjV12o2Yl4mtOmzr77WlmG/sMajnyxEltVNAGZ/KBtzXoU/o+qUUlzdSPsfOQ81
+tRfUl0ZnpRSu8NUXIVj5r+5zZxzlZviHyVQLizngBHeTkYmi+I2WWFUF6T6pdgm
HhAI/0+Bdsk1r7txJoNPytEbJ6sJzYx1VbuPCZ9UdFgaEoTAZpBShJiKUb5qlB/x
ApT8htjecq9veOIOz6b2THkiP7Dj2vw5EO/Rbxho0QYsNIF5sXdLIOtyyfPgwHd+
duiPcRgGqf+USpp39Bw8VzeHvvCxAotFq+k5jWd8ldXPMuyRBjRcNUOy5t3aNGui
dEDSOzNURzd0fRNoLO6du+2FOGNR1DeG3BRvz3nTLYleZfO1aCPMpno7AGqkE6Zl
agTsNLF1XledZ5c4QSQcEbGgnS7C4YpfkG0oAtXs5CQobPs+9q2N7ImPNAUhnu8L
LTRj2xPWsfCmUbVlgX4H+RuBAf6/urKBG77/vzsOjEfJya40WJ/eI1HoTtnOC6JR
U+WLgQ9niNRtE/rHbtd7nCh/7sXqP8KLePJbs0BzbHV/hyZV2GSdTGlsAdGfCf8i
S56zmQzeqbIKBwYTiBg5JsGw1QiDl+InYZ0A0dSeRS/WACXGQFSpB5zGpy5kQ+ro
cFvhZEN/lqVqUTLFCPApuKiDPIGI2WYEKqXDg5OeRqs4R9Cooayny+YHp+X0GfyA
5knO6eX4ZpekpeibLX+ZIOsSsEm+vYR8XErcBq3wWZvSC/OmVCfoIpKN7jmkTK1l
eCtSomIn1/YRWY9jHtUR4dgG0a4Nhd/vgMHkH8trPnTz2UT2QRFyLPVtmhicDygX
oRnFkmd/hYe9YJfjW4yhRWRKzQEuXKVuuvfe/5j7GMDw9Ul9vBJnhMWlICmuIoDh
BqOw7xUYqzRMPxYBdXA5I4/FvlZ2c/8hexiAYOx6Kc1TkfSF/a0TLtH+zBpmLPNy
2IIFZnacYIy1sx2fYgZexCPvi69adPwkA0UfJHwygiSYvetvGchRGQUxLEU0fKOy
0csUY+aUwwqURjM2eiKYD0OOe/4LTpf47YSdBKOiDKfbgBAw1L4RTV6N2uoEfECc
81qYb/3sjCKV/4eRFb+iJXVxFyMc3Vm4d6gbuOtY6jrv+nKE4sZxwIkqzG2QiqwK
hICIypcA5aE7k0CBT5BOPgP8uTO+4Vq/Sf0jrXl0u91dZbuYhrypUr06scaSBgFX
XNc1QB6jRRdYntlwPVv2YRezqxli9nj2h2Irw5ltxbXpK2foblaWWwUxeY3CeZbv
W1xSKB6i5gD+mKljJbDd2hNwKFyc+ZszKlJ9BfMFcx8EnYnfDzyP3FNGnE+gFW+k
YCSfXNdAxO6swwrVrGle9CS9U2IlvAcR04wj4Q5jgVJ1QXo+o6ZeBagFtHWmwX1T
FssuiHhdBG7b0NdAwY1DFHMiR1IaWnPjvDalgrUPbxiuEda6CC1+DGjl5JeUMzTF
88RLJuxqtvVksdPjwNio5CQ1puuQKHtaIrYegyUqUbIrKU9UoBrRsM1AjNc98uY2
Y0WYT/Oy0NFV85CGOD7PxL/yMh6aM6TeHTM9qxE/bUWG1b2ahHDwPxK7AcO2XvpX
ggZxvD/NE+XPZbk5ltFXLGP1WlMRaN23WjxZp4cWXkqSNmcb1qC9lJlCru2m61uJ
ifetHMdnc9AKlms+cjcLJAqKZLkBpNyaFtXfi2n0xSlfKmK8uvguCxV3S9T4E3gF
mfVBECDM/11oeEEe9BhIfBgIfD3/hs7WP2f4Ua4jJ2w7BhBBSRg1Bq123SsfdfY0
duSH1JTxdXmgpTeGFtDeebVr9cDA5sOoj6jTi3b7PftFjiuYfyihBlrEQo4/p0rP
CIh/A+bCWVbCZRqmKHn+C9WTzZFO4qGV0OyV0v9WnGiZbid7UUdvkzTyCKDxS2JU
wxDR2sfcc9ZpIzQI4qnNXhqAa34mybDTC3reMY4yQJA4NL569PNNq+g1KFAV6c4k
jxt52m3gt6DyNQvv8pEw3zTvXdV4Tuu/T+aZ56PfcTcurLQraKNHwSkT1xVRb0Kw
3FB2tgBp6g3ctAVa/Hzsv1EAVLlkq5YdvQgFBlGTEKzoSBX7srOQM71Y4mpV37Zo
pVVQLSpnzpqcAuj2L6gn6zvWKqUu8HyO+fCAMLcjnDNG83e7wI3aCz73zfNDdFNo
khwlDbVSaVfSjcS7d9O7rSOVsHXkfhgmmGuMGRWdJIziHJPf1IK2BrGmw0wB8LSj
BxsQ2D9fKdTo9IlSDnIgl3bThCYGns4oM4rr1cuUNyCoj46VhnwSDT3qbwwKVq+Y
3CQKvyTo+uetBL0m8eMjuy8J+OmQ1VzW9RLdKeEdO3sbIqc3UPhC2x/S1pJcyiYm
lpuf5sND4Fr/li4CJdIjUhso2dZIk8N+5L7oDF8499eOUDaNKEakTfjJi8Opsmzt
ok7JCKzowJ6OFRiYxAHal1l9Adt9rXHkjjUf4ZBuBhgyTgjUTdTrzQOV3lo4cfpS
Ee4FYZ/zjfU72Av9/nTEXdp/6zfNDw6/9lUvNSTK+V84stLkcNlR76wXFK5RvB3c
a4nGmrmfUpF2CFQvX9LMbv5zpbGkvgEgCL+wxWeX8QigFfUO3ZQ9gAhPl/nm4r2U
ZW/YOjkXSn+fklfOiCP2Oo8R+Z17Nxmc4ze5STpgxEpRDD/kOB7aXOV5v+Wh1omM
f7Df4lqYOl2nsQ7nBaL0pmS/2BOSwFKk0yvUtot6dujAib6y56acXdjQd6ej4IWy
nUQQ8ZBTxlZ7Uhp1bSvRoaEWCbFbhumE0guE0gNMr8Tk39wQh8a3/LAvhaE5mgyD
MFG6ac0qvPDyRPNncy3hingx79XiaDf58RQV6B0CquXTHdE9IoGlNpRhbzIwLMh+
v07MKnjKciSAgO/btEq/Yt48XV1PYMqjuhYJbMkazKdOsyp+fMithZQ2mkkmr0Ql
vl5Hfhm3SBDVLa8vEqCClKutiHKNGS4C/tp8lQouDO9eWteKjUCoSnIZX5Zx+7ok
Nvqv9kdkArgMRxMiCcZgF5PXvAyqKCWqioMmOA5SoZtyC4jb6T2uq/tQT0WnuGTD
XApKhmu9kP1n0MPMmOmKSI7klGSeBXTa2g5mQaMU7nBJ8WaRHLazWuBEmBb4gCgT
EawEe8ahzk+uaVkntLjH1ek9/srRe8IIK7z8HSWDaZzQjbJJPKbjH4ekYwDxkuNE
KB521g4LgEkmpUBCgAhnNKni8KBX0lw7WXLLrM4QJzETgc2ioz435RQS3/pbEk3s
qc7NV6TrWn7j+Ie54ui4pqEiteOe8n0AFoepOJ3L+ev584aVWqbGgPG/G2vEg6hH
FvscN5A5MEgCndV9YJfN5dX8CqI4egOn0P7ItjEwFWsSZjLvYJ0SD87IY6aSHLXK
E5jn7EZjqcpsLR9jyQUq0o7h72zDVbToxax7xCJayqX1FL+VstUoio5+qej4iZXS
1exQperqa3ig70FIOuaPlQhSbcMfcrQbrHU4E4zAFEtUKT/N2ZUCqQXKnYnbohwD
fGqcUBm306/drhb0EAn7muxKlRqV7ecPPtKd553MmqQMiuQudfuN0Qjf65fwe38n
G4Y0Ugew4Ts3Ky5RU+jxfV5AoYsskxuOmbDqd4QnoON2zhHra5SCgkjmW0Gjwf5a
XATV92VFX7D4F0SRdscQaEgFF4TFwrN7dBRioHmXXBEWjc99RpX5/EBTaUIgRQQe
5l/YoAP53TEFUS1yMarHXGT37dUGSVMOCJ2I7kCnoBwxrMUb2csBmdpuIvR09hpZ
o0JUGIxqPtP+eV3TurvGiXsQhNm/feqYXmKsHlw0aEgh+nMcH9GNOlVXOoJtgphA
hCOg7thQrBCTVqcTEHrSbLr50vpjdgX5okvU0sKgGiFAbFEIkbUQYNTtVBlDCAfw
8h+vTRnJeqsn9A0nHUyH0gbNAw2vOuQ1t9NXvZcO4ipswGFXBg8f50z0ouwqdLjK
bylJdi6afk6AQL7C3hBvJYpzp8pMiDhnoQoRYhiWB4tzXoylcUsv/rcuXK9JrmOi
4YQlKKvbixgzLJyCpuPLjPOYcbNhZnmHu5FNUqH6rjLeCu676QWhiq8ith7KVMeb
lQTngcdNhPA9fI4uvEmbpIqFtbnBj0e4TzR9rhqeZjJUn/tiAH+3vYqoZsUqVTEI
5iHApbHpplapVDypPokPUCwrdFglCEv214O2GNqiM7NyyAVJeKMrbnpwwV2Uz+zZ
VXDCC6hDVLXwnm9GI1Yhh7m3oCN0bjQqgsrnWle07rgXXnR0vOph2oRIxp0CI69e
1Vt5CnCDfvpGz5J7nsBnAtDklpuBX3u11RtkGEftOCLtuLXZAAe7z1A5maEKCk/V
lCUmQLtzWzgmJcPo2kz5hFfRCqb3OHcdfynWlkkyIaBlKYBF6OuhvpWYfjAiU857
BtBYwbbhkwUBWalvCVhHPzy0IFCVVMkHDEbIZd4DALza9YR+Jr2T0oADtgFwLFva
B6JlPNBazL9vNkBzZq9ZdT8dPXJPOCtES1yQl0BiNf4MNmNygNBw4hc4lnQsN6xm
v0kZqZvQuVjlHEbdkRGNFIHlN0L2Q4ek9luucc+osFqZnDS/A59q3gdTcZ8O59pe
LOWCCCNmD7tgBazCtivRRRGt0cKNfDPT7JNF1j+f67920TqZXI96NWgwKcMPyZdF
keVTMHlDtQJIOO1iQYv3bfvkCG6MklHhjSMdPMXunpNDfTtOeISKtqBfkmXMtKBe
NRVmpBKowXGWwlgnt93joN8C1we6F4aXscdPV+AwTmoKGps9soF3zFgN9DZxcJkB
uoE/VOMAbA+p45z/d+AO80IgA2YrwhML3yS0QMpj1Olm+vnbITDRUOmt1w0AW6SG
OajcnP5zQHwFJxSA2bQe7Q/MzesNn7Z9OwOULEG3yi9kl0V5XWUTAUYvlMW50EFd
J3wpcB8sUnt+cGrVbvCbeSPlBF0GhWkF3N3r1cVzw544Bj2CcI1nBmu+Mu0CZmmc
TUXKWyeiDD8YJQmd+UIMlrZQGuLcJknf1LrSUr0FKihrxYEmTEg9mtkUvb3nWloh
3KdVDj622VspH4oXLZc9C1r9FFL+tg0qZWXYFqLDPgsaYyDJhCh7T/MmWoMcd98/
vue9I0EOhMd9O2XGsyNVc5fxq4QfqG4/YoZpSyPHg+20RWHr/aM/PSGJB8FoRCO8
UOl7FtFXaonbLmiM2X2/8Foy6YnprBDiI/DnJJX2ceIL8iVgRUA2s8hHpLR68FUF
Vpjip6dbKxN+nmMQ185ZcwtuVp0zd3FAVSu6Jk5gKAr6p0wfP5oh21xI+m1gRGYn
PdFD67APuhP3VBhJ1iqpE92Sm2QXVqSXtBPcS0Pkmc0vqtODIlHoRmRP3dSDw3ec
+IMGBYZWv+FkaPXeTpxvdZ3niN1PnVG7CmP/KUcNdY3yMVpYGw5q00mows4Hq80I
lNOpKw6Nhbjwoy0IRyj3KLSGngd3Hb0ujjiuRo4dVnYC3IFb9wqhxebUyntx+jEE
PhZ/Kh6I7KFMS8IHJVtcyOTFuxKHkD+f10kc9vGyc5acCQS8PTI2Owx//FD2jdNd
S67x9H3naSmsoTTWEYl+UaLqiHzH/f9IW25xr4yh1Fl+y/pGe3hwaEj8QmFHyN60
zcddPXKLcweqm5YSqqOssxtI0hqCKsQ0ti0W7UDipS3vf01MZ/FcynvT5BdsClRK
dNNw4gjBaknrMhD+0qJEsaJJsNNhe/AZJrIcIr6N6Hvvr9S/mYe6zosox5c9l1HS
u2jDRa4w1Z07ldsqVKb6bvcykONL/95WouUU4wP1YMt6Xyv049wF7ZGAm60p/p43
RdWwKZJumQD8fsnQCKChV3Tj5utRmN7s2Xb0y5GYXfPGjVeCVUpbWhKB9JvaD+/2
c+xRaJv03Zr7lDuzOp9n0Z/sFQIsSLgR/Gs3NPi4U/O+3rK59/kbwCnMnW8oUJdU
RBnZF0LEsthkG0qChfkA5i/1D1Dz9bWRul0Wwwd3j44gpqoQbWuOevvGXOXqPzTb
P5F14YRO/VN3RoD1KX1wv5t9Ks1K5T2wf2kAFLQuvTnQ6rEU1vCGCy7yRtkpZtzS
2zmut82WPFc1yNeCyxPIDhQerslj0ZiA1Dy+jcVjKbEIZtVcv+cgiX2OZUtFY1ev
TIpfTIWxRnIu6NC9mndP4JOQhaDAN40RHRFYXOjARglDaBSw/6olUYjCv+ulXFFY
vGflayoCcPD2ZPivCECXhZVnv4b+ao9GAkm0w9hwISI8mclz6TzLw4gMdzdpVbIi
vDXDDpD3rBu89XxEVet8Svq55nZ8QUJYZuy+Pnj1Af/qu/wUXyIvp0OwEVwM25jf
pt0cPMaDr+p1sdSkVlf/KpgMAdiDdYH9vrTZ8xVuzONt0oAl5Pqv3VBNZaecmVe0
J3MKBeL+XVSTu9GzGXYK1ldvOI9Jp751VQnYyoACkNUAjRT9A5jTGY8f7KgCIgsB
y4p8NoN5RogERWbW00Mn4Bd9esDLvr5rnfZQ7jp6Mcm8D+9mrBvl15l20cExiZ9q
UuIJAB8H4VdPW4epRtnKLsz+XYDAfk64TsLzwH66cWnuDXKEYzNlrTuH6yNgcpEl
fzMMPykCa3cZOIWT8IHeeNtVF42xFC0/Csskag0HkYmlyyKnvxKBGPdW0EbIs1xk
+I0evkN1JwsuG3aEYNiKi6Ggl5TueWy9nFCMGZAORwWPE37/K5u4VeU1G4g+ainc
e5NGxQpymxqntbIlzqRVpQZcddBXQW1KP3cDBeijNhTYJmdPaMqlYV0P48PxayrV
bEFYM6w8f7lftb7Up1tQI5UnqI4S6VklfLA9AaYVbafQqGE1EZ9aca8UvJT3Bh2v
M84ZXhlFFdJrXHsiLukHjPj/G4X1JpU37Uu5kDW0acw4jtyHWXD2fXNS7gI/G9Wm
zqrfkMwxyQbgdTgDEVJdGb44xKqV4+9+dkx+ykL6J6d8eJR2h2QtZ1894Eh61fWQ
jrf+Y4QfQPTHIRsotULGpSLV7xdr7QLCWPchoU2MPzGD29QgWxg9tUmM+j0Ul10q
ktBCDG8LyhV98PWiG+dlwt0oqMdhS1vO34Ya1R6EJKFpSBlYScr8Fzq5P7Dyv/BU
+fnpamRKjxQrP5AAEAhhu2QZvGd5XH7AdfGlyBuzkk8Kan/G3SU74MtPWWgTEuJI
Mc7W/MsPQ1KXhNNNFQdMcCzaMQo1pKh52fJpyK1pAB7zPkyJqvzhIn3eSzBgRufJ
A84XI+4KUF3Bk/nc1LuDZW6bLrFrGNnOEJEm74izSZp6gDCm+25PNjJuNOjsQ73Z
Bzmy8uYS0IsbrIORwVQFkeLnQR1hsn0eRvdp1k3vh3NIWbsxOrYo/3xVP3UhEcuY
mUJxJAzEbF7FgbKG6V+4xGVrRalBasWECfCaUEmiTpiCb8C3cLwPnnDyxmq7lZnQ
gNcdU3Kb59l6xt3ofVWcXzYS/cGroWiA8P+J3zIYDxrl+8tES9h/mCLCE+I58A2W
VzA2o6IRL/QulWAS6/dWhHa6Th2vgfp2Uo3vVxeNTL9NGTS+OOgtoHkyc8B7EQFM
5v13aUnYnqO1NJCMrniX5RC8HhMad3FJ9ugLl0Y+xX3ocmA+DSecG3Iqk+fHE6LG
zU63Es9JRujTyoosDJ+I1eZon+NUguT4HELu5JDUoAmHYoL895rAsYjGae//44T8
4XL14OjEW/j/osJ7U9LuoQ6tDer5QNMWj6eHByOYtsxK04qdVRLr7Mw5iHuaKnRU
`pragma protect end_protected
