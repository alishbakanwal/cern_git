// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 14:01:24 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Cf/C6dGZ7+NPMP8NdyfQv/UDmNwWtC4IO/Rya+90Vx2ByjBec8H0JhI0+7Guhmgs
mTvNQ/bR2mT12j1Wag0/wgRNwQIaNF7mTIV0os67agSuKgiTJE0pW97c4ldLfyXA
tfyVh/N2Eq5KWqOESdJziqt1euQv0a0XGEOSePXFyXM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 69712)
XwidwnEWiWAfS12bzMXBvt2C2Cl8O5sKTODx76eVKNJYi68F32Z+tjbpU4MNJkqY
z7MUa0yyrcXP6GWH+mccQqee4CVsc4dmZLgRd1Y9o3XKrXA1h+4HjqOF3AwrSEQY
3PibNJi8/K3Rz5QGxZi5wfhsrYJj6Xp9tdOuzkvjI5rceDMEqGXmAqRzhgWsy44C
rNnkK2hSBlfK7qRAFuOkoCHn5K0KXB6rJrP42Eyst10v9hTz6Q69i7t3manBgb/X
kqBTC9np+S9M7bQiSXL8he14VYUQGGQYdGtFgxdP0IdV9QxctUX9gljd8T/oVuB+
QCRWW5ZpQQpo4eep4Jnbip0xOUflbms23HYwHImz/T1YasROHTgcvfA0Fu74sexO
7adje7MZCMwOHLWCc8CS1fFKpCYtrx8rUwpEQgwmzgdHVj239aAMcgUL/dz/OiN0
9iRBW5/JQnmbicZ/yzOwuStSk1RBWx+yQp949y8jiKBZCW/sVFqN/3Sl2fgsfvDV
R+xbD0cUfyin7mcF4YHhbdi77jRNiH8mImqfMyb5qk5IV/s/ft+HptSIS2R0mvA2
USd5pm0szfAtrYF4QmFQzq1qDxxOJJgIh7H01xRM3wrm3OrY1fYtTWNpOaW5/l2T
B3q78C55QaIcb40Eq2nvp4POYW62bvFmUNEN5vPWda/0d4uQ/gtz+IwMl9v/arYT
lsS/eCIq4Y+q+GqwXJtgPJRjtmEmzprSZnGytyFyJVVmdPB1ZCloGsrnz/xZASB2
ErRS/76+JxkDorquj1dZFTAXSI5dRwHqA4oErw0zq7hEBFjd+hSPtA/0W4ZAEh0g
rb80+wGOEJD2hCECLlpHVazeS6rv7o4y7vSqDuF/siSj66dKgMMroNVVAEUm4E0a
1RDss2NO4W9I8D2J7NWexKvMLYfr/eXoK+Bz814xffqIACotizJfcLs7NmNCNEmi
s5QIR7oFaQwKzKuo1EEPR+ODMy+SHcg5sZXfQiqlQ5ZRHgWOOi8vpA1OD98HHeF5
zm7hQFHZ4r/wora9X6rRU6ReKLCDdlFWTycPsP8tl/6ArtRiFhtCKob4kyj2WuhD
H5chHbXU3hM0CDmTqpbOYj6pxxgUoHugRO8KSvezrh8hCNRVRUuuMbZbzI+CLU52
oNOvRR2MpwhjExMt6p0vz/1/KpK4vxMKosURDgvzgO6UB5tKov3nCu5O6bvRnzPH
7jHVgfddfLB38M8fzBnU07xvyPJAow7715uwrhzBAdks6VFFVnuSszp8b5qspapb
5fzIpeiDtDEltV4vUGkVnwfAiICNtzcf8sq02TdhuGHFogSvpx20nokU33ZuRKTr
edfmO3P5gx6F0vgXgIKJ7Iyz0Mf4MSEgqDfcY0FqOHoSBvAfo2SPIcJGIT5kluIU
PZTlsk72f+3Z6N7XBcDM5mGfyvNepJFkcto0Dp7b6+bh0+SIC3RUMQFb5Z5ZzvQh
IRiEZiXpqWy7eXLzy4ihCPkfwaHsz81qmSLp+SnLKDSlFUAc8bNpg6AVWJv9Vyz9
kyiDuyN5O7LKdQaDMgtXHkMFDLBOmYU2nrtGaqgWWY1Al8127WmcWkE+uvm1KUBS
9vJcuEvsZqU3GAANL/2qqKxYq86IROLxTFFaPlldAKuJwm3Dt+XQg70FW6dt6tH4
Ic4bXDY+cloCQfwEWu83Wp1y3aNnIrwOPHyH0TX/J8ymM/wjFVYrPZzcRlJRMInZ
/g+YhkDhwofoj5lQxW6BwI+hY1egmSciJijnbocn9qtgWPdkJQdkzjuugdwaizI4
DlN/BQkBosOQpkaTKPQdJ9w5KLiovLJE/cMnp88CzErRMtbYg5T3CcXe+q/KLBOR
++ZIesCSXI3HBF2M39nDgtT7C8Zr01dSXm3UxbzyV7ziuIYE7n28GYFRJLJvEUpW
AJGw6sWd+lpgVAF8mb3hG2zViceZWWrpjROthTsM3TrwirqTe5uDjX/SchEmegb7
cQAumQJ5s7enbVyaARG42FSdJCzLH87QZV9F64Q+R/vdNlfA8lZDVESBFDHnhKZr
XzhDjDLui/eDG8pN/J6UKZR5TeUqsk1CQ6MhOVGMTWiJiqWfxi1iw3CNz1di3b0T
14tMIYHeRMCLxJSslE0jMkdKmS00QGCajxkwrH+PqjlSb8F5C0HhoUh6VdLDI1ji
GblHrDl20K/SSo5X2TA6TBbnKK8vrIN18sTX/7anzX5ahtmFiwhNV8Fo2nhXa8j0
sbnRyaB45Ns6oOC+7Som3WaT63sSERZ027SyWKElhacxwwk2oK6N+h+gVg4MkHIL
ifxfbH6CuND57/P+w+g/tYrVdnqO3NsJHqmiFCD71W1tJIxoCgsooUdfklEgzVHP
cyQBd+xkwiHiKdso+XkptRg8fK2h/QpF+cDp3ejHKnBE/HPRSrTsmacZ1duGiPMg
v31dUqJCV4yCyTkBJQBwdJR1B4ZGO3J06+hZhSJhqMnlEp1hlrfFfPBj0+4S5qXm
Cast7T0SCC4N0WrHiHSluioJXasrH9t01ttKVOojCnlcVWG/GyolkFa0k4JLqxdk
n5QgI3X7Vv0P2QAnvS1BqHbK6Ya6NH+BukVCRPiew97BiYDX70I67V19NBpWTsmU
pC0KjiFxS6RvYruXg0PDrmHW6LJh7nMQQBv5sPIS9Js5Qm9WXt5f9mSoxZhRTgNU
u8mFMqaggoFTPa+uElgE8Lsqa2Qm6xPBhBCWSkDsoAUGUmt5OHpuuH6JagUHoe3k
BhJBr4o8pR7sSGWRX4HJZq1uIMJsD9Oi7p4vtlWp1+AuSaIXdgXzpce8Zcur8MbE
ajGdlTpZsfFBx6yDzMXvMfXzAWRRMxGhwVFCmgYqMgiCXwWcc8YacBh5tABsw5/A
TqVxPm/dk3AEnPneCsrjY3YHKK2I+Ug1dUYmrPe7W1fNb/DS3wFmIASkzsa357j/
qTU9yVnC/RqS8sZW1REIaQhgZRutULcO50bcB36CL7KaT1WKmHs7i1Ld+205tO2F
GnQFoaGzByQz4uSEx0pTjc2xgv0/DD/pUaiDWXP+nBFYVuJe1PQSpzBxa/wx+qRC
3ICB4g+ufCCVT7wRugCEbk9uRzbxwpMPmdrmvoR6bREpUVjFwZ7CH6w+r6fM7pnG
tU4/k36M3H9hxH7pNfAIq9fEMy/8/tXgZDYCwXf2H/TMMXZHcdkZyRBpUKE150Yq
HyncLX5tlOpJIx8eK4pqh+JHmENVXfVPqWVN0OYTqmRxTL9uz3YfOgtTZUQK9VUx
OYhezMojOC5DEaTqGHdD6VZB8APotfTUqVRman6deH0q3b5ztQ2mlOVKiVlQmEyK
qUOwZCU/JpbHB7xWiehZCRat6WsJliF1AXw2elH3irknyJrFUZDWjpOajos/drtS
5hIBK6n/5j7+UdafQlXRGPWP7xRTLsqR8SB95Wf01w14QSj2pmy4rCX/GI0jPZdf
RvhPrOlnlr2gVqpDGWW2xHhcQB3sVWYqA/dsoUP+L7Q6yFBmenK8L0ljmcI5vZMR
pIatWZVmuNJa1X3J/eTKF+5TdaUbfeOsuu3H73ANeHqmmpl+HiBcHNjCg+QFk6iM
AeVW2nE8CJqw29N143F4DyU4MRz57eSWdUv6jCj07JMJRxkqlvQH7rK8+mSrIPyj
49cb3XDaOyput0PaXF+ugU/pNf4qlIBNCBIotwFElirbdxpeKwrD+cUvweimXwmg
p3IDI9wBOxsDtIm17s+wUSVxcGP1jIiMyu9juVLm54zK9Xg7XSdQWvzbRXp5RDTg
s4MH6Iz7QeD14n8QQc9iwBvcZf5cSgeincPm2X+ut82ZU3RAZPbgz4ahuXc91u6N
fWZJtFx1aeGMzuBbCzZRTFTOYlyEdpzkELrJy1AqJF53upceeUCZJZgP6QoIlutv
BGAwOYaGDtqxiKEjEYBDNH5k+uaAmOinTcZm5W121LYTJq1HCueB0ji6/Hg6t3Ef
ZIMZ09Ft0i8Wo3gm7eoT4whCba198I/gkAczpLdv5Ca3LvqnvLfv2/+Y/AFRziPY
zGHMlaE9V1TygB/lHEY+iTq5WXrQvJ5TI8oYhB3Q7LOiEAziDeRWPpBtrOQ/q1N0
9pFCzYHsobSkITXNpbPBYpvZbKuHanl0c5K2tjKKzxc1H/w/LSveOnW+inxQbBnz
BR7N4VwOu4vUSJg57qhX8Ysbe4Z307lOtKencUtQtQ+o7+nTSw68BrhZYr2b6mnz
PdD82D/+NM2EY95MkIW5FTbONPnu0lTT99GvBVPcRas531N97CWakkCUfMj0GaFW
/nHnM7buOAKyeWZBpenIUi9deQe1L5ZDyxr1F6pxM2ctvhgUuahJeCN0A1m1M4MQ
4uRd7wX1HcUdKdQbKXOEHsW+qLsbBBHZobOrGKV9N0B09N1+bvE8wyK9qCaN0MT3
zq9c9f9hdKRt2TK4JfOzh6BKNhHh6ijnWMKREc9+ahkQtSPuP88WHy/EqKb3eZdQ
yyf2vg9h2VD5U72vKEE7vHuZGQJMx6gACqEhQs2IgW8g6lA6yZYWwDAZ913Lik5y
mzPEkedV0ZqOhska1VIK79nFH9nr3v/kdWUAnkfqUvWMEJF5mTHPttuKFoh9Yt4/
YAGNIIqyJ+SgIzRoyTizy0ouG3CPeeK3BUc7oNd1CeaORX2T7AoYOykc1RuAjqA9
zDassuWQOHGc5ALWPma8tjX0YTPeRv2wFQUTBom22+7EXuFMYHUT6JXgtIMoLuCF
beP0+W6e0aCVtJiJV7KF5KfnugFyWb8qI3tO1DPFoY6ss71HRh/PhitzlPfMdsip
3+wAxdZoBcWmxHXCPl0L3NHRS70elZo8oXw2jFEMlvd8Ke+m1mc1Bz+okmuG5Gv/
6kv+1/jQwnbqEY/ckxC9fa6ox6w55jHd/E5pAAGQSfmbO7fhC8a+FYds7GP6nQkW
eHjtrW2qzzHd7X6v8RMZnPAwEGMsIAM7MyhQdko4DP+cO6VKXbzgtctl5VPVWCeg
gvrSnlFaizx64mbsXEZUP/Ivx3d0HWfgw+1NdVw0OqKYyTnXwg3/hefGWhU8iucQ
A40C4koUin2S1NTXurD2OrojmUKJvd7LXa7XpvBsSRZyZXeJL6XjILAxD7iStzMS
Nw/GkGFpklZiAo1YZ5djvll7pAxRu/8uAuXiML1D6H9iaM69ktpPg+dvogqIBv1/
Vh0cV5pvo83eswS7cOyvq0p5u3VUbF1jU3VyniYNKsmrfj/GXz/omjE5PLQZjxtY
TT7quzwgfYHLDhcr8RmC5jx43LXWKYkl1p/BcvXI8odRqa7SW7LOntRZBvEi0z1M
VLgWwN3vWewGmcYtf1AsOpf+FafCpYDvRFgJAyyov6OnwBYycT6mamUbuFq1mvsR
MmIktZi0Yk8z/Ynow1P7lnh0n4bZELJJS0XQFpCt2QzPBbQvGFm/8J+nD0aj2wiU
fLwF8O8S/h/2aooONoNq2CYMICNuos12yUrV406NWaOiqKTkqef69D98G7Oatvll
7bVT6D5+gGToEDouNlCjYw4C9FUc2TPqkT07FwnoQTOy/QvC0ofEqKXcDZpQwMNh
NjyAPwB2Vjb2R2w3x7a2Inx1AZW5IHwpnZHJ0xdsZAk12OwnlTSBHcMwSL4IovKm
qxbwH8kvdVEVXF6ybSK/zu4s+OppoP5yLPEyP9KF4FV//3tbX3q+D0OPzjN3s1+l
F1aYA+PCLuRp0ElxcbJ2BHSLmzYkrqi7qjWHZMk++17P2LwiP87NX/6JViiieLuq
xQYDMCK+XIAUtdEpg0OAZci5yywUwAk01YDipbzGoNbEIRzmIBYYxoSVXBJhVeZF
Tp4+3qQKcVJN9Z450fLeIoKINR9nxQ+xR312pgRpEt2NkVP649iwF55bDpUKpBxe
Rvp+/QntaMeaNMJ8gcAQpYM5XU5MZ1BWz18aEpeg0GHwW68ict8nyvTfjDGLg47c
a7euhXHl3IqTyaSxS5DqHExyJNdWpLEjxeMtCThrvvmXGBiUWTTPYx8GAhkAU4IS
/dcximF4WhPLjirN+mJEFk0HzU0jQDiSexCOhLmpuEWLL6LI4om3zpdjhJuh+Xff
99hDFMeuSzlZI14AYIYG9i8r/uOydfQfR6456vaEmNsXEl4lL+otMLRAYAO5mJZT
YsaQZfTfjLRlj5VQBOBsiONQuajr8wIsUDTSj8TkuhG2nhZpINaN7ouxdei9WGCl
NslUBQSc6L77/+wy08wMjS9VBzchZBOatRoJBkF7C/IYJeSPQzchEEtzq9XnSxYa
vulz+bjo/KbT+kVQRyXl+1sSrAW/YO5Ajf2/qoL+FFzdqanvQ7bPOR22E4e6zjb5
gjDK5eblZMSh/+BjCNjb4hVjEyax+n3tYGJQfeeB2bHR7ZjXHJ1CKH3K1gFHXwOB
okzHZArA6hYDGPUkbZKBPa+Rw/sFj93uVfIHWilrEqGCEiaEWqcePOVnKz5xaDgb
jHmumpoiiuA+TcerT8/Ev0Rt38CpFVQ3LsKmtxPyuMckVJrwq5nyd+AsJ5ALjL3k
h7X9qobO9vmyHmA0PHMMn+md5N9DcJI4+xkyfkONVIY4FCyOnb6feVCLuWRG35tr
M8uvPL+Gwh4kOzCf3GYIXVJ9VkEDBwkrO+uu17owd8CmwB8ZoSi3gxV0tNLUi1bJ
YoQpD9jRTc2hMIEKLKsLovfDNXiY1YrsbSkILoPy7+8l5mIlMTdkbS1lcE5Ziyqt
6gtQIVUiSEAj5rKEkNPZ6VGA/iuzkIAOH78SeFnuRh/CjgrnucyjylXWeNbdqnV4
d5VLAiywaSLxZggK2h1UpRTJzkOXY61MreXaBh/r+U0abmSTL9KLGMtzXpkpFOZQ
YWQNlpzScKOUEdREBBgI6Xrc83L524zBqoxLUQ0TgREr4wl3wXN5cC074GqAy855
+l9bb7vQ+qvLilqWaXsUEBHRt7gF9/7qfnxWoUrjQ4+K6/kkBC2baBCgOIrr1RHd
lD1Do9ANaDrQG8JOrX/YFNE3LHOD8s2ZsrOH86H122D4MIckfwLyQ7++wjxnVr9o
QkHFhuUJTcGZslukA/9GEugAgRldcxDGZyNnk/eyGfgS5sHLKEXhX2Q2sqDkKmLu
b4IjpVsJmprM+yMy4ZY0VRkUGGyN5DYGddQOp+lyzJZwLlAajscTXWFYnWao4waz
nASp0LSO3r6xj8hnNQzDZ9j0aXOv+0bmfazbAfYFmWbQOS0N3Z3dF5nDY0EcnZ6E
OdXbIGQbIlVFsoURIZT5vbqvGVsL/kJF5Rl5y6pUM9hty/3K6CB61dWYh0HAvozZ
lzm38Z1GbvJL8psx7SvOU5veVCIJLHj4zPAYMoKsrRqXGZwp+zc1h0S0rPIAqAID
B/jDMjEtMV9184ziQDRwZ1kv3Tuis5GCNT14gKAOmcG2/8pKQzhBPKG/Znzn6tUF
9UskxgkgyaEUQd4R6nbfSRszo8loPFObm1DlmgWpyMykusfdlpTXqOw8Pnu34cV4
ftazwYWna1xjxe352IAau3CQKTviIJRl22bNFEEwSDlmT82yAgFiVDhg5k7DgNaY
8QN3MPUNXyviFH7AkWuShXz67CYVr/bcl0336HEDDP/MaYgrjeA9E3LuVcFguadB
mbsDoI77GyQjHEckVaVwfeo/6IBNGgD2CynKJbNrVLWrA2yKVjg/AaatZmhqbKGG
WRrz+tgldvqOmVSE8iDLEiiDilaPq7XBTiNityt66zw5DjLuJlBlNSHsLXnK6Dhw
Ru1nB0JxvSjipe96XDKy6OqrRkfOSz6gme2OBT0RSnmlIiyrNTM3ahvBMdgzPek/
fPDI3Z9l/uSQygEDqAsG5Q6znIaiYZymJ1nJC/3kIz1Qm/cbO8Hr6NsR54vZrgbl
6tkg0ub494fRpHBqyqUGA3m5HqqRzqgoITQy0les//pto5qJlDWzjwNw58s6+aBP
EHqx0Dy3rqH06CDjr8K/Hf1TeDaGRb411KJk1eDuQgjh35wUxBiuPkgjJrqim1LU
5fahBQov/KB7YtQ591FpohbgZqBqPAQnQIGQHksb2AfOzcHGkSPN1GPIUljhEXDk
9J0wVKywIrQjJkRL4GkExlglmeH2SJ2RaGXT1P3JFlHRjXGFIMxiOJeTGCNv1hBk
zqOQq43Ed3gYpUvJZOJYaq4B/CUJ+zxtxkOyzY5nwb6sNPEGNb9Z9y9AmEZ1ViC1
UUg7tS+yPhYts3PJhVNP+KYQjuKUjq5OxNCStaex+SzbCKm+c7aRKDALXVruz/br
L2gznaR4jYC7O3xI4PojFBumaWpnzeCd4WV335YM92bd9j5urfmnoz3+9ptBDsQs
Z2ys9D6VcdD3lDekrGjV0cYNo6nLLm5ecIfRhZLKwF0CJRL5/BRQvAq/+5BKslWs
PvBHrmCRd4hmWRY51Mjih29eGa3sfOnIoB6H5ynTO+Wm+xDr+WvWa5f9RUbxpIU2
Gt53NfUfKmEPoX4tzzcepTnLgbOXmWsVSPcODM3+EgK3YxYOJ4mz0EpwxIzd2ny/
bSoWmkdjV5AGle1SOI/Y9NGeff+Q2WanFhpgczjknHGFdo7EC9x71kEJCYwR6sBJ
IiGr5UlZXf0ZejpniN3tc3m4S14eIgZs5L4AhSFTvT5vjRPanHWwkdf6SE4NWqwA
eJZA6CKoFVCFaS1rgTkvTYKB+3ZpYTGn0Zdarw26j7GRzqixoANThjeOakW35PDd
2yS6PfUCUGbcQuaxUkhiGXGv1o/wtoY7BolV4JPamHK6TlSz1afIpuxvjCpkTHvF
gfFf7iB/QbGUyDQAJvdJBRqJYT5tL1sCZP09O4MoajHYnmX5S2by4NivNy0QWcXE
OuxdWuAdA8dzoisE5iEzPShEDVCuUh3TNXS8x9rTn8mNCdOuUX3YssJekRX4v/Gz
BzAtKvWRhffa3B2R26dl29m1c6tesRtkCTnkAM9Kq0RnPUg8JwJrxE2JjuowVVGH
/oCAv/9li0LPcD0YWZt1T+CSfhbWufjNzpx3LPrNYPdN5Jb9UcjivslFOcDte4Y4
A5kemmMASvDNGaxdn9lK7uSxhjjrccV40la7J5sB0BFvYle0821qJnLXNjyBwCkm
CIM8gmUT4t3Rv6mQAK5AarUgCB1FtKA13RLtGCCl7QAW6WtXboouvoLPGiBcGwyB
Yr+jACxh7ALuD/w0fWaVmaoUvgeM0R+wExOf1WEIf2eEpOrhSL/Qm/ims5XBGDk4
IZn9in0vER5R94sel0IhJ4TioVbnF5eHQDGdtcEZgfGxK/nUrcEvW/6Y8aFfpvNs
LXCum/t+Mrq7XkQF0ihH7M5Z7juuaeuCggMJNvenjIqd78HvoRpXAExadumf5zId
TnsHvaeiCGOO5K8vj/Oi0FeX4wq/ujNRdcTaUmGK8X110AGjrNnJ1l73Wyu+cYMz
ehwmbhrfqeSPUo8I3CUsfJ7RgQE1bDtPMxbIgxnpX9rZy7/9dCEGWP4RbfQXXhq/
a/arZAx4to6zWVd3gCEzn6BbFg+eU1pDThscPSMnongpCXiZ4Fl67ox121M0XW9G
NDYiDghYIEcqyms8FWjHWcOVr1SiiESSlKrDZNYnkU3t1Omph/a3/z6/pcw0gsxr
eQ/vJUzU2SZwa4pKwtHHjPpFaB8zDL2DloLmXldDundH1WwWk6vQiqwDXUxeCKoi
qRhyrJXPPSXoPMrxinzR2K0xDQ400jWBKgrb/H7noFGySMUOtTR4krJkHWkCHvjC
Z1ExK+PM69gKulywZ9dpqvOxdxw2/rnGM8AwT+JhynblmOXWJRDrbsgQM1uNJQ1w
5NpgG0Gvdjo6MZKnjqRHuEAqHtHdXsoQitrfsEp6AaNVYMBFrsywOcHL6qBv1GUf
d7ZDgr1p3XFN7GBuhl4B2gVYwu5pmmLJavM/1kxFb7fP5nY+qflPkWk98ItJ1xAt
WccX7C3c2eJ4k2ovyia71TRQvmPFjT/5CWC3UhpW7C1vAIf+1ICDAh7Zg+k1G836
RHMfhHHYSkxU69YCAWXOfmiuqY9BDNVkzQ0TsLkO+Gz+gvlg2HYqwyeNw9pskDV8
AQximVLb/HmTh5plQzZ2hR+wL7jMv8Odi1U+TjwvNJvl58tgSzMqB49yggYaDkJq
1drOhtHBHYR/saq86rKeBCICoetJbxeOzN22d9Nv9wtXdPDQTWlb/ZgRkGdGZCxs
iFdHpmXImw7ci9nf++eYSxCtuXfP+OrB1dmwbC0Q2JbQ1kJ7mrtB9jLH8FnXzspO
oXhUKr8jCprinnhVBNVaC/Jqnr43PPhnwFCCxfv3TEQxOetLukQdOUzQ8gE0RLho
dZvBRoM6OVXH9KO/lOQ6ifYeto2wv7EHUZEVfpAbDHF48Qi1exsnTjdXIrIbWbje
X2ET+xjfPyEj4bDXGjmHDbNT10IoECPZF5WnLkBrm1vMPReJWhBW+liH17XrtzlG
ahlSM6ebim3yY4xa+DV/NWmaO8ZmluLBNYuEfrBGkxVEfKko+x9Eibqpyj8m1QvR
jh1IDRjd1gfH1Mgy9+jTtpuimgqmAAGu3rg4ajsllUgwqF6BhlncB5lZHQVcUncE
F5FbL1iR0dMsVoh+qBQ6kWB1qdjugkAklnJP64i4Hjs6x9MrPC8QlYtgfmPI1zdH
pPtNUaoyS+WXwqRJIhi4l/9ZzA9A4t8uXkEIvkYrsjjFUK0rIh5XjwjhUUtRF3xo
GPzKbAsGkLZsYVn+JDmQKgb4ZnfGSxDT9RknjUplb7ptuK5qSg7SQAG2NTr4F/Jq
iwSdSrU4LEDaSYIiSdAaXsoaGAWyL5tfzEbqZj6M2JWHvnC7OR3ki+nxNGVs5yU0
03bPaayqJZyyn9ZsglWUmQL9FSlj0K+Cm43WNdyxvmNSkwxO+g3Bd0PbJfZ/akir
ffzRbrXYkvPR7VnJnqU90bq8K0VCVlaqJK1GoAXiyR25fvJ5RZSyXAUkxyxYJLXP
i2mFWaHoYQW9GscX/uj/jzipFTFWxTzUSW+biGyJApo47Ih5IcUIiBIcNo/vvCWt
hzEkeHSj15qgbpEbcgZF62HiarjDRyeU4gQ3ysTPPW0MAo7XiNwFDbuI4+HO76Ph
VXC1MiP+Sa5AVnypnNEgaDGCo1mUc1SdHfJVsugiQTttckZSPSObUUdyTYHycAUA
40Vg0QhwatYg3nsyR9/LQgWcshHnlPkh4/5Vo9DN66WiE2KRhyzQTfuOZds0lsgz
3Lj2uBvo26JsCPwloiy0+p3JvfzAowQswGEOAPdGiq0YjizmNlGmxc+0gBNmyrwz
zjvy33bd+BCjfQ0MTHUlPmYbW1PHnzlatUkGC3Sy15KN0y+NHXV9/TUF9gTL9lVx
sofguLSClVsQmjC6Ngad9hCzkdnHPeOounsmeBE0pAbApis3V4jJ5jlJlT15cLsK
LoT3xgmGKnoI/DIChtgyhlu6621/bU+Z6LYiIB7Hl4TQFd+QzfgVOwlpV5mghzzW
MJoEgzkgQWmFnnfEO0pDUJK4H1L/2lHZ/6IF9Vi0uWzp5tp/O6gS1FMKLidQV0C8
F9wRwBCk83kSqkGBrrURoU2Z8fdaH1c4lj3quHAJMKmG8xiAjsZZkCAED776gwuT
GF7kIPbl06gw1+OAkciKHPyoByDyThK9sYmz1+GjSuPDFy7083T3Q4ixvED5HbpG
KP1BN1rhBhlQa3n92tUUjuw8EOw+uDm7Cansi3dGvgxGzUcNk0hdOJZyiSleNsvK
hqORFbMpbDanVA/asRnQKb45h9v9Ivd7HXMjIJDmeMxA9gb8S86aEtEjK0/PMbt+
gmDQXi4y+TQnOyVisQoQJ/2Q8FOlc/aBs+U9Kz/+Hux7gek/Bmc8jZLBSOFMNKL+
TJ+XQWsNwrgpULHKOXuCrzPmsy6SZrEl7KMGAK8tNxYpdu9cFRdHFB+G5g1/8bZD
zH3sXZRyHmGmEBFNc7L3JiIIWwtzczoccY9zlomvsj8KzEhntErDmwfhIIiSha3s
BltgbZlDEKxMrZdNgCjTXJ4kQwAfKtWEWWYtdJz31BY8NVpH3Bd3Tyxl+FMYFBpF
XM/C+o5TzoDtkbyVmau9FTRgd1fnQVxstBChhXFZdwYJ5Ze5uLhUl2fH2xtUC0gq
Hg7fFw1700YvY3BnmN/9tVVgqeeLD0+oIAZCGW0c8kcKQG4o/76i634a1Eh6Wr9E
gHWWFj6nd7BJcgfGJTChQXeeFORux2hkjwFLS7YdDxXPyU6S215p76DZIyTi6RVx
rKigJHAP31aZhAiNk01032/iKBSJMpTEh3UCDU46K0oAXaSNJXtUrFJy7mSccmYS
aFia+eGrwQeN39dh7nVl4MbzJUTnSL0uMX0ofl89Wi87P+1mv/7DLTUepnTXMajQ
Do6cqbaIEs8aj0tts0L6k6wRo5uYiyLoC0LCp6oO5AVtdH0g8JbInxxMhwkrTha1
gYUxkxhCO7efOpbkS3EEkLV/EycpM42kVy1Dm1beNEhBlBhYwo8JkFNZNjd3w9HE
WXXdU5ZOZntOQvarKNizhv4KtWCqoX/RhW52Ss7QGpfeDuiUh2tT+EGgn5yPOFqb
wnukJBRvvAe/v1kk5jvA2KR6Lkt4wywc4P/5sHy7Q4qD1m14p9aRmvK+AINYWo2S
41hHs/JUnmOHQGM35p4310aUJaxtIExDSMQPK1vqzlV2M1Dqd+F4zl4pQGCeLh1X
WZtApaqrtcpOMHjoQqhgxfSMW96rPLc0fJbSerIlZKr7tHFp9LnykZpVaFhM9iD7
CD01Awfytgnn2PLzNL+73pt09oVR8jyJG5EvOEwaJ5evQUZnw0hVjOWZ8crjUQSm
X3+YBDsn1gAsQdXvnNboAmFv9OyTnu2BpndyNLimUGUzNGj2hnBXYxq11DWnApwp
dxyp5GjfleX7EINZC2u268TgXFQYSGqEP6+puQpKSs3xSBQ+HUmKU5dzmUlrfjTN
ofKaTcn3pHw95XtA6jrXRyBlyKxKcGdxD00tQ/5VOpQAjujguFufFtsFSv6enHrD
3Bj3cMGIOfOdlcApzbpc2CDaf8R90Ssy5MRz4SO6+xFPhjxw8iwoqOLpBXDEiyKf
Pd478zf0KYmzjY0Zvcw9V2vivCtot1VMT66/heyLhdQwiQ4Zv0Ay8uestaG+xN8c
I95XiCvA6rRWG7ROFU742YDapWGuXJN03WpgbMYcqxXfTJLIUn5qegoLWTJhijr9
IzT60EZwhK8/JtoAHNKX9wTMYvGkwjVo40ZBROqenoFwgJCe12DUcjibp7wiM5x4
KIrpQIzlKfeK9Y3rL9bJhMUeJvYHtOvZAf8uVhC57XBU9JkCQiZnCk5y1pnCMpnO
vu0e3y0U/dhQOfFX9atPRTtXxbG7idw3kJtYiKjHKy5EQD1pZo1mQR0RfyV0Mqif
YuYRb3cATQXMS2bHoQl34xVn2FLYDfkWwQxY8EhcfcdYHLQd08ua74QAJZxGgug9
45SJI/YX4IdLwXhVnQH0+Vqu3KlUKnR1/bYhgwqjHHe4ZcUeend1MGdmbdMU5TVS
I5qtnTx09DY89bYPzyrSGzCpp2MBFgOU+r14diN4coCCEam6JDiDpXvQLSnAnK1p
AFv5nshtdm9dgi1XuDk6bqd7Let26CgNaC8Ekt5WXPI4SuyTI/j8ae4m38gEcHpl
WU307A8eJt/IDowtrcS5qO3Que7iH8V2vvokqZ8E4tYPmD9rZ8x3lMGx9t6REER+
5uR8eNZlw9rh+UJyTItWRZrdmW/Svq1n1fv+IvcJ63lUMm6eAUEj2MWrUoWUqGgv
LYpFJ1LfEJrGmj1PG3q39/sfqx7vwdYYS4DY4zUferi5BI2FD0jm+AbdnrfOqjv5
odE+tbEhfgTH0Jx67/4n5LWTfKUNFLNk4azi6dtkPRhpBSD6TWIhjkPeU2EeXKnl
5JC90mpSwtGXlPGZuW1ZR5wYpnjcgIuFCV3NhzLMSO8zc+0hwDzLNaXCN6Tl0c9v
KpBH4gbM6tSw/8wAWgM5wHIZgT2dc4NndiwRvy0fwFoZRmPrWQrdD41Sqv7SufDc
60MTjEv05owBVPZLolnje/aBeiq6g/4/MiSgLrJkJEZ6HAUWtVmEncJgg5rzXluZ
4CVDC1JJpI5i/L0oSDiMUFO2CnHPBnY1CvtXd7hsP8o2YPKrA6x0jb9LeonofhO9
nMr0Ozux7DAUMLY6qx+Z5CPeGDHrnwppv93F8f8GT6wA5PpvK8kRcZruzQesNGLY
RvH06dYewePiRYwoZnFJvoaKaCN77cfdh0/I28KIQr3uAhqXIIGnQjsq/SzMCeCL
H5FFL1SFphcHW8SrAk/L2Cb+dNUtd+JqwUUMgoSfzJBvlYINfKGonM5EB20WXGzI
+Dh98An74e3TETKT16yGF59jcVRHxOz8VTAZN3Bn9/LKjYgDHqsBcboFMrtaVVRF
X41mp758E0bd8ty4gjhlMOOizRD04A+M54kOu3skG/JVtyHHD/iwKKhkRoQ98hZu
WF4CuaA7A11eZgD65ktDd599wNqIMpaKYl+lnr40jL8cGEz4whGskkpFhtJUFJgb
jeu+WWY61GYnMTl4scAXQ1jyu/gZvXzbm08kS0BlZHgNJcCvgSmiMQ/svPzWbKf0
qH5Qj+prOv0OdldjTfwlxY67xVR5OccFW72YeJJDAGM/f2M4WikNIBjawXMQ8jPp
PpOR9Xg7wHMd1toWFIjLDFm3nCa9C8r6iu0qt4AcI9nhiInZOnZKqECa0qaGb3HH
At4ibgDkv+uXh9s39SxeLvE4O7lKIkaq+BhJaZ0AVK9FVS9g+cLCpPQ+6Fcpf+4e
dcf9wieMftYCUO+OwatJQO+DWFMPBdcytgKGYnct6eKgNdfy4ZCUOAOTRnfpucCH
gmn2JN59Q8zl/JxZ8UI+ePFBz/qZwEC2gPPDSj1/psq4GpHzfwAqsCK22LexoLHq
8moT3OCq8OqMhV5PrltDV2b7SK4QwpVX7czpoaKO27yAGMU+LkdQLv4tDwjQeC+6
Qmn8Fnx8UYV6DEu74pR2JTjK21xUdK2PdOSxfGJLZDBTFj1ElhivqK0eXuWEjYAz
6t7cbvJx8YksqDXOupmDu2RfXnbmsROv3OJEYxL3idHHVEOKigM0iwrBrRfC0ghj
NJG9zgj5FkwNQh9o2GgtMqWzJlMvtiaHl2rcNyOymIEvhWzElNN0ZlTJ4799Rp82
uSATFOO0XFMH6glbmJ7CXhhJfxvEMSR6C7wdV40CeySMqPnIWpT16losqPZcFAsx
VjcmSjl5rYsZ8A+12zrJUviwmgJTA6nuYw/UKawowEgqFpEwNVUwgDPJw63CEDuj
FQFZe8XGezN7dj5owjiVAMzGvBZVYzWrsUYPiobYjEfDXOTfp7WC2BFHLS/8DB7u
TRAgcai+pynZhM8B2ctaUU2yJ9YYsPq11p9w3OBuhIKnQ8ymCFa6zM+pILXmmNpM
ZRT1dUce8eR1xLPZHP8wJEOFNVweBfP3iFd1v/fLvmNhdmecPeYRCBt+kqtYKJRL
9TEV13mX9Uio2+avYOnOTGgD4VzmUkGnnxAbdY4sUPS8j/VOKhZp/UUBOYLzYe0S
wX3hCDoGBI1q8PNrZgwPYdYXEJRjNNgsYN16g+ZWMmfXYrtKV1cvxaJncaP4eAHt
0465r4XmXsjsaFETWnmCO17cBBDaoG2dQ2b/KHQn+X9aHaL+9bI1yXK0eC0q1mpd
/Hd3wSb4HMioD2hVdVGgfprwDmYAOT0aYQC+w3VbSAlhim9zL0QQ/tx9quwHvbGN
ON9FPqEUHQCZIVDtRohBOZQZ4OHiCii9rMLtVJE+gxlT2xkGMu/eSD5gyjejL+Qz
Xj/KW+/Bpz5g3fOeOG8o0ZqjtBIOvqELpCAK2CmrYVxwlbZpgqF2b3xxh1aONLP6
jx2U1IgDiLFRPDDwFFG5xtKIBj388GKPKnVTSa8TL/BsBFpxfVVqqazmAeVHyfdA
bZ9F+uwzVAMI+yXWl8KXJh48KI0e2CWgcbRDyWXD2MzUHx7qy1lpEUi6NF/is2Pl
VzvPghF3mR55qWPs7SMtV/WJ5M+vHH/Z1f3ozop6Ye5YdVc3pWoL82QLcfHcZHDu
NGkKrHgTvZhHQoyEIqfcQgsw26EnNsna3AkrNi/ca0isrz/5l6mz5RJvSsmxpZxt
hRfrujMjBM3N5FfDhkC8Gtfbn+PblTKYDV9HVu0JfLph9rpLzaNBOhzTjgNBS/en
gi4e+zOYTjNydGEqG0QIvlWSyUs4dZsZxptyNQBSJ3F18MkxQmebCAXQ2RCtQf1S
/Uwhn1XmQlml89Vs1Ip78+swUgyI5PNHRBh/Mxmw6zqOvMMtSIksRGI3AEu5WtXt
P6nPOBiTA9P1QNc/QTAWVQixDt2oVXQJdO0ea9Fef4C9eHQrcd8S1KuJgKfo9H2/
BUDZvKZFv2xybp0w5SqvH7lGsOSazSFmDELN2CmSGprWjOCcOVHG1DbviLrpFzLr
ZRJgc+an+UD86fBpJKJDXb6Lgj1xg2dZ66P1f2N6UEVOW7P7u1A0WciL3fjagnHH
7jU8riT0AE6QEJVlehgdSLQmiC3d5Cj8C/89pMMPKTVRYR4+CjFnw65yWJ+w0QdP
z2HH+2+4XGtM6OKxBer+LSlKfgVnW1ZxiCX+tsVocIeEep+XxOcQjpWiqjVQQs/e
PSSAYugXaM8bpVGxLAdWpRVte/kOQ2B7jip63LHEJCfphVuUvjAulZlT8hgEotzq
4qLgqjgHdTvBU6aL/i9VO6uiki+MIsWWaCRrCckrYNt8/4+VjSEd6S5vUlt+MhTA
F/5igQJhJiA/KGZtZWlLO+vg6TR+08SuuhxzvQzM9AOKifcAQFmky8NNF/M96jfA
pYgKPVX91nd3iXpTiQpet/jxM9Zz2emquwpc9R1coci7sAaN63k74VJDi0Hrb7j7
x4FgnFGomnPZ/awHCyVLBzb73ZPqxolEX2r+tvk/FpNvjyjdikgoMQPUp4aQ+E+E
4/oRLr0HiIZXeCALXyQHK4klst56Tz8IlRKxP37a9P+gK4iFMHGgVb03PM9APNy+
HXGOsgpcsYEL2a5I2Kvn5kCKYM15RQWM27P7jHQ/W3f/35k/ESRB+j0cBGR+zgTa
Ed7ixaMXHg/hy3HfuJMbWIbXK+fFvcFb5RfK9gLG9j15Fu2fFnB9BWFbspQSBkCj
DGx5cs/umK1groToOyHjuB17ByS41azqqG1SOpJBubfCQlv8O0jaZIJbbMTdAiqg
m1YQzl/6MoPHrKobhLtp0Ujx3S5xevIJV5JJDs9sx5l22SV0xNPJmHIrJrlqJwMD
OScy+ll0/ME3qn0jlQFC+cwBnyayTwbEEX6erEpMlib6hl6JAiZII6DJ7wVXGwu7
ke063Na4e0GnMl6QifjPWo2dwoJQMYi++YDzfX9RVes3dzUZflVIBAVeLCjnGSTp
5AbAHqE1r2CasM+sUVved1EHz1WC/4DpL+NM4Olic6zhykruKWauVb3Dz0fn4HqT
jzvOJdgOov8WIaHFyTtLu9filGnDNbl4dB7pOANgHvhY/gYO5ppgEQe+KGwhsXnK
JGP0RvPaQiBSSSv1KQXQHgGhvoTgtWvXN+WQJa4HpzEhe95wHQaPE81duiIowGCx
OOMqxtp3EzGaO39xxf5XDFBYOQ/xO2RfqOIM+arMfY21TpKBAMYpj/6W/xvPCteZ
5iI5B/aO+wxG1D1qtFREzXkXWHqTGL6Gjb22yFbXESwgSbPOALCkwUEiWcYyUJQc
y000OXiw6TreTZa4jJQ9Xvl77ctPlRZq23GD7LGabomUcxAPoKRfKp4cCidJpqYY
q3769CLzoXBmru0bJThw1KsHl2iCej+KP4JaR9xcJr5HAqKdZN2flEQBsQ4mH8DE
njtSkM+TJzPaXDx3wmLSo2+IADoub3WF6Shk+a74dYkgLeIzbDVaIWIbOQewteZT
k0hyzsxlBwXBDFbr5QFZQs2IA65k5xuqUGRBJOGKD1sqLCkYz+u6Yp0kLjxWULfi
86pF2mrIP3fuPB8FeaYqcJjKwHZD7bjD34i9JlEk6+4VG4mB8KK03feGFkd4j1tT
u0DDoT5d0k1VHjVroBpE+vvPVyQnbfPQv+vNS7L4dmV8MHgXbicIgbEJLMWqoPW0
2yEtP/KaPxmMgDzP0ZPLS+ru1rdiF/N002tev5GsrsodsIQNxsI44QB9abIUEAsq
gLN90WHwtslwnE9dF4eLsIMRjydJR2/os4Wd+9Li1o/KHfno2BQis2JZDIi3CVEA
Dp69bnbYsfFd51Qu9AXZjnfOzYoACZtUwhsOz27VeTc8XEtilkVQIQ0pqNeaCF3s
MdrDW3HCDG9ZTxXy+R4wtPeCWpnbPl61ZXPy895KFnKKxfUDoHIYm+1JQa2SoQID
XJy+UNd/hCmFHaQc5f2D6AM5MgFB5FCzj4qzwkYh6wO00bgm5lJEw6qCGxMElSb1
Qw1uPh2u2olxNdPYpXol1NLFRQCNtmLemmFejuQ4NJfH85KaB//3SdT9jMx4XRU3
H9/oJl0v6z3cw1kyPGtQFd+fBTijd+bGv2w7Vqro457fZEP/JK99TCBwOupCpCiU
f+FG3U9BvfetHdQ0ykLAfXlpAT0cJocz/Zy7M/5Kd+Cs2Wf2sg/y4vdu2WpUMxUy
7G5WFazK9zRxhWXuUhEXSkbbwLvrQWW3jZmIbCbHEAZi3DkBe4JNsIpLnxIY6/kq
I/DU8E+2Lca/Ee5gJGCwGIjh3ZFCKXJfQNRFM4TKwx7BN5I2tYX6p4mEToXCypET
Rd3pHWhuJKGpKZH+3/8YFPAcK+7vGsD7Uwy7zSXEarUL1FBw6MsIY7RYKEmHyXEM
zv1OAPw7QARtzMMchorQkBiXQ9ZJtGLTg20daB7wm2SLtSn1CQAxfkOVX1ds8LtB
Sreft50HALYs12kHeCx6NGAaUuOGxOVGQ5SMjlekCdFm2Clhj/i3BCuagQkv548F
IlY1H3cN2ze4h6aWrs/LJDkh2806n+HzkemRoamOqcfH40hCsIJINq8oIjJe6l9P
ijgt7xPwOAAnznJ4tvkp/BUZtcEt2ai4pcYB7e2kOXDbQVLZ9JodgLvWeKt4N7NX
TmgtaM2RXWVt4Xyo0e0crwa8zatrNoFao5jkDV9J7W5GVBdjYwO8vAY1uFTFCOpn
Bj604iAYzLAbWh9z1CEJ7S/+s/4ntsN1Y1y2KlIalvMFzVZvsOAjLBQo1US4WJFC
XGvcxnsDllLvwsR3JLZ4P8H2rMqdW73R//d1FSPg6StlDqR/JPTuMSWSTq12O5sz
pjPI7aJuG2qJWw3nzC2Aj75p17UZ7RZZKAeloowT3hHyEx9eVVkSdTxSaH0elU2R
V1GRpIPVHkvvee1x75QzFM1+lh15mjVOkuuXPDJKTm1q/Nn0cTZLm8d0Dt979RZB
4mfIXtltdVpKPBGYvUEsQJh6y8KEFNnHnn1mguvfYld3tYIyvNkfKxdQgB8o4lmY
r4qHF/OoVlzo9Dr9xaKRQwAZuSgR3NtG7ArhrIm5wpc87rHs1jSxBrWl+ow72cTP
UUP4jSMDKov+Xvwi1/bcpJC5dw8H8K8jWoR511uiWDpKB3yAB/fcPPSyJwer97uB
R+B8kJ8qJ+ujnxs6uhyF9H5MPKlNP2pE/KsRmtVn36VqnF/l5YIqNJAlcui6QI8j
Hh3GPnsxEqL0tXYz/QOuiAGxZI/JiR/VAP2aUT+lBtVdd/1s2JKdyzqfpxruwib3
pUEL23y0mMPWS+Xi3jhkKHBtQrkxsjEBHmenEku3kBMUChnlt+R8YZxe+WUN0O0K
3sL/YSw+2Pkv7g2j4R9aOcu7g90kIfvVGhcQ7an9Ah4FaopVftifath5tMpGlaEB
p5ufIR+4KYjSLEBrC9xQa6DILhMPiMXKNYPTEG7pDrBVQ3qkQsY0a5ULDqx3JoY0
rx0yOAKwlQ1BrEutUPR8fIydp+KGkCi3V2M4ImieC/ukCqk72cKxwpSNO7ZfR2Md
73AlT1GJ9cs8dXj40xHe3Q1VMz7qrHMQs/jrS6NM54PtkIHTzxCVz9FkjZkDs9Uc
ealtsQM9G5ahZSB34HEAIwzj/KYwBbExfTx58f8BcohcAVhKCdtP7CDZZgzRTkLd
w1uOr8Yo3UplpYQscvqvQqgFHaNTq7nBdsiM6gSSP77CCi/dlf8GwEagamsO56ny
57VFZJe5mQjpklrgcv6AOI4S/mqRMNS5J4Dbedr6qQd8ThXIeH9BeUG9FzJ6d/a6
C/qGV8acPpe+agUQ8PMHEYKPAj7TaG8KuFFK1MkMUlVGnqCgdUWNUwwS7eAQfUkl
M432KFrLGTdteaLEW0UKsH3zWCKIOOnZXFM8cqZs8fR6CVWfuICMB4tvImRt5WpY
LlX7MWfqPCMGSxdLGNfWnbMgRV2X5qB577dXB3l4xrrD4lhvzE2k/vhQ3R78SlL5
paYX2W2OrnTCygG4Q6Qymiz9WheoEiQ7yjLMo85O9vbNj6kinClbL1TiroayeiMd
qy+wZogiF3tRK6hFGmaPShGT0TW1D1xHqCowp2ouCS5u1MbzMFnbjQEFUerlqiu4
lp5XW1FMYaAgwEYVADQYasWohTJwCbVPU9xSNcrbYGhTCZWKUTPr7Ay5+n0zWwII
62M24ahFiL1wh0qRmIv/gERewnsBBv1RDIBnwlxpmuGXsZoPosY96H89d5MiTfcU
3Hb5yWGkPTE2wq5R3OXDSIEWgCFeoh9oEfk4OURWr6t7QyiQ4BnH8YOwuJak7Z58
tztBXfn2IruAAXQULtKHFDbLdOH5dnj4RbDPsL1va0azSZysEY2iAg7UftD5QSOJ
82qrDS7j2EQvMD2U1AEjWfYUrl9NYIW5soPaiH4xMko3/CnwOwYuUzUaRSNiBJZN
3QW40zEf9EdMdpK3VczrgPXODm8EFUkXKt8cY2CKyR622AlzvHXFZ3QGCTXhoPlc
fbaBGx/JozFg89AjKbyvzM7O4OB/lrYuThmWGgZf+hHsXDkn7ktuCnyzeCB+WzxX
EuAIGDsQPKN9HQTutDPQO+obsVtELDIOciP17+GTzxMAVnYUW9Ks1Okp6ZLP0CFg
s02Eq0twWD4Jg7j1pBX1B9hNEH41ndamx71Ioz5S8YQBRestN0xt5U/HbLcyD8cx
RzkXvAjOIqJIcQ2X7hTqfLYYT7chTLqMOAci63S2i+mERG/fjv/uRTKvOkgRL6Gq
/fFNtJ32UpRBEiSjNduK8oBnSKGYdwwiK+L3oXYLAnXvb6PLS8oewyir82ENA13h
hXmWhZ0IPrMAqBgqOg3qG7KNH+2zQYnhRWFWSpniMg7KiZvwPe76llSGRyw0/U8Y
f19iDi0X9IdBxJ7IZdcc25XsL9NjYWwbQHrsKGE+i9Our9iH7rUbqTkGiZQ3/XDl
OPzPL+4XT249LOLC/LeH/ycaL19CVFnKx6brg8Z5W4hS01iIGlAeU4ZY93se7g0K
ljgwXAzU/5FTHR1IwaNS94pjog0pavBRpa5elwH7u8T25hiNIlzudsH7AIdiDsGU
fCQPejgAKPUBUwMVpI2cSlKxU/vJZhwEZuJTXTYJTqpqmrHUTzFT8WZ3HoCajAng
oc7nxq8Qixl0BynAvVpFL1SyJJRZeG5dh1Aoi7u2MFsSy7OV9g2MvIXSCfsdzvSb
jfO1Byi5VB8hRXSr4DCE/wfSIrb8NfCmIXJZseb6fII9bxsCTssND5Ub48kku89+
nfuqacHdCDC5xRMRqCc1J7uMMRBOMmTeL1BJVedyKlp5DMKp5hNAvqoi8eZTWAbW
9WKH4la8ICCyLWhPs2iSB1r2dDwUgboocNbqc34cShEiyptKeL/1thuVF7aeL67o
y4NLr4T1hPZbQmLTp1AO/8O4UmgpQzc+7CXIvqwHBKlxozZw91h7cBJgyGXaYbuv
MnbJGCyVYH3LDkUJ/aKHqd/oyy/iFZgmIn4UEbDsh6cGus4COf39+UWEPlbxMwKN
cHwQDZE2llH6niCmcQq7Br/3p2L/5qOcyHBomAnAQbIBVQku7PPMBwMsLqQulN4l
iQRkOeMH7CGhakZkXreXJVQjiq7SMWNKfn+vWz4rtTL8k+TM6x5tp9uLGgIot+/H
zk01oUxpsT0L6sRc7VnW/FqxohUQQ23o5Dx3Au7zFC39qHB3aXW6BhCRYgsYFDVW
rU+n/hsWKcd4Tfi2ws9/B2okqixkRQUPIQTQzC4msAoBHFON7aazJsOJTzQ+FOAK
DRq92a/Bl2nfD6nFs8Kb0PurxCL19x9Gbh0Ep2XG0wxIYFGlD2a9T24wcYtvaips
Y0yZ5ArU2TmVdhj2m76SiithzwnWkczrrM7uNHHelTFp+6p0H7hvmqqldXFhnEyN
YjhHvbSh0BELTy4/fNjycORvJBr2z0o78L9nDqMRl6Msm0qET7ZWaZrqh/S5ht4b
cnH1SEgUaIaBYlB2UTFtR756dAZGBR024i0LUq2dVAdWIG1RoRAKEBgHrRdU5dNm
1ghj7Pu7k5CWPnc9ducv/8nkpaQzZVf6XhSXg39DKQcuW/w2J0teOfoclWI5OoGl
oSp21/72Op1e00K5hMV0YXjU/zcKC8YINpN3JJFCCuz3a3RaDFnAwSOpDMfNVBoA
ala2IMas8J4Es9PaEVoI7xzQeizfay5Wn3GyhpO9/rzQ4SrDmIka3Pft1EAtYmO+
LEJ0CfWjUqmrb9/02YCNZbAxBKQ4KfJjxfkYEh8Nt4FmCHe+e1iHss48PJUdwC4m
i+0KjZfjFAHv6Vwjni1XdbgTOonVQU93WYiNg2ZDFa0VPnd56SB5KpKkBG928xwT
H4LKazixDca1WLXRUwP/Bx0SABD+0vvqhq0UIFewZjTbSzRSKnm14Ncp+jHI5Mm1
c8oEzr1GJREesG/2ioKMse6Bzmpi79hMy4gnHu1bO8O3zQWNQcsnKoyCOB/qjVr/
xO9bxWamDgyqrDQtx5cRGuEzz/2Bi0S0loBAckkWe2OLo8LYBJOQ7T9JCkwg32Tk
uL4GojBZ8LAmKdm7yZjoL5+4FmkK2GzEtKZGG4mtv7sZb7vG0qUdm1hOKOqkXb/K
8N6RbbZEROGOfeakKOgvON/Icd2zCYVLtieO0oDTbQF2o9TU7Qou9sFwxAZ2T0+J
v2VKsaMnuGsiC97oWkhteIDDmJLpnZQPSB7JPl4+IaGQ4Tg/XEuRcTgJ2R+NQxqi
AzUW6Lrjncgt1MjPNlr7ImZkao2MVBrqyKUQYp07ldcgGBUCVE1i3kl6NppSIXL4
tZRB/58ymtFRAh8p7obOOFd9P2yeTIlTPutPpLo8BZ0paYaS+KjTZPkWHM8bY+HC
TPx9duS+2hrfT2qLJ0GEgQcdWU4/6m6dSxzeR5O+lOXcCJSJBPKrVWZbVc4JpDv1
aWW5aE0HePF8xzLdtvu92FGQspU4HMOv5J4z0gjPOmNs7nk8HAxmQxcAbJ/ZIUxu
LRfZrcQLDXaNwoHJdFY2X3xi1BT7XjQqcILCIrC0kEwkdR+wNmvbccsm+7mfrLz9
0hwjz6wGqve/7EjFuzzRFwoN++AZ0Fpen+MEHoAhKLxVhCFhIAzd8xXPQ7nRyQFB
Kj9/aOeLPKKKx15TMKnNKVQxXtPp+B2Ez/3CMqQf058VCY4MTH66okNOBrRAUz1Y
l+8D5cInI9RFRSNSF/2ndcRbnIotMiaRzWc3+9JBJdz/gLOg/cXbeg82RbJC6oWH
x6mXMO6QjuwTuaxp1XoUyrJ6lyy8f8gQaHLK4d4Aflyn3ygWDemQiv95pf81h2h5
+2eo0UIw3nsn0ulLzXIJzZigQWu7fQqeBBZh2vCPLy+0S+Nmx2Sab7CzecDKMQp5
fwhKmX16WW1ESKsLn6Z8fW3h4rIABuOPNGOEyfP+ekXv15pXpJyXzVWDVfoGmGOt
oiJs3Rv3Dptf0ZeTTNvfQCGCVT3XE29dPi3XZcK3DY3jisaEnXZD2zwej1Gk6foW
xMP+6NLpb+7aTZ+ntXhO8qKePXcocBpb10+33i6i5atiPsrJyx7ataUscSmSIqoQ
uDaNTf/H6T+RmuIQq4Hf+SUCam0OeKul8/WXxCxxYxw78qXOl4w8KWvoa9Dk/A1C
eKmAMnesvHzjdl1adoAEs1qD8t1ORuLMXsqTyuXSoID3dcw5F42NemmB0w/iw9qg
pMHiv3ZS3B6gHlzJ1PeuxotTVU69+Db2RYpbqbTPN4jZN8JswyTkW4jsW4uTamHz
w9eHviUdH9VPf5VG0v5DXcOwgyXVjiqAjjpRGj0bBYl5loMM7W7yXwt6pHLYjhbX
Dq+t61AesjaWqXVAt327Gqxli1b4F1ccZF5SWIUZopd4ZAB+mm2X/wjKNHawaWUs
EmUzcTuTLuHem5gsAo8fyOJe364xwybhH7vylvbV1Y7s6AdQDXy4uyoG1LcT5DhE
JeiX2RLVjMzLNEBGbJ6TibiHofcep1T8c1xwyyBIVvPn4udvzBusf24QdQNvxbVO
9Z4En56d+zHZ53hr5NzrFXUDkAJjH9nmJWtLqLPHLSCHeJkST4MgDXu0kV0fS4yR
qPz4x8pXw/4qPrpotvPP4MFx9ULiWSEwwXAsLu0Dft9Zf9WRZ7PC9ZVEDCuHeFHY
OKYOxUbRKrZp6E7MymRMeEnBUBwihKQFYa2d098uktcnXUXwMdTANOqRGB9Qxo5R
/wAWXjy4AAjmTkzPDQtrZf8A5CvmV2yWH1Ky79jee7WrBlZVM0rq2/HozNrLOVtO
0BevtruRp3dk8H/5P9UlP+VCJYT2Rqg7KACcjOM6+KbT9CRK7l8QaA/74PWMkPFk
KRUp0OMU+p78OXAtq5oHKG/zD1I4gleSM6Oua4FoitybZY2/GPJ9MQNS16eL6syA
tNlt6hCbLOh81S1HuQXCN/8iUE+8O6A2lXNJCyAgvU2AaDizFT9q6L4PcPF2sZXN
EVErz7gEnYYn5tuyV2wkfmzcUzXD93GCyDTG+MlVCbvaD5yb7KPn7uggJN3gfopM
l/m2hrFMTC5x1tenVHQ2Qq1bsrk15J9kyeWb5kF9HOvAKaDv/awcyib9yoDRzdyw
JNAr7l2c5HxnhiH4ke2kShtKoor6uR+Vw3ifFjG4Un3U9YPow6bfZ4rkRnGdg7q/
kZp/0niKXHOIbDUoTCeSRBTHLm4z8PH8EUpyF3sjwSPDRQ69JyGS7WfGvNNig/sZ
vykETjO7bkL6+NCxCUxRmniNyNgCV2mpBhDhVothJ4dvlv2JQZTJHSwzSw/OI0Ja
dzAReEBx9M9SRgNhzuCZ7Gekrg8QI+EgA/UFSuqiF+iaDHgsTTOXbJ+wMsjCoQIp
vfiaHQBe+j2aR2E1lICLHtHbB+R+UZYV09xWCgL2PKiNWQ5mFpqKg/AwfKjJ9BWX
TZhzZHzU7xOUQ+203uQqQqcts0duVcYqMIeT6bpPwhbO3szoyvseQ8e8hFo20+RH
rWAzwKRT2WEClULDzgTqDmFQlvneeDcbdyp1T6ayxD9Xu+uq3Z+va0iEokerZYD9
94Erv1ntBqke9hhaUczN1d9reoKBWP+X5lYoXlJOnDEZHjwQhDnR1d/apTEMNVsT
Ljk+HRLakOZVkXBRNyyns/5jsjKAqtyQiaecRltzl2Gve8FVT4uX7OWZmC7ZEav6
kBwifYAzaw98vYd7khdudHSfxfuRVFoasgyZNPSditM3Oi62CQmzCHIvOT1A6EhA
xFaEwePmf4acGBGNhPNZHchWeWVJ4PUWjjpOFCdkLmbrV414QpXx0EITfY479yM0
HQG1OpXreC11+0yfwzcHR7YRwY2NQ7pyWiZvITeTeUQ+u88Ukkv3LtECojrqEwXP
nDCr31niBP124WwCqc9iA2ENR7c+P7SD6sWpbQmPpOUNcxzw0gRg2+ifJpsIgUQi
JoyY52pOVA8nqUaWlC0xlK6ku6qtCrQTqqAptI4uaq8do0QypaUfNUyXifdCVZ+e
rk4AJO9uNwohLkhiMWFa6RmqTs04eBq6et7hBjlydVnHmD3NvBB3d4KkZ0t3g9Zf
xvjA/CWN4qPMutwdJZIN35ML/7DG+MuPaaedtQzBrNLHe1yqWZTPhvbFOAvxBcCj
eZKJ4Kpb3xcxc11R8nN2KNuOslru2EHnP/+A36FqMV4sfBY3R4FpMzgtW4JCsEOO
v27mjxfTWh4VrSJt5Xuz9kX3Ag1w9ZigmLMbpEApUQ0+ebzWLslqjzCFQgDbkCh/
wio+vMrH8ktcfNMGXtHamtd7c+3NtDU7rB6ZOzD0yl6IjEead0gWRMl4THNjtmN9
/ElRsEe/7OWPhX4A+zrslBLv8b+od39wgjbZG6cXLZoXmcEKLhDLVr+4sWeEgLh2
SLpGpZfSloJQoBvoHVHrJcUdviNuEEZhtvcx44mtF0fkB8BahE307IFJ+3NYvcVo
iGo4QlqRHq2sTBOwFz8GnTpqfJ/9dwELwIHd8TstZiKU+emZzIcjVFeMWMKCCxpP
5y3ZtpTEapkDscDC2mBCQSEQqFBBZfM1yhpOJ9UumNCa3Ay1c+ZWVuksvE00E10e
q42I66NrOYV6cMXPIg7HbdIPtwW+Ba1062Vh4JG8QCMyorHfIZfd2PrhfJNZvKmD
knV2JJJvOEwdoiCjE8vDda/5qF7l3hpr7yRJbS/gGiIjMA6HpDS+/ds9SPis8CUX
CpPhM2K4aTrHBvBYzziajE8u6Qaf1bIHkOoDG7Htfm8FY7yGVrQj2Z81QSlCHFp1
nL6hKBTQXXwE8QXSp1oz8PDPJmmu0foh9Hl5GCXgJMvs0aoHdmM64ta71jfwVz/k
gv0QThwhFbA1lzFIfazTfPAZwD7s+wotcwLtjHDlBh+U6HXglRI5FOLbg9ZJMewt
gVIxVcQIpyrep3viBvrkGUxOG12E5Ehcu8/3UWB9mv6WdaRJ622dion/uHJeuZ5m
WP9B5Cx2BdxKrHnR10IRD1CZ2cSuIjSR2ZalGOBl1OjhcK6e9/bKz3uQXdtdcHkT
QML9LP/7P6WDJ1ageklabSZkKcbdnpk26Q6s460S6B9356QAKt1dJUujyrJMI0rv
HtGQLqsXNJ4jPEL5v190os4fbQQuAgoHqR45ol8nnIYTV9LdqUk+Omn9CZb66N2n
NP0pMSNW/aJDzO84sGSJ3L+c4GXwWO7o6f2CNMPlqSK4oQWo+S4MPdZUvnBxQQP5
VBI2H1VEEZ0pqK1i/KBuRaFvLZRFG+kTLIw+cudkboVYs59hsnHIboOAyI8cgDOU
XF1SBLlho2aNRo0DE4bETBL0TssqdzcOu6d2LXM6XzLKuGvIu/59zJFftS673BKA
41zOSBsO0U/i77i37Dnv1vc4XptsSVHKs9xl4d7Ay+wdToVBZm8mh3S3CXq6wS2l
aMfYMwZVwtneUJldeCtDmDVEPfznQFK5p9KIWuYhc++gGc+sdOmT3fp4RtbLMnD2
uQwZYFKnRVpAFdUfVax2JT+BXktqM2CN8yJOYchhE7rtAhWWzQXeKTgPR+SJuZwB
a2QusLAaj6FKtdg8ImvxWAY0b+97XHGxAmiOt6VEECPbzM7eGFjT7b8dZmKWDVz6
qAT4x+d1S7kGeG5XtAmD1+HdFoSE9qPPdKrWfUZabFxnUWTmzwv/gw5rpkSefGOv
zrKyVeEX22i7wjh3w+1UHW7HwnACMZFqri38yWzTtuaO/W8fj3kSb+5g/WWuOB9w
ycfCJuaWnMzOqOVs56BIH+4fB0tG8c0D1rY/JKLCW6YGITWyEhgtB7gYDs9so35m
YLpxIlYSLyrdzK1xvV0o1bbqcnKZGLVpHV4QUnMQG07ByxzmenZJNXyRxtiuDx9F
SMGKa+QhBRD/g/DrrTimwMsTB9P0IiCN2qSTD6bsEkWtaU8uVGjtxXpdc08ibGU3
CAvE2Jk+H34qqRMDsFINzj9r4QjjQF1sac1w0bduK21rb5eCLpTAeOcF9QTUUKp2
jXejN4go1RtnmL0rt2cL/9pY/IwmFWWhgwBqmeu6f5OD1VEZ74yRgdEFmbhj2dnE
zScEKLiCgpOGVXNbJqMpQzA4Q66Qpm7JE11b/Lqi3BxSceII5sF1aeA0fCp2s/fv
QfuzToxWcF1FqiFTE5qgxLSLSMCOOR8eQdM9PHS2sbwwxy7asJfFofUKXjtnMhXd
M7+2cRGMkZtIJAM2NzCltBmf8JQHvPCGXOW2Dg9rqCN7V2mKbhLTMW55Rgeg9sJ2
a4mGCN43unxiUBtZVqff7K6DqqRAa1T4Hr0bU/0rNpMcdCKU7q4hRKl/pDEDH+qV
FDZYlGWMo1xpRVf88BzDi3JA6g36+YCfRoG6zTcVArWQ/j8WQ/WsFsC8GB7nXd8W
52pKsr+UL2EgHj0If+UqizaiAE1rd/2ClvuvY6kFgsN932LeoSoe29HWCGHiXvv/
rBh+0C6iL2VUfqe4mrQGmHhLzT2eEZePr5YZ1goU6mu1ZOaGWHUVP0AFHnVV9ZTl
ljpuQvLkhg1UDl1adw4fKYsjY95o7zt+vHi1WZoQDodIslJM1Zu/nN+msEkZNxWg
p2aqKWaSURygNmhFcRq/jeN7U3z66HMajSplGaYYniKTX7QQCmQBrDuJeH076u2u
QzZyJhe7Y8Pvyw9Falm0spmMLAgJB5mvJv7wn4Ut9262xNbiwmbQTkMAwUVGEbfL
Ualdg/a0ctMs4+y7TOv1jG8M2OAGnI7AZXk67ScP5uwV+rV8/aHKpe5Q6fMRWh5y
PAPQ7pvFDUEPPRpKz9DISl6moQ75ON/QagKswj4iP1fEz1J7epAW8nYk8udrDftx
2R+AUSUnukSJPl/7tmApeAIBnmZrLJFkrgMPiWzjkTIG1WGB0ZTB9cOZfI5qrPVA
GKf7r4BK5Pqqa2UzDPiqEi+QJXSK1md8VyLhEyP2DkYVqcjm+oBt4TXMgokHPZcZ
HPqdP2qnB/fJqEcOfItsNSiBFNaYLBBXDYKoJm86mtpjeGnxcAm+H1xOINiDiwgC
Qq132PVrGR+VlPd9vlJhKELGnHJDGJNt4KYMNAb4rX+rjB49vtTeGuvHMIN48uFq
60xc9iY6rbpAr/zbSKUzqb0Sbb0YdY3K1tFQs61leYb1PRrmwxARE5Wbijc0LGPe
JbvFjrRDSkwj/czZJbFdRjin4gaB7WLuqoChtLvNnjjONlhj5CmwUspEfq4d3opX
XuW9hqg+9Pxe0KdkQBLKYS6LMDvWOy+fuRM/4/RBgSWQxcpj1havCZhy18xkTLSe
dTr5G7nQOgvdI7bzKcP/ovihrmcok9I93nlxPNmHTQdVFXMn913gdC/OxXi38bbs
cFbNjGEuOjIOT94EX4j3NPyShzKzxrzJ6cKhOQZnhXM7B4chRRQ92kU1OyqrXTpV
XcCqU+f0brCOJp5xqmMWabHTu0zic4PbLOIhO0R5JDXH8ix9lUVegwRhL/nbRmr7
qQ0hyX8sIvsKaFBU4BAR5xAyzfEwgzbiRllEFVdcaUb7kWB4Kosfi8sxMnxUzFIp
y1ugy9u+XCMA3sBIxe9LwSLsxzyhmf8eEp1cMOJ7vWVH+r3JNH/i0ixZQspSy6DZ
24/I8zaec5gCs094G4m9AHng/ZIqoNbqvvP7zNFUFdvnX/omX2UVuKdhUI3t51JT
jvcVMUm5iYwxlF+416Ycc55Aen9r/xnso3069RU9mpJYIzdUXmbAKSoO3OOTScLr
ROpt88SJMgee1HG+UYm16V7RKMVBvBO2DuyIZgl1a+vlowKtN2XwvS0J9jxDeSrk
bMZ5wTvzmORLXz6/jnb4P+vILHD7435g9X32XHsXlpXEZE5OnW/ZpuytfRNiyf01
+98f6spyvw/E4ROfP3x502iWU8kBPx3grMUBNsg2UO/4zfLIenKrH3Mw6mFwTib4
r7d6k3q3p1db1Qn/Iiho4Tub0LbJ/hIRWND3WRRihl5sO5vuQAKWEQunkl/ZRGPr
OVU8h6HCu+DiKwU5yyNnToagnNjvW7r7ISOP1gyO7PvUXwI7q/t7wxP0M5R0IkKs
mZ6jG8dLSxUSxaVzUgkY1jVmSrCyVXXClGwHvKHX1ndybx60PqZJhzghFbDDHWmj
pbTQWv4KVPExP0iLSEhogDesZmYlEagLPiONIdLafQMchh7hM4o+kI1jcZxm3GCo
HEmgB3MVibj+mTfzh9w7VU8dji/GM+aNVEhGudhaXyOMY9hziHGmdAPZmGVQ/5wC
rTG1CRHQJtsSOw4Qmk+yWFZVWx2yy8a/R6iSErLxcCcxEy8U4tnEKCHIOXCjI1b8
Wnwa9zQa7K3NR42Y29vDKdj7vmu0dL8+XrLIPciKFVlmRxvHm8oGrjlcwLPm+kSh
YCoLxWNsq13/IKaR2YJXMeOw/WtG/ohEV60pb3Knwr6lOh64BgfDH1SWzl2gm27X
j2j+jgkYUqxqP9PjRgdI9G9SqpxtPGWhAemdJV/IWeciwkh1vM40yR1Jn7GF5Rl2
YLgPFQZfvh93MUN3aasldaWLY8wuEEQjLKsG1r/RnCqGxhcQ7owmWjRtKeTA/j/U
3FERLBIjzPYjKv7lciyhNAvFME3C87PVSDc9V5WyFvnyGJEJRzVkvBbbUA5NapBH
D+SRzvXNpRE2MWCtN70TkmNvuSEjmdqmjFf/Df8gkHKNtgLlD2z9ZLnYoEwsEsQk
H6A7+UGmbDSMqQJE1kfz5QXITOHyJiImUOSY6Ptr6fJEvWquSh1ViWi1UYits4H2
dAKOJEqtwuiZlQ67kQaDT1XHeba3Fvp42Li2nn6WHfd7flPTU1yD9JroOmtLEErg
ls/Bsz+Hz8XMne6ARMbhEGQ0L5iOyAstQFXjJnGTtq2HN6nivHZuZEPpCJ5bnQxt
ec1VG8JnfmjwOqAALL1pR5JH96y3VshuNQ3Xf+7vjlylK6GZsdypG4qJ6xzMdTtu
Lu6jlgeMy7bSIzzg37p3Gkfrr4CuWIVUCKvlxel3kthj92LkqgurNWxHD19Bn2fV
9G3oObr6wo+rOMnSC/SChE8Tn5mtllKrrsqD1Qa5+vWRhKO4BaE28CqnSmyBtXMm
Lk8XV7PR5ag8CY2aEHYEnN85gPbcNyE5iG7S+Mn/SpiDexvzwDl9xRv4DARnZC1W
FALy1kE5IkBSJMWGfzkVZC8FfDmI3CbUKFzl/ntHlt3F+gkU3TIavpGZcFcfJaEZ
KVnlk3msHlTIo5FJZdtLfnqsv5fpncjydm/OTd2aIFmD9EEBWSPPsODHFESHggga
XfE2z02tAL/frNfTkCHNRI7vgty4gFGmLxeUDHUaP7mglkI8+ogAKffdCF9hoe35
brf5mzJgyRKGuiCNCIgGuL0NHWfhxL3rwZtbGhBwbgs+4NjtR5y/xaWI6h8OgPFB
bRT9yYs7fkSKwc9xNwxCpF0BXYVCT5uAL9icpROa3f++/LeEfm3VM5kNPbqTBPFk
gqrddwP8RkA0AigCcIC7LJJi/igU/gSCyOonxSFpuu+TtxjRnBCoa7EOjyWuU1bH
dg7pdU2BOewxnvXqj5rYIBwLsZQWLaBrv1WG1l02/kS20SSVL3JCecFk5vveOhbK
nvKz+iO/WDCuy/XfDovDwjDvm+twhEr2X/56tA22bFKaHVvAtea2zlqFv8LGRqvX
hbf5arvNnF2DuUrOzK56LC1XVm3U/+zUnOjpPtkpE5p187m0RRb2HqYSGwmP1LTx
UX9a1Z3kIrp6gCpsIJI5Od1UpRJa9GEmpo9BE0teM5EDPfUkaNdyG7zkXQ9DKqk1
fE1vxGZ81oOcdel2MNUR3R0FA1FujxgWlIBC7+VM01yIoxGa04p9v+KchnwixV/z
ZTe7PHrSM7yNa2ZuPTR/N6AFVCRth+v7hMaZ1jpsvnsOGJ6WjDV9Kvu2HwyFP1V1
+7BkVG+TWSbkIOfjyPr7l9XMA9TPcfGiO9piX3TlhJyMH+i5Oc/iOWjOXyGSAaQN
iKkK1oBYo/H+QLy5BoitGQsKyKfftM7eWH91snO2+1NaPhnlnKKfUIuyGSFHg9mO
7ydbkjPkKES7KdkuP3G4K+7Xaboz/KNkOiC5E0DxtGyyUgjbzetuuGxIK8pjdP6e
Q0yILxulaJ0dmpv4anYXqtOHCkLT8doDZ4jhWqpc/tNT41MlHmHgGYjWqgLfUM5O
d2K5C8jgc+qU65WBhMEykhKDKETVIYlQB7U2KbM4AY2H60oyb/NXKDqFwnhWA+w6
78VMM/Ng/nYyTLV0HrbN0/wLggcpJTZr5gsCC5l1qdEKlNrJu47s//tGZW9XFO12
Ivv0Wiu6Z18aoIrCqCBlYcTAd68KFlOWPHpHy5pp0NRmYVl/4aZ6peHwPjHhFuMH
W2jmIVnIqYakvThiZGucoC9fSJz1SbHxycapvggeBI+10mQRTTduH2/R+bZbaQo1
342p3K6x/3CN68eTzErCIWlo7VOgVKuRfxV9oykMd/0b1c5yx02n61cNLLwONmSp
2v7KwXAte52IM7M75gBOx4+ZlGMfrT5Ma2pGxUNoClW+a3GptLzG87y7N4Aw4mhv
F5j67P9Rqua1e4+fdXWzxicmzgXDy3VuofGsctiLJpgqs4A4I9luJzYaqu+x91EH
Jc30AvCNOBPvA69UFoqWcHNEiLtSOJP6hOfmZKvQTwHIjgPtil/65ZTe+V8/3Sk+
O6rNB7hpxfRxv1v3tbeXXPwjbW5ZKUEJGh/RtYlw6BIZXsn8oPwAvLD8twfgBXRP
Nwc+UrxABp/JHlOURipUEwQHuCDCbt4pErj3F50iKE35/Y1I2X+41Td0axNg0LYe
AtzfZNzn2i3JGI4XyudD/1xgykgMRdTldLM7SCR70Z+xaGpbdQW6o02uECnrVkSI
gbDvat/tQFZ8ILtxfAetojVYvel75dHkC+/0Rj5YcXsc4zflFOX8IL1MbKs2iRyG
8k1u1YIwR2BKlEJFEtj6B6MtyNY2yPH+Z7L38LsBrVOlVbdh0SsY8GIyPHDxmczY
F+utjveAu+EzfGY8/Ge0mSHOl9boTwS5fYui0ZyrDvfsSzf669uHVtHHhY7NoNOb
UKgQKEhO3qCJw5ebl8tAfwqwx/2p9bKIs2fPmJbeIeZXeEcfJwwBeUbbBgnkWr/s
qbdE1rwkamJJid9cUaOzAiIE1tWIEtwNgiF0fLfkojaPbfObQC4LAd5aDaLkzWkm
DP0BElKPHPQrd+CL3Bo7UmD433iPYjFK0y9WHsxt19gNUtynrvBgtrB7oB/CCaVW
Q61pgnMtfmLfCfa5ZgACwXmuSrisjqITOHEuD/sq3yVB+jdjVH/IXuCRKL10wPod
pGKZYZedgPMecB9EkrPNztjQOBoDs7TtmZgbb3QRpcLYFHMfcw4Hp/lVZCnSq/cX
j8wOxZXfgC5G14RdQNTfRwtRHZjdqSXJ75/isr2H6cWdMsERFyauX/4dOUfH/c1a
v3xInpJFqa9g6njASGqrutTE+igdffOQg2GLk2i7TQMdZcSx4Rwqqb1fehEtrAPi
lObNun60L+5HH1IYwGabiCeynDQE7kcCzG8OEvczfGdkUalX5n19Jwzf4iIK1xPM
+Clr1QMrOTTsVHZmVWpUmWz4W01rCuH73DbIv/M1z24sEc+bV6X3yUhkkIeb1eY/
BFdRzlXl0poBfUwhj1pYMUhKgLCcuM8cK47Y02ZsAoVXrOZGuAXe/NSX4GADsn8x
Yfu+0Qv31wBDmcusCfRrzwY84uwePdW/tRyPHMWiqx8WTtdAzCEmjaj0TWqu/6xk
VMpyh1dBdu2p++lrx7gogvEYrigv9XYkvnLqEq+Ab3palwr/KhKhfY4a6tMWWhwR
k5wCgiq4gMvj1XxLad267CHTOYe2PJUuBwFtwDzLH7kPQwuC8yUOsWDwETPvGrLP
4XZOP6RKKDhzyj4yvwVJMTlW1tPtLrKu0VyLySHYtZL+OIS6ZdJevMdGIa9AVntA
gxcohqChCDFPPffKrsKD6vZbom/yMyH2IeyO/p44wiVNpPHHA1oPjm8NaQF5Bnio
acCoZ4VDiAGXsK1/LohJHI/lJ6H3FMUmQyTbm9rWv4FoZK3rpPxEwF2Uftbc2O1p
8J8PHmkxpkV4zG8dYk59N3gRv1elDw0L7uoRRRjvL+L8owSYLtBO0DlWIBTxF20Q
c0311v3oRyCsCBxCfTIotvl1fHHYodMKMdSRbmENUmM138VOn1bv++CbxGAoBikP
cUvtF0JLfm1qi702P9BPCwCHZiZW1uKib9+3b0YqzfvcXSa5iLptfxth2PrexbAM
BtXIkJrnIBE8TgaNoOEzGgw4jXcf3+JKWetrPPB0exhcPNx02b44jO4Q/SSI/4b1
1MhaPD752j7o87VOz9xoW0BjyWtHqZCnJiCU1qUqU39dr6BwagPYT4DI1rCi/0Cg
9YXjinnsOdQ8dSb0lftnF2FZqLBgCcifnhw3PXkBLwS0lzUH3MQinZbWp2qbm8Pe
meTSAvUg4mGxNg3D2PBpv5c9Q0qOcxPYxxTQGqbvVzKOin3+RO/9Aec6XSiEWxnD
+dPDUffQqI75pXrL1hnqqzHm4k+5a+vQLtqEZ7yUNyfDtwmCHbX86P4T4q5iyzRx
fPHqcPQ0/TkkuwVxOp1QsHq5dibzoDxm6640m7vvpqZPiifg4Nc6SQcYemeScQS4
txsip0oafAR9gNZjArz1CoruQFSPmRjMdjrScMuk03ps+VX1kRTReQYjQWahp9ou
fHeRw6+eRDWfDt3uEsQXzNRXcofkdn2FGNy0WaXbdbBiYVuvgWC7zfU0Pcfc6UHh
22Wm30xT3ohhSti455a5vPcUYo03cb9IJT+LlUhOVNYRQxSm5kdA9siuXCbYd4oE
eTc0wSX7GsdovUyAa/ISY3P+fAOCkDAxDuLkvaLLoMeon7kAw07NocGav46RWnDU
eDYFlo5afFUU/t1eeE86yWTQqEj/pczzt3eyTpEALv9plnoNpEQcx8wg5/x08chO
vZ2luouuJYw3xMag7uqsnY46FSZBWaBld1qVTc7KxBitDMdiSV1+H47tW6HroS/q
apUgMpqNrMnqy+PkTYel9Y6ZJh9xvsso4yiSwDVTwdHDhwfmTNV4DvOtgL5dt5AV
qlwnBPyK0H3rkfeQ7S2hkqDTyQ+EPqIllbG9grnErQbrUe2QghFkX7VkyJhcpAyA
H4Wfo3EYHmzkIrLcEnh8z2FT5PRlyaWlW4ZufzOiq7EKAf5DT+YXiLsM/8BLE1rw
3R7yOL7W5I/CDEA1pdyAkLkU1ceVAqsH4FdFskkgbZCZXvjaHSI4xlBfkvWn6weJ
MUGQgSlGVnTewI16uUakC+3rQppbGgcX0u7b5oOGSQ1/hdSRzzD2qh2N45DY/qrj
SF1LiPUV7bg6V5qdkQkjEiYCe7iE35Wy3Lz5IdmY2EI8RWRPOVk5LSPgVsnFOP0d
8jimk1hGv8gzxGAV9S4v9ooIk4FODKQD+WDmOS6jnKLeN/MUiIfuvF/ClOT0MkBD
NQrnPwWzI/hmwg0eLsr415LniJztOhuMFMFIKmyOmPEauCmBF+b8V/czpwz4t8kJ
e6XSo0UtfFlBijyhej11xb38upOAWjUKuYUx4d8+WUEercNxgysRKh1+0SGAAAj4
g09tsprjgsbFECcJkllk2HkUwu1xKs9WnQYxBDnRBJjSi2OSDUZqozNisgy5/CVH
gAiLpDCP/PSlpPWJpsLffgKBsTPjY87GTvN43U5rg6Rs5GNjGzNxAnH+Lu/SpZgY
0HQJb/lrNpvV4KdDK8XWx2xZ+C662cR+sFev2amwG1QOCE2WGOgdtgWk58BRfedq
LG9I6SoqbZGz2l/6K0hu4BuU63Q7g0xIEoRjs25To6Y1bHl618tz9KG7xvRcHs5N
wktgsrIxmD2aDTY8CGiEy3r/wtWU+mgQKyvaT97txDcj8LeUQX0hqHpWBiAVmj4O
X4Zg2FBA48UuJts5EyWDHRB7/80CssoJTToMv9uZcxsu6SQZQhU4RpIXb1kGQWoy
nPwL+OfudIo6IwgUrZzAOKN1yK1dMHfv/PCWEVtGXetvLGL2Z+6JqLvJMHTofu/U
9YEXZnuExjiJzdsJ5j02Frhc2dRPYRWcKlj8fC6ZcoNKK8tZJtQM2dbb7fmh2z5I
mIcq2bDBQxHO7Gz9M+tYR7lOapQ2lVIVrDx/z9G3rnOarVK4f5oFU45IDYvsEiOh
FkPrAzSUkCiTWsstCVIPz7es6hmrJUOmKgJ5dtXgkdy9dA0JcgxKIbdDErIAGSTf
54uvPKQgQfJkzv2YdKD4g5anR0NpZn8JRHb99iV0BL5fV/4Bon4hvlci0smtGdlS
Sbc57HKgvakbikLsI47Z05pVhIMpyx3fkoxrRQe1UnU72Pbw8Y8U8F+JWSsymCpZ
riMf5dxdubYLIHRdfHqbt4RxfR58hTy6Z9nUMXdFuSuPjemtYJ5dP5/Cga617slY
VNHeuq6mvbtk3wJwPMaWfXY17mIKnvpjPiTIZWhXrqoxE72b3Vz5Vaqa+aEWIzpl
eWo28YVJQ2rK/wvgMH5V7nbQ/cc6iRYa0e5hYOV83HaZkUKC9zpriVsgJLT9qAqR
fNgGVlqDkXh4cfqMfNCTVsfb2ZNRhl6VmNRWOQwV7x7+SBZsk1Y7hD5oI7+kUtT0
dRI9MeJpb+Qwtlugd1leJhP2fJKfeYllGGQG/fZ+eRu69PgrH/oVI6Ue/+Niw54Z
b8/Un6VfZbFeZeAy0OLjHrYJ+lZIgxr5sHSzAPYhH2t1NRqaX40ZN8zvy6N0dQ69
+tuCLc+jNnYfz4mBPq7npeZf/UwmBlLfKTMS/yQTlYDNZTxTToiYj4nspIvSiG/9
QC6TQqglKnWScV2iP1fE5ATVf3oWwqIYXmDWbpgtCb5d7R5DfWfWMyXyMSJb+zPA
5MavGma/2I5SsaPqL/5Zt8f6Cr4aNrt3CWAKI5FU/FzuHpGHPhGRCHtLzAxBz2Zi
Y4w23aPUWN1e9THvJJSVForTIZQ+rYim5uC337cQJyut2t7Ip1X+Maj3IXCXInKM
ZQJtICEyJwK7fc6TmikApi9lJItDvYBVFo0ym2iPCac7jf/paMhsmlImJ8O4oe64
5LKjbh1t0BAvvkSM3+7r0rPbY4hiBAmAVg06j2NwZ98RL9dBj/arLwYh6Qp/Ll80
LkyybDJ0w3PPENmVlqWOQc4rrK3/QyaPXnmdbPitM8hMqSQww8+PTSB1TVLhe4V4
zfPyJAOME9F/5VqRK+xgTXGfVlw0lmkdb4s2ug56bzbrgafU8TkXCTP7W1CLh1cd
Ekk77+3Q+CTOAifHKvmOGdsWQf4qgl9YV2OOUbrFPlalhzZh3MVV0ss6542Z3l7r
6m8GRAAqTzsu126z++ZEsbTpdQ0MCaghchK2+jWhsbj7W/HgOCVwjUei4tFgm8Gn
jKQu5DRv8xyOAMf+ckkD5WXn9a0YmRBlWnJ1un7uTsVw7FydkVVh6qChYgAXgBxM
A7+v8/l73kWcZTvpwYqjWQxsLpUzLSrE4FcvQ44eBsjJ8NnIbe5qZFBQVDkdHazW
cybzVKtj1LYkyoKvMb6DwNuVK+v7bQE7FfqMse97v+twpnKuSXDHp6yJ81ETm1sv
HXh+pX8zdOQ9Zd7YzVlG3JI5gOHz30OWeBpNeF9bxAnGZ3/yEaBhPKVlkn+TcWe7
Y8bwcmswDYxDtnBQptd29G+a/Ud43esuKfGtxCeOkbdlmMnddE15ijIvQPA79Tis
tFVJDwdpGzEu24bcvZT2HLSkU4JC4vAQhe9+6JKsoS1DxTx4ksjGuWVXTqc9p4Vu
J82YvoquSVYvXrH+CfyooEdF4SZc9sBHVu33/0Db2nzvjNsouCAgTfqmrG1iJyL5
D3kwTkhrosE13cARnb+WrQT/APBUC9SUuNphr6OQ4axqlcdECa6qwkHRoO1D8ie5
P17A3gNvP8CjQAz5RiaUn9VohPvrmoeWnMESbV+9zBplzUFqKKBFdNDU5QXe+V2c
GurBZqwzSCx5ZGgs2X2at7DdJBNNK44wfpRI9Cog+hBEj+Bt0ZWJb2v4d1hImzWB
ujWFhNCgtroArLNJWwddDHvo4Zyr/lztQrXEtKHyr6/NiP+W2PnSifjTLX9i0pW0
XACK+7NZ3UKZ14uap9bl9PHLjTd7kQ8Qs0H3uywP4HGUlmOpVxMYEeg0y+C08HDw
xsluL/NU7guqSy2N+LOswjfl8kwPiL9IXx6/NXscwvPi32mYDzijfoMnNab20cpx
EkLpeBRfKW79TTuZ9sYue9j6M5u2fbnSXkWCRrXPAdTOlmC4wYrSstzu365B7ACF
drs5YotCtzgO5PCrDq/dudCxQtvzEuEPovoqpV1PnLf/l9AvLFBI4GZnpIrjbUBv
edTPvirvKoVfFoYLcOE+oEUJz4Ebh6pqu0VVcsFdVcpxEUyKGU0qpgXvLoXaBdVy
59L2eV0j1Qf/R8WP9WMonY0FVciG7k8p1j22eZg+TIN4T02cH4j1F05pPN1pj6Hq
G7qiS4367hg46b2BOPb50bRsEe2zk2aZDimJCrj7Nx0Y72S6vuwjH3VBk717YBeq
Ocp0Kzxa8vbq3XdGdCsLbH35K0IFvPHud9V43PWyXpKmOG1NS2bN/M+JKUJ8m63I
hxQZVswR54rfq4yyI2cFdM9yD5ktAhaWh0x9uAFEyTkgh/7PS/GSzjLEVy9TO2Qt
OnKamUSpK3EwLmzEjcFdIGv72JdICpvJvVcO28NHdmTseUQJdegEtibgUzvZBL3B
Z8EIvTvRUPsp2zR0FYZvey9k9jZd/wS09T3njqVseR6MgrSPMnAAeLlx29W9dZE9
4rmx6dbv3IGwTpBZxTD2HELLp0+H996bTN65hrk5owPPJPliKuyJTsXpcLvJ44Wy
zmBoKxwmKBY+5trdAaLZODNbXJHCsvB7x26kSxJgMmw4Ku9mj+aHaxO8oTvcNBq7
E7rbOaB3nG4i3P6N8c+w01S0wCHfEfOOVSqEB/y4GZqLGACk9fXOlodoR1QuA7R+
GG9sVMSjr4Mos+ujn1Ng8LAY7hqOLSCa/UL3r7kZH79u1z1JVynlo+kkQ9PD57DP
2AWuYU5xA51e+iPrd2O0q3kcJSggVHT+q0nYcvraiAfXfm9sl1LGIEf/sjdR/onY
cYpypN6ORlyX5JUxogR9u8W3BM0TgaoVyn+itBFlC23UhGfYC9Z2Q2rzgt7wPJNu
gwL5tnf2fmpUgPmU/z6tEEXlZVFjs4y7RCVwAb1pelZPbHuPTeuhpd8JiPQTtQQG
8OS1+ny3Z/YqUhD+i4WrJLAjamShqiOnSUquYDkO8aHWriV4jFnFpx+cpflrEWvj
gAO6Uu8+2U/jDOHHU7tpo9NMLCGl/aOJhUgWLu6o/IRM89+updJFFHwclI0XE2uF
L/JUApGU8/CqkBwHwLahydQJGwPwpyyYVfGInXTmLSx+1eq5/6qxWvlve2Dpw4Pa
JUyNg8CvITFcE/E/rFA5lTp7vVZyr1Ralogc0bZi/K1iAoy5i91kxsaicc9A2903
WHhssw3WPmct+q7bA9JjPLo0Q4JpaaeZVypYJKfqeWfpiikqhRj8O29VbPC4Kkt6
1zLdUOuU+i9wr9CZZ1FJgioNdyQwMFUhkcorjcYcHfBDciT0gxD3jHpnRuhdeNlh
Sc/yHwi8ibZ4qpeIxSvBl5KPE9hh4ogxiOgV3mDbhWr7qPi02TwTPP6+Bc4/XPv2
TeYGIypplWoyL40kkRsiQWyeGvdnmy49IYgwBKa8HDmSzx5OQAM6AnXrIAz9HKOV
S4Mkg7vfrcFLCTOKCQb+bMBZ+stpzSO2J+Hgp0J1OdIUnW+jhn7gUQ6cOydwFnUU
fn388oa+xgaGiH5iXUiDr00HUxMZAkLEcwKeHmLvpcK83py/DCSzdLB0l37sK6cW
JM2mwS2UZGiZT521Z5KRzfORCOA+xLmvLu8lolj/PiLfOAhFrG/wvcoib4wlCS5R
fkv3+zAq6Mqp7c0ZfbIYTK5K34waMBWGc69bQBrwWs6wtsUH4rLZpQIVKCCr9H05
8iIDxe1lnkAc3I/MtCStAlwuPgxmyie2bi/E1jQugTLl/rIxLHNQ8cTkmvSmTVNr
auL+DWWhgZYGODoZt6TdUSbAr3Bd/AKmN6ilU2BUNzCLH/Pg8W0Z6i7XT6hkoqfi
nxu8pjJB6TfKrgIegQnaSE60IqzVWcyfvjSYxayhecYj8S4NeLcJybXEfphgedDx
ossMgRBm/VVDoPjOVfngza1b0Ore3m2XAy5F8LKAdN3PuoTpMLLhkg+DNkKvd/hJ
y299K1ZN2X3XpYYh16wJvxKM53XrAVqjYsn3ZUzGCD5TpMxakKpYqEVPB5rqyq20
+IBmglE2jwoDQi6o+JL8cn9ujWbDDMSQk8/OXlnqyLLbCG3rnhkVKuPi01b+cU6G
iaKnha3S0sUSh/qCsv1Lv794YguQUaEKeRKgBx+WDbFr32wztinl77w46Zv6Pg5g
JGO2METCAJs4OwJ6i4m5MOxjkFje29eqCpnyW7/N1UwwYV4btqsbqGsyzy1xMKyi
Iu1W3S+ESDocOdlTwf7DUgG7pJcnJ9V7PS4x2csNl5Qwrd7MqrhTtPJgUAYKDhzV
pdygYI4UiIpRJ1GfQW5oybxYytXbn+cBmbj0Xvdxv5CYlL84rdWe8W40UjaUB+2X
eQh01TnEZa/or3naREQxquj8gOnVpnPvMyx0clAmLGbrvlW1UQD/DPDfXZlqF4m2
gcAEaC2EnRnPYPzALFCefgoH9P9MsZ5G5ENuB8NlnWcbiH6iJowenm4YH3qRrm5m
6pEb5kYzl6LAb5T/nyztYx7a8HL4ltE/Eq8ozLSa0ImIlBrhq1Rk4b8Igv/DAp4Y
/mybHeKAr50xIe3X3TJasxPoRrqTeSCD7WrrReQhqp63Ndl0fSt7arwc4edTwnUU
h8bumBIJ3gih7de3FXP6OkW1CIInrlbndD4CSmTRKF6k0ry3GwFnFqKFvVmQ7AXl
szESy38WbDnzWvhHLHFdk/DbUXfglCEsK195wt2ouZimnrFUfnlfGT82A0nf7pST
bbycFtiIUXX3JvzD1zPFt1M4+Z4ifRi8JaqAIrEjEMWRu4sw4qp26Tqzi5XxLaBN
HsJ1nReoBNoJINzGzkQPdgFe3r9t8I1sSyI3z1u3vEu6EznMeYyLGNIuvBG4Z1OP
+wd80eG9yRK+fhfFoRqsJ6UOkP1JaGK42Jq20N9vWRUIJR9sZdYCIyz5hjDpJ53r
D+xaAgSHfuZTGOB6Fp7ujFGvtNlC8rn6XmvYMYrnqXYlKeYwlCGKpLc9DXCUQqZ5
3fNq6KlPFheuDhZth15Olhr+l81fPCCZoLH317aBEN4Y3+jHD+d+XkDMEpAmcmEr
tZ3kf8D3sACwk7B4qhYj+WmwkQmNrJzue8MMuNDMuz4mShQkQ4MYH2ozQchLacgZ
X+3n6n7fxUXdykGednI+9IA2+sPmwpKHyuU+kFYTg8dst0wG94exHPQfk22Tfyd9
8XyRopIemzoYgs4gNvwYwaZdjdtd5Udi6M3+Ghtc9PO234/vYuYDqVFVGyzj+S8/
RwgjdljWOOT/pJaRYBv00Q+pTJbYIhIfTJGJ8MDnmFQDjAJbM6yu494kx7U3OEq1
CBnPBH/inQSFKDtA1LGhYyNA2JG2yFx0VzTJCSx9+rnOQJmV+6oNijMMGCGF69yl
sholBp0KPVNMtFRWQuA8ttZ4fuEyn+3kb5c5dyW8HdR84grsSImoCQ4HoJ/89bFo
g8lHAQs5QpwjoQOPOfvw+TJ4nl9XgOxt5JBtyeZywFGxO/lBUQsy32QNqs5sjBVn
mCAXhnCyiNIXJImjGGkkQsERfj6t/QjCy+e+wuwiXsY4SuuA7Nif0IRXLolevMws
GIOf8jc+EZPgr++YuoHHsq87BGy+dKgDJhZutzmaudznUfa0ouHpKJ54dftU4qfM
xaYaesB9LfXBpfuErVxGuyIBwdBiCkNStzlx9YBHP/9w0SP/siwm8NKMBIiwY3vn
rHyIXF4Igb6pUvWAzqjh8Q1baH92IOTcxRTsimGzeA0mZaZGun01/0uOyKTDMwee
zuLw8Jtp1boQQ4WTMwY+wZD9Yqpr/kUENXh9kQu+l3nuLu8bmjC9fxmD+vGG6c3M
uyGw+Msud0Mw7hz1mjaRMtR5H7UWx00Jqw7h19fyUZkaMmKg+sdx5/JF6eaxDzuY
vmd+Pp9On4wfeTYZokfur81vsfqzfdxQkqAdFF5N7iLfUyjzjCZmOMweaF1auLad
qO9J/N2ATo1gBQzoOPFW8bqpIWwNi7+zrXCfYTGB9yEfC0eapCCrIA0McFJ0ER02
KcgfAazXIWT9NfDHudo/fzXxVzGxiJp/bcX8P2zkcX7yP7C10l5xgHZvHaXjbgRM
uGbWTNGOUu3ywsB6hDdt58wjUqQem8vDf5wgMlOeRoYNjgiLNFScUUO/JUeBJBOL
po1hquZ0OFXm6QbI2ZdBTe4QBn76CM0xXX/5jK/qW/Yer9+8aYDZn36s9CAa9qLa
TQhhrqqwckT9uLhwRiSIehTTNXdPb4Y2DXb32g4Wxfn4l9rS9fKao96hbb8fVJqL
djaEgIL1CuzJ2nhAKKkX86ymp5beqUfs7S8kTHIU2aLg3XUDyDnokzvzheuFWZu0
yIto113ardy5JuD065nhhOKBZmMjVxistlJuwrloN7gmrC+KB31h7Cukz/mnNxcn
qt66F1I2Eb67HIE2IK50pPv9zGEAwg+Wrjcb9dhPUOp3rYtoM0SjbilxNkSwK15Q
eG0Ixed8cTE+rRnGMjM6N7ov+JqsnNco2HouPqD12Zo4ERn1/U9kgd0QeSXmVXkB
e4TY7bxsDftdnHf1Qo42gZGVKl8AYmd6fuk0jha+uHWh/IzAF80V7L1iLLJONeWN
UkYMnJ2E8zbgE5kiTuJqwhoub3Cvrt81nZBwWf/l4FI1lk3x0EobgKs8fZu/7/LV
WRcgOpZBSbhPOdRHREOgca5b7YvRrDgCycns6GBAXh1+0XrOneteKv6lUD8zWIl3
aU0YlSqzJfRxtkXoAHjfZptoRDNFNgswnQV3ksi+leaFsXsrr/pUFSId6M1Y39JE
5nK2Ilac57Ch1nEm85DQACE23viatX5HGaojrQsqsIAeOss7n8/43FIUJ+QIpPQu
xyviNexccgA/sk4t1R87jSqo2+a/NJ+ePnmyoJi8cBu6VHlgC773X0LtXkjLOYKU
5mT4X5JvHelO3bITeUR5NZPAdnPaxpX2G3DVzRht0eOg/k5o1UkZCGP5NTFoj7Y5
XCKkh7TxBGzLdZmZJDlqrFFxnqgubYVxb/xCn/KgJIScOMmAmYA3CkYuczFwLNOB
1sfO8Bj8uMg0x9vXJz3l2wCdAA1lfTB3yKhCEjHIQmPd447gLwJQbqdU9w5O8vqL
GM4EdXtOyj0DgjFPUkclU1wn4No1cGwHzlVJZvr8TR1JiZBU/ZZ6BvMAa1t5MJNa
Gpaf+5w69TK1bVkOiYE2ucqMlkjgbPiWHn4nOqb4Wyc22dU2U7k4pri9QHNf0QZS
IwsSOslSoyTv3nV+obnBohJF9Zgc4aXN/7sKQwA3isKuVAoX7eQG4WTwV1xEcZub
57UhEh2PBMezqMk9D+dUc+EZjdP26Pc6aOKDNUtrXBh1WG88I0fXVlhpDkAgdtSE
h3TD6gcYiw+xtepi63lJNcP8nYYAOB6fiuQ+vrttqBFq3KMRjXwR5GIFRmi/Nbhx
ozeGC/NVp6M4zmK+EG9QDMEFiJ5Dsw+rv25o7BiYtgiVuszo0g96PBWsyxE0+Ktc
UP0srDUD0qR4qsXHhKlU4Ssh+yFEhVn5OHesHjDuYtF5Vg65pkmrXgqQmQ2npREW
uMHls/QVnLNtcw5fMf2pGj8rOBEGQ7gH6oPowHDInmatHLYH9vYv54Zgr4gp6V14
V6Db7ZfBh0Me7oRS6pMhLAwmZwpA9sY2ZYPrifrJWXFhcP1gufQ+9vMDoLg+xbOe
dH+Ub/oC/fgXo7/EZ6XBYLnhHE1egFL3hiGHWSQBrUX70cjhTt054W18xEeZSIgj
LvB6AX+oFWYN014/SHT0guKSmLpPgg5bbJ4Dlzpemb6zB1sBwxbFZfgDDzvDZPx3
PMjEoGuAI/ImciT3FsjuOgPObuOLYDlvM3vBma5+44mqdmSPRhdWHaRdTpVbVdeu
8lPRd39QdQJhHZHtl65/veGRdIiaKRwgTF/QAn4W85K+NEp+MXHBAeoBRkAKUgsR
n3UWmWyH2xAsbHrlndPkuITv0JFXplNVkvM4RRbuVOrmpN2AGW6XhmU9F5BLn/ls
c36eBUZmP0G2S9jCaje8amthZid/SnsXEhozgBM2PKzkFGmCRhOEpyaJs9EF1HAy
ORg3JmkLcATbkhkJUlSSLkSW1SJG3tI/doXIdJhtBiMtaXm9Pi6RLLKMXZ8gJfVL
sSIvrWqrrtLmpHH5dcomXwTfGhoZfgz5NvQ0MV1R3Vi0a+y/8koMTYyIO0sHKMqJ
cTw2bI4Gc23xZXA2PnLsmLz0cDbZ5ivFcnQcMRb4HUC/ViGDW+a7BoAeinlaUj1C
KN7FrrdeUBPPayEdD1JifXBis9oBwRb6dZcxYUc4KnUw8sfddA4mKzsGW12/FtOy
+6cLx6m0NoH7X/b2yw4p6UfvekPqhmS6qyhwP5emPtuZd3NgRSXy3Io1Sn16tsm5
lS0UGfWE+XB1zI7sn24EoaMoh4ukScTJF9yMJEiae4dZ8/0z7cv0blbWHXUv9Ib1
DVGnAMtxODSxz1SNHjCIKANpx1m0kEGXcZOTM18Llz3qNRlEM1CZl+Quu+p23wrl
tiUwBxJFWX76d2d8F/r9bOolswTIKQRMM7t2w4vLCh/zlWAK8SLIops/hb4itnOS
Q8uiRRnDBK1zUXFg90GmxXfBRCY6pSWwgOV8Ar/vkiwLwOgkhmTtAJu6GGKssqxr
OwZ85Kwck6UbrAxBoIQhiJXr7+6ER/X2jv4dtxpII8Ig/6bTzeAzJVIK8AG63u7+
CI84nDEmeaTfd7PnUK6Pr9ceceRz965dVFOIfGVtbiA4i2obAXxXERzzL+ztCPbS
HILUSs/qcIHEWMmbIAGiyYPdpTgFbCim6QIXqyf8y1MJooy7z+/wjnyC+YWjF71u
xv2dnxJCq0iFUXRSi/9yGOkLx6ZUdVeiP/e01H3BOodanwxV7Y8IVJGNOSMU1dYd
MmZ45cz0oBmXJ4b+tVgbcGwKKji280rTG9O3me9kHo/ebosfB2qE3TapEaWYf8lW
IyVUyUWZbUP4xsk86lN7A8oqVnCLIfSNB6cpaUAbd5xu/HRgdZed6Cm6xYlvAb2q
dVTY1iembHcGF2tpZzsP9C6TKCXG4LmFTcjFX40vTeBE5y93epCkrZU/CsJoibHz
cDZqez+hwzSL/yr3kEVLCuzZY6YDJ8j8eQEPu0YKZKBJF2uINgFiysQzDpCTHiNE
RVpArZnh6vjqcURJdrPvznNZwPh5wtWXtgSOPiMVdvuriGfjMu43XrGVOrQiof5u
WKT0/u4NAX50uOUPWd49lM1xPpR02ISkK5W0yQ8YmvX7xa4bpQSh+LExkDhmYb7j
12oNtJ+y7Ds+OvOVSoNlBlq6oeHnMxKFCGP4kaat9BPy7sFGMX5cShqGwpDUOBUS
erlZhN93lLMu+vEkhF6kPvD3w32eqpKHEIT44h9C/9Hk1GWFLjuRQGamF1bZsmFG
WN8ZSQ+dM1H7Ehl+C7Bi1jK3QpqlwFhStzw01DGrpbDnqaOZJRdze8iHhRHsr3QP
pYWoMtwd5iJ3wQivFrsKBa9l90huDSNghCnJJs1/WRkVigifeSNmdj7mW9VCsLUQ
M0fzbgFVp/wwwnBpzHF6YJM8vi1cHxV51TheiVyudxJqcKxxWNtggDQ7IyEyaHRr
PTILcb1hJJYoYYEIRP+k0SJBHYE8uJk3jTUbjO5gobtvVOK+SGI7cLsLr/G+Ay7t
3bOtHQ6RV1wSZaxSnVH9HrYnE/bVNPBbZ5J27OcuJIjmyYTb5y7VvKCpOXz8k6OM
NrT/zV/j0TBJpZtxVau0wLSx8PKmqhGEiLv6Ee65ZOcTotAZ8E84h60ZbJ7SCees
blRua5Q848LMAs4VlQsJPNCMXC2adhVzo5cj/kcOZEUYut4i3iy0X4sYmFyHyXHE
woKKOzFcaG68xX8jeCHOm3JeVCG0NnMuXDYmJApSNMkKfpoLOGKOBsAIY6xkCh9v
VgrO5PHGIGeUSXG2Q19uTit8xL1Eu6A3597ug+sednTL/UjeCl6aYIEDFhyLje8D
MdH7ZQAej5T5VYGKHbFVXr0Q+eJzetKIbyHVbDTp8IISNIR/s7t1k4Lq/2jpFecx
R84SuBwK3Z1VcCT8C2D4xBWz49z0uyFOcuQwnYn4QmT3dfCMbGcsQW8/UmZhz5KO
wRWGyxOQKqEUatClxumQqdfw2KU9CB6AOktGgUrSi2tNPY5XORBpBQeKCOLAmdye
U1AVbpe7KQml3uqZz/TPUTkxZZMS4x8k/HsBqODEw6xR3/gQMvtA+jPaINOuRPAk
PDdQixNR/s1Eg0UI7HByIcWlq3/n87QDmHnV5TFdblmro7gUxBwlAztxUrHsMvpo
79hF7xtyzM6FkUox/eyAlbVZxdJtBoW3vulzKs0xQitbKiaGv0GJXuX4XqJ6yhHi
JyreqdJO5+zC95ddLDlLGcmQw67bvH0r14oseuGeE5haQe5B/Woh5C2RW61ag4QY
utOs0Zr/CKQ88rxSbydTRAy3GrnvNqDA9siuPYcTLUgJpGWi502Dm0kluagrXhQt
BRo8vxzwGi/lUNqT9+xg78dU9ka9Fn8oNGjsiT0hhRsN8wPrQDsqhffiaWZ7K9yk
6MT0rMkGv693sOZPJPnqBDj1nGB9p+GRRrqJDSKQ3KriqMSdF+m9DmMn3B4XTjk3
RQa04Gepskav6OQiMC4KXEJl8e8cXDyPMN/b00L/B0oClnkWwjhkkp1QiCsMmzwP
8tk3yUalcITUUog5YduFXJl0LYF2YUEDIU6NBI2hEvMqBU+c1q1fzYybFRY7fh6y
tO3k48dinulzUzaqfE/+vCD+qy2x6YMT2Co0UrrtOnoARxNoOy878p9xWlWP3lD9
EK6KCx+IuxQvmIymh/1JSDKwYL+NbYtjr1gsZaviZioYs1aXVpPBMZMVPGZcdU5e
bXZRCXAaEO3yZBhsZ2fYINZHgDrexg12AjeQ4L+c00fbesN/UWudd/UwahmIoE05
D9uGRB5AqRzAc1ChyuW4WapJClBjVC6skh0KOUyq5vMnarNGhi/Nk7WxlzLvxkZ3
7oS+aAk6jUS7PX6PuagDkY92M88SrmXi31cqaUTY9teO+NtJpNixoR2Q7eybCtZp
oiaYfaWWEwnC0/wZ+Fpdxn2Jytu00iVcaGJ58BPROB8yidG7U3cPk/IIcsjXJtdF
vAKEK9Ggjvl0psCWpd+2ficSmflwvAWaahAejM/tyOT72iCYXsha89D4MIkeHlb6
5qL+DJkKFwmmYUOG6FzgPw+usKRDQd0ujvZxwhqpqJ9Hh3C3qQlP6OgRM55DR971
qLSk256Y9WO8Xhkg1FNQAYJzhbgQNDqalVAZ55/lyB6Fm09uFofCZ8f/F6ug3G2a
gpMUiHB9v82TZWyqzp8997YekWNLqJ0YLP0XfASVJW6H3mXSCgjfvZWbXX3YuMfR
+NaDneBTlXkE/RwJXZWHAwWdoCtKXAnKZmceq+5regWmuf/e+scU69MUyIoFmOmn
iwico3kztmxfL6OxtpJ0aq5pw/lwTHa16q1uNQ2H7MY75+28KZSzYLKO+pQpM2m7
1M0vPpYBGiK9XwTIgmBaClbMtmTfmpgwjNrslkl4mStCRulFPtghxlqoBW9Mdvsm
jVEfbBh2SW4Kg7Mov7SNEmjWov6QWxRqtTS/bzj7X+dVK7iT1iikv+LvABid5XyM
V0vRoLLqS4giqMsBYCtZ9Nf1MiViX09W14VuNg3RRF7gZyqvZGqNoPrWrf5aFOgo
QP3Kst700F3tWh4gMK3iolyqo9/D+3C3xzFCH0ta8gJiNd99332lTQF9dIXTnVX2
lPYMInbUzFMJ4jM5IM6OCOxIAffSEY/Ol6AdXZpBgllfT5zmzhxESACvDdwqP3Z8
7IdpEsWUtzJZ4JiOy1liHJkSmZczVzl2h+HiU72K3w6c1vK/mYdZzClcJF6h8abP
pNe4d8CqaSVRWQ7Mze/yggLRnEDJpfrhFNBirP5lB7Nu0GHGBBfB2NGOTlRU36J4
TiByopOD4/6pXZjGRQdu3D+MS8WgyhTMHJlcS9uHpoJVjXON5Ic54+ZTGOn2qZGT
abXtKbDYZ3hT/fOuf+HvpUP7zvPhyBdSpmQG0cxdGAAJ4+z8bEpbR8aETNN9EDnc
LQoHHeKibTUq4znPim8Mm4PDSEFJeFlsAplqHRf1E/eMVtye+sfgF2mnPolPga+Z
LYYXCgNo+29doDHw+Tjj+RdJtkZKAmmKWYobKRxFbXMSTeyrdtHuA5oVH5CyQP2K
gs15bvmU1/HitL8uEaMazt8Fwl9vnBjCUESQc42UFaRdaoJtVUH045WcuZJIriXA
8iuSzShz5Le9TnFUJWBetqXZHgAdY8txZPk5wIJfQQeMZ3XhlWQOSQa2FTGE/7Uj
uPnDtUziM0aOGA8wzjezGXepxa39D2w0FiETkKfLqcuOTMNZ5Th9vi/dcyOlTvzV
CZkrT8f6w4i4OeJ2nQMHkIdhXMXPrO3y9Uu6IkVshBBLSEceK5RTCopt6u3twNIe
sqGZXIuUXm2rcjjbnGiUfFe+AJIbYPco6JNBU+9essxnTDJR6J2IdZh3pH5XahzX
g/Ko7+D6/OG4Hi84ozRPEKkEPKK//nb121+cTadywypjPu11uD2sJnej0zhYqQO4
Iz2l/ufc32Ef9lb0f79Druy7efne10ipqnaPojT/1YqwcGHgLTAOYgKDBCMmXNe1
cRik4sOnTZLFGE1PLb+NiiieJohz/4gutPWgsfeXk+FY6yXTLI8yY8DprAPRbGsx
DLIxNIYALLacaxgQmS2fZBcjYlie2o8bd6xQ8JU6FiAwwD/X7R72tt6oZGDA7Xs+
ySAIVs6iV0fNWun45h0pymWLmK6TB1/Uri1tAX6uKlFKuz1tXzuAvAkWokjafz3q
aCOQeVmlZZa83ZWePE6RmN8aVaTN/a3WECkecFfoQTvXNOwFNMhn77ywgw9tpoNG
nQsvzYxD4WMuuAiDwkeV7ag7bw50lUYJdCB3pEMZUjChfdMGVS0ONP6uLIBqaA50
yZ0Q+I0Kdsk5Pov2c1IkT0TOH29g4OZRq+wihDz3wAXa8d8KfpXjtr2CquNKFZfi
kJgPdmSHQ5t4VmWfhFST6PK4BYsfqzthGShc+fRopeQdW/HNnwFXz9uNbINzBVep
lORUlq0ndSuiAaDhh7ehybwgRFMIt2Ou2Z6IbLhNhHOEnggNk52gc1nGYJO4C8NN
im0WSFdjy1/Pi+rWSGdjAZSW9jFvCQQe8HPgmO1N/LRSegCBE5e+iI5hE+CtZu0P
3OrtI3oOtTznYqcXrOW+f3ncx22yhwMX+lUTLooD2OSJHVa9rk8CZHbqTnWIgf66
6W2fGY/y85L9Yk/mnGjkXyO10SGrlPWuPcFKgo3N4CByLSv4xYuE8N75Rn2CdLi+
l/yaIGIsMOd51wHkuvGQlGhOyCMZtuaLd+hbjkOnP3umWlozg+90gj7BGkr9FgvD
Nt6tFYrzbTpfzYEasK70bfUScVOYQ737VifD8b9U1IEq7grYSouJSgf5uFQBwMp6
KwuXPyptSJgXl62uEYIvhLIptiZpmocWfSIV0BMKDuqBrrB9cl5eoWba7OVTgZ3j
jJ0la/XAWcTh+iArEyFZ64FTGoCju3UF8motthl8rG4czc+jffJRsYGerwjh8U6D
fEmJy8rUhbcHU/iRHOmJoVzAkMzzYxnuvVG07zBOeNUi4cLRTY5Y7fFf3czlHCd/
2nB49XQTmINAJmwcf6R9DV0ETBSp9qEvfZYoL+CwL3BSThivFDkp+WAKgFZGOZSN
eYKRVTpZiiFyWsIUTwwPKDyDt8eJ/Gp6WU4xp2Gt9LHu3vIX6ayfdDz+rsbT7cp4
x3geHy1U9XiUyzvZkq6mGQAGdFuodOc925Z9JOc1mnpZ4XNo6sJ1UOd3Vw3viIWu
eL7EVYXTYQM5o89FRzN3bgP/rSoFgO+GdTJNbERvaQm9rd3a0VEg1RNfgfLXSNsw
neYJmcyZgufTwfn0RmBH/d7MPYjK3Lj/nL4boWiiRYDWwhExDOmRE2SFnUTNnqIh
rwP447ehr+eVNmaKljHicA5T3YrWAS046DbeVUkz5mwgB+mbhVk3FhkfpHJ8DrWB
bi0rOsXrm1hRQaleRz4DYBk9PE9DxeD0+n5KR2VzuVX+Y/M5ZJCx7gHvuNGplB+S
+fzx35eaDeTkh2UO11k4fMpWzshnZ3Q90ixh/wWzSUGd1ZvhdEvPOX9twnQtByQb
5E5dEL8gIiES2/0BfUrELtpvA2/m8yNph+sKQrU7h9pKkvIwlDiyhncRg8AYj7wT
0isnRO+mNPalC+a7/0sKTmVOxLM4JBR4V07XtsEoi5+fYG4ttUo2zMtpLxiFceT0
vbgpoC+JgjXxj2VTT+8hkzvUeMzeTTRgTG17xeIz137a6JrKWkXkf6eFod2lij94
0gVGQ0YD8Phc4Nle1ZtGbE9CFc5cO2XwKweKNioKcOPbX90JjHTxi8dbZ9FEl2iN
ZcBZVo+Src9YCx3mnm/bOAFl3Ebn7Ble/uwlwXVw0q2hg/I9moo0UjHfbdJpmaH/
vHWctWr+FU0rshe+xD1g6jcSOXBlO+kyFKQQpyGq4NrMJrUXgR87pTKL+8RYv2OW
aJA4YbFN/eIMOrMgRPgvrrxjdD8HzElOr/uMIHPLJQTkc2bWVg1llSHfMG0uyY9w
S3l8BGGt8/pt6sQCXqccosEcEXSpDtshta2D5Dzllf2ERgNQHkGv+hYptL7DkPRq
HGeu1Pr9c3X7u477UenTngPBoobvwTmCgZGrHlrXV4etm0Lv+0wOa3WFjJ2s0/NJ
xPZ95KULsh1uce0JhmOcEPuf2J/c25fkbkBtDIvjD0PAdyZeOEZX1fSu+V/UnqBd
D2oX1PFHxoHllotcMDn1pTXFYPK+BeK7rawqD5XCU4boHisZqAr9uSjdXiItOC+7
eeDQCDcMSzobFABHfWDAAS29eGyTRFE5kiCzE474qbFDICBwPpsL5tIsghqdO0ow
IvtgS5T8WbOpvR5hUQb1RKhZG8/ht6477YEtOm+tZDMlT6SuZKVT1MKg9sOzZoHr
YDI5YfSrfCHA7HaOTZBpmW9BxV6GRFKthVXeldmaBErIwMVuGVl39FVQicCdxLPa
x87BBijSKzxbrfukaPJdIjfS/2O3D7rBYEGVzzgEl7S7jVXhWOoq9mcjhcMcyXzw
PVUEqC2DWOcmA/tGND4bFGmdiR8UkA5dGTiQwxscapDv8UQroSkRUzpjCL0M3EIB
sk6UTvOojqCKqFAojnqJdyYEd+IJje40Ds5INtpCH2KkcP9PnyqiFagJqQHpZ3HZ
3n4vdfYZQK9opAgwP/1R78tjRti58kFDXPg50gH77hj8F2lA42laMg9W/mglI9Y3
TsAwO3NtaqP4D/sWbRrvEemOKfJkXVuidEGaj0Vd98XWtZi4MDkGJTmdk/C9qVDZ
CSfoHLtKdneTaF+HUmcY8Y3fhh/N+WP/z9zANgeZojSAiS/JRzgzE8SHPIP7BFZ7
mIVm058TATapzwaeW3wnj4fOu4GIpXnVbyehc05AVmjE7EBzyHnHZOjwt223tspY
MVm8IsRzwIm2YDQ8yStqb35dujiuIqEpVhyTsrz8ny8brysxCsS6OIlqAvYQ3Qbx
nRiAcGKkm5F4SJ0eTpB83IJ80nIhoQUhIgy1YmXKx2lfvVnwqgyBqNG1CRb04sfg
SZWhCNSDQKLcGTWLUrIUKX5ZYU13VKmwCog5Mbf1gWjXKHfhKbFMcA2i+R3E221C
D9CYWCqskXDgJk1fjkcxgq6T46fPF068dyTghHYDcgZqnXfOID6LY1ATUSMWIywP
Vh9Kc0dlfZUF4TUGbrLpGWpCpk4UV5ilsIza9nvHTN26iCZKtbcBRQj9SyW6E311
0JOGwHKg+CjLCOwdlCP98NYAkt4yuRbrPzBeC6kkUYW4vEpV8mTftSqiPGiS27MR
kEPPYK8cgXGgDRQcr03SsmdNcGidg0jcFUTXs485usWinl7mw7NUVCrMpFqv9RFX
Fh1VAaqUeIY0C1N62CVrL8oDNAkXX8jFVzu6Ymne5E5YcEZZDJP92ixUmIJXRkon
LQPtGJDQGDZ+leuHBVBQ9oPzTX8gsM3nTDJwA1cNnHXfqjM/w5bdV4bBZUSeMYhw
XyBHO5F7eEx41+U8seGi1fa3RBZCSGLlzPI0pUlGHfmSWzWgNTEdY14Yot98iflW
gWLsQmaVEnYa1uq1XH0lirJxpA9VQ0sIocQ4ev8fcasSTuWJzHWdevPI8bGP2T2C
NKeIvTssRtO/pLmMuQ3vLs8LSG0EeAIgM/pFEFnbNnAchjctMqI+sSc9Zl43UvBm
qFIEBLSTn1bX29jfLHPFtWVM0rCyAS5vjlR5FqLoJSnHNaEPxkwgMFM8HQp5TFE7
TqeQKU6fpVARidSf/7axizmVOVdMEtyhjUYBtJjAw5haTfnNScY8e8giosZNnb8/
jy2Kvs18fCMevB03vguZV6HdXxt+yMX/eY0udsbdEZw2B2UtUlsgxQ35VAciaRhB
2+44D+bpdPBcEemLipR57PLgkBQhKIGKpQ4DU/TEj0b5ZyztH4c8ZE8GqzkC9oUY
nFslJm9Gzt8/t+/6Pmt+PUcoT1xWg1UNjii+EoSaLafFBcYQPxj4Hiee35Ffhefq
pkncdBrunSMdgYV6sKcyiXfLqPX/2n6Ord9KsFiZnAD/K7zJC9T3qg0I0CVK+JRy
8JOA2P5v7ylxx8dieY/kp38yy8GzeatnDMCkT/tXuD6xzpQjNAAt/D1JrStcxyCi
jZkGz0KJPJwAHNuz0KUp6oUseERLIEiUqOta2RyQXbSHAeC9ua/fkkD5C3jghysU
eAVxhBgE6Ewz2I7QIpZ8Pmv0Wr173pEPKAeJd7p5cylWJcA9585dgYNMFSGjXyHz
Pixo94LnZ/rC16V5An6dOgc58RTr50HIfaF1uFpgDvNMhv0HMhtUdWSHCZJzLy8Y
6cLgHjFNU5K1qs5B2qf1HNIgvzuLKbjJ5XinGEha2+vk6AXtCQZl0cuGAJWYdfYS
Le8nLvBtDbGFk/+s3N2SIhBdQQFvBu26IAU1JsFj4hndrd290dIsfswFjG4jSQNC
t7FPcsHS1hUzUgDBn76sE7Wxf8nWbkmuSVUHvMZe9p4Mj6vWugUH3DGGBDLdo2tg
sHsQHLvJ3Ra+At8F9rv6gTMsziipcLjGYcCJC7oA9/Mtc+RJTjQRQ9WCRuOdyv38
3x19ygM2kzhlOooDf0WZkMR85kkxIhh4k559mI5X+7uNebCXlLKRpyFJx4vtciWS
33VYtBTzI3fTffFVYgHJHjdUHtgwTfnnkI+D0u9v22FYgzWloIseWEZHQsMJtgd1
bPhrh9TrIa1dACNXojyqbTzPoQf4yf46NxuJGw7kt7SNgil9nYQ/5WjTrn5daEWv
qxMCpK81AkUo8LgSftbrDKyjsP24ttwR/wNThH5ILEyNjkT53lU/VVW38zY0+nVh
BD3NhxyE4BL1jZ7NAmdglQjgWgYLlWWjxeJGfm2Jrub4HVG+zBrgVIf0GkvSLubW
9r8BaOVtLF47gBAKPGATWcX8I78bo7tAtwgnGcj0iJTvoAMW89W5E27ES9k3JBnq
RN105o6XdbJffvMjJz1fL4cf1TWHZQoI/q21pDe4zdm4rHFyV7CGna8N0xVzRKYW
bUCIvq6H9m5bTCQW/T4NmnX+TTN225k3gtcDAZjXNppVfFoir/0YCr6jzNngdZeJ
TuE3v2N0Wvw//mebYU5oNdrQuSCCLNGScy5AIpDSbBzr0BNcJnmsXY6lyogMWm9x
FNKhrsnnqHberHruPUqN3uGXr037Hi5Gy+SIC5LsLdvGGnO+bGcRaFzW8vp835CF
mnkG6z+sM6+Le+QQbEm94BmE+QsSvTBwOpgU2r68Y9+kyZ5Wsgmy86osZMKY03+F
M94Dn+iZ/P4TCTg5SoXZxy9vFSCmJbtcbdHB/OejxUBibwbtlFA1txcatRwyRWeO
rjydKEbC4+l8E4GN0XonqSGDq7rvtOxrGG25nvgIp6EQayXySgOD+euLU+Gtlkft
wHYFRigH4IQwPen/rwHVNcM1e0FWTlnJfk7fq688yRRIXpaihu/EeeNY8Zja1kn8
Gb/HcDcvitpFfAlO4FHwK1DKYepXeRe69ofR3l50lnlBxeQJdoodrmyz6gfcjcxd
6DLYlChgltZhbbssbZpx+lm9/+R4xfhJr011uY9xZF80i2DrkAx6ayaE2/QQJgLU
WRgGjE+GhwAa76ClnMq/eg4lsJ/EqDO9VCLcVx1QmnKSxpBxDvFOaXY5NknTiMPP
vE9Omw39/jHISC7I5Zo/OvoMSg+GAbc9z8UdXVOKZDFNJxjhokBh0GnusP4lDw4u
GYoIAoRMDn8BQlkG+YiYr0tPfIvBin1MptfDyXy613x9xX8xmGzYDR2yUPBuJcvV
Qgcku/vwKW8CmHuy6GartmwxpoUZo/+XP6x7G9xLiCMuADA/i0mM2glhXjZBKRls
GmeQbd6RSeYI3P2QTW2oFrkaeOL/6t+RH6a7hngUVkl0EFmk1UryDK3dxeruLzLm
hM5hgaWNq8B12S89xUiWCDEe9JXtS9LN8AodZG+zylwV4+XbxMH7rswip91VaJOE
Qz4JAIAnjtp/rLbFI7ujxRNSpCSEFuujnWt7RC7gnbLv3hGSGisGLdxGD9j/Lzqs
L9325U2UCwe9SAcdSveFslTn71KYfmWZP9c1kXO+CFUiJ7nawFt65DrD37nEPegQ
bg6SISk01mp4s1VoMoxZLKNr5FTnV1N29fl0CJPlVvp/5K0DAxQ5M8FawtcyMaJo
8srmq7cK/voyTlv5ua/6nnXuNRzvAhfULjiA69C3AxnycvpnEFHQBsXHPIz+x2B3
clj7GBTwANTwV9sI0HJ2WDKLaWYsvEB60oweSwRGdNHLeZMauVIKc84LMx65L46f
qGtYK9I/PigrD7WEK+poSfVb05j8CvKecBfnRx3SwetqysYzhCrSd/8KuTKkzZIM
lJ+/WMSNmW7W4+FRw1TBTyA/kd0xI+x5FeTRkSVomCD+BxYk3RjNTTYKzpEI2Rvt
Eg8Lj3QgnfBFumJQfcr0/JNCpYtu2+x3iWzvgNdt6lNDZAE6y9I0aeXBzUOkMTZp
/yKjg3o2nvLgQY6aL6UbbnXkMGzIZGbCGH0TBpr3Qd6j0/ecHJdyTrqjsMmzfIo+
tGopNW3VWIpf8HX10nPOQIa8i5hlQa4ax6XJU5W8Ld0gw+abnOJsVFodiJNQjDPN
E03qmSW1ELgXU0c3ZlQeBnZ/pzmrtJb4mZDUq2dllN/y/gpvOaqbD3l31cwYsWvM
exHX/rJqOhLatgjggIznBFAW5DR19EoJ1BEX0Ad8dmK5hjPaiBn7O/mL30jcxjs6
k4PLpvSwT5A4ZnyuJTDVw49fSJUwFDGIWzY5V/Sz9AR+rIpHp65wYvshuyWxGU55
UD5RdFwO0jWOXJn8havj8hoZUcw83mpMFREqfbmzxB/aYZMCfgiIwBXnJ7yDmwhz
s1EJFilsVI7042+uSkdgAF6alDUtfmQIK88Q39BzdkT1g/LB9K9pdim3xfusz5PD
ARq49kubwZu61i5KioxCDpXSiDKNPmdfuvR+FL4EE2c7ImlhdDdhLnzGG9X7EL/3
hAhG4xwxrbkqNYXEIJGkC0ID5H80YfYLaFPKzDMFmAsDzO4Xc1JQFgUWcTMkGIo5
I+tLJN/F+yxQdfkbF60wPjYlGSyDzL5BwPq910FjAwoUFLxHHMsSGFvfrZIuTr5D
sW0VI5AOHcTfxX/cUOlq+Y4IYAPw1ndmMc4n6I4KV8kw8QT4APN42kduhiPh0n4L
BmCgVU7SA1Dw9L8GeNz5PCA7iBaaGBixwdrXxJjLFjWeH/EWMBHFm3Ss5XxBapg9
cSE4TCe/2UVWqKPb3BUUAIT1h6V1gIH07DCLbS7rpYlguSi+BLSWDJtrfbZbvl28
Sn5NUpTOyMxPp/wkjIpbamBZQOmThtT8tOvzP1ur8zkqqJS+NmVhgynMaVI5zz7q
ryOjhkWoffzjvt7uRWQF8k76h3mjLdAqkYvJb9HjJUGPQf+c2S/3eF5PX3nz+2c+
tVPU0mCUvh8/zE/WoM8jzpEQfzDqppYlaQxCeDD5rph+5vNVbVedWoPZFp0jTtsS
OWVIlweNRPSxQy+DqErLBIdGnBQTDmp+s6k9jNuPP21M1Fd69tByjL/g8wZ93GkE
NLd/mxwjJRKfrnV8mGsECqAIMT/mPZFRIhE23GnjEMVm0xlv+Cey9l+sOS/QT8MY
Ap8v4D9HcGpqOHN3dxZwvZGFCjh9bud3LNJeu4BTK5RKvvLYfbLPy9QvWhiIB6HL
HPHMGVlvhnIPu1HvA0ikkQJDhDKduWPA0mTdJbQ09Qo2aBBKxlDXs28JLBdRNs6U
FMbmpUvR2JkJf4dEpUuPVXpX5drGQA4ID+RJkv+qmFSQil6TNZuhjl5z9mitJTsV
bQEaXsuP/7+Ce9q/mGBXFsX9sbuyKqHHp1FIoN5stzJyM8ZERvbAihHJyn+0+23P
uZ3TkJQVJvaeEroM+IR6WhOaXg2TQwh6JTLhixnmTxKWGE3Bg/txcOpXgsmApYgc
YLaLAftSvuRVbu3q6Q1CAeyxqIRGflfj0ydzE1IRQdcRRB4/LQItFNlDMluc5BDi
5+0eqsH7EHm/Yl/JoFiXc86NbaAKFXT1mJuD49haSDQcg9LjEOkDhko2pQpmGbFG
XVqX3HhFgej898HOCBFdcotR38pVvywBeR5Gusyo+W5/T8T8jnrk5lponEa8r8rD
kl2sZ4xTacK4a228C+ywAlDrc+YAqx6KHNc9wKSIlF4Qeb/WKRkOIT49xnp7FoLU
Ur9bJTTnbOZeR+71bQWPAU0IWDmIj5rlNwB9Jdpi+6isA6/mI837Djj+H69vSHHg
kJIxCMnypAxNwl2QFMWqqnetIS3z/H7+8aHGgkx0hyRGSptcZGpZJ2RlaxM6r+/N
oSo5CAMfr2oOUXHBLjiKZr+dl0E0P1IA7bf6/cpIk/ykfbxw+X+pIk1A2jPJA+zE
h4EBwwybSY2c90wtPBqaSJtohL8WYiT3MoNE86nuDal9SwL+DJ3I7/JaEbi59U0l
rstuHvCkXewvxXLe4EEfzjCPHLzDH1mNPqKmiAzc2RMzVDyRduhxxZJHGHOdw3YV
xEhAwXdEYxqTvLh4zy0SO3sBDktyiMHzTrmujtQaMmSs21cyAoFw26UKHqNfZGN7
dy4tmxWFxdVtMH+d4YVmRYGRWuFKxLheUK5x7tl7XQk9PdansUGgFHXGuFQdRtLS
mu+Ik0Siqt6ZLjZ5LXZoyWMQWGKFNyED74dKdYnm+rAFTt8Xidu+amxwPDsTb9T2
sKvIh3AKDxtsmcr7WmKEXqAgGQ0eIP/fOnG4MTQwACZFLsyRsJi4jSzE1/szpuYD
YwivfXQFsPnBFCYm84QgSLuzeZ5eoEWdqVKaUbvr62E94aCmxZEZcYxtG2Jj5rF0
rq/JkmDuJovvHjI9OK1iKvRUU/hNDcH/OrgOe+wqLHOpgm6Rs6sqaW3OH8NNqx30
B5IZ9A5E7wOGgE3035Sx0womBZoptPbVYketgZMqrUKx3Q1e3mMV1z+eEOaJT7M0
W1dYvLU2/bkvMt26Z1dgHQxMArwnlk6ZOFVd+t5ShW+kXUaImSTXYZ8u39g/2aWQ
Wqhlaf9EI1gJJK4zubssfyYNbT1am7w0R1rC4ymPfVNgr0smJ8bGoaAPx81vMspa
q0rdjnG0xWbAco8FidQM6VWg4KiMwSOD8IEM39Q2eDG+hG9p7jkrE7HA3zbOgE0R
+DCFkgbKZKrw2noYSymU1TtD1pZ692VoznxCPObpVYItfPVlP0RNxQ11Cd+4S28j
SZONg6I/GJ0ohcDkP/0LKomOPYDFtSaTWEjGyoln6Hy+ZtPG/HT6TOLnWgcmA1qA
AOIyPrwFsZ0I8vhc6xLU7DljYyZRmiE2ksZuBHHPw53zLsCKc4GQ04veW3rY6Cd1
rMcoMBEb37hkCxQzEI8QMMJrSH23ZIS5eJE7acQH1QJjBNTG0VcHfAr3xkSLn0RL
VuowakVaiUuK14927uPiGkP7tR6A6NQAZZPVakjsGZVVJB3C+xYBxv2M9b5TXBsB
wfz77tscHaUiOU7I+B1gyxCncNY1lcS6fQ4Pwmwu/qhoFh0cmZybd3pLa7YgAn1u
7UDCKSnKjGoeWyNZuxyRLryPV+U16AiWFImKK0E8ve44WU3QxRTMqn28+Be+Y7lm
kPSULLDiWaOWav107iUWVxcLqgoMhYIW18IheXMlRIdOXzI6cdqBEXM4k+PwkBT2
K3dUZQfut0dBaZbibjTdI35odTTxbkdRIRH89jfvez9pUDgdtprQ1m5WbM0hzdEa
Oo54MGzZOSOOBb76sPqBwvTDBYo/8pF/S6au7h81XQcAEZm6YigK6C1wtciBOlQR
rowfxpF9xsNnUJKYnzVxIUvmV4tfgZcuOWLZW281DGyGfEg35t+C07AR16aAw81U
FDALBTD2j3ilSs7ajDSwZJfe48r9+kz4o0IyibkXY3gjq+j4VIcqyGk//+/kWc5L
/Tbn9BuNAnVPe/UXGUgmGLLgIj9+A/p93Im01FqbmytHD6lfXhRlHOidaIX07/7q
cVfQCuZDsz0VyolxX3pURU+gYL9m3kd7qPapIgZ3tqKjoE5ValhhHiO5ClCSCfdP
vUMrU6XQqjhYgg10t3xGWUS8krYW17qQKPyKPUKUK9R/WBC1RqGUegjtf0vhKmv3
XO4VpVAmokHJc0u5sgD2XWJznuTmAiF8O4ZZX5EXx0nlGEZJmILwpRmZd68JVF4/
az/mG4oaRd5aM52aOod8Pq6UQHGtmVQGl66PTc9//JXGmNXmXNGzbw1N/1DJo3Rn
qz4fV9yGFragzbd7LT8qVxR69xGEHFuG/QKEkDUpqBOQPoRkHR1qtcbmv0zrpxlv
he8lFioQp6Q2WUtkWn9a0vpJsHOvE3X3obWwA52wnhvx4aWpFp5ZG6/VeN8+FBZJ
NeakYxd/zjlVSkXmuji5te+WC/w9MHQHCU3tp+XzCPi5iLocxR83yCHO6UBOO2Xq
Yfb9YIFmaGNUHf5sOb8OClij5twsFysvyrZHcZS+tvHOl06nc9kQ0lJVCp3s8VOF
0cJRIUrd6Cr4gkrYSoMvZzpOsvD4gK2vb3LKNYnM5Iq+Vj+RqWu4JFiWmdIDWsyW
qysiJY1+I71ea+9hGqnC8XHbrL/gI7ne33Kb4jDf8lPodZ+5MCYe+xVMyd8n4/Ht
F3fLggDZR4+N9ggcsYXEDTkRg71HVe/OqY2ncbFeo/OssmKMDR1HkbAynJXUywaF
otiw00iTICBeToIbIMleVCB73pTGWgMGjOi2WTIW7Ekr8TOjvG8CuljCP4dTaiBc
YNmu9DJBux6C9jtH0meHDoTfIub9KJVxKOm4rpNrZ2W5wFG6VLj/UtFrKd9vvDqo
7LiW5RChhzB8pjVysPAcUFUwWmWMn12Csnxgi93acME3KyfgKOvpwAA5ZaNQwRJk
cD02n5yCQbQFJUlsMIMLFgJRW1OcvmtF6kChS7EB43RsgoNdY9w1BmoPLQ/gEFhU
EvMXW0yjYaKCrgcPhukXm3vVw5Wa7qHzq0acMPeNe0K00UFnnd5cKkTR8TMAJGLJ
bojkPjknMmlQReUVqH2nuOFhhiKWkWM8Ysunk11RbOZ3Zw6tRz6y4PT8/RQGq04g
X7leSj2W6LOdmK759lgZJ/l2NzdRLOwa9jj5tveP5eVYkJAu6sBGcVfd+4YwCJEU
m/MimXFcLZef+G/sZ4tfs9kJzWzpcs5il9MfWcMRPDksFOnaR6929hTI2luSPX/z
ssKChHmKJd/4xTFuDYDhsB2FWWXPCxg5vwH8JMi6qTkM+f8SsBvHij4OY9+iqlQh
YeOP1XY9eJvpKkPHgqo5PhCPtzmaHEMpwdaAGljCufxh/jiXBFt7gfSD8sK48OTB
vs3oxFsYwCcteumb1sLOUIxT28OI+OTi/VCongIp/39cat4qwWLSYwz4RSWsumDC
AH+YS5bmVWFKYhZAi1kWxIQw04upHkGbsWYJDfkIgFg36EmtNy6qIifAw3MkrehD
OyfJKX9gNY4mab5jWxexPTf2CSd8PCPdRh2k+DSJce0MtbNIG2AD+2FffU4hkE1A
BKV+TpOV1oWKvYAdzRZSkmVnNX3PKzYYwybr3WFKxqQVv6P40s51TCPrwgIpBtys
Z9ArQAji9ING+Cs7bBWldyZdOT+ZuCrAVLe33Hn3GRrTY+JEz1ABSdly8fadauyv
ENWeZ93kkKEgrpL1roM6MVAKvtUhxB8IviokqdxPBaaEM4D9k+MS9NkgoBjWDBzw
spvcd/4EUVfHURCtFyjndomDrMG9qk+ZTD5lH6xjLBYOSIbxqxQuytuN4lvVcc5i
6mYF+pxc2aZXdzbLtdntG1mKaEMddlrYXhtoA2GjuAhlkY1CBf7gveFo411E2CVz
XlefoHikI1S7rGOGiMDynVV63Gp+I19UFnQh5WNJLRrrBn01mm3w87bGhpLQmwfM
F8vdIala2NoSBoAGR5QXd8n6wAw1h8q3/avPbjR/Ky1fdyicCz45V8ehdYFfpeMs
V67O/lufyAPKm+AyhTXZYK3/EesYzoCyGX8+AIHshZeI2EIEHNjUvKsur0XFDc7b
+MoF28IB8sZnPTxPG0nRnIhqLJhllOnHR/9VeTX4jcfunsk6qfjYFk229CTZUN6g
kGKkd+1VLW0CNKOYPax4Qy5XzDO0lfRNZOFOpXNJWq5OeW1eakMWTS0HMzA9p/4C
buZ5yxx1lDbHSb5oOlLrunIEix0X3lBwwjVF+CB/cDTh7BKl1hSKlkfc1AbgKizZ
F6XoNjV1l+4toZDNzjtWP7cLhneKQxzx7OQdIWM+Me78MKtLuSWR6/HtzAaprNYs
5lOBLbY5fiOSo+t8PY87fy7WTb1JyXf6bbmPQrl7CpkIvv0r0GHd/FSMArFwB1O4
ktwdtJ6f7HZKLp6VdzInvwxtIVx3afQyCivSZpGUtUuZe9+DOUuYzt6+YY4Pqsmb
XJ9rGGFlSzyV1WBLE49CQqkWR5pY6Kuk2ZVqJiVwUJKmfcj6q1uz9WCUbCW9BOaH
ua5UCk0ikhqvN2hYVPjnf5d6bImxY85qDp6U6LO0s13xPDfQLkPHMkahQRateV0D
nQR0OSdfhJPdCAmbphYthNcW+kquvLc6d6m6tn4ZUM6hH1LGm6yirHmwy25HRLgH
7pZ1t3OiF7nnvF7QZS1hYEPFr3oYUiU+NBRwuq+GCN5X7Br3paj0yZKNv8TucqTb
p3HREFryj/u5F7/n1k2Vls1L07bRwQeCJPNFxwAHi9QjPlBSIus7bbDsjl6zhIi+
GCC4mzIPLHdgvkrZ1Hb4LNBjo8wOMpR7D/hGlHpIeiedZy4etV0tY1HblZMZ36P/
qaJoMVcgqPCHNF+eP3aaTYauMKzSIRgwcMd0b+NDzRfGvk3uUl71l8CnXAQzdMB7
9tyypikhVCUxBEF4BtftQhzsm1ET1B7zJOwHBxQJYLxaIqrX/h13gFC8JIxp/Cgg
7sKVGh388Ewoem/UIBl5FzfhDNcOeTJblRUmBiQnBxjZffzj50eSMptriRV/gYGd
u3DJ3hWKQm8rkwyNnTSLt8ALwQpNlaSayUOMkUlLAVBb3QtQHcsuehT0IPOJw0cR
+RrOVolWTAyaTDhKG8OXZtTTcxS7mE6OBS/ygK+BXKTX06srjIptPULcLjCsIksV
R87RuveNUHWxXLUK3sg5m9FK90GZ60BpNyyV9PDEWna2MyfxRn3Demx93L/PYkYT
QTgpCdGbdN+aV9A2Ya+60HA8FhbyDKRzG0ONURmIAnlX5TwyHb/AhTfo7u0lOFHp
B2mcgvadAPT/X/weAVElTxZoZw5TyX68yZysRCiCC49Ri9uHvsFs2m4uB1Q81kKp
RY4Q0P9JpCefDvd35U513ZwRxlnBnQ1oEEpQnt8EZ+GxoROnu3Al+V4osQDbS6Fd
uhE89+2NgeOewWjC8EHZ1mKlhKnoT8BJvVxbBttZqFu/jVAdHX7ObDAyktWVaZFZ
ZW5r1PdH/1T5V3cx2YBO1kjUVJXdH7OXShpgKbM3lbZpD0ccCGGf5jt+6EhS6cK3
m3yBAbYxeBWwwAafkcLIXcvNDPwBa8V6SDEcR6rlzoe+7CBaJS5OHx7MNvmXLVBI
nRN3t+bODJ3oDMQVMCFH1l5YG5WU3OZRZdu0afTruUCcs7yYVJFm79ebq69XOwuO
roI5lePNIJviZhmb/yaoVNovCwfLepRoswet9qASXmKCy/iWSCE8Ne6cYmMSd4ba
wJ9t7L03xjcn2uOPK2b4us2JvMj1lAYVB2KA850QtvFf4sioyq4brFwIsHN7Qzky
peTFnpzu4QAZNbcr54fUcliqV3YnKNlBAsz9C069UFh+MO4pKV+AnJblwyEI+rJz
AP00pepl/OSbD2LrbRciuQMfd+g26ECauEhGsqj6b2jA/Q9eaYW4lH3HQEXiWJtS
9wVv2SHcWiW7Fj9MLi1MY4pzEeJEU1XNO759xwwSvtm948TsXGn5TUyZOQIrx6BN
aX0GYtydtsxBe0v356ud4FYVMnHsncWnzvsl5woe4NamBazfO2rzn6UtWmRVKby8
rAka1VWjeQP2Sdu6V/RawAfy/Sd3oG7Fe+L6GxM2vpsQIJn6F/EuLm0cVNzCEzk3
zJzu1B2PKb2/msARzs04PbKwPIIA2IhneuTv19Bx/6Zt+qgQ303oSmdMdmlxLCwT
asb+guiTq5g2NNgxtnRGvlNljaNomQcTxX3+Okz0Ks4F8fLDbDPPgEPBpGB7bAJ5
ILkNrEdSqFVe0/Lm2jxSN/qPHyNbUqr3wBZVOB8eGRmMtnP5OU4Om1OLhTiUPlvq
hkgy4bMgZY3PTYjJdBwoKuz7zaxYMZqSHC5dGLTbHdGxFpX469BvZuymatGYdWcj
dFfrwbw4nyw/rmxrg3hZxr+ajqezo4uylZDa1+8ly5ErNXTJzbhCtyyvv7hF23jV
nE6FqsXvuWQ0GZUbKGCMCAgKbCwuMDtGZOITUoh1qwocwjJIOwORLSj2xWGU1qTn
C98OVxPp+ajub6P3L7C/DxFIm8Mj1yI2N35lMYPPpuVDgiBaZKNmNvBEn0i3e4rI
DgQGAng5L92wEFPVMqYfz9u/J+ThmW8qri2GVf1PHNxyC7d3LuW0ycDWSb/D2xm+
hEo3rWxMAZOgQUXqwzOQDE4/hIW0A9P8SJ5UWmXLm7+gSo6/8Zb1ZjdHPT0mVwlb
Z3Hd4paGPYZhmNru8Lz9/mViJDAnNmL3sGeGY4394VgioqClM58UXBzwkVlwk8qL
cfvqFw4HUGqu8KcMG5P+XTPtKvYrfMhfkoXnKkyypTQ6HxUzvyXyn22iHO06wFHX
h8L24uXX7bpdo4NwIm1pNjo5kV2RUyAZFr4TMKs9EpHDKTxJ5UoR5ak3Q4UNEJkq
VMOImUYV1fEdCOl9ihoW1g6toYtaNWjJRpnU4SXSgHub8zW2B9rI6RRfMlaHsO52
PINyjDZix0V+hi2pLHAnO2EPttBRe2dhhxEshSvq4FeaO4hDGzIb5prsQtW94q2r
5agZhkHfwpLlolYq6XG52iH8ircmX1okkcJG8Wq04sPJD+pFUp+qF338q0y+iRar
yUE2R9+4HpSPnEjRX1BrmOAohDVpYOoIQMeIlcmxtStQqSZOPW4w5UwkEx+eGCt/
yraHrMLKsNXBeQfAD9UOD0o8C73RuPMWs7YRrediqrHS7H1lOf4YPmcsGKcDZQpH
bO99pKVin7O30eG4U3gOyydF8PUkqQMjNuhA/I2Mz2LY7b3i3n1PgbLw9LoTkFsT
Be4bKVbUTatQoqW6NS1NF6KVGal9je8mlW+fgQ4bRq7u65i2sd0kAu89JYfX7WBH
51TMBnogSojMX2QHTD+Yi7gm31FP7nEAv0nKd7ZmOYP0zHGF59aZmJS2gwgsmvvm
PBjNKw9Lv8eCYLk2GGcqqpRLFltJNrPjXUZq9FEijzl6B+mzkdK2gt6sK9RpCbvQ
/TOdO8tmtFNq5yqRiu3+xAMX2JCNtKXuNzgau9vc99F9ivyEj2NStULcjrVSOht7
0pNcMY2SLOzhJ3qq1NWDpxdPZ+sD1lekY88a6M4r9kqDQ2weRtaHcPtbdv9BLMZk
fyCApGx3F/ky+KoS0qj3YlKxTzhGQFjBh13GZA/Tl0Vs/TZ4Ky4BRnHDFvMhQbZ4
yysS3m9NN68UNfGIh1px6ZOu8zXCSELDNsc3XrByxTh95nHshX/6SZbRegnTDlOS
y/Q5Um3q9ocjSawz1C1sMl3U2W4GfL+56JXmQAZur1fhS3jX959a5GmKgfjKSvuI
8Dxl9F58GEJx+Jvm9gnvCaiyogZmQzIgIGwepOTUBWcshRmEwUpdt7HhWWfSH2nz
NHmmbL4dxThH9HG3gsuYR3BsJdVR15OFxkyUIhL4646qCvRSVaocpFaD7OJDgdm8
MrGbNdySz7ETsuB54Y8cgKnDMlWKwwM+29kEe3RUBjBkY0hTSIIy6nsfldyKYec+
qqXMSlOsG986NP82fTp4N12ND+8RzQOHpAVdAcp81lvoiF6d2+EJt6UfQMUNf2rB
xbNmVSW74payCtvzx5EyL08sMpOLKInbmBFRtz9TyUj3/Y5IpKbZ8Yb3ckhxigfp
d/jzD5C03NqeDW7MJEahhZbeWpyI711t+Qqf0pAtDcl2P1zivoVD2Fqyh7fTcQwl
MwpdmqTpWNe2GirGZfw/zejQgvhi3mjm1Wi5D/ZmmTv+tMX0ocDMpkeIraEW3Oj5
GU2q/8zVBqI6yxHtQ/sMe373b0/+APymwPdOnS97R59QbUcHWdaRG1HKtz8L3A/U
rAprlGUOhO2BZV1Racvk3oyCrN0FLB4+R/frFE9E19e2XRFbF8NweQmOmTU4s1Pj
J9nSnuD6nguuajd7+BJP6vGLjQjVNZZON0L43tbTRutJfQ/MMxE6XKnYoKprJ6Mo
K9ArTyAl9tK3wkGQ/lmf5IoYx9wa9TUED3UaT20x5p56iityUiOspM1ylweqd9tp
jaUrW6yjnU4ZZoC972uftUt3kMKvBaQfce6/mBL4VpWVdj5UGLIqUzk4YckOCuYI
DoxbN3KWMhdhgndYhsH0QXPZU6HjkAZJS1bYwlArlFqvlTdMQvNIEjdlrVGGIISu
tfs9eHCoQD/PsstPcNcnx/kwFYZiCzuU4gXAKBZ67VbW5WnlGYQVmzYtHbiv+r/x
hNK6l5b6XIpkjsBHjyfdieEjdsrSKjb98vhVJ556H90KMlB3pPPK6P8KVHdXhNp7
6qMfVNfZ0WxoHN4d18ozS0+zuGxTsAIgCOtmCkHS4tYTwOvk3vEY7C9uZ99va32+
0UTFd4UHoq3Z5jLO0aUEZlI1wFThEVTikR++w4qlfTw1kd6PLuEKZRGW3a42by9A
6wsgvBOWM7x53ywDF+Xeok20vYfYaeej9MbDcszTl8unYeFknOb0cGFIBZgbTwdS
TVSeY93Uv7c+4ZHxa9DdSwWC+23o/I240Lh2kp70BgHo8k0EZa6Yhiv9u3u8cDno
C6D5OYjQt2AfiynQiGBDx14Z/LLhEidf9DK+lCtYYyU7WYKGl1VUs9CBlQHuHxff
k4Ist3ngXNMGZIIQSVhD6sqTV8tTj6sAHWEuhFIDiUNyuxbMgQV8EzagOevSZ1zi
QiwHCq9r/t2d8G82gcWH0vv132PFtqIc9/c8wbKENUR1GL4ktMHM9pM7yq1KLRKn
vJHfuMfqZjezU+5L5asFujLFpA0KM7Iv/0V4DYO4bzE47VEoy/IhY582xh68urjN
2D98TElez/KltmyQbrWIy/gY4JWdoUgFTJDQJz7yhe7snrNcEAlXIpjxScLVMLE8
H692sWXxUwU1zieXvwPBwQtoUUsW7v1mlql+ZrWtIHyaeqsudibt8w0PuMnsTypG
s7FJwP2KncvPP5w++7VIDPZx8Cgxpbtt+tme49CRk/TpxiK3g7+BNPRZpEgTGBTF
5PZB8IbOqRK9gvi+vo6yyIcVihI9e2ZZVWhE/gBDr2+dMp32tOT5quO7yW2ez0jc
K50SmrOvNooIeCPseKarKLZpUnmR4fxXz8Of1o3qch+x3TNd9Te3ubQRPLh+fwa4
BlemN5jRakYP+W/Z5cJ5wCTs+6dpPVzTRrQox7Bw5hqr+V1wvsOY9pUXjNbneT/w
cMBdpqfCe5gLuxBYTA6XFJmo1jz6TUdOVKtjf6StjUt+Hzx/QU6AeptCREkaQKCv
GPb/A7qZUtw7Yds2CZB6YRMvs1l46mydyua0rNZbkp1GFYN0U9chWrhqctOfLDC7
FxOseOsrkoWmFXuRxBV6nYVhR10MY3sELcRMRCuQ9HjTvZkA5RIHavUTgFUQSeQ5
NeTB7dMxO+uVWPjCfzuoP/fXfYrNzg3ecpouB1+Mg9gWUsl8cJY4+bD9si6ZSO6w
nLjUi8tLUhQP/YXEilboFB++1Vqo6iwsrGpSe8vFuuz0PgLyeJhiFGWXkZqa1m3u
rYLiJZGAJBWPZG73He9ku629bnrmE+QLLNXK/991dOX639nSWuq8tJ4PqXP1JET8
+D0ndB5DKHtp+A+QWSV76ROqfgtSO96AAwYCA1yiothr73f4s6H4Os87YXMbjXOX
fhplDOeysWrpbi1Y60wCBfXA4mJOnqD62MKWsBgqL/kKy5F9PPAf8pyi+RWXlObR
OTjUW9hhS/dEZncgM//hp9+Twe+KnKqDDxKfGNGqy/DJK4Ip7t7IygXJDyLtKdm4
DomOdGzOtUy9CkZK2fz+XUtn2woIBAukQboHeQoG+NlDvz+99j9Xga0hVh8gdJn0
X8WeoqwFy7zBrOwe1EX1ubdzmB5bc/fDTDgQWXW8Nt5jNYZQq7cGxzo76oAORh4R
eTb+uUPmgeO2ZRSUXRD9OFnCNAck1dy7dDvQ6fgqwEk9rB10cedHzOHp0kLMO/Y+
l2OT9hkgPMqmtP4YYQTcaD4P8UNuqkoDFLIT9KXDj5xxB7fkKjp8B0aEYzBfIXhv
s5RjhWYjRb1WLV5LLCZ702yQOguu5HOHgNQy/ekmdZ+f5Rjs9eB2MyXeaoZQ7V7R
TcpFPsFwkauF73+lQer6iyP+zDomVT0uwD7a7sc96ML3qnCxaJZZ7ewbEpipGNN+
JIJ63XMCe/Cf659JkPCCOZkO44O+YOgGQ2IFH6JKvIK8CNHDaE5Cx20hamkqNJl6
JGvRAb7h8IjvJEPlVP4G4kZg9/Pf4ihpyX7O5nqxAz4/osuTIJ9zeZEfiqHLmE3N
CSHRt/c12QL9paparLqPS4vPE1jLKOSq23XucP3Nkl9eEeSjkNH5xS6rXNxQIZtC
TA63sM9HB/b5kFEcwW/qS3MZ3vwcAk4GEg+6w9zdeQMYRirhOX9UruXjT0/wmLQx
rUA4puzBfjxMvsu0hd4sv4Vc9PTC+UclDtETKD46/v8nAW02OeanY25yjM+iyROW
ohqWBbOcpRhyUuhO7UMxQaWXa7wQHuUzFXJtO8i33NLRfDluoK3bMGTmOJ9cJYz4
gg+cWN/h5b4P5YMvv7FUtlOo2c+NCXomCE9VV+KblcTAmChECEMaODMvVZ1qRPr7
vcLLeQbxMR2zRSUcptP1y3/y38DJtVxVcjgaXCaUPVBKuwbUYvdeTkBWLG37cde3
7yHRO6SKA6ZZ4bN8rRZ1AaR28UPEdN8ZQyAER9tcSeLsGyn9lkiubNRtP3FVLAKz
Bx9yJhxdxey6yp8dko0ZKC5HDYeEn5p+v9KB0JcD+0lIju+WmFKST7DoZ7SUfppm
finiC76A3uDHtbXkPnkkf6/eMsB3Xwg950NE16jglnaTBS8eRfUZa4R9XiN06p87
6fn7+aIj4KyBuE9DJmmaSj0u48GNEXoa9HJa3MKIlQuEK3sXXEJtr9L6eqOgNA2P
8L9OgR4lHVmrORKxBM/huz9k10ZaqOPahYvwKYW3VJcV55WECQZPyyV0JR6M0Xm4
sz+z28xm4+TTp0kHJO7w0NZKsSfAa2x0K+mWkRTteDz3fLs5xGakFw8hWzikkfqR
9RuGKBNJe31QzBx3B172E5DrcL/vboHrLzztPPeNqOz2kZgjI6Bm/rIyTGViOcGc
3IT5W0GcPFXo4z5CeGlXcQxBdLCydeOb9Z8mFX4RVge9KbQZB9t+owjxZTUeUPsZ
dywkx6Vc7gqAAhXqaUuPeInzV2LvpfbyAhk2DvqruENMTq4NJLbO6oZ0FY3Ijq2z
+6ywVA2Uni2QRorFau9OtNOv28qKoNEPpNIsiMifeh5FX9kXvBts21DyFR4Q99ZN
gGUSeeDb4TQu56YoMfauajC/Vx2vfWIhH8wjd4WpWFfBnm6vY3zFUcFQAjYcMgBf
yExPerAEk5PkEIpkaKISHp5zK8EC4wfekHKhcSY3nZXw1VSWRaXFEviAhFeua/z5
cI9FONywRvHLhU/CMImMWUKPbg0GqvVtQgDXqDGY1D4pT8u7ug0SsshzQKYLXGgf
EIx7dMoQnDWEw5tkxz9elaXonXXPImybdhxdBOwxA2Zlb4JjVuIyOwHqC+hoUlXN
ssyYMe3a+r/wUfkJ6Cp/iS+wrCK739FvGVDcI+73wHIWZWt7zbqFdqNVSjJCU4cf
CbWpktB4rjDPVTc7WE60BpSePqiIpKgwb/8rEncE0BttxgrD0inA9/Hkhr97YSfr
X8/RhDDfaGMm0VE+QtbeokGi6WaP3G5dXRhPifuIJPdd6D8h1GJh3g1tH6j+y2Dk
OMGiW6JYqdg3k1asG3Q33/7WVCZUrHx4KCueaEIU4Y73hKPEWHRXWC/s3SP0Q9Qb
dXSASWqO+4RMAUqyF07h/7JyCOjnOXyy/9NxfN+esiSdvSefkLeXq9Ob8n5+9zHy
myeFs5t+nlP1GThnHRWS8CJ3zzeYPpUF5Km5TJDlcShb713RtCWMXVABS1qNSFgr
33sUt3LdMlgpze9zntxE0B6cNpwEO3u01C9CcLus+VdziWiVs+JMftAVi26ujIpU
XOaNIWaWUNVYAE5CT7BD4k+TZgP/yZImCOHsF954ImjEYFYNu4sFa+5DEBWOwjxi
Zetslb+CeYbTR3Ou+5YC5bBhHYBh3haPKD/+fxHn/xfCDpWhVEMBk2KhdaCtaAuq
VvUnzHlJ6Ufscov3j8RSMhycLsKL1zaBJ/yfkBVNATaBhNAfr+vB3HAb6OG2E1br
GIdmh3hXwGs2YT/pPWYwCV7WjCPLB/azFkh0C91nBAnjp27AvG/fg4YqcAz5ghrZ
WEoEqy61Ca3usSENX0VSJ6B/APQj+oe9k0BTFczdwKChn82SIidz0aT2dqauK/DY
4JbrcamqXJVwbPRZbKFeP2jwzKSA0fTWQJtbV0JNmZHNgWRPjTSE0Zs8VWcb2Nw6
/o4Cqy7ptxMSxvlzrFxQmAYA/MmdMxdStjJXxMgpCiKRITsggMiVQ8OaGoJWHp9/
wEYaQ/alo2+xMslS+YDkQFN1HFvggvLAIPsSkonfr5dZMmBrOARkrhhZs0onqfJQ
sUi9DLEEsjEKaBXvt2UXFURW8mMt5uEfn3PuDy9xmegsPLqJ/1vB6/GqunzW7Xvo
tRvx/h2N84tydEMaHRTE+5RbDKHe3OhoDMolfPBpzoBAXjDiBMGseaP2x/7eqKBo
30+nD+8UrpmFu5x7ZSr8sETXVuAdcFax6Vd6NJzHmkDi4WwOujXd8AI0BQ7a+peG
fmfmNRcTaJmb48kVMeVEzoKlCY17dDj+PB7iyJNrkvtWuKS6UG5r/qY9xKZHdRL8
XBe8+AGLTD14mxicckbR3XDPJ80b5BBG+3GW4sEZv1o/1YJu4aJ/EziJUsSmG7pi
3W/iSj4vpdx1Opt9hNph7KjXTB7/iZ5SwoQBFMDAqm98ASMeZBan2VHg6KhCjuSQ
O6A0XDtpb6zwFSM0+2m8FvdpVaI6pVC6XFEDoVYeR12/44V+wZ0bHDe9A6aDnf2J
DVvzaqFXVMBx0Y1dbUfLmSCxe7tZZKneVme2SZT5MJUPiJs3RJDccd1p+IGlzHz0
xqqocE9SwygrqeB7rGR0epLUpKQp39fehm+AbuaGILv2eK7ifDaQ0iKLpijJYCh2
8K4n6j0Xlc6L41W/wuMAOM7su80asyFP0i4hAAcYZbWZ7t7HdteibGY8Kk0Ne2jy
32zxBh7jMe1QPqUjuEh0p09DJeuT0G2lWlsj2yDUWZ/W1/PkcCpeXcLRKK9I163r
iIvQKdINDwgQG5ehWnR0202oPDkOO4IHeYBE8tbJoQuH73lXesjx+crF+6GdU2qS
Lpy07deZLQRvs9MwOr4qmgffvpR4kpl3RtwJ9j/jOKutsaDAo7UIAWLrrG4eeHu5
Nuru48Z8SC7LGBTFvqXNHXdyEfNHCh5mVben8J/oYeW3MpR0LHYDwMoGI8b9WDbR
RKO7FYLOJpyZmpcpuPTKpVqtbXASJ5zcNegbuU14D3iv1k3NF//3pa51ZEk3zsBQ
SX6kQfvXXomxTAkJwzyPg4+6Dy3LpzeiBrTab+MSeA/guJeFn/W1bkoN37WLAOxU
B9kjjyJVDnfByQ4zVHvTCCRgVJeV4rpOAvN/Z33jF3D7dotmZeLuysqkuc4CJMKV
ELV065RQd0hasCW61OEmG5BGIeK6BfGjGfa5SQJyY2r8tbYWK+mCj48oG4MS/0gI
mX6lqV4S0GA/8ZXbTmsKoMAPziwS2MNeN3FCOb5U7J1WHL7BfV0lv9fWXOVJHVuq
15i+3vuXGlfQDaS/dp2uXKAoMxxEUDB75R/UsRzFs1gEsvvcQ768F2YRv3wsVw+L
ULlDCopMbTuf7m7UbnoQJhqW0oYqmiqKmK/C4CmhPITMh9cot64UKZ9EmtJ0hBuX
bg1Lg2lNBsWySKWahuTgzuKZY9Ux13Nq0rUBb4raQDXyojBFYmpIFuVjr9eULdiE
Qnf4KVZGlE23KFiiWXEuV4967T3F20TkWkXi/dhzwaXDHjl4e5TVgwGeOeWjTf1X
NgCGgV+18xX8eit6LBryOBx6bnK9HT1jrJpzzGkw984HW9/8BKPaeDaCAdaS1DOO
K1l2NzWK/STc/oTCidZxZxshcjDBFTY65mlBGgU0iLPXPguQXqYm0OyvSClWBeXp
6StdbGvohtiZt3KyISXciodm/aybtwFcMiQQLv/vw7el84KdqH6HkP6SHdvoiuWF
izhkRE2S6UVKff9Zc2KV1T8grYuT1+dNUa6wu/ZaW+AlGfWeVuaL7jKsh3B6fODD
+OVUVQo4KBdL3DYtdTbnOtnxQyCfABENt3rKPvgDOorRrsdi7JzvbI0vetn8AeCD
KMPw5owpk5X/LmROQfHAuBLhLfmQrErvU9/LCNp0GOSFqh0W/5VQcRrEh/0FuH8S
ADVPM2b4Oq1Rn76JyUXwmo5fm48M6D/qPZgaiiLj5UQFTIgCOwS1zxYvwqa6Vd1l
9eKEaIAo26rMyOAxjChhZ1UfnhzUAgsazuPfiyU7/Zo0II+yGMVqqz8rzSUTEZuw
SRlqhHtSW2qlLtiXE2XOR7QOyig2OPx+nIJUEQXkBG8MyGjXFJUIOLZmikK3Y+db
XF7b6ysN8O3AeaNRtSk05IQRajtdJPhG0mW1Z+QEfas0Ve0T81kkh/USNucFO2Dc
TP4bAUfM6P3gTjBR6pTHIamt0xGPBZjExdPFtJ3fX5pWxH7es/JcIRNZYIs6zoMm
MEvMWCm/AMhYVKchIn1b+CE5MtqQtbAxrUmg5N86kqrioBgb4+6WAzOf3FYafJwg
vc67dUxA6rjAGXcaBQKuyP6rntbfFW/cng975nFU3xocEeeanKxUruwypx0hSFmr
RtRKPenKKPNxBpRLUbhoG4pH3Epdy7cKoOP0vM5YvP0gkAQzKn10Z6lNIgtDiE51
lt9qcEYjfKlYX8OtEcmUOHapCYU6/QT5VLube8SwWnxL5MuMjavo7wVrIQ6s6tO/
oXTM/l9VlFH4Pg4IjdX31DSXErlkCwEBU0kiPzPg0cxgWeWBXbWTHumBWJj82LeZ
ADJ1r5kvntRT3EwIXEiUd79fSUm/oyw7/KSTC81c/vLbcWo8ZEGMP1uD3AAfwuxi
NZ/EM1s2Bp4hmXkis8aywU4p3aZI7lbx5BPstPq4+vAtlm3LpqOuFINedAu40lRR
CVnDoFFfov5fHH2MmcK+Hiloz3Dv+ywGGBl0NZxHWEKCl8vVY3DzOAN4MBlPEpUz
gUEBjugzpf+P383DpvoxMfAdpkz+dEar3T1v0S+p/kMqZXyJ7zU+PyfJ4DSvOPlA
lkY4iJbKtPHb9LkQvk6j0Nzaa/tbHqrQ9nRSImOseZx9kv0GXGRJlQSQCoSKAY+B
5rJaek93K6gmEg1h0pEsk8CRAtvV7MkWrB9jPyNtTk1iicRPuV9Hieq0ClWdc3hB
ZRC0vs3BHIZTgMWQuajRdFgrXVAKXhbQ55hdPo1Sbohmq6fZW2B85TfAAMDYcXdt
O6my3SfqB3xT4lIU/n5O2tm5X5UMIbdBd3Qy1cuiecK2d5R55CcJf0O2IVHhJhxg
+bAs8V2xq7pdAH9V8S6p5zpbnhJg3oRC09Bq/4sLX4gejAjesmGhSPoqrAUpCh29
HkKIZlY1mE0lCI8Lz1gElssghlA6T3pvkVGiUfwnBBPv//KBasYr10pmjqw1Y6F+
nxjyYwJdwZNnZ5FyaG6JOv9vVEJLmklQ9o37+frMKll58SLWyLxQSeTESDyoFIvv
rm6scVJBopXEAop7q+PQXVNbV6PzPWzJBpdWq+EqGA7FmtTp4dcqMXNdzuGZuVWM
HslCeMjHP8yLR/jfqZ4ySro+EfWqqw9JRFP781SZZJQnQdoQhO7SWwbloPMm6RWG
/cKK2H+W1WUV3lfBUQONn1EzWqCqh0hTwl9BznsdOwPmorZiqNlmFSWXgs/Tsdxb
//LcGh1Qkfx8iDbWTvannFNh67cUVM9BA7AZ7GcW5APS8L2KIdI3RIf/NXT/tHVO
odBshn8n+WXCHbHGSgBoKMk+AXxPnb6jlnmRVU8pyxjVz4JpUmN+GvYYy9r/LktP
hV9toBlk+yYSvxPpXG46oVkyGdumyh7JVvmoCnfcBzzHL9rW77Auzhcrd/9wlvhU
Ie5UqZOmD46GLRdkpFdakIDvNIsqSF1/jcjzRv7wpVFNHU49XKmhZsDcvKBPQ2v8
x0JgFuI07ad1mkNAnIoTAdAQPZuqp/ERc4FTdTz7LgI2+qTsV4aKKEU5grufDB5Q
zcT/LOsgLNbsjBFYyAvBV0rbOnYxglfDsV5LoCIK66iufWvI4TtOrpPKsn2BCoWf
/MVza3mu6DmiHDfX9Ttj6NARXCxnAIXY7ZtqrIvlYhy9BPiva7JgiBq07oL4oYTV
MU/duLCDypEO+Zu8C3hanbDhPmb0gFlVfid/c0auk5V+A42XuuMccxHRVZnTaPPw
HFf+WLySaeVuomp9+UjRze+0QKY3gJ4st6ewvn30jw8Yqbz7WqcU5WJBw+umUiW2
BVWkH2jsX24MkYN1gBGo9WY+LPXuYvuWCffgtXXfcSsulnWLezvNiLQiDGpG0N9E
+UjUWnZirIuu9wEVcmexXmXexgvEiwfXX3gzdSAQjNUpQk5TMSlh/I31jEYsQ/A+
tn19G5B4qsuwAR9NrjSRwed4m0gb4msLQ1thRMfIBaEzgkCC3Z0FWqYrhKMObjaw
LPwt3Iq9j6VGvyzNLPSsF33ntn7uc11gTuudEN79HHxQQ/Xg/suMH2lr7a6qq9ak
ffGaibSuAeynq+5hjUn21pSPasZ/zYr6UYLRtbjnIOjHspZoDBjtUdHFUTxphi3o
fdGSTQ2baZ8F8MrLB0V5+jvOXA0eT8Ew/korQT17BhCw9OMTyW+CAxqmTcA91moS
ySXwKf5ZDbp7XAk+0jAeqJCfuWz49p+wpA6KjopJurH/ZpX7xngK2yTQSBxwLvhk
yv+mBxkK3g0Zby6zKMruDY/6FzdNArYMhlJ1aMfHj8Y40VGMWBIq+iKW/TuGAqkn
rqw5HT47sIGmzNaWD3T/9UNtZTrBpsbFZ5hAHT8UTmANYcEK8T+q6Tz1eVfH+Nhy
HHKPc/WauBlpPe9aqf75Vgmd6BLnMtwXcaGfTCHWhFy/JajHCP6wgVmpkYLa6Y39
zaP2EfA7tMVsMJ0T5gwxtO6jCW7BIw9SaXB9R8S2qIKO39GIxzR0xooiCX+k9Oas
JxGCPQphqEEn4dIlPyv+KrP8lm69LKBUEZCaNQxQkQL+PEJhkm5ExvIi22H6FOoK
gngRO63tf4QREvzBsioWyonEnfeQFOAXX6e5eIpFdswT/rzyO4y2iR/ixwxlrBFa
KMJmdjkdL1KHSsmfpSmVggVL3o5AS77pqQHGSGGWarbAGg3VT7Ubr0iGma4u7QUy
AIsi7XLQlI5OMRvnB4yGwYwWY2P8icNmDhGJ3L/zWsFYkjUm3Lvh7Ru7sfctaULi
aN4y5cFnKOwzUcr07IDUteKYkfTMfVFwnMhJaGKEbSMMVG8KLR5EplAVkve9ANoR
w0Tda54o/jPQhfIoDew00w8cHaO56XWROBMpQmq00/WgIdbpZDvQB4aH9BH7vtSs
oeEnWySx1B2+qokB9a47o9H7Xegt8z8Q1nFyO6MUFFrivlIdb6ff33xMnhdMEeCg
w6fJXk4uGttp0neUhwDQrNgRmXYExSByRtybiA+6sevC0iyXymSI+BEwrNr1AMXV
+3TeRSiKwmJC+ezOGu7fGNn3drQVNQJlgT/0VYjgIG990Gsf8kUvsgUjDcvOXeLQ
rYLFBF9Pv53mHjyjwrzPOEuJAihqciHAkT+XR09C0ZzHhojk3ehQ8VMYEK4zuKOP
Uie25GHTJQebK+5kiz899irbkzFmMIkYISXrwasZ+pc3Tdhf8Gv0ui39QrcTlu7R
fxuQ00svHZFOC/P1voPcK3kTmUQxj8gGsNCUQH/wvV9Tzt0knQXE8GOdusOgCAVK
O+ZDQQVySEIddSbOgGhu7z47OqFHC0fuzRbi9a0OXb/HGxGeuc+nvoXTSSTcQ9+e
+Xhk+ZKOupcUBlDJ0hNpLdSi+sF0xG13VD4e8VDoZzIEivNrNXC7fgFYu4AjmTSR
5cMt3B6HaAPg6JlnyN1ARUd1eGKiuDFf3So25kMv91e44msdgnHreF3sLKK13m53
lrQAMNlaAu5rxPGtZR7Pig/akJ2uDkraEc1cSFA+f9onKuAPI3D1j1gSr8cxPUhq
Uue+4zYbzomEzgXFcjoyKbWj0x6jRI9CjGlanA9GJZ5lwz00z52hUccUTkI3SpAR
p1qEGfvZdAPJONHEAea9GG2vPcj6XXR0ZZpibx+fi+seBt+p9eYqYPombROZjWB0
PfwDcYxDvxVhgiqpaUjjFfq6HjHxOYDhXL7GKeZ/awB/WYeIKHpPfkGM9Gmre57Q
VxL0kY/GlEQtRMHu6oh5i0ycbYUplfZNozFvdqzYdrC8Yts16k6ozXDFEt+AFf5a
slbYHcLNzp0WpwrfDSMskT4Y86dy2wMvXnON/O/OGCaZKmZNevppR/hcGsrZ+f7H
/HPzW/veUzgGNEEtYpW93MN2qIwXZtE0dbfE6uFLZngHI+ZYfYpd4MJGev62uWJj
aDro4Wca8IozWKrpdeZrN308nP12eIuIN0WJuYTbvSRRa67uUnw2CLjalrYLgBOz
0G0pKwXp6prglRC6np0RgpBmbNSQW6H/4Biyd9UPIBOP+e1T8263QOqd5ffmGEs1
SMCkTj3cbCHtfQ7KDHKpc1hyR/W12VNkttalo66hyWvIbTzERvRkCKZ0zNRGn4gx
MA4Ay+Yaev7XtaQAEV2iQzGQJmco3qvmnsrNipwTBF7Lk9DmzITlj7BFlJRCEnwr
MiDF26ZdTD5A+hYnLMt5BsGL6qKOjE8ga3cMnw7DYRDdMta2cg8Hu/L2xt89rWaD
tmxZh6KTdli1cpcOlLMbJVsiRF3e0dFuvyCGRYWcOPula0GZYwsbNX975Po4kWp6
pDNXqpcApa39F29ouFg8tKm6xYoF9234+D4pU+0qSranAr/3gREojXUcBIJpORLl
o3gh0he9vc/z3//4eF7AjzNoXYQB7GhNK/WYe3GvFcuQDzjuv7Kkdgy4o39S2EYV
ic6IJbWgX14AKlRjGFspidQVBZEP2w/NIvVVAWPW2O5v4mN65J4ePv5T4KRVdJ85
j0JcInNw+BifFwhhcCJN8GyAM4LiBdPYGmMz4QNnExitPVMxX3hVkmB0rWE3ramD
cIRhsuqyK7jRO+lnNOBtPG3EkoZlBEmhNWA1+Tg+dNjQDhztURzL1AoDJbTqgkGB
8WrSC7sE+JveDIFizO8BluL2D0G7BYzRWxwZ5jsvWTyu6UoLXFUTT73U0RJ45Qm3
JDYbHTFGrd6HCyD1kHdyvBXpY+mtVI2Na4Ysm3z9GYBCxO4S0f9j2snQA4MCeMrF
CE6GsptdXvtygJv5NrbDLKIrsKcR0lStzmRkZ76hcTcDZ+3fOQcEweRPiBrny63L
b7jOeeZLiQ2n9S51xAa+McTUiOKR1+3IAK400lkOAQcjx04I6CDa2UKbD2CWjlHt
WRyKwZ1F2iuiTdc2yYh858j93gxiMR0p/3Oms3l3PcJM6zC5D86d0e6ePkids8oZ
CDsavhZeedP4SblQDfwYcZMaftVh/5R8kpkXrXr7116xm4O15W0di1bj4MUWgk/9
8dIXDAA8KVqcW9+5xz7B6YE4VWnszCBILniSgP9jFSOdaJKaf2Tbsh3CurJPBmBd
eN6zeR+6ZvAs8AeXm5uLd19R7y6kCISN9wZ6lPOxLA1JDO9b4es7Orn3aohxQoWt
/19s6ysOBspqil/8jZF8A43axQqdrnU4gQnAUf5e797LV99RuQNWDi5IKvsMmW3I
ycXmi/ve0MUyEOnE26pVVNCXh49Nw/C8DlbvqbYYy05hJZrAr178uKKOZFPwbpwO
cbmRHMedhOoPlInFSr7IobRLM61WMiNW8Lit199kO8MF9+sEwX/mxi7BMJgRtbQC
i6YfnnRMthORD1yhizZ/DQ6wUEsd2XJ0TBgWmkpLHZsAI5dSmkG4nQjk7giN/49s
lZe2wniw6QSyJ0BEXGR3zZWtmTSS8k126O5Uk8YAF8YBZo+nce9ucyefvhihx3se
Mk9/FPcdhHvBocvJcXglxVTL7cpPcpO2X/OqfNi6pXp9LE82FV4C0S3plWQtSPfF
+/Y9TNWMn6A1glxXKPBFCa7gfcfSsHNhd4ixf4m9QUMJh0nO/O4f6OHuK3j8RAKA
/Fp7V2JDtU9fVgSSNzvUV1dhXXMgK2VtErLV6tRrrqYSRSJeICyqQxUhms2Qcze5
9fh7HzjzMVu6lxXHbdI7XvYAzMlqYDPbHwqkObk+YGMvZE/zd/fF/AWpiJNVhriz
zDmznRdkvCDWuyz/LQxL92qI7zP7PSUGBO0eT8RVhZLsUGEhREnPTgJkyRIAMd8h
iijogjvl3Kc8IxDi0Y+AX1FyufYszX1gRyHrqpBBKYzcyM+ySl2QsvqUSTK5yE9L
ciT0io7lRmnp2JWVemVT8xW5Wp5Io0m7/Ewvd2PW4k1KBjnZgBqeLbY4JlkRRtQI
pOz9tK2l86Px+mrq7pfFZZxIkhlQg5KFbBPF08m+OVcWnScCfUemgdKp+ZoPKgXC
4NOzlgE3BDT0ybAKfecfQ571BcofgFTkU8jOUYbJ4gnNBiOdyoxMNPoMlz6RpBiA
JALuU9X1XhcM7Ypraiv2Mo9qD/+JuJbUrbO3QStSU2uFV9iQelDLGGF5/0HPxpeQ
Flq0eEX1D+ocSYQyw9yBx61UanHJoUF/d5qGtx9SP98X/h0Kk/nn2o+qcIY2RWsV
57j1Dx9Q5wWqdNi4vUdZjCwMxGu5U/EOe2NLqbYAg3g7Iv+343xkMejTM5KRnpBd
c3UFvy8Lpw8KNxSG1rkThVWRQgU3+AivZC7jzYp+vkM7mdNkOc7BIAt6l4C4xAbz
XZ9VRdJUN0hyEdDMJS155E5OyUj+fVl2P24hEYXJXKdUYufmtsmIpD9+ydFqKWZ4
aD7zeJ7Wgcu2wuw5xzfuuflXJk3Dn+eHTYu/S45Wby+3ENFPlGMU5lCGqqNeXtWP
+cXpnEgYvfR2yVT0KgXRNTQsEH+YF9ASO1YzHxdUniwQihvfpzAleqn4Xf8WKGOM
7hUSZaU/uui4LfrYLn8dFSSt3Q8ho33PGTkKZw4oJJTg4VbRWrkZlAbHTIVEaREn
iXDPoMRvTbMO6i4GxvZ4D1pZcN9VQWDWypj7wtY/75xaY/QFhA0zFOu6mZz+ycgJ
WOfzftAMfa4kcEMraPW7a7iccn60BCUfAK0T7Da3KosCJnMJdNQzWKqWTyex+KRW
j4KJhvH8vkx8cqzgTbwPQXw+jDkkOBARdHn27vAad3+SwAimfLdR2fs1yGotuu4g
CBxq7Ecc/uVrjGlFzs5062ZTpOdlxc9STyZR3zNW9hJeEwvHg1tLIAVh96bq/8M2
4rZ1V4oNV7w+Yzra0/5ycb0CYrkyP3sYNLCoPssLJVmzUeB+dect+p2o4YNn8j3J
pxu+1vj++sujGavUQbExvWfbUxkY4Qhbu2YlF1LxGsdR/CV6oLBUZ7zSgevHMaj1
bQQh5AKZCHVwIh4v1iDIudz79wY/4RxfUhSCwB+yty4YwXKHogXnnIU7DtZCrQYR
P/wWu26kTBR08hR13tzmQmwHUrDkT4CFz4J350dyQAbVkpcdc9dBL1jyxCVZrghw
wSXM+JB74zQHvGU/FaB18WBKzU2d6fRy8zj+JsvJXIYnd0+bPOGZ9MCieXBQHu8j
x0BjD6Or66O8LvCkVrc4anFJUTMc++eZCOd9GkuyjFjrSghRyhO7jvE6Eo7vJ2gk
SfWN7sfPvAP8hGo7//kr8Ggrj5lkTcPhMfS7YRgGtxtII2loxOb7oqQXxDIR+RGa
qprF7Rdp7Okj5SlMH/+sgsrCAPi6mH/5KMxHlOD9UoiXrBZXVrg2JOXGfKL2CUpq
Rb6ne6hhvcQs2EbYupH5s4oyc4B+8dv9AlMECmeQiTKsHUJfh2ND3r7IuGsx1nrW
EgEh/tHgpqhp5tDLgSNh38pPLDXR01zfuHnO/MID9oU7jyVTZ/atIO53oBR2nWDh
IzYNvgeRBRPybvxmPLcx9eUafK/iVMofhuOo0fKW/p13MkVYQYV/ktxJY9Sz+iw8
kxKlIU6mtN5CiFCcTas7NvBLo/4COnByMCBQaFs/NiFy0ukZrCft3RpUsvwE2xKa
4G7GnQiKRiwR2XvvHlRA0hcEHNtTXlWiD4Opmyu27+HNM363uwkAIKmM7px8jknO
iYd3LuXniJJPlTWDqumIM3ppugegSkA36R0I5iGKTgLK8FGTZBM20cHd+yUrzzV8
P9hwtyhsPfyF+wzphkMwasTj8GUXqUfxYF2NBrTZXom87223BvQv57gO7uw1SOyZ
ECkrzxKaHn5oZoanhy29Rr5ESPS38b/0Vosi/7nd4MJEaS32C0YkzINtWF2y9PO9
9/wUmbmYcFJteKW76wO4JrsKOMMEIUu/T26KqaNcfZwS7bprhTT9Gncs0qUw6Hwa
WjtoAQFiXECr7BcZIX+mg8aaVerS+iMLHvkIJ9Z+ivaKbipqqe9nj9iBD6yuTB1B
NRx8lMMQzg7u+uPOFz3/lYlslwvaXNk3yUvfL8ILmkfdiP452oqOSUDAQKKvgYyZ
QgDrYfd86f5RmYeXC7PIBjhuZhlS7BFZLhS4BWsZDsb9rjozn06aBu5bwxU18BBP
wd+z0bH+MALHbnyEX91jAg2JyzoUncAsC7AhJtS/6mJDlS2Xrlp8AtHTX6sbOFJm
M8Gsue9eSLoR63MhUMsQnBm9lpSSp5ev7UsrEChfc00rA0TWpPhiXR7sTZfDUPve
YwHrC3vlYD/P9CW/8C3ipFLvTs8o4I5s08Sdx5AIM4BN/xgvBgWNV1Z/h4KjPruM
GC3ZobzD86B3Lx76eTdVZ1bs1bZbQtJvD4jSKE94iD1d3SUdqjPIGzuQVITXW54K
MJd82I1dL5hJgXuAyLoe4dwAx6lLs+Wcr/RHpDGQ3l6oMgKViVka0IveE9ahukrO
puxWbjEfqicx4OLdv/BDzUIXuuZ0pRfffYJaggjA9/u+iKiiOTq+EnZvPnacl6ID
sqH7h2jTAngA5aWV0L2ZYgvfGrsDjiknwy+6GK7H1D9hAI4uOWAvKqg/d6V3hEYe
Kr87bezcDrXdiPhesKXYmbYHmFkspMaxmT92D5GWqi5whb6lCzVuRDS3ypO7VC9I
S9EoNEIf9F8Lqg9kyXV9Ia9W8YOnJtrkdSDRM6Dy2Ao+O9shdMNBTtR97ZZ3blo+
d4fWVelwOoFIBOwZovl/Ph0tWoEh5UwhJyESd3aG2hjwVAaQhzTnQuFTuO1mL4/Z
HH5JmpeHhFOtf9RtLWf/MD8M9mV67MNsslD5T4QM+rzA10d3aMsK5Wt/3m6OoXzl
C9/r5Cq+FwwE/yT4UFPVlF42A1d6toUJjoXBQJnjWdXy9/U+LIeXqDSc2FefA7Gw
DJhxZ+Qp5s/tOUs5sZLLvgrBFFFNb90qSEp4DOTZ+bU/POnZQNEAR+qn/vwHteKE
bPk4yc6Mml5aHSW/YF2LOAWjRYx8SUlUZ3w6DCVEvyLB7kXwNjls00rynDIujk/1
lvkVeosTViqNSqWtPNWSqPDb5DZNEeYhD7WnPG2GKOprNEQmi31JLKAckMMHIRlG
Rd37ulpTBSr6E/1+uExuj03mh5TI4JjodcPQjsSvKYxPZhEcVlu/ZTKLfi4Ujz8p
nqjgb/+IJ2Zs3CgI74fv4HNHq+FSkX9hpZQMaCjSz2NdiQ9QfgFNJcrqv0uowGn5
gHQybe/NWBJliEDeUHoGKXt7Vy7d7a7hcSNrHlN12IO4XEl+PKrzwbbqQBM20uUx
iVOQ45qcEUZVdqkuIpkM0mAl7Bd8V4AQdsLmw7/vkRa2XUU2zc7BEKJ4e0PC5E4L
xiG0TqlF39dUbIZLtCkdBGyUjsiOuMMKTEC4O1GCttacA5N//1DtrxqczqKhmEOd
+R3eMAkOwapWpRuqeK8Bzsxc3rWMta2hJpIkMlXQ4StXce6ZB1K1avHieZ4oPvVr
xQLZ7vJFysukHImt9x4F9cyaReFCL+BHMexwSTrxtiZSq3KbabGLYXaqrR3oZxEE
nEOTrHgMsVDEszfTKJVhVlFJRfgb+IWqxeMYF8eF/Hd1qhrIMXMWRnwq4H+9/tpB
XIlFXagLe6KzvJLZJz8MAl56zqV3fgHQ0LNSKVLXtfLUHG+L/d7cvp8El0dUUgkB
hPytEj++0uVKJZdXq5qQqcm5P+YyJXfbkYFauNelFPj0u3nua30my6qI9Qu7KDNB
sQ6KC+sF4qosK+g1ahQaM1mQ+lUqsgbbRKbsnHjgCxZ/2vhikqHjjTkO6ME4WQah
BLaWA5PAq7AasqIjY0fCOKdkNenY37xeLpousFOWR1sg8VlUfdjEO+CMBkpjnKZ+
Z4KC/B6PPjAf9IzdqRJyGqv8JBZhkoT1djkmSQ2QRXzfbbKa7joScoJEK3vBXRLq
ymJxXiMq3S/vfvwC7oxUKRHr0RzUe+GKM5FqnFiVcDPDsI7H9P74BNvWWn3/Nj6r
q0nIb0iz0xog76oT0gxvUmevQ1DmKInoZ+wOZe2TMkPULsl9DvpKOnh/4HZ3EoB1
VKMrBISWmMudLH1PosdC84tMH5Ap/KvEIhKbxhHJhxAxD8u7IkKKX4ISI384QebD
ohGFwz54wWGlVWbRnlGE5Z6Fp1cRAbpcBQF2q7a5KAhzs3KpkeTrRf4sPaa3vP/t
DGOfTshvCNSTGJ8O2FI/ZnTh26Aird1cyUFqs8rgLU5wp6I4oY9AGmyCybG3bW6b
ldn/esz2I6UB05HkFgeKnRQWlwESY2hmh06p//FSeKFmIRjTXRfB7eHD2ba6z4xU
HkCGowODCsmlwHFLmhCejaZRvFYOfGPkIxixQ3eU7trpiFAii1f1RFmO4UJZPF+P
WToNJHShbNCGow6803pcPRMSqSHFhsNM4zn+NYhQF2FT5sDXf85F10B1BGCxba92
pzS7UCq/HapV9r59D/O03j2wSL5mHzOzP/8wbm3SuwOG7zt4ma0GoTjT3PF2jbDC
BNOPwFWAED0IKE7CjGD6YKVpOE1XrLkDIu7WgnHg2YudSkIj6N9pLc6ognis54RM
YxvJwzAp4Jqmq88p0vpfh1kN2kIWdFWf5qF9omXcFdSmy0QuhNuBvk4GjwBjlqSm
9ITCpbkicybEJb/8qRowlJuLmfiW4ALgTvwMKiD7FmW/4/G0BH/c98Z3CNn/KcS3
S5OKNuTJaDNz5tUxZfTWCrACtvaAr0mPPYuChw9oyFHjIY5PaPcTs05c/H5GpIif
21aYeEzN2y0TMlZ7Hc+gVctEJEvPSOP1y3F5pQnlgvluTbqdSovoTAOTcCmQsVI2
hzVjygp+/KCon0UL74n0kep3sskSzM2gBlk9lUJku9NcmRrO13l8Qnp3mqToBCJN
pE0NemQdqqLOGr2QPditQHdVJyeiPFQWSwX5jcajaZWTfFCp1zeSKy4bnN4FS//c
hOwpmZrM+jS0T09qTxG+3oEnsSDVUXxTIcrsYzRdMHSR7yNUVQOp+QAfHUH/dkFw
8hIBCpxBGrqxKwxaUldPdXysqJmJbL98m6kJaUtBKvUkJE2JpAKOH5lSI3uIDmLH
gt7GuZBQ0Y1FoHUj6g9yPrI4kUy9qQbVs0F0BakEIm1yaqSKwSR6VlqWCLyUXIx8
R6NXLRMLjkSbLt5h25bkTSbSQxp4ICoD5XPX8mB9o5EwS7xXQxtAInlzXtCBOsk2
SbviwUDkvEP0fH55xeiubtFC7tVGcu6uZtP1/31vFytx0q1bSDPAV4Z5Ps1uhlor
MI+OsnigvKqjQUdTLQ41g+jRUpIrKAHvvQXnoG6jN74bA5vOd6RyKKHOSsPBBHpH
Es3ApsPzIULnAoZyL2TDIQCt1T9SFCpxuGr5kNTG7MhVS1zdICkOwSp36EuK+uyH
T4rBfcqrgfEGJi7GGkyO6ECTBdwPYhQiZ/4CbA6Z+J3yV0Nwu1eiSgAvoxGubh9p
qmzSHlIvBGMUSjHmm7jA42GXVtnX9rb5AKtpYUHXyWKsOy/+SXEi03r0iAj66kSh
2cRFIIc+CT1YOfmCF1LjHSdGzGGLbNsG2PXODRUqrLqtKmfduo/yfkkep8K49TTA
b50oEjMKOzgaSu0yzWLKfoCjIVju2AFljJBmUtQ51RdlsDkLflNXX3bzK4qr14t1
Etmtm/BfkybMZW679HE+/pysNnxBiS/mAqoPKYqubtTUTxr3lvUE9pCINt6w1exA
sgqjyAMgkwsXzJs77iDaLR6xickBbxRGmoMajvReYOXWBBnpFhoV/0xAPtaOS29V
McEsvbsvse/WnvrlxShTc2OD9ATMAZS93pdmmz+C0Isy5WycHC7s3tHuNRQiRPjk
rrylVmSDfAbjl/3bXOoBVOkj6goLhzsWX7dNbE4khb0oxg01N0IxpZSiBHiIARLr
RR8NDmyBuxlFgV5VZwHyadqxy/6rR7MabTwjvT5qqOgOjdFjHiL8y5UWj2V3C146
SSYfNaWRkC7eSDYIKtrOunlv66V5w+6pwvBby3osx+TTXZUi5GqaIobqYsKm5+Jq
5jRp6NB1Wjdguyv2nsCNmtQ9wE2Q972UMBsHBUURbdQP2q6Ey/4t5fgxAWwST05G
0M1O/dHXzCzB8gL6H51TQC+jI797NcoFiCTu3ugG3X0ZENirRV69pmHSUx5mXi0K
qoeHgLyrSn/9I91Jy67ju3X+Hs1zgC0pdrIixPuX9ys7S6yZv6h9XjlRZh5/h5zn
9VOPmkSqdZtuodPMkDjHRQEap7beLmi6tASe7slTv4HZ+qF7C6eulJ/f6ZsmW2ls
q4E5V4bke5BcQmUT9AuPDGNAgWKsHkta26qgNvEHGsa/eIqF4yFr3xKOJgtV388U
l+kQqiGzp5UMUF5iewG+S3/p3jYKEzG5R3wwvsIfZOfO5RQ3PeYrw/N10RYQ1VPV
qbyXOwke/hzKFPgNDPai6Q4miITgQEwgDkxMWS87/dRBFDBBfLSDJ/vknZ8mBuVQ
bTizYwYVj6SJXBsEaydCS8Bv9FWq2Hg+Q1/BsWN3Y69vXNibhbeRKrdtohiubh6J
jKyr9HyMtSd9vakAY7g08Xm1LjPGs/MeZ0dqDYat9OO+0EKUS+VznNaZdrVduaA/
PDEflAinuK4FCEeB8+lQUNp0WnsJIMffnV/r4jfgM0jY/koRgXt0bcin4aGJp9m5
syWLyFHyJ3rTsyUR/j3XB+rVqbJfImFfp4mDMNBIkwUx2lICjIikO1XqzavRMg91
akodbVQIObbQAVTYI/O9V2cZIBVev9/LvZJzcOH90oJpzKTfUU7JjBC/V1xIPa1J
oKQqAsxuYwBCPdHUCznXBjCldawGoMo1guzBH0G1xsjvH1uOMW93hR4375rhz75o
AhAy7rwAWxSVsD/Wfmxmg5WCxDTS8H/aW3S6cnpfIYT7oDpFATwrSf0m+GindilY
bYj0znIGzgKMilBV0ikpX3yViQ5vAYO7PnuIjN84kmXge6MFYNKI6Y6ofJO5Llce
V0gKIFfDekPCEaUxkopTHSJLK1pBlCfe7VXqWbDiw5tjc50Zg07uXzwPbbQOZMvQ
eX9PcCwMEftkp7nCEO/7VY5aL7i1910qcg9pnQFTFMDSI2XpLerx5yY8/VH/tlpH
4ERaIFWrLraKtbnVaJs/S3uNWzSWLRst1/OuiEx0O+noTWeaZF+1SAIeLZdGIFeR
ln0MVPymzbryBWh29cQRB55NoMbnyv/lJgQ5Y1CXSPeHZz+ZGzTyZK0+C1/vdv7w
kQ+EK8gi5Sfk+Hluhz2R4H8SJ8IAHSauBMfXhRuhDSamPJE/2dvSKC2eC3AfrkZM
qp8MaToOPxr1yB9oQMYQarNaDMgzsUc5snh9CuPfWiULsubwSXnT/421+CeUVyHP
1zD47TzNoyT+YDffs0B37wSh6spCqmpTPt3aRUNekZR+kQnvReYk2ZeY8gUxrkli
I+tlG09iWCnDvvOaNhkOoldSjv0pTGIJrX/83tfKNHVo/Vu79gQiuFzMsLseqPTx
SX9RQ/lc7rI3kjYpb74hSHdQAwBm+Xg6LMtVgDFjUtAadoWkpqh2QBousUAQf4DB
Tbw18EnMVrQP9+gUgJUaRo8K3eORK5v4J0trMy2eUlDvGBniVOxwOV3PSMpWzGgX
+T6AydTjfrlRNabyd2lBQIIm0hemyzWWJnEWhSUvXlyWJPtIJ7+/3QCXjcFfEPe7
eElQpUsZzYC77iaf92ZvOjtwjPCgYE92eO6uLHH2qpO4zkbMPqAENXSrqiIQ6S5G
HZk31wLRVrT5wuTkc5c/0q0U74YynaH5MYW6xgnyBHk1KCgS7PURQ3i9rw8BIHM0
9UGs4zA/X7rSVC/utAvnMQGUsUT4dWGSPlKwk94aLKXumq7uD0ViGB9cenz3+Vpe
G8DwgaIyGHQAD65C45SHClJ/a6ctHNU8Bcxw3XpAxFWHxGK4lNwuu0kiSxLcXels
AS/d3fpPiwvSDLUCJT3gAZCkU91We2C/0wMAP9g3w6qTQJ4Zs34ZU5xYKlu1HJwT
psd+zwajO41WWwDj/rizQvT8jgPm9J6pA0IJ6/eAUpGOhJy5SmwpQr+Tuw6Tm8BH
wI12uC9Kz0FKMm0ZN53dZO90RL2z+aGoLB2AhUqqqIhZ8GB5IzJ8rYILaGSqRJ0r
CKJ6bY/GzWuCzutjq35e0yu1xk4Qw+pDxvWDOAfOi2nJ+l7HhD5yd9MhJ3aYjEJK
ZAz21CQ7cY2FSPEwE9P0edgo7DYITUTB02nU3qydNTiA1XGWAWokQ6NmYtK5Zkst
CRMC9Rmdt0ABV4WYqm+Ht50l0Xwm9SBtawJBvSpWZka/HvDIrYZcLd3mvodsfNdK
rV7cHUWsF/VC/IG68SJZ+82WoQlxxc64yhmphf8vpltSWQJ4obi6O0bMcbSkVDOz
3FnvHtIvA8r9GsDehTDmn7svvb1JbS3V5P9XTNDgEJTJhe16uyWGF5ZzhjCaYylw
yVyR/WvvJJbciD1EagcrUfmxpNKg296P7jbMLivBpLwKSymvoy1hyIZ5adX/qZt4
6yEv5wGTryLG8O1KRqtin6OyTYE5J7I42a8ER+cHXqo2fAj6zeu02RHpC97hH7PZ
haS/1tVNibMqs51O1A9oJo8r1Jg+CkV5MnE3XZCgVf9pWilNee3l8QlAzCGC9xEE
nupFUCCmpEBO4RN5ulJFFBCNQ0467Fmi+cT4imRA0Cvk7+4snlXmyCEnRfQEdcxl
lKSd4Im8puvtZ68z/YUcpeG6GRyhtKA4lCXTreuR3FllSu/1sEdv/69nNWlkAPR4
EIFkS6C+D8w7vWfkArdCgJjoE7MsNPf/o25JDmMOE0P3MYHkS1Jcm8KDfQpOuEqz
sYv/dnAQHJB4wNCqwUkg4u4fyzZ4lcvOY7oRKCtHXsyXAYGZBratzwfIhvvJbWUM
N/dy+68c2YU2s8iG50HoO1CDzak89x5BKfme8RvlyL2jn7O3uQy9KuvQ5bilM7SC
f/0sTY5+wK59eLuaI0Rjq3VuefxDXPy+Fz/k6Is+wkGRExzsJCyj037/ohEpubom
Qtoe9c+/sGzr8RcGW0UvZtvN66iDwJNrFKhIvwkEB43ffDGwyp88rcW75zkpZg/P
vZ3aKuADyDZ2ZxQ7RPhC/dlBOV40XQbeC2qTcBUjGScwt7DOgUIDmwC96CLakpQl
5DrO5LmMBa6yxBs9G21D3+yYSfIJksq0xybK2QvKuk9xYn2M53Vw7YMSDTyd73at
oJqZfAOp4hbw/gePtbzZ3iR+Ino+kyfh968Uleqm2ndzh1fWV6p/Fiu62s89h2oa
V30cEvapW81gM17fjQTSUm/v2mIgzNCrpeGsRpN87M+yT67xhirGejF0x2Aae7Wr
8IBtmYTlMeOC/ZRSvG8gXEsJGomOqyA5tDVtaqbFko9dbzqzNjsq8V/VZ2rgXMY2
2+sYqfRqQoTHO4JwAyr4zqmwera5hER1gxWh8NcgkCHJ46bhoPbxXKzUqUW94IRW
z3ep4+2VSjNX5XY6wmg/8izhxWAMDg5SrrxB1HnhTR38r4O+RvDRBTpB8kcZv4tB
099u0p5SNXYim610Jssuleh9msY9NLx5cuTKgc8HgVBoRWu3hd0hl74381F5VKzM
3uSNTj/HfCVtP69x7nufA0rOkJCxl3j8iNfQj4Zqhz1kfaVHcbpx6kZzEmNVfN+Z
RwfMTuP1vYKl6h/64lJZvpcTHoUNEL7S+F7+NeB0A9x8uoSDDiYqm5bGg2naomBe
I/yhV39uytWbOdfHBpb6LhkXY12XIYAdnlujA7UzXHBb5KJnpz6PywX1nomEinTH
qvf8jjFre3WQsn3tnghlUck5N7UehbXqC12dwJeL94PtNIBmxoEM9QcsNTTiBvt0
ebmHCJm5NFKSbiIPXs7WMQJT4zBFcauljdBp0ZKhmxFk/2QjGDsJTIJjYbX2BVDv
jBnude/309Isoe5rOmJMrT5uX6PiE21+VCKB44CWp4P8wT0sNqndr/+nzVLHUQjK
PUfTzlwbZE1taD5RLGYOHldQ33LasoCrVrp6Hf7rU8oQDK6FHmabcE733PMUgCub
87iRwlpUaMbvsvinwf5H9nK7jfaWU2al1Loj5QkUrg4E+ocRTsWPunDTgPZJrv49
vv+jZ+WNWbmSiffaM0ZzKTisaygXx6ROoeGxjyuzZouOtMdCQumvCefSgtBhDM1y
gwJF+tSNq0y3tnOzH4H4UdrF85BWGEBeWbxVQkb/i8BunI4Ll85YWGEWiwxww5he
Z6n3EcbQ6BF7bfXe0/gXWCQQpVKgXPqUEH5Ksbp0vhj6mqymcs9O7gqAiHiJ/PKl
552XhRXsSdYBcDw8fbmAivbSC0JeeS6imnY2HS3StzO3UOjmi6pEZhMb9qhSFc5X
bSYBicLbBScURhhcLfXZr+Uu0bIKz7fEhrkA1XUVdWzEGG9+k2MzzDGSnITtqRAX
EXm+T2kZWOG5yVu3UAIXkyUYn/o7bv8BfskMoieemsc8CuFzDK34/IrodjXnpJEI
Z5todzKU3XEfRDzQ07uU+38pUr/H5TwxMb9+b/xNXNwl0r0y0prAUryMZF2clggy
C7+LjX68OPiYYlyhMff05g6Q2KA7Oaa+QeuucAHvtVDwVDbeDszlxazkew5CUdKH
4tykJ78sBRORZfAWSaQbztN1S2J+TSj2IyfEV7UGlnCGtRcopymO9MxQsGITUNvJ
UNy0/SmJ+QKwJooZEO0ytp76k/uizAJyaLdU6X/6NcOShpKZLu8nuetdSAzMHPnB
95Z184O3Bk2bvJkGaIfAK0zifslSu92mI/vW4amOIDn6A1L1vlyAJu5nUprMOro+
gbAxS1by9auh/WPPJrBoqLZbU2PRP6oGcy0sFz/et8VMZgJ8/ZIiOjdiiOCTGkee
Uc8C/f2PAijeBqN42GT2IKy5VEPKVuIyLcE6hsCVml0F3ei3/HfKXnLI+p5H1ejQ
KJ680YE5GY3QH8M0DBUDH3s2OKmM+jpsix4LZNDA7nXb8xgnHmzzu4SV3QhkQX67
bishcsTL95idRrICi1RWExSzXKURIrgY7vj2lF3ceau1M3QNK1hHRAJRPdynkj+I
1o9//rKUTPooOQpTjGyWCW0foJNHpaXHlZq6sOOB7fFMjJCd+wv33aZaGnA3MXOx
2IJJ8Q3ysp5z1aCoDzIA++Ay5omEeMU0oLIRZOhFOV+ey4UJ1fct1dPlUmbzhogU
57sWDrY5fn5cczCwGD/b4sZTLRg/2dW47lM5G0K2OjF35dnzcFN5B9US/XFfdWeX
JwwhceDUg0qEinIjCyKqSUZZNlVRdeXndbb3gypqBKQynBkAwRI61wXu2KZdQrf7
uUKpv6araZbV089FuY19nwb9fLMJSvYlyP3FwSsArhjHpcWrITiNgRm+8VXTk0nY
r1ObMmQEC18M3IUdef7kTiJz83O9b4bKsOc6HFLg2e8dkLXUW2upYwLAdhOGOvxX
jPQwjjoT7bD4qzOEQF+mZLdgOLBpMBLbIJ1AZOYHhKA/TUreqVRfE9PYt8ML4Jxo
fM7qnQFoDc41ITIZl12aPwWqnDSFYjMvY4kO2Ln5hKk2u4/6zZtOqPSdokQRySPz
WGbknzmfBTtKsWGwOt23R5fK9drNNhB+msNpllXqOWa/rddLLfBtPCu4dyRnj6mQ
t1MvrfHRQIwSyNh6M7YXhXQ2mxr7v1opHHXXSEKiXRQthgPIVhmLoiggQK+LLynq
IrgEBYjH2YtdYBVuDqEvMr1WptOjF6Q/HugP96BU8MPkccPC33ooLNWI/7zjK8+N
zB4YQp4pNpra7N20sfprDYTBo41y3D2Ma+LcMWbngjwNT6nnSLGl6gnvKn1mZOZG
WI1IuT7eVXrF6V/tqrdR3V1vaI41FyDXew3cjzoU6vnPhfFzpVcDPBLAenRYx15i
CvXWwHhXLMDyqWjwNRX7rqjj0NfMDpPp6CIQCx/HgoCj5eo1CI68toVbTFtYREBW
tf3/TtVk2Aj+2StZLLGf9eQe9bighsyedG0MIdMcXUhz/+YDgVQleC6V5O3N/ST8
Lb8w7mQHiTwobgjM/PyEzEzgTaC9tXlemzoWeJQQm5vtYH9FAIhDih/CLzwo7foH
231RESVnAQABt/iK6hj3t/ts/BMxSPoawNBaIVw5WCkKeyBXs6O8kUArRuDZ3L/G
kZCa+q3cSkvL1nkUWJxuoINik7mkO/Qwjj0lhuCxaiWz3hdM2P5tXLsgFFv26zQS
+5flRlIt2+KL0jzhU6Tv/35tb8cxkMJT/Ah4qDfnOx8KIQVWT/WnBvvkhDUk7nuz
TWRixP8RHLBd6MRProiC8q2jTMDc4/e6JwknY4g6PPljyjVrBpoHwIUcD8c1Kx0X
HP9uSmXFUyvV9WN9M0MluFk/13Ymy6stu2K2V4FP65eHx9c6MVhYOuv56lYygpOQ
N3hw2P7UlP0j+ZNonxu/mWeytwE3x65pfps8N+dV+734ngU5AJR+W1NhhJPuCgH4
dAvUULnHLi3t2Xug7TFEgGff9L573/ORBelrG5HISCxcNpSjM1CX+lVM8A1pMcvk
5PRN4N+ZjtVcL2sAPP7d3pFIHXFacVg0h6OrtVP0rKmohs34WebJUMx74bOb5cCr
rv3xOY+/vcl4W0omgPa7GObZEkEwfCN7dnAc0E/vuGE0JCN692nJT5j+rE9P9q7m
95WmjZU8qyliiNp8jkvYtsRgv4hVcGkoPDuJyuuVNIOobRXHYz3tZ8SMu7696lmP
cMd25OSGsc/hTbeKNLQYv++3Opo2Flddm0EUA1fiyvMQ7QqplCyRKYOpYDomnDPP
ddm/+Tqzji+ACw17IXJCM1jMbBtDY+MrhC4QAhr3eqOpZ0SHX0WlemzDtDKsizUq
33ZH4FMGLSPfn6wByGseaK40tG9mlev7RVUBUYcRnLwtJEnAXHhviD+xG67nChXZ
POuLG62IRyit0POkvoRQ7XjW5AkKdtvu/j88uZjcMJTiMobUnzQkFeaRhkI6bU9r
vKNpV8raFHLiQ7JeG4Q4xpeo6dzL4dDvPA4g30/d8gfXSOQeGnBewM54StZWC5at
cWtUKWl43QJxc7s5Q6rTgScnKewyFt0yjkc7yisObxV0qJAb3b1noLk6X0hclwZF
cmy/vwJLcLZPe4ze99FV6VwZNmU3E3ub0GUX6RMfazkCoaC9Z/IgnRn7aBqcfQUB
mQmGc5eySn7mxpbu+VKOSfBXqO5pNyiR8w0wjHtIl0iBoILlYHI2eqJspTTVoKQ3
xLeTVP18sSs6b3xaCHC4ioGJ+Lg0a6EqEzNQJRxIx8ZOkRokoD/VWu/wrZJfvPAF
X3Q67HtmZvn0H/SgVZPPyq3dBbqDPh17DVEI5/1Iv6CMTOwpWQDOyEKf1zlU3Aky
K+R1Byix//Md3EsSIEe37QUrsi4WrnoAMx7Tzml51v6+510PxapXn//jhk+NkUDr
JYXDm79JcRw7VHtPlovE3QcVq2dCdG+vIOrdw02XdByjaMihVNFRJvYOa8ZD2QX6
mNueH2uwbT01Jr42JAU2wJBCN8WRHjIAWi+YwPXYL3bcgtxoSbdCHvS8oabZkAjk
fRuQZ24H4qXQgOsoKy/hhiP8dwf2aVUqh9GBOvPJdYDVkJzACfmUDbXz3QDXejq0
Fwrwt1/jcboWimp1LyAMjKnqztoTJYXtztBI6q9h7zsK2EJHMGuu2ynkto0D+hb2
KjhIzrwmRCCTLDXtbXZ8/jSN2i1h22AUnsBxTxUOtXzBJng6ZXZaaiHSf4a91HML
QacGxKbC4BoFmFY1dYp0zXd0M2Zv1Y1bnpMQRQpgoSX+Efhyo7hy5JU17SWkDARg
DfjWQEpMTsRTkDBKuZfauQRnqCjdV9ghqoa/h78K7kEW56CQyTOah2y7I20X7UWU
2xc1RvtChx7NXoBSMoRh0OryaewkDiZp/UI5ozAYmbgYsu42DpycT3F6xVrEV0cu
uBpZtQkFV3oSRTXaocfoXpuNy8vora1/wwra6KRyeaoYpvT2MVFZJqeSOu6Hmcn8
U5dn8MomTFdhh7y54jHVa1CzEKxxfzoHLVA+KinJsFT+9qY0q5UtiBijuJiuxLtt
qlgqvH0M5yW5dWvzxs+qhARrDNYG32XA21Cuh0HNtnISzMxvzPADMAVt4dLDDYQ+
ldN6YuklO3PxHbV2iPgMEZcCJvsY3F1MyBeBksFoqgi+sAlvW/U6DlbIbj+CyyIR
a1AebgDNfdciiiYSEmYnugi9w9R+9ZjENBr950aO3lfW/CsXe3U+pwTPjwMvmsmN
inYxY1QfDwGN20Ar4sLJ0dyYjWpxYCIin5T9MtWvZ5YLU/hNErEkXbCds93lbjnQ
q3HguOlxEcj3UlVIz4RPdzdmSG/WeidSXjTrd+QQloOUWL/QfhlogOWoG0mOmtg0
NACYNcvjKM+5p2P1YPonTIlKWEzfHb5ndayehxGnCSd7ALOPyRvn2sC6WNTovKNg
fScMkF7B2E7ioPMIIIAdSaKKQhStNg9QfRkUUZDKl61neImZW89LrH7wG0RPX91+
PaHaFJ/kGRH8KwUDsL16RW1gdUQzfd/L8LLzZtXwB2kgrKSkqBWnhznhJ6eQOF4d
q3HG7W52o/GA42m8afJ82FIq8wWaYakcALMQuPhKn8K1yzW4UX17ILL15uMQ1B6Y
9fD/EsWeeQIMZZ2Wc/AuZMUQLfImbBizrR5XDih8z1ysebJIKTentMGsu76UyDX1
hoSxt6nHS0qYhCbIc5KZubnHVQQb/5luosVDKUtJVYEuZnXnagQmDdKq0bPfpt6Z
80mal9lMUyd+IC3NPtDuLLXBnwkxgLTA93TU+U+k0ACMAYYh/7YsJa3QaY9U/caQ
dpITlDhNwJDUXEFN7Di4f/xzDH2L96Trsss/nzFf7md2nNIe6crSWKfx+YLok7md
O+fiGOG4TOx+HIrFivJx8JPTqEQD51gplSVwxsxi6YGFvPWwsOvHSsZGf1QAs55L
Ip3v+qrbGJYxMHEA/1uQIA==
`pragma protect end_protected
