
module ax_issp (
	probe,
	source);	

	input	[14:0]	probe;
	output	[8:0]	source;
endmodule
