// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 13:57:46 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
hSouPGt1odv901jEPtojl5szqNgSZjc6A/cVvqdWGKcRTwgOeLc/keX3+ylNr6x+
3EVh/7HGtXn8oYZlwRqmSUZR7B7JjPem+9vEK+8JEVaArfpE3/8isfYwNZ/gidww
cc/l2ZqLUr03uHZAv/ZLsQKpSPWQ97eXZyV3s/Lv4sY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 30848)
hUUMJfS5iYvhd3ULuRdEwQJp4S88gOZ6W2bUPY8pW1W7d/ADxa5YRY/0BgJLkY2t
9Z6hXEOto9pX/sEJ6lpLyGyEvRIVwtj2E9oZV/ObQ6bl/g35nHI+kJiTAIPXC2EQ
T0qqprhf9i0XOuEpX16EZUwi6ZPzKjnGol4A5cUbxvVz1o89zngTy+XMiEkCJTZE
zsrH7x6ygzAllWhwU7BdyP6hUbAqcDNt+h7Xa3wnAiFew+6+Zps24Ru3u15pfc54
W81eU30gQbGLHVzgfy7g1AJ+XCzwiQeyGuMyGFZ6mE9RjzWB0bnU05GnIINvK+OQ
A3E9bzFJ6z158wNP4sOBUT/MSPEGJQ4FU7RlYKSzSF4i12d83aR/1nh9liNDkkXN
mLyOcDSZXgSVcaWAogAcLs53S7hd/N6ytyepoEuKK80SjlUCguaqYnOy3ouo/GiB
IkDQrPDnSc3KYs7iOyiteuSWwKBBFuOV0y09WhJylO1Qf1nKVK8wB6elmz08LsG+
SmyIcVY/UiB1Hb8fe/70EJSazml6/7UTAtEqgA0+9P7Z7Xa9St8EuSLIz3j0FAAZ
VWOTWNAYXuwjr+RzMQKOZUO2CFp9OqXsB3Z0ufi7mVYt7DwT1Qbdm7zVt+2g5go8
SHhKB57fcrHoJqLQ6jvPY7z46dQeKdvEUJmXHXb/n++sqv5NUxbIkiX3pxvDPx6D
uVxB3XKXpuj1nWppDJTGGYZeJ1F+++HRy1/WvkX+7Z1h15WYgjQCjK1T90pzJba+
MCVrty9NonuWF2kE4KZIlxASJSKExWGbui1mTrwa5f04CfRssLIXjV/oJeiR5BC3
CdEixxDUTYaeyNOJ65yCvwJKnrSaRMmjeFplKrrJ+vYsQO66//2dP7bwPDL08r+t
qOe3eluAZYoXOHm4r85/Y+cXZQ0x8uatnY+/ZB8SUnS9JLrhEqLvZ8cms8mNYW/w
C4HxVdv4k3gWYTeCVw6aJU8fhJ9ZtW0VIhXYYlSTkxbcRtWuTHFwUtCckBChRGWf
/Qatmk1OBYhvTy4lL5PZaU8JwrDGi0OuoqpwsXJ/gA3oMSzekbfJohOY7iOGyCVy
/FBTWHqFokMXyBoKWG3zVTatAC+DdeEezOG6Tmsp5A7yVNk1yuWoG35clM80KeZ/
t1mefBD/i//xTLQbB8GDrWmbRa5YeRmejYSlc0EAva4m+g9v1luZZltTi/Hd6Hxs
c4RppDwad4S/qNMFwdT3Vql0kRzu+eEnxUrrQwACbheLLi/30gVLvttxhMhxH/LK
7mNF77JAZVCSLaNd1JYXZnsZc/1nK64ggxmoTjNF1a3K2f04DQ8ypBDRj2adk4za
492AlTDKtKJBJrLZHsGZ7xOxfm0Zypjo3KliNI6rJiJ/OPuri3FVOYty7/XODeOx
Ahu1IS9RFTUMOGyU7VjHjyozV6U4qvR/TVZkddQ23xgDCuYLwWPgOs7vh9DGEAb0
JoOjOCjpuFgfTA3yvuYYhfc32/fxlp0eW62oU/D2acAxm8q46Lu7K6zAGe/s/9LT
Dr+s62sSLHUPN5xf0b5qFo40NlXuO4//4oIathIeJd8ZJK/C9PLNCQt/0oo2rsaW
iJ8B4f7Eooy8NDWSQewrmBuyAb3K/hBy/cb7isZ+fl1KIm9CTAiJgmxlLlKKEJkY
mzKz0iR909dRc+Ly7io8qr2gCvTCQm6g4YWqu3nc6dR8wSPvUOavJLPsWXmFDxg9
l/KPCyGYKRNQgaQOSlSDx/r0we4/KKaNksTNP9Sb1iqJqbknMJ5+LvOl8irDDyY/
/iF7AsJqDjLJIzYzKbQIXkKndXxcxi8n5xTndWSww5mjnaN+L+KQ1fBENwXLx2V0
oq4LCQAq5oRowYP5m2CnhMmrbbKP6b8mnYm4QjEbdMNzgB78RoV8BA1ljsUOMuvU
bilecIug/3lVcLYSJ+U29EVFdHqtG578Ndugxw5OqBZfpeJ7TexGdNae0i/foTIP
2ykMtOJARKLQuBtJRM9+Qz/txpkxVJ7G3aFpYaZeO0PzFzh2k5lkhFTPX6yjRUV+
zpuIeaQxwBhhJ+gOTLhG5uOGv1wrk+SiE20ldMtAe2z8sBtkYLxHalKYZO2+2dS8
hF9K+lkITaQEOfScskXv8STbY2lXWS0Na7aS5FW6NUIygl3drKvBAlm4DgqsS13r
uQG933qWkvYwrPZLVD0VHFxRJa+vmNbcNEnYIQUeaB3M00fzIhzq2ALIsrm0VKzx
zpCoHJLKFlAxHCEWMMwdQvS861OG1l4J/DANaNSv4y9GuqsrIuS4SzGYQHZZxq7L
CIkmlQH4J7vDn6DOGfZfbAuqJMjnzh0ZUdZq6q0anxKcXzKPT8F7JWLaeR3SoXWV
tev4sXZQNeUeLvfHzIk/9wQcd67pv/eChtVsVJyFhcWsWSpSgOtj8XkUaUONFpqr
3LA0SEGgf0U5907JTenEqtcXr857KjaJ9ApwmzPIXITvaotIkGD5n6FzfE2kX89s
6z5TbZjOaZtdZW2aUoSCQ3y7ts3iU0hc5T93FUJ6pIYdstjtxVTl7GK7YCs4OMlO
orhrvRab6jX6wMOzERAx4bvDmlSPLRTbII7vaLW1nrhTXoEycuEWiuSiFim7FSec
4lqO4e4wdpCqaY0TwBY0Q+0CzLXBwU4Ky2jnl6eEwtibAIlJsWq+qQslj0Vx3Q1B
3XOVPtQVRoFYDfyHjFnqYTc8B2YhqltMV/Ini4t6SVAdCaiXUcs5R0QNsoFbD+gd
ywtmPfXrkYZ/I/i39iGB1i7+ZNTWdnQVGwt+UYnrhkYCr8iT5V98nth6CKbaovXs
efA9S1mDy3L4+Vnquem+PR+B7DmxeZ3uV0MqyWb8MKbh05/Pp8PP1OAx/gysCdqe
7XhHOZ0kFiwqHpLdSmKIp1X6wSz0L/UfHiPezniqWpEhl/q1N487Sq8nObEQr5nV
m8qPnUfNG4TayrA77AYpP4aVBaXpaANivP61aQpotu357SsxUzNV/YLhloBH2hhb
GNK+nDHRlt0oRoWsTJ7Nt8xbOlHQVnxKMM7jGbUY/2YVnIqa9HHAoNMCc435Gqy0
VPmVqdoQy5UZLnu0KqaaWoXcWAPhecrOsoeEatsyrwilRNrw6xjzTsCiKe1r2ApZ
t+WS6BSRQWaVDnMpfWdfFvMlo8hEKk0ZJwhf+4PiZEvVvwn6c3Cx9g67L4j5T5EG
V64tp7loSlHra39LyuK7QtBphqDORjYw6yMAK/LLGxbzacCz33n3K2RQLRAr2qMO
OhIkyIsTHjyO9qz1aq92QlmF2T8pR6LB7+MiVNAlMHHFey//Yi/YGhX5xa1p75rP
+w0pUqcguRz3kzzO6tImR0cvNUR23dciYFwV7FTlidnPgvTj+n1mvQKTh3B4Y7Ll
u9S+GjiNbwqUxWf74SbrOc4zzdNY7E1YUFru74Rds3ZWtc/pivvHoy9zCm/cyIwa
+5UuNHc3f2Giq2uBGFiAqrIAueyQ7UgJEKk9Q2pHE98olCGd8e1+/btc5hQLT8kh
h+egMzABWBsHXoQChGhQaZGD5ldtfApy79dHk18rF9AX2hVr9ZgswGECL2rBsIuH
X0Exhs63Tc+f8hsQKzYNcYb9z0XYHW1w4ecI9V5qsQCMELbUyRSAdy/hqVUsXPNw
SpP9pz436hNBQphTgVOCgd9Lb/7yptDfJzNfVlIFfzMdeq4iP/R230ONYn3q0Fqg
HO+SGsPkitt9UF39nYPoTlxzlIdaVgVhCAeN6VVFf/mIiU5P2eWYl2v9vk8Teq+F
/TupYqCJaMLoazcIEvbL9H/Dv3Mq/KhMzNqfGKlNIWHetAgnDKPwDsr5jlMoF2PC
CJO4PVOdQYdF4K5oVeCJbZEAHyZqiXTdm5gD8ldw+nt+FlLyUbUES97lDp3+DbHI
DzhmWDf/cYY8wPRduO6xJaGqUtwK2SulOMusSMliBMS2bgSl5+hoTBNYBwVj7jo3
O+tfQqFLyOHtCyzld5sJjqvm6Api6acbj0VLHCGoeQLQPAO9ZyCy6Jms7E1Kikl2
MBI1blriYWzHTdCQL2eZUfAIiB9txPePWjsjwK+A29M+pldhm8dOOBIU1jLTT7YD
TkA0rfTeD6apeLj+ttqrKR2sgmHhwTQ0QyFKvbed5pZ0fgpofSd34vlUiNrF/8ru
h3ZWeeZH9bweXUakJzhQZrl6fUuTr0IkhUJMsXMaCatXISk3BopOXeljXuDGT7BN
tpTRUN6le/3RXgvzomgowYVXmTf7qWFTwQ/TwJs76qIIdSCWHyvYc54rqDIS/l2z
zAfKZWutIDLxlIth1YI1MHtHL0qPgt1lTflEPUukmjefnuxJqPUOP3eGbtZm24cD
d7FI8OzoNposLukzkqMSvxIVWSwLQYBLBYuiYrzkki8rBxMTVJ7M2iMzFwFW5E04
ifThFSIQZst1Fc7mOEPnVoit2yphrM80962/pMH6AHo1ebOXcovRdMo/nd8hyBm1
G1JWP6NjQP5n9XXL27wqeC/7KbszqfU8d93+psM28l/HRqrE3CSxZbOwfX9wP8pg
7bNyg/UnKzZvze3kDK7y0jnB8IYHwgj66W+auda5kf5MFqk+j+MspxtQcFnPznkm
i9Qoxb1mW1bTH0DlOCS6vKdB36eHNoX/3K2IZdl+bsTEQbTA4oxfutg/4FbOKTzf
NmyicIJuswLhB/Lxe4bE36WpiAbJZmBZJpkMqqMijndrkQ1RsVKP5ITgoUp7ud8z
5fK8vk6NgBWdDgv8m/ljnBglz321OR+fA5b6yyiUeWt57pc6hUd4RmXDZ9lgLLbY
awmZSdIqe1or7ki6wrQ4vqtW8hsOc3IsmeZUJXiIi0u4LgddN59Xy2Hhpo/66w6E
kZU/Xn6rGKynAYWkTMtnpzqDFa7tiW6zdICmJ1iJrzs4KyHArCfy6jXzK0rOuRRJ
bEK/0pFR9qiy5yoxtYiyfoHUodA9B+/aayqA1gkhoZ7cVkI/cCE4H9iig9KbmNFI
JSn0iwiFQUwtUsTXSoCt5HXQ/e4Hqd7CDZzN3nYHIQnscaw0WA32hUDtwQqj5wC4
4d6F5lo/XpqOPD9i3ZANQHp/KPav/5BUpV8v11FdaNkgVRWWhFP6n6vSfJ4fZBQC
iNoS4pUe4/62UjEVfrjijwtE7zGmdFlBo0RsvvragNX/BYIi1WLNrhGhBm/8xb0a
Oz2lmF3TBTxWieQdky/N8Qp7iI8CxWXEIJwQFSf+r31Bd86AFvqSB3jtHu0N9kCE
CYwQX5OuweHT3DPjj9so/USNQM4zzLdgChEd2pkDPfZ2nJhOSPuy8ZE86LRMOBOi
wKM6iQ6rZKCuwXGmoIUeczR5SM+6ctfyrFzEr64U40F+CCG4WM/L/fqzD70ZxHE4
TTSgWG25wy44DFaAAajJKWrRyzQcaqQK5C07/DNmdYzrQpJyI8XuJHbLuDEwb/pA
oidM2PutkcAx4Y2Hyrz2ktNNsv8b462rFgbyE7AZnOVuZClOBWxKErBocRUiyxl0
Tn1W3xLgkeWm30aY59ra44nxXv3LyFzn2rPe1Qahuf0TVtp0PFCS0HmZ2+tJwUmo
cjx8cFrd28j1Cu6h2qecY/YxDKQoTkWi2vwFli+pDG9m4ISZt5gapHhYKsgE2N6y
tw0SvP2ykBGAKQPnGw7iI+UaotZkjJLs7p3mbj+xtBYyrkxzpYg41U01suNh9K9R
gcF59sn+TkO/SsCPfET2UsBlxO6ZYrTX87BYexIXkISKZY+jFMGX29ltLG1UHgrO
9hr0nrQGZEd2lfqyqoXCQhXqAnCZDF64DLUP6Zaw6ekpHuidxCY/gJIMUjN9DMXx
IO3Ywno8q9RIPqKrmHRsSFmi5sBUJF0aUXByzInCwObDk0OKniRs15WXjQnXzaFt
pH1/7HbI+9KWso74WhIuZF3DYS+mhkb4cYutXqUYfI4r9UKW7R/WicFQ6B9jNrW1
dJVzecT7Miwcbf4jrOotBRmN+rIgUIJGI49q/X847jFNwMgOL5AbguWwI20UR0Pt
ljNb4BVRB+vbaTNl+yzHf6CzwbgpVZ8uiM3iZVoSjJnaTvqGWgky7aM4yxu+lBg3
PSHxh1dHyRq/hM1l4ynQn1NqfzTig0ObP/cUuQ05AOI+llJrnhbGt8I6qqz00Xbt
2ATL2P/NiMIAYegzAGiHkl6n6I3eydOVppfCyc5Cqo5VXuzEM0iiJg7059wgzrHi
9/JnMZaVnB9d2ucBwUYVdHO9fELTDM3lAMj2cZYSNd6tsb2M9ook5PJWZC3Cr3SP
5Rdi+MQg0kriOZru159wMHU7iF5XY5NSGx6si2f7dB4TU1ZuQjIVnQHYR6RYJWH+
3PaqZjfgdf2KK53R2n4NulJGliA6oBm1OBmuGThior1oddZE1ODNIbGaJAXrktW6
YpO+HdoTcODzA+i8XwO4wk/74W/slwIcE+SOjZu4XzKHT6MGiAb0sc5LPMlnsuiI
HpMy3gpAZkZstWS6XVT/RrQoBZ47cKyxMQPqr+1s5SqnkOLHFoH7YBAhykO7n4OM
DQNgjENDtTKL5vnviGqiB+XDI1ek0pawVP6GxV1veeMlxad2G28HcXi8bJzMvwu2
fQdBOWYyQG5szf5K2Y+xUazPYaxTwK3KutLnYaqmFnLW/rmC17b+NCPFdVB1U/Cq
PYOPasRx/MBe+kn+cvjFxIyUuxIXUu3HY+fBq4uXWyM1Y04nmm6B6Hk6n4pIqnpp
RGOn2+lSa64S9ZPFwE0XmL2F5vmP9y3sUoDL06jlMmXFi3CUei41N8q/S8plzUlT
LQNJoGAIjA8nYv7VB8nzZl+jYRgo6yu/CAOMV7BCGPVCXHXGCzpTVx4rYE20i5Ao
WJvBsLSwJdbMERcyOnqHG3e7DK6sjSQ9Cei8UTQpvifsHCUBzBDdkzDUDGk/Mj7N
Dwd8MM3gZBLyvAeO+DbhywaotIR4qK+5mC7544RKaLVG2s26vwDIaOxVKcaU/AwX
utp4+7hOwSlLeD542LITvfDSZCGaTF4JUmPdyC7MMqeh6i7xQ9T07P/pli08K3Az
kEgQsjpvxPk3vM3FGzu+UmH21RkluVq3IScvIsb20yyHLeB1AEcWYFqEemWxAV4X
07s4Hhvt3GYhorVVgkOICoimty9l0aooOZGc4W6O24DWa7qMwQgM2UbOgyuLl/up
xTb8RvAuSoe+O8MtCPsbiQ7oy3aMYIa5S85SeOf0g8oatrEAAbcyDVYAHrGwp5gn
kgdYQfnYpe5inyTk9yEazYYu0bunfr5KjKmTkR7CkETJd3iE4U3f2jS/atWNb5xR
aYyGwmIW1EaTXti4nkE/gtmgn4W2txTr/M11sPyf+3eeC14P29HDZ/8HWzFkPYJa
k6+sc7uYLYGF1lSkh+/oPyIdPfXQnG5KY3xNjGzsuXo/gC4UCmcEM6fSKUGxqwdZ
q1iQCFIlzFJ2tOoHguwsCQC/vReyUAJhICik9jmARiQJEMJSHyxZNwKD8ARUgsQ2
wsUAtgOmiC6jgxbi6JSLKuMRLtb4CSpUlym/Tkt8WbmoHEX0aHrueuVIdouE3Jwt
zf0f8SQFzWltGuBeHT/FRdPQwOSmWITS/YfkueejFrT8xijVUaeRHUvcUTVaCT25
Xr2LuyACz11yhksk/XO87JjHI7okme2W4G8a3tj3YI4oEQuINRdg2QN09MqV21ao
g7+0drZvJkVzq0ojCuNsFj0euw9P/UBKjC6z4oRTxJanxw2gOImAC1FNISxdA6Cx
6L+RuUvc1fNVy87PbagxVdK0EF3AwN73P7QSNcOaRgkglKTxZZ0jH91JH/QrNAcG
Ws7k1JMkmUvg+OhQvviRbwzYeJVClrfA4hU7XKLpK2I+z4N1RnZLoa/Ht8bq2uSP
Z1JXxr4V0ib1J704PyivzEe+mi0kMrTJhLvjqhnBsFgWztDQtNUSQTbmgHSp03BB
fyGkL0JSa4BmioRNLErGUGnEDwbyt8MRkwquJ48YIvj9aCVdqpxseLCLHSOR68Pw
mXpCgQCP35//4K635y0YF62DSpjF9qOl7fn0+07PO1gbQD6bXvudfORes0Zw/gum
f93XNT3zf9PHDUKDiLfnv/8oPMt7oDeEYyegO8mIYFSDGueL4GBvOk24QrRHK1A1
iAte9uI1p6VX8oe98Q8uwZkUI+QEwjXBWBH2pT3P7fPQN0EoG3HBoO3yffWZGu9T
XC8ELdlWTEPioBZBdFsvjE5/lIQtTNuE95Y3/CNb+qJArLfVk+JVscfs+JP2lf2j
OE7xuSZhK5AMjnlZqLatsB/47n2MqPnbUiXjPFERUtlHPNqPkIpD6MhH7lhhI8w4
3HkFufz/oMF+TiYFAIBJTFd1Lt023WObp2Hg1A5UU+a25bAJbQmQmWo6sY8Nxa7a
zV/FkF+qIaiYnsCYAPVmtSB9X0txkjF8rn8ZXqE0hk1gkIpayFjmNPKatMjNfZKb
XG987zjU2gIeZy3GGjJMvIE/HIA1d4hweoztFzaYoffd5XaXPGD1cYrbWXr4TqfL
DHixOHFiHmNr0NP8KwZe+O+jXJg6rOq394fQABscPZ/QOiUcHXhz532lfrIA41zL
JRizeFE9GefMNJy7u+XdAjWzzqFnrxbmickYx58Ny/YhR05BeyWiHOEjTCzK6OFg
l8tUbxFxINntnQvY7esVi41NOxVsX5ui8aq+rcdmQVq8kBHlfbW3JI5D7/6KLAPM
YV3wRdIvrnbFlenoZOGojupa+bmWro7cxMbUasPhKdj85bPT/OkdBdgXriFO3mf6
PnGVADD6iO8LqR/yBqUFf6cmnkbdjWlO4TOVJrNhxziyVa1Ruf1enBaMUZrmB1we
rv08I2H9ZYjvVmVdv70asUA0/i7Hn4RRhprqhel04EYfXj/k88tSceymovBphv7E
rABJFpn81pPZF0MTg84vut+gVoRTqzYe69RJXwFn+OYMKFKRw3gRlkVu3tjwwVE7
bYkmVqtdZY+aR7m9H5kl+sZLOtNhi5UbVMmm6qXphUdm7QLYSFucDSlto8JJh1kA
28JWgFi2LEQpE+hxMe05obhGi5a7lHKjRfhFSzSwVc4BFu02Al3azXl3qgTCgj0Z
1iYxZlErk60cQMleivt62u75rSDglUqkGVeNn+2SbdMz9a4vKz83/wK7DCNcW+Q2
lCJEajb3/hikxyZDSBfh+NFXCL06fPpa91yFk5P1WhVLgv63Phs1NARl3LjZlnnS
zo2Sq4kG6+pEhYWfsKXRH+LtNhJAd489IDa7/kEgjHSDPSli9uSdD9Wg/x8F+oRh
o187TClByCTnUUdaqFnHPaCfuVCfhufelSSahymMbSdOpMaid4QLfiJeI0ZxBXVj
LL8lhqlGRVCnfIpkmYcCnv9cJPylyeD9Ivmqbs7CuO/c4u0T7Vl5w/Kb3gwaQP16
fMpqCM/P5pg4r4SP44Emg3rtUCiI80TWL0YJpEkwkT5gv6wJg4sl1RFghtr3EHjW
9q98RMjlBZB39yMtgBvZv+zWRZnqOVCf0tM6W8c7Mr5F4eMxF5BJYEyBSB1lkDta
g6c4wohScNxymIXuQxjpSFlkKIyDM0LIsGdoJV5uKYZqQC0eZHP/F5uvdPBkeKVh
uo2svbFqyAOtmNrRkOEpbX79YSdACweldGkQTubiGR1I2iM+tP7eBajtTYOS0WA4
N4w55pM0W/u71iLRKOVGXhiRNdZ4BnZi87149FLOksFLNZzblv6j45CFQ8r1js/I
wTJgLAO+KsRNYozlBm0Ac4hoKtq43FV5hVVSJk+RlxDN6tK5+wnYUOesL0qRduo5
5OAXG2gRuZ9+47ny+LMd9+FIzvU5GvNfx72hlR5qnHlZbKW2svAzw/Tv8wVDGfG/
PtgMiJgjrkAHa+A4dTic/V3+T6hmxmn0uNoiRS8C6cA8JCqjfBDFSMhGWV7Omz2y
3YNaIGRFe0f6SUMGQMm2Wjkj27O5Z4nth2IgeL90NcfbA5qi0HeW/OTIpUn11Crf
WdNL98bbM1B0TVYJOTeBdjBANqbKf8iq4Y6SfbeBk/4jYC0UAJqEuC9JQgiNZSYS
dUuDuxiXIvkia2dbA2XgsimfVZcTngabY8cPwjarHQ0N+FPRBM+13Sb0pe1JOfPe
l59YIzr/VL2yCBvonoOsnWkPt3LNvquDu/CejfXD2+1hNp0Y08Bje8ePUDW6wKAR
kfsq6j/pzLu5iVl2rwMPmC0f8SiOyttgATGkUIcgd+7Orz2uWzei258oTJ2xPxs9
S4oCVm5+AqRXOQ4sp9XDz9NKbCCUryKLEbZqj4GXGMZS/kft+LYM5GVn3JFhDMOY
mfPQgBCNKzDKLJFcA2z15xeTTgGt/dEHUTORWjNBCvQNx0fKAWjuOO6DO+htm1sc
5yvHsgjZpzMKKWtSUWYA2Ua6p1LtLwy45Ft4p6iTdr95hmeGMKzlRSuNGwgAJOfd
I908Mm/7Qb5syVycyz2FqNtqNAdrm8rOKOFFLPUYRULEGN8dcN8Fg1TBbWUSZSPy
ixzasf6RvwwY0oxIJ8Z28eNrKe9MRlEPOczrU+4K5VXVeqsNL9c4UuhhJhpjV3MF
xEYKa0Pp95oqZyxrsM3QipNk193cLJMpj5DmJT4W2YVhlSrfJpShHfpTgwupUXnI
QwJ0KfoD1BkhhtIyDxwMszWiTjDVowdFgd0SXolHHohDidfgA8oH+eWUGNUN7ygI
6EUtMFDIrvT0TU58OmG8VplCfK8otHMwyb4mjiwt9jVTAV0lep3qHbutlrA8AOMK
lFtrgTHF6GodmVnSHrgGlGlCtk/8HNWtKuzqj+TpGDqIVICMmMnQsb+/nQSPIDQ/
imqNzrrqfdDgiCH6Q/QuDzb7wG6hni0nH1LqQoIX/NoBGuLY5RatvLqdW7YidnAG
00woPTg/G4dQT5LM5tkvcWQFn6ncG9TO+WvmvldPnWHYiAU7JS2UgKQt2HD7p2IG
YoHz3wZH8HS82DaVInrUSBicJtJQWaNJml9FiqNCRK3ubjMDhFjViz8h9T28h20S
CVTYRbvxsWesASUrtsneeKQHyy2Lr53Vf4CDGELTRnlXRgpJywHEohfYISQG6ygH
J1C43HuhBivv0XZhAz520On0Ut0onvq26f01wHdFJXk7s9rzuFXm2j0G09cpH9Og
Lyx9405grdV67gjAcPVVPna2Ajtcs6qMGRJVsoTSEWRA8e/Pk3GqXlsPT6nkJW8Y
n3kc7zDejg39AV5pXsol/VwGSZgfAoI8qVmVlznbc1NNjb9rR8JmALNGvFgkJrSh
ZcC0L0XdlEXnNVozLLA9iV0v8rDxKmYxjHWaH4IdOHa7YQ32Dzv4u67ypUNzOw8A
M0Cx0Uhu53d3Bc2iS9lPuh9Fzfi99TP9k0XWCjmK7biSJ1sGh1KjC42/1o7txsvz
IwhZat10Pdzj52Do/Re/sm0bEBPiKv+AqgJ+jihLuubX1jmgyKKevpWcFVIB1YJd
AyVgGsAKGGeF1HC6BTUdSQNvMQ9yuS2kUsrz6WSIAHm4ibIKZ8zy9ti46cVjvaUs
pBmBNV4ETdH39RhGQ2AHqpfHHGFVSZ4zyzZA55T/DbjpDsBEWqOgwrLZP7NjUlp0
FX8K/YgceE4pdpAlePEnCYtBlHTDwciHSXivhyQT7HP4AbvXLx+ZcV5iBLJ5xT31
wzbtajDLSFAKTXdrx5jbCDso2qfiHaIeISjmevKJhzYnwh7AB7BLEQ5ASEWvdskI
XvB+oveParutCpwUa6buF8rT6FR7mr9uwDJcP8vPhlQVVBfF1uucdIEjgOivUMNo
c2vPch8/NEtQBcMTvDgnl1o9adKLG4Z97sK1l2MyZ7mbkK4lkHGcQJt/52ztBS/l
iLQI0uJ6Zx46BqFirsv+T2C1K0pJ2mMcKRbEUeyyAEsfnzoWHeWdvd5VQL5pHu1u
yWXA28Wv/BxzGtWjrnlxNEUtz3ysWQDWblUlPKQ2/CEOxAYkAE8ADtT9IC87o6k2
XExFTY2GiK4B77HjpZKrYw8F2LHinRQyZlI56hVC2vyuJJdQ8do9tQoZ+bxiR8JF
avdZQMET8eaZYxui39dMoSg/tHRDdN2UEyuo9MM7vDB++l7zY3l0NlONvl+J03+Y
l4vtdgqugHM7hLvmi2oobm+MI6bys7ZBTlR21l3tj0YKypnSzq7wbVKPxUcJD1UR
YbaSTFfhv+eB0iVMpc94gr/846NoePpxz0o1b2BuXAi8RJlQhqPrl4R8goplZfSQ
v761VF2vdgEKjNmOR2KrXQ0stjOsCH9fLiBlgfzlD1pj3e6HChmbuyrdcqocTb7O
NWVVpcOyhbnEcgxYSzOg40pEe2WxQ2KgH+fa+VNGFiJ3VjssEvzvGKkclqHjP3vi
24W15qXFZJ8hYgd0wRJ8Bt61cptbo06focdB/B3US5BVjt38Df8P62qRiY3YByb+
y/cTeRQnPSD7QM8+c9/SHN2QR2bJCZf0DBAg2nSzAAmdda8oMQ102SLsFOUvFS1b
APoqoBKcMXsi1+XXGaVK1x29KbYWUhEm6q0NhtDoD59uIv+jMVuYj2vYAiSgoh7u
1qv+heAJf6bCn3+/iutNtsraURE79N+ZGHg5FiI5CsfZ28AyDThIiLXQQwXKWhDJ
TtM9ErR2Glp4psw28RzZY4fLiKfGo7/8uv0iyPB8NzjiwsjQ9bbtjE9hUoIQxj5Z
4ST3uoKZPjHaM+hpOchP+a5hq7AA3cR3qlKs/IvHppgQafYL8ME2IXDy4mDMjjh2
p2N6EJeKDokHvP9YDn9bNjwYN7dZxP7FOolW2U95kK6nTMrISTu3SXSDw7fAhEME
kGZ6Sx5j8msHEHaFZsDDXv9eaC6lke91P87H8GI/fQfUIV7Ne9Vfv0FuxvlUiGMI
uPO0MQDAO13FXRvY3WFcB+gTSwwF1J9MbWi+1P9elWl6v6AKksZJraxprrXYEk1C
t/Szrjv3FqkTAHV+mjB6ivnMVHX3BEpngs9P8SlRTmVZPN8Fl8lSHuPhDdQjHz3I
yb6luXOfyxdpu8+LpcrFuUYBTZH5uGh+z//e/wzRVJ8HrI+XO9tdifWnpQ/3AMpY
L8jaQWicGyizsnNXC4XdOvAkkpvyTQ2+MEcLIdaP+a/ujpnFIQTdmUrrLZzbby/v
bm5zHTch/DYJNo41r+EF13Qzx6ZQj5E1zriFWY3PD7sRpinEejbVl9MShBNTESbP
vuOkO75U/ZWuKjnzIOOsXjNe0Elc78PQY7TozxEU1SManBugNYiea5UIjVtXQz0H
YZhfCjgsS1yYA/TIUTw4AGv9j8H27+MCbSsB5GmcgFvy3h5EmaPk333TeXZYxVF9
y4vVzF3nZ05kIeiuSpXY+56EmugeH6Z2TwBsx4xVE6glqO95SdKhstrrp82C4138
ThCeyReUA0M9QVDpy3qphR9BoB5Lkb1TgSZFsdtYb96J0J7oCzNfAPoaoEc5UDy0
OjQqiaV9co1U5fIQuB/ljjdcEen1mUNwNMVAUt+MRzZi+Zth3GlchwJDjWMYwS1H
orBZ8StHfBc84vlFZNXuQlXqnrIeWWJQf7WRA0KDMxNYomb5yYucT0s9SD53v26w
Vmmj41bb/eM7v8TcWaGG/P2kyVjoj19WWdKyqrJMNs+YQ9wfILK/QaGA+ESKiLG5
V7dx3psHtsi8c/VyJrQL6YNjgyTgMaAgUdrnOi5WAXuqEJP2pf0biffAEVjSG9Mj
dJWNRoa6hWyRFB3rpc+BAGtJjXACoWEq7wllgt39t9IeLtYceN0W2y19W9ZsRbK0
pxNeIECkB9g+qGqgEAQR0DNOoIW/WTlwub+A+Ug82nDfvqHAFaGdueHzh79t6X6W
kRXfQGNMIQng8V7e+Wk+3/YpAlJtt19iBs0KOgfNoxrKf/hL1qSxd0lSB18lxdz5
Gxa0I14S7m6iUUNY6cNcig5+4KTMw6DzMSipJROEt1p9SFes68fpOP5jNlGUHCh1
HDa8txZcVSjSSthRyXxm4LI5wJfaO3P2cxKLZILW4/q2/f2LH8lvzDBya+lqPiFD
zAiOeWutyxPhMsyxxoERILOIk8ftTnZkbHbLA0pdOHrlAtlsBPUhmhLDhQNxozVM
+XXVE8GPQNpdEFnlBP6sGHGN6uIdYEpkoTrvPjvQ6gK1oBECcfotBl137h4BrQHL
YsvzqtysDvMKVYS87yAl/WcwrpIQF4ZcxjKrt+kC49Vd5NHVaB/HYq2tzlf2Xz8M
zHTfpqk47V0UdG0zixs2tTwagvE+BpUUIohexhyW7O3K+TZQuwilp3MOEQEqjv+M
uMghqzxiCQ4qZe5R6uPi+9v8BvvZmK8BWmmN14/3PsQXcXwOc2uKu5b3FZCjzXQO
UiEbNbPEIlwPjYUrJb+UHy0IoVNoBWcBv0rlLSjtB++uSxccMOq6x6J9KB337Oqo
o87MAxeUoX0JUlAI/H1X5IroJrP6gRuCrXH9NdsjJnebCauNVuI84QfSU6H8MIK4
cGjCmJFLjbrzdwZ8bbUJeA9oOecwdIbgClALWoFeinAjQdpazJXeXdudwWUxQEQC
JxNkaEz0bsrYZqzrWYunkXIBsHwdZht42P6KOd4q4TxhFRPCgUL7+LFwTwtKj2pv
UMFl9T8NAkSW//2FN1+tw0OQmMIeMmsVnSX8tQOHLkstkfcurvrpxJor9W1CbftT
FW1drgCQ0fsqIr4PKrqA34RVvHzQ68FkkqamFYIw6k1phfU/4Y+PaK6rotvb/GSs
O8f+typ9EkKLrWJDiFAOJWx1WyYIjRUgj4hc8cjniymAhpJDMabukg/1UMKFLz1S
0870BeQunk7+7N+pogSyKurkfL+SDhVkwhwbYvW7hOdYjVhCZpWiIyArr70l7P++
nfuvVpcTZWVy8oZueEFfvoIraCUkEFafksRT5e807elJbepB+sJY1l+K9mxG2/fA
Fv8SwE+N+WxIOJ/zDMPouHCFOG/y2Q1EvvTSS7liEI5rV8Cr8j7IgdwbbWt+aVO4
wuYgVj956mOavCMBCwHRsjToWDPwmGOutRq4+FJqHue5jwHqIBqTUgoSv20IgdTY
QmEv4mhsS/jfcoR5FT8DebWdwh/0TPft+Yj3yUqK+bndInU4AoLURRMRqrQAz7mu
WaFslB1LFzdJYmSwqgbiHISS/QvFxSAnemmtzXb9EeEcIy7Sm2iMLnDh07uidGid
8QpE7PDUPrpEaNmxFAjZXd9b1ig88h1Ujw2eG4vajC72aolvcCNEDESQ9Bqy1rUF
RhRpaFV64N7TT/oXdJjsuJweobOTYCKVvICGYRqTsKzcKJNRa6/mN8t2iK943N/T
gL3XovUpxBI0s0gJeUG8rgyo71uETiYcV4orOj5wmVUCGPlXtghnB9KMfDBdL4o1
ZFNXcjkDiKVRUEOPkG94HMg8mGFwPkXL9BjkoVaWpJGsEcgV0ADYgrcHN3Ls934r
+RQSY9l+rtHXGAQQgGM6Ma82Sw4mwkBqOZEr5r/VisM1lxwVZpDj61X1odr0gcYM
x1+hqA25ETlxq+Nclj8zrf9s0Nla7aIclAd6/YXbF4xCkdblRaFznxJc2blKPgKB
jIfwTALjCqUTytPREG8YWQosyTSb8Ej+wv8lnqsNLf7WXrSACvF3IZ+YtG2Ptfok
jnrXnfaBwIV95OFKGE3KBkgnyA7TLmniGvYmo/TqB1PfQgv88fRRUkJM7fh5PEts
mPNlIHg5VcnGSVxZMlqFbKJo3nvWy/1iaxT05neR0z/ImNpK7tGxoQTIpASE4Lwt
Q164KAhlQ6p4ctPyLf0fjAie5PCKY/t45lQqRxXI1ZoT2ab/HczAj538Ajwi2cOH
UZn84QEZhisWO6rV79QBqst89fJK2ROqS0Ob3PnlSt+F1qpxGgYsfrXnrgGZA/HO
fwQIhfZnvX06iVZbRse0Ioekk+YuC98zDqLtPEz+Ugs/xZ+FxnSFXbH7Iy/UanmH
r6IG59RXjLtvojkBsPNF2UdhFrU6ZFRgj6PdEK8FljVO5WTuE6iaksIufZFeHa50
IgTzlmMY0taynvMC6PiZ+TT+BZnNhdhzIXDubnPXeSTW3j3mxZYOO5R2nZMI/Cez
cGEjsEWoqZYOg4rH8NVuWle8pZDGdiuqr9W88wuHD5d7FGBZW0/Sut3q9+J9/p0S
7U6nVHfZIKmWllmQrViwdK5gOjdTSOLa0W0yFP8dDS3PqapM7dHpCeRs5iw23yVy
PqRfv14M4bYENJ4PgiFSMMPMLLIsRVKVKPgDlDrIyDFoHfbIa0wJHq3GlvwR7qkb
KwQhb5OJCWIdxZDmZ7hZkzyiS0Tqi7hGHT/sRaezJFYwaYPtLHd36woFGPZ+zS5E
myCMhJMbNTO0BqIvK2wZJRPOxO2sdxOCWfhQ1giZqYLMc2tdiNLtHr+BKY6iBlr3
9E39X5B0Ot2lbW38+H7onHaIq3Qafd1Eggi6Qj0iKMPxnieD9870OXuqoiUkKtYb
PdW23FVbn7ykIhloRq4PgGzc124DjWyhgI+ouu45Nfazh2EDl++B6ZvciA4SSgS3
V40Duop/ArCJreKlaF64inkM1Ettpomesy/3wC7t1B9hmyqfDcYkkKflcV5d87JI
0LlradNREj3pGOtSFKvMr6yCTiBqXI/GmWfZp4YGTGdtOyJzYAB2jyXlRD9h9Bi6
9m7aNkYmQ6OvmQH/g24GkZUs7RWmID/rdMlpIPu7by8TTFLLiOjFD9MhLP5kD0/r
W71rEG+AZ4LGLR/dZf5Na90jUQPDhKekP90HLq1bELjcB6MYVETXDFYR+noJBvLi
YFQF0BTTJUTaiAA1+2nBxzFRWCqAqVFyNv73UXp8cnPCA6jQ51tOXXTXOmCOP+Fs
cLdmTbDMRHvTHJRyvBZwGMlnNS1dG3mG7v+5wk9b3YooOTjwHrmq09di4SKTA2T0
VuswKgfcrrnMvo2c9Qt20Mx6j8pKXUu4ca2COMTs9MjAuVFIdwamdSBEvNWAScy7
TRc7q/YBcVqBJl1RJVuo1GVu0r7iCK+Q0lZEM1VW7doZfzAFQLYOlM2zfkK69ntl
GOYI9ekB+5DH1LhQXw8nLLHDB/17/6xgLGFshX/tcFoUaG4pqYlhECTyUAhPNUgA
mIWnmKpsI2EASqIfk/hBu6QxeX7qHt/fuKnDyyg7HZJ372WIOhPRt80IHiaxwPDo
XxGb/ilwPQKJ5rsxzzYGqYwHsdFLRC2BHGXYFHlRk/OsHZHvBRTPV+DUBT+5zC5T
c7htFi8wUdVaBfdZYnhYvnWCYanUG5g+DaLbrS0AlU37r0MULjMb3ABl6ZsmLGT4
9eONEe6Om/wrgGvk5YEBt5pd01ZiskcxzlDoRQ1O9DRCdfUssHNcK6b+Q6ngKPfh
XVH5cfnNeDuJx3ryb6EvmWJhEZ6RuxefAi8SK1VPH0EVtP48cEujXaDG/zYwNB3J
VC6bTbrK/3t7u2SZp5ZaYTc7glhIjz52h7Etys8zpLa9Mext1Xg/wCqZREcr8WNf
YIbloH08R0mfYvrFApWeGmMplbC+qVEB6GLEW545tf22wfuTfYiKLR6keiS85+gx
C/nAnsazB2loVGyE1c6wiqJcQrTMjNwIMSZec+ov+UZWNTRxxFG6MkXnNeucA935
w+GBcNugw/jRySnD02OqJbJruLyVx5A0EcYNawrJ2iXcK068v94LE7uhzGw8ZqzT
dqH6b5EAYrIGThTN/Ehf5T8yESOkgTynWiBmXTC8EnH9FB+I0R1NlFAwKSBfsSjA
IBh6krlhbQxkylSvPP0C2M7W8frnQTsF12XFpoK4mNtJWtIoXKJFhUKkWtziP3jA
swin3O/19f7UUCNBB/+k0rJ9uVN6G39WN4jxpEHAy2ThuE2YEwmWaBI73h34v9rH
NeIK6MOHngNFAu5Pe7YadEdO25vUGM1e22jWRWLf5JeDa9M16/tESY5V0ATLfoIW
VXJCYFBfKzN+pR+IphkT2DJXt2ctPI3g3YEJNquzOT1UUe26x7mDlMJOAy41MbS4
oUmeEQvTfAgE4EsYV8R/1M6JQI0pi4BwMxoKKBimWzayx/R4MxbQrbaZE13E4qc6
mmzwQ8tHVoUiT4I306yB23Dp+hMJDquIG7DfmyFOV0Cokl1I4F0EsTHHqGUR0dNn
TYaQ0hzT1ZcdmD49nx7OkmAECUNL10ds3p6u+OhMMEhFEGJoF98th64prNjGtuGm
7OBFXH7VHNmd9bNDVLH3oSDgjbJYABb86jkP3ZiJvlzM+VKK2WfRbCjicBACWIvS
T+TXvecqTZEeyKXZjTMOtgv9P2NtH3HbU9efBO0k/n7Hi7bBZzKz+5j0WRsbbTGP
b1168OoRkO1omllRN0/tRwKG0szSiKDc8YsltwoblqLVNsxbTJeJ3CvdjwwdobLI
LGep30ealEhyLWc8yPq4rIxkuyijyvYRMGeEZjUOjdWcMca+/kjA3ZPBvPVioJF6
q/HY2zVLl1uvZd7sveq2LcYnTiqEpNZBRI9jdJNm8yamy5bs2WvRTcJEoSU8t/82
ZANMRhstLNJ2uHHDYBLqjplzaDuJ2eF6dr81J+eISlRqLTwVN4OSmm6wy/vo9HOp
SrROy4wKAIj2ri+GBVA2gsi8RFqamlQevjq6syBjrlW1CEmI5AFsXXo0ZW0UqYb/
wBIGvT4LoyKkhRrQa+HM0FfvvfMokzERXtkUgSFgO4Z4xezd2odclCjZ+gI0UnTQ
9ZLrZZCRwTeBj+K49TwCaCNx3p5x+xT3qHY6ajnTGUHC+fUlroUuECBuh0Z3dCUF
vLXR8eU9mnRQxIDr67HbGrEnY2Dn/HnWacYO+tC9Po8iH6bBVYCDxBtzMRHTdE79
n7czytyFYUByXilPeA8k7H6E/0m18j1Cx50x6dnf/8ejWcMyVR0CqlgNPjExYCfv
tjiNP2wucAqthGexcmhqjoTJIQmeHIQLSEssIycz993v0Z5XrYHdHDjbg4sIX3kp
r9Qwj0VjxISFdoAgXHlPZpftR5LzbLNC3wjiC/OE+85Quwg6S2C0RqvqviV0qU0D
vb8hs4/H/GInagUpZudjSrzOA7ilZ/0jlUNfvdl0gICwmCuY65+sKeu+Sg8QGrIt
0PBsG9ygnJzPiWCghtWV7JNDgtv8MIM++bXPuxQ8GAITPMMQoZrifjpvui7HI1i5
OKvPdam2PfVbbhvjJkrM/E6a1ZVkPcHS2gHhEXBbFnol48JHQfvbbDoB+YaCMJwf
LvkCZsflQ06PdkVqobUV/yyJdpYMopQgDKHcgVGOHb7pxSKNfL02evwoMSPsiYFU
xHODnIymc4XiPWdjAsIwQ9YeBLTo5ryh+38YlycEG97dl8R+ha+lAVRaBnAXh5j1
tt6sgk/p0LsNIWR2upGR8pCLFcFM/NfN9yUo97jcG4bUQhHWjv4IjldoPWQHpmQx
PuOFGqfLuVIOCZCcFD8mZxFAvbHtV31yqzxj+nREZ4RUdPtCXZEUZ83H4mdOCDa/
FoyF1aVFOWYEYMVmUNK3I06DRDaI0YHsKdlgiJJdFzFl+rmWxn8CB9Xzs2bBrmoZ
qnlupTc9BgxN8odqEhWKwhgDQuAejzJnP2uOorrclmuemB1FtcECY8WWjtjEG885
iJ4e7Gav+SM6bwdiF2cG4HJQJJnX14qwimNKKaQqKB5oNm40F9VZIjpc3cmgTQPg
p23H7FLeEFfUdBlRv0woaQN68qlkyMlZsUieqYUnfAQjDleB4pDMtzjZxSOKoAdJ
UXqESN7WIpWLR2QJWx6AI/MdW+J6HaOKc/g/B+QZ+6gO0zfBjbTVno92WIApoG1m
LZjhJTsmBPni9uBWt2N3WuSVI6fKL865r9yyx+ZBAUEhT1qdFqpqGktMk887KIdB
NI3ErQ4kk65ESnjjbEUDwiJ5OvCejJE2Irwo1shEEZY4T2Z44hFjwUQ3lQwHAzRr
0Gm2yteFvXPBe1o/A9tUbrcWdb6pXtX+7zgCAJR2IFmBaAubuybTmXUySh6k6k5H
hWNLSnEsKAaPM+yn9MX9FlNibsOcDQR9IEi1FJRav9nJW+z1i6et/cTc2jJ5W5X3
6+Ibw/vAUVWe+XbebgZCTS4T8oWdCBXBaWbajWu9R4g6G2eZRv8bR7P0ypLJiOK2
X7rs6agom0SnI0Dw5TQGhO0yK3r03VfzvWfzPoEA6BazbQVlw74gBKVY959ukYOa
kM4M1TH8QlN0hLi1+GQ/jHRj+ra8XGUnSsWPWEOdO5TOymKCYqTmmcxHCipwlY9A
opAYOh/lW7ImRIYW+9GqGaFm3d3hmI5Ad0VodCqOLYNki+cn5z3Mx3WFQX9CTL3v
jSeQvVdFxqIOXRQoPoMNUd+q2PY9+19qRbc+G9iftq846JfSoDtVL7ncvoFLBQr/
8A9x3YSny/U1cWUXnekF52YMXcr0veio5i7/I6L+Dwxpib1aAXusbwqg+CAWd2Um
k8XCMvOi1yDZ5YtnB8ARH80M9ADE5rg5gZHTEp8gxlyH0jpoXPP6BfY12nYQekyX
Y0CL8SlU2JJgKx2d5jhMS69lZcqMQZVOUx8J3tpHD56oYiK0W4dkHDqzsO7qF5K/
gb1gnzdh4dWyZANp6Qe0zUOiWbQ4geO2ud64uPfCClmQ/9INlZ5hmUMm4iN+lL+w
mVtsW6ydH3zHry+IfjcOuq7XvXFsmf92jS1K4SQuza/Xypqrqi/V7Ar/rqtwOJBz
5y9CNBlqX0i1ugXafLPvDQmEEQYK0PUGkviBOp99PFS4H38QV9VvvnWya435b9BY
VElMFRqenPxFI7Dc2jwN6u94JNXA5/LU5n7KKKsQifmrY7k5odUGCaRZ8Ga8sUJ4
NEG9apcmATZ1w0Dld1SKJNcBW17MSwTG4U9IxC72YrmcMYO4ElNptxpcQQm9c1Vq
CXBhMjcFOceipyXoVrJv8cHbpMq0ERuzLoXsU+OgAA2TG/TEBi2AwRhVhIwpSazR
A4cONakWCRXvIM6W7X0Y53+7jAK8QYmjbFJahs/TEIM/mno4jsl+mOR+o02NPb7K
/MgyU6dNdig9yHnb05ZfxfU7+O7hN2vlD0eWZJrYzfF9C53kMZlO6mOtSOvxSN+P
We4ZBBHV/gF559lK+CYEyXGKF0XEyb4F1XreGgyvpzI0m1htFKashwUB9oVfgg94
k9RrVrKfsVmrE89HPxiNU3CuefeTKuXOd2cGCtev7GAwJOYyRPJUlxQfvXfc4JNa
PhWYBzJBXeE/i2aAaYfOuCLRY4Tc+AOdybZHX2CkszbqBaLFEBXI++O4bLWxN1kW
BWNmThHkBwaIlPEbmjdEoUjdhE+5xKtMGwhKhhI9B+SB6MYJEs2aaxHWQyI4AoR0
lydaycn2+hqoMRwMndDYLQCPqxL2M8q1T5ymm1eqlv6fLmWHgpnpAUneDM1+ddbq
2DejAn6PestShD8mTLRpfIg2DDZvRZaibhrpj59S8SF0e5487NE6luuHEfJdGjHf
6ZHjpVxA+BQPLv3LgMeBQGtVhuYt3LAHijbt8GI+DDmxQH5wIA6kBTrTmYwgDqRg
NoiMYNMtEPO8BnIQaWuTwaCiVLmXSHFk3QM2eJg9vukF8MjcUWyOGNX+lvIExfvL
3PmeKm8EpiMtuXmFxLFEMbFu+TYVUFKoN5yBHoTR58VJ8JPnpGk6Lkeg2T0/hQ5I
HGS4IlBtvep7Vwj8w3dyRDQsHaXReVJgGmjQo3HWS0F9irHff0Xiaou9y//6EaCX
OZBNEaU6g/hC1qShHVoArI9yXpYFYlzAhUq4gIo/hhYulcqlhF5iYnUKieynjtqH
fl33AOXl3x62UKfSfhwLQq6MKmwGn+Rz5mC2+KrkdRlqXFQuE4IDWok449UKpi28
E2z2kFgOl1QtnWRFNoZp8eU0LsIsARhrHpN6P43dUggg9KMmx2F9iNR307zg/lgC
qAqf8HBbXGElLJuPy2MUIs8SnHNzYSABr2Jz23QJzF2XQWjuQ18fxYwyxEErTLOw
yOEJvPwuVd6W88pvSGeWAeQ7HtMMsEu+2sWeI0Zy9upkN4AV7sbtI3xHpRBA0hX/
zhYRhL9ufxk71cCQNYevRUymYkLQleePVPhfD/crPEP0udJGdJDeuN6kyOLC75kI
nM7qbdBh2ZcTW4S3CpMswncacXmPBoEAf8mn3t6hpZyMRsGP+678WHi59yO846ZS
RnCMkpRbNJk6fywSXC1DHYB8eSQP5eeo95KjRUC6VDBoJDtu2B5nLbXi9w28notA
EGaqmK3LgKmAuwn9LdpzRwVQQ+zExW795T2sJF0xW/h5sLwsECPmxMnvv2dMzu9E
HpZEpBu5jMDY4AoGhfrdEOO6Eoh44/VINdZY7L0Vbr/Eg+eyZZWcxDAfq4xfUjsa
/kYRdUA6nVuj2S5aRiGHc967H/CgLi6KFTMketXJ33WhrM9TJqDT+JfkMFDijxp4
+PPTi/o5gVwv1pJC7B64PWZVd5oiXeDfdjORC3/meJa1mAObY4HAJGaS7S0FfJnd
7egTfp2PzSxyFO7ZkOESTzD4Td7tzpuBMyoV11Ipv9A7OEK4tfzFikbGBAbbjQjn
3dgfe6czgy4+oJgMiFnefpVBtLrBwh/OtX/+SLUyjZQ+rFGASE8OKaTEFq/PWMWM
FLmyDaoKiQ30MHObQS1Suv4cvV0UF1goTUzFLFaFEyTW+3v3gjEqzKEOFnmKXFhG
7q5/wrLGzcbSYCCMiEKHXOU6tiJCnHxnhPS6AHk4ISQA+Xg1yT9d4Fe3AD10bUbE
rWnLXeU0sLpvRvY86ABE4OyN21kw/HdPQDRvLJYu2FMASt8zST9rxpe6wLYAxPUw
59LcRbmOXBtNSb6fxfvzsVqEke3XkpPtgvMsqec/grpWNrePMYEogJPoJs2EiOoF
DvjwD8JeeM+sTll3lwH/txyMwAI+xnp/4zKwQ88wM3FnEdj8bOFmzuKDV2OQIcGA
2RR0ReYJQD24XBgFw2kulHwxXKKFt4D00SQsJTD0RKSUWSXbsVhzIaxxGjwqmZ2/
cu1ojY3nvstR62SOv0YrsgMp0EUMMTo2lmFAdJTiugzhgicUA2EIIbyQhhhXYqqB
sxkVrw/tCk0i0t2ip2jk2huhlokfMXcgOwSpKWhymR1tZdY6pWy+XOvdx4U0apS8
z1gmn3OOA83YK6KWwMSKwHjnrT5tGE13SoBHcXyYP2FAMUltP+UyYaBaeaOyI4LR
hPfLQIwt259MbUgrp1ZaqaBXGRUoUuYqQyawGecEwm2ZfuAGWkJVmYV7W/BxVlks
CpM3IKilEpch8Tt8l3q5SIL3wlLN1EjdA/vwx6cf36XeUKY9CCmkXQI43h0agNqi
Bf5fNJIKU7Kt4gubyoQgKi/hqayhDl9BbiZEkUM8hAzYkueNRdQnoP3OMtP3ySfn
42yVJNlPdIk6nLkgqZ0u39U9ER8Fw8U4M2ps5j9K2Yp5dQZRUXrPvIpksB5YUi9l
iRU4U/h8ZkAcLVPG+kdSazHRq9A8wiBevK2JD9rEmWFPmXNKuk2Ux+kXpvSLTlA6
VA7h6uZZ3zqGJMj4nMLf6I+9JCeG+oGFdT4GNNYORvDbeVtmf5KhdcGF6VptFJGA
ahcUZKHd/bUH68876f5PAcCJNEzuIAkXrKg/yBRQTH3oiFDBPLoDu+MyBu/mDK5z
DS4Vw5J4CoD14nJ3bLknQEm5CtfOSHtJtGIv48Jl0Xp4YaTpo/rZm0jXoRy/N5FX
9edktp79JP6CG1YwhgUTnTVWgMDX0bXs0ptmIjc4ym+eCYo5xB/P1SnPyV7XDBts
d0WFH/3I8vTXG8qrApT2MbidGj9bTXE/cdE57yUTts6s3r6GuBIzzRMSm0YnhpHq
mbIy1x9HwznIox0j7McVdHtkj9KZ9RystAlfL2kFknxIaixgeTNff7y2fhZh2pVO
BUeLvDU+Wfk2NgpQT90i//C7WtUGdc4uGFi5pnzLsMAXeGH6mtwxDY+Y+mrIa1vD
30eeLHTamahWvrgXD3sTbElg7dXI7Hy0o7LT7ZeMi1euRPt+4oFLel/NODqBX2iJ
L1hyIfjWzgNQq/UAnk8YqprgsRitIq8deSagZRUOhP/rmRIJUt7tQBBHZ+/UN4j/
IhK6H3432zhRLP7uFIqha5LzdHp3Wcs8gvsuO7WvDcqvyTcbP9OGGUFSUrdAaTT2
Ke45GQTPc8ZcYUYHtnbNg4du5TVXriMZrwjy1BGBtfWtRClbDdRYyIPwYhzUO0xm
pwvJj83Qp4ih26BstCgu35nt5rj18tMAJEQF0hXam8P7/oGPiEArnBul09LELToi
qHDb8IQznl2Ltd6oOY0H3FpTpeBbYem9/Ftg3SmGVVIZCALeNo65uoqh7keRlmCQ
ISHefhZgdX5XJh9Fk/E8RR4Q+AMmQFpzVksP+pk6doa4tat8xJDYBNFfM1fidYp/
e+ev2tzxt1F4AM1pqUqcrZnsQeVy7soAgyMkgC08Fw/Z/apB9AbRDoL4aSAU4C3D
C1j7m9y5I+oZV68YHlK4y7/rOUVA2Kt5fk3giue60LrMnHkKhOskdPj90lDR4ZTj
NFsHVs2m2QMMA1VTNqShJxl09dT/gUOyoNalGGacI/qBaERvsErOLB7Euld9RGpQ
YaylwABtrI9Z+PsGuoWIgzvn3vL+YW40DL0t/N22j1xUWbeUZF8ldIzAdmI6ksj5
ftZwmI4MumpNA7SeSbNBmQSNdc1060dlaxc30uNTfWn/UpTnWPjoKD0j7umsxGJN
w7V86r32Po4cLN0mIAWmgu1G1Yo/G8CQBVdxH+/J25Xim90qTaQTDWgucUwgQ1RO
4N3VpgWF58XgzFwc0LNv04dEiinbD3TsSvLzSFGbUeeDmXkFNZSCE965/08Y04eu
fiN+/JMjfaNqSl0QBSjLaRU1yWXISj0ePB28iy3NyYWtfN88RZtMgCUDPkPVyzFf
+FpkIFkI5A1dqdtqc3M3DqyLdwLrZ1Myys6x7pu1wycOIdEuFmqEtEuiknEjHD5T
nfnPuP5CW9g5mcwOSeujcZu6R9tS2W3tw/ZwBr9UR2cPTevpIKFg9AZSSiX5DWJO
YJm8Ip/MitKIfsm3ckJhWVfTG343t/r7EQBfF2jwerOdzvAIc+x+hhrDJvVLBJdk
8FLo/2YfA/a6q6lFXzdW7rqdL8JYyw4kyf74lMhsI/I7zkqA5gNewzbkrydN81cm
7TU4NHr8KNlaEBmhOK2/yE8Q1EZQ7Apm35W+L2GKwODJl7uDWjCKL5pdnLPLq90o
zVPTIv5E2ZpS2xOJJxs+nCFIvp1Dq47da4KZgJabApqI/eRCQUtbSRXe6a1vTRFI
jc6ZDGVwRYQs+PhjjzfHJwwiAAraSICshXjOFDja3m284ZGXTUtkiUaz2j927kUv
j9OEtu2lHvgjY7Di6rATt+JFn/IboYscaBk7cVfM9fsuRs0kjemMSSGrxTx7Jvfh
uSe3j8RPSWSXh2kkrfpRHd+BnmwPIpFQiEX3DbhcsAwuIUs/n8jqEujffUpy2gym
xR6HhCspevOzuZQ5YjOxu5BTFrrmyT05fqy9CWh6gMxCdLNjcl84GkhOK8MaHcoD
zeOY5gpIL8M9TRgvHJyyifuEjA8SuSYsyZzOkOdgS2L2cG+XKGMuk8V0r96t1FZZ
stF0e9rnkf2V0Wy7bICkbfsSkkrtxqr6QM+6BTjRBK4OVgiMLM58T9OCNMrhS6bi
eJf223v1GdTqi7adopNju6Owz0BXAH5FobpHKIFy8wnI1k2A352f+CyS7NSMpX45
aUm8E3cMg/5+LfwLnkL9szCUynfJu2oibypUkDKR/lUoVnhoL2GqzQ62eGOj/6Ts
4WMr62tzDi5bXFXt7hepmq41kKGztIkQcKdOINOkNXQb7Ygd8Dx3SpQShvtNC3IS
DavZBux1TpUtuy6e14cBy4dI48MSxpoV92FdEMyeUCNTJC0PumfkjkP8pWVJirCX
Biqwjx0dIo03QWttkEB+yOd3OIoQ1e/se1k09c0+XnoM8yBa1vIv5XRhP9LkZZWb
PoNg3ZCH0dSXHXdCkiRnM8J6ZxWVxcYfGydPZZxkUwqtw2xTWWHDJ7T0rTpUio+a
7BkY3c7Z+BbHzbRYYnHioconGa6Xv17UWpMrNWZ6OiPUJ4poTdJgji8FM8sm1DOn
4nCJ1E28iyPLEB6ad1rOavmJKhXZVEWs/NBfM2XSDNarJSBeRjGQTaQvisul8FTF
ve58HrWWK710SQahiVExbLRy7riNh1YefsjUV8+h46jiCJXTZ+hZa8/uyjIEwh+a
fONgaRbViqrygw8g3frYMX51OV6qn6qLXEpOnLeYuDe1fuNxYES+8aMoD1RzbHB0
WnrD0tPk5+4GYQkCP7RtsH091krwbu9fyoOhBhW00THyxz/Z6tj8o6Xjnxi0CT/L
1aBQq6URnDSG4ClAwmQUf48isQr2B7I3zheAyJ2V5+PVJMeBAB+M4YXH1NKS5Zup
KYURNi4gAVRU5QdBSgnEuS0s0yH/LAYS7BnODRMNeu//zS3GMHL8C58rGNc8wV+D
vIAutSNFXKanUeq+cPTliRm1DKgu0Gp1T4w5GYi/6H1qyiNXV+qF2wzLe5Q1s6A1
U9pgvQ6GVJYAhquLOCCUlOkrHc85zzLE1iL+kU1s5eJZc67yu956sx3WfLVx3EHB
7Dg5ufH61oGfNyl8zbmalWLCX+2bDG6uBfO0J7LSAXfchF44a1VDIhuzZE8TbQhH
z0Q2Pixvb/e8afZMXW2wvWoKfKuy0pObRUV++IRh2esaYga8OaFse5axuU9+jEKa
Jebzx22ghORCkaZV/reCaJomnNzqO5EB4jsGh7rgznnWUdeo+mVPwDm4ZJz0LFOA
IQX68S5ZPe5iVSoRhQyb3la+An14nOaGemrZjFD9CgydZmBjcPAShGyAXWcwjsOO
2xQnmprKAzpsE8zwzpZCAKTXI8EyO+8VLYCVN/XQ4vCDJmTCJci8E/h7hGI5hv5R
dmIWc/z3yjUwVFMXNDD6LAR+35PgrmLnM5jySvn3KbBKH7b21DazlK7dOMYyEhCp
LF1uxPS4DjvkWHgHcv9+NXcv+GbrRwnVkFFOWA/zh3CppJTdxVkgGYtsRP4XgN9t
xPwqNfhCS6Y5ts9HrI13j+mnMEX4LE5jDaxCIsZyOPdyKUdFARrils9EyV6SsQFC
lSNV9FTRMPCKh0dYZbUZYzfXZ90poh6f+BGpf6uu1L7FNjbDUk9ALCeXhX7yr+jz
2HZ3ZBdkVSNfCI5kP8V4SeHuDbaqFBr/DRpdVWFIlad9p5x/FeU50Vno3TvbMxVe
q9EXvcwXiYguaeeUqKAzNgCngp8XChB0kAqniY2IokgG86HAaEXaDfkbPkDsiBE/
03yJOiqQkpyQ3Hj43bWPTBc5FnI2AgL9YhUZCB0ACVGfzM8DDychGIsPI7Ia/QAe
P7JMLAswhfcU1pZRYvRHKIJzhDTKX4qt6rdxWWvynB3hTzi7SWBURu3SX6KWNVua
bKLpvnCS6WG+E/2O9Rbx6yXNLn5qV0ddJTTNR/DJNxtBwED3dnCgMpSxU2hXPvge
AGyTDHZSqhd83xXZ0k9agv2XJYG5aMc2nLpBYePNsEZUH1vHZiyOKC9a+Zn+rbae
iipo0/WKIhHbZ1tGAWyQQXATkDvSsrpRY1RGJ956bscw/Jxm55J0iEUeePpFw54J
6ruwHpPWOIJRRqHpw99qrqupA/nk7FK17B6tkpGCiUUuzttjNz7XH6rIwdyixL+1
7Yh8T/GHukmPF2dstQFyubVwrx+nkj2FqblZhRMl0LMF+cTeBZ3lMVShoVevdasg
1B+PFDO2X0Yqn7L2O7EQbUo3kRuCxW9ZpxMWZ7Sm83yB1H54aDTlwvvcZsWn+61B
5XeroNg9RruVZX2Z39nE6GTPQKTDnqGxuhDiCkm1VX7qPdV6EdKqM+hsfPSvbVOJ
qMWgqgmX4ryxBrKf4jc1Qv/7YviRX+E86HzzRh+HGlmZG12i4EE8+KjDWHso1xhd
qkVF5JE8e1Yxxd3X1WFtsgqpk7dEr4NeAGK3kW3EB4zNQwRNuOXCJOgB3n8WGiTe
wGU6xiLMryCHrTAYhYbTs/IcuJWywx8moSBaDXtXqdvuOFmKMXHyfhBy2LNScx+A
fG3t0VFtubOznWixK+BjnK3RKPyiyZSaiDYOFw+ACR1e837ZXIj8J1OUOGzGDhDQ
+bTrWfXMj+9Ihh64jgEgVD+88uALvywaiEcO2e5U3uoDMTdvQdJ+t0eEFgWr2fyZ
b/yNBYBWQZFb7zQ38cAE1mPVsJby4iAjxBVNGh16LDvaBJ2ok5spEBuBjbbBv7Rq
ZtEJYEEYcWO/NHu08NI8r1LdYa5JnNI6oMJI27yyXHIXL4lggAwfPBpCRLRswPSg
pRRuoofbdf0bHBWrqTjuhjzgIae2iiExkpGMd+Phj+48LYNIY4afZdU8NYyoOISo
txIh0sSJjh/9/n6YZBHZeBY7g6N1A1akRcN8V4oRIVKufqa3sqF+kVXdrkFFsndm
zSSWrzMhmTtT/K/8MGd2PaWgspYlU+406Zy2gHTEgxyZl17Ow0P7EIlOsTKSbnwK
zL8b1xWNoCXo8NWVNnO2j5d+tB9ORnWCS/bsUZuoFd8j02WSEEwLqlAvvOV4g+iY
VzZ9Gvx4iPgDAZZ4AU8U99QAcNtuTTbXQQhac25NyHMgxMtWybUFB74KdUIyLl3y
Mo4EGtjEu62SaOZni92cP/dq4SXE0KoNaWgx+oVVfoaS7TWRC4X1RGuGNTIHKRcL
7Fv1v77CG+B8XCYbz4WavylehuSlKl6LjI3xt5S8Z5YnwjRUMx+Zoc5W00b39cJv
7HP/ZMnjS8AW4Yj8FtK45r0LuCMk7Xt84X1b2Q0he/hqPjYd7lzZpjPpV/d8uQ77
4b0EMAnosWPVfRQu+D0XLuuNXq978m7gG4gkGs+KTpGDp+WWTh2qFVyaam+j9/qf
hK1JlO7SlrrjHV9ozLxqG34prT2XBfvSe5jcwaXjByEv1K+TZE6csnPreepJjXqL
YYA1KWTa6wXkKhZknd2OU+Fr7gdxw/kCiic4sMvPrIB91mvbFTtws+Ygh8fV39eH
2FABwsoMov36pdxcIJB6g0Ix0cfiDcocAYNtoWmK6HfFHOoAn6+fTitAJ/PJp/yd
/Xss5sVbGmU09V5hqlsAksx1R9o/Jyoq+eDdBjiQjnPe0YHRS9n7zhcND1ptxeFt
ceGFBK2cylyFPpVGmrlkUzXUmsxwIBVnIRPO7h3WJVZ5O2BMQL82sNiFCBbfODOs
WsieL+LCtzrMpEU27CErlCgFIVfJSYGaunNFJEBEAhWXl5hjRWvsanAeKDJ1kG21
A0TI/kTMOnF+Mly7NGUrxHWK/K8TVkkzqd93oxfVxsQH8WvrO1RLAlj6rjxjZdhw
xW8u8YlVkzOACx/fGN1z73DXZOrDTMoFCsURcfMhzV+LYzSd/QwvyyMQDtKxiF4c
+0N1kL4rP3WbatuwcalYH4JfH53m8uUPwtxg84CMC/h0tBevwwbvSEg3BNabDhZX
Wh4eK6QLmI4ht6mAhD4nZPWdr266y5Dty19807uSnayG44I8vbG5Fipfg0GktbTc
DfgyLaWVpa5SrGASdQFb/zWhT71ScF+EebcpiYIDx1ce6WjrJWtShG60924vxp6w
V6n3Pt9FZM071mF0vgBMOrvRkRLivWoIHJy6a3Whzm6QSwZbBRCZiQ/uq25RFOFn
CNX5W1l/GX02YPyjeZcM46ho74sDE3zua41LD4vgm4T/tmSssYsr7nCoHjJin0Os
p3WI5mF69qHe2v4bf9hMPI+CCT3plu6QsZl+S5O2D7mxNEQB3NePT0PX5n0TVE6T
WsLT97r0V/P2FjTWcG9PGR/xy847OxOEUx4aZyK3465cJmuuwHR6OTmkAYnuCi/+
idY5XhLGyUcJ8UPLXHnqxwhJV8iEynZdWqUoNzJJu/mg8Is+BpFovsLEt6ElknZ8
BIJ7HL1EihKfX5kneDhVKTOGBevogH6cciKVKWkl7TGUPnS7r6sdbizSM4YHpaU0
0fYV/ixzQZGge6mPruZ0yiRuZPKP0Lve97cKgYDQBBBISPPq+neGXosbTbxrdFIU
VLMq55dXcLYqBAOTnC/dhjaYmngI36UJrGqnqOglMaJ4F4FKtIfQt/uDrFbiIYJi
0ISuoy/Hges39wUS9VvH0bQueEWdsW86YJW4/P6OUW3y9qp1qaImGrOEjTs2j5it
DIqEWlIg9GbvIjpXVy86H3CQhFOuCdqJn0HGvKzVqO28p3NWsDKEgD2A61fcT8Ro
8REO9wHvac6z8Cm8y37RqzEsejCcfrCT5lewoYDq9XEAmch9UYxGZOYtSBcsgFtd
zsQbFHdKz98qIizMIFD1ckurdi4oeHWCdZxBwm+hwJMV5gq+CHgByy+WTqHeinr1
UOzkPrSnRmR5O124S4LV02VikA6lrxFwzRYV2BWhmWhGfwUCiGVPEiXfTLI02X7g
uJf8Z+uwIrjODKQTDmKkgORyuuXw6zv4HH9JdHBSRzO1NAIX1H7UqEzSmdjVakwT
v98qE5theMm/Qfg+ht6UyPDJKsJE0GxumDNwDVT0p76gDU2CTgoS5kaahMgMQz8V
mn+stZKTc0pMsTaL7FkjjlThYYVL8rHbYH9hvnvtTOJxg4rX7SC5tRdZEH181Gkz
HngY1OSClm1kn9boV/TR2wmHG29HZOm7VHly0lH6JD3Dms1L/9p3rFs3cfeLwjHp
cVqBkse6yav9d1QQGtbMyL9W+95rnU84GodB9PyZB3xgAL/ST35kf6sfeCIp+mIc
iLJxnZvhfXQfbBT1sCM2FK1Ip15KIVqzJoM1LzOh2f9BgVcoRvreBIfaNeJ8d3fx
NsBPl4mokwxoHQ4UzK5ZbTXSG6OBkGl/ZQWCjVakj5f+v3E5xGvLJUluTFmRFwSc
gqYeWunTw2qV2oUlLeaiB2qM5xii+MpLGiABS6mbkLnixBBY5CkrRHhn19ORcQbt
ktKXXKXGguxwoNymNTqTHN0sPPq071vfQ0cb2qT6ze7oyZvnAoPvP2ua5E75+YFx
rYlTLKYOTzJ6lYjXmGlU2lQu0wsjWd7tTk6ViI4t/bJmLE/t+QyHmwvaqywtenyE
twws6mXFGhSur2vMIlflMrmueonY6Tdg73Gswmu3vKRnfPFXtxqXUe2kGZd9Orah
LxyqZI1dJXlOCYhMxZdG29PiyFGch7q3C6buPuq6uLLU/phySxXtlmcCg8IUY/Io
/cTA3XQLGQZD4V3j8CXMYN3xwPgI/FStVTrNo8vEvEG3Gy2wZ2x/o4QDziAxbhaQ
A6Lx4To2+TwcCROa2psBlbP5uTkgsTqUcikI7gCga+WZCpwruvxaYNcLH/+KS9J+
gTvVnttgHAqAa2PaYC9tyrYK7ph3ULj82/0F6t9o+Ly7axmRReNaIjCwFxND01lW
fCUTONQGAopytY8IgbII9qF7rFBQkt8t5c66AwT0Ckq2qArsfP0J58Kyrg3xIXOt
cFg851SnqZTbuXPaWJENo2peGkLj3ZhBT9muIx3+LLOHYTU0cMWslz/GxFbIb2ha
cDD8nslJw1rLH9jYly/OqMzq1D2nMcN3V4ct3MGuguCmL3cDttQBzt2MGGjW7Ufn
aIM/s11xyaFKmeQSvoCu6pPjc/YfIdFeMEwcREKoWiPrgklgwhdlCAAXJgstRrI0
YC3s44IfMB0dVsb+bEGFzOKLnYvH7bjub1+RizMkYgW3gok1Ptv0tMECu1vceYiF
Rf4pczymG4oEdQD4OP1df9DBBEonOyiU1sFBKVQhOEQm0owaBaV1BPFqER8OjZDy
1+InG2B4oHTjJ/xSBHTznwr1nMdelwOnzF9PwZy4q6AqwXxK6XUz1K5XBA02EqYZ
E32PWfr8gL2teWhaOq912QL2/25fg5Uyp6SpLOCdIXcipD1CBQab/rWbAIWUcogE
c7y7QbKBNyl8H4GbFX+NkTQ23frDgNHlF8VQMeNCoxeivQJPYIk3OWZ8OMvKwxt6
V/Ox0H1PDW8Ze7oOiB6tYmieEetI0f/Yjxnj5d/K5Zdr5fewAxll7heBPEm6hynN
sL+X0V+WxZR4kHL329fxrGEvHVl8vZKJ3S304I4OddxV4B8qtO1tHliCeUg/XGkJ
Rhtba1Ql7uVjie8BX3mLBoBB/193FhWL8XLcUnLNqbGjzuIuEyqISUjAsC55c/Ez
AjwOiaX/Murv3SGtCAp6kQMZEJnTQos9GwaaHmpLG/90q0rUVzMHhdovzornWnUF
uvsGPN75/SG/qpqJPudrjmZUxTddxVb7/OG4dqr1vgycP4XCI7jmCyxAan4/fULf
AFRzlmOLAVSOYdFT4lANFdfNkgMZm7MvwIMhX5eMXs0bLukMU25/4TUC+NE4hzJH
XSoOq/zidpJOP63yfS59kEa+qEMqAwPgRyiXPMRsb74BaFjhHVb9pSX2KUjJFiC7
Tlai5dhLRw6xBV1o7MHfG7NiIwtxe+X4rteUmGK/+qe+ZNdX9Hqluf4ifl+dhdD3
3fJTcGbqXeE2jh9EOZ+uTceRh4PXO58DSJ0uzSpUdGTJbkYMZiv6lOn7Pxsk3leJ
pBoEiMr4BDhYDAUGtmbv1cdMLpkoWvGaZ8GXDqH47PCc7e3D7Dm+LalTPOWgWbHF
dJmdFXR04tFpD/133xZj5GxqJAX1sJGu2hYVA0iL8C0ylL48tBEdKOk/mMoNk5vR
w69JwAGgn4xhugT+LUBvttD1iafOlECR60BJ/w1nMNy3bdVo1wG7ZpX7W+A8TPC/
9jAGaQkMhGYU46dZ9Q+YGSOW5V53k/5L3Bt6cF9wHNQovCWO88mApC9EPeVUp+K9
UIYu/tqQ9MwwsWxSlzJ6GeWlf75AQuM4tz0DH5+ScBGUP9m04C3AvZS89bHAqhtQ
9mrHtduOgGFBxYuViBUe0bkuV9MRFsXG5Ys05aJLruHBfv2ANTOnevcXAicWXZ4C
QJl5n4JpfMANTeFsqOFSyT7jmR4OTI8UOoWcLrTzuyV6V/CdSkgTGhVB5bSoB6BW
DwuE3xpCnXbcs1YAviXu7TwXiXNbV6GhT9mWKssaOK8rOKhItp4w1fAj2JQpFBiO
eOMxI+/aPMJ2BaT0rkQF/Qj+SpeSRIAhOFmxLcqrX9foSnpNOMst0QdBSdrHW5g8
jImy2GrNtwECTY8TnfZohrbK5mgPa1gOff/n2UVd4cucro43MZcm04ae4le4EqG9
vKeiFV4fbm+Ix7hiDimtjEumt/67PswlXzzdqqf54zP4dlXT0kTs0kWihcCqwCuc
ywemW/gpPIXT4KJXs3cfRABwmXF5DSNCDQXn2K0BWW7RYvvlUYH+evglfeku+qqR
NqCVbDv9HFXWhAR4KUZQfOvCUo8l/eLZ4xv1TrCpmYIfptqe1aZ4HC8SBwYulJNe
OTPfrg1X+xeP0Zp+7DYmLdC0oZnIeoPOJOYYSENjOc1zPzn9nR9fNs/xp5EHAwDZ
BBUdMR41sCarG1Upk4CTAW8RNnzy0iah5Xs2tv5274uTpZjpOkmQxa05twSIpXt2
ZRhRAcPGSfQVpc13EcWruVY5eMC7Vwm5xsC3zIS24xJBG7uwkbspmXN1h6E7tHsR
gpZlIMDw0OeHSwzxl/6/NQ71FHBkkpOyfBjcMYquit1bEReHVWgABrj5M08D73E+
Qq9wrGQ11MfMReDuwEngDl0P3Q36GM/Q/ZxQyu9imqmhQHOEdkR0OliNE4YEHjM+
CAXRHDtPF2U0O99JamV5ETFImpQAu811fMdv125Nos7Zbj0WuXyFclL9opUX4AS8
Wmt+GDSnq6/JqpZ77Z3qI/h7CX71+tUTOy8MJolFA0NLvYMn+6vncD07/cfNZbZG
2pMTlb3YzeYAaYFnXgN9TQgVtjmbtXz7wNyh0uJ2eVX0rYLxbfTbTiDsonFA75SN
AAZb+IzGExaMb0DFbzCt2WwiO110QLP0kptGD+nILNyNh0KJavJGU+nNzrytmfzJ
ijikh3aQjmkWt2f2wfnaZ0QtKhvlRVJli0FY4JDa07T9QeP0gXpL/stTPDTQaVbA
bXcoQkP0kqWMrf2R7CSlngGKthjnECngFYwiah9u88mMh34cxCxLdr9e2HMOwq9L
ISzCrI2IKHz6KHRm8NpZxLFahUJMHZMFhMf4l65Z7NngSfpXYNQjH8fqSVI981Q4
oTiBRuACh2O93FyQwrsFqVCLidLrkdeJAoiXyofGXhK622lFEjOd29NRNTCmpSby
nO3Z3wHV0huvWfZLEQrvHBP9rAJwQrei2qsN+g65JMNjPV1Cq6Hq0myozyrDGGqG
KnCrmeF5fLgbr3Y55Lhq/XDtu6C6B0X63+cwEonlQOLpAY/5kdbtn4EBlhPOxHPP
Fid1vYYHcihHuy7sAXWEa/S4HVaarjU78aDiQjDY+0cN/iSGbbOodJyKpkNT2ux/
ngUTlkIlKhtLYCgI8uzRg8HH8/frYd6NsncoBXZZOKUCw4iJFY229XdLDxnFYwDF
RvwhlYTFV+VYeiQFt0sci1qPqgaPtoxYpBJisE7btTAQFuTOmA532/wVLcGDhuHJ
ND1hEZm45ZGRLzPVqUETKKznmuDxsyHCTgE24vFNFImJpY58TCnxMm1h3oBqKKyE
VE0pZFgIo3iM9KdWR8lldK5Il5ihfpeLs1avK9bU/rdzsSrpgkKXIndYfRYAmyCP
1pmwD3mCt7VPfpdeSYrzMVaY+EOMUBeUwMT2HiOVcbhAU5W9co2IqSkwzLUK/uUf
VQMyqHzg7LJuccYWxy5rAekLLLdTs4DOTo220Sz1IPjYJUryq3ya7zd7QAdgmwhg
QEuQv79ndAjzE+H7uD61fW5gZXS3mmN4r0IF5UkFvLZXcWdcEYwW/PxQq+0H5N1d
CN3yyYu66oG30xs5NTP/JXxeyn0Qk3fUrST0tv/ivyunnLfz9q4JK2d/E9vQLtBH
DpCKrClgtphm5NpxMLuduvWYGBvxOVOA8HlvDBqCODAujw2RAiN2IqLcGUKUKQPp
pxvS/F7rJUnN742++HHlpJvasL1cyBhDP+x0h9Kw8qaq9INCuvcq0zU3uvpsR86S
jZLvXmYz6lUQFN8nDvqDOtA9yfmP6+8c1BBbDoLew0WlBEwMALn95DGmEDlqD5Lx
4JUc22oHzkJwuwX+ZhW9oqYbMVyT0cvqdmyUS2LIwFRiRNnyOZBF/xHoOe2x7Zab
Rtqd3r6QVuvzgt6uyeC0jN2KZTDvnSg//RYij2CxcKeSLrkkBnlG7xRY7CgbpT9L
lOx+xhG70SYfQRTwhB7CfbM99YI8GwPbMQ9NaQb8eW/0ngvCaS7lPRqas10+WgXL
YZxmMOAIsKTnI7vEJOsvjZigCkM95dRWFv2iRF9BN9fA9C0rUwybaXIJNkxP6prR
C8023MSVE7A0bnIJC4FG0Ipr9HkEj7XjeAReOHD5bbXPZzZ8BZBb4p4SXzk4puyD
W/qb1rK//knHwU9bxrTFfZzNhBpaDya8gcGjGMY4S2QpiBO7jWlQJfjS+3IUVo58
i7+9e1FSl9ZOiqgZ0pQyphdyu3PjfsRNxZaw7jQRNNuUBo2y+jnEQLvbJwoESPFt
pOr3d2KCcmHznMaoReGm1hMefnBsgcvllgJppHUQho9gcsXkmRafG9tSBopT7FLL
pt0vHCxQyflZEUEunR1lvj64ls3Db/LQ5jbnc7MHdCAzuonTSvZyQHRQZJE6ipec
0qkU14yyewO6Oqj++r9UF/rDJBf0oCp4iMOvPITo8vOHbvwRnv2TB72vbkaIM9At
j2K4/v80pC/mjF9+gJxcwyARJoH5CIg6RI/IU2eCwBPKi581ASepMfrIpH2UZV1p
FOiTCWOq4JTY4Ndjp/T434lW5jGAIOC/Mp+GQsll50HGeZzPCoSbl1rcN7PFSkqJ
g1ws8icC8O7rY5wChE/n9oKRMF726e/BYz9H0UjLtsi9dSkojCThMYdaNktjikWY
/v+y+X5BQXYTgQ1RZS9oyUsXUG0wR4Xpq8YekJGsck34gWmvidzVgRCCAhJbQqKC
xfZDpg4U2eicAiGc/6fFJs3sYOU8/XrP2zx2AgjODI+v7KjFyvV+lmE0m4tWgoGl
8PLokB9nol3JKnLlp+0+ZLgUJDpGoQL0SMLhpt71sOUCVvEK3SmTQYrre6DwJwU+
204hYSWc07abkCJ7EcsabC/D0lzFo84M+GRyLuuP7BAypS/C6dGmvqMweN7GAws/
czbUu+hGxZoGzAYH5lUxmZ20sqHnIJkg1pNXpIfKUHOXUiS2XWpNLr5jHhsy9gQo
PMLXFZ+w82+xvnnbwsO3oOgCw/xWrKq3U2fdWQf7XL6HwrxUxqX5jbC4tLZSyuYc
W1Ux8GdpDUZUDYO/muk0gg4c7P/IYRUAHEw3nX4kijaWx1+hTIw9CUKD8QkmIj1o
yay6QI1lL40c/4/FMl4WV0mntl0G5NeURBah+kYIDCDjxpp6VF1EYrP1sPJ0n60B
xhfXnfg2k6oES5Jc3dDyktcWGi4ym99/KShLIok0ru91P3Jg0KvD9meA+H1nrGl8
ZFh7LZQXYWWeOrN+7ELxRRgDU2A0Eui6BxQ+S22dPFM6u6FwK+qwyTKVJkUVcpyc
om29qVX1r1d/bXKtI+1Ie9uiuQ5fghTvcpGtO78e3pw04CkhCLHpyMYcXi61YWjb
ZY5SpWYFWyerJDcdBBoqmcD8A/nAh4d04472Cq1LL8Z67IKWUhmAds2UJNRQWddj
oWI3661h0MWM4gl6uHFukpH3RmPuUZXV0sLBGCelYHFyYAs4tW9jTy8PTI8DaGGH
PhRA1G5di26bi0gA06+1YWho+0xuKBRMVckp/dB8nCgQmZX62iMpjUvlWeUlinJp
8Sst6qA/ikwv5i0fkqfNioppoFbjcXUEs4agEShjqVN+p05ZUPTkNB615jiRMOFr
Z+/7Iz7NaqQ+mETmGZ19Y1/bVprTW54Lie0IuEsidaegZhuiIBLVtr1OxyX8FMBf
4fjdeCntqxmM060W1so5oBmwVeDipUSros2FxjphMEWr/LP7onxlgzj3a9LK14B8
DjB8GUm3P3T+RqUl7F/SvfnsaszST3nfzoAXkYKRJZe1j2EjO15wNIU76c4paT2O
uDGAKDCnH1JpE/wg6dAttzdtpwN9a490iPVDtdO/5YouAiMLvyHSdl9cShUjojJW
JRT79BbQ9RtUsvp6gc65WKgGQsk76KH2FdFSKNzL2xnTvwaClc5ZVNaGW7amLCfn
IqFwmLHeIcR4WI1ezS5j7+vQf/z0cfhsNEf+V9O/qt3h0mjXn4tgUCU8GhQW5EkV
BNanEHVoeQocKKTgO6buPC9zNC5eAjs75G2yFOF9kmHV5aA+dY8gCku+AmmMpsDZ
GQNbQwWpPWW33n04N4Vqd51I/LlHHLOOHIen/2no8EhZzy6t1axHa38Y5M1+/tEg
9GjLL7dVDivck/DdZxlRuIxwzUKrefU4qP7Cr0Qw7gs8EdGwWXpmUYdI5PnnIN3s
LTF+zuHCUQyab9hcKdsPUuXlSSZHOeV7rsdvVM5hBeO/X6dlvZKbGFe7rhLMQy0T
J1N1gEfTt/QwRC9bT4cgjLHWjWFm6kxfL3wSGVon8r/TwOs6Tn+6cPFUZvN0klF7
FjSoeibOVJ3n2+qlRKah7biL6hI33VMKGHSEusVvBY3KGjSVxqiKr9K/7CftBTBb
W1VSuU5qpvZkrnbIK/Fw3GwPTVVR5vsqXrnefT3nPqFUQthnWfDVJ3JpfIccPVPZ
WeZVV/swb6OQvsU3UttmOc8YNmVn9c/2IRg0TUn2Pr6JSq4OW2Iksd/P56OvWbLH
NUGtul4lD+XnA19D93fwLo3y/iSccRrZwBz/IjN7lVNu36h2ykvQ1PDpj4kougLN
cdLruw2hQolwX4PUC38Gk6pJfvHzrciZBpRVRXWJrAVBe7Vtg4wGcvPH4lM1fwr6
scTNd2Xh1/iLYeypyULuVWGQIawBwVF/l96FmHKomJCp0cbuyJYqNDZJrUYXtDzu
vLpD/SROBwYFNxHh0eMrj2Fn0fXJYxqpT2StqpkTthjqSz9LqaoFlQsxPopr+2M6
N/pjtiDKzPhU1VjVo9gsOZvHybZI+SvBbt2hKXKGucXdPgknLQLzZ2O55KyGuN/A
DmeTKAoqpGoSQbLSHqHAbItklXKZkZi2dErVph635uHjE9pdi0PC0hDR89vyUs2i
dZsuOhJoej97MiAZ+COkHYT6Fa5ieXuBt3FIQtoLoxjrtxvnixdIOkOrTarxjGN9
DiZAiKBFd+RpgSnLvi6MSKJTrcrTtbBE8vKxdxJJq003QhFK/uWpdhACZdaEviM3
C9U8qdkpcmsXfTapIfa2X64BeorrSMIdMhMGken9WDfydfmn0Pd7ss/Kvg3892hE
/OuAJyKGk1JmiNH83qflXkiab/RNV2TVB6g6Z+a/3SfhPOHRAPte6/bzwibLdcqd
4IN2eymMsGuEPv6Gxhzlo0SKg4ZL+hj6N+a7+r0BdQHWZS9tYmaHHKT1l/GNYzzr
fWIVtjO+neDXPo3KBQI4WlN3QHp+AVZd40tew5+BCWY/5ObGYT8fC40a0g75ybFk
jE33V1XvS6/CJongIjJcJzsYG8Ks+MjgE6tOOPW5mAobjGVzIF20RYKC/eWYh4ZC
3+WZk02xFI5PbdNLb7Gft8qCMO7rEoekbYLxhH+0EkwAig4SLjvprdscXzeCh1s8
aLVcHhVivBmBEM2lHsDtD7pZRyx7xONFAYFSIkMiTP0twVvbaRTxBwtjD3SXfiYw
g2KOUHXsoMl/Sthmp4bYkJWoM6oF24K0iVSKmObKMtY+t45cGcVXoFoEUZrvELux
ibo1/5rpyar+lxt5xXS/GRAgKdwYSTM5tjETb5Cu2oOj2C7bvwHBTh+9eyJaoYMA
ojncPk8NoS1EruiX9L3yARySYx11ZunqRKoI7/H13Mt2i7tunjXud3Bkj4tSCIfC
Qmr2EBPjpfDXsv7Eqrxl7oKjFGYv2zKP5p0WpvT8Jyta1L1SIC6nCT/YAltRHKUk
9X4BhnPDtnZxmWWxDPfwPPbWmhikOyFggS+/7GFCGdGX+/4xvQzUWXJbOmtrOjYD
y+1+SV+UwtL4w4dsaZWdvTrSXqh2UahpOuSCOG9z93MjmoamGQRKzekAl+Aa0gUh
ta538uErVAmCbD0aZkTRnpXYWUVzzIHXGaZn8F+AR5WyA3hcuiFdUupn/ku5W2DY
36XABw4VgfVsvfjZwbFtsk8d+j4EdycIBn8wA5bXcsG4bq3LUE6tRHqm76NbCvxw
b05fSeu5RXzDd7O7tluQP6sk6+FddZcNMEKBZV3IZDxpWs3CzXdJnnXpsgosZTrL
9FfKVDx4vrBl8c60ZrVJtu3DhztGgxvOqq9F25Wp+bhnVJnskTfQ91o/EB1W7Kx2
zAwUcPp+P5z2QrxfzOJzt5qfYw5p0VoLB5ZTK+dR4JSyQ+HlqGTL6B9LM4evHpgx
/ybE2IqSnnOV7i1BQV9R4+SCKUwQPa7gexUq8bjBS6siJgnQ6pmGYW4mmX9PUSA+
f2vfjHKqGUJwJqZeUJZNI673fZaV5q7YYi1h+0sJw8+mbGjDYyUKxir4exHqr7+b
3G2g8HgEitYkzJ8eBf36PJFpza/N/Q+MSCAxqzlDAKG5u8uKVza3WvnjgLzpEGA/
FQK/yKMc1eMKANgD5VaZu/K9mIaF/txZhGo4rPCzHfUc3D02R2X7cX4yatzhAYgQ
F5Zoq+yyS8mtjHZ6fmsXUcBT5kuMYvkSb1JGHcfxs3Ag5btlo0HcGppuwU4SNq5T
N4l97dohGVlVmBU1CntrYfsGjpCEobCp9wfYOsNC5Irx6+qtHOtCAnjAkZaP94Ig
Qrpc6LA45xJMf3Vua9HJU6BdDEOb8rxaJrzrTDEe4GuGpAd/Dhr57PpSXEBno5bb
cn3iCtFX/3ABNWWWvWH4Iyi8W6n4Z/43aj+ytxZAUw+5XdnASn6TCh0n7Z10h7n7
b8pOCTsA40wL0stV58LCJzRCpeIlvwLxPrEm/Z4dNQ0mI4Nnfq0Y5UgJ52Jkwjm4
/SJ2+5kx86E7EjY2X9tvJmWBsTQXv7737t9YYSfATNOAQErxFJrjxnpcBuyzgerN
HGfLL1tjZlRZFwkXM/aVhZWjHM4zOdfYTScAw+hTGGQIC/uzZYqOe088DpDSgf3V
dA6ztb7AHoUCWVAKwijJBz16NbRU5KYpP89gXAkkKPthxrS4hbnAfYYNPNVncSq2
JMZwvzSSDv98k7GsCbIqYd8B/zOYFEJ/384vuRg3FQJPD1QdHH24UZR3rZt2SylV
KOFwCASmmkyJ6uQtev809RscJw6ifD96rj+eOYJ7ftn++2gdrh4PkId1KSwyKOIk
B6cwE8soZIABx4R5wvPlb3d4Got1juLgCqKvMEJu69VyZ8lLxqsAqYsBOjUTUfs+
irWQZ87zRmVKvaeRm2QEvR+oLnJUPcDrDUbp5snMSmmElLL5AoCqytl4X0fkEOpd
SLKB7JYZaz6MQ2KbyckoHPCK8QhU9Jj78IjcW2W6JIga0SsXKwc3/iWGsHShceth
Oi0sLg3rnSe3DmjdnpT8BL6eBJ8JxAv3AgAcvUH2VfkAFJBH9sthwj0m7PrxfDpH
6LVBtkAT3t+O7tAZLjCdn7cbkrcOjQdOzBjKGaV7o8V22A5L5/OAN0QVHhGdHQtU
qd6qRE+Sb05CEJmD4SUFACxZdWTnLsYyTIJblr7y/hAYoIRD/YiA1WG02o5kdBlg
jkjt+9IdZlxNrjtIBls6oFAsWypdkrUYwyL7tCGqA+9tSQk4GIL/NWI/+n5cVqpx
aa0HAvYUay+NAevXdrKZg2+mbbGKfcNG2qG4ZKKZ5WBMAqJut04fHnOl6nd+jmim
QI2zDGy//2KdM77UtOO/4BuHm38Lo6TtR2yrG/ul2nnUQL/hnWfGG1oeKTB4SD+Q
2Yg5k/Y3lN8dRpJSGD4+y5m6HBLwgRMiF3ZDoY0sAOu/qtkOI6Sah2xUcEniPt9V
mMhw1A16ZIhj4lAvvJVesl9WGTQYbazlRn1kL3vuWrrOsfPlzJhsxhG/b7csiopZ
Hr/rpFBp51z+9bMfRXYGQ4d0QDmo3sJhyTGAiVJMGIg=
`pragma protect end_protected
