-- alt_sv_issp_gbtBank2.vhd

-- Generated using ACDS version 16.0 211

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity alt_sv_issp_gbtBank2 is
	port (
		probe      : in  std_logic_vector(19 downto 0) := (others => '0'); --     probes.probe
		source_clk : in  std_logic                     := '0';             -- source_clk.clk
		source     : out std_logic_vector(8 downto 0);                     --    sources.source
		source_ena : in  std_logic                     := '0'              --           .source_ena
	);
end entity alt_sv_issp_gbtBank2;

architecture rtl of alt_sv_issp_gbtBank2 is
	component altsource_probe_top is
		generic (
			sld_auto_instance_index : string  := "YES";
			sld_instance_index      : integer := 0;
			instance_id             : string  := "NONE";
			probe_width             : integer := 1;
			source_width            : integer := 1;
			source_initial_value    : string  := "0";
			enable_metastability    : string  := "NO"
		);
		port (
			source     : out std_logic_vector(8 downto 0);                     -- source
			source_ena : in  std_logic                     := 'X';             -- source_ena
			source_clk : in  std_logic                     := 'X';             -- clk
			probe      : in  std_logic_vector(19 downto 0) := (others => 'X')  -- probe
		);
	end component altsource_probe_top;

begin

	in_system_sources_probes_0 : component altsource_probe_top
		generic map (
			sld_auto_instance_index => "YES",
			sld_instance_index      => 0,
			instance_id             => "NONE",
			probe_width             => 20,
			source_width            => 9,
			source_initial_value    => "0",
			enable_metastability    => "YES"
		)
		port map (
			source     => source,     --    sources.source
			source_ena => source_ena, --           .source_ena
			source_clk => source_clk, -- source_clk.clk
			probe      => probe       --     probes.probe
		);

end architecture rtl; -- of alt_sv_issp_gbtBank2
