// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:05:33 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
NoOWNjd42a0eZjQt+8yV6jeq9+wQbVcaYolvsjUpMqASKpbBHyFBSBE+JlJcxKAK
xk+7UoL+nmnUb0dMZJk1VX2Yc8EcCIduw9L2XBceaUvnsxZnKU474TCtxJnW9YPM
6+c/dQDpq399JwMYXi5iijoy8m6itynW9raWzNLPTgI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9216)
ZkWK6OwqUFhq7hySqlldi/zuxrFsgkzUcfKnt2LgKCD7x7WH7KT/WSTwcqXafHPG
Izf56xdIyeXk2AvZsnIk3FJSwsJLR5GqeGS86kgZ3T4X2b/ba3ilHHzHiMxMsByV
4vxN9wG5YaSnbiKE6c24faseQJ2k2cL2qtTts+mxm4rfsfkGX/m6aOVqqpey3OEY
zVVurTauZwSOn0zmOpbaQzAJ7CQFLWVALs/Ai94vPYf1JiTHVDiwHXhGzbYbcUn3
7ev+I/pILoUDXHGkuMVILINmporoIbmTOOiKPJzwpeB0c4Tp4FuWh8TStsMWCxOC
ViqYCJ5Y2aKvBVmpdeBHdErpZSnKOrqGO+rzHEIhOJ7+LFX+LFYA+cz6Y4xrrrE+
SstmZIMdTE5r8sjMGps2MuJfc8M/ot27kEk21i9ZoU5HJXdmPx9inl8nJx+ExC1J
dD+JmmfPkJCNEruUEx21Cixw5aTw8bLs1T9ycg0oEiNEJboa8euaKMh8uxffZhlE
sV3mAYlwLAxUCUdXo7TneBy8+Y5nupw2R8SfjS//CURia8fD3HwFAdSQMqtGAk/6
1FDGNPE5WfIwUWUBUQiFFpo2lL9wY8qSqazWnzfQKoqFD/7c1+k6DUKiQk1t+O0O
GajoidqR5jKgCJzjMgFwsR9YJiOzP6lUMKz/lRz+zIl9N/simSP1/sf6FwEIvM6o
xcXjk8iGHNpSNnad51FKxlMaMsD2Vp75OfVai3zxvPyihRQD9uQc2HUDsPjmIxJ0
UcQShlCb8CnUAhkd2X84iq3KvbL1Ul51BJGuRdbLM/7l4ZTm39S11MRrul7bYVGw
1oQcPjdnXKZXMYdfghw5rA6VmiV9bnwi338SwCG6h6MWS6qgiVNYyWVy2iKOzfso
Sphj1hHtPaWVIVBLNCnOWpuJOzTYygpx4HMZHp4drYOenXHmw0ceNpO4kQe4jfSX
6hPoqLeq0Ra4T+mOonV20g9QqrL/Kh+MTJU/UC8ZgZUDRH8cdX6RI5Umn3aMHDeR
X/2NR5DRm8dG31+fLpBsLrtmFu0BgulqXeuDslbtH7CQa4/m66gR9S6Q1ozZBZ9O
9AOggUMVifm0VEM8QaZ6wKqynwXBJTNd7C2IbSEvCENbyYzr9qc1Bzdt4+i6hafc
jW8hgH3NvacBTKnHh3ZsSStp81vLmiWu5qjv6UGeDIlUZtrm+HhalGMYjcHbGAyS
1sJ4SO6EyX6xbv7lzfWm5jwdTUljhIWdH+X6DCqeGOons02DjtW7Jm3PsXltJli+
mT5wl/OumRBMfQ6qs7eEqQK4KUVbmseaV+jKnyUT1UH7SJZQedXHOWSqQutFe6D9
1ydFznI4sBNpEUviVuINyDHVa6204S0VNpN5rmFAI8l6EqTPkx1lbNbJWfY5p6il
MwoMUojaWC2SO/zZzyw7RtN288Cprlnr+I5EhyhQMYwD6nBttbI5dF4WBAx47ftZ
J1DJiIhwH0eharf3203dwqj5l6240lUWz/BR3FbSSGeYO+sfuXNPU7oQagoccHFz
cGsZVja6QQ+uHfH17Zstz3QZoRnV46Z86Ee4wZAyU8/SXLP9VZEge/uLg5J1lE2Q
LTEkWBZaVnJUZeG9YWQoWlsnH7zyaWJBu6KShU6rTHAvOmTg2eaL6o6JKWsKKsJ5
PjsPpZfaYGeTZdjHXbrQw1EWohNGTZyiYo3Vt6uqyeyQ53+txIKQKRH9p9zJ794r
XvJJwHrRv6n/D4zhJJTaj83N/BiWrJfIriOabrwcFJv3RW5AMwYgvOO5AYqWf41g
OtkeU2Ob9EMV8ljon+Ylt6Yu640Q4qZkPUWHFRg8GSiBBqhKsHYfuBnTbU8NPwzJ
wvTB9/gPAFCziP9l2RASb33je8rrVBUmZdv/m+gC9OrntwP2rv2kzBOI9vWZm8le
hc2pi4i6W2I66sMNqjtFhKKuvltkqBYywgT5xK4Z79IQBzeWM3UsjZ65lxkNTbJ9
TgB8gMcFhdwdNLHbQXrGI88sf9Hpp3gGgmg2t+NH+duUKay63olFanobZGfuW8mQ
7itayRaEC78EbYvbX3eguuAjR80pbyqsByQBMZxUV16u85NLz6FLO0M1Iv0R6kfe
0Bq80SDSIbWn4tjulkd/NChuwIu7gu3tBiGiSX8ikZwdeEMw5YL0JvpOttyuIjxN
0plwbPAZ5MmtYQ8bKKj6e4Xdb5CJyjU78hhTWqw+Z6sAL28GyzeOhEePyj+xRvl6
WWS6iQXGjNemYNUHC0q7VZjHOfDUrRr6V0pkG0ea75BGb/mpub7Xfg3eqtNt9bIM
YmIE/+qQaojiOFVEUz6ibzL4zuCHIUOMjDt0fKKYPFI1n6wXnCZBrSw5FKWYJJCC
m+l6Xm8qGxkjk2uwOlLTiOfdesGvnfEk+eGdG/tTJD4SeqUo3C5ONRrOcRYJKZPp
83R1kAwNNCihH9c9DzFDN86jrzGw4ECp6ZLv52XHX0Kej92SMZ9JnSAHmab5+qWg
O0LFPNUWVxUq8673NatNAvmFHD/Tl0S2E9SmICpIZjXaP6y1XtwZ1izy51E3qs6h
fyQtN+GJhToVSJaEfYzEtSp95foeRI91nCypbmd6G+UfBKqUP+gLN7ZncRCjCG2i
YNc9Bq8X5IIBR+xmgo+L1te+J5yxV7xlCEfZdWPw3Ir5zr2GPAS5TtqAuLJIMQcL
Ardm7i5BHFGugbDmw38n2sHuX0fKoeGj6A7Oy5FdUMTpV2SS3fN+rd5NDDvhxM4F
ZS4bk1k8vHhXvprTRNRBECk9SekmgqfLlx/uXAn8fyZtQHz432Eg+i8s/42tDFdr
3QU2nJcPf/HYv4z8wb4Oz5cQlCAhCAHjSNIXq8K5PBr1B/1y5a7MrR3/zHjV/V4Q
6oMV6Th/YrZ3uV/ZSbYu+IuR1qkGSszcVGHhMPNylGEdsaJxkeKB3mfzIOVwzzBz
4GRnYoqRAJJjmvEBHlR9yZAprHlaZDFY/prghsXa9sCVPJ+LKwGj6aVPNDda3ZQ+
nE/vurBtVkw0tLx5uwhy0ZtAAeI88oCZLTs+5DQLHltg3ZVi05e3OPjImGXdfDW7
mcwhd8Ul4lvGLhRym+Etb0pVeHwCxv6bUBxhcGtDnUjklDQMhyQccXC+PnJXNaTa
UjUwTBlidqAguwOnnpgvrSHT82AAbC2Y4VCiavRnhAGgI5aSufs6LFVafKG+s16U
V1oTWwCIvPm3IHGQuGg191y4mHmGqR+rSE15mAY6UE8h6D1HdRBlrc6MjE54mYR2
nJnoGIKmSwPa9UvIbgKRO6jTdBAR3wwnoDpq/jMcGgCxg8UurXCzwcnIgidjGN5i
7qvmgh/jM2bGA7zHf4oqXy3HBLsKY5BhQdr083fq+6JzArzHv0b4mTdcl6+6Lip+
5AdzwszFrH4vdC4G0xhtKSmvhY7svI/kF6Kty9wxgyegJIu8udJMMOX47J42NyYw
EL0yWwRltwxKYCpqFJ4Oj0OQxUxf99ep8oWyIWfPgjKgWzM6SqRipwZVp1sFl54t
Jq4Jvp++5y/mwxASU6wEwJIpxrM214+7ZwUe4EqKkeTB5ktoJIxJUpGgvF9KeNxN
lPAP7vvXvTLoRgy5rqH9DFxXwp+q2w4moxI/uX1zlxQ0h5SBOHGd5TbisXKTL1Qt
MfWiDoKRhLcoIAHdTripGqYftS9kgZOCoM4SrvCMJW4EO01UYbAnpwlpCNjkQwl5
OQao0uS/QYuM+ZAKhBdxvG4PtE9FlBrJapjESlON7XuxyZ38DceY6Hl3swjVeXDP
MRRoVa2G+2QBKZYeAaISh5yBoYLxiOhkqZVDTXt27VnWlYJo3QOlRf0dLfJ+PJqE
Esjlcvl1G+I72Y8QCkX6/NQIDNQYdBxBoEEMtG4KsyIlaPDfgWyv/OywllkjNbgU
ZDJZhLkKd9GjVui/8yQTst+vONi2PkGHz6D9jcGsa3nZnMKg5si+sEkvytFkcINE
T5bH54Am2HwL8WegMZkUqNHDlPdGzPLzzKqYR8IYejHlZYIVAQ2EtcqO0pqqqNSd
2gMBH4MrcB67Ffoq+mvAlKwAtIWfm0x4BP+P0ViMdxcPGWfAbVaQedlWdrm0N/be
EcphwvB3We8UYLn5/RCTw6CCPLbO2aBbdV+bH4lfBvlQF3thAzLpQElxYDQKI8sS
ivJiRjcFQBzsyJ+xi0EQiEozcuzlbztJFpuY7NpNXx1atv5VMB7LN7N0zC2PFckm
isJvLNAOHYXHM4wm3G+4YMxP3etLDy+WmedDFn4ccTQ9MmO4a1VIzuuf3Rzp2jb/
/n5y2BVh42cbFxMKmUPSYj4tMNGMmYOrvePn4cbCOsqUU9GQJ2OjD+citSclWLxu
zJLP2DpJpZo4vZFsOR/TWNrcSmWNo3oN2JCY/ihqTNlhwnagxw00h79PciIp8Puq
rlDFRKrfJe8NbIPZa2U8pJX3y+DMIp08kSqP4oCzAKanoyCyoXSOftZNTSMJu9bM
cGG6M64gR71iwJsgHVCv+lo/ggF5OaXlPQHRfW032kHgc/VQFPNmyb7tJZ177KYS
99zPiL1UduTgNB3gzg3tFVitd42DQ20P5W2AS4HzAFzqTmgOL4k5NXM9lhLeu3wr
KhYfWuxOB3p1p9eMYfzKr4ZrZFxj6H6b4v1l+9MYT/A5RA7bYpi5s9jJsUBz0a3t
DGfHi5fp5kpX2o8AoVBPZQ8SCuLQ9rIqnQYJv3EL/eqCgUEe8CSLp97eAmscUY77
PsClXkfLlAMpnMWJKhbOyyj2y+YJDrLeizxSjsExCAX3iENUrx1CVsgA0xIdjfTW
Dzh3nSTlx9pFp1I+VulXwerwx4Nh+7lDxIIvVvB44hsrUQqnw4rL5E2bmEac1Rsd
fbmprg5wWYASe7wrMDgpw0jHQZygRaAbLadPPwXzpcBYO71NaTtlmj3OIUJBm4TP
4xj9C2CWBenxlO6Mf3DVv5DsBKpf+zaRni5kTR/UX4P+1gmo3S2crU1obLP3ejCo
1WQ5L8m4z//nBOIj9ZBSJR1GK8V10OG1RCNg5rc8TJfbdIcemDQXdI2VgS5H2BHK
1U07k1Tx+MjKqmtY6ddEJA0kK1XKVxS//dgdKocwaI8j7AHb2TrG5QoPFBkoPH1H
YBHBw37fKtTRD/3/8ZMTKsRLDhTMCWmtFfsZrj80GRKSZ94bMDpOgNjqHqpmj4Il
fexkTwiniycgaM3mTqeMEZ5LJ3WgGnyTPvM/kcsXVws7gyRL063KeHH+SQYteuot
UN0p0ZdgD0PsgGIn8aBoEu1GLhOvEBC/FwvcsrnyadHE+puUy549Ad+4bKLxT5oW
lSsb+mIdpRt+LP86rNo+/vqQHxYB03+mdpOzdGNUpafr0EWV0+2U9M6byuEbhXUf
Tqgb45Cm/2K65oiWDk90plevfXRJIEwqR8cUllzvnl/Hibx5p5TFyoNhsbVHxRKO
3AksH2oCdk6EmVaygFS4PfZlPPVQuwXizYPSzLyoDlTaM/HQ49QjxBs0m3y2QiTj
Cuduq1WnyzM19vzxuWu1uThxxkGhtpBKb8HyaCEHjnNdNwFcz+Nc+wXI3Lm7IqhD
1Xo8wEoUFqBAENmlInQVFNY0ikcZjrAKW2DJhZiaYMZik4MtuMqLyqFgAs9lu7I1
phy/+hOLFoIepg+qn2lpEjv0VsW4knXl13OSZbq/grGafzDCmahk7a1SzEYrvRlG
SYxOyBqd347fMFwvcmmgPp0YXRBrC81UWgeUaMVhf4U64V8AsAEPFSwjB/f+PmvA
0kpEYPC6HZEJX4hU/a1oTEnGj7WYvGyBE24cEP4rqNb9mEbuBbYtjC/XkaZRQ6sx
kipk8ab4sPnfFUf/L+5F315OMqwZsdlmnGKTS18wOf4A16lIWRJY9f0S4YwX8vAm
G48H00QVMUK/WNIkSz8z2FaQLQ7bAPHISW2wEK6naJj7ekoR5uIdUg4U/xBKCTmW
Svzcqx0C9MtjYAss1LR9rjKi/148gzyPQqEawlokZ+ieuXYtGGDoKvhE7XjLifcC
WfNAa43Qcd/6nJSSSBS2L0QcWT3ByIIog/mMyJ6f0++6gSABxr+zcxLGztpCd5y3
qUBRVnCjQGEBmfAbEVu54c6fLk+wMvB+sG/fMyMcvjXMsatLIe9EnsYwMf5xW6li
UgLIBLuBxB0N6CNZONcbcDUdQAUbYZqEDe9jhnCsFH0w5RKnwzv2JoD4mHsfKr1Q
XxpPHSLDdrZBIfJ54rd1YOaZ8mf4IaEwBz4sPmRT9OWq983pedBpHHqAC6owybes
DaNctYtlgv9lb7v3IEjnq7LLv/mpIo8dsSOAw5MrO97ApCAtjzKrfJVnDJ/9ge5y
3mlkbSnzlrsF8coMIbXC4yBxypkEpU76aD68G40+5velUn6OLuMXMITr0THIazPS
a6viFwzn1AVFkMpoCR0f8SKuD2WB5TfF/QDiHLy9RmOU+ZxezRi8q2r+lS9Yl9wP
yJt3HyQvYo9qYrZzLv0T6YJLvRZZpmXivSs61jpiJxWZ5t9Xm9P+082uxfHT4R//
KoHhTqSdzGDK8SocBqgEulSi3/LyH1c43YuGoY1ccAcq8ZAD15p8QaT/sG1SDslA
furZBfUq0B96cwTYLV3K1RtpYoxzCA6YxlTCvN/kbBZrXnl63HLely2cJj1ZV2Kj
r6DZ+xAcd/vvVMqr11qPZFHysihN3qom7b74ENCdH63QUugKV7+iwBaHm66mAPwa
pOIxNWeU/jNfmYYy0Hiz9i6pqZG+0ZmHdPVg438jWG4sMvGV7+WCZ8jLX8tFuOdE
tnlEPc8vHEQ6HmVqtEfBalifq09ca4IdUReEZWq5a2kCCrIOzJiR9l8trwhh7q4l
pDEe6Y7toMdf9RZH3yJzhUqXM5OeUiKQiKo+RFa+qp0kU+Gj7uP4FiLt6bPpPOsj
7S7QixlhsIl9Og7YF6P0dLy8r9qg0RiNkVf8ax7H/GZcYiUv3P0wVmFS4L2cDUdf
YyM+gpLeuMFppXVV7hbj4F4Ca2BjbbkcHZiBlHDyYYh613M4pEWN/xfEhm7mjrHa
I0PGYNoIND/eUL3gXi4kRxm/olF6PeHVW5M67GTTAx32rw1QlhXpjSb9N2teTBAE
x6UDGgXBlAB1P3VFiqeCuURgRyZP2d0z/eazWBv9/TRH21+vzqCBh6YEmd3RBXbH
qV3uWVCr1s8XvKFkjLaAl8EE2aVgn9eX8TquwMs4ylWIwQd372Yv92rzdD4CMx5x
pVYY/WMQueK1RyWItp9OfWRlGpFZNl2vKKXxiczI1cwn1t8NCwc5OAdsYuC5aNmm
GHesDhyaoq72/tvCUILLv41iZXp6Rsq/LdjQbmnxQfzrTnFd3S2UBKUNg/65QLIn
aWGt4PccduzO0+TuG788kyieGfaDUyWRx+mWtFgiBJsTIklmCcC2WBNvuTTyH/Wt
uD7IE3Uqr4+DASeXdh1gSopADscs+kQsRIV7KyTXE7WqNfq2bAZat7QE2acmYQgH
Ibkzy+yaeDxVch/17d8gqUw4LYT13CEf1ded/mRDfpQwI8FUDbN9twaiml/dDPHd
g9UVO2EYcQSG6+zjcy9guP4nqAhrFnChg3Fwx7saD2Yz8Rnu2yUu1EPhn69qlP3Q
kVspIK2+n6EvcE4H8Lm1vCfNb3NqknaLDQaDsLnllUG6YyL8FKEMeKCEJ2lohm07
4mktu/FYgjB5JdRw0V6wxdbdsWRQxC3BOHRnhfaiWTXq4hbVcsACX4VBXc0aedoU
Anps9AlIjhwcQqPuVL55zguCR9Omd2S/b3grxTFH4bfmbNE49puYsrcvQpLH+kt9
3mjaNaGyXsGOGEH5LNBz86wWknahKnxCbgT2eOdPbg/k2Cuhm/7fG72DPHnMmX+k
afNhf/ouAG4/PCDGUUtpqmt2dkcp56JM0thFZUKEQO20lRobVeXkr8pTMK9V6LBV
X4rWiiwK1B+7XtfcnxxMAQptJnjAjosCxoVJbEEDodnyi+pE0KDdi7SCypbP6ePq
AJ0C0rXKiSahbtl7qg70Vy8m+tMh6bTTeRCVkMBwK4xg4WoCNZeaRn+ZDCvMe2xi
52Ry76LNT7eBU8QeYRtFyb4x4utBoSLR/ih/JPYWVwAwrFid/+T/x5M4iKgJMMaG
6DHGgazqdQsQG+eZuJUxfdIqTn9XaX3o5f5RyN9xsGmLGEmv92ID9rCKJ23GbT+F
V8accQmt3teXl5TKJriggj+kao8RLI27CST58ZG9g3DcKI8+5pfOUlKozfUmTgOZ
76RahRTJXknJd/pN/iYtAH5oq3Y4qALxsnbTx4DJKanDJcXAhH2pXbJkGRFCPPkZ
BCmjmW/hrY6u7I/bL0K1G1hpbAgM11ceceEmWDnZIVgrctXDeuEvQ2B2k9YfwYjk
B9+w6U0wsxPOVvLEZgvHdwwR30WfgxepFamOVOcCa/h6yLQXiXXpMCqze9myX01I
/DGJkajpBjZp3OmL972tEVjX2gnkVR6ajALHMZV97IKrXf60H1NjalKhXAftZ2mG
sqSBlkbJCQMbqx76+zM2bVeEfHA0pxBsG4zgkcI8PvK8LYFnpHyucVOcnMaHIv3X
Lg1m2Ab/SkETc9Oe09cw8Yw8l85dQaDSw3lN7c18V/svoVAGlC6x+J2IfwkVg54r
xF0KtKnT8WvI/8Z+ukJU+20QuSuuANusxqirc6eBUPR3T7BNIHOSorPX2witYMYt
n029s4MSOfhfohecLXZOSujt+tVVl0lXmULP5RWUABbTgnrNC14rPsUAihYkPS5V
OFh4dVNEEEzRPd2Vr283seOtOK/3WsLYbWQRyCuwMYmpWKyQCm0TP5dt40X+nYmS
rwyj22I/Vg4kA0ef6t79ZWDzXcjgK90U9Y9q05KuN5/z9K5zFr+t1k2pWEyU76Qz
7/T7XVxjWrzPfMOjgaeAdsG5kHyPjnla+z8JkNXWK/vgYkw+4DYwzE5f9cHmfrJY
QiZm1eGqcfxr3pXHk90vh4huMjjUHFxj8ETkGahT1ZdB2SDamowmLV3SGbpzFa3B
sz/BeTvsKA5IH86ha1W3pXW5kG1yHB/9QX4bcoogajnhgnCdaIGHhGzWYPiyzaM+
58us8Y7dy1ePY95iDZiDkwA2txuygRt0Y0gpiXiQ1IuDD238XGhMqVxFUFgcqxn4
+wk2eC+4XJOZnkBrHopULRW2qHkZlrMLFEHO9+WC4DUbTBr4c6UlNBxcJfb+U9U0
JVojHwbxzWqUiR0mK0mNCC8kUXKYrTZnK7XfwSRgMhC2p2RuduBfLzaEKm1XmHtv
HqC/Dd1/D3vUAeD+oVHkgoLG2DbRjnelhyrBiCqbzKxXdTxJLk1qxh3M6InP8min
GtuOyuStv0M+hMy72WsMCrRhoXCUiVvULSnkQz8ZX2dZ/sRIzq/PC5CtGHX62n5e
KiRaakaQ1jFBQgE4SRH64I9cnH0AgXbZ/UMd04DzCvDGe60trxFG9S+0j7bQyqFO
He5kBgvx4+TI/FwSH+SVkzPoVc6b9Qjdp6xTTk5ICm69HLjhy4clvTt7WvJTCXWA
h8rkMJVdyS2ovpbkt59YvEh0SUpjJY59xk+6bis5qWNVycuh7hanm2RnfbpJjE0Z
+APU4nnwx4h/rpn2mMjC8I5xTfLBlzPeBSVMa0QIOfnLZMYa8jiJ9es2KSMA0sz3
SveJ6B/ciGaYb54lGJcI1owzLli2gVXy37XenSOPqt2FH43TAoWXflnI7hj9l/8n
REF+JM7V0JGxK3eb1QjYBUKL3XJPHyjyJzA74o6UbN7KxZTPuX1/CwHJ/8E2c4oy
zCDfJSTarsVAj2DKKJRa7yt2COYs136CngAXNCT93K10pdIEj+RY8yQTqZuaM8lK
3C2OyzemsW3nrIuAF97My5uhuZfh9jktuP4LwicXI/sk/JAOV2pDowUPXGWeJJoK
Cqci+ucqQH2izKSIPON2Fb8G1RPxiEyRgxM0Dhm9gYe8qIkbsijGcCxVfRBlVC7J
Cs0s6TqnQKxNomTi8SPHmV70wOFDs60HkWkArtcFRBRALfgQEugSPalnCjyenyy7
UVBp+/l2Sml3LNXkA2NXTHVKJYwBK8zMA2BBou4c03MbrsU09QMBAtAa3M/oXz3R
iB1YMyzsSC1DFbcl5r4ssB9gc3v7GkZ/9HIXVHAFczkvw5UDcB6Aurpiv2e3f0jz
I8qa3EysA16rAe/2ioDoHUuy93PFWTa7J2ey2lAWnXSXtKRQdl627vL7FToGtNJ+
aE894a55oHmrAqW2OdpsqHWlHNCVaFLf80ACjJU1hktGUzDlO1CbEddj5dFcmAZK
8I6cs+vPLTy3kgH5AA//jyCPljzZgFl6DUEy9Bm7Gyovw4zgQmb24gWu/DvdIbHz
+k12/vBchqYtMSrtGnZVy7dcR73ddXstVx9NdGpEsO8KORhMjX2FTVqyqpBPuuYU
ssemRIr2mUpV7CJhoClha2HqrjHdZhDbNN2s3GXxpjKAIFf94f+iUZpVle3213+g
8YODDWqerB4xT2iHWnXAkTLl6vbTEI/OQHwUEjVYHQCqByzlHwbtFIXNGDhReGKE
LpWNvgTp0NY15Wom+4EA5CmSjbLuE3YNgxEimQVURgGphhpx0R8lsBd26gIjoua9
1rbYfTHVKo3+xEEIWMpBxdFekuoJOkASlevLZTr0JL6vrmHrs6IPhRzmCyuNpYys
Cv7lQBo/wQqdkU6onYToYZqADmC1+T1I2CjNKn6Gp5iTv7BRsCqdbGr8FBhiI7Q1
YDgELEHZxV3j6MjcKJJ9Z4jGaEYVDFGuRDMB2Ee17yl1M4whk++cEDjXnuCXatBM
xDfrwLCHJB4zwJ6SWmdD1w0NTZSWPbr3S4XzLKo5yilDmzSxeOz0KMFBzeD+v2Ur
nDveTP3Fu5YVcoQL+IdpgbrNhvqLj4SbbGM2aCS6e8Ad46kUc6gTxdvNfaVfcTeO
V5WWEct4LlGCcyWZSn+ifM22d+WTdYbrJTxp5g5eNM5sMFmlERcoCW1v4CgLjLu7
pViwZxGaCYkdQahuHd9G0X3ivvHQyfmimrbN0l7MKJMjp8GjCvXwIJ/PD5dgLMti
tDa75dzJWxVMh4W346LBnRBRu32DY24ehhmIj6XFRSeunnu4Izd/i+nLRS0AADfD
6C1UTZ8k2Fg9pVe+ufIfXNLit0XM31hqoUqYAID9JNG7RSOX1GkHZD51hn0aM0+m
tlFSilkr6W7PQg/368crlyyHXOB7LMWD/F4JN8Hzp+mJEWEMaY4PYXe7PHw0uzZM
Iz1XVr7tFhDtJTEqcRjkq9P2bCfpa+exmDZQDuEZBaUkQSuIXcMZ36vTb5yJghH4
pFv1jRR5q7WQ8xp2Eu+OM/tLJBjRgwuyaMtITq5eTlidoVvRtZmQaWSyOXcl/da2
wSqMsKsk6oJFZvFc4gaUnpySYBPtt4L0OhVQPHeUPR2XYz0DlaYXfGzdRu0GIoA9
vTnJgECfAP/kO0w+dMbwYhkIS+Q55cigb7jscu9mCQRt27UYApd8WKwAlt3Gk3EC
3nIUknmBiJVleWyeI07cKIuITkh12QknNSRm0E/F5/6ZwqsSwCBhnRXaKW7/ZH8d
ycoaAJFYt7ycRzS5QTYwza1KcqfsE1lX+qFnIv0c/akRDcEl/7iuDJtcOjnZGcMC
OuU1WJV7IT82dEXLtQbJK27kRAbwKx9CUuh/HNERMRG1BZv6ANioqA8p8z17oCqu
cLDKK6lGGcRL7/vBg2CbeeqQ/PhsziqixmqJ0jWOojdD3JcUpxf0m82FpyiHyDA1
p7iF1mjbSdxOyXKVeAlNBWrmGvYw/k17TwK9YxlJdo20GONgXstP6UMWTnslgiV3
erqQJ+9jq7g6OGluP0sCWJ6C8SysD+5CPj9DmonOkbLc85rTD8iLhW3+mfmTivq5
wBjhUEmhgkdxcaMRffzxbu5FZLknYTUqDeZED22MrmuwOrQgctdVjcOV2IJmHmLk
xxHTta3LKrlZrhM3lQmAtkVVWRbT4aT6Y7oUWB6oLX31osRGHmIbo1wte0+zUXZ7
p9tfruUOY2ZO+AJHlYZDet09FQg5aQbiQn0E+3aNwbmIFhGLzdFdJ461ul5+xCK5
fI5zEESvJWAHgi/QGAX1HeZ4W/Mu5wpe3s6Mg6LFBZP8HQeaKJ3Gwlk2ffMRlvmJ
kikUPMBRk0enboymmyYnymn+oUlPkdd1xsCeHMza2r4fjqbnI9RhDhhVsi5XAEti
87aUBlr3P8cXLdX2XTpSxL0vN5a2yWDrg//7FgFXJz3jTilTU9xCqYULUEZ10+A+
`pragma protect end_protected
