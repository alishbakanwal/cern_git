// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 14:01:26 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
DsvB10fg++kccoaDmDwxZs9vPX5yoJTUcToxNJTw9B1l/6NYAFnG1uoThE0/PbHl
wLTBgs4I0m0VdhZGS1HuAEr9zn1jKnf01GkUSTI6jjnSr52HT2y23PGM9GTERJ58
2YPXmnEV76NAGaV/GEI81+kmtooeLk1mQYIiYRd/scQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 32176)
FOXX/DE1w5Fo9cekmOtUz6CbSkC+TEYnhDpRnfQp4W+uWqMgTU6aIhA7KFwWhWl9
7qS7yxDeYURPV5vOsxDZcmxyafsOBNFVMi+Ig5GBNGsjOKwd/HQwBPoc/3ze6J0T
Zseke/DnIYGa68AONbaz5d9Ghz6gVr+8PrnAYaRfnxIlCqomp0bP9gWiBBPpYNAC
SkcQtuKTObvBmcHlnfyHBDAHnJbK5Ws10OIC5D+kjwQikx96vI63aLO9mFFDxji/
41j6d/IFYgRloov7y/lJfAnsrhauxJhazQj34NFVQpUM9K8eMd9H28cbrdfoKbFT
garzL87bduekHnnvj1BhSJo0qEmWXYAb3CRlJ9wlGBL+mKPyNjSD83K7DzTxnWoc
1iENHPxrYbE8+Ak7LPbgcMsRo/47sJhvJztdSGxu0+8wZoeJWKnpUKN4eWm+mziu
EI+m7JP8d7YqXhwNIXuIZfjm8Zb8A92nWI2p2+7ROxYJZK3UPB7GA9K55Znjff2o
QJk7/UGfm/oddw48c73TtEyEpG7JPMjJ+YGPnJ9N+9mV429x1f3/sCDDsdHpEuJH
Wr7Q8KAtVgAXLfcWahYGcOXefa0B0whgZmNTvzwb9CY69dOr0O6lAPg+jcIjvLSZ
HsjyO6Svh079jTVZ/krtYHDUtxDTyB0v8tZH14etWTqCRerRif4gnw1jTFDUp0Ys
XZ0glZs2WDpQdWjNo5pydU3166Sdw4u6oxD9DK57g09xH5fkasBw3JkgYviu3CPz
lofQa0v4oEkMoixVA+ymJRkeIkVgOHPVnuMagjDioX0xsNPJt6Vvhyfv2IF1EAXg
tVAbXfd/+VMskv9GdkcipA1RIYJyb/D7JMknDyckAa2cTlDRHZq7VxzwJ87bn6l7
7PEAwPqA1+ZD3dZ3r4L3+C6d/2SwkiKpZ0VTxTf7Pmf6qIt27H+xXglj/8ncuzHQ
+GPfVaT39kHQjIz5ZmLWNNQwc8y/yxORJGk1JW5npqtSSeJ3xreDqmoGnnX7wEeE
RbEq6uAYKP6X0hqsQ8lELpGqD4neg0ht27p54+4Cklk3SXe1+92GQD/SPUTS1ocI
TCppsd8YBFFPQhDDC4V6PoEt5DuTxXqR0UVVww1sSqwSqXaKDxNFHrXa+f/8RkyG
XfFSuosyEKFGibAL3ri65HM5BoIDTVixgak3/va4c3Bkddd2vSHXiZvwMo+tOHNe
m+oaTg2hM2MgFDdT7nyR4UpEU8oVzIXnYnOV2pwTbS5DGxcopNCI59ENG7VKWyPG
rXtcP5sSI9Q/8Dv69B0djemoBS75Qrh+6iTCOrboUwlR2FyD0BZIJ6O3PqWpRoQY
RQ1FB8EjknYF/YGtVPrP5s+wMfDuo6Tn8gYyEUUtEzMFIV/2zqs/SrzFGiU/sXyl
lVnqN//65EWIXnTiwv1SfvYk4IEVrWuf0CdHcIbIdTzAY3pXStQbqAxuLAOozFzr
mXOKTrpOynphfc92rWFbsBQuweU84ykDnclaAQfy5dhaZjcAfarQaQlwT4SyQfMO
Huolr2pmA1vRiUO8npo5Duuc+rXlQSOTIsFQg/fff71oRj9E2J1CzOR8wr8+dq0u
50GZrkZipCoR1vYg2aYSguy7kfmBCtTzTYXYzj+FRfjP3OSQ7pXW4JEgN6Hoyzij
YawaDWKk3vOsY/4KTQVXY9ou8QIgda52rVr3SaSJk/ViA4CwhgVfRxuwrnL966zT
lk82vNmJCB7mVzNRrfcwj7l9Ugaqp77wUV2H99wudHj4c7VEw69p5cHNw8ck2N52
lFqZcm9QETOC7e6LG28B3uMPLzkHhgRQvpLLSwLlEPJxVv7E/Zo+X7ZQ+B5MqtUU
J+OY9YexLRV8T6er0ZaNfx35Sj0FoKRuQiD1kGIRnsJHCHoyy6rDBbMjn1CVi7ky
PHWqVoLL39lo9khOtJ1B+pMcgproB2kG9Wa/+BOHw2EQFSblWLkD9YNZZFPmbCyw
uhsUIltziPni7SF/VdORCMAqEhHA5//8RXjvzkKsLzRTCdiXB60z27NTI61GyBah
ZCXKmiRQ4YiFibHV550jb7PdQPVlEZNorcYg9+Lpm6SHNvQnDGAAuemUi1BaYiiT
qBEES6KezvuqIezRxdDuBslChdOXtrV+YRA0W0MTmS6ObhODlmMHeDxCJe1UWIQt
NnTvyDQ3XQm8lT+ZklFo5OSBkO98YzeL+nEkm5uPO0ivk95i2xInycBYOCeRxDTn
PTfZ62LrBcZgYDcLpiYKvvzequ/he5gOQSlZN6m3o/x4YdJNd6Ma7UIn9pWHVzDK
gkSk/zPDhwpIwecHfCwadxgdbZ6Asf0xydP5XR5u67HVUz3HH2Do9vL+uvChWilt
uZ/tgItv3mC4eoCRH3Io5jpEfJ352HplrcHol6QDGEVi8JGIyoYEGqitvl9hSS5f
sPInncz9UYXSCTDu3HGrmMwNI1JTFp/Nzysf0/RmFHvKtVG20PKFe8NLr2HmFZIo
REdTzq1AZuZb8Aq3a5U5lhWOZJ2dXTuEBnIGIB6jahiBr6dPbSeYuvujaMtVrLe2
aAjEKVzFYPtiLaYaIXiUtZ/0PIJ+tjafiTNL0Yh4UJ+d7xbfraw0FyQi582Uqmf3
kYwG0wAaSulia3lYQhWKqYH698IhnpKvgH8rrbnG1cVjPILOshdQlGvxlJYrzdfT
Vv6cIzWnKiihrifGFEy9sLlakWalQMcOsg5Ntpbbb/M5ZTe1OyTiBad14xtLYtmJ
wQyKmXcxD4L1yzR1raGZZdHmuVstLtaUZ4LXuG1Vjs0amqv9YDE0b4y3wyiwEyYc
8Mq0obwsGGLbnX3ZB/sFKUkT8x99/S1fzDv3aRA2irUCCpcfXyvu4jycdVBXF/yR
IjGPTsfTUQ/JJc6Z371AdywR0IrXAjmNXkkj3qo9hsCbh/0ztwvsnDVvgjwtCldl
FkcU5he4EP/B1cfthU68NFnVZuWBMO+21dbbdBF+XV65FrYSC0tUb2FOjYnG0c0i
OcCWgKKevynSKTpO3OAUvFaFbtzApi5vdxuQ2ijDBdV7GssH79c1dUdKjs1HiW1Y
MUgyPWugBT9HMOPo59JYuJkLLb0UJkb0Rmw1dnV0G/XHfljVTkESmVIkrziE9q3/
LoPruGL+QjgtEQDrLn1q6DAz8bpC/ECULK2Yy9gIkHwEYWVZ8Z2pxwjVnhqiUe6n
LbqouMtxJynOyFT3WfpBupMwPmmeaOPVe6WVbNXV4qWrDsEZmBn95Pu/yR9cWYek
typEZ1rLW3ibBhy0udelky+mvU5V82wSOA3MEeYwSoaS2PS2AApE04fDtJZ36Loe
hPHgEDulrJ+CDqCFQ74s+BLXbjUkoKOEIGwfbspdjnBkUE7FLRsHpIlj+tt/TBS+
sMpFpvgpJdBR+64bLEcF+40+jsZHZF9e5zQ2XsryTjGMH+GW0P2l3KFhue/MaOpV
sO/BE5HKWNLsx4NKfHsCN6VoANDYWGWYICqP2mxNzcmyiLqBsAG7fBBuoF3eImBr
ye3hkaeSI6aNnnQCBobtdhUP5bv9KdnprFQMrp82OxetQHKkt0dggcsOfLdGqJ+l
pkeuMD3LkJPUcZhlq0JfSYgVNlSyCWRY6uaIGvlonlQ5TGeUL9+IJF9voNOj2/qi
cmln7HihTLesiTGYpnJAcP9XTkCuWI3OikHMjJFerf4ms4i4ZDOwVFFoKDZYtUOM
C6Q8JhGgJFYN7cputTzR97FADN47Au8Z+lBwk4F/weRIAvmF4GYw9hhnSAOoQGvA
8pCGpS/KGThRihh6RTynkdAVCKvP7cU7VShoG2GvqSs1vjkEWBTqzsSDvMOBCDs2
vMfo+qNluHxjrMJmKwdiwcVDDg8CTtQ+cDE6ITnzjF8/8g9dvM9iup26pxfwH88R
OBoJB6NIaisZYNWMlpnTsYiMbDa5ksxroocH4pyPzC1Xd/pqGKublbdHYEtVCpri
vdJIy0DRlAes6K/PLg+RPUB2CvvfiJwrb5a5f1OV7+wv2u/9usGkCbqBeLlS58KZ
rpYe3OliEIPmzkFsf7J5rUWMkTjJl2ltrIqWyxia6oa9Q521G9XT/+BzU/0XdLHF
DlegzZVkk60DF68vvSxh3t70XzjxW6q7uzqgNqzaoYOZMNGS9Ad2ho/K9P8/Oxjj
wfzEeqmSnDCfBP6rwlVPE02u1TbeAQCotSgKOArjKVcewZEnpn57Lb4T5kcCKZ+G
lDeye3pS/5Ni14pkSCIqtJBzkrGxuxeUwMx/rBkyRXkC1UKTwl/wD6QZQZ+HESlG
TW5VXM8weVLVq1qA44kMSXL/uk48IHvAv411klGCrw12spBVL4/ugRK4PVuPekEy
kHAUzCGPYatdByLDpoziQqA6reMQ2NdwCvLL3QuQNTzOu/s3rIPsCvPMwPw/7ohp
R1vBIjQ/XChrmVzZDtDPJUbcY1iISJFpsWe4pfz0uTnwvyO2ub0O9IhsJlrlbRuF
7OYaDrJ7wLZlMRrzF5kXWRpwOwGNeH43x/INIGssjAEQhXytmx2pKi+2FstJZEr4
yHAHNFUg+9s95YQnoHtIZkC5t6fFq2SkRsdMjblfxmi9M4W4HhAmd9DaI4ta6eqO
WY31h+P4xw1xdedPlWVt01FHnge3DG1IXzlTbPBd6b4zySrGnEdb55POOHVsa2/Z
EKr8TV3ynFIevsVsDcqMZhM+GcdpScjzoQmX/KHHhe53spDIEWYiH6a3++pnLyeE
Zh1e0gUnP6Lsf4TZqmwBU0HVRJSThspsYjFUFwXFqaRl9J38x+R2oyWv9gGklquM
NxKFfLxcgLxn4LzzZb/p+Tyv/GrmKqRmIqMSpIHCNLW3f0KOV1ar6bbcC3mc7A3U
5jukt+mvaGO7PvXqbIM/St6T96yAoBrphPP4im62E323W0FuAvZQepreNpw8FPUb
LI9CucjNRhFVNVWSS0LExe9mL/Qgxt5M9iwCzZrk+ToX4YwgSxJc+iGnwv89P/m7
iNe7YPohIcwBV0gDozDFPtULN1eKOeKy4JiRk/pMQIqGtIjdUVuaUgFhV/UPMJPY
WVKRwUs1Pp6tQlwQ/KKdGmO1WUaRo51ZvjD4AG6DPUoXi8j+1z4TzevIj9tubJB7
jQeonLcUvyZVHwxODwAzRmB1VBUdlj6wVcbTIEK4j2bqnyFzJiHVcr+CKvXZNxwT
SESL1+nfVshLPXoCqWx4nScR5R576n0nkpzJUZas46Vc8BPUKOfsvzDrWoVza5Bj
rc1e0hIos6avZ/ZWwGkyJJB3YKq5NonspJ3g3VXkaDP0tvSiHDduShESI/kZWZX+
NUKawUgdbRB9VGlpmkzFI3JaYR9+PrDhZV8COllPKwKy5eIqBducMsKut6A+X8/t
OcMcs4gM7tHZosK2bs91vRFCM7gu+S78+l9aOaiCclLJqBAfB549tpCiKdThfo4r
jt6JVXKd3r5w6KNrOjOAg7p7eTq3ZI/xC3sUAhsPG3rRz0bPVkwOA438F6yn4YJK
vNwRQbn52mH69v/am3MOUnlh4Bpc5zk4ulBtXk2w9x3daN+cWPw30769nLdASIa8
2O5m3PN/lkg2On2jjM9xLN6qlG1MCYO2uZEISzyomsCT/y1rR52x6Shc0hXb3UfO
e7OFBM6sqT5aKMrMTn3R4F7CQah6YiPlBx0YNRDLsIQlGnei0qhkb7BM6+Ph7+pg
TfF9BkaDRT08UKnEKCh3a/Q74snuK8kVnCz/5W7djpNqG3LIm8wH1QscezkMKo6g
Ys/9ahuyf2RMAgeXQSxXaRQKaYphDtPIu836QRmnoX0i1UuFS7NAL6X2//CYfrhW
PuZ0dHvyBVxtfZEvYk/IsNrXCW/U3WFwOAMbg6WhMy+XPJDzvCaDB/xXkAo6AkSe
uDL52hB4zNvQXfEQq8jiB0jMikgKEx3MXAfGhNv3tp+hbMW2Yn9rAouPXwNddz3B
IT+aRKkjyPGb6lXXBSdkR3uoqyxMjA/lCgOwsDWQb2AhdW/QVyQ9m9ui3tSOGnw/
fftfr60YSXOjLbNWW29aTUklWQkwRZG3xt/AMPBHirpixgjfkSXMqgU01Eop64ZY
so2QEs1U6KhhVi4fgeSinw16ujeV8c557qqK26oJBshLejAhwBB1VUqOIeicHA5X
L13Ri+UtDER7azkVT1a1QSh1P/1y3K6zQZ3V6nPGVRUyuW4c4qHquiUalwWTCTps
u8BXvkGnk0bWOCh167jhtGmy0S1qM3iuLb2SAsVp4744R1vv+a8/0EzUG419P0lG
vwJ3rf7QpH6Glaw+y91G0E6GqbJ7v+gOHeO/3zC8cjMm84MWrBQII27VSi5vSuF1
ZfRxjKzsHoMoh66EbjHBLKcoKDOtRGSu5Jh40dZi9V4OcYKV9oTw/3vqdt0l2Cmf
ZxS2ztl0dwjNQ0h/hR6nBDjiFIYVF/QtDpD4YWalzB+CQgpLN3onNVsP+wd1f0wM
kuFOx7tO4T9IzXBuzZ63b/9efk8c8Z30wFCLGaOXeUfVp+1J2hYbOYtL0jPXQwFK
O3xi3gormYdLzDtn8uqoeIIfHdeeDBndEb/lXqxnmRjLJXbN3ndUs3bltaIDTrpg
l9pc+OdragfYe7cYHGbYaIVpxsi+azZg6lj17fSQB/m38s5RwzZex3TKfkdYJBCF
SwriLM+nxSB8abAC/ZMyAk/IzbhU6aqeJCkreT7rIXYDSCvr4YbtQH8k3dL/s2q0
VghJ2gxmRlp9qid6oNw83QLipsPRt+teamlPXVZ/Scf36JXGqMxK2Hm8yX/9H+Y9
IXkBV72/gJhpikF1B2xSKD2BnLBllte+/DMWjBSajI7CF+SxpB9TpZv/+gNbRYie
p7FW3Fkxu38vgJYzYnAEj0gnSWQrofbHara4of60b0rrGQyYrH0G157H16QOCNOL
TxafwCsoVxCR+2FUvDpGD/NZTYLJLfwn9IjcuuHGjC8BGIbiMA7o9GfQ7GZ2KqBJ
Ah2nWWER8wPjNtM7cX2x1/+Lkb6ODmF2d2t8F9IPdflUbXssY+i44ug+pXct7xVk
J8T79WewA6B3sAFhGvo19R9vAqD7a8eiKefCh0yJ85d/G8WJcrzhHBNaRFbGffe7
9+W8EhxD3T6Jlvwpu7JrS7sCMLzM2VWENt3BOkg330Gappzisr6/r8ojsKFTBZIf
Cc2rG3TUy3fMA9Bo0ETPkYr1U5QBtNg3a/V4QAsXTzqKTfuYaS84mCYma+9pXPTY
RR1z9a7sjp8nMxqHWwj9vgS1O+hcGkEYdKAyZCYeXzHI/RN4+XdmR2mQ4anbBLGu
zQvM7h/Fr+WK9PbamwDBmMFP1X1tubpq9ByvVUZnqlyWJ8ObhHvK8wmDxRMEi0QV
7soRhYQvBxh914cSgv3q/0UhnVETHZc/YuY6UX6OyulxiSy7kZ+JQPgxw0puA5ct
GyoaxcGwInNG/GmYxfT1k83OGcjfD+FguCuhjseplw/AIq48qB0kakeczh7z3bZY
dcXXWWmsktWYbbzcqFMXvqfTNUnBOTa7kjWvMjMA4KdVHXKcr2AhE21Pl1thWdjV
9De/Co3dlw3n2E0fPmpCET9j8sDjyE90yAZn2ZhrPPskXN3RkXmOXnxT1xhOLQIM
abdCL2YwHEbzwY+1T3k+B7YBDV/S1y8TAN+3iPGPZNqxs9h8ZN3UZ0f7CwjEmLno
iFRRlEtWhtSmKeRYDCpapZwU9m+HtVjHr3LblCQMhf3/+iH48QDC8h4dvjygYddc
5OQ1B/7G9ZP80k97UmpChgfoP+E4jGkoEijZW0BhdHX0W4hugzf27/f3Ide5N1P5
3BiCxMGaXP4wkzbJmyeN5GwLJFb16cyo+4jiHufgedfodvUy+KxWJz3mFg0ph6Lk
9gA6/2Gvk4tqFpY2nIUVFz7IJVusFY1joNMmpbOHtoHbAQRJAhWTrFQwF+c+l1Xs
VWaKlgX6UOzZokTulb44/b++J1xpewHV0iPZGCLc6099UCb5E2LjIkicsL3cX2mx
wzDcqoHcJ0wgbpKdNhYQk4g8ozbWNTw/v0bQyIEqJaL88iQLhA46FrDdAbxJanfE
dO2mmyK/tA1FjamKssFTZlyK4uw/d/K6iL48WEscIKpjDjBOvnJH1Lyr94KwRZxN
Ybg56nibtaFxq4cFC4H2bqFXPBQmgNYFhiCS1dYdt78JqN4gubSoWPuqZQ+L36at
CpsjmIz268qdV1AePsCvKa5/oGKWxxM2qB2f/2e8PELXzzTS8WJzBNQa/8rhejPT
QWQGq+ZLnJd+jZ1M6iyrEaYW5u+ntMT+mvUaU5ALUqEfw8fy89225nUQRiG1FFTZ
PfdAYcv4jUeUyxRq/WrpG5e3K60P0wl40k5HxxnmQkVSrNLzqLmiEiFubb+2t/Cn
q9jdUJnHGX/P0Pso6R9bEOTSwzLeqHrB8F6mGsFCmHusGdtq+WxfjyqFG1cnirzK
MIcRP6DxVBmR2fEjSk31Mi3S71+0BDIrMg+gERb2kDWqcO25pWU8bg1VN9yQY5LS
zs3pinRijywsmVTGKy55/gBo6ZJinxha0IWAO46tZrW9NrK/N60DARV6mvwbCxVg
FNZFz8A2Wt9lJVZ9UrJQsDtam5MzbVjwNLQaV5N/f/WNB35SuxJcfC9NM9gw621b
d/EFDafsprznvE29Xf8jIAJUlcAM7blk4InPpRfn7vhSrA7Litd95ONAsvstnUyW
Wg1X9rnIGeBcWu0i44+L3qtBtEcUGbOqFNF4X0H9vWBQmPYukqEoG6xMXb8lAnJZ
jsOMaLacE5bZH+YzlJXVf2FZcgobAHDTADXXANy/BDokPLMXs1ZxsWyCECezRL03
WTIW2Iom+N+h2JYDpNFsvscUGqgS9uAX17byIy1BIGWZurqYBYu8piPT82reDspd
GAsvqA+MRV77t6fRQZg6GYEIZo7Ph4+YzUDXnKyhXkTOxK2o+QbtUSb/x9yblWxd
2T30tq44H1aKRzI1oY/85M4mZfinQYJbd8qDb6w5oeyB5Loic0GdQnaJy9tS0tmj
G31cCbCBnkqajXBb0RFZ8PAGKGb9WlEaaBZvsoP3tDjJ9wKT3g1UXU4ofKIQwAs1
DuawGC/JrOiKEROtjUGKeLAygnK4Q/JS6bq49PqRpZ4RLDgFtNSWDO9vfTIHUIat
EOGUEXQwOWkSDZN/5+xQj4KKUU4tinH3W+555hNdk1oYZYNfJ6HpeJB5JPrKGwHM
koYfly16mhA1R5u1j1tnKBKcvMSimXnlCCfB5eTnDyxPa6+IZa/lpdTz08MKOCzj
xxt+7TUBp3ts92PM7vbiBiXwBSpXPmT/CnMVgAl9yX8Q4ZdkGoXeEKuPmF2Gkcsw
YDSuWsoHNJ7ZD5MHpqOm7j9yinM6knT2ZuVYsFvQMfSIdUjefga/twDBs9c8dce+
RCvPR4+NSMutMDM5MoabjNA6lKy88Skd1yHpO86ueP8+shrbOELxPxafNrS5gxVz
U7Ng4Oit3AM1W3Du+Ed0O9PrO0z4++sCb9SI2c0l3DLakrENanHX8dgSqAguytoA
NpbRi6qj0KbJTx6sXRvw7xdU1KHKFKfFIWJFlnd4/0+KV5w2MaLJrNdr1EK+U+Zc
V4T7rilp4Gs2IPWUFP9N2OpCFJz8gxyIyWVB26Ddze0u+GWYR4Rnrd/KkXXvH57V
9fNFV3iFudTSNdiFd2YT5I23MEXtAKHfIUcfWLnRjkV/hDTwQ5PDf3FlpdRXZT9e
SymVhS4eZ5JJd5zcDLrRZ0/GdnRZCM9d3XEMMjBc4P/360tab6pWBvp5KRgI63oH
gAjcpCDrAiIn9tKoSiD2KQ6ykMdT3TDmrmJF1auEyMYWYe91vWGRjXlHqgap/WR0
HOICjEfto2LMe3NdJ+b/A0zSd2zi7jnwr4SjHxbqFO9x60LtIzvNefW84AGra0T3
vy2vWs1WtY1UsYqZueHuL72X6Td6utZsD81Dfx9NCcmkvZwKzqQ/UEoZ8AOu+0ot
+E2zgjCoTMz7Ee0yHFB/zIPSAdS8HQtL31K75upQCYtosFSYl1t3NR2Hron+ktIh
Q+oKKiqkXLJOeqh3yb9/KviU3L71rMB7IJiGYsQ8sIhYMkjRBhg/xVj7MZtU8Fjf
Ck+uRHkyaoUKluDxuIa57U1sbXUIoVN58EDA9IRsxqKNV6LEUGNRopZdfg+2/H2A
xGyvWG+PChXPP7K8PleIuDDf7+pyl9wUSTpIkmA4S4gCpWrlmV1o31uU5pf+q3n6
2QF+J9OehVKmwsAMIdRopueSavRU49vujTjbbHiFkI9JwjxfVFyJam12Seep+wYQ
LJIL40Z3qOrF2opO3ouI11DbrlG3PJUBIgN/JJI+g71zRdSuUQHn4LOo4wPFwggN
25SguVMuMjWGaCD187bQnbwXnibWR7GHsEeygmoVRSP7DOZtDSloLfsVJ/kifghP
20vOzGUso8sMW1a96lI7VqhGxtryv9PLpf7DXI0ce2E3ZgwCwT0Uk0vhS/pJt3J/
STFyXwshcruTr59nmFFZBcGhby9wltITcVQHvr5M5Lujh5BzAVK3HHiuqzf4j334
MFGxV9+anLqo5BJOztJPtktDJRSLFE2xXgy1LsZOXpRME2YFhl+9y4Ib1EcSWEpn
yY5UItoI04JKx7xFAZwhB9hF6mxbem1aq01LxR3iHhuA5M03aYzHl+ALLk5zmj6d
+t43MDz/4b7IIXoX1gTdSTzISHdmpV12ZmqAMd1kVAo1UqLNJvTIeMXeoUE4kpaZ
698s826Ofx0DP2BKPS6EvGkGAjQa42YnhdHjs7gGgrPViUt8Qx2Ns+36x0EYwgiR
nPTe0qkFJNgUGloyeFi9/fktLkJp/sfPdPgmZzXj9ICP0RI2F9aRDc+eSKWo96UJ
H6/CY10lDRlrbOVal3RaOdW2fBrkjO35QiE1Vq6877KQhI6nj27O3uUHoCPFc0mL
MXVIPcCHqdkfO9hO/2Iddat3Xp9VO3OMVYMxK3Hpp80BvCzeYCL1xak93XXUgi6N
CfDb0N8vXlMRVFwiajt5BMlx+04ijBu1mjAtQFrmgPa/zA8u+QKPNZIpPsOLb6hW
UlHMsrC60sYxwF2eOoday23kYBsjzN4AOWTSIxmG+w2kXn4kX3mf1dKYqcQ64QM5
bDsmZD+gbh2i6OK7n3A0tenclOv0scQ+QZnnKTBsibjtAnek38dbx81nUJSvRpBs
yzph2L7phpdlWLOPgioRyoUv98FiOsYZLSXVT3biZB42BcTDnNIGW8hy7C6TrC+X
r/MwvKB2xUYW4fPYBqWIlSeFCOakKijHFyjvbcQocLNORUJOE+95mb2t6H4r1IjE
X0kNaQov4jh/uUEeSD0ciT+3gxVhlpAul2QxN0nmPpuUYFv/UtNKQoXyDoTb9AZk
ok+vt037ChA1+9qGODpqAVIKIDEnck8lOIlflfVkvi7JSxJBGTmxuox1Pzxgo3Lz
Oh3ymUqltzoiBtlhJLv6rlg3umxD8Cma6HXgvQFzu12bT5j2LhlTneRNQDWOAtak
GKkY5KRPmD1VI9koEC94a6+2zY8q5IpJbmUDZlj4aOVXnrf8N09A8m2Gg0cijQBm
dcoaxSvtM1rjSroNztu4dirtVv0YnHkt9jZfUlrUwogv+AcZFlvLpWBhDGp3DvCM
mJMSJb9vQLr7SDR782g07HpM9IwVKeEf2R2OoUK1bO1vIoxnFrgItIuIGNILCBEU
ZUwRbYbOIP40uuBP/NjYQyNJruT63nUZYSoiMk/wQC167n0WEJOACia4bdME9hPE
tdMms3K9GE4lMgwRXtNsL9oVsXGOKyJovu1C63CANmSxsgd+YfpjT//M4EKoavIb
skiQnRE8+ayFY1ujZPDPwtGTN1Q6NfX/cEoyuxJiqhvT4HXLLi5DhvzXrvXW17eb
bQ6WlUkVUBnhEBn3MIVXhXmA/NXtA4Ab90dCWRtYeBpVEn0XPKErjCaOR5i8QKzB
XVWndyYYjzae5XODFV3TcoMki6N8W9vhD53HwezRBqPNUkP6Batw2rXM2YtK9U+C
vgtm38Ub/xOjnKax91BfMnkNOuutJag6+f7d0sbQj2a4SBXI28EqU3BiAoaHV/wA
09yWhNwUxwep+jRiUm5dQ2cUD0T8nSBrP3XvqWwn8nMLTmFmZrshrhOnje6OHqxy
bitRoYFvza+HbHwhxj4Sozo0ZoP/luwxrAgN3NMt6XGf9tLiSR/3ZZt/5RbV8ZgH
6VG5fIm4bSv2UbmO/cnQVGuQlkSnlhTv+DW4uhCH4lgxXgZUSfbXAuxqIkT3MMqp
I9dhEMS/cK7vidlWbodHwFmkRXDIOGSnqW1MLErOPC+oHV2VxleGzUhC8UnFvHzo
9kRG3p8UrdU4yxMGJfII6XRp4/IQXb/Emd59ukqwoH0bQQyr8AML7BiWPf20A0vw
IRPNhsoJwspYlxdR66hxVoGpdBHOLaOY2O7nuoH1vPum38aCsBV0CX0IUGRKXbsL
LCKQk0b2ta4U5G4Xu6wpXD/ov9Weg2aAwl9e3pD3tY5urHRb3IdOxOz5gdTpHMeB
NVTSJ5dwjV2q+OXAwQ/ibtZmsvL6BWK879QTJYMGiP0saXOlWtr1GBswaN0ZhLqc
R0gnPVFptZNoJQGT5UdZMAftf2s3U149xB/zg+4eNkK5kdyE0MxD9LpmZDSN2iiT
xdvsyguIkDZbCVN5Ei/6gFVZVZTJ/l17VfpX+m/C69OKQQgGIZDzuU3XZH2koJTN
C2gSs7zRd/jA7mwonqSXSPthhKk8J+qeLYdqf2sv9SRuVCnFlCq/1lhPw/rpBPi4
noYdbctxrfd62RvDbW/Iv0roLzjzHw1RMIXqZhWPeq0+mKfpsBBcRMHZhVnBRhTP
sZ1A6ne7rNGkJJX1MEx3nfqK7oLbi7HayPWWlDGgG6G9Kna9ECrhzvbmxFwAkr+R
a9frPQNi6oo6NmKPgF1eijRjE5FAfBKIlTR8mSCg8ccEummnPV1Kl0g1iBPGChsM
TVCQ5Bk61b/80HcsEeZ7qV++jaGPNWYwZU5dFip75tiX/MoKxBWxzVuP5LHFLWvm
jqG92KnW4Qpm+ZYPlo70tZtnKyuVRv5F7ZGlxD5vx5mM6T1JReTgKDH/cYX53U3t
v9Fi5zGcUslw2uPq1Xh/09K9sxQTEQCQ1bGnYK8yL+ejDCRr889Gu5beqA1zyVZB
hfHZqN34viqA+cDq/bKEOzHIxwQd2cflWTQxcVAepePgYlcpBGytS6/NhbjjV/+d
Mh8TrX5pLRJwn3l/i02psh2DT+s/+tYZcCjr0vM146T0aZVCnYDixizvBf5iXtQs
dOrHt1ssyfJqYDfdccQ9iv194yRV+NmWs51XWm2eBpftktxJAY8sly+o2PqCBEe3
n44grN8qJBXTmc85g/3l32uuK4r8C5vefOaupqAiR6YUBPyCd902zAxEv7OICWU8
cEzIU/QxnxOPAFoj8Ek+P34DaJsIPP8dPUPOdyKtecYELHtMP/5PkttNBEWNM48l
udcdLWgj6F4DXReZT99e/UJYPWHvjEbTeJweJQ7MM6ydf5b9NIFtq64O7CWdEet8
MgFhG9Rwew/nkYGVUkf1mG3XA22agc8SoxdBcisyJtAzQj7TnaySDlUggCPpRRvb
TVVx6v8pOnWTAa3NmTn3AY8/A4bIW+pCfE8AxjgjCG6b8novdBqVQmFgEOkNDmL5
46+bVuGXLhpmdWGcjxLTuGJIjDPMM2iJB1rglI3KlAvgwoRSdO3/ckD2dj62ejls
vLTMUho3Cf1mr9pA9oK/72NkmdCQb6/04rjwVXZlOx/FQo8T74zYeqp3S2yhQmdw
BDkTn81k9MKwZqZMjVwJ+YdknMy48vbtHqUmxxicEY9VUeKyr2A4RHhiBiQ9pdvt
yucP80IzUANh+KmhJV0SJPr3hV6hjbsSYCiVOFeQjovRQQ04Qzhb8X//xpEibzWo
xCrMYn3rcZh7o2GSd0NjcSzw9auhfel5/el33LMt3nMvvWjdpLTInqgWy6uSt1Z+
x19saDfmFclwSxzVykNrdg0xlzuNhxqfB+SIsgzgFelmqq7wHfpcnZjh6aNkYtr/
3yVFNL6bQNjhVvxhQU3vbeM2F3hKvBd6MgMyGl0nnLMesd6YRUz6X8jTZt4aaJz3
sYK4aTVff8o8btDLzfs/sp4Apc+azfOMlUQmWk6K6NKmKj0gVWonJ9usHN9ZjB5B
7Dyb2xVcW8h8oUCzw+kOwI/22kS1VlnDbNqduaxhGNThg9fgzU341Hwv+NchXq8m
QFZwa2R9pZYx4Y7ChTW+4sbddt786BUYQYKVqMZHg3Mzs3R7HW0bfOV8kOA2Q0uT
oPCA4IsHTSXGv14QeALJIlDtthgGIpxUThbXuC6LwaiYRBXJPDzxkET/y96kCrsp
QCprdDqKKqYDjb3fyJRJ8tLdu6bJQFDBt7e8ogaSwcEjEZZGnkop7jhwjZ3F9RGU
QQxb4D7KkMlTmMfvPgOqCd1k+mSLsn48JJPPJaX1w+HIA6dP5F9vrYNWFksD+VFV
z77/oFmA3+Yosgqb+FkfrMjvSqwVIaiQgV5lCHf3FrWmnp59jmotL+FYbVJEOAtM
nI3h1QRpEwn3ogDQVTtSSVJOqJgXEa1Hv1mSIxzxp8/F4YRkMJp5WsHAtBuOMR0E
6nqKgl9tlYN9Qld1cYXYWMPC+5AyUswJWMxk3jT3xfetciMm3yAOHWD53xCyLyei
dsKROjSr8dHdwsNFLiwmdfx5lAc0eihOHNxFplwM4m9HVCyY49sudz3LuEdSXd+K
fy9ySOc3QlbdUtgyVlr1c94I5P/92yW06CUb79rqWqRRVBXpbYyf7vEUZyIwzBpH
cfz95WXUGPM4eH2Ps2EDC/LB+GjPbgN7b6hBJzHWYCC/IVLW1AJzDpeXDm06wCVe
lgX9jCUIG01GdyoO+NHrIHL5S1lNdLZ51L+f52UzU4wkPAAyRgxN+5MFGdR7bkcg
FYuZxh1YkKh4f7u821sLUnnKMhhzadSHKO1e5ChDfZrW3oNYpwkJODA17AN4xtnB
roBBQN/z3eteXmlpxPiKaPIMEYw6TSWCeE8YI6km3gfYBRz1r6mh3qb0su9jva8D
FHz7H1sUGi9gigGZ3g7e8VWKKf45IrUH0NTHsuwSfblGF0PA58tEvbjjd0nQNiqG
3jNhIH6X2OCyzWwfmZpXOrOREqefLlYlqP4SOR1BaCkZXb9671ORLYhSnTj/c7fc
/52yNDz1/QYlIzziUrbDt8y8iJ1QBGLQ2LeWAwuVTw2RKUtlYTIGhL9J11o/l1Fz
aaceZbDEh3c6Ks9ErEtZ2j5nWx4mQVdtBm4K2V9xev+yAveddCvuSedT86vyffrL
TGEmFjubhl3tZ+DuXY7GSVdVrpD1sc8JEe8uW3yUHjXJYmKDpDuQC1vwcoXW/Dex
D1exu5eIDjRcfMQHv7r5btW/oyvTfZ13LQayK1dmzcVxa8ZEMp5EpfKek+Gy+bPW
mj58sLchc3+vV0CBtya4nNyIk2iapFrguekRzbhWigP1TqSFt9iOBcru9oZQgPIk
I7suNNzfbEEkO0hw4PzDADmQPVxAfFWv/T2w5fTdVBNOOgUwidzp8DB4xaYEeMOd
DNUQ8No0bnjBGw3fd5Bfo8criJvJZ3VpdrSoNOwhNUVjYNUsWL2PvIi6K3QIveIL
JkjYKuh07jMXYcp/hQgtMe+cLM+R1A1OMwAKk7DMrLoWKFeRdTiztTCtS0+y6GL1
vW7CYKWg7NoI5CNuzgm/lfinOb5W2HBhKeoxcJR/BvFZ33ZIqHDQSKPgClH2ULzr
c5tMGcU/HUGjqJYWhibTc9Nms4f6FUWok8Vb0rbU+klh16uMGXHTFDyReQ1dtlk9
zJ9bV4hd6hwUSYqf8iBGHDmJvyoKsKklWCncWwTwC1ujA9KW8LcHo/CL8uSVeSkx
9gPfPh8Zyo6psceOmaQ2wgGO5HMbnqzIV95Se7gdGrf/TaB4w7hyohb67rOHVkBf
Dsq/HQxoLjmXT67PQNhqoJVUgUTDqCxVGrZhJJQmaW6YfGeLfFlxrrrQ0VJ2mkJ/
Ro6spH1zMmXVUrFN1e78gsL/43Zg3BnhcxYEilM29KtgZdXrNyHoNNfD3V6YIDE2
6kCgWy2/clkq/MbftYwsP6EIle+QGt0MQETxPVD4wzirtQKzgYOxtHZiUKPPemLt
K8lTdZNpsLYsGXqQ35dglzIXxROAaraOL7cKaB2ZZFbS87RQPGmAFvamNbhkVUJk
iI3ztyNQP9LMizHWckINTiAFvfFUcp4CcMS2Co75GIcpgYF3lAwLTk9MjI0OBnkX
IZEWuxsbCEgT5fHd2a+CayO7HgEJ2qNACnIfIulKmTI3yTwNkKSlS5F4/pMszsAP
TQeTK/pA4aXmG2FkPjyFnj9aq1r7B2TG3mdAPAoDz+8GsZSLoJzNlscXeg92NGGC
9zB7tEnisYkTAOZAR4Jx05WuK0GSa/ez5sLjryRYVC5RqklhhRovGFspfI+YAiXK
FhHWJvD7OSCEa1DKfA5JDnxNPxxLuZhpOkof0Y37rLlYzSrNdLAysbcGh7J48g8G
Xc3E/F5ddXsH6qMMtVf2VfFa3rUn99/4q/7TeR2ewYHiTgBa3NTPDhEWXD3ZA/Kd
1ihKhhM1Z78F64nX6efrZ8CYSQqRt7rwve/oXYpRUj9pcx4vPPZ+DMxQvWlO5Slx
A3ysoTQfyzsGSLEGHeBfLSD71U6uFO9oJmmmj1bw2RiDKExpde8NTrvjl4TmH+7H
/pBebMxfpNH2LZsN0OwLLZKHktLshkSFMz6FUTtMnAc6ddgqAddblG496Mh1Iuvm
vXlO0HX/s+C0PuiZ2lnYd/+5jQbm3vQf1WvEysB0gQm2kCBFXnRL93qcwD90L8m2
8ORPnl3Ngz++11ZHJshPUZ+z2HA1ueKpMCTDsdN8ukeK5+VAXFCtGXgRKtcz+K7Y
imG4312sSyUfnD9NmExsGTgCzDTl9BZqVBPL4AqLLkz2aawGrJ8Qblm+HpOKoJik
6jic8RVMr+3BhyF8qc7Tilc3vlRRR6viTfFRKPe5OXPvVD8NrRhXGktoGkv9H7s+
zvwSVnf1sLwLmYPSMAh7xM2kmHdBLwF0AuFZeugs3vbDh3s1gdVkO6dNtrkPvIhx
uJqrwpTO+DHV9V2bvcjCjDD2AzWPY8grB7BrBMOpo5+VI1+gZTG/I8TsCHhL1e7Y
SStskQkaMPPPzZb3yDhvShJQJgz/JsBi5/cb3gk07jHY5z1meu/5adlsQAOGnB/B
gvXh/SzsZ9a7VhJzfxulHJsSNJKrMvYEXo74e/lJeuvt0/4NJe/SGXFhJPrhdPZ3
Q+vqCHyXj4U4tayErhL5xZwRpz4nT23DADUmngw9RzuLofI1lLQKQ4QANnAvoUoq
OutDG2YBbtbFgndrXCjK7Azk2S/QX4+nWdymwJsTqjrgDSnmNuHOQjf9CTPjzVHI
Tn7W3VBwmGQbIdu1EcSMF1a1BaVLJpk1xtbgY/yQTYZJQkR0I2EekIzKU8j+XM8d
rnfHKuJAbVQOb5OppNl/2S+U6I+4yQRomdIyr9YDMe4yUWhSXdv/YBUly/E1bGgm
QAL4a6wRKiuDEuyvyfuEXX0fZalnbCkLnnBbl0lj2xhjAdRosqZgDHqSUtfQdNga
Y2fzal2mXCkd6fQ8gxAis/uoD902Faiq9h8cunDpQuHUG7XZvXgitfJWQmNvR4F7
xz7aF/xw9beJTGyrFygjcQLukZLK7h04G1SomJ3kJ70MAIsu4D90nZ2buBlRsj7r
l70qmWS9UbCaAkALo0WRx4hWga7WCtbkpWrKmkL5WEdrvKcZg59qpSVxQpaGuhuY
V/tWlg1wj0K2shrzn63f5SttICzxJMQ4P5sL7mn5RNt9KJ/2lHKYCZN8XNsHzlC0
FTOcIyBgtHfbJEP+qYLUnjW22pCMUFX6ru9aB/x3+aMxzXKPdTDidBgzLzT+YeUh
lx62fZxOHwXbzwuMKOFbhkwpvQiNEMcyOEI6Mcfx7D5XMre/mIv/lNp7oBXk4YKw
cKJR+LCRKbzonuGWRDgEpkcZSLJhikrPDAf88IjPdo0ehPwkJnW5GXCrI/TewQmS
lhOjQD6dPlaTkkyBPq0xbJuKGjPkxDdZ8DNWRhoxxcHEZdi4GfepX203egfJ1xdg
WtiduuZ5TwN797+JdI2+OIPrVTNz05LKaC32SBoxP5lwWUxLjj89qnnDfVtSmUTO
AG7hiFSU0i8hIcKm4xvBMdua9MhdaFpbQwOl8tqqnSP4dD8jl6zL1BZHiAG96Cxt
tS0O1u1gxQAUdDOIhboWGujOnYiFVIFQ/YfyeYCo4k8WDKjlyeuqeNPLjG5nNLw9
mNtK1dVGOC9gomgamdomub2FypMI/cm+H685VVjfotmvkthGBZrks0O3zmlVt3t9
24ntOI2DfX75wdSTBVpU3FWUUKOEBhMlWpPbo1rX/S6IDelYCnlImgV2UrlfQU7I
AH7bnP4U3xLkOuoYxmqVfyOQcHLY/ay0557qF5A4or6ikqkiwGG+aP6rRsiP1jAf
ibvJ3ZaYpfeB5NHXwtvaMabk6PsiSsmrGqTqPSBmnIQvyYToVWhKbYIPZoQgA22k
tVyo2+jEMJbK0E4qG6WG4ajyWBQ+W57lUYpboDLwnmuVM4OOTZ1fZY7CKbwyfZoo
r9wdLi3DxKYNkznZ0PegS79pTUaISoTEITwVwLnjc/3s+Od7WQO4dP+60cjB3YsC
eDc9RK5NIDe+kSVRNMGLmfne3MJFT744NjTNfz8+k8cbxrkch9UZS/krEZy5mIez
Nmiqk0ErbrK2DH0fnpcL2jLEvUSGykXtAiQasQO7uM627yZ1YCd10AxLCcbLvKMz
aoY0lcGOw5/VWonp5q2IzdpeKC93U/FnO/2aeTpO73TiWTj6cWo8sEMMESr/noei
Zujno8zFZh7DH4JXbUzPIYr0AghXl6ASW8eGO4dWEsj65OErhUK4dUa4Xh9VzNSm
1jt5l5jW+t9KRH/OP8B9J2+y84LXFmsuadJJzxU/chBI14eVnNbcsQCIp3Niv6Ly
aobTELiF2lK7QYJzkWr/a9ZX+eXaK0rAjHAhORF05fUpOoKBKIwFCYIDMxUEdm+2
X4DK8p/KukKOaaYeLE/ejwcEPuC56/ebgXh7E00hbiwxpE/3r6+KZTUanMmiKXXE
+WiDGmbLAmSq5nuXR7LgFNifvWW/GIJqxcNSLG4nyTlsD+vNj2kEqXMbO9BSVz5/
GUJxwBVLN0kwcGsSWHwtjd8jDs32ey3KWP21xpq05tkFC2WRo6ZUgcC5rCYrh1AD
7ipyrNfLogjutIvTTEYZhs/QHW4BFhOVTM/HrYsMmi/T/OWaQjThTWczNO4czn5Q
M0wAjqEP5bno7uR6xPg8UTT/BlQNyLOpJsfhlcIFJxTppb++aasLTZLVcoyXD0jH
bBgauuCxU7X9aUUy7qbH8CfJCztVwNbX2gj/T1d+ceWVK6lfwooQrFCinJ4ekQjc
vYGXVV5SU6Iq3Xfbw1dfAxUVQcedlMG+UetUqXKQ4KqK9WHzfBEs12V8jINo8M27
Yt3KqZ4188sU75pAEH1xkgs4Gw4FX+ygyXb5PhQ26L6U9Q3DkzuozWIkPVZ6Ag3r
bOdheA8ERhlBUx1BcSKg3u4ffnXsgv3bKad6dLezV9EXXZX1/czpZ19y785ht159
CliUsiHGvBVZvNUhawA1KL1Kbi7OaJAVZz25XesiflCg3VbnooMJfUKfIIlCsOoG
i5+NL++EieGi5rl06j48KF3jOD8JKYSKhnsp1bCQw00JuyGepDOL/GiIgp9Ykn0C
67t7k65DU9xJTtyL4mFtAgGvnxchw7eO1+l6q78yQOBZLZPQ50Dx+/+j8sKx76h0
vy04LJA1uGzAnmwn5dVfAoEXHN0VR3+j+LqZUkJnDfBWPYu4sgWD4qDMH9FeF6TT
zjTHFKAfXplqbGPOgh0mgB4pPoJqD1pINBiOPaqknkcDj2AMb2wdc0loqjaABU+R
Fjdwezia7nWAU7MwTxxl7nHAohoBiyqZk0dP2sQ78uAvULuKUaFdZGPAlRo5Wj56
pW1dYrbgZwus6pmGWBjWDmLe8W6iuz5vonI6yb0Snqbn6AWGr7UKNtrNoRTtYQir
IATjVrArbYs7ku1sHq6qCJIabf8SS9YOWJHa+Tsb2SkM25o7VZMOLBJ24tUYKFDH
a/u+L50r3/CXh3qU9Qz4yaCq6SO5rtQzl0lN++3EjaG1tWNm/FiJLuqxhcTi/Cc1
mQlrqrH/CkuaPcG+NmpzKjhvBmmh4Zy6Thy/H3Yf9LvCcTV4hK219Qlr9BoMoiHD
r63KzuaCpl/aVouJtxItK90hSYFEjGTVgnrlgrbSqLgk8cYV/aZ2HtrRvntuY9t+
gvyemQ5p/nhKId+jgTcMDLcZwZh1hloKaccDd1h/op8mY8M5JcqEKB1Kx6Tb/U9F
b5LKnrBxxMHGAvmViplR5mHtHWv/ou0egCBf3kVFBMkQH8FHgkdtM69zoB7s5sSL
plGi42QK77rQWXts3ZvA2Xd8wgT6pk1mNMliYrFydB7g4ohehjBU2k8gQeUtJzhs
Rv5Op5pTmdkowmnfF6hBOtXCUsa7Afo3a2zkENlJwoBcc7/1RcBMiaJE8CapQNh5
thzUrGn3Enl9e1pjSxd9fBaPf8eHNz+KE1fbYkhEB/snPBbHo316cnhoeerawI+N
ME2FheZ0FaUZHEkEG93d5mPgVSiPKq+PUdQo8OaQyeWxsEjIYMgPJB99Q/082/xL
bYuEOTEwrkFYlot/8iGe+Hvu1m7oF7a62/FyTK5+JiPy4lddMKtdLMDaOGxBO7p7
axnz8e+tt/mqJRHVnA/upj/9t5o3WSkYgQnSBT49pwQPvNELz+SgKg2PFVJpiX/F
u4X2one3pLKbnJGDh6bS+ePuQloZBOk8YZkqQuqJ0ROA/UErf2K6Up9lVlRBeitU
SDQg+ch7hl+grjIv0WdsdbbkIyKhU0TFyPozhgbouZ41RzAQS0oVmUB654pIh0g0
Kdi4kaNEXuGs1uIuEO+RT1hbKMFTe/Siljd7UbLBmpJqF6LChWBu28qIwEEbWRp3
AcRGLylx7hqY7pL8k2Jwu3UeLNAqwJayA28DWRDYn3KqP3Nuc8kzeJ7FlDAO8Gky
E9Exw7F5znHmRxraK9CskH2yBCQdgkAvWlSveN0z5oKG+D8ru/BsIosx3Pinpm4P
JD6DLsM2mluaZMTGDnC5sxgSw20eiUxIgCPIOpJdTnYpx1j/ZQxxKu/yqHnGdkYL
gqvJq6jGQAZFTSyh9HhAvmazrp7rENifB28gb+cT2aFfXms/L30+uhf8dCWseTQo
ndyScvMhtTPeFyzJ+pPiJo462KyF70A1R3Hj/J68r4puhzePglYFWT7AHWdKZFHq
gATVFuMfnPdxbEchWOA2Lq0nF3gZpws+Yt/BLa/Y6v6FnO/VzKjlpL3MHhNydVB8
QrtFyp1nkT1p+DMDrAcL+esCwvseXUsWDuONtwuLDGjwtuBxPldtHXOlYxF6X23Z
+AvL+w9fn80FxFMTYD8Lqcw/efQyiCK+ANYK8IOGp8S7OmTY4FIWyeYEhIigmGCq
6IXmVE5Fq+StJLOZ7j6KkhIddnKh0DBSSC4RUEwCVkgLfOIInv/UkusRUj5cPZYn
QG8XYqIUIuhfyxUzA8gPzZ4sG9S775GbM6W8ZhNlRXlCutHf147J1u5uMAUa6cX0
IKJL9Z2lh/iLyMjuCCooUdJRDYca4qf8SmIvnJe+eehmJRclrE4DAbRuzBWLFr/R
Is4GxpXnm9k2WT6yE7+6AR0i0lpItqnNFZKM/FTp5DVxZY+GcVWFL9voZMq/xgtr
yPvwDk8FiiMc8nlaRNveOZm5UYrZjga9U/zRgn2M3uvE707cGAfrAWxsqksuvnPP
lgras7/TQWzR9hhCSFN7vW7zyiCQsb673NThN7AGznSuE2Kv8RPQUPGyRr0UqdFF
0TLcAreTep8ZTFVFL+XptuNy2ogZR0W2+zh+NuGwFHAIJRaJQMzHqqxfqlL1qPao
kSZuk0JnKLuHgd7kMCO0+fFG25AECViHCl6M/tlG8l4xnVfFTP9nysY3NRJtVEg4
9gUDU1nr3ApO9vTRUBcG8OBz0i98w1szg9UUtw2mUqQAcgUtvLR1/szEbYhm3/Ys
a7XdqKbm9f92j3Rfaq4yze00QJ4FRF0WFoj1/gqd2wUe0Ktbnp2TVv2GNsry5wc5
00DR/r6nUZl2yN7Heb4L1f1U/ZnVAD4Ilmp+4NnO9sKV0xpgF9P1EuMMQoxQwYQ9
xxvPzfX3Z9GSAwoBbuaUb8+XqhezielsPwSmlUM/UEDHcLxgh15Q2PiOra4bSApW
zCk+Y4b3oh0ef0NAojH/A3temGHgNS6S2lk/GWIHxlq+Jkw5DKKDbIRP5GojwedA
COyPsco4WLQsmOos6XM1zteKCfspuJ/yi4yDcodqrqJaQqetPI/IJPRsUtwFkfOi
9UWpShLMkB6df2eoT5gtFgQ49B1iBAoZ3QHBU2tPhhAuj41TD8qMJnUD000TlOKa
tYVjISBZ07yYp1JJ54XX70I+CUudMGwvvfAsCMDpi2Q9bPSVV8POx3t4DRjfOQjh
75laOPNHW/t5D0ke46RvfpspDLiL5jBsiUGw5lO80ZXS2t0fooFv1RgcG6KsNTYT
WJrku6MXsaN5GqnhMvW9HlYCvE7EfcvqPLIGndy2Mzn8HvaIsPPhkzzEDV5oEEgK
xoYvx+6h3rt2RZChD6v7twjuWmc68giCdTlt7iUJr+BV2U3ejuDf7QIolhxP42ol
IYpAUbVxLsPRhWFOIqETe7HuWAQB56Pwz7Jl5Xnhwcf++9LEtQnUaopSn+BteZxD
K+lGMWhTKCO0kA+iA6ui2ai+jrkLfqSFfvbMX9QKmvC6YevaXgXIxlsB2SJhb0BH
mdBMKBwO2gM+2EG6lsarSdorWf4AzdkBrfPPFRkLCeeU8qlTy/do5ezuNx1mlR7a
K8PZd6jnYVBpb8IwGOVQNaaisdp3YkLS7Ikk0/JSArmPV5vTZyv/Bb3vx2s8zlzh
hL2Bvn9VEHjbaYC0NW9kguQsZB/6t6pPWGCNP48tDIw0AOxmlunhAPB3Sl+3yGmV
OEU438HqSmf1uky1jr/MPvQG76/JolbcxEMWaEXMdTmbg2s9/r0/DfiTAKHoKQ/7
XlIrnxR+gPitRcJvQMEjUHWN7UvUkKg3xhCDWmlSaZjfxQWuh/6T71jUkoMatocm
jt7Iinn47Sl3lrs+6JCdT1NR4d/HnGGlw/lzysrrWDh+JMuyByiTn6OXE6XVp0SJ
kWGxdAYgr2/Zs2PRE0lM02SCj9g3MtlsZO7hDAYFtUe1HCbsgs0x7rKnikFOzagh
+wAuFK3uSW2Esvm5HeD5kchJchXL92eYnTTy3nZCqCRz9TOb23F5lklxXif/BFr6
9BL8cpR/0STPLR2/db69vO5aIAdnIMeM2atyW9sEoVvksjN1Juy4ofEmgYgbtn8n
QtTs0psXeGOhv2w9+ULp6YaBu/kuTbwx9ncRVy3tREr2pVZYwbvm3h0IUvGeRMoo
7yuLCuLYR51sXLfefgpuH3vOBvw40fPWXBJ+WsjAbGimnOy+SDrKCxP8jLPLLr7i
MIfkWKdv9nK1kRtbvHbebwKP4YY5IPSLsyScvzDT/JeWaqF1FrM0UeKQNVg3YLyN
Mzrsg2n2rd3QJGchJfhzKbWRMOVGOb5O3zmwzPNSf1LEyhBHhULAdiuLZY7kUyeD
KLcdeZSgxhaQD9mCXt6iNrGatPksvWRGoOHbrW+MJtALdoFkOgXizGjYR+X74skI
7EK2uTEs5lb6v93eHdfWd5sYerxNd8carv+jnPlo9ctNN+YbXV7UJOy4SAvsPkt/
EMhDX+Zneyv4z6K0scu3C/9m+9TEsU/nJs8Deu36W7l7ltI8Tb+Jz5PaPL9JsoMU
vu112ZmJGtaSliSARKYaUeuRtqt3s48GBEyjwqQrbfML6nMgQV5ipzGmVwmSlgPg
9G7+60Km4qjWSzt3u0vQq/Q1brBqv7fdMXhlKwToy3/mApvoKZLZVU3Hm9B2QyGV
vlYMwjUfyuyE+sKdMbZaU2gA2BJEuP0Tespki0RRhgwOY9jNVCA7aukRFGrpYqXT
MolfQ+vYCELTr533f2OcgNy5gJKIdstFoOZPCjXufnD6dEUl0Sedj+HnKJbDywPZ
2banaPcVD0D8Taxstx0/f7kYvS6H/9K0UbP/BqqJm4c0aZMvgzlDQUlYrfHMhARs
XHtIv7Sg9x8LF3wpGAAWllrexaSCg3X73HKRbTz3UOFeJrcIa9WIRBS6/LxcgCIN
zn2wkhp83aoOIz8ZXpDxDaT0BDNooTDx64fbgqnCyry8xn9U4NFMB14t92i3CYSy
GmywHi6GJzvMTaSwocSLTAO3QoUTftXIUtOKXeviCVOAM4CElTVx0DwivJmcCcVb
Ga+PM8qPPhXPzdO6FbLhf7Dscf0VL1mCngfRgQjLUoK441UeFkQEp0q7+50q5JIS
IxnlD2o4Rmxe/A8BZJDZhegVEsVHKmCxX+5CqpFCZu7GswgnyQfDZilXtHhJm033
2uz4JENGPSQGeRdCe/VcR2D7G77EBH6VlZ0fEDK6g3ncIwYVegIE0eEbWC6kNXfG
cyRZGR5qRXMgbtaqOosgL2Vy345EfGieNb6EF8nv0uEZTPCp+5R1HgksakMp6eOe
zyea1rI9ZRI4v1pdcrcZmEVE9/R4cb7TETgA7/JcdXfSLwcAVpqu6T80kTmUULab
P4CGU7vIQCCSQGTMBJ6PfQ8FHg9Jp1EI20lyZZX1fXJXe0c+PPaUpmm3whOYXfsp
H+/B9y8Qp3d6Y4bUtzGHgG/MblE8ZoBf7Tpl1b7ac519UgtD7v0qCc5jm1W7qFDo
QW7mukeTVpgIu7mPStgEJaDJo364NF5GUNx+GDSwp1cdJYvtr21IIYB/iv2mtIRN
z+ZD+vC2SlmNvTOH78PIBj5+rZsaYgIMYKsJGB3iLksk9JlfUJPiLK7XZopsnfbE
4Nj3XESdO79R7amfG299kkOLuZJTMoiXGZd7oO7+spVlQQz184nfX6Ldiekv04by
ta80AH7jTDcODyAju36rPg3NrUwPWh2PdWbt3DfweMUzqTF6edh8CgDLz2kP+pjI
2Y/hoBdihDFn3Yvblq9OWrY8XXYGLoXpAcx0jGqw4+yk1crDbx795jYe94R8eJBo
MjSwADgOFsAmoOV2stTLWxuMGzmRwVNjRoFb2O3H/tutxxsdawHUXSKpwS3i/Kb2
Ig0pLKuBFPWTSktD0D/UdDhgMs4OfT+XYdWQCkqRPV2JyniPaoD+PkceUpItdy15
oXBlK2zBzDdyso9dYGa8nI00mFESjpPMe5LaBMYAO8czi0oupC020jVb76auLTvY
hJUpi/pO5YpL4ZFC0+S3AIg7HXu0wbH7466/ijydOI19xf2AAUydO3yL47ThkSaU
CEtMIuuqgbJb5g/ZVPzZO8VRH31QPSyuca7YJrj+JskWAkgr1Hh+Wk3fhGNNJFb6
WDdse/Q+rzecm3CYW1ZQAfWQD/k28fuGNCBzpVmJR/i3apktd+p5YPultFiUGVr2
njFRg7PWMpdS+UFWSdv1ROqHjrgvH+Epv18ZBMYnpm7K0hrWR8wjCxhZZRem64p3
6r1y1TquwvoYIEHFaxhMLpupkOBr9caPFbiUf4ifdXwaJ7Me1ibaX37a4JqR7crz
Gp6iZ/DVS8W/ijptT1bF3dcfR+vAC3vPJs5uGovyga8m5Fg9UA2wKkqIZB5Vt4ij
+aJoQE3ekMBlLCmbhlBPS5dyXQ8VUaAyUN4T5/92hHlthfccPFBOVNK8FAlEr6WR
C9K+G8p8mV/772H+O8LHRVOgloDpZVa1z0jYYVNT6UHUy9tcZReSFOacJ0ia3qsx
b6LGjsD5i51xHk+k7IUyJg/HW7a9KSwYdzil6jJ0T69HONFghdDbPIXIuTOfVCUk
tb4KTwVt0Fq8R3SuVn4FG8Lv2OUf8hlbTuofpd4xnC84EkeYFtFn0NTj0PmIEOZe
6oKZT42LHAxzd2s28DzygNsW9iS5EDjfLnPSx9D9Qpug8nAt5GbZEvOoatUl3lXd
xWzm2oCbEK8HVfC135SQDbvIHh1eRVeRDcqjQr+AMM5UKSPmso5qOvznVcGo4qbt
mZrJnS+Ea0jzGtic5DtCf61dKSo63TAH0NUPwOzRGr1v+aaBYXU2egwDuqf5JqOI
io9Y+wS3hUqd4M7/Vats7/FXdaQfZ7FLmsbR6r/Jc+6isoWh+x3oFfywNg8UPrks
eSQiMq6g96by96KvH+ZP0oORsa4EyWcxwB+Fpd7pTLgPvgjpkt/E+3DZHHtE3XtS
QAj3WI8mM78Zbj41JwEH7gsgIpbXcSjVExdFMNy4wyaVT53EsxvBeYh+U/YZfOi9
yUnp7XKQPb0EIT76jSXaoe5el3RPuMcUXvBkB6tMsVUeUiFePFA4Xo5JLXgyHzfM
ANneOZcDZFAGmaBR03JfKg/y8Yx6cUMJUdl8xIdbf8bt9sDJkV3PKWZGAxUxaCmY
w5yiWU4AQLxeC4mLjKc1F8PlYz8Mr+a6dxwrz2WIRFML3GJOrLEsPjwGx7n4Trxv
A/Sg/inrVx+pAEmFoPkO0JMUdhsS1XfgnTn1WpRiUUNho1lV+bQLRoBmpKsAj1d0
Jzw0GhiNfM11fPrgaSi9m7dXXIbX/dO4TseTj6zjeZOv0pEsbTIinv4U6pOLI7nn
gyFH8+PZLxUbbvWLE7k2mOD6CnTfOVMqE6QEkXPhDwjTs/DTExyuKo4J+vKCjw0u
xlhlqMueGpgRcdewNdXvYhM0Y0HR9lGk+4j+a+x8Itcqa6dAHvpjJKN/lLJA8PVO
G5uiO2cTS6ZumIMQq64x8qllghLolLPQiZN9kJGmRpG8tDlHktqyTexWzkmkFbC1
9V2DU3ianfqcMqVySQTTrm6/iV6/lyx9NdpAWH/HdbJsvqy7+kxNrJhfmSmmA863
z5GuuhBHz/h2P/nCIh64/itm9j0hdmDkuPPEWFr9uqNfBocnXB5es1VNiwDCzI1g
cnj0fEjQDh/oPeGRG+l+fWIQwbAUorE+lL3do+8NCHAEKK3bm/SPN0AOePsXsJnT
ntDU/b8ZeDsxDwFw3yNIBAJl2xEIsGuJCSfS3fjsJVWhwcZNHgiiVVjPG9rZpcEs
aNeQK9yG9J02Y1D4KIojWWbJrwobxSIICbM7cTecFCsjmT742FKt1VABvxmFpkZE
hgVex/Jz6obaPeBCmsyVEgtG2kr1r9pK5yA5flmLHsFFvd6ImWqPyNCLQNWr4aSC
J8LDHoA2DNUqk4YLN5TSJ9RFhqOnij3h0YWMsx/l5OGl6fqdVS2hNVxsdojOOGxm
Vz6BzxNxI7HFzYsdruslHDZ951SfzZogWcVB7mZxbJwo9hINJUzfGI13tOr9Nx5/
x/WSc0Sbqb2pDmM8eoqayneZKrsGJB7wasAbC4njhXHjL9BmI+/Vle2PsxnmQNjy
A8ViffR4tcYj4OkMNODP86yVTG6bxrg6lBU5ckIYPm40vOieBWehZCxzzPNsKTdS
d9vxgVFMqR0CbRxg2DMAxwfypcib+O/4DJU3a4tvqk5kt+E5aXgUbsSrkXcX388D
4aR2BDyha9hmlQ/yzCF79n0LduOcekWBEf8nE+SFUFXBBXEz5HpmOlwRtL8uCpAW
TA5Q1WMJWHnPXSe92o6i+okOtUVKi/tH8MQbBHuqEANfT0p/sfZVfivDyFrrVGG/
CBB8jLKdxrZDJdvnQ4BrgzweajC0zUB+dQ9/yAg/kDlkbMm+s5N3AlGn0VSMLps9
12yAtV/MvwapMSONFyKgQIDgUgk8Jb/oPMUTfNjKr7UQr45RrO6ZEnH7BaJPIbPK
giXkoDMWlOM+re+706EtkVeuAozrNXeePlC20qgThQ9xRnhlW1WZf1UXYX5SNQYe
zL6aQDUiNw/03V+jPPo11hcwog2X23X7mrTZUrcauJrW31NWnDkZdmTpAf/38Sqo
nXEL03PkOKQk6jJVKsoA8ZDAybqyf4L51x+TDslzrjpIn/ce+qSULwnEKmZN5Wgy
wWj0Z7oV5ucL3zi/dN2/dNIX9ZBYS//sZSvL0pAK3nc8A6Iw24u01JT+LC3Qfdhv
kp+F8BsWPylpKF0mc4vTq3OT3PvvCRL27Dh5tRJwdNrW5RYlJDWLmJGLIdSZdpkA
HM978Oot4WMQE1yALSRuz15ixdK8mgO4OhHVA0QGNbirNqU9r++gONeOwdsxjuxh
WoXjz1dyr+nX9zfZxM+2ZhhagJia3YEi5KKS9OFVOkSi9qxlw+AWCdPUQdwLbhi8
hPeCPJAyTGdn/4yX4d9RHqYk8+CnxrFGtJjt1Tb07PwK7KdziC0j9QhdRmNdI/54
f/Ap49S58qOH17c7/KIPnJ4FyfaNOsX2uiVZiUU2LGACwCqSTyxKurr8qJXJaeyX
Jm2acplrucdzH2d7kKUnAkBLT19B9VTrVz2q5Hgs0iitXHgOh4VFMXlrfVpMDs6o
uppyDyhM+47XpQjpbLdFfC8HCvCoe1TKlOjh1WF5VYIK7o2m7HnHePwAsBJ9RXIA
HahZzybUhcg8S6o4FNal3DvUkRxGWlGQWb0KcW1QrwTT3PRAtlkIfv8Qk28QNf5b
bE4T1PnvjybXqelog7qUK3DjcUlLwoLJI7xbgLUr3yZtrderNtLFOvQNCEKF9jVF
TwsxbSobrHJbAI1WPtvkK8+LFmG2W2+8/aRkXISAXYGE06mlTnmLjmbgOXNBA69N
bJY7KK7c0eKu3wo1kDEFUmVEDKMGnBt0VPSIlLdgcsNBKJqXcsg/p3VcQznAHY+X
XOhcDvcGFrfLK7jlRbvNgIAa4sIwGqsy/FrMtbmEWsMoCcoTyqR/8dgpHjiM/Hg6
1zUPFRvryXpEvuP0c5EmZ0K9Ns1dgThCsGrhCFeNmCD1mZAvNmP342pOivzOb0JI
/mJkxeCkejWJzrPDTXFQnnc9H8Qnli5WQoQUXQ1VBs/CaXZ/qMHYf4pehpuLzfRQ
v7ArBROjOLlHl5n8d1jMXXsNOPzfTsQtPJxbW89DsgOHg1HpHgpTtdK0CRv+SdSZ
c1U16u9ByGSgFk5HAuDK/WnJprVXQKxUyjEtnAfjaLlXQyWtIjJGo9j3txXzDZbJ
D8QMlaBoOED2p3rRnCclOgGKiOtXqiF0kr0DUs+JicTXcRVRV070/XaCegHba96j
poRzXaTKeP8NXfCFe0xpsr5lTjs/OJLC6Rq9855yzw/sczbeOZlpC5BjdH7MtpNu
cby+B78MA9KkVz1FSaGz8wGZ1yKAcIIWsrh0j5VxtzRMGHc8rp20TIBlds3MNpwA
ZBjMoToiIfviAW9TV2+jdnBPuGn/tz/5r+fzkcQcpYSbMKN8FZidNm9fO+t3i0uF
Dr7bbD4u23Yhy4D5muqh8GF6m8s4ojxMHzJcDqmPMqr4PyNkhCs9jMbwbcimV6ul
NvIU/cMEnOJMJ+CEIDiyoH7XirVOhOmeb3A1AKJBWJmLx5rsPpUm1vWafQLsAnpq
K3Lw1u3p6rtYCncoLh2A9Tjsuomtu0K7eHtRR6vtaHuQ2g3r4SxMgP6J+qvOP6nW
328iF1gSKWIVgVpsgAovfFhzZO9eRisPWY6FB+7blXBlxcfwLaCmk4JNE3hCBmQ6
opxbw7tXVFSYzqy65QwNi29UHCn1ZuRU+gwGntlSoIX86PgAIRvgYKMe+M2Mx3yd
oaiVcxRb6KWiLESb8I1SdxHU7L9Mx/pJ9Rr14X1xfGABSPjS8+Q2UsEd7N1/S8eN
CFf3LuwWv5ENhWzm5Hp87P3t9FLRaukuemTVcvd3yiOMFR744b3ufG85rIslFBdw
YP+EZyHfpRw/Ue9CiGoklTotB3WSOUEWguLOVG9NePtsUBcqg1wPuTUfERNq6V/L
2sIBp+4FbBELVZqwRr5E+8+DATvg7hfG5H4GKe4mQK/Fp539WS/l8XbQuEWQtBEI
Bc/oHrOERMOydoNNuikh36vh2j/w7/g/8xfBL+gy2iSfiA0Alp0Tdm/s4sH5ufs3
YKhYvpGJJomqBLrc4TziTnSnyAbFsrAbtBxT5DN6GsCdqrKO8kk7h5qbNCZ5Tr6T
gC+iStU8mIueZOVUn/ycjo4Q+1dOb8EyCLeddbloUFJdl+ZOJQavcrhyKk7ffQwN
1EC2xnIrpIdFENqvBcCAO/LJouaQ2dGuKvBKxDbY40dl2MCHr1XLwREy4Iwh6y5J
LVXquA7pBbWTl4Nd7E5D89gp5Pw1vl2bKXmYphd2xrXDc7J+qtBZNZWHrETXGZ5W
RfnhLS1e7EzfBLgcwZtj1pA/U6rrLoJOzKUVUnqe1QAIbbIjEicq1FupUOHGLu07
R327GDTkCCKEy0HijoZfcRkJ5p2uIVcwAMMFvjHoQCRx3nSCrjBjgs8WpvP2/G4K
qM6CZRFKgbGt8rHTMliEEgzPwtlqPuYejRi599DZLAa16hgUIaK7xiqRuSxOkkDH
g0zFANWTLRTAgGcHGhG0ZxZYJSsH10MqdMzQPTsBamSXHvVtS2OuUw+HC1b8Iu/g
F8g4SjcTk879XGRUbBz1miAkeTGbsBaIXX9tA7ZK3OE0o/ieY6tmFNDn+5U/tCrx
qszP3f/pzq4kziTS84pCsGlkXBjzZ7TurioKKgiz9n2E6SCA5VUzDwzWL3idzMbN
cao/iRj8AiyooQPtUtk77gXLPqxzaSM05OFOvDgzsHyvVa9XmIuK22G0+UeoCqR/
gYkrCUfNYt2G6+qzIZk/kdFdYruWuX/lH79KK1irfDzC7LQFvvQjPe61hkJvdn1m
fA9F/VIeDT9ghtIoI1UBrbZbvOvv2VSZ3buoSmaV0uOV0vHPl8+LGu+aWWr7CcxA
hw6BryHVkJqIFrPy7cDB+opp0yjJqvNKno59o7BMWYqfjC/d5SV12tONXEuN0J3g
yHrxPHHEE9IkFgYzn0w7srPwpGC/R8irOeSn4qaUqzS649hLbsb5NWC3i4weiI9c
jeST1nIgTb78uD1dQ4FW7a9RZ/wihtCkuFF4gjh0J1TDczVYoxnAnqNJ3180WmpP
SSVCqIJwYVZoVxF3WmnYC0ebRVtLOv9JgxT94qjp2kidkJKKvdnK0xdRHE+YEZkk
uqRqSnbozmDNfik+4i/YALjuDJncQgkz22FHIauS9Q3xms/cQt7DLCGW6/z1MD39
tMd93IO7BtUjFeQR/X7p/PsWITqYL9CvAglZKIlAoCIeXdXLob48ubDA1e8dkvs5
zXHRdGc2D1xjA7R8OqNfvLsQ90yvf8sRQLoU2zUf8QycdFxQi5LuSRbpF6pbBKPH
970gFjpqNIf0Cqq0HBwI1orrfimjkngHjb/D7O2z0cia3N368l7zK9oZOMxns9Ej
/R4y2dwmd6UIPn8CAVbKiB2NK2R5ktNPrXPgTIt0JptiDdFpAryjN08sKti+eNSy
aUIwXXhJ958v2Rg91KN+YJFvlVS003nV8zGg8OOI4TxOvAqzfZx7SC2qYObS8a0Z
sKb2+f+S+Prg9g4dsAESIyBbQuMnxMKHHRzXlU77YSTagwqzlFXYZ3c8RGQbHQOV
MTXkvYEQ+iAtJkOVr8F3A0NlSW/w64LuRkUHZdtUM5APEVY3BD3Zqd5G+VfpRcsW
7PwPExxoDdKteQSxKaYAsjjQjNvGVO88zbpfjEPFHcnpEgrvtCzJVIITF8rmn3ow
gMOsuxNDQSk6GLV/CqDl3VT+QUo1k7O6xiG+1n2ABQHcOJho7uhLJakzTfr3QUB8
vVpe1OBHVME1jTk41YyFoBd2wc2Uii31vbC4D0RcBT5YnPbwipy+uQhi2wSZEAbm
CREaDGWlvNpOSpkXinj/YujPbIGbH+ZtXH16YX8GE+CTuvnK6xGNO3/bBVW4mCA1
vjZiZKFxgbWJtQ0pZtBj6bX42BLL3/6y/khVw0Bak5HPGAWzlgJL7LDr7Cm8ges6
NBeYJlpqR0EdrragtrsT55PkAUwYXWb/5e51Zrch49Pk431+jd14XKm4ZaBA1spi
Mbt1N9/oqR6QTBJLC8Ei/ViWHY1Ijv+wTDNEXtt9oRepnMiwrx3P2Zx/Us+dH0TT
dQ7GgSS3kryvYavCP30vqRJpMkZfWRGBQJA52HaC5dgSJIBF6lSmEmGG8ZNcv8WY
j0BQbWNpxm+4IhRbqte58NVCZo2YaCGPSkZruZBfKhYPrHJ6l4e3E6P/avC2VF1e
hXHh64EjXDgEPCgisHiZaHjjDT/bVI+jLJxF8IFs87hNkjlnqXP8Z4yoRDpsdQ5r
HufN0OhrdAkjW04rpBHeMgXlZcXpZRV/GTzWDlhqaEMwEZmWhKYTxkP7Oe1A70t+
CPZ5lQNC1bUN7/DLAA6Md7VhhMgs1HfpnLASP3qX6ElBWBb+SFl+PCt1gdhYvovi
gYKm0UvB+5LpZxEXq0kMW76IWpHq6X4YP47978jXOT5YHqM559lzSCmMpjf4p9/U
KNTnnnuJZ9tHoXf02iEuTF+vjwGu2rV4+ELn+MrUgaVk1NvDP38e4P6FhzGR7PMk
WxUAUvMw5/F6Okx7vctXRf2EQvCcrDBVU2geZlQ1mjsO4isQLK3/fc0AxMTiv4mz
b8uKwPOZhzyBYbb5/i+dd8kU8sYVgrtJtvCEv7ub0EIIXyBuIY4XqGnOs4LcNOwl
RjbaKA1B4CrIFsgX3k4FBTEoMgwnYwb3TMrxepkHhiGn5N6Y5JY+LBzHzO7iAeNe
vxZze+S8ftriJMCPbwXtJJP+FUE3W/rTlGa2vOIhq6+YYJxBjDTfMHpb0MP/kR7g
nCH/wuI142o5QMpvtGSPPE0FrG8o9o/cVkYjbGa9EhNx6ez7OnP4NXJNDTN7+1ct
0g9n4hXtPYoRognY13zBVoSY4B+tZ3fGL+/sO99cVkx0qWRg69xmIBwb3aQGnzp1
LvBxSAiCupG73TQUNxPii7rzfM5KBWPG8gVQ5MNB5h6NyZTQVNZtRjASpRexquy6
Cha82X+62Yh7OyHhnFvfgHaGf8r+vW2Z67MjCUElw87N7LNd/4s7tBfxWhp+WoOa
vps1erJ37xVsgx5+HldQHBgZLu3xwWPgYLT1T58A0M0o5fT/9l8VqNbF78usWixv
N3C8DSdYl0BelYZUOw4w57FjTWlTEnkWiIeN268kom/ESb9NkFpkDRd69n+D/0HK
xsw26pxS737bH9KDlCoL5C0yN76lcQgzzfnUeJqu4u0gtfsQfMPk7XbaGHeGPW0X
3a4ZyeG6rXMb6tTOHGEtj/nsuAO8tab/gjKmI9yNEoEhWr0NLqU2z+mCcFL6cAkA
Ya+K54lJqM28thTyh1bcR2Le7kr2TfefwToyHmv05oJ9DYQJodljyFGfm5oCv2AC
2foXCbUnQPZ2npr19OZmeaUwmRRcIvZPHetkoRjM9aPuLTEslfMayfKpi7yWWLb0
O8gyfkeF2fjLFQbra2KXuodggMs+jsNsDwxws/wrTKYjL05k0zfHTxxm520v8eTZ
CySyl/XQaC+DJQVKqTxM9ar1aEg/mgb9Vbs322+f+yYtpUb0Oi1/7QV0L0/UUC56
1b3z3Pf89d6dCY3WfRUHDYixGs+CnbrvxP8lSHrNbrpkfMlL5NkHRbPXhClAyRK5
W3amqwTDPufrRmO6WgBBQWKNy9belcv5MP4zzgAGNlEe7nZXvOWUiIGIvD2eGeIq
J2Wadk3kfJQVhok91T3DN3sWsS1jMZ5gGiaSrDEcocQhWqwCMjN0usXw9wMhn0jO
YAUwYlKqNa9DufpqvBPlH/gaNoD59IVA4HdrBqk3ClnoU4d6sEhhpcYkWVY4NMa8
bPxWpZTBqEE3+YCeVY5P8qDQ01KXTfj+Ba3GJigaOBJ9Vb/ECNr/qqo3O9xiZwnh
8sU7X137OiUzU9erulijbvx87VXoce5Qv5i9dYreAESMJa80Sfsjzz4GWauLDIgR
d0jGV4vq6Y9O3Tg+Uv+pq2z9OwvSGovK8nJ8MR8GGRSkAyCDsuVMAp7PhdyGnC3k
SHF0INdEJh8apBfSIn8/m6B/0DbUKHtBbvmIuDEA5faQgmYoxG+PRgEoIRz5mpEh
qlcki3gF14G4ooa6bBs4csc5J3OhL8pbFw1HxT5D/hVE7oeSzPA29cuYoUBnisp9
GXdP4t//QplvBaFQKY4WsLj5fCwlYNJCzXaOpKRKBSellfewYEIZXPHgGlwkoBqx
JZDDVGmHQ6sa2H3H7mhnx5agWblSt4H29sy7t7kk0T7Vgvnar1yqc71MEvai7l95
qM8a0SnOHHUi293UIM8/s0Q+1HIACHp6pJRxOt9iNgBdRQbmApTBelGRXw9Lltt/
paRjtmSDBWoak0wp43l820keWpdHDvryc1uLYhzTgFeJHSMS7klfLFkbbnSIYleK
Rde5VQ2RWf+2oo5G1lnXZxF/hTURYgHv+0qxr4Ad7OuhxelLR8OaBr2ttx6lf3Gs
R4kYVYpsu/l+vIuy/frBQftIHex2vrVyxf5V+31mWR61qbR/EQ3ni18iugeUoVMB
1vgppU8ObJQ4NPXo9/OeIfb8KZh2+tV2JlCJRP6MiRtPENYsC93goIN1BsmufjMM
qmZf8YDfOiC8HQBsg8NOogWvixoGiQzYiD5fnaXi0paJd9Wx+y4iatj4I/oRqfNT
1zOGVB/u2RlSgzlOz0goiBWjeaa5HnoSexAU0zJk/w+EofLrNyXszvqia434Bk2+
Gr/XicBIHfKCKzD4olQ7uN2S/Y3YoXGeKm4sZzxLGQDUoEI8PR/syBvqxDc/3RPT
Qmz5sI1fATdC1QiI+4oeeiyyVQCirKa782mnR9ltpF6yD2dUxjPFbPlmmD/DUaaf
eNXuKYi5X7B83ahrafhCpnfY9iUK/SA9kyLapyXM5j5klTTBMc+L4vQbgFdoOo9e
ptK6O5Votf97K4sBY32J6NHDifkqxoSaXNJRGsL0Z9Mtp/Oc2t9WeF/mr0i3HZLi
dlAlNvrWQ7dl9JYGPlZz4YReVkgliyog/4KbEhXRvaUxbuypelMLAOwe9fZy+Y+M
8yZEp9BaElN1aVMUnTZb7HlZF0P6WVfyOw+wgqBsuv33Qnm/Mjj88M1VgdPdrbls
ho7A4cubVS3ym40Gwjbrz2gb7U7t8x39mLKhJIK5cRi5upNHYPl/bT4o7/K8ex42
JvQnMa7naGwvicMVxLTUEZVSLOakKX8tK2cNHLMib2n7tBubzhB5zYaHLmCHjK2y
5KFw+IjtlT9OiunJ6LJGivrIzkb0qIiHiggqSNOyJbCTrhLp/0JRj2DTinnYYghE
d48OFdMloVgb+WZvMf/zdSBtk2YdwmvMx0ED8xKMYQKCJNNAj83L9Vq3b0xPZsxD
TrbRprnpwgxs1bIA9M9gCRcDXwW5TqI+9qXexeCGkzJMErBYoNV2roBl3GgdcDeI
YCYiQ2yyefjD7LWwIDqdj9tP2vqr597SORuGGQTGP+Cfof7Rg6PIQ7VGLOL21lzd
OEc3pv/wK0nr/5HDZ8aah+DOidUhw6z9uS8cDmKvWyoIPDJfOknUdzSDkRNjHPoa
2TarpWV/w3NM8AdcMj7ZDgPh88xztmwKqx/zUWICiz5D5Oq0WBVebPElP4IxHxlG
kEeTh6YbDPov6Vj140Z8AOS7FOyCLUFomG6slk6tupINdmIlP/hOvVKi+iU/op18
HSgNwLdbeBeqzXChoEOdk1RBhBG8vrGZ/Cd2XBORIUb59WD38uJOwjHJk4VlZp2g
Az2xZIOiGUDeCXwGHABvLHQSulQlI6q2Mbyh97qad4O2vmwhF/MGXH+9fwQOYWdz
R07qD6oQ5ZmKyrYDV5dA8uH+DwmDhU4mKdDHOgDDxZO2UMPYSC4e+7F2Xmc1gj3N
5+J6DlofPAECxn98rmMdEXFki37bmxQRPZuL9g886Q9Fgx8i6SJZMxR5lb5L9TE0
BH63WSmp9gZZ+/X+iIi0DxG1VnXVjBTHxqCzPVSuGE68jlt5S2gQGnq1SKoD0njg
LLla1E3O0JONMRrN7vxnBHPja8FQtCtbItvhkPTlV+/rKJ08oibjNuRf9M4yxwZD
i7hl0RPr2ydZzLIN5+rdX0jhcMLXZypkuvErbAzDR0ACWYN011peG1wsBxE3ddXx
RCiDe3Wwv2/fef/QzyECG8RoVpEWH8bJt/h/ze/2GCwBoC7G4X6taX+GqyD2p+03
uTmc9cLt/olE315XLvbTvQxxa4OUU9awMAVzZylz0ujJZV1JbI8qqPGv6fCqKU94
9u+ijxkhwnB8qqkqYUzqUpuLn53/UTrsZvOEpeXoKhS/z5O8+wpoRBC6pGKaPVL5
bJ8hxbT8jnDdNfi+OKfCnzFyCbiR1PUgnO66ZGGcv55mZkoB/QqdC32uX2Lq8WiT
KEgbdJmAYbo/LGd+KqXTAOv4A9uGg31J2yAHcKklYQA3fCiHJmYYGdJT5f0f9mp9
SYM9kxw9XT8Xkc5E1ay7ljakycAcMx5bK5NA3rjoDyM+lZU3giSXneCMQvY/0yHV
IV+WR4DEdVcdSVD+5EdsmYikKDaWtMcMeOAB33mUDS4IxPF1o6X+HeWx/svIAZK+
8U1qmwHVeJpl2YfkgakyATOFpacr6FTqi56Vbem6MlSL0yKFtptoQJetzu3P9M6q
0MxsBwuSt4MeeozXUI0qHSiSw9A6Re8t4+/VbSixWjw4j1K7NfBVIZtPIi+we0me
O1W0ec8eL2nU+tW/w0/rQOZDa1pj/wePNgfskVds43nS1Jl80bFBlU8Gan4uSrEB
iJ4MWn4RiJoO3yolZS7TxLCMdLWBVaWj9rH6+W2YKlmLvgHNTqi0WIkmMmIdPxWZ
yKtXxWi1ZsX9ZGIvv1FB1o1+t2p4ulntCM2wF2EPRgdZePqJf4D8mZb+2jxgu5va
9bJNb3kfGioP014xXhuky0ZSI+5BEuo6nWUVQsBhv+YteZUEuJNryubDShpcSppN
+kQ3Sy7hReJ79dAV/Ocunc8Qc+Vo0Cz3UWN7TMrfAo4rvV7+SA4urvsuakEbEJga
wd12j8FaTsoeOPbKQWdUDBXo2tJnFOrVU7eZaSvEUBlmACtpRg629VXsKa2Jp+Lv
MGFcztIh5JCGrxdlshRzCpv9I6xO0wxrmVYlplaF4wDOYb6abPXQKJwI5zTCTCQ+
49dWmSSfI497nuaRfxg1SzcaGdQBzIi/snnOcxIabLMHEVIxWU8WZToqiwP0LtVf
3fj5TeXg51H+dn+byXJYSHRpSb/WN34HIUoUQD52Srf5M7cIZncdGQWNfhz8sUIz
z5yH6IHwfOKdsY3+GcH6hiim3/iC7rMm4KnxRu+Hv9J/Xl5k9GGqbALKv7jLZee0
ydHiSPxiwPA6pl24aENlwQcpa56NdwxiGuUHl7POAe+TDIpu9w6NOaM+LeSSqWw9
c7Llce8LvT366ZmXDYS0SNARMiKyO4YaxqODEBSVEj9pGuqeXh9mR527EHwdTlcb
AY37pgeADGDCf5DQFHGRzEPTu27k66a5U3BamC1l4ykA7cdgSdKz9s8MMhL3vdL5
LQ2VWfWurMFA9U+HUuK7VDNEZCaRmyTCLVe9duCdhAuwrracpkRZo38pZDomc6zs
eeK/sxMy3E90zOBTYHH/XVS2qsSyhSP0Owj8oDMjLsXOuHd5P93uDR1dL4dMxKaA
UtD9ZYj7t1RJ3hOFAjUPRZ9l7R9UiFfDWKgXJ7F6S1q1ucVZvO1W094R5QC5MM2E
RTdhtoJp/OT7LYzIkzd3JjW7XbdyR5dBfnFvImwdFn4HHgM8FdG8BtvgqjqVsgqK
FGsWP1e/nJyCusLwuvyKUyYHWimZpSajOg32Y8lwfSdPNKtsXwsSOkb+0xNyMvgI
WHorpe8KCNifRkLBFqNQZOBxlfmuu0nuJZHmQqTehLSHDBsTBcJ3fk/CZpoefpni
V9RXUVwUOCT7+1NjSWCIhPgKv1qzE/c9MuyBlnzY6bkdkQ9ay2UG3eT5PNFgga85
NrBxoAjjZQBRMtOIDIaw0cOwDc3u7J7goNJPqo1P8RUC1Hu8v4xpql7JBiLeZhoG
5Uxm/uBh7EOEzQZwudnmFaIDaIv9To9tQFEo1pG8mnFs4u4nSCp0/5CvvW2Hh7RW
VMbe4irUcYd1f5S1UqWg/Bs3u6QF/nNScuBWqn7kNWgFoLislb3u8IdDLEEusV58
gUWtU/b4yaLhHiBqnsslzvBR8cZKCkL2vkp7/8H5gVGzcOACuq1A9nuKx39cSfr6
k/se7e33ILqzn69LfZ2H9djpEKrwDOJ7ZVKDi6Vxt/RdZOwrkxLwgsHG34SzFquZ
SddclKlM0jXIdH2SLntP9qmckDLXFD1DpXG158wv9UlfyGDBN0FwGhN2+kEkno2l
Avvf0xeCuyBStMYiVz264ULuS/ubLkfliVxOdlo8DwX0qkJuL32xnd2acnowKBkd
nZMPCZoYt75S5oh7NnwDfKpl7t68V/A/3Ikc5HKN2XF/MAAzB6w+5BboegeKLgsw
MYXF10jp6Vfw4kWV/u17FFXFPguiSRgWs977snyWtZikdqkURdR0uqZ5CodO/L79
58hGNydhsvyw0ben43m3Zkc3atIHvxa0Fg473Oa9PHqoxKgt/mwSuD4VlrYD3IFn
lofyGjE96aH/qh8qrerW+th+czRzWxPBW2NPzT7rdpzAlJFzHRmJmi5B4BpuQrYn
ePLmqnb6tYnS9er1jpnXS2bpewNLO5WpXXizCDDjZJWOC9S9bQ1AY6YhCU2xL7zl
vEKqYlHVoHi0w0v/NU831YhKkrb+bJueNGwux0H73OZXpSMj8e+4Howy5uHcrqd2
qRdSFmsVU/lImJKDl7NLCgWDJUROfSmtCbWPRhZHPpTpCD9aoBT/FhUKrxgzUOtT
DF1XFZEDJ/MOGwx5KOenxADsTO6pyw6ihkmin7hSYIltdwDQwrIs/AVOzRAIYcgp
u5kvqV8/m6DKJ0daLuMW/Y00XC1hm4+OcWQz6qwe5UZxrxF+kpiYak8CS3fPXW3t
CvvRZrLDdW9fF0/56x/0xnAVjN5weiak3Ph8nw39Ww+00rpM7g4L3wfg3d1HW78w
NwbwQHw1srZOcb7d4yr871tttZkW+G7JkKO1shuVzwv94u8adp/k+jQaK3Q41IWJ
fCkcbY067bxuocT/gevRNYIAS6cs+oBa5ntB7NX63qLy8Z2beRLh/z3YVv5axDqo
PkmxKrjIlS1dH94km70Ho6NMnqLn2Lv8vLHVglC9yJ/+wX/AKqdWgGLxKtE2ZunR
YJk/GMDYRHhOBIHxko1H1bC3EgMqlgBoyUQw2htfVWF9STGZb0qGmehIHdNxpS0r
fdppICeYgX053QAq2DQL5sobGf3mC9WYv/O4vcoCP7rd1uCrR+0ifdOJVVQN4yp8
tmE89PNV+q02OOZlczi9jpqYEr9csJrHOKyU1xcowBAjIFS/oFIYhysFRwlktCHz
SbU20fgjL+xHLrYsSie/onWkOcoNmCamyphIPjN/O1IK7pG9poDPZwrMePTx/yFO
YHqVfS1r9M4RnKepji3hWMSAh3nyVlQO8f7GTkVzc/8zIB4TaxcArMI+0h1HtEpt
Iwl8gQCBSWKksgtCcqVlSUb2+NaeQ15dBcP7AivJZupWg9paR4C5Ryaa7BFFYFCo
w1GfluSUQldEbwYcNKRS/Ha+mgWsqO3W9ZeLjYCwQdal/ZSc73awixnzdPDSH0V8
PBMFrT0UOTBrQHl33NZ7VkOwg+fch1MM4vaTsjrCp/UN9B2ZT3QCyvLUt7TLsqvk
X1yW1BXkCZLFC5QIAb9Wx7CFfe1mvbFcY2gFaoVflVS8q5XWEvYwlwhLk3D48cYk
qaEdrAWUVLfnbPaQHybKiaxBcF7I6MIoCmJlxha1HULnZK836Qxu1KDYCiH8jLIm
hrAop+QpcgprMdc1qeR26ysM6vuJKCbb3hCgmYVQv0DO1bbrJbF5bKAXKtjrVoc3
GtqFSXLxEJRV83WinxcZ6JfsZSZxz2y68HpCoDMlIncKGkO64NMJaWwMEPz5F9fq
xqsaO6GBhgw5N2MsNsEC7DOeajy1yi02MIRMqCt9ZX8UneF4CyeBXpBmddMutPfQ
qHQ2spdgm9oO9w30F/51mClH4wvS9SjiSJ0BaLQSdaNuWZd9t+wU8SxTgOctMN1I
0jMLTHsNYlaSxvq/FLEjWbU733B6BIWpn4w9PyP1E9hkptbtKP30pK/4jb9eqXTS
QBVUni8yB7SY8XHCGB8k9jLfzrfrA60ou8vZ8m5JoYPKWw0ywMJ+ExuPdYPtF3+Z
d32b6OW2pnif6iU2ecW2vxfza0pddsu6vTE234qCgedaGOSMLhul/G1JgRZ/IKqH
bjRhil7McgTkgBqsiYkR/c+HKl5rQLqWT9biyEhXKiYgVf+q8bWRegDYM9UQpLpN
4FfBmCdY6pdfMiQGvYSW8BWs88BYSNgmgYzFRKkIsyceFi/6DhiKkR9kYHJOhUp5
csSvrtwzdJk89GQ1HXhdRfq5c3wPceDQ/irclUtZyXfPCMG0FRPiDHfDFtWJanTU
JBWTRsJFMUcQrRZL110z738P3GRVvXLPEgT918Nl8rqoYorNf1ihJrzSA/X6MuO+
RRf/mHiA0pdIr1OEoiHhrlQaPCGLj50DlxabcZMZOjESeSGeTeR8nuBUeJzGS1fE
unqAMy/yZRzOqPXmRfvM6nXK4ZZadNyflB4+KY4Ntz4VCDUmYRbHodd67G5qfiW2
bwqhKBYprUGWq5N1rDyiqxl6djQtPM2u4wslBoSZtM+j3ruWqNo2dav4G5Cd/zeK
4HawUKtdP+CHYJKx8gQXInzZ1jzwvwKzXawieM+WTmVhe4p2tDK7J/vb8SDgirFL
KclAWubVQHV961b1xUQGldFLQq+MQ2LVNDnrjPywGny/f8uej0s5lvumeclf8Oer
sEqf4uLLU74G0YRFPGO25TntUq/P/JQjO4/0sr6VqI1Ki1jN0jeADzahcmYKX9/M
PVEIsxJTBm0QlX/yVMDKh/gLumoTk9akDBpAVDib9MF7rTG6SCPz0EbuGo/XJkhg
nH5eYlkloLX6QJOle5+BOz6hhDhtE7e5I1y7Dfel+ibZoxf6/qO32w3jWI6x5zD7
cleef7X0XukEnJkM4sxIplh8u5e/59Igkf3N2TvxKRzkv3+LDrBfoLlaFVHhxjDC
iLUxZOmIN01b5UxWOeePoXAQePOYqGjdfgwqWfXrgb5KuYD6K81WGr/BYLTvZ4ih
ntfn7I4619gzG1E7DQYYfZks69+31HOnhHt8dBCYiJsqTkfFepZHxdfcHuzMtMzG
IjbcIeY/3k56sb0d74FvRgdUCnIc2n57a5E5Z6UXN/+8rgrTyDeDcN+TRpC45DwI
PQ8P+9qExf6kAO5P2uZukPIOrdfQKw1SG+i2a3QDrDcic43/crM1NRFOO+CHlJI9
gBHZwKyhrVKH+IGWvCHs6v0EDGcqyM5bF6wd/WFRCF+ipihrsrRrX29nX2t/8ITL
95JTF6xnZc7TvG1rCl2bKh+tL1pC3xrAhT2eHnefSdoV8fbTZhwlv0XmoqMR6wjb
WgLLJyXNon60UlPlmY26/AebH5sERQ3TqDsapABZ2Dbfe7oMQhjdH4I4wZkuaZmm
U14lsP22jQIbjw93AAiy3AgvYNzBL3brk2IRZjehG9dQlhzfXNi6fAYAhsT40xSI
U4GdsFcI3LMx0gi50TTUwhXBlx5qfFPN0DWoZxVzOeYZKB5ib+jH4G8ZmMV5mT1k
+mg/KcWLqFPTVk/FYrNjcrgqJxl4EQC0ldOKTuKZvPuDToPNcobVAyieBIJlDVwt
kdZNYzQ5BLbDsnwFkFUoQWFEAbbMlyB4fX/FDZtsYRmTBBIrKWkxzGzWZbylPAtC
P1PVccSJO5KJKeD3yPO7Cg3tjvSY/QYuZNTs6DyI5377ZMxwIEQ5pU7bcUjAVG+P
uTS1oyRfgBg9WptbA9xYgSK88DKnpejqe5Zd/iGC3HQUP9e7CgpLQtToo7pty279
STq9M6F3p5z632+4J+e4waI5Ja3W6ObD4hcyj6ozrwP7YzxHVBLx8T1TFSNn0xyy
tmKg0etbcqoa5y+Y1rRFnBjNLtlON4y3/FRI+kNP8uGp653XgqutmB125XXZ6XG4
+SnqNQKN9wRpZN6BrgECPBY0l5Jw3dWHqGXvcgLKpM1yOC4AYKHyqoFw7/lU5twm
+3pBeQG7v4tUs7tBnPiIVk9T61e/3IrFl3flswdHo2dujD8eiZTsDAOZe18RX2u8
3f/n7hQA5RG6u7XA0QTw8lgsYXrqM2sj0XhWpiQlRArjIPoozVHdwUIrh8Ozw/Ns
9nD7Yos3KJ024PuRR6fM570ZeE0cJyyBz0XVNu5E8sCXi//Nz3Wif+qawcHgGYAd
c+2oPaU+OL3kQfdNQXXbGa3gm1pFbIT0XuIb1OT2uKqpxjLf4/a46SpGW/McK0VJ
waOgq8aYiLzg2MvAepINWLJ5uSxCy1Y/JZbg9Zne74+/dF2SCpjgusI6etoq0I4/
eExUu+0ERuZ32aFtFqBZNm2HGR93enbkbb3mPlUp93ZUpw5KHmCoXRENMO+s0/fj
7+/1eQTgLu8KiiHcE/lhcIDXyGiXL68xumkZ602W8ua9n++HjnQ4Q9fOpDn4zmCX
VIy4aEUJFuFXuh3YuvHH5ry9WIv6hJY46KbY/NdM9JWEoQFHSyoywe0h584jPt2t
gUiCFhhD2Y4XPgKl9uvnt0XSEZCNQ+SqYgS4I12wdWsiT7FHE0f2uttuAt1emMcK
Qsi7MiC13zCi8bWyIrw8uw==
`pragma protect end_protected
