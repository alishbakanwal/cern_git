// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:05:32 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
BS2A4yaPCrcrHQfVvur8LmtqczU0E/98TFJEHVDsGvGjZexJU59Se6yhYglUJD/j
obf8jvDpmCwsGSS2XqX34SdOSvmVvdcCXt1mC+XevejbBBtIrPTnvxI45ePFWYem
6sZFXV7Jlf58wTPZ9uwAlzF2XXF7untzEF6KFAX3l8M=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 19632)
s6bOs3tztvWLm5G4IwgKHkgTDBZXARRyJypvILnOWQlhUbLni1vP7ks/Zqze32fQ
O2MRYeilVJw2+3MNgifOBYhAIUwBLNYBoL7qmm2sOKz0W7fOSJKkbRpLTfnrS5JB
/8c6b6oYwe5FuhLD+RdCRU0klltWx0K2Q1V+dNEQcJLxYMNKi7MNKjnCvxUZfrkj
COxfNMQXrr2pB4W86s0HNlk+sGz4JGqkXvoth/MwuRzTBN6Ob9K1PCN2HdYhXNKm
+hkAlcg2aZcHynjvCjkq35PA9P5aIC0dQ9CeBLk1eRXerJfSk3E509EooLFOUFFW
M+dT1fDpLSw7UsUa/TEZfTO6MO1jVcRvvmh1/FwTYjeG0lzTMN0qWuaeoOxULUMp
AW3eHaaW3n1TLU4Qv4areCH54YvUkRZ2jc4nSR07uvmSXpHdHO5GNd1pWba0dm5O
ScnYlEKpEQOKbDjZhPvI0FLosfmhis+qtB8Zdaax6m6/7CybRQlT0JQNe+O9SLnJ
1N/tMRd69BARwjoYACiW7oQhdApvEBIq2TJDiNgyuLbdwZhdQ35WOMLYZE8xzy8j
TF26+iamMhd5JODjvNKRgUSHDX3qIr2q3Xq6wELnAoccZQgHOmxuZvGJfpVjcjCr
52hZTLHZR+EXwYRGl/muProBNyigD8dzP4xAutK32SIEc9ohZ9UVsLr8e3bibAj5
sLU9u/D9Hw/YjhZEnbJCQfGX557Ksr9xoU09vHbFPue1ICdo5uWTOlCh5rEg1njw
gbV1Z9mmyvuMUsLxMhOrk41NFt1dmnRGnmXW2u7APaLMrBLSaEmQR52UjkeEF2bC
cHe5ou8X5cDN25msUzekam6pwsP0htPcauiumZyN48KX++n7o02Owa2HkMSzksmX
kyzXNPm3GIjmXvnL0ULry+62ebdV5YP7FUrPo213H3K5yGKzeTmCMMYwDS612Dt3
+DSQXeHWjDGLAJbISUIFqh6NanUgE8QE6SasBCMK3zeQ1JLCaL/vT7zP+11fEFGi
lzPMYgzMLH9PbHLAPgcqH1E3ynf4C778XSCXVvcJqhG3MbXXJrky+Y4N5eFlK4yF
k3GQ7GE00kSHE6EwYHoENJNYcnHV598Pyxt5XO8MTee25gYduLuW4ve7cN9LpeJz
xTrTfodfASWbikfrY7GhB1v+6+c1TVLiLFEp5GOdb8T+QA9DpyDr57FxREsfg65Q
idsQU9rbjz3Yv3UOmHt8j8hbBrmKdVMDVWrLV8w6gdoMaw7o3ckMAVvYUURYweFo
RxpR37kv8Xnd9w+/9Dhnji8ZrrEe8sMUdmZnratDekBbGmZsiCwm0Zk6wBeoKFJN
Qm9dyMr50QVAOJnRrCiSKhdoHjm0ZRmor6mw2jtQ9BwUiib1tUn+ky45W1RHA28A
LAbHt4gJ6mhLQQZ94Ls4/NwEPNWFBlxKyd7Xmpgl6YXu2Du2phh1jca6ooM3Zu3R
NmVJbvw3/Y27WUwr5ldz3Gd9IQM3a/q+xF3ThsyQd2MN3ov5jykGKpY8yzT0pF9v
GPF7+Vv+3ATRfrOpSnsQ4fFO8wVYvBp5cyflC+KYqUyEbbsS9tii8e+qenW+xC47
bQnGhvGW9jtjrjlm7u+IibkJd9kMk2EBBMUgd9dU7jlGNMwmyi1vlS2dex0AZVPK
wM2CiRVgKY0san1aTrz/lCFoSrobC+CGCBvi346hYtT4oWSRTSGxAWKpDJWAWae9
7De3yLz/szYhIkUPNpE3GjLaoVmU7NYJdKLJvcNmHV6m1leQnjW5+WrsRx9QGM1W
9CxzMRregKd2g1YqfBrbow9dTdR0AVnGPfWEAryTRFP24H5swYrobAs/WzxFp6BW
10I1sySBID/qyd6oya08/kh31PSQWTMgD1YfakGWRLRzfckOh9KQ1e//M9A0E6+b
bWgzLY+tiDXvmFSUQ33JnZAmW3m4jdf2H4edgA6nYV3S/jrx+aOgNWGISI36N57O
jBRredPHfICyD8Tu2zC8jBvSHkG5TxkNaGEEWNj2PTjIk9299Dt0m5kwp8PCph/m
YRUvszBzkRnngcOpITQ7QGRe7ku7ZHUmvsfDiZXDKcoNvfcvFE2bFiO5uNopyrHf
n1pA2fHdMnZ3RnN1qpT/FEMtVs0msyDMV1OAVlLoLnmdzhyT89euI2e1QGNsZ2G+
ayBFb+x6hGVCa6E2HqALOP6pH0rYuK88QBs5A8fj+09l8dctWlBsD8kHLjBBVICB
U+Ahe/+ymYYAlMiwu3l2bRf/aryDcboeIdEZ3XM+4sYKJS4iFCc6lpY4L1/CpMRL
NWNyeJE5mNxCG4A3aUBA1vjGiIbDXLAYSH+QLfn+RjFU0vtPh4+M+Jp+LvTNLQJA
FbHQiktKweYCm7Dl4cJUArGCNQAu6sYpGeubbtajj5O0v/p9DTIPIakzZhugIETw
wvhi6lvj2iZbBOwRbQHww3FJm+z0bqBBmYdorlFKn20pKq2Xt2MGNOQtpgna9RV+
S0jlou2JcyMLfP22Da2vEsIQasRAIKGiiGxM4jb9OLwucRdXwxdM7U4buKhcGljR
KBmLmBnb/j5sCUZyL+zd+0QXac/q4cVUCs6XJN+9oeVLU7Q13CifA/NoVG1pP7uh
BQDvsd9Kv+TEFg3rZW0huUVQ4kF9G7uCBGK5oj2YLr6IVpzU285GHHBWGI91hgkz
ejViESYcBxMyt5JOBOMoo03IhCsPGZJXX/AOaKh/Z0Frv1KOHuiMLXOfNb/Ppu4P
lQPEVnsXewbjkw8OsrR63emcXnwza0Z6w6PX3aUaiA2V0JDHKyb1jtKbhFilezd3
ycLck5k+p9dxBUdMd8rL2gHxTs5sYSnVAnxbk7ArCO3dSm6633x04BF0lVatCTSN
SfhmjAeVl8G7RBQq2dopWvaZBtrBFxrdIS18KCqXHFA0FJFLA8npK/4slPNDQvIN
Ug7T43oq1KMyZprgjj0SUiynUasPebM/JiYZZtvJQkYa/MryeSuPMW4HLvvic7R3
8pBV85m9Q1s1XI19gSPiCPHFBI6YctQPTERxBjsbb2hlFABSBYB/tIuIFzAGxFq2
JuANvaL5fCs/XekaGS4dQw73BXgpZklVN7Iu8DUus7g771fCIB8jwdge2m8qquev
TeO4lwpFj/8naqz5drS9ILdccN8JQjRIved5QLaxoh8lS6F+RkUUbx3ag/VRQ58h
p1kqXUcNfZIPoEMVW9/nPiBkv3nXXNaFbvuPqdP4xgFUVBAUZ7vv6ZLDiGRSYqSZ
pbSsbs5c0elIg45KbRWH0tpk/VrVSFLd3V2v8zj59+puolClK8RdpW8OJvsVqhRk
a/835P2oZuox6k0J0xkd2o0NuxeWG/igYDztH7Vgno0+kOTcHtkny/cz7Wj6llO2
zocmzYswV/1Qtn2jkxnGt6rmRIpk86wib1aZFhP/vh2MvS4HSVsItN5VRxRewiid
ffoaE0T5DzwUMwf+RzsBnt3mjLzTU7KFh8pVvjDCQjOlkNpBukPTog+csnzTmxvR
+N1dO6GwnZGVvaJeE1C1uMxAVtdJmd/8tg+7UudfSHDHIUQal1fCAnSoWlccTA6s
L64GP2rdDYQNsN93RQC2jPDSHNPRrkH0TOmj7/6FtV9fjw/zDVxEIMtJcRlepkIr
7N4mREU/nZvVqqvS/A7OmIBLLFbM5sADzjjm5LOJ/5vX8cP6Ljp+jkKSqEJ3HlWJ
lnHnRFpZcbtK9srrymvXAaZyHN57lBCBLHSfQrGT6KxtddnQwxoGm6K7pxQ9/j4F
u+xYNXh1k2XjMjLaJdOPdADCwN4QZ7ymD9leV5xfBHslj5SibnF2z4hxhXoYFsRD
EJ3ycHR42HNXzw6HPuY99Q7/Ut/cejALeEX+5Q8NegrLty1HVemnwb11L6vDiFNA
FfvPOTJJ+Yj6pZ/ro02GXLmjceYObL1iWbH+/F/l1OwtgSE1oDVhQUfRpVOCUckl
ex+oQqMwc2Od57LydHKL2spkKIlkbHglaC0DXGbG+ERPXtPXpracIMDrzojGz96z
4CZ+LqePN+uTurmN9nqbnONMqW4j35gnprOMJoJ5Ul1Yma1USDzVTsFJukr9vtbv
eceaHDJ3ZKkMw63HfIfm9InVQqtbfP9XMdDeg+0o11CzGWTV0IDJ9jq1qSMK7wvn
Jus07XQyhfkjw983BdEsYaZ2N19ddEFJL67oAK68Ra8Q6FuUuFnyPUsuHAZvIJSC
uzzTuQYZOO/tUbDTUaa948N85eGMTdspnybpTdPt4DZxj4Yc5Xovcw2N3N16Wqtd
z+oSYEQqgNiSN2ejXy6ZkjpCeTekH9DuyEjdV0f6cPvb5jzGwgB6S77G5TzCjT7h
gpI1oPM8fPinD01oEciCNHrlo3Acr1cK3cD5aVgyB5F4r94EeC5Xc4VnL2ic4Mu4
Tf5O8haA+0PLkGGJHT1gt5a5QOjrII1bu7wZM9SEsZyPS6VTbOS0nuuZKfGf89nt
olGUMpApb8PU788GEOen1SyE9diRlS6PIZ+tfLs/qgDM4CKFanz7I7fqMTOp2h47
vWHO3XGE3j5lWn0HZD12g9oMYafnG4vZExyMWVzax4YoD0N5KQMAUcUVCUd+Bfa4
B+WmVtQO6Kn+M0xJn7HcVOvbyjch646UvhSlEcbRcSdb0VSqTRoSZ47cml58IbCK
Lv3LLiQ0IfJycrMINXCMLs9+38HWM81r7dbbP9PJhAkGQcgn2zk15kMPMQO/q94t
eHGEbVIEPEC11pDveIjR6EqaIOX74jmSHP318VhJPFxGmXmwgOluaTAhwHw2FmHh
FMExyEq/SF6Q4j20AqGDNWtWbqZA3ANedDbBRak+TeVXBz5NmBNmU2+UOMEaMq6q
fMAjnTsdw7ixjvhVZJLXayWNePsk8knhBU/WZ8Co+Pjkq9c8yqbVXDy8m2gkyHiL
M9z6iSkiGLd+zqGz/yeM28iLAn+zRv6ZPDPSAE2wyz7TZMr0E56LFM/7ZNgy/w61
N0K49rHKRUd+aQlT/SjGKQdF+0ndz+n235Yyxfwjt6TvIyYN8RX2OYqph5+6q8xj
fc4ewBHVo7Wxjfv2dJmPx1CxVZ92IBHiLFd45NgN71ex9KxERBTRKMDF05vbNl6g
SsO0P549YZ5uJqaca8Y3Mkq0FP0iZATCv9cmZqgztYFxU6BrLqJFtTEApyYdtdV1
2Iglw1OXv1ashaRg4sIYf5KQMSOiQPc39m8DD1jjFwyXcndzoiPX3HX/yVarjB2r
UIwDExDhoNM/JHKBTwefE5WxU+/XddPaBNsHugqbf9sFeqMhb8sMU2rysrCB+gKT
hPY+ZMIv8C5i79vWm6ZaVLqGA48ZdngE5CieINoX5PGR5lKsbJifgsUTh/cTt65c
zxvsNfzerxyHC324ZzdSaxPb9GZWGCOy20ZJ9VMNNYSFfFfFlWhvx7MnjaZ0XqBK
DB5d30NTTxrdk7onIfiRu7YZ3luzNtVlseQ8gZrsSupHJenXEPJGRswsicoI+azo
7VeErszQJ/zt89h4ddvD8455j7IbbUZ2hHIDwIYNv36lAQfKKWxtzYfjIe1q0OA0
e4vL3viiQ6NYRmM7F7Hqgrbw9pE2Tu33P+bXCLJplk8ZaXVIcCnEI270Te5sZYTV
GjzZhuDtuzoWZUWYW1cMPxXlenH2mAKls0XnDGHCt1p2XGRaFFxv79J3MO1fPBoh
B3sUnbJ2SCi1g+pzogBHWmYqC0IAIVXHGr+O+OWZv1rs2YH8eoBS2EdM5/AwzKbB
KQxfDhHRmGmp2iEXjPOfJm1PMbDQJ0I5IcG8os1IZRIebM7zjVEWw6//1XIE8LIn
EXYaAgEQeBBLya+4XLuW2xD4T5SthPbn7Mc1scXIzmcDUttMcIa4UuJVmcOTHbLY
B6CPPXi+0708vgw8sC8REULSaxGwJycqsEQkEPEhESfOcqq2LKR/YDYcL1Dsa/Ac
cIE+woxdSpwO7NR1vOpx8/jn2SYf/ETC2JW5xziMMm1cZ9N5viU9tj7b58k2LN3+
MSUJJw6zs3Rqlk66//yzv6w8f9WarWxljvHXrviRSnfeMySc6zfsWpquZcBluWo9
rLOeA3gvWNY0396q3npdOJzbaX5z31i1MZBULSPPC49O861B9v1ZfOEjn7JjAYHT
JMp6CZDP4Cdr+Ahdyedk46ZdOCCnuqFVXbQ9JKcUHNGtfI7pjY10tfyejdb3SuIp
cGyfIIzSF8hUS0Se/7kLp9RqBJC0g8oM/Xc4pLbbFVyUyjBAf/8APKIOznRqiV71
c5aLN5h4K43BqEZE8xckgbrkMc38wIz0jxvDSqqkorGia+74r6AAo715VlXOh70G
YodYBMOffRj9yU8oMayunvlG5YuBwUJ6ygapkkfhfZgj0TB+raTwhk0/EYeGSX+T
dhnhKS40HgXWyLbBItbKJLKCg9+2Nd7H71MT1Zi2hFDeYYcp/vLDs87G6P3nxs7J
sS+swsBy2iu/MC0k+isZkZ86ZvX8hMNmR5cionJ11KVzleWjMkiDHZEN8mG6A64q
6RZsxVUPWcGAWjn+IMYjsiEiUyZWdeVAcFTeFEk4gJCCzdiliqaJLojKabAPt0sW
fOZ+YUXmD1hPS1czyq+ipTGrujo2VNeq2fU4hiWitA1XicA3OrpPxgQcZ2OO8DQD
PKZ98+b3jny2AQEKmt0HT4dUuwINeVqQM1je6d+vP1+qd/gVV6oivBRwd/lhvaNA
dOw6+wnhpLsXKSIQu4/u0XIGsYOAcez3onQn/wkLKx2UXKz1m/2DDa97C5AvZYLu
0KHuTYFVPYYdaOja9hYTXD1E46NWHfRvbZmypxuqIi9xYUMMba22Dfb+msbECKCf
mLQ0If1gYx6RaVVWQlNobFIHab5cTQvIi7wq/VC8nxyPeG+NyLKXJNimh9z8rau6
1ZTCW63epDIeoR0ZY8oieVy+rP6BgQvfPsByPd2P3mjyzz4HbhcuwgbIaQI4a4+h
jwDajOKfdVScLJR9f9KOesR+g2nusb54sfBlUn+w/3zw1AmTwNKDOkbWdkDjEpy+
RbJczcHuhJszENMcBQFFGSvkr/d5fLMg66G1f8YXtoJGgBE3XzysW+sKIMBT+XP0
UdZpBLS8nVhlmtgX3jzYtrk9jMRtBiPiyRgckSo400D+8k5NVzbjziswjkBzUTe6
VEllJb4jlPGsFf3hZV/RNLECv+S+bPMLrGY9FSTnLwq21ssBjNgSoKKDjM43TMWC
tqPTrBwF+sWQ2pyab8LpMXsBisG2xi84ygOr0PbAqcH69Pad1mUKTHFcQ5otVic2
i6S+LunNvmByhhqHfYwm9i5FACt83Bf8xWSMOI6+MW3md5gJgx1Q9NdhXmlO9TKN
/CLJcEbkTpQ4QwGVWBV8caAoNv33p9+y5zfyDPcEF8SbQjkpnR3SVFK8P/kN5BKE
8vWf569keu0IVynsDEt15BLv90+mWVZVnn2/5MQjjG1Lj9fBW220Ww/AALVjX72U
A4BEaJkceB94Ee2aO54ro1DZzcz1FSHNozgwsTB+bPqHYIyA+ODXbIwQq/lNxzAy
a4R7Oor/8E+CWs8pc1ze5DIze8JJeLvlzmJvBfIhRpLipHly7iUSYVTTfMaO1vzO
aJ5ahw14QuHB1VGJoHURYyMehYYd1LsTt9yKRZIthiKLI8TqCXvaLXU7DHNXZyfN
vdYxO6VwGsH87UvFbZNPReEwkY8ar/wlpcKgV6T0g5hhunY12yBuSL3+ei/1daCq
Ijfe26Av70xey5DJRYE3IFWKNWRyJBMcYMGbVVk+G5qHgLTaCVgiK28Ru+Xi9pa8
EhOe7ppAS+vFPNjWYAgVwuhyOJIQIvMGCEV1nP6/2X9/szYxtD51aFOmPCDeHQfk
vGFBAYh8b7E1CwRrDyXBlO70niw/RWkrKFOz86ynzcrqyQ8Zf/jusWS47tqxS97D
MB2wPndmJPFIdea5UJO+ZEWGatB2W4D+0Yt4UKcb+Vs/Bl0NJM0eaOw4PUznjRPJ
vEpRjcX06cFlcewCX3cEaSanka0JOH/rWiH73j/j9y8eZs9vJX8lskNS7kQfQ/ei
EBNNQDAp3pxsDM10zL1QnaF1S1z92DpY9qBDlyzVrA2G8Pj1HnXghDl1ergzMbum
mx0Pgt96PqBGbQGlT8ta/qqbsBEqbAHeNUckuD3Zqk/3/1lH4MeNzDmclq4UAYV8
3yfCo3u0DdccRHS8Chbmjm7YjlJQjBSDgcfhx8KMBfoYk5DPKzaAzwIpN5zHqr+m
C9pwR96XHVRnmnvD2387SxfKT1YD5htBlluW+Tp0mppowiyFtNjXtYB6dDiqZgHa
cN8MpJ84tbNuUZJCmTVOIKt3LmEOtaY9yX4OupjEyn2pQ0WJNmG30Jduko5rzCwg
ZAuAFpsqUMF9oGlkQlvk0sIqke0w+AQzBYy/ISa/9O03F85somaYi55K/zS+ubfo
VHx4Nl8/iUwg0+Vg/tKxq34VrC3YVMjiAPuLgwnaa2t1hm7abaZVOZjoGj2cvwZS
N2iw+g9AERu4+dHEvzhgXfxunxSODgPhAqCJj47DL+N7J2qX57NfV45aB4fUHyz6
MooCEqBFtT+mvxhj1u7azcKgPhhG5PuoHJjRXcyqINNpIbYn7y/MebQzMuwM0c1D
bkj+Pzk5La5OgzOfM5tNEBTCxg9tmep8BCx4Fli4nWXuhzbM3KImHzlueDxb2hMt
ZSuYM/Wg0MBSY6k2ZmZzu/3QT4P/3SmhDJoHwCWMChiDqfzitCXl7eIKWUQ3Td5E
BWc7bLJC2suh/q/3T+vCslxU+VzBFhsZPBOpuw5xnA7udF4Uob30LPKUSp4vvopd
87Rhf7vm9mJYgIi5DB/yEcXLBihPnODMMFjj4zBxnkE5TirHJI4dVnWR2hRm5bdl
79zSqZASVFzkGreZGcXgfp+C7wF2hScq1/tkMFDRQPGa9X/bdFrLzY+wPdQCg88m
YOY2NTjiedPyCnr6lXGN+dEcnkEyLa6TwaBo3tK3rD9qBvSRlS93OFF0c18Ymwb/
QwZyiijeGXS/CBBmftA0RsqS+ofMLQArHi3O5UystEMCz+IByEo2bMOaK2zJEx3u
xoNob5pmXtcXpMEvTySYc64F2Whtf0m0aD4JpEm/mqJD99ar9UhqihTQ9JLzJGsu
BOlCCI7ITvHiEdNHhMY3TRh8idwRc8yUY9bwCTdUGmDmbnJnTUe/5MFgrYVuZm71
REx/GNUgBeMnSTgLU3D57EAxKjXNUj7NVjDGOOrT7dZwTaxQ/gmplzjvQKAjKudX
xkQ/Bpsdnig3AMlZ1nrBTcJdvuRSOXZJs1TlinCB+ZVJinDoKJat0qpFyUbe4Jwk
oCIfHqBaf6Withdk7UdKpYFibkbr2QfYGR6oqdHPa2WmtN2eZpzU7U8n5sXryITL
5IND1b47ApKGQ5nQq1rJ8blhzg7BklZT0E+aUYFzaeN7UWsNYtpSx2PgNuc2tQtM
ytsNRgpvceORKuv/XOYiyjvq0gCb3bC6c8H07DWTrtwNXQjvxyF23uYbcWU6TQ3p
QksrcLMWepBCdplxCxcah6kOE3C9FlBaGIIbHgPSJRO3XSG+vBU+pWzD9LxIkwxp
bYO2fGVNBJJPsOoYFB/yfJnfZ2kEs5XBDBBRafgD4fUOEg68mLLK44hWQMGEpUCE
P56TsAduitaQEbYvaIoGxawduVM5K44L0fBkgSUYxHxkl/3aPMxxk8iTREkUIzSc
5FywfS1nibKl+5go1Zq/aRW/sRxJGTcXINuhcK7Py8ynw5twGKLEN8iJ++emNVrD
+YVU8N5AoMF9WaIiUHCnpWZaSu3pJcXDDooRuUz8o8azs+sCXHJ3wcDF/SpokZKb
QVEPhwoGeVHynfiGzB31lYme4WsY2HaOYbdhZy5y1sl9dtSybyJwVkNcOGr/03ws
gdhrMG9VUQSoCrsqiWDFD1RhgPFS9nlbjoXfxRlW9tWIGT/xv8pbapZp+/R8TOLz
VFEz/HzG9+dUzFtm1c9EM9QMs3lrcrag3N4MBUbR+XJ21DQjlC2IyxAfQN9YfDkc
CUGNEx4m/bjiSVqDa3KkPkZknOx1sHdVnEB03H/Ko/rssIINNOnzmch81e8a6ZjZ
gfULy8YqEoZPgxCbHKlIcheAr0cq32UZAYcEXbq7XHZErsgSpoGIYzsNmxpzbmJu
0kWRMca6GjC556MlsUAuk3OFOXPeBQmPPB1Li6qyJvLCFoHWrWUWNeQlt/5LNraG
UAoLrHexF0R5u69YYc6cV+JbGuoC3gbfolIxBaWr/6EdrzWcNJjrOJWu5Pzdp0F3
wA+2l5pCntAq/LiAQgOAehN+PSWb0px8OWfeOMZRcrV6uqIqLHJWFIa1intOE7xw
FTSy200m8cNxoJvvVM1rXN/+pKx25nVbPi+O/pbnXo1p9NVajmKLA8ItoxXo9eIT
/mWRwFs0Z+sftCCbc1V9W94QmITpL8Z87FrwKYuOQkFNAJQ8e3l1NvSmKwCMFX74
7xh8+VImUnd7R+xa4/couotwCFWNW9lbxnBPVp8MVCgn2c7gT58q7MjgZWE38PcR
hV3BAZLAxNQzbyc7rIH9YvaJwjJBstMhNWV2HHdd15AEdbBXabfCscHS1qBsN/Cy
kTVROByagzk4RXUHv04wMK3K4z/ZWlAYFvv3mSpSj7jCavLrP36Wn3V2jGEP8R48
dt8eDhxFRxPyayxdd/AvGZtu7sjBOpNHjCu2gGEuTtrxCxK8U1XxsVLflxdEJK/w
x2ZnWGCmh7V0kXYxKIdhIEYgeJAyZbJwpB6fjp2TOcv8CA6Rgo6193lMFGi2XcwO
jKjPERAH9Fbu9nXK3FkC4GMZ7QLjzWFImIQgNh9FJJ2sEEg2M/sVhPnxuJpzOs83
CJVWGU8a0EA9HhMSmcoleNZLu8ovGptRRmAyA+WXFn/EuNQfle1yJaIMjp5Gyoei
O2pi9V+zSrRQkPC70IcItCYEJquy08+KVSwuvzF8r3VO2HEwkHnjEDmFiuV82s02
X7gKSfc1Gw8kKQwKwKAiQKGtRxQxWEyPmMP2trrapuLt3TqnPoSD3VB3grCVI66Z
UMVFCRL7YY15hszy16Yn/pvV1S5bK0h0aEk3kiJ/ss8AYUU2kl78NqPDLw95c2o4
xABB0o/N59diJJjW885jISRDF0xjjfDy6Rtr++x5P2atqjwhUK2fbayVwzrB9g6/
MlIScpwmTV1738kjuf1yt+bEJO1afU4iEXO17vu8qtAbeNPqNiv4FM4nn6StYAe+
54q+ykOJjaVIxMNKOK+YeqGNE7CHbBmRn26n25kwvULmtazOZG7w2R0x9o4eL10E
yqs8Sz9TmyM0cYB7rPVxOL4J/NujoDjSizsvsoXJqXHpRUP8KcEEewb+hA1eUqTw
zxYI9qdNbULwcwodiCWwP1qPdO8h/Vn425COonCLqbOSzze6vMjVF8g8Jjv8NhFH
HG5kBga/nXJ20uJ0lsiWYiPmAC3Lr46wi+jiU2TAXC1kU+HmCWCf5osAg9GuVjKQ
m+Lt68/KpIH0K6Cr/zWARuTWkja+gm/BRuTTs7UdjWxhQMA3CvTD8U/YB2dQk64q
Q/JBtp6QMZDBHRbYsI75uVZtmmA5K5tE3fMazBazYlm7TAdRVpdtGECZxUdgaB61
zFdY1YtrGtoIYRqsaRWducyMfhwfd0bdJRXBblhXODGaILtr6+gyvy51IaXe37Fy
txBbkf87eudh+nbDF8XqMcP6vyxHauqaLBS5skP9sPP3ZlERa+y9MEDEJycaPqUU
/ph9e38cBem7m8vBwiMNgwdD4j5OumTCGKFCOcHFiF+3HLIP48Jn2aRSvmBVq1vE
ioOBCddKbhavG5dywjGrb9+cIsiDmNya8HxEvcPKbORr03TOz7eG1J1Bndmvgi7Z
nHRmkvuMizZcMb1FoArdgCKQ00oAczf77RUW22yqeD2pmZlzh72nLzDNlimu+CRk
mVwtQbfD/mlOHOsRBPXPkOFE9ccAd3OEadN1PqL2uppPHFfSpL4fBCyjM/bVaw/w
1o//vSIG8LXXgFc/MM2jFxe0Zizlb3Ep6rwEv3Xv4b/nytJjKU2MIZZPg8i2zo/T
BgkK3UqKRzUIo9nOOogwG2MF3ncgSOUyCD0RGccxpeaxaqhYCppu792zIqXSxGay
dpeJtL7JPZy0Hn2MOkDUQfnqAcVxt0NC0sWpbNdkC6aH6PxNTv6GZqsN8ijbS1FZ
BTFxgbA50MowXxUotgsOoGBR9Hmp+1nvS66ZFWO94Lw88R3vm3uJGQO+8sKC7FWN
l55HzlW4QsWsYrSaM8Bd0LONAPJREoShIZg4pEGlfGs6GxhrnHwkdC47OeotV12R
ajWwi+P4PxWxj5BoJHZr1sBz6kgu+FV9/RQN3re82EZWs0fgxY4hu0dgLENCm1Ro
MUN16brKJpgzZL1uLVb/njwBFx5QVomioQUXDPRtZ8Z4mLX9yINYnfS2PIfa4cK+
FXFHAZLPOS2TGbYsoHrbni0pn9v9Tc9Fmf/lz3pX9BF+IegxKQkjXQgoU9bHcxMs
DYmg1yZR0jjVK0nwi6/HwH7vEGka71jP/yDwvmMBxgP4rpMw/Ba7wroE0LSW6lrT
zyZSTk0Kdi2iE7oNw9kXL+5TSrvFR/AdXmfMivJgD/kTq9mpJFoOEnyPR57vHKpb
yrGMLS2+LO1hw9y0DIg3DpO0j4S0iIdHOArKqSufvEp1J0EwcQ857JTagtXs9t2L
A1+bbxrOVi3jggwQsUOT0WYfGUJhnxHf9f6y+BZaxIrFJj1WYFlQCaTKMFfhEBUF
nDIsbaftgTA6FijC1YZAzfz+YSSMTor3mqZ9CBBtiBmr+pFcP2cKBeohKd9tfPqd
XYJ7sD+/pQX3md9JUNASZ2peiDV09rssAdEqXj67w514ks69N15IufR6gifjENz1
Oi/SYU15yyu2WeLWZCP7r8U9THLX1rgyTsfe6+1oWcMRPXl++pbJmNm5od2zVTL1
GQJ2xPH3mzecEUWtTZ2IpoBAjtN5H3WglNTT7wsCmkguF81daKAAO5kxGu8clPNT
fgeCZ+7sBU0Quk0AlK7FpZk3VFz7HtAdT8upHP+K3co9SnSYURfdzwOrsupjQTd3
MCZAPvXQiGGNdSptQpgvK0RHtLrwOTVS2jaDNcglik9nhfJpHl71IH4in1fYs7Zu
Wgtdi3n/M91wNuDd1XzHUDallxxPLisdpPXY2wCAlRqG35KdanQToLy7wcqSCfWL
woEzZddvdm/KmjF2jfHrgDKV2zbiYAflirYLDzMQxg1A6bcwZDlo+y6kR6g7/uTp
E75bhQgBRYDIvOx5LF0t2LhR9NAlRHB84eLHTULK5DGgKkIGFnCWV+RgKiM2D3VC
zV17SMTYT/xqGy+LmOKX4IQmFw7Pl8Uo3Z7ZlWxzhp1i1gpsiAkxREdNJaG/V9bP
gFbPlG3cjsFn5gEqtI2uq1HxVkCOiIgz7LjvjMqoaFHS8n9X2AuLB8GERlCGAtc+
MbXytAOxqqQsahwcfQiZXeshwEKITQqJTzh3ttIDfI829yLsY7qAGw77Wc4P6/v7
b9c3z9ROYY8umppvndJtVL869h5iOro4drqGSQ/mmyuG9lQJstM28cb7mT/Imh02
6DhKAObQPmLEnOONau3tXcRVKduFnd2Gnt0rYqEOoeuLRNysdM/3LZBMBOSxBML7
GBXdnrgni+oUFY0PowNmCquaqW5lgBupBDWmqVSHzC4lrCT3S0MmMZV5cDB1fNpb
0YLddR2f9PfHtdniL6dsWXaUQf4gcGgcMPaNpqqOikxWzE4UnjT/s01SV7/DQWGa
SkBVCS9WvlmdsQwyCnr7mayn0RR4ddRObQpl+YuYj/eSwSfxumHztD/idrQI3j82
Sckaz10TWLCgE4OKGhVSBcramVyb/Es1crDBvMatPcPHw0qgyWA5Arl9EYnY20Pa
tq4rqaOqkzy9+tEBy/oBIhaqzh+u9LgpCdVjZFCtybaikw43IPx5wTBUSj/3/T3j
EC8MaXlZd0mkCNhM93oV80mPRgBinN5qa04j5txnaoEDogxPc/qoEkL+oF7fYcMq
/BHHXSakEAIsZ7G3Tg5ZqLM+3qBeXJb2E2Je3R9F/iIEUV4yl7Qr2dh0VXo+cJfh
gFz/y8YLgrZ8hHYdWviXo/Dhqvi85SY4x58RnaSkkVG0OjIAkQBCCcOeYfqotWlz
iDLaezN25icnGIU/EDPPKmtmlg+QoFELT/JdR9cBU27ccD9D+A121I0xt+28435A
srhpja/m1hU+7M2Jfcqos/qyhFqwXkxpegJCf33kQZoLJuymdP/Gj0rQci2FxX4L
5CwXQxCb22HsOimchSkcL8jVerfsr/61CORNFm9UUOQOYUc6txREjZNjVEi81gR7
HZ15Cphr34p7xyC6NHcxbHOCHEx+7As37k7agGiPkQ0nZQ23d9PTZHZh/ShzbTh1
wvyphEZXsno5bgktq3p9nBdVDkTA6NcmZS7PSpOMUOj991a9sfSJBySfnwkjqrzD
EcAGUIKA//Hyl9OvyITAGVlmNhyHoHq+4yvmfDh+C8tHIKSkDHK6xaNNXzLqb+Pl
kli4FNGRWXiiQ1p8ObYAqfiOQbvAfdrlGus/Kese45C6UwA19KoUIKMuDSADKFx1
h2oNQxwlmYxFT3CTFY6/h/h/2/mxTCm/4jY71uNQNT2WICIeDuw+2fB+tB8sYtIy
0XB66ANoxw1dxCaB6JpieVQL3V5TNeg7kgCC6BEa5oULGYaMJE0+2pn4Qr0UkxnS
8CYvtzuaTa0WVfjBmDoJhEWOui5+X3A50jUDzmLnKYhkG4UJInKJ8ReiobW6NaCE
RuG1ANyfr2C9j92qP8zkCIS4x9EBJGn252HF4R4bXo83bhpEsd+Azl2bKyw+x+z3
H1EGtUFdIlHRY2+sC42sfadf/sf2UvXk7tMch1aU/EgXIzLN871WRB6E9IFPHYF6
nL3S5AGHn8eaU80WiBDmVIznIHd4o4lsc9xCYOFWAf3mJXZ14NxR5QpGSLs18RL6
jebtW1wmCVgs7wcdmoT0m8IXirI6YJl4m12geNdRXfFwf3O7llNO0pVlyWsIhDkU
gdzp8tdI1gHI2kMi6edUY/YxVKwoZDX7K+ZggMNvnm+bNgLHuI6hAIsO9DTFnqsW
gU7U3sO0Y0JpeZylw7pK5+n8mJwKL3WBWlzmgkS8Toiquu8dpNhQ/8Ywiq43BsY/
sYH2I9XxiD83yMb4xeAljBTH+QlMOuTmA7JPKOby84msp99l8vyYdLM9M9W2OXtX
f3IWURVeHhlEUk8gFQ2icau0HL2vQS9lbEbtjP4KZKag9kuF2OCeCSA5HfD9BgYB
thXiLwVSGT4VKHveEDV8dmGK36QO0D3IgzpFFDG5mryzg0ILYFJEbn7/6FnZ1fKt
n/X3V9w9cLBEkD1pxb3GHXgI1W3zjhu/WEYJ0e7n8AiWhthoP1LCnKxcZd8dChQC
H9agcXRkajkfPlgD54k1uVw8wJJ1WL59tov8OVBEtFUlq0sYABn6fEOCqxoY0J3u
N3tsDGVzpUaWHYVsoGiQ7XkO5CwgvPIoGf8ZdgIuowgdulzFkRvqzd/Et1Fk4Yw7
hKztsPRjTewL6EfodU1vjMunv4qxsraNX4Z7lLQjoQ7eGEmodQuAoCqsm4J9IS5C
J0t9279QWlMYH9VyI5IRph2mI4ut9xZWiWQWPxNGzgiUDIhqS2JZplrHN9yOKuER
QZvRtv8auI0ac6UmKmv/SMUGVZlCDbevjrt08yJx4giBjWvtHj5oipNPzHHHIP7M
vumjWD4Ur7JrEZSnlYpBWEPmWE3Ti62mDo0Fi3Mnws+XYTGJyRXyi567kDV5oAQl
fApHCUf8rNfPQEElf+yt98xVw/MU311fQiZ7BapXy5Ap4Dfw/NeUK2UlqSTVW84m
cUzN+gqokC6fKKHoQtcGXMbPcun87bSqvi3Co1/SSf/aiVu4tv9KyIn058cgpodJ
2UqrLEkIx+Xtb9zDQQaKy2vX4MkwLg2L49/OvK+zz4FAN9P+YR1jJHmOMnv9wo9k
41WPAlqSIgpT4v4WL+8UsMH+7yk6tSDIo7rS/gaWocmiJvqN5zUAPh1dd6CZ+Q/H
ANg8M16a0UhtJTl2fF6zoR6bjY6NZlPjQuxhCfiHGK+E+H/5rMtRzYH0wGvh+OGO
jtFKenPOuUobcORGQZDDyOmdejBlWJOx8dLKDNL1wpU5nCHIclNRnysQWT6pCm0P
0pLXPIyMfyXdkBTo1Y0WLbtSnUiVxBrNpUXC0H9OKh1pihLQNEPjTcniQ608Gh/H
Zk3RtIqQduTaPP+nXUe4zhJm2qtXz1gY89QXQ9Vp5Eii8m146nvrZfbIPPmRo1L8
aEBYy+fUbq7Zm3ilndQHoBuaoLuVj2S0ncG9yNen1iB80zoh4re/fcCiJEuwW655
EdOCjnTtJXenoVpfNtuliUFT0QjyX5tsCBDo+AbpgnXGzlEc8XY+AOG24u/GFcgR
KqgfjUTz+uvRQugqxzAiBK3CIcHLXyjeCmhaOAmRa0u9rnaoxt5jcbeEGV0Fiwfc
G9WueGTcrhcZ9iGl5AzcjABBmXY4lVCd26fHoN8DnDhpV4iPd3ViBaByQrGORJZh
mYQXM3XdM2tL7xE2VeSDbC+B/XCQf/eica+F3ZnIMs2tUuzcTBRRZsARuC0vLVYO
L2Eb2p8bFKmjP7iYFW36X6jnmzD5ICFiAuPMCc4dLiXI7LQrzNc8nTcVIHQU+3TX
fjCWpA4mIxPLtf3iuLyVIFBaV2pLTFYrVAe7TzCHAd+nxFp+OHIRgYd2SVKR2f2D
LxzT8oOVQeVuGZQtzkmun+bKmdAM8fBQIjyzIGE+a0Z+VHIbQTDStqVbD6VB/bOV
gWIWBsAcR1zXY2n8akle7gmR2mu5cvBH93i3n6vDQcLlm+R85CQ07bAAzMzqO7aY
cHQ/cAfJ0pe4uMEkh1mVwsBaHXJwh1fLNJ49ku3WeK8AcT+t7SiDL5OKXlcwAPdp
YB9pjOxbLniLjBrLiEeHb6LO3i7xoUOtFTUCul3rYsyYjG39QOq/NGPlaXHq+xJx
FkemijsUqqdK0qMpIByaxRk13sZQBHEwaWEwUbmWdO+LHdok57IjZTBppwj5LKOr
0I1Wbj0b9eeI74+iFc9rzbGd6YoIC+a+WDdupXrq48JJUGcYP882udb/o0fp7OG1
23udlkx/P8Od6gAebLcbdnUMj/YJbvsAN+aTyXzm8kAQAYb+FFvloo0zauP7ZZ8z
wVOOGqjdPSQRJZlQbuk37e/MzRum15Em2LCiBqbcBBsUPVfUXVDIlmD95XwjlCdG
b6UcNKT8oVcs1y4/DsRGfD4FDnt2GT/9fa8SCRbWi35vJPDJ7SPlZq2G0PsdugnU
jSUTWVVfDuNwKr+XjLaBGettyVZL5c/BULrctHkLyt0j85w3Q59X9NtPrdHr9AG/
/e4G/K46gKzYfe3vSKexR+ExFT3LO6mabTxPVWC7Dg8A4zUGmOW28EnUcMTzEsW5
fj5b3YVzx4VECiirR62uXlAfDn8aGlAMo8DaFpXMRp1peZDmiqWvM6uKCzVv6+VU
Q6A8NMu1a5pmjkfsMGhY/uZSqElUKFPTkVsF+YNL8oF2S+3rrVOAlzfHS8CMj8ST
a1Iwpkwg/YYE0oY6PitpClRJoPOmZQJOG1y91D1Zsx375G3cygidkS9he0PJUeUJ
f5yDzYzRuijzBTklzfhvmC3EdBZhiMYVzPvfX+1xhge+gNsBNfp1fMKTkV/JMdq7
o/4zrAVShte5bPNbxQEbzvW5Wi1IXES4CHYYiieSVPuwTydc2KVmimeRXQSkCchR
98y4dsbpM9Kzek1FphNwK1f+XauvrtEW3S/sQbr+DcokVqnndggzm2jQhgQ+4Ukr
sQDywqKkH1EGu/aE37nFPHH1Q/onUobkPtb308U1IpFvI9acKZCTiccIeawmVdOZ
BhTfUjrNJc9/ixPSubG0IoGEi28qZP6jqK+QWrOi5sZUVQ8/Q7tVO/0vDZeSStlb
OcKqYs4H9LnCWRVm5RES/sSnSsWUgNbnA1L6LfzkMGWXFhCNkAD7rVVecXtm12eb
GMUFeIc86osKv1g0yqlinWEtIrrNfCNdtiElU7YZVK15jd3hzkJaoZi+g5WjaApX
8tJq6f2XWY/kbkUJMLOQoJ8GJgtlopUPRJPJ53T3Re83ifnpDQ53BhQvWGnBgIxQ
Z1zWYXoXy7hDlx8X92AjYzOxII5lCwEBPINObc/EKHCe6LdanTvA7b5D+P7+Bis0
3gDyK9VRRN0Fy9uyGH6xvEjaYjUtXeOTzXp6O4UP/nbmvJr+/UuEhTOpkoS00nBi
bJDb0+N3hSDNzwjOU9BodqeAg2b8Yk9kW85UOOLDKQ4PZ7T8q+j+eWktF9cTAk0V
ews58etVYVUus5V9LK8cxy4GEhAe9tN9x01iRUAQVgZQvvtLevmpTAx18syy3DlJ
E41Jku4luxbTkVNbl/dVF6RYFum7rJNoKMJ45vQSl/wmcbkaoxt5iK2OEMq1cflx
+LgIzWcyNAoQwHGOLqulATgCKujIu3MsmZ8Xh5u27FnSElOHAUdan6jUUVW3ry/8
Q+Wxf6oPMFQgaD4skXx+tQPUGsSL/wkhKUnPNBqNxcCUgz0Pl3XOt1P74gH8vkfr
9VUuF6uT/aG5stbjF+cP4+R9TQh4kBkopIuqs6GQTaKrD5fQ127lDrp2TH8w1RK/
BVkJGryJyNLMEkM9dcaC6KuMB3tnnIArj1cdHE5BUecqescPYxksx04FcxRrMh2T
9DzFbtSav9fQ5EsHcVz0/3B+8ABS17PDjxd0MbTyv4M2WuLmLBzAJDJFDQtOt3kC
4eQGT8ZMoml5X+oYypxDxvoGdFtBqTaaYKZtRaHYDG+W+2EhF52z+aR3lbC/ntqW
ov5rH5zohMX6Eoxjfw/mv4s0XB61PoJFQNMktYoXj8q6o87nKxXldQbXqaEhGmNl
neq0omxvgdUWrDdQJ12qzqam1V6eYQtL4s/Zmd7mU3XwxVOs4hzikK0j/laMZJL+
1IVUEwXGRYupU1TSk8HtqBs6+PZtLqU915t3kWiiip6ICUdFhO1y0kRymGhuRfcN
AFuUBwt0CApAM4UJLDQSSbUVFiAX9b4w3KK+kQ1/f2H5PQ/CMcvwvK1ezCE93Fba
FNS+VxCRHvOKVpPJ+V0ZdILS5zPZptiqg7Z/kZivcIAI8gFtoY0SAz4/uUpOqeGl
k8skKdzwKvSlsz0tFrRJVDY+ycmwO8rM2/E+Umw3hSRxjxvrmpL6tpfUSyVtOoZ4
5ftvoKA2CWqkhZNTmvS+qqDFFkEZO35qCUZNywtj9A6z+bdUFpWYJDqKI1Kurwnk
Elb2/CaYEQkjOgcJOX5wmXFwiMY0U+pkeKcGq2zj/2tvXJqaG5MbPvTCaDxGZfTJ
y88UI6gUpZ0VFbAxSt5z7vmoesRs8G/hFZKRZ4rbmnmjgNQTjcqZhfTb4JI94ux0
e2cirNHxmClFFp6YYkm+dXTTIc/J/2Wa7opZDk9KzESwEnKruwKdgs2C8HRhhWoZ
q7kstmqhI3Y7SAViRqr+s70N6IFjwmuz6DStkjPRIk2W9sVA4+K4wXfnL+99Vfm2
WKx5yHi8doDKQTaC3crsa15zZyiJKGsZkABtegBF9V4+cr1oF+5wdKWkzMYeYf8N
WHJcaG4jz9p672jf7cwCx9/mv2dddMeqSNth/usZ43QFk6JxLglZ4hWu75aebT7m
jiaVrq6XGyHi4FGCKuarrZewESp6FWlovDmi0u6v6ifhogtq+elZSH+GoDYFl2Ek
u+pJHAfSKHvCjkQDlSpij56FDvevSvWuJq433ak0CXcmfy+CAxIw6O5UiJ4y26lq
h0DLMCV5LpXNF4ex4V9JNRdzQcsaMoOVH+HyvANQ6vxENyY+qLqMEyB5g7nv2j3N
qdzZU6hf2qZTe6/UedDeuZbakUvlQxQPJ05gvfLtbi2R2AhJ6baPBnvBoVMQfA5J
dXNtUyKzQnBn21tSU3j7zUqMGV2a4Ys1ApITEVpM2xVJxqGEV+slIevAPucOqdTB
PYd0DY++J2DMTuEMdbNeLJisAzH64s7vzQAe4TqdVb7WhlZOAPBayrchLfWx4T4W
YlDONSuEczsnGUopVfmC3hdwCrNgke6QWNC/JdCYGPcDDeJWvcc2hbfCUwLg6DI1
PwvDPnD+ko0tpeo/DRq7yC0C3nSE6BWZELVwVQD4edqBLWPlpVbnRqaH9xEkanCR
N0hLvNge+wg5OMM4xnWsDs/LH+R8KOCM+ThruvewFTFifjLc63VbyWtTAsJzUi0N
oSpRxOZgPlyuoIgH/WV6DHJeHq607mSU1UwX6QHZDPyTjWK7Z2QJqYntdxoaUAeZ
wBCqIHe8L12tijOAIr6EIvJkPUzF9u3ZUZqL7+4YSah4BHs0Rc7VF6lHguNyMVeE
HPtay0cidZMDfkbV4ORy0mUXoz4XshA6aw+YHAMdBerIGpAwwFT2W0XTxhOxTxlN
pmZZKluLnIs6Gi6KkGlhYg+KXAiwGhtYxhUoNwD9dlsp4hujfhNBGuihfOM+yvQ0
ljJ6jl4SU3sC/dHVh/kj0Pgkcb5Z6X2YC/Kb5gEGshFSv+zafti8LvljPDs1w/Tn
jZe1NhfnGdyNTOKZ/ocvy+3a/A1rryhzoSRRMONnfQHEA0a5qb1rciZyjYA0Vdnm
gi6zuYpaATpCyPcjHKqjl7JaD3UYvBO5whJzBIivPkeVUdMXcxA1cdqsIuuc+y1J
eLlCIL1ssgnVLR1jg9tJ5CUgFNNErKXODP00bTh18TW90r4HrekIpscuM0hy9F8x
dpbfezwotg5FCdd84xwaGf1YXkDAXaExh89sTx/bGj1B99dwlJij8nxWsNoEXaGm
niAkGEnPEZvxBiGM9xH4b6pFrtgOKvLNjJrWrDcsyLb9ipbbhfgzGCtDu9rFBPhq
ohw8/QRX1J6vyOXgIJlNHg2b7ce+wX7l58gLgFKRD/oxzkvaZvep7WLMtyOQZ8bp
hh+s7xtoBpgC7SbvwKq/sQ+UPLSNm6QO3YLUxAzZ0QT/iNLjS7Vw6nHxgIyS1Duc
27CZrwUp5Oxtpeo9rZq+iXGL38T0X8BcUo53NMzJmiZmcdUJKBjR6/YxJUODN9dO
plz2JJrqBWBXpqY9oll9EA5Mfi2tUBgomc5AQJA8iyt9XcTXdo7fgqHoAOp+95Cd
IxKF3kmTiH+6isP4I+sfzfpExNYrzQYKyhX/A5gmZD40sCvvp/ENZpbRLdGom9a4
S9z53HXET3veTxl9Z6iXr0DrEFLK2RcBEHjjFzxnYoOdVafjAEkIgKL4eoSirULE
GYnWb9mBf3/ytBfvJVB0P81XKConeeQpyGXeunFaYIekbl61ljY8/E0fS4DxxnmM
zJ1v7XU4ueYHwUFoDifA1cU9NgLAP02r+JRv7fzJUG1X04cXLSPeY0Q6jwhbLmLc
MX/9Fnf8yRbP5LE10ImCMxWqOIRUJMAzkES6fFe7QYpXOrOFQUrnhXTU+N8rXBIe
4rFaj5Aq2GPO24PjMHwssaYc9TDPO8HX9kayxWGRSKEWRKyuz67jmR+S1uELHNIb
szc/GAB5RcezdIYuf1f+3TZtSSaMcuQUfRDG9AgTsPA1OsZ3Ts0T9KHsYy19vwBZ
G9ZSvzx/jVXdnLYVoW+RyBp07AO1cCeseoVV+ZXGNW4dF7kiVQ3jr8XAaJLJjU0U
X46GhbmhIFh4e9zq19GINxB20DKopaglY0RyQLATSmhFIX0OBFYS9/fd6Xj3EdY5
jOdzY8rKkCWg9DT3Qwkpj1+GXshVcRS0//9kOpOJ7url6ZnxGZxlP7+wQzFlED86
8PPikQZU9JVk7xg5XRPw0joTDxDo2gJQqRQMKu71V3ONPGLEZ7jvaQ5tQKg4Rtmu
S2WN6ntvu/Bz2ovXJClbyBJwW9TrUjHwc70lfupeB7dzklymcwnEZ8vRpJrORDzI
x92tgqE8I+9tqGllOdZQkAron1tV+QaRx/Fd0Pg0tszMP89dlsLh15nGbrK4tPbA
WnVkR42F74zG1FMki7o6bhKYBKIW+P41TL/AT0VxakOiOdMuMgqzQTXjpFKLQEPl
+Bid9SKWvAjeSuyc1pAK2UkwMbkQ+604ZMxWzSbnN/VsakluSrchdyBWJEjERTOA
9N/MPCzv5Sidlu4ik5e6nyi+mwbsFKLIzddInPH/UJJgQ0+WV+8N+z7Pzrn4p14D
bdg/yA/uKHFTBWrXs3s/vWmcuOeO0Ejp1o5jKsS7nqu91YBf9Tsc5y28C9KHtEIh
gKb8loxM93hNwr6zW3LtfvBG6hNkr2DwGcfbU62bbzkvqZWNJJPRnineMw/4B2FH
Bqk0oLOfR4A5gV3YS+hqvGyoh93b5EDke0PYcE2AMDvj1++mJR6wy0mFiGb0RBsK
GI7KPI56R7H7n23RsdzFhKF+mWBeX/YkDEUmUTtq+zq6Y3iPXp4z8lDHHFV1zbtg
FRzHCeMLlCJ82HAqb+Ii+ZHu8kN3rIZgY6hpvKvNcBJ3e3x3S+oc08RwHNwHpuow
B04C/gOmlbkwcb07Xw4jNbMB4XPHxzRSHsrt4HxqyiUXN/B45tu1Q4E6OBFArwlL
gZGd4VBuQIQMxf9W7mv+vci6Y6dVvDPBmLaKqyP2K+mZz5+WWfGJ+/4DjihM6vi2
b+wdczYefdLpOuE7I5ee8LptUgj7AXGGh49RzNAbV2aD/vemR6sGhPf+frb/l7mA
RSV/fT9+YtyAeWSD77hh3ohTICxAI8SmPmLKd+K0i8Hbdo0sS/cm+FztU2M5qsu0
zQYCQ0Lp1fbI7Jrwbmc8uBsR0Q+dCqvME6oBe+Dl1pUUX0akfaGkq1jcaXmJB/yw
ciK0uCuj2hzWH0PNz3HDEmskWh2lj5ZY03zdCPwqceG94MS4k3aAThPBhwk6UTJG
Unefebv3lKHDCDVIs/fsoaju582CC5HJMGG0Z4NesdY8W2nKUCYVDOdaFi1eeImK
49IZSxkyPIDK8vulK8I20SNmJRhRw1LwaH9E+Mc/rDTJjJjqKQAZf6nBjdS6HT51
/18lX9wmFrxAJ6W4nIxNwT68hn0xwtTBhbFBW2eEYypnqhILfHhhcAY1cgA1Ggj2
5OoEtDm7hXw176wKPhWdwQe84zwY/FHBbzKP9yrOWtKHOArmaWR5SdkR2OBFWBlp
D+NtorW/LJEAvJbMgcr4JyHjKx29vmmQ2thrYElF81W66QMGbS7Ae0SUTpQrjf1s
M+3w+1gvnDMmEdErTQaueux0eOOW3+NTB1fF1IaJuiYF5omtrvZiw+aU0SVqhcAE
XE231bhBKtenRFdRgtmny1JOP4+f6tAUc8Mievje9zG1GI8Q/WIPa/lBQ4pOxDQK
7fuIzAq66H6Qmg6qvgQbsHbkJc1LWHGz/CondYJEhAe7OGmbCVPChBrU0L8jDZSJ
JtwJbnWdZBEG81cr1er5vvGw2nNX/nzQrJQxfPG7jQ8bMXOhkhbRtBkMe4MSTZXI
lC2XEyAv/vJsK1AgBL9YbMc16XXRxNkhpXfGuZDU9fjBaOb6aO4Sa84lGdfMbGPb
pkdnSakmD0uTGW5HvMb8HtE4jO87LOdhVwYF+4SzSK3fZm7CYS0lrhWIQQuAsAlT
+VGS2Y6ZVBCvXq2pMtHlhDSYMHjRWQrXI/9nmpnBUNYG73QSw/x+ksGY+MZH1HzW
YLha2wq/S6404Po+VsECr6orxR2DjE4GbeESnGJOx6htk1FbFBfWSO7ZWRwcBYhB
Pfva2P5ohqM6gBR/2GsIL9b8LRmQo5GCv9nDb7RvB+0fftUbMTY9+QNMV99IVPON
w6tAhPO2dz8Oq0AYTavOwsuG6wDim4+jbWpA7mEBI4V7ZrLvTgAO088fa/1szctj
egV+aUOXSIs5pmKzB/hnbvlV/oVVYCp3vZ5wkvaEyrNeX/dsA4pU05uRRzu0WqSq
FV932b8GpUbwHNNdjaIivprKUZG6wX5Hekm14wtxOUN9udyWHNvE+C0bR1SqHptu
j+keDny8+q+n2m00IcB+jK4ew7f6YPe/CUUKkN/l8bjJjhvZcq22OhSIc5TfQSto
321C+m8s2dnrkaF58GSBmZrhKUbgztMip+w2y8U59OQAmZR7Lydcr1hDu7L4DD9v
7DP2Zkrm5Rp8aPlRqLa205UXgrLMr0OmVJXLQWpg/v6liHerIwrkQOP/egGO+eER
ZfRulI3mZRKD75ba4kIhfmGANzCnMtLAVUy//yH9u5va+Vbq9MjYfKNt2KcHnnRg
Ms4DcN3bTtf1V84UJAqDIKtqrMsPWAmcS4cmDI8HFkMLfPuC/DH8mlGO96/4gT5a
kmqqqrEhTJu/2bfv0Nj5MospF6NMgkunG5avUQyDLPb/9Oi8KuVptlo2RdUmGGdf
+q1jUSLPKNCXPRUfBeZdJLb27x7ZUa50EFWsdpEXeuD9NxxFnwCOqZ3Q/1GrOXbK
Q/gj4IgvzmqASBxxGXeZr1QHp9O2v+rsibDCYkY1TKksSt/uE+AIJeKK7vUFGf3K
K/487Ggq8nEQIYGc6tUUK5mxEz6o3b60Zj/6LiziL6dX6pSAQ685ZgI2rivgr6km
5uLhLYGgZtXYr7u8e02OiWUWO+nW09eOBAVzOqES6bppXSSYQ3Dp3nvlnfGQed4Y
/bUXIsPlOMmqmEZdN/lfYhZ0HRF+09YsiHT2DZuvCEMP/90umvvoBsRwfr9zYVhl
o8W/BbPKMbKPHZvwijKIPwDjUrKrCpCWjEhw+LHR6PbA7MRQPNT4LE+dPp6HsWRh
0NNy5EVr2GM5z2FgcoVgcxRTfhSV74jo+CB1EoBZ1IAt1eJRawtWc/6M4U+fea2h
e1/ujCx5vnPVaTAz4Xvy1uOVzKLnGOLvKoVElXq3yUTE1J1MKYOG2v1oRyQZYB4b
iC0jchs4tu6X6H0ZRXc14iIFcAeCr3QsHmok7/ukOA12fQbTYTWlXkxCB039LwxK
F36q8Z7/AdXK4PdFTIBXpHzy9fXZjLNt9w2H5tdF8CaDgQVnDVSsGupGph7DK6Um
0LjOs84KX91LJPQ61oEQfYICAYYjhHY/UXqMwKhGTGEiXJJ6DqWctcqcxKMzp9oP
fBI2Jw9ZSxeekJZzRZTRkB+uGI9Bk3CcSvQTs0BGpkMulb0whEv+k7N6BYP95mZc
3US4i53JRv2234TnDkpY8iB/Eix4TsxPqvnqgEI8BCcIKcCgIfPnBEp2430zjuO3
9ZsbuPgOJvvrJ37Rpg/AQg5fCWKIytrgL+xYafAp9qTLWW33Qe7XonbT8Og86Lzy
DPI7GqYUApp6SSX6LZ+cK74EP3NKL+5V/arnmcApFt8akto+R8tLwkXFpeea1Rat
Lb2bP1hLtWx00BpqZsYMgiS3bMt3T08PC47moUrCxnRM0Ur/rrdJruu0axD0VCR+
0/w7zRYVs6m0DBOZZrF+sOtrxEIgG4WAER8pVgpHEuVgeCEoS7p38aUzJv49iMSm
WC1Rj7PE5MH+vyRKDvTBQ5p6FEpv6oFMLiBW8v95Ye03GfPypgLXrqoaUvmhJIJA
KyBm4w6XIjJsY00WOh4M6qW5fNTYYwipmaMi3hD4jiXY3Dq/obVQQylN8ouAMkHl
Yx/1iPtOMVjgG9lp78/i2+CL/6Y+rdJv79v4ZBxgUkA82q/5GC8Yl6UUwq6Nv/Id
P85i+wo5dvVP+/yJrzFFYzZn1IzNZnmP46sdS4w/sCm7HuuL/cGfeFLHrrn/ZS8w
dDGAR1d/cgqThJr3UcA0cXJ52C+2DG5AZ/b3L6mwL91/O+Hj2HlsXqVWrbmej3/4
rfnWR7TL/S0Z4dFZmyrvwvWNmRpTQIO/QcYT30Cq3zw2Qj/bF9YZc3GBbR1gwpza
54GIMbfJfg0Z+6LrYUnVqAPG87bYLFi9lmXKjnUR5my3wNJCkmhoMvKiCT2dYbj7
LT7yLfzqqFLY56jKlCIsJ2O13BCZx4IJcoJ28DujcjZ/INUPCbuHyPjbQUs8FSs7
dJEidOQLu1Ii4kdBUusM72ptdPeL8qb31KDsZxOBPb8vowsgUQKmGxQGOBl0G+sU
ihkWNtqx/LHypKVg9SXfa1ubaovK5Nx8Zb6v2TaRY5aUV6I6cjl2PhulO7TvQrp7
`pragma protect end_protected
