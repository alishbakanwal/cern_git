// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 14:01:31 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ib6J6nl/bBbR9iVYPJV9qcDc2/BkQGuA2DRab7LxoaTiF3iGqPCHMI4EPvn0sKrI
KXgQhxPdC6gIsIYxPIr30P7NcWtVcO45BjQM5bCh3G8bD2Nt00Rb34ufYgKxHrOa
eExIMTn51adED09jUI41ZXJ2pmei8XeSmGJfWBFf9E8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 13584)
Nh5GvWfPsM04xK1XEIBMcxsObjWRwMkvPDDRko/uEYSK5vMPl8cDiaXJD8DsedW1
6DuHhb8dgLbiNIrpIBrfKa0tw6f0V9yYNxic/zylN45dhoXAs1QJ9/tkySzNWO8P
HNrfnAJdCwkcxPTIjPGgTZdcbbjcIxW/pmCz+i3ZOSeDKStvWBssEfhSw112K+3Z
R6SSQF10HrZE0eXXrjEGdea/FpyaDhPICbM2hiFjkwrFhT8+Nol2k+bdgxkmLhSq
SEVYw4zWNTgUJkhzfalz3AvOqnKZWVfFM8dOTYuVjkE/Gazv9hn9nin4BhMx04jB
eMNoiSVcCQQ96HCSinj3iALm1BmzF/pWcixYJGyi+gv5r/+nTV2tnWwCpGj90ZyU
gZ2PU2i0VxeQMygpmeZheeUbwn+fBY7qji7injCDOXkbanonDmem5ZmUAyo/2Hig
iHfoUoYETRwDdd/OfyNq17g+aD/HcqijdndDuJOWLwyJbKqBONfgNutwa6ft+HWD
HgMWfOSYIPm6A79DrFYWmMLddaVTZiBVeIL7BgZ6szKcZM1KWzu5u4D7XPgxnXLE
OIfReA6FWwowKcoosGSIUqDBXTQum1JGZvirPwOEL6KtG55vyZznGes4lRqli700
wM1amQLn1uVwYW9/u+e8cWlihcoA68XQDCOh1DfYuGwCkfuPfZB4ELcw9NBx2U+C
/sztCAN3GtN0uxSdsCYtDnEeoAZxPtCWHfEkOUpoQEGDEnKyb/03a+c7Ixyz8Rht
yD72IaKwtMxMTRh5PSXLTzkjEdMWqAiaAdFUOe35pwi9TouV4r3/RCkcA0tDcRgA
8HW28TaZEfz5OX5yeXTMVak8ni3QkfRCzO4Uson8VgrfZv14BuyFP+tf4ey/053h
y30tepglQYQarvKomk7XCxt0TlJaK3HAFD0Faa8pO/SH0y7NnZz4pZLPCOjcmNDI
ldGra8WmUkoYyh7MNIP3Ms4pe5iWORXqHXTm1Pw/+EXiivT2QlJUuSXfyJc9f8ul
7wie/RHd6cCMqe3iS0J/0gXya2UEU9pRv4D74OL/b/q3eKpuIM1OlRkrEtc/3z9s
xIbiumnNqA2ff9cUC2CP1+TxUzfsb89kt9YWF+A6bOOheUjmvfqcU1yga7Bw/SQ/
JLeM3UzXLn2WwwuMz9AXbowy38oTlbHssH3A/fAwOwxE9VtEkp/6z3sEzG7NzxF+
ig9iyn0sNB/K0QEcyiC9i9QS9RasVKouAT+C646nRqGh9cCP4firi6eYPqtdIpCs
0ttCpuCqI1kLQTRDbsaU+Mlh+Y1fiRidx+mpRr6txn278PxdXp3TExW4oKbPuUqn
dudKIL2/A9dwlyxeDB7ExVmvbEIVtuKbD/lhnoWwtnGowkcY0OEUzX6WvcaG1NAp
j4mWV6vBzNhn9CzpI5924fA3uPg3nMyh/iFAW6uIV5fNCWejvfMhjktJ957ciNr+
J8zixQE/wdk1ug+3B+Ba1TuysvHXIgAp4Y6YdEHPo7vECVOZtQaayNaL/x4LvYUq
3WPbdWS0BAVSr6JqQBS/cqMs1FRCNP1N82BUOp2dy3Xjlf0Rr2GB0nwLwde6O6HY
MgtAkXFF9XxvmhFPKb0+/TssmxfOYiQJO2n9bT1+mWoIYLt3MYE3a8feO/5tdbub
EYCtBc9riQRNjRSOSYyMv5jGYffAjlhU0J1IfYi10BZK28uQ60N7lJmnLo4w/CLV
K2l+Mfu5CIFagwyI+oTZAJzfbvToI3AyOTfeTnBT20yo7tZN1w+DtxhvBi3IWPSL
OTUQxpE66eS39EXtGnYR6d8vElFXgnWLkKQYak3br18EirEvKxC9wedzwbF5B53I
Du+4QjBZkwwR8y/vsltk9K1ydWfjYJNiWeFgeF8P/ho4gdlPAEGzxYEbkUVMyiPi
1SOgj1BScKYNOotY74jI1U0ET4BFrzSC78rXhMnCypLpFVo/ABq3hfZRE6fQyn57
SqO/ocDRIwsJ3J/8pb/i2677cFSK1c5qZ/jZur7p6G/VuXC2vrCiskClAT0PWY4M
gLYBVdXFq/8p8Bt7DGKwxc893VGvDMYKNxb33CGXYmOL2w6row0U1hlSX3VCVvvf
oSliFcat6dEKFqa1fL4V55C9JXitE5ALb+B1Ss+Y53Wlu+XolVHFGPXW6tjB+nbV
FCFqMmoIX+NEZnSLSAr0bY+rTTxrJyGaPbmlRk86QUBWpjtWIL/bZd3XLfDStbB7
VDPdyDdY9KoMf3LGdkAsK9b62oQuJkB6aF4cpoMYcuQS/KOUFBH8GwXN/Oh09hlq
u8iiaFE5Ndi6aS+0yftPTyVgPmAPZ/0y5PADx1nD1eauNQvarEpnA3Ym/n2BjdSI
Cwe2oQJkDGrcgUv3cHIuL9BbORqtFkUAouwKXrQ4HRJa7hXOD397xlF209Y/60U6
mOHY4sTU6OFn27rAifmprQVNDOvmnF+G2qHoTWCHiatKzt/ncAi1+YTpcosHZu3o
YDK9QSpWig832uXmA6phlsdE/uoGEc4NShOfH3ABAQZ+awSq9yDW8v5sZv9d8RV2
/QKdrYakAlrWxo+tCv91TY4hTO5w7jxyWaeH4bdj9DlnLWbuvf/8Dfy2OaC7iArq
FhDIIZkePv2/qR6ehsR3hVe/K5i9TLZyOIx9nbDQjNgLf5LaNT1k7ZblIcl94yGY
3ljyI8dBYKtraOuW4W2E8Li/0IdR29K1C0tcKpegtn+mSGPONHHSH960bzwZWzeB
iBLxkLZwyAzxEmaKrnuwFIim5e4eZh3sp3N44udI61w/6am48WYxmtljdHNSJC4N
C7s+JhbTM/wDxb/OgosKF9QIjEEyacIeBA2H/3EAMEFo09vM5Vg2DgM0m8VSLHxY
TCfBXzLx8gIibB5jHSsgif8NxjAPdyd5eVKsPZUImqXW4rJdsQHqg34MENQvsd9B
ldQavcL2Hl5vHJZtC2se6yDNaNe+6X7gMEFRKOgZflywNKenP71HJSEX61zZA/Aj
ExDBH62MUKLjP9djqcyfkQpZVmU9trglvPDD3wtrFvm2VNkTxPEt0ucXzpH4GWOl
sjPb4U1GZLG/QX4VlXaz96T10vrp3RCm+OC2jYofg7yVPG7Y3jOV9ZBMVbXaLmiU
1on1c3U1jWEoKXxIJYl+7Rm5Sj6wZnXd5vvqswtOC7l7ZAC390SQPT5sVldME36Q
3+XkIsBxbee65uGFtZ1gFH0eITq5RpJq75iUt0csuw8l6soGmqSYNP48ER3j4mDy
AHu68sz1EDZt+yjsl+q7OtTQH5cK8egSWWkoiSHn7vcRf3mpXaPZvvEcYyooJzYa
Esh5JBAABRnRX/DNupfnxgSiM1AlufcH6AGzI8K8ggrfrSmKb9g3M++lWEzR3PTN
KN+zd68ZRnycPOihqr0lCDziL2pYsNZ2SiYQmzPEvAVfmhmy7f5DmJFub9qwxv9V
MZOJgLxcMWr9e9e62QEh/YHBOdiNJBDXA5DFM4r8aWmfRhhG6Kcb4kAAK6EnIilH
SEqgxwGLBZk4zuXLaRUgqbk7jTroMfqLHZj3L60koU/CKK18154I9b+rE/DaCTEp
8DdY8CO56KGu56uv2+vadJSQ4irfmSgUhW17Hn0Nh+ZvkruNfJaCNceHTG2RZ/nw
QEZ+MDGGySZfzYsfIScd5P40K3M/fp8+lmWjs3P83z2vfupUWfSId1WchB/b3806
k3wqhQBGV+j/1ixdMqlcZ2ZXC5Zr55B2K7i7uZyaknE+XPawyB+PEja9RaUewX7z
e9wl2PsftCCFoaEgbXxZlM/FUAa5QYnTYLgkJwHbumEkwEidZwLnyUnxBwHz3IWx
po47MZ3LuDOe6O2cl597SKYuMKa0DloXYd2idd6/gDyREPAvUaRZZs2gFSpkwpM7
azl7XZK58v36hhyDzvt25JbZiVdlDxmGAYn4apD8FJVk9tgpqu2VRIWQmrs7HirP
ZZK7NRAZBiy5ana4AzGucKafMo/Y3enBhzn39Dre2J1AbX+Gf3njRg/XroK/2vTK
o1l8Cjr42tpHGYpd8kBiO8RGBhjWgbPB4A0BnByXrY800cwL9lZiKiMtokO4cOhG
eFMiTvPZx1bRNdXtyVW/ilC8H7+jbmqbDwQKZWJzMWkHVhqKsFobndNHRRpPRVSv
nkzInhJbKlzfDieVkTP1hL2KWPWbn4BArrZsAeKXDz8td5Vw6mx++fsZTh98pZjs
oEZVTNEZeSy+B4HsFjTk2/yaOANOk1dhbVNUky/UUZLKXNRZmx4SdPbZGm8NPdJV
TgDZPzVrcD9MtZKxhzPm5SsXXqoq1TkCtasWXyaChd+GlOoVS6kln1UN6ghnHnYM
T+DHgZ0IPy5QpFVh0wLn0tqeScnDGFLAhMepZUXdh59KRtA/SMVOJNKUO520pXn+
/b1VCJl9Fzns86os5DH9imihUHHUImT/UGdyCaENVwHunYRoSlOy+wQITPL46BGY
+vYFPJ8RIcbCuSnp2FKlMHZiq0wDQ/Jlv86B+5KIsAiJzR1IIT94o3xhSWuJtjaZ
cxuuZOgXx2v3zBfyVpWavbhfpiWAdIHlF72vhhmOKW8fLGKV2hwdS8/blxZ0Ybph
WKxT+RG80OIlsXePvbInh+FrSl5x5IfLBNOGX4YZHaxJcoGE1BTbt6uHTXBMumqF
+ru+9X9J8/UzOQQOPk28/lOE/FSw9jtrZp1nIojqeTITOABk09WRL1F21foFyt6l
NZCyVk6Dca/uWROqR0Kuv71dsdhoe0r2STlLHEdpXZKQyF2Wdpsu2VJmYkh6H2WL
NGa6SbEwT0+gbN6hPyIKdPRggvXJn3uitPXSEJ1y4LYUXF8acz9pFxiaemQUsVVW
O2Dn8+Bce1yL3JNMmf+MkqdPpJy7G2mz6DJtranNUp6i/aj32BKR+HDKseNVMiEv
A29/vPQAtMu2eq8hrpqdMmZDEFzfFKWh3pol+AFW5BcT/50LQA+aumHW67o16bN7
93YSUm5Suv+PjnPVsyg7yq3B28JgM7hLhqz7d47Optqc8GhnYknGdz7aLvXoDpp/
6pGmi8dbJQphik65pNpzvkvQP7kUBPnpsC0h5yvrfWOCtB3Bk0Nx7AjyMjtwaUkK
awNzrA4kXK6dcse2uxIvuTtW3hoKPCiDM6LrwSXulFQ0gdF5v/iXwvSwYqx5af27
m7XSnJ+Ba3jHHtHrjDobSx3sXlYGPUpzgYCm8w/+qLeDzUJvGkiabNNVhyV4RlsQ
Dk+3P3psDqDL5IiYCi9++RJYBJm11gNktamBkLL9GtbW19BCBaEJ4aWeVre8IhHH
u3QwVbQ/mQ+k99WQpjNTMjgFeYWynkMYcCD+ylBzihgL493GwohBLQQtLviQoPou
W2JLKmpeBvXvPNj9txDdUp8dbPzBGnsA/g+uGnJmub4TRDcjJndEFzBEQ3dkFTXy
8PSX5yIcE2INr0LQeHkNbMP1AsL9Mn8XyBPRaVqoiYFdk41tJSTLKwlrBpazzg/6
KOPqzu921VxXmz7tRuHQRLOecizg2l38MLmdJVS6zxWQRLOjIjkZtZmip09t492y
de7ZPvFvPsYbfeZaCKefZjvqOxaLdZGcP6aqrtdhbGT4fZTgd0SvmKlj9OwRpM4M
Njn19lX/hH4LN5PIJ5BAA5NF7uuTLgvWYowLLTm/wqpnC3maOrj95a64U6w8motv
K1W4UoRLZ+/bmCVSLSzRfMz3zwEjMODRL/L1gcVG5XnOIGS9O0CTE7DmWEM8wnSL
4QhdmfVYVGLlwBvYm623BU/HuSxKa/6KDFN1G8GptIq2QfCVYN2ogctrn4RBFC3T
geV/9jpvxSfqvdb0mYL2dLdcj1p9d7VhBS36Z1ydDZBaoILgRFRo0gdQn5WN5Su2
b0VcPJel2oH7gygzTjiaM+kB4d0v4zAXsSOwXzHh7gdNxnGHubidlDsk9rJEaShp
SytWlDohCSRIChi/914k8gYbBi4e8kUunNyWcGXb4ASj4F6zUodNtDkRDHs2t35S
QFtrZ7oZVObRW6Ac3sFn1NmTmFb6ZmuvLsfIzkqzXrYTlWaRUTs5aTWy49ugnOs/
PBsM/kXOIO94MWYQzJIVId5Je/hxeYtOMm6AGgN3lChk3cDkbhDan0r1ZSWgc8Fy
lTT0eerxnxLIhczNntYNXTqNApC21VpOR1a5EfT65k6WmI9AyN+zGsrp5a5dBFPU
niCU5vId1j2uqXDiIBU7EN5wfjEF1gD5CViHxkHRnUw3IdSXA81L5F1XT0HBEZbD
YfyFhpNfIxFS44rnz3nufak9c/jIKgOkRO7pJ1/1kT+4nbbsD4HIzhrAqmxEO9/f
8Y2oSZgSpg8o3qVhOIHzCdDJLJYxdzFMTKoKGyW4+bTdGpQYcpaFo7U/SEy6FF6p
YvKJuDH/Pv5wxxBlmZ//vBhCpkxtQODvd1xdAzvR1FDhwDEA1846j9Drn6ombbPf
/4Dgyz9uhEuxNefgWql9dkb1tf8a4+VybLpbBfo88gJ18sMfdZZVp/dLxMei1ayX
yNCa982I0SlPTjQCbz+6n4xN4OYLykZHGJCrJGkoNy8GyUD9O5tmqnIgxjn45JTW
LDExqRW5o0wqySWTz0+PsZ2+NobSELsIo4/UydbxRnCmAbVxMTJDo/eB4IiiSO30
+auJdbpbpaNQzjuq9EP1FdkmK7Dx7q5YiDRHgHy97ffCbAOBLJqPe4QXL1XBv0GH
Tt67L2x2rpRTsQYb6FFchW4lN//KSsYJ7uTZjlVCwZJCyYb/8aLyUZ9t3UaNeVpX
wI51OgUSMv3QXskbORJY185PoBRFK9j6bksI8I7Gp+oDfItcIGXRp7rYiTKFyoHr
ZsqJDo2Gu9QvvDkYT2qr5gb6VI2QVlqb7O8E4Mm+nA7EWnTXna+xBYEPK0AE/5El
FxTpOT0cGf8AN5tuKh1hnIVLqJHASy6hghWE7j+Hoh3PvNiFotxkGAnMGRGX5e9J
vjCbxHHK9IO9o9+ITIbwsj1lu3CmGwuOVL+DxNUVZf2X39AZCEw90kS5wL+PICjh
zyv3k+q492L7MwbTxHPRaa8HZhywrFlYhtFy0IlOqzpeUcgeGQ8OWFhPqTMhYEru
VBbAWdvPqSyK4mncdT3yR9nF5P1OHHNxnFoB53uAcnGNtO1N7kP9RCgUO5Rk61lI
1R+ODrMaSsqdn1p6wx2HB7godq8SiuHDzoBm6KCWPByloAxBPIP1TLpu7oCZfPeG
POvzfRqBNZjE/KsqzWoS1lEACdMnXKIZ8DCrEMLRc3rG/OPCBdgWayCun2GjFNha
cUiTMrL6S55qr+hY5RA5Jj170mFdRk7ry6wjtjEddemDeg1BaiUaOZTwnnR3Q6tR
U7w6edmlk9Zv8ye0qkHoAShauEhYeqvXxUE5sYeRMcGo7yRObZGPqdpLok5fx5WK
GRV6E09iiQ1MfU/9xXq1OhfpoJ7te/JSTVUJHCLvb8AB+jdf6b9/mJGjwaT5rhU9
1LssXB74FcGnysdtxiFHSgLr25YuEZCfiuUizhrso6J7TsRUfZ7kCmzpQxiRb7XA
btp0P/hJNybnSH59aUa8yat1PDOuT5iHckN+4OWQ5S6+ib4PeC90RLyThw9Y8dVV
bKw9tFzBlrCNhZwv8hkCcaDH3sKBjptbWiu6tQ7ng4E0Zp/fN0H9RRDEUEzKHD+I
pmGer5iuNgZL+MLNgGYPw6YSvQxaZMUnbpUCynm8FSHjyMrSk0Dh94Ly/9V+H/Uv
2CcyO/xTrEx3cXvt4Cf6hI7w5a+hoFtpgDl+wP8Ox/Un822A5iPcw6HyqcrubeaV
I98tqQv3TLfJQTw07+1Hsjyg0i28PHMOZXUB5oscgMdm+szB5Iq3s8hI5jH2I3LW
xbM5uud3TLR3ypQC7RLF5hQ5loXGGsomhG0XUFV+e9QVu9qNxGlONmj8tj7ddpyQ
LIAGL/xSQk72o4Fw5Txp53HnjeU9/OXY/PA2FzUsHpv1o46jafWp4asVGEVN+NoB
p3yquaSI/E1FKbuBMFJq9Bq30pZPgvfLish833Qd1hVFoSdYRKyDCqmI/2UQkZPu
68hZjc/B7AxfLFP/22mwHUZRs1b4MkmpKSFHmhX9+ltXL4YQb7Yf+garda20+Gvn
d1s7+VyZgV55a44XlrkR28J35dhPfOUB6HxWRwPwZuQ1Hs8mGKfhu5Irom68AiDe
uPZyZF8PbU1+aYErWmt5QE3msxKpvomt90dxrfpSOrLy5CtV9xAVPsohtjjafqy6
4QhQ/DLQ6fy8E6sCLBR5OvPSQD6/Vbxc/bpoR2sBpXJMoyeIVZQBdBry6mlI7QhV
dlzbroQGv+m/kU1MjZAsslyvz2DVSMy/y1E1CKAz263SJ/RPIqZ4fOHOT5s4TsUf
De0xuyYawfGtcjV/f7HUoXkPO1QVhSM0qvCijYSStWOQnW+2LVDXFbRLHdaQnKHY
Y7d9lOwq6YkhGgOSAA8dZrtmijk8ZVI+rb1X0sN4jr5mXVvE4YVIvxv/lWYcKV6g
M71MlKeEpqzP4FGdy0DuMK8WsYhn5rUCza/s7Yq89TI8bHyNC4wESfxt+ceLUOgN
HGM12013GMfpwRjvOgGCwmeVw3FEHaTvWAs7fPQt0O71zLxWyaHtW4YoAWAsPD89
6zeQf/LjUvmc3paIN+7f/5xp6GYJCjpJMKfdjf4Ldt7lDoZIqbRZ5qJyys83x1nG
ACZP8WnV83UfWS0YtPmHYDGwirKEaMxsBsqoOMCWZT9hM+3OcyWbEUbpWZj2clov
We8AwkRkEVGrYDyBb2LaQs2sUSd98saerbPLkmI57gYiF3EwjO/KOiXNd5Kvpj98
5ToSfrxaalKgWUmKw75zZ6RAgpcoyWKkYZopLzhdCV4NM2ULQ/S5KGXA6MnN3iWm
4SrW/Eg1mG+d71hSrlnPRfmZS2u0S2zgoxKrgFmM4CJX4DkyzJ7MCoTe0e2FF9r2
6eDRHZ62V9g2TrAi7/gtSTI9Pol5fp8In24CmjvNhs0o+vNuvKP4tKbZ/vU+rgLM
eu7v3JCXUWKM5oFyJLvBI4YMr1Mvia7nZdFoN4a2lUHlPgBJKlluY0WNXncxi/Xp
M1Z6uVXkvrHe/BuKQWCD1Xp75svvdROWKEDbflmpPQIZ9aQyGI6igneJsJmSzbSv
9//rzv2Q8xYv0L7nT+MC/3Fnipu5fqboRLJt8dfHXNhnN7W2rTxj5cbi6S09MdiE
QY9tsuzfOImfxjHI/N2td0mtVzJak6qyEXNsgVlt3LCVGQkZejAT4fTvcZqDhhub
pCq/04zIVn/nsaqtv+V8c0ariyDvgjuCl6Ix72odeQ11Ug32zhQdZlV91podkffd
tU5Lzqz4orU2FE/lQx5z7m61AnmBtfpTiFD8Ve7fQABzU6+sq1xpfxX+6uRoxskH
V2ID3jCQ8tYKlzr2Y6OgMWN4ALgXcx6BHlDC39e4zcuTryN/9LPWaKIhiGqYz2AC
hvrwGCZk0Wj6xIQE/AkcO26E3N9iFXBMmagef3eMGMx8Vdq3RgP6GjQzYTrjUsxR
a4jLxbxDSJ6vUXCeXszh/ZJ7HsEzY45gQW7H7e6JkYIJBIUhbmd+bwXUInru96wA
xkkDzPDqP07hmdzyjBHd5nBVoeZi4Y3TrmC/brp2tAOoPQLlRrmjSFWSEGVZOrt+
dWQUYDz7zq6R8B2nOIK0MYKY5PBlIKbsYPQllgQmOabD7JO38VJzX3PswujVpfsh
wmkniZP1g3PdqWiDJoHwaVG0jeRLl5+YdZnEAK5nWj2L4ouJXHawoN+8yfX3stkh
cmYQm5WjLiab8VzCg8638calgK2uK6HHF+BbEPG9g+PsdvrZhw8mxWnD9LkufTBT
vFbfoNu4wDUQwov7psjWv7lSsPCgIUS+VERSPdHJ+1SfpZhuu7V7AUbMo4PFziQD
m2OjCUfUkIqRTj2m0g6zPjQww9vfytCGxhEiIPDpjMNMITB5peGoB5E5pTW94Z0S
HsNnJsCX+kau730TxnyGn6WCLJrW0hHWfOu9wWtXe0SmVjdpyfVVWvwzzZE8Oiw4
Zd5JW7ywcRRXX34B46OfEiPUtR7IOyZuDJgR5T06vo/QnfwhO9zC3vSMSl+jN2zx
joCxEEEL6DZorgajqkotBVnXKrcuYTLRVEWBu8l/Qu+AYUcpCHKzss5eVlZY4IDb
B5DVeim8QOItNxxiMJXwXnWs0xwtKLl4SSD2LayAxcqkX9jj5UPDhNrve9ybETSK
6zkOntrj3m8Oz08mfJtDBvsYw0GOPcglYhA9v9UOhWwUM5DkplVKBhGnw7gbGEUT
d/VLmbPAtN7nLVfAeZfbGev6fWwnlAwGgpu6IPTnqeIjNxDdBR2HsbeV1ReUbWz1
dmbHxeGVvcGIRPlCEq5WfXkqTnjGpwWUjiE7CQgZ+sN7IX6Y9lTJxFytIn9zrJgm
J0wHTc/Knb2QX1DL/aTPC/AtyaRiNq8zfb+XLqAn/wTvV7+UY8fCelTpqEELGp7v
5yempjokzxLsTKaH9DjZXAq/wweuNNcG+PlyMelpBqgXR4IzzrDfD5Jcuc2/hsyl
wnEBrzeplA4pZ9zptRvTQRfTLofZAlBcjve0I/P4SsMnFBGFTgmalhS+E0ukceJt
2UDeMAYYO/nwesHth0+E29jrjGB6QlggRf+SABArkbl4vPSxSrBvZQ1t7Kc/oT9W
BvUgZAUeuReaPeHhJSGu/1NCYlmFjilu2qg0DfSafafHZ9Y1GKicCH16Bk9OIx44
ba9Gcj5xU6vJZQaSf6CQT4iMaDF8J8F9gwcCgkFjNru0EmiFuOhv8tp2XviQLrsd
/c0oaGoYj3BOZNJ3qqStXbP59RPJhu0+/IdFcrKDhkNMfwQADDORB9R7fF7pWhHg
8SJppFt4evKMen33nApcF9np0yJhXHvXiXxqhGmi5iPG4/SthlEGKo86WwAxaWtD
dlbeihjn4l2ljeiZ9K5W0c7NlO726xZqyvCHzdz8jJtqjRTYejPXuK4/9Cl5H06A
pbBhRyzB//NdOsJM+jFIVshdNTV9m8JCm++eKL+gND5Q06peQPKhtNH8A8P/GihI
uTf8ecbSEp9owqA+a6HukT3egDuATrC+FIogavXw8HYaFE5To8ZC7XBp8/HhsCFq
rwd0BKNFOdjwXOsH2eJ45bLkODLox9YupwehZa8WSQwl/pEfO7TnO/yT2VI1chOA
bRbeg8wAtOuLU7quG+48mLg5Vf+yb1dkMAdM9XVZs0aflOIW7tl8OImyGIsiAyrd
nmRLWrOJyqpXlwztbYK4xLurISpX+bSnqKVgtn0AL5Gg+0L3rK901kGQUHqmCX3T
ty74+UhEYcvb3eLJUuknKScDCX0L3/NXm0lE3MwOpBoPu3cgCWMAPFyk6e3ipDOH
Pp92/dPHOvCUYjZ76xWvrBZ2IMVFpQdgSpWcWegHn9xgG62WAn0TmwdBN1mEFOh4
9wrrIgzGGDhhMyDJfIB91iMTKh6jxzmEVvZfk2CnQkMTcUI1AQ2CwriMw81RgJKy
QUfrl14YO00+d6a3v/bodkBqcWMJ9tK7tKXKcMCZ9FIMUma1MXniFv9FwRwYBFdv
Gm3QqX8yffepMcIIoRCbFwGszRenWuZ0L+3J7LX5HwpYctlnkM+V7ahL+Za72SoX
x8vSxDB73oKYE34CnRvWNfLA3ag9S9HsccMf2qK/4+pMuwDOfO+8RPkAyCDtS9AU
UvnSJa8NVaBa329T4BgID08q0IY00CZywV/R+05/ceW25h/0YeB6qeLS1rqUBuAj
KE+1Mz2/d1vPb/6HTAM0KCxsG1YHbJkQgMIuvFd7sOFLbaBQIMnS1Qe6t/7wkf4u
4ME0t+NQFEuppp7MbsSGcwyF0ux6vpEHJdNgV0YyeRhPvWM7RGVleI7DaPTEvsSL
cCEUcPspW23GAdanC0JNazx+rtHUlreB+bNhExHHnwDYqhVqxN6ausVg9tLWqr4B
f48BCzfnr0FVEG1JyYWf767aLWarZ65i4xfWKrfMG0Wtz/jLTRWKWD/ToK0BcTTT
5/C8Uob62kGveoJAt57qdML+rWDpm8930FIhM0O8g8dQtkoEkkycPj7li1zDf9vs
pYbNPJTqmr+RnUc/D0Lpw/AeMGz7gM03lJ20K/l+65RtYLK7QOcl7ogVPiyGJegb
NNHPIkfS/N+cYgP/uxH7Uayng9I1xKmuUDcYQAxo8E4WJ9lpU6GfV3jLR6656gGA
pOJeonjqq4ErHvQxu3EzGrue8RRHmFeNnzj60idJGLEsY37VUT95rj4BzhDjrL0E
0m/8Wdq01UGp4E+/rvFGuRvMxQJ9B0EwN8/7gb2EhU7NMIFmwJyfOKHBOWnAU7xl
yKWDM9QR0mugMePZ10J6Wk8L5b7pz6T3TSj/VwezXubOduZMIBrT02Hp4ewQW8tV
nLBofHGY06Ff9fTqUHdq692lVDU9jyD6TSASNWKrhKXKFGZChYoW1uGjQPa/oXJh
Z4P2ye3dWEKelndk+4j3CLtpUZNQVzI8+4Zi0crbviLhL78zk6pex03IyvzUSA3t
y8o0SR5i3ZwgbV7S60empqRIutz9/ukwTMdLwMgOQllVeYRkyzbQoiXBhq32BWpm
a9G9HBXNZVvKHW0TXyZvnb3lRnw5ZMph7FY6xBI5JIiDcHWtmWqNt1T0qvueSPyu
NtlOmdCdO0Di4NOzntwcZcn76o3WHT5LF7LNuZTkBaKI+s6tZOg8r0dMoOmHaxS/
yrgin1kbyQin5eAousFGofE0W98bkNr2h6Sw8pYvdoLC7bPGwCM8ESWz5JkA4BGx
sqNTEYlcsJ4FF/ZVwCiwsM74DE9NNQ/N2u+Pr8EAMGDdvlhVsXAVCfZ/FejmrjUs
r1c7r5FkCbv2/qdaNxjud9tHMeo9JE7p69bsgNLp4TXGFMKQGuPPwNBTTRtPGXPT
e+ukcojnwbLEETOEFCnGDO7K7GZlsxQNWibvpWldLc07QHc1e7MFNrZrYGSITjii
tfoYG6bf1BB2U+xXwDM8/x3NXhP7VemZuQZH+UJBmqM9hXdfbDiCsX/doCh1bEMz
8fT1sUN0bGTrWbWoYoqKmw7xn0mWVa12ofzgDcq/WKmn1NmapZzRFCJMgw3i3ZBz
j4YJnOVZcf5f6MBHDwVkmBHm1ZfC/WYUCTQY6A8ij+o7FFq90cgD5kDpQK72aXWA
j9u9+Htjhv3DuwhzEZnCr4F5GnjHTfFDG0GJi5wCwUEkUC6ny24oVW0ZLIN2rKAX
ZGX7lUf4R7tGRfR6CpISw8/NHHijjxnNcAtIih7tAnLkwryYekCTSaczsjsHmoYT
SoOd0a+7s6L6tnSm8VdovCRC7mfOYwvc9o1Z8dRaaRmh1ghQb0wtpvyHCL077T5+
DaR6BchBKPn4zuD3XQwZ/OVmuJR1x59twGzRls/Z46yoRXVtSqAmqiPAOJZchVVL
fsTjBqAY8VsYXcr6fGMMi7c7EIs6mAns7qxxhQNvT5PaIqCFmBCSm8vZfno9IuGC
DBkvLp45xaY8vh0cCBHlPN5y/NW1FD/npGQ5oOJnFnRlq5jp3aBnRp1zqZTR3alA
pPwBncs3xQboIXP4Wp58pO09C5IwtY4Q6hohGCaiYf99KNbhVUo8qcqRra5Vr9+G
KUpemwKCrL3DDjamNYh5p5CgI5NmjEfZMuEGnqn/Eho+FKa/YwS7u/lkex1h0mJE
BJVNv8g8wvmO7Fn0cSFtjeir5PwUgPlpZyRtV+CpbIMO3vBJDjqXWBRc2vOD9tKD
lOb26bQV5FL7G4+v29nfbVc87c2Pl2ScSfYSEnWQ86nuW/BhZqmZ32/yZWKnixPE
ohh2hXic6gob3J478VaGKPoma6gTmE68wJ7/eLItlFaE2aLQJ8o3c6yStt0BVtd4
C2grIUXagrhwBcbnHuvIn6Sc0rAKd8fbmNzVoyODMx31NYh5F005SXr+5utqzT9S
xjByRwM2fCnufmftzX8mpv6oBKAVGuAhvwekl5UlHUIx89keUGTGwNG2nq4V9EEc
S/jW/IO0WhlTLjmRQv22ZmDiOzZsJkUeH1NBLKB1D01GVMpK2Kt55IjZPka+bMNh
QfF4AYHgb8XikowqXOw28eNFi5i8x5xJFHI0fLlO47cHkMHrTT+eCRgJy75x23Bh
NbSUrE1KNuOgpc6iPZAD1aHwH7xeZsmNWvd8+9Ng37x5qBAQiveAnZ4dlrUTUD9N
/3Kk7arxASenBQf+Ry30N+F8vO/QuIFp2F0yzj4sTs4cRT2W1mC1V8Aw+iw1X3Ve
VIb2N/+MUaQ0PWY13q9e5qebzeSZ6xLtGZ9OyAukGhjpwrqv3R15aW7tuwGjaM6M
odO2F32+wY2FDjCv4XMSdtQZxycxih4b9CK0jF9PuiK2EPfjZtypIKH5X9oLSNhT
ZxcuAILmo8kqEDFtZHEhdT/3jDYysLdoy98177US1tPv1Bk2cTuihjibx0LHelK9
orguIGOBlQAxqMoO4HDb1jOrctuz5yt1vkSgcZ5/MhvQpyTJIXQ7OzvLiT7rsExU
wcUB+QwPw+tEb7TAkxFkmEznJ+4jfEt3onrVMMhc26zoEEdwtLg3Qtl9KdxkRuD8
ZbcBbw4fRmbTeOwT5WX84kRusNllFI2wbJp0sR7C71yRr6VF/KFRU4oMMUvrEgnU
NulDUw+Rjv1oJACTLLldAyvOf3TrML/5vKopG0lt2stePmL9Z55rpTUiKLkadTdj
yeCWixBWATxdGoxd9ZoQqGjpCY5YC0HvPW+LLky/wtwyYe2YiMsfCrSzRakN2fi5
yPaz7qE6hkbHvd0HL55Z+K82J/wl8vBUkRKxX57qc6cYWI8nOGV6Xw2EsOLRGxkh
tcCK1AfOeCi+NuN4UhCKHKH2R/xzDl7a+z1gLaET6FKQNFWXK1TLddEj+CIZg0On
GN5BvfHxrcLYiNtGHRAcABZajIuYgb2DR0I8T0hhqluE4d8QoB15/nYi9o1ZMFdF
DyZgGb8Zh+JKx9iQPkoqEM4ouQRWlEa9BA3oymclYkJge6TTez3c6zMhnNDoJ53I
aJsIM49A7sU9CbxZgqzVcYtwRGbLY+9jLal98mP9AEc1ST3kHekluC4YLPpMaMFR
PrCyTB4kwaY7+I8ghpBqzKLOJd3rQN+4TWorLYweNqJ8S6IiiEt7fHR4ydcw5d84
07ZaBnieybGYIbWZu2qPhs4xSsY039+UclFdWqk71CTcRckRI6K8OKwJm9A63AuP
EA74tmITc1GIJLMSjGqk7hrGceCP7ZV1/rOY/WCUgsEh2leEB2/oSvxU8R3xWUpv
aeMOxtWaUnC/665L69Ewmn7s5CzbUdUBOJANSX+pzaoMdVzcqkNBwDO9ZXHvZsKI
gBpNlTQjzSQYhCG/3fW3kFcRM+6MueCMWoVGxwmagqv0FXEr4xfiyzaihuaMIH5E
UBdhgSj+U+tqvmP9KNWJ0Kowi8yMgoHYSdBgjbrbrub77h/GO99MhU6Wznh+TqXS
trC5SXWzdnJGTphKVh55oFrq6CjwtGZ6weReA1LvOs4Oz3E0O0fcJgYyuNLX9oKC
jqJSTykts+IE4WEE2WUhLcFTGgACApqk2Cb6plFZh6ALwWZM1E1DVcYA1RIWAMNY
GQisi0/deflhFWCdZVNr9xYPbgGx54JZ9zMCox16x3aczV/wlt81bFoPVYRAz8wf
njVwWVNGH5Nr1WNtUW2CxrjkDqkJcSWbUhV7DpN+8VFHexZICjid5vOUID8AnLgh
+fbZEQirBHQH8aolIwP/drUyBh/eZwLO5vXinfg7kGRxZESU5Dl96GceK+fQjRXW
ZonZJTm/h5IpfqudxXb15WbzYbSI3/kmpSmsN0rReR47sDzH/q3D8Z6wsbbL2dvH
OKKc1M7R9+YSgUDagCiM+bTqbHKrKAn5b+frT7vnQMCAl3RoVQRgR7SIO7NJx5nL
V7aDmXrUTpl1t7tGLH7Lbtf2v+7euI5Firhv9toAN5SgdCgcoTZ8JLcT8q+sTy6k
ImSjZgj09Ysvqxc5VMBiUXxxIAmXaOg5bOIMnTQFnlJihoVl7bh/Yx27e2mf683D
SgZLDzFORBdnOiY/Iaif/gtfQyjF3hhMGUpEgPzLrzLIRnhkotMjoXKP1ejT3xa8
9sPer9Ri8ZpaDvgqH59eYYMisbSbwDbo80aWJ+Ja+yiYCIaFIRON14wNzkN+GPaN
/mIUUTwBIyiSSZY+SKm/6ebfly66HlbMPzydLw1wzfpSAtoVqJ84ll7/zRQ+o56H
FM761zI4NunGYL8K/i0koOT1IwrHdXH6cqZbfUydJk58xgIuu8lOTbmFra2op4YV
hRehWo8AdVB5Bulc2FyJ50cYy7SF/V5359RM3ka8cykVMX9XTrrWICXcd9c7MZuk
/2dtxsPQ+ws+X+cXHa2XXslmDuqIqjC7ZapKHMR41WkrQ7xc69XA0j7cus+m37ke
fEUP/rCr5ma0ZsYce9YQWqR8+ihlV9n9ktRGLhiBr03AfYvqG09wiN1k8tu5E/fc
KLF8HzxdVkQ3PF7vu5fcJF6MYtbcXtS+0K+TK1dEYcaQJFUiZlCaHo6PLwjFp28D
XebiTaQiSaAckgPKhoXJzR8aZy0T0p1jQMnIlGHjm5C+D2LbKJp6LNhlFHTk8aN8
UbX+81nMluIDpVNeezUv+jMhr7SXk3a8vqbvR/8nVIgDnxThg1JZZWxedP2YTQbO
ezmFyJ5JL1FmIBA5mBu8uCXRLMvc3kJUKrNW7xaFwVWgMQQmBJW+1rDCIOyHY8fM
Vrnm4qF2aL/uJOYI4z95cXAZtT0LmnewFyd8jnR1iIxPW1/8EthES6J8ODulMu5F
ZKvZe+Dm6+6m0tGo5UBMx9fzK0reBs4Nm+0vhPGER0oGj4jk91uvXmHcfnTLYL7i
Opfl+49s76BKJVq6X5OjQ8KPHq9tWxFgKTJ0MTdjVwFB9MFesHeCxY6+CKk1wdB9
jRkRAG697GQ4hm/VYMyQ3x3R7z7RquoRRoN4yxScd73neyRKKXNwtapepGKwSHWH
nsA/limmvd4rNm+i7+j8sgv43/XUJuu84VWk3kyzZ3I1FcwNn8n8snoVz4zc0mVC
jyZ1RWRctuvhInJHVgAG67rGhG1KNe0ZB1fSY6wIUkHHTNJT1f9d6Qxe6tNCM39W
8QiZAfJimth/yxoO+z1VQc9vmFP6nlLzTaqT8xGJdI/ZM6ZeJmaLEHW21kpWzvL+
OxPcgcQ2HtJQw3hrCtZYe0gu0qBlr99YRGvh2A0Csd7edFDqAaDb3j49xd1+R9cl
SwKkX2Ts0ZWEV023+XCOB07UFfDqdTc/u5DTmMQydEVtinTLDzZuHp6/t8U9fQYo
QLyroCfzEjQWbraTM5XdLAzYZhjXyuXCg7tqPwBTQEiqKngxQBtmf3D0mxUNzBFa
jFBNwslwG/5nHKPlURp4EBTPiFbtpGhgRqt0M3I+JK6Glu+SxmdSZMHquHH1jSuU
AK1c1r4tt8Ij3F7WSWbLCdmy9eP+6Awv1TyIZJjOP2Ry8cEx2Y2oCOoUeGQl8YC9
FX4fdMA+1jbp9fhZb9kn55ZeIKwOUGzeoa5n9DkiK4Z0dAQkUMcJm2n8APWDL2qD
sfX75qO30CvAkJB3T4bl/vlhBuAMzZiPQUW4v/naoTYXA5zI9j7x12eFRCqtF3YM
4KnCZGguL2Rbh3rDkAY+zuPPWTpd4UpLNLdUlY3fe3/a4+Lx6fyMTaw9o52OUsdc
4Map0yP9aiF78KjxGRWiNVJsVo8M+7EauaoUK/hgJVvZUd+WVYftLl4/bqRepDqW
mzAYUmP301RmPip90IC8Asy2L0IxTMiJvULO6GhlX/MK3VDVC7c00rIlOXEH9CDI
IS4qysFOYd1NreyHmZ1czF6gkINlqul/eIBXZkGYYRMtskZOzDDdQrJ+nVEEVI92
y9I5L62NYXSNkdpKm9u44PIy9VUeAqT+LZXgWRLhRk5RiDC1cQo03um0TxWEHP63
BfxCjQuhwDaJJ1x3s20zHDfxgYIFIs03wyqkevPeH9H418pa+NVS73prcDeyDMze
RKZvfpMthPZ9NJnHnJMXQAPr8OdxYsOTFX/YhqSbSM2HYURIDnE3WzbwHeEqWFJM
`pragma protect end_protected
