// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:05:36 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
W9/kfLzvVP0NFdIoifr+LM2AkhygddX67LZBapFoeU93NI97mzVxhn6G7qvlLR5f
iWfPgOVMMuuDid7RWOZKV/rUysnvYe6fxeRjFJZja/4a30z3kBvGEuScTxf6KpRh
SYUu+q0ogc40nMLg81rydAa48waDilpo8ZelLgg7RHM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 22624)
8eJfLTCrYTk+vlOZo4SAhHoiJ2y4W8pVsrX9+i5vIY2he4fYtXesvrcBVjQ1beWL
1SxTRuEsKZTuTEW00pOPGck2uQgTi7NI3o247yElB6g/DaBhuA5dMx93xjQIKACx
bfME1PHFsS6cbFV/QJ/NVHiGn8DiZpbtUejroyWvnPaT0nmTg8OgL408olDfwjCK
RNSYa1O9lLBrpCdfVecSF5Cxyhz1GB+d8cJsE9rUgAm4q1fWIvTuF3zAOhApkkOL
jZhy+OBshKZfUcTI/WK7vNhGynhvRN4EjjoQuo8wrxVDkR9tQFgBYuZhTX2TsmNb
tViVC5HXs0g1rQYuvXypGPj6DWsvkHwwT5kzOp0o3x7cVnGD5ZrRlk3q91Ezx5Qk
+bsYCuHDSCYouofrgS4+1JfhA7QQzVgMngNIDi4YEvcROoYTS6XQ0LLg1BQluys2
G/wxod2EJr8OUz65czP35uVI6XFypcoZcj4OWuxLVSvbWIo7zNQFPdOwKnbjvjWN
r/XdxCf16CPvTPzziqgHZi0q/Sck3MpfdJzlrfdn3xo75/iARX2D+Ay4TsAFq53j
yBgzk/ywOrzmvAxFy8UgVX5lngKxqdATe6dkhbohCrDCDt372ld3ZGA0Hue1iaDw
BacrGQ4Zp+87V0TCXg6XYC1wEL3ZqFySrjv7hgH7c9FgNpERLkxlqqOM1azzVG6h
RlmrcTaN5wfP/xEbw/dWoYZ2c759FIzsOrFemCK+/YxL4dBBGdUZN/MHJ7KBnNJP
i5+du400gzePG7vfVGFp37b8PMHA3Qvf1JHDeRRje7OKOOXO0tcW7WeAEa0wFgxZ
CYmB3qjkcZ6i856rnxnrMto1suD+cc5bm464/J7XYJHxEy6KjmHOUEV0bx9lT/o5
cMSKIHLkD5ICJOmtcIPgTafh7glU/h1tnsMeKJ4ZEm6ZWVWzkoeStKe4ZItDpAQh
8vWTYAseTBXYPi/CAZrokl4S5S+oP0ShWP9z0AK80KVfF5sakzIel1vYGsQtlIx7
lPljEOJzEbbOOhwZpmu4pYci0xeR2cUM6CtXJRVRKG89NtCm7RA1ha0HBjBGxAdy
tyiwVh5cLgKsqJc8FzNtVOI4vk1KsAwYFygL5PapCNL5LOGIltR0vnnOFp6p0rzg
LdfpzDnMZfr7xk2a1PxXn720magK84L097qMrF1reaPTgbEvBP4iE9fXiwaiK4wT
kKM5gaqDXrlANPqh+2sqCwLLMtHwX+bz6L4+oqmPTGqVQkw2NZrQH1AZ/LDzNw0I
yfGPCYlMhVT1mBrUT9NxqyE2FDh6n5iqSTlvS2feBDhnZWWwAMTlXWNTRuHpqkeG
kOA64bd2LbP6lYnGmG9KYCYTT+81U0Cx2F4kwA6y/s+fl7aFqoEJKrO2LbCumgsO
5Q5DrKr3afEDjHP6HPVO88624IFCfp5WCJdRrYGJgQ4WB4p1WL9TkZ8euF3E4ent
NdUEpwRTSwWBW2qKW1czFTGvGwUHlSNZnPtbzlu8IOqyGBv6F4xZYak6t8IOSurm
dYeixPY/A4UnAKPywAHjc/3E+5xGbILru9NIFhc81EnXm5PsparxPWaSMd6PP2z6
cuiqf82H9Y8ofDLwgDORG6XI13j+dYz1GUP2W0ulPWirp9+feHtqiDpjy4c3bCze
cRFjvHkUFvqjGRBJWGu52sMABkCmsNTtqEQjphsve8CTAzY9E1TsYvC1U5/yrwEG
BiXdblTiqCFllYc+xNsjC7mexMJiPp1I1rJcAgFG430W41WCFQixtAP5rJEDiSJE
6tvivUdB5tY1mr3RjQfDVUeyOL4iv6MttPHP7zIGjacQ+fhfAxgRhvRpUACCVGMg
Is3Q+Pz7FkZ/nZWMw5UPGdYxRJWhBbo0bMfiC2kEFZZjJQadPmiNThZVNtYeHN4q
BNLdM05yngKBsHWChJ7f6jI3LBuOzu0a5wTlO4tNG/SoiyRFqT26lIQncA+JvtE0
xv9bA713/Ze7XMJAx5rnV6ZSn3k6nKToiFzJDvtRP7HGeJnfTGqTrsMLYYaaLYA/
/GVUtOiBq3et84zgdAckHfZJl4s24I2tT58AXntEnuSobdGR60EPCgbxD1LWZYYf
62VhWyKad7yYiwW4UuSLXOcnu/q1WijXOSY8HEk8g/uulYTOJrxnoSavTMuXA2GN
53N9uowaAbqwihjjfU6xgaYIabDQWbIDhpU0CAuwQGVRPV4xaZtH/JdrYZRjcT9B
vO/7GGABY4DG36PY4nBiEYg0krzjAk0vD7SlQlsvc3RVBnJ0nkVlfSSSP1TLl0Hq
kD8TOcPYY3ZAbFwVL9AvBN5PDeyzUn6dsDRz9OnqUP7WNhUskGX4zOEa6+dnSNIs
JKt/xWw4xB121a/eXU4QdaFpy3n3qcYXUXn0rO4b2X7HX4StRkWm0WysRzLkMj1g
gucZ++Nb7UPTvJuhGTOwvn4jOeBR8nKJ4edLKNWYJC3UPGHxodna/44zUFrCtVlb
v4BlRed3AKtMdHrV88vqixAsTdYBJYNImj0s06O5cEj/U1G2GTGl6fTHU8ga7pqI
5sjZswnPzdrzlu3Nr3rd4NQsFd0dIT8MTWPfz+m2847iSmJumWrMf81weuqS7yfP
qub94+BBsAWWn40c3WgkiF8+jS4ZRwLGXy8HHcCoCJzL+P2JbRlcieLxbmBqSsjA
icPU0k4tfwq1TYET5XZxVsnxkZgET16BsTLl/GskqcKAGaMf+wB+5vBX17DVmo6u
pBkPjtLRhYjsFcbPDOMpgrRF6xnY5rUrvgIL4/S4hZfCyuVsOZd/vQKF8GIp4Yd3
/8i42CyzINKs9rqiL7A4pIeApPVkiwzU6tDvClk+8s3P6OXDPT/rv4rs+BY2KNqk
jCvo94jVPP1FgqKOH04Y6+aQMrSZobau0P+PmzRCinmUZ3dAYkZTkLR1XqDHuEWa
9thmW5/uN660G71W90IRREhrEYIBFmL/MPTDXeOhrzIFvU4U+9nm5mxB9ovD8ACO
5jjcTTZaBD9H6pPBVS/pIuDiNqtrwB2mhqc8KijwzUx4/PC2B+TcIcMVkBvdRUOr
UKUCylIqhZ6x9Vi7MHQtfJRuRSMSulS5GU5SY5a0F+xCqLpbSS1I2Dx65jnErLvt
WctLh6wvATPvVZbeLYFS++5wc5V9AQUGE0CayCdGKANoOA/+cdTsHmV37ijmf32g
f/wfIGv88UdcTGDfmXMrHkOsECmPafz7ddBret0UjD+84nNp3DYStDN/m+9KfggP
X/oamqVP4Pl78wRQ50TMelvNT5/Yrw29yWQn6J9ilecjYZkjl6XNZ52Ok42cPX9J
gD5thi3H6YICz2ZinpA1YmYi4bASCZ/TyC5TjLu9d/ZXoek81VsYoj9JPNzod60l
FQIj7Kq6dxpT1GGdbjGW3z2jSvPXqNYfV1/g7meh0OoW8JaWU2w87COSwqIE1FaQ
xjjNaIhersxzOftPtKTdelD5FH+6zwDxcr76ob4d7WLK7qInawir4jwxNlid8cDL
VVn2dSc4Qw7Rw434MDi1TR0dSxUPt0yWB0BJ04LC9wdeMIZQLbqyf1xiE541w/96
AgWaU78fNS68q1pRk+Y1sJcQQdYzQsGWYuy5Ik3W/srVcLD2bGjBznT+hTTmjkGA
OEy9BrR6aYkM18r+ejcDB1kvkbEaeBgjIq+w/5P5zl4IlY7sk7oO0eTJkKXFeo1F
mnGJD+c2LLNztMYK7m9kzEgYDEOccXNeTM67AC+vtr7X/iPLhdKixNj+C2QeFCfc
QOW1r+4wMB/SqCcdh04X0uZbuwLJVVKcRpanCG96A7gxLKSIML0hPtKpA0UNILsu
u75+nSNuMFKkmT5fHZh8MBrPiIEqq+WwYEk1AzyVjBZsfzSwlhWn815aDTquiv5R
Jehk4rZJP4a7NuPQXZDltWvv5VtLSLFaXBn9Y+ebXjHAqYihCZzOhPkpBkmUxHkl
W+c1Q4+YXQ+hzMePCcvb9DCRsLP0Z8O+oBogZGGnnpJ2jw3xG6OvKn6K2yKIwKmx
G79m3pDuaUh4sJujS1fF0Qiiy7MOJ3hotGZsDGxlq3KcpVl1dagF5lqLCtu2jyKF
V4h8O9xTPPxNf2zndty/PGUgLaERIoVaLR6hDy+XcFAMnVb+6/VofiPW5Jsb0UzU
6mhVb49VkjrG0ryG/SmdukEtiKDwNbDisDFhq2y1Tv2OJgOt6WXuFWELR3onQa6c
KQXy9xjenFUwcbRCai7h5tSW3lPJn1IyBo16gmCsSNWlgpRE6pQhzgh3/fga6Mvv
Mkjp9m8t34llZF/eb9cm9f8tsQlCuY/7i6zRjD2sUolWaB4bRWaa7uGFuVfQiD+h
546zWIp4MyudM14BxvaE7KoagZJLdZLYQmvhhWCzYxWkmi5iNtPgc3tsexop830M
OdrSEbjUpiWnUuIZ8eFgMYmpcpGzX2ObirHmAaYZuWL7BiUDIi2Mm59MexVYW18J
yz8vZVF1164mB6OYp8T9vupx6VQ/BzQLHZbH7cfITBt815COIN0pxnDxSJtrT1Cl
qA3yZf2BQsZ1GVMON5dq5hG8SnmZ0R7lXZudh2ZNgwxJlt9k55s/8ZxUDsFqAZAQ
BKPTYBK3QrxVKdwAd7uegYBB1Gu+BN9GaMWiYFUQPxEIVmJbYpDcRx7B5+r4F4vT
PProhUNCuV7lnl6xMT8AClTrXpOMowScsEHKx1Zt/djoAm51npRcmgOn3WHrbul5
FcW8T70HSfAjP5d2sLP7Crvcj85g4bREDYrnQokYNnD/AnGIJpbTOvVYp+vkHIpv
OMYZZS3El3Wj5rW3n4QWdzE/X6MdXDaqULLxokd4beV02WZXPShworCj9t9H5kp6
z+z7v608OsAlyA8pznTqh7mHvu/yCmDPxJqvBYGXDav4T/B5JNTsGg7pYl8E4rO/
jkziNvOUvk+SwuxWu9eUFkahI9IrDCj6gJ4KiZJfE22TlqhNt3CFXbR+O6JpOAoA
mvHwR+KzJXeeiRu0q8Fp/TF7JFE75IAcAgDDiROHMOU7cW7AmT7IMqkfphehzW+L
ZIo+CR1fm6uXj3F/+cGi/YWHvsjH5J2G8M69dORXmEdtmx6+XF4CKtsuA18YwZjF
p82xH/xCHqKPTI8cLXxhxZu1mXna4uwjpqxmH77Q2EIw8ZGQ8fP388Y5KpC4TJPJ
N/OYMc9vTDlZXnvoj/P6dPRLI/8TSz9nkAJAWFD9c5umgmB6W+AYQbvFGNTzXBEO
ojSBj3fQWwGHjgOMLYTdxgRJc10Mzfakdf58PsH6CvYTAg7slmdAiMEdswS6qhVV
3FJV3YanyXxm286/gaAo+YrrsdJ++1gmPwLVo5064ClZD/us/Ye3Y/lUdzC/p4tO
iBnY7m5P8oWpJOvva4PI9wm1INtZDyj5Z/ufhhbWSModjr8Ix/PQ2WUuFFnx7Pd1
juHRmuy0b/oHvf39eb6pOXWfs0YPd0/Je4e+eILU0C//udEuad2rx6oI6bwkrWyh
NFbYVHI+1u6fbbNiZr69PKn01u7EBYSnCqxRmqwS2aNQIDGg8sKYmiNeR8cVDTCq
IdKxzoOLWDWfWhqclv/E5EyXTz3jsy1gpRBRPbV/UJthVzHzN7oNGKnykYJsOA+l
vELxYNB9aEKM+LRWiG0sofKUOjaZ1BjbljBPxCq6H7WKJQ8YqVzAN1Fq87Cz7BNP
6Fck79xm/jlI9e/D3HW5l6rJq8qdaKvq12EsHozj3x32ac/jKf8gxfB3/L2M+ESA
nGYiR4dhhyZbJqLhmXYOFTx6KoNK7s9VDa9wH6u7LKYeGOFOEizSXKjZIVdwkM8E
+FqbiDTyI0azJuMYyOBVRlwrvTuoh7iqn5QDGFXNAOfjfQxNOttlqNros2wwHSjY
wj257RfVlnj3KyrcBqNbW4Ls9B+tC5wc+pYovQEkraGHfe8fPHkgfzycdRlMhpMe
j1pFc7r1kqGtoB1SXNONDYJfwmT4lt+C648semMHZvaBz1B1B7GT7y0Rp7n2gXXa
GgWLPtXsvz9cwKFksw8CGL6Zf1izn0Utd29FHXg8yG8O6iuH7K48EDZ3LKauwKoh
qZNOLpuc/y/ESuoGtBs0FpExMHhpx8meTOkdiM33MbTfVg8USg9G7SMHATcdyJbV
ar1raa4a9o2NfW9wHXLxrR9DMytRiC/yLU67O07gU5yMT6URrh2cg8qOw8i+gM5m
+H5izKRfsD37y5m1nkxePSL21ADsyhhNftte3ZeZ/E/9Rj033aiYMyG+ALBTcU1q
COQLszfv0/KtAPGmusNg5I3qfuSrham57v/vN+FGCTOICIUmt4DsPWBIU5Rdi4ka
2lJwi1OrJx/wGQR4McunKx+p+AsDO8G+4PqL89PEvf9hmQcEfe82K+gF4u6khorR
tXLHTuHjnK0MeNWqOM69NjTnrMnPqQ9BQMNmBIn2V3QwUxN0FDUcO94ngEZW1SiI
ATXVjPFTJPJ4pERoerbds87A9gK8FAXZr8BqGCG7ibqNFaz1NZVvdfhUg0MDKbuw
jnypfKEuGTstcJ7baWUzX+L5zjMzbj2ld7urtH/MUNxHNcxHbv5Ss5DQjqRQQPA9
IHGQKa8yjdSIIJlTR1ojNNyjPI28OuFad9YBxhDtz2TX+piRSCI45L5c+M11uqmv
0hS6ySjN6d9bfP5YrnOE9u5PqD/r/4iJMPoaZ3nalz9CcofX4EfhKLm4qI4IUtKf
ckShoZYiHJmhlBYl9E1RLfjMNbIhavGp5IT91/tG/4JlmBq5mUcjqJcGw0rElBTI
VXsHFxvq210lAOjPr2Tz2tIt+v0t5gqCIlGKLNUQhDX7A1HaQJnKE/KHF+J6UzBz
6ozEk9jEusWiSyjixCWFczVXopJ4HfNB8sAfI/itHMyr9QL/YIw/8LblklMRgyBN
oO50Zw4N8UWNLtUHbkcS1M5ZKvqYQCL7OxhxE72f9xgLqtXbBGjISLGdKtIIgYHM
M0yy4oXr85Kd7nGWsg4Jdk361H0m7sNJ5nUkBRHgkNAEPlgXkwRDJkTs1ITkrCRN
MQM77K6QTrQA6v0Rlxo2or4+oMKGuZKhCkox2GK+c0CXHe9ZPgvhec+2xtBhoa2f
Z8CyFb6o1CUUkPGyZVMUtJjLGklHof6Us46Wb3mZJvL23BW+K2SvNOXW/PkTuTDl
XQgiIiwKJJXZenyNLZeggOjzePl2Y4ZBi9PIRfa366js802K+wDdvbZdaoZxhXct
fibzBun+/rp8v9DZSUqC8aaDl+IVMOiblG5J1ItsU0oRgS77GG9kGo4oMQXBFd3r
abPG7TJ+9SkTJ2XyswDtt7Wxnw7u/DlS6MnGNkMN88W3ypJVhYpqTG9uGFu2SYae
tgfqg2/NKylIA0Z0cmxCvhRsQspbfOE+QgwgLZ11lLTK3EnUoJ/16S+k3fTNkWDE
J4pz5zax6iR5M4K95lm/yTLK9/YBKVHasSzANgi5FO0Lr8cbe+ZoNttPe+4Qpy6a
k3VCPuyKogSQh7Bj361bTrjBB5Aob/ymTU+Ih6SZNf+Nkgg1oVHToP44KekkkxWZ
akiiYYArhiDdIh1Oh55Cxw1qXZPrN5I5RmPS/YQglqtLxLiCk7ZO7gRx5IsQH2x9
OlAuJYo8FgcAcGOFjH8CgLLEZ4XNZJRQ1zKsi4r7919s0xmWi3+qBvFpTfWNrbGy
kiNrka9jRVAdn37cRLoXrevkEq/Cxhh8DFRLBTd4oyfWKuW8M8jBjhwWVRZGiu3I
TtDXQtMzagLhvS4SEYPOiv793wVqRDEJ/pVgnLz6iIfQxX4C3usPtsMCA8cvjh+k
f0oQFoNXg/UDqmfmn1y3Ouv1orw3mfnaTB8Vg1u5+EtvrfZfrvgl3WqJhEEtWEBf
s+sTKzhWgea4/HvR2irH8O+0Ti/5vw2HPG5yopKeSfrlAO2ACXCpP8Pt+PlAidUT
99nLjdvIRmtuXxlEzRZBCjhZGFdVm7Fa8WwKdGGcPH9+u05knO9mvH05O8PdCT0B
X7OPx+VFA77KIOn1ovDp2jytJtiblHUUfhpt6m5mWza/w2MaMql3fRrbGmirkYqz
qVt4FYqweVr+HZnzuBEWu0q/lL2cCvbHsMlMQ3/dtrt4mqhad9JbhasH2cUByOGG
S8TC49mC+acfjkL3GLNupS/P46hukRVxwQG8XitnjdOttdkjuEw1zgAq/sG0dtne
xbYAPANPrTruJVH4zPCpCQYVOfrV/zb8hvOL2068s/YKepqCe9EXFbp2CqAO1vtb
xrFvr2x2IsF3JjhBLfuDqGvhCsyFU59yNtmhkNx7ZgaKp3T93DTpWfHdf/Oy4kDt
DRPbw+RMaLdqwC9HktJF4LZI/JcFRj3MDTae6GYSU1+Fxb4frDxTzPFSJAlgjE1W
ig+QQvBvsJ7gtbPUhGyidTyu8l1WAr/a3MGrLlURcgwGCIQ2hva6yXAXuGLWlkaJ
L1IjsIOEgC6PvBQ5toTCqJmHOBChFgvoVB/ehjM+wbeacB8JagP8RzpMsn5hUHsX
wN1WFZ0FxiM7OHm9HzIIaOYjkAlBCYi2AK2k2m9YeGGpI5fiWdq9M5fXKDL1hUCF
QAQC0UkZPrnjquqltVQ3U0hQ+d8Y00lr+yuGfSfKrYHyWnYmtNq6ig5DT3dqm+vV
EM6HN64Q1TBEma6ilhIg4QVi+fkdNRQclHv4orK8NBwYMVCtHhPFXNyYivKPCvp7
+asBy7K9Fp1Qf09Tw4TEfRk+/j9WkWKNK8GsjrcHbb27j2c06WarFSfLOIYzurns
7nkYa2ShP5phVJ2btd16SPla9ZcnhI+viAUmSNzVeKOGC7itnfYV2yLifYXRiLbg
dZdPN7ELLAX0Vipf9efvNEEvBmHiwOtymZRQpfcs6FqTZQ23IWnaltMcknhem8aU
cIoPrRdIRlgl+XqeQ+3oHY8/ltgbWMuI0DUPz7Kx+PYpg1QegYD6ljMNB/f+v7mg
N6zUI9jKogfhvWPmvvShaKCRXC/gxDeLBCkzUXUi3lUrXU5wDY9o7lQaMvoeYSvX
W9gazqtcndab1zG7udFndgileX9o1R8IA9KWS7nldO7whenugS2AdYeR5m0Ngew7
EtPyuoKl+asducuTkTcwbUNYeCWW8TGOnLs1NYXmtzKSTjqKjU8Xex2mEIe1l6md
8Tt4pnJOvNmIweaHzGJyT12ueVmaY9tZx2ZTcpKg1ljCM9LTO2+9VnmuESmZWxJw
IRcNiQPjiLGJoyXO1NH+FK12qW3duOY7hMmBri3xoayAev9+GLv9F7R2EBWG5LTb
NJOldSiBD6TRZZjzED/bisqTnZ6yurGMbnajMpSk2M+fsQ/zzR0Y3ZDlFZs3Ftms
TaDeqtOjrP6XA7uDR3xPH0OAcfJWXl426poMDTwYmtdLBLP8Sde9ZDQYjgxtybTF
Am12UR2Sst0aPF5LPuyC/NPokyrFCQI64X84q2FCHsdfDTAe7ZB4kzZb7TRQBqLm
q57/tQeMzWvZiNz++kTTW7QBxeLV/VniDgwlzqRyH3DcnoWlyDP3GCCZVOcd6V8J
Ay2IOMVDvAt2MjFF6PMHluuO9gLEb/1eWq0zQenN+mbrfRtiPo58eS7wwPrITaHR
GboYhEx7oP1bn7Juq9x+eZDzzjyFPjFEDOttmSfqyWorPrsyiDkKynHtut0BB5vO
G7L7XBlvwX4vyzuDRAUqcvmLFy5rqaw2qv0vAiw9of5xZpY5Zct+rH8YZVZC640e
7++1fWWmvtC3gQ1nWfe2/FukrAOYO10giMmMVsT0tgK2CXKt8FbAskqhQnAcYUgH
A3VaMl1RuuVd5g06HjR/JhBsj4K5kM97FgEkr2BxRC5BbbrFsTyzCpS7uVqC4UGW
x3PqxRMRlhQUPn3OI1kyMK+1My7Bls5SzThA6eDSQHJGWEb4gQMCBUkuess6xvQ+
VR5dnp1dhXUoUjlk3mXlebHz8qws5kcaJkbja4MxnBjpDeybh7+DKRuRG8iaAT8M
MfXxmMWYq8Jno3kwQTE3ZfblW4zvGhwBu5e9HkfbcPd8EJwd1ElnRnLI+ek9Kp2S
Uvd8N7bxgOsF0P3hOzorcGcyhGNuD9Ks4MumavKh+FBK8ceyxNm/ysTf0GzVzIu1
c/G07kaIghnoypVGCBO4/Ww8t/Jg1zoWdeiDnbVlhuiIMsAJLlZUag9T13v3DIO4
UeosSPvOyRHJSCEqYbuB/g6jeGo7N0KVDVbxf3tyhHToP3gfQ78IDp3iqmE8FtdG
7LfTZTHiiCLz0F+jZ+FGa5geBbHUzaWeb0QOJFPa7JG5r/QwI7B/iGuOgXIWEN8k
05T6Dc2shepSSDmqKT+NCkJJzacP93FgA4bFknslWHKxT1ufH0w5NjhxOxsbJbuw
xFsFRyslWn3QqwAM2Dqcs5o023DU4TMqfLQ6JidZ0tlC83CofiYYwhrBt9MfRQFf
Is2Waf2xuC0Wg9AMjprXDrZyASN3iU6/BFWz0uA9RaOB8KlZsdliPCqQPSAyfe+c
rS5aBfEF5cVA2f+cy1ZV1CPlVtq5jHTjAmZurM9NEwGMGb/q3fAYdMBDgs1lKZuN
sVyqx/ulRxZjTCT59aKP9SFnUcwJQnNobRL0cR449WmOit6jAplE7jmE1JH6AgLX
RjBBqQ4XAHcoV+2Df6O0alegBNGsIxRPv9NsvuuuvpCFiE135exg3H5ERd0GsS01
VUiakRzwV88TTKsaMIY3qo44ORaPDPdXzZC4dJHcOJ6iM1/WjFYp22TlFjJnz+W0
Lz3Ufds32RBk4t2euufrpoWN8sMokVC9wBnpLlgQTtRHHEnOyxUuXPaBNUrdTXVr
yWCmFWei1bcKFeaMChpZfATXWF64FmjXJ4h/+dkASnOwhHfhT3mQHLUUKifjctKv
b4WDlHHyNOxXJESsrghxgvRTnKEW48RPL1v1wTrle+Xm9wz8pNHGKLYGyeknojeq
ZziaN5OCbZxUl7vuoXapZsfDkqhdDt6efJTV9ptRGdmHfAjGmBPMxTMbMCUTsSXj
Z2DtDKdiUy7x/fR8SjIhjRv7vogmBZ04DveMNevfJ533+U4XxV60KPS2wdxRH2lu
YsQ9QjTp9lxXsRzY0Zb1WgeHSSQykJPDEezdttZujFLyU5y9apm7A1vHTySaflou
QreY5ueCjkFOuGBT8tQebaFBdKJmbiP/AIwNFrX0/TyP5FmDuXv27hwi1JCnkQk7
WSk8/n4n4k42hrJxl2WsJ3xKKxvo9/fQBX/moTcYjIMTtXHkzsh7lKJw6gNfFG+5
c+cDs5vx6dv59d6yHTPbquSZspQOeBPf8F9m9QW3658Bh9yCdFiTx2TEgRSI+3J6
5H/NhehFhd588ODnEw9ut5HQJnSj/+kXdDawX7KF7V9/bErlQqn466OOh0LeE3Gv
7gvL1UZFWe2nn6aX7EDQhyyJ5dMu+uqnhAclmTrjSZRpuDkNgwNoW48TdbPPC+tx
k/FUgwUVzHiWehFoXPUaW7E+ysbuPASmjOIEF6YBTP1UEFpeaF2/ws6794hTirHz
TYndWqdqL5kVJC+ZA4s95Wj8CsBlDDxN3m0RR33ja1X5ncl1KxfiszUJ+cp4J8aX
8X1388Fm3Hz5+Fjzw2CKZAtTDt9Da5rEyZ6PCbawMfDuyAOWLIUF17B9/BSFYb63
y9QKdx1f828CiqXdWQFOn/HGxDiqD3cUISNa8wpp3XRp5zcoCXWx8Zvuh25ZDcHh
GECR1tCbvQII/t0v4J0LdczZrEn7YPTfnhsfv1AYN6jSDs7/YUCRi90fWAn/qKXj
ZDI5Dyjy82dDUWyn0d6oIR1qM/P/F7t9vBklZZNIkgl4FPnAwK/LouSwjbrMVc/E
djoQintZ79tD36sMB41gDoSwl2gXOrcTAu9ckJtLbQFw0lsl0RYra+Kq9YNE4atg
uTXkssOBXlfEmBf/AC2Fj9ni/dNMtwlwsjBofMbswOEGwUumwWUAwDFeUNq/L2Dk
vCAeIhfiyjbklTiwH149YhBvn3A5R5+NJbnJ8ZkzZ07l7KSWBYWb+8yCZJUFkKnk
wVV/JvgLOmsS2t8BA1FFO+ALy1UEayzPUOSCBhAFeUPEmkFeChMyb3T0ulXPfjqn
Z7+tMBFgyzT9VMotGuouR2PsjBU7p2g/8einVaT4SaXYEz/nmc8OIromOEhQIYRc
fKQuBa3hRatwTuWuWs58DvIdeLbnC57reXB49WF4gB0VkyLRJNB7qY3FwxSWzx5M
cFENLPuk+1RBVX1qXNcUvzygYvImvxMZ5DIeIRJpk1TzXeK3MNQ1P9yLkdHGcFYO
OjbCio0LSW7Kx3U+zRsxoGlpLdl4yqmOCAvIWK4ss/9n8lw2YO8riRnMZMk70bQ+
X96CqIZD9B5FTE8T6021LDjk/4QUIEfdTYWktzQ0g+LyHWXOxhbWwfDVfgd7dXb2
DWdnU8/bdRajiGOwZB8WxpGNZee+gPe1K1vs6LObjdzMv4rtg6zAGzpKTClayzLm
uEMGiwRbBYzh3xtPigkFENW6701EuTEM6Cyf/fCBb+akYBuhMIMPSf9EqzrF9krl
7c5EYzpmEcLoAzf1B3WbIMiqszm+g8j6KryrVuKq+tAqCngLN9tiJmcMhFOUCaQo
a5l8VMfAWXJFdOItJhwDgJ0pKlh3BB46RJ5w2R9UcPuius7ugy/td7BAfLmDDX3h
mjpj1BCTgfjoqBFf0DORr6DmjijgHJ95VKjxhs6qz3LFAX0QYLlvKZDMW18k/l0Q
lA9swFsloeW4ygJ3lQ0ATE6qgBQuAiFg6nzKCK++hRi4P/Zz2kOo6dPdLqzcxhUy
bHmEyhnWDNPbHra+OijJsBdZ5GVLzHwBnqO3HQ76lmaqRPqXoT5zDFbxGDzeNYAk
LyscIsRKKsN+iV2FaVa43GMVNmQk0j+rZAHk9BpPr6NQYz3+5r9uC1cBZVVYLieX
B+T7BQZ/Pj3GfH56Iw1+Yo5vpMpnbEOk9j/cJFbrg2qu7uhE6W8evn+YOYx9KYWr
VkjjG3wDxmAlAlpy1uiIkt5gXIgmMM2M9vtTrTRB1LlV3VikMvFr+TrMU2rvWbtW
ryhro4YD3UekP2kP1ijJ5CyQ3ALsODfu9VqCydAH6PgkFrw2EALueu1NMtx/jC84
eqxW8Q1u0UI+C5afGKCO/kA1DH7xGtJdm5G6JCZuk313I7bzg4yk4IVOBZVF7v/M
dKpLQM6nDifaKGzvPoZGwWm4VLDK9Vtdy4gtVt4HF75I2twFZ5y1rcgV3MIc+1QH
1iPSmHgse5QQgSew7XHjdy9y1ytOKqohnRAriMZY+kjYkti6EzUvEakarQny0coX
qQsOnEi067u2y8fGbWqb2MMsmX8T+pN5MbtquqlH4uTToN47VDFgwWXSZZg+33FR
upv60t9rBI6l6EEK0GjKbL5S7fStLCj5pXme1dfUq1ySYL3UL5yRSaUA6//wYY01
piGV4iJX7po621AlYc1iB1cAM1ZGgOakssSjVgQmDTYOMP9WP5tS65uNo7mB2Rwe
tQwnW5WzTgQFLXx2Nf6gxF3H2dn5aliza7HtK++snZR6QK6q5PFS4L5UxIlX8nNf
geXOtvLzWLojJCD6LmKgeNKVp29XB2eOpjhCNNliGWJdbtyI/ZeRwt1rkOAfvWnI
gBVP+bqoCyeYMWY6KKmpspf9+69VOnWLjrhb9ctZC7yyZHze5+154CmC+8UfIVcP
z3EF5RvxDrR8fNLux8d21LeBSCOFnSKBtrFUh6HKtJbHZ7jq4aq6vwREUIfWs2XB
FpmtJxP7qr3hes2O4Wszmq6xbDsP8yQu9YgbcrU84mz20jLEduzJfDU93lOfCOHp
Pc25vVb9n1LiszUSDshouPE6C1KidBaOqZJEuARozNESW3Ri3CGN1PMrJbq91Ajo
o0az9RDJ//1UeeTxucOlOYTcVXDDqtfIddump2/Syc701UDe2iQPQAdLHcYG270k
eH6Spdoqee0KgeFj0P1MBHxq3g/uJ5nNIrDJI4+9I4z97aDJBuLsWce3spgNIwvK
5Aj3rHvOdU3mKCs8dazT560WmDwgysOtK16zrSS6JxNfBRE9zhqbVqAbVO+bwwlC
/najc7c3fzsHh9cSEeG3cerYF8kp2cqQedd3+TjJU7HWkTuHVsQQEEQFJPaqSDF3
H9N0v3erokVts6Xwgvvuj6mftu/ZX2HeJL6nlHub72QLALd5wA6gpI2loMkxCczV
/EyMSMFpFWSnyld8QQIzVQAXxdpDdNrtX3fnW6pn7YInOzVFuHdNVMuhWeFfX6Y+
6t9LAcT4gr95Y/dthaf0BpsS98w5DgR+QyVJXB3gH5q1pnSDhKKbs46DRsPAFiZo
wBCvXZ4BjQTv/fkTPodT0ugdbiRxCuqKWsqAcTEH+LRAEXlRkiobnGcLDuRsySMf
pTbRGT8tqclwmpo2vLMKionR+E51UZRQKrrtJ76e3a9SRaR/3le00WHXBd1QI1BH
8ob49fKPcHBBqHeIJePi0yS8PtnFfJ8Y1g9e7mCCLPy/aCtjFm92sE3FFIjSNXrE
fH2XM9wM5kaJMM/Z8nHFBOegUQ/nwhjTAP3/m8UBBzrQpJpzx3fBnfme3oVVyL+V
voCnPBYFJ0aX1S6EmPxNX5bQBB/+8nc0CnLNqQ7aI4TdTZdUnd5YIhfYbb21xKLx
91K1w/1BpXci4PVfU1yxh0QUFCBGWfdUmFz2z7RegaG2EFDlVlM/oP1AbjK7klMa
ULAmfOhJwtUcEeYk8wK0x4PEM6kk2+XxAZo9cu8WTpC3sFy6gn7KOXBni0ZMo2CA
Xt0LSv3IBx1Wdrz1B+ONVA0RmCdSis15aFYAl4NXFYQUiV/ohWqeAovn3sRET8w2
EwsM9w21W1+K7i+iomTWQWPSN0KIeccjj8XvYtmaw9IG4WcY2XKRvphbXA/e8efk
20hqd8uYX48FSzdKEGRwLxtHHMpGKiG0fap79v8yS/sZXTRUBp9FzqUza0yHS0f3
pbv4/hchLAGc23DrKs+WVTY26g0kFQTnUq/Vyv0W+wpmJNODnFOLX4mJLwSgCTsh
QSh8zz2/yIte/s8P5s/7gJqa0JKqm7Zb0I0ACUC5eI9GIT+LG0KbshYHFD/2rRPg
BeoIUlbAiLUcdP2F/2VwyNJIKb8imu0z3usuIp+zG8LIkeQomesrc3FsEm449zsg
Owo6RHragcUv7Q2j+T7dRo7ufEpn5KD9eZWaTEitJdT6MFXwJ1yLE+J6gPO05qS/
5EbrlnLmAahlHOIV7A3uCDBrHZjSPx2lwkO8VDCghey6f/HLlxUvbA/QhvqQcCNd
sUxRHIikoJnn58iJ4ryu8Zh2n3N8gZb6Hg1d8DvTxwc+Pthvbn6+wbOaIoqu5cUi
EX04VqbAKRQ+FrQlIX2x4NhfW6MwH7/Sd+awY+2ZaXz5CfSP2iy7JUuCB4VwE0hD
TAzJ7kyF9jfkYGMgt0BynktW9MsNdNrIxqfxVe5w4WGSbYsXYLMhLlYKbHOVc+fs
G/3JqX3yw3XJIC4kEl/3apsoOzRfh9xA9w4aJHrGEtSZRhdpVJ1AhlHrNX5P72IH
Q99sxMA5Mncn8sQejZ71Hb/tRYKe3bN9y+WaYwrmkogaipMrRGptgma+FSIcfHVe
VUU2CNjkUmhLAwKsJGmH4dP56TSvkNllIVslmSn2FpZqOPho56P1KrJhE0YsJkvy
GDZNXaOKZXKDH+T5XD8VToJUEIOgioSr5fyWsihdzG12a5SSa/B5uNiXJELikosq
OJOzokYenLAcM4jsTiBeOgYHEUy2GXT339OWn+D+i5AWm+SczeBkIYUILnWZHCFf
UKRMLDg1jpzf3QAgG3E9m+u6JQz9te2PmuH43kuBYE2Hec+GWSO30wwnhhAj2jRA
ch0CfkEHhoV5CqPH8XVO3hDsj5KdtZJkBnpNYh6LzYLPAMcsbJMA8Teki7GV/hxw
/hKhE975mtHYZ7bX9i86wSrr2P/VPAFUM/YMu8uiZdUn47zQaMscayoKvYMnWRCe
lh0cVBKrdr3OPqUlVcS9zig/eZ0ixeHN/tyd2yCMezSA+ebtAsDsubM/AxPt689D
KG18042XJTyBd98KRQsjB9hZZ45bVrSGuGJxOX+6BvSF/nM0+324qAMgmoUW/QlM
evjL6/aD7Gkvn0d5b/3KDrV/kzHGR04JMfSZBMIx7Xm1UrYo605JNgXBfkzoAyK/
0gYkkw9v6H90yIs9JopHZHaDUW3a0n3LMs+MmBiJos3evpYxRQNkmXuXpXUSKTmW
ebH9TuP3/OsrYK+q8GoBgCiKjfaFVyyw5aNHivmzCqo1mYAD3NrCnLEGoMF6tqYz
wInrfs+khsrE8P0s9LTw2r+w5u9lxfg3Epyg0rtsDobgofOs1sP18NpjwLlh3ipq
YUJNhYrj3OvKN+CZZJ1lHfWguSOKrBJUELUSLeCtU01r9XEEF8YxOiVx2LK74NAI
hKL2mC9iNpMiewaEWhBASgVHSSSn7l50mamiMN3lcqAJWhxsMqv6YYF9E8E5z/Po
tMNzND7/it84vc9pYGN0wKjTns0yCH9u1Lnv7AJohFWZbQVh/FQSp9uN5Eq7pEBy
ssEsLdP1qZID1Gwp7PRGexP7kjIZQCcF7nE2cKIXVL8anuGiTfE63Rl4kCyfotEz
QcYhvVklAjSKfv5Zm7W5u1CzPZfIlJGVtR+W9TFYSKm2/UMgOtx0+Atz0hGyJaJC
dkE8oQf2c+eHwbnoD0TWK/XtMhXcwl5N2bU8ZB1DnPsgDYeAm7tHCPoxwNLvdJ8l
5fxfeB5yNs/j03JaayTC6uFucvWClN36XA80mKWAyovoiMS3UVzTE4pu9gDEHcdB
QNi18WVfnB87oN+HQE4DWBbOOg3HlCFBCl6eyT+k+24mNlT52PyMqGxY9pTPdJAE
uuOvjLxKdWH4v7EBWz+o+CYX2P1FnkP11RmXpEr6LFBnBLh3Cu0+25vEv0P4jmej
+oB9ianfmF3YWwd6muszx/MEmkEEYXxQQEt49dKCIoWE51KuB98BzYkhTKGep8AI
77aw5wmc5jV/CC7ZerG5gLNk1BkF4y1He73fNDaBZc3l5vivZxmJ/ZD3Qa74R9yr
uhMYf5sgaIKJNvVFRYcjQwWjSDJkQMKEPWkIGOdnGe5VuNrtvb9jcrHD8IaXPrBQ
ABc+AGWM2SutO/AGOZjPkPhl5IVArQuzBEJgZXfn+aTAyP3ONAL2x1UPYN6cK5wb
+d+JkK0okdtFCm1HR9LNz5Urbu0jfh0O9XQu5NXGZ//u6WFLTuNydJ1K9lDeSi+b
eNZWyGAknWfi5aNE7Lf/64sXH6h+gnPcH/mY+OQhHNaDhTKzd3o3ZzyCRub+g5jS
Wmc7K4Ez9UM2go4kEpF8TLzgYsv3vUTCqCeZwDORJHfngUlst+umi+i5ZqlEdM1V
3mZ2KHiUbhMNdl0Q0lP1qtPBz8IjAe2sYzpA3ZQKZxRWBWiwLQYH4KCH3Pr1CMIc
em63r2nakcijtGCSUi4i1BdNFHP62+kuqysOQGEH7DMuu9BSZ5+QWllzR19yvUu4
of9/jev/LBBExuRBpNWyA4+coRTedW44mqGGYbuEC97saH8E9FhRAi9V7AC/Hs3Q
+fLND0pb0Cj7ygyv95xdsLphGn9X5cNNa4MIM1dNPrma9v1U22hFKWXyMni7qpgp
Qk09gvvy7+/GPEpcHFHAzzgG+PZ6Lf6ZYI/ntf4XQzoJMzsTuX0U1XGoG8DLoifV
8cbwX3QKaPE+w/SKqtqxUZuqfyS9IGLgCN5cqNzT6/9+AtXING1NX/wcDrfzNMma
vEpz2ovmC/ibKUVrGBlhKjFZqDXzVXOpGe5fS415mvEQI72Kv1hpOxP9c7sRRRYf
klnJgMKWAclimalv7E5zLWEDuLR6ibGOpWx5TkGKoQ/TgKqYdF8P4spy2kI1wmcq
tL7eoW6b0r4cSWrJERF/LZKi2SVrVzsE6+njaDJD/57wv34b0wrFeUAakeeflmwx
0avboMEsFGEKU8HfuwZnRc+Gv2E9mt+2wjT+Mnyi1oicKq1OZZ23oU+fowIKxjim
GuHS2OF2fJ/TsaBm9otNVmWDxRYzJUY7tYYVbRqbHPJpCkO+MGDSBW1XRrrRvUl+
kgWlVWmpkfyasMG/mCAmt/DdFEH9jZgM6KE/HAW+dOphcWRgp2bKpEf2HEq5a0Y3
N8a/E+3viN3Xld1feSHK/aoiHb3eKHHqaRYBi7vhhPVFO13N+fOpxHph1QrgKaKy
ZWl68IY+Za2zkmGoUiKYyjQgNr8q2xbrGLK5d4AJ+ZktnXrv/yMadxDwMd4BibXK
9hF+RZKETFxfh6alRh3TQ9RzP1mdF7nY8ZX1Fs/nU5Jkx4Tl8LQVbHm9QGk83Z0R
pTvZUD8r2SnkptdvGh0wQoUy9atV87v3Cgj8U4VBeAP37pUBkFNGfCIvU1wwKcG8
mkH74enU+qi9ffesP4ZNVlZYB2W7VERGz8NwyrpuwqTOszAoxRG0trN7iGuxkdwz
DJXsUOpg4u6vdA5yzq0tjkt2RMYDYrS9ld7Ze+yX1zRGELJb3k6c9Oy22VImlfch
+2YXhGbbxwV/uzUiqTWhXGoTZ40rACLOKdhnyP/oCxpjECzis9TZe6JqD3FXYZaD
tnydC7sCz5xTOIYpSumhaT9HMfJ2wxcphLHPSHrDLFe8x9GdYtsaVD1AjiuC9X0v
fXPFcIUBdGZ6tTIJKkWFIcsdw8EZeO9SxwJ9ZJCNHO0EUbIHBfrS2wN7IeAhjlDH
UhFWg8XTlUdGxdgByrrnb2FXtHSOEdze4xgdsfAaFrg3yO+c5IX9XEpkXieTUAn+
OoVZ7Jb2V7dDTx41mSKw9TMRCQrb+IA+VYx+jEKxNmqYpRbhwuPsNsLkRYiZb7N7
HDOpoB5JOzUnIzdtsJ88BFxxvZ+e9mGNb67LcNg7hXuiHrnher4EinvLypyrfphZ
pEmyT7dc+uSteqLQ2XNtSvjbAgvLMG2CtGqecZQJUHqUxHvFPSlCyX3DVHzBQ2RT
efGuBHCA9ymoKEN3dl1B47D7tAAUBeQ0ReW/XGwx5L5CFffcs4O6EAkMTzZgRSad
uDM5wT5JHZD4BB0SE/VlnVmbYJkiFBJg9LrUSN/OHuDdDyv5wuoBKR2QdNIOSBKl
cbtLghC9bNv6q4f4ENJkubNyY87oCATcmErk2FLEUUF1Ep1/JhtorqzFQ8WHVGjJ
D1VN97ZqIPKiwBpmWZkpulrLaIEvbrR59c3RrkZOBeSZFsdzYWWPxjlRZclB1MZH
rqbRVkz6PElWw/8tJ68RH47PVMvjGEdOy3BJwe6AGRuHsSZB0cOefKGBsCjRi7Ni
RJgMoskIT98VaCK/dP7M+w1bCrW8qsHs+ntKodeMxcTL9BPsNIFnVkTa92a3qTCv
BLU83VDAlsMUD3p7mP2w7fKGQB3A873CQa9FBouid+p8XMWDcgXCKnj9PBn/xZYd
IQebYuPBG6NjT4hNoUIuVqJ45A6xA6Uwvg1wiTvOvG6Zav6eIKMcqFTGAn1/r0M+
4yNWqYnAeQcDNYhjDL/tYAloevzad7TaioBCVKkt4HjYqdkI+/PDUwIHrvg5889D
T9tOR9vBkqFq2koy6O3Zu2Jv5q/87bocnG5rHekb5ENqXZSgT2p27bDG+T8UCis3
LpmQ0GvS7eXhjI7h7yVCC9NN0wEmaxn68mLRiyAzgHjJqBFQuFl0uv919qQWmzxG
eow5b5wqBlFb89JypVcGIF3l2AB+nGbudySH1NhqDnV+7yzI7bGVc2bVOmtTAAQ+
76FCsbgzFlkQgOwHOhZKJvnA/HGnPJXG45taxNZNpHu8Cqlo/6SFo+Zeterzqtg6
FTiQymGABqxIl2PF0+G7gWr7FI1BAyZeCA1of4OkUCIn5xa5zOutDREM+GNY0xVf
eoEgtXroHVhH7gLexAsUrtxE/q6jlUVjSsHvEL+D875ksFCBZvG5HroWcm1zkhh1
0bvLt49nClk2xIrgH0MwwhjBRwLnX/BE46+lgMtLWYBNIoVqLGOFgMW/af7t3UQa
RCHNTIXhZGiU8oTlOgUBs3mpvrUO8UzQ5hdPcH4A5F1m9rlj4aSYswz2+fLgU4j7
rZS18U/ixUAQoFdEJpyZIAW6N41vtP/wjIGSzwUn5H6vbh6yF2hDgozBYcLK6Xoq
Ra4TTsG7YGNaC/YfzH6pYUD6pgc7gY685Q3c9GT9HwGjRjhOA3xtClK1VIFo9hy/
lgMzTBrbcQELZdFkYjeL0P+kcgkmfU6vzFE0I9eRpVlqBW5PveTYkgs8GaIdx/0c
p92PLb6mtzhz4RGda1auxdgknm9UKvMjq31gNeu0eDo7QNAlqXd19iCbdDTnE46s
Gr0gI1HfZqMCG3oH+wkEvA7xb5nOLvPhcFQ6mZDoVn+ACN6UazqM/Zd2Py4HgzA9
pt9natprI3Gx6/MxxbWIG8w+bpBjc+K408LqOffNCr7/eUx9+fQiKFf6yPNyn6rd
mbj6dCgvuo+77ruvkFhDzFpGyBF48hDYYXDczYY5H5yaHnYFW3aJ1FN5AWC+S1e9
UNChiESo30nMuVCmE3LzMdV22cVRF8oxwsMEdmkiqOQh1ZNk5VRIgzj0cG6DgIRo
CY9mV7mHuEAFETgfcK37rINuEGj27iPCA8wbI7Y10wYLHRYKXeWdi6mqA7N/MKsb
OJ3dA1QJ1zq3UafibImzDDAmBrXnpuG2+Ann/j486+V7JChhpgAe7kBvN1RqtnBx
2X2eOX1qd1zuW2T3wYUrV9x/EYM0OU+ugt1l2yFB1qfYsvbCRC2JxY92Ev507kKM
YOpxl85Z6Wd8DJnFDphQfJEysgEOH7risAUhhT0GoaLZ8QZP75WGcdEykEa1/XOV
tWnJ9oO0vqHmTTHCAWgYeTkxqzTffZOdnwYLgiSc/HHUWQoC+WMJ6faP6IdQUPIw
9lFl3oQ+X02yY9WsQG4orlutdvyeVLQHB5Na3ygM6kFhykUlVolmPmtEn7G7brZt
yXabgFecLyWz9bSq+H9PyiMHQUq3ox+BD3y3Gum4qpzRg8C/2zTTsKwKSWCdf8wP
iKK+Cp7Cr+jc0LQhH2fUolgGsYHiTYI+ydlQVSIkJCOwWDFFKlhH253+2zO+q8NQ
I/BuRKFvk9+Jj1yoEwIuzBDzwsgZbg67s2bwFzovTm07dGwO04dqPnp1BDZ3Qrel
mz/VqOm4RmYX0yy7KXMtOs6l1q7yMhDGz9HY/yrQOUQ6Fhxqws5ZiA6hSO7G7Dbj
KQsbWn5O+RuRSW8trySR1aTxh3qI3DX6QIlI72Z1WREVYToG5lgggXtVZG3m57AO
dIWCj+TqDdggHcSYKXQ2GDutpzs0Rw/u5Ita2UShXx+cF8KekqhnLINSQu7JtB/n
g29ROeCMGtoUhtZm/YbmIvi4j0rjk60p6r/DjorFmiIz4aDFtHRJ63Uy+lDSiqxd
6nkzIAjVkYj4WQsquQRslCEvnb8wp/U8SbkdQpkgBwO8yGYYs5RC0lWmVBgNaVfe
RUYwpZfj+w9UsYwUZNoVLiYjUaXgUVJttb0fPRkbxkW2iPvPCrm2SAbjwPOy2k04
+N3+uhRBJOl7OOpLKp/m3HK3J+tHyn1qJm8OfkVQD6ygKEBhOJ9oRAXyTdN2xxcS
K8qWCVqAlXQC1Gt6EacE57vRhvCCQnWJ0kA7HtKCKzpOrJyrjzAZEEeBvrX5fsH+
ebvpEEdjmWJ4YJDyXorXgCTM/Yw3eVr1MZYJDWudD/SwSYZR51035FDOxST7gNc/
8Yx4Cu6nojjsjfeJL67JBP5Ldi17/2AEUgMGgsrc1EDAnn4O+dEBfRXcSK36Rhzz
j+NxkBg1rlg4yH/otv0BlWuZA5ofPVZ80Bsx31mIzD9VF8c55FR9ifIk30BPf/Hw
tracF54AJLxVu3d/fR0tj9QycoGEi1IRtb4W+av8A351OjiQjGbVZWI/ETCyp6BX
3tdAQoakIE/X8bmv6smDyYuIbKLT1EJFoDsADRWpwzZb5RcKxMKRly7G2FLjWwCD
eBsyv1+IkXEv1BLHA01aK7129fRzoXJLXGnBN22ZPyNB0MKaiDpGws3wZ/l3Y664
xvvsjREPErf33jtkykNyiwI6wLLj7Y0tqA6gyhwATFQySfF+LCzhUVEwFh8FEQlr
QYbpNDzngJfYcyx2ms++s1U0n/iCMjxkAOi5abMr0Fob6oM1k3Fsm4t5b43MD1Xg
N15QXW25BQmqtMJwi3FfrU7v20bySUBLgARklI2TL9HxoY0ZU+cC6K/fiFO37zMS
A+v1T5wymvYMEPu9KpLzd0Shn3XXEB7rtTilJ1ZWDT6bD1yyGDvtVns/rdM3aGU/
8+uI+XjzVdFIJWqVRLG7EN8XQE1Gj5dFCdDsbOyDG3t8zAygclw0BHX6bDYdUon8
xNrI51gtocMqFmaOivGG8JI0DXJh/3ty12shknQXYL9odKcGECzZxuQ//5miuO+b
9aNvgJYMVBwdksAk34snyeRwSxkJRWxIBVSx4D+5NjWjUnJxUH+/M8H5l1UH+8EJ
/EzcLVds2YfSPcF6MPel9fNxS5ruWoar1oNLLc27fxU6i7EXmxBs+13OkATpWC57
z/n7d7ruRYAXJcgFWEOJOL9EexGIggteJKwMjgmp/ig6Cru4QxlUGM1fn60/jkAt
7v484YZV6rIYojIetxXyS2sRjnCyEaxZyuMqNUcsXREzhgVUkuEt1IoW9eFyPQEm
p0vlIXJ2CIinAW/hFi8hhYvaVSJ3pPVERoI7hixQPDX/ph/NMHCJDn9HGaTtT6ba
a/NBQ4JCpWuQI67llu2aShtKtYUqPtgN5y2Z2nJbKzWIyZitkAx1THXEXU48xCC0
WvoFk3Cd00HhPniP+OnfAOamMKMqoX+K5gOmZnVo4ip983S5APPQUU9OV8KINhSd
sUSoe3Jb1IIQ9je9hnAkQH9s+/9JHY5IUMQ1oW7NWSGHzNkgYnboNq6zACCnuHbr
zowiDXgKCuu23vYGati2Z+0vE/ZJf+wnfOc+qsjOgmniheben2YX+IK8aJHSB7oC
ihlRXVk2f8ESVm0xjeNbhjxG7uY7V0mcJdmf1m2QVbruWgFsRQDhkye9108jDJJE
JdJvoCcSdLKMijbAETSZh2Tu9aKXh8CKpvjPgjCvYlEMrfWYCgUTyW6zD2+HPAnt
0kP/GetC43DRYquWPV+pOQw8ltNYnhc6SIrlvmUyg0bESl4RQRiT8C9Nkkp26ujy
ecM44VfSpvA4t3/qt37n0eihr65i9D+X/lFrz4E5SUe+MT9VqxJQToexLm9Bj1UP
P75UW+Qwcp0QatJNuX4oJkPNnt2wPXewPMEorJtJS9TvUtAKrQiPqZIr+drTJ0lx
l8atqPQAr/ErA2QR5lDC8fM2uzHyrX0/TiAyNVrMN5l9H0bWOBLu5eAosvL7cv9M
EeCbdovCk+vzv/ok4tpehpWmlule7L+uDp8PGFWe+T5NtriHsEiS+pLp/hpwxN5H
e7Fs1zpKNaHZ0jJTUDJp3hx2rqmQavgIdP7NDYAIKXJMYM6XDUO6v3+teQbs0s2z
95/YeNVV2Q9THRpvUaHPWIOaSOcat05YD05YT3imBvLH6+38fR7H9ETIA5EDmcc6
2bvslJOKGNtVptnmzI3dsXc6ENozUiD54p1vPO3B+sBH0TKnrZiJmeM+QxnjhAz0
xseh2nbTwogeo7EmOo1ovkk7c2sclcU4T8/IT8/nwypcwwL0lKYagbtr2X+SS+Q9
QySIPDy9kMSMyOGHjQ/c2uH/7QU7931dFeKc2hO/oOvpup3/1yUY479ToGorRtJC
luIe6uDGg59M3u1yg6VJOtxaxlOT48M2cKYPorCxueTaTSoEYHA1hx1F8Ium9zc1
BF2qqMKODhNhWOJkwHASgOQlNO2NseROWpo+t6ItCJM7qE/02dzuLTODgjr8kwnU
lG6aMrPg1szA24C5lrx8zs1VoWpA2twFdMQwdl95TO3ryJp5h+Noe/Y6isFwqskJ
tWmDcmWizdc/e/ffybTPNG5bwee5fTb5J1CA8xRQkHeBXq6gAOCj1DKwTg4Xjr22
+MPD1q2UTpFn+4H6t8g7JD8Fs+xZBa9IvalbaBllSHK68pKmVzGOprjxK7GKsiB9
xlrSuKqwFuKEJ5prGbv6X5WlNjJDQ01axRRYxQDf9GNj12Mzwxwy0yWXV3NSKDxL
WzY3AnJ29Bu/baDqmWg5GcjvC8sDD7YHIQYxYwiFODY9Hz/DRuhUWiMA0sRuk60J
B1jLuLv+UP8cdUg3HnS3OpYq8ktx7onQpzVSBOaAoio+r8EmtZlzBELHzsFcYxsv
jNVFryFJunsR8Ro7lxn5jTxyznOCbKstv0Rh0nAmnZqvOSUSHthnmaTwdoBjGGnW
6xmNN8b+I4F2BrtQWkmHCv0ZZxvgwW4/KRSLykZ2iH4K7xkQ8wfx81mbChIZ0Uh7
PuXTe16AJiSrT5TZU3SYK/eoX6caLl7GVWnwd/ERXSG3lXfYFYCeevz1Tt7Bzn2p
qF2caf+EuLLEsvB4zfODsnIsgpRqVhZLZ5U/hEUQjRM2B73RKzjlDJsP1+utucsY
dqAVMejdDm/Gk0MpFk67b5dRmozW+P34LlNlYevUXv0lHvsrw28EWd3AbV0BKPQv
xG2kxRYnB2nYEL/2K/2BP1mMyef3aD96ib5+ok1fDMONz3lSNlCdlQJZmNUr+98G
3FzxC60/eEZ8M72WundY939xfRAFJD49wLMwFNWkz/MaH+V3ydr0RNlJnq0J3GTn
FXDJJFH7f4687dIKuWdD63mJcDAU9bdsaI46OYWS0gRB/jdavXVRyCJqruS42iia
Lb3i/qMUJWC/yWa4FS7uAuJDIhSFYqwF/Ut6Bna4dBqxry8JjU5yVEpErwl8X3EA
R8rsu4OU61wSxggKCnh/53fNeHKm4tR+3IRjQhA87FkBzF1TyuSooZUCmUPikrcI
Opg6RYCgpqz4lZEPj7TmrXy25vhReyLyfzmy/lRZtdWUawMPG6uesHxC+OProF1Q
NMXjF1IDlC+kpVyg0RipHHy83y3J/z6JgBM0zXfBWFc9Q7mdYsuazPl8HiM94oNA
uhqpgF7gMgYPi339x900zg7Td0/Gj1RTrE37OXrTg49p54654Zs75RfNsY40LXab
BtIOxnfKu6LYsDkaYQWDS8l4H0BVWY6XXYHl/8pzt9KobVOIuMbmfPCL6xxrHS91
0XePgajDdMZcRgaN6DK+dKU0k2RxjfjkPKBb0+sXn3ZVAeiDGRFiQ12WoexRdLi1
jGqGDiPTM6oxWKgqNEiUD56Qc+Mo+8ampVFtJJXQlyMCAzX/a4N2ZDOAsUU6i6ka
1ZTz/8MQgpiTrx3I9Vxsauk5ftsONXedE+9FPMsKbZDoWZx48laQZobNUCUgFhuy
xBkuXxVsPI978pbv8MmuC9Ek4WPkhlbFOdIHjJI0qnXFH0irbyXAhbrMb9gBZqmU
gr+95lQglSPgJLv4mR10Tj2S5lS9NEdTm0L+kc03gkbz05DBsIHQ02dekf12jIRT
VFL61wYWZWwDc3E8m+x+fzlJVfoDr31Ku2FsRL3QIlmkkNEpfZD80u+H+2l89lgv
+jzkBXdKqbOTWeLoIzaA6IZ9Ws/XczqylW4pZ7egRAuCvQuX+/ANNHo0Jzi1jy/L
Up2NL/heeGFxuyU9/0f8c1RGfohDG5jYJtfiVUE5fBIi3FLYxvEM9QXwEwH0uymU
CajfZUB8vy9lmY94dgxZqUf1ztQ7Vyv3SqVfr29h+jHS+nXJRQc/1zQWODYAgN9e
/I6albGLSLLq+5TrLuZuqgjiJ0KeFxMr5joQWZGAOolA1K560Nhf1733habHqCJ9
n7yIcwWuGajbzRs9Nmzl+npvugieWvnTyTiuYkhADnYWGshtnk3tBQthbgd2Z24k
obmtk5nW3T0EVC8G98sVW6YxQlpeJoDU3TC2HT3lY8oWHHhp+yevdW6Ae7CVBRnA
CGpge6RujOFh3WRF+U5RMmafRK7qf1aJKrBx+BH/nJW5EfUY1xGZk5u9W5Zfhgqs
iWrII70VHVDe6sqaZmrVpnpayrc2usOJ/6+AaAaMkHX+ym4KlNhNck3ojewxk6w0
9a1e5z3PsOix4oPSmZalXo5i2A8bhD4Q1nJEjFe+htV1HIsBXuD3lxauDYWyCE60
sQunM4audX3A3edcMYb0L20VvUyk/NVMm7Sv/XpYV7d7ZffkNMQkihhUFZIA2QJF
Zy3shTY7or/tXMYmcgmdJB6V4NF0GnBEGejdmRkdvS7Vgy6jvWnqc4/NpOj4Twhd
DBftfJPG3ASOjf2vtCJSPq5o/osFw6XU/o6N5FqOtIBqi1Y9nHO1hcw/P+rwn9sb
7hLDfXppUU0mJqpxHUDNQweLJqtbvTPSUFHav9r3TcJn/D8BqyzqjvFzDyOP/PGe
xPnjFygj3AJ6OTBJtxDuJj8i1qMxgrn5M6/t3IrOSeHyJMoNx9OwXDNBHp9PU3pO
o0VncJTQiGkSgN+vRtRq95XdeZPKfNeS0B0bZ5YjltV8fhRYhmOqXM2nUxUoeEM0
gYis41Q2M1Fz17QOENfl0NHwf3D358AaJj8V2fDUEPjsgzraml9z/INETT06HERX
q2f9zUDmrFJUOPZ3mXu9nY6dpD9e6mf6XLakwdU5pzfwIDepadAFMJAlPqUGKRZE
X9IsUoOXcGIZM5OCYdFDkKItYX3MT3b+Iawf6ChtOb2uZNUWT6QtpghrHrROTphk
W7ecOf/GjFz52t75bGGbk5buSEY3IZmRRQqOLpLxY4WBa0CHM+yg6OzBp4gqSLnD
bCjnMt5N9eIONqnu61r+MJ8tVrXViFLn7Tf1RHERCUTxiLOlrI3c7cYV7OGIby7w
5ioHNwn1By6r6WALiB75IQGXEQIef1i6+uYb6enPLIfFF26bVVkQEHf/cRhZph87
A2wy+Py80vq4i4e53r3J9kbU2jfTfixLUhM54Vph1hKxeB09gIOjp06eKSNk6mnx
2006BE0Yi9D3aUjlyjc7cMXyta7dDPC9CVEpqSrfSbp05+KYuczKQP0b5b5dNN++
xiaqaPqa6jwac0YphxVJCEhwZp6l3hpcKymPnEVvVa145cXLNHSRbuJ/Xpq7z7Lz
iTGPAeo+FzxTyPjLcgfxN6zfRa2GYp1EY0hHL+mQDlu5siThzrQ7EGysDghcvU6J
VOmoSisAjU09/L2pETAY0yP8pGvhNdOaEKM3tPIXiOTq/5ioQVAEg8P0Bx9sscgs
AJxJFMO/uBnREUfTCqZNgC9Jy2h3NqFPtdDOcyPhrqyZPcb2fRsdr0YSy3aa7eGR
NCOz6NQ47MbuBuyUTtzuTWf4+Kb4cidj42EtkcP6+0a/F0e1y3xRyPBwogxl+Jw5
OTIze2E+H1VSDA3wW17yst6yYDA6ZkvZ5BS94Z9JyN/voFyKCHUUXoLeCT/mRMCJ
DPpseXap4tJoVGb+bnexvZ6RjxiEyrkWpNUsf8+Ss/WEuqeU2Mml6p9gxI0Vb04g
FAmreCYVxP/QmKW4QWWuwH2jQJ8di9zK7FpnKi2l6EQFa/a7vRSHFDqK5/l550S6
Gn4R6Kv3/9Urfm2Te5N34bFLffECUNe+RDd5NgCuoZ5Wsni3FGU8XJM67s56GzKj
m6ilyDaKfezKUIc04iuAvqvqy6WrbtCAdY9azxcMZc1df5tSqS5MHP0Br0XUTD72
KsVUsaHLkhMKYGyork1cLQmXCZzuuESun1fHTatMRQ4oFOwO34Vz+au12mnapt0C
bYMdxMWCBKl8Nb/4mdDckhE0e96zqlwj2dge2NAUhGIQDjOP1YMsdSDWwAVYrf9K
rvWuvdZR3eraUYDXXW6T8hIT47TQp0wj8vXjiW9YiKCONkcZNzZxip6lwNUyImmK
L3iTjskqu09Zq9YQjo9sUemQ+04JwFS8czL1np5GdjLXwMFUCd6DcgfzfnnXZXmA
gSa8k5yT4ZF/Qp/3Uzqud5H8KK80oKedFusudN3jAKPXA12/cUEfB7zSW+P8owFG
0hCjKohtuEZPxPMc7//Z3Mwf95hwL2qyfljUc2m3b8M5FiZHU9px3WEdc30+kwG+
moPaF6dK0e4nXyo1T5m19yuntMrxcg69zalYF6JJsM3p61Xv/aZFUeldPYR9JSa/
2iOKwFhg8Lw9OO0FFeOKLITvK3ufplnNGOw5u136sEAtbdzc0xoUQi61BzolqA/I
9Ff80MjCT4016cAtq5g6nDsXe2SxGrMejUULavh4bbBvc7P1/AgGuhiQpXZN6TbZ
1xwZuZP1jo/AioOzjJDGwlZlWIHBsknJQ9YHnnbjTMaoTaLLkj0vkVUxFeLc0v6u
THg/MjlHJcZ23yBZnONJMH/cN46zblHKUF4BhVCKEHbdPQOWvZSnLN2/UtAKVP5I
lTsCV2EGsbnAs335SFcNUDukfFezOJOFeeT+Ff/fzD+pxSVmHNVOm+MuDBIcn97F
LdAuanbX6q3nU1GGRcBGVdG3lQcZJpPq+cV56TkFZD8ILRoqDN+MONw/9el3GgEd
PJ1h9vpEMWnTpQKtFaimdBE2rU76w+EPF8cYN5S5ETIo0jrVr9uGhePGq/sGzD+l
CUnoGDNnmYOnuF3rsStpR1VUBjWjMjxK4u73kvaWnWl+GzLjRwQIQFQQg5aTh/8c
v9SDYHRQo2SqL81U2OEtFc+4/lGPCjXbQENZkfxN/7zcsg/FDMZj47gxiZHIVmWB
stX8QCFJ8z53eQ8kbjfchxl2UNMg8Bq6ciQPRXVvXAIYehpiyGh03IHl3NSwP8Yx
H1krdLAXr6Gbr8Az0KsgLcWLAKifAPSDXAx2/sMRrOcCIRex99MQTFWRnno+MlQW
R6Q5rEZniGj9elYslgrdHEr8Q2eqZs/Cj9UOASjrdRKuuOyb835uxTqqovmut40b
FequBQvVFNt4bPX57xoMJ9k0Ti/qIruaNltGamTxI1UIlQfxd/PSB480rJHQJMZD
OcPr9wjN/yYzjgV9YaVh7G5BllZF8S6sX8EoU2cjc3SAqsd/53nCix16fGijGFKa
3EzEDel6xnn+p2BTLszKZDM8T7+qxd6U1NkJU+rCQBomlU3Rwn4xYru6QHEu1oTD
n/Bo4eywby4UT9uenr9iXMKsKwEata4BQGlSe4GBbLef74EpDLSf3ntnB9tYqdET
LzVEybjoi0UAlfHf9ynmSedJe0VLy36HaZx6zlzfO8UezMu4L+53vEr4Xar97nkd
aSOQgpG+ee8cjSKCWtNno+p87vaWMUhnejILdWelOwbkzaYdO3UgGVRvUcQP4gYb
p6AS4mpJYWs2Kn+lFpAPXQDB+aTl+MP2s5fy3rI9EO3ohKgVHVPJNNwwj0YZ1dZn
f9shWaXQtl0x5eZuZgXttHtwIEhwOF+0pj7EUGduHnwXMh27qo/wNRmimFMrxpPu
tiRCO0xDkK26UbYwnKBLqLDoeQZ0wmXjrrGVJu60O1W6hY/Ui+6ve/3eaRdOKwMQ
MwuSiC/2MDIe38Abmja8pcKjyp82uWkT18fnzP8QqBC/vvQL8gEdW5mVLffTxbfk
0ru0/of5ytetaAaa1ZiOh6S/S/pAXhtXX8ACoY2RVgzyTCmBTdkeBgKdYZaf/aLI
lFCZLBaYmaf6edW73oS4VXQcELCQ+82xUBDU8TJWLoK7ZHr8Y+Zoat6G+CGF5fH5
ppVqbSsDnLc7deYk0Aobq+DoEi/XnPoyeDAl9S7AVp+M77v8df8c26/WXeS942b+
gaz9VwWqR4Qs5F5gMKOTv0zf8ZBo8+Jh4tUdYn2ww1hCw8/EvRN61MqKTAcP7g7u
ST/SXjBxmknmZ2zqyPYOtLX9tVwqPJQ+xNF38eEsQCYrwuLc/cpBUkbrF9ngYWjd
gzyz7Dy1DW4mojqwe8aZzSbmLaJS20Ley2ovM6iYwWfE5+538yZVVunq8t4sUl/d
2hxynSBD0POeM7NiqmzINuzOsL3by2fkJyfrVLtaQNrung8Whre+ABYDVDxZuOYK
wesEPSHy3GwNNmVoqGcDL7/qrmMj/apmEYA+iycN6e4LJyVJVsA8fanVZmP2syp+
1wS+QxcjfUBFBTg42w7UTVUTUHgarNDIz+lRr/onabxgFwrKXPSQItmrocnANf4J
5f/qydsJSAIT3Ch638KGDg==
`pragma protect end_protected
