// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:05:43 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
AtZsjGeVGXyN2C2AN5qeZSUuXjh5w/aJ1nCgXr4GpSQ4qWPDnxtvsRdDUyv+WmIh
NgZBCVW1z/T69jYq9OQcaxSjW08A8hgFOEPaRDc0BHekt0jwNHpoDCnt73OZdLc/
54jvDwF6WbJsPRKjF1DYEpOwR9DXCNPh61+yaiUEhEo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 32800)
Jcloe7nDU+OA+Al18xSViaJaRuIoj5xBPucKrElXZRVc/fnGx1SizqXsJttgzrU0
bohzuCu+ecbaUnrpDKZknMAJgcj2y13sA2st0Tdwipj17Yw8XDLaM2XgIHcTFTBt
aggipaM5zACm/uyIz2qtZKSP4havyE6w2MAyNWEknrl4pYAoOeEsm/+XZemTI9Gf
KcLmytxh4ab78e9xNxNFZ3wgIOkJmQ8eAjmEZn0ccbIuI/0Y33ywOsXFnyJ8hkGP
tq+/U7Np7GGtLyfqTg4PPRkfCjpXD32eZHaJvP1XZFST09/KcNNX90Ab6o40g4SG
f3HOqoMKHm13px3WERPepZTjVViQYTSOZ3QLwOcyNeX/halRz+1uEdcJwhpnLTfb
Hi1sBZmNabVuAdHK1esIMM2K2TzTdnjTGy5Rb8ZqAA7iadyWo0I7gx6VSZj05OPI
IPzE6XCj7jhCTrmoB6KLSwRMbMxWioIvr9uzUWDQKz6L/KvTOTjZdHdNZompMozM
XjHjxxbwiEF+yLB/sHUuvCNapaGu7GQqu/BMz2RosNJpT3dUO5lonLA/zp56WeWl
rnDJfZR2vXODvAS8FyZSwc7yXUvajZxDL0znCZ86Odc6vgiWCvfTtZDc6CSrt3U8
3M1jGPGFwqqa7o8HMPYBEI4eNawZQtooUXoDb9TVtm/QzB/DtMkxfM5n8+6h4MV/
d/YBb4LvbtNofPVlgw92KIJUYHifPCbbjdCzduSvFvh9JcUVGdewYISzPCXItdHy
DoulIs8mr8EvdWP1RP1/QAq1VzZOekl779KVRmRZHIMhAxCYABqO0R2f/SwrDNt8
EHIVjFO91qjksKFj989Cz75A3HoEMWn8oOXq3IMvNtVmtkGvYYrBC/dWvmth4jgc
1Ao99czu64wspoDupNVB+Ttgrx4PD4pILQqd/G9eGzgIpNY8GN2kwBUDTr2ZervW
1sClLRYUFUDXVfri3cOwUvzP3mJEP74A3LuLSJSQUz3n145tBw9OpoFz5hpncikG
oiutyxcEs27dqlUSVqhgJ0SJNvKL19dWGtbq9IPcDnIU+L5dr6anmTohEYzCqsog
zZPMjgRj38eNXRvBByth9BjnCGh6nbiA6nTOVvnZv2AKGtdv9oP3YHldIe8/gcy3
LoE4sqAstwmKak+BewbWIjMckgYsySJb+v6Jdd+xZhlP16N1DdJy2W4QFaa8sUvs
BG7p52Vp3Zgek5aywUe+9AzJSsMP6uQ1SGYOwX9hE/SErESkvARZzJra6g+cWt0W
CI3S3mdylepjYBun5oBncFZTsZW+hvlD4sZ2HpOpc91k42aW5Zadszq0s6lXlJos
jF3fzn7Hb68LDfwiCGrCmj3FFAa2EWx3fG+aLHbS0G0cuLFMGWAJph80SkoK2nmX
5W7dG0gXbZrGP3ZBgM5L7sNikMbWsyKf7Nq10elDu24MZawD/6vveYXZkPNbuv5s
dPkaHq2Es0ct3/NjcpM6lkNnuY5Joqs7CP8Ou+7ECbU+k5Uf13jiryHTJWw6JGpq
kGi9EMwcZdIp2/wbDgsyjz16jG6ML3z1MOV+XGDTHt9yVGCt6tnOs69tBy7zfqjM
7hO/G1M4iBrehYpz+auJNTR20CTSKgWDj9xLc/nEutXAfuIt2AWryrS3vDFuhxK7
POF9XEDzANF4uMI/nhdwo/N2fvTWskHKdNDEE742zrrEp+r5Tnw9W5rCUyjvQ4Re
k7j2HKm7nStdRqYivqAjzmqJwLCjwrHloJ74r/QujHQEuYm2yBCvBuXfeQ39MENz
Rd/7tgUjyfWQUHtvR2y98FNcX8lNlphIArCG/2BAsBLWh4VJtK/XRxgYsAWhlwSI
gMAAZmPXGm0XdtgayYlXdrG9g2oWLD0IUf6zQEsWJcLIiUN5oszSOf1Sz8QxWqeU
HvSYkis8KQ7fFpa4QzQVA1SpI+cA5JcVbMoTG2lKVguG0YcxMrux/lNIZ73A6Yul
96aKcgjpp4t6LbtLry/BIg42pSaUm89xloJzQ0qW+KMCnmky8EE+6nLgZ0fGx47v
A4ET13EuAJNV7qwdj4/C2Ypi1oZ43b3sSSrLNMiGLG94oNdmA+9HBbhvm0Vp4K19
FP0mrbzpjyUXwVzDNqlSyDerOsvYNItj9rq3h3iFr8HZcZ4LDayTTn5nnjdBFuku
y9Y1nCbRGly7La+5gmdac3qdvtMOFV0l0ERMPG5y6hX3gHJliHiGGvRLoIPV5ll2
1ENyJHNhXwXTfQUfHpeNHbgecntObsvRKVH68n4mJmXkbuSbBpcYW0GrAhMO3uXC
a982EeGM7IuDR/a5EjRUH68GQssTTQHBWoBz8Aa40t1RKMcvC9A9lALRAoqJ6LHP
59IYey5XPyoKcBog1OSfEgyxqp0p5uWdmOnddOjaRDpp1369sW8szoaSF27JrOa8
RpuPXA9K+Y016gQz1h2tDQCdWKzvm9gUR+13TJ4NtPZNFu7PiitpIqVD49OTqqQz
A9famO5gWpivlL1Re1RCmLPjcJJf7GqpvlhFdlHCuEBtBKK10mU+C3JtjnC58R+C
5At2ynvf8YGF+eJfEINpR8VCXU2u/wJ8ppXMqDPoQQrIyH4P72DWTdczRIPUPX1p
OuULyHlcJlClkuadu3nbhEkWxCtIqexMg/glyZ9+Orf50di6lnWopm2kEOn7Hzav
01047a3TvTHNjxsYunT5yz2goeyepw5wi8NHS9PBvWZYlGKRYQBDCBcUS/gkqO+2
a6ym6c4sC7ozVmusTTSo6EpR42/Ne3qh0EvPEV4xuLKz4XRHSAcW3t5rRjFzGxNP
KGTj1pECkemKYtBJqK6QuvuyA6/lOIory1TmpcpSusuy5RwgCIFs2Pu+03EfXGRh
TqfTCj5nbwVT1yzw0KajYNusyNBcY9ty5fW+FEB/MAUZxaYGsWHJIbPBx01A1fna
SM/i2jQ1ZP8K/R5WpzoPfNTI+X54YRfZYz8cEoI2NuN3bxGRhb2IqVOXDlMpyKc8
oW+r0Psfca+4/rr5BFb/keaGAQuzHhP4jOP9zoFte5yzTT04gC5/N8JQ6jAq6iDV
fJp8BCLUBOpzylihGooS9XEvzafCbaktY78DNdcodoynt6xDF40gEMh9Gkt7HWZv
0aMnPM740SN62Ct9XiWRBCL7MW722cNoGAfVdn1Or1tOjOX85Vt10sjFT+BfCEz0
t3T1qL+LNWHqKlS9vapYeA5Wu+vZxmHtv6WRGE7PWTQGNJaGUY7fUyvZxHf/K1pa
kHl2Pzr/cBUkA/nNk9jIWs3PFTrSo4wpOIXSqy44YlQW+A+X3wXm8O1/qpeByPCO
/FZRf8KxweR7ZJ6UIH3n8O8jqwv9CM5FWf16Fpdxkl6X6IR+RANtqfEMDyZZfC8f
vHWQx5su6ZJgWbjnYURDdeVRLMv6tIJHnB0X7s0VfLXL+F5ISYa6ba7uGs1LuGHS
TPvGe4Nn7k5ze0c6nq11Q/Vvj9GmoPCZpVa2x0LH0wNrqE/zmGnm6phj62/4s6QI
NrrLTNbCEcTOHQMr1DK9nqdh0G1DmpYckOXksYYOgAkebEodmuUzm8tRF+TThe9I
1R6xj2reeEoe5JxzOo/2NBh9GLUnL+01p4ikQTKVLM3gzxqK5omxi59Ob1kfYnvG
gDobGezKTa7vulMZiW1b8eQ6wNqzYqr2OsHVJXHrfLp7b9bWcrrc0jjB7xyERLzA
a72gxeYeQKmTBH3vviel5xUuLKe9QWciSurVbgiuvKNcLN2sl0yHKCTqbRsIYtV/
PM2ri5UES3tr6i+HRItLNd4ATYR1PLXayXC2BhXnw0DiAJ10C1ZhDXftT+Cywih/
aUv0BOzBj46hsFEDnAuALYKE98JSQL+2bT1WaTnaBW+/E3RZN9MX5q8S7b241YG9
mdSwkuHOwyjU8N9gM0XlvqTTYfvxbBFDdwXEsdz0iw4DAvzOy4qoqHgYnEobCZ5d
isUKehrf3vVQ+38eV6NgjfrFF+ke6NmxqB714Z7b5NRiaD8OgD2KNkjcYdK8MTZC
jq6M0uxqqvUvLEp9aVCK5x7e64OOOp3VQ0FE3cuSYp5ko9Qx/WQXRY4jrakqRNn7
BMT1bNgd3dgabfT42pn+CMZbb4yNeFSGDucnwgU5GZQrjsEzvKrrrxdvHaiKUa9K
zbrCP95e8orqMEjltuJWAnX7SvCjhLBhY3YA9PIFq3w5yEWgHGg79TyATfXNTK4R
5MR5rVztDMIn4SGJ7vRiPdd9PTpjLAdh7ubbsapFeE1VDmS7ybpy3f34X7XZci2y
bGIzkVcrQ7spy6EWPs/SHPokPnQ/kS981sQwg0EWklm5qJs4bT61SRLq14FRbTU7
8l/hIqL8F9q/MzFSM70K7B/Gyz6qJiGfEpDg5bsVOK2YnEiYrZxb5P3hyL30nJri
9uRc1MTGydMJumLtnpphJ2kS/Qc610zqvahXGpm6agNgCPE3LdU4I/TDPdEgIy9H
qrOqXk99npik6ZzjO4pwfdLlc5N5T3JIyf1+nTQguC4KxN2a9y8+6KKO/1mKeFGS
+wRgjD5xUbeUgJIyE5y3srBBItdj9wyedQMv+GOECDvqZ+iwxOYldBOuEp3xk8YN
g+yvzMjh+yYvyOmIEDXgjUEMwiESOHMvTG/C8ri36zAR87Eic+4H+60MG5jIbvAX
p+l53p0PBLcq+XH3cz2GO7gPTJQIYVAhSX63fIPuDbZScRvJzhqnzy1OQFo222Ma
yuJfjdrTX+Ek4aucD0H37LpygyJoHaGDtf+WkFCY32CJJ7sRZ47Jb6UyRsysSJ2L
c8XnpdaLNWsRZ8hH8q02bWPcuxfKFvQ/qKhdMwAkrEiK9crrTXX3kAcg/MHzOs9R
eofB/roXJwBzJdgQNae3H8iWsMvMxcP8cGtxwcuVtH/0gw3QeURlYwT9USuG5FQj
sZ58u/rmeNyVXWZbnoqBS3XCuzu20Co75v0cIU4rQT6DKTs16GgVbkM4PmfS7ANR
8JGB0lslUQPUqTHWOkkT/bZa0jJrX16f5Jri6Ju/+lkRJ6ut6nxBgjTTMqSRhYZA
KUdRFMCNRjcPWSwWmel4Hd1J4JFSF/2lmpCnxZa6Sq5XlZkfnynVDUqDWo3hgzEn
KcZNlb23zJ1nnNILJaPyoU1+ZPUx4SwBNwB2jyhA9YTh8H60KuVCGExAcwTfpFGS
4I7Zn9gYF1BOqEO0dlWx2ELDPAPJrzRjrwIUM9dVXVQHd9yYo4eagToaQygAQ0dc
cyjQtzIdO/e9WyUGaFErPSCUaSH8MwRQ4DMX1ehvZ3R/c1Qp9MAAdY3BNKJ2vkoI
Dc18kEtCMLHnDEEWMU0ayBYwKVK1EUp29qEHA8uWOOmceN7Ff3Ll6R9uTaZXnX8N
dLOHyNP+oThktWEEyqqbKRyNB8m7F2ySFiZoiB/7vSA1FNgmmP6gelepjrX0O7a9
iIx8gwghfrhdbleoHPnMDlZcG0j3A+LSu6o0Bk99VjDX7AqccNL6XFp0TFHcj/1G
rOS4V9wf1ngTbbcwTHD0X0cXwT9sEnUrQqtqysFWnUC6s4ORCuDwX6Oq4UYrLnM3
TXPbXZGQ3bemsDRp/PMmf9K64F9RIBwfaUqdamL+/AZW6fq0/SL+d+Psbc8Re2Xc
BCUVFE4NagchQxQLBedh4ZuA56vRLGbzK02R5LvXS2/h1G9w9fbx7kclSTBZ+hn7
iMv/FYHUi7pzCtiSMLKlNzoXbqtnuK0Rlpc+WVn19cOm84xJXX5tCwkILEc11tZj
FkCoEF755ah8+BCaq92Od1b1YZ8aZ3NIaru4gUY7sngGMWtDnlpg6CTK9W7Ur/5n
TNZs0+QLof8/VfXCefayeemcI6+R8PbwbkVsPGzZ8a2rLLoHjW9xw1QG7PWQK3i6
iQBckDTUP0Y1K46LSqJp5SR90iqx5lftOEvjjssbMzqbLBYigEEOC5FAfqXthMI+
n/1ZfSlM+gTQ4uPLoG5mKkiFLbRawWa42QZ1NZ/gL6aLvoxvdlqoiARYeZIB9tNU
sUgNYc1KC6rAJ2pQuE0mV9tQpiB0GZHTDjMsKad0LGoBJYDA+9P1cx3b58z2Fb0F
tALEFEtZPN6T8C8UXiJoGeXiRn/S6JKynM41HLrTrsRSN4cy2IBW0stiWXSs0eFS
dgDhAOc/KvJos303uw3Q6byflve/jfvf8mxg9OGP86Ax05fdUwtgt5KPigKEKUor
CTLJAjO/TJnnP+pDfUOriV1P5V+R7v4BMGIGMOCC6Je3VdSJ0XWPIi3yNv5NzqRi
tjRjfNpy6Fs0OGg11Zy/cXeVjIztPoA0VPvN77ILke4hZhR2MaCFOt/RFECzccSd
ghpU5SuFNDj4ycBpJeluCmpxZsAeiC4oekkcXzQu2r5GaUQ/CsP26uMIoMa5UQc4
w5UZrK2gFLfWqiS3z4RKHEEc9NMG8u3U4uI0rsgw1yV8d52K7RQebC7gORN7JOVs
Q8Cr3A8r1UafgiXnIHGLJoUi+1IW50MuOfXJUGZ/fuYtLSJC1c8PkngwwouIp9Hu
HGIiP6PKkZBprfKwkmS6azves0CKjDMAUO08yU1QHQkc8eMeYFTbRVbtsxce2DG1
zxlIFxYjzSwUpBD3d3ERnihUjGit14vCUpzCg6JOWndRGcAFsIY+4og6s+Tr6prx
QWQicYSLCA9Bmk1ouz5zEdXLG4I6XjcLeQlm3Is577R9gZPKGdxl/dcI3ZpAL1ei
qhyag7eJbgxWowVY1uabqm/rlWFDTNS8y+zAf7qcBPhZGzEpAOR/V+VeZYtD1pTc
J9CARYJRVCt694DgIEJ8kbwosR3Md0voyZFdxt097TJo9+91aPCM299xuB6lxImf
TdvwFolBSi6JlA/7pfgvsLGBZbPZuOe0150MOEojdC40iWsw+NtxHbB6Hn0kmJ1r
ZWyHm9oClm7ysUrDcBiK3OzAlX/vK8a/LVE5cdMsLAW3FM5Mg3uE+8iwkToYckuW
Bj3M4tGBZoy1Wcddt7q3h5pm3d7E2s5JCJiyTIRd0DQstjdmwehQ7VMosCBQxHs/
SsQZj43yUfB1CQfv6XRs+EKXCMbi6rKR56oU6b/JlPp5Ipywe1ECgzd30Xgnphgp
OWuwyUCNqOc9sB8JLDfjs1g5qVR6U9O/wmmAv68nkW7hoIxJL6aUj0TLVa2VG5NO
OBFiNJ9UQ+zufEr2DX7muxsOEZIPa4Ng1gDiwULero4Jj8JsK5j215SGXt6u2UD/
3/Qi4J2pNtTmCtUSAyhU48Hg0EYsFeYd7GXuRZWutngg4D2MgSeRK1VfvRGLlagq
fjpCjeXEXAN9VkYIEdiJHosO9EyLpkVQfMQ8d3SfLsETgrdiDMaqtjn7elw/ip+e
xNjMjM6ta69VHO6KvRTmvw4CwZbjnVd5T6m8HJEwJreOdwD9D+zVJNFinIb1nhjK
7MS8W5V55ChefiFmbBgap6S1egMf+OgYAog32/VccFW9aIjY/t1moJCIfLtDqUZO
dU4Q4/SPQLrVkV4wqh4NOCbfqk9D8rfdRwhVIrlvvW80s9PGiq26oVuZdq+rr598
pq3ybCUvp9tuO5qZHGulBuYU/iMkpsmpenb7092HxGtEZmzMkf3Ubw4THKFR1bNr
1V/7po5j8rzIYpntJd3k7i7kNuhCpMeuxrV7rtlZFn+8mjGTkJeXyY7z+Jr/oroP
s4Ns8H9alF5Nyei6ObeZLldTGfFCbu3zFYijvEDxk+OP8ZfTTgwS5CGvzKGlb5KG
KidHOm7r4vPwLceaN+3gJmKnTimva92ff0+DqIK6nfL3Z4BOhcs7aMALBUjQmiPZ
cdsdDXXb0whi++yO65rUfP5C9z8wbsmCgIHmm1W2Uw/CcxDkT7C6VqqbJfN8iDNL
4o3+OEi0hC8Iby0kKxDF9BPEod9gdkc0RhttvkkvzMvn5EmLYYxETpxm5QQ/ow8E
GChDa8exws2J9qF+6vAf1nZiGhw/7iMQ9JtcEIxN1dveBxFUFPZ5vta64n1aBhlI
xFlZF1oQ8k/Ko9Cbm2xDHph3x2Mhz0Dt4iCUE769fUPL1HaIDZJdedrGTz+Zs9PH
vEnmeSD4H/bXZhHsUtqXrC/KI/JJKlMNoL/+OC53m6lqax0NGRZajDU/e/l4wAzd
Ejele0wkIHZo93Mkbx73zGd0Wq8M0KQcGReX8iFwiJEhW6pS75wrwxUtrAroQ5jf
v0WBs9KYS5N8eK2XbPQxCW3IyvRTG4ko9pNyBToxZYkUmnSh6zFgBSBPMYDnIoA/
3fJLmviKOwSF+s2G8E4vX9WxJFgVgYHZzEVrMEV6Ig0qM809WP/qkaQ+SiDWJIce
99e5er+O5Ihk9g2l4fM3B/31to2d/fiTsiTyhLc/xieWI/aAaEn6sdaTza77fuJe
6Dq+3l8UpQiOXj+v+MX54LNa013Fowg3B4uiTfub5l7pX020fhsOo/7tZJKtn/Yz
BYvvagDQ8Jv9uZK7GxS3T8kCECix2WiK+c5TT3UVMniTcC9FKaG4qtK4a6cfBkQY
/+WHA3Uz7JXSdE15ZS0S3Dv2r30FE986hxLnION883l5pSRmalAShfSI8NRV8eIS
6h/QTfnFsUF2NWTRco3TT2G95HpdvO2UihTIp1bcBR6MEdII580hIBUIovkeMo0M
tB5Kn9YAfG4vV72e1QYbeYpcq61SVICuweL+4ZqV421YPps8Bx2ZBHzH2N4nu1S9
DrmIaT2InD1NHqs876mPEfTSX1n49EuD20m4kblxJyIxV2xU6Q5kRbKhoj6iOtXV
0WNATe513C0NgNQ3r++qkUdbHh+6U0EJ0sSVmhDb1E4sOiszQwl7xNH6o+qqQ1Ae
ojhQCTFKP3cSE/cKuZ1Vx/D7LexMOfZc9GJqbGXnInqe2DWBWZ5edeDAx/i6soPU
eSBVEpvQLYL7WqQqV31RPGvTNlUExmqG51BqaqvT1FmVvmJ5UxhOKVU+E4mlfZfF
ERFVR2M4ZMsLy6S71TXKTn7778LtgnFgKyPoYAAP44r+ITFWMfjB8T8h/Ijd4j7R
liqNiSY0dcw6lVnUkGHUN7+KsMZLc0TRRHGtbEhGAKO+YsaRRqTyIEjse5F5n27U
W9X7dj8YheTnONwJ9xebqjEJIWPKuzQy8911s7goM6o9fmw7hfMGnVOirnN9OFly
UomYaKUO4IEgDPQpVsXLG1jNcE7E7UpDTdxt0EaabmmXrP7fjTtQwqDSypYHue+I
RnSamtjIXOh/AQW4NuDSIIvdCRN/g94eK0CE8G/Aoz7Fy4C0naSNxEIoQCIA7sqC
BUGpYzipdx3yvwPyPeWSH7QcZ9k6me6tDPwUAF+yzjUi1nXpWFhLDWMI3HwMxz4+
gP2o/G5ufVjnT49biodSEMoFDg/zx3WlGbUY6+Sezdex0WlnQMzH7jqgm2uvqiKi
pTWPWM7baLgDUzXBtHurqnG3oYhA7KazeG4E2qxPBiiotUOQBGBc5UAqICFyAeO8
9h3MCDsqvVCunrt2STqTyLs0QwdC/qkkqWU5fQ6hn/4637qmu9fEe0LL9I7kMzwG
hAAM8ZoEzLKBI89jv0gjG4ufAtr4SDq94AR1+AR+IC82tUWO8HshmaNN3RM6g1bX
2Y5fS2iYI/l2z42EjkZXCX7/NdGin/P2ajGF6S+tw+g+TSh1Rhh8ZE9xY8qMARgs
NsFV6vAlvjg8LovFZumoltl9xhCdUxfXFBysC3lFIHCtnXNQxnaAOu7N8YEktJHF
DpThSK1dBSXo6rdhAyl9JN34qfygqHsCpJe+Ug7j/PRWmApF4IZV4bBbGqwOyCrs
Ubqg2fO6KDK5w3eIsDKncsIDjmz/BsIMP1MRyLbF7imWg6QOBnnSIpET2Pz02Kik
tzaXGF8IGpnZ2pSTySGa5MFy6h2BCcnGr15o82INUV4WsCvKn8yYDIGDpshN9MOI
W4mkcqIM6BUIcdTtIO5E6JsfCrPFoTAqOhAvzhQ2A9K23whuvroDCYBubeHs90Mh
EtfPo/E2RGnhS1nlExAhvWJOtRJOOAGFR9T6/xkEWjzqOAkISOPX+kiKm3xa0+EZ
NDl6TIi2NKE0+E/5c3XTZbey3alDmQTtKxSAYlah5yIusP9ZxS2VcfmkfrdUHtS0
QF2zDIzHe46woIo03h/MZVLfFCIRM+7RawvDfUPRSIpInU2OxXjB/Td4IY1XWLnO
rn/Tw5/ZnLLzQTrt+fvtXN0hJAUc3QhbqMAt7pMkVQRASqEJhjrKGI+29/TIHYC8
yH4ckf9i8bn0pTtwGcYMv3AGSpXKcu/oGicIX6WzGY1Wo44NChtFwjKTpeDSN6Ei
oxwO48dan7iy4yBf9UnuqAh/PV/8M1DhEV+VTl88QtRghrhveaDkbWX7nXY6cq1x
G0X6T8e1IiIMNS5NmxWYwT7pPdzFvPXnxrHCIMXGMBdZ0+qICAXbOAx3Ipi1ihZF
H2+O1Z8+a2BjCk9BK8D5G8natiQDKm2BdKFOHkVQCftsqUULrEBiSaXBMMDSg9cI
2Khns5Z2TybBH/kcjm5LnpOP7xIraDIf9xoRbNCU2rUSv3tXlszZ1Uu8OF0JNj5h
uShpzVZDhpeSURmgoJhpGvgop1yST7i9PPwBMCa018ZPrOeR33AIKNnilmjQXptJ
F35aprcltFiQ674Ee3UNH6eBL7HBwYREtm+cH2Zr7z2J6e2jwQ8jOD+U1lTIjded
dIk55fgNq16mIXJb5MQIwFJUTvaJiPxpmLqauODgEgTDKmmEHMcja1/CJxOPUz96
QoUYOut6lZ3obo9EF1FrU/+pU8VEAFnYy5lJwvonZayT0aNupPW1Nr2ad3Sa1EXg
K8ce8N83/y2x71+v//gEInSJBV7SJ4N+llUCNqjG7X8aJUHZVt4hv1Z6cXJrZ9hE
HxjH8084zvrPC72DDSWPXuS/VDDJ6LIBe8X1BFVIwMEABBcArVAzNUyLOWNai0vA
5n0tQsJ0scFg6g5/AoiKlyNX1Z23ZiEe8NoJ0nCzZpDBbDX+pALmcuzKJKPz6LnU
9/ckbU7IAZgkIqGMggcBq3SxCF/yXbUbfdoHEnbUFXHUnYTZAsuJbptiX+DXlVLk
sq+A77WDa1PCsXfsQEqHDdOtqUuT0BeJ07FoUYWv147MpJoL/aHQbWx2dmT83Fqb
rDpwm4Bdxz8q55tA6RcqL+0+ezsdbkLsOp6WCi3asTP1pVRvlr1Fmx2Cv/KHjGm3
Qe0bOjG6my+q8Tp6y736kf81+tZrR5SmLWCDz6jalMrunhyXAxsOQZvnAwjVzdGE
qIj1xQ7QgOb+lc/Q2aB3Rlfkzh36UW4FN+5gs+xhCs269bStc2bTHDH0rpU91Pyj
2HFr6UkTt/at4GxkYU05bSxM32o8xBa0QU/BM5Sz25gUfabR7Us820AQB1N6FiRm
5xvjruXhqx53oDUt93IxRJrkCZ/N4uufse6CLWDqk7HXfJtYV6Hy7UqxBynMJVYh
M9CYYRmM4BjGovgZ48KCSyN1bCgDrdl3POKLGhMTcKmoXaxwGMz+xYtRdWOOHR85
DEClRotWfaY8DMqkrbmSzzd4xbR7+4P9IRkCx50U3MO+YlsCljUHdB3ZpD1gfmMy
dyYEYh/fKeqD6V82Yp0jUuD//tz3/Duo456xVOYJy5Ok7uOuCdezSG0Bwx5806mB
zgHx7ZAK7TOef5EjppnHhfJWC0HZL1AQHwT2uFHLYrK67QzfUXBZf4Ufcyc/tz4B
p8mhnCcEkPTVZj1s8wz7Cbn57gsjWvvIozirPtLtXamIICyKZxbZuDFFXZ6vlJPy
sHIY0bJNmqtKKQsrezu2wJ4JFmvYGrdq0hCVrc9iTpW20cx9SqhcxIUzQ41mbtS3
lwew+Bbi6RIQJ+4uZMsTXTvg6j5Uj/Spupcb/7qFBoVBuwKVEoDNs4jCvATIHP9/
8OmB1p1gXD67aKh+cZlfFNncag3h9stezpfn932h3M4NnAtaqdt5s9/iv8PLbylX
fePhZSGscBLU12fUhZ7wCCIWext3AJJOoI08jtPbGckrfJrlKzzuzY1M6BFPizno
0Bm7ueLYVgu+aI35zKWZaCJ43I7txVNRf8/VmyuNU7hP5pxrJI+B8rvadajlf8Zn
kUGfq0bZV2FEbcxhZiRr52bspgtijRo2hhjffJKq3+Iuvm36qoaQsitb9R2YaRWg
YFNndnMURqqpuGx+bTPLcuZxckja4juVoVpat+2N1YEUnpAK2IWcmpZv0UBwMIXT
0+8ldC0BafCZf/ahbx2t9MLGUPqU6PRDTSl/OSv9SGW8Kj0ytQwHahXM/zKFoBfN
vAjWa7HJy2HtqlSsvZNUa3otlkLq4MsEzwatceIe7bLDSu4JbLNkl/mVjbiXGERF
zEfOQPWfgobfW1iN7YBCxc3AEpthgqEYaQx+dp6qPj0zy3YDyUuK9f4QLsFE3gfl
pXtmSn14gnBC0Qa8N+cYGCtV29lB8jvszhjtn0OAOhQubIrDP5UIwZk9MobNB2WB
FECiGOd6g9yFhNST1J7ldCST7NtowFxgDXLdCLdDnU7YDN5oHkhwgfn0s708evfp
S7mYtLp+0JI+nvR9QmfkJAbKOB+QU/wb6KFG6K3PxxL2RUQvR3rxF4pWcVzrLw+L
K0Kzj+WbqgaMr1hI7P5UyCDpVG5EDmjCActs/BHnitIxPI0b0kMODAvdIeAjziF9
PfzMMo1h8+CfSvUDStOEWnToqFqEl3UtcGU0tiYXPxiSYQZAbOceSS4jcpseDrOI
XmbsZPPtv8ZyYFaIxR+iAKPkOUZtwA/CRyJuCZjVDgN7AP6Ahg36I6zFL4BWZ3Ga
NFZRbGhjML4oLcqDjIWwPVsBvOmgkcNf5N/PUv+ZNvBveWeQiFZaJpW9qqy2k/zX
adtrQmEv+yNQ/KbGeWER6qct8g+8uoLl6VGc4Syku5lCCd4f00KhwTr2GRFSF0FA
TzMsNOmctC6f/ljLBmGu2aPECNn5VXpwL0mFpAr87lfg9UCXeAMGC3aacLZFdmWv
I0koKIXfw2Z1ZbNV5F26Hbd5Z8nC2Efr5EWuxuxwxjED5Z6HEGC1sOcds1U6XKYh
tZ8FeHCXm4uu7A6Nk+JRmpc/2YgVlvmtFPTldaUQpJQ/ac38jRMtLDiJJznlaX+d
qsglg9oWvQ/ZaVVf8K+cUYgvvIpWPUByy9DaOjvfMEthCpaIBrQsSWMPX2h22yIq
uPHmm9wdRXuc15d+DQ5U84M18Wcpr4sHB3rLV2zWSUkI9yFnnM7QmVetbGWezaHR
dMS63k3xc3IOcrZguHIYM2zuXurkys466k7Uh6N7RhlEQLylDnk78sWRars7j9EM
49bE4Pd4DmS3yhpAjYIuZOn+SdFpiSudH7uC65e2uzQa2rRqsm9xlI7MvkCdtVwL
20E+ElL5so7s4GMIPowsHrBmIpoJ5zWIW26MzTowqyRs9i0O2io4Z0zn0JWc/CDQ
Rq3cGZThM+zBujueEtLr+FNoOUFC+QtgimRIfDiVT3f9DS9u9FADJJFMRJnUoAn5
yrK76bGUxP8lhXhvCNwfbL8qQdY/ni2sjRzlBgheP44FagTlab283/2W8VFnWaHk
2epyzaJteEMzcFcwCXddqFSOcIQEgf+JX+2VrC4KqUKDr5Iyditxg5sRAX5Z1DAt
r6YmXINKBWrOMGSClp44ovWjEbZm/cQw/ZntXo1UvbzEp0zU/H7sFNk5CX/nlF+F
n0zY2HfjRqGpGYk5555MufpiLB04ybhr3Ufi3XEL8xeXEtbZQCIpHjgrT+XyOy1k
s/1kHho2I8A1AVz3ltHJnd7jNZURH9BNglCmI0/MarIiyP53Iwt2MINbe6ZX1kTx
sL3ftErJiuaEGfhrZczbswDSHZs7FU2ss+fyg5mMs3n/atbThdLIJCkojpaJVnna
nJz+Fv8UeYZNml66Z2sQCRIY5c5jyXdlwXYjhsrZPun5UCb59aT+FjWrrdaKeQOY
OZ1cL0RSUsSd5s48H91c4Us/M2/S9ESScC3fNRdiDVB66Ao8jo6tRV8hGDbJQvxR
v9DQvjG+djMHS6iYGEF2ZIc/wMdZcm5HWvrRkpE89/4P0UbLc9ytIFgFX2vJvdXW
Um6sHa+z+Cga2rirRmUxOrPI/h/xYFfqWqrAgurX/wsQrfpSx7yXAwJ8fxxkEih7
PC9h34hbkPfcBi9Ye3MuHdiI/2ob1ne7Fq6rahACApx37q090T/+KTYkzIrzsuj9
V+W+k73Q9ZkiqoUmyIFdzBQcQP2qT9kTO8g40H7yyhxrPdNJ69/f9PchngFNCfPv
oLAxl2wd8YwZ+BLf3l2vu8f7WIZe8ZSOHKY+ylh5xAjydqVHEvLOqNj0sx3gt5FM
/eHrpVinUNERJaOzQ4SIRiYtVxYdMskaUV2vIRWJjO7gIkoCRpGZITIb0t/dGnkR
PkPhur87jp9hkDY68QFzmEvDW9UAR06lnWOXWye/i2WYnAMhf2ieNk1O8hJuJYSa
F6HaDxr1fg4d360QY2ZQQyVsxpB7t2+iW05AaEvtTbXir/1SmqNaCkmnhux81fCz
9wqyRAmAkPHr77ol7Ejc/mDk23j7wactpdQnoxuHSyL1AwhgZt1twE32iDUN+3Kl
/H5AeFVEkwgRAljeU93tmh8B375AsB1Ddod9ZB+vCHtUGeI8jF7b+KW8qo2Viwb0
Q5rLMtp4PKLRw5Is7JGjeCvp3fem9ZM7x2QffsrxGeFDgONyLmMNQVvo593WbW7I
+8A6gJfNK/fILgja3iVrg5CFJwjBrwjXoJkCH9Tjar7TZ+mW7nCsVseVjBClm+yb
Smq4J2gNkJHmOxnEYfmkBCW5Bp4jAWGlxFnXu6CEqYEFMagfaeCrc/i4ag5IpbDW
A2i9BZ/R0uNfx9wicwD4hPc5Ut54B1m6F8CMGfB6He3E/EJKyFFsukQ/fj9W+wSo
iGZX43Pt1H9/baJ5QVNo4xI1Mq1yU/oR4sIUoJL9ewlBbegmrivceL6745yHlpV7
hmo8X8ygWmYQdtjw8yjYrNtPEMl/BvIXTv34mH9+9rN1QgX4i8YlKJsFSiu3xHXi
Vb4RjOyn5NxUUada0RyffKhdU0wImi8W/JfN1b++60bLt7M9IsJHLp+2x/BMrxiO
QNL8U4sijjdjn7l3JdF2xls+KpO6EZvr4PObJtH7NRlxO3F6KlE3oYlL2j72GSJ9
RyHT0WLUZeXbvAXHTHPxgUn0glPd2V9bsHY+kgSzOva1uXmlBiokcbuuZ6aMXSaV
xnp9NJeTQg5FgMxfrKq98hZTScEgdqgengF+X5H6G4caw9NAhXTMSwKz2X3UTS43
kdgHztOCwcgLiX3vHa5zx7qOmuAAZasR27IiE3HCIHWC8BniG6N+nkfFP1ZqbWIc
IGZEyG4dx8rmJHBl+5rlEL47bN/5st2v5ZKZPo609z7uhADkL6WFDfiJtiROyryg
1+mHcblljfZgP2lV2EM02WIC6Hj9Wa+8PszHG0vBzaUc12kE6s8s9NXgpywN/mRs
j/PZ+NVmHpBNik1BU+YJLxo9dXxjTdoTMMHsEhQZg5YIERs953rId81vaaPZjYeY
p8j0riXJbXOO41DxO10YwSMagARgYAp14DUXhr+8YEHqNC1e3mu9InWvCq+IyWbp
XXZ9rwSUnk3ZDpPq6XQx8dt/FBPGU+AnmDIQmlJu8nfofG9wOoGhOMolVMu6Lgrx
gZQxhKwoILi0sixA/F7E4GDHBbmOLeHfSm9QTrKWmILvaRaM7J23cAym/8wSNi5q
DeEqCMqvjsuOG5uUHs5cSSOh3KtVnyqmvoyBgT9GiC+6f7nATJMD4wU+GC2fQd4u
2G1mfUKuzsEyK0KFMZODt5ipB9NVLPgF0Z3I4ATMkx30B+edVFn1Qz3z0Mh2GhvI
lCpW/lPLvkMIwTwBV1PhbzI0TmJYxq+bJRFRbZXL41/6cymr3L82nbzOQfkz3iGX
zvkiT0DBQkwYFMwvxgmetLOkHb9MSajxUwmz649FCyE9/yWXnbWjqGZs1CUXYdsD
eircQ7C4TTcf1+wSOvBdjWW5az63fXy5OG7mZp5mUE0/TVhQatNS2c3HeTy2FpC+
SbhirsWgh+NCsCNFuTzhwstlxUyXqIAM6dxS2WBWNDkNer4KGLIjLEPb2Q5TNLTe
1oISzru2DASdNv+VVjKbtAlBcJJYHrQVxEHrBpS3Aa7QpKDGR5bwdChSDbKVk8e8
xa5f8QIME2PRmRVw2bGzBbtFBphKJfSDh5QLr4fkWhgzqoId7dYIWNNRk4eJsINt
+BeqK3sJcSVkKtMLDzuGV+PUQmhe1EoEkepCcFQKGWePxMgAZv8IoGKCQZyYnV4C
YAZcq3pZpQNlApCK68UEBwpsmOmOxPAvzA+K5H764pWEDgN04qR9Msdomc3OVKM6
HnomhvI5x1XiE8HlcECN2qIE6nO4qlsrV+detLz+6GH4nF6x+C2It/59rz0UJvvR
0ECWF8XQgpQHmps312PI+mf0Zi6DIfdQ4DwWA5/xaLmlWm2g/zkoBz5cjwgTNN9S
XeCtsOCuhy/PZxZmWhcUqh56BcGi1ViXwRiwguV7pDXsr500Xj9E13VihNj8in+O
ruiH93hDkeQTSZIEigvsMM48dlrHEL8ASsQE2S8WlEmlHJCdZFpyvYLt5yw0tFYH
hwqnlJs1QyjDa4vIMm+yha35LzSic8Nut6udVERb3Z6KbEqIWxDOpEo8QNZWwtb8
rtg96hCYDjuAhk0ytgHHHJWfOXxvc8hKHsPQAp0nCDMAMbCBWFaCljKGkuj++kX2
ob3Rnat5eI1YkM74vYxnf94puSGfP5C3tQIzjra7q+ORQRURQP6G7RqlJuaeP/3Y
DFtvXnX7PVc8PDz/eKQZT2WYSCTDX1Z2qC+wJF8+AIl0zMGZ5kftoBmnzSdJBvDR
XV/Irk7ha9ht8iPoD7ZPUACdsiN658N+kTsw/yURUZyrVgOPkxMBsy8p/oLixzUl
Mf6DzCKRG6/6j5hWADxdW1m/7210Gxt8/30nNNmIfJDMXhIQNvhFC0528knzrhiC
Jvqzi8mJhJ624YTjF+R+G2waf6o7gmcPa/hZgKup/kkOBNIyT/AukeE/rZIr7anr
H2vPyNMvzhjhjvr0KLZNOFTtlD2aJR9K5ScoK720Wp+1eG1mXwTrvcG2V6wyatAq
cqBUNDj0cU3JjD49voQ5/lO59ZXccWaXsMKmreGwC4qMpFfeS6eeKDFgtBHP8i8W
yUmjtDWr6zktYpsA3EGH0rSBcfQDZuy66183r0tGNiD61fEMLFpR5meXVlXKI8eZ
e6vrAxKFeSSwtNsNh8wga6Furyuf6uBGcohyN7zLUr6gNOuWJjRAHsAj6uHUFxIP
+nu1JX90bVMvyanIdbJ+bTm9rH12NMayNY5PMtfq5RdkDSEw3O1tA6J56/mXUUgN
CVl57Kwf+5o7w24oPgByMLeGSM1WznG6+ktt14AeVWDsu5ocSyTzrDiJLCayCk4f
4hZHrzH+YYE8CXCUsEowKexZ8x/i235heBFdViERqVLmgvjosnfSqnNfKbp2D+8y
SDQ5YZOpzWJ4VAjLiMLfdxk8gBvJV0cEuGV8TDBCVt1xuD25obqywtpcFyZgE+kz
avdA5rZWnX/xXvpDnAt0KqtoZuRJiOex748ZqAEF8dslB5Aikaul3eyyNYzn2Kvk
Yh+TDC3ltCxwbZklAzExVQgIMpPcbLszagLOye+xieg4fbGfVmCj+ycRxTlAR2zt
FryH/KxQhTECAzQkQeDdsqDUtZCJJp4S+ZnUvjy+l7o4deylFXboFUM5YnobxR5z
dD+l3oi5SA/gHvJyxI42Kpq4ez06VYPIhOGIkuvjTbX4qsMzPORSMO6HQCcO5W8J
3UWsapnP2sshhvJI7/LwVFHGMgZTM2/RoGONyod0cW0NOGCR5qmfOHFo4F+894UX
nC+RmA8OY1p9dkeD7330AxJ+XWJNhIL9mXZyGcjmcavh5oKNLKxD3SWxUUJaaxvh
+BC6ae43ggwZnnuC3x1Q6r10i1VLKm6LXSx7U1Oh0Zwb+cf8FwyqK94wIUmudcXA
n3ba5ZdpVrhMyVibS7ejh2XmVOAgoUVp042M+jkXA6yRIX3ouASwkt1J4CGG4vqV
eHX7DAaAuAx8906kKpdUmClSmTbwoVOM+ubiLb2B22JonzNVt3p04wsJ9bDJnYib
Cti4dsKoEWnBBE6YT4/eh2ynWIHTchErH/Vk6SX+aMv5JW+KYLywQ/EoaZ0PpqxW
NSXHyDwSQF7Aluv4IarhgesbtsBNxJ9p1s2ndAbmBeW8ZuKaYLB07THujjQ77sk1
qHM6wmfTaIWnmYqE0peYtzIqDkfBtPbOU/I5of/XwcaI0afFCotPZfpiNwT9zbil
x8JY50mOxB1xv+ed7ocuQf3iSw6Wb/bG8etJgS40AOqhJSVuATBXEfqvpsJu6Haq
GVb1DvVedlfzakHW97kT75D7RF8Tbi9cEG3oW4G3uR51V5laUsG2v0FIGr4wRnni
98kTfX6NllJv6rHYUtKyfI8Gm4Aj9c3OwolDSvmNkfNEshfN8RkLHI+oEPwbTx+V
5zdpaxwIzkpOhCIfTUt2zVfT/F9DolliLJmUpjZg4Wl1qUGInWpjGPTUxaxA4qBV
2GSioobVR3sd4HgF3dcyzr+1DHF24aCqlZd2m35kYKx0Bt/UsGytDQEu30EFIK81
srt10qa5G3xbvSzzT+xYMlv/tBDyqOrcfnJPrBDY8NXeHE4sio93t23J6hTaScBf
PJF78rLsnsUKzeJKzo4ZuOOE8/3q35oAfHpDGFLhmUWVSDWnJzgGFqBwoNvMhEKZ
oMCAMXF71yakUDV2E1dwSvpx+gDSGxhFvKjhJ7Ah7VQxDR0JAhq9415UeHQu0WPO
bgieCppXdDzGJLdYlV9zD6jsfsc0ZWUthFg3GCTawAdQc9dGJs9X7LKQeN1jdQOp
b/1kUfEwGpLstjiAKDtKWYwf2zn4kCvINNmIl6aPf5O3Yc1cONxAjHQ1KWgOP9mR
rSfzMNQrTZC9gLJLOWCA7HzjaKvUiJwweCAkFWTbL4nNYfo/hLYzHM25knPmhh16
z96GdeL6hUEJG7s/qcIDI0/unrr0O80eShkUB66TkYR1+NJW76n6wYqULbPSaEO3
T+GsGb+egB0Z0aJLAwYhgkf4PpHw7puGXm5m5gw55thsHLLHM9i2+OwqIMZ2TID5
/vQE0+LpTJ0+K0MNCE6DkN1NRhiIjKGkE4tZWCxShH3k10NRoIkYoDfQKZUAd7zV
TzNUOU4vj2DwxERIhKJYF2HC+QRoSt4JTjXxUl8ODAJDtrq5SP4/6/iUke+Rf3WJ
LlrfWYhuXJvNI3xL5F2c1hm1tInEu8+m8SEp5KOzQNjHTuofdX3vcHYeC+1Pma2K
hboX4RmUmFBXrZnq7x1GwPviqR3e6rUkPNSnrbtEZzU9d44lc9lWFdWAlPRJsX22
CoF5JRBQKTT+BAcWM1VnpeRWf7xXvXEqG0r8Ac5Dpg0zfg3sXW5jT4WcIT5OL6p2
94JuoJpF3Y8uVIIRmQ8hxLp3htkBai1Td+tLuOxKw61YfQ7VUzs25VaPRIhpzj4m
/g8WCcshql2uwCxpv0904zi1hvDeyqOvKbCsT9IpSH3cCFPG7B8tQu61FpaBHmPy
iR/Ieab8NNvUkCbSzS+F8ecbQNWOMSvVSZF+LE9afclbwLyjbWYAoRdHOjsLdRme
lAi3GJO4Om5hFLOUvWOg2vnYqcETgpgLbA/NLEdda6T0+WsxzR2aB1yQzU3Xy2E9
8tJWQ7K+JCqzzjkW5mKxM+617zfVI4/DrlVGGw2QWILY61PiakVZdSTmSxCM5zwj
aYkh8YOInZvpIZ/ilpMKhux4y+02DxCvlFI9z8qPq+6d5MgDRberOnopZwl2t30M
oQ4IvFzkOCf/A8l0YBstMaOs7hWVIL+VlSHvrH+5nGYy9n2uhF+9YdR6ty8TQLcK
uJyLuhSC2cW2BU5FCgo26lf3GueLUaDjHbJzXe8l9ucWMufqPMSeTZ+imiiyJYMv
8jowBDhkV/ebf/PZ7z8g4eYbDvLfet43dayx0uhMTkxk4EhyPHuo9n0O0ss8hmdQ
45vAyLJ/pFJ9CNtx23Zc/yoPzEFrjZZmhrWOCG2Wm2e1hSiirhcEcYJEPPUEVleo
cpZ1InWyK+WMGWxeMTvvr3GrPUC9qYp81FDx6xDn7/3v+VxCrBMWU2V3O8bxNwVG
zwwQ4sy7g1TTPMokEDC5XnuMrLV6Hhw70a3xa9TOm0TCuKyM7DGY+voHlKKhBIZS
yk+OI8iLrvJtdDAeVV5Yhe9Ozrznc4jFowBkXwclHqvchM+qsHxL5xoT31iMA02p
+ANVd2G8ztmilYz8Tcx6Uud3pX11y9JtVUY7fN1a4JJZT4gbJIamFKEjVsG0vlzL
ydndUQ+bi94plN7YPOxYGrh0+3ll/BzyE8INKZ6cVynp/qXLDJ2iNwxbPafizqEc
c5BcdoibFfNeUhfzgKb+F+1Ii7PQ652oqhEzV0UckbOYtWYeb98TPh2502KlmBqU
Nk+DdKle5a8NJTRrxDqk2M9hET0bunWDpRzOh/OYtfZJUSuwX1DgG1eQJevUFoxN
phh3BBQbgVONA4zM+O9mlePKb7+5SYaa/EoGfT1ndWOpgadgk0/wedu1rRoelFkw
fxNWHw+O9MoY7YUuVu3aQSuhlvDxYZxgZojSm/IRQfSjUj3OdfKdsFssRIP3TPkI
MV2o34R5iZk6YiHEQRZ0wrC9vQ/u4YDTVeKugxyfT5bYpVSeP/EEW74+278fo/M+
nJR8aFKflrRUEshDwsxQ/cOqEtYSm+O7EkelmT2skW6wfzEwsje6QO6z3xPlCwe/
wX2MnvzwkakfNsCH2VfztHi6X/ix5I8lOaXLN8DNPMTczk6CFef0DLAOjXCMn1zX
1LAY1thQuc0QF/tOQXJxAg0whffYIgiYUe62ajKsgcwvCM4uw0tsAs4zdgbIKBSM
1lEJ1ZwSTLeR1hij+st/gl2RJ4nz7pR9+6Vr9mn7ukdHXDgnBXufZEGO0CxClV8k
p/gogkFap/dygS1ObpsLSGC7rSHrib6/c5N7lTDd5rwro7i/obOaCd5gkZvMGe26
PHoSSzi60OvbZghcoev9pHnEYobS1ZlWjoCU6nvdbVVOEGmQKPoJSiyqqY5fnq0V
jTruHeaF9f0zL2o+8S7n37Wod1K/L9byemB9TCxQOFnPYq5WnSFRFohJOTqOSqHE
tgnE8RVhmQ14CijxopvYDIK9sv6xZjX/ir1ie0ES3OF8UrERyDz+Lyyzx2DzvutW
gWVCSMYtmQzwOhMIEeJvtMgKp+DpRlgPTUpIhj+RBaAnb8+dvaLPD17ZkyfozrDN
J34itXVTcMCrruBWUEdNRnlOKDU8ySnXRn9TCOg8g5eA9Saw5HUqc+ZePmUg4ZJO
CIKYGx/PduI90fl3j7Shcc3pLa8ivhjocAVBpTiNleoX8jzP+TbQ8z4Kh51hzM1L
TvDLiqw7iBWR6kCOUOhyctUNOdOUkGpRE4RRuHPGkp4bXrvT/VcEi5Q5AykdgJOG
o+e0p+w7Jncu6AVdi7JV4zHdCzobIwNtWt1VwunJ08NfR5JHt1do9In2EXleeXJ0
g2XoyUcwh+ioQc/JCJ2UeKv9XbMZHwMrKVgL1csJcviat/0H2unXnTeC8wiQT8Cw
fP8n/9T+ChiWE5sKjE0oMzPhaQTkjjoExBbG6aUTKELpOubJAwctmNU6NN4VcP5s
l9MPNeEnosZrCbM1w4ZdtTKxBNk10hohsPsJONSnYaTi2I/t2ObSf1hO9IXBPG5j
Ry5FH0DiZdAh4Yl5JJFj/LMTB+5Az/y/kaY189mkMxR9TvO8JBVOn56ejLwVfrOD
xFFt7OFyUNH8XGmnk019CUkTVAZP/iSi3pEsP4urOSGCX+SGxvMo82fftxRJxIgP
+h3J2xKzgzmIYp4Nor4wWze0aOTACPhBNoygVA/3u8DOifXIKY1LScfK0xQjsUPe
Ui4CObYih203j6GZakjAA6ySMOczIuuB6Quo86j+mHY47f765cA2AtC9QKMAgXOp
NoocKQhjA94Zc2YSc2Gfh/QK4ElZAChh1iALyeBZu00tyunSSBTrg2/pfWJy+m7d
PcIESyGpxJEkgnGn5zaXp3+2L5POX3hsESYktNXWZ8XF6KesuPwG7R9ewrGIGRxD
UJGtTuPGdVFXurP09GPng5opoWCMKaq1y0IgF6pmBnFvSrag0SAFOKVg6txsfHY1
fhUW8KwPcr6efiXjtRgqZll+aPF2Ec998u5bnPNDMpHV8041G7aICN0a0r3pu5C5
GXSLIYanSWDmvbUt/C1tDz6TlY+e0l3nyDJuCSiKb0+/omQmhz//6DgASlrC2cxp
o/GYzlJd80ni/v5DJ3g9/oqTTAXn4zD2vGSWDFkpuozAE34BxgKF90aJiz8F7uZs
v5THriQjo6z7m3E4otNwfW14XSNXy6oSQnhlKJYc9XJ22Mg+jVgFRqdOcH9GTxSx
5TyYDKNQiGat8BlOMorZxTw1MZY9EgvxJDi5hLrN8Qa2qgj8A4w9bTQeMQh9Haj7
BKFcS7F/EvBzy+rk309vHbFMLTZmnn5siSY9dVns5NahGWxfalGxAEeyo7eJQW1j
ipQpVkNvZEOkX40PIr8UFktzi72mR3+dXZcuNldBywXcsXWuF5BRhW9XovCWTjHR
XYiBj2Mz4BNDUVTXev2sh4u6RiXAevmXViTvsqkQ0fc3lP2b4DYN72f08rxA5WC/
vOkp2wHSbGveotEMg4NqKkfzQiv5ppMVq+Hak/L8tUvLSh/1GHkXLMDyzvgygQSn
FqbFCrC6z/y80euHZhC0sXIIcPRCd3Jt6VQbnqO6wxLSyXQCl1ykS9tCdxraSrfU
TAFG3SvCiSieyiS7vbuTPZJyjlEbqYmmb+/e/bKopjMvhKv47UepdQYywEWeuGT/
WAkqem5ArX2qpU6lpKSuBXFAVTcprSkvDaMtEGUSqg62yRR1mMXi7nFGhPu2HBrF
GUloZiVwYgVse4CUhk2TzB3hgFLlU43Y6fyn85QcfY1hf6Y99MCJb02cwwYAwxag
Lu7IWYD7WPNJ+wNzJe5ELNo9rP9Uzn8gTpguoTE1569uUeT0oToC5N2MEbtN+tRy
YdEYBA56BSnloetZjNMtlHBxDu4UtFYqazwKYHKOOibg8L23wdoojxVM8Hwyfj0f
D5qexRFErd3qjWBzVLDIG7ijBvKxNVofcmmeDljiMDJNUOaxoJoyQT6pFUxj5Oh7
Js6Zguf/5gm03HOac+6Ph8NB9q1xC0JTtC2XkwQMGXQ6x9sRmauXXFBhX9VYPRQP
Gfo4eBHhyG3U/nzhlfgkNt/f4iYRMKj9GawrxbSRVdIttLWZvvwjnVKPeP4l1hUn
FkVgSO2iueHjHO7/iDX+cKpD2D6OU+stIKFgPz0T2N6EoNn1OYkhLFT0642Z/4Vy
DmCDqYsnph6XT6n/4PbX8vid+xJMDwRjch6JGcJobN6PGdf7zoKnwe8kwvoT35j3
EiXb1ZVqbGjq2qp3pF3f1NnEZSDnmn9gWbjbqzsm3V4sNTbJPJvk3vwJHQ8z9EX4
3bfOVVvpj2JDZLpDsseFYt20A0x/CD6E5mms/4xKYtDlDMQCHxmY876SGGGBg0uf
9RCRPPyt0sNzc8PtOlVEqrJzg598nq4zwVjrC67Q1R1gbb69xv/HEF2fWqKzzBJS
Sk54MQCQglFrGUGi6nRGatFuosudQ1Ovi0mXXWifBA/lzwV3V52dZQRvoXsER66p
REDAfMaLYmI4boTgWE9fdePfgMlOq3t/mMzy4C/9iEQ/VudhT4WnX7MzKsAeQ2Xb
FOZFAwdH+eEteBlL64ch/TBIbBoFhq8iJb+ydAFBCdNrok3rboih2DCAMwTr8xMi
R61C8GKRShEsnTqxjxvCiPzqaBp11BW1G1/U26p/IHfmfiDMi7Z0pnQeJUWTG2WE
K8Eq/zKxwn1AdoxzsdgFepCjdBH7tHp9VeqK7Y0HTMRj18xU4YfEvjTBZJN6nGS1
iPu/weX9SwX/qWrSrk1eoqklg5JetTmBQCmYgWhOEYfKixtFjKOAd+zjtIHfCjX3
o2IZLp0M30NLcdXTWQ2atojow3hVVyvmQUXZGibMy0/6rfM/GXvzY/QK5gXvLbyQ
rjJXlg0T9nM58q5RUzQQ/DhFhAXrioQFoc1gt/9ndGAVPjpyYSrmH1yGcqd5ovFB
e9UMfZP5OquzvbhJxE3DWelFq/Di9hT6UKKYzSXRVg6fp+UUVSPtwjen4AI3LEFp
6r9u5YwMBlmXN6lzChGFj2bSuPCxa1LMDv14QZYu2Y8iVMKqydSfgbiukDeeMq7x
U7UwRPJf4uMG1cm1ZyepwqrUEXsal1h5skJiTTR5nQW4YuYy2/kkY6GEsvHjv4/L
ZDnmaUw/CUDw+10afN8LjiWeG23bA2+bYqa7ej/wtLtlFGON7F2cpBrxPwHwoKnl
4K4tlmx7iT4PSKq0EV4Ve/9W38ucvFav/rTu3gtVj4jYFPX8j0S7NGJYjjVPJI0A
FpCeSDqFY04nY396x29oY9YpRB0K2n7HZeOKRuB3CTGJRtS7xrlJyiES80hZle7K
sglO1uKvbx3APfBjgRXS9BEEZHqe0UOk/hbd2pWd4v8W9ZQcbkDrpKRpCXuJpwCs
GnMhzBcDIiKlAYD6FaX5Gkr5qTPwmhaTEfoSJTtPIoH7dsJwxRGEkWX3p3zrQyIB
6mw63Oxrkn2MHTDAmCtanSf7krfmmneTT9XSBPByXJatGBv96fFYqdX2HQdW3RzM
az3Yz5MJaBg3fNy1g8j4T+HjIjkQ2gwMZKivTpWxFRK4wmXmdevIOWgAoZM7mG+S
FENlJfA5foHP7zAZGJxLAhs7lTOE7JkuZMJXFpiP9Xg+pQeytHH65LMsbrVoDgEQ
taxfOnV0ZZUJjCHqsWMrOhqVGSGzdLv2LPYGp/wNuwOn70BnkZKTq4gHORIEoBwn
hjG7DAfZCM1EidAKw7+mKcKE3vHH6ZRNrk+Ovqwcv/6KfyHK8/FoHxl+JQ3GkH95
KRVc1WSfyEIOKz1J19ZZ9AqO5sgAnfx/e7S22z1IUM4KgSNhoBO0aOolVHE46W1I
hcyLbf7bra4X4se5biH/vLXYREL1STSVi604ANbsTYlVlNL5OPjktB3v7dVEdN3x
Isfs34x07R+p66IGeX9lmikDJfslTOWnVrek5ilFtW1Qe0RQbZDvWAJ3dMAhCzol
eUTYrmR+87QXieznSjS8rC8imgxHYMVAKa9VHB1OUvBF6zANilkeJHepO7svrdYJ
J172j/nuG9HN4Kqy9apAeIOCuTwz1ws5g2pbwHCXXlhPdnPyD6+auOujl+KogbOh
+TOVyqi0xjBp5XC5WwAx7Pj9Q8RSejvVb0cibOWg6mX8glFgqjSLlQAnBLd2BCLI
vs00Ozqk8j0pEO4SQUzOEp/kG74A3rsSxkD0PdRvgD65NpXF+EZweN16XcvoW4iH
w3XltNgvtoaYNYWW3A7Z2kAAw+reUvgi1XAUEPfS90nReyYcSniuRKAAjkZ26C+U
sFXmZoUpA2SwEcdyS+3BZGbrGS874A/ef4mdr3G6e+xtzw3bhMnbjAoPY76+UqEf
xFAJTI6CPW9Rq/8GuX3U0wp95nx9NMcJH5k+Gt51HRwwnWwo76BTRvfyDWIjjj8x
ouQQfF1gQRzV5udiuChsICGnI0I4vkzunajKUgad5+kgCMSMcxUN3sF6vc8X7AeB
6HjU4h81SGJTmRY3olcPgqGqxU8FWSUL0qS4zwlnqIeuC/bCwEJ3POeFBMU3GDa4
ZuFtUHEdcz+nBUB+JzqhcR08SQkaguQUhmW/w1edFO/D/rFUF+FzIfIRmBjxZgHW
LeSlnrYAntZxBGZRyX49X5wH3G1fK7vfu+OC2wR3nRKtC7uieMdsoZoovzBBaw6R
3apV+ws2rzrwwk8bt+qPwCY03bPcw9nacyZxLarog3LOCfK2Wv4VGwK2EGm+MKJa
d5mWX27r+mEkesMjHt4DW8ofyV3IE9aYwx/MyWNFGL4bHkNI5P3TXS5hk+eJ4Uqs
QCZFbs0C8CP1mQHSc5pdPrUBVlinV6lHVXzRPpkLCWq3zLaX/+RWxC4WQOMfhf0n
tvCtzq4C3vKQ/LNXYOoPP28kFv9rOvKwfZVV19gCq+bEruWL3aOyw5Q7wuPD+Pkj
fVBWE1SesZHPlzhNpvLkj7IKXCtWU/O/Nas9czyxmrcDSFmkeb55UI9dOKLlJAbp
jh1Gz6zqmUJahB8zjMwkan5Fl0tdzkD235xyod5HFADh1+j89M7O9tiI7u9JP0B+
kRQnrxyd0pEBVEaUpqPQb7R99F6BKX1BfZotG9GIXlZLnEkKWXsc9ElEJ3ciehZD
jJJA3w+JLDfxsBEWl72OYqnIwMr2hGFf/+as7ldQM8W0Cu9GbYFlDY/PWRKToMfj
/5BUgfm8tc0v14nG5hSHXXZTbW7OJUI7fvK7fBafPkfRYoDJhBCgMbM2jtT6Yl90
ZuND0J0t4JlIXtT3+W47z06c8XTLS6/GLIIpvwNLRaIliOh2xCbDcBjAbokvC+rG
/0vYclJtxaY7YtQPLMtZd/v/7/qAHjCQFiRXklLUOGeAnFqSyiFwVopTj81S0JVo
jbHNg6GcbEUebHbEmaa+cIHmxHrWqS1nvAqoQBGpI10tVdoZyVLQjaZqMUOT6B0G
66J3SzKyU+c5yQlTlvnZeOvLAQktshWn23Zh5Cm0NIRdxdh+KD/FqM0udvD9EL+b
28xG9b1WriBU3qeEqemLhFw6kRk1g8I9UYysHlQPpOb2E0rAcrGj3Cj3UMNvA47X
RZIymIrQvoi84Cin4oI0MT7yPfGNy5iysnfq5VPyY79oR/rPdRWKEV345QYK06wB
W976aX7v7jj4kaO//tzWQDUBir0iCeAUFjZY8SN0iotr2y722IikRyIlg0aSbBKD
tmyCtpCDfFBcOnXqiFBGrU5QAIUh1ALiSFVPvIi+A/vqU1o34a/Xmi6NnG0weXft
Uir3LZGuoYqDJLZqWM6S52D+lPRr++BwfRRXwZn9vlsftYOsNvtkd1ly9U4e8HsU
dcfbayE+B0uF1/HqPmxIiqU0dFW9hmKnDmt6i1WBKOlIlwq/cANAipVzmN8Zea76
DaYiIDsIcrXrYyAjjEYEHagLtEoW1hWXXaI1ShI+uIcp85rfqLt6PLGzs11C3ROI
iCGIqNjx7iaczVhPswDJMKGMX3SISSV7ipJtFLAPpf92akPJpLSGNEFaqoa0vWay
TH3vyxRqgWrz9sUXhgf1UFLFPs9X0Rt/WAnEFPJyUVHbU1zLzULtdh2UDxbzM+Hc
FgpkGWICrA07zCYM8YX0NgoVNBYfsWFV9GlKtvNGOchnCfFGifrjqXxlJSli2RVJ
PRlXKC3xbCBwy1q9iFHortuT2f0HbVnWsCnOssw8X6XQ9GYMZdFtGQDRjVWA6Xnn
iSLBF12bw/29BTk18cDQMyPUajsn995N6XdEJSTKaW8YkCVz/cjc0u4oKYVCjbp0
Lov6j1a0l3Xf9rT9oYeehg6zKzGcF1WO/T09sLoz6et0MY78DgRY0VzTEBZIAsxw
7paAbp2cqsjUiR+yAbXMREgOFS0fhRoiEQmoP6KvZAtiJL4Xa92O+TPa8XaQl3rC
eUofvF+e4PACOVnXTc0VB2B13B9966UMM9DREshuhXOMA1cMvBSzzIHi9p+sIiS/
VmTiz6a3TSOKIDITnwxu++eOU4o/R9h9YeFB/w2jRuz9zvvh9nd6+JpRT25f8Fy2
DfkgJB29WRUH+iELRF2yPZ/yw6pvThNYpUHprJy1bv16f8qwM89MTcRTP5RM0Kz8
X/g/3odpdM133wfULH9L26hFYZdQPHA5ElRh05JmXHR+bbnJnlAiEfG4Seen/K3X
slci4CZw8G3FRKsb0Floh4Wi4efQgS0xzUALg8PAE7OUEU/DLELPwRF5OblsoVs4
ZQxUfYit0O1F9V66L1GpDuqelpjAaXaGx2JgSw311AwEjv41YOa/O82+J3p21oWF
N4wjTCdhQjX3D9Vlt0clQ2Sf85ZklgHF+n+qm8qrtDdcivDZ+KUK4RNsWfChdTMn
fK7TlHOm63YryGNzSWcFR5KymBN2zhBrbIeducT1UkVgByUulaWwrYjIChOwgHqp
L1Zn1wqfdXEYhZkFAs+XlhJ9X93yV4V34bDzdhrXq3iHKOsdmchCVX5FhrCobkzP
/vexUUO5IFJjNYMugn+Cj/xjJqAD7ZW/ZoR6ukPg0ZXGLUfoz2dQtTb0Le2ChpwO
PDVgE2nomZQGoIDioegXMFmD2Y5TIQZTVrtYzeEHbq44G0AVIgbINfdQs8t5zOsv
eqUsdShOvyUl3GvUUFO9wQTXL8UNKT3mB6IdsgYBOz59YItCM6XSGeen+T7H4QWy
U2Ik6AriWBF6LkWwEBUiIiAYmiA8ixwMnqKYUr4PYHY1iQXpHIMtRf/DQ6PqaaDf
B4Xvswwtnd9+duWXAbAs51h/hH12TfExZ+wqDLsuSilJGa+hDMyxedXRJJ5kwruS
9B6lgaYoBz2VYQJpSrtjILHNWstjclE6xUS9seE+TWgjaPGNObH6+xJaFQNs3Fkf
yt6b3gH4Dq+04k1+eg+lAMWVrcM1m0eucH5kAySCK9/KTlDMkx6tvHqCb/ZTJq6N
78oao7rCIST3xF7vQAhkcKH6InhnF5N1S3a1Kmtp+wcRMxiA3AE0VyTgi6cU2WUc
T5p58pSWdByipYRen6DKdw36x175RxhSJM7yI9gJeIU44whUzFY3EEzLvaVEqzww
+E6hZutfvJ5ldoholRwhXzaycnn8ap2pQwfS8IW3bHsFciZiO4Rg4ngLPtlgMJPT
7Fx1AZUNOMUM4YRn47cPdGjNn1haS7EEvKoRWbIKemoWjDJ3DNGdPJ4bOv7Yffr8
H2l6ux4brJDG5bZLydf/SoZCgkB7NfXuHm+zrWaBKCIJlM2NO8k7eMIBPrfnQx5U
YhC5VqKf8grDGnmdARfAq+vbUB7yh3ossBdO3XyK5B8UbxTcTCZlTn3vGy+C4FG8
IjnfMRr/xeUVCUXtjzFM8YTZC12dbtYfFSWmog1lCim6KCZjmXAX4aT8T81pTV6G
GwIJjC+HW5qRYt68z1jK7dUSWFxgWgSLKp00K1Pw+VPUnPT2QCl2vbN+xgI5LEib
c30da88qtfXJ0dTvvOTEhKPgXjliqeMDcSyyhuAvRMZpe+oEY6AJov3tDmatMZFW
hyvdUz1afotPZqt9C1KaNa3kDfGqWXllF09teolbdZ2Z4g7Oni6qgFDJ5k639WkK
6BDCAv4/LwjJ5wv7SK6Y9MLffXmjN5izdUHtfuE/ffD1ZXttdm3XOuOibv31NTKy
NnUPiJJtvYJOQTqVp+dmDTgiRvLallFlsMSMnE83mtIVT/pc9qwtIoQau+Cduf6u
c+BFz3JfGJeZDuKzBWpKw3USdcgwkjwsdM4UP+xp9HkhH8izIKwti24KRxv/jyvz
QziRdJCUTkmdyaHho1t4BSvN5rm5plVT+P1yeoRPBjHEGx744B+dFIg3coud4uZn
vHU9FyVfSJC570LeAmKQbGkcY+tRXZ90jJe7Rb4/J7R+OlnQtsBDBlTR+c7LdBon
XByk87JoOIqQoB0d2y5wV52ugwYfXHTyaLeFpV4lTrjwI6n5ncqdbcVAVldG7kfI
f16ssfv4JX6goP4x/VxydkSsi8jtftD+ZJrlKzVPKDSNBS7RVdS0KllbSC2ca/KB
3axtHLN3pCh6LBMxy6UPmT5zqKK8/sSZLu8Mg0cN6oaXTO3Vkwyqscny8nezHW6x
fHJstJn75oDcUt5JtedkpusOOgdGkXzLfstqUO2dvor5a3i9jEg7mZC9+5h2cRv/
sVt+JZZA2SbrbkVM93hVA8DhoiiIEMw8IQjZsvLzgzQEAT1Nbw18cCLz1inmCMmW
a6caCNyurDyZG8RowiEjrNBAlHrRuSaQnJLQoW1dJdo2hx26GQrM7jwuWLJ+aF75
C47vAkBSKa5z4i8EyhIVzR47lUbekKT8Q+/FYqtn06adwv+tBAQim603HE/BtJx+
T4vqJo4D//WtbV/B9Fva1fkn5Ykn01zm1PVckkVvW2hsthMoUymnTl39Ft09DKr2
tjb4VgKpqiHay6LHnPpA4iJYDIzhoVODknfDj0WIvtoLYItCA3pR4/H2QSauxFDA
vpqPr4e6i5kRX61JIBIZRsrw50pa77LuqByszckto3L16Vc3c7g+MEKwAyG/5E9D
JQXpd53Ign5kajiB8FS1iowUQQC2ZbS80wc5X/Sicc0vz7kLngLqfEUSb6HUXfre
oMw/JIXGK8oYTsuySbZwtiupmpRabm/BzXCBFNhSQA4AnKLIDmcUHeni+Q0JybtB
x0ggKy0dO7H+trcdsQwtNsclwdlY4+0ZQ0H3OLqyFJmPHM9wV4yC2L+x6B36MWlY
mezath5NoI7YY36NfmxMrn3ATJe3kDdnnWsGK9o3Q9qbTamjLkeX4xTbegW4ySMx
L3HzIQ+we+iMv+xm7bibrGdH287AdPy75vH/MnQxAycKhVOwfzdvsFYltDAeBTgr
QdunKmNWjCsthiOTrTsHYJVWHXR87oG82UUTDpm4JLle3jSV3YJM4rUK8CoqOBQH
rHKeUbldUUa0WhA2bHoaWeR+NEJNXEnK1sQhAIoaDn/y4rXxUNdLvwms4z9A7knn
r0lFehpw+RnIEG2ctF9uTXJqB6KOigN29gMfBFuamCrCwK7/+uSMZ9uaY88rha+j
JGVSLfQ2hmVg0O7ctZffQbkMcetLqXdZHNuanm4m30QSFZ3iAxZnwBcQ5PFMUdac
l1MFdD0f/1rxY8WlKhKJ2S7H6T6iegflcPN4JJz7sXartkICWW22Iz8KSwutmGVz
0aGu2/oSBQEimS0akzNY7uqfyszpRFWUH3c7u6nuwmEa4k7RwOHQaNlwr0r44MIE
HfLe9aoxyMJwVkVoOYY8emp+uNZPDKJ7OBiut0bPzkBgmsYs/N9KbtoZ04sY4OYf
6m5yxYUQ0Mu2s4l9klSYxE5bF1Ggpqdd7tQEvDzMKI9wZHEorxli05QKi8MS4n9J
5qnjntYjboTUkHhae56AKl1XGqmGHbBJcd836x24aw6AtUOEaTAT9NYFj1e5eE5p
0kbshdMmNViPgqX2MA7Uia58apweHBdSm6jmfO7v971jMip0dGAxnqeSe2nbIFI5
oKUi0XfglcSjW5RwpZkTr6yXO5RTi5Nkw32JKJphmPyoCTrHCutKwmt6r5adUFWC
ax5PbSPGuAS+LIe5fUG+lEQ9+/IVZY0oWo2KNOa/CMj7EoAQXbCktK6658JIeyN4
Wtr5XjQXOYSmmvegH7Wv/1um6QSNixUK/Ep9GKG2/GAVXxX+Ic+AaX2b9mk+1gpP
f2JIOUZ6aYP4WqIpzUoqeZGRtq5MxDyhx350kAvG8X194hSlQCYxq8fb8gsyMtM1
gSy7Aha323hkpikGXh7ID0tV+Po2M/WxFG/TlgOAi4eY2sZZwaeozXqe2+xepetM
l/eWIbM3tmk6K/ogBqxAg4PHA91XPzXNEJjmHpo/qV/PoUp4tvR5y/5kPfYnYyeF
UqsJZtike8wYTZgO7HPTqkXDCwK8THegEHDXoWOEv1NDogzDoMjX54FoBaZhH905
7PSNqM+dcSpx5FDRYVLbqk8krZjMBgRMUATTlVOpBYWiufExl/WAfkIK+Qq6yqBm
j6ofYz18Ge3s71ASziYIGblzX/uwBUl9SLlvoXKv3bzR76sj83C9Ne9uTLpL+WaH
sNpeviCi5ghHA+tEJMRQ6R9i0PKU0ARecz1I+9PU+y1RxQs/O3AkA9E6yPi1Li6/
1VFYeLUoUc3yETbIkrNj3KIhNuye6Q0fdfNKT3NOi0r3dIkBPNnzopn7/OOCfG5z
NdTYFvzQfGYBfaJDZU4KJeqNpQJnl/I8aBhwTUVL4YU6P6e8m9gG+VDcwzLT2xh1
yaJfRuTZrXvF9yCQ5aMtIB98za07mBWv2N2oz8EzXghFCUwreWsJQQVfXU4Nrq3D
Cluo4Zkr+bdiNHpeqyt7eErpTxbYW7bdURcsre5wDo+mUPKHjyN65uQDRvKnhWs8
drv1ADQq6eaxqUsqAjnrMs/Mluks3L5BEIeJFFr9J2UTs19O+LWo1LwUHTXYtFwd
AwtFVuSNzBT3Q1Xt60kyurXVP9kF/AjIQ1i9FkUVDJ3cBtvkXkXJqSD9wENzAqyk
A7t/9jLd7MzucbE9FXZ/Fog3OdL9JJncdlNR2lCTZ6aUYs4w3VMgfrRsbi/ecyUT
WmcfY86qYKk20OZtL8FZ4mmiCxUmpNVRv1k39tT+plAIwpU2loPVeGZ1ejbJDiFy
vOTXlkcdXb5xHe4rUxYubFcpEqpsJgot7voKKRqLTc2Sz9LTmwPQv5d3Qd9IC12A
PxSjIO3LrF6SK18ltgLOMJrH/nZVSRQjhAaXDdOoXjAlAXR6/IXuXgYdC0ca/n4Q
OPhQrh6BpUxR+GkYsq+MsFPm794HLvvmmms5X5dDkbZpzr2iXuN3ugAHEENJIGw0
ue2N6YbFtuoeA4Z8wWizvpblEdxGNdsJpesqn+KT3MLycQrxkn0s7bhCMAc99Srw
8TAYadpwTC+qD3mrl26nxGPbhhjfcbq18R7rVdDexTe3QkEBXUY0Ro337PbzxMD1
6qpflAhfPr4vvL0J1yJea0jUCZ3PVz12zArOnFrPp2lkwgm8hF/1d9fEXgGZgGlb
maX+fC3i/ra9SXMueNKKH7JhZ6o6GkU/mReyl59PPlFrNnynoqsk8isl0jzU6qny
t6EM+TQXKgz0g8MDw1QhOmDC2ZorIl7bKQIuagLzY5STCDj4Bxy9GFToVubCN0f0
yZvtaLU6Y3Bfhc+aFsHjn3aIRTz8Ha3aPSr+kV+ReeW3rFXWGzEB8ZjmAbPl0f/j
ZUhYqdkJmlq4QL6HWniaL2MHjc1nl5sK7JAJ11vq0cwlzM1ueQPNGrrjBYIImZ+M
+3ZttBb9A7bBa/MaaswraGQq+2xXAbhe78XvTjSWFqJesJZagoRiDCAadvGO6WMA
E1z5WBUlpU4UMD+ijT6Q17/obr3PvnrbWiLoYlv8gBPHSmxKwfENJlSHnQQNvA6U
oecsQmKUZhLFbZHIRhiFjnYu+7OBppqUwHmJDYoFSrR/bwp1wPV1SU0NamK4yhXz
hZLWm2JBqo6xoCguO1hcw4Bg9+21HgTqejMSMLfNUeLSvBsF/avRCIc2Xp0lBnmS
cOSo+dMLg8m3WajPITz12F5sCP+Zar+xdQCj2ckNmcwgELPTPwudF3+Z/pbEcDTW
3e+dRG5PKKLrwcERT/TT+PmqO6HPML9aKSoR83xKYRLQb+llF/w09yV5/asz5ccK
F8BSuRoblq+MMSNLjEsFnyin7BituA7aB1HUA3YYyiuIx/Srj38pX+it6D81J+Ko
2V9gPE8juXP19hV0ssIyhekQCnibI8fU65l/tzYsdjOFyEVcF6qYp+Du4MhVK/Jm
Q+nWAYyfcHgJ2rGl/wDcVEB/nZg6lhyKuIUECT6YfPgqkuI2pt7ajj3pvZnQtRIV
/ICUM2q+S2aF+SN7XOxQbdj1sqXqTCS+H7wOxsbV878ZfSffzBpj1vsWbFO93C+/
6NRfWN9q7Ld6zYy3Oa45fU6VinohKTXmE6qvf7XF6FfYp0mABmyWQhBipgyyCXsF
h6fS0RrabQ/fPhNgaAJkhIi+AKfbSg/kh92kOnoUB+TFRJqVuQZKO3a4qCtxaqk4
Ok840D+jf9EWeoDu9sXIFiXV6oUKtuI7T9hrLFNhiMPzRMs7NUexu7bWRX2LxSgI
J7kspE1QyW8A4tgMTUx/CmuSA62+ZshSMqQV+9SWQ8KKYfz/V1SZ6mHqEX/EpBp0
J5jdA4kchoR561COa/k2K0ToW2+gvrSxalyl2KrPqzqw1W6zSQnqDox92ueA8OHr
Y6E8McZK86VRM3KLWdMSoFHr3hJcErLZ7+Jen8LO9rQhcrN11a7ZpRP/8PnEdUfc
lNI/RQVFFAFBkuhwbuCcupU5cCEi4HxTC1NG7r2dR/h2fbuaO2mP/1IfXTtFYMQw
40fdkt/Zy5Xz/lbLMoWXDLyZ7uElqh0s9LthKUJHHBREKKNRZlhwo5k1mIzpQibx
GrImHaHkUXQdS+ceZbEtFDxUvsW259FiCX0unVNU2ZIj5uqWLaDd5fXh3GOgH9hD
9fkAmth9cTiwNtTbhsBLPBts1J6DPvhTjyXYXj5DlNGGrN/CwGccwh0SIIEq9swh
ezHVoSl/qJnsNgsm4yJ2zsR/CR7rSQYeTTmkeMaSjIiThPhpuaDpZNM3rYGpcmi1
Qw3KR8i1+guFgbs/xCJOvDNv0Y0oFAPiLKzueI4BsS/LS4Y8MfIGCP5UOAJ4Nzq+
q56CREkMCEPB/jQJ1P0mQCeP5OBUFWUBz9FbsvPQQq4QgYaPFG5fVs9fvn/2yiGE
cCSlK55e1N/V6zdyYU2yqHwgCGrSFIynZTLANAowOBSfFHl/CWRyOabzVHKifCyR
OODlg6SeLcFp7PCO66enPKxreSYKljqEKXdVMeRKDpUiPq5HlnJJAUazLCZUX+Xi
dbuqKZX3Lj6BWOCro+auTNQjgzUkFKMl7JhnCn3OIICXt/KZX48tUknbysslb2NP
oXzkiz3KzS7J3pSHhL0KQppWmLtqU1KZ5qngF5pkMs/5biLA+yMFHP2hOxMbt+/B
AhCgDIHdc6ABZ1Lhm7dyAPc4Tteb/9Ueh7J9rYMly97PbrJSf6EMl0H8KIMMtSzE
4yET1DKjJfFdqIwAzBtw49l2laB7BEr0a54XHKo93yeLke4x7IMvmouKxyNkzRfV
UU0DWdlboIVXIZ+aIl6yPBCqPlb5dsWU2zDBP4pB0hihAHtdZVSgcjjWmh4Yq/Pv
A3WYKNKYEq1hP6FOCbjANGCW1qNZ8KfBqgaeKCYbzu7jkAC/FkpL4FIbHTovy8D/
5sUHyl528yW6MWlLF8eD2ejggn1BNZG5oryRw6OhiChArf9elM0f9hOt2OWbUiH/
xzFc+TNGloHyVUntpEN3UOlOAjd8vFZv2/5Eb/d//q78bppI6tVDcO+ZsRSmjMsC
yc9qk20BIy8tBV6fHOUva5fhdbnyWY2M62d9q+rEwHcKRQ/YAoDrU0LHteBeXCVX
fk3n3zZvBjQFoCbq+kGaoUxX1qJ0aQtCsS3cYr3rdT5Lz48c/oHx1FZno0WHERrQ
eWbsr+y9rZ9avRZ+UKKIPHds+3l9xMJlMCESbgaBGQ+ziHCfleWZybJ4wN7Ws6FL
rDu2FsGnTkIL/kbjeBGhl72Cda76Qnk6966mflRcHCuLASAnJf9tGvFuUIu3nWoy
tDNUVbKXEcyk8NfbU1uBD88npdJbm0k7PH3SmN6LkFwigKRG6RAN+Rqtdmp82Naa
2a3MJCehlZGb2hQhmsnTpyKp1AJIosvzubwBJoK8skOK3+bOeaNLWDhCFfs6wcEH
IFJ2uKwgxHnLDObWuRGbgQHroaP3zi7ZnHJziJKYFjXljYHzRoFsnC0emXbyImhG
ucrnKGalL+NPIUhswD8fxnKFWdwsBVe2aPXiEVcdTdGdiMxeRh9p+SewoEyx1kS9
Pd4thYYk2lhmBBXdNyzomTlKDdobUb6z72WEikCo6o+9PynrP8BtUoQlQJKbRR4N
t39209MMs27jKLxYAR8BGUy3UN0tP9OrmtPZw4qCZ0m5w0GcsM7xfnN/BVWbCad3
1TIgt/dTpc6UkLQWahOxnlBmcBsBc0Q/UoC197VjwS+B9z2DodtYTEOvQLyew6Gt
lSE5zISOvpGS0upFdCMskSsZ190prkeHYTkBC7pNXmp8vIvN4zwAPJzpKJWGG0dK
TxmlYnTXCmVDOmZS+5RP7ziJ7Wjec5SNZdJArAv2/6fCZzexk8XulQhBmsGXLIfm
alEZPXSJ2QNz7cgYLuPYYk7V60YkOC1NXf3WPqCK8viVxQocA5a9sX5TfEUA7mNA
SPU33JJD5zYT/UQiXP7oOIwlYg6xIRFTJ+5K+7M1kwQZUDZoN6MhUpV7tlBK0sx/
AOqjRRzy8AAcmXATM5I7XHosxIBAwdvh0OU6WJ/lW9GBdNW53u4YznAm5WMgZNvl
xsZQjOn9fIzcM0/4wQfvK2s+ol3Jt9rQeAEVdopBPYAx4bY+v+3fLfZCc9m0rma+
S5av/YcBmQ8365K6eRJlgg9Y72d5vDF29RC8Y6W9Y4OwOlUkgm1cpS3TgwsEPCLc
28EjXBO6ZWAHQJTFGTI/Pff70EiD+F0rdi9LYgx/ZLI8/0nQ88Tehuef0emFjs7i
SNNUMAEQK8M+zkQA5cq3kXsKMzmJ6ZL/eg1mutySsIf09hHgDEibyNLCdPmnPgbT
4MAaeuab/cI5uijtwuvwLs0Z4Kp7iS9JcEoSpDzsV6sJBO/IVaz1A1oTcQ1W107u
j49eN2YAjArxi1Zk2la51hRqsbV3b/Zqlx5pPL+vWwkpOndR7MRQM7cDMZbJFsfT
+nUc4q0ahhmL/Y0KqicdtUZjInzJmzJh0qP3cOrkeFfOjahMV70/Xy68Jrb+B2sn
TY5CH1EW/zcfV2/H7dSjH3b0mS+LTldYRSSLcMUJAYNfr0XFUiNc63/pKeucCZQU
GlhGwyNgCGttlsp3JpSvDRXZnMGOhoD7VJQTQFxVdcvzvvKgc1I55OdHbnAVexNa
MBdlkXxt4t27va8z07rZTV1bGHLrqVLcTLya4Iy9uoSVJaFebwRUPFFKdsYG1MzN
ekcpii6XZdhrmZjSH/kNUanJspFWh2JKSWpVgbuNCt4xxVTKmvJoBhdRQYtDHZP+
XDAtMSBVUw9T3E8c8hv7eQXuYabIEPJb9IrqWhQE/4Tl7P7ICDcpZAxxWolkJqD7
xGLZE8q4l/dGa0zeqQ9QuuwMF82Rx5BjVFFfQFozUaa9F3eenrRofxtn6DPr4Etm
YS4B09ykS0CaN2SuQpZ290eeL6+BULxS32obPgBSW9RaYG3+ZSa3kSw6y0I2Wi92
cppd/06yjWJegHJjERRxhYFS57clsQRpoa91hmw+PWFCgzyIVnvjEhd/f/pEQMJK
77Py3P5+jdXI6jlcDXUJE+i/ntLu17vmJlj0yVhkowqYWbTTt/wHySKYbTyecv14
G1q+Nz0AHLCbzeqsF9A3DtiaD8TzQgGfXWm96s55opXPWWDPQUFwQe2kUYI3clD+
4Bu0/lhQdaJzIhT9y4HuRV4yu96mzQmUrRnf9XM7bwKRkJaXS+uEnm3PxHp9rjmD
UciJWBu7WuDy97BM3OpIR0kjd8PEDSKSAJTjV5devM/tRXvJ/cRds5dYJVBYE8AS
xg9cP1H0YBYhTWfZVKDXqTyqV2MKfZn/qdaHWbGh6/udheDwOjctCyUz7h6GB93i
QFPNZujdgxNwXp6spFjynJMd56mjE2bpZyTlzzOtO93174luwKI8uyI9AX49vHtV
cSvPTn0C8lsESi03vIcBMysJi6y6vmKmkYsaE3vnwwL3/NItg4oS9diuD7TEQknd
tceMe9Dn0iaa1+8++sDQxJ1QWquGCjzfauM+MxqISJJYSFGPO/AHi4r6mlsL+1rG
i9FLDuKCgE2tgCy70UY3Mzauq1a71njr3dPGsEbgl9tkXXfgcSZcfcNT1+9DHQSP
dYFSsBsKrZxaqPTvCJ6UMCygDugVYorth1HJAQR47dDfq7vU/UyYOb952ksERYYb
xM58lny93gKnvbBjmkg8Td56DpIveWEovDYuv7h1QAtboCqqo0igDVKHVxPkkkaS
yUPdTBGfc+Dchh1CGOwGkTiJ7KIRSk/4+zqHhzUYZaFl0qs3VcJvhDfhFoPegzTH
VTpJSKASvprI6RG0uwPPYbQO06p2+/YwZsTErtwqHcPx0j6z3L1soV2b6aiO1La4
RZvSMvw97sEeVSb/NLoG+qqoSSYfFftZtMug+VFmZ+8WQBYvg3iT1GqJaFYXhZRR
VPCySbZKAxqDahktF5mA22XeAR2KBfDQGBGCu5ZH7T/gJgTU3G/a5TCt3FRg1gp+
7+f0gOq+MchSuXXlSLwqmrv/aT9gLp0wwN+NsUmc112xfyo19J31gGVa6jQmb2bO
oqgzL9o+U0dtkJ6MslRcCUH2D3jGqSh2kO+5AY0q3Xex04da/OxXUd+38UmPvFtg
m1x3oTUSE+WZzrSgFU06yu/CFrk1uyfl1NFzJG9Tmc/Jcag4MIq1HOxl18gHg1Ww
uvxxTgz8gDYrsFfrHLoUZ3m5KgtNRye8pbkXgvYxAjtymveOgnVzNlo+a3YdKjNh
/PiZ/c0DMGIBUSxIVq2IZ6jyyOkz7LVxvaKdpETvzY5uHmSKqBGT9norMvvTBMvT
qCNfekO4sHsdWqZnbwhfBxMc4afhp9SlhYwY5rPqzQet2c6ICV52R+U1cOm8XQWk
0ryzlLTUJSsNvjgMhYzNapwYtipYrMLufn/8NjXVPbXxNlkC0tJnh5WSQka3G4g3
G0QFA+hmmieKBQOoOquG1ucWoqLblmrWm2wJsVGMnMx6mRkm3fN9EpD4HCKBtndY
wB3tFQUChNoFOtzlQbvDMDASm6wq638knj1Y7dOHkqLO1CsJyRXlevHdkjaPkaAp
dW1JP1+7c+qt/3vvsYhaX0MmZkI5kPxJBrpzMgQubo4BHQ3csUkDt0c4BqkNj3Hi
GWHUqHVEZKd/5VS5yXsWzsphyIzn4FapU5vP+0YPMxQB1lGIXqfy2hBfB0Ymkgcd
E1/1MkZnXzM0SMqUAKUcxcohNfMStSKvEfQBHYjKNIfetADzwXUoWxDKSd9yTEzp
7bNO6yrerffkc1UE5LNa9bkd1pHbm0HLN+qRFJAGe6EF6fPaw+lAK50BYt2nHkBe
k0XgCLftMRCOJ2y/xEah5Zha/ZCkR3EauSnNTwnJMnSQbFITjuyDqquue50nKNWe
2StEFf/zBbZFmDNkbQGrYYw+QCVbrhp5ytEL+bmeCoSZkHuIzgZC7FzcmG995Tt7
ZtBTegh3u8G/WG4CDoefjHkZRI9obaI3SyJjrrFv1FADtWVWe/23/hgB+qWe6SaO
fiNVOIBezaC85UxuXaVYNjTRNqSp1MTuY3cHngYLwXe/BTATnhN4bpIkjdxU+Lz9
l7GYJGoi5iccFuO5r7Cek5Vx9Y2yE/AS6ZKUXcY7Vu7nUjlzauVWaiu3ajIIg13g
8EO0yoKozrgcb0y5GbQtSrJeab7pCyZpIn1TedmNWQG4gF5a4yGwYDs+tHzRFZpx
V/rx0KJkrc9Wpkvx3dDNEFJTrLGZaMDC2tAe4qkBSXOV7K3bA809FUEJzgHt9yyn
NeLNHwz4/oB1co/F9qdl2Wdv6/tXF1MFCaHpcfU4nM/cR7SB/qnuiTraDRkLa9DS
9/51nwb+tSolHiK+SgDGFDirkTKdthoZldoYGwfIIldCK+BD8evhUoqFYMZpFW2v
A139UwM3Ku/fqBh16CZq3r7yGEu9IzDkml8FyzB0emCTXG+EEc5PHXGNbm8GOpVA
jKqj1SRifnsMkRfaObD1XohmMhS0i/mrZdblICpIacQsHzM1vlXQgTZ+cfQxHv86
+inW9eUc2q5t3uHT/yISxRVf1833SgjJTKSs8fdYkRXB5mXKqPMk2ug7lUra19Ww
DqNZY7SyaJeTdKBXcT96VN6D3xSvsafou5+n/44MjI5zO+2otBB5fIAg2CTf2yKj
6yd1l8M4IkW3YyiIIQ6r8HPG03ovUtI1ZBPPqtmiqKRw71gPnVSZLBY2TSeBg4cq
miNvdtfPXsi74wzwB8ZPyTN1NIvmC5S0Xgx6cE3ve++MjRbOjQ8+EYXRSrO/Yptw
iLg2L7EN7S8I4blsb1YE9VzW4kIV9gL5r73fpzmQwh+PuHdOh8gv86zrDIl9JYlU
ueofjm7hhDnZSz4e1fWWAKRHcLMBdCPMLfcRwiYoIFoDY7Wfsniaxt51AvCAHvCZ
82xRWl4B98nI7yZ1+xyeaQjqlTxcqrpdLiMD4fjDBDY5r28ePfxUr90aY72jrLg0
1n/gETOYVJh60BI8J/Vg21RG6ryu1o8TgeHuwcALLPrT5S5f8+46QvDUWehgBCg6
6brYraMWdtWVCAJjgjNOx0lfXbM21dpOPqXpZNx9+xQ/pe4Ir5f/JdHma9d5q3MG
4PtwdAFq0Llgxgn9ap90RHpxpj2WPI88ltJj+Q3iJwPnKmRTqLR0jezifCuBT/5n
/spuctdbSW6YK/LXWPWdig9hOabri0UdLxYgatBbs8kgmbGOctT3TpNklAIZC0Yu
6XEa0Gfgl1gw+64FoOohptrhSJUBsEyNsCAGU/ZoW55+FRVBH3l+MxFLcxg2+t3Z
KEPWryb8ZHFnVugR4TtXNb+xu4s5RWzru+TkjvXP5vIbbQjBS8+KkdfSLj58taHT
rbdSOSoT5mCWOiEiMluA/9VZNAemdCY2T/1947Uaid0cT49LFmEiY4jf3MM3UCHn
kK7zUcxVcSTXpLAE65ja0DTsXS23CJgQB0+lRvIsRcJzXdBbR9LWDpHs+eksPK8v
jATpz/Zkb4IEvOJEBeHopdPoT6gLY+lwpsDK+hAOgegZSILMbeXo2txJlKemQuXr
9oPSUgvaMgOday0t1d8HL3mQXeUDEwBvOeoLnMusEsoULA1qgsN/NCchfmtdR4lo
6oMLNQmX1uuTmAD2kpieNTij2UT0DaXu2EcQkjnjOe0EE8w8R+GhPA8z1O/Rj5iE
PDEmJYWTdcZext/sq057sgfFx7DtUngSbpg7myGP0v8UxPJl/ZNLcmoNpFmc+Miw
A0KC6VaHPAMcAAcwfpMuDlQUJpsZ9qcZSMyMnfVAYeCEvXPvlsuO+nCV2BxxVA/Y
GYHTLdpB+c8l7yAxsjEEqm9kfDe1DU4AeHlcat5rzgou1cjwb+L3z9SBseFq2zJL
0hbm9UfvtsoNxzqjesJsduWGZtm8CH/pEAXyo/H3FWu/HokEXideWVKeMZORXp1I
ckrx2u5wU2sGFTXfdnZNdDmdN6MCEWsXt03Fhddy8Kg1Fe5/JW/U6DaWVU2SIDRr
uAd9Wtq2kLei/5YJJjaqjnj4j1N2XlcjJWXUHcnAxrLzPiRDAaY0Thyvf626bGuV
XDjL3J2YwIMCWPTtqDKCUbUdddC8vfB8goyuvP3gZ8kyAyeqVFUQYyvZHVBulRIl
Xx8MTOEnowxmfHQt/YMfaNJdb13HE8aEN4eev/IqKrjArhvth7T5WZZCt5vH2Ocd
oEXSSafTSHe0RySz+ucPf5uXXYVsIOgRWZFXkB1SmZhf32g14WYppqK241gGr6fG
39bB8CImGinHB5h+AnbjLyODr0Gr/edfIb7sMMhid0A/TlP6Urza89vfZwQL5yWc
CYtl4rgYeNpwqTrf2cm32mxkfYeK3ndvYmaD6VMP/jXWKGweoJvN+vDkHr0SyxJa
PhkJ1ss0s8cBu5A1ipp/xggPbBPYeB0wsQK78WnDOGNd7W4Xbb3uKIyvXYHxDZkT
BMd7ZStstQ/zE4gn46PuyHn39KG4BgINYE0SuGVFtWEJRH83Biz86er4L0rXaf30
CKVsvrKsvwVSQFGoFKwW0+wVmYso2D7FBWTfiX9/r3rl9MBcWWQhdllLiCKzR6Bi
aM1lJXUTCN9etmPUnZPkjXZwP+p08EonyZH0MYG5cRGi0FSdpzYJSvus1TFqvwS8
4h+fkfhQRBMe3B0XKawdHuKgKFtNtPlSz/jcx/DdA+VyyDGEerxMGeQOng2iZeV+
Qbb0kh3mEpr6pPjPl+xM0xV7A96fdTpYuMx9B6Kvc6GoBjbPMbC8ZsVKRl4xrd6l
NL0aYV0QC1V5huGCGlMG3BCV0cmhV5zZMtl7t2dCOdzYN6p/VQsHhRap4Z6nYBbX
zQL6GLb1d/VeQWptC+MMLE7bKXdTYZzwR4S402YTTo4mdaRlnDp5vqhnXTu7xFxy
H4GQnFdtinxJxGostpACE6O2/9wczEg8ihLlu0gaXeJBgiGUd1PN+TpAmg6+115s
4dQ1cRpCXNlrxKOha2fczsvdIWEpp0F91Oj5DjeQ8olof5mBqOXYkFha9yjQtcji
A8z7uxMYRLqxfpjyW+HIGbkR5IsOV9gkcM1dF9WcggU7jaMCMxXPjmbkXxiUoWla
CgbV8ffrotN4EcLZokf+2Nxc8yXgp3PUzAdS9Er1SsW9J+qPacSamabz6hjbBUry
3Ge10xnBoMl6oNCeH3RafwS+7vUmQZZHd/BPVPhqXgISMB03XeTnqmwXNDAgJ/51
2J4cUXWthDb7SOLkk5ta4NLn3IZXu72wD23rWfvClxvb+6VDejd+OILYnbbRTReN
r62wHzBNlrWl4m+nUROnRackWXhJh8HX3MQyTo84nbFe7bJh/t4TfHO7L4YRRpwM
3Rq0CAvUbZNIo+oVSz42GSHbF5BYoO/TTQsF7qRwxd9qetZGlGx8axfykIrKk9nn
SZvlMCGr/mKnWSybdHBki32zMatMs4pXve4SBpEdIQEk46D+m2ycbDvic835fYbb
yUU3xf8wwaosc1kD17RZGcLs+x9rYiJumIz9WxaS9kNWfxlf3XSNzkUWoGgsDGzX
NdlGRXNXW/9nkNjx5eetjZU1S6WvCT/kvWFsUo7kI5/yXBbFDhGlFG1kz9FMdLmK
SUzLnxb7uAiSFcILc4SxKVSnc0wCIeSjhp2arnc8Ziwgr3y2ZoF/7ODw29IcvIAY
zghYU9uKUPgvZqRO5HOIEuWYH1EhX4pOBbom+UEh6k1nMGAn6VtIej97x41URofw
MEbLM8g47GeKmrnU598/zlOJz2knq/qedgFjlSieVqo4eQDOAz6ziPBwY8JKY3Es
l7j3iIgiNioMO7hxgpE5P9H2r2A1qVJ129Ny7OkxkOoiLVdySyetTAGHv4nrllTx
0wr6TBmVRTHJ+p22c2/Wky1mH9eUI+9HH47LZNqLYZDazGNTyItMBI5+dqi9QHwe
1RySo2ej1MsGGWyv82gXSYMH9baAkoM4G9tGm8ioP6Hw2gyUjRx3Lj3QkD4oBOFj
aEbOHIdU8xNZKMRHmOwB5vS/u963SwwlPvjewNOp3C6cP26B23FKK1qkknk7LL3D
DpHhokYNlYLWrtLwiPFpE5tQjFMjB60MDGYm5J98UZ4xtCXLnJOD+LvaIBblwIop
KT9pUzHgjY3wysbuBqrfRGOoaSFsStEv3Y8RgBfqOTx0Y6ENLimWQt80tlMYN7QW
dc1OK9bfB7bRLFI1cKNjppLgv9ohkDSHDbmqzeyoSExLd6r1WY5JAMwfhiKNcYRB
1/6sCZ/dxWAjxBBmeIYQI6XGwC7JoMpENlatiYOVR3TWt9WsN60gfLhZ/fzmUyE0
ZI1CPG1Zw+uPB00GCG4yrsvIrqmQsIqHa/5I4+6rlMpKj1ZCX99s0GQRwZgw0myx
HdCbdu2DmCcHky1ynEGZg+n/8VPPZexsV649bfxGOjJAjXOLACfEQ6mvwrVTzl/a
9EDU7+aGwdoJmIby+zmy5++lJrPauPn61Bt/emaHY2WUUn/5lqCmcXO5Nv+2bLmw
n/ebab7eo5qEzrotnx4MH4TBdBKARb4VhaQ3a8TZMJCr1gmU5oTvdsni1qK72IOq
OBOsjZzmQ6dze+Q4xqj5/A==
`pragma protect end_protected
