// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:02:08 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
YjacVlUoj69aZlBFunzqm7en4d4Sg0yNdtpEC0YMzloxC+dMyqrlUiOnlk9SyAxe
QXAhlZhqvgERn8eb+RIPQdP+V9+iFwPlbcLZSpPoPUYDQ1sq9hdnQbhGtD5rQYC/
kKSzJsHln0XmZnSllzYUaqBHDrjdQN2cRqGdYJzHfLg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5744)
FbU/9sHmqIFelfgdjjbyOvGTr0dLcwXPA8zBH1EyqdDq0ycP57pb89RAIJfrgyj4
lYZC+XtcnsAzdwTZF7iWNJnsSaptfhX+TP1KgZj7IWYvbLOS2z3DPd7/1zEAJTu/
B18LHZrsRPaQ3nCczgPIxRkpj2w7wFEukXNjHIHWfMzNhZXK7JfdN1r+Cpegz3AR
ddKtX/+WPlOUCwGuXa+lh535lbtAv0Qufe+Jx3eAgroUV1lDhnphd520tFqmdOrW
wCbMDTIwgyft9ivOQqs2gUX1t6oiTu8EYSTUZBQwsMJFFfFbKtM+CZPbIGIGaq5A
LxXtZF5+JQDfbeDmF3tSNkXWwl2xBpoF54g1gDcMQl0+zaFS3VeDNxVG6pMkqdZV
ImBYfnKsGY4VmIjjl/XHeyqiPJnSVhfqi1523bWLUNe622KvHED/rfdcZXy18hnm
QqRT4JOs+/4xNKwYZgIf7OZDnvYQS8Xiajo6St8c7oGwkrBsjQaR+ZbiJg36MEh9
Esa95333kHU99Kp8FPD5y4kT5q3sftaUq70N8SpH84kdSUTGdw/5QiRgbqA/nxcn
GPGi1hwsqWLfr7gHLie16GAjZ91ksWxC2Ojef61PTtHD5aSZBaNY+en+CIBCkvhX
uIb3jaDiGPEe/d5s7BOhOdSnUHv4EHUKGYcw2ijxXvTo8tI3bSaIQoJybe08xN5i
iMG1VlmQqFwf5F+1NFnA67rd9U3Yx+h+1ZkkBIRVXXON5WGnQhe60thk8Rv6TiH9
bK7SSO01VugIYKHj4nP8n2s1/U4fWXGgJIwXobTdwjxG7bepGlUj6AjPFe1te+CD
2cHIND4yezuvUWZOLzNKDRQJZSFmefQcge5YqZP7BWo48tZY1pPZqlPxL7MQwFpN
9zSwd6EwLVONTkksGZy5rAmyg9EynQ53wTThM+XiaZmbRBi2lhq1dqZrx8KY5PFs
uu0RIe1HiL5xNDa5dZM4DWiWh5Q/QpHaL/YBTcYkO1Hv2oCsekXZvvzmy5U1lZnH
xoVN3DnaU4LL8t5ucGk0+3JxpcewO4Chb82FdNQaHRsJw7/7AG7W9HzIGlNP0tm4
jP26YeG58y6JhP9ly3P2zPLp2unK6V+jlZCa0dCU8onEWkuFpuM14y0lijp0Sohc
6q+lBAO+jQ8jcqxT/GPBaWMCUlzcPig0x4nIf8RbVckYnuvEPUrOWMt4Iwp3ZNRZ
y0D6bw4MA/BqndTA5/oXS1YkxC2znBg+YM70Dtyn+Avjz3gy0l3/+wZiLKMZZmQ7
oZle75FrLlN11gCAVhIWKT2ugWbesUUtn7iakGNbcIzYHz/L/D/3/46OG5tIQIWD
25tmP+zELEDcVQtGTT2zNsb9v5zAB3+2rE5DXYtzqC/VDANR8Vj7qxPOLRoFcl98
RKNRKuUgkWOG59I54VbgnZ8YPRtP0guEbAE7kOvTe4n3tyz28NbIQ8mlSP2q/Obx
Nd55BTI/uMqOJZ7Rh+ZPQF4zm+NnxbLyWPeI1A9dQABnpbtGpJUWMgLYPRzGztfV
I9X22IOf7kU+UB3iybJxt2tdHg/F8UQ82KRs5Y5YY3C9pa/8k5As/yDoqwd+4Wu+
Zd72pNojt98e5voR1OYeJ7MpA6/SPb05pYbFfx4qwKmaBm6rIJCxQwbsxA01SM36
fTcJTKQVBP8ZiG1+rotQi0LUrZ1UFLO9pynIm6Ev7mXbiDBbGzfVaO5QO1PcyiTW
Tk10cKoitzOvKtgFKVTo5fylJWRSnkA9hHIJwBbxd7FF4GtswkV+WJn05wGIa1jQ
LCNG7kruiZ65FX1wQ7Hr0wP2z8LBvDBD6nvlBgkvFSgMiTkogmFAN5M4yngPc2Yj
ZSox1JrdEk1JK3++PROz3g7ghJ6OhaIimK6jJH6UvfEffk39ippVxFtskj1xOtBH
9ySUzwY492qw8b90hQoMqLSybgCjiQFdn+p0dbsK33sX+5zUQwdqlfR+/MGYGF8h
BDo+SQDOybj9WhJNy8HnfkFSu/K59fwMkJsFUbAfl4gIy4hH6zrkJyu9c3wUa4tt
pI30V5bWXMuya5y3wE3Tttajkj/Y7suuSmBh99au4YK4XIbMbavF/dC2s6O6mzvg
C6cS/h1CkxMzUcaBmXdwMWefO5sL9TA8j1/S/XEjHiyq9MFP+Wkv8TYziPca4gaA
ezn7wM7Izh8bwoDcYazYICCDVtJ4dG+B57UGpVawNys/0hg55gBwjBW4/+YcoNda
RvnL4l7gFZEp3ZtiSOBNs2MmOr0h1VRFBJjCpIRjV4mfeTy6O6Z9kLBpl68p9vR9
25m+SETAR0JbdUsUoxLUeHiIV9iBq2MioP7vT85kg6155bLzW6xoxKMxu9rqhepi
1UwG18j7rt7Tys+VFwWuCGqdTkg0ZSYDF4qx8XvyS7G7MGgkHkNlmez3zewzK5Nc
cOFAMNWh6ZpppsXil+ea0pVNeDVP7WFKcXG161H9pp1QVjOU+g4wtAfuWuG8+LMn
Bp8a7i5udqAHBzlebPx2H10Ka2V93kG7nCGNb1rsNffSzzWg3oeM9O0yTxaK9eKT
n1rEWF9y2qZcUDonJ5GVi6V1Ft1zlIMyB3WOlxwtrSv5thPUT4KvinxLBLbJZSPT
lr/oZUpIXSd5t74ch39KEdgVIICrVb4z8z8NbfKJ4XJtFjHMKTuXzjO/mlsTfAuI
9OJA0SAIPXBNAj+ByOfi4AU1tEPcopRM7J1L2wbxn4RgSqh6kfaVSUskM5EntiHU
KVizSLCl/3Rl8Auy1mFJpeAPWR5ad8lyDliEjK4YdjQLx1t9vFh71C41bRrk92AO
1ryKOPusUWseUNtCNaScr5rMjYiP0V05dh4TUM35X5gQpC8ZyOD2/uXItf8T7bJ8
GBjSelrAD6CDdZTI/W2IRDd6R5CA6soEvGDEG8E20WzWpE001m2xEYHfnuwLq+Lg
fFYzK6a5EVwL9ANj82ZMlZz1LUvzwAPtFGS83lvWaWC+76vtSpdRHj5okkucq4pb
ypfj1oM+wWE5jDPtIh7dvS4DRqznCOY4s/fEydY3aTMkydXpVkDfMwGNUeHcHtxG
2mKWGGdFL/tWgr94ZTFHl/9fLvDe+2cT9zSPPTHDcnTMMHJeGlKpBdtVXWtquso2
RbuiCYJwkFuLU3GYtq76MTxjCdg5SECLrkEwe0NRAVZI6CMb9Lm80YW3wxonnsPL
71ctJpQ9hE0CfflVUvS9kHIMDN4YZmZBXVMZc/nsIDd0mz9r6nPLdBFLDSqDIXOT
m8d2A1AtB1uoUQazmM0lg56PjiWoq5xNJOEmGw1bdeK+lLic0h3k1WgzIbf9b0yt
0cOm6JCT1kfMSGGWvyoEKfU9loiPSedpyw9V4XY19/5/1NCa68XQcMGzOgdsafP4
baHVP++A9B+N1i2I+dGmhkXcKXz6Dz56z3zb8V3wn8lIf1hxZXnz2APxyQTgzjSl
DDMRqMMsecXwIUEi+e7E6S6qV+h9+RS/gfEDLoYC6T9A33wh9JJ0gSVAMmes5Ytb
d+SJGJ/fgLFYnWsb9xWb05ndP5Uv9uAT/nDrkfbJVSicmwcVe9msEaJbzvCvqfAZ
Y6Y/H4/Z4czBww0/x3iQ8AQUnScjmEMkL14pGjkXLAtNNOx4mz/7BE1EVv4YkulJ
tKwP1V/4KJHbE6Hb9h0rPdU4wSxXvSvNPqTEnn5+yE8WFlIb6yc4ir52z5GjOgvh
UfvVX4/MV5UD715SxcCoZcHXyoM0JoXA2I9Xjx7mjIVg77J1Vmx6GL2Zs2+QFCJx
nOZtKckTaQa243SDNbbBt2nBsjOe3ydJbxxJVrldT9h7b9GcppGU2wNGgW6mendz
3LAtNZlm6+7UB4EsdmSqyytnStKHsaD3NzxvIuTIWU8OZl4fWsTO4S6Vi23zKDz0
VrChKuwOxLg3IUpnFLay60+CI+1gkHP2tkxvE2EOHK6vYEnJDuOhsnJjEvHTOEjV
LBNfb0kdAwP+93YA8JG+DwF0t06KtqHiiyIuUxrGAy0kSQocr1HWm8TBYirn+1DF
kdmAftUuEGp+4pokCAFos0V0GRtouk7lzCx765edff+yQcH9RQI+zn+gR7eijYI4
lhP4wmKo3/Cl12oIx41l78XL+qDbEvvoWg2M22/uj/SJeehRfmvIYtM8QCbr6RE9
fIzwnUmx3iBaBQxhzwl9PUlCtiQFeFMVlyTmFcDnQaLLDwEX2U1UsIXRfQ+Wj0px
t0GyzAVLzR2PTMKaYaz12RjzHKDz/vy9qVb4+bNWhf8TCgnj1p4kTSnVjg9Ah7kG
He243WbRmBpsW0E0uSj6p7jMDv5i+OdVG3Uccq5v5IjjIOJwLSQ+6cSSLLU0XCTJ
xM1gYx6+fA/Sb1OtZUCZomMzRo4Z7EazXJtEsoOKM6Q0qhux4Ex7SWtYQM9CK4VU
gZayrTXpdHYqaP74Uw/5RIhYoqepzbjRd15XPaWLnR4o82GDWFvrHbUQ08f/NuXK
rfKAFpjjn/xHC/lWhofalOccsPIOidsB9ZrtCMM+OwJ7GzTTVZPdZm1boamHuy3H
SJaYsdI9E8IQ0twMiAT6o9EwdRrh2TAXGr08gbIkuWYHmE0+mk8qOeCMGQl0d06+
sJo8MwRA9Vjug02WnxJkkNhRZTyIQZoifFy51y8UAKYTsvTDerdU7epo3vuGeGyo
TINc8tIfzuRoE1gVeeeSM9gs7CGFtvoxDtMvCpqRX4VWGi01DnIYfwJFcsf/rpdB
cLi+7A7ZTO1NyhVEXBjURUm4UQhNBl54jGhvlrbv5XVeno16QvQlBfWCftYsX0M8
lobMVOfRrkld7tKUtlQwJsRrmGjh1VWW2x7LNlA36YZXp3mkNVppBxmqx4LUuwly
Rc2X3P6OcnjZTSUQNk6j5jMQ5PzzFnhUCOBw8t6di9mDtZH5C5cyEiuRn5HsVD4j
VYTCbRppCY5OORyRcfudJsWrx+m3MyHkmlJIFcKrcKCDxJosm4Vq9QjJixMp6mTs
LC18Dd3e7DMQoUlYMYbHXQr5NXU2hXbME2eMBILI0Hoc3SxrSamAzwfFpf7ItLqd
NrLh9eU8jaNZiWsvSq0nsSjL3xnh2iDJgBkwTFnaWkjh0gBZ1YCa3LlnfEqlwhI6
K4fYt9CiAkM8qtcymf9C69uVnHJGn4Ql+ElrjqdkVC5jTZJgzwFcARf88+RihVC0
IUoGR0shZ10vn3rlqhXTcrNRESOhnsrfSWVp2PMTT5Uy+UNBx315APIYXS19WeAk
uMZTdHYHml2/PS1T4aVTtGkWqUxz1Svc22ih/ucZtQ2Z0+CJq+RqbYLWUg6XpMXF
y2ImON9Krf7jtGqqKD+YSwwLCTeAb9hNVxQHgmv2fT6jOZf65t6U0DSJk+9wGNSg
ThAgQOAG8ZyvOTHxGuh+YAu9Yr+rcqtKVFeFob8alsdK4YxvYJ5DyCo0lKpaVlCq
95Kg8msjJI44QjyJSGjjWIAyTI5XPbPgshyIqaIU5x3f9FLEiVahgbNmTzIhR1dK
XUcdBY0PCLOM3JpAPOIEoYmfkoZiMj2KijdnOoxdNsbAntnRlOxxqrAZTfgH8KMx
pGMt6WnmpAsd6Av6R8jTgDmY+HHL9kICJoLaiP3bf13inxQeQnhrYfgphha2oSl1
OVqs51wbBhvmwksHXyqpnKedhtnSgqogmqj+ISXOrDM/h8CdkXveJgEdtZ2lyHNa
tJehU3oREA7LYmfBN+CN/7Xs9nvIuaR7wyJewQTo5Y84olJcRxiUWXsYo2UCOaT0
qCWuJ0md71esMnqh3IzGKujb2HKbxRtTTB5GWvlXAo2qN3Zcy4yhhslWQiyKFvEP
5UgUDlRCueTmZDkJq3MYH30MA07/tXwM3WXxBLlRzzg7nxnqRXRhAFuzweIVNojY
CPiKvpt1zitDysjiHO7YZeH2AeVAziFFyU4XEjLXMy9iN+zk49KohiAaMz/U6dXz
EhAECWzZgyrpTpbtFdrl/Zrlde4U+3bYGVlHl53TlD7Y10UV7zWXvVPAElH5zFof
Z161K4j5mQ2S2yepHkhtTS/e/UhvgWs7WSYR2FswCeu39cZEHkDoC6lIhZGSH2XJ
aOhV5gs5/reKJtKcReGnGgs+lMlpD67sOe5gnoVQ+FxN/6CzC9LxsLwEmpiJoldn
/ylgDsr2FJGca4cUQ8EY11ahUtupxT3+zH/tY6izRz35bMHaamyjLoedGKJL9MfT
pWMwfEsSsyN3WSOCevYePunVyhqLZXhSdoUtxcuIoF/6tImrTXODDGu2NKZfLPom
EMVUhvjaH/tHffwGexAfi7hw8k8bQtyAgh6lOhgc+twfZBidrq0g3uYRCh14cP4r
1nk+z8GKwSgYX+WJjKNlawDimi/bR+dH+YMOs2dI+xFJhjhH6KgCib8h6cJEeQWs
1LNhuE0yYMO1WRxpMtHtzvqe9eq/45VkUAi8v3wSM4HQV0Dh2Srd0v+1K9pcMBhn
IVPQ8guS+YUrHEmVp0PLBtJyHwbB2SkLl++6p6iHqq1eLmBT2BsRtyLGTvU9pkDH
+5IoRCefwAkieGw3K12TqY70ZOYBOdbeVmu2+K5fWd63NCgqkWoApVSIccPHtIR/
FAR2B53eXXBiQ3gGwJdBgF6VAJHtYB22o8Fgouk8qe06zzpNOtDSbTb2pdmWuwfw
5VbRVYPVisp/7yYAX1F+cKYWesAmzW6o/NVfoHBCLC5XwB3LyNswLvR5ddjzCEg6
ZMZcrHxopTdycZ9Y/NJn9l9PCJ9Mn70oc7Um2qnHDnO4GA36TvUJdMW0il6p42RR
PN5lg/FTIaB0DdYBW1og6+kOHWaOeVSITfYeBplZh22i/MkHoHNnyic56Pw7h63i
Pqp4bY1h1saCtRNskIPIacPCKL0EhiGL9L8cgetNgBX7c4NEM2kiZNmcZsgD0WfS
3LLQY5KdaDzR3dxwKSeaN7jXvgLVVS+/CTBlXX7f/PGN45tepN/WR+oPDtFnaayK
qCZqEpuI58s0HC1QJQMYjwDYK5SKKCVMgtpY8oTwGOYiBWsn5Z3ysoHFu/GaQ1c/
QjzbLwA5lGqG8EKFJE/h5F0fu/RS8KplAf99NlJT/m7oaC82JeTju3mkaMP/l+6+
i/TspDpnBLWsPb8ALKw8Pl1F116bthMtYwNh5bY1Af1PPupdEtTbVv9/MXJTh8y6
SBJJQpcmSQtSK9uLrBuYEqqhd5nUr8sPqBp3TLkjbRLlY5naSpORxDMH+hWXYWGt
V2IqQ/S8pTxcgg+ClKAe0IJGKqyP+s5RkvLmt0/ZO/T9gpTD9EJpLp7nDw7UnT0E
M8rZxZluFW02cAHPCHOl+giFiUOtVri1Iv6PFh1mcQADr/nSyat1bS0yX+S0Tgqm
G5TtWBZuVEcQdcFv+1B9WCNucSgxcMuvnWzbazGJyLdSH7tTDb8GCAOeIph0rbJv
oHPxtALZdLGs/ZhNzG4EZuXw6rQxKCLZ/O332EdNj69IWiyv/Dzvlk1ztUMsIKA3
Sqn4GGdMGS3ZF8dWmSFkzofSXer3wLL4mBDjBN0mUnz5z6p2AIBIarak3s6yM+TJ
nAAiCp3kR4ik3oOlMAbCbUOPAweo1uVfGfWnOz96vqRZHAf/TTPb+Wfdtzxaeck1
a1NvzqQRNUT6EnBWWjCs55X2jjQrj1UZmuKcFIpR2uk=
`pragma protect end_protected
