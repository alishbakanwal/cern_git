// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 14:01:28 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
NnCWxI2D/1Jh4j5qw0CszTZTD4QxhJpHfeGzdJnYeBxARENMXmF7RhZHKCjtrgZz
CQnFi6rcKm4NKyDZNYx3OywdfwxvMuzWJFjWseSg9CyS+GEbAKpQ7ojL/97QmnRb
9/g7EwZDaY1RiD2mkUkX8FgylwmgFh4LAVo2Ts0t6jo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 4416)
TN9F/3kWGVs39WqQhW1upN73RKVJtgD1ZZ1U7VonLDbcEJjE24TB6oBD45MucqAp
JLSgg4zarDZl+/UMnsJeZAltnY/oGB0fYL5YuU0EIMbFw/yXVv9w4Q2bx5fQgw0w
UjfGHGz/yLeEFTvUDFJ1/nGmNufltMZvsm2fuDQSa7IFun7TtWytSMAXK2aQllSL
yI0tW7Kc7dcz2SyDQuFkjXmypF0/hWBMwe9WLaz0Oket/dO9PbQpTCsmzvOB14O0
jGgX7j3XelRJ8dDg7FidAvd5HzpdPjNGG++Wjn80JOkmRiEJVZN21WrHSWJDBBf+
CyuFm+JNm5X/3lVVJzjXK0ZRVBJoPEGgOfAklHCy6J7Xd52IaoqPsjh4iGJiWtIN
gXg9/DnGrCdMpkHOY0DdXABeQtDd5cmAAA7R+QL/BPxZ4O8r1SgL6g76lsXKOPwu
87G5LWXirwBOyr6IoCfeY9j1eTWQDTe7mhWXrcG4OaR5pivEwuoZ4mADVhfdGUDa
eUW8/LXN3U3GwvwvtAwa+HDhn3x8ioQEw/RRmIpPv1EV3S1r7HJBfcP5pn9IwMWj
vi+JisEKybjqRBM/eIRlTBF3Jjnlk13AqEj30gyJegYlFGQl86d+KMyp7nNoQW59
D4Hnn+DKi1IMKuM0/RLWZCZyMy6s7iSFvarINIMVEB9gD8J5FdeCmfIHZMcMfmrU
Beo9rdcgJJjv7SqDdrhcC95Ot1SutNu1rZpr7BL0xWmY9NHGFu7Wauj01mjd5MmS
L+7hAYZTgPlF9PXocu9du8Rru1wBHNEnKGDgZPSLHLvf4BjonVWPyLrQQLJ1WQt2
IO0vt1hzQUrUeHs2HRaBWA8bOMVlnHRy+6LJ3jXjb4LkpPGg/iEYvj8hxElwHnpB
z+bNCk57avyFVAclfor2Jf+jkrOw6MOEVOlUp9QUztUs/njAojl7wTzrFCPDI773
vFONAdDUbD0JFqGdKG7SzEAmLbaULki6OpEbTgWwsELrFrirUTaY5b5+9tEKE1NL
Jb9AXasY4dDIRZ9eKa1hT+emYTdfwOZZsbfmW1Idp/D2AbPqCY+h3TZ6Qy7Caxxs
ZWAliPSL+I2Di2JbRnmBw3I6aFs7fBfSrvJKb1fp9/zEtA38OIN7k7HnP3/aTI1t
pyqEDX1BE+JcyWEf1SlwX7UlPK2MAi8w+/dCuwVwR8RNPzbr1rkSrHsa5ld82k5D
zOrLoVdL8fR3+W5oofHceOFhm8M6o9qAgQ2fxAX5e3J9cbTBSrIgCul1pe7aXU92
g9x27U5ZTiKcHOMnlitMO8H/EmFa0cW7yHcYik6cFOzyEQD2Tm/E+x8pnmnKtUOt
ndfGG1PjU3UcGsyFp11XdAYgIXBERZ4IGsM48jOs2/0NxpB2UWuDHwv5rhjSm/SY
rQby4vTXa5OZNqSckeJFP65ASpp37obNM0S6FCoOTczS1cTqDAyA8Vx8xCMXFmkl
+bnAcuV43on8vY8xr0BmH/kx35Ii4v/Dm2P/4NhWUlGoofV8zWBnQI3y61iNY3Uu
nLr9JmYNJRprRp5GYSE1OiWV7EOjWsXCwoE5tuDQ+cyxkN7SHBaBDWeFjOL5L3fd
wlZ//xYmMOTfeaUUQqXojPVqenVbW+LuDBlBJhiuAu2Z+WV8rXe98fQK2lQIkjrd
Y/W85qoN4AB3ZnXqV6haPIiLibKhg1gnhZObcU1Zj7nofevgN5jfMubYrQbH4wV6
5RUk5tTCj0k+uetowwCJ21xHxyVl69etLXa21nBAAsHX32KhtUSVxYAef14P6RZ3
PjqBtNyR+EFZDk3Ke3For6sAWkeHkHjvMN/ab0QJaec6NYYeRJJaEha15uOiiDl+
rLdEsX5ulJoF9wiD7TBS0UOLCv+gqNA3rOgIbCToog1IaOGopEIpEky711Bb9I9B
IobW2VqINLobI02DwzTBPmnUe87LnRmKoNR6FXIiWug1gFAX0gxsUNLjXocLFv3l
LPFemRyJKuAdxN7QN2VOFC1olLHaC0C0zAVclkXpcfy3GM2mOR5EaIg2BoMC7pqp
z3t8RDW2qNI8UrfyV4kwFuFILV3QBYdIye5a8tDE4+CjZWFZwdBlUSO54KYuCOWF
PrF357uXEk2jEVdZzhagH5J1CbwvNkokIWu2sHR925M+gfoCYadRPLWWSVefLlh9
Cu96IJqy/SIC5vJ/xb6ySU3FfiKvmZAPjCC414A2t1yT648nJdQavNfkTkB1OyBi
YpSMeNMOpRx0Hs4GhAej6YlNT6eOe7oA3hx+j9JJnegu68V1c3P3WlZltb6cgD6N
UYzWP9lKayB1/vslxqyDfXWtnV/QRPf9DEb6sCijjh2TPFVxT7i/JMeXbq62xdzJ
aWZNFZHVEk4Uocexeuwq3FjlxKDkRN4uAm4bA4LnhYBpZyeb+bB7wZCvm28mYlZv
XqNxh5vCyY/hpLb5lJvgy/8Ti7c8YWN8TBTnsQYIxetzcEETtdT6o0qld7pewUf7
CFNcxhNx2kvxNES3y0C7kyffWlmm4DjqQEzzAL2SGSy6Je0WiefufjuyABf2zNey
4zQrkQEwf5bvLACkSFKJVCdIE+LCsZ9csv+j2n/H4xYvzVj1ECP3cN47+HrUiCmW
jY9tdjYs7xn1uCqvNOLLm00mBWU77jXJz/75VzFZxU8NJspf295lqrVpLE7qEm5H
1hBa53BdVdLVMnhUE8acPDdO8V8Klom/Ix7jcThnuDl5x7snE1W7fiWTUFMXZVag
nVZi1oZGNwoGUrGov/1qU0avyqsb3DrZbeYZl7y8ebNGs+k4+bP0OO74PooYzB5U
IkNsdzHhOmEHaXVjZ8qBpnXUEZoCV3rU+HVpf1q1XHSL+8CawFa9y0cRJC8I9qvS
xRVe8GEc1utk+aOWdxjeLRu3LGUdJLitBpL9lGc3HI/gSwIBOEIAMfflDJuB5Aqs
Je5Pu4gq/vWLJ5VTyrMX7Vdbr/u/+YUDI0SpFS70v/v2hp2JwA3hFMjuUe77hcFp
ThKEIwjK9RELCL0bvv2hl4fktoJ+xiKNJGMIYeBFatdv6XxtDTU1rvwZaw9ap1qj
pfopHyouO7zRm8HJKZzzrc68tGfxV8SGz1rSyIEpOOO7yH6qupqGj5engOq61p7N
+NmzAks+xu/t37K+EGgxS2UcsBpAeg9yTc7Uv7mw3t20zKTLjUPjlDYP04dzrjIq
VQ+kqX0SB6YRQcctVuQl4bgPRI2g4FUKeguvmU50SeKyWiDXUx4DlnPe6MXZks6W
LziILVZMuYyFZcoPhP3uJb9nykwSXbDWyevoQCXBd7J6968TCHsQJnZv9H3XPzUn
cj9/7E6xlRCELDifvSfcWI7zBLOeejbGstHtvLODvg8LlT8YXABkUJQ2KK/T1CFS
2IOBZbcGH6kWV3XIOeDhrFmyyoqbBugzuYw0w5nXeRkYCmECdklqhZNiLw0rP8LM
83Xb3BW/oY4Dne9LBcsR+iHfogA/rnxtE2wTS6GNl3vwJdw8SZhiDxs29VU01WNi
BT8TzuEyFOsZAN6vIS6OQGogsa1Hnut3BuexARwlTHSM4Rhag/1TWKoIpPWUBP41
uqegNktAZZBrfydaMYxRw5r+TCCVst5drhVi/fNefQSuzlEySSykWyXnjhPtccTZ
W6saYnJCzDFGKX/4gJJ26W4926CDVw4qwfwg1/Sa4BDn+DvPRq8Q5v9SPhIwsgaI
NOwbmJnk5V8ckuchhab3y5CwszykS6Lv4Kj0AaLTlyg4ae0Swya/i0SiuM/x52pi
H4s3thtsjD5WP/XnpexjMkmVP64BeO+pqy/CA79/oW61Vf9TIjDEuT7uR+7KZkpc
pS2AAZVK0FlD86/fGWXqgUmyWm6NsWitZEK9ahqdd5fcuWf+9mmzitZe63bK8i0Z
gEA0z/ubzUX3+8Vm/Am3QmcN4ZM+mgYvojk56FA2+lyzqEyjgBZdHJVHMpxrtcuZ
4BhIV2SfkaOfen3HvFx3bGTt1Oix5nq3xTlVKcI/FQsVDcb+1r+Wx1AOuRj/CCKm
xsLzaWeJwredpxHma2IyV8MzvuqA55kH68EahRxv00eZonRTKKREJsHnU4Ru80JK
5g1tryzX6ucOKrEVHVXhFaBMlsXy+mUM9nS4c90aqR3h1a6NmBT8fx8sNa43hJX8
yVhJ4EBnv8RzT1QIYa33+bhf7ZGiTBWTL5caEG/Mer24hk58htlnrFM85TKUZSx7
E0AxNk9jOyAll4AYRhTxcBS/8qBq+H6PkflQS/I++Z4dtBtFer/1EVsVsogk4Uk7
82jKjZXuaMsPyGjUVXWXJCi02k8P5DgNpGMjW0g+Ot0H/vy9Hx7giIo+zp5kwhCa
yV55l6ylmDQ5yX7Ve5Hx70NXD+XEbWA9x0mTOtGr7yKm8PfEpqip2iUf+/8XV5MF
JwB1YzQCUA51jAOdxyrMTZLTs3ilXoqC+o3p9Jq7mTXXjXnOkXPfk4gpSQGrM2vM
SzQoVlvnB+3WWe3KJb/3ZQejlt1DBy02pLS+jtLYO+UgsaBe75gxDs+4bWOiy5jV
XbR9dKQiqDZF5C3XG6dY2ixN3BtQFzbHxgsWAgv2jMM0Qpzt/hjjUVAln+769GeM
8nm6Blc5NtOGhG6/uVyCQn+cocIRyB+8sQKNlpiFnMTSlRJAT2buhRhT4Pag6JRO
frfwh3JjvxXpph0KZDT3lP7WgLq/Zwbb7DLlYU6OMR3RzGk1M7g1tvqwrq5dltAl
MaHv7RfBqZnimGUG23sxM7fU1cWTq7RKZzcTTnctJl1/MGsKQT7bVkycfYIqFFVi
W2hjfj5I008UV1j44ZEmNz1/EtGLtdchpos9RCE3XK2H6pfIOIbGwfSyfDagnkM5
CUatPNy0ljTIX49+HbCVL4u34RMSrZdr7Zl/8B8WR6gpFqbnTa5wKl4+eoa3S8IB
tyjtaMh4pvqaA9JtVRQ2kIOOFLkpvNOxjXJzjJcXiOf3Xw1VVbP+F8ozHMOnmee4
sLmZ1Dw64hLnmxYrvtfigkXITN0BC5Wimd3TBLHZXo+sUBsyolc5Ay9g4S3OBVAs
GRkZtgAGI1iBSLMa3pokQJlrTJzUHyv1TS73KZse4YzLyd4j/43RBJV7WR0/Joz5
IcbvbVS2un9fspGWStesUOpRdmvnmeoogJQ1yD5juPSGLXBGsv4f91fZwvFl0pDx
5/fOCGu09gL8ZKfPUC4m3AtnjMAsFy7cN0/wWqrVRUuxnpnM8husb049EplPTYmg
nvTTxuApcK6GJyeEAIwbQXuEzMhGMV4bE2AY/QmxisiiQEPlUQMtOREE1/uCsza8
zax8jgawUKNOpB5A3USRgOUz1B5Ov6rxwoxgYDVRsrDt//l9Zhnyzsvv5sricm+H
ljN680R8N511erq+pdrIIJuEE7OjNUgzHw3rLY1lrn9YPvhyPFiDojHioD6jiTRW
asm0nrvq5mUOedbMeSLaPGI4SELxhDVaRbTmw3KytRe8N1QtWE+DfL0CXr8A0/e0
E72Dbm09bTn3mpTfi5rlucjFmr9CO1IRaoRB7+wPevPgrD0i4a3fM7lQl/SlSXvw
xZikCdNnCQjE/4rf5+ap4Vz+/gYJjvQW1z5bfNDUSzu+rfpQcrGqRHtBS/oh0LyY
3GjDrP0sryu8wdifPTXR0u9S4Avd44izny6cF2JTkHCsBDB0jMlbL0fDajtHN+Gi
ASVvf+Dqt2LMnX5ZxoUBcgp+/hPMOUUqLfLSsWln9ZijObydvS0B1r7Kje/u/jLT
8KWus7cbmzWWDbrjvXuXg/gwV1g8D2zTnvxzM6oUYpGTUx+DmL1yz2YwQdWsUtwd
jZ5BtHNu91oVGKQl4iriGVVbBhpbThm+gS5x4brRZhWBwFAl5y12tckNYP7/c0P+
`pragma protect end_protected
