// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 13:57:49 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
mOE+esmBDSwzU0aKeqt3TcxwNnl99X1Ka2qGH6c3BIECdm/apRy9yLoO0fvaiuKv
EhLo2j1/KvrrYwM8Mgcg+SNfXobmIYUUbpR6ijfh8twJq8fJk+ROgGAKsX2VOkZg
N1d2uW+B7QfdQwwskISyI/xv1fpi8YSkB5VIc5E5rTA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3296)
8/aXjThHvTpA0RnNOrl9p924fWxXpeBPIuJki2oUFvG7Jh09XD4X2s8nuOFIdUQE
YmXK6BZMBZ5SyvRflGchd2plab+zhlFRAkf8+ldGq5HxxGV9n5YZtXzys4Wn+jUA
4iLFuLrlzIn6CdoV8MjAfMgCEy+1Y8xZe+J/41HWvkgZ7ISmAtFp2SG7PORWCinL
baWEWBjQGrDZ8jderknEXWDQQ61je0C66rtc/reJuJ0ZcgzDYrWx/1Ztdav0QAxD
hhVz8iUlvlk+JNez8T0sKeI7d7DiPexvPBbhrTAglq2EZ/Z/dmAAawGGYfIGQ9ZE
12HiiOGQ6tR15ry33H3WQNG0h9kMy1W39NUSlEgUpF+X5Y/VI3md7DsX55yal4Pm
8J4owI3knJuKnZR4IHCkiwMjPwNJPNAUnTUSMiJwhwtHUy16pB8PsYT7Rq/ED/8L
nXwCS1sO2NUsn2TDNE3gezGsidM2v1629R69SKEcAHYztkZVcsMQgGlF7ZiDFzaH
/tF4tjC9muItmVzowBbAkiOAqOuFixF3Jq2pQN7jLk1wEABUFi45wbOifau5A9R+
1dmSDkksLEDjp90Xf910VGJSwSvJxk+6oi//Bn2bMnj3N/sfwmT2I1SvYeInO9Vx
DEF1Ev95hOnIM4TEKU/xFQyLOjEkLUQlttLH/7p0bDYAIJmZMFEgn5lgj37zOlnL
8kWMAtAt+MmQk16bLZe4T8MWcDp9RkOyjgsCuM+PgmkZOovOAAAfsouBTPKuJRdX
QaWMA825G19d+9ZfBnrowN5wxYml9rgM09FA9eZtNXMfy92hviNmX4SCV77fLujT
AljAl3QWjeLKmireL2xwBocmw9dLjGQ8c+YhJt2WxFmP76KEaYwIXDTds7U0cp9Z
pFkrgdKWpG2AyN5PvXZTLhCVKFg1DwZM3pt0gfLeCUIZTOmDimP9NWfQe24hIFOc
mWlGpM0XhzyA4zrXfxwY6JUouiElrYAtIrxZ9Dg2wgvXlTGQwJN/0Utnh5vstMbt
Ir1UPt8vd3Pa7JT+mfV3NEudPR3fSAEWzz5VYzZ6p843313t+4GMWYRYM4vMDCB0
ufpRKBNFvdRA14lX8nlt1hpKXHxSecQI46oD6QYzZNxhYtVw7bLMLJdsHmfVKGcV
GADLLV0iLVszENIf5/AplCEP4SLQm2c9OvdljoEv8j12KoRqq9jAd5iOyACLSA6d
S7LwtPCxJnkQJsM+Gczh0veA9a0f/0bCwtM/3/gA8J3AOZWo/qk1CAySccfeN7lh
nC0iANkWJZn7XSxilC3OYzRsVRH/gk7rCLWcHX+7ecaQflp9qMiTKVUluSVt82t0
Ty0YOX0IJsIvdqwa5EMIpy5OXqPtV75zngUneKMAOBPbRDE+6S80RWyNBRuOF5AM
nUu491wPz6uHEVM9zxHfsEAo9njzJcVgq/kNlXUTXARvR6XBGEJfRApKE3Ke3mTn
T4OQ/kHLhvn0LvGSTYVG5f8YUmwZZOPkLrqa2MbqXLadU34zGNUATUgE/jN+LNV/
oDUy6MBkuVzIw6wmk2h2cg0qnVvTfmCnxW1TDTEZOpgSdZv86qRFPHAUlRubngRi
gPYmD/xHOh7aWlsR9ZCTlcLZrx9HcJxROFVTT4XBfrKyJiNuY9X+iWkS5f++Vj64
BYeXT/aGfKzbZxA2i2puUdId/JwxLT1N4yj01Wvno4R+DaOUDV+HB2exPCKEY4l0
pob6TY1aQoOQ1RpFkWx4zfAVU4xuWiAjHIYtj7tvhShcwJahYtExtluS/E91jHgy
nmeqXLGRpZLs8lULQ6/+oMCV2J/xHqe1p+PjUpSWxXFV+wbQHktfZYgK72dj/2ul
cilUnjIAcDR2d/kO1Oi1w0Lct93gZoWsgfgKdkLpMCe3ertC2JDQ7cYx0p9mHVbS
ODeogbXze60i97Ljo5esriQ351Yj6/V58osKMKiwTVHYj6OdNvJpY9NWzjiZ20E2
yp24Jpf5VAfGG0CuTo92FxHn2cMqYCB7dSCt0hmrd2JxfhaTLxjjYNQZeYsIgTYz
jNUNcX8ccUrUVZCC+xfZQ8IwpxGEtIdZ24RC51PXhvnlPPYRJ7ZZxSAQB+tMmk0B
BjPC0U1uBg/z1AJFgjpwmXidwCe+As4KFmN6VMjwP9Zbu938za7k5wux836q/P0a
VOr6LeIlchxsP+wejqJcnhYBxDjPkHi2hoIsGYoQhCtPlXBaRjxRWh7blgiy7Jd2
OpUiIXDATmV/tgN3FkpEaxZT0iGC5M/BZh/EQIYIADUvAc+aIZKVSwaKy3GMhhzC
Sk6cYhv6Z5aG482NT5AixReUA6xc7GsM+Wq2IRT+ZmHX0pUh5fNZrrHA6q7y+Ru8
MEIVM27X9fOIeDZmBTvmuQOvje7TzPPU5re1+G/sYWA9+l0bgUnyPs3kDrUQOAok
opHJbppODJfmE0Urw0Bb2FpUruObaawyRGoJQaUIDMz2dlve1C2Rg54vu8N5YAFC
iSMBARA6TLC65nIRHJCO5Z9GHjos3863gsPpCZUgdsP4p/u6LIyi2q9M6h3+iHkJ
772KSRxoAGIAg5ZqsJAvc6mWH0m54SSMbfCFjvjyGpXLaZr1kFh+6aWUwQSticTh
y2FrM0l2UEGmo/BDB3OIX80M+eW/G+/Jw9gT5s/4CIXeQxjJwe2KzV/XpbWfw02X
uQYko04vFIj20u9bsGuJmCbTyMYlBjPlQ/LAbpalIaP/LuSR3L0Tp9A3MxzDbUDP
xUuMc/P2FzfqHt/Xr4coqR40wo5qerWRyn4FhGCj+ey4EORKBnNuO47OiWt0yEDN
eRh1pfXrC9aftGoV8R6YGmV+lcDVgpd30wR3UDQVi7Z8ha5Ok3ue5deW5ekqb/1t
lwI+e9tLjQBEKS61jPQwhp96h/y4czW5l28I+cBwjAQKo0x7tJoMUICD1WCiC0fZ
MjEJw0m3MIwIx3ps0PVaa4MajJdyRDvI5SnX56WPxcMLoX2DQgnq0I16kksteGB6
lnahNSXgAz3qzayfpJQzE8U2ka7ZiRutp3taBSjFaExvm7N3zXIOI136JcLBdaGJ
lrs7fgOo1hyiDhawa0jW8GjxELvwAbXokmjei9YIM6JuYIMUXnIVNNZ+mlR1tRel
V0eMrV0bifWkpABxL4rvOaMQOixrILQQJxJaVEzQ/aIicfbQlst5qR/I6qvMp/pa
FzPLi8t1BDGgG74+FFqrUy5As51Cu7mk/w0RipBCqFzuj1c+uyxVQCvd2M+RRoMq
67Q5mWB7AsQu9dYM54ofzWE0OEr7544PaLe8+jzLwU9UeCVdRfn6IJSRx5WlSU0u
Ak3zEEmtLdFfbgXlKwoekj/p/aekh7br6g8knP3PbsioecWg+UuGvK3Gb4vo2/eL
lyJuFBewD4+jVu0jf95wBIQIbV1hg51amSYidIy8TyIxS73iJ+4BpWwWdAlKeFIq
z0axtK9uWIoiIyJ/6EBecDnYiFeOoA/d4D51emBpd+ElbJJ3lfpYC8+l5NfH8SsP
RbPJS+5TqtLmSfp356rHygVObqG/iT1SjjhmZUt4poExC0eXhMSiBoqR9Qkv/XvR
3RRWjscOE1zhUAjyCTVKSTS16YvKoZwWi+50b916FCiaFbnNMLvZ+x4iyw0a8OnA
CxR8Oi0icmp3vpX7Cth/jNGq9pDizlzqIRXoISCJPd4JYmXKUjs3SQ5W7k6Zlit8
p0Qd2kHlT5Pp+0rUuQoajbm6vddouv0hXy63ZsOGrlSFt31Ye31+fTvgzP2TDGEx
Gc61yc64ge7AY6pS7XD2PJGZ59w/z5hBBMOhbDbKDLIsB7QXG/Cnat3kfuvB45ZX
90TSaqaWdbJmD8w6dHBTKo8vTJohl0IDvJK+/ToqjIUVpFb5x/mm2nIempej5I9q
CYd8yXxCXF2rxepJJy/A7L3oPRXy6+rRJWuPlzxnq4I1WrG7vZrD9Y/GcTEKA+NA
6VnIZJjHmwZUw9tbdshPaIhy/dxP8PqdfXsRtghwldDJ9qbzEbwOTZbKwvsy6t+I
bIcOtLWgKAxew+wsFMC0KtJPuaMo3SRh+WHrWRqATvEzVzrfBegTnk+DFl+siqUw
8wdPpNE6XxfvbHA2spSlwzR9FAtEnkV2kG0Q/EA1WC159exUahT7VMWh2NVGB3MB
eIgTl4+VB7W2rCRlCmxdUlrEXX1Ku5EuLeEsp3yNOmMkufVAOfPL+gbMqJ3kHDIF
La76YprAMnxW8h966ixC774WbE9Dm2Z9Ic9XCI0o/2S/ln2Du68HZ3QFp4vSREse
2mz0Cg4xHro1rwWcFfXxZd5/AcF2qRsBeexfv5jh2WLfkRNHLqp9mNyfhzk8R5oJ
o2MiLNEp0Y5g7/wFMlr5+SYzVMzKqesEdPwMUU077so=
`pragma protect end_protected
