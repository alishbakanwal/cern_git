// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:05:38 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
SKWDyao0WbTSPYXAqrHGSOs+bYFVVn6e7Jt2v+jYuJaOSXMo4qbIkKfP5SCinH0m
TmiyH/V3Uh0IVk6o0McUnp6JQe2eBlAc009MrqBx3noZz+XxUz3sBJfAHXKRsUix
TOkrKa9E4QsrQVz3RFKevtY0zLV0viS3znnn+nes+Iw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 10480)
xXelVpir8WsSW31nXuLVbd8ryTxlQUaxYuBjeSwRHbMo7p/CtL4S4mFnXKO/F9wO
qXaz2osYt6iDMbi9YMQt6XQsd6HQbuby8VOLbjQtCQclIuoqIikyRVCC9AzhjhEV
fGyO8/1VXSiKh+QUJHhg354QnToCNG20Y0G6FfDGU+AUXh2GWZLohONwlbr+AXC3
bMXM9N0rn1NXIdTqiyrvQJ7TTFywMhzsD67FAXxezuWtoXkUWSlvD5taFNa3/qD7
i35upBvfeuBzg6StGFnt9hm83Lq2JcKoEhUuoFunhaP9U6uxHGRXEkt0VbZ0PUKB
waxeTtp3LCJDsbR2jk2feagCUKTnlkJN95z884tMk38os1BxxhPLFKHOcGHXNT3n
PQV1EE/OXgvTUBu+PEAXz/fxq0MWd+3jYvvgtSwI5pq03IYxrXbWhCOpYfyHanuJ
RFownW4juPEOei9axOLxbdrmmglucysxTiu1UqxzH4j8vVFJrTTsBsQNBpB3qmoc
/bXPoGlg0hvcVBeWkRtgjdcU0tPJtEQx8YkepjzoLrCWF1zhjGmqoae9MKYf7Bt6
vjpSE0wLeli1Yv2ZGkD6TS9vHWplkqualEWWAqzMACbJg0wB1lT5frzQxl3u1eSR
9RMfMwmtqtLavOgJidvNN5JtPE8m0mX2HGGPjANUSW85/siPTJpIK0UmP7nEiSZE
HgAvqcxXPoHHa/8tq3qqqAKXzxfdDGnbvouiCHkH+T4hmI/83FROmrrHcaGDKC5K
8fOH2okXD35sptqbRhsKemAaYdl6RuhutEU6ZArnCcUZxvPS0qq0a2hrrVUguW7N
waowPLZBHJ3vLln19PRqnKV1CuN157hZY7zYnGyO33ob0x4b9UlbgiLFtY7zs4mK
eeG5uxlOAOusNUgUeaBFDbQg+m2v8DuDe5omCeFvUNuMPV17X+9+/WfoEH27FD7B
Q03RsRQ48kCsb9OpoTZmd4bxOJ2yNU6j1uJpzYubRcwrp2Xpoh9+S02Wa3mAmIyr
tDgzWGtjXevKtE4NlyUZ0O6qibHCYbzsNWpPkvPl+rNLNzcbRUAf4baSEHb50DuM
BfjVsDenWMjKlybtvWvDc2qNwEdYuA5Z3pLi/flBpR17Ixn8zwFG53p4pQe6zl7Z
CL2fM7YibKJAIfXKZC/XlAXX3AXuOK1uqEyu3vQACoqgJ5OEDri10VFGQ5VXKsqG
3Gi7bMbgx5msE/DOSNwPcEm9cCXl3iQCfriPPwKCtReUHvNPbSPC70X1vYEyQ8sD
jfplHkJs5AlzMZW/T/WfpQNoLtNDoQ0/GTZNeeG8qiobTVHP6gCCrfxaFpR5p6MA
51jEJUXCEh134A4eIY5hLi40rh4/hne6Dcdw+dH/B2J5f2gUr/RZgICMS3j8OGir
w79e8fDUhvbM7k5PuJVAI7X/S4OS9XyWjMXv5RW4Myyc/Eu9SIfsPoaJmYoRdaRe
ujEpR/O7zUxCaT2h+mG0xDKxQnptBsvXewuk2veotr7rZ999GVyDYmzdePfZR4Ia
tDJtwa4tX+peHE6P5tXIlLFQR0QI66lbRrBCSwd9VoCT7MeTleIc5FUP6QnwgrmU
zCfgBr4v5G27phDzP2LNtb6KzcNgdFUxjDA3gCBCFERbPTRDydb01ndY7Fgv2WMe
ik2+VvFiZXhS+vMX8ppBfzokJbcEcOWpXoDEaBz8hBWhdUjofFCpZ/Ya/FAfaQMU
VvCNwVRHPWPIHCjtYQhWB0fCyGpA0wT6IUQGnvmk+j9a9lB4YG5yYR3JRhH2gXu2
GM3vvrhZsHlTcBE9hd/3ptI8oBVyXL0RPcHYGWLxlywJgfRrWFhtk2NTsFYuKOrM
FVYgRq6Q1vNyKN8tYTs79VtMDIdBvvw4JWtfyQ2AwBzvaTNa3leZezt3YrhYYQaU
5K8WByODgxenJkbi6px9AQNajoHJoes7i3U6XWG6WTAKx+7KqbpLg378GCalDBre
OpSSG4tETPPu7xU7d6b+potvbIWTQQO/iwwmUJO1yj06IchjXjQ9DouoFourgLaf
Jvep+GLKXSVmoiBR3eTueup2jbA0ty0nDvjh+k7EylQUGtXRRCu5dsQ2LyuuGVNl
JlDQ653BjqyvQ4BqBNpEaM3d0z8xtEnAuHOBYMU3qDkzfYkfZAg16io/xyct2OK2
pzWv5bOyEbrwMJLUJa2gWzQ7Z2X43s4e/j7QK96TveQsx0XR3N6fc7kYE2GaKUU2
FdpIOpnJ4tbhsOn8nG+kHhYt5waJf1lUxtPitLzH/yyIbaK93a/vnuR8FzKgYj1P
TyFO3jb1AkzsTNG8LMSg4Sx2e7ANLlEBfIMGH8io7Or8Euk3xjh6N3s+RQsHPAd5
necdlXCS/qVx9Q8er58Ka0pPt3mbMlpqvFIts2pQhCRIHIzOPFo9aQYSRdBwcc9d
HsuiW++U//mB2+qtfu6YHM/Z6uu6rhxK7eykRy1iZBz+da/tkhDY/EQ7aqZneKPO
BppiB7cF5XMnSrcv2RfW5KuQmUnKLemxKznw3Vq+XNIHy7VZ34Mt26kGqH8CbL83
LSMKWyHVIUSBrJGEkMUjjRrhEhKZJTI4Hu1quTO8s9f/tTRiHsycNFsaK1RUvGUO
FPXOqhHGBBW4HY5alEn7ZU9/d03FpROyPYAtW6HM45Ebs/9piHxgTUSvh4fnmnLw
AyK3Xy99bqS8b7tqF8O8XHf0bCUdjNnw6jjpI9Qe3/2CaFEJOfD4gdD4dZTaXc1V
Tchvx0riJ3gTaJuY49Cn3jGjxTL21UJ8gowxaax60+IIgBaf+aVSagL+W9MhyE90
qFC77l6oiRxhgOd6Gbtnlx93A0Bey6AexBRW02UeaChaFO3kPCRigVNGM7zxUJw6
gtGmUXXdfsIZ97cnP2V7mm29OPNC6oYDNKRqmPbI1VMLX4yPDiAv11ocu1o99n2X
EQQpePLHYxgcKjAF00IUHf3/5TfU/sV09rRPvELkAMu5t8FnQfai495wxrAZc9nf
TRvi1izZ+rHh30MB2ftZFaPaDAdKqIbo/dBajvF4eAQRhvuY5fu/v89wjMQ/fsk3
DNOlYrec1CIzkQtjyXxJQPR2k6m0f068bDW9b/zWSZsyMjGvbTSXeOWkaICs/Ha3
D0vpNk5gl1X1jZp9MtXgi05Z+IvOJQzy+N9Q/6tpPJcWnPmydWhDICCKyf9UPGTH
I0fkXP4efcRScYkovHFjjeP9DYn1ORWcoC7M4Ykc50ChsOz+RIjLWQ1lE+Jx/9eY
9jJ1+FV+CMFXLf7Hof9tgdoL+Bss4h8v3uQCU0n7mli1DuzTDj7sy+hdGMrkMPCz
ekOnC/ff9ikr7vej3iy3rKq1ci19dA2CIkXdVSKwGyxC0yqK6uG89yBvsZp0/vhX
6ZTJHoTZh8cqFOQSESVitTx6NsVv5IBTMcBesUdU1K7dvGCqrtGKfxf6AcgNOUq5
rEuM+uHVVmrUVyWkdP50i4hd5aJV3INo7lF/r4P/Ox7hi6Pxz/BvvKS5e9mYT6xX
gjA9kONpLmhFP1lg/UzMfUa1+NMWC6Q3kuLEB7zAs05MY0HzV9RD3c6NG542XJam
F7iUEtFV2JO+oYActcUOTExhNJZQ2tcuoK4SNzNj/UHVsK1S4fiBPiogiqDKxkfI
w4zTABsMyrJukXduHFUgJUQDDb4LLmotL7y5Q3UsJ/YFheSGDVURPKXg/Q+63TV6
rFjObbCxI35Q87NHsHBlEgFb/1TiHSiGc8OzGn+olsqZDoKWOQ0oCw2PSyn+Obk6
8dQAbNS2v9/GgJaIwzMA8qaFCnatHn+6yt3t3PGZgaNEuk6pnwXQW5KUmUPuhmTI
j/e3hd1Kq98lOQmM1Vy2nS3ORPR2YPFxQJGlttjZZIG3P4eb62n84qLdQLo/0YPf
hlpkXbMdlzEe1TCBuBPRtCU9IK3NQn5ZJBhAMlExOYUZtHTxIf65+DfjySlUjo3I
g8uMzl7h7I7CQrp1KI/W3jSuHCD5tHi0pt/Puu5+4pP/gcPd7Ir1YQQ2y8dDccPt
px45wnxajJxGRAzMoqG9aINvS0gbep5MnfzbntBOmt3OmWLhIyysvDMVhwZxPEB0
sT6xttvoj6DEJZIInaqPJqJlp6WxcNlRLL0ZOJZ4xjyLUvPPsqG/S8+j4jzVODuY
x7I2/EOcosxit/jh9UyjzBbJ/m2TZ4zbI27nQuOCKnh5bfbKNevReG+IKAU49mIo
kVSpeptY2TNRF6U7w2HVctvfDYXIit887BSrX0azpTIPARkEXCD6ROksdng9/7ga
uFR9H6Ea5OZ/7jm6wqw1FgmyAFLINqwHc/AXxYX46s1nNibDeFJvSDE4zpOwC7R5
KjrsTY2epEo8qb5NxJlvAIngzs6Y0mdWFBTOI+97kqj33FxLio+VCVKoXYfzHzok
2vH6C6h3KJzmPtM+9GdbKWc0hWeQYSBk4t8qDZiU/7+IcGetWy1G5gFleLuJKDeO
oMkGsoXGIQ0FlLgSj7ylAJ3PXGdQiM9IwpwOs0RIvjF16He+EwJxw7J+tlkf3D8O
NJrux02mZ5BEzwP3W29PVoDc03dxzwQLTT12Il/UMsdZgJvxvF0p4GrFyrUcba+w
toQKNY8ZknmS3YZ9uZVz7C+g+GqxlAJwJwnSqtlStguk0/tCFopRclwfA3Bx57eV
wlLyKt7EWKD/g8C03kMyR9bJF+SLux3WcVYgZWDdFXaS2fa1ilc8dXi95WfuWx88
VRMx81AS0VLH26FH9NwzoYL1kh/5I1+loG10CNourZWjL7T0R+Uk/kt8+g+0Qux9
O++PZjsp/Af0GwX3/JBONvx/sJY6pPJU6+PalSzxwzezbS9RQPBUBaVLZmOYGiMv
39NaA6+rp4dcg/D5p77VSeYLv2mZsQM7D+5dRzYOjtU+zrB4wPjkqEPyn7kydM5k
O02B8ubkRtUfDMeFpT0uvVIpKgOTa+12MwDhgeje9NDF38jk3rILekAX/uN/gM4l
PUBTWj5DzNYFyQPEzGsilCXAKgKgHHRNVEkpKHprXvDE8evf3p9407xAET1Oyplx
tQ8X7L1ojjOBQMjVC+K10QgJNgt8EVcYoOY0kO9XbqglLS15krnNOGbjpDzT5txN
3Y+NGAvq0yXufM52F6SYYJS+pSyF+QCeWEeIXzJ4KKDwxgVCJKi5IRcWPwFBgyOY
6ST3m1MFugO+mMiH5jesrgPnxIchSBVWMkw+vNO72yRUXbISUdU9s1Z+S0BIt5pa
hc43pNGnq0Rb5dNXQ5tz18s/FiH0aQEGXxfr+wsbHwLBeiTWwFdvrMAsE1KSCnCc
xpQ6JvjcJrGeZMrSNcov7vQ1GAHno0GtCE/9Z/qYdjWVOUMno3LF3hPs6Yu6YDE8
aDkX6eeGjr6jjy6Bu/YxcR/sLcmfSJsuFSnZPbK5N+VksQRyGszeKwbl+/trHBVk
SvAPA4gEtUeJNJJeIIPZl9Kk5UgWbnJU6OmgBAfFU78V8emM0rEGhMkpG/XA9z1B
TBslbcDH/P8TdB5UkakEacUx6HYlISrH6jEY2ZeA2yM+P+nt6s/gOH5qYaHyj+4T
I/8sAgs4M69zsh0WZ7J/DKv+Lcky7rBMC1gr5GGf4DOHgH6CdLElUAtsCVdtlLz2
//S4LDwiie84bex0i/L2ruvAZfkBlpvXowkaksikS9XyL0RCrta9UzIzoQ9OzcdI
HqILxknLluJZN/A7MSkIrxneK6OYpfuxLbuqIU2Clvb6J9L/N9oLYvYQJPL0YKEA
zcvCFP7hLvTyzQo95b+9ShEmSj1WlKlN3FZn2t5v1PkmTh91qwLiz/itkjwmG8Za
80AztCItHWpjZ+0tfb5r09YWGOKW3/eRDVRJDf8dx5HFOpuLoSeLytOQ/RdwZrBz
De8xmlCTDswBc7PK/5kfEsUmST0QfCYE4Z8Oslc92Hk2Kk4xkWRj+fBg5D16mpyv
3PDhqFa/uEhlxh62XOTdaHq0TgzlAmZ1tYKXDx3dplNJrQbBs3O2h5+F4osV5Aoi
s76EdZudt0g2V8nXPVU55rrnn8lY71US58y42NCcrsMjFQyhT6DZDyvvuPpMT5Gu
8tDeDE0hjPBlsxd6/klyCpe+ltK+UGqLMbeH1QNMEcqcsHSfHBBDFZZv9ZrqKLqj
vYZbc3kt3NLP+zBNZN78kUzaOwWP87N82LEq2vadxHhAc1K2JhArjBZC5GB9wCk4
/qKZ+rN2L6FwJRgSUps98edgbgM0vwWXZpD6A9RDhcF0AGw4itIdH7fdvpcobvM/
uFYB5v3UrcxoboOxXaojUcx5tTAMI+RLSXMxShaxB+uHMSZ7y3NyLM5WVF1JDhQt
pLTpeXubMU59b5Xz05YOY5lGb6kjEHDEqW4TwnyhxLbXKVktABFKd3q1lZo7ftot
CH3uCxZRF+oC/dgos1HIt7rvSd+d+qglc5C0S/rT4ja0pdR4SwYp6DV+luYA4d0V
cR17g9FwLw9GPIqNgNC8ceDcHR/O66ooErE04gI/CfLBjbqS53V5A9LaiWAs/J/7
CcfAn3lp4qHZ8c3ZocKcTFcX2etsZKb8CafOWlGOSScKT6/dinz2s3Z2cU80Ly4k
7HRk5WiQEHO1QYBHYgcFDdetu5FAhkHWb0HciIK+0ToWx7w+Eoka7GYQIrTU/9ZZ
AAQsRF69gdUFBMqSwd3A0ESaCvqwjtjRHRxRKX4vsP1kHGPk/ISP2fd2iJEUwQN5
k82G6GDZVOuQBL7BpU2n5+zTlqWVkyFqNbH0sawk8CxLF8qcrj85tuM9kAQn2Ict
HNtCENcFKRSsIufTpksUze9SXj3Sf9VzRDsbTLQMRDzzJaQhE6ycWaDoMatDgPI2
C6tg5pF4r4APYuZgUCQwMqUqx9Pq2LkSV+N0dAWnq+VBk6Fw+cc5+2gP4yGkvx1T
WYFchBc6B63w4u20E68Ij6T6SxU1WV0anyKhp9FoTnay7SHWkmmXjd1iiskWTWsC
1wdDFDMdwgcrPjVrZNOmaG6reX6JnP6lib+4Hn9zhpLsTuKWXBWGse/Uay+1mDA8
fh5ShzgFZI/dldsRCsJhZXpqFyk3VFIk/s3ft5spB+kIKeX83+j2dJpKXY1bdC7d
jfJqoV9pyzq6FnzF0mXD1vWuCaLO7j6wYcJqTKg3kK9b7L9giWzOT2s53tBijFg5
EmVNiyd563GGMLcbjn4QivaLilqfsssf4Siq40grNObZyAdFWp2VT2BcfSGAVX8D
MYo09akgO3C++i0wEQl4AUp7ms01SBxgLV+8cREZfGL6g/WAK0mJs6mFO4izF8T2
Kkr5l0aK/xyoISC7Bj0GPtg/xz+W6d+G6/fYpKpnPOL8rzTgN7I6890USGgw8X69
BXmxbGniabVUWQiOACQrRgPx1FrxwnoqeYfHHyjh2NLqLMNVii0YKeqDduzUaxXb
GHtrjDJaDvqHL6UsgdJJnlNV8Bb4EJX2IAI8cnUngilqrkEePDrIhJbhLeRJgQmX
nTsa2BWCtImvcJrWEOMnLs1p0JIyHLjnzJN+bTRDlvwD2UAt/8mtC/5exiZKmy7z
eguPo9PV0FBUFIOEyWzBarobAlmlKJTa2wtYm5ruBt6BgSpLNt+9Kg96/q69NL04
gPeTjlaDgHVPoulhvzD7yv45WeP28y+HLAJcjQkBoH9RIgK9ipOUgA9TxJVffAVO
EZ6r/DFgL0/k80Kq9Hz0+f1Q3TkxPnHnQ0fdmb33D8seS+uCGsj41sD0buP//2am
BSlI2qMMVwQ7HX0G4xienBP711GOm8sBBL6mynjuyCfsyfAoe7VQHu2tXrW3bg+4
prhDR0Ern0ze/+Y9DdgE2wcbuljGZb9FVGXIqP3LHY5e22UX3kSnF4l5pXsUxbZu
m0/Ghp0zv27TmccI4FCjCgzP9r9F4m9NL+NBt3Abu4QqWDWqN5yj/lUOI5hTGX2B
22bUM2//ffK5T37emPIlhrdWuzpjDZ3QezPFjZx3DMP8N3Kk/MMRYXdexMhCXRP3
3xkxdOpS8Iq1ATo+ErSKLXwVqac7cKJ1dWBQ+Vex4CAeDo5yv86FUnA4+oToyv8E
CIajQODOt5GgxJ7JtSfYGmw0e2zOm0TJKQFwkTveNB7j4sTdvWPmaqkr7rsG+iqd
fNc8BV+Usku/fk7Rf7OXzrBbsOu3ec3iiX+ljwzLi7fECtZJ63yTyGb2/nq91jAQ
sfcubYuoGuitaNclNQ0VNZAyI7QcymGOh3/DF5AHBGZTuEuzzkg+LfPg4oLh4n0+
S5gviMkxVmlKRH+wZXkE3Zvr33CyZJ65qLFRo5ernwMp/Vd4pDdbn/2jJNVK6YNh
fBP6zm5cPkr88EPDBD9xB/tC7hwqjCMtJZiej4Lkt2E7SjbWscmB3HC+UM/MYDf/
LoxN6H16Yc2YVdqdYxjtqUDyqWDVeNNv1hJScQfsFss+r1YUEHcgxLTe2dgJ8p8G
/qlcaz8FNNtMCMZVFhxolFw499s595Os7Zh04Sa3mm3M3oxoGkznYkgmnDGYvE6S
h6mXTP1tK3zEbPrwQGlP3mjwpA+JXVU1ZKGoRfvhl6sAqscoaadp4h8yDMfp2JVR
C4KvUm5z3VKpUdrR5pj+awU7P5WTVZ6pYLpCU2ZEqbOT3YG19YGWx03vuTYpgXhO
njzFwI9bxxSEjpV6wn6JJAEwbGBg6uNgGgD6PEnw+4vH2o73oTIEuXzYhOpprWYg
1+ZsYDmWehyRFMk+usGCbN55Oafn055Ue8kzNuHGMDjSyJDeRHL3+vLSGWNA2XOi
avOOCapZyTiJ1x9jsNlvxzvenJKvX9D/shNnZ6SW9cBZFXPs/2Jzsl3FjN1X9LSP
sYnMADqsBtLAquhvMeTt0jpJkiB1iC1Ik9c4R0t9m0hcGI51scQN9a4m3UOXAbHr
D1KGFUY/cm67msYXtLvKqXEKC+jJjCMMX5y/hrMr4L3pb9JWvqLDfrDQMBwgOZJ0
q4TGS50U5Kw4vd17f6JW8Lfz+vyfmmCUqIuQazfyYXdjvLHh8aRvtGInAMFL8tFl
KqFb+/qpzjaIk/9CVC108cIw1bfp8v4aMsEU/S3LO4Dgz3Th4uON9gcaUTxBxrUh
c5MfQO2T3BSxXPZH2EbGjn/GkK3UMPr9UaucVTIE8c+I8xaPqVYjMxT+FnMm33Ip
B9oG54jum8Uvq+D+i84ZiutlpdNnKXU+SywnLb2rZUzrUsKR1qGb2aVlE7JwkZ9W
tspQ+jn4U3iT0+9u16OMHL3PnKl9dAqyHti2G5SQJBNC75HJzgaUN1Iu3hF1JkVY
OOQbJs8IwLPL+VH81uOXG3J85/5xjtHZd21WpKvyiaD52PjHQzwvs5NmPgTQFZEn
vfh3JrE43GHm+ATehtdssdlRAR978DoV9TN1sjmY7zlAMBsdIUbCPAKi7CI90XIk
J5zmIP9Wi4nBvfO4A06ThpqO7HKNuGfFeDWSzvA4LAkpueYzOfwMJxEtcARgmQjd
2SRjp6T1KsaAYQfyg4U/sepWD6xpTg3EdPqHQ+LULFO2mUyW3rGzXeQeeHTVFzCh
Hif+/nDe0Ql63By5aiHxnXVYm4r+cGd+oXuee9PQq+j+rbO2t+u1BDoiOx7S7eFk
fFnOnB+krj1qXVDswCWmuoim6RVEqu1pfW6LQZcEDeIjKu0Yv8Evb2NleKihS2lt
NQIYw9nsg4ojSbs83sYg6qO6tZ3yK3eHId/2Wg+CoZtN89r2cxYOplvD1Vp9VtmF
cqWCTHAoRXwP63kUAaM4NM0R0+aTfxZzmWpSjJ7HkLqDhMNOvFfNQdVcELA4AeaG
/Ri63WkzGgU28ZhA2fGv568LfmjPfbKhftGt5gxMASodwPbLA0zjRuE3yXyadnJT
krqqjmaSKRPoxxhbGNmFJlgE2E7YqwGKPVgXAk4gCdCYJ7j52Euz7K8Ck+zWR0+T
u2HXhVb7huhj3YWH0gxr4fiA10Gp8DvCr4RtMdfBpV6aMA4OI4O0gNkgkmGPG+zP
1M6DtHo34+3ht0zxfeMHnhJzYY69nj6RWqVrx77JGzIcbID5efBm8Ew1L9CKPTlg
1U0LfMvK9+/FTucJ0lY61DO3qfsHyraXLHGn3owK113TAfh/r191MSDQ6aSCO4q4
8aTi22F1tqv2OW0B7fDnh5USUNCRfCXVuhV538391ozWg8drpGn43IuSxvKhuJwP
6aAuoZAs+DGv+ZbrtDQWA5Su8N4AIG45lRIG15Ca3PaqnUdenlehnOTJQ/1WPWqt
iNljYc53TH+dIYC9bH1a3rXpTUpXzW9YMPVAvBmf0qGaXb32xPAOEkoiWUPqYxUT
QbLdJEcIZBoULe+MhFSmlK5TcgnIbLc76l4GO+GtAtD86bVrU8dTuGzlJhKyN7gn
gCnY9RePhWbW75osYZn+fBWNVEJm+GdMI+lgvc4xiAan+atuV6JAz79Edh8/ZJhp
kRNMEgqEL5PB4N3ePasKZ4AcXvY2DrxUs5fdHoXJhkQotkewYkfUFmqYikECpX7/
5fqoQY3sQsv5aQ+euL3SknV8+qx4MrtXmqq2dL0zLKjS3oAhP+bhCWonhej2p/CH
mmraqV9SKMD0Rvcz2XU+bkQBJqgWE7TBq139yxyC6DJPuDA91y0MS05kkommNjVK
/LNQiCtg0iT0bz3nScRL7Z2hYCg/q1Vq2OSiusqcUKXJYTE2evt/5OP6S6FFZKhy
lmW3AKNwr3V69dp1rnEBZhHjNx0sAUlFO/mxYd0Wtqa0gGGvZoio4r+Yb7fQATXw
OJYVfv68aG5rejYBHgbxfF1YT07i2Vuo3qwxLJRdcnHJ7Hwy674V3Dpby00TA3jL
XjbpcUH10hNCJu3DFee1Dbf9BUjsBaWQQIB70SWO+DMLbJe2RQrparhxgPapOJWg
Q9SO/jDNqJZ8kmuQWllojl/3aIlfSQqihQd8lspo3ti+xQiWQ3SdM0Rk6lqx/m1a
TXJV0q8Z3PQZfXHwi5/VdQk73YCN4YfQKuA11bM1LPokBkL6xdpxRfiJArDViWyY
ze9ifWbSeGF4sQf+EeyanxER00EUd8hsFUsrtuYXL3wqBGUezizNv+Nmkwwozq30
yND+M/MAAI7AxEnZElkfmlbS80Let1DYiQTHNQhv1CBSFm4WBEz/ZsemGsqBHMUE
Eiq6EYhrJnccBMGq48AGdssj2evme5kLYWVtFydCYiK5I8/Lwpmg6Yu3ecMtCs8Q
8XCxdYlmBWzrsoeEKD6GETHXLHgc3c/4yHJ58WBcb2Uud2b34Wrr0fOCeQyEd6F3
gd5KEQNzxpEfFll7BIGkGO+iD1tgCThC1Awef0mSl14fqlW///AczPCCzV9NuBo0
Qw3weSzibROhLBi27VaPLq+p7xDWcyc+o95k9I55Jv55c1XBlrkY2Bs8hWgrQULH
0/Gw9+VRSmk5nb7K07LdfpjccF30Y4+L3QKgnOdqvE/NgXzeyGJinHAFc94eh5zu
6OzBbktWJ0Uo9uOyQLXfazIyAZgljg543hwADlwnLsP4HH8xKvOw49+Q1bp/8B4l
hqqJ3NZtYs7apfkka8CPVkc6pg9kpH6V5GH2O3V5ksRppaT/bY57cKpOS9JGigLR
vUZ0BlK9PAJkOkY0XaXwL9zY0QchJ/Q83YhlBPWMyTR/OhvvpOjoZqmAHuXE6QR8
XvlxjkjZSBFmQW0t2La9+E7rgsrDmUiKdrP1Mn0K2z7ftaRe+P0tleVqhosVt3B9
6NakQLKoW0QeVEsf1SYJgmE4aPfozydJiu0OIZfwYlnd3WSzUCZKWiIt/l5uU9iO
LBFtxN/IrozkA9bjpmEIRfG2J6z358REntEVdkOKAKjU1kwZrQaw1u66tZQkWYdE
AdXFz35QRXipVTk1ybquQJ7l9ptFweZJWQsniWA+MrpN0vE+JzP4o+D5amJTq0bO
V81R0mKDbW92aPSa+zD3Gh5phnB59SD/ODu4nI1Zq6zNXdrRHw1rOEZnf9N+DypL
c5h59pQT/do0OEjqLCzmjRy7zsdA+RUGjkyJw/LMZfOWd7MVHQ8gM0LBy499r3rX
rsAZm5ax3oO2ZJajx6WuggFQ1HchCl7OBQFOekMoe5Su2AtxauOskZg9ATwDlt2Q
cSOxTqhb0XW4zQfg/fMy0JtUIT7V9/2l6c1YM+azf/PR7ycT2JoAb8YAGeAnV57v
3k+NVhxhSWrDn6C8QvYIzjkurjc9BORlDyr8gD8x5Nj20kJLx0PvrhSj2zs5GDvM
EZlMq6I+5RigQqK5HIAdAsYGpR9WHWKnthg0AlPBZ8MoZwMp2gXhkWGGkw/oiLal
rs56NQOX+9OQkC/VWMjZ/3yG+8dpdZYlIV3Ul9DfBH4ORF1FlfrEfEdBElnRkdNu
fv3ntT850hy49cFOG9m/WG1HnmDkBa8gvgi0HwcsLTA93Gx9quEl5L2VL7VixsiB
MIN2ML/gJrz3wecH2+MYp+L2W3xyyf/PfDVsYuynkEn03Qi243YEEUPBwvQwqtYj
KEPW2SQ0fPJpbukKh2ul+pFmJZV8Ujt58JLgVOXKWsYKYTzMBGykPp43TAQ7EgBC
NskNdYBbzFa7pUupsAMo+ggernFvAkizuwWbfxW+/6lHOavSDMikvMWU1rmZ6RK3
RsdIoWolROsafFDK1E6HcoD30AQ3xT3CeLJ/oJsgFJs5i191S7WhiOp16ibXb9JM
8zl6S4LWOd5qyR/8DJizKL2csRgNK8MXayR964yl+cezzGGqwAC4kqyoCs0b98LD
91x58jRda4fhyJIuCqIuaMk+WTqH/7h7aR89Ny37ib3Dtl757OOBr8zh5OSk90sA
TThq8TGy2d5W2VEK7GJl441bwXTk9vKuNR4/ZiZThannPb5kirp8gOJDl8NY0QNT
davAZu+wxtlpM4TJXd/eaXSUUwaXHEk820MbxFroVtE47wgMBkMkHEw+GoIGtYSu
OO+4fenZaBISAsXv+fD0gNj50jEs+P/tsbatxu7xbk2B/Hj/rMicn1u+nxE2yDDx
N/Kq+6u/pppP/uXXYSeH8XoT6VwoqqRCXRnEyGHgnEtTpYif6UJJoBObrM6WkGKS
S3Vvzq8DE4a/aNQvHC6YksW0tGmI2Agx6SH5lx5DK5WZ5yTPHUTMK2Cjwhluokhf
OkdKueog6BPTmO9Gg4IsvnL6mTogu2usRxWCqtti5tiR7FaVKUgaUmbOq6YF0BPJ
qM0MT9+qHoNHraM45WCdb01jUaD7sYDRzKmCnQbECnH19hM/kELBrNBcNIEsHYnB
5ZAgOQ59ZqceC6dRU2cz6rOf/JNTkjdJvXeFFqgoq9vCErNRwDmFUe8Qzb+jkbeg
N5nBivduXBe8cH89SmicgvUEnrJSllzLEwLqRzfVBC27ih5yEHuMUxCFfu5saNTn
mBCglasr/GYWOt4Vq9A4VqPoNoV/POzhbyeKCuylgPQokgy5YbH2+bcPiVe/JQEX
E4D7Sl1iCfHtqqNhsL5MqEzZoFwvHyArF2SSjm8QOyzyLGeznfxvsTtcL70B9gsm
4EYekxWXs21kNTs+hmU5Bs+Qr8wCmNNfVtwlb5p6YISPhwQ0SCBsvFTVSsSeAOln
uLlnyKG7EZwtvvO/jmyMtwWaMFO61TMW87gR4GrNIVlEkMamCwrzCM2Ds+DuUJwH
SkwvMRiumr25Gd+S4+nK+Y3Jm3VAj5Qt5cxVlv+MQn/0JWS/HnmSJKYPdmdppe5W
BAK9OovB0REsCCDPDMkso2rGPpn90nHorUDbPzYey9xH4DjLsUk+5dR/4J4o/Cqi
rs7Puriw8+Bov8FviX+D2HEELAPD+PZq3VV9ybpyseA2XHmsOZGOvPXz9y+v7ela
7vfAJGx2dewgcA17PdXQmnmgfHBmq/mu+KN1lL4EhnVJ6c680ONfjUEHkVfIyX4G
IOkJh+JX6VUdNg8vKu25lonoAEF2tcAF8GuVvjrrupvNDx9rnD0ynszIUxVVzgwL
QijoBySXl0qvEAcFHfs9JQ==
`pragma protect end_protected
