// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 13:57:50 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
D9r80VoJ8ffCzJWqQTrMyfEAh2+rpYIT0n6GOK26I0oeiO9aZkIIgSHk+9xjFsyU
mRnPl4hkuL4og9NhOGHNIceCLv7YQGnSdtrfUIjOjWhSpDSKFSxVRwQ5FiNB1OKs
8hzB3HGS4XPukQlP4Sop0xaVxKgUeO0UG45mu/+H1Bk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 4864)
kjqMQ7wp7rDiPi2vMPyz4XABD0lva/qvWYEIttHsSXTUAEoIu39sAgmwKI/LcxGX
nJyMoSxx7Ww5Y2X6YsrPWnDV5sxEMZMiMCr7ZGZovUfw/SvhfCs2qcZsmmkIs/I7
Jc/yqLsuCjfVxx58oLdkYex+q+cqg6Sw4NFvJdwMsIvtyz3zJTfawciunjOrlNOi
dZNOSJx1oM7PZyENOLDMiReeXcZ719MsjSExdeKi/Y3p7RWy1ssDsqENGeiSQyY/
mZboQJ5Bs6NYhHR7PgGbo0noo2ygEIW088FHArPtIdTm0heAd6ziEzJHt9hxAn06
j7ULtKv3UPXMK2JFZs4HTmKt4FGHfffV81PTJm3gCCD4oG1P7zPqTu0rJ3ksiEOs
fcFYuE4QN6wjfNIi84vjy0ycuNX05U/jfQQnz3YCI+kXB2JL8iJVpKN7YaKv1pY0
QeRZgL48qWBDxciXBqyI99qFvuZWy82BzFUUKMMGmJP8fBUk4Y6USk62y8Z3Zhug
1w+VKdvOUPpuFfN4rkfeIzvE31h2VXtCxETkaKmUoohY1Fqbnv8/lOWUfm8HUkC2
EMfei0Df/2E0k65IHtpZgvtstWGS7qWiviwhRyqemvfjpiAgPLpAmgriw5LurSmG
IngXb65KVSsEOE4sL8gvvRuIP5H4TvRxcOSRVJrXueHHfLfH0zCnzBdMmQyYpRLD
rEFwhlLk9MSVSWQkeBapMWYNS9Kjel2wL/L2wZXuNa4hXUZYAX9vVj0R152g9MOV
EWFXiGcCXWeIxCjx6FOjxcE2Osav/dbWDDOnF01CLJ0iOQlji27d8eimUmii5ZGn
8IiXq+ppc6t1mSaJKcaphy/cIWwpRL/Z4tR14KfKxaNU1slbOUcE+2bDaVA6xdc6
kXk+B2AhAia8XPf7wY1gLTdhcRiPTT4KWhsVw8rXuknbgAhVDhnpQNBSNZdhoY1W
nXT9G5JrHP6eKQEOQDgW9QI5okvBFxND4v6nhXTcpsSVdLoYDy0qwc9NkreVXjVX
884qDYXnbJ1dJe0n5grqvwVaXcT1SllWj+87o4GQ5ki54L7P8HKKGAHEBVm1KY+/
5rztXHVDNKGK4meyMH8Y5mPP3r08xhr+uLQjvwBTAecNNozZK/iRlEHKPVAJ9rAc
DDSbhirLK2GAOlUVT1L/qmbXOpHmeqBEMwBdE1cUxNOg2iCq605OPa0ocfsiiZ29
ZLPK1lwR1uUbjk6HQ+LqKjtPxD1j2inqUroZNVRB3dO9VfvbJS0CcNoO8zVb3w7T
+0yk1yr6w5GXznNHWbL4uqp5Qg9bw4x4duhvWQiMUdGJBE2U0vbx5ArDRJ5IPa3Q
RuBjUCUHvXMm5FuWPiAoLS6S1IIefN4EQ7SC6ml2asrhpMeU4U9aoPyo81CjAGaD
mFheIzVA8d9YYcsVwbuDKZCnP42e2CfJ7CUgv+1c1qK87mLs1N9IiGSWrDwiwPzs
L7wHDT40m8bh2g68KBUwGuZmeFYNv6VA2BEHWKLrtwSCGdS6K2dZ6t8Olz3i0zmY
XnG3Qjbp+hlkS3TW2i2fRaBsEyKW1aVipFINlM1Vsf8pRGAnSnLUuRiqnKKuywRP
RJmkSFinWOAB0LKcjyswVve3FiPI5C+bh8uTKFDEV98MB5aqrTUEXYDoX737YqHe
2sNMcP8fNGkCGlkwxTTvU0e/7tsbXIuuz/tpm6HJyeINHGfaAmGjOO3qvUseQoKu
RM93BGEPwqtgRzKNqkWR6J7BCit+ykso9jZ2szwXQUQ8cylrWC/PqgGYm3eVXO7T
cODJzvpomaKNK5qK9slZWhTHf7Qm9RGowPym64Bx+nCLjvpoB+eBFnLc3l3Xs1iv
kdCBRMhWDn+EITG0JPSfagWwm8zYNu6GZC8DG+K23DhgDzyTfvZO+sprgNv4rAGK
h0ExyYyuxxJqZ0vyu1CPuwE2RBYaSDwtP36jtk/2npS8DeThZ72OoLfdiPOh7Qdr
TufwxUay9rBjVLQcpPIwAZImKwusV7go4qfcXnXq3eRKEgtFGdSM4MBJoPn+wSox
9ZVPqOG2sXRjhDM9ndIH1TK4TpaACsXzJjtk6aK/ns1pHyUVYdCAOGVcjVA9+t1X
odg7d7asss5ImxnxNWCcvzKg+rfdbSDh60D9m6zorilTQ+JBP5rd07fhip6l/hAa
PPrGiJ0lKb1YqjgZmlU9Lt7GJ6Z+vLCekld/bQnTiC5dxC5Vj1pNyGWu+1MeQE6L
ZNYKcxvUA7X6LuIqsRuUFOfkLvoIg+t2wFmvU9nr6c2ZugSq0ChckCr44lotLeDu
Lwm1Nn+y6yFv8/mHtTquasy5ClYNcBckVWCLW1IUwx5WvoKWhWs/W2+me6VUH2n/
lGXXkqG2xCAFg0ZjouADuAJ+lWOQuxg0sIp6iHqzGY9FcIg+xZYo6M3a25di7DA3
hU80s4j/eQGE3yUNwxjM4H7kzJg88auL9ijchZLxFXy+JRsCqyebJBF02WcHgP04
Ed4mziGpeq+zpzi+cj9b1Yrb3cKYmID/ee507CdeA5rM52yRsai7VOjpgkT7mZws
/bY/cdH9p2HRcTIky8oKbpoH3bJO5qdcr7vnB+vgIcb9deVCxp866c4YS1qC86HS
P61NLCdjIALYc5eHf/GE/fHK3EvUgB/rFPlvdWiG/C4ntMT8GDDVll+4wybT5i/p
CdQ976p0nfd1/i0y4PELkiL3EGnarh9oyDKCi2pIEh4Ale/WGx/aDjAlsHL5WUrJ
Hedl6rW2q388WmkOOnJ9BcU6fpuR4ZGrW1BPebYI0Et0wkOi564YOiEw0mCymX9v
t+yCAkG5YIv3/3mutz3iFPMQ9a3fP8dCkMRptjouShoiXKDoh9B1HVegShkkXgWq
CDyZiXtyRRUHnIXK9aBPLLb/hnitUhCLCEJOkrw/74WPUMMpF0whDHVyR14X/er2
4Ls1QH+1TzXUsi8OcPpV9YF/Orw4E+J3t1MRs53/rbx0dQA7aOY623kJeDYJ97Iv
4Pu2gguvLxRwfOqk1p7a7vjSbpwa+izrJdaQLK1y8hymYAubpoX7LBQQismyN36v
b7rFKyE3JdmFWikG/v3V98v//vb7QI2B6s/R1Wj/RXWrBJOvaLrRbRT3xKYFol7+
P7Pd07VVoVf8xUdOgvfus577B4vdeNDYsLcN2kATGr74fixg0Og88GIdwxnjV5by
NfU1HIQ1ovvKGBgnz1gNtzGM51B2KrsB5xw+DpqkfVJnjODiucQw7vp6HVHdEoP6
q/5OG2HtBvTNH580z6CkROKZYeU0UdmyyEsqUHebVrG/+7AtPJ3x03EszIUss85P
ADnV4YWN+WqD1w7H6GAKlsfSQQgF+QXRhoLbAbauCNWq9a+Xh1VLHkfBHhtgMx/V
4KBVlWQPuW5zUScmm0NIZnVMSh4IrJ6NbNvLBxEXY3MvJNC324tVOSHYRBcB8Q96
D773nTPec6Udpi28evB7ahqsea4GU8QMl6tZwsUntUHYcBtbSaKkp8COEv9JK7fe
w8jXs5+3tM6XQyJv3UvrzlxO7HhUyfOLrSG0+rV0MbPTQxP1X9aCiy0Qkl257het
5+ZeP8laol8noGIr+x+eNB7m1xP/5Lx7FadP7uVKuE+hBkBaE8KP6IVXovxcgBqB
3NbBQpc7qptg11WswBKiqiKwo1vzPUNvtg1UVzMijcb9TfSQyFhD743z98+Bd/oM
o4dYYM98nmtyc9A3z6XTRI3sc9VZUj4+dC5SPTpeB4L/Df1UhjlGicmMFMTqE1mf
Q4CNL9vg3uuOkgQGl1v0zkWaPe9yJBUNqjuQ7cV5MiqSaXR2dUc9uAvHW+ATMs/E
j3XLQEHXrJLzW0b0mhFaXovQfUdOYoJ9CGLUGKzqpPjEdMWJv/rJxTIpn5U5MO1J
oI23czxBNrdlHPHw/7QmpEF0Vuolh0Qe/lh+n7PGPnEacgogLOa/Ba5STFytOfIL
seG+gSYdyriHb0wdm3LwWYzV5EY/u9dYOLY7wCwlYaM976dRohZvb2OTg7hF12tn
R1SNKMzMtqgdi2qlLFkrbKKu3iIITBiXBCFKtwBhjxd6YGZ1IGtHgfsa+vv9c0iq
YrUHAMJzhB7CTZPVVOTmo1TkoE4aVAxJLJ4Q7C165ZtvdjpFB2xA1+gkTCoA6EBk
O2LjJ/xBMp73PAr299U9o2al0OQfs9hYKb+XjQ+bNxOXm6oMPkdoW54rfXRjJq8U
IqBGre4+stHBH0t3cXmEIFsDRGf74cyw39VqLXFvgti+vWEjelG4h9lZYapf5S7/
mz4dn+FRwoohNNjcWzeO7cFfIhjpCWLBWyLB+VS5Lz2usOErBugklIcuunsGZmJ+
geovKDMMNdxpGkAIID3dQUo+xajbpP/vwZNcn5YBJFQjSsMuOHd8g8vLwKn7mYDJ
GLzOaHHKrDfBX9bnxVkNFnsPp5hm+jkkZdAbYfT4ljY2rZb6Q0O4XpOFPg3EOd6b
RHXwsAKactVPDv3VDHkAN56imFclnl79gxaVs/2Z0YVv5EP090WKiw5X9lZM57qX
uCuZG2gdVjjqJoUWqGkVQKzCkA78y7UJ8iMhmHr7LgY+jpLZnQl84bJSxRhLBZuf
7U6u78j4UUaFbODDFIa2mKoSQ4W0iem1Dqfri7EdZlF/td6dQTWsTZwkSo3cjhPg
qvpLc32lPvxJua1EYcAVwcYNQejycm9MGLshp1E0V4aB0fpXIZJh4U+IrtX+v4Sx
H6cjF6PGJOcNYAIZAWaqZTszQYy+hKfUoNsSOn1xi1YnwYaWIcFlmTbxrLOxKK6H
6hO1kPh8wkM8GGwidr1Uvsububuu7whvvPLhrYla0tC/E18FZIhy0mjK9gSXiyDF
Zn74YS6o6fBpZ79llyphUpRY3pQIGuV/MuqV7bokf7jWdEMiZiZ/BH81cP2px2Ry
wlI9EYqtDDfHiot26NgYAhdUkmeqEFdrB/jsR7NgThNnwOwF8mSOntYhlBE0kCSo
s3mNCneAQM4FvukkWLl3NuY4XbVLXBGmq0n0LG+1syJC5jv6ckWiC7T2oG77DsAM
03qO/BcVlQxMtgpBSQ7lU2xGW+PTeJbg3XNK5XAfrPBKv0mvIo9ljfrBnwFB0ZvG
srm8Ii6Ez9V7ugZCqMF8Us0aUsP6xOMm2GhKEDhNr4EfSaJvoZoy3BFHiyvlqqge
FmI2cfYy+FgdS7ausiF2y+b+0OXihX2wWkLZhc+M80gy6R80ehNN2+vjgJpLgOBN
UQIec5UfXvC91/ves4G3oLp1AkyRIqhYCh9HPB0BuFlMZEpRWPr70vcVDzkgDGQ7
sXtpph4zCLPdClG5yXgjeZgg7MYqtOFg/e922YoogHeUcM0LZuGqBtYc9iOsvdbl
FLuhyA3Rkh0bTl5xM46eAK+/9Cm6wEu/rX0yRNcwqaS0rPpS+ScKSvcvY4CeC0CU
+BUbREOXSdkeuHfikBQNbmuidwqjgeUpBDGSMpAz/l/8yyQoymXcl7ILZYTG0uAM
rMmGIEw/cR62D9X1qnvQT1Oy8ff6bAM3YxGsyU4H0iGezHldgpMtahRYZEbZtgnW
QLB7VRz2QBaBDRrJmomf+VQROW/BY8Q8sdTCvWZ9P9TyKA7EMKOYKzxlKMn/jlP8
OHUpThxfhX4i8rT5izGARSlHxMfwqGwow9JqEHm+8cR3GRJn97RsX/x9JG57Xv96
qEncAeXQpdxTshJ9I+ZCh4jq0xBLacaQ/7AlJ+wv/AMfPW9QqMfpeJlxoEGbCRkg
g+YH/hDbs/+YMvVfI2VYtSNl/QeWAdEkMx+ssjapnvWncTGgxVsHK10sE2T3h1Iy
k3+jXnM3TzIFdLc8F+NUBRkBsnyndo2DvBaAb1vH5MT5Sa5h8R7GeaDPL2vJN9RM
8JCQkwXx8xMWVdadH7jQ7Is9eDKDgjm68GE71MkloGOSge/pTQREkueZMAV1C2gp
KJqStnVb0lSvSq+5GFM/GVz6wPdrxrfvDmZwSM80drNB7Z8f9cVHBpT2VHsrxWYc
7WBHB6uG6gSGBN/klKFENW2xDHsZl9Pg7VB96VrDaa/5oDdgnrpJcsIFL535bf5k
4uUpXFfo2pLDflIjPs7sYxS+zgwWXo2oK504Je35O9j9gaWS/lj7ATKoKdqvPZRk
1LdTO/BwS5TqgfKzsHyYxQ20uiZ1xkr/0CCviEBhUduDUfscbiB0uWcF37cNEokA
aDeICLNiFWBwKl6qMCTnjrTOHkv0hkJDTkIY4VgwAyDQ4bEt9kQT8A0BX3Tca6Y2
xfTIHgYhlX4hZFfxpfo3+O0vBd7DIxY2KJWMouwkpIBrbSpxA4olYkIrr+uMQENV
4MAQYT9y17RSfxMi4B7PXTcrLnHV8ijSkh2mcHwysZnpxRSlB08YfGsAGA9X4/1u
dvGa0smtIX3Kn92XD28+c39BE31aQ0vSEPhABTwSDvXaXN4CjsCqJ/eMOEmklDdh
d1Q6uERngD8AVaRNZjIoKQ==
`pragma protect end_protected
