// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:05:33 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
rpItERR/aeKc5bKCjKsfv71YmA6/u1eMB1BeX/fOsuKmw6SWLnC5I6ZJTU4vA+0l
dQigjDarXtcfsDlA7I+AWVE4Ls9IEvvxdUq/SqyAxvsGSW486NTnZApOFgYmqs7r
fe2q87yX3OSGNb6GyGJpF5fZ/euyA3+QBgqe9vMGlh4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 26032)
JsBGksDOfNRrGBzSt37wOZmavsgf/ik7cJfpsfdSdgdbjauPrkS0lnImW2AYSd6w
On2v3ZyYYx2oxZTJZDQ9+Y7npYEGZNGhG2MLKzohAp83YmFE4sBqniRbkUjDDW1u
BOzr6twEEq6cOnIWdHcvs/SNK7tEM3DEIVs0ZBFBhr3wAz2iZ7/uHISRrsZI9vrc
xJGe0hUrsAcY2Al1S7uoDpdHuJYb44lxlGKNalhVq+XnSATaZUeGFgBwTdgZeESy
XvQjAoertIQDok3+ydqKxvxeUegyFedpKoshu3pymG8T1eBtBln6gCsC5a1ECbwO
7lz0t5eA1TKH3IN9TwxkwWMmRINuP9hLDutZwilPyoA8+q0W6u/vrE1O8DWw2Ctv
uInljxLmsyJyOJTEwEpXpudfnaqQaOnkyOlDANfwo2GaLpBAcjo3llUtmQsDuS7D
mXzq4+2b185u+9myMTZm071qqXxcH7m+xB7lHOEApHhaEvuKAk31EZRVMm3/BBW1
7bZh3PlyvkuKvhoVCBKTx47YQatB37qusq5MH7VbFsAC9Y0HkhxdZEJyjoxv8j9I
s+nJentyH9YdlBagNOGXcPuetLk6tP88EY6y6PfnJYcblAJdWXqHuGue5P4gitnm
1vsyJPSWLj7ucC9ufGgAAPjQa22qBTG03EBtx/A0qOk2btzuMoSjF4dl9S2QrzAt
0EqYoywIP1ryZPxERsWR67E5NdcvuX9bWQw9Eb8J4CCRqQJ9jpyGa9IRP+BI0xBH
rittqn4DR5ik4M7JTNHPa/+9RzRRXlpUMqmRM+xy/fmDewevuW6Hq5jmxbtxs4p/
rfncIfQMP2KW5QIK4m4Tdk/1dEq0Jkt1Qwdvsx9yTAaGmlOJuCI6sZQ9uyI8PwV+
5B9oAB9kxs/hWkcefRixLl0bPT8N6gSaM1xCLCDcB9Gf4NWzZ/e5rMv0jfzSgtHH
LSISNwQd/9d+A6g0ZN/93XAf6qvQpV0L9erAKCRrTfFbn+4oQWoZF3JYtgGfRGRd
bfPYcOLytMMveYUh23CUkqDvx4AwO4b605S8zlB3d6GgVvHnL/0F9S5Tmstyaj8N
eRtj6PGe9fB1PptH2IGcBgrVpqjBfhgUZKuFgco7fjUIOHJ4PKFzXjVJReipKu3o
B1bQY1VkgPrB1T9WSxhM009/CGOiSmMIy9pTi3iDmIpOcqwOlwhEGTv+13L4tZYs
B1bmhpMmUgXxMYhEg9BJKgVQtM2XucuEjHvVKU6GJShatfCXPtfdCSY0W8cwEpFb
aQCE/ydx6NNevix+o4AVooMLJIDqeDtf1gdTPBd5TYvhdHKKJx09gC7VqVk9Z/ek
6C27SkpeZEHM/gLF2qNB5B/1jYqGPLL6lUeMQwMpEfVeBssE396CPpKIL2QdKQSW
6yFJASFBoR3HG547NMIH8B5ONSSqCnjWpjLE24155rIHa8q+UtQoVmzd9nAI2OPA
3Vbmb6X/WL/Coy2iI1/ohAI7PkXJ6kf3R2vuGg/sl+mzAvulL9erZPON5S5RuDpQ
sXyxA/+ZO3KZYD26zuYafTlR7tVlPE8WRZIaLvrKLyc2zs0jCavCCB8WW4oQw/lJ
iiAqjg9U2y6fNOPvTk0KRp6gH+hIDtmgoekvRnWrj8GPhrxQoc/Dlx94DDXhLPrm
Ve88Gm3nb093+hQX3rb1Hwu6gB7H4hDR/7/2EqQDlVQ4HZ5m7Wgs85uCMfo+GhJ5
OnHMh2xbFCZAU0t6EPotRlstSVSw3aAshJVZ1RZH/SobctX2IA8ScSPcowoAwuDo
jL0KMo+QEeSQ9Sfq/Rc0Z18PC9xl/9ZpRu4mHswtHVWZ7wrja2/KbHj/mSyBgfCe
ja20vpLn2tCHZztUG9QQU66Z2H4/bMQN0P9MAxShEzbo2M/lF+vyIb+oqeyWSgrM
jOByG5QgdtmF16nt53cjRxINeukqGhJO8v4llfxrYx4vFAavrJuAax1d6xroGa3L
u2weu4WSZ6qb8zF7HijC1GAi5Z+LvPBxiMzKUNJtuvvxjnuUtPkydsF7d8fBdL9j
WPFSc5tx830FAROwIlL4uW4NA9vpWcRV3rwiQl+DrwjyzeMXx5UsCpQ3MPgO9tQV
t18QQB9K1pcVRs4r0r/AW35l3yWGct03QnlXvINEDm1NsxOhkXo2d7PeiE+W+6Fu
KFKozoV0HYB4g3WzA4sIVYHQhKh6tYbegTdsQ+b9NHJ1BSwfJN5G36FON/eg0S+3
r1lgrJu0R+Kym/47piCBrT0+MVGFDRS4C2VJd8X32sSo5G9xv8xidQkDGfFmdSe4
Te3FXs1ewQA0T9XHwUQ11MrnXTZy09lsdQL0SOZiSigRvbjrKxA4onYMk0CE//Z0
mw/3roll3ISPa2aGmGIESABQ1pl/k7ZHu7/R+niu3OI9KKoJrgOCXynYeUB+5hNU
7QKvocTgXxrApUvYhRXWqcGagus6mw2rkDpEFen5Q/MHQaYcP+PIn+Vy7F8dh8xi
yODD6FMzgOY8DlkHGTzLwlUjBy69WYvvQS0INO3Xz0kxpJJ+QFcI35ytk9iiCAIP
MdKquGE7DgDx4Md8sEATMy8qrexypzlyS6VNoMWOuZitl3E5RVAyoGA78C7MYBUw
jGAXfbl44B2RjZnSC1nP41WkCKSBJClFo/lmhzgDPfRIOdzlkJGTy1ZCsyIfuAGC
oQOO8ZzStHFDPj8/8gUSC7vdCI8jVYCnzw4Z+v8iT5aLk4c55nxhqyghtP8nqz2K
C778/1VnDmA+9J9nYwSBt7BfoQ2iyvsHq4+43fpvPeJSA9Rrpadjo651mYWy5M3F
1cXfWUY1pTShShmoG+HjwWCPuV/Js8F5CK40xSPlIgXRx0+A/d5ujYWFK7dcIuBm
8LgtQiW8WMZB6NLWxMAX+nTr8AqAGviqK6W91QupTAN+OvjnjtpMp+28UioJE64B
4kaFsBV3oIqJEjt00UkdJZg3Gyxd5if4ks9v+RSs0A/zLJYYORCWob5ckIbzjj/s
wjlAUimv9sNXJaVGCTkI/MoLwCsayfCW9ZwbRJIIfgKYmr2guJ+Pif1USJEzf8k5
VFFSLBNLKKnpb7e/2AGWdjXiZcy0vBAbioDqHh8QSN20wpBFcnl9gHhNRaZriZ2f
UoaetmJMzR2eoNfJhl5dodb736P9ageEparIp0IRKj+wKcYw+3a6qMxyfo3Tc/QW
qXxOL1YqmEuExzbLpRdmYVyoE/pX8E5mWdL7pcphpl/KKCSMcW4NZEViZNP0BRgg
3GON6dLm2iK0s2O1jqO7IcZyrDqVPrGxyHqLM04tMfNvCMjD672sg1qjpTCot60i
jX0RlFCKkoLy8RTgMiJJNh4Al6DpAfmB3sq37t4Cz7fN1lwl4FTLEHpA8JKLxCp4
AhqUBVh6TwOem+8JNTboEB2HQSoxTyptwStGYGvmr8L5KwuucH3a2ERImlSHW7q0
byrA4WjxSl6M2DcKxiy/jejRayzKkb3w+v3npZbJpBGMFkq0/T0nvz/6I4ZRfYes
+xMLXNce13uv9ZBev7rnDul0KZnQknF2qxKRkJfIIQ/YSw11+uZB7AzZzkyoLMX5
cCKrp2cDzJu1n/FF/P2B4IsqIEZ2HR3kJtLrhFP3TeXf57jaQUWeEW9A4BfGFKby
rT7vRyT2uX+Nb7ZVeHj6Dx6U2gB4qgSaJqlGFhcWA6Q+KQBM/OO0vJBV0rXRqkdI
l4DIIUJI3Gt/KVg91LRTe1sCVXS9h+nUboDmfZ6ESniyuaVnlEZRe1+sgRAk5vun
7kuy1QOs45g51APONq5zTr5knbgYKIrTTEdnJw6hO+BrviBLN5nXhpqDR1HEi2yz
w71K3I6wgjV0pgzi9qO4DF/qeJpMXi+gTce0mHxI4xVFQa5AtbZ9FS5zKIh8abSc
DMr/7jBAMFLCuVljPaCcJABSf4q7u87JlIqUJiXwx51COfBA0BK/Ctz0+diUYBK1
B1ffPjKUr4v5EIWiQsFyciBu3UNl6VVinMfaNpjAKZ1fHxdv27C7c4IrgmRYk7Ml
m6Jo2rtJAEFGNpI/cwdWFlS9uqK0i7LGIH6JWS7H8cpmgwelRePNiJykNRuDTSYv
ZXuP7VBWE5Bvo+MIg7cSoCBOjtU0m8yWmvaHjE7QagG7j73jshP6yAN1lHl6hTru
rNl8dPsd46eELP+9aHMYeLpZ7FoB5VxiBhCpZdw3dbLbvnwAazognt+umjwfqIjG
QzaOoUJ6qk0//FbNQVW/sYCne5axpNixF3KxgTjk7xXu7P+TiQ+XNPRpHekHP4wb
/99a/OVd2+Flk/0bQUc6vZEfVTb5jA/ASuVDOQooPz5s9oiqAIaTghdtR3MTt828
956bjbO5H4w4MlqkmYGYIjSmNkyQDNIDmwFFWb+kOhwVLfQ9AmcbII1H7UGAUHTZ
hr9ZjRQxKMGLYaRLkT9IjgckKQUsNB2mdODihyvJNWP6b2c/KVueJ7ObCb2UvNXq
SYn1UE7/qYsBL5pw1mbGNBzupA10ebMn7ksZ6e+Gg1yQYsXXhdH77uWCV7J8gE6u
tSHwMkSrbJLH8J6YttDU1cQrD3c2lZGWSf5TXP6SGRpYI7UxdynR/kpAFoxJ7mdE
b0N0uMsg526Rn/eHEEc1542EP4onpz7pRKztNnllXE4FcKI268yCRNCwEBwUhA63
MjESTevW4vJ3PQI08/SUNfIvVbQhuBLbuoVT9ELfbTx8xaWEIZ8H77Ymit8SN7cE
UuTVvJqy5ccYt6AFMv1VkBw4YHqQxXDVEAXRYjyJ9EhU3eSyDQzVzKnKPIsD/Gn2
wJQi5DRisQ1TKTP0k9zYNMV5VyCFBJ4dhje7lESfXynKuhl+d/cq6ckIkYy2HyYk
Ivtsk/LJCD96r7TBpgsasVAnQqXKoJNHD+Utq9MbdmGUxZgYEWKtFFho8b74dFr3
CPI/Ws9KDPNqnPBTwQDHZjlzr5eXgKBRqWvxB4W6I+ESwnkpmQ1bFhcldrHXRBu+
fXdEju5UvkJAlLxLewT1C6DQR24eep2nsbtl90nVxcFEHbS4fDyHc4SosH5/qm9y
BIC6oW72BAmibvepa+/2KX1I3eJG+Febi20GR4FDUe1YVUqWZPnv3sqcUxTXhI/0
CbgIBPafERSZC+p2VoeLjwKbyNJiiEdtyCJGuslbmQt/OT4CF0gYYrUJ7kfij1nF
3c7vlKOA11Pa6jF0UaV4/lsxbn9WIx4vLD4Pb14ygjK6fRC26d0+zRlGKRV45YF3
iZArlJknlG7t/UW/GsKAY6GE2HBpnJGzszsiKxLpMQ153hr6O2h8pfZ6X9N71+Jh
S+e+t4MQmynCBw/5IeKs/DmjtHNHUtBWbeb7rrxssk2PpYToItL70vfJFz7qMqGW
KQcLfUPF0Yfve0YNr0SfbCZh0q2il6CyFDcREuv/J8pd/xtDEnFZIn/UwFe8JZCC
z96qGVtvcJr6OhjRpovuMHA6bHNpyzJ4xhd+K+5Btoxtk4pRa9xoX1KhYS66j1kZ
f+Yt/q6GDOOOqhUpi40YdbYuuhoQPD2dcMchlr8Zdm95QNNKaQ+jivZT5D/mkAJw
kwj5Pt91RNNItImrTQcNM5fzbLrYT3Z5qOW2shgskxyNmVp2jeS4xz1WVpCY3tEO
LlnpUe/HuE7De5S0E7Tp/8xsxU4duPdIlPzmTf4XYzUg4G3u0ayE7GNVOl7gNuzq
2obDXA3GJTpe5sv2EMBE4KCK1R8u2OTrfmFHgmtEgHYRpe9Pqm3YoYLMzAlePR81
D+y1B2tkmE9sKqKh/zWxtXBZrjnGgR0IgMnky80qQ1edK23pOiTan+DcCgkiSKMe
odrcrEPNn6OZDnXwwzrUA+BFy2JOIbAOn+BhIqAAGxBwAou7gRu6oPnAi5hyx+91
DqhpCAMJoNEinshRBRzczcv/t7ppR2j9l4Q0gzfe4IdsJnhU99KhWfymxCXvHuLX
eN+k3loRaE0IZdiwsMFwgHkU/NVhf83XMmDyX0QQnAw47NAPFdm2bEIy/nL5uxZn
IsPf0jNK6rAVekXnCFPvB6m3xfde2vNLRX9hBs+yNkyTWnIa9dOmcEb96+ZRrofY
hi0KMm4X9OqFBoD6nE8uxwqydAQr92W2SImzefyjQzeOxwRNowUdWK/hvYDCUsF9
pGgnlIt5x8dj3tNC8pUwo8O9RlIdwRU8HSPeqV1m0x/I4rpdHIzHN3Db1KqSLvwr
dtd41nY+gaNUyE07XbDRqL7Iu0OrxrExsTEJeEAGtT4shrPvLrYAZbmw14qvUmNC
uDvev93m2aaodAqL64QEjljBcdz5BotJZcwjZlFo5I3aM3J2szmI97ipvHiRjF2z
H0iwCvhS950zDgcDbiviLM2zvRISK3dcQ1i+v2proageVQhE2mbRyECxogcQ9I33
1GX3LHQwiD73XxfLOU3xfzOmkiSFbTU4rwgYKYf8FCUZCSWfNuKdHwQd8FTRNGVN
ggRHQSdHj7I6o0U7zbu5eK5pdKLuUc1ypSoPkQlgPPAbXidg7+iXyfOrDrLeWTX8
3uvWldKqurAwn+k6LxTBv3QTtwLGa7zZEW7xURw7PTZ4xHqCaXr6o1dci7VPtMHm
QlSmmD2F2+8OKlb3N4L6OvjwZzZOkRvzlkDlquaDHgOi2j+BCQDahvdrJcJaPpqr
vhI7pvOVduXGftdXENdf90JnAEyM0fG54In8iKyWvNf9NJqWbAgcdP84Ofq/Vv92
Nmu+d+RuCary+/Pq4fNb48ZE/1YlyJFbcVGOBiZBg6neoI6adFS0JxUeSldTwWqN
vqFPHHe9FnDhdSl7jEoKz54AcUB9hUl4Y5zS++E7nvSqJFeFPabP26d0CeKqx1Sv
CqfBLjguxo/4DrU83aW20FoBAjGY3g7EfIqPaejeLIyLX0x6p1C5DfiKt9e64nMJ
xWE2vUi4mwQp9968mMC+VYgA+wdXTWmq2ryRIQVhOqTL8OCc37A9HR9p6L+0Ln7D
p00VQQ/GbQ10zFBxFeCGHcA3cUb5MV2nKwutbPVCgg/kSAbWjg+W7VE8dUUcisXe
217NJYcChFgYByyfGYIY1R4fuFOnci4QOr/A8fjhR3KKhvTIp1w08jD5QKf9H//F
730YXZJEMya14z7e9R3hW+qttJrIxgrI1m4mzRG7CGGpjVKq0P+/HgYoEaFEjTv7
4NmbMRzKDLfXQd6QwqVBoip3CgN5Y45gAT9OMc52E5EYCu/IC9Jt0PpG6kspeAyF
ZTAloTL9owvZm0cFcasO47ObOt65qOU3/tc1pJJd2mnHiVeBtCWkAy33gYYg1nky
Cxb0BvJx/GXWrXImBQ7zJt9Kj5DF+Y5JwALuuJD9WeQl+eVRJykASX0R8QKzGdut
HwJMltVXdUk+tN6uMZZtP+mthTM7wZAfXx5hshsMkgYFRUGAw4AnlootyyfS7YWU
jVkxxRX5upYmF55YgOGzbLTvK1xo1g030iwxYFEESDdcI6Jo+nT9F/XL+roKct16
5/CHaDQbP84upRHY5ITIHhAg//tmlkBmW5DXN/t7Z+cmh9Wp/oeuK8Y5EJ5e9nCD
j0EVjMoV4IbpMD7Hruzn4OmrdLLrorVDqIwc6CAtGAnDHhOYDifAZ1Ys6o6tug8j
iEYjfQ9NsZ98gKgrFYuIUzhfQeudUwzHQ1BXTNI8mZ/tUfW7AtgzLJA1BqiiyRXf
6bD51EkshFqGgS4RFx8CIbyuv83F+RXQcVDnbHyRRKEvHprLs7UzE9YpCbpOZyOx
TQrfsveK8SgogTu1X1QAX81vXLMTklJ+ScNF4s3OPeVnIbHm22cYjFpcCR7u3Lie
kZdLyeEysLddgRepl57aJEFL2A8BzG7TuL5rAMWWAVNzzo81yfQjCu50WwuCU57p
UoH6ylC9n7O5XZZH0w/Gi73bJngYEzxjpC7JoMSmZPuC6rj9j8g0Hbb6MTzghuUy
yDK94lA5mMihNXOG8H8Q4dfFDojSMGbB1+Zm0PtU6DAk9l1+zxL+vil2hXA6rXbY
xP0QGFzO0LIIq4o8jR9rs7q/+Yf+H7gU8Qrsaizr8EmEnhMZvPkRoNYI187bSTVt
KYoEC/sBh6MAwVk72sdLevt/8pCo7frKDoQdhXh6qWlQLz5VOYGupPsDmM3MufG3
CpuNoYaPiiuNLyxtZM+Ah7clklOk/TMZwZTzvWmeBY27yhEnH2whDZ9D3iLBnLeD
7CGL4X+MnB+zSt6TGJKq7l9i35gBFW03L16zCafih+68qYfrozo91dfloOE9PfHe
nDnIY4h4ryGokRiMMHpOsqEI5zyc8bYN7BX83PB7/lTWRpLzEwJ5a7Le/C5jlxgK
wipKhlvO35Eexo3qlYusaaQUbGE8BPe6nJFouCo01JLrgq2VV46NKZWrX+1/fMUr
j/XWpx0UiVNPx493RdRbg2r/vwDI0XbONjxm4uxwUCyf/6pexvjuFH7zXCE7vSGe
8VSvSkeS2l0HyogzavrmlIY9ljnoz1A1dTajSYo8aQMQhIXLRSlWf31FXc11n3NG
DUzOGd2RPIHnd5L8Rwo3W2gZ+nHchzSfguluaxW3fmREYOdPYTYr49CA1N0IgeDR
Twvz7T9E7vZ3UrJghWDuLw1c/uLJRZ7YI0GqGtf/KP9Cfad/9rD+rl4tQ8cXyOav
f/6IhV3LyKZJgfUvzjFwq3gzaE1hzEO6+x0fXRxIZONaCdA/03r1mhtb0eHquumC
7q/0bOLLskOVrfJMnI7HOFGKrK2HowsjycnDzev3GVw0Tm2zTfWBdoau/ttgBv/C
VhnuvnEK7eikKNX6IYnE7WTTPhHI4fj6n4JsO13nTWOf/7L94m2HJGf5w+RJLUYE
QFgj3PEOna2GUN7+87DyUw8+oZeK+UyXF+4oAfXs422lIdXBwkuSMQyUqhaJodVh
xY9L3qTd4rhyW6Nq/CmAsjjzSllG+ZgP2KV1n5N5uBerqUHuXEA0RWjXiBN1f6R0
yLQEceFPPk/+zJQdMmQgFewBd5+unrrg+BrL8hQ2ejsBoBl5PZt0q2abHDOsbXtk
rGHRAt5gELp6LQelzwbtdFpf1g0tq+Dm5Aly2tHh7yaFuDHNZmcCcGczfeG7rdOd
+CC+wkPkXUAgTG1buBHV7IzKYhMokZ7D7qG4fGTKY5mv6PxbWiLyIQ6QAgH9AL8F
mM3F2DuarEffaHUtdTVnewwLAxZ6XozwOQ7lD38T8NOA3R8EPTnNY/7k9jd02e+4
wdFEC+1jugrk4Qoio8fjhlillkZ3U53lnSdWOQMgDCOceyZ3/vg3HiHQQPh9FIp7
yGLIJJnYaomf4ce/pshRDnZoCYLtuybJf0PaYgXOtEGVA90ARdxFRh6IY9it5S/U
t7gFf45phyLnV8hBW8WEtNhqH6Bv1n9cbX3z1WFIzsbgbazxPePwlvArB4g6JhlQ
JHmok5nJrCx4lFpE7773q/xxbQoX5W0RTH+sgTvnIm9e23EgRg4Hy8KVU+hVb6VI
JiYvTUJfGQQ2cO8nJ1yE4MzNS9TgYOiupTlm7eMOFKujgo13Op8nEUM+fxqbYsDp
lR5TWa+rPAy7aaMudlyyCXw7eVgJoTeC7imoYrAzJKQMxwx5k+HQIJwZ+rLRJyiZ
QxjbawSmd3HaR5MLaNY2hYKBg6Al+koLvne24+4FJugeEX+3pYN+hABlf/sp0isE
O47eyzYtQtNYrLLyxC2rVqBOFISQS56Ivrp9tzaFG3g2IHW59sLR7mhOp3Ftewo3
4QtXSrU2q1FkUZLIDSJFqlSyd2IPiRZBeVVboA6tK6HWJXekoSd2rQB647QGLJkf
OxfpTaSyQuw1hnzw3kRvF2/RHMTTfZgWy3xOtSq3aZ5L1ywG3kdyYaD5aJEP+EbW
9btK0y1XHosHzGsd54zomWAoUxjC18wT45xzyMsAku0OHuKRcwB3odBg7DjNTvEy
++rVdQ6E93pV2YvxRXolFGBye2WbUVYFSVrY8bo96qiR/ZcpAUAOp/CfEePZow+0
RZCyK4vG0UHBtI08issgrHtGnE6dBspOKAbVZm2ITaTvuH8r21k3jXy14Z9PWGMW
Gq8y4vE2IiCj2sIz7o6iXkcD8oiXfviaQfb7I/SnVccouUmTJFSrorvO2lTjV8xD
FYQcDojJ7J9Ngs7+t08N/aEMJgPW/5my9IJRYZnnf2cgPC7IQsUw/gUQKj+mJg3H
h0Bb/I/x3smu3AetnlXKFnugLvRS1iwNIT2IypeQU/f/1WVijnuZkx7HNr0FKY0c
8NW3WWzAC9GJ98sRSYgBuuJ/7RxJpvcMwg2bLlz8PanrvmQ+oFHMGAodnnw9B7Mi
M/l+KB6U5EJ0Xc8Dhtdpq24a4+/716DeHKQTZy3QFwtYPaSJ3y3+A8zw++BMBIZX
7EiJqMlMC1b9w9CD2Y+C40Gvh/gTZLdUaPTdESTOKBJavfVREmkQ8GUPdn95Hodq
2e1PAKupc3nXKNBLTKjui5Pw10be3GOG9C5p8utMvTp32WrXXQZkG8GncZEKIyn8
ZMXo4JuHf3olocxzqR26gNqZzL0+EsvOgv6f0ym73fwWzL49mCIpuTxH3a6l6Tdu
90QiaUT5uefrmfLa8Bl7Hed4CWDR0kwInpNt3POCvoXHk9Vu1k5NpkKzuQaiWXsR
Lp31SeDXs4kU2qyQl1iZHfJKNKBvblxg10xLg9ioxj2VHqN6qHYeJBx9mc4Odi/0
ua1Rr6sBczIpkA4b94SPAjMJfFIe+HZTXwCXmOWeFtCfQ3l30Te2W1DJ0EfvmmuS
A/PLBECTOuRN6nBiovWkXnZc3wY2hZfmaEcMZC6yT5zmvY3HDMEk6cdooJs430zN
aU9A0fJ8Fgcg5ahn7DCtA2hdvsQyECaaiQpAYH7nRbijCHtO8pylxfXq2EGQ8lsA
1HcPXeWQuub4FyfPMKyag/HmnWm47NU8Z/f+1Xd1w1daYB+frL0uYf2mNtpS/KMx
wpPkAlX8rU3V6Rc6EXByrJzrNgRd9R3RfVXdi/sh627M7Q34mbCZitTK1FbWxbIS
P28YIJiorzVxkR6a1FbkQ/jBVnKU5grVAwgs+HLpokKUSjI8bfxm0z2739IgBX90
Ys+U7saaIh5x7Auj6x4emQnN9k47TvAObEFqFkebZZtEr1lKlR+K4cp38p5xEvV7
GsrMBmqJ7t2iRNaLI/z65NpHEZZQEeEZ2zK4NNhne8/WgxxhZcPzq/muMIv9oKs7
hIJbCohb7r+tTsfdnqvkrOC7m7SEDSS/Qey2d+5bUWJX+NWSj+NMMHfznaR0hc/l
gjgZERTvtXOuq4e3Gl7BfHtVAWTkxsg+FmGW7AF+quJpxxqbcjEFEO3NzNL+CMFW
B7QGd5SYDHyFHFA4CF0XbcsYiCAVR0S+rJQznAbRlrE4FzO4c0++SSQVQpaeR1rr
KMnAf181pEUVvw+KsNWwBiGcz6EFhf2vjl/imKPuC4o/PzwhhwE0mTtCjnjMwBED
pHsdnAFC3AMQL7zWjoT/clfm2tQNyHNByzVBCEyiYfh2D/emOwLb0e9mFUFrMcz9
OlsVmdlJ8v71OmeUAPlkPp9DAiR+d+5EzWHr+AopTq6r4Xn2rh7ZYqhzI8WmWB2T
zum/3OXzyXyEoA7963X5Sqv0lGMai6z/udRt78NoUUaY8iUWDUeoyqOXK+gDgua3
wE37wpf2E5qA1L6o1qWRej6MmlIAKSov0B73fXAiErOdlmK41JRHsI334MLG6MnK
GRWhYIt6EdjOUNIG0cEYh552JdFaskF9/LVGXRUF0ycvzo2WUay4CrIrc93u6EK4
5UF0X4iJ3tJYTebkY795Gq6ERDTWDHPbPVN/AaWQ9rSlUda35Cuts3tgOmmVRRsT
ZeyiNwnAi+++UYf4kL8XVmFDE0QCgtMYwYc2LiKNit/0nckJScYFKrHe5MxqnLka
XCTEP/boy7iof9HJjuOicYeGTHN5KB807MPLFUuXste4sLDe5BeA0MX79fhuTV0f
dml1JSb9Cgxqk2sp0dZJAUMZz8F0fa0SlVxwlawIn3Ca8oAGpCqRwP35npPgHvVA
C/lnX35el2wAgc/IKf9fMXMJdiJbh4TxOzbzGJyeevdfAdeO+HKGQmpyB+th4og/
GJxogH4kXE1nQguOkm1kqN7DNsy+wQYgOa2GuiVkQbPXnznoA6aZElGmWLrdX7QZ
6eWFpq8uyx0GwGsh+BeC6+qqwJz4zv6ECcjqKsTjbMjlPSPWUZ+Gzl4i24azW2dZ
V59kLlaUdYoPm1UxBI3aJ19lXgQGN9Z8pmyYMIuK8PKcSO+nD+GpR6RlmeMZGyWg
dD3YvZNxt1IYDG6+ouVm88MilgxZaCzagWdWBC3mvC7N1ttCptgz3EEWQFfWIE0l
v7+JlK5yAaYcfe2H+Fb1YGmFmwVxI2o2oTOSwaitOf+TIJM2pkXq+hsGQmGLT/pv
OywxaIQwr33/vPhAWiVtS5lvJzRACDNg6vvPyWyHbuACDl5wVmg2jCEx+DWsf6NA
By2pEc7FBLcbbHJcneIBh4kYALpCAiZ/vvtenkmEY1FASXBnLUhgXTb7N6qR9BYK
Uj/QT+4m8TzYoNJFGCQU3PwmjcchTIqQwFlkjslM6cTZxOIRRXxWjfQIx18KvGuK
zB9OsGMQ/8qHq3W8WH1uT+qNZGqmyO7CdzZyGGFtgSXmoyfLyMliP5NQ8ChuoIWP
ba5+SrSalGIjn+4n2ClGmIxnAjyktfBBxylTpTzIUPWR9lyuf0sIwergT4XRNtxk
+NIupFu2V3k33jZWr0JIFC1c18KZhvxq4EIAjXb99CltlQGVwbNSfqc/Z+0GHpBr
h57ZEKm1YFVhrCtQrLwY9wMuAq8JIzZNAkuyidXELthFoOMEwIC6v7NwpJFIMFMn
rIywY4gDzT7TRF2Eizb8OJ36E7eOdBEPfoGi8hcmthZ11AhyLqbSPPdAWl7W9irK
WIP6aPKUIV/4y5nH5AfZr06n88dUWR+JwH+KDPPCg0jxa/diyObWois6oi9p/8jC
ADqGPTw56NAO4V3auJv631s/NQu9EIUy577aTHJTFNTKPgz/HnvVsugRJm/HePKV
goGMvNXTd9WNjVkasRg8FmAUldwjyzB3DnIJQAXOEJ0gFpjf4hqGWVCxlDKD/K/z
rOoLjxWvRNxvxmP092XzB9bRKYGLwReMGTNwZcsmHa2I5aS+h8ZQVLK9HWY5WYBU
dTPV35vxPRdcazrN0wYEy4fkUb+gE5tJmtaSn1qi5TMfWP8s6sKiL4d5F1ZVMZ6/
KYLkFsv7p0DGf2QwmUnLswMLqvXM9SafkvwCKseM8F1CAtBb7Qnfy0/A0O5cyUku
kF+n8PWkMkVPbzAoPmQiWxHtO+4fR2Is2GTKn2nmdcghIe8TP2SK/c0mBcFTAE4A
dRt/uFj5OHpqrn9oUA8wKa7KO0iCaJ7AQpRPAOJTJlOmhdtmvWb72StU/jEV3Z9j
/D0hu3o89dcI291Qbpp8qf/pfs3yZKa5YzJ4aAT/1GNcbwGVFLAe2UaAeAzwKWge
B+qiciQ6KGc49ftENp0zSu0zsLrAycQ3ZHbbXN6rRdXeKfK3jZeZBohUVphSrNts
NSdTeVsACld8TzecLKSRAi3T8Od8JmDfFXaxM4CAEfH8AoLYVgvM6ssVSue2BgCd
NncrF3w/NcAw7LDCHPbCtNr7p3tRBSxetCr6GUj2fpCDD1KHkREyOA/QyWO/xTTR
F9mXlR0Pu7Nc65fL5ntlRglEg3CA1ZPlR9jIv2mN1STtQUVK4A4nPKlQe0/e+6cw
wuhT0cJSIq3fUYQD6bZReHuLkywMN02xzkCCY1HXD3KsGJlp7rTclw3TtuRZF+Ze
XhViezmsq6fYXbOn1lzoKRfA8p0a8OuHXYvdADyQt1dBh0Pqw4u+Rl840e2CKOcD
2F7xR+CfJMFdJg1hI8JznQx6pYnzvr+8CZEWFpvcaXwn0dxucBAWRdJiN7U+7gF3
OtjOs2lZ03W/0Na9VFOu39U8NvKc5YDWIqmBeBdGHI/rS2FjWEzl1DpCM5tIcjpg
EixMZmY9qxuNbFAFGCGn/bEV0t1LAtbKbUvVU8QR3Ofp50BA5Cwm9/PONtNE76H/
4hOmXdElM7ZF9icWyNtK3bo75SsJoz6l/ehyQzuDiLphfAh7NKeZb3GNuR/A5LLr
6NzlBsJt2XX7WcEumfpkMfkGJ+svD86ocEyHLnSeT1W+KdAkj6YftLypPwZZ9hKP
gtgEyhlbhCAz29psYouij7bGxML7Sb3Pm5Y4aT4HFMwG4UtGTmjmEdgEGHk+Me3n
92u363rE9uuzoJP4fSaI/swkCfkthZ2HWctB46JRmfxdnwrqgrHbke9pdtfqBPyw
/WJ00YWR28kzTNRlBDj0grKQ/gNx1w3oEF4SxU/KVYpjpbBk7t9LeDHj/zEf/aDC
QYbLA3lgUUG1aaW/ZR6T7RGlW7Kgmv9UOzpSYLjNIOzHy5N9yxJf8FC3fbtuiMea
DmLHI3/7ZnhEQLakWI81F6G+dRtnn3Rdt3i7pE5TigVFAjp0ZSo1gLAbY641g4al
ZuVtj+NEP9yp7CyycLMil6i6Tx0Cq8Q7bseEQSjzcdN5qbebKRMo7Eg0xKVh/ctz
9mF+OovQtKFr7Ri7odCXFGkZx0na5Aj90vRJBKvFMtvxgGYFBJVCQwgO7xOI8YYs
QIxvukHzDWwwps3s/XxZQeyZknE/GuU0PGylyeTe131nd2lK+rJbuFrhv5EoTyJa
r1pJ8tTCzc6UeLWKrlxNxZ+3i0AXYYFHmmntm/1wzKYGql5dciW4quu8jpsN0ea9
HW2HKuVc2nNPK7hbChXFaWUb6jKksRKq0e37qUw1dAwMzDMMZLKh2GdpPaQoBhmm
c9AqdcxVs0+jgclpjs0Dvarkd0bJxFjy3McwQdnNtgErQeunHWvmONfdldhedKTB
LD20+wIIgzsg5t46Ji7FCPtmiyEARN4sWxU5P09kWUaBH7had25Qdl+uGV5ExSuR
RmL3VTBd0oGB31etNan9YCvk1cBLyW+OZmVOlPZa01Oz/uB+3Q/2ZKkBELSDJell
3mX1/SLbz2kl6nVAoF57Bki4O1A2tQzQt9DIJnY5VSCnU3VHTaRX+hrkrl+tdH7s
oF2dcUVsi49rzOkzE104fDC8MQA8m9Qs9HSoaBv/g5oSpCGxtJBi6VRKy+vIN4UL
wYoPfedeqPPlIPckV+W1XKBeM4DDdTu2SgI46gSJWg1YH4z6wxk0upGhqDGs6LIb
+ZntQ63w6tmaMvtxxikX23ZSZmzLm0joGmvKufq5N650CxCQqkrjaU3XWyVDPWJW
xxDgF373MjBi+6V7wSN3VAqt0R5zPWtK7BK3JKbUL0CnX/TkX5alY2KiIGjjnaAr
Wukv9L8mQhD4hnowgMgXOswsC0KQUqz8ciVJAJAvLRt6VQPHGJBFjJxQ2cMAoe1g
AYU0iIZsHIdh+WCezWg70H2PASBs5drMszvvL4QbYKBLBgX8k6pPonV8+vGgAI7J
3yztwvbVAAiFnlgXxCEJxzTx9Y6CLKDV2cVOqGdkwd9u93xJlgHWqFOou2JWOQUM
95J6jXO/cuCOLPD1Z8c/zGmjR0co4jIkw+mpOjM8ORoYPVcLOIGzj+gxKVR7Z0Av
RYvUJTY+rZQhw4ZSRuurwL0AbLeDZsYv6YCKQkbv91b3jhokBiJ/X0neiLmx3b3O
Nu1cc/UYumfMkl6mNPD386QEXq0FZCQfmixYzKfD7mmny0Rcdh8J3uYLk2lrZzHK
PHQrbGz7hFHXUXUk2PKTk6n5qBuAgNS2HE4OfavvZG9yn7tpoUMXVpVrdcK5fOOZ
Mj9XrsR9bJuSYtr5QVrKMJ9mOW20JPPFPnGb1hcDsc7Vv00sQd6d86kzflx4QDqv
8vAPGqxBWGoUIfce9OiQ2XWTf29m2P1vM44JTvg2uT76z6tzPe82AmUuqh7+7xed
4JhXi3bvsu3QMuulrmpVPjg4r6snfpraS7SCwIMIeB0x9x4RPBNFTZw6PAePvTiq
dCu9fgLJ7JWyzgjZH003vDatjyV9f16auhJhUWMdmMsvWAByv4bh+x6sAN5taF4h
AlwzndCHSxsZZwySrWJK2QcxhAc2xKG45VtPYIejESksF2uAc/hiEQit1+zRfkHK
eWVWEVjno/z4spnSSFVNHJlldAU2SVs80MHrWgOlyTtEWkgQlsvzq6o6LvmEsj3t
WwIOTe+/QLLwAsQJW4GpcAdPCD/FGu5swdNBRcEw7ifeKl98WYCa81O/KL0N3Jwn
KcqfkC0CIj5p/oEFZDDP/c5Y5jX68M8NXNRLjkWvjyj5lYUu4mFJvaDGTWfqlT05
VldUTZcKpeiFbfPDwHKQR/o7vcIzvnLxRBUXR7ljbpwoWn/NZ/yOGrMVGMn6Rdd+
nhU0u0nN7qN0axR8tDz6rwRCHX57TWmo3cdL/ihic/zj7zMhIf+Pku6MEVP6XeaE
jyOg9N1Fg/vkE249ygyfhjyZrPcsrjBhF4LMtZLvD0bf/50ZPSkgdpndu23VGFtH
N+lxPfZQGIB7owOy7pSjzNaylYr2fffGS1GUBuuX+Kz5TvXAwmdpr2OYg7nNCFq1
aY11Y6gYgL2ibLAoJDmVEso1V9jNH7LeR08xhmgWFqd4KiXMHHbvC84o38A5fnX/
NzTQAI2a4CYAGOnWmZLjbH6m/0pVUles8MVzkTu8M8ZAZtjwy7tKY/pFUFZKr8Q3
+Zbrb6c1DMe2DFu/l9Ahd3HyCMtiy+YUmPQsDXRWE+AoaSzb2pIRuXrS8WjnqaQj
SGWxWZiIkR1cQcwQRfOS0jC6YpVFS8/VFLmC8jmEr4UOPFCb3jGBDCWmzEo4tNaG
Ff1T+8tYHfuaaZ/iECKT4Jw2t9vE4mIaFxqQ1aVyuN1xqaXlk+YF3DUt73gOGj6X
/1B3IvdrviUA3AYxFHpikT5D1YsIAlL6l+2+jIw5YxftkfGIdxBa/BjlT6DJOzRq
u47s/HoA15x9eown8Dd8a1ht6hyibBEbIiVuXmWpW/JTq0KXKMbyJgFAl+vr3ym2
HiLVYtfCQ5wdAnWKIneWC1/0WYNMATU8R1idIzW05GLuQo1oHcUCYUqknpjVQhEl
003+gpBX4OL7ZEFlD3K6+oavMXASgjiRuc24KqThwnU03vnyan+lDzuIBYpILZ9m
f22IWlyZ4lgTnA2fNX46lPk0IelSut8m0Gik8YjR809qHpCUZGaAlNiZratQa/t/
pQrrs10wVePV6Os0aYg5Ge0Pv5mXSIaqiWHqGl2YbO8barEdYIxZ4+TcPMxxv0pA
rmW24WxQHsp9yznaB943ao1GMN+KQxppqdBHbtVg4x1eudk7tBV2Y90Mu+mbk9eB
gmAfGrSbD8nmpWR7Xc8vjd99KGk6f7OztscWq3h6745tJAFEN1Qk3BkOWOjZ57Uf
ldYkoP2PS6OrQBW87hg7BCDBcPsZHAkC5fNXZOBvIAki96kcDXPiCBNpXEA/MEpv
ettIrNNr3dIfu674OL3pKnF7oN5j+ZhcMWK17tzRQJOlzYwvL0uP87WtVZqpzKLL
0xF/DLGtc0FmLV1j0AoMAshKNoouHmxE/0DBe57SIv6+BKz7zh0xaupGKATvDo0h
MJNhDSJ/GmiomvM4YpzfsOsc2bjMBE32GSyIfX4+vNrMZVcczSm2RT9yr54myCQI
9lrp9//QDUGmeYexZ1EWx2vJp1tbxwZrQyuAtgZ+Uwqf9qMeQ21h2/IGmteiaFko
QP6z5z2sgwZjgMUCc/+XkJupeMAVf7HTEi87P9XOaquWyyWUa8Zp/X+zqcGlJF9S
VrkY8uY2tMALThGhGxnat89EsSQN5o9tPt3KHjeEdzFL+Tt/LqzJNHCgE88CMHmM
eJrrs19mtofhSghpKJSyU3JFlzgxGwKLIsOwwlXkulcJ6/GRw8ZIN0QGtzzTuboa
gWEmXkdPASJNDgA2eKhgAfhLh3Clu5LmuQVvl3MSPB6ChRsEaizLoTz3SSoWBAXO
YQtTNR3Xi7Jsvqs0j4XN4croCxmvoxgrh5v4R+9XPjfzL4AjCYJALrun35LZXOuk
coWOEP5oQrKdLvuajFCJNd8jM3RNJATBaAzcNpWQ0g6cohIruOnvG/7QjuP9EnUY
sBkzjs4womp+0emb+RmJobe3s8o8MxDADp20JAEzGkw/TkNTiYIQew4VqlMDWLaX
5tkAxw5DnOLbpTdCIBC+7llzpC7tiMoGNhUozIc7xJFV/WE6lsnceg82PDy0GoTb
c+Y0jLDUWamw7bBV6OvqKqdZYFv5Hp3rM/gCkSeXgyxdqgUzZFUQeO7LyHQ2Bv50
osNTrMeQOGsPuprQL5L9mMFnAz3+u2wXpqHerpdHgWZzaWFm00Sej9VqgAcdC6NY
x6e3k5CfGFpwW+wT4SLohg3yQly0tkEpSr3G7MNVOd63ND2Z2fpq9Jil4kkGs08f
Oh7vD8TJ1UO+m4uzkts0soRSlCnzlqgPN1BX8ujAmlEmGOoTqRBfguOXdEqzB5R5
7uxpkA7/iTRgK8ZFnVvj6l/uYUSQ9xa8Xa3KU498F+1MvlGuEH5eCVkw3fZde46c
C3s2I00+l6PIMDpP54kGasPBreruaXLQp0Q2Ga3E/MpEStt6d/MM9lcSqQ/L8sM5
ICAcLOQd/MEpgZeKAWIpgZIourjZZsQ0YB2ESNWFxITRTKCE9yHoAXq86lcYJDMn
r3a2EQU+porHLGSYj0lmQGDaBDKUmLB8THFtXsTFd+OrDVkCvLo/YtvEHWAbMnK7
7JUbI1ONP+JUyt4IpIp6ffRJyzUjh3d0+fcai/74feEFZhbBoVUUHkS2w634A/yU
VOBbKWEYSZoDjEImDyhPk9LMT05WJ46CONa6oK7Rvj445qf4Tn/xEH/KqmYRGZra
PLkYAgP4fE5uZ23SfN+FffReQUBp74aO+ddsPb7tFUdzVa37YUXqq0kOk9mtnbBS
3AjZ8rPvHWk8qU04/BZfkZnkArMyNrWYyhFVk4VL9rQpc5z8Q8B6G82fOVXb0lbY
GhNvSlHBPew86aM/gc0nHZhdEmA9m/iwBcz5iYeJDh10GGtvMu10fiMMytSJKEGT
lVlCOTPM2v7QD+oJuERQRtRjj2Aclon5OCTW+mJJmkddT9KEvWf7ByqVNeIhmZr2
UP7NVQlPbH5f7DKfDN5eIGbkVCCE5LQ0joGC7nj2GsJPA/iJ9a0QBGd7eOIdbvzQ
qXhqQkum9q34f/dCEWQ4PUFLPRUW2GxHAPecBAnSVjH1Q0UUoW3MlkFFKYaXcVGl
pULkSmUvJZTjZSa4M9h4x5qnRUuy/NHjB+Tex9/Vr3oU1+eNRnZZ/nzwazF4qM5W
c8TEoqh/UNjfn6sUJER4aUCdNPjUxvhw1Sv4bQfZTdefJWRwqg2KbSMxSU/gqgaU
B2fetpJ1bxoLAEK/AkTydgz8rc1C6ag69lh7czsO9V6eB3fOmfFbspB0O9EmC1W/
V/gf7/ODmHg1Gc3irObq7ru6Hgpaln2Tfqu0sUS8G12cbA73dsg/bwkVNuqQPbvh
lax5uxukz8rNVl1K7j7alQl2dTgzGw2uUEYZMlXM11jNoCeaD50ODie+EsNdmZD0
V4ZhgtjrbFzEx/tF4p8C/pynSXASQI77q67FM6P6P+jUa+i5RQ3kwnW9wdIh3wot
abOVlAdBtePpJhNae9D9g5HRzDPseLMAyP/7NV/dApvNCDtiDMC32hLW7C59MAtF
FU5z1uApGjprSlUNilUzBeEMSidUh6a+JiLJn+SoTn5wQbfKmhFJ/49jcgeUX7YV
98cMBfVgb5nfuWrNj6uM1Ju3IO9uB2p3WFtN3d1N1mmNFhnu+uR0XvGzeGmV1uxA
vJtUxf3nIgS6YsAzQBID/BQbfIuCUEPFrb0iNMyl80fuioTEknf1B5rrokspj7yu
PfDUqhebon0G+1HImjjgwdqx93TbWRekfJ04cPcaeqPlVaDH59/TD2oy5PKVQXb2
O5ML97d5u0kDD4oC78nEJ16EBZkJrChW7vPnr5vXipxwwiEyQnIagGda2TY22u5b
1l5KopX2hZiV4uRyOPR21YzjksXHMPipNPq0SSdqxSh4fyNmM4V0nroc8D/Ty6EF
yKp4tCuBwNtL1P7RPMjl5DPIR4P+2GlCaxirK2g3vZb59dL3CHdkWOOCrtNNwbYG
pDxVgyPexY2V2aGEJPbqx5ZM+b7Ti4AxjIB0KJUcou5HGXosNDHmOTnF6VlISH1b
lPyHkVUyoRsGPjntKcx+5JlMXcgVAN3Dfa8XHjzZQpGjqiCWCFMj5Pve5E7uY6Yo
RZPkQdmr6l0cU1Ge1IsZqw0G/419FAhu4zVtoZzY+R567J8ej60uEKAfwaM2FS7T
m3U4oaM7p/Q5CPp0W4NY1NtbW4quFHz4aNhAup6C/uKJ9ENdEO63Ubut2TcVHFyX
iB2n+W0X9wPz+rPdQYtM3eIaH5PVI3bRSZwY1dP5ou4NYYmtcEhP9mGXd2xHZkpl
O6ynNHorSwV7En62aJnTxLrNtxZxHKcT1h8dECi5WUGMPd6LqyQuEPnKIYFsCse9
AoOgpQl+1est2BFaBRsofn8U1GhXAekHFMZOIfxLZ9U7tIpnoUbZW/NJW2HHmPTj
MmFGvrZLixOB0igP7wDfKUALQbu+1BLbKBrxiMfPVYRnIMyx52MHSCO8ehvftP7V
Ju/8fXV7S6vCWvGnIC47w/aLg/hk+kMmv+snFjaVa0oV+2QePM83r6jBn0YDag4E
bj2X+TH2W/lCrfK6QPyyAgatv++vjHQdHO1yYKe/wO5P4nWoQieEqoIpayFL0RJs
hgi9mDHgsbu41/pq58dYjAYB/NXpGurr661GXO9suo2mBPOleFUzm9zk2KFjLn3B
/w3HjaiFpOwgb4nklNOOIETbyC8J/9IAzWGf6HfIID/yP5fyO+GchpwfjKlthK9m
BQHosH1JQ3vRt/mJ9C54hbo7fcI3bjbOiLDKPObi0YNsHjJTrAcMbupmw1nboHHD
Ft8oVrKisXGQcug1TCSmy3B/yyXB6nxRKPrnjw5wuzqK9Fk8XHtYQJ9l7ePvO9Hv
scW0wtuwYeRGDFSm+7KEVy8aYQ6mJQcN3e42HAdD7KIICJUsz6JKypd0EHsiFuGj
WFPeM5ouDKRTeCea+Twl82f0HEhmC73jDNKCjEhYodPLgV3XIe+/J8tfHLe8grdO
K/h0WTdF18uBKUQiy9XMoWSMOzkpkQBlreobI+kE8aCtAdHpfpjm6Oi4DDtm/pDK
1TzNmN7OOueuQUFqenuDXcUyFdkHcg3PP052ZECOZuaZdmNh+UuBFDU3fUaIx5y5
ifYaoLi+SIspyjmcIpQhOuB6DNhtZwF07GJl5U0Tfl6zVJpm/Ek4IcZmsDIrvGZ4
tEqhmfQrAQ7yyYaDf0mScBubvLEAG1HNDk7AF42kRxGSpi4zuBiIbl/MC+u/mhrU
KFEMsn8Vrm+Aju6/Qg7iTZ/nUziaCSal52FewB1g5WwAOielpLWYV8309DcaJs2y
23VIFx90qb5NbtjxQWLXvqq2o4njtfuQDbys2CZVq6g69qbLJDKTS4NI3tJ7kcsn
qnSobAShQUXEM5S4Fq6T+Vvg5kETgZXXDQnCuyknU184KKckBLr5tqubICLKTc5/
/3kU8HJIV9GdICgffLWz1INU6Oby5vtVD+dBb6o89E80cf5tSkrj67alJrDqCP3y
biUeUw7D3jIyX58x05tZg2/o5Tp2Ps0bthlOERvnJzNp4AmZaRASs13G7F8dUGOR
hMczRNf1DJpSVQuu6k4ReaNH5NQbYx9EQke6z4fdVMx/qWfDl9aT/8xipX6zS51C
Y9glEEA/eGoqJqn0G18VSVUJc20kmY592a2qpI/qBMowgEYgRFsfx1IF5Mzv2rDD
r49KBhVjvt93hvpo9EYGtbZ86uj6TcElQZpZuUaRJd+edGiVa80bzAc9fmfsOzGS
J5VaqH3gZcLM3v5O7V/OPyqLLazzG+9Y1WrBECHqz26R4qi/KVF+Ka888AHFnvy5
jVlLNoL/egUYq9eENIfRscM8UKP6bXW9WQo2JCFSRaPJeIwroicJOzgTJapaxT8k
jj6r0GFsvp5B7k5W1AI+nHmIqu82iNldtjxRXuUY14tGhY3ySdB/7zDA6UfYqxfS
XeE6nYClS4km5/QFFWU8FwYZB/jmT/AVuTElljp/BAFH0Gq6bcGZz+zJtt3T3e8H
41uDgpt3vGJTnEP7yn4NRZWpc7R9Jswa564vSJmq4LniAj8xBhovdrR6nqg5qfkb
3dPievzBDqw5fpm9rEdiiVS3eFGZlIId6o6Ch4Apr+7Yqm4LxYqMCBSf7URv9G1I
ReFXLr2ETM1kdbQQ9NUADfW04maXbJKLkiG+kM1+oxe+VCufjIz7VAQBPv8CatzN
1/KIwrBpv0WPdpwGu8U2xhOcYsYDIV2+cW795EWcfpWVy1wW8lP4lDGhmo4p/kWz
HANZ2upP4gRZM01CG2HEYhGlI3ZJU6X0QzDzoZHPBGCbjKIqkt3iBBy0aoJfV5mF
60eOJ4XErQ720gG1DHEVTIf8C84QWo8Zap9zkLYchBjZok5Q/7P2wamKs3jShUrA
q0IMtnLYiPggoxjjfbWbMm9/7P5bjOf3tpE51wkHWGEdZRlA0UriTBv+pED46xxl
OtLTR0WKG7zC5rVNUx83Bl6UAFEWPzIX4bwJNJJXQzZU6d3SnfKEPVBeUmtwRK36
cD1oh7K9g0icJJtQxulFB702y6Rsy7wDB9hOLZBHXiWFAa7d2ScyuW0nYIjPSSDL
xsx/p+LjTi2qGOgv1QEKc+ihRDFDLKH3DiFjfBQ3qpaAJxGldAsSFesHH5NuzF1F
p0oOEd1RqGjDPcRbc+aKthMENIwcRrQX39CoCjoMwQ/Y06tyMLYIOhpleNpnddpR
vMHXZ41Z1SHMpVb36je8ejyNz7tURu7XspHIJY6GmtflcUwrw5kHuwBJC9ynEww8
DYJlq9blkV5lxXjDsfJOrLsr6FBjUwCBkmnnVdJO6Kujt9KiK4X9FzW16CPF/qzX
3yvAsLuK/8EH6miENee70576khBXlhtDiaT+NhAHfaemwW5oT6h5IIZmCLBE9frc
bEe4SwUyHtp04NNAr+i9LxI0lGwjDEoozdTfkNGyA7FJ2ZnlKc00/Bu3kcfDBmDL
zFuf2v+v7vQ28tVMz3ZAaLNukz8MOsZzqJH8RLNhqUeMoBEoQK7XcWgBO0PZ1xu3
DX3j/dwnVRFnXr0jADroNR07u2vYq6YpX8Bd2e9CeTWNylvfVMq0ceLCPN5GQAKS
6M26Qz1/A1gf7fLfjJiM4PMoKAmfwZQo8CgM/HcfP1Yf6namvpLd8wu1DytQhqP8
sRI2ayN2vibvh25Hyp6jPeIn1IF/DD/BU2MGAG0BekW37biJipWYPPWl0ykjbjXi
Wlf6To8ZtVEJhxUG0S3XSdvDv3r0YD6J78eljTH/gg5S2hriFYoLZzwG8n6Iwlca
eWhnz9ESGRTR8XwKqFeuJ1dm3qwEFIg2xOo8S299ngGOFoVwYn92y5x8YzDa7JL+
0nHL2yLruZV4LZwgnD98ZY9VgHd20be/PKVvotRLLW8JbElORekdT7Y0nOSx+ldp
+9TheSb/OPIDAOFCDVZoWOvLvOubFSi7lOg+Om0kMdZuy6FoGv2AkSJS1rvFGN5e
uAxrqsEMwfNgO+Sfz8vElQuAGVjFo+etdGPQrF9TV+mcT73oAA6xgZLwdif0jY/y
TAO4o6xhiuVc7VrY05Sa86QaXkptyyv2m6rNAzlBohRajX/63XOH3xng47uOSN3p
tHeLzQ9aIUIfCH651cw27E+dvu5zkSHBgBqAUF9jrOZYpU5EhaPLCOan2/7ylgIw
CqDd0jPDZSoPYvxdO8prJKdGU/rwGvMlB5tESAYU2xh9EZDoa8MVQ2OK6JixUvHh
saMEft0HG2MHn4RODEf17GR9eSNwG9QmZZWMvhCupdMyGdp/o3O+I7KegFRn8D7g
sVl0gt6d80HQERMmBBkuoCvirooQXV5P6Y2hK1F9FzOKRZK4vPWg4vuyr6qIRIxv
OiQsnGiXmMn9j8pt1VL7SiBr1Spdug0H+kcwCF69HAX58XwefKMDeEk75nMEa8Bh
BQpd/r1RPORO5pUCJ25PpUPORzgtadA6tI2yNMnSmlyHkvYcz23weU8r8NgNDk64
S29WdH7C8/gEvbYBeBcAyCEAr4X/qrmjsbtKPNXWLlEjUCeZ6NN49ne+dl4Z2Mhf
TP7iQJoKJUQn2xHzDkslSL/75piKw2N8vkAWkVeamDzDbKXRE18tePltvoHgfWid
qWsTlT7ofrpGb128Kvg4dG9Jfku47xcWK96yEAzs9x/Qvql4SZmFUf0IXx0ce8/b
sB/4QSaU5/EcMTVRq7gIB2pJpRzp3xlRjLBZsEN6oFcs/cqHtuTSDxdgANWSpDl4
EqLe8SxLdSRMpEiSWPnS6VbNDzJkG46cxCZ3MxKTXpnERBoh+EgLJonMQGbBls4z
F3QjjhB3Bxe1AAWwcrRei8NmZ1e32cmXRM4hrlPZ78XXoZiNc2QiP6X1Re7oAvew
z63dJ3fcrLdKlzcSwlwZnVRG8f2lREXCyw80SdvvA2URi8dGnLPoph6POs0kgxuQ
6qAu9ALpxb07fl76lTVpvnB+Qw3STWKQKLpv8lo11I9Ba0QwCWzS60rVh4kN3zGv
UQ2LMTyeB8omqxsQpK9nY6EWN8TUAVhe+QfYlZqq8IaRiVkbJMz0ndOE6D9m6yI1
5uGpk8/8jDweTLwFSVj7eGhB9tJNxjWk9XgACWSDVAXHxF4FTySGVq2LmSMVUaPR
Tl+b5ANIBiHCKfaM3OcFMAGoYxEH1VL6QaGDDk7VFru6othjjEjquCYy7/VjzEoD
SM8a9m0shFPdjbBh6qg9tj8tFolkMfXlWMKi4nuRXhrjpgyLOdsDj30fQtsFeFky
iRrKvjabBA++qKmPc7xbtrJtDTq/crrajgcxoFjCQiVQbjIT4Q2f25WFvKbdf3dl
DWqgj6PgGTNGHx2MnH43AMVY23EYZ2qUNZgGP6Ay6kDTPwV72pzhdw9b2vt4G3qC
Qar3Hw8mYgH33mEVOcWeT0N80gwYDKBxsgTCdG1loHyYqWnLnBkkWiopU7puHSGs
bujpWonq4+9Js5z9BAh5+rMueoAutTBtRlfvX4APh/JcUqYbNoRhJWAlFoHi2rxH
IIGsAbvYc3m4GGlwTxoV69917Imi5ewQNOlxCPsBcVa+Q7Ud6nZx8xDZiTsvqJUN
REIvJ/cMOD9fXStj0x8SL/VO5c2i2QNEfpa3Q9CGu0eXlTGR6iKY51ImW0DXum4Y
HjxIw/Zb/djBQnCnVSipUD17oky9WPNkdrbBWoJLdJhfn+Pye71RnRqsFrnnaFe3
6rlQ+S0xoz606vFbaW25/7uRHk/lsQSQ6tSM2GdHTYP/z39Jr4yJ3ntcWX0ArKEd
JngFaTe7viz2t3WH7VNRGHb9B3q15nUd2pdtX82JuXm5YQjr5O3rQ1yjP87qLNzl
0/92gkzNfRZRhtc09ao95if1+xWqe0qGbx7v+Q4/T9pW6h14++uQVgo2B9UppuY3
HM81YagjuPePghOd1U4Wqzto1l4te/v6WxncPVPz64NKNctSgDYP1CzbeDl4g8k1
5jD1jYiD/5a3fC7/mMm4/OhQTv85qySW4ttqN6x9uYulD0bwznIzMyWlTKiDPdd0
/a67+nwHeXJTyqY7ggDcYRX3nIVXVQJ4MNHyz+xWRwoToJwvDAu9rUxapQJYhywz
OewsykOVgkby86mXNEOUMHVXpqByy7Kj/5XvZDyESqQIwtmUezs4uHlEfioDSMY5
li4ew57fc178U/aVSue/PHdTgfzbMuSkXTLtHLkvXWSmUPyeqUWrpnez/af99NzE
nANWXYKSkdbCE96YRaA7oKGq79S71cUhMlARsr+sBuNKY28/VCE6s1cMvFBrrEI5
bUIVJlVsNT8DqZ37Z1WKWrvSo5pIdZWcbD2kaBeXnk3n2A9vUsfhho9M4YkvrfB1
hcs7OTfcbopqqL47Zrde7h4zr5irDsqEHSt1b2nkUy6/Z17tzYvjbyyoQeBhJuyj
eFyexWkk+iTIRuX4RY3k6X3jPoQaHBVRAPOIAmld+UVrx/SLF9NZ6fuspE2iCC9b
rt1JxjtAwWXHMXdluFIcfsxLdQhrCXiZ+LRyajD+xLW/ElgVPIXo5dbdKKlpw7XS
AJSomyZBawLh5gJoGiT4ZO542QHNZm1HY+kwRUMpW0Q+jJ5SamN2UytQiCcFi5kT
nR1NnJ8HgQ75QBIOlpDr+sH7QbpFCQZJ8UL5oct4C4oQFqfBEtRjMejUIAjXnKee
/IXt8j4sNllQdY5QgMj1cwKSeeQah2zoF1fQEJ/7zx0K706NGR6U1W15VaGcXak1
TOhteV8KmptEazb542wL1hZD+950oqAuA0gK9fty1gLiFl8bk+L9ZjeRnRxWTy+U
zy6d2N/eIkjNP1UDYr6wripuMNeIW/HZo9rS2xvuCUYaCdkWiEZgDWSSAByHmhkn
+rDqKIJHFpxucPJ4u5LwqUOYSC5ItAVCfHpxQhKfbMCgRpK5++TNfj/Z+52y1Ahn
h7fOvxrN77QiPUD2vyCN+ieGuTevEWQxWzBcsDMtqNPvtkAZvvQLdv8FZJZPYD4l
QCP9TtUAU/3rotYHzI6cXH9u6w8taObyamoYuYSTSq+XqmIwbvUtqT3suRh8r9/P
KWyuusaAVcxHVz+MQmpNvblx+lSnPdspYI12Y9p6kbjS2vsHD68h31rO2Yhn49lG
lB8ZxgTZ6LdLP8joFjoNPs8ieBnNcXElpArGtgbuxaxTCpicAi29wFXsdVdmXzct
sVQuiPpz8O9uFz6/B2AVQDOVg2npf+VpHRNvKj+yDGoqKovctIibHoOI6Awncste
+3phzJhsbjOFBrx9OhAAf56nq6ECxRx3RS2LZZPe4rvf/uv9S+VBptZ3hg/aksFw
UnHi1RRi6wHAcS1LOyIWzqu6pOk6RTXruxPloDKz2xK2AQ2eMUsVHMVGozmd/Ro8
5XPI8yMU/CX9p+HD4T7TpxJN1foH0OaFRUMBFc10eKvkA1LQtxLWaM7zRh1o6lFI
mTMPDx3GpLf+9n8OWR/vrl3qDrxP2d6cBzYS5sTpogoFzvW7aW5tl0OdEx5Utfv0
X7msnfQWEEyBLwRX3GYMrK0B0aHgQNrWnbuPvoYRX68Cx/BSYS/2nSucPy19KpJK
z6pUKCXIlQvEuiTd0Uv04Z1L6RlUxJURDLYbQjxsemK+h79s0dhsV8P1P8HCdBfJ
vvSAF3/GWh+O+bCAFkELB9EYLfw48ffk71OyZUTGDKIMIJy868/Pqerkw9u0Ga7Q
JiQA6BbPmTFNQZQRN9c/ukC7QvfY/wS4sMlJS+qhIJ0zv8ZR0IGR2Os+0kRedZig
rXHI9/OGuDFxCuNPqSgr9VluhHVWszl3jMwb7BsqFGKNDR28gSJVwIkakCLTjtFP
7kdn97f98ie0isF/us1kLUB5GXEs7CRPPLoLT/ZYvS1xasCdV0RGctXIbuuesQRM
DOeZeMqLMPZvmdCfBr+ZuaOjkmbAkcxTm2ANXp51QUt0vBKTIUmVC58e9uP9h8RM
tMQ9YetbTxDjwzedX3pQZmB2mTHkSNCqM3bF8XX9E2cFW08F7+BBLXSdE3P9nILK
D1G09z4j9J6+tIzjDWCbLmYxcvnAVEC0qtN2iasI2iKJOcqEgbStieeOmGHoLATb
NL+JSaJivxZlwWEBkKcWWYEusKN4xEhQJ/hzUIfwaZjRZBtvCTJvQatiydWyhSfF
luIH1bViJ+dyMCQk31LQPiT6au3soKc2Py6tTbOioHSXZCqOK4wwyE6hHoS3wrHe
uxSDBcNA9NOF+l9g3i2mEhElT7bBBt0U4MO5gDmCm+q1vHAZEzJ/oxGMtTXNRGdg
moT3JrmM+RH4eOCOy3eIBhcbaBuUNB2iJFuFNsjJiqjzKxNm8baacEy6ntUJ9UHD
7mschjkwdxVVsJmytjQRYCf3bNglaNvzU7NSXa4joBjxfcUau0PkclMIxiqTGMGy
oxkX1QsrBEiHqmswYPUh6cbxoCNO33fKggcyY1Xkx3HdHr/Te7r4l1PJUqPmQKUL
Bw2QvovnPolHjjR5mKS+PQNTtz1uK22y+fGXQmfk6FYkLPFWFoBaDPQqmKFg1C41
nex3zjzXRjNPw6/CM5BBd8rOr2RvWivA+F8JfjGB0811Jnab2rVKV89OK+oS+O2a
9M5FOXexAUzxvU0vzQiWDVBo9mCglpb86/Mh6VfO7v1UKJIjocmbEtJmL33BIenp
YXwAbf8E9GpLkX9iXTloQkLfvJaGcxunkdNAEgqzt8Sp0dju0XaXK8rvbnM7QS1v
BVuJNoyUamh+f4Ha8iNTQieDGh0COVLV1zmYVPoe0Z6Me3WMV4KvjE02Sd1gwLV3
zt8KBzu2dVJrGcxWotvz4QkLUjbfbO70wFC0mLoDd42rOYsXtS0+Mm3CKjZA1Y02
yMBSJyi2iy38/UwqUtfZQzb3pwptabZAEXwS/rfBMOEnQj8cnk9n5dSATKK15nE+
js3ZLQCfbZHcrtTESkh26UeoGk5MzBlcq/Etm+ujMT4/m7YUrwOleCCYzQ9ltq52
D8+heEmBLth/BBxqZx1GfyEf8J95avM48NjoMEg4BbVzrV4ywJJoT9OGZ/ozg1ZN
0MokFa4qSaaBM1ITFCjaO27X8xrZquEAI2v7NXOcsYi7x8TKDLDEGtwD3IF8uZjA
ck0wyx2LVQwJtK+eCTbjujMgN+JWg06QfRw1Vci8CucdmW+KGze6KW2o2Q6/jCnl
ykZwP1pA4Z9xSQUHc6o/pxoFSPu3RAXVHUgUzINfkv9/zahRlA8pWV/6uM9DmMUW
bSfGOrwjWomywfzHPGupF+ijK2AW1V6vV0wRt/mjjGc+6fA38mkDy6CtXeXy7mkE
qNIoeRbruZOumarqag7wbPu4ypSBGH6C8zSflAap5r9ImDK3Qw9vKd+X8krHWENM
P+U71aev8RUMi8wNjoqzHa1Ia3Ooqzk8+nlXuh7JI8yCf87nwHT2QuV4Y2yhtv5S
Vy/uSZsjVZaxdBltElAZM4b+WC6TtMxs8Co57o+tXOsik6dihBMsLLPjXmWIa4R8
RDffsDD6++iQbVVJ+TuySNwEBOY8Lu/ThxS9eDwQpPR8uy4J4xlJWDD2Byn/IXtX
d6n50+DHTdOj/ZDsJInmSOoUqrE+kDeqEG5FQDhiET5491RcFydslrKR59MYf1t6
XfCBc4XmlUP80qJr2N5J93PDBFkFixeHraX2xAgJzB5nhWbJ7YyqPlwsu6606pnF
FS8TPVkYMWCKBBZhr2OmQY7DwC6FlpAgDbYqHOiZzpeKsw2rkX8Ab1TnkacnPmQB
viTalt5Avo9wofZMSlPqsqZDO2j58grnNpCNK82KYuk9m0TDVTk6SZ0nVx0NlNQF
vCXnKzsnTEXrP9DiQMnc63KwKp4yQQZCmNEQvVKOtvTpvmQCUktW361yCF0fWovj
yRm2ZlkmKwS+7APggK+/tOz64B7St1D89XFTsBZHoY+KvFdlm8WruZvkiF9i7VMV
NB6euIH7UuPSNahU9vnQU4OveAZqilrKKze5+lemQRWIjpH79mpVc+Mw17vGRuBy
R4XUcklnFJwUBlGFwA7I80Th8QZnycHHSqg7mMKPM2Y32tTxDE4v03y6+68nce/3
IZtBu9L40ZCBHm3xBSsoDYDtdnMKXxEbGhG1pfpJbh2FFx5H4FR4zfRu1PDFe//Y
IhMEOS0dWvjIcqpjdH0Wqx70/JAYYNCq1Y16SZHd3OFW99/bMu0GnctH2qtbUhur
ztpgEk3R1EyntSoOZmedYL+Q80Z3lOp4+WTP3N1RJnFO28xmDvM3Ct5fJVSxfpjC
bEtCOw9prbVAO/ayzgOxMTQJZEgkjlS7ow/TR2js/4dixSBu0HeEdVcN8+LY0Q8r
ZMZSkeFPFYG4oo+CYTHmb48NMRnG7+3hJzNHorfnUNsG3DqIIM8hwuA2vDM1jtai
w68U2++R+OLSA1x/s6h0uWB1hXQKIb4QdQH6aUZ56UBCKDF0SuZE+nxYLgTOkfUP
/qkKeOewHdTRhCzRPYf1nI9uxNrCiQvBITvIsc+IwUXOUA6OR0gY8L18ol9fMgXF
IkhuisnWt/XTW07x2eKRL0Q5/7bwYBSQ10mT89IGdeSzvVMdzPDtVJQGYsUOPe1r
VNm/+Yt/3J8zjP09vXmaWsw7ZQBNN0S9b6J7BvMBTtGW73hNpH0it8RLET1BhS5K
MLPxCwTjoxRByvMz+wt+JU0W4G25ZX6S4Z5jnvV6f+a16TP3GVKlN7Mx9256JqrJ
hZmltUlMoWpAWB0HwIWuecxhuhayGqt8GBwZ/+4pKzYZLzHpjmbLuGcSZxLJ/hjq
jSPdpZqXp3EWL1v7d99oDWJPW9wnptmu0oAb9fi/dSebExp3cytOOsS0+HxN+xgS
+NYrnx2g8o0LYD2zhxDdV0EMyelJhCFAzl0Y2dVa4fy+cr+j0zBvwruMJqn1S5Ug
nrXfvWNX/7vOHyyNtTUjzRLdwkmgYr7U2Sa5Ype4UR67QvkmyID+R5R0bkWCx9lY
8QibZXiBw7PpjHdN15DhbtJphqX/sVmJjdWJv4xKNWwR/ad88djpLQM7EHqndGYG
XIpvEXwfFEQfCziaFac+besRh+orvT1hirMn+slu4N/CW8pb2SzWtYgOuarNM1PG
TXDNfLmzM7lDFBugEXCoU8iVsSWeIgEEdwgWz2UHEnfLB9nw0v/iIx1mNc920tJ8
QPIUn3KWLnCMNyR4AB2JC0hTBgFhDMtYNv/w0a3iONYh8KIDZHONrt04uKrv/OYD
iV6Kdoop5M4K4Y/JC8wgGXQInsyvIeccbNR3I473UblkLIhgg9Jk2od+hyiMB9ip
ETL2Cd3kDdP28KxLufTzlzmld0gkqhwHZrIaaFXCx8aJAV2QcHIq/hzvCKSk0i6v
Pn3RnOy3BitVaK/Nupcf7S7NcElqh6N/YM8tDnoxqB4vQB5Wq4DE8M3i8bsmCBqI
ywuvTYyrAHkSw07S79JYZ+ahaCIkcnsedh7Mjv8ReTzaYA1RoxzjWboXaGCMX+Ul
0KPSvEuAfG+Wd7wcj/R7X1bD1Zyhtw2uNjCsBafCXQumrnBQE2btOiKGHGNSamr/
ZSJNiObngRWNGJj2ZkHhr+txwhpemomiilAbe43x5isaCg3fSdoLWKQfUJS/MlAX
NZWHL6oi4qsKk5ArzklwMj6ZjMZH++lzXhxJ+L2CKAhZYYt0Fu3H/PAtr1r6ndl2
EtH1P9yAjW98yQrLVjFcFmVq3+LM1BbN64h+4X2AsJB+I4tS7kW2V5fdr634hGbC
pZI3nthS13pmvVHPbcCEhHPfg7jrhhlnTFhJvOuFw6tuR7JTILh2q5d4lbtrrsl3
yxNkSToChJjKHwtuBvHAaSf0Fhz7cD7UyjEHogDPJKVPScTizTG4wd1Zi9IsZ+h7
REWM1ZSsaTP7Vloiu3iexyb0s9tvb0G2AvpPtBx3ZNuCh1adpuNDQrx5/TC9EMe8
N+acm6pgaoJAuVMnfPr7lZeeqscrSFpOINvoUMo/ZILO1PjAKhUVdeP1ShBTslBE
smfCEvaE0rNYGq6wOno8WGM9WVUjWDn3QYzV23eH80O0EhcYtaoIes18KxjVJbPj
RAOCoGFBwgqzqx8pDtTexPd73WNOdQHwIQuLna4MOfvCbTA3hFUkPnUnc3neI5v5
5pYTHhBGgYfYlB3X8NE2x2phtLo/DxQFbjG2F2m35WMGcTACRSDzyplAZNUiLMai
IrV88TwRLiUpPOkMZbnJpadV9m10JiAKTySwdy3RBfEoTbx3zRp18nfslxPfzVBI
Lz/g897KSkZzDBzBFlOiEySlHlHv1KnpuKnQLg6VD7MrQfdYixcOFEF5O8KJhzEa
br5Y20YEQaa/eQuWcSYG06UQhF+4zKaf7JXVOOHS/8KSbg6VlMKbj8re9UZKoyRe
3985gwp0MAdtX7s3fQAwq1Tf+c+pbrA/lT9+QpzXbJ7NzyeWn7aPlXJkalnwW/gy
z0eW4T2wrVr2pg+NaXj3XwWIzgde+ksjoyeVtg0aah5Z95xwg0Yg5ebI5Oq0vv2T
Zm+VSuGSxAtHnyzujWMSxtIWRgaKmjDnOPpX0UGp3vPS2umVhYA9ty7QzbF8VSVj
3PSgpEY+m9bO8YdjeMQyVKgfL5va1QYpoFipHziTQ44HacV3WksmzP1xS5041ZXS
lP0crcX6erANCzXYSLaZ+Hp34M8gzjZ4CwbrOZmrGnDK4FZLErgi441/oywAEmF3
RP/1NcnX6VauR/gt0HlmRqeWlMcFaxtV3tszV6OCuY/GZsxnRAnxWcW9ZjwjH1di
Z7zLZiHClJF/z9q+OpThoYNgwbuKMdUc7hUATBfZDmkgz8J5J/F2y4QHZlfUcFgN
S1rVdr62LcX9ey2SYFjW887zA1pw1BkJlJkcN0NTzV5vDyNObKW/N7129r/jBgzv
TKbM6TCqY6flAYrL88MltTdwo40KAvRYloUtRb7oL6A8rX9Db94+JhtIGb0HVC9E
k/22uiZqYIer18GMX3RRVMd3Ai5bGUmvWqvo5zbDjPLq5CfRF32+pcf7iF8LneL5
dO6sIPMrg7kGSqx0Hj4JzPFCfLot3FBN6ICcnvgTFl7dr0JeRKcQVrs5LNx5xPQR
Hp3jlPGKaH0eucDaDNFn7peQRlnCUl9gZkqZ8+U+FnG3Cgh4zPGFtYgH9QN5iRgg
CunJQs0bW2sUzw3rHv2ggWpo4ecAaywG5JU90CenF3m/OrjQzWFNUKul5D/GpWBo
k5q54Z+0XmsFKaNAoKb6at2864ZUrO2lkM/QE9pcaU9hJaSfSKLnrsl5/8cQkbVU
O2bWgVwdXgUKfdMOEUSNw7w1F99b9Vc02rhbVPZHbOV9YMtBV6HLO9/7fjw6Rc7E
slbBcZH9SKTU64PKNN3vewnclHm6EoRLcfdR+UF+7yBxkaKtGhtd5UFMARv4yL9V
yRSFV/jIRfiTa1qAy/0yxAfduOxEGa/9nTLE0Kb6l5+sIPpP2jcbQg7ccEyd5n3z
h0iFTGo5Sdu/JlOL0dgDrlRm6Aq4dmBOjK2Gg/eUS3fQmLjzZshET7mhmYUDx+iU
fWABjhVVmDbta6rWUlo6aTcoHfE8In7Yf5XrepislJdFw6lqwoJ5YE/UKHYaJLgM
E1OJ7c5cSQ6eYGVmV0B1SeBW0WFpenm0NtF8DF/sDTwWi6CCwfmY5kEojYNZrMFw
z6eYYaNSMfcsZsVDPxnPjwUPW9OswwwCkPSNKXbNf8NVcag8PwMfw7cqOCJ5psrm
IvdlKwgEoYnmlKP5lMhdxvpgrg53WukWWSYVsiMFsYhZz4uLXDKQt744ybOAcAzC
EsiDSLd/FGGqnSOeRfDDYNTcfVENHx/Ju5oE2dKDYdxQ1s2pDVEkR7yqz7iFQa19
MND4v1fWTJAkrp73koKV70k/gS/T3B93Wsj0QQWlV11FY+I1HMKsEuWlOr95eJDP
RFeWAq0IFathCqS3oA41ixk4ON05qkaF0+pRPemOghFFtdfILf8ejSn5/RFj/12w
rBP0pVGnU21+sWR2WadPfrIaUuYJbNalWx5fkOjPrsub2x0kpiUf6tuYrX4vYP4R
eiDrUZeeRYk9H1/hKsLGYNzxjEn8mv4Ah7LmJPSaD2GvFBC1aKZFkHYlXZyuKD3d
9VOFhkM3BzZoAx6PAoWHCJLsTMBwZ9aj6m33UrczGxIE1ROYu+CLjl874T0yCih6
SwWOXv5S9UAgwbixbQXfPNzMfPY59d2hizu4fES6Ry2/srfwpaavUvo01AN5Z49T
XcnUY4bwfTIURca0WNAY4Xocu1COIVzHMrV6fvGiYL1/7OhbHnSnTSKpk/ewxOtS
hgYT1JFaQC4d4+rrYP+2/3m9dKl8uzxJ2DCfE3+W98f65oUkou1w+QRcyzgr6WbT
G1S3XxsWil+YG4XEuwt5E0fLD7ls8XIax8cop2mMQPdpdmmkPAqvkSv0xEE/opmN
/C9ICjBClcpdC/LDWHxfzXKPc+5rKcuISt367M6qwz1Oj6JNZY8EOSX9zecG0F40
OnlI5L56tVVQhUxtX0p8EVHmpH/UkBy5m4Wr6401mnvjC/JpqsaNpQHoHse+eNer
pmnPCPGCkCfa/assBoCtPiQDxH9zWKVgDstKQEJ9PDIJMwFTSDltbOOXByp/MF+j
mH+X5B5gCSDVAb3clPFAWc883cQtRXmavHdl7AxX/ElvhAUlXLl41MjdzSnXuFgI
fVHkIkMjRK7F6jLM+jiWU8KsQMjKjjBnyFGtLvgoR7nrEJR+dtKkFGPFH7cXuPt2
Boi63EWQFLhs5Sze3KyiSkHCmoDCD/NoNBjRJsyOLur5x1QbHdLuVCpJMubVgT3U
8ZSR4/J1bpdAeUkV5R3ps5D3TDFWcJka85GAzlt0H7BWzPtrgZIuEmBdoxK/fIBs
u/9Np8pWKH9gzv9TvhO1kwMPzDxG/vLoe9UKJ1bNsJ35+McFohU8lkhPVp7A0HOq
4jMDMEUBDmYBlA4tlxmXdN0ymM+bFedbFGDatF2oxFJM1joqqg2yMM+zfoRi01vZ
tboLQJqm1WOD20USJLmZjQ==
`pragma protect end_protected
