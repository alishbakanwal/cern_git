// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:05:30 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
WsHWhWOnuJ2h24PKeew0z86CHom8Kqq64hoI6+RD0WEF2afbpEJKZFV7HUnnqmEh
NcmmSreI+OdvjQrw00Qn2XPpAd9YfoO8U7DVPowOOP3jC44FLD9oGryB2+P5GKUl
Jj3AZ0qySH8fEFQiCSgDewxYGU0TRQ20rIkabVoxqYU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 71408)
MwNQd8bSPFKKZFoCAWotDwYHE+DGguxw5JgTQ+cg49r7chCNCm9YVrgyi+oi2a34
/sNLSpi/hL3MilSnmiv/awGAZJKzC8SQ+iMk7touHbGvEZUZBmENJ1+I4S+gt3g1
9A2O9WZjeaTJOmHhoxJIupT8J3mPofiA3cMc7z5F3adxctStwltOjRYr1dwi3Sg4
iebLbCTvj5DGLP/WXsh9Ndzfb24M5Rwmhd29kSIjnkB+JClHcix32La1oou99bYi
rUtj4YRbUm2ap2j8TtmZ2rBj8M/f48lVNW3K/hMKM27afpEJinaqPS5K8e18GEZ0
KGyA4n5wjz4RRn2ZM3K7rRYKha0tZyHad6svrSpS+Jt1N+QnDMx9F+8bqHq0iBDa
1JjWU7CTrZUmh+iKmdRrT5JY3MrTfP8tVSCKazAB4pW4OCv8/UWyOT004pP5y+5a
Cil6ZJ0P0XB8AEyqhFS4vnf5FAacKEVApp7AbfO8pZUGgrwDF2NC9YJA+zN71Sg1
fTqm8b+EyT2ZBb1bORCcvMWCro2NT7sgODqB1flyjJw1pIw31McTLhceO60eph8H
669ixjjQHnBam2hsWTM9YoSDjenhgCIk5Fv+VczQ26+QCNkiLDulNJbQifBSiQdN
zSariQWPqxaPelGQ9g8jhP90ixnuOQouo7+whvoYuIwa+53V2rqTs2AQv6vhcbDc
lGzH4HnGFtUJllKM2oh8Anqvnxv1sBEJP4ZMww/ZiGLWuwwGyNkuKU5K+6PRkKOA
LzR5MuRUYwbTsNBvRyIQ2vgAcyIbVkgIZpu+w+pgkd2VSFafwqH08suPsw5VgTLz
miKFHt6BtvarJUt2nhdh9z4hfPScEHSjsYgx08Hit7HcpHLdti+/Lp7FkV3wafw/
NTNDnXCUTSYLo7nd1xmFHP5tv37rvv/wCQJnpkOJ+eJKKjyyHeqgqI4FjH6PWWi5
dlsKxpJU5IDgFXDelXErTsrMeO1xDUTrLH4t7KZmFYFwszPpiZDllqnbjFJWrg5i
WE6eYg1wAS3HXwWynl9TG1a1gbwvyo5Spcth2GJO4hBbhVn8gALQTvTRp88yWZDA
0UFmydVL1WmaDhW6HLqVtk86BqZVPhnMIrJ3gcv4sNdcWXoBgIo42l9I3sHbF4Dl
z131b8mdekIU+TbTVROnSrkd5khwq3xf2a/ZSPffHHsH0MWZBgLnWLiwDRCHNDg4
08zAiRzUWiAx1VNuSBmsK2D1DUMzT10s+PB/h7ctb7SZliReLxl3L+S8t+QDSmqK
d56tnws8G3U/TFw8gHR2xVvdxw0DrSXaPohC1uPiwtoBUcUfS2zu5HfgzWz4wiXe
qOZlmWRgdP4SFmowQLuSTLitaGQtvjdcDlwOHCb44bEPrl6XxRYNbyY3HajhmIoS
r7B0eKhTbK/HUSwRDgp/LCjT/n/NTS6l3slMv0YejY2Ou0loISXETvFQIlnSnKzO
3JaNA6Fn1IhxwrRC3r0WvLhRefa35ahXEG4stQ6sALaTcjCzfukT25xmD4igmNFL
EAu6UTZlIU7Vytg71jrFA/c5nMDkvhuqzwA8hOArqkW5eIbqPIbWtMwUGJZx4L08
oZFsY+CALOk2nlwMVyixSvpncEOuunuY/xZFkt8lQrBc39H9QrQucBFSyRXTbFWW
Y05VB3qum5HRkF38TmSxIyH42R2WQ/x3l+daU5A64rKlANFIQiXJG8gs5bRgzfY7
SVZlXQYoxkJ6Yz8T26VkWB2ofYlCOZjYAdOScMKX4O7MLTXHoS9hQKXnoXCyAZdM
dk0p/yfSxhu1RlC68yiZ0n499OFYBxh/c++sO/bJZm9amkn9QPW5oHnNBremHGBj
CRrlK2pEP3B8yikN5oQYQVYkYzabjxqmosGqcXjXzL7MJmn5D1XLah2pOLhfqGaO
7hhUfQa7Bk3OQikhTCHLJyRptaVoOgvB3nS5OVQVmMNjIjA62d0+v97YKImpSPKo
jTguTPAw4yMEqZDmldMMG0g8vClTTFMynIBiA5XJl+2QWev7F6KytT3k/BOOvhBN
W5guQBfvBeMXtB9ndd4oGxjxS2NPxF7udw0bqiIzZ9p2wI5vKDOQgZMrLQwfkvnL
PqalfOEUxvsHC9GFg8/pqqYAmOJJv5M6F2pVdxMBb8R8argBpBvvpLt/jlDG363O
beS57jzdFS8zoLHVckFFkReh/uP2+SgJ+t537NuaEFWV0zku4KR1V6wRG59cc1bF
3FE7oIn4SkNxjZZULw/lwkJ+EQ227n9ybdKP1r1pVXR6LIc0PqORX8FurkJUAud/
9Qh14uqLX7MewV+ODliyOFv0X5RpGcFyT8tZZ+i09fB8p1vfoifLHFW+A7ZhI8ko
k8M1m1fkP42SqzvNLVmT9jWN/j/NNj1JNd3ss+0SVNK0Nfgraegab4qLuACh56Pj
HL4eZNFO74C2tTfXLi3bg81qBDSf2tDSNUFLN3zAtLa5azMesPbYj0TBkcAwbc7a
25ZBxC/91zNQdBqO91+OtN8UdfihS39JnFtfEcJxn9L40RuYXXgYhwSO1TbBi9Rv
/D+6yKdqRN4i6ehKOs5S0ebY1capL2nZguQgaLiUgmS/g6s5wNe5P2y9qzv9Y8qZ
q/EDkduQs0xog9GlTTuDyq9J049I385rU4f3aPFGM8WoDQzp+6gIQ4h1T1po3pL9
5zugseG6kAvg8krF29hZBW0FdQZreQC0bIMJAuISMmGT4U+72nn03oDEOAeT007q
AILvWFS8WzVdtM5egVrq5Z+ClmpiYyph+hb4Cq2rIhF98LfFH5GrjONaAYdH7lPp
AUdrk/AQ+tZdmlVv3Uy8hMp0lZLdIfDUcklwii9Z7FBULfJvyo13D7cFi067unfv
jGgVGhhq7UViWEwpCi1phwjwJDEhb93BeimvB8ajiSJHkvbM97vS3g0oi3Su5eXg
cYceLNMviWacphnFJUbD9PpbdBDNqMviPqkr8vUwu8T94qZuytR7F4gNpiho4Zjm
6XVGsP+poIfGjD6PDQ9upUdD03jvC/0DUGIIM/H7hv9eXrs7KkekFshYIjV3Z4ss
D5sRdHaeablKr2xLmsml+MRWV2L4UWpxYu0EdA+5AiZyNuskmqB5yrs8RGyqmnHC
FZn/NOydX8WWIgpLZTibISmzq+wB1tOuDrmPKnv5T5pLXtaEytPBdZGBSJchqL2e
yABcDG2Df1efz2NBJDTgL05L1iXbNZwODrYeZ2FZ9W7ISKToB3EtRWtJfgNX0DcX
Juc4eCGmSxctFfxnGgsNhjc0h+dcGSODDnhDPg+EXPUVgTjGFGsjxtfbQGnd/T1W
rW72rXS1gN9VAqDsnJ7wOtTWJK+IaQMbkUj4aZsyK7DFZyqIBGT6r71DYKUA4Kvf
mYMfeC1kXAs/6KVLx+o17qhY3sbodme5WVAys1//cskmUBBgQ8sRXDKIFSpOQS4o
FBgqaBu7AxAoH0SKRjn2P3Wmw73JefWycTbS49bcowzUWjPHXTN7DHZzjq3Q1djJ
85ehQXibT0hPyL4JS/ctn+bUqbFYhSKJ8UoJ9IdYS2UNfxxXlBzyQviJIWlzFqpy
spD93KLeOm7q56ab8NTjK652F6ubujZcgkZH8kJ7tkHQGN46shmNKALvacLTvvyN
TBR3P1AE/qfYktDvt3qx4SBM2TW4CbiyDC2FR0NjmT+TJCTpZo/QSzfjr4h+ak99
4WLglvTmNu/HVFb9MF7owko/6V+t81EsZyL8QRqu40U1UrXKpCr8ZPKGS+Y8cKw0
X9t15Lixq3NqTpoloWCBENxpysQpixkmDP2jokn6V7y4+X1O8Z7h4Qn+CY/m8GZt
0hYU4rLNq3h3VPyDnuiPu/cqQy2+moE6ypyG7LAPTFoSiObGdUvNOLYbHwQEsmG8
H1HhM2SfyE/wdc/rFHIjTaZyEh6C7EoG+54ErVQYmBlgmNvMWy1oqX5QhO257x/g
2yr0xsG/N3MrrBFOXgjptgVyY39WZNRbnm7lovhI3NaRQPNPh9RrOhbS9oHGhJL4
okHOlb87FbctMZ2GMIkeEZ49H4mOw75u55iCU8R/nb+YZTVtf1k8vCalQbXBQPnC
hWNXXBNAQOQPuwHIZtfZEb6Qmx1uFB5UIrRWRqcIuArXzTyKbTbDMhizwR6fPrP4
Be3E8jyzz3/MDoRDDyOFXUBiSGHKnzORqGyALroe8oXPuk8qaE9PK5/BGfGEABqL
4oZ9okJDM8AtK5Zvs3NBPUqRtlO2boEGu/2Y9W3XWYIIFPxoH3ZaTVb5qUYdYBsH
O6QTtiZsqt+6jLZzY/15ZspGxX5xyXOpxbHqMEzZPZ3wkiWyIRTF0NMIpMQJ4WJI
ThK6JJHTDbYZpv2H2SV0XkneTlKLvryzDSxXG0WPle2ftLegkh+GGoPAOqtoOk2j
E5P1KozsoQt/bAG9AI1FERHgmM+fLKub85+0VpBTpYpG6J4f/fVaGAKzVeRHekVJ
lAfaimhWmVp9mwHKcuJ3couUkr35B0gH6Ad6Tj5q8kMMJFvAp7ayrROMp3gM+/rs
kiUSGQoj3GterBamT/6IhFawoNhdEDrMitz82ac6BpJZLiIqxDmOsqxcrkQRPpdR
KgHXX8UEB8pD7X9+TnIY2lMGuN8R1fVxuo8a9LHGuSH49v5PJ/clTRbE+T2F3tA/
Hp9FTpfLUgXj7RsN+WTMG1u3iymJdR9Hr+nbN49TMmKnUyYhtpP3fCqbhaGG3oCk
xEJ2zHZ0D1yl9usI1ISZgBCsdcNiLeHmrMNU2Xt7bbZVks9sd2kW1JZX0Jj++Or8
UGJtLHQyJdg5TuagKk0WPQsyI14RF7upjBq9AUYxhZa5OBst8jsGjdZZka8HLYSz
2W5yA/XZCNIbwk8TWqwreAcNyhyQOsIBRqB8lXiijmR3fKM+7w4fjHX1fJJaOSV+
wOy1RAwzn7LesUnchzPIOXu+GukWu564x8XW/+YR3ZDztyIH9EUmepcZ0OIefAFu
NwK5T9hid55BSb0R7ILRAosVy2IF1iqx0v6IYVzkT0ol1C2eB0ty1x1jqHMKOMYY
PaSjgsAu3LF0XLDdZ/o2bdBRB9RVSA4eLT6jPRsOkS4Bhmh5+le69Y3QFH7DoHUp
qHeR7LdJQVYbGozgTtRvGzqKMQ4dNoug/a2S/QiGdcUrAQC75Sl6wov88F54BlEj
8plB8bF4uLnD2gWgqlOIiTy41r+fnKSvlNVuP2kVxfcwh1ltxIVW4nV2VaQoX2qu
lLXrpJy1mdSZVMYBtI0a1gQjFFWiHelYite9Dz0B9uowCdLs8GUJ1pPi8DegOrkZ
utLkCTjVTBkVMqxL927phXYg7HOh8h81Wc5QqMleQ0EHUqJv80VZqrlrQ1t+sMzO
EV7kdiq/Vfz998WdO8SjS3k6rxg6J9dh7gIrHdSAH0oARc7sQo8cs0BTawvdJFaV
fHBPs9XfJgfFwlOnQPRtMaRkWtMMr52JVOxwRvJr1hMmatuV3h3lDYShMDdOMVtn
KOSAH9RiNlRyV2mRBWGetVZd+QrLCqIXq88891tdDmdIt3tu8bbrKsttnQaBFXZ1
/nCGZamHXvRc/kk02DV8+dhAaaSqzEEZEvD1w2X7qnLaihcXo9AYxeJdu0nO6qAh
m/R06CPJgkOCyhfKdvesHaPtnHKjaJaURPaM/Yp//wCyyM4rNCCFtR4xq+Nwcxel
sCVJg8ugZcdJWDmk6fIfCjuswPtlw3uKaiAOS8/A+PEpPIHGm7OligBIF9JAAEah
bpdZ/mftJEZfTi4WFVxmYnkebq8A/Kk20Twjaug+/HJ99jRBDRTduLr4CLK1j3sd
jajHj70Z6hE0cyvdAOc4IBtwYAIFh1EWkb25tt/2cXWDUZUQqX8835syd6kSzUOr
RyBDpeIrLx+dpuOwIb6xIHw3qYBCnGsgCzjjwXmfjcw68G8a5sCHgj+9+t2m9IPJ
T2bknBhQqXI1bw8Te3rKHf4bh8DNJo16YHFgEKAdQd7j509qWQXQfbo8zfNd6A8T
ihxq6Zim9yhhVbvqTPifpmqQHCpJUZTEqdIZyPM8IA4EPqhteqVa/1WikK9Unzj4
FDRk4pmr35jQQtUddJA7Esm3/DDUknVl7PtVrDCR++mzyWteRM6ZxMKgUoV88CPG
ybCOJHzNePI7T6lU6SJIUibTVOXLB+CQsprJBeElnBpyRR7XKlIzs3NFDYw3CHQj
EgPWUXbX8sglemX9B4I21c/Kfnt1Qn7SfjJ4H9RIUX/zjZfbso6t7Le7zGMNHiD4
AmWKmDSp2omigjs8wvKN/LQw5L4wcdLPibtEOaYIwfV+3MFabPDmtHk0JFaNHX5s
QmyOx4ENI6l4FVT3MpZr8hHQFtDivEs6RW1UnG03SkAq78uuSkU6vMr60hWu3o9k
y4kD5PRRBGez5W4tDv2oi++CrRS1fOKVrOzZX/uiXxdDl60JhMqROD4lPiXFw5MD
uNfkPyQ6b2DVMyQCR4pPvkLPd8WkL0NZzup2spw1jbE36gELAg/pVh41DGdhv72i
F4+oogZO64U9SIqf9nwpzuT8QZqfGDXRXhFn/SmfOGfngJhwippTpUbClo+Civae
GkB1a3686PhZVvAcT9muo7yvApKN3IsfMYSmixSXnhQuuGr+tLlmKLNA/jwgu9gD
KSjW7ZYZffiCWTPGwiwLMEoRAiij9YSh7FQZ/HiDl3+X2Mx3zrOonNrQcN6/W6y4
BXaiRsRdZVz+GX0Bj74c056aaxkTyXg6oxS83ZhqA7nJcqJeioQ5oKqgcVZc8MMd
aGxtHPwSXgrRSwWd9SqYH5sny+axRdCYOWMO49C0hNYNxpgS186LTjuTuD65tkSW
7MVZyqed9b/G1ufIU01hwEMCZpQO2oXOjg0rhwAV2J3lSeQEf+4kkT6P+HQa3B/6
TZzRImGpUrxTdeg6z5lObLFFEkcFscPgUhEfHfUFXM/Nj59TqX+gAUYmQKiTaHPw
kMeYQ89ohByBfnh/xOHRmTlOGl8oPEMWlDY1x+HVzCUTpdVpqiTHfDXf6Of6tX3A
0GUjhDxQPQWj75OAjFmjxgcvMQjk6uZoT1wtukN0nYuJaR+Y+J5zn8J3Bi4gAFw/
XHKtQhZ9v7o1FuA3jXh/kKyUtumOf0ZYc7NBMq+ke319T4b8JBhZI3wRBlqPB9tp
3/z7XKuXSw2PgX9EtfuM6lexobmFAWNpaYooDyu0N6oLltd8PhTsNT8PjRPxpWBi
dAFtGpzezhEM/QQmh7j5JqsoEgMCLJzekKMbPUkWyOfeU/tDxsN6ALQ5nbW6XTLG
g4tLQIY5bhyhXnR6sfItLDdmz316bum7t0zgvzlBI5z3wpypee52G3HzxmGCgVh+
PUZspPjOAs56TNZCjcMVvMUz0eaLkCRjhIyDiCX3F67Sl230Zk2ffBtc04+MrHjb
t5GqTDu79SBxEUiua8/PAGQY8nWQiLTY2pwCfCVFhcShWyh8GDs7gd1/WFl49kjv
BSaSA62D23uW+CQkZQ/ai9TWAgTZfUc7HTV0sw/WRm/Iwmx6tK5ztX6C2z6HVH2n
gY/KRlwQwJ93dMLmD5paFZWQXeubFOu++UG25VKdyaShETUBZiaE7iLDpA3PSLka
FY5N8E2sqVeV/L68MbuHamJfzrfJVYSNoXs0WAPvUHL/f6ohTQSK+oBZUfsuT2md
ALlSDJOc2LXYfCC7qjUIoXkxoEnBfzAWrGkTGjdsLK7cfA9DoY4logKE6sihSDRJ
umqV1xMHQhoeHeylIWJn+Bbxq0rDmxp3NYPYfhAl8pYJSwh7CmhBpQXR10aRxjzc
aXaONCSG5nhj17+o6O1Yk4G7pLJx0yF6nxh0RAm7il/+nlPKsIRsznIboMjt4+v+
sLiWngX4NDuJ3YVZPW0ZvZhD5TExJPDs+Fx6i/HDn4dnkoPKc8H9PrIb5bbTEux7
JCzvX1fk0Z+Nym5+IzNoq5C2V9X/0fYIdfU9Zzz87WsUs949G6FjVhtmmaVonxMk
gbmdep8n/fbjGCxsUCkZh6PCUdq9p5IZ7wALTz6hu1dBKfLDOZHXju1fKSaJHw5h
D5qgIf3aQxwyxZDXvLeOUuBlJuQxq8e5mn3CNoPVAgIN0YSPuTFJAxJx/fs78/Du
fhmoI9gGHNY46RiTdvl58hXituXbqIQ9zRbxebAzpHn0Xn4DCUMYZ1Zo8fOLmgVT
ew5k+xScI1C0IEWaTmAU5quOkb/Hy2POGJuneR7Ci6Ve4ULXguyMVf1UQgFZYZV6
twJb/E/LdsQcv1B21M42xG7547IwzVBfFS070O42b/m+vbLo0Ma/z8dUYPrWmpDd
W7GcStlG2qOpAjwtt1+X4lo11MjmU1y3SCFeWtaLYDlilno8WqcDTP4e0ib7/lHx
ZyctQ35tnYf38MvHZb1Q3fHRnPWr4UJKDASu+WEAMPuRlL+Z/2UL9y5Jb8y/IWFL
HHd3RPK8qKTChY4UYecNJUHiWlXCs9MBfBE9vTnvj/qoIAZGGv+QMYam6nPSSW+V
4vXqK6XxqG9dc3Z58KPX3bnJeFreDYdQiNjdlxCT3VNC137Xx2tko3EyIM0wnFRR
5Kw+X25++HWppkUyAreXZOjiSUhQn8owfiVRAUAWzTGexc2VSF0H5pgq5Nd12S+2
vNfzhDLn2m5mnmML7i3rCkKzcoNx6GhS4h+XoYxoknU1k7AbVPi7k0xW4mdPvp/4
oJgN3cuzacI1fhgVsj4nP6r9zivLTP5Th31Dyi1XUNS29gFHW8wCiZzI0o67k56o
b3lt0Tl81vMIZnsLWeP/zeUZv3sxiXelA5XSUXdJDn7YGWFK8Si/R0+mGn4YYkjA
bVjOzGACQXP3Yi7oq22cD4IpZgUQ7mfGjWRBAzVyabdT5tkRIGYwbHJNkcwzFD9q
UO79el/Lj9S2Wrv1hQEoXWK8RkLn/mr1ioO5O18d44YCsx/t6viF7XlsE2QVFW4W
p7g1iOHnRZREqKM5ya4hVp9QiDsrZxiotBuHRqHTI3n9AYoKcrxLff7BZbC/nset
qJ0GoCSwELJrXqBRjbcjwB8wzV5plRUBtG9pTIn8eABzwdeMktbMnKIg/kHZa+tV
HpFi6qrFY4tdjJsg7XcFL/if866j7gZRGSPiBsrRjMhMVIX3MERDty1eCzbbsa65
5946d3NtorKIgXXF978h1h4PhzXvin5d6Jryf+4BrmXNWoNIOEcVxyGWfvgNoTSm
Zuxr3TorKZSqGKyQ66Acm222RZBvd4Tw18w3eUmomjFkzv4DeahRpdpQ7TuJ6vFB
bd9W8ydcK0xXZbBIyFoZ/lPfBWgt0XOoSApyX9iXDK6AMLVtvPUycG26y7cxOBQh
tcB7ayYVNys9t62qUI3liOHgoGA5MtFBMP/BiiV5DBpR5uvCJLez7eYEaNmd9HCx
okkWgTdTPUdnWzbLBhmSoJmb4vnRtgbULRcOH3TK4RvNfu3hvS0HzLMRuLkw0HLh
BfS7IkK3jp78gRV58Uyjf4a3HCHEKnxWc4am3n5K6EL33VSArNetIWdwi9Td4AmQ
n4SecZhXwKiuBnCdKRB9zH97+8MQcXmEXd5SualrpxSTIepkh/d7HPo51FFv0rUd
SSE1XmGZxvGz1YP2HBSjWmqkMbjWU53TfYuQk7Nr3koRVLlTeppcj2DGUem4sEf2
5Gj/Y8hDzvt6kkCN6CArEW8SrAVDgXryLmgkLx/jBiJjPbrosD4XN3i5FVGzyqy0
5q4s4PoswCGMBePZg3JR0hcKrrKdRbPcWjLK9Lx2nCQeNn72FR1dN35dHofLmJRC
RyISeprfKGiAK2ryh1FU1sFwMDswm8un1KIPls6+QkvRtageStam/qc8wPninTJ9
HpYizg5nH9QIWWR2hINWorxyg8kVohp1+qk9R1F9sJD9cgSRDStjw0um5Xca4vUs
I4e6rGOqlE1bVIB0X8BVF3/esbMe1CDMAsw5RGqMUaX/1MiyJxYP+lR4p0pTjzS8
hrRt0ZHIPGnkFNLhl3XIeopFzCGVjrqWpwQS599niRyJd9khhJQiq/UjKgf/PdLz
qDlUECmtWip1S7uobn0j+f0uGvWUUb627S/U7lLUBAPse9JduoYtnbPc3uoB1KRB
YX+xPRxzg2knkjuf5+RD9oy+9WkYFnA6gbNtBgRCO4cDr2q/oPbwr+yfz0nBpB7l
7M+KAISP7vIM2H4Tgrysu9a1MneKobSdwePLah6Br13JSCkJ41shzUFnaK4bCO7E
JEnY+L/hKKjLrSvSHGtQU4+lDKrFqgeoV3T8UTMEPkR3WqKIQJOKL2Eg+1txvFoW
XI/oRZv3hdAd8O0k64w5cTMDq73w+WOEdRFiO9Nt1C4NUCb575nAEB/lwWwUem+I
Hk0YFY41ToYiTAMiCQGqqCZCv0B+LBbmlTGNuYMUXFjSMQuJMtftQQF5LywNjV6a
5+1AsNRSTK2OmN/g51kYKzcch9iz/QWgyXRsJKquRLxr9IZmMjf9mciIJLixizsb
OZ7lpK1d9OG/zI1eHoBkcgQX1IzSPREaqBRvxkL86r2I5sPtasF04ZTN7cbw2E8o
5ioXOpvc0jGko4MVKtRcNnsgTK0JUWJioRFwewS2A7VFhcoEDeeo816qlvs2qGbh
ThD3Hpq+eEFfzqldmaT6bHcCL/HY+tVxd04F+7SwnO3A0CMA+/dH0w7ol4TEBLv2
P5trfpI7yMwAcmatCdYifjBw5pVuiVy3GWVrwxH1hRGmzj3xxyeT6uN5VvW9A/Mp
7bJfy53RYJ/mrj5h0WE2cxaWuA8e/H95y/hNoqbthvEfSLGJ7/OiD/wJczlVoCqf
pUrmIrixj2rkAXuZqU8rns9vK/t9gxa9dyfEaHtKmKEsVi6+OTQBaCEur6WtKafj
lJqzMo5kySv+8TT/bZodrOyQqyaGzO13zNfpz28qdeF0V1EPRnKz/mgoSSKGhMzj
igA3q9N7r9xUtcvuoa2Lz9Y7gFcsL2dBnG9u6VLcZaX0a1nFpa9S3Th4gUFeJ2xd
C7rhz06UIOntYvQ8lqq2gNrSlMSSF5bSokDo8OusRPIaCEBnpWt9SCB0NkXikkxC
Nq0Ip0TAt3+0TEs+jkrApF65wIuSnG9McK8Zg2LE4U/DDgZ7AGXZB0zlD4H5vlST
GLgU4/mqsep17jzpXQk/RT2+ODY7SIoG0HbGLVXcy+FeRLASnQZGGEGtasG2hvqj
GZj08ajcMRD7kXXaQB7i8h4mdr31TRQNd7CRYisUsrh5+KwbI0bIgMOUU5eoCVfB
JPgxVxjvbJB8COKSj1r9fJEnLIpO9bXulFIwjexX9blJAgtbQvdDX8M7wkCBv7+P
QvhnaYL48Sk3GoOS2DSlx3gjaCmb103ZlPEvbRfa221UHCVhaF8VGsEFV2/Isodi
u/QnYt7jzux+VS7QUbjO4mO/ovPoIIkyIttdE2vnK8OzUe/DjeJqCeohFiT4KIol
JM57QmoOZe6gBiL30RUJvGY0jv/hEbFd3sdQw34WTgRpsCjbVqZ3kmi90M2Em9H7
ABoH0VgXXcagFrng8SirhNq9cyckMzMOs1mqPTqYRl8xmrNLxhzkM+V5K71TSMMh
xjtfORzoscEsS3RQSDJQx/G1KOYUomixHTuvDLif19aUJiApgdWJskdWk0u+ni1b
AgR4tPXeVrKUi0RjTql2QNwDSJiQM5OC11dLjGLk8SFq2Fkvfhn8F7AhcttetjBJ
DjKgUrjhy3gagjIDtTlqFdUyH38OKuVMvSZBrldL321/Iz4c67pu4+255c4pLIn4
Ka4wDO6zPRrp3oKlBEeiM72Mx0bhZuvXD10hjKdjrO8kKTdqoaG1ebZ0Hx6pSCYa
kKNsLhFk3qXvZVVwwvzayKEiA1fmHEofVEQD0r0EdCus4bLXmidrPhQOp4TSHpQl
SaRtxQJstSZcQ7VImmR1J2o9CO/rsCcAAvKtwi44F3BPOZmMWYXYr4fnFQqdHjUO
ZXyQW25neR9XlrfMVwdxzPaMWvd1bJ1e6meMAjcMDo0hr8r0mtFwvTfzUWZaq6GM
fLJqx1E1NqI8pzXtbdV62mBDSnhPumprX1tq71hFxT6haav43isCkfvqFNa7jObT
IYarQfXueWZXFT7Am9QbiK7Qn7JI+5TvY/nq9Lisins8cBo3nBN1qG0GuRmzOsgL
Z+ETDGx+JueJ+OLlgq7jy2vAq8rzDEqo2ypPc7FInuhWhQaoOnw4NvwoTJYYUOlK
aZ0BO7OQSKP9ZNGGEPo6XDtXAIOygLu6LuYoUT2tiRL7Mavi6Hajyiqd39oFSgPT
X3mX8Ha9VuiMh1O4NfcSS/EsQV/B8isMcGMWk2Zk5fZjYUKitItBjJ79jV5Q1Bhv
XIAx8S/QpVNIWn02Tpah4Cc+m6R3itFX21SPs7pRdCpLHKFc8Tsag2qXSscDZh7b
Wia1khimf5GVYfll2PAEG5MuAcAGC3v/1Rdg/+jgbbMTLU6x7SSXD0UuBSeSFoQh
1lD0K58TFBrL3YYWChKY2xu8KoM6SQRsWLO9GGbUidOSaJLimIeLHky7i5eJCBhx
iAMQ5w7S+bcxX6W0i1VlBZFRiCMRXGFDg90j96JLn05s7CGrT773/Fr2LJHqECxx
aOQRruAu05dPtcG8KgUWwLHqsSp6qDJUuPDOn6pQ8rO9CdtrCCjBSFxbmBJBHHkV
dKwNqmpJ+5iIcaccibUyMZmUAVlteRYmB6dvjyE1E7fuS2+9JM9CJedx43mZXSun
evMNmOvDelA93aA8n3etxyJNjFqwEIneBCip/yGDPl7ljyoW8PbjRKr4o0wHcAjr
k2YLZO02QQzfnZf0tapP6FmSPoW8CJ2q1WVenzPdqvQ4YbfghaTgYrik6mr9Owlo
/V5daciOlR2QO0crSfzEtzhf3FBiZMiMiAxmgmWtk9yn0mAJw5nRqbWvH5ahsgsU
XyxLiPDBzygRdy3kTIP1mdycwkigt9QyERcrC7H3Z8cGKR45ZHagBNXn9A3Eogt+
X8TVMiV89wjHjZHYfBnS5hsZmBA60APf/XsYSOkUt2tWekiGPi9Q51S3onQkwSSM
Glgig/ZFl091IVoYnyViIxvlABgardDiwS9apDXoDsHaJu7W3i0Q0tDhqrjOOeBc
swDag7N7p0v3zWn4d2hz66cVr28d2Ugw3Y4lA+MsRRZBs/Pxg4EcV1gaXtgEPXWE
ho6gKztv8G6gA8QFsKUXPHJNqKWTbr9zQS+C+yu83VEQUNI8qssxg3PDIgW8cQse
ZXR6darN75jBEKOPZzVI/oHBd471J53Pz73LN3hWJJgdCDeU0skhYtrIqs6BYlai
fE3pExSERpUks1//FTiYeObaiUwKkQgBv9jIcS17196/CV+rXQNqZN9MpzPfKDUR
B8k6eqkqaNAKXlL3QNSRbbUTeBFA0TIzRdFMqhHp1r9rhoInDaGEELBPhb2UxJ6h
NT9ObQvoxLYapg3v/F89IaCtp3kR/Yq48U67RE/GKv8WQJZk3eMrb1tjeTaIs2cP
vvRhUdHHrNt9YF9IMS9BUy5QnAaxmjjEiKIZyy58vE+pN4Gd1DvOinuAi+Y0O5Q3
Eb2Eui4zO1SKSUWGeUHz6f+UdE8jkYtHeGoL0lpTmk6GM1nrd032g2sXfkr7YyvS
IiByzDUhhhQ+3cvXJVUSjo/daJ7ZkLmxDogMc+whafjdj5BB8HOX/cUt/kefBmyD
BRDPty/dQl8NiS4Nm1BofQI2FoozP7+aj/SFTjnzJ8AD6p8j7/WUkUAuTuu3uncj
5vPZCcWcYp4jgYBvmOrONQsQ4l8XOOFY2dvwMa0P5XF4YP2pgTBeJ83JplxF6aU+
VIgqpc3pZ4QCq4+1/0CJLW1YwIVaAUqu+dOdujYhvnvPFQvVh7cfp9dowNhXnOnw
iGc48AdFSVK1M5L+pP2Y87sD2UdIcfse1XfriZgMSGBWZqMA/RfzUmkgP2zTlhAV
qtrXlqe3bhF1kpY8Z4vjO7WU4bI0j/aEB5dVqh2A4Z74vET1ysXge2XkidsJgRZf
sOJoM6BZWr4iNPnDWwCzkV2ZGe/sz410CEFssoMz5b7/x6vQsX5kLU3IjvOj0JeQ
GzOsdeAYZng/RuOzYl8E2xdTQrssvlGd37fLaFWTQj4PWFLOSI2+HQH+p/Rpdqqo
r7io5sSf1G8kTS+kaMknsxPyOT6m4cgh6OjqneBHplbHwrU9Wm9D7a8goJm3RYmu
0257AiaVzsC+ZFVn60wiujzVmkkmywxRw89ZavOZiis07NUWLCmUTWPfkh11FXsj
piopBqnURRDSG/TR8uXY6CWjgBib7bsJXFGNZ/83K6rPAxVVuIu056fAPOSuwFbZ
fe6zfEHMaB99aKo0a9N01ud03iq4fTXW4M+MxhVEQb9/FGTiN/TGreuONkyUdIRg
b4HTso6rJWHisEHxaurvPSNL3dbr+PtFLj9AKIgzdh1T420Vd/wWhxDcjgbt5mTF
luMlNYHSHRAKekDYuLiFRQII2mZlWKCdHzsG27krz8zrN/bA8oY0SwKQgO2vu22D
EcHcL9X+ByhHr4Z3I/EaoR7d2XzrDElPMQNeSCEuoDTKDr0I7ZVbpXHo+qS4ZreJ
wsiT4K5gutNAo4S7wpZNvPivJ53B6E2nbxuAyqetAhabQL0iymVljPwB2XdD2DYP
h2YkR2vSeamF80JIyrq9QvlP+sweZDfa4B8ryBTTPX/FCJ+FmlxhpJiQm3TGq4Mk
G/OIvt9qhpl/QZSqcfv0hGg9f8PJ4TF7r0vb4TkL0CJ3ffJch3jFtjiFxU9JiF8i
YrH/sJIrFHVtVc88Z+As3yW+Hs7DKJW51RPGtnn4gRPsS8ppcL0tno4xwcNpmupq
jXIVn9ioiKXGwkfiY3ehC3g3xm3Gv2DTjy/3+V2LNHaG+HXH8nLMdSgtyzX54KTK
unIOB5JIJoo5rpJdBIOTccZlkvalaIT1trQTSFaCPO+cWRy/nEdzIeiRF/LlrTFJ
rAOwnLu1ytuCa4xuzjixf5Y1svj2Kn2Cy6i9xCt1XxHxv9RrcvU7qjWmfPc6LJye
PzdhC5WVpCa8yonFE/NX2yX5VA1cuf8mK07dZ82RXIn2enDXzrHVVUqBYVpc0ZvQ
FEl++lbqLRnGCSJ6HFFlbTtNZHAwZtVlD8N2EVMNRspUPpYZvpUGHvAfZUgBRV1F
pxR/7k5Gx2V6SsXa2l/2kHX07iH2Y57UGkWoj3s3rAEXOVi71JsaU22rlkuTRxp/
utwkDjr+o0tLZNDiMmusOkVw0au+l3i6wXAdpwpoGDRMLA10t3pIoOLYvhPXKX56
v29twPs5H59M+iwOndLuK8V7h8XxOD2+6Kfga0dVMQSBD3YxsQ/g+T9vLns2xR5T
Q8gb66u9PD+a+JGC/qsvTQOZjnh0xkBUjUieFiQV5ajLE+JtfFwNwvpeJDX4LEe8
QgT3igXMq2CfTjhVBp+33mq2W7HxYPF1gRd/zomjRiuId2zZ7ASr0cplvOseNI4t
8HUKni8/cYIJrmDsFme/mIWKlikpynWliMMzZ/IU7HTkrQ1g8zwrwupF1EhP/T4E
/eUkVOUpQUfeO3FYEYDljgT0Ji8/JFkYJx3mEL0+aO41hAEgAm+YkEyYiyWHdBdP
nD09dFIaRBjigJwMKbYNUrI7nuTifhbIkROdoRaWd1er09ONhTQW+09inCKQhEdd
axS+uz6md6qJsubfWBY5TUD4uyu59EW42zvkYUg31tmG1KevCzB0l1H5HSDT5lvR
+xh4k/G8TJyf9sRKBpWKZsNIpMqIMzQ8Fp4OWoGoryJpoe3pGB+WXkiSMRB1JeLv
8P543+53aq2YDSC4Lp+8Z11D2IiYNx1zk+mhExADcxLhyUNRETaclw1QRnczRMN6
QPaXG7iXgklRfgBxXrvA1VjMH6O6x5Ap8qouSv3nV0Cn1Vd2TlmDzdvg89fIhp8B
yMrV7AroW0yRmhw9i9CInT9zGUW/HRA6UM3TGxcbCV0ytQwSX+zkg+CL6HwQ+6ur
q3obiEgspTNBACFoNeAexKSo7ofe3vlu2aHBBxA550NdBr/R2/x3Mw/W3T7ImoIc
7Zj/oByCmz6YWnBv9fvlXXRFTVv+nYdZcUrKkQ9ZZys7v2kYQhB2aEdmhGTB/lv+
AX45+AIThR26pq6iC0tc41gDTIOZga1fmEtxxnPedxvhADXSf7MgauzeXLRDa/DL
2g3mGCH8zgIH/2lBBzatVtlOa2CK4ld5niXBGKlrCJbuH5TsQwzZBRVUuhVbRDC8
6cAme4Nt9S6qSEuJ51H1c26FC99YgQy6SUDhthxNdklNSAT/xXTtLC4RRmyZ4gxZ
fXp37elJmK6ayXJzlsqlGOLe08Mq+gWMQ/lkh+TcntMGthA8gGub5Tfedf425iDG
KIZQ/N4QMVcCWBA9CuYoKxzSpUKX2JcG8A2A3OINBZ6BwTUycuakeXZUtzV51veq
/yomTiUbYWLtNYNivwD7pzVZUIiT4AF/LnmEffmFvWeFp3xrIQ65wNQw3bnlvmPn
DCbN09FumpRLNhEkEuwBoo6DTK4YvwMvg1zfBbBokB6/r9ygnNwn47Vajmm3kSNX
13BznTvwMf+tLvttYaT4Qn28OusqIjefzldKT9BtXvUnr5ugJMt3wiQdYUeT0iWP
qlwyc48AE8pI67Im50bJvF/LaWCmsvas/CZoE7aHY0ptqaSdyXR9ZAf8xcnPvgs1
tyOSVfmY+3Qn62Y6cU7wgGp0/gU44GqX9LQJU69cNRk/X/zDH8JLMpqZXoJ+v+TD
ASDjvzT9svjLt8KF44Xlq4cZuSNoGUg21A5ndTaC+31RTpZnEyj5LNFryU2vPDmx
QMKw2CiJpUB7gfOxgUS5t+ZM7W+AuVnSSBdarKm92VRMpBP/2govZ9OaKzEU0aqj
UEnb3ZjwMpsTVK4WU/bbDuaR8DPyRRWEzJCH4vYKryIvBLNxrvkSo85dqHiKRSj6
A+fG5vfNO5bq1dht12w4bTMGxYSmJMbOIqQV6bNbaog33TynPgRtoCM4Gb2dYz7x
DCrreed6ynaDsVQohqbWZvvqcPmh2azi3J69IX8e8q5x7+a+hCEKXE+OF/1ztjN1
9egw3ILZM7nif/5LQKI+Oy7Oz3UXWeJgHOVM+6UBF0lX6dOUZa8otgSVvF3sBlE5
KVoeqK/eN3eeILFJuTjo9IXMeF3pO4+cXRyCpXxfnzBKYSlSOwVVT9JFK9SW/4NM
pk4wnuWUBmq8WhLr/AiRCxJz2YNHc1rTiSmIprFs67U43WJ0wTUHyKwjtd3tFlN2
VhblkiaU9HpOX8TotrqBAVznvUWJSyEdkuMHSDveFfTovszYXvor9Wvx9yc7D1D0
SsE5oyP4s9AtjD8MxptQKqiChhqWYF1fKznxiRQpTBNwGSvfslO3+9+ddFy+QepA
u4EFLwGLByungsksNNs9TFZzcR7T0eOxPSuZXFqh7tKfOrLjtjLYQJPoEwzHiQv8
61W/b1Q1F6qdegRBw41nZtlIbM91HIcZHdPP5xtcKZG0wKUxFcVkgV0fKvZUIvQ9
c5DLjARxkpsyGE3b9N+qnfgC8t/1Ei+BjDviN/O0L0rY/oQUMuOHSuAS0zgaCv9w
Kbc8ut9jW8o42BbQPMxI9SISzXuo7jog+K/JEbQct2+eEag2tGLvJYAX0upoQu/9
ahV8yPV3O1+pvel/aRzS54YuAZhQWxMFNubTZ5DDvHd8VB7yKpVVF+JXbqKnqQhY
yd3wWQzgs4P4bL3RXSWify3xvMsNruO1nVwtcNzg96T74xUlAy/ROnaFBLlNIvW3
mebdKMStLooQ0KRB302KpEf4V50j3W1t527MPlQQHDmzCKtgxCvLslZO9fy7UyV3
MtrByNMGtSa4EI7Ble/dOlIU+ez8uka6sYG8RDDZO/sq4i5uLU3/6zOiDUTIaj7c
Dae6KlUhptBMTWgxBlD5SyFmdfYYe0N+TLWKaMoK3JrVK25AcqQakFnz5Sjc4SWw
/wmx6XubqTN1DcIFWSCyvyvsUi2T1li5QJa1sqwUYTXUlXFOcNVWeynmJq22o1DX
0DMztCPXS4OzM+W/buxbFwBG9yh1sJbGN4QOnI/7aRp/MHzFbGabpI/yQs4Osefz
KeTeczbxGUxh4rLE9X04LbAUHh3jiATfOd5WowiS610YMIIaqTkB+XIuh7pH3Awp
fIhVbIKzj4t2k2vp3JmEvj8ffEnOx38Sb0VDyDrT0h8kcDJD3BVgOyGiPitRnlB0
BmLynfLita3q8Esjc1Y7eeb96O9Aolb8NmgKdOTaXErsaYu/LHHtC2evstLmt5Xw
LaTWzvwfmb3DmX3vc09u4VgqwfMUlkAPZYB5VLVdN8YE5L7U/yA7jS5IDx6pTLFy
lK2Snwtm2GJqifYcf2eWKuXNksNeS8GGvabQU/W3mcrrs4njFzTFgKemhiOV4/d0
Kr78LbXgVDA+xreARIcSrOePJ1vaEWGmMtqTDcyPFbey3nPFlOv6eS8Sc9IOS8S7
R3nSKQn9d3K7VMhzv25N8HIZZ/tj9XEPj6e0FORZazZBrGU76d8XRJtVLcietngF
UhmWrvhYV/lf2d7972+ai3WYVqeehzizeuhth36JQPEJGxAD9IGEws0Iihdv2wD8
Kj18r74qt8+EE01IMMAiESHvGRKIoMuaGE/gKGVFoLvA8ejjh/hbWWlMJbc5XQo7
CPIRgYMUem4FMLeAre6cJRfsjSDj93BVf36Fu9Wr3mU/mE9Z+MRgCNt+uKI2Sm+6
H9ntoj49iCB6ihc6whQefYz/+XFz0vNPv3fwJWSkyGRPWZRdZA2CrTqEHogz55FV
JEtrLbfBYbOtEfN6d98LmwGCYWuWQScAh0Vei7nqGWQ0PmXjt7/lPTz+YBkP291H
oirDz9tal78EOH1tfMNMx2IxILh4GIzwPnC20hpxu5SvGS3qOJujIyog5exxOhvI
vLw4i5X/Z54Vr0M5tyww7j2DIIq1fPuJdTa8mCABBr2E+6tuy91lwMgJYIybvRPk
PRwW+Lkle8hX3e7DPDG2ARVpfL1/mo115CI18A5wTfsXnoN4UmolI/3DmR3sSibA
1KEVreYcPUc0x/SPaAWXJ1e3E3eCROmhcshWgNGI/p8j8DHCkbqFJ4FqtD2/tIHa
1UGaVPXMIXXJq1/yHieB9phGQgm2/gfu/ACSVrPYE1Y+XcizTidQLSXYLepDRel0
beg+kt+Ioj9AGyw7cy8ydQTqS0SusvFMYPz3qBidqwj9YxYHH4XCYextW3rieoEk
x60gktLP6TAmUZ3c2WdGX5DF1U7Ct/67XAh7EaoKOmxX7sJBliuzt0UNoUBkRIzT
iJRHdsqq6yie4Mo0SMZuYfHB5wNkZI2BSJh5Qpu64ZaiOjqX/3eebG+sD9HgPuAT
UpCGSsSrXRNEeG6lLIJrHoQl+r/ePDNHn2zrriTR1bGdc3TPpTmHYSXxVuN+yt+m
ww1GtJrJSaEWVDJmHhjelV/IpmaBlLdFL4MNY4hQjOneJxD+XdwLZsE1L19MWDm1
J96YUc5KFTRELeV3dgO1GbiN6Y7C7zHnmCtxJpe327CWbAUFwshRqCXKtr20s3Ju
MxA5JSDvJ380cU5v2NWmpRd01i4ZDV8hYco5Q8OO0wLvUSjmJRNnnW5DaHPCvfE2
PGpBh3v6yE6UwvINRkPii7UAwzCr8NEryMeMzChfJpObuNOeAvt1nxbRiAxntQMv
ndtISv+yUFEaSBEy+EgsOzQDCwUwz8EjQiv3SYSeYqrnnab3wjTi4L1C9xxzlFVR
a4Xi9TCS3i7YGPrAM4IVKiBzMlFPfhsLK2gPMeiuoNWJq7h6bIcvM9go0/SeQn2z
o4M1RVhwo9bZjbgfPJdQDC9caCd65kpPmvX194/qCQFLt2I1pa0DvpA8mHd82qCz
oz3EYUlooonP5SyRUWHbdYAagipePk+y927JSKW5vjDgxo4Fpolggl1ZkHiZCVdb
AkZPGhYGRZZvJZbr0WMOo6V8lo46ZgYbf4DK6l3Cqp6i6Sy7TUrgl5RjQOpOB/p3
ZNaYUuHU9qC/CFIWDPmil4kLoyOofjqE6sJ5MpqbAhmNUxAeZSiCErFk9s0ECGrD
rbC18kEvRSwTntjFguLCc1l0zTAnrfr02Jyin1ZYHCp+Vy0fEXB4zx5HXlhXX9fi
Vaof/+ebxergNKbhGeFhGTknI+SU8yOI+nSYsKlhtFaSfq7sM23ffrxRElLotVDY
tlOEaqOvtmqVl4aipUDQhJ1ON8AwOrzwXIBfhlnQT1d8tzUu2tk5jaQx0H8vciXi
vZEijFZy3eGiQMAGPWqe4XXoHf9DBKA/ggCDImgkt8/PeMVLCVXyPNG4mLByVhUE
/7Vwk/NgOOLPy7c7S+bdDYECVK/Io1hVtUjY24kbz7h4DzAuHZ9Y30uwSxmp6pbP
bYpia+H3d1bPQeYG+TPpbUdMT6r10VYdhv00kJV36LB4gkGI+NGkQRNfi/KDklxz
JsE/wXzJkQSI2xoIifw1LlJyCrkXd5NdcdVFHSyd/JsMOMlI5cPQdx+d1dp+qPl/
qR5eXTh0PWW+hl0haYIiD7DS3NMlG7ZutOAvLU0FNL10F6MVmJNDKJnS6vFVELsV
KLQDRi/AgRww/RjV9Jr8whkY0M2QDH67AuZZ6edt/gfD7FkECZNQ5178ifbP5QNL
a0//XE3KSa7tyntg7vTmD3gFvqObKKt/cktrcUnEaV7H2VVrh0pSlccGhCEXuCjL
f9+6D604rG5iPJ4WdxUg3Oqz0wkMlNp039AXI/aPEoRseHTndTavUIKRhhWcFXis
dRPm/zn1BHOQVaLLOhXjlUj8czBmSXuvsOLJL3hTsnCgT37hHAPiq1zv2OpoqKs1
vrZA8tX7OfzE02to1Kvy6bYHQTY2jRlgH5+sBXgJ83Feqstgavz9EKzz4MJcypcS
hRPtNsjz7JrZEE+yRJjdAPQlEDs6c1Qw7qF8BgRY5u4Honh28PkuNR4YEZMwkZik
aenQ/SLt+tHFjDc0f+5dXASmy7OyNPENIyPlg6Rs+f9yWTbaL4XeGHA84rMD0w7Y
JjnH6CTxPmR0aTAnoQGTHpqI2B2LeJoree9cKTULY1T9LBwHi/Zuo3ZQRcjZyqHE
j5zWiQMxty3uqP6RbYyOlCZIqbgYyidSylgrunrh6uLLECtUNn2/cD+EAvVqHZW6
lM6Q4qYAKW2uL2oujP5fF9ixVi3r2AjuGPzKJwoO0zlO+4YNL7ydAuMhoOqUxPe4
+HZZX/56wbOL1z39IVMbnGpj+NhlPSUTEeD4yqrdtRDY71hMOrXYgvPO0TaSViKP
2zyrVzLgklOEjauPcSihUnN+WtnpdYcVz67Le5nboVpr+P4F9REnxiZnEtImHdu0
5a3LxoxRSPK8VS8T1BEaigURdvMEnwAoihbGhaV9RQPG23ozpibICTNx2waU3cGt
bQWuIYQjI0tnmX2vyLfyhtzWDpcWSp1vROXg7ZNudCMtTeXdB47dd5Fx/AeqEbv4
vBCX181NuwDZLI1zDDgt9/iGOpcRGjqQqNHo4W4JP3vGHvEMJAdqzf3ux1UmeABS
GnoqqiSgl95RZit4hDP3z1leE9RNBtmLC3h/gPdkcTiMscqzE3/uhjylmITCknI7
eVRuwAg7VqM8VlGDw+02rMIMc5jQPhaM8kfiAAnC//E/cYSpkHY/77Wp/deQXTQc
JE/veB4i1/WOJDlhTUcEr/Eb0kQlVFSU0zjs+LH32041QHb7443lzPoLAS4zu1df
iet4AfHvqSheINjmYOT9auidrucxgbxJYhznufcl3AFrNVpa0kchI2wuhJEEi9Fd
A1o7IZInXR14zAW/yHpyeffDnsbsxYIFk+zuHUzhPEqxK00xkLo/Wsc3u7JMkczh
HiQEAAFlDa2wfFGkwfFNdU1vE8B/Sjic+5HVbWuzuGHNvsgaKJW/Dn30fyfE4cTT
GvIbTlQHTSxPzyi+aUFxDPALJD68W6axeFNtsXXpj8VfV4jmSKjRg1L4cP80EgyV
kPc16lGYiCSl+6jFYWv5mn6pq8gf5NrAAR48mwkp8t4OmNJhPVFDOZ6UnPTfuiTT
lYmyq//EzlPgJzB3tHbNTlpQQasaC+tjWAefftkwmA5lMCPSZdKCRGJjn9ekAUDf
1MlXq2dQerJMtTl4oeZL/MqrzYO2wDgzzTwFxp4DDTjpe1Tpy/unAWtNN+rILMM8
rjs6WYfGf4bdMTjzZvrf+lvOb4Q2n9dnPtIDe2OVMm2ZnQjygBGWvTBIdfSsrgXq
2fqQ+Hjxu1/ONd7IQ5J5K0BBzn63DQEHF8puo5XGnojLRMLKF6Y8Hoe/MKRWs5xs
7W0zf13WNZg7hlj+FATb6SCyTbdtwit/Hr8hQ0seioWMLgzeOhJ2zq2D4ShyzJC1
bHp47VqxBaLHd6Jl7XwSaSd+qDOLn75zUoEaHqps1ZqLM3j9u/XJDzsJxpPNQsHR
2T7I9M94NnvSdLCTwoC7Vd/lAEDMTOwSgZFZAF11PRec/Nu3OdZ62CDx/v4vHcSQ
3W/oNeeQ1qUXHp3PCCFBQHFDH3F0d+puk8KR8ECZ2HKkxxwfRCatL66bF/UyLHaZ
BzfYEQrHe/NzztiIRcb6CSAQoo/yyR2FRIUglx2cFWUcFi9mZvExhqL5A+MlBKdq
uDidFyjGVzksi4Uomc+/hVfShoIemTfRfP6mZP61O/oTwjvBqR6CYvygZreHCSb2
amjL+carAkqE2nd3otXB7puiS6wLLS7u4CJ78WUrdB26sm7N5vq6sZ/bnBPt9zWx
N37lf/XGCFoVqxr1ybfK1NeKrFnjE5Ib2SIrNA2tHDKpRSoQzKOXHj86sB+LcFP+
xTzW6MFGn5T1BGPH3g38iLa3nCHgtXZYIgpkRcSBDnSrrH89eNz+UruKo6HWYpw1
uYgdnEjaM0UZsXokrvM1TDn9IeZLDyvRQdJ5QiaWMLNbe3wr1hviBQHaSB4lpyQR
oTSm8WylWAY2bSmXsAye2gXLS4Kz1bhQRub6SA8mT8gZ3jyEvgYWLK2OrYpK5F7K
aV/BNZKdAlx+4HL2c4xe/nopbOELnwTD424x5ygXS5eJVVClEc8It+zzY6vzB+qO
7r9A2hWMl5PM4TkhGJpDPlzlhxHbF10trcW/QFEvBmBgxqEQNiVzDQCTvua+NWwR
Iat6V2U75Fk39lFS7IvrUI26sqpHgGBsH/Zk2GKwxqFLhGqLTmBUZtNtwPzSCnce
m18GKxdYQXXzp8QshoDqAS0g5Tw0CBc5d/dlYOp/ljxrgcPzAzdOO3a8I3o20wOK
4bNP1p6RBp4SD5n7+ELw9mZmlCdeTe86+83FjGetfZsW2c3JNUQYpTJJ8m7Bs02D
TKnsJ+Q177/qyLjoKv+1II8eFwnIEATfQD85mTPlTq6rNrfpo9LkbdONsKoi47qa
l4MMhsRNwNaaJZk4Z9ycSQThlcilaytO1YBtLLPGXOF0hZ5gCoLQSvGWsa8n/zcC
DPCVsiCFwU92TO2Uxul7bsC83gUzn6NV4Q5Sb5YUJuXSBL4ZrdmT1xF3/OtZseLC
i//bQV4l8jd0ijB/Tpe5Pto+bSKSB/OW0BxtVOD2/s/uv+zW6DHSnuxoaXRefF34
eF+Kqu0GT34P/+YuN00Y7oP0KSnpHpgm0Hgj4xIFqvLveSglOiJbRvDkHYmRsLqO
ik4ubJRu+8rGTFeyHFgm72kHfut+iG2rfCkLA1lMlujY/q1yKAorsUbFevrMVPlU
SKU6mq1s4DJPFX+TF0ZBlkjUAzZyjAFHzlGwrzDrcDSdHCf9StlvaU4B1FmIFGTG
oKph2wrTuD0rD0TEi4Cd+dPn7SFuzevnEhB6E3mkulXV0GJa+lxlu9yxcCIdvPRb
HDdgX23kckCQyNseav47A9fSep6zhOELRs9grnsjBTJwt1x5MwANWUq3egtfzBRE
0yD9ip1mYdzKmLXPOe2yWR6Z4+dksy+jW+mSgC/UXJLvLhMWsepoytGs6tFFLDLM
KKE8MAczesobbskLFAtS40QXKk4xyhlfsYIK8etadOlR+shZwYDp/DC8pOiam1BZ
rYOZ38i1DopMQNTMfjjvYZI2AFURnXoj7gUZvWLyQHbsYZHzy0buQLKfX+X3NeA/
wq5B99nxSvywIQba/av1zNLfCXRpEwS3E29vewID7OMWVYcbt1MSyeVEX1YpavP9
A2gl4L7uhwMLq2Scbf3/D54Y0RebsxuL51s2gJdbYykZH+AkRguE52Ou3KPIygO4
djWOq1+caTvOAE2CgWdOapYy7BUfm9ShkIwx0GHoXMDbja+GkooZz2v+c9dDiEZJ
Ml4MJvOdorTh0Yq2O/UBfOEf+vE0pclyRifdM7/beKV3lHovXAw6JRuknNEjyUwC
XrDqOlBELiD6VpTHCBJ/q6xs5196lWUSpRB7/4IpSilOlrL0hVAovZgVLmFfTdsy
iBjsaiqx93azwFrBgd0vpQS59R5ibPEnSiwcTtuCJNLWX1NPWepjmbiibLs+MHX+
ShLGwVenCTXSw7m0y3HNBy6fvT9eMe5v5pUCmbHxWxR62Q/fRprOWto6PWFQmeyd
tUmj31U+kQPWtGswm0pQY0ss7p7QPsbVSBQobhNTstpr16OIM1ResUoaCWH55Yyg
AOgmCS4nMy+8e1BwyVJjAhkPmcsRKflLN7uP29susGvvue0tmGbGrRV+Mqo/rNEt
lZCi4jqoq/yhRFnyICeuOCxbeoU0/kXY6DeHQM9WvZutaOWub1N2Wl5oAzS5lRLV
Cb4Ph4VocYoKy5I7ftVibISkB96DtpcxSi+dCxCzFyjug7/YA1S3n8aqsOgbTa5J
wrgBfKDDDmI7ZiWhkwRmIOGTdhu7grtQQuBZLw9KO80MtYrSasbA3TyJvTL31keP
SoRcgZP2xPK0qETF8unOhMUK0UpJzi2TMzt7/2+1f4TE/uUWa/HFQrs0qE2Mr0/I
+Tg+LMuhmfSzE9YCmS/YPj7nHcPAi3qoz0Z4cB5nCd1ouT8kvtqEMaprx946Zt3+
n/ReE7crrx/NpVEw5/90VpGephr1Gh3npL3DZj+GcJxla0ZI3S10WhQjWkPynljN
BNkl2k4oYgk6Jlv5XwlEYkKIOuBv6AdS3HrM0Gd+Bbj6YdZ7Bt7uYEt3SU5Mccc6
Px/MNdc7neZDAW3y6xGCnrL9KnRtQ0HXwbZ14g1cOeDSamOj0pvIRRKCz8XyaV3x
gWOvAZL22hBfKZxMo3fMstYISmbK0aaraN84OAoWNDYmRVMDL+vY6ju7AU5HFNYZ
yr3y2+zD2alHqrLbh5QdMUrSQK9a4BDiq29kJXDvVPjJPs32/ShfVXZL4DtNU/zJ
LvZom324OZWbXWvy8wGepI53G02+zqMq02bt/1XgQEt+qDR+1AyqfihQY/Epv5Bo
1GdT9BcKC7dPcqzAMDydE+8PK2tSB6Poly8ludUhnySd96cB0X3MUIVbKT5F7mPC
6Pa4+DTvIzt1eT6NZIZWznehkgBxrgMWxPbMInE/bngYTkBWtyKD4JxmoLcimNxC
5IeCToWxWNFHeyTYmlc+z9zo2exL+AMyAKLwBWAU89zVnHYvowe4NJoE90sI5ARj
oO/uSWoBIhfBnIHzFAuJ7WUg8hgPaAc68vhbTY2kZ7WgZ1AQoQz/fqGqUl7Y+sTO
VCViuD0UozKN6UYC5zQ6SPbZjMld9sJsQmVeBYICXbUeh3oQCNOPo+FIkmJ0onwB
vyb8K+OXpM6p1vV7g8Ybpeqk9mTvIRqQxYUclI1W+UTSYXP7/XPtT5jCEpC0c4y6
mjdUeBz+MvceehVgRjeSolv5n0tCvBOOh3vwM1Kpmk3sdH5+TJ68S7shCMEXEo/x
5sYmIpDqulcqLgyftkE3cbEURs5nf9qqk03Drmw9vFZXxsJx4Vs8zp/0CjicdgSf
AgujHfulccS+p/zZ8xjtyspWplPgEnQHjUvzYvtQsoeZZiRGId9sscLZJPJzrLFD
CHQdKpVNJ/zgTZPHaJG8HtrHYEF8xzo8IhDjOGUWb8YQj7i3q0vJiYz1M+Thz/5n
ALDsDdlw3FfkDZyhN5Ijw/3t7EOyMlDNrkCQWAZuqjjRgyAr1xEySYIHg/iFaKiO
oeOQ+81F/n0cd49j4bjxMhc1qTArEQk01BcMMIPQU1p+k9rC1W47aI9VlRdeedjH
9m78BMGdc0lj7GtE8FsTvskRpPqd9SmYXZ1IUGAYP/QXwBkuCIqlKV3Q8LqXLERf
urtzDdwYZHOjf/rXQ06E7vWctQiK2690B+gsQ+OzZKRymRQQnxmTEgWVcqUYcrNk
BWorZI4LEULGLXMGv0ERRYeeRXd1jCMf8T2bcxDz2L75wvSjdPRtT/UkaxSfq17M
xf5bKReZyUf2cTpaKDBfxqLTyd6G3Z3qXPQhXmf10nYbrIPAJ5X971gJq2Hp0zQP
CyMJW6dAPSguGoOJ282Vdn274OoOIke09wKbEvblTEIjxWnzhVktoPEiaYlu+QEa
ArAlYXPlTaFrwcNAbgIpcePV5NcDi2nXzkR+73akGTRG+c49cyALwsakgYYWPexS
dSQLNRe5dAHAMNQXqPMzMOwR7NnJnY1Z4PKCErnaJFBCaXoV3PjSJkWhVMSfwlnx
kpOQ3PsnsQXUfVgTp6JFgg5J9Dk1gCDbnTTMNJ22obKwJCBTHpAavnjQAPpsjMjc
IZztKpz/SlXVSiOa81oTiZhBv3v8TmsaI1sg0Mxv8guZTokXVtJagfauEZNTOpuP
xpB/AiE9Ggc+6x3MDqE0dx1aVZti4OBI2vZpt58CWOpzVpdr3PfzkXgG4nUpPAwM
TalGStNAsYnetDizrACKkgJqUl/QfOX2/e1hgeTOBCbG0jZHSVdE348Od+uVBbmR
Yrk2qwjT9vW/w7duWwGTBfqUrNNDKmADoggDXzDl9lJXu4hl51nSyxHERNpaNrRA
SQxP4yzbGyQ6HZpbWYzPXpjrDmeSX2ZR4w8dCctMnOnk2jx1Vr+xJWReGkf3pAVf
CPoZaVCXzCkBCeH7vNEJ7Pnv9vhtkUx8/5zDABrIJ3FXYreDbSapNg4qWRWv7oX0
tDWkQGm6Uyx00J3jtIbxJ4XfXr+sXu81P5oob8MPPk6UGxKIsHE5oeTvM9GwVzqI
U4KfhfZg+oIqssNXT7CH+/fu8tnakzHoav0oj/BprCEMRXnI1YZgr+BJr0Gt8R0r
I4/bTqXzIU9ncmilXzzsLA1eyzs0SPqI8fXEZk/hpNdsV1c/VxFTCBVPuN7ssBVK
KEUFCPiGx/4HSut3hf4OVfG2+sSAH0AXdjLWZBhqhjPsH0bttZB3Y7xWJGxzV++N
tenL5xo+9uEajDOBRYKsREYqsi2En+xxc2Yv2aTzz3LYDNRwIp1Q0k2qx5+3MZBl
BJJGWS9SBJYgnoYQ7AdscuTNMqMBzjQTdrhWUGxu+Vb5DHbUvv6x/igO7Lwzsu7q
5+IwCBMfDhUubeiiPl+RpeLs1GuiHFUMFBtn6kUrqO1phaKYT+GSEu4bWTHV7Px3
ZlmsTPhxOoVbSb7TgKmdogOUjSE++PpLmgEV7j2V60lpzhO++bE4wr2Wg/Goay2h
tMUvWNcnsqM9T0GB4x9lkJB30doN1pAYQcPsLCT+djZDg/coqBbVuUw5log+aOBE
X2iQ4FvYnITUxo1aGchFqOCYhmlaB0t9qlfb4MIC+wcb+CGfMlTknj32HSmbj7q3
0a2HqsXsEN2i+dilguohSiRjYFX50RdyT8xCNru/kpzkAdDs7iV7qxcHqYdciSA0
vS0X20BO986AqsYT/U+PNU+jYXHJXKWaGtFyr0cCVYw0WCVq7Hn1RipsuDNpaJIB
hS3QlpZf7U8Ig306KxmyxHUgHWlgIy8jbtZ7mzcZb3RS+QXHodwkhdhEP7JbIfNq
9uNe4VGiXdB1zrpac8aVQAkrlhZYDgXMT83vTEmYF+peHezBXtME7PQ8BdDxDmce
2Ne7YOfCQQyd4cvH1YFx5syeLGai9vZYCSNebCCsSgE2pKf4XR5mCw0I7R5d9CMw
jUmgrQDkakW1nu26jQAOlVBJMCssyI/EgbXNTaIVds0c6v6HbZFqVn8wd/eeTo+Z
YZYgKucWRuymb0z5uAu4YH1Y+tr9Fy6p0WoxjZSE1+zA8NJ2XtafedH+sTr3y4WB
MvPnLiZWlHv5wcVZ2+o0w7HZe8vbkFooG2AWqp6zq32N5BbC8x2oMj1ObQNUn6gi
+n6yXhvNOubME9AFgPNYW2r0XgzmiBdGBZt4L5jCsJd2+FhzN3LuQ5JWfP9X4Ypq
HE/+zTyMNQI+1+oAAX0MxvpUN/FnzzDhQJFpX2yVoFLPA/YPoo8DiZH4WhV9aiqZ
kLjPRrbtMR427Efp7sBhpcTKipW4lCGA0hZnCdtvXZjJfwhcXWVp1OUZtQ0KC11m
+ICTAIatdiT9ThTXmT+VdiSLderzAnkDy3u+kYFly/6gy3dUbhbr1trYXz7gDlY0
Qbp89X83/sKNpr2NqWtCM+1l89pAqU38yMsyHSj9FoykDdI6je8yhPUwm0i+IJrz
bZfQOuzhiIpo8Ee5ZRUM4m8Dk0j/B1u0tDVbLmQ+ALBnGWGeRIVVqNbDdFCVj0rR
Ks9sebQoMSAQ8l0+W9m3cY010C29DEfgGAXH66xeLa0+vaPX9SXB9G8v1A3p1hc4
v+3iPY0tdypOSwHuJkRLRRS2d1vTlPdJweHVFDSjPG02DCkZGOuLut+w6paypq9c
DBJC8mwRRMbW36Rey5L4sgz1xiMIPAoxotyKJEMaGeEhUTuaa84eI/iIT9iEhRoj
s9VuOEGm0zw3v8Wn2VRCEvD1T3rJR3Imd+cXrRIfDh6HORuxY6RNyn90j6MhEB/F
LWlLUd7hkx7yaBWlbE0AL1/YTOsW9uhnU/JfIh4DXWoj8xuUHI78YgWTM3OBHxl+
+01jAlDz2qiqm8QeT7zNVnoyJazDQbmO65aqD1nTzKqemqUNJqE7VKxtRYcOJM2q
Xa/2lgdES2mcnhMCgJCYHfp5lXp/agfAl0SG8Kzrm6/RMNavCavqGZhpiqbF3Ade
2XPXadEkzI/kWHIfLz2DW9W7l894RrwV8LWpeMTpIddtvp457na9Fz7aYwt1bPd7
iACfNkMlWjuNWjhPNdYxVFyXY16zRfEcLU9ydb3WpIyB2j1iRMS3EB6OCrPEhHr0
GDxRKWT3Jzqw9dLJ9IAKG+OY9SpqEk0y5HEOoiguTz4qx1UFwMirpCGg1Lz30bvb
vAt4yhCCL+BV5f361K2uVQubH0D+BT9rc/hfXZWkpaPN9UpvKssrfNxxN7omfqFN
hl4mzAb+JSHNJny9w8idH4JfFd9B17mzoXK07FxtpCtJqgMUe8zHxUJ2w8R1fny/
YUdUOIHcsi4d549BPiqqLF3jesXefblu3G6fT2jLA3/X9o7cZ6gSsdxSyEwazbDf
wZnjfZcMEYNaYiX5mWUDIeeW3dTck8QdmPD4drHWSPGoi/TpHxw6eWpIW5xzOWam
pciR7RzCQZMODagIZSa2D4e23SAu72arEnjkGhztdmnQ/6O6oF4u++YsMxMJM4pQ
Ix8vklLY+gVC4lN1M76jecppokMSC0RcHjcpFmO2JnhIHQQR2ZiKv+dx4R6Ffxc4
vK9K49/t6Tj1QugQw7YTfYbodfMaNFjNwO8HrVydWUJspc9UT9UOgk4o9UQKKu5t
ddAItc/kqcf58+JWdJQt+Ozcro9/WAm2aHbvHtVWUmBNg3+p/s5NHVPt3d3TLDQO
+icjx8m0CoGZrhNmJ3wYNb5fjlkqXalfYZoIvJDCusT7DXQq8EQq/u8VLp7zS385
DTzHo5kVU6EnyxfEgqfmlY/Dsnj0W+D+pWYyVuwcSGVBvrXfmKmJ0zkSFHHkvreB
zAM6aUe82VEp4o0SohF/NRzJ/p8+ZZpCCbecElKvVzXYE29iPbTADKKTv9l8lYaX
z8Gi0ibxqkpiwIFbzvkkwTvidpiHONlSHDRQHZkklqev3ZcDdd4cUgul+Bf2mPnm
fy74v1LAFfejykJCV3GjIYCz/4Fu3LGp9pVfabpqbPjNs0lMD01EoCzErkV03MLQ
2VXTvVGiIuGLK2+PJUPOCUj1buYfyQyrIylX40FnvwqKI36/QItVzjtcXKKSg59r
ng5JqMzqbkSTjo9WZiHdpf4ItftJqATNhiC0Cxv8lm/1UNuQSDgFlm9O68QNo6b0
3kQKhVcgXK5Eqa9t1AAfc6WcSMklwJajfQYyrTySffO+L1fqLesRab87H3KDRuX7
Yq0c7Qo4FvvS+8uxo8SMPT1cCvks4OKouKWpdTa1SXR/hfYBbMV+H/HsemhCO+QQ
kv2IcisMfki04Lx4+Nv6Htm9nzGqd2uxJQ0RJghspwzhSTTStliKklHkxJn7/JYN
QKP7GlZvO9uKrWaIRBLwibyEO0lW+3aOpcA+ArYZJ3LDZSFPPT+n1Gm73gd+YoVf
fM95FfhrsSYgTJCfgag/FyvHM3gKNvuYVxUkch8sReNJJnAMdYbLjaFffrZ6ShrF
z6SDl7OMDr9lbUgw4FELVtDEFENuknRxXf2UKjjRkPAroZhGZ+ofV5+khvYlpsou
KbZQA7ENiaHTlxuAyKmNuRkV3t5XTnxgkVV5grqMORueiDHAo6lMOkbvLa3sYuJA
G4pYfNtrhkFItvgoymnc6QQZllAe6MmJ4d4d4qqAAW29qpiFzXb8EQVXRh5gBUro
y1pkz/PHmussU+hDu9xZ+SZpBhl8GELOBdJNk0pSw3F8Xj/c0ex5ZM6qlNZeTlI1
keGpHZCHQwhXT5Et8zEPUeeBl3nKVOeYM2H10yYPnsh6q5Ok0dW/85rvxerKfx8J
mlSEx7ujV40Dl08gIUnTWEHT4UFxVOV0054AIMVSVMOWOsYSTGfSM45fe6UCBYnT
Hf6zgNt9PbmKC16g2nRBWMXfIu/5eEiIJSUqrcLqazfttkuJi0nAJiihUtM8/AP+
aHCVUBrPpnHdrnquXglD+wc1YKr5n99nUb7NPTzk9K0LgJAPTdcB+7uOJh72R29N
lPmx03KWP9/o/BMTcIR/bKhDMgVELdjWruP+79jDsZzyoCvNHVDdBI7qu5F7onIO
JvTrAv0MDFVa2+7bMWcL0FzDrGAsID8y2wl694ZJJQ7L5jC4clnWZ58NgeWtLgu7
OiKK2idVD5tmvOnAuBYcYX+68qyKe4maUMfY1V/BS0fQ1M8faZ0gOvUaTbYaCK/O
nisV/kXgiw9BdALcscB8K9bkx+2pC/F6+AU5soB1o6F9wd/uJx6MOnoXau8tKrQf
RZ0ENhfIUuPW9RcNCqs92nT0bHMOUivGCqDowu3tsjKa8DK5pJlqlxRhc3nnNpLs
V8dwfuS3lXgTsxQgyetghcEP4uf3mVyVEnIrc1jR3NbHyCt9USsjvyuadWSSKY2C
qWLzQzyEtDh3o2ykTdgIjvdRTK/nM28vLx8bGOt7qYOzh8NQ4MCkdueULs/sVe0n
UvbiKADON1R6P+SN5UXye2jcihfmPfYefa5NEC78vSkw27kQOo7ij58s46bJz+3f
MG1xrVIu69+7TTyMvFEvCrerYDP3qGmAjIcTKQn9UrKs36sO2SK3Blmh1R73G3mn
e2di/K6q4xj7OHfOrFjFO156LKx0fE5oVSXzcbeIw3Zsuy0gL9KNvDOQpKewkJ28
poE0oMvqfF6rauo/wsT3EA3fQtHnidaWABpmBqu7nkMDzX7DujpDr4pIk+tgNceo
vOIy3KIcSDv0W+QavEGOgdej7TRvD/39lQMKmF0K03v9m+pwz5+kxHUQ+4bYtbDp
2bKqR2JhhGNJyK/9xtuMvoldFvQdgcfvm9txRKAJsfNS8nd9rY3duN0G0nDpyoJ8
VrjsJ5GmFq9I1ZftHSyxyrhnpxBrN7a90ER1rUtHp9ZElFTJ1RiL1j3OC2vRONcr
ST528MfW0s0SZ9N8gQcmPyfHGMOf1147GX1ekHL7eJcL4pGoAm833qdqtaRiqhUj
QYmn9VT61CcwihvXHFqrS7n+DVhMA5nM0yMrHs1ioQkpkjHvPNYN0nZ8Q0uwN09g
bxTHOY3O4DYFgfF0FT9L6K4OteutExRXzMxeUTIpMe8I7AxPj6y27d55v4Zmc7ep
JQGNafggRPXpGtdiGdK9lXVUIAfcB4+xvsQRxH2RkhK6E01Vrkhra7ZUgcXCYlfL
yKoo+Rg+mt5ucbWefK8Xsd49T43UlzGbU6qcXuguRlecqTjHsB8xad+yOgtLn212
fjRA2bx+d8XkeMwuqpCTUikBZfLQ3AasuLzNaGnHLWvol7W5Ai5Jh2GqECRrx8uw
iAEPlewCb4LchNvyz1QrSIRasl1z8KLwU/hfDui+Ln+klfZIua4+5NuYbKVH7tqh
3vPqOo6JkV1Wa5Nblzpu5QH/rYof9jXH0i0r6yh7qQMznUoRpphQkKF11BQYpIyP
Oerx998mY3WJWNTSK0i6tphPWxS6oYU1+H+wtex2jGD+vh6ddzzjnQA1hJOEL2bU
Li7VpMjj14yA6ULBDkFMzpXacCY23iPEKwCvLGrFv/X6ckfDvID8jb0FCdZpa7uH
z8tbB3caENb9GH1ksRTkzmwqscozntRDdP+wZtTXysHLEurEqZ+Rs/ZASe2SzL46
2/rFSKo1dqHzMdA3US52QquYIsMmv5HBcpOD1I6e0Wtt6LSGg73ECTiVwxFLdf60
ztDElHVR7fgQHowdeTVM+lT1py9KlDVfGGp07vxY9kku9O890SRprwlD+fmEUJKr
nE8yrsBaRUqD7ig3ff2MiEzjF7OKas/arKJx8XN9VD3WxSIQESz/PYFDJmO/y8np
p4aBGg3PMEeKdhuyxdzaYQ2kuAuRlTsLTLGYQkuKz/SiTVf5Y3OQjpBTR7TJBHLq
b8NWPmkdHNcENiuKc4BPpB028ZuDtwT5Kvks3VDL5ExkaCv0Lj2QlsvkXLo5wTNF
+huwVgb9mkL5h5CKuMh2ZNKp7otxCxuuLTHCdWm0xRJVMA1nQVaXi6ZHmnJuVQrF
PTb/cs4ZGhwjmxHnJzTKT4iIduhWF8fMAcdRi+sbkiuhv3YDT8bh3qhQBMvVG+El
WcxxEv64i/1mnMnTdWdeeA+0e0eYiQMS1phN+ewdTzfO6ABwRNLbixCkYg63MabH
+OljwWq1Bz6MfwQA77qloyzuzxEQpmYRpYcRc6l21ZpegD9z1T+e+TY/87fv1+BK
pvT5dJ1akw/Xnd/L7ZrrJBe5WT7HGYSU9l58eAprYwEO1fZ9GmjREuvWSsuw4nPN
kZ779HS75fz/ESV5K0FFs2ham4K5/y+g5tdjMeZHNP6L/AJwIYHQorEN0r4h00du
uRQ130b0vubgdXn1h88crv4Jl/eWQO3oSM6TgZch35twQLUj+xykgpxN7IOz4on/
xWV60q6pXpBEu2UC3grsQAtnTTMB70bynKEIIfc2PLmGWvZE9xrfL8fjacfZT+WN
IvU/od3ZeqGcwGHc8LaTwmbr/gfZbWx7FZsZFvRt0riRfO+tDV6jHak165CNdk7/
VnWZvanJ1dZ+czdsPLIDs9OnHwqt7VtAhFhZCItYW251g2kgKTNft+YCSUaytRPo
tBk9IQRgCqbH2eSQFEa0sC2w7VhD9Cunbf5C+tjv4Zp/XeYfnJyEYDs0qQXOJA3M
+nvOYlAOpljS/CU/H8P8DBtHv4Q6vi3/6BqurvuVoigmnw4W3pk7sQXPmaoyNeM6
bICOQV/z1hIoY2J4jbxL8xvGJazIvhuGvKdCgQHq5uZYOPaTCnRq4p80W/WPbyVr
N5rJoNXYZ12G44y/17GyaptsH43vsmBvrNGghyu/y4+8Za5/BfP0SBJaKmUPpX8M
KyVebH5ob/bHmiMpW8eEDCcOgfZJypNIW5OQ1CXJ9jmuBpPxHPi5TqhQc0LrdRte
uhqfkxC2M+J1ewMaXZtO7Q543EXrXsPJS69vuQm+Daft5XFhNsxNWKC8OwvsBwZQ
87xEU2XpirB9SMKX30kW/Gj3dYrAktIY6+YMRUd9LYdo5bbF7Z3JLjB8TqgRXO3v
9zOjmLVGfIgd4TV4+Qgr2LU6GMtghdDqCjsUaReDav6SgB1pMo9B8W7hPj87aYYh
Moa0jiZc6gPhCFDvBp+rtMR5tjuh5CONSCyly4SRxl4A6g8YVNWcHzMkHYAf0BWe
xljCJxA5iUCkMofQ57kamI/Z1Bjc0dmc8OqJb7MapccBife/i/yqz8tMQEEuEXw4
7ZPsRr5idOWvuRTysECQ9fd6I0vxPt1rMUGelUuBEsefjUsN+iTfC1BKGK9c1t8A
wSgEWfupsUK+31MAqsZ+2mngoQ+SiNcIvMxFx5r17190kdOW4UrdLQ1DrOHRoyNw
UVzsvpMSMj6YssJ1Fz9y2ZO5l0Ygs3b1ukPT6NlPpRv/sNTl7V74LJAxv4QGMS5a
PaUdngiv7aMQD+egIMHq+CzzsREU6K0mHUWSIuE+O3y479LaznLamJJw2Q0QCtQI
ECJJtaEtPIj3N1819sjdMB4pQKfilUYM1SoFB6nHq9yYmSkjMZif+Sm+iFhtw24Q
F/pmlXU3P0P4dDj0td/bM2H30W5lcJ8ISIK1kizLRKD9Bn3+U1w5A7AHXGapIJUk
+ZspFVyCdgKtryHQuABBc2Fs6XRCjqz1+0yzFxF983jGJpbQXoA5yMKWwvbowJzu
KbDIqPVEn8VM5SVbQYc6nlaNfeniq9lWvJPFX2vRVvRy9tL251R91h6gAhNra/aj
uUCi/PKYZe4P49pj1k9cKs3xrvqAzWC8QaXmmjmNaAIedsE0hWspZRLH5+g0eExH
KA0qdMDMjEpUgYOgkesoCHxS7UmARBsCSwOFziS15bKpYBJ8Kuxzsyl75704b6+Y
hX6uji9oaeyHm8no+r2MdhAbsHS5GKvMvdEHM7QEdpEpUTvCmFRKJJvHGfHBc5dU
I8QrggKucud6FwKHI9Dkfz6kq1qvDInOrpy4NURJHkQnda7oQlfJrXYa5yFUgvdz
bTnjVDHLlRdaBRKjHulQMFjuvuIOEeSpDUzWJEQxSTVQwvrKFhICSSjO7lxjzs8M
tDEspwx2OAUIaZlWNBwV7MRQhFhlCyNULCFrSV4oP1TBShw5GAI7EXH+loHxjWBc
vMjBandicR5q7e6mZ78TWW9eWnCzEo4VBhG3EToGltlWLCpxAXMR7XHahygaj9Vp
ZMhLUboCMITJCp7oAda0DeAa0GiKBwgQEEhEjMZUS06fBAbTxZTC8jwJuJktGUAW
x2rpvVNkALIUmOIe2wFSM/srxGrvU08lp28lHzYMFuLbn4IQK3m98b+k2bDp9yJh
sYb1VIGyPUyohKX1umqJ8eVY0A7UswT9bJ4aVqNWp1c9EcP4hYWbLNvcgBlXQd2K
rCmvf+ugp5IVM3vf915NJL1TEneOOilHdE0vgqI92eln+lueSqT/YEjjz1C8i2BC
FR0brltJRWbFe/WP3bGr5ZXo4g4oMHbnE2z7nkzTij7JTY5IpuaYlIVmjXzuVXo5
9RLvPl9lE+ftIKdrNArladS7K+CsPiWpTn+0p8FcE+VXnVeYAbcq9IKx/4A35/bC
yS7+aG+ZPIZLqPUxyspTCf/DBFXWHpsm4Mwv+zw9PECi24N8iYo3DkVKkVZBmfjk
Qk9cY74YTgVo1bODgJjBc51JckFBuJ0esTHKPt2vUNF6NNt1RuL2kklkxXHB7Wmq
P9eKEaHZhaYA+yKgB99Onxe0aHyKpmxp3lqa5M+G8MSt2N64GbUKk2nxVk08DopC
6m4iFDxDlBNkYF55yUXGfQO9b++LTMcMIDzNawYbc57Go1tqpUkn03WXczNdgrAk
u4azlbwQy2FqiLj0A81wNpQNuGiLnihtrKcZLd1tYogy56W/r48gNVKhSBOQPVVW
AwkpSfdPiAu/EsGOCcYOP3TCOqH9uwk9eeW6xrM7Syv9Dc1q4n+WLLXNO8GfGV1l
O4hFsBW/iPKd+AtkZu/9IlKa3TG9aicn+M10KuVOpuWamH1pIsmp+KssPUix+f0J
9yxSw1WDHfLgrJXu/pS+G9CclnVYVGaui04gbUu5VTgPwmxnE46bMZKSRB3kZO9n
RxKD+voruRnN0RjFUcrKuAy53lPl2zoB20P7HT5NIKDBKVW4TiKnGUdAYp8TVHuE
4Gak8UhnfCjM7Ljf71JDVVN0bKLEiJeZA6YwHlox2dzKnGKFXTBn3nMUyubJJm8E
Y0vv4PUNdJ3PcIyf3vQZ6EJ3QrjPqngA7yC+lWBcnzeIOaOdo5bueyygHR5Slppa
WhuetZNmlHHBEG0AQ1BK/w9h5XNJHXMVPtVGOtv8BoKdkyAqhkL3c1hWGMFdx25Z
iIIVBT4H1KBzygdg1pcxZheIMpBvVkrNYYedmA8kDFLbAEA8U/ycXd2hYUHzfBMC
c4+tWSgAwqFUi5rijFqe8t8IAsOVAZh+HXVUtFRsEe6bjWVfQeMxbd43swvyFChP
hJ5UTQmKZ48OsVuq75zMYoxzxPQRg54F62qETy05fJCicJ2BD/Sz1m52WjAgqkB9
dI+le3VuHWVuytADbatmej4cp4ZNLPUEoLSt/On6guiwooXgWP984m2niOz/SrQK
09Hm9H2VUOSKm1jFu6Wiu82ojB1i34eYhXRG+suDkEiQ0LLdpA380bgXnDTYSQdw
lhWxxNQSE/Tr2qwZmwQCJ2HFg8hZHrqZ8cu/0CWYbZXal14cSMRhn7BdlU5qnaWA
zuHWrsbbaseckYn5cqajG9QttuigNX6zS7+7iMO++9g3KhywEJC4vcZyLp753SKb
dh0t8QQOD7SXqoqXGj/M5+xsKp1yG+VcVKS3Vup9kzueGqCOp5us2TkbV3BxDtcj
Pkp8i9R1d5s3DKjG88xNQUOmd774QullHfsYxo4hoFbSxHreIk4gXPXvpg2JgWfn
EGDpOZ7Ab83WI7PlI7Hq66gXgFZAOu1dAOCSiq0l2gsCVTUevPR9mhFPkdPoUWjW
kidUg7xwQw4Yci9dKa/WQUy4sv118KGfQR4rrp/P3KaeChTkzJD3azsRqkvp0qux
thioLFzBp2sM49BitZ88JAL8p0AAxKI/mBm6j8AWrmfk/m5b6ycMYDdwkk2hdWzl
GslvU+sqkYSYvKeNN5r/AKStt95sEw75nII03QZll9LIVVb9RlwzJr444yjJLtvk
wxeimSc+dELC9IFF1jMUC7h0I8fJD8BQ3J4GksdbySquJLstnGxkAG942ifTc1XE
YmsmcAJYvZkcY5OsvYpD9UZ/dyx70Qqy70hW1aBCyT5mglSbKT8y/1bQzDbH0Syr
XTuJzIL/Eq41L9ckHU+08XabyTZMaTZ8xAs5WZewqT/gBsSofgoomFUa7vAIh6ff
4I7GQRzcbSsiZL7PzznwD6JYq4BQqqJxl9aSTDQm+9rELA5+N0Ng6howMw/b8Rtt
Ea5mXxXYQa7Loi0LIg9gC/JBFJgIMFZtWTkL3oZFT4aAL6BhAkZ/YfcC0FHm4fSD
/VrxGxmA7WnqicOc3m/m5wb7V+ErKI1eLwI+H36gtYYc2Q1uTU846tt9e4mWOMY0
zUG8XhIFo5KW1cj9pxHtgGsg/xj1hpHPInYpN+iN6VGrVPddPNGOYpArr1FklRm3
PBNNlSepOiyTw9ldNo1ffFpbT9uCIzSK1hk265njprxsURhY2P3vHs2J6L/hqlG6
3XnrrbSx45p7i61c+wh4xo+aQz1ZStojxuKb9J8ZMZJV90zPbV7w5UriN2SSffer
09X9IKha4GpWR+SvtG1J47/I0/5Tm7T5dVS+Fz/DrMV/GtcWqE/p3IsggYeDT9xW
T5wmUEb45OLW9CJg9mSvlk2goufTJXzOCFFayX1XFhyhKWP7aBAVVpfdPQxujs+E
gHzDY98cRDsiNq1GLG9G9AQgZ4pRStnA9Ux3YQYR08yYf9q9QkBP6YkPToDnnhEk
2eZc1BNvuzJpk9ADOpUAWM8VDaQ7Jjf5lwszrGf0x0LCQPkvU7TTbS08YTkopR/2
6miwweL/uQ/1J0j+w3heZDXu+tnDDgI6KoaL0Zf2n8qJhkbhqulcud33RWgtHifU
eJp4jnEx4oOPFk4wOGrIUJjWIOsuqPycZeeFmkLvtuvBD5sm8WT1jZwa6/QeBE7N
XWQw5j73ex05PWGI8kE18iBrz6fd64ryrjt1aIRFTXyOsk3t5dmo3chMmToIx49U
lHRuyyi7uNE8UVFKju1A7rJEMKuVCrne3iRuDgt5KJiXzNttt1pQR85CU9p9ZLcs
Rnz2Bv0t5Nm/+N6G+HJSoGf6HqcsOn8c9co+2easRIzrfgSSduQhRu8NT6AKDi2k
EQ2ObGbIqHaeD8ITMz+d37sgLrAK0kTrF+HR3uSCcCckwgFMRnoRehE8Y038ax6Y
nI+rE3HLri3pjzmv9R61guzCOT9c30IA63S088LBWeSDknQaN/Ga5hdnkJ0m/TGa
60bqtlii0HzZtvQAqNCxN6ZbFO8S8f1V8tRFxA8J6Guzz/ZI9ZtzgHZKpcYjSi8l
xivXheDcWiS96N5GO9H3C44cRgGI8UKfsVCWO+uXOi+5AAYQ93KgQdyyUUk9KpS/
QYBF0BGItkREHGosP9o/RW4KWL5O3G5tCXPwB+AAHJqoCddPbUXcM7Z9RI4KMYU/
HqWwX4Mu/scvhPHX7YBMNAT4Xn3rfbKNgeH1IcUX+z0x75mjSgXkqB3Zzwws1ywj
cCht4gaZztMcrwZ3klxcbOrGaf2mgmEnRZnfSsXX1duZGl2uSfBGB4YgfWH7FdxY
IYevgLqOdUcmJJkS06DaU2JP1TVAmS1y6Q2FPzuVtsU3szB4oV/ci4Qk1atbJw7m
svTfRhr7qoNz88AuHqE6O/6S+Ok/DgoWk7PqGbERaKdFqK4OxTImydAPaTzygGms
bE9ygwpODcpU3IABhDCVGeoldSp0AmFfJR/ehCGtSY5mSB8e/9yHsNMCQ7M29XZN
CgaHI6Dx6NGEHY2DpS2BfImC0vk3y/PUIxlegEugTwOcFWH46gYk7XAN3KOaprcb
FanPRwfp1bY2BLjO/wbGura0NvGm7ZtRIMJmZGBYqU7SJy9ayCLbQYmWSNsQjEkL
U6vFXsp8UmHLY5IIulpbPnlgVrx1bOm0DjBIaZtOHEk4hi04VF9y7S0pkErj7AsN
u1tQ5F4MKBQGl0bL+znfcbg3p4wD2R9HpUfuE71liTB5okH8TY13t9smUvOMOgFc
7wi4myi5f7+xgAv4go6DBhq+7iirIJTHfar0rpIJDLDCBjU3ZtI336RCHt2CpvwY
0HZJwwVa1Mk6rc/w+7O3X0U8g6etOlIfVtBPfhcFVkIropxFhI7VDD56e+S0OZFR
7j8K2l4+ysyIPQjJdDREAa8eGFcS5XYkuZI3xexwvw2VCou4LGkpHGy381u6COI2
m61fQZ5Ng7X3L58qjHF37zjMd+vzAmu2BBaA8OlKXkTuNKCoz5tDytj1aCNFE1+9
kg9fVI2k9DLx0F1JMd0DJ4cPD6CHcKKLrDuP4q3sqUV37WcNEHD0p1sF4xcf7ZK9
PHZ0lGA2U2jF1yWQxWsFsPEeP58KBfAstvF5Tb+PWcLqSMn/K7IP3GJYejwyAB2x
SwpFyP6v/IFAId8OxsO9RkvzxE8ftlLzVN4QurGwecWuL0CMkb5ngdiT/C2UCkxj
9rfvg14fgWTKLcsVDsR7CZO9hOAg7TImCtDFaiu4nW4ZPD9ZTN11oCa/B24Cq/5H
1iUAVb7HraG7tyJ7cLnFB7zDRW7DE9vd/nUTmPZV9AozseomIa4VB72Bo/uMZiMk
gqshjGT86jshByz27dKgYJ8io7/2nVklOkLsJcGJyZuoH9U8McgRgX4IV8eWd4lK
3h1/heplg8LTQSe7Aj+QRJukl5yTAtXIEB+GMrw65ulVypitRZj+dEPfjNLeiViE
X3MTaQB2dj/s31blbEO008zTeHER7e+4/3JmDumQ00zPy5q820MsIY6GJ7TXaVtH
nGqTvsTkoeN/TTW+9tS6/OcopDUh1se5Kr1QWlV51+s0jYgZdf3RiGcm9//5LjcZ
GHoWwUuR/pRPlbJz2lCMlWJYSelamytPSIm4+bB/FztwIbn1y0p5o0soQ08ciLUk
WFj8Nca2ZFmbnQgog36Mhf9X5oXrkPmOVunX02bi5QM+Kf0MivYKw1TYx6yQtlny
QqF6gfebL3jldKYLnGVdv1hhfEU+U+GjHpAvQA26WHUTYTFNHLVW4XgX0GmAwegX
QLeWPufPs99GP54/vnLnBMbdsF+CFbqtFE4tiMaHNdXTEkChQNryA6kuqcVUI2Uy
jDn9W8VH5oT9uK19tCM6Tv0SDRn4FJOPuHh2WnoEoL5zIswuu35R74Zp85NTRzco
ze5fEIvf58JsEtqbT6snDYhRd2U8sSjHuxbw4lSs3is/sZa36Fdhzk935Mjuj09i
o6678+MCwLIxGhoDfZFcy7eDnDhKNqMTBCttFYU9lucInS07cuykHr1XArExnm/U
GBFH0huKRdeKe0pEIbtjc97awup8wxA+p9xe1cnU2SRiqIk2AuE6uSIlMeNGXnOc
m9oBGfNSvbDbQR7YG+lXrRO1Yaib8IriBzQO6aCQXrhjrYxM2To/kyyNzbyck+ME
dPCS+kLCz1stit6sNkgOnkhv7khTpT/PDBZpTO9Mr1eqaLjxG/1zBBCtI5dIV3dn
JbA9Fe+9gbl17RDtfpaaH6+5P/piEGomNwSqYIGiDAhea5HOmLXiA5oLBI70LrRm
19sJnB6uMf45gD6jpDGlgJgM4U0CMNb9gSRgUiLc9wQQQThV106cB+64QfXrVqnM
CyET/NE7yx59RX9TPwNnSv92SH0BNIZAhRennRqA0v2mH9PC1FmiDSG9yKnk4maq
0exzuDwENWikzRbV0+LrOxylrY1lx5mjJh1e5qxD4E2MclRGhoS5zbB283tyCfPD
yQibVAM67o89U3fT9iTnWkpNLFzaTm6tCkIiH6lneBxCVqECXA9qM4hambcUmmHN
EnejzR1lEudq856OD8oJMZU67hmP/Q1YE7yV5r0Mp+NIPIR+2x45c+HQ3HgnZOHU
G7+dXpvjG10MBpiHjOAUWIMYHiQy9E9fZGjcJcM4KAA2ikvGkTyH3tHs/doM3tX6
RHyDtlcWHs1+1zFawx+XzxCrn/wvhzmXO5d1fI+hUSwKuJTvIQKG3ondlRq+KA1i
r5MQ+wGR4WgZoeLTvga/N4e3S4pIeKnkUmjk1i9Lguc1kWDl04c8HINicvAOivoy
1K+j7977h/DnXOXwaHxOPZeYWhl5SYzbaXhd+jngN+hJF1hYmCCtsrnyXBU0KOQt
D3j4lZqPQ2S7kqT0923qTohDzAVCjdca2phmWnO93Bli1HU+n39SIUTSIxYLzc2J
iSzb4yrZzETCo2ehL9Wkn4alHfYeSihz414/U8xfT7VoHrmgPI2xD8qLkfRk8lKW
pYl2LixKJ6Xr4MeoHW6ZkCWpZeuMJ8ApOWEYdOY1I09oxpCtxmOdyye4G1H5Ql3f
tDO+zAesV51zVcUZkGCyVKlECgZJ/wkb/0GBPv4HiQOGT8pDHdccB4X2BcttvMSO
d6bOrlrGh2DeaPtw4c9VHi/XmIKvugoVr5h3FIPOBGdwEGrwjRJtJ9AEVafNDxE+
KzG79wKIPPHIS2KvB3viFTPuyW8YWIPL9u5OHsMSdqtzbv0ZFbNCCYI2um8o9d+b
8ePW9es1H72DcMITkik8oPo02Ofu8Kg5j3Yqfivf6nwiMiKGAh/PaIxHHNSPkCaB
ZNap5lhobM3bqd8nOuLNVKu78e/oD33VwqzjWNgiZhE+0FrWAoHYBU2GU1Ghb8wq
WcmOfciAIoNTBU+5hNM4UEgVWkVIG3jI7XipRgQR1Xd8Mu5hYx3TMX/IS3Jr4OKl
YqML7vm/fjm+pCH/rAgKYXlWnA97Q/8GRnOHlhFn9hZcV9OP8756FaZ+GodRfwb0
LsGaMYIlchejDyQqUxiuam9khfS77gxkSYhSHaldXbKPDd7ySKlOPZI2NWfdYm9n
ks30Ix9eQa3jgjddWpjRz/L6kLinGIMJCu7v/ExRhcph3Opo7Xf2aIqn9xrMgh4g
D476xl6XIpgpRsXY0dlNui9iVQ/iEKuoqeEJLM7l7DvY+iJwcA7Cwbs/qvzpZckU
ZnJ525moB4srIaGatLohdvzZPkGXbuEApdwC8Arl/b1ULri7H+79Hwpc02Smd00z
6TEAS3qI1eEY3VkgaiIV/LE8UvSk4dTXkSHHKQ7yHeYTBQ2TFS5BGH8p8VU21HFK
wsyPBU9uqTE9UUXbXLXNsTQ1vLhFQrh1DqQEcYinjPheYNPn8xBQpUZ7Q2XPc1Bp
7eIERVxnUXXyl74vdkDbMKDufX1a7OHxk2WK9tGdDCifHidouHw1SoA5fzURd+2t
ZkMARksZyThCOWoRlV8LoBpxOJyexCq1hFCM/CZliEzlJTNLWcTjNIC9/Fqs0ESi
ycn2ZgheZ1T4lx06xc5Ey9OtsyNUGfUDCWjwSJiFTNRz6jsem4QcZNr1qqfTecBp
x8rAzDekt2iJiOO3s7jfNKDGV6ToGh1Xi8BvvlTl1CikPofIHB+7UeSCcGoVtxsy
Odsga8Bzhhaf44QFVDe+mzeMCVzfGBFCN/du3NkjAHZx03m+8qprC8pVqTUZofxd
5JqYDL7fD9/tM5Bnun2pst9GRGi2n2qF3ws4NHP8jTpTPZavsFGE38e+LqD8Y6J2
gy82qTbYNv0SUxQ07EP8ndalxtZMsoXHXJ3v7VthWc30ASs8W2VlVJz/hBxJwfhC
8u0VuVz4fyL4awhLuM+6UPckRYCcLdD26bGVDZPcBsrRCZesM3crjIxA2xkJF1p7
Vre+3qc64HWKN2EfqHW0kubI403wt8Qt1boDjnb6cTFjxZDyw7VQOMkhXnzIqyCW
P98mMm/T2kIATThf1QRaNH0RpB/L6Cr0+SK0uT+ILpN80hCMS9ZyWjYKmS2qqnzO
8eIRhYIpZ+Jic1UHYyaFuEGc1fJJt2abq1veg/kxfsf8JoOO3kWB2XLDsYUddlzg
TxYNNhTNDUo6PKBUzutZqrkzy5Jxv/03eCjOTiYz1uNf0ubMdNqfJWlxq+i7nFZm
iZdMgOFVl2BSCVwCHSVlDowf+qMGKOkGBPu6e6NDobAH1qbpOTo6MS1grytmbhvg
B6AEF+7eaM6S/FwmMC4JmPXTFeb63CA/HdOLgW5tPpPZYL7OhHZX3ebSS1LOenm1
Ph5IbfhHY0adistvYTueoPar6sWtT7nIW+F63B3A8MRS8F05i7vyT7dNSgEOLHHb
10kyRihQavHidYy3GasYLbRp15d+Iyd8SJ3a6TYFuP4gDxOW+pjDONmYxzK5O3jn
tf/QU4M1HbbJucFTTR3iKiK8IPSviGsv75kR275Aab1oOOfIzXj+Nhmakj9N02s1
Dky4PDzo5hegoR1l/wV4lCQfvmrIyr6aQ2BFwxlxleCHaG2CqBgouvt4Q3Vft+oz
n5oWnjQPgsNxrtHIkFPRody8Z2JBcIwd/8RrPUskGDj+pP7W44yUGz6QFDvPq+i5
AKmiWWpRF1wRxS8Zix1mz2UCnPJ+mUTmnvraiwVyiR1nwK0FpjUloa7Drzl2jCiK
r5yzf9NiSV/pBGUsw5l9oOM4coZE/2TXZ8UT26lVwKr0eD62Dy8y6u0dwT1mvQrv
JPTGRxAHgn2nZW41I3fPmkZPnqBkDCWkEA1i4+zx5aPiUqQpwkc4hUpG/4tTLwJS
LOiAPQdhkqphgMkmdZSEbAXF32vOeCRJVkxR4tJ6skGsaT72OvWZVBK87D+a1/uH
Fq7YTE8/AqreBRtWTrb+bWIiKSH2Lf0pKy/1ajHSS66P/Wtcp+rVnoIjH/6Sb+bv
I0T2IdkRD9Q4WDMeYko7TEyQDKFFBlBGrC0Z0umt8bkIl3TlnjD5l7C5sHhoSrp/
FfFS5Hk8037au3cBXc6lP3f7hQ41lMERy/NeJCqBvzZ2dhF64hwVhfgvH5rDLsMF
RDrDBkJWCMftxZwx9waBpfRSSkpNG6XSKjY0SvlNSkiv4sALHC3CKHBp3CksLweO
hxf4gdc2GLZlkeOlZoqaEkHCkPfkqD5e6poMXlKg+/llf8g9cxfqG4xJ403FhfiI
VHl4xMVFgMPQYij1DO60tIe2fLZvNEzx16d+Lz44l5rwsWyLwWbJI50u6mjvjezi
EG/9kjPQuTyPQ66TOGsjw1Chfk/+uz/4Xb/n91xw6xkMj+eZ6C6f+TO+ZXvLxHwu
pFwINvuJpzsOp0nzCUNazXtZO+DE8NST2KtO6/XfXrFW0XfuRsBw/CnZLpUxeoLC
0MY25erioJb345/pHPkYPYrfF7EkiwiNxC92jvAyxDq+EPSEHZrFIpf2QgaV8UxQ
n2SqPGyGx6n6SY7/EvJSHY7Akew6uGRNhzCc1UuIit0/82xpbNs2wdU79vvGMzt6
Hc1aWdMW1H/BAF2B0ePylP+P7YTH4VzizB1QztqJ4t50rHgSpUOEGrzxSTf3JGve
t5YB13JaxTRPpkI55LtbZMR429jCh6pPQhFKUoyTG2GUIp+Qn++CDqW1vm67yYtU
jsoNqrf4enWSsBvMxu4fsgKHezxvwk6Dek3coFQQO9ZeTnR8QJb9s3Bteau/m/4P
4V6hNhEGAkjDUcbIkEucO8FQ8s2koVgvIkFQqfvyflDepqnl38o7QB3mgUbRjPgL
Xh8UM4+TeJ3BdlMTjGasT+RE4rOq5/nTwaFZpPG4NPbzn64jzuqytl46ZCd36Nbl
aDL81TrzX0nGH6ZDiEIwJ8qMzZBulYJ6W9wvvZaLwQAl2afI42OQVaOuHtszcVr5
Ck+xstlCcW235UvvvnZcSgH1fsJwvdOE2jAXeoVWdiYcFJ4Wti6/sUhXB2uM8DEP
An5LR2YljS+hLJofvp4IIs7NffMGTPMOqvTYXf6Su4okQ5cEg1gMWh5vnJQce6GU
IlcXbb5J0OQOoUALZtzyO8/P1WG80bQlk9MK+9D79FsnlIBX9YzV1JGJzCovrfgT
Ec+eymbl1rwWVBhbD7/XRxiD2GCqai9pYt/07b26ohRJEcaPrwBAEHNetuvcCClC
aYcTNYawZrZEOOOeEqyePu6b0Ru5mopsDkEbejAcpAyJA5UNSv4aU4X4U8fPONTu
QgEAyPk1kt0kXd6alnsaR7z0kVca5COT7vt+hjEAs2KEw/PKYDr3TgoANCbJ329j
Gx6k2lkQqfpIZIRuTgzNr9DBmTPbLYlNtfEVn047QlxWxw39ryW53by9x89Czxk9
sHGAQREnElsHnkK8DrFyYyfdH19Et+7jwh5l+4Ds6rc0OHT0Mg8Cgy3tJ7Nap08b
TQOQIXgfybR7IfnA5ZRZGw4CxYUPPZzt7DeC/WdYroKIGK/yCeEPfH2Vl53fRavz
3qSnGjXE2oBd6Kt8sM1M+URnvCoHuohSRvwNGbBDZx/dvymnLGbO05Uv7M2/C27G
2xEAGUkOuoD3uSK/Uxy0cUVl5rkBjb6P7RRsDHDTpFmfsiWEHCi5wU4EpqEj136v
X27EPvu5YQFlbrQ03CYBbdcDRzoKZ9994/8PhH1r7U8mPvWAOE+y1KnNfxTN6fh1
UYjZGdxPSSI3ASUMOXmILDxaSdRCQ6IRKO4rSpHABp+P7Wgl64t2uVCK0opkUAqH
zjZximJeYgViVUAuXBX9xC5ePVOxkOBWaO7FBokTTkn5SQdKSCBrH+33C54p61q9
8oZNKV6l9o99SZNJ1M1rxZ4MYZXbhnTGLG/0A+Qezw89PcfOtB9TWv9pzxtRxBev
A1PY9fDColki0tMSMAfT9TFxWMwHPJhaGLiLrm2IHKanTtVk8LWOMDUoTSUduZh7
2OL4aYdHPpDMXCQXZXds9q42zJ+vr1PFRqOFkymFutoXctPy5wL8+Ug2VKSecolD
LgNp4eYEyT/SoEyUd6qVzb6Nn3IlPB2ZNcKA2prDjQKKYrAzMejVffb54L3b670e
I/2e6sL8ay1iJi5hnORH6xODa6QIjrqIOF7AhHfe3eW6i4s8zm60329Rp6P//pvj
nAdmJ2tPQ4hipbLf8DhLpfdmmzONaCbMnd09uiug3qnm19FhGPb9LkKGg9fpoiy/
U80neKGZt5jjHser1iXNjFFTMY9PlFaHHY3lX1LMUckiqV5ZVWo75rRRrBSGSOJV
4JiFLV8vbY/QpUKcZPNiTYMcZCOmB5lUcoGmbtxVa3XmD02rTFM1SG8rnolVxSIX
jwBtUKdqtfO2yUawV0ioxQ6dxTEZK40n/Sm+Amyc+dSivPH9y3sTB45P5Ep9YKnq
pOp2vXCZA6Fp8qlkVr68/3msph2Zxy6pvt3sS5RaWmkwa2ram8wu7JWNaWbXbO1d
+cCil+6o8Ztow76fBxCTKmWw0yiBeLATb/0UIoFiehxhdTlX4fNgpm5CwldZudVJ
33fc+liedPvu94NPdUqVcG+As82O9M/KziaK+jr3PamlmL4Vi6yXMhyGSSkMGy2w
UEYY2Igo3RYCWR12Xmck1Ou5JXwcUyLuPBCrrI9COqARLmCxkm6RJlzHQRoCm6vU
NI4H9OtUrfmFPPfNESxEDYIuFqDyd1aYsLf/rFDnKuIz1wfv7ZqKiQaCXb3rlzzO
p4QehWJDVSlqh9maXYcID+0CAR56wMrUzTMzXyMlg3qHVRVoqQuYJs9Ti4G/81df
2tjg+PRll7VzI7V1YznRyVYafGwVK97rJJfBinvJmZAvdGAR4KFaVQ+oBGKPSBfR
EOucgCUHQHh5CrNUbwfTktBxlyHpRRSXbDKlsNA0gwplzfaiUtyDFq8LiMG5/abI
Dj4gyLnJ5rd1dDMhmNVi62lwpj4+cm53eAiYUCretQNk45LGIb3+t6DA2bqmcJ9v
1rXSwG+wHecOa8F3aVpKgFeqth3YL3GKt9i3Th7J7ceAY5okB8f3woZXjRIre/i6
47Qubl8biCD6nsMB5gwLsJhhX+SWoKIKqCjsUsHlo8buIAvzLu3qpXA7fwi7eX09
CQ3zrXjCjuJNfYr2Wp0Upm781nSMVI2LC6lXp2iKh2EAn+poOp6OiqQatrerefLn
f2WdRt3p5UX6v2+Ajdj8IFvECLDTsjfp/4SVuuvF5SGSEDzoQIYDxfohc60C1Ilq
DtUWKlCud2tPf6AHU2hS38zXXeHZibRihZCj5gDBvet/xbmxDVCQvEvOqE497YM/
/YDfztRGwussVCC9aK6o0Edd84yhVFz0THRABYfOrffUYoIFphLkSiSEVeKBNI64
fWJAzy6RLiSseVP8Y8v4uR41v06dfL7KS0iturrLR9tP4TAJv7uPaGYijjxNR6Df
VYnW4O3i1PRLZpUlNdDfquuPuioImsk4jYTnfyLfWOiAgaH2bkT1pZ3Q7wQ5EfXu
0K/8bj1ujIZ1wvOovUUiRF6G47354lxK+ENQP2F+d+2KY+wzFXJoQxn7s7rKPVx3
5QDZsX29lVN8cz9ndR2faObXZe6U5K9sXJi29zp3QJb/+1FT6J2IOtjxqxMOrjrT
yzNbQjtYGizPiZ6Aa8b2MzUKApixnTAasvifUg7Ecps403s45l2X2bxXjp+rsJ+f
c2Mzu1TUdmxo0SqiKjAj8yiQ5qm07iL3IFSrDMpolLpquTDX2FGVmjnpr48w5ftj
AY0jCtqnU4G+J/UaLbQzXPpKqvhzw8foKbQSP9Sh0J+/Nd7F2G9SKnkEW4051diD
cKxwKJ+vU9qR4ynRlKp+EnvauRFrcjK9yCMtqeuKNCQjsdqooIcotnjFuot0d9CE
wJnPOetdEcp5mj8k0m87brxFIrEX7gcS0upW3TTlZ2SyJombh7aZhRozcbK82ZNW
8vqKRQohBrITsYOswVxSom8j5wGceq1ef2BHO/PNgsjXX8DGlZJWTciYi7O0v4EW
sG18QOxp1DvHiMkHRFyJM/8oa9F8VEnXD3pPj/HrH9LCFW9OQrBMqdKlTEHRgm6j
DPmAH9NyTDw66vRCt6hjj0fDsFL2oMapniMbLu8MLB5KTld3UFcBkdSAo13qG7Ve
hpV+uHUwMdTUINXq2axGgB6ylRAtR3VodGHCAfSH1K2vHDrCl2oi7/Ql+8cuUump
md9cRG00ZMDKJwuB6BlHBu8mDMnsaT7RvnYfLkm6knNydTVrLWU0X88LpdVvybfa
TCRg0nHr20fmG1bOphDNbIB2Sgg0C3vEIFCLlnH0V5JR2nJGFKLPtTa1AIqh/ywQ
ItwPQhMH3MgppPiO/YsMm/0VsICrPaR++X8WOVzNT/7GQABsGWIea2Y5oAw3keyN
8ToG8n68mLXbycL+T7dt15p3zCN+5pq0M6xyPIwbcuQm91kX9cxzL2x9+b7ikKHm
abA+b21k/xhm67Eb9OhxJkfc6sqWTRTj2f/2JH8kgFy/5FXaDR+wWRE+dh2s3yq/
Wifcv+JKomghFUP/HyLyuZWFJl3NwnaU6xd7YOhxMVNB9scwR0xO2iXjM/8mCWhc
c5Gas7WlAsAm0ibPtF3uGcEoPXXcb+y1Jr3+7CjszR7VayQ3+awyjn0nq+qvcGYw
fc2RQ2zCmPxtGZRmjfH7F4QpzyuDfo697Ub5ZbsKaac9dYUPuXtT7DZOz4RlO8Hk
Rtx4YlYtHzBBtjSrUei2fnLLZFwl5tXBbay74rPQpbPNsdOdxKf3J7v6ui/Lx7QO
+yW3v2MOgSdOlpiYmeMv8ZTQQilrNAKvlAisjCvC1GLX3cRq58nHQB86+NcV6jIk
Yir9s5Od4oqJcbqIuuFE380JoK2t9Dx7051+UhyLwPE1QX+adklpK89/5pFp7GqM
drSZYv7mutsN5L6PYu2Ron0H+He4xW1SphM0EenGpZsvuIzro21KHFlfSCwl7f/7
0Bid087xPSJYwHQW/sQXTpfbohESMESKjZYS+qflyGr6SDaoF81lnW8mwLeC9I/F
Uzc+SMkXcNaydB9BaNQ7ipn0ub+628befwe0lNZJZ9fUTDvnSkVwjT63ahNU7vI+
/racZlO/BJGPfKmZHB7iH7OQPggw52ChC1EzrnMAUXi2t9xsP7TKleif/HdGR+I7
vLH4R/pfJeKej0mmyiNbulQPc6tuXfabnibqHnKIZqnnPsXzVCTzbqmOArMV7GYu
fWTofqxnRb6KR6TbUtAKZIxeLssYuOMIrJ20B3qhmrnnB7yrG4gyWa97io7hbU4p
PjB6USIRF0geGivoSTS90c7YWRsMRm7Alv4fQisvKXTPYRfQSi8NEYvCXQHoCJrc
oaIqT/3efcaGgTbwmj2EY3e8rdWfM3/KXRuZVfWnvxBOxObNIHUm38fiJ5gtspmK
EnkQ1gfWGC2cbYezyLNyvXqONAj6LZT7hwVXqjeEt1T/sc4DlPrSjtDdNhSKLV9J
25PwRK50b1ntX66goIFWYxdsmXV7R3PgOhMJQWVkyc8p3h4PiNZs/f3ojnNIQSLc
9pt8W8VxlP5E0XrXC+Q49Oi9ayX7vEXxUNgXYEwgYfBm5Otx2manzvgHCnmDkscc
T0RkVwJMCx5DJdDJgDfaHKctiID+VtdHAcvidPAF57fcrJA0h5wwWegigem3QDE5
oiWhhthPruohrHc9XnUTm8kBtnodIIqrLy4CuNVT0BZxI94333QrlXvs7b+DT6R3
MDsRA+MB6S7RKkEtIV9q6kAorET0lvGHuLfQ9rcxFJzsf2r8reIz5MAa+7ElXMHz
BGybgFt2V91cPJ4gTb8nt2oMwZQl6a4LRYdE3s4G9cOTIBVBKRh3UZJ0JsZ9t5bP
fxQmiFGAMxCIpA5kAkLABxLrpgy2rSHpt9QGeprdGoKZw1LtFZkFF92lQvq5DOw2
RTP+a80VH1jJEbOeJoW6/9iuFo4tVVKfZ1S2P2asKyVVtV6V8TNhUoKRYmW7dy2+
LD+lfSgevAQftlb9m2I4x0/xpkBo5jgznmZm3H/jIAKlSo82BkUZNtg7JnUQpHbV
XuTd8z6bkcQrO7FpS9YtcaG00QAes4r8djK8ZddpsrYyM2YL8hQNo+5wh7hGO+wg
eQDXApRf2U6OAdbHHgvodJWb8h7U6HQbBv8Vzdp8fpnwfCcUe4Vi053wi+pQ/8rf
Cd6OEnxv5Fal9NHrLggL2zDOjjNCU+ZcX/Ono6eUJtZpAJ6JkWAfZpmqe6cbV6HI
XKrn7z51b0/5EEKpUhY8JHmt+r9duYuW5NySx6IjpqnzyqnqgqaBemoJSnED+Du6
hCYfBSitxAfGwa808PXu9Zgo6GGyuE80hvfTSsjsRCFTwmBuVYxCT2Dpq8mj0n0v
cwTN61o5dRTcYTmuujyW5Sp8y4rZ+c+K87S3Ke5SzAqhr3H+bvv3ce5KeMdJxSYH
rx/LTtHFSiT2VTxbVzM4rOGpDf4pC8YbNM+ALQSM433TrAAU5fJu0Cd8MI7IBo+5
jyqvh0GdQfOF/PBwPgnEP5lkc33uf6it99EO5pD5mfj/1Q6BQeqGWLdItzPjF4x5
FFLj8d+BZUDDKlnGTFZVHdY9TO8MWWpfw19KzR1I/HsLd1YZaAUF+YvVCKEFuoVx
mHLTeQLzQ242VeQOJwomOpD7sFt/MIa0jaXvjj2I5DmtswDUlqhBfPdjMuE3s1qq
PAHG1OGdKLMIM7x2wj9HH/RP7rB7dLWSLSy0jm1KKglr4VglQoHFpWeIOD/8Jh+8
x2ZWT0KQVMh+lnwxx6D+6+srtCsfpN4wz90ODX0kPZVj1WJg6OvQuJ86N1+zrwba
TbX4CoPA1arwfZUkEpVwvP7JqZcXUzLjY3bikk5FS2C25AZ0n6+aKUiDPO8vNTZy
hR8vSD+/trrhj7w0vrZkBpuT2SfOhGPN8SILCXxtjMs72lxjHTpw4D6aKwM8nw62
P6FIhU+6A/Ot78vTkpjUSRGD072RfkQ2/jvNtco9oIIA2XSxC76JNp0uC4u1U/6a
aKqcAL90BzxCkgAaRhr5nErS1EAjPGIMu02FcB3uvxmLPDIg6I54xZvvBvAFuyXT
lAX1vVG56aUguMuQcGfXJkw4XjfJ/eyx/+53wTK6Le6AW3h1Np2taeYbaoJeBa0A
iV/OYVCscGT0LbsA5EKEGomw4Tj1NIqg/et9Ftw3cppMEp8v8mIIxWt9ZxqWaRoj
U+p4RrKPUUGpmiWWNpJXoUUlmJdGTlAwWkgWoiTVyNyZsR01C4jfi9j//bfZ1HFp
nXH31AC3w8ZuDokbz4cATzCZQ3hZbfryb+OT7Hn8uYn/HFSXCMoF/BNMHE2ULNTt
EpuA3svgVM3k8kyY49Ao21zuSqwpqjwh4/zTQUlZPSfdo4LDB3cCtSV42dWzk363
mr3X/drScxTQP73/+l+muCPNzGlU/8dwB92HHQNQtIXgb68V9zOmMAW3//Q2GJTp
4mn7HYgpvESinl5A0WZ1zLQ55o3fCRq1U3DYgnxKOLR6QSaBMSQhqJRLnRu+gVc7
ZMGas2h3u+PDTQK71/BcfuC37XfTlWTiqoDUudl7m9uTZKS24uH5IaOMXQ3wPaiQ
v0BvlvzWfUR8YUXd+CShok2MliE1rsmil5Qe1Rj3L/33qbnOW+USGp0+nTUwDICS
1KwRYnWJzkRXldS6EQQkhnmaBFh1r3nFLQawCbZ2VM+Uec8vdWjhB+kJI8s6obP8
jw52rr/ubrGbt9fVA9Z2JJK+NtbPtIR/uhMxZcgsvoOPPX23P3IH7j2VmN4Nixrl
LmFN+I18oiH7x+Fw/CzcdJtXRDPWgSRXNS8+MSjyyue7Wm6lFnUzTvcRnA0vwwBP
Q1g0T6H1LVCXqQt1gX8d18I6jneaJ1Kzy22F/j9xsV1C1cUhK3jRXpXFRWk4FKmX
ywvlmXUgivkOL7poVVhUJZrtFtrlUeFWK7XDHc/uIgtbjomCjqhConRZacNFEcUW
T3fuILUfmYoYTU6/WViSvhb07tehXsMjm0uW2UBMCVvRL5pWHq+8WE221iRDaYmp
bm2cjt2Saq+KtJ9LXHB+Mdp7yRkfdzYEcAYdBtfUEhVJnaXIpYH9B2RrSEFi2vqb
rl0HkGfEjY077j+TZos8sfCm92EIHPrODz2TWPiEjktPK8vfTta+orjgRXVxQH3f
lB0CwKPPGoTv9X+I2zYyLL/7GmovCyaH0PfatuXFrpeRysRC3cQICACC6dRNwwek
U3NocLEVLTyo2MliDriR6S+fnw7nPA8ULFvDSjRcQMh3I+xU8zopQz95XTk8ar2e
1DK8YVl42gq6AESTB1HdmQtTBLarCPWDeoBXxueGNKPlPvZM1wkaeYUDq1Hn7Ic7
yp0fUJsMqciTkdIGA56rhwJo8TuEAhUTVHCxu4V09RJUCqg1G9b+VGHexJXMuH/D
dRUe2w4D7HNl+7JOZ4msOmdgkaxS3zvKU7ORBdyonXGwPtAPDhV5jKDMaBWrgnIv
KeOM8cNbBnbIm2/aQj4iagq7qz8GzJlFN5XN07KthoGMosfiJSCoSPrnQmY43yGu
30KzKajlt9nDBeXSytRyy4CsY5hP0YnSr+rbt0UmAjZp2OPzYW6MGLYTdkj7vdNv
xxx4hkXTVxIFGrInkdRkixS27iN24CyIC6Au89HeFp8aX+b/46x/5cud6h4ScAbE
2XL6HAb4Y3q8lT3IN0LWzhi4lw9eZcGUpdO5ILyKKZ5RRtzj+5NrFHFKUp7OKsVG
autF3AGDeM6xPoxY8lmizQ1nx8wLZ+ILou19ZHCDlItWcv3IgKkOUuiZoIv+coan
T/1dQUyZqGOw2m+GqwgTo6Dw97uIYmo5fa0xlY2dVihiW5khjkf+D7cvjOQ8XgCW
yvW9gTlq24GiqGrZHbh4NxVGr/b85erKCpSL2EuRU+4VWt4DhP8RGhi52nKVHCBp
WK8EdstgckbZUitwtBd+tOI6szhmWqvl7UxRxsrQc+suLDlQFFogRXXIqvWzyA/7
7u+ItkgZajuW+xhLRSGINkFttUkkz6xQjXYM6PlrsVtGvFbuYxxA5hpFnWFCDsGG
vq08nv0/k6CNOmeHdl08NFAygzJMADLt3VTo7Sbdj4o6wLtPakWA5ZRxzDw3bWQd
h8LB026UtQR7KUoziGcLZg2+XQuKMzbiWXAstm6HKUzMx+IHiWLZ/DniKL3OyiP/
dgZXJoRltlHFe9X7D4mj0Dc9gNJDigZ7dNfGf/PFu5WrbuCepW53SQyxFKE83AXS
Bbb8zvkWQkzoZ7Swv2WlacLJatIYoDKD785fEP49vjRGevbu4WD57ZcnX6YUBNEt
sRadoFzRl3TGigbIWkSzpriosAqLNs8iczTD4eZFlisyhvV5UzDh3LTr+UZJlwDI
mC11SBCe+rlgEjR3X+kDt6VoqJ8RI0D98ApEVhRTCzh1QHRAmJ6vdf9eeV9nKxiC
x1YXV2GeTPLSwbocv6YiUMXOiOLOe0Poba0Vk38jmeDA5phKLQuRf6+m2lMoxzlp
EX6KVanFNyAGYGoJe80GDM0HTOiTtXleSuiJ5zwF8tEnTfvD+qXuWHJW6d+62kgd
58xddRiwu2/SjEo2dcV/z4QKyGyyoj6VjwWEDI/4zCtiXpUyUYbLrWbRcDw+r05R
VNMej8dVWyC+lF9udllsCWL33JNV9g+fNWjAKzmM8RnlCLr9bfHytrMq+a59WKUf
T0Weztch4+J8sCQvQ+Ojy8GIKP38On4FUUgFCcZQPkxS3soocbw+/yjKb1t/Bhvr
oyLr+ourI7SwNvHUc1rJ/lQMqGrtPnMktl7K7Abo8gz5K4xNzFeb/znPyDPJiRaE
fcDkgiyRScVd0JdFZfNn6CEnAKMix9KAsG49sd6bR0lXOwFwH/YCtkBXT4kvnvqJ
DMSW4e5cJIG6+i4wVZxhGwrHZRMou3yQ+JmchIo4DwZ089XlGdMV3bB3X6l3Ex6G
jpvXL78joxSaAs3Sak+S/yGxax78kp8gv2Z/oA5egclZ3tg95jNZlb0Rm0u2lS/H
7eSpPa2rQLX/e5PtAWoBPVoknok9k6FT7zlaeqZoPshFTwV53C/TYFzYC/i8zV8g
mWskHxdbZePZEIdE4Vb5696mwlcUV87NcIPWWTCDBONQz3C8RH5RHBuf2LlISKJ9
Q9VTT3vRSD1nOz37PJLOW2CiXh0hVcWkctQKlnaK4WVFdvVtZc9yyQuDMiub4t/v
PgSfLBkBKElMfV0qmgiEb7r4qYOy5WjrBCfokUBXl+eonnbMjW7GLMeINYYggkVb
zSsIpI3SOl26x6oa52k4ixVfhkoQloeTYer0T/rLGakj0y2iT1Ve1hiHh86ShRCS
sgxalfOmfMPyPjXsxmfU0kHjSJUFlxKJnwlA8IpFHaDQontMiKD1OJe2SXrz/Akg
e32eVdTVljBlSTrbeC6hXlO8wFmwt+9S65jZkdAq31xIgHHapr9d+FtT1k6lYVfs
EX3Q3GUsw4xLACDnHIp7gR9nh/8frBYftx9aDR/OOsMeDE/DrxV/TauxZA7Iw28O
WpfAh1RU7/DxW8HLxsWjEOTVE22Lx3VyKMEV3MbeBhMpurvAMsuCSUx1I0xt9n2s
eRXUGoqSKoH5ozSALrj+wRuMqHPi/OiLBOCwwVcPs0T/woaKJpY87mA7cfXJxoUJ
Kf8cmh8mMK/M9PqD/PvCosNi8PejBEhVCDLDHGRWxDSSOVNklqc+XnvQtKqxfTcN
GyiN8rNeUNWtOlzutQiYqR8ID21JWvInk1dejW7XE+JVFUpUjsZ0Mr8qwyXu7kgT
sGZYtAmLJxBr3lUC40eVKKylY+XFrBzGlDM5b0T2YDGeVynyzJxnpGCnhMW6ci+e
fZBfUS9psKGQ9IDJLK7ueU7cyWcct+mkZeDUyq7ehYTeH0lRlQX6OxRwKGCsQFuc
saAC7n8kI36tcuY9np7AITdS2ZplER9Ed6YZWmVcBw6x0Y1JFxKfIB8jOXlvNmTP
jHBkF7J+SgzO3SqjFnVQMy4xAPwjsKyiY6NR60d+HxqcxHpMw3xlOqIFb2i4wzap
T6WlIZwgBj90PFGRFd+VIMyqJw8yW7c2z6ye/F9R7xm7NMPwxsxw2IldpY8Rpi3T
4dvJjRyyWwRVQ7gJyleP9TrbHl13i+On7NKKkm9ufpXbM55iP3Hu6L8dR2e8tATI
9ZQZnx46FF7zghz5UxQHzss39jNhaYtN5EDjkny7ok2LjR4LdaeqoJGKH41u8JHi
yjvIQ4SmA1uOLej5gj4XXwzgB8zk27xsdT95IMtutId/1NYwOKvTmCdsXFWWalpA
TnewQaVK4Q/zsUW+ea/D5CKkLt41GiVrdQ6Ox1SJEeh+Ni/d5vZKDsD1Glfde62f
kbB9kGKVK9gAdZRt/wzVdnnm8MM1fUbSdTk7SZTitMEwu2KwMt2Wqd/2iFf4e7q+
8liCLZKfwaY9WRyRelYxnXVbbhI5crU9Gf9bQYctkxmZVbba+NYKLfRa3GqnLGBs
G8KXjuXM8IV++qmYIeJltfwMvsd5qkic9beuhfMiOigOs2iUmYc7DhKEvHC7MAEl
ghqkQx+vWwisfKSpO+tPTEIm71SzS7HLDFm0QsPJwJix1yjn45JnC4gU7AMjNgCY
A9aRgqQNtDw/2B9c8zBf9BQ0EY6hqnrnSEhtyv70yodeXPdVUk+C2wtTINnZwxlw
DFzlK/yBzbiDSbcLbEOqZb/y2Gy3HG7rR2NEDgaH2jqd9EVK8HmhZwqfXYK+NhiH
zuy6+jTWm+ng0FgnmPcuL6znK+3uGj6jftYOCErdvQBaNvW71WqWC0jq359Ez+We
TZCNHOBZGc49PyA0RLCu+zQdraQ9mJzCu+WryJ4yx1X/OFjE/gaaErfSjfmWdlvx
00tmJA1BGBs2LNDko2xSNKeFuTesucf9iv9A56n1TrI8UcLZRjFZFMgE0iWPG+3z
p3KwqLLNJ+IFLDEeta2LAF5Ko312AWwVX1EyZ+Stu6K5fljJ8J9NbxiYtoDCZ+0z
B97UsT9v0Toa6hab59Ja9//wCR/ynZcPrwlkcrKD5MDuEWLSJrqMN7CnsoTr1Kg5
iF372Yzo/JPPry2qvoVYgyt0LpJ1GB3IO8qnT3lyUey5jkhsbA9bmIyB0XGRBrYH
aw2h2hj56t/GUkNYTxsNBsRAxLUBQECfJJAYnr0GntPtYgWnRbGjPE+54pKTu66b
MNtV0Whh8X6iDV10yNv6wgk6GuJ8e/xgWu6vSOvPiSDvdOIlQLJRplpwOecw1ldg
z/hgGeuftQ+ZltFcgKikVunTk24zRBRjfv93Z8uAaKsIOrVPuPv7Sixx+5+IeDg7
Ra2qqtIoYqJDax9aFyDc1PniTa2nekI5NBZQh/xD5AWmMJh+z1oo1SruRGeTntFT
2Lura5bGRgAH604dFcGXUwUPEPtQHgVfx4zePPvF5oLVm6sjb0yEx9nJ4xtC4dNT
hCfggmghqW53jp3Y4p6dDFgTCJp9BILhKSr3LdMFyMIlY6KCBGf6UA4R+rLuACJi
0f4LLy1i4j/UlG6Iut2x8kgWirgJL6eE7PSvIhXfm4zY5CbKfVaBmW4PfFSKbup+
wA1ryQIXRh+5CH7SKfpjdEqGqZoh0g0NpY+j8YpMKmpAvJb+efQ1fB1cTfMCUkub
aNQoB5/2OnI2vEqFAF45eARdKhL7pKDoPBsGGDGq+DGUgMwCONPjUPYMuFpcc5Nm
h//4ezRdXeGIdq4gizFtYdcxExVz+MvekGVUrfrHldXPgEpd8m7U6YEis+rLkSlW
1WwIenk/tiOSHAsQgSjRr+NSXYVD4a8nJqYer5E3tT0uvepC6p8dBQb+4hl85QQK
c9S4Zm4pFP4JBD+aPcr4uplRuOOZJwVxJypD5TlUZYxBBd2IdZN+XUXfdBx5ovE2
flswnaFBVEGVMYfGWro8Rhz6Iph+sgiPGqpfdZbdx0Meez8X/HJAYoQm85njlWQw
qmk6neplOrw0B+NRUPePGMhV9aRbtwal+VhGVn9XacaE2PsjQH3wnJLdLPUIniTW
hg4B/+1k5UsbK8Yxtlx4cdHzBM6XoODWaEjSej03kPRHNQf0yrTk6wx4hgHSrBmo
v97fHR1EhU/+d1qNnU+HqQbHSlpBtqfXKD5fRTOpIAWZbXhIpczDqJqNVlNPw0ka
ZsRxSK7c1Y9dvYCwf8ml6NUsO46ib7KnxwPtCvxgPZVsstRLqyeDzjm8rRCywXIA
zPDLr91L5HSlqYP6U8Wt86+++wu4/rxjFru/viccfKauy86+b/SeBGlhZjb5Kkzg
ts+MJwGBs21QTVF5MbaiHECC0krL+17iEHpPJvRUBtOYQDYC3FZXInJGMbVKKYok
tj+6aAhA8VGwymAHDGN3gZryit7k4BCpadae0ul3eXTueSP4yUadbPqcCsVdb0C7
DUmCoXS1czrzkgztKLu8B7zNm/UcNtRR4paIr+KRlD4qwH+o11xwWS07+4etIXkN
tRgoQ8QKG/OYYwm8/SfOzHg+bJOtEXY5Q0kdZW9EHq5geOo0HMd2yDoPNhLEbsqQ
w2dcom3yja/ou/mAme3i9U09pRe57diClNAwpIJG+cXeB+gQax7GSbCWmFNVc+fG
CNJ35jAQc71YG41NiItUkCDi1r0swq4th23M0dVvu5/WymaDnfb+mr4VJ/dMX3cx
DvnX+iAsFbGZgteJLUtB8W96tKexpAMiPyQqf34aymfCPqvxJk1w6bEwvIWFxfer
2e4FHY+4dHRO6XU9LDS3+L3IYiDiKB8biAxcBizy3oqJ3jie4xUAgXlKIhhaPq2k
zFrjOdCHQNN9EAi+L3XsFbe7/jKLryt73NMe0nKXeyEjTxE+nliVTCV0702vKEZA
NWkVll4emPHouhfOG8o3OruUMgGWrIAewG+K8UVvY8rd14pubWidrsNiPjwPsUsD
CdLY28NNjt2NF4uR13Q3nAtJWRTDYZ+gm9qV4oIQwGOEURbJ9HFUq4Jz8PPE3r8L
u9PS/NdY3IGSHRXUwZlsC9iQ8mPw/NbNEWzpFxCHxkALnBgjE2+e9jXwp62avKbU
gdlz5U0X1KAoQETOVLFUAHaFYUH79gPjdguEUvGyQM1uqgeb9l0JDIhXAdJ4wTjY
6zQdn8CgKBSvNUpLZUABigffNX3fzfs8xGH5MsSA2ILQa/S/C+HEijdv9foV595t
FMsKWOgc0KELuJ6Zx8aCMvV0boaalTlrxqip8Lo78/0IHAfY0M0z1bI6FWQ98Way
RPaPvbmJGGDrGorC4uzuhbIcRLJ8uwt5y045MblkJg66PQ+BECyPzPhs43PXRiDD
VLFp2J4or1+hxo6DsA0zqAnbbyTVNZmIJgc6tNta4SgV2hRdM0L03juYYYQNd/qO
uhblVbY1cxNFxokp8aQsXSL0ZUiY/OOC1qi5+VQOgITHg6DI1EMy2dB5gk/0WgHe
IcRrzWFDx9x3XfjW6lWUqWJWfULl3sm178Aw2ZrUdcvyTtQsp5fY0BWC0IWvapVj
GwfnxbkVtX/Lhcf8m2fjtgHvPgLEc7v82Q/rptdiX9bmcnMdz3TWtbGQX6q7dYpf
ezzGXR2OJixMp2FZKJe2angawCUaQjq75DO+RqA7RzTUd/QXSbEmjErds4iHBuoj
P9OAGtX/anETg0mUy9D/l7zzJBh5BaSb+ESb466MKcg24tDAoKwxVUh+A7nTzMor
Uui7S5XjOeN47afmU7R6BD2r42Hj7auUucLYQQR9AbqyHGyLcGJB4RFcDiJwmy+5
W53jCL958YgNfQ6IqWuaoPSlqIaKdcSt1mzyFs58czepkzxFfTUJPipEKhqCnrHH
uWKJjASDcY8oxjRL3NP+VGDYT4iqise5/EUHFuiuCuWNVSOapZYVZzc3/yK6xgUe
UywvBhUM8Y1NNJwL4JkAzgN1Wop+wjQYhXP/FHjZtBKGBUqF7dbBYLm2JfneIlgR
JRD/20C4mfS4agAjuIjYb+aVSNmnPR0MyLdtPnwLiCZSO7077x0sluJVneIcf7cj
/6Tk1iJ2L6Ljmtpd1yTg3MQH8KIv//lF5NnS7SDvnXbIE6F4XzhvKv5Ct1U+8WRG
FktxPRTKudQD/gV9XImf6suvOlxqj6ZHC41yE/n4Si0otAj/QzPYCbof+tAHCnj2
mNmptwV10XPpAgeDd+ODubSvuIx7+X1aXsU1vlYo/wbkFouzgwXraph1eeehs4hR
fglmYwpui5/x0L7f9p/u1fyBVJyNU1i4kCQpCN98uKti9IZ5N+XxXnNbcn+5ne37
e7uX9OustanmEkN/J4wu69wgvQV1atF/JGccfd9JAWE8hdkLotyHNzpKeKvF7kyV
KT5n/cySPc2SmM+L1EOm5EezgCgvGHhOTD7rpezwjCt691WyOjdLFl+qUyNcZuXz
ZB3RUL0XJgR7a+m1aR3lHEo57sc9pvglf7pdie4l4L96h2rSL7QLHlUXC4j2L8fA
YtwCg1wbyiw7mEb2M9eKK7jfpx2KR2jr9zdXuqqcGGnNcB0VmDb8YvbPNHK19FYL
7/RTeNZf9d9/REQxEw05uNrNvL6ls9emfdSQeEvi46GVvivESVRN3smlfzS42CiO
Yeggy312+amGqTeAgqqIiI2MXTgj+D8PHN+AVoQSmgOPNUfGr8xUHgEcm3scz8WV
AI0vB4TWmfzNA+WVdv4HfvdGv3zYRCSPNAc2hgFIIJHA7hfjwaqhtj7GcdgWQR4H
Et/YW14Q2tZgRyFm75BL/QOUgGHcr8IvXByrxVt8O/2OdiYiGppGGCiD9DFq7ws6
1IRfTaGvIsy5y/iwcp88WMZESVZuy6qQiCOweL8idPlSBFYKIFAmgWmGsQfdp93W
1S+FNBJQnAAEuu6gn1AwKjrVc/d93zlpkBlMVlyIwVIPsKnLiexU40NeOLEMOIn+
tvndEqSXyjijlbs6Ge8AZWeto1/C7pYN7TMH4Pdvur5lk+Y3C4vSV5nyudKkrW1e
7NiorwqFZBmALL8v+ddz/3J6x/Fd+v2r9Q7IUj1qg8pXaHA5bOxQsa/eqhAnNvVV
c0Nj14qpt1gWbzl+fySGiH+ckoaJ+r/ENM+lqHh8Aemj66bQLO9cz948CJms9SIJ
ZbAI8Dl7dDUY8K0THsqVLzx6B+2iKOgxg9rYDDFEvhV4wmCedQNShRuZQYCN56L/
PbIthS7PeuP1Q161SfPgh5mEXPoRbM1eq7THAKvOdY9EM82iMTxtkYxkbEoZ9ysp
Fb3+QrfybrXpzvWDWea3NVwkIK8RAUa7vh70bELZq0p0AZHkIFnXfcr4MRtAReMI
XPXvjr/PDaeg3LbXvbDhBvjougtWaMWqkeAnWMed8PxbcuOZaVCNCInCtUNKgsfS
GtvozSAgXyy06dpSGdOZWtXT37onw6BJ39ZnFzL9qKfBXhk50RSCovLGMtK6/sd+
o5aeSsLDpbqoBkUjGF5OhR014rWqsOoBCYX2KW5OKG/E7KYsu1h3oGNEwWjsmNy6
kvdnBA8NZMkM2Yt6VKkMcLbxnHcdmn6e3499CT5OEUfkz4nLcxz7TaaHV7Q0Sdh0
RGEl7m3JzfP71q4+l0rSsNXZ27/NDTMv2JWQ0DFaTEQDwuw8cRsK8ZPA0VEcBVbZ
iMfoF4z/d9WUxQs3z4OXWBRgFG2DAucrbaLNLoSR65Dv8EE1T81hJpeTM8U0T8wZ
IWfE4FvjTE+PwgHNPzTnGoq3k0BQmKZbK4RwrWqUioDIVC60P7PjMfQIQDBoazkC
wi3GU0DDgDVuNS7yX8t96a5UCEZrXi6QOzZyHDTY6oUyIxoX+uveAWRZs0Y/zuAZ
Q7lGzJLRponEQUlVxslHrg2ON1zYin7Wxs8br4Rhe+Re+/OBJ89QXSRtRGSsH2/q
zjoRtWuTsSabKQ7wcf1st81n/Urf2DD5cTAZwELLgE/xe4VHP5uPC9+nzpNYri46
PnhDqURt/1GQ7VsH8tVyDviUSJ0dlZNqM8jCdErHRvgDcbvOjOYYoB2Ehkz2fwi9
RtbwOFM6k3bIdGQbRPgtfuttcJSd7mcjuS8sIzRZaVKhdvleoEf6/E3djpph0f8n
WZ+eues/S4yff+XwlW0kC+DcsyFJQ9BsdKq644HXoTnCyNEkFElBv0DK4cG5jd+j
AGrubUIZh1JgagEI0iTn4i6cpHdRFm18ZdkAxfDHxWN1yLC/jwU9WzQ3jqHP90qg
rsrPsJOaNIzbbs3/xCjLD7XSGqh0sGEG0GucHqzIFalz67HD9+KE5iVoI0/2d/rL
L51hRlBGDVfGZFAxQxvGyiQDvC4IgEXhW9v93oW0jne8dUSjSGHtrWZRwCnM9B5+
VAgsiEvVAIPPFmmgG5C42ndS0eGxBStvpNK++pqIj6nSoYqLpAXAztcBsNpIE9HU
L7Xz7uyMx0rLBpO+YqTErTnEEOF3zQW+4tsJqty3tWMipFd6s74acJjXj2Kif8D+
I/A5ZWutIt+yFqu/nnJW1gl5JcVJmhCt+kBHbBSR3gjoFZ+cXQX8kESkCfrZ0SQ/
kN6zM9qL/IaIA9CQh6sbaJu8tFVjvEPEeci8DhJ26KYeJxxbLBz6MjQcFQlsqI72
+su5jldBPCyNkc9Bjxuk+oZaOw9RYg26Yl5AF96v06hjhb5vd/AuMsSE8SpC1NjR
mdA3nElYIHGmovr7FRhT56/ytftEVirvvqQIFMpfrv6iKA/fTBVvZU/6fel3n2Lc
nOncrVrGNn/3Y1fkaIdSgAkgxf2WZVI506IKBbdynYOdGxYLzRSFyv8M1yFGYIeA
OrukzoST0f+8sQycd814BFWIxd8+Zk6rfnIAwsFmJNC7+I2IqcjEICGwc7mfk4YB
HdwLLVr1waRV8FrkCCfbhJ8P3o03m9o545ZCI8zmRKFRAVREeeeb+QwKqXtTe8T1
jhsEFm4weBsghgdyp4fArYD83bkiymvtOv57uhsmeP9H4UUPLj4JejoknW/n59MF
sN/n/Ij4b2UA96vwViaNIB9tlyf9mI6flhL1hjd6RtUzxkQrHlYeLe6AF12t9HmG
FbMK1KYRjC8LEviAYGCopTAATjC4Oa+Lthn72UJAhEu3wDHwxyZ8TwjbXuuIQRCL
FbEhsqpnHNgL09mzgiOH6zfw6eO4RPdq7k3rCivtC7b8TtCpbnx4E/mmnlBXh4FV
+MRcaeYJHwa3B7Xx7PbOryQ8YU6cGJATU98xPsT9a0GyaTXpgcjRQ0F0amwohwJA
TZrdid0devQKgkWRp1SMh6XlDjCRz6yYBsHGOWy1Hu6GCYCQaYsRDpK8Ic+9wSF0
PDyvAAYaDwYaKQQiozWejwD98c9S1esA0SNi92o5SL4B4pKxvOBYTJ9BuBQX3gms
4WDkPTHjrAfxyKTL41GA33N/52cq8ko5PFw8M7k4RIsMaNmcnCB23TGlcbDHvf1g
QgObL7vVHXITmM1FNuL5lFPAb6vKc/XqoXPP6VNHFUxo8B65UA4P1WF54eD+1MzO
F8+3/wZuRHtCDOZ8kQIwz3G3QDHOLJ/15FQ57AAN1gUFz/PDK24YdszqVo6bdhKc
1IzAqq/wSB4K6gpOz4z74eoycuuTSiRLc9y+ZtvJUDAU5W5vm1Run82Lwww+C7dN
fWgbMDWE4BYAHjF5KmPBQ04Q+7l3L6aRoUkiumLouXNVpCG0r8kGS2xel5bqz5bS
3pi9GIvbmXIthTxIgfmWqIXTytNNvGBRtGMTOYZ/Vnr2TBoDdjyJySweR3lkCD+E
zm36n+0GeNIfBnn/mesgJGxgc4oR+r0NEpyf99nMdE2sIDBScYCEHlAdyDmgjL7s
pFFfVu/DqJ3Kv05bqCUkvv3LFx8TuXVmQT3xqVquMkUpPb6F+WHbWXW/s3sXGfgN
Q7EV1hh1KqWkiQHTbj/fb3WyUDlWDuqJ7Nu5ZMN249E9icBl5/WRk2VIPQcQxtet
CPESmW2HlvMSId1ePLigzMAgY3JpJswkLB+U0BD5UmvLg9r9n98+exDcVLSiUVE9
JaAolfSxnO2UelOdx6oD/O543JH1M+zeq6BfDkKX2laW80Eo9IkXNzpTieX3fj4y
NpXOfhGzpmIAuHih6usBwOHvf+TVoOMvU3wxWbTQEYLYKY/eGscfC+/AnNi1rqhv
/WREkKzT/Sa8XkA3mtAdWknZBOD40RVTcCQdOdWP2PSyB7VtlzOae7aIU73wtkd5
Oi6oS4T5CjgmhZL6bbFKq8GIPgiUBQPljvF30Q/7MOlwmKLNq29PnOQhSeixTpRv
ZztdbZ4qo9+MjIl+ggmjnXqeH3dZLECd4UAgFa3s+48dl5avgzmyTp2KIE9XQKgi
5d+UIJDjRoIw+kj3FRa45R4+QfSm7C8TXneAR98bER+frV3vNMYHju9sSaHkh4gR
Fi3qmFOOncaUf3ufGnGjGgK76UAoT/VG7q3jJZUuXF7IwPRlQyJLiIQEmObfGLIZ
gQejJXb7u1EJYHF6JXn+7uuGgDJF19rK3JcufIW8zI9DzQ5m0sMYmgDvCWyZzly+
bI04bn2HDTVhdLQOTnjN7WAL60qqIOcdfAyPOo4qqXaH8KwXQALwINK3f3LMqluY
6cvpb0vuUGo7zHvfjb1lePMpHK5h47Qsrs+P7PHmyJWgMmVirsekskJncZHQChR9
3KX0P3I+1H5MMm/YsRXMdJBPj03mXy6Gy8wSeLsBrGjVJdxNIhFeGqjz/zPOLYMN
Goa1w1rINohSvNyKFx0j61qW68IcI96wdjfOR2NKeHNkhe2OEdtG3TqVYWqf8YTU
vgIBX/z/BSHcaouqcBN651aH3fst0xaTzO20TRS6NNy2Lo5UFcwYEYhn6ZDe+Eev
7hrMijZ6Cmu/3PmokRafR9jDAczOPDFCb9dW/LX54rFH0X1QJRkovhEHvz3JkslS
i42XsGdmGahd1bJ4WBT4XNiotdtB0GaX5svcbXTegBTShj2B67rcG9nFTPgIVITg
kuW5ujZHo9yZalfIcnotMPOXgdrGnbvvkb63P57zrjuMSunf8g8qvK3yeLfJCySq
8Lwkx5AlGR1a57AVmBGjDrpkeVGwjrMXnQPc6G3lmQx5RszKXoUP+mS8Z02gkhX8
8jTlpgZXaprSha5k8ieZxFJxeNfYbMzhzY70Q1MGzNMr1JxlzEwxzDOagzifkzAI
VpaAncFKAfndniPlwO/f2gEdwdaQD2T4qahwLWBRl1Z87yebMmso5RFUon1JZkUG
Yet8OfNtvcqJ7BNiYomLTrgPmZSkf1/48Zfdx5DR+0foFeS1fhBUy+KHARNmiJGg
7jbxLronSFczSm2q7gyirK+xDVRoSgU11P3E6ViFx+wD9ySOl68jk40kbEr6p9xx
U4mLPwqtVdWxQcTzfBSoIHdTj41K0w2Mnkic/SXjJEhlpCeM6FgfxEAxOqvXachY
q7otGb5ejnicbHFEe/jAvYtsb3Sfk9Mbj16ZZm4UUdASmEpbc0hNolLLLBbcVZqg
KaloixNW0+M/+jxBHvdy4+UjcmaEGA+ZFZs226FgUujFc8VbfhhpqDSNi+P+u4yi
SIfQV+fARHVq7WjEzYLq7dtTnb9L5TKNBWLQGZ+X+z5mmtIsjWkvoOTI1rs61Bww
DM0znHOmftL8Ptwn0d6uAbIR6bxxsgtjgQ/hxaF6ii018+Vn57Y97dQKlAywVvNh
hbx+MKqbGolkB3iRUKSHiVbP7jP6KK7zdOpe9sHKDhO78gA6uWg1ptRZu2T5TxU+
0Ss0hhp4MVmctpga04049tEzAwkv/cUVNte+hHTlIeEwh4kYJP8cm2TcHzgB0XQu
54jz9A1PVMVEqkvEQXXIDPdecA0N22AET2sX5A0XSoGPpXsw3wSBrzcMudpmy5sV
6RSOmGkOw8Aobfh62eUoKAyb4CfspmTrI40/8QGr8qg/3A5NEKVbrN+NQn2lOUiz
CkRTsaVdP23ewMxAAKt9vgb2WBzPPmBQIOUQ/pyS4CA/aHkj6YPjZnn1GadDR85q
ho3A0Q9flgGlZh5gF3pnLTl6/Tkh+nwGU/RHuQ3m06n2gnx4u6kBhIdZ11Q8a0Rr
Nh/Xhf/+6z0RCy82pqXeWitjWp1B48AFcAi0qgXuE/5B0qMKDxTTNMGAAf9WNL52
MrXWwhR+TdGhMewInulii0pL3MGPQPwTLHKU96lo12wkapOXabYED2Upg3897sHE
NhHqK6o4Ct2Nf5dbmZbaeB+qv9oepq7I9S/YyWebt8rmOvIBWWgEniS+TPWGMtMn
tqH6ciQU7FdaPceA5r65fUSWLTR3D9+PSDxLKTbdQwzlLHtqd13R1PxnZr9656qC
7kS6pL9LBSmOS/h43DBX4TFXH6ymej/1AGPzDztMX+dZBbcSEn0kT/ed+aodxs1E
gPvPd1N8tRV132i1guF+1KooefxVFlQPWmWTXmtEZrj8bwU5oEj16so3hr4R+/n8
9pTaaIzv8BWyjIYrWxNNXmd3v5C7mFJbQM5dC6loxJPFNq+2z4alIbCY5MOrotZ9
OxXFuKG8TQYXi0T9YhmsUDRxQWyV7FdnZWjARhudCETwYQlKSGjahXQOT4XYtOGs
HynNH1FcP/aGsVTOP2b2GOAtXKuz110UgD4tyjJbU04Upi0pQEsooyIiC70qEZ6A
jKh/tDYRY2+kVL8AwsTsGP4kLm8Vc+JfWIsyN1XtFR+QJQtl2pOhyMQKXz+MO3cd
F5sZcFPjYVtMDFNpekYQ+ammLSyFEDcgKP5CYNSgiNcYoBZRZzg8LjXhp175Sz0v
DTXjuDQVdJk/HJ7UvNQDDi78ZfBdr3pPHVX/61nojLRs9dwiydRFHJ63DaOkRHcm
/DujdyETzJNIYOv70laUm17LIeFzqNm2Q64dC0RMZTmLhgzX79NykmMBwthcf63z
811ZrN8052rtfAxjE5IPoBInKC3l9pMTXw/nTExno1ScZ5wWhg2ykhMeveTTyEQp
4GQEh2MV3K1/4TYQZLYnwLwLAF0XdtkeOYims2TzJ2DOj6Kl8uknS5vPe8mt+rwM
AZ6cjyOM2GIRw5LU9QGdcY4O+R9rqxtZeuwijMb5w/X+ajqWDW03GdblysDKjZhB
q+kvyAEjihcjYrRU882w9bJaOUqfI+jy9ltSMXnm6pLTPkKPVg8SsByVDnXUhOQ1
y2/ogntsb4gR7xROncYGFYiS3wOyMNjRer1fBrjqGDoCABF1s67kLB7r+2MRzDQA
edOCAa3Ng0Z9qpLuKSiSpJ1SastN9ncG85WcgM5ELMPEa3CRGt9pReSmuaDSrICT
6Ip8whk/9j/u10EKPmbXJG/xJ/aadJuxVdzHy7BuVGraokcvWLppZFuxIOavBB/q
mA6OsnLPzMj81rKWFM/UGBP3GjVsYxRKtSTflGc6YLTqmOna0Wk996OY0tJEiLi4
jWxIOibazC8KVYmlQf0x/r9extGCdAKyzQVP6/FMaYbzK9SraBxVzrIGrUCTS1ur
MMp6DC6wcnCNY1hrslHKcZRjNV3a2Br75qcGm6/GrMqWPqI8iGUn84JFc5HAUTBZ
frM5yQqMNdaM9CsxbAUv2kc5bXKa++jCOriJ7LmfDgI4TAh5h2JPixEc7Twl752A
/K2ZwTSDhy8DEQPgOQviS9B22Pkv+hiXJ4KuWZGOvxdhDne4DZtepO/8ra9YoBHh
8AhvFJKQTTbq8zwvOaRPS1RRO0YRIaSZ+XKE/xqznaTcCSeqh3G3fvz8Zf6LAnBQ
DC6dccrC/GWvx7PkIn9LC2xLR2tMG8GFmG4sOK3jUGCXB1Ga2r/wjvRdPp/H4BbE
Zo/rETLaD9wHkGeNcigghshQTwd6NQ7DaCpIdij4EOXzk7aR83Ku8KeOR7ptwicE
on6nWOGVUIDRGbsgQliWoKFTv65hEsWHhP4UNugXg5u/s2R5ypFg0tq3bXvX3dXe
+59fQ05krv83E+ViYhBRHKyqpenaGLiuVvi3YGVA7v3Y72AZCZuqhcbxbtJAKLgt
sqXt2J2Bqhmf3TZIJhoqEqbax+qhhOyZt7voipNkfAZae0wQY2+ZJ6bFmQ5P+iy4
EMpPwa9GVweCS2Bt9XS9vNon+z4sWU6Ib9ODuHFpeB1joRoLYz1HyJycPR+ZW8Og
qFlvuNuZ8bukH+IVKW31S6Zyx5VQ1hmyPOMUYSVF6+IpBuSEHa9Y22J/yd894oFB
K0bI8nMeSEvq3FVcEAa3wA9gn8Gztg1YPZpFsuJ4Yx2KvObDak/cvkCRB17aFlcT
+mJe4JTbHzjnBJn92T5VXGKjDnJinT2z4imqsVuRL2PY+nDHCU2qI0meM/2l0WVj
OiuuMrXwEgdZsfSXQf9rZH9mU0izLyFQMhflQFwcYjSFJm5TXVQVattvEqDfuoiy
Ud5GxcmPS6PAhl8XxGGqeWJSpUXTKqRTyUegpMeV8DwS+ji98g+Krfda52afJIY2
QP3T6w3TsKHbjrZAf2YrqnYttnCaAqHmsq6hjYgYNcb4Z5/8YZ1HqphdUBB1ipbW
o7fXOpRnxd8ycwYG03uaIO3z/gy2/m6a0J5WEl9X/XBnvMcNUfXsuW/B0VDasBJy
rycaIyDAHXN6r1mH6hL4eI8eyPab2A09J0D9XstfjzJd5FeL8DzDGA/eY75TIBxV
KQyW2GCjf2oFGnuZabBtLuiAA3XVVtDavpTw7nb/HuTIPvyyRy0/loMVoS1u5Dwt
xcv9DuAkew6ylZlp1jbPX2vbtBhtjNQoB6I6KcQ23rGNb/1C7oiZnlufjUmxqkTv
CKvzT4KYi4C5FEwN2rr29/XxxtdcbNM1rhzaAHW+1DhWcU6nzE28JaS8FnOI5bex
W3/3NnCBMYtI3eAWhPszbOEQ3p8xsVHzCv5q/cYumWq4QtIvBZp1Lrs3uWCL2B14
H+SiTA70/qh+Kpl1hdiyZDzZADLJlDZ5XV2hk0P9fWj+8TUXZp2aMo3nqtVNdOs8
vvmubnf8V2cSv+nj/Uh1s5/r+pDolR6tS00Hbz92nC94sS9iC3uLf7qv07WPQoTV
eJU749VM5i4CR51r7JV8ksdQnopveFCEIUHQ+SF8y4w67qqeJGR6ePb9Ou3TRO51
tmEqCGPeVYabZBWsfh7MN7hPqPweXb1pirws8Q5jALR7eUykiKYnErtKyphOZZ8Z
kqHVXXhjJsom/DiDyVuv8IBeX+M+sZc8mmeM+oUreE9g9ueDC1EvWY034CO3CBtQ
5iYyzGtyyLazpdtFUjrbg05msx+pgrLQwiXvITxIcXUygwnfkzjXhwKg0hfipspF
R8cMP1z++ej2ZXQkACParFXHyi6LvfILEby3HbembmO9tirbWtpjvkXOPvjCiEnP
GXX07OPF9rvMGPJ9c7rjGyrboLLzsQ403JCgjsJl4k7zB2pEXWUuHR7wB+CKp/Ne
vcK3t9HnTQXzs3OeBB6dN6b+cCVDsJdk9xS9WxhpBR0MuDqtvyyapn/3678KcvIk
z5zP5GpfLUuObRaibyKyW1cSKGVk437xwElwCK6LeqDms1IRGOzbN7b7wAakIN5q
weT7zCF7c7gzAygdG+fHktjG8T/OB1VCrqci7kzRNBHYkim4tEOgzKNTaQuJVOqs
Zl07AJU3xme5qgZRc/Si8iw/NmJeXvzhqTFS8s9WkEM/csKYNN3hi8gG8YxHs5Jy
rwSOuD3xIuttS8zbhUhB1Llg0imyszyhzGg5p8wRa4qlavDbwdUisKogqrMbsbNi
S6Zc7o8TSv+KxwKPScK3Jtzi1FATQDDqnkXoQ3KLdHPKdtGwkuo3z+7oZW5NmM6D
86EHhHH7KQC2oz3ZdzhbFOrRF2VuOeO20Ks+BPVMqHEkpp/fX60wyf1HzYN83d9e
iDmnkeiHIzkkVaxX7ObGaA33+XbvRkWGPfYZuQPspbr1so2CWNvjR3Gln9tJUn3a
J6VVJ+9ZnsB63Qf07gqWoj00g8i0iGWjsPi5jakRN/buguPc8f61LNEbo4ZR+GlR
NiYcTfBTUrSr7bK9JTI921SS15hoFu8yQvq8SJvJXIw/DxPaPlZvP28PcebbMIhF
IPXuKFpFDyLFTGlWvYoKgZUL0p2nhLKTxFFDtKR2UdWelb5nCZndYqU7atDPdIJR
ay+VQuqkHg6SPaCguzAJhYz/mlHb7TjE8UpTxexzGr67gSrX/1vDn+5HfXcm4WpO
EHFgJgLHBxwqpQnA3SEYuWpo8NwVCIY2x87kOtFlMdshZiqvW7uU9O3A/lKYi+0I
ccuUIOjxznf3Eu6KzhjR3I1Bv443X0lozpZUoYxoGIBY1h9/Ni39CgXNNejyxaCp
BFMGHQ/mCdHNNrT5rBeclNk3ZnA2fA7hPQl5uLVRQk6gtKFW/I/CyD1EWgobwfjc
dCmTMjNIrty5wk60yFGJArlFCwQkLrIt/UvdK0DkZxTJ9bh8fydW2vuTRNs0vUN0
ftQBdyURBVXGCoHTWq33qxUNkgU/xIp9H8srEdMW1ULZB75b1kLf1/eKpnvNxG0t
1f2NX+Dm2vnrqmjsqWHZmc4qwyje/lppmXbSQ7HEHCZMrAN4g9KHz26mo1oEIlWF
quoha/7FZC0vXKj1rBqXHfu7tA0jH8qPmj760D6MYlX39k8ivkQWhou1/94755Fu
vmPke8rtuuSxCfHphgyeM496nGs8ZLaWb8437wA5sSITFHY6129RnC3H+lVj3u7Y
/ykmT7JGvYnfkjOqOHvuZiKthGfJywgELeM/5jn/rSRQ4CKB7qvK9SU+00Xg6vAJ
9+teTsimIY3yBl22+Sr1MaTJarzkdyRQXXGYvlT+byh6zxRdVvkHGPxVA0r7PzpP
4xneLJ8z/+QiORbGKV4iTp69P4C00/kKayAcB+Tn06QBoGIRM548tQmC61Vixg/7
gGDX6bRwtTSUvAxRrBfgZ5sj6Ecivd1gbkeGwI/To9yFQ1ot6UaC2Q6Zo/vFsZu/
marz65nDap1YWRYz+NtSu8qKbjNihwJugoIfO1ItvP3B4lZKu+58ZSrXlQS5eZyh
jCD8UrwKsmzBB5wBky9cfcqP52fHz3q/tTQDXeJl4M9fzwR6qieVvf7D9leIwH13
382XuBNAYw+q8aV0IBLW86CUxJ5MelQhjQsRzeKFVCWJzsidLuILGJTgruNKoFGA
6tAeuxBczqdV9rPUQAtjHQDLldvJZ6EX+NxUGniLfE++WBaRoCU0zWKL38DmxN7p
5ydZ4WSCcpn+/3wBB4Epos4LWRBbBrPLXc+7W8Rq+Nbj4ScnOTe0tz7Lc9qXVHWx
Rl+PJaL91qMA/W8egChlaLs+OyQSEE8Sd4zg8WsiB/MVekydvC0w4cmGZa8GZdSI
KrUx9y4gJYxGaBEjD1MuOgPRGpOREL36u6uv2Mwks23R20n/UW7Lc5D+0PhH7SbI
SHTAUlf0H+PEb3CEdIA9EDA2drXv9WyTqGK3dJs/mQ+s6EJBTbncLXb1ExbjaSHv
ccKRIkAqMGZpVD0E90R+N3ThbLjq8dQng3GVZcVw3iTFRvQ/apE1m50VCITQH/aB
IU7BSZhH2cY17YB6CuMuXpupbzR7B1XDVSYrliew3zAJwxZBKSrzGFFuK5M49AUu
939BoqWdbhxUt3to2m061vuaDsP7vvNMZ0y+YTbFVjfV1omCMWVBTKqUcDOwRKxT
dk+/05eYehS/pT6CL5osR9L4xEFmnjekoMTRNoQadvxhtKDhN/VU6gLYTqDGvx6J
XPZXMJe/WWqHOmqFyTXHzilIHu2BXxfkmfCPd/kYZv5AW7hQIK3EKOiB03ru9Dau
JQmtm7oKzGooqCcQWkOq0XrLAxPqDs0fxJXZKHRjz8gVZC81xUyfs+g5xzV6LqYK
F1ZBAV0MmcJR0m2bAYr21yjvR/QHRdeGginuGW4hmGGa8s4x8KklDKEwAyTszTUI
Cy8szAe0Rk6ZUWQHowRHekWDe4gwJ92Zro7NWaSZljkZ6cJ9tQ/Yin60SbNnx57N
1u6cTBQ2Mr6Thooaz1Mw7Seg23x+DICgSOsTj5tyR+U2+DLb1Qb4e28zRPQ24nR8
1VslX5mbwfK5KeCdAp5R4nZrbOFXc5z7Ami17l147H6YSHT959Rank/XWgEHlZUy
TmL0uMNr8ph+sGeq3oRihZPkCM6brnCBaBCUPtfXPerCvH+sVjiB+aWPNPSh+9Mp
4xojcWNvwbd8cy7x8lW2pOIxNLO/29G8EuhiNhlxPXLW30WU9VIYmCIaVmBzU0FD
iQOWD9wZ9+vyLVPMJAm5WdEUZutQlIzoFMHswo9897l7t56derveKlM8HtMrN0vT
MF00Yhxw+06QzBWbfVAwI4TkUcvBDZP7QsxynmilscoP9a2fKuG8YEQ1fl6oHUGY
2rwdyj/pcC0ZTE5noLkDjZ2FZNRDfbT6/Czii4t9crK4D/4qoqXJ0nU5XQc4tMbA
1XuLKL16fdVa1vN1Iy1ipRBH7PywPg8VLgY/jtu7Z7WhfOIokcMoPvwZgBZCHoSV
jrXvX8UOJZIWlL9dffkNLfG/TC7O/1u5SwrSgbfCK1MPWN3Ns7qjLsl3Q0iLvujN
ToocKChbvHNraBd0V/xqLDrGtCRKYJw+rN5GwfZYFIB1w3lMH4fhEJuk58epFr30
FeCHZhR0m1NoA2XhlSsscXvoqi3/0Iye/UgMwPyo6fqC5pzaEM4wo8K4jOpdydvD
d1T4vTDh/PuMCE+8XHEz5kASanDBSrseG26ZXbrYFbmwaU8uTuPYGs2ECS3zFxgq
TWYiih+ePniTzRpoXplJ6SipYrdcB2cNuD7bjdjz9FvBvdY5N7zRhzm6BdCSVfzY
Z9VmLaQS7FcbpysmUPfxC9ttgqnYsJReyxZyLRFrGd+g39zqMxs/+QBVfJzxOtSG
JcR//eW+oVgVCEGDq+BYW8ltIri8IXVU2fHzVIk6CmWS9RK7GBRGconuJ99bwgNL
ikylWrZc2YlYHNTI+X7bPcPUO8v88W/Cu9YNhQojADDMr/ynZhBC0q6RNiFOPucc
LlvwWnocbk7SdgIyBqHl7oHCEX7OGCzVLFSZGa0+ZytPoXThlccM46MS+UELP3n4
RdPxtDq1UGjAJEePxwC2HvZjSgVPpM9bqS7tzWMIWkRPbvFRjObyggcVqvkg/KwK
/v0q8gQogmQHKqg1JfsqosSSGiCBPEMRVLcpokG9U5pbzU6EJGoIleBVWhKeu47w
1XU7mBYW+kF0crBMr43mT3ncC/VcGqazCAnVzqdxZjZUix97wHFPle0R9AyEt6c6
9ZsdwnHeXP2yBNErhWMMYID8Zuzzq8N852q1ID98NfOCsVIufGChMy0nlr/q1DpH
nfy1q4YRWbmX6ZodTFdQFsmlB2UUGo9vOCb5G8qql2cEg/2zFJRuJFD7iDo0NyKY
T572Uy6EBbEe/pzOeTfMPExbXrs860OBnMCVSPWrHxyBg8lcoh59NACo3YhivfpV
toBwZhOop91jI/a/+5qW7YmSmSStCPErPJ8N+fSrXZju6qAQoCpmLhVe4ty/BWJe
CWpdrTG0noxTDs7RanBMnc9zjzef/dfjptHvQJfv4F3qT0tJo8NniJ8+RLOsTj8P
+XiyNY/BVgJfxVTkjg13YiefR4Bj2JAO1R3mDiNzQwFbY4h6RDG3BSM8J3wEBXVp
vkO6hZqQafbmGrOoWb/SYn943mBuoUzjOehSTdzEWlh0BWHfyGk/Iww5ZBFUaA05
LvFxSnz1H7jvez3JJ2EUV06qrkJyzuyj3v8qS9xAp1mcQd65ZXuJfmf4VeGqEdy2
EW3ReSrNg4jd2aYwfyqEB5g1cDcDuE46B/qHuAs9qAE102W2BjjASyqDIbSSYDLz
Pn3vdT/pxjQDJGFZ4Et7qRz1RZmCbNMlFVW+rMpZzOBKP1abiSpUveghP+EnCtHA
4lzT3xHusPUIGm1szHEIo36HCClun4tXRwCI177XpYpFrQrLebtxvOuULJVWnQX+
RSUS/cOLn77uTABnr/qeJfp5RQF46rzNeA0dDRz6OXQt3eULBkTgkQOAI3mb2UcE
Lsb2u0UDh/1hH24MQwCBylnyK2O4cAsl9c6hlrY6uxnPd4s31OujEgKHVxhVqZ5d
vz1pw2GXrT9cTw91PbPDZj2PGK0vG3Dd9nLzsX1aYgcc9W3wBPb3cLV6hSDdZhzO
/l+8nEbwmYtsZ3PLu8xnKKTgJ/Iro0eEXgqSl1N55K7laDgI5TuP4R8xPj+R5i1f
iSQdS+peM5DuqCxSQTlCOuD2QSTcFjLn8WHZiGPgAdsYGx1PojjFp41Qum50IyzM
zYfTBIEJBNseepeu3fm/Np82M88i36bQZ6Gqc6cRo8yfMv27Xa5TsYMIc+f2Rbbi
vMwmXLNAhqdgqxeBWrVnOtdHrHuZPPGXzNaIcjh5ry2LgiZYgCp+c9GI0L9iQUTV
DMdSgOUUEA2aUkupBLd5ggzR0BXU9evLW8xRzNE1mTuvP894BkkF4xjK2g24t4hr
N0f6Z3NxerDWoUov51Kz99HGv29mjcyf5rm7RO0PUNlbZvWC45gqmdi4gx0wiGpE
c4jTD0c5lplQpCRkjE1JgBYzOY5rEO9yXKE2TzmOip3nTGqvW8mzB1udtRjSJMWN
GgPjHLdn/IjryQAieYzS5G/CY0AmYV6LKFEaWinDse1coflyge/FIm3TXYCYAQyL
FCUFblzI+DalNWWEp50Gu8Q1Uk8oNhgpr5SMspM/rRs04QyqAUFCOfvQpX8Np+yl
Nub/oKDxrUov826s3XdUwvc3bF2CFQo0nLGvuE7Bl+36mm0vw0QB5xqlU5qUVMke
1xmOvpWoiqArbhprYRK1oOLrn1euxU0JnrNIFGTvqOEVKek+BI7LmEPuT4LVgtpd
V4JguSUYMuy0UZRgnaPq26WIVFShso4e6VGujSWh6zvwfGJlUoc9iS6yh5Fv4sEm
CXWnnR5dsXExKJ3q3IVj/ALrauADM0UyP+HT2rDpry5WUXjwXNe4xFlukVy4TSjg
ZJEN1DAvtz2A+KKcbUODUvMoql+/CZpZlwrC0GS6QlLi0/a5iaI1COt+XsB2HZXx
FbzRTn1XdH/h0x8iOWIaCnnlwyECbsB7x0NUg6rTOmM/XWAjfJe8CblqGE374aWn
TCXxe65RR7J9VEFVBTYtIqHKqiT7tjGIvAETugtpVcbzRwH5YTlP3OFcuRhE7a6A
/udL66wcjVSWR4T4TA/Rt/A+a+MTbtHJrHxGIHcjuoRaBBiwyFRmaVmeWotj86B3
5zX1to2peqx7wRVj4BoaX2VkgNag83SWFvyg3Y2UyXoSOhpwCY0kFfvASMBxWDkD
ut1gmK6CNmIp8TuWIV5BJ/wwSDZQP7M7uWeEF5CBGYLbsaZeb74MAafqIPyO6MnX
FzRpIgdqit+4OLdDfOMUbOkx+OGDB4Uwu4VzyQxhFdb8m2JVxtVC1+USZx3yx7IN
ceh3u3QT2dTP1XVmTaL/qZzZhyZTQRohrklB+PF5qC6Npco1V64cdmpLXGjGmXDs
FtI5i+CimZ5doOEAs7GoEp/27r7VUWqYQxXIMxkv/4vRFjSqGBId13ypJbrFVY0m
ueO5wwGUDRViMed6n4QbTaKYDRO6aaux2peQbVFKYvwYHEMRCiUh9Jwdrqe63TDA
gqX/rvksPJmjtTFSB36uaqdijtVjcpVt1cJDdnHoNAVQewsZIHEPWGJiYmj3oA4A
cpzOOJxKyoRAcWAKs6US1UatBwuphb4MfjH79C8y1wSGYXyyWPmmQiVY1Xvng6n4
tt2CPKZ3HO+FHfzhrm2DTX61nVgFfU/H5ycfy4XGCp5BViy7ogOXeFADiC3iiqkc
cVO+M2r2T4QFUJ/sguSSoNiiXJX3EU9DvomQneBIUYz4IUPWtkW2+WytHi2XBXCB
GL1pt3cHwlYEe5dA/gvLUIIBQOQaNAGxEuGwl2eBMKUDGS6Fv9C6NwXOnmvEh85N
RBM6rXWi+u8vPbcIUqRugQLY2ELm+lNua4IVV3s49WC7TVe02ifhy4h0tQILShYD
mENhtRzzdv+4ZhbiwyV1b0r/AG9SJcQRlOPX2lLUhh48A9KAElFxMAc+jwHnZCGF
N2OXOZERwMbR3CIoSnut2qyl1LncqNQlIARAfHVc9o/Oy/iLrOxHX6JdhAKfH8xt
F7RETDztiojEe+nYjDPOtSl0oq3t4evaF4ApCRL0k5dB43kT5VBwP2uCxu9ME5CB
0iKP8feCfBQyhg6xYQasZlKxRDQfymggH6bBO676w4durGlghaVfImGtjs5bGhVk
FkQiOaNlYM9p+CNNFhB/enVIXaZOuuHaxgARbt5MCidrCNLYudLTi9VxrzxR9Qqj
vJfDO5DMOrz2qpXjdM/X10e7Zya4oFHBNni6VVF4prs6NsEr0dkD+LnARWXx7QWW
j8ghGHQ/1OW+IsWhVulCJdGXxj34DSorO+RQasvSc4YpQZiYqaC1SQNJtv1SrW8Y
XJCZmfIWxWfDUOgEgrDZ/XCcjg40t+RYt/5M3IPxDF9JnHvJZcYX7RJ6bE9MBpC7
InURDCUnijfF2BpxT4FIdGVjNkeQiAfbcqmlC2tQSbVcInUYjN8ej/9URBz6gEgG
EHw4zPyJD7WwWRvEHmOP/KcVkwZBgp561+RKX7ZTFEbzxIvI2vtMj92KU8qLbezV
qmYJuXbqTtxQd7mcDLnT1ZZ6XE+xUfxPf7k8PKzkoxdcxWfsCbQrhz7ldwR9nf05
Kms2Oz0pJDYvUeENdj7B49jtCXNNSwbzbwztfl1v5Usia+GAQcs9V9NewZd27wQS
FjfoS51sZ9NaN5ZgHxXdG+B/uKzLDT2Lfh5wI0JgYTB5RaEWnO0dkZF5tBInHYmN
1TSghq9TE1ptC1UI9ld8q+npUVWZr1QNJYbI2AytfKOKwvOMWPwD+i7P/JdN/6NL
RQ4LA1iU668uotBkIN6OpEovhPPsi5AMqk46/4a1nac/SleOavuxa/HB3nWdfl7P
68hqRU367yEutK++xMKDFVZpGEjTl247WCv/moZz39yuZJUWdMpIKL1DHARdp5up
mhgk9CTWGGyZLKfC/wUPFxVX/Tf21VksrD+yF6tG409mqCiUmNiMvne8xYHsLNLe
Q4KU+dItvwq88EVuBSCut1Kh0CrKBXidl4b02cCl5L4wS6mUWuBiC7dqP3WbYSvh
yBpZVAgsc7A3WM+Um2RkJcR9S3e2i7te+nRhDTh8m6FrujB/CftZd5Hml39MJrRe
YZnUicyK3rehtpy/C9AmUrryfPX3E1O/MYEfr5J3sl1Ig5sOwCeF3M83jv5PhHL0
PpCjqcIfmSOXcj3NW7HjykDuFUWiQGmXJopPN5WHZbkoeZz5WdQWEd7Ndmx/WvyT
pv/dq4GVS7odRkWUprEHMDtXSN77yOVsItJ11/iY6bG3T6uCBH4QG9R35h9o5TFy
JKeVlzXJAeUDw84WEflGqpCtIx5tJdzvHgIAERlGd+zS8/PtXkQ0sywjVnzPKgtj
ordBuUJMQGf4tBQKJ2GZhri1avs5mHTL36Dk0XD0SH/vlctf4TTEy81JgMv1h7Gh
qfo/tMKAEV7RCq/b+iWLFm0mxMgEkDx3R+SbysMbB9+wYgq2brI7nNBHXGPuZpKj
olCLm1xEiHmV1Rm1B9s3KHBcokLNCYpUzyzPcx5kFoNyD8StQc71J+i3k1OSeeVZ
9+7BVuKmD9Qb4BsukaIEjXvQveBQeaVyCDefkw0ZDuZYFLV3R92+5Oq+48T07j4f
AS/zySW1cyY5rLZws2JySV0mEGmfL2h5I5xICaNjiidhTcDK5rcr50E2KhQw3p2l
cjXmeejJNtqaLocyzt8uEesUQNU6VDjgY/QK09IV6+XAd/TkneBnaBtdwcM0qnVo
F2zcngLjOufD/c4GgS8NAamKnz+O9Lu5MneQkIZ7rBRyQ6yx8OX7y2UQ+s5Nv2cM
PQDfqzF5YY8MTOYv9vKC2/hReQ+gJrTQtUFb1ZcfsVvgu9TSP84Z2Pu0K0U5NRNg
9U981lEeKVvvvmTlSr2EYsKGPAys7XD11iBprfODusRE+LUczS8+G7VPZzGJxEhE
e/yhBP8RZdpai650ZChbEOPKE51Xo/E2UEHxwhM8IegxC0zAlmYARWZ2+//2KrhX
jmVKZdIPqsYweMt8dNtY8aC/pwkO1wR+3kDTpZlIauWyTiDUAkaxh/lW2LtLuJaX
EQP+jx/nmDA6uK365D2JUrEtma4Hemeg8yuVzn65lmGFHvd0d0R72Hu5WCz4qAy2
gg1N0c8BGctXJAVubFoltg7MU0//yFBWFGevAowMwzQuNzkXBU+r4zT7r/JLiFYZ
tRze7sPfyamEQPR2jL87/znlw7S4hYXRgdB7xehqW0qA91LlkeLkpMeE13w/qtod
Hxqhpg0T2Z0DiWQXbNKtBulAtr/y9QxfThXHEKVaHuOci0JjgC0rEKtT5agXHVVA
W0oV/9H4PEqZy3ka/L7m80o0N9DB8gmISzUS8fBeoTeTgV8ei0ApsxHGl99/ekSr
LLquJBVo7D/mPOQFUlqqWz6oy/Ttc9qU6mQtPMy1Er84DMatZ9fLu2BXiNN9/fEP
b93pgZO1yvi9h6xvjOJ296vLcBOQLKBW6/6Fr00nAci1FovYE4RcS9PPtj+HM3D2
qB4NonlFvBdVPM+sVeeviBlfHIAy/6tmkq5D1V+PVGJ92aFiqexlSZom6ngzANyl
evsuC3lmZmF1DRd4URxDfcsYEWtbl0Zli+33X8NUY0aqvp/yki17jbFDaxy/IiEM
sRmMw/z/QP/RitdWYPuyuAiVKrr9QzOkpIEtNFokVlBnpAFLYTVbXgw7Hq3qRkW0
PaxwbPoP9gTmIXOXlb0CBmULcUWcsN78kRPJinmrD3wYpzp6KWDPeoFPYznqQSHg
PqQDGKqbZr0/1dVugCBcnAUP4B2Q4QJ2s3Hl6wrwZvdXrZ9+qLkQG37RLoSWHMQq
qmbL6DifOovUKbXjpx5iIKBVPdklv6xp6U5ucGOe9JqHVA8abdCUgy7FjTy8/D7O
7EmxN6YJubBuLMmZwXuzfyziRoSsjX+h0CSRaCma7egbDWAhL6QwwMM7p6roEe7l
szkAM8TQce3243zip3D13CRFBaBf1yfry92MvLOqD0+NbeJ9vTBM8WfcIP47xVrF
Q46lYCB+y74SreSxgTCjU6B+OkHVLh9Hn4kFuBcfowPVuDK0tzEeTALxRlSCl4zw
WKb9oDQa0vObOn9BRR3D+WKt55T7f3H1JsFDg+3ea6qKdJCDMi+2/Bmp9suTA8yU
0MXWBEr6ESeISNN7ZM+Ao8N37ixqp+wTJpcM5Mulhh91djaj4yp0m4PQHq/D7C2g
/95WQqhcQwBejzuXq3HK1NWLZMeMJJ4oPKNYTJ5H851arjZldqknWHPEFFLFYT11
t2jqMVOGozTI77VyXsOjqeqNLeyJXeOqaGXpHFHJinYPBZNV1RtOuVNN5nQ+bfGM
0Ska58uJy1mevO0MYZ5sm5CP5ELkqpXraZZri6xHKLLd+y04ZXCBKocMJz1cGj6d
9TJDp5s0i5b27ikSBMa3cnb7qjtokgD0P18zMuQzWsu0UYSiiw02z+i/Fa9hT5/b
/exOF0W0CyAbqJKe26SKkA0dnk6uhFO9KKwVC0gDu5qthhGlw11NnEzD2PQWYQEY
1wSBaya7HKIZ5DJPDczM/wsoTJKAqG2RJ8E6spwAw6uVHZOMeLAZRiuGDUCrKenL
c2zjk1Ta9GZtJyVMatWfIbFCX0KBpszZFpwsvIPNc1I26ovImh2rrNWlgTyxQ9Pw
Iul8SadbMqXYoD+8Lx14mP9N5R/PbL4WPPrlph/F60ONl6/b0zli/jE5by2KygfR
oeOG5JlouCeFhZOrbT7hKemlxSUBznbkCtmRgXsll11Qs0YLeI/tbqJUuc5ONXdJ
pAMp4OgOYlh8AA6vfNO8i9etGy45QJkhEggzM0OmSy8CKAwZZDo9onkUr5iQpRfm
olGdHKsTNestPkfBXtV55i+YIYoCslHvvfRWEoJsXvyS0r6IPtRkQukMdODeLOqQ
fxgvmobonWOYayCL9cUPNGNaifrwMDUHGVgxd8rUsB1T8ApM/Kq805kKooHDhcZp
KQeOzi4LYm5GgoJLfX+ipfz6tnkTpIDlKprXA1q3Mj4DAbn7s9DQKiN+wd5FkLpX
rx9nPSKKJZDm2ZxEdLNcAPoe2+XfEp4+8AGgsNbgDfUAhkv20k8u+zQI5h0KfPZa
C0Z9lO/09kIsyF8zhHpLMSiJmmi+lkDlFvo4s1v9ix1vM5qrptBX7Cz5y5zsAg1t
RSdYqFxN+Evv8gTD2lU83Z2hmWyRmQF4p+CIqTlNJ7vbGVJyzE4dxKuPk63TFr2v
qgWchHYPzPP0MSJmCbOpR5w9ItFIOuA6CueXZt96JFQ8gneGH/AO0EXT1fTVyKl4
93GbuOddb+gRsDinjWu7rrN6mDRRosH5N1lXyXCYtaPx7LQUbVp8fX+Qk3v+Fz9i
pb9YTSdpUIDIfnfhvYc2gqvE4NID+NYONrA6uxObW3inRIF0zkagXMkS4V2miRMH
Hmm3F8zxwTWnHEqah9wH6/civmOTcJupO4WjyTOKYiJ24LICNR6vhp5ELKVjxjg+
bFGKe0X0+vJhgUp7RDSjkMXJ3XliSjugoDhHSOrLxw+li2wAuTXvdSVJqY4vyvp8
pumr40hAJjtpAJ3mjqAs3yrmBZUriQbS3j9LJegRkFK3gGjJh42dXQbM9gH4ci8h
HeGG8engmINZe16t2enzFiivDMP+haUZlZHpiNMi+48ylSBdUJ7yFKmXojW6R69p
fnmdbXpMjoLSqCHLYYLQr5qqFovXIPAUoC3eRL120VnM4ynYNmjIH8kj60CLL5TK
2ARraNFRFTJL/Wwu2d8Oqk1+XTsfkd8sjLNHasa/FQ9gUip2ex9V+3bKxlm4W0ni
FpJyvSu0bNm2evcXgDnpnoSzVd4OJN2jLxjgxfIVu9LP6bppg4IjAAjuW2946I70
/eEapIH1HAwMwhq9A3XDeJQaKYSQlEBPLFMlrKtQ/u7eHGUz3mJ/eHpBj+PJCDkI
JJ2dwkSt/VvQcGB+Uo0wgrniuUZVLW4sRyn4JmI8qwoQJzsLCWwGk7u5eMggH12E
jLYPAUAnGdcHF+4UFRYtl+ItKisorqYFFplxWKxrcS1Xxa5sJIp9w4v5bQPqkP9U
hL1zTzjYzRC1noX7Ukk8f5HKx2Bi0drfkfDc2z1ycbC/ZmEzYEsxjhAT8i1ipKAi
TKVv12nq3Hg2FUlyT/GUxSyk/RlWQqrfLigMXy6L5+LxV93AexlGPOcCKj+uAIJp
2hsgSsy9qEE3Q3gUx0962JJFgitBEC6LM7ZmvuNPfSSkDCkkgt4j5x/AKSP9+vXP
Y+jRGFnzNglPttUvwXfS2UkW2CreWbP0YNnTFGIs26CeJbMwhRr2e5HaUmlaLiDT
FTxrUEelWGm86YbLR+efjU2WsYgqje3e0sPpm2qU+IyRkRokIvvO4hAjRhyrxj1b
pFDDYaXN7H1SVxzPbTVW+19zpLl19PPtXWiDUOhtFUiWIpve33vWDhOt7QVp2kUA
pgEdOsN+E24MFJqr3KQu4paqM35C6/urb2dHt8bVo32JRhPU1tcvdVm+pkAL4rDo
Rrm9SWtAiDLDQ2Z5CcrQ1fQs5AmGta7Pl6xyw9R58LxO0ypJiZ3QAECANN552cyH
NE8BMBCQCyj7V02kfeHrLSGcH0aycdF+44b31smu34i2lyS0SIWuUo4EU/7ZArOX
w8bTTgOzUH8rDddZXTBszwtcjjZfaID/BXT4N198NxsWMPuv7nZ4USgGQAxDUTJ2
9pzFLGWdGUrWZCQQjTgKUByvKCxujo/XkMjcZH7iyFIP5wbtZ5x0q+CurDjm7K2P
izr44dsxWwz2CCUfrsc9xmspB9Pr5Wg3QjA0PPCSoQvQKCwGDdRL5AoX05k7znzB
ITEDXjtTbNqCA+jQf+mj1i+ICWSaLuFAo18Gs3A79Y0cbcT0uRdvGD5fc+wQnY8M
43XgggOqlFoxYqV+JvcXUV9abtF4UAyhBahjrTYPDxVfPW6anP1dF9x6pVA0Y42E
h+c+wbjRXw8Ff+T1S5FButiIBohE8aQfryFou3C+HX3CVIZMy72LdDXxxrK/PqI/
AMkPNXC2gHOuhVqVMq2pkryNITL38nB36DKASjQ7nd92DCSGLusYW/3JpuxROgrM
4PVeJuw7/EQxutZyuL+jrxIrcUj+5MT+UnTXSppqC1mkwhG2d/gzG2Nhu33/KMMR
L7CchmmnQHhqzrXXoacdmybVGxelqLyHkbJBgf78HAX+tubNnPt1SFWXhg0wVqz3
HVnMoWooKwyk6BaCVubXiREBff9iuqtT0TsJklAQu0xXgVivTFgFzMAKe+A6ejNX
6QIaWnL29CBKRfsojwE+iuYoIYVHdi9/T0mlc16Wo0/KSue959KuSKrRlMBJN4NL
btweA5NTLsFNLUDXoC2r1cwzPo5iODfbK1PVeh+7+PJffe0XbLVC9zLjEnh05I05
pgmhVZC1rBg36uuPzdOxs8k2lfZBUHvg39vjBFxEwzBpghuR++pLcrYWzRBSjq1w
d29ds+HCTRbDxqispt14guhdwR69SdT3nTdNKqdNPAgHYS44BH8pKhfK5mgC1ohR
8ayMVex10wNqiz+wCMhxNsk5mI5kikXjtLYv4QYomEFbuwnyL+1K5fFhXd+hmDi0
/y5tsuGdUHqqJBtkNndfJQX6kFZcpRAUC0jIDw+VsOIpNvYKI+1PO4tdc1AsPnin
CtC5UjZtxohg6KScYFP6v9gTNlsLV5DKTVn7e1dNiL7Yog/tvhJzDcsxwUHRnMsU
X5OKRsV7FU4OrCOGdP+gb1HnSgVZ4HTy5HfHvA4xx/zR/143r0F6knPt8gSUL+2m
H4ITsHOj9nWqj6yJywBYz0KuFi9N2Q7GVwpwq/fjyq6ocycZgIbl116nJrHdxm/e
uSlxo7dld+iA5cA4q1DWZxQO+5NkAdiBicSMKT3vrHfZu7sxmypBsKRoRsvcylw0
tf7djNoPGrojr2iwFBrQp7OXdyAPx96Gv77cVB+st7zL+nJsWD1syiax9jiqEvaQ
FLVeVm0J0qPgdd5i4X59uc87L0YSoxdOGdsrgh/ukR2AVwbQYcMYZKWhWZmL++Uo
RhXb08/1fxGQbxoMksh5RjJolTtSwhKPtT2rAbJ4RMslCkka1yuqjoaqbvPeql6L
8phvMPzikWsYEYJpXP+vrPNT1F1ainf+2S4/I7Vz5F0nZHBQgvPaEsTEMzSj6+fE
r01Sdz5Livf1I/RZzL8a+7IIF8W2gs/mwP7nsETXELYqrWzxa2TRsX9qN8ZqK6p7
K5TuAoiHgEf8BaKRv2pEQYv3dUnZhSQE3O/pLQhmjQ6QFjnl1l3cmVALnJJs/s99
odI3PGbs25kkiciByzhVIFXkDJucEoQ/Ez7RBx97EHBYVdUT/4GfWeEy/h0cnE1q
lzKiBjaAyleaUd/4iTGrflWigKx1+5QWJlhWk3kMgvsixh+OiM1fVq8bcU6K4Mfi
aL1+MW7qrnOnZOIdfZYDGqG9EKRGA5EDB7hTib6UcC1uUPNXoSKWyaR9yu1uZ0Ks
g1wikxnZemGmwKg4O3w1qvI9c+g0PwRorno2KLd13ayd3A//ldgCkvcfI2Kb8qnz
Uz1kyLBaIPxIaa3/2+jYEQRuGkNoKOl0OKFWMHCrkZHtxIpBE/JppTkI6oO3v3dG
20rkPpUW73h5PD6Upmv8QnL+73MmeJbUtDPUzBVdfaG+EVyocOREZsSnJn7Ql2Wg
HZeZSdBpImjfnDDHnJeIU1zt0Y9UxdAXcMogaD4hXw9ZfNvNNE/9FU+vyJ4qgK8M
DI4FQdMjZT82tFOWAszv6fP2pV//Znjg6+COQ4bLWKqKoDknryr8wCFjJMzWfbDz
IrlLaeIcRZs8l3tYXn2i4jzymzupZGun8KvDXEXu4SvufqOUbZ8pbR7iX6tKAVaw
lkOkYHr3VIUik+uah6zftvxBYXVIc3yzOmtvetn/CnlkHLBQWxto2NUpJB6sHO7R
YKUr/IXKh5i3adCx2PKTsj45Evw7Q5r888I42CisRZG42jy5JFSXMZzCWT/7CYkT
FsERsWv0QisgAdayGWmVziE6g+Ly1kZNSNhDcZTwbvwRFD8GYIbiXcXCmawEmxI8
yHxwVErxTKH59UoUVjkD501PtMeiRDrkUaI/1SeC3mPXqB2NBV88OjXeQc/t9BYJ
k3BmXD4GhqPSC4cvIawIOitLi5/rj+lvsUPhNQgjjUyHK/FqgE4wwHpp4ZpyOnV6
DNf1cZas2vgLMvK+pn9SuuPr9t9+UM09V2jSnJYVZZU3MhYLgC1dIUBTp5+2TtRX
dP7SSuF0pR+wkFYLy3xq6LD1BDIlRQUmJzh7YAGSNQGhmPLCWikQxHW0MKGVXymD
f49EYmI4XMZlNf7Hw/hdFVeDt2fJ8OfKgdfx4m3Yrf4EU2e9exfkvEw4HQoI2d2c
+SwhkiWnWVgZujuSVGNuARcdYARvkL5EHryJ8DUJIEj9KBTkNOBanbWybWI3OqVe
nKeDeUXaBcL0WGgqsXiXR3hzBMll4ZtRT85/1Bk8E2F7ltQFIxCjmT6YynNVWi22
f0S+PnfXIXgISf4p/QPiiKVQejYiAygrykvqdV2IsRZxsH2XymRNZ5satkUkV4N/
U7r1ACRE4/usyT7ruYPmSSRTfbWkjMjiSicLw6LnuwdB0JUlEhnOJyqyvS9tKpir
KtGGVXwRzdnZW4cpETUsPynTx+wZBhcIguEDgAUx9ohNRdAA7QKXNmX+qNT7DFf1
XUnYp6hoTOJF+qRtR68WaE/TDWDPZpPnFF6QfCZuFcz28RRwQUFDHzZkXfiO/CI+
FHmpsLnNIj1mYZDRQkh7skJ8yN23Iz3mK7dbvHpfrP6OyCuu9qD7MBe1n7xwGqNK
JYcXDfNaoA7RMk2/eMFnujKTY4DJNns391ttGp0Agrgsv8+9l+b8ntosI891MYGJ
C7NrrzRBpccxmQq6lW2n63jVf3nEOADCx4wLI8+D0+bRqduW2ciGTIrmNv8dDUZt
B/lE2hp1H7sVXIb0LUbCbYMhuhALnma1WLNlvBDIVK/D4O9ORqL4ApuQwFeBF41j
TeLJRlrdpsYTDzybhOcqWBB5z+l6ZFxxWlyBaHzTIs/b2TmOCQAm5FWLcqj8DHcl
BDkJWNc0OCa9+BjeMtS/oG5GmiZpKSDXSv2mPUgVs2+Z68+PThXwhII99GP++Z/M
5bDV7cAws/tapK0ItWMn6ga7X4oyl3ccPhSyayQMGZs+50ZzvB/0wqALTkw5GFDY
VR1hVQMxk2JZk/S4fhE4I+Im9mUgOmTSIo4rwWSzgauwZgKG0V1+XtceNVSIgZa9
kteEAV0/B8RDb34JGYkh5VQAs/+EoJfDcDmGD4QMY6U6EqE+nbflktARymsLkGHZ
tpV8LOHXaeQRot+498p6lK0PzPKZvWT9EYpvZwv2obA8UvjDfWpTvuKInFk1S1Fp
4PjFvBGh3fVTduJo3DYWVD4Lvn5rPqQV9JyfISBzW+5qky76F9+hDtY5aG4u286h
swVQO5iCKWwAJ54OP4l2e42P83lHVaaleC0juE5s/9xRlDR8CREQObSh8Q1IACRr
JWkFR3HJFKfREebhWXvsvU+USwN1nI0gNeU30SM0EQC+I4FbZvsP4ArvTUKnVAvJ
2U3PjYUaaSIldpC3QsdfJgXnnWD3LJG/sI4BfJiyHXk+95uN04m+7jLiuyTCUzGj
XWkiRKfUjokJUkQWUKnE1E3E9mXYkyeAsV+sEzreV2+X5nv4ePEZ3iI7bFC1Pkip
Og1RX6xdmRl9SAFDannwocZ8guq3fKylinX8xImqSQhUJJpKr9TXGnTgLZPtW6yh
Taz2nM9Q1DmCMpYwXg/BYBknz2gAs1jbNluwYsFYTwpMfPQ5hdsvBnO1iqlLkrsX
aaBiDlojsVG7pAPayduukdTjs0FfaOIAtaixOCyvycPGKfGyMHM58vdQbDX1uCxD
o194wib9ziIbXh9QFchjUXzQu377+70oKEMVRLjxcPgZrtM6t2woTTzvULHNyarZ
gpQud5rvuPrl4dt4Tqc2r6/DWHGjRlaCE+SGqKM59yWNmIG3SDsPVOO4Ix+AUujq
Z50komHfaKNfEFDOrX++ykYKcFlMDGEmu5VCOMSbZdTEb6g6FekUf97tdsB+K1hk
htfQ58eEU7YNUr58rcq+i2+sZ5ywwAjANjsH4TSrK4N9rBK2wWcWJLXS6BZUt2wO
3l0/PKOrUChX3esukFHBqDIZHha5syA232U5I9MEUGBG4kms0x6oeLSVC4U6iEpO
CbUXFI2azym73PjbbpVoPCI97OQI1u6CTvz2U1cmucUdHL+Z2ijvQXg9u5p+LxA3
XZ/35ZHXFmYeQUT9p9gSu/1TUhH1radZsk6eGPrgr5DGItL6pApbUYwootznc4Ys
GaQm4DBGBfFEwGvDOO+GoFHDo6YdHXn3ZjCOH0L5QdOW9TTxepmwVbEJX5mUxdlS
eQWCG5+q1OQkDiHo2IKahGBp2+DnukYQLYK8UnDoTZioc0gmldFqzNGRkzdI1E3h
I+JbwHg7mRERYLIGsG6tN3srR6goeqOjW3kjA9Yvo4frE3oOIhmEEP8Vj10V7obV
sPRKO7r9fiMZYwGlP2Nq/Hv1OSv74ZrA4IMHms+oGfeyOAe2EEICLgoYajBQ6XQB
HvhooWajSODoWBSv/IImJJxcJxBdGAwKowCCMwfVFR1U/oWxlHe1C1XmBGeIuhss
CDUOxAuo/PJuG2ez5yXoagWmInnc+J1FYSriPCNh264EubiRXVRkewmeTIf2smWg
IU58X8aYPK9LOXxZncJgu6IeSdO9w8khaWHqICMeBtFVx8tlEFGL6OVhFhVycMPv
zH3irnj+5t8a+MXimsl5b8JaNlQK41QEzq2EMGop8l7scbm3k0/w6WmOlIpvDiTA
b54wH0MfnWBJQxvhqPCpy7ImPojs9cDJERYcZlozgPEFGV3h9N3mTAiHKY99xaDW
OVg26MANEbweGEH3+zzAp6ARNOXbpYNT1UvjYq8pR+qljFnAVfvtDZ2MFkj2VuRb
HeWm3Rd7zvKw9etnt06+fM6CaiuHEbuycCL9r+H3ROv3CFb6eEYcl7IhwBopdRwd
wX+X4jASexHJWHyuY1TveTLSee4wvZhe5KbK9XN3fNPCudVaseM0TrFkXYBeuI9m
OKZTX+IDSysCUdEmUEUcFv7ImG79ITbPp1oKTr8jmbbdtmd8vxwxgaq+uqxPU69d
1EQe+J/5h0K8L7UkMvOyuI1DCjwBuX/BgaZs8DpQISy41nbR6d9Ttc0WaWMZ1R9q
hyp+fH8tGY8TFSudyJhZUgVJhb84X97vIGHqWjjPEqMQGOMNG44M0rJDpBvEUdQU
3KnvV000hLKtZo/AxZrhaGfuYZApHbcCaKR5b7gry65Gy+EQBVayQTqL1zGwkOyr
B3H5rRVqohzt3JwX2hJzB9e2a93562oedtkuU+oqTiM+p32WYfhcosqK5Dn3M0Il
g01LTyUtNWHPVyOXoBmL1iErMJ2ioNrPVr+ov692YG+ZcbXqmQaw5SDZcSSvy/gT
UEIkF6cCWTAfXXM/3ZK+HCymW5ER0EswUvcxGKFokCoJNuz7SEixnq4K8G4q9PgQ
h51VbxYmvcvG1ypfnAocdxMGsZ9DSHbMHQ/s8wsDf/xULrkGjBM9wihNb46pVI+a
fFbnkySkYsTyapEzEEFhSk/vBgjR2NKQ47wwpOtr9qUOiSlJIwxUpycs/AkYewFv
DbzI72uwdKd4JhSbSkKWQ/495J57s3vTFk4VsYkkENnOECtXEzyxhCnANqyIQ70x
D7dPKnsngDEbZBjliGNKjcy2/PJYdaPlymYiizwgSVNicrlH/iKWABrQFUxGKiCn
RUVr2AYZDTTHw+JZ67auezb0DgsWXUcY0AvujhqhZmB3mMDODN/6UDEU40q7m/30
k+589zzuyUysXhIrcRWAQGoeBC7mBGQfY443kakqRBDx0Mf+K3odd4bfAZ1TrNVu
+8qIDzEHDWA/S1LRBl11+aAQELA+BvvuYIJunAbKk4d1Wh+6dulS46LyxuXMP1ty
9pG52zOrXG44C332YX1nUrT+NFIkyiqOkmOpOvA7/ta/EEHxzc3gB38yxCRjA0Ut
LblOOJUPBYjUzAayMn3YjZn6d0WWYADosXt5A63KE3Uxrm+Um4InPS7b5etCCHFw
yfG7JWEwPBwDjlZSfczv3+TFH8wYn5/zt35p30JORFsjud5jYK6C09N+tNjlO3W1
jfvgnYMeUGtRbNhnrPspOAslKD155ja9UaVS+fUQ5jBNK7V+PsNDIL2ZCQyEWBZm
WD+pSmmS0gbmhUuHzYecsyqPtLAYq6IMBvrJ0Le/E4A/XJ8nIIqErm41KbWglEQP
T7/+jG2GfrPGHJoIZJbvFTDRsGBY1Zj/HHz3eiidd/unzK50woW+34MCcKQZF9yv
RbZN17FMdyMusSYInqPHsNbjpNImC8NG7oetje9Xw/sfrMW70rcKI3lZbdSXMeQQ
+yMdQFHYtb6H40yqJWSi7Rwa0JXe6oK2qo1OaPDcastQHQfVCMU4o9L96uyX1nDi
rNlvvhS4W/cAhpEO4m4NqxSJ8n0C4+yFwKCvrNd9OVlfujXJsDsiHdxGnWrtK0oS
MfgRYYVGyxddK1PAmr35qTsm238vwYyjd0W93NpRhEnhX9uFNBOW1kANRnK8PnW2
0xiCXYxIRK0Y5nuWcvui5XNLEO/28KOzKZugTWoh3BVIg8KREvENXgWubBH5o+Gm
/uL/DqFmqD14bqmlCUevIgUvO48N9j50ouMB0aHh54ge+LmD/7o95AY9cj6qsgAB
KWuwTkxuViCygqX78kg1MT6O0hXEvKFObKoj1Z3hKaPCeBmPq6+jUdLRgkIpaWwF
sqYOnYcinPOjvBdfKbaHCerdCFc6y133HFCsll+pO5+eLHHZHK+VajceW4Ud2DD4
MWZKwavdWq6Nc7Hwc3MwGqTYOiqaOTXDyHmvn8i02N36Zr3j847e3qghadg3dYdI
ovQhh2ZP+DDPbwhbWBAZxJvLE2JnDKG4dFpIcMCB0Vik+xM2hW8z09EYSbLDie8u
CCujQ9l729AodoHOGJOU8y+a+SH+VY/mGt1WepKXolX/LgINxqTPUvNp69bvEMS2
oYxPrzM+zS+vzX3z63gEDby7MBshkRvz7pU6pofPW/V5hx/+SpR2bY9icc5WYBdN
fF/n0MyL91k8VwZcetaNFIFbLX8WiDAKeB45jm1UCsLwH88H8A/ocL5SUWmM0k3k
xhw7lK2RzkeELdF0FkZToHHa2oPe3p7SL8DI+TxUvzyY+BTCbNLrRiMm+1enOyrl
/QX6AxlYBOsZOHkNSp3G/5tYfqQbsjMCMdytNrnnJLlkUC8OHRUZgy6xuCIhN8mL
QbSyPPIafmA6SAkR2c+elOIX0t/oDH+/iN9k/eaRrXtbJ/UWI1aWOOwoO+UKAdpb
UfpXNB1gI5nteX6KQX44LFrKEWpBTpG9kURdRKIhQaSXXkinDf41CqaDXvXakqvf
RQIBv4AiwkSo1ZGFUx+RN+unozcU4X0M117JjhG5AEcpivZ08Xgjh2pXxbnjrTru
JTYAFQtQcWOuVC09gYgcGIK9XGyd4nllO09tgd7mZW0Fie6N4iOSEl3mGGRR241J
criJo/3DtlgIIhdKvX6hQEYtj37dtk9znWph8eo1LDtniz7zYTkNFms6ruL2uC6I
198HGyV8dRB7YDfcUrebzccNbUJDrSpRlodgT+X/JjLKqUfm8BmStU/m4zo5RrHi
qG8wLrfwgKwtpiy1NcPCOoCY9AcNuqPR4hBdPBnSgpMn80BGRLYKLNVBlz60nMN5
7JpKjpURmKeIR6hjsU1oxF7MJkwQU/53oTvFRWQM/17KqVochn04WWvNoowAwKsR
hwuxcaWC2eYZwEuLwmk0PfkdskuKeZl4DkGj/ypFc8ZQqlGdFZap3wUquRbtiD7a
vK02oziPemdziF21Inh3XQM36BY1TqtlEiT+WDL/j8cMhC4Uaa1+4dBVuGi45gP4
D9z25nYp7WHozyYxyjPTJ75UNWYrdjOMnU5rV8cnwjPMh42+uTeaI6I2q1farHYF
VHe5QP7+k82496fueOGFEfZJ20pB9d1OfaDUapPDBdnAGheBk4WDOxAx0Qs/Jj59
vnIfxB3tDkNe1tKxUFj2YIZtln6tp4wzb5oMoTw0Mr5DkUxL4eBV73CXtrmip7Vt
wz9KEd4kvc6foSBbDg6tWsKIgjI4lAf0sErSMyxEEmQguasAWA0oTpHuXwdSp8IJ
Veu5p2V7Y5nFh4LmRwlxQE9G+j1pUelifUYonbIO7TzFhpEN0TFfa7NEPc35swjK
hIs0RVbWOy4ptXcseeoQI1CUDL6eAcTF/Qu6yvV+sRjkPWVexmzSnNJrTFI+hV4X
a6J58E8K4yuJLZQVHS7jfMglIiIj1dl1Z46yhIxdXDWkhUWPUMPrgR/qXtV5L2ZD
wlGovX1MBb2CqHZWNi2KfmZfQ7oPiz6IrfcuPUNDQRaPvVzfcOv39CEtj2ho5uER
5LBXDejOPs8jbdxW0XUxq3WV9LGy0S0FBpaRw8WqQOBFyrf2tmCI4mLiOei8AMiP
jhFANuMwuFjQRZ8qWPdHPMTxJtwX+RwelwF+bK31mFs7C2bn7a8BnPor4dYyagjN
1J+JESTQlHwkmiU2q6TOkQR0swGSElfVCnGihzCM0l4Q/PXLtkpcyCgdGwnJ7oZ6
G4OZSRF4E4jkuxJlTXOpgNz6+JbbgjRpE/WwICpj3Lv4UefEbGuUH4u7aTW60T1N
lBrjKCa75PYnhAy2sUDm7bgJHVsmkamdA22djhHN3uU7YgZsm9rxkE1oaD57N/52
Yl552171OpusTvfCK1e/oO3Gux3AmF6CQLyru5ETvSaJOUyGOLsnz1sx4j90yiTn
LYH/1vR0EuKCDWd0anzbyEiAICitKy2WLJkMeUukQ2j02VCufvf88P03d63imkfz
qPWQMydHdilV/KBYtSjtKFDvpWmgurFYSgdj1OxxTtDSDuDNW0mADxZQB7Je3va8
+xCrKHpfc/pXpBwszIbdAtlxiG1/Bc9wrWrtHaUFLyoFAsNyFFg2V8un7LM0rGKp
T44qieuQt7zqYlNUHAleO/ZndYdwJr6X1bBLK1QJobpdBFuDJP1zDKsVVXHJequ0
6KFQzIEzD+CgXxF13y93EVBv3dd+fn5gwNom++fP4i+M18ZvSgIecBjHLZtb+xJ2
HeK59b+v6AyJvtMt1PjyQNvT7p60VO61WFXMACFn7QP3PH61vSdOdV5bFt+nj8uH
/KC9++YzTzU6d6ZiswG8YvBF7AR1UxlmN8FxWVCO64rrNXXyqzDCFddOD2BiJF7N
tkAY/EpZzajT6SK+P/4z1qCYoEBFsjnBM9iR0xyOhkqxWa3hUS23Asq5iblJQ++F
e332IZLdcxtrCsNMY+mARnMapKUmRuwckjpe+sZD66BQ+SYGr+DQFkeTT/7Bqr1b
MCkoCp6gJIo+i/lLNIA3yf1uTtxsACiVaRTTn+jlSZHrtNA5u2vcTUd1p3MgF5qj
wNeoRwfkwFpDIZpqg6Ekdj7rNZFq1rd3hIFhzVE9bzzGEmC2EjkdpfTtyc3Lzycw
q35AYPi97RrY8LiPja7nChmbSdpzxnHU4HVETBfYUqWrSFY0kzD2uXYJYHI5BOHw
3kuQUEKm+rWcnR4I+9L19q9FSwFp8ItVLACmcgV2mzYq9BABZiCUbgUmT3nyV4v9
eNIHPS6xiDz44QX9Xzi2ayqA58QbyzuTltkKNlRpjt73uDLeYV5VKWnaAYuFkY9t
Jmvoy5U8kAvI68KUAJA+gbn9DgwuwtYoQbm1rDcoRvXOw7YyLnmFhyaSLyXPIXU4
+fJelWIU6OtvsMdoNEJYKvOfiBXHzvbtqwSWPpVFN422VBCgdUap4mEs2mykCE+W
qh5NMv/INHwyYA3otLWXRZGOaYaMhO0Hq5LU6+V5waDiqucPg/9O7lpbtTP82Hjo
wJmOmham5RckwgjjGawaeMC3G4VJ8CHBkHXFNjq/dDdr1nxrpksstFsSaESLmfTf
vyrDOHexVUhPmdxRfUvsTbIDSbQxNk6g3Fbvzd/gCnFctPN6kt2LIQczDHhkQKoe
Vv/gY8OrxKHVCaCQfs0RgObuRvENbs5UcP4g392SigOUsmgFArNK5RZVLE2+Xj5b
6T4sfMttu/77Y2Kp9AtE8m1yOvVKcPapvlNmJwsTPtLw97SJbw7FGLjFAaBOQIqC
zFo14nYNpz0TVZc6TVIqPoNAuHaUFVG5T8xFat1zOGdCx3J9TxMwcBUD7LuEyqXG
LeOIHMZMcviO7gc8LlVgJZ78IjO/P8oD2x+ZV6LDrlqOxzEaUAJuYj8krrbK4jDh
is/tA8oIkyKrgRg6wjaMElfVJieo0jbY8aS9aSeqmm+voYNonPeVDUJcTn+5We28
mg4HsYWlnU+s0ySAvb16pmsxsJl7UGMIezDdQL9ZKGveJ94ovrwZdoP4nsKq+5cj
kFHxtaq9FmUXtEejTjDdeUs40q49R1YmwTINF3mzF978E0AiwttI5yBB044hZkAV
77WDQG4fRX7SaS38in7Gjky5/Hd6YCnvIWdjW4jK6o+fO5970pKpH0PaQvkYEPUO
y6WQ3AVS/3MlzYIa370E3Hg9DL8AZ8x/U0a1m4G2nMIUuyVWnhEQjjuCWiZ5qXkV
qF+NNsrThSVAevir5CYCAKmYCXUzfcRZ5co/z9005a/pf8EJMt3cccQjslBUIqWi
TYzAO7ZRgrQhM16v+Hyq8QkS2brmXkdr7Tt4SEJQKPcZsObziXKob3kp2W4g4zEG
0jaRgVRVpP8YBnJ8B8EFQJl+XGzVuCN4XTsZSXn1EbiI8YcDb5qXMxsjXuVxpQGo
PVzJWpJxw3+una/CUrZYLECB4Q7P4mNxbTFDO10Vx3J1ctYI19Bja9Q5LRL9N4LZ
HH3lt7rAxaooN5kWc16PLTeGhqcDWisIgNxR1kJ2U/ohozbP7xNF+01EACgF2NDq
junXH174braA9gejZpseQaEbdjW/vbhIFGVyDMx1lhTaht6og6dQKoPNPkVSkTU+
04OEhAoVai3jkAWOUfFWwEPdH2GQFzyHQIgS0czsZANLO51MZMxEKOtMz7ESvoDB
Bl57WtXliB1aHFvR83sn4ufN4ZsFxGMs5pOn2UK6x37GnY9KeIfCydJwdmMYcCv5
aQmCAa4kDxzun/KcmsYgY0rAjq/toCAmnWSokiEL6hb0cSqMNFe9nXiJgRkKjO4c
Dnh/lkgnPuyvmBG54kgL/xJcU1MwdtK6blmeeG98d5wfU4CZm5pV2P7bBPZjRGna
j/faFDGBKr0vx5rWfeNQ9H4vjXCNMkNuy8HWqe6qt4XuJGolLZ/KG9Mpgva8QOPc
hiWTvLFdRkwTo7FNNxhdJhLrgTwDLylH0rb36hbKkoXJU2LfDMXU9UtVtMDkZJre
9itoRgR263SpMP9PmBonerwI3gdiWVbcALehb43BT9fj8lhh8LgO2/3JxtuguqBG
E3VJjz0jMxSGacYN6gtxoHw9dIwnZdchc2t6xxGWwbeu62g5Bp0hR0AYSap010by
PTvm0Rg5dE1ooeWXXxJfRpNf8RWSyeP49zVMc4bdnIg3UPCfMtehxL6AXQtUznZ3
D3YaPohsoMdo/56kMsi2QSE9KnyBW66pmqHKoSXqiuIhec5Yuz4s2zc+99Ss39Wm
iACcs/FMWHWY8L8ebGnrsZbuYEjjr4GwCEiu8OOoqJmLf9gAQGN8KYVgbgcmPx9d
b/fmq+B2Gzt7FXQm4MMesBV7/vyf2qy9A2pEqojrs7I9GQju0bXRo+d8oTJ7uMto
nO7Q2c9Pz9zDl6+uGuLgO+n4Zfl+GOCOs2L/Aa2DrUXKSpdCgOGWhgg/SbXUumT1
XgKMFrLCkGW8uJIsIjO0i8iPBUR1hTZKzsn/T9NfH4/qNziNR5Pvw1Ufvta0Tv7u
C+jLZwmkms1wjrnXgQi26YnMznaLOdWxsmJc3/48bNhQ8g/V8JMRbmorMyHmNg0d
JjH/HV7Go4HeXPB2yx8QY5lYPLm8vjTCEw6d8WbF6z6+bGRZeKIQ4dvnAb5Fzi1s
RuhprGEJcFDN2sQNcEkCuM8/JLN9TKZ7KA67U1XgniEfhRRCnnCRpBNql/JpIImV
1/0E8kNvlM3Krk9mab9iyyyO/4zTLDxrNl6pGXjAibBJ6k14eHQfKIW2wXcHRyGT
e7ViUg3l4e80AvRyOtFMG8tKLxj+vDcQNiTBQohs9xYZVa0wWsag7sz4x+V9k2T/
IfwsJShvnTVN9TenEJr7ZlSZxlbjf5mqnukHLYDuTjykXDXr4qFKfMqven2xhYm/
gPrSI5WLSTP/eCbeMow2jovR4bMkXtOf097pPBe0+Cg9TRaUjaYBxymRPRt+1i+2
TtqxWYcabfFBzR1VlnqHK62fguDW00h0LKfle2owF1Esg4b3f+u/hi9a2M9hheo6
daCpDIPJ/TiG2+Kecx8IAL68HGEhv84BTL3dPRQl1KgcRlu18Pwl+aZ1ojM46pry
GtdrjYriBVMi0CZ0N8bsRLPfBacjHNPgxzyzsLMPXPlt+pTjHmhv9gVtFzL04utE
ReQ+0G/s4RXCqkWrGYJ+c2nZ8FqnS+yl3LnmfRiz3pI+GQLb2T1hPcehVDzWfIum
cYqsaUuGcb09ZqgAsNnmkYdi88kHw48TwVUssNQlC5vZEknhE+I9N5Yoz5qeoi/G
Vbh2v7/ckWRAwzB+FRbxvwpfKUgkkRj3FRR6WIvZQ2CnJWI1aNK5XQCtAYzrkw0F
d0jxHEO/mLcH60eihHomxvDolMd2DRKpPhGS4ygvttPuwNILhk7beENjm657pXhb
xpaVn2aUWR3NzPHXSabQZkyg304uhpQkDI0WCVkW7w2Rinr84CTeU284FH3+wGMK
6PG0q+0sNb1ijk6CkJJf0GyVp4hwWGESZQZdQxO6EBisC9WNB8wPJAgw/sFo84sy
zRdpl0h7x0ZUDx74xNgAajIMTWnFMc3d18w5l9666WLqDSzOLPZLZVwIaCYBNtMJ
bcFmlzOdS+CNUGrM0MAS7gEiS8S/jYhuMwZ7zqzi+EwVGAHpCJvaeZHqsUCLzKz+
tP360k2tX2OXg/gk0NnltuiS4qcArg6DP0a0OBaGPSuL/Qc1PKtFXJ5SqUY/zKY7
nwkLW9xT0b6JM6iHjYc2WrxGlAzfWQXSXDC+aNfhyrbqo4Nz4Kxnm0HN/7J/4hTH
zIHqr/lGbL7QW34mPWEAykiOZHiTVmdwRaIq8Fiy2dwQtlWBaNiEtbyCbOPr4W8R
uU5xUuHzGS7V6CXMCVpeLMHWvbGj/ugaJP8xbW7KTq04RkZ4jv9K+mZa4MhxeXVn
BGhlr0fWuxoG1lLoQlbxOipQ7X6SgPcM8KkWvTWlYQsxz84rT3TzzHQ8Fpeygxjb
O0yu6+aXH52/ZtDAUf7c1LSHLuQJNOm2dWfs8/JZde9rURN+E0Mq7DPYfOv7viY+
17yNYXCHvQdKktd+H9Uh7EEuMDBvQSvsnmEExbmVgP7je/WsWxoJtcirNFkJbm+V
L1gfDIbE3qt4j+g251kcdv6KxyHek3RLD+TBu//pZNIL7rIEOtZ6REkyD5/U1VeW
BJ8+R6LS3UtwIYapGaFHIKXe8hFJ5yq6KKF2Ow4QDU8VawJWAhq1Zxrpl9CYbPBk
/VBP6nmO6eugVz2SfSm8C4IX49UZrlcVJNQTckoMsoG6xWAZQf24EjRkGRthlGfd
5K4ilKDhQAZUcgX/TbEh9qYf7r4dpkHO9Ev4nifCAHL6zs+veRhHqoQtPNPxRsAR
x9vut2uVlhjnhMuENFfDCRwlF7WHESzC2EeQCEBWtN/bCD0T5S6aXCPn4XMOl2a6
WO/rsFR+l2dWKK1UexFrOPs9D0Mc927eWNVSZ+LvTz/Ct+7dYG9ZBl9e6WY+oXZ8
PfskbGhypozWufMe8e+kuaD7Ar1PA0zirqG5MaQZXfIHgnV1IsXQ1XtQrGvfrMoN
1KM19xDVNgM3dKkNwQI8uJnAFt5EzhPaQQupGz/fnYxoKu1yK3tMSq58QTGL0I/X
z3v6znb3wdywLN/d/5zDqaKwqwEvM+ICV1WfqmP+5xYVlV6mC9+yQwKS2PCUzieb
yCilo8K0Q3rWulWhcMzcBY6cJ1wK+4GGu8IYG9Y/f+k=
`pragma protect end_protected
