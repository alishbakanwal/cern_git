// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:05:27 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
B7rkddhVJnsfe/Xbx5iVz3BQHxvnJuGaY9DXL+kcC1aBDPulgWS6p6Rhf9M3we9o
tWJ3PGXcAocDJ5mYzelwheI2AtQKe4lwlKRu2SnPZLypAXVWy6ayr7NaVnazc6j3
QXdU05yEI9EtTHM1F+Apwn7Ikwm1gaBbZO3igdeRJQI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 15968)
ZgdXWuoxX/KhK1CQByCM9/0xDe7iXP4Mfp5veOYpp6FIveu+oBU61Qxkxqiamm75
0x5WpEHFDIyk1wGIp2Aavv8Xkb5M4ON0NM2QNc+J6TZP3mFK9IhFDtRqWqdUSrqV
ywhruMD0wsunUM4dMYpLieKDmpesIBjCBsn4cJYRmUgu9cQKiwtyftU2PgPjMxX4
Ml3Kko7R8b1a13UCDOrp+YnU8/r2UHLz/WT0XUB90omz3BXSaSHjCmRDpQvkFYsG
KnNs3b7NZw4NvO1rubIv4KlAnEy20Eluj0vk7x1+egVPQ2pxv02TniioRZDJa5dQ
ydbUCVUh4dxa4mlSe0/NUrS9qCbTzWJRuYAxH4ABmf9PCsNSRxFaV1gKvgoz+vgQ
2A9pmtvuz1kNkA180XPmqtZ86VJRKqZaj9ykCEebPMUrT8Zu7J9swFPEodnFtbTL
2Zww+88670wNQDAzhLTRQfLDEIwMHzDgONuydy9nm0u7GuAVbcAHRx2yiHpTdPua
D+Vphd1UxZIFPg5qKvbno64JNeodradHJwWHHcuSSolIy0RnNAao1Sh6WV8vinCb
FoqTKTnffdB6YBKsjpQ/hV+8tVhZ6IF/CSaeQXT0Un+jynoRTeEC9ZfqX/l0ZpJ0
OVwgP/39fMZI8pKndNsKKzQyGNxikWVWeA9mhIqMQK1Erphj7yP6bo8JBGa0rNx8
zAiHLL1Ga1PZy6XFJPoJ9t7SGTEQ/J31Zy3XvboZAlvvtC8l4tVijp2Tk41tGZCM
yDI00DRA7ZL46/nHaLErCliJzH3cihnanotiEmagrAL9tAgBNnAntLwyJSIdbanq
/to/X1z6MnnVPlntop0z9exH5CGahTU/IvbfWV9nXV9tk5B7UCIefmRrZ0WUa7ZB
PreXwO0EO5cLhgPtXehOLNvMSV8vOqt5+SH6h6JOnfxX8Kf2eFMox8PusVGQWbV0
B3Rpafx/bouRni5h74pGv1svP07w3bB7JRzK9olL4xOexhUvDd4Xgq1kZQXV65ef
KOfe96ArnArT0+pTjpe6VkULAYFbI79QCXhBcGn2RdTICNH/ldKk3snLTodZ/Kww
BOklz7d3YWiMzXk/cpFwMOjPKYvtjH8pstYGNXOqGJrVWd1Y3D4jxt27xH2xXWEb
MhRnaMgK5zLy5jb+VU1cfHPElwL6ekYCrvQX7OEzU+ynm0sDy/qmdlNy5m9cnLu+
xVVwDyZHleUol5rleQ2S+SVQ6Bk0s1H383ULOrqgYLpgdLdW573r2rQiXHw9+Wj6
gbXA+kcG/m2S066DCxIZX7w3AQJZcIqVl7KibISGyk8+AnGIruknktZRgre40Hmn
pWDBqfKiSNdfVSR3HiDe108aNKWlIEt68O1avuMDEjbhCvlomggekz4KbVJm9bdW
L33sWOXnbeFPYXlH6WUsLwL8VicdVF6J/HpYeQE4oMFt7pwak6rvY9Cyog4hmygY
dy7EPBheAMen6vDYPKL9/KFnlsfOlhUXhupkLwtTip8Beu8VYSyf+rTcBcTWfyTn
vqW7wgHedTZpWlntdWXthEcm2eaOCG5cNdS5JexG08DrAuWhZER9ehXnpZ5y7dEV
HOW36AzCmTMHkkbyPofX4dE2x+0uG1+8DsrLv5D/w7GqVyWgsHi1I2/w5sEwOjTI
4JpExK+r0uPi8/iOXMT53S6dYiw9r2AVwkr1kldFKE2rXM3IK9wi3vE860VHinIn
dEXU57haFkmvITGa6YPdefEDXQxsAzTPtGYgbHO32MSSgOWvp12wRpy4cBQ80GWv
dCOIxhdm3rpxAJ7G3X0Gz59UFqbeMUlixr9YLQ9wFrxlZMP5BuKFUKKaM5VCRuQj
d2ASMAA/bIPrtTNLkx9m9FlPtHgHQ6zAp1TzcfBUrZqtkuOPAFTbiKbESPEtBFYc
MZS4Gs7uAlEUsZHPAxIKTc4vveTYu65oHpB3UzabL+e4TlxECvDNw/gl8K62w1Ir
EYAJW+22lgojJVCkX9ejmsQLwbS913n1WkcLd+MnpoVpBCUz/CI8jNVIy2DHiseY
6sSJA991ca87xALZYu2S12eOhDkIn1nWn6c2Z2lu5cCeroGTKySR4xeuKedrnwrF
5ec5xHvzkUsiQfpec8TLS4prP88KTKBkPezl4IuWaPtZSvSuuOofcFW4tl4h28bU
Bsv3JgEURw257fBAydPTeHR1bEnv5+zoKiOvkHlqKn9IatG9bn81GgdtKXJrzG3G
kgaMRzU2nr6vp4c+fS2o2tI+a3y1mDwHoPWeAvj0Ivan9rfoTvfLNRnhGFP+2uEj
1fgWU38TYhd3YjB/HIZdVqPzndU3Ep81A09h+2qR5H/AU81Q5k6acOhXYvRYSZ0y
EQ86HYSrk9RvNIg38Ga1Ksroecs7q4TKgwe3E308ct4cBHOQUgf0IWRol8JGKyZA
Wm//QV0Y6QvSUYDWhFmuQ+4jeoBtuuNTcOivEV8kvFE+5jjGQ3GQCFKCBop8tnoV
UqJxQOQdpQXej+Fnh12ZNru0vX/Cs+l+rFp4PlcBI4Eemg3/DRO5miSH99Ts1vBw
tBuk/u6XqYJ0GkMxqn7KCADJC0ec2eonsSw7RBY3BFo3ERlcSoDNg8KXXGvmA6K0
Imy45nrMmCVxlLW3suYtbsU3fnkwoBIY8uD6Y7djcGeb85XWM+kVUmRhyWyYNdDU
jFuW7FHUFkQHo1qmxC6neGXeDAZ1I2HD/as5AqXbT1a0al1ZcvAeF0abUWpPEXmp
f72L+HNpWGCzJ+HEcpDnbyVEb5rob2WRkPKO8mIvlLEfJ4unHKJJ7ikLFxs7Q6T4
QDAF42CLvmoxRpwYVmbdk0Uhz9z4+ELKY2sH6CGL4lP/ZBPh8xbEpo/CjPk9LJkQ
UOsJWtt6/7xTnWxSW0a0zEa6LUghW+CssyHEYDGnjAZMZxkZMTI0m+CiCih4MDNA
1eNHvjmKwxhyknsGCld+gWOlYFBXssFvIu52HVDAMLqqhJNeFHSLeKlrMIi1zjMc
hsGaqbcdlC1tCU0FG9moKGex+YOg261BMDeB5pBKUk/sdQna7deTSE2CNSpnuVt6
eD3M7sxovBgHKSFGNzAatM3IWmh0UsQRjlvx+9I7ob+ra4dgKOMpDT7S8s0pHToT
mMFyjTZnHGc3U8uk68e7/TRM7drfNCtuphscFS2bvrergaTAHeTil33+tM2hf5wk
5FOsYh31SDaSyt+yapC0uYhAPqeJjmqb2PiSOD11NN48VbWnIULh4TvYw7r1GW1P
cJFaM/hr0NdTmTjkEcsk4wqQyRW1DRHObYXrM7qJhBFu46Jgy3wblhWrftpalmwz
IXXJ9ltN7uIWhsX60HEFaSDhEU+fvVDpjctoBKcKdJchd02yTrvKGn6guBGQy6Tu
uk/CipEdWHTLsOOH7F1/UpPemkngKe8PfciqoMhlzCXht4JyD8OnHYcLHGeE0Ury
TfsAp2y9Cyi9M4kuIbRxZJYIkRvxXm4VuSsPrYkxgsAqvoEZrxCH6S4zN5NVbFlV
qaJWKsTpu1AI2v9RKQfozTc1YoTitIQtdkwclfFwlJZWFcwvJUrd/fF8TOFWXYNT
I8zqFbtIzxk5LSyqXITisdaijLfEDT56ge+A5JrF99KCRAuuppC7znV8zcwGecUa
KD9ZEyUWfe4KiKI8/W4eFIO/nFeb4k93h/47Cm85NoTs7lC1dfyI/AhAunzDaTnD
RpuTUaftKaSonWx1TvAZ4mwwwMqCV0X1Xk0JbGk+07d7UmoNhiXkE1jVAPog6evd
DiOK4qzerkU4SyNS3JuF+MtuTuiKMhrlDDxrOiLZO/IVwNcJ8RCoN7fNWd52/dAu
F0yRZaFxs3zwuveOURp1eKvDTNmsClilTZJ8ikqtEnXO17vEOUTylDBeFSxGGTdn
K48kwp+ENIos3n09UiOM4pNbDEHJAePLNkCYNyPcchyNzTA2JsQZCaomB6sZdVeC
qMLYIjmbz+rG2ziLt+UkPQjp4zr5k17Y9pJUBlE4gax/EjQ2/Fi2TQYiIni+J/Jl
zp2qCYIRU56NwZZc+dr8rUO1mVvAR2ZNDa0aZnJlMxJZKdkDn0+3WRGovZvb8yQS
f4Vt9UsrC8OZuD+Rfh6OAqhlJKB0vjfr41WEX0H8kyUVui9dqkMabC5erYGQv+Ig
GoEWM1Ooq5cDiA7BeFR4uL5ibvUAatdaNO/N1P82vVJ6jeqi8LyRmm+3Mk/wjsIY
JztXud4fIcDUja7p13CTjnmxBA61g95rh7n90/iWcA/kZx2hPpfd8xgeWNlqrBQZ
o04fiflKh6iFxCrTjTVXY9A7z7SOqwyZmXtyTkSXsunjhOKY75+AVADwLuC9+zru
24bWVl8kfyt/Bj6fgiIXjxfMC2xSTywWn5DETuzx/TXxOkWZ6P7EVbCLiL4KgRX3
raL62BtCNIjpHYoeq3IbCAA7kYjodJNWrHQNqVIlha/MuZYoKdv+R0eAiGVPJccw
bd1gRLQKxfDmRaFgOGvquG4iIuH4ptMR1mi687KzpHf6PX7R3Q4HfHOKwcKnq8w9
54qLMFntbo+0Cfd9rltesW7X0IxhYuzzZCAgfTroeUmgrGRP0Y6dvsIzxSVRntQF
x+hRNewZ0htBcQc3iZeF4PQzePi7W/ZB4V9H9IKJ4hcMMR/j7PN5bSGZGpGbx94F
BcLyYcNf39hp1F+BM+HfYpp05pm+ZngLz0i9yHoAQY8w7qSRNsQ24vIrLRB8EcRN
SPFSapUxgbvKEzpLWwTSgDRPYaSHjmSsyV5lFN/PTsSWxe3hnOKFe1AgM+Xyp9pk
c8npkrXyGdcDeP4wLfcBj/UBg3i2qfPgLg4BlYh7nN5LlwXihjFLcZ9ZPsgOUmpU
2EXcx0E0FeaanBAQHRLaSUuA5Wpp2WOfJ+gWci2S6HEOgezAXeNwpSP97dRrpihm
5mEswYxNcq6e9PaC6ssqgasSWKGHOrl8Bv5qW0lT54aBVOIdoFQS01ZG5kb5vJSi
sJu3cN4K3W0yWkAHw7KAkeUcsrl6gd9QA5DYEFgWbq+ZV3wV25MT+wpMrxW3nEKQ
Soj+Pjzupw0/JC2wNMGUAiaPhJoUpZSAVW54WOq6i/sQplIC/9qoHlb3fSdZ1fgT
ajZsGeIG07Iv4y4T9ZDpH0TP2AWLHtce3Ziy3WmRTAOxbLioF+/HoaYd2Fn4a9PK
DKc1fTVGIXL7qYARgOrfVrxL8ZRi5nfXKVV2HweOZoGzdexaIXbFM0SBz/P4jZ/j
q64yN7T9kv5L5xBR7BAu1ZK7HS0U4OQuZh/H2ZRjbpf8H+EPIHBnh49XIIc3jx9N
DULSrjEVeARABGpIfB9gefT8iQqjaxhODqsgL/PUJY/QkMcEO1AKC8q/EBAgZKoh
5v4/aGkTA9A1SMvSlznqnQ2VS7aDhvwDhW+U9LISD/WcayCUFXVgUeQgHJuzJxh0
pqdOGF/d0SrdMrwyoqc9L9IYXQbW1T+9ees1l6thgRImSCpmWiBti+TFUdsAgbKe
QCRsh/pMIaruE0ag1nMjO1dOlkaJV/M1aWk+KyTrRefrpCN2cg2H0Bf/Gt++qYuv
ZP/nqRZUP8tyX/cZd5dTmg2Pw6WACowm/yFFHSf0N2GWmQ4kcdrX2qfNxjpg2Ct5
AHN5o7pUL+EFF01pcAA8cI94nCYI8sEhb7p0CdixErxvMf0SWO8VU0Sl9vfYxvJ3
fFnAcN85J3QqP9/ev7BHJOord/3iO8+wk5X2G/RYk32/Fss1h8OusXKOWvM6FbjZ
R+Jf31umOVhLzgDpddDcIT33F3GHWh5wDgUtKGLKBL7WOMIMo1iL3b6WPdA+BZxX
wpbEmYqttgueOSyZT0yKiXhS56OMA9GV1sVFbXGbF9b8koDLwg3eMR+WTDDd0nBz
XExiPybdx+Pksmh1XCC4RDW/l/SfcVP32pJhaIguM1LNUdjzudMI3cfu0uwIfyI4
px6MTJdKK5/JTaakxiKcm5sbYdt1uiHT3aWoORU/RKpcOec0YS/4QVVZEQB8wV8a
NDFhk+4tsO3g8vketKoQGTQaOItAw2QFjTYOKvY29OYsLOA1UUR2s+JLc229lPMF
Kef2eZeobCuQMi1D90neQk4CZ2WqXKY8x+TntoxNdr7adi8XGOkMGajpzNyk6eXh
/leZJvlZ81BW6/A4iGFZJWQxVvZEtViHyo6rX89DLaijfc+T0ajKj6GTtfBVCZLR
NgqXDZHC8PLkoTIi1IHgZzS5TVMvf2qgc1dbygKUQLhaIen0HqIEdxK+wniIe8ux
3I17MeRxVz+MkYmWReLI/bbZe9ejt0+D9WSSI1RZWc3MBqYYcb/QMP2ftMw0f1fs
GQcary389wowLDGj+JuKntz4K4kXJet5CYNKetaDplmmf90gb1oeFFi5zUQugK/b
MT30c/FrnpKaEi7QRxXkg0cwfpAuPtbVjbDw6vR/mOrj3fDj/d0hmwZBd8NQ9qmy
g9WHdydi3TZB9XG8vhO34gM63RrAPfAg5bUfalk/yRN7Md/cNGijTLSYjL2bXOQC
0m2ySSr20mGI6zG9jMWr6APgs4XiFW0xKxwTSsmzN9IKvVrPoytKKkJZhwwmiyxU
3PcbJeOKYceJgHlKOKhHQWY/9z5iMw0gUPPzBl5tK7NLcaZLvf7nVSA4m5U2tcxW
TT+wu9tQkKmaM1jaEtCXJlvUQyTpm0S4bTb4xgKSlAeKliNF7l3HNUi+LcqkCiOv
DG5WDv8SL89HGZowTCy/h0HWbrgIaoOWDKCvpuFWnudA0Erra4jM/03XqLp0SMyz
hTIA5P7x5QaikR85QmBXDDnn3NU7DCe5Wj7XbvS+YDi7LYgoT9HOz6HrihupRpY7
Kc5MnyVMOZOQXwCrTryYSuqw+hymb244xZojwAgEBnLkNcfQ6YTpYdkd5jHYgy+W
0T3Fp9qjMDSSxDAEmhuuu5MvDMXBu1Iww8LyaU5J8iQT/FZgxJLKKMW3/ZUgi+Na
c2y166+APetpaBdFv/K6okeKj3pmQtuvEXqwqknYy9SngT7mnd631TAR6ohrQUHU
na3rV3q9t1zQ3UfEVEKjtx136AoEeEDepzBn0dv6W4xF8csrn74mLuas5huh7LwG
1K5lTMBzKMcqNZVb2ESpSXYTa1/qIdxKn7ec7Rvo+yvPreQ1ValbEu0sfPXshqSd
Y55wDPwMcknOPPQwJ+moI20ZA2f6isdGUBxNQK5kBHcCEhfEaVnLUuNQeLg5lNJb
6Z/ijT3sDY83RcVw99GAsEbKuFh3GIjojD10VeJlRwqaBTFuSeaHeA2p6yX0iWGQ
F3XjPu6851irtnvoWY8zSxLNx5MMYX0oZUx5dTuqixRqoOVQLzYV/5EGj9ERIfet
YEj3GwdOYYhE/OE3SQu//6xAz+XgRvlbCBxE1hFmN8wlAbn019+E4m6aOiYH5xPS
lnqq6jcXmcnjozdGFP4blMQMaOVjtEjdEOPz10RsU4ivaAeXDDg4NGfCnWhId8EX
fk0EPQWrVj6EjW+PbPS6boret/qQZ0i3G0xztoPsFunXPkhCw49fIundEDcoPrES
+ESJrhRoj1VMs8iD7J/oIiFicQFjjc2VcXFdj0/+srmYAlkP+rgSjRo9/NGDyGOA
Z/tH2Nj0TcdklydDCRiDroMv1NthGAhNM2rw27/d9kR6QsiBmrvZdeZzyXw9PNY2
XDT4/ERCUFdZIVNbMccDzlk/KbSglz4/kHOnz37I7nF2xLq9vvZ013Q+YJ1c99F+
ht2s37Scuz+Sv8CcNvxI4PAU0ZHzqI1hx6v3lAbzbPe0xVpgZLbZwqlnn4Od10Ta
dRcrIchShziMmcXTwPTrkhuS2mM1SpfTFo8svxOaW3vzht70dogz3mEyXz82Nw8H
9RB7u31fBlXhj/Kpc0nFHJmjuPiDfR+BoM0RzpEaR7AVFenj+HrZNEzQehu14xy+
dBdPpSw+EW+T8A+oqeBjGl7PyOxsfiowVcmSdpQ9npHitIgPoI47mwCkHvMLV7PC
UnxwtExh1IZ/NFeZHd/Fsba38rfM5REOsp+Qv736eBi5K+MqemlezyhFgVdWQHmk
7PjCc50AUm9855irpj6HYvluKgAM3v1H1ddeW3Yzbpwlc4tCb0MrO/YLa6XekbJa
CY8FJChExQotDjyH+C50FEyUaM4H0Ajss6R0XhqRqmX4bxchYOQBn03oSIkm0EIn
QR6x0DuRb763+mDZa0tVikJkL/MNbyR9e4AMgtXTkaEzkKM6jVp1PiBUIqaq3CbN
+fB6X7dxSuCoE9z2sBA5xpOjNi37TwXq8r+zQBKPkXPhmL6DQJqCiRBJ2pcc/KIB
DydqQ7THrRibI6RKt/gL5dMRWG2C6ujyaWRB8KSqob45y3QA7k10NB46M38LCAg1
6EIWFFbKcqmQtKzWCCEpyv1+AsdvR9QiiayRQwu5YcHltoNB0yn69OK2XG+D06dE
Hr0HgQqzaIoZ5S6TW0BbwuGWaNzQSyvXRU0nxBJkX9Gkm/KdnpIdPI1gWGR7xbsp
p+Gh2MRCIrhGc3aed6rShDqhOdh0llXht1wRsReyLvu0ok125NNMrd3Wij/OaHCj
PiI9iSmbTrFlL8rOvzw6kXUjwR6DRuZ2L7nzvRQPj5+1szTSnkgCqRDOKGyKISRE
Nkv2rFoPq1m1GoDgjmrPM0ZkY57Jhm9TdopP8C331LW2W3YmUDv7Ppflmr9WM+sl
/pF8/kr/PCSucEZRNzTaLdnBtnb2hf/QsG4gpyRJxKr5Rd1cS3msuLVChd6qPuYu
6tCHAEhjJ5DC4Eh8aoBoqgdEexqpppvcZpq0H5sKLmp6LnAiQWGqxNDFyayB/ogu
hnDGKBf05tK01DgGWu7bieM7bwajD4tnyIhqgEiMuMFkkPpiY0X+FM+hQb/GCNsH
Y1COCBohzWARbJsslY+WcOxdUUBSyLFg/+Yhuy0L1udarnt0dUE+4f5Gme4lKxPP
WwNOt1UT/6GoY3s8+LOT1eAqpjuJWx0SPSg3AADvwFxhyrYXs7NgUcl9KOjDOclc
yvWawDZs/ZVUMe8307Sa0JRiiLYhz0zAPK6QQdu6Mnxv2YTEHPl/dAp0EA0wseGf
ihubRASKxoQM5WD4C0KQdDVjAM6yHCfh0hfsXpAMgZdPb2GO29OfRtSiQRty1nWA
rakJQ1NusrFLWwdOnsZeuqEAinUVta0q1JR9OecstRgGNU/dGAwQ2qJR4gMO3Hla
ekwQpqB/fyQWQspMvhsUyh1lIX75EoTt2XEBWDSlilBk/Vb4k4RPEJhfR10WSW5E
HZa8e/bR6xIuFDTpEEOSKt8nRlcV9pcqot9eeHc5Azz1zr5N4UZRDScixKSHOkFg
0qR/wiIkMoSc3jnzqLwQFj6yPPekQHIIrM+Cpj7Wm86ZzpfS5NOS6mw6Sb19gIPt
W3qf/zzqYH0ajhX6FAHr4CSOqK03iuDxqYp++f2KpiSJ4yxJO+8W2y5AaKneOhyU
eb55HNQdiiYoFbcKgOu4MG++r6mWaobL+nW1tvznvse41DtKL/V45JxWaRKGLwDF
6AvhMubVbTJAhdeffJzly9M5k0vbj/ZKq9Ze6tIoKmU1FhNpIgl4F8Zn/DDLu956
9nmBWmRb7BDFmqHYWF6DfEZlKuNQzYkV/l3T9D3mPzbUuTHd+IQYRTXYlGW8YUAi
paSouIBnU0ub3KlsGWLCcthEaLZpCyn2/lxJ8yq7CTgAPcTTVFcUsdOdwBcAuhoL
2gByc6jjkjtztjhGfz4vwJgS9I+TrvJdhIVwM7AEdRLWNhHV3wMLlglMdmC3ErfM
gsfdciF+OZa3bnqBpQGMQ5eVgaVvZiCim8RthMmAAZnYuMpJSGKb4CzMZtomx4FP
j++6+5VHgbPE5Qt838KlOArQbFAh+AZMPXA+X6vTXn9t2sbVgpB7tmwESFS5beMX
0rHIlLYWPbifoSlpen1jgoX0kVkfQ+73D+jz2U8qqicZO9kvSqmqz5GYtIho2QIK
JSjz+azuqLu042pkMG18wyqCE5yb6z1qXQxKDVpz99BkY/rzgJKhGsRC3cYcqNIn
Kw0jmbyGmf/0vDY85vygXjNDlISpbDrmUlRIBbssVGn3eIG/P1zgqlFf5Tts6wxt
q/415gNGSBowCx5f5mYwfFoSJQ6aT7SpIVtenx0L3EVIfRFWa0PzlsTdI/mJlUvG
dpB/EHM9i/z7h56K63iwESyznDvn5lcxW6eNgBQRwba3qWgvVL1EBqxAY3mRtRuc
vTyE+dZ2yCMy1UOt9GIvg8KGnttLApZ30dmdwAKgqEVlBxh3geXBFLA5/aJUjE8I
TvpP3qs1HE71y7Tf2WouHMJ9OcPYoVnG9E9GdH6/pclgBWcfM9uOmIUOMYBzC54k
4VR2ucmRQuhoLBSiHF9kSkzyh4a5VzYyVHRIKK4S9moSnBjej+Vr3O9OJ/Lnii/w
/WS7+6tgVq3ZBoOl2HxdWFM4HC+IaRVQOcLJirJlljmptKmmrnApuyTFO8Cm+6Uu
X0Y974+srgexsDG1NGGtAnGgY653jP/gC6ID5BdXeDidYn0DlK9dFvDVL1giocUV
SHkYuXBh9faV0eNTNO9YdVgFS/lnroaVN6HXZ89j1MMwZ0U67qBaSIh13gaHYHwS
Au83K/RmDpg3hH+yEd8mA4PO7TY9A+PzNIvSP0Ht/242RBNQ19wrW+DcCnNJme5n
BjU0p+hs8zD5zgv/J1+6iZYUMA5LkUKw0OmWiuBQHH+3Wyq4pfT1ZqIZYTCzveqE
AOYX3YiV8kjKBVqbGsYMSEvIHx6cqT1FOH/HACcy0rwF+Z7jlWkp6TXuqNmgorkh
RHIjfa5Am1Oww9rLXTzSuQ4ziAPUjl/DDuFDCFNkiclGfOqn/SvADPeyD2bzhkG7
w+nmZPGA7ufunuykRYVwhbb/kMWyKgr9j4heNe1H3+pCP6t70SrrBpSbD4ZAoCnt
iWDS4+gTh4aqZLgSwwiQuMyR+fV9H8wElJduofTrw0tLj8WAEE79MyZ5Y8GcpIZs
zc3BazBGSh4V9TanXjW56O08TUzhk5rBmWDJ6ECSTc1KQMpsCw2Ea5GV+Wo2TU/F
w/oQPdstFjdOunc4ii3+WxsBIaxVHaZxi9en1WlUU/qfsrx1DfvdMwphef79d9Q3
SfaIO/+gXY8iREfQOhFpfRxyJyPV+v5+BjMJxHi5qT2xyIevCo8YUhcuv2O6aN6e
AGS7a/aP4SZwsJZzru/d771ipBQqCj7bbj97G8nOV8/2y74p6s4W0v3jPofk5DBb
1x7Pnh8030plYpHZQE/4ahvv2ZpgA9zws1D52N7Zyex6p6URfee0ekeme0QiZxmj
uMkfYgv9WrvqnRDpFfFTkviqSu0L3pSZVpjrBbMHbvhgzERInLL9Ok6vOH//uKt4
yBse6a7AFlNXRsSZAe6IQryosjWFiEO0Eu7LbhvKydZPlWMrkRDv1F/AD3isBiBN
lh6Nt8UbNBXOJutN+QptHAt1whCXEHWDPjLmaWZ9I4X9OjdZY3cdh7qaoh16a4l/
IfS+bVFSUumagPRcbGfwiUP9PA0ZrJKngdUpy0DfLti6JpwThGW2wamepSuI2WD1
I9ExIEGqJ7S/HTTiOrPjdRWAOmHkbD43Hf1yjZ/rjW73bCqRv3a21u+LGsak2Nll
JM/2j3ul71iXnAzkpZCwZEUpczOomGylnjE4IHhULjtk0/984EBWa80mABOgq72g
EopaJCo4YV4MsCPWkpx2h0S7FjTX3fs/bvydFQ5ftxazPD73PiU0gFyQA6NXjD0T
LOu9KXAkDL4ObwmsMjRrVLb7HiP6WL/M0nB/KvKmOZCYB1w4hzpzoX/t8OTENgqo
VyUmuXPjPGYnhgI+ApTtWaaV+5WZSokL3VTr8ZsQpcqkENyTICkQM5HPPXdghtKo
5bdDCKTgPpJquBXMAuLlvJ4VBpjeaW007svENZ/qkfAEs+tPbc337dR3eI/JFcdm
DDWnlXn7r34+PGcPjxfvU3EVRmyj5sFmdDz2L2IEzZ4ENj7FXi/5EXuroQVJINZQ
iuJjogIymQWwpXig+wgA5ZjH/0wGe9gBi5WulFNOmifYmsTI14COE5zesRPo/dWS
7QshOYjoONDxO0nQsCpV381JnkFy/ih/aEYCpBQ941ca12JkyX7KcTPYUuuzkB+X
WarURtIcZrWQ+nFsHzPet133ElPQwNi+ySvX1N0wQ+RI9kGr5fZAHEdHGffd2KZg
TQmZSbMuYyW2YmFSGjoq/k8xr1I8iG2wC/fwbVGu3IZcT7TzXFucxTxom0JgzLYY
rTecK+sA179+oKEjYQzUCCCrc93i5SNTnNUqBn0ZG3m+k1HmOI8HiotkxaCjpQuM
ZBJ2rIM2aRlVd+f1ZPG79E6XE/1173Sb5t4srqBmyzzShNGD3bUc3eUhXFkM8w8o
1WoAyBi/smxPtbbIEeqFww1MglgTQRyFhbxYC/2zH/G8Zlr9HdJy3pTvY8wNVYMR
FK0IZBkQSD8guNMBJrzBfd7CfcIchI5eMJvPH4tHDK0ygfPbgrMG5QiNg2zmf7Jp
amcVHKLDm4OdAAU5tdg9t8y+4m7rFUpdhCai4OD01sRRmwDVaHsahtBbJPEoxXEa
xrJ93XibEWodgsaCI0NM9N9JBtU/p4AtiTapEr+c6zdZaY8xwqpZI6WkgCqpy7AK
7v5yUYugmjrVWttMnwXuU6ypU6pSokX4eTQHuUJBDmoSTzSveAwX8redvyk2VXzY
tN2aJAVmZRf+VtTG9bpE75caOEnucWHokf6fT6LtX1lL9MwiQlWipBGRh4bUwUnf
rVgBbl6wcptrXmulIMRpVTCMHWcgz3KXNPWnnCPZ0q6+7pgQaVMX1iEt6cOvU4u8
+kPNT3EFBECocRehk2UKQPw5Z3GKjuygg0c8HrjMY8OrF2hQVEkDuu2bHoNz0+C9
s9oKnAgjD+VhmElcbcAAOHI3YfahD6YdUl2J4XY+U/iK6a1QKOof9WIY4xJ3kYWO
6zninGpxhHyz1I6HeVqC38ULOv/jxKGVWOEXkkSF111hVptrnDRLh7nOtKzCCLsB
48XcyA83cAQgQjpZm/m8x6Scw0bEx9x2IFxJ1jvDnE1W+YAOCTMv4J+UAg5WZaUa
6dwGp8qQ2Lk7M4ausZKKRgGqgSKbxdsEfM354xR0kUIToyd5OlX9/12jtMDRXf+I
606bnizOC0e7+tDxhYIrIWAUSaEJPzRokrkMszL3F6N3zRbby/9ZmO9k/rBDlf3M
/2qB5pEBVD712jF3wIu1vLsVFgZs9RR+gSJX4g73AZexSXjROw8XU6nVsm2uLRle
9WhUkZkeMaz5CmPZCZwuSQ7LwxqWEIgwJB0rWUtolRARTlobErhQ9qJxQp9KSqAn
WdFAUW6gT2t3h+au/uKdbibauGn/EPtd3WhKgTTkq3juBowXl1eC/X6tyw+0bf69
qO1ti17KgqYV9t7SauqSPtyerRsZdFslo83HljUkZcDquiTrTe94I1xoDN9Z+X1f
ziW7INYskmqVFuESwB70CS3I2LfZntTvSGy6C+1csq2X43mMt3/7bDcRd16WzbZl
UAldPduFQ6MrsQFxIHjOI3fwakae1K3msRWascfjeUxurULRL8urJhU9BLtMxuu5
f8O+gP44L/zJPYhxfDLp0vPDFwI9orz8De+o4XhWgOPzQ8LvrRjcDQYOKrmWfc8u
A6TRzPp/n1UVSl7dCb/564vNULOH+ktkVFNtrwbgu0IE9VS6pN96puxOqP4Bq0Q8
FER4pROwMYXkJ7gcCQYmd/vNy08N/N9rzOQK3WH48tVvo6DaKnvQy3paThaYd722
pE+/wNzhwxz+E8RmmupBTHqaFeTvWHfRhOntjQNxuyfsfUNch0SMhEVAHpasFOap
XxSB+EEdUul/y20evhw/xF1RAiwpjWNXZXAfOKZzS+N2lvPnqgCFHnXbaZ/PXLIp
i0VCptmD7QZP5RToim22a76ulIdBtVXVFe1cUyVEwCPK1YsTMWQbo3usQenWJRSF
tRXpm/WeJAs0m+bt9D/WR5Me5gCQ+oe5R2IF59dXp2rQutFaEc/9YHwbSk19oIRF
d55AGY5fP2jY9LbNOYjtDyrk2LkMhN/80veTMNykhdzAQWloPPTs6yixTrckr9GR
1S5EDqcJxROCQTPEwpAkZupJcXUEQHw7q5QnryQe3ULfVcWqwtc6P2PwC4Q8Q/y7
Km36sfVJBSyGHm4E/cJHutUiAfANx1bUeknQPDaZawxoVJvtsovRgqO2G6fglIpd
jK6JCFy3Xcg42SWpIDze+HMJGmcLaZpV68mBtEPL1/vm67xRObDKbavHOMSxO97T
CqIfuh+RD2/Ly8jSeWut8GELjcNZfEWvPkTd68uUQpUSWVEP2kXwxZ9vBmVecXWh
hfF0K8GYABm3wwsHmiroqpRbqmqHNyl+oLHBZWYfSjOMwnpeGT0mEeH9h41+zhCG
5HrRKCBiiNypuxb+p/Zs+8azsVkgHI9eGR4matOkUySQ1dm1AQ9wP99t7guYI1qT
f/RoFLPGFL5HkMfEYiENGvUSj2MQQvtQjxgT8R4g/DsPhqfS23Mv6oYXsevktOP5
thrsv8RdixMUqCHvFjDzjIFrbHNOUZI/km+eDQ9ILHKE+gbcaJQR2FtXkfDy70bS
y0qjUGNaOH6w4s9R/gmlR765qT5/a/zUPu5b7k8xWuIXdrwxw9FB3BlRpuvduwUu
tUZiPqVh381c6Cp/VDAkcybf6lTu6HAKBaAU1sKCNHtmN+HJxURMp5lTx6haax9W
zr07cRpP4SgTl0wqCpzvAUZgTHKX1/vjqASSrOUggVH5ZA/m7PczkgbRlF5ctsU8
8ZloqMtSDnQQ1oCdRGeR4tUmD6ngNuqTBI2VYEHYSeumRnR9RnpY3iczCcvlcdW6
sjffCxgc89VKZyikLwwqUOgz2rZ9/yJ8mI9RmakHS2ukRoKz/+XPSO5XSgrWDuXs
faHN/ss4EPI5gi+eyYzBAF2VrEUysL52+hriMnz9k9BVnaLcTUqQU/lseLFUdtdy
ySGPwZcxb8h+4hLkAheCGxLsR3LnNt51sqHo0i6OioenEj4zYvVGWJ03oJUAFKcK
zKEAFAc/Fxl/JMPLBKwIdA5MDiZL74U51e+rUJwiUuoFTefMsaHoeoq2a141TKQ/
/IcZEn1PQelfpSR0z3bTrzff8u4M6JdunZaqlMOvPhD9NhaC5RwRTjaR0mVQH1xh
jrudBW73Aeru9HljDwSf9sujbbdow8uac17PfbpNTDmDy7zNTcBJwhq8P3KX0ikD
668TlXrmcGXqcJTy0OFUGKNMUaafQ3ac6Ld7c4nr7M5/SBN8C4jCxJSfvybIedDd
BvI+wT4U6Dh8GDE13sh1ELo+Hw5pCYA3NQEPBZHlqJfWnjKj3aOhydFmgaqBUVTD
jp/gypF+l1UnEdwF2mOdpvodAxe/XPRvtQCxm2N10ROiLhAxU/9RMolQLg+KACQ2
R7XWtBquDK9TuGWlMigSJ1nXw0OQzJj84KcPYhveFVSwvN+JtftxKZKWJ/HFtI5Q
IydKDOt0gy0DAUrdGldHjMursgTiT9DDWNjP1Az2A6v6xpT4acFWz5/IRrcMEzik
X4Sn7jfDQv2FhrqlHECMX19xjSN4adR9FOF4/hYciNqxk4j9SyUQZV7hBnaFF0k3
s2q86pT/FfM84NzwqvonxS5gKsgfpiv6ULJ3XXPs5xo/oG2fZBv5X/H2jb16p9yR
Bkg4BVlGecNux1pm/9XkkSvWKeXUJAEDb2x5EF3jg5PZ7SvZxoUIV9pOU2IBPvNc
+uZO3YeM8HdPjVm/+I+POoZnlY9SFHgcV34u29DdOCWZOHps5HY36vG3Nh0SRrQZ
eGY2osaimHyYfTloL8+0fXA1Pm76urY60wWZU8eDrVcjVct8yrR74jKL7WcKH6R9
fCho7lg8ZBce1r0EcU19NSkSGg1DqoxaJKiv8hHNa3QdbU/BJMfH6TqbgtnP/xBF
w4mToeQc+kNgI+J7VgcvMWJp8nhLS+oldcl3gOTwrE6/ieAlyXTECVf0CxTecq1M
6mMFwnh+tv1EW3/6rdET2l87q/l5QnIoHr12J8iCaDbJPljFgkNCUpW3tVUrWATt
QTryGvu+vBihXqUJ2TTzlhrmgpMxAtiYAA1zjeOo+pE0mttcsmRSpOdQQASYP6KS
6QBLCIeHpKFWk88/mYS2BlxwhJ9mNLjj+GGUinAHZY94BlWboG5YnndQsi2yrCYM
swQr+41A9VpaYu+Na2mnrD9tmA/hpVk48ei7uwN7k3z93Quj2QQ5D2cUkOpd1yAC
x3H9lH8n7NwceopwA+Cfgyw+l2Mhgmrjn8xDpzlrxstM926FmRNTKhvHTd2O9jN1
JtisTXapcGx5TqOvIdi5BYX2dy9fS+kVmLK8DyRVKSvS0x6pu3XLcGOuiuYWnjUG
lozdBOOOdnxyHgwsrNyFHEET2b1tqa1N+O1+cqJsBdj6pp5yxe9EgloB3FBLR4tl
i9lMcNBrk6Bi87DQWMN59QtzoLpmQFKFBygkdDUeBo7hDZ+21ipUdQrq7PeSQtoP
hOI/O7uKCLoeYMPaagq4sXQR36g89XKR1JjhAhytgIu4JTrN/j4BG40gxYez71di
ucIF8rzEj3V65K1/N85vepWQZfX2MrOcsCPGkhzStrP87HUu+SiJFz0zdM8GgsB0
2bflKZ/hnmK+R0+X5UMYujRYGgPvGBrvP5j70nfdFykQKGX1ekK30GaME7U8Kczz
4P6K4sbTOWHjoewHlZhslNucxPWOjdAadWSj6HsXhfCn6MPvCYHG0yp0kg0OIj73
FU5eS8s8zO/YhokjrNFU5lXh3DXLOULRpQefzP/2JFhvIOAgMw6j9dpg+4rIyQJF
bmXT+TZlO6lq2Lae0JbnsqDZOQ5AQiRtXjY7LDIFep/uvCv9Bh9wQqI1UxDDdA9t
m5x7W23yMSgkDBTQDSAh8dahKksoD31cd9bW7ODVItWfHAxRwbPdIwLKZ6/y4Vbg
TD8gODn5aNGkwRm3HG/OTepvy5Gg9s/Hw8EhWIK96McX5itskZC3fmsxw+pzerMG
/QsuBJQXuQmYTfUlHn75GCCRLstQL8pXPdCduTVAaZ/Ho2trAd7pqfGBAF0j+jnu
YG/jLDsNRCniIIRHrKGy97q7w7SySGPkGgWAY8BdfrLoDMAfeYJ/QjtXaZxGMxY3
1ABP3ntm8UYIas+TmBZKeCzS90KeUTjT95mSPUoFbgMXsbZ94e3/YJeG/RvoRSIc
c/im5thvZ2ec34Pt7X4ARxR7/ikqf395xZde7SQfcskqkFA2kpiArQehOz3Y4Rgv
GQmN6AwKM0ioXajPh1qGXlJ7VGliRSZUsRRE/2V5r9S2ZcDGOrqTRQ7bkHB9nnaM
cofwMu/SO87DFFfSTslA8zCAsYoFKoTGq026AM/iXM6Ut2lUXDCRpSz5QI40McaM
9D7Gikmt6p15Mw99+z5bg1O2jFWI1q1OHgHIJFilLN/akGNTxhN9BvpvdCdXe4LJ
zzcOgMu/ZlykJP6wrxscFewUB6EhnqqKAhcNGe0ZAZ5EYj7zgEpRJ+RiVe/WD4IP
UHWpLtqR6rdGfy1CBVX+7Uoxe3XKRFzJUC9Bwd2xCJeOQZXuTDte9loVs10mhwNc
9ck/q41yJb44LxCVJrXo1bsEB1PFi6FupnP4Nr1mLo18rMPIKVNhkjLvAp0R6tW2
lfC0ioVm8+4rAfIlHTTOmlbOBvcyjzC0ajj3xMrSd8ye+FSP2czNfNxZsyFfNVSm
Gx9TkE2pYnrdxSLVnvD0ZgOwck2gf63Ru57fc2pdRMQwzF5/DDaLjfaUCMSJtF2j
WmVvLvZe/zO9ik0DFKgiEKz3R2Ct+w/vpeSum1uiJoG+kQGGu015j/5OjuOcVbp6
BOy3K+eVqHez/sB4P8C5MMqgwavA4KDbvCy/nhPiu+DsuJkl2V8AEk/ffsnYCVxx
ypQ0PcIlE3P49scUma+QFKt95joflaP0V3mq81lCYkOgGm0Ky6QHNlb4/zxGOkRr
d+HJTbucxL4VwkydlTo1w+0fMl35+WYwSebqPWiIh8KKjcMl6rffY+B4iPeq0K1p
qlmJP0Obt7YibkPzgAf6batMCQXJ7NDzbtm6j7mZCZwTXA4RNYlO69MNctJ76sVw
/FUmeW74yN5YrH2pypOGDQoOqfCg9Ae4yqPyBOPYRoflmyxO7c608HGKvGjIHqT/
eO1CelguukIxAUfcMMFhbofTG4Sc4ILv6S5OTbVP5JYswAwFqN/MrFEPYxnb1tG6
Xg46YuASien5mkGBrya6ko1j933zZEcuCHNpgAl8vy52pndLymz4q2b0KebKBORV
dsRo4BTH2Ut2bRlpQul/hF2rfIOLRKbAyFAfv44/S02unIyb8Vvbm6/Zu1m+bG4k
56tmoSPHWWitZnf5oPSxzvNhcPoYgf26DwPHyPEDNXKHwnUT9XREgH2MT6KCWEjv
t+X89DfdALiWfjJDpX+SMvigr0VfoWUV1XePUwC7ESU1Z6jie0Pt5UJOEpNCNgjO
Al5g2rP0yPcx+DwBRDibsMpdo0NmyYqMcyF+2eLXURp01PDBvqtBXksDh/hYj2Z3
GUqAeVBPExJYTRMnNQ5/1fZTkhKV4eQMlf+Z+sfmUDra7/OG2280I/rrkOITxqpQ
JaYrZnyAarkAbMwlS8OIQjcW87VbdHQQIiZc1Ie0UQ1f+6bSu8zXY32w4BnG9VlG
wrCldg3u9HJzc9tess38R5Isgavv2GO+gFXStkhItn/LifrSNtYXnvOheTZFt3jb
qg/RHmjw03LYNn5RG44WA8lFspHt43ysFBVvqP5dEsZC8IwjnGaytUSBZzgcecGR
1LXlVC6JVuD5rjvtFwrzST8MbJcSy5zS+KlW0pUXGkOmoiPxEasKIIGqYKFwsykC
yCAnWg2RdVn1Wa8Ujcc2FMlWYlSSQuq3rKf97elLZSgxRItyRlfMfd4jHfpAd6Gc
dSnGZcNnYZ0V5YawKE7c/Ugsyb/7Uwwzquu9a0ioE/IGSx/Y1ivanaVVQ+ejHbp+
lc9llClIlXyy9vXGrLTPjYoMAw4gQO0GYGTa1wb3iiPZ/GwvXMHjs+1YVXorsuOn
OB2O40fhMClX+LyOEWkM0lb9U2M2/gnW36xI+qIRgPu2uErGY+AD59omiJ3XjJ0R
92ezqlwJC9ulSXqiV6HxD9+5kYPLW83PVH/hUjuY6N7SXKYlRpQN/ZtCuzM6inNf
jqt61wT9qO1dfbXGCi+SmZD/ZV+YAlJ7uqr6yaC/izYDz61pAI/y+Zqu+6zQqCKZ
kjt2z/C7j9xbNjqfI59JYcbpY0ZaDPmW/ssMbkpG7LSy+fbJzIxtdvjaFPBCVn3k
c1p/2FPPNPgSfmA/h4sEhibWBA3eQCAy6VAS7ifAUMolhaVt7+yogwJPq2bxUTPI
vvLzutnOvaf5tEKRnAeIgn/H0cimdak0LFHhkG2KoW3SjTbg5Ux19SUFA8RH5QYW
kRnJbel6hWnyQv/wPJCTB7gcseY6a9m4pLp7ssudVpeFJ18Z/ZjUlZusAI2RVqbV
Y/rB2/pkpEYXfAyJHz/IC9AlB9DQxDihyfNk3QfTVGq8fQOPHUF/KbOfvbDMQaeG
PBMYVacHGqlFZn1gor++UOHBbh/mW4ICPCsPym0Ca94LAO3LxgourD1kNBQWT9rY
pkZtSiK6OEj/oJaWgUewmeVptQ97kAPX443ZR+1tfoILq5u0uTDR8BB9C8YxIG7l
erwqiGe4/SfxAunv8jhiS63knWthf5dcbeJdzTFKdQLUNiriFAssJw1E+KPPFFfK
9x+2JRLB/abQKkfYkE9OPLunv7XC50UVvG7Tx6J25zj5dMz4W21hhr9WIz/zVwL7
ttJNlQyY4I+V37ZkbRRuK1H6VPBm+Unk+FPsrOxigqZIRQfRuoBci4TuRIwbzpSN
r+JXWgkYUFj6Bx39a3nSVITOWGccDBUsgd9XcmEdp5Qhk5V11VjhzTkUtJTt5xcw
XyLV1EWUGQUKCdjWTEfpyWEUpDiJ1nvwfLDlh+XFRbVXOFh1Mh7xrhqjSOU1kLfD
PaO71xU3utuEdcB2pRqiDNTU5Whho9/MpiFIh87PrTAqQZqSRZQca91HQ0qEbYie
5MQy6pKZQEGXlYcxzbvnYgydq4AVRcIZz2NmC+N/86LpJmAKcYQfXgJdHB+YSoij
6f5KwPRcUsL1qcZZFwjTg0/YDTztKHsuKqx351K1Qu5z8yjuJWQ2ppFcy69OTEtb
FnGZs9Dkag7w+hNJo9eugRx9CSPfLy/Mk7vgbe5pwzfcNANalflhfoxYUV/BVPH0
38uZmu7ElRVmggJhDUFBMWP/rZBnm0kDbECTMh1Vd49w3rWuv1/gndERc0RjdiJT
fq6FIO0SAnP6F7pnoHlHQedDYW0iV83TlnDXIMqQCwxsHud62qLtiT/zmPB+Bk2K
aMhS+RJgDCnKZi12FKrHaLHxzUZtquawYA7wLGs7yKOhm9T1WgDTL+/F4snVE8jI
rs5tXdDLIiWETU9i7Jz4e9wCTAsrTEO6Qq0yo7o7ulcWbtE1dodqtn4nA6i8+4LC
y2N3ZoJXqJ42/xniFkcKY/AX0gKvxzeS6QiL1Ay9F4Ge1yU1uuSJaIHWLIka/acZ
meniZJzlDt3cTtrVtguriXDNqtYBiKWvCCD9utSTCnjVYL0BMsn033Vyr6x2cZmk
gaaBZWBjrt7nhiuf2qp3F3Xp8GokbjNJHJ+td4ksyzW5Cxw3uQx7FQh9uWkCmi4a
j8DtpA3LrU8zYK6x3jtW6otMejI5dM1Y9n1ZQNLhmKDUEiuF5tItNjbfMl8EBOrr
R0b3Zs2ooQ4xSleTgSx1fWYRztDXFNA86KX5oSx/jci+ZQ+o9GXOI6KTPQ4A/suF
j/QD0kMTiv9pL11GCuZQbCG/ZxGK4RaBX+/FS+lczaHP/ErYwq6fstbpzPIVEd9i
vqegiURga2DKP1qr53Zaza3l/HF/Y78ogoT36Z8D4/A1xvrC3N/6L+QnclPAMSXJ
IJUEP950MVPTK5LIIQyJqhbefEE/qRAHMNJrwJmwR21Amep3qonIPK791QgJqxa7
W8EYg9HzYnyBKAHKj9tNW2/rurOaI8dm3gutmWLoYb8z+Vl0lsPysBqGLM/GBoNL
cAJ7dmSOuYrzVuGEW1QX9uKcYAhgGELXcaGsaHgcDczz8OqC4DQ6gL4dO1xgyoGg
dzveceZdS4ELFFVurjUd7KKSB1jUBIYGd1YWtsijaqs=
`pragma protect end_protected
