// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:02:18 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
lQkChATvNaBkf7nN7yS452MyTIN+kxvQwBzcvR6FsWAwt4a5iqAl+8nxK2RJ1HCK
w69t/UtVpbrI71RogtOMZC6SZKp3OJi+S6FLdk5mCx8AzYfJDMuO8K+58EboNQQb
GJrDfUuUZvCXxvyYhqGYEewqdcsad3jN93odPm3az5k=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 19520)
MfgOluyWmoq9kLzMMpViv+T6iPaO7urCIvgxvzOxb38BthqWqgSfue/J5lzp1Qtg
GH4yUoJoxEfYGVZpsFm1c6PSWIgkTFn2Q9KfyL4NXNI80hCVZ39aAJ/YNbhXi9re
PdBLIh1A2cb4BelFZiP4rpJoZpb0yxd8Dn7dLrAAnaRa46SEME6BNVSoyfeNN8yu
P4IZzgWgB6NHdxNjusCYmtUrBJIetTeXlFcssTZwwehFws8XQtZ2SK46QjvbhBT7
f9/4wLPw/5t/Hi29VE7+NXVyZiwITIKleRTuJ3OZ2f8qM/b4PKB73ukWIDFTuwD1
p05NjUnul22NkqoF+FYiXS5brIJmhN7N10brhZiuGTLLuF7N2XO5p6j7uElYWZmS
TfrCG/qWOaRFSb6MK56Ar4Lcsi2mfkdUsdxM/a2SuVcp6TwhLCVVd9GQP32psbrS
5DUeSVnEVL7BdEiPQXUgjn8bIuwjYHsojRrcG/+LPbtDLAVxrfg2zjs5xHVk2yzC
tCxzuVzCTjJc6QdBCKKxsJEgbuxlgSmkX+ZjDX+HQTwFhNDkbYxGDQr/I644M1e0
7auQ/AM+jgZ2SY4mOo/qERADhm1vp8o83BW1xZoUthWYqRMEyh9qRFnr4VSYi1yE
HWaTdrMRAe1VRORUxGbtA6b0cj+C8uNaseIeyGFWejz8jaZtR8S0XWeWnUGBJrmT
6iznuVvmNALpMNAgTQSmwkIEoFfyeQfqssXaJIppNC4VOYjCr+t/dLJaqkV9U7oC
taKVlJ4JC5mYKpt5QLyJhiOslg9UtuDu4UkqxMKLUNx7ZAygT4Dh8Fdlai2noaIa
BUEB20FCR5/K1iEVWm+m/io4tXq/1TRW19A2MPEA0Adg/kFY8B2BWFGM6AYI0RCr
1lWL355V6RpHlf6GZhNteF+blK8VZrxH0LZlfUliVPt/Oux8aYNt1J/BLlbMtCHw
zAPY2wla2jeWbo2xJ8ppUKTeCbBIruGxAFdqe+F6Fy58eo6u5/c6SnQszYpwpWVt
cz9j0V7jKNfjiA0AatyujRBzoKDPaOYqRw0tVdkSCPBtDwh63yp0yrEvsrk2sZ40
Y0pJJhMEqxoVaYTl+iaSpPYyT/n4qZ9uIWGQ56xddBbbEXCWkN42KpSbfiVb6yFe
upTtTE5Sdnt87xBHEUL5P5zy6EUSu1noBlkt4pHEWMOTJEUVKeYOJCq5o7/GGwDq
vSbPkIVipiZCQtK+tqRnI2Kp9HA4Ucblg1Bdr4Sc2eqsrOZeYXmOmonuuoVyncWi
JT1Nxzs0xeOwxbhD5cUoBtU5Oi5Rs3XUwQp/muZ5Ukp1sZ6PPRCOZPB6zrRnxkzY
LfW75qXNC24rASjgPtw9bsiacdsGelwcfFG/hUVlK0NMUB2llFfvtBCBzyp6kZyy
zfwzJjdeZ0eVzWM60ENgiU631h8ssFb/4XhGiit3NuXoi7Mycmt5TRuZ5ofWej22
X3KveOE35mhrOKmAZiExIHs4zu+m/xc7DM5w/TxszgmWIjlQrmykejq4/afMXS3E
1X2jfO1dKjAnSGX8ReLhDUvdbUP1i2AvDfvGqgb26UzFIKfuMck0qrat6E4Bv4CI
/TcI73RNwx3SbFQ+CrwVBDeUzupl/hbCCgBvwC9lg/jJHoXc5X4LVRzpQQ2Ek7f7
6O607ECpfxv2a8ezfBPYKDY4moiHpFxRe/xvnCgzHJ60qW+6m+vOOQ9JUIGjcxa6
5LyK5vQtwxKVmYvcjLxeesOb8JbHOHPmby18gUM/YDuTF6mig4y1BBrYzSukst9A
pCWb6yPJDxa1xbxkZm7XsHzvkeBQrEWBkwWtyRUZTrEbwmcaLDpFI91hTGRBHaNw
cGQYjxaH27Hau6Q8rwUxmdzvuxfodfA2SjSBdY0G4oFtj1rupitgwhEEbEvVat3Z
SvjlR8bZ1olUNDkViltagzQtilYHQJ0zD49r4pa6t7Ka3nn/FwSV96ta3yJEftKK
cwlRIBDMg61QQqqnZlpT43zRKvJbtpxCgM63uyDEk4S3cxv6r1y8O8XIU1/fdYIG
/iJ6AGIkBkgO1ThUd519mrvSwYA3euTvNQ5jl6BukHZ0P3bixA0smJHKIWa1lw5R
aVuh8XP26JNy4BhzSUr1OpNKZH3B+IZ2eGLDhFT4iKZEpCB0bdUL5nZ9BKdXB+4J
0jTnBHI9Z1UXMR0G1wNh3QW03D5tSFoCz8/1BDjWKnpE/QAlWLPnvxSKGNIlaPLu
bOlbZBLeoWNSZiGKA/W8Ixw3LV3Isr2OWRadXZuJhy9Uwown68x+d3YiPRERGNS3
3Di7MM9ErCwiH7/ZTx8QTqxDZ041PVkLPbqItyW5xTTUZSpkKvK9S2tTi6JkXgR5
hlSwiHZt/vdCABwnoQRNC67LN949JkqKerHUP1h+5T7rbn+wSsU7PUJVZ+v/Hcvv
1AOEWIbuKnzo1XbXZAW9dx8D5J5IyIqJLMXEr9ZRjMRW9x/Tbmn5lw7J8GMpiw4O
r8efDZ1gEfu80dAFVgcS2Tsh2JiNQUK6Zknuv1j+oDFn6hklSO9GyVRzOpUsRcTH
SSVNjhyiXRKMXw5nPrwP1hNb2je53zQnW+4NcrpNt0PA4mCDZHdtzDPXzAu/vXFq
SwrcH5908fTPXX78Tt7XV55VwQiJgL0sKXtufXpCwCY4lKawvLuwDzWcOi1f0vOV
HpPM8ix7sYqmWaLRd8HbQyEwpP+nQdJiCEvApTccuBC7tIbp44NqkWtaWGQmBcE7
SYQW6AyJLq4RraBmmsfUsAdhWvGE9tKWrklSWxYBMTojKm0fEF+w9u96AQRLtd5Y
Ag3FRt/03Dzj2fsl7IePWtRE8VUsG7pSK03JcNZlreR85wsqmrB7BvZsdoYaPo4X
tn67ueFFV1SqrmFTclTRUbSzsb5N13ogrVnkh/hB7+f5vLe+ZzD1nIeXHEykXlgb
gIMWDaovJESJwBuqEBGvowEefGF2DUKMBlEovyzdgg8bbhFzmw2BFvR6QHAfVvtl
r3vbl2PvlGGp9VetojC877YoAoAVgj+L9tFEzTOTaY22yHF8nnn8QQ2rKzCjVwMj
7bRA6iorVAg1xlZQS32ZZlmiu6dFLdyZONzgH5kUqPOGB2cw9NyMrNFP4umphx8n
IBKPc2bNYr+EVoq/WXzwA7lnLYoqdKIksRTGacTPoB27ACv7obCh18R/Gp8d73Cq
HuV0syfJOT36odZXGU9mQO9dHLBp2xEjh4dNJ4FElL1izBcTwgQy64sc7a6Kdrgo
FrTxqLasVd/BmBHEn1wpbQ220X0QkBLrehG+Gx5mgwbaI8ff3OUBuX8KSKKZgOnN
Wnrj5SGjNdfwJJnUoOEmzXYJdqvo59uaeSHb0Xu89622nRIqHKBWBhqEItY4J9xG
rPDf42o9o68kHGSWH6nIJaiNV35hznG7BoKrOvjDAbk2OEqgNMaj7Brme1xMoZkE
L1VowmD9kHymyQB/GRQAA2CHCY9Lh4emOQ5bfr4v5zfZmCzlZD8jEGM5Gwdk8PrO
zqFksc63z/tIT18xsqkM4ytdUEBZO7wG2gL6fguxfsVOHtC0tCkJtuWaDcijANMT
356tYMfJ9EFf5jKdFC5lN5ETPpcFEQyX2XrSLYCzi80+C82bYvv17m/PHg7uuGCg
DczqgSECk0xfTO4vgzUgeYAfi7t7coUqDHMYsu3KbptQI5PLAKijuVJgvQ37v3MS
K7RgNDY7JHdelZYHqyhbYAVr24lDVpD/noD3SHIWeKM0pC+RHB4D1mHl8D72Rg02
AA4SLupBVeV92Zt44UDwzdu39Izui5/ht/pAwQcnGAUZexpO7zEw0OZ7xh5Vv5BZ
KWLja5q/Slr7/vb4NALESmvGY+rz1pGasei/SyteYiXhm4VvBouwaRWKt60tKASt
9z7jQ2YR0NSD/KudoTaWgAyHy9P+T8p+R2/7+vb9KEjanogp4+SC2Zr3b6ILXkk0
hRIZ0+j2xM/N9R28NrKYIPiTbsETU1BQ+hhVjUwC0KaSWqD64VAUy/HAmTWv3uGz
VKo4A3jQG7CSISxZhUmiryONSyj6K+5TXc+ecZvoC0mOoMueH/tbcBrtgd4vt9YH
JveXmD2HeorxfA00Qn3EKnr2vDBr9IW2fnDa9pi6J94UGdPIAsD4r9/P36GIqGIR
JpmWrQbvMvTNVZKj+gg6e4WdM2H+bU63DRRy8O/aaOM7pHjbJe5OhkJoqaO9XCAo
0bYtQvQNEcIHhKgVeKWoK5umIdws7ZASAe9irCacm5zTe67KEBRldIV+Oiy4NPmj
OUtBNW5NFavRlUkfE4Y2i7Z3CkcHYaz6Wu85kY08Qc0Quhj5JrEYgjQMelDXJyZf
rqTk+Op2rBUFOZ5BFD9AccqntAhmpwcr97JUv3Bqbqw0a+dJedEnUsCsMQ9Gm95D
nONcOfMjvYAZUPLgkqd/Pucj5UR8HGwZIp7I4TDFfHL2zmJ8nHQYo7LypNwqORX/
8ExeV35p7R/05wP7A/5gQYss8Tc/12hQxYrdmTfTCUYpL+No4euZCpZ7uBvid8Y8
WVfBM/+MT1SROh+8+bc6GjU05qB+IHlRdpfODyv+fiKWYBxZsXp74SpKwSIvfU2n
Kgl8/AeOp3M2tCe8sLlxKfcPvMNkJ9gBWQ8iFeEO8PaBS77XwbB8WTJ+yOSzwNXm
xHgjlFiXfU39m8PmfxhTZzKyYf5h3P+nZOlcjwx0zR7wmCJjK6QXmdV6+6HKqV25
RZsSSTrlWpJdTnzj5QAB5Aux4qE+2tO1EKZ4eqjlthaQ/zkp7a/JLKXxz3iKBb3w
aiLaNhKc4msxxGb2jrl/ipEbZpAv5QDRpKpigipugDXhz/llEa74Zn/sNtu5z2ZY
ZcmXEQQpTABHyYptGYRvUph6cbZWXGPR5oyZD8VaKa5HEn5Q6w+S3PJbhejdVzuF
Rn1IjCmNTHpZFfDKPl28aRvbfj54FDB1M7S4mYv4xDJpJzA9RMwZJs4Wd6OAyECu
nG1J7FxQfz7+CZaO7TYg+sAbSHEsxt37DrCptjeMg5c2bc+mJDp0m2VTOXUGvMS9
5TiTlYFJm9gGpPp0BGiXt0i0b62k9yNi9anGIoL4ubHTVIv2ve1ou1O01jliply4
9YgbrdxE46E5+uhBE5XxB1oU+IdBneODI/BpkFRN0yRmocjQQVcXUTc3EBIACzFb
jK9nV3nYOvzzefx7xHLJFFJMmVIfTwV48R+uZ/WUGlZsn61msX2KWg/WSU62T9gQ
FIsIdBUelRfa9ZvQ2ZusGF3et1zwEXLBfcjkfDCa/aeTByKI8ceW+RGaI7U3yIg6
0oHbpBl0+vnQOb+TGh1aM9olntZW9HddKxWccfFqdnXJt61/zQRZuj8RGlDpctUZ
G+eSyJoOjB18pvnwjzVGAdTs9Vmc2tppswMTlfhJJ5ycVHDLvRMMxFCdiwx54Yi0
0xdYbnrOEuMXaarVlUiTHgkd1Yhxtosr69OxhBWjiXhaL3OjtVGugWSSHarz20yN
AwrxlvwNojVbtTSnEbjuXtnT0Bx7xY91u8CmdiI9rIO+4eKsrTiRK4jB01rvL8hN
JFB6NmSdteDP8vjRduK42Ox0dhxcm2RIYfg32QxrhMj1b5jSZ2eoKA7/x83ZIPdJ
eo1fZc2KKFFH05zEms66iHa+ID3ry9Dfzcty8gs8nPiwR+fgvq+COe7tuDX+OZYX
5OuRb9DINhmdGwq3vk/ZumOzjWk52wT9QraXFt0/qcSvGRQMpvn7CJdygwg/27d6
i6gYqHoh1vA9kxabB7xUKli93S/hC6gTsQqJ2nJRohkMIFMDc9xiDPCTfy42h8M5
f9zAPeVwP5VRbsHcug+EdHv6abaDV0/QDhGdvR+cpPMlkpJKsws07gq1docMMi/x
Kx4MjY9LSWLubNpAYKMy9b/PIdAY/KA+4LB6VpgbX7bcS+dN5AawfUAk0DOQzHwV
pVJwjxG0Kc7AlL3Xn71TmN2SLnxrbkiMYY7MFx8/OzswxXVt+hyMTlrbtrY36YAw
DadB+mM3fLI/hvQSthbxXsP43QO9vwxvTwOz0smSjB6gtbh2GrtBS4Ev/xNBIMD3
PiziH4GMeXS9dcpTO1haZuR3+lZGU8kZX47cSKnucbv9Ku1Oi1abNRVHcKprVElA
TSCBIh7jL0glLGr9fi3x3WBXJVfFJpJwIKzA+SalrtEomn0tGwK7jderFgm1xK+m
cWfWFHRaSRTj+acjwZp8Q7Xi+SXKVeCO4ih1GNwPtjKfpaQvSOaCz4VbSjXTWNPf
yRUPUTBZPF1922UPpyWOeHLeQADISdw/xiYujF1fXFpudpcgA8EI+5WCU8Tl8y4x
gRzqsZCNHq4KKZ6w7u9vJjTClyDkpLy3mnoRyRX/V20APTW9z7NUs0DFFeZ/BOPd
1S9vZNN4flVR2LY6JdC+wTxIeQMzH2AEFwiQaQmZ/t4gAq59w4LF/A1bCyqQSg9S
G3OVwoNp6jYnAt6tWom581TWpqy3toIsqNHWGs/JWxSS0RVk4APH4cbsX35OheGy
RSCy6APmw5ISwYfYxuUdmXEWQNZKzFVXgSPjz7jK9eW/IKkQ/gQgE0amYMEyjpHe
bwGzRrrU5s/biedCTC0iiG2E5tS6imDlvu7Vmw0PnCareMFXQ4dfgJDKPAGpP4EZ
ArP1GDoE5alLXypMVEoHonBV4pfGyQ9DsYcOI/RJNmzX8245zXsTYOcTr324ME1y
fm1Pyl8FdsOWJXL6RlyrouhcfRnmij6yEO256u3P37f0pCaqEbh3a/M8jUYQg+CY
QJSfcUofOEMjCWo79uHmjzGvHqXEJ21ersY8qWzrNEgqXxUegFIK6BpR1RUuXm1C
BPNhrWOzyVDRFf711CHFXc3qlXGWBdoripHKRjLqn6ph68Od/Exvzs7OfImLBw8M
J8YW+gHJVdlW4JxYbgOB5DIQ428Qoe31E5aQINL4ReS/SlBGEOf67aRRriU/sbme
+MNzKyI9JI7qmo1CMB7KCqE2m/cmxVA2rN60GXvy0cQB6eq440UfsOHffZfaofEH
XFXq9WAVFKzlO5AM27vbCmRYCcIP7aXk0YqN6FtrfZYOuHGYrXpkfc+mYRHgQ736
3xBYF6NQHOB6nw0GkhfAvhHd5N1FVLUHC+Idgc/GmmTiZf9oTViZyctSVRD1qa0U
Ho0K+R8l3zeGw6qM0hzdvWnC5a9nClRUXurQArPedmwXOiBgGY+So6GolzjbioQf
e8nAkLyZMyOQn/efnTdkBd/cri/Ku2rIOcudebqy/o2nJSA5zVdZjo/tsy8ByWT1
C0LGMk+MSH9o2EYAnkGc0PNG3p0C+gKwJ7RjDm0/MAsjpX49bRWYNSpcD4RwfV/a
9nbCl6tkNtO9dLgHz4YAHlvpLOMmcq7+6ERNgnWg+rBJDzGi0HLeoFdCgId/QNQk
edCAEeHWGOUgon0ywEymlEC4fQHTBoN3H9VxDjfKsdEoreCX/oSs/SwuuyWYw7n7
4dJGbngUPGrjfn1Vg6xCe/Z1ngOFQC5nhj6SLLTV0x8m4brafLdFFoDYCB4RK7+B
D4bFVfYcy13BAdZAY1seRPbPUcXlv3s3z2wyR10vnlCTUDIRp6EAZss98jeylKSB
bHQZgVgQMvaoprWobbYCdOk4RPfUAOZSUCKQKQ3oO9Y/8alNv757+g4cu+pYkY7e
OxGxbz4h88+BKw3rEdJCoovr2wmVH0DKWG/bJuv0cv4uDM+lXRU28utbRh+ZwcZa
pUH7AfpCFhVPO0zsHWdNKn0/aiOtsdN+N5DcNblRSGf97ymfmqQEL8XzjHuIzaf3
EFK8Dw3te6uX7Zt0ZQvS9wa+oAHCxamVpaxpuuUD9OVStd2JpdOIAcOaYe+pGgYP
ztphXymRzMUlQJ+qCnwc2y5VF1Uw/A2jqFhFEnjnn/NT0xDeOc4gKQHwpbQjp71W
3OtEml2R416qaRTOBIJ5n3lnzfRm8/ZfyD7VBxnmFJNCojV85mbg+Ys8/k/tUV6o
njD1DdssdMQ0+H3ZeXCdJsAoz1MtZIKwux4gVHxFHMz8H1Gsy73jYbui6V9f283C
zbIR/GAR1BzOgzIRN8aWOtiU/ArcV0gpAL0EN0Ww4p1/CJ2+Ktjg1T3eAI5C1/KD
B/h4aADw4oXlZkYKfKByrQj1s+RzLDELLjRm1VqXUsNlkH7W9QHNwlYmEKVzQhGh
SaOSugOM72cLGKAPXpErbSuO49G1PyT3JQTEoqXd/5OK1qiHWrbIEKjLpwZ2ZIqs
D9dGb7zY2HYx00PcYbJaQl0Itp3iOgl/nIqZCIMM+k6QLpF9ZYEaikNgXKvimYtI
zSlbMdXee2GvRkSgpzm1EytEUTgtTFVMrflkcLmwRFhaqZ9uE8lhDQ6KXuvkRry+
dyVHzs/b59FAaSxyya0Taq9DDrcnOr8RODixvA3wr465p0JSOD86hh6kvkp23uxE
be0r0janrTT/Jek5pkq06cITRsRq74GqnCZR07rzJC5E1z44YAU2mrcIbmQVNpea
AdNJvGhKlG2vofOG6NTLUIk6NABKlvhqc9DJIjsoA2xaycKnHoKYiM1oaIVNp7J1
j9mBYJyw4ySOqVCTMijkvOJK3+HgJ8mnDy8KGThgFXmujlSIbE6a3v6B/MLsoaiZ
tXT76t6CgeuWH29XRu3wsizSUy5qam4WVvemgBOGnMp64KGeue2/SxzN7s9zvkh9
mF1xActKhQBcWifxlO0UhAbE/efl3atXUb2Kif/OtHlFXdzc9Rz4vjJ+6nBmOuw0
1AgAagf4xS2JwHXn0xDHHm0FGNDUlLuL4ofVvUFaifZzdGq4dMDKHSbDg1y0y4L5
FmItlemBfBYApzg+v7g4F6KGnlCn0KK5P8Ot4iS+9saLO/DDk8eqzVjAMPzJm4aB
NuTDCU4DKTwFz+s2WbizSm7Vuo0MzEFs0UvPeOOMCr1EelMVDYpCWEY3AjvqilDG
2tAwkuxLEIr3eRs6p7jNSk9Ycpk2WZeb36Rc43lCXIcLm5OQnaLGmUwz0fk82knO
tNxd0fdbMPLeS8nyjpFTPtemS0KLVFwtRQjSrJUJrYYTECJx7RWywMBo+dn8jLO+
uGL6EqiahsOzC529PZinmaPSDU6oH0Oq8eAT2IbBEnWewtwHjGkEqLQrzDP05/eF
hcjwI7IIbFbGFwzDmgeyO7uugX7JpXTaYhrXTLp0Y9DlnbzYPeD/+11Bl6FdGno6
o/LxsQ0lP2DMBHW9BeMSdeWIxCC1cI6LbzTQ2OPe/znr6EC+aXoFs5DLhFyE5dFj
eauxld6+gF7lvtcPymChDsw92owkgKQZYHj0YGovCjWzGiykIM1+DLB3PXI0dx1l
zDh8Mo922OLMARLS6ANl2+Gh6MY/BFNs9YKbg3TBByTXh61/RPoVCX82F+hnKZMG
Xm1bhmNMedCx66dbfFXZfCocJ1UENgnYEQsnJNtKeUIlLsbM6xSH+wbgaT0A1zbI
MSMjTpS+ZMMdpi8dObOBTkuj5XokoTSTmJxLIEvXnsjpDvlb230TGfszvJ2iPrb+
0/hn1rxZGZ1Ueuji+BZRJyVATCZqAuk52PqGAf7XUEelefi/puexg6Zhmo66R7t2
CSr/0q3slyLSbdnaGq3vNjmEJ1gTQjQ8Pg/d//PFCVnyIojKM9BW0aVh9pf5VEqH
AsHVaailpAMY57pCePHeUk9CZiJLbIU4clXracDb14l/JHRfDMxoj3NySqJqVo6R
5tHCFlMoLeUWGOPdZeTkVJlMUP29FtmPvrK0hiR9Nbo5ZJ9aITxDJV4M30h1bknh
k/NYR8MU8zEblgBz7kUvW7ekh4xYD8N+QV4zeDB9IvzW+j+8ttVOlWyLkehaMCiS
Z2bkNoUmPl0aIehsEJ1KIS3zdEpYlVnuGlz5U7PseMh/N98ooTZ+eJiNGjdmhcO7
f4V91nHTunV71HkzONv67lInzdHJlG3Ej9Zbvmw+taI7OX3ZK4Pem+DM0gsA9qwg
p8yDokhh21ivBC9v8sbvbfHskGBPThYEwh6cFjJm34Uqz7B18ZqQlZG2/fB/PiyR
onohY7sHXfFpMEKuCN/KUSo9aNtmBHnyPr0R70GrGoHNIPM+n508wFw1cNdQL2eR
/EGgtV5QUX2WwcMBFqDFh++nUVgAQA1CF2Fl1CNjKRaA/sjr90pNFK4221p9NMgg
cmD49tTqE8o+ZSBslTsi5DHGIRYBq+i188t9t2kdYmdtkfPk8ljoyFXRrkB/+Kaa
kHx2TwzOIMj+sfGpcWHeo5zk4JhrjHrPyme6lOMUjIRMnR52zgw0mmlGrILfQ1sO
YG8uTpctJBmOJNolO0IKbJOETyAypyJkumlpD8k95XBYZJTNKjzNAbltEqlrV2VG
Lnd1qOgUkcFgrHK2N/l6u1Ac+idLksnEGiO3JKcLvePMO+FXFmucksZdLoEvbab3
RIpbWSesJeDMvW0ZpiRXcBeuD9R3cfl2SOv0yoJj/svjy60EQOTeT6LZyGLQEEmz
pB+oxFkneIhlmD4wR2TQDtIwOSRezl4gr/jIYbB+A16+NVpNdiY6W+H748egD830
5ICLv9KnXFFtow5aItkd+Cew5PdBzF5s10SM+IA44zAiN67Bmmqzy0ZTnNMAuNny
YpbNYh/sB0odaEctlxhFUGQ97G0rXkf00KdxWFiUEDfjqlkupM+bvEYTM89g7CUq
51bkAyxjkqXG7ECIxyMP4vruAkE9LwhHx+U8+wif8wgxA9nZyFQm3voPUzoBy/sK
OdBffS/hk+0+EdrI3yj2hjdXIGlt2cdEV3nT5pYsaQfKbz5DGNCJTVcc4aHP/WRL
0hiLKEQqj+m77WndOY6NvkDEnXBwV1XRm1zeCiHBHvx9vOYNh3r/MMIyIRC/AyL1
3y7gH3ZT33hWamQ2vhwK9xPGYuyzhaccCLTa7763gRvAIbWB6HiL4MT3wCz8K8/2
d+1Ut2aYcz42/uSQAIl+PTPgcRJ/Zt8cU6JSX83pE+qyeOoL3TOlkJ5AiNLRV62J
uzgfq38UhM/IK1ErsstFPIf+hKtji/BAGBCMuCDYaosmRQOHM/TQR2zOrPljZxfa
nb5UvabM1m2o70xZjemRFtXsiQBOnvGQ0eOrk9lfTE127wNLNmM+yF+MHfIi3e8K
m3cWk5/5wm26gQFX2ps96Z3FJrkv6kBS31+xQIQrhH8h3/QXQgjwdDd6uUVoaLOU
euAM/k8CilE4BZ/+AZ9K/Bc0BkzD8vHSA8pJd56UMF+ZVInfN1qqB6Yp+L1tv5gh
TSNCCdtQDh4WPRrDuB6owKJhXTzKz0mMRrZUQKXZ8biQuu11XaOeT/uVvfqDRnh/
+eEaNGL8vBAswtHaCLf1NiK+Zj4LFvh3Rb2RTQg48nAasKwZB10G+FxaYXdLV236
bCgtlbuqudhLKosO47AguIQA2dtuAT77QeArCB0Jp9hCaFtKa0EI5uTIEIuDqK9o
2hG+93VhPwcjd/SidcjHqQs9kla90G5u+vcc5Mm/rB7Yzau1ipjCeRWwzd9EsN0b
TXt044b68zmqxVv17IS9/r61usK0jQBY02CRMiOGuPB4L1nH0l4wNvRKfd2sQYC8
zNKz4Shl7fj+OSzmXH+gag6oegYfXj5XUgAcoeNh6OipaeCquzhrF/0oRHr8JzeW
hDCECJfLmxT1eMXT5i5l3LkKbHSwmIajsJI36BHb4QMidKlUtR+p5uTmQogCBvVK
wOM+Tlqo88Bl8cmGrlBnv5QlyB1y0ovoIpd2kz51gdBtLkdr8Si8hs99X+ygImpD
sPNs6m4VhS+4Ll4G+iXk7uHc7vOafSJTjqnL4n6MoXwx5o3RU3bCnGvnfJ/gs4Kb
m6jkrVMEjjQG6PwQlIaAacygqVh9zqem9NaKFSwRLk3aipmPwaQjRP4iIhIFoRVr
Jpnjm4l8uUkftCrmRiZQnuHlC3yJdm8qUngBnVLSV+TYduZrgzEF/16zSSsttXND
nrdFfkljkQdDjjBC/DqD4AYOcV8H+l62Cdcmp7rn6meIZTad0qoomAPSZxH1UEJB
CP6yZtuvVEPRGyuntvTs0Zk88QDw+6ISSyuh0IgUblgNrdEu9siuN02d7WAY1tqA
CMccEeLUC9W2GdBXz0W5PBVE1Ahb+WHbtygxkZvwfGtHiS96nWKHFRiHq2wq1tXR
hQaK769LT2GrxHpuZQc7DdOyfP30Fp+GMF8jrU3QWtQSrxHYvS8hIiGT6guTg0Qq
XVsE9l68qkseJPdskGDAkOgXVi9HXphhVGfZ/9aKkmaSHBqhjhdCu5L1yXXDHdAB
jm6GQM6xKupW63qZTXeoWzsGk+KsBmDu/VwQEThPITLOiTRPm6db6veeZ+q02xy7
Ijo9EG380eDWxEI3ynSkr6/hD4LZDxd1ABFG4hQzB3xqMJem08tGHEVFJPfihHk+
mpC2SQY47Hr32ag19aRpDfd6O7E86L1G+irSRfMraTuRhZBYN3cNLh+Gr1sz4qLr
nTsElaykUiv03LiTmYK7iKoApLR/ICBdw8fPZg1RAhyYbLiqoaZhRu91VrnwG6PZ
zsTBX90c59+SQV3yo0yI2MY6yZywfzRVt1Yp40FyFLd5e2D3rHUf6a+ZBmULPLRN
EC04U8PNgDOKvItb1o5idJs25/6JaScDldpwZ/Oeaoy7WE9qaZVox166LrLxm8xF
a5YAa//tLDXGgSEZgaxCLLM6TH7Jo8iwFZd37mXxiTyCxxnR539M9biDQMAqHGR+
JcJQi0JUBaLM4H5zrtg3t18qC8hmDGlz+HqkaoCx1O+pRSPpo7TW7xDGCi5xml0B
ClgVQsUG/FEremzZDZMeioddKn7dg93L7cmdjjYJM2XptdzknRskfHXEYMXcS6XS
QQFO0V0HVxwNh44hJWe7ybAMAGlTNRxVXroHoqmMw5as0Kf/D3Vh+F5F+695GK9b
ft/4gHdrAh8QkT0SFB5EFbCaCpOi9D5f/qn0AQlcHHmN1l+in8c/9m1mSfmSVSa4
81O1mDuwXs5Sl0wlTm5XVSiIwOOm1Aak3FXjBuDa/RNMHwYmIr/PnzCt0AfwkdGt
Hg2JNvSLn2v+kf9loiavohwxZ6d/1/PGAJdHvTM6VedGkl2TbusQwUAmAJMHjsdg
TQ+xv8xd2xXxNYu0QF3F4d2D2D0ywZIScxLkEXVRAy2z4ah+nVeEhDQvLKxuu5dR
sHGw9QkfbXAO4lym2ITuEYPCM83TJW22vVVKlnVymBWkm38fP1DfqYhoDpb/V/FV
i7Qdure9B/Cf9Xhhd6DlBcksTGmJsHurRVvVqRW/rDOaBUb2fi9Hi6PyjM3BimIk
KFXzM1+Cok55t1LAarOM4XEFi+H3k3JsX9sqP5zPj9RbD1q2/u28y3TYw6rtwhAA
o5J3JddIWl9aeSVvrejajyHQK3PrgRh/tbIEIHsJJA9ZDAX0VxLli+5KzX/zwd/A
h7Rb5xItg/jjz1K6uCb7qDuylIKd7PwPW6fH/CYPSGToph0riIXIbO2L2yQ6jj7F
9zwUTmOO8lyMpXE7j7/SUhiAe/c+hTp7TMRNw/NiMtodtVf6d+jzoq7i2lb5dw9N
Xeon/PbS3yCxrTw3W4JhkNMpTMJ05RPcqErdJi/CHmzcNSrCiYtTmkXCrWgd6y+M
4XFAaMHzhW5epasWMHIxWW+NBTuVvawPyLf0g8NFqgK2XzClMCaYb0WeFPCnQj2N
fY0MD3Xx0asSADtUWlqtJYP9bZuTQa0HvqKSlKTr4KuWrchOZtQWMQpAo5/fW3oS
tqjGaq3ZnBferVr9Sbx/Yhv3W4guv9vsiDZvqOYzqHii0/RD/a03VaPI4huhzwUc
nmcoibewYazMvke7bGUUcXACeBG4UJKpU05NtY7jRktJLuNAu/OzoE4VF56BBjSZ
Bd4+4dlE27sPqPFKBOHsZrOkHrSKWHLNk9t4TXpPIY3WZcY+Xb+44mCSPj97NVSX
XDxj3xYZvQDQh/4x+CUBj8r7Kfk3nZczUcdD3tlelh4zGveUHt4eQeQdzHvnOC8X
iEZOgGWhBrUXhBechC8R6OmCZ5PQcOF6jnkrUkw0UHoP8iQyKhi1T9Dr2f6s8qWh
cEQEQaBqok+vEq9Pf9kJjDeR1owyjyqvlaqVpWEyxbFOvtXIgJXj3+qamV9cjd8Q
A7RPuUWqbxI05w+Clpg0TlBX2LZ3T276aG//DhBik6WPtr4IuRUsEfkRp608dPUS
XDb9y9t7vIzta9wMOprH4L/hRe3BmIQB07xP5dkrJCsEFdwNyRUnoKP8p6UKqP/R
Lbv24VdCKY0gmA6hZYe074owZfNtzaboyUGyob5j+ePo+qCzBcvLWuJzNUukKxRR
GkaR0s5f4Dkfvjc+tOCqxMASeF0ShFFo9hXhm/fl8m45QRy9FKjfV/VJ94KLPZDg
2kteJQ+5wFuwKtUrPjUbYxIiWsc3uk7/4kIa3TNYq275t2cXdZldCypT3OE61Mv8
KW5vYzg0Po3Bppy2WPBAzpat6dbVCaVjW3xmuNvkr2Uw9ybSsvdJk1gVI23b+Rbh
otu/aSJNAbA+InYPw/Ou8tZZLZHQfeO9XSDwQGdSoNIfVbqQvoC8SPU+u6XKgWug
mIBHzXFkd4cu+uk1hHG3Y/m6sKjp8zfDgKXFCdN+Rts/X32oDCnDYCY8gG+JmOhh
nSuXfaHx/NdnavgRcXptYN2azW8mrXxMqNFKuSt1/5VA1QSp33M6tgKSb5YfHn9C
+rEhCDBcLPMLYOHiZAj5ToZcakWG00u5xXpmJ8xfyrLFp19v33MUK3EftuwRAn6z
Ndknsl1BncQVH0Su0YGfOp2Gilorcilclu4aPuhEGEOXy4tBU9uu5tb6J/nmZQmL
WPVRB1JFdbMtGA9P1bJejE/QOgdGNyd4qpo7Nx2tc20h8tZOQfZBOS4eHYlb2iOg
pwLnRcD8HXp9mb8rsIXS6ugbGgq2P6iKGWYcJ+a7+Xq400RF3opL3ix4sWHLMddt
qC7FGX+uh5FMgQasVN1Gd4OeRRWWs/f2WpVnOsjbFweh4QXXRahTz6+SNNtKEk0j
TzNmn/LYy5mQtzNYBFNBqHt9Mmf75p0cFIB3C8M7M/M1A5gs3/rAiP/wyE2C1sBx
uGAy0m//dwCRBH1tmcU79vdIaHyoof5NjG01uD8ATzMK7trURyvgRm4yG4bYWDK/
x2NOvLemj/1rsiFKp96GjkXNbmtJNxGCFV2XmSEXURXh4ufv3GPsfmhmhys6CP54
VTvTY9HL2nJH/LgRVi7GFVp6vrJtqkMddrdIo64Yf+502zQ8hvwLDI8Mz4yN6dQN
uYVgwKu7ffsmGl5tsJR+MZNcO1ph0WmjwhsbwhI1Dmad7+lTiMDyYNlwNbj+QO3i
FnxnwvtjrLZc+NvDulKgaHPbmOsWQa1whrT5eDHyAgHyLzAcfZIBBBbsSFR5xaH6
UIk7UE3onrcMd5QdnKfxQ255m2AOxJ/G5A8zCSE6VXD4hKAzDDKcMb9A6l2kkLGB
cSNt4/7C0oNrLyo5NWK7EuoDR4MhPuy9J4BbdHnVNAAwOh12mkMbfE5QLM3I+xSh
8yPG4uhVB0KpqgeX5ayjCeT6mNqivx5ByQWXWCnWZeg/mK8of9Eu422i25/NkXSE
OCC+nwS63Q7IWM02C6Io/7+8v9TPDrrtGYhoe7lTIa9Fhtg9ogMoE7kdaQDZcOri
naS+Z8DpT6M6Vx0kWmVRO2erUFh984rzMYiIeICsIRIhyPFLMV/81v8qSa1+e34G
9LCcA+0TAPm2fHqAdkfnJnOM71DxqoA/W4sIavOE4HxNiPLoDU6XddT9CZQUWUAA
5Jr8hXlKtLB9qf2Zg9UgC4Q9ZPpganEPuqknNE2bwHNxgF2dS+xEHwFm/ZBHLQUq
eTkl9TG5xdNVcn+sqKHmUHETLaOgqaPe4uu9iEA3A6pNQIsgtzmbXnNiUiE+Agn6
URZv7UdoQT/4ETTjU+35c8Bn8azkZygKiTWyV1fDJDBMIbCbh+4hmyFxgyzPPYT6
3t8wVwGZP+vHo4du6VBTAUcOCGPrlzHOrtt4Q4j4EziBc1wsYutqysuBty77EP5s
LNs6MqVLKE3h9BKYQ/6Kj7BYvQMae91GGP4D4XQIRhu1FfXmw6EkaQDwh9pGRk+G
v2LR8L65XyfVzPUnawAFYJCIFSnNv5PQOE25HqpsVQQw80rTwLnwuHV9LoglejBl
QxdNs3N9jA7J8VYOUF7GRLM1UwpHL0a0630CTyoJKpuSdBfLGjEOysB7ddcTumf8
qbRO9vejaJCA69lYmo4vxsqYc9fX+Ankvz5yIIm7g/ze9+NcW14NGy9zbG+OkrST
7Ovzuv2P7UqLv06u60Z4wb/NoCQx/cL3P1mh8+cBKWvPCA0WQxquCqWubU2yiRYf
xfghl1Fz4UwcHV1Fn3r7osx/B98Yrp7Qess17zKTjywwJpv1hwsfPHGNe/lxqZiP
m4+rAO/eXYxKIV9gfd0A8/sZlY/Yd1kAHVSy8hBx6bpifjbONiX9OKQSjg3Jz2tf
yqPqNVaXSvrS2PQxx9lOkBP406deFS2+1l0Djz2/r95unBObqF/X15wPpABQ5hpj
rIg/s5UffF68q54SIEHdYOlVDMtXeNsxXBnavFxyJi1O8hPBNSr+/dnVg+IOQgnC
0VYFOHrtcxcUkt40jDwhUpT6eiVMoODe0owJzZfctr1yAejQ+uhnLpw4N/bXn8xL
ffvvfNFfSoSZ7nv7QnCC8hdklDqNOotSC/lHhzLLBJVt+bXLeqErbV93BfIPx6EY
B69ccs0JEaXuXie9JglbARPqfTTmmer4M9Ipo2jlZXdAsq6rNToNjK7/IWiaOPlg
kPuukWz6t61zBVUs+PpBgELn2qceb1qWS6qMOW+5aJ/tPMDZzqXD5Ak+3f/9dWN2
KfsiswEkoBBKbCUTepZv/sjSEz54mxGmrKZumL8flsIjBpE8mJTIzwKKkRVolY0e
oKrrJqGHicPO6iktFh+3QsiGblEiQ25/7xOkWpmXsxPAAwh2srkDEQ7pLHclWVHb
W82vGQknCc3oWc24ON4suRnjSWtM257tm9dng7Y/Lr2U7lmgTb+SOyxgh/bO0oBg
wAHeBMzze2u6KD1DYlKvLCbE2EEeBzhG0WZDJ8R+b7tnfxJFTYrzMGk8SQPXHaOb
S+gvCGtWIYGVbAX/9dSoO7/A7jsC/RVCZKN5oNmIBt2YlwxQezhyGylMsadTSXuQ
Wf1DGppcyj7dFPc/BAYgOqGXmCoNJLL+mjkZJ+akk/T0I+SdUbVj6pRywPjACUpB
zEu00CTNUALAHfDMFCbM0yagSXq0LhAKjY3K8RYBS820p+mT8UzOQEmKA9hQHjP7
cYbv6Vo4L6w3Mbtr1Vzc7+VLs5vzArpihCWqhIQfhzFZyMqLlG0zqRbdVnOVphUj
uyn88y9ySyQEs2kDwO0PkjXxGuQgiOtAtgTKPcHtK/2GsnefhNFwgvx9ymeGU9du
JtGXTjZAu8vvA8utiyy0ulshq+Oj36MkOPiyaFd65C38ONJVOnkf7A6fik6evNOe
oXWav8iLlFDQqFF9/1jeMhTl6IoYkrkeMve9qSlmJvVyoDTKwsCJ/CWGvnpAQtm8
KNs+7BrWxOkFNp+KL/40HZ4ZW5ZbddxF3AYWQ6JpGQGvItC2Q3bou02zD0vXqarG
gpKD6EdKHuk9ZlZSz0myF+JEBGCGFUgFG2bNJwPK8IoNBa2Rwe4l/ItKK3L/YVO1
Tjye38R/wwcp7jBzgsMrQzWZR4vMlKRCkQckmejuVL4+nOFrxmf3nopXNReGglts
1I72w/I1pgeqrvscpzfYUwfg6nie1AX3009NHJEvbUvM++BX8Nkbe02tbHSsSpQx
esVDTisYKD/oebLhfQzyUDdCe9c4eu4pBXwR6AukJddlmxbhKhP3pBfftDZWqC0t
zdWS244ijeDn0EQXP8VS8zF9Tx28tlrXgdhAr+To4VXU7EsLSmXzpANojr/XyyvS
bnn/VLni5ZWg3suFuQoHCbgOOAtYAHcsVTEoL4v7WpGMqG/IcU2f12edvwcJP+OB
oKqOSHzSkxGC33b77gYN6igCdgZmfJuUclg4JSqxcX+E60IZYTvlGi0CSU7ROaqn
kgxGS7GiX/aq4WNhcyNMDLmo9PHhujoU9htl3Xz6eho13ZzGBhLBr5NrnWu7a8c9
I85ei0sx9B20z4ZyN1YNyvJT2GS19Wc6Z5QrW0LhKg/Mfqv1MS0w++OKhcmqxyhq
sIKZ97WvUTlUxOSv43WQ/XaBtX9pdowfofLwTH02cieiP4m1XzNhoSMN31iHYNE2
yobr4Y8IBsmrLdiJgKn5PA6Ymo1WIfFjlQot9CvUYC9oBxGesY/bHV50uLAz00HR
WfmjzOhVT+iLcBq+a/3fl4kmgZBidvD6PSjgMekHYV55u3rgJTIqACLNBf1us4NK
//n9utX5VwOa+ZL+/70k/c1dMSbxvxIpyWO+U3+lKkaD1tCdcSEn/gmnqM0+q0or
EeiWJS2jm1LD8mZjpBKLla+fUD7sdoFpNHmm7oYk78m38rzKDruyZxwe4V6fsOW5
WRG2M1c5fNm+HfpbWT7nUwvhXxvsNyp7P6VNXFJHDNJcWJOE+8I4ZoDAZWNVjVP0
njOe3rqUQQFP9ZUpvew4IsJZH0VvBrylCg5PlC9TC7ThTs2PVxPg0Fo1mtrePtY6
3emXO9EXrex2EH8Bcyp84ZONxea7TUcNHGhwu499TJUSdkoMfWjEyyeyCX20cKd3
R0feoJupPOPlsuEcCgefV8QZ3tShhDQasRhZXMaybhPzbPaY6ajcYePdnMLhZU8V
j7ZdKSqIDbNAmJaKpYDgS52Okq9LJIXyL8DXD3KsXFy9NqK0B1u71qbD/JJFm5c7
V9Go+tzlUt3csb/qzyE8aJM6slC7KejARYhyd7QNWZ3r+MUu+E42PeFcfoXvYumk
XS/Z5ZeZFw+dnwouUO2uOq7i9E0v4mslVJwOEr/7bQx4pH0FUXeKgODNRkhXwt48
zHmNHMZnMWwosiNPg9QP0IsYWCWNvIPaVrWnIA/sa8xusG84hefcxlmJaO4rafQI
/mFlsJ36JDd32RHN0iaFXyumum/pTFnX9uLlKDQp7bdG0cxlH3Oi9O9fLMuRUP/i
A1NccCsGC8aA61l9JMIdObvSDdr+cDi9kg/aHIaD8lsU4C+GDbknQ73O+IVwSXLc
5HN6Vo/VsN1UAT5uFIlTTG28E6zWluFOYTLUtJRUrbHDuMl6B1xUMGbdC+2M5cn0
S5zyLwJDqa+vlT3C/7z3Y55bT3iZbQiqYrOpqWdWOvoYIKOfCgXqtKMpYjsU4BSE
LvqKJICtySxzy+monvGPVmfvqp1gegTREwFQ6QS3opANEXdMaTycwqlVWR1fycrU
u9Rs1HqJMuH1vo5Tr8M0JT72hOtpbxDgmqnBQM1kg0PCoUZAPGvBmHONNErWAFJh
egMZYLCw0W0cWtNuO4FV9SM7KeRiahN7m+F9N8j2wHYChs8MUj7hDy0mPp7oH0GY
KZptGvIvqblZ/xkpAFSfVrdgyOLFwQnufXs4MGq94w8TGMwgdEhYLtou+Vf8ifsP
HpVMMj++XukIyMOUStxUERIXowNXK2+Xxjej7dIaNrG62pT7FsEqnDKg24+mwYF+
7a4SHeRRN10KV2kmiZhEve7ckQw0L+X19xtFE3biIsi8pEhV6SYs//SpNRzypslr
78/aDyfBQa9Hb/pOdt/dYL9nhCJApdUkeS+yulyQdVyzKKwJPoUZNWI/IZgPgElJ
X2KqAnRm5qM6nQQi6/Jpb+kTEemwXNP9IFu4hHNXkuNbQ1I6p1jq9+HUSmGgQU4X
LDuRoADPgRla4s03BRJyibdWAZYU2ekAsAaa/pFPg4LDQk97xx1nUQGpxGSN4UGC
B+zpWn1dIPMbu5ik+NaGCncmekH5d5u9d6BarPp09bOJ2QnjC6gKzb4Qy5TbZGlG
j534vwueQNn3gcDJW0/oAmRpmaEvdL1J0ZAKd4YljSnmLx64foGBPd0sMcNyuDEH
Qr4SmZmjU+kPO+HL/CTG9h1NF8XSnQJpZ/hOnrQxmJDoU8Xwd6pRQv8L8pOR1ym5
swHttPqVsm2GX+634yodepMRKcz9Kw6SGwDvK4DeXPZvQxqTD1sqOoOjU34VA8Lm
pBlCEgZvcKfTL85teW5nPm1xxkGnXzWY3yJFjb/b7NFPXUrMFUI3n2N9FBUKquBo
/SEjsd00HWIV9Fa2tHRxhA2adcc4uZ+oH2RFGb9A7DYrBUN89/4ECT4WMBoopO6y
CpmjzWQStgXhdimnZ+whdvvCqsK9zmjW4I7VxeIOlkTNpyNK9OhU1OAsoQRTYngD
oQ09I3qg3Lyd1tUPf4GAcyvX5IEftEJpQi8dAwNKE04/yMQBQR/sNjibWzXsDFCT
yJHUOJQ1AoXsfZ7yS8Zb6+esiLT+jIjBXZAQpXM5wG+ReMPM28drdHbgydmjOBsg
qkW8S791+ZjZIdNyhNBoghNh1yytqDF9xPgri+w+JuOm7zL6tv89ZpAMym3Le0+Y
/Jhy2ZrkhuxkhF41l1dhVSmKA93sXvYxCj3PDTcgLAAnmVovBalj/zJbb+JfEayM
5CuYX0I+FwJ+O7OMeg9sYfumvhziYFLXGKXTALvUyFRRthlyhqKXvRb/Ilcx7RwQ
gFUzHM28a6Xgi3KAH8zyIE85IJlTCgwuNS1qDAcGSDj2mA5rNlktkxPUjKPEcnug
VVFmsZSGJajnjwQkxbNDL7U9ogeacGhKzT+kbpHD+Rr07rquzLZi/M8EbeYCtH1S
p5880D/lw6GXFsUqCuMj5YFcNohO6UlUBR35BAkOZzN+7taqpE3diHU2mXDZux6J
djn5Djh1qT8KbABI7Nypn18bdA4jANeN34iMTsYj0kEeflbP760txRhLww0h/5be
QKk1r7fyk5piVFB1Gd+/mJ6I8OP5dEdXESzDeTMGmVcHvflvm2ie3hUj45nL2RCg
pk56anfJvSe8ndMTYuTPn/JGVmcvPMUbrVVU0GyPNnZHRZspDYDY5B2NAAFXbMZn
C/J32wRVZWhD4UJi7gENW8M0jpUX800jDblZM+06w/FPM/P2MXOav6W0TSmB98nw
Di8KEtqjz8S+KxAeOjwRTBRIt1berKLvZGsbVv6I2xKpWaQRcZyA09E+Jemm9coO
zTo3y50g2Uv5ZU1bmIwvqmhQhgoanRg+CaO6HFtSfCxDrXfKQTXLqpHQQo3fZ+h5
cpTaDmVMKN+Pq/vtN2adXek16VATd42H5XwEPTXutog7c4w00k86mEmmQOsX/40U
4I+gl7w+T3DcVFAokbG2uPhCq622GXyrIRRfJ63OjiJDFkS/Gx5EN8Fvb/GlGXj0
/1CpfeIrGyT72krgOEG52noqynRZtBN0ij0Re5JGbQVnsiEjJgFh2hHp0p9ShNU9
x/8ACG0WAA0cBalLesbZM78s74+2Hz3k/z9eSBhI/tJlGcUKbFeG5Sco9gHj4ELO
nt5nU1D+KmR2aIaTLShGXB8/lFuJVWZ/t1tGF4jci/qp/qrZQnUQefpRBdcqqlJj
6hKQRHkpzDLuULSnc5OqowYrDB9yiXnPhw14JzqvUYlPLfLsqw0pavc24xVvYNBd
2IWBY1z8i7S84xGWaFUwFCYJ+yQ4ecVp7nTQb9fH+gSOzhM96QT+3rL4gd1dh6Iz
3RwxJmtmO1rz2bqlQzScTUAR8xvrOteLkzVSCoqteBhGR9sEL8TuJ6mcRYctpduT
s2M5C5rE0nS9uHRmGl0ElYzD/w1jEkpnPihKqIEer6d2AFj9jwb+svVyIipKEcwK
DkkbmxUKH81FS5KoTTduRqgTpQuvsUdcjwel/MgaimwQC4Me+amauNyaEGsV5Nj1
eMGfptppGBOeYbVi5AoyD0nu96sFahtjnUOFFOc0ouJDS0lBwgLH26oKkQ8sYJEf
Z760q5AqipDLH5WCwp2YPojvTSN6NsRDPNfTSFDnCK+nDiZg0/himX/SIOrDZwrg
WJ5Qke+RwyvQwx6KVRkVbfWN7yi8QEHMT9BPKSasvyuVHUqfeEXMWyLFqBik5Ems
g5xBMl0pAxc7HElRsrAPtokPhfGaWUNJsAnWNO4oDe7j4ARXwPBziQWsaypCHkkt
RzSUau5lqOLhDlU6rpAUOP9eCZeMGdo1I+aH2fSR5Y4n2UhlCyUvTUBJtBPACIpI
XLh6UxxAvlzEG3q3FSNvGKhVYI2SG1rwpXn1/TFi+Wl/XyhbIv3yosUmz4l26POF
jY81KMRqNKvDRI/9dX9+QZVZSuCX/UooG5xuC4GgYEFhM9+HoI/1ZAPfMAL7eQ+r
sq0WNfPoT13rTP3A12y6T4c4eeYw3njJuh4SB40GaxthtrV277LC/enRbpXZ/Sb3
txdfVluAxdZzXGvXOvRiSBdo4Gbg+8HQl227OaDOBeikzO8X8jVGwF8JB8+kHkib
1f8KXQK9VS07bKZtHwYnpYRmr4ZnyW1KeRlbw/w+F6ax9B5+rd0n9FdC+rhC/YH8
HTkzwQw3Y9V0vGoQDMQuDorTvs/+CrgSeMGuWFwVuNBHZFHKdADypzrpvchcxDyz
P9aCVN4XfWZNT+osUCNP2vaUyfos5Qzw66FmwaYJamz7whoCriNPgc32WXvVUWEG
2Uxe7Mv+IO6RLEQjlDeO+3Ud1tLKIq+MFbgbpHblC2qk0zjmo8eOZL1gkqlW96Mt
uanhhRJaCk+PWSp6lXq3+G0Nq9KuP8vh0ndUPBVrOUVnXnRyhd1iK7Porz+Z4Jej
4Yp1VF3+FvPkUUM+B2GqitqiC/l5TDeU4yJpuW8f+alB49jiiiOBeMGtdRYtjoLZ
IzD/SwJ6xw7O3r3rOsjMnsQlwALOsW4awxTsIdYLGLHWJNeQhBPazM/4ZP2rCSMd
FEceojoUgEZ2YX2hftYw0xCObJ7ATda1+VWG7celoTNxhYP9YaVZLSCBnMviCnXt
F8/ZUmRHZHnpHnKCGgT3hLU4UQ/SUTSMaNd30epe+w38eApUQDDA8GQADCCBTSmm
5rFnVSBrPJrQYdlP+voCK5yTT6dZRChh0iz5pwFg/i2weyZx6L/LnDFM855h5Hwg
yr35yxdMHzM9RwHrVoB4L/mUBOB7t1rB6twUR9yxz8U3JtwNocnrrnueY2pRabMP
pPq2EQZR/eKXyJkaH3bqYtxgayBvItgLH7sWf9mjL2e/bYgMj7VfyaB4BqGDki3G
lNMcbNSpzw9jjh2QCq09EijxKfEdwxrdheHlEGT2meyNqIBaZjBAhQo8vqrWBYIL
K1Vcip4xH+j+mFPZe2PwkEM6PPCSyMRYH26v9IczZ5hwc2rtph3ady3u7PYOyjh3
5QJAOdS5fzZ9vfLWkKOHOsPUJOj7zRQ/oNWlt1cgLAMpKLEnliT4vsE7UhdNGEu4
MmfWkZFWSHYgAnsjKqJZZZB9RNoZ6YlN7rJ77Z5z2tbd1WSbTnXaQOt5J6HI8f7U
UG7Cf/k87OM/z39IAQdc8eUyu9kI6GcnU4MRQ54eUEnA1e7n4e+3Y+lQeCrPPb8P
pPTi96yzpn+qLZdzxkn9CqrQNwouoDtWvlz2C8ztaFpskqEZ1etiNqQcD17ZpywM
lB2ETe7Rv+jzQP63/2D0yUzroHGRmvuH+GYU2480G8pM9tz8EcjCsMqHgHtELCga
+NPigejT1d5Mcwf8JNEPadDTDGB1D8Te9RA7RWjGnMIt4nQvW5GRqUiX/SIMoosM
tbRmzl8HSZUo1IFQkeDR9E+A7hZaid2qrKYZuZjWYtodkPXpxb2hYwoau5XDw1Cj
uRz8q8O/MuIK91kZ3lt+9+lbWCge8ouy7BTall1qiUmsAv8GQkMKQfxUKHEpqURu
4bR8vAp1vrCyE3lfjud9yLXxYiyedCZtbRgT4Pw2Jr2pOi+x9y9tSQ18qplI4QiE
sJM5rOKbTkaL8eT4FlufvjH4axk2Jz0Q2RTTHr8y5YyMPA5piLx1g+E6OqLAYlML
ueos7EYfxMb4+UoK6pHiCKooR8plul6ICV64P25T+x3tFeFKCXe0W8uXhDTv6VM8
aNLjBwQpXb0dPhS/VSct0LlD9Ni3+8jMLEYzLbJrrulP3JSWw3jjju01TZsZNibw
A7Xc0cmJmZ2wA48mak5YKTK/jXLw9ByeQaRVjC+dsl6kCsfnFVd46J4Ti28SUPbA
joBMzHWZWwmNCAkCCIWg87FQbXjzXS6fDW2ZU4QoxAPiy/ok2sRaKm1N3Lh9Woj9
GBUEpsqiQEUIJpMsz84HE0ODYnht9BnaUjUyZUKx0s2/bm4f0ErQo3KXlqjuomgL
z6bU/Oe0/Z78U5RHOowsmS3UVycO0b3rrz9yF2z6E/5S7XNSNHz2PSziLTw4DfaJ
diPqpWv9Z/zQ5v+jlCvwE2QQlgXhGxJSwlmq8uA9zkZnMdptfXE5PluioxhAwl2A
3Ly46Sh2CgiA/5h92m4zJojDaqgeVGpW+R6rkoUsGTCLPj3vZAY5XITLAtXJ51Yj
jhwIqkyczZ2vvAd0f6LGodk0KQXWtF6Bduh9nJgj3Yp9O65pCw2gJs58O9DnGuGG
leW8HpDKd4Wrs+8oGQ8U+Hp0jDOBu7tH+f/wKNYcttE/qaMmYEYdZRWgb4aweHS0
UN2UHOIeDjZ3zM+W+sMe+Mj4xsGlOQr0GFm2TDFOVZosiYySEaFyzJTfIJQNLCPd
tfYWTegKUWTOpXPTsr2U3DfPSBtdZvB6xvEbQxAEZ7Cm4KmUT0okkLyz4Z2qyB0Q
oOBohnhNKahvTVJPVj0zPvDVf9D+QnyTSwhRsPmxqhG1HmdyoRSWxx4/LYyM0AX6
6OD1EcGw3GKfD+4e/G9USp2L6wTSNI4hvbKhsb89HJiPMYC6sZnDBrJ1W4WjAj6L
FKRtjOMI0iau6AHNhA3csuCMTCaJQQtEoT3qG/0jbFDTI3EyeAKzjUOb4HZo+BRQ
O8dovg1LSewqVMSYk+hDnvQBiN/0AHdgWX69MNKjwuk6vEopndlRckoOUnChlVq2
qJnWHQSTii3DRoCz7O/Q4hDKlmOm7gGjgJhgdw1IfzarsyLuAGgwMJouiJZmzmBG
vLwNMPQhafyXu6Pj9W/fNWUP3cHxdojvF0lMFLEF+EqGUEBg3sIpKzqGWy2iUZiG
Aw0aCIhZu2LtPHk5q4XmFnHScVHTCvcKBANpErSwSUaQKphKNoqs02nvZrj48uDx
umjWhJkIkWHKwJ4dOLthHBshacaa2eECSV1bGIM+6VBGs5IlzMmwDMusw9OVB/q+
jlAh3domdcH5+WIzDXqqNwZ8idbODxGb3TjKCtxETNHd0ECiOzhmrGFeAxPSpwH+
QkoHXuSPtgIpOZGediddGPbAXlmOxcUhvF8JYVX+9g4VnQfSkAFdysE0cz7m+M7W
unlXtdPB385tDryBcAc9Ynf96po+UOHahcMxdlkdJdx+YBIgQQQUPP1J6eO9RHYn
rUE/p+PDYw+XlhhB5u9c3/9gNI/B2+rOeLcTonvGDuxbzTT3fBOceaI13ZiSRUKa
CCe6xRzj5frwn4tyki8GjjHe+T20qKQ5+3/4qYjyK4BfMQjq3kVQpeBugbH9QhON
EKiecxwgTdgZ6Z5/7MLXmL6c0/iJZXgt4A63ulFQMv+ApHCea5KYhogc/zP6pUfK
yTqqO/CjBXkKjaS89Tac7eE59AQjCn6td4WVqfbjV6uVaJxE2A3wHrCfLpqxA0FY
OEfPPDSxNoJ++2CrD0KcUb3vzuTj3RMfd/X0JJ8jIdam5pvpAb/I2gq0triYfPha
LtDHQhzLIzj6+88m8qPo0CBs3bEvPzlCh5GBJw4QVHThsYYYwMFF69tTstMBjQ/V
xDupIULXuVnb+e8UZzxqHQX9VYMCCsDYN0dM7qOCXI6frBmf5Mhyke42eZu2ZBmW
ENelzSrHi2wLcvvF+PA3lcVlqZiygYO9/sze9hj+wGLoFAQBgTBGdh7YBdaZ/DIf
lTQCHkj8kNflpAFDFZp5uBBspxO3MljCvZNsHdDEk4A=
`pragma protect end_protected
