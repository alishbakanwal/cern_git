// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:05:42 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
qxil+JbJtjZi4GI4zRmBjmUPmm6dmnFb7Lf7FNjUagQRikCMtTRzo/f/6VWtJoih
AjwGBvCZ35Q3+woTkj4poQxO6s1PDKyBSLQmucV33TQgw4Inm+RLYOwOZvxcrKA2
W4oNpcvvBN5mEN3UjGFQG3HOxDqTw0ibMD4TC66ZLGc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8272)
lb99qhc9/65XjPP9jBJZxgD1oC2k7Nsq0OQoELpVFlB8nRW7hMcFOjMIjA64e6gA
l6WRC41BrXycb0fbOhkAJivYSC5oRX0rnaybBnES5xb4SzPhxMnwnOlWIgMNdvAM
xusrEfml0zRTHa73i9Lt5F6E9dteMwQ6FkRA919sGuMXamLF+yrPxxvbbawt4vac
CMXp3ia+qxnqqt8uBB0JCQD3eeO4+opeQmQrPrSYmIl1m0pE1rBXIqT1Kce/Dbe7
sXlYvtXMZqNkPO4+GtfNBW12q/GnZ2q7R3Wppx/m2VwlmJ3rCDuo3xSRq966KiDq
8HHEOQkVNp3MIx/bw3yzF6aguOMr5PIiRVi9KpbTRRoPI/ArmS14Oa6XvpfB9xOX
VK9ERQSKgqrbu/HBm5qBSJbMsQGl4ff/WViih5W0GpPL3XToazS87S2309jquQv/
wnwuPB73QGNy/7cw+r6l4GphMstr4Wa+vRN89Q+DibVR2Si66sXs/VOd2f2AsRGQ
rZ12//9rTobgN1wrr5kq6YL+cXG4GsXOlAQNHtcadNWTpXIo0+poERZX8XDmMA2E
HyfEMqh+KNMEycysbl46bA35aTUh8OTcXs9cMPTNzRq41Q8Cw7hoPCzVkdgtDaux
MHPwOuiOpc9gAjB9KsXefI0mByK19g6ipAYfhFsaqTRQDGt28emaC+ZyJ8ZYVzO8
pVflIARD1SHpUzShbPrNocz1Cey7kOktyEWtqvztA+tP9uMaES+9v10C/jC3SrDv
yHcHeM4/iDx07STdhhasmEiu9E/fSpARiaOdsh7rmMyxXOj+dt6VT8i3Bo3c5g/d
dmhUxj1UYgmIj+PK4lay5ZJt7nkKJvJjDPx/lEfBUHzMhx5eL5iqhFPcLjF8KniK
dqk6JNh43t0sMZfKISIpn6cvc14YQHXvttEzZp+WC4fKGRAaSH4bLYqhzFRZ6q2z
joK4ueZ37D9idw5v+v9MvZXtRpmnLKMoKHBStlSNK3LJexSsWLKL9lUgOt24QI4F
4yYN/Xwm3MKWFmK2wJNQtkfkWYQRd0+MfedTqpiZA+mQtk8aTfbWQPMigL2jW2kV
/xhxJGwaW5xgLf5szRBsW9C3JUoXc7wu/JjLVtZSI6hp3jQBSjY8KcwxfuvfT2ut
ZF/AidNssmMyS100GaM2x1I4/CK5RUZ5yvUR2/L4CcsvDkTaqnlh9XAwUUYvFuzt
Vji53gIS/jlmOn3Uwvem2SPC9WSqZ+pYMCwntRq5h6Bz7MrEyQTw0Cy5KIT0m8yV
UG3SH9x5+WYuDSE8iVS8mctxur+wHogbSHqBgR8+0E/xjiDcIz0e6lUx2Mz7fsDZ
Zxm6sbd4AoDKYiAJ0jH2V2Jhz9aIX0uVV6UUeo4XgtpQRzA4sbUdcXJ0ZtwbO+0E
t5FPoytQBxU1C0QdtLbgiE1iV+koC/3AHWaYbh3OeRAulXP1IIrJ7rn+ImCu0jBp
AhpezvAjf1dg9aGVEBGClWB5u9YUiVDPURTC9i6nvHUgAGNhOTS4cRqT3SBsme0s
+P3UFmMWw3vYkicMHyg3CRokOg6AGr0+ksXHm7MTOyMp2f4a1UhdN+4ozdZsRxoW
CaOOZ2Pi+aSXGs/dUOrhBjWulu4LsAYdEb2VT3/u8TzqYDURuBN078ZXQ7P6pgDb
0LR5cadQ7jXONvxhZaWzfM1SojkRdPxCQrcDy5WhaUCXHCu8wOTyu4LNCfDKngL9
ywG6t3Zno8ytUM+NxK0o6ypV8YpqIiHAMHtbZo/NkCmyNNSR0cdTgbGh4l7wxROO
Bz15GGN3Vc0BO6GxH9LHAbo0WE4UDjrxItasonDrG5LKrrp4EWRLOb6KTrQgbzDP
HkXHz/72CybxSue/wAgSyje4bqhkcBVK7nhVnRHnItdRxp77Nl7l9jHG6DvSQRD5
QZAJds0Pja/Yqy9piHV0EJju5IrhwA6rZuZLI9mz3LTYhw9QyPpa6toK2fJE/4Mm
F95ONP00rCW8cKF4Yat0YyL9KL0i1+SN/f2WW4bDuHDrmm+qVvW/K3sVoKiIDvPm
/7R1DwpATmG3GlrdigOb8f1OKqgfU6ewQQjyawtEnTSIid7YKOz9WcZVQFuJW2Sx
ZrkRJBcqQBr9/8LvTFzZnaDhFSG92tY6MF9jXeZm2BJLVhZ8UfvLE/c2darIMWWt
Ze7DDW7z3nt/Vsb6VzWrP/syFS5EhSKP5SnKVoYmpekJDLDX2kQf6BvfxyE51O9V
W0R3dKJF/8GYBUFCEn37yMnsR/YVpG9MjIc2To7qnLVv9zrArrFB6XmJu9mpx8M/
igIkLIgVbfj7YIuiQSQ3o+nlyENPW4vccpgsDMsjFLXXVKVev2coaPM9DsUxTM7c
Cb8QOEZtWhZjhgoVYZ0hdZRKQNzYvr6j5azZ31dsiYGNHIEpwu7LfbhRb3GI9tk4
u97ycSgYFPVGpw9H3pv09jJQMs7yEl0oTw7TQ70QGneogOr6wymVtp3hVAORo9qC
A58eTmOSvtrPDD1NU/Tg4xQma/v+clRi2T/g8SDGxHiMd2wIMmLOccS8xfWlzSlO
9Rx/yx1pozck4aS++p6xNK7DCSlUvb39ecvObQVjyp1fEs6Z1GbaYoAj8njGYdWa
7oenEO39N3Gpoeo4tu2KzNE+JATsigCgflP40M06UuUBDPIqQT2v5ZBsw/g2xvkI
t9rfrPKpGPrjM2BvpHsmNdL7AdvDTf2yyTAo2FLW8TBkvx8kMnF4DZI8Qw47LpTe
zgxkpbwG0Gr34fXsVr2HcGtlPCtCuRi6Ei7z06QewVk3cMyjHZS0JKvFu35JJB1g
jvFMnCEK4j75UG6NVfRUOdpl9SfFTmdb1yF2fvl4uuEKKX+8WEhmOnxhKdC85ZsV
ZRDe0dCcffR3jTFSb2BtNhhAT9AW8nyFAstClgsV8yzplsAKnc4A0AF2uyQA55gk
Xj4MHt58R0SiDnsvkClBBqnBAkd310MpgN9Xc6rozx0OolRmmkupdhiiKf3gVM0u
BztpD/g/ElquyzSaHFPJjffIYIVdcmYeTm9kkPUuNZVvqbPhYzaT70cKQZN9nL9P
YDogEC+WUJWJcmcvIBMMueYY20zvyhAFcB1mSqj3MCa/DdpZp5PmTVh8hb0zClvU
BhUslcHYO05SNInV6WosgsDYP6uLW1bQ4fAV/95G00B9ndodZXC137uLc97D/8Pz
hPi1lzpyA195gRAxAi/hQVP1mQLSUyMwZM21Yho0u3SEzFt6gEvb2JK1BXxCzgc+
uDKEeU6tOp7xemfP2ljDZyyufHNZO5JEZ7U3YgOyaof1L6FtToF9QU+JYfIJMKts
JBegd3EZYZExCHOIVOen7NTWb/0hXRWIgAAaBh+lNBkHSGjE2ufbcCR4fecVgITC
QctV5ZJYpAzTXE8RYwVryJo9HscRiBuAGO8iZvPSNwZK9rsjSLMRG3ua6AVw6jeX
yT9BhDNfUL7EbYhR2Y/YK1OJGiM+Ayj29xyN/ctsSp9FRLMAmqE6HRanQg2TTYUO
+2SNbvBNr8ZbEpyoNmEIrQh0iaRBkYLdV5mDfz6o1AfJ39mrupzSgPNxlaHtTnsc
wV/Db4XzBYcrNGLecM0Iv/pzf5fQ1q2WLq3jZ0QW+o7YD5YsAen+dms0IneE76/3
3B4y9UDHUgBuE3HtXZjNB7XAJ/PoqOCkfgmJZfAo1oUf2fisE9KCmtvxggjrR/oM
DVoO9VH0WnYmq8f6qCjX3p63F29no2Iio7xzDGtsGyLZrCn0ApCxVoKotV+dPDJx
q460gA7Q31lo4b6GNwGv9wQFLskVStP9BoRjsar50tS9ni8+gzSg2bXu60R48CVY
ty4+govk8QW5QHuqHFbM34sK4alUij9sTaLDS5m8fT87li4HBdk0RgQpSAnRUj2V
pHfXP7JfdoWt2MjXpAx2CpCnvFceUlmrDlFBexgLTnVl6K6U1hTqJtjdu7lMpKSE
g8dOLezSdKZD5A/vNKNMEwyi9b9Zen0NXlosCVvQcSLNer6z2SgoxezrQ0RV1QG6
TDpsForJi2PEm9aewiin+bxQQwwfBkTx3zs/V31rC2HBRljqXm+WYEoQgVS3inBv
ukzUAuwvVG7cuIexb6bMWvkA1BVs4Xctd0yC1C9wbXqHdKM8PqaTJPqOhnORxpbb
p1inF016HUYYePEWLm99UoI83PIqHJ4K7wuzZJYXABJ/EP5ytit/7cns0WE0SOek
FjtrNTuHHVKcDEd1AZC8I82wECwARANn7sXBAaODxloKi9/YyjMtA7+CoGBlZGRb
UVWdU3njdyHNCQVRBnttfRlK4PxxFDmv6Cr2XuAIB+TsLhxdY/PPoWm0Mq9EeJCp
30gbeUb6OP0DivnCoTDywFG9bX8jgws/l1DvfuFQPKGNGfU9Af/46bEDr3LDginX
7/Cz8B+GG91fl18jS1NoFvtSy7xZ2BMKnuXOblN7sRA2k59lAgfbiV5wcIJy/XjB
axcEu2k/DcwInXlAbsy8b/1USU6umfBlo6grl8rg2sVq3ay2p7V9mEqRpkCFq7vl
r0+jWMwjl8vnjj3ycjaP4tWyIEtFqfp76h8vtUsYUq45+XkPBdpw4oJPkWQhZbZm
m6PPvTg7OLr3jkSxpZN0L/B9z3Tq3qSJut5YRbNmPHa+lN+9Eyae08y+PVi8NUG8
f10sk71LUK43tSij1EOKzmgmx9x0L/Nrgvi4TI4ZsS6oDa9jGaP0eBc9EbFOA16e
jF10wY5aj8QDugPlnSWpDo66zuNQYeVjg0S/j5w2C0hl8ugw+kdy7xihSGLCquoJ
HuZy8D1KJlQmQRqUfZX2Vk+6ROgklz++N7SWwJA0vYoC2CWMo7FecDGtyMJTN3GZ
+cSTcJHM28+mrODjPP9pljzTGY6k5berKiwN1YHZ2mpXiTcRupwdIemdhX/dmSVN
GzA6y/Xq7dS4kchNzE3N7QiaLoWhybVKEp4wgkNKlzombs3/r2nx8B4pF2MTfFgs
G18uHMPx24Je+kD1jLWCRzZU7Ewdl+seyrFb9rblMnsCqZqNKPGq1FaPmOQL888R
gGRHbdgRXpqy/uaLczx6N7lJlw62yUU/I2z0k+WX+n0U77/b0ZXxXQCltJHd9gj2
bPvenSB2EI9Yu5f5t/WZfDXFz9o67dvpTL/l/iQP0pdF00kBuFnxH1JoLvOvSBZv
yveLVa7cZ7N28k3ry2qGMmoB62bR1gA0C6PtKFPkIMBsv/gDYS1jVyEjDmpe66rb
4BmgiRd74ExUtBQY3x87OLXO368txqKPumCUhUQKk3vGHGN/1fHRerkTmiQxxTS3
RNqoXn9qNniN29g1d+RucGXtN0oqxpQRoKMCbWuXdl69cfEwJmqf4gsvFK1RF0rq
+tqj8FxGp2+olbrqboCTn8UT6CXNTFj9Q3KuAD5sf98zTWSeWQUJMxJ1jPzgVkRN
WQcN8ZvJD5Sl9yeXZOj8q0FilivWOREZJEFMacTM8mhcI3YAOM+O8rHQM231jdBt
hDGw8yJ55DA+tKrt92lGVgecvU4k41ea96VUzlREVCWcKIIMH6QI7errrQiUtHQw
QIz/p8Sm1Fn0JG0FB1a/h6/DRCjN9jI4P4yTfmwt58r6q2X9MFZ5V31Em+TYIt4s
OywpqLFX+PH2AEDe115ciMZCwmCMOrr95T2sRsOq8UTIW0YKpsN9ab9HnPa6AKb8
glveXxwGBG+J+rh6xMzOtr7XbtoqhosQe7raAt0XkmMj2qNGAmhDzQUNzI4GjI1t
5L2DmmvOX1SvEspM1P1/H4reJa86BNkFAHQCC5ATt+w0yrEzRa5UI7CAZ69dHLzK
144MRPxWdKyOl+LUXU5jcCOGJxpuqdmy7DjhK69rCdDV3AlCWyEwhlY45rlFxHZC
i0AdjNuz4lkllFM6v3g8/kEN+Zhux4VJTR+tbeo1GvZ+3ErymY8EBVrzWNt/oYQo
5kIfjBQXYDvAueigLJow+GjWOmdWbQ5hKy5XzeiMlch3+hIfSH24kupyOT1PPJiT
Mj2Z22Lv7dQp2yJmQk2BX/DqujCkxOQNgyOIKzkIyomie1nw5ba7qNn52Y75A66O
lfiAawhRqj0IvnkUlNCs7vfCNCyT926R2LZX0O/R5im3LHK0UobZp5r6YEDWnk8v
29AcoxS1X9PNHCX/vTztENoE8uM3cSTDr3IYZJtm8dXUZMtaYkAk9WNEoFvVCMgY
LGzcAg04vb5vgeN6w768KK9gWKVcPv4TuJD/YAA7n3qNLLlzwffOC+JRKcu8BhFt
0ZfFijFrHjeHdBeh/7fT9l4/HnnuBuMUDK1clv2r5BSvx3IKqGW/IcJ1ztN2ZuSE
mKENLQOlfSQ3+FhJaP35toLa5Ub4/qZSFRQG0JjeOfBUolEti609CtViFdq9uu4w
/mCxBiCN+S2thzLKEBd+3xlgI3GNc8oEL5riGE0EW8/w2bb8JyV/fOwSBG8frB6B
9wxLADDqD0MRHZWjG4yCRXspNDfz8kaGsVLkEfqn6z0EguGLFxfpQkHoK/Pw2idD
shUw0DbwuHgZ40Q3Ig0s++Ba1LBRclGmgc/68eSYO9LzZBPY5nydhslMb0maprs7
KbRS954KZTdvdWs8PY6Ps9fYn6ltzVnWqtwm2HAwNvE8edudJkFI5IgjnHbAbEah
y4emMHGikgTo1MwuykKn0TDSc/lM1mVuIkeGF/b4YElgl5hSA/hrVyfrdzaT6IfA
YYW5TKlP01MuSU/dNqYC8HV7bzAY+7BNEHqlyzT1wKcroPM7Fy7vrEdcd7lV51FJ
RV24kwm8eLE8PEI5Xk9hslYCC3ip9urIUjzJLv6VMjC7t2ly5wcI63hJRCPGQKM4
jWJfbqrTvD0pMIjlpPSf3GXIxZ6VKVD3TBF2ti+cp/gkdeumk7Act9FA1MxTGZnU
cwREfZaSTwSbGznW1cT786+62T6bY6pgNwvydFrxJb3nnunEMahvMbjSXA0ppRGD
PR5pzqZ5T0Bk+nwmFudZ5piPCHjvdwju71RmULuJ7eXG9mfzB3Hgza2znzBLTaZE
oIrp3AEr2YfpVbUrA4zadROJXWLIXfCTyd/4v5l6NZsmQvOtVa4Vj66fgkzBrKbg
wLSuwbPFMJbAgpz3Kpaxc0DTAR2F5k/odAUp0XNJzsQNFZht6pqxHTJmPGkH7zmK
fW0h8bCIJmwQNZMx+o41ogkj7rhrSKb13YPRWghvWod5vNa3lhfHSfobhD7A/dnK
0bx5QmJPNb/0/wOLXNI3w0xmNUOGSGidmuQFDezRPemzAxa1UkRP0GFhN1Ztd4Xm
bkmvNYDdSsiunTOYFpc/rX8sv5g0SChPwOpg6nchJi9hvy8xEK3cSjRyonsNh5X5
r/Kft4kzne7h2kQ+Pqyx/evph1T0KcWYNnK6b+vFH0ubeFBpjFIFTdUJ4oJzMSUj
XbDnKFXOxKpAG3XoGk94oaDv15Z3ADoksyvlNkcMbyPGQoWdRl8ypUVl533sYSK+
g/gai180qSjTjttYOuWSMzvVIGH1Qu0jHSX7Ns9JozQmvPhtxo6iuqTbTXrWeExf
WwFpN/H2gSTL6p3idhTEfqgX8CbY5VV0NbR/LlQfxGyGH8JhNsezPVGzv6FSRBRD
iQGeACtzKdFuBYhUmQXqackxGmMwDUz4yx6qqbP6CS2NCvGBZqNhaAKenBx1EpjT
Q28P4G3aI3RJxPhWK9+Dlk4zq2XOQhp8oCELJ/tTEq6+AUxcZ/gv7saRxpz+DCRz
V8Harv4nR5hy91xkMk19J/Ldk9qZnKtxsy5HJ8/tPs/le0r4rgWH5Ubn9zHbuAyR
kithplywqFYUMiUafmqtvOenUaoqgBmiXegp0eQq1emM7IWhmOs6a9l/yQ80QZsT
uZNePBIVe8EgkdwekX8JWxg9AbQDK4Hsy/HpIL8A9NhzGmZ9W6kfA5tlJYBaFpcZ
gGXW6E2yXQxW0/KNkCbtXZIE9tiLMqT/oqmXHsCTo87FIxX1oDnQmXvsdllj99Yl
E1pbBLFxn0gmjSJlICiStw1Ab2rFgcYPV/Y2PZNW7aDY0VbMV8VNKzlKyMxQfUID
+aMrztnNUW3jctGsu9ZD2ZpcJVbmSW7ZEbHCw1/WN+bAWpZSW2HBUB55mAQ9O+IY
kO5GTlCACryY+a5IYEdCnzRk7yAlW4OydcjXlrqEsg1PfYY/FV+yOLHaYXWgl79g
iFJtEgBZOj1uY+9HNe2rdZupgLCvelhsuA6iKIseUFEgHk2pvy7r6XBp/8BNqNUE
YafzXaykAa0dmHJ2/4i7oEmrgQF+gcuQ07pDIzFjzEWQJnMNrBBdcKhil4rEpHXF
oaa8Kc6eZEIf3g/8m9iqX7ZxrOS/qSoXgbm7fGL6l7/y2/f6fKUnA1ATk67ZHXJh
2zgy4dCau+sgwr+ssCUVLMV2E9SLjWZza8AVawc80bL4F5refqyVSUiLHk7sOsYz
IQc+lufRlMXeH6mgoLaaH6nXb9UiTSLyHx4v04ZYtnVJybMztKUSiWgcMlgIFfJf
hTqIJoeZL/ev1mJYJEJAj+j5pfv9lTfWnvuTnZsUtqIWkY/WlEi5wLQIMkHVm3/b
GpXmWoy0ICw9clJ4dQ06645hY9FDLvFdhQnbk0eh4KxEU0hZost60XTZF+qbohDR
nO7Rjt+1Z3qogANWvZQQuSLZbbMcBDCDU/lOYqLUvOXZW8UBSfKuJszLA/5UKu6M
GsyxcBIgN9U56REYyClo6J5QSQsMdfrPAyFcq9MLNHSRRJBt+uwDghOndSseO/hh
MVr/eWBORAsAcquprAYYsvhfoZrucXhm1r24La15wNFojLhkWzqOwappHEOEVEfR
PpJmaUDfMC2GZ1HCT9yR0g7gwG/Ax9LF+e6fTNCVVUasEaXGfqu7HNRsp9WfKJUg
XrJAVAJUIMRZLBTS824GZlvlOKKkgYsG2UUuF6zpnu3ecjcZXdejBiqoLQubEnAp
6umTAh4OplVw12QRuIhbZIrR8qdFHXD7YeFCuB84hKciorwNFKRm++9s51RBvb89
y+a54tIQtLlw9H+i8k70Fb+gQYxY0XUXXXMZlq2HHbL7HVbnyIawoR62kWw5QsiG
VTkBOrtgGCMTlEa6oiRX7i14wTzCHYeZR5t5PjKk88W1XJgYpqZj6HrtQB/m1mS0
gO98/Z3TqG77szU/0ysF2KVYLQ6hkAntHoEi+AhYo9aymJsBXs8EIY7TS7lXtEDO
C25z00gTpSxQOM3dfSjtethkJoELcyk6HsxkF1CKeK3PUZtZtaj9RPJxhspQ0kbS
YIQc4e7DGilXBDjDlhJ01xrH9xWbk1Bt7wCMYC5AnrSg1Sd3d+CcNuTCfNPfN4bF
Q4qxL5gNDR/uERBIMX/Z1IauAlYJ28L/vE36WsjBb2dkV/NLoHvU/D1zSwFvBcIc
I+8RuNOJklSy+uYFhLuSewT9juJaArRc9aThrMRnyuD5qX6AgUKfYvnTUVsatT0y
6NNg1Rz/qncufaCBV1GpwKm4ofphKBXfVDwTpfOJ7sIA5vTta86hOrH8jMR9FdJJ
3NPceHicgufI2ZaoeKDkN8kp39HP8g6oPfObSoKH3wlpMo5iHUUwC4y1fYi9FK3e
zdljczxGcmUrRsd+4KVc3frMg2Z2zvUPVn6ruNiWlAlMOyfYMNIWXsaj1a9gmtlt
ZU44sGAcYXXQorYm+uwjVbgMBOcpCsE8Nu7+Yb9mA2QW17k8IoynOCaSXWEl1yRA
v/yjqc7W2zWkf/ez2lICiNT5AFgsPvdw4xa2mC/SU9pw/YKZ0+JQ4fM5tlpSiFBk
SyC2v7eP3XG6eLjfgTAwuQH0jyQthLT66HU4lfK6weAaexxjnWyvqQAwCf4skmTZ
NNQxECRLbgrkXLaxx3pJ11vyEFZiEZ0PG8hkZL1rpW6or67Wn1qanWo3QVQj7xAT
2xDYZqKapb4aH+Uf4yCdCiWvo1jK+l8XjAN1fsXfneFUPL6Q/pWKpvj6crwKrwU2
XJLN3BvqhgjsumTFeqPyDdSMl2pg4Bkqn+gN3d2x2lNU5CuJM8Vu2B1G8AI8u0PA
xGT8JlREkJzfmKG09QHWXA2c4ZtcK5MxlR5gkEZ/vCYLIQJlOmUpF1n8HRP25ONz
SpxZMrYY92r2ifVNZiYx8QcykdiCk9ptirn0arb6e/PVZ6ErADszqG0/Z8AUicrQ
rXXoNquc+w0rBe2HTcwe20kuoCCuF9BmEtplMmxUWKkgG2Kpi5hVA7eqt1wjxlHH
5znnTgOHexQtUZX+XKmpQfAn4oXpmFqGW8huYnxTcFYqgipVUhe/0NLxwyDDS2JU
qMwGrtC1Y80Acaix+OHgtGQ9ra63rqX3+lAZ4kvQWKUK6ekrqZ5NK0DFgSaumRN1
MtbnWw1mbTtuB9kBVqzHBJUzL6IBbnzSSsYsAa/dfM23VPOiyzul5cgaoG7gSIGm
BAkWTkXh2+dD2UACzJ3V52EhGtbnLi6+i1Gtp+LFdd3H9qPjmc2Gd3JlVho9cGKi
uub8LOlTFlBDdF2DsutXNMxDbAiaRuhjjZSRb3sC/2put1QQ32TOnsJZLK/joyJp
knZ6zlBZ6A/Oibt22boN207thcvj9vFpKQwxEx4pFXGlmAX8eTdxFwMbCkiSNvEz
nvyXKoI2sRp2gkkc7qxT3+IUwDp/gV2pd3Edib8ky4atICVJN+LCAPU+w3UamgCz
P9rt2MhmNEIE7U5h52I35g+wROx8/TitekiB4jWBY0QRp6i09OFZHLIv0+gnMycG
l5uOU1gPgdOireYCLLxCwxoGjuywyb6eNgsgMjjCSkgmvJjLMw6z40mkEwzrdUJz
IoJXl/W/0iq+f5MiU0duz0STNnKkVhMroDDCUe/Dqqas0P1FNRrLMxjoHK6bP5rn
N+HpPCwUQha3o42TRiaDuUTblvxnYgSa8iKDHJ/5SpMO56GaLqG3P0xsrRiQWgij
O7Y7Pu3nh2o4JtpQHR/uzGTTtTvD4i9ASoQqFH3N1+TBJlOeiqLWr47KE8WPfSS+
dRV85rarCazD6MtcWNzfew==
`pragma protect end_protected
