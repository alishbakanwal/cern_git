// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:02:10 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
TmUxviVEA5tRe8f/0AzwUibZ7Aw5JiNKRbFDuoO0pzErjL9R+V5Lv3SkyhENVmF+
3yHjs2thvOs3lIJR98kF+aRysw7ZQmJ0KhgfBtwu07LYWj2Ge7k1b6NPw47lc436
WV8BuSY8QZa0wdraFzZiOowEaRKFgqRyA23aYtpSDi0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 19952)
wlRl3x2zMwFvjYJABXXgvjx1qIqgZwUlEYRgq83ibjHOllV2ebF5/u1uF8nEO/2g
dCLzqaXiGM3cTvwf1eh4q1cvZhb5sJlOqiqcLstFmswDzC6zCJl8laKsTUtFu9+e
dlewbGYrbmmuJhH029DJBxL/0RKysDs7OCu7+22p9RTvwtSqRgAkbzJ5wfhjiyPD
2ipAWEl7XPBC4nE67/qiirvPehId5i8ut/nLp1YRWTFnDqbTl/NeCNdxM38udwBs
sht/Uz/Id2xpNawvL3XujXPzjpQ3fLugMzZZqtGUCYh/WjIku+2V1qRH01ycrTlg
C4vDlJ5tccrVPe36t6cIsZs1oCJpfwxABKr8xnY+zoDkZGXUm/7H1LC9CsvX1T/n
FDV/vWXYvBtR4xaLWe0FdmNvx0a4aJl8KqLySxMg4sbKrvklOK9Syedl7ahV7s3K
V6vdGQynMKO207YcCT6jnKASehcDhpPxTaAMKw5iL62C++zu7crrvmSJCS6aBgwg
lsfHmHiK/BZrVyaNJiGYL1nmSjinIYUaxXjZ8ZugGTdcqoPwS0xd3Pv3OVZncMhS
TIx/popQYH5PQG/KlpjNiaDex+yIv/fenMgHSk6OT7W5R+jennOHw5eH7Cg/EW+8
TSkcCIxveqtumhcIIExESHQLN9DiCaDyMw6FaiOFrUq1zERHEEz40nUjDmLqY2KG
WBpntJG7QHZR0HupHVQWS2GMOKiXxsXSoxS5m7JOz05sO++YoIzQXoIH97WQPvfM
oHk+AEdu2FL6nIz0IOfzyQ1ZUxUhGap3pvAYRy7C3y+WQ+ZGn2nHJwB8SJzfSR3O
GRNzQz/Pv3rgGxJIWYc0sPn/S5vUTsTknlc9oBjYMQbwiVRth7Xme9kW/iFSMRx2
20L1UamNFQiKVZHceVTKKNCrbXfJl0KuA162NiVta3eO89Kmu+TjRj4BADhTJifQ
DV8xVDMQ9+ocj6xp0VsArbb5dheHWixGyC8/ywpWeZ/Mn6m1P//e43EwvBPrfOH+
95bcq9dUHe1Hs0B4krGz8adxo27j8J6rDksqnnn8NRuTa32ioz2CwaHubx3wmQpF
A8Qywsk+fghR94FSdoSOMQYtIYC1F8w7rdmZx6/fgK3RYwNHgYhADenoH3U2RyrW
rnu5F+qJ3VcS4OtXaJaex8Avl7LF+X6yR4baGHc65YRVAO3LrZDhKZFRp/5lWV0f
/hp0So1sR6C9YCyKnTUsY56LLGUkAOAsxMWF0DWwD03R9rAfHNpdIOtNdxFATgdl
XhTM6i+ySo9PBSGR6ucsKw9B/I60f2sNgW817CXfHpMbfemyuEl9wUlNYaCblHCH
McswJs0bSd9IulY+lNaaTA0B42ieLKD/ZKObcKAkp9hlFkm/GLP9/4c0m3NpUVwn
8WAGp1/XNQJLEDwRb5RZiUZf3O3zv5ouy5aBg/3U9z5CHDvWcR7Zt3LW9+E1TY3k
8v37PWZsSR3U8jubpPwDLGHuFk7rtrb4B7C4JQl4d4NuuBVBq/coD/vdYu3cJD4l
wzBr8etvT+LNosly1fanFk7yuLDyAOlkydmkVa7VKuKXsu+gL1bxBkWVp2eRI0iy
ViTJyzQmBL6EBSUsGtXqsBVKG9BkH1hhw7xp/PpgTSo7yG/fP2D1hpZcFnW/kXKS
Dq1VK65+1uDclcf1KhtXq9oyBaMBTDG3sxKsFIY2J7pLcfjwU44wJmZh7AzziqOZ
szotp0vAfQ4W8MLkTxBl8o3n8QbuV5IQTiokI0Dz4ROiwkqrburz6EDiLzndxl2H
O8QXBdEupdRBoifO4ovaki7rmaYk55mZp0VrFgLT8+QAQzcmLt9XJfBt2+8N3cxv
vHanbGpXwnMD+0Jw0n+z3kzNYKFS3envBbeHANPH1Lh8zHnnBNMAu/8gobMDLSUt
mg5eloJi9+GORn940KCd0EXZRoHZ/LuBuF2VOAv+qjTQIvClqtcaxmgelj+e4hRh
7QHq12EicNUTal45Buv/xEP+LoMEER7V++Ospph1KFnxlGMJ++gd+crmamNwczzZ
6ffo686PXS9X4YWyhb1sj6qR++fBfn18WcpZ1lJ+1XJ690xCRoVptCuxzeU371dR
dKkP3zEVnrwbyxXOZP/zHOcK3tFF9N68TDk5gTHEpL3Eplk6p0no/lpEZzhhTOFZ
cwY7lADWQPJDbcN4xHCyLcWXdCgixt4NnkxfYC/4UBbGdJlHOoly7zqU7pRt1uQ3
PaqBJvnJQo+uuPAv/KkvTGyQF/5wwwS3zAf7711y0weKPq2NeD30ARdy0qTgvKZ3
EJkdxc1YP1bqeBkX7DQ3DdpwRKafyp71yf2FlNNGlWmaRpCH8QnkXRHBJV8D6KnF
3hFwJFL7TxQgrCaNlf41jH+CH+PlA/fhstiXOd+iT7zwpO5ig2217j63SpPFQy0T
HErO5hrmQmVSIBxCQ+ggj9nGj2di3gw5hyNzFp8/Hr+xCBx/t6cwwp+sCBwVc2jh
AR2EcbwtJRYbGdHB1IYhlaj75AL2tpKzLE6f6nHy2qrqzHrV7/d8t1SEU2ETOt3N
uBijdkAvmlhTgHRDk4Q3af3BNYOdejkrQSDnkXlApzZ0UOn+9Og2jsE/HINHiXj8
hE473A6WXtRn5EuYQIqHZHNQJUak8WVAM9/rkpNU/FTAX1mkn7pFiV1Tv820Rdvq
6Ya1VhNWOWFlQhTwFglrlH91TCtSAw35jLrlsDyhR7TklZzDz6vvYeHDTeXDZFpE
r27cqpmq2DMto/6igsp6K3X8+p85rBvM8yflcpFPWvIMBzmDnxhmGustuLS1BQv9
lQlPDbIJT/0/hHLuk7kmWDSPS3MCCMSQ1A2ASkd5RscNsRhaaCuZV9+9eHSElgq/
7gxIOLdS57CctCis1amVsmoBG9ibmupNs8hHoYS/DRuH6iCz2eg9VKTqXaIjRhUW
QRU7ejc6jFOd45QfPcXomPM/Tp/60ef1+U52PbD/W2HJUl4t2jrrdvwmp/w2hC47
MuBRG+lBAIZt3dZoub09gV1YypPvAfVYssjC3Ys+LNXnAXTcW0qa/mVYOqeXld3j
gQ6N+BAkGikBc+Ox7IwhKJm3nv7n+X5E7zLLEx2bVMXXW9aY9Jvw8gifqgsM5YHa
gwiBHbRq4k/cZCJKpC5YtDFPcsAoM/jkQtt17Wfdgcq38anz0/hbiyWHxXpZdnbG
pOsS2VTFY9PPF88J8KYIuUt6L51Fejldc1Glk5ZX3pIDxaETZIscZVgneEVoHalE
jGQZU+eql73Uzua+DE9TzjBj6WWyFIUazg+QMHP5yw3/hJiMSrzfF8zLSNoOcfhD
zuwkHU3w9DGbZTQwNooGCBEValxDLM1zM3EYsu96w0dmpK84j5wrhLP2J0AN5Hwo
UcukmwUU171A41U7cB3393pvbMu9onHDNDFb2LWqV1k8UnjgpK1hsgU4j3xMyTZB
JJsUgifCpQojEwrTnD4Ccz2KZxR34LdV2u4Qi4QcrbIDEPiSbVd1IK6hv4t7+Ea+
ThgbYdIH2wdE/2AB8tdmDHk73lIE2gEvNtjW+LHcZ4DEyu0skGnHzWI3IDsVcZQR
MDPGuvNuptCCEW2qAgo7TaTC89JwYccnWml/jK0V8LK1Sumf8Q5ZWAKBW6V76mkN
MeaQeEwd/T7D7jBeoJfNmzc7K7zSS4Vdi50PgDiTio0Sb1+1yRugBWTKB7JqaexV
VLmmwLX2ff1a4A1/NGzYb3+L4ELLIl8j0CYmZ2UVC2LzYueUG49ra7isuVqdd/O+
XZ2pbvCbj7wy1Gk9N9jOcC7kFOVTvMNdYOHEvMNVO0fxPvxPUSpD2wQSpioHxcw5
rkAuIJkdkODVrFD4cG5PC2odHMSfv1CbarfetFrAy+GzKBm6upWQ36uuXDvwLMtg
MYQpRPmgwOsYlWsml0dYoP1b4eHJskX1mjiJ8R9kyGsiQyfsw2jmlwak8JJcO/Ul
1PUWisbRLXOBhpUuOQluSnnVSWEooLogYh8Dkrcq1a3gbI7RieMqOWAZnbWcLgqT
ZKejvjlXVkwrblhXIeMFMLnSdPE7V5c6kuiBmtj5b45L820nFtg2A3RhI1065Adg
t/suScNGX6GA5IHqhrzPy+f07sGFDtOAOSnkHRWXYF/kQqT8ngbYTs5iXmzAtxF3
cpMxl9vCD61AjFN9hBcqHGWopP4w8pAJR6rwlhT3ddXJxTIrqBPUjjjDq9MHsdLf
3Gxgjppj2HiDrbt2x/Lfv72koxC9VXUUiykpM8gUkd4EBeSQ7ZuuW/KX7r3b7zX3
rd0wkI+XD/AfB0VAibObX0GqKtg52LPsAx4F5gHSCI82z1r9K6cDwAUBcQu947oL
t+XZy1P0Bn1rGNkA8k9nPPdk9l1e15KUIooV11Pb/ndCgUQsgF8Yxt1gCT4Jo8Qj
oxrqamF1avmn2r+4TbIkahCq75hVjfNGxYs/v9m/RXg+WmSaCi04IWWKLKBmSRBt
1oijNwUFk2Y9+BZ0a09foxDLYrxGpWsNktcwUgfPTkAGi/J3eYWkLh6ammKdvnHy
GMz0zuw/coEi3jCm5vRT47ASufrsCObEGjDeq3Ou2ShQaQKqheJhmAHHvjWL6IfC
b8FZ0TUCT0bitcvbq5sfGgjKrLmrdEJdK9YGJjh0xs2/bGynPZaHhFDHb4aZ7Ma1
EjfFiH8Pmd8U+i2tHmXp7xSx7w6srRH7hhIqLjdew3Q2FHuhQ/uTIXIKU/xZpr7g
guVPiTP+rnxQZCAk3cyf8b10IcC5zAguK3tJNX+cNkv2+qN3pkK/uTaBGSD6uDmv
M11cHm9QoSdv36PJwEmaGS+BU/TA7wuYXjAef1BRW+GvH1OIS/WixsUGNEVznvvF
sDo9bJ7FdWZ0nSwq9WWmssEkIpT3YR25WppeRk+jmp+VZT7H8u1+tD/7vJhQLIU8
U4Jj9nsmm/qHWoHrtsy1POdZSyiOhI2UwGx7+u7j3/KV/0ctRhrKHUio3/oUMTdC
RiUlSOFr2NO25y2EtMbAGh3Dsa/gKJNuWvM3CjCWsC2XNFv7Twbo2OUZh4/XNhug
ZyDw5SCAQmbzpuBsSQgE/VHu1YN5oDv6Ie+rtZo1dKCoHTLanpkWtcbe0YeKgtlP
E7nG8riXjdBum/W0129rP2OrwAbkBAZ9hHRXRtj6LbS3BUMaoxYCXUZFXTmKMUBp
QbvODyDtT5m8YWx9IQDO7OTyMdyq+RuiMOMKCwMGsAvywEqjvg4zoX+irzkjCZju
ccLDqemj3vm3/z98diON46RG2+0ZsF/ym2cs1tG/2Yll97UiIr+u4/UdU7x0Kpr8
ryyNeKpL3tuLVRXUp7i3ELYA1S8KE2w8rXGY3TSl7qjnGcJRgAr/D1wGfsQxKDK0
9U0YsAaqhZrX+ZnAySRW9tt0uB33/9GC1Vv8GumMEsRtDoN2RSVLbibVnfRLD6+/
6ToDYyqiIIvS9q9i1C4hZGWTvsJ3zEqiMcidBt3QW53yrqHJWvaXJc8L4jrypZCb
RDpKoFMXAv0MXWrBlTIPoI2PmqZWx2zkrCY647Fm5wd7vay5AJ1SA9FSZrs9B7t1
xIGL85l0X7JFfAD4fsZrxb0CTreYJAwU1peIils5iHE4FaW4zZvoyt2SD0x0c43D
+ELocKxWS3OKURG7TDUzYM9s5Y3CSIkKZKk1XixLXvQVEIMqcF/s8TINiKmz5R1r
1U9CIXInHUFL4SSmCZXDXXs4XAl5HwZa93620eXKNKF2vleV569qq07Wdpga6Wfv
pI3opfXQne1/jWR3zxlqpMiavxiX8ZJ5J4P/MBGub0vjfTsq5OFoxIM6V7p8gHiC
B9xbyY+XvAD3NtoeQTI6awVqU0FzThXHvBGqre1d5LCNb4Bdk1jWWb7G2Ws/+995
wpYpklVToVPx7gkaDd9JA7yWWVWOZG5WT8EPsArtTUKZf3jGLlP9usUh+/aVE2OO
WD/x6GBxEbtweHtIT0jwUsgUx0I8C+ruga47NHyjQRAzEUOcFy3w6ko5mOVna+wT
XzK5VwZESssg6qSUOfUO+sck6Nr9HedX49lmVEv3l0Ry/aAfH98vOwBCmI9bseTM
t8Bpwo9OYt0XPQULcQcnWkdqcLezHZbqgXiDwe2JVPkLEP+B3cdD9bYA8PrafeFl
4stvnTHItEPgze0FQowbxEj/eajkyAiO7evvzYCcVSoJCYyUOxB4Cv0YO0Ngku+5
gv309PFT5YyXIb78040NrOKMy0y4jJknI8LHMiNUPlAhnOVss+mjiVkCYHVvJ9zk
RtATGzuyBkxfMD8YPIN6WPHDqQTN8llM6xitGGuua3BNL1XlDDxfgo19a3B62f+E
rJsq0YrZ1xVTJyc9NwDnhKIYpQMO1z4Rv/bIVh9sfxUYufc27FWoutk9y15DSQ0Q
KGy4jlmmWiin1jgRYcKSD10VqOHUNJivSG9vuGa7HXaweXfOLqxGw2jj842j0n7O
Jna+cl2kpaxpEnGikS+TsuzD1IdoEvGIM1Nhr47b2n93QItMcqDKKb4eVw1mzB9+
Hbvl8mUdIA4WzfUwVWwe9uXruzgG3kIVVtCnlJhmJ6IdB3/Kr9FTdqHmDZ/TYlTU
YOpHVXcaEkBgK6ceSRdKJ/ZSEkL2PDNI2nO+QXQm9bzgG+S0oPbdDXKKI4TEM1CI
ZvENs7iKsiYfIo+ztD9ecJIa2YxSDKT8qv6cEpLqD1wOroObU+jIq6/tug7ITfhS
HyAQAkpOD8OVGJ259mQt0JmqKRGKCTZUTsoCVHEWIY+01VJTkkgEZ9iCy8GPKc14
E8NwIY0RnPnDyiRHoJkcNi51VlYqLAuhDKS3IZCF3A+pECLkZMDTMuiAX19dbMtk
Mnr2g5ogeL3ZJFjtqui8fsqVO4uSp8gDdXSQLEdaxlw7eZLhWjEzHXbAvOzp1o9m
wP5sg2HGyoqmiaS91E6Q81YbprqxDN9NqGxWIizgtpLzg7dkRR8foRTE9prmZASM
eZsKzQW3uDLtIBkcko5EQ0B3eAMsFEUXhmoY0BuTZkF8OueBq1QQZmSnlbU70/je
R9NpfJjjg9wo+QKkaVq560PPGKo1jVWiGTpxKQ8v1oYS5SvJ+aiYYLjQNdHKfVg/
YljwooQqTDc+3J5d8obP0tObj67pTUJN7cRqQsaeF1kxa44hufza8XLqH2wSjEAr
llCZ9WA+JwTr/eBikrZEVXOtmEFGM2vKQes8VxghDzr64mvFdeaco6QvFkXMHqF7
hng/tHZ6kju1A0CvK4ancxOhANpRC6pT4LfxnSw7DADZ8Ts/56b9pZjKMf+rkGr5
zvQ3zUM0cgX6YAI5dGrgQrWozb9Bl39lllolrEgHypeyfPmS3qJh7e+86dJK/t7J
dZTgytNZqHITuD/rAUDl5HmI0MoHFbFGUZfTOqAoW6AHUEX6Kzt6YLGDWEwNvLzl
Sxhn6VvpBnA2w5c+477zEVb92yKhJ/cBmuDiUY89G5q3uy5+TTd3KwQ+r5gF9SoB
qJFUWwCY28kpUX6cHTcu1N6va3QhyYLvZjVQSZjpEzRPinZwnWJqwHpAACJxDbGY
hJg9I/Qfb/qEpwpZZdUZ4la4ZD6HWLHSS8N64uDN6VcNbHFi3qHdfc/dLI5a3pRE
bmyhhmaQIA0zKRvZ5cfCQXH92eTqEiKfU96YJa6hJ/BRq5PudfLFabyFLoClso66
n4nC9Sbkj53MnyUeVhtClNDJWc2TsfUbydYEt/ggtVv5x3xWjlOwDnATD4hVtunQ
4H+BKxmVBZe57OgssLEiGRyy5NldZY68i2HY0VFHvMzvm5F1/QpeBzYUGj17k1eu
mnrHxfi5jM23r2QDa4u+DLEDUJ3MSmgNHxfOJ8XhYOMwP7+RFWp9mDbglfFOgmDQ
wBetT24UVb4KsbONIr/xMEuLrMmXFHoDpKyfr5nffusyMgboNr9hSLL9IrvQXjCD
3Ixn3kox6mqpnTZNLapjCsTC9k79ymRzzFnDbA66sKwMEc6oYYbd0Xtvfb4cvsHU
RK64DZ2TKpM/PeB1uE3PQFKxaKIMkYIMt1c5857chJTkUcpZlY5Gp0reccxIhUPp
KsFJQgk+/DbSV/JWkD/sgZjo+STbZ75F8imBGB4NKQjQI/Lyj5t+cLYqCy41r0Gf
O/aEt43zbV0/QX4JFmIACqGyJnsAb+BevfTWUBgCsC1IEBw01rFN3g4lQNa9Fopv
D4RvJ29hbJVJW0QThu2G28cReQksrehhEklTQQeq5PSuxSm4FHyeHskIN9DSw77L
7y+21wVgzj1C7Il31bSU8WS0n/xkFl6uQQ5V/3rZ3jlTByWQwqY/9oc3XEXRYhxy
SPlUUEMvgttv9yC2PjGuQRZGflZLf2VYoT5VNTz0318k1Mn7zYfiTLY8tbx+04SX
OlcR8rFKjo4bpTA/pqJWPvJNluPspxOqXb+GIBN0EjCzwJABOo46ulbmvaRqHCWr
W/sn/Ljs4I0v7VL9PnG6zztpLaFCVIuGx3cLpJ6Cvu+Y+s80VGcPJOzHjNeL3op+
HEXFilarOk27ZCTUBPtJg6PYsnT+g/Oxgfv1uqAlaZcE+X90J42mkPilmwReUs2n
ps8RwjzjeQdODIDca18dguit0uwMe2D4mEmbk2TRPNthbLZYTAcb204501NDrltZ
XoIteqiKsFRF5AqJRyU/q9qRIAffIZw10Nsug85goe5qHagCERSacOojmODb6ojm
pnbWouc39WCj7jIaI+E//ApnmZfQrULWz9SkhJo2841cGZpy5xnvTjmtgbljD4/T
RctEfWu3J6CZio+xeHu7oAWdDbtIWyBTBgwut49Aw/+8tkKD0cvf/jUwav6OBUWk
DlfENe7MMAchBYJMiDzM04c1FsW/EGmZT/j1vjyd2Fmu/uky8IJgw1T0HbPbBr/d
DpEh4M2dBRq0osrNSSTaWF6bLi9Iw1Sfwiu6yMcH1GosF+SQzoV2O7v7hqqr949N
YBym1j9zstYraR9vKYJvTG1WJpwFQsbGMwbstBlk2Ii21Hw4DVksuGw6hfewesxN
51RnW+p0UiAJzUQsZkgUjrlMpZ371FEKb6g9W5okiIpS3njn3DyvPGA9l2rZcNYS
b6d9W/kwCjirNoJ0cpT/WxWNQotdRYJ52avfJwVzTtpJV0RW+Ho0a7thcosKJw1M
GiUr+MkSUobqEm9Tr72s6agAQBI+pN1Z9iNjMwwrZEgCnwTabXksIy9Uc/aTveLW
nQgIVCH89OuV0OpN8xEldQWYUI4acrBGMVqa30dFjEm5Qc84G2aPwh0q8+LuRWf2
J9LbG/pdd2s3gwm12jc1qzYUNBtz/BfkenoNNa7W2LAMfAy3rqQMzSZcYfIsEYrZ
m2WF0Y7Xp9PBZfGtCPkTVXTEiUzhaH5uBGmvbsZBf9GlvDiwbi1fRFl0+Kbsoy3p
0MYrU2UQyN0nwxxML4ktF9vB55cEVeEBv4YOAhZMlRP+ysUpLJ42uS8wf3Lqaq3y
XZanzdHvGvYgcI23XXbU53+wDh8H9vju+rM6qL7R0hoO/vrsP2JWODWr90WSHw54
mHGevEv0u++IYMeG5boEqfWqXbD7hTnFl0x/5h+kd3h4WXZU5nTQO47V9dcTqqmE
4LVSw5zJzq8HkLeK+MZIthH4Z+g7XBmt8R8rU5EVh1KxlxQpOE9ibjyPTKSd0Bu2
4VcZ6/LeIxIoxsHVmGmaHr4gVeHhU5Cp8VW558SWEzYgphwiLAzw6Eme0Vbqy/Ih
HLKx4JVG6YBz1xufmBOZctq2Rw0kPcNM+GwUdvWPqo+Tl5IeI1ASy8cHeI58TeLL
XpJPqWe+ylqHE7DzDWTZR44BKZ12hQcYw6EJXDmBNZ/DwiM0wc3BsRX+6jxlApqB
sZj0ca0H4lki9XwOFnhamZdwmztMbReXshiuN3Nrsxe1RTXqScY6f3g6ezQEFl/I
nU7rJQn7zFCGqcrSE4qirnz7ZYg7pD0+1aU3HZr/ugIJTDDzbTe0MNseyZbQnHBh
+AQA6nVcKC6I3TgBDox3Y33ilcHVo38kEroumorDRfkUbh4t7GlmnbwQCTWVGN70
b1/bSYZ/bLYx4AxkdiOV/84XRwjw5ih6k4++9i49ML3kapnefghhAf1lda0HtWwK
gpb9t+KL7uSL8/FQ38xii+MxuaATsUgyYkByVE0q5SOC4t8y2hjyYUQ20G6nfJDp
NdZq61TiiTCKYhO9BX/d3JaUzcE7mBjegD+qs15GGtd5EcDNMELQdh7HfIVf0ULx
Lfx8TTNEHMMLnHQWlbCCrW56tyrM/llMRokM69CgoQGZes/8CrZUgoy+uzpgQtcB
GcNbfv4msABohWvD9nqZ/b8K9KaUnvtKSay01stl7hl3fKxsHGTKSXHCvJNgLp1S
ydxz27thTdFRihDU2Eam6y29yQQVY5irhdJBpnUZC+S/IKEquhu9C7tbk4HVBF9C
jFnRmhQKXKg+zOxRYooBMX6FL4FIsqpaQ6mJh64PTVMwqaHN/TXBHbHYM19V2BOw
5j73X6QcPQEoYCayk3mzQu2+4csogij+nS2g3cZQFWQROyPzOrFQ0RxXAqk7ZCEa
lf5mRwbO/NVZZGbLQoOss/+gjbPtcEeGD3owRjWKhEpTrB2XirDMin4T/hzkgHRK
jxoX+4wvBhCqpMEga29HyMHthq3PqmAWPUpSMvQCcQODnTLpdTRo+iQkbySbnCjr
sCHKVRheFZTU/lSSvvt3xYwITTnnpb9OyzZXnX6QKUdJMOoTtzsMNdx+ahhttNK4
sHzgCHm/HH7L+Cg0PNmjKD21W1F3t8u5SebfaasfwDU594oR5Kf8hJHHLoV6aQ0r
FymDC/dCUT773zRafJPe7Pc/DdfAae/xTRJwkX/EbRNQIk/4yuxZOTlB7Vls6xrP
70L01SpgZBAPTRZTQBr9kJbvOMPp/xRx3pqEr0hyfv9MK+15iem80QJtQR9+BpOD
Q9AMef9u49jKNBK7kul1VJliEnj5zFKQ4Gqe2ZyPcoX2PUGeD/lh75aDqQ5zKIe0
UhOkaTzRMQBdGiUBDM7ESMxjGQffMZgzZEmaZ+fmbOkvWedr9sHn18vtLQTvjVGo
N1jMoQMbDpEnMfiz2Akif3AXJATRvWfW3LbQ9Pw2SXx6awHIJfT3gPNUiCmCS/8A
efr66GGk9O6DUU5uzKWMrJA9UvihbIQoftRSxvcASE+UKIrET+0DhwNF5s3rYkEN
cN/6MJMKvQJW5SdIzMezk37c/fsHcEg5BrdJbmYKAF/78ogmzp5Tx4o2jEnDg5kt
i7WjMZSK/Y/WY0GV0QmQk0vj+mxcnYfUWiu86z80aAIIx68J0v45MDfsjwEBcCQR
Qv8VMvMIvGmxAPnGFAxlbBSQd/vWmhdYa5WBU+uMPgaiROvk2vQNs4IF56RVtAmr
QRbxi0R6wWYBXqzDHvoJRJbLAjG/RrPaeHF241h/i/dLAhaSJ4CFu1mISQfqNUmy
SBIgeEBrOS8mzi3dbPFB4RgVZJjCOCIQhiUlGL6OW0OTSM5O3V/7xoafxl9pT5DK
96N3ondKydABBHP8scUEhOsDBVPfGFpc+0yJOC6lNW3oh0S+5JMV2Xn7S0HG55Ip
KMbkj8/s8kUnRqXGoWJa8l9n6VZ24yKAdVL8Yw08yB1TGGVyocHde0L2KY4SryUH
g0mwH7W25Gjd+u9fD6buOGbxaG70UHVmUl/KyHM5vsbt7+64G5Oi7vVbU94dpXs/
TJjfaz3vR9R+LTPYkF13PBR1MvgGWsB+4SFwyWyUZvKN5XjCtDv174J2WaK/qbUy
ATmD4mfhVgKQ+Ol5lZPb/PssET083aN407cCVyzvA/dXuITnXe6nqlVljXpk4TRi
oG/UX5/M+wOaTRFBZhmP/sc/izYLS4hlvK1SrBiGC20q9Z8GPtWL6R3gAIfbwbMt
HBWrv2LxLcVRnr+SfLs19uBtUqMh6MF8o2nqE0qGeZxeYFTqnINJcCVsCSAVPT6P
6TNHOhk9HsJkGKOzUs9bIZaq2W/5e0AAnoMpzeRgCQlrtWV+nO4jcHqQruY+3OLb
isBxIsBYO43SN0AYKBLP4+ixR/b73akT+zdv6IBYmeuuMf0U6jzpCzhEn4YRx/+k
6oIMMplG6TzCMlXR1cbIBPv30zpyPEHq0h2nqWAmTFS2liz6hEIyaIJbQlsGY6MG
SL2+hZKSpeahBxyijWCU23+V66Zn6tKxpR3YIn1dGjv7YAHXC1TWTPEBhghfyRFq
K8bNEpVhCPYhw7+c1zCd6WdFYTX36YFaUfNj9sAbUlviH93JHdBodSeD+W0MG13Q
gxblfx6RxqbQePIathZh3N/kvcGKAsLwrw1fe/jDwsBNCLLPptFJPEtnIM+wra9v
A1JfEVodW1e5EsaSFfOF+vg9dOWhWJzyS3DasVhjwwzR84pOB7tMhLG1bMH9swDd
QdaXpOgaeXeGTevSZ988cqQFIrg5cSFjcEUjPiAXPbO9QmRHsRLgzSULE3Bab0mA
/uk9Lvab9kcjy4nUjiQaFdroz2onJikEoSpMh9W8VV9YnX8U1MU/wTXAwkbbkaj0
iY5zgOk3EYmumU0FO2VQrlH9rlf/BTKcJsAnHbzn5NExUWqf8pp/7dHufvK1v/3N
4utpGBGOZA9r+ONO37UYp5VAsI4xHHJw4OV/2eMK26zdfLxmwdsIvqBLoADCKk7z
B4eGFCT8/iGx76YB9429WZRZU4Hj3cd4UVJwKDzAzPotZLuUaQ9BIO2csq1lItCf
BY+rHTkhhYQCJ1uYDLbxDty6z4jMppvSSZsTa+zcdzX9V8S1pXvGZkHlfkDEjyBs
6sdUImOQEPqa1cpz7QxlRQy4HPD0Z+QcxH9etw3OPSkDsM8FK/8QTcXGqW5PFbm9
JhAhjT/HgSvcVUKDgiHO6DG7y6DSQTABIo6hRbzIRXrhtqM2e+cSJnJLVKEgUkT/
697WmjlXJUc7mOk5MFcTe8KH7oPrjs8Y9cp2XHACfcLTZwFtSRsOmtwR2CU+uQUl
fN8JgEJ6Vbbt6HdO3iFc690Cedqj4cwBa719QeGG5QjZ1Dq0QGpf7UySO1xs+Xjk
RwWBzhYtkow1URSSjhYMjV2c/+HpVvLvoQvXjczOHDOX4zeYx79OG5PLOgU8xwcd
VGvA7igBTzt3YZ7kw2bb1cVuH43wSeawyigXNEGdDq5xeA3NPadza6MTaQXtNIqb
8t4V79Xw0pvfzqS5r294lH0L7jKF75HDwp4VGht3TzI+DkR6Pn0BUP2uBST4LPlg
kjiMXQuTLTpdIUj+kYxlUpVNmlAoG0fdVOTefnMnKLsBa9bAl57yC/G2VfN+51EI
+jVPlBr6mmZYWORrjnqpEVMRaGRsaRwebReIzsKsKwV08YXiYy0o2s1+coJ1gB3R
WsX0iLLxmkphI3/ePlHCNrGZuK77HWxe6ygfOtTf9KKZBv3KPl8CGbbF1mBGRHwR
EfsSeiEi+dY5oi07RKYuKrS9BvXd+OoD350StvAAWgzx4GwPPTz6+IXNya8mongn
SAHelDZoywJqfZkJqcKvSX3nrjDdEUr/W+uMonUtKKdYl+my3covMZiI8iS2NYsv
nLSOQvvAOikw8kxZJMX7p40lUV4jESxi9P+FSHf0JMT+86caLU+lYZF3CbGz3EPu
bXnZunIpDpQpVINfcWCdVAk0niTo7BA0lDycE1mOJZVPYqPCIOgzJzPmoQN25AQT
hCSXXH9uJ7MgkxWR7UcZVHsGbHxChHG5k3bYjR/xvotL2tphF7QcVpd+scQ2XTuQ
/U/6US27Gw3mb014AqDfao3QzSvYQNdC1q8ro5emUWxuvSpFiIerw2ZHdQ92sm7O
uI9KTuYYvLWHTJenQVD6VK1CJWzH5D/qCn9Tybtmwz3ZEyHO/ZVoOphx0fo3Of4+
yCL4L7aKzHxd9sjUPDcDdh6LluhTD/KAfJkyT6PqFaGKRyaw3bF7lEDhiEP0hCRh
5rx3LsBYXn6/R6Iyb6HOOW/5t+Afi4dsVMFaqUgGJFfBvUAEiibB1PZj+nn/cpKg
Fh4TlGH8iZo/tmkfYaJ5e0w4GK4VTb5fwTspKL+Kwo1BKpT2gvzXzJWy5nj8h77s
5ldEUxnT+YvKHDFnEaVovU6kykeO8luzTTIuRJGk18FlDEBz5cYRTTBIBnP7VX/N
n64cjA80N4Xq4pLijyM7YO2ZBMy+Cm2g99+T4tXnX6PHrcSbRwESJxp3gcnZsy0p
jYCRjrI12MkxH3gUZcD/VGAg/AUuF5z+yno71Gut6kh94bmkIOQRajYQkQrVp0Bt
jEd8Z4V9j/EI9oS7iGbrSMN6ciuM8K5zTBFYF+CZD5CCGCfAitfQh5WMrkdzfc7p
NzxgZEiC73d2Vv9+nkSGQT1oetNx8dL7pu81Tf5cZTb/t5ydSO8M0EqBg1SF5bdA
EPsZ/R6/XF5mzeRj2b+9gT8xHeRWvgF0XUlSM2YDMdDoENHWfuE7NeK6U0waJ+hq
9Azzup0jukqs9/316RfWGPyDGGCR0pcBtaJL6swNNKsrb7Wkm7v5o+aZyD5XFhGo
RenyDsEc92/kwbbOLSBonxbepgloDemg0Shi4S35ljAFmAqmALo28Zx3sT7agRjK
KTbo7sUnA/LH4cF7WuJYBmxUDTKHEDBKyFU0kHbnrqkUpPN5tBLMF1tATUFnks5g
dT7px7tzhgBc/8YwwawGFn0UABB9zD8fx8UUDkIZQPqWVIK2mtLqt2L+tzw2vzs4
2XbvOIjLhtSxXYU+DbFwdTGxcKYd2vPjArBbT6uk5PQMZto2wpcQGKmWcTUMAQqy
sWNSLCUcmnzJO89L+xetX5W9whcA4dXZEbrh8VRNwrvCwLLEDJqU4tFbAVg3GqGl
Z7dy7L6yHE0jIZGfxankfOFgDDdGgPIBk5TaIr5nSACQGNrcrrJrRXQPTPGa8t7l
7UohqWWCOoJ3Wy4hvePWjADB/MnLivjQtfdKxv1ILk7gO3cbFzx+Ib/VnfmATn8/
BJkPZY1gwrW3wjZFBTJ/8ZUXUX2RGfdwSX5b384PDAroN/x0tKDJdJKmzJ0ATF9A
6aUoYTPrUDb7X/F90i2NEW41WnjEJHRZrH0cEHu1qZ/vsKfAQ3GoFuZI9ekEjmkN
0AGeIS5QqYsZ+Be4EYtnQsX+QhBuzDDGgXpPWHLYtLprXpGQZHimQIYBqu4pgSdf
pKEz2xFz7G29AaNXi3Vs6J7XKyHfcD1u4VRnnDDSOvdzgqUwjXlTij4+puUoZJfg
ldT1Ljg4a4m9W64JwBuB8M5kMuuLVBYULKyoeJmlqlp0i5vFC3d/uguUMgdSsCC0
RGJyHPqSgNWSMAXYdX3QlvNRXMRhelyvi3uCufuLBL/TkSXwaeZWgdxmS1I39wuM
MwhgI23bYjNYBSsOR+N6Ov0U7h2+yL0sls2BKvhuyWTDYYMZANyZWuk/FgcBX34J
xww/AHPZbN5l7sfUZpO3w5eJAof4Kqs9QtI95MSPtvutHPxHPLwZ+wlYemO9CU+P
xzWATOh+L0MGM0BxEPv2h+PnuXbh5bSWzG5IfNWALlmAYG7xOrVvKk1UuhEKhjr+
9KnHvv3iGAT9ciqu5IafwwEK8NHJSlH1/ceqSkdwTSoYZMNVSYmFQRZwMgdGBjuz
iLf4DLGdBv3GxqTiZ+kpc0n/EVlqWpg/7ZINKcZzgGx/hERMmRI80tmY6VDdTz46
53whG2KxCg3bsjfyQTNs+8a9dF1mBeY6z9jNUWXem9haJP+QGYb+PNr+wd86aHlV
+EUk3EAmQgLd20Pe6TtGtB7COPSEuK28j8cII82Ae4p6H3Y2NCE27vYctjo1Agky
WAuOrWuiUuSECwEQG8ZcITqnx8/KNmCIGLaHuii6cXcg5qMds8k+sY5p9RdWzaCH
RCZ1S1zjqL5bIj/l1gvxZB2dCTfhyfjjCFuSCnOtU1eZPOf9GtY8xXCWPrzdPm10
pYavgEBVbN7/g4kHH45WxZVIQLe+ICr0rr+LafR2KsWFEV820TK+cnq+OOaZ9Nkv
B2D4Yz2+GttUPmsjwyrN+BHyQlInSZOleauCS00olJTB0Fk/hB9dKA9+izXzU98N
ldRKlEgkTWPD148ia9w/JBcBN1cYTcJXZ8cVRBkRsnIdD9VmB+4Vk4ehh0twsmny
Wrxj8yHObKY0cQHxgnUVQVNExgJHC5hSm7kJXz/42QKw0QX0JdB0UMFVRYEE0DbY
I4hnmdKWGQkYNXX+E+Y+NdTYcvLESNuTYcBl8rAE8UOisjmZS/km+9i7Mosx5Xui
5dRlrApcxM4+8cMNuzu2cPVsdZgFYQpFtsnwUaVhnk7cs8ZQcPTY7DYjTe26Fq7I
W1c6xvWYxyH+gpgWxO8CGpdmahH5VQRVftS6p0HhRh3cJpK3BtdSFCXoFEPfJZ2m
BSAvtFt/HMfkWDuvSu0blX+pEDhLYrmT6GPrrbQd7dT2Jb5M57F1XNvuyhzFCzcE
aHQbWDsV6bmucT+RMICGh8wFut3qmF2Fyf47f1AC+n7yJHqtigRUWxsOoJXUEjYs
MykHGVdxsctLZpe0Nl19aOpAFftWmK8clp2SvW67t4JI02heBrxPQC41FTg1zDAa
HQd3DohhWdk6NXZA98gGTfRy8V8iWCXyYakP8nwK0hgaHdKneuYHkI/oEpunJThd
TgnrKP0OY13zcVLBpD9a3HjTXjV1wptDvJvIZGYZBm/Iv5wal9T8kAjDs9Iv8+/H
vwPLDO2vLmmRIYWuWwXoXihrxyyK28eYUeOf6sj0pCBL4h8393AJZFQDcXXUpXni
0oIFWROJWFLSMqhKlfeyJG4/5cUQ6kdGXJMOXwC2LDA0LKpzB8nCD+SqOhwnfl0a
Xhpr52GBvL4nSoEga/8EEVKEMz0B/56XiXqBWt//XEeIgZNjUQvISpWZpEi1dHeC
k/wWxLAARPKOuRSXSyP2Z5Fy45FkOvEN5Cgga+uPef61Q99ayUIzBpBatZc0eOty
3qfSQALAldrpLmTzUEk3wB6ss2Bmt/zA7crJQJuezxM6cwxD0+fikj+jyUU75loo
EYypQqjmklF+JZkW6B5WY/Fd6Hnc00bnDMSPz0o6yQz6NAP7lgEc5Vlm9haLoYWn
7XQtYrDY+1Lh169Ad67+6ZEWSuZqLeB5HOOAmYWGRvp4IIw2/hzUg0354iPPpgq4
yMOYGRAlGJow9z5LoAxAykp18ZJeJs10Tcn5x9z50Et/EuJ62xXMqn/Nwd+moj+O
wPT9xi6c+R0QWHVHcRkKpEwTRjZiTpwxDXuR9qjwtoaZuEhlXi6A4bNiINIP+zRs
HzqaBqgD8i3x8XiGBCVV9hil0+g1DwbNXdVacQo3Vyj5lDnoeCbm9G3mxkyo0hT6
z+FNLnFsJHeyO3t1TDct2fhxuwxlmIS5452pdrEU1n9hLGWuoQl/EaGE4enYBhP3
ovp2929hFHGX3zIYl7sEoXnLVUPwX9OYmZGUQn/IOOA62c8UkoDd8pBFQVKt0VxC
Xm3POBsMS/C9wajE00zXwOY2wblC5GpHCsHb8Q0zfvVTf8NBglaPZG3KCIESWnFL
zvQCVGOCqdmdnBIlN2Bm/coo3BerIEC7gxR0s7jdfuBzrfINRdyDT+h81b1vwTYK
ecN6xcYRBXMRfuzmztTXRR4S070xAe9aSecmm2usDTJh7ESkLAtK1NM3J7Tl0Jft
om4WLp22/boS/B/jUzl2fcXYKn334m9HAahLjknx0ESqsVkfdBDgY5jrj1A6DJYw
uJC4dRXAEdsb+PjQ0jpuVIS0gJY/LDvvph7VpFie8BaKGSF9KCFMkK4pKf8wxjE7
TPzJJJZViZwHE5yZrUn57QiOpYeSakrAi2AIHGlb6UmjzH+xqrCqgrpcG1ZmyTeK
+ViOHMotJ2P6dOkKYVq+bFgjCoyHSOzOAT7XB/oPZlhYs/mS8xlji114YbsuoGpE
vyoa4XcPaioo3RowzV20Q++6Qt4lE9pMLGjxsAC0+ea3dIlD9Ofn36r7xhChj+nZ
RBkdvPByDSeL/WlP+PGG8dwFwUP0VI9KDP65rmjQ5WXcHfGPEIw3u+Rx+QTGpdkv
DTzPcJgOvR9FeXiJ5pjklrdGqzlygbeDdqv4B4+YNcr1GhcEMgVWG5SPIFy04/1m
whyS1wz7JxJnCWvviA4dJS5U8gd+8vcuo9VbGzyppzqa/40RA/oZb4ErBjWc6y//
H+FFehkmpA13v9CaKIjTqlvLQx1eY0yd/oOLQCtCVQGrrMDEcnbEuH5ZcNY3pofD
LyGUbiRhnA//GsewKqvjuN/q2ekfaqIbaeMm3LFL/ZexNU/hEq/9xlaPFGJYI8Uf
WRt/Lag+cfMO7Gzrdh3TXgcjOUv2u8eU4E+lb4VGCnzHVCvMDHKk3XjQQ3vOpb1R
yK17++sX5jFNuUNcVNOW2w6Qgf4VmRIaHT0rtIPxeWkgtSOReBm3Yr+CPoR+WUWP
K16K+4L08Xsy5HYIqwvNacO5DFyrpq95mpsfOXY3vKSGMq+kvVl4KgcqaawZLzmo
MN8ilPpjJXsw11nUU2+nFGh1+mJ1/N0eOWff718YCOplrDV+qY59ArEjNKVSqDJ9
deIRGCya3bosyGpN4RfaXp0mj19u6WAsZ9+YNhGffHA1sXKANMnGzBu9QSYro6GH
BehsM8H8RfYfD+A71mBCoz160A6bXGcOSDD4U3wnjYQE0HZWxH/KDQiDKRGb/Kmm
OylNklyLKzeDWAOrh7FfxmG8n8c5ujUi9hN2QB1hQ2HDqNes0acgFrJpfGTGQ/V6
xx1KQoWOsTMR4FEQXLLoHyVJYHyOhJRXf5CSH7vM+F+CwdKs0FwfPoT6Men6NELQ
dKH5NYeaNV/D8mYpjMqIVZq5nGcLQ8xv72XgO6LJ8cY5qQCbDJ1gnWterFWYiWDC
IDb0Y9XwlaSEIswPYZcKKufejzoVA7KJvg35XtHY1JEy8/11RbxPbh/e48r3I6c2
9yAep+AEy17/RkI1ZPdZY4ZYgJBsuuy+jAxGBm8kwpaTOMHaEz7zZUguf1nd3Er6
sQi2q/3eCPmF1adBizb+vkpwbxhE5XzTo6CtFSiVSLD4bRlcxW1q7om30dV1oLh5
7FpzQiFzAB7tILwAg7EAkOne6HBPYVP/kE0MlUXvAgeWkBpc51ZKsmuB1D7JG0+8
4uKJTtVo6EpW3FGCCkao8stZAlWPun/PGDyxPNHP14ANBVggIoe9wzQfZAoiH60a
AOq8GyWl+rkWbjaMp5LQqhyF0F2KcWrUAxc01a33JdsorCFMwDALL2SDTaOLvU0j
kvGeVtTA62buG0r67+5zBxZJuMNXwy7PuTiTiQ2VOVFSpAwelDLcRft/7qUt2lFi
NGR8oxPGeAF43o4/cKGWbdKZQ4xSBjEitc0cb9m2CQGHbMnCqrL3Jxn/bxfBebD4
XkMAzKuV2HM8jsJqWl74xTBZIkdGXBAFlmjZ3aSKihu47ey0C7aM0X+Aw8i7xikE
e45dfr0I2bvm5peCBeJYyh5EmVEMXR8gGPqOud4cIRxx02alSAFkIruOugrufB6y
3WtYMYwH19DVqlnsR80A/PKItUwiQvEfzv58aHddU3ZtKfVsfMJXC5Qed6yqotYb
dcmiJ3jaRfSQ6wu79//vEpev3tbPjUpnFQ4+RuJ8WEQBvPcjgHhJKFLoPT0w+KjQ
r2Qj0H7AkG1iA1IHDffjpSenTCUfvlOLMt4qYqqulw+JoX98PJfPAah8G5GHzdWI
UATETThKeqz15OGrGcU17/+KxyRoJq21igJAx8/2vNSM3AhO5Q4LshDzP/MoOuhn
CQt4KuSkJScaCLsP2JPYapHnQTj63FGNZlGRT4zCBARsLsLHUiQhEEw5WwvS9fw+
hnPBxlOKMgiVaWCQpPfPZjGAVifWzhHXj9AmAwqXeqUx9ABhe8nE9DSbdkHUREjV
Y/AWb0JLnGoppiITJlk+v1bTLhENCuqyzqjUuajcjGU3NUWdCDM9/4MrdMfq5wPQ
v1t7Rx2q8sc0yd5vVc9kj/URYlsYkl7j9BpyyFcfrYCvodFesvaggQSej6l1VBI5
FHcQWu2/PaNQm0v+g0CrqjfrlhRrisAEBmH8pWIRL+KOKrMOulFvL6GhXB6pjvAE
TYG5ptErWC1AMTFAFb3/ptXPh2B9NXGu/eeL+fejUvKeaFpx+plFGl6ji6TOOagc
sg9qqNE2laWRe0uGryAIr0dFu4z0NRogqZSTwgxSPrfC871uzGg4t+SrhvYeYv8Y
xqJhK3/t7unDmeg9BwZ6Yxh2t7ccz6+VGJ05R8jPLMJG5Frkqr1PcxDvDS3U/oc2
KJa6JC9rqwYWMqEtVCvWTpN6jEXhlyWk35PypIgofVdYcekAAV4asJm3rePqnuWI
AdiI0vtpDxVJrBfcJgXGOSDjVxZCRKrLIBcVS5fRiejznD1KiS8d74oSOd24i6Os
lZv0XnIqHpnTmHEvRJMlgnFyuVqBFgW5JtqaEL7YotbrjykG4QWKTIyKN1F7DkAH
xvQMoXZ5pq+3+/nU4p96wCQ62VtQFZc6l3lmlGL3cE5h7zDlr04t3+PZuaKeCIbD
PH1hVPL5A+oI3SDGBnRPPkqb90iSsqoXw60qPMZaWBKDletmpg7owPYuTkAsUjB7
6lMgb4zWyuYV0/hy6athqQ4iLcPprujDN4Y82yKBi0j3AwW03k4rJ0E0PrRixDb8
8CaJ+zjIZXIPh3ji4NFR22GdBdMpueppSHa4mjzMb/A2QCkrpY7PtrVNmSQDdzJ2
SZmLrBaNUn7xXewsqbol9749QBL5eSoGCVKbdQltmtzvzFnz4rUMmPCKCejkuqlP
ZDi2b5sHCmiRpixqiGc0SehMtSQA33/l16IaIb8SOQ4O4JFVEAw3kvTct7nPJdbG
8XXICg217d998SYjy8lWfC2adSRq7vSSN5GL2o8Gmk+cm97aUyEPnJjjwKpVoCth
ZI4lVgAGR5yeY/Ab5xeaWundKCDKXQhBX994Fk7uRiE5jQqnSeXBFxeUGmwSgTRV
c1m9cTCP95Ujqmoy4A3TXh3/vrgMbH3Cx9toxba42zBoTT+7Sx9hvYdirWBe3ENX
OQRMAaHPjRicHCz56cDtO6bXAhTH/0sCaduUel3HHI7KsDMcN2JLvYT5VLkZxpOG
rs1alIm9aV4gJcVK5TRd9JqaqPMKlXbwvuqAJjiXiF7zlEseXaxWlKr3PYuF97y7
Mxctg2InJ4GfGVK/W3atF7MGSvuV4jA5ZhwmGZC7hdhEd99OZ3ODrf9CzNRlpN88
Eitf5fhx+OZDPBdpZHUdfmPWB5tpy2DRxX/kqX4v+8XsHZVujHFnhi24GXwnMXZL
70wqbuFaeo7qVcFwpLmxC4vBcg5//vH5pC44712w+0YMeQB1QjsYSSYOZVemxDhg
FkBgoHxRlSMXHhmcNlJbw/bMB+2mH2HSYaZTk2rt4FLEsgd1+QG5H+5sLxZGm1qc
w97UZpZnmW13BdA/cPRV3FsIqKjRiSiwQOYJNqhYbkcR54auQ8e2Ubm2xqrN+EOt
D9bQmf0HIaEg64wLZFVdI+lKuTJFJmay0Lk2Wla8q0loBI8zD+fGs4+fq/MuI9yI
mMDRJQT1EvK2lHow4/lRf1KCON31vFTlabBNuq3lNaB/KqY46XuaWNyowerozFxU
zi69gf9G3qaaS+cqXCXh8seMexMIu6/YDU4TDk5ZBzML1DAQLjjtuwqX7mQ8eJo2
qOexgZAd6E53W23uYXdEcMs/pR4UjQ8rmrc0AAo2AZVD++BfYqTSVq362vcsHxBv
o3JT9QTC80uHyBCN+aY1xPa7EJvpNhIVhQw+fFapkVbch082ut8ZplqqOlplUvEx
F/bu36b0mzdX3wFcA3VDB8sUTPSSebEiua0UnwZEZotPh2LkgYWpw7w7qwhlcqHm
BWMPwSHRtcMJulzJjBrfWMghhIxtHcuubhyBHtPUNhVm2NhMnMzyGkUrsPxb8lZ8
o8GrMHLizhmfEkg3OyL7aecWQBXbj8Slk6wUhoZ78p4HU53/WsHspcnIfezQ7NMh
b1nrt4+rZkwJ6zmiulObFiRc3Pkc57ylBlnGS4HZCyZNI6WT+BgAfDQQbv91sRma
1jb7iDknfUYqzuhrg/fXL5t6uQKCPUqLCZkbkVxOPSa76MxJWLCEdJtkMg5WBSyt
CyLclWy+NtOlDk01DGqBups41PNYE/XE/vdK2oLVdc3SLgH6hcGfhCX/CPyhIV0b
4kxeMcRzmkliaIPZDrUonGx3fD8KZjWgjxXHxvTsJ3No5JagZ6KANdDZn9wZOgRU
PAKLQOa88ucw0vttWKbs75aOc+GqznZUkl/v3FPB9BE0fh4Anf1iZFWc5blqDtGy
3yz3z3p/fMjAm5fGY3HnFAudx/t2MQE2i0bBgHPG7XxfNL5g4zSG0JAZxFCSRWEO
Jd6gJ1SMd/VJpAjIXPSl6csjyAillgEPdBe4ADkhpAknXsWX6VrBGxefZLaWccC0
qHgVHdttVxB4up9cDsnO9U5f2RPZJiFQmCiC9HUiTPUxJOQf0Z1l0csC1C3QJalg
m/2kqu7rn1gW5AyJO/2z8ELzSMtTp51nH9ejW2D7tb40hMfKzLr+xEJ0LfIpMDt2
HMH1DqfWuI+vYzaKgmy0zxQjT6RHh4gv2XXmfPksR4ZSeXNNvNZwJqc7mzUkLuq4
38AxSrY6iNwsuYf26GSdRvoCHhZHP2XSjyGe/cBK+tA7TC1rAZxzI1SU1tidzrhE
zI7atVSM38x+iNOnUegYW4Gc1pXmfEylJ5yYdpVk6sGIiDHYODEdN/S3lO/e0pH9
AINoyxjCprRhUtqDFf6dkApN+RB4A/Bn+xri+7xQNostgezjHNjTa1vhvawOZr9Y
LM+cp2iBZ7Y7FQxcUJiM57em60Gvy1B9tILWYIxZutNE5VZruXywnWShmfsNtW5F
ZPDnP8Be/xz3gZ3z2Qz1/a+67FbJF5MhOGYU4NOF6T456GFqJrGAH6uw6C8iRcFl
XreFpH7Y2dJQOv1eJAD+0SxSf87kI0ZjwIABcVhNCzocbMxRym3gxhr/w23qObMG
vmtq34siGTZIC9Klb6j54WopArmnGRaQdFFL222z9hrpdGt/ee9thYdGJPn9vUPl
MwGWqVKOfwk0llEqaga78uYEH3t1p5dqkBC2KjTCuhJXXJANx8y6RwJk+h27s4x7
CzPeuVWYJhczdmipZOv9/jKHJKi68/WZRyIQJVyMc4CgSxtMIh8XzLrjKp2LJQ5z
uA7BGu9wIP7KE77bzCEYBg2fhAxUvxqo71uXxHjiPjam+9S35TN2NbsODELEqpy6
KEtE29YfIKUWz+wFTXXdQTSAB+arOAEmGkVke2qYb7wOZf8BUd0JYT4uA3EqAlJL
PMrmhp6cG/BUK4fmnyVqpLIqmGX7ltae4WK/rBwM1EtQkRucQ1kZJVUjnVW+4x2/
2Jsozj/hLLOgiBupak3YDDGOyC8ERjWiV3pDoSpZyfzhAKiXX6KCI0qBHhy6y4jA
YhUVFHbbvR8Pn7s0rErlYedFpLWl6XC6dxlVp8JCRD+K8mUK4SM9KJs/qsl0JkOM
Kj2+YmQdEzktGlIQZHBiY2Kh4kBymjqlGmxgFehEZ41Rabr7hhNY0vW878P/1c6e
0Xj2iNqZNninPFrhMcak2FRclQhaE2EZ7Yl+/VBBAEoCHA2rAaLhmtdiH46X5bro
HoKNbzmDae422MzRq/2QaB1k3jkAFYvipJmgtcx5yimrS4aTERXOOEm9sLuHwEkR
zXoxYt8DBQ7yLCxkOggXkQpEN0QZrgU2ourbmqMZSnWy28bbXerIAqFL028Rbg3h
Ql1opaW4qKF84qcTufcHgtI8+hEG5W8EdyK+1CX5DDdKIq4dSIa6zNmDTyuMZWpY
vQA5iTr23kfhSTr8RmRln7X6kMXLyF/iGntfU5Pv4FqsrzFWH7/z5BO+7Zf0azXo
hwkxQWRwOOytwYz7INgelwjlk/wGShQGvERsr27gm3rF9d2ZIxdje2bQy8RFuy5B
DzP9+gKNalm4vlF4oeddXFGwD8/Ki5SXQMdbPcew7ANplFkrzTwxdcwA0Bj8e6Kx
/6KtgS2N++2s7nmXtEYBqKtJYMj5oITikV11HByWVm6P2xGPTuxhhAk6IrJRgpyK
uyO4IFA/4M4Ta6+fZw+uiv+IvpZSYTsmZPgPSV5ATWclg03waYEZ2pfxmY+/P909
5GNVkoe55hL+GV4CMgQo1jzur7+YoRSL7Szsbtl8eohh29MFpH0t/W3bjVDTYnGy
3CGjKo4bRDk2OUdi1qqjs+zD/+4aIaYJe6QGh69wnDdruOi1CsV/OAaV1SkEPHqu
Y7hDhPpPRhNEa6yhtId6ASF1RP1oFryS1XmIkbeZ15eDc6pXWgIMP+wl/J1qtkB7
Wl9769Ik30GcOXuHAInvohu9vyvdo+wDmxFeQmZh6ZI6hBOG3oArGnB+tK7Bh6Wm
T117S3U1btCY9GhXaKEQPvbGAz6hqptRu22Qh2vWRnYsRgCg3toS/Yh7K+UmVRsf
Sc5KSRAtUOXGALDQzwg4I2jDv2d+bc0sciGK7V8tuOOqAWhuJh1fgHkEAdVgbvvd
HRPO03fmYumziUyZ8Il70fR3qSjIvKBbuzp/SmwSfCJSeue2dfonNySOUOWExieT
BEGytuV6IS2TPERUZcmj37iphgdAy54SjW6vrjHMvWK6DPTiVxB7WAMPD2bPhxAh
qaDVrA7AVdMzn2jnMaFUyTYlA4m4bGYd0fTXqazLW3gGq0ky7OvwbL54tkV/1JEN
XWJvkX0zjKukJBAjLIV4aVx3a6mkw4OmGCbFpXoTlQtE1j2GNqsC2aoDRHefSIkx
IqE4gLiJqH2+A+MCBJUPxcztDJOEo3KXCq++ZTT/tpgajaUmov9UHLafGeeBUgQ0
pIKVvLvEe78w3rMzkjM+pq2sJTky+41ibiQTfUn+meDJaR16nF5qTilr5YwwKhjc
6MQJT99+zJYT9nz54BSQ+NMY86I+3rGCGMBptKjYpeu49UDCpqIpH7aFWhUSs6sS
WI++XnQhEoF5vbEbRIcxAHp3iboyMGGgFHtQgQcT9z51Y82nQyRV9OqgshHvm5kz
+Wkkpm5rRi28bPcd9WS7VZ+Km//YxwKyrtaFT5QtZJuLRsws33JyV8eKhEkxYXZ+
z9EjLwbLb/yX5+BDj6uCDIBr4cL+xMlqmIx/xZJv55UNO6FF3vuQ0q76hRa0kYca
Z6oxuew0bYLtelxN2jQqgLTfE8myoosvY49HpeDU+gpwHDXH/BjsQUDFHlU+I7zq
ftLnzMH2+jYMoKcfRcG2xMLOmXuIGYIy4aqE5VjK8I5/iTQ9LxVc+jPBCE/XASqR
2yY5VV2arktSw/mJjl9xdGDhVDQx7gcoI7d+uioC+n0yfnJBW6fYjGOMXojmpyzl
AjJIovU8aZnUQbqv3RXsmAxcTSlWYO2oRXBw3DlfTUoLP+zQZOmmDmhqXYH51sXE
fOWjBJbWYKZtIyKmRSYZpl5L9rxVBS5aOhoTw925te03qUHjrsOPqd7P/6+TGwe2
MHFCNZlMSgzfyWYFHrIjGUKs08lWcxphJUw5sqF1x2t5rObS4rd/oCmzn8OX5C3f
h2vUYil4tHFJrotN+8kKZzM3/97T6xByLziE9HbJifJyY+aGhl+H0eFOnqSyaKmw
42VbfKPwdivm5MPREFGb3WJjiKn6ETxH9EWs6XxB3vjzjjJlYlY0FUjgACWxiOZw
rNZoor0x6H8txKq4MD0KmW1sxEo6BKlFz4zPFiJlW10olnXwIpsbko0bjRXDS0/C
9PqK1Ytyute7kshHDbAzYw7aK6VUhUNEutyUsufuPpIp8tNUVSeDAVNdpj6rNbz1
TyaJ3LjaD+IkmUGmB53omEwz4QghRtSEndKqMb10kKKTa3cK4R7faTaWV0nd6jJ0
c/0by6Pe+ZMiZQla0VANW3/f5lVufwCGSP3hgtSruESq75KC7hzFPGSJIozxTTVJ
b7S9GP/ewioQrjGAYKgQ9sAyYaT550FUHhpv3iCE4Ro+lRpi+20FSNbAIsuYz6U5
TGXk0vu8NAX4qkb83ZjCeSII9Pj8x2PbwsVoiU6dbxifei2b2AXb3iD0d0kswU37
UI9Clk9z0V2JTB0SdtOyb12SIo/1HSYWBC0UHlLCvqkJyDWxWdSFV4OAAKz/+yAO
Kj+FyQ3it6fUaK5vOpPjrQam7TS94h6yknzZCih4H2yHXfD0eno7yDDo0uG+Kttn
B/7egYtqSJbT78Je/f7Csf7nY9CjtNi4Srjjw1vMNcUR2w8WwsZRGlcXbcHQPbbc
vD4olIRuxud/DxJ5950l6z+bjXLkOHc1lafmfLCM+nipHFazz44w0xDJ1akGH7qy
sw8fZJk//BCGHkaFdHBj5hcByEJG34HzQ7+LxugFRG2jMW8242imWeHzdo+yE4uO
eArZ/3ffkxcvCXJ7d1CbOaxEYf77i97WYmJk06Tvb0XtH5fKv5hCNmg2N2LOjrKX
W9g3nP7WgRhTU4uekEYHPTKfVRQYBMiWlLt/mhAReGP6tBqyRaxdbwEqz25un45s
YGGqXeBmmRK4zgeyDU+fBIuzVsAYqdqWNZHgGN8v0cg=
`pragma protect end_protected
