// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:02:09 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
pSQw2hsoaQLC45eDmAaj6x2dablIC2MgeueZuIRIy2n7vxEmhgCHGVhyPm9IvPoI
EfQJgdVaTIc2RFLaLq272WZd8BkhMg373okBdEbRn7utaxrokK28wnbVUjZ/WFa1
OZOY5XETBvUJ8+GvTF+yUplPiryWd5PI39n/K39WsmM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 12448)
xWbr+z3NRk/UmrjSHakhrSoq2rEyuuuEUB75apUMYPRPOc2pRlXehLybYEEKVSrQ
DBuwpkTHrqDKyKKG5DKuwqipMF5hOwaYZ1t9atSwE28fMVJgNkzGCNmla85hY8hl
g3/ny9dqYXYHWYwVLbetDYSLUMm2zNOnhlGU2PKZdVdhhy8G85fjDqdazJqy84zV
2MND28ddhCal6GT3ka0NxvDtkLiKgpgAo0h7zH7jm/+HXIFKdIV59JYDXiSX+XJp
RP1I6d1zB4O7xOojvi7PI6KuJOLdg5SWMX577Rb/zUxEt4KJb4FiNPj9+nIuNvQm
NcE4Oa2PZ559eZoKWbo1ui8DvlcXx+2VoK0LZJwe5HSi0cpNCOo2YBCYv3u9hR3y
QGZqRawGvOj8c9790E0YvnYeniyQnEOGP3wwoo1iLqZwM+u0SjxpzMGtFoYweZk1
Glhxm+8AH73GrK0Q3Za5PgjCBVY7aqNbJaxoUqY3f5Yxs5bmpawoQ5UEPjvdlM30
9XgvPM3j9n1h6UCzB8KiZLEUEK9FY9gM1OBAfrDoYIQFXY2phiBDWH4yFANNtMgE
+5iY04GF7/DDrZ1SwnUsFzXAPq2D+R+cVvuAEhQwoMKKKO1nk1tgNL8SztGaAWVG
Wvv4CO2jyCgHNzPc5JLcaSNUtv6RQJxJQY26v+wFtTyWSBvmeMrfzmmAHvXnttlC
imTmFztrjFS7N1Mv+6RXBX+hYuIJwGhxTiiBb4oWkSBzdno2mpkMcI97GJBsukfb
aqns78WTO69rYh+W7kUq0wHS4oyZ8b1YX9lmjWgx2UTjig62CHLb/juFpGmMIS/H
vDKsiaF2CE/6iyOZG7IomNND7NlpK/yZnC+Df8tF3dc1MH+W23QUQ8rXdbj5iHZ1
ZNyz9M24rr66IhHGP5AT8YpLX4IXKYJ4WCsN5u7sjYSinQkNC+/x/AZCWXXRi7eb
FaibCDlRrupLGHipkxRJLg5/yEcIKrDfFXK+4hFlzoLI7hTGIKlWu3xHp+jSDmPV
Vtj9etYMMDBqVz5hN63KuIzqLEKQB/A9MXybJSq7ORG/Hy5gksLuzm33zCxDCGn8
69lvnMxSAB+EaiaeC7DbYjpiiGnpl9WuvDB1G4+Ru87lxvOADDtZU0lv7Z33XpTO
9Pp0GaOi/+H9HuookndZyb9UtFsUoXzw8wBzyDZ7YyQ1ZwiyR5z6EmDNmXFhquGG
jyPkPLvuxDSKKZ2MLNs/OZn4A07m7kYluN1VSBiT+IT078CfSBJAPeO+gjC5z4sT
AJGzbRTrVhiO+bssQEXg8oTr5gOgCLn0UOSAn10AJvsgHgFiNSNTPXizsxaG8aoH
VkBnGPhrJPflxMuUOhVg7r0tWz+Hx2LG7N4VZ/yxQVFQIdUvrxT3M7VHZ53Ekk19
OID/sKyOF9e8TL+RaNYLcwh/KnLdY8cgL7DntQymg3ydy/qnQsX2twdIByJZSzBI
hpUKV998y7OVLa//ZseetoS+su7fNaYcggf+Tk/saiGaMrqJlj3yUmRJZ42H9DzP
7rjDeQHoeV41qQUuYnehU6B9JtNfgEIPe0ew493zx9zCnnP6K5P/zU+vObvcYnCV
79ZqDsO9naroYjODIBXq+gHln+VEIR57jwJQsOeZFfsXOHwHEH+uSiTj1SG1J5eD
nN1rfW1Qr7HWUrDHnQ6fvZDp7hePQZd5yA2+l1BGsNVN9x70PKt4cK4T+F83NqT+
KcNbrL7bIrW8jBKhrXowB3ZF0wKbqtefjiCBb+DxaeA3txNH1Fs8lbP7Z1SFVW27
zqgT0ToclJvA4p6KPzSMWMVf4MNEcj+O/53CWqW8/nYsAlmvnOhfdMxnR7F0UU4I
kdxQOMy8iQBgCDsC+GqRDdtHdevTMT/V2nZ3C1cdJZiNJ/oub1nQXgrvNFCARRob
IdIvar9Q6rJdxkelFC7+DB+C3PWZzneYtu4oUZ8lm7vF9AyGA2Ou+YpqAl3waUDU
AScV3Rja7bZTuyYyu104aqNpAyxC7PNwQX+6XHfnPfM8HGhhH8SCoyZFRUPyGJ6k
riWqga1jlUdSZjQtctoUk0xGUaLlGIsFR9Hs8w2MMw2azvmxNiEskN5MHwHlsaw0
SlA2oohmrjU2kJvQCWOL//QuxL1oGbhpxa6hwnMjIJRvdOuYYfZ8bFniWmazF7ex
P9/vS1CcwlbcD0WWkHbAgU1AdZ2zzGoYIGsZQIEbeG6HiRPW4z4pDb5/iiE6BdNx
FQuCvH2EIOSydzQWKvy0vsJvm/bTqPkkKIS1f4nK/4q9Lj8/Qqzbt6NhHF1eKyY4
XrSNCaALQDfjapMh7bFUH352p6ZjRXu1cHVQwYP342C7bUMQzztkJkxs3jYCFiaS
ykSGV/FKC1RLZ5rlCsXk1Fnb2lNtib+pkLc9aCCesVOxL+9GBRQSmnAwiUWZTTRO
ej93zmlnb/JKw/ioqzUq9iNviOdyHE3GXe0e5GCj09D5cNm5Y0W23lF/W0NJxzLn
WuzfPY1akLgzPvzMzq7lFmuKuqopR7ysz6+0azI4V3Tr5IPnEEZAaHodZ0AZ0SQ4
FDkLasO3UifkOq9Hx2rUpvDNOiuD+gBWbZKSltN7YeiNbOFGRkBRaBLZbJfyavXz
ZAmlm7sL5g0X9ILALq0NKv4QlY2SLWmlSSXO4LjMo76EWVe9j5XL0ieANPEvbqp/
bJLRBC3SVPgOqvmZCViD5nloGkdrVQrzNHJ5xPumkwWZJykbEoXY7BdLU1iUL/oU
+Zs9IH1Lt7F+BsNOBIGJiP/TTedoBQrOlnrGKNtMKtX7vJxIbZADuUCkSVOn2qBs
T6c4P0sqoxIVa5aNqB+Qkl4gxtQ2K6knNTuIoFYdc0fCXIGJ8JhOiIHjL+QRIQy6
O+eNHIabc9bhutoC9BYco6lS98TaCK29+WX0fDF3fIinJ6CpPWqVl5aHe39qIunS
zKOhkyd10pmeSYeC65dYv+KEmCadnHftyrs7vyD3NWzj8di8CKhCG+c2yKZuW/2b
11/sldG1reZnqjjblCSLslsk0/dqHe6ztyc9Kca32BjmSDbTVHXCnklH+r47v3IE
rosTLNgkr2QwTE70DaulILhocnuPcOwOiTi81VCSa9n19+hCPIwO5pgpQdfqDImn
bIoPhMbT7PwdgaS+nLHUHxFwwLEJKKaiGVa/gr3CstI+xAJfEcLsUmcoyWY+4ru6
fj4Rq8ndF3HCGq/OsUh0OfsfC66U00uAWjlEs8MDLOlMwRxd/N3fzZMwRBnNdp2H
Om/WsZtPcuFtqHWAjwsErseUKmCafQ6kdVx0Wj7bx2d/oDyWPiSgWpppswDrxA7f
K4B91SWfw9HYqFaClrWojrikXEcdEImxP1A5hQ/50XJdFKiTI7xShtQY3q7ikeW5
Xddc5OkudWHhvKoPteCH0LApFecAE5U/yxZT2ZZIJ4yCw2lUYb8MGO41rdOfH15t
+VuBTN/pS4qS5+LoIB9BMacygUafhFk6jEYBMbrzgXfK4fRIAJwyzmfGg/K68nAW
TyelKfJQKaLYsD5uo7Yt39jqOPBL2L9tfifdT2P6PmP5/BABTzvgjQeHAgapBqG8
XYZo10rH+rNLte0B8aJcJtkrN61BWeMSpqFRk2qZvh1YH9szjvop8nKGkwS3nQHA
5DNJecEpRqqRB8V8R887Azaok7GPDwSlGUJMowMw4GcYtBJX81ZEuTLOxVzdapJP
B657bW0av4knFs0ot7hHi8YajRVxkctpqZRO9rRTckuav6Oggp06kaH0f+mYRxjd
Or7LmBL6UsHeip6tj0A93a9qsRYjIiDOslCuZ+a8tTxNmu8arXMst6TDlpeX+9hD
Aoz9u2dtkpElnj370KWVot+CQ6EJLq9Xbem5Ig4Em6/sFl2gi5i10Ag8orEkLs+w
UtunKmFAIy908LhQH6WmznBShPwqk97UMX4mNp1Otpvx9QJETPLDG1dB6CIdnZPk
/f/dLW/vR4zrj+35SmOXO5fDQtuRz8O0g3cOTdQIXMr/sYzQUMIoZ+z67J2dDt5o
5t0Z7elW/mRFp8QBSAsmpFORQDCre0nB8Z+2AsIVQ80kod50H180rwsKD8C1GM0P
0DlaCQawS6O+/478SWuOMY83s0l+VLNdgfx3SKMcpzqvJCOcFVH2E71UccGCKdLB
Nob7unWo9b6buzHApLj9Ldb+5cK+51bizeHoqKmMRcEl/yv5yZ57jl7UZtg2z7w4
wepJwVxYAc4rSx3Wv99EQs8ALODyKW1yd3gEby6rgBapa2CiYq1lgq5mze6KIEcM
bZ5gtA1uQgZjvt9a/cahS9S+AI93M4ozLJchYZklHhQ8PqhnJw5dL9EXBx3sq6gR
xzV7CrBSdHr8FjZbvX1/upVeADrwpsGEfIR5Fs2hQFxyhmz6gnyfzqfi0XBW2ylJ
rbqZjpIaM44ye68nfXDIRhGPPZT1Ha2IuYFR90NJ/rPZ8QX2oGdSiKGSqvLQSWHq
akTPrDPq85WozfBPVDxHknTzuyPN/qSFi5Xyr583xnp9MFNrAm5eeZEmLKnsRl5w
F0Pi+S3ZGZ2ADKzkZaPnxcwTANsfOXKw8RqERxbSEzElyZaJCVbfzUcfwBxqWVyZ
TIWri6kZNwCeQuEmTYKLqtwFaGzsTI4nd45kb3JM1bFf/OBG/VthBXFWNiTgg0EC
tucbFB5CHjgFDEiX9AO4pU4iM8FF9myabZGSeTxy/tVX/3rS1vXEh+qav++KjVAC
2gf7MsPwzqBIay2hSNF5uiXZed+bxiTekQW43sBWFH35qkHHTpj+Z/41alOZ3hHs
7MNH1QmtoaRIlFbnJedeutCXtfRMd7JNbNv8tdj31meVUrx7Y3xtcpuvMno9qFHB
eQp82kBC1woD41KH/mdcUL/QdKNf3k+Bis0xw2DQCXjJPpTNVT2bKm1zzrkp/2Il
9E/aIu92xZRzAocP8RSGyxRiR+AxHGLdki0ujkbaJB48ityrTXP5xlBzwVe+jKB8
wp43ZgYKSJemZh7eO7vNoKCK/K2ygVTZJe38CJszgTnc1dlEexgK6619ZuulIrv/
jVQQvRtaVXXlsEgvm2TotX5PuzOi4+CgS+eVaC1w8Uvg+I9q6cfz3OSXd/HzMGgh
VB5F5yq9TLMGkyxBU24EKIojLaoRccrHSGWV5pS+nCY1by3u7eWOYzaUCvq/VKFK
vPhmsDwpVe4G8GbUHIzvbxrlhWUpQ1nX5vRIpL8TlR3JtG9tLlnHbL49te/Q5TPp
gpbdWfADK3XS7acimNA+5Gc4rp3WnS16DwOfn6+xnos3qCHBFC9mhgX+C5f8LQWx
RMUGLTOxugN/bHEElYNT9ZnMmrAXiNZufNVPfeqsFgmd1k2KSFMbujmJGSc95S89
J25GiMi6reQG4kX04NCzbGiCrHrCefnES98LJby8R+pOPba6EmEjyzN7P7DO9NXM
PFbHFfYGsfsFU72cIBU8JCAAp9kR7XUSFDHrKUJQb9vVh+d5uN8u6X+Zp+kWRBeq
SSop1u4NWJ5uINVcJJkvoDoJIToIm+o1i/mGaYJbaOA/v9qJ3rmEJmUT4bNqrWOc
Lm1htsUl2qZO/Hp9zWeTjV/82AktA+qMuOQEHb3XbNB2/nj7QNDVHYtXhJTqq2LM
ZItu/e9+N5bLAgHF/ujMKWH8vZgBO1InmGhQbCOdaKcPSuIU5PXgpW5qcW7KL+sn
QGTJhbJQ0egR9KgVGas+4kp2lFwaMuRNQ4WqJoB2cAWyHV3qdn/ITBkd3MJzFNzf
K9Q3d738aa5iYMgEDRJ98l/dvfgBw0MWU3Dqf+KckwIIPM3QR5PmEt5m74ZxuL78
aFbdWgySRTK43F+6dkFY1UqVrjeDNEF/vWv90s6N0KN8ap3BB2Kne9DP7z1GLce8
n0rHVGKO/QLi1BKP/xL1q3X+DGLRvhJ4NGX0bYLbamHWnSu5cCY3gsAYY4ZM9QhY
xV0VOc3WS0GPNmcADl+hw+ZdDuhQYTSyDPgyBNfukfgtCCsPeoW2g7WDJfzpWcE7
5e0EvNTcMT2HIDJ10gS3TLVye4I+KWJFRj5hF5468oscNqUaplf2F1WRievZ8nEV
4hkcVokQkgG8QCKadlV8YNQTU0ldTCjOXqPj8/99j2VbAEzKDRUc2Gq5MGAd+2zw
ohIIwVXb/HsPedTnMdtS2/HGj9bV7BnRXu3Zt2wxGRaWJY1yyYr34vx5JcDApy7w
ALy9WmRlbr8Oy2DUbfiGrqGtdoLuAn61umx/09mPUF2QHR0HpCxuF3mC4EKVFTRx
v8fBNIw9PAzravUduNeb9MC2Pp0+9WugYGZiXYZVl6mNZAG/tEVIpwRYSUraGRAJ
MggQ0ZUlA4lapty02mfaas6qSGFlD6Tu2D6yGj52SWNPuVauaK2xVAXo5QIGITEC
a/TTHPuX9lDPpKd9jL2MYAko+4lNTGAy35yyjoI/gRyCE/ACWBrs27bZJGATfcKe
IIyFL7vAkgmXoqBpzuX52BSJ4cJWJaxZaRYO+tp95wnhj9YGfTbQia0zi10VgkI8
5lXiHB6nkMxdFwcg354Gnhg2oOS5a7JI0F3xJ7RAs+D0UNRLYQOyzcAA9PQfjsVx
Rs64/wn04JhnFMUpFZpttZ/QvC0lJsIfDSpBl3NgbFpdn1pluf3yY8+0RYlfMN2S
SlMrPJe0WCyJmzzENv7OXFJHJ663w/BaugMHfMmhpHAtnpiSoQvKt1rC8dQ5LElf
b5DKNqH3WFkwCG14F3wpFSLxwdsiYhKfnTtbroapuv8o/XJxj/5XlpaKDhDzOWrb
qrNVDXV+Hq2+MlCTnlB7ZN8JIpeHCXU6mBOiA53JJhcOMC8J8sB5U3SOto2iu/0B
/TX5c3uCD48CZq3gT4e3g3Mk7gOipglClCTWs4NRorw8ZeZFM66uXp6bDzQ8nYzA
Mqlk4hxo18T1pHU9hSxJn/SibR2jHnVqaMn+b+wqtEHrbnCQ7IjJqREHaBQ/a6ci
MsT12m8Ra7/jY/IvbvUujbky/eMLnqtnP/SU6fmkUdGZUn6XaPaC5c8YigIGdm1J
tCwPu8JvKk0zCAsQKHJXnUiHI0hK3RSmT/p3kg5BFkoQ2GerW5NpnhcI6UHK+3Gg
FanX8mZ47BTpj6vxpbk9/L3N/GSGAy0q1rvfu87vYtA3w326Ws6v8xt0vNDJr0K6
nU1z0Uz8BgTyKBKtvm1O/6q4KKmREYHG0tIeaMyQm3nD/IWS3y0k6bXhw2rSgZD5
DwFCIe79KZpJ8tieOTM900dPZDtd6UYci6Ouar64vyUzj6FJJia99qKI77mrLeCk
i42jw3ghjX4ESt4xxKBaLQkDpRiS7f1qcZ+f13p6NaDHcFPkM3II+uzMWdDegdwU
R2EJYcXaWUWzmWAfyU9+ak0UF8Z++2HWH3PkEfjeQ25PUhPzWQ8V6hZzvGBaiEAe
YJX+qUIb73iim5qEFc48iGogNl41exWvLdcXCh+pkeSz+cVecdiMZix8Oy8zLuFk
Q9uYelDLPs0fFhlKQvubs3ePEV8+eqgGZJMVxsvwjU0glZcB3XYYXPpQPoLmaOBI
anHXh7ri5sueLlJQvSIsHh80m/G1iDD0V2zQ2Z8A69Y80QJVPuxJ0f9BLmJruJBX
hMjBsSnPnR18BEjoXbKSSczlWbaA+3r8nyT0q+Tb5vmvudfiT3JJFPU1LKYIw1gn
DuyoBEEBeR4pxNp9J4SJKEKPKePcIkoxVPuFZbJ9JKEa4iNZu76gH80UgPHC/NK8
CoFbFeRvcXHBLuOTCWXqIDGmHKTywzSpRUJaFlhbBPO0THdhqhYfcBDHnORw95Zp
oyIsLsk5o21QkOnrcAZ5dOBkGoXopudXO8z7cpfwHtrKDncmXglTd7/5cZZBrlyx
Ggefq8DYDHLmB/WsQUe2wVJAdu2WAVp/3/TAf5qJCZbFoGU1QuMCeRTle2G/4vRj
yFjl01aQdhYeuLAO+483YRGFtHg5VgPNCd8jO77tMtBu+C7XfOWmD2hUDXSGn8zC
J1oHZQKrLfOkgpKWMITA5IUdiHMen46tAyNcqEKAIEsfgcYnMFH4NOjX+kwHocpW
LGNJXKBT+2I9FooGb4j1pXvKJgmGVkCoeVHvETZQL92sbwmvnkaELWV5EAvY8eec
60W0/FuJ6g4QTyreRAyjKGXGbsnV12Uc6B+AZiIxz1BXx9WPzn34cn+i7+Rp8CZn
WZz7CkHdmI7uYDPzVhn40AMbBYUeycGjnb7o8HW+WpueA6EcoBqpqs6Kk9NOwdJg
2vQxYe3flQLcMT0l1L+AzRO3QdHjla+wm7ofbqHmKx3sBFTiuRS21LqyHaqJGLUD
gg5VUfRP5GjopbsRCMqfYJVSFsYjkBDmOdqvkXmTcvsNMyFiFUZjVcAa0z7CpC3j
ghZJE4es5B8LO3koxc9HHBDR0+WemEzvCzCjvhgwGgtdsEeQ6KeYqYJXscPPyifG
joYxcTzlaVbdilFcdzOUD9LGV1xydNjdwrvEqPpxGhn3N1fOZYvzarL2H7CmRugJ
OQXVfh++iLR4kT0rJ10hnVs5+MlbtmGAmqLvpblqfDfT5ILh05vQUVt3XEqy7EVu
6y442XexFI6RCFpV//5FIBH9QdaO9P6pdCJm4VOcXRGNh4Bc50+Gqj6vVaPJbVAD
CUqKDQptuUKXcReyxlBhgnZOkJE1TkIMlIh8+Ir8SXbWyMr3UU61XBsiLA0JGPVw
mEdXbekwUH0tJhEUsMfZgR4WK/HWZbqvuthjDO+OW25opy2MUA+PMEL3r8DW17gB
PFXsPz9yY2xzW07EXLoKfTIQui6LvHjWEREJS/28e1jCvz/FowJpDLHnB/2Zvx3L
RYSzyi261R7lyeCrZAjfArYMxrkGyiHTtzW8LBUy9KOo69jRFWqZGpwOFJE/MgeX
jEjcK1eAGWqMLDfeVK0g4vb2+CGsa6UJpcQktoS4B1pJaob5q1z6YqxIrrVElLPe
S8t1M701sLf3p2k6QGXtnmD9cLx4xeejnrUqvsaID9p3sN5tdDsgUGs3z2GYQKJ5
2L3+ubUycs9H+PyuzE1pp+pqDi0lfBNi7HhJSgjgzOTYaRLZPVC+RX9y+ekp2JHS
d1K/hOBn+hoNr2xEFhta2c+kzbbMxu/v7gmpbh+S2ArJ7/eu/w3jJ9shZlvr/gvC
wdadQfcmY/WQj0ZjtSFXgFOUEXOIMdodLwKFYuNLVcn2iTgZKOPG3DyQT2YFiAFB
zmPS0UjkulqSYK2Tx35eK27xd6DwHlMMF9IHfAIjdcj5cMPhcNejgHkEB5n4+aLm
nyLtooKJHDYc8CYdDy00lU1z05rgheQEsgKBmGx4IUDDirYum5POvnRA1nvnNuaw
2xvFNKFbtFiAjSFuUNc7iKVxjtHyF9WtWq5MF8zh2sRyudmMs156J3LP/VQP79OM
QKJ1BKBM82k2IkgeuyNijeMfQJm4ntRIwvwsViKeQgFr6LbvzaIVvOC3zBlidiTr
HWK0KWGAv0JlQHu0kbD3KxMu53kYqkiQKY7iGOVYcAnWtEw4YDRQD9kc21APWcZk
5LVt83Dg6eJyrBQDiWWcNj3xJ2N9g6HVKqGmR4CRjJiAc7dfGoW0Q0gTOkrOhW2T
s1yfzpmB6n3GwwRU3wxrCSsCq8+gOI3NcEMXg+5DFuERvTIj6KU1BSj+sd14yQMB
+SqRSPo58hkJN6OmU1jlrfMgXFTZKnmMOsPeiYv9DOIM3H10AEW/JY0ymLGga6En
ZFTzJgsEj1Vri+3Ob5Dbpf3oB9e8ZXzbIsEEiSI6JKPUhwn1oduo9IAC6G3n0qeO
4WBV2ooh8O/341+ibo/3mE0iyiGcozYDWpabGnjk/EbyxksexvBX7eAD6dA5CoSM
/DceCiPS1OeXGrVUnl55sG3ADDKamq/JvVZz9bZbXBfeXFV0F0GRtyNpmFP9V+TD
HWv/f5Q7lWOx0/nfbDIvCfz0IiJR7ndESdMm3U8Ui4uF5J5v8VEoTyAx4ZeLg3/j
/Mq0BkRkOrf+UozfluyR5g+i2riAt11X/WNyxasPgr8bsW/PmWnT9Mt+oIbLVm1l
9D0VeXYK3zlQYLg1FkxULXUW/zrgLz3wPhNpj1G9YCtBu0ioySqJhy+vYyT9nCgI
NtbPtMUHMAJWvR4KmHg9ze0sQk+cwi7oVMEAUcKDhnGoEr7hxD/X5zEk37gPK7KU
G2vr45fqz48Nmc8JEZ4UoaOnckewdanI4CNKqgDSyV+hlhwQ1zsGbVjzLxTH8Esd
ehgIZ1OZsl6tKuKi2HZgFUKIzPUGiHHzYCsGflo/Bhic996aYTb0sZdcTt1ixZmC
q018tTipRHNcaiw92vrCK5kiM+5S9K9bCIMd0Jk17I2EbgYVcbWxi7Frjly0JHdB
68AZGWHK5dvutzm3XztWOxKAoTx0Jm+VR4Ex7Cni2MsZoHynyVMYdfIOLmVySLU4
mm6qX330DRGnLtMrvmMdBRCOCO0g9gx6UoNI61JB3JquZ3oiwfXvQINU8cvbJ/xn
FpNTvq2E5eD0182HcmIXQ44Q7lX9ga8XZWmDuu4vF2IlPKf0nJCYXOAW+UrqSRBe
BANZVAMu0gcjCs2TAz1226URW+bLxZkFlZ6jCuMze61wE6UKbfSi08SM43VcpcSQ
WBjvYR+TeY6QMdagJbB3S3NnVE3dJyJ91DHirHva3s90VEaqnqkM9fE+CFYxSuIs
x6oL70LcZ7MHTLWFbmYqAeyA4C7YBmHAXnxjzQUGgfZk3pTSurlKKq+VOBMA/Pdz
K/yXv5tas8wbyF+UcnIDbYTJMN+gQyrrqroCDmeS/rG+jFvE6bt/B0/evdeOHTF3
rh1XTFKuQBc9e4L7SfkFjW6+SpjIKwG0KQUbx+7NwYLx5/wfajVFlpScDrrtiJoT
xaoPNHNW//Me2dxIa3ZrcaaI7vnSAzLfx7TLufDJAuYsipjz66161n7dNlyJYnti
pUnMddBSkz1xZ9V7ku2/7JLIII88KpkBVby/xfbgwx7bsIKUHSjNpy++RBxBgOHT
EPC7u4AcQkoZfTyRsHA0dO0eWoBa3uNYXdDZZrgnulbGFTOEGpxZy3VOVinUgldO
4En4WDhRdZfLx64msrrk8vbZVGs0Z4X/9E4620mCY5xOzJlMS4CBGD08mV+4TlOb
aLAItzWz+UxOQMzq8pBsUvuz1ETDdCv6ZG+ER5WTAVqsdKuX7RKZQzMHDWNHvn6y
SaM7OPicRhWWOhvNkkqnQDLXRUULoFvXYppmRiDQrqxxiOO+Bpb/uWGlybTyb42E
p7gLh2U63ciuztzUmmFky0VG/FDwAHUGYRvrK9Yb8y/Zl1MccVvvF2YezEggjRck
lUtvApaq4JB49iEx1z9UNjLPP2eL6shVI5wTVA0JT431yEkzAjroYtEEfG0ewDJO
DaewAYg5gndk+XDjRAjVMHyf7GraeSJDnzCmmVD2gu2ZPfPrOBuqfbsKHQjEA60A
ERCznKIa8DfgFknfP9c15Q3NMC7kad5Qk/h4YAjslkwbJkiFtum/okh3qZ0GyJPA
CPkCvqF5fbVUzO3PKfgOW4qJiMulJth2LI3RFwOIdFZ+3+ZxRNUc2KnuSNUQ+1Io
KPDDUlEp9pv9vZwHqkStUilBaULo8gfXBCB/1JpWEea7Sf7caeQ3Cx/RgsUkDVhF
SHxuN2tWsk/ePlQfnN/G7qeNglxP1M79S/9HIxlhiavJcfWPxqiaTQwjRcjMligj
GqE1Iu1jA+ZlnDFkehJ4ehKptqiwli5QQzOej0FppyVTO8pHFShSGCIi0FXZNhGd
L9Qbh2AXAo7b6uOM0AoB5jXyS3K5Sk2BdjXaGpEeOKp9aVRoKtFB/6OMNbUB9pwg
S0qg3iHZ60LLO0O1yQuqLeTKH50Y0ItpTZMxiDohkfUQyUXupgdetnXo2NJ2T3Om
idWw5pinSirFIHj5Mq1pxEgkkg90FGRNy8gXn6rHXlJ5iHysI20Tcckq+ONQQKzJ
uRXeENjaJCpJuAUqCgyALXdKg+pFLsTa6x+ZaiKAHp03GUcWXk3mXyzz6DUwCcny
syynjXjn/Yj4zf0PA/Ppg0hQzaMUHdhrhQ1klsFTqvMfth63KPvfRDLEPVqO9Qbf
MkeejRgrV0gyQa08mcw3eTVz+wafic9XOxvWehhOW0bvF8P9mQHduOxkRYCQd2zB
wZrVRwthmo8jihAaGeplzAk6KnA4i5s6KLaDznPVYcDaPQ+AjijL3fDxwoNQeFB0
5MZnw4/Wpi6HnwPK28flMqJ9KK/kclmdXevJ6GV7DdkFXlBzpSGUV/3c+PqdMNFF
H6SDrtbi47tGeMKFK0VYdOufbREwAxFFEvUXPg0vJlfq9HvzAPYslVhmRFbCd4HQ
qN6zdIRHz0EsjqdLvODUMrC8XlJQ4e7RyDW8XGGiVCIhxcBw0cRGB3cKFPKvQ5I/
yKVO+H2fWrSV/zzPa5z/37fEwt+yxOemV9RC1inIe6GI933dlRCJ5j3Je8xzuum/
qeiiNBr0D1v7C68L+cirJ7DFoG+FPFpLSBnQUjKsQTkXaKhYC01wL1FVNMBGYtze
NYqMTtu87Ot15Kz8CWqq+jVDRlrLt8F2IuiK67+mU2y4OfohlLp1HFchUj50f4VI
kppCoUV+BI/iF0BwTpr76SIj6iWcD3GcSUMtFWlJC4npgcej0+pQ2GKktlOmaC9S
YFMgWSu1N6nqPxJk79fWCM1Vyi1QJg9G12oeGTTFJnsDDIf7wyyJKhBWnHHnyqhF
k3U2gXjJd3fyu20DKVqEjVmRaYTqMm+87pf1AJ5FSzaKe3rhNzeBK6hsHq/nCyP1
z46RE+yHOJSjnxVmItkjBafQQVtvCX7HJi2WesOSTiVL4WAvh5s8Mx4qii5vHWAE
9lHFQw2Nvhnq8TxuN8Mow6+BnTyfZTw/Y01zl/kEs/kxrBEa9dleXeVKHRQ4Lf5e
HLlZGT6rbpTrOpZ0fSxgNQ0jNS26kQY6QMdLe0Dkt0MCgbYF7oBByWUUL3nmUQnN
lIA0y6jiQeToHgHdyVHnQplJVD4Ho57rmRsgT0Vjk2+q4AVGOsBI7Q9HtFrZ0gqI
fhG/ODceO9thu31T5jAmYRLiYl0iDrtN8EizCw27jN9MlDYY03eurklGu9kealLc
0nwoCpVOdOqG1iGqyMOoET3Ot4Et6sakY1NLb1RCKfkIPJ8rBYZULQJqPmPDROE7
3CZFleMtORsHCDbhIfe91oJEP9jvWryArFOqKn2cFYX+Kj0YWACGIAdnBADgG6Qo
RjuhcNV89MGjfMoLY3sizV2t/JNEd7AGi4W8fWQS12+k8PxTOlF9ixZn9bNOH61p
OivAkqihB+w+Cf/a7RvG0qej79fMx5JxrlaV/Gsn2VdF/GnhsYaKH6gQ5sRhrtQD
R8J8HmLJ+CYxlAnWhY2QVgn5sdLv6/qCz0uiecPOKDw2Lrmt3+4lifRHTDU9Tk5L
NRlJiZiCENz38I2+6o0MICx1lJsgxNU7YuY9k9GXu5oR0KC/Sw5K5swVXPSWDizP
De4D4d6xSOVCFtGmJMcxYKFyNFzxzQne4NUaDt3bIzdpJO/uxC68oJgjvN8cd4tX
oLfP9sVeEztXeHdyQeD1nSTsA9nlAiKrv1za0+5j9sFUnnAe2padf9hGUuaTQFL3
taRv8ylrSBQsNyQMZNu26XP2R2det7gc32uCnyUxNCT2jFaq/61LpliH00ef4oFB
Gb8BfE2LpLFAm+3Cq4vi9sJ5DiKMYr+wBWWlQ10cgSPs1CfIgczId6Ct36AY2oCp
AvSSciypAKGmIds2epdm4vf8Ww/GXIyPeebnpMpCU0pL1Y3xTGwW73YTrCDKBKJ2
ld7lbQ248nHaur30eOsh9hQGmBj+wH9RkT14Cerla6cwBfLgoQeqC/hoSGjJ+hG2
7CrmsACAzlJ9A+DE/PC9R++mk3961A2yYz7GInbTdlFFjCT/Lv9ozJ6eAbfM+Qrf
zjWaOTyVMxIW231OJiAiHczOBZpm23sm17j4Eb9vHVG+gWsRS9wrEkr2C++EvpPZ
hSXjGjj8Y7z5ZxiuNex6LAKStGpohiCNvSkXl7Rw33rsGh8fDNfvI1xTxkYWkp6u
+Yqz7RkxM0FRlillEQozv0FclSitHF1FYKulDM+mR58bwuhyGsMqDDt3kx+APj8m
Hee44GK4NP6+Rflq16GaXctyVsqYu0zuWriLdyL539C5yZpsSOp9go3CBlzU85cV
bhsTTUn776kCoJh6I3wyWGrjsRzvBiQEfbQJIXSgKbpuR13SIQHPsG7cTSeeWKv5
wq8V0TSIlKJtHzRVSAGarU9KU07T6lv+uXeyDS04cBI0vKibrCl8Jwr+LrW80f2f
s1liWhFSUG/41l+xkijfM3AdvoJyGBztwWQFdulN1gGqoIP/C+/vciZXN7ADZj3X
1XelVxTUlyz4v/tf4WwFpRqJwSj3i51ouYidLfiwtJmNSWZdCxOyl15cHuCTwyhL
1ZKyvd6V3m/i0dNxOoH9nFF0p5jVVATmweuIZB91ZZNsWgBn4pVyz6Ij3BniGZnd
rjvo9YSTbN8aFbEh8t0SULv/N0lBdR1vXMwvNpVw1yKk/77oIXRvZ9k6VirxSXUJ
13GAfHhle/fjWFP5NrJRJhO4tWd+BRO7n0RsA9b5d9DsYr4TRuPY7AOJG4y1Pp5a
fjTYKTZK2jv2CKnMbnywR1dN1DkOLDCG769yP/+5Tz1geMyvz4um7CFD6qC0hEMs
4qrVJpiVDaUQ342NF1Wl6gJvDCiabMPj7ZNUmPVBtC+pmHZc/Kb3UPWwP2G5EZWS
XNflx6Ijd5+XQZD1mKiH7YHJ3CRqnQjKKQjgT4aWz7KaZGqOXJPaadakH8UKhcgg
XpaX3jFgZQwm24eSpwlSfbVHUXZ7h2/OrX3bgjQ3riuKy+A3kWBHDNTgl0XUDvbL
45DPyrrupjhHdOepd+nmSLr87jhdUvXkg/8DEJCLikxab+4AqJBH7zlnGENtn7W+
KYShWNnGF2ksPd9nrC8zLYmuFr8BParxdHC59ZCojGUuXspAENqo47jUTJsnZqGN
jQcFBqWzEZE96a24zsH4aLnjYHJQqxx+c5yVcjJXb1Tp/VeCJ2sNL3FimJaCnGDH
KG12XBtgdW/r848TSfkbre7oQxBvevhebOv1rzz6tu9/+PeOIIfeqtIFTlmb+K9V
j/17klbIFs+/nD0cPyS3SnuX8a6V7zXYpNi8sFWcAiF88uDoF9D73jzgNSAvD2Ri
K/A2sZSutMEoUwF2Bqer3bfCJXCDbsyqH1LcqwIQbz9Aa51rvMC91L5YWjxe9/da
aCARatcGdyyP8JJKOLwZLj6RzO3ZeFMEDlbTcyNFc/4GPr8GHRleg4pSWtEsH4CS
7fkxr/RvNHyC73eZmPJ4armjM2S7ExM76Ltv0ENqelMFBTRvt3puF8QppjH6ohzm
IbKQEMn9s5P3YwYaDVLjmAGtae34z0vR8Sv06hobUmPVcGXNtPYZy4/NCLyvmRye
SHUfyN935pnIAVprqLenlI0hWeUCfVGeW0EXGrFCFMyrxAfnEjYc+SRHNDTXPyak
S0SP//t2NR8uZzn7gk4P9AeVOGLvV414ifPaPiwag3JkvsoCMJn/KbCjd5++fNEa
kxsTnyhMncxWtYq7LOr78tGiQ0ZMLM3AvA0HujrK97QyVg7u1utMKwKCp1IjbgiO
JhfIZ6u7X/kpAi03IMKDwGMyaFtzn21Z2tl6LaitaGKdK76oXfp5oOIfudi+6HZH
0lMmEArvLPDMf0wfNeh3+4G5+oBJHkhwlq73usW5UkvvM5WW+3PnBeXzaAewj619
Zpx/eDIb+TKj/p5HLsAEZiRYFgXYyYbJMxQZi4CXejVVBV8y3DpDg1iYBKTozqsw
e0QKvLJKoNaAEY5t285tlAhaFLYl8JKWCJPIAEjlSHQULjz3bQW2StTM8zLvEmSc
BhAzJhQhB250/a41cQqRMXaVUZPGDQPQ0VGOcuYYDUq92OSAnDa/qcwI519ANu54
G0N7EuAEMb60h5KdWh2efP3YJhKqLD2EkdU3LK7GbQSkfuclzut0n4I6L4jIMU67
JmmndJU2Nb0URXEatv4E+iwFeP1VAa8TmoWjGQ+nJKml1YHYFz21YA8eV7Coa6+w
UkyFA+f8P/UZq8giFayh9ZlrMBAcU41p9nKv5nbMcx+l4kJuZS5JolON5Xr8Bro5
VwKmJnkrI8uMDp70+Ysp/oxAQt2A4olSef5/x2wF9LawBTkXUWFBtHmGSlSKNAYS
KAnCDYDI6gJPU9ecAfp6tZrW7b6q71+0bvXdrw9aSscfDtjNdqNEI42gFuYkGd+P
Qcpw60BsETKU5darFVrDW8M2nZqgNMTET/hvPt5cSIVV3Ds0mnqoPHjWV+eQ92Os
pEYVBeHMVnb77h3gAo3L+YMO8iK1WaWluVFdwvG3wR9TCV1b0rYib9+bvqO/k6Gk
RQ2B5FOxau171+pQE1Fzorw9JIbPlaZvBV6BXvvoLjSv0lBjrR30PfNzc/IOiF+r
7/fVRWCmJXnp9pIqn4t1793+aRmGosu5/o+oaf9imJ4TakKlsgYUku2dwgCIUQHv
VRVD0zaIUomxmhXSMgr6XA==
`pragma protect end_protected
