// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 14:01:31 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
TgU1JdsjnPwWHlaZrzmL1w/fcfiELQuKiCePbn3e76fMPOsQO7z7kQC90VhjGyow
XXy4JrVTpMrxF3hotWEYFk2zNDTYe6UUmkmm9innxg+5OkdD9b1+B776SfAJ4t9L
C+xQrlymDFM+Hi9G23a/THBaSrCKShvjdIj/445ct40=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2224)
7GRW/qAMw/FgeiKUKYmrmteXvFhM41mwMvHMmxYfDp+mxzc1nwNZvn3rIg6oNQO2
8fAvB+JF9TCbvWdRG8fbZDcNhGocemNLlf0CI2l83xka/g2NExU1BCz53wzaXBnm
LKPwn+4j5+qLG/VYfbuIZ/j1PjNjxWZK+JaUtLvlazaDDbMPKfZhHmFk0cADx2Rs
jloV12aNpGZZFni3VD7aX8S+q7a1q50GUBo+r/MvULz32gHcaHU2RBS5PnP96rIN
NwA1ODKx70dtTTuBF/WGx6h/P1xlYWXHuRGntnB1spbccQB1OZXDFBWz8BEnY621
jRX6MmgyMgvkW2Y3uS9Czbi2bCuOepcG1/8vbQKsFTajJzowJXCxTU4J6KUluNJ9
roTQSnxEch0b4fviJ53Md7XaBxy6BDN8CWgIOcDVMHfrfPsvKJ7CVdfOvk8q68IR
xIwaJkAhuofs0LmomxAbfzS6uI3nGkOCLxs8pBZbzPDry5I6nWrtywRgLOLApdU9
A4FBK1hqlACP6IXS9KGGtU5Ij80So65YBeIaKpdOKq/uipaZpfPmMwnV4GivbDOS
gO/4HkVsddG/VbiwpFsrxPcFNiXQLrqKOsyy/G5IQRekiRyl6rBYr0a/d/u94H+W
bwVhyhMKMhTmFaqooLt4517A4avFYSpqLTUjcm6YXw6M+U3BOiVO8bFZkXN7fz8o
FXYWJQ7cmj4w7rZfwBHxgdfbY5q2HKt6gJo1mnD25ai9WuRxlZRn0MpL00oX5i48
r1xWsCRB4uVo1rSxHV6k+EcqqugdJboGm2KMk7BB278vqzg0C30ubVqBPp6lMxjW
DacEoSl/N3wfX+ZbtGw5fHRhEdHCYx9dj60xZuq2C62c5HfibqF7ARAFCfM8qQHw
STjR8/oFV56QS0b2XK2eyac7BdPaJU8JWF10LcGPR9WPYcHEJS7mCdln2NnYR7Ph
GI/blqY8xcjr0b8ksRvrDVls0zXYiHsi3nmennBiiNSKPjXEcbqzt1GUEqfHwWLi
MlpajMCya7Tl9tVddcnENwCOyHQGaKfAYOBneMn0h8haItdoa+6cdsW7ASmkmaCq
YZ/xpwwSXwK1GGR0xIVcFwUIFUTF/31E37Q7pMe+PrFxRfAI8ku1X5Vte99j+79r
qebIAt59pwzDAR2pC2ekHQaiIC3vCSzOW/Ut/TcnWfawz6yrABuBr0ESiI/dutpG
9m4q5I7M7h5BzoMgf/mZp06D2IWQH5c8QEAA0EZIZzeSOS6/55GcpSwKICk01i/w
ffJoBJ9/gGhhZN2ai1E6PtiYiXdqVGob8Yn82OuqnSamM2y1uqlr4BpFs45Ye4OQ
OB236TI6heGxO5BphJ7qERkzeUR1pAnI7NQQXbUBtT0ledordS0PbGB21eLhsHWd
aFc5P10xIF1fLUjvilipWgaXLxbh+6EY4lg1qLXgvH4K+wscEjXSEoIcXgIgXwrN
nQCF/zBee/YeI9RWM/33yIaQRpxFtDDoOXAP5lV0MioE/QrTyzf5BMpjTjGEPGdh
mZry5av39FcJ7AhS30N4sgs5JEZKK1O3CWN4yaP8llJJOw0Pe3fpSsLrgE5Mlzur
kREc3abjmIkeTP6Z7k4aS2GSUr+PVWX8KIp0R55kpVBUL1sn5QcEqwHXwebu4HXP
BvKLC4YnkTFtqBtWCIRIxuJc7BK88jkJXwCUlD3SQTbJYtdjJnVHn4e9+D0RCBbL
UpZdT2V4H23WX7I2f4FLqF9XgQtZjwQLxb12F9BGpMAjZ6IwWuT1XJrFDQ5Mqadj
P1ND/fFwK+Suds10+H6OcgOOwLUZ1TFgypv39NtLqKQsdaT8mNtdsHl/b7MWt1RD
cfz5qo16Ki2k9N/tZq4ihSBm/V15M0fdunojQW3PhVcPmKt5/6v32FkcDzI5//GC
xJt9XClj9/5OD+6GGGxAWUua+xqqHIhocHUKcsMLFThhaIZRb905/3M5PxhyqeNX
3dbqTx9fL3zxlDjcqWzwiD2FeajnkeeYhiqoSDERjPlxJ1zZ7ZRyg0ik/NU6uu4U
3ZuuuPMzt443mInHXHkqw5KRZKZf/r3HoO045zh3Px8CdIPnvoq8U9Q7l5dHJS/Y
AdoSKNp7oqgzt+0UQtmHmE7zNQK53+mjuFC7rT/VGladL+6MwjYXAdjvGozALVA+
L83R9pkraX2zz/35yXXlxp7d/cdcwGnTP2lR6h6Ss0JpM3lKUGBR6wWcuAP90lVj
v4E/Jnx+CWrKzb8144FPZHF4PwJIwz2zx2QE6jNou/55YxWqfl9fcyxiS2HGfbIR
Xfwc85Nhs07ivENRWunIy6d1souWrX8/a3XOlsMLVzi10rC6B6MySf4fhkOJtqXD
Sa6gRndbjfbRGK4X8261wY6d4+/5pcQjPTtgsqXlYqa5Wz3dVyxAsQTqum9ZL8FU
wZnnQUh5YP1Ho9DiJdXuucfBvJHARFgUdO0l6FtPgdMYXNloNo7ArwPupHL6ahtM
U0OnWyiIzxa7CRpjkuMRC77OIM3/U/Yfmt/2sge8Bg1QX5JzD6pU0sTJHXWRlLBE
s5lDKvdes9E2FhpLu7w9cRzEfrbUYf+mxgJD/PJCti2i32sSBt4nnmTSHfNls61g
2jOqGjLgneuzw9YIypM56oHzsJKf/ltzFjJZVj9PDcKhV+SE8qzPSC4m1tANXIt+
7jlQzGXaqBLAeatjGJ9ZR6mzEziH13xvvwsx2HjkuBHuUjb5RByJLCUbaaUIWfPL
J/tSGgjF9ZIzm17fwpWg+8dc7Nr5sCHmbuJqBEt8SvTuZOPc3ozrgIYS1XYWJM9T
RPThbdBgRr23gcY3SkT91vcwgKBSzM6Ko40qPPS9M/fiWq1L03abqu3Odo0Vf/th
J5n5pCa8VhnkY4UwX/QN5wNbZNlT+WZyrc1v0XFsFk6WXcavGbnKA1kzErdcObg9
6LpQL8MPYkWX0C9J5/XKwA==
`pragma protect end_protected
