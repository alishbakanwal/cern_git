// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:05:29 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
mwxgiSPM70KoRaDSPM4PjYOYuN+TYty+nfFXygWHm70km5+6hGlHBICqiLpamvDI
1XaL7EriQsB2lo7iCALz58v4IHc8km1uvviLE1izyHJNkgGEAMzKlRsQ9GvXkMWJ
F1wke90YtRlDdg5icKQnlrQcqOZFHD0uiveNuNpxVTE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 10784)
vkW1r0LsOmCJsOO6k8SldbPcrdyRlYzR8wrQGQZzSCtrH98NZv5Tv6yGiggAn7tD
KIDXbkB6ZwCgWaZcU4cW1OJ/amqR52XU2tQyyZsWjvxQpMri8tgkd1sSG+clxBOZ
2U6tPy3rekAx5f7SMAC6UBK97kOzWoTg8kHznsLrR9AJ25B8nEDCSFgvdMHWAq50
6ar6LWXgWe68Q2vS1qjiAEW4Qv3e54Q8sZOakU3Vxam+36Q/McjJ+/BVE7J+MGxU
LzWH2dhgFf1jHrUl6ncn4XbasRToVmFcmcg/2Ngd5iIz71JJIRKhrRHRzwbvU/uz
JV8AO0vbGuRkhxkAxwmO1Y/Zt/7vB/RBpIhlD4Ytq/6k18X5L2iFtcGVvN46iqDv
OLfWouNHmr/kjsMiKDBaHOf4a/PMwCaB4SwA/+vPR/iJNTxaNMG918EvYFfUJskm
ow8W8dQlmmbEDyVYjTxsfWoCOil4uAU+qQJBc7TEp4wJx8lt8n11zAHviFJbuxot
s14Bk7hLhyWbFZr9G7MthxZ4pw9+WNpJuPkrHnMv0njjpKW6p8REPRAYyjH9bSP3
Sb1JAETv3TOotjsddBorprAUdEJhKfuG8kwted3ideJpboIScEJ9MSNoiLwxQ4yg
kuMXds8rAwlDVBDuroKakmFR74nfIpRGawMA/X26jzamynNXI9kmYJ+z+TpAt1Wk
d2nZnhpssfJnUChPCMcifpS57tcvNMh+FceYIeV2F3Oz7Kw3VsHV4+QkWH/ob6Jf
RBQnU77FFuIle98a+Cd/PK/oFkLs9GY4cMOsTWggavvVdbjpvza7xcZUxCVf3K3O
hxYXeGVREItIRnjVCTgO+MCx6zzXhkxauQ1dri9gNPlVaRl8UBqu02eB8IHhJS2R
+rNKUSppi0QoCCgSkFQAKoJdXzwu5w0KCh0tdS4LddVD8MgCgdaGvOd98Ex/N9MR
+Cj6cUKlWxfdg8AD0v5QHT1jlSBqQKnF7zqjn+flNPFxfqNZwVjUXxtXGWW3vuSc
LcvfXjY8bTR9TMBEeoeD3JLzZ4mQiOZuej28PJHFuFAo26SVk6BrtP9IpKb7QZPU
AN1oscHTUnhWVvpN8EsrB7FMmN/WOhgYxB6jAjM5Jz1UCKsTQdwNrHV9AGnMzDfA
VhhhvV67KswUgCFutk5tqBd+Mijumg6mitxKe/IPd6rAnl6KM5/QWUn2FL4mj1d/
1tmQ+2GgCe9yYaKthGkx4igYx6TZLN/qZvJMcEFouRDO8lYZON2JpIFlGShNFy+u
lW0E8IP1yJylWeP4AfRWzuUU10HYr9bUIcoXR2vupZ+/krqoKILqhUk4sSlkK9PW
2Tc6pU6NejJtSCBcD7Fkr2aoIZUWKeF25Psh4/pqvcLE7D/ZnGaudZ/+UoHyk5Ve
tImqxHj2L7t+eqxpDitrofv5tNdgcINJMR2WaMgVoBQWZQSKbwdaPdz4EoQkrT9h
ua+pY5OY5vC3p2NB1aYybF3d5CxCKKvNBsKedNvSH6qTvZ9y37n9xVsQlVD6tkqC
m5tQ2AIwzxfCxMlm98vT9kSNyiiP3ILWAfsB1ktRcerdybsZGlTtwGH5Uukmd5Mu
gWfEYRl39Jipof7mGO68nq1hiN+0NK3gfkzFKQrLUJsvMP3oM0Co9xjImh4PkxL6
MinPTTpUKhuDONCb/mNYXUC3KplyKETw7ud8O8PwSOg7elYSSszw5TTVeY3j1g5R
ofXGCgXf2X75ARaNxp0wn2bfRUe9z6odmr5kiAOAqferrVsAKBauXoJpaNwST6UM
Ijqjj1k3vn63L1ASNr48hjUEWFdEo6RMnJaU6BobHEzvZFkkj2MhyA2D4bLqTGYM
8hqSQAkgcnryubMN9QVrqcGF0iq6DV47MkrEcaDIWmCub8sRAsQixUe3Y+tzcudU
hHt1Mpkdk57I/jlWmw6+zb75QCke2wfOARmdkv0iZIpsEufr5ay5CYqtLsdOip+9
C7NGUmOcKTRtmnmein3GSgaFGSx9L7P3lojYpKEJad81UjU9Q4PeK2KxoL1piTo2
2PoNGQMHDDJXEaOv6ekAVfkYz3PMdsf0kQ/2PAinXpXF3s0EIoYR+Tgky1NeyEnU
T6EAeyHpmwj+bftR9O+yqvMA2zncuYp34D++iBIvYVbCG7s82ayuSFHn3rWUNn1p
5XdzW8UI3Br8JDaxYjsbIh2fUeDLMqzqZnekApr6EG+aVe14FUGLZ+ZVZWMzZamO
KmU0hdCofzQjlpJBderjO/IAXWKP5QdWQOaTp5Gj5u3MXqbZ+6jtB7yBTiIOGHaF
uEG31DbFMVF2gLQbW7Qp2/3/mUci5FO4iu+vDieoCbuNspq8xztTyCu6r2KnUOls
WN6O507iFQwWYVdWjX4qq20wqBSxsrr74J3oAsYQ/o5UULxMc49LajAmE5wgVG8+
CSBnwbJF8/q4jyi2LuVN5p1Ov9fARL0k6sRXuE/vFIO6A/i40ZVK8eUunvzO3p8S
sJgdSLERq/lvp+9NtGDC4T5YU+H3b3yr9zYYt2brz2QrZU41taEOQAUL71+4kjTs
J5VOUhy5CO93f3XQnZgG1s5gWHjOBONvtLDHFaxUd7YTjMBNYQhnodV6IAf4UAem
eQz3CE1jgmFEVP4ZP0yyXbWgVdl8DQXBWTY9ctsIQx/BDXnUEVWfvCfkg5bT2WkK
m5L0/f3Ddi5dJlnFwiqC6KGEFoOAjbK23KrWbD7H0PWfUbfdtoakRDLslrsLt2/D
D1SCpdZq/zlU9g2p2nL57QQuk2s8LG3Ab4IyYwyksst4iaGy0vcNrmRmw6z9tP3n
0mg4+xxo4M6PR2rBe8p1jEGT6k2LuinYwZK+bCl8WMG5b0ZXXUD1j+pKJ3EAEGI6
8pAjCqysGlxosKJn/RR54dz9nwzlDRkdgOdIHX6MUbUg9GcW4mxdV/nWufWbWpV7
PcoAXaRwr7MvEbzTT6dp8zsyjW/xlh8F36RXAoY3mRJ51Dk6F/n5CBavgbUNOmkT
vCrLI/Y8mAgKTwMk87Uws1KEtOWglF1eRMw9vmBMSYUStnDSq8+3n3KWL/6klcc1
XUSJWnTLEmhsGxxamE2tO8URtZjYoIFCAx8vm3H3nUPM2pnrxuUvRJId38FRVApH
e+ySpDo7SbMISOYhbHEMz7J6Beu86XndUXrI0H4wDsqCBsb5ggScUPcNhRnNs/OH
G8a32H9N2JuACB+h56nEiJ628Np1VeJx75Mkwp3EGPkRvUMsL7KPwn09Gp2csJKD
ZJPkjtVt6X5GsS19wwrMYA/KZLMudHXT7OL+H/BnsVQH/oGb4z9lPoeCSYQBSPXU
TIiOddx5z7HfIgM3ugNBvYRGSN7INEgKFMDuJgw55yqDfl9EGxHiL0znIkJe5Oom
uTCCix8l3tHCO0bCy5WFaafohafP8DKAZ3hBI2IfTtDdEEXBmbKBSvbivxDjTQyp
Fe2jA9nf5Irg1be3SsGNtcis9AJDso6MfSqaDHUIKhoNLWVBQ13hIkLjok2/EG/Q
ANCLeeGReySkkoVLu2iVMkMWFO8ms95drYQ7nqM+oFJLffTEhRBhGgANuMK9QEaO
wRGnUsclHutTW7i2Fw+Z126zJ48tv8mfxB2AWzGGc1EO7a5WPf9i33PSHR0wHumI
1Ifo6RQRA/7A+VN+Mj0z/0bnX04XIP4bt3Hvwk7/iQe0dZz47mmXwK5Nj0weKU/b
xbXHz4ZBwtSmY+o7FsxkyqTPamDnfoMRnOkdoxisMoVNmmoASK5x+TXbQ5sIuoC+
eVV7kppt5ytkVhqgw1TD9lU/H7j87XBT8YG73OTtlYU1EgGwCYPgeb3+1OeO/rin
flUW/XRUexjxCtrmO6AFyCXQYVDKNFZvbkEWYeD5iMwHM6lxcQWVqoCnSL9+NHcl
TS0MtCFHHchqsGnap+mrGxQhZuIUARh8vx4YIG+5iV/aT2tbS8xVhSYFdLTFQ0Iy
JLyMSuJOJ9q9NtzJ27I7R2qaHulAUMu81JGykrOekx4AC3r53yFpJdh3HhE9sMDW
eZbjJC1tFkMGWuMMeIMkpWVOfhp6uwx6tucz5g2qvA+uZ9ET5Wh0COvc40KI08PX
dh2pcUrEzYCo6zNPamGIm/7dnbFQKc4WWRJGFZJEx5Xq8mYRNiuvaBCmvgAJb+aH
YzxOTJs7vKv6Wp1+U3mWO/cLTGfd2XH1g7OAym8G9KCJHwB3sJ/7i5yOnD+axiUh
qxnRxvMKe3xwfazhktfE4ZwdoYcnE2ojSvVVT8+ksGeZmSR+DPeEAPISd35qs3gE
EqxCXvLUQy6eaem2l54r2a9yBgaotsM4uLU5tJSHQxN2UvyMxQBi6JhpOty1jCqB
pfoK4RnxsXXZ5U2OsumyfAVLc7BsAWajkdqaKk5IZ0t8iyKNvoSvan8N+OtbbEPH
40F3khwE9uqsBNCIMf4gyojzt/8Wj/owb0YnShpd9zi3s82nM7Bb++xUTRq2ymhs
zKrEOcwmqyUzt8kFyWkKnAHDvL4V8B0R00YQnzlrIfWJBDsSRqygxk0+R4OTmy/p
q4k3vcgCgNqMZOAcTdhOV+ogfvJ9FEnjfS0zT2+8t+m4P7zyf+3nN7cY9aJy5BT+
8GwtuVEBPMI8lJE0sVxgpHdfA3ZboawOqSIMN5j1KYzZiBa4S7So9M3RwXMwgE5K
OqToDHnn0UZhrrP3UjTbkIoFxNKsvcyo/o/E8xxguXmacHt4BBY6VGiN1FzyiN8k
zgWq+rreAfvNqer9Ym2YkuyxH4hO81wK5RaepzuIYrdELcx8phhtJ0W987pn15hs
lt+9mDzk7dzZyZZ0fkgUBACxvAQfXQlEF9quaif9D7cF+DLb0Y9Z/6jzAXhQY5j+
0VQ8shXN6GzB7XQZDcAQswkNpelds5/LCb1jSxv1TlFXtwNroZr4+omRyrOAm3bs
jiQbvby/HKzqz4a+2Hr1brWs6qzPiKjoXnzwMCdnkzV1AwmOzoQu7KmJpPSWdE/t
LQXQJgOXlcwrVBjSATH5oZAqh34rNdF1m7xf6jTYU6WKwu8oaXdJlzqX5MgG64yR
4LlZS8ZZU7PkOuEZ2XNHZDdR9hJY9VcWTQUpu7exLMrhqCE7YFkzn31R1XCShS6k
+J9t6weFn0Zg0u8RPhGEsY4Tpu8txOjahUOav+hRaEd1bWVQHHLXCwvaJH1sgrLJ
YnLSORI+bUx2dJZILUzRzVZO1+DzpbDjoYWz9H0Im8KVNCzx0D7ULivEaWwGAOQm
waD5lQuV1Lr2R+BsPVQRwRAXmY+/pK0rgrnBdh/bXZOn/4ugWBRgxc7shwS3sdAL
ok8ZVBwtDr/nZchZ0jx54wlZmSAWyXYOXIIlfRlTemckEtHfu8KQn1ALo4QO9ktL
93kJ4zkLw4edoBW9DIEZVwKBUMG1ykc4Ua9WNIH1oOMeW3EvOxtx/PZf1jesp4Ys
VCd/L2lnszJdsuLbDGgPSunM/5TAg6utdliI+efMxS8W+LimGohVCGKIncxxKV4A
ayOh7Rsl37Ob1MM4KTZMPNXslzgRr7H9RBTAo5ZfRNLjOXDOtLPt/Sva4uoRBmuy
DVwAqBMlW5h15D5FftU/0UikHME6PQiA1HvVW2PGxhzaYCPBCf+s8oQbj+xjMvZc
517YHNjvOqk0ZmSlu9rY1dqhEmO7ktm99/aC+hYfvXGnt12C3V/5lsWmy3WyoA5F
5TvH4soCQmkknwku6zrXlQaOiXzsiceBYhNxRerCIJVY9XrSJSnCV7O6bT3yOxNG
UY8r7/FfDiI6gbsvsMBmp8hRDI0OlsYFui6o3AWh+33w6TGDznT3xebVcSf9yhHQ
Frkr2ryq6FT7KtZQKGdMVni/X7wqtGu9cKLllmqAlZf5+aLkf02VM3sFClVQgjmo
AFsW6NMhDYie/WH8YmDutbZZAvMPKcc7ZLVOdEHYuyP46LQa5y6DvncTNKbwOYFf
kK5X+lrwX8J8Sbl3bGHIQpCXUpkY5vjyKzjuoBATty1Zvi7BYYPcZt3OxbWXaV0K
nqbzdA+t0P732k2HEraEkjB47s4f04ayKUEAgGg+8RncTIkUl4+vO0DpzOu62YCa
VwI/bK06OFrlZwHQ+DxvoBAJjbYq2q76/cUkqwvYPra8OJ6X1NSwv6Cc/1cBFH55
kOv1NLIY88RYY/qt+y0YbaSI9QvPn9svkLcO+QC1e/61CV6T30fZgPgMzcjbZ0ew
QkoIKSO7NDYlrL3Csh1aQwwN7FUmWThLE09K5YeX/WLUbwVEYrpPeZbmh47eWKSW
ickVaTp58Lx3JAsF1rp3ucC1ITbamUXcCOwQudQF+knrO7Vxz51SHwYlwJAm/ccE
nW4D5oul6GGASC+6ez2zmXf+cYO4i40QM6fLPGejAc2Xvug76uKmmlj3RN2NPGc0
/BSlREStk3tGoxriCxeP8J2t5TO8rPs3ePZLi5Xc8sEtZLKBjoaxilSZZ2dS8fcl
ijkMUAcUANxArm+fpx6j9sVZapPfC7l1GdyqPS8X18YpcbyvHaxG4uo6Nu4G97C2
I2RBzBNSyEqHDj8xa2r/6KKWxbt5IBKnRV82wyM/3X2cMGClTeEqBBrcmAQpfE0s
a78xGc+wscziaNvVJBhlSA3DgyuS+DkuBAFSZs8CRyHBezoujBMmNIA5RFJC/XDJ
FBWZ2lwD60ZIyUTnIwA4LaK5nvqcXUdLdpLeu92uDJ8k9tGTcPZY0ZDFB0Ls9Lqr
YB+29pT00USyJ6H4snBNMvECGnvGfH0dVoax1G6tte+NDnZqHQKk+Or4AXmzqwxG
5i6fA7+sxIg0/vl6EkK/PcpMPTGqVokmS2o9PxH6l4VwCENKr2dolslTszjH/Vaq
+qAoyoonc3tfDhEDq4sVNhUfKHZQ3PycDpmBghKBFcAQ1MV3K6i4TP71SbI9Jfhj
gevfPHUB2pADXqiiHrxlwSCQ6a3daAQ1vKA6/KWRtgXaxNeZ152zZJ7e/CUHa4xP
YybzhyZ2CrJWwlvkV0SjoEG0sZGYjE5TEId77VnSjt4xu8gA73A6cVz01hZvGlIv
TIiqLlXEo3QYMezo1/1mWpBCAtJtCWVM1jznxZwdSfKUKc3pSIu2CyI79rwYaWj3
YxNVY940RY/SJGrRfXoazcfDIYCyBYhcYW2ifsuV+MTypbDj4yl4Bi8TFlfAvUnJ
2G2A8ylka63YJq0eCsY3rp23fPIDP/TYtkXstHDYxkGe3nqIjscQMmLhA8xLbq3k
wcvHGXFfXrR1Pln6QlxYk2jlszJBU8szL4/L0EpXypwt9zZCexpEkz9naYET+SMS
zGohTFjp/8ts4NRKalExFYBdzwtDRDqqU9l5zAvF1XJvn/lDCm8eHUG+3MFjCdKo
AJmv4LyjpUoF584JsROIyPIQQYchggNQGMn4cLlH9+7JrOss7hAPnCEgVDXt99jE
GKA6gRdKEDju1mSWmorK+u5voOluLLqJ2CCgMPbMK/ZLPXPMWiVb8N/wUoivMu7z
XWr7BtqB/fvZ9eq9PRnGgFDO+/CTmnEEGmozfUKAXqpc+fdKy06S3xEDFR0e0L9Y
Htyyh5B8dTat1MwxKRnFKeCasRns9ypOt5wuLvPfLXl7r4DqJlo2ejfg7/hs5uu4
6Wo24MdqDrZhl2/UBpACZcI2RBVQWHJX76XBxAyNCTbYzW0IxNmJhmu0q9ZDuAZ5
QmqiwuFJ7o8LTm1FNJskrZWDN+/neZeCyOSBADqymekixcLl3YlS21TUJyRuuaaZ
S7jHImiA3lkrX0D4EAiOBtoOqX0tHyDiPR0VsYi7NXsnnCLApxt4HXLN6Fr3dfkj
By0IsHVTwsQ2fTdA4dPWBEawSNvzHEnsqyHYAq/xmPyArmrdCwJTRLxEDRP2rU7r
BLhXgK9dpDCFpKzwoxBw/8QZE4F0t74xh+VZxqhmCMqBKS94YZNQvvrO5PCHLLYZ
RYlBrsa9SfxJkEKT3MqY3JNhYHSUeJ6KNdp+yV2oc0Vct5gcejZk6E+YywNe32Fj
3GCt4TOFd7WI9avX+r+MJrxpf5oA7GLa1U73Io/O59iWJicgGLu3ADf5r1Pv3bya
kI6eb1NY63BbXO+pAShknZSkH3z91vNbrsJdr+CY8uJ9QMRdn8jY8423aCzoKdcg
Iag2ayWVjSxfxhsr/5EcrJPypalxGleF7TJIg2RGpRAo4CHVFSU2F9N4fy2gG1yf
HxxKCa1C5hmnyQ7Wj6CPw3BhRaOF25IQh/p1bXtApfWp3brMn60fgfWQYGMv3f4o
TzCTsVmWKrROKVZFAXjmulcNUbdIxIowrSQDTxNzjk5MsdsPdZvBVO1BNSPxDGgV
UNPcpIBJylGB++P9PLiF/7tEnSC1J9Z+FL0o4UyTWuyo4RlJen5dOVWB1bxV+Elu
OgS7QJWUH8WbVMvlTix5EcFsQctt0OZxKM29wMyITCDSSgLlYuh4F0BdzIz+1MtP
KQ7AYe4sqHWAW8/ekHuoX39Rc5hTWgXK/hf7NMmehSv/bpe1SqXLWSV5QC3NqeLH
nHWM1rDEayuEmvt5EDNoholIKdPhapelm1uJAaycNPFEJ7+GGJbujWiwVnQ7H8jB
hG3JXOpJrZryHbi3WB/wHkm8sB+B7Wt0NNloJNXvGlwdZ33YdxPtO6Cps5ImcVUN
oEfUs/D5xP03ibZfdkZWgWcnGW/FjXDtpKec9GUGfXw3Y9jO36uVm4HH/gFKAby7
5VDKkq18PW7TolJ/jF5e3NfvEgFpgX1KhO1PKj/xlwFcIc9UFVCzLh50I2v+8Wed
nmkRrvh9+3oLIHmvnTp38LWUmXn01blPcUwbFhwz2SYEuOJEW1vU8PsNzBw0SIZ7
MiYhGfNqeqKgu9mGnrip5JGsLWMM/pke8PAJL5N5twfMgd64q9mH0vQlYqLBwrV3
VU6bcwwENTf8GbvFR1zS1uOxhDIlP33sSWpgZ6xF161Ill6/fekEQfV+KqkDapjX
ihLlkYTiMTl9Vpr7/iDcaoLbtTG30o8+aRibyYZhFsLnvP42WvvzU6vR+VpKUU+A
ELibkDwAAThEWIaRqmMvproDFYAzBjrzY0euVbP8hWtpZ0Y0xztlMlvUjfiY1cn3
8+gTeB1AqYu67xf7tuiBILnQH/nplMCfOwqA6gStU+noZYMJ9IyW+u8m5m790M17
IKGXrTS1nIkIsEX0aBNaU08AHXcQgGp+h3yTf94HK6ELdzFilSScxRXk9Fc0EyL4
S3+3Wpv3ufHeAa7KrBdecdjuwyo+lnEXHqwxVGusXb9g53ETs2yDztPeZxvJYJHk
mLnc/J+9jNghjsFUooO2CzDVdEe4QZXbmA4LUd751vzew3NWva3aqMGE2GgCjwd+
O14XwHQPDojaZj7YkY+O9jVlwo/hjnIxH1m2w3o+gzv9pF/q0yurSNOBq67+qH7h
GdgW7bQSdxLaYmZ1WHC6koT8rE2I77ocCEFcT7b/BpXp2gLjd8iGjS//2zGtGZfm
14fsz/cgGpZxlndeeigOh3RWf1rzSDNKuQEqXbwUo0ahu0bKxCqftucSHEr4Xzje
s9mV3Ha5C0qXG01G69EpjS1+kCNP8PKa3eOrCLGiFT27UJUofun1afXiY7xVkvfZ
W3zu0ZJg8G3JaBkzH9WnqjbuyLVarlcLOyLIL1TkK0lwTJndpf6rD0fgdB0kK47y
hR6l3JzB9p2Xm0UnNYqa4etEAjf9E7xCVsJys+ftgMXCZMiAgc/3fcOHqhNqHVCf
n6XNGtDHzs68ctYsIjf3ykh8cJTk6fO//2ICprTKToOzhKu0zd8Eel3JqwhnnCsw
Zfm9GzdwTARO6C8uUnFAbg/m/CbTZyVK2El2X1xTU+L3mHf7szCwQh0B2tqSSLmc
Jf/wzWmDYhXqT4PmwbudxtfS8+qgQ+i83I/ZmUvYzmWhRBDJYqvL2X/Tjr6m7G8H
F2D5+jKJH/VBDsuhjxHJgYh7n22GmyFDrkGaOIulegxCi2X5lbmoJbhb1cvoXnc/
rCvvX0Y1puqOYH04sJGsHy47DepNcuhXsS5Y2yEZcIFhuZ5iq6PcJeMAv8RE7DAc
fNkYtumyMjYR1NwdKjr/7DAYdhpWdTcG8HxrMsnNkEz5KAFRCh+O2u0js0heCg+Y
ZJMv1H6KMqgRoxrdyDxwdifxdAlKSzOPYA/r3LcU4wPsiFThLaene6upuoRvp3O6
3yHwRzQ3dtinPc0E40adAOMiDdfuGy85NMyBfEZO4NyqW/Y4mL1CUjPx4d2oPwAy
i3/0a3roNT2fk9bY9YeqAW6p+3fsO40JO2CntCvgiG3zz7cKWw3keqFI81Oof9U3
xqLWH6ueFM91kY3lCpAGz83pP2w3X+m46PXY+wRCeZxhthnnEODKCLbrYVelbsPb
JM6jYsBBL/xPRR8XwIm9AFnhZ2qcoFY4GE7KfFWwIXhRV74oTT9sRWIzxEF1mCyB
E/GGodxMCSDIp00AniXwLdYK6vFCbHm8C1XpABsZ15QXAbGl1uY5rHB70+waVmeZ
3a9QHtEpqZsVhqKvaP0UjqWYJmSQ01iWSErcYIe3FsEfzCBQFDLGPIgjvUeMS+K5
c4PWjEyDUiysu4nBX6E39brbjmDMg9j4TNmJCZnt9F52113YtlSIgriC6QZC5HNL
GG50+McYxKUHhZUmvHt3SEWQHan/85svXBb6j0KvVjeZ+05p/7DD9ZF5R1wKT9WS
tj4wJI6BTQMkH6N4ifqocic8OwUkKjjvY7W01j2kEAvn2cbNzyOU+urPT1Puj+TZ
rYUxUNlfaJpNkIkdiScqZnXMe4MibOqvuItLmTahZ7/pkZkqAy2TCx7Mx4H0GjHr
FTLBnh6qAz5/eQ+ACadfNXP4hGSUPpXERZuiCEteNYCXcAhhx4ukYmnSV9T/0aJ6
pcVuUOkYULphWUPdpwsvTMK80dk+Vaitxf2t12059wz2yn/8/HHpymE9xHpFOa0E
WcwSXAq7P9HmG8PApBNsJoXXOTrCn7bhZxf1AKhdA4r5SgGeVU7yV74pTEzAIKGN
2nvV8/wwGf7DyErJzXSXuuBxOoiAQtNqWr+aW6JB8MiiwEIEPJUDx/B+Lad6dgK/
sqOQTpmD8v4flsrXx8FGHUQhtbcyL75idRCuG0v9ScHWXEneeuzJp7dZrcWO5NsU
iegvuy8+P+zihoQBT2Mpi4i3+vDIb/lX1h51boKPu9EH5h/m+9Q+3Bh2cfvYeDy/
W5koGYVlnCr3VbCrm3WXOOAli1xJLjmvHaw+S3tTgH6gYR69SqQyYe+JKLi1F3++
ECR73B1n1yZQkOLRyTfWs+pmB1hgL87l9cykez5dMEWoPtm4ofJPq0U+SSVEDN7b
qK0ZltHTE2qGAc8QzqMgWflU+qzr5RjNzmmlysQokJp8MPy/AcOsmRP9kHolyubR
cvuy4fdSpZFN0vkLBXKoZqopJGJxmWIWnw9kzUjzKyEJXugs5SuV1ceuoKh4m1Ln
k7sMhyruoYZgn4fDSoyd7os1xkS3K1Wvs4vhblBPzxJ/kqBz1UDIJZ5LWORpsSyb
96HjfMaU97jpJ2Aan6LQRBEQ1BV6ctJgXXzztB1nunDeKDVBCJsXFFDFIaPu7kMo
r8ltDhD3dFraI8627wria+EQ18Oe+ZGaLEckiDo7v0sCfWsEFPyhJiOztigy8IRm
cLuYvcpMc+pyKyTrus74LPY9xnQPQ6pfPgwkBBGWH4yB1UJsBIBVS3grZCOcAAac
cMNsbCWADtFTe5ROlu/ioFuio0DHzczXi96RbqMBokJ94E8VmlhWUdYDj9nhcMAE
tkqMTDrkCgiipM588BO7B6pV7QNF+cep3Md/FZhbFfO7W17o2HjGNVnkp0M7U82u
wzhdgHF5U7p/HZwc6AmakTbFLX5rfgo+3RDspLp0Cwesab8OKetoxBXp4WxjzROz
NqWvhxOAMJ7rWrBLobxQO0qHcSlvtBvnGEIkB6w3kQvV9EkByW1PW+ml/2kWRer4
/bVo4C9PhET8v05Ed2QdGjMNvDtXuUM2fcHRKsEWXST0KNYVmG854rBH6Q6ji2fI
IY+KKerlUXPLYmYNSDKhEI4nndJpG6R5gy+jP0krDkuRwieyEB49gpS3JOAUAXKs
T6j0WUKVicJP08UQI7wQaQXHAEsyt/V5oXFmNWFUbxxDvrZmYj9cLFc6wsCSPNra
qDHG9qFjQ8IMaWwwe8+EtJeb6Cy4KISkNEwA4htBH0jdPVsHo4bueAFvyUX2OaB4
RUlcpkSqI4c1H0IFxmZ26NT1X/23hNgp64x5XwjZmVJmo+5SGCLY4mYVEqUnN4Jy
0KYjAiR7LkCt/aW4Ox+iJdAEU6M2T5xIJmFWD/Wy0YA4BuwfaPRXXpl46igEP3ou
q5azErdjAMPjLe7VkaBuEkUD1SPIDI1CPMGZ2LTxwvwAjKbP/EsCdTCn6jZ953cL
tru16Izz8xQfJwsbJ0aIs+BZZfq8ioF2EqO2aGEDV0Ad5k669jFib1lV6ie+Bbu9
UaDk/HGXSw+h9DVT5QL5VnZGkiqlqH63g2LD7ZpaYxb1szXkoccSrGuIb9SU2EH7
0RYWQYvtfnc4khqKxX7fbG2NFftAW56ZcA5WjB4ruPcq+eEcG5GKchrHwtRvZWFM
1JM69i2UuJTyLeyIiYMweZrQgBFWSln70IXSeqiXTZYx/ScY9IQptMHxEFHoG7rI
1WZ1SpqU86cnt/NIxXDwJu+WBXrS0sMlqaKweLbPjCNlXHg2ZwKkTfFJoUZ+7HXp
0delo1pd/p1B0evi74L7wIfmQnspoVUT9Z72eU3Ev3uALZ8PhhzjzcX/vgLaY5zr
xKF5eeLP6GeWGnXpiSvBFP47cZnfWk/1c25d0fJtrZvyIJY1cMg96vZEK4Cu/9Im
3318B9w9+BQtGaHAAcvbxAiZT7b9VHSoQeJ51oLb/zEsVwi1A/0zpH4UUEKaKhch
aKTZQ3RLoXuHxYp0vF0u0o3AvNVha4CtP7iXjz8ehMy9DAT5YvhViZsnu5HCPU1C
LpW1RKW/5AwH3z0QL76iCoQuE/MRpMcp4UPG7DHWNrWih4J13DIbduauUgqcdCqE
GThsrnu88bo/VzccIdO4Wu+4ASJ1lM+bStOwYBs+pmJZtjjduNcDbnlew2O7eFFU
2QKlyMbOZtdNs9aKxVl7RP01dG/G0aKz1DfxvyLtDyN7tfZnXTCmcFd/Jaar4n/r
PA9cLJOHJrUVKYSOGZ/Qfgtv8a9ObMfGk6RLxvAZds9bz4HXZxjbiIRjaPTHWLRk
mW4Dgy5eTGRcR9fIwfe4ETvGmsUYDoEZvfql0KGW7JsnKnI+IHJaLcdUv92djI3g
9EPgX+gMpJW1NnVoJkgMo7NFfqdzty40PH3cue43NaazmigsFocixSPlB9XBaqXa
Jj2vLKifbK4lPTzFvMYuuj7lGypk1bKUQjMUuCwn7/GusoRPwNDDaSg/Lz9JOiIg
Pttg2EwX7Go0kWNOZcO7kBg2UV2W42c5hO6Wva5ptAOxDK7UapGqOawxfQhoDsTY
jiBQ/5wB88eiZT2VzWEnbcxja0CvUWqaqCVjC9sMTsETzKTLcdINAP32O9Le/liq
tI8ZT6Zn0pppTE+m6RrZGzWd/79PYUMVEppj+DJXr/10NJ8Dyr12/cZwc7jxKMVp
1jvKdKgVTsaw2OsX8n/J0n/q3RZjThWE/PwpdmXHUbUz19poiURKkLUj1jvtWQZu
z15o0gzFxtEJiH5us/st4OdPSDTEu5w382e5Ra2KppbHDYdjS4TIBlR74NpCwmNq
OEcHb8I0LA7Q5Ya2VdIoylZmbJoXDHoqnZoUKk3PrA2xdOesB5YBJotTcLXUMQMI
PnqgFzxzFcWOkSWRivb3zu4zUEBJMFpJvKwZkBSLkc60XZr+xoFz4aUaCNcvjqyC
yMCoz3Sxy314ly/FW2wQsOiOaS4ZiQebMg08PUs8BZHeDHVtkm70FxUeY1jN1Bcp
3gv5xQT5VpjVmvZibA1rANCPoCiE3b11fkDDxiBX3xAPYlWxlkvodgEW9GL5Yl4q
GvXwiVON2xvfksrYayd8g3hyp48eSvACbO0bbNzh1IVewkbdpLgaZJEi9lyrYkw/
avrMJnWXrMQrHl41e2ripyQvgBz9DtnNrTz13uoQrjO7c4+2dNuMOKAPNR98LcL1
paT0mZs6GVy286uR1HYj67nrsrLz0uVCqJkMaGhq5QmGUww2z0mCTnqB6kmpPS/7
furYZs2msD0vLJnefnuI8a0+ZqDjI+ekooInyvfra0OuzQX6XScPYnsCOvefWCAu
cwP+FT7jRlA/v/yUXT9LUiihDYjojR9t0SFIUGXY1YuedAV1+nDNlMfZkY7S6uTZ
d2izaOR+ucRInPcmNXyXLSSulM+nbe6G9+awS1OHBjc=
`pragma protect end_protected
