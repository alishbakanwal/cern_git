// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:05:39 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
AqG4CiRd5a74F7G15CXt3KboVhiFYb5sKajTmPwfvJBSc5T4QTOJNaqLy4Mq47Gp
4XUT1mmSoD7FSZtQ2yTKzt9O4z0kje2PugR1Cmeo1EBDw9PD4nMEolQtvmBhchwC
EDqJ45I9Aov24ak5iq0uGAcflITR7S6hlTUACeTbXt4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5216)
NwhDGRO34ffvHBiEdg577/q+6/tO5LCFXJ6NDBP2gzxG2lCdvaqgHPtHkCUQV39x
noWtpJMCz92Etn68Zo/YJFyVFI4+D8O7szIQorkkWKQTX10ccxz1Zqidy8u4oIg8
jc5JhEaGe7EQsIUv2g8fc+udXU78JsvSL5X+2ZLYOs0DY2RMmieeRphi0GhU9ZS2
jqgyNOPyRb//ZeZ9HL0oEVaiNXzQZHbvp3Eg9yJmafoo7oxwcVCAwRxhDeLVpZbA
ZwghWCG8QsaWgcCtF9V9wtG/FDGkVMBqLN3fMFKw0u0yMinnEXLuhKo1lVtUUR2n
rEqhzouWBgi/oLgiHH5nudPUKT/X1hs1d3h5agLSjf5sLqrtpyA/PmtOWI7Z1TnR
jVX/HQLXjY6LCMknMZuuVAj2Kr1oQdk07ez4uC9UCPUofJ3dxJzVyGzflMSPjZMJ
b6/5cxgonQjOwM8UJaWNVHkfiZJBXKxTKeKLMSDVAQXjHB1aE/rCsj+JSG4aU1wP
qA2BTcBaTrJAnNcJncClWn15X9P/sklcG/5hIL7dGREY6Edo4uAevMb32L0VqDye
OHboy8/LGnh5JsH43dWICQ8GaSG7cPCl3PlZjqo9Pwrvv9TVTZrMlTwEyr78r82O
yp5ohUgb3wnT5dUS90XTXtBiJBLDLRzjLAcM0bnYKnDbobJ/220V5lImzpmLGWNj
oV23yXY7kUxFbImIIBjqj4pyZ+Xtk1G5PDzy3KQwsd1HGs21hr5liK1lwv4CbddS
7LshLGb3NNS/VAqGBn0+FwutfLFX1GGGK0pODk1FlnJFWGw09542vlJKBCi31NRK
eeW8TndONHTag4PKBA4JOIRx29ZPx32sMR2sEQzdsZZ3Fd5DhmZqHKrCLCHqClpc
lJpvE+tvHzxcC1NH4V60XV86s0shfTcWW/r9n7o98XxYxhDa4hLXlospCWS/vapO
Er9eyH0IxWhNrFO0THvAHwPfkmpEexRzepFiIHbi9nx72R7NwOwUHkGa+jRd9ydQ
SGasDhSo3BXd9nIvK4c0iEGOKohEZWO+we9jx4fylcGTP4z/pYDi9yLBQIg7KSP1
JEHfxMgPQkmmfm6qpYZMVJdH7N934kKlpgDNUghpaWueP+eDTh8gQFuCUqVDc24M
vFD0PrHPVLEva3mke6obE4WWMXy1sHiTgvZe10h+Pn7diutcSYlJBcVk9tvSQVjC
liCvuPYuzM/xObRGRv0Gdtjm6hOPDdIhm89wxGQEatlcn96xIyApNfECXEyvrDAC
CfK6bdMiE/Y0HJjAk2SA3lud0WBNMKyoOaoUtVWLP/an7m4zJE2mvgDRjAg93TXr
+IP4GNDZtkiaDxSKVAM6zGajgLBaMnbjJpYIEGZgNH2ahFp2VMytM2zjhMnvCUnp
yzTkEg6r8oikKnduD2dN49/suOnq9osgqPLdAXaK3HOqoQpKYZAsBmOnBtVsJveq
iXoVlbZ70d0fUrPXrkcM3yFIPARomCGlh1OPxl0F0t4r2CD972Oro2tcBgE0Rt81
u8yPssd8funKtoZL2x78Nq6zoj2rykwKzc9OffzbPJ8DfhTZiHWiKzeWtDJ0I09J
LWVIYa14GrYASwXaF02fsQVqVBYj0XA0RAvVa4PxHzeXYq16Cnoopx+bl9qLUMxR
/PSrlrme9YY8zzi98/bgnAOrwGVJxKpHIxQtRliAUlkRDO81yXmZAY949DcXpJoG
WP4RoE2lwCWMp+ANHQH9sjiRKOPu399DEx0e2kXItj4wUHKjmGCFXbEterxZq+rN
CS6ONzb5wLTAH8fkvw2IpNaDemGtVFwOfvHWfaY+uelkNrtvzCGligu9g5eSeERm
AzUOVo0UYLxXmrU7DX6INjD0ROHKqly0gbP2ddD8Tgkq/ljtNap+Mk1w7SSfZ3JM
89NEwxv7SQiYKu8aO18YF9fVHyqeOUYT9w4lyDy8FPWRy7t4X5AS/pEvnc5WJ7l5
8I5+DlSGUWeHCf3+WD91R0eS34SL/eQedmNkKqpsaaz+IBqEOdhTu0DP1jBzqWVR
KpSkGLcum/kLTK50WruMJ6M2SUG+uzG1fdK5ckkpKC6YDtaSu46eqJtWTa3M5FaU
voXQCGh1CarWFL63TNt4OKyQ3Pn3R5Rgi8C4sFOyJ/XdT/+4OKStf7O3xs3XQ35M
9PyUjS/bb/MTw7h9EiJxsRPnNkajnJiBguyLOfv95knTsdU2YnN1B6MIQ7drMOSV
FKeuXAg+5aLnQTvPSqmNLQGU7s/mdI2wdOrkd5F+1wQTWXxqU5kutUOM/N/iQAL1
mM0lVhXAUQr66cQsa/iwVLHe9BwBjfz+pH3DI+8mIRbpZiysbInhHam/BvrOL/wZ
+AsEBXotL1m1V+ejPrt+gtgbbAUPCQNwC/pkXh15GK6A4UUwibDAGlXkN6221ECF
3xFpn8qzqyxURUhp/ArRRRP+AS8gNCK7Jdf2R1vABz3w4VggIyunRJsABKsQFTUZ
4lK1yNv6rxYWar1xC4BTqB+GumGdT3TNvxyJE9xUj16luQH/mtU8LcqAKZoN21Ww
HD9I+PyyOjAwccyuROJlnbywIj+LEw8O69480NOsgx7PVYyX+fw6DmQvMNCvqyum
GjfXj9mu2fYF+h0+4tT2bVfjMhkYqJt47Brvw7y1ymFwWJiS04nEUT2XfrlCZUZd
z8CW+Q31U0m5Y6uLrboQUJcmNJ5ymJBybZoYUvVYB84ZXOl04Xc3gLLDhOiMRiSm
fdxIbEoF6zMowqcKCyZ05xkMr1QsrkIfijm/SBvn0LG5KzweBnGhst0HGfk/kzOJ
pcBolZAz1iEbyX9uZSSRntO5vkB9t8TzEchaJMSwaDPJkY3vmB4WAHcQS6iWsI3X
Ag8dqlxVAvqWfyJU/UeZYowx0PrpuMNoPom5bkFQVUYO6/QY0LL6okGxmIu16GXc
ug4isuy/IjFar3NG5wxnCq+538YHhlH0iw2APOhvPCjI8Zj+cwcf4uojztSwBVUA
a0XzAiJAE/PnrdT48KF5YStvatwxWMcUj9YbMPU/M6IwMqasSl0HgkrSOCio4uB4
tGIRqTaOl5axRt8tdL1ZsLCqFUG0Muy0J3q8HfVozM1qxRnLkA31Rz6h5dv8P3uJ
+2ZCrlwUQ0o1AJLSnFzpYgyyz9MftnCqs8yt/Zcfy9DUFP1lfbkrLp0p7Ouh9aCl
hqbVmu780rYDxYM1LL8iSo2EjSy+yq6AZUq8M+OU2PLcesQgStvFl+7yK1J+88dM
+BAmYSEferMfruh46v8xBI1ANYsJbCn6R1JFAvvoVL08pYocY/ixcsQp/QF1UrpR
bCyEuOb7sCrak70ktMhI1TR9RM77UpbEVpaXC8vlirfD9p1d4f6K4Ol7Gw5rFHOk
uz/K3TI/X5CBbNy712aWKJwvoKdxwk+egsVeicJ8u7+JF82E38358N+dpNTslRCi
u/D+s38KvM87Slj5FZ9+5sD/PI2q4oRqikdsHhh4GEA+X2s20tMVy4Ji+qvIK9bP
poRPNwmWQH1lQYaH+O3iigMwC8JX4BA2ZjYr9ha2Fm6u5y9wS3P0/GiH6015ujHM
bcDroilYmBvz1IiKtwIni16Pb6LF3XigQi8+pTOZ3tD5ecvIGzBgxrr05jS2szRQ
fESe+ApQVIs4u47QRdsNAfZLWG0zePMFH4+sU/U7hEV41RNnTtlHikOUygtnj2A7
o6c1sNMEOQFqlaZnpSdqM9RS9oO4GVkNGZgzrlDSHpoPMBZRcBHvRE2NxBfpCMgF
gZr+HJx6182iifxUcLrtDWz33nQjtGbBTB/7P0X6WPCEL6cO5LzWTHQv9zqJQ/cl
3eo8EAzRCKuTRyanoBAmq+5nwetEjdS1O1t35pc5hg92QtBDhN42dYBxSLh4VHlk
lOwn6NiNKDm4evHNxrakxF2pcpg98haUDaIFKoN1MrEvgFjVlWvizhF1T5ZVLfyj
Q2D1m8foWWRI3kKuqyLB/q7YxFhAAx3TOXEpgKr/VZOjimFCn+5/1kMbNiOrgWym
T8SHtAa9x2TeutJpf/BhLe7iWB5rdEfeOz2hAdSFbL82aKYMmfJz9p83Ro129tQg
0LeVMNfNopKgs9Bn1BntUx7hoCBAl/NUxVvlY+qBWYEwdSlqCl0kN3lhWFYsYYt7
DbspfoVi8S5HmaLaRGzGkxf0FmokO0gAqlYjUVnRSUBtNdW2x/l9OLR0yY61sPio
ZvVPQrt3FqRfQTKFfApe52Y6TeE3HZnCZ91rEvsR3DP/w3DKKgnSkW2PIB8uoqWX
ZZN+D4zkFUAu01cUYgfPDd9dQxKxOEpHMt1yxOxxXprnCt1ay6VMyxNQ+nbMJ4rR
jX6F3h/Xvjm4tHQ9wOca0uFM4Htrwo09+iKpEHKsACSMjdiEHIEICclag9wIHx/S
RxVNCvp5Lu373tQmaruft0w/jL+KGgA4QE7qIIws5mDvcaoB84ggDxisLKleMq/6
1p0m1boIKmRri4DzOd7aGGn8oXrt8XuT8W1/qfnbELXJL9+8EkF28J33xaIzDAHS
x4KNfwFx56xaX1BCUvg+3DhojJ7zKABKU8wN2sg/jeKY43rHIkIn1lzLSfoiV2rH
6WrfxzVVRlQVL1j4xgoo+CP/GQ+x6oFb7XvBYvsZkmBaqXZPucCzIz2wNA4BgPuY
YmynmbsVDLd6HuJV8vlUfI0+zd++xovRExwFnJlHbeni5Hzd2LEfnMToACcM1lja
0vNeoEXq0inY1DAi0qVMj6OU4r5v+ggoJljQskdyq7kbsirlrX8EMGDUk6GjEQea
7XyGWF/gLx0h3u7sHqYEkFhDryhkvw9H4P5LOAQidBIBc5qmP9sdCI8B4Cmwnh4W
Zw7HOMsU52o76NZbrYV/uqfxDxPIw14K/zqT3SGXGLWGUL6/0255uReeoKkkkraF
rV/L3u/aqk0FsIHQnIViHyAF3eYMF4iS137FMcRpVre9glMVKhmpfrFlrCHxyKeP
a+O5+4CHi6VWEHjUSuhH+Tl4+pP4UbSeOnalOGVYiGbE5B/hd1q/U6ct2hFJ4YqL
GT62r1hyxUe/zm1aeelr6c6cqoWgIZCQUwBtnEMzmeCaHjaXMf0IO8YLRILUT3ji
XXkOQ7OI8CeD6FvtFNGA4SNNuEQeyRh26RcNQPKCGONi9/PrC8p7w59dJubbyfO2
BQHzyzePZEFrCdOyR79+K0d1HQmPvUTnQKVaiUm6UFb1pZ0fqf7cmpHPZB2UyaKg
rYJno5Hy24GKv28j7jmMqLk90ba1MICsA59NQoDBxsZSID3l1+uCr54zF8t89tBK
QrANmo16vYIfyojT1yPVeHISolO6CmxS3zp7kKEOAxL8NSy6WFCfqgGUYSnWNj0b
ZQSgOBBWI+RDLfCbcJPb4A8Knn9Fvf3nmIHw7p1twpXLLDR7ZKpChxysrqan/6rs
ik23tJal3IR48JnrvH6lku8PkHT6GTJFDlcfi9/qkNERHrYuJ3cTOlnGUvEWg5bl
Xuz+0V9GzJW65UQd4P/v+/1dQJcP5eEEBLfQEYt8ibTdMFkTr6uuSz+zT3I9ePOU
5B7pV0E6xkdWwNxOI8pv8Vm8Xd3n0luLApDDPSvUvta/wXMlWR48h402x+yhxMTe
yMgblZBm0NsZ9++PBSbHzfsKeG8127uUuL2sipTa/ECusnShYMxtJde25I6SFSvi
CM4HrreOBDv15l1K7ZFqsW3urvfovuyx1y9vBRV0paZi9FNwTd5cAN4Yhh/zfZ6Y
CYUpQkXPSbrz6i7TXD9p1o1+r2jX7BXdGxtKaElNPtCobP/KgxB6PVn4+u8IcAZ9
/F+Fm03lpsL3VEnJSHZsZVeMOlG1JSl/HiNLkHiPtFt4v0W01i16obK5wWR5kolz
JAlrH69zhy5h7Jrt2m8R/Ad8islGiyFzufOvNJz2yiYAje9Gsk157wDzpmIBefus
UbgP4SU5UtqK6+wlOcwYVoDmZBaKYEUKDWYQX3sy+qxdjbgxVCSJ36pltOGBq3qt
/Zpd6m6OK4ROz+t0kPFxmOq6CPa2XPq4JWz8ypvkqVaWZsk9kXeMqX310Ovs8lad
AjiRFPFiFoIE6fSlAu72eRcSUSLRMC0QjTvZvO8ntrGnMcsmVKmoGI8MzkpfeyQf
81Pids1by2o2TK7aoyTopOCsUMNQ/f665+ndT1YRKqPb7QLVdc5FNtHX/YClHf+3
5YMovrcNTU15dm1vf5Fhb6npe0AVfHQwLXcz/Wy8CFxmQ65+ZeR5qywt9V6h6yVy
QPwuQL7TMcQ3F+vyzGjWdbkYjZfu09q73DQM2NIrRYeHX2t+0gdH+clLQsWTaV+j
IPFroCzuqBWEH2tS/mT9iFPSjj6cTwuGeEdwaNOhwUHMfhWw6VJgqg3fqj5wF9ex
d34AxhD1KhzxbiQUZfwGOF0f6v7+BJKL+tmPik2ZxpATTBY+6Iu4B1eaRF1OWUYH
qglc54tpmEOcg8V2rsJ38SUA6pJdvJruZQhc63ax4KNiU2qBuOSjkKvKQaEaTMls
F2GELwDQEkW4CY4zcoEXdv26TLAaukQNbpd34Ovc3u+XM896lMLr9GTdcdM7lB1G
IR0iZ/5zDYDVUaxRdmzwmnPrxlDSeMRw+pb435dBSj8JYA9mLQBZbOhfHG3Qy29j
x2fa3wifvzYWEI5q6IZ/v4dMiwYuviM/w1p1AauHWTW1b8PX5z0a5TPMXh2NvCSk
Sg9zptR3iZhfLvEaXlK+5HVrLfVAByKYWnFGdxjQ46Qu/wDjILYM1X5tIcRSzkD7
cH952qVCG7h+X2OeLsfOvkEPMgu0va5Wp/cdhWry86s1upLsAZqHyS47mk5XnXRf
+MOEhteT2rl0m5STvyt8w28G9DYjnzv+roH6znoN6UGj1P9Iijib3QPRa5zp0yc/
XLw67O6amnNuEQoG71gjs9cy23raik6fb/YFEdEuHfY=
`pragma protect end_protected
