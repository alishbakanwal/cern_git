// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:05:36 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
fFuhgF1cqOOp9j4C8IRm+FesBYwb9pEu3g5OKJsvfKZ15hegTGYR9VuBmktH8PN1
bDg1S9H/6611y62BmDQlVjn5YEpfOnJcKalA14wjQagXPsWh5U5ynpethgMGstJX
W1eE7KLiIKO1VxvRnqjJsh6pCC0Vkc72dK39XYcSpGk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 13184)
ICkvcHiJvN6m87D8xdb6IU29Pm7Z41jZhkTaDBhIlI1dMTEgzBIs5dMRvXxNrIbW
YZ4a1yfz50WY0amDjMF0AMdt6fBG6DHu5+RY4QTRWO9R3Ez4Aqf4j0lXmNhdMzC2
dHtYIwFQwNg9xCI6jIpVyQu6JGQNaRA9ZsPjVcYiBYS5Ud7dt0Y1kxk5P7zF8O1c
DABixPvU0Rr3AiAnyaQ8yCmt36evi1bYxPtQLdj3jTo4eoScDY02s3GszVavXxF8
6jA/qgtyrCWyAAmBVPxtaX0rL6RTSYAlf18BIMi6q7vSBsRKBpRqzea9HCb+2F7C
SjEaAoxKAQJWNGYw49ByktHO9eb5Vp3iTBhLL+xgYF668uzx6e1tBohasRTsvWzg
N6GsOQWthnz6qnY08Bf+8at23xlLCPLRfn15ZFNIrCM8OkeTyhgIFoPA7F6po1nz
obrrcdsRUqN8OWXt/cCblvAbcbXNeTc04hk2exR6STxw3QDKdWHL8nYqiiKFCAtw
T5IRXuLs3bFLgvvoZVJS7e2JL+orua8YSqgf0RPBpoW9Rf+gva9McV63fE9kFfN2
640+hSdBw+GiYpI8+a7r5lJ+srBvXrFKzDzbyImBJIvW8FnxNg3Ely0NUlWKhxs+
KvD6ow+xW1fYvkp09WLxGJvzeTV6+kV8IxRMBNxckwwKTjXE5/j4GaxS4kSA/7Yz
IzcrU+IoJ8thgqiVCDjbNvSW6QcpMYC5fxg577hrXv9izV4W+V00uQ+kB/EELkR2
OOzL6QEwO6t0ZJE6njTor5gGA7e4+DX22p2Do2yDlVdaXiE+mCcEfRbucGWFWcq9
ngkQh8HUYSCKUITB7myMjzO2UlTHrtB+KgD3ZSaYQ+hKiw/uZqAyZrcF3ukohmXe
ORilfoYELJSeRoRs55U6Zl9q8V5xfcESM6VNz7PqGTsdnDw/fyKRL+Mkhpk5QuUm
1N8V5VLxXs7gLXgyNm45DZkgoKrYD4ejb9+UJVf7d/Otx6MYER4mq4veCtpss8FP
Q8b8DgH3fG0PJ5ClEDeEMj/QxqoFy5wZs7Rxt9Pdh8fAy/fvB+VqBRHKbimwTntO
PUE1kds+rAoL57GyZIpcZqeXyx0O8lQteMLgl9uT2pNkBloPYQy/WwPo8ThUYfD1
mkHx8oKDbEXHbRB2PYHM3S6dGLns49DR2f07ACVo+JgAw6aWHw9R1d4ZboN2T2NJ
KjvvNRr4cFfCrKxbBma2gXe3Nbkv14jtQbx2L0IAWdHZCXJ9dQOtOvC1fTNLW9dL
VwSMfeUtYnPEAVtXNWzYOCgbFoG1pJBJ0eaDXr4w3FlwzRoL6xVn4vrc9td2kckX
yCJA1mduZ1QI+sGLhzxDKBMwMJSMR9VbFEWYWZprc+o92WYNEoucstH/lOVgkmzZ
hpLNqWlPFECdPFk4s39PIh5h3JToS0TE/Ms3mww2LTBavcYxp9xmfo1SZGqYTr6n
wa2oEFD3Un2goe4+S/lX5g8TInUPXLh+AF97HsDYU907ojFGUoMW/ckv+QTDl2sK
PIPUo4aIQP/+eGSwdhP2vsvgVLs9FLU20T78Lxb+QYGztyQVBffN/Q8pQvBT7WQS
Snnx0hqLGebV/BNsFNu+PzauhME5DwXpqdE674Mjzhq5ntHwfyqbpuMMQh3Kn5/0
SuucG/3rKFJnVM/0Vh5uKXFwKcGd0e9aN8v53JvWhf1OdTv1Iq0aM5b1L3kZih2j
emGalTwl5BtGPA0UOk7GWsC20vAJAfgxMxS18lK8miWpqzYCK2WRIdyZOVn5kmdm
Qa8arXjOMWVVzj6ZGopT7eVAjtg4fpUf5q756pL3gRg7IoyWUKx5sO0B4Q84roYJ
qRvasLMD2tZ7x4VXfjhHTyP8BhR0gKNEX2lgtlqeohZ+855qDmjX5L8O7xA2b744
PIIeTD8Yc+s5ZSChfjBIF96rZ7wCGHm4dKZ0GLwFHzOZ/FSz7pZ+C1fDNxrT3O90
twTLjvJ+zsqqCyLujx2QNa2T0/ToWnHoTPNqizko0jsJPSVntCalEM7FWfbuWokA
yvO0oL1BmduKyVsZQDPeiYerU8MZ2dX75J9BMP6ucjGlTUFyq8xZ1hasbpnrqrAE
2oAUsGRhXQZMUmN/IPNLo4zjLNSaCRwLCgGJnxw0j1xTt9es1kSLgJ7DinyGrUvz
l+89lA91vPUKyjUro5dLKdOQCrYjiRUYSAabi8l7y2sPGzB4KlUoGgscMhgvOArY
Rb/n3isHfsfUIen78heLtvnW5FapDm2hDyT9s8Sngy1mL4VEjCuWMSuIMQG1Lt+L
QQuc4lZmJrgTc8ah7J8w+sUhcdxpNp9ZdCdZCmndz2smg7U+fgVXqSmPca9L8wyt
zPs6ax1KkBQBJOo+JhnmpWtcZrOHU7m0I/JLmNw4FZWkBYHMB5wkXTRK2rnl+UgD
1w+4NHbNymjhlvSL0mHzLQ37JV76Sv7n1M2e70oe1aTMb+3g/AdvXvy1KKZYCMXI
icnY/8xvsjYLA0yHLznzIosUIEzyGmhBHEt8FwhU3o75Vkbg1lS/Aq1+Al/GaofA
tbfD71xtpmVSg0bO4f00YNp8v3q/rf0s31Re/ztz0slJHzVodGyGsFSoQ/ukWJXD
48xItNfOwmRXDzUdPzV4gTzKna0lOMLdnti5sg+Zj3TDTK4Ut3rQyu4RnbBq8FSl
bL8EAPoFfDoqF+LyVLDvxl5kVV5C+L8vvmyb9frUp4/LsQ5fRl0mTYQ4Sb5x5U+C
AI63DmBNOfiEkjF7N6W/zLcLd9qM95Y/w13kM8ChV0j5gYjiP9Y3ll1AEdtnV3dd
ThJhW3K3hTuG3NL71v437koAFuV7JGrV1GW2JKMVR48niJ3wAPiy0MFr6CPfY42I
TQMMpm3atbQHkbrlo+j+O6/V3FDkcvF91LaI3OkHfvIdIHHthN4IQwJIRNSI0Az2
BFBfdMOHK+xe8w84IcH/bF4iFlu7AExgxh8TEFstpakU61RYdy9XfDNYYqHMdP7G
3d3+33V28ApZbRXIW4tUdunXvca3Rh/cB0ORkl0u6SPgUfwm2qKz+gm8IBwdjBPI
YikWu/HZ3ObZ/yIP7eIcgbFpP8tiQBadDf7kuLA75dk/2YxYqMz2Guwl3ZO1ZcT6
1vShgAa35t7Gd4eNOVqdvSEvVWSnOh9NfG1KxxSuQmDWO/wGjBHrDM9fYaTHhi5k
ztfcWVM5EQyANZ3TpOgE0j/w7pQLFATBwhL4EHayF9VsFVMUj/ZhbjYKILQCoY3e
rgyCX4sYx8pKUnA9ZNkaxz9JlrAVP9M86w6g8xGkMWnRt7TNsoiIt7XUMxKMBTMI
0Jw9U5mIsngeCd8NP33aTTpltxPBSYAK5K81iVKhO1OmUhGjxG/ZwClplsHmGX04
nnCmbn1bdOpMLVm3b788IFm3qDxeON9nr4RmVO7PWgbJXNljlaiURc4moOknscQJ
0p/eJYJsyff/x3m1c8XZl9voOS+1eXmQB3zLfuaTeEByWX7VUnTtNNV7Sp9C4W6M
LalFqUds5fturyXbbT8yZ7aYsvAMPHp1Ow/koqxVC8BlertDOoNYL4GJLdgIOwC4
iQYfGKBET8f8uwjJkO9cFavakIyGHxNdJA4r/AY2ZffMuSHeJxHBpHMgFPMT2m7M
B7fFXql9po3287jN0C7Oko1FddthI+Hx3PpwJVJuBUWCG1Gi+hGozXaFww54Cukb
0EE/WOczgIV2VqoXGaClatwFsJvXBEkywfZUWkkYoZxI5U5eQfHwUkeNUdmSiIMH
24nhOXtTvBzW9EUZWIpKuuQ7fahuEFiaX0w4mT9KTbPbbRVbtM3/NwzFV+xF6xLy
JN9S9Mot/eEz4n876bmaXPhQ6fBk+Qv2IOl6iWFRRrzAsGV8HEpgnfr+JiCarSia
WYMGUfDfNeHMdNkcyJbL5hZPAtxFhew4LSazljr9dwQvAc56rSSvVVImnPov8rmz
rgrPnZwwdYz30DUurC9SZlmaHGKL52bwItCRgb1L4rzlzuTfO2nwRVTZVHXjANP+
G98pSXpeRNEfyi+6DsVbS1JucIwUMZT06GQwAyXO6tUutBdLQ1lzn5Td9BBaXokO
8yYiWV2qGnjWYgmc94zaRB9X3WL8Uh60gRqGtnThq3g99HV5A7ZAm7ChCNc1oojV
qwflAmwZcNWXrrsXQL6VVIWMVscYLfdVQy888NJMHP0txXjM7JMZeHzSRuSqGlgh
EzC/tt4Kd+dXjSYDMwIcf8aMljcz66BBTu/OjjqiVePUoEbD4wbinY33XWAJCWyV
OIPmveTPReaVAn910TrtG07O5uiIR1DlDCKkF/FkGWVcIz47i6FySZ8Xq8F6r2Gs
Rs+dCI6CCGxR00kmjYJdgch4wLXbn4GDcjgIfTHeJdi6YhvnwpOWIrgDdyre8FC0
nJ1ELDSF4qdn7yAcdw+DrlITg6O5Xr6xbAkkV4FSH91bHs8XJn0NqhnLRpjZNEcU
rRvK1Mvxn4om6DfQID/4Wfn5oDWLezfTed+9l0GH/wDTJVvoqtLb9HOF+I2dmgYX
5x/ztnKsBHlgDorE9oURh2rvgsFwTqOQVO/2qqckbVYZLEQIyCkvEjdtPXl02jio
SH5LvBr/W2osFZmZIk6E6nR3kKD9qH08B4/I6QFoo4KF7lU/DxP2nSC8MwczSqb8
smc9A20b54kXrDOUg4fjhxQX2naArsrMvhw7mXHmZP2DgW+xYswxSjn0HJvJl/jA
hMGPGJy68M2f5jI/5lN5VqEl/V5K8cPvFm9I+UjrHqgG5pcolNVx117GF2+vdsbk
TMLIAOwgW/1W+c+JAcy8H8IrNMfI3v5eOTyjwWeOAVtk00tRTuizj6BENWp2mzZt
Pdo3BnwKpTAPk6sbQoL75ZsNtlyjJ+4T8mWIHpkK42jP2NjmCZTEDfyjBBEOcPKE
1uAaLiwrbgO0ABcTzJeml6jVdyPtQncN5O1blnbsah7kAng312OoWW5FDEZ8uAzp
A9JdpvT5a5TGl+pyt4pQw8WCUtJeU6OsqtWYIOkVXF0IVXH/X0SCEzS0729s0E8G
t/qn0wWOSSTUHR9BP2jFiwhPqci9/VdsWZzlVf96RiV956l1S6w4ZfA70sI7TIoc
Oso6aF4Iby0AO39yIKjC24qRRUePFPEI09B2VNK5G4et3/Czt41F2LlsvWUYDPaI
fdhdW+zBD82mnF5bi82HbFT7KqJSOlznL4lUWGoikYWfU1cudMm1TGBYG6kjUm7W
BLRhbd/KdXEqr3/8hcOl6UQ+UeMJ0LZqlEoDAifEnJ73iJNagqMtHZA6ZzEEUdj1
Xor9HU3jP0dhz/aLWUeP/vEvjGBIj2G12QnhR8IRI/fI+hHdEDijCRegit07xDAC
UmJZnK+JWiTCyqUKFmcWIRjg0XMGdStDpjUuo0Co0GFDAqGJq+iEDKCUmy+a7BS8
BbmTYsxo1y/OLgV5+vy7p/8QnDab3fbOH3/wnNiI9mV+ZULEIDNMg4yOBv7ma9yG
4CY9qdJJzXuyaxhh3EHBpltD0KFZiGAa6AooH6WxFL1pmyiBeU1ou4GLweS7UAi2
cRsAuRbU+NAZ7AieNKRVX9YTkNZYN5BQjO+Niqwn3GJP/NVDo2VyshT+1ChBmffm
0Pw6wLUzGx+X+vdfEVEKRVy8obwIShIEChvUwxaC1IbVyZBic9nx7M8arlugzSio
aB9CReXfbK4uf259lsF2afCFT2dtqAHQKqdsP5cZwB1ArViy27vq/+hYDTJ81oaM
Hd2HphcnuRUNxhRgZDxBfGgdpsOu8sYTvs4c07u1n+n0m/TdC5FSmqjwoVMBeOmT
PKruiHiLk96tRSMMNQnGxZSTClkg7n/dd96YbjZtCta50o3Nr0ZcQI2ownZ2KIKz
+o9yXAXkWd9BNPUUJnl54avfIhybVug3KtZNjTJ1XfyV3f1fQfQFypLmsiDKWDqm
0ar7X/aaI2Jyw3vro9g4+cqFRwwV0Litv7SKbLIT95aggMIgTgYNRn+44FSYd0P7
vgEhRqfBVCQ49NzrvknNTiFUK6WJBZV8v2dY8tHSTrqt1O3dWA0K4ENh/JY/YE9V
1hC6PWKiqdpytnZ0jOrW+/Eb3G/GhDnqJ/CngRhrLagvKjAhsSNdcNoNqub4FsK/
o2aWANkNpXuWnWzwRkGQ5J2TR458Mpgzl2LEvlxY3bGogW9NfynTJqz14Roy1ewe
LpBglwE8Z1o/onNdY2yAOKU2YVuf1cIKZrd3Anzy0luS32WO8LSq6OjrmNYQBgi8
+lvvxD2/i0aKUmmg+kQfvVZMfDrVSstITGxfZzK4loXFMmnhqeZUIOiAMb1HUMCn
tLTDtcx8rbtXMPN83cE841Zxndnu+DKSQ3eMWVzE5h1lW6i6LTFreMq+tV65ZmYD
dwPS+jtMtgRtjZegqVwaVpmP01S6LNvvWtD7XQbByVKHTWH9zXsOUtxushyNtSJ2
qsB+KAx3NDqt8mL2QjbXkD+A8LcFitpV838+yAhZf0uhg3uc9Q2ZDUhc8oiSnQnG
+G9t9SRCwHzc26CBz8NMOth1GiSWdnNP9117ACj/FX7s+EVSr/YSyvs1bIzeCKa/
Gm4WtktQiaKBiUW9sYc9a2KMK2anmyPm118pNaPzIKAsLqGHaHq5iJJqxdAWOCa8
f8WcdOXa1FTYginRx2Y/MvHTZv6tzw8FF+IM+uvs0rV2+ID1PLjuHG+aIz2qXmaG
JJvv0Iyaut1+N/AZkrvbGrMOocB9PQZxba0KIkhbWU8QkJHZbTcZalNikkNFkXVh
85EYHoOYwgZep/nmZmsEb/IspZeSd5qEOHn9x2MRMaOhc+47i0Kd7V112NznO19W
P3P2vqUgUgfZ//AFq8kwH/LYypTjqDqx53y0r7q1q+n+BtkIUtjp21VoOD2S7JJB
zudQe9mSISUcxM8Lf/mHNhunMyeVOQdy4TQGvx3Lgs2ICICiiVRiLbuxmqB+5Wwi
Vurq/ra58R+1cOWpGy0Mi2gyMThrFpszw0dNVSrMio742q7NZxYD1JRNiRjp05p7
B1Cb5POcF2xa/HCofdk4hEZQnN4Reyp2FVYBg/LY5LhmadgCqQdwS9gD+UWrcPfi
CC3Z67mff3NLm4CRHZ3ZMNTODcTDxVNEeEvt0MHwcix2w79FteU4m/+sXgV878Wu
4Yxqazuob5oWBitzYfI3fFJgoAyOa/i/gxe/CIuNzbrrYw980mY1cKtsAX60UIi8
0H/YZ+P9GAuuLUutf7MutP6pQu2HS1lWtKDQb3sPKdgT0reO4PePdp5nwMfMKALg
uJVNp65bfrRhBlzMNhAwKq+af8WfKsDakZD17keE+hksTZxYDwBc53HY3Ux3DOkB
7LeYwif6Pslq+dO8JCwguA4nJG2nn3ziMs4wD//XlzUwjrb2ZOqJzxgnYKLoIFUY
bAOBWEE74IA3tw8X94RThduak2VhCiqC3YfAcgRnemaKsDUcCZS0RWBZleVlkngc
ZTQRicW0M/fL62ybnclyuCKwJwWIa6ubbLt85afKynTacTgvMerySqMYSpQo6KtS
FpauIM989jZM4yXDqQCkQFgZhWfts/m9CJ0z52K1wzY1yz8X3/a5839DR7HRRhAC
PFi7NSSgmdJGeCUEJS96QXRi0oldIfCrUL524digFAf4Y/8NtEWMmATSDvfYHsqM
EQk2ZR/pR1m9TRO0G/XX/Icvr9EKJrNHvLhJydv1g3m+Ws9C8M1ckydewD3UVQPD
4YnQhJm6QjdkFm9wdefJ7WPmz/r94LjhHDhAIDYLubMAurtA/hdDNYMpRdGnVNUN
L5AQD/ea6WkJYUdJnekOGK62h4scTObCVPKjLTVKjDQ3Qp2EtMDbJ+7J6fXgqyz4
dZJXzNI8UwrNOu1RkODP+HoymTFmkHMveqCsc3G54AM7x5N9eOkmU45nll1d/5Cr
oyHZ3DQgJ0qC0MfGgb98UoWWaev26Bmfv3uNpnVmw3cN5tsiQP0veU/llKOU0DoW
8uP0KgcapGnFYgqosdLL+P9xH+ILIEEH4Lx3rGmOGSNlq8nXwpgch5oOKckNfErY
BLEKeMml02T+Ag08rWoz7QCb3R3I+qVxP5xhh14WnA36xJ6wLj3SsiE8kP5v/ner
Q92HeuCuj2un01MJzfQNlzK6VtJ/JorsZamknUYdYb4YzZH1KrpO5oKb34cr4gHw
ecbNa6zIzWCKuPnshuJwgPn4dNKfSDtUptiZ07aF7XXOiUcSqKxSt58fSWjvoJkm
VM3uc1OsGuTgra04l3RkUeC0figUpIeoGI7F1UH1ACrfGuxJTge65bmuSqNmIGQX
8a3ppKjSC8li00Bs4dk0czgH7boWLDmW6wx/2zhM7VL0YrykNUk9ZS46eB136MDP
ftebBCgBbg6m+uCWODDmZZksamTebF7/XvVIjJh58B8bjGYliTsg9hOs6BQCJyLs
K2K+tcN0ioKuVlHsOqOxiCYcrLr9WYiIdf/NdvX0ZQZeaayzMdIGT76O4AQ9uGc5
1bTfW2bA3UHj4cUqF586R4NRZJdEI9KFC3dArSra70+vsAXdkimPRj8vZOPyhXPN
3Tf50OMh5+hu/F7JB2thB3ZBMqO6tbxrVfPqe7l4Kn1ibLwvbj4LsYY/rzioliKw
CJ/UtNfuyvdS+hxmM1qzZUoMD6ubjEbaRNh2Ofzlp/jXPx7wcLK2HNmoziAl6xZv
5/h+bqghWKKDrmKfFwsC+T0MabDklH9vQkCx7dn/9RKuYJUr0spxKCGRDkUiul1Y
17INEzRQ1ZkgUgj0cnAdY51dn9NurIlzCScn8Hk7140nR7iisETWtbWC6w9TI8G7
+viuoh1sYnXA/+vDWTUYybXt9d6sBKAnUiYvNS67jumW5GfzqCmOjxlhSGiEyGP+
0q3JP7znL4g+YPGNk+PWLQdJKPnO8YgAi3pqsLoq4Bkl8UXUu/XQCBVmcL5hna8F
lldvGqSPgQHVI30jk+at3vnlwYlXMZEBGnYMdgn37fHfwKH0XqSFUSiEWxJ+TXoS
Xf24ABaWcEfH2EcTVaB7BJH7HKaH2ACcVrkghncl7RXYXlZOWsS09CUwHXq+5IFS
xoXiY6YL9kiaaDwW4klHA7Aq7aNoxx17gsTSO+gx5GnqVnQLyiCrQf7HUwQH5sii
d7aZrecFA7Y11HoUF2zVl0OARxjw5xh0IG2Jp0dggvHukirD29/38ozYHK7+3QKn
v3eYVAckVtMsEb9cxRxYQFIdPhaM4skjrV2Y/uhxSGhmwqgnw1AkqK4ZGShIXoxs
eVo6ugL9pV+jVSvjj5x8jVOL61bAAsin8L6f1NcsYJuqFGJOY7fkd1dQ2Q052v1o
C3d6shWz8kUVZ7HE5RZCL7HYLZbrU5zX0/9+F8dRC+ofXlMV7AuRSWgR1gI/addd
iXlVl3QMDuG0NJA/YTfOx0RFfMfpg5k8k1o5UtWqanM7QYJlkltGEq8y354vdrP1
uIgLXppUmWR+1+K2RFKbGN3raoSncGCLM0U+qZp29ZhzVbAMTV/2q5pw/3DEwWz1
mrtYp2T/D0iDoMyvgemFzHKRbeXRNKBe3ZBUTRiW7Ttg22X9ywNkrXgwqp7oGZ8N
6luJ2fLQ7FRyiG9ehPixV1CkT91N7lnB1hsgtR8p0LBfPVqyFdPG6A1dkdwfrEmL
eRVmRrKe5oeeoRhKA0n4MU8RNn0GMbe3zUfaLVX3q+m4kvg5T39oiaTYxsdXjkbP
H72D7kqHLb+DNm635x730V4sAk4DWo1L6f238NPFO6gvrSJ5uiSd1IRM0yAVAFrJ
RujUYdy72TIIAB7dRAgKFyrlyXxbJJiti+fhpUXDtBG5nT2OsGDxMdkjl1w788Zm
Z2VLirDlG0D2DfygiKzZV+phSL0txO1zf81kFkcIEVXH1f54LjNya6qdITvzAxW8
QZMjXki8X3AqNXGQCOZ134l/oF29Fn35QiWVwXPPixPcaJJEX570ljRsQMbqidvm
Wvt7FUyvXvwsoNtppgtaNtT5zkooJmwsYnnBEOelkJYdpfNhU8WHAKR7EuBuXca9
xSrrLjI0qhV/wfLWlikC1p8TqIvhkBiFi4x8IFXgnva62VH4KIOYKXzitp/pPJfO
K92o/Cxmw9YWgVUXo7p5bTJbmnyClUDFUWmb91yye9hAwfCn52Me5W5C15gHSuDq
/NCQzOLu4Tg+dxjiCjmsdYx2R+5/KnauIdDvIjMrxNVfsI7Co5+Hmt5kkhSDndJE
aOcQ19TqV4NUhjo14UyCPQT7qb0Ys+AhvDV/Y9dZdP+ftxO8J6kVyIf+Ln124emF
V1mW8NBpJGVdfjkKmYhQSXsPf1Q3B94u0GknDnE/wCJ8RyNY6HN44TcM7etOa0d4
eMHxaAKJ0GQ3JfE5ljxJ6dyUktjCye+27UXZ53YjY2oUIDPeTCS2XBj4FzmVbk1o
t6qAe9ntadYlFbIRlJNdO7G5K6aheFMOphyoUt17jvi0GWENnt4vHqb6Jcl4VOJa
T6lkGJLg/cuedniODaaudUw0kmZsMCwRGWoULbVBzAuwi89UHvsxv3t4H5oK9cVc
/5RD+NVQQKH+ScxcKlOwc6wv9sIYSlUBR8wlBRTVU+Pij1JAbDfk7A2JlfhYmD9r
2T/vUHIwqde2z59L6cZTVf2Wd6Gl2dZlyb+g1Ln17h2X4uzZsAv4YW+seNINacGc
2Dv3N6Vq/3xY94pq74RxZw1viluy+ARRP618wzKTN+3FKdimEmSFv2Nc9sk+WHZb
ryaNBvrFtQ3xwlYH7cWWM/lHW/TEenGlCWiMP6BzTzL3YOZtFk1G7synX0iJwNuV
skka5b2yXt7+J8/+NBYBMsHIBcIbtAoIwGfO2vaofL5L2vF59jQEIM719Ih2GDGF
aIvWlZ9EeIWIPbJyGTpYFZ6JmtwPe6osyxtrEQgtLkUG3iWznk0+k5oRC1UIyauq
IDo16PNdLM1jkcGLsWKp/IujIBXl7wSO1lNhuMcO4vXCEmK+oTvlV85p+GP27NvW
t9YDtRlDEp/PjT3E5P/vm/0jEFXrZf0wMr1eDRr6fWd7v4u9rnKKkNz0opNrF/Wz
q1Lx+VYdbZmbl/JfKaz/14UQmSKY3UmXF3Yis9mfbKFbo9ew97wolKqM6xjZYjko
jGehyTJA4Hm/8YZTk7scJEfmfaN+qDZz1BG8c///z3704BH5nvA5CXcl7hgWCpPF
2cARzG1v2kHcuyaxZCEmX9gp1xMaf14K4AIYeHZmKfoTixExSSm7TB5rMDkhZL/m
l9Rz49GqiOy2bR5fRwXEEvLw3tu9fpPjbnks5Jl+5TWw9KsI6VI1csfd3/x5kkP2
F8m/RJzBsCp6Iiatsg1kQ8F8yucKL3IN1P/by4CjacoMzFAU3Pm1DenqJoFBB4eA
e3InreZUx0eBPgFy37HBuqIdkbDiYGwLF1NnrUY8ZgsbxGPmRbA0F4B6NhgKDYUJ
EIO3WBI+LhgKnlhoLVLqdpMIs3usj6GPayt42XtvGAgf+HOyTUeQXMl669Kx2AY0
uRKKYKRQGLy/Dv0l1trICc3NOQV5SKQSb9ddIe9M4Q1b0FbakanRJHzw0HMioDY2
FbL6VcbSV2PHqfpVjXDzaW81Mh1WVL0nFSQCI6aFTNwn/cy5Goq1Mzmz+jXyg1nd
97LSphQMJ8nt/6o8LMKT71NWw3nBcQhkRr0KG0A5tTSvRE2NL5ojwdkjv/IEDQ0G
3xGJdj8ZLPTEcW5yW7ZPzkj5jjm2WuTQc+h6vFnY1rZ4m9r17KtnDHPNJsnbVmcA
GR2M2IG5tb6MaMDYcwYS9KEC+ppkRjGmO+uvxuXJmSFQp6WQlof8isKPNcjsct1k
yR6GB7dhuGtgU19cyPQJ8zNX+3dLLJHOviYD7Ex04U4SbfkyYZ2LBsYfVbdPQg0+
uqhzBzkPK5WUuMy6jPStgsAeOKcGgAF1GYoA6NrnE3/9pVVVjTRF6lSGlxuZDH76
n4nmM4+rL9UNkUeSkGtih5gY5fMVmDiCL6SDapHD83f2wL7cCrE+zNrpeVHeXrmK
Dv8IPBsURQnrPJkvV+DuNzzT+3+8C/Ysf9aHhVVXxtiQbSXWqKvF3B/ioy2Op85M
IRPuf682YsKQVIqqINHEPZtcMCh28GehaiMs8Tii98HHoCn/FuNURqByGEhfD9Np
FVs+JPnWsWR2+PvCgr7MpeY1JGvPy75VAb3mIujGRrRVUwE1BrS1FRpIHNrPPZAi
dY2LWSvEERURkbqsossq2OyxfiJeYXWo53Q14Y3s5J/BpYSpcnItZSzoRlWr5Z0u
b64rgbq+JcIMgdcQs9HXv8g2JQzm2DnZnXJJrUczubP3kyTgk6Pve/zzba9ircWI
JQMpsc6w/M8CWC9qVsZFRdxShQrpnossHKjMP7EbiGyuUk4MF5KmpRvSim8FzbTk
I0L/njhEdHwCt0q6tGTbmo1JbmMDr9UBNsS1zu/lIXDFhJqW6sdtv0uvsjZYIPPi
mD59h+QuEZPQjMMxVO2cs6h8q2WMhYtK60arPeddtbAcTqXDS1D42K/t3YNQy4Kl
8UK3KvJ7Dj5PJo2W+QSGdJNu/jNDnew30TLysVp0qKxHA6Z61hSdHd+OSIe63JGX
GOwVkr/K9MJS77QxOyuJVm91byYOUI5T7Z95HrbK3gQjxHQ01vhp3Tw5TOwqQOgY
e/HaQBETTwvU6Kd4sYDIESxzplfn8ID7fkcR71gnFuHeufi0vkRccWbZ3zkcHB0z
3IB1sVAV51mcrN9lKGE3yF+y1vjUjNNtTFPFNQJBdRpAu0jG+EiyonpiSq8cjIlH
+LpZZjZx5gk0k9iLeQGjjl/1oA899iwAie0wqNymk6EuAhvhTLzpAPi03yLFlC93
0H70YX1Kc0HkWQA9mnA1N9AxfoXqfa1aann5gklddJdkaaje2pIhnCwPDQAHNLWC
Nb5G02RwK6L4vRmR/UbAFMQYekeaflbu/CHPh8+PqHk75MdmEXcLujqgY8muWRVm
LQtlDa+LqkjMmXHT3HIuUM0pVpnBeJ0YaH6WdeUnWhh3EQWUnYta2iH+xTifqheE
nvFVAecTcOv7iRHp5A8BGjgz0+w2b7rInOOkvjVDHecYSRF4aPu4QhshP+Oz3o/R
LJ9Me0NgGI1X+r2Q41wANRFhBd4ZPiND/oqWGbnJfos8aggBaXZe131i1EqCFM3Q
8I9jVobdCcBOwysvSh+ko8zTSGUvE5VaiRt2HSkkPWogOPzR8FpbB0iRlgdKPm13
PqGcnS3EzHg618YS0vf3g4IAx/V48DZrtjld++MqwjDb51ZHkTR5fk5qPAuWupjw
0Z2lBT67tyi0Qyr/IpzNe3q+JCmeU7XDVLQQ/yrO6ptvgI3ZyJSRqPzyTB8pREJP
YOmk15KxAKKg9vsbVarO99gnpEIsTJD8E4l6Z/wEBOBBhQM+3mWxftKk7wQHeo1y
1AgURswmcP4eR4UXroRIDWeyibtRfHAHQtA+XmcDl/rdFj+87ERvxeU42p34gsDt
8zsPU5DD7eMC2lfxq7PVyO4o7Xe+VPk4/wS/RyCW06IMHsvx7VXjgy8RxSndvXhF
QsaYlJg2YDEySG1hlRgeo9Lxk4Tg7/07rTN5jMZB6yAi8BE4u9+sINhcT5aco691
7OJA80eLb4fg70/TAYZWsxwLjOjqxbA0jVPqzjQosFs8r6wFCYSp4eKhwpMFtdC9
klSr3aByvQ7betJ9Yuomrv3UQP1q4u9iukjvC/hcq9E4ez471I/wfcm54REKj9v+
5rcqb+6mWH2A9I+/gTXXbdHpulJDEqYv2G56lJtmEI/s7WHlcqexy3D/QpZHEuW2
wSL4Kl8Go9TcERnNfxP7uorObI/jfp2WsYA0ZTYu4nNjbO9aKyGbGEusMbCXUcUR
VdAM52l5CXH3yBvavtkmatdl40e8mXhsiOpfV6xCV8tGA/knK/ZHPSZcP/C2ovQ8
sSfJyd/qyRCQyIye+AqxPFLDEE5AG3oVKQ0OLaiU5YzHEvlhuuOikbH8qRGwGWvH
FRjIjFGZbom8Xxa1xdkynC4bGyVLqtb3FHXBZmQxwss5Rw49izgbUU/Vt5SskhxX
YwkMq+RsyIGPXf8dmHVh1QeBaxjNz/tRXQM49ft1IIohI64q/8LYBYkATfovkIMD
69lZgPIBZz+fI/y+MfYI46xBt4RpkhVs9omdG/ISMV5IvD3pPRv7zqXibQ9IL8St
VrRZYEaLOny27LM89ZGhjHEjI5pCKrMeC6Zu9IJMGhWqEMkdhtj+0PRJxzqGcS7+
rVX4UA3J/x9wNYmKr66OkqMYIEo7DmWN2aDHmr+YX2bAx/SjlNDcFXrwNIO6WX5H
IqcQKEOSXfOnqQnleGxN9Mg2db0U5zvwuqgbcy7umDvS7BS4HkW9zWUsABXjm+5Q
4EljupgEC336RfAQMxxT8BCgkyeMDrBXWw7hIaeVlD5vH1utclzZOaJfTOtn1X4D
0g1m1bSxUyOfLaTWj2dV+EV8Qv75azgYekgXPVgxeWRBIiS1jtq3DFThpBDMhlAM
NIOCQpYlZTW4YBtcsH4MbtzYrs3T/+vCd9TVQQB3OEqYdWahMXFCzfVh3lxchEf0
cXrtGbfQkcEoRGbXsDlFHI36hgOlgNd4XMkB5ziYhcYvK4UqnwSeIHzq0kihzPl7
6SAOqs20gwlSwsT9eZBRxo2455ss08Yi7IE71YxECLD8T62cKS8y5INZRTm7YCy6
14g8WiBhNjFiyxwONwwpFQDSF+0I4+3PPbQxjectOnjTOrNaCd/71QojfbeJfmPW
SpYUVqvfDG06JqB7I2D8ciR7lfp34ukpognGIZDqhr/ysruwQkjVqr67rBI7rc7l
EElncR9BpKUeeOTFwFPdDC3+WvtySEIw/aXOU07KCEdLfd+xryIElg2kj3QLhrIx
BPwNg5Aw99awGT7OT/E8wmJp3bdbkhTPEAnaGWGJCKEAAwBpHNnzYLqvux1TmmUg
lByUO1WFC+ZwRu8ezPTI3lPyin1wzpogJg7pSF3AjXLbT5VcmP0tgS/QO54nQ6Mi
EWLz+mWyNMgzuhBfyY5QDERgHpIHe0plGysS9S48ljEMwAlXnOkly9o7Sr83ouPd
WvXSAWM6ZtsgCfWcc07MxzskVh73FPZW77X3ttFVMZiI6fnjGrInYpuNyBen5ALv
OxKDjKch2xORxGe0m2ypqfhcCg/nL4uc4pHotb03UfkgrH5R/04pBsRzrCDeBDnF
F0aTWBxMFTQHA4mfgZa7bUq6EEDj8ufc9bng2kCgq/JPVCZCH6T0l5zGO4GemkmX
W/zamBiTeexSTglICef4YbYBjndxjM7GuzfUJbj9lP4U5ycQV0DXRLd9KRunV8xr
inXuAuVHkbm79Psl04KBi5yk07gmedrJs2YlcnekgyHq3R1fMl35UwrcWId/Lroy
yfs1/kYF1dQl0NfzZV4p03HF157vf6TKmPG9b1+jIhdIHoycZukq0EHr3nVEU3zX
yYM0qmYq2yNOAfyqg+6SBotVDLmzEDHA7BBSEacACqD1f8gKPGz+1kcFihzOOesu
EUjYN0n5ADSHcfnyFoLRoxndyrRK/HOKA7Fca88z+PV0XPndwFJVM8fwn674NsPM
Dzf3YFsnkJ1SyaMEOLQAt0/upFrXiffVdJ/1lecL0Y86iTJLKK4lHdzfZDllDwhy
uZV6NYEiEektYGqlsum8D8zQcsph7aZ+b+4gsi6L/5Q2idzhwhpHLwQrIQVcMMo7
f/ZpbvtKaXwDPIJBXZDZXMSMtNXjHKT7iuEPy7UCPYYlHOAwNe8cYC9FS0+MDX2z
lacFx2SDHR2PzZML2YckztrLmYrCy+2PdO/22HF/zfH+2vIA7xDTijVP4bZMi3ja
cKaCi3z33UmBVN9oAWo6rsNnTASgEg1Z7vjsZeCGSUhkYvm0okjBPTDJtBkjdnjv
ZbmWINCyIQMXIXo020woG0k40vQisr2gClML4vwdcA0dvGHtQYgHYfy3dgoE2FQO
DQP+DX4xnwM38NL1WDoF4nNv5AbOFEcfPUhYBHdqHe1WvigPtpOrsnU/ROei8J8E
PGxpp/8EZ/mqGyqaBln7YppK2J510up2M9dvDkMZwfkOP3qJ9yw+8IlvtmBvO4ek
p+9xBzH815BufG9h3lHGqz1PG4WcEjtMTcj9H5RblcanU4mLFtiWRZ4FqV6ru6lx
caOYo66ArWryFiqCJ2m2x0Q6ku3DYex0/+vguvwAJhTX228exa0/ESH47byy3/HB
QGj7dZR9HscY9Pn1DYmUJTjaD1FERMyQVF0Jd4XugA72TX5fYqDG00eeO+h2utWy
RWuj5VQcbdtl8KNb0e25Gk690RDnmmdklLuGjDuFMw1vAvyuVoP/rZu7Nys3CK4V
g7vKAWxYp8Xs34TSDMItIrjA5lqzC5yLCKkOdWAASne0l6Hs1JWcC/7C57gNUUqD
dcDMtlkdvy/g9MgkRJcbqZFd+vSBxciMu/L1dNWPucZdSvV1QAII1UbBkjmCu6YY
0dYX4MI7kwzqDBvchYjqf5FgGWavnqwNlRRdGwxwbAoe4ALkaySO8gSAjL5V435K
xPpHXjKN/+vz9dEOsJcgrxwXcftGC9EOGCQUloXz0Om/vTDvDJl7ypeFCBKm/3D4
P08VP8jXKB/L+OnDKKNqRqCHhM5JtIYNhC5i8GwslR8glAbXdDZ0zNFRV2Dyajd4
ktCyRTlbVUdIAzSVRTcVzHG0UDCRmmFJJfPXSO6WQ4zg8gi970wN6sCmIGd3ZzUG
NRyEii9fYlF44J9GdlWrHMWmdOPZTODyOiVBnmGvyFLlCqDr4xZnjQsHLRBLfUgF
nrnqLfwRTzJWWzvftPqc8rEQOVuAUwOmJztOtki6oet0waVT1zJppBJHyOmvGOvH
Ajyh9Nhm2IOSljaMkrDi5wNJgqr+YZBYDSIDe/lH+tOcBPgOEfJ3siqR72brv4w+
lCGyH59CBwRPOw46nAMB79TkozrOuZ2RknH2OfoqbTIB0JWx0HF+r5hxNyYwUGYG
3n3kfuEmnb6WnERE6qtZ4sj7/uFbyVSroZkAVpZUc2FsMw37NVlIA/HN4pC6QhuH
LchHUU+K+vAC8RwbbxuoEfwNazLCmVecDeWhsBlkbztwy7c5dkxYufy/H7c4+hFm
yXqLSmMMVv85Z3X/aAnVfX7W8N68yVxQEFuhpJECgp38F3CpDLm8Q2lnPxKeZOEc
jY4cPJw2jjZzWqI9AFQTfq/gfuA7i7WX3eC9QWKgB5TdOwoSxZClCvVJv8QbGZ5G
zdvZShivSX86CS4t5x3nN+WO/VP1BI9BhWJqD7oMXr6rwqvK6MBO2075hK8qJQHP
VOkyRSFFJmIHks/0dPAyUokUyW18sepEu8dLvwtz9f9HQBCpHfOyZmuisaaZch/L
T27MCI8fCLBhHMPGNdmNKOguJvC4MQWn8SRIoM/580julq0c7KlY46SmUOvtlyZp
l1VGzYG0zKDbf/BvQi3vyD2pxL7DjNbikxOT23EJRJbskwtlS6B1ZVD+3tt0p9Y5
uj6CR9kcSUahb3tEQtloO2uEnYJP5ypZPU508n9flLw=
`pragma protect end_protected
