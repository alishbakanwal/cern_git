// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:45 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
b4W+wyibkaYXVW+UKiysCPlldLvw6T+MqumBq3SWhMGI1JVy9kXXDxZb0sF0AS3Y
4z14K7UQLlrLfIkpZEDu6AueR1Beow16sCkjcWM9v3b8x6P98llJq/6laI1B6fPv
uoNdQkHZBUpAcoEPTNvUEHvBRKv5sEdKc/JRrMwh6aw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 74032)
47cER7wh7nNpG2CJogN2HqqYjqhz4ilj+I0Nmo8rmGjuJleEPgpQ3uR+NApEIMxb
4ceM1Sa10C8tj4JECn8xBxEfQyUBs+h8juYK8JWSb/s1W0ZA+01VS52MJ9fNOHbV
JX7DdCNknJ5cPZYSglntuvepHzqQcrOsLx5z4sWMpPnmTdKv917AiksIxlczBJWH
wcCCV88XBIdnmatphdYy2CoEW+dx1gINcOldpTyplgxDXehYiGFA4PQ+jGVeCr8Y
LLSCewgbAT0ufQP4p5u78ZfFM2RR38ri1ML208AUqMjH2Ex+bdD7gekwMa8o3R4/
jM8tE/HviF9Kzb4PTMqlkb6McrC6iOmv2iXCtuCg/JG2lnJatCymBWWBb8z2P8mp
ykW9nu7WvFLY48pD89cRcoSp1wwB91OxdCSgJZZH+Rr2O5GM8cxBCkS9f3mG7xyf
JW7w7ok973MoiCAMmC2tEv2fPZu0MrpHdHa/T1Rey9ajg7MAo5fy+HkCxGsMihNF
I1im2Z+C8IGVmtwDWLP6pM64OUAmXkfGXM1pMNggn02X5CGFT1EQCJ/RQKqcV/il
tFq95JMkPlE5PNCa2IWrh5S3yU90dw9lPc+pvKDpCMiAt/KQqORMXV+R4oNbaWux
Fg8kiyTTRTQKzvIRZLRRH3FwyEvp/kXSEE76kCsVxocXcCEVjfNxgldx778qX66C
SJ9iZYLdAh+PG/uXxgBzY0LUVjJg3hO00qBGNxgpLe7W4cElbVLh7+NkMUxCXKdy
hbz5buSaat+b9M8OWO7WpDJCYLAE4DRlZLNrt8thov0bLRRLkwuLv7+dPskq8Zkf
TjN71Sc96uaUzU24V9iWGH58kc3q15RoKEedXkhFL5kS0mI8rD1O5EKnWO3QtV87
B2BL58v3Zpwa7IRVBbyscNgGXJfBZd9+r/OasyVFY6BfZj/u29GzJ9BFzMI/4Vgl
3DIIbTz25dbqSmctU2IlJ9bY6Y5f01NhwK0UNgWcW+oZBvfNPDwg0kvFsfrXVe7D
/cHgzKweV4p4ghBA80R3iNpNJgfM5wMovI2ON5xI5YeqMUM81YkqG5ACGzZ3qV8c
ZLkj/Qmr3S7acPaJGRgqG2Uckq/fxOsyUvyvt/tk4Ml/QYZ3dzuebd087maW6XJy
cs/x0YlDLEtEKS1u2s9NyQbNYShBTixv647MCZWD7ZetUj9f+kTr/dAZzkaUYs+u
051ckX4YWiK6Mp1CsILjRacY5vs25viDV26+ijKo6zhAnUbW0zUshk3GJ4FcItTu
0N5wE541EBRF/WfSb1qRyEiGr4BnvM4CxhbzGoBfxZj0B+YVOugknTBvUjdvKnPB
6ZejgKkzgmDCSFYdT9u90pGCx2jqrU9GDxvEjKzfaU80aAROB4zx/oSpT/IqQPVs
Q30H+eqhUgBcmRLJ11XfejzP8+2GxTn60jkjJC61Y2QtNYO34TFjTr4//W5hH+jP
yohkn0ZK64oTItUCzFP7AuDvbyQZEh8q7mf2GZ0zSREqceAAsNRHDdIEgfMW2xQT
EKVUSfUsdeBFZjBPSCtsvlf24fUXmdKxhFGTuBne+IWN4Jww2SZJMCX5I+zrj075
8j2v72gycLBeHEM4c7rktV/UueqfdaJQX0cod3JOFnC2UnzPOC3Sj9tykSa3kTBs
+jpenkKLvnC5unS0eZuOBniGm8+hOHJrok8tcxqswCwss5AtFMsEr6QDq8jrj6DO
A3EpAhNc/4ArEHA9Ftmc5PJx7tEx+DA/thUB6WrM07RERwbSLmRyMcmffZwGJxXJ
v5bbjZssKBxbggA7tUELRGZ8QIECO2utyU4x3v1z+QiImGmf2mKPhXYWYj2APZNp
7waMdAI+7HlCar3aKgrFBTSXMme9CydelDG2cB2FbTbj/Ztvw9+evndR6kJF7HZW
zVs+sNefP+0e3uzzymB9TD2tYmvSeCVnHvpvM1bWzjmekuHPduOWE8dcv+xZX3dG
9gDUU3nFnHrInbsRAFoUssjexacyqFuu+4m/uPFqFowe+KAEUDQlJPniKWLz4GxI
wIT4dI0NUP4kmK8Of67iPx0IwtEi7vDhOFQd/qtav16CFpPDXAoFLuVQcwTtGXIh
kFWH/nkXz622ggEjD0Vcs6gZm/vxg4HDpfR8RNsNJ8MmSWncQD4TESIJGm4kt1DO
sJmA2aSfcQ7mVVoy/qp9GjpW7Fj6c/1IF59Xalpi8vGFa59hVj6XycXtc7TTjPvT
DovwEU09HTIYgSNLZnhLO+XE8QIbmksQwZfPv4Cuk/759HCyhX+thWKes5drvAYY
R0Q1m0fvzy58ARAqZfvUf3zPO6tACuyPjR8Wl7SwttJPKEQoIF9nEdIxu7+kANly
BIOk05RNvogVjGWL+c0e4AjhkYjqstJBNy6mK83kR2M+ux1Z3KjcqbkoEdRtCmFw
JVj6gZJbolR5H6su+7Mw/VescPSty+IPBwWbAZ+l8Hyi3Lzc+i4lj9IUFho8CKDG
Q6GRbd/+IW12nhJNnB7tw8YWR6+kOVFiN5hnrGuRrBUumVshpv8HxLCACbOXW4d7
LhqhkFAEgWyiJGb7Vg0g542DJOH/cok7Fw5TSdC9OYCoSmD+RJwwawrXsV2Mc8ha
caKRd7vrE+QPvh6bWPgafV3VHjcFjxFbUZn2VJs4cB9jlGYeQh26WHHihtIhP3Qn
cZT0mqHzL2g9MTKeBBBfECZ29iQhXDXzuXe2G0Oda23X7FC50/mRt+THxmq2xsDz
37QpDOsiq+0u7DdaFR/I26zGwoTEj3115Mmo40S4tgnscC0bwzOP3VR2jdwWHHo/
L8tj9WXPh+YHwcaTgSWX+z18AqcfKdTy4YSOfqLYhbpnnhMtNzRDs2RGWAxBpaWz
Lj0Ej2G9jMjo7+d2NVw7jXlgsqldsKYx8I/gDVP8yyOBRLB/wbYtH+sJj2Sp+uQx
5z7hptAjC1yRdHBQ4eIgSaU3E1QSVLDacaTEHUPcUG3uFvnTFpxZh+kkKC+yZewh
iApNgcPq1U5GpXOhlkiNDfiR9ciUHxIcZAYi3r6lwPFwh9+Gz52A8oI6LUsb4Wg0
Hdy2YUnTyFcXBLERRW21XDmeu3H7nAP61Jf1gjtCutyKSwBDmL0W8n7/mWk7fFiy
aljIUxGLr3r2x8sG4EePxpzsjN2hD2+X3CxbBaWIZExxM/71vy/KfIANNZIrvvF5
2sitVHcLQnmj07YSzPUClGP7yKy1JNVaHlNOhiCm5EO6Crsu5O+VJKZHTOL6mAI+
zV/PUh2V3P/AGJ3iAsLbSARqyIKm14zX8W6Gw7Ahe+g+r3LKw+3oOailUgYXcBsL
Xy0Bl+vqCiapY7+rxPCmOC66fwhyFogGEFANiSu/mwv+wbFv3J0xffFyvJ2uWCMy
6bWHAOBL65OqkW8RUJWhEI6/fdPeF+52EhEkeeubRhFO9/ralD0fPbfcSGCpa+0S
nAdvt8fma4+PYQdzJ9jpuXrQmIyugE+x8aihoS0Lgh53qNh3JlESck6W+hTCcpI8
/GPd849IUxudFLJ9vkWoiJVewbNSgSJDXGoPrIkdSL3UxMev9r2wQAXXkoZPLGiU
3VtC0hXz0frrjTvbW7HT5x5tNrM8iyLSmmuMirr3cQ6e8AjBsQH/eTibGtUJvklv
AKtYO8Ryn5kY7EDYTwcz759EEH7Rv4P1lLhPFLliYcMUubAVhdQ+xy0B3Ttl7hHv
PXy1Nrbni8daI31z+u1RuIDDbMKsl7qYiXPRX9Qu8AMJLtQ746/GFS8w5bc7aasy
zoXugw/dUC4XmY3AWcOQ+60ZmPzLn0bAgIk99/F/DonY4ZVCQz6gmeGSmHCZZlX+
w9z7TiH0s25nsLt8YOQOGwVPs40UZ+ZKZ7vN7UXY1W6ZqMGKM045dd4nVfoUb00l
VkOFLEomqTAcTyfaJFvtywidGgUyBOR4Pc1DoqhKvHc4pT5kJqaupEo6eKtwanrK
cuA2n6IamU/5IYHbICotWHXLc6nNmZqMp7beWtiBxuxjme5cIr/xAU59pRcXPaXX
B5pxynnA0s4Q5chUmj09AYnGZ4UVImu58Vyhja1i5w1YxL1LqEK3nVvK5BQ/wh5a
uEeiax1fIdLi7YMdRccicXPL/jUm9ws41RqlYelTlhvqgfFeSR11LM39bNgm1Cug
koSBdlf7gyfE8tgWEXZBpBz+vC5jeBZB5T4LBNmCRhGIFpeoXEqIEE86UQ81PQJP
3HmGyqAA8EDEi/wyYI7BWr8Za+DgAP9FJMvA1SOrVjOWt2Oa8QpvWHJx4HRpZpY8
0SZBStiYBpVO2pBtp0dSvcVFsjEeNVf51r6bXWaP6/T5k1KZJPxeM/XsIoGQjoc6
u5CjgNRUcSK5sGem6kRjkghe/KHYO5gbkcKNAZrfFuqlfVnSriYYq4mLOcH8Fjaw
ddJc9sNuMNX//ei5joAAfAz7Cgz/PVishOCw5tZzGITETjRzE3Q9737Z+R5VPk0H
jF1B3H/1P2Xihj6AD0MA6gwO6G6IqE8vANeYK/tOGEAbDxRiAceKaF3hVClI0b/J
cxva1Ri9QF4GeaZ+CNvjKPJFLf32q8P+MO22VhMl5aM0tlgxZ1QnOvA+jMJEdRHL
i7d476HIEmLelJn4CX8Nhvf5G1uyAo3Lf+3+in+euHr4AX1L4I8yI+X6DKaPjZkN
h9O8HCCrutZKW6C8W2BRuImKfEz5lohJrNJAtgAXxRUuQPZv26en9YjSspH3OMOx
M8kVoYn58GWtvrUuUzF7bP8tEH4zckHpiTE4octQJetWfb+RCiXJxi/fAmQeOcrD
Z0Gtx0Uwpsb1EZ/R51kkgLb3b9ONaz6ot9PL3FsKinaMBvGXZXMda4jGFR5fKcBf
zAhxrhGzNQUwwHYvgEKIWdXoPDtgq6/OT1Mz7dIdc26oX3iuiN5JKB9/YIHOWNTD
N4m3Kdf7CApQjceU5ZCNote5qNTJOuZLUjr1E1/CXIgP4TbPy6VX92yiA3lP+bgo
5B9WmUJ2rqPOz1Qd/bguUxIxJ9pMhO3rwivvNY5OYAJT12LVqsj7yeglkOAKPXyV
6q+x++6Ij2sLhXvRHiNgO2+2aAo0ppIQlSxoM76XdVwdpfEJrXXCl5dTXjDqNLcV
Lob6FHWE1mp4mXu5CyM4dne6VSH/6BPE/f4n8RAk9FNhS+VAMeoGPM0o7GMA8v05
DFl38461ApPRDse1x7HWciCqvlzPx9W3NcgdFB6SGkOzod0Sa9E4fxUumJqiq+vL
EPkYh8x5Uas1fsHHTWYIMf6iryI6gcGJLNbuZHS5jiRwMtiFJL7hlT0ZWT41OqxQ
RoiTvLvZ+YbJ/rph6+L6ONj6nryHl/91aLQPnJMwg/Rx9wIMyrK6W4KQxYtUcunS
TuxfVXij4wH1xlPCuL5+8ollizVbHus0kjWj3bedUwAS+KOXXaWtohTbSqTj4uZl
7PEIQsxAhkid1jGFWIPCdggKw1vN25uvBXbpOgUADjc5gS/DVGwIdftWF2wdcC9I
rt0sYhv2gbt6gL99PkTBAYYYNBCL6MdPMXN+f9tHk8rtQnLKN+56hISoc4z9Tehw
pE2TRZww9AN2McjPkKgaIKxTboa/sS/+qjtgZo5eVIgh8TeaLqb8D2eSTkRz5kY0
dsZsj4MsKwHNDCnacqd4SWZ5mP4KclhJwF/f6aV3gNcs1Tf4OMVU2Gblxaow8XCk
Sj+ztght0WWRdYDahndhtvFZYcKsgNDV0jHmoz8Ke1GcBRx0w66E8vwpNMT6eoFx
5JgDYnTH/0nfT0x72+EqeSA2Kq7521MVk1+C/l7gJHvnSBwfGPpNPS9bqRCoeUj1
s+CxJcZOjGIPYXvApRJ92qb2UBXLyAqvo/f9t0qgbpSNFET/h8pGminoA5aIUCu8
IjB7gO9FvNMVjaLvorusglXnECjRO2SXIFzTD5bde0Irp+097Y/nnAw4dCctqYjO
Sq9kn+8seGGk4wLmEu1Tbi4kduQ4F7m/iFVey8bQk0jzWUAtN9L3ZHZRM3K1kEdN
2nMO5Iy6c/tPKmKv5PVPaLxtSYD4u6+Bw3X8JkOlASuLtcSf8SQ3gdXAkYGytn0N
Okbb6tzxSRUhxyZLWFbUWhQIkG3Q3hI8tQWPYDrakJEa5a6Z2b4H2gEb6qpwSnmX
x8tpqQFGVJKwmYHSNRwrU/vxCo0SPQWFQSDY7I8Sptxbe1RBKUfwuLEqeaQ09rZr
1adiSKItmAOEeE/74VUMQ/A2P1YKy0dyVHO4alUlgGdo8SPoch3XRkNbxHaiQaVa
ihgF16UQViuvXR2XTPIF45OdpNcgspoIOV0HNmr+9Mn9eSIwOTFLm/qkJG/OkGct
WpvDCc4yOwxxs9St6XKM8egfYkC3aTV/gCYr0BWKLcnPuslTapa2dqMvo+Ey2CBo
IZmlD3/1ctSn1ZStZX1TWXNaKtnpEfyd6N5Sx7sTb6YDtoiopI6aYzZQVf4Aq5T/
J5+5lwJaiOvXQO/VrqLOz46oHyz90SVbuhuNGl91nCkItBZ3aLVpS5COo43Xoa6C
dMByAB7pzura+nuZaIfpyGM0coY8+NPwns1McWuD0QoDak+0MMSFSIFFvGXvFckF
cVPoQUENHW3QXG/ZoZTDuinTMzwkO4EDfNPUPebw5pmjscQj5R9sYZnDaGZF+SLD
NaVBrxji080Nf3/9bYvUCLUY7+8/Yp0GrDN+WM4fuj+zBmHiuHJ+KiPVCQuk2Q3f
ASQEylGnTFkI2lo76lmwouo2QDU0eEs8ziBCiM34vim5pA5eanpyauC/yrrC6MMS
WIR0h/cyAhXRJYvQoJvUldlnkOOhnktMzHIhH3Q5w/tx917Ky7bJGe15cfZweJAM
Ok/bueySpNYfHGRiZRkRZME+n69Mm+rGlubPDKwZgYsxWoLW/QaGBn7Ip1Eu3sv9
Q+rYqbqXAWKW5OLpbHYQwJYXwSGvRzyWG8PX2uchtgjSwbHlk1Mhza8hWoXUUrn4
CnIxk07tQO0TrJtTKq0UhaTVy0w9j/TtyC29z9ATR6Zx8FMm0aK1y6uffdgjRwRg
epo4aWBv15VdR5llhaU5CHc/wAIVa2Lw77rawP9UuI69nOg6WYVSsCnGtfnC/ZLB
z2QbElTZAfgM3P58TaUiFkLBbyBl2OgeCGgdxScMj3610BHWN+XCWGKmxYNuAgu4
jYQ4B/05C0ROvo+nzbSdxTCm8ngvp6yfP6ET+zYlxGF/lupq3/ZwiqO2zNIrreC/
Wwx30DhM93tvzKVva1MbPWaHEAJvmAdCsu9qX2MXCWzeideS/ul6pYYeKB7n7A35
CLS6HdUAUfWi3bjOtHFsHC9qfOIVFu2a7yX3UyU1ei0j+izvSbCoYrrHNSMjFVxz
M43nIYabxvW3lKLTALUAiK64fEBsGihnS3mGTApEBSEo/vZLOk+/4L1EH7uZap7C
1jtubzUP2d9dSJBaOi+5T8OShhyJR3B98lbpegGWj8CA2CMK/3RNP4QOzbt5Dj1B
Krp0PUmRn4Ns0v7QYL9nbAU2aZzrQuf1s3QMh9hIWReUrPyfY3biW7l1FxBXp8ij
mqXNBBowJKCaEIhQqthzc+FXyrDVQF5a3cbTULCKUEFwB71/oyhM79SUD/sns8Qp
6HLCTalHiiJTFNi+VWs8hMvhz7PuPES+kByQZqWIxHkuLoIos5s4uTg/K4sPIRPX
A8QDMYNkkU6d0NQ8Q5Kb3mzDD8vcIqhSUlT2McvPgRfDPs1eD0ec7t1pA4jWWLWB
vl7c+1RvOnMRg36ZdZmz+Jg3AEKj9tmNRpsFeLPdxHLNW/3CeGGuzSCUscwrAUMG
9ZlkYGjBb2giKGse37m9OPa4EENshs9e4hvUybvtWk0jbpsKGliEL2pyCgLhgnRm
dOL466YD8DYn+J5bhTy7hTdSMAxgvAyD0KZ3jhILoJKX6gSwVuQly6qi0DbteScU
33b9qh9YZ2mMa316NsRf5ikXKafiI/v7zNhaVW0s9NfbVxHYsq2kuWic2r27hl4P
k3tkc9mcFRJ7CSIsf6d1ngjRFIzzHlBGrDFOccZzSsrMLSInOSvb0r1c1AKKtr3F
Y6s7IgvgSo48cC6kdLkIaDCu8zWnGoxjpzGb9zKKcEc1nJbXXO5bkMgaZ8wctUrJ
Q+/SXFSjOwEJlV6paHmTwN28LETcifT+xTgj1AqqEzBmUZlE+TMQU026GPINE5h+
xxvQLxlRNiBDa4YDqEtFaUdpJNDOyvftxRRCRFt//v6a3ejq0PTy20HR5gsPFf3U
Zs5uLr/FTPasw3gDi3TR78OTAJpf5nDnMjpi4uWsJX7Lxq25R5O9GfOciCx0tJGt
1pcTWtUjcnd4sRz8Pb+elAzDiVd9v3CRhbrzkLg91w6vg/xm9+4v6QXB3F6//W7p
BGvsZKvKLUyxUTZv+k1LobWO5nWkPY9moH4s/LXDAl54RJTSVfQoSRrx9EKSBtND
F5JKHvxRfG6HZZEZ4l58ftapsD0xeJEXMtjD1k0vef3FHbpYsHWTfVTSPGraBpC2
6HigKlMAUOS0HETvKGk5MDqFqUOBlSjcskRaZ5xY0GO4mkbem0po8rIDDxzUTvwV
oEPizpMlfftCNMIYW/X9dAPjuGmU7WikQaYAYcn90XVlESunQv68sqCRfa9lj1+N
ujBxcteyDOWX+X5SEok8evPMSvBwANSN5eEuskTuPP9EoKfj8H3BETVEcn5F/QIG
2CTx8JogHODC9dSp+KuUGZqv8hhnQzl52blHIvtZBiihrpN30og20R3tCJD0i1mB
h0vhN7n/gr/elB8Unt/0ihGO2fbnL1fXewuk9uRS5fOtat+jF9VmXeMqJTQMRTp0
wRaRONRcT+kVcb1NOsHRtCjUSh3ivYZYgeozVcwp/OjDW7Y6Epiiv+L9hIEsBRLB
WKLXJgUv5gdIXS0axdoN7Lu+BIRAyYnefX/kLtBzVPJriThWNdB4lXpWU/QsR/gP
IOwhmt6wVtmkmNaaGPHV8YPzOnUzOIs7VdSUMqdG/YS6i63nLIzFSajAuNPG7rgf
Y8fZK4pIRui/c4Y05cj7rQs6KU+UuDhbmAhFFCngKKPL12agBRRGqHLVxB0M8Fpf
ZzACbDKN6dCgKrJqexiFAOvGQOSl5PAIH9fCwaLFsG0HA36DHYS4AbBgP5PPJ7g1
N6jqoIj7H98yu4gi2mneNcO4JaQbLmhndebdgWrR1ptdPURjNViPBvMVehH+3Wju
QYfAk4WOF6dXgcu3O7Ccellk8vYMYzA7Gf44OmD/Xda26YA65YDUkk0+IHnSabDD
9vjaxymQf/XX8OKA/sfhK4N6ZtpIJosC+6j0VOVTTpfLm3eFfha5SymxGVU6zaPu
so0cpuECtHcy9D+XhAW0xMsnGvVSiOG9/CjqCiceBuNZSwZofBpSIrGvBiOf7OTo
iMrLrcvjK1fNdMSQSP7z0sJGnjGqL5GPN9sBAzSb17fu2+Ez7rxJIi2pC6ZzjahN
2nzpso6qJBCF1WWkAzEHH0xdk7wHOc/h7E0e4+QBkP3VHQUl9N7fzCUdG7gCxqlO
tzZgI5jPCDsqqDWRW8C63o3tYZX3MixDOHejJgmPOLTXz+CxAYJ+BNJZPrAdIzY5
0l6Kc09BIJ/xQkBSFJy8RIK9X5EwIjf98Q5mrDHBsT9iAGSUBq6W2DM7hQ1hVs4S
keUC5c/O5rqfVoijN8eP3QJr+Fww62GRzqHfjI+hMNDOP2nEeCjS8Pt8QnDLKECR
CIrQS1y8y0j9aN/Lo3HALbzxabRzIq1U2rZq7AFmJsxzRJckHr04AIpAz2SE1RlM
YQSTuxXaoP21Vy68Kt4mCwNTGDHwLrjRvtOv3Tm/jzr6yrbiHUVyajL1nlSlnM9G
Eu50oz+IRQXkRwZgMs3sXH7J0Pnz87AZm018VJj8UOVyr89IxIBTLE+cfquSYfO5
n5AFi0aRbpr2xdwHAk7WCl2sGF8n/mK/PtV1IOM4fAyWr+eul6wb7tsjqgtbprQy
OeFLckb8urqvICnyFNv0H33eckY6vF+4LcKq7aCGB9qzcYml0nHBOgPkbNUTz5Ic
N9FPHOIWa53nWXsOrDOKEn8+o7rXm9WXMsWKWWGXGZNXRwXwcPc8qwqWSgbA6YKI
r3VgTATJ4OGtConIinniXuMaFs75T1KhmxrnZ/604+/WnslIMdCKYsMyH7LghlSC
GasTR1qDMKBWh7pSIcjfbTpqeLIKSHqfmr6JiY4WACni2VesIW1X/Emfk1nvk7h6
9fzGS8bCiKl9c9h3dakJj0K93y0XRqfzQ+PGElUThBP22sjXxjwmE8nIzCmIbZUz
ab91I72d5nWMTZMpGaUgWC8XDRZdyzQmrFfB8h8A8LAHvPj+RE85QnjnQv8VEx6H
5uVYO4YxAAwWF8qP1lqhQZDNm42tcDLIZNn7XYjAfBncl7uaYm+BGjJVwn7BeWbV
R12Lna4y+0LU5t6VMIYL5E6VG8KQcVj8do5t5TjgDXENvkdv5unDVouZqbTyWdOX
tu4nJWX/7RGfHGqqXiQA29rcvt2YgNoaOrxVXJx5QIcjmOMjPXzTwFPd7Ge8UsEf
nbX3pVz2Kln5XU1X3/AmXidjwJn8JxHVzRe6zh7DwCoWdyezn855LC/h+6S9tUZC
ZfA+mZ3z5O+5Xuz2Xzx6ZH2YPQ3a9TTcBOYy5HvXBiuq7xFUu3MPLIP8FnDwZsat
hgZoG0ZTeOeE0QZZAD35PZEKt/SThMRAl9zwddItaH8I2bVj7Rw2PtkaIw25VUr4
+IO7sloE++gKGtjNT5ZvKPs6lCdEeSHP6ievHTnd4VArxIfBFMNMieWF05/sZry0
fOEa5FL420UtY9tjCiiGOy+R/PhlMgbBBDjDYZzKM+6B7/uUG1u87fnpqQia78SN
LMPj42sBoacQ7G52G6iZKf770OG9n+LUrmWAVO1YPZOUvfmtsA6YQCarAlLHz02O
7KmFiTzIXyfLLsyTIlE6gSzTlFjP7fSkRFdDD3iIJl24G18ADLs41Rbg60MIr2P9
l0HzL4lrJYGqgsaTqcJHpqz5HsS+eo+QjHPcXPelcZ7XtSKnFv5YFKus/F//e7KS
1Wfj1A7yxH53uubiw3Ag8E83jHFXPQzKBxbVw2bsixATuC679M7xxQohEaoVJqjf
ZVF/rp+MIfLXWo4T8sjNA4TGSPrCBK1d6O9scAWVeHbDJRm05WSWaH2+02tHGVvN
NeNduU/NeLFMxF6sJzyomezodkqU79H66PseqCLUcLWaNSoUzOoNXI0pzMA4L3OY
BIwptO/mKxxNNmRB9qZxLct+UgflqDDOakYXfTHu4fx4EezCq/tTSoIx1HTznE3u
nuF+sRtr0a8tN3w37km/1WnX4h8PGDYz9sOx68NnZPnI1T50Qvk6cTReQiA0ktMb
LhkINg++8Kg0hErrJBeabKP9MIBKqdg6/agqqjW3y5gJlt8EjvmNv7A9Dcm+8bjF
8hClTmrrte+FFN1MsHC/CiGAIMbNVZHxu5+s3hHVPcP696SbCSPtE4Eh5etR2hyv
V//9dBmUABPKqzdAJaB4Eg0gN14eYnhnS2WA9RfgNTrENu6+t7REX7SugOfLyHqn
zH2uDrfo9Pzd13Nwo/WN5NG1/SccDfgPw7zly2rZoFpNq0XB0g+JZBSe6EAenhg+
v6RF6QfIRdIP6ZlwKGzbFF7Iktus79pUGT1ZXtt4n/9kO96pjBCV+40YyLF9jEZJ
Dbg5PB2gy8Y2FbEsqRP92VFB8gXpRROMC9uI7DTOonqC/aZgJjqtwH2dCcuzR26n
it6nZkiUK4FjJbPTopMIWtNi4GCUkThy5IpMgEo5s4rXYe9Mgbz8xsd/jezPJMs/
STRdWjG/boWKfqkdRVp4sVIuDc7wYgZAZ3tGAng3/532eiDsVYuIqC+sPCoHiwUB
1XhuI7EkDbgOqHwz3rm5Nxwcj9RI3luin6EjUqhme/LMYcmSkmM2QnWxm+dWd/Q0
h0ZywlVubY+EmCIRZrp6IyUuH36yt2cwT7FyvI+lvxDI7AxqKxWFYPtU6+XwIT9j
cwIw1j9OnMBfWDqZSgm8RvIC4cMG/XyG3x9dMNXsN4544zN9biSl0I5SlghP7aLC
fWop8SFodTwG/vabI3iDBHNxPX0fR0g8KClg4hScEQlLalo9q1YcdzMBa8XURQVK
J6z3Qu4tvSNQJ12BPAIH5lEXWIcIFzj7kEaon8aHgPJqwG/lVHF4u0JE0p2EddtP
gYFxYRAdkFqKEJzzca/jYvV/eDNQHZy8U+nKQE2iYaXAFCD84KnTcUQzRP+h0oq3
EuWckavexsBsuhqCWzM4WcrQeexj95fv0bnq3Fph1JyonLiZbxepOXpRZZGzCB9c
rXAbikQeVDtWhxjM+wseTBEjmdj+8Ps6+YToBv1n2FJuVWy7PD7zTR2BzQOyc2d3
Oe/v7wRLM6LNCfoXnTSr3+3C/n4xx7cdVE/jz+Mll2lOOiIW5XFmLjryKTqaTucv
TDLyAIN57uP1HAWe3RYjq3lqnWpIAUJKzB2mnHNPrCog3E0qt5tPjZjMsbGUsof6
CUe7pCJpK9NqrYYssY5fLlJpqkZcIJlVQm+4wvd/KW4FbPt4REI3q5GKjSOtIJp+
FTspk/7xe9e9aLEr5w87oAhK0GXDA8E78gCBcNYoNEvk0+qgyR8kH50m4Z8thfxd
bBePo9JnYZZWB3ufbRSKwHWEYJfRkOzywjxqb0znFKjuSihrOEZ3WA2JaO0XSwhv
DA/mpTc0vhwBocxRiB27PWNN1BR0+nIkZOR1uptjOWi41oCeSbR5PwhAkhlWl3pE
V1IHRqVyYFfsbK+3ct9eqhXhxNi76AD8SfgKmQAvVjDoa2HEzbyrWMQuOAnwPzTN
HRXBa8wQ1H9tondvjECEXFw9Nvh56XtW+4e6mriIXEfaVBpMPCq64IzwCrQm5mIL
Xw9E/8vNVkKtYHojruN40af/i/FsbTWC/JqHjwy9tkzri/zateWqHsmUMnpvBfZI
FG0XttijW6e2IBEQwDzn5BKuoq2YlycdMaQRSQ97LYJXN9R7sQ6KKAwatN2c8QZy
ex7zcE+m2g40IZxmmMpytouUSVn3qft6SisKTapB87va5rTqRPb5V38RnQzrvvwO
kT7FgYFbNZUREwuGu0HsH1lOJftXNbLmHdhyOP6+USYZmd+CGz0Fye1/FVl0mP/3
ctyFwaiVhtiQE99pp/z8RiZJ9dyP1oPrQt6yTEhaOiauo6cst4aMSn6GCBxoZPK1
9kvsMGuFRm0iC4Qq9tCyBFWNX0Hw62NzB03B+nKCFQj+FAeUHBVheDYldaegQU7y
Hq/uJC74q7sqfz1F9Bsmivu0kaAohcR1fajeZI1S8kLjwGsAZeX+ayoit+dODl4n
p2hyE+UPtuyn06+Vc74AEG53R45J+EUFMKflv7nLuOuzpnftvQa4LjntENtiSFKe
Xvlh0pBwHwY0yNkG4SxkOtsxqiyov6gE3B8zqZhQPdAgfod/I9syPYxbG6tb81Gt
1fkpacJU0gv7Qu0tOsRNB/j1FzmzO0gDxD2TDomb8dwL28T0KPknA+PK7MDxmO2T
AzMuh+HJD2UPocbFfhNI6HuT83TPTfJbIbE23IlkEkmj6zKaVrPEzgfeU7UzjshJ
ylJhAQs968m9anP9cMcTtspAP/xKKFJlXNIndoduyZTyijUCVrntP5FpWb+3a+4g
SYurcylU+XqhCCLCkWOSuQG6M3/KYOz5XlZluVy/n/RwTKsL+WzCUPBMDo2Ns7Mx
VEOGJABY6Mx10ZThZuYYaUha2W1db/ehjUw34Ux6XyWFARQOaewjCCBPbRkKgBFJ
n9IsaTDiya+H4GNO7i3mZ0vJysGdqDTkDdxc/bOZ3YMIOtBiP1UMPFrYKkmjtQQ4
49fIc+1goEqdcM4e0es/dtstE8W15Rpdgz19Km0IzVBW8mEmYeisdleeWiQn8+Oo
fvjUf67StVh48mqFiAKGbgTQvnAVSWVNAh1tjPutu+zxsETnRjz5ygLPrASWGgxu
68LouorDNUKxz17/zOuzgIrfBm1qX1P+5QbDBijmYVO/4ppJ6DNz3dn2cH9soh/f
saf+uaG/qcOD6X5x6Ct4I3ibjG/7nH8I6gyYqdbPljGllhNE8B2XkW44zCbf5Ao+
30otvwH1fD94unLeLBFVrbIorZ3aTpXLUBo5iJMM9SAWXnmA83/Mgk1gySL2Q2Sv
iTVqauOIES3yxk202rKSVOWXYwzjBU+TssJZNldHoqlCnRGeApkj0Qy2TKVi7od2
8WoEoRrTu5apdjN4UCIcasvstC7QnA+qvUCd0YQH5ABLwGFuLI9XuT9/K2ds380U
o3QAA36rB9ppZtg7Pjk1B3wYdCHm5S2R3XDTR8kZFCBHgL5HjEdSZKJq1piw+IFI
HLS1VIjM6Z6CdzdcCphSPjxAExL6191gSWaaBUw0LOImreUdhmdxgJfHcYoCM6V8
pJcKjI5gxqAyDk9MNg5i777G4cxU8VCx+YFcFQg3BRgl8L7Z9ibji63XccvZcM3z
UNVI5t2dVFzpOkNUmkp3Hj+WiUGFVmMFjcTGC58E6P9llwFCUbrQ9/hh9bnBLnJo
ZQKV4T9D6Ea3ArhebZ5mNiC4hsOPM3QZtkpKb3cSFEPx7xhx4mJfgbLWJPF/ulLH
kPAMtnaUGXR3PRaLsVSmaKLepdJGHh0IFzJhAn6aGFMPXSDgka3ZZ//LSfoyccDr
anyLfl4km1qNnjO0tBF866J5yyZBAWuxmfzVSEIaOo9E1cHV1yATx5o3d8QIh2KI
yNBZAyiJKYrGB/ySx3zUb+0l50Zjb6A5rd9gDNjQgbyHGuiGZJ/WwxZ/esagh0OJ
7kTWll3ZDtKrsg7/9xSU/YMrnbhTeduRuXB9GkZYpmuWq96JkuH4+reid80wG8Cw
ruRnqVXN4aZUKqojdTvrU4Y+SNIwlz+gCjAGkjusQ45clwdCf1fSYt9wVdD8Bc7V
rZFpPJWIaEWIg6pLdvs4PfRroYtFEgBAxEJclTtnvMz5j0CchNg4uJlh8vEYoTgp
j2dyh8k8kty8ntoKPTctIvo0Pb+l8k+87HrCOsfGpOUzCjX6zCPPMe5cCQLR7ygs
77jlEL/Gv/MM05Oofn6nUNxMg1f2MrlfqR9nBOjjJvO8zZajdqrbwsApubZOIdNT
qrRuRl+7wWnNf78Gdv3blePsGSBKiclKwQvaCQYGoP4WyQ0dgBbHByMybM1PIgPX
Yu2eA9w8thX13FYnrvi9GRU3d2/XSQIROCoE+p3fp+tVcgPYA0rI5u9dEPxdzjTK
zRGWdLV62hNVMrAV6fxjpFNyZLlffW7sG9gDr5X+wzz2jqyWpaDBj6jG4jpk808N
tbebotglxX6ULryCb57w986EE8H0NBWZrAyruNAGfk+2206bcd2lWeg3MABqngtI
d2ferf5G6z33aZrj5XizalfNT79y7Z0ejCYVmQgvVmprAAkFSfUvyEDQPhxdbUCH
P4QUoXOnTmPvPCwiVnpp/4z8/TicyfRBBN4LZ8fjqC/826MtGl6JoLG6aKV3eo2Q
rjCNfO07vnPDtgd1tQvnN6fZgG/B1GIL8ArJxVN4oE0HbRKEBFsUYmTc7oGwT4z6
i7ZEX1HSWRwXA3sI1sn+mMLi1Zob9outc/bt9x4y5QfI7LfAAe18OHThSw+UGi/K
hNBivG40a44e0X3itmP/udpgSr+0NzFn56WI5PtOh3wlp07gn+nwXpYCoeAVEIbI
RAHKSa+7G4HEZFWE9CSDOuBkCxEWtFbDnrehtBZm8NIUMUqq/umP+vKdt3t/hFUC
Cbm9WJ1KSdX9LT/dRSL2D/eXAMA/MQFNy4IXjbKrYVwMCsfbhLV4v2A+TVDmUAKQ
vOuKM3pz2tQWituq7wkd87xYmf/G6r+c84w6auyqhhoSffWJu5DN64ov9xDVFWeZ
TNOct6cijwiN/ny4iykz6w+4RqC+8Sj+B+AmCl8yYGFEgJj3kDNq/vlA7zojnIrK
U1WkIWeRWPiFwaubORS6KyGBDBjNjmBrqjQSRs6B+rNhkroL9rCFQNLk7XoIDCb3
M4EyqTmiWw8i4B+BRsCB84Pex4LYE2pVnHFZKVwzUp4I377+dj0XTvrnyMR+N9lB
O/otRevwCS8/wc+gsdU7EgnXN1RFXcJxWGVqvRQrCYPokEVTcPqJRdSEJpAc3AtN
cFxGPglGSfVOVGFE0UAlo+DOnYDufoa4D3AEbiarZzNpPMz3TEUj9Hh/F6vQwLDn
IroHq2NFhRVxYC6ObGexBYZbNp7Q68PQpXz8BYBIVKfIEwK1Uo8PiplO3Q4mH1VQ
8tpGAAA+6GFUEhgIqEuh5dLZLRLk97wiavAhljcMzyneU7sKChqFszYcl5Iiv7Vc
Bm6lniToH0JKIE6aiAWHVYqHNlIWfrWfc9u3M5vqb3iTLHe1xmGOzuVyD8GtRdqw
+Y/UVDK6HUG7o0NY/gwF3Q3405Y0AdFXdKQ1ntRiSMN2SyDhI+iWi/GvTh3/pZ5F
qPh7IMJAkmJObQmbwBNdQZLaStbcHcIpFMxUmzSHRLuYP8GYL9JH2iIV0YiOzbSN
GIaHb4FlmG55uVj99zeok1d2hzg2HGUyqnxx9QhMgKGFX6kwcPdiq2ouXAZZ45lb
Vnd0odBynurGUjgqXl0jg58NpCm+5GQ0S0GsJUmgRM6rCZjp0P5LS+NHzkJuxGw/
V5PV/M2TVnquPR4ym3DocXkp30Z5UKlK/YeO2fYmlCMBCsKy7S/mS/alEUJnIB/a
hsjsfQ3JkZJ9kasr1eCLcxwsGw+8JhVQQob6cgFnZ+jxcIhnnoSfXhvBHm/dswi9
41Ju9n3Gky48f89CIppda2rX/HkOZLaobnGIyVcUv8V1rOemFciUwGRCg7XVpbRX
6GC1fbiuwIAAIW6GbiLx2OOSlsB6rI0OkqNMlhpJl8imjkKeTF39INI1+w3KiemU
U5mDxPD5TItEepTRWpI985tpY5PV/a6yKsAhrnpDPEbyavqidbf/WzNPilkw8D8P
IkZWkReKWGEK1ZaChqZd1SQM2ZEh8OzfLbkuiRigq/YxK9GS+Mv+O/M65bXfw3Gs
bUF10NSrPENfhqjq8xEBfqzECmGRDXX8C6VL+TBFGpBx7XzOyn8bUwmQYbOd3/LA
IkDgH3gggZRK1TBhE9TFUVAWjH2xGsPKrV7FoGNhFn129pWiih0leR2Rl/WhiCdB
BYZmbkIKp7XYLOcLmLCjlfIpoVMJnH0P36qlWYzt0iKmD4Zl7zttcfoFRryTHD9u
kihzk1JZmG3z0wUvIcngL1rciSnsMI10BqlCrunV6Jbo1VpCCEex+qSaVd+BI/JB
XPm0a/qcwD5IHuoB02riRaiDMaX7UIVYSPs7m5zBOcDf798OTL6CiVMq3x+KS3sJ
nN6QPXrDT1w9vRXF2gT5o5n6obKvG4wlJvfMWwalwikL7LWxQxt+z7+px87wO3EL
VHlGhYCp7ZPINoqacLX1rY0Cr7VxZbNA2b4vTUPeMyxFWhF9brxD8hX/Wdi1XnfG
QNcw3V10vB24PdvfABKzSHwaAY/70+A2qBEXdUKYRmhwSvUQgwcQ1vYj2MBJ/+Dg
DgvPhO2jMfNPpjNLgq+Vn7HrtgC32oDTaI2W6lY/RwARi8+BgwaBizH08Bl+CaZT
FE/BfiwoVgaHs5DwgeJ0APtu1PDtLjx2i3Ris6EA2G2tVuS1sidtQo6FG+YXB+NG
7TYjDqs9pwj1dk0ZBcWjFHDzg9uAT6gKvt9KF9gIBRJH9pO9yIGvp9fXECHZ9OuF
UQw+KncCnnB+wUTYxpYJgQUxKxqKl8ITQTCL5TR8C5DizeOn0Y9QFDEuR1zvJlE9
pNu3IVzyK8hhva4iTtzUK09dIPlkWsmC3wJLaQnn1OrPSE8GUSRdY9P0RphH/WVg
lRSZc++/k/sJ7ADVHwvtmLgOdmPiIwQsfN+aP0uMAqX3sPPqwpiL3b68dviXtuKk
c9ZvmGYOWNIepPFhRQ5H51pYNkEurkwgDNKzdmT1C5k7TnS/lQCEd7OsQlS59JPH
9AuMbP9QQT4i9rRVMWL+3n5PXZdhNcgy4j+IEwIlVmi/0GmQPQxVCGW2yhd5bO/P
VAwq7s3SBOObu+bJ25NrVDv4RVlsVFvPQR8nVSd57MtiOllWf6c7IGHE5O7iP+hh
UiQMbqRwglDcLkOJogRhhAop2AiOM7dXvuuWfilaQZwD9pu6d61dxrr+urVdR2s+
6FT22iP9Hrj18nKeeGJzKwPkdXaO9h+tblFkvJXYAG2n3ao7NdkOrqLxtLTS3k+d
0dOgZRo3rBhkFy1NWAVrnLERQU/ZxBz4YJDV0PaZbqxCcjWIcc2xKCynAa31aQMc
AibRLkjVcgYmC4+gxN7J7fL6vHO3a33iMOGlVKa5ojkT5ZOOWjILhW2mEJgmgr3I
0Cdam7Z/FLa24vCwLxf6oJqa8rslGy6UpMo/FbMByD68uZH3MYN4GYPMwocDpQqP
mfQmCWrOu89y6QWBHzePrsC/yrcYGM5KKX6W0jH0u9WAgTFFmZgUKapTJUKlrKus
IEm5UpMuy5zWdn/+1Jj7pAOW04edD4I6luLr6WahO+gzYAnYWvGgjVk2iPVDE4LU
p5JUCKacswpOUjXU/LKKnNmU/oji4fh2qDS3rK0fhxEISAfJo0rWRyEoaADAIik8
O070psEgA6c7bEQTK1aNte/DdcQ0+Z8q0jrKWDoI1bqHu03Zsy9TZD+58SlPS6Vr
XJgyNuqLgt2IER647H2uFSzgZa9A6OltLFlks8XOl7iIhWEHn4jaJeVlyIlpIZGk
fdlIUHwRz91krPEaykcHS29nEgp3mXtNrJszegHni1mnMZqZFuFw0nu8sfwTfXkF
op3WlvFmJ0NydTeT6j8yBUtEhx0UpMWqdGbBj7ZnanhLKDWchxnCvmg+d+KB1LFs
RHM+JXrVo70mofJK7nPMQ5AwgVPqts6deDsHihkiS3E8kLNNdK4BHlc/5XQpf1oW
zBB70yF/tO5AmBOrHzlKU6q8Gd/ZWtVhXbiuknpB14fDJ+fuQJL2M9HbfDBg+oAQ
dBzaZj99FUDvyoVXV4xPSL2BzQz+B0GenJOJrD4VDDXxtaQHBj1b1fcZn3yRc/Ow
3f9YC0WcY0wGu62ha3s5u6nMTvn7a8yoEdhqnbyn0YSnIohyGtXDWegnJVsdB83c
xve79LLBRKohHBC6haRLBQDj4mbHAGStmB+eUZwwoQ7Yr50XdyNx90f0zsMJtIhv
XWMTbcYSyP3PpUEY4MuRQLcYOsLyy5R6P76SdgjnqTeMD3ptUOObqMWjUKeXeh8e
bg4mY1SOAsKRSE+MnyGk+cIPPoVfLeEccjikZqZ2hsY7OvU9E4w1XtijZECfQ/Eh
KkPTctnkYRMwGGdMw2cJBHRg1MEZSStoN3djodBrlbMfBu6XBpEbLtPMA62QVvf2
bS3Yr4JhGPd8AratYeriF2+1nXRS1leHwd/KIekk0jQiwMVO+eFXQvdc3OLUPC9W
u9ptJbdjGi6b9NMsJsQq5G0EDyfUa3Vk4L3Y6tj3lyFL3ByVkbDio6+b99Xl1X7r
ZoP+inMT0QAjz2TsKTZzBhB8Q1q8KtLq57zn2nIBqXMPa0vSL9RgkUf8/Go67hWI
eWVeUtjttAe+PzPR8wRcESwm7NwIzrGmhJca4d69lhm18dIaO8hHXohbJOmPTNlk
KuMu9RzBomDOKrm1HgXqg/DP1Z/+NBvH/DyivTaSYPCIHTFzDvAy6Plc3rU4W/aP
znUfRnsAOz3gYis5XiU6qaTXGk2ojFslLtEHcMFsJ67k9Arx1wvNJPYOPdlYrUmg
lxBWDOeEl5Vccv7Q/m783XxbWCqF6uYEf6jrYpjyw3+p2Y5TuKTz6/sx9ls4OZyz
ZVNE2/Q+nM0H76estQDOSRxIR4XkqH+Ts8RCuum0SN5GSWFJ2BZTXo2FFGChcSU0
Jnhf0Yd6xkYjrTHAU6JUCP9ev8DdU7gosGzniwPycalPYejOsmWIh8+buFUQdA4/
sQJiGI2AAJ7QV7gvhCjj+tzH1aH/EpZfpbeEbv6cVlbhEmw2ndLM9MWGnsvDf7La
AwA5eoRyR4BTVbLSuGCUS8YNb9V3XVlB6lBao82AXOA3hsLDaDEmr7qSVnpyythS
awf10MpLFoIO2eAx9Nl2tLHM0VJ43viBZz/ZEKorznHG7XVpxLbFk5TtSL44WHlp
tQIzpPaxD6RjO8y0jPQ82RxBdTzk0zhzHNRD+PpJDF3Kf+kDxB4T3jvneMeqrARh
FA3fYBqAlxIlN2g4LTeXkPJQhrdjMTodJq+QBy1AMZNJshhptIPfawkpfU+Kk5LP
j0TeY14j4wNBzEeFK46zWaA5A2v5fEPp3aRlHpoE98tCjVOUQWoYg2k3/2L7rc6D
YQPj+3k8UYuYh3VP37EfpAHcm0dWi3GQht8uBFhPN85K+4qMfz+6TXy+IDVVpoNq
AnX0zNVCRvxqJN+nGYEWNoiq6ZejIwtHnGzhdLltiFTbiy32PSSPjFguQMVFSo1B
MZBZmQYrff9EocHO2+ehrbWawVYNBHtDCyWWAqnw5yiLI9tVBuci/C8KJXiShCqM
A3VrH5hucGPvD4CY4KEjUbP/wPv9MWLIuY5XS/XziV+1FxmOjkKAWTNSgVzVsPcA
ph9Aybe7ounfsqBoCI7foIDrCXQsSeqmKeVMfP5R4FhyNIf8ot5TGCsQ/LIRjzv4
3sIVWVjenPFyWHdIp7hM/Ii3IoWTvkVsNai9lQXmk+de7EJUiIzDceNZUwlrOGzi
QQnJrc2wHH4zjBEptM6bLbuXBoQ7FSSA4B45m0oDjYvfCUtjZssIBwetbEfzZvAd
M5FmSKwMb3DJeZ8DUrirSsEh+oZZ/SkMGUwCnufyZ78p4zEsJ1BuM6z3TuvEg+Dc
iqxrmBzZf/0B/8fFQQ8nD0UuEpUq9vkzOto0D1Mq1Cll2FfNhMvhXc0fxTKcaHdJ
DGn32kfGejuMT81/mo9vb+ttdcHJb9yDRJLbt9SK6pIXwrCrFsWPc4p9hUhDftE+
Zu7d5/8Ui3iaBsbr4ynjydKgbOEh+JUtKiTzRKo+Csr9BErGNXVMLmx24nPFqfDR
44poONllZgekw7JSaa27PdxsrZEaBirntDHr+U5dl1YljuIikWQNElaaH+yT/S3J
izrgcXPBspWMvRSG7P0GgrXZU32DH1277JhZyPD3oSWpidFJGIpmlcp3dEM9fdBn
dsueodq9SleKIWQTPOEsQoGS5cKB2Fa7FT/VbaBRzNB2UYdBqRy2uQT4MlsdSS5T
4Fc468QhrmFqYFAMns7Q4Qpcp6JDMw3N4H/uHAzhtzYlkn0dlKernDlFgcVLZXFb
bLZ0Pr1kvWnxOhVMzM0cTeYivU0e+LlR2QLpC4OlxFk3hcAts7UO0nBxYiLwDXaK
j84T7FgeOM0S0+LucoU/mFoh/v8ruGfEuvYbQdHsbPShw4OWkwhcJQIfQNGqXbCR
EdXxQO9JPXXOEeL/1jzWIYjXPiCUzw4S2+jLYqqRtp5Og4FgfrfTKCdkvlE7y/rM
qVBvrNfDFYrEPrzOipWPTjvJPtoYFeYIPoyXLY8PXTRmXa0V7FMVb1bmeWlHryjD
BR41P8ZSmNlPNF38c9EXKxZon9wUbk3DxAoZZ0VPbwh533Mk5Ll4QStjX2f9sru6
T3LbFSu+xvYUcUBxeRaxq12f6HA+UPNMhlUzSMZqXvX6fFkdp/vFREbORgevR38C
ct68S5IQ7cNfDCtcJjniQ23GTA3B3ndy1Rmn2Z46gmxbtVPpbQYIbAi84BkjcnSB
9e9CDTHkU323alHz1Q2BzQqodOHIQUKDOGXF6KwckBHQY5G6gwowL9iEAAt74GW3
kxeFjxIU1j8Q/+YUkSIHRITemflejNNB8tit5WWNou6ftxUh10ALH9fNsP9I26By
VT3FcIZzO+O+8NuXxM0f/17mUMrzvomMMyqXChR5pksf1p9AYMssusqrCWYrorW/
WV7AkYVD0Q7iHTGaFbapI/IYwu3+xhdmynA9N8ILF1YpxmMEFWG+IEhvBbjKY5Ch
YEx0YvLuoobEIhk5hOCoHVwLjvYAgzBPpK3xw3Ku14uacGbWAIm1e5+MCWK1V/3Z
he/4r4uTT2uQUL7til6mDM9Vpdu/KqqQHtz3aHJ5pIBjO9nsUo2TwAfGS/ROiVUv
JqLhfIfRTR6cYHIbNDqY+E9QPUGLeCPbGb73oM3FOzFMSB19Z0k4tTq9sYLLa0bc
bht0VhDxhL/cEgmmJUXcN3cNr2PZ22XeJrb67l6LRwTInmzYQdqo2DWQ9hHk7s0L
UQUhGYNlvH34udVL/2ceLPKQu7MBPSNLKANIyMiBxAD1HQ/+Uyumj6Bf+PppHJHk
Eh9MdmYY05Rt1kCBNJkIv5S+MRhRuVqNn0tEQ/FApm5u6dcOqnbyJCTcj8sK0OwY
swvA9upxfXU66M8nHoHBIQ4rmtl2jeS81AT+8R8BP8xfLJ60aZQ4JOVDa7uUpvlD
KDziI45Rrq8LRB6s/sUgaUer2EUNMvssHJBqXoceKykUYbkByBB9naABADXmTXrB
kZ+FSVUnuBcGDA3gzmS0pGLXaxS6jjepnBd/aob6fWmnZMbGOmNcG1DF07qjt94k
6t9iVYZJr9qSoU7+aXLRoFDl8tjMosKARBNzPCyd69xmoBOSu4hLB1NY/Agm62Nc
o/9zWAm9sgi2FYWCa5YqMkhHA9iHCwYN7jDAAveZahBHq77RR9A61ncn69y2R05N
b7WWFP7FeBHOSlqgRxoOsBLkJtksHaNuHiSlF57fozJGsoBOmuC/ip+EofBqpZQn
JQ5d5zANsLFAz6SYB3kEAOWkp5sBzd93BGnfxXt6b5hpeKPJIXrzAWudOkIdCYBW
2eMK/3s12wf+Xtz5BQ2dyWwE/zmlyTgcDDbcktREOyRl/AUcPyDWYu8qtXvRGb2E
G9shTTidKj/gUU0ZMw+k1CUmXL9+iecFd3TuYU1I65gwanTusqeye4tl53yTASGK
+vtI/nS88g2oGrUmlxTGEwLtZHQjg1C2dl4eAp1A+iYwtuxRbKPHFqBBzhnBYVhO
abq0+1Z52Xz38BmZWUaxmNFf/slsgzCDqH8HozXoKoueV6TWvcKCo/8pVQuB24F+
3bleC76YOcHG0tdCwH82+bPUQ1xBrSJ6f4vrHauIvDhmfyp6AcxLqmpmiUnZl1rg
wxf79l0p8sWXAXjzfEKKFmCqumg4WASFCcsXgqAT3M+pZYPdoIxKz9X1DvewvVux
I07fhtu7yVb/UV/xTKQ6qC0pDASHqKRgPhDU2wrAqP3eZdW1l6Pr/JiLryXoI4Xg
5f0EvxuFaaOjh1yfeB10YqjPT6EcwG/Lgl+swHKdKRuDuCtyvtl7aA4paFVISRUs
VN9h113rGKLFz59661CYTv7gwLt78eBWFrvHl+zVjYYTAyoOh5S/WIWvvncGe6kn
ytyvLcJN7MUe29FuFv52zgHZ26fA0ywkdH9M06OXiDkjeMYxRl9x+kY4TMGWkwJQ
l53iQZgsW/SIFy7gkdYxELn8Ys2qzL4nCdWzVz1PKQTzQHSs4XTgjyVYd8Cag/z9
RJmngcDHNUlWE2XAwxtX+dun1k/0A5h/0+6C6u8aJwsnwyToUXrtlSNLIUfTEPYM
8Z93RaqaNwkCHpKlTcw6gnKpyGPgWr1WqEVCTzdpk3tqmYXMd9K11jfKrGQfl8T4
6FgjFOlztsAYgLvVx3jPSF8qhmVlWgpLon7kFTWfZbRUnXRu3L7311fOOl2PTUMw
HViFvtkr51LTkxu8x9SPUQaJSCURQsv2ajn4w/hYVQpjK/7i31sx54W8lcTsd380
s36bEWyYSZxaYg+GA3pAhZNTBznZyl8qBKjdWf5bf46Q/pmC2apNowlaDkm24HjE
cgwTvZlRX7Y3HqQs4aidYQsIVVK4pBdXHWjy9NTHuyfyjOySiQcWQ9xl4FLwmQ5Q
yY9mpZkQ31k/gbf9oykvkYCI01D34DqlnykUYwZle2oJvdltR5UsFTiI2RriO0kS
Am70JEzsTN8KgTWkkqJ9fhQNzXbeCc2Gq0U0ZpOWFKKhkZ+AsVh0+zMGbc8NN07j
ml7R96uYbGeLCb5S0ahtZkK7OmSyk2ZpeaonkpK8+YfgCPiHHbeNlPSSlCx3KnJy
VhbJSdECDY+0ckvQ/V36JRezhzdXxNZk7ka4Pi+/lLciUk0Bygrw4VaY7v8ifgvf
HG0uOZLFKVp9mPM1pc6jDhS1NAOyJXba3/X0tJwvNx+IxTgGIZSqb224piHsPwmU
mJkfKmSHtaGjiN80CsHPg/AdGDl/uXWZgsOeSTDWcsPf6ravQQ6pMiGg6yTWrhRc
kibYxYHhJUaeNSXnRfPOrRs+COOV9yCw7Dz800HnFd3XNI2sANZez6aW84yuCvok
XscBNeUDrgBav4Aq7ZHMQWvJxi4WExmPljaLq3c5EsiFGOKwuS1bG9Eb9oUznZkq
riLRCbqlYEAloBepJMTtkTw9rdVos2AiF/emiYgNXl4CLpcHFtGfJGNhAIp6Wxhu
TsB7Vb3+/R7hNQJopzjUQIq2MBUY7ObNh746fPgJl6q+nDd9rRy9LvZG66eyPhDe
sq7jXBLJHMNgUfhOMyzvTUI1tXNYTrHFRWT7pvTVhtnZ9bsobstGbR0v1THRuTiv
3O8VQAn/iWnx+834FjamBJ3ICwXPAohHxnp45U9V0/f4U0W/SouJkT8H0da6sf1T
kl+cxv6cLfvSxjKYk6/B6jc4HGQXo8A3wr2b9CznOcfI8LTY+myxHNQlcpgXaJ7V
SN4FndMytOdjXzZY97zeElELEhyxdGoQGE8C9ZWu1kZZcgQZFSPDsKV/tA3Fj4IW
//fDK2fs8ZGACIgiPjD8tLb/IKPeLa5uDA7aXgR3yJaISr+lN5dHb+Ch3n6nNnWC
S93N8Rm/uhRX/gJ5nP+Z4E77AiXqBRxfO/nxF7f47MJRQlKy6l86jWmQciC8ChDW
OMQr11M5KpvE+fSGteZY6Mgdg5fXQJe7wR/adK6oFNuXOH7ml+8Az40vYwEenRF7
B0Ggnp4/R5Ti+XXW0aHIM3pplW9Pe+55cYDnL0h9D8XyzDJd44ZghNtop8F2IU4Z
pJJEJWqX7Bb0tvO7T02EYMaMwcjN3LsX+gz/4JbfUgxDo7xqEx14YmNZl0Xb4tHw
ZdgCs3kRhFpP7m26hGxH9B3j9BlgH39/cv0bFAxMYEJt1mk9fjLIrh0qwB1ux3Mb
G6Wm5cdH2XI4zH3tN/66wyDe0GdeSMqcWSn4gr2MXbfnLG/cmcsz5sXiWsVxx7pU
WPyPqyzGeDLPRubAueEaAsdkSUVsDkg1SsuPIXToqCNYHAJXqbvhJof+eps5VEu1
EC5Q8neMz1dn3k6WwcpMgTflITaUoRwnAvbj8t4Zq1TQ4Pau/BCLPS2mXBkoI4IG
maCcqi7Sat8R7gekzQmIhlZs78YkJkmapto9XAJMJZaoNVc5owsrN2WfvzGnIHTm
IxwyGRVqHR+UZbW+LpkyFIc6BuaEdn/bXVYajvqk7niQrfbY0r+KPn1wc4DLW/m4
KHSzX10r+tFd8tKZFq7hMQduMhAM65sPDJ8Xnx8impzCbHoLoCjEMgD3hctAjd5P
XM3eAAS03lijzVHTt6hY+yG4laMpvTUTaHGN+Po6UsqZXa4lmHtkbubtjNPb9ADv
wvS5t+Q9s78zFmGZG3R7cWM5sKkiZc1IoFXx5/ztZGBFokJq8i+xSkXLIAerdfjF
zYaJXP2F3T57b2n/DO1GFNC8FFF8LtbNHbUf7iEWrJUSJ5hR6fNy64gYPCaLRop9
owHA3oc8xOIqo8UPwSai8nbPy+CMUmWPBm7rabn5nQ1exJ/RafLMvvsECZk/64Y2
X3kuxm5aloiyJU4Vs24nG2NGicYEL6gtSNAqt32jMAgBoaCldsVk2ACteeK1U9zC
QOSTIPU5eqp2lR57IgdZx14OhUBKezmYVvzIfIrBlCj1cdDLmi0QYa5IRUbB4K0n
Y+qUeXqTEBvOItOX3wJHrvjvlusXKT3wWW49tTDfTUHyKNY7Blc0d65vJ1lxCEni
4MLmYwHKIhVShFfFLspgNLz2lJYSfb+/cBwTtVD8BIOiuu1oFAqXosz5vYuexkBc
wWEJki+xrgTWbeZpD5FyrbrtxmpXEljuow7DcypGFV2jU9xoY3rWCrFB50p99Mvz
paoCOIyAytXdOoq1R7VCBW9+i5XoIoBZ5LkbdRQywUXDvcpRx9B6TmhAXxauLV3q
XGAK2a8KMeZIW8gA/Sx9P+wNTFyyFQ0FivlWP3UZZHctBKNwqe7gG7V3DWuVm+gS
TIxDvcV4zxZOeBPgaczYL3lnk1NlMrhOXjZkOsQvvosU5ezRJnneUGl31L3CVTGv
DAzLennnBla6SRXSnOtyAzPQ99nC+Nx7tDMa5hKRJB1iau5FwKPLYWbQe7rLW/nO
TccglTb/y3b4H37vDE7bLzBYCBG4oeJgGJnnQFQa/sAT8O9uWneuppmjRc1WPj33
T5qO2gOCk7N7LpQ2r8LRs+CZxpSC47eh+Fh86oEOilROzdaVYMTkSD0KMXPCzF6M
5qX0mr48t+0mHOQrl4OiCXrklWRAkuh++3T5p0q5M0vpJdi1g03Fs09+eJKfdKz7
YR4FnSEJUaDNtc/IeAgL92XtMDZCbU0Ctzqjp8d3CcGzfezAjV9ubHh77Zu31uZt
PSkEGZBpLBqiaRWPMneYGIX4c+E2J2fYw8XK2ts2FVB2W0Drn/e1TVabrT6CrGG4
ZU8uRZR2jQv9DO0oS0GAiIpuB5+mOE4w/BejaSG2OvBLeVDhFercyCjj7y+urlpc
a/Ca9INd/+tDNKlDdeslRWjPIpG2DiN6ys3F9Wiayj1Ovw/DjnSQe4JQklB7Kjqr
hd6sOlFDola38hWRS6yuhHsdaV5jmXKCI+EAJaLwRbx5DvuTIFU1uyKkJ0yPGZYW
RMkvRt3QQrl7GWRTBS7H/BKLO1gXbOQrnBvifOONciek83rmatahVFdXWZ5Jh15q
bYGRuoOC+KQot30LNixRAhlUwn1extq1XrQ74Z5oy6H/bEYLq0hmLQBCGvk7244y
eJTEtNklEPf/HCn+egZLoyC9GwhW6QLLhN0oYXFtAGyd6ZZPNhFC7ummEbbbVnvx
ZgIBV/G1Bjyfsa+ME2e/kXtKUspoQg6e6q9DcD/Rx6Na3RMiunKfm6bDzfbm/X5+
+5FddsVGv7ovjfSGgcLAdmgm/3AGoOjUGDHQddMmqrBBbAvkHRJo08Ztx4thDvQh
djiqkej1lDRUzXldkFHt0boE+UmtV054eaWfVAfENJfOTQMcY7D8oxNQhuGYfMZa
cAMlEJBVjDpSjgpC5mIqt1tv1M9KFlZXkI6lE/cTdVnUCWQhtZoZJ+26J1MHFfIA
5BkdH/tYgTY2cI6PwFD58ywTx/3KQm9y8j+oqXN764fHfORkJ+lcYIeJjy75gW4L
1o2g9rWFzEjOdCjyMPK1VSLE7CvaZ8uAFTnLfrifEwqorkJnDFn3jc/bL00Zuzth
yJxKU2M6w6RFaDTiAaBpgbidnTBxR5FOL70lKqNG1BsdalR5vZR5/3d33+YVwkMr
sWOeut29LZ9QQRrVQuQCPcfwGpaQjlhxnq9Ugq9DIATriYkla2zNsSEsnC6hwwCL
PLvYDBGTy1m8mQVClbSX49KZMXqno84zc+nMJUxzeXIfBfBspRkHe/1y6Ly7r3Ub
iQuUjR8gawxqX4pevrypP8F9ptEfuQ0NhETfULv5z1DYGKnp54hfOn83FyfK6B0g
onvNxWoprO2WRYhXBaM1Zzun8vRj+fXby6CIpYgSooWOiXMw9or72loVpCoVF9eh
M56KBJWb6af/vafGjiGPLTmJcxxxDVcdJwqPA0NNRo/vwDsPSKPAysq23CUV3kMm
m6qzePKwxlBapxUMID0D6ulchQjqIU1XMJtNvgzrdcE6YhcuEeTwSJFsehL4DatC
q7tXvIaSS/c5JoMWxxjeIx0aHokVuXdZrv0u/25lbwAH1Y+HO5dJkVky1IPGue8f
TNHBE8QOgV+3H7oZX6uguD2jQOvvv9lc6a4R8jusaj3yx4cpZmyajp2PLH9iDP83
5J093J2DOxa889XwyHn9AQgdXBv12KwF/RwpOzbglGZIuvHMffWc7Vl/aiem+TS4
9NnhxPp3SRkZvUsTwrpzTwcK6W+eeiR1TkDJiXta9CA64FmK6WMdo1RgcyHg6FbI
k8eRo4dbDdnS0I4DSSoIWUY4+M+UoXFcQ48WKUY008QFO+n/Ei7yGzIX9qsiB1uc
IjnRNeRiR78qS7ZUmDwHP5UOXDuSx4q9IDMO4IWtEvv7o5XF3i9PO2Ia0FGgpw9P
lsvET9stRhfrShrV6GoO+V8fTQmEC0ZYDx/95MW0ARWrj9lj+P2rviszYuG2mAWJ
J29XiVG/vsYvfixeCJRbZ3VNs5qroZnL+XZvdO8xFjnSl/2H10juMxee6HFoPXOJ
ZwwjKCxWwgW9GMGIztd/Ux6Ucnt4xRyrgMWdc6fMOdRUyoT9OTxQ76vy7GCLiwkF
cVfk1xt2ktezrWd3PRk0Y25J4SFgihs4ievPvUANb6gHRItlBkEV8/qmIqLZ3btN
//TqoG9wS/HRioOs/65Gu9TUVxvglKzJvJ2J71qyvc96U0GyqJIsS8v+kPIxf+L1
840nJobIvebGQyNbRM/5YNGEIErAJEfAMQ5ecH1rY6LwAeOS5VxqT2MZFqzPZ6Rr
xQq26DR934fiQ8rfGXbB8YPemykH5DQe5QNFUdxJi+5joKvbb1RuE5VpIeS380C6
3JOHoOpptKPHgTpvfPX5bq3ommL9g0v3nINCkiduU7r2g7miJZucWSlIz6MBnkuV
I16YGIYDcTCvTQwV4yPVRfnmecnwbmzg52UiHb4qNEwu7id7RxvVIFSbLbU/UZRD
+kNCTwN3f/VTxmvF4Y1Sdp7CS+Ndxc8Ofv7rbpjv8JGCFrsoFrJd9ugG0ho5j76A
SBgxc4ytGbCBhgfn8+DTKUKTxKCPKXbprJl1R+r8bSrTJwldnHBaLco09M/UdlcY
cyuguUdRJJyyo1fOp+fxHWm/0qAT5sDc++BXs2c//3GHDw5QNmFaS4FyprKq0jyF
L8o+VUhEv+V7yy1HaqU4MsFI7yDf2ERkrg8nGXC1sVHb5yIL1O6CF58IT/73l1C6
Q7ULw3Njwf14uNYobUWObMVnD/Ds2jnicuBxVBpdG6+Pkj2101lHhwyZIgUD1sGK
uWa8/iQEcapNusk3AmBPegtBI2W+vBy75dBHPYaCYr66Lu5BPiUWd49lyzu1wwdI
KBexCrcUBuRKWBOlXVZeC8HDVIuqu47dJA2aF0WGRqBZtla3eXHZHNmWxe5CzLTA
U3tWje7JBn+nOS/SP0O8qnAuDpAjx71xu3cMduOXWIQTHqzXrRlBUak27dF6MSlR
5Jkjet4Avnp9Ey31fxLLPDWGZEdog5aNyrprLCCiWNARif8Jvw3F0Bn+en7r3zCq
mNpRuN7cSYtWqQzrxKhioRLBzsOxfRAfEzl3zrESFyv8zcDs+DuV2pS+D6guPdrt
bdBzrefILNf+ZBwLqVXUxgKFFiOfCaaeybT+F/YIZNYZ/ur64raLpzWshJI30WKk
g50o0AfPNWsF61lFAFuLyCKVHqRE9hAQeaa2PFB2jHHbEctr6F/D8GaqNviU8Nwg
DWJB+x1qShoh6+6joJ0BLs0C2h+ma8rfAhkelVdZoPUVqigecg3FFotuYgDtPm6S
O1QQ5WM9FjwVrY2J1YXBC4+2xhufu8FomennO7Gt5OasaLZLFkY59KcdKBNDnpCC
9jxKDTh0kXVEDS4Gg5YaTN75x6kjfcLPSuHyELdWdAUOt/QivyhlT8R5gHyVE+25
N045RysXLjjXEaS+WwdHBNLWGVRKjuk7aGyqW0s5Ep2v5ObiNeoZ8w66mqjLmXcg
jG2ebpBGaOuMwrW3+LvYjRekhbe2fyQ8YyxlMG4g8R2tFiGbxYqSCiRdWKxRZEnR
tUiW1gF/UsheaP1aWevEP4A8DS9LzNFKAYfPTHrpeWlTSzMHX82t8nLSgGbfUMOT
CRDeZWJefnXiQqn06FnPAWOHbjW7vGswE0BgMNTipSOCadC3RPFDtj7/Sr/eCZut
+TQsTniM4ME8JOy+NdSjL9k/gC6FR42dYEsu3hIHuDlE/arDfXkhSOgpR479RQ6k
7h9I8PROk0MeUafQZaygm9nCmA8wRuYSGlPP93bkGRquHyGlMlwnRCUOCHqKzNcD
uBnf3nhMBoLsMsz57ZJKl5YJcpT5ukJtC6fijfaItReWiEQPR+7ThsM3bJ08M56q
OuiBSdNqIAExr4wdGj7CGRKnb8vOcPf8B+TyPhV0ilyeWjk5UhK5Ci/A6kCE7Qss
QWb7sbLMoa7oYOr22LrEimPwByKXuxcovq+ucMD9DzbvNSKDe0J59kIGOJXPGYBA
4vIDQQoXCrIv7mU6uwYIczaFnRQlXveIDG5teBMVtfMjg5QUqJ4oA67Q0jfH+vxc
KfLT8PE4frHihD4J6ru/CgFLFKLXpaEbnN0XFAqwzJu3zkXKE4Ml9oFlJu9e5U3z
q2TTZ5JlyDCk6uGuSUw2VWenSpzpNG05CaoW0hdnvb9CiJ2XkKPykLOb3l4EyWZy
MDEKpeqls2NYdwtDH7+9PAfUbELXi3buz3neOXivHeLOpJ3wQjxvAcbusbTf6jbv
oyQ4LZxpWjM6q/8NU+yD691uoR1/Au/NkjjLNY2TnzY+ssXgMyYcY6z04gJl2bVQ
KAaUcCPSXjG9TNV7h+5eH0qlH47a6aedLx5zBSJbT95XpCvHYvvfM6xBzmZZdEn+
qm7kcyYSRrH7NNMUFWWIjJBcTlCPvMykOX9Tcis2AVVXd0rEmTyNAtBkIGN/Hewh
4bIv1Balxy9g/P7Y80uZw7bhzpPBX71m0TVxpF9omarPEpuXQldulia4opzvb23x
UAaeBQ+Naec2BfSG/7S3UsImLMa/2HPDMHmpEwdibfum2nO1zk5fJtipLrBzR4xk
xI+rVIjNhKEPfon2kTIxQpbTZQs1a7iEczsabtdqItJ6HzKYFExa6YD/A87UfeGZ
sz8tGlkAgzILx5+KaDSCMSa22ILO8+D5izxjaRh6EoRZywZdiD0AGdyMCmMJLocb
1aubaaOyVwAuoi9r65fT4xaJ0bZ62mm5jHxRFPT0KNDQoySBzPSeuE4V20QWkUz9
+TeKM9Grl4lGVbxhuk4raNeuuNdAijtZX0eLn7dsavbJFFFf/vq5aA+IL70rFp1S
HTDWboz3lUnWLU4EZxdjJlI1J9yUS17reA5JX2b8ArDj0MqXwI0+ZOIMc3sg94cj
7LIRzafuUdTsThJsc0XpJXQqJtmrc3/MW4aRu9MiKq2u12BYzqKnp2ezdrxPE/2a
G8ajr8pHOl/QbLUlLaC+ubsaPXS8cnEynwcGsQ5OK/UNvdRQ8yDTr4prClvc/xFE
EtK6CXQgrWtmks+jh4qCAL6k8Zn5uOqkbjwEp1EZVAgCsycBfsdQRKobGWR6F2HV
W109tEvLgY3Iu0NdRqXDJmuKS6Yn7zB0N1yMi+Luy8mzoNSYJO1jxoxF8xZfGEsh
ilmhpU5cDfHmE4i7yy8XO7qlwKJwlaV+723olIZXZPe2eqntDi32j+RTYTgzZrnF
a3Zz6LmrrCDh4U9w/EF+cLr0kknZiRfbbirWppyieHahr2E7LIXCRMIs1QQ3tZkJ
8gjhGQOpaKegdB+kbCJQ5R6DkJ9aEp2f2FHIdKpQ5tmlyQIwERtZ86YnpbuOBwWP
IjIc6eov+3V6/8+7UtnzeJWTydi7dTwaepQX4dK4Ka103x8sbnYsL7tfqQcjXido
K0vUMbgh7gkU75JZRdhE0Iaw06pwOJ45rx6atPhfubfDaRraoy/xcgyoUT2LxHQ/
Cjqyy3JjcTlSXvqohhigNjO9D2hg1nA29lHGHixF7qzsCkbgSNeUF3ys4PwSyE0S
q9HAPW4zKnCi1jakEa+TqnpGTEorFP0w60WU1KhgRC8gLKNraSRxImoEOvNuVFON
Y0a9mqWOgDcEE1aWii+ReSgg+7FzkOU1ogXW8+yXPpPtjJv4R9lzIW9uVYN7+oBJ
zzxTM/zP1+oo48bkveGMtogXZffdBO9/oQUYdpeH1oNTFP4iWDLTYxeH3noiz6hr
e2K283reOrdQWXovJzYZ6BbcoDXfByiGIEdp1rKO4WQh8bhzXwlEgZAAubdq8kzj
Yp+mr7RLQeUgxJZ0uKbp/P5fzWFT31pZLnBKV6w0pkuPWLFiROtsYs00lxEWEWwn
kx81p31Fb0LhdsOmFpihhh2IT/7q3EpWxSVS9LmstW/2/Y6XxqsLxyUXXU+7pzSA
jTjGBWnIjTggqcMYaYr9aaQh1AbVk43Xma27cz0hAs81W9XOhe+pExSh2T/TAFIt
03LR++AD8MmspQtOvIPIoGTW4MA7oy3xE7m9l6mvW0M76frNMP/wDvHxkdh+o6gl
6qLgpoVOo0mhRavyVyU4+AT6AHWNb5VrGy+5qgCZEnu2lEn4ziuBXVOJh2OWbaba
ZhPexsSOPCfFB5TwGTDW9ssLqW/6TkP2MWTq6HaIkhaiSX6FTAjbZUF3NNhX+oW4
1Z3LBzZeE4ANF6DQB3fLkzw+Lb6zP56ymnfExaDhTwFTqhS0B79/U4e/UbWSHqfr
CODk2QhsYDgQm6GfSy5TqNH6DCMuaNN0SkjYDVP7wbiNrx4dRmAi7D7MDEU7g0ox
/aIU5x5NKDSRb9394pJABXnTTAurDJyNw4DLfUsrVKQX+ykk3kjF7WzaOQ7XsZx4
XdDknwLp1O6qQZfF+xHBIkjKU/DmK3gluNjLhX75rP3fgn0oh52rW1KWHaRsRTiv
1XbGm5CZQX/H+gSkRNb/dxdfC5xL4lGRlPX2SZUIpEGrexQuXWVZGNZlAEvNwn3O
BopUTcEfJpEMDp7uRgS3OHQhrON7eZMbJjm4h4uq9/zGj027QnsJ0lzTAGm2UUCg
iP+cMq92KxtSlc/eeiirOOPLtT/58hsMYwOUsmS9gRzX+uhjAp4hZ0LfqUl4/pvw
T+k7svktSPDTsGErv0F+Jx5zRZ2UehITDH1PdTy7XoHovndLWOAm2Vn+IUhP+SnZ
5/a3EBYf/uxK9G6mWS4rkrBvPc+yjJ7QMMDEl7kg0w5s6lUS0xWIE9dpbysxREFc
njRutkop3Xavu60HeqDeLU+b6Rl2Ctv7zaP1oaIfclwwvtWFoh97KBEvT7oLyHBv
N+zn57Y2w6GK900LF7nANaw67O76/hlXsxvFFNRWxa0ulTLyTgKD1QLw+xjVLwLc
pUNuB/mj78AksfTcTNn8Nk1K7h9jHd+PrMN0+Vnu2/AmmowfMnoK6Lf1C07wGVpz
1JspIIm+AEegRATXqh1RNGjjhgbCWrH2z4wOP0q5MboTTnTs5BNFjQXPdpQqOSSI
gLECc9ohYp2KdiOIIRQTw0TN3BX09S30xTgxqRm5pCmXhiE5dpDjNvLDcKBmiOpt
WMUm1bitIwqRuzuDQH+yIlcOPwnOUzRiWDwCJSoU1LPzbgyU0jAxLCn+2T2kP0Mr
zj/6VdLYov/INJU6jB5dyyzvYxNw2HiGS/L2Ktynce+NgSnVuQYtqvxBahzU2jlR
XHo1fETTWMOPj7w9sFa03kOb/K0VuSNE4geUt4VOSCRT+VcTaH+5CWIe3tSDhvIo
8J28jj3yTrzGpW04za+Twku1fxX14v+rQXFV9Ezyg87S7bEdfHEHB5FL4327YVzG
vgXtQp4tBqZIPBFbyoqRwQlZL3IgCiAmw4pmfTFFx0o/HGVJrUKGyoYZBXUYjwjG
Xz69lSbnALWK/Xw8+xi2EGFxX12skwEIX3EPCgoSJ0Q56a/7W23p8IT9uS4h3Kkk
EJM/gTWUnHq0gub8keKVLyp1osaUN8S3qM3k/D/4fNm/zciEEvA9Kg00bSmvrHrO
oh+EzmnGwzmJYYiSAyDLiq0ayORTJZ/Cf404za0cMVhsqihSv9jt+nJ/PP+ZjlkM
8PLzndDwaDRKX62QCBr4H4+lTmB9nKtVJII7/Z9jl++hL/MCBRWKJ+qF9LGi237W
1A2rNJUPsHk4OfBZ3E6QcSyhott3IPpXjVZ2mHO1zljgVYxWLKku3Y6Rp0kZPf2k
xhUIoMiDSfhBNMe1kZSOlQYyNn0pbQrKENh57CjG8q5MPgWOrEmAtRh7GwOliF4T
nb/qsPDS7dlkaLOwiaDzFu0Wp5LeN+6FFCruVARxtA6qYU6hnnGcrs5i5xp2h+A6
dZ/BRVlXIyV7m+YvsAUexafvTrvOXI3mHA/w5LPbY05OyGnozX7heA1GCpSjYsHy
uhdyIstKQjJ2OolGLYH2PBeIKktUDvU7ncUe+7Kjo6r1bAEkIOHGZ0THwxkPHKP3
guqnd9151wiaH3RuNY+6CeR94jlFYnI1+NUj38t/144NB1yCuhP71DlCufsybi3f
k9BpEdxPqnsRSP3WV+YrpPs1T3+RH4cmQVYpu8NpvHvBr06ixU2ImOJFovsdwmLi
grWcXziyrTRhW3LSnx2zo7thIBqC2zq9N8DtJohb3dgh3bBjTQqHI6f5Zy66SCKa
Df+WAH3okxR1wCN9WCSk07n5w/ivETKhJoTUlOBU9RUUr41kle9rRrluMjmPLaDW
icqs2+E9L1YZKG6FU8Ifcsq4ZomhthSummvVzHI7Zbw1nm4oHy9pptCvG9bYtmeG
LcsOoa3l4BIhNxAlRD5UqDsnNihGnGyU/oZSseLtdfZ+o5HNFHTYQfdFFmg2ApTB
O8U+9VXMsuj1DihA+vK5glsaHxrRbEf9aCvynxITeaapmKDSpyJXb+aCOOSUfTww
OHTq5MX3ERP0cbwiN95zjxlvF7xLATH+YNKUx/3MkWQBd8ibQJBUL2YwQBvSECYf
sVMVmGygY7aK/TZw07d9LIArro2lBvGeKaG8brED9j6a2BdPMK9tdORaqx7dmbws
FOciMLP1nFapJGZHo+67CewVL9VwyuYi0N74XDofpHqCJ/K2yNImgYpqilN5r0nn
BJ6QJoVQQ1W2409kKqAwie1yTPQAYut80oRuF92P4XUCc3WupAhvy+43/XKM122e
NTF0Z/Je6A5YFetHaNZ7N0AE+75fzcqLEh3/x+1i7lUnLurBAk5puhlCQSci3MN3
aTU3HWZS62ESvTMFRW81CvutM/a6JbMKFO7X76LjLEc15TjNBe89nANwp0D6sbx5
S1shr/1fcIQArDNQuwZp4uOoWI6kcrL5T9RllarzWbaTwrNdHuYKo6TqNzBzvC8l
CuQ/y9NgqMgU8iDQY51iTqoDSROl9mk8FJeLWbBw6nKHZUVpOjkSfdeQ8TBECxY8
EuRO6NVnNA+o9GQC1paEw7jmXmGieSLNN2L+1HTYt3M+3Pr3tCeYLASyG36eA+rx
EG7D6dCnqq0rCQpmKdVv4wUpOcP7ZLVL5cm8ZVCsgRhL7IhthAvkdNBeAq1C3vpL
kDjK/hPL5yPDK1Ld6I1api1eF+YvnvOu5stGwDbGEKLZ6a6NNa+yLeJ932hXSA1B
k76Wb8tAEoeFAwBSzHau4wu5KZXsMHprrXligjMyVi1Zel9dTUs0H+tG/AWcS8qG
vqI99NAjfrDWWiR6un0dnSEEbXXr9MGpxm3hWafy/XbCpyn37UBjOTXPBJoLi7Q4
98um1m0ryMHGWGsf+iU3AZo6tiAk2CGIdyn21INT1bQtuUcZlEJ4eG9mVFnW9kPm
Kj2/LgsAX9eFSXrsIbUpZdltnRSSfNvxkbTtgbYDx9f2u9fCXWn86ojFMxaezsmf
qoCAhYyH6oip7za0gr3hHSHLQl77owW9HVdYOuluJ+eguyXKY4uokiAkHyGEpP1K
EDTfUwqvBjB55zlW9GaxsOl13pvBZlSvQeCoE5UpKejy+8PRzoUEXYm1UYbqr9MW
ECIZCpB5MTkQLuCokF5t/QXv4+5sT+sGrKnbA9rdQbRwPM2lzmjoUefOhatvdeT6
o33/uZxKsiQyMDLMmYkIgK5zjxjKicuKlcp+jRjRhyUJHC3L+AdlF6AkW6oMYKbo
9A1L5eeV12LSOcy+vWJH1+fDvXsG2Mi75n76YG2gUsckEmWjvGOH2eJ9U1FGna0z
5Dvd744t8RVKchShITWFWOK0+fl7EN4ydbb6KTol+1XajUX2yEtCv01hNH2q7fMu
3akXZGH5RIaQWvAaNiCKAnBiagooTJ1Q1/tpAa1J+KQDP02qbaEV03A1jbkHYx/e
jPK4pQpQ6DJmxKUlPrPQOfIej3RXTpkqjNF5D/vONyhtUMbbOwCKeiRInQLpyRsu
2Qtu4OHQo5dHlTP3PvK0OpFyMCxjYWWBJ+dhe9OWUpAxz6wWndUzzWjhylsPmAU/
RKBeINlpsvrejK0Ou5IjZ7tXIUaUH8NfMiNn7I1O/zcOit3vXEiXj/g3y1Y2CZ6U
uGATPihpzg72p6qQmj4AGor4EGtzAzV/khIV0UuDN2/1NqfuF4EFTSwV2oBP9dEH
06DQYU7+POHYwYUY7Sa75pdiY9VJmri2Nvs8RfxIGQGlxl1EBKnIaotVdByvIVjf
yQLZflNTswJpxh4VQ/tNlZKmj/ncgDyzAw02LuN+tn4u0la8NV8uuJ/+F2PxATkk
l9GLPxoIhIv7HgQ/p+j41m150WcTptJfQBs3ipBQjiYTZgiQZp7StWrwiMB/yUhW
wjDxz4Y1ZBH6Wp0+ioIlGM10mdBG3QbcmfOJyVAr8fU8QHcjDe1+1xAgebw5JUH2
Akwvh6BSRU8Yaejfb8ah/+F1nvpVPHkA9EKJUY8IANEpBa7PaHCMAJ+qpJhqO3xt
/qzu0l3QScAJ3pM3g39Q3ZRwfYW3Xrleii7mjwuY885TZ0C928VTEpg8xjsOKXcj
uvqzSA9KaR8E3tAjVd6tOc2FCSlYW9ieRrDMP5sD7Rwg3QI9MsQ8Ma8svEI2FY9l
OEQ/tzt9pkZFTIIG3tSD83jsle7xBUylbAtGRuUQ8e4pXBOpQBMvJAUzz0QPTPdh
cuBzQLyc2b4IuZ6eMSfU47+sd67ZQLKAnRt02fNNH6EL5N0U/JhsvJGgK07XqfmV
JCojEZHgy1NkZv/EaTd4acTcwQxFmffq+8k+8eMd4tKWor30aAcghWdyn7ASoEoB
DPToGki9jI5Z/2yTGycingRGc2jnouLqVF4RExK19rcAWG5kJc5m+iI/D7/GncJn
UzfPHNYarV74ixzxnh3zDjo/17CWWy+DHRq5qNz1QJaXb4BRjiGGqDGkDG4wOuRi
eWPlxty483rwrcNokmZ5BD9dorxsYGkJgXHnCJxkq8v9C9NAu8CHZraZ5JS8aim8
eM6LRKPytlWZVX2OL2x7I673B392hLBCKUvcHcRo/hvsnuLMEVAnH7XeVy8QFJs3
S/oot75NE6QapHFkr3ng23bEsyzA7zMQFUAsjpfL+fLEsswTpgxhw58lo8kuXuVH
QQauSyYGEC0jbuweJZvbhtFsibDu41SdQNMyL0VX41L75h6vBs6inal/7FiXjNfc
UrkRXIU6JPkPzM41B2rd2/R61bO8Z0414ZtCxe+t25lhL8Is0eelR3qgPo/uBW6t
WADdER2lXcgULfKHgNhajP0qlCTok/L2eOUIZl/aZ7CVtGfmVII9tciGARHdhQq9
AaRDtO6pLS7eJin77CSocxkhISbPoid+DXRv2H113Jb/eUFKXHOJocddpVi8dfcX
xLoAz26y4Qz3Bi+BMb0pazU5RFw71pE9eQp3wXSzfCh70OLzDmWKHxRkPSv99oSv
iUHBdeyEq+4BQk3gH9vcYAxq6XeCbsYINAzMOk/3+aHlPozBqrEQHSMCUpgGpwme
S+MKgBXkakf2c3YnwsxUJob083Cp4228leHy5jFeeO5WlfLlu1xmsxDMBp/Xb422
bkMrKKmDFzgz5lCpan7h1sN2a7P5ldzntygQnK9yevYZQOz5H7bTU9qco8ei6E0I
zh/v4VcTWijfFRzl6pcnqTi4F+2qZjTLCx4FThAoGBb56aFh1v5KxXF2WDz+ZyrO
45zbHyR671ugtvCN9EF1MvnUXg3INwKpDX9gx1KdYQiEhMrdBk/piRFQxo+HYyqD
2/7DW0hSovgj2fcH0n6xxc2rgyy/5AOkpouPUTdbYm1tOJCWlkJ1TIBy/KdHy20K
MY+9IdQ6Rn//wV1Utmb973bxZlTq6SyzSuNtq0URjK0DKml2Ozs1pAKzqTXFFe/7
wzJrtluzuO8LLpyOqIwADJcqUGsIY2vBEnL53EZBKxt7csVaEgaGrRtZbYZroNj3
hAiNyXsbZPNa/bXfumcTB5eDTNZ4WHcaGqiu60eUz7FAFT9+EoaxRNscrxBb1yNO
zm8luTUN5qW+nV9jNwmNpG1DbAmiZh6RL/8QgFer2Zu+9QKO/p50W9w5mpwzOiDY
KkEPXr2Oh5jZcSCse5WqqzskGPRIyPQz7DltNkgPHq8cXCqGkaTPQzinGiMkqW5+
EjzHX7s4/qYRVFbu3y0ZmV4vlThxLpjHL3tWQfzNhZTT92RdQjgigLyAlv+jxPs1
UOUhfbfBm6qD0y1a8GbhtNm3ie6G/bZybWwh92trP5Diba6Onpi++xYdt6cCfnPG
g4vFhPc6Y/B+Z89HhuNd9eKcMEguwEjdNeHG+3EImMcLyU+g45FByQtAtdX1d+Q3
xN+TPWQJ+9RpEsf8XSnBcT+klGAuSXkLp+DZVG9ZFfp9nyGPFLPD9+i8aj+mVVZS
uOVh+42tKonCCIg9aECyj3bA7EV0yTJXTeQ2mDprorhkqGOukBSyBQ1yhLITQflA
/r0SExag2F0PJd/5pawkhsuEnV9G1MyOM0O9u4QQBHrUNVZEpTIT4tRvEdN9B82S
aqza9ZvDxxLhDEjpCX4aSf+kqNACw9HvIn/Z5mhnd9GAhzZmcmhnV3aPIJJcma2X
B9iad5fQ10370cLzlKX7sfxQBidYeCj2H8qOu225xTNOt022RY32JBtWIT0HUUgh
X/q8ElU0c+wSLnrI4qKNFnGEQoY843w6ML5nhwPveuyvUD3N5DMj4oJ6ACAhnAnv
hXBaI5xMv+Mhe2bcf04VwcGoO8ikA3DZTis68h/oepZ6yvADytVx0pPRFUqadCPU
A4woXeIhRwMT9R1YgtDmHkVUgFSJniwLIS1nizRDAekJ1yKPPm+HzrSKPa3W1X5X
Wtkey4chfoaj9Q12RYgr8KnPp5+gnMa47XXZKpJVUABZ/RJl5shm6/n2yxujPzuF
YeMZiTGOSSyQoTR5M9WHOf4f8GG9GflQo+eDS0ffL+uxBdupKWTaLzW07CmdgR6f
OCNrBM56iqCRUnWC0FRLeq2/rsk6sv8TKm0Tkwg/tvm5gcF+sxdxZXbOhhwnPNHp
qU8awYtM8qgvxGe3eUQxwUp8HYwbStBEy2bsRAsployUXgPdHGC+0aQ8NPG62EWG
gx7LPI0luKgV8PyF8aA5ldSoZ+hO4Hwxb44NnMUPBJcYTU316rkrl676lg7s8AjD
swWalSNEalpsGPUBDzJpbg7EEBDYTEzJtrRQJ++988emsFgbvByvH+hC10vzrUeB
LgWIyqeyEknkJCE3YfQ4/bG/ZFr0Ehp33aPx+W+rpec4VRUkT027LK7S6+YalkbP
lbADKES1a23lEveMbDZkuQtoVbyNPo+xxKAIapOHm5UbzPZlx8QZZhbxKU5XHjOD
2QEuZgFZBupHQ/MiGaJA+bzowNcKL0qeVTnlPkbv4u0nvW3X9SOwkD2xPUMb6FwV
8SC0VJ/tZUp0dxvWp1g5TvU2ubtFFQLXNp3vRfamLMOK1kM57MF6OYWPxdHUCMTU
NQRx7+ufNRXR4MRUpgTtYlHBYdzyGpNP0wUws/SbOH524DZTPzJEShTlXV7evpDi
lLQeYp8miHYGj3UaQOul8CtlcU01aMOdVf2xdWnQ/WamCCB0a1pAoYgmKO6yqBFH
k7L9oDhVhBqblqeR3iIPlUq4q/t1kD8xqgvk5qlBDmyAcXX8oqJPfeJOgHpPuzTZ
wClDnq5fxD+0RNukS31GdkV+6g15NU9+awHRxqKEylD142HW83M8Sem+dfDm1DAv
3rVoHrjCkBinMRdwOJJP0JZtKb8JFTZ388fBnaA/SaH9/lJbRaAlz3AA9doDBvJO
+r4mFZX08kKN2nruwV7mFjOVPKrlOkkVA69BBBNbKxGe8uCHETMm99U5xNo/9Wb5
cirlXxdtn+6OYRtKJTQi8jkTB83h3In38REDCM+R5ZTr9bCx1Y/4tAFd4qCxOghp
QsMaCdzD/cIpwoVSKIcnME1arhGMq5WRHnuwbVj4GwjloH6cKElyxrOxK6zslEVg
DXSYJVIZS4k2YOHO0aM847BXhHn3zviZ27uMEomBRCbi9izpXYjIdNJqkBhjQHcy
s9SjckN4PUbYsetrDPJbu6aFWW6G5CquQdZlKuzNlX5y1VzihgGtA5U2scsygMt/
McuWVUnbwKh5+SgisPoLN/uM0lQhhFSc5G0uMLBQOx7/sUbcClB14uWty6kJx7Zv
kps24JAtrWw9MpOLLzdz/sGnYiJcxzaDp+MjO+2N4TbyjUk5fatNxfXXFgftMbzS
Zhv3zAIaqkcogS7bgfi9BVLFfJKhJaw2WFpMWt9gHbeJXcrVTtVahizQs4D0jWHo
HOVX+PGQJna5t4Gbq4r5YMR0/LtHScTdca9wAltM4n3F98eopZ12ImONmNJE4fJ/
Hv5zNxUpF03R4WKQt9rvdWrRrhH4VgUr2sXS2CQ4psjBiGIanHQ9TKwM5FjodsLA
oof2vw1TmP71L81foxUapCD943/2dNOR6XbM36gcaAevmc9QbGho5vKOWC/3WWQA
NZ/PFaJd2wbQktGMBR1kRJAsk4+Rdeyrup8ZIXcc5jnPGn8OruSvyh5Xgdo3hVTf
97ckvcHwbOhe1x8hrtBBngBzXaMuLnoZpBI7kgls5oRz2EIZW7tdYmhy+ZnXaPDe
mTChzBoAjIOJkp42f2U6ASzE9uqoc50esu2K7eniE6Ei/YogYBC9IPOj9WMpEHFN
Y1VqGMWYecJO7FJRUWZ99Hwz2PBMVbbMn978kgAlGDnXHrEpES3SsXJ6eaKemBAE
K3TAyXp7GQJ1+wI8OLrlUHuP6yFu42ckauSXYkz1FuQ1Ugi8etzxxcWQ9ARKFOIx
1gQIgG4IIXP0Vf5TeUPjJC9TWPxjnMm/mlJHg33TjStKRZK7fwcIyCR7edppLtB+
HVdD45ugrkPIHU8Dnb7wNoy7Emc1hOP+TLglqSRcpPRwQdV81ggCfwNRyxTEmcEH
qQ02QVv18TMyQDSsix9utfKPvcaSzG6RRiCReg/9yRWJOCXob0JbtgBPrRi1reMy
odeG/+v89/h1EVvOR34pKr5UMVN2VlNEh6JMxx9r+eLJAdxESLYbeDOB83g7Hr1A
V9SNqjhnX7V/vrhI3mCfYWcr0sLe59ZGBOba3dCLZpg+WA4Gltpxtn5RdwIOgTJx
FyABKUSYytI//PKzUVQikw6qpcxnDPAvgXJR2j0741upmK47DFjR9EjyMWerxN/7
3R8faa7GWZ87Qe9Jy5hqhgmYds4elXEsjdprT1/m1GmJYS9Q91ZSxp76iz/8d3k9
Kw2NsDtxPb9ExIRIRRBcmN4uwLIG4myKHm24fbnpUasc3P/QDAadnxlO8bRXwB6e
ZOMar9NWCizkWexH5sjAeMo8ZTn0MyuC5eZbiwv7U+bRG3Qk4bE0YazLm1wXa2CO
B5VT7gIc0KKZyw2nmDx9138A7sSD0mxfbCVW0QxwnCZ/5zJchg10ybXaZEJiiUMM
WOTvvNrdckewub7UT2klfP0oV5ulay7XZTR7dlrScfn9siGesx/4yjbR6QvRaMuN
ZutJQuElSVgCqmbFgwJh5sm08McO/JGalnj8fVe/MSX/jSpzIzXHExOuwwbASArL
D4aQM4RJJwhBRqPt7ygaYbiZ//crG5P+6TMCVBSkYWPmmwkBAwlWR2FEk66iGMIE
EbOWepvLD6WhInYfdzIo6GFFTq/sxf84+V3vd5fH9u2VFj9HZSrAG5beZ0BeC9Y3
HXZwyO214VbXVKpWea3vbqKl6FO/uGMRD9tS3khHr1wiaEnYva6xGLpVSrkQtYGi
CPn+nQ+50S1alxSXLgi1Ow3J4vZReTO4HfXE7yh7boY/nY67+eQfsM3gilkbzD2t
Xra25/5/lhqsizhHN3tbuoBX0n0EilhmLaCE0zfWwn2sgfvvjg672f5rKAjVMYrx
ZrH/79ZOAecM+MrCHIC3weewQxV8zOHZ7qogEMvknAcd/MGm8jQfUW0HPUKMUUkI
81/JLnPYyA1CmWmUsFtsHzdzhSNMwbPy3CoiBISR1vGVXttZWYpAufWskqjSgG4k
W3TjqP2bFU11+lSFdxS9NIKyS2St65/s/j8n/jbbuaEUNbkn5KoP9lKeCYT3k8bQ
gSzEACTHpL5XUqOK8zcNGFeU8WsOxf6UhdXxtNLFDsRkRi7xiALGl8Gewwm0WTXs
gY34SDyNWIqVfoPy+j0x1Fvhabr1UgmucpVKMvE6d38REHkSs0jAKxan0slJJobF
QFawCKUpCBFZxEaJqXpZVzrA4ZVh7HfBKm6ZOjUu/Rvt/lwEIfViipkq8HmGTnnp
uB394nqOBHo681/cv/4+gAdGgZCTUA3fEg7rrlyM78xZ5gP2++katfSGGXRHVQE5
Jq/H7pKxpA5yEbijqQiC47fR90QQH3UqL62tHicrFaXbHuBTWNybLaibPTdN++69
fN4j752BNw0VWboFXF+AiGTbJyDEL9Qxu2H4sFlogrPcDEkp7Ah5JUbFM11SPJh9
MuTyJur2ukeAvNiTQaYGKdOSSP/avDto6ThsfQToNCm/LLiHgonr7botNesNFFC2
e4NZywNl6Ag6tbvxKuzs2/wEXZIGdRJjxL9V6OzELui5ogKnQGpGSe0Ea1CPhW60
PN/0zbVEWfE45C/ejccovl1vvvqvd1Hgef/sdWpMKrQ0N4NX2R1quypTDZGbJqPB
65fejbfAyhWCPffSFf3+XaDB0tR5LLA99UtEpqhuuTv9FPpN2i3E9lZlvyC6C0pN
ai+2tQF18F60ovn7bK2KoN6WBrykxzwM8eHYnqC47rqYdVM/5Iq4hO7OryvOWCmr
Dp8NZzDybE4axxPhtHv2cUFv10L2M0BGZu3fKZ5utmH22XM9OeScXDhZdgRStv/N
p+1WhucLO7jV1aa9k0MjgdusGps2xh4ThNEe9CAuIxPa3vSUbPR2jkB6TmDyBNzX
UCjWSuQ8G+xBTj+rW/H2XpgCPmg2YQb/zmf+NgECpweJPE4P6W6t3g1boL6UYBcX
WXGT58JxqTdv45WRhL0xcW2wzxR+MkGjmQTc7OA+O++NlMmmqvX0dHa58zICf+3E
zDeGTEcRdEjbvI6r+EVTuzkIfcRoKgDmw2OcJhZ0JC8frnIJH85u48LCDFbuP0Ob
OBHVlCPcZCYhWt0GquV6l/Rd6RBMA+TnIxHFB9jjHXJ/J93W6QnZ1tQDp9x7qiKV
dzH6i5rtlcubUOD7nPuNCuqrKq6C1uPD61bqHaWADRA4SbMiC28WlEl8YTe7iLGd
x0anQX71lhs/o32YWuR6ZC2G4aK58Q/mwEdwjYSwJGau9aQc5gGK7FKQik8PfAL+
GTXPuiiq1QSRm8Pni7rUC7iw2nHL7IoALRMxutvDxmjXpoB7FKQmQPd/uxnnVZSQ
ARYvP/UqH2+cNmERwiI3ohFfSUbGXGSI9g1u/zxXyUAuXN/BGKbUdu6RiuA7aZIf
zQF+0ZSeMfWnK7cGmPTofURnukOqdjOFocHruVM9qUzqqZQdytAlNJJSvbaYu8Zs
ndctzjlFev9HLXy7iFT03NfkHv1/Z5cwyZl/LuGFLp8ctMm12YXzYKtec5vQ27Wr
fqJRRMouX4Zlh794Xs6ihyXhd/HK8HxZ+10wSVxZTN6w35yS7LZD59cCl4wT1Y00
bQJqktjDSYUYhDf4F9nWM/F9efwei9pD8G03Y5iWEJuYUaZ5uHKHhh2uIahScNFM
6MqkaHQ95unT+nJk0bTKXAh6RN7TlpDsV0CQVQHTTQN8ILX1aTv5VfTq+iZtF/MY
IiI0DWsBoM/ehUXbdRKE89qYO8xQdYHZZKzzWZlrvH7Bs7FxiByMSr9eCB/Bd4jL
qd4vRqhBdYPZ1NtSwmmcN+7WHVJDmneKJC2MRyn4o++Ie0UfDaEGjxc1W2JwlyhL
ZHbWxdlmo8lWA9gmKC38AXVkSd8USvN0siwcIZWJV9y1OiMoPoRRl8ZcWK1Qzg2x
PkixMXH/740e8jto+A6mPMUkuyPcnXCV+P33lmLlB18iUheQcUz7hQ2HoeunxFZv
070Y8uqJs7ZHYzVvNOzecRXmSxPqNP4vhf41EOOtzE/G8h69DP6FHfFUKUzo+fRJ
+V2hJ+cn+bsX4qGQV7fHztOii+lVMmhC4reV0SrtwroynYC1a5BuQvdukN1g0WUq
F0/lbhSZhzrm+CwD7gNIqmLaDVhEUGgUHkUUUp0XlXtpJR3Of0cRPRgHr4AqodzX
xwHDYCtnOW0Eh+ludu9hi+VDzylN/FfO0xs2DneMLq8tQ2CsK8yX+dW0dRsHJxyB
rLxz8o4s75PtyJ0wOkGaCHlQk8xhY5fAet5l++6r7X24v2AjXNtyqc374M12FaDf
n0FpH/cpRNkagdnhROBLe02E/9sfAxb4asyEnxvi3OVegt0cOziHB2mkymF//Ujk
dV9MekYSpBMYzn8usfjDGTgSGONh7W4e1F7XI5EDTXca9u3JxRR+/tFmeoOfNWKG
Y4e8PEQYyF5Xw7gxIGYYM0Nay7ThihoCN0SOYP5L5ILJ+cGIAK6hN8WLdxmr2xMs
wKi5shmzG5U46Dll6Jl10A9Rv7jTbIwp5SoikeVxvwCxtBB1Fx2cx3eb/ZONEdew
yIiaEVzfxLPN69UGWbdfmKYHC+1KfLhIsbAoIqmX786uaQHsxr8M71UKMVFsCC15
1MUUtAHTfBr6lrmrFgUKj2bCS4cXENdOw+m5tDJSTZDw7qPSq/hikfDlIOOr8yqB
NwFYG2pJ/h4dNVhrinUDWbmwhmeGdiw0Q3LG358pv+Z8sKCNEG99t80HQ+SNJy9O
JrovkcaJ6m0v9cGd+2GTiAoj8C2MpP/AkPodU9z7s86uXdR4D31sXE6XmhSIE5xd
0T1RBxklLJilmG7WJgVVA5ql6TDLi7/ArQyRN8qMXOluXQTQK5zQlIi85oBm08ud
0NNBMtKn7I7PYQq3x00w4Wv75GRGCoQpJM3DS5rj+f4jswI9zfadNzrUaACnOwzw
i2fJj4Nhowh9cZmCjgwYbqXif3X/PymwGiZOafzTrwBn8cUIAvhiBKNvbPXSArdX
oKGYfB+Al/iDputCMdK9AM22JKSQG/XvXhFuiAQ8GJMmB/V/HlbPGrZE4nAE/wOp
WQbybWsJEJwov/B+lheM1+vvpEeb/t+X1NedhFGqWK2UnNT4hfFrRhh6W9hTtd7W
kngYh6HbCeV9BSG0/KnrHb+r1ZdDeFn3r5uhu5oiz5NWaY6d0dl3BUZt7lZvadDq
1h8oLA7YbPD8S2hEq83naUXzH6mjm6fIC1iJGG2JtRqPpDVKHfPpriEj1Gf5XLaT
HNx3/BUtNK93tfc+rOkD559w9zPd7/VtBAwZVTrTC8F4phg70yKQq2WKIVD+e0SC
P5L2qDVebuk2klfwzHub5aNIgS+pf+eli/EfAaWjDpu0M0GskaPYeiyWYhkgWzPS
WR8Wna9iAEnkznHbTarJJ5Sni3tAs+um7PXQ8N4SjxyNJwlljzj9JW3Cva2a0e0B
QH2M+0+qOEWquQ/GkjVQIRudPptqwhmNrxsCKTSQ7SqwJvoi/Uo58qtr8PPJlw5y
QuibPVb1MIDFrqQZfkgFNVo2ZKgDOLHV/xJfoNCi107xZCLVw0XODdZi1wlQdJ1e
C6n8YTr+6xuPrMdsiwI5893EdWZ1Ah39AJSCopZELOEJ/PgrcwDaDSRSunSVzrzc
OHEnTJ5aMO2tdPP3rH0hzEFgaXjQ+MEDxfzJaOahx7lmj/bqyzcqT+RZ3rWnj1Yx
/9zxrjPVA8HFHIzmoWKsqg5KKeKMYs9Fvi4MfzALxFFPv3b8pF9TPhCyEX4yafjQ
sqlpz5pikkCfy9RIbdlfncnix5XgabQMVx3QWutMyu1mkSnjJ5bGSzniYjukphxN
IDLowCgRAHLvAezc56uFEaw8m9rdtrBERuNhPf7kdNSotjBsPSuM6npN7yS09nuR
YV1MX5q22WMSR6nVC10k4IV08nxZ5csrM209NaPMTih+odKtfjJbCQN6Kx6SOKpd
FnLnHzRChrhEQH3ifo6k5X//cKtsABEUo/XQ5tfV9Lw8tOcPtgMMjFBHqANKQNkW
XqomNXKpHLcuXyFZ/nGWMQRKzxlNMlSQ0H62VFMEgue1IhK2Whg28Uh3TYANmUTn
wGygOXRbWdYUpFz9+UMnTzXFHh+xHQaDekdHZ5ee6CkB85DFEIQzeq+IBSfa7AVh
ZMPUdP4Y5JSfZJHgjacD0GtDK5H0nKOxFBKUkxfnD/L1toKC2QUyvB0+pHtPsjVB
Qt0cXNMVykxK+2/htquZRp4XUlOcvW0dHe7UjpkJpekVxLVsJ2ypAoxs2EsQYfR1
8DJZfK1Xb0fgh2JaDvgHWapB2G95mVsWUu84L/bzRvHA1/1Xoy0IjloEY8aC8Yi3
3KzLNdOpC1jSDCVQtldi3u/hmBGMJD1ge8woKV8v6zkGG5q6nuCSLe6z68dRbnWS
z81HP6iwbhbzLzl1KS+zxRxfW1EyIK/anHH0IIM5onNweRJ457etJd5nRhT8CLx8
snvIJ5d/txD+Nj2ew8rbosOM0o18eTmLlok8yc2AooHKtAck48D18+2L+CttXEAk
VqlZv78JVjLi7FwPe9xAgKr1QCCLw1sFoAQiYZ4tvyaQTznRCrn4Hr3Nts+P7Rm9
szamOEfPqQwea09BqN5OEi5VYxjXgjxZo9tbrAhQVMUAej+nsTck/jz/oXKkx5vr
nYuMhFfm9t2W10AgHMt8pbplD0XtFT0Z6egY3ISur/6rkucMifMAZp95Ag1JyCpz
gKhBjBd/NLYlbaBVHd8KowVzvr9/EYfAxr65ZfyCfEWqAXqzlCAX7xT2s7OxVlg2
IGrTcY2gdJw/DU3kqBP8Ln9MmTW2TmLDKgGoR+9pJstkYeX92TUzXj4bQDTBhN+p
8Xx08LhHG/BSXhboBeB+xKHQyVrv3uerPCC7IIs6QlBi9VxFPzjJd0s8S4JFRRtJ
H+4UZyArqyUObgxSS2YuTNmjjDceBgUQjMnovDYBamGX/gde6Y3o2MN7ozjVrQSz
04wKi8f8lSJ1nLrXLWP5HnFvMv+46u8XQ1KnGU3KqQCLKfwc8j/R8iU3VC4DPsVl
8ZNdXb/REp7icoCJf+dCnqUNPrG3FbGkuZu2my3uK+VZuAXp4EyL+wcCj/pku7op
TsgfUCZvtiy9+/026rFydR+qR2x3mIAXlNtSTFTaIdrt8LsqFKA5+TC0IQxqYDhD
igITYOQzLg3oN36kb/WiCBU7JJbvytW94NKy2cLbBK/08HE0cxuy3QqnU4WmZJT2
iWU/Q9F1Boe61usKpFkQ7IFywKQpybKss/bUgM7iJe4CpqctP5e/obpJQAoKQ3nS
yaDf+73TcW2zpVP9RX1kgQHekok3Fuwc2dYlhdpn0uH4JsQ5LRjFLV40JZzPZooo
WXXtZj2Q2CIU/rbne/MW0UTm18R2mkFw8fSqk+i/EXWc+zyYiO2ePIzv3ik178M9
xnGOcywSOah/ihW3VgJl0aj0+WHw3DhH14LU24hgoP1dh4XxU5boMIne7D2HER/E
tGGwjsz5zLG0NksZVwVCVbePmwo1Rhs5OA1X0TUdYZsti9efE9snXh2lV2QzzOka
CNCDTcMP627vb1W7B5GJRvFzJeQyh/2CTqueZrpumEgjCiVXscCBFnx6jqv3HfbX
Pfd24lr0nLSQayUIHJ5OTb/v2GtRr8FKVey/5t9SH4FMnDyFesY8Y8nJ3Mh2Unol
rdaAZMu4ksj7bb4vwWckmGesM+3YH1Z9RlSQhGFi9+qRdeJ0d9p/ojtlhGvXyetZ
2Vt98r8UqlUJADU7t74TZwEbEc3Wqhg0PTo/LcKqcOHis9MUtOPpOjX9CUIktDOt
taBoar5wznKHY/ibd44fyWjgvGnZinJXSousPCF04dScENqk4Of6C17Jn4wsAhxX
xaGYQZ/wNOtHmNUTZZIpeni0dxnC2OoQMsS8c0cZeSbwAfuSyYs7lmjltjfAYzC/
tO6m+JNV3sm9V3PgyzNIr625y9XPDvR41DSyIdsquw/QpoICDwDuf4RUpd9pzaLY
s8PBChgX9PVxtkfbnPkNyd4NH4xvmXjcnxUNUh3NnOWs9q80TPOviwEYCvAgqt+e
qdpU/2KlhzPqu5lJLiqVK5tE4Xkp5FLl/Qhjy8ithqOTjt2BlfyO/6RWUUUSearT
XhrIvgjyNT5/ZGXPz4cZwOMeEGze2FW+/DB/vwyGPjfr/liSky1/crezdxsoFMen
5AOvJZovhgoFo34Hyeo7d1IXLYI5DI61UKtLa2qKZ1TGoSzTXGW8VcVNoTWcF/kz
zKml5U/t1XeeOfC2pXZ2+7zfjy5urSz4fRZG9zPAi/+1ihC019pad7c0Bk3TcUgG
W6ULBog8/xLe6lMlFyuIwJbKQYgmK7Msmuk63Gb3za1iTWOWhkPlMwJKn+/MGHpq
1MYICSgA6NZjhQ13z8jRN/o7L9oRH3RChP9rxugxkdeH9BuUbWTejt/uGxwWEN70
AZG2gOgTKqS+xxoouA2rjCg9cZF/nh3nHcQSAyzi/P9W8U8Fw+0ycoraGH0f42RA
JJguqRCMXfaHJCLGNRwkZyKGpCa2zvd/lxvYhvdBlfR4j2cBqNBAV5Hivws8eXax
S+rKy9IRKMFq7oU4y0uStwKMon/g8ypBUMPxHVH02zqFyRSMC5hdKja2JP0264Hp
u8jdI9R1nG9oBO80thfgqN7E5eXwL3GSSLTWdNgjRnqMmxs8WBKpzLUN1pXIgBLa
ddC8mhEbWr4r7BvwwmxFxVsLfUZZF81xNKWFCB+HMsOMHiDvpdEvCUPE31BBCIg5
k1CgGW1tndoIqob3sEBySHXr+QuQ9SjdITMwc8cK1LHRXGF+EbnOzic9RMZtHsQI
+9cjbb+stpr5qDq/YDxksNojOjy3B+1u8MmU0xkT7Sk/iIg7l1K4jh6OJJo7dOJ8
7jNyasGJdsZ9gx0isW0Brk0K1BYR2V9TWyWV6lYMaoibC+y2QesZjZZu70SRA4VN
6j5ZEwioK/O4hnkm/QGoNeq56z1j+KsntRgr1J8lDeDZAhCxYB/3HiSK84l5B47L
QgfRDemK1QSDqsOdWbdW1Fn1XRkSFX2ittMbcKWhpgJmp0YvpQndGyfkK7Iy/SFL
DdetZGzQwqSbL7BLSn26QPcUmS92rVOly7MMXRvpVeIrvGnENvbbnpx7Lp3dvFCZ
flQgmfmEKjZVLoGP6+dB1+J2kSydLUciT5XSJgY0j+aWnawyR8cLTO9z8nZhIzQG
4pba+85ous2pLja/MC/P18OpAGhNVssRxbAdScU7jFZWd4iNxNa+9MF/u+pe9wq7
lqE/8AX3XlFRna1orDTM18qdjy3zRFzIJISXuJu0oc0exw7nE3ot5b43YTQ883+S
7IMzj6dug8q8UcObNtyMgSQ4Av3fwYTBkYxNqApoRcOQmUNDnVBWRR5yoquI+KSI
ACxKPj/qYPSvjZCtX9aiTJmJTOMgzNQkiKP0pvbm1LexkNqBlMb7Sez2aBYBDwu+
34L/e8lreSc8+Vim4hzr/fzvJA12R7kUyPqeZPLT8JniXljsSqw6ZnN983WzTG1b
XzH1uUXyUCJBhuBYuRm8VBahl3GENzafIOj3uRfSAeLXdMVvk4lTL5UdU1W+BwyE
iMdyEAM+JrDEkGVm5S44GEhMiMpdfzSVo0d9N0OnwdjGvUgh8oHAoch3rbylvcTl
v0QhzYvu0sGrtrdw3LFdy/dGXeSDvk8IiQWsKI5UOykeBsQohvHmpRoRQT0BUrj1
l63wR7yUZ6XDDSh9CT2I7IiATWOcrNHvckkTc1F8rBZ/1sI0CtJ+VwG6HQelNW6H
mt6j2sSHGXuPg+GHK3r5SQ+Fm/x1l5amZY6a14d1RSkN4kVyY9VaQzVT73yCpOd5
7mYXEELnxmgDSbFOUW9VfmBCzK8u4+tO9XYcE7kpx9tjhjBnOqUByEegsnontS/m
AUNNT4yUlv5p4yZGcyQDspqaAZd3mBSMuAJUWby4AcdppmaiLo52mf6ZcPdBn2tb
tdA43gfNf286JcSGqTDjV6KyLCVgnDtRI7TtaG1uoTs3Vf2msvcbq+14EKftTJHn
/wMyL+D/iZz0ifzFucfThhbdKtWb2UHPejR4cSkZ2kZQsS+vv7Bqq6xJI1/PxACM
bHLsbn9wdbfos0A1Fi9iyVf0P+12EojdtMgPi+Q17LSME9uKSVN9Fq+Ts19U++1w
Ws5eCagdADCZeNiN9E3ASABPBqtdpZwqxEEYMv3XPI82ckmX4ttRoPCfYAX4QlOr
fC0KQ2cHCVGs62cWyfJFV2HUosIlUEAWRxScy6rnvC0j+ujmcgCHQ+0Q06M6Og1V
4GFgbrbsZGS19s7BWsphHbVqG6oZL+JIhdborNSJ9emyAph9XP4bBivpKV6ZXg/G
KebdNZuR3YaVjbE9UNMDytmNQkVX+tO+8YXXj3nVXhG2l4ZF0QGgqaeFbKMjMTpo
ojJ6QchQAy/9NTmfo2t4veh/JPMSQDN6Thf4YQ9pqJ9+CET46cUQfxdJyu5xoUP/
Xe6IqfHN0tCoCZKmu+eAZMoPQY7D+uZz4yWdQEbmJIHfPEGjoZaspBiWk0My6QC0
BHqajLvFh6UAW44L3STtiLgoDEgO0mHNWg8PI7UfTci13U5U1HbIXxabOUKvJjEc
FLp00Fci/RrY4DxIDuf5LN950At3B7ePXdehRs+iIiC1I9IMGLZh8uj+ShVxPOQO
8++GBT2zBpcKfyuGWzzQXRRfcbsvFoXaeaougQKabUlVzfxXS/ZcyF7kV7AY/nZw
n24r4S2VkNjFMdYUZIuG/vjo/OVxpkXruHbrXTQGPghslGI3cqVtFZ1Zv04/aMqE
9c6KHcJIUE58vbW5k7UOLsvEQVSod2w+osNawvUzAhKQq1XZtRuKH58qvxwGUkQH
giNEpyeJNvv+I1BVvK/uwiymv98218LyDQ1WAygSqdeNYT3H6ooZnbfvObPF0TaD
vXTs3i1mrLs21eoCkUpQ7PBJ22nX4eKGLsTSXfkZNREwRTj3338C7AYldIFhR5Yw
fGzdO1lLERwp7XTLmv8oidqUwhk9JyxRlShrNe4hADBoq6NgZyK8yfrAflIHrq7k
YDQvp9w0B7AxXYie3EbWakcWOSld5MpAkL35yE5N9lGPf0fArml3QcqyYBwudJRL
aQtaylHy78QtWp3342gM+GECzj7cEtXGhO1YT6t/5LXxMKzfEdntwTdNFuYQZmrZ
lcBOs+t1G7xaP7OhdNUxS1SG/FWoRwDD6SKwzLBReYvClXGuwFfaYplp5oD4EVHN
ZfveZryKqZtMqNjdUNK3KBG8ahznkUz9HOD8gLwZy55U9Sw46efX/tEZr/PtvTbO
94fA0hGT9WBG6ZSOwYYQLJbpseOq6BR78HI4kePTaCkkh13IsEAGRfTglmAuf98A
HmqJLTDfToDQRjln5OeUv3SmDyxFja/3EeG7EkayyEdD+s5nQUr9ZywIrom9zwuM
btuV+zYdznmgbzZO/bisjIOZIHS01kpaHUHeCpxyXYXnIqhQ98FIZsIS8Oa8zSog
acbyvccJVDT+7X7arVuRJrnf7EtqIL97ip39r+hylmLg3/UrLLv8oPUE/ov0oOEZ
vEYwHcuWkQwUDjBrFFVVYV1y7fpIWa2Gi8CFu3DVAyKhlWH2Mr/clWJe+JWPqS3U
Ja8D9bgb/I5BtJzjVqs+IiVw6maLWOjsKQR82FcOCwVNWAU5GMVu2TqZeNdvq++H
ajsFrWAUHfrg4safr692vEdzgRa/kpEqo9OY8KFPYMRCGZZIWLLU6fEUvmd7nUE3
TBY9h/ZokNX0BxSyXC3DRkz4ChqhKCTFt3MzjJ4xVKjXDban34zU9XGil75uWf0S
DlBzRpC6nvIi0bDGdpEvlADq9l+qjaSGdIliaZDKGuC8UKQAGOsxORSG9tCoKyOu
ap242GnCvcR72pndhb3sX8qf/lZsbEkRYfxSGIejgonJiQWmgQDBiLBhzxyw8B5j
ow+6qfGeGhdRIZCq2xevcP8pv2JtnqH0bwoH/AbB5dzI4mj6BX90KxFGBn1BUc3/
flAiGI9KQmgY7B8daplVUEWt73Aemi9LN25PZbtXrQR8kBswYpllkYMaz7q3apJ5
r8Dm0nBATzyPdMxtMfjhiGEtZG0SQmxW6rwdXxM51XuRypkFZeXxZwxwNO8FN3cr
fDDAZAyQS8zROzRqpfnMKrdz+Cp9/cHoNDmWhOO44bwuZXlACHMvoQdaGBDUyq1Q
ylRxeBav0IzECOtquHFTuSGOf5rpOUaX96ZUOiYSoZdjde2MC39pCacqtscnH01v
0lPvRDo+5csdsMWk355UzKjT9y6RTiIlmxRvwAIXFyLYfZXdLpAh5PcxoSoBnh1O
+DvP5w5jPo82qgbD//T/BIY/LRgv+LFIm27girBCRecCNvxb4jRujTqTquvKVT+O
JRGo9YPQKa/EzKgRTx1taqh4uq6f7AInyp0AZ3k9rPxZgUCg0WyPqGu3D2Bwt0y3
ZQ9S84p9Fb2JMIHDt7ghjjySPnG2gNW5oCNZFR/U2tcs+c+vZ4JjKuQL+dcWySvk
mJlOxgbDJ8N++hWnpEK0CZ4NLGnZ+nboP67tAVS3mWf6zYi/GowCQRhhCpbnNbQl
Z4BrjxTEylcMW50hRF+Gs6ibBo/RxvclgzSSoM6GWuPm2in2h5etPUR4CuZmQUT2
xQXMspaQ0outQj2INFRFK22WU6QsKf16+uRw0tqbwtI8xDQdLfTQl2Q1+BQ4k5ml
mVrkf7ABybOmbHnFMFZG03kx+/SV5mCTmQ3BR8sZ3AsB0PYia71ysjaet+qq9eu8
tOEDVlB33vIMMapxdLWQR2rO0lRRG1ZIk3lBy03PA6Q8OI2L8yhH1CF3+ylIPx6w
Z79LGAr/y5aiQmN7G9AfN7is+O5xsk1Jr5M8p0otrQjbuu54uH5UvNxa5E1965sq
64iw92Cxlejt0ec9yL0ySxCixCL+ptoqqBHsobu6ORFgqOQfHBp87tcvECzt1MaM
0dEEsNtUapYGFzhG6c2BE6RzH2zyfk1KYBak5ZyFx96AK1G+jykngpa9Spj5aH3D
ZhMcCF4sJUXmTVls929IdF8OkLyQB24zqBdpqUv2XRK5U4S5ZNp4PmXG+MjWS5Gj
FYGEY2x4v/d/bY8qFpBQVypemVd68SeEnJwtnzAsv/fXn0Rxv176KJ+tAjCiJoIi
2efu5Kxyrnr8iLS6prWmjzHPmAAkpZqTTtZthZPq2f8Lwjx6efHf/ihZf88Ceugy
ssd/76dLifYUHaVYIJta6KegzVAhlXD+ra6bELcuJ/whivfye5iaVp+mJTbQG9M7
d+223o+8nfYtoltxIwZfIpY1MB+fpoP/PBXqRMNQrc/JgFdv7yYN5VKMcuzsvLbi
000ODnqJmnUqO0Bq/QlB7T55a74Brs7yUStf/Rp8jS9u+QbO/l6npKW6VbffRBYM
6EUSotZLdjsQeI/0sUvz3gwnUFnEG+hBKkMl6gGfgX7zpISTrhmdPNMPvKjtH8lV
LDthcA/YRgb8hu6FJra7FQumQht6y7XPJlPCUoyKEaC/wQt1J3a/i+42m/qZmR9w
jmM0uRenbOlo+Mt1ZEyS3v2le6lzbuzAls2bsI3TE8nxy2WsO06E373xZFr1dMNd
3RCm7aOuCptUoaSrfZ2tT2AcgGQckjG1CmT+7lwxtlyfyeLdc0s4BkO1i1THTqmW
BCSPfGIIHK3hH0la/L8jwQIli0/FckOu9JvYaSVhVXKXDrjQBanHIJH6JlGUxvGu
11DfUpSqrjMXhbaNcFLxkT06mt5Zqd+2tJXNt4+NcWcVN5v9PkNySzfyhA2c7QVv
y8knL78VdWWe6C0f8AezoEshTua/u4mohm+z3e5j5Qntkx97nP7B1+TzKDcPlpOW
Vb3oeIvveNga9oxm+a+n1eiqpVCknmrh5sgLwv69Zi9m16k496MHr41VI9vwzaiN
yH9Qxvvc7brORKl/z4stxajdoE+rO1NuxcvPOriRk55Nnpwv1S4VHas+9IZsUwEH
6eR4GPzayZ3slrTd6wdQ3J+H8sEQM9UhoFZSycDLTGJCZK4dljSHvE4mTV8Xqy3E
ecK6fPxzE8+/JdWFylPRqbLxal8jvchzv24SYUnof1WYuTOeL0tsivndGXmKkKmN
M64upDwRzDWqVkk1r+Fw30+Y3/RcbqhRhWKc7j3yr386Lh+Gf3rONYQ1ob2nI986
tA9boxpOUwM4FE6ZBozAxsccA4uj1ona0v6CfuuLbfw3h8sgAUTD8ToTrkIl5sVG
aTelTatAbcs2Wf3QUcRoLiV0BGAzwzlXb6xDj2QGnxnvsJWblOaw8DCSSeKNUBNg
3IA7MJ98QmEBqJnmMbCoCaUdWIS1XREF+DNye8zUfpGoseXV0q+ThtceMZsHlrBj
uggYZl8X88yGo2l2qr1XyC+GeEjG58mSyLFaKUi6leTjTPO4OYesKqmyikupYmSn
vDtG7+y/lggj41iNMN1gC4EB0PJeanRZU6fAQ6uuAjuHKAdJzkdttBo5cZqqDznh
aFI8i0dsKSIvQiV6LnmXP01X6SYqTAm7yzWb9LUl3Q0y4KZnJgNR/2UWbx5ZCZ4Y
C2TZiY+UkldWqxFDgsBmd18ZDic4utVeg1f7XIt2w7qikulDGinw+OBGeDkdT5hS
Dfwi6CmIny67iqe/rgRhL56fYchr1OpbIVP2ajByP52DpcJ9R+dCmBzgIWpMdl9m
4iJDPY6TdvGwV7DQ3nkwHLOgkjcjaGew8y/GQ7XKgLtwMvjuqhP/evZEqXkARn6n
Dmaa8yNHL9AfVkiP10v2Pi6TEbY+ZposwQO+5Q1b/GelIQRME3uJiJLiWq2upg36
9UNRJeUor9Q88OcyjDC0CxxcDw6g9FEaZ8IKDsulsQsdNPNgFurETNjNu/saV2PV
RFWMapCLSJAAK/8nRTJIhk88OGUr2kfbh9Un4freuTJrPUwVZTcZ9Ip1KUyBz/BA
Wd4xFav07CPIhqfdW7Tt92Su2RggBWn2QHA/qsUd5PXWnCcHSzzXcJ+d2B0LNciI
aMLKOalbaueFaJ5qS37MkjwM16TmuZhjg3i0j7MGxblDpB27EjoeORELEheQTHXt
ZOIFVTV2VdwOh/ULauQOTAC4DlOWYilaIS2Zpzri3PCrmU/8qA5vxoxb1Dv7cWbi
FyCanqz5/5JwdPhT0tEN45QjYX7zQ8Vs/rUQ60z26CIMzBaG85sVgYGY4/xYeuG6
UmY5vUwIKMJN+bwK2qf2u3Pxtt19GYvwF6/gtdfHMP5l1U3Nq3cp/lUf+p3ZW5si
qE7a70A4FdHkqV68ReM7NNLv88YcyGUHluQScrvrW6W5D3tKjT41hSnHoxpNc5d3
dRZ9blb5pNIAK9+AWtpbKCjdQYWpLVJUZyMe6WaiDIkbDK5LDElyjOoxA87hIni5
9SpWYSi5VMtHfYTzc+SyurCwdeYco2wv1HOlWWyRKdfm9T6oF0dRR+ZCRve5OUGU
mSIwSjtneAhCOHLY7P+9+X8EDpYo6c3DgKarv6jhH7u3dXJWoaLOZKFJkZz/vAt1
s33crzWudZs20tboueFbmiwkDxrUnbr3ULgQMfFsy5gMROYc+2rE2k4tRtb/nbt0
y+q3U3vTvTkHU5zg7EJi5Ia2pLqGjjUwVZkD7NmblDo7PSK11x7vH6uVdTnjIoiV
uUxAy6y4V5XJWZrQrXoD/LMmUbP74Qg42e4Yn6hZBSJWDyjfc4fy2FUK/QMUeSW+
Qdx6C3kb7RXmz75By7Eo02pKhD8Gv3S3U3xkBGqpqla2nNfWVPGBkMm6qdNUZsPc
Q6GYXKE5oZg4wqJzZVHNewkACUz5D04kPgybDiK8vM1eKb5GxIClvrmqGqZJjE+E
NJTeTfC6pZ0OI0lLF1rAwadNPSMnKnn5dJp8eUjP+w4Fk3VvyOPG2FUD5K8mIjNd
EsAOm43dWp3xVeFwGReE0Rw3gMt3yc7UdVPX5CRCgTSOQdyfk4Tioe9RfuVcLrnp
LS7J5Bvuji3F6uqSK45oBFm5eEvfIKj4nmOKj9Go2TCltzl0WyFKZ/WOROn4BQzG
Yw4EYIwLUP+MUteeZ2OOJhOFWRj9PgkY2VRq2hCM82Qj5fxUCdRVQEz/RpiMtS36
zFB8+HKYKhP805KAaBWicjE8ybxEZY9dKe0z9o641C9jCblRTF9D516N7VqZWjF3
34ikaTRaaojQZUE/9uqFM81Y7UoCfFFab9f6NKbXJsqVqe0Rgg8AZS4HVVxRGE/6
sFHtY1sKmtFlw+fyfAMeNzMpULhADZkTfOshAQcEix/cs/rsnGZ8Hc82uGdlPhcc
oLZ484Q20Cc0H19dVsMqOo0G1UPDkgQraELyZRMcjjP6ifncPdOgEEgJGSX7M6ny
LE+t+9X4yKvLzDXaIsvpoM19SnVJPOWR1ZLIQpzz0+CLT8UBbBCetXaxvTJQddSJ
yJ2NEnHuREUj16EMe3UGWjd88PtKDFWLNf+oUC1Z7FpFqBUETMHnm4JzVMuJ4zqj
nBjpBjU0LKbQfdzHxFnlJMTmZKepqIAcJRYJrc7Gbvjqb9VfxzjqgEeKDucs2ASe
F1eO9IsAbbeWGxOKh9ImW+EuBPnpyns+cdiWGoz/WXVvry5yPKcm/yQkWl0eVdWv
zsK1atVl5JkgFMSNiFxxFYATFNZ9BOBqighA6X+a7rDDfOSGbU9CKY83KgPciuH1
9IFNYg0+rgfSKItGrk10tC5iV0/PNCdDlD0c5ldLWuSAx/hAHEDXoOnFkGzEs1Iq
icIF/M5A1kTHUzs4wCingWH+xyNpn9+G/u+gar96QtNHb3TNL5tbIAjmu+h5e5hp
HLpekkp3qn8ezYGX/g+RNwkGJhR6umrvfVask6MxQ7QWONddWFJ2va2i1+9TEPAD
wP/rtAhrM2ULNdQNmgmZLoecht7uACM/l+fyi0gpYXvjH5BADoKnYZVrsVQnCwDG
2jjOsXkctjpJd+V0a7nnW7RqvSjwhL3ofd2rigzBubGS7BfDEQz3tjS5sUz0mxQD
EErdl/a/6yEQV8kf/J6zeyYcmj9bIg1Ds/Hf4zM5jigbTNWnO3Hqz3+CnCV+w54o
wIJP2VjxT8Jk43RJer4QDBQtCse2KCaTcm4J4CDqyGu+O8cHwW9BG10vdCzkWQNy
SljUlo35Hf5NVcC5PI1H+3MKauYYFmQlYObzpSbS78Pov7t/Z374+AiI3VuqWISa
TmW2Qr4SisuWM717UcP/kaCKOpu8b+kEj3rvdvGngWo7hwZaa4wXrMi0hj2h3cSx
YwarbMWAv0gZxq8wDywuHzCIP5f8LH6iQ4ewyI2JSSg/lNaAH5LP5EmcXQkD/wnr
HG/dqG5WZ1swIaN+6qmshnNVP6KCFqa4DRpdyTmSBAXF4oDvzIGaXXlth2alHuHj
FMyM+PpeI5xXtY4dzF4zMMouGcdWCubfpd5yDDeI9BjMz5iJdBBn6ebQ1EZfNfAZ
jYekWtIFkoJXVnE6yLQomDa+NZ9xk/RiwVAXZ8LAUdpam4BOEvPvJn70jR0hweyj
Fp5NvCDc4Yho8TgJ/GHAZjqZj7mLHVg2GYqO/UsAQDNOKTB3RRHzx/llWT294tGx
psZ3NmLc2SgKVEZJR8CcHOpUqe9Uq3FSLtN9uC5rwUs/zUsY7cmPT0kxKu6Q3cJI
V8oN5J1E7trXVn09pez41OtTSwFR5iw/fGVaxAgs/zdhS0LSIWRzk9zenoC9fb4q
MK2xWdao2Q+KizhKnL5/ETbcMjno4szt14jWTnq5vIDZnXwSIu8ptNJQX8ad3WWy
m36b7srgv/0vsZf5uA5PXNmYFm41Ezp0U5oagRKYUisl4qf09UKS0v5c7+HNXorX
zYCYc7vn8OzYwKPCGsnjFN2jaxUuapUNNH4D1Es5QuBwN/SuA0rN0z/WI8M6k71o
raJEOWxVY0RvjHaFAzpfyuStFCJpGCrms08eMpLxNBRejlPOp4qBdJ8RamPnVSqz
y8FF73iQblovRAm31OFnnoyD5GT6tKT3+/aME6tgFTQYbuIA7ph/kj92nWx+eX2K
53QinnAF8cQ8CfE9AvDatMolt2Smd6uVsNokbMg+0Yx+qfhLkMcGdUXTqvyMWvoY
z2vQhip0SXRIqkMNfiZ0Ag5i4jglfxd0Gx9XgoS44SBfhj6aUAkR9c8DO4FPGESi
asxXMJSsiGImXArqCt4lZhxbOLSyB50nRam0OAowrW+1M9uGdLionCBx7B2Xhdou
TvkWHFPi4rU0dQFSHBM9oD5g12UG6cIYoupYP8np26fNrjqkK+1/8TQv8qNELb68
7U1+/Z75yTq4Q1Wp/paVkw6E+wIcuNOWf5pHeP1gDqyePfV896bYAtg4mApHXdKm
2nLFoey7AzyjmiywiTP+okeHRNZopxhi5NPHPS1VOnpLMa+CkOAqvYZUjni2ghb0
EQe4rlq2wJC7VwlLY7R1KpRUoYZu69dNR+5M8mFsQ7Z4cLzEHpa9gnsUcf0JfRN/
9anU35KuoQHya66o8+TdLpf+hVrJXR2cMhT3BwhR8+C5PxJk3oN/D4NltyU2R0K5
1SBg5TbEJlfW7p90/ugAhP59aOcYMIW9butUrhS5TSa1Oz/NLTcfvR266nzx1sOs
MI2g31Iba4Rj3Q2nkMeoP7bRV4GRjSu+qwksO/ObRxKa/2LmS7hrg2ICrXTKR+zE
17iVd6Cc4uYiwoAWt1VqEdFW9rlF5HuUhxLRa4lKKMrIM721zbDT8ThI8sW72B8b
82XeYA93lTV6WyeYVtEWB2H28Idf7LEC+iq6nzNQYNBwfiRRg014FHa/fp/DHBba
gth/XmJxt2SXKI85phQ+p/7yU29h6qBGoaSmRUTUl9NQmdFPP4saI7VYD/4m2nlZ
V5qsUTEM84H6xb/YCVvhyQ0GDixAF3ccub4DUVsn8Jv4ot3LpyJgCmLw0aavNjGF
+3Y3IdVkmHhCCYQTSRxi4nWPTw3JzFtimN2XQkBgtvle2xJWyKL/ka7034Hl4wlY
qiS2xq4mUGcnkb/v/CZXK7PkFl98MMNnXtqZftPH3ph2840PLArjlJ2j1blCuvjX
ZuHZJb8sMdnuegim7ChCBvEbdniEZevR3GbKcDJIpDz9xhjoDjF4Uzp8+mX0k2Nw
8MMKliAHYybFqUcgmD2se8UKSP0+rq7TAf0fhtpUBxnki8nG2ZEnEDSumrHE+PCH
KbF4VBnKTJPIssPxyzK0t5W3PkAdyyVVDpN5uoEHemw9qIXc8X6Gwzfe1D3xTb/X
WWRQ6YsxG4BdpldOEqRQGRwmQWopcLlxjQsQLjz2CG8HB5QKMzJq0+6tqEIbG0/r
kWVV9Am1r7c52Ds7zAc1IeNSjWMCV/B+V8+z50OYt46dA4iq2AJtEcMQzQiY1uhL
xBinwfNafmyLXsQ227nE+3cWF8hEEZv782UCoz6W0ZFreAw6GhTuPuQdkppjrzHQ
M9YPBaCKncAL5CULKLQE4825CF2XRg01aXjBfGWfcgHKH9MpYS1iKqzbQ45OSlkp
YjpEnMsQ+/h2b6b4ubKZ3kaA6shf/h/3IVaNMPKnspPNGw5sXM44Tfi/Q6KX53/H
IXAvI+VXjcLh4q3k7VN//XSEcFbmuSjvLFYpQ91RPLWzSFur9Nb1OEATZAUX4jSk
KU33j4ipl5wj5vTuyyov74ainLsjEBNkk+BeQlKofLfbdU/F5DHwGzii86Zfik91
aTvmkK+QflvLfCCvKk02hPrYZeYEEasm0u1tbo0LLwWDBsLlg9TPzLm+5OS/lQPF
mua5sB7qAZ76elxHadzHZ8nOWC1KGI6B9cL0hFuzExMZiA+rRhbVc+B5x84WfLn5
cuQ4VWvIz9dyEeZIGWaX5aJ9efTKIvrGPc/iORB8Vxj2ufCGr9uk811i0FeILREF
B8F/agjCeZEU8FZJEjTj5TcviivO8ZZpC5/FXH1rn2yq6g+SVqMfW9/0nDRy9QyB
GkTPdabLpbuCcbCwuO9fioCcGKeTFu9nYkJN1v714VnVypC/eM91/6wgPxzO9vsQ
/i7mvuKbHSwLieWO73QrVSXWrsrt6Pl7sUA5AaDm7cwkoIDfXs1czND7HejY66nj
F9SU3rWjZTaccqdZbS0zUCtEfAxKentfOnub/MKZ7RDI+U547MGGlHK3IHI8RN1V
Y0+UM38/XOuNve6KUkRYZR/Mt98pSLrMc55x7+5K5661gtninbuq49BEcqs/mwg/
tyQk5x/z1ikeggV+8gbbfdnU7cCGuZhWFFCoI5ZjvyP4z0t6mEVuFL6Qpb/N8Asu
9hjydYvF+fwnObSHT1IOyPjT4pKIrwznNOWvMKfGryUMmH2+D4lA/ZvJ/LYI3MIO
AQpmhnd7CdoOiHpKdVLOUVonnGVWbI7es12FO+dFlv4JUsaKlKW4PCPQTyleyK9O
N4VCaHcbaNBoSSkJgbX540vXs0umTs2VKKg6nREccyLh8TINoDfizROL++JH1rGP
6q2Yzkc69suK6zpTGwBkmyfXFA4YoWiSoXTZ35FqTjlZMKZRpphA9Fl2zSoSMAt7
yXpWOzUPL8wH2Q0m8rpRGraIPpi/coZXDQ7KZyupI9Es8+xLbPqvvFhcf0/1ITIS
E7Zgs1r5+jzOp4qK43UpBu8MSuEeAFZKxxjlLrKMont6RwswawHXNKnIcamDRDMq
yPvLYWLEx2SltI7PyUeeYwXbZZVT0C/vxTDQS4iujgHzohYncBKCn1mFRZZxQLFx
JrJgtWPz5ixsuf99L+/tLE7SpuqB4+n2aei2qKvUe1yTBbj/qgrcH54LM9SfojDp
Y+J5J2W2xSZ2Louq+OLQ0qUD6QxoUyejj9rS3xKXSOmETo2i9nm59jaSdEpf7AHN
po/Kr2QsmAFzaIhzRdFKqGHkvQ8Ihir62h/UbSL10cBnl96JNRfnu3DNZ+79RdvW
UZM0U2eFNNRRGuheKLvcbPQGeQynNCHjiFWA/Bvz7XQ8xMa/l5oz7AHfXaDXW5Fu
xkIz55yP5WFyoBkp0Gn4cdf4LCeP6a7lhv5Tji5wwZTtSHMInMrRq82ie2QntwIE
79NolublSKOVEPwSDbmvgayeej20JifOkzKa83zONUVJhr6f3eOeJDEXR0a5ndnL
4aZrdSAPr+a3OXClNxl9zFxqHikyq1Je22/Ony2bwp3XucsA7PNF9U9aMH6dLXod
T8CzeM5Au3W/99aSVf1FNyp+eprhot1WBcVGy++ca6GsEmiCoSCA1ED1UvvDbkpG
YJ+4HJlV7bUA+qF72waFZStb+VewBtMEQu4BSG0vQX00xzXk6fI/xTFahYxHGpsF
mh5DlCaXsiNFyNdKyxcpizk5mC7lMCu00QctYrlv0K0WIzqWzKmyNigpcxurdZu/
vgToB7ssfaGF+cDyZGVBMvFjMZq3Dr9Jw4oMex2x7cb1d3w7C3mJownaMwc9PsNz
wPxbs8jZF12BHchZEFBhs208/q6T93rMUQi4KgKgeQbe3ZgepDh4FN+GDXr8iTrC
o/PdfgWtHT+8Lta4t8pW4u1wzBn66NvnhfwXQ7D2/osLhZlfh1l8zs1p2eeOkaos
/J9v5Ixqka0Mn8avvs/5D/q/gscWvQUtovW/IM53isiBHWwXOrQjef2sSEI2oh6/
UetPq6X8j4ooNrG6gWu3Z18ZLqyhlKNFVfwmy0LMKc7c7mQUayfMkzTwsp+OlE/G
/ReV6nquM1v1Rr7MZ7QvXIgNHRhucNUcBr3MDrJVoMA/E8V7BgVNQzLpBrgNc9CI
p+peKydZuUhGIbZCtzTlUvCx/m5+/GFvgpNo5Aw8lTNm7wEGPlu3oTHByr07kP4b
DX+Nq1Olff2bYzr+zv5RKqifAmRDRVdpSB6ZNT1Nw7UNB7oPXyOP2a5l+I3RfhWK
gx+gD2omBofOZL433vLPS+m8EvOdm8VqYgUTfPGCxBMkVCN0/UdK7DiXe46Ab0I5
1AmyTaPagVoOdHSv/F2N7p2SKkF8TZJHcI+W82ZlaJLRT8pAIZnMgawTdfOMGNPq
4ePc99KZtyzDDi58ocpElSfwm3zpO0Pdmuu70qi6a34UW2hAvvTEdz1UPplenU6F
kuPN2y13SP9/0GDm1tSfe9BbGYJDVYHMRAqfkJ0TlUGYbxwzpGe6NMQwOryOGOKF
sGrPMVqc2J3PMZxedHI8L8ldccyZWm/Oy8egeGeE8bhcrY4qB3f8UrvYSrsUDAgV
9dQbevaCzxqjE7aBKliW3ACCsGqRI+ZL6jywE2EZNl3xDx47UU79QqxKyCzl1g3H
WPRAcUvxHkLF+ymDTvPvEpk5k984MVMANAXA4cBVtym40ey64uu6uMAPLAwSgc4H
Rd6I8x5fiOomT4KveFy/XQ2NHAe+XhjsjGm3olEiLFWzwp2I0F1wmwz+NQxluq+Z
mn4QI7OyVZtdMPDVnFCxZu//2/IPT6GBuFdFjSTZnmbHEKR+4JP5rybPXKc/6TNZ
ndSpHkF/fj5kDoLl86o01zpVcGaYCPwITXoLrKeB+w6v8zc7TNdiVBO59cuHdb2M
TLtLCz/iw5m7WkSTCc0wDjR3d07wl8hbM74fRpay3jhgmmq3URKKxRfASxXZGNrb
XinCi56jBtKI9paeS+XQu8u4tjvmmy59iLyWY6tRr68lO8wSASFNX7lrxHFo7xX7
vaBRWBmECKLHnrButRbjJuxxIFSme9MLlm/flZJwynwRMS0z6H/46wXKHbxOZH7X
ugjESExQMOxXF1AI+9JXTcBrTsz6ah8SIDpiv7FJFZPYZtlwx/jXX7BNh9oPZYYz
NtmRg6L0ucZ6TT9JapQdkLMQV8Gmc3n6+CrU8Qljz552QuKnpo6wzGCvWgwNuNge
A2uKif6wdT301CwdAgU6wvcdyUZUpTrhwmSrO1iUNOMeNui7vDjI/6x1PmYpYNtn
70E+nrFD9oGmvczx8fsIp83EFxh1xAKNbsS7YZzNK3lXFaoot8p5krAseGX//ui9
rY24D0BSL2mPEyc70bhrMsovNQ2yTZgitcg6I8mUarJD3GXD1GcnOE/B/LAlETQD
f0wrf+7E/MQPpRlDXB0OltjdD3mZ6C1bIy1+f+rwd1i/RXhpmkkHLIVs9lzRK92I
mGxV0gdBFps3ZuQBSzgCcUszAPJkVWULu8oetdthMXKRDSDbClDVIOeWjifKi/bu
uTvwd3YrcfmfcWDRPTwSuNn5Qjv2h0Tc4hpe4qs8bw1E+Cno3IrEw8Cd7x+09d++
5z766oPhkw71l+p2Z3HRvMkMu2rRd3y6K/jvgoGYrML4eOouXFqlcq3FTXyKiPd7
fUHSQPZAPRP9YNTzwy1grF1xInx7KORbZheGL9GsMjCbkgv733TRDeltni5sY7RB
nUDBGP5ng3hL7qy/0fiGWzR/183h90x/cGQ82iFhESAPVnGImllx+/iKjywq+9V8
5OO65kdFZ3BjSiiL/3e1kjR1p4q2bJ/sWxnzrzh2Mr0tChkAlp3xHM6KCNAZuhYx
0U8Srd5Yv/pEiHZoR2L9zDlcuvAyXclBPr59+S8QN2dMzZEqFSsT49jr/z+Gb8fI
Ch38GXMrWyY2zE1leuytt0+iD/mfbZvglDYkzgPOYcL8xj4tpfxrT2OnIxQ8KeBL
dJr60GNdS4Z8A0T+87Krt00nDuvS+A54aWc/o1DNIMaFwPhWFSOprjJWi6OuorFC
9+aunpcGP8SOu63y6Pwt/G3XiXlJsukrAMTG9qzUScuEv4GP9fn5fK319BOoxOQZ
/tWLOz4u0/QaOCv55jkrlPp/tfnT/ogsz7yW3m6BBsOMH3CHaqcM/b4nFwEHxcUm
Gsi74cHzgWXJ1N1E3kiENIUcfgD2EpzmCFhgKSZFXQcMgZ/4g1BHMCg8B7/uS3v9
su/Oi9Fbgvy8X8pfiSKfMqabl5tOpGs9PHrqgijeZWHuquAtnid5XLH4rxDCd7bZ
9SwkN2ZNHK7pXBwOCd72DfL9RnTP3MIqe1WCrvpI18Jh9DOQHiUrpvuVHF/GJNkq
n8xoyDYd0w+hAPi9jkTTO1oWFa4Vcky6nq/Cvf+0kWHw2aS8rKe8h+F90dPJx8NE
O3YHyIC6iVAq+Ju+YzUjn56qeoKTZVQa9ATujxxZoi2nKGc7zykbaQYU/1P1PfKm
OE3Fo4ss4vKtZweM8j1DwOi1OccfNMxRkUtUTEZ1eD/yJS0tOXFs9JSuRC1KJoAR
YKnNiO6ooCjKi+JINUtuFkBs2oAD9uHWzW0WN3nDTiDYCT8Dojyrns52LbHgOLl2
h0Ts411Knt5bG4EO78Y5JoXqf/kF5cDTcYdL78qPdsPBwgxgswcjUbylHB4BVFE0
Nfwqdk1LC0uS0kDAGh4CI+2UDCK+sI4W/phHeSiPG9NTIMINoATyjXM0NhufSr2Z
+cTGpSrZ7p5LjjgAv7MpK+OEp/Ld21gvMxuGe1jc0mNmhcqVCGBmkLSEQzUypOuX
YEeoXlJYRNHop1rJiuSd9VAXMoQoZWwgTftw6P/p9eWRIn/o8uz1Dx/tc/HQA+go
3ozr37dmrXs0XadxPV9Vrp/8y899q7PSjTyJ6yhYpytS2R113M0iY2w45rnSIoYY
HNMZgIMLGuN0zuhDRFd1QDFwgzznm7+GGHeJGzrD+OQ8fcxBPFOv5AwYTNErHkPU
WpxwKqbUD+BXZ7KI9JnCN4GpNf7tsBlHgMRtvFPpLP9d0eCX1R+OR/vSrJKf9TSR
bSRQ5N04crBldAY7CxJSFNKPtMgHQ+pYyVpu+94V/d8pCmvpdQhgU+DwMqULAQ5u
aEcIllkjg9yqVczGSU41Oke47We/S6iESRnAtH6Y7Svw3X9tDTpCWH8LNjeGt1Nt
EFT4ss+BRxaSR4iQsZKJXY7B3ACdRsoWQ7XeUoAEQTrxp4rK3d3nZ1jrVh4CKqwI
JqwM1ZUsw4nyy7UTIn0U3OblsyJAtELEwMW13GPTRUrx22JjTyZt/pycIz3qDV5d
2au9PNpR33ZjtA0+RVz28ue1efHjFpAbrqBGyfw75yLP9cQMXI4LLGKWhCDPP0bI
wvVwQY9gP0j/YZAcBCRu1vxIHHPZV9GAtQLEeDJsLYg8sDJrpdeiWE4es1RJyRld
TfHRZP39jgyGXF9+GdjNlwLXVFMElTDhoN9prwlHSyksWdiuBkEWy0IBFK2LKlvx
k8XkB2GN68uM6R9L0mu0cLMmS7AhoBKgM6op7m+rqBjzYJPuPn+la20xfFJXidz2
J12jSPyztSC0axiFZg/8hJgy+nEF9GqXm7NrY3LMCw8xvv+ezMWNZEo86dGuxUkK
j+iA6iDUEjciDA0G5Cjx3b4RiwyjEeHGt7v9JXumUjaw7FzuAlPl3bluTSgav4IN
nRPc5JcfHvSQ2DgBENQH7RsaH/ESnvMDAkFlqfDMsMKRcT+hWb9MotO65Ru3atCz
0zd0W47FudC0jDolCaS9LHUgD7PbmNvSv2zlihAdL22HAdVAhvsjUTxk492xo05u
DFIzvO6bf3VRr9TBRYjAYrQquR14reuw/n/dSbIBYiYUQbkl1JvO8d0AQmYe6KxA
ujrrcOnCysmTU8i6uv8PGiRbxZ+kJbWECTVcrhXUBmtEwIjrYRgbyyVqC4s6owkH
hnTZh/nyFeqwNfNMUQu4i4x5Zo76AvMkweHXaHZdDWH7IzkzDa0IJiQjE9MryUD0
Dn3tYHqnq/o7QQc9s+8puEpVVW164UqZF1dYbq4stVCreEYPRxiqq3KZc3U694j2
Hwps46UlBDc0cCHEQbRsgbUo4i7azIDswsfv7oMcw7QAq6hsWfd7spOg87nNipmy
X6J/BjTr6rZmgKjXtu+QZ4W/1tKa5TNlt5loHhTX5mEmNH5G5nDarJE7dVxUs52h
joSVAlGpTKr9QEzrJASN4AohvsWOn4wKU6UIF2IwUeMakAy5BUqk5MrFhshepD1w
b+RnC3o9CYo85LGsG/fFEkhGfHNAaIJMFEJg9PyXJTOo+NuRmczMVXSqx88ryR5I
FRbo7VWplF/NE4Q6BuxhVZd5rHIqdJm+VNFClCBjRk3t6q4vkCcgPcOLKE5ojo/F
NNn7P4697gXnWJAb0gT4Im2dNuXK4u9SWsc1ukc3r6RUOXtI2Ih/Tu03dhu2aLvD
P2bz4phqeNph4VRKwBvNE8kylMDj0KwQbyVxsq05fTQl9X446sTzbhWU/ntoVLX+
wFuy3Ks0Hh4/crw5IXYaU2o8djKJFfWovFUvEi5xoxK1gSlMKHXSWk4/1ZxdcfQf
DXfdWEhvHD34iLQiq3S05EWpa+F5HLl3CGtBQfltGBDGVyCnLMjI6BBFkMeYIdlH
0i+f5Kwns0HB1fdFILXMIhYaDCS3Tcv4sIUJn6MNGtLaf71kypwjs6uW5O5GM3VO
aZc3Uxd1/1xsdUrOTCxvd3xObd/OTiIVU6NzRRRDJBUBFttnuf9hgBcLaHYr7CRK
KCzcxnX/JpoA1gRKO8G3tvYqQrC42n/Zh9fNsvg7h9cPscyI7o+0WOHGsehtMJr+
y1quaPtS1LcWz3hpUzEw071MJbnZy3U83vHzvXAK3jVXB/rPwVnmZOSaj9UhdZoe
4lI49xiyiX981PYs0kPr7qffsynr7tR8Vb1Xv+3j4FURamVlGDMEKNwt2eha+m9I
i6KdEUNG2mBunJ1PFIJ2WZ/W6VjFtwLbDSw+nz8NvKlgYA9CsTcqTtZjd96gM+qr
Gc/jRQmbP/E2bHVYjY3DGSvUF1T4/JvHgrLMegBJ/etiwz65+mQaW4YbfEAfFXx8
IL+vlbUIDHMjCFAnGnxRxY11F+C8qVReoPC7q3yD+5oltBSk+k+lbmIt3Ms4hf7n
4dGEUWq7RkCTy1ig07TozUv99v/FwhJqLZ1l8EQNsAeXiUqh6EYzyOl6Bsa0YkKx
kp9dbcTuihByaJ8NypHTJkJz535/8gjYB1SkINuAOKu/a0gFx3KpJLb7GYzVdYAO
6gj0gDQeRrQon5s1hveJ13+IkN/4+NzItNf/qAdd0Uv6fYMiQ1iI0/ogsBU7Mqpt
Wpcn6f6DnVpRSAQhNc4aWOqZMHkxV7bFKasDX241rpgFaXQ/zQzWw1qO5HLAiMEq
g+IdO02ShBQKdWe+PS8enQDRNQEBGmEjs6+iQLMzconRIC4A85Y1QUe+5rZRE+MD
N7aq5KmYs/aROsRwcvHU/iNHm2jlas/HGmmenA0+84NGL6dTyXmRlLIiYOEsLEDN
lYmNxYAk+oK/vstAecLZY/82cr/ObBiXaBKFdJBoCd78V4S77QIWlGvmYxl7XZe3
wMwWM0XmiFGnNryjQvIcUGqrigZbgtPU0fljr8cRTIjMf52mmJ0omzRseZNr1DIY
oQp+tTsSJhDmfyBpxtt2bGaG7OQfP6VGAxPKKZK/TNP6GwVyx3aTzC1tdTCML34y
izu8ZRRL0Oz/9jP1ictZaJXheCM4jQp5o2Z37m0l4US0TkqbliN/RQ+dfep05qKx
ZnPohZH2TDDzVpzBgFo4/eDx2wQTT1PgVfpQIzkGJ6npOMJnkT2CXFnClqPf3JRZ
WQlRkzhUVCz/3zQVxxNaY/xOe0t/gIWtiUw3flh3ZkuhSRakcHWFiKV44sGO46Fr
DFQABgQCBIFnoFE7mYIXandArnBx07kKfogCPe1zrz958E2JGy+wc9Yz7Dgw2bOn
3ZlEvMbT9n0YoU1E6aZaZRlX3F0bAvIvgw9mwhX6VLTTJ3PkrC8+dIX3MKCgraNw
dNG3DKMUx+zMSgzQgDXAgH+Y/j3m23eY5AAQGFLjPTybB0Z49hr8i7/rt4kfkjy5
+Y7BGl7GGN7L4PkT6j864l5N3H+diPe7iKuDBX/EfGfFUQV1zfwFyEaFRN9aqMKh
ZzvTx0VuLaZRoe6w7+rxe+mu5sOvWUeC1uhhJkmc4+q9c2ngpdCJMTprJV3h4hdI
rQc5YcPb6l9ZayTnd9TAp05VGhMft7V2+0B4iD9ZXSDxlK4aGasXEdajjRuGNYPj
LHZyIytPwAgFuSYG0XkhSwb6GagBp7Jq4ZktM6l0zTL7DtmqVjtpPsg+x2tVl38s
Qy/JCWoRo8GnwrNi3hAKuVZNgkPYMjZjBCUBrtxSjxBz8hbAPxdIZiLkeKMUE70l
iCxun0ybTr8PFKsGerg8YO7B018ysoSDniLF/tYvB+5AkhgRo/4bxHdA3mVuO2CQ
q0uYREhh+RXkaNvcpLJ1DMqvZ64cDRzwQ57KPvghvEOFRkHNaGk5QstyOTM8d+dE
Qy97Expahx0KrLw4NWtIu1hesA752Nanki7WNLUmOKJ9WH8yIoqcgFQM2YtZavHz
SK3gQUFadDk5VWNHHJfa7q+h0r2KotqoySXfmAm2xcCFJZEk50O4uRlYP1zL+bxs
2Hw61VN+EVEryv8pAniQSz7mV1+WEVeXKVs+FPxUPhlzgBuQlQjFGNSiRqBdnyNy
dk0RZbjWsvXUNSbRVXO3q9vbItFnQsI6nwo769n+Sas8Bd2Di9Ln7A0QrJdB2KJC
+nVWOihpvZujyZ5IxjBcOFg+Lhfxa/0d/hpXF2vSb412/zeKuBC/UDtIfHzsJwvy
jT1YkYNryhPL8igpD0R7SgBUkd4HK559drmrxUHEMYNsJDetWzPZQt0OChkutpqf
0bIqIaNaBsN24HJh1M94GtsOWB2+o8p5/f8I5+WqhzPLTpaWmCJcjIiN/Kk2DmRU
MFJlo3Rv9PgbqRpJV9VSUrTOVmPdkV73HTYwAJnlWbRlYoclEMvqv309s6EtL0cB
XuyjBKCWOrn8xsuA0TNdo+W493WfOn9MTeuxlDCqJrM/l1e+ojFY8PWqxGDF0F+S
UJHoC4U8FPVWzvN5SCwwAruZ/55IVOieeD+aPB5YPZpTLTPDI+/1vIPX3nZk905m
JIfz/I/8LzXQ4A3EuIpiekv4QVbra6RnQf+GzbBybIVIYrZKl1m/UfEwUYHvIT19
8xgiijKl2z5+fRQAFEfIb62+kZTqAW0z8Wau62a+PLD0L08H7e7p3kJFPIcuPgiC
Bl/FWESQhiLc/fSjBO3y2YZcFZ8uIn4z9NQ6MWzguCsDdrOwmw4RdKx3G72IG4Mu
WHEeUj20Owdik23YuN7M7AXyaCurAkAPpLX7446zSbvwAbzG5BaTGldcrBRf6oqQ
dHFTP1dfV/ZgY9qudOepdQKBJWv5NcKF7TZnt/Q8llwdBWYlyFZ/itJnwPDW3sUX
6TOXYTnH6Su47WjpaVcAx1oFGW21BZZvl3NuH1KpNTAniMpOfkzVJCIO9yQf9T81
XYpGSXbuq4641m7H8mnR2BLJpSGwLAN3dPsgGl4UlClehh5Lq72M8f/T6ItjUzWC
RDGagkVk3EbYHy5UxuO1Az6lm41o6JeXK91bjkY4awSQ5UAf/AWtaZRgOBYHaQ8H
l6CWbMXM59vJ40P413MwUahErnH2Q6ZdVjVDS+NUPr/1gPJmx48mfiGa39g5ueZ8
ANa15BP32cRVsmELcJq2V8eg+RnYqYCzTPedL8SdKWs2IL2JEp6ogW6VukwSiMzK
rlB5OiH5HjFjgf11q3Sr81JHdudGi7fFbeO+i26yKv/UoaXDPeAc4+iuW8xQIfEr
sEGck8Xaui4VNJ2QAEkyHV+jp/mS4zwSi1HMi5DlJHocAoZTq+AJAhusXdtNeF3y
Mfjh5N9DfVJ7xu/ysKA/0KnzdxHC+RV11tWFoQRjCUbVIAP6pA3ZbZK6ORnDTw22
06yZdB2LUhoUIjdAOQ64cMfJiHcBazki1oasM5AjXJ9vvW8a10xBKC+xIVLYB33q
fB9dwdBTZiroGT3+tk2UjhGE4I8TgFpIi7YFvEbzv5QdBzVjwvdvux5kw2OAwkso
9aTN5+hyjZpegQQMF0yeA+g7nMJlnSpCRaNCijYZ+eXwh2Iq+j5FBhLfoImrxe4z
ot/Axbew14zdg2GKvnPr2sUJKNjJjlu0vS014K9UEoj/zQ5gmZ9AV9TUvXYPzN+N
06id4RXFmFObj3U6ewRk61hPDMtfi6IjCkzP5X2mNoi+XyvNtHojNxGMfrO/sxfi
rIbJvajvHBXSKT/Yho5Fku0lwRB+0sUNpURj0EZG7hJ/WH/m1fqO/IJP0IioXl8R
CqqulzPNHo9O1l33EShy9/GzNCUgxx/HgrMGQ8947EXEuIFh88r/t50sw2fx6nLQ
Zr2kSQSTD/L5dLRT8Bd0NV/gPkvGF13FtEucVsk31v07PZ0rUo+5Xc7Ck0jnDmdU
cELzwhJBBQSRtSHCtcPboe5cjruMqze8CZWVQIjFp8EuLIqYVCw2i3NavNItFl7i
ZV8HFep61THrxFICzU5gsxqq8pmDD3JX/eFFBpZoWOLifDA0n9DRcht3DZ+HHdWG
lYOXI+qc3OeIyvWcJh2P3kpwIxdBvQlRVTWvM9rRjTDBJTNT/LZYSUdB/VJz4UmN
TDGT8Z0QxxVHuNSfNWZE+lFi2d9RwkJXxeoCCVmg5GHpbLahUanmeTameJr04INJ
zd6zxZoXwU0lF9Hz2mbBkuIs7HuOLHzCBSNe3XmBgGOvD9SmTYCPy6NvkoWfBnmz
mP18UpsoF/s1N/sADM9oSRW6HxcZphFN7QcHXqeicexcikw1txu6036T+fdgaNr2
HrTDMPHw3z+3TOVA5VMW3q0bVkkOm9I3XM6zJgCXQDQh96aNuRc7vwQI9TJ1LbUc
T0DDCmpAcVhjOYu3cgjLVgtFlUfLMwL2Jcm6jMgK5B2++MdWrf1OsxWGRa954rOV
7lpDECVfklByEgyUG1pQ5LbiBDjq5fjeiQT13nKGFyiXF+NcnVFN+h9PFzLY+MEg
3dyDMJhn6ajM+00278cjd84d41mBze1cSwmRTuDYeLZ2NCvLzluiexTvHTtCM0ni
px+BJUYsWMsupx/X5XXEgY1XMR0cz4fkw5Jp28qBjl8LLxUGf7XGrviRVB7LaWYE
+wmc6bw1si/bvcA2SmuL+lLkcqt3DEdXYxYCKg4Bc71vEDqdrf5SdDMyt9Q8e48h
rwSSYN7MVdfqnlJcDJsKhLlU7RRo7VRZVeRJcQQ9i0Qal8Cv6EbGnBHv1oFdEC/Z
+oIW+La6k85oxv0ECfmatUEkq4+D80mvOsScBEIkoU7/9Nlm46VwUQdDkWaR0yWf
rHO5cjMYjXxxrSji6LF1OWnAKQnrO+3DZ8CsH80/0UUNHNd09EdrV8xMSjPd78j8
Wur+2Hvtawg68J461TDGNO9Vcy2u1tjbdqYMDW5EoYpg59TeWjVB1R65u9DeMF5F
+7GuiZliKxL6T+ISagB+Ni6UJxrUy6IiF0zHTqa+hE6jKAS5RUyb07hIKV/0FOw8
Zn7FE7X+N8sNHRgQv5GSQ9+AFDLkkMxh4TlycdqznwZ4VRAq6r1rcaZat/r5tZpY
nUk/9EGrbhJdvIgbmPxy2frwd3TFkbnOI0P4/t6StVF7yCpfGh4mje5jWXZd0FOP
KBjJKt1KO4HZA/iO1ZxksEVbl4U6BfnXxpbPvzbCOam883xdeag99+uTsyzJOm4d
h6AUf/nX4tLr1kvWKjzmL6XzGdBPoJhu6R8/R5JTiEFNsg6t69GjYnmzwh5cpWCp
05LIcWGJczW8kGs78EJXwJqNx6ijBiz7gFYWXXIjGwoeghbUh4lXgZpP35ccZcX1
jJAj8csmlV0h/SHa1kKQa2uiGAFELvOFXSAtkTYIRrg9vijQLOpckH7JFA7+E8ZL
/dVjILsYi0zI4Z7/myDDIwtNtr2DqY3yr3XlhRuFZmuiLccr8KCMw6ZxO7OwvDZv
nXM6d+xSChb58M6y9F/JxmCc3gCyU6kWchdftjOwXDg7jLJQOXJnFKE8lc0Kt2On
royQq3z1ecAEI7bsq8do2Q3m4l+QBLXEX4NnunGN7V46y230CuVJ6nHnXepeAWMy
SAN1ThtAxMJ25FvpNmLkcF9Ua7gW7g7vJTy944Zq17lIuH73bpqpqzhX5Wai0JOI
UQWES95KinUSa3Sg/qhAQKTg04FcmNWKCDOJGZuZg5Zzw32cn2cJWpjVWpRFoS1t
ev8qaptphub6WF6xZOIwhkZ9nKwe1ot9ArQb9mkymCZaN2/BcQkNOWoesOLi0UAM
sJ2bluRLuj4PfeWAPkBY8cWAcPcvvyrPyqzbSedwZD/EuWYBu5PGJAiuDkTmlMHo
fDqUs+Eatka/uT/zTj/iLusBR6luKG/GQMN/MHjgc0aj1/DXwOe5dJBCo2be4QRS
DPsfNFg6lrs6HyjL2w7hz97frUjEZ/dHy2bdQabttbfM3173w+kJcKvYXJhlLnZD
uvjubQ3PaGhBukiAgw/doMqZ2M1WqnCG+0r0wiT1dl6WdQXca53jHWLkxl25OHqU
eyB2l38FsIz8dkqfjCxj0wQnHqJcdEn8z1sYQBzgqZ/xrzu1Ul81EsAfkkvYFw43
zogUyvs7bRJDvRHOeuKHyAL/uhwYBclGImgJzUqBHa7LowCCXz4wlb5TrzANjppV
TXap6YxZ9IYuRpY6Xaah9GDaw6NcFI+EsQTRheSulEqhRPx+lBEVTi92J5PcLtbL
u4OGyeMKJwod9lpPpZHWxW4WwjOJkbXgzjlyzYPQl9i0NL6Cs8GTwSlE1qX3bVn5
D8b6QXvjJIs7+DZabjPA9UwHsIUOROgFjfnvWNTY8KZIh7QWdyhdX9buKG47RHKa
iIkFtwFh+iCYNh3C6dxP/istBIrQufJ6bkzz2xfIyhVqc3unOIYEj3SFXE5r7hiC
Y9QphUmSMy/aE+K20JHFjkpFrRXvWJo+UIoFy1jaxLiHKRBv3pK+c+LXy7jgGGCR
Z1XTT4nRZQO5C3TW3JZ02XposcV1+uWz+35DvfDmiAC9lQhGY+kVPNEDNAMni9jh
XcTFndWvW0nHggX9Eu3mzCtw0fttKyagmEMx/m+jC/rc88THrlmms2f9lC/p4XGF
24rH7h+8FZAIH4v7/PiHihaBlGgWKMaasvSK2T7QopqcRfqXqaMplW6rNen2aGQ4
39PmJTgtXi1WKnYJecICuRigCysFudIfG4FjYBEfYPZnSwdDAWCZ3MxCmlFpjLd/
aqsrSBRL31PzdzyvijJ2vtVhhAggIcvgA/9aQUmQVqVz7CHb52iJr5BS0sRsh8um
Jlx9ISvVAxKsi0DGpzkNxlgSdRIQJmZUZCTvw2CvAQAjUBeCwyNlvJ6p2yYgAuzx
8ePg3agcZk1lowE7KVy6ItZ7M94r7iF9dNpkM965aFAo1jvMBQqY8NHU06Umy1IA
e45FqEufQ4fIywL5BSS+U6ye+fI3NcvKduQEcjBrSPf3KBLGZfUX4bSwdUzSoXdJ
Q763rXJPywt9e7Zf3hpazkO8oZMsie2HGF5/Kqaj331whfsXvkSNV2+TzhBLm6Hq
J5X9coAwrCV2edEOoP8y4c9dUsVyjs5Ej6NFReCC/kQF/4uyVIFjT6Seb47DaCeO
WnQVJUjo2QpzNaPdan9xON6bVi5jK5TWnkz3fOdvTWiJXgfXNnPWv+6p9Yt2I3Ux
J/rPE7k6pbnWqh4/wJK869GLPUQkVCQdRCZg7YlAcY38cAw9y6mr2GLYTQ2hMCnD
I1uWahrzx/+bAk2a/J4E9XsHMDHYlZu2NLR23z4GAvGIW7HWRUqvM/G3OFhvMBfn
ZRwCFWd2d+WNIzqahG2bw+onxuG631wyLZ/Ss6DZkZibce76EcoklYncZ1Ky8tWK
Myb3WbjyzCsyfmDFPkoIJZJ+FJdbuafayzvCS1lAF5LV4wWfxHDEOeG2mHAml7zG
glr4zdUE6tFwlJgc943hoh0F/nPLvBdPAa+VOwCopP7Tu13qMor8T9/1yhN+jPJx
Ysz8xbKqDlRSoAoTsJD0FJI45bcBS+yNyseIvwfZEldqU1nrytq5685Q4h9ieYAE
cUgFbVY/e6tpSH1lcLMnMCuuS6ON7zWiCjNk7YpUYNu2jYkJs6K2KjkkkkgcpPy1
8NVrkOb9ixaUr+oPa+uiWxosk0eYHtsfKxa5/bd+82k1T8eo2QKgvzd8Qpfpckzg
ucgcxOZINQG+TAQ+8b0UCXT7zHZM+WKkWAVTSkFo5X+6SN2NiDsUwcm9lAldio4U
o79pf/Ykk8209tunOclQE/UMJq4g30ds5HRqSMV6d+27B0li6ha5RaH049bJdcuD
CjFlSTTKpBM17Aw0oXbmuBvA3UUWBfv0uKPXYFugmtlu7O/kIFL6ODPylbSzpmox
4u6Gl16N64GwlczRqLHvv5KiOI0SD5QoedWgqd6bUiM7GZqiwaHsolrP+gAy+VH3
/oslvz3fYC2T+Z87mT80cyF4Gp2R3rcp2bZpaFjKgevrQco6bgxU9vFpH51sslaD
uDJGwupAKWE/3J5c9rhXKdUx/ysdLQQB2m9KgXOx87Ay+BTFiUPIbYtWLmggjjBn
28sKFcM1PNniDMYk7XKHy9bmGY2Jw9Q0Xyiu2a0zad2cp05a4SRjCUgeO8KzK7Xg
8i2+ZxasgFSARB5esKmac7XK2MQIou8Lp63XEyL6bhyk4VvIN3HNxBiaJMj+IdqT
KkK60TbcgBysul2ecpKVBkPRWTTBBw0vrEKHRV5LJv68xVvuxcbNm6DBzsp/pL0W
L41HRX0kC4j0iPRM8Z0qhK16LB0SkcR1gk7taMbGj6SYHHfRe6uD00YpwLsRgPgc
jW70EyklAqB6lnhteXJ0AHMhBsOvUY0xewsbc7cqFm8Hh2f6m4eEEVDNpI6j8Z66
sJQ8HqJ9rAHp6/AqtZLSXS8Z0FWwlehdsFs48pUrG+NNwgmtj5ShxM51+qE6fXm+
+Urim5YfHrUY0sZPAZGjsBRrFN9DovLKVoIITISA6QGjc++vQyu7//0vxGsKTK1h
sxxldIlcbfFgu1yara+SokgAXoHS+aUDiRHrZiNRVyE5BG6e9cC2rvTqRPojF3bb
/5pIjKY28rzg7NKllOjg56cpScWa+O1Bw1MCCC3QaHzdiu2QKMxQHTAuUlsOzFMF
JePaLw1JD5r47fS2KeIqzC1SeXewwWvIjsY/tIjWo2XX1khE/YMhskYJi36uxYwn
boP9Gp6Y3tDdvOaUDPBbRhWln4+KOu2ap/oawwJdJZcHTLptVsAk2fAvojFHjYxw
oKdUL1MPONuPMGo1CW6G5/DNGhvmj67pq7vuAL8kqhLpSOL8EsXOYCcI9upN4oWy
UvP5Xz4031HrPxa1a4WilJPPqcBsH+K50c74NTvLTvzBBMDCpMrQWBI+bejxD5wl
jmAhFlAA0TDjM00iY+w/1M+gUSKeOFpxZQ/9TvCwINXJ1YGX3y5vcmhdGpyG3HoG
YAbHVCYKoIHyDyNc2ff1wIU2dFINldLA9rL2AgnJIduEjSbwvLLEK4STTm9pykGB
eNBE0gb943sfF5Lb/bcVj6BGLy4Bu8MX8m/fVfBIpFCXErw/RrRS85anUHvsr8zQ
LqVcg47ycjMNkgd6msft9uxF1Y7vH5y2+Yr+smwDrVLRhDJd5jzOt5HevWBz4Nj1
nk6jPt7in5gC90RC/smODY43+XiuS3OmanE/mgZuRHLK7hD70bQoZlBbUlTjvh7x
GulZFpnurDXbyszjVxrmTMZ06n6LH1LqqW6xg+xcpsfpsBeYdeJrt5Q4XmT6hQch
WpXvWsEPBEcY4SrU20HhgPYTaQbg3XeRRdxubRTCtC6+1xnGfT6sIvFpWHuOE3dd
3jSP/i0s01X5TZU1l8L5KjiUSiwsotLjdU21Ox6ozqRFxHEzeL1xUfYs3+FHaOYq
6sj3YkaljrS6xiZhX9jbRBRplwQoPCOxsBjoqdKw66IsrsSw5UEr0apxiHnMSejS
3rK/EMwLBSB8Ab7YHdlpiYuUANfrlhoQ3Hs7lcUG9DO/h7Mee/S/gAypmK3WSaii
xIB78EcLahl9p9+ngAUiUJmo4XXW2+rJxkLh7++Lcu9hXgkyQUC2diwhUUjCACZa
M910LeDxD3zMWvm8hEBBznCDkAa2ovkglR5fRDT395CFXLZN0UWovCy4UF8qhGiN
2a7Vza+0oycqVT3JNjkQ3wShArYYgmA7L6vzqfaeu/VLx2trK6A+LbBHJWgFxhnU
1VzTR5kJcvZ3lbNZsy3CTIje2WlQWXCTS4y/JhsUYCadKc/2p+mOyfcuh//ODIJG
5rUFbs78lOeNsj/0qeVCeeZwWEfkOF8bU/tFYwNkFkpjMGvjNKFLvgMPuf3RnH0e
k2o4zi9rHLVUc/clT0ILd4yOhIP1CEAQ5ccgHYKT6BkLHYX0Eu3HuZtXHu5aL6+W
VYapsrKKCq++xARyn56iJjrxMkjGHcHBF3seRstpO4E9HzbfVxWvPcm5BF7miTZ/
H3JYjUCvSfCxYEVkudcK+JYApxLGSVQjIa9PUcuF8uyflLYN+Vw97r0QRVc9ApmE
5LmRDu6iFRObNMSCBGfQfk+oFa1L6UdF3p8G965zVQcT6FQ4MqXAHBRH7Nn56k7X
JhuYJEy9ehmIPEpwxqXtSdttdozz/2ne6joRE+6WhjlDXF7t1BjwCSNM1XlFCemR
howeb1F/8lYAkNKyj9xfy+p9OYGahp9Md/j6VKHGDOKS0St3HKKA3BFVI3vk7slo
eicA7+tbgStH5wDyCx91cWjsd5tkk44YDw5QF8+pDAR+m4cmKjU/m35PqbU5ia8C
TtGi3khEwfUOhWJIkL61IFekDdV5cDOGVp+CmDVU8JDv3oBY3Pm7ELdPb7JrnLzF
eMMuNI3foKlqWWcVBQq5CfqDCFDjxyjsgh9ZV6LEfh8IBM/wk/MqPcHFPJvcaox1
MZ/fU6QYxoCS0uE4+hM/zabVt5HdCrTJ2SIbgvfiU8Q4Hhvzl1vy2aLo1/sm/JBK
RjkC5XNHeISQUESRr8d0he6F6M/kvKqLxGJ38QLuUBlq+iCtASG0R2oFfJAGXNEJ
ZvnDLPO5hEedCh8uwCsDBqxH+AVA8XOrzoCBdc2Ekkq2KUT8sBpzzzRYYIiFV7HB
des8G2MpnnF2mfDAvWlUVcBDcOF6268TXkzSa0JK8vVjuEgqZL7Zw+pIOcYUgmQx
xuQpI0ZvXxRWXM1/Z458thHNmybvkNGvypg1ocSWlAtqPlvrW5MMNyHZ6FgFWux3
tKQBUsA92MOmO0mlh7yx/bP8p0pq7au7rlKRtx+6LjlUfSPOXKEGSVNAPf6O6XGn
p7KuiZ6x4EqylAT9+fmJ4t9I71ZVMXc2yptcWOgsOYlj0JoOw+NYY6B8PCFh2vH5
hW/aEAVTOUSizsTQLs5oOWE7SdcBd5DaM5hiShcrPSLXPz3wO29VQ78UoI9Si75b
f5lrMEn3DXdo0n5s6DNLhGmKkEZ7c0QJrPSeDyORmnZxjlHaCP7vht0Tb07e0LY4
5kq94NoG3qs3NSJUEF82Pi0ZrIj/Uil2lwbpaSPbOP91o9Qgs9ktc2Wf3OUhFhUn
UUieAvxIp6Z+Q4Ul9Nr4nbJr1Cda+2tfdGT+C4ugLCyxf9ZDMsm83dXD/QTsgdba
Bh+tKTAlLDeWy7GGGe65Z27+0CayZBgfSmriexDQJJ3gCQyUFyCa+2bGAsWULE8z
q6PQP0dasaKUYHIAKR80H1Oh44F7zL7sWHU2oDmmZVsYLpB6TTeg5ktzMtFXVoZM
I3WkipcVcLjkPayp81f3Zx11UWHt0nYEHINeon5YVSFJmVu4uaB7XvtKNw/M3hm9
MOWJamOQ8vunveJ2qnuOz4eKeFjgHmAnSjJ9HLUWLXBNOdIPoI/u64AjfFenM9tm
vsUBhARQ3hY7t1PSqF8iuAyIALtQ3DwvJL6cPHvFn0dO1RvBoc73SuV73vX9sBpn
Qz2XhUVhqGlFHYJTH6BRIZAiu1L6Qh5JLvcRIyE2wi8zL/nOGssENOSO4/stY2OC
0bZ142Jr//N3hf1mgmMZb/qjRn5aynuiflF1+SmyAJJIGRp5TV0SicNvLCdqTa2W
X5frHkrF1pOBgpuWfs8pn8zzP9mBry9V3NcNyRRKDrA3KHTmf6jSuRNw/mhUir4c
jW4OxsYxXv+FJ+l1oK1OfkOobc8SIwB8xey9JxWFyGx5srPh3MceB1NAR0hpD1Q8
3MIg9bbPodWtHWXcdZoRjxDjye1VzqYoBoXYRWqeM4ppLNNlYUkEUQVmWUWo+owD
RiQ01ORqHs+5iPtQLkIAer73g+3JLTanzcMGUsEAvJmDlj2CnZJRExkj58NYi25F
4IjfQ9yoIgDurOoti2NP+DzqwLFHRPPKs8BcGJWpzv7eI8rv78bcprANjBzxEd3d
BCcxId01JwpN71+23WE3HJe5UC0RBkN9UEsyR8VdZp7MfmFSzafAvRmzFOAgUVxi
S0D+Sl6BpBmxT/b0w0hrH1DYr1Lr3Xbfo3qFomk8Fp5wrUXSrrX0PJBE6hKWlMvb
9NVN4O4mN+qe/jVA1V3oOeAwKCcKN3wsHku/WRq5EvrwKTy+QLAwBb67XIsjNneN
/SqLjjUKOmJ7cC2NllKpdl9BvJBcvbPreKLmkteEAQlRkA38Cy4WkFOLU/GMwTG3
1SFWvRLBXwGstVZsbLZ3ChzJmBFOtahTXqjTY0AgRJcspYyymYwvPSCsJ4ctms54
tgYjfeE4FkA23/PHmv1JZ0Y5BcnG71FXnqDBCD7YDoV447pxApTMTgDOu1VQexZj
KdJXd/5FjHxN8WcyGL6z/Pi9oflKRaYAfCH65mhqHlboN0R5AIGR0nDpwr0lystK
yGvX63Ps7Q+oxcbenwG+ONBocEPiHOCenmv8u+q6W4tD5Jw4SGuGsICtwayvDwe8
de5jdHIgB9mNbZHzNgxMLVFLEHSNjUBAAZEbcotQEllBd7xHiQaKH9nCHz1qE0MU
XFEIMRMRypughHiJDf7/T5Djxs7ULt0IxNsoxV+o88kYH50/SpDc4zwjCU6y1RL/
JIRtxJX/6CageryL4Bg66UD3Xv2lhCZjuDGdOPwGa5KRHlRweC4PuvqeaZZCHQFT
ofvdnIRb6eMCtu0CeqSp9me3JVlCsOUqix5TiGkpSOv/EBqP/ToBUnLmgzRfl+Pw
/oLcL4pgCINzZUwKBr2fJxA+APO+ajeNb1pXJFgsTNpPm7iykcPtnULqYwVRQ7OW
xeu5GPnkdvjZGO2YtERG4DkamRmsEQZrR76RBq//wttHsBh9Km5ggntdX8NaPVAO
5xm91Qt9C7cuhHlMKJuIPqAUX00HzDSk9Rtfz+Y2VSdBWRylwRDWjE062sWRs7dL
PK5LASqFl2bu22jdvssjPhVJEFfG/Yxd1LBQIjXsGwiJxfgEqFcx6yxfPkHugFCU
kKZOh4bndvlenmy6mhIbFfnA04jJRdgGWkJmXVR/iu6T5fZl+C7CNndEydWDdOnx
0mfy/dsyMC9MydJGbLBuh8F8HyL6QWy1pcj+vDN3qhE8V4p9VM6TzrxkPsZ1VVfp
sFNoEYSK848TSVWqSqfgCUUwPWED92L0uR6G1qlPgi/bGsdCqydRnkVa6Y72/ERu
3jRuSUSFViQltAZmw4YrsF/rqEu6vdE6k9643sZVLj/jyKuqFqI2ajIkDFsNsSra
HELbptV1+ACu3LDSqcLj7AsCmRjDl6tvQvq1g7jXffrw2OVUuvZQdg6zqtJ15fuf
aLo7KBLzA6NZVIeiGMjz2c7momE5p6nG8NasDALhJzd9Oeofghy7PcFB5TJnNZba
rfa96oE4prOqMjmdXsMmAL5zW+uuyGlq9q+kV7YpVwKdPXLLLm62UuEfSYE08Wfe
hfKo2RoNpalM4fBq0953XikfLi2T4mwUF+f95c29kT0U+pneDnqhg2BYJyLvvSDl
KHzB5BMUB1H/ujjCheVeiyQWoFje/OFFmxShjeGwyMW5bqobWWklEN5BzoonSOgM
ROHugAsV9uYJYppC4PDAvhPmckv6hjIjUSmo71+uSr6PIdJQz76eiTPBk4/3R+Cm
x+4HH4Clo1m4c/U06rai8G00mm62oboRWyYtlnJbmIbA09UY7jjdtXQLDfJSCfJK
9rOtxzzKpnHB4JwuvmVsRHi5gQ69mKrSltNHO5WJk9nKZxzJS5u6QkzWVqAzMsBP
WRHdsCL642Lq9nSYTpgykXjgglc+HXYnieV8V7kDdLOFP2phoEvsDexPdrWx3wk0
b27hUghNXc4M1dwUKtw4VzsDS9VymY0glmNmVg1fza6SG+sqQtVmSBAMLYDgf14f
exZ6KW+bqtdt85+rG8kyDsrut3pKJFW8zQZHdXXHSOVJx2TnmPeEpGjIjd1ai/+H
I73qrrQSqpl4FJ91Cpzrl5UGw4ejI5gjxWTWZDSifkfRIXPLI6yJUnnpceQg2aRb
QA1MfCELC2hk2fbzncfhYjK61KIz0FZqFyMKbRjYCp+T+7gLCUwTYwmglPYqzSmD
RSVZF9bnG7KVvyCCVO9QcXi8HPiql/D/4LXL/xHCLvq7U7gxjohQH7Y823ss7xn7
q2TtItqGhCvfyR+cQ/4Q/jzzQzpvfF3EEbN0q3yyKFL8gj3g66PAuNzG+fP89XdA
okCJp/E+Xd2FdE3+UdLHPqSjNo0ZzW7JIIDql15SUx02ukvBEf+i5gvIioEu8Pd5
c69L9Dv1euyOAVK7HuXmXa+xdjK2jTrCKa5rn+mvEIKcCm0+VhZGc5dRLdkg5/f8
5ghYANu96U9ruHo2DwFEbAgcbFcLWKhc4CTNGsNEybwMogDAJk5TkoQL5NRvW9fq
iFhmM+YB9mTIFXHIyS8tClQuUT3h+D30TALPNfYEpklPUJwSbGvQX4SISxluU4k2
zm8X6Tru9ReaqjXbh71iIiPIsOZevAOT4DuoWJUdFuWGhqs+JRZLWwKqd+mE/yDl
2XdumWxn8KUSYXWZ7cppPz1YOi7yJ3iZZmAlU/5D1JR/EysuNXepwygKkc7hN54N
2m1xNPSh/IFETtN7bF9UmuTDgaIJ4fXXR/o8GbUXPpFBoOxICcatzz/laOhiQJgp
YNkAU37eQeUC3bxpekL9riSYH/wAbvy3ecfIahrrnYdeygeB71Kwm0/om+3q5AcS
1jriW9fkQJ4F/FCbRS4LwVfJLQsJmI2ZNGEPOVsRj3gFTzTFrhoBzhPTERidem14
f1iemlQI1INeDxEBMNdbr5vBXrUIGKPj+kOOBjhNtkObjPnnVmDB4jNPDRQLgoLh
CHm9U/bgRdA1HfGLJ1tVdjFpQAvr3VJAVSbTh+wxrnycTHkCblIcEA4cELPE7GOS
5jWS32VLQ1y+hsh2kGL4w2sd+9xWnG0R3hrCtvw2wN6N1/5Ra7b8iOCH6W3UGXRb
n9RWw/1p9irgtoEmClflGx00SdKHpDA7vPR9vj/6kbUEaM4gbhLBdkP/pIdxAlDU
B5R9SRC5jogAlmKwKl/HFdgkL7TIX3ZRV5ELRaedf/clVnWGuhs5SRU48m3RUeQ+
6PHoug0vdE0CIMfcdP9KQFe7wJ+UARYXc7ykmnQLKr9oa/zDcIAUY9P9WoZN09/h
8yA+ToVEClKeJzVj8T3VKIISJs5LTURIb6ADtNtBaMHkT8NBOF1aSXMjPC9r9lfk
YsLMviZiZE1AgzacZe+1Fpy6EAjkAQB+Wxz1WNTBal0H393hjXtVJ8emqR9JWvES
rrciSu3/U3vfU918KYX/BARIcRb3gsJxlOLAwEB012r7IQ0wx+aIHlX0Rud1syOF
a1H+I5Nt21dL3jAvExDghtgGyjsxOd7U1hfKx2chgaW0+BDvyRP3305Ye+dLIUyC
4xWyj8MtUUp7KGTezQYKlMTffDEL056EKdyGeunZjSE8kI91l9e5GQoA0f0vz+2v
pY0u1Q57XJ5XFEo5qOxoyqH0bZamm9U3TbjShOUiMh8+EIbNrSOP5+YftglTOvrN
OFsYyAqTIpV55xpgm5AtMGaa6t9abkt+QbYVH2M77szGZhSy2MVOA5CWUEjfG/9t
wfhRvL7qN56BpLWW8KrFFB1ed0hsglHK9q9MinzSeaUzyymCanuLd/KNSHqb54u1
hT5FhujJvM65FS2tfL5fyYfOY5UqPRoSmA9Sg3kBKYZCZr3f4D78jv/3v+AL7FOf
+DTE/FmZu5PHNpgOH6A88Lea4GcBk02WSysLgnxAdp/G4HNhdlTxPrdGqfQH73bx
192DXfMGYLvnd9UdV/8hFce8aJGbbbwmUyoGEP4Suwqd35+XRGbWRXYOOJpEmWYm
0JvR61Fz4f2zwJBtwKYAHlWzn7sfRwwDBDhLOelh/6hrpMLqg6UfUmJ93JC/f1ao
tslZACXJuYWQIlgB1ig0ybWn3CSjBJX567O81trViNg3L+Wi4DlP8PUlZHh8ocJV
vpaOdqMH2f7AwNn05Sq/27oJSB3KvKDS+EZDq98obMavj3ulONpbugtOhGgT0t35
ZllZza8gnVN8lxMmQX2Gbbvoj3POuUgtV1gKpqRKafhppsBP1Ul0kZANYNENBG7h
V4DZ/Y6I3x0ggGrV+b1zjwCKld100zsMjSSb3bLY54ifKrMGJO1a0Bx4uQIKTcqE
m0k1G0/dgxmgHqTNgM/pdz0Y2bQt1epnEJ1J156DdQJmhfYJyObsvh14hiKWRWV4
Bp+USSOnSAitVGPYLQB2F5EHtinNtW7FQrzoophYiS188N7i8/58luC3TKX4Ax3F
QdWFvFnRBBw5yMiiwJ9O4+tbj1oIk/FSVnJBYsq2xwSpUCrcDb2fnbPNGuNsDWe1
I2zrjrYCTnvG5LjjH7BFkY5IeDW4CKrJGgZ0ejGoA7VsfFpWYpe7l4aWEQeTzIk5
Uvx1lRKtNMiy5ZNytVJbyKu90sTrpOS9SFoUHlaXAWi3UZOAdAP/VTlW5MqapasA
wuZlMEHRi4MDOA8xXwjU0BosSmGih+XZTU7STWXk5frDXdzbJ6FmvlEbMNJ3F4ig
nCSWjrlSjGNjykikxEfxMJemyC2hT5mqaVU6tWYOXL4I/WsjMtH89gN+7kKZfpq5
Rb0iwgqS3uUYkfLQAsi1gdIf6JExqH6DvX4gSyDwbGkHw1fpiXnFgVFIoMQE+3OJ
IhCrWyvu6k3JtZ4cIDsvbxlHghWZMPik+hrDjpnJpHAIum2mIhT7+M8TWglxzsI/
687Ietnox4lnJEXrI5RYJNcj3IMAGAqwaKP2dd5DCQIQC61+N3c+Ja8UgBntNphB
M5vOzFzD7/8s4mK8XqB9DW7u9R9XO2l2gwP+LUtGzwm3MIto7Nh9bRDEW2AOMupG
8EURF5h2h0xSqcW9+waRvNnrIuiGRqGiGUK/3UMRQv2O1joiBU28juZDMVV34foD
8D5daZNPXxOmrWZD2LovjOO9MagJglH52rXr9tWOs9uTQCmyduyJQkxTi6HVuwCp
yROt4PaeqwMrZH+KEqa7WSAmcc8CswWXytegnalI8gNLOY81hbo4Hhgo58YlaUJK
xnzjIRwTz6sMbbqJzVpjWEdk6pSpNg1zZV5tVXD7E+Kzm2wAMbvseM1Lq2rdouu8
uwGKBBvbt6Xok4jCdaM9icbDJbfC8lb3Uaw5AZyq3HNHxwLgdNxO/YkuU6zaXqO3
NQ2eMts50wGWK4373zqSSUsUGPLVV7L6q78Ct11TFknGiS+R3wwSM+w05uXAzg+N
/+bMoRU5PXfLIzFXmrehaGJvNBLruxdsS9pf6dxCcGrkiJ8Zu1xBDhWcVC1OhK5w
gLc4fEAG6WdK8YO2amSy99xmC5houb//k/5JTn71Ak5xKhWdzCMKl4+j4uaYu+n5
qQweWardJwOCISZiTlRcBkNBt1ZO9z1vTgzLryoICYiPUVozkqoUMoxtsxL+9LVF
XrjXMD4ce0CG+eR4dZUjH8N+EDZz620WDOIYpw1sFsHrcswGGWzBIWQbs15peAsH
XCzf641kTVvvwLl8X2iRt0hKBzYk+VFiPMVhgPe6dNY5t7KGBioKu9m6WcnBNimb
NXYMnI+Iv4YkF+507yI+dX4XDn/ovVyVGnY3kqlMUesYRF4+NZWZeBITX4uIW6VC
VZjI7Q14xmVgwGRaqS7ZqeNg9QQzwbnfG6yiZIPdjMqM/H8fZwwVfbeoVLAVfcHC
4po6MB7630q/QlY+WzA3MQKxJ+fogyBee7RZewOoo1LkVgALZ1gsiq0a2rwLinbj
sbjxosuTi/3tW3PnJiTeEVdgVCefdIw5Lcgj4zQ81hEAyK26X9eGbR8tUMOG0OOn
5aczhzxAlfwcrbzbYA8FGWZSc4Xg0gkyxSMkMb88ediEbDADVHNXZ+eckF9Fnx0l
B6jxfJhvlIvR3Mq81Dmz/fMZvt36JoBqAzR+yX+jsZtFOkwbhBhEKRaebAZWLk9R
RPxMI4nDTP689xEFHfO9ZlwKWZjDB9eW6448+vZeBOWOuKMPDx3F7QvBKD/Z5hly
F3MmRfruyUtd5RwXL6NpUjEIYgdRmvRtH4aGjvjwJexTwQaD5BzxvItjffPnFD/a
fjTttGW+/f3vUFtsz64QkNtLIlh6kM/9B2i/6A1ozddHpAKaa8GErNbsRQ5TT0eI
5JTbRND16TnFaWW6+ByPEPdQjvlu+8QBlI7kA1OPNrGnVHTIZctIEHEVFB6SYaAo
8RaCqb35OmbWd3sjaPAP47ambz34q+JJNVFR+H/vKO9EXj/LyDXRGgUYTbUfEahk
rcBW2XfgVO2RjUqc4vuQjoxfgDuHoKOarOwQn1peL/tV/E1fwzoE8bZOPO1bdcaE
YcKf89LEBR+ebsMMSNB3HrWggRSHna9T3JyvTS/HFI2X/xHn7GKGiqAVBdF/6OJe
bcUlPd5gTdI/Bv+GduVD1BGBOu7OveB8GwkYm84ouYiSdsQQ86qRrsOH37LBiWMw
JXzd380P9J2nW/uwhMPvcpFI7Ul/uTnqIO+j7zQPEYiXSj1zjQ1HLVLfmj8S3HLK
jLzs4JkGGOvf+sPVYS89fSvUQm5p3XgYNKQswppiNX0ZDqIT/0Bhmyh+EbE581EM
ICfrEGOFy7bZLOrisQCRmhi3Ut7vaVP79LEmw9DnQV6R/15DMYY3CsynOvpULOvu
FEqQrUKAAG1foq28S34P2UEDBZV2OyIVxi2AigqLwOMbzxTFs652GwNrSJ9bePb+
q3XBW0d6kQUcTR1/o4ZoUoDMDK3qI0Rn1WKB5rhxiidQZHE5bkMKi6VDJ3mk2+Hb
80XIDG4VdUMvVOi8XuygxAReUJKHZuyGXE6gBY0VHy/VzNViDaDZqb72mpZZQpjF
nx6q2tBKJwaPEf/06C0cbmttjx2daOGJMtnezUEnde90bWctWvbVcWtKzlXaaKsz
RQsJ1XAfm9rPYIycIZTOl3eNs0XwmKP85IBQPJY8TpmyaskzGbVeD1xFpwVc8mth
zRZ4oKWcwgw3FXkAgP39oIhc9OutLSlf3zkBXkqU26lNTkdUzPisF57FmntDOM2q
o6Xa/vkfNz3Vgas1lsxvjKd+MDUL3YhidmmMAZ81KZ6UAjuLT5RZzp8pW2w10jEQ
+QHwnXexhQWEsZIlpXKM09FPJ1NIK5034bI6zs8/fChaypGXA4Dh023It1tTWCU+
ePvzFwQq61G7wgvvga4c9YHa2UB4iMr0IUNGjBFIrdyKprmWjkRPhm+SngXe3Iaf
wDIBgcmR/7ymHLkXmAqOK4z2YleG/HYfoIcYsnZIjjyzdJAncj8Sf2OTU6f9TF4x
PA4ipaqqB3aRgKhkvq2Hmss4xCaa17AaB2lDR3MZB6X5D4gZ8FRR+ANk4vRK8bN/
wj3F+4vjSj6Ep5E2x6264MlvFURF+MyR2iqMBizNvDTqfHzvxUOADo9Z8WKzZXpC
TPrhg2XyhcbnGAMNQwj9u4D3sF4rJyzqnNm8N+Pb3mRCYrkBH783/u/6yozfg/rF
x1oSvl4vXBez4kZvRMBteMEr879RXnjTZ+CduI5gnXpz9zp+LxHURpYaaGb4vNOC
ZmNvpdI/67Ay4hc0MRv8g5afltmiuyliF1yN76d9ilFJvrV8pQHOtI2BNdFcDvuT
l5dIbB9Gh8OY0jqDF1nMOEtcsYMUeXUkOyRPK0hMxUSkW7MoLhx8o1OeMJ6Awgcd
QPsOBhGVwTO+gln71GveeYRtwSkqAkHj/L7lYISP+kVOY4eyMM7kIN1y+tGFU4An
TUMbAX1JPfP3SeTVuI999VhLBNmDBV3lIW+/SQhjQuJSnwHH8NIE9g7bW0RufmVt
AXnL905d+33cVI6sLOvvZMpBqSJMALV3WhjEChtKTBVAMqTJjQjmCbmeyHmgQ2NB
EVLziqLV+TRkFbUTFoqMYgvcTRyO964xBKdXcxsO7Kk58p61W9EI8zRWTb/tzqY/
CejKcxjuP+VFLRTeVcEPNeY+X7mDu8+jVv0kgI0jhFhRA4CBVOjgrOipCiqqtR7e
eyQzg7JPfMGTCQR9wbADzcaQLP8hc62Myx6GUuqJTDTA3Bweuja5HE0iLU+qsl+x
MhRoFwCemlptMs2UpUoMt6rSsSczgCMTwyAf08jwG84/biaEDTSc3zRnmGOqJgOZ
9jlm70CiM7S1fiTeD/C+uQwF20+a7EsVO4qBiUwjibFSRIzzchyB4NFV8LS81b7q
IjkEhjPWJxdy7jEW1JkLVCIHVGhu7qrp+rczxm5PXSfztkXfna++hx52CwFCgrVt
zdlqfEEGZbuYXVY7BE/lZJY/Q38I9tSJWAwDw8rW0Lx5+9mISX/MzPqfulZ7rery
G3sd76+rQSSEeuLPJA+xrnbLSBG1pFvqgWyeMMsBH5HAut0C1YoCCzM9fC6cdFc7
PnuQEWB/fkBxE+xowUBlzGiojYLTSJMDIxPeEVYMMaTSGyON14rjv8Z0rwvt8soA
jiaWwdx+hCJR4aK2piSuyoEBjsxZ7ZoEuue/NnJDxUHYNIwrjCdmopHLZo7zfWVx
QkVMJbUfckW9eRuUdiccOOYEtdBfrZ+fiWZ0AvgpwoCuWtsW+Y3/NdeFAwoRbJU4
CiiI6E0cCwiKXqkWTyUGCW4DhSwcDC+7ie3lDxCxb3WqnkBzE03aWh2x3YEl+8S+
ZL1wVewU9nDm/OWZj2NTvd0p6nT0EWTCdfcs3+GOoFkockwkZHDT9gm9YDpirJYo
C1Ss9h9vJ7WYs3Nvokf8tJuld71mBdWHy6ylsMYgQ6+qN/Kkb8GiKdglxu/jGIOn
e3CQjYM+Ch+tixwGVqv+bqM4PdfMlGWRufxwm+t/xLV5Nv+ZcWLgfDQIO+lJByMt
c556nAikhVSB7Yj+rbue4dXjk9qJrOAmac56PYWHkLvSYZmr8jtc1bJWST25IR1f
vkP1OCzbf3D7yJA+BvIrNMItCqH0q3tovw5gLVoXZEC5M/CLQVZsCUf+DasrtVxa
Z3PLlxep4HU0BysI7FbRl/uTkOukHKbgZ50NbMKQE8fuWbFvn2tPfkmRoLWaHxja
i23yQ4HRhH4Z+WFeYZDHCNTFwgT4Lcj2X+kFhxcPQX/L+f1hVlY9tqnCfhmbeiE5
n8AemYao5VV2eeBux4cAMesVISVIDD6Nx1ayjdYNVCf0E6EUbC1cdKplxJXCf5Sp
KxoTprsmJrKUuqszWrPU5+LKBQNXorW41/FuM1f/jTMR7HdCxHO0OO4lVwL33icc
9+x7cRTSHeDJQBDflb0Ms7970AxGzoGFtWNbuag1+Hz0Lu1SPdqVDhwIhKIvoTs2
M7AWFuZWHul1BUbKCYCV5qXC5ehzyV5Myw0xIM6UyRURFtVJCW5npA3vbJAUNLJg
nLWZmuE8yYl0dHO4rmGR/KXiG+4KdF5ttPcU+b5vzE6T3SZToeCwsD3s100W/R+G
JxYi7zW085y4g+KOb4FVh+gSNU1G5XJAsmiBmc3wSs9q8l/zJ/TUX5OeMKJYCRnZ
Dyf9KMRd18s54UsqCkmehTNFxjYuR/kilBuF0uIAwAZ2BEKt7Fs5nt738JtZaczp
z63gOq5YE1P3R+oyGPtUJExwgtYjFaFfAFPedpckA4Wg+j46sBTlNhizg1R9rxFJ
nE5iSiigTgkD8cH80GCkxcbTp/SBZbihEBax/XRAfHFW+6FruxDXrRMKvuohwL0M
XGtVrKAfPaxqXEGpkhadOtJJ6gY5n/pJke28nKYhlcxZ3pgpWhFXO/f9anW7q/Od
sZTKnVUQQxKgDerZHKgtdmi7wyiKjreKiDrS7yQHnVGbjsaUrxGYt2TPoDFoyp+8
F5NSOE1XIxRdwLEqZ696XmiyeT3cYWnXMgxeuY1u5diJDPDajnNsd+ej4Y3eYXoe
e13Gfbut+e66egMKsXjNun8CqzYclV2MqO+D3j3tQB70RLKa2psP6LNaE8TMGhi5
JpgBT1f+tZCedGZ1MTcfFv23ngK2zMAKP0Uj8jZD6/3phZPJgMIKjDdnN5uovnru
NjLSaTlzhN6f4pMKmOLOPjt+zuERPNQ2Psw30XtjTsNMUP0A1sPk4ZgmmSB/sG3t
eKNY8MO+Rpesk8fTHBOqkTpodDlNo5dybPLjC7u3XYr9zQuYIQtag/4RlUyesaso
hXY+qaSruKG7gRiy+8b7u5JhBHpXf3Lbt02dBlXCZxKIQmdTbS25tqOMdYoJp5CE
ZjAzYlrk7US65NOY/Q+NimyS3M7srzW4ZpbEIccSf/kic/+ODM82VKUS49DDkmS8
AUVvu0GtAxM6WhZcFJ44TAT3NHCjNOBfbbMDI4AKcgXsXq54fElZGgbTLSYAgLJB
LjezIKMfnBaMXUfauFfUs1LAZAX6BjMxxh7j4eq5cD/oRP/jBS3y1BageOEZgMIU
Ba3X0pKS3XhxhKEpXrlxCtdQ4K/pyX9uM0Om2peCBExAWwEYAzcYUPviShrdPRec
jLD0J5ALE4ga9NbAqBY3IZi/8zXX2W+qS9jY6mLJPvCJRL5Oaq+PdloqMYdoecZ5
pCMGtW3YLvgR/bt/V6dNm8rUeGB0BGKj6ljx3RhVOgvpA70lgxR4BJsTPxrYl2rI
WcqqPLhq5XMjqIIyBGF3dmUXAHLF0YiuGElv3C+NgVfXbn56/Jd5IyIjkNiuLU1T
X85tXGWAn73ENHxWQe9fR0ty0pG4ePparcqLZi5z5+5VF8WTp+UUj0pDaY3A6YV5
w4LjH7ZUwB5p0OdoaW1xNlDWNvSFFjNgryhvkovm7XXy0c6V0c65Yv2qxwwBJQYV
g7iiNqM5NuRVD1c5ShTY6rJIzNxT3BnXnKQmgaElyx5QsluHSj3S9NBJk7L0S13B
vsqRgd7gZK/d35DF5G/ImPDaaAi1zkiI9CWiSc3DAIKjbcD4QGBBvhXvi5pqsOJ5
D/P+ccslsiXwv/IdlzMsAQfaGd70gWoDN1VNis7Y8BLmhyZtoCcsVLQe8SGLjpDl
Wnsxe87CWDO/n66MT6ciNRy4OtpPLsXBrJuSmHQpN2RrwVizk6UuafVOVWvqCEES
8pmPHVtoDqS1mofjV7P9XBTU4MlKugWHUQ8cNkg9cwGDV7Oy+S33CpnoKSDc9EMk
uWdnmoKtmVs0gHCcUJFhCsgJ2m6vb5V13pWcFFG3O8gSat+zH45wKGrmsDpQD7WE
75g3Jzxqpo7FZJd2ILokz/LePp2r/HLwiRO3kraqaH1vPJpbTwIacZb+EScph8aT
muDNKywZLVPHCoz6Fx8F8jslL8op3JxYyBa1o9zwc4jBfqXaGmsRnfXUeLCpaVRf
JwCdmjND9LNqjSlwqGs071xO20fIWXEj8pkpHeCZBk9EQ4kfn5CHgV8FRWVnU6ma
Qoye2lyfau8AyfRSR74p088ap3Nuf5iL9Qpmf2xniR9kJjURYTE7frXUtuSmxV0P
XRz/dig0JkUSXQC/ZDA8tVz5N1iw3zidhFHVQ55vTb7kkpZEZPQWUCgFGr8yTZy6
noFpF3KUry04mqyZO5kvNJw4vnUPpPpdQuytGQ2cOID8PmgXjeVuG031bUSDTV5C
JB6DTuqzDLWr2ODYYeCTXMKiXB7Le+U/igR2jWXtOqXH4YgMcFZCw+scicLoGplB
EI4L4vK5Sk9ohybitCnUT/sdUiK5+yp1nX10Vcn7p4lCv13VyIZdUsNSljEzdUQG
RLFYAMn7Zat2A6tZiWYN4esTKd2gJNfFePa+326IojrQlSAYh6slUdmp3fvw6QNT
BCQdBiJYc50Ra3eh1ppF1ZTSA60rJpbwgNd7sRU90az6gq2gcCnlKAPtXYOayeXx
2+tqiij2UU6fci1anwzptZi4nBEJtLbFwfKVAmHj1UojuSHArhRuQrj/ayxmmbVI
3uy32NMrp+T1poeN3hZrXEvmg0eZWGJY5OzJ+DoqXgewHa36D5w8lZzu4bRGQ1gy
O4ty1C9u2HMRI5z4DmzL9gdU4c0TZRJXjloWZF1+6bEtbSz6dpFRwH3od8UCL+V4
0V6gBdFQZ4WmZ8FsnwR0tYTf/M0PhZ3NEnTJAA+r9EZIvHUxNpb3mlpHtRFoL7CT
uH7dvVn/TLO5W4y18ZGUEM3IIRcwMdxUEKYe62SS6xle+65Hjc9JEiV5ZPQuLjoq
2lEZ9vpN9HRD+XVHaOG3TubVALbgn2QkOJDK/xYJQco4NhWBG3Aj/ofnWnXYdVMX
qVlduGa/Oi1k9ybbs8faoYldwmGI5ByNwnC0V4ADolV+S5DpWe+MFyVqs3UIV8Rb
9uqBPVdStogjMOE1qoZNWmTor4O2zLv/c0R4XjGDZmcuqCJGPZBzDGyEJEyBKh/2
Kzn0kEW3zoXfXI4zWczNDpNDtbMGByXt1Zr3+97a6r1s5lpoJEv7OCCnT2pmgmbp
VElHTLVqyZ1cRuKq17k3F5VK+1Jf+QlgOH0pxqmvY1jpkCvsdxy4OEpyN8/rpFdC
YHQxvXxWDtDfZGf0GQDGzSw4xf/az/eItovHKpHZMWgfnTB30YJynJoO5chkIWym
QbnzdKr0kGC0o+yWHKz3nc1yjxXr8SSlJ8MsoLEeU7Z4udrrNOEz3bN/hlwfkztA
ro7/ryOP3+W9NXeuXOfkdalOolE2fFZJCIdZdiaZ17iEghjT+LnTT6TTpXtyciT0
vLQOURrnofTxO+rAKCINHN8n18h5cc8JDgNFYA3jzKrfowu6SfgujZ82ifWR42Na
WYA+Q+YvqSeFo1TFQ5dIe3HMuRm4ZOOw5fDwHLhymuu09W2qN76wN1efXnz665EC
L3V2C5rQanVG0XeTy17rmPlBDv2GtE0PCjRfMjw5pt4809PTrVgBeOBBsPx272D2
1EpnFCYEs13HlGhi2wMjGWAAQUSVAiBtkQ3eHuBAOU29g/rOJ1O2jmJ/R60CifwU
OCZ9bgF3aFxGuQndzAyPo7XAFXdNSl7+ERSjGELJMgNQBrQZmhEMawj/bdgRVNDH
Oli2wy/FeLNZ6xtTruwUpN7D+8izazBiCIzyn3+9EzlJxfKZf1uvRHvqvirEY8T6
2H+1zdF34awWFjSjXiSgKhPgGAHY3+IiKob/PGRp0Lncm2XS94w5Fx1jBdV35UZx
UxRqksgorgyTRFH83BJWWx6PPzA08G/NGbL880Z1ZgymQqq4tPhcdhXJAiZ/+4Fq
acTtpneN/95E2Ji8ZGhpqZcZ+i75M14iqE8taNc+G0P6aikXtVJfrv6QVPvKvXkR
04aMLVyPwNtecjCYjF+UiL4waHlm69gkO5AQzL0kGzXHTdrhFy1IZIBCfF2dR0R3
pvsECeJZuFOB5MItJfUubPZr1V33nRfVFyV5BaFmDCQVb4RqH9EAnWqyPnUjA5Kv
KIaP2KN5uo6MhJhJBka+3Yr+cM8b08/XbkZYVxkoa2bcH8LRmWWlVMlBkkr08LV5
xjxO9E5vIjvh/F5Te0utWrK4uYYEaKv8YlN5E4LHfFvd2ktzprhqew+fccDvl3Jr
tqce9QASrawttpbkYaQDt/0yjWbvk21MOpOGDOUKBvdAzSBqCuZCZSqUukic3Ky7
c6zJAGxY88hjAkZWPkQRoyVkzLVix29dMQQrsqHsPJo9F7+/IzNY7okkcj5UBklP
vbkP9sstQz7dhEvIjAGjQuYplLP8oc8xdF+8ntFAU4gbaVJ7ulqoSjsfnVyLa3jM
kDelL84wTv1VbBaSQAxkZuDDVx0jISX8zari4dXxTc91UZpmoyjaSyhyPbjaD9nq
I5gpcMRYg0YoXIcbsAS5445EHoDF+ozyXFuTGkELeOm8l9BLcvdz+fC9ZeoGu3iW
tycbaOv/okhdAAEVIQ3fqYOOCuv/4f50E8x7W/tnQZ86Y8uX6eysbQ7zUOMc4U5p
VEwG7UH6fZCLiN5MwnEoBxXVC0rGnP3nmOsI4Ub9K3qlpiiuCWOm1gncxeUCmC4o
Awl+APwbphuz2dBXQGR5FCFkQt+fzk8rGwb77kVG3BorcY/aLBFcjTTy8bhrE2W8
XRjw2VrsK8/Gqv797YUo/mDdKY7ZHYNWbtuuxWWJaQlSWiNDHAkMiD7/Fid0uAbx
vVT87S3vqbZtupR6WflIFwP316cPQiGKMrfzjEhtQcAmNFjS0LFM9YS1Zg7fdRB7
kTWJDDNleBX1UZ8iElWv+qzOpZFh1JUVvnc8VXIJDxnzUH+2pVBWNAQBzLF9yVP2
VSATmj7WagSS+2zZX2vop9E6SjxlrOasdcd1jIh/xJu6tpuMLAXpyxNaQb+uB4Ex
0KCCccvx1eZivefHj9Xc/npj3UhxslP+5BWIWvRtLqHIBoXYXl8I9OOYrN8xh5JP
8Up81/hEKTFSDd1xOpW2F93QtmvXn/Jhg66FztYHV1Fib7omvTydrIhN/rcxK8n6
9xS5l8oExTKZJqJ/N5KJvu5uuRq1LhhrkmgcZqD6tlSODC8G56Q347QNRqPgg7Su
Wd4OV5LHgFyWk01kxV5DXxXPXgRp2WmC06/jBFg1d5Msoxsr1UhyfMnO+yLGv4gf
M/OlheMgfUkcSU2v9a7oxhJ7xEgWSd+U4Qk/S0f0IdzYYTBWMK/kBuHhfiaBg41Z
Yp0czHYTxcNBLPzQpuXj7gnhLD7ChasgKmuqcSb1J7RhJlGqF7Nu8rAAfMXgoQH1
xoXIMFKfdtiK2Wc3xvZhAPbVS93eidr2skGswqTg2aS7olLMMl3bfXHM1LOL7QSG
Qhun+81zYGSonNbSXf+XVSRGcdHMzhWDIRw4PPZzV6YD37M8ERFfysHoS9SWNGVt
tZMQ+O4D+Agrp9JmZgiN00VlIgYStb3PBJOzmM35xn4tIdEy19G2Qoogbn+FV0nR
QaR24d/jU0BlcKI6k+QO/v7EgGIjDDeX1H8f7xUnwEZYNG4FWCcjrI1CCz95sczx
J79DPaBnt3GsmryuYRjkkfYW8sriVGHbnquXNAzuITNK5niQLXUn8Z3pAOyoyM0/
hHDB9nDoQc/Hm5WllmBSksPm1QQXx4R95N95oRvGgKH/4MtX71aPJ04KICVjEoiE
xlvu7Z1qReAI5+Wg5AeBdy7LonL8m1HKpGH+DOdZDHV7bXrYhnHj/S1mM++o7VLa
mmRJe9OUfUvUxly+zFS4dTV3cljYSL6M9/1gAxoXWutpJbmPzr6cbRfd6hoXqItd
k2WZrOs1HqpTpkQWSdciMw1BZAMx8++5v8BQfHTBQsab4CiOffwYsHqca1lbjC0d
TnhM8DtGuILm7yjlbnt/gNknJNdNnnujb+Nnjz7UEelE6iZc8GQAHobIE0Kt9eht
6GNa7bgc32zSDxomUtvZPTJ439xvA9QRH82XRY1yq7ZGETA1yLq4EMwDgMiqpldY
6nwMPvoUsI1aR2SN+SN/5zj/1jQUiSqXFSicd4kxrNcvbtYQTIQS8fDfXXcbS0+A
hr7mUHCc3qdAiaYfdkFVSZCrV4Q9VP8iMGHNc3wlT89VlasT0Hus/OC+51X+rLKh
kPyZ9OlqIzzU/+EdCnsiVwdb+1poWH9ExGbf1rribD+DMnkoHgdixPQQekxArs0x
KlRoPV6bFaz7dYQ7RO47lhPcwpQpXF8SewI5OqamYxCpoRHA5Qwee6KJp9b58tJ8
b92qayBQNmSqo8Lf0OTvVzvp8ZAYgcX5F+SfQhT3nNpw1f8A0ACme82rpGC0bek6
MOejZriociwe+TK9mlyr9jOrcjF1l5J4KQI2GdI2n+DO+KLQJFx2cK/IO/2zNwOU
wbwYCDBSG4lA+not2feaW0AN8J6atouTn/MBmIgNGIXk2Dk3LzfoC+5ZIzVoPCl5
/X5mjppQsCgtrdtAEu182MZ3SxUefd/GQo1YRAMOHwcoZQpiHeVF3oZ/QRwnuCCJ
CsEXshH/enm7YhJ8AOS4X2aS7HiIG0Y2UYGjWvQVAiZo6nK02dMtNK+vSpHEJFsH
yOptcOMO8vIv5+ZejveWaxGZxjYPBpy5V5mdD3+p8amLBR1kMci+xS0X+Di+bczk
alU1JPdw4x0j6PLKpKPHUMRrp/k31wsKg2900zeq/xDcLhBM0vJTn/0LqzYAL0Pf
1UzHGn1CzI+5P/g6I1I96ihy77SJErZTzoja0PD+cgaI5KhBHbhf7+NSNpxRnOXY
SANM/Tt7ZOB4nrhyGLx/bbw5YvXURgoJ6QWEsrBzDqICbFd/4wQwDI5mnmb4Gsko
/d7qVdc6is4Z6hD99+6VQOdSdi6rz7uXSkHd1OSgJ9mv9Hnh4k+TN3qtTbHJkCZq
AZRB0ST6C/3eEWf2Y4rAdBmXY6kIsJYrNwr4ZTEYAOENkIiuQDHSfYKlgtsKsY5f
bOSxPn1LsMomC7JXz0LOqflRjq3gsl40PMVFzFqDnpjqAcFrmZ7u5cBXOVjoyZFF
opq6oV0T/cTukc6oMtY/K5b3gWJe9BFc9MkbCUXwKSOmQmVfisPVpVfWYA1zZzYh
IMR/T4iwRbwnrWip2ddFOWhlbId7hQbiZB3wi+3VEIfXibX8k8Ti2+o6orqugdx0
AznkF+v16zIz0mCPA1Bq4hV8sw7RQk84YrAcFnksdaYI2v7q0BSOqdZ9J5xkwNSp
Ene9UCXUyldaC+qf2xDxW2g7uyeGRhfnEgRPLzjrV521FDR2Rhw67KrJmq/4Z+ER
ymgY5PlFEAY3yD2j5L9ZTVCJTFkMyMn2nVelqfLhdp84okiGm5PwHJTLJWp5CFl1
k8/T4a61OMTshJeatURGqXr3ig3J2KehOOakZKFFjskeI8yg/6bfv2pkas6PN3GR
SxNMjTm3wr0BP1EmOFL4gm13WnG5mis7BPVHyy56pgC2bfkg1Rd98XAD89MMWVea
aDK4s6nRcqIVoRcdXg/HdM9mTt+HDbwOmywxlyhDn50MoWpHfpf7hqStEL4DtcvL
9GW1AdpPj4j+4x26ZpUfoGm9EcUAxKfyWho9/n3a7NB3WlSKwM6+JJ7uo6dwYeln
BX0cyZqx+i+SxkWJT1QpEb1EzSO4co4pn9BIv3A96yqPd4B9yhVzG3p+miZWLX3K
7qHWN37ZfLQQjI0yK59laDOoohDZbf2zMoY3c6cXsPl/Vr32RgWfITN+7iBpR5/W
cJHknnKQxgQdePYMia00Pydjm38ab/lNlVaJbdDygWULt7ArDQrDIRa+T5e/IufX
1sSSjwoySxRDNs+1n3YbHujjABWDxKxKdZ3A+ha+tXaRgyxeIUQw1jEjwT808z5i
HC1q/Hz8MFQaon0F0bOBbVYCN4Adw4ZdpqRp03oGF8CNOPXRqRkoEO58Cr1txoUr
qbRhQJmVG2CSIYy1nD5RM8ebgMll57zXESds5VTWLj38LiQpIKWjMfjMpQ1GyTjX
6twEKPZ8FKbLuAVpVfzaR8Mm4mBQdMWL1hri+E5/ckUNV2UndAIC055w6GOOLi18
rdr6yFvXyB9e8G0DvYp9UPUP/YOFl3jXPUbXfvU2abi3Re6quLYN89qbP3R3Fntu
ruicXabdQyju8tFOcNSO/LTHlTXIEPAUzFH6Z4ZICnRffLnWcXtyvUYrXCAk0ZBi
caRmwvhBUXP1+GYbRTLllmfBfOUM0sIDQ10iNAbh2kLe5HX3Cbn+UHgGKIPcvxGM
Qb+hbV28shqp4LEaTp5BT2sZQWCDtn9nnNeUF036xZ64MVNSfVTnVz36hqjAZG8K
E/43rhPFPDDYjPuZd7XUgC7qubwEbLq4h331fayD13ImZEkL2IFG1xn5pLJrdliQ
UZGlxpHJj7Yu5sPDZicgP95JfsO9GQkMrew52cVPW9bOHRUG+DxoxRfi56lD6ryK
EJKw6me3XTbVx2ZJs22KCQ6uOWX8NQsRIvzixrg4ilZN14wmwM8eP1X0FEt+mnp+
12Y2NEX0r/w2x97cMGAm+DwC5FcHs7DfEnrYUHyfyaMmMhbImawDN/ofkhEjQQW5
cwjVffwg7X7edsEoUaknqqnTnFz3yRineojAgN4a8whh4i6B60tR34kqvYGTqFsO
wSH8FodA1kNrDabWpSL4OtireR0/LVk6CUJlYko5X1xr2MPzPRSYXOoVU7vgpu7w
DPA13ZUwHo/qQQQz7ndS9QaBdyud+DCZU6D2WvajstvW11Xb6GwOKV1/7eZEN1dT
Bkbn7xw2Ww5BqqnPXeNs8HRQ1I5PDW+G1Skkrvw73dERFl2L1alcTn3hfDknZK9p
c9XhrvGrvj2CxxZlKpGHIT0o2tdsiaB9FKmCVE6QZQL0O93G08o6yqhe9ks2FtHq
WYIknvL0kx1WGDU2WYpJavLuZ2MAEH4Jc+OWQXdbtsIPpuPN+hamGe90DNyY+Va+
doBplpktVQ+z68nFmIWuC707zDu3t2ExTaBm5W6xy1uamfxqG3SSPj+fMoFZcIfQ
B+qA+WcAvSrxX4Q5J9LZdtEdxR5cFjQQXf9n1JZSombnz/rpFGH7Y3BKf3jTEVwD
Fbbvo3Nc4XPIA8DLpGMhmF9E1l5HGuBpsuU/PJouA7VAg+JlN7hRHWAKB1aanKts
mzxeZGUWiR3jbqNWBIbvhgWtLrwADonUr0S9oWhwQpJOpcz6zpbxEHjrUGVJoh72
QBuVOS2TOx3Vha9TDaLdzl08L04ChHdtKLano0cBOBYUTM66a9L4l7DzKot6FykN
PxpPErX/F/CEl5Jld9HxCIUpwrfcFHmIzztLCbMo/7ft4PjmMJZR0DVeepGF039R
FX3edlsZxOw1cN6iPLO4E0NL9XoCb/lrqfzLRLYsznPAwPioeCVJ1mBm6TOL4XN/
dw/9tN4Se19/5nnBlvUiTVGiqkkOcClrUUfbrU2tQnTJgagnQE5TOb0JbG4YvPn8
e9jwaBQFoYIyrgKLHZm/QM2jYxgj4zYpdYJB3lUTk5I2BIUn1AB3iYKMpIi3Uea0
UQNYg2pa7TnQlwOsaTOI78RTjzAo+MTNCyYpUoq0YYnJ2D09wzB22ckiZTy3fuNM
KsQmI2r40H64UKPozJpXaQj5sGNKLLPhONA1F68vaHEQIShXjNxjRcNrlEIQ9Shl
34/r9FxaY06vhXm8Pma6DfvSamVHwa1DbEWpVCpw9Cmb56l7lJwgqcRLRzS5rD0V
pHRQ/D836tecHontvUYS9Bw/qcmcFQCSelldBBfZORRHA+Ns3dNrrm03lGEBJ3h+
OqLfi8rW8+p/eTIqkfubYPwLhYxn3ZrzUbQcUnFZw9U7AnhiJhjAhDKw5w9vU63t
eufb+6BeK+o/Bsm4f150lvkF+g9G3N5yaSpNsbgQhEilrNtFzJrKI1PzWcWeDEQ6
JYqO2PBhOmfmoGy4qRWws6HiZHTBKlpoK4EiiHE72NRK/mScSigYywgnq5a7wzfx
C68yMdYicQUKNcXuEAIabK84OX6wzQsYjTzDSNjFh2huBjGRbEiMmsRxy+mCtyai
K4vGGmde+N46hTuKwCf2dBerSzeepjWBiRJZHYOtqb92ySfJzQ1r5cIXk03XDgkO
6d5O90Evtw9xkBe6k7CC+ec7+CdJ0IJXHbO2MUDOLzoWTIn9u5KF/V785jArilol
weS4/kEl229RLrtNkZIeOoi6f2MgjJfZ6WbjvX/n4+NEwNLUvpKB0fba+oD3GhVL
m2PeqEM66+jjllKguRKpkd1KCIVSzWZE7xjfvk3dKaNuKXtklbuLU+8SEKriva+4
tAOwgBV6XwW1YIHDl6ggqtpIn87IphJ+GHKjdNbODK5RLUlFLbNaT+96PHVnwL/f
QacJTcOMf7qRjyP4OU/mM5TVyG4jmQ1JyWgQELHiE+ChDhCEO8QgvnHv92+3/Pne
7lgz4GHSNBB9vzYPFdssyKy5JEgHDMZJKyMSotPKAGVtGU6RzR3Yp4ImdSvbGxVU
Y5hFuyoIJydEWazZUBdhQTDhSWJUg1sZxkASZzU5XH4C8axssT6Gpf1LQAF+YCX1
5SlApdUo5+QzWnOCMlWz3ZZwZlZgJBQl3+AJ5mHzZmRalsCWXox3wfH6mcz8Aho4
IX0XVMoslmOsv3y/zayFxA==
`pragma protect end_protected
