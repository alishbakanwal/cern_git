// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:05:39 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
MULioKz2PdJbyCcNZNqGTNOjaDyOfEUrzj9bMG10L6iD+m/MrKS0c7ztdl20BzGh
UydrAEvshIDSV8IFDHR9Z0MR0bRuM1siFkvaVbA7tHiaBRGP6eq3u6PJyOPimudm
Ov9eeRH62awXETaGHz/c2mOn1/TL4/ydLUn4Z70UkGI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 16640)
BzSiv1U0XAPva8+diio66jqdYRoraOCMzHjTK07IvFwKmp7UA9fdmxw7MTWH+mz3
XCw+I5VHtrlTvt9YFzti5N++xHfEKzAIoAzZFtTWIxr/Tua8VeNBIdSwgbyZtyYF
A8dEw8p2I5lrMZ1m8TafoJ0D0w2PJb0LS1xLctgIrpzRhVwjD646KtYqRFDhONbG
vpQilI5+hvBVapFEkBldujlNnLeNbuYEW03H6TLeXy+6hvP/Wir5MUrv+efLeNZw
6m90NFbMyob5Y80eYKIs4uGKRef2gIxJDCUAFU/FRHDJtErls2z0eCczO/X4YwT4
YZchupqt499QA1xaGcdgpk86MXvi2zsVGsHu1eIYQr13T00MsFnmhbG8bbfrmtXU
LtE0aQyWx5e0FrZU0Vsbs8lp0KMmvym05NgvdkORuoFoBA4P+iK1L4e0CjmCUYkQ
HR3M2xS47d2zDXCffdoL3bANWw4rs/evf7BvJhJQJfw3bZZxmnYyy0+zTdDJzY+s
8USh/2EVjhu6gw0qE1T70K6ZR1071vCPDtIygf8EkXceXiW6vdP92LrLv7/UAsFC
IWHiRxrdpdRmq4kIVDILcvbomasVqcqkjNP4vFHpUQPxtuot7PZGotPFtYLK9wsd
5d7twZUP9ej7zkA4Blzk9INpdEnkLkJUnCwuacN+/mhACOxLLY1YLb8XxxVBUlQw
9Qeel6BbQ8uy2/rig16uzNvUCyasT73nwKPFlvc/QfeGe2gH2BM3+GEhrTOT4In5
nJkNnhKKTNWGbC0RH6sWoJzfsK3GZ5awJgqCSZNhzub7UjnyhqMjmI8dJcCLgAD4
sRkTvnAQwOLI6zd19AIbwAXZX/D+tNbq5o+hmIzA3UlsnpOnhIrcV7dNj53GxSuH
9fxbIZf+4NCqMDIkto3z5cMqA95z31PWVfoItXxyNJONHRjNjNOGxTKh0CYHMcGw
1H8Ygj01GlqHp+4Uu7ImxyRYzzfE4wgGGisgNmrETpAoPwToaqrUQrCM8yJnefv2
nGMAKASdJcy4v3Je1qTjZ5RjX9uXe1behmjCXih0dLFbHx+HR/iESSNFZ7aTXGFR
LYYiA2n3gaCUAVkmWMtPz38C4Yoj47FlWdQSHWGk7RfgxwTBV8jgtHuI4rFIlAkx
MatAhrDTr8VRuXJC4g9XCYJsNhuX5/dDVV8fDoZsWIwE6rsZh9rQOMXFMMrTGdjg
8IO9e2UmPDZBU8GBaSs8SXCnc2J0ku1m7u8nbz5HTX3ncK7Pzq86HKmsODCHThM+
RoPlfpT9H/cLPQeBAsyBv9MzxoC87Kky3d8b2NGSLiYbuaJfDoCtn0WYIfSvqUug
Ee9rulDwLVAl5GaJkCrkLAnf2WyFbxZ6zSjbj5+84Tyq5I5Lc3Pq4kw5fx0zYNPI
k54vXFFEB79Frc0axKcbeKVZESSMyQLhZ77vwR86PtGwFEAZCZTW74wc/rqGjqvW
o4CU3DEwzbWMPyViQzGo/silpe3mbceBEPz/coXaoJNP9ddn+W33Pdc0l1ujYtzG
jwUpXT6Zkl1OCCwHAt80CcDp+TtxkMV0fUovtp5LpOsSxjFBTGaVrguRy/Avr4Rw
mFbciCWAHBkbyM/iMJZ7Gu4Hk0D9fX5SvH3jmLaF2AU49uJTZazagygv3uVTD02I
hgA2SwlAg989ooBrLR/GMzE7CcmEcQpd/4406f+6k2Jzd4hgrhOyF3/qEQ6N+2I/
bEZvBsaOqNly3PZOhCefXsc5Bsv175XkqedGDOjwIzSbQVIS4w7DD6g7mQkWxd5o
xMCXfbXb6U0j/IdpggaE17nYdqAEtwfEoyGYswMAWJxZMPPiUMFMrAA4KwXbb/+i
RMKZyw4hHr/3heHBr6hJTAVrc9nS2mBCZMCPy5xC6EDaxRFCgXGCCcA7L/bEAq2T
EF/1CR0LUgWknnxAsKn0wddn3guhEnjT/IsbYft9nAnNb7uiRBWhKLR7owzFsk7F
Q6onIFYlrgTv4PtFkc1NieALhm6/9mDWD96idZnaORMSvhlPzFhLuLzXk7XXXraX
gZpTjzFRUHsSP6a8KRs/QvcgH8hmaOkUA9DZXaKcxccobcToXmb3SUnLulo+0TA3
X6VG0j47u67+je2VdhQfgKdfuXeBDR0/mJEbK9dPcMHYpl3uR3JgnMZ87ScmZY6k
6sQ7Le3alW9gRLx8FCzwuLLCkA64VohPo5Qk7JS404vF5YsDszfMgAz97yHTFTMQ
lukOPJ1wHkblcLEBLC5AYKB7vKjASsGRaimS6qfbIPjqKWwo9PMYziGnNnzP1DtR
OKEd6ihIYAXkD2GvKKWgTxawLvKJtbfMHnO1k7EvngeGoH3C9GCKjTGCxV7tY68W
CiUUqX8Bn4uGxOwNR5jjUgB+O6MxO5ITWmA6sfeK6yMeC1xHNOOAITXSUEpPv21y
Z6BqcGAsdeFFiFHtAUJoniFJWbsADEn/mMHKy9UP4NA6LADgRZzWSZwwqdr0j6lu
U0h9ounZM9XoA2Ggq1gR9lpIVsfNxWdTp1Q3f0kRhklqdd8IpEDwySaw607CNAl+
8uV4gpYWEPEdTue49R1zt8Jg/6S2o+OzeF+JiACTr4Dj5ciebmj8Oa/tktO52OH3
E3Ce+e5vAu5VwIyNDgks0S/TFm40wQQt2Q1cDjNeQ/sQ0ZOrXQYekW0fPl8qNST9
ABcYHthNZK+VJb4QHGpoTsQzR9avvlW0m/MN+uMZkGJOqXD+hZSrf5nQzqYybQrK
485zQql71E3nAiMxJ7eMO2kI4Qbai9brwPIMOUSNXm5Q9N74BV9TFFdlVcJcvmsT
CnwkemzZkKXeHJ2rNWsgCHSZI2VkqpGgd8De9B+iVBlh5WX/MBWPsh+Nx4n4xkJs
yto7CvWK3N8Nx3//8LL7+qMJPTCcCwTiu+LW16MZbar7pmnoV2H5WkI0bdaiVT8r
wKoe/Zw1ZpPZJxiGMVipB/pgp93DNDx49DJ0+Kb48xXv+Gx1Tg6xr+JvI9Cax9/K
a9Z2cYHyYN85AyBZ1QVM/5M0f8L5+Ej9UWLUlg9OFCPNZkHP4RWmGwYeqmsp3KVQ
ZFcV9pz0MzJ7jiQMC6j6f9m/s5hqsrUqNjUfNL//IZMg0SBRPNlEXWCLjVwrod0Y
6dHh5cqhkzId8pe4qaIXX4T/qE2ojZf8RC5xQFMyBQQDRw63Js7FNib0pGlDrbDu
imsvR0Z8okNsqf03rfj6ctgcG2e+5Mou+c6C+1hkbqUf8mZ5IkeX7vaLuqqowQHp
STubLJEqoL8eBI3LnLr8LHi9o7ZJaWkQ8DRRgzGSzuilv8xSaPraGiQEvcRmbaRD
RZ3FG/j9K7xROGauqFRY92/o0bD47KPO4Wfk0nP8FdFHVup7gDfSQvHh9qoJ2gIV
t+XtjsK6+2XgYOq5hpUIqX8wpulW5m1hRrRWyyxsRtNHChEXHgwl92xonrOyv2CQ
PyngmGLSYc7Ydjf4FsjUs27Dsgwnb5bJgbbSvyKIe7EQVn4uJ27jx8iXA+ixdi5P
xKFNnNBLjHLrqadHbH7hrb2ZfynhLCiJJGglyCkAAJnd57nBvqOEYk9in9rY5icR
D/IznlYXR+h5PRHRGqf00X4nCUoYMXko7IQtTRVjFMWBWghoAbLSvxhSip4bJQHK
0gw9M0Knob2ZXPkh2TrJlvK6uK3xbBJ28/9Qvh8X7Z838oRPLMNArMUwWKzDqknG
jEwjJZSB2B3x9KTQgoJfwd0ZeJhDeeSARyBjaGogChASFVAM+T2O/jHUS4SrBfMf
WWFX3MpZGBOg4AK4yrk2lJdzDjr4BpVZhtQqVuu8hxZT8AxCob9aVK0rBlg0SllW
PluzI1Ocr+c0BE9fvByPcCppR7fRFyxJt2vt4UJwSJISWXC5v5PshbWqbA6cpqmm
dxGQFnifiJBhUaur3CSH+YQC7WF/UzY4xGOE6yK0S85YVeBk1L54H73uDBUh36Sz
cbeOky3u2rL8KufVYtMOK+ML2pqh5DRlf4cDY1WBgqbDV+3wGXH93oaRNLdx6cyo
eNjdskPdbiZp2JfI9P6DDK2WgGWvWvyXBmAAWVjDi/AUygHEF0PO0Vvrf3aKJXUK
HDV+PV4OIPWLYkZTg/Wiy4oXBQCabRJ5ZJt5tRpIfgwgzxXMM+617nUcNlXPHUlo
YnfQKrXOdnYscTRIoGh/LN8QsfbX+oPD0j8iPWLPW3Jwjl97s4nIjIzupVHTIexK
HqB9Q6uutqVal9Rjc11GBVGZwu6e3jZSLWLYEn5Npp42yczkefVKulOWFc9o4r7G
Uza8tp3nbrsyzy0zSFR45KA27+1c/fl5XaIVdPJL46untRE7EFimCH4xoXTsn+J9
brtY6NLqqKRnvxSK1cUEDdAwH3GmkFdB4VsaGveypgMr9GJGlRP+ZbHjSpdtGx5q
1VrsR+bK6JYDce+Ehb/lqUOURxsfpOuzIv8q2wt1U/7DIWVFzgPIQaW0b0lX9p+G
II1ZYPiaQnyI+a8QKpf5fzLxtVj9R2ZFlGlaLlTPyQYK3pK3WyikOvC+EqXhhECo
fM0nBrr2lYFVL9qM4YcsrzKe3+bUKqeKpgPCJK1tC50+Jxnw83zWZgvWilM06zR6
dcrGehhmu/N4k3vEBw/fe49YFnfeS+kvYlFOQBkvLlVSIWNcLX/kpaMncJWjrNf+
wVKrdSS2Qwwdme4IE5KxfbBfynMAan8cJkVC0kGtFMNbOdddKwMEWuyGNutqN8/S
uGNFIkh1A26JQMFL4d1HN212Qxu/8FF29nGM8hJXXCTbGnS4vXprGVwMSGD7Jyk3
HWlTLVwtCRRp287VPKAQKQEZB5KA+cJL7qOBo0YwbCLPh4qky331Z1J8WD5ob8xA
KNrOlH7DtxsYRh936Y3Z/yDE//pkQCspp32d/ULgl0N8oPnoFafk7AzdbAg6OL4N
niGvsf1bW343MW1e4/HtSmxsVEEHmzpYCOuV5PCa1QTgq29T2+ewxp+N+Z3saFLY
cVUtJGyYnpujp6sjed8NKIisF/e3/+MtLu4iYT4+jJzCnn4dkX+nqBHZzB/7nBB0
WTFWrprxZD4SQRjsi0Bxw+4Z62xMW0UZRgYWcjjaX6wGE6MiBEl9rogO8S3wvD8E
dXnaq/l5+vMa6iu3tdvL97Nx/nBG3JJVU2F10TTfJ8tXG2B6uA5/xpIcFReGm2BU
+mv2NzzIMPF2ymwkHDqEcXcot5TACszODjkNvOrCMrCLh3j1eCf1l+p43wv04T7D
TeVUDXK6yG/3hpvLEkOQMJblhC15w0WeQQPMiK3miCHnfDCCenv5xOgNIe4Qax5O
COFTGRFzkiBRE1+dGZMdj51+twfIML/R5ZLGLJDPzxTiqTdRszjVD3MPg/nX77Dl
dKaN2vBEZAEw03WHC9QzDX0RSfuoJEN4VpdummK/5/HXHwJxtvq3kpyQgdy4GMsu
21X8RMis9caKg/8wY5BbJJpAxosZY4AVgZVq670F6wgoEEDrhLVMuaGpRfoUlpdG
4lXCZLkJWSL3JizWAjqrwj/3c0SIS5OIAF7U9znQT5j60bvN4U+SmOnYaDGJQjRo
VzWIXx6ZCiY04gFoVBZ2pYd+BivY8vdZkQDrsNc7SNiN3Z+nWANsCIUbJFroQkrJ
nMl6z8qPmGN52F+Qr6+uwk20AxZR8HicBvlF77DiZ4eWOF+/x4Zw2WTEfVGMbIqe
QJlVRDFZZjxaGNa7EIs5doslbVX8hwe01CwZReTMzLAYJqEqvw7t+l2j7kMGuPCA
waIMIbZsEOFKEw0ukrDO4JmLmANpnw+telCIcKytDubYpyOIV1zIzNRNSIHv0MDt
leoqgqUWEKOpAnsYzIaLPohFCaFsN+AZbovvXlFSPC4JmwxwE4NDRxhI7bdfx3i9
FA9Tj8GNJD3gbQvlq0zfRPL8XN5plCqmQi8a7Y5SGwb27Y81QmhxzhD+pqu1jpBS
VOBR8MY2r3NHstckuLVVfTNEV993xJIyv6SxbqfBBth/hHd2/qtCMoty0fSMpshb
KgjaHdEGL61w3Aci75ZpDYEceazDZ06V8I4kcvGvxRIdlIfysC2JYvjx8xXK00oT
8lvkV6uMHJ7UiTsGLYIVp28HmMexZblhgOQTFxDjSP5GjzJsgCxd2NcgiS5FiNeC
mx7Lza7rbsjPhmdL7Njaoa+hQlS/NCI7Q/1kJ9WS+J9G5N7z0SvtKdQVmSIFtUKr
zyqw46uWB6JvZ6C9xWO2/4Dr75wjk652kk+ySttlVAgjguo52217mMFmXtjUa8cs
u8QSN3yW4VcWM8XgZad3+4wQmINcUoVTCGu4EWfgUy14kSR/ktHdZugpbnDEYNd9
LNK9Lvt0rCSxJOV80NDa7IYg2S5ArjDaKGrkuViHZn9Z9BEprHbmhqUDS7dvdYUf
0GlYC+D2qLvgvNLMk4rV/IB0CCeuTNiALZ6UBH2bpCV+uoRj8dicFzMkZU7142Bx
2p48/1td+nkC4kvtnRPWn6iS18zcO5vfQ7Cu+uEBYxT9/L+rHC/PoaH6KA4NdJC/
dpmzvhE1jBxZR/IkgSKq1YaB+hq9Zn6Jh6FHMmxU2kfTbh+tKExcGT6W5O/neU1f
xblMtroV775ZUj6iVcpsUMbYMrZxruIQ6dOboeDUo01uSfBK8Q4K2z+eoxFNCMUS
AfMRBbW+G9UiOFcIB8ORI3nzullaAg+CRcKeLM+7X6f9pzfW7Gr5umCV7LMxzXq4
bCtPvOlfk8kFbjgQkv97TIjL65KJ0C9KJjyVF/xwtav3jWbqz21TroSA3WvC41GU
DNJ2Xj0eMCgsQalU+zMqJVVwCuAJ7S4yzuSshRHcwyO75YPrnOrKUO6ZwCrU0cTk
E40sQvCFZSOs4L6vdnmyj2VBnO1i7kgX7LOgbS//Gkxbf6Rv6HPUx8iI8WrIZcSd
xjxGOsh5Od8/cxmkffupUQ8yiy41EEdh4KYIO/ebLTGpDTXtQPsZmNdlz0y5TxQM
uw+XV4lSWcInLnuYpBpFWJ/CNiqcphapn5oLA8+6Cx9a2GeUVvwSX0W90oK6BPDb
CBopd3GpnWSzi4/gnq2qNjm3u3DyDxYbAHnbqcYDqTjNoqoY1/bZvSvm5tbKMQvg
+OlGZEkk+pye6oYuvJujXHGDqBcy4jbi9LI5IqKjOebbf07vNpZv89UUa3H2LHrd
jgimrKzv7x552zTRhOa7PHaQpj20sHklHIajZcESmJmNt+oA7AuZ8IBH4V4v2gNk
/BeNF1pZUPUKqFKQH9/mf2BBzxzNZkehKxXCVnBflPTPFaKsy07XOjc+5B+pwn3u
zRLkGpeKmxkekvqbDJ9f04k6cp+FHnddCFqrJqJKzdEG9PFLZG1xeJtlA6x7qL8D
60LCO0MowoHDeR8+vuektSHyu/CXSIEiQrRB34RzmIhho9098Eqfy4xvK8eBkZ3d
GXig4wnS4RGrwbkPHn2nsYfr6BcuayT9SMrW+n2SYfbPk48rHJUsFtO7J2HCgync
BVFGP/GDIvqbwkt7mUqNWnZXKOb7Rdrl7Tjab0EvcbLCD52iksmmYUQ1+othsd8s
97wbZHJlNEuF/U6QSWWwK6Mi9+Rp+DNialGlbrngbHq0qEyLmN/Kelb63Hjxa+W0
0IWoTraJBuAawK5zr63M+wrwSKfKGKdGKx0eATCSuqYm3BLhnMB/9mlJ1zgtDS3v
vrJ7nO8HwIVprEDeXISWWh8d2XPZ0+TIzScv4etTCttTyFOr2hJELq24HbqXdgTb
EVPz/eHdZSzpzab4j2jyDJzioiLKG2WJJGWPKMiBBsWEDKf8SWU/zn7BqGRCIzMt
HneIIJ//SAMUl3XTs3I5wLJHPpc5Lbli2OlHGEy2/3+clI/btm6jg4xDz6iLOsk2
l86QfzMCDfFFul6PgfNi7CuAU79uqis4GNNoNiLg77TsmQXs+TxHeOSJ0QyC4s0z
9yFKp0Q8YV54yVaQZR9BUuhsZrBWYBcgUnAXanRW1J81UvUAC/lZOCOpQTp7Jc8/
jzqN4Wb0dx8rkup4BdHd5Rz5jueJs1WWmeKJWz2bJkaEZJJzkQcDWQmSlqQJ0S72
q6vd781PnPRzdk4SPiRCz0yPjfzKCPiOo3VC20TjAG15xUmFx2fSrdAZ122xRln2
V/OxQdqc2w4Xas0drOgQdZryd8AFLOnLAY4NIa4RvMMcC3EgspkrqrrE+9GDGoBi
VngjppFb1PkCKXflyODdq/JiAgwmVvBBeW472hORz8Wuxb2LjErVw5xz8CK2Vlkr
+WOmwswI3OR0E5/dmWiL3CkgKThHOO9MUfuVj59NLk/UQAMCgUK1RjcHnuSrVZzi
KjOJ83TYpho8Gcakk/FM5v/87VcLgA41hqMz+bxuHwyTUB+DwgCrLXd8fKoJgSuo
tJTTuIcY5qIuU/xFqor0Ktp/JiceTAy0nh+JvFb/Q72zeZFnJDijbz1xHegwxVuY
y5ZrWt7FwWvbVwPV54XLnrPSMMM68E/3MUVps8PA61QML+GhSJdQ/RKuh+8Y8pwi
8XXR+qCJnO/+zLzBF1GmuC8/5TDOJ5BJGZOh1w8meVL8bZebioKUZ4OR/S1dwYsa
Xf6N7Jgqe8V69ktRomYIL//62AnJdaX6FYLd53hga0gU23t2QL3N+xrp+EVF+P55
WUsTPKnl6oGcHqxj2jNvigSG2TT3vaywrS7SXUq8jegLKQyOcvqfQUAqbalf2HEl
iucrt3kfU06UVUxrpgjJef6DmO/5LdzqjwEmJwR8xvf8vKsOJ2FeCTjM53LwVOgw
7dTRv4HUXgfeHAaevfdW9MFfpxtF/os4SKwG/IviR14ZsIgysKKONL0izARgb8TY
eMytTVnWvb3OmPsNs+SZd9FTcYCpk/iBSTSd4TR+wYzGABizl35vBgu+gDStaciU
foGJvRv0QbfxW1L0z5Xv7lxp1qm07bfBpeTDbcPotXlKbAz/iTaBzRWvLGSu834A
DAhgVgfIHPLLBqQwS+KVs8yRjUyasI7NIgdgQYgUrk0OdHrSGO2z3RTzLRmKa8hs
mG01FxLdZ/wd9WbFMz1SLZiL8Xn5cdH5dOdR7wnMiP7jHnLp1uZW0wnbw2riTBNU
uFzDNlRBDgYOyDrPo21R9xUDL5tcHIpr55/Q2U4OYSaqtEql12+ZBYcAUmLRk+7H
mIKKUrcDF8Jw2Y+1GgcK8c5piYcfksT3x2s13RfrHJh2wYg29FmiHMzkllHXoWey
IFCq3g1q8/eYLdFnFxgsLHpQywXKR5489zX0oUCaEoVCnQ5jmO2PhEK8k2F0JVt9
wV7dP08R8Wv0FctBi3L+KjVWCq58J6U824q24xC79gNcJCw0cm1QPAnq77lMIMuM
mzH0tF/DrYNd0nQo0mB7MB1sBVopMBGKxOXV9sY/OG6eAtu5dkb//zklpfqX/TwA
bSHISwcHT1BPFltO7aVTLf8dHrmOi6Yz9CLDgPTwvuBQ8Hv6Szx9tiLl+cm3sdVP
KgyaetiV4T+WxfzbWaDRBRZ7nKxn/QiIoyfTO/JODbRgO+UQ6KREAhGiHZBWTneb
1XrjeIzsxNAi7t54+8m1JzFrirEirPzxSeRStejfHthIS5sAts1RBZmyQGRsMrj2
XdPTiWDj/7WrgSnS7qDQlil8MYnh5Q44A7XNRjPAixlQMaK3wmNt2Igef0ZrrI6s
jZnBV1IMwN1S+ltjT6ecUG0e5+KZqkNjk3JoBIdaMNRPPOeN75rzXiLXQmxJRaO7
EUwtlQ7XUKuAIihp0u8uaXYr7SFgazGfeFrkWPyFkHUbAB6bIzKDKduD1j08mqhq
qgFaWpf6MlchqEWb6q3BdDnM2cdyCtAPJmQBFezJPL4EOjZRQ+C74T48qzyuEwnK
DFamlR8MEjuxuf47XBV7Z5GW0qHZVfLI4R8rMTuZD71jtJrMykBBobTOriTnbJdg
Lb0K+8DpEFqnJi1G72iRLXhXSRjLCYaO23mmXzOWGdfQFGObA6zHSzO2Cw1CKmMh
59llm/Au5nm3jBetWuheZI23kogi6elWyoZD4kQCOT6voyMs8BKNPi6IGkw4ykU3
k8/nO7p8rcwf+m4Drt00J3LIy1yVZfkthWUSlTk3zYVaQzou3KvQfH9lr7crJt17
e7/9h/eD5e850wcZp8TMfh5E34RD+yMPNsG3ISF+SUXwpVJ9AEQatRCO60lGsAUn
NGbIs7NrF1hYz6xHN80Bfay+jhPuXb+tK5C4/FsU4nCkw2kwOR2AsNjsO3cqU/O7
3KbT3DpS1tvm2Sy0NWecpnn0ji7eIiN3dE+Mul7WAqb3yVjjrnZj64rdPhl+f/ii
GzQwMQoRrgyndehmxUg+68KGEOdS772T/naKKuUYr9qDS4pr9eP+jBawGClCu1nb
G9s3LXx0L3sweHqHCaM8oP7TWML2or4GWoGB8RyZu2nnTbDB8LPC+M6XXM7doDQo
xrCmKeMf24rDzJ1oH3bgrLqWUKXEz1jK1vt76ifi5vlOZF+Gv/in/wyCz8G+EFh3
zVBhCFwkNT/lEhhJENpJhDr8e8x/GQ9N2d1tnmQ7DYtnIKe2WZVzWc1T2Rk9DhdW
LTmAWqM5PUa5p+jTiN8Bt/cSjzjfsepzPxeS1XTayhFu7fsrLaz/uJNzCXhvyIj2
6BhNH/ywz0BdAjUJSs8/oIJVjVvR2lD8P2Q9gM/ZX4c0YPLzwpNeN39jxSDygFCO
0mrOD6XDJLP/z8Hdpw+fq2Ei7dq3xpwjLJOm2iGAibQlJayqQOqEQTDf9GeCEcB0
vRb8JdVS6/MPbPlfqzWjbPuZY5lhbN6+tgsAkywMoidLcXREd7pGWhuMtZRnPKME
zRnLISFmSj21/9/jPerPK+8Gnixkw7h1WkytIlDYhFyRqHlfKsqs/QEIZdM+eJil
X6Mm+yxO2Z5jVFRTb2/rjEw1iyaX5Ka7HCsW0mUNQEAacXFs0f8qNchAV3o6jSD8
CUxY7T4JUVMv/RVcsn5mll3v2FIQzxWz01ybymNAdiDZXMasFggdizidGbsoVzRS
chNHXiIqXGXfIWai7GgYRZJTM60us/raKrR/ckyjPKh6aoys6/YCpOAMqbo2A2bQ
2ycydn5BZg7l/DV8xSl09+B4zdfYA9V6n4z1lUWq8bwGXYGfBcMS+dwtdbesYaQA
3D8cpb0HMNtHkjzgOQqtiWChdzWwMp9DDCdD3noQf/Yr8fJFUNjsQKNpydgeQSB3
UtCnBPB0+457EOMOgELpUDNyjOtj0+EnMaBvX8ms0Cirjye6/WR0oWJvEXILrG6P
nTpb9LjePZwPjynv0FZifQKU+85rwoVMgvbvPdenOwSV/zB8502+fanOVyS1NtAf
CBEM7zpHg2Fmaw3N5q8VtbYjWpqbOW98Evbusy3WgjbCMMwQh/Hrpo6WtdrVqyqd
+sha/9EdXiYC2NWK3Tbh/FQrq9l3DST3W4We1/I29bFetJ2B4F+DOR20rB25Jfy9
YW+SjCaU6BJ5ifU+3bpBcaaoM3Y1Rog5pJiG6mjkxSfO8bTV8pgQak8vdkdbyZiQ
Q2AYVQy4Lx9vOgcwiB6TeMVcL3merUrKSX51nI7wsKS9smkxXBsPoLKsDm7Zp9xa
Ja7+dxwiA7pHp/QNh5hfJ5ubx3TB4xRpedARFad4hmkKuMJv19rwhmOMqwK4WuPx
2gnI6BSmQsUDQlDrfAYKXLLk3IYqmqxBONfkonZiARr9av1o/rp4gLRvsx0YSyWA
zc1B4K9hXsz1oNl2PqX9hkeq7wgXi+CKEJBzFui3lTAVb+vfegMfuXYcurc4F4le
Z3Ss1kcB7ZWoyZw22Km/jHL98slAFPw37bCeQMbEhsJfa4Bk2m0rf94AIASWzGKh
oAlQwZN+t1zbfaIzfVJJSzBZpFkUecgsw3KFPZKK3pPFfm9LMFJQic/jJaddZIIV
rbcrI3m4lJXtmCehsbKEjjqP1aDIJQLXJxQRYQIp6qRpIHBn1fLha4pV+ysP/ePg
Ko275uE1diQpyWHmyQx9AhVbkifqJpS52+/5hAcpj0iUb+ajvUrAZD+uDMv/S+td
oBkp1HkFj2J+QHsU1l3SqFmc73729MJEhEsh1anzOBO/e/NwUnOAPLl8ZN5iWyRS
GS0sOA87PujcF/Bsp18hRn0+FcgzxNdTapw8+TRYyxrI7Q5ApHtahG914dTAARfu
Jbo9pQ9+2CftifB6kh4mGEfwfQpOeOC+8cT4T0JXMKlaKxCbW4HOZAUG0ty4utLQ
aCVqFhIXhmH+a8KYXOM/9jOThX+EKkZlhejj2Va9nCTwZXdDJQ6gfBReAMoNblG0
pz6myBnoxiHApT+Sn82ctdbHbkcmNYmMn451ICXYMsINx6FAwroB7Iw9OtUgH8b4
3R4deUckGrigzbvk4rScqCxGvEklY9zQgYpiMBUzBDAsQpHMXrPjT0JPuFWobZKI
viIneUADYGr5FH+u6pB6HZ4CNNATlfdGesZKoeudV40Dsch9UaHx/Yqmqb+bquGB
uT3FxobQKlKq/GHKdxqvhmecl30/tWAEcm3XdtIAUfMLzxKbRf1Gnou8ufAtV0S3
JTdsZmnmqsL8z6/gFY3ptUiSZ0pKLHvaZdoD2hP4Tak+rSWU8BMIKym1+uQHVuK2
eU0Y+x9W4ZqE+GOEaajbfMTRgm/kaEY8YaxkWn8WZ4MSJZSO21HCHsZYp/VwBbW9
YK5Y2RnznRNQ6XYTLGskFZGvlSBvWUsFYi+lzgE9QmMw173jk7+mamyfZGqxVnO0
74csl6S2C4WaznNv4Uxh7lLxhbHNB1u/4hYu4WgoD9Ggvf/pKOu5UFJGEZUMqSIL
nM2KiQKQYHAtwXID9h6rGIXw+UKXuexfXAZ5sSbcmW6lwhuRl3RCVx7Na67xvFro
oJk7AwcLoYvRahHV7hfLYoFBcagwk21ivgzfZNQB++B+2bkQqvRCt+E+2LAEEW6m
woPRjE4BFvQ8CrXVjn+tyeFQDkLx6ljN2CzxNEUpMkdyo3L9+93MqdD4wXmyO2Fv
YGibyv4zramdojICJ/bQuuc9JGeRjpDqe/n/jVWX4PeJKkin+jBu5kWYSvu+UY9f
bT1+HwZ5N1XK+u3Jas4c5PudzK4ogwQJvdZce/uPmJNhwoNlNybba0n5fVVKhFIj
3tAzoUFo5iKBnX+XvXe0k8wUwfaWTL5ZTeF5zctxDTuVuRsexY8YaDxYAUlUHk7G
m2rm+lNZYJGeXoRXxZyn+yBRVnxY8Gb5iPVhe+TR99Kmexpvtz2D7Y8oR05U3RTO
dZzc1m3eT2DZGVYkLxCa2RukxCpkgVi6+MHNrg5SYKaGdbrD3dj5AQEhYzEXVZOT
GTHx24OTAjUytYIHsGJCt2IbIuNqyBP1nX6I0m6TK6bqlcHIMFH8HndW/0kfS6cj
uD1lWnnJBuX+2+r+iAt0YeUWN24hBQcHHScMeWN8ujUqHPzzXFQyE1cgXTqLBo/5
ZkGlvP4Smjs1CEylLHX2qV3i3U4zonPU5K7si6MJTt+x7f+cRNjmLlruvOTM8O9n
zT9rLhGOIbXXB9GksCkpiZqPU4VYAVy+qbOq7xF6yabsNrRWP1zxKEaFzUl8wI9n
YTnmnyCl9KYN5MBzZkYF6QhF1Wszcb6EcMu8LNow72FA3JvLOoaETMSaipsvRalL
qlDbPgPXvbTNZ5tm/NUNeuDTytFxlkT8AV3yOmEkP4K2Y5haoOFATttwmj2szuSa
/UHhzIJ3Ww6U0L3VtrElvsdcBnjskk3G/ls4+35VUUrLYMZ4+yn+AAVxCMkHuKyi
cei2W44hK9f4SH3WhWXUjapyNCybhGRRIarei3nWAXhe6la3FOdak7RsRhU10Z0y
FjZO8XDeOsUuu5cHfunewA2HmJmrGhqIHnTM0npm6njgs/5pXxB5Zp8tX7MXPJ4N
1ELAlHm23CnpdYRGmILV3A0heJUWCtt7uN9XwBH+2o8A5WCFBi2oO+yeNXDaq4K6
S/JR9yXZRkLhJt45vpp+T0T8a3SWizPuQH4mXY70X1LpYCZjVm8oIJy4ZKkcaF3F
X169rTLI7Xq1Jbaos9lU81j5q/5w7OCbXkEer17lPWCDKj4a731vBGD4Dm/HttTJ
fb+G/c19uM2L4SI2d8YDu1a05WpLNKHq5WQy5+UK1YR+DwCrNkcaNhEItXeGpTl6
1N3+4Gz/fF6K+eAetTLHQdf3t3ADItIs2h7SQj8vMpFG5u5KCedgIrWyMgDoTvQc
OI/Ran3OuIGMTvdBLbd5aRbPRR4+yYhh3+26+XNo0IUnnBGLOFsfzUXvGY56NCQU
9WXKqlbIsRX4v99RHYV9AGiomL484XajGVG8m19IPbWuAsgZ+JV8YDSziCc5EYrp
paGvzIsRRexvox6P+qI6nr9CllRi1t90iFo5I+M2X8gLi+zGWEMGkhdmLDN/JnYf
gBImIzVKK/4q0/4A1Ob8df4q68oJSE/p+HK2Gt+i4SwmXZ+pVf2jguBlNIXlz+cS
xahvoB4oP7guB7mzVyFJJMOk9AB6wTNbeWJqZGTnykwbWYH73eMh/i0l5Apik0q5
INE+rjb2hx3zA3+KD55a9gC2fNhB1elbHe0G67sUcVMdIncMTd+0wRAFwe756nJH
5foJenWJBJ97Kcc92xOboGJ3ATp/wCmFiO2yCywJBwFjnlx06op6HkHsw8YOQ/Ck
cGTiOAcVYU4mw2tFFFgp811h6R3pancA/U8VHPFwClpT54bFBXcpFwH0ZbUoyy33
8WHAKGNXsnmWU4vDH44L+RLpowf6DIUATQpew49bMD8mj1n6A2bvacRudJsOHiRa
S/ojTI57yQqCP/nGd92uLx30zVwPiCBjchZoip5QomUWmQ0bNPFQAEWU6eJNTOIr
aNIqR9ZJjUX8591SLeehXlGIO7ch6W/BgdO+Snvs3I5Z+Dom0VlUDtHHvIbQiPlp
Fl96zvTx/ts+1Rv6EJUZQcMxBjHUANQzQTo9P6gbJ0+9LIiQaC9b537sF147PYLb
IVDvqkAy+5apZKh9oe2PzPsznHAuhHn5HgY1Wh2QurgmHFLJAoY0SxqCJr/pmXmV
GxO4BfQehZ+45lXoWKHwRuw1zC7vBWwKAnb84dmWT/NiKvJq2vWC/DyC7lCH+MFL
AzvvYO1tX/xqCIxRuVicCUatQXpaLi3pUZF3iJH+lo2+7jaw7KfFucFJNL378nfo
az298UNptke3iOSQ+4QJHBA8imCllnEaj7OR1kAAwpoLXDnqqjSAHxkUfEwuTV6r
E8PBkMMU7Dgqws5UUCNiGRwXr9FJSSIHKLjoINNuAdURK2/MBnhNGXOVfykiC8Cq
ePvijDX/136Pa6+H8c3N9HypAXxMtGIAu77QzA9/e0YmJoEVwSv8zhf+TUkinvNo
bfqC172KDc0OwPM7ilBJkBzhkJH4e5Cf76bWKaTr44ngcljkgio81CwHqrto5gPR
LqoYsrfdbDlebl11YBGdaxdn6bfOfxrM1ft9p0iA2twTCELeS4nnTsCa/voBFdvd
4ra6lxj9fzW7vgO9AJbs1KCIw3HomWeUdT1gyaqxzH6ox+7o8QgCauCdlC+NirDH
yYI+Znar8wQ7H2B+5n0icOdbB3kTOoYZcX+ZHyGnzwRVU78IDziOMKa8hDoLeVA3
qZuG7IXpnpxH5+HQ2S1Nqt0bSbxahJFHcU9y8wS5EIR6GJg37f+qXMSo0q+/nbQP
qzDVij1Q2CXozHquQF1hsjJDFQkB/rGoZ4n4/hnF7NnFJ948JgG4WJVV/HTjzcuh
BzZ6xKQbRQP/W+AFjJ7ihsWMZixq5xBRSvC/ueyk1vZe9oZft6A6NQI345efaZfM
HI86Fqcvn4fzBFLMMikdq7UWmpCJ8x9X1E516BaFmsKwujElIJQkWfmHU517VTo/
ICYc4QshhWK/d/wUkVJJ0XFTZ/90rIpwWE2MnXbQELH87VBhloa6HNxiY8UtU+SX
e5nO+1c0NS5eI8L52ZJ/9zJF1cdkVABytMYupCvcoDEnHDVMo/BaTy4s2L6ldp+o
VKHr9GhxEU1RNQwSEdKKVnen2IKm43B9WwAiEpLizOexZVUVViEjpgP5QooywyYX
+p2i02Pn8RHse4hoBS1HbkQr9B4SbU55c95RR4yKw5I0XDFDyfGM7MVZn/eAQd0c
Tq/3/rqCV/jMDC3fLtRdGA52WMFHs8O/YtBpp4XhLAMDr3JNR+zM4oFiygdLCs2t
cKyDNAoOwO4TclRoqksluQr70FGm2OOid1QDG9GuN9imkKe7u/KEu3cjFoeBTFVZ
S1dVx259npqpySDdd/tBTfW3nBSdujS6HE7U+FHHr6sB0Ns/Du+Slc1fcuocqbme
GLEeok8fzxDREeIFTGjOZBKbodm/LWyx8S3zpZXhTWi0UC34mRnBw/gMVfUurEA1
pfpHrQ9q38C82nLsUnwaPygBaQjcxNtbj95rGNUH3okNXAG8cOD8h3MziSe15HQE
v7pYOApAtj19adcsfRj1jp1Eryn/kHuQtgtQrqO6XINMlK9WQKFs/jWTJBmZcR7D
YnALVx/xjJWYaNwlzWbhimBclxtIKFEK8XDJznucjhLu9QvAs/MnQ/GX2r0pMpit
SEUFrRxGQh147q/6O8nk1acfD822JgkYNp6AWFIcJlqGzFmyWHGQ8yncf5n2EP1e
ahO9xVFuRGTs6ROBP90FfllNp1tHrvC+a81nNIYn35zHzJfY3txvP2eVpD14WWA7
4BcI/8bWt1KXtRTI7V4IUJ8EaMOK9PdIakUAGh/juKaGZwtdl2A0Ikzx0YQWIiXW
K4qOc6LJPOnEZkOWHp/25TUs9kxQStjhMuJJPfSTXul15ZDIaafrOvspjukJDMlc
J5oWTrRlIl51dNXsN7fAo1P4e/U9bUtoZwi8JMJ8pY6betsMqjoaJM0aooWK9++Z
TVK5yrdXrq2iZ61tATlZcBXuQZfKb7bN3TM9G9P2To1Ggs35K9wLQUMbs+buhBkU
7xYGhGhbO0IsFshX0TYedCg0u4T88A7cg8NB2moM9MmGdMd8bta72vkODv7vrLkY
+yQQoZ0wpXclE3MT/OHW7hPjTxPtack+qiQPi0D7lX2Gq0vkHSOvUO2J4xeBQ+ib
TEov1/ng/WYXpl9YnVsPoZAD8+Qv71w3QRM7gBdDAFSFQSYdqdWhACe5H+hisHXU
bR0pIwOvqO9F0fi+Vg5B3Gn3hCXgkUDi9BtgJjHLiIO6UpUrKAC83GjRh9Pf8g9F
shkzXG/AvNF69xk5mrLhNPJNtV+CtQR8Jlh90LE8L+RvVHqc7qMSwfgnjZmUp8kO
o1IQjLve5fsHYJ8XQWlo3bKF5s5UpWGY5bD5tXRXHI2v8TGxbnryxx2QyT9iOg+a
jNBzzY4WZTTgnF5T5dM/ZPWVFbBc8Xe2S+u8JZPgwiaDvJFao5HsuZT4O78jcUt4
EIlyCFPmHEdR35GoqZHFJ+oO5eTjnv1jR7bd3MsWxXN75Dbq+wAN4rZRk17dKOw3
aAhBpcLXHkzDZqNXAtkvKJCkGp1Cmq05wLSwenxgwQja4dH371OcJG5L2SamZuWh
HihJeaHszF8GWnADxW7qnKgUmhAhgIQwr3vLZQYrUAU29UqJt8iRdons51+e+IRT
ANVXg3sY5vz+8IWqYC6DuiFxYFwZhNuzIv6fmq4Wi33+soo/CAYUwUHLPjhRhjuv
0pgPqzTAO4qSTRSJWnQxOMCwSE6R3fSKYWZ9mH9aEvlfUQeKHqYMuWDtzqilpYmD
jNyxcqU4UfGg6aekW8KqzB7mttKQMO+gZwACQCeAI/qRtFwNLOWlmdrrKYwfGqA+
WWs63iQdQ6RBtE726JsjnGY/exAfxE1LnBXeYYGC7fZ5TMohNMwgSTpj88WvXUCj
9EeMCxk1naLlendQTdKCkRj6jikdCL0KJxF4iEbv6ry1zeh2ejEoefTIKpHW+iop
yuMsVcQ44cJ1cudvErigyaknsMDqCbO7AADku7uKIhSWSr19DsYrHGnTUJ0zzoGJ
s3BBB9G1U2CpVdIdcX9n34nBGhJ0I/mcTeUITKrtti3U+52Aigz/d6hWlKu0VgjH
6dch5o2ALOYIUJASDKshccU/JhiynKn3CGLif2BLP6WJnv/iGnSGl60/AaIYD+0y
rNkRdHdAHQj7Ql42j+CUn7szvKKHhT8hpEiVmoVnoGGFUXC5z43pQTEHmZ0mIwXJ
NIj8/vwoJyRlRdTFocKXr1YKt1JQHDqWFvp4L4nwovhtyqeyI9N79/aHQDBN3QNS
7oMgrUTGRU1wFVss1j5qlc7Ev9kHPkBJ5Pc9FUcMMQNPl31R47Zm8FziYXHeR/ml
swQLxZJiBUZba049mQQP4GsxsTY+wWuihWhgei7TMJO6ohRxeCuwsNZtNPjfJDg1
xen7t2cE01/q/F0FXv56nWy9YI5xUTqOpnob1wldzwjYp37do17PKvq2lZV0qCIN
IpS2K9SCeEJWQnAIQtd6EuxUcJZzUlnLQvoQDI/xp59NzNCoZPDUD+ZyiPYRi2nn
YodN3w2LnbxPUWMwKHRu8Pw2W1mU75AFUuyoSd/qGKB201NxXuT745oY9wNeblHp
KIXVk5+g4mrdLu8Bdwirfg5o70PSmDa7yzfWHYHWNWF6t0NFIJx1A5+0xKZTbJU2
GU3HGMcxTaKd2bJS3wbwmlWnqVVwJ5YfYSzpzwotshl092inKmjAg5baFCQ+1eDF
FhkVHZjF5DRfkdYkfKOPCjShI+FbZj5jN5eeihgETiGBCPDmjJ/G0zC0Tr9xqtrt
KCQFfMb1q1RYGgej+OMkPozh6wDWxzEhjEQ2iTecjCvOQP1FKOW9aDiyQV/1xcH8
0lWGn4nMNFBjzYEb1Gv9YYPAl4mYbw+UkkgPEu8KZyX6qR3bCYGG89lyvRoNv1Qd
A/PyhxsypV9siedBMFZyAsq9QZnKEbm1tzFm8G+bkr9Z91JfoYoz/ikpPS89qK0P
evHNm0DNFjOW/eBQYVvmbxwcr6GWMpdEPPZ2JZlkAhKIaPdj1nu2hFTbhYvbAUni
8NVSRK0hCT2mE8GI962Iu4cf37icZdcn+X2tY4xdjhEpUKQCGXAXtKJtYgMjoXwN
9ppMRI8kKJVANHd4vDqKnJlo/vMfLg4Iozop+3Bdm+sh1noNNmxRjbZPWJgFDKFA
OId8OFFQFtpr1iYUS2TpX3SWO/2ks1lgDzF+fl388IJjLOz8eLXwFNA6DezUGNcl
JADxrnv1EXc468iWxyspAmiS6Ucg6+Oo4ZUDzjEKnAo5Rrprat9fzhoTusslrJIo
br+/XGU44fZJkLPAwRw4cx91ZI9dX5cGZXk2SOZnGXMqH7myfTWzRa5MBEfZlbdq
uSfrGATfJqVCKwtjgiZsPAjV8nvU2MHSNNAVJ5NV3HoKv69Qjpyfz1YmtilXuROu
QTJu6RfoyTtr7h5zDYjY+wivSBJN9nOFKzbrm/GBSivsWZ1+76mdEXiUw2+Jq9j7
ASmL2sJtJ+azaQwU55CZd4GfM5oWG75qtuBU6YI43ArIHGrVGAsBjIfaO2vns4oD
5AyfKjGNIYlWz31yK4nLg89GlSArDFBP+M+2KTOOu2IG/1aKFJlT6oX159aRrgz0
7BVDgl4oTQfSc2W6fJ8Nj+vyMQrG1eg2jfUfzHEx3olpUkFwIoIWXbF6ChcTvqXd
BZzj5l70RPdQwClQccddY0iqH1cEEkpwLxbUzfeVmPCAZOdmlKtJ5oPmkG4ZjsLq
XX2d6VzD/3WhQkdhajyDe2bHomRlt8fy2t21TlLDep02fHYFaG5MRWkjK1s4a6gw
yfmQqSQsRMjIK+pDVHa8c7Zzc45yQ69nk4YJbRODEF1WypKrjNaVb7J21lF3IklN
8sF/XtHHD4tzoE7LjGa64FZ0Wwxj4J1wmuC01xfP9i1urLTrXCp9H6b4PU2567RV
eADU80Wk/Y+SiPJkWQzhsYlNOHTCFT6UQXtrrV+dhFTfXOrvt3GD4b9XA8Pnimb3
HzP99MP0JayqjWNv2Ef7tJut0VebeDey2fSb4EWOyf/BKcxA+etST4+mnyrgU/8X
TohpxXFmlXMz64ucbd6/Mv+whsaognRLvhDkrXLJioMB+slZA2bVBeNmhPLeMSb7
S79pDOd/dIP8bmBsduTf4nBCWHTELQHw96r1hIVFXU6wIKKK2el+hpbAtbYTyVPU
/BOOm4p7xWjTu+YoV90mshQBYb6B2pPHlvBGklpXw1wUZeb0f7QCvOBvvv1jfQhH
GWFEepE8E6X7LX+0XYcL6JKBBymtW3mGJNneLjS9XctP9vRBChUEXreocekWq1RQ
RNoHYQYHAIN0V0G3pZa9YzKgxVWH6I6jKnV7tZXUOvldEugNopmEAfPqjfV1yccb
WqbyioM6lx0cKWzLhEsnbMu0LkO2RdyLEK8mBelVmsB6FIgqHx5GyxBxv+iOL70P
rvpJicd30oo9TvKH6QN0GTWyik64nKzprA0BcZiGCIrHYnfwpY95jZ7D3Lw7OAIo
Lgg2LJJmBYsI7S1Ucjicx+VSN2qGOpPj0aY+VqjRxWGEDYUb2pq/ReA/zPrXEmTI
KicVC2Yc77kBWKH9wFtsBWhKKU4NjDyIpJAldeJr8FGP+6pdtziZmDj/9HksDruQ
hs6MnNlIGpvyohtRG+385+r0WakmczuGBgs+370Rl73Bj2A0ePWDRXih2Q0q2c6S
B/+Ax+wQDSKo73ANGJDCZeZomri7vb/2uk3qXZMszEJwErUiyH/Gj1ITy/vxVN0M
HPZw/+WB4/j3gDzGTcQFkGPMfsH6Nm8vKjT7T7BHEJ4If/5zf6yG3AjTYF/Ekr8X
9K5gBnvkJbN123380I74E9ZKTmn6h0DaNfdvTOTAKqsU1rwUXp4JGelLt9Z8VjMm
7QtutFEqUxs3+Y5qW/7anh8EiEiSh/f2co5C2HA/VOhGBNX9g+7hY7XYJm/3i2le
CPbO+BlECBtTBVE3stbAd0rztNNAigrUZHz9braO+vKrgnQJGcd8x2npYRClnRpM
m3reyRi678rw+vT0k+S52TMlG6yWSgpcfbtsxM+g8hnA0BEZs5MNzSJC9Wk//5aq
if7X4aW11a/23o+1eaziQSqtFnG5/FIIyJHFwxCL5+GIhlvjte/vs5VCpj/c9weH
lDp7bQdtr22yIDFY2gl0jO2dXsQapmM6mRZiHU5CU5P5h3esGuTJkv9Et6C1etCz
4EFFs5sisCXTe22JhAiiy+V7Hd14MqDYJeSkruJ+rlBw/y2kdInvZ+EdS7iXByzH
jSU3atnIU458znQ8hGrSl75jmVM2OThDTRaE6r7ujfhMX6k7CesN2C3/EX8xBDJN
YWeWtWgA5Ir0+PhHtNrHg4gRoH47FivPUceIGNGHZQ1PRxUMcDUr4cxDHJ0lwd62
xhRgGjAeTJ1eg3Wzgltgqga9DPxb4wluXomDqpeBPZRhgWD6RPdUcp3yUMVWFrWE
1c8xwCN2VYOI5Q2BqL3nAS2yEC2AQaE1pooh81P7gVzs9FTIMGhpWVqGegz7PzLm
MFNKdtYd6iOdeLmze9Z8iS2/FPSYgea240BVEvG/m+/JhAE1pZRHS1dnIZDrD5TM
BiRUN/ewh4gSrQZM2LWxPWr4vlkVSGwFGyFWuq7llYGkQvJTdlDUqW5Wvpj4B5Qz
8NsWQTw3aF1XYjgHuUeLvmUAknb9FOGgecSZLM8oWMfJ6LJzNQWlMj9a8QzrBXsn
xE6yo6kV0uE6z/uXI71VLO9S3QR0NKCD86d0Sjc5V/BcOju83hS5kFagV5b55h0X
OghSY7eiFj4FKbOfwjxvEakgYRotDb5yOEgT2Ud+PLddrQl8ZHC8mbo9fG+be0xm
HYkONonV2LwuxCrZGW0c2jaPpDtI6+SIXzMCid5oCPjURncsb3UZyAzmyPdTMthF
fU5jlUzzwo44OJ3J5dqhEXkEJnPN6L3Wul+4ffioE/RNyRE7AqupsVlH6QQ1pGB6
wInxbbIExdczHimuqhNU18GOnc9wnL8Qdcy2g0ecBrDKdeSZ03Y3d6Sci0WCXySh
oHOXPm1+T6eSIaE6Dczf6j8Tdq3YtisEJ7xs0v/CLkjf8I+75jSRG5Xjo8EnyMg/
kx9YTVxpWdzjrtNtHz4qZZanQZ/YqCo9YJdEHUA8GbFXcx9wGL0pyHIASTMF5O+j
KhmGiVMObmrOb6AXpfLN90NegHInDgbdmwk3WY5MW5E=
`pragma protect end_protected
