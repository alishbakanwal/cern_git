// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 13:57:46 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
P8A084O7BPHY/ysFi6YPIlWyecENSaSbynhEfMzVolUC7gOfzSFMfc2kng2rZTmC
+75oPoQr9FJsRBuoYSWUenTplTWLzASAEMJwHViuZDUoHJ6WERW51YRqTt6rZLvC
ogtarUqIKugkGf5ULZW+gwNUw+oA/bH8NumfQv2SRW0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 22080)
ZF+7+8bO842wH372oEIl9LewmA9npYlwXUgggJUHNOiOKvrJZQrpaItVo+37Ivwl
N/nRk94DTSw51I/jgSBZ26Xl4fmeuSlGCfyFcX5niG0z5xPXNTYn+Vvjme7VLpve
ErKS2RwtYwIhTECCf8PzjHkuIszuM/7ysi4IItxjhKO8lYhI+CK5mBiJmn1sBzUY
dToK3lnCGGmJg2z4npZW/vBamcZBGBpc5L2dT41MIctyBLprP1+Dvf0xO8tdtBHK
C3IMBaCx5KOcjZONxwvE+qPtHR1RKezqLiLueP6USEe752xzeHoDkS2/X7g2AUz/
KwBz6P1tPi6IIPRmwcmfGd0ts/kgJAYdAZfAcRXLvBY/f9vYxq5rHvx9Tk5kHta0
rSjG3pBAHrmkMuXwI2O/GE5bP9MJs8w8AEsrABAVSYs3hxsamcDpmDeLA+AJ24/+
v8TSsicf+y8PErwiQNNqCKB2w5aaJw4Ir/0mX1W6BcyVEtH42WtJEYjd5+/IV95I
tehYBcnW0vbGM+zlymW5TPBGvIPZkupprAxIvrMwaDVHKZ2OCfhm7EuuzioNeqTc
QfhoT6uNOFvQ1f3VQ8sLW3r9Sv5SwfcREd3J+HlOJDDHLnduEZI9qU0HOj00LKn6
TroeKA3Ru6s7/Iakr0EcipkFcmQ/qLDWg3HTXIQFTErxCdDPTZpVBDM3FfKv4ZFL
eIRyEPUPpof847SHBKfy966yuY6KAEmqtiDa1fzOXMs1NdbComU4rgk1WIU+pGkL
RO76Ls3py7EdATdMPNQWaIhCYG9U3PkwNhlLh2jIEIji6nd7RlziFLp8Ey60pWGI
mjck4f+eQAao9vRAoPhAnbgULbx7PFUHrX/CJ6cIvMyGYNrfMKZaoPl667f70sQ4
WHK63K1EbQrh2O2sEEcSWNnhbaSa/d/qGx7DABeWr8sj0IdSfB0z4mavL2rnBznT
I3JDep5nPpdDwbcRbm/2rlhwy36TDDKguCYcPXjnH2mAJchzh8DzPowsCd3xMvs/
cs3TZtJbAXWgf+4bUAoQlikNoGGMJxWx1I3X+c3U2ImhjQaOc5mbUHm8mYvsA7lb
sBavZvxwuc4KfHNJl3RcP44/giQAJtXNpmro0bt36XP8MzxDzFyoYihEW2UNuAkz
hZnBE4+IG7KSugKIJr7vN3+uwQqf0H6dd7GNZhZOQ5hvsMCreq1Ym3zIO/IE/aQz
YihTtySuY1T6bw+0ml+JaUjC74Ky0wWDyJbxoA3ttn8vOYbYhKOI+y9ro31Aj21d
EX78WnvM40q6RI+N3mrQqwO778qQHxPYgkAVmi2YqaFULGOtyO8J3YPNAfwMw2fi
D6I9LqECAfsnrI5GptvElwNtluJl5/9KFg4dH7ReGbTtw2wwZoxpFFG0UL9BCER8
yxeCq1c9TAq8tFcjwYwVzEcEF6De44bHDJtZ2VNKQ6zdPe8DMtc45fyBGml+8QbN
RvNamUmsDdFolKmB6Dab/V2tYG2S3/3VktNp60TNUbB/DVjbJMfsO7XUxfSOtNfj
UuHKMLD0Q7EANbHkclyZcXSDUGDhpOUZGoAOm1c+lzQrmDp3ZOu1d2LOaQnNerJt
BcSHCW31y6Tpay24hUyu5XjynVig0e+GHQKTzmvK6E2VJTO0i8/EeY+D6S9NZX3j
IifAZEmWTu2zPvm/GA4PWa+uJEFshmBGewbqTQfGphHtUgUlWXlcogfLlgZZmlDV
80udEXmTv6aV3MrtVnH5SnxsWv89kv7nOqvVnBlvuCK7ZxHvjBh6JM7j6WqlCR1X
XUhh50r7X/k1dSGYfSrf8aCzxZfjDlMdLY8ZDOS0hjihSdQmwMjjB5Gnj+NWPm/U
jWyu1mbUAwmsZp/kkLqJq7Ap/miQBxKZymP6qe7AFKJjtteX/aDYnARukkRwZItX
r38GUArnBQA6vTCB4lpER/OIw/EUpWCAtJPT8TDTC/Z/QP5DQbjmJJckMT1beq4r
O2Wim9b61tCciOMH6RTQMT7sLM3CRRDZkdCW2OzKrfEX2In3kPJqNG3JNLP4A7YR
7gmmy+CxZZl0KsXCqQKbbRwGuH3yZgelA//kk4A7o1bXPPgLSJoL8kBcJvhzPOUt
CYMhxQvOmU0iIA9o/+wQSOq6QaHE0rxtT3wX9KnUea0Lg4sv3dYRhwi+SmIvveDY
WQfq/Nkcu7JTOHm6hI0tJGdaru616vNjQoTl9F7aUIqw02ieIQKt8MsnsayRvjwy
DVZYGc3qQ58Q6dt3v59wZdUbnDkAthyi0dHUDI78qvj3s90vyz7oRVbevlLI9LUr
DM/U6YeC3HYDdXNkIqJVPYD5LK6PQwrvrisRWOWIE41b6O9p/+Ct2YjjAAwxlOBW
g+blY7PA5ZtNT/5k6YGJz9hHl8+mQH8sShQtyaloFElJSeVJbJpF+709bZBPTrdR
nluqK00qiMQEaT5ApA5f5BZuhOBxUsvnPI002w6E+XcB526hCXCHsuu6V12YRwC7
4np5ZuvrhsmOkwdW+Q/ImFjm9DKRzgzNBmpSjxdf9zkHFnJ9zwsddaggbDTqdEWG
ST5ph9SaC5pr5OSlLS+CjTPcvctkTijcwsxIna7HSF03YPAuhnT6+Ag66Ag3Sff/
Rn1FNgTOQ4lW6TARgMySSajaX+jfmvJlnJA88wxMaxlu7OCZnCOADLEMn4Ng8qDR
uaBOLSdMcCJ0kG4zHu5yD5OEuvtxHewDO4cAGulnYfiZOlLIg0Gre03nUJ8LmC8n
/LbgM63jwAdAzuQ5SsRF2xXwZczi3k8KA50IyPz3VBadSrZYPdrWkQTRYahM8W4K
cZA3BFnoFT0pTMqXWI9GnUetjfnVFom/vGn6bApmCWGw17D3NfI/dqES37NNmLgd
ePP5y0Ps3OUy2IoQOhCCizMzw6JGUGUIWItI7STeegU6J8JRKd2ACC2RBVfW3dc1
iLhjDGRSuq30puBbNkkYhZo0NQG0c09lsBvt96b/V+7/Y4FAX30/10bs4yEegArV
PaJncX8aaXVkihE+lAPy4lASxDrt/n2MYT53S+BNW/IaSBKHcBw7varib1Lgp2Tt
KrWiIRziL2Ue/1Z50wGPDtQr/qFQc7yusiGuIWI3dHwpsyGrN8GC39gT8MXaBcYj
4NCVjx1a4ehHLRLNWB+/7kWTiS3mF0LNMGrBnLcpaoJgQhaqJh16DCqQyYNdNr0t
4puH5ZRirnDySJAw+Opff/e+ZvQ8I60K1a3kTQuTPE2ulbeERkx6tks3g5Yy5w+h
HGRO0iLRGShurt7WJliY1yYUtkQgp+hmmD3w6LLgEtNMrBP6rEM2cSSW28k+JVek
ydSghEZS25GrPMVPqS3LKS78fGaLqlJbvrKqUlCQNYZAF+Kjrh24OxtUWgkQDEMG
gsaZ12V4iG8OZJvCsFjW/7U+4BgD49WXQD3Nrd7EnfsOCD5Aa2TGbqwCfT4EcU0Y
m0po3dP2NHiGI9lt5/MaZ8qmlzvafgd+Xp5vIK+3z2V6mZFtCXXJHhG9Oct9J4rB
Go8aJB/mtfyKkOh4RU/0rBRwkrq2OozuhV0fxlrd41kZZZpQNT0OZohlZ+MRMA+M
2uh3dLQfkgtuKFFROH77Q45IGgpCZUJ93P/y8+ehkAdUvaNS4oF19S/8+Hf3iABD
WK2ForN1jUahldMP+d2eMYX6bP2EjctH3SR5rcjuzZWDzNUOBtuSL63G88LnteSR
acsCpBmtqAYxZXwaMMYDhrk7xs3LLG1wkdzzYEfNXvzXlfzoFxEDIjWWhA/C/q+4
zJ7CD/3apJqiTeNMYE+/o2HmLRo/Lko+6ECcWb5LDac1XyZUqnZ/R43Vb3FAPyL7
wczmgcZ6xnBBalOR0QSM3ewecD5lIQbIHRchL680EcWu3CHkxSh74fq6NZIsOTFT
KCwhrFJBqIbv+v4ARlY7wa8v6D3qX25QHxEf1G+Nl1LHWzKW7Mt/neNK+N8BdBnp
kuJsePfAz9x1NVcgyVR0y0NYvQCVfUkKQ1ilZqgoJjgZx2xuk48bfapOwr14Z3ny
jAbJb5IeTbR/LZ9yjVjVwMO6r3GABeIxWRmZ0HR1iDiZdlhYRjZvMb/pm/oKGFp6
kwRQWmXWtD2PAg3SJmfwO+beyBSstGBZz1jRX1FoiLnQmEj8Opkc909mEArGxzIE
3hMyNmDi2YmQzw+vReHWa0rjwyvy/mja7PO5TuUQCZdeEnJq0uVRCuWgkV8hoUqp
9M732xU5jfDKOeiZTPbHvL2nXM6oZb7lx8NXWzvA5QNzujsQEeUVpUgblx+yHyf8
hscUdoZV0fuJv1Dw2CTdoGNBPy8iy3f3pRfs8411jI1I2YOZUwqAJOaoeK2Oksv5
fo0CWh3Xgmnw5cz9PBDikqubeXYcGawcCBIU/OaZ3gVORAv0lf9NsqcxLeggAOG7
ufBW8SmkNy7Qb6R2t1VDS5okgqCXnq4jm+KkLxNM4veRhvvebSmmRlKLbfpQz7VE
mCHgN97MPF+Y9PVHku9cqqsqGnWVfARcQNAb/3d8G5nNYrh6Diy5KP8Two/y+YjR
BCuIsHnDmXsRm8e4ckzlNj2tDh/mroQQzNTeJmtTczp/O4p4Y3bPlS6ouP3oUGMd
UoWLPxIoiVEXyY/IN5XZmUqLF1af9GNxOwY5+wJ3MDWoLE5PveJhCMRv/KZUw6t8
5YNPAV94K8PDckzAq71UgtjbO9Dtmm2LcembVsNsMH2BEmv/ZAfydIMTBm6JnyQl
dzRKmaOStKcUj38+kSFxLrn6Gyf/OCcgfb1tQDQflGC3f+sN7w+w5RByoqdb2WuV
W/rptTSY2mQUdmpzQCSRqbHxnH2AGhL9qaFScapf4urt4i2Fcx8t5xF5Ha2Tc9Yy
qrTDVHBeeRmv97UMAKpe3qjwSbz18jOHRxU6PDda1hV7NajOXONrKFYHvvgpqSgQ
BzVMkhb4B8sLm+/J4egZaI3EKniO/wXfdLRwBaR/LHsIVdBccuY184gCr7ZWzf9T
J18CvBvFIyKW6yy7Ax9MGvH0XbQ3TCNE9A3BS3WuwDcKnEV0V9J5lZY94vbYyqXW
m14CxRiBGXTQsvJxrcz7NWe2wNtpjn7tBrnYYToDM9yFsrcDB/geKFk8SvFhzbT8
Cw4ZQ0td3+iug8Yf/kHzYoTSMas2+iCbIShrxKStCGBR/k4BWVxsuXCTnW48Pfm/
H6TSdOt6UyRl+PTShj2mNQKjkl+4PiODfh3DvChaRIGpEF71NZoclEt4anLkeu+D
y4GnVpMDiKNcRWVnZDqFP+Gg2WnnyE7VmA0e0AJcP5tcBD6c5fkmMT0IlyAmsKgK
EvnjdAgUKWESnv8mdBPAe/D/IHhr+X0Be45ShNI/tq0d3Lgl564EoEhYR1faR7H9
b0D97v/k4OW7WzHKQq+oeSn5c3CciYD/83TodxWpNDC6ECNYdOU1naQYW7m8pXk0
pWYh8fOjmJaRYdnYDpVCPVPIxroS3Wp8kY00RQhY8j7P/NdbLhfYdzWi5BCCUies
vOvSZM/8bHhg7VUL1kZj8b15YsX+MblALLqFYmEYBvz/9GHv0Ph5zjYwEfAAh9KW
SdTknfyBiUfGT39oPfQBTIXbMlttV5LuD/FYOE2INvBNYNqV4L0klpMGdWMgX5q+
iuAhp3ms5UORyqlEle8Zf5ZdIHvU+abMJR5C/uq7tMGuShsbzBJUG9HVkoLkSoUz
XbScGLPIH/f6TrqBx5ytkuARGUZqs1dQ2FmbLgp4MIUrZszLBDke85VP4SzrItju
zPvsqz4fqMWPfkmwj3jDi/uKU7v/J+4wazxz1Drj1o5ohoyzzhy3ltsQp08Yz4fQ
LKHpwip75AgK2V6zOfoLkPtUPYBYTu58tf0+3+vNr8U4IAZhSZp6I3T8ZPaYuKeD
JLi09NPV3WOm2vzKcF0cYJZofAdLUkGJC6/QCMYOMY4erwf9WcrYdsJl6+85s+9v
JKJy8QHpRwx1KTagQjG+8aSYhJk9e1mqW0XpbENxsrj+mSqrMIPILZdejP+8rql4
5WYhmi1LC0OtsYUrNWKGNvLsyhwZKMwqseQv85dvqxfvLpGzPVNp4pfryoNSz9Fq
94m9rOFCb8C8DbuhXX8Km33h7RWXq8pFHF+vo+HVThvbif9x5atG3yViDcRCSz27
54jt6LYkGe5wZIJUS9D5cRAApd9r4CD+ntQKe1QLWqZCQcz7oSN/tr2fqKX1i7Li
zyP9tIRZRyylvhr80J7vxRDkal9JsJVHC+cQP1GjmSLEnRoZZDtN5zJ24smKs4Br
fl64UTzvOtOFFTN8TKi0vedCVZYGu7l59vKqSQ8OLqV7oY9k/RrxmyXBhJVqK3kE
kL3W4mnBZ5KLMU3cD+0rxR+J5tPMFX3UkvcevQcC+IZsysV+oCs6F68XjIBQ6j+m
cZH+tN3SMuToYAm7PKwMkDCyEorhTyU1hk/r/vgqVIzieR82wsoFIPHYfSom2cGN
AvsGO0UBhU9b3IKp0GxIUnbiXAiTVsP3UdH+GOvC4tdpiLp5Z4LKDkEB+Fttfy+i
0E2u5s/J+ZT/hziSGyUSpBZeXrv+6u/Lp0hnfpUDjQcc4MOGIpPvy5fqiAO8i+VI
a3hLAnfoGEBpGkEa6ke19xN2SxZd55QsBn+j5cuz4aftlzrrpEeBHVQJ2asVAp8+
y1lVvOyGwKBzxvKz3FWSAApSSJFT9sBnLvn1ZPjwGEROyzI7LtCeskKT+OYSOdjT
goYR5ZLCjlAPOinJn9V9htsNhRIHmlTkn0jHXhtuuAn1vZ5kuf49yMnLVzxTmpRc
LsrhU37a5ZQ2l8aBRZFc230Ld3VKstB23e4e4HZ1tBVEHHDvoBfzHI8/oVf/7u+R
4VzqCdFvMMl/+MWG6stlh9WeH0pvY+zrjCuJJElKVLdSL61/7mxyTEfbNwWBrmCk
tdlV1b7DSlZzJSkHpC/M6aq7ClskEgG8buADiO0plvtpC0/lAeSho7or6FUrvt57
F4OTDJgkyz8SnMD+WLrF7paCwhh6Nf8/1kWEcWkXxQuUMTrtTQxt6EBkuXEnxZgh
ScD3C2ozoeqo2/bb50NzIMnQKg7DWbtUKzZd6zt1R/rUBCyFVwVGh4qAo9U+OgAl
X4WPSR4UzZnFNOhELpYz/e0Jjky4QWJLsPVJSjAINK2gJSNQ+VQNKg3rvCJ8+I6N
8dl2fNzXS7pGSFZsflea1gPjykjzyCtnYYASJd2IQuLFCAOOlFskalf2uYCt9Ire
2rtpkFpYtnhWRozZZiOGW4pEiepUftxanyzieMIdzfWjsL1PnqQkRnfmDeuEKH10
z1NDaEch+TkDwvEuesEfnez+zkXogtzwv9tYadHbeir7VF1grmyJZQxomDU58quo
eSjpinrPkaW0aVm7gKfw3q903giIRjpdupWoFy3ReViazJ0bya2yWKehTfgXWWqG
9H7HuJY7anZd3lchny9GJGSfMwlYHv0xi5BluzWkTcg61X5ZkUKA1MRx+bhPofv8
+5ZgbEgwTXO7S/EKl8DtsWDYI2Rho8l7fQVIoBFCu1tSKmdEmLPNs8tYG1Sl0z6q
5hLT7OZ5aItHj9QbgJs8Za9/N+gVCle59Q717503caaijSUQSac0gMpNt8pkxxtJ
QyUVR6RYhHoffhvqu5lhYTXqXvsSbhGVgbelw7arUVety3IxPFHUV0ntNLB7P3PQ
XbzlAdTMmfrhXT0jasWAvL9zSkCjz2vypYJhSy2yCORB5z8MgcfZsU+bkHdk7oWP
kv/c0GtcXjakM7CuRVn7gS2FFU/+f4883SRQRDqhfHy0h5yd5IPHevleyomX65Vl
2xjxVuzvLgQuxuvuPOvYA2+0lj1uyCnZr53nBdmXBLtne7aaqFYUc4wlXQ0gMV5R
+0m/vcZF5wyZziHpUsabepsKtXH2x/UtYRNvVGBV82nbBITv41bzSEjtVWF2wlWO
CR8wtF6g+zU0o79i5n9Z7gvQXPEWr2mUVqiYp3JSxPc0zCvPJaVsIVdPHdtjn6xv
fFOAc+cVDviN6SGdjjELxnI+RpzzT0nvFLaSTW0fdyOfJH/hcYKnDWpc035LTzeX
pJ3waqNLaBlb4a2pXU7IppC110mzY8VshSPHb8YYBWcHxTpdanKSEmWA1LJFCYP0
ubDfvn5b9TxzsCCyoQlWlbm2PvgqjvEKkq+wIXYN3rHVb6OH5+R7h9Lv+ysft5LL
dj55DsV72Y4FvztC2RWRs7HrUmV+FdFcpc5SZNMs3SABonXeT0hGgXKE2ies8/UO
J9Pj8gmd88Tb5pJCb8B566vclWPIPSb/zAhcOkHdDo2LK1iomnYTCF1E7qAN8k2K
R4A3hYtMGPlwrWpf0xz6mqpsRbjDHL2s85AoIDUDhhXib9Y/rJKgU7KyOpSZofh7
MxT6+1TpK/vaCMjjf6NtvJxOu8MrxPvnYuHm0woGVrBlEKqGCcIS8Jb11gi9oRx/
yXXwF/dyAz7gqpCJIz2l6pbav/NoRDTUBJUcrUTpCYcJlD7BrOf76LTFZ5P+SIq8
vHOyBORMF0RHbLz+xsBmW0RpsVwSo3M1CRB98kBHh2Ktzf6Qp3ObgNNt892JAPXn
STMJG1FEmq3X/MrRjmkXVjwFqHKk28DRtUyAP/wGLVB+35QUP3E6tbd5nDUhSIZX
UFRaRU8Ehw3WBi8M+0m7YZB4rl6Fk+bF7UF57KWO1AdNenktG61Dua1TMRg3ROZZ
KYrUCwFVQfkUQcl0R0rv6bMZL715koBgmH8ts9mQVQr0xadrwRt0u4ukZTFevoFE
iLANaR/ocEM4gfa1QoTifPNwc2q5e+TTAW/qak7UYH1DthoeTO3TQPMJwCAyCevK
MtBSO0S+1bsIfGlgDEanyfgl0c1BG4lLYlXv28bCJny7llG3NudOWXGL61memWos
ty7bKGbgqBti/qdRjfrS9fi4aG+qFHS7uObOwJ0tjDu0JqZfi7OvEIKzoLH/QRHG
PkEtG9muENswFupsB//0oK2VoYdTsOD4sMklQB/ixH0MkK153POVVtoTbblVbU4K
jLzXkoeT51qthM2jOZH8VF8pVYv0v9JU0q9LeD+jqS50fxt55eKMTcO+rkUGKhdh
8TLpso5PNSnrWsVe0417N7w/1LAsymoK2Wr6Ama7+JYujtu/Puu/OyCNW+ckXpEq
8Psq8jPCyu1L5P7qqI71uJXYlouITzz7ZEJBBpZaZrsm47QnFSIenHNU0EDYeJFg
uVmbDB3Fd7yB5BOY3yoUnQ/mO5iITqonVRw9u3P1XpGRVxC0l7MJA9yo9/JTpjqZ
OCqeQ+0J9A7xhQQNZszNQpQlPnKZWcutgZd8T2NCRA5Q0DL6odLqj44RYu9U6iwy
22gMignOuqTlfBeKCe/ZQl+zG3Ll9pXoqF9M4tJ8hAcjJ57gyBfQJhR975ZNQhq4
fq1kWj6O7RBPXwqMnj7w+PhGQBJXjKDC/1oS7Iya4CSN5vJ9mJIPsyX9QrcY7igz
9f53d1K5vbGqQQejQsBTvG6MRgW3K+iInfHtT6t6H2YnYyqycEVJapI9qFxl40Dm
MO6jau0lz5NqRpHKR5CUNu+ZxqHHBjh6+lKdTo5pl2s484j3I+Hw/iFYnjtGAx7b
PulkvuAor9yFbE00usigV+NRJfE388+ttlhYkxMy8JOgdWM8zydViX/FLyPqDegc
JTVhbxbP89lRdijxs1KdIMAeGWoZaN1XIZKsNxkYB9amYPiOPrf0UqUEzz1j3HN4
0AgDw+aYeCGkpf/mogXtLj0GRPfeQn0HFdjVgltxQqgVt+bHRJm2fpmpe6kDzXSp
QRq6IdDZ9I0EW0Mlb/0P8c8Dqwq48GgmYeagWrRAIeMA74DVAlqzcF7odinn8HAW
Ct77+OgR/tHlaqaT/SKFM7Vn5CPQIpAo63kscOFNUtde3FEdJDbZ7FehBYF+gv0C
Qe1wnpQN+FO5MptPcQJtn7QdXac1jHcW7hGpLC1LvrnqYYp6CNkF2sAKjlRuFKaN
K8V8cC4rU1KwUg2j5aknvTIckCK0q7hCm0gEgOWsIguQufxPnTgKyJRdm/0ezJ/u
Rfeao/CVchnau+dBg51pZD2CjueWwHdam5GapLCGAiL1ZcgcqOAMfadMN9jwsjo/
KOoRYB9994dyPw4cIO8MYsg4iuKtmBkja/ZkQEO0lnePIh9pFqa2uRUZPuteFJPc
pRnbEFi38SovHWjt5ebaWh8dD7PgiUwkQrTsMTOsOenABI2DfstKrl0qNBpn9ewH
o1HBm/HJpKswfjzqebGQm1Nt+Ji7LAydSrcYVQueWPhjGtn7hW8f1QKjF/FhAkvy
6PKbT97kc+zApSMHWmbdx/CO9U1LNIkhFw5bwQCDUge4HIksi0qcwM4hKmCPI+5d
Tx0YYXOYzhfVBr+zJJ6G22YxGw/uKcUnQX+/sUDFJcLdLEl1ZVIfSgqEN+wCJVvo
mrN7xMbnBZxBAvYRHHpT+ycqlhW394ht7PW08K5GO2TUCp4b5fKlnTtJ9uiLyU52
RY/HH4CWU5DoVGEiyy6Q3EjLqlBmb8avU2ow4VihaXpQMAejMAII2rh0kBWvz9Fy
JC/e2qH8b7+mUFmS7KcH2ymbP3hPmWuSfwEsLTVqkfwlqFjKO7FeoFCc9H54beTK
yWqVeA+C54LjXpT/OWc+Z8gxuawQO6QN7uNOoBhq69JzEFWOnWlKRl/hQQ+egXhG
BNLFqpBmvF2lE7Dhx/IhGAKkOZ5JTUvn2qfTI6Vtzq5iJRg9WSFrENEFLAKxuZJO
XJj8Ri4CvBJW3699YTpHZaRanpLvxL9vQ/y84HRJIU6IehbSt8gLR5OQ0KZAtaw5
EuNHJ8h7jgqT5/VQ0ldUMEbLBJun13Tg2NirvqXYsIt+8s/ifdJBFTidjxKPHlEW
YhNgNO1sFEU8PUTh2Uk8Nu9LKT9w5l3fRf9LwmTN95XcGHGXsyiK76ER9U0f6ahz
ag1+4jdzR2oO+9Krlkw72NKz66Hd0CyEPh+2+sULuh8M+H80nr2XjnH8lEFel9Lo
HUfoi2g66ubN3427OlyvXnm7kkrmDy5OHeGDu3ipO5XDfvFMuv+GEyiV5eMi9Kq5
rKnc01e05Ze+66AFok7id46FXq6U4aZ0gkSiN9pGgdCD5uHUzhmISktajJf/IYMT
C1oZuAxq0QUv4CL6hy7I5aeF4tAsB6Sfqh4s6uAQ4bs/PhwNGP3SQ1WZzwysBlHy
KT6iXvQImBVR5rTBS/VF5WB2LPupOSVIzt6ED56eKW+pOy0mKRZwKIBI8Gyi565Z
ohvClmWoEdPKQh+X/GHckDzv+thojcvyMJD6eLrOkmI/ujOcPOU7BFMcpU8c8P1e
dHGwXqE7zD25Rh0spmyreFvzu5/yJyqTmfJgBHPXRhc3czFh3kLoIcNAucJN3Mc9
B7ub4/Vd0L5wWG/EoY8vhOoUKIjI0el7tOBCrUJteNvs/H6chd5QK9JNWgOv2M2M
WGQcJLu0mJXn0btDIbs5sO7VBh2SjgeGp0MyLn1/ySLP090BHQbB4cXAhSsbAXZu
G83F00rWEuFPLbSBwv3G1iq0uhvuOeBlNLm2bUQHJGRPSvH1lwHRMl6u1pgKUXef
fzdMwUeCJ1AYL1qahfFK3H/YtKVYdEkaMriyqpVLW27UxrYl+u+eDRIbndNSeAIA
4cGqaP7QEmiUxIT3h2V5JKIiWblHE0E2D67RxjibtrSKpKKQN4X8wn3bPalwx+iN
oe2eRMOUTiN4a/F8JHQIXbRjSQgXnuVkES9NvEwj2bBgapHs4HjarpW40i4aNC7G
TQFWfGTlqnBoSF2t2T05HdGIDSD5A8rWa+L849W9YzDPp4lHfQ/oiSWlMNBvu7vJ
Mg5zFTmn4t0LIFuDDTHVf4z2/0X7uJP4enZB0DdFGKkyalbQrsPlxBRcJLPhWEnV
axOANqbksAf9x3cfe6A2g/VadikNfLnZITf5MuII0usuIV1EvlOXHz0ly9FGHAyC
72J+CW6E4Pbbl1R4YACy+X2bhaIaao/DRgB0quUWpNQHc/20dOoKcO1pPD7ZRQwg
pXGDXfr0uB/w8HyobpV9hVX+VWWzF8K3aqOQ8N6QMIqaloz4vzD01HWV0CJINrpN
Ir72Qa4L52wvhUv9CdPCBw9huykZTUR5qdbV2dbZlIRBhddEETd4gw16wef+hm52
1/3gy/0cQ/Djd3sWzql7B0ngvCGoT140eY6+mj49VnUnzmkI+MtXWxx2e5wSiNO2
e/ltTCWLTugR8OkyMFyFUFogXKfCs1WGnfU0OPD093f/NV8Q7SG4qMxFgWEGpbQ1
MIBi/fS98UDvnPHgzP3gNh+tJDJTIWI3tyzaXU7ksg+XSwkV+71rsaQB4StEpnW/
9lowh1YmlpCXwtjZ/9IpQy3bNsNS3Zs0K6061r4hafl06f05CA3aC+8R+EQ6PiWx
pLISILoFoz74UrsoSkO48EBtlYRbRi2M4CaxJFRKxi7xQ6pbBPgJFo29i+VQ1L5o
rF6GrPSEZbB9cVXpT7bsiLSGW+s3mmIWc4/4JZcPkcRfQ41JWH47aOGxJvUH2+Hv
ARpp752p8PdSnPYm7OGQTQN0ljJsUEsLQlFiQEH0GN27vcqKfhTAge18pxgkJaGI
A2AOm3m81MfPUMC51GMCl2IgDNvhwDJhk94zXE75erNKbFT3MCX5mCSImKnqMVEM
btnb/I8EKNdEEpH3AUBhcAHjWGUYjckzpXAhXFpdjWw6Y3Rc5V/7QmR5ogtpG2z8
FYV+q9nWIjSO/vu7V0wXq0jHPO1ihM/sf6ly2ekz1LBzSTx9+rpSty8DEfDYTUTX
8izLZRYCOXaIK9bL/496CchGJIHZHObaiNx1HhzqZp0vIqQY+yuG0KgwuAZ2z1+Y
EVbh8OuTtEAAjPO6PAF8FFcScIHQjehG0EiDPqPXEuzB1hVtXROMPDLZm88tG+/k
IBB/IKzW7YNBVr6P2qUkaMjjB17d2ackD7Hm8DvrYgg3XGkzCMrWtLG+VAmfjLhm
EInoxLcXzsaxBx2UwWdtHHPopHT1jDkE/2w+iwXkWIUlbuspemIUYwyBivH10xH3
3T0zyyx6Auypf/4Se/CyuxNQD8mre8vBAYAdT4ws4hHcCz9A4Vxf1Oy/Xt2h1h1U
6mztJ0YJz7IyLAZ6AeFoJqycKDxLGSwKRkVteQvINzCK2PjJ7GrvDRSSnbcrAimB
oP3fBOcdpV+2HmB7z4r4jQcouWJh8eCzoTb0mWscR2Cxw0GzeA+OQHNV/1TrCYd3
S+TpfLcAgNihdsGl1EOV8+55AefrPp2EPpX2h9T4pkcqdg/XyoPIjgRqKc0djej2
wqGugOr/TjKIJaWrY73jqzRW8a+zA8vE8s58ZxwW/UJIdUfLXOOOaiIOorE3tD18
4slEKQ+pIhCMOewqiFwRHI/bO9pZxJdfgPRUPOaBLN3RS2bgnMIkYlgD6tQq1WBl
IkpLeQiTBfkfF6/UqAMB3ivUf3OCqYw5J0TV67FDyTmpZf3yoV3E+PUO+1oY2abr
SWLpbkkT/H4XZdMkQcC2mHeDsWv7D3WL0/lZbzVmtVP2/IPJbr+BBBmexFEqYCjG
fYZvzbWKWsIJNYS+6qYKtQIgGmWiXfNWfDDRIEuAoQ1E0665HkMI9hPrsYvF7xdo
M3Igvv05uug3SyspF1/1mGCYKbMjRaTRrpOXevylsbzXzDLiMAnDzb7asIjLWhMs
dpqFEc+dzlA1K3bszHooBCy9XAbdIy30TwnkEVvNMS0Hj5YF0COdXwDtF96cFuKe
E2K7hWdOJf9snIrAbJUIYDkjDhqSolpTqe7ITsL/wEPR3EOkkGpDH8Si0pBfsbzt
lGxYW1/VRaFOLnKOpRJcC2mvUIoYsFQlC0l1/Tl4mhFFSjQxDV7njTw3qlCIcuWn
Q2BF7fdeYCOV8T6G7AV71U29dtzuRkbNapZUUdcqTfUHDp0AVgUbyZoR7uk91jyo
vXOn4azmPpFvhGTfbB2A6+kmUvNxuxVPYkddODWibuynmPtc6ksMM+7xNcxGIP/O
9yKAIZ2Vx2Hu9U/KiXRmz1eVu7gCoOR0fjlENsz+54pw1FF86bXl+d7TiR1GR/pA
xLBfzWLWYB+3tHSkBjZHujwqd1mOd+NMthYEHC90KaRkKErxfad33ZWj1MEMqGRE
Wh5pon7VnUoprcG5FQpD2DsW43CMCDimBVguMSnyic41o7sLLVtaOmfsBwL4aNSV
IxkvGkGDPtyi744VmJs8AWutt3e4QTmkuQsRKJUhwdJBUmEzBEQYEr3htwVgEWhP
nSZfFcz37M0w0jBYxLxJEqz2HnOYSPDaekYRAklzd7b4RdvF/Mnz2n5eU+O2Gy4Y
1KwtN+RtZYmiQpWinwM83MBBAV6BF1nZsRHkSxAOqbBMrZG1Zp5CnbxhlJRzbJ7T
60UtdTrPY84uoP8vZuyDJrF9higICe8v0GGIXaveMX7WVLglPF7klsnEVE0dUxrh
NdLrNzN+1PjSa9aLBJfbBqMSqQ3a4AJ3yrAg1knjMVSw1iztGGpPzSTsdUyHenDV
mTZNnxn2Xue7+GhyFViBc99SENLDEmfxbvBMm+1WhDB6SWnx/vfl7P0eM3WUBHOE
9WzOv+5hfgcwVZT5cvXYrBL3nlN9g0UgdtXvKglg8Q2nrl/xJOCr52jbwByvN3pB
6w/q3V6QMd6Wdzij7Qo6XTzs0NOSUk719t0wjGYEVTN/z8hUJ6H6MXWp4drmkhYx
IUtLw8gO3QbbsSp0T/wK5obrD8nRFP/OV0eu9vCQ51k8pxJm4ifeo7OWQ3g/rN9S
In5rRb97/fgJYde1fDOLCwhMEwJyJdwZEOpHvvQy4NmuapSWYJvrwpOLrVl3TpJu
uPcNR0bkXueWtEqRrHoWIX5pEPa2k+CUVUGtAkKxJXjGk4UjGqxYTUfYC/tpEDPA
dx3in35b7LHFIuHAKqAw2UxcTOvjI0FuuRDIAWRgJ2WlG7smxvMLaok90a/G6T6A
tXttKNiT+FknRHisjNzLQW2YNvQ4rVh8w0nTzvu6yNH+mfafi6mxn++CgAEuLGMN
ClmhVT4EQwpNYmMDbvHr8OGMavTveEGWCRyIZAe29+Jlw1N5/MOPlCwfSxtO20cO
cmvSrLRJqJdEk2FbY6Sua+chG/eiXzoorMisflj2NsIkxLegqLSpDiyUYdKIk7sU
YFh3KAXFsFueX/tUIJBCQhnV9hzNNctP7ATbxsQJtZX6eGGhNUuf7UBnZpVcfQ1s
uiL8oZ+UDp0bqlzE1/VhWK1qHBFi6lJGnzp5nx30al0GilrRiivhN1ga7q6MzX2H
C+PVe+JemI5LER4OVYWCda4XtichLxsge3XK2g5kfOmWPm0VAz6xjFXWgRihu5x4
GI3jEeCoOFK9CkMoFX3acpfu4ZskVKo8wRS0UGuR7gH3B93aQcvO7fcivSc/vDUl
iGcYIZKHxS3dFCeZCt8Wt7pvLe28dXKfAgChl2sP/8h57gP4XOzPy+Y/2jtHvwl1
S2kp3J6I25kdA9x+jKNhSEka2Z2LxI6v6o48Mn22+PpRVfMhxqphduqh7Ei65O4m
P9OunGt5LGCtzJDZHWzLcR8E0tJK5zkFSzk8/iyBfL2IAs/5adUwDFUq3C6DFypt
d4BG3jkf/ssE/UxfsmzekYfVQAi5iLL/Z7mjNM0F03lqHJnNeFrlQauTBPTGb4Pk
8LQ4/CW7V1JSrfOCvPNhlyZzcLzBBFnhikHyltnK1UK4yLx05TXKAvtai6nWFWvK
t6iqR9/VGMwS1/Mbdsj3EL97kvIGRsQEBE3JdvDx4xSvLIKi230EfJSp8YJ4+hoV
p/Fk8/HrGKPiznvQGemlfpL2Zp0C2kj7dx8s9xwOUocHj7I1Etrae+iO41DQ5V4t
Bpi09zmdfe8WVlN7QSmCChrXo24uh8lz4pdJx7Z1xL7w7O7qs9QS3MYfS/Y0Jr7h
svUrctPQ9rlZRwz3C2u+zhz0D3Ddd1Trp5k+1a5UozFjqbLpjPJ77sVv3wlbwsgB
ce1lZWHluUbMYYErrlkMDnYIQYK9M1DilUIozt3G7SdowzuEJcMqzHpleXQzGTN/
GGjN5JUaYeEtE+uz4xEL85csvwR36mPugUO9147OVOLTqUIVOIvImelOx3vfIj02
WWkoG+jdP1CQgwon12QE5PIQGbfUzIYwPUwdtP3m0eqLnRNXTO7C7BErzcFlr7pL
3SgnECX0XN2YZM9Pa8n4n6a0gglrXYLSkrC16ei/brYMsOSdHa9REohYG4Wznf3h
zrd/0ji8sMcqp6zcAKliVKpM9Osq3f0hQJ64rMSjdLBZ9lm1hcZvlIR7LADz6dFr
7QJwXNZtSjjQfmsoDT5pmju+rkJX1q8JJYs85tHV8DfljkqIuriyk7vZg+2JcdJz
Z8P+hBDDUrvRc9GJj8vtXA7CIoVJi/u30ge/U3NeLrErD+HwpGn2QGGJb+7xLgm6
+QLv1fez0EWaoUePKpjOgw46ippK/0yryVxUmOS5CMDwWnfG67y9Ct8MM+7AnOiL
poO3a39Pokve32JqWIwJkMPIaYvzRBQKryKRRF9wFA7jAozW5quQi9oX6KblNxk+
AbhDdvfO2y1WG3Kgm6pTImk8Opz3M3nYTPQl3ut6t0P+MUUPsdDCLwqVyGly37A9
AjyG7BOjJOvtsbNVQ8NOaSkMYClY+3xYUxMgSosMPQPuDiKkra477ViNIhl9vNgi
ADwqE13X2W4T8V4JQNmer78aHtHU6xN53GOTKHMF0NCPDei387xReR8XwnGujXcb
ZCL2wO8UnxDUyIJwawkDXWUSD9PcKM0Hwnm0xdK5SjLGK2vgoRcbrXWhusSSxYct
baUGBeZVTVdsNk4Xw/hR+0IPZPd6dWDhnqyzw94eC85QkudSTw9N3lP4IFhy2opz
uif3tE9mdVRfaQO5Ln8Cn+NUG/vYMuPnHWfbaDm4BVrHvEcS2vMalysA3lnAhK/2
RVC2klH/PQjpzmW396zXys/aLSKNLAXFpN/bRWofJPdksL9lhzGnmjEPR/Nb6iVL
3nrGOE82ED0Rv1yClmOJ80hqM9+JGievSU8lAN/q5+qHixwTOXAr1Gcl5O4+auHG
nF4KWuTfULiAKnj9Npk3J8QDoIFKsXgjnYQmMdivG2Rs5q1GxCYTPAHwNuqDqEp6
/t/EeNtpjbIlcFTT0LO2xcxmZ4zvxupxZUdWFEIVNCRnIFf/XdKGBL7Z/Y6rWx1B
OiPE4+LLkCK6eiAWe7eRWDRuqLKqEDoCzCmtmFKmDljYLgewtaNGcJboQqPlxO9Q
ZVwSv7NZma5pklF0pLXU5aovsKLz+anp9ggTOPMva1Bv+H0Mee1r94QHmtq9yk3c
z/45Bj4mRhHfjFfwyPZmgMS+A233ey04C3Ib9AL6eUtSeIgrcA0HGN40xa26BlaH
jxhnoMjXi3jbcqmNeFL6YCozYSNUX2o6oADe/fxp58M/1lJAxQX7E6sxHnfROFfD
sYk/6EBxKcta8wh51dyHisvPlUSMXl9Ol13zGWiSqYyj61vO7MXmv6jYLCXPtUHd
cGkGmmu+vTWYdMaxcehiaCSwHG75eFff06JUsV/ATYiNVFhAiOeDtOec55kT9Tfe
s6ZdBpOBBgU5cE5NdlwaQUSqMSze82YFXC8F8yV/Kz8dUQ7KUiMPgU7VvfRa5SDY
Tz8piB55Zu591uu/BCtMnB37k5THR0FTH0NRU8b/pk99gyVKWa6qODBdNzSmrP8Q
S7ED4HGFH7EzG0WnfL+O0mx3RDCwr2mF1H8o9c6qv093BMqiW7U0s2C0+9YsGX3/
ppISpLEskraxbHzL6UVnxq5cYGWe8lzralm6Ug+qjQXB+0na09FY6kk3xOdolgV5
u8qzDbyqLFTK0X9ykHhGc+w8rdqUnk4PhS9kn8zBcVNzlh0Rvygw9/cHcUjK1UWl
aNhJdabY6UbssXqQhfihtl79hhVDSbZwW6hYlq0H1pWrOvljI8kEdShVUoBmj3PJ
95cZ/iPaRq8RBSspwUhC19josH20r6vTYqzFFVeSkqKyCgLcsKrImcjyH+tQc34F
b8CJl3ZFgEbWQFuMI2CyBLJvvXC++Ciwqir83KtGu52eAa5PcGurnzTcIrz84Kxx
BusQ8Zz7Ky8lXTkdTQ9V7kWW22KTKeG7He2faWWIgNJrhuz1Gv10YleV2zVAN1tI
SeSVYIeDRq0T015LKibL0PAt3cUN5jpPiP/PJgS5/ZnHBfJVEXFz5PTgSMpaRKef
FAnJiTzXhkZNAbAc6ipq8AcAgODASmvTtQ1cbujXSwhFg2KC5qpmKHzVg347qAOy
dKfCaZbUtaLUrUsTTPpxFa+vNRqyn0JeZ9kfqJ5VFduvW/eTp1oAmv0dL8VvToc4
INbGi1WogGq5ZaSbjp1Os40YJ746LHDNBx1Zwlhp9Pd6i6AT941mS0i/GYbrTlW+
alYml51+TeB8ViWTp6uxBYrPWbHixbiShT8HJWYe5zOo9NK8UUnCQ0g/fG4EMHxJ
a2WvaGGQM+MS+9pwMF69RxeQSO16tfeAzfY7d9Z82sdeOLHAG706m/0qCIeEfXr6
lvY5udtcHE6fCvLUfjgjm990LV+44CJjsyhcm8gOcD9xb0B+fP3xti1/eE9Ik57h
QcvdL+TX+y+ShNWJw6/HBKy1QjzqoM2OaJJxmqmC1fRqJ3nFO8k5qsJ+OxkUiP6B
IhJso37mEldElno2LrYownn/nRlLvfJZxukVBVNZ1URdMAj2C2eALcoYAgXjhgUv
WItb6clvvvRiqZH3uEU1ylKSGGCcBEG58CX3nWx8X9yIzvqA4DpDKvjiEbEcc36D
qO4OL3iYJreW+WRuCiBTBarf54jN5sO77G3yBHR5hc+sRDDvnAnOxxMLk+ak5Mwl
Y4S4Thc3OeC1SBEKKVybylb8q5jVOXiuW/aitW71zBwLgkE87Q8NBFYIO7/GpOX8
gSILRSkkNPbF0lxxSgwS+CjDwIDOVRIYLiquiLguyHJTP5dCAvpWihBK0omC3Td2
ZT6nFQE62r4YrL1LrTEYLO0w/8Ga5rBMtgnXml64pbticTrAzE6gGioIoYaL2jCX
fkVacj1FG1Wo2ITDUA53xr738/lP2qRrTH+yhP1BAgK/FtMh+pP+LNxhOgALA4oB
Wiy3VIod8h5/WhKBPlZP7Ma29RU8kP5Wir+RQO+p8Wz0Yo35QhfQ13xHXI6Jros8
Pfs5KJXoky8DL3b0AWFqMvZlKPWCm9AiOhtrpgqDNIjKL10Abwez7RKIjwIAqBXx
44JR8hcSksoJbDDEn6HlAGNxmvbiSRMkqfpU6RVYy5OUZ7QB4FwsjUxta6blBmzB
w4gDQ2NJSRvYVc7GTZBq/BKuw/Nwnke5UlO5+oPmQut+yCXonX/KfQ4gjf+cSdoH
rv1Uzm8SPYEsk1RF7j5KNX2qmqC0JbV16nZyngIcqkFOiqrXPHB1+Je4GkYaDjp6
HdQAUw5P88Pj0BxCQq1JigmrNeSh88ZIzVxZD5dMqx6TKgRtaSWv6kRHH0iTKwqV
YRSeteib/r0JrFSkKOfHOYhPpla8PRM8j9PEF3GoWAKF9UcBgv2BLa7Z8AZ3okJ0
IY0brHb5xDeai+PFay1bBIliZiYY/hrdw0hWmW8WA6SHjft0Wli6+uwozumXoogb
5Xycs7tXMK68Hzu03TlscbMB2pKWZtUHjxtE2HNmYdb+H4H55mRvAU15hiMVVURP
DJnhaw94/KnkTmH0mV7+aC4CfGlcxREzkzCha2nsHYfAy8Iql/L8ZO//iqxRq2AM
+YopjokdKbH7rRer9zR+YM28hbi8Hwjoi2IlxhBprFjaKniTC+JDZoqhN0SsfUpM
iYX7RrwKJNdE1G12lmzLq6R/6dX9tGzyrJHB6k14H9bznhr++n54uSnZGuGf3eD/
TAUkZ7Ymp2XKxfSgyQfCtn3CnQCJnnQwMnB8uaYBGEpuWMppLqX09vYPfkEOajoR
o/FwYAyaVq4Sb7iWpClUOZiE1bLAryKyFs37tJ024gCrIzQM9zRSu02vMaAMXoEw
ttFzSRbZq74r/xQsazbFY5rWpldRUpUMbdFAIzCLhMTxAmR1ihikhfRqVuQlAIoA
WrY1TaAMKcyJqVwjmJnJah13D94oY51yBIQBtM872rUF9pA7eUEPJIt9w7tpjedJ
bNKyrahWltO94tp48HnhqzLy62ER71J2R5RXO3Pk2HjTImbkaq+kv6tvypUzCmiX
tCD9/Z2toxBDme1JvbUfHKY1DhmWUxdg5X82rgI9/OHZ9DiKI3crC2rcMZnF3RSJ
aFX3VASvb3IjtQNVLoNRMFRX4n+oV46hl3EDDzSfdxmy5MJ7qk/wt/nokyyPhS6M
Gp/tA+JdJG8mulj5MeBPBR8BI4E5vH/8r/J/6pCetQW1LJ+op2iN1E7v+hOV6Ubt
EbNj89E3bEjz92qVYKrljrlA207CGXjPy/nHy1qYeSjxdJo2vTAkBdYVkk+6cbUE
/WskBgfsnOqoTs9jjcHeWIR7YAazHo+XYKdzVMfLy+2KntBRj/cUcuQ3tIF/kj2D
fUJ0bBdLWux93VTpiuVIOR+u+7ok0d6xzsIiSX4jcLVHJUTbrrshOnHv/gT0PJBv
/QUBJI+qW/ihLulrTmPptlCilYbhss3RSIyLhxUsQdGBo2zg1Cs3KtNS/padFHpI
zXEgy6yMgdH0D9YkQZKHWO/+1fQ/UreK/PC1To31mGBu5pBIGHF8fQe+WmDDU1OX
NRHjGD7C5wZMIlgblvPoHlOsypuU/rs4TN9fz20bRGQkTvBTIKfegWZHW2p5k+r9
YTlHk+R4Qy/FA2GqKFI2IqIpMRGc3QbtX89n7nwi2O5gzg64GPCqpmRX5mGqnd0h
Xk6vUjGRbbRrGnYQXaq8z3A4n4CTOQeViy458ytJIgJOYDeXq4JL9pPovtuAra6/
ZogizZMO6v/IoVnUE5vLyhbJO3OVrgDbbkGEAa0c+K1VsDGGzT8LGpXucvoAHOhF
9eeffaW6iyycQOYfGfomNUinMQhITFA0xUaSU5do5lyXDI/eFhfOEncLvytePsdM
ULfQ5m5G4QX45dtntBQtKLyoVYyv3/T7RLvRRqm44c7Z9oLiX4dAYiSFlozbKzYE
5/HaCbWTtApX7CWQ4sEi8FN23xxMaC3MxXLg+N2Jth+zEBETD1CjP+8C/KIX8GDa
tRgrhaDLEXQ0Y+EbEws2mq/Bp2g0OnPl0QTOUKkg1FuEMfsgRiyGxQIyKTVEcIPv
8xPo5M2sWQ8xpqa0ekKIn6xNQ69L1zF1B65PHIa4ZY+Ru+xsu5gPyFZuAUmMoD7X
bm3dtltPmg0cCH2f0YEFdiZ8FPMTvHsIUy8o0MNyRp/NkZqynB5DkW2stcqtV4Is
3xU2XI6YkYcYINpLSucCwIKfZFp335zI4bBc2zY9uTlQb7I6lYflhI6Fl8p87ChK
LYKGWi9DIwry3R+vApWOhhbXkpsyZ44FrABW66k7yV/UHdcjOS5vs8xOhm09Fzni
1IJ+USg1aOQjd8xtcsgaC4JgEPxAsbydPI/PpIFCztgUabDOX5bubfzy2BIqXiLr
V21pE6/+vokU4EmggqI/IJddo45YDnolHhj144c2LnYmHagC8+nv9iL4KMMTQERp
DGbeBlFsIgPK58ZHnci1/vy4c2Vq2ETwoZsVqTKwKzV+Ifte4FWVSiIq/0q74eRU
yiHmNhgxXoNk/ap3eWcyYWejlgx+AI+NRlnpfBtDVpm0BGbbYXZ9BfioM252elKs
HBCRCPCp/gdgh/eYp/XazGqUGonMcXVLVZO3BSNjwtY71WwrAtQXXGqbDnoFu5dZ
n2YHgiOfxqzjiR6rFsEgVm3ISkzJ3Cz7l9mv6uLRsMkl99gVdUnzJyFRiVpq6kjV
iWh89T9iqNLFMWL+B/wiCs44PKI75X9aSrzMYfrm+aQARWKdn0SINiYn+53fbmu7
BbN60CfM94ZFatw2JmPkiukzOt9w3FBLW/b8TydUHrL0ccbJB1NPEQMlUt4oNkOx
kOtiVw3tfX1ZDVEjO7opWKChicDISM913j6OrPKQ/7p4e2FHrjOD25tIyfVF1QTG
YIz52r3aZzp5nYQeRTkbf6W1OB64U6YsEpKviGeh+wZyT7QY+SIochQ8Vy9Kr8gn
W0zEc1vrdg3XfjQP0SjzIH04HYzL7LhmN6XA+rNwR3zCgMyDhUlqYb2W3eSPmhIj
rGQSk1ywHJao50vKOWvX9Tv6GGGeuc4Mc3s1IR0jjEWHMYsEpjJGJ+tBLSf00msY
7BU5RnUW0EfYgK1hvtmIokiE9+tP1wqbm17/CzWPCwBO5cIXhS09zWVsLKw6afwB
aV8nEs8nQLlqiFaxXAlvW9ljujypxh23NkbPGswByYWaBjiyXMKdOttxQlLIHFwd
nZR77q4AkmjTf3HZ6As5RDwKlLzZiIpztLXmGMi3G/kLIBHOkr85YdkvZOfCQMQY
dKgz+Lr8lQpCdFqTwQS2SN18tlOlyRV5Bl17tX5/gnmDnx3aFhAe56zQL1tNk7rY
AeXpbnka8rIm5KiXGuYF7/Du/xzIpcICuebV0VghayzT0jImLlGjih1rofZi0xRg
FfAYeNLFU1SHQY+/TxooDWZA9nPTwF5Eo+V5QVTgwk5tMbfG69n8SwPF8L6jmnMZ
t8Oih2bU0SStokwhbC2oBY6x+5CYcQKmEXhthUJHyfvcGTvRi4ivro3qT8QarJIO
eus7J5WZHuM9A3t6Az2wznZbgsIjJGriGcvHXrOWnLnCS4zNmYMxctEnabb0hwyg
IK/W8TxU1PvkOE+obOXebZbaZU9bR77nvRPdZ/UMdoPCK2MjgqkV9LgUiHVYUaiS
6MUzX2Ck1sdJRJSCnMH8EprifVOjxPV0jCJTUVRrCJoWg38tPjbpzcUpkBy5xTZ2
nzA7Rg3cu2YpMJkN2P3Pb8wcfCYg1V7/UdLTCVXI3s/nbT/2EIfMM/djQqlgeDpM
/Gt9O+2jhBuYcjNwfiyuKQNt8fBNe84MvdmBTQdnW+XrFhJlYpB4xAGk14de4e2L
iMPUps6PxrBat+rEdXZpVF0d8vYru27WTCt1eEF0xh/nNkknEzqpEIN1nlMNWjui
O3y7/bmlPelia4L4AD8rXYFMNOvG0H+27sKJfZCXFl6QxvlTpDY5GpfkBEW/d1P8
Q7TqMt1EqduSf8/ob5GKkE9SOQt5oYQ4gvefqJ9KDQxDyR3YfdMCg9NLa9CZwtuQ
qyaOOFhYcbeVV+6fENOLpx6qaKhkzjX8B7zW4I2lc8yABMbk5E1Et901jkKKChZK
LflYne4bTKRpoU2hQWPg/HPcCLHiHnR7U+tScNyyuK3Vlvo5LesLok97EpzHNINv
42VhWB7lucU6cZ9Jya82Uly8KDMHJqIo+PTWlSScDHV4Qe0/dPa0f2mGAS56XqFC
c8aL9eKPEmxwrvuAoLuc8Z8hOF9f2e9JrCtWkqAKyqRlyldv+tveQ/zY6TA/JFhN
fXYAualQb996nnoXNo8w8fQucvbWarvPNZ3TynysCI4va17YM9BQjGZTEAEbkW1T
4tYcBvQ8D68ihVoCCdjAzqRM0JcHDOeASPoirDN5ONFpjSNHHrmywNgD/LIIJ0Qu
Q+2kNuusiAIwfqoz2sMXSqk0jkJ7tyG/L1D531sDjOwMrD1ZSzVo6+5VHomRaBSZ
OUwiNwgeawrDOtOiEYk9gZcFC/WLdr+trQ+j48zbfKZHPGsPKXV5/zMfRWq+rfR6
dxq0Fqlo2MCXvaMM8AX9thj/tMtV4YF6COlZ+OxE5q7dsmjOrnrJaiMiXoRn3G0G
Tzks7clALg2kEIdBgZO6Km/LYhHmPJI648pmHOSeiBytiW47GDdeUHiycgt5igPP
G4oc2seEwdjrMjUwFkWNEgJ/5gQSQ8SGD/Hpi3HM7Ia9fZ0QTsXoizHIFf5GRFDU
8QPa3f/Bk+W52dfPen26LJoESvy57I7+6TyDYtJu61DtcemQkIXsFPYhhYFjJ/mA
WZYs5yHv9HTIA0Mhl2sJump9CmPE7Px19nK2rdKipGPJIQkEv/m6z8ofso9Ho9su
9waVupcbpswXvExTmETGFtPex9pVLpHfZIVReNorLBejCjMbGCGBStRsCVdP/fFR
Z3VLlcbMRySgD+GKV+OzYq4jWECGBG1KLyay1cnD+oPKzCdoXhp00rzwWxAEmqAv
LKkzpqCBmJgIa3sK0FOApJ5e2xgY7XERD5IGqxWeNVeDChed39CB5pCej3J+oaCX
eNcFN/J8Z20UbJBCyawP8HyLOhZrGLIj3BxlBJMWy/8XGXTSOowLI6KJi/XWLMsS
rSLrV7DUaMJihp5qlyURU7dbn8G0TfC4lApEeUNnvieq6lB3J/uKr/tN9FvKnptf
fWndyqnWyMf5rVrYIM+bElTvSus2drHUclM5I6hcrh+vMkD5DKDHXVGkI9KeRB2o
p8uwK/6tazVEM+U5q4M/+w7+9Gq5KE11w+lwbI9ZlYhr8vZy2ch83WMcHoPp2IzP
TS0UqnAYvmi3q9lKMgANtbYTOzf7H9smwgiSfTtMLWiZcWZ9qD3UoR9+mn3hDOLS
Imj3ymQhhrGpYOkdhFMrWKGQy+3uiCzbpfKoXC1YaoYJAmywmRDO4bLqkhL1ocE8
Am2XiPoggYG0i4JnUva8D/iWqKXM2TFw70DTNT4/NQuxzb6i58ED7Op0iORXS4ap
LN3KmqEXiULV5QtMBY6kvaI8KNIUMtBHGjUKvtj5s8IDQPnVZ4Zh9qgAYbQ6NW1i
54quvO1x/9Lk3BXjIGR29PwJMg6mzBuXPSF3CfwXliaV9lkm/KC0PECo38u28F0h
Wzl8qGM7fS1puOtchkdXbIuovCdSLA5MsWx7LfVNewd+2VaL9/JmtALNOjuDxmqg
u67JaoS4xhz0ucEHeTPa6gSi5ETJqiI9GczVHT2cbnPtqxJXFYz82v5Pqrp2+W1H
JkH0Ru9ttoZWf/AS5+yYkADCMpo/uD4PA/y0lzxMNn1n77M/jkHDlfYeHWX01Ga9
8O3g+HAyiOzo0TLEc9kIhebHl5k/Rr4gM4mlpbHLGNwKZJQfyUBDmB3eHjfViq94
ZnApP72MTR2pzlJ80ne+le3ChRD3CTleNoKubJTMwPWhyn8Xa994QFneVSTqTucL
dd6bSKXPJH9WdkRpla6hiBDnroAqqXEtD1S7Be0PGJi7IjrV6e9AyWYrVhVlk2y2
F7Ga26xOWX8SSZImgaYsA4KYxk8JwIfVFBo9m8OZWyQgjeeXhb9RUd6C3AYL+s9Z
4Kw5PEsbD6z09liYcw4o1SnqF/67aEciY6aI0t+cBTq40psESENkt+mkWClhdbpe
KFPZ4dWri5EMkVqZ1O0pwA6xKm68gHRVNcqrv4MJXxqVEnKVUVOOqCTBOVhLIBXL
u9d6Y2Mv1HtgTe7fpk+hHOdbCQySBEO8UFiS1viuhvZBrHrafpYM7qXHUgCp5LPk
zhBb7lldZFI7ZJ4DuAGaFwgFPZE5QY4f+S/VN3t7LiKr0CBUZZEBYfQV06OvM6c5
/i7cqTMQe50kRpcTLlBZ5MdllH+32tIB1geRqYSfMwGkX89Cx/W9yu762lrdVw5m
bTFaeiwlgBZxUzMnV42/sHeRggFpJDRTn5wAhXpThwDmzFs4/5srKIZ+fJ2JjD1+
wHlRbJZMoCc/+Lc1w/GSKlh6ub/4qKyLrUSYVI8UG4xODR9VCsdpUHN55QEcq4Oy
WqyIxClq9RMH4QsOQcaH0ONN1HLFPuQtiLpneWCv/FO3yKbg6dqp2BiWU6wxb/RO
Q1Oi1J2zIHpRE6eBhEpAZ0YU+ZQ9AVtkHVjv8JsIWiGP5NyFA7lZXJm08ovZNKWQ
y2CmIAgB/coNM1YelrWIlrl1Geg65hXFL6anjQJKJq3EG/u/9cHxvSlXLM+KYDWj
tZxkcKXOu3VJciwF16ZOzrXkjf9aoc9C9WRjVsiqMn12RE9NvZViS1IkPGd/3s9z
0HdHBCfNRGkGotH0T5wnXkn8VDIYzjmH/cwZtWf8oQ3AH2IJyYzWm+vHx0lPnvU2
pFCfrwwrP4dSHlt+pA5uvab1WDjk1l/0XBnwrbKFVrv+VlW4ztD0rewojB3yUy2G
HMbQHJq42izqXDx+XbH2xSL2bHsiQRRX0JTDiwsZ+r4H1BGZBhy2xqO3nxRBYvRQ
/Pgkv6YVoSsAQ9ZdNQlEBQVkKiPWLo6be3KBlzboyNHeKagPTL0XvxlPNSI7nTyq
NOJq1P787nqXNtLb91WS5nNfg4JBkA3GFJE63EO+mUY2Jcp8a/lTBRkOIR3Ryg3C
Vd3EoA0BEYOw4li5VyXvcD9UQ5ep9CPKLaM3huPn5HFsT2BYLiWZnaJdcrH/3UeV
4XSTaqs6h9tjNRnBq4MjlluPR5uJYBShaSzG/SDLeG7bzWzB32+KpNBLuVj3Nr+e
xrBDtovcWuznNSyx3k/IQwOfGjA13VFKb9HXgHojTCCiHaENckR73flFX/9uwJZ4
dVg1KFkOgdo5lzUpDK00hdI4BM9KYAUy0y9fFig8OhMhSliDdFxDwl9zomS6fty6
ELu5Ur0FWO54+Bv6J3XBr+xCBqZkhBuoSiw5adSCRNgIiwKuRbaLe8DhQd1BOQvt
mKqhYo7Lvw+FdhdGnAIfmHCpMx3FcYCYdTACk0It3zDhWWEZ+HnjzDhky5KIr5TF
ZCRan8tap7vTFp8QnsX3lUG6hvzG0NbXzYSunyqbXwz4XqZFQID2KS5nDfQW1vDT
obHWx6EqZtZmPbWyHNnx+3cw1nuMQSLokn1wf4Bjq/79c8WVZmsN4gj1LU13JQl7
o9jE9K89wVUUkmaWiXO0uLN7pltTt8Aguw2ena9POWN2yidpaNrpFa5u/gh0MOYW
prB0itm8IwKxSYN0ERGan8yG1i4sJhOaqrq5Vb8zLFPNtsEG3DnRS2gUMxIsba6b
x2TtbAIAfPvbW+GjxhJ5iAccsYlKfIcl0saF/m0umjUoJ19bTyIWmITJOtne1+gr
Jj+5vBmTCbj2YapDZKAgULlV+1HRSLlJHtaHKLEqQxpVqwKrKx7fvHseZ3G8zupo
6d/MCBMuSd3It9Q8Tpwsa1v6DxsbwIOeGSY81sjT8Q9VuI+s8ijsmFyimZzjfBFN
DvZV1/fZIKzGuJ8ho/Kltg2XghKjXGHHqgWpwS6SUOdAOKwtN9p1Mn9kbn2uFL8n
3cBq16I87hmxqseiTmKNbxzZcVOz9MkSzyZidZnDFjlgE3wjWc+KTak4wOv5JLHi
hF+WBpwlR+M7qFB6MfclIDCbXruJfsLFBSwIQ4/3n2nxxltDWKNBjvCB0hZxDpgD
h1WMt0sUPqNbvgRAgNzUfpTqteubioQTOFuyqF6ZnA8Ijpz8H14aUAgpECEsj7/F
G6H+L5GkRPEGHk4qcQz3ydlmzqgB5tXLVqtvjeRHCsttumwqS7Jat04UtZlF83O1
rR4FqURkANo+rfBksr73XdhU2+N+OvZWe0tVjnr27vkBS551fIxF700EBQAQmECR
6b8yNO/EcUybhjrzCi36Se8MLs0eXxeQ5kFsnkDal9XU5I5F5IvVs/tt0XuS5WAB
F4mtVTMNQm8BixCDd/B66i3q35qGZn8MAyElf2CR0ZI176oQI5qasI51ld0RjeCc
c14rDAC5zhZr72u9UuCCTrtX2JvAOgYzGBbpDbjml0RmDlGBVZ/XeKvgDpDFVvSt
WPNORhAbqcSRn7+F1kZZv1IfzGE8aQZwe9kz4N4ePU153Ug/JOoMcRb+wysmOxrq
XLA2DkTME9VWhYZFUwVFwi2akQT5LVr6ruRJe+bSClIvHau42z4GyouVopZlpHLX
9RmspbyB7rw31U8hF8i5Rp+G8flgX9LwPBJVV3ALqYLAIl8JRIobb1bwEQMl3Zqb
qZSd36frQoHIRXiL4eB3DGea/4CziZVofeuulI5sSjT17JJRIhMfx+p3kx4qMrCs
90b7hVwhy0fduuBA7fxOcluAi26yVjaU8C3i/XRDrz2TKQrLGCAjRBibq3IoxSwp
MxZsBQ6tnTt9Otdkj/nBmeiUqOSvFR4un+wRPNslsUAFE440PC5KF/rll+z/3qsz
AhuPwItFojRGPbNXLcDxZSkHnPesrx/OSl40/Xmql2AVmZlqpke3WzV2r1XUAkxV
/O8yREG40XVNoNQkc8JeP5EEWecBCZCeR+sr5H5avokoGWNy04Qmz0UrNO3Kon7C
+e3B0w9rvyDnjV59zYRcUIKCwZAn/Md0/68LDGhNZ3iqJ6wafqETK5TAKnwdUK9d
DEI6U9ye5dHXMJodwD1bL+a04SCOgrfSYVUmYF1w/qaxFn5pgm8qy2Wb2vUOsd+P
yAL4aSyvQMc2FOnN1+9NKgWXD+5aoelerR9001dGz2xoRwGMdIFBvKszWCoIe6YN
kwKqeu2sdzwt7pifhZod6yr3bIWxX46iW44AwOGJqqBewNgpHaWFFnr5ZGDUNCDp
vB097mN9E1kvR0tFjvQ66Xp2JrkptaPqAi21GEH44DW2VtDce5OZ+6Joha0SObbY
G9bHsUhdlbxB3jUtue3Tm3E2ih+z63AGWkTKr0wmpD8zXq6DUyOAoCSN2jxwDf+P
PSfsQLGQyb3lSbK1hIjOPrliAYEFziNz2k1za+CJfZe8a514gBg53t8u2wIt4X3p
7BdeqfcUVO1rJ78CFJng7to6GQyakvHn51PiQVV8U2mWH8os23SsSqp2S20EiqH0
i5OwwFW6KOBXCRkBO0m25WLviBhQgX17OfTOo+tqnpM3qCOL3NNDWhA0WuCb3Y7m
I3rv34IPkyB7BVnJzvkxeg6lC9LwhQXjeWbril5NXLtwL2mpfgEPMJzCqur3e0T6
tjNOCdfZNA6fVP++2XLPu3zTyuLmS7/YwpEhGfOJC9SwGdnSeS3g+diukyj4pjbz
qrdfG7ktRq0CZ2DoNPfS5ESlvNBpUdJYQLqTliOaAmivXQ4Dqk12Bti8shEj7OHG
acHttMq69X3wClbKu7/aY6Ytmmt4MM6flGqCU5tw8ZgtyKZTxJ2busXZRxKQqJK/
WiIg2NeHZhU/b7lzOM6tr7nYAbw3J5pt0lQbvbg2+j/xCFRKxavCE01tr5yzPcHC
68CMd6cGUPfzNse/h22xQr0yJicG7/mxV8CSV3pskmQEdVTJztCyrJytHhq+bHyq
QPygBYOaZwHSdbxRxnxkwBjJzKJrYv0RO1hiBUEjC0BHviDJj5b4nH2dG4UCXaEH
DmKYc/9igJTF+D2UTOYmlhNiyT2wtEMtQLRQfFVtAkHNsKLS4cI8YArNsQxhxSbQ
KtEyJMFVE57kXQLQ0lie3eIyJuLQfH9lppy6Q/ZhskZowXXsbrPAE17nrn5MA8qO
tTI3m8x22OJSNfumJvLYtdBKI8LS7jYmNXXRd34OCEgARVAhTF2oONHVjBnWh0+E
`pragma protect end_protected
