// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 13:57:48 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
EOANbClqtB17VN50NPkpoh94xiUvVK/9XjIrLsNe4QLcchlz1/OE9hsZTHmmuEQj
5tEGUrFT9TXEL1vOP7C9875pD9LiLAp5dv30hFhUcADkejmwibgNorhDheQ6HGrU
hbYpiAMwj8oqG9sem3+Gh63byw7tUzyZNtzV+uHvz3E=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 28032)
YVx/NOr7U5smClFSABe6sEotDljVFfPgsd6HekaOhb63Qf7qrJFuPknfhRGEPKp3
kcb1HooF0Gd8LrCVwRCXLocfQOt1LCCzD/KxXtrXw59CxsyFTTJFNhyQ+vjn73et
wcNy1c8L4oyIkcmkfTt1hB+mLVHQF58bsPrDYBhe7CFV1IbmYsEBjzgazTm5NRl2
VgeizcX5YeYPx5mxi62+LH61ZNP//TXrlSqWAlco+Y2UsY/xyvdpIXiNdcTMYzfb
k/iLpy2q8f6AzFYWZgbLGAwcYa/h9jRSncy+m4geHsuabqWDJ4RsEaR4FbxAieJ7
UWgxm3t5akXoT9ufQ6vJ6houxawvSwtAAf7bhwwK0jYgxHxtFgT+CstPQOplQbpZ
7dIIqS8pqnaMJitAKiWjssL5+u3vTZGutZikd4ApHPwdTqD9qDT7tU1XXIwEeIOj
FI4k/wzdsQiNCjJm+J8KSUa5yCHDuSVTBPAtmGc37+VPtRRBo+cfZmsPy4O7Gf3d
AKSO+ZP3agNrfRfrV7zhiatzKePuxTJ2jrnAA9YrkD3fKt1m0N5dud+CouVUTMO3
CujDJUC6wYMjrwhC3G9IXeKuIguf4TCtxCFUsSj1ZCV2PywAlXMJM7JGQGqofpqf
Z5ERTjRfRrX96G54TaSWJ8EmPo0y6MGt8wc2u1JUba5z31NMW42mclGwEpbhg1R3
BjuNsICGyzdwD02RrRkEHs2t+My//Tgaj0Bhj41Rg2qTelX+7GP01nYoOZjOQio4
zrT4eaYg2FC1TvFTjL8fA9Tfv7zKtQanVC/rovJVuoR3vpOXMHj9c2hTVHo9tcGQ
4ns4BDOTwHnO1JZLVnsTgTngswmGE8VC1CXxaNU8fIt7ySQeTkBoIdntCLOEcIzm
A4e40qNVsbofXVtShDEcpxAck3nFVKjf6dTF8eCXBwvUhC85Q4z6FEuonCPwnuNx
4WiJzRN1gBbEVa1T5q/trbaq9s3A2g2MhB2hr3LHrADZlvtxsAgeypkNfzC43NMf
Vaxj/yXFPuB0egKn0orox8pn3Q8q7Ic9AJihoBX3YLTelshg5ZbkVLcUxSYe2+Jg
oakXSgzmT/FIPjpd3nViVPKi2uQszxm/OHblfmd0dSewhOViyj9c4xNeQMzR3ksN
G6YOdkCAGjraYxXfjkt+GTMORMWgu9OHu8olUUI/M/Y4KAZG4ogHMTpLM9VLCJi+
W9r7Hmgv38+fLkeDGOAeEeG2HSj2r2L2FCI4IgmTxBvVNqcDNBN60ou6h2p6SJJB
AvYh1BjeajXE3DIrsI/fbQl4MS5dpYF8PuTx4pe5vU1xSWWK8DwonY0VDpDFaZle
KKF4EJLYO1wCrwVkRTAf8CAQGBy3Agdb0JtJYLKaIbcBjmAvMjOPLgVRP84n4O1r
PNRJfm+h8s5KHxv3XziUult6lV7JiyaXPkMzjUdl4jsFjUZYgkm9fF2P7s9+si4z
yzj2RYdwtMYM6AzLeEGbYbRo2cU+4DqK3uMDi627qFRiZLCQIAr5X0/39W3P5q5S
BNzXQipQ4MadJCG1K59aHMSPgiUmqhYGju/os/OUs9NVI7Plug2FONlVtj/abWyD
mqNDWSVkameoHJPAnwYNyeS4SqP9FzEzIkwQshihuRKM3ZSLb8rMWZecF1wAxHbV
cD6VUo6TH30BJhdZhAupXwL3DSkF/CSjv0nvgnZ2N36uszDB9tGfGZDV9NrUyp0U
h9veFpTpFjk/MDmMq3eFBp5hhgKFXSkB3cy4p2p6LddRSW4VoNaNswJ5IYEWPFV1
hpzHjt/pkqF4dtrv8jrnuxoTrKArMJKv0HRum+UWrIKndqfskMfokO+NwXwM20nI
Bc7TTpGgxwumNhrr7DIDBhiLGnGM60lxV6OyLIx+Tq1J9vU/z+IuatfGBIdsZ0iX
5OJkIq3p5LQhccZwZsn6Hg2/WSCk/AUiwtOJUMP9H986D5rJubzPQ4L+XKhWCqyT
70bna0L4CsNrc9yC8ngVqxHy2Bjc4q6t1uJ7QDh23xxNVVMHVr7BeHAA94R6nkSF
DwwB0QW8JHZSvT7ofQMudknnsQCO095HgDgmQ4A5jNQ7EreafLF0sZeIRJTxH9J/
KZIqxyrXwSu37sMLUoyJxjeWt2DbQgmWu5NXCe95SRKopY0mXSu3/sBM32hoAPx0
+5quEV2LBqeDtiw6oVbiYWD4cWbQtTFFHvPct1UiDoWCUIaGh6aHzrVwaM9xhFGY
fKDWzSiBh+oeDXZ5IJJCBL9xVOFMezzLCCKmPvpOpffkUFhpGzrX8wtF/0tl1aum
L+BDtMcsskpmrhNeo7kJEg4KO00XLhHPJWMA0DZpuxSecCAmmMrADjWJeujnIgbE
6dotECkls57eQWpDh0AiC+fClBSnc7PDbGbbtkT15DxcFVLojH/y4iVeXlAVDCbC
G2iRF77HRyboTaxk05tyWLDf3SZMPpu05eoEr7vBYj1K9hl+heLoxUcAp4INvtMV
EaNP5IdzqU/wVhxRMWXY5nqT0URFcYqJQpesKxkxNl5RKyfoBNMoAN7YpsFd7NEy
BQE3a5J86VOnif3PTTNDXBXO1xJXNG4ZtVpEVrEhC+AuB98u1lknsTDRuXMrenkP
2kihWP6LTLHosM8Vyjn5ZT64ktDk+9KFflT2q4Satlve2Pq8tXYPONJNX1HPyYHB
cy1BkfTUNl1G7v9pNTPr20S+XKiglGeE+E/toX2WrrsnhD6y9OpyHrAtQvbHaf1P
OCAJltFSDx7Jhzoj3JmxHg8GHu1enigx/NBgDmwkzcoEPrYcKJJvd56Xit+NSA3R
hyrVQ21m/ueDXUUdMZ/M92wTHeRmW9wzR9ERRJBinuSod0vdc1XumERXn1BYxGOK
9oKpGbPoHgJntsXIdUYINXDfPvuVS9Goz7R47CfQDAPMXpjKP+INdzE0eNABiSZr
jfQwSyPVoqY26EEhWdJwIXo5cCmcY0jN7JuzGdEo6dVCJIaEV//hgkO6NdFxkIXX
cS9JTp1H3Xa/0YlGHZVsgYqRKkYyFSn/i6hT0sUYaFgcwzbT9HNxlPeEcPpYXC64
SndAMdii4R9CU5SUBgHYZdU/ayaZC/mOGEILalTBO4RQLvfcY89CCgzU7tbyTBR9
rqtEFIHDVhdazkFMgVsL1kZ9pqFwIfbvRNa7KKmpMG5C8PH6wRatBTkVeYUYs4Ef
NfTWwAAQcM+LzLlgZ9Q3lxPuCkWEERHn0Vz/33wVBRcFC1ptXdELoGPuakcu/0a0
GtXokdglkdz7h4iijTNUS7Z7+o/Z9W+hv8uv7joU5FRCkXgefbP5agk8EH7x3jlf
/Bo8ARWUTtH7lVjkLM/fouJ2jo/nY8p/5+v2dDFTr+PYd31IibPFgo009nGrnoOC
dMrbYiXrc0i2H6SyBcKiUEC8fSAWuKiHgD4gXwBdExssSKnVriIWv/0DOBk6unT1
s9fC1/gHFXXPlLnsI+uBARd3pU7VVqWEpigLx4ziJbtkctZhgaPD3KgrIB95R9On
cl8D1YA8WTQfZgMT4NbKhbFbRcnTLPwlWnwx/WTp4fQV8PxxdlIyUxgPlK2FazSy
3kv7znaice7Q1aEsaMKXAFz9ZQEZia79VSEcC/AejuPLYEKK2PdMWr4CL9TMoC4t
ER0G5Cyrg+O8a9n2z9/JUqGDIC3dpYjl3Rcd+m5XqnsSvD+e0+31egsbm60mLsiR
ZBM63fkwoYrIZY03t9b3N88srpvCxRWv966fyggaGXyil5U2nvC2YHBD86No8bVt
6HgQymPFS3IHyqo6axZDYdNKq3eY0ZugsS479VXbcMVIhFxiz1Lulst+euLEekUo
rSo8iXBWCYULNbONewS1sMe+UlvSyqxoGHmVRXNp4qI2kyAvYzeGwat5HQjuj0sP
2J+Dqn4XBkQpiJoclG4fGJ84XBny+ExoShh1rkOKC4DCqn8X7aoUPRiN29ibWCEh
I1BWkGGSd0qzrUq7UJwU0OveI6zCzBRb31gCNRRXEJgOi92pCsznMJSbXxVALLOw
ixg4xL/A+HX/Re2xcLP6iFKwdQWYrr5Yzjk3mXmdMTT+JPtsZFvHD8qVxuUYaoyn
pZlPSz3qQfECWZ+DjmWY7yYSeqsFPM3gykIHVRvZZlFqpEWN1Qk4YipBfGsJzPJN
Ed2hAb60O9c+O26JYwMRyZKk5RKYIhRsAvZ/FDU12MqOtc+YJSHR/2jfWFGpmuoS
rAiWa6963rZkTNcTRkwJg8eJi5UXIBXLCHKKHJzllbJwlXQ1FwOZ0Bov3ejCnOsF
nciWWQU7Q2lyZN2SrDPp/uKUvDBPZAKiWVI13P1OqwO+LbVG4wt2uauf5v7uEB+h
RW1IBZCoCNN8i7SfN0MniA3dpsAKtBzWAVjH4Th7A2wToO/WZt+UUjTP4sWuQsgL
5BrTJAHBhMAZP3abW0x/+c87hYUXQdwZvr9OEgbZJI9pyf1/41ViLqIxuz11fqSs
rdNoomPUx1wLX/dEk15IE6DuMrb8GRoCA5UKkjqyhz77pOPX9PZVDeRLneGaU8yi
+FH04ppI/zqgPq6kS84s0HYTRPsEyf6yoz4Rqt+kxZZBD/5MP0Q0reQvly8FeG5a
HnAtsgTGeNhARSVQi9lY/7tqKdEj5rQeYpPbv8iKJ0z0LeYOstStDjOQm0O6JVjT
N5YS1VxWL1KTwNdcIH7pLrBJ+4aEMtr+y90Wv65xxSYfpxkvDTZeEbrwvkIlDBLF
UhVmhE9nWKGNAITp8886fQJvtigTTzojfzut/7b5uPFQtjA69HuQCT8cR6wMzGYz
yAcQknr6VVpveotrluTpCfla8iVje0xSMdLr5TJYoSo+S4W8MWZBpBKTF8WO2fBm
ynJ9yLBDXS8AqQDe3NvmsRwCn6dQjLcvx/Jdikx8uiLwzIc6w5Kyx+NPBhPAypjz
K7i9w45Id0MoAtqZ2wBsEZ+Y2+MCEQIJTs5Qvsj8ux0ZM+Hd16reo38p84+Qvsfy
knDrBM1V6b+er8TXppmMu1UHfQ/OA899uoFVfcK9DfduyZCJUGu5sTXyXqyTKioI
P8yl4eQ/N12049DJbyNywfbsCk0IbUCMOeFcU5ztuteCgQZzdXjFER0gEWJTkzaq
T/C7Vlfn6jVye2tIk+G4XT8t4v5tGdXuSKKZu8v2xtjJ4qkoHKLzTunwNWx/mm3s
7KFf8ceJb6hTKfReB4X7+39R4V3t6WJb2MBbMpZ+sZAmGDlwrokWlQfp28dRF8iY
7X/eGmLImfn9Bke2cPC4ArPMosY3r0pHwOvww5Tqt63B4vN9dEOb/6SmDDajO9Qb
NXUXe28rsQpsU/dj9PwRI5d+TYzmSK20Yfr0sbo9edNGSetsNgXZwxDwyJf2iqq+
ThhyBsJ+IXz/I3YSd1i6rDOgGl8mIa/svm4QPkG9u8pQVqzcPgF8M5+cGbF1oxWI
QHOvtjRLEPV0PYSkjQL61SZyuT/OZJXFmmmv5wlCuaIsnmZXw+LwSPbnK5sf32+G
9vZZIdtn/choL8mt2yQMnCtBjdycR8BpFgNR43fdj192GDwsoFy3Z+z4YLiBxSSB
w82MCMDWrfNngiMj+AzwEawuc7RNvt/4kmgYSIxIyFSwOyiJV/ZKsMeSNj+jKzqy
lR8AYaQ4+HqZhmwfS5C4c0alAbkbYZuOYd2o9rPvF/dzyQo+uD3RA5d6hGeUGPQm
sGMnN1nCDvZuuH287D5r/qpfLwJpgltLEVjOQEEIQiqmSkwe5vrVmPrSCLke2KWm
TK0gjRAAa9uO60kOhuSfMARVmhXSg/Uf1r0/tpVqgzR6JBfbFB5OUlYIj/4oqRM8
z6crxVfOmmoIa2TRIuYSgnEKl5iAFgUhVVgDhnzXi9HpuaT3iLx+bOOTG4I5g/q0
m04hkDKrMEh75mLYrYkAZAIsEarTZ7+RUVnx+khr5gdKjNua70btZd0JR+GX3auj
2H6Gmvz+RBzjGE4xQKqe0G3SASZvSK7hSUf+bKFkWuuwUX3KZBjgv2iEmiJR8SNh
GdU0dwp+b2m2axKs1bO/lHsFv6jEBwBZQhvdRiR9nHsF9Yj9z41m7Aux3nz/MBGA
XsWrmdYgLEyekKcSE8G34N1ZBSVkCoc3Uk61XsGN4F66PdDFw6OYrXLqUoyUVBCV
KAyIipGNw5XQ2RJkVNk0BtHT+waunqyeVerdqB8sfrlQ84enyrGWVBEr5bttD618
Cv791Tf+vOu/r4lr43ydTnzHSepXQb/1mwm2IN+x/p+wxtAgkiJFDaFHUDVmJqPY
D61sDKecQuDSbeVkzvv1PcdHOHBNKY4nPdvhPYxZp5ktW6a6zV6Dkhy5infoD91D
5OoeJNKlnpAnyuXeK0g3WIeJOpuI9P+Ptyvcm5x1z5Y/l0VsSrQvEoiUo2CZ6mH/
FXf8pUH/S2QWJ1wkgnfNHp5Pesc9HmSSi3YDWp3bYk4YjoHqczaX7AH3RY1X6NCB
qy5gzJ1j0KAq/v9mXPnupkzp+DRnAjjpKbkgmX88PhCSUZl9b2ZXWw1pOMcVxURp
nt5b2hkBFkPyEh8JBKmxMfJ3PQ4zuEsqQj4bOWuYFxy0XzH6DkA62UZeRoSNRk8O
2Nh3hwkPPnuET3oQ2iaikqtYdzXKRanSKh5tx4qY8ueDT3+e6nDT5aLqa3a5SouS
cgNWq+lcyNFYh6MQiNYaaGvvFPlLSVyZfaEt9Myt8R2ecBjIc8o3e4gLLQYVyXcO
dPRruIOggG71tY9i1DaaOuWV1M6tGGnvXC5XUT/TuZFET75URyRadPBHYn9psOm+
oopZ7MjDNLnm+n7oPj9hPOplPQdsYtrF8faAO4Ld+Olj+5CwN3mVHcvKc/nv3P0r
9rxVtrRHKwk/ky5DaUAdEjx2rvxUDmAihZj+sRwyxBLN12QSSZDASkSNco+qnW0I
IP4QtV00Ap6zlZv9cJWbwLaoJBPL2sWhQ8HYTN52mbI9nyG/qinBcCklHEGlEMJB
Jmf2rRR2PWkRF3LevQkAiRNPEVoCRbOS0eidc51aR2GewkUMk+A37/hhwogdIH9D
nBsSrpfiRF1ay1NJQ/V+oCtjFANMNWOPir7CA4T7BCdT+T7QvSdC1cqOePwDt0fX
eqtKFJXs/wZ4TEk7S5hKhc0l+f2rbBTYWWI9xQFBMHMQG+k0Wgkc1JwyFXkRQPPT
f0lktaG/b0AYtPAL4d1rzrCa52jeHZluD5An5ZuEI4HwKEeQd3BSfeS4cw31ouMe
yZUeGZtLlhpNh2nA3Z84p6koRS790iDC+uY0PsUGiuhkaGjmHv66z9PZRIaui9UA
M9WC8/VY051eAdRBAATjgEXG9q+nT9HNjSk8pqUcY9upgFZCjV/6aY4WUyAgQvm5
GBbBR4+8CfnvMEm5DJvcSC6DL0AdRxQm9ggg5y3mrxo37LS0v7xgQYGCZK89lkCk
4mmlDK9co/ziUVRtzsL3v78lOzeqGyjmxDpFRsxFjO3CWw8XVcm/N5Xc3q4YDBgB
VolG/ar+8UrOAUCfLh/pyIfpppBmTbhithK0l3Ww5Q7rOauo23eMpfPZTL9CURk5
drO8i3SQTFKgWkpmXxfQhlXDBFojEnyxYu+PHWDA1WTGnFWReI7NGO/siE3Ww9OF
HvC9b1HLIPM9WLujWHz+HbR1kqB1W0+KbkqBBhBeMhzSGV2KrqmGDwfk1MM8Xns/
VOc6yoMSe1Z9kHfwccTBw+Lyo+T+sd+JzXlS/1Dr4aziWEf1iXeQj7nOZ7GVn0qW
QH+6tYsLQAY8orB8b9EFi+V3Punb78RvRRUnrSgwqjeoBbTVv2fOSKhmx0+5ulCy
i74rVy3U0XP5ekzjmNn/tCqPzXlBSKc/leUdqEFM1e+cqPr4xAHhnMyqyprGv8gT
F1oIOxyBy4psWLRb5PgUkkBatogrA9itvTqY6/hvJ2Ws3+fOqw5B1pcji3ZQRKwa
XJb4hDEjxqmDyfWrlgTERyz5oU+dKGpV8UKiZeukM+TFzftfsufjKbWaK8jJ2Otu
ay6MxWqRHFEjn72Ev2VPGWEFRSeaVgW9yXT8tMkrJfgFOrJZMXExZWLyxhuA6JeD
xhwYwFc42d1m9BT/lf2pvD3iOUcIOLK8r4nAgduit8RRm9B0itB52HATP/EJKa4m
kuhpdT3XPoGZ8Cpxhvhe9BExnqjglZxCRKRglI+zHzwhEpsTrCuNIlPcjS86wIhD
STdlzfX/mzAPd0hg+XHQICno+CFp3scol/IO9UcOJ7HabdQI4b1NgDx4QI9gkMsr
eecv8cqvJoaXkMjFhq5mlTWkeOgcw34zeNkn9RX6h5EHmAhn1+hyIfpTvNKgIUfv
6bkNb/BY0llW+B/A1B0M4U0HOgmFrsvjh5bmgKMY9OtgcHjGpdy3VD7Sh9NEZfY9
ysho8KX3iSk97q0uD4ap/8uLq8d/4rx8kpFryW1r1JEm4bBZAfBqV7d0RJTOOkET
gXbhAazYtoHurwQghxIl4VKqNoSzIhKdJ17m0pb8xx08ZCTEyaA9v0+gzbvhd5Ql
4cpxQEYxtwvM8S8gpolKliIFtnu4rjATGy1y6xRsRu4QmWH1GRz999FVJWn0nyJq
rUziX4I0kuU0AEVBy7X5UoAPqPUj12HMghmFV1UOl1awRyxRod+WM9jTgxrliSuB
OAIS9NohVhgaIksEh9j0tiXPKa/Z2dkM3V9npsuQKflLXziF7hbZhaKYNsQ6ctXH
o3HQ07psPhZhVzixryBEAyOr/DNKMLvCQ/QO+8Dn8A/jAHTzYNxZMkG9xYA3DvAv
wPSvyTfTFYzJfr3iG2JYmnhU4iM7kTCUQf7r5fveI96ieDm8+JRC40OI7YFckiFv
EFud86BauIJ7C5Wf69VWRWUBrcFsnEWMD3FHpmm6RfeY9CU95s8+hhVOvLNC8XSa
OcBnmFstc2fkzAOfwCoHA4meOuriJdunlXuwrX0b7G/pJhveq0XN/rrCtrQH0wby
yg0uRrgOnwLNZkT8cvHQCXswp/AlZJEcgI9unXiJZS351HqKHKMe3Kd/WwvLqh5P
QCbR32FhPKdRjEXGMTSeB59WaQIH5Ylm4zPpCxtBv9iRucITJR1icn0QeeVZkCDB
R7mD9AHL57yOyDObTLngmeSADbWYigXiDMZGLF4sJuckOjdKHBdADNuRMOm6+2zi
HZEI3dd0c6XB3AK1xGSGL6iIsIMmhD04JuOcaGO+6D/h+JvcN2jSUThK2sgWrU6M
xE2XPn07mrNKNx1GG2yZ8BSN8E8sJbsExQVw6zST7U2rUYkmBclRy4HCGoFOrJXP
AWYXPL1wBfuX2H5TShbdn5NXttFXYKruci8cmNHK6tVwZi2ahBDRY0LaVVk9MJuC
bf1IPLCWejmJf2eM3lDUHYmt3K3BWl5hbWp64sYijJHphm1+NJb5rCOJ51dXnW/+
1X5bdCKHM5b6z+zG9POXcy6x0zrzR0WstbZ6unhtAvK3CM3MKl6eVzABSSqZflWx
4zA8IjxsUNbacQfhPkAz4//xoV002BgFqxzv5+4STVw0B7EJQpyvPhKSPxz1dJAt
3wmZTbR7o2tI1zNrfQTyethHBem3fr3f8YrXF+r+vnsPoNUAn7D7ygv++SXW1ZG1
zVCz5zGTmXWVu5le+zPvOGsbIac9QeXEueCrp4tTuuPL8U2r6Yov4sRhOUkT9w1s
P9bHs8CPgUM9F4bsXc6Keif7QzX5V6BmHsK1S09yVF75DNmefTVU88C8OtvwJa7l
TGl8M1XN1UaCQ0ZEUlu3XTtxoKKOdIGlAcycRvoq8/ALzZhWgPmFT/wQRBmu84u7
Bw72NjvSqO4V7Io1UtjnZ55AQI43E7/u0kIDiDtq+Ay1pmnU7Y/M/yHhlXbzxOmM
/I8bZ0HKbsT6M/E2uB/mRI/6vlBJDZzu5HqdIis4aFVVu+PJwDLaIu5skpNJxbrp
+8HTuV3XrmvB+8JVu4EWeCKeiO0+5h1ZGwtkxScXxT5ow0I5Y9hgCZGo7O0iRT1t
c0r3h+ltT+duhu48L4lhNLLBQjj+yaz/suxSiHGQBGjVxQXXGr5MmB7CezO6Fl7j
TZF9hbX8261VzhfgitCbrpzMKXNPoK2iWPl4ywwYOu1bAwkOwHt/Jfnr1dXEzO5C
OfUEU0BcAG8UZ9+bYfK3bBUsru5kVYog6waKuvVAOv9F3VPtMlpVycE7xLw2hkND
eZqtO/YUcNNRXDRVvxTlHQI9nHlBERHI8BsZWpk4c2tsbUSl/6QMdu3hbSQEZ5pt
bxhV3nTgR0Jshg7SQzmwgbTaMKmNipbByPgLCntXhJh7NDLKYCvJnaR/2a2G0Z9K
PoL+tY83ca7TCx5qMz7igfudi/LBwG+GOYSG0l/NbpGkiOaadxmzZOLY2dd804J1
CDBkLtkdd25bzpr2wp4MPS07IoX8zGBtk/wXY4J/rJzAWait+RII8GNfGNOUHWsv
/47CAaqNl+hfrRrwiBhqZ9tJcZe0VW20e8OWh45xuT6ojUyNUjnVSnGuxR1HRJ4H
kZ7PVZKcf7H5os/3167jP3rucvl+FN6qVO5JgypQRw5jYVDP8m08XR26KGTZdOK3
K03A6xdctKiRyZ0asVAbYnEihvpRYk31tT7tQwT81+x+RCLKe/d0y39dpHUfy5kR
HjNLtv3MVh4eXnIBLh8n1d/ilfeQo0KSoE4u49pniAnKuajDDwok3pfLr2dzuFYB
ZfDDNI7ZEdcgssli3Vs66TS+ZB7Ujsf8bDHOTHb/KWRpQTjFlXQDpH3ECE7aYfjd
34xpCiuh+kEaG7+yAw4XM1t0kRah2AON2SXUmvi/8Bv5dbz3e8b8e4QiyS9gB6f8
7k7AMRuQCWINm1GRvwDXEvihGUFZvxGdJv2kpQH9w0Y335U48hPpRMqEfyIvT5l5
kqanSh2sjBI3ceRAdRBEc/sAdDUdUkj1FJg/rDos1NuYGkdLNLTh02labKV73mvP
945s+P6buksqeIi+cHZZRzyy3sKiVNb5o+tpePccNsUO7T4x26Hclr8esOQo+WVJ
GwEpg6JvjXpuyn2cNjFqbLzAIvkPv8ReXmnm100R1hH8Sda4lhUYpCtY7P+CQM0c
ZzofPBZNbL+zTcw+9K4pjfBF6HxHP4VZbqCBXPzqeMnOQnaQq06Ddayj+dTHgFwk
qd478vtnFXv2AQlf7UpSnm8ABY6cgUpIB6YyjG38x+zk1/C9gfhTHSiTfA6QWVuQ
JT0Cilou86kxq1Qtf0KbEaarMfd8E2Q/aX53K2TRFB1XyFNYlE+dCS1O3NPFVtzQ
wySZRaf5L9E0ZWaNgqG+LvNtQM69z2r4sWSsBFE+lckNVQ2Y1C0ClD8OEcQATL5A
1s07fL3UsNe0wi7BRiXgtPd8IlKFI8KZk5v00zanRboXBev7Lpec8Wd14dsQ1GZv
5OzPf4BY4Qk1kUsGWYK1tRccdYN4h4aENyPX3iHA74+7ic0VNU+lHIpzyp+r2ZeX
/PT8VHGZGg3+LNF3Lgxi0RUC7rykDZ9M2zJdIZ2kQ71dC7jY0Irgms31MPNycDYo
M68ddXSYoXeLCIRTfDktN04pT0IeOvAxV+70o5RF10sNMPjcoZINdTB6jBxlE6V/
Kb7V14/3qchhAN0BbYQgAn0p6dBT3pPPl3aypR1yoeBhWAfRt6HEKBt0FAmDEpt/
lbwpSjMxZVl1jGe9OdpjhbMRoL9FWFqrZ0S6QGHjXjz0oaUeU8lJSDnXZO1tubes
c3gIgis4Cf5eGkeHRoOMvijyG68dZMKAdDzQOgW4LmgM+Mj5RyhB5uov2xVnwMyk
fNVc9Kf8loasU1Z83sU+Y4SkAhAL1mqiWb7x3cm79M4MRKkkn5leg3Pd7/O87ULu
bMW8jqAQyEkrJXfTjwMFacfJZVuJ341af2S0chuUAkq6Z1xQm3Ro2/pnpgWVVj7g
NpnuO4wIE6nP2epjDvKIlIxd/QdzcPjb3+tHpudj2fQQEHx3OQMd0sPBgOepYKap
02qlp8KvsCR/DpZFjqk/s6DoGB/Ce4yswMopoHR66hLG3sMI2DhaTrqr1Q9OR/nr
RUpfjdT2bRo/sKuOat4byVaYQiCckERrJAxecnAiS4Wp+OFK2JaP3UBEfuDlkSOo
rNomxziPTwzk9Y3a20Hl/zczUvH57uUD8btWG06ccvFSEpAg6xkxkjohVE0/C0oX
zp3Uued7pW1JXqW+xrdjRYuiBlY+dl8TvoBq9i9gQcktGuuCONmnMq4GAeFlRNxD
TcgJf4YvvgVvwYE0i5yOges9uqmdadYizRZj8I5AWr+o8qaq4AdHzComNNvJIHac
TQBLF8cQD3i7LiCWJS5ZE7ejoUNjNYcVtBv7xOT8ILbH4GdbLQ+5mXCj/3yLTKps
QCqLoCbbws2uno8E/NLeSDK8Qm/p8+ayTWPj3f2p3Ow0E3dKj6N02PQRJ5pC5Mnj
48DU6RoMSgVJ0ZY7rLqEWjVedWfNm+ot921gptlbP/rKqvyTAQV9mNGt7Ah+wZ5U
tPFuk1kGTdmZ8l+EmqRaCNbuW35iDLwbTQNXjmCyBA5M/avbSdA1AQE79uKNJLmO
YekodRjSXrvHu965yUphARujVL69PduvvtoZU/bl7r1ZYjhNfsk3LQ2ZgL6hEUXi
KH32X/J6LJ5C+OoMQPAruv+CGNRgWK82M4wOkhHaSyM8SOYoq5TyHQr2jpbaZRKM
aTZeXr65U2/pbu5JrnIXvZCqmCTvsMQh2V1RgAWJNtfco5PeuXEidgrR7dxmWV0/
a8ne/x0U6SDM6yWL+BKOCHEXN6qqDpuXsI0pq18ZnVkH3pvbG+KlSdfxjOOcOXE7
DDyWzTrNtwBAjNutH4XWrS4dp7fuQIQ9wbKu8UCWQPKGpOavE59uz+GawxsX3+Fq
HbOx5a5G7EZ92dKdVegMQVNypdwgT7th/Jm0IwnL+stphR4EgK1Xtz66c/PxBkII
F+ECPcGzsFsU9grbLEgDJhKfMDXHBtYIWgvZ3NdrwNnp6zu+Q7OXbUmNLBDf7UiL
O4uqqfYvbEQ/2ci2nAmAbHgrtlshSjqx4PM4hAEN2KR80ZGNeByIH02E4iu1aSaE
o0NYoCeT+AYUPKLwzigJ3QEiXRL0OYiDIc1u9FIthWEPNEG/qQTE62Ko3oNSKbhC
FYelaVUtAxLkjzbg+cPPx7jAVB5W7X42xFCvCcu/Ptnc9KYZTB1HFMaVAUVJQXpr
n/NdS5eSkhPa9/0P9pk3gKhPyPnC680u58oZkQbUBsQBYoOeptdsMk0uIVLSBiSb
J6doELELYKR2v8udYLMqCsRM5Xbq52mhfw+YVfCw5oS6tSonr2ptLN4E8uV5fvw5
ULesMqsurQAzhb8z8Ihhb70GoVpBXER//gxXRT957cEB/w1CmmyAYQvarTUqNDci
q7aCH1HzEPjhVlGUVcwjX/Xz3DmqgPzFwlIAlqSAa0wLvjX1ZHT7qfkSDVPntgsS
BFdXWVEhLsBY5QLpkgArI8yqsSEHbjlTnsu9TLbRd1zvkcWFbbFwZ5vJ8nisuuRY
156c/F7uIXDqfY4dUOIskZprTiYSytKQ/jkUD/18a+lAYzQSfFR10h7Q7mk8RyP8
eZKtGz5Rl0QBLqwH6FSahZftM6zOKI+7oonmG3jA9zvjhnuNGLurti3MiZIHwucx
hysb7KTPj0yLZdt+4znArnLKxZLEfCSmtfrjJ91WbVYWCRFvlQdIjfO2gLljWpCX
DkAtrqIdTQePy9kh9omZCqYoWjOKdD0756q8+V/dEZHYjyWe1CBYa1ID34O7zUVz
sEQKtUaIt+LNUzqBFiSX4RwNfKvK0IvBJFR3anB25zJxYKpbVx2k1VeMz/sKcPiB
41i/tcp7CrldrbyfI6imcsbfKBEpwg784OaLKho+jlqN0rOez182och2qbAzDvPE
FvJGqAZOsgT/+ictbQsU02gQjoEa2OGqI8F4zgb0qhJCilnrTBu/tT/F5rmpTgp+
nWJOEetRBbDOIO34LXRKajh2p+uqCCyzvF32lbpQtUsxeWg1YrC0DZvS+fqCl5nt
FgVVZce8cCNM1rI3HHmWm48oGPZw5gujJWtSzvGgr7UY0deiBFT1Mjc9iG39xiuL
c7jk62/OWi4dx6fD3mUbthVx6Qu+PKqEnQpmOmk5W0k3BWstDS/bFl6PTBmsTRSC
j+3eJ868YoUhAMgTL85b0xP7hFKs+9h7QcheLJjR2xNozvFtpfgWIQ4b2wrw+Ka6
zA48VX5BS5ObRN98yWQfYvu3+GffWpaOxpwo0NDmJZiD9FCOoP8cQnxFy5o4eD+b
HNApm7lUfeawf+DCoFyP2650x65Ne57cFWMgNbl2hVu1U1wjT1ArlknUTptwLpH/
BIatuMftcADSKc9ryzZQCvc1e6aCpeGyEermQNZHgyyieavfqr2RLwNOpoTbIbjH
uLABDoP+QiztllZL0ny16iRz9nLimowuS5ujooPJ5KLnkrFOdv/OIYmscjRaPQW2
KSaHodzcDT+1Ej25ueYlWKkIju++wW5bGmxqbVM4zLZ4v4DQ0FStQRknhDXaf8TX
0WoUMShEtGmSs3qvijOEkGZnit7cJzovNBUuBXtklO9E3PVfXXagJXYs0tzOGpRE
6oXwj/SEDkpN7l8Abe5c/zupbeFYHZxmmfqf8Oe4vEx/fesz0WwasZqS9XySdgdy
wJCrYGNQI5rlFiGaCXOvPX5uXdMnf7oCnhoi5FqMWqI9x5jNBEh8HMbJcPicwX1A
2wzxH0aWNcM9NBWexYtlmo+268Kzw/pxubG1RbNLMa3FJdVnq/RSwApYHCEGRV4O
WnOsEns1Dnh8EQ5oygukW3piJAuMtpE0msXZSJ1SBEPNY0eM834uIU9rW1XNCA+R
5Iu6srlaVh+kLG/LwvP0IVBd/tkLEPy18EB3gKtmEBVz8oqtZfzD7E4eSGSelTue
LdC5MxEp9gIqDPHseIhZxalxjOCetIO18qhbiiHlr//vun54FKo8+wQ569Hb3Ahd
rzj/00Hs9vVKTpqDYftgnXJIPVDzzcvvcQTziuZlvky2cR06QbzPzJv7KlSQqYdb
bK36cI4+rITcbx3c9IiricCeLMK5FIRyXeE5PMVpSQWnqbCIC/Li1S2Gnbsuwhej
2PxUdEaisR8Om9yQH4ZBXQ1UbxwKZUXYHoFMmdiUE84H5nGkPYbwOkltpFZl1kxv
vqW8scb93xamzcDBpvahQmf2Kb9Aq+JQO+/Rv1lyaBj846pdDyNbGuq0Lq0wLmN4
kcGAB6QBho6NWsafVfygL573MmgFp3B1B42IlBEfpy666IY8p7l7teYow1V6wPb0
BSRRnN3VMdCAh3sChro41d4jecaapiRZUxtEU6rLZdJUKMVcAnSWDwTOY5sa4Fp0
RfT7P62k8r1cqj9SnOkjtLbpLDjG8EPm2ZyIajX8uctiEzBwSh6SmZWXs9NhtRSc
0XghMfjIknbFEdXyHNzd1vqxUKQg1a9GGxp20njW3ti/OMtg1nqrlck14XVAgTW/
Tn11uLMXVTtE/SJsFBgiJbena9o0+82NtcVNeN+Mj/s5pxMcCWtIAtAwskuhVxWd
//GyipLXKLH2GgzkzK+6//ZYo4DL9vYa4NbmezArpt2GzweLbXiH2hWIEb7clOkE
i600IR15QIZ0h8TzRcoK2ipEY2ZBVXxkfPeQK+RTlmVL75GxYr+kjiXOXLf+KuE5
aUaljRiuxBLovKj4Z4r0VrJB8be8c88F2lC7xEKbJFsInC0UFeWYxMFfC6QMdjge
OAw7dY7NQj4k3EuFK7vDTEjNVEm0k6OgcymprXFZxKkEWoBSDhTBUMDbYM1JgmPn
YytznP8Zw71vSjz4k/fgvFEvYgPObFfj+j/9iYB7+c3eAaWuf3c0oetDPsH9/1qj
EqxmNZCz3TIa8A1c97Zws9BN4hLg6jBRBNHYq8mZXtftRgY/6o8doPZzKr0Pzu2i
Yvev9mKFLR5aht7BoaM4hSzaFnvoxHALIqzpWUhyys0GDoKeTTiZiZy5TQHpzOa/
x0d4nkaT9YKow3xqrOS3YXe+cY/2oYgQHsdcnosVGVF1HjV5CUZvM0ryqOkp8kPo
051fETDpX4djvGaFP+80gIdB2/tCmn4k7JwRKqTPEcUJ3vEky29J55yTYQqX1QI6
D6ZTmrHsHfFA49TutL3Bi+NBhQDB5eeADTy2U4B90kFk+qbi8hBno4wuKK/wkLg5
hdT6AFaJGdiAXmF7dWrslrOHkK3AG/ub2VstQCrVetiMN/pAQWhNS03npORxgClK
HkP91STYwhj92IJJFBGg8g9zd4Jki4e/14f0wkgJNUXApFV9rPGqMHaYelngomwf
7Us4ERwSO7kB+nFoSGiYtJr3uiNB4tr1IQsoMEzcEFbOsRmD4gKsXBY0CgyHCF8+
Kh15+llbd8+PRo9YRru6MuuwY3lrNgONgICRFlO93EO0wsD4lD8KTMZdZYMV1Z1b
0zXvGXBhNbQm7OxbKTW9itPqZYZBw/WwPD9kNptFtkAyuUe3nLfqRF4vnEeEIx2I
b7fqSCJgtlYdQbkrIpBGAdsZkSS9e01zY2VyhCn9QdHJE0LyguxEIqn2AV/L2s5x
vgN8b9UiLmGElhEpGdJnRdBFH8QheEFyFCiCI49R/2I7Nmk2JmbYrUq19j4tplL+
cQk608abL5ywS0+fLtj5NC0wx/jNUSVHju5qN3JAxIalJs5p1Cgzwx8cbAZb2LAf
0iTAaWHYRI8xyeVbm4GQQ9yo+XVXdMtfUr6xMffuCM/2DaM7YYjlADCAbJfshorW
U06tOzFdSNYKNseN1oHsszSACslB136oMmKBHkk8eo+F2TiFHueOfDnUpaK3fbIp
47oI9KPWOnTk7O4ugHG9Mfi+gI4LiXMlz9MR+FPx5AVVN0niEizuAQB4cqf3eIRg
1Um0kZVGucapn4MqFYWCXdzcn/CBEPpZpC8W4xm5ysqx+SvzJRukZt67WxvuFbME
3b9wNJ3vVoBIDAfFSTqCxa96XDXF87TSyBcBzEMIcEF722APa4pINztd0cwIOp3A
tHrRpM6SPOOXfE3pCM8l14aHrf9lGPPQc7BR0F98qGZ+bBioGOqMRm132Jydrvio
+bewpXhEv/aLRh63z3NofrkMsoyhfsSuaF8cVFdo19kRNM+q0IrlfYN9KB1DsQ2F
3S+H3lij9RrepmBzEbABSneFtl7YSyVCC6TOwFg9NBlrR0LLw+kFQ2XMEW0uRPfb
SbuINdUZfVMGL+QK7hk/Xd4Uryjw3JViLDqI89KLZyMvyIeBbBUWb/w24rBO6ex7
4E/x7d43B8ZHUxwBrSE/nvL2yvD0dWNG2RWJpQ4POZ7PEiNy/NPUl6UHlnGPUGNh
ztKJNz1iQmwGQGXG0EzFE3JM4K9gqtX5BHpaI38YEZhHMWPXiBPmaRcXgLI/ei+4
S6DaQTEroVLDNJk96QgbvHZ8hLRmAbGA6rXXr1VZEzfTNFFgmkHAN1Tm09awb3FQ
/JS3j8WbE1R4DFq8HquMJEcxmBBBu4vuNMuY+I1Bhq5C1h/YktkN9WkVkP+V7tys
NAaH3a41e6uENyLrY6fPtIchT9J5bVIraVsvgNP37+VwTrS7X6YFGT/fBwUv+3PG
R3Oo6+gfZWlI0x0yRMplqyBAWLghqQzDRGZ5juxFca58L915XUfypwzP+dsVYOX5
kgDGunjlkTUKANIee69fxplZal0yiEM78VGet6BDrVqHArBqZi4lN7BuxVJYpKXz
WAVMUF+FAPrzZVuTiEdnI6/SDS+0iMTafpKwz6iPpYCIoT00j2XZaJmCKMjCTFBB
fPgw6mRyMjRbW9C/Wx7YJPCXPZxU2+f5OV0eF0nyMfuJ24ayRPy9kcmWLA3H6saS
Y36VU55mjdFjzdbmA4QpMUKwV230oWiw7VmBfTFwiOoKtN5lCq0bGUdqCL5RT+GW
2pnS3WL4gHce7iAkY/3dDlQ9U0yMf8KCmIXDUf+23P6V+qsHPmS6Scz56K++DOuS
/q83EmqM23Hcq2ykF61qplfDPJf3FDLSVhtoi5g+i7uYhWDVZfkwGJZOuj5PnYsX
/QVMWgs3FtHonQXwSoMkGdApowI/8VBCksTQLUj10N4+nTRwELca+JdELMwd/Hk6
TpCJcMoW4K9Yz9jpIJ1QgHy6ZHptOSrgRPx1TAFk7gWh53T9Kq9CAVgTu1Q7EEco
zYoCxvRfhex8XqLcmJ1HnEOo1YFOIkPMCXm6n7dMTuwkqjD4xuW8eaXcfCLVIOpv
K0c0nDLxFel8D/NtDOrlEYxR/IFxRqDR3zA1GxPhVVCLJeBPV16b1QZRJIyw0ran
1ppieuHczs7mLnnI1+WmcqnAO+erneHnTsrvIh4KGXxXiE52amwn6iVno8TBvx7y
RskIUHFjGVOoVo67ChopjFEclol+0RYNHxl9TqPk7b49xqujkRBRuSXv6E4WEBBQ
hGl8S6Chwh8mz8eQ2bWiQ/OpKejiKcd0Nte9nrXME4Tu3ky5/2X33cmugXIfS5+I
+li5+4hyVSrFYH+sAoIJaCiEtRwTJLv+XWqvtNE4joSu4x1IB7xeZfsoSKC26gUn
tdnS64C5iaZPDNCrjZiLTQ1g0jPuz4GreXf8XcUZKyMQfMWCzBiYpHMiZXxTJFUw
R1et2Bp0ZRafNJYPC43hj2eKDBwGiCFU2UmFJ4PcfC55IfGSu0QbErsMHMztgHGG
BLALdeqoTcIhCrdF9BfCoWqEBPKtdi5esPqu9HM35RY7J/yx+D5t8sHxX12yYz+Y
2WohlJ8Vm33SXzzQ+UdYVK28PjRv+4n5VA43tD+RhH3PTMDCsOPiUC7LUYwelTzM
dTAReCUsOtXJcKp+mul9/lTS7BXK7vLGG7P8ZwweDKviiGnjwsv//A42w0W9G4H2
OmjdcCIFfqfiOZMd5LQmNnRABnovOZ0ufRwIXwqLMzXtCg3jF7zlfXOfPioyCf0a
59agYRG7jbNfvQTjYtueY+79QLBggDoDdK43/pMrddWyB0zX9jHiX3K+ebk0RWCX
Zik1HIYzquZgttZZF+N/uhK4DLOiHUq/aFtt/djM5SOB6IXXaWq9Ty4XPiDxmQ19
ssEdH+i90A4M7P0sAVJWwQWkUgDuoFz3zbWPFAhCBgBzzBl490u/nrBtyFoFOc3x
kUzQD5nTubMpBCAbAWe4w6H5fv1WXRBFNIQpt3j5Xchjc1AGl+zMsjbOjjSgiqyC
4/4XBufg5/ovIlzpGqjWziybcc9QqdjNEUVpYFSRaJQkTRpxVMuS9TlE1vpK1x1t
91aNK4YytGvPB2TWpgzH7Y4y0q5oKkhqI2G2eIE6jGFLaVKITs6ofB8ByzBdzWgc
lrkVfPYfaPz6gXOegyaGVUV1FCujWygjk8xBpgXmsAYkme6P469yo2GPZiGDAkYm
VRKZsAFRVGudFJNQqwX5yVYZah+dCi34KxQsRSrjwNP73bsXFADKlR/oGKshyjTZ
IgXSAGl0YIkyCtUiiNYO6edlAdcmnAZkSXvRH+JD/rguF0ONZukrQ4m2g6pUJCiU
YLAGlsWqR6dWLIb1Vy7jqcb6/XiFnwXOtSX799nX8nVu+wvEa/7xtzF4rOo55VCI
Ca8obYp4Vcbl3b3f8ROmqo8pQ7xb7dr5fkgpk9kP3K6NxeauEkFacEyIAhq8TbI5
bIYz15bWxT1eGzIFMTesLCIVecpYzQ3GPUIoriwIjdgUdTEjh9RhxbU/p8HCHaNS
hMHSpsbScsA6U71Ja0ItnoGIpXtTo9HTeEJdMF4YMv26qLH3cQrETKYgnkzW+f4E
XDNsin7eHjawv50to0RyoWz5bVdS9ZI6Q0hhdYD27vAog/RjdMZqw/DSr/x6Xxor
Us6b7eH/pEexgQJVfDDNmR7FN2/sHD7nHH0EN0O7NoPLq7QR5xZHd0h2fG8YERZq
xKEYNRdZv3ZasxnI6FPJX2+Z2tyq7vFNOEp0UWgAEkY2vuGNKi7+9D0vO21RzYlG
Vnn3HRmam66aYu3BJOEF4I1guYErp9TH97uwtWvQS2He6zpwtzI8mPCco5z74qjA
jRqY+eHr2KtdOqDAtWTm+6mnaFEYdrZD9WZRqtshNbRFo1BcYw0ElFbnmY+fEMIY
0BYTvUbJPOdQf6bqkpp91Ydusa0ShYcQ5E3vtNOJHKBZAXpfpOEBU2gwhyyOO41v
XtzOuESZEMHFYcUt+3GkqU38kumTvuRdq0WwHlhuGIT35Tr+tNORxRe4HT22BLHL
SkQvAqCc02FztJjwSkxq5lz36R62Dq0fcspVMgIHFjXKDaKk1VZ077CwfXvmX4hT
u5V1b+N5fZiKF1DJ/D4tVN8O9aY7EQkqh2yC07kZgls1/63xu1aDfXjLSaVFsxxN
Vy9Frz9C4908ppc7Wra6ZO0zkPCT5uwzkFf9sN1N/D3KRbkCzrz0bc3XBTFdlf89
kIgyBiRxaFuBMY7fiwROJH9/iTCfCWqy67iUWXurqRlbT4ok8D1EXxs2rimncURY
Sg4JYIWAgNSACigbe2YOPFBqrKkU2Ad6Y0abQ7LCfbhMGdRqOjtWBVnVOFSwJ1wh
N5blh5xTQyqD9Aeur5oMzjwACYNOdxK9OKtKj/NDZJ8yBmJt+0P1kyWBlcV/1w74
Tkvuhph34i27zBYbEms3Ttnpyr93ufWHiIZrWft+D87FreQ2vyn9Pzt7NN+86/uy
H2yMfdHkA50RgWiT6XYqE76+B2P8EXabBvC6Qn6mK/uRFW0hfGuWnxXIoIS/B9o8
B42FVqjrubPjYBvTB/qk881Bb7ekrgTJSdwqofCpiwXuAgDMeGR7uPxVB7lTRk2u
zzEzZyN/mioB631n6JvsTz/9a+ddQQ8QefrWa/qNUFMEKiyPmovQFOrwnmDUHB9R
m6LfgLi44qifker0C83a2Ww/9sa0zx+K30C0WC0si9J+RUAyrsGQMuh1TRT6luH2
ClsDdoDvQUPJxiYW40Nw/Byy4Ax0YeymPJoBxzHh/AQUqHdVhwbJe8dx52eENzY5
RWHM+KoPcrvpA7QdMY1VL1Z2xHn6VZimmfts/+f9THksvUcXbZjQ9HJFmvbAnjaL
Bz7VrR6ugsTbXghOJYtUd7pQp/TE6WCdhWduz+BJbOX7Q6Ps47AJvyAsI2w/6Cn7
UHv45vGzStrGJtElloSLuhkdV1gRfCq84Xj3pfJ5H/tnFnpfdP/Y7LeTOWI0GiYU
bWAfAFDVwLTsG9y3EP0IHnrOFYf/+aaKkED+vVFwhPGLTtF5N9nFsQGGxgI/2YkN
8fBVpR9zH66tPRtytjkwsSmaZD5v+N9DjpkHF9mYgHXB9aiabFB5SFtOdJMilbHl
kx19W9XkEY4gjol59SSzmFeYbIsX/Ajq5BuF5oZ47f4rU7qeQHElN5t7BKmgqVmc
FDKlrgLzpferISeebvqKjzF1i8Uya8hFbBkK2UK8u/CGfx0hzz7cXmztVaW3saC6
hXFDFsj1RwV6t0bY+XDmDTznSHdDHQ6+ynCfaXxd5KzFSJbTsKZZplSputITyNwW
tmvbvlSdFzoj5BphRQK+BA4ZXKdtyMN7YRNcwj0/MLsJd/qjT9FQB6FKUS4ZQcVX
JiCpKbeoj/FrOU9wxfezbtt6Ov8xHMRB9UvwfxEVx50oQXTOkA1HuA3AwT5Jyfd0
ebkxY7Yqz1C+UIr+L7d715jTZ/7vjtr9ygQ47r8Lx0Pz74lSGbsKI3GM4KB+MUMY
aFgr0UwgR9tG6Uk0fG4036zGtyjEPz+dBLy0L7DOzDjZ3hZQ5IrWRwWcT9g6VDrU
08ifsVdsdFVRCKyc9Qw3ivfyY4MY11YjDle9Mhv7SVxyx8dCZrQuMI3AXSQinbDR
bFMYsSKDoqR5jjVZCHgKwJZdxcnM6ho5+v/7f5tdzzqZ833PiTFtev9FmMROy0OJ
1pumYIhIhlcigHN8WeX67PGYedk5GI740td1wjdcp/xyGGTz/L6jFbx/V7VOtkDb
RHxq8Q9MJ4+cbjMfbLhXkRh0vaB7JVERxJD9oMucwaiQv2Djs1XeZ8j7P5Lcc3N1
XFy4mFNJpgPNpKitVuCHmB8/FZvq6FXSLNclbCbLecSmvxL41tb+mAcKbmCbEEbC
lLWw/aPRpQYusuXJ9DqGKCpa/bhQOeeUFoEdrVZGxn57PofAg0mmBvNUjdNpBLbR
ymMqtQodPvgFYgNSKGbuBJbvEARgndid3LgpWMtmn9s6n1Hi8iO5Hxd5kx8m9Aik
O+FHX0E4KovJsNHHAEB+4dz3bYxgjnOOHS4D5dB5I5DSPXNGfa2Qfr/vkK86JJKc
0p1zXYCRYtpqEbVoVnum2YhKpajN0hTAMj8wowYEO+b44bSk5K3eRj7fPb5dniK1
eSV+ZBlFR0e9tRZRHC0rOSYDbprl89pZu3RUWKOA3NUsbfc0mbjH4QjmAd90nqiN
1devXj+BciFmNf5Iga2bFvgxBPJUehEwHpNnWFe89dE+afW9LfRVbKus0ycU5Sn4
rS0j8UGdDybeF1TSmz1BhstsG1t2rwyxkqeWS1CBl9I3opmYM+mTxNqih1VrioyV
kHMzWpihmUQKpLJsx0Ur+DjlV+4nGji3nLAD8yYLmJfr9D6UfQ5ffTmbzt9mfRfV
m8Wan3AJwNiJbtTKDbMWbjkQmP56h9ftd6zVBHir1virFFGy0swHpomQNgLzQk9t
IvpYFkRG5gHBeWsg3fGqMc14okX8IBDMb/lh8kDKT1Y9pWN3IbI8V263viifDAAS
g8toSRtvi/3++I9qBngMwIdOo+q50aj0r/fsUFSR1W69ErW1LvyXIzpKSSrzn+Ep
mWSWQJZAuyjZDvvTiR1bvQCrpN6ZcmeKTi1PMz1cRkBDJqg9q4njXF2FCqQI0OgL
lBMZ8M71evqX5lOiojyEbCP9+ALdtPZfnwIh/+QzVIlzZYbXvzGPXQPdTHxWQ3x2
6kHO+TdP3LuRRAfACH204EGrX2+AZxY9ZEmKh6AYo0OGQexma9pwhSF1yUhuLe7j
JTWU/a5tvV/JCYAt97sLkd1cbZEZdfIZU4y/SsVwa5x+wKJ93OFIwYwUKZlEouA+
1itjYUZb92VLBXdUU5JoMlZwKz5EHTKlHkk/LSXCBDZkQEd/louL5p5Pxl7Glopq
2upANKa8MxG0BR/87Lru6ZJQ34aIyOY1R8c18I0Xk5IIjQawbcgDgCHDnaBWJHfC
jFy8bSAaKFj7qBLLU9Q6inFon+ugMS+jnjgJ6H80TVBDfBTMqRjHQK3hHpjQh7mo
HTZlaihGK/iBpEikW2ChwfOM7DcIYdT/KxB7eZJ4otsFskceu/WAr/OE3qrns4nX
5eFQyKDE62XHXMtVCezl4WxQwpa9ttDDjlx9hhQ5gEJdJqV6obvJ+SR/7B1hBSTI
1MKptSLDuR6NZ6zwzqQOPo+mlis1DYuQuKPFPoXEfbcx6y8uxNdAAaliE0QlAqZK
saShpa4YJcosi+MjxW9I9sr2aj0o+53+caPof3TVmdSLQYS8qVJ7Wx9bGpjDg3q5
SOMbY977VM+QSJ1vJZfvpH8VFd0QkLlG4U7ZqVKOPp0hGZ6Xetjb8KSiPwHvc8x8
Tbgm85LB5RGvf7vcQJm/vtlklPXStMZrP5v5ooD3DFiqlJAEICq+D74ldCqV9WPO
LG1wXoBgqN61t5VbCigDvPF4Ng4fOSuBeBruy/TuTxqYVIh7dge+DmyZw8Y0MRNP
sfW1g7U0YYwLLyrD30LeSIE0utBra+jSRKXEuc2ZZalkmSJW1sxt7lhso20NqUjj
bH0LzWl9MbtchunvC8A5n0zboSdl5AhcgrIWgQU05HQFz4Rr8wvycITgKnP+5fVx
3Iv2UBsV0EvkORKP6RAAul71/Uh576trdXBewvBZg3npVvUn/T6SYTPjQG8GOHP5
4HAdprBMAJ6MIudep9L6xolvA99yTrBdRX6D3REHdo/7TQmAQ/gGf8xh1AjB5fgc
JHdggWsPt+pM5cBpkrq4JbINjf8CpwBi1KyMfg/2aNJb1Gg6mR9O8FS4CyUHM/lI
cfG4BWC5WRn/xt6MGUNkNZwvpyJWsMg+yxG0P80yRdoXBjsv0iPwFwZo+T5Ff0wN
E9NhJMgdhGlLuriy24Y+rtDOlZIRtRaJLGWlVBzPqgizMC23Bn5xFa52i+bpiDs/
u+KKnqqqyUB57gPh6BOvTx5CziiOZju6bB2CeNDFYyIPmBDPsN9nsiBge/PUIp1A
Rn+29GjCeZV7WQ37w2bqGJ1HjLnN4XBVYkCLCEswKSHP4SWZvLYT3CMpIBegflqe
A8NKTsfK2U85Dcsk7LGtwuCejjHtUlTmue0hnbHtGHbPKG0CVmF9drENUZoVyAAW
96YP1hOr6nMg9mQS3tMFAMN+f5YXjH+9VgUJpb4ep4ZPt9p6AOW3Jhp4mHL1ejd3
gHYvjyrIOrjh67ynUBDIT/cN/xzyMOMkmWTqZFE/awZLXKYIr5509/k7z8v+t1gU
J50h39kYmVpsJzL95m+LBp1KAZL7CeXd6kjnlBAMKT/74Hrer0yiPE+5shsup8g6
XF3sSiAIAIkCGKk+zcAjy0KFUySjSZRte4KbOUBu3diNtt6WPb1gp1eJkD3cPwIx
GX4UpzgLSBHfnRcb3H2wOCmClO/KVFGz0/Ujtu5thyAYGHq6fzoNzapA5Og0i6O1
M5gxfUIJ2DjdckbjQ7vVzAux2uuOi6VcPe9MKqxMXCxR/f+fD63hdv7Jf0vgteUd
L0Gkgvr1E1+9eu1uDvDfLRf0NKDN7zJVrixghWScdsVkf/Vq8C5au2HpHhbxveZs
ytdnscmfO5BTqJXUHn0u6OfT8FTS+iG+tUGPiKyzzS+M5g1nOV3EPDlYVYvjQdex
fj76xSdpxO4j4ceIc+oaoSmyrG1TeF6V3sKk2OdV1WWgL4CydxKzm/bQu0ZG8DGg
NPdQhN92BkxfjCyuVxhWFYuBk0Q9IiXvjeoytJsVOb+FwnVhdQ9QtQJNLVWV11Od
IGhhGvmP+hYIsIxl5IyIiRLxZNb4XqYCzEnhTTfRBO+VxCegeO4ybDcVkUItI5SM
b0xTRhyWi+6l4lM8rZ7fOXb7PojBwGbOXdOkTT9/lwBvyEbQ+NKdD4iYTGVUbHu/
80fsED9B16f74MRAXx3zvpf9WU+PLkZ/yIlhm+Ee3w65TfPEydPuTXZ3AYspX9QU
Tx3f+fZ3/TovL+c/FF++GLw1CIS5i26SgZZV7MQxrZ+pwNCN2WPSl5YO3bJ48QXv
hMRQDSS48GNr01/+eqSKoI2fM6f4jpBzH72gEhl5vlmyJypx/VPegsYMwTtTIORn
QPW0dbK82kYsndXWFBd7FdetH/XeGK/BkbOWSssqqSMnlT9W1/UdVIY6BvGHcYiH
i4aKmsBFkDZ+g48akwSvjkhMlEG95gRt+3Ld39Ae+T8BTPt1RrTq/ko487KKObm2
KgisPSfTBeMIHhfHSaZ0oiuYZMPOZYNwkBqamy3C9cSbiJCaYQ/PD6soehbQpjhp
9ChfAA9Lb2B6D+4FpUpiJM6jEnLTVO/fAgOfKUnqXUHT4XJy4X/HtPozoQkkHwjj
S6vTPXE2FG555kfNPZ/3GW51stgPmmX+IJ7do3mTEx+oUTce79fp/4zN3qs2I9nB
GwX88z5v+A4nqivHqNM0i5Pjobvqq6+5gyNR2c+0OgiTLSLHQra8g5hDVLQEtXtj
n0QpgsxXdOBNaWWrcPsDt3+1oUaFOLgYP/qvtg+eaP0HKXtZ6A8A89LF1DoVrwdZ
yAxG7vkDK8xQiKbx6m/w+YcJ7CRVEPGG+Gjjc/xCjhChsVoAD20bTTMHigt0zaXW
k2YccRECxFLHpGfKDkLGLRegckGQE8vJdAKKiEdvDqEe8s3niRW5MbKhmn2rxLV3
HqsL3pkUnVMMw+ILccsasmHOJ6fw81UMdYgQyp5B7jpxf245deJxI1pXuMxjjQy5
9zvdgAGPG/8DpnVctuA4HU2667jf6EclaATfTtnYCEgvau5MgWTQmCj3ovwSkrEO
Ykbh4X6MX0hOg159onBoJQed/MsD0cjdVpkak73IUUbjOLVddFw78YxPOxz9dBRP
J/JwfAt1SRpgtrH6u6Wxp+2zutpy6FoYQZ6GJSVjC49nobHJjIBf1BezDfb0bpjm
+QpdAnvkwIkCN97XKYZQsBCKHP7vidfHw2RYRAPNvU9yQsyIHwAaOeSmji9e76sc
jx69rsYdlXF23n8D0lsTjgY21OFo54ypQ5pkSuX5FUBznsil+5/QiWhY3EjyQnR0
1N+cy51BYMhjCBLwIdCwzlBURSyDv2IWdQoxmf0z0wXevJNu8tf96/j3ZH2Ekmif
/DMjwDwAgF5o+n6+5GZjED8bHczmfAPpcOZu5lJzo0hJxQd5diR8sZk6PA7/ZqFn
RgG7SYpIHSK1H28Ia35wpU8ZknhNY7/l3oCM1TJGg7iPZ9KB45lLfLq+P6TWaDUV
9kg0dBLhsm5Y3kthSqJDKGg+RY1NZiXtRDum+62OLS7JmEXz3IWEsNfkL8bxy9fe
b520Ds5pdJ28+PShteCQYwPeUMpw1z8qVlus/T+ZaW14/G8gAD/YJTTn0ZaBF40p
Gfc28HjJ5cGB6dNJBP6C9xqMQ8Mj/tGYAiomK3oDhF5mPErccv43kIxd+PoCXq7Q
r75ftRs/qxvhvOTSgU5SNA0/N0LSxFeJs8sl4F73FNAek1bDJK9G9nPj+Lhh2CSD
n/S4oqeaN7i8QL26ODW8S/ykp1ainQzSB0+PQo+34Ym0ePz+5qqjBXQRouDLiqYc
b17voO5D8a+m9+Z1p1VGCjsOQ97/oJ/Ci20/DhkMRkU2SC6u+nxoEYXDM0700FtE
i4TxH09XUwYG6uGx2cM3dct9RU63fzwwdrE3ytOhqc15TCEGReUqS+spD2GkB8K4
NcpgXN9ZrkFb6OluGZog+WEaiUFoUgu8CIXOTveq2o1Y6p0CcA2f5Zw105PdXIds
y5VzOT9hVdsPajW/Ie0xjOt1lVm9ufEDF2OspvA+/WbYAB3OFvnd06ERjyNXJs2W
pGBLDgQgL93pZgE/b6DzlDgBhUdYwWXDY5b8rwsqXQ/zAmeFoTsWKtBvR/1kzYWR
8Zdszg/3Wbuqy1IShCr8Wc8qnfhj3EMeLv7Rttv7HuAM4WAQD6cATX9NYPNqoDTH
tw/pKYh/TyyQxx6SDjav/IwS0hGLJ1Pz/eB3t2OlObiC4PiXBi6V1xqicpX62zFj
d18pnsU7EWu772PlwLUCxSYiQrbFtdXHC4aNVoOdaaA2W6BbNmdZxP+5Icl3i3oZ
vAXGfhvKzH45o9xd6JzKYhI5dVGlV1aFoe1as79y2ZvW7xWVgqkzjOzo+QBhO9Xk
LrnDRbtHtfIU8R3U8jAPpSy5MOFca8F8KqhNaU5/eQPmQP3So/CfLRjhIFmifdNI
HVUI4v5wfKerbDKheNIUafNdIujJQsoFVWPlolqVIs5A5r8xuBYIWvHhXWsZ9uV2
a0uhpP8aNje8efxQzDySfBp63uZobvgOxOB60UKPLVKVNpzN/evMNdthMamVkDsN
+iyHeLvbpP8tr3TwzfIdgR81oPJhJq7h4HNNKuAg7Mstg1rux5O3cgsG+Ea/MZxg
uOfwMLxQk5K/ap3Jx6AnJOgWRLUU5MVd14QETqd7R9uByEUK6uHaMdXGdhuRy93Y
q2JAegxB8Kcy2IOkejr1m1kP9arEVzzkH+5QWsXXrwfCmmDgYit14+ZWHX1Fq6hU
wIKhaPOY3TO2O2nSYFTfkUkJAAbaQHHm1lVrigj/nJnvBV5q8ld11nxnsDvsQq+D
F4sugncnEo1XJDtm5A5QSpAGSPqrXbT0bql/WXaTkiZQCMz519rOKC6z8UJ+Ldy9
uB6ul2fR2moS1uoxkk3COfpWi3ADU5J0HA90LQhugcwl+hj36pDqn+YFrjUQlxwD
zw3pJ5LNyWClzJWIqpUDKrlCkua4Q9WYVKZzV3uw6FEzhE8yWfYAg4AZyUCULuFC
iVFDFxtoekKVhzNGqvOcv/N7X0fi3hyhCrr3PX7M0XsGeLlWXyp9UvthFCKFAcr0
Mi8wGN6aNsoLvm3i0+iql3GZ15XaUawH0fh1teM4GeR65UcMVYZrB2tkX7isH3Fx
HGFPPst2dvRwWrPm1Xmwv8+Rd+e/VvOeTzA0Efm+9deVlYZHL8zi3v5u9GanhO1t
2gwQO20Ml8ZNmNBQuS9qWzpBGUgDVCxblre3tOilFsscXLyyL9drYVzegfKgbAnm
EAxIhyp9AS0vmrNejnq15Aj4wl/xYzyVKNoIsppfIkRt9NyzZp5JPWXcwxBMZWJi
RDNP7WvalOypRpB1VkRJdqoxvshO6mn8bmnhJE+5ihf4aXDY1+VYs2QQ9mVmlUQM
BCclM1RbI3pMPMCeIU6Asob4WksF8sllEClvRSN4Wz5tC0/GoT8eh6YpXZ1pq9KK
W8FdSXiXzbmndQng3RR6YvmdzcvMInGM2eFdeTH3WGJJiW4dmKvaErBFSXFAZ1/1
L4VOKazjgmK0rtdOhF6glIqRlTRlHDhysotajo4GwR//2pARR2d9DPJiReqxqGI6
4g+zyppDe2KNgL2IeF1jxnO6VT+hSWHpYES0evvXGbPm4kMu8ahT5yYnR+OvUwb5
zWA4qcNRHR++fvAsT4fSwmYDADiioRJI8HXCvqBfwTVtn9jQHzH1O657OrsRASyo
wKgWLExdrZQFXtSQDFe88hzdPhq3Wf+J15myEXBXUYH7HZZ8z+3wN2tJD2u/QjCz
K8WO6RqgS5zA3K+1LCp+I3IwaBytPKkma7xSoLWB4hAbMBq3/LWH5uDdY3b/TOis
jCSN9rHnJIbmInrK66BK4o3ulWDTA1jSVwnk5SNILtLSWvFnKIdBJER33MfH8wOe
7bmeVvPdJgeh6OCxwVX2p7C3zEWKOKXwCYt+CylPZmKcMwvyw2HIcvtFuCxra8tU
QX5gYtd+zepJLfDBuh1bYNQAiCVIvemGT5BEP17DMRomNftDs6B7BtmfLRV3/ek5
U7rIZtpX5VQrqjPQ+dvN9G8wiU1VpVx/xSzLeA6Lu6gd9N+tP2p+4aDGn6goirMf
iEbh0gcNir2A60FYG3s21c1NQacs1PWysd/1O7HA5gsATcWC9m4kt3wnp2HF6ZuU
EtNWq/2/Km4F/0pWWywtaYRXw7OMhMV2SDqnimA1HAYKR4FsE4a9pQQTx3hAbv4B
ZzuVwTrtyO5Zp3Ezr05tw+d505kw8K8+hAzkuZ28ljdnS9ddhesMu3c1cJSD9515
7fYNDkBeNWJV+ImtE+I8f14mQnWWr25bo18liztRqMmD2oOcaES8CFQswCyoDWfE
dolWZ9ikgRjbt+eERn2ptb6wrghMGZ5I1GFEADc6Ggwf50gJ6QFy3eYE3vRA7eY3
tELpkCvfCtOlpfWlDvucV7Win/NIqyL42U+/5cZ6hg9NZ/O+fMxW2zMnSVMZJvdC
KddSSFzKSQFj/r4FiGCy3CpDkFLBczEDyL94pqbM4HURhWGILe4yPIGSfLLi/VU/
f96OQ45HpPugZO+Mk4yGygIRsWuP2adnpgpzsmPeuySDBvBZm7LbTjGbVxoRsUc4
SqvL3AonqHGWP827POwTZifKbLftzIsingIZYY5fxWp26u3++HiHIQDA5OfxTBxb
i4Of1HbJrwK+XGMkbisL+vpDs5r0YaDnmcDI1VmYK2iNP2ypPtekeBFSLKCyQN9+
bzkwJ+u/dmye1GA9a21PyQTf3NsRBBkHNOS9cBWV4T5CMKFNiiIqi8zgCje/8RCQ
qDX2rzb9ELWNFXt4/zjtEa5Jfle12Ay8/15+n/sIfuQfwsOhZ/+0M48GXPO1tqI5
aFA8BkHWhdRkD1bE95c+w14K+RYRhyeMidHW3l3jpvSHhIowPQxswA4xO7tk9qTI
w8rJgVbIKcmNnZxym8O8qrTO50NWiXF90nUVwlTPvG8vwv4Kq2LSPZMurdkOeLfT
0/HQWCCkil/5BIttzpDR3tNfLywEZzMdyVD+JP9HX2+zQ8oQIXcshLQGlF/2cbud
8lpsVRSJeKDRQvaf3+o4RXlDN5irhVwy9D9O13sGKj8PKrn2ihWhqgAw7r0dHVwL
sH7RBr0zX/rqWgyUCHSk3wHVWKdHp4axELQPtm6BzndlEXtOnbJM8ggka7iJ2Rht
5On2n3Hx8oY2oZq8k5tzruS0FrjAWONEPgzsrMcf3tycq/2+7HxT+6He35g5ZNQR
n3EtWymLo1cM/fGZvXraWMuWJeSaZGsuwu0jcF1QhT+mYELmJg/4niD33wwj+5lJ
LkPgg21RsY3jFanPnuvkCMOyMP6RCgqafHViOgFB7/AlgSLILD3M4IEMSFYQ8Pjz
qO+VrprMPM1v9LPZktshmKOzWAlMj3ghsTEUCE6TLgg1uk2ymioaYt3Y5AKyHU0E
f8EyAGw1JojfmQS4ARFec63+eRYPeR2YSpvOm+uXjqnqDXw27sT/rF4jOdvGWwsX
Lrp0pleaoVzRDSK9Rmiic1ZKoAs4nCau7FsUAX1J0Rb6uoSdmITgZ5H3SbTAxmX3
SDz68bLzgsvlWFx1ZLy9/OQvTsHTrj7vk0xxREvWv5VMnOOzsz27/ShjC1q9uiy+
wCUr5q04aXtOOmemsb1tEjtyJShxpM0tRNtngjzlpENuAqNPUr3t7SXZwt59cSgF
6pHi6G2TksnVw2MqeEMJKiIDBuONiBq6/gel6FimAfZt7KiqG6FuE5c4y1S2V8Tv
FVhzxNA1dMX5y+kDxWNFhmUgYriyh7qbvlFsIo20/ZOZmoc1K6sbkhjdjW8ew5nA
OWauODzZYtlWcSIMfB0ZjNY/Q9YSVY9Eu/jtONlAA5YjjV4xDrDtjtRNchvBgi0c
B00ly1nWL/jM8+d7oriC34e+bNWi9bPaa8+sxe1xbvMzS6j1E1UgPDcLLyH9FDRW
nySTi4qZTgr5lOUOF/Yt3ymgz23oOYN/TQYg+JaoUC01cMqrR5ginz6l3WZ1BCDf
KzhJobYWQQE4/mkCfwmTz1h211CXbRiI+RSLVrF+hePXmr68MFpgppqH3PPfLtAO
5JgJw3isNrbEoC1+2/0m71A4HLopgJAd8F5bijk82wcDKM8xKpmJ+zK4QEFY7ATb
F8f5vjT7yI4ikEuHx2ubAWWRWZIqn0a2oyfeo3oyhgYHbu0icNECNVNAO8iaMh0j
CRxdmEN3z3+6vKa3rjywdiHKsNR+nGF0sYroGCs6jIkLnOKB/d6MtNryhptlVfrk
ibxDEu6baRKprNsUA76CMfVt5dJ2P5LI+QsoaTZaPU9fGNCZ0UOviEZghOyxJyfp
FX8isJX/ZxMloG/TxDf6RXmTwvwGMS0YDpeH2+sSuhkbjHueWwgUkFcAlnhe9+OP
2QMhV89n4yfG0m8yyO76avFY4QCDv1MyF3Av1GjS5at9B1lPpu2fsxT8weLHel8M
m4kbmYI5DaJARClLZv7CATOV/GSt3Ex9TTImuFPjA16QqGdNm9H6pWCUDLTglCQo
a0ImcjAcsEuQ0AZohNVgG6C1qJnwIkLuDpDQbK5o6PBOyYkaET+sKIugCwrHBHQe
BId+E28VCCh4t4ZUyc2iv4OS0MB+qmTNbX+1Tq+/KLdSb2XylxObOLX3MGGQnE3T
JIX/irNWq/8fpXyF8zc9KhzEcruEw22yAprfUNJbAVEn+mLe4InxHEgNDj9rnHiB
VVq853/LPcXSjdXE76ycMW9cmvqLeE+1QiAgtnel5bKPi1wbu8SBG5y6TWjD7OkV
4AzWBLMJ71us9W6ED5tAwX7wYeaYdROFdCjrmPZBTG8+Y3RZ3WWOdY1zXP7HCSi1
E259QGvoefbJENoXFNZVy7iwzNeGYm+3Tdec6hlZwok10/xcegKPxXHA5J12S9U1
w1YtmOTPvV27JzZVVPDomFhIGNDYPFmSTvdqMhnp3NOkJ3mNGWZmkqmyuPqhcQ+5
K/fuFATdmVcycSHRYJsqWjBXlA8IhRfj7iW72chOZ5U0T5gTlm1Mt2PkbdpEd3ZX
MnQuVMkMelV5NDVFAunUlcwBbdcJBNc23hBR9qfYUCEvXXAyfFwbzxQhp2O08H3Y
nVE3JFYO1IexKnCI84xNBNvAwO+5CjImmeumBhtU+09RdFSWR2gcU8xFOONIpXco
e/bGSAkvpW4YomZiPHjZ7w7A2pvr434MCqByTRW8DsgBWHFnpGEDWWXvfb4tEGVu
panSOotcSiZNyn7Wx2YPyqIMlLb5nyQCau5/KaAfydBo3Idx/vNtWV9JOGjfO/Z2
ozoAFhUxFzWINc3Whq3/BoNxIhNSQ7E5nRaHdoBqUG68zQ+bk8Au9kyhwDrMn+2R
oTlJLh8eRefoQOXmESiYIje6BVMySAl1i7ejZnW9Oj5Bw74kDeWJzMb6jtWyRFxm
sIHMaDf7QipI/20GL9KOulzFCE+wWUB5Lxz5ygO5zPGnKLdJuyS+MV33nkBqqTBa
gtHdxPw0z0fhIt6vFFbeG7oexncn8DMh8DDMKzT3C6jWpQcvYbgoEXHMeB2fpsgt
AJZ1fYSBm2mWgnqicu3TyfIyU+SxuZF0G5dbURV3Jfq8cDzKTYFKA4KI0py8zh3f
H5vSx5HSEg1mXNv/V/e31w0+W8EHqujAHVgR7lAFjng1BK/Gu1wtIfRqpD1AWhn0
DiEb9xsCoeD1czBN+p7iKB4VTPJ27wj2N3N6g6WtucpI1VuqWjmyau/HK+ElARaS
3JkpL4qhQo38+tR2PWLQTJdO6FlaTCy5RqcV0MeMYgbsMNu/1hZFXaCEu3J9WTqp
/Ar2IvbVXtxNNWdYKU0c+iNRdNDhZ7qVBhFjrsnJlCorFTo8hkbw3PGOJe7nLhdv
xCVeKZpauxDRHeITYw/zaLcg4clNuuzWw526+oqjRmuJfHGwWM9nRTp7rYFNq6ml
S6r74CEx3I5VuhnLebHoBMCgHc/J4uvoZ/VUJvkadm0p1HHuq6flRvrLAC7lMBpx
nR/qa7JTC9m9CjlRht4BtPGwcPIUHrvxOr1mBvYPMx3OWGX9glXtHBtlFNT3IPHY
+i6agoUaoWnL5QJvy3Cg2WQFpnHbTL7eV4hlEB8uskcCtlnm7I2xKjCoNYhNbLTG
VYbqls6Dn7xS0R4hc2J7q5dacrn67DE6AfJh6KGwo7VeaE4fsUPnHjCmWQD3k20W
nN6QGYUg74smgeDlGgtFtx3n0eCE4i+d8H4+uq0BLVuDPmASbGF8y+Gt4KHielTw
8l/ZAtBVKvelZLiVW2n5A5sq+hAu9ykBcWtRRI3CS1Edyx2EKJvngsNP6/6SbCWT
DuQ4Q8wKczHEh5w50PCIUCKlpyTwwAxJ/fDPNYvqIK+VHemJHcfAhhxvAQe1TwpM
9CHQlUyHC7O3mNrEDmDktDVl8F7yNhXpGIjCSFH5Nh0B7UWOLfez/GDW+fmJj0QS
/U4rjb/yNFCvEQlN4qvVJwaeD9qSNKENsruH1OVlZbzMUl8CA20jy27gbNkm1zCX
inxUrSOIPp/8N3itikSpOoeoGcJ5dKneqfcOdc6u935TIwKCVoXgvnwWdRonfABD
eArmKHcftId/m6Sj+QMAGgR/AQdSPbPideHVGDRBKJv0xSUeNkjpXyZ98972vDXR
Iv3s1SisAklv1hsRjs/RdPJ1VQbGKfI6+ssGm3+FYI7qSD9yG8nmsYIkq1uK2fiG
pdGMQVwQ98inMiwnYzHEFz3B/0B3aEtiNNxGQvhBKd3ax8bZlfvKZBVlOzS3bbGf
2w9m2BytagEO10fnmUkQY5PM6e2FseDlWh7IZe012yJq/UFmxS4DAttP7lGzk41m
PUKghG5gpEhM6xbw3FHDO24iejbHD8OELzAdYjsVZDrHop+yeXDITWDAwA95tkeZ
8SJN6UODnJYoYJ005W9LxT+V365AC2tnD7I7YTXXIky/Odf1iHsnkxlb5xZkxdrL
hcZgky1fljE9ge3ujuwGSEd4ro0RRIZmzQDu4z/4l55K6COHZDodoUuihCcBG+E3
8MJbkAv5hYQCrC8G7inNpwnU7LYX2NLjUoLLuJ8BOXL00MReGK+L67WeVqrFi6f7
t871ZK0jN+ajM2+jy3hcQb8KjsTbbyjjiwmwvDpJkXbMYFob19EwvizigXYIws6I
0VIlopxUSBAMYezrq7cDjgQh7gfiJFUOuVj29EsoDxzETsm1G6mzCkUSbGLvIA99
7CqhMZA6wsMYq8p//4kkTckgClFSzMt6VUIWztPp5VuoSyxSRL5SejyWGg0ISEbS
S6sYqqg1t4JbS8vmgzsBb+y6+qCDfyiqn6q6nzwDF2SJx997rSb1huie+/Zb/PTI
QuX+CaWfswHimmDD+eNisFKJQRaN8IZXJL1WMygXHswcOYqCPb75FXoLfEgcG8ZX
Sg23DC5UGynqmVEGRxie5hP9LdbRDPNQpVspxt6KTZ9PZwIGF5LogjB14l/WKfp1
uJKgVVYHlZGWoWynX5f16U+kksJA/nxtGCIX1+sSx+5LRCUY+VcYPllIeOCoKJRU
cE+CXVu7ZPzwFTDCbnYwqiEVtqEiIBc21RDx8S3XwHi7y7uv5xdbkclvCApCy+E7
mCuERg77onMD6ya7Q8TRjGiOedzuf/QBKx08Ts9V+zzzxBEjPel+p4rsqTfbzF3x
spT1WO6fqEH5CW4Dteq6J1gpLKS/KLvldMmb6EzRihozxlaHkyZdhCQcRA1EcGLr
pfQkhT82khOF4dtKDiaYLUCK3ERk44WJPpjCRYWpqAiVLSTczL9YSbVRfG604DS5
G3+hBQJFh1Koda0l6lSFHNsk4Ty9BU/oR9e6buDQQ8rMLSyqI/UjzS3EfpsMjYYH
UHDVPnjCr+ZD4CI5A4CR7JQurSpJCp7Kg2wHTygS8PrND+lodklVssq/FTxKQ4Iv
HTJx3VLRt2HTkMzxXxS1wBeHoaCcubhveMArVtVpoQS5wV/NTZ1jC+jLjjv6iNZI
AkpvkXsB8aeIWUSyrke4t6i/eMTlde8p80lgU40d2IHDUMapQ2Vd9qe5/y0qeHhz
C1T4jZnmqv+vYerBc7BWi7lEfyQIL2/jY3CExjB3x/viGCCFVsQm0PB9J5bBFWdV
ykPA4cryvlUAw6rG9y4KlG4P5FPg0jDq76KReHjiuz7mFxkcCAIXQ6h9f4SXavjS
wNRdiRIfr1s1k9Hro9YiP0aOlNl6rN8frR33YtkUU9OEZXkBoOLJZV7ETgsvw0ze
Rs45tgla/sCZfGZeWjiWxIlOLKEJMf57a00ahMJOYGA997DG46/3j/3cbPQLyllK
Wy2J6GpvTAM4j4Jq4+kwWZU2SVfXLL90ZhpRTqhKaIB1qmDygbu981XI1+27gEs4
SYJZz+fi9+H8JX/VkPQ/lepe+dyr/B3xNy4mujEXk+yN3/GXb0ksZBH3+r63WpMZ
bz3KCNI1Q5UvRQAwTYPCO5IH//pY4uWJONgx1fRLapXEBaGWvVb/+oOPu0VeTQJB
5Knis8gr4yl2HkKH4ze0l0H+mcNYC4LaHLpwRuG3fpyefObo6GVuaqxHtc0EtYAC
flZb+wIgOIu1TFWyizLJ0ynz4hdWJc8fK7/AD6f9SF33+6A3DvorjcaqC5vjKO9q
Z+DS7/W7ucOIl7/wSGu3tHjaiWTIZHiRqn72ynm2v/ty7x50hQnskOFleoYh643g
aZPpUvMpHGMVtcTP5WYe2ngWldqH3XRgUoTHJAGoWN6n1M1MJHKiKOjzh2i5Taw9
6Ten93RmNOcq1ESNkGEIHbVRUwfQiMPP11v55YG+8o8TRM3zpTrmkZ3nF3B9Q4D9
IKe/aBaeh6pA8gC5YKF+TsJBr3ruXxaqDp3YVhQKWgVQlHJDC1uTd+60pv6Xtu/Q
ZXKxQ++1C7nw0A76/J58SwkKQv4uJLe2SLGeLjrHGINsNnxUoV1jzbhef8+Tmqh1
8M0lwFLLKJNnBb+z7AptNOLG5bmKiu8QYtGEZc+YgukA+KNqXm2TK01iN0K43Z4d
8Tg4Az9fqkpWHTG1nsARZDrSmrJOS2zx7ytKHyx72Y2K9v9ACdnj5zyaLAGx9nmK
iLrOYVOb8BWVhW8ScOFAR3pkMh7CtBDWrp8Uykut66hrqR3akvSYefII2AJnrbrZ
7P7GXWMT9USxV/uG7HNke0xaWkVz3wG84vRUH/zx6Upwd+58zGgZNvkvImnn4aPQ
RAlTi93AiSU1Ip4F5czbGOiEWOkI8xfsoLWzcJVQ4ywt0YreesaVT0wxEZ43DxtY
HDUYxTdHSZMd4UMPOcB6NnJtP3QcZ4F4Bw90sM9LDFLDSQPcn/Kyrck89cVHz5z/
+NsyKb1Sc6aD/08ZYtzhzLHKWbawD9bR3QpsLXXKfVxQlqnDm7pPCQ27DYAZspD/
JkO0MArE6Ea8X/FOdMshHcaPMMOPCmBKgClNmqGBPMtBXmn2Ne3OrLKd76H24mui
ddJAX274qmSw6hzgczo7zLMuA6B0UZ6Kwpq/xyZCfyvfdjT0HC+eFyzPA6oa7xKC
7/JrhURCRNpmMxyC+mnIgc89JIQhLrL0CtO5G0fSUqfwe6X1zZHMt5mF7bdRTzhV
n0Ndwx02lOC8/+TbPYXNbk48G6IsDcb5uc27s6e/deR2CfBkVZrK8g446xfAz2gZ
eojtHDH0G1Ez92+EMPkjj9bVy96WnOgB5LOSv2ONsxOiqLI0zNbkKW/3EaMqZVPO
e2yDG24VbAAJlrHUvNUf0ZwfBkYIOXMBmfH9jzYj+v3XLDHB58fZLkrlkk1Pd+nl
WcQCrf9IeTdVOgP0WTrGwp17bfvSCVFL3BRM/hYgFtQ5n0VpDOZerg0AdaDuYCan
3znkq79kf6UIzLvo6iBCiPAHECvFHbcNIjcDdzIHIfdSPKQad3YWlfiyf4sp3RgT
Jfu4sV2RTWYIfL19W2DeM+++sy6aKyrdMU/8iRWMI06rP1XX/pion3C7ostZcpGU
mZh+etWEiU0wHbcLEoXxoU06VgzwiylAjet/Vt8x4w407e6surxiPm3RzPtQIry9
yfv5i2SgolGqclmZal1EQzWTO6IQCJ7Gu7p6OWCpzAEYb43Z8WwVGWsk/QVRySGx
T71Wg/GcgChWh3mcvy9qawwey5k/+aW87xKl38iD/TTQS8ytPy225JOQhQWgxWyc
kr/VJ0pvSoEG4qzFyf07zWfa5elRXvE/UbsXfIeppe39gfEl4+dfrwA7cCwzk9J3
TP0+nsodwhG8WcaExDR0bO9Ujet+8P9EvuSTHJwFtjJ9a3EUmiVEa22my5copgXR
h45MaBPrzItrV/fUt5IwhxE7x92dsMrreRTFP/tUYZZLfLUu3QxT59G3KrAAr5vU
dO2pyLiZVSNF6GJ0o+9WbmzXHHsXBTBc2HjaHBZ61v1kRBz7S1LanCsyO4QX6Gbs
`pragma protect end_protected
