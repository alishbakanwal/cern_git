// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:02:09 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
kvRZw6EGyxRIo9nUjc3kF1tSLkxOA2bwXN/Sjn1SvuYQ4fcmWWovlhPghr7jue+l
eQCb+w+URQz4onznF4st3cH5nvTHibXdGUM/gcAKBmtKKyvdpZteCQYr9vnT5pKT
u1SJloQ8fvpk9+6b+1eJP4xGKt/zS8TefXDK3OXszl8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 22080)
Wkb1nUAh/KjtC0wj9dw+p0u4xhjT/ZDhTXal8lrJp5PUNdpzlWRndzatv0U5lX/y
/5/kKUjYvD26WsLjv98mTfmP+Rmhorlwb6gQfz/T+6HhNNlAdqcR9JtaRQRP0930
SjXSwvzGNuLC/wDe5Dw7CI8YvBUPMwatV/Fj81wWuRySao0lHjW1fXXTV//z9ibf
OzpPX2d7UPmyFnvBedCrXaPbx0s57lgMWXcg4Oh3YjobcGw9xmFPhQL+LqPeDDgV
g1uXQyFmGghcHNTZZA4bsdQY5UEqLs381CYaQloL4Bw9EhLgWPR7/AFvx7BEgeYK
zMmUHmI2P63pG6UCIp9J2PXSyXzxQGW9kktZydG9+hpVX5eMwObjjYGiEaGayo7q
G3de3yWtfC4cFHZ+dh7NMTIpwx6nxJXxzWOl3Qw6V1VEf95RoU5DXbqGnfweNsci
davxiCKxkMWvCZ9RGHdu5z70+SktGVIyPFdefJ5UR8aM5ULqa+ndsSQTj4LZ8eVz
mOFBnyb42K2Ws8Ne+HnGHd/gjseXFzb2VQWnvKclmYkzvkgDHZo1usJcKLS4V15W
Uf+sDzAMUDnxHL/Ptzk4jOdDP0kYYwik4CQj2GBrWE0M+ms87WcttkqtEy81DZnM
IXh6JjOc+D8Cbmn4c/N5e41GUf/3ShhsiWHQc3+MUXr3XArtZHGB1nQ/MAgky8nm
q9DjV5ZeHCpgqjnLcA2Yt81msL2s2jf5dljpmXLUKhOw3LoZv7fvOkGO9fM4YCav
eaHcNz9WCm1zKAK0aS3iXnei+ipmqshmHAE5vDlN5gCOyFoTkqL7v8I0kMdUs8DF
lgnuMpnkggPmklXuvXeNur2P609rDzhIrnH4o5Z5aR6JvAoFu2b9t1pdMbGRdeDD
mZ7oCzbZSxm6HzoRt1ZD022kG3BpWx3gxMj+BGx/X2BNFytVQkCcArT/hGqWdytK
VH9YAE+R9JyEWgu11fuoet1Lr4T0rZjxMPgK2DuOwd9pO1FPZvxvbeVqDDM3RnQz
qMugVLZVUhL87Km1/kxlx9aaCOs0V2Hl80bqibGCI34uDMFxOQZA4Tze77OHLc97
94EtNls9n0UvosLKOj64sPn6T8JGSYiSKgNHoqFLIO0PWnU8Cxsky7ZsHzJzCFqU
cudnMoLEzFU1pbwzPmmVLNHDDtVXhS049IRCKO/CeHPC3i4pEKB05F7lZay7XhYn
KGQgULbEAOgjOVX/9H/cP8z+ZXszp5uw7gmf2aOAMOYwL22PfdsVwPWbAXXKiVgv
t7JShkXR9wRow1x4w3pRjM5IfPfo7xkFKYYRUCe5pMuBwChqRMzRCGAMfry3EkHM
vZSAaIlUCDq9ddiPEZSbVdMBKUro8KyPERZrItwoILD67XeKNflvTJ+rgo4lpisg
RyG+30pUR/ETTt+rADSxOjhJNXdT1SCkO7i0aqAwYio/ekvyVjzsw/jUzFbd2Fcd
MZ+Bv409A35fsmylLUi9b3T490YzfvSl/yveIf/blQIuEpotOmcsYWR4U3mVpStE
IsmgCU7AP9YEwFkhyzknExUCX39J1UXZqnyExYzgn5r0aco2p+M3s3YUT8O88t5k
ZI3FXJ+d/fh9VPNjXYJs0LFlFNugu3UG3lKlZtTAidNnWWMc47dWPLj1iHa8806k
wFfmcaLEP0XutsVM0E11L9jyic7MI9DFHXPAhzEakMqVzbH0NXFUvfc+17JISYwf
ewHdafWUO2RuKOHsqFiVStQjOvG28YWy5Pm71sIyEkZcEiJ9ea1lcyWBk+gB1b5h
QaJEb3qeWarKQzEVOvmR3SRWRfukiGwoN8UnAq8RHabpnFkq5m39xU4B/xXDom/q
A7yDTCaefbzE48XZxHDRJiHuEZCbYOqvwjmb09imvKOcfmNKGIfDXqivLJyjIELv
p9/ZQN38RfFctx/5Q95WG5wegE6cbrMRyJxEZXOXWgUEAVImQwwm4Qcw8YwbfYEC
pd3tWojuFtR8aFEJY6BJSThcvoWSaFbOfmOBCQIEC5pn4JoMOCnBwD3S+SvF0dQz
zibDoOi+rUEZZ1dxD2conVydkXadLIpkNmXTTv5aXrdhcwS7GwDqkejmO7iPPL9A
lH23MdCPLeniBsRv+XM9hj45YFAVszmbt5rozJzhY/OcMjkrYwbV3f1ZMYn83j4r
Z/B5c/uPrHbWhsDCexLiuzTJPJjBw7wBnTW4GSFK5A2GUFjSXHSpRLz9ujmvp+Nq
NFgcpUw69b2vW5boBsLOaUfPjtUcBtghkhoXUY5YFfRIxXKtUY5vRVhUeN/z9av4
ltnoIgLQNlfSfz3h5rcB252nJuZvI1de8GiuyjMYvmoEZiuC5WsOIk+DIl/vZlrj
IJ/CbvA0tqESiVc2YPlG6GtptNMrFTbEArJumnIt4yluA1ISNuFlcLz13jtTeVtH
VUSXgvtpp0E9SRq3TyX1FRX4y2kBXcqTcln0HNTmXC4B0ouBi6kebPdwrElbkOB4
Dzqx5VyIGw3SZ2o4pvm4xZXdB4Gb8MVmEtrgj1jqhDLmh3R9fBA04BeXCN4qmtDs
W91Q9ZHlMxzlmzsY0SvXRlhVHev9uPvCi+lHnzUcjrO8X/N4qQWkhbzBf+tu8DgX
rNW+g0K+ibV6w5DWejLioxQbLtvNl1Mgu9eFaGEZW4+3lz8nCGQSnp5UZAFZV22x
E7OTbZKDqag5H8+AKPJlSb6YML36J49TOqNO5vGCN3kEmgHSrnGQOhDoVCz8fagL
4c6QaaiLWYb4jZQ/NFQm16bJHI5kPjeWSUjD7e4UMpoDvw00p8CPSyJBXCC2GtMK
RIuJa1eOmIaHLDNuOnmyjs+AeRdG0B13sZ51nlAOOq0oPJ0NinnSWpo+W0Yxsqgp
FJ+KO8rfSVs3sSVyVLgAUQ0eh2bIOagh914X3rpIJVLVk9p8hqn4fO41w0h6blTq
JBcWADfUUVspbM0K8Z/tBpAWQTOt5sN4J/BzJYVDfU7KFIegG9cetZ6afCEXDeh/
x7LU+PfJuGsTwaqRric4XV7YGU6NQk+OFA1sPXx9Mri2PMvGYuj8gHoogv98wlEH
7erSZ3NXGcVFRC5MH57Y8VXWpYPhUf5iwjLxce6WmvjHYmZsYikgCZDZ1upsdTUn
WlD1PPDWmhGNp1i4ztAFyOpT1ZDYpWWRMkrOS5zaj3r1h6OTbjXG1KsH41fl0DHe
xOEFVsqRy1SQIri4iitqYzL08Hlb0D2vGVGlEPMUlqjs+UwPZd/6Vw/w/IinP6c8
d5MlwmokSBUoDEvLmoGvJq892Xu7Ge1rLsXNEuNF7M6u4zRJPTODIJApWxJ+QsW1
fEDydt6Fh0tSGUXaj+K3meq+TA+fZ0nrJWnfZh3pFT5nVfTu087TQGoSu0STrAXw
88OVUKGH5Xdbq+SDFBonYm4AW5s9tPJSNW91QeW/at8ZyubuBtJCEq/Lktc8qjUM
HKKH29IdmRSelQ8dcRWXjktW4lV05BRZqGcjRVTq8VQios++h2cYXV4BKYdvbYhg
NEaFMZQCYO63fwQqu1YPZHDO3P4OpI7tnMSYNNLBTkHAARn/+bV03ZhI+n7DrfF9
5oDP8W9VGc1I154qkBpJbpaGu3fOB9Ce5zxTRJCgdOrizTNZpQBm//DcYWSGeEjZ
YGC0Rgu5zJz4D8cKDfvh8tZ5DhaF0oFlsSaVL+Xi8XP74WB81D3alz7nVU6Qlgyf
pkwGRuUy2xRy36EX7WMoHB8puS2MaURn2TyYRqxfZdE5PmLlBShY60m2j/qLfWgR
DBipDrV8YXgWGOe5cZqRHKJId0QA8dV05txZ7LiZuG79aoo/0o43yLrP6YhC0Ggy
a2hEMwr0PEiKSElAoyw1npkMGUk4FdYTWCzPU4rR6Al4dOBHiFxOfNAVDhU2wnZp
yOZC2hf3dX5OIFbeoRGYXs804lbFyLwGDA7D6oD60e/+3aloY2pXhH0kUUhBshK7
TtKwzw0XW37BgA9mYJnTy7xSo7laFV18FrImpyBLaj06Um13IXU0kpxMMVEwoKuy
wxdNs3rbmFWEnr/kQTO1AQbSCK2uVHd5pPhCj218CxHoJwHEBhjSkNU4GT4zwWXA
btomsTKu/jIPhtacgan1fm8E569c7ts2NZ/AquKc3qDjq7ntrm/swwAIvkVX6G0F
NLQ7CD9ItQLvixsBdtbHz2AMvTgybVTR6Vhyfn/IVQLca5YlhKLOH0WwzXh/LCFQ
sRiXsTjMIHLXOnxvnOgX/pG5HBzk/jGbHCwNeGJO3CtOtxZmb+rj4hTm1ZsaPZuo
ou/OhqbgX61oon3b8nZ1qWw2aQ965GzedI3FEwliFgOX27cGNMM16/t4PLWbMO/k
y9oKhEJtMS87fFy2lDAOgE2ILld2AdCwNcocd7+pmQ69zHOF6oEPqxMj7qb0tpkY
I23a+IX7TQ89ZBfvjR+courrJE1WnrKWQX5iPSlYHG+LYto9Qx75v7KzPvuUaQIh
mqybIlKQr3jtj2Tmx/P2q3aGWPNVkElovfUij0QfNuioPKQI08Vxqhr4OGWegrVe
M0J5WgYw1iXsZn7ZYGCESi8manRQG4eCAEe2PONYqg9ps6lDFtln047PhbK9DDEP
MwnEybje15CbTocM9qH9aiwVgnGv59Wq/V2QUTkCWd1d+XQSStMFIeGM4QvxJlUh
6sqR+XIRZH5i1s7uVSn/FtOBxBP2fJavh5VyMCUG2ZdDNUBODVrAz+bXbSpaUk9O
i2BVrwjckmOP2ruUE/rjKqYBiHool8Q94HPs7ao/i94+tExRmhNefHYK5QguHPFf
pnNRMbGMKOI7DE5m85040u4YEW3v97BkEN0R42h7qSplygFEtKZoYWKdCsEaxDXY
smk3WcjuQup/Imfn7e2z/AUVLIbUMNXc6yMDFe9JLHoXNHl3ITqKD3Y+TrakR7UJ
/9wmzyrwietZ4xsJ8sQbAnl/8J2SIYjyPQEQaIPmZWtBfyLGXNhA+sWYDx4jG54S
CTccyD79STl0biyWSlzMgk2ESvVUhlt7P6/vQQLCo5HookFDwgPr6jGCOIVM4d9F
IgEzGY3odfj2VX0Hpwk1zU9lYaw5sqYPX6tBN49x91JxyuPnp+Pjw7wzoJQoGGjn
VGv3VMmcnni3GYEb6pPW6ktHzTHlnCYjPJ43i8pYP4ERSKPxmGaFHY71icW5npC/
PRA4czWLTHOJRLjiFsOhquy6ESx9Xg6P96t/yIKVC7XFof9FC64qbz7o12sMZK6w
T9JywCK+y3UcexPJLX/HCqBonH/AXcTIsMlX/6TUHpErqFG6u1RVzTY9eo4Rzyfq
ifzoPAJYPK+LUM8kC8vBQvQSxtMDc5nNY/JuyZFHamT47tqi0SIHC8dW12pgchmq
1u71kSPny5K0wu8O++V2HZg2xS/YHecV4KkCHzTcol3Y/+pVTBbWEt4wXA5Ayqnu
46gk1eHzOMKIcRDSOSeJA92FR5tPe/30Qtsj8gXiZW2eG/b05oO/gyejTIQkAHB+
nSPF8SIvUqNoPawWM5Q73DFuidPO2Z9ekBZJEmdl6IYhaaXJ/r18UTEuNGNs3yKp
amcXD6r7agVmdKHipcqP4QwG+OQ30Igz2gECyVcMgfZqyQ5bow8fuAJlm6v2nGVQ
Rnov7D/CRk5nligxFc47z+eiMvuwjeeYM1x58F09rnovWzcxVr8Spj1fkfrNDSj7
/GO+yMOSUd9MBU8QB9vsCyjUQ/iP98vuT4gNszTrtgtD8NNhsAq+kP+mGFhRlRu0
vQk8Q8DzM0L+XGkJHIVVTBSWdD+SgIze0FDQQaj6HS3gRP1FgF9sKYzHlXMsyIDM
MJ89s+XeJVEg4DhNlus0Rrl2XrGjda4CUy5JOQ2sJ1siX5noxri1KWNcpVdYfL+6
9Qjqkc3aodGoCTH12dPRsqavjPGW2Tz+wNhW92tEMVX4mavIkuzxDIEHLm2I3mLg
COJBRPJ9Q2MGabB/8e9FTpNyhDeTTvbB9br+q6WmR+O/JU7hQ2ao34xzj6g6OJW5
Ex1O2bWxHa3wDjxMFz6fUZ/RkdpCztmNvXnwGb6OhBQJsZDG56/gtxurXZcmy8h/
ippVrhcd2q6Lc63/TB60HeQMNfXdZ5Q/GQhyy44/4D8yS/TepdNPfGCiQ4IRz4YU
DwpbFyte00iAk5A13CsGVwwkwcgb4gf4D+3eKQsHYPPNP8cvFMQH8ezia2cWWFGc
yy6+JXrV2dom0BWTPWx0wet/ubAV5D3cri64BHDJoStbTTQZf37KLTrhP9VXMkIz
TEGN55tq9/BxYUr92Fq8U6tavMZXmm4PUdXQj+5+rbH9b/INrQlsEvlkZlstiqXB
/lcgWVpXChM/aeZp5a/U5UAgTkApG9XR9PTp79X7yQUk6t7aS/GBN6Eem7LXUZO9
8Z75bijTmItYXdjaJSOYfG0VuiozU/0Yciedix0VIQ3K6DImoZTudYEJZgGiwyUB
G/yiaqqwhcRxxd8G965Pngpva/KD09SNfSrnskbwbQqBaWdZC3onmcFBv7FAM5Xa
vx15rbPtC8RPW1mWLsa12c2d8VDpEVIhRhjypgnIWiwoyegO8j3sc0usGrFiyuzb
ZSNkWIidCbFaTRqNE367yoqEvfzW59A/TvyxvnBQkaFIykLCmH/PKU1QWHZowTtV
Aw919/DY9vL0dp5eownm5iMxJQgEgL0nmwrpRG7tjinIrTdyOuSuVh2bOLrdJbwZ
w9AmeI9+/ip0JTgvrNEVuAcW0skvDZpC9hc55dxq2AHL9v8CHFm0OrFlz+tPqExh
Mc83ZzM57pyHHES8n8exDHaVd8Fnuh6QacJ5wBKvcgwO8t0pydeuDBDgcpA30fDE
19/7sanNfhMW0ufd29EHS682n5pr4mYHfUunAapFc8O4F5M+AsWX5TmiBUYTg6Zp
1Ar63DFC3ybYyisSLTG/+FG08ygUVqc7B8tK2oHhNaJ26WOmsCq5WBcT96dv/YYF
7CxD+UQvVa9kvSRxpqiMNg8V0ZY6c4mXdBY9RThtWFjAEaQcWGwZZ6d4JJEUQ9Rz
6KzpT2gS4PYs6bC3hvObqjKgPZbzL/REcrU53KzseZgUfVUdIrvktPpRwATFqJV+
pl+d5F3Ou+i4TT/t/1xFa5NeHy3Dq+ZYE9zTNJt/gC9+F8pxrqm0nEOg3yXQ+BLT
/3DTywoRh3xi4KCAv970cUQnR60ix/1zQlUHtGXA/Mue0GMhstQw5/yb4VR6NG5y
AhUZ4CnXSuM9Usxsix6Q3xHhynd/HTFqE2uR//XEBp7p0RIP2nztJqmyBnzl5dJq
+f6R7x+6w3KHVLjjQZt75jZpe5SoAMwb8FaVwqrLRyi0vx6A3ibzAcWctfcpbx17
thRXVGYSqZsamPxOKh40OJUNROBoHTDJwP8qzkGChjk2f6iYe+H4vW7oB/9zjgdN
ucHDoi53jGK7LyqwVZBBVNgZ4TQ6JTiqnQ3ES+LJPRvVmY6B2ZITH4qZ7bn9/i9h
9BP9XGXdLpwJ6s8KsvlSnvOoflsHPR6L7X4ReHkLzqz189tHhgbQMxUERLM4tSSq
8tnxbKTnS3H+eQ/ixJEzJmzSh+mVZz+jKNzgyr2umHz5+kFiT9++ngYXVV4p5kdI
4+ohCEwy0zuz/zN3UVvbchSCiMYe8uqpLk/NDH68MiJK/H5uNCcWs97oVqcqrWrg
mmFuKZNyDVRuEEmNQA0ScnfhE5MDh7eDdhUIlBzYfsZD/dDwU1D3NZx4lUhypyQf
4j5W3SupYqHulX2hBrXnEVPRp44CLlVMdpaa8RG573lSpn1S9Vmo+OpoteWhfJ2c
nWPNQ9W8Az3uA0lfjdDMqF5WBbH3pATKs58YOMqJZdrpHGRAHZoD3zTlSilhBWv8
skcmkKBuVTT2Z4EI7XGMt2I1S11vLr6hMWD7Cr5G30HN6qZiqWq0AAuTU/Tpqy3t
VP6QiBh8e4iImFyOHFtFp+IU8O/qZOyD+VBAkCrbmB101gR7LVnz0LaWQ4VT4Csh
tYMgYL3u2ean5hQB6cLm/iFzckXKue72Nre2IQT8YqbDuUbCElq7V1eLsINbHML4
6twS4X7q0OMbvCzUNcihhxabpafdByE7zVKXqmf5Kq8yTLfaFjBHxd45ZaXM4n5F
UhB+mKQmFyxRgm5nUXpE4+MCJBx6xN4oOY6bggce/jRDnKpENYUvBiFfbZDSZx+v
IzxFvQyO+CEyUjRbsJb19uS2Y0gO8b6tk07WvGDWmXIRScKzt5x6lLNZcZccf6qg
wD2R0tiq2xpSGslKYg2K3fAhOn/HdOMZyx/zXVSotd0zS2+Z+BM+XwxsSJ9FRDJt
GLoT2vmVuCsvN+17B1MF7rpbf9H2yX0AfjXksIT5rCGxdteqmnUQV7iJZuLnN+qO
gtoIrybljUxU5KsY/69/afWHjPtklRgE7e1QrTayLH7aWvhi1HbZi4avbkb9MF/2
70/KcgjY2lZPagMs1iprIHyF4jgPxj5nz56BKidEpUyaHiW8cupRljnNxPe8rqqJ
b5OGBA+E+jzLWEpp7GzcSCqtMxYo7jvYKyu7hd1a1vbpSPzjLTAyCsQmjjSmXYSv
AfsMkeQpyBHFcXte+TEDMT4xTHrQas2gWOW8/7ef2PQn5PMbozBQU7/hIkDf3TAF
P3J+P/gHc8Fdlmtux/X1F+3o4Lwr5J56u7/xdrbwDrsqa065C519BXIurqJI2jjX
+IoP0r7ZpJIEcJiY2Y9v1TAhoAhMnlLS/GUyQHP1ihg8RBdoXtyyt46K5pby5pS4
VSWT6N0jlz/Z4+OoXXFcs01FzS0VQpJCuneVznOWkcqqmCSZl2mMU+06nArZ7nc/
SXPJtvzoO/z2bGxiuKlAnVmlKlwQ/4Mh5QyF0dsmSVsJYHPUGQK0ZQhAVrPdVNwZ
cA3oCekhKwqAAkKGPnoVggRUn+S0E5nG3of2q3d/FL7IG0tLLpXV7Z/1U3RJnMeq
dKfvc7mT8dtPZssQ8QaHkNKiTMyHy+zvW/HFjazJXgLarlFS51eRK38rHb2VIh5H
Nov1LUZQT7TSkEkGOytvpv0ZA6vybN6v+WO6cHEE5/f2nYRrhiFc+xxtmKUQ7zEt
IfsuoQqF0JyUTGVlWXYT1j1FQ/SZf6h03Kq6eE7H1JhVFvqpQ/afW50nrUoTysXI
QG6fGX7qp7La//wqVsM5lUyXNQELHl503pI7zGvIs3tJCSfnU1MwLN+f4Q8Aslfx
Q+sCikA9mOHGDKwfOZcLkb/qEFrG+Z5RxG9D58RhUvdVqonyZo0mfkAiiPyPslI1
hD6gKg0fC1BjVkgvLdk/1+T/rzWp5M/fDckEyoUflba9BDHKowDK0WesAni3y1LR
rkZ65S4VvXrKCAxZ2QMOw8P5bUyv/o2jXt9ycCFgZF7fU+/t7jzL0HNIzCdrZpxK
q9lpclh6nSjfxRDBlnIPh2SFqLwQdSYAE5aTPFUX6rNoeZN1m0dJUy127D9/RmT/
Ttyqm+0zCsJfaArl8RkRqRkwvGqQO7ZDszPiPuzNN5F5+bC8g3xDaW7yqvVkE4LW
xIYaoDwKUxO64msXfdL32iNDOQKtaXCWFdlJBAEfqvkLFPLSpyuzHS/VJmhKLxKX
/CSjmxSc5Lbl1oUO9SPs++bGoPaO+7Zrt/VjiQN7LaVg9IIzyOCMR3kTL+D/7pGs
CMZtYWHzNskHBKKM4wcuBFcs336RLdDBK3oCz4Ff9pg5DxfyjXP/WBHBxBIEUa6v
U6V48fTjgUDZJWo5HB2HmqgF+jGyIOT3QudPUcg0xPyE0vDLWWSs3yjQBprid83z
WmWXWhVDnAvoRD6Q0LIfOXotYYDj7cxBTlFqiRORXaIYt/cytcqIy9j0glPqKXmk
qYuRG7ZKdOXS0P4G/wuYoNBgWtJv6JgfHVkrl8CCxr7TeJnsxzMz6MH4TpZdNb5f
8Ih4DTYYB01+fB8KERh6amZcrfELiixY7K/rJiXZ4MdEe7UYHOXEjhMW4a3r9H9T
VsIKcTA/I4L5GPB4DRsyW4p1U3qWw+1CmAyj9e+KJsYVYBHzfoPWWy9bQhGitWXj
z/tI4l3acz5qnkwz+wh6DkwMxIiZ2+YXlmrS77AFqPKWcqd741s+tdfX2BYiVd0K
f5C9PSVHqIVxuTqM/QjaLYdrgmSX4gimIUdIL0yTWeHVjsbTU1v2gczmuAi14h/O
ckqovAEnmVm3Lvz1W54u1nC+F/3t+iW8IjOw+e3sN/Rky78HqjpSyLdXgafaA17Z
Zf2xd/9iy9spYea3tQgfJ36LsjEH1wkX5b0sIo/jsrArWn9arSYyzSDzXKoZye71
yY2UtZka/qewIvel4jsSHi6SwMnw/loXyXKM5UTnmHh6XgET54fw04sr6hGm8jsR
gB0P+F2S1MWX1MN4VyYqtCT8u9B6V1dyg6U2kaI+1XyEU2D8TTZOiTjW8Dtcu+VS
lJmiVtxNPTIbuNmY00XvILEwTt2fAVq1FFa6B6qo/6yF0iV+8LTI6gqpAyAwUKiC
vBWXXje0VgHS5oGRCRZyaQlP71NjdbI2AEiaHRDd03wZh8L5XC7xy+gVdxAn6cVb
0B34ve8+yLny/ks6LJz+ijJNihWV5e/rCVR6DdWHmoyJXOTHd6+iMoZn7yDkX7SW
ujIU2el438Mbu7yaD4cwW5Cs/p2MG/dtLB4YQKmfE2djt+Sxy7Cf5e2R7hGIu+PV
uvjqMKXzushy6ac/l0lkxP3SRdi2xA/lGXHU/ia2epvWFfx3sl191gl/OOmLKu9d
oJ5kYiTbJVQZna3sJtF+on+EE2QWrweFokkzGRRdY/0LJ7XluUHpG/xbeOTu8MXk
wc6nPzMPVfvXJfOaX4A9BO2zIU9qw95hfLMJT4nwNwh8EUQK4uOOZNrz5GnMYAHL
92UldwKHbnTGQuQ4UUq3pQ+3BowdTRzDwZq0iBMqGsOzjD63gUSFXVpgvpK7JxLM
wLOzV5tEaOjOTTE8h9M55NVciKEnW+uzK+KfPcmnLLxsA+EC8VqHmdTvJyPKbRQh
bGV5Je4fBvpY5FkxXCdHI42ss+0xjZ178FQO1lw9EX2lrOExVTIAZG199C4em/oL
dPLEyYskINyn/6vFOGNu0p9sg0q1gdvCn6caK4oDFgtM21rsHPbR8yAb0SBYFiF8
tuMBe+uquwz7wRD42wQ7r36DNQj7JLdgdrt3Z1Xh91TgDiGzGKLDhSZ6nC60lRl1
ubeaXWJT5/NyXp1I9uXo4QhFdc13rLe10qzpggkur10Ek1zmTEr+kz9jjLUxBccG
zwrOwR/TWcT6tgnHrVrEYf/65mDp49jAaFcAS/WcJvMd+HjL2IduArwejyFaxaMv
dRqT49MxB4uhDiUvb1bGVM7RekLBU88r0490IO0FVtR+ZofTA84xVeWbkAnheuGp
B+LVwv7b3SgU5dKtVaivLm89FB1k7TkXBMe5t0n/8fq+z2rvw06j3G6/z98Cg/sC
CA1VDT9M3PBe/VwQz+u0jYrt8kIBTYWpe/VceHb4mkgxquAvQcfhHqy9vlxG63xB
4Tgk4tx7ZwzaQyW7LfnUFMpAgWrXfpppkYrhD9bHSYeVGUiuQbF3v+BvYMolUGT4
1uZnXPTCUDBW+1y7Z5OP23h0HOyiJwxQOtGfffzkHKSR9y3VO77FOjLnDYFgQIhb
gJUvGrMUo6vinehoJ+x2V7M9rYdENi4eEvXmBT3cIJqHiCy/2+1qi9MZ3y3IhQRu
MVsh62Ws8CJL839JopzmkR3eurS13uE4ax3PD2Dglg8fY74jAOWUPnipnxxxSnSK
TSG0B8o5rf05kSSs8c08M/mlnXu9r3qL/l20XeZLZk5w8eymj/unz0B9Od2fd6IN
oONxifcS+mLe5wWw1kLwNZLd/ENaNGMokdLf3q/Al37eq0SI3yViiBjyM8s9j8Z9
UoK3S1JmlKAOE3Yy945jZIJTE10jXGNJ8wnt0sOcVYCzhA0PZPUyTVA6zsR4geG7
TVC1IdU6ate2LqBlpFq8+iMfiQb9hzzFfh2NuTrhrh8/KfBRx15+vVY1KaGJ8Noo
lKU8qKE9pGodiLhGDFqUJOX4rFvrOyj5D1YdSaSp3mQqDbrZq2v/XGtxwyC7f0jd
DbST6yxD0wenrp9v7vEVEhTAK9jFbTS/gPHxbpKenBQdk1eo46JqxZqUgr7yc9RJ
G99rh26DHEU+FFh2CQ6FUy/omOwltQAbyb9U3IUhCWxl6sHEPCQ08EKsy5i8stm1
P4ErnDlVSQhUUpX6Ajjb8UIxlPIjjKmIIteLhDRgdim6Rwq+HcYLkqoXgz3MBN4K
wmymJL7wkqdr82vrf8IZqTHyirasvn3P/iDznRk3vZhAPMhdnOjXqTCSNa/2ACHb
p2NsOKIfzZbXt5WnCHm8tFaGHfu1l2SsW3JcxMDSX3cEL09vSDS9Wf4G+TLxejB6
G9UiTzF9584ropGWdJ0tOqk3eR5k1YHMsSvvWrvd2CkFloPH+54F0FupaEfc8kmg
QXs2pWaQgN6HdCvnasKRpWFec6pJ5WXwa2D5rbFxELY+xbKgtebMShR8L5+UnNK2
Zu5i3ft/uN/NCzqy4o3IlWecCn7YgEijTot3oPV40VU9VOQ2cz/LdTJ8DR+2TDIG
FS2mqemuyx4O08KJgUMAXoU6a2Yg6cDR4LdXZmgAHw3rVuVxpIb/2Yv9BhNvjyBh
IuPgxLA2naSjYd3YGXGrgDL/RO+JOtr7+0BFz7CgUC9I/hhCKa/BEYRnwI56gllX
n7K/44zcBdyP1WCfpCfnBBONwqqy1IguBnDVUGBaPcs/NwaSyW5owoyURiejAwkY
PsnF7tPjKIMzihQeV3LQR/3kgGKBnju7k8ZUlrKNeOWaxmCsjeRFRSQLA1xpQEGL
lh3BM0j3Gb5zMD4JApvGsSXdkN75N7zMqdxFtcPm3eyJNFiJQlndAYqM5L4WVlf2
yV6fAEeHHuSuMfz/g2Amq747y3DdLbUeLS6vflBLjfNVNPJCkSwJOhqp8s/6RPEo
osNAoxMd8D/5gwx2Lz0Vu4ATSXN7o5HupbVkyA2iSMdKGGTlzAdH1rFLHEwvk4lR
LaarEMzbmsdDJSc/KRPcj2z3bAhsLD5Q+TWp2gcSzz9daiAU3nJ5Co/WJ8HNKEuS
0nW4fPw1TfRow5pDyzRk73Qc9fjOt0yvgmKG1vYEc9mDQLFTWat/muD6jimHCrZq
Le/9ZTQmVO+qFt/VJvpU9HWmaRmIK/YRpBSTWXAA0V+x3G8x8mfj/DbVcGKoag9x
mnRueugD6MNQJiRmnkypvaRMnpBT9N2IDRkzYTb2O+nHUlM8Nyy2JgUsFaJclewS
jriGDHsDsgf0Awz0wazEtk9LgafukpsN+jKSnGfUwZpUy/vmSReOVhNn3cJA6sfs
35OnZExFBWBItU2XNyhULBy7U9OWSOR8v79gk9+8GxcyXPmiArOhFYhl9d8wy1iG
EZ0+DWmUqF/J+nF2PaZeA+i6mmW7AUOptCINVHTX8wknYtcNBZEqdzTHCB2LuVve
bQDVnVS8MK5UDERQs7RK+VRtLPwKB7JojSDmmK1pmgBdiBQCwAfIM6fDdhj1Wo4T
IpEofbc+RuOI7ZFaCvxVV72JL8F88TIRmRqkKUakZ9DTsu++SyFa4sudz/GbJdTL
ciYlaGPWeB5gJcdsxHoJVpqKlu+ZISCERkD/sgMpYbPHuz4L69ZxvvVFC4013Fvv
fKbB59wdmvF4zqzNINQ3yA9S1jFbXdAqp9rO+SHd0gwpOP2rdyT0cTW2zySniPeY
TWizjRNa5H5y0GuokK69IGgeIR9xFvhNiWS4MBsJ5DDsdR+ehMec08FyVaBRz6al
I+ZbN/HE76kRjooTJ3Jsn2hI9vflOeK/xQfnbDW5paaUH5RhJ/rPoE0LaSk2EJhE
/6mtCBgKvONX6OuE6XfYrI7aYesy8L1bnRh9SOJR4rR1Wl8+WMSm0VcNlW6I5vkQ
VX17zRT6DaGdJ1/X3EMPjaVu9jCCY/ebdYUvVDZEMKuwQIH3bYHdHwbkn95Ch+Wb
TLpgXK3/ADDu3MHv+gRt0zwJcJAHLw0u6sX0p6eYFNXgbQmdIwxgpZdu8ajLYlpj
3Ho2rToD9yjcB1ecafC9Me+B5sizA2xsaXbcIVFN3P5a/E4hlKzNt6v2FJ/1B2vt
MMaFj/iaBf16cslMjvVYCihMOwfZzKi2vQYFk65yka4WmkKEaH9EauzdTho8ewmU
Emav9yaXuJoL57D4hxQFueknLwAAq4wY9amJYRs7al6V7y8feGRo2vcSPwo+Buss
M0WbN70V1KdUl0XfcE7PyacZCYwn16O2rz806xT0Ql4BFqjtb+SFpxz/hLy9xLcs
TVac6/XeSzqLf+jZKnJBOjJ4KB6knudwunDa4TJFfD7RhSkKJpSS/1AVA3tcagmo
H6a1p01WqCY2S3HJ/pJVXRu2dIS5Iby4ZddfEgV8nxtKg+GklDKKBdIPHKBs1+zd
rcXtUryY75GFK4Ral1eSdGjl4IIovJf1WuxwLJbNxxRLJHo/Mw4au5JzGXp6dxKM
cmWZKLnVw/7qDWG7A0Cr/wAtJte8OObtSH3dUK5SDbg1C2KjA+ihAYbEtKYIvXpC
LTI+7ox9mBHnYtH//pYx0ShAXiTbDwHFTlJj2myiMJPhkERB8oc+LAPbJwg35dzS
DdwhmK9T2F1qm6I2u3feLCjON0I3Y2Pftzum5tgU15uOTPuP3FKZMCHCvF6uJAwa
yT0c4x5EtS/6JXl3UXqWYzoc84dz5Ag+zcbsGM/NRWT/q3eMH5DMRQpoT1SIyC49
n433nksoTamH+Hyxq9USVsV/fGbftlJXy+F/5qj796bE1l0hZe0rH4l5AM+BQ+x2
e4hEMPoQRVeQuUmxLy+sfzgfDA2XVkBpzFfZfuzxHY+DlzUBYuMA3oKdZeqqo9BJ
66L+YEvrr6okiieW9eUqhA5+enoIcB0LVEFz96AAWI2yI7iyb1Hoa+AMamip6Kh+
r5OYfhUKKZphqAREplNsOrHxv9vPAJYFH/gfSNTNtPRMQ5o05F5zZPEU325CCKU8
c/DFA9ksy+o7LDTGPZxXrSdNl33+OXnLOA2lMM3PXdij543TRS7DyuNXKp/lImUQ
1S8xVE4MgCL1UMVK+wk2l/EPlHdRv4i/X6KGDgv92faBJy/pwtww4m13+Gj3sXur
U0Zz7NRtT0l13Zy9iERzumwlPvzHnNcE/uw4bIl8sCXR8kYnb9Sv49/m+SppyljN
GK7IsaMSBa/ugUqo1KCCh3/GZOxSLwhTVKDvz2W+PvD80m4HREHWVSvn/359IhGI
wOPQGGFqBIO6MnQiN66ao5RCIgYnCN/ANC1aOfSm7OLty5RU3pdv6tBOu7oQ839K
JYfqdH6FnprjUZT6BomwGqK6fwlkHkI6434f7/WxRcydkoXeA1lrkZNORKfD6crR
3RmgppbjZJ2NOHuDh62nFeWrapDL1SuKENl8mavgBH9LLCbY598L7qIKXED2908s
yCkpCSF8jgMun6V/CTcIKWiVE7ks3TPokFCgx4nsioG+7DnuX/bZmzwvF2HCk9tL
ZD7fhTy8xrv+re/NqvGibcjsjDDkgynwlVzIZ3sKNnYvTnobUkeVTAOnAh3yfSjN
9KrI28f1W7cWDp+ydQPcaxNfQfAu2gWVkpQ2pHgSwV1zT/03fTvfsBOaTj+nbmtG
06IJ6wpYUSusZ72JMdI6GsvhX4ZbcfszRV2kbf4eWRhpFKon5ZV/UHm6T8P5hh5V
mXCwqF1zGkrCJ8SQwAr1EqmCgU0BZ4Z8Ml+kj7OkcEcq9mrAULzEw/m5Xa5ZExz5
zO2HMB2DQNECshG7qduL7+8uXbItz5aiv5OfqTkLlRluKygYwjC00Yeu70YGxH3q
JyNcG2fZgHTGvD7GNkWapQ6toMq2zJsvuX3/378GYn3kOYaIJyGevGAYKpPfERKy
yTqcvDd5PQvVvJufN3OvoAnSFMx+vEES0j4+AuXMrHTfSjRUpM6ffT3WDVuYdhjA
6e87nZHTs+fuuc9D0tRKX5nYxz8jwvJC89oqw+qz2G5H0sjnZmAQxbKyBJf+WM+D
HkLPmu2N9qlBpLM9Jc3YJSIt9eV5JPfUW13EpeqAHPVj6TfttY9BHGPtLXTlJ7L+
Y3Xo1Clt38Owcm2MiCgeUMD5mO9CIjjuzktCnohWovsmHhk4fhMh7KUfHpc+aJXm
00WRDRyBhINMPtqrTfre7Cm2tEvniwhT1tR8Ua8cNHsnnTn+wgL0rNQCbwJYOjPK
GZatZYkEQs80Nh1nvDpPWyUVsdNN2ulyeIj/pRgoGDFZCb4ysdvZJMldQM5bstSw
qZz3yrTX9xWFd0ZjeZcpv3LyRgHgeJjTHAHJo8lS4y5VUkrpmRZ435cNtsxoBBAl
pRSwLQ9eqdvCow6Uv4Dax8eomsfG5egwPCl6ov6TDV3EXY8EQ2Ou6V5vA7TzfToY
mqiXAK1WBtYgBdx9w6CSYVM53G7fINDapCiuTuDNPW65xDey2KrwJ/CEcP5iFapS
onhcU5DuLWlNJ0jlII4MoDQB34JRJCZh1byWqaUKQiEYGbcfgOB1QO1CoDOJCR72
Lo9t2geWm2hnSCeSiXP92tDtjYPNZHwdLTMHaba5VJBe1aqmMI6ofJFu2CJSN3t4
Uo9cKtnwvg2ONdiMK5di6phU8RNPA7JG7ADoAWjNcTW4K/GEoF0TMkZFzKdrSRuW
vjqKv5lHqMoqdYQSiX2jRNqP9mYKS+ZROLgSUrVU4MseRG/ITS1qDPp+N80maeqS
r5rvHFM2QWUQPjxLrLbxf+WcKrCIo0meDjQp2f/qQyQTb3t3Zy0llDRhHylBXzxW
Mg5/h0rVbcK1l1DmGGBPeAD/Eo3j6CEU0gMcaNK3h/PA4YjJas2W0IBOEmId6FvX
2CbrnSGlmDu7NMnsAsHcRYq9Dip7jrIuYr48xNK17+qFG/r6mp5Li5ZLKTVaL8gR
KYb9idJ2dUV+2+IQesoCUHabB2/arOpy/yYgvtetUficFgJF7pmRq/cejV0DIlQX
Pcu13/X99r7bEMsGkT7PTKJ0a5K8EuIB6E0v7mQtnt4rIB5fNSRakDkAQpxEBvm4
1OyxxWoKU7OpMaEWUgQYQGZB4m1iy66KPlyDbBxfQ3tQZpO5KCD7PTW188jOnM0A
BEJTk2qwGA6P5YmgBikE+eGXNv+DzkQsPuANVtVXeXUkwsQZX3ojG4jirI3ww7EB
gsi74MvTm4hsxzF+1+bFzRKsgTJxsCQA75uY3706829sd2TNDqFwcoZzMEKOfQFM
JhBYdT+/0ujMH4XYV5TAK4uU3/h3x2BmDXlKsBCF/vuqJAmLormugP8qcLbbJERp
cYJQEwLcI65UizFkd5BsEbSJ14y9XJjUUHGfsvdZfV1TNkF0t670qm2P/1HpT9rX
xeoeSRR3PiIaZq4xzGfk9v9vkL2aWiK2F4wOCl0sYDJbdDhEgORuC8gqtj1CBvz5
/aDffu/oVH1t7dRXtnvi0tUPoKXIu4U4Gby0wFnQhjZV+wV9gZe7InE9iBbv6yqB
eIJgHXKyCWuwv3He1W5c566ht29UoKiCGOzx0Y4EgvYKFSl/bDoQGWDsCsn+zE4n
inTQ3PmDu6k9arS1BBKkG9ZhoY7m4dj5vXRLJTPyHNkC7S00i0+ijuvZYMlF3Zj4
suDWEOZ+k6GLOTixTWENujqQSIJsnn/3tTK0IFAZis9Ri6PY5zKKgqHpqClZcf9R
0MNcMApqx7utnScJtSqYAl1h//G+Ysm4R6boB/1r1hl6TEl91zsVHHTygW5q/F+0
qx1EwJdciBpmRl3cYTNdzRvNvkrDi7bDjIHWVY4MTScufecfb5VrzGRuI5m2pFO5
S/OUgUpmqRFsj0oqVGBP41PASX6USS35UQgPsc38vx5M2m0Bt+q10VlSENE7rlHg
u/XTIY4V42rVvEEvI29oFhvZIbjaHW41niHn+to96wdSysSJhzyH7/2Nwblm7vZV
a7Y8RRdtDdVqxy69leVCNRuAcwqbAl688asf5Cr5zpasROSckZ96hItBO8KCb+nk
hgtud2hryM1sbXapONL/fuF2x2pKYkVBnfd7toqOztMpPpuex01LkWxhH59eTS27
NGmo/8Y6+o1LBdnbMj3JKV9Z76JA5lPpUa2HXYnA7ap1qz8chqFEy8tky2WorU6E
lLmcD52FlEXg1823Ka9vVxACm3bgjqYyQP090bKgrbUznJRSdjgj6orG/wNSM28P
LsGPhDCdscwt6KILMC+Su1EQUL4MSYzq/9j76f/+HBmRfICKaxMhJMjaU/emMILV
8uPu3LEtziF1KZQgWx5ib1iv5q4w1d4vjbrwAiqoeqUCuZTYsfZC36z5bKOXAJoJ
iWQTqUgYgzSVgzOxC/vIA79nKG2s3t/KQtjdybIGnk0DMAPTKipId8PFPEqMCMGM
Uqxz9QafZV2pw0RhmrVQBXKSDAVLL5aXKpfoa+eucQ3Ph0QsxXw3oE8Ye59FM7oK
sJvFznFVIPtZywt7w+5z9qZf6rwNMLOzsMb3qShb8f4HNJ5NizVec8BT3MDcVqb3
ogbqKQDEQwfiFB78jciAuG9wTm7wZgrXUiZozUTYk7woBHYM25VlraqglB4tRQPz
t/h2rqtxkbx4eZGR9ikASoiEksDhmg05qN2R4KIeKDJkDx1tvqKPn5fqhKL5Rgem
iJSfuweEbyRyJ5eiEd83Ia6aA9y8ltldY4YWkJcJPZp+jx52C+IV4F91KLQHG83R
C1PjZaYW83s3HCizkXu1T8PPv8objTiD6bTE/tsoJFvnfZtXsal+7fUgbl1uYqfL
QiDLuJ5fX2f5Y/lGHzzYE2Nl1CRkhKC4SYiXO4LO1xwVlMgiBtRcniMoB+KkVLEM
92jybXCOi1Z5yxGSavWRDyjE1VoDMPn+dK8y/v65gUehZrqiC55nJdBjXBEzAaBj
ri8Tn1oKJAvgW6SvdlKsMORpR171jQyLVCJCBjC8rNS8kSHz8AadJvWnUcuJvQ4x
kfuH9OjqLNCF/PT9Q13novrMOEie8aCvn6uXPH/oqc2rBihk4828CsAccCTBpU8v
5Vet9g6DbHyV5mXiURiXeL+75j1BUFanoctWFoOYrIH9y4SoYksaYDMExz8kIk5v
y6PsEO4F2WBVv2ZldONl7P96QaT9ODla0ZrbOMK6GqoVad+AorqXpReDZg4gnLKp
QKvHRwUfuOBzre1X8eKSywnn/rduHMOHRvr/XHlGLmHHUFYDggJRR0W/YMGpYqtp
6U7euVSwJWklA4r2mPAEooSTWfExZ1fg8PPTNYkaTX6Tph4Bd5ScDQujfaTMIba+
n+4lGRmkX9EkKM2ZqQbSQ41V0ywH0Byy+IK+dzr9p1kFsDqJR9V5z+MX+RRBipik
jGRDqadznE5hdtDDaUNMupHFw0B8Kjf5z45+KspVYCmIP9Gliy+mm2csKmcxd/lS
bGkJvjjAV0l9aYQPExkN79NFM/85JI5NrLMookfqdA+E0biAwXYPSStunkeQy65v
LYXV6dDcGyZ7SyJUaktHhwGiGrjs2UT45oiCUQKXhIPoQvP5F5Jfw6NWHZDkiTH6
WhXc3LSQ8EKzXd7SdIEu6wL76zmPmawjm0wlFPOR0vNWbplwln63nfE1cWOO3W4l
T1og3bD9N1oBNcqN0bRnTjO2GjBYjdK7Hh8e2nFPgu7ito9RkKouhH1a4iKvLK88
t5+mO0pl4GYz30O9mb55mKsqRENZuaDpQ4sC9/ttoDJNwtcsQSmowA/FycfpzkMq
uj7wPQI7vARR5xYgzZkPsyDl1DSx32sKXYDK+h/PNhScJxnmZBz9xInIWW1qYw75
Ra9Xj1kupp7k6V0zFBlfT3y8fuDN7XeU7XcEw2d9f695QRZE05ZhpdCSwZD5q10m
+PRSdEjLfYeFrwClxUzY4bTjJ+ofP2+n7ZBKj1UdK4XHMTxDnPngABWVlgWBMVJk
tT/XFK1XHQ4NwN66K0xkMeIXkOHfheMGrXR9keDgWwgEquEt1nFCCMAC4SmdTc1C
jW1Sdd450JAL9nwJTfdd7Y7iSOP2L9j/pZxiGJO26nvc7021lKObPmd8evTGsb0o
t0vJQc8bc992kGyEBeusPtlwYFJcxEm6BptNhY2ldv8jsFzm/3ovmgp+AtM4Edhm
lxTIxTgWkQ9lJWVIGeA4TJR/l1ISHK5a+k1WCjEG5Wy9fGZJ33WIqmuBHOGTG7EF
qzb/DxgWLxoFXhsRThhk6uEP15w91c8Jouv4TEqbgbIxy6sGzu5vLa47V337FZYR
xlVmF/pHC+AVJYT2B/6XeD0OD90ltibjQoCa8Br+gHJj0oXIpej5FwFsOTm0fsMi
cZn+P8qxgiBBXEUhvgnUml/re2VvpiutuGzDT1C8W166Pdd0leRO5ejlml8FaD0q
BVWjjxqrYLSfRcg4PRr6ibB22Huk2wMDTHK5TnJNz33MVwDhIWQ8wv7Pk6xDjRCe
1oXwR9LbK4fkvVQ4ST0ynRInbEtkaMF2bUoTCkMQakdTJHjjbwHxjTLvpCTkVF9u
OiSPAZ9W8+RcW0KT5mXwzCyqSa9A2iNDt2vyd8mc8u6uT80flTNnUeNnPtndxzr7
RzpRK60G68ruU1u8XRGEOS+NY1/A2HjczE29ZN4Io7LWitmzciGOD1obOFz8+eUs
xhAUtx0cuv8lpr7arSDCDzFSQ49qitzugha6tDXr9upVZ04Ord9sjyz0epx4P7Xe
X6Em/7evUnUP+imCbzbaLbpXOHA3qFgX0FlCFxjqyyBFn9Rqrgp91f6y7nGeDdDw
Ej+QrrFjhQK8fpASjTGEn9cSRjpGEaV+u/A/JR2BECV3c8rrI9+9lj8JHn+t2ZOo
PeU2HJ/nCfJ1bAtGyCNzc9G+zI9elpcK5+6KDbDoLWDZ8JcqHr2tMG2GJAtZruYn
zwrRXv9orb/IEwIsMdUDJ51fkAzeDXEBy6nWubguGlk151z6rPYWRdWxDGGkVBz4
nXeJmfGLM1PMu5AdHHMAAVcflXCQJCm/kpkXhdlKwb6/mIet/IY8lQQosRJp3SU6
1FUFQaBjAkL7Vh+k/aXiJvrkaWfxt2ULkq56rdr3CDY8YW16rWRy2qmnWz2UJpAI
tOldYP/lVdC1KzisMx+d8t+kOwZPMBc36cKiiR8TOopKMsZ3ktsrg85vGpw8d5N7
iRMd/4XYGflBHRfAbGBRlruFf5kaj1OCCtIFns8E7KJ/Q8QhX1Ek3yynMTfkKJTQ
rh4LJzEpALLfJGYxpTy4zmfLiSnXIJeo88mgphvvxTvgMs1Axl3W35C/fXV9YRWg
Wrl7+DobH46an/I/WSVH9++6I2mKi859CtxM4w3+z96/st1Z0Jtyf5l5O4rJWA7j
l6bod/rpZYI6paBqY2oO3EQp9mv9K1RFDFnushEtJVUVGaKcRp60SyDqAm2ciOY2
2UNDLWLc2GXsFu7gNnYDoRPZetqH0I2fohQtYRIoOboKmK6CPpsQenGIgNW5Sth4
fD7+L2ffkxce4PzouotzAs5vGV/3chCnF7UpuExPRwOZW/0EJ06C5OdC9kzU4+UN
E+nymKN2GylwAhCPdoKYMh30/E7Q2WwsvYBPz67APEhP5MkfKPHF/oPuQHGFdJfx
7fFBNsodDUAhgWdCtSrU+qSwWwJyt3T6E1Ml2DyGY7z/0n7dXd1EhDnteJJ6+hCX
sLqiIIxSsXYp+KYZZLqDXK89vKHmOEo6sD5QqxNw0uMlXCTJBLo5xr04+DZqGLuP
hAYnEPaBP4nN4cLkW8rl7CqXXulr5/j1ltn2Y+4hfGen64nsrtGXZ0hc+kWfzSGJ
X4VSD4rjK38pohUcbG3E57zO3+YTYPLMC7armAbgB3Z7nccGmiNGfUw1xyX9pV7b
1/PIV8YUh247d9vP2iLoWwEsX8Mh0mtVUfMJL4h3IprpwBQzs/dxa8zFheOIpjOJ
Rq0vOVLd3LeiRPQ50fQmtThaEPouB/VDYk08o4RIcq8CAAytBFoVEkCf9wNi25O5
j0L6FxiVllj97Dq05gTq4rdrHLsprkCfBCBWXalOOdyazgH8z9sR9wzItAjPBzRG
XCfm1ZUh7MXWXsAaMmNMwKO/7KRJyoexNyrViv8wAhwrZAXYiqMN+qYXvnJqDBxW
JMT2DzAyhCVBAVO6Fo+hAiJk6G9i4T62XeKGXb+tpceBxBKYyehV/l2TxptLJTP2
uRhJcni1V3OwSDH98FrsWQOWBAKbo+DaALaisEJsG8SQCa85oN8yEykx1lEZ+qf9
tIqO+9ymDK5ajA8wl8ZBq0YxAtDPI7ZNewyndbWhniPKMbb6I4LjUYqfYK186qqd
ujZIVpv4Zt4LMdgK4M7WqcMeBzASCbDNki6OGYvWSfgNrmWndil40GTjqQpgTpWo
lBwBDqwGkkhqcFBRGCfOStwEkLX5Y4IlYiPYBijdZX8bvEF+J/3afE2GI2c2V/Om
n+rhLyr+gfxTs/P/lPtah/XlFCBHICE9McaJn9GoNqsdSJFyEDWvY2F/88cl5eKH
6CgGV4CIqs+dGk7ym5UK/vgkSmIlwfh30urR2tMG2v6UbiKRAuekYTkuIrdI4p+l
8cL1qlJ5QupskC2luVY10yxwJBO8HT4cLCdHTbUCw7A/6EihXn4XVDi4HlXR5Xu3
kluFYqDMqZPHCncy7xc0vLqnuFUOCjbUstY1Lz1Zn0jGURN9nNkApFnsJBwcgcBp
1iJyYmIPFIQmyrwUWf7Iirhl3e8mjKnLoZoGqgGLAXeFzPpNG6MWKV5J8kw1s6PO
JPG7QKF61qaxJiq2Ctp6hYaoFNN8oaLy6TtH5L5ybqYlw+ePZQ7GeF+snWm2+Fxk
an/KCrRaMX3h0OzOzuaRn9931HVCYTqq7MP9EVZHksdtkl6E8WoYr27crKHuHmor
BlNeAOAxQ9xeZscN2GIjcNdNyMElIxiVTi5TUFj4ypN9Qc5+7t5Ui4nvc90HlqD/
ZCE5QzyY6JBcsv8U0xAkreIUcR5NY1I0k9ZzgmivwFdb18cvR+oS4xzjtQ1bXb/F
su6OCyQTRKeOU1yF2I4J5DvbdfJflPXTtetMaZx7x0NkLFqsWffFCoBAZO2nb1Nw
1I7Ykf+KkJfYWBsq9RgJXNpGceGAM7QzrJ0F+TyC0J0NWNMDjQqvbXQaergKl+aN
lTp9XAsBjM5zf00e8oZ8aM+S10srDD2d6WJBAVOlklaTqX/m2hh8cPbKUhpkQ1+j
EfaWQFaG17TKAxFtkR2egz1tutN1h9vTepnLig7GCakDKE69FvZQbFBt0IK0eIP5
lP6Sg/73/r7fsHNSIlWVQT/VcosnuVo6DPBrJCr30XDopa3Oex9Ln3oWJchp88LS
Qa6Y/V5xpeB4FD5BUtnuFZCMk3/52eFBJtlqn13c5UmB42pjxnnVKLM66CpCpMSe
zpXyw89GC40wmyXX8rq2IdBg/IiC6X/chQNseAwelp1b1u/omjYYZgOGhJNuhnpV
ayZQg9Fve1I5XS5+H9GMa41DzxfobQCOGbh0UiBDPCzaf4k6e9Rk4IZwMgGtm9vM
l1yKrZVBIMduk3UTgO0GPXbGHSmdN4V3LYnPsL9jkjgvYuh7Wc9Lf/p3v5QMUG1f
Jt0ceEkeXGvv+GuwHud3w3GKoZdFW0/oWnsWHLjmje3sEqRaKnkVQZJlhOOYXXmc
yccbJYt02quPau1FO94/f2Kr/+5ciruKYO9+xHZFR7ZiPtrDYpiOY+s4yjvllr23
GJ/DEHxHUGPy1iUFE1EmRFYbeijXK/Zx2lGSLXgE0F214Z7H8wSMFmVBZV8kPu9k
MhNxNpBkqzjtGzTpQJO8ivCr8qONAX239vGn55RQi0m/aCKNQsEma6hpqCzcLRjA
TcCzg1wmcyUM6IR/QSn8WQEsKIFob0Vsx50jMnhOYoRjmGEtkOOirq94QScX8tMY
wd/3i5P6x2Fni9ENNhtWpLer0MzE0am5/K5SglujfUlcExxgZFEVSogLdUz+zsim
ZINIfFJMGm0agIPlVTXQKq4A//1rAxLQy6AC7F+oKBWAyp7xS0gD20YTsifIoFbt
eDnuyBUr0XQDLF74t/6Xap82NOMSvLPNHwZbyinerdFF+KqTLcqYMffDPM3BGk4D
QCxyfs1tyw+9oaHIEhehcr9qr5rZnIXzgtEBiEafwSZI1YFfV7JU8ZOcSsRqyO5U
m1H2fvRtwmJVRJuSsEN++VvPBkB8qYMx1VxWaN2wxI12EFU8YGRK3/TbeQjb8NGF
FDEc5uxbDkNA8IZasoHU4TZrrSi9fCfNvjPHDn33CKs1hIMAag+X2EV0iV0BYeJP
6Z+TUBtfAKhWm4pRM07QL9379pMTwKnHLhBRGE1vCl6JNz6ip0gwaQ9I99+CKNC0
DxI2GbMZSE8oHd43VvpO1gXW1Cvau47nwhVId9IP4RCnreTmwcywo9FMOAFxJn3Y
5oqjAn482wIZAxQv/IeCvr4YD0Mi/Lcd+oMHpFICKU6tNKWaPTnw0VaYBONZcisD
yC+DCVFLthkW3zBI9gVq2aMMfkTbXsrRymVFnqsL6BKMFwjgHmPfMhnnJPiz4R5s
1OmAx+DVAEJAeCSpj0d067SsXBAHVRo4xZG9XTR2IAeWeshPci5Yoj1yWtSq6Q3S
pHaar/nRGuNYYPR9DOLCBt3hok4miZZN2iSr0MzvfvuerLIHV5UmvW35CvN0lMXV
+skRHxmtjqdA31mMyuYnjuEgan/j2XsqAhiK/K1UhVqDpchJXSc8mczYvxAXnwLt
0ZP8mHBUejYARfOZQv5EMkXEBoszpKdmISbdb9lKXmpi7ctygtSAv5yZWGE9UBpW
SziyJc7PQXzwNDmFyDpukecXCHKh/w0Y/7AjevGcddl7kx6Sy/QMsyPisUC+LDRa
6w8j/FI1EfhGmNUT95KB93w0ezZG8RnANOYco3DeHPRtrxDgsyQcoSGfbNTV7o3N
bDG+FttL583ypU32h3/MSpHRgvVEuBAznHhLfiQvFI6Z7LbQNKcTxQ4mzHYP/nrO
Rn3U7cXUOfvUVQ76o/x4IgV3VFYP0eChmzvOAdu81gkqG748avZ253pJbNmCH4+4
p7B9CKlIImeeA1waqLkme5HhIwsGgGrUelo47Yk7rW2CMOGwCi+UIUjVjQ9S/GRR
X2Js4+rapbrjk1g7YW30x6f4YQCbJIX9rCYlurlTKiXQ/+3pvvExPj9/J4VWErOd
kiO/was599MTHAg+VboiYwfckCbmO1oLm8w+I+ZHhZjI0TY/+zSyy2iT4ydYW6Ts
ZTU3QR+dJu9TGZLIl6l23RsrO8t94YC2q9vgCKQrtD2que8nkAFfwijOQ3X4IfGF
RQeJowiPom1Ak2SCQ+jDWOICH5ugXsWMi3w/HsgyeXvMkm0ELcrKrMXBITB7mU1U
EgaGruHS4/KTNLhJ6azg56tC7FODome2LDXWhyQiddN3KmqRrvmqIjvPmFMEk0g3
eSycqgtOfis7caEXG2Fapo7oKrIq2ntNpTnviRTBt+JH9pOeYmnptwFviub6Cqf4
KezmeCLgAfAk7I8zXbi3PNDI0/F0jwtcd4jBDcXcKZx/9Xdq/iNFiIMzVBOHCh/D
R5tjIlyZRJNT6lG0E5Eb8yRuesURysI4Pjr70KTNAu2ihrTbyH6P5U+KChbnumuc
voTEqc3ajxlmDdCbCeIrJqSpQcnERyZ4Tr1Z7FgA3p8EG3kGBqv1UYDPY81+H46v
XzXcROGTkA+z7bv9XT0qn39HBxO1S+Tr60hfRiDIazABbKOt9wykyQmJfKiQavpy
qgEJ1pxVb6eLrbv/cAcsJuFr66+o0WcnNJjDYccOgPCaI//NSrchhyAJhR4sCnVw
FWSJdTN9g57S6kv/jV70qTT/1CeL4H/RHvY28FxnUrmO3FMV42xWzo2T41pA1g5Z
ZYPrtI4OlzaOEiWbkiEFLX1dd+W4fC+7MlQaGbJKgCes/wXYcC+JBhzBxruPHsDx
GgZYvoLm101s01ud2S8UEygrOAYWeaoPvn0N0KCNsQT+lsSeYndaE9v5D1SV1KVU
IfemGBlI3/Z7cVlABhHrIqWkO5E399zaQ4zT7rsxlPJoodkZBXMmdBKFRF2witvM
7LuybwSUIyPl0jdAmGwzqTQd3C1snC5ygQzyM9MrhdglNxEGU6rzAwDpVkJ2WU97
vRIqBVZqlU5ywtZXkbFwMermPzkEJ+sXYWTXQxkA+u1erR+04em8aG/C6X7ywByJ
HGezR53ljVrGRtHG6w7IKEnV74ndmTk4OABMplzegbkonNMOmW6uyaw1cVOtESbs
lxzIpXONUwe5PkJ3Wwe9Wy44IH/x8dJYCpiabWNI3Ad3M0WF8WiNIv63YLTYaLS8
0E2XQaZXDr4+Vo/5jgYTP85tm5ys+N78YDeZiSbnW4lM24Yhe2YsVKZpXjN9cZzp
gBdfDk9LeASjIQFy6dOnouptIcF721x8g1DIyKVUf2ptKcg03AK8JFr6JKo0gvOj
rCMoywB7nrCWw2FyBVTpdTcuPBhSrcOEX/dKPtDL5XhIp6KUdtnjsNS3cxlMvHSk
pp+XJH56zpLkF4mc2azqEv4ImkW94FhE/E/svJPnzD9hpyz3HZ6r+lGEBM41WXRo
9CAvHbc/TdwppV94EU+6Rfl3RFr3Vlpm+gmCv1IOcd4a39FuaUDAad0g+J1WIgJd
py8DdaVplFyGD1HNHRY3Mni7du9diHydrsnejlIVJLxJjcgD4pj/j1haFJivmmpO
lldCCfvTyulCP/eKYReHtmGMV4Udh+f5lIllxIlz9H5OHCA/s2qTrQe047nNw9TU
Q6/h2clyRpXKqSiDYc6awC9HkDNHlBZTnL9bblN+U1rvvDkqhwirOIktk9uYaLmd
hwYbCZuY1VpUzBAMAyEYrIasoMQW5JOsfFefgdKhTjkBjWhva5Os3lhV6M7GNlFz
DDAGKMQegS8GHOIyScLQXtO0dB2EcRrnpUOzluQFHD/pWNiTPTJTqYJH4/dp4S7F
A2XMC8ndaR9snsUx8kTrZn/RrJ+/mJ3ltM0TXU0CKyp9AKbI+2V8aegnMKSNB2Oy
39BCHC6NU0v1J8rUCovQZQozsWcmjbPtOFDcCM/p/S/ytZs9zaildJYuQnLf/++u
CKYvdiv5KFcop1P5eZIH7TRFgXa1I+2qxwJl9RLf502pVcqHyblqPusqaypVt7VK
0rB8JDl2/xDOZuOct9XX5+JvTjAzwSwJwN1DHaytRIkdk049Kj2wA5aQOfpNDbBC
SvWEGNHKj9vCUwlp29wDkDZLmVx0rk9GVI06L4jo29FSe6Tc+62BEfRgWA/N0kMx
dYGiZgqSPeoVMF9Bj0Kn3XALXACXXSQvc7rD22qflLzAwkxHn3OokfTipToH+WOR
Bkm6bxWZpMpQsY1tfxUoUZTC2NEdZ2xOIsyywZO63sJ9rzo54aX+KwtW6uLwiWzI
mapa3x2/qfCoCCSiryGy9Yp8MWo3b6xqsokDKhx1WrrFCGvJPGSNtTBBK5MApiBP
vvwyYrDcGLm/ucZNzm4VOp9jUBdLNR0K+RX15oybr2qzLD11x4URPUkokUe0LqVt
GySRXQHH06cDEgj7toQBXvxT25rwukcuYq8IXcTlrqkhWut7wAK0zLpJLywVfd8y
p/oO2JKvREDN6rJ9LVZkyNQUvGGtawnLCdTT2BC9/7ir0JGMfwFkaUD5BvdYThsR
YMMv+CH79/2GMUSySMSnVC9YJfcdOUvQviNlB8l3NL0Uq5k354UO9bzjnZ7bPWpE
jiMCKesOqcVYcD1KiEzEV5sf64e/t4yEY7mWEWGURXOgRMZe7ifhSG7cIt497e+E
tsPsn/ql/+wpWnXVNrhqbwRRhSWzWOZpa0sGWKQxnS9b8urJuJebW/HBRnnWT08m
P9dzinXxCtaz+INn+YrRri36AYDxl59pV2X0jwfmbBLeDBrFzLp4WcnU4L85XoDW
aLZrdMBy0h57iajXgCv/Pw13dvlse68nB/oT+/JwAQQK2wwffkBdRV8qoDqztRmI
lQJYQKxBJBSSP4cmLH3/SydXoBHg3z5RPcoVAebBrYSpM9OuKOKYAXfAURnJyKQf
b371ZniH+kxkG9PEaFF4nQFVirfuwwZhaHO57u+PLgta4QCfH5y3/u1sxyx9CHNE
KnzNKowvpSqYLBAuG51FRfX98uDeeTgBkDmeKjYMDgs3zMWSUlnX4PjtDj53LMeN
gEohhZcKRje3JcQZZuCHPFEWwnecDJ8q2aMp/aDbYUkjDjZYCsVQIad2JWhpLBxv
VCu9yHutx1pSU0H2ImvOLLVWdOEYKFtQ0eeVU4SrrRMrV17u+Tpja/85B4g7/ZIB
HUknb3ZHRhO+HSdNYE+F6XsoXqhQMRWjuMP1l7VpIRdzAqr+RHFuJLci6EIZ0Nh/
bAMj0uyD/mksiiK7XsyNClCbD9gyqC55UUbQ+nrFGg1CZ2nBkxwMe3O9/TNCAxND
enAFoHKxgSCQaKaeN1BjmqA3JCVRbSHXh99Xs/Xb/QEkeh2kjOIzBLoKLNrbSYTK
MzVEIm+CSKO+jsqS6dxagvGpA/GL3IwpuJgXnZer9mFVYc6hyAwCenoL2FI56RI5
NlsYG6izRCac8d8Fo3/fZPnNyuLhvDDanGq1mYouyj3olU/qyUAa92S7aBwTXjdx
NqsFd3Gpn+inW2ANO6MGAZJgu9RZGFnn5oNl7vsF7fpLgkoGizv6ePcky8/ivrMO
f3tnBpSHnLLmybtolNbpM9zBjCrVxpC83OiTICxbXL08NmL0zPDHAfa2ogqZ/6GF
PqTkPxqdTkt33zBIVT8QlDJJWDvdjiR5I8GZiFVeHpLtAEDAmN4EuFQhjUPsveDE
L/MZ1cY4SW0VnkrJ0oaMYrHyFZoNC6ja4BHqleqYcsYFDgLKnkOvElFQNVNVLtzk
7bUKqiWOsDboJq7fXySTWxthnBiIZlA1Tvks85CGP2BBb+0v8vxfesPOXlPwYV+Y
x2EYqnBXR57992Hxm4VP2WkD45Pz6QeGD2qE2n9uQahll5mijajV4N+MhGH1fJco
1ZmVZ0UuorqSSrDiRcAmNrgdoJh0/MMjkpvqdEJZDBiZEYh6Spt+/K06U1gv++PP
cl396NvYwUQ4Qqw3yjS9amsDN6t37WrrawcrwMRg7Z0MOM4uxfjhvQY18TlF+rtl
xxPuYGXXaS4rychdS15xMJNF1aU5b56D1lkmF99GZRBYjImL0PpQgvgsQKLeqfOg
gxyp8TBK3TxnUNdu25KP4Va2OcGqdtGNF+G7s5rqu5oYCxaH/DU1bFuBxO8E33Rw
B7lsrm+ARTk8golbOJPT8eizHLUXqVA4C4YK2IScDoNJ/JE8EPY3YJ+axw+kDQcw
yhMOufyFuECTZnYAksU7pXKvl7yEtdlP4Z0peeM5Wy3qryBhdMrE/KxYmC74Qkrj
`pragma protect end_protected
