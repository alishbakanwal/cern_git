// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:05:37 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ndM0Hs6uk94gWlBp3dfxqNdZyutXBuPUE+zOk3iZEhLnmBCwmy6pI+MQasaPtwNW
xk5AGy0ML+eNNS6cPzYTr5aw8KrbU4QfuTvZVw1oXgtohhhJRs4PuEQEc0lYvwTp
Hl0eIu24iMAhPSTGZuLzThJjFJCAmfs4dxr1tlTRSP0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6576)
4aKrcxHKD1k8BWTJk8dbIujtRD+CBjnzQPROkpCLRbCIiG6DvZ9lNKFA/HzCgwRG
gCyVg5ua2h0jKbJEfi/3085H8RmgsZEx3B0zPo+mKXaNioFqnr9xIP9E9i0nHGhR
B3IRFVVLnwRNivbmTU2WoE19joJHHHCx/usF6uhYmKlDYX6L0aF57dR7X2S8RkJd
HuHCI0SCLySlSnGyI77JNnpCfEi4z3kk7DVVYGrKsbziaveX8osaImrmvz12qxfU
hDC2p2ImsdI7jWcFLrzqDo7p+q63Xi7RWuxv9uHZHx/SzsA5KqBrYWv5D5NW36He
4QxWc8sT33EOMu6jnoq2o9J813OQ+CNu+L/0exSJpZCl6I+Kj7eFDxh2Y3P7JfL3
1crUthBzDCrfmC5P/FozVdSXU0UT0eZ3GaJ9iJQu8kx8X4PdGuwoY9nYFh6HDoti
MeKJabuZm5c0WlnTLevAdNwKyrJ87zkOn4AQ0F1r3E+ewvhKDlp0QVWrsmotZXb1
J6Tcdgju1urz/BDbN7LeSX6ouPsS+iSYEMdp1P1IDo5fsh3fVOExEzhD7+KTV9WQ
nE1l8u6BtS7etqVqm5sR5IZ30DoZmgr+qyd3eA8/c1w5yDIRMtMbOooNTrq9kpR/
FSSTkqHB96lERj+9klwswLJmqMo/AzW1ulSk7q+gmwM/YPL66o3R47PExHkecBst
icQT2oikMJhh0Apff1BcAzAD+MEz4GDir6oBGFuHLHszf2yuCMnqkLQoCAd6iQHo
lnyK53BXcjx+0LsvlUV2m1JCh68IpMP9WW4p7Qz+Ui+gKN/oY0jeUtqpHh4DGG1s
dAz7AznMWt/pP4rJ2jz/BttTIJzbi2LEGWNaVt5auwkFI6VQFAfOfjD6ZOQyo56S
p3lp0L/b3BKyen82B4GDIjZiOJ1cZnkHIph9pfHZFn70M0voWdhoO77/NPu8pJUk
ZDfwacMM8vuqCZyKJyVPQc3oPEVZ7CKBv81ED2ZcHZ0PaQDvov4XgyB6acUUGGLz
zwQJ/eRpwGHhjdwsv1kCbuFQbwZ/OcZUVdLc5q8SI4e0SMn0cabTBwF7gBNwpvZM
DKGEMWJlR28gl3lHMoFABgjaMB0GN6yT7UbUdRIsDae5cfrwqenRxvkjwIkcnQ8V
siPoiXd44wrigJa0uvyJGIbXbWb0Xoq7bcYqukiSaS8Zc5mkdddgZoDpdSVab7PW
9dbNxrGNjdF9leQo3SMlpKaR0h0VplItbiCbni7b9Fom6Jbmlzr27FyGWCfihfW6
lTjzlkm4EDzA2nf9C3qWjC/btcFvw4foFWXeAQ5FNarTUrrpgX2qj5YD7BEd6/Uu
bI98Ab3jD4lHrfVh+S4M7acJRYyBplHT3vdwk9WXIWARYw15y75MzUq/i2+wb2yB
jbvXenBm/YWlSvY3/qmxKibzElMKXekmTTbfoeTGvQ8tDab6mrGK4o96iAPJzLyK
CblYuj4DWJ1VfeIMR1NdH/iJHXsXnuGDcaO6OwycAOePwI7WX2UCeZwCcKcRhqSA
67VwBDIyf9qfhGxM6kMA12u0pxGdMBJa12nq+jzYLyVGlj9pmw4aZqHMXY9sSTF+
z+g7BSQhSz7h5QFcivVdrHEapfD7i7DzOxAzaoOkxkFAsNzny5eXWiiB4lVqVd2n
aD8jO/lrhCrvmGqrmQA3h5kLtyeRXR2NXJ7WraEiARgQ7IlC0mFhdm/0Xy+HnJgs
arq9gCkzOmRIhKbJiunpqhVIYZKxltREjjdczbJbPwuuwZcBcL8ulVtFDUFsuTk3
oUSCMNJvR+Iv3gSOI8cQPrUYXzXk6NBQ1+r24CDfO5yb+gz86VYPpjMWD6+j0wGf
2SaQmb6JkDbgAGOn505YCPLRAhr/LJp5jFkhLbiJ5c4gEyMRI9DnUkaf1xo0Uz0K
t9wg5aRzRuYr8nMWRVWvTzSAOOZ41+RKRhI4GgRA+Ntq0/XItcphT/FoGYRvlB1H
L06QGiXuBMAqHELLV5kAT9qO9RMG3WYJgE1w3f6rbSSaQMEblIWQzHxY+WarTDAl
hxvAO4Z8Z9i2uwQMyModk3YQ77qQozW4TrAn0ZQ69ILNawNm+q1TWJSu3hqDwjcF
gW3N/LiDE0IvdBzvKq6wbaP1xLGF5PS8Hrk9Vk+VaOhxsF9T/ieBPn8areXTQjWy
dIK63AiGkOqTJaZyNpi4cVnIr72uC1ExJ7qAXOQXsfJg87hA+0yNcnx+XSpR5XDM
2FE/t0Up56aVZnGRzQB0nz86msIBxvQJ4rnrgH45VCkD9xGXRoR5VvKoy/C3JI6p
l9v8IjlhJx06l/63fLiTgK65Lzb7tstpyyHd83VazxQUuPVDB2w2rTykTrWcaEwB
3dJNc0rCc3Uiwt/SPLuz/E6J98BcJ6Em3s+XvPvyUUZTJAYqC5ADWr59QWlLwGHl
/cf+/CFtMekZiLPbc9f3raqkLOeidHEDy+h+O//T+i3DcjWzEJ8SPJ5t4I4gF7tv
px0pGbwzTcDQ96SEflC/yFolxn6nJyMPhvHdEiZzZ2EKhD+n5V4EiyR0NFJTdNYK
JeV5dSmG0qut28jQBtmTnzpBCha3pq0iJ8jQ6SODEbJWBhBvj9sMJ6W0FuGB5rzq
84HFA8MWksX2NKkjGZVYYAclWHEDkEB5rW2eI5r9SBcRMTv4qEwMJ2yA5n0FoDvg
en4x+eiQMWsxQ0pp0nE2y+H0vtOZQJoqiSCMn7eSu7uBAJIsXtlKKFXn7trH48lp
Lbf+wWN22KSPPKfmC+56cJoTsHFOp4HdHaE03WqZzEmHHRDYBggU0K79KhH9NOGI
XjWFgHJK7RTPnLMdl7zswqfR6n1RbjNK2AYK93PvObwuNMLnODRvbqIejf+Cx7Zp
r/0gNtSEqkBM0mosucPy0mlQzyyOkjZCbNpnpNKvsFjvSZr/010LdnYOTOjUsdch
Xybw4+f2q+btkDmciiWV94qV6X4/yHsEQvRz6IPBPUPg3/+e3/anJ2UPjOhW9Dg/
S+kG7XAr2lSm+el4FJrIkjI0zFYHfoQyaF1m3caycLI94TI5QW0b94SHVJUi99Ap
+s7LgVORlXBm8mdrHCbgYi6a4lJdLCVSLhohTNk80WHL/QksD3FjMaNc75BbcSTn
r6Yy8VSYD0geJG1gW9rIYEcc4Ampw2Nx2hd4MoI3U20LXdnSNJ4wDhxqHRcjNAEK
uj8HH3MIBjCuWd6qdzuYp3ca+aMZgFcgBi8GlQpSxL/r1wHZYxjN3fUQ64Qu9PH+
yrR7i9kK4FmYyAGNdYAE1DTMluimUoqSjR+xVdlK9piSuQcQlSUQPDUpc+t/rNQR
pG5exUFcXj5K9mgEmJeNem5jJ0tBcA6Z/dFMDnO8q4rM+Q9jrwpco00bhIevxPav
kewTCfcSXHS+Yc7jn8JtOYGA15aT4BV/z9fHwQsprxHunZMs9/0T2Qn297xKmneB
Vp3OczyLYZNcmhMxx9k44iAjPxkiT8p+O6nv4DUzmewpSatghcNiBSRk8JSYBhSE
Ad4Fm7XaScdIcjxocCcOMwctVTgJXtYu1Kpx7RbwyDwgiUdyLyjDvFdatQs+GaTj
PQ/ED4hVkGsNNkoOxlETDtbVVFItbhURIHhZFc6SS/Y6wzj63CyZG1d4QO3pc1oA
qkYK1n//QTjbG2sE6N2bomvLdtNjKz+cPSwz6i7U+1zCz8G26vyRlHBPSEdTSiUf
o96t7KdyQlEUmta5FNpI66lwEulASnRbYfADiUil9LbUP13pGIJHBEWs4sOc7FTb
oyZtv0gPP7VPJSiIEOgrDj2SPxZ1sICM8caWOE5Y1H54/x+7eegARirUW6EZCp8A
8axuheClSR7mCRpM/CMQ76t8RL1NqZVUqj5E8DO5H34wMtR4SiVotLKg0x9YSt/A
Rvq7x21qyTbUyPQfKLPoLGYIEehd7SWv16aVfNRkyTpo7lOoHvK+Kr2EvEbsOkub
kSlSlPH9qq6DDYoYRIk9vGQkgULjrfwB94iqhGhE3Jpvlzkuva48BeudI1qXWxgK
/IZnmlxJLGeWnlGjinSyIbKE2dOvpncWpNM+QWAz5lLxMm9d8PcDMHAt4BxR13ZT
FLjmpIP861btHjYW32v2Rok9Uuh9VZLa8nFqEmyIyv9/qxpqj4eXdAqC5m/3oOGa
Vy5pfSaUQzx7soDfpPKcHkfaJATVQpK6vF+0sSh+7fvKcLxfMCW8yvuoCLQsB12J
NX8LJ+xpJsRYMgk/7Ze+p/QHDnETpggv2lypcj+XiUqUVeM3REEMuPuvNTIjAKkv
omGgZdl3gD7+eP8kZbL5phQNApuP5KDxo4f0SRNmUspsdFPNAAhFT5QdjpuD6Hsy
5QHeZsYzHZ2n1jBKwjP0qerHOMxMVCkmCjcZTLzrsio8PWEsR7pLOvpH3dl16gLC
zkLyS9lndA0wIeyuywBArDY87fSD2GmwJfPSXxCuSjh9HuZbXBs01JCEGbX/spa1
aE0wsI53wLYh6FOVSx8zm0MYp9HglwyFzH0pkyMVJZGLW8wcWLSKD8dkEg+dVjkb
b0sCbWSsYjk6ClrTaaVymV5B8BQNBnPFpbHDoBSj7+pYvhW7j0PAmjyMKw8IbXoR
pmoP2um3cTNLVRPviTH4CBRFpbdnCKfmEeOCqCzJxIOojjrUFNV/YETTmwr/0Wbs
h7vDm3t7H5DfifQof/mqFkNXfB0TsiYjP8P/1MooXZ0dPkdN0dB82PBwJye33yLh
BwD3vArDaRwRZkPthmjavJ4VEFv60DaLiOjyxJ94JoMtDIWaxQSd9ITvei5PGwNX
YDAY99ackPhWqwOiMjBYzIU29GTrpIiXUhDtDzNScVyCplVYrbjbOhTiDsyHF+nY
FrzENvd2a4PLQGaz0RmLJ5PEO4hAxYzDRMMWbw46o03QJQ7oklQOtiD8vErxHc5E
ER7cdB3dKSSv2sF1HC5wjMP1suzhN8jsDFMKlnKnWY9HqUausvA85jnIUNsEde/7
m40nYs9Ahmz6CxMWIls0zqc2xVo2lofGxo6M4tRiOu/YcJB0sa2VHOblz13RddCH
Yh/nnbf0ZphEuDk3xaWbKy2yAy3EZJ5qJXW7K/PoMrhUc8zbdxMC/Tc6SEzhK/mz
bMiqgUTfbJjhOdPoUVmOWt+SHk86wdAPEMFJY9MLbk54AYXtmlCOiqT9Vm2c6+cy
SEqTlqkZUn88BOIRpH6EpX1r0/hTypytLrh+cHv5j1p5b4zrh4I8JApN8YkYGax+
6MsT0fCKqBIbORgdfNFsoeY9BNwKuoEuxFKTdgbrqaptwj3cCm/GpXI4Nt18pdM7
v4LbtZu5b69PR0ifTgju8T5KSam7nc6jwZ8Ng4R1KDPSLqov+EuquOfSTf2qG8Qz
cNcL5vtQHM/cz3k4Jt2hznkZImAZ6/u8VC+ai7vqmkIYYiWvNVvRks5rSht8lEj1
qyAuSyVAbkiEveMugICCYhovsB0C/4Qiywg7tKeunHAzmdDWIVDF9gkGbJ6LtRei
K2pKoA3/2iKF2EmWGQmLxNfzll7m9afhoxwxGC6yXuVsy7LjoeOPpsEv9Bd1cl+t
QgwLBrylJOdv8AmaCPatpA4+bV98C2I6IyH/m2AyMR4VfZQj/VdDlpRp26od7BHi
wUqVuMdtwY2tzMguuJcUUjC9ptVOrv2TYL140AB7QQs2WapHNWwm3YegG84u1/1C
dgo/GVW/42bWqrqHP683vo/Kv6WjcQ18MJ5DrvXe9lMDnroIPU81MJbmLJwnJKSH
nGLLgpDReZoJ7doPvuL1AEIGUPA/G0INQXZb6gUIrRGEQTykqEGCR9VVapr02Lsr
giaAx1PlNB2/jGmhZcb+a0oUEb+wUwT0JJPzAFxonn4VorjZ7HQhL1N7kZLU+rn/
QF+VQUWiUx63IwsHLj0TVOAc8qXgTpAyVlfZf4XJDbCK61bEoyTaBFFDfRdVyTuz
Oe6nQTzx/tLe0rJ7G2Bd17Xc+ze4r4jB5tkESwd7h0cxBpleUJyEJpm+HmBrkkSz
XESVeXElIAaEgVmjsHsMwfkCRJoXccAoJlH5IK0Ukg6jS9VyU0oQ7nKDnuDCz2r8
iDwJYXkmomhg616FoUhAo4CEyOs/klewl/kIAidBqEdIxHdyz08GFrM9CA1x8unl
F9K/KViAT055qOO42E0KK6s36H3fAQ+p3Xf+v6fK8jA1X9A51nADmIi5XFa7IEYk
/F/zVvuOFMEwszUWaqZhEtMzxa1JcxN+3jC3ndVEMW4LnlbrYHbN2JIP2VOUxW3O
7Nw6yM8bpVbJR6djgkZjXXO4VZaBnxIv5Ra6ajK6zGSj9W00gCnuQaIloXRGy3p8
Sx3lSHcRdka8iIRI+qjQ7CYdhpvB8AuyqJ/ZWnFXPSR4vDuhzeNS9sOvlBF/c1NW
1aCLEp7JA4YKYK+Hcg/2n8caooHVhf6UPKR1sQb4V+SpItexhGoJIUsxwxqayBod
SzTxKifpzZokmT3DZovjmI5d4aaBRd7pBAgu15CnBSzK4ENZzlVznJpsNT8+IraZ
UfTkXQroEMXptZHGrKWE3eqaKs4UrIavqiGf7njyZpYZCT6ned3KMbV8L9C94Gla
khiy99Ia4ktYDZNM9pRniBdQu+wr1jTG8bvUe4AF1Y2O/zmdrRivBinqP5sqAeCY
aqgYv7ama3H5DDykZaG0nWbgJO87tN99+ISxwcABtes5W1iMtFSI7wGMOSkeKWOF
T9+wEZ0Zuc3PGqSa2V4fgWob+qIRJIWjXOMu86ey5cxDI/ftPiUH6zqYQq2PhduJ
tm6Tec0mPZ8RBQHDzodMC2wW0LbG2IgP7vsZrRhJXnFtn3U/URPch35Odgt23PuA
g0vT6pEvy50HPngPbM8uQjZYTHpuGT3a5c+lYlnAxZV2rR/xbWt0nj+1IyWWxRog
Wy7RG5m1DY4rGksZ3XdClUYk3CI2XUjJ3iislimPWkciKphvNJuKVAcW5qJuoFB7
7Syu3ais91iaMOOaMuQITl+Sxa6A3fFu0SjG84ezS+XT37JHFzg8mV/r2lyEo3Nq
tjG/VVhwGyCY60GLx0sDssx73QzwHZzgp+39weEzSq5bebYkDxII42hAmeQBpQTY
aIKKDAXvvy0FW5E7p/VnR9oxXrJoykVY1rurpSogcA30f5ozkBn6Rc7X8D2pUVEJ
J42UbcKmW4phd9dUOqiiQ+6ibGq3g3cvImQPIoT8qLupAeJr0Zni0oivlM5sDzp6
NhjMqhWtZD+VqX7Iv/8OkYOOaNJ4djRKIpPj8DZAKLXQGjn0jC+M+sWNBFBnN0YW
os62wmBpnlj0J/3LlzVqJExYMQPHCNCAuNrEdjPoXeQXvu3SZ0/ipj9C/RiEnMCd
uWKnlWBf1nNHY1gdVRLDjo+hU3plDOl7xRkjxA5TfqRQFVHLmVOId2c3Lvv6TeV1
1oRUOOvWqR0Li4VaUjaXcO7bhW3Tu9JuMB7jU3cO6kRbDxIpcToxBUdkxyQc98Hh
e5o1UpzSAXJENvP1VEyVd197FFOHtSlgWk7PpnKmebmSuxlSFz4SOtCYizUHnSYU
5SMOMnorCT7QjvDXeqvCL5nX2eAjHqVwwO8Lt6xYeqT2rgghfblDGZwRDJtNH63r
VaPaiWZr967eqQEO65rYGpyXORBd6ydAe+OCOZRgQnFqMVuzmCdkBb4mLQWylUrp
uHIi0vNN4UqMPzX0XunwsS+I9uM540S/fZTvq0VtDDLeJ659Z2CKJMXi8tj0Iipp
+PgGWDJWBo0ZaKOP+JKqzrqezq/dWkWhjWx7sjXfij6hiNlFo6ukz0TzMux1uOF0
qzlZiO0Dv44JGkWbEj2zVLm5lrRkGYgl1FPr09l9jd5ppodBd405yMAKvcp88N3z
1iqY4DcFKMVQhasHPXOf5s9ey35uBOfUh+Zb1vuxpuMGDewYl3ryChXLjD+N4sfe
rDvw1KuiIpNkvjFziVSiE83RWMqpIhwbIiiCQKkjOXhEynUFDZwULnxXxqAGteX0
6PyQg9iQNSKjfMTNyBIyALdhcBNHPqFNT8SE5lj6hyZ7eUMoRUTEslLDe2itg0w8
mf3kOlBBB8PuN7KJvu0MS6qOzWysVnCQ/yE3IzhA65hDX3QFHieskfEqSVcY0Xcc
wKlU9YTePJc5ALg5Qcbl/gu3XdeX8gcLLx6kgycGXrM2YRFW0/uBmf6Ak7E5/ZAm
1/eVFmBpBnJL6BxlYPXrUDYEjQ+T2ymmnHYTzM6T9MXY4aD8elB6ff11euyXvo7s
X1HFFCOQljl+YUudTN9r1vJ1akEiuj6V/Wk8cf9UvIbOuWIzC4w4sZBwA8b9H0kp
tLMlpI0bqo45KQLJatLujOVFW6gMfUhUDr41cZE5bchkffUN3lHw9SkSAjArUFQw
OBCDt3I6jIPU63tEal6N6zsdVRDYN7hr9+s8mlsWy9UqWsTtBikeHc9bPkph8AR3
4SL2titCFAF0pp4DEXP3wNfoL6z22XbBOYaFKpiS3MJJVbTNV7nXUGphVctig3HC
wskdYeWGqr9no9C3mAqqZQZYRfrCqACOskEVPhvf3pSZ+BV3K63A9G22dl0y3Q1g
mK53tHqyJl5y6ypAFaQrsdlMQiciAp1ks5uLnu05INri7YCHLsBXegbb/9TOmrAC
KdbTeE/4FXZBfqa21K5sH8lxldjOsiZWSInO2hhakvioo5vdjZnI2ADY4u8plu4F
D6XAo7yYP50OT7KSXqjVTOikylHcRShNV2Cdo/EYlp0PiCnlWX6ED/ilVglvf6LO
`pragma protect end_protected
