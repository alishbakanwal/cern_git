// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:05:44 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
AdjKTXrHH+rQtj+dtqv4wBLZ97vU46Omm84prH/zxru7ubQwfhszJDGd/FsLCrRp
PztQauiqsAnQbZDCx8ZiF2zfeimKxdh+DQorrjK/zaLAgY+IlrLhsd5WxJqenxVr
pqUN35qjRvps9wDNSixhqqExVjvwYcrKLDrGUpSN1D0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 22448)
JJVbKtFNTM4+lpHV0mPsCZyh2j5hwKVlXDvaM1TG73pUuFKLk+mODMeqVhdaE5LR
P0VHBQvBHs61/UrYdvXU3W5vYAL/hQPEL4s2meHSze16ou/WVfkemrPuLCzGFXXu
jdpUv6NloZfObve/s4zr9ltqqaDWUEybxUdMNWQB/jrKVdA7lw+3M/Lv4el262wR
ra/GL76LS4syoaFT8/2/34RcqtlHKE1m/tFj7ATgohXZ/d/CYFahQaRhubPZ2CYU
L10A32I5mjnOx4eOvCmEdnuhIfo8dfggNpyoPswJf5rnNL5N0L1890CutADvs+CG
pN5ToiF+arZyFy3o+/bPa5KhPyLXp++lu4YAQq8FqwSRk8/EyE5o7nfxCLi4T03q
/pS9ZNnTlF7ojTc8fsNz+gN7H6wHJXSOPRyHwW+tUGAKkMciNX74Ig4kZPtpAhjm
sNd+9h0mShHidbzlPZV7PHlpPRNXL+gQxkF3HS2UaIF3/kIEFzPKsYlYJ+JrJ6QK
MCAgid78LLXG04OH890lpT13ZIHGZIjnGlgSIijQioJEaVM74jLcIh3dxpTXAbjJ
lbcCKaJ2Klx1Qvm8y0L2R0lgDbZdOstZ6caCVHo8KY+K7UvHgjdHZIti2wI52if+
AzCJp0V1RaYY/TmZ9uN5zP4K0XOk4FGhgGlrWuG/OKt+FXM9qdLd5O+ErL7zMHEo
uRPEh8w0ToZPlpYxnEmAiP5bcuKAYFjJE2ebH5z7fxXcuycL+LuhNP6IDsDySW+q
OAY1RzN7rJZXlIP0OXN2jirwTJJexYywisn0yjFjHnea5k2akveaD/5+XbRRZ399
DQuMlbNyuWgUQKgJMrZjsiZs7A84YHd8K+DryjKNE0t9fwzHmejrXtUZSkVnChOa
j6Z0IYbs99N0x8zI1olV92gvWPJVN7+11XgUJm+AWz/coSGBPiE23+gzSwQYxT+z
yBIMfOb8EyYkVKF38ICX1oWQImvKqnxfwpYxtLn+BcGoz5YJiCHyMRz66DIFdc09
fjSB94HjLwMVv1QRHWmEzN5bSasqJsrPs7T4muIQztu0Ohd77fw7SJQbhq31ytDl
wRqnKHBPJz7/FOq5ZDCdSwVNywMW0GA5W4JiAxcLjuKVQoLoSnrM4ihovSsKG5W1
p0kdoixuwTRhk/wPfPTyrDeTjo3xwJDvdrba3AFDgqqWRRa6Iw0xPKUkLB/B1Xo6
xgs6gD+g82gTS4A3WG4Odu6Zrx3FDm8SZ9uN621mnGKDoQ1a9mxJRY9FjET/CugV
TsRKjp5RDaFlOmEpwP+O4H4GlSXINmTbNB4fKy6nhI15UWXAcMze0MpfBKiRGs/M
mM95BWdcE9c7D5S6t9A5yb9FL7LJV7EMkNPFFB3TQBAAXvlolQH6RMUD1pBMsYad
M4LCBdy75SQWQ2YKg0HZXxTjomoZXX4TdcfgIFtSOrRJ+JnyeMZAzMYhL9cdnsHh
LMFM6mjyWvsSCq5V6QGbjLY6D4EB30bI18RSUvvhp9BkeZ7vRjSXCenIRwzh64JQ
nvJNlsyYB4RW1MfEklgV+qFISqxJdaC/sn7jVEXZ/I7PbLeQYSogGnwy99N0NXXt
JO8g3oj6P5pq9LB4bZ26kiXOp6xrHF/kXTWopN0RwWM1km9y/HitjeS6sPNzvTup
XhBhY1dcZqQAgeiDMOQOcIFsTLnA+isx9SNeGqWPC/lhhewJIrmZJvnGK78lvvea
ZyOld7FEUu126T4fVz/LV2mRmPq6B8P79YqSuSoLS22FEbHYMEA8UOQz+t4cLaaA
+23wL5UKGOmy05fcJNvpQYRIes3W/q6QfyQ5acfcmOpIt84/VIKh2sOrt6Zh/dF7
a+zF3PdvuWa+G19F2/ZfncVbbBWrF3m0B0pAGBOOdnDujkl3Lzd0PsOxeEBOwbkm
RrEyqlEUtvEzkOclLHrR3DgF8jnut0Z1yYJuke4aIX/9sJsjH0N3rMgV3iZF1UzA
pObp7Toxlw3YYn+iYQQrJ7d/rmpDUSIJXMWvnI6L/hlT2tJg263EA4sA+mOPpVML
0r7I6JfZtIO6vZOIKYHpaAO8PSDQwqg9KPnPDcYX4+VOHXrMbls49iCffMb5DRY+
l4hQgmJMYwi/wb+3EjmMb1VWW2zvZ36MlLbrT9Yp4qbzXd5u0kJbuRdu0qzTewZ+
eL8UWNNT63otyk39OTpucvCy/GDtAR6mNaq/6uT+q5FkD5gGj4e5RodVZRtUBx5f
sDp2MNIHHt3nTGhTGxNZ/RR6B84GPKwv3GmOMshqwatusfSGHlZYTtg/c7ECWYW9
vOyXkM7UU/m1jeNKq5wkdcc9lTDwcDccgRA8dE9guojkZqfr9XS9cgTO+xBXk/Tz
g4IBm0Gu+XEcTHtB0AP5osB/wEMedNvO0Z9McKzRsTn7yM/dntoCoximJikpFiDI
xEyRJhAac6WMKVqADrbLPRV7z8IqupdNb7ZkNllQZsag21NnZMVtswIf0wtimqBF
fgTGAh0oQcwyhxex/IWM7gbhygX99ayjqvkB+Ea5jUsZ+vC+EgnEI0nSf9GdPiRc
TsYwI7rxUaiZBEwPryNeXB8ysRTs1HM4F2XnKOkqQBDVqFjRIn+dgGmZGOqO5/q7
Rfs/tRIFYqGqyrT0O6K7HB9wRKlIKxqgLnCaNgWkqX4Tvsl6wIzAnmOPzDF8g6B1
JpySrE751x2HSUKq2IGIXP+A1QdNl9RJH4LfuSDMM1iNgQ/+Un8Byq8nSZVyAedG
PDmedo49/H2/yYMG3hjvmeLVnvrmK2qBjOt6wTybDr0lWPIEOUSRKUOHRbm0vB5S
uymUYPHIpkpMBMJdqsy5L6jRPqgoPGWlcfrBDl6lQkagJMvMP3ecI0fOgDokpG7A
ozGN9A9dNfr9b0ei14STIixNBg/ERMJoWrrKw30nc6kRAU0V+TcAz4+sFdJgAcMV
RbwL3du6jCc10FBM/+u+U1mfVSaS16IGVwRwIshFaZO2ZyKVJL6TQPjnGVI4Gqi9
FkHxQMXr+WJBCJP55K5tUiFQOGwN5CcV4btbEk37OZLC76KDR5rqfxbsT3MbG5C2
bVj+K6Ajg/D6iFpoxGvJ+KqnbSwKYxl54Ly8ro5igQa2huR0nPiXZDZbv52Nyxtm
c5eX6/2N2cqrdeHl63s8j4VfOsnaoKuzCyF/Mjangup9eoA0PEd9QH4u3gZeC3lT
QBwZRLwZ3OZ+cFWY/yCe1aFdbscWoDP9ro274jNZQ2UaawerjQsX/P80VWoUPs66
jQkluL1NFq5Q5QQSbhgeUmvd9mwxR5p4SsHSlhqpByMoUKbxYohxm3X6467mFT4N
fybpotyyp5Y3SnWp9fXg4c7MPPd8jaLbVs2AHCG0L2iGYB6v2s1Mp1HfpoH9y2oZ
AxnX9NInjoidSHP9lRtwOqmyVVOADyfOOAJLa6yeaxQS758zeupopW6B4MF7pC5D
ZKt4gCcyh2BgGMMAJa4BXYfmcK5hbqXjjQ3Sqs0RxSofVXidrnlU0IvIVsAyfZPF
P5bM8lqB2WSKJvEruMA+YU5v/ME5NRwLLPghOSr9wZ1PtolVKMtAF0J7vIjdKhPY
pVCu+6O361XMy2Ewd5aZlI3DlDimUSph9dOYJNP8Kv0Qn6S55UbiejtVpBV0twt2
G7BvyZT0NlaivuB5zGq6Jnyq/1dVzVBCsFwTTZk2Xe3tnSUKy9bMVc29Vp73vl+0
h5aCqpzg+dgx0kfV4HvBm7OQ59VAA8tOuWD3aBSZYYQn6eiZHhT/RelNnUDBWWBe
NlMHoawC0Rx8F/p+GAT6lW05oAd5EMsqBDzBjOEfHCNIrqJMEy3meRULxOGRpjjm
D+inQCOZH1taUPeqzpehyLHVUWIbe049KlRT6GCdja8oEj5rGTl4tCi0WOU8W+WW
3sFPMdaUG6aXR4ihBBsUbmZM+1iMjQ9UzY1GB9FZALW8CvRQkfRswR43ocRhBGBl
+3M5CqhI7lhLne2SXr2qHUIckzTK82yGCULFoqy8YLZHwjLLp7v/O0lqpmbV3nvn
eV01m+1/c8+OC1w6pcV3bYoVGJOYAS6mnexGUAXTfnAgGPGQD6vnrW+l7u4ePxxP
4djkg/9FKx7xrUnPghRDLZgAAAD5BIExNpKDBjA25D769GT1Yeyl1N2sgZ+6oMXV
I/oyHi7K4Ltykmi0cUMJeQaGtSM7sU2ZAH88sTxEnQCvZ/gapsydJgShoYJLdTr+
sYmUO0fKxaMk6Fa4uvXg6Gw8WkZ2qbjRwVf76tQkq2OuxsIlJDLfyh1n3grK8E+k
hsBuzaFlXIdM2SHr/3BIMV6AxBc+Aiv9pCmv57h1KUsSeA+Pkz8iMWWQu6KV7866
6QNb1OUwmBG1/1JkrPaoyKhjmVWe7ofjZzY/0Lvaz3qZMmfAcC2ZHQkW20QRbk5l
uMum0df3fEGGOZEEi4JjOp3hNRUrOl76EqD/f8m2MaAHEs45q/OidB8FcL/GKU9+
jjb9emQn70WnskXHy63NsYchoNuqZHugezd17hbkT405V2CiGScV4v9vi917ath4
3G7VFpbpUm4KOBB4FfMsE6cC8BVvCpAkrUD9ofahHIdBdj7xDwZQKKPAy1jukpJ9
fppK0p2SSbGUfpkmF1Xxsyl1K/12+699rNo1ufNBwH+SCDucyHwMdKigu03rb8ll
J88GMw+XJiTWzF5CcBYVratgsSCxH52NIJNXYmBwYV/Ehz+lSwf9zKZcyyYWSBoN
LvmpZvRp85RmQCbckGxUqbSHBs/8lYVg57m93OnD7SdHsm2p3vL5YffI1d9w1y+m
Ok4A8lU97C/uc6Y0cZlVpCfm7XuwvbWtR8d/kRm5ApW1Wb9lxtba5FGyWo3qw3P3
HER/mrIh2VMKtHcDtKzc8qPj+1w0FjSCPt+nOerxRWqT83CqvxCOSSRsq8pW5oe8
2m0FyRZMDYaoZsTvAnM+HuHOjzkB6937RMKdZJAt7IzKmcY9IS6ysVVhO1MNcuTP
SGERFek882jakzcbe98jZK/ubdLOVEk7fAb5sDY0ekfZWHBITMuAd9jh223nZoJA
1TBQkDonQDvb6Q+CIhZy95XWEE36/eVaAtY5oowmiUXOx7dC/S7YVfMakIDPIUCh
aX137ohQbezIBU0RAlJhgOuegbygY0fKlwHxQ7Jir0JNxarLRaRgYG6zK1WMqs2A
h94iU1S4hJuDPnq9bLLCI1q0PC652SHj1TTbzaN8BSIa4qOamqLVEu1LW+Q9rDrD
upNmUPEGc2jlBWw1beYpV1E4SG8wpOzb7hPNf6f1+wOYqNDF6ukhNn5q8eJy+7Nr
sEOdwk9TUhV7XiC0qcxUSFuGjFmENsniCh58+MYwMgk5NCj0+KbaGjg8zmHruMfw
DHW2WPmI/tRE/lVjRh9OHPmgmWTYUGlIWguCXxLgLCo2kP2SNM1wS0A+B60eztJe
iDm+/OqIb0/t1LptoaSOexr7JFFATKg7O1TJlcZnxoEIkyU+6Tn120eN1B5Yqtuv
T86XK/+Qz64Lx0ysTvc/ij87IA65cYk5pfMPjp9ujfjleohiRMhbDJ4UgSrPqTf1
UCqF9f5aSouFC+feqoikwVgO/ANgF+drtoLQkyc4EgSXyK9OAAsdfTDoXSj6jBt7
15B1i2ZmhrChpRgUe1TI4YYsrWz1yxhgRBRvfltNDQAY0gE6XUJXLv0YwP4GNpiA
bdg9Eu4TdTr60XifBmMpLFkijRe2zcnTeHvDkbAnmpmHj99yISdvVUXTOF2y9OI+
LObDbI9RAsCPu8mFzJzGLu6LucFdYUEBclQs1gpx2uJjykh0glVLPMOPPkxr9mpg
iUhceF5gX6RbeYvS8avEvX2EQMedL2OJxHLkCeqdlX0atRvwSr4rGKtn2l+8RA9F
SIkAtwVT7WADHezBE1EO6sSeSRDV4bNyCEqw12aKK6VIU51D6bZq1taHhledIILn
zu5FwBEZaYriVa0dIrXFKeL7ReM8kZ95m5gq3mLa0ndsrY8E6LLZ6n3FMpLBG8mG
Yua+XfvDZYE/AXWBUW1lpoKODh7phXB2WQN8kfIunF36u8DtSPrNjEBy35RcptcW
955G/Wra3TrHLcYM0cRynJkUJc3pX6p0RGDsB7hCvAKZuuV/7/shNBHRQFuDoGnI
QRVtaTqMC3EUmCsJ3e0oeIZ2Mu1DJUaH7n4sxvZRZ4NDhFR5pnrkLEjy/6YnEBZz
lHLf9bGueuRgyJOrKqHZPZy/4Am+et3HA8tUZbf/qGtn/dHvRGWK70g8S0zArKBg
zQg/KeYMobFIJyR9oGJxf7PZPmE12QlVAhTDne7IDDsL+TD3I3WqJKr44C6X2dZh
m7i69mXRUjGpUHZsRJlqKYbmB5q7NIHmIxIYpIhTsSM2rbpaV/bzh3AI2OLWtl2i
dQJUypMdG0zv8oRZyJwqejaBVcTpzvNEelsKF/qjaNLpx4v/3UOBkunOwHZU4sfd
Al/OlkVmFjz3G3JMawV8aEJqP6kc2KTLJofkKeEepFaB6e1WjGQfBCzuKL7nJdVx
wB3PPjNyFSgUDDVBMcEabpCykobEZ16skD57m5OyZQLhRX1xqBlHX6NiKdAFjdnq
RHGZxj8NDsiKNorEvJuul6yh1pKJBr+jcfXs98UsbtO7JW2BVdpbsNcWDyNVVZMn
1J0cnyjwlTfZFZNfSIISYHi81wPrDvICt6fq8oSCP7QfciYOSpfAlo+TCHSHjiVn
HIWXmCIf1Y0vWk8yxOMIIe+Tk3T7mijGdNlsM9lh6/IDztM3nu8+1Y0ba65tx5kC
sVjRfsw1ZlYaKrwuDmP+eDOt3rkJB45yfFxSh/l4FHCpSf3rrvI+BHrmAdJy1bkf
nKegK3uIjTv7YZUBkd0g+HOAW62XK64Cfc1LEmvTIRSitYO7mds2H/8Wp9HQAx9g
nk6AuBfKacfUe5Qt7G++JXW7U5jQDdDtHBx/pwQu90hEL7m7YXNDjplDgeshACrx
YLx8+EW/XJ95kJdE1oPVhsOGs888r56DFqjsNL78kMzetPuIb2dXL3Z4G3rud9wo
sD632Kl3I4Zhmx6araEGNaFF+pwhgdijS71AIn34e0mOA/9T0k1T6WJx+qMAXu8H
VoGZTKiTXKoCHtBL0OkP4P0aS201Dl/aSjFMdE9Z6qNB+tn5pDGxSjyBQ3+8TFUo
RYpZj0RDmIYKUSAb9/VeX23naNOkDZGwOc6b92QwbPmzkb0BM4zsUDRG3i9oeNMt
v7xFFEX4CJkMylb5lkAnfXWauacPAU7lcTa/iWFRQr0r1A7iyorks/Gno/9gM1aP
8I6uB6rTYL0Ft+z0ldtQRmbzKnd6qIuXLILmpmdp/b0iz4LlUmSDVJbCTyL2ndu0
jLfU9jtrAeF28UYFO4QBTzLAcABKkwg+7RHD/2qaTSpZtHfb7V0J+D5sijqZGr3i
oK904m43wWLpDI3Vpi5AhZ9/D5dEdkg8Qw4eRXMc/o/ovqCIxxAufDPK0eUOygaA
NYecxiwPbXhSO+yCUsd8WC+ZHG7k7TJDORzTvbA/+bPuiRwHPwE9SRX7fgDvtA/X
MlL0WLbKUo21hmqBWErrC/yv7ZWozvu/FqKwlwzeKddgNAf9kA4qi+HyNHXdMrI8
MTkmo9o2zcXhxQ4ch1iu46BfWkWtkQr/GAJpgZkkkr7DqtJ7bs6d5TD9w4YojsKy
w0yZQ/7rw4h/CHTOuhwLZx+1mWv80lOBxTVUYf6TqWolCLoXlipygSVf7e0DNKXf
Qsmz42SLDMPYCiq2+1jDdayGq3c2zV4+Eifbd+iHGhtx91rLjT5QYcAmiTilKeqA
yRTjdf32TAPozIWrnOVvnPxt3wTXYzF7oxDcHPdsgZe+RJLSx1gblSDkuHV9E3rJ
tZfKYo8Ve4VTsHtwK1e/+1W3X5LizJtbhNYng3+E/Skhb5BthL2t/V4x0/gUoP6s
4FK71tlapE4FtsjrIVAUvpBcwNCR31G2tkFcWiCia7S4nEDidKwzRLlmXlQYEZDl
SEgTO1+8rkRgcivLDcZXhddYsA951+SaH6DMrxYYkTRq0Tl/YhKW363zIqz+TruI
1juOc0u8WlIBMRSvGvsSFIpa5PlhqIaaSrZCKLVSNBNc5V9UiFb9E0+lS6PvpBjH
g4CI32HMdWdsogbpczA0TaFwieqjspaKY77OE1jfnTdx/wCYE9b1Pn3ero4+VrUZ
Bau5Nokytxd797W0FdAVJXgbkXL0ZLO0wiUkNr0herf9Sb6EPWsPJys3piu0IT/x
ctkZ4LzlqLVFe5XS6lLN9hX+D8l2+hpR/ljruZ+5M1GzRsJFjz3yXlITjXVjcvHw
IdR4Yg4eiNuAu2j7RIWH3wG+AsOQpQH59Ch/CxaNYpd1n/D5R2Lkh7kGLerDl1pc
6BfuX8hq2WaN/YR4No89EOiBxAMOgQlTsD4Ab/NqXqgbt8FybS9/nuDNUmKdEDkM
QtMIC4X2id1qvB8jIw+mzNoJ1rVwD7EdyhgnmjXA7Fj9REiBKMgPV9LzYmW0Kh+0
ykZ+j0nDGzpLhzlRfSCwvvVBnWQZ91m3AFBNMiIP7qJ9gmHJLe7UvRiTOmAKAfQP
nO0A/DAMb2OjaZsKasZOlFvUfUP3JIuZ1tDGr4WEZsQ1CFZy+WCAurMmyWjKG1ve
URxQtXTxINTjZ4wgo/7ExhTmrie3LGX3OowQTLCpCuxpeeC0pRC4TU3M76ZpJgSj
sbcLxsolYHYwYfJIjwDNhcbGx2oWco7PYpZTv/H4RU/TBE4o2OEyCkHyjPbR4ao/
moabEkfslfo5n5UqaY//C+PXRGH/rSKvRY2jUh5A5IG/K1dqRa9GW1EQIpNkEkI3
dqCvpDkoknGtExBVZtP3ByokSnNzoBRoS5w7K+Oc6gJ5PJVsC3pyB0wf/yPv6vQv
Y4EK2a3Fbhs8OOF2VkpR05pdLMDCd+SygV8SPk8hcVbk4n0w2P41WmZ91M18A+Lj
Qr0KQKYXnr+pXXvlybXtpbXPmQQyfAtvG7s20022OUfsFngHdk9G+lJbl4/ztHvQ
BhF+uu+2XaGwfX7g+bZJFkHJWY/oTtLX1mHGuXQTTc5vZF11LFcYwXjOHenBv5/a
13/PVWhoiTr1Unwj4yb9P5GIHeaOPVE5VjElHVf/Sn7a+GQrWzY+MNYfARdV16AQ
DTF49rfhCfoJosDBXWL/IZDqdI5FLqG4yVBBTSAXs44kd8u8EhxSUC/muWo1LeNp
TPsvSvy7PnbjTKgXrsMenRLGjQjl7lpH2HrrB6W5s9jzZmowvcKEZP+9lC39DiHG
m55j8bagYREFNDrtatnXauHUH06hcI8+cEHI9rYkilSUqEnDvNn5oodSK6akUZcd
rHxuHShJX/cer7QbRIT7uXE7wpesYGKrMKMGMV1frAc1ogXOqPN1HxgbK5SfVoao
ht6aq/fY78MXy8SDZs301S6opO4rnH8Jieynj0vxlctircPKEsTMRYLU+14jyDMI
woB3BAbIpc8HZVnvVd9R07NhhAbzdXY3/YN31vp2PH1rwOS6Hi81KuajPKUWq9Ga
6fBfAX/CwU04Y3Snr56lGzhmiKHtZeAW2cfVE7xpYdDgSYrwTawqNKw+N+x3W5qj
M+CsTi/njvAgY1eE5Vcj3CtnlAF2i1km4AWsXolp4DQIENMNfuG6Mjs/CZjUXvsF
bAyWsljsBiQT/GvoYKuI9Y5lAEW5w2gwgYgzocig97naEB+nORvFMLwljZlFA8d7
rjnaYG5iI2bgFRItxewkBAmB+Kh9FpVTslRIBUv+sXuMKzmLZLaP7LJNBVBD08lt
68xypr+xOA6wz/KjL84DqnWnBD6SRg+TfGsadkpmC3loDEAxqjtwV95mBNzIA16Z
EAc/vOz6PG7vzYo+R0NEiHRN/7o+IhQry6IYPcbwCCCmtCUK9UslyskLX3gDA3Tl
z2TCqfJJu8TU8HSkRkGQaOB36TkjJujuNa5SK4EMFgi+LqCyAlDZpj12iYad4GPu
QDgqWCb8gJH4QLZfg4tJrDYM10ssJ3cFvgvtYWfCR/QsZ1Fa1UZcIXRAQ7NOHrQt
cBJbKB3AtoSCokrAAQrkB7e0UjxiSAC0pq8hziXD6THZMKgCROze34XkF1PmZ1+0
DSdXc8xNTYzKJma2rFhBiJXnX7WmBiVLPkAgdAZpzTHIQhvzlRPwY3CPrikZP37H
5EVRpRzrVMxxI4N34U8/b8RB5dqHw/6mqW1Yrp/PTTO6xtzBVvoE9vHuBSaeB0t9
5/KpGfsxmGRTsCoe+wyanuFKmeR6wmpiGrDMFerit7qzNYyqgm0nXese/INGqu8u
Eb6QaDO+d9zdH42gR5b2IdmEsDPDx4mN6ujHJ+DockLQ7rorRrlCdDbrXhujRQ2d
LJ2EnKA4KdQiZPW6z8L34P85YTcpjVs2VNR5fKMa/iVLKExDgnyPJ9cj/TP94+WZ
Z1fftzyq0f5tsIp1VmLBkvZE4cjBaQkK562BZ9wRbgLvEhNYOM26RTAPAY83W9hq
cy/0WCSvHF/hxw96A83ip+y3UO0gOQtW4Td5eZzziBDB4LkAQwferVNEc0Yg8pAr
0xm4cpM71QDviksj1VLDAIYtv5cnYgd0xZf4IutoWvAFLxWOp2K1UHjdYID7n8UE
9QQQZn0BmBrREpBMMhcca0/OBUh5DTpj5L8WzXUB4fWw6TswME4cFhQRRsx65kUq
KCb7ugEFpaR27x+lTyZ/BsUWClph4vJh5g1R2q5CQpH4V7RFbPv1y3bnkWBau2/9
4VvhZTj/EJSgI1F8+n5nfX/A9LU+K/BUzFxnICcuY/dq02T3DJhuqPi2uuZqzSWx
IZWf1hbzXlBpemvBoHds2d0Ttt27fN9Odvc/15vzmggau2d1dwW0AM4nde7VJEoM
wvVkBon0BxMmASGBF13VX+IQ2SxJ0zwEygWoS1/IvzMa1Rikv2Z3M+Va/hDgl0h3
SL77aQaijDJ0FuZKP1IcFjjLEE+dJSk2HwgrKAQHE4QDEsMeFC9fSzbGSb4KhYTO
Bk0byntZQzxZYTtU0CYDfhiQHvkUqbPHn358qtmKcGVpf8srsQG8Obb2b2AaNm6o
TK3D87KK1T72L9ArcqZsfu8aRGipdkytDk5xZxMB7TkABTapUzixgCR7Q8JGhHGF
/eW1aVPVPQBr41rX4i8xs5B9hovZh/N+UNxjoakHaztoWYXTl/CvEX/wYkvEj1Bg
+2t37LflNFKQV4ZJTsCIZztpGvSpS0Y9RhULtyRuCTVuBq9dUrxpFax+TipQKj6y
ap+2omtBiy45/cXYXs6QPw0bua4FZ9qtJsmiJJkWSKtsb/sYvnJ6nvKyPDXM1MtG
XJuFF7ibBcgKZFxzBE2pi1GU5/LKFzUF7NRIfzT/WL+n1LdXDff8zpBJmJ5MGU3I
z4yzk13B8ouMROBAxqDqUi/YIddejVry1gx8PZj638XIsjk7OEj2fA+PTLyYmkLY
7O4aEGNxS0F/cESz/tpgmVcO1LmlUvWm0HgJ5qdt58fxvPxk/OOHu2WYmBG6zPLH
+axRb1voo7DLannr47e+9TFlNT+LhrDyMN2imfmnpa2lY+ZEpkFLyMiycmch1zfZ
OBZ8TEI59yiOhir5EkaMmM+MNpvrcWumVD57vC4qYv9zP+hy5TbNDKmdwaxcYR5O
9T0EwEq8m73F2/cpn+FfpwlxDE+x8yBON6NCCYX0UrauwJReLPuNh/3+Jkai+nDb
H4nLK4QaNFebh2YnHUs2nm8RoBt6qahhpXr7dQtY7ErlZajH0MuG2GGRrnLWW9Yx
Q6KwN+0hHKEGGdNPBfKuaUtfP8AyEJT21K/2eQQ9werQFs6m86SbGc55PucHCcsU
NybTcVIGEHxceOm39cvFkM+EUn8buqQjvNyF5/qTQBhGuH4sfoQTDWPDA7NMjNgv
6aZz+u/z4LGV54QCCLtMto92CzgMML0r5XU8RYQnaaByOY9FkpY7fhanyQyPjX9/
PSJtN0G63o2kEhdUs9aw+QLR907QKT/Av1FDOU3Y4Wj2liRnWaKIwM+L6SdQtkex
VK6DYgpslHuTOGeUF5X6njurwtHMuhzjPPBCWQDYwFMAVAcnX+AR8hU3DCQB42BR
kzQ0MIHIZ214WhC5sdX43AqVOiBGz+IWjr1+3Yoe0jwWh+O5+6XW7cZKfcUOhQMn
YJR5WuFXN7ZGnRgT2KRd+jCMXW+f6r3TmXeHxTYBPAK6qS+zqZIzEBfYQ4c1Kjou
jEqRrT2TRvAugPlDGMh5+/v/MXoEBwfouHj16F4tmaOt5iVwHxUF+vzPEUh1DHLr
JiCoSNoQc6Ho4TznmN97/MCa21yP+4PI8T3Qz0Mxdbb5gYqFVrpX7+0sOJ0EB2x4
tyZb0sBkdEjzT7B49bc9SVoulBkmomJa0iHrqP/AN7mXWp90Abnc3WXNCKoEAqxR
qw+QDYYT0IzH5HuYZkyi4XbLwcJnm5N4wX09L2MvqfVBYHJ9b0mG1/WBRqDKPyCr
VQ0/PqshXqX13sHcmus1oWG1pEUBUEIHxEkExk55v/yr+LoTuH3vSanlCFGJXBmD
AFhyzhon0AORl5XPR3FRrk9qn/EUtUhdDrO7N/lnPuFUEhoncupQ0SlFr0kk2FD2
VUGAohSTgS9sp7PHbzhTlwzTpyl2BO/OfT3DAN8weOCuxyEeDJC2dxFazQiWQkMF
FwsLlt6KGN0sGrWl6qM50XMY1kbc9Bx/NA8LIGVtWtt7iD1pYJd/+JXfjwl/K5rw
KgZwKs+SFwFaVS7O3Sv3gcgmuKKwSXYJjQk9Iidfrk80oLXwSZ4OI7idEV8HjAIE
4s+m/1xx0obDDqFuan0wDcOCPEynGzBwaO3gnb5HJqu4OAko77UIXXYEOlOLV/vy
Tk9yznRFUF6ytrFyamLI2TjKNcU3J3qPtE7wWBjVfX6pUdEZZg/QY1FOGlNlEIYx
F1Jyi4dXefTe6B0UHbDa1fR3eeGstO0LNL2vHIjwqCXVSridGkK+4N6y3VflsDbL
LzVANzs6Txd6dm0XYHS5XX2sRzX4e9ax9knlL3wBJwzcke8ttNeA+u+BOlez6TT1
gHwk9vR9k0Em6jIeBPsN6tpCbhCmqjhf0BA5onjjZLmosgRc5ajL8OZ07WEbMcLS
QWfAEBV2vEf/ehLJA/wj6dm1A51UCOAeXwNxJgnj9HEqI90xRerfmvX8Bj5WRRqu
yppGK697fyKanO7rKReYfb9GFIw8xsMCgJBYU67a94W47xMFxzdbZCwNL6HNI0x/
lHT+b4UgVEej9IQskFXWXBPS5jB/eWCtMnBgAoToYRncZDP/eKtb+N22gYu9lSG4
nGDJhFc99ZZapLTcfsCiGXmncQdYzICgDN3Ys4eyn7ecvUb3tmdITjt2zLEtcnej
olrBAOsn79kFfLLAwl1xBlY73IYMWJhEXmnp3wGQMjr0GhIDpeBinXkMU0jXPJtA
zymxI9NHbD+SVoceKNsOLZINvGUEXPxG8lfmo2STqMccXy9ZppK/dhg62BbhL7pG
WK8aRx7EjRGnX0pPGMVvNhwqvm5ZyQWIGOCggw/XLEi2Xf7GHDRa2r4KJ8ePkRA/
O9zMXpwXT/vyVRAq/ac1CEKh8BegbSxPI9+UTwKm5YWTjphqp2OxbaAOAmNMPMKA
RbSh9590BlkSZsYILH8vitlu+tI0GnlZ7sORgZttiLZF1YdM79zPf7igXQFnGi5l
6xoSqW/BqLV+b/EUi6vUtwm/dQ4C20F7EtXGmcEp7JLyEe6ERuYfnb2c0PR2u4VL
KxQ4tSpWaGlBmbiXcWI7atIVcPsGGDVgmneOUzok6tC4QKN4OzXdlL74s3zSXeoH
2MOr0qO5qyf0GzAlAWkvoeOHvEJtiL4lYVlKrv7G+uKm0ZkTPy6/Shn7ZQnj9B5L
eODW9OVyM+UxtiXLanwVgJVFT5uLIQODDVfjrtbudHi902Zra+x97ui3XDwLCAFk
YkapPQbZlNVn3o2f/rNesBaAmqyytRgWY0EiX/0efJcSTEDxaIL2Z1CUcz9J7G13
8h03EjrPj1WXbxFL9xVaXSb+q2LDdmT8E9t0q8sa3H1qpjNx0gj6lHar3cyfo+wA
oTxNe7PuT1mTl87sX89VFcaGTIgtfAtDeHTJG8/KqG/nU8McfvwhhN7puqRdeHb2
nIywF4fV/UFUbbbBR/k/ZuXBmNqAf/FoBvGWI0wEYnDzfjNZaqYibuifk5YtmITF
Qxa+ozCJEzK7KymWZsgeItF0Bgepcu9Z2L2Qos0L5BwiBbVUCBkIuYBrTPs6SAI8
gFM0kEtNDAZ7jnKyRO9rOXbZoBTYmnJigClALBRqgFJGgjE03jq+7bNWjhbCaQNa
pPymsArwFRhJna7TH1dTxCRWXYyDDhEIMdb+ztvAEEWEfACiGXJ9k4BJfzPoaQvS
C8BQWhWvp4On5pBXgJ9Va02q01baKVJZXVixkIT0OYEMj7uTqzpV7XNDW1GhAAm6
pAH3KgkX63peutDQ202lObQG8cDogXxGMNV9TA/yfpupJ4k8gLX/urHn9ThTZGzx
XMJSD3lP64kdchnUpGuolK9NZR5wRI72XAWHLQ8Scyqpi1eYg+Bf4Zs2qK77aaBp
aoekM0kF56UxL6ocmlrEO47P8qzspZqKVYuG/F7aP25vpLsnywp/We6K50E7f6L0
/spIqshcfMzWkQrJ1myHsJPGAZIk9wygMWIeVQ15yHR3S4y608PCnBPibShSbUc6
JvIbP+0ZufoQ8zN1lOxMNbnbMxgJCzmjLf2gWTsEMy3qpuWgA0wQULH55ZebVd3T
VHaDucKdvL+5PtFFEZeMv45B2GCe3HkEKSfzLZD8jVwi8ZKgIK1OPt7qaiM/0/qo
64DC2iJq4tVLtRWgF08OXFv7XhCP7ftiibqKVprljT5rSJNzGjisKSMg39q0lXWI
kGsbPCRfU+XCfCWXupoaixapuq7Of1/ry0NekLKCumz4r+Qpy6VUv7ghsJRbc9hX
AOFZjGFXU4mb9Y/Aa+UfvqQk1VA/m9Iku7JGLdNDWkG52I2M6RQ+xUwxgGvUaUWS
59KcB8K21eRfAwYq6mwfpU/QJaIwrsfTcRbWpcszoQDPTdhzDpyX5GSY2L+bdYHF
ATORwXI07ZDK8IvCqxQukDwrytYtbKrvoD11DrVZWc2fjW8OYIiosYhmealRyBak
m6+UJJBNVu+2rJMUbUCaA4X7uIyQnhZ+FKfjzPC64Jz3UgbAokWpTYy9IqmxP17k
60jjfjgNTU5inbN5bP/rGeyg7sPUnO6tf1d0OmO5laY5gZ/h+HOErk0CBsmrL3V1
Qg/ZXrM/tCzV+vpMiRci/rEilTjWUUS+XlARjCMW5rRycI0QPVYQ4guIDQx7zhRz
sqYB4Ll9zOclUTj65/GCtPujnl3l4qkIsORQ6IN0w49LhKfa8ivEybHoxDNHaC5E
WPRBCxqZ3rPIIssbaXMVyLJAQeYm8XeDt7qXqHUlNLIrM3VCHm5nDIlXlGxQQ7Bl
+pXAwW2etGy2wbtkpxFQNScSyPb1aPUFjN6NIpbUzG84QRCP9YJLRpnlDTMNPR7h
tl2IGu/cguSmUStdZ79SylgjcmckqWzdrAYIuoN3SuxOShyi5Ip0HU3pyLQMn6Ja
aOUn5tgNvxQlpxX0LabMNAZjHPih8QJH1YMTPvMJwj8zHoEjWs1sYnD+nps4VXSw
C0cb+qkeW+0T1UpkWV1fPoVNQtjNGdjYPbkhf69kx2hMhwg1Bh5V+z02SJVmmjFi
oXN6mSkFHNO0Mr2mJj0iQzPn8Onr6882hof3MRhhpzzfn3ULvdE5OFRe8O/vA9v+
y/Ez9hnl2rdl0d6JTOCc6yW2B2uqqUGQ8Zc++nk0fFZxkaLtG+6C21MRKnudxzwr
hlFiuC9xbKYMgvfSw30iXCRPSPDCruqKzTfgfjzG32eTDC/Y18+IVqwe4mLwA6pR
a/zWT7Ze912UoDmHa2cVpwPspb49H277RlbLKfYgpftGL2hXwYiHsX7kx+KmxHvN
iH302ZQAeODQbXjkcaE/XrexF/PZSXLoB25DEOVigIbvgsCk/19UT3w9mObtwiR0
UOb9S+vcxmGbVJ7Lre+jVF+KQFe8Qy6D7o9qDV/ry305WNYBvXXxw5r9sOUlUcru
RJ3oIiYm72isJXaTY3fb8wA3lHOVygpF7ogYmcZngJJ2bMU7wmvTflCEDjfpZUiI
mTkzKJGd0rpMhf+3WQlfzi63eWsI052BarxQVT0ut7z7T/aahoMsTS//ALchTbuW
Vsr2510rI7aU3hkNdtrRW4x9DCf2YBIfzxLFHy1A+xSlMkbB/y0OXwepiaj3Nj78
G7Pj/SIFDdKSqlfMT9jV5MoUECyfYWf7Gl3PQ+nS4HB4FEhc42LL9okY7qWlOB5j
B2BesmMoUEgnBCbW/C8dn/c4RHgQ68/t2WjZjsqxzMvLaOU3Xe2l6tRCcx8Wsty7
hECJpYNj26w9paWSp9qu4yFVYeZk+mo0bR9heDgxkz6qJUnfNnIAw8MrCMhHbya3
hjabVjZTgZQ2tZuI9/5EiC6cPVHdXxSoqBrk7S6Ql4uCe7kHtgKsds+aqC2CYKmZ
n/Np8BG4zDj4UgtHxTGkfxdPgjnAkTJAaGloR19dJDiJ+FnWkhjZ+/ILGlWlez9v
kkG7/eKIfZb+/tYajDyBU7pjTd1bcyXYoGs98N/qkynx9Mr8oTYRpfLg2MXYu3eE
y3dlivQQA2pCnjkZ1D5VSqEILKbfwJhfoNfPqHHWySWldqCcTS4qt34q15KK7Y3v
7kFhbysbZcE7FM067jqGGqmesSDitqM0cUxo4uW2/nEkYgPtjz7dQKrL7tojx1EQ
C+ApcWVlu2Vc9FqKeRbb5uln4+h9Vs8nQM2zqwjzhUkkXGhl3khR8OEfwSkJeMBD
XlKT6R/kN7eC6Ug7X1oDO52f4BoSk4wnJN/dF/xMehkixKITTr8HqlSAQdaJsqMf
XnrMR5Qo52mHhECEyzU4/qYfTVoIxBTdAonS98RxHvJXr+G9Fb42xddJ930SyqUS
0R7e7yF2T0UOTfmq7Ix/n9w7NdUBL1qEujC+lGh0ObK0Hcr0ZYOLP/qFFNMcskL8
L2K6N95JJtTwvkpE0zHqaByFR9ubEl20c1BCwIWI51Sif/bTJNohS8UO/DYyvPeh
LPCi1FqfV3Lgcpd37hXMN8gVglT1eL3bE08oYzwoTp39KJ/9IsWDQKOa5TopuUXn
YsBz4oPhItR9KfhTnrhppRSWpJlx9AnFnZdQt7Py3NZEoLCfZhfmLQ11Qfjg2b7K
71z2Kokd9QW/qd0EhIP/6hETI4EZfVPtRTUxYlaNn58LA15vppXEKweuKBcFrTz7
0gFcOJuXbTIKJK/WtQtgsZ4/bS/a3blIyaNDWQvFpIbK4ZXb590i1ysZIksqmuak
z4XsOLS+EqN1FniNwdHTdO29xo9zDMzn66f9sFKPDInpsO6USD+o77Fa3UCJWYZv
mvA02IuNKIVnTW56vUiBBS5d+l7rFPcgm7owvIrEicDJ5ra8T1lAU7gsnVsg+EAX
b6iQzCpwx0N7HIWOc/mLY39koOKwZhIm8prkEhhxYYrHorQ5F9o0zWF2ppHV7mOz
n/PUMQCnHmYDkv6tKvvx82GsitMLuqtCxN3MGaNRMcEKiMgZZvFVPVelGXNCaGoW
uyhaQv+Z7eu1HFKeBTqaZaazMMoI49Ylp+WqiEpr20Q4oaVlYukVp90LSZkZ5es3
7R/Y6WxZVDnnS0K67RF7pEZ+biAgm/1tMXYHb7yAsLNtNGcX6JV53HWfee1NVCO2
kYpWKWCwdjqKq60A10YkA6nVKa4CF/g0WWLe6rMhxMOEHH5YoqLEMPxP8ymZrfuc
l7hrje60LwIvjs65/ZGCh2oglq9JMWt/Y3gFv5ttlfmbAG5UFfQBtVaqeGfFtQt6
NuTxRu35/k/b87gCOg5tg1oC4N+bzzTzZzjuEespoZD94H8L/taEtBVgKgb7jrhL
tbaHgMh3wZxFKv4pzfCoNHCYn3Mg+tOxf4nDxEf7wQqOWN9xOH6dmH8i1DemPxCM
4K9Xt6MHq6cgFl6Bw4CR17q7bLO4aY7qLRJxpM6u3Dol0WINl9eFhrbUyO3ZEPeX
sBnsvEnAVryiGk599k/NEZ8222AeHmQq3G0LyNj+UkKTYsgMy/fxEUpsg30wHliT
3I6KDd7hpOlpfoRXsb0O/iuKfyee7z1GVvQQ3hYha3MK5ZplOEi2F+jugp5vPjLN
TqpqA4E2sk6QVI7jgfBeqP7f1UXiPlFPYoyfoACU367k7IeZhXvPhuybgJX8IwmI
peHOOKzDdYmDb+cM08P66N3V1Eh/liWPAe58sGQqDEsjHgqIOlXg6ymHMJT4Jm6X
bTNYDGqP1oUO902zh8bPY0flA5JE6cTRL81cdWT0GnRiNQn3OGSiI4zPQYuG9Nl7
r9amegCp2N43/6q+c3X/amGByB3Zji3PD6OCpEwuRsKDycniEPrWb5FVwFrsNk8J
rrsDpHKuZKXZvKFaIJJCRAbUnkgNJvXpinXkeDJLgB4jxOuqI5hDm/jG1PpRCiH9
eQgdLkRjJ6R/Haqi7c13PBuDxYdYdi/f1O/6+ZB3mTGNIa23orTFHkWVM6Zlxv0A
f80K8/3CAWUvuVMliM0UQIaP3iQfayCY0N8ULYqF5uFyMpqtKjXBOuvFkVkF2FlN
28BydOsYy6b4OIfQsLAA8iWaa/IhuVFLO2qT4buoaueOU1arXwLB1WeVojF8IVeX
vWRNNenVgfT2z2cQLzDLBmmD32pkxsvvjJli/oXu+c8Lq8SUAIKtBvSVduhoNTtN
lTx71miOIOwIanJ5hHmKwk5VDj3Rs2Rq284BmJ0UwlqTp3cIbh8YYsgVQkZdKeje
q1GkK2uL5lUiDvi2fU6+BCE3xZnb+7bkzFzkmLqMsmvJuO/MQ5yuNkvlVD9YSm0K
6Mqp4/l5i+c7CL9G9ieuwJfEnuo0rV5xMRXdsyQs57ojljHhgOTlNoYTX89mQLtC
QyA5rh02egGTqEF7I0+EqKOwNt8SzQu/qy9ZJNh0u3JjNhYW9oksCN16QQSiJeNU
lAPIGKX7IwKk/cpRA30e2mRzBb4cShMr049fmdsuEsuEkPOnBt4mW3IY2rQ3AU7p
uYo+teq5c+55vuDTI2ZcLAT1itM8dvZ8DH9NgWYSph89TdvSJXQnJNhhCOU30LPA
2geENjdQbndfk2HIlEk6iesvRpUZBXLrfpCH6qJmGppyN+zdggrCa8MRondBp/sW
KfcHuipQkMwRpMJLiNaER0ENMAYdp2KsSNqTiMvUunvz2/VijbaGzT/8YGc8fOxl
xy3OPsmb4ikufksRnIYyau+dQv9ntkdl9ByI6zlIRKMoIzV/EnpV4H/GP2vkGjCT
WTS3P571pOE4nk6pKjMFCXUA7XeILimGgRfhMFgQyir2e5rac/tDNSqztWzmEBzu
lPWOaGgImWNayrVFPEjEQIszivkvj1Yuwm2hza/LbfzfhJx10kf5/WJbyoL9/26V
CSmbfTTarVUM8USlJkOCzyB9MX+MfqMrhqQXwHy6taixNFSYXCvyNfDZXsrQ8UQK
htZqxorphbUScNHRtXD9lT6hPGphIM7kBJnYleJrNZrB2EHKAahDTzLMzNXrWS9p
C/NqkKar+1LDpli95KGsJ6mYB0YGPoLQDgsqzCQDpTrC6a8OfqtiQpqgkcPJtUNp
EmxGIpy5Hr9N79wf2PW7eCyoPTPLxjMarcZhn784TXJ1qUY27+jOBylAgTTdeqIP
NJ23dpxQiPa0kJYakNrf6aqCzaWTFyj58rWlThcbItLAnWTOo4oCvOPvuSJsbdIh
7v9CgktNP1A8vvb5QWzzI/ZcCElBEKvKztlQH+pTkCROSeGKe/oWvwKeUZu86l3I
vRkm7t2V+WNbRK5JjDIY925tvC0GlPaAJOvEQU0KxcwUhofB20HJBgG8pL1U+cKw
35FFT49UXtJb54onGMs2SAVY00dqIE/Se5dASalRi4yQ3XUnO4A3sdFo/Egapnmf
GtuV/aK9NjUxKDWRcZGBorW6iiFBn8J6TfDZZCUNMHJn5sslDXu8fwUq24+JWagx
4S2Y/ONlvYXeCYpnVyiLdRiTt5Z+VsqIz+Q20zlui5ZFyBPdzR8H035YF1itq3te
4fykoAPy0N9mb2XbMcQjXe6Cpl6OUrhCeyBh7nts6vUrtBkXTjTWaUYJjgZ0mpIo
XTydp90x0/PE2tE0sNRfI0EFlQYlvhivySX7RvfgRfJHGjlS8BGkiLATdno8j7HV
XfbdUq4wW/ARnlhislqZXyLj+1k/cp+e+dgZxmc8l6AI+VXCQhWMwo7fHY2v2Gp2
vDX5DbH1curY+De1ku+p0TbBxu7uhRnXP4WhR3qGOoqBQCn/1j3Vv0EYR+On1i2d
gS8KuyVnHzyrBfCNxJ95IXn8jBpYWeAaxm9Oesk24/tJQfGW51985pOo/p8Y3Guu
HxBhO34nNEE0fZjmloXx4/dq/727QfMMHCG8dfWZXLcZyuFZLO6Q0PwGukP1kCVY
q5gDlFMw3W06Ef8Gpl6/Gt3CZbRUE8nRKABDIOPPXVvlkY+3prr+8BHPAGeu0MBu
W3GPww4Qn4f+TiyCVNh3cCScnV6uFjowYJoR/kz7l/tLSTN0mXdEFPgJA6GOe7J4
f5lO0Qk4XtJKIYIR+HBJR1k6pqxzBK8t7LCYn1ZSnQUlOMpYOhc5ffXhoxsiDEZ+
P7XzvA67lGzLldwz3AWy74uZ8czUYtDXKdMhc9G/wMP4mH32dxUdoj4NhcBaos5w
drCYb+7E2/irxQHg+dU4yfHsUn2hokY4II2AdMxTSjzpL3d0bckcey7hbU29kiAg
rETcBLXI6S6OPF0JU69jwFf8dP2kjsMZPzTgtc12VERTrT+zhR+GghcjsYc6Y6X+
WmHljxcA2S0pvdicc75+2LVCneJAuF278njpVhNHc/v2j/Ck0HpIBruKbCFJANXa
Ob+7RL/jx/mF5ns2xkwNSBTlZHK0pLxF6TCRqUta7MecNH6FQ5sMtD3y3GNYEQCW
A6KHWnILXVLuiv+onVrFRnkrcWecy2U1GgLV93qdb+zsGqImy8L0DVQQjcVIKwqk
NUhoMh6mEzKuC/EZZ0iuCMUYY+N+BwR3rsXZ4N+S7SqXgNNMAEPkAeFMZpDs6dGj
SQbssfcjXIdTFSNzm36bLQ02KQ1ObDo+nz7wchhSRgGZOrq6Vs3XILDME6Uwo5cQ
X/T4WG3EUT8JbpVBQBt8ccDgC5UOgJxwW3/sHLwuFUfcZFqbE+jS66xGjVSE4sWD
/qGxhT+Vphuo20yhmM3p1ic0NbZVYNETktK9+gebHRf0zlu4bVKtjoERUiScc3jg
zJ3iO8GfithdxN/ti4ysVAwvrisZVvGzWIpYgY8a9/8mWlpdSZXv0CWQ/Tu6OJv5
zJxQcqEz9Qshpyi83KwLUnBJhsmgzX+GxDiEVgLBuOZHtUFg6xxiGkiVGvd0lNgA
zDcotJ4NJ4LdmBeozrGTqU/bNbBjNfj5H9uNQs6tgD7mEBXB/eQ7wW1BsLVitrRt
NmxkNj3jqs4vIRSMUCTRqorfUgpFGutZnSBc88KAuyyX7IHK5lDGbup2gAi/agDt
nO3gP5ojNn0Y+tS4uKr31xa31gas37hnbNZturHYWsF40klzmout+Mzsm+gIUzuL
OSLFoIKPoA/RKZ+QkWXDslE79E70g17SfsbuntWWGpadpwswHbHiYYdPO6SY28dV
a5eTRwybQQ3yW6/ZcEnQvxMJjRz6489mA1t/N97ktSCjQk54a4fF5jERgBY5NNDr
sTdPyryIlHEuZGJgFQi8t7LK3kMN5NjVQN6JavHWYWVRxmJ+DoxnFmZmrKFWGnMe
lq4mbtFw+MLjJyhVW/C77RBRzsLhWuE6hRmAPup8HYBY7LqatVf266rF+iDg9kAG
bUvDBg7/dVb7UyZ7Z9BtQj6pa3ylUW8A0TS6oQPprN70Kri+5bYGiViTL3Gqn5Gz
ZRX3W+49XEhRvywBcZRZqotPFNwk3Fv9DIeoRxYnkxGzJMos+MxQ7KMD/g0nJkxQ
YOYDVLTj7TpWq00HGKwcv0/iuev9pXfVecHN/KOyVCAooi1lGowGLJQbWr1ZIK6l
XqKpZDJp7cqNTgZGgwmpBaDNOueEudmN6XEEsubRi5TKcRTNmOO1OpavmUFa/VoV
3ByJGtjoiw8PBJ1qi9Kt3klqcr1NZmil/AMFUHjzeNNRJI5ICl2NTkjLTIIRsvVJ
pV2DA+hNcpCV99KNtAkozkHfGj129U4iLKofqQNEuCxgWxjZ1jLF8LgZFERACBN6
mjPtAezCgM4bXz2SNd3YbHIRr6kgTJx6S98BJKgDer+8tnNNdGRgK82/PGBx01bA
6hPG4AD+/5YbJ+N9sJ9mQ5HTVlZxGqjuQvZfJ7LNcJugpMMXYrGK8GhSqH39ll7d
P+PsjDchWtKvk0Eozzy2WTpSTtiHCFHDeHtHyl8d+OEXAJ5GJBMg1hZroB+jy5Q4
TbFzKNDJvmSlDM4dMyx48E4884OGrEq80hPLaVRuhSGxGY3a0HhDoymOhutyfk/7
qAXX1teLcRcYqhW7TsN+ga33ZcNcbTGk+ajAY+vPkLxltbMCE7npljREH6+KXt04
fYrzZ6RY05d/6PTmTb2VTsTcQjmaThgAtuHqM6A9BpoXj27TwmzSyJJyGiXk1Iwc
16Bf6uD57JRKTN0YS47u+WCkx8+qRg7fyYNeF9+6xws1d9H99TaRsrsIMtQ+EVeo
QpsGe0U/1fmxfxvMFNQpTwwEX5Mf0MrTSvA5wXAY+OvW5Ihi72mBLi+Xy5IE1Qnt
UaU3WIMRLBLVkiROdLDlmsTwb0/j9lyb1liXirWJWveoqnFBoQjA3mEp6nL9sUde
DoM40hTFreega5NXexN0Hph8PHwq+3dZuNPn8gL39TtY3QeBt1+tEJobX2ouTNAW
QJpGvoZ2rYB6P7QKX1bNTtbfBGgmc2MHes2aAqJx5o0Z1CgKp+8mkPV0BF/e7yEN
8okZlcM1W9kphtk5P8hhLd0aBiNbMcTooX7BDFF8dPnG/Uw7ss/iiJp6KM5hIBV2
6wbUrQ0/fI3jGKfCPNheBopssm2Ayf6AoVDKF+ykRfMqG7ZFqyJ/yN8qkbNZTv8s
W9F4a4o9tW/VBMkr+eI6eSFIq4pH6ia8J/bHyU6fbUjFk3zmQV4g3sblSzicUrpJ
ShCdRyJHPZftr3DvFNQNXFKlcYQb3Yj/Q1m1oH8d4/O+pVC/bUnhqQfQ/E+SnPyS
Z6yTc0rzajEQQGrnDTY78Gl1tYWMj6yX1LOBsl7Scso4gmEhqtfAi+PXaEY+CB9j
VJ4TkRDH9+y5mrdg+raPuJWxzSkwfIyHxTiM4Y2UNHenCFF+fsNPerjFpe6oAbOc
LaDFOkwNAwrjJYBF2WRf5l3vtojG3EWBpvDcB5voaYTIPLZNEURj3mYOVF/V2NKq
1boIqEL5GJbh7z4iKQ82ugqEMlKr1BapI0cmTbszAI15EjZA4YcxJjkf2YNdonvm
3SMQcu0F4zuAIMBcgNNLD8nq+9q2eoEG29VV0BXxiOW82juxj4xBIFtuLYPH6Ffa
+YoeSJ5hVxkUo1nPPICR8z3ncln7chixDc0GDiJACEWgG28VC3+c+0j2zhwBsnvD
mIfDkpBvNi0mYoLpuFp58bys7/hovasKwEYlxaty/7wpQNyzvm7dgEbFO/Ytde4U
DTkF1qhr/r7eYwJAwVPeGyKVA5ZOi07JMhdhtKwIepGEwoD3AbVsgqgP7n636a0B
4A1b+9U+7WXjFpLy11x34P5SwwT0N1Ky7sclUGfDC/hbZyqgfToDHIoptIDoCV36
HHc5/nGh1vf8K//bKF/cxXNWSA+RshEvpEZekN6wcLGVGtPIOGUFuMedbmtptrQS
IbBiss3iFG9sZPL0gkXr7oRQRvWyRGJeTir78SlvWROtHY/0lgAOZnPrRXfbHF37
ShPxvRsz6sQkZS6oyLJoMfA66q4m4uopQyah6ySQkw8jArR/IGZmFr1EvKX6y8hV
A+/XOUI3Y/zOlZvjyDvaw/Zgeze1FclSsJ7XrfcLZdX1k+Hfab49kzThR8eJ+VOo
6+uMEdc4XzYCPR6nRmhyXRuKJF2yk5ASUWln2aYKkFhAfSZ/RLdixzjkxzUNvneC
GX/8StApwCBcU9JQ54nC/XQxRwKyJFNmwmtNixuLkNhYRNw4MjISonWbYILsBvyt
+86YbK90ycm50L3pFnStv08h/VVsMTvVlAKvkAJvepITEWRYG8epN/+9nnDwEVgX
ON9E1sFGVoOpJH0WZa9pDJy32mJuaxfJsZLDHmD1lolCP9tTlf9Yjmtqmkn00R5g
80N8cUZjBXyka1lGrVczrPgkGHvZOS9mKEhTk0zbgqitB6UHhLWIgKTiokiRijbh
4ous6T6+i+ZkBE0IgG84McqIlIHTAhZCd1psl2rwzjdD51DAddJo/9S9f1aCLk2C
i3oTDhPF11LFVmq8ifyRgt5NDIhNmp+D32h9gknKQqH8aHVfCoZatflXz8Mr9Mmy
JRQUuIVx6g0jfzmgSfnz/ZTnpbNAmwScnkgwG00jyff0Da3Y7MY7FMSMbJ1So0rz
+M5rNOJ0XEX2rm8ZtJsswACZ1+vBEqT4ea/g+4+9s2JiAlcm91TpCinhoomcwW2Z
CMpnDWqqg17Q71r5OySj9iu5SzSmPVKozwvgdcHTCiytTyNo5lrP1hbm5EXksrO1
WGo7LXP7oLro+D9W8JdKayNMu2C6mwUjFAg03XGFe/8AOTU3shrAVHP2sAGT6/TL
bm4jvUidog3L983PkA9hsN46NVDdL5r+6Hta2J4YrSxTthXyln+Imhgekz3rRnpI
+PU26w39iSPVhqX5xy8RrdZ7wKSdKmkuhK3kSQuGAWFczASQzsTSVI6OXCXGhPHI
ArWS0SonG7PWvYTgPyNmtzk78Vu38Y3JZGfIn5l+D/e1VrSQffruAnoP+PIfH0FT
iXojuA+oHepKClMqpzeNGrYr+dIEkLRDdXWePCO+O2xWzKb+KxxH/eklxnIRMjqs
UeEEauR5mn2p09zeTCOPFmvhxlYgQ5v+ZwiV3RgsNrxasy/Bj99vyRE+N9nmhium
OgLr4UFtj4mLKmoSCSBLH3NmuXzEVEi0LHqAMCBbHI8Mn9+1dBhCe5+fo9Ol3cCV
4nee9hZKK6nKhHsztyCl01kYCyZA+hZHhqhtczAhCX4IPQRRlhRxzC3B8JrYsP4e
LwVEUrdsjUE/ukZzWpef6Q+PwQFQNzc7scMPH0IUwpz0w5meE1FyO1OYf2NFBVY7
JS00nAMW8cIe+wehzY6gxInugxaBiKdjlMlc9y8pEdjEeVSpjQ1HyYwzglWJFXVB
MHruXlfaaShWcBEtTjAafAARdq51BBT9ue6nrZIYduGZ7AQ7HvETHCdzw4wy5195
jBu0fhatvblQv9T9h62BVgXxT5zh8IgxdTvFA2MUVNI/SqpOlrgAnq//iSPIjTZm
q8liUE2x9781olG9ZAY1r/xDd6XMyciXGWQ8B3YcAZVbO1KyYiXHp0yVRcDwqtaJ
ELa1HLVpy6PdriGL/jzCkpSxaBLndncbypgpneXvYRfvUYjofQY/beIvKl81RcCC
YnfQMydtZ63nuIH4d91g01SjIj7WFv1EA5ucpjOFpew4365xDA9ERXZPfV/xlXwy
YIJ1YEhGM986B5dJ/On9YEpC8yZ0jGsEb3LfQ0HGqb6CfwirL2UIMGDSwz5NnGR4
N1U+G3mJwFyQPllZ261xM09EOfW6iEU/ZUfnVmfbCfvgZDoJyHWNZmGRdSWXzb+r
x+sq4nuDJNY8EjlOyMEkfcyXnknYZCjNh6F7E2DxUZJOxvxlkkIriWtaj8EBzZL2
yhhs3ueOSr1PhOinGaGDfkBCuymw3WDTmoKCxT/S0LT/X7U/RFqtGG1/P5nO3Lwy
trP95KwTeCXBopoTuKEfOqq4YQiAki7GjAnG+PklMRL0p9OzI5fnaAmvwvHjuySY
A3krqB7BpMizQrBcqt5H7YnJSJVB2wKvsmEJDJD28b3GFYc7BrG7UQmCHVvw0HXD
ozfHcPJs2nCvuplGcG6utuJGUs8DNHEmAezL/GZGkttEnUIx7i1Xu7rluLhCoW5R
cmjLd1RO073wy86+Ise4FgcPdsVfg08/+zzTE1ZztmlMR97dLug/g0WsTukIs37K
HCiIUkfBIDCgjfan9B6qB29Y3mqV8qoiuh756Pvf6fZRFiWz9n9KJHNsIGB7giKE
GK4lFrIEQiM0eH3Rbhc8qBorQ/a8EGjG6tS5pnWKknfqFPb/tK171tvk8LvELgkq
EJ3REaUu8QsxaPocHUlwiYonOV7dqwn0IiNpiQ6BodDdAvp6XZxji794WincbFTV
i5raZTzfCZehIjdaz1KspqFAIyU09mxFejkM3bCJrZR3fkp7PNyWO3WR1mjV0sNf
Q9RGXfU/PmKNMNSTn9BCENNfIhAKZtjuElaurl2QQeQvbkQDNKcJ1t6lDMh1nUnX
OybgztJwcZMwGxVCDyPaWQ9/wT9XXiq85tDduyy2eHEr6qlBanCOJeEtUbD6frp7
xXt8gvwX0yeUGnpFZqoSDSSmQPQMupOUHlD9G5W5/P1rCbq0s8FznDlkBZe9Q7j0
Nk2u37V3JJs/dWp1WpmPFYm9mL7lFzRXySjRdiBnug3tXWu/nXxJrLiiqNL758CY
mwayOMeh3uaPj9LPXIah7tWK76PwHloys0Dv5lM14XdTIjlCupphjja18GykClIu
YN7C0gDWdBL7WSm66hud7xSNPucte6SfcpLqHBRC6yYKR1CDnpYb2oTEQaHE8gKm
3cWobQiyz9XDB4tUsEnk557in2NG5c135PD8odIRuA+0Q94vW/6JNagDAwHK2VWc
D0TBVV+OZyLmMHllxittTErb26ibG00ViWosjPjOVQHfdRF03EJxUem29+Z3ReoQ
1uhcrvDVGV89D2O3KjVkIZvTjVwslEaScFsZ8SUiByLti41vR6kmi/+qgagNwxeD
Gpj8zesDKaRksO5HpmYj6DXFHgtpXNLU4ZeenEM8Q8cdKbp0Zm9kvbsq5yKOSeOm
wdLKMv6DAM5J/RfbDCPP9fXpC022CRbt4aiEKKWGBcMx1sJDk4w2UD3F9Ly03p6D
u6ewH/nZSPhAfgmmLFUlPNRdrHFrwH8RJdSOU9p15tt1I4yW8sX0LhASB2CHwATC
eWiZXVLroPB22yO3mjH7NomAC63/ih2kIsSmEpGtmvu90UCMhJ3gaiMp7KiKiVaE
FK4f7x6tGKlNATFR/R4xKQb9xXFTzWHtizu+HNLP3l5nMvurEoQGp+9GdU3o5oUm
mpZD3H8v1B3PUIJdreuKLsXu4uo/ZpTkf2MDAvrbQJdHzoKZtue9jLaOv20X5ZVs
/lNZPMBgWkovkhMu+pXkQqMDW4S17NUBJYT0tX9Y9kcVuvRdsLHSUiVWAl28MA/h
nc6h9cwOOJSG9rk0zfyW9jedG3ZsD5Karysh1K1n1ZJfRB6GARB+KBDKkv7OM8uJ
iR4WhnDRhtXp38+3jJvZSwOVw8BPXBbtRnrIvuTIz81pZyVQl0zTlkhQJJLcSEYv
zIqWps4BaHOd98N9tZX/AZJfkGVXbXsN3gc5hzV3K1L1kp73l8mTnRNoO+P/0DjI
levZksoCLeRmI62zngEhKiVnUtiPIJVvYELOonyWuQz/GBOUedourLcP0QilGlZp
wapIdtKgtSo2cc+y94hoUMkeYoY6xa9kfpe4BlZEq+QefE0DC7mMejgKSX91pcCH
JNpxBPfhPTY63TB56PcZtO0jI7PmZbjelLe59CRg7ZD23Ont/hVkDl/06g962S2p
lcp9H8w6Ynhi/vJEA7cUhEZCUbmaW1JHB6ZzpsXN7cUxqYin1REOcJq70kmNDEoV
/S5ELrc8gKEZnhl1KVoF+9wwnzixk0Hu4w4PtbrzWtr7fu/jl6g0PvxNcPXWuoMY
1cuYj0eA223NVLpQ4UZIft7j/oIVTWYt2YTNCkTyvv7wzXE9gnFaR6KwJIhhnrN5
jkBF6144sUFtNsjDwqvzT7n/lW04NqP6BbYxwJz8jRuuLYXSoMWMvQUY1SwQg5uC
nywsS8AL+2AHuIFHXPjYcQ3AIhDUMIzgxS0IqGWS3s6hGzkkuApW8rHGYt5buKU5
J5sf1bKMTOg/GOusfc/2MgKRTUv4jr+vyUKcp9M6YH/ifh+MfdHGQ0+iOaX9P+ok
MwhPbu3y4SFx03ZFNJVLXB0kpyecKxqCfd3bETJTeOAFOTELVM6i7S7o6JVbPSlU
8Pchi+0dKvlSeoYg3BcB0G19d8/8xoOcSxHcCZ2hx90sVNkEpt7iMZG3zRt7ZeY3
uk/KpPiw4r8BcAI1GBb0YUHM+cNTbEsv645Yc0uopaDX6l+YEyOpGcV4dVQa5WXf
ajIGK1tbQiwmj0USQv05mxAzaDk4KmepWploNJ+OZIZhqvIevl/UOSZj6By3dizm
76J3gx8HUDVNXkqV60YGkzSftYTSq//j9LxycjlGwj12YCfmRqv3621iP94Pgoep
Pzy0pbcY0kVYRTGcXFc+VXkSmHtuHmUU40T0k1Y82ntNqNdX0EjTDPCRkM8eETrU
5NjMMWIoBx/2lzIU7NNBELp5Wxc+1avpvTsgwqi+YMiIzL37ZAhdgvJwgTSeF3hE
iF+rQwKvzQHwOijikKWQbOs1muleJ2A1qkZeQD4uyi/Sog5soqja3hy57cFCY6oY
FPH5rNiAl1W1uLebNYND5JFTzvv84Mheq6EMylg232y6CxzMh973afL5irECWQYb
EFKjgppI+usyN7FXNN/kRt90d3vh2NidWQ/f7leHYNJuv9Brte6QuEc21cmQwC8u
YeK+PqlaS96fT6ppjn3FHDACF5V1MmFGKT3BFPcIEtnGFBwVVCrAtfmTMIK6g0l7
VfCO8fH0j64XYBoy6DsYGagBaqpaeCGaWXo+WVUUJmOmoQnEvt6FwdGse5QC4SdK
UDnjW87vmtIaZishKh1pyOP32qz4DtuQJv6idqZ/OttNSbHDwMS1Yru2C26X6xeP
NcPOznnsgTrQQPYOBH0VQ33xAUFAwfrLX4DYsB3ZgzSiYNqCEFjy8wuvN0nSUGZL
oZqGAmIA8dSve/Aufnb925KkMMeb8v1ShvGjxdv7N2czjM5MPVcj2Io3ObpVPjmm
APoyC7nQT4BJNzIp5JX6G+HDn/EI4JWXYNjEI6pfkCijk4SkT19RT32dQPa8kAnm
nz65laPE0NE0lln1tiOn65bB46fhBqPP8xGIdE4U+7H3q2/xY7HLkBE0V+eCTsNN
BA7VpSh1VKjRXbwT2cWNV3q5f84DUdnVKIr681+YqdRbQemhC1uGYgy7GZa/gd/u
Wz+r5VbEtINKA/aLnfxw0D+FJV2RF24HShP9XuXgJctIr0qRDwNXvR5lOYGY+bzd
iHFxX9ib9txkKMUneQZQEVBDysOElRzIxG3Q7d+uF3RBRPDJpJ0XAivJ7yw0U+oa
SLTDqkp7W+1ca8PlYl3gd0D5b3Z6zrCHod+oid3QXu67wDiuGCtkKMwmPiRHys9c
rBIga4IwF2u/f2/Wv/3UUPhAj0gYlM/Q/eOsPIcUr3Qta/2EDYOeNK5geuuVUXsX
hG7PDS041Jh7ZFJPszWeS8tw6zeRaGh4QTvucX2JCjJj+CxXsgbWhj/g0Fs+39QG
1mb1E2Jt8cjkTJsXyglUtcLXjgb7ozwbxFByjCI3IfAyY7UCvfvc2kQjvzVfMVO1
9kBpCx92rEofndu+8dRUXQwpZMg7+JH7YR6uRgi7RySHlT5cpqkwLks8OnjtZZSe
y2EFUwYrNiipqJRc36c2gsLT+3Bds63Np7mJH+vUYMI=
`pragma protect end_protected
