// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:02:17 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
DLoEGZOHnP/PQic4yn3/nDL634Z1EM1gOAdLnYP8/sX1tCw7JqgEtxM1/4Xmz106
7PmNCZBqo3FhHeH447kIUt3q3SNtGV0ksmVSuJBanqQRYUHBh1BpxANh6LEeTrM3
8jwZzx1XNE0ORv0hbGdHP7K6Qw29+Aw4gSthwMxb9EE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8480)
yQ/KGPl4Yxr9t8X5KuSHh8Vjnds18s7a3jm461fnkv16Qn4OZMqrsuKCDn7ejPKE
klnrP08BSFZW0hJdnk+CCxJpW/nkSuChwjYDmuJFvKpgRp/zZ9vqy42YuMQkzMM1
23rMtjCs/wkS9yQhFnxqaWpx+OzbV2RecRtKDFRlFVO7SpMCtkS0tkkGwyLDk54j
Yas7ZSTbDTlU+QOy+Amre9IVOSqPXd66YfuvIeWdJIlbjqb/qniBSSAInKwSf7SE
qy7GUhE8BPtc++8iXODVeJm6xVgJ4zzmR4Q7OTtqreEzafkpmAMkKDldD74sFOJo
gluuDqtN5xgt+Ely9HfAeZUsdLj5WnJrtYMxWtP0j4WLt84FAdjg2IodhfHq1zso
KHVw2NSkK87WJVj3SP5q76VHfg2kaIt5vWTrR+G9P6QQS27Agtj6b++ymmXuMqtC
FBNK78eoS75qbFQVa1JuZ9RJgHfhh9jwIlf4vEDP1NsGw2qL5MQxyXfERFkCi8fA
sMyUMlu9H+DRDJ9yW8ZS4IyzyqmRc31vcsAPkVU/E9gnjYxinMkozVB+h5QM5/AV
IoT8x4UqH8cNa1Q8iAcPQz00x+pUdQrkweN6HxziOwzoQeqqDvUy04RiHHe8DP4o
kpC3v75mzCRk2hYO7maY3LaJpB7puc2/oqoIAlQlOHcA/5W9y2B+9ISVA8Tjqn7y
gJEHphPpQXD4IFAzBHYbYIkfnIZr4ScRHmVTYpZztRgtFF7t1F5lGwdVdZMEkNJk
HpK1todP4Z1zL91aZjTbB2dnmhEFkYQufeOdOgEjQTTq3Li6mXv4KPY4ZwIayxpN
E9HDcADQ6Wknqe9l4t0/1ecZM4wU2G6opcA44CNmbmGp/4BhdWs454IGKZwRK9L1
Om+1zKn+qTCOBZqXSVU/rxrqYsjkagSsZG43rUrBTPP/oT2d/dZiSQo0XvzDqq2e
MdqKKA0BLaOF2CHtQEH2hZOe9/h8LFcza330ewXsw3EzIe3llIcTaL0TOr7XK91n
A07qUW/Givmw4jtRceliOtEGKc/ZUU9e6NY4vZdfagY1Gl/iOIXelXyRk7kqM/XX
LmHQ9JOtyuEiA3Zra90q5QGOVRJb3GrdCl56gbnVAgzssB6v8CYgiUq8rp/wx55K
saPujp8fH/LlJVlfgv1lM9H4+OKtOwhVwyoxZxosT/p3j0r06GvnzZPMv5KB2wAv
7VuoxSV/yuJEEBYu9GF1xo4sYHTsO2D/xhVyLwPv6+GVN+OnfupBCbJIJOIQb9sv
3Vfx1eoQwbILNYVg/+1OJ6oBHA4e8lh1RW4QWfHD6jy8f7HM3SyMNVxcno4pR+s3
Xitio2GvcXc2EUdfqG1xj0AkzaR5vfGkWBga82RjlPHL5bqwViedmnfZIumKmSVb
0eHg3/IoWILcmEdh6Zj9FzhDBgf/jajzA8g0JMK8/M0ODxbz73mCtf5U+LjPoQ5o
buJpalOQjUr1coiBjeoy0mnYioT8codSvFmFGGnJwe/17O1kFF3UT8RDzrkK0aLp
xIPDgHVT6D+KhfkGLulf8iLyL5LZescOJmmN1E9Z0fCNR6Wzv3raMWYYQqLftWwf
dQhtFBPYn7/Qvr+BH94d6XpinsgCW0scRgGHLM3svdodBv/7ZwrIxmi/IvTw6LI5
rZSI3KLkXtPoV4Ej0mgViHAGlxx+brvQNQVjcbHsdjyWb6lzRFA59OeKd90s0zMp
2NdjCea/rouxFS3fsFbyzDB07jaONkE70ud0ngaGGCIjaIhm/LeQEWMHot7Hb79j
YMlgwre3aJDGWbCRkELqe9mjtQmc9kW9waBTd5d+v7pYAuHCwY8XVHjO1ussxzbJ
S+BVErsKyrOKvQc4Q7JtP6JMWizuqms5Fe325T5F+EqheksVvBWb2jW4P/smKigr
Lc1i+tVtsIzzfmEqjemDuoyGmI1j0Hk3opIm5El/MGPHsPlz1FcYiOu81bugIIXc
pkFAuNkqPSs6YOlWiOH+4LKV1+9rd6XNT4+labOrVO43uaM6aYz8zyHzf6LVz4gK
+VMpGen8xpEgMyI19ULYR4RIzdgfORivyyAFm8IGZoAIlhhGM2nS4i6+e5FswxUP
i/TZFHAc0U7bp+G7uogtn5YIsZe0YyP2i7zOm6RaKvVeoDSLsFdqw5M8pIXWaMu/
k2hQBsm7nFrwq95Yc9ZAXMiIIv4xiih7tU1/Q1cqdge5NRuZiJsLRwYfmshEqYwZ
NCWWbD2bSkY5CO6CKTcVlmtmvldrsgUBLazf0dK1iBhXTuJEKE0LMLWG8ig4/clK
6PRb4mv18ZWIJr2fpdvlB0kJiZZ366VXBJBEDwlULacZ2s2YJuNGpePC8aIJvw9p
fNMzpREGTvFVt96YOjjlOQvVzcIuHaOQInv1ClPeGQs8WCT7bV7ReZH7Bthcsf1F
55ZBqjBCOtmHlS3Teq9iudsvpnVECiUU9ntO67Kimwv7gyE7ps9bWg71Eo3WAkX0
r/f+HsJWHhz8nqKBDDaM+EasERP84gTP5H0zNash1jMgiVIBpR4cVtbAaOx5+o7P
KGN2hrbsfV0zQWttx5JzeRQEsnGR77l/clZfv2HOC2amA9rkj/1QnLPPrQL+zP6w
PvDYmOd+6ArSssSZfrB/6m1SiPSbZy1QAo8l8CEMov6T13qiDOXPi04AW/SZovlQ
hHMOK+5MoGM+lhV4lByjWeJEKfHFg7/5Er2OIUX1/VB0VofHYrfrh6czYqNjsUSD
q/tdZacfw2o9Tv5KF6jzSLnro3hamXJd6UePv9DzK6Y4LGFrdwr5wXlW23ZpBqZx
9loES7jeMBlDD8nETi32tWMyE12k3CPWmUaR6hXw8P6Dcf8jSzzS7VzW4VCAQ2dV
TOb10gHSapZzMNHzqDEOy4/MmZCq5hoFVXwzAaTy4zFtCRW6s8z0i59DGK7ohnhc
DVgQSAOAthXkhw3dpOHhVrj920lFRL/73Rtf/rDuB902oXUIpgr76MFmHDiOMWem
YNk+1NeFOxCQCpxiPMfn+iapvuE4B5sIYeduGxxj4oq55z/iaelA1wRFBM0taAmK
esSl8WjJYUgYTyUXGzoy9LFyPqWvnF+H5zLx2rEeQYCIUeujcpnlw14hwPN6VIKN
cLLpPzBby909w99BUEmnACAB0ILYvt/DpZnrUT+WZVfR7SSvDaqIFz0kI9GrWa3w
uCgHcY7+u08PMdgBC4bX7J57fGbyRVu2VSzUKdtBe1s4bu/LqfaR+SD3BzvCt9XN
iwU/fPeAG/r/3O+sI8A+GP1GSnrq+GIYjmFdBq6i1JHPxv+hAysG1OjkZ0jDOxID
sW3I5CeHuXlQ2fFNjMhr80dS/B0tkFDd56/g4xFdUeXcZ9htPYERpoaynJvJBMKY
iLfly+YRlfVAUWFcOSsTenYKR2n0jK3PW11uqNsA464sVU9ApcH8bRJKTVSP900j
DUthdZnAjVLayKEMd3qGzySIxu8flaV0UOrRkH4Nd0xjNwA1IguUydeZi7+kNBSy
/hQv6sC3t6wPLom++QUHLwxS4V8btm3g1tp8Atay6/NvNnmHDODkhPzAuG6EJIZ5
Ebw2Ln6Cli2rG5Sz5lyivmHN82hlFIkeg65fYTk+pqAJ/uNNcAto1bRRRydtiDi0
dpGpiud4/Y9+JWEKO+keAkj8pDl2hla/XQeH+8+aoKQk1K55WUKxugKOMtWxzw/h
nfHAl+gnUE78XBBA28eiKmT4rpfDiGGPMglfRGShmvqX4JLmYh0BN9wj/qe7cQFK
CibmUISkUYF0VSZZCW1WCH7lQLwX0P1+9TVYrhiNvH1i5DZourv9HK8iiyZa8/NL
nH2pSQAEIyrccVF4/3VnPEfvnt2d2YIVEChAClZP5QtRpopW2yhM2phUo/qj5urx
kx2BwboU5UlVdV0dr2ib54p7QQq2pwFyeM7hPBMvl2H6n5q0O8EYibXZeliXwjBV
5O4OV8DZtcIvVlTfGEZkVa+RLoNgNSh1TVwZRmAExtIetvHEDAxYy/OtHFVuWAb3
Y26D7MaWrc4eCnQInrk9VwEDRqT5whdMLmBKMX7ToR/294rOCmVp3kfRyRNF0zjQ
FCEW2Tv8II7W9k0WQ1biCBZEAeiYpgBmPHBSfyeRLp29A2IuG+zNKO1oS+faJnUv
1m+/7MDpm6TsWhGae6Qqr9Er8IDEKshE4PoAfM720pobPIMK7QsQ3EervQ8lsPp+
Wsnm57YmthaEGB8wJbHmb1wtpOA2RHUaI9v8o3c/rehM2audW438JnQzmUk1kv48
K3prfqjKlTAnXR49qI8JOXUDWIGUY8Og2b3D3B4AZ3OakFdV1fQTmnvbRo0DMjHo
x5JUkQ4loMZjZHAxHWi+UYJqSjVpUolMQ2W+bkcSkSEEPo72HSPlqAW3qg/p7L5d
dqQnYmFc+Qnb0tih+bzqDvuUF+sGmXYGJe4fNMoAQnTT7rSB/E8X7YvEJD6j2WwM
tnAciNXrMilyUEXYgU7jCdEnmMRNJx+COvAMhh78S/nLP34J1exJkE00lFgdh4ZS
AlppcxogaTTNl3bzmtSwA+aPq3Rit3Z+LmTYpEvmUIjY5KBLEg+TYhGtogvHaHjp
EtTwXGxQjE1DFY1CNE4UUsSATF04X7S7D7FJ+pAetM5qhLCRyp5kiY7OeoR3+6TS
gbqDjNzowDz/cky1txCDX65sKMu50azAjaidZzbzuk4VvcOSe1nmMjEbQzTAu91e
7w3Vj6TZkkJ0KnQGckIX3oTxKz9wW/qJ7yBpDGaoenazkX+2hQDGtOeP6v+z4Enl
QGkCdsmdoLLUbd1PUO8h14z5ORmSpZh5I7Fjh+VFpi0F2woxR6K3UcllbRwA4p2q
4IvTiErE/sgyXQ5b1G1/rmQ9hLozuRD5Zj0fysDnOYStCvp8hyj+ezWGFPP9QlFJ
xtW3mYw9wHl+slkO/P3tibR7r70/2/FpPeJ4n+aFT02/dzMPjn2ve++mShUvWIWI
591UU8LAa2cVySBUkKMqAlhbtC895hxHdlf4LhN6WDmegfWU3mDPxVAIZ6n365G6
vFU5EXSZ/m5jqRhDGe/6A6ffZRPXJ2ShtqVJ4sPGByMzDxmU2VFZ66PmF02z++yk
k+swm1Fhiyz3WDEabFTWrt9HwNfcm2Gisvl6XOZOtUFI0S2QE0JUw5uK7fNZPgrb
vuGo85ek7KYbxpYyI0CZfIvQkrXHxk4AlP+FFa6SGfNatI+hpxXJrre1cwtHTryK
SIJu/aFzgR/OogwYI6Ia6KWKeW0ohs4K46xL5nbYQVBug98RPcXTvK+jZ2wJDwJo
e25/TbCaTRP4vx0jcQQ4mWEQsSPxNR7090Pm5ZqR2dKmyBmJc7R2Qno1JVFQieG8
NDy/RtO8GC7TuVks/nW48NmaZ58u7375lGuuD5KbLHYg4pdN9TYUy23skrMsnmZQ
MfuoCEWAO02E2rLWxTSenTGMAYrDWGebfcE5H5UkJ1wCzY4ZDdW7E0f/M/D9oOlE
FjC7bx6wLHffzAUXk15n43InJ0bX/Kdh6Y2DH5L2QX613SHdE13ZtxgkZxVUcdGQ
ZQwgKUTAMZk6aCcyfbBRmVn5IeEDaa8GQl7PkNNrDvpYS2/DBLJLNNwemDD+kbQE
O2cuUND6BjktZ1XNN8dMlmgZgeOhPM4ir7qIbTRXjwSc0iGHXlM+UFKE9ogynzM7
rHIu5c43QqJ2I0B4JunON81YAPa9sYZ4nbA22tXn64hwDky2aF9d7aGjv7JWaGWH
ilc7nghKePPBXZxNyy43hf2YGFmeITOKatqFGQXgOVyZ0Ap+R7l2cpDwNh34GYS0
1Jt63zC/fJGVgrTDM4/7MKr3bNErL3YPpclCLhJGd5+OWTFwXWZLpxQWJru07nEx
1IMIcWezNjCRq2cfgbkrxabv/h0HYSomjb1NIr1+bbBMSAc3mLtTL5qxCS2dXroU
6yOrkwidalEj5PLdbJF0cTu+svKjZuNs8mh3fqQvcBPj74NlBXTaBmnT9jxLtQJ4
GKEqsySo7mMlcyGcISkjobSG2tEujCXQI8YgeyGQ/TFHxFoQLU41GmGNVZHv2FRc
saOwrwe6DNqgHQR/e3HZ1BQlWJsDpgSDcMzleDgBQtB950RUjMHmrvDxIDWCphjQ
YKEgl1y2/izEe01MnexdDCTg4PrZKn7GkFXRCAHObb8WF9/XbTNEd0NO6m2VqYnw
l2tzuuPWPliBcePKeO8eBcJKYdv7EOIBe/vMmIMa8uB5qyVx57Sx2SrqnTg4RFlh
osYSx39X6057STgFMJHPUp00CkRs/4C9DyxbA6v8M8BJHvlxnOrOYszvhzUq6lP2
6Q/+ma4Bis9wdHNgzS2UheunCoTawC/AeqegbUQIq93oH9mhWNCWfwjZtauJbEzZ
6H/OMAW+zmXnuPLZJndn1lfYaM9MpVj57915LLKEiVdwLo1ssIjGiuEUFcEEpdfk
mGVSflz4BUqCypcCck8ywUuKUvXYlZyYR4CN16g1XJASdoiDpZM07iru7lbfS+nN
C90CJIeQPN93DiSRE3xyMFCigCAok9siRqXtPENuD40RvibDcpI0PYQbQ+N1VYn8
irbBBt3ABT/dN2e4h25DeVKrPdlCYwwILUVW+2StWXVGTpOeeSxPPtMhmgkq6MCt
6GAfPXiyHK1BZy60rjnc5B40uPoJKh1shOIyyuAF+zycsqmTUiSVmQMR1YklHE6v
ciwI7yfz7XgeXI492W/UaaDVZFqsFhyf8acr1cGxvNA4yG4fSQmPmt3Yx1yCThZl
Q0eFhv0X0pClRW++ujMciPaxVsZuDwSj2oImb5B8+UtZbZ/xg9gYCdI+9d0tkRrc
Zr+rE/22xTeLtgRcnxE95I7iqo1qD8E2tOsAet5Em6G2pytDfwe1/EWFO1SVmoAN
xHpDRAb7uximrYQePLjjCTOp2nD8U1y3KHPQSs2k86n+4561HxvPapZpWW6LmIv5
KIB3SGGu0LITN1Z4+4AO4QOh+tquLm67U+qj74ETcL1ZDYjIyMNX1lFTenQDMHs1
EZIgxUu9HA14pakweNI0vAzhyYlyyVpZqAH9PmG3nBUzEQD4ldEAhDEAPtxYzQts
wHwuYSjGmXwd3Cw0FZ/Qk9cAb5gksUTIYKQQwgB44u+0dP5UKCNk/3mZStQrnmZO
PuwbgAMuQbCxKn+u2QARV0P3WbeDVKDlpNUkevgQxEHpZZkiDgsKylzA4NYqhvSo
ktV9vKNFV13BDjMAMio1GXmzlnxyieQppDBzIVYJZfg6M3AwduU2ZMsgYXgonewK
+eHlPNWFu614GUbFSkZHCCQMtGaTiLTfBlgIeGLUa1bu78jmWcYw8KZzQLg9cbVe
2VOvcHNyJDqAGPlrVMPKlL2MIjFU5EyrSr1JzC4Ko4qLzPxo+g24dzPT00Zho+9w
MsiNVZRBtkwsNxdwRahBfYVgbRt2JMdF2+ibbtFDyB1tv3DRkOFzg2JqGD9TVEEr
g+IeZnp3baBqRHr7FMtKssORU3uioSBFKBfB0+Kcx5D5xBIpVPqF0hgRphwlmAss
yT334JrOIl+de2L3BX5FfJxp8nITaltMC1sVScNOtY42BJ0PzXfvSsfukVrjF1pS
qLGw0iz0oj6rV5VI6KhTlTo+b9ay7Dc1ioxptQCn5SSB0gLPCbAMBFUE/LCT6Zpb
mEbTXJQ//9cNhNnG/9TEbL/05ELyOwwJqeHjrx7XIY5oMz112bi7I29Xo6gGDMs8
Doa7nw7Fqa7OTDcgEwdNaTs9SvBqH1istR6xCWATu3bH8eFkWUPRIjlUekfFesS7
bSGimLbHeu6EAYV4jldLRVDGbTLOH2MjfF23khPVbLx0rOKWbG9Q41nMA1qPyHPJ
byUqkpfFvXV4dNMiqpnTuSTFEs3b2VSG+yMg/ckEYO3+Frlzti8GI3v6zxMMImXp
VnA7OXuT/+gGO4W8E4sTEaDTQ+iI6xrYRtMe6IFOHadvJSXpap1jTVv2/qxKk2PX
cfovKR3lwB0q69Dm0B3fEo1IlrLltIEtIUqwCZJg/Oas75MDy0GxYwkEx6N+Gwos
c8Hq0RVr21Karzkc6gYUvslfgrgr50jhThZFpk693JIpZFqtb/RyD95iZH385FfW
4NTOB5vz3WjPdtr9VaZzuWtIfz0/z8/P7HSdrv3IZDg2ER7p0kohNtYgkLmtABj6
ODe+fNbQ2A2jX1Uvw3fOyuADPSjLeNKNtSljG797OiO1s36EXrWI/NJEtGSpLxKP
R9pZn+7PRct3zBunVSkBnl4VcJpUqVEg5wIiv3xkmMFQjaFKApQi4GvTbrzVHRiG
OZlFtwXDJvDxsnTba4hIMFN/xM7NdVsApsrPuE1C6/53zZGEGEOEZdVmAQ45zM93
zxCmf8DyyN3meUQuSCXeMnlPH2Wnv+E7DirJT9I6gY8i+9PIj6jF5TFck1B8X/rL
5VA1c+gZhv0qcpnOCb18cDX3eOqRa5KGEWXBjCF/DkCyQurQQpDasWunrv4HpxyT
8z4fUVQsp5Zinp1WMtSiLWnJQ1/no1KyYBgn80k0vE7+asXz6CS6MA9X1fCF8Pbr
APo1CSSpm6tnHaray20A7tcvw8ELkTIvxeg4r9SnYgkHOQrKuAPTvUJhAYc0loI/
fWOyAu/+yaVlWfxCxm1mMfWOv8OdQrzZNwMd+KUvG/pK2h5XkmRlANDLw7MJ0TF8
nhO4EHvPet7iOWGxrZ7FEbJ0MW0luozbZvv7Qs9pIffbavcexFzefB2He5kPE/bm
4l/xxYBY5mAb9xyCjmizCAQxuyxB5UdQ66FVPxTYdCQAnB3JY70GcSSISqja0waL
FjkxyfLLOsBjc0OZKL5SzafNktioDNkZkltMnONMQmWZttks8WLDeoBHKBHKfp+B
vK9wZ8c6nem9RZQQ4B3NXrAf6vz95QHAl5DOYDg1v+Ul1LTKvEMKk1kKLLnv+xVW
kTsqcKJ+G83lKt9hhvD0MsK6iApvk6AO1aM9d96cMSlpvERbzHZtugF4iyh8XgvN
TJAWmED3KtRapCR2ReTjChstaHi+ItYB3DI77C1+DCLd9wGEni8VmdfAdc8CN0tr
0T8BSiYzfXUDyJJ2udc4RMOrQWLBGWKgYTZlla0RkQUwQqh1F0/Pquw2VQkqv0AM
Ez6HrM4MTJOFDmAgFUrpDz8eCEpg6nc0BtNzorkRmt/al0Q/oVcCp40rvwAyEPTf
ziYd2pj7OdXeUaRg3YuxjWYiZ1+FGo5US6pWBcWoFynwHu+McZnr8jQLGgw7sC52
/EReeuYQoHrCYTEWW603zKdiVEMkA1AiU9RAK3Scqb7bNqPeQ6G5k9M1bDOpeMBY
uCka322USZ1fKMAN+BioxVjQH6yh0z+J3+uub5QEQwqko9FDnEmhBmcrdHSRdNaO
cB5Wu2BSCGVlkJUenGTgDiHPVmFLTV4pe9s+WiyLTBs1OwS1VIJ1KFiaL7JQElAq
ByAHEK/BToPXf3QY90sm5b+nIZ7XUShYkX0zDEjodhq7bQh8PHSDsF7qx+BQlNQ4
YgSfj8mq1rG0+tYjV6VXp88sWi33e/0ZNdgSUgS8YdTWxW5dyCNMl2tpTKuNRD91
U9+vpjySdw2mdMi0f+RjJLrVz3u2aqL20GGnRogFqkJFUKMkFdH6UoiGhIvKLtbe
9pksfCZaElni52KADPHhhLIkb/IK2ZK9lc1iNow9kBJlzQF7txBj5HYKSuZgqZ8E
Q52XEU/FwTBhasVpN1z9RI/KNZtZ1Zd69k52y93CBqtjGHkXq1W+0haJ/4iYXy1I
9hkfpGVaNPUy1tOW6MKrzlADjqYQ3tF5ld+eHnb8J6cSaHL00AXBgzpi8YqE3/l6
oaDDeml1jYtnOo9EBAtAUC8qM6p+vF34Y5cu9fFM9n/6Mygboqj8cCWUuLMTFi8U
uD02oigdXadF/FIddh9QsclCz8nUQc72P8tyrS1gyNdHOmMIdVKRKssMQIsZFPeT
Vd+JTfL/W6WL2DwZcsDz4Baw+1GpifPdWC9JP37U+kbkF6vwUe+YnITEhCaymF5Q
bLzOEEIdTJYyp2/M5ZK3vTgPEqi1blXI5oKUTTzlRxTnLjxttFGZo2vWNp/s71qm
giafU3XwTKWC5EatbzZ+gRWsl0J3FurTKfdFchkqFabaxE4E8eoSyar2XMt353YQ
L0knOvsGhyG3juawuSyyoK8U/u459N3SL0sJFrLc5DCm1UJ59SzXAijxx0Nk4tuC
jBkCzsoUyQS2GVqRqZbLuNykChdFS4BTxpsh70o2xI906UH9v0DilX+ujNOGy2EP
AWuKD2ptvyGMPfySxf07pob9FA3V2IkRNI6PBLMYNEjU6AUfrF3XUd7DquNVryo4
4AvLZ1n3siBCEcuwEFdqPJRTCaytlWBkxBHFF0pJdJDbQVRAH5gwlV4BwHL//46T
rGfG74U9cNtrfW6O48dDifEDSAmjWEBWHdmKfSS5WC1jxILelCe2fFVEe5oCJewN
wgXz+6w5dj+Tr+UHpzAAtszcMTWy8RLly0z01MuKZ45lRV1KgRvtJRSCAIMmO/qv
DxVk8xiXRCgy/X8E2szM7uRdWtFvWUhHh0e5cxmMugdpy/yCaDdpqpmwHEdRh7OR
Kl/F154J7T83TzYFwMJRgfiCUldVkSUN4LN1wVXdrklNeNSJpmRfgIqxmyYFvb0i
XeHB2RduaxpRAGR7RrGy61MeSZdait4PUmxBui+Iz+eHoj+G8iNErJxBX1wD/9B2
yXcsPvg59+v1qKo2yag4Uya0QtRuL1PZyyzQrzQMJRlzeYZs9wJx2mPZl5iU2U4V
AUzYMDHdrXEE3sod/067reB9btrqlLFKqXZ59/ZteTQ8jeswRNpt9N9LzWvFNtXc
d4yAQCvK9XIZ75fP8KXFNDIV7hmnYdH6k1z0dVQAqdcdsIPnsWI/P6QX89w4wRyz
JuAvBlg6F9kpdeSlBUG9fQ78LJb2V1iKN8O8pPigr2Cg2vbCDLswEwYILKPwJgpS
TkBrUX6ziIOfktozgZ7hQok/QsuYZf0EDKBVULLSlK5Wk+J2SyTxuqgun5wrv7kq
gpWZjx0Kf7VTbNTMlmOglAYbUZ3wVLvhnaXK15CjGNg+3AfNLybMEuwKEA9RBcJT
pBW1DdYkeZez/hhGZ0tSwZ2QpA/L6BwPZNf1HYpygsagaiP4EQjSwCPy4zwJN/yF
vSAZhQNWDEd3P5ro2g/wf5hOzC31lBntlLqiESplQJBGA9ACM3VUqrsX4dMEeEv4
rBkc/3XSZyUDUd2TJn/Uf7F4pvopA4ot6nnpEbbvduQ=
`pragma protect end_protected
