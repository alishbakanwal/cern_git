// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:05:42 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Se0ktF6GRMfdBP3wpVSMnyUfIni52szCAbAbcLITCN3QssxUDNWuonVB8ysy0jkf
739JcGaF2iLdE0Uwyef85eP02iV+O64Cr96eJRQ8FiKzCIqXlh1qhL62uoi9Dw53
XHJWGiHU+Pq8ozzB8ONtdGFgG+cG3pOfYKfaWT0C1/k=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11488)
gi8gvf7m805kc2q+MoMoH7+nkAmIkSbBwntlKhvMGOrbZZF8YHJd++F8TzQe08zt
rgA1oPrwRCBtOYVWgeSQ3jlpKbNBhb9C9htZmy7wpkReWCyaicZzTIRtD2yOWzN1
s60ZoZ1Ym6XDqjbQI51Bii0gaRE/038m5U779k7SLwTE/EQHrMghGB9LPST1xMH0
WZ6XMPhBpot538MjtOUjQso8HYzu2qFd6E/pb0rjmJzhjSWlQEU0l9FjQfMq4t52
SaL5Vykql9SM0c5JFPpLC+80pAwmK1DxKI3VJnxzqK9DKIZ0S7E6y9JP8grHp+A+
yGSHyxnf7FfS4mfRDmvfYn6CC2oZFmGmGDJKWNCNVKyZT99Xipm7dz2ak/6GcjiU
bU5YTNz9CzOu9xrsNRBl5vzr7VNsnYOuMQ2y4wWzonK2uGBm1rSmRGMaqo8fKH+P
VOl0lpazP7ewWQEGGCWVp3BIQ+SMA2stStzxpRZnaK/VSioEsDU1yigqR5sH3KTQ
twqSHZCbbWKLJ/zvw5O3AArgl4kmSuJa92cZXYyrGbEMUjq80xMJZthyb8Y6f4In
zwJ+6We+Q7U5bhzBYq/jK53Mx11cxF9bv11yzEKyLsjmd7LFLrBUcBgFkTzNClbV
7LrI5zjaTdHFKgqOOi8UTSZ/cXa+jnXIonuCTuro1zWgwomvtufQ/nzjjROshSFs
ueSe+3l+Z/smDay3z9UhCJyvIPHrbxk3A8oH8ekuPPMcP1xO/+SMM8R94UtXjoDt
c2vTAm6szwP6Q06fBGDwRTk1PWdFDMevuEuUSZabpSy30Jn4hEcpYejN6q44TwOq
nMmS+ipCohFueA6398EEsxHuMBaUcpBcZTHCmKTvCp2aGEkx/ZH8WTsyLkdC1bQ9
5APcGizF2WWJqwFTJcZ5hffEySWf0HviQEcNj+cTIYn8mVOtVLUlJeWpnj/Gyk8A
IUMkMPTye71+sTOKtHRxbe2SKANdBybZptsWlScXaul4o7WBRKK+YWwXujDT5K4c
BQFzttHEGx0MPTRdek5m44Z39MSgFW7V0lKl3BBSQrHhDEEA7gSK0raKoQR4mh6m
uJVvWiMEcuPUYfZSoQNBHl4mj8NWRYJrth59aAcCzctDbT86X/vKw3asMgZUgg3f
jgoyGAgoE3M84RAynDkd0iqASqY0FABIZVzX1Pp2TA8aqEV/VtaKp91DeJGTzm1T
6hhyxE+1KuiyQkVxJViB2Sn4kc60oFhI4qLy+0YTDbUnpCl7gXdQrZwmn+BgSYDw
/xqzw01q7hcZddnxHQ7RRMpgJBCkNEVVGTSGl6YrFL7jBM4E+3wzFmybbk+ldIPK
3MZdNPEYu5ivc7U37TqbQ2jcDBh45uAS3GCnHYZz62c/ETtt0yP/B6h4z0YJNLoQ
4PM4PRzZbQuu3InXLTgz3k4W70qIecQOV+xjYN56HUBjn8TwwDpUpNjwS8+VXfk2
XW+X08mer2FD6Mbq+juaLz9giCW9XYanBQbPDGct674NE85LdvyRah3m/YwEshYh
PTS5ve2tQynH/knIsndpvabKZnfjE22xT4Zg7YYjkQsvAKGyAXZFeR7QQE5hqQ62
ZgqZOjRv9nOmTv1sZKushZHk7Of80Fd2Ll5uUge6sqG/prg/+gWRiv/oLyHKl8v0
2HvGee1PHU9Wbc+Oovwn6T0IeWv6xUSflo1aZUFO/xwxX46Dwh0HpnyZHUO/02mp
d/J4t5bF7vyhjPb3ssJDPIftZnuz2o7tsrr/SiN00u0A7F8Xk4NSkA/g1o2jQ9Yy
wcNhBOSsBFz7Wob5yMZdiUOs3x9zLX2rwg8iAdr3xuXtmwLkfKb8awl8d01OHlVP
bUneb2A4yq3OSLapmBqHhcA+rL+bBh0F579RmfOLYyl75YYDe/LXScZpCkQTztSG
Y0xlJT84QLj4EvN04Hew8RaKc08O4IuMEsGyMC0cYotbrTFuemXfj++kJ/Szzuri
UdLWAezM5VE+Jg7cESjVFmBwEwTljxG3sZlOia6zDRENAsRVamzM07V+41FWxeB6
T8hHwGLdZ4NgmtAFE4W4JQRJLZuRkKV0k6j930X7i1iA63+thhtxT++h9wkQKThG
wInKPmv1pMTT2FGvLYDuH6tXM5mcVfDvPGafXu+I88vNWdziKLjIhnRMmsHKgjn+
zh0irwtF3ACXLVqeuKuHjdwBqL8KwnfknwxWHh1q/gOQGNPmDvi0PwDYhU48qckp
Omyt3AocRFBqtof0ua3fLc/HQQoz8Vz9G86dr+rMph8J5VsymW7dWvIckLs6fPog
WCLkvMm/g2kuG2ViINhZ1R/PBwW3lzUdODbe25hIE08IsbS3jL98eS5N6t8Y2pJf
Wn7Fjayb8s0a3cjRUC0AehEl9WY9i7EQnxHGMxELDLCwB7FFne4FgvBe7no/Gyba
iJsnGAMKKdjgHiExPzx0eLPPYmPSJLJi5eLvuYhUsWp4j+NqpekJx6JWv9VMQN5J
u5hWH0k07raZWkZdUesEYDLFb4GdekSq0zwdKJEtngLYFn3ATiCBQCsSD0/qXLpJ
1O05EOE98jirdY3IgkC0GwuUiXhB1zzpXcnxYtZSneXfVcUYRU3MoFyZ4VCmBlvW
IYPKztUc6QypYAa8pUC+BHciKlQMoiYLJ9QF3OFg9ATgK1EeB5W08RJKOl5sUF3e
ffQvZ2StLL1+XHalS2TqKWqT3YvGy+Lgi61jOb57Zdql+V14sIkeWzzPhUJpdg7q
Q2lNOVJ/KB0ve/3NMdhQ+MXavwV3n0tByliHVUyefAKJiQolE1titESMgI7Xc9n9
M/Nd6gSHkqCV6MM/t9sf7lHGbF0k4xLD0VRFdEe+gdqMOKo41pjXuUzCZF05sjhM
jOCDyjploFqJHgo2tLUFaFKDiNQomXP24g3tYUMIFH3NuyQt4AUU6b6ov3lt9MDr
gIhhKqkNq3NM8HgARHLOvaAUuK0sgTsmfu3n1sA7Pmy/8D1CWodXvvfgDcn6vB/L
8OCAoRSAHzUX0GsqUdHSa8OjDX0xDnQL7oQTxsx8ov4SbHtXY0taFrqwRFsepNkA
c41TutJh9GOO1VMh9mZNEKYjJnKVn8047RImVuhIS+nSDPzj25RbwLTs3sOQrx0v
i3fet0paykTrnTm3QXqjjNChFpC4nXQufhZ1ll860+x1w/+iMlJQqiJscV/KNAs0
MvpaYZ1Sv9yOjIn78pSVZw+x0U5ATEXMCRtSqjYTeIM8GXp591X8v6T08SFrITDV
zZqDZTgvFpgMAwwTApGeD1a+cdpCcoaZiE87SsygFP8CMH+TBL8v1nZxElGh0JWn
hREEIbNHz7/+1uIbhZ4nUME1Lp56pmKwnbc0EpAEBgUyGo71/8c0J+tnQAhMRFzB
lsUrjDDaT5hJ1MJIxqHyfWUhJNZydCKHzroatepArka0vG78oFZI4RhF3ZXSIdKd
l9D24ojXTVS8yMaA5619kTq2j4GtKkOBWUVt0tHXeN3wL8Sl/dixW0LKqeUuHU9K
+f8TWXez1+K+9AFLph+rI3xIwfYYWmOixC6/sLS8A4ePI+lSZ89BHLgnWMYGElm/
unDH3bx97kPNes1ruTsCfy2D4GBkMCE2fog6gmnwDhwlOi9NLTBmQ7nB0SpQXLmH
5deJLRR88SwWeswlcKxMr4JE51vdHfVee4A+ZN6/TzEIFS6ImuwCg7wh3pdCfDU5
5cLyH/4HfwVUgc74ScpPlqvA3DX3Mr9NRsUmJz/7/BYUiHo3O0AXRs7+BJWJvq/f
VYbeefyCs+w7MjlkaBRaHsNcFwtytuxSFCZIdd6GFR9OoxS9g6HKcdlGabM/d9vL
Fq+m0zQpqT0CJZbfYbawA9VnAjInB//zkgqKWAKhv8nJAxHqKC0+M39CCRNTkpe6
ky0AmqRBcwPqCmMWVE4FSDu8mnkYuykyTTt+afJRZG+9620OTPfd/qacjQRS+ObL
JXGQGOrIkopqgXXQ8eZoZdoyxEHfZNytcb0Q0p5acxzfYj75PfMgiXVfj13jBSdX
dpuwOQgM4Ne6KjlA3BwaVcwmGK53CPKnCReJR2pvVuZjWOEakTfenEsi7jOc80+V
xVy8F21EW38sKh+popHoW/j99TLYdYRrBiX6IsSiHtpnREPmpqS4D+Ri2/xRsV4j
KuFSxxVMVA5aJNNodGSDk1/ixx1qHtEetdAct6GLxJZz07i6vvyNkPKs68yxj8mn
w7FjX954Ah+BUWFWSSVh159XMPGQWufzqUPCpgCJ4Ru8cemzX6amYQkNv4pfzYJS
mmOv8w9Z1sYrlJhNXF4XFw/Xv7QxIHReb0AMNHbRomGX6ExgpLFLHjOkmzkC5JG5
eTCXwVn+LaL1K2rJ57p0P+wVE9txP3fqu0uoZbd1WtvBF/CJBXHRQZJEWAi5Mkcg
jL7gQ5xvHD2T1J7FOKFv/ODRaFWyiBTcl42EobCDCK+2ysTUL+CLjnw7k2rlHf+L
LxWTFDLS7paSGKvNwTFMwhYTRPjYPGYBUStYDJCv9CGAMPUnLcdpfZ7SB/2i8xH9
vjAAno26w39XyzAOgIy9/v4UvhAK61pFmfcJil71jb8cKr56AwPAdzl8KFYZ3RCj
GD1GzJ5pkcF4UMDaEzNdAtG9DIYOJzJI7oK/qf9a7rYBWVTsUa7s6ytGo6uP3FCs
HNfr9omCTVJf1s6Q9BABOiMRhF1bU325atFJEpdMWPJ86GBOiDJjf35Q9galZD9W
VkZtpUMGfOqEK7IelA3U60k5bTOd7UrKekvK2QJNjCM1ad7IMFHjQWfikpFBDvIN
X7o5enDBHKjzX3jGgo13DBIOgM831zseFdbmJTE0JHKDmjeKL4cFvZ7hfUaMLY5G
MNtPvhJh0FeRbTyU1wopGqWEfzLGJ/bhLmd6VCz8hUZweA9H/Vt+h/WwUELzx4w1
x3xAHbZoaku8w1DZUoRea2Q2yHaCl4NDSF32EJBc9AO/SZudNFv6iuVhk7m1oKSh
fkcPvhSQmTBgACPZHs3uBAkbIA9xQ/2ZlyTD8XZpPzBGsDbBo5fjijRqa476bej2
986Km3wJt2MkVhtwFda3KoulemCluT3gzrlRLJoJTst07e/I7XkyC/1G/A9z9am+
BsUbo+O6RfFSNyKhvzG6t52xnaCg1wxjUnLfWxn4H2uNxBLMizYGGw2CN3arAhkz
FH8LOOqk/3zJ/xDx5PeJoKzAiMSamciM+8crWMKMfDKe0HCSoNYmL6+mk1k3OQCY
Xn/8+nviGTfOLhZk/nIPT119dKR79NkGei0sHBnerRk/v7O0Q5AzhSdzznH1qZIb
BQOltcPSUZAcHirIqzE8Jg15LtOv1GPbuCfgt4pTgWmCfB7keiJF3w8TAojXA7Om
siLzWC/z3ywqCSx9YkKCszm4uqY5MI6W6j1+f2kPmX8YkPeEPNovqB/LF9odYCP3
IOOGVK56elPyyAEk6ieilrvXtIJjrlCFrTnIhGEOEvftPVNs6AIPaI3EfIldRzjM
wl1zWWaSrAyDzc5D+2g5ZFNWW9JSWsueIrRUSGrGDJ6dRiTbzB0HumvmnBuZKxNL
tGM/hMeAk1zRxjTGmiGLYNulDKfK+E7AFXGAfYaGHIqvRoqvBah67kbQ74P5R79O
kbbQ3FCZv4IKi7YIt23927iC/i72Ae2VVK9cOiMKTZp0IYmECOxPWCHf5hECNoJG
aUEUeOfupADZel2Hf3kwc0wGqtfjiFGK++zmzvrw0ZtDjuQbwk+3+QERRV2T1XsM
PExM/DL8ff2w4VylA+HHWIUPs70uEzzsaF1+WxNpKH05sgxa70tJYgyCZSQjyzSB
DHBKfyMJBHSoPmBzwaDlWde96dI/N4iv0BFuC8imMYTMbQkYkcBdOzaas7XAO0IQ
0IsmmtZBZPOmswhwdp8MbVmBrNmmcjvJxtUKQI/NVH4ZVH+d3PWi5VAlMVvs6HV9
JBhBQ7x9C3PnY/GlzMvdQJZb+D1tehrLDfXqThFOV6tVFPaTbDh9dt9tVF7/hWcL
hxB7jBXM6qFuGwETM5C76ceieG1X4rBoZOxzC/gl+KohXjZC+N8Of1W4A5v5n84i
bp3O6Pucnip0zDNx+W19x+7NY1ygKPtU8op+9p3SpBZnJ1A9XbKI5OjkU0BJEJ5I
lmY7Bgc1xbqIbHGjQa6Pdctz+G8BC1FuTpuwUty3Jd7Hbc/6FwuNe73efGEOJquB
9WmMlO2mniba1nUSb/A+gxk7oyFKVTM8m9KAlH7BN/FuMo+10kDWR9Xa8i0Qjrg+
EcbEAchIOFDLbNdiclnRTTMLFm1itsqPS842v8GYBOeg5FrQR8m3R9YWmMvBkh09
a+y2NBSRLMqvlBIgoCnYRt/3jaBGbs/T9fZhCqkgEnhJnTUY+dDsUqkHTOqcqZoO
sB0EvrLU8YuUvoiqrsXmVr4d56m0LANSN+LycqGSR5pcX1YE7riiMdYqY/iGeril
UgEZ9m8aoKVb09eFdhHcQfk9tBcSODHYeDX376Cln5u61+2E+us4h2C2VU1W2mlZ
KflZArxx9bdDat0wOaTUZmP30OIlPUfvl8HGeQldhWYNfSsXa3bu9AGWZ6R3gVIc
eFxIyMyRy5qvN2S13GvAPf5hKy5cLKAd247F9a7gwLNHIiFzgOoN337J+HAxCjD3
YKDV9YpSmvwQZpvI/PeAOhccXE8NfCDE6hBG+vXnNr/5/qbiPlmv6oeX0Q4sfO4t
2AkPunFJsS/+a7gtUKwXmDqjsJG3RPJCMiWU/PEPpCzjZoWXbXAZjFOUxmLnxDwt
YEpsilhoz5j6DovNFabQxJDlH76um3Daj1OrjHeLm3REZD90Hghn5aFeZ85ZC8wn
CXVhVUfIZ9q/30YDB3gqLAqIoZPtNvrC7y7llg2XH+gbyl+tiQKlhthUEv/+47fl
V8RKwgduuP1w+P4kiwQJwkggJA39kp9aKDSw87vDKaetu6rQssB7ufbJx0AbYzQ1
x0erzGTY+pGUuWGJKjahjAtUhm1F7RtHZjgYoNVFG33i++ZxssICEspf6fMLaIvX
w3tzHheRbAmhhK4zX93qqpeIT0WKmnNNDQhH+Gg6P18/DHXM1jrpL64NtEuFwW7y
nVnaN/xzAmUejU5FNVp5DAfs8Ax5HCBZWoEcPX8pjCRXKbIevTDCKFSeqLjJzGy5
5q0qRs78+hAAsi5S0uwnMDTllup1nAyGfDtQ4BOjBSNdgCh+UdFt1x+rKdaYvYj8
6kRzDaQenxXdygdZX00EUQqvv1gGuja+v+wOxTEW8wkmHwCkrOEx51r4PYrrYGY7
XU/aeft3wYw5aRGIlKWgcQJvEa3/iXLW8kNMpOURiyMWJ3UmZhHlDt0Vxd3p0m36
7bTMXtU+NCKZSP9jbP/MpBehxcovSWK9qChLo8KkqjumzCX+IxODm9Yc5eeQdZHY
Fg7pN8qoq8N75KbhnF4suoupYQezCC+m5+7ZKXeYa0Yc+l9UQWqLNV0VGQDb7ANe
LU/aL3SnepqZYpuO16ltf/9CIzrljTpyVorfqOPNlfbDdURk2DWyBLF0oY8+YiLl
mm3onIKenOdR8WDcWLdXeDZxNwATlQOcWuloutNcBfkRWhgZ/Qu4q9ywWf16djkv
QBoO9BpN3X/kAKL8fdH75YhqOHf+tx7EFzr+1rILEkA8v/NSeQOIHbonSLJHuh2K
M4Hm611tgbmDHoDU+A6nbSmRBoAQXpQQDcAKUEuxK+ddtM9/AT7gqMZZuZcfF2V3
b+EpeHPHmwyAJjKYtcZh/iM4p1cNI1cYil+sJyLCR4Pyw+MX7Hmxk/nu039QjQtr
CnWQde2nOGpW0+EGYs7m4hJO7VRmBU/3vYxwNwLFEMWiQ0jSELtFhmIPUkWdVjfp
PyE1zEHVKj+COTY/qewugkDNGiItFfAAGT1PFCChawJxT5C4IOmNOzZA6wHJRGbe
0L3Asru43TP9AOnruqSwVzm0ynZXW7DIl01Mw+mIXcT31KVzD7g+8TsYH0g5YvQq
kRWDCvUG+JXFyZk3rvDevvDb4mp07WYu783M4rjBdV4InnZ1IXQ88Wt3oEK89Z0H
f9QVu5CVnMrhHn1miqEoUMxumJgm2dOr+pRczgkwaQOLaTxQFMogQiwm0rYYZ6DJ
WJUCeLlQ3GxBnmbmimnyB32u46k75jkUeeDyJu4/jMXaBUSCOotvFF/exfim17Kf
dyiEZnkTGa52e0YbJ2afORvkRZRoApzomY9Ko88mxvk9mg/41yQmDvmuixkzrRTe
sgb9iBuHfaIjt1TquV5sukbfoLgEoybgWCLFCqpzrblZ+vE/R9bpL+Hb/qdjhMSU
0zEjiR3SZFfNDHIFjTR8kNOTTeH4dR8tmAV+4pnfPoq+QXdXS9EVTMXB1RUthJTR
mUl9dQb1vGdPUvrGpMp9fM9o/8dBatuX8JXsI9Lvcr0Rh/23jxAc80a5JhPCdNgu
XYTDPXEAd+6UhWQkjrdeswvJrmM8JoywihipbiFIP2JmYPBA9yQIO8FxV80ki4Xm
6wb9wODL5RaYA9Egp92aGqltiiR9u7YEdegMGoqoxt+WCsKuhUXGThUpvuwtxafg
mx76DfVtZimtf5sVP7qnOAqyrze/IqfBBk7h1NliU604h883oDyrZi1hK8Xp+evZ
ozMjaTvhDCNKuKRjQ+Mwawx+vJsAUI76m2D3jERNGtQy7fU4089mbD+Yh9zAMEDn
w0oXYvliRuEDA/HtQFnOj4tlOXiYDQzy/pL/UaXR0gnBcWDNrsfts18KnKqDY/F+
70WBgEYrol1pMbrTklJ1cNJrFWS4lVeBVC+I0PnrvurPYqxEl+Xfay5VYsZvkvGs
vUgbq39SuAJSA6FwVLKqz8bo9I1zRW8wXN3n5T1XayNhrHzC2qlGjEcoCFRDp8K5
wY0skQuHPDi5F8J6GfylfxoIFgQLsCfaRy15gAWKzaHKzCf2ScaFqyGiJ1muAb+M
6rq3EDfUuNqwPQ0K32oxqiaRIlIHnJ8emMvYOUoqkGRYse1iXCKUEQ3bdfvQNWe3
5574XHlTo6H2WI6I9DwkrssUtxZfz0WdfyNAVHT8BWr3etlQieEoFMUyY0ehFKm7
do169S9/8bRH1LEo+6MKvJ49mlaMdMCk4S20c15wIfx5yO8d4/ZUBTHDcG1mdS75
kG2vsY+hm+akoERRZKZdIXC9FDP97UvWm4yidnngsChJtW1dNWnunv/e7B+0SAgl
0QxzFM9qHbyPbcIkxOpZQPAqpUxKe1HWrHdBLoJYeFyZeJLPUV66PB6zVQ7Sq1bu
o4i4b+sD9miJhB/h7BXmT0MCmcDAHNsisiTu9oISvEalBPv7tVmrra4D77E3pZoq
0Sb0/3uFgU7MP6WmdwnNcaHMEE6ld/nVXVFdH5T8OdA+Sq3vrYaVT7HWmGLXOlcG
T6m0McaaYUMwnvK9src0NV7RUpC8Hp+AYqNC6sIee8jgnbAEhv/b8GZZrWBgbJxY
VbVXjm+Jfq60g+tlZtMHsTbTacq7epEiM08U0fMTvpJjQ9/83OcAzTgZYInKnFyW
mz5cy4+xXKK5rVg7iil1zJ0PntHpsv7jBbTJk0/hfukqvjSqodgB0OQkRhyXwLyk
AAdKlWm6aXp7wcqfeeF/0Zxn93e2VbORdh2wGp+arEn6tiTRVEN45HPO0jQksvj3
5uz8SnywsaYiQG+pkahDrnc4bdiiCdWhCpjhtJ3AoDeQ7CkkBtCNhCF2M8ivBZSo
d2gxGxs1PtorZsgVj1wktDiR9M4s68R6dkK13Yq888ZJHid7dSmv5qdM6D10hECS
KAYM+7b7m5UK8E/ADrlFE7YkbhMylBxL0ImepYQwLReCkAljgUzMg0BE7UnNf1nc
B0bY17SyASWzwhagBJbdyLINuRoZJNLZ0i2CFM6eixBNXJ5n/xFCKqjH7SxffwfY
iDeq3RiHWJv9VulZOG2MkkaGuzX/4pa8iHpPayjH6hePEglRfUClMNBKvT1Ued0K
wCMkjjlHOLAyAN9OfXIeH/0PNYHapr1fglPIu/Xa83PTpYfpjGhjI41rNRreGtgx
cs3nTyNyKvEq1f7nvqtUvCtnA/FLDfP0nF7rfFE6mCPMH5JktiQ0kZFWIcXtvC9Y
W47dbFf6bnuxKvfckzRIaTLJJE7qPLr9+/Tiui4xhvCi2czF6sXJUjObrjEa1UJu
GkQptYpwwnSzdW6frJXX8GwniuoBu1M12UM92nN+Cpbq7gfvX9WSMpv29aP4jaXf
p8uSv6N9VULf5YECu+gX6Dk6TL9ZOj1tzR0rd9Kp6LFIZBTO5Di2pz2l5XES2B6x
5t3a4cSKGg9n5LC9Iqlu9G+hMXdyJSvDK1LvYjWoZL0Ez+Zn2Axb26DjO7Rt8RNR
ZQvo6BI7ZneWeU+13Y4ruvOSAvKW2A+GeCSOkMM0B6eSBIe5DP9VU/vnwNBdblUP
sbxGuMbrzKTP6eiH3GBs1Hi4ghEL4ol8JIoxXT/5hAGdZql+gSpbHpae7WuNZKXX
xK8DqoaYcJfKNytXN8kQki4mIb0WCCGQBsjIpB2IP2+qs+zGDZh3JrXG9M37C+q0
GiAwkAfTWYBkkuQDU9Stv8cusKoOFnEl0Yqh9v71Vc/VSz9eo9dw9fGG1ClfLQ7F
qdAe+iBln8djpgPJXjMv35Qf+tgP6GJdbskHF9zOBVF9uaMEDVvNXGK7po6ZSBFE
ju6tvah47+68sMyjofRuvD8F4TIJB2OoHcl/yvBNb2RfKXGVE011adxIuyDg/Q2D
2psIrn1BIXI2tRcMB1ugXXJenjyQxykhUumAqbHSEgAsqkHVAngiG5Bs93Dv5FDJ
NgKs/bfBQNgVACZVx8ITirIPV6N/zC/MaR1/qhDbfNDYeQMhdtByDIuHHAqOwt/g
l4qoOeuyhWCDLN1XpfvbNOrlGRXSFEnQslDF8J8picvTdwJLXrXKePaQPLITLhbg
6cyPjIJQCB8FIf8kB2omN+E3+DIeuUhvSrk+gWLm22bRShv75Q5sQMJyIdK1YzVt
/wle+v+eVw9ix74lhosT5xsOAkAJEkwF9cRI8Hy+h15TL9u22OWa4WzQkB1EluAR
/wqJ7a6rSbzLMDaMUvH7U0sf2/XrC+DWv4FYJHn9FKgoIG07zXBL6qDr2lVeXrAt
P/UtWCvZyNvvhpCQp4W6R87InmJf3VvGo61tcwFDEjkraIqa4b8UTF5QX/n7r7z6
6MhzgOjLpE4wRdtizpSm6g0acz1K7+zozpA7jhEcAIh/aOPSTbPpaDb34tXrT11b
vnSsJschc7VG9Zj6SMV9Z3nm5hZxODHUT/nrvqw1pLdyKKafct50obMrruJsV7O6
iH1t1CC7QdfPBBc9jrGV02V5F29jwr1uSJJrkgbqgNz1SwyJjORLWvqxYgqgQJvr
VPzpP/wXECYWDQabhjUjm+gkM27nwyLkmQShT3870K1BLaeYWXRnwpb5Hphcv23y
5r5F+U8SN5X0zqHj7PUDX2v7NQGaDNPDOLsvt+BOwRbNI9vx+bBQQUJI/zCKYfd9
IQOQBVWXNPTly02i+NDqlPTUJ+LzTl5Q2Hfz7o/WUsd8anne/FELdtOnWv1RduQA
HIfQiU8DfAR5iSG7rSMoV+/kSo6ZDPAaDCyWJeoPTjTkzF/JSNdCXHCH3+Lspu06
XFPwvntVUNq/95XMYdzk2NJzn3vH2oVrd80qVzKJU+P/iKS4umeAzbHL9VnmkjeS
vO6PxvJPNpkZRxa0mDM792POltsP4Ldl1eK+RR5diA6ok151vVhRWm9yJ6xryicT
x61RxBvfdgUGelFqG8OLz/GT0NPHJI74BQlpIjPP+/Pn5dAWbxC266xVlKURB/Sv
ZgZVeHGPEu26PgDkoTo1pTdazijbNahWaGkk3A1F/MW89M70xljKSFckDDAfN/rX
Ed3PUhppPHkgrXDLbQPtAd7ruiAq5u0bRFzlmp6ezswkiE5+DubENeYv5mMAcSXd
tBpRFpU2a/9XI8rGVQsCVpCv42J05I1SfrXZ9dsHOg3eftxvFUzvZaBuPCf5wDss
6klf5ROcgWF27GxBdIX3wd4VT0vpkj4pkUIXwyTapDd1xKLYeNaLGahzZSq5xqIb
mMWPX4q6c9VTM1Dqrc1xOk8pkf7APIua2vvDf0BUb8cga8GXYybXKSqfBNTw/uW9
ifYR4f1WpcIPjCSdy+V/n7ncEHYz+f7hP5Pgmx+hD4umHJUb00pu03E2VifYrfDO
EJp1HQKv7r0+bHE24dLon6/aVslsQbGJUvUNXQfEqMGvLhseHrhzFBYg7EUuVUYY
1J5nDO/X84AD6ZHjxhq6UXMLvQNozY14+ziCKb4cYubyMH9P10xI0Poj0vgLbmzT
ycfOzpGbJA2p/nA6WbNFjAMi3txArIwV1dZXtdcwKafoOTQn1F55FBm66ZY+hOfy
hLz4ssMpSG6an0PCGGlRo2nOLaFS9JCZcMh31vguSivx/LZZ7V59Nbsy/6iIETet
z/WiM/Z7WzzRftP1ZA9TcU+eseyw1+dIC5SNv/96Mkr73QqG9LrHAQrN0kExT0hH
WzhVfhD9TfoF/vFc0OF+nGXblzctycquWPWBrYJDQcGQ+ojAvt+4eTDHPRwSNj9s
i1uJ9YaT2+ka9X/mWhA8w3hZjDKxF7zuV/PGKxg4L2gUJ3NFYDhvy4sNPcvU3g2X
PAdJGCgAIXmbLFK/Sz+ENhnogMa1JcjyA901YS6c1OxccCEGWE0dKXJu+xiOFxJL
0lAmAlcxU9U52jiOT/khwHmZs3CbRsL4faDFXTJjmyek1wXgH4XPpLW9RatSqUr5
QgWR80VaSlGjdIZL/4GeMcBxf+GKUs4wf5/mLh3XOaniu4FdGaa1N7cQiXPeHH+X
uUBDOm1qcqdIIIKZ7YK3v6Fo3prdLOAT2iqSJnn7sthc7XsidUGS53i6y2BcPe2t
3ahwQKBlIR3x10BGoQLmR2mNV+Vc/2NGciLHVFKk133Id9btc7AE8/nAsr3pcfk5
rvuSbBDfCI/ECZhMpyLkabjcSuEu9wivys7cyOv0mlfpynjzqSfY80KllQiZsQZ7
kgTWhLPAgItsJ90sG0fN2pn6v7aGg5NElr36yIWaF10S0bzrsCojYZ2bsTmFidbw
K0wohZ2tuxbQd0JyFVlQ7YHDOTT3O6IgQbmtvWyBhZMoUu9P6emCEseDZTo78Ft0
lO1JXuc/LotfCUMXPqg/XNRruaQTcDNvMngyLmx/ZvU/irl4wuGnw00p+80qEfGp
34sBioMeVdtgTIWk5RFp+/sc4PPkkVXZZsrZvc4HdMC7Gwh4meiquWK8JsFvzvvL
teja/VHoLKBXQnCCLvrv7uTpaHAlIZ94lEljm528ImmqF5s4EEhtwm1ihXjqOyTy
EsxApsjWcEFNarJnl2T6BxrTrQYSOsRYFPTsPjChowH9LZq67j7oP6hL7of1NFgJ
yiA92DY7Ud6awMih/MnOg042g+6Yt/f2wyZH06xlEfGJfF9d38nHg7MAhvnxZtMr
MkNO4eQmNnWw6pMv3kU475PzCe2ObsMOo+hb0i+lwXJVLpFvVFe53cegkYv10SAc
M6oZMs7Yxa7vT6TiDz3bFmeCbR1JtFRUYD4j3qyFK5c74mwBnMcLNQw9ZFUvn5yx
g7bID+QBqty2Xsyl2ERdXVaNq0s7RNkXZ274iVaiTdYBs1istrINIOoUZdKN+Auc
anfFLojx9MBCND9htNnfMNAHrPDYvFUfiWQPyyYVJcNdfYWmV9+jh/QCSPMlWoMT
5wh+o1x8yg9CSfwmpQVNxM7CrWYK54p/XhibV5qH2Md9QrkPYJhmxE9EcpPdryHI
Sxe87tzQpIyqwLo5QmTodeLuRn2W6HNkkakhX9RlTIsU93y2wNqaGMHnDaBLAf0V
9o5KTxC12NYlXsDw7Gmp5MQGZoKcTG+968yMCZZy+qw0uMGZYJtl7w7+qlLXLlLG
DkaXheLerdL/Trz2azKy6uyNyjWwL/QxlytMt/LXEE9Lglm4wmI2qxMMly4rRfkT
lMUxvb938A14VZ80mci1V1ic/r2+tHIRcifkeDMHLLP+NDQXKSWRspOpGFWxUlM+
vDPeMWM0sUij3rRSPeRw02LVb32bUB7zatbdwwGDrjs9P3dstcxx/bDfAoBBp96V
oDMxpggrt9MLXwDfb0bXgRr5qOlrPlzblDtJhSB7iVdi22a8a7b9OAAQqovxvdu2
tj/qwvzELEcVBEX240a4tXU8iFEqvfPncN9FAzV2cgt6O0QyejXM0tsN562s1mmr
JG6cAjGNpQ8hqpLskVE64GD3ixPU22YPRPzWum2HpDVbDfsoJKijOTx/wWZwS/aq
SMz+HAheH3y5a6wPH4UbFKcHy8a46czfrq79q4QO+TfuQB9xnFyg5YGMS7zefMYn
UILKEr7T+A0cfdVUv+dJ3KB/fxF9fHnuZvUD5f7VOhEd54+pkW1jWq6sJXJEavuX
MYyaA73KzoHUI/RFDGJpg7ific4AhSu9yAsXjziwiY16/9IN4y5OihE0htRHPven
/nK6SQxO7542sgBIqTTqCC2MaYvodVI7gsMmGS6wwtMXn/Vt1xj4GhbOTQUN95vz
yTCP4gxAt0hveDqFdJRfNFTB3mdA4ppZqByEXBtm6DRjfKLfKSxhcIMChsHqq8hm
dUn/xhBT8NdYKEr05m5fmSiXF447+Toht+KKJeOnjXDHSiRXHUdoxP6Aej9WLcye
GJe9q7XQhpQpqVsOmB3Pdy40Hso785KgE24X1bozJicz3tfS8rPMJobzyEJgPOIg
wyHsD4A5mpNduXdae1ECRIbHEcowUxZQoy+1R5SOU5yUkf9Q7F0vwNF7VNU7AXlu
OjA0WU+4h9eNTnVj/8J39O+Bm7Yn32FgPmA9PnKRyksMSBaqh/x9r/3uEyCxoSYv
sXx0TcvgaDS0hWlDGWj3ZYc1I1Vi/OS7+uWzaWAInutFqLTaYbGlHjHGFyG6QPSh
6MSVIJVymiNx9my43Ecp5SS001YAlw6RPm63bF1HTrM3ViSC64XVRTT4hnWV1eRc
ArqW/tkq60yFZR4/r54CNiwTp+bE7komddi5Wkjy0g9TftuZuZAS8UH1EYDTKMai
9vTqv9n1fV7lacRjC8ci9eJ7BJF6N3v6Mw8NCUg7olJ1y5ERnmxjS6CCfTnXL2cl
mxTcOCufyjG4rnpVHYZM9JEQJ8pGd4yG9vlBaWNWCWxNFOng5J86j/nVTatTo5ki
WtQzlhAGdgbDfrughpScATEZkVTBmL+cen4Ertwa9XmCr0W5mLOXiwJFnrhb5VoS
4OCufa7+0KyHRYv7CVzFLA==
`pragma protect end_protected
