// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:05:34 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
saTFNX7HFj/iZVabhIM2D/LvxxI//9OdBqQ9qt15pJ/94Kckz9EM0lrQN2Wxj00C
yKHVk1mkgUbn5ZDU2BE33H671qYAJktb5+EV3pQFh2CD1O/168l56tYpzjMlpVq5
6cInADanV61A5q57DQ6MQVkHl0XL2APptQly868AS50=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9040)
6czRE7TWxH9MhPgNFd+PubqtR1rGhdQgvb2evnmlEj+/fuQN/oyNLeG6lA99hVMX
56dfpiSe6q4C9PcujIgZmSv26bBYmy9QnLpiELyWytZ9hCP/GMjOLjtFGkBSwxdj
PzhinsKPj7PPgd4a8DpAQtFkJi9uDm68qhHTWREuhYL0LcJBzdqQ/Lvmofq8GpMd
HYS3CCnHHTuROaHt+UvGmEH/Z7gg5vhvkgoKTCSDiLq6Ov9CLDlBbNbjtWREakDO
FobjOo7cQBEIS5Ik2LqqEpJVge/G8SOYPg3aWAlyeDSFLS3vpcY8S4icDCZyGBPU
ifb+bfNEHDlNHJinia0Q1HiV+tYU22gDIunheFSHckKVx9Nxw16oDxyPESxajJr2
RTaRwzgYCTC88TrANfmpwhfumH70C8g/X+sATlERrtkbWPUVcYXUYrrResUB4Z8E
6q34Yvt3AoJMk7/kObUuKzBCifY+VoBvYSkHjqDCPdiKAegCR0CaAoTC4RmtzfiB
01JhDtjd3A/DlJNPfk6UDeML+NxSrlI8yyWaB24D8B6GZkws/rAcoa+tsF9IzNrG
g65LNhyCEOxfTZ/3c6olGaXC3HFjY8a+uj+PsOFjYbIrXf73ngtQHJ1e7HwQuYCB
dPrEMCiz0xgiw2+2eIwD/lNN/Oy9kTmc9m0kiuIyFu79TPy8B9Yq6rgmb8AJDZZn
Yhh9vnW1NaYALWlsmAryWO1FluCZuy0TNiLoQO0CNHHzs/DZx2e4ouAZINsRpPxN
rrIWj6JRKKSre+ap6higxOVzVZTqFiZEzCMo0nHrOVpRh08cTDoI02NwhPZQKCQZ
C1BjA5zetqFCr+wjowA22LB6rb7PFEK5L+5haZLt/pB+txGQdpeMsK/t7bMQFHh2
2g0hmW24dw7BG2NFifHB/98dxn8U9rG8FLCuP5se5PIWKJdwdYfIn8bUJ9gwdTxz
oIkf6nYs71hha46F2HKaKsDDaq92auH+Tti1kUbsa0xAucegVnj2MNU0/fckFxP9
GSvzomTr1aRRNphdNxxSh2FLH1wOVVcv5kSR7/4KUpJDQYSYMEfHu80mW9UwPksA
2G3fODPPuzEfjJYp1nZ0vnVfNTmKmgvhTGRSDfKOjIwPsHnFb+A5AxsAJ2fcT1eb
hOPwFdIEoNm+SQSyFMiq6AbWy6FQEC49aGNcNzNZNKyanGyMwrBAFJZXech9+UsG
Opk7ylhf9hx6wUyrwdxXfZclLdMxRmP3iLwmTBfnywNyhS9w6TBFL8Is0VYogls1
zuUzoMN7wx7P6GEuGN2RmXEeF4AIsCDMZQekk3xKHxMz5RvZJN8bw1RF5RD5RGGG
T6sZT4qNTxi6hFoT6VkE0kjdxj/4AJzp++BGPzc1Zha5SrBZagSmIVtMvQsgyIxX
ZFIfW8fsmk9kyFFlyKPJQPnjbOMgM8TqY8MKcvpD6gWnWXapp2zES9QBf/xMkt1P
GKwfz80kE57JsepYwgjHPD1byoAfHR8vmjrmRKnLt/Ar856FhVBMKaCdGg9Ey+p2
0LlIIOMtHRsuPEkjQsGQCXA4dVdmjI9KgbdB5v1rVQsaiigzaJRpEsUJFyop3Wl8
T5YazRyq7nYX5u7ixCToSju4OeHp7qhLXi3gO3pJIsp+ZkWECqYDr+nIrIrRGR9n
JlXiDIhLJgjEzw0epHlYhaMREwMPLPDWUbu68EWh/R+vRXKVOAvgRqcWrGQBA9kO
QiXGwFLIMoOTA6dzBY0Ogo5cUrIEG+VqrcvBBQMgOrNsVlj3ivBfuxREnSROnTqV
UW1pDKKL+BVcaQTeNONPakKWiGsaHD5r1MQhq9FMwJ7s11qibGDei2xTEVDnw8Hi
tTSJIGspOWMD7D3KlNFhgpm5QMRtIXExdr1uwgyxdeSOr7XJywRMrZ6Sj34vR2KY
E2XOPueFDKU97xqwEv5E1v7l32YWMI9e2I8d6LZM77T7fykplOrFTCaSS4k3pf//
G68HkzRw0jE2mNAbxWXAmr/5vyVdpZXSEWIGVD4SI3Al3u9W4JTjZTn6N++u4Pof
pj9Mz+t/9/qazXvNck4ARMVZh4W3emhim8LL/UAnuf2IzA/JVAhGOx+CU/Ztl/C1
6zNZSZqQeY+7kav+h0yilpY2LtoEqW+tYVxk7n7TVxRSkl37qthMKRlMOlC3J9QN
ijgnYkGAtvANFBly4Kl7nAgkM5n94ETuqVv/ejLV/CR7AEIb9FQXA+6tQKs74h9O
hgYt1yTq90wFFZH66DA7Yws73Zh0HHD5nBYjN1N4/Ipt4jjxZgLB2jSucFIhH5jp
j6tDTJny1BoSkY2phc7FloqR+WmRyTDrT6ZnXgsVHPvQMLumMMoAtbBPmYiJeZSd
mAGvCp1Lr9dojNHI+5vX69XGrzGHfUH04qoaApw/uCE5DIZIeMOYlMBy+0xfOgOV
cXsyii5gsa585Z1y3cwHvepNNcqIZKukdW4+B/F+o4tWfFohei3pd5da0zBj6HO6
mXHVyZcnclbWHyliI5JqhEFmOaKpqYB2FidlCDJmLWyTxvXLgktDUQ8Schah1rcR
xyrbJYEqMnKmDhhtAPfJDiPuYWp8DbmzRjFdAoNj0BM57ajokI6DOp9r5mxwMcOE
zL8bgm+5QZH98nHa6SU0KbPILz/m51X8shkTXL/aNjQpd3vb6yFrJa0aUyW6GRrQ
UPSkM4qTLGnP4/GOVKdqB0satazYBJbqMa8djyUqyVT45JSzUKWlzWyKaN7xbRP9
PSUV4hxJqNIyLj60UjaXS67sTESovr1lbk2oYHPH7AhB4xg6/wZRnMMW+sQb1CPs
TTWtx788iCyInG+ByYb5bO6YKhlUNNxttNzlFQRldp6+Q3v6IaWwlian70ft66tz
RsOE6NPlk8naBmjhWn0F9qIijMHeYzRdt/QV/z9SoHKmjOsLkpR8m+x9BYrrES1b
6fPi8uufFBffezffjYjy81EaVdSLrUpwTlz9/8asdIXI/e9CTnJX4zaPK6gOYzL6
6+riKXpgsHD1Zxw703QKv3n5t8dJ1gqlqapGjEzdSsn6n7u7zsGGkqfbbLnrWNPE
n6l6JHUQUKuCNyp+FUnbnRLNNOTy69FGaIpBSxjaTFRJp7VbBJp6vJygrN369MRK
BG5xqRHhEe4VsVo/8fbc6WKwBu8wjdYaGhJDC7bFWXoLGfgx9XJBILqF+lhz7+KQ
NygPzCo70NiIHqcl4LaaKabsC2+myl1scwralX4leigXcKsI9tUw3fWnRpRicHW+
q+/RBRLwmFSS+V7EDtfGE3Rcl5hbF/INg2WxlkzhD6hiWeiow4XO/9ofocvVgcuj
n3Koaxl4+XolFajn7r/7jOZFokocp9KRRUlrmykt5UrcUY5J7OiXdO29UZzekKMR
b2CnRU6c+7W0jBC4xmdoy4CwKNv/3fCzKnI3TQararyrfwKWySMnw02rAtue209q
paws/VvWoNNuxhvP9AyUK0pwJdnOJzOsTQazdAkK9XQC0hXI6QHPK5Fp1IHccmqk
1JAMQ3a0MIZXamu4V9/3SK2acDxlsNBDGiLQr2jf4q67D5u9EU4sCz3EthDQOl8O
q6WMsL9UZpnzAecwgo9BBe+EoRWbn65ZoEqx8J+4WjIqJMS5eMPyOyzZW5efa2R3
wCXaL1hQpmHQyboKeSf06M2VuYKlL9Px+wvxAJbCCUJKZwEhcK3aQpDJFn8AVT3O
kdslQuwmja5MeOY/C/UPS44n8RobkbDW7bY/+Ra/BEUij5fR6ytFkubLunZQ0ZOr
KAza0WC8pjbegTKbzG/hI0DGqteWis82cqdUZTS8YoREyEvIiJNvKcK4dMFsrnyp
jTx572DA9aADX7Hs8ZFvgKji77wOEgB+L6f8RGtpdTcPdYFJlGVDxxznE+AQf+d5
O0gTzgDPV6cROi061GgkMK0+okUvB3+9LmDSFqzCfTPTPx5PDJzqGbQpCCxVHPt2
6DJ8zXuBGOPcbZOW2wM0Ce64FukURCZmADuACC/bxv1Nzzt9GxuRD8nxU5bYpq8b
fYKHHduRKBNZS1QpAxd22eJ771H2EoDtSo8Em2qw80NaUDvLFzbiFrB0+SSoqWZF
ZYb0cMJJv+KrxDOUQ81vH/w9CdOyOTp1wWhEPUMVba0kVGQtJyzAWUEnzi4XxjpL
BBxdaRMe44JpUj+ZZKaHsHgwGjz9TpudQGZrITzz8DVH95k07ScDUJPdB7/zqs50
IklUc9dRM95oBzQTVfIYG+JGyNEyRlaDiClH/YNXqV3wxS1RVOF6bC+7+2UWRdzE
aUktoS1BnSMsuXvHiUNgKhGgTAmEbvUUAgDOM2pmmu+8MCzgGIug04tE3sSIa7Pb
UiOpzieEnbbAV5sCK0wUFQ/wr4n42rHBZaTZAKpvD+mj1rlHOqwwhBPT7aX527fZ
ZfzEPX7mLGn6IPIVBTRnqnx00SjgSLIICCKhS6behH4j6b0kbwNeJ68dbIUaJMzv
ConVhHax4zcGpLnzS1vYoCwwfsoXs6FAHvC8PlRT0IoRiqkD32lqDrSUJVTh4hfe
J37X2G51+aVIEcewatp0DFcij5kwXJRr4PPWAv62fqCvN+Og0VIfPPOstG8Bhs3Y
nA3tC7rfKhhpW4zryHuVcXBIqfUcjiBH7eNVU+BEijrjzg7s3kEEMhJUw5c4EhCQ
jJrOQGPZFKV6LntBMYOgoU6FOrb/OfveFQZuwCSSV66ERbvPCAjQ0CIxLbFZTL+l
1DBpb1oPcCV6iFNCfbpEJKSc2gV7QO6xOjzfEcNz2i2ifuz5nTQUTHKEbIDS9Bwj
YySJntuLr8b99EHeC5NQMOoWFgdw+xZ119MQnQkE+IlNq/Zr5NmRFLCAEIniN49l
iTcPCf9qRfcxUWS+zHb1REMygWotnsxKzEJoL4iJUOAtf4NWuxsVJSLtjDXrzLs3
eFjk089GWsETdEe347tFxI73Qx1tlDvJF1aJIfqxkVk5ueCRArbrND41MKbcjg7F
hAR4wfjXtPFOwy6hldp3+gSkWmyNvVmtdpm31sZtcidlIJIX2kX7KyCo2Dv9Qw9X
XlCAyLV1xcdxPhCqxP6L+Xk5RrFPOdHZjoDyPsHLcbqyGhIQbyqbdWe6ZeZ/YWHP
sv4wzAxlHXJdm3HmHONp1jlvKVSOSFlo1ODHLs6+yW0dMun8u0u85uVGavpuV2+C
kaP08MTgiAM5kZwk+UaibH345guhsvf9+YFTpKHY1zoKInwBi0OVpfpjjxAQ/BKc
7caHgaCa/DZSsQpEjsBNLWh/z1iI06dSHjtZHVgKr/kfpY2cP1hUe+BxK79HlMDn
QzIMZiwCjTWWn4fxHiNyJvZ3kVEA3xzBbyvtIErdXczfPkSAfmXpIEiFSXDLwxRh
rycmvIIhpi+0jVYX1G2Ey5B3z8vXuOJSTnb6yUyuP5TBjbBui80EZLBjv1pmhPvf
WJIGt/bDKaMRR/xbTV7+sE6DHDiFlZze4tPlG9RLicl6/YZWXvp6qLibDoeCenjR
GpaifolYeB1R+Nq0I6C3UZRwg0xqUVu0VuUr1Y3nXmnw7W04J+mHPLGdkun7lWoQ
EmnMmFt9qCQ7WK6mI9fFIyF7vt7DoqH5UCFADn7OEeVNZp24gqLvC5D9FNMVRhNb
Gc0OWr0CPU0xVvGjseW8XbrgMwDoCj9oj75BCV2BDE6cgfT0k1JKCYvmwqTFus9m
tLw529f9C5SV62Vci+WCorZS02HaiaYlj5ATrUCdFnKwfeQwz2AYzxTckOzeaNaf
1skvBBR9UrSDDxjNe70Q+5fd1TxdhdTNpz1QCUQ1aRPbhEGyQMa0Qk4/ripKyiYG
dAadBxlDmnQqsoJn5JvFSvSUgxfiTO0wbfL9YGpTs4ufdK1U9Lsf9DC68I9KvQmu
opLo8OfLxrPwXltzfyFd59K2aFI7qw51NxejIEBLlIh/03JfwovPKoL41w4wT6Jc
Xzxo/YW2OtqItIg0XqI+7T+E/16iQIV5bGpJDOHCAmYTAtljgdzTVb/35TX6yXRM
pXQgReSHpM/mE6U9bgwR/GIUi/K0cIzLHCu8aODk9SQYeymw4TOI+ogK6XXg/MQR
tk+FaEhXdU9FwAqE0MQocOCBQASGAc4+zIC9VbuJS5r8W1mP5U3zKX6C5Dpnsj0D
mNoUxf//kPD/i+rqJta8Aus4IKU3Jz0O3dWIBqv1EP0pmoKMKLYeLMJKqX9v3srx
lG06SWezzJEfXYpnCxcb4QE4z7x6dXbW+jHUUKg+ZPjisbo72EnXrdFF9IwvLtGs
vt4vCF78kuGyUyQChgussN4mQ2/71/Nml6XTP/42+upImfUeC22L05f0td/GTjVd
h42d1/V9RZDQ128XCVDdhDRsTclWL89ZSnPwAESexnnXjpqzuVllwfDlDZGJC5sh
Jnx6jpfCN20EYM2qAimb0HZUmrpwft8hc2g+uMWTCFgGZpPRqQKS+Y8IpcKOGho3
giYZOc96EgSMf287xbePa14Uu4FO+/faQ7mAqFYh80NLzy2peF7TkdogVxCbxWql
Uhai0QPxeh9cG1S99A0wLln7AE2b6SezNVsYl/wTbYIU/8b9e3BF3I7hE6V/YTbg
Zc5Bc/D1YMoFAFPkZ2NDefySx+Vb+OypZ/yZzeaj+7zqOJhfYf2VeMOdFCxhoaya
xMYEbNcsVS/DbCt5dDvhrTHfttCZG8+Q7latA9TMbZYEYHbfTuKlpsQQVBymHRAS
LiU0N+pbgkIXf+xIM3K0zRr0hrAkGfHNGCXN5RqIpvp5+gTjhrMRiPyFKvzbonMf
eODw4iwCzZtkKMLc1s/UfM9u9XVfGYiJQTj5//rhENtwnTSjW5qolI0GtWCyp3wJ
g8RoaLzPOZX1LI5+shdPWaP+h3QgIgegO3qITX8AMammIN2bK53l3HvYs5wV2qok
zDa/fLiFKuOdg3fR64Iu1F5hERYdppwv9hz1Dqv2euK/wnZuCufYEGole8XZHRiu
DuibFerC013xUguW/ws8kKGcU3Q5vOyN80Ii/Rw4kkXGFtjqsyPtmMyH+rqpM5RN
8kWkNTP/NYtTIpom5tGff7jBTLLlA0m55NLTZgO73QLaONbZ/Ou6ZR+4tTcXl7AQ
HbvvfUoglfuacGIImHxXHm4PFrmPl2BdHVH30AAySrUzOa2pnIxHCk2dEouSIiqc
ntHi5Vml2yGpCos6ROTQNDlXYp5C8Q4G7i9KfQDyMKycgNxmWcVRX1a59J/OtPO5
SvdXPqjN49lTWRlfjQVVmyNL6Un62nn5OKXbDt5rdsRZ5Ub5WnW2CJiSpLi88CJh
GuJJkJmpbs8POWi28PGdBYbGXj6BsnCI/MajIFVGPu1h0ViMjeteg9O8TsTNEYU7
s4UXg1ulVWspvb84n0vXR23ZLXA3MRVlRADB1cEJ6lyuFVYN2icthj2bXl0AG5S6
xRsxV3mZCglzVzgIo/sw1CP42HoeJwCfZOj9LzcJV1+BLAI5vsJIp5QpAG+T7n3k
k4dXJJY1x/uyS+h/kBl2lulzU6HE/zMgopYLU2SCON3yj5Hldl3ojxGjAfPfsrA/
KtUapWdNDsLwIMKrzCjjvF30z5qK+fMfuJC5I9wWpPTA0UlLx9a/1oDphXm6LGe2
Q3yDzRb3AVAClk9+HBBi02nmNVrOtCX6Uj0KQgnV2VP7Tg/2LSY62MiEsxVmQbWh
8cpxlCeY1n398TYq8QmXZZyVrrSWj0J7nlK/MChnmuulZzXe87sMbgwRpVwJIPWg
EhWY8hYcYLYJxzAP1X/ekLe9TEw/Wu/8wKgdA2flYkUtXtmX05eaTfN470RvB6m1
hl2C+UuZO6O5iBPjdY+1xgsQO8rIHqmuPiAI+9xFD6wK0tRPl5CNFTHqy/9mmIaC
iBVS0HIkGNvWOS8WM94dScHIgo5mXjsjn6yNzZJ+0WJLN3HzGjHFAsKlcLIkDUqf
UEvjvuajXheF1dUPGbw0nBKglWcNFRxZqu+cR0++ixLNaKW9+EjHT4LM0e+bWWmy
5gqKh2aktUYJZuy0WSoNrgJSdhoMpuEVtcyMF42i9sH7XBZArT8Zf9CxXeLMEDpn
UrFAX0PMZ+qabyQq0nLdalDvMUFAwRu1l1OmOXLNmrGPvTDLY+Nc8tYtjPLgRg53
JpejCeGnsDwCOgsr+7RSRzNVjOlp60MwEV6u9QB1IiFZyR0eCC5SLFlcJ2UCNoBj
YRnW3Ps/VLkyVOrrmbwU1+PzkLEWU1YFXehHmU5LPZ/tQbbQM8GCzp9SyAsIks9I
nHqRPdQm22UrPgzzS2AooCMiXf9o4zgbhMbYe40yOHqgVdR2D8ahFSdbqS+mKhM7
m69FQG1LAndOARNPrn30aUlBDWB8TTpSnHpGbp6NaAQbQ4wwR4mVOg0bpDjcMQwV
r+Ld1+w1dA3gPkXKl164MaHuVzaqxvNcOaYcIc1376Ii+eo7jZGbOLHHXosFXa3E
XywBYWgkc8F6yovE/zT00VWPxf33uWs7tCMiAWwrbeowEFJ0IjXiin6etI8iQOzN
Cat5cz/xXpE+IHqOVt+c1ZoWR+YTeOZN2rWqivmw+rd3uZ2vfge0R/aMuy8CJRX7
R8sGSqyC+2lxDdE6WXFkrFpb36L2moltLAjJc1BQ/XnmGx59t1ZYJZ8LKVZj4S9t
F6WB2SGsS6DmuqAYD4CJTMHw6cBKjKlo4+YI67WN0jpH/5Svgl8sHVUueErgctkr
wfF9whc3+lqGDAAsB7BTj84MtTAOlXrt1PJH6q7f5tIaCBXKq1PbO60u3xAiS7Z2
6kxspCqQS4QIJnhRXSKCrZsFW6cD1JKhVLJPMyAts1VO7N7t/Nso7v5f0xINVerq
6smM3supB1vt9E9dSLYAL1nhUp9BiP7M7b3AomROUiFLK9z0KLTS5hPF5R4YaFF/
B44B4zSflARgcX5gGss9EzWb6+R26Qle5nIeMjaozbVKNyAlj5hgKa+itt1doIli
pjJiTRl+duiEaxkZs+d8qKVPSyVK5wQSgTYRYKrc0CCdsnpad8g9ExABnmA6mNLS
A68OlBktC79emBaQuozZ0VrRMzCnyfIh0Ginm8VORsa1PfrALd/ErUjcCmsLBuK6
KESN3LF8QOBKqc+hKMsPwC8GpGIB5TPm5+28L6Fzt5/mE/kvPO37rWdvwRKraK9E
N5sNWjhxUsq/VNvdD/zVLMsJu3/R4UaUuK6smyLKdUZJIsP+9xY398EjYW/1LBx4
IFzWFxm4edmBtLpF0dRU88JrI3no6nF3aqrQ9oDYsUCyPKiE3MQwUwSGT1WOWAWj
EuZOm05P4kt6gnM1fkh54spSNV3HUpZ+K13jmCYsp3fGatfiOE0f2xLtotyxBakc
EW4Vy6i1yiGhVaLAYL5g1LdOcKCBfhMuAKEYJIqlCF/oaUYmbsVx1XO5VKg03cut
e297/H4FdSIH3fh3NrjfXPbUmOdEPcLEndg9bWRq13fdnZw6QAxVTV8q17dSHd1E
yQyW2CdQFJrSb8559OGGBiR2M/ByiBeTKyCq8eiq6MoZqlN09LTDM97HsJz1siSf
rje/71a0uTKLBytvC2seLcjvat2cziQda7hjkHByjKvAK/LMQxhPrCRFiLnNKULx
jHqdWGkd4hSRV9gl4z27svo8h2K9ON4gss0WD9Uk3XXY6z3M73RsZUJ0X2GihUW/
TV+TsdHQAEF33Z8SCF9IDehBvkv9iG4q28SK30jpSybQY/n60Vz6Da20jkuYAo85
D7UMHD+S/RLo+/UoEbh8icNsAIxH17QPhM4GoF/B3kbvvXOclkA69Q7aFKChWFV7
MSvNH9kbZOYVsbBUifcYU3wj8ESy87y4pf6kH+MV8Sf/IIcO8pmo7imMhKgsgBUO
sXJcZS59E6QcYS2dlpOOnuEYOPXQ/OPVIxZE+70/ylljUSPWbjIFetZWAmrGE+P2
A9Scmiso3ynqsfJ+xtu61N3Hw4+XlhRcgo9+365JMGM+xU12IRpEu2AA0pEIF7sX
lYIuWEF4fZWtoO4pJnsAruLVFrik58nMuNi/8+6EMScaSOb8/Fv2Bd2jA7ZoUx2/
XQzcPbfVuBbqpOu0Gn3A9yAv6puA2pVWcwBG61qGNpn/EbPH+yzA7CdW5leqat4z
4QuoBMJkeJhXVUGpZwpUya0rTEVLEPt5jSoq3CVr81pOkh23lEqQ+mNW9tNK52XG
hqp2n+jH057AbTLtgkUeCy5gHIXJ6Vm5Zs7FY/L/dSdtB7LNcBHfm6pXG0IfD5Dq
3nxpVWp3o1negaCCA2ZNHjwGJJIL7z82uf+PwQNtY3MVBpl1kXWPCwMVUMi0aXu3
BzZeofkL9CblGObxIMfixi06ZixKPXuhHLGa/ppJ2cxytT8Scw/KycHX3WXu4+5A
YoJ2T6Y01NB/+gA0eIs/Go5hyiWgancLIeZNr/ZAeEhMbarY0QSOC7DDRA6HrdaW
bzWhmfis5uaTQ+7I3KbNELfU9vmDrGgQ7OrOLKhoa77XAxpYzFyLhd6i6PER+V51
Q0TahRTg/ztjUaQvT+OOKrG4FBVlJEPkttO7IgNHbJIYUYBptHvKMQoC9Q2ToLYj
9mJBVfvXc9u+yEwt9B4M7d8DYIWP/3MMuGA/G9mIxS5Je10yzD2Wbv1Hw1uZpJi0
hCV1rvuKUE/rOosSTDWI7Xl43Pvjd1YjW3F3ALqjnkjCybr1c6nHtEJYLMafEA5N
2CpaX60hCMntmYva3txfz6fZj6SSo/uBeh79Up/kxeVRIsbcQJGy0enCjRydEjVf
WWmAmFKx2LnqPr+FbAqwv4SbEaHt5KSDEU9fL2i4v/aJTJAmpoR10sk6niXaPbLO
R707p3DtlFmgE9VELb/pl2qb5WYjGeCdfpY3ssGDfX1Kqq+12hpnbEuuk5PnWhjv
NLElT+s2zYybgLTb7Hdfbg2XrctxlVzsaOKLrhzRWGVybH5nGKswrbji7m3q0E1M
ApGJln3gruqynMI/ggCZE2mkyY8KPpNmJyuihQFXgk5Pj2U1tYlhvv5HL+fsWLXV
Iod+D0fYX9WUxKJ0Gu4WRZbMVCG3o58BblF8oHExdtYKxzpL75dmHGfaIINA33mQ
wZl0QLuVMVCOghmhPs/yihcr9rGdB5TMu90ED4viBE5VHKVRgH9Fjf4Y02wmWMGp
uT99+6rqrd/OgFqyjth/lt3XyiroCFFkjye/95BoXfCnB0ZhacxXcARdM3VmX2CP
H8XghJADxGhAqA8H1kg+viadfJ6J8oGXxcE1JCp5T5aylPPUur6ukQwi+/Xk19g4
7rQT/NEEPCWw2jZhSAtaoeckYGtxutKQlnLP5EvU+D0SXIaKOKyPqWKkaGjCpQlo
v/RBE/ESqWYBfinx+atmlUyLp5iFrvlbko60MAXG6Vs8/aRpNm8+FtWjkF5w4Ejf
n4L1YWlGbuC4qVFwCwE2ZVWKvx6K2g8mISVTgNixXjrxYmrGewUOd9becVr1bzf3
wpBbY3gA4gk2TSYZC+WvMq0L24aDRRDmF89HBQLuC7a1L+XmdY6dD6SURhKUKmIt
kh+3+l9VxsyF6iPFTmjJuiDPOrz9qZjYbTZ0N3IqKHKRX4uUTdPQW2QqO3BE9ymR
KQGjoM6cyQdkXdAh/butPFh04Gv6vdwRv96PUQygMFSK7JoKMKBCAS31uOEESgAP
h0EyO7nEUKEG3Egxa5nBSbaNB3FsvmgVFakEA+B6Bc8acZUU3n/VsJIk1AuY6VTk
OLgh1F5CEfKW48fKlLKuInn2Ex1yPlrwq7EJEt3Z1OR4RyjjUIKn7d9o1bjur80i
UnQqFsZ4YieevtzPFrBrDOKV8T++9ZgwMHAd57GsRmPBs6tuz3n/Bfbwm+yCPJiB
HvorrgENdG+zoeiJTbl5gurb684nZdWJQAxmCbtEBZL68CO+EIM1qZE0aByuBpcX
JQ6ifPGH75Wk+wUHgcbMYvJCCup+54z2xhIZ02xDzC+AEYkqBT6iDSgf2rcxwN16
HnNgLVbmSGdJ3eULXob+a2jLMs4XiIBKnwLwv4+uKy37yZEHUuoZzU3fm5Wj7MOR
OkHgja31rvaq9dUaJRcg7Q==
`pragma protect end_protected
