// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 13:57:45 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
izMn0zp3B1LFBqOKfiud5BUY9gixLT+P5oicwYxtav0A3lhQfQeyJsZ+EYfP7nb/
4XPHzM6NnJTDfmkzkvI0o93Uqt8fT8Ur5jfmtRaEpbhJo3bZz8BPEW7rxj3fGBw/
xkPaMqlWV98TuBjGqymzfeN47yuDVp7vzhZYpdctTxA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 35392)
FMmrKq+Cg6tZQ5y7MuATiCjFfUE+0i7LJSaRLV09qmxbbLN0EzVKCpZTuGR2GUfd
t/g2I5vWtMDJxUNt6hMRbrSbxV+wU72dT4DoaXGDgQ96bflD/3f9HzbHfXOcTjVi
30l5tpZWtaKTHbxlo3UgZDKk64MUY97+wBpLXfaA6sq1nDjxscf1T4tZELkSpaAe
2dfoCqS9JyLC6j9ViUWbYyxb/RO6rRBLufLffVVzvPI60vqM8w9sPldgJkkl+Uqx
IGlOmbl8eEyKLl8K7MwM4MIyAHN0+Y6JqTBsINqpRN615sCKGhGfCXwNKw1hu3Ga
Drf2Y6hCHl2oniPvtsxSrkI3k9q9iBW0x71zAhinQ5fhK659hjU7DHPPuQCUb9I8
WumSRGL7q+Rb6PEWXLEAiYyinA7bOspJQoPbJFB9cQ5wQwxdMewNwfiGAy7C60oF
XrCD4DMabe/5cnQDsE9SbP26gBt+VaWNMw0KwNNu0HHCOP+W2+YSf6bDIUD4ciPa
S+g3U0/j9WaraeLf3BlGmdc0MExxagqJnqr+SCwLQvsoh8zVWBPmLb81yjc+933H
6ISDP2r+GzyeuLk7rY1Ah8ydRtWQ/Toh/dBvgF9TaE2vpanwNEw7G/MTzqU02jt9
/++9hqfhCFgpZbnO2mg53YEcAIxPRVpoOslRV3sqgcOOsX7xYcr9U1CDu/65VRDW
aPY4wT5ZRBbVH/7r/RIQmaNb3nZVM3ibNwO1G+zSTlQO07NhAZDfaHiqk3hK9I4o
2dlDG+Z1LgKqnmztbVqEJM7BE9JP75+oa0YwC/NHCR0G7PU/Wb1ZWZOr0LKHJc6f
zCv8cOZ0Ab8ruvEBfmnPoehe9gF+jw1Ejh2BPWwTXKpnWedV/yb41NyGCcAO77p3
jGabMDEpzraz1Yep3h1y/lba0t9dx1rWN2EzF4g70xSxoJxmASAUQgvXu6Qwhtil
nm68esH4XcmZQtNBJ1tGdJm+d8hAwN9ZXTIza9d8o1IWNPZI0CyOrln8ZCabgF7w
ZqD0BxrOTcvaYQVX4NfAWuLwQMXtEPjZC3EZOmEZ821qe/azSxNHX0iYLY8fBgMW
rYKz+3wcoAdjCg6mXLeKtq6gVQw8YVB2x0/55f27JjaSt9JTUAmmBUDMWKDHYDHO
ZzFhDeBiSafLMBUOc/fG7QxHWbqRu7OH6WHKCq73SrtzvKKSW9eWWykuG3mVM/Sf
KT1z3wUeW0qmiQZ/bnPvMOr2gauzCyTfFssgHpl8U7vxXV2x8dqAhRch8aL7guUJ
IJEl+tl+R8v7qz0B0MKRe82/Gr3jSw5Ar89zl4HZDs4LpxM0QyC8gffE9bBs6jep
t96ZHpBxRYM4E5N4ovI1hRVTQi7YkfM47r2ev0YPiiYf8P0lfB+xB8SrZMCyBTyW
lI6xoIQomqXlht5WPJITSBr9RAsx2ARwVWs2CzyhtHV2wGIF7T1lQX0lgMkLYS0f
FEoKzkhaO7yYI30VeHrzTWesKCAYyV51LDjy4B83Ct0lIf55iIeTvO/b9IHyKks9
Qlu1dloJhurne0TCVWrEjU8DQCcazrBKpgcQ59oRAmfK2vXM/3Cnc3o7jWIhB8JE
iUbwHJCtHPiR+eiv3yC+NpQZ8WJTTI0GM1XR0+fVEurpfaT88BcPpJYqzKYKUH2n
b5IhAPIj61/5n1xQJLcpteu4FLlIwUjeS23E39C4VJztk7ZfU5S19+BtKSk0yKBe
IZYSusIlJNcyeXu0wxzBEuAbXGS5i4OmgdU2gnFqajRfiqa8IhdheoggDWLYei4Q
tOxKqb6NlSvtOOwkBJ2Wu2F9UP5I3aS2tMejU9fPAu1ZGwTGtWeEMIGSePAECaV5
S/CEtQ9PMfFZbrXV2jplGV2QJ+mQKCfuEKzvhN2LUYK3xge5X8vYpTvD36Ov8SZs
AmDuONfl6mL8SqqqkGnAka6yh9rp285TuRJ+6B7L75AXogLIErYUqojWJQIhoPvc
oidq2Mwg6wUehEN18tNiq35vrdOhLhUNA/907i6ck2tGwYJ2sxUL/ccsb/UbUiNR
PcJHf/o50fX1Yoz2GU3PDkkl9BWxdamTsxdNsks9t50xEh0QXgYVkcPxWjbXt6dK
SeGK1QpxXiYIPt++lgSA3xrIahFhKzVo580byClpV523LDjHwKbE8MCv9T8zsgNk
BWWSom0F5qJlOa9xBKE03LP1wibyts2EI1TBWegprvq6wnq4OC95QeeyZmNnAMp4
Op278D0hxZgWWQ+gtHP58kcIEFYNK6XxcFby0E73IC4G2yCKTamcCZJBWKTrpOVj
jLvNDoStP2UcXVDd6QRX+cI9g355ChIG3M/9jgKckhCY2mV07U2LTKuckYmuITuc
d5LdtGTZDkMqlxI7Jvp9Au2XnlvenRFf4ZYH6xnAmPPXyzs7sRT1CeIS+TelXn+E
pXtHBhdlacaEb7Vc4oQHujMeWjuPatVhzQxRZfCA8RaKa7CA/1EyGtOrCkhg77DT
xCvpexRQOv+i+nifDzfRrdJKdGDYQNPcY161DrA7nhIPkqWajiJdUTnYv012/5Ul
WMRTtGFBHfVKOgpJKAgvOgxEGx1M7Hz7wZ9RGV/x6LVlUx++5ts4GwDRzycCdpIx
8MX3xhqFlVgWmdyjIn+PY4dNNxIGve/BhCQOyrRyK+JzqqgHYX/t2Vx8MZP5Fnp3
n8xIIOj0Ius3IBuMJMeQymSe++Z9k0y3vdUpuaR0gHiYFgA55Pspm5qDugd2zwB1
ECFpJFUTp5SbT8FvwHbSoaYF6IzIcGkZdoI3OKvp4OFRHmesz+PMSRZNC6/nrAbh
RpZKqkInH4pkKkEok3OjuTL4J6TZbkroS6WxFZywd2zaWPVnVPUEpYV3xwSk1STh
q3qUeyq4f4B7E48Yhcb+xE9a4RO1Pj45qTEtYTooklGZHeuaBIbVunVkksPHf8qb
8lTH+BF+2kWY9Wi82pFKJE1qq9ynO47jWeMUwjmHuhHHilsfKq1DKbNrN5XCXkI1
s5eIZ8h0GqCn1vbySOPB6Dpp0hyRoVAl83cT431g38dksFoO69bPZ4w1ZzA8ppd6
iy9vYNrTNCRDT1EUZWiZ5PWR/eEam2uvU2Py6oZJJQcrg/JpHEsSc7h8SMl7Q8Qt
7M8DGM9G1Hdo5hHBmhg0/WbMryeOjBTHe4oI94SpuJZYHrwI2jVMd+uyBjmJwUxH
chEf9XQUF2tc1GW9bxTmVx2hpBUyOOPioOXGNYmtkoosvEtNBz2VRa8NFIPOH0SM
1mojSG+fBpJBdTam7tW5oOdKlZlMekt0RUwSmiDP0fE2nxDwzji4nFtugUhE+Up3
MrmEwcoTDuYmGVu02WsI+rChNGAhVmIOGIqC5MXRWASSjG+iSb+u0KV1oHntZUwi
s5POusq2OHWf4FRGpN/vCa1pPEJ89SqKaQeuWf5Oe4Cvg8XvswyXH+7JKpZsTLkf
0aIjQ8NkqZzHuYDa0y8kOCA6vX79KoSilEYrwmho1XzTFbx1cAVQ4MZUQJh9icfF
mFPn/RKjTvT0FA66vH+p1G7RFmuIaoO0tygh4wZWUrkYEkXcg7ftK/G9RGUpV29Y
jQHIEUjra48zXeVve7Mizuk1UQOahP6zRtr19/oC0ZpXYFFuuEa0Rn0QNkWKYxpv
E7XJSx6XmBf8sHUlNWKdMN+m6/1A33zCI1FA4ZV9jryz7rXRyAfP/O45PEkk+mVT
r8qCYPYPKz6Z2hZWeUuYwwcuRaT29hRo91DPNtuWsucCFw8ic9sX+gn2udiMijmZ
VERdqeC9YfPnVOeyNCLYo+iO5r3+9aUfwlw6HTZ+CLDYjCzrPskeD2fWjMYdO57t
vi4LSE38Oh7E/gHNs0qZ+4omDZToFPoWSAFv3aIVsrb9E1NUqElQtCOJh8L7bVCI
AEcBDYIG26K4UPUavhw3h6GzVvzNgQ3XWG7T0S/DrdFaZnat9trPJUi78UCpecJW
jJKW6cG84G7pjOK6giPQiaOtFA32YEaKw+C4f/Deg3hBMyFP5rtriDc9rRauZLPU
r3zLCQCQcTBI8F9jr4IfoDn5MKDSYrSfNbQKLXQOD3ppIvHWhlv/8oXk6Nxxd2PG
DRlPgrrREBu+KZeclRh5bIJSr2d7upPw/v8KsnyxoyHjKtfAwbcHcp3JZiTR4iov
QcepS7NokavSEMux0DfevBAypCqTyXwb+RQ+F+AB8Bm2gcYgEu1LxshM4E1eACmp
Amnm5aIps0e4rskXFaALgbQCBEXXzKp7gfiolqfcTxddBut4vkZPa0g1bC1Cvr3S
rRKdwZGTM07aMRPX8uiwAxOcQvikcCQV+2yxoiTA0cFbdMS9mvz0dbhRxVdryUgr
Z+/uF1wcOH56HDethwSc3nfUnWAkWiscHPsg5AhSVP5Nd1EP8VCj3r8MrbJj0Ujn
ksNs1tYcTYmC1XVzAec8nGX4JAfoyMhgpoy5DVWTSXJ6MZ7qKhgUCAT3iOWhpcfZ
7Q71tHipqHicDAi516ZxozTfyu6OFnyZUcbIlUgVnuWE4TxWC2HwfOjvvPw62cmw
BcXiukcNSVKgHmwN/WQ8ReYDj27gro7ldqguX9Ru3zpkCXxh+5DoN7krFUlUsmpO
4H2flY+DyFqBfJdNMBJdZBK6xwr8q2sRkItQTT38kPU2VB6S71ZkwkEfwafJ/SFp
HhblndSoCa4/sfblZKgn/y26h7mQ/eQVhZSUEWc9/S0PXZlR5jFN0TLJHd2eFmLt
4Bj7PKmO9KowEjeLCHouyZ4JvXJi5zIK9KykZpVZZEukihf5/y9wJEP+PEjwEIKP
Ws2Dp//hANMTtGmAXsAOqidQWWnR/F/bQtZkofwx7qcyR0dyc8Ii0iXU5l2ygmbn
aQGZ1d0ckpMJFhjygBrPSvsF5E5jAgB7aEA2KQ9oH7ksbTBBy4+vxcwUbtZULj0q
ZaF5hnMECYOw/Ft8ELfoPF8bzIhsI8w23KjAvZYhAmhyW7pSVR3bGvBnMUy7BuBl
9678x/nq1KMyRV76xBCkga+YxWNSScM4T3ofDHMlpWWozBrkS5rBRO6zajIUzy/X
mfjPYiqP4DPzjek/ZcLSpPsAlLfTTGYQmzncV6/aukKOoR61hs5kh5C1oRNVnreS
YfAxJk5ZYHPWM8sU7TTI6zXPZHp8S94fdWyTNS7qKFhDGvfVQb/K0FXM8btydPvL
GC/xjAkDHqD8zaxVuNdOSPGXj1GB4gZH8/I2Z6zoKpHFKsB+Z08FfRa9fzKAvj/k
s6ZHLJ2IQgApY0e69CDTRHvXa9UMDTP4h7b5fbVyyAEqGyFnH/B69hdu1KngDgVu
uBh09GadaK0rJfsen4gb+gVTYfPDc2dxFDMGeKt82ZcV/09acBGz2E/GpR6xrmmI
+bL6T3zkT489Utw+ZjKUDJXj69rMT/TyFGSJxXRJr4IvdYaTGH/SkJ2i49Rv6Dc/
eZPTaoxepr4hLZErV+VlHLjLgRnmkFmEUqJTGkueoTobZoht+hCRtPX+GtzShul1
OgdfaHtx37Dd7EdwcCFXcVzBAIKbgeknhjH3RM9QuaQn/ILHNx0Es71LTpOdorna
LF9UvHdRSPF2Rnw2J8Ww/7GV+4U3jUVvpN2vH855mm4oBMsypTUEpfTciJ0hM/Oe
UmfU/xByK1EWllPbH2KQyKvlpTOK0lq0p7C24j667oOONJN+AuPGUzFyLnIR7XVw
8e4fHT6mwccOVtGxsLaym1XlzZ7nsGJU6DL32NL5tDXq99ouikH17QhVvwNNNOHR
g0tNjkvSWksyQra6GTC7otwqWn4wyV2hBk9XYg3HBvEzfKr2ePKOcP7uEIICrcG+
Z/5nttfkGVGtROHuP5PhoXoKB1eeNbehGnimBy8UCpA3pqfYMzPi2pLaEvpFyLaY
+IBw1GK6hWwUXB3AwOWUB31L77uVzw89aVP649IKDq/Q9sXm+R84DNW6BvZ8ovLI
myJYgGRtkjlGxkpj7YpY3b6SmtLD+XWzoUcOPSI5AN7zEar7eYeqUYWDZkX6yY/C
zQHKt4O2FUNZzyJaqlBlOvfXpj2jBYdlCSyQImUfTwKKUuFkZfTUAmppqv1uQfgu
R+dmIReVIsZ9h6SjFjwnNsogQ+18p3VOcAeGBjo6uC2Qvh7L7cqc38K63BcwR0ZD
E/at3rc21I256DZCRXVN667fcF648ftSt4ViNMET82eAb9zVoZkQspRQGOegoy2n
p5StFk+decdanjLUQqKb2npprxqEkGc8dNMzNhHl8X7S2By135idcyAp+7/rWDVI
XKqKgs/RCK2rkSwAqO5SOTV2/9zSdZdiCsQ/To3/MuGCtm1wCfYKcKqdVhp5L7oD
odHxc8cfURHGi7DkGq5CJnP9zlxgY5ES3/WUNnkzGpYM37BRI3kebZ3+J+RC4EHL
PiXZqcNkEiqVj0twqSUsgA80/rP7PFY64kdttTBznZhydtRpfbSz8TdfNops+Wjs
eWenJ4tgUJX3xv3PLdEZBbyIJCcuoroAhQrc2EGI8ToEU27D1AzyhMth9XfgUk56
nf5EjP6ZUcuFZ5Kp0GIhNcPMcXKD/ITPG4hnP+BEYK0NPh+gJqzAb5f44MS/4aL5
NxvoUyGeHSGTlJ0wK591G0dh6fU3NEslvhjB89KC2ADMmXgQgv/FuNAVp1flply0
Ds3RoMTQ3Zti8Pfm6sfcPVTesTAaTQDwtlqqEmwBtA+EN5PVnAhaS2RH09Fvp0dI
3BKWM+eJiUzpDQuegqA8USnEtv/JylQZch/dc1tBYh3ofbzUKKPfweFgT+7un8wY
4rBiTyLTsB++bYG98PsuBxIqn3zaMiBAPa6q9n3WQznv/zNTgnMEDA/mpM3BaGhQ
SJCy3E9HK926IxHk+ERcw5QjA8mIPLFqRfaV2F8GGJM8f8RziG3rhuM/E1imGteU
yQ7SoZ9HorruTe4TxDt1FG3aLu4eIwxCLHr7EXg1HUWhoQePPH1gWl1cUIjQ6xQm
plSsx6fXhIYEOShiNAMhdII/qXOfQsW9XTefVJZvcFFuvqAWrb1yGj6cp6uNLtwM
KGyhwy4fdZ6E1MwBltsgFHBqpSMdgiaRXhfOZLtQS1RxCdjdmp7k17oavKm9PCkv
/wewG++24rdy5ntlMiwT4GlCJIAXNoKCKlttEKG4ShTuDdAdWiaw6IsxLKkoIQbg
n5F0YV1XgiIiNp8s7MlQsseZUfyyUXOptWtO1EH3e+qP+qoNQLe8z1VAf3QzFgTD
XAmWvzwN0fR4qNiRxV877+rtM9l8kuTFxRprHagku43REgJypBE45fs8UWtpYBHS
sa4bTgVaqo0wc8Ajlf6HqpOprwX4QtXFAmkXOmzBI2Cn5pHhdNznCxFxTC2QxPN/
5eKICLmN4GgzKXGhMmFUPvzLsXLzMw7BcLbEjKXezO3Av8DTr/U21IXn6bLI/vzJ
06rSb0ERilOUgOJqtv5yvcOZHygH4h6uzVXZjnRsba0NTsIQiFGk5+VTa4GRHSGE
irYvlVOwGI1i0CV7j1WReyATN+ovSLzvV2sYns0oVqKeXbaZ5LSJkUEqsZdAsaVf
cLxhrVUeqC0meZOFqUE9Lf9DRBnlJw7CeCKqT/FZeS0n+o+FvffcsQffXAhXz1uT
K5Ev0+uBC0D7kXWWjlTUKN+W9NJ+/QomGuQ8gzt8Q/YjnY946TBFV6EK/I2CdQB6
B8zUYOVUcTURRm+LzU+pIYwtTkTZ6q1p29B9KcWQKGbTNgkOOenDmXpg2Oh2BPFI
GsilaXM58f2hJ/ogIBG0TX+pj3WwAfqDyRgVO1KymjDVPEftRmGRU9wnbG3+BGi/
GDlyUXUYfJnUX/D51Zmye5LfhSTp4+qr+WDy4gI0Z3+kchk7N9AA9PRCF/E3F1hI
a1Qp8B8+tR/EywFZKzyPr8dgUR2rjssnCP+S2NmzT/oM/SmxN9WY0HWeH2wBS5hX
RMTeAmYlmMtCA1R7r22i4lxzyntR/N8go5/kf3u5KtG7yT+kQnGnnVn7y+sl17HX
tuSfjy8xmWLivVEoKyUwyZAtXHp5/28iWbTYmZXALcDpmKC64FvRPV/O3EtLzi59
JqXCqNSudh/7x32OW8z2WKc4r79l/mKX0UWlRU/PAoQWHdtoHg2rtfzn7Fi1yWKb
GHCnLr0SQoxJDKfKfzEo2ocf/zrWkmp2beK82LXtN5QbohIvEUpoJ3+ZdzkoVsBG
N0Fxr8n6cBwMHVUHJsbSvnEZiUCvRtoLCEHbZs2FpWpDoDA95gWhXOGFj5JrfMUF
dEEaHxvNkje/0opHb01F8deyewBKfyQ9t0sazSTKaOT4FC3StZIokqP4cz6vo4QC
ajFuAxGTKB7VfU1Hs4kNWlzV5dcMupdndC5tNg0opXMzzZENMDsp7etVtXOgodR5
kXy11nEDlSLX9TkklJvNgduGMGNbzcyCLxAV3MEnJg6cH0OHsW9kKOngzXsB/vF7
+2wnN/8YmwpcsBckruf7QRRu8Myr6K6g9rk8zQNvQFpsWxKCWB5fZkC7IIhEfFcs
riiMdAcRGxDPoLqylbWte6NKFR1GM+Mb9jmFv/D9oZbnE1u0azm+XpiPckUsewBf
5mkLTDJcVZJVIDQ1oPDcuYgCTxPSbv5q4Uz9HML+Iz6rW1FkhCXAyfLIyEr4Q8wb
Wgp80PR1rRNbr6KhiBU42/uooV5CkvzZ1TWRIKbgTHBs2jpjWDl3bm6A6wO4XKEC
k5SHw6ZMSbLD1k1lDXL2qdorVtuht0sMLo9GcueZp2BAI53I3rfGKucBqi9ymYh7
wsJ/IJAXyU8ci9ChWVSgOAoI2EV8ePhgp3sDFNPMeXnH0prIB/1Uaov/VlPgmRpS
197ZlVCBIa9TtfvNPKrMaWZtsGr0q1HYBqgTGErfXF6y9K7xrCySEU0vLGJbw3ar
I7caNnlO1QrmZcGf5k9IAbO96ija/71Y/arjcmN4tPeegOIbSFq/tFbVBQUV+fmX
34QM+q88I/CIJdhe6JvwEeUZVzD9AbOm6Rvj9XnNJYw9Iq+SkSnmG1gIrmm5094Y
05PUgqIqYZmVtJ3z46bxbiN2Zb2RSYEttpFgTiKIEk1hldNKXYfRAV4gxzy6CN2P
nUAidX5374lguQioq63EQ64Wi0Qyr8XkuT3tXGOkwKhPTsqJ6b7vGCIDpEHUUsqo
nGOCVsT1Yv54fn2dPNdCOyuOt5u4oQaso3R8o2+vMS5IUk3I7J+sZ3RgXHjJyJ8e
PomEqpt31p6Ri0JHCUDPh7tFxBJplkMX6kZl49LMBLBnhMbgYb58FCrDJ07Pa9gO
53bGbYpESk/i9NEfn3MpyPlLQKSX21FdVFSVO2u+mers1J5NdslWAmamR/cPjkts
kuvvcg9cpBxlgd85xAPvyWGQW6vc7XYwDOj36LH7KONoGzDRTE4FweBMwt6e6QEF
wuKsYBhVLl7ohGikz/kJgAQuIqS50QqSEDeEFoA4IQdOFoiTfaMsmeVfI9tlTf3+
UrEqk/egG8T6eWoMchOy6V3DjJdnnzrczdZBMfpDpzKpVYCBqxzHlo3NELLThwcS
T2mmPF15Q2V7v2oYP6sa0QhAKWvOJWk1t6kBMyt3hIN87HR21rK3Cx+wQ1ajQUPk
oa2VsBGtJMo78srZ4oNGsjFViRAzwt7ibqhjzekrjD7KbEo9Yy3MblmewxafHm+q
YctfyjuSaiOv011nMSFGQCvMOBBUOMkT7T7lN6Pr0LhkXC3VjvwQsagiHYtbSmnd
piKcmUDv+pq3LiZgqaBj9e5ufC5GvSfCzfg0RxHqtkt5/vRZTwDLGFnbiTIj/kaR
TlkTukOmZpLxBnTNi8lJjT9Au4EHADML/g6brzK3S68p7wUAa8voCEvs4p4jB/Ze
lIDhBTdX++ws4OzK7b8k2dvi/CKxb17TY6SGJGScqeIPm0Rzcdchh++LUeFnxQxN
reYKWvY0msT7h7rKz6y1gaBewPfFyNRRsh2h1UBBt2Vg2ks0lhnh8gD8v/aHdxu4
oHo2nWSl7fap8K/P6tisti8UjMPLEIusNezn4jx52SM05E7A1UpTRJhLWeq9UdH2
PK/0zL2jSrWM1gC+NsT5ezZ6e3q43aJT4Auiiv9AmXMVA0QVdk69DfgJ/B0H+seb
fQhGTtxgo3ek+MNaRxBgaAtn0sPcZIjhWpZpSprSM4JSb/XfhAmm6wnSCNQBMd5c
ceMSRwEOXC4k7kqaCTTMpXgH7+XsWeiPigjXOk6g/EdxWBWjtfpkVYqAAXdCEuBW
OTsq7jsf2CNZVt7zsebujc3EgXuJkFhRlF0+g84EKqNdh2BDAHOI5fzY6NDS6TlH
s41e85zIdnyZuuNHXU0NudQOK+8KjeRcfmPJay+erFGODbqDwMDB32Okn2hNjCd4
sxQAbK5ry4UvBAFz1ozWezolmPuBBShKh8UU0AK7RW0bx7xVpfxXssmzrwg/g9+6
GYzIxkJdmxL8mqCxihbO9MY2oisTvwpcnk8EmAxgm1zf+RqTrJqZ9LLz39do5qyv
ixiGew+q4StUqaPp2oMZ7iztMp8idJUbEKFBr8nzHu0WpcTqxjsDzqT3STBkkBTi
LBy5LQjcWyDTnn+fgkfT/KqF8ip55IdRh2zQo9y62fo84saFa7YzqWvWKDx4whLs
ds60QyGoaenEPkN0wvyduWyLND9Ewox6tI5Oie5wo/s0xtfF/ps/7y1XUr8dVunw
ZwC7PbI40zbhO+HkXoD+xjZec99yMFnSDe66O3UTXtW6qPsxof/fumqwsurIPeMB
OlbPHKyK3UAcF4Mk+2n9ffEbVbWr5CeJev22N24WXPKEPNmBFIeMIDDavmlM0rA8
y8pE8sX2b33RID6bI+nO5r+gWkVtbZ/skH2zsIzJcZY7EeDXFIiEJeKECLVfylz8
a2QepbJiD+AY/GvPhZNiYOC2yHWMBWPWZ2tU+LTidbUZJc88vdCrNIGzKYiFXAub
n2Q4GxBP+C7rZtdEJaXQSBV1EYCF3AB6sYK1xwmTtGVUnKfY+84vGCl3h2KXzYhy
I//GnSLzEUVOFJ+E29wLPWkwzRRO0+sJQKz2xh4YBKM7lxSEfVVwLik5cYJEk4fn
87oyju/egyVAvg3p9/VpDg3O6CzZDtxfwYcTZrdXqd4opcdX0DeYsg5etg7ti56a
X49nzsobcOL0pzgzktTlzxBXrnmXTZAtrNSgEl2Puj4dzus2+6Ka6bsYdQnnnL3r
s3hJEDufJOa4+V9TQDkwRK5pGJMQGNIWALaK6HIDBBRKSnkR02yBHs/Z+jA3fmaW
9CZlQZwbGuBU4afJ7CLQ9TgIWhQ18WQNlkasv/Jh6GMx3OYTgFn/H25KHC3ye4Xj
6Kc6tRcVX1ON62CCFuQSBfkYsv168Nnhl6qyS8nrFVCspHuI5f9gktmnj5wIpwZj
4zwhWhWH0OgpiYpdRifMSN9eMo+a3tEL6RZBtZVigO9A1usE27MBMCsncIpSLgLW
M+xQLhpmUzQYuR/LCpfmEoCppARjAIOtBZyrSgt/bU/kt1xfYnI8QmDaexp8HVyi
SxTZBF2Gk+R/AkaQwbg/kQwdvGpb5oWgtD34Nf4AUFZQdCCDJHeB2AbARphzYfKg
32S0ADdD00U6RQjs59ymVcbkmDFRK7tcB80zjEfgTe0012PAlHrjqi1YvoVXww/D
uHcCr+XD7KFoQwAiYdLnjolJGaG0UD5uTQid7DienYgMU10AxVOYXoGPIlb9g3Nq
G+2oBii6P3UIivkxkec3OQyDuKN3+wG2INxnvUpTPsvZmTsa08qwJ/39nO6bjvKz
SoskLGd8hFLsekjcgrva6AzTmCjb5UMKPxPjPJ3fTm+1oVeo7htVxasPI9Vl4Vq6
9IQ8Dz6NEgIw3JCu2n5UoA70d7+l19rYJ7Mv3H8iWI9rRVSISDAY20H6fgz14MsW
w6DcvEJVA7IOQfkQ25dRR40/Dej7Csn3VswF6o9cF6iAiPP9cM8f11xM4O3iVolC
ij7of3mi1z9h8CvivWRh+RbNYxg4PiB9ER4hlnLE1zgWqpgWFVnBBEdxZS/ANbZl
bHGEPDIVO/z9o3VWJP5iwxjieAC+vYzcuGkCjxEuKdKl/jqK9tSN0Nd5vM6siQwT
u5EsZegyv3kVEMR9KpL70CP5erAY4NQ5iSBJUn4BTb1ga513XGhiz4UbHyt44ms1
P2yVEN2d1rfrCbpEJAomPWHTlRff3ydY3R9qJcxxvr8uulQfnZhnEqFsi5/9bsrH
N74T1btbBK4BV2oGFtQbV1eZSz3ZxeozfTBJITd2XjZtJzlC9EBHf6Qnib86a55D
R/fHF782TwRYZsL3KrV/FK+UMdSw34L8LDXPT6+ctq/azLPhqJjVu5imOEs5ycEl
GERc0Uc6E2tq427NptaoK7523+/M3eGzN3yF5Q2eGpNZ7nloW5kzqlVvyiEKKjmU
meIlGfh26OVCJdd7Huc6xyVUB8bpcAkpK0p9b6zvCbiVVEOuqn34OgIQhpq18S1D
jl6gLMdrB4knT8QR1SZERr5W7uw2A+ItqYHeQOqT7+RgKPaoiLsmK2/9MuuyNOpR
lh1mRu8U5OQpLVuCLDwuYZk+h6g6O627BQAnA4vYQoqmyqTR7ni2b2lIfdD6FIZq
HZ5aTumTyEChhNo6DDGujP5I955cEpzopQldGR4xbZw5NA1xLrqwezv6DW6yww1V
5KjwDvfD+OoXRTC76Fx79JSeqhvko33rCsowbhIQkP17fYRMmJsrokrBU0gHAcEv
SdICfKcyMDrtpxiQD7ZOMtlD8OLby8JQnww27KZYpGDSBsrNLur0oUq0EsoxWAvt
p64Cvw1QmDIPrawsBBC1rJAJf5A/GGZmAO4iCLSK3F7cwhoWbCGEVNGOkulvv72L
5fIzHVBkKxkLjU4hS06K6UtY2qzf0a22mGIWZ1od8g/6C1HrhZvO7sXB9w21v66+
L395M4ct26u0xwduVSwFzAnGuIVt+lxbb7eFRwqeWVroPYKHOio8m3v2EHiC1xXb
b8wNti1+TWIHDy3qBZ7wSKcLlz0+NfKx6rRdsaCynhaxUSTPbp342yBntG31WkjX
NXQxhA6y3z8OK9K7YfkQLzMWPg+M1XeWqT8wP8ub0cnD54HZvJb6/5a5dHPQUYTa
FDhREC8uLmt56YEJBbZSktUKkQfleTU1WCuCRu0ruLQiaviyQRic8IVKRg5tON1o
OdgYJJHhLmlPxEb51Dfk51cbkUgxTb0OeVQB2Uza1lGNCsrMXFoEikMR5LP2QcG2
8Sq1PbSeBGmCvli2/IAj5CNrsheuk0s+urx7Tq9C/25vkyVe2lO7tU5P/t2Rq0c7
N++3ioiDslrw2jjeGUzoLOw17xWluRhtwke5LN+ySxJ03IHX9c8ruHSQvMsZ0KKh
5/7HURGv4b30EBgll6Yrd4lBz9Gxp69ZAcoTep2pwszY8vMSVP7jSOAS5KwPH/BL
zZCtNJxBOsfNEVE0Sh2qtZDAYJTxG53crgvPB3ECwplSgdP5yBJMDrRUwiEzjY7a
XNbvVlobb2oH/lYmMX1EIWFeATvnZ6+cOeuIssQ2yu2choTs8h1K2KjkTuR4Grin
ns8HcMSfOCNqhOEET0IUx8hGOY/lYkTKI6yPmU40TJTso7reGSh612RjcbWBK7p0
0wzINl8iTp2ovwnYhy0dm+BjG3AdDGkDI5espZtwpXMs+c3N/P5cuWjDiOzbdhiM
5ZOrzDa5I/HSsNnUxsSmEIJ22WnO6u9eV2a6+YIgP69xTwdQyzf28nb//jPGRLB6
oh8xN8V8DdFa8sOnQ3TC9ihkHU2tGwIjz6eFy8APUSHXr8tSdU1XlfgxDrp/QyVS
bjVD7vzldCCFz/0LWxU1xgoswy5yam/t9FgzTOk3LIp0uw7iRlT5r76LWJ6j6ecj
ONOyOyiP4nyXy+yg7UkY9hLkzcft/yYL51SViR5Qniw7qosDsJx4uC9Vb0ooO6Lg
sYJiikEORG3W616Ji4L+E0MoVgv2dj0izKwvhwqhnjBR4f1H5QYjtbv+L3IpRDhx
l8IQJsnhRw9vYXmBxv0o6jWAjqu2n+4hLmCpwACmApDWgmNs7VH/yBx2hI6Jggt5
KOYBKwuDfO9c/gUlFtyM11LwMRfMSP1/ZmFdvqhupOik1sTYzKB+U0zZmumdB7x5
0L3equtAFTo7i5y58AskE34UAg+gSkuusHyRTDNrCqzA5qxC65KHby8FlTIrgueR
kmRQxKajGv9xprl4R+AQV6QKQvJy0neI8tqnd8ryZa8vnIPQK+vWOxrc8yH/H0Lj
jqP/VEXxrUvQRyt35ai26Luiw33uO12zAz5jUshK2Unzg9Unz4B2zCP/uebz2kGg
fv5j1xUKItVSEHXX7uIEzW8W97b6gEyzl+uqxuM9f19Qep8xFBryRhGmVNV1V5+T
XzH/Ly0A9AWYk3a/ItYHRKC5yVR1eurj6CtuiIwNBjgWe+2GyqKw74XyH8NEOkjT
Zj1AHtJwuh+/BpOue3z63jxfSD4F6TrPZn+Sf1cQNkTvTs+GBmEZpTxa+iFtbAwK
AtJ/2f8Xj5eJ66O45WW7M6/vON10sbqqXtoF1QTg1vlqB57Uge/uWPhKnj3L7ler
sl+brnNdarlEjUKC78MCX0LwonObR76ZnqVhhEJwCNPpR8wEt/auvp611bzJCXHv
oz4/n74HwjYaFr1Yrww6bi9rM2pUBRtlV3ob0+vK7+hR5EQKaEIYuNi9ISPPtj+P
O8Y3E6/Um7eG0LZ1BL6NcWu8esb9E98fEBIGXeOlRG/dyEARh2BsB2AKLCIn4EiG
LMcR1L1fYrKwliNNE3pc/c0JNSkSgq8gZNUawLjD9dkO2zZ0nuhSfKDIaMw+x8N8
NF/Pq+zE/3/PKuUrqbNrhoRz/m83pf8kEC/yreTGWX+T8jswVTc3vR4J8MJf7wVw
HO/7Z/gyqEcW+P7x0uhY3MMBqvn6/lAgpoRgprMC9HcenBGG+Lvy2g13xvVQ1SCu
DCJhqbchwPHQ0FFsGJWlUKqn60932eSZ1lIvh9PVLUr/WQ1vLb/FOpyqkHZCVolI
gh2xVdHLrciJGlA9u91eenCPuZeJ15sjUI2Y9+1geKIH3HSmJjpjT2D73wFTBqN+
LdlsHgEYkEpLDxOmVunssKO3ED1RpwyxvI6U1LbYbs1CIxXCMTtCL8QL0kHvY+e0
dJsueYGGK6ekbpDgrgedSwQFiHeAUmI+KgpkFnAYm8hdwTgrHqDfp8eRxRhLRX5X
kMhGztDHJ11UuHwNKUY4oQwPmus1mCY06mV0YX0Q6USzUsD8N1dc1omPvZbw4wwF
610O4Y3p2Ror7eGMBOJcISc4GAZW02xYujH80KqdbchqutdoHR0Had5mgSwO6kVw
nQW9HEDO5e5+O4KYygMd9KElPcG5IcXbqFeqrdj33IxFkYo+pwWS3eUYp/NQf8KV
+8lHbJFCO7wiYLAMWST1Ax+Vblvudn+FztsyQ5s/44wQfV2baMdqwCQnFNOco30C
FX5L10AMZd/Snm1LZvXWr1VFkdIStRqE+QeD1om22ZY+Ozjj9lixMj2FQsTZmR7w
ZIMHTl2Y8bTFZStl898PEsYo+q7iYe/EnuMeGOra85oRc2AY/feBdXCZpZElrg6K
OMck7IiUQQ4dAVV0VpaSu//K8NCKviY6yMV5vXIZL2j9ybDxlcrXghgxMQYyXS7k
8MzeHxrSOkWbvrAMsdeHwFAcjU6piAfeoqSC2SWy4QIgcNoasgfP45btKiv3vvni
JSgBMr9vnjj7bqviMZiSsMPSKsn/+allv74ZnbnncH967JoAoqBryZ8l08DHSuWH
bJtx9aZHfyRA2GC/kGOkRO4h4qt8bEgN/S7GeRju6/AN5US31fjWuD1krj43Dn2m
yzQQMtRhMNTDBXhV4mcBYPoVO9yPBlGZfu1BXHXDQLAd69QJYpTGYN7WBphVNy8W
ocqte+6xXuYn53/PXZoqXRu7xXLwYHyiOHk9YqenxpJUTF244wh+uLH5/hmpkDbQ
DP3Rmhk/NXtsTdySXLJchbda9VqBYdwadVd7ofRZ3FZ09i96d/PW4XpADNZJh5kj
UwAAKkrjXG6M1dObzvqGuq9h99nXB5teqHiJAQE5E08KZptWoM3QKWrpyyLxNH5w
Opi6ALlAyKeAzr1IHPjHIKVmOQd33MzrLVcy5y8/CAMnwrfWR86XuHxevkldk83a
TRsdaWkLjlNLngzJ2rKmtrnZbEIPC6RxzizxzGOMSpWLmX7prOWqRFgHPCgcq3Dp
CxmK2wRQLWfHTO5VuBSSVJWYh7AVuBLjv080efPPsVyiVB6aquOkdfmHlj6XC9QZ
USvjQc0sz6twgLF7Q+YX/lmUWnrwdoDgAnHToFPlLDvM7p6qFUTjNvqeCZRvolv2
EBQ55MZkRKw7AsAVlikK282sjaxXMph7/matmGMVOYXK/uEMQFpX+nvcOfu+sCve
AjDkhSArByXwIMbng33iSxpdiZMdsX41/nVDRsRzbpEfPG6Dya8r8fYr0Ed6yBZY
CoFc4U3d+8Z6oEHVge2/gvI04Tl6i3wGbu3ZNK+cfjUp1oyWBJRSUY0ugZNQodyI
aUMBTbwV0rR/5gcRT5j11S8BwasCBMdJ6oYZSu7tu5BNwdvSl/VOVCIeUegCHVoa
UIajnZbQJ19kdYZtSNYEdfW608n945mPqBiwsypsLAQVRRBvum3RpGfmookt8HKn
WIVu3LAQSRBwsEMtkVwUJfkXUCSbuShHCVfQilN9s92jtBNAN6Ev7h3hNxauElWG
O8Iy1OM9NrMNGYQUx/pOhQ7L55Rxun3cTZPmzqwBZkqCEhGLex5vQBNA+N2q0I/7
WupjCybSogH/Hp8SrqOdREbW7q1MJPRTS0DyXPGE2YezM49w9+Es5x4s+r+HeSxD
VCW9urkbdWdydYw3Y6uFEJMyJOza9C7bqpKDioOPugtAcELLZDq2MNeXarzMMJqB
x5EOgG8O1SpKOQc5swRm+kIjgg5ayaAN0WC5eyR7eeJXsRZgahe8Qc5flGdgAxNc
DLlLo4fP23SnRAxHy5nrt7kEWiT3kin0Ck203fGKQJ1+2FnJxGyz6+3v8Np03JeZ
NYDeytmlomDhx98q6a9L/BFDz5xpAKtwORLoZoocOkjlpQFHpjwQrtBFC2zMh7fa
aAbLnh+U712yjM72VpYbtKwMEV30WibKwVjuzUSa7oDHBXytD9XRmGEWJtvVlApA
io5Y69RsbcTboofJF0jhhauj58I6PSbZPuxl/dHgp7sou6uBGSJATLit0gG8RIQ7
J9muWvsjpGBEVTXL/sut0UZJHwWa690US5X7tt6PzUdfBoYvx5F8ul7zCO0NCKOp
H7xbrfQ/dimgiFbDL5CEpBA+0MN5A0ysxqRVCrWqWAh83cpun58npy/3DtPzSNQL
c87RgfaE9JOPY5Qs+Hx+TVbWGLoQsBbJI21gusZnnP8xJpzF7kTgXrjc9m4g1WgX
xdTpQcY5TbJ85Z70I5jdimaTnRTkgXeFj8zNwoLZ9nHLNlbTEj1vQVvTUS3l5kMF
oiGtJObV5XOiix+WtnFv1sed3pY8SefCIMVHTOAThGl1AgxTdr5OouNStVcOeetm
BDUVQfOuTjynk8biZn0q/K4k4b8uu2qbCisBielTW6ItYt+Uzy3Ciz0qHh1BcgnW
8k7Kh82rx5q7zp5ATF6cuyjjELaNXDjO767j63aAXFU1DA8h5lPChWlEZAB2TEqI
/Yd3w8nVM7lqUQwGimharCgv/mw0WpoQ/g2s3Nzcz0UizL8Hr2fDR1X3XjDZkaHp
82TLvrPdCHIyuwTE3HGhrnXyVc73pyNhXeR1vrJZw8BWURSGkY0JHkYlHUkA0Zai
ZUy6fA822g93kz7WKMJWdhDSXQSDmQdktGSz8L6Yh9QydFfElGUg1nuq6RfTU80B
Qfpzs1pMdTmhz5N6CnA/lmabE0TacCheg0ocgkzNltyZhiGVlEik62TNqDjm8eAC
z7kayXAgsqVKgUEWb8WdNQAwOX2ebeetl0tYQKF5APX2dYSqrlSJWSVYuG/zlQ/B
Ki2mMLk3lySFenNdyfED3ECza3jzLu0tE9M+YzKT3g5d5MV/7dAxC2fuGGih1fLV
aXCmG4EbIna7d+y8ra4Hy9XRBHfA+grTHoEyaShDp/SrGR31uaBAVQpyQkc2WEYI
zIAQXS3YSoeynolKYKHyCNoFNhB5KGREOgg7G1ly2kML591rGBC181UyzN7LQO65
u5ekC2dK+Kek4doApbRFvqVzzQngkC0WKKLMu8iLbAinka/Di84Hi7iC0/YymsVf
Nv9XbnqSRENkq6fyyrMFy0UtAze/EMR28hDkODwH8FKdoGr0uyBnKscgHm45V1Q3
en8evxlgMjk1HcDdjRe97NQQg3F5gn2dUvoi6Vkm0CFjTdsyDVlkVkn8CINZxL+7
CxvfzgLItwzJ/lAjjWVGDegnVcZDhW2ul0kRmJPDZ2s8HMzri/Dmhj2vJ1qj3fpF
w7AKc34fRhRwMDfGAvYiOEAITPAEk+nnCknnWtn4wcsMR3D1PKGILuCTJQpN0GZb
X2z5Ro6gdwupOnrcK8oGmPxGsgCfHvPf2BzrdMWkXvNZEBfXrcs72BO+JeXGIT3c
Dpxxse7hSajsNQ66yUOMA7KfT+69t/EjzipXklHJY2jetw+RKLjQ+l7jIm5FQi1H
C3BbZ5nOwpnKdfHJ8abYfOfW8CBAjrGdjCb5uprSOv4C+HxhGXQOCeK7d2J3ZiSc
ZY6qsk3nEwDomNki5jJzKwxub7M9DH95KdqakXRqIHXVXFPKP0bG9C6bMJ/1PGR2
PrRsOr6RMQzWnEJIMGt99W0V1gpglkg40av7OyvfJEFMrtDwWvXwqvPFehOnI1L+
7C6tHZoo6M1OoxKwkoSs5tUmXzJlfyWQ34PxXNo9uuDbCjBaeL0FrTqJCt4T85DR
/gg+ug1y34LP3NKX6FBC9kZGnMJ1dHd7zrwUlKdT6D4fh76M04Zzrr3km+DQMCUT
ibX08pKShFw2754VMzfkPRyI6bm2kvvz2OojilRddT9JOvxRt8etFcimmIxc1mlp
BnKNVLzOfzU5HELELAW8pzaygCl/NNSomzR7VPfxrywPCgMQ5jWjV2tlGhpu0Q0l
waemrDr4bDkYYxY55YfTM/uH+ROLnMbgKDmvXlZ2GMlV6PtSC5YY0K+TvgTAS6ri
ZtXENzLILibDb33QM9JCegIjmzU+jj127t+SOUpZFCudv3HbzYj2tERBqQVBZTn5
HpAQ40MZ+/NIEACKV7J98mju89rG3gCnfQJN1hOrS0tkA7bNL4NrmrM2EMRubf7+
sxLZnp57iwwJ3BaC/XreRFGnuHCOJCFgvmsw0zqPF2QYyHBqKdSCd99mzp2sQ1sE
MYMDIAXFU//u9oU6tsKS5jw7vqj8WLI0c/hxafwNIKwaMzrQd56Uig9J3GeAJ1e3
goKu0fc1UC3rL+o84UiHcy5sOiUtJpC/NzKcFWg6LtLpnAHYSBfxdjNlvSW5l0Fp
+HHsu6W6SowP2ztD7y6a8Qsd7956gBWAtC88xf4jrT5FR6BZdrre2PgshOnz2f5U
yA+BM0bqMq1ZNi37k+V/T+Yvmj92IskZV8Zj9uk12cwy/om5mRerWtAWwocAuGb7
zF//BPYZhdv779TBGNenty0+TlLp5pdLnuEgfYdrtERofg+z5iVlZ0UhxQ66vmQD
/MqDVxIrQStM0ciB4tDRQANcJGhE6328Ru0Raw2wwtrbMOl2/ewTKEVF10ehAEJJ
IDKtY6pG2rDTMAG+TKWoQKx9mYSgUR047ab1J+XhO5IEtUJhOQ6oajR479NKj2An
w/9B2IanFLAYLAOT4Ko6RVqB63n6jwYcJWaZXie3GELzSHFF0tGniEi9O4tB3nRw
I8obG13HgZbZ8RhYiYNo3daR69Lcr9sQ3Kud2VieSZWc2rioj1iWe79HoMkA6y9/
k3oLAei7LzLTE505hmdr9NaObuRWYl2BCP4/sQI5wll2ZkDO5s2ZoOxA98Kbz0In
NMUd3b3sQDC+r+IpQ5/u+MqABggeMzmIZWLL/eaPEw+/hzsv8yrA4XlMmAOOHusX
XA/NyP4mvLeddIstO+XgrRqoLuWcXUO30kIV/GT58Mh0LLrgShq+MLHhhh/hCtDW
tJCLr1i+JbZeNH3KsadnNv1qeRjkJS50J22yFY55KC0eyPIXHgKVGQKYe9QtMl2Q
Mhqytjo0ToWRyNeoyhBPlIdkVpzK60ZYzNo/YGveMIQ+KA1HzD+oJGpQo5gUTZYf
H/1Gt3Fv5xqE6gVpxrt9T9AOldCGIN9Rt0croEAo5p9RNPf8C10ZNKVKe7OzyKYA
9VlFjVfaprwMaw4muEAq2jrOyiwQUH0toiB/TL+E2F7DgMY8MKZUcJLDRoCFIAKY
TDwVlWukwcHqS9oOge1LK2vCBtgkm2jkdu7N4IIzlyY9C8T+baS0cHsVAdMb4D+6
ImWagXYYpMXN0qofxXePrw9iHqXRnY7JnEtlfyNpwcRdyASkRo390GU8M12ErESx
iSCfVzQIykEPt8ByUYGWNppBML2T2i3+n9F588lAwGRwV0B3HdllGeGucXYW1p3g
8zF8PWNhbBesqBX8BChfpbuPxhk7+ElzzmgU1JtvFNM4IAzJU96kX3ljHlewgYxv
DssV/GGew9psCT22c3r9t3fjQWSq6CNHxotJIW3Ae4sH4B6YaReI4x0612RxkupD
BoKIQ1tsM8eXZhgGhOG+Pxb54fji7saUrcHulZL9ikAdIkrKmwoBOfZpbki3J7qN
ihqcKlWapwegLthNwXTNf7b4m3Vzp02rPXQr74/I3Ehz2LEIacWEFmlTmRRoojEE
rzgyYSGhtEJ7X+WNVxw1XtRi8VqWnRrXu1SctqlNPer5XEYbWYql8g7tmQQVzAcw
bK3va9S3QH7QwHGw8HKrGYjGBDjIw0HuBaORUKtQAcW/pQ0yq7x0wpNKEdJKUDPY
rCBBC0g5vIylc3ccnJBUA8ZbPatm3a/ISPS+o0ZuABEX7V7OwXt8eRlZ/9cJFpXh
pCUb53eJ5t+KGrPePOoSVa+BIhMeT7zkW5uLT6UxB1d12dOeOAB+z4b8oGd8s9xX
GFpKO4/NSunyzqSlFXKlxXkYs4gQuUkBHyNWiYllOsRinWgrpuGCI6Sk7EplKp8s
lmu2hx2I73eQ2xT5czClQZ3rzqFcNC9xqWUof9eMUZ/ghslTJ+s1X10lPMWZ+sO3
ZpwGqRRSaCopnZuRmZhVwKbK3zoRa3PhevBMk7cqC9S6dMsKE7fsq9I65rJ9bcfb
VPsy+Qf3bWydMD7S1QL5p+yRmUs/8/Tw2yZrNWZiO2Pp3UeRDMBzqK51699u5ae0
Mp1RtNstmFf6aUwYAkQyHMVNY/8Cbi2KWdzmaK8I6OvL4c8vssPhn9cyycnJ7Tg7
qfbMhfobsy+++Y3EaZbK5kdqxAof2M1KySsEkQmMyqBaG6HuaxyV5p6dQDwIy8px
bhCQQSDIYwgIc0EkAyp/VbgEvM1HDBr0BLY0TA/xevpiOyCSFvePS7GaED4LX+/1
IDhYhlr+CdzvLWzLrv2EMDcs1INF9HuPojU0M7GvJj+jz4SKGdbjIwWHEgfHvOdC
bMrDrzCCeJms364dwlaLP/Is/o7GilVEsnsQQ8USPHvOJFGGxaEVYTtTNeS8uDCM
B/QoGZohfqe0eHg/H5eG+jssFyT8aT9mLsJ9d0I+8i4RKUnz//u47LXWoJVAZd5w
yoI8af/hy8As40WrZrKcuty5E512IPYtRM4EztgLojYr2EtNlQn6TGrcZneZBNYH
7LFWH3uBRiBch3CZlB3G/lY9xuLF513fAjad0gy37hjf19tST7yMFhki4V0EqOHk
0rw7XSwJjCvRBptZiogiIZ6oewa5ylxBWde2cJRTm3rE9aaKNpXr0IhlInVEVPBi
Nme4rkU5Q6uEEiQTeaV4zoGFlYU7vnjgVW3QwwCcPKZ6ce5AhmXX0vc7WFaLQiKT
cNVNyu16Y5Vqs3KShURbaWXwqpLMTcU1w2y9n+Ygdjs3f93AjkiaKRv8GXmfL6Dm
D5jiY7Rkt77INHELFT8GdBDhqywugOWyPP3/ix3tI1geRLyz5v42vSu7y9wj9hZU
G2FZKMue7xWSwA2210eQWqZXUtr4XUfUw+WsX1z3WuR9GAH+oT5725NNMBzjrokJ
+ET5wlBZuXYWkAwAAS/QHR+N60ze98di6Asqz/5HH8XeS0wsBY5zoRtrnVw7GTA9
wLDAeiszrVU8E1AjImSX4cijgf5Fj8WNlr1c+UMun6WIi97UxMO9/zjyP36SdZ7Y
0GY4/YDTUWap4Vaq9d4LwEokbMPQJB6fQ2WQu8THYXKi0Q7Wqw1jT3xGn1pdIf4F
4mfDIyuYD/D6Y5QJc2UFAnKBzi7NQPTK1+PYiAt04Ppy77kzpnyq5zJfcRUsOhVi
bf1ZYRJlxJvoYk8ehEc00qUqV/m6QPw2qNThSxSnTCBJhKEJsBNiMypxZ7361uYv
xGmSlsjm5s00nZ1w0uqlrp0PQrp7kWbgHn7sCNb9WcsP90IKAte7ZGV9Ux7ZxTqy
pu6CkcxlB+azkuknhKLaLv0btMwJEQR5QUkvtuva+RgdvaooA5mnuY032Mkq2011
zCUFeF1v8U+8ozV7Qb+SZvYbphLPlcy2fBK7Zi20AYuBNeFvyW0kqDmFGmKtrRuK
4Bp/7jaSQCNbHVKPeAZuxkyQ0ow+Dgi4xbeU/90SLdWiZhLyFZJj8QSX4/n/V0UV
/xkKDQyeYxjVZHFDhn7fG4kO7r3QH2ezpX7o4kILvfFcmk5jWFe5KFUxgtWTDs1D
r1pLcm8iwkFbkelzZVpfFsZJVKw96j/o0rNS1slP/7dsWp1fmymoZbfS93QcBPqc
PlQYnUNpHC0Hz+mIRzA4t/0Z2h0fU2bFIpK65qbgMeebJGG89dnAIzSYsuwlKakq
ZGxokB8fAls4/HVGNhnN8WiPUYleYZ8QjnaT+uSFeRJfEdcbKJclXVi60z7z8PKm
qQCdf9q+gcnws+a1tRVMo34CYHDkNy5lGNthY4cMGcVpkoiXq7wHjtL/pKvhYKxy
EzHfaeT6DcwwcbRQHYG9prxXT4fPzni3AdR1H45RURfECTWbUQLjHr9GYJD1P4QN
nnesu0rIJk5/mwDfRQSkPIv8T8N6AjQM1MfjmBzroL3DuoYmREW3U956yTza3/Xf
ncnZIrYQEbRBWyw5UPkp8EZzOU8Pke0+WTO9U/awifhcCg9ahh8C8WFd5yPHLjQX
ZbiHiYtVrnJo8U3Kl+cfYJzE6c98cAWMAg0iK3H+LAGzqk7z74reMILpMcQ+Dydk
2oc0yAL7VMtB9QVdHMw2iIEBnO0PjEeNAA1sOuwN2Y0k6QmWpYCxViXoZMcff0UT
hJMHZmb7cCnWv4R7IvOCEjKEzv5Nwv1fu7mc1s/1pHPooELsaKQqwtlCumeN0KD7
AfyLhaJSASyKLEdRzUDYGgp8Y5JUhCBwGJv75szWtzWhpg5lCFBUDiWbtWwf+ZL8
h6DWopJ1ZPXpi5FGRO4MgDE8C92nQPbPpDncDgkzewRhVbkYv+EWYntm1TFrCrAu
8t+HcGrC2x4ixwr6NFlJji0MBya0zhcHWjDzrhIrgPngdc1Hkkph4y2KRKzNMDgv
YDc/yjhqF7wEzFUBjMGmsvpxB8ICPyu5SE7TthAvV7vNfk6XZPHKV1XsLK5GbMKw
aEx3L3Cb3tJka62AgkhlvumJBAnoMMdXms0BoFlQjbNuLfIwFs5ivNAxS2vSGxvw
b6phf/d9cZ+CmlDmUgNNt+MQfZoXNHVVHkM0wYVs6l0EXhejAr4i4XT9ZsMWbk5Q
rJxjF4QNcwZfYhowphnUKxiaU7iGEsP3CWi03q/iUkFRAE1RnIKH01vTkNzYpg/A
FPqrYsdEJ/F/LBGCzMNhTmFxsHJ3Z1Gdx+Bp2d6l2ziVo53obZMGaBFzK33yJ1Pb
maOu5ERL859uwe29LKAlik0LPd+kBR8kIme7B+x5f6deHnWRC0nXrzYZPnUdZ/Wh
uHLPLKdQHRUGK3+iwfFugwRCcC26QrHz2wYwmxuFKUZtWlWH2p6pLIZa9fM4+S+S
mYKb9aXVKmDJYtop3T1BBs31dmKq5OYsbswqJyxRCrL8WT/Gjrj6PVfHnjyiO4VU
jF9k8WEsgp3I2Ms777VPasKSu8YnNyzIVnvxxPhgESv7wS/nlN3z6zSuPXq397Ka
r0wPvM/lPm99dne2TNLWBEmxyaFFoohbRGp6XN6lcG40hOkS7zIIt/G83CWo4lrW
HbZ6wvmvau89OB8cvQAJSSoHbCbLU1FEVo0FY5jFLxOlRryrA7qsxmEaMGtWS3oP
cMDzZUyUzyaPBEKmRSjJrlFnaHmffmGmG/ZrDrEfcoAMjANu33mElSHGm7yLm0w4
mVYZ8Ebstz8Mi4WTzU5GKjEBDfTRqb12OwOrpsmYWasZyzopUrDf+6HVcpQyVKYd
7/3Qks1B7yguoiHOn/YFKHbToJRebQ1FydQirlPmugla/v1+3ujfAmonQA0K3Do3
XSUU2bq2pIOqSg0Lg/pVxvQcNH9U3XPmF6faMJIIyTo6UUgdo4cFrSjU77S7Ja22
remkrgqeiOa+YwTr9rpOwfswKHpnNzUoFvpCKUAYOBG5cwE4zlWjsmTP99EFtrPS
KFtc8BkQZ27zQ89N+xMVgXJgldkMApHX4JGJwhIVknq4NIUssN07tfrfEQBrzTiD
o2pnYXT1SQj+HFdlm6T/H6EUkLaOxkmOe2z37ynAHHYGmNnRgqM9Ic4KWhskbXpa
08NbKdCLUVupNrZwVWY3lMEZWzMJ09TMLgG9r7U8XLhEMpTyY25HS+777xBKgqBO
gMQZ9ie4e66H5f+G/Y8z19wjaH0FwdENPDL8+uMgU5JtWex0p4pQfx/RJvR5887e
5L/y4PCV/mg720UgoBe2729/JpDPHAmTULRZA3PUWjhBv+V34+93RH1fVCVR36aC
Gj6quBNi25ifPrl/WNxx2uLS0fMijfAMVH8sJ1eogu0qblVlsUW5v4ldODw4AYDv
CfHQdQZG3tcqqenrHErlAPK52GAll1Tlp/b+lAKk3xwFzzvIBsamOJs9+ArHRdtR
Ub/5dA9++IoZ+Wzz/w5uLIECAS3G+bQemxsQaO5PCBamZW/AqSTTHM2AwbjhD/Yn
CsDCprP6e1G6YS9QhLiIICig7UZZ9nGBBXLBrQSgJqrob1mmIFKR16vux5utvYhX
k8C7YD5s1/6u0tkbrEpsUjASpzgSDqc7UxehRDLbFFFdO0ADoqAC5bmlOSOl4MMn
Lchng6rIucNPHbZuVMXdm0F15vxdGpfg4hiNphtjRv0CUqP30HimUq+cBmSYt7iT
KT9atcLECti/qlWOftusGp0yuZgO2127s9CNo5yMxRGFP9Jge1Ec8d897A3b+mD5
Dh062YBb09tmzqrZ41VWqqdkTSxlPYT4QBVwfAt3xA+z2xHGFc2GUjQos9oKYFo6
AY+I4vcSvbbYxax46i27BZlF5Z6w8dWTDl4LqSDiRY6JPEXyYRuh9bK1diYoS2Xd
+bxJhbq3a+wCdF3rHPC/gwBXlxjzPKtoTWe2ZDyoBjV70aE0kv3OGQA2EAtXcYix
qvc1yXKVG6685UfiMjqGnGmLrqspmJ9CjmNOroRUMX0IoDCg/6a7lmVJyUuJxJRF
XLCtPsAGa2QaEv2RdsUwjwl0M96ncyJ0hdWHkgl/oNo5/Q7IXKTK2gWTOfxUmPCI
Jq2MbZaPPh+FrBG1Hn596AHDZfHd7xb+wPA8/HtiZTcB2azQUy2pAOlCOvQEuJTi
gymdl0YI8IzOcxXeqgK2jE1rvZzoq2dWORYR63vvxf31K7mxxuZJ8XsoBDFMvH7n
KjkrUlzPc6h/83hF9L7Y7OGZSUwbQvHhVYlx6A8zELwJRhqsBN4rPP/al0uYSCtC
WrXs8dWPZxLsSmgyh5/sL7RDaucRtPDxafvrvT7aqQ2oYmSSHTbpcTg/kWB2dBwa
aijrY0J/wvLU8TNE8CrwRIrTpx+HjNt7sA+0pxuxni1En8S8V3fWLnAKEyWiRBS2
cUfm+doKXHypqCjfLhN2zO5uFNJkGjwGvGBgEPuOxTWPkjfClVHe803zyLr1ZrrJ
lKVddlBopIlZjMC2OWt5nOgNXy+oIpg1ivKPNB4w28NAIc7b0bbYc3d7vovs9IgF
9V2qe351dO1kC9nO6Wr6NezB9+zjNhrRYS4/QVlNPvAU9njN7XgN2CsXHQWWjaea
LBRoybt9lNBO052pVCX0xh25Uzn2ttIxvdsyPGs0gEXCAUrrU2IUHQ2fu6ZiID9X
ib3YfUE4IzqzYMXPtgQ/VuusmLLXHawQpdiN8Yw6PVBtBG9XE+mgbFu9D0dGHEyg
ZrdgnKmZeJXOhBJFf/s8QoXv61TNI7gOdc0Ih5LS9cx3ZyQSaYCVt9Yj5WPqZUz0
r+KVj+tnZmoDp9uwdJaH7yRdM7lqKI9nrYmrlFKN03L7ssKgo9CutHWqSLb+xR59
jxN27QBkARVdEPIW3f+vqpYwmpSrFK1RdMw1tmwhlkQHjUIMhEQaw00IHIHVyAFX
3ZOD1jht/RZXBV4/qyzJVAEB20vNT7kJKGuLA/irP2PaBomKQ4K62Y9JuZJgUeFu
qjLLUeJzpGihMDKk7xXF5YZyoBDsESYxxCAmnYUC+zk7anUTw+NWcLVE/6P1+EFF
r1Ree+8xfWmzkikE3KhTO9u/2HnSZYeTizUIvISSiomxWk9S+8JXmunG6//Lxhep
0bphOXtoETFJG4MnhkqVHDkmgnadrClX+bum6mC1pEOG/fBJrPp9AuSy+Jt9y/xT
ND3ROuEGpn6FME1nRYpWtBpW6g3qusb9cKi4xsLyUB9SQwgt684aIvgZ0AUD32Wn
0agiDAvjJFrbJgXpAMCHFtQkpIvjG7a9cmYVaFobczFdRPu7vj/QE0VYfr8nidow
izh/NsZNM+WAkZmEuwBu1hYjeHmmEmHCRIx1JayZS7triZB/hdOQlJ2dLjs/i5M8
PARb5HrvM19AoQHCDhXzbfAQkVQIiif0e/mYS2r6dHBeYqsjPdhT2BTleZUSiFNd
SmNMAOEoLMSqHIakO3eQ3UrkmKpSkrz82ZC6vJaf1vnGnubnEDBBMLPgosoo2xoP
kn8x91+RUmrgFnNwOWZNgBgfrxT8qbQLm8htrNkyXVKOqvwhFvp5L5sos/gWQuY+
5d16J/uwfPLcx953ayjRuNZJf7OiFhz2c0FfjTHXs0d26uSAO2FvtiLdXHUQPOdI
HHKLPquZTAFKwopelorgGWZi/Eaakni9DHL9rbFYKqmJjiAv/sws0Ag6jEqfTGQm
r3tcA2X5rINTkEHJ29SA14Yj+8dwsB4Y3D3tZvzGwbFKJx8MxNsK8h6YcIz2+RKc
5Euia2N6I4emklxD+F0WdEmJvBOHPrtXxpDlLW/TXUYjmsI7JhERWjQe2tn+0TYX
fvpBaracdPYIiSrCil6JzdQXGF5+Ft2qrD84HrXuf0tTlVyGDUJBBUD6y7Yw++UR
asr3lh4InYkvJMN6PlTldpuUn4kUXOZkWhkvtQ+HBxAuqsAZCP36KvUwVclyLbjP
/6P+FgTluzj9IBKqxlSNLWlHtzUMsGHV5B4ctWbn0O0QvKFHnTCB5M5nzGW3MvC3
p24frtu+srpBTHf1XcNc48hIWJRm24daPxB/cnM72GCvaufpYrzInFQ5QFunKMCy
2tLP2BdadBJ9yHf4ueTXhHExMVEmQf07wCwp1Ji24MtGyoMCDs3RCpk/uKKFsXnJ
Hr7cBk/giRq8n+factUcx14k1XOIwZD18HLjF1gY5Hs09nmOrttArzYTQ7w0JLYC
xX+FTl6gHyOpq2UUIJNqPN7faolLPtADuvnxtu+IvdoEi39Zt8A3145+YYJ8lkG6
vD0Vx75m3qc20INpXWWGD76K2UlCv5jdHkdwjrxtFAwxauBmThhU00UnIcKn5yPU
zgn07COylasgRnt9D2X1jmvUL3TSxfpbU3Kx4Barc34xBvw+wOnkfMrKR00L2ziQ
D2aXICYT5zEvIVdZc4l84XoK5eb0B2LS48BDPpEdN8CTVxXPoxu4ul8oaQs3D8CD
Slh6oA7h5bHlYOE49blbDoDSHwFpmomV02EEoTv4bk/ZPzMEEDIzpMGgQhCNdZXd
K9iBq+G/DRkavN1f0PCh/uD1RZjs4FhSmvDPCbgiSsDu7sXCe8toCM/DXPiCtR+f
Hh8mktfJWXhgCcg1olrgHJREZ4NmQJcGi10um1WXXoifgOXEG8wADCMvP/g/lQRh
PRB2lb+LZ6Zm4FPKTZbhuBKbIMlww5u5twzDbZ3nKwqo2YndNG7dKHDfZBURqdwn
HiykvGMcZpvCISq2WSbu/1f/ioaVweQgcZxJ61RCe2Seqi6302TGngs6niERe8y6
L8SM7//E0VoFAV6VSNMhDZSzAqCG5lHpPIZGQZ/9bbdmDh3u8k7PFsS1f7pkJA12
P8aq0SCR3xOBKGxwSUpFSQX82u3Ert248AZDZGHp4jgXODwlbYV12bcEA2CHb7cD
8dijCOTFFEmJA4wfttGfiPQ49rr1XAL0MpDd7gQrT0L4BvqmD1P0g0xXeHKKTC/v
H4Rd6yW2ZrpCzuWYLQoAUGYD2ueQFhqoQzFQTDrU3kookozWmQba3tHOX7lny57w
zVn94rmlMMYbBV0DnQBoYSMh7n96gi64QsVkcpdnZQYN396N6SEvDI4YH1O4sQ7a
/keLs2fL/Qsz2GaXZgQYtVfkNTe7ZF/CWUwOAVWXNOg9hKiyaM1xGip98SH/lR2l
1pkv2d0jFbHj2b21aR2N22NWu5nigPJxkuQnym6W3qONvnF4EPrP8rLuMCIHNzZk
ywxHiGOtn8LtIpdQpQLXatLDegFDFwNXiUqGm+3tXzq3iqWbPncCNnZ6ganTYKH9
awz9eg8Wck9JH5gdjAWcjkPcdGo4JtOv4EJImX81TID92azETLBHBlpAUjxn5ncN
NeDiM7YaLYziXjPhDLlal7OyVd5EYfSsuBRJJEvl2/IPfCw3XYSetwj2MUVJqGPt
A/VYO1uw0GA3fSArfhslfkq5Er+b665P+PhVUZcvr8bs0GpX6Od62WMXAyTP3Q8b
IOF+ho7odfirxxXPFRnt5iGyWu2NzMk1UTzAr6bV2i9kCZglf1o5DTH4WMEk+WdN
3nwdWjDsqGA+K3+aUCGTocLaH6RuJ4Su12p2YDhRmie/GekTqn30MHpu2ca1VWui
7nFgGejIVgSgeYVMjXLadFP7YhcnB6JJbhXtefdWVKbrbrDXcIU2RhQMf3okI41c
G3bwo4NYPzvlkPgdM9PCj0AnFVkTyndhcI/Jwoiqk7ExwnwBux2wCK+4PO+ipvl2
qaNmliJsQ7SdfBy8elAFlxnIJLfm+qz6mQkYq0gbhXctpHH/tqddjzINa6aZK0y/
pwQT550GrMylASMl+8jA/4I3c34v78XYaTEFR4rnhdn3y4RgrXF81YJeqgLVj0bH
d2frtL3jAnU4Xcfmh9G0kRqkTwHC/ggKgT7Znf7MzAYekelGg1BpN6VrUtRpl2Yv
pQvinScFRHXeORMtlWD6wiRNAJwq6jjNwyYE4kOMKdUVXDsl+nfwH2mwo1fguNXb
xBxhT40wGMGtmd9tEKSTLrMlAJQVOI1tR/AVmg3IdWA99Kzadcf9rXeemKsgT1QH
iyWGwVfyUpaq15zXUb1c264STtgnlebxBSBZMrxRUXCUeW5KNNOnEATiIW6RV75g
GQ9vN2JuNJu77zT89A1+AzQMYo6BJjrADH0hk7vUowylO1i3lQ2dwGiphYGD2wtV
TA+Ylj8AoHiyPVZEVxemWWFAXyOnvZxk/VZ5FVz9gyFvbiHCRbr8IsgZp2CT3foy
cv4Xq0fZoe4V2/jJpoIO1KXHJ5qhAih1Hr4qW7sN/mPv0Gi1Ge67589YJb+AgG6U
hbuKS0YOrpQU7AeIxLKeZ6EnzCMdCycnhHzI9eMZ5Kkh0O02EHwPgSjz7cEUnnL/
sMH4GnajrRKN+RtTE+N2V0yEEfNEDvUat8dtoZCU/ZCpEftLIxZyDmC8MkCOyjnW
N9EQ7tWfzBAt5FKl5iFmYvnXFsT0HP+2qu87E7gIDEOW4mwftcMrvLGZ94UA/+49
I9Qm/hSwv9qVjmMP3nI7V8GCL/qJ7BiDazk7QqoGQE7l9TzKiKSUbAG20jTnUoNQ
Grzsdh+7B/ux7hb8PQbZHULwF4iv3IPd65nbWeW2Gld6dVOaiaYioBBplfiHMxUx
+K/op/uoNdi9Rd0zRnFc/VNd2aH0QeuRpeEs6T/oAfOd1O9Ywm+eznY149rNSzIY
8zGBsFmyoyvZ74qNPedAKmnbV9bIQOQUskuDchcQOvY22X4CZioGSvAQSe2UC2Lu
bvs8O7x1sEhM5FxlunD19whr2gIBiMbiaG5/xVOqWzC4wQHK+M8LWG6PoKIMJgyp
vHbQi91AUJrIiaNxFojI1JWE+fbtj4Ngj1g7Wbv/Ac6r1yjBrJM9JPuEQX5dOAaG
tgE0jYrssT+5n/fBWMepsrUEmE9ebd8FPFtpnicG+zKyHzQU6grdx0+S7U+OlEAA
qbbOwYc55c7GObcwoRNADO/Gzi8J5wfzei/kyTsjHgvqAoYUEgBe4MdcdKi2YM66
Ae97XMV1jiXTztxJcWkyHJBI1p0GKoBaqWfA71OEIJi1jOnptu5PzNPWCmsbq9Os
en7tbM+jpdO+1p66vBeqcwn/MJpwqefPZySgyJyFBWpFVXJUGZneyQMCBzetJfV1
ejjM3X+doL+v3yYtg6IWMSa12+Q/F/K47rJekk8YTWn79GmIeIh7uhRWSqYqe5Y+
9Oz9M2/XagQFHN/jeLV+zYqE9pXtavaotK2GoLRYbg1TbyN4bpOJHM6L8ydHj7mK
VdrMB5asK2snsgObTfY2FTK1rwRcRx48xlWa0kUehf0oIfVlOkEN2U0AauhV7+AE
mFWY7On5JDiMiHoKLOEfnZzWNuNShwMlOIimk2owjljVO9nCqAzVwdMs8obPO1PB
bR9qXCw3n1v3chD0xcxnaG49NXk7HdGB/W+CGLpOopeGFzQHZwvVcRzL2di8uohF
ONi2OeoQJHSe5YiFXnwgL7kc9wWxXJs5gCzhJcvD70xLHc93qOWzLXhv/w9Qxpz3
ie66hLyiq6rIDpfm0M3Z2ZsIapFF1vH7vr8mrRsDIAeNYILZAKLBsdZbOmpHFYIJ
mKgUVr87NqjyrCsBL8tYUSrHsrFNF+BwCWBBcGpo3L8pyXyLippWrEVeVloKdyJo
5AO8K377/srm+YGVnOz+DiHI+tn0LzXi8t79g6D5YpK2pss5VpdtwC0pTNlJcsxK
Sf1t09pJb2V8KD7jhAW1Tkbsiv+34PwfWnQiULHzfcSsfP3RKMeMmREyuhj3bwES
aN+BeIrAOadc+vKLOrk9SVQn03Vs005oTLvNHuqG8rktIV5mR+ohRuAqsxuRq8JS
bE65O679Nui7IDNITJaqBtQk6eiFTRHDMHcFrxp/fuBRVg2BqNdxP4d2VcUe+10G
eUQ8AuPTsbIIpsPEoiWypssIxuu1+CJcDxpV6RpOJGj/AB+Fm54tihE1AaWAYMfl
jLJEKcQ3nx3uMhAVzLUWrb6NqD+dxMYbPkS+3bVPa+C4vB6hy+f75AbTeUHBuRTm
H7egJO+p6yJWYuJgGo2m/jDI2WeH3O9PnWynbXYQtLVqpqYFbqePTO3W1OwSWtwh
VOVxvpioWmaLD+wOWTGOg+KkeSMZnr8eayEZeTZr5FrVfr2tBlYJUArTfovxIfmd
6BV8o3Ct5CKauBv69U1iDrT/YvpGeJGUPCqKg4oKzLgaPnstJ0H2rhEh9rgDaa8P
nZvR91v48YhfpWFPf5TAFeQDb7MtSwIHEHNQLGZom5D1eG0LQ6bctYGBsXBhMehS
SG5KaeOaN7UYvyHiuxvR+XNWNDBC4FqgJlXd5XuScnmKufge10dyXivUwOTccQrw
H4Fq46ecJiv1K02ONMYm5vfK0XjgMhxYHoux0LisnDNn8GwHR4/cf2m1lZSv4qiY
EyP/XfvF2WvfRA0d8F1efA47JM4jIUy7vLP5ITQ+8HUxcaJJhkWhHEnkIYCgVV7V
vGhI9nP4X89aAWVK4KWALjMNq0TACssszATFG2D9N4hf3M6pYUTYmaMBpPDMeYRF
o+9/xFT68Zqz8ez3t7+2oyj326B2bwo/TzxB44lS7WKJUVgsXX8PKxxB2aMbhrp5
e1cAluK3KOujoqWk3LYHgDkRbRNuTH5gdpTNjMrxZDwlwFluB56yrsvJ0pnWkb4a
INt8AjRKjDGQ9O4qXHbG0Y8jV4gX4u4do8vUQMT/ydnMFk3e7ezk51WAgT/YdHXW
iEN811K51+hAp2CChm9G7cFDlaNlNzfxSqNUYfjno0tWYPgEn0smIJ6nvbII1jyo
6qMv/eg8++SVmJxTuc4HwzjpidNVCKpQC2gBrxF8jhxT3Khsmv81Cuni68QnnAH6
guHBxGmKaZ3CSTxhSvS8oC/NngAaWbnGkMWhGcOwooYxziXJfpT7PWan7Fum6D6W
zK2V4dUNJ5abw92+wbsPv6dq/yEY68HFUMFktIeLju6+EA2WM4KZFc2LIwy+ecKF
7atzYYoiN7miZ00wJQx5Iknxz2G/3dAHU3e81E7LxzZPKP9nP4YqnE3J8akxoPiL
wWPYWixUewLIb9GtJijjjGF9f3GKShsxXXcZuDSfNqVJAmtHxffRGG0y1lWyTHdz
7HlBeo1w19lTqQw5owTO/Eu2socR+yL+1mXdsiH9CqduihpVIeFEIXjF+aT18/fo
gx434TWnPrKJ/F7EjRWSqtYAuACkRZr1VIqEigo72IOSw3bwtbs7bZqBDsaXzHy7
pyEAp1+f2nVPkzE/S6wcorDm5tiWxVj4GIPsbcc6DvLUMTAnFqYPV5mqvoSTAtfy
U2yZM572sluOEdEhym2jRPgXDEFx4Ql/f9X+DQJmulotA8dS7/f9mt1H91p0psfb
RZ164AfMReiYGfbajJBTUWWZQbQ6wB2XIK4BETaYrwridVnDzu/7RQ4BWNpe6MbQ
s/uyZWX4jUETjxlqp7Wc5k36kNcmeHhocgEz29YoDEALGlurwCAGuvTMpM77ouZT
e6L228LDJZqiPbAdKooaGpHHMQMWd5nT3wYEpLuZSZjenxiJ1uJh4fTtV2ZcdBYP
wg9hUaqlXgAIz9cglZ4vr3uVIoNq0GSZdBRveTZU4Vir0Ne2hg+g5nX3VSNgcOTs
jiedp7RIZVZBLrClFwlo8RxqTmFQJuinCgvQlMcWWgXEdhZH2Xqyy5/6uvPF7/xs
F3XhKK4d/2J1rJAk2WkWLppsdZcdaGU90aEyh6m35pGY/2xuVD5IAv5JzgCWT0vT
J0Hxge9EymxgqsbH96R7px5XdU/YjhsVv6rONU7cXj0b1Fc24tDSKQxeTrE/A/9s
kALHUUy1fFZ2c1RopL7JLMBoAjVIcxOKpk50yB4O42cTQrX/qs3N0e8H5jB9DXsk
GA4XYlW5DXGHRxP3tpVvmiaUu/l1wggpX+E+NgnHsk9eT5wbR8OMhutTk8J33kzC
KwgZr6N5naOJQAacsHValFE24hP8vqE5ddxw+/xXIrHSYEaCiquL6PTQ63mHUTwR
FDTuXeFXch0oSyxyNNC8MW+4jF//O5+vsy1zBI3rjTq0JLy5aNu2eKlHNlT99pnc
NQSmRIIBMWe2dtJBT8FWfYhe3Q2hlCTCh0oSGeQV0dI/AX8bBudDdb0i+KQt71j/
XmM9sDfHsn8ZiJQYev8nJehK7OeeMeegt12yDlaUdfQzuBQP+RE91tkEFbcNLEgD
q0pg47FCyEvYdnSO8cxH/46dH3AT4PyuuM6zD0ed42OpD0TBhxtmm8RRZRkIoYtC
DM4B4k5Ah/rY9D+k5IrdtWpwXllMwVOZFUFwZjDvzY79g845pk/MjOr0+PRhlsde
JEaTHfDSQOdEXixY8qR0+uWqyFcWLjSs4m/m43KcjRyc8GEFBMmPzaOGngUOTtvG
bTif5vLzVHa2EaQPfJ6ReTonxL1hJHd7CjumerNbsdPSw972qkAD/0UFSDuRP/VW
z39zF8QIaS0TDms8r6XqZPnkDJeuwhpPJGje7ynJnTK8GFa60r87+lYAKln05SVv
DSezC1Asz4+Bewy+nAM1Ic6Hdb/bIm3UjCCIX/ODTYz6TehlehDRB8yHJITA+6hA
dd25juYlAKxn/tZBOpPwdqkP76qxFoGXW155XhHw+EJATvujaG2lZ1LdBxQ818dw
7AdzexKct5DVz97s20bPUXAyyIZ9YwacYRkEvp2/wUGlvA/kXMAf09ioyog+KIcB
iaBZRYwWeZMeOZ6+6dKiH6eSi3Z7O85zcNcnBcWBLkwVctgX30rH9haKA7i6ev1w
chPcs5SZemfQnb3BWTkC2OOzGfkkcu3a9SNm4piF35KaMqW2VMWi4kjKD+JzS/BK
PQbB4z5zKDx0PuS3jm1Q3XYmIw3XXkRQhsCnxTMRY9zS4/KE+jDcsg5y4lH8iOZg
UDdzKCkzaHQYAE3MCgGnC+6ngn7HjJ1ewT57J9Pxh+oM/NfnO6OVqTwogj2NV8gx
qXCFGUHJGNeYzrdOh9ZguC0VomkZJ9Bkak43MQDbtMCJqLtSJkdjfQvyEaRT115I
fZAPTpyPDls4cI3ZNN/LA0ZOSr9vArd2OzbE8Y+xF1YSGFNVJPPaSBwfRlLalvMZ
5fGff5xhDH8mav9RI6/E0cS37Mjgp9ExHH1z0HSl7RYYnviWuOLyPoqxppP65yfa
tzTZzPyTOEYlprEBSVSaJu5egb3UCnB5FeJRvVKdi2u4OeV1rmyCISiCAxgDqf2G
Idi6TgMfLHlEeJjf3C+dBIl8ce8DZ0sgvTdIsfSuLf6ssEthSjInktfidJh/AeW6
Q2kAsr6yHBx+NkVOUizW+KtmQkPzV7S9Gw0+51Qk1ivZPdePvjGqBg9exRv9QIxD
+2nH2eX8bTP0mFDo0NEoTGqnY48Hxq1j0HKSwmERle72YdBP60rKzyV8i7S61+8d
aPEVP1R6zTdVOWoYkAGGrFIssSSv+i349arFm+Lpg6b/wrQb7erk90u/PsMr1FXL
FXHOuS7fvEPgqdplsvXdDi9lovz8auRO08RMdK8Eoa8bS7Uz+YXp4w/ySMKo7mYC
Y4UZQ5cSM8EK1/Nl7pOcnEF3Y2K70wrxUm9fE4d9y+QkwVr4t72/QRvbw/poTNIK
oPTpjbcha5SNZIliFIvDGaA9Vlza62CU4P6db8NzoRuGXhoP59TdeXbCEoXx4hoK
W4Fa6RzF30GXON2XWRbJIt5VMeoCSgW8MTQrpgOvQThuI5XQ/c2tnhwHSNSu//x1
mlMqgs+BzZB7DRNwGWFW4GK6THHJ4n6ju6nhAX6o6xd02nVuM793VaAd+gSyJ0qU
lKxrwdb0QS8GcYlHR6WzygBBuvZKPUE6/Kd2c23OroqmVQHkIBUoUPIgD5w+nVC/
Yoc/6IMIDCc4YJ3lo8qALF0/C4V99w9BGNYr77w2clvYA+jSxrVRg6jiOh3MlYtc
e7296TQYi3wwpU1njwzY6dkiv8m3YpagPAHDG650Iuyuvx8Ws/K/3q0JPI/zD8Bf
rSN7R8FPDLsbKq1EqhQFov09Mdf0d7LyyI2qTkrQZssW/JuQystiD+1p8rS68GNl
mdUy7djTD1zUchpitiyWK2QGDVBXgFK4p9OegnXJ7uflab3LFIcgChdxwzPYI/Oo
KQ8vp9XkRRCbhI64XUJNAvN/QStUtwg0YggEGExgx5PiZv2y0Dk0eaj/2uZ4kQnK
yDodNqnvJDaG2yELa/WnlPytbAlcv+IkCF79h83v9Imi/jUujZyfDwNzxQIKc092
wd37ApXM1EYlYqBcrWl45COq+j0a32gOleFKDBvD6jck4BSJzcq/Vv06hOvC7CSc
MXN+C7wNepnxju2womtXfKXgPFXv4aSdxwvNwnxW3KhQM52UXE7T5BI4UPcnThvm
p1XjGChW9ruJ1T1/3N/o2AFys3g8OqlvtJDRGquL5zh+To13oyuGlM8xGxAe6sz8
/7VqvGhOihm7M2qHM41jlQmD/9tB+iB/t9OmmUn6Abr4ekRUbVYPHYYMBX5ZQFVq
MvZkko7lDYLGCuYaczyQDaDgOd0tpQa2Y9zhFhxot8eMYa9aBnVsvm7+VNJoczsR
PqJ5AsKWsP8upmDFDFV76Z6WRbRUJ2OFCFCw18MCrV/AMzFnrNMnj1j7vI0v5YJT
6Yd/ukXPDwn/EO/pS0gFsNe+7tKrzIGKqwbu+57aZjhyIpx378p/mr/hocCB6sdn
6NbZ/TtIRfkmBSHYntIwfodB2xST95uEq+VijOLC99pAtVkX+2IV/w4nF+3CzYCu
UHtR9Ebo28clKwtxaAl4hdLIyPi5La9gcA6GfzVCQevLwrVMzK0+dGTgGNGos61f
OK+KazbXM8YK/DnPFTLPZSHUNMSqDwmCvMrB9auijaA8g3F2VWB3ekLatSQQcCzm
xXnq5VCfItvo8w7uBGj5BNTbNVb60eHFCaVnspq0LggJ94L67glp5buVUPXU+9Vc
m6FkuVzPno4tQcpMiLKiTTjyA234MPB6n2tQNB+Gjgfb2UfsNHROHhC3tGrJ6ysw
RCHBbfTSBpOvBVZjRiq7BIfs/M7p+RPMaHWkUXtkZapae8w9lU7Rfukp7sBkfegl
FOZ4pncvMEpSQLAiYBgAV7OIxB4JFLzcFKm3laUOaQhVi6LoiBjGIFp2vKJAWCM7
k5w2pZI24dwrrZCSF8qMhCVcURFmiUfkgHFUHsPc5re9vAdj5oaXOmX+2/pR+ONv
rnGGjXIA2dLjUmxe6ZRI+GTY0r4LTqFh6p/TR5mX/Zw7HNnsTRcaRkou0Vjr5ftT
gWlvND29EpCv2sV/oZ1rTx3OUyfHlabu3MoP9sZ2AXZbSpzUViEBsPG8z5T/5GoW
bOoXqCnM7H5HBPlPPxm1njZFEW7Rm7zj3p53h0dRQeH7KN1Ij7Qosm3kRAKJCTeF
0GBCFlWu4aarfstSA+mZZKVxopNQhO+u2gh026RAELLwaXqf3qlpj9XaSqyqpyDO
5Ju6dcYlmF/rl3+DqRFDh64XpkUVRwnKp1Fykaji82DdlsaBOgvuS9cgkgazVvhI
Rb/VmnRMofEer3UXwJmdE3T2rd5BVdG2zs9FMjqyFCldtU0gueeBmlA+McC8rSDx
Rf2F47++LrQJsT1PdXFCIs5zxj8XyI5s1crziIklHkw38CWtS3MwDM7MccZPyQxm
NcLUdIoZ6r416lXb0AAuM3FqdBu4mznywoGgwODt30puytOIb7XfxmDKEZSg0zO5
Li6q5Fq69yBueKpZTqLF4LzOGZ3xVgctfd71ovmWS5w6NcImNfya10DS4TwxaQcP
3KSBkzr0vvYO/4ZZqKGtxKyj2Djf6R6IHwHDiK9ZUls1b622ImH6HM4Yy8AEgZNB
V0LEp7AkV1xDdEu1kJDGiO8BgJdeIbl5Mv1OxKJICUUWyZTYFOg4KGNJAnFEd120
Pc7SioAh5H8U29NOyXGE3dxScYZ6wjjowhdjNfjobfQafxB9LIsJyBdJiCJdm8XM
lwddtgBQmnUFfODbyxEHGAeMqF0bBZfMapdA5/J2R1FY3n3stij+i01JmsVw0TXb
lV85+0bMWeq+u5qpW474g9aRYS4yioWoLe7RjPKEKcWeRlvlswlhKGL6D9LXVgS+
RT6JwpjdSs69pVNCIs9+nGxhM3vajyNaA3fUXePcTUeQwuKKBnuJ4wXUA7MNJNEq
NA+V2C/ReqVT8aIcQYfewm5CPOePzzc1hZlw9XylMediOviMUzrtpGR58bt+Xlc/
YVu973zGu174WIVMe82+nJpiGH+RKylE+V+QAgMwTBAhiW0CaPdIO89kKaj4p+7/
o0h2KgeCxjASGfDHPy0ztlKsdHSJzvBsSucLssAQ4N6uySF++O3r9+EwzS/tMYya
0eE/FhswXmzNEaoI7CBt1+eJ8VaeZZoL4ylF7NPGOcrAu4+1VDIuucwAtRxl4K0z
isQR0j8pGv5ZlXcMUoaLKAoOEfhGYUqM7KJNXDIfCfC8Ql42H0c5RywTbsWFnxiW
1ztPX0299n5McxdAYPlmbi/opdrw5Eq+PfCQRZRP3GhmT7xL8mx4g9LexCeUbwQU
YxiTWOmmRYofNAe5BUsxPKq6qh3dgkmtNtpzJU/+GYSZSHeGAC2/8nADDffRZkor
q16ycvssIwh6vmw1SjKWsEF0K1p0vo2f7cx6bFOHF/yn/l51jrO+gC5/fjtz1JH4
f9imC8jWdQW/hnOes+NJk1hEDR2eh5aY/oYuJ1bh0TKOcCFSGb5em+ZGqCi4sqD/
YEAsP3YvGlkz124PYssYRGP+rGJ7Une/dADMjJ8Z2mM0b4bmJAIRJDXYbsVjCTUa
LvE1S9+90dh4DycQZO6YjGj6Mo43Dmq7+Ph23yw2oV6gHj/4BCtofPomwCJFZFTd
ijqRimXninCSsm8amz9PJH0puXKnGdilfeviLH4XdwmanMZ9vjbBsB/SmxcrHzBN
P5xh2erfrehH7pZzWjpTARh8KMskN3RJ9/C/JAtXz+WpBeCmY29yAcso9GzKJibe
TW3xDX36o+/zy8aWKd9jROriKUzjycQLLPO+v5A8AaXrw3xfbwaci5/ChfokO3c/
bbjXjF+mQW44aHBPkFMeU0b+MBwpbxyaQzzLRVuqY3YrCkcLg3hck4z7kdWPshEi
v+DP1CrpSv0yTqdb3N/QY6HYqx41zgxZCh/aL6KgbrQkMT5QfyfvKPU/ktmJnqeS
XsPZ53D5O7G5JRGCKYV1uXtxkDuIKeYMbMJhQUGUl24GnQqbEarfJSvezuaMJP4L
TGIv0vYFApJ8tawcmOYb+glZWL7uRqPza8PyVrJGaicQ1nphkjDbYDokhLvJBJxP
Z1mCucTwqLtUy59mU78WZmz40XV01CycP9jJkXrehFhiURPNEQkn9b2CHSai5s5w
arZM3fmsWUjgMTSG4cdxlvy6gECbeLyNvAv3D8eLQy3wy62ohN0Sd2bTm3HiHSR6
wVyExdLH89serRtWsUhms6j3oeYijLDInR422YN5wD+tJEAII9jMpijZfXnfAo78
hHv0XsyBj+F7BJnPIGvI2NHnZMuWiKhChA8TGvSarGCKoZjAopgdOZNyCqZ6Co/r
OfZ5gkVUy8n4etsOYzs86aGQ0GEtDXCYqIU5Pew9O0tsF7kD5gzpfU1MKsz54f4i
YiK47YN27ezoRCA/vrZoe37yx3RCnDyyxsdVTzNlqQn40u21xBWat4ZODvOjmohk
KNPINNWlYWk9jyZV/Pi8YVifOfE9ieEKMOPb6xQWbIxdEoOX1bFRI3wx78o6Ghep
nmIIcvg+U00QNxpWONNlhgE+QLJL0U9VZqHwWwxPKtjWJmFBQaoxH96K7eZx+8I+
OciOkmfK0nxnV6BNxGhxmrv2PYym2MkAHLLLnTRVkCldcNR1C6g8KRbpoIFDo0XP
12paRpYKmGjxicg3qKHJ8sD5aXd5KpLxleGh3PUjgLY/hxeJgMqG0npI9El8/B2d
hLZNQ67Vo+V7d4obzgiGmlyXGZ8rjaKWxSfb2JJXQEb75e3p5kvUZlysbdAjKoQX
/0j7OBfd1wcBYWrxekcOxYzZyEZBg+UPf/2osq4AC4aSKah/7/vL/dsg91PSFLuk
4SqWQHc8BZdK1D8e+RN6EliwxAONjYw22gdkmWG4eGf9mvyVxgjU8ia81t1304Py
ROYYxXmCZ7FjXbQsLXR0XTbmaWhRKpKbyVq+4mL0mwrTlGyRb9uPFAqOIvMQbv08
LBg8n5M7772Z195Yx2eDR5+IbU8jkNUSfdDyPCkbvmcUrmMyjEPqkiLQoi6qx+Be
DKmgmTi24zxTNzf+2WL9wY4wC38BZb9Jki74OfEMuT7WVmIs7+IcqjanqSqOf3fW
mNkFIeWMv8XXQSrxCJ9Xn+YQnHJ4SH9tMp2+mrmXhFf7vJLzvMupaCmGQ/rSb9S1
VuzU+0UnnF1YLbOYiSe/B0mwBsIEBw5M6zKICS7/isI5gZrBdIwttUNuddCBBoKA
8/1U05Qgz7yIAVCf9mUUxv3/mbJcoE99pbCN4pkAmwZ0uXOwCVkGFOKJT2LmPbYa
73QitNbZCD4YFxsEt+1qbA2L/bx2dYsu2vDkXcZymh8816D7PdEd6ESdwkjrRcDr
O9OkGZAXGULDvdfLxLH1eJ7t8jDV1f9yd97ciEyQdrOWaXxB61N/aOZSSyLSuUrA
svUq8OO5noGkyKI8XrG/ody5PNaA4UOkTMm8UCiHUMXytC89r4JQiGsaMI2XW/by
86gTzhoL5hkaTfYOMvg35a2K5ZWAKQfslg8u7uCzO4jIkJIg/ZZCs307mGfjTdOE
k5fa0DwzuNB9PoQa/LMhzl4VAfCS7ZvjnrZ4pK8sg6CvOemTh+F650Z9Ma+WZfLL
OwGK77Q8PhjbCXwBBshvJWACX7Z+bni1wr3waB+LhmqAVSK2aFatowrVB639gwHD
/x7j65PPdJrqR5+gJmlPnm/mrAFX85ViC5RfU504r/ioufShfyZfm4cDqzYzwAxx
AGKEO9EPVxBJNMPu2sDNln6b8Nz9cV1zoxdC4G0Q/DmP/qTgAryTqVCVCoatCHyK
pI8wmsoo+YRKGaE3KlO+IErvkugy5AXHVMN6gQoikqFVzOjNG/jTc66JLlUpIUFN
NaWNH8g+czD7Gx661BISfz9bnh7vsv6Z1wFFoO0ggvMNMiIBMS1vRLDWVQFMBi7U
AaI6qw27BtmBaE+RKmrYd831VcYiQ+X82H8FkARK8vhHEkF1V7/WJXloHEkiIN/4
7jOsoazIMlT8j+8gYgU3swz7VrMxVUNRNI+uiujHfp/TSTmyDlX7ZoAXBP09UKuu
KYS2j/DKWV9uOoQbq2Uco4vD6glQdb+tAHGuxgvu1sDR+7dJ67kHXvhbxQo8CB9T
PITyaPJwRBVgqR0ZFw2jf9fvpZTBC8CziPOb6vf+P9XQTOD/U5oAgOTPP1AYM5AG
Ctjcv2vn4rlZbG8rYH52Ss5j502BrXuURCtT1PP/oBguc1L+jS3XmBatF1NCGGIi
TLA2XFMqkuRd0BM0tF4LkxNOj5WWod1LOJf0RypZxdHtD2mv3WD9PQJUYJxnTuir
gzdUxbcn/5VQ4pmYwyXnpGs6eWoztiq/PxtyU4fv5HddPB/nBbgE2WkNbzaYr1hH
7XhJl0KINm+/131JyZJYvmC5s+Uv9YAH6iSFaVwQ7mmLMw9Rx/L/PD5r1rpJEKXG
ifRKLrwqu7688QQONavKCatxY1LFjL9t/mibbHOVxzuIivhZYKYy0rGxffoM8nKl
LplPwNl4GebL2ocH68xlSObMzAvWpjDfb198pw6a7Xaex17+mMP6tO3VDzBUZRlY
ZxrGWxobLE7Pdt8LZwlS1klM9N+ofxhINr+DgDOSH/ZSgGGjkziAvkRBvGKiaHoe
uUT2JPsTe3P9JSAzqMkdIdJHnXHTP29FXRr2bCN1C+96sK14y1pcWO2/95b5z3JP
bCjDv9jvba2VgynLBpEGkBPI2R4H53FmvVgJRKSvPOXdvAK8itHNQb76R27YQUiY
aaUwgq2M5FLneOEVyTUsJWHgv9qSpDwBTd9mPYXc+P3E0hpn7MAz5TzYrWyGluLQ
sUlS6YBDzortsfi4X9B2O4KvO2Oizd+RiANsXWWJ5unRwVF6DdAdvUqODlGTf5Md
nZ7XYGaNec13DgIXyt1GOM486Z+85Tw6QIp5v/1Xlr4O2zVdNLJQf7ITpImmSr78
E1eWAkghmPplV8YaI61IanNoSv/CYya+CHdTX57fEgyxEpfIhwHRgUHuzVHrXnrX
myk5HfW4zFHm0Xbf4HjjYwfgX3PIo+GNg7kQdbVXmaWRGkknP1uxT6GQBMvtumB2
FvRQ+f5PzDOxtJrTaLNDmKKtZC7J3wTwxENA42a5Ha5TH6/KYnuZnT9Q+pbwSwPU
qEBxABS0u61U0EIr6Mc9kesYApbpJs9Ni/a8mGC3/me5Po0bCPkqu8BdIBV+ajcQ
oexEJelX7QBje0JIInyQZwxnewyH9CNCHVf+TCexOb6rTflBfiVPeWUrS+H2I2vN
Q36QSyChTakVvAbowfSYazwtqIUzmLw/L+cx5KSyAkL0IOBuorNHZx3ogpL5nhp6
2UKnl+xglgB+qpyzGS7Zm3RsaGPvPJFjhUg2TdsocVpyXcfUH0xxd80POf2+Q+Sc
YPk6vVgMAyE6cuewERu/ZZGG/zULT1Yv6k/xBCAIRmR6H3/0ry1IlhykioGQ3Y6x
gchhfqMiKW2KafkHqo5g9C48LlafXOzRGapweXli4pomAwuPo9EZZcJkqFsM9Vz8
A6m1GGIEWMrv3LST694CMhe80nP88ccj+VZNoQp1xLu62pPGYSfk6xuhdiX/KYwx
UUkGbhKgAHb8VNr78jmE8GTdbwsZFLn3RPfwIaB8Rg3mz3XGX8NpjI+5MgGMHuRc
nIwpW9o3Qih2s54BKWHrr+CLBAYD67hhnWnB7WHsmchnHnHQ8gh2hCA4ZR0V8r8A
+Ly45NYpk/mOp6FvYQm+2HLvVdw34+QLL/E9ap8L78oPmYRfgWiHfadF2xhuqJrI
e04KcBREjy7np6EMYxVjdhbIrrgk1bi9W74ZSCbr/mCKRnzjSGqcfq9dGhblncdD
ite5nqgO3Ghg+H+6Iq5PRImtLguMNhTl/hBgEWGKOjASyrym0LJJRwlQO1iMXYDz
A+ee9T9SAANq5dKT88pjlylINKC1hkkCfcTv95ceHe42Jz/N2vxN+Hzxo7azangG
e9tMQt6pea14/Ht2J08C9ScSLmW1Uaic4dmDKW5Nh0TqUELIDavrCfHkVbJm5Z/d
N2Me3JVRE9dA0tp0ugnna1suqLGhi0EfD+g0k08o//EkJ/aNIqRSmWRYby3acyIE
KVxDVcl4bztxa7QZ5aCwKH+UrfHGqjXjRecWEqG07d7jiuC1HmMmAETy/NDhIBHF
CXljC0MGbvuDzgS4orSuxmZPOgknD2QTxCSaVLk1U+ZhA1VM/yWmMY6C8r+8AnfA
hoLDGTDbuF6ITlCW9VcaG3+8vyd9Xr5Eo6COOhJ0YEublH9fR8Lav24O8Pfgp8Qn
CWrGRz1PyWE/l47ZbzjIMQbmIxY/ruzJjDpI3zy2eQgQVyUrcsY17026gwUe5eUi
l8wz8TS0uwju977CkBpIl4oy1yfu55Z2jTfBx3+y+zo5XRQEOZ9R849xr0MowOLh
inyj2FQ8t2BLkdKUqW4i6vpcTWZpqkon45mWf7fByKJYkpM+wAaNLPkIdIF6qqRR
Ew4pDJIEZOHpBOdycrawv18eZmqDCDRPKjq17sOaMDcZ9JHRhTXYmUsQ9U1HQ+R2
y/m5sPiziPoUXpgH2WG43DSbZaNRK7qgmxtIGD8FbPGhuHb1Wx9g3lkhQFQWNAwy
NPwBHTsXCr9T8fPbVu/dvY2OVLi/OFx+09OtfWTiKy/7pL4aom3CzfT4drxbf5hr
FhjSp3Bg6WOxVQGSwMRNEzN7k7bFHGj9CNLy9nzShx+fy5MIM/CBAxF/OE+QIRJY
SJzPImmS4R7O1LfuF+PmmVtDBAVxT1ZNgE7/upPDRRCPczEG9i676s2q0IugeY5h
TCPsilI32yeiZkQgMBeHpiNp5MZkek+25ElbwqjDXWe4DPVcFFioPTqgrjIelE79
1/4Mgn3eCJ7yAuJsCyzPYV8Ow1Pch+Veo/1oZjYwxloOKPWLD01SAmD8UWyan7PR
r3hPHdFswRJpBjrYpvBucX5mNxqZ/zAmhesKT11kVuITTILO0U4Xh8YzpYEg/Lru
c6HpJqMUITyXpalcvmODQMcSI0kBL+lyO2BwUSU8ODH79rTRALDuhEGG15vj7aSV
C08AqTh5fVTO1sub+DUtAOAG+kd28FI8LFbx8KoACXq+HJd9yCskIKupGcOkvwsq
2sLcvnIJ4HhIrSwZkusZxjtm2SaVCj5rehOjGlRERizyc7FZSy8DsCCBnoctW0i/
d7B9gzh88CpRVpMLxmH0nXBgMM0lJcZLEN0JlNK6zDXJot0WjQXvJnet2ZRkMfuh
arxrtPVoiGrfw/cZgP0HB6mDDiov7aUb6/Pwo1tRkua4u0BEOOcDzdUoncguPbvV
TGApgCNn887sDTPC67/GrqGFee1DpoakMz/klO0yEx4QONobz4Hb0PU6QhFuRqVw
T7FqmQDFS07mM63SnoHhuILFUzcYL1Io7nS1pzJQDrUUqpFYgftxvA5ixEI932lR
jFRwJ+XFibccbwr07tJ8zpstil7AVJJlmnF978Q2RISa26SMIsNIFnfhJ0LB/csh
LpnZ/JZykiAP+kOr/X3N8lqRgrbEqEcMqiLw9jk2hpFVRYIGOyXWgLiw369Npjcv
O0e+zTHRRlbSinCX20k7njBfZ9W3OuWuHpaRSp/SpXxVhUwiddhU3CxUq32sXejk
CJB/DtVOp/qfwnK3qiWk7zzUexqajcw1daKPSDgyJ47tbm/ORK4W1pO2tK0BfLIc
kMxc3iwb6PRFWM16qh3qI/9JzR3OcyhYrM6JwQ/QfVoGaxGx/uz/A7cO0oe9B6Vf
g3jhop8iipRPQjvLUGkQNZFUfBl2LK7W+HYg71Gsnb6z2RCpQ6D/Q5IPOYzw77OO
ivwA4WEe2oM0y2pZcFGq4dGPFC//VIucwKXe3sFjsBONLGkp5MlZaKKscBXIuD/Y
pDdjazwZcKTNWHW1gw+KJiaQsLBsje3c+JL+DSfHOGEQ+QR7HHMbUkMZJZx3G6XP
J0HUJTV/sHusMJsPDAhjBl4Y9Z3pcZ9+Rv5tK3DCyws9C6AhWM/dfCieyqjLK9h8
N1FbI77xxrqsPOd1jahv6SUwvf1YWCLos3teELXEzx1BNOkUcgqgEIBvbu59DDXY
bxZGPh0j/io0S4Wrpq/w5BOrbbumGOz0sNu5+S4V6shykeOXSVh/e9n+IuQ6C7eO
CLZKjacAvpvSNsKCE7ONddiaca/ywvR4kpfm/Ygq6WHnjJfKYWsz2WTbBWZCn8Qz
hPZSoKZxRh15zaMMVG82BOkX+pCCBwIHHrKyo5KKUBplqj54HbZW9692ucLqRxdi
khcOMMIkWqH1feLNzN+38kysHwJYPcpowoep76h6qAPcjN2+0PqCmTssto1+H0dx
rS2Rjgnu2t1V0IBgqjrQ0xmglJnqV2hCJuiExw/CsrbOUwf5YsZNy+GZYg32k16d
Dq+4rYMV7BEwPHrH5F5ccjrnuQ9I+C5kivKIazKdElGiJbvUWPQoZRg0qTnKuW5r
nIQn/EM8Im4hM3Daauc946TK1AUYLPGdnoYoN3hgeJhBCrMjPLUQWSexKq4K7WyN
6RhkNRQhKxLG70QOe+GYIu7uvkirWiuFP/q6E/9o14SxEAm0UiO0/R0A6eTePHkP
kIoIwHTX9wExieKvIGZnSvNBnnMogwOh1HdRw+Z1ZCnd3mEgJV+X0BXrJPaHj6w4
+LjwTlsdh3E7FfXTY5sWCfRt3T7+NaDgaZtFPVYK2QLZphaOsUHmdt1R5qFouwMc
lXioBgez/QzcqL0LWO7GyzuweV0A12aH8/mfLH+95Mn3Bk7YohhPAG/gtieNn6IQ
vdIjR+jfVcHJXb+uAkcCd8ul6TbxONGuqUVDE4g2D8fbrTnc6P52Qm3qjy2JQV0t
7eWvd8IOR9cbUnKhTVOgu30K+2hc9U7l7HBQG6PAdOYFyeS4qwm2hxEgzNzs1b4Y
3xKyL4mB78p7iGbHv1dDdM+McQrw6mWOO24L52yPzX11dDCXX3oxq9CKf5LY28nw
efzq8l5AWS/BoXnfnFOtu1PoU2cYN2KgBTCOJPjExRX2az1FKzy4WucQSoxqi5Sh
YoJCQrH0fhpYy/uMzpbtGT7SvBJZX/KOVo2gYDqMwFzDXT64q0auXYpOIIGPObK4
m1vGCC9JE0QhMZDpXi87RRpp0UQmVEmkit/1o3qjyjimHNjfww29P13+htcxtcfn
2DdXW3nTbIlWF6nL2qIb7cYYQARfocyVpmz5F4OsvVqsXW5qLz6aJKzJ8l6/3lds
rQkwSSjjEoZhrPPVeq1c2mQzqlum+zpp9n+2jdOIUtcMxZEYo/fFsQlEUASqGHF7
hz7BKkaLjm1d2VyjK20gfCqoMqMMn62Sws8I8WivGWo1KNTh9a88Wgodp++jAxXu
tZ/ZPb1lstEOxblVf4y6qw5FDcDqdCNalCh8XeXQH+vVWanpkGICoct4yoD30OSB
mYM75JiA7J4y4ls4D6cDO4ya2BS+03rDQim+J+QiCONU95zbsNnhdtM46+XHoDTC
EpHAPPJ0CPkTHGf+nDDcWjt4Tf1s72NVE4Z9NkSmbCKbCT0zzegCec81lyE6nBqB
iYg6j4EJ5zA7yWAed+afMCsvDy7UMTxfgXeX1xbaWAv8o0mECajaG19BEupl7cfH
hj9VUSehNNhlwiJ6SZY3qdSAHD4PV94Lov16R9QVmoqOKvFbnkh1SBblzeNjoyfd
EWlFMtmP4eHZs1o4bd2YKEvUZp2dOWGJtotPrl0X7Q40P7QUopOPIO+sF6O4THJd
hgH3GrQxCra+j3JNk5GTX8gPmLRFrjobLiRov5ZGMyZNIp4w/Vh2YvF+NwTWtwAP
bQHPJwWp5dqIy+vdLFgmZ8+hlda5yIspyo30OqY+i4if+gHF+HovpJ0IYs8D9ElY
KnYtpI7RU2WaQkcXRQbcecjXIqGp+57nOnpLv5WK/l3hliZAsWQw8pPHP/xiadj1
a1oabReXe5fLSqPeb7gmWuHrnDERbupodvrEsunlnXNbfIxIXSY5rW0/q7EMcD8j
p0TeqiH66UnT5h9iO0rVgH+jKR30+91f5UlRT655O1L+63Cr8OZhoJlJIHnThVtY
IlDLLzes5DeRgCCGvOtgZWHshYOWF/Z+g8XNgidRMUua71/3U41OfmbOL1LTRfmq
cbIXJ97FxEGQh3HCJpIBMEIDN+VnNl/fTf6FnVh13yFX2RWN0FZoFOzRcqoZHYHS
M8C7ZjSVPqdedoSYGWcHEg==
`pragma protect end_protected
