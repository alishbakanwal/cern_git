// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:02:16 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Z2lCHhQt7Th5wxYrWUUjvDQz2lRD9W7D40WGPnywC02xhdwW3Q2rPClNSpkvFJoi
s//gYdtpF8gTe4P65DF4etTDqhk/hNoQFNF+rq4gcfWSfSljad3G6991mBiLfwE8
aZqDgb2HL8Tc9qXOOc408Wm4v7EYaZ6V5TzNHOwPUAU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 46672)
QrMq/ogjqWPUe67A1zGcAgeUU+SUsV5m4sDIjLdRSc3dyPmjvxCdiXgSdKRi5MOo
Cw+YZcrGM70LLEFh5abiWmhoCRwKSMFROo3ju5om+esEJKd74qQzGdhxivW96rnN
ALmzKDgfe0FCmWo94k5k+4E08rGEIjmZvbe4JB70kn8XkF3uxBB+ERLe3+UTPRrS
h36bx+n3ANsL7v4Har94bpYlaEZnfTLRp1pEGtCdeZTAvegqn17hiGKMutEIYhZS
NAEONjC/UvajeXyanQqonCjMy2Jhh59PjTOnEHdZ5R95J36FLzgDftlQYlYG26zM
+1vhNpq0cdDaZuU6ov/SPh0c+BsxmwemeCKymy2d6fEd12u7Ee7kk6reqfGLBF+G
c9YOPHAuqa+QsR6WInMQPacPiGuRrzu3HCrAYbnsFgkCTYmh6g486/rqx01n0iyZ
Y3Q3+PMuCRmiGkiZaAYo4gUpoE9yVCNAQSM9/F3Q0TzeI4LiZ8I+B9E4p9DWCQ7a
+h1T4fY5TBBj4jNRORbBafkwRDH5HCz2g7YHgyzJRB6dKoG/3iPbfLAwsCvj/L21
arwYJBmcMaSQHPt/y2hYKH60BBj8nVDpRrhRKRwfECGTZsGB7UF5pa5ap/yg4/DG
arxhPOjJFeGjawbb23tLxDgWcLh+PnBUK25Rut4lCPhGOEUL/5P86nalPWiaH2kg
Z9C6u7Wgf8MfvREaxA7Xe6AkK6vOwxLi4YEhpriBhnt3Kt8IL5dQw81sy2k2plwJ
ZV4Aa2Ec1k02tJyBIjzvvR+4X8WRQm/Qu7d9xm/frd4/SgVn77zrl767b3MimYH4
+7+WttJGKl3200AoGF8kYlCNyy02eATXni2L/TFNf7yqVnBwHUJrg2plwN5X68Yf
pufbKreDivFEH1fV4bKdZGc0eXjc6J2Pbc7dZoiGaH3jU9ffLtLM9CK/N1myJQ9f
LNHAEN7SdY2VYBAqqFRTbgvCnVCOgfdpXj8FJfRw8T+1MszbwXlmoU77+i5Mc+FS
ClAo5cLHwK+XQKcLpirxYbiZBof7lvQi6/19QW2VUKBrQAvAENE/w/3CNfDkqX2X
tcufxXmczqB0oahJY8xLuJr8gNp28jioRn8+4q/d9N5c45SZvf8IXtn6ZrI/2S4Y
QerlSXlALko+4sBbIyvYepfnZR/21K38rER2+8fT4MvJ7iM/q9OXBjequ6J/hPy2
qgh937fYh7hekA0xS2JH+ftWng9tZ7gd4YZfrYEoyn5UwDvKj1geO+dP3LnyFL0s
VtJGm//ii/EXuahkdH2kDZziA2KzwF5koT1auWx7VIFytaRSnM0EsaqUxGh0y1gM
P/yFHZlDYnGI+zefp7YJsxbsnpAB9V+DYJQB+H/v/HuEsOp+9vK2MBlJ93KBvnya
qrqN77r2W7KKbpzKEFGU+H3AamZfMkvqUOORz+ru0CreWpy3iAiS4KhuO9/+CEEi
hGRNC9gGJzQAS61bAqjM2vs68tNZECR10xuqntzNTVddh66clbqBjoqxOdfSs1JI
mU9H940ur6EBsFurLWGjKwGcKeuwQ6IstYyMW0B86wp2L8lAfDuRhC9eKj/tKris
UcPQsIffEs4XoIPZBTN5UfC5QiirIoryS5iXtDXkB3recuIYQOeprKzqvuBM9H0x
+edoXcvBq5iPyA/iVUE8AslHi2rjgeFlMhVWoYVq3Y6uZFxZps96pc5QqEbrZ880
kU9YzKPIl+SD0dhSKKbMNTqLTAaaRA1iuAWF8QJi4qH/B7ar/xyRYUOFb5FD1wXc
S0mK3IBp+TikmUGmxAg3CP3emq0ZTgTaoL5Z12zjtFbwuQdA6bpFnLQ4NFx7Weqe
2Ao0ownXbMfTmhrf1rEdUt01rsZwCNTXy//F7JCtlFX+2P9rJcnM7vj5zUzVYioS
luAhXdo2nn171uzcd0Y62PuKrEq4sfWxnCM2eZ7aXN9E3gLYcpsRjJPXlzyE5F0x
h4HVT/7L0Q9m70fg1z/ShQATluZDCNqlCWpXj+4upp61bJBAO12oNSlM/Trd30by
S+MzzL9cvyXVfa+JEgdaM2D2PFfUsECyojbYJdYx3IpH/HaLEuDDgtt3/ZZyOQDw
PTBBKvha2vyrFzBsm466PheYwxX7TAAGo2dbJDpxICsEGwOdlBZtvCiGLsnBJF66
QgHPpHl8l2rtwcMotfd1s/c7+b5mBzRsaU+KSxuXZTsubZb/zzPkAafGDHcHZQze
QcJ7G3OmPP04zprNAgztHEc42axHtlFfEl1KJDJtDnUQKW/UWkHHpJq1w6X8Z9nJ
r9ZIJI/W3nq+R5Lq3MFqO8uDyBBeR8FqcN8nKdHuuHrJulLP60sDN6uJbXon9EMk
d7mytAMFuN8mPbx+yXDkzQJifIJ+wXuva6debRBwvkZq0jbEV9hztJsoeOgs4rxS
W3eEC8L5KrHfdw2NL8kmp+qIOKtKAoglBaw0ZPjV/2KLLo8Mi77QV7tF9H3q0/bf
42q7cdd4TdOxMue+Stx2+aFZdygsdPSd3YeXz1iE10kLuZqAe9Ko6DtF5JBVzDyK
Lbw32BY/VeArXWNOsao5fS+DKKLMV1+NT3jiXIR19w7+r3mCOXuqh7SbBWNPmlSy
iyJ5fHV6TwN6VWeFH/tNUR42qVG3XQAGXdwA40kkNJO7jCnjGplhwAaAhSkGkkEE
R9ay0gNv5j0cr1wxUWKCWiJM+nCihXjkT3HFPYcpj2+EIB+jP5ClXVYY2hv1uwh/
vdlaVDp/F/WFkyrjJ6J/hPW5YpJicr2tW5RLBt1OH4dLptujtWj/BNsu7KSQPv+S
MjGY0zhEUL15GaFzFUvQtKxEk8hb8Jxaoze7Yx/KVKY9K9mU3Due/iPmihGEPOTP
oyfK3GOwzC87jPJMjyDEPDgu02wtC2FqYJSysHlX4Dh4jSEiECscImPoHxbrljwH
zLw0aCZjoIGSFnOCvEqb/6W7D87me8o5leolwnUBMqo+u10a/jbMzOerLLYgCqSp
EPgpZ9f1qkemEgHUoUAcn84UIQz+vXn6K0xEU+N32I19Q4DmP4XNAO0cs1oprclb
TAldgi7TAd4XE6vbYhm5zuLWadt/hKakFMSboZ0bTW9O7bu2uo54SiSzOQAtR+V8
3xwHBlEyDJegPtOt6MWIl0HuZwVcm28wSAgoogHNAsiEzCTbphPPd2xhC/GZiUnH
kih2N4cMpb2kZnSura0Q3V7qplHuot4r68hduCqmkAzCXfX3ZhqVc1KF7YwbBqH8
ejU8njingN7bDCRXUs7/GD8jvaj7CK4qmjR0ipWDMhZwUNcNybIr3+Qu7pjFqZk6
l6ajnE6iKPWnlTDw570ti20iOAL7qcVAKlEavJuiRzeFy1+T1FI6kZ9mPxZBSoA6
1JzDPBkqkx7zjoL2XUHPKAATcXMEyOYOhZ6EgLGi6MHt4ROWP6ZJ4vbbTH8AMSgc
4sTjVL3JmabMpNhtxZc6YkTyCZ9GKG+GM42/Aja88nudQosMqR+1iUNYdSzAypiu
pGlweIBIgYlJRCR5/xdjzTCGVeLHW4cqMoebyTqW5NRr/4UUsgsJttIGzZfLVS8l
ERBlojbeMgKm9mwlmqa9XTWai2+YvVkPfjJpjzKeRFHxPa22hhV8vJvL8nVJOQSI
w/36E/Dkgmd3eBWRK0eWPvdYHdcf+0rc3kLeim/91xckGf+GBkX526swDVCcvJsa
3Pjad0jZepu2ezq4kj/z62c97qxyh9lIrURzXOL8iG8+nH2Wz+w5dWr1ctGxYvRu
+B8Y0SMvCjyqCzWo0s4MXZtI4aTwI11/KZMPSHWJf2fdCQnhPhNq6nNy2b1lXWhW
NNn+4Iq5GKzJRdxoDXeDRtgKWEmKNQnJ/BpOG3Set9p7DPoTm2e1+r8oXau4qRLF
+Wu1Kq/MT+fLLeh7LGLEJpd3Jr39M08i0AYm89yzOC1HBAXZqU4YicRpydf6W5m8
hQSMDQXJtToqeJC/XtBCEZSg+5yv9yXJy04RD1HoTjgl7wxePnthveEOFDuc5cMP
389qFWD9/NhNbgK6pgI8J+X+0960QFpnpRyTp6ktprCUqnppJbi24jcc7AExmQ79
NpW0+Ioz+apjlPLBODQm4PoffHMEhbOKM08bzmIzZDmEX9SdvHodBcPrTbGeIMP0
EZzut3WHOhmahnB3MYOA2oZQSxb1Ng2XKoXp/Lw/9fZPB2e+QreFJGcpcLpBv5C3
Cfyp0E5c7aY3h2P5LTdiPSqO4y+M5G2Fqnts++qc5YpQ6A05ngCc+MPMsLFblJEG
vwy12pIE8clH/YUrejlY8OjUtKMzUfDG/K4HvEgA0ukYSOxX3lZQzCQOx70lHtJm
AteJtMH96Igx1worte+keY1bolS5gIIzFfiY4VfAUr2yYPPtTZSeKefsolOc12/M
cIJP/JBLk9ziuFymQhV9dv0FSaAybHokmcY6EnadlRGBaK4JGug8URVbmQUJb0PG
Aygkzn/Gkk7m7awboYCPVmzEb6aWOwxmSlZTUDHzetXP+OmNVbEexGgoB48yk/ij
wgxce8jXnEb2/qpQBBbTpRXyjUsRkReUXpNxV0pX+6aL64tGWto/hALLsDscSWJK
2OOErC0yDeEZLjDtcLfn9rGPR9LKbG6xMHiOQyS0qcycwqzKj7iwZ9r4W14QabYC
TqmGx181HlRsQfIDsRoLpeRMCzPHFBc8Q3kTuDu9ctaPnVzjRU+algzjqLDW1koG
dS2eH2C91VQNa0lnR7+qTMjSLCbyVFzOfgebOBxMfPdDW1BkTfnKaRu7CqGdTzcF
XY9W4wY7MQlEwJxUBKpKCUcd5Udr/pbXiXa0WitHtLJNJWvUqp8au+A8V3NQV7N2
9CkM7OagOp6NExId3qNiWCfznL9zGqDaTJ+kJSdbdGfAA1bHK1cKYP8Vr/2MEob8
ItQhaB/8E2Fn5QuhqBzzLoBJuQ5xxeAWqmSrumpAK+fH3v0EVPriIIYc1bkNNJTM
If/b8O8q+1Yc3PiiLaAFiYZL3fdmj6tgO7p7tQ0d82raCZkzN+9R96V4FYdqFSqW
X4ncZLSx0w7s7+OPUosy82H3IeQO2IVfYRVs666YdO1vd7E5FHCFYa4VO1btjrex
QU+VrtyIHyZ8QO92Bexwd5qkFS8za1i5F3Xf0ywQ78QjX/AFazPlGkGnhA31Ydl3
y09kqPbYyIyrzV9T5D8TO6EwpclHUqLC7fiK3kG6KvorN+NX3fqp3YUBdIsJEeeR
+LLTSt+VpUdx8iWSToD43gG6BQqUFfD2l7rUCzdV1Qq8vY49+yE4dVzmiNrh6+fX
8nqi2MYwEVFHgTPOnjj7ChB3DLHATittbEtsF6sLOOZjlK4psfuzOELthQKhSg7H
vRa5mxzr3x1PyQ2gS4RgAuzQWCh7B4l1jwjIGQScKfgJfd/Gjj+FvT6/5ZJUDTqB
Fl5Es1Fd/Zzfh9LZ5k76/gm1Jo6KzAm4kkMfCSzsKd6Na9ykLXPO2vqrgCK1iiPr
VyuBQNBF0mmBKwWNw17IWieRmwk5Qu6vNiv8OKIqE/xW6LiTE0hlkyqV6bOKT0Yz
tlKam7A2FYQfMg+xyUMcsWPyKlt3Zc26niBoUqStFjid+7ww7O7fd9Iwa+Syz5it
2fMo54s9XyFHJEPazgpbaUlB2/IqA+aaapqB+9a59NoVHvh5x0pnFnM4TxRNTuQ/
LyzMHfyOJ3xQLT5LHPtyF2PaZYyJ8Op3aY+uJEY94mp4xhbYRqmnsvhtKHuDhmat
SClqHlCRZB9MCbxlwO2OGgON3sS8GB2EaqH0bLeFF1hBe70+omQpSvFDph0u62t9
nWXG3K+gb27xIVv7BWE57IW5TELoL7UrCW0K9vNX9xKd8xxs2GFe3I8Pfw3BPsVq
AVJ0ShluReSLYGOwQJW6OY5ku/5DqFvl1jh9GmzUcS3QDuMNsnr97ZPZwPvnLv0W
prY5gYx/PX1wY9rUfh1lLwKIARfnVkk7yKFEcSBkjkZ9qYTuIf/+Non4s599Tni2
wxv/AwEvMymFhns8WCm2RDAjfTBEJvwc2N4r426Q13mcF2whG8b49FBFJLR5q/ee
86pst0qj3I+zoEuHOsbJuZqZoSzuXubjUp4upTbFrNewZJSxBHvNIK0SYzA+xXKR
9DJ960o+WXV/AzR/x7vbLSa9w0/QxUt/0IVHrI1D/2zvuunKA56LCGghImR+sIOc
3LJhGTfanGGiwraEsqr5RfSOO3NVlDynUXBMa1TQSqtID58KIBmquPo9a2/S60Aj
Zj5bBDejGXJgmZ/CRPfthNO1sQdOqD8dfz/vuxv/+j3FCVDdCbzTeYnPKbkzaI8d
9GG8BU1EL/1MdKGvVGbD3oIrVo6i3VcIPCxPGdsUuxCB1qZoBWTwgJBwtGc69LSy
whWAxge80ODtifMZLlfwevnuSUYCplVR5OJ1LDFY8RR0A/7BNE9pzPK5gWYft6q0
8RB+G3/BZS9qpFHhsrnfsQ8zpNF7hko5PwW8UVQ/H7y8Tze5B/uw5dH6203w7nK2
fULGTxN6qrWgqGUU4mkopE3+lIVeUe22XYXyTFR+fzEWTVpfnCRLDGgR9p6pRYqY
27kLnHLrJkAjmiRhBG/rKmzCA1MsUsT0XK0HmAGTheyNSoucu9MpMPrkJqOcutXh
07Oqk6gPPgMTHZJzKAUeIQZ9QIEW5VnJsKO3QgSRUglE9+ciVJwZGF5Yq24uBC/0
RtNDxRVi/6j/zMBtj74FD72n/+IRgY6fUMCBQ+vLmk/2UU6Dods442pa9H9qrhhJ
88yFCCV9vB8z5LS7+U78ecwJPtP/vdt6gzaZla9RXXytoMQvjikKr4C5hmFOlTw8
CjxLAp1XfbPjG2gQ3/dudI39oG9RFTkgMjRKXwpvlyhixciZBhQzD6q7184CSLcC
kwtGjW1R5OvP2lnDYAJgD3O5KW8TTh3ClkaYWB3AzGVzK9QRW6Tae+wIP9vKy9gw
bKS7hWpQ1KAd+hdgbrMNiMWptpCXyP2Can5md2/YPt1lAbCgyhJyrfQWQfWYgjmS
D7oN6zVM1uHHuRSQ59JUkZ3Rt97Krqh0Uva/CdpXMMSArj6iaYXxYruVavH2Ozgb
pxzvy35z03dw/DCCxYpR8LmevcvO8sflZZDXwywQSIr8fbkIgmfHD0Ljrj9QupUx
N09pAAlAvtIF1bXFe1seZ3VT3HzPZ5hZfTQcSzIs6+AlpvCkasNowRMU+R0MT4+e
bMc/3gzenW8EelWNskVvfZcSkm1cEkyj8vtLFOSbRPHOLDYP94ekE/6RMeuVmmvY
Y+SwjJgpCuVJYGVCeS852Zgtva5H3sJL7yovXEIQq8MVgB8RRMWoa6qJEWIg8ifE
ufOe2cnKNu0VR6+i6ztja2yd7wwARwVMV6E7k7ITu7q88tTkpFFRa3jJ2feg6sgI
w8PqPaQi0CZoJS9xkJkptwckYluOhLRTD+fNo3dmtBgnDgfkN1FUFDm73gtexs0G
LaaMDwz5uflJyy8FMkBmY2t5S0bF+LKvN/DynciJyJRk5ecYcAMBfhpflRT6o9bF
W2JCa2aqM4KC8IUjeKJFBFEkmLaHHTIdDhLDNDQKv61jR5JMSF2zDdjV7OoGJa9E
QrP8G2tSpUhzzaXWUMi0AogV+qa1mGBACPZqUSOrWVS7lw4RJyZYgeTum2/o3iTy
xCycOXnjkXptqYdiwwbscguWiEJYPVpML2SijC1XQpfC/E9DQVbVK1LcJNcYLFEL
kNtxMo2hzjChZqYtDxanVNJ+hql4zlBfbLRjMX4QU4PJIah4yr+8EDC3s4m9cY9H
nsSUDG5kQHGJZXHJvj2Zf1uSYJiuq0bejgYFP/kjQyQIW3mZeCHM1BykMnaBv9xd
NeGSI/Zd9w+yPphLso0PtYR4cuWLbDSjV3o545XLtJfSY7V4F6I58YS0H4vBzZ4g
Qpboyg5lmPimLF2bjoKXE3jWNMRM9P7nvf7WP3W7mPauLKKPwbQYSksCvaJrvXAY
680r9MHRzKxvgzrXrIm12A3ZGbm0vxCtk+DGBRvdTXXGoYR1A6zOam8I3NcsOxaI
HaO7tBs1PuZPGLM0keaQcfetNXTcwD0Mb+XbecyQkHZrcl+YgZXgqNzutlhog7wj
eDzNY1q+brIAF1GzA9jzDtFuMnopQ/+ZE5YstC/bTtu3+xXuwF5v7lwXJUkyvdlM
FOmPr5hHlWKbnd9D24I1bGhQ/4PcCTf+bBWZ0XrOtwGJbB/aNXzEtGg5e2BuyZSE
O4zoKbxwADO46jUrnkGV6hUGpFNYep6ej/aPxh1qRlnVSHgBjbU1c7lmzaGkrgaR
fQwb8SpcNtQF8+fGE7IDfq/IgXpSVBGWD5M9hYh9/y5ZDZK/8/DlAGmXt9xPygDu
hTRXVEUPqikFIDgQE2/IE4KhA3c85JDuOgs7O//u4qSeRAPNyyBiqmzNjS6q40qS
6jDOydR6t4qEwqmntoVegR6b8oorDpWUCOGLrw2X6Fw8XYuZ8kYz9c4YFw9coQpE
wJYrFoHjHumgHmakvX7e+kmwYArYIeTdTRioC16Y5FgEvmgWp8D9whUu0nwjnYG/
8nHsV2fphfSoXMjzZ8253PdHK2WgngsSLGdwLwhdDyCE+XngfwdZRVwmd1k4webY
GTRc4s8k06DFpJBjVc8S0Cx7G6MzfhNr6EkT7WGrkgFUdurLa1KQBilftbmQ74gr
9XfXHTEWwhw5ij1Mgw1oYAnaw6yk7fxajrq9O5TuU9MLVptwTfDVbBijBrZWh6GZ
0IrkS+7ULYnt3bnLn/ZmzEkqdfy98Gq8Ouk3B7j45wpGSyhnglpAXTAeBL14BadK
f1gT9JvMPIKcRljoJF2mdvIwm6mD/OxA1w1AEFwGoB5+NnGyaQDKPvZL9EdL8Wns
8Qo/VH01imGI+bXOR1hQdZAI3OvofNExXA99Pw6kW9WZ7okL70WgLSDstbqMN2NS
b3cOaDGVernGytRDJXJDKy5FnM0R9Q9L0YnhZazktXoGWFj5Rg0P+vHis5eRPFMU
lCRYe0beSKcJXiDFvlh5RugSiK9mHFFjipXPyt8MLkchJhmigGujWl1l91AzzkMM
83eI4ufecfl4ZV2v0hPALpz1L/MUyGA2PR9fVzWATCg1+/WNBErOZ2G00VCYeNYd
vOenIGfb/sBQMkRoFdmDN3NUfmiee4wtPR/B3IHgYvT3NJukIwpFE/ff8DdLomTG
gFoLy3wH/bDbcKj8KUl7xCQWXhFpVLlRScdk8KvZ8XpMTHogRxbM5TH5K2AknOpC
i8/W5wbLUYbHPbo4fH6e0gZ5y2k7RqZwuWnhaeGB7NErtaFh82e5mmYkH19QCE8n
HwXR4FPD/AsD8ESUVGXNP0uz9pWB5ISJ2ozPe0rDzKS1+/RQJqqPR/rE5Z6mMDFq
+5Wzhri+6j5ODI24uCeM0jHJh5n9MnEDo5ZXczozB4s71zGFSaGMlpxLjgfokR1O
X91RJYoDjlVq0EhCCpIfzl4LpwmNNDuY2Z0ro0z6hnTV632/KnUSPwqtgfnxvjvT
5VQed2s/iKf4JB6oBxwPmo0XcDipO+HcDP3mVpTn2vO3ZPBGF8SUEgfDyqjPLTMG
SE2e27C3/sdekRkRJ03u0k14BjRHewOW6T6uPUOPUDPfRA/sDy0ll4gnH8W02kcR
hWP528jBhqMruoDQdjfmWrGlvIlu7hROn2bFSwvLIWtMHxevvuCHk4QdMPxtbCaO
fT/73D9uduU707xaonj2O7eMklj4Hs9AKnZZp8PF8GbH+7T1XVVNOG/M9Jx09TzN
R8VkkFiwup8hZRYz8WfCmbovUUmg/anWq9QpechDp+WGrCF4QyiSG8KFM2S40pos
NjWa+n0Otvs+WYQtCiWeDoduvtFNEp2WeyUX82yjOOs4tZQD9ryST7xA614fBHHu
ImMM0Djb7O1ioQjgbr6XHEQ6c/dgD+9z4YN2ltaOcGmq0a4ABTaBKRaKw+sZrw5l
J/Cbdsnic4FblAZrbgT2ffZwp7dmgei0jl+I/tMp3Gx2YCUAMVG6TOJSiX/CNwJx
5NwFxUdpWh87n3zTeyVEMk0ElGKsapunHoj8Ry0Ac9BBJ7tLRJ6faNvWhFI/vMXU
d8nbZRSiBIixnnE66ORNICtcfmD1P/cQelOY7vrJOkULRKxmVOPD4WbrR+o/mW0n
bLW8wi3HPdbFFSW05D7fCchXloOe1vKmn/XvJ3PTgAKr/11Ez7gk1kjWHbCwGaE3
q6ttn7+2Ed6L8c+W5XBkrmUp1zBmID0K2DzwhQTHm3O5FJ8j1fD6VhLPHuWn+REL
4dED25ZYghgmY+e8gMJxbbTwPKzUHYCjMFoThfUMrXiBu/+6grxs7g5eOBLoRecV
9Q/z5nC6RZK+8EjzRRVTphtsV7pMZkOBdCjm3JLRl/RNki0ubit63hu10jwUVsBf
76ttmjZpqGdiojiIZqmZ+MrIlvULJXe/eTdJB3Pw9+xZ5laK7hAULrhcffA811BY
9FIhB19QgNyH72pZ+Cf6b7TdxP4Ui3uUjH2wNgEtSvmjs6clCJWmJCuj5tSevR26
AwmIj+fsSp8EFVJjhofPs17fdOMEnlqzqLYwp5F0+Tc36OQsJnshA79XL/0lEySl
sa5rsIiZgzry/cfqaATBuXGhKx4XiJJzsx8/AQRzcU9a+Xj+5FznLSzowYkTWkkM
sVt8EOafmFWSx2N6oPnYdD8TeE/60L4pKrkrf73qLkwLkWEQzyBRnWooCG0/htm6
Nup0Wbq/jOa9PJuX60nSkBunnrMpp3qAfCdl5ybU4SeAnLBSJVi834rn6RyMutqX
7w29mTJW7YDC0Y4qbRcybd3FTyYDbC6GfXsPSkeM6ko6NLi+ka8KCTu9eqVp3MnK
XC1f8aNgEzHnGHwZQ9UQ9P3abWbwJzsthLmQQrTvcCLZwQ95Uc0u0aypO88JxSqG
PgVTwRDDExj7LVASD+Kpb+ZIu3hTyWaD7h5PzEpd5ceE9GSr1ZkSJjta2fh5pupZ
t+Koo+LVtv585JxK5QgFaBDQkMkpC7/T/QLmAMYG1+7h+g4zAvvpTZS2w9b9WaKq
jurLzmRK733HHS7AT5fbYgmdmFDpGa6D3O9hClMuJJ1bmgTV8AYjJdzO2VSBC1b7
XYzpzqAkwfIjLhj5BREzbj5NTpphlDcgOccqHeDnfDIDKfTYcISRLyJUuQ1BCb65
fqJ807H4u7Ok9uTFPmCMswwsAvjw/8N+QbDhnqI4Oyj322umTPtwQ/EIXgJYZ+cL
xuhI26gZNfnm8UTdpfycClQ0MHcUnElDPODgaC3waD4RvYeKFU4HiMJERUwSURj7
XlLa5Q5nqjhtlFsdkmND6ymy20VWLQVtCqmYjGIgXDC5/j8eq2yg3h2VJCdIDMJj
ALuJrL81WTNLrP36gJX9EbWSOwNuNVqg1laP3JcXaPJsplYXtTHprLDzoGtlM8MX
zd4s18fvkcrzvIhBd+iZm53Z3/TKbhQ/T26hK3FqrJOPiVlLT3xS64uZ8Xel6xPG
JYEVLWgf5J3VRI7NfoLgYfqjY9HqAirfon+6v3Aq4/Rh2b5CI8Y3KG5LGQKgq4Uk
S62hbKTPx3rzhQ6iVgWnIn2Rzcmb2NkS5A+Oa5lqqIHalDSdWU9t6VYLK/yl2uyu
6UL2AIErVwFfdUO+f7Ps259SZyXtwjOU8Uf6U8Q+j0viTtrpGgsTzQk6JaqFMVmj
IRPjTUBCXr2SmCFyQRdvngCXnjsVHLnrmPRVIiG+74mhKVO/LozIasLyfqMNGbsa
Ijv6vQiRKvDyvcWdpegiawnjF6jhyjFz0gLejH1A1LcgomFb/J/KRACJ+Xm9y8Jg
eWp/VsVlAhu5ScoYIY+eRJhG6SYYgAV4UfFo8TzJi5/swcOJ7xIFgVih6hQYrbtE
THgmYJKUYI5wEuSrTTXIyqbdGCB3smuzzhHsxxSZ5uPloFhCgvUlWiai2kP3IH6p
OTlfN7gL3vtj7rwRqbz4hHz8itC4Kdphi1jP1AY1PojLzzZEuXX4XUDjbbCp/W4D
jAuUT45otVX58f2irVwxe2gr9/wu9i2HMS/QOhVrSds7zv4OJXd4E/i2pq+MMCNS
c10S5jLiQWKUWd7Z3TxKxDwoLpa6fSd9cdx50//BEXBmuVAVeDyI7XkOqgP68jJ8
EezhW6qSnA/02q++5CUhVpq4If/HIDNZnkkaeXBQsHLRZ1ZsouynndQKOrcdTV5P
0AahZUy067jwCZV2QK2yWvNoRpfsRwp4BtQoLYTjkOhH8EZzQQY+1DqloSg+aZym
ulhA2zT4LBBl+2wPZ8BYHm512Gim0GhsL2XJnC3o83/QXnwz+px+5CjFCZxOVPsS
V0PmiR+EKN8BfNPkU4+lyISZLY4TdxlEc6HYj49CtZUFez7cz02TsmYPOUkU5rPn
ktBOFzCEhmwL1qgZLGlo5jocTeQpE31jRnrHreCOxz+dr1d9OYkOcqFRnSdIoGfm
6WPdbffu4xHqCmAgvSrGxPHGb4MMJSqogXq0sOx9/wEjm32v+4lBoY8MewQWrPm/
9CKLat54uRKi8b/rRFqUgpaq4uxMTMz3NnpNR5RH0adbXYcYcE3JxeFNpLPuWBVO
YderuSYj9vWspUlUU6ZEiE2pzBmV7tChdshraASHVgnEkIVsmyQoLZyC49LmjFH5
842oDQguvJnGBaH5F9jsN55DT9ckqNFyCrrvdOWWGFOwG09JXaEKKmEPHwxo++hf
JSMK2eox/BZvntHUb39v6+yYa+09wkFiXbXLWLh3rnIo6F/Dx7gZG9PPNxOzVGE8
HVQN0UgD3R5zd19f90aFhYMq4KD7cLXyj+DgIEb7BnfNe2gG1lDF23BjOHU1JJ5N
dMfvdnyajujKvA+Kcs37UGqhlKeAdu1G0Rb4R7AJoktO3GyzvYunJ6pkR1m3IZx0
SojpYI23rBvWO7jlys4NgJZChtNtIxa6NgFPye4UV+bWkmmqJFHqdRBC4MGOWQ3e
xUJIbqOhEYmwBwtYA/Yn5DzApcpXVwl/tyMk8GHtOU6tN5akJT0O/ATIT+Dra7Wf
rt/IysZXVu2+QpPxwLHILSNkf1vXdcrmED7I0w75og1oJ+35Y/tifXb0s7i+XWC4
HMQf/fX+vgJOpQmdSJ36c0UJkMac2bhtN3EaHK5JlOmkNssPkYwq1+ZYnlUgjj47
tJBAAjSfQlN65ALJALP7RJPkOUjeoqs4+MZdcGXct4+ZFa5RwecLqYW9RTa04EOd
Y+8uGvXlBoDghN27YquDjxhi31TnkSw8KsjtqN2GVHfpCpUQVveX9LB7j3HJVDa2
9UBfmwtEtE7U/g1yQj2haCZgezaTd7GYe1xiKBAVCGrVNnlfdUTJsCIfG4DsxrUW
HM1u1as0vH2fpQzBxi6maQHGGnC/n3BFUG9RwqWGsXuFauVHc4jyhT9tKu2XiubK
bT/c9ZYyPFSAOOxwOQURptrBMPaW6cJikF/abIp1ZuLvgo35JcpG1jjrYTg1zrcU
/rPcofzdrmDj3Oe05uW1Og8yySOPjXw8y4BHFcPnitNxrZdgVSOKgFcpvTe6Myy2
fDD9Sakl9CGC/IfxelxNR/Q+X8TIY4rRgZ621WIpPxzi0MQRhqeJz8POOl0CHnkp
qJAaRQ3bnDXucu6edNnjaPQRN4zZD6kxxPAlBa24OX8A6BAM/7AoUl4b6mxwiV/O
+Fz2A6LBwCxFHt0AfjwrdiSzYbd29BswKr8/KSKzJesIuKQVj34e06QxNugHBpkP
Xsbs4o1/VUvkekew5Ar5F45RxtVIN6oXuzFrS/ly8LBXZluVYfII3w7VgwzmOyUB
VzX+E0hJ2nCrMQFGikRDHoMjlNSLbD3YgeRCvscD7jOrnuvG6Ui5BYSSn159GB8H
v2m65q0kF295upDa2m0TWjhdqCY/USW+JcRtCXtwk23qX6i3Kdzoe+jk62hAHVJw
XGAVVF9FRolNYBlEVaMQiwf7JIz5i7/oPNUu0doiTw4P7w11P/1XFHdJqtNp+qq3
KvGlj58xPzmnghbNtffU5HdrlTBi7LoKmLFWsgODs/XsHsmagavzrKIyBcUJqLPX
WwUv11KYb2pB40Tq2Sgcwfm9+BNBaLpKePJbYwTRlpyujhCM1t4zUYKqZm/DJ9ZK
P7Gnekz0OIcNHU1uFaI3nCAevTFgGmEl/jKc9zbtXtPM9x8cpYWZykY6sY0mk3LK
zc+twwFoHGp0ZF/fFSDFNso2bL98x7ctbkW73nZ7f3XtOQHb/+og7LGdRMLPGtC1
FqfgTqhkErA+WJKYBIkHEgD2CRHT9XG6u2gH/f2uDzLkexC3+hVGqD3kPLy09pPB
TLMx8U8zt3XoPgD67pA4v/JDSJJO8SYKX3WjYuGiAX2YFAOFeQz6hYc6n3Tv3wXh
9xb206NxaH7eUUigpov9odMHoLDaYrjf5SnA+qpX17rWNRfULsOtm8G6gH42ptUD
Qhy+J/DEFbTUU/01tOFil144e6M83MQNwH9hx4U7TzdQOCNR8OVuPLpACyMS4kTZ
nn/CDudbqt4d1gRmwt9Du17SOA501FCOQj98B6/V8Y9SxYH3isP548v95uaeM9FP
sN/yTZvuhTY4LQPAZax6tu3aesK7AvJ8uxxZ0d6DUT9HOdDuxRS5m3m/bQY03OEC
tZiW19bL3WkfnSn2aTqF8WHJN+SQRK91fAvRF36bgxb+E9/KZGqpWyAEc7sTamsZ
zQCA8VMDEI9monKLlaoLJ4CkGn5GVd0MkhUAlGx7ff14f4Bi2AGdm0MXQgXl3kKU
SKCoQMkEaIp4nTqynsLWMyuDdfUFxAnwkzicfIoDKYPteAQtgi+bc1zPy9MQV3bq
r/GooCQomH3slZXdriUnYwE3Q1ENBzPGjO/MInWFa+C+pXiwTqwKMyOl9BMxX7I0
5KqZFy/3nRZnUkwyeO6ugKgC+t54EuIQnNUa6X1SsocNuRxvZz5m2s3Zj3zYFiOx
FlBSh4/zdW5xYTbh8XJw9QZEmnbMQ2J+FRgNni5WWKx8EyXDRrzTtCuhAcbOFx2O
t0rziqfR+PMcZ486/93pb9eFIhScYUTIohEBI7Pai9yjx9qnjML3X6AlrPJlkyQG
ElFbseDkRPCsrZWMwnsKHvYb0CgMbMmQNBSkC5Kt83ROoE/mMMI5mUlq9Mdx/YOU
wNV7Mw/tNfIKo7RF5NEJ0g4p9XP3hSdSve4sSpLQ7XHN9QZr19ggsWUdbosd1Qjr
Ctpy8TAn9iE25Xvgxb2CJb8zL5Iq+d+UMMWyGtQG68qdTEfGoFAoVeUsC4GY8ivk
5Pnk1YdEAecg3KAV0UHVDNKD9rf3BJtdbASWirkYaN8CzijVVYaJ9yRUD3Y+nlGG
N7L+vLOaQ7bSugb2986omerjCfv311zxQrwXb3cHgbC5JPA0wJIAp0McVa+bLD2W
q+7BxV5fw6kf0A5NSvAUXE+wWS2vO8zjaBSwkDQQRWafymm9RlF7eMr8avGV0L0d
Ab9SACeXQ/rnyE2W6wc3Y7Tk7TqLnz04ZnwbH5aOkK8TdheDAte1rgNqXvmQHLTL
3vvMG1f8+/d/uaYcMVrcXHnaamKAquwjxZJdnXpHTONAeUCzVJ40sQou92zjghSR
QQXPhBpg1vf65FOKawJ/uhUwwLrCupiwJdYsfekowsAAvNdzrECAdiNO1wLi6yq0
952mRhHHP2ktYtRets+3FKvTj4s3Zk01SWf5MEtdruQ4CQMEojEduVgFFuBvU0U5
GclVNPpslIXLEP+C1h+iG6lkyslfzs6LJaPehU7R9uxdq8tQmLQLcETXRjc6vlxP
mLIAR0nEjEfJkkYakjJLJ/PDas3UyQ3QQdil8LYeUtHEcFiT4rgEBbqS2ydXzOUd
iYmauYbn4Hhl3/qg1rgAS73xzREyq76E2G3MQ3Z5RL8nJvEXtQJyuUWnEDQTvpof
sz/ST84/w5ZVnpB6MXZsuD8CFFxRVlnfYvt6+cKHRg3cLoTXMXlnLlKnH5+1aQWn
0HpKPISLU/6LrBNB+jgoTECoSKL/6tVCw95bMmlU/MWnhQ3AvTd15PgMwde287ph
p6/xjfQflDAuSzrE26wIwBzFORsLZCqHHMX6PfuBj876cH4VR4IcanO3WGNJg1pa
PVC53xZ7Z/baSo3k0V5LePqiqstwK2ljpqNtgTucwD9reSAmwhkBtiCp5hWGzXqF
MkwkVdigkMaYGYMbpG9tgyFgBpXWD7uJ4r6Vi/KkWDKZ2hfqhErEodwdTWEHKecR
0MGJxdb0TDJj/2VmvfSaa5YR6aN8/1iqU+KnsDUAfgzrefzF+F0RZVsklpf427vv
X/JfkzSondGunxtvYU+zI8W+l/4F/eWMv7++VvPW3b03DdjH6w6VMctkKH1/Otop
dyq/szcbSg0/YAS4E4wKi7J/vAFZFgJFTfTe78yKHlktFbzmEwyV2ciVH7Cs2Bdd
p28VWi1gLsgkfYLnVcZKY8QETg/mScjW/eEAKCKPqHNMPHKhirF59JD60AN7pFea
26ZFsTvBn/pRfbkPxaeZU7vD042XSC3xcCQ08ywrv3JK+Vo52kSW4eSbrH3YPgQN
7IYx9B+u3rSvnZR7ZhzXGdCAkt8B8h3sP1gv90hDrS0Gmjj3Mq0kd12hp225Uy5N
01VmKOvewR3i0V8gRZUJjjjNcn9UANoqiupDneRZHqJyQ54JfxyKLL+OaXVo26tD
5o+C3Ztwu+e3ORRKmBHovAvyn5qq00IDWbZXPQdvws7bpkzmLx357Fre//iSFXgT
fBRE6Wvu17JQNYkuRoBKoGTdiBTdui9ACw94rkf5RvuDffqjA+roAjx/Jrbuw3GG
cjHd+y+gs5J1YRkwBEPKZ07dZHAvBSm2YhTAv/Nfp2tRsGbtQWTG6NuH+CHG9Y8+
fQ6CT2XNuRXFyiAlwcXPjpPnXimXbUEb37VsKnW5/YT/mv1yLqDUWFu6Qj6SrKTh
rp6QG7SsLiUxfCIeBp8yzr62iuUAeCBhljLf545iEsAXe0ma0vx4sdcGd3FwLkaf
EWbpsS8q/3aooqKvGcMhulO0CDSkW2MNMujHjFHslFLuOBaQSuP3WEceVSgQKiM5
nWO+iPEekIwJIu+Oc13GaZLSIdbEJl9/tQi71plCUG3EK8dWy7k6eVXMNwm0GfX6
o+m0ReV8s+5JOR8hiAt9tSn2T4nx0iddoJgp3nb9Tgm6TrbHF2LtQeZzZy9W5LfN
3F/qgVoubeH/3vYshHo2CJazaZq1Hx2Iz9GJXKD74H5oR0KFh4kZDc+CofNlCAmJ
07khUTSrHvA/WkdVMfqr6isihf1AzVP5mtd2ecfzoeQAZr/fgEsDUbM1ro9nDRdh
M5ytQkzdYijqojgwO/E7bkfz9AikILzKVHY1rOy02ZWLIyAlHBwvdd9iOlsUxffJ
Z3UURHhrRUwahN350tE2HJ9xHIlDVKnxpDCDFctpE8TS8jWr30uO+vstWPA94iWn
759xcDjsiYKa9UMhbcmKhD4lus2Hf0DCrSNTfF4HVA1ituCVvGcl6yFZTZhEl2Vb
Mtpe+Kq9IxMiWYxJJmkoMIZwght57c30bAOqBp/iHBNw9HtIkCzm4REwUcWgsttK
916WdNTOp1DFqDBHsPeSnM4TfMA86gd7lJWJfOkV9uwqDPJoLrQTXPj/mgHhAsOg
ejpeSK18yCtolvdS05jNT19Wy/snXL2vcmO0/Q6WeYyGpMfxWqafw7sq+b8wdykT
hU2/eJ8xQYxW0WGFIFdm9hQlQFGrvF6gpxvAMtFU+kNmk3j60C/sCYYBartlbdJD
uCpxz+tNYTTaN6SDkNgy3V7++ssYmQaIfMn0TlrWXn4uYVkzN1vOZv7r90aKUj6c
iV5CB1Rz4MjYyQGv1cWMULc8RixIOgjZfQBI07qciBrSzjiXVnV0IF2unWWT7v5o
+Jsv00MvQkgC2U25jJOo78QNO56YVhZM2nhcy6D8QpvsKXDPqF807Jd/3UPJEAyX
CRwORTx4yn33VIsSOqoVttiNviggVq+eLrUrx2EXYWy051R7xM+BIofPVDcGnN/K
d0tXRimwRfcmnfl8pU74Tpp7EfVfDd0NtbYdNtkdbZpDl3cjX3d7U+Ya5nBklfXc
E1QNDjXmC03/oP2COd5CzH/F/fY7iPGfLfGICyariZVLMEkb4Q7aWXf7jOQ3MeE7
2lrBe2SZC+1SkNyNfUO5ySNj7a63UIa5Mt6Ju80yJmi7+EiXatpX4Vqbq1B0LOqh
7fylWJAHi1lA4qUkajhHwte0Xktr2MMB3/XPb7dYatauYrMrIW2cqr+jXBw01euP
GsDCMQe+y+lWTClbmksvyFhzcrBdFpOGs4J/buOsMBLSVPRoOItsr/lVi4MF4+ys
dYcrKWls3H6Pf/HUY7kr/I7lW9SZBWJY5JOY7d0nWhS/zo6RejYWPDtNCn6xk+gK
msE56owQ2I7HSsBIy5DcwQlbLYLYZ0NmYIFUBlHQEKkr9Cduw3Xox0mQdOouVbCk
hURbFP3jLkPmaM4PNkHtSoLmmzZbz1AcDjJBmndI5asAzgYfnU7QE0auS5OUaK2m
VyJAlhPynxD/gPCiFdJuMYSKglBidpE3/tPfYAc+OVF5nssbeDWaamQVg2GC0kOu
gFQ6P7d2B2Jsf8mSzeudHD8snt82Zc3jHOxLLJxCqbpWB41RjZiwThaUiQ12XP91
91prSlPUQ0Ld9KCb4V7bDJj8DTSIKt94WOVz4Wbjosj+FQPI16Xm/cvEhKuKvJCN
NlVxK7PkuGgjo1RXYSKpocR72Cu83dFCI7rnK9T3iDm6aWaOHsSPHKxMzupe4Ya4
BY7evh/xRlcqgBysPJE2d6pkiHP08DNNWsZw/fdz7GKSsO48IiTzxWtjlBsWCigb
rtJZ6D06VKCTtebPND7IMeO4vrnTTVlgGJ0KsbBYFlHvrOXOoC7aUSqlavGxYEep
J+6mOylNoUKjCbJHkOiJ4jkE+yD885VX7lbXC9mqURGDY/rLrTgWrQF6CsMJ3aE8
ygECa5NaLi5avk20RCxqUI7f2G6qNtbz3a+xuaeI6L2X3D38fpy+pURe56IJmyJq
DhJQFKa7gMt+0d2tCeB4QqgUqT8nTnOJcalHOU+/BHxTEuNj0VtTOqFnscncMbDt
KRPNpWwMlIpTPNUCxHqiUt6RHrymr5BzpONvoxmxpV1Q992Str4FmLqR/VUQdzNq
RZYrW3vIu0EbH0LSZHISQ6/Y7WsR4Ktfo2aBSWVSyar0y0KKSYffS3ymIOuN9Mj2
fP+YqgDYr72b8jGvL8vpeQocPRlS2X7qGB2rZVhQKiYA9H2wGOT4Aype8dOczcqN
0up/L+qIgkDWr7RL26YOmS9jnoxafejv4hepxfWFBtvKKichwPPWDuHeqvWW1UpA
sjDQSgQ9d+kXookP1nPYyXstJ055WX05dTpgy/aT8+iMIbDfYpeJDc0NTmDZWqJk
bd6+Zrj7XJC7X+ggmU+KyrTF8+zikyTxGOZ5KKdD+pTHEvbq91ppuEdqohOV90Vf
9VqIzD1MgqT9PNephtVxxSxBXkDd+aUug4Wv5NahvLnqSeykPjIeQ2fkKC3LPukq
/PHsIB5h2Hj6hNEQMCAfXYkcAb3hVzs5Xk8n8EK1gLm2vNQNmSw2C48ayrJ+8TNd
oZA9cjvqXUj1fHCCv5aq0wr692VeTLQccFnkohXWzRkZ37ecwXZoTNfeJHqTrq4I
otCMBN38jEO0QQJ49o7mgvyTiz0LohbXeiFzJSm3MEb76vEjzEQXSOBOrn0bj/W8
CBsF0le2jGkusxy7FTkCtfGiFo12jGsiIIb430FVgDb8AZ/5GIesKu7Q2DM3dGRI
an7fJcc3WVge+LC7QDnsKkZWC7vyNYP81LHn7D8A+jdV++BSzubDhXyLxXnTB4/H
SreHfDcyE2zMme+dNKc9JD4T3OfKXm0K9U9P0LwvbiBTqxQaVMRHnJ59l+lt/x5t
Jp271klnnPwuWG2Pg7qmRyv1tiU2rQMw2uXyw6hgzmM3aZ1xBaFqu5u8TJih+Ypr
AsiDrNq/iaZI9al8w/I4hPA7QxNb9YOubwEdKwl0FdhBHXnuoJAioPcLZnp1F3X3
qDDrHPPyDq59synQTYatcHLufHHz8wNN6SNhdiJvMXME4ZqiPxJvmfzyJRs7Qznq
++0zpkc37krP106REYabRVGyytB0zst/2oDq+fcnojRp89Slrd+10KFjm2NshEa1
TyzLcCXWpiuWmDQQhifoJWXZtKrcCPg/RksefD54MuCpZnJ2M4BQBvgmcr3WeUKv
YfhLYfW3aBd50oclJ/h6+K6k2aHS9zhtrlA1B3HA6gfUv/VDfvPWzEFuGysU5NS8
aAfPVac9/jy/1K6O1raRmxkiyLg4XAkwVTvEjwJiOLPB1TqXwOOpbyQhpeJJL4+6
qn7/MvzJKpF31AuEGyqRX4iYIT2o5xD5AsIDBLJd9GBTg+ws+2bxhMXA5tPjRpxl
CjSxhFmMFNP/PHvY8lg89knvlRQFWidyqZDD8WWGsOpoiEjEzAEl97HOzP2cO7D3
2OghKOdYmp4gyr7olruz9BllTJuoBeiRU0LStVzhWJJ/WT6GQjVbWvLUvPTaiPCt
iAVWWHFm9tGfpNJGQVmPfMCUI9Znx7k3UCD+dj/3aTYqodmY0kmtgj9V3gyPNG0Y
vEJISaFgW2G+gNK1S7uIIGJ2xWBNnoebwRfVKY0JXXKeXY0K78l+V8qhoePTQnYg
yDL/QM+KXbtbGknBftoecIopg5O3t5Wr4k/K2R7L9EIh488fe8uVytiMZJgZJMxV
R8haYRVPqKniwW76qPNTih4ehroN681jTGMVZ3k8nan8D8Py96zfBU1P1Aq8qjy3
aRYzxnJzEIcHzMxdwkH42QzWOlbqDbpBvSs2GbgrbfUFvgRgD0z1BJzE8UXIoqx5
pUdnAHPFTX/roV2+HSv73uMUNmpFa/gcuUm1bwYH/rhCy1unmE5AAR/ZOCsSy1Iy
0qReCYLsvJERNua3df3tXa0t6Tdw333EjEXe9hmVxYBSUmbXKVY/oQd5Zi2hyWqZ
8p+Hj5NwJg+jsUILGtnlIxxiVBYPCEAoFsUHfWhp70JKimQ1Z6S59IoD7aWoLVae
7fqfwDjsIMAhfbBff5vO09Uq53xq2wFwz2+tdtkWSpVUbjsM84qagoDU9yjrZanY
sDbaY5EBQ7IftECAJgnFfQS0qajXbP0um+AdK2rLdNZ42bH6rIOCiI4Gy8/5z/oV
nwePGYXpBvTnerR0WFJb+P6B5b8JxVfpTQb9u4RiczXxAUA9ZGvhQGflSebz7oAt
rx/4mM1OGPwlqOOY5t/cVdjX1vuviU9KRFmqAOOqZ6wVOBiT2IV6AD8jsokwcq2W
msJ5prrnvviSOINA7IxJGffWiz9QWG/e/KYyNUAEPoMuTTfUKelnw9yIH1b0Gqf/
QFFFlyGzO68TDc4EC0rQAxEQqQzBgmo5uJqZ0QaWwEx4rOFUR3adA944aYpEuFdG
UdBqudrvfBHqAnakqZIYoj0vIbELoycFM+7MyyM49abOK+EJKCjWkhEEag5j1Je5
OVOkLz1FO23ljDTbHdl+AsrBeuYTA5G/CXlEQ+39yzPx6G4xlre80d4WrhWeg6vE
nAHVfcTK0goFbtt/5P1d9a089yP1gEzv+RwiKugGVPAHUem6i3w9aH64a/SGvH1s
2KTTNK9DAFv/TLwL3owWe+ut77XbYCMAo7rqan2EtaHkMjqU/XRfDRNabzdtsq51
9NpYPNcjy6EECiZr8Wr9Bv6Tk0a+Kdp63Cz7v4dZjUEAn7ld1YhVH0IEUItkXxnh
uRe4uyJonP8EfKF5c7oABu9dS7FtsDIrbU6TKeWbn7D1ExYCTWbWz7tzrg/1ccZM
Riox9Ma+yJwzP7E2Q6hWHGxBLnPVGMSXlc4IBPgldAd7nIzfO10kb7QlGjz8pQ/B
gw/A7mpiPeAFA5hFysXr4FJiGER/J/gY9cdRrBblRk/kWq8VdvhyFMK7m9a/ZE73
tBCgB0wDw99lgfr8h0UfSHGfxyRFgd0Ac2P59j7pJcigaBQlT8Wuq6OXr2dWMTS2
6x/QwXnkj+U9dnCgqV+yVmW0nV/7GCvUML9uaizHEycwn5CiMPR3DyziGl9zkgD4
oeRYC1b7zS71F/eXbWyX14c3r1XkYfczBcW27xe6jTz1gQNd9n4TU58ONRZfeYMh
uiodcAVn8n/oJLIORkGy5VCqtXVTW7J/dDIpf7AD0N7EqYMzmni1coFyLI/U2dxk
QkbgAuQISUgwsg9CBpNbWPvg9DK3m/3EEs9Ul9X4BDRB8UfPOqOfSaluy2yxpi6o
xdFp1OGPTBI+q9SxskDeML+ycIwJcmQW64vcaH1UUC4kP1Qs5NWKDrMiFzqMIntw
EL9QaIEbiBxyKUAmrx7ekA3VBKIAfV0SEKTMOKoVs7dBqW9/ZHw6ix58iS7WAt+J
toJ/8eTD6FKHLP+aLM3ac9J07a7LxoA/6VzGTRaZ8k2udXvXPBMPhpGDNgATpf99
b8k9Eoa4jagP075b++r5ZYZHwu2Yeyim83/S5fewtsb6DsA4kuC3Vs+rOL8Ygc1c
UIJdnvr3OQMHYy0lYTltKBEWnJcFstuKbk6y34lcFuqdLdT+wWGFW/nDagq/qGCF
zg6R78ID6+C+xAuUH4pI/C/Id2PrJGG190mynYUezwTs5TxR+PJQj/HMArtko8xp
2R7J0YZlMTeO9q4aYYW9oNNtJMdJpKUD2TRg5l7YqyW1ffnEnY6PWGu2046RsvnV
VzDq6M66kLuvt7WEoNlpxY1e6Cps7jdyMXKYp7ssi/WVqVRIF+DRUJYf13YdS1tK
UQhL9slOaUIW3gLuhGsfE2f7lWL6ky+8kCmp/Nlh1MmJ6CyxOKosqsg1c7v1ib/d
asQXAghijbkBv7V3xch9O/z6fo7QAC4K9d35/kCrqeBONbec13LSN1wP99U/tliB
8d48E+4b+bnKhEQtxR+hWUD0MUo5+GCKK7mA4HlVthiQ1rccG093ZBPMkBCaGPgZ
CHtm5KDhIdDwAnjisC3FlCeA401qKDkFZqXlseOS8xqr8+JW37p8XDAqe1e4SvAG
PCK9d9GI9grkuGN7TT7Ng/cO8zpbRLCPewuLHmkFY+fe3qWTayn+h5MuV4RdxDPG
fAeOARHOe5U3tfpQD8H5yCYe5E+ZNHynlNjKIYL5Z8CvprguVqrw4KkaNYLH/r/b
24BdPVU9Vn4tQYpeI4OaV4MEka4CZA5V3aX1a9iKGD4ZjWiXy9USgeAOJtbee+xl
P9mow4j7BW8wuyN/JK01SyoXPhecCbd9uYkFI6VrpXW1E8qg/qvqbndEBvfMnElt
KbTGHNTXJ0LymARYPGJQUCjiPLG4sCis3W0T14TnX8o+uX3d6iZkR2hKAivbzkfK
Ijr8qKkEBfV3OdeHs3I9Y/EuZzcK0YCeqHw6PrKMnal5CzjkJSrqCn5LST+Sbhoj
gxg1PUYUOfnw4ykEmbaybmeSFxAbJZY5vTQK4B9JmWGag++gsLnOYhGDdf1HhdMB
WNO+3VnGI/RvYfTKDGcXVvfYGlrN6iHmcIFg2qTLK5Sn6fJ3w1RcY2MJdCSmHeIf
uPhyjyR3IqOxBTgnixQTPmsAl0PzVcvUJFuxanpW3BFH1LlTAQL91Js1WLTZcmGO
bgPL5Gw8P8jgPoXDhED4I3268mLM0qfnZ1rpgcwlBhnPfl0sHVKLDYG9FQf/cvLg
qCYD1LsWqcdvslDPBQ3ERNQXVuE4MmDf6KBRpR8fpjjORbI5McvCbJfGgpQ0kOBu
a3FH6GSGIwrhBw2CTMc2mUQVnyPKApBPeeEUXgPhxFz4WsshsgpaPdoYv5/PC/A6
vuLcvJ+pLthbC0S+T70btMeYHzzykvqGFTypWaA8jhqZjxoRlmHG2e1lXmts23Iu
1GAgf1ZrbVZDKWYcr3mdwFB20U59NeyY5Gj6Wk9aUTO/WRpkhI6LxE/UDMVNo2ae
UltzGHpQa1LNzn2sf0aCKKl/v9y2Orr+2IHoXbMKatU922YHaJsw3GMCO+rDat4w
xB+iYkNOtJUDsCrA5HmO4nJ+iiMetXcy3STS8YZli1Sk7/Wcnzo5tmWEVMaBR72f
XCvOebWigxUpRSqxsTx5M9QNELYOi4fYQmOOlE8rJxi0XeOEJvlS70npO8loLZCd
oRo6yvArG1jiPoPTi94EhEtuAZ8w82xvKLT9sY4WfiF05SNbevT0uNxFTY0PKBQk
KP+hPHFCCoCoeFe9XscdHEN7iysd4LPfz4JlzdjJlBLumt3rLxHtmmPku0KJE20W
YmLjw+7Q4KI0sWSkTsxDwb4iYWxtgVxYj93s3j2I1rAQ/4GnWcgG+pJ+S+Q3y+EG
Kd6UTOSqTrkNdz7hKXmVQk39hmqdVmgztgoFZXpfPLxfRsbjiNVsXNvoZ4hoMaeE
ugKlnoY/iQodtlMwZrgEeS0JRJ6/KJApdv8uIskN5yIinu2bGYg7b2Ctnz4s6DlH
HHUK4nnsDk0PUckKFuggKuOmyel8Tk1MnwjpUl4oWKBd8K8bhMhJnNgwVDR6StXy
bKHVoGbiL1Iy0Jd4QYZz3unSkIWq9cv5j/gAcKm4w+bF6fPJr1hb1atohk4hRWO7
IcJUsJYs6Nr+xOP7yDH+/lkSZF0au83vyPEozwDBh336lV6FiSKVkGPrVsXyMT9d
5/I2OaeWaBJYgfSrVceCOxAVaLA0RK3Z8XqsqxUE9WHxWerTLOmjJVIxzAhBw3ZT
U3jjl/yR5TbYBUSWjqQusbJSTHmjPBFfbb/csgLWL2qWCk6aVshRDs+X5BOTQfVU
K4vfrdEiPIuYIDs0/ZTxCyzrl6vO6zH8DuFq2BGhw7/uyfjbzvgAQ4mEwWlpTo44
4EBDFzO7Jj3z5FZE6XBDiD4ch3yJQG3IvmVg3hRWpejmS63WjuQFwH2Fl7D3fp1C
vbf502MtKcoi8SYiNF8RKKZkl/IkCyyUolsh44SLlJPjYGE0vrlt4tk8D8KCf9Io
mWRs7K6SJrp0HOtwMWBAK0PLhHjHOu3CiBG2wjRfyDQ5pmhRSeTrlFYayplXtCKy
uyCBddRc86aC95hrH1e4SDu/LYEUglFXfyx8oHlnbVLbSqocL6sc2t9ED+DUyE75
Nngrpeltile2mQYYvM+SpHPDCwq7PKhk20qDDpLWZZuwa0UvuVjaGXzl+ZIc4pnc
PeJKfQkCl+lqjHxGYiVf4iTOUWSmkzCoGC0oKXZ5oXCI9QOq0NJ+6XP+0JN8JEJv
dby41ClRFtJfVp0DdITeNS91uDiJLMqyBmAiODr86gT7KAEKAMacxpQ/fx24U7VD
hQP9+3jAxhiyGj9QEMgzEoKDAbsUvJuO4TsKV8SpbQ3tkUv7KUbPMuPPTYd9G5S3
YJhC8QQl6ujwoP5T//wG6DYSbLq3jtSSHCZRLTdmdndKbEkl0YIaj6mPlW6+zVsa
WZ/AmDDFmv43Qwge+vaNd9tAznOZ+rt8IavxuqAmTB3X9WWiZTw004sRPoFuK+P3
8xiCekU4jjU4bym2RBUVB1uPOm32a8e3I5VgSKG1gppRHMOeITzBiFD8qxZE+SL+
F1ykYdYhnju+IdUzO67OvSz308QPaojyrLonKhqNPS6oNbYk9VVMwarVILd7Lbcg
Wyo3OBjDGLdyDJnclZGP2WkwOfYCsjLSSKqGSBd5XImp/j0JNUkWLAO+NS4j+ydO
YZZUMd0NnLjrxeDFG0kXWH4r7ebQMKyMV+SJ6pttLwcUw1lR99LfIpIay0w7zxoV
0QcBAsbC64wTqd8+HPwku9Wf4Wcb4X8Uo2wG/Funf4c5qU7E+v6CffuPZqh1BCYb
7XJH9aylHB48bU29sZqPtnNkjVJDQWhye8Wi8lbjSs50LPey3F1tg0tMWiu/fDx5
ATwoAspo01coMdQ7b7Fmc4U8F6x4jsuuZH33AcAxQpb39cZ9ZIacZRdhYWekG0v/
mJsKL0HRvkLCVeBLM8Hve5RNDj2MerNqvUIClHlYHeO5Lc6EemvrsA77VisfQpYr
1ACfE8lfMOhC0bqCRiHV2hLJ5CNRyIeybcmNN9ZXitdHaoNNU7Scl3yXrMZ4U6yQ
uwlQruTeIXULuqX3hydK56uPVE84hQs1ipWD9tjWwZXqdq55tpgqs1XlmIK5nrTD
WWijFhvEhpADmpIpezy1R0ajUYlNybMGxc6meI9Q+JPfs3TU20HXjsfmTjuLF+qE
zXXWhbp/Bgd1TGaSH1vJ98jZMX/B0xayXOQx9JWSx5yzS7Y3kSSc+bTb21RQQnAz
5s/r9xfxONmFdo54nOq9InOzSI4m27DDsjRSdP4IzF/eWNRZh5uxbi5EMdw7N7Ld
7QJRw3Ie+K+CfqfWgM9Riam3n6ssDLkYR6yWVc1mzhifrvvdCHZF2iwrMXmPLab6
2UBMTQmv2K7pjMKAiqqVNbXEUI0F032jCW0mKZMIPhEeUHDeFmxO/sHG17MV9+xK
Onv39RTNpRYI7QBrFzPh47HPuzf9ChUGOKQwXeGagqWNPKyiXrkqfo8+ga7YFxFy
6YLXHiuYIqHeI8Ar8iGUAM9Hx/UwR9cT+aLPhpMc7q2ZirGJ5dkRfl3fD869Khg7
xmWZPtgTUlPoorY0J5SKQ3b9goyXxhucRixE+GF0leOKhXjaxrVnkS9JSBtrXkIP
egfiBdP4RdGD5Wb4bqk2rgLjSkOvjCgN6xG2gej/+X5NynHbZSyd/oxRPW5HJmUx
MtzQACHdezVnC08LAgvK3OGVmlo+z/GFyXGy3KPyE2QMDWwDM18HqJB0i8c43Ukq
5kBK8yMY7lhL9LHE+6r2//Z1BtBQGVjAKBo0F04HcssQzdLKCZeJGe20dhq53s8/
HD35psASmANvPhvpl8kY2Y1cIC8oAWXEO4VaoxwmlxrV6st7k78VrrHssaZ83YYE
CIUJVBMn2GR/Qf8GiFBFjL6wtEFutgdb5uKQFXYDqUy8HmJh8DxP2fZOZaDXIuMz
QHF/CdupM2Zv/8iQ9VCY9BrECNoJyM41O+wkA5qNJCuxbesC9uL4M8kVcQ1mqdKI
qbqBUm9p+1FFoHY3UMH+Pg9b208+LjAyR6kbjF54Gg35OdCVbMhqQ8Rm+UAzoRYR
hyue02S2O/PmE6doAMpncInlyeMTEM+eDYa/5f9ny5w5in316GHFyIgS2p8T1DsM
nJiuS1UehJYA2Zn4cWP6Yx0o3DOeISd5gKDfZ26Wfmy5FMpTpxkUfPoV8qBpWlxo
knR/0FLkecmNvWqmyAMq5/BlhKPUT5Ct7W94myK+tulUTDFTbXZwZtZPqlEHFt3C
8bWkApo8GmoUw1E+q8OlGZczWhjAWqYwbfnHZC1xcGyUcSffUa2B2fHpX11oGufx
jfzo+GJuC4kxuI3ISgfivm6U14uGrNQIG8yytkhZWWuiAwgQOB1eH/V99bxq59Ra
wWszH5qFe/R9Ne48ntzJoKS60+sxAC0GO+63wpZDIUZe4+pzvongSG7mnUGtunWk
WPbSwXSEoiCWZtLBr+0l2Bjl79a5hafJUcwoYtmPwThK1NBGUILRBlb1L1QzoPJN
j0Jk0hF0hJf1kU50xcI4JcwVgMkv0n54Szna5sUI9wo8DhdLlD8SnkdXfiutIeyD
AfzS3kbslqGm+lH5C/oKxyvvJv7uYm0dEa773VKha+qfzam+d3UDo1ASEJXVO3Xv
sAXNqeCrt3lp5+ZsJ2KilC+59r45kGS1mcTsvVGklOK4LQlOGoqP16FJUR2/2dJs
LW4YmRJwHP1S3oXSLMmcvh3+/KxsIZUiXfX2yHN2xBOBmLKfJ5oAyhdu8ijU4SWu
Wb3Xwgaggvx0KPKi3qfpnfDWpDsFPHkmXUQM94omqzHBiJT4o9wOmj+RUOP3Ugp1
CFaxZI+exLyWQaaLXgrUb0cVevmxEBQ38vV7mgIwWshtgDZYXirSiAwfgtjHn4BN
r1BluU0RaywTGnhQeh9xO9OmHsMUOUSKNVW3cSTvfZ61eCutrm4Yd6YYfRUMZKwn
dibqUJlx9jFc6dQh37+d8QlmRX9EU+C1ugvFVGfMrWrnIaw3QGAXPJ+z7DYuiPAk
CSrYvMFYmJufXmPXF4VD9TrUjr1K+QGEzLGo449WyhfhWCiZ44WdvzxABhSDAXOd
AEHc2r5cErLeFp7qoyrI/FwDe31wAHf6WziOnENDmgnEYsFxBh+o1Ok9WEGe2Vzx
8j9UKjMHKtbKJtvzGbP4A9umvOuhSNB4RP2MY5hpqajZsfRsKc1JS7HQNCcj7JyL
pVjnfw6IjtyrkMASxZvTx3hUtcXmAuOQT6TWDeo7dAIJI+II2twZT6/EwipSrx01
PePYKev5SMyaQvWM0x3tgBCiBOc7PLODrdkpX4ko0JYGkpETuuZ/Ic8Lf6ULNb/z
JL11BYdJgueVqiQF8kQDT+aKJDMCyCYpGzQyZnI8+ske1tYtL4Azgp26lN3BvN5z
w0z0/wZF3aDbX2mWdH4rb6EmLWyQk6ADc+x7EJsyrlGkWlQayjWHo6ibbqsxnC7G
igRk5+xZPVWPp5WKz0Wbx4NI0EfgVk0TPlmIKglLp2+9mHpUjWVvqV80h9417Q98
n9L/GtCAo2Mw2qRsBifmviZKMECfLM9rk8BQSnkB7f+sZXW17rFDFrWFh3JNsyv+
NkahjM8fayjaqQvMjdwBlLUnqquXCrIZIuySTcs/ekVWHIaPXRD4x6vQJqc4PpSZ
MUYOqDQGlniDNg5PQuqnDPS4DRyuNfqi3KaQj1cHfslYA3nERDbjPxrXPL0gdq5O
519erplv/HpUGqSHoiw3FQ4/urWmGWOHtvFN8Ub0PFVX7Ddd78XPfKBsES7B0HpT
fMGt+dAWligLX6SJpr78EV6uVSrCdmvlCW9g4RLc3lVJZ80Zys4wu3I//iQP2DNF
aqILbvnBYDy6KCLvAdnMqJ6+mHd3OB90nsJmy202wDn2pRScgmVMbtWA3wERuEM+
P3z5uLd2ufTVwCR1f0xUlFwMOOvt42CbAh0AqkR1NGyST0BKcL0klPlIoCLZl/hh
FJvAo+IDlWNGZc/adEd3SP8MYdvbIg8OPjPGEZ19uRRHyM3hwbQBoOxOIpHu7D+7
h6R5lvjfLvZClK7DOK6FLQmV+BD+3pfsiu91zzqLElTX3roabegppuT0ZBHes7Q1
yjnD6wiE5mi7XHS4uhjA9rtibFATH2DRDF5FuoRPIwF5ZrWw/UF/vmmomL9f5A+m
npAUZbAbKLC2Bu5A2BS76iONObbuvwW35MzFnnem0w3OsJ/NQRYreZ1aHYKNyCPQ
kTVTfzqmp2OUH0IOKXVlbqp27h0W1yN4vneejml/AbUiZaH1ALfMBETm6lLtZuTG
2nwbUYdhpSKcx4DslGM1vRFLK1IY6evp5Qh1B5+BSBZ5L9Ixifmha0InH7gt+En4
cimIIXc2gfqUOqKtlM5dWjLZqrASkIsKLgtY1SPP/Ex25Elu6MifL3QfbW8Yk8PC
sw0TSQvE1Uhy6p6q5Zfv+ArFzqd5F6fm1HXvkmvClRxtWXYuLeJj7Aa4CIhxUhN9
nu++z0983dx6xOg4xbEn4kj0dWPbSULqxSmYJ831PZr6cXxYJe/KiXVh/bukylcj
gmm1fqhqHI0nj6FkZ7Y9wjHhFlF4/XBawXW/+BDWjA7Uq2J34bI8+HFBC7iswz1W
9SMcXYFzycj84IFBxhA4oM7ltOqq05dgCR3NjdWtRFMdUJwxxYILUoq7ie7fjrnU
JIJrqGUoivcDDrp5YONPCbAe/vy7qXG4+x8L+x0Sq+25VGhyoq/AOT4vV7qwRDio
ZDTIOaZX/p/5JYzEFzmz6w2SRDW8OdMhlFCX62l+b1l+mjWcYAmOo7wZlQ+q+Mxe
rugEVARfJUTl6fP9bDMSRTwQGclXI4Mx2WGe3yOAjyJWeX37/JHBmyztIbB2m5G2
p92j41JmiArnDPceH2PDsZbzDD6VWEZMIBd7kA7m1AO1H39aPfpiMh+B0jKeticT
DpFcvvmdI0kT5dvvrA6KEMhFpj4ZN2vs/ASqA64TWU1pxX1NT/xvLt/LYKcELtZP
coFv03kHeCeIM+f5E3B3lDs+bnDSyy+clyOffJskClCo/q/RRblS0+da4w+Yh0qL
FzwB+roLOVdfxRVWSrRa4uWa93bny1fRkMD14OJpdd8HMAFBeAbKj6hBUbg9vjSl
ul21R87tVXCO3FjGo18xXndI5AJsCFFbT84tgep1/ERtWgHkOxJpM7Hy+g0k/zq0
dlKD2zDc/JIguWeCUTdqkObr7oURXit/aQVGqjTB2Tj4Cy3jcLtmT0UsTOKemrFC
pG29dra/9Iw/Ei/PSv/S5qephAl+L7J6z0eE/sIJcFo+N3VsBuJV7RTtr23L9Th8
p7LemZkPJWLQSgonfX9uC/+G9oL5uFBcsgQ+KRT6QOzpmiJr5+L0nQofYYl9QfW5
VGDxsGIxUOgwfqaxKnwXLFt6E2tXsyoU9Do8HRfLJPWHqQOF13miOioj90/OhS32
z80EAdgWpG5/2iFbdc0ZMpSwRQnL2lggjEE9kPwFFFefYHNDbTdmqQ5d4X9K2o7X
wIKiqHvnlqwK4G9f3Gt1E6BmTa2paIclwiRmRhfx3A8JJq1mf64r9CXSHgY3nZgz
X5GHKG3bv9bz3K9ODuwDivXPfLEAfpT1AP4ntfJmci7xb7j8S/cOz+6SIUyNpKBE
0S6OiJHpb2h6OF1FP27/pqXXcOYByw2BhW7JnE7SWb26AxFfGoC/QpGmAc/0YPOj
45h48xLXLxadd1Sdw/DKYIclRHt3c0W7NPmODBelxcfUAZVaiIEdMHMGDXe5pqjt
3LyZhlb+IdUbP7v2Nict5uWOeFApnt8KIz3CkxyffeX8S7TPgorOofDkwnsYWuUj
bjqZsiNLDkTfBzVvxV0TxrkRat5tRxvlX/x1YArxTx8W+/GS4wE63Y/4H9Aug4pI
/0nQwld8sUNQlrvM2X2HkdYB/RPqYWqLfJRthM8ZOwAFsfUuiQbCe37bWh7H8rnp
27pdsoMftszbzbtaKz+ROc2OK0RA5O86Cl+ZCf/aSoCD9o+g4dQuHeMF952j0gYk
lBvUJXiEjg90ALpHuEQV5TghfWmCmX8tIcLdD2BqitJSDfMlLpTnawcfnjH95Jcy
NCG2wpfnSP5Nd7dGwsaOe3DbZAGm7MJ/96tp+/yovNxRa5oV4LQO2l9yon+R0S4F
Mq+iUOXVrvkERHpGBONDJdxDexgL+0JbqxlUwEgIulA98X3sFV1N4f8CD2Mhw+oX
fVTCkZxRhjJXB9WsZVypgcsVi9xZ7YOtFgtz+GRKH4NZ6e/NjraJFPADw09fA2em
ZI2qLLHDlkG1LddKkVxNO31pQm7xfK56v/dvFJni3L/tRICMZjBN1iFwViR1TvX1
uwpNdI60WHiksYTw3HT0IZ4JPcLDxUa/UMYTJ5yKapWOtmN9RSPwUkVIslZbycql
mdXHVZLdjJPJ6ScSnnSDU/Ie3qh0YzsMzogshj65I5NmMFzAf6Pmlckpot+3rQeo
wgoTO72RDfnfw4b3SZV/kMivnlBX5zv42DD+5fG8/iG7HLGIK5CLxntRJx7kXHSX
KaasaQnAAqusXad4gqIdnlj724fgtTXbt/m24gOhHW1JyAtxMuJd0ur85C8+KSGI
ZsxR4aRNI/gdy+Q1eoZeOpjoh2UoXqDR8a16HTMsDwE/0fh1gjsAgN8J80m69BWA
2xZ7KkdajJl/yT/j6i4XoKf+XFhqo7zbgyypUuDrbbVocuFv2nVJ5vI+dU+ybBCo
S3gZIB/W3/qyrJhOue0dsCgybMvYRk3J07JtD+RCUveoKBpvaspBKtV5TFewUXDE
i6/P/lXtTkFn/gORY05wljjb8v4onH4H2SuiFomm6YuoUINAz8oG7QDxgK7c2pp6
X2wfczJ1WI4tm4vhBrHStLn/oGAs+dvs0aFAaUqgSpruU9VuSzky+6W8nSZpJfGk
9bwwjcv9JGXqUZyv5B0UnMZ1lMk7ragU32OoaXHJi7PDSfXZjYSCFPbJx7Ezo699
RF1YEGT67bvppqVnq+vD3I65tEhH2UqikN+eK3QaOwYT0A2n65Wn9zLVJvdQm93b
fZI7LyTKrkpBn2QXBe5lR09S9659egx2+pF9QMCYw7sW9rtdiKonRFjod5KVS37k
D3GDXgCgQstyHnOBaYxIcnM5+Y5Av997WRsRO8pG3hPbKmWRrS9kfnPN8WEFLt+l
kBYh44DZTiYLvTwx9fp3BL64f51wFsaRzlFSC4eoM4qrWdRfhKwym6iEjshWNPlO
2Zeo3QjwutRNB6CL5dVXyTFsXpvSKpbogkcT4OHQwak7Tk0lNjAg6sNSYiuWc9Vf
ZrdmhqpkiMnrK7XFHcufj/TSzNOvKHRCsTH09PeSyD0vTtg3ippPT7AP+TZdG0iA
Zt6rJMdYrmWb71OtswtnNMn2P9obipH9UMOFe6A24fb326sO2iVHdp2Y32JX7cqm
GS9OU7UslH5Dtt1ffQ+weQmz3rKRsPJyWDnhwnSyUyWxANoBJ7FaF9oXGQoJNPNR
0u+PthoHTX3ZkuNx5xSIHREHYVCit7pnp2agqTzhjWeLojM/4HdCpZ00cbdHGTsS
YFS6BUQ/WKX73HN5UnQyUT8oP34xneOxs8TuEL+fMO5r+iJuE0EEizQHOTUYRvYi
WKGhj5IsIndC/s5+CxAFwQgrpaVNWxh5/dRGIbFOka2jgtUpUI+oeiCQlb//73L5
Mp+NjRVBXSEWfeJfRm5G5iMHYGgXSEE/J/xSlvOzKo9M9heKRE9H/qjBYYy02iVG
eP+Eg5m6znHcWVnpge+lYvvyC2qRPIAFSL6GyBVOIMs93Od2gRpe3lozVmd9llTg
eWbZpU7hHxs9Rl5968Q711Gy6/5ekdLxk5XZfqXfzq/2avPp7g00XAVi2qmvWRJG
eoBqDsFgFNa4PxmMutXtYUoQY1O6wS6MFLshIr4I9IyBxc7AGKuTIs3TgdO7hOlq
2KB5xEwe8oJgDo2YOrdeVwdWbag6zlS+YponkRVIcHlEA0S/EPtRjmhVYQhGjBUE
8kP7OlROAJMr73Vmjl65YnKI1GgluEsuzDwLbbjkGJ8y1mekv+fb34f9uMuN+qyR
hrii0TCM12DGsWDkizWp33Lh1cTdtjYYJ7PDOvQ8egzUHD5ZrIkE74zqc05zPzSo
IqAFy4WT2AA8XUmBKEy2PW67Z2uvdNGQttm7MeHR8SSTG6+L6PH65TSWKjr7smIe
6+HpWsbJRko7CeCIQSN0yDayJxl5baggy0pS+Ebo8R32uvmAjuxb2RYFu/Zoy0Au
eVB1CO4Vj+ClvlWfCmddEmY9NQ8Ul/O+YTt3vJsR0bngsDwoeGFTKIwrIR+ODlCc
vn938swMbE3ET16b7tp4iyLUwp3Sr2ZT/ENJ8+TfQAMf3QG/nRKjFxLrQm46LQQR
OYYjhXIkK+TPSNX/ruiuPlvL7S8jwDwIJchcYVSnEoU8HsUDsVCzKy7LykjEW/og
7i1PZZ7CLyuQIvEGn9a8Bj3ndxXWcOcGJ+JtwZjs9bSHIlqJCUudmMAvRk+4z060
FSa3RraBN1PaZiyYKkpaPq/hoxIHDwdC47/CkZ5OwRpJeehQjoSfVulmgBxKV9sg
pOHUHadOp6dwa945B+GlVx+7Z9Ie6L5r2gacROrT7Ip6dw9k3fkU85bBObvMsMhb
TAdqUKbkdRT3eeV21hmzyg812X3viMAuFuYR8sPAfJ0SZeLQvrGKfFqgOOfLsMcQ
/uvhMfDcf9jN4jvVnkz37qGDc5MJUEAmDwOBMt0IXB+XPDr9HLJQgPsCxTEX7Plr
hu1D3MBufAqXJLCU5R3R8ufPkcFJ7c73hZVV3d/anVoGsWqpHuySgRyuHyptFXDG
Z41z0Dwo5ekKadkbQA+wp5WVWL5Lz8LryD95KxfgTzLXjZP7lg6CMkAQGuvv3kIE
2WLmAyTkC+LojMc4NDoW7cotiLfL3JehHDK+FBXkEYtxBOmMvSV88kMV5I/0emWt
OF663moZTFma14hgnarUqyeWsp+jDP1ikmt6X5rDWFL1eWy8GWi4BCiK4BYvV0jW
VTjZztk3LDIEg0J+TRkewG496P7hcNqB3IG4RjiwKmF8U4PXqViTYWXE4UDd1fqJ
Is+2nzUV090XSgxVhcsGPavnmxjMQ1CLORp+PGp2Ubpe+vB91ckcwASnE99w3o6j
JSQWwN4GmBOWiP/MwuuaeIcWSG8NZqUIp2vjR3wx9FUyJouSIiwXRy8T3EgRBbGx
f0WC1OJwpxuCdjkPb5R8uclHfa5yxi//2n1CJi79gw5lbB0/yUwiBj7DGiuVqGHL
JFvPnVKA2wYP6Svr1w6CHyUqKc8yBnyZXwh0aB2ZLZ/sd9zxvQmw5yZpyKOGp242
U/0M0raVtfY7ky5hFYM6bKEd0mxonmsewWEKcfUDgby12tj1Cth3tWc+XnizD5Cv
+q8M/EE7ybT/XB4uZ3RMJ2V0jpuI8Q4cKFyCSQwZXmYbPTezkuEs6R9t3OGfXQpJ
O19X3hbEVTYoOhvveWUeMEsTf233+tsd0RdmuDjCpjVHzhTfq+Y7X1QveF8/suPB
3WWLusWKmEEtaQVoi57r+Xw/5PHnfoTtHxbMYjzwOsFFqzPqQOfTblAvHtpMJRPW
lcXTKxwT2JxenRZ2nXDGMDOEbVUYZr79CJHfn7zwSk1AqNCFUdukAQmCJFkWq+Ns
2lnw2/WwuXA+gid7lnyWfOn4ICMrdW0gJR2Ct0lXXPIwz4r9ZvluwJOHZ49T9pfZ
c+m6PlaXIx0MCCtPN2ZUyww5VX8XUKniXc0i7OINDLI+rgj3EHG9ouL3zMCjvTbt
AYqresZUwyUjnYw/wRt6gTRrlCDv910eQmX9bINdzabEtVbIW4k4SEuLBEFHLrXK
J26LJN0IX8pRO86hBxsfFJzefVHhEjj+qqJicC761UStx9PAbId6i2QzUpumdZw9
9vwIsnnQKJ4suAJV0t/LjX3IRdeUrLXWZgPqkKkrMaMbSn2/TRK+QjAk1us2qIzs
41GDiYzNu28fNjIVJv9w7q7UP/I0E6rCITaV62kQbK1LwjeTn4iV1wikQ3gYyhEZ
8e0TEfd0Jw3ihgUv06FyasFwDioF9OpT4IqP88NN8uTIj1XBzhhU0tMCHewtIx+w
qVW7Ke4EkE6/qMB+JmEkR3vb5WT36ZnZz8ssj2baby1tN/3pO7d5IHYJDTRCD0iv
o+CE/uH01SICyNWtWEf06Tjm0oFMnLEaWHLlKSeQlhKHSu/ZKA1P1Qx8US63aMM5
cQfV9Mkuu8YWt7bL1ap5ZKYBDxdvGSpvf2des/F061N5/F5z+MfQgI7wZh1TL/BN
6eWYbaHtDMNWQ+gfIQVppJQoMfUCPNEGCOaj87lQeYs2/JX5xUL8rXJVaorplAwZ
Ti3IRISl9agVM2/748Ps4uifS8r9zBPUgpxmIcY31vEu5vH8bzi1dRC3fAh9v4gS
Amo1EV+gJY5+ZPfX5vohELw1ZaWbsSG/nDuDaNLwIzvhwG5sKpykky++k+Bv3DPY
IdZKqqvmDWPA1LZlQtqTGVGJ9kOaGAp7HYzLnzGx/ZFsn+jMr6S24YZ4FFePctLY
hV22L6arcatoPXBIhFEKEh3HN3uEwYOi9ry5MzM1UJEYzy4RTW49b2HhDRz2Scyh
/4KoguRdm7WXT658OEojTSNhR/VS4OJWv4U6gYBKJ0BRj/AXJGUqrsD3LjS2iXDb
QAX+MXTE7o5ODrJAm3X9t+/e4K+RhOMRG1ALjRKO/cfJT9VmImyo/RnB9UpZ2aSq
KJX4Vn9fu2sCEm5eHbxlrrooT8mDfLokS1xvxBHieFDYwcnWNmN4qs7x3Fco/DxL
Wf3kh7f5MYiXq5KYBoCyvF4hKjDU14CzGNZYBN3GsIQ7ZSmY8j/JiIcDHLwGntmB
Ofr1BM8q6xjHEZxKx3sRmOi1LFPsZ+09KQkkLoIIyJ8PE3zLWgL+QGzaTFIByqmF
JxH5Ax4h4PBQnMjD0BTSTftT0dqkZZvZLSzrGS0yy13U/O21FKrNvD6swp/IT5Uc
fYo8iM6VLIJdHYoOi8JD42SFmU+Gu2/8M+4wzdbnA51ouKgYy7lh8AkfqIk5WXSH
sh/9AkeDtWF23ITmh8/wj7n0aW6FZ/7B2JnotgDAVGqGeJzBGwiXMr9Mk1s4sQlG
OqAZSmQ+YqWWUvFlqRacBjZHmJFRIbkqy+9jyRdIRjSt488L/Di/vIk5t17Zi25j
Ccauc3p6QRydbEI9AkFJYh2e+TRkP+C1KZMm2FpvD+csM2WVMkADP95NYjsXZT5t
mNYm9SHhwna3OQdprO9/yDj4oMlAXZYKtGSFTFomaRfO6xGQsdUIjQf7bewGEYlk
2Lw2q2q/0s8ChySOHfrPK2vGJnN5g/gfVeEiFgkaMXOCjXzJj7cLBGCAM74pw2Wk
zQ84b6mEDNgXuouh1Gtc/v70/Ti9LrxsSEdRLmcK5mdmlTEFaPUTlu6j3t2vlkiC
G8ag+6/q8ZuubWfRZyxkMYbupCPW60+ZzZCXS8BHQII13lwRInDUS+e9JSVrcKr7
noFT3I8qU3iuPZaYq+ONUl/p6DOIM3cVo2n/FTjz2+748KY0GlrYn7JPBwRJT8YX
Wv+Yfh9qt8E3UnHKpmbqzScAdulVq4LWBMHfo8kmjBXUifm0surwV1X6Zf/X5og7
+/LPn3SbtuyMsG9Ttd+I7kql6NzrK3O1VMotX7S4huN4/JidU0kL85zfQ/7497om
G2vYKLBSUOSnreUYPZgt19IqxtTf7X60h7/fwxo3M6Ov0/Js/kh1ePd8iPotKLp6
zQDtu8NvQQqiaenAv6/fIDEx/rXZmmiB/eeumPZsCOROOW+Fz9acA9yrfJM0Q8Oa
oEiOqOF6uVG72p7AW8w+PdTOPqacN4mBt0u4AJSmMiWWSkNvm3KVuSqRjlcfzAqG
3hPv/IGugZepynMkkMa2vnV5CfalKgcR4U99264TOzsappZdUlo4EAAYWFaoKKN7
CD23IS925iicf0DbOfpJN+Lm7/BQoVkCHDO17UvRwBkXTGXkmRoA2LYujKfiSuRE
IYIGvPfGIsRX93a3iTaq4g/q9iePXs/fxcbJGBLJfk2cebxX/D1Eu+pB3HWSfteo
ACdJpsN1/4tPIAzm4wWwF2Y1VQh9CeXy+0idnHbxRrfMnwhT40oJnEcF0a06O8g8
hlhT+2RJQt3HZTBk/AMZ2o09oUJR/M4ERB0GaxezPsZ64kBdyGGbzzwKQe/334sM
9ZljFWAVLDmTUIAVd6FT+XQK07GrlZavwdPj2TGJx5ImuOf2TyV0PUvx4tQPWSa1
hhsXiu14m8eAj4Iw6Bq/Rh+rc7OBKjCtH7XzAkhrvYY0kAI7uIfR/lQAiyYBTJBk
5Gh4Q6UJTKY58C6JvbRmgy5SBMJ1xoUOUGfuKFO8EDcdTwXGsmFhi/uTHLSKV9UH
CusqXIPmp7jQvvW3GoqB1wLorIN2g9OeD3wLgefzhV9hPRI3Qb+9IcllUEyYGQnR
oO1rjQSOfGJYLag43vLFEeH2OTu9QIdtoymNbzTI3U9TnYPLj7jX5RZ0OUoAiFNT
e4JzdGaCkzsCeoX53LBwX00mVsW6LaV9JZ3XMPWC+0bcGmOr04u2n5C/wCiCP/Rz
cYoP4qqqfv3n3rQS9aopfn6/9qauyulzJUhuovcoUwSEFWwYHT9dbF5WtDVgSzAn
EqmRJVQO1BYIZqCEIR6KHli7AV/R9dXbGB0DO3CgpDLXBfx9ARVh1BSeMZEQ67V3
EOv0LPLSXB1HvmFvggF3Ua5s0NOah7dBECdjoa/esw5KIxvrI2WC8RDTEYycUREq
zkOR36gh6HXne34H8CT5Xx+B8ID88N1XG59d/XEGXJ/e+ZeV+8QZm6Lct3AduWE8
O/5GDr32q9dByQW40kPhlKctAgECcHLLeGe5qTPGHrzYdRFmrH0NHFaZe0wcYg8B
ODtgvqQFcOKeygTRi9PLjGNrmDcdMx/FwkkaVtPB81JK1dyJMokqYLKBXaTdl3Yp
IuvpNeja2IpTp2JkbRFlqiKLzmCElajVZd5bdgHR3kFJfmWiheS5ClTtv3g4VEUI
3paBeK7zDpOOWQCMVvVGq+r3lBG7Oujl8cUNXbYC/SEcFb16GbGi8VG+bDbDqgRW
ZmRwUhvXmM87mEvu4s2S3EqQOatTM2p6cuxurxBviIg8rXqd3yoGW3USPk7UYSNx
rcHyoQaP7XufP7nr/3ht7J4qp2fXtLDrXfpDaJIB3GuJ0zKWpZc/duZ8woDtBht1
C4Lrjonf3/6qb67rUx1/GYv3zuHaf5S/pzstDBuK1es6SBNj2jc+ws5cMJJWlerk
5ciyNpk4bskLYvyd4IA8oAERJWQEEQFa0pzCVoR3CMAP8nbivw9A01kyTSbXtDIr
b6W0KTEpJ6cCK1k1K/aheZc4PTwOP/Rv2dAbrkOP/pTtX7OupIUVNrMwTPeMk3KB
biFlhDDhDI8ljYoKNVoAbXRV1i4UruUiN61jqS0fHHi4JsBwGiyCvr4jbE1ZQ6io
uZv1ziX0HR0fOj44me1waqyHaNb1uqxdl2Kxbc/CqPcv6z44ORJ8BWnunUCDA3mV
Zz6rWK3K41lE7jmF2aVv5aAKp+Z9UdKJAsFolyjDzJA3G0r9rKLiaQdjWnuwWG5P
D3984VFXMUArZ7CG1cKWBYyfiWLbxBk0Jwy3wzFcD/ck4J2tKb3hLvAWByUyyY95
DtUWZoJYvq2qWhN6eceV04c4Y0nv5u5neaYHGL9QPdRJa8y4I58jXqfCSF5Fn5rH
oAx9AtQTWDDc2RwQDl1pgDi/iyyagtq7nS5RhPFR9Qtb9f4o5nUwKWgu9HzRL0bX
7xl4ix0FzUmYNFs0XDan5HY/hOWNeUZ2sAsxlMSaeA9Px23hgJ/JHuWnlAGbribB
UHZUPmkUqNxmFrUyktqNHJU9iHFAlloeseWHtidcEJ9qXPPGRcyBX3SWhgP4q+ew
bNjdrtEr5S9wl5MLtoAsRvBQPlhpNx3u9tyXJxhHCDqZlNarLUqsHcmqovDKzEbN
KsDclVvGK0Eh5z8avEY5EIcubs9BFw5usy3tpioHsnmgNMp4u6HlUNBkoYsV14Vu
KJqJGdcaXwaGD0vz+u3V9/r1W2oWFHIYY9dpYzpHE83vvevr21LgDYRkABDx2fFT
JpgBjMIY/gjUxSQHL9bz3zDJvxLB5apP0+0iQlkzjBLasogf0lYiVEfZX3qVryYI
bjRHFyrGFMS3pBhGht23PJTqhtlJasOThNl/hl3bcTcbemicBUQxDplkcIh5S7ks
bApyX1DXukI/h/3xQ2xRYWqUyrVLnNVbj414WGY3NqZOAbayV0GJg3OrZuMP4g6C
D2ZkQ29lDtLrHURTmfbk1CxJ50hxvvhzcyHVZrLEeSKkNsgcAw5lH4NmunCiuMOY
FRMeENksJUapOqsLITk6xJ8mCHdI3sOr/4d5vzfDxaqcgKwPo1PUdi4ca6Xuh1fT
1VImhQrjlY5WtfBm9aNCFRoq1Q3iuxq72vnrEM2mhYRljDka5MmdR/VrAg9Lb9Jx
glgufvlDguffQv6T6IErZAoWvh3E/amS7eU2NoDYZ3UiK9ObiVhpW11Nhd8Ec6HZ
HrM8fVgvJdPoh+lRZLwf5kRhalxGF2Ga97oZW/+Hstm6+1dHuoJXC2QVeRwV+eZL
Jo2SQpIe7an6hdx/6kKoOhRmRL/Sr7WIS5rrTjllMuQ2JYV2nmd5gP3NJjDXLXa+
72nsul2pJwrploK+hgCi071NrpwB84KbehqiGEUYJa/+UXctFHtcRd8cwLh2iE38
dBTk6iLdCiJnlB8/aZbp3uEWMkeWh4USCS6g7knaC4pD2JVaCtlfdZLLKyoYbSf7
ZExE9XWj4u474kTtvfbV4d8bGTxqQ7FYitYehh3AjaS/fVZ17hDOqYV5Gt9PHhcR
fb2XN6OU+tAjfzxYNx75NLVObkbklKaeaK7gGn2yyM69B5PijkA9uqfZyiLZbaRe
Mk047EzrHNKXkyzV9cEm850rzFoiQbgLmLHYOOi2ACD+EdAjWG6KITatwI4EiySX
xdL4dPYItiGSFuwdQ1fsLnhVGuCcB6I48GJe+k0DH4ITogPI5izG1L9gP3JWsNiX
lNFAhQDmGcnn7Oc+mlwTXnsrsl/u6j5fNahgGr98rHFzWKLwnEJ72lWRzUpuvf2/
APnkLA2lWNc6m+pb9hswH2+yxWkOPHxTnrC8SDeLx7lhUpsk5uQOyM5A9JK9tk0W
5fu/Ng8KQz3Hi+ipC2dNN1jIxlAXyVOp3h3i/9pdb9vob4+TW7/D6iuLI/WkRWSW
lS2Bzk5k5g9TfnCbgR1SB/prGsVhyrCnp3RT5SmtaHH5y+iRVCTba6DWNixD0yba
otAWAAi0NbiVWDHoriPkahbB1AHgoHqU03mHmqHg9BHxJ3lqChwFpsLBILrrxDkN
rK14LiyhvhoSzmfInukDl88KSsEYokDXqhX0zbJLaLSZyX4KJ0iABXYCWIuguYJD
8pDPSk03YL3OiBE0N+JJmg+QyMYguttZzCpxojz8KgGq3VdAH7F9dYc33LqSS89T
ollBlIkyOIhEqVSZDufAtXJocjsuL3tIr4HeNlCvPRiGD0SKP3AmN39x8vmk//WY
yxi6NOVaID/NARd8iidnfterZb3PJfitEUeA0VaNflhE7NFvD/230BAC87u0Fo3D
1Y+iAfzcWTS4Sexo3rm/PRgIX8phwVohn2i1p8hFl0rpExhGg8csNjSUjQYNvPyT
X7Gbsf9yKjLlD3fUirCMtCkaPHYxrF9rE0dNlh1tO0O8h7UYdfbIJvQXOriOpWz8
ojvFPdR9+k+LuPYALzW7NqnS/A4Os7zMGqrsvAPKSYUt36kAOotVvRxU/pHueDQV
Gh1bxxY3S6bQQ6GoPgR2y3hQiJWHfhzztDzNMLwBa34VIedNEZeP6Qg2d5yRpvlP
6+i6tb3L4c47VoIuRAB804PASI7wFa/ztTe/QDeP6B/p3R8TSNm7t9X6A9bImV4N
IBL+Cev3nWj9wlwIiB7t8a8mblO5ZQatkdBG1FQzXTVGPKp+NncXmbgASeaSa3j2
rVOeP6DyQmu8RJP8JUnOIs5ZMSdN8+X0agrEOv64dmZ67Sq2omdOeWsxgLSiE8pu
8+fTcNLNxUt4x7/0MsvLbVneVI4XRALxICSOzJNzCaFDl66BseQWkmpN+8vbbhv8
2Q9aJm8O/MZtKVWZlU5DiXzhL3LLZDMiJ76QYVxF3NXor/YmVNigkUGezwYTCrqE
103Lhq6K9lvqY/cScdwPhZTEbMhRV9R7I2LrXa223QMSGUfroqCnUg0/cZYS88Dl
rWHKyHEEcFtkoY+ZKGSawTgqeM4fF+keS1ilnfQpcdsyUw703zTWDxpEWh10rnQR
5jUwjQ4PORkfCkbjoDUifdnn1kcV2crVamKNqGJn+l5AjtuVmu/j6Zo/ofew24sb
RlpRzHVyhwRPgK+ik4kneiPvSZ7VdYGLkDiBmkFuEW8j28rbOCvuyL2nACpAUKBA
n5weniNY+TBEKyLR5qLoMqITZByHfXfcIp1JPxhAAqhY1Y9PNR54khQ+ACHTKx7J
VeUOJ965XqXA2J91qz9EliRad2BiEfFmxVrPiC6aLSVvVoJLb8BS7GayjjUodyOB
Z1IIsGdQgp9NE3XbJ98Wrl2slQtXXicARAAHfvDlwDTHt6saRDL3U+3w2O3nekUL
bprzS/AgSD3gRAh0iX/ysSuR7om6yNgGYDslXHq/S/wdBPhpB2EPiYW9f/1LoFpH
ITs+Lxgay3ouHYjAOcToRiYKC2+v46vn5D3falzFFL77AkPjlC1Dg6nPb0V9GQcx
1otKlsV1aYGVo0PgHbs4J2wAaWih75EWHbF/n1AJdGdGeqwyHzOEkA7dleJA5O+p
4FTIkhC7gFgCGartbHgA+xwqgMG9adqoVo7oWMrPHGNKohqRZPJIl2SrfC0sZO+6
C4XcIfrRSJNoCHP/4jTT+UCYdkP865rrEJHFCpaPXSQ3wvPnze5cdWwSzaBM7Cd2
e8AGcNvXlRrFnDIQRww8iePNEjIgVfel9y7hnjpn/FxI3dUR8GWdYFKZBJhjk6wo
VRthcNznHdeEBvUTPjxqvy+JGqB+7rSRE34mLJCGmYb+yX1OGxbgGUT9lo0Nc36v
Y/fYM4yuAZnY/2dpbVGm0Fvow7xv81tsxXBlu57HRCx86q3IElkR5DxYG1/zRIyy
BKgnI27Iu9udljWDDv/ICUfpzjple8BM6UZyjZnE4lkVt2mv8szHf9n/7BL8XI4G
xAxjS1DjpSN9QSPNHc4kECiagD1DSlddKx6LyOzYhmMlaIlVhmcw+LJAUxkdFDsC
5UYSpZr5SluD/mOvHDSEYBKms3cSM6JfRED7B2XZfJPqN5Ez2et0KqR6eJlYS6Tv
9ED8mLtFbQYGbBbd8UndmgUTvDVMjEcNmJXkKFluFJL3AqISNcT0XEza0khP6YBQ
xcmmpRPM0vnWEIPT5MVUgUCVUhKwBCgmH3IG9YY4mnUZ5oYQzXC6m8XW7S5UBgvw
3YvRoZvemOiEzb6/8NlLNSKlL7uBal1Q4WpclgyByFx1yBpb+zYldLeeMXpwoQum
7TAZp91SrJjBZNLiqZdVFLzlEjkG0U/t51EhT1NFwXUk9ub55OD3cKtUgsm1VW00
UUBzTWE/PtKVK+ZZSUwYs0XgGYueVAyVVQdrgzM8aqG8LuHkQcu2vwD7Wh9izSYh
+uRrbAB/lZOeN6i9iLY76uTKw9vsK5ylBVjHk5HPlEi9jKnn9qrQnfQZk0lCS/H3
nSqVzkXjV1HgADHN1KKG4vRITIRocwHbM6Q8D5CKb3TvLI8SEGv4n71tc6SlB5il
nDAgtQOyrw7Sl54Qae9GOM0DfiLaCorlCJkeR/hqQa7dif4LH37Jwthrp8ekJUYw
q3szHXh4qdQaoZGnHJjF+mAXV8LVDg4LYOL32TLAHziMV5da20g4wMpoJ+HZJsPd
hUa1FXQlrZ5ntQoNG0NZnqGzsQnHPNRtFx1K7Kqhx1kboYHlwchrJ58F10fnmnFb
TR9zceQligKKnnANVGgthI7bz/WyKq6NYDV2sToXLZV8mgkIGeIP8cI+mgGs37XV
PNIV4H22xXOAR/+uIRj63dHILPttSDJN4AcjPAGpgVhYxPp1F/q+MTCCQBpFJO00
8f91hJ7qtH4l2xDfoIbt4bVsJZtklp9o6L4SI8Jl+aWu1nLt0tYz3wOSlEeB/IQd
7xwJ/V0oDwKfyK514GwdmadtPQlnKMMrTkS90hf4xgPqRY8Xj20CRyq0uZrtzRwC
kr5HEip78uuXIgXog9bbKKkKngAZSoV5jsKuSzfC3bK52a8B+LH++5/34uoBdujV
d1B1FmRBUMj3yJirO8EMVYxadFNY8MbtZaJxN1R9UAB4twfegyhCLcfEucAYo57R
9wal4x3o+4D/7sBUeA6bV+bUPP5ewrrogCQUlQG8B09nnjC+nhczrR6oW2HuyV0g
qBn/y8JGFZfus5mEh8Sp2vv6IFyWd5jBYV2U24qRHj9kE3UqeJLuBezd/cl2uIRB
t1IdaDFU4WjcU8p4hqF6TSC+p8WP0WGON1EpPvw7qxK/7qqw31CYFU2BxTR/jJyB
16vBZI25VukX9qygpSVFRveSpqgQFa/TyC519mqwe1fMKzBWRqZYXnzF1EJzJGYK
DD/wpvcaS0Jmo4as2NFA37EwtXOZHvGIvJ9i8AYEvNyFgqS4MzyNkJ1YDR0iV0v9
K+pNcrhI9966xmace5lJVc0Qi5X8UGsr/Gs5sxSZNCiN3dKUwEJBB9ARRKj+Ve1B
hEn/asYPABKE/+tQKYaotbWUXjScme3+DdUid7tkmRSc6ExnCpE9DqZ2wXMjVGXU
OZi8CIp2r8x9DfWr2fY+T0R9nW3XaBRIA1znwz2/fkvAbnjtl0+sYHgCcth/MN0b
5SOeNe4BDGMQPETLaXPv/Cp/0FR6GRQbDy/Btrx9bXYgPebgUFSmPB+DTOxxDDl7
v484vq1gyxXnpcsveDNtovvpWEogKkslaashcam4ijiv2xLvUeZ83hctPlcY/0cB
xYRNSS+uapgJPY3bf+uFaPOmmolbp/Q8iY+va97NwXnv/C29+X9I8VN/NEVnlD1i
xmD0VrFU51EYNekj1IeDViCqT7j3TalITlk0yJ70PcAmYuTn8N66AHMxhnR7vse/
Vijf9L8kRP3Z3HjcGZQRZhmzE++5Mf4VBrIo6aAKU5LA3mmSba5jsg2A5ObjAivk
aJIWN6UilNT4MY+l+Wj1xa2DznVWiy9LaqABlcFc70mpKkVEvDIJnHIypLhYN8UW
PQQ6nKA+SuLueQrz3rZZUN/yZXxVhrSULR0YO87/nnAOan0nrwfAEHWX9Non8BK9
2uDZJMc3zRKd2hV51RO/UJnu6AzNeIEyh/goVUJvCXDA6X7qkmYtVnUkOiNw9sj0
vdRLGCxVy143XCFDswG9yvvI+4csIIXpLeA50uReTVbq82ocPSyslGEHpOBkKr2A
ehrKlsUwGIXfFlP/tHh0jRIZE9BDYdCVzdBA+oCaNfnflZoC5wY8H2w/O4UtJwLu
+eRPp7Uff44Cto08fxzswXYy8rA4bfkaP54dWU8xpqKYp+dA8pt05IMV5L1jKt0Q
0GtVsRfV68kza2jaWMPl1pMj3tbuIlJhfLAgT6iXvqLTdG9M3lcGdoKYWK+5Dmae
IdVG/zqWvRf+Mr0SqJtBu9cqJRMOTdW4AfK/8RBCRNOv3umhyj4TIbFf/b51P4Gg
YJI0c+WaDwfb1XOjZMu5EVJib1L292PlU0pRrC/3AMCCzOX1mY+DsqXHSp6n26CY
iobARPHJX54R5bVNVJA+kpMDewRY6uZRlH6qtBHcodNrY8FuesKDEa1gou3nuBJP
ZDGfAPT1NR6G4u2vGJaE0Sw2TaRxm1LNfPSHRH7ep9Piwjonb200o3Mc5YT/w0S4
8peVbVuq3T59Bq8omPbN1H49NWrwIl09tqEt9SquqkoIzIsW1F4TJ2t7hwAEEW0S
OB//H57SnfauNAwDDaeYRVh/gaZ9OEoTGZcGcJxwvMZmrVkCyhRFzE5VYmmlAWd+
EhTLkmubEi+QGEuKI6KJx1wYQBrP/kmW5KSKhAdfo0ZXxsUQSffSOIyeraTUjTUD
DaYdEX9SDPiaIiyP5WbRDfnCCSrfK9qclCY43ZInlopmNaY0rVsyPqfefNtM9wM8
KbKMgu9jZUrUodU09RfWs/McA5rrJIA8j22RBI89guz5/Mf47x4Y7akMvTeC7FrL
SfbrrDHczDcykv5fhkxGggdg9UrXdu1luwzoZphE6651VucqHldGyaZRTV2pH9Vg
hLAV3P+Ldcp8HxIJiPWpDLxSJ+CA5fH4Sp0/ufR+QWD1YAF+2PLH/LuBOwPjlv1D
Eb0UGVRmOXKaUyBEIOoKrZgzD44aCJt6jS605wB6zvDNkD1TrBpMIw6d/FJvNkLc
94xtThQYKTr8V/CzisiZTjcDjZ+tTyWFhu+rbvPv4ydG8DH/jukVxcJo4UiVKOxL
2a+GeK2V/cD+Qz2PA3YkwtIEtFYmWxPcLUUgrIDl0uUiK4v/FgyAjmgD9rL5aXA0
4iXCdAIb/DuAo7edod87+uOMav+jddtuTvqNYhkEISrdLPUyb8ODSt3ZJEzq3L2G
rFnFQyhHYvLIKITF68rBRceA0zKQTfCt1kv7TMZ3YFZPy9R5WLUxPIGvW8vEo0NR
HvZ54SkfppOptEJ41lUXgsMNORITR3SRs8lA3G5OuA3D0h9E8lu1C+TIyXI9GUjN
3qkYBf/gLrQ3K9QnBs5ejXaxcOTGsBSDyJs0vwshiIYl86ItTwYQPqisZl2tJkzg
dAcvVO9GPMYLclmat3mwdj3zGPecWuS3BfOU7y9c+hWgGGBdwePEur+75R0g6Oz9
JG/3JncZi81nbCY9FcE9jEZrg1cS7F1damkRNCJoqcDxCJXoUl2gJJRMqO2du1Nu
J8XExYFuDpYKn/V5sgFD1PHZ+cH86RP4YWK2Ua4IJsM6Oz6bH37aXif7bJ2Px14f
kvUs4mS/f7/8yiLCweEpqIz8KAiERZADCXUHJY4fN6dbDMMq1P3hVirEuxj4glvG
ZBklJd1iUfscXNYvb6UtrFqp3hssvc14mUXw6OMt5qzrsuS8yMKhU3YOpRM8Qu8H
q21thEhi0uU0g61nVLxU9kuIJkfwp/1gTaO6pHK015xv2Ws04kOP6pt7woFZt4rj
PvJotWIK1HFupWpGsaLZYDSkOJCsdhesGV116I8fiG5gC9zEcUZ8oQcEd8ZMYNl3
DujS3Q25jfAD1XF2z9E+dkTXAnf/zPieEzaFt8TpY+YWAn2r0RdqULip/na4X4vT
HL1Zb1ErITMGaaCKJjvsgG2q2lpcn3+hcrx539R8oe6tYQTU453z1yZ2zEI0fKJS
BV/va8a2yTfRGbJK/kOuvGFeE76TdPfvCO09sG2vSz1pfV0FR54E8q8gR5JgwKVu
7szmS/YEn6vNjSTY8OLJ5Lgw4Lkpz4mxSHaQRdFhhKcLM64ifdudzRMFuy/tQ0h1
WdelcII6UCj3ic8acnO0gn9K0/wdQ6sjgjMO6j3Daf138bE3oUxyaiKPAB75XhzF
UM1oZutpkq9aHFnLf4f9OeChxfISDiYImnMdkIoFpWzLsE6ncB1+xZg0WsX7iX8f
enKrPXAlMXEm1eLmaBbSVsge3vqnoWRzqYSLofhNQ/mXBfJJdN7jItOP0VWGgcya
caapSh6T8vu7VWHLmg1ybbKoITai6h8XpZUKH2mVREAtOfLddqtnrkoAfM+FtcoY
TFEgvIqhlvK+ud22FG2sksw+UCGCohj20rxXN71vKkzwSeeR9gv0/09rwrsh7Dh2
RELkUkeqCXJ2qme8ndgCLNR6iuegGtPjekoow9R0nOOGTg6+ocbmFVsPqWnuy37N
z9GKfGNokk6MQAzZ/+zAKgAW3tidXq2PCTIijHRzIgoSRwXQHDQv9wpRUlh/4xGX
gTXnqJjuHDXRMbhBsEkAeHECnRuIn1FVpni1moBok3OjOa+KoSwYMf3gGQ/fnKX6
9Wq1MEitHflsbS2kJe4N40lphUquiTNM8jgoHKXhHTsxjlBUhIbCnJTP1Bmh1PmD
2M92dTd1pTUbpTGVenusLDuHdSf8IW2Qg/gxdkbdKeWt5Gt9ojJqCh+LYb06UiwS
h31IfFjeU91OrA8wGDy14SAcrwKhrV2EiUcf6S7HzJ5EU/TYbRzWge7GZqu2jvUZ
9zC49jAcZikHZsRM0miRxZIP0yBlY5EKSdbMrJyzsCX6MICVYPuDUYs92SImxPki
jc+LLGUfxN7/3moRDO+2FUj1r12Xg05u06hgUTBYro8yhqhn7wQRDbnX75SeL5Ff
Uba6OinwdUjJJoYAFbxJ05dOCih/4lJ8X72MyLr+/3SmnT1WjjNCw6MO+7WUOBn4
m5q6hhLQVk/1aKxMPAHP+++b74vP6HmS96ogwAs+Cg8kpLP4xNPP1dvwuClmFnxY
Cb0icU/4R2EdGvGb3Wdr/Y63yk6fai3AVIBDs6UQDX70bGluWAECbGcUv26mu9cx
lhQRybOpdgdalOYXu5qeF/oWTvprvggoFZFtTsaoZua1lS5+fNFc7efohnlosqCp
HcbyH2FUW+tdQE/xQM0wBRVe3ThHrbhWCZj5BQoTcic4MEpNKLXgh49FIz1Ow2w8
J+pUx3IzV9zJZ/S8zQBJUxVfyhf7EmtHcUa/y9nvjVFpCYpzPjtbJQBkyjDLc0Z5
3G1Yr1Au1kynIbQk20w2i/ukLgPe/5SB9m/XrYhldg9c8hzLUPD11bnnf1+q718m
JrPdabc+vyxMcXL0WxCJ1dja6QV6CAnf1gBDYA6iUr3A6jJTnpWhLrZzTPoQyF0Y
RmsKqsYosNx0+IdzdAOFqXt9M/zqr9Upp8GcxnYpiYWj0i8QbxXh1v+h/laUyY0X
iGKEkqLt3ggzolscL4KlIPchonphhXt9XHYGSP/m5a5u5/3h9Ck1gpdSWadj6iCL
VF31330ZUXyDkbbOHR2v229xikdQUmjFC33KmuQ0Fi0S6ll6v5AbsnvEqwUj7mS/
7W6DMtWUmHBRE/qD8kqVyMavNCD8Y+SUaPuSIevb187Dv/HS2TIBxHsegN1/5bEg
rZWGUe631r+58NFyCg3l9Bu1TrbkCIFy3bpj9rflFNcf3UGc2uYAYnVQcbNXCVl1
ebVbt97su/zrqATs1+Mt0lAueOMG1J7CDncbCJ0dkHYyL4YlQtEx6QwmGRwfE9hF
2H4ZJ6PjKKtppzMyFla4skxnqtBDk4uOtbG0gS72++dPUM5tLkLcHB5JBQp2cIQY
X3OUtu6ECKSAFqkZCjppW7YeBiZNOwcbMmEAWB3xRRwRezZvmPg+LZ3t5MHB+Bw4
Y4MpF1kGXz/jAJx4PnVeXfPcw2bTsnzsym4zSmaAaBuoJpehg2RMt/xDUzSuc4iA
Ps/oOgAMTtKCaohkwjHUpsegG6GRhilAEGdcSmg0hM89eFIfDJEf++Us/GciypBc
6KEyv8ODyKXIjiur5h/I8hOITm2uhP3+5C8Ox2p004GaybXUpV3x7PY0/v41CfKv
fQTgiLt4NN7GQtbOTAEa134oz3JvDtT2mfF37hGx+IDXffIPBDr8ur1r4AGaXpaq
Fy/Aah9eqRcahll/KhyS2gjMe7a1AYHln1aFHOU8YowLJijFy06erbR7HzzN/1gb
5a9vJJJF0Yy5AoCAAFRs+UCz+Im5BXCT5RsnERkr+Hfwal2wYBqzESssuDMB6hq/
sInJvQijOe0R8LyrhmZlqtdyIKzPMrKFJWiroTENm1HMZHxk7cMmHj+riYeo8FME
N1GS4xql7i6I0Pfm7fqj9VLLP7iJsOkkTV8Oyz3fkXB/LVZBDl1+C2SpdZaaNS7s
Amu0cIVfDJ7dZ5sr/kzB9ADGZTb+TMspyTtZV02Am2vfoaRV1eq0+1S8A6INR80L
VA2KeRIQmdd1MK/zzjpQuSQljpR35qQOuQVL1KteD00DD5HfgRHYbznmxVyDRByP
G2stQbSjJDOORKxFmNGUe7jN+ncvvu4650RX6dIClQRmRpbF655Gw67ncNg/dwkP
hpX6YzecN9e4Yw9ibdORZKw2e7RW4Aqnb2iglkwJenYJNd7mR1Z4aSdZy64P/RAs
Z5kHmOEGGgFOBdJIpgtRSIe7D9EOO600/K85sgt1gpxLgWFNwxudPvem+c4x1uql
wT+39ssb6r3T1Kkhfpqwl0dsyiWyX8IpoNOsFUx0jvBQSeA0zyJUg/ZxWkHYRdng
mbDxcg6rFx1pJATbKDuqHLAxMaDflfjRxPtg0O4YqQSQ2u4lH70gdVz7O9iIMgND
eB1xPQmCn6pynI0x+KSGOmHiIrmY6iPOTWZtO5QjM8P3Dfctsgu+rOKLo1SNA8ri
4sh6dZ4Vi5BhVJpDF6jlO/gDwjKvv60QLh75dR3x8lh+LT37yfOLGAsf/JevHcEm
7t9PnSXjtKP3I6TuRcsA2afDgNm9xgmf70R1jTT03M/+7fmQq6tUMnEi+EQCsWcv
34BvBsHy+JLAPhX0hAjyuu+xJPS0a3hhllZbpucamZ/g6EEkTrv0USNSaZ3ZCwel
3V9KbxGDUYW58PUIiEk/CIcPSQWsV6or9tVuVAmCXGUEQT59p5XJfDd4n3skoyQa
Adw5ZbpKrr1KcPij5WKtaXxgkAc4M/+BDH4S8VE+etuHNz/OKDdpMOAWpQMFu87v
nvo1BBWO9JZ0Sw4oi+FE3/FhRjAFxpduKy8gkVkQtLByujwogJn0C7Q8JJ1UxZ4s
iEphrLNcrNVE9pUO232OSJcL53cckl1DFpuzPMe2Dnm05UlOO15A65Ihd4DQwAvu
nq8qev7jZ2exkNRDg/2aLIWakafzJ50u93hn5aNIwXnE/jBkZ6LCclYDdgVjVDFS
//U+b5PgNqWLmH2efuHsU1wj6/gEmeYYF+/6QxjyxShDZaAIx6VesF/L5ybsddkC
4KP2sqW9OF0oawRx4DeAXUAtGhLE4y52dg480cn78TAPnJhC+vcBfctalNqDwxz4
shH+eMt7HrKZ5vXX8uPXeYF79BdWsrSg2mCxxWV10q8TOmrwhaihTSTHeG9uSmZn
OXvj2tIZsmywGQlRog+tJx9ksFluPwFLQvIkhIOTC5v1GO1XFL2g912VQu39QvBA
cE+lJGkz0U88OLv6Rf+EEqssG+GQfi2AFoIUO76tAcKkFKANEqzHVgqaA5iyEOKb
hDwigyqU2hl/ijFF8bgfcbM9yW8d3SswTE+8l+euWasVqZ6zbjs/yZe0zJfwt4XS
3Ddge6BA7SnqujuDBCGYz7CNOt7w8unrCTCBq5GbPvD27iCxuRw0epX5c+K92dKP
xqr5Lk2NYeZ7mXnRfhY0o/eKYW+zRYnJgXOWbqWQ+kavtM1t5indk3NVP3w5E1bt
mqwy9hBEPnDkMy2zXGdrKVoKxqRL0QO7c2qvAzY0OTz4y4eQGYNmi+FSpe0bhZH2
dnajaZh+OO41psyEOdJqfCY7QkxsTBrDJNvJipZ7mca6kM/hOtHazaRaaPPGnflZ
KqHhQHZGW8lNn1HigTci+kfsi1h8iqwKl/sEUWM9OdAWPEXcYdgZW2mCWsesT5kh
wbfK7YuXHW+d44IIgcLALzP3oJMdesHhdhfapEeMpafl7n8We0JoWIZshVrJXZF1
hlg11xvPH8hZO9PThw7wyq34crSo4HLFbumHI9Lhnk/dCM6rLgqHhEqnyFai45yN
gX3qAVcoljUetTCX/gAeG1FqxbHgbHW0Da64uRofJei8zQyMS7tXnS8RIMl5VZ7h
mVUTP2SWXcgOI92Cbrz24+LJMeepHt08hFUQ4ixNkKgw2FpZcAUL+FsUUDr3wFJG
Xb+nTqu5bCPO3NAblSYyKLD/K15mwLjiudEy2b58xkRUTGxtI6rt4BhgXeCUHV+f
e9oExbkH/UIGrp6e0iUuABV+rTqc2j52ARMPXNwM+WcUWeF3sUAa0cvDqwJZwHQ9
iosYNOluLJyBaWbaBnrH9a+hZPnDdajHgnhJZDl3n8Koh7Pea69dUSS5aEYo/6YZ
w8BHCg0peDiloQ2dNBObvpZaEujOVP0Aw/rZ2nyLsBhupr1PnVRBFSdz4+TVxzKN
SiZAJcwq3MFrk3TrmcG99HhF8Vu6pBswvfWQD6uXbgAiPxWBXScVbwC+M/QsDS2A
gsL7iiUQ00n4XFIAZnA5jZ99PCm/hVrJfmpCxhtgiLDt2GLFDHomsAYQ9owSW4Eh
GxL9H3WnwKBllMKvhR0a7KR8uZhaL+ViUy8U0edasUFp+uxB88yaOOWIs01VkION
qWCpCsP4lHtjWIx3ppueebzYGehzvYwo+Tqe39vvPry7Gemepl8rGF13dwQgQvSK
s1DAHV3vohOaiCO0MNmRm9tsHVxw8AN7wE9jmsukCg96D9OgHlUTcPEqVPiBMRcY
bpTWe3IUwPcmqn1LDgMZY1klnLuffZlsmwFeD2m5FcWLbfcIyG7f5frLdWYg67ay
J6RtcADNE996gtnGsW7S+waM7CnoVEOwr7cdydiPzYDYM/OTLh5NfCehkTGzYtqF
kv8/IFa8ljfg8eiQbps+TaiokINgZrDzWd7ktlpMyn+/pPEhAkf3o54j9vRtgBwI
d87nGP2wBiN+qR9EfbKCVJgTQd7mS4aYGz6HMDnTfENz0L/TPIhyQHu0yfeAkbv/
Aj1ZKAjPp7xATa70hTMvy3qXkOjnUxgJPgSlBMXzIM6y5yNXs9jd5DkdQZ4l1YO9
1r26hsoXtP5S1nDgNq4qeFty5LZArtHA4jp/RbWW+rTqgT6JxYoCbjvxNljujLlP
hwR6QWoz2uZcQyqpnr5f41wi43NJH9i7TF3sjyVXw4badnD/vVy65LBXLkF6Outx
p6muDAxl1IP781JySS82lFC9aOQgjFqg17KtYJN8A02L7poL5inrE/CMrSK1fSB0
eLvIOApBtYKaYcjMswNGrsZp6rAvs4biuwqVmjEvqzSeMJyWNATK9d6EPMre55wa
bLxixkZcIdzOKPJoH/AQ/1QX6lvfz7p58wHI3VcfQpXxRHKATglf3tMDnO7xqdeZ
0KlCUtOjdLE6ZlG0cLHTULlpWBXhxJGqvcLAgnHtV85YRFFI4YSdOqAu8x8uRLCg
j1oD3xqFvwG9MTJ7qLPoQykmlLyZeBVD5Y21MKXHhqWWLCtR4kULSSi6a5FGcIln
98Nj8g0h4XQqpXuYmAfisthibRmj6i7c0NDtgxgOuB5RPOYWW4CgaxpSpmtmVV0U
qOlrY146NFupmhfvRdQpZxI6H+PN0ZA58Em8CcImdbg/2zlifiAYkVlKbD0mx7c0
TkcIUs9piMTkPlfspVxjDUu+FlxAxh1JQ/ROCOy9qykD9nGhukrbgTIH/lczSAEU
f4jIv3vr2NjSFIYXx9N9Eq96Wm9IvZ4XTF2el/QJkM2xpvWKK+xIdPaeFmJyz6Ck
7gEZXjNpmx6XPk0+cIFLpUvyIKlf82EUK8It0pPqlMtjnEG//U2g+r/dNy3BIZWs
x+9DgOgmqdq6mpszDaZc7w4rAIiIQujz6ETQh9ZNsi3mjOBuAbOBFC8FQ4MOTmRG
rHTdZBS5vbNjLDaG2luGFdJq0rJin3bNshMVHBAZIQ3eYOYwhEoax05tIFfnm0CG
NIA3JV/yMOHRVoVhoLZpOBk8TIw0jfqkD1eJa5z9A8y4s4wr0JwebOr7gQsD2Z+/
V4ajWQWUQRbWBUN1OdBmnbH7IeHY4XgM9zXWjvA7HERaiEVD2U6q8XR7l8LgKCXJ
a/N5awT4AQ+dwOY6qIcYNqNyuu5zYni2QofS9wpNXEqW/rQvEPywm2fvVQ/0OWUn
ypufCnwho/lNZyuR3Zsq6E2ZCZsQ3VM6UlB42ZmuhbhVcStS0k1XcoAZCpjcdDDs
T693YBH319vwbWQSmQhbGx5hW0S0QDnXoS1HtuIxkiJVcEOlZ2j8QkmJocNwXVHi
v9ra8DoDrTzBT/PjUWxV79mqelUqHTK2aSfwiCG6Za545DVoGv2QM2uj43W+xmSg
oh4Jtg1tvM4izh0bta73KqYCKsajP7HUe8McuRz/JF5IE8DMQdlGS9ZnbsZh1WAl
YRu/BgUcDiYOGzLUYUyrsYTEIPMXqzxcwmgogQjTJe29kxM792d2oTq3FrgwkiBi
+UjRyA+WtKHZORXVUiW0++QBKzjlmGjUN91DUsxV21a9+cUPIKImrJLXNh2XtRKI
Jj9XfvdvQ4nt8gAI9IzLcHTLWMcLZoXmisAFO5uy2J2immq60pRg+WvQ4QgUDFWg
Ng2Gpse/tY11scyRF8YnhYNDdrx7ZgExDIBI25LvL7w0CxPOU6mcPIKYCXy8owXV
V9dnWLfz7Lq4/ymYZ17tAjbHKpoY20EYMGCOZXQZNiMtf34MuCHHvSGaMcC/YZ1p
9uNDzWJXWuQELzQahzaRSTKKQHnWvkKHYHtYNw+0ArZIEHoTVKBql2wQ5IdngNtj
fPj8Bo+nMuai+a5j9VDSTpx4Tn97kbSso67cEp+rynyvc8WNuIk9TDwK1rjv6qJm
svL54UV05ba9Y8DfMyjPg7WQQIJFh1qbkbUhUsF4OGuV+D1jYrUNKJ/53Z5Wcmma
PrnkbN0pW7DcRHJ48n9uciTAoG1u7PskHTj+Z1swrcRzseP/I5FJldnh36LfeC/0
zeon00eIaYDjHayADcbLO69O30P1P7YS6qFjUv1rpUzmn4P6jMks8eaKgeteYmQJ
gE2dEZ4+7kGZGu6IC+JwaurgN0Xm4T1gR9mfp3ahxS6+ZLub5V4FKnWkmrhEe23m
9+fvEBnrQrtlUMlVpb8e4jmUyAEt7EOQaVXzFhqCoXfOu59zMK/LjCzHtYCz+c4L
0taFCE96eiUvihzmX96lfkST6bkjIJzBUQBd6CLTNeNm7EpkKadfCOTG62Jd4MyZ
zoynQYhzfsp4FPrX+YNPsgk2u8Hvd9I6M4zUO3NsxDlFhoq3YQyOqeuGNXmnvxNS
JYWNyHyKLsvFdKz/tjuttdGRlxRvbBjmmNDlHS9yUQEwWbg1QLq4c+4piji94m7x
JcW+wmmu2IdiKZB1k8HTguNw6A4RlpoaJFZFC/3MM/6vob84r4GeUAkB2cv2bhMC
yuVwCetUoablGA1kgB1Cf4TP9NpZdlBL9srg4e9kRvdNvrEIeFYlRgAiMIu2//Nf
WaWASCt5FeW9Gl/PrWPRUZBEp7kfJ1Ji7Eb/FnOjms7y1c2/Mq+60Gka0FPbAv2x
R5LZJAq1hxy6iFOGmmT3r6lWfMt6/9cEmHcE+qFPF6aCI7Ce+qoB+J4WDegrzbo/
ycjKX8jNtUx03fVQD7ZeNd62zmJDzbAoMldVh3CVRZqQvqp3jsn53CJ3oERaQh4/
hDpxc8V2h1ihsCBEk8N6+mpTdpxExCcQ6VXz2fL/j1od/Gl7YFQh0ITIn6XZngYN
gJkOJpPdCNuHdM5GaEgKod8IKEr4BruZotsl9c2IRO6ZH6qUozOD+/HDlGVUnVpp
OWU7/g8jX1yKdNVQ50BB8DfaV3Z1GocA/Nisj5qgbBuaE2rqF6TNg41snhn02q5F
9IjxijKGjLbxVNdIkMB3slevNAiIUrM5Go+Ih2tA0iNKMVwIv+8tVMELNedRizQI
hDegVYaYnQH0Q7UPx2BJIYqh3q1ijl3ITqPytQD++gdTLVFzORmnbcjT3v6RaDii
/kOGfKlgRPo9ODjrcp5BHc8ilJnvMJmKS7auWFlPKvY9WBupiwaOXWQ16fn584he
cmynDkAZG+pBFvIIo3MPqnSVIgMI2jkHQhqUYwkpJ7uy6LTbf+QT47hQyvL+X0hs
sMLhuCrCg0EPdsH1UwdNXmrYv5oxANdSbq3XXkIhbupcIh7mPeSoKJqVXdsXzcSH
pCEv5AKuJyaEIShQqoYnfmC3eQLaScJEgI67RIJT98o4ayZj4Ls+IaQUXDYKcy+w
xGHQRwJqac70xQh84brRMW7h3ZYF6klvJFPad71P2wdalK5yisMDvMWgjCaRlIL+
AofPFrqDSzrKxzWIwQKhKHlYkRatc3dAzdsjSfVXLZ/nUxbumD8ANBZVQCGhTklY
qawtdAFoBLLzraQB87rtNkzP0Z8oBLuH40i0buMKHW1shHdlSaSS2mv3pdUPTIa/
1t3n9+ajH+hcV8+UwDeZPHVi4ozvrpfaKR3XepmhS3BDrl2U/Rj8zMFCVCNo1Adj
RQ7+ax1IF8/OGmWKfTb/rynE8weL+ajl2u5bt1TopvcAWUAbCW7fBuweWDwMPLsR
m5f8zw//t2AgU85kg5XeFrfuzXdiDB/XTiirrY9omLgO+4Rc5MBlQ8aNpNTdeVmH
2ryRDKDU6InXjbbB/7+LNXTmifH0G9LesZD5X6rXA1lEYkt9eDUqB9ZfZ347CbT3
Aae4i4AwF27WvsprKyCdXnRTLMuV8ebNty5EJuK1GjYAvKxqnPIgZV6kzgLgqy/3
NHdO02imX7KoWBtL/LX5QG2Qi8V29sA7l4dLW2nG9xyJRErQ+q0tEwPmXuad8B/n
JcXUabvh3qJiJZGrw5KFhiEzjDLTNOfa5kiYNgeKX9kV0vMokecP1InWZEW7lk6J
DKBC9nYCju7cLuZkSjRkoMvrUWNd0tkOgv2dxBd6SOI9E5meYkklMocMTnqcjHfa
fCMKOA+BXNHvZ+sYvJhv7gWLuHMYIG+2ncrRbZloteHol+PWIKTV1VQ1x8wdv/vm
kXpt7tcWXQxRJCODMXOH1zQcdEzr2GrEWWs616OHQGz4x2zs9qVL5AkPYElEVxpD
ayYAecCRgcCMbhS1WLG9oJT4AcrgsxYvr9emk9hokhOTKQgaseYvUFbF23Fcb/EC
3ZKVyrMwWTSo6LNU/igKAlwXIioY+0kXhoJFAg47O+InF0DqHGShpJhgTboBxqJh
x20+iYgvYd6Ri1Hz/zV9md/GGXanNPhbcaj0sZjq4c9Rh/mjjg/5kRRyEvwslnMi
qW63pTv3yOc08Iyn4s8rySPxNko/bWwL5nSKkhW/h7KGqZefzaN8G43NkQgNi7ed
qW8V2zEZzu9FH8kVlJlq+N2CoeDQdyt8wzHWcQi7Nh2t3Ik2V7zsf5If2OwB9bUt
wz5uhB1i7ENQDUh5vmtq5RzZfmBb5r3/B7L8kN+YnATURgKLr4uVNSgXALfBh0SM
mcgmWSk3ylYASOIO8c7U/BmBe5HHFeOtzEldidgbU77snQiT8bVJgBnZVbAdivg1
gmS1QQ+IABs8miHNas7Jp314OLGiM/wt00xtUvDroSesZwFVbfw626/EZdxT9W4d
oaOQ8IU/GSRdGj9r01VhAEMybDSpmc2Q8UF1PS4lfhO31cMCDGdrds8xwbNRGirn
l4dTLPN3YBH2+Yi4uZX5vtVSDlC8Bg3gbLvWK7zmOmedAgfVdUyrFlvB+hZSwEOm
0svbIYOLRUCkpURdfuiQ7YaLLPE6sWpmNpYubgghaqTKqvtXfY7f/8wE/5V5G4x/
w9zSjl6jgyPSGYgbKHatLlJPnlLFHrebwsQcz/ohu+8dkrJC44q3sSdfNBrWJXSO
LctI9wUWGDDYa9hYfnx54kqcK8nDWmRqXRNGKoXLlKoLvKmtRrUrvq54yvNfklBu
QJ7CyqUblLs52tHLaBAtDcKzsQZZfnu5g3joDi3QR0zb+jFT/H6KNNM21TfxbI+q
Y2g2sQbh1G9a3IL6hVONX7PyAlqT6544UzgDWQZ8uKilMDosK81Cthjy+ZxAl/Ec
02UpIZ/8Ug2r+9ZYvuKsxEoqEW/NgnVYjnUIxv5TiLbPVoRcj3S9q+nQzFD2bT/F
MwqU+GADP7IYVUsktHSpM/3twTf808Gs6rYWPKX8rtF5U0nNW5I5abBJzysyZJUK
sOxyeSuMr7++W+s143cuHErLi7wr3PTWVSZ3nnKHkrouPh59HKlSjJgUAaq4HWug
lL8IFsu0fZUWAfFFiZxz8TEQ3vsnGF3AziCqEgBK/M/jxxAcjwUI2KzmOJrTY0Sn
H3bVZxu2WT8KNGOAL2M/dN1TmL5ppV7O0R0+AY2wYHW64rYvAVBbH6doDBg9GkLe
Hab6ZtidPOw5lf8l1J8zaQvSPN2F4ofD3xZwNIvThV6wsj5GU8kBEgu7iUXfjTAz
ZsoxiYNXoJVNuFabp/7shjWiXLZo4WEgEjNRlHpqS3ogGq3IJOK/sMx5H+zzIBpe
RcVE6U+wgA1DjIiArT58LVg81sro+HaVpNIQSaWy/PfeOfp4GS/7fLBP5E1Mb/tN
xu7PokOw9rQjL3UlWEsupPUrm8A3eMk3BkzkoKOpiOXV1Wxx/LFBdU55/sha623Q
hxEky21ZzRT7aqNZUmpuG+Bns+VXAsRlxKgiGdF7pvu6xPKuyn8AgJmzuyKv054w
nVWnjb7oZ1QfUBPjA60UuNGCmJp5icwPT5gQF3fqkDIB/E3tYEmm39Q3n5aoFWk1
yz5lM8ltR11Ok2HKu2HO8GFkPtdBno/LiOY4W4R/TprCZQAfEnEJ/YuBX79kpJIL
UFlIVg4yJRb9u2b+ZmCWeXd8yUxAc+Z2uJEefvHX5tiCcqSDm2nu1L5YMlh7Q9sS
lt5B1hhPhCrRy8psZs/JS9/5czAYekaI8sNwn98DGMO+/X/fbBlwkKHtCU4+/VNo
/qTFdIGSV3hICzs7f6Nj1EU7OQC5d9+n34UMGAiNU5PTwqVItfU/atLqz8lB4hSW
ZPHraEDvC7vwRx+2i1PIL2VGYjNYauzqHLRCxbZ5YLuh6XOyVj5JUo0ui+xuODVy
s/6rPtO7RcsKDzkEMwwGIw7aiYoY3bEnOk0Kkt8DOnKqhO3aNkmodSMGpgdpD4zw
J8kT+ebXOfJwNooIl0vmzMXMHNql6chqiPSk+ce7adTOeI9r60tnUUkMwJFJp19V
Dw85kJStnXTYRGlHdWGkYVOXnD5kajbqIXwkvA0/AbT74aOxicHnua7NfenoMOOO
MjXwKnkF247ydyGspKNsYp/f4hZrBrNpHlKLsSJxUruyXsWG5M9OhaNwbY7s2wgD
sofNKrsfoR3ldfQjlaCfQ5IKHGv/WCqplmSvRxHdpR4e4/NcK7XifLTvsQzk1SMZ
dlYJubZd7U9qXDbV++Lj1RIA8jfOWHm4y+SYWiLUbZB5xpj3ZtZfNMUzSyeTE3vj
f+o2tLFtiKJuEiD9C2AfNaU6B5CsVt8dygea219w8MB29aytsgYVuAUkDNF+TL8e
HjbfbXNnEVDYlS7y0d0jEmSzx4MiSh3RgOntqxaDLY6rJ5io9F+WrD3JP4Ve1sZQ
EQsP16W/bcdrHU/gcs1O2qwBw9Vi0QR6Gdxb1eKB06rfmspP/3DJKus8rGqJYKfj
BD4+Wh8PpT3AlykKxIGPxTGlhGLngTJWO9PDTtJIYc039Pwcu1xCy0xKjP9T5AOs
m9KUbRBr1zCrj/aTfsZogSRcwkJ4JF5thYkwp29FSX+K5vqdUp1z3TK8tNfDf7VG
T+pZhWXAxrivB812zXwX94P2wIxcK3ogfpFlSeMKxKnP0twha1p4cEQRrw+vRPG1
gcDOaJE2cIcZuA43R/5SoTnYijHLXIGBpLbs02egZSc8jd7lVItZQQ86zASPlo9y
jbwVkLrWjr57yPvSi848p71hXFpW57n2ttJkaq6fsrLOAf+DpbaYnR48Vr9rRU83
vQbSM1GpKYnoX7d0/GQ9OwSWgyNyktVDcKXveExVB84VtmlnDUBa/q8mM1l0rWFH
jwNB5+wvMkYzsyhyu8+BA562/ZKws1eSoetYl7MONWk8qHqLrWe3kli9CsJDjzzF
UcgGMMgzeOfMcVjdEMdGHA0fWIOWE8zFKCKD9SlZZCOIndVIC/DrMcKbaTJKWHru
Rd5lMLh78d5UTCIf2tkrt6luT1wg7fsYb3mTLsVSAnRYzvsr7k1fiK5E3gGs08Y8
KT0EpEnaJTwgGZbzLfp4Jbd6n5cqdRQdmX4zfVlGgm8Blhi+DC6bDQxPtWj9WLVy
qLFxlh4/NX2e4rhu4Icck73F9kIgGpgk6m45wI+NOxZOJR9voaLV53piaN/2mjUm
6ItiW/bwHNcPrnD0ktIakLhWygEaky1TLW/TruJmZ6r4RV4sw21D7zZKqCImX2gq
SarGNgENmjQza+CsuRB9PxDPMRB+/78gzbm8flxN0CoONikXfDtpfAAp2QFzh/1Z
DWv7sTI103phyI069IIpv8v5Lb9bkQl2Vbh8wPoTkOl7xKC6oX6GYN+HLqxMhWPa
QsnzmqxIw8DgCHGFcSh9OoV64FtFBrT3BwBTcwCrWgojRZ3gvuqxhJJLHorK/J3D
wFCrLS/5o8PivDyOIJC24iDuuEDFexmHRwMutv/dkuSjeDpL9SgYLup2hgE+r3WZ
hu+I8gULlf1wVPfiko9JWznS8xtZidlJ/px5SRn17eBjL+IC2su3tIJhp4tisjqb
oyZuNDJWgjqlUzU+OR6p54lI0qnAJhNYv20jS8TBPNKO8mNtW9Fht6bMzvHznWes
T1If1HV7ebcRd8wIKaX8kI8Ykx3dSzmG36WUCuYZiM8uOcq4hf9VE+HuJizAoanZ
iW0D8iXbJMG+tNXpwoxFWJbC/g5InjEIbDSQ3SBl5xwY3l+rMuwQea0WEDkHlmgJ
FSvkY5tZAQahkBY0ux3i8v59/WtFsU2WDmNgy1XJk+t4wd3HhVt8rEkorbhmaFYz
fPv2Escid6G7sM2I2qMWcDrKAGkzMGZSPGQcS0A1lhph1LzuOUXxCgfNYXbyM4KF
6vqEopvw0c8uFaOL6Wqz18Bn1bQirhtKkK5tw7ezC17z4LFK040j9bPdCyGoGlc5
d9KLLht4Lm4q9z8Q0evVfRNgl5RWl16Dopc6eFPg9VdMUizh2iStyrpV0BGJAVq4
bEvaAYrXdsqMeuVoUh3wz93WwXONgm1gd15fjICeWQ2Lv5bGFMaREQLiVNX7XNeW
faxbh679h+jei7RyBb9sVsgwud4Ohk2PjGcQAl6pZHtMKUwSjJZ41R/moeqcCiMm
Do40m8jj34MSqVLgG0yrk88KdupntFLOILZZFk8nl5CCqEeh3a3eTFx8U/RekBkb
7n4hhHJdJNJ0kfj9Z8qX0wmTfCRUDRuCd4vmT9wDsvnM4BT62nlG6r9ym7svMzhj
zQRzWFOvwZmdLhDS9Ac10Jy9QN8lN4FFqtbKD0OnrrThJXKr3EKeuykRgxxqvsN0
xoy5w1hdBU3R9CmwikIZTTOILx3BI22df6CqRg6NEJai7V4FuczJ/4InfWUgBXui
5uV2yIKilYKdy3dJy5Ae1+bcciN+br09mFWZPQ73RAib8dF/MkAHuMv5lgQ4yDPq
qK9JCFTYJ5pafTgyie4Y51JeKh7RbPydPoiHs9EAXPkBchzw0idKxR0UXbMV0xGJ
gRkpy4sYUB0xTsGxEnZLY0dF7jfpkbZ0d04GGjed+cjw2pJKxuZXntrXUb8UmZrn
+4XAghz1EX33+SWA0YeVKEw1CjKtKmNzj98o904Cg7OKs1sKkkAx4B0DwqMaLgos
KcJs1ipbSp7JcT4vXC/KE4yE7jbfQabEP0/5XwLJwXn1g8GR8vIEFccbh10T8xqa
hgExpsrKeyrnzz5wvtnDbBlRXZf1alzTQY1yfxjgFrMtn/MmLovA0cwkchrTF2o3
MxNT3Svf3Cnb2ZXR3JzU21uG32ovLDEhOdnbYFTWV+WTkTQBzdB0keniNnO/2IIo
T+TEUkb26lcF9tud1535BXnvLP60kA+tjimznySLPIkExYmkZ7r1VaLaKJTuz3Bk
6u1Z1ASlmtFmtyswoG/TSf4CWOE1ylHi1Ss8l+gRxQGYhP4s08qIv9prhs0k4zIX
1ofMYRAtU+iVg2FUpYKVDvKC2PkNeP9bb6FHWrKD55DwissXpmjdN22w4xtju0sd
SQXX1NyFtGDgD2c8ganTFno160oeAAwKaPWxrOlC+ZIdfaQ9JxFIdiQROVbbwsHs
z0NoB2kkDCJtN0nLWFkBr7qkEt1InQPshBCYKL7pYBQzBwai1CCQJV+eMSVAUq/W
DLXMkm9HqXpkgxdEK1DZT/bgmDP8abhkposw9sQ0dEBaD8F+Ocs929laTjUjh/sQ
xq9BSehXYrirBfKdPepyyS9hlZuxN6IxPk7xstQbBmmlMZiu5Gi/6EsCP1DshgPl
/kbz26Q5OrA0vBOhXR0sOxx8e8tqvmnoYIykiL5BpVR+th1Fn/b+a7OJMqNbmHFk
couZNFjIxqTvqaRjf2+fkq2a2ND0BplVoGmchA4g/OqV1I0OpVox8tgN53+D+/GT
B7Q9dKoUTejgI4ivBXB9JHadm8e/bN3+WD/0WMWTHANT6uIFImpXLl0yZ5LweoyO
TCGe/I+XJJ/L+4iwdba5wsPegAegfQLrkPuNK2kZBoWVq0yP2SlE+pFXG2mS+RVr
F/xpN5q1l+foLQJqmEJFjcByx4zjPWv1zB1XmBYURo4XAYkXMnllwPQcKezxJ1tn
PYxLnPPyFcUuiWh8+dKYBFBJQXY6pfZc+Ksv5ZdlW4uGx/q3+Y19M0ggqujp2dBo
2S3Ee8eNtDX5YYbTcshMMLyFRZabbQQkoXPwXKw1XOzZegoF66XQvbY2G4KJRy3w
XvKSCC1cZqKIJnTjiFXt1eRcIgQehdGF2pTDal5vOCLH79yFq1PkVFzbMZ6rrLrD
aHL6+LGgCNUHTbJZnr6HaK2Uf32ySMSCbpxpDSo6DjcaQjGI2/q8CVj63tCPqjFA
hGeD7pwVj3xuliuU/jTPKZhGTt69LQdA8AqKx+IGwNkE1GStMJp/EDeNwvc+S48R
WXlV+/lzgndpOVrGoGFNLAdCv9z9IqGkSnxuzuEi1AUzYLNTXZLirf3gAm2xXA1M
JoPrn2N5QbswJkZ/IUuuVJA3V/9SeLJDXQPZ4XdXQpyhGCGk7DkEhhNG76i1Kze7
OR4jDVP0UNtV/qdSlwa7bPXBBNNJRY7jlvtxvcBPIxgFpKdtkE3YTrwJETHFJin/
sF0RAttRtgsNMw2UnpPFRhYTgHxxkJOLcqYLwfu7O1zEh8HZJAGcqGg0+TojJlQt
ydJQlSaWppxjZ+YN+TmEdA==
`pragma protect end_protected
