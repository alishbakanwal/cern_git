// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:02:17 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Bfi5TClJUUziP/xS7k5VOjbCFyGP+K03ABOklhWq9UIR8leZkbu/5uV20uX3Iz9C
AEr2I7WNWzFKoKu1i5XsEb5acJ0Lm0Dm3sBRmJYcmA8mxowBnpJgIDAbVaiM+zif
vKHfjCzZbIYkpUGv8c0j2HQNXH4QO+THov/yyV3tF18=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 50816)
0gkFAi6oiGvn1m6Zkh+T5sU8wQXAxcUJxZQjmutygiwZ+F5VgW3bmv8LOUF8bG3X
27fH7ZQL0yYEr9yIdFdYJS963UtKFI4h7Nz44lomarIIb1LQwekHZRnJqwM45yxs
+U39OJv4vQgfHCg3GbwojF88dkEf+P8tq4tyMvWbkA1MKsc8ATD9ZEEYTzLeLepL
pn27ftR+UecLSqPvRxiNJMsVUUVGSe/PWnSlqIwgu7djJL1yURP11Fzxh6NskfZQ
9txL8FVJzk5mItsAIr2DUVDTCsFsz0xMKL4lPwT5qFqxXWwW80C0Z2E+UlOTyo49
R1SkvxjFWCtKxQ6M1kV1/3OBKT4LnUGMqOmf7UMHeHIWs5+uvDmI7JB9jlpDArEe
jqlrYhDkPlDYSZPKiQYstdOuzINab8vYkGrm4tVMl6In5rIQNY0alzi1urquhcKg
1bhz/AgMu5Gm1W2Jpp+mtpXS/RyG7yPfMcpx5tMiTjQbnchg71wCdFhkPpaC+yQ5
qbUskQJUDEi1qBV11lvjAAfzN2NWagfjcn3Wn/CGMgV8plZPn94wICnowhsppRP8
1ZwvLlHr/Ukb1wNV6YOzDFNlx5scCIOro2DQh+U9qIf0VmjWAXMSegN/i+Z49r9M
84hjZM3QSA2Mf5DsvP33F/XIBC5FHyq1ZkJXoPCMQHGKnRq6WZxayYXKmKeKwVSo
QjLZKRbKrLtb1oMYK3Un4rJHULBhF5Ct0wOU2RhjhW2s0a/4yMwMBm4lOK47jLF4
gnsiJG3MbntqADopb7R//4LPuXvnLpvK3UbDfxC3S4973Mw6EaFeXl+/wnM6hPGc
sV8Kgev7sDDX6bMb/2rlLCP/ypJ1RTqjAH1FKvOx3w+xsqh3bzvyOM+KuZ+QwTlw
kN4kKV2Jw4PS0hHSkYKASnlZnjrWhmEIXjqjXf2h947w6O8jG3105HaNQOES2I5l
qS5/goep8MfKnfomWi9Rm+fenlQ1wzWvpAgX2Cnh4PXM8T50Zvgl5ElB4RvVh3ia
5ixdMVOxB2+TmuutHCD7otL3PHsxfoWA5tqt0JWz4rTV5dGTh3GDVN4bF30RDZFt
M9etMDARo8jQJmVaBadx1P5o0RrU8e0kwhv4ONU0J0w9jdOABipBmyspK2zVTJSp
4KdS3GZqU9ochpbMS+IgElm+M8dvby1GNPgHJ9IpJLi9/nir7G5o9qwrklgFRvuG
q1IqVKsaYV3vHOA2b+526Hme/Z1IEX2BPABh8DYX5vFBcj7Ex+WM47MwcuGBvQAc
+LJwIRrvKaTTWJcYXeu/AlYHwH1NNECBefu8gkCyIQyu0YSEIr5wxkEXcMU2kL4A
Unb6SpqfR/Fv/2f9K64sba8WVFi4OsJQ/2INb941yW3Qn4JgDSVPOzpc8vBmG6Sf
a0hQQP9cL1vM2G9Wk+XS/kb5+Se/qdrYUnKdIGc77t3s8ZObe7Vw1itfFW6CJdle
q0HzPtTr8C8rPU6yEysyxQwmGiwIcytqtjP1/ECllFGTzUSpdEWUN6Jcmd1IyHzH
HFH1ZbIiZBmeyIohS/uZVQ2NLCogMq00amse3sKXEd7+rdMbOZgmQXLs6jtqRM1L
fwjbCR0UF9hc73JQ/qhSNLJC44dyPpgYifdU5JunSXJ3wVH4w6nPz/ZwNV1v20sD
SVTH9YnwWFxQRu4vOA+70dogp01F/E9xHUzHJ8SD1nx5pKa4re07hWT1Uc8gsX3Q
zcBxBFGOX2u03Lz5eNuYUiPVLLKZpAB7DcQapjGlxym4lnROklJnjwKdxIgEMLqp
4rqmEbIfCOkog6Bung4f1X48YAuh0g79bMvWQ9WHeZDo7CQbznWGxaWJoAQACv4z
Ow/DUZZ7yTlm1Ohu+4C7i8up1h8EfYG4QIKkR6spLcP3Nbq4DcdE4g2Me2JEUG+i
HZvcWUrEr709iFZOHRYWXlIAcTPfJ8GPQWuTN7IKxdI+gslZc6kTuUCSR21/ZOtw
wcnJ+Q9V2CUKPPH9nF8vg+kv+I7FnfCJSstoRFadIuGjVAaDf1FuzrwyNQd+CQyw
EtxNG/2unyjD8X2IYO8mkVcZZMbIwFGZ9RrYbiMO90behjdWKUK4GV8jJU+mQohY
o2bt4ZB0VHT0WgZfzS5TF9YNtZUIohGnDs9fpQSJ1MRKcBJwy1+G5Mj5QCuODvQR
J08WOKsMq6I44lRujeFDlfOffLhUlKF2Bfs5p6TIti+iuUlsoT724V3DUgqC1KXd
oTM3D3geXmOGhfOn/nPWvVjgiEBmFuTl2j1AFmdGi8mqWC7DnDBj1Z3UwaqclPKw
JKvc06WdqD7nS0U7dyNAh7dmlm1a/kRbPUYn5kCcTT42nS9QuMGT3QeDpL0K4Lyi
FznbyLSwG8LAZ4AhOhXwXM/Au/ov5hA02RIxXPCKWES/DM1oU9jmcdWKrXTIAAUQ
GWG8vReVWBtZZChotmzc4CqzoubFewMqkePc8Y9GI9Ez9eMEJRYhRkXhu0vJmwFg
Ykdt2ELq93RBYJlGW3+5Np13VvgSzqZ1OZHipbAhaUIjCtR6hqb+GVJXLebmpTwI
tOkR30UfmqYoIch875fERELG937OnSj7bTnTu2G5queVOM24sOrWamsCmeb0znid
NTWxdTJ8MaKcwaAQho+O3cWwwzoiG51l0/wgNttTqrY/lVxKres/9BLl/3fHTPjB
W8a5gMloJiRsa9HnnlJ2TzwjG63/TIxEV5w9iNPG0HZBfpnnjBf9CZnvt7r2Qbb7
tPOPuz7dmXTFBrr1T7qQNDzA+7VYmxHag2m/nHkm7TdcZQpqv3cQvk3p5ULBncgC
lWaeBS5r0yVSFqkzUW6GJ6WREbFVlYhZHLUwQufoAwtZm4SOMZhCL57DaGjPAVyK
cFpMNT4ef+lf0OyQD3TNV+WA3K1PH2jPDxF1gkd+LQnM2DzYhtmE2mKIaHlwCacS
d2jRqofgLvQOrnMjinkMwKxgKSGQ6OOWzTeAC1xvxEnU3ah3RoY1KZbcUlCtOx4c
sTS6X9ieKI7Sfp8DXNIE04yiXH8SCoksJUFWhYRhX/uIHZibhoOW10/0UE+sRqty
aEa44hzqXPOL3W3g1Qz7y/BkqbdkMtx1M4qdbKjBq3qjAA3kG5mZ8xxCmfj31po4
0ciJSjQqWP0fNMxPcWSIlBlnOHGNQtrCqd7K2jNcHN5aur3EjRbuUBWqqwjILihn
JlqGtsxKKXfRatfjtZ84p+J+wUOd6OVsOLPDEn8I7MivEyx1rOT14p38MVlQDBaP
jCLpwqcg+2kgqCQrvDnCMvCJ1cFPGfH336prYbUtMmSaU5IKFwuJUpfmhIyV4FqR
xIN4r+Phce6wIyb2bU3vL8uGam4hGtGR4zKgnFPrOaiRmfZGWGwPrA9zug8KxKJI
dfAmQ7L8RoozZGPLJK/d4xm9KQ4LLDZvxyUJCDx3w9ZJj/9SszqQJOuz5NEXkxYJ
lFhwwrN3kxKMt2Np/uOoNekxb1Lydx7+V71DjzUsULUF7Co7uMBK+uBp9ry0jhiK
04G8+ppKeN1IvUWQkNeOZ1662u34DZhtftQi/TODfNq/+mUbNZySBpc/WSsxT0Az
ceaWqPbg/UfDTu/mYmSRT3T9R2hAMxb0/nOAvmLWTi2WPAdYXP+L31nzpCPJP+qV
oYoebk66tvg8fnrADCFNXnnug+5XbibAaWO1Dss6fxhFZdhfsaYKh4zvmRZd86NT
ODKGZDbnaePosNf6Uqf6g+Q3ufHASnrsllXP5fZzxOyNfKtrikhRrYXsgs4MINo7
vdZ/NVdnO7yeb5/OdqIYiR7fELEAsCDsDiIEpZ1FMH2Af1JaEmiJH5cY12q7vGK/
htQJ1gREALSemjjWbgxJ1408cD9jI3HxpM/SmDjRv9nCFwZsMmzHfOUr3f6G9N76
Vhp9XMG5lKWQpk25sZMhOTKtM5HYUlFVMLJ4NuUUYvsfX7NHQO0tovSab7oPiyDs
h5xI2KvZ8JDRckhmZ/zm0zT/sxDJu60d20+VPBSeaLQa887BSOUW/af6HEb0sH7N
DUsuzhk03lGepPlxHNWBBsvAgMNybB7hGyC1/JIt5/t00tMgsPIsUcfNPFaaihk2
kUWBO/l7HV1OZ0JrzLEI/iIJQ9DXwFKnXwrX+3ha75G8zgl5K/m3wUY7urcwgtV1
TSBtTu95WMyg7wB3wUsT7zfQoGMMliOyjjqZDpK5TUBiSvxtmnGwdIqV9uCg+RIq
mCPouQ/0IeypvcQfZLCCSZY3WfMaVWttYzmoSKEhDTSJrlIIAvBeCGQXzKI39v12
eO+Sk/CLBIITcY3lbDiX3Ycgj4mCv7+x+aVHlYgTrBoiNk2WjAehHcvYhCNVkK4T
zBzuZ621NLm6jH8/vtaUPFF9AbbDSGjJwa8fZzb6RxEmXqLtGIkCQ/cd15RNgDxp
YY+r2rXNOLuK8bpop0ijmyM5Q6NSRpAfgO4zFlpwoxQbbFCrJwE9TOMpf815Fgbu
+HW5ii5fnp8nlBf8n5GMPOe3h0sBQwGc2fUu4SDM3LftlXuGFaCTcl9rZu+r8qqR
5i7FpP1GJZZowfRjaxx+VBPlRSNrj1YIwfYGgruZPZA/rcTAinqYmRn17w+NE2Jp
6jtS45oVU3dUYr1ChitUKkpryai7/qIfDhJER90/UJLJU/v2yAa0UZ+p3X9C3/Vf
TV/04esh3kPGJXcKpXg6saVvzaSpfyLRyuQ8vB/lk1/pmQamrEtD1+/NYr/ilw0R
r0kAmTEwjTgmfVDD2186SCkLl+ux5t8s9Z7scd4eokBGB8xtWMPoWd7Rv0sPCt/D
+DO6tgPjmaSZZSeTB+UNie5W/IIAq9DxbikTgnVUKo1g0Drt412Q5NVw4biWVEXm
P/t1Yl+igy0PfAeSeVB/zitD+zo9i79szzAKWLDjTLkQimWtjxEALYABDa0U3IDV
O8wHmZjur8RN+Bbwatjt1ICnzjL3mM1kFuVhuyORZo9EY33Eckg0UI/9g2bghfeh
iMVuYKWfjfedwmg7StivcAwKSIAqJPmysV5uIXSdSW0E2aRS8wNkBCwOgvGsp19Q
u/KWgc52Hn3/abYxMhgOoq7O37HYW4Vy4VcaR1ZYU3q8/DsLgdXmnMAPSbndGO6w
/OrsLH+qMDO70xJdJZz101tS91flgpQyDAHT36cuPcKvLvFCqD0SL07kjqhM4NO8
aYpcTVEMF5mIWCmmNpUcRAiZHLFjxGsnzYbYzyH2ehUdxsKOwaKoVwT4+W94eoRa
x8PC6hYrtX5DWSybbCJg14W2zkTDKO3jRAiBuc9E01znSsNE5IHMJXfmA4BCITL0
U2bIyWo+eih7QvKR5p3L+8G0D0vnxz8wTwm9S4jvKw5MFdDIwzRb0LZbxeVbV9Lo
JKwM6/E6PKwtmvWexog+LiSIuRLG/soFrjhQSJT7kxe8F08D/zdSAUiqPT+U5EBU
tecyft2iovQb68NrhnE1DZj78fSt3MFGgUiJje10Wbm6ShhIXaxWHJJB/UAlCnGW
GadkH76UUNCJNh+3kNXYmM9z0rITvAlVx4gYYWRVJefYIpdymDnAepyFS5ZfH/Mu
bGrmBMkkpqAbDrlN9RWoKpEH3B4Ek1ZE6BohJ2liyvhHDlTRceeToGrVYZzP2Cyk
odK0PeQabtZ/+x1mxgY9VbhKffi3mH6VJdX5M8OAuN5TuSVvOornpkINetQ6/zNt
+/o1e2VsYhzKIvtJAF9PjoSF/Kv2jTWKgz7VcNLmETzG3n3DsOWDi4ZoAxa4ktXj
u0tsdr0dFUvxyrpN4iwkQSGY5EkZ4Ow2nzZB/pwoUwTkStDDbhs9RTQNML7Kdy8k
0oBSYtEiMhefrUL66tORBLDo9Vo0aQbI12u6oL++4RndCrW6qBjC0sbmpE4SyLIV
iO5zX+OMWa0qYX07y8lrsmV41D6Bz7UiBQ7TXzMrBjMjH1TUMxFphODC729J9olT
HLuLfym32MQNV0xSp/NUwwajYzVaPD5QSAryML3+axm5i0wuG2MlBEpiA0I5kRaD
8ZYJYDjYx3wtAIG+0If03LjIUPjmh/eMp3MebaLmriG9TnFS93BaIAH0tlE8Fbx2
v1QK79fP+Lt2Hf8gBr3WRUl2Dv8jvVCyP2N8tZip5HbOBbsfIT7GBEYq475Qi4Y/
+5lTKmFjLNNSeXczgp0RN+MCm/udJRqqkplEeXcNcTPffLQAoJ1mQoJgB4DOyoKL
0b2Q8zxUoaVZlHzoEze8XBUZJasg/KdkjHhI89tPESDklsDVYipMOmzAAIfcQMsr
mR8jpMF92lMGqQcGSl9+uUCzeeVkD7lgoZMEHyEiUcbUNPa13c4kI026P8oNwUvn
UJxj3Bsw70R7FPHcBHghaUEakD48wI9MZOfx65/YLw7AfCGWXnLL34lCEMg1zcaP
/fR/KbPyyIDdkBDwT+1iVeEdNevTiMPJ7bEDfxEFxAy0mN7O21/1E83kcKOEs1sK
I4XJj6LtU6+gzstRmBJhe+EfwBnFEL6rsvNA26vI2RsTVe5ZO02CDd9RNsy0PeLP
51Hq7Rs79XzwTeSfBda4dwWuLDzj0h4V9Wr831EO/pdo+q0PWdmG9m2tkGFRIQn2
nxEu1mqLEx1v8vVhy8wk4HWnsSlZANcTTLMIUfWa2Y2/b4JbpKpgeIq0LScA3JO9
QCerS7kAUAhPDhusmOM3pF9S0HSZyB3OHlVAGg9JpGrsQ3CvcPislTsxUn63burC
G5QtEAkIkpqvEBjEiE0sJ1s9vZEyescU+cbCg19SwQ3eDqLjZd/T7JYNIeeYY25N
0BdLK0JddtsvNdrKIwe+n47nAo66nbDoAFhGFatsm0V+gac4jehzCSfBFiKkx+WC
/A1rusIILkkyn1gGYQPbb2aXb7HumFzoCau7Gy2FqCxnDIBhFyOxBKnkvi6+rb8n
8US0m4X/QggjzsDwTuUwCjtuCdyGezepiedM75dQp7oFcGLYqlidfvj8NMePp44T
p/SvdukxHekNSjVGLNd+Zo6lipgw6aIaB1ZyD08R3Evt4w8UTH7BQWhYhlJeI7vB
3noMNcn04eXY3JgNv9wKEp1ToOkX6ozd8JCtMBiwQ97FLKk8JXwf90ku6PtvwfUj
A4Et+n8msbgInckIdenBSkRa71GXWqH5vUPqrNV75m7GY1p69IqVkTgk2CwuJa3J
uQ0rlxzDg8inI4qrkJztqpy8wAIA+3mBVctrKPfvPoy+0KQovTqm4QD/DrpSgETN
Z5ylODHz5WNbZDVFu0oPToB3+eVchmroqYk74q2O63l1qJ0RQZwVfYj2KenxobQs
PG4dRA1DX1vCGhbHrTxnwCh1nnEvnRe9yk6AbDfCa6ArrOO6fPxFc5qmb8ujOlyM
6yVAKGYfdU2szvpzJkKIVjWuqGYBp+sSjrJpRgrZizVr/7YDBMX4Po3uDfQUxzmw
+nRguFCEdJCNFyZxZQ4WZnAu1e34UO6k3MnJrgsKRfJaoyJtEmn7ZmJr5QWoSv0U
ezpm9H5p/+mNfOAGuIiNhqLjUARiXlo5APi/5b1/7qEdeNCGOAFKnrz8rxoXcrqV
OtSY2O0AYnn42YUz2mIqpiYX9Ozr79ofFQxzL3ePE11UCEhUWTUymA1ILiHb5A4x
B2MOX33FAR6pBiNG3pOvLCrdJuPLL73N8QBaR0pVRumrdcBrwMQ0CMqcsqgurguU
vfGWuL1vnjXmnLrRNspvIYiedoX9aL4v8EaQcV5fZEIVWPEuWb7CqAbK0z3rHpzO
NoGLnwy9CVGPC8d9nd0ZMYmwJDKH9apMbTDBy0uESWwGTBQm4pgTELPfOjPDi4eP
QzVw7SC5AQxFUutmAevr+Ypk3oShjFOGpC+2BlKO2TUKwvbn8MOmLIIrFBv7EZHO
D6T+pHaF/ErkFjZTBnf6IRWRPO/RijlGbwe0NT8UMOQ+/DJwZUlKF2fQ4gDHQkdv
vxhR8srrLeFd6MLY29+EbGShcBpdEkCzbsnHVUqbl7xQfEWCpK8oHVt1thRfyOs2
zn4HFy4WVB1fEYiPf2ReILWM28is4SL3ez4WOyhu+BiHbdwjB6Mfb8N/zX+KjpuM
lk6tkADufag5Ftbrbh5Rer0/RQcY+jHkToR8DJC3e9HmTYoYBjU0+ZOglXqgQGAT
sylfaGKLLbUiu6eWEQYSd20a5PqcxDrKVfPa9uJteOUeGcIqmnIWt4wFFH6rNkko
dXtTjfPyL3x9FohsuAXsIUZuyis/jp8UO2dvfIURP9VwezmvTOcz70i0M2C0uqBr
txNMKX4uM6HP8ewUUC8N/r7c8VrmPV2if7eBwXtkx2QH1An2dVNgGjt3YC2vH53T
npEEQgJzrQQjarwfinuYux+hpGDJo9pQ0MEj2Ka5wjy5zwAwZutZkSXcJLyFdTzN
v/9hBhN83cbeJsEGtTMFXNgVODFTVma6jk282d4kxuuyLJ2KyiXK6mBungwNDzkH
YFoWDDeKhucD/ReBCyNzaV9qdXC9m0CtKBXICE75EnNyCKJt+tRuuF/bfdumlfig
IPIRhdFFbpGqPX82bq9uMYYWfrreA7eukQd2mFsPibbWxMPJkQtdEITV3JnmUuuV
EJH1mfYUwtqo/gOsFe/VSwR6J9joOPprwWC2KQLaSTkeurLdCmJT67FiIpAjyE8p
LcnhBbT7DTOnUHO+ZsxMEMts/lVym0ppMikOqVsKyAWwsP7+JHef4MD7WeIe7rWe
eo6YljxyXrN4Ecxoq+5fc6r6naXOhrTl/gEw5jhja7bTOwjElEe+K0LpQWim8Isn
MfUPuZV2kKSxZOO8KGmT31ozPAgPl+DbgxJxWgJfqvFxB6BjJk5tQYjk0UwNS08A
EVedQsWWPCT1VFtALZYduEqgWAgI4bBKgaNg/870RcjWFzwFWnw/+ZbXmEZOnGQ2
QzBdWIRRzii4sz2NLxQO96sx+C1doJpy6JdBXurfzROeVyKF04JHM2/Q9f5aBi6f
lBdKFcLMkZePahRaYd33fVlTnl/xEARRmRV7KKhYZO7DPKzNllrPTvX8RfoivXI5
9JM8nFnAlas7sWsJxmKGTaIXme9VRgOvfRmX5i8xSNtTzp93VBJ31QTKfr+eKoAG
MY/kPQIl+CzyMkYKi6VhcvbnkrnTKvuCUGIEr7j8khVo3unM/UNrRUkBSVOHR/tP
/gAdxQGplDp7cmXuNus7j2tbi9s5OJ0wF0zAC+MF1JWufK50YIUiQmnyaZlTFGRk
VImFkPIktlQXT9FzrmJlTLI5v0V89xD9pf0egS22JdSl2q6WHCslkqAe69ifGku5
CmgWCFaBnb4ejpPPHBYJfAAlniNkEpteIP1aH+hKR5UBuKuVY/xIvWCrRtp4+U4k
ql8dhBKetYoIZyfhpRsJ7lZOV5ecvkPNAVwsz8HQY3yA7dzceRbSmNJwU4QNKsTU
atgU/g1kRZBpkBFFiXB7jfFCGO9x+jjJoe7fpuOBIt5jsG9+taXFtlE4Yot4wD7P
AYuKAXDs+DVc1Ww8FNAGA/cRputoIF+LtMi8ixYjFinFMwLq+w/BRPhWqbSWzoCR
L0MOBDkJ6cwWj14vLX8T/eFLeAr3kxs5Sf6L0e2Z4dwuzubwXYVD0vsasfYmApF6
c0PKrjEM+MkzYm3UdXdVLEm4R3jYf1Rts5/R2lA5w0lq1FFmSQyy8Q8jkNyTE0Be
8VkZTMgBjqowxh4dm+BC82vtzxDxjFO7+Gcye5yebpqjsuJ98UPoaAv+xMdX/dXF
xSl8Wr3OeVAs+wUhFDTV0prObm8WCC9g8uXbU+tivGD43icGaBy/gAyKgEwwCPR+
eTiOwQjbu/d8pfqkKsulVGsO4ixq6c1e3xEQsHVYORt8BLZ3uljFkB3DdRlF18tG
lOdLR9jmJKGHxU1e/BzzEkXaA7Lm/q6O4nguLjI8yKvVWbQlKACe6AWqzNXD7tnh
2WlCdZmrw89hy3VNCDGg5ECY2Pf70RSvv+hhi78DQUYX5E5+qwE80Ukr3oEdDdmv
Vs5AghZw5hxxppn5FWG5pEiOC3hIvDD4vOVHBUjUSmwiLy1rIljRcI2Ymz27gDMr
JhCHCUbGXxZJoMVJUn3xyBWRRYPx9wYehvBwrRADPDynLgWks0N3gzLA1qkylKbl
H1/QqEeaxtCpOI3NlSPs+goMN6VUhbNBlwQMaj1tLQ+chR3x5pH5p78NvgU/n0yj
XoDcMLX4HTffhrWtHA+l1XdfWH6auIlYiFEFOPJHN/U6VIxZh0kuXoRxpSgpbRVA
elzxQG4UNinZQgCeWKoevHr9Iy49AwsxWXMhbl13A74fFSQ/vNkg0+d9MJeMNCVH
XE0Q024YvLKUBKLWaZZSEGGYFG6nanZHFV/02HmDaWVdSb12/edOXwhfXXEXvfm2
yqukLtXcajXCLEvwFBObmsxd2bCGa+v6UAQHTEQGKDwYLokL6CPQ3M/0EKin/B70
KRdh8TwGUxdwCTG3SCNABDY3p/OoV2k9W4UA3bVIPR1XpnbMwp85/rlgN1464flA
CD6tnnfGbkLv2wOHNPlqkWwtfDTmwsssef9WRGb7597A8/fLnuWYCDY7JEmlce1Q
IaKezJ5X3euagjmOY8IRyD02rghXqTcGssvg54IS5bJy5CFBimpGFr/g7AlgWy6i
j8LHC9qBxz8/v+Zo0+Tj5mwRBBy9MpgrF0zf32xqT9UUFZHV2nWlFG5nMMs6Qd0M
2wepHNJ9ti0C3VQjUU6Z9uwc/nyZpuQs6KHGyfLHmH6DOnFw/1UTWStk1O8Ktvka
XEn+H9n9C19EaELokYbJDq9Y14j2wjgQAQ8yjpx4lKpU2fd8tPpaslKmtmyFPT4n
/dNKgM+6KKZiHtySF49uVn//rdA1iEecXmdrae308WA19O9w6uVHM3d/cZx2EYYi
Qul9CiTmJQN8qRRX7qsPEHSI4/sMmxpnZag9IyveROAHas7JmINpFNnOvW6AZQzM
GmQ34XlkIqFVcoGW/3Y0dTDVTP3QNOWfy6FYoZqvdof/ZgOad2MTQyZQpBwibo1u
MJXHiTb3jZ0rNHk6Ifo1MPQOSKWUn5LRZjt8poBT6Ady091yZKJ7FW+moqfW8OHy
HlI3D09LAJ5Ee9R3dXPf/Q5Z6Dtu40Rm6jzUKVnEfQh+5mwEDTJUCcM+e63Zzapv
Vksn7ACdIwhSXKEnE7ELFp8o055/mCTezKLXCtMgTuRUb3tAQHJfq239kXrbMHnD
10AUirvsoTn+VmA8zQrNvSc7bhnHk8kkDuqNrCTYfpaRc2PIj/COB7qFS/ZoT5Sn
yZGB/dUOIdPMeGJ7LX502Q1QoIMSuCFxiI/t4oh2B5OH9NPKJHg3QJuQy1Pb7NLf
XwJguOaqaXpolergqV7wFfgUSpblwXUOGFPDerg2NrZVgyVyVu8HDXH1NtoLd+ia
ZIGKigZ/OcPALbkNWszCcFKfMCk1ALdR41qnTYBCORmOD5u80+Els1iisd4jUoSu
Fey0e7d+xPAE3jkTVcaNHDdEDOET+fqyKYYAL8qN1YRvGRb5PvPzV16CUuw2LBrA
+WhsjVRXcxMWvljIjL1BG5HfDLHCytrArnJUa2LIJxeX+W3ODSzm6BEECpE3v05a
/o47jiHuegc1d9BZdurPpOtXadjAXpWtonEvSMxiL2jG1mhmzqUPuO4pBybkysfu
NpcqUFa2YZZvHE4U/v4ZAYQAmb9gwaaxqNF0dZONFw2bz9qGSbegHVdra2pwC/l5
brh0Pj68k5mahU7v5gD50eufQ2ITU5/+8wrgV0j41aERWROc4G67K1jQSbM6SAGK
7CLLjGtPhLi2aitmyQFvy7HIGtKRIJMjif0pAiN1CLIAWhs3MRPXNSuFt2o2dqx9
/C6ezE2hZAhfpVNInWDjochUbZkrFqotdlHxSsey0GmEyjpR6Tg3BJr6PjobI2m8
KLV64joKku6qeh2L8dMq0slblnt49P6b+t4qe0nU4ZrC03O3u07YkpTSc3UxC94L
AaWxcYzWa8/iHlCIOSriGtDE0j48LRRzS3x0H4HtkW7HGLC6SXZPEVYwiUS8D4yX
UjLcuhjkkKUHe5ZtwciTBLWGvSdmuBOvI6bs0OwO1o+dh4bSMylRUVjLBfO3WOu6
W5qm60auFeU2Ff0MeMlfBl/HbhYYG2AvZdKLk+n/KugqDgJ4IzneE2Fui+4wvWHJ
rNxxsjHjZk/FYldP1SOZXrcrNRVgDwt+FZDIUOul8unKwSXi8xJ7DxguDHTFnhzp
jdcR+87NXgqQCSsmhWoiBfPRC+amc38M230Stj6WChqUXPSnNqGo4GBY6MhsYGKk
/LLtNbtPbIMX7odJzXFcwGMN/5uTYwb3SakJHoFJL0C6PHJucrzJ0Va5jBSO+7E6
Sblil2OpwGNjRfQ2gsdNxsDhEIhn5uMczQHG66B5pOtjHSyTIe1kx4dknLYdhFr2
bY+NJ7/zBi6HYR0N3Cq/z4hEl6OoVDXUYT1ZAucAzseiZoQEQrn37lqO6ehI/gu5
RoeM/oKSJZo70j4sVo3L80WZSWlcXRy3PrAxFaBTg/e+RPOaW0/BtL6NzYXIMerE
EJ5wFVP8jvOWJbUnJ6KplP7cN7O3PfPVhuX69UyC5dwaBXMnO/6vcutVSnrvuAR3
xFYuDN0bHaUPutZvTYg0eQI2Po3K83b8RzrUTtwoFMYOflsep8F7cNvomzpu+2ix
SKwjH4UNwikEJZJKG7NRzSNBbw176bVXLxGkts6mNLhYaMWTZVtx3EJkDR2wTlPC
mTlJys5ECnZRXTz5RMFPUX5wGZua2dY51lMDCPz6I+uoGA3oFacpzq1WVsdKkLBm
6A4NNNel2exTIfP1hNnp+ZWGXQZ3+ND0eIhQGf+Uy2NCabXlBVi+ygNAJN7nASh1
bvU/+nvMtx2RE48ssg70QcB0gxy2D8XEASM4nk7YyMb/9KQlmy7UQdSTg8utE6IX
70VRXls8iPRxW/dmCNPN5fH9LtkcsExc96kfhgs2RWcgt8UswXWOwIsmLXHroVpu
mAAfeymi3AWokjceaFYQqSXGnMZbZE2ieoTxKhIOSWY2iYe2o+iOvzTHMhTd5QcE
ylrGpTP2gp5QDCfsse/BfEwJuMTSvh4JWpEE9RBaAKHtW08DTY9WEEZMYpHPiNNS
1Iy2KA1aY2AXuiwXmbw3WDawqp+iKHmh0L4JwL9aEc2wSlJ3KPF8ddG84qsa+Uf2
c5G13zhXEWssxRPPlWxR4HdjkgfulKZCxRnYHTX8LSnq/vP2lcLJYKVvGjvh7BPt
2t2QZV3GASPuaIQ4m7BCyLt7Z0+NoqtFk09L7mvUaaqDE64ndnpnsbE1Ep3c87Cr
/MPQC9fNuCllduST9Cb4gXwbENmiHqwgCNOflvAEX97ZmGHFlNSVGiGF5vctpsOo
5naitediBq1KDSt686xvb4IfcuLs+2585leWUDqlc7ULPndkYdycxuh0hhag0fAX
kJpW7r74GhkpXDFZFHJWzbZrN3ErLVtKKwlLeCAinQMpQQWlTq+VQtNpZOJLg7nl
/2YFuXW4RFCGX5gc8z3DOOrOQy212AcX4JaR4l3zzoqaXy7ps8qEUXCARintytkn
b0wI900IZB7O3lyHzbVcxMNTIrenbfR3PezEwNcyunyoBAajmjlc1YBQpXkf6KZo
DsMo6KDMPrDgqEWS1/TEemQ2VlDwwBv+DcGuGydxn/t1ff3lZ2cDGi7i9k0PogS+
Zk9anrXGQY/Pr+V9eJg2QJ7wMpjrga0ehlOR4B6LnGu+7bU+bfWluQWuQIqJfHac
7hDK5d5ffrc9vCUEIylTYsO2S8wnGlnM67sU3LtJZl3JrhyW5fj/Phnr4Nl+xFeM
GEj9A0hppaiHgj0nYjHM6/3I2a7pjkOGufKtWufNCFs8+BLwGiuJT6CK0yTH814k
yNg+nAIIDsLDyd52xmFuGWfm48PYmy9FJ9CcvVLn+P3HuTL0Lq2l2cx26jQmocg1
GhbrYCVpT0Yo8UavyZ0WGZ5LZewfrINM8PlHYHLOEBRRnk0LhvmANWGc51JoNDL3
TDJALIOV6Ff2ea+m8rlObAeO26ijljS2LTFyZTjpNSSGRnbU7zZmBZgrRlS7XM4v
50/LL+UCik/VS68JDziN9yLOGjs/qcKbmEO5V7xv5mQEnYUTnuCmLVvzIJ+wgZR1
8qj8Ct91Ue4XVJnsGqvh3x9kucL8lIcTJY7Jg1LFEffgUmgwg7GYtamJOG8Aklyt
cfJYltockGLu2U81wvVEb06hTzSj5PTYz8cWIJJ1JNXQVp9LAsPgt6EwFzgtSBRa
M8gAG/jNZqzKGnu36pINob9t/Iw/5sQ/9UFAf0N3Dj3kd3cub/O7Km1TrDxoqh45
gNhGifpTtM4VV3yBpGdUVUm79GSDWENQCTkFcDV2vysbhZFAIM6jYaoMJJlBOHL3
/6mJsaMBwn0vT8XL5pjY3cdpmYWp1GS+V8nOdKkvh0BXQ4C562gVzOZjM+MDTKgN
gLpeC4rTB6yGfzQETAB011sQ5AXX5r6BClgIsOQBkKZVNBSENrBBWgXQUSl+qbYx
FCXIlfJis6dLbNy8l4VbU6DF4ZfVsi6QP4c/G5+P4BD3G6FZ2F77xDe7Cqakceku
UEkouILzvcRgQFTPJbaMCO6fxJFfg7z5oPM3MMU5lzLgbCJTogNzNh0T6sbEtr3P
4SsnOkN7BOQvFdj2KNMWyvqHwLuvMIuie8+snVHrx9WAbnGypYacw1Cc9oNr/ApC
hrqoXCc5396YNFH/rISoC9w/B9aLHCElnbygIfWhsIkX69D8VtjsKsaOVNmxHELg
2BbTQJTvleEjLaB6mh3wPIYPovPkpYC1VrNlawQ+GCCBX2XRyD/cfsLcCqI+xere
DLFTvHlCQcJrVCHRPWFNJdUXuOI3PUdI+bJRCKD6b48jRe2f4p0U75NhX/F9Tyd9
9s0DkYqOeWzLJUEP+E+p1FIUMvOghb5NF1X6Fl0u1pQwDDUnmDn3iWaBFi7GIPQ+
BlJBfC8O+rsF5Fib6bbc5rQT/8DVtP2Jzym3fi/Hm6/kBsZaxHFiumblpZ3JB0iR
sQ5yJO9PPKw6P+bGZzwjh2sW1qDyU4br8E4e0SqUhZaX2IuR0eoTFAysTUoSKoa/
TUE6ew0BOI2ti/XOf1M74mr+h58oDhjmq+9A4GE/pRpVYcp9nYQoO2IBt4AzzVvs
RQPYVzV5kGvhwEELG+d/LpBltdizxMVcFL9bcoOSRCgFZwI1gsUn51nxacigqJr+
SteFZV7kmQSxbsN77jxWAMz6+RnkOriPePOTll5r7kiq9FqpmBmDlvRlALaedz9l
l1buWGgXHJavozZXpUAkzHZMlpxO1jwQc8jZHZ8cSXfkykKNDCK3Td5LStxZI3gV
DMq24UqO8jbvU7X7NK83dNmpIM0rDyy4p/rPUazkq2iWM484G//ulG4UL41Th+zA
zRddDqQe6q9irY0o8n5A4RtGGU0XYn7SICYAkbGrcnfsxapPwaI7w5yifqH1nyai
dBxtHm+7WnjG9h3aao//V7MZPcAEKSa2Rk3z1vZ0zc1cymEDTHAQlAduXmcHq0bU
szTxDOCVWSXjFjINTQ7FsBA9NxTi2G8alq2Sg5bmuwBYHPSfOpG8j1/6VEWkQ8Ix
8y0Z0K/fGufhkr6rmFZvA+YKXQdRCXU0RjdcyJqwiSOsAlDHFPnt4fEYmJaYhrAO
WAMXHxaxO8+tV8mIS/FHOzxfeRpT+rD6TCvjxxV9GGOgte+FC+xBGFVUT+LcMH7o
aFDEkN9V6R9bkdYxmACQAlfrG1UukOEdaPUdXQlh9xgEOPJbv7od8Zk+ER/QYqJJ
Ep4loCRrwhptvL6fSv/roAUysALw2XIBQUREvSAcbZBpoitc/4D7trWuUeHZmmOC
+10aMyN/HlStAkzgBK6wY1BM2o+/9Q/zTf7W50arr6St433DI2XbgoTV9YCdLIla
VOHbWRqWQUKlYFE6SSpfAVh/nmprYdsh/OzAoozvKtd/lZFHePt7TSVYmubshok+
+0yIhgBv0lAIJ6EsXHGt39jG4GCfM+ChhI576vaaO35CwJOKH21muMYpXC7JwQKM
aR/lwsE08I/fQc9lkvaLIV0h6xdQCnl2vY8haQYsGoPCDmx/qWJDExJK621TDE0r
QsPEqeO70wg5hXiDCGxGyQY7VuKJMzxlcPxTMA023wL5Xe/WKAAEKEpyPklf+tq8
B0L133NpQIT4NFCTTwfOVMof1Ix6LhCeOfjdpxvofBK2Tkp/TfPN2Ad9kjUu13Z/
3RcbPDqc57MzJCusQaaqEVaqnxJGnl4BiYBUQsqY60A898niArmOdef94+zNdOXC
BxYGBya46wPPyvAMEPHDroapvCIOkr7aVoUMJv5tLgDnY2PI/I6WwEkzRNJ6jRcL
MdS1TIxI+NRMycgQn7ie/3LaCoG8VothM/Tjmgrs9jAY7JFZqMweZONuHu6kf/if
pAWCFOIead1XeftBoqqh1fzxGeCQRGkVS22bSxx63gT0727RPHTZ3RrmmD52Ok2q
pk4e3WjTahcoiN4t0BeVqN4p8/mwfJZQliUjAeLdtgb2DviLXvcDt1iZkn4VcTTP
MxK8YSpQTF49soXZJGlmW2HcfQsArbCon5ZtyoSx3NtO8chWhlMYPsexIaTb1G2o
YH/4rlbp8ETaxtxPMGfaBcOQ3pXxLZlGwUPCj0ZUPu8tv4IpfFpqkDG35WlCUqSq
kI45LFBx+0ry2iBZ6Wsvl//Bazuq7fDEg2zzdhU83H3jaimkPKh/T2fbFZLfbkeN
+2EGE4vk99Vs1zAa1dCplbPjv4vdqRdoDJcBCvsWiIfgshw82pNAjvcxGq/fnZPo
OUQvL9YzQQ68K46Se5a2jlqD0DYHax1XpBDnPVJvwPwonuz/jkDD7TKvVMPlb63z
geiKxa/7KngO1PZ2tv/g2NyNlFJKkmGdVMp72Hwwt+wmbI8/TmaJfME56yO/qPXb
7tCwuK4lsa0qrBViNGKQ9GnuQS8WvrNrLQcUAb8g4dgJMRl5F6CHjAfBvCW58VeC
UHN0eHALtC24OlANUJutVlB90oOGWVnMSCjE8D1evku+QlqqBzcBdPt73j0uZqrW
A1P/eJjC5/95ZJBeB7bJQ2eUH+byPznpcXU5TAsgZP9MCNFOsnDWo7zh5jO6yW11
x3AeM4DgQkH9AoEv+yEbu1bTP1m4uW/TfoN0iCT2WrrvEOeHEYeVozreASaBm5ig
/ljBPjfkxLZkgMs8+1rgFvhDEVPB97lD+vY2W+FcAQk49JDKcutuOtIdiFke5zVM
lm36B2OaQJjRiHcW7ntvMvl9STmrbbjt+v069jTDtEFBGf7dCXNMsc2JAwmcBXMd
c673pF28jbKUd5NDifGpAz++uqn7dcv1OMBOfgt8yDsLTmJyIRrCibNFjLYprPjd
KLLQlpQTaCtRIjKR7iXGMevyEn6Q9bo8GwxBE/kn9NDzc9X+NU8im5KofKilR+k6
XWHg8clXN08BZfmj/WEDigjMoDo3aMgaFi5KBw5Sa7ZMjofcpgAs8bXHAPo28G8l
fIv95rTUjL3MIE6z3jwyQiRRd7Lx4tzagUNPQ0MFM3gejlmSdXSaBxgtE7M4GZWx
lHZQ9j2ElQjOs1iKmlvI7jg2gHnBCBfXkI4IU4f7+6aRMA4Brdb32ZjZwS4C+wGC
OTPmivZb6XESvFfkdKvIRcaTo3JFUrSlC4PXlpawhsuudKRyMfe8cWR+SxfHTC/e
WrEZ1Be94HvyJ42KCepGU+5pzZOJ9GVdxTOLh12IFfUmcsh9bBnf41oXRypV8v2j
b4F5MFzqLi/tRAZzFEOvBOR8nh3oCu2u2uGSxqg8QvzAFcGnlo2w3om8TkgYQa4Q
zjJOuk1XevoKeis5MPcvT5z4ujxf6gLiJsYcC/w3utPsgG0S91JkDQZkgg+EgVa7
54+E11OM7OkCGTwu18zNwsdIQ5ePoWsbS/CH0ARGF+afrLnAngZPVoz1gFGa+65F
b0a6zKZT9gFLh6DJhvMiqbtXMnyN5beVxw30pCC17NNP+5e033n5vyaSBMY4G8SF
Xjmiiq0N7GH0cThyeEMiELa53Oeyuaao1A2SMjQIJjXOruwQZtidqXQ38Vv4p/PS
ycMdFgjq35Jk3cF0Wf2CJwtgwyq1zuTH6twUVYatYb7qp/Bn+U8tmFG6DTs8K5tY
ZikChc2QVuWK0zg8vjV4GcGJo2n3cQL4jLOsOFS+HFeLlyZFlyFALnet7VvbEB2l
kNN3UXEp2miBQX23UzxiwR/hkadG4zkMYBcqiXYN88xIskTW7U0LcviDUDSa+E9y
GicsudqjDQ7DEUEfqX5D4wE5XjQchRySSnt+7ldm2Nd2Ue9C1BtqIA22rxq/AxEc
Z5ODnlpb6NwtY3wrSnd5Qlf4swXfHKVX5PoI42Tv5W+wAI+11hGn9YgNtWJdSzhI
DQsP+jBs0bNhlweFJ1vHJzNu4NynwO5xtbWrTAHGKs3ARy/8vNIPS+Gq9CtEPCt0
Ktvvjzvf3zBUYVkbjRxjSMQ+E5r2CkRNFkb+vb1DWQ6qGb203h531S9Y0y5fRgcO
FRs7WZ5RMtCavcZDp01TDpfBqBPu9TGfHfnDbxhD9wBOLiDlMDaippwkOqRAGjA/
L+M5UHDbj6fQpFZO/aWLbUdf/1pt3mN0gjKecrfc4JCFF79pxALX6Adjt/k72ig/
/7hCpkq2j6ijCxOw4D1dlEIzcPxY6f8bxYPh1zeoeNZlCIt9vx1oMZOdSI2RA+KJ
h7I7v8GaOOTc/jW3KpI31emguJH+yGNIgJAy19N89AFje0JQX/NT6LuHzJ7NuhLJ
089yjDD/TCSFoW6ERAd+PRVadJgpyV/lz3jMoaRE4C2kqSzI9laSjfv7k975wMEM
QQ0EVliny8jXK/pVWdQiOF4uX3BBod5HuXVRPDOAnciCpI8r33hJo55FOOh1hTfy
D3Afe7OaYVOF81KmLG2B46D4Xnh808IlOTz3IRjub6HFdvTHZ0WMZ60Tr81OH4Z2
ETpazJ6+o0xbiJh0T5AP30Dssl9B/zYYAd3agFRZ9NQ0puoOUUyFuwCP94Hj9v4I
CZARrXUoxsLVK1ZEWwmUqthTl3w6y9TphiljriPLPJq5lIv+FQdCmHrWDMO9x4CK
m9lj9cDExvm1CQK0puLVA7NsX+ZpSQO/iqw6TiU9cLnBMKwpRSX7p4LY1E+Ut8YG
8P9mF9G77OSNgfRvp9TS9DW7q/5lsmpmiA4XlqrqZJLFIDutg8BoV5fDOzQI5U1t
n/L28sH5L3d5efEuslZUwokwROqKehRD/mAYBuENo3ugt+WDFPd8QA0PHhXPztjZ
S2kXk5qDXDQmdKftP9eL0Aoa1yrIX7OcXJnEIpDFm4zdFx50AWi4Og7to23ngOQf
YJ8jq1YbM/ONQxZCjA7Fm02B18J6lNiIredAHq47KOh/Ft3WmFg6ZOhzp9RaBEP2
sQFeEA4V57MpGjafn1PHLGeovn3M99N52sj3+gTe4lajyoXJepTd3tV5HNVgjCtk
C47Ajjxd3+3WDIZQpXf7d2jURtZ0JDCwls50hx7bbFk9xzkw0mftZu1AH8aoQDiT
ROnRhDn6IwR/S8bPybb4ANJfUFpB2Hjv6r/J/0kP1RjOl/junVvTnK0wXSc/sSL6
M0jdODBv6VacFQVZplwke6V8qLM9iGpt3b1QJLHbkLemSVBQWV0aTgLO0/jgVRvd
Tdz5Q1sOjy8yd0c5s6/C9pbdLeOCxeZrXEZhh+YClZZ2C5Sqkz0kiRxHIeWaYJQS
91o2SkbnlnSf4js1ZqGlblDlv8vhtnoaHA7UQah0gB5nEfwjBDPku64dd1b5yI6R
YeZVy0FW+2OJBY4xr8VdVkXxoj7F1SBTt2SQWEI9vjZ7hT7qCa8i7Zcl+5AVk6WQ
K8WDe3EJRUtPSgpIPpCDV3VZ6xiMGpzFzjvsbhYZ2kOzF17ECo64b9xqUJtqLHqH
Ivrz4HNzzdkBFkS5onB/6SyRuJ58frFtKtDGXVIwBryogigItI9WH0yryKg0+m0h
7MmbRj8F8a+OGuMbsFC5ChOVZmpbwXs6qJQCV5tR96Hj1r75YBQiUi0N0bQkFaYK
W32Mfj/aYDLemL2SqYz2UMGhJlv96fXIHUuB6qMh17ER6llOHSc9x9tQY9Rfd8/Y
vvrW5v5UZpHv6A5OGN9tSbjoHv088/mZU40oKyjiK9IgAeJHbTvVmFgWt+Rl0cyS
3u0d3uwwNQC7FGiSEEng2mKeZDK6PIYzaBQKy+pO8dPqNciQ4OwamwUkOEviQQ23
JQtCF9JsMBZRU3lQsQ/XsKDdbtfW08/P3vbMiAOL3BKnvyDq1fpdJ/IKDNhJE+7k
cWkartdsiDUumBk8Z9I04tOPBCFIP0uU7vUgMQQPBYq0JkHdCgLvDs3TmvDlU4Gs
jUAB7I/vke4EoyEriBZGryPj89DdqFqLI20cqzuozcecYvPzz1jj6uboEE3NVDd5
WlqVKi6BApteE+EYiDGXmqbTDTUV68iL67kwU8+xG5m+AdNDaqSMeJbQrmuRNj/o
y1kvTPGdulE+Wn/IM2BHENmDbD5hh6onpRYGYpQBmN6s9I3xdFT2VsaxX2UTJxVJ
HWynA3YwbKF7Cj9FISKsLi74z5f9/12Fd3gokmlxVPWqe/PewveuKxjGj7Y9HFGM
AG2j5D9G17aNrIx5jnAUoWDBu3ohI4ZYBsZZOytKbwBs/fJ/BM8jHCtg0gVt4AUI
fWD0j1jpeaaZcu/blyWWU3smtIK7hGBytOrKQ9eoDNY+scrHft5v9nZMVd+dCJio
qAfivYzvSodZnSRo49qBadKKfaAF149R05asUUZurd+HN8iWR7TtMGmLNmtPBvv5
7QY0GpZ7s0ACe21Ph2DWBSxS6cu9AP2+UhVRvVVsTF/izc5epvQqJow7ZYpM8jBE
MA7BnaoJESjhpLI3Zd3G0lfNT/xJOshFqaTIvip99gXk0aeDr4TSRaa6Yov5xq7u
BgRrRj2332TeRXfM7T5iT1pID7N6jjBK/eoPeB4hAmxQ7U/4kerzQXYQJMrsPo29
neRV5jPNPeGPbGPJpL1s0jfPeL1cNTteEKo7V4WbuYym+3OT2Xe1YfMSnuRthOQx
PJob7aVsXI9VFfGUoq5guLyt5XovESnkcPT+7L95nUgi3gX3b4Z/Cz23apETbHUt
8Q0BBFSk6uzMGxzpbRammUJxIGg4Q7OInZQbn08RMsO4K/4PU553woUToznStYIS
IsMa7+AHB67ok+V2tLOwHypFOihRgK1y5HLIW2cMyrM1I9AQ+OviumnDP04FQySN
rnH5SK5ZX37pNxnbETHkbMypbmHWvOrhVf0tU9cpZTAJvW6c8YGhtK1QrQjH+yVQ
SzEMhJVMc5zCBWoyxBw6MfAM63x2dKsBLe9kpE6g8r7Uol9EY1JP2vsMnxn383VM
7qBEgQS0gxTgDIUPO3OmtlSz34mg9ciW3rW3+DeZK05U7oRIERYTIPZ02zHdhqF7
+b+OiValucX4eIF7d6/l717rZLoSDmJga8ovZStKpaxKrZsmIz0uIUg+HmYUuciP
oMwZL8TTzfNh7SAZrTBtBjBwqtOmOdaPHvw5PLHywP4ef3Nj4uQhE7YhJbLh2Z5V
IF6BiI6VJhFcH4UIb/IxAFyEnM0wft+zKD08Gn3TxCiFsYH0poiRIY7jrVvn5zPv
GTpihTXY23dYtqWfMuDrsPUx0QihnrrPDSjClB4f9tWLm0/1Wcje9EhzAYOgW0O1
SSffflPAeOIkhIt+WprudrPguJ01uZvbHo1zdWwe88RYSdw4v9xfvFhYVOMatFYK
vXEMj/RswXT+TtQtH3Xb/Sgowjl9sqcHttjglWxmpE5vZwa0rywrx36mhdQYloSH
c0Yy4UGREVFciJlXEgb0ZykIdnSjLumis5kkfo4qYUelqsYsnlz/CX0s6x4LNNl2
+w3ul7EulhttsFtdgiKQ9K5pRM2oNRvnPO+j8z1NUyQjk9OQVwHuK65aWce9RlcL
DTccN1j+8pLascIlgMdtcsDbmv2q8QctqvoYm3iIBf4R7Mci5affE7OMCEJzGMMB
GMKq6HABpcjxivu8jzUu6CJll5ohL+L/ZfP3FIv+lRVvM2xQlbhj9jys38pXjOMq
mw4E8nytrSzt2yy5Bpwurl5T5HGKx6xDXUTuu+wUroZxPfujcXrDtnwyyhJ+0KcM
cctZrQB083oXAOjeOsbsc4wcYnAcxYFOwRfrQDbtX5H9oWLzLvSZpANJ0Ws3v+d7
gjc028IX+gmEzFhEqlBSvj4Tz3O14a6ZjzMU6zWigD6VF3lz4ET4wSZ7n6lrJVM0
OQLvR89cf3WU5loFv1pYwDg8DmETXXMFE+B73YFV6FQE0Ju5oPTZ0h2xsMcdf8Vt
Enbx0+4wqFUFzI5h5s+OPiQ5vgr6/ohjK9++yG0Q4VA6l2cwDsXgguhQZEYx4qwH
OyYjnL7qPNFiCK8kVK6GdKVb2Q0J2KbysvtONj0ZYKmed0jwFpbYHjPSgWMtlYu4
p+j8Vo/8K++BtvN50+8SSSH6+0GoX4k4yFRorg1TPzLko+mdYqtarND3t1tRsjdx
gi1As4GVBoNVjeekWZ71Mx1I409ozTXPMfvKhauEYNEcCpjqJYAUdE9Ira0wCvtI
aSiTQPOAkEwRObws/z5DV61M/wpEqeoJwJ7mN5ZgyYZs/iFcDTOdsoL5ST6Por3q
uRch+ZJLL89Fa/dh//3RU2MM3KbDDearhIMBb/f/hT3HVI3+mvnZADZZJ58RjwGF
RVMiFhDX7VhKkx/H1jR09zdpwdl8QcnSGdWEmUWhApS8ix4NQ673FUkkU1KXHV3p
dPevbqPjC9avevEZ2NntHuIzSnPNAcJ5nocGSq/LVoFnKKO+QTBJKDhEtHMBrimk
iW12ftVKQ5twNQOYn+WebwD24hAHo8vFjuOR0I2CO2PdfLHqmNO0WfUxYoYTNF7C
iGL2Z6HeqRlL/ve7zs9+M/qJZ2jnGOLDFLMhxwjUb0kIw4wndDIyZJXAWM1x+tn9
DNlmff808oP5xP6QLhxGTVB881RxqGbrQjreqzYfKuBED5AivG7sS0AV3m8HgPoI
kK+ZCYPAumZVDJlUxVzwSh4oK5Bprp8ShublgjU4NbRMIqltSp+EduAxK9sfWW+l
F49AuYbO7Zyr0xA/kba+saIyi4fsWmGOBIpyzyAm/rS+kHDTH6x6VeIxpkqCgVMo
jxx+XTzny06vXeKMe58PulR1loyIDchi+zvKCZZcnKWYr4RXfnzM6a92iXqY1FyD
oAab+Uz/uJvILGe2O6lW5Vr331GQzRrekXEQHvfsKZYk+0n9nHr63i6p3Tnc8pdQ
Xwrbkdq/AKMy60gL1yMKVM8sIDiPKJBhczSqkXXB8ZVk2eFEf3rsmUPGXGw+6EXi
xP6/NYyiFoEjBMfyfAnenmaoiOc7SxzvGsUkCbObi/zovyxGXQ/a1FGV43gKCwby
9zgYRxh/aWRErAGKKzLcdJh0sYc0qw51I/+BRYTZWjDjRWh5goqnHxr7TIzg6g9M
o+kb0yRz3bMfMMgTMlHJBJmJlti+QV45Yjk4+/+oHFl3Zb2IdS+TAxJU1rlABwaf
tJEZVkGVKilSyL7J9Fg7L7SeHth2Jmz1LCOa1KFM46GwHr1RsonMo4E+8xrV2zTI
+5YP+NSdgiNSq1rjya2XHF1E3Jzr0Ncxajvf5/qJ+/GtymzeoJxc/o35V275o/4s
7eco7lZxfKvzs/kelV54Ug/n+d6kshzEMN+hRL8UNn8xAVqwReqKX+gtnpEv16Kz
JlvY8YxeLJDBJCpTZoZFhuJF2X2OtA0kuozLuuqwyX0VgjBUuqWAl/MfnttXsGCE
tE2f2NAUBTEHvrupRLfr+P0VMLOdbRJZ15zfndcoL5hj61MM8svbgcC1+5PK6eee
I7ZV/FwnEC9ewnm/3nmgy78BHO3ZeMyMDqgrheuAxcc7+GYFGGUeqm6V8Qb7uZ1i
ko8pmHOGbuiFaDSaJsUeDD1F41/ePl8bW+dUGq3cuRd/NFiTDnAiAxasmbUJE8Tk
xWisJ7rY1vxMiyEdwurpsq5Vc+8MpEf1v98erK0jVKJlW6CPFSP1Abjv6kLm1t9O
+r0SaCb2lsgHTIyafFLZm7ztN8jXeLcYNgK1Z8iWTmGYcgFYEKg2WqepEicDiXC2
3BGPqJRTSrLys8ooFHrKtp8JcIt6ROLrce7SdHoG1R4jplxSGKOyRMotWFwJX6FD
NYmHc5r4Z8YSvzZUiKCnLzI5RaH3cwTu7E69IIstDRAjiuC2/DK/acWncNUXxJfD
DxmkAeDoqXsdICZKH0/I81nosqhnFsk8Yj+e3OPSbloe6qfkDUHf2/98RDYXIUjh
kGmLNIX3SvVFbyQCoQ9xnMPgc+TkblQf+D+uZtjbaqiSB+x4IOIF+k5vlh39keQl
5ZHV0kqA4Pe1SXvXgTeM76RK08srzBbwkZgvrlOw/egUrIMlC/ER2stGxVSrsa//
11wH44vG0cqOgtoVAUZruNntM5xAG83Qp1qNmZDJ0nbhGgCUg+qCg9WOanFirg1Y
3TBV6SnqjUND9++Q9mOXtzCq2hY6VaZIBxBY8AQ57nW85NdtnRUvg2lzmQ3noH+9
ivENJBsSp9YaVahLR5pTiS1HYZgxY4KTLLprW6rFaE5ssG9h3xBRgBc9NZ6kQ600
Zv7m4l5XQ0aaCAIAb/g7KdxOGACh9u7fAx+4TjtgZR3mIsFkpydARkQmvGKIJJYx
N+ZiVpANvj8pWDqCNy15Vl776PSp27ty2U0e7/CfEcrsmC20dlOv/QFLIW+PH80/
PMBe/b1e4r0mBgnGaSsx5RWuM7qXgdGFJz6E8+F5yEW/l5G7+nYQd5OOzBC9GCr5
OAGEentXJxIwmZNxCHC7t8i9UgzNmSiXrRHFx+nF7T4wY24zAheQNuLPr9BuLuH/
hahVmrXrOh9WFmvdyyvIB4QtzwwMX/zActRVSP6102y7xGrjaI3+Ztyr8ZbsB0xp
x7jrQJkCDZVzS1Ax7/YCoccd9Y8jKqFPjkdSalOZwXawfODuySDMEYGfSDz/l7W3
RSeNZalLnSJ8mEEkATQuqOwNx2IKrPQD3CyzafJywxROFA+CSOWQcIXCxU14EdF3
PfMxkiI5SYzB/JfyEoKqbDZi+G2IFok2/wGFCV4GXmdr+j3JqLnn//z3QMdtJ0rn
A2CDShlWsxToIIe4pGN6xH3hXKrg7P7k0n2JPo+7c97OMxXDxodNTa5GNT792T8X
9qraCQv/N87glbkd2iH6lsPeAUUI+noe2PCZzoXCHoTNk7zH8A627RfLWMLUslnh
ykqFnUHb99DYNb8w1z//BlQBMYNetwPbxWa9lE0GBYUmUmAxsGWGZcH8L85p3DE2
/eKH35Afq/lnLbePLHisf+KyALGAfuD1v6tJjBmED/tZq5g5VJvNfjpFUwsN7rfr
9GzfdhsWUIz3pkaQEolQGVQjEt+2frCyAJS1sA722U+u+DMTyOEK1uNpjqZdAUOA
+Ornw9LzoEUrzi5xt/oGJKasfDrgqS1PT6mZ2jRug+H+vBleB/Ogv4xDViW9ua3A
YuVgBYSWCDJDfZOJZtZCsCbf0qtE2c210sIlFi6H6md4HO947aWMyPHzW6JlymNh
04Jy205R1aAeF8Ly6Vmxt/IRR8BR4JPe0NEM0+CvUqoTHak8PZ6TkcrdJZzlCHVF
UHozQu8j92V2IvjjjFMr/J4TQ/LrtYnYoCVie6S4UFuHXt15LXaud+RW/vND1Sf/
WyjWHKMGF5Hc9xZnMRGOeN8NQlseStPzFNAB1Zr+d0lfmOEp8gdYmcCAZuq/ZMGg
tag9LNe2zf3cH4B/nXS6jaH/m9X+OMGzL2u8PJcopiV1acmY9tlvW/zAmp3ckFiK
L3uqdUdIZI6KxoCHYF2OcQa1UjR/xJrwHWUjPe6J8fpNxsrNIYUxtj+yurlIEphS
e8Q69Q3UOt/H+pEPGUGiie6Nnj8YspwaiDTF8QXh+973RHZndGheD6OfVQnv3VEU
MTY3wc7hJSDTJ5AouhDZdhU8ianqrQ/Pnph6jind7E5BgMlHBhOd+e0YTZCHCQRV
Z5jZty40t2Gvmhezw62P7osggROp9XCkXlTprBUfKqa4wPvvahw6m4UlVnP0lXeV
KGa07ZKulj4zpzaKo/QvaKmNsutEOR+ChzMC5APIzotgL7hfPWuxFlU4pgnpe8d5
H1iYtnC+ypYfkV7GB4EBtMGTWffHdKWiGkvrNZarv62TtQ8Ob2V1kBcrD97ZZQFy
KcwMhmfmzi3COfuPQo/TLHxCUJAKDAWw7n96e0CAR19edc1yzRIbv21VXz8EN00T
aASoFDwlxVBhpwZe9OnwuPC70I7rrir4teraJ86onzSpzaSAJ7y/ftS/R5RDoyU3
duvTJ7z3bjDmhOxHqjEJWnWrPfY9t/cm1G8Ilsp8VW0cG1pC9iRnbR8VD52SJBku
f1aIl7lrdOnPXIiJLlEsW4QiIhvLxKb45sxn4he7X0BLG4cUkDLxCKT2ecMll95Y
CgXG1wSNBeeAGyOtpkaAnBssXpJSrPf/ay20I4F6H9I7PVd1QoymW0vOnhf4Zv3L
Vk+2jvCbg4/d+2+AK+1ZSX1H+vlWHGaJWNH2ahjFZ/16mdLG8UxHNjHGI7ArqWc8
RwXgZGmuBOrrn4o/xU5+ru0r5CegomzqCucFdz/sX+8v2HXVgb4onc4PMjLD13Ry
t7E6QtbjMrD1LRwEwbuZ1RyUyA+1YcShDNgjCypL59ago+R2ExDEvloh4o0Q/6zD
Wk+KFyRpJA/PQN10bQTT775czS0kHVvlLBAXr+wctoVMbh/NS9D/HKPUV/txkujU
jSx6WKeW53OJjoZK/VaL8ne6Jyok2zObQzYNjPwoWv6OC/8UAvx0fvUVYZ9tkGyy
4IKV9mpfqvj4NFq1DLTFyCCh6f1K5ntr0gy+tlBONO1lq4U0Tt1F2VuKi7aGem9o
RGJ4raFn29fjKjqNMo0zGJaUTnV685GHBZIP/yScBZRaJSzpcdVyAmu1L2FT9K21
0hPC9chjSS7nIRSftlhCzLjg8Aa5XJyq5JpxXaLRnpghiz98RpvuTSPzzvpRNTWy
M5r3hjaoeVJOt+yi8V6JUx5Ncp/EPhP0bto+B9cONO3IiVJazvLuAt5YhWzjVirz
bNqzLEVRWhCjWyy/WZh36ZUYhEgZwbzWvMIClouTdQKa3hJ8kjQ5dSXQRxQvDM9+
sUJGy2b9mq0YoA3uUhTtXUvMNLLMckD0S8Yewn8ybaytGr6RQyNqJMcN4gSkoifF
oeVspmjZ7II4/vuSRoPGa2JR1W2vFh3j6rjNRe0Uch0BkD4AL0aUxb5JV+y4nOzv
xXMtw1rlBBFlXskJRE/iQnjwRLTI73wRZHuj2Pt/R9fs8A/Kl3OwgCgz001SwAMT
bpge7hSIOpMIZcSWVwoSIFObnEK5Ea1DtH1uHnBbwWetKbMGkJ4QPRZHUhxfvAqB
7Vi2JbdH81S+UvMyYCVvDjYLfh9bS1D640k4L13m/0qpfRZQpbbIE92NFpd4Fy9a
i3coMiWWDdZrBz7+U6DMJz+p3tAcc0XpnVXL1pr6f+PhQPwJ2uyFV6Q/j79L3s+9
cBoWp9JdIbnMaVmguvzKF3TZceW3hWvIBBzHYH9u40+C/ipE5RCE6DH7lpN3NSNR
B8zXhxj9Z7grclkI7MFTSz3S5Z+pqa55CrMQlMHyj20YpRNpmyiP6PG5SqN2zAOB
Hb3atryv2JRA7KGQOrpuAWkcdNe0P5G0s2XuhpGGV1yPgBkrfTqNp7UJx+YMfugl
SLlDhzfUptg6dmBbVx2bBH04prvSOOdrea5w/TJrr7BPvFFz7Sg51VBjxM1Vmj3+
P7IAalx0s7iKTbW8120su9Ib58FzWA5/pZza+qliPYwkxXGcKywjyznd9/uPsSOu
bknrm+ZfHR2N3ninvAKHhaODp75t7juQlE6bn3Jym2JldfEcGJsPWodVU51ohZVC
cbCe5/zO5tMknQVIn9a+Jfl9waRKcuGc9sKvj65txVNfDyl9WzGGR94TvHGruKCU
pJalyiwfKpXakoPRJhfRf9/IBQLydiNr88GspX8DlbPUCMorWeZm4ljfWLcJO9lY
wZCgGWvSDou90gsdSomLXT122ER89x5g3SyFmyOK1Edyw9WcrEsHWtCwsJ7uPojy
m04tJ9sbfKYIAhJLD87vNRQOXxxkoHT4kbxNPHOOlJb9uy0emvCLUP2biiQk3qLd
O7mrJ0DcFiE8u37Rr090k98KErFNXrrraF4QcugwRJ9eYP6Tn1PFQYIAQUFALHxH
Oh1oTYqPaVserXLduwK7QpjuyDxKmNphtLd6ITBGkqovV51QnMLeq/Rkksdi4h5A
iyxK+ZL6enyfdSad1IXKpafigcePZw4uPyvaEuV3UwE2SzjdGEUj5vQeqoIqHRe1
+6TeAobpqfiKIXT/GLs7SRlpBFuqjnmd44iB231bYc5pDGyoJZg42HeKb8fJ1a39
7y7Mfh1TrCfdBC5Qg71xJ7ditFPcOF4zfFQeSgFPgHGijRG3hnuqhVKnZNI5vjEG
/C/RvHwkDQujjhCf3JHNAYDPfT7GNXpH53Mt3JB6Os3l/n5nyeht6+QMGYifpkhu
6TkC18CaLCEDYk6Jsjkqr5NuE6ucSWBUaZyEclbi3syagodkxTuL/fJ06v829cxo
CFylJmpaOCII3acn1Dc7jYuxKG/NgtjAs273Cul4sZDRbxbqmcmBaivPoNOCCRPj
hRbWVP8v7+ykXDpf3Zk12YysYV9ybU6QOH2VzIbfHc57sQxYo8OYoQTqHQYcA/YA
lWyA5xQDfJY1bpxqNQq29Fnc+gNPk0kPOaih+PpUCLwl5JGeH5j5YdXS+t69LWN7
WoL62/jVla9vQtMhCJnfoy7cPFCIJffYqcuLh2au2YfvleUhUUCQTmcaTjA/iE5K
SxioT3oJrgqMekeRv6k1HEcyFOb1ThD8nY6Lpg7UMcjENq7rnmaQv3LxSqgp3b5Q
GfMAoWmvh4kk2fEmwkFT5eWo+JAA51GLWDQlkxitrOJO8hUKKUsHomYYLkPUPamK
5ShgdCqR80Z4RIzDZvO9gHXQ3Cpg+DsGzZYo3kJyUvdhbs/Ep98FCx+IYFCp9LUT
xT4AOPh1m8kAcH39u6nclTtVc32yr1wsgN6pNItTLUhSYlIVKL0osWP2QeTLI1+R
hKnK3tlRRJzVAcuHk6XtXaUj4rAWO4KR3i+9nfZCfZCwKRyfuP1f09I974IrlbXW
uG8UA3ycud47aFaDIh79f7IckLlqXSlRJ3/8HBkQgnBMBHzzW5ASamYEgjHEomsk
6lSn1mGYFwUU/Vz5RQtGMtEQZjvbNRzYH8rHuBkohAexpHEMm5Bg6EHQKLlBHK+r
LoPttvMI+0u34UtTLvTJl95MDILw128zyOGtqBH1C5ZX/FS2oQofxqiSsmLxgjJK
x9U6j2ah9uo7ED5CM+B29pFU++qly3GRmUK4M6GAAFuIX4BDloQu6THtnOMJNnvg
F9oNUDVGve2yYp7C3h1cxjpOpU+TSyxWZRgwSa84P5/CJh9ODKVBwRx8w/voWh0E
QP2HnDBHjXOX1K9pzeAyojwdY4cBaawSpR+6+rVxy+YokyAXAlhuJrXsMU8QTK/N
gOruy9G0DnUiBMV2mZEvo9+3gM+UoPoo7eKsT9rp53UdUrPim1bTEMrfMlj3pLda
ZL3fz0E0I7kyQkg3MtnSAv3FKt5CWcCArE4IQXkC0hBd3IU6sRxB/9GUkBXzJXvh
Ft0+FjV8zMknc6EB+GkR/KouSQtU37qxyiwBX95ZRgOMHMN0rWtUSvNT5ks1iMXi
m5LRcXPevbE0ki6y4ic/kl04CPespwIkBsP9dFdZMJ7rjQid50PMxQh9YL8C/bIY
zHRncBwLTBmWqBSvHlS2/VkrdyAi+ku2PijxycY6ohGYx1FElAITnZGEoSe4/v27
uF8ow9EQBrH9cHtKQZK+GFBzCa+SJvvjW+OQ/tCqfVZcaOHWOIo01y+QiC2EzjxB
IVXdJ3X4QXxjHgdv+ql5iUdj8CApxQq6BLwpES0pw0KUwytup2OVn3bHBweFmJYo
7o64AJ0EfaZaHiFXwxzXmIWjI+pgDBJOSWLYnzmwa9skLsw9QE8GXBm3QKG3qoG0
2YFP+tK2mk3gJX2p2sS33Zi0aCl0EB6uCz9PU5CoGl3esftMjQDzgRxubw3MhhvI
KysBJa6QJ4t6iEJXDuLal7SUvZQ31iceAOBkhszfR0x0dLDk+h0TnoYNde/4Ofxc
HbQR3AgnQFHowsJLDWgQhujGS/ESne7XjssqOmFezQrM8v6YYpXewfQPjAVcWR0Y
YMAysMaBK/AlTRiF6aiIcmKXBNBMHbCJ54R+imQCRgcnLF09WvHxGoP0KSyBtLNr
XbQ8VWgyZQhRXD1wPQ2PIS3Bg2EwM4UBuQbVUaapKW8xkXJ0f1Pm6kBOhxACAecs
ob4ThaLGk4zDJN0aO9Oq3Nj90M0j/Z88aXRzKQljT/XsPskFBItGiweCUJl80IZG
oBFp28YYnFNf9d8VXorTJiy0EZifpQuRoUXXF6teca/RZUd2nszopadSgZ4qkJgw
UFzAt/554F+U3LyxTmqlaIJzLMF3DJEmfkXd2VvU7bkuETZP76fQ3O2GP/HDyxig
/k2t5fEg0/UMbo6CjpZhitNgZhpOZL8dsWKmUFrcnyOFOXUjI8+Yt3bVV4ZCWs8O
B0JdByc2Zp68l1wc8g/wWHVAzOleQcV93owAJc7zhBkqDJtVbvyzT44kZpOYoUCQ
3rjbHw8qbWbBs2OHdy/Qjc1FsEYdGPQULmThzBPeB3RJoHGQppMbwlXRXkvWr8BZ
hBbWm/EFeMPaeiLl0syjRLevjj7FtxfhvaKYmmaVHfZ/MpCjubXxUZwpBRjfJTrI
VL1WAi5Fgz3HlVERco9NaNH7HIL4h6s7M9MXj1tBJ+PP75jinyGuOv1W1WXM+yhp
LeKHc87aUmpjnTgOyn8FiejJzHD1tuRQljh3ts/Q4WzO7cceqAR64gsU5yR/5Ds/
LZGlDTP/QWPJSzOEtW+6o9M+4mqX1HMTvSLGS9loIzWlkNaI7mVoRTNF9tLjCoHc
qpG+RyqQgb7TDOmenau20S646hT2GXlwY2xJ3G3JkX9MuSmcLGipTm19YVw+3KGo
2Ma5rkXHNhVJ3NzCvKHmxghc8fZUU7zqiuyYuwk3HkvQknq8/no6k7RK6vC+Xm6m
OPWZEMpNb9NsAfHbmmQLbuLPrPtVcEDyjtd4/ALbaOjITmorE+od7+nWzhfqZPsC
1+tCsyu78+9DpW9XG51EJ52iJv2g8GbmI/eNj6an6vzydnyBYHJeB6TFoIOY9NWL
caXjhU8D5Td8xN7z5nQfmlo/40vjVRvHp7LQl0UyvsGEuHmbb0TzoqFpd6NTIP5S
R7/ECzAPvTIhbXxbSJKhiBDxn9RW6PyCs4Nr3y8/xdrTwVAX5a7y214JkqtTla7W
7oxO4Q2UQOs0ZHP59C267DO9MuLQH+FFam6L3uNyBZV/0N9yO/6yppeuBrg7uLtv
ailyzGK+hG8lIaJZsPTWWSHS3sY9ong+4/UuV+xvPLD0Up9lmdHf1Zg8UHDDEnpj
0cTj7M3dxqzO7x1P0ZMjCxgcH52XpPfnclxCi/MXUKUOZqttQcUQ/C/CUq0iHl/k
LqJnZYIDTwg8HT4tPS6fIdmgwtZLt75xUZiTjOr3Z6QVb5/SJdPOMYGVzGgpcgn2
v3+fUpt+gMEFVI23ExjMRZAsNGfxCjWtXLdQBb/yY72cNzaxnWD/abZt4opBWLja
dFQOwFFuVnhLWRA6YJylOw/gWbim6nR5wEhXXXc/ui9DcvbQx9m4MR+SBAUR9hMQ
NHmzY6VvXcAeAIAFExrqcieIxffnTiT2YGl34a6iudRKk6WE9QddbduZfo36Ifvk
OB1MOt47ytNCza/63OF+J6Z/uFYa99dYTTrA48+HjGW6zFCvGyZ13WtOvcTomNcv
M1M5c5QqFF3wrwaBciFHBwXwMQVNLo98uR996lZr+DMiwCtVbtoH/UsPC+EZRGUW
iRImljYHiRNzHe9Vbj7R51/6P5VFQ9beRWDhtxO6GAd+b+q+F2ReGWMbTZkMh3w9
b73Rw71xBOWM6o/jl5c2GURMY+Z53Qx9pjtweZfbKOZkyS6ugOZ3VcSM9OhP2EXi
MSnv/gVuYTmlj9YlriZdclNV5sUpha1zPV42IcV6cpRDscDLjBdNpVpXlsrgfG41
KXROaYCNScnvUspsCBUlFG+0KhB9WnXmIUQRFMsn2cjQ0P/VbrpV1C8vDYLU4vax
5LMEM/Ko64OZbce61xpY2OvHkoRB4YlqBCX1K9kwsBTupB+Ykv0m64B4C91rHoze
WE+RMpk61lzHVfSMgrUUxpvakUqYUIBarRKWGq5xFql8VDFfCZO65eAO75WlBG7J
Kh5HenTh3W1jOyJ+TGF6vgV6sMChsYaj8CRJ4QI+ewDVcQJ+DFHy5FHvbEhwpyge
8gd6T2T4PIYYsCMHrVmyiZCclOHMgYzbUYLEeqAFNMYRRSxz4usuTvxUfQAKhSun
RVl5UQBqqNzQP0TCgASvQdsAEV7GeVCYWQHxTMLa02kboESsaQu2jEpcoCYNVyc2
WgNoFgbmpQLpldcUsRcabtA44RjM1OAHYToKMW21yz2tSxsiZSskCsHEsuN18SJ+
97xvE1wENYQOHOE29zFQCNdgW4eTU4GePjidCVJCfBPkzaJhPcldGIaMRCCR4Dep
i9IjkOdq9Ka0vQKtFZXVMOw/QBgKSJ3wjlQuEViFFl2Rhm3gZcC28ZVF7CehwxSP
XD7kphhMTHBxK1Gby7HobqKvrlQ6hk2Wl8XVDEINufmZ5weo++32VxRNI4NkSua3
hVTTnAj6glMEWLVZ5+kwBRUMVxeP3zlrlCK0lVeG4ou4xWnT6oHs6Eo3U9vexdAg
iZSsuXQ/rXh4SGEcSAI+xzy/ZVv1Jx2cSTq+3NR2SlXP8OSnAxpyV6OcmQp9OjoT
F5GIBBMhPVoeQXr/lBYfJ932LapyZ7od83fBqxoDSowJZw7RgYzVaCn/N97GcfOy
9FQBvUBfJf6k4YsI/yHLsDlfNFf7xUuD7sbarnCZCeKW6cwkiIzp/BFDCDoNWo1K
HqkE5RfAqQqQapLhcRenIUzzlUJwV1ITiwwe7zeIK82oTCMryh8A5W3MvKGEXKeA
2ynaYssjPWA5NIQ0cQqswqbK1U0ujklkzXTklDkuK4TjYPLeYItgNkRH6Xv1BSNF
M+ulcTyt+3q+8YwV7WFllgHTQ1Y0ffAS4+AlFtc/FWTorPs0PpQbifUoK8oDe59K
AITuohB32POr8ygZFEAp360OeFESsDaIY8kwkx+VUhBYI1Q1/i1LtMgFKYy0KJIP
oLnuS5MrU0vJQCLhIg2Rv5UyWrlFUwJlLHIHdZWDi1ZL3zI1gBRVSwjbhv0lTjyq
LtqUrJCIMLDlKix6ChWObou27KXJvvp6fZ+kq/geE3yGTD5LwXPZ9+d0gYnP/HXK
ZIpJ7XKW835EISaXCJze200000GN4SGwLeU6Shcjc/FIes5fEx3209obbox8xrGH
K0M+97OdAUZj9IcPOHai2JaHbWKpNDG15dncuwWzthE64UVOqIJohwsI7skQrYq2
/8ywwFQaYH5t2mHocWO1OhuGeypuH1YJ5dS5jCGgQs4SDgGqDU+Dcfm/wnfxJvNl
SpkDyUJx8VJMGDp1AM1foXIkWpYTTuysi9GJiqWwlA2WuHu61gmo8D1SPLmS591G
YspgqeGsWWyHIRbMKzYdhxQKskhK7PhkV0tCK/AKgcqrXtd1yPUs8twdIc3MfBpF
sMfZceshsw4MBJYgP59p55PTals9rSNsun5dXsEcXqcaG9GlWu99zL5H5FIIfebD
6k4SVM/nyN2VBtZuyH+3i55NPZ7zo+kxNmZXmWk6qMXHSz1yYVorn8DGNpcHtRbM
xwxnnW7a+zUxG39xnd9JvMlIEwQOVERfHQEZv7dXNLZLFH4RX4ltHIg2yeqSXsWT
M+1X/DHhjrIuSFxJQXaWuHNML9gJ07w5r5NgqHgmrOCeDhs9w2AH+HzSS7kSH/v7
GnJAtOwgPbnxX/zUs4h+AzjKVMZUwwBUgFvr8EVn+4RWTNmX9K47EGvBTOwMOixK
T27vHOALxM3qyEu6H6sdFwc8O/8/8RhzH+abK49YKViS8L/Z/1rsZJ9axda6Lbmj
k09W9RThx0HyYNeQ+avyy6+t5JSuMqVZ7RI0ly1+8gvVIpTSBveI/D73/o+8qN7h
yF54h9uy16ckuivlMLSH1VgETXxTHDSyr1TzJCuiaB+DhX63jM8FAMSG/QcwkqEW
FyeQl+0uYHvAmkl/YLmTWxnWQ0ckgw8SXUGlQ+5cOHtBLCGYU+jhE7RMDd+jujWf
5ykESi0FLC0SlFCGwVy9ocCJjeVCif27Lyj8htLXuawXq2MAfXLJTfhIeL+8B4B4
itIuJPjBCdsFqGwyoqNmGZyLg0Pk7qHyiVAMOf2xGchAYow+jt0fDh+Ds6JUOhEf
PlecMgYHnE4J8289oUMzlaYjV25qRHOF69bXFNTfQDfImihX/UARp5sh/7o/y+0X
QA5Lp3uiU3s5YY2Q8h5Ru3R2D5b04LsrfNFSm61GFfewMPXoHapoBpcZ1lJWThfb
2wKRu8xpMksDyzx3Df0cycj2uC885LPHH6Cbtjrvlw5UCvRrMztTLrUZnx4yxYgt
gnWkoyvKyz1J8VczYb0t/WmskVTWsjKdl0mboJIVzLitoumwjphTlyUCHkEVqIQb
KJFNzu8sRIhnMenzziTMXlbHSqDsoMnliRiQ/vxt1T95ILSEtnrpucYvzUnPnZ9h
p5Taz3vh8jeUtRnbTt38wYraFvs3lpfEQzhFroiIHrC/oBC+ECsAVLkEYzElTpTR
0HTE1/fzJ13tyCwW/p3oIsjb/zWVt8JH5gJtYfmKqpFzKYKinVe0Asrt5My4zBPJ
QRX/l0cgFFI1tpZ3HdQmmK+QnT0Q+7AF0Hcme8SC5R4K9U6ATuUzhDTzmQOCWlbW
Dp1p/oq6CSnZlqaneG3R4034DFGhEyaCHPkf+uBaR9HiOZHCWmr4wmVdb33qh9Is
iZKawlyiLSVD8PTi/rvuEoR+olOgCjQXkDhihTIMGDHboil+XlXDXs7mBWKKk25T
jhY3efpDrYglJNnn8AQxDbB7NhilI2IXccPTfqI2L8DxzCdAFsVa5383/cvdcIZb
9FULapdRvxE/RDZTCrDfi2bzfbgitXXSqBu5xSmthFkbYuRwZV8Rt6BUkQKmbPtR
DT3no5l5TULo1Jbpm35+EA7/cH6WbTBch1ucH2z24qkJuvQU6GEW1/rTA+D3wXat
ZLgGghYGgYKCYrxSUKntqaFI6m9M3WgwjW1cD0b3oS3BQaLF2AhrRYz8pZ4vyTrD
/ABtB//y/boNtoQWCSpSCa79SKpkrSIs+ozk4tLRPS00wbOHmKudQMP/rS7bvGfK
xIGU3+5WPAHpyvt0cSGxah7eDRzApRXuNN0wycMulO+uG5ZXMNVHsj5FzyKgr1Hx
sYs2kHgovfiq24YU3zGUwhovAGKLbzXcwXPIzchBUqi0+oyduvdkLHWR3eOYwmk/
OdAiJTCWaRVzX3ry6g5S0x31hCsq1SglvqHKxeLzsUd6yDF1p7ISF3UlJhptkQBW
sWLVXIWG5IyGakQ/gx5GQBEnHdgCumVv5EkRR15ZH3Pv3wIT7iiq3mQRSXysRH/Z
bzQoESGsi3XoxThyaHW7SvOmBoVFTSmbyuNZQL4gzSeSHC84ryMXIFpCRUfX0zJR
1tXakczgRbI5fFU8PezcrjBvaIP4W1Wbw3adqSnZ5bS+f0YCNa59h35WThXMl1or
YqcVaDGC20JRg9P+gNloL1+eqJ3FlZgSUcW+lXmPEzKRKv6e0wj9wMJBSLo4VZjn
aT597HJ/NMCrYtydNQvTSW185GB3MTMnJiVSL6E4Vo0FevT0fsfsc1cEdbLXxJlu
FpwpDZHYuB9Gr9jbBLZQNyS8Q7koTi93JN+lSAewluxd64xJ1NOvm7Dqb8S36qww
HGs+DZOlZXvc5uRMa3n9jzHqBXttKOh21FLayCpsbks2jvc9JYCnCt+4ysVajKbQ
TsC6OrTscARKh37GBRAdyBoOARkHJ72N3pOXJGgnDwVFiLU+/T6zOn9NHfrTLYjL
rqUwfuXjqkn/W8MPMPkAiZ+oF1whRl3VDJswn9pIaPoYxBxbESoXk4YDfAwrSBaf
GjqulkOgrbspBTRYlhRSpxRc33UF7AXskpBXx96XITG7kN3YGw7SgqhsKCuWWPsc
eNu0znREt8NXuN/8VzhE9urdex+WzhUzqn9POw9sa7Cg6Rh8r8oo6iKJozaPNlvP
/lyhfFbvl8E43G8vTzYRgGo+d8dV6MZa0F/fPh2Fojz6d2NZyLwIIVK6UH5nPsk+
+sMSAhsQNOZSvFVo7V+H1x1sRZXUbNJfOP037g4rAztbCv1q0x9PKl3rqfTUG8v6
NGydXj+frHJyCB0o/TS0UIvuvRd/EGdCyFbjglHjubPgPBvJsiTQojZ2p7vWGHpx
i7UMFbYRez5B/CX0qV5C3si0b758ZEpiAb0ynwTM42dUSSiVz5gCNPzJEwK4tgyK
w4bMo8UwkZHAiVPDNqHTQQGZtdh8D6lF8Y/8pGLLcfVenGML/eFCUe3S0DNkBdIa
4uBT05uCc93ZZaxzwupbrId9WrGdicrbcBYCHxlIukOfTzA7j07jOHzjSTZpJb2t
OdvTOMJwD0Hp2Uhq4+InxEfbNRCj1UK+QFwfO8xzj9gIZKMS8neI8om5VCmg9E9F
YMbtTiajt9RcpVH4GTiWYr/woZlnc8Zeg43Aj3wNTZJnS0eaOQhQK7yb+MqDzwci
+cwL3BjoGjuDQKbkflXqY0WdKYDAISh/di7dgQKeYnW/krcEsF/Irkz4JeGlRx+H
QhYraSjrkLPQDDixRDJeTtQ84y42EL8jQseM503ae1pEWCG1lu5S6XLsCMvk5tHn
QhEBAmWbZjVJhb4tMF++r3dEviSzRDcElJinWuwO9kVHZKkuFpuTH9Drb2746hGI
sJEP1hsjTGticdf1uwci8MFzJbwulEV8VUqlE9rgUlDt2olWhdOC9SsDTpnWKwyl
l1Rz+tgtKzBM7tU1VOgBryLf3w/jk5KsMYZqKkicY+QmnpytXU/7VtLN+E/E3rUH
qxk8lZ0LtlyfJGX0a7OMTOmYhbpWwsaTbY2/FULwQoYXez6NzkLQpIu5TcpN0Oa4
X6c47WtCF0TQ2TCXw/1qUaPKaJmpGCOXLK8KElGpXGg5psaFI/JW6m2/k/+UDupd
zLHT2xD+g9V2WLlLKmLQJI/3s+7SBXZCJdkb5ZD5jKonUqtKYNEGzo3GFYP5iavG
2eaoz5lChP5hx1K6Vt+9dlkad9NVQe9KxRyo8rpXriwJ0meWj4l3Zt3khxes7tFm
NLIpkd3vTQS4z8ij3CEMXKWsQqUe85SjbmtkEx8hgorFvOxAezzhcmZzZ9xq56zf
NiJn4ACR1LdHtZqdki8GhUb4eEX9m/geIMLQPcZkf3kobWqwIFP4C+1SkagNb70K
2+EPIKN3KP7K7rd/GwrQe53JiZHJTnAHMAJZ9RhUtbeCN7tL8BnkDc3potRfxMHZ
LijaqwcROC4e4ZkmV/tgyDiJE9+kVDxzWsoFYYiqD2Xu4kiZ6zMi42+E8ucGdni2
Dvu5gHkDgmEQV/Nqq8p6MtCcDjR2JB0DCWMyx3dL8uKZ7CUKSOeu3EWpRckJ7FCl
RINe/82yEKb/MCbnGQ5SxRECb1dsD6UrRDuv2V6PVomteedAjQw9BnY6lQnpEkn6
euGWrDPm4dXx4HoGuvwEKHb6RPqi6fFqNm0FcNDiYnDRgAjqdd+HHxRcY9RYw2nH
wmhsRb9hMYLDEmQYnmrAB1u0rPNsQvHifR4ghoS+s0iDFgjBlfeGyMFPW3lgd57R
HJx1mYHTzA1kkXJZBEonmhsuIW9Q3QtGVRdzEcv2YRpYCIC3qlL+/sLZGB9LMgNW
Jd/DXlDk4aPP4G1GrIHAamqzTYTVs+TiudBoV1Bf40csS8uGVqIYQta39mqdNUy0
ZYGX7Tf1pSWdDpxvNH6tosfiAYGE1dzlbGbajAYl+AuqYG0ZAHN3uInu0ZLqhuVO
HiPnXpqfDDesN/uqP82S902L2bpYFG+qDtCS9Dnv6lGvARrw5XuwuAk7rq6eM7vu
HyH4KutOAc/Q3DgFWdm9FzSg0y56pn/CqBwz4Prg+g+X55iQdF8HXWQv8QpgTQG4
0Kglysr9JVfYvtQCut3xZU0A+bIjhhyg6ekTklehj6VJMyTS0Qix6zjuZkDsJ/9D
CpoePgP7IiS3Q6yLVnHhtpE1oY7uJRVB6aTGlDguXC7tie1CrAy2DlBKTPpirIyb
OwYBRqei2/CVdJbNAlS2EgY0vkocoCgpZ+Nfn2nx/FOKFsnwMB8X9iay2pkXtlkD
AjRGKkU7gi01eLoGzjoTo9IMVwPz4UXBmNFaiu8DGUhKSbb4sbw24NfBGziTRpfs
J9imK9QsaMSYIej9QrqPWnPoJL5uKVoStecGE7S18K9hZ4mDpn1kujFvKPyolXJg
yoSeVmj575JeHLxr8eqQdFH1MqiwBBS8PzHb922wkpaBOaShV3CdqvW4pBylc3jZ
ng+UIrA1hy/QafzNaRna6r8swvy+bmUUq3wU2J6Op/pHrs0B1f11qzcNaW1QgHML
1Jep5UuZrez7VjOQeTdd1P9RcRY6vXqkgXJ2u6aO2p+TMYYsYqwEZvH6b0paGKe2
/4kDRGqqV97+bkonR83Np8MAOVpvvySAn3SLb7G9+mh5HV32LdfR+nXEPhp+NguL
U+Dx7dVWM21qI+GSf0f+fwO0r++IO1I7sEQuTO9csf6uG5z7Ny8QMZgOsf7cQpAU
luTrV8QSiHNGNz2tFpTYqZ/njDyATU2e49FU/54WL/WW+fSuYb4AA7YkBmnVH5jQ
0a/OjEbj27JcKyu8dc6GUKMmGIunuEhzchLMV6wso5/giMpbgoaCu+wjxbdvn7Fp
eH7PlmAeg6CuT9Zh36/CMKypXhGnreW5Ulx///h6rPrUsk9JMZOEUERs1rVXL7s2
hBR6EyXmGzRKMkyy1as9SUXQj+XuKwbfjFn5f/BKee35gD1AvtzbAcUhM0nQLv3m
l7ryJWpbP6cHoC5arR0wsLjOibvQRIG/VfSWOromwbAS6k7nweCcza6XWUBkfV5k
XDoh749ZoprdC1bhVd9C92JuxYUshNDsVRuhHg2Fp0AyKwQJBEIgYylb1Un1WaXE
U3pA7xnl1+cDy/od/FzW08QddHL9k21Vrb/1mr8suMmG30BZSDFa3PAtgiwlvlSs
RDRl08NeYNWDt8VUg/vtRxkGG+wgQqHwQFyGfNkwsKJEG5QhChjywX+vY9z6EZwS
ZLkCKyK0jCt3T5XHfeWDapQPNHjaUID6tTY3n/68PI0M6csMQ1nbWH8gcV7Ub2/9
/dvKPaT70vdjdF8qjRICzLo566ML3fMbVStDnDSLkHTl18Pw9njlvo5Sj24md5ut
1cxuftKkBW00dxTPqyY8bJy3SG4oqHc+zYCGTfCOwoHRnRkCwdeUVR4D5A1yMZWX
U4uz8D92RB0HCILDXpsXin1E4dzr5bJx1j/D86EaGjaQPykz54HN4wYMvtOs8uZc
O2P9YBD4v/b2EByWCeXUjJBtArRU3gc+XlrMOqrc3L4ulewRPSvSKgribGsjs24+
3FAKOXfFvyYQIaOtIF/apX9tkuioAv9M83fn0DQau9Qr4B0+fUYTzZs1bx8SntGf
/t98uXaWpE+ca64p7ywhihbDiF9zcoh30rXS3/5cH/EMV9d8HGLLSuKzeJFcmwM5
AI50f3piVrAGDUyy/W7/ck9ZUx9hYDazS3Yc2+U5ljuAkVMO6hx8xTMNUE5h7oCF
MPnXpSaVXp9gM8gymTOhBPSq/7A6qr+O46oQfJCHH3VWyI8LzOsvMR8WLhAyTxzF
joLDK5T1zwnHVKZKh6OjCkOzjNGY4V2FhNogCL0aFSecRHcce4qKG7N6y0hhkyeW
FRcVmjnWWqtshSy1SAqjtAvJrNBiyoHu6BbwAYVHnRZyyWhFTDU6wYmiG0DKSh8j
7cUnw01C/4RYjOgCGq16AkklCoetePPD9HTsxazp62eUyCrARRe2cBZsLIFdjdpR
kKjHcU+Rmdy9/YFlWrLCPK4eIYpg+jDtJorLxdo1+av6wfXlgRcX9+XFz7MDRRyP
V3UMKz3nhC2it6lJWj9GKE3HMComF4kyUrAgYJY6mASrh5U131gestsjvDCBuVkr
jTuMsi57DYTDtr+ynovb4gwbCvXpGhj5xtLFqqap8xTzRg2nkUz6X4Mdx4hNKKYF
kUDx0L/lJk5SdqR4L8C6vIjuodLOeGE/5E3MQ0XwYpVOPTLUcH+8lQN9E0mVQuHG
bavZA0O0geuaD2SdkynSC665cbWjamB2H2BaI1W9YRw/poFYOmHZRHw6ZgEW+r5t
I3W92TKK5kmcZs0ITXpY1EOCOKWlNot9oygi79n+JzBxeTxOiTEvBYw6y4yDXbrw
lR6NNhORcSESuGAoph6ePfxdRCSWH5S+27E8S6FpQZEWjKQwmy6sZZVgDOhv5ATi
6rIlW/9lDR+/+yw4rbY5rPTTzqeums3QF9ZNC1BJAGchtsxecGylwl/Tb9od5fFM
Y45Jnlc1t7lTXpYVmBR/QevxGgRFhggsbnCGzLYCjJtEx3GgpsC1uKtyKU1HBefn
EZ72EOpy5nx0FCCLj7BEHJgF+9sM3Z27PpKW+CXgq+RhhYdNL++o+G6KpvZM0PbZ
twM/NbdZ1ksvDvcfCAEiqB5X0VTHvtV0KeWx06nn5DLmDk22VxmXwUEivvQR5l+J
K4VKWARUy0zSixkzHWKhCspakY9+CZosTPfiQ+SSDGdpKIQxSS3YzOPw3EJMnZnX
07RTG5FmpX4A7ai3EpOTnRVt2K2fj5KZ4oZLAWc/h0PTwkNSNriBtZICT0ETPUSH
hKL63LSG8grzVAMQCx7O1Lcx3yg+p+XDmEzKJSafG0W8m9qSSBo31DmZeVUzhIx2
LQ6pypHYd/ranyYmG91gJFYV4abYubkBCQFJvPy5Qq1buQ8dPk5sIxnT8Sf5xvi9
c1sBT6WKJvF58UKLBXKXg7Hg8Erjh/boBF0eqRlCi/XLiG5H4W101433JgTYFmRB
JlpOLyhNgxtJq1PG+BPAYZX7XzImjpQnl4pS/Pe2XaVBl5SRXXtkFhpcZh6oEyfW
sVYeKGL1DhhXlpE9nZxUTaLWOYNu2P46wLfSHTgdaP9gdk7LXplhiYFklzv/VTFU
qc0Wm3dbPVFINhBeYGxnkLMDGEPqUH1lq8DQO6Uq7wMAHv6YvDKdmlAcY7WvdFu/
fhshWcpgw6iUwyrKnqcaE+xsnt+nCIGP5bvOUQN1+3e8TJ2grRmnLMhsbzW7SWRA
TKX8ADwrIOon6URA7S0B+iZwV7Dv1KO7wvEmWIVXmYGY8YQZFDsTlFqh069DT1yH
lIzmpzFzFh7hukajeeCd9q5MM9F4IwRK4CywrJQO8YB42s7cNm7VKJa0sp63d+Dn
lqS5/1yjSTMwRvptsHVPIanVsxgLawgw39oHJu9mdLiVLqGSdTLm0v+you2PMPuJ
h4sVJS92m9lqnMHx84MDkrdB5ya93zjyfDH2OGpb9UavxeUzkCeL2Zlv+obzELaN
BJPEBa88BgPW84dpQq1V+xK5b/vRMvRfnkUoXgLh+YrIphMU47I1wB+IYTX3ynkR
/npJBupUFhWrlYk0y8l7nIDcPQW21PCjNxdxYXcWlWb6M5G9mwGm0h1YOsKUAjMe
np4vdx55g8QUPt4DTdlxVGn/UsSnb9RiBfaDZEvii2FOVVAnzDVXVURy+tf+6gyS
Gz6CSoVegAHGKwb92wmFEByBUI2Cc0Q93LFYPp0QEIti+D3nMsUfQ7uU34LgWXgV
0qWrqtJUlxYUoSdJPFgBthpDX7WOpwWaU3E5aQ+BaLNFgDf7VRTc1wdfhSi8tUTK
+7HMVYsTcDRrep9yYzUnzmflyD5j3+PcX3K/kqU21DghR2jrsjD4Av28PwEXD6MJ
YCf4WXoqCIpfA9tmxgSoEHTda7uN1fJtv9EgqAr4/eVEReoUiswhIaEzTRH0CM68
xWo8b872Mn+IJL8tVt+R4xWkUuZZce3343hAgSQQmshRv1mCDYUdXjfRMZat2xPB
1J1IzEwb+REVL5JqR28j+Z5fNMiDqk8hIxIWKF7E566h/R8Omi9r4JUHGYdk54lE
wte+J1uW0r+9Id/uarTgyJ9U4jv6kc39DdV7clxB9HzX7sgJ7+OINeLnCeDxbg6k
EqOjf9dGOYIMhChQnGgLF64+oIUilN6q66Tan+W3A4Gq9KNMS9BxmGTfYw5lL/FC
dh15RPBAQKaQMarTgADw9+Xt60Z6zPITQ0Uz7mxZ5HhUdF33svszMkG1GGK268gD
nENu8tR/Q6EKfhEu8tho7G/FZkxsrlWls5b1AJQOgdSJljeFVrTLLmyrR6X9hkyR
lpnGVmApXYqx0UnkdPLk49Y9Ewi4b3DFOoVG0Y39cYtOHF5Ewod/muYr+7YDTrwl
N46/xNdJ/VOCgXK3SkKarQ8X1UtAzO38fMch8rUOee1yjP/vh0I79MZoc8ps0NI0
D6Y3bWHRWP9MJbSZcnlL3fXKzyfOzw7R9Osk5Fxe7ssnUUPohGskvM297vT/g8KT
vaBiG8Dfhimiknmmmf2q9SXmREdSsNPsdUiXVLCuqxfsdwiVwU09UrQxOwJVavOr
3PmV26kPyr27vHUw7Jzkmx2ZEqqfjw4zgU8L4tdBu51TrC/n9y89sCFnyXgC2ShK
8Bx2tCznjqQtCxo5AUqPLQTS6HdWtiRp/cnakUyv/yeaxNx+6W2drJML+zqE//Yb
2tDch4R/uOEIXdTDNYgfvyMhstbFmhnbWrowEuA6X8wftp6jYJlE0sZlT6/6yX4E
R/0zyg6ZWuKH4jYGNLO4XjmnGaEQJovByucDznA5++SnzZGPycKi8nwxgVDNNIHN
kPARqn7iOljv/TyOQrmmvpuQ38p5N0y9tQR5iPlEPJ6COYoQgyS31GX3Fi82XFBv
9kG5wbEniiI9qY1ttReHprLH9aHAsCAKTKUE9qZV0XZhCfd2NzYSDhL8JOBhXmvf
DFkGfITUPfhpI3RXcidaBWZb57mhe+RtRuaDB2LY7538FN9xmY/lUh/jfGMfp5BY
BcLKQu3HPePKlxnH3rK6enCoJXXaWy2608HFWVX5SGACz8yZJkN8PtGBS7zk6af5
BAI6TBuP2zsajIyR60p5VBr2P0OFB6EFKWAtqG7nUS5DMi7qjtevoIbyXczrxEr2
vzLGiSvNzonCukgTal72QNuxFMvJX2YW/qChv0OCfFQULDBKMOTJSh5UvhEUaNkv
1plArEZKbsxOknqcDjunNLabZnLjUBtPWn6UGTNuyYyjVBj7Uc/VoP/4bvvZBALZ
bYi96CDGakC3C6qKCcITGTQ8X5CFa3Nioq52c5713cJC/EEmTW1sahsWX+LESFhC
rRDmOL6JN1kuolt3kKxQJ0t+4W8WW2TwzBNANBewCF9CALMYMB67t96sZzz1k9HB
CuCbK+PfBMPwqRebfk7YDKdn37o/w86OT3ZgmNtASzjIPkACx8wnCBj3uI1oZrLz
65zbcMa2q/42bY00NHHUSEWz6+58tYp45AMgNoLDtuWDMyk56FP5L13buDRRafYD
M6+l14H2lPuZeuOJVrwPocJyXRH5E/FZAZe+Ei9zsSW+lw7TiGadN2uYicyVS+wy
qPa6WiIuj87+wnWCkvToDOlrlvOPpHpBPhI0vaBs03xh88Q19HOkCSkLlJChu2fm
LG2i+vQiX7uL+XcvhY5MHseY+AW+6rlY6Mg67IhqT1/6cWV/5D/cabee2FQl1IMq
+SW5+oFxPbRYC7IM/eDB1xJZa0bzsZxVAIHgeI4Bd7nXXFHEAMAXjiiUz3nb6aHH
IxD2rJkUThPVW19ujLY5n/4GLl1FgL9vHHVP5SVd+drVspV883ICjPwMNarg9qEl
Hg3EywScYoJ+XdDY6u9arVFeZBUgYN/yHbx93CpJ3gCxZL+/Iafv8sYoikMyZD77
VLFvpF9u05fwD0nlSnp7SmU3v0MHmxI8KwudtTlhw/Cba3SyT/ZFbjaseZAPD+L/
Ep3Iug80bs8ujh4mt1C54AGCJZ5vnqwFlOzVUEZFMEDlLovEPToYBLvexdcH8qzf
0N457ebC0OyOiuScQabURjTONJfJhjPtxcl9R0k/C5qTKRGwxGoyz1+XBFzpNgk8
0a1N6A6bsRBt49JYendHJXbbWHNggi4BKRAxKA1kJxvCb7D6EfbRFeLjb5HLwU5F
+nCi/AO/aM34mHKKPwuXNPIoOQTjqoQaG6/g59cvu4KASSbsZRsMtntLJj6he0k/
63xsQZX9d59bCQ1/KygggZA2tgkHyyYT5j6YdxiROQV41Gkg7xiBpJH5R5l1UA+d
1sJ1su6AbdkZcf/3xiEM8xOec1NBwgwGS57Z+z/RFN9m0ieD7ANSXyR0ALPGJqPm
70wUzSpquO7BI5F8GxblkYLkbiRP7D+K07TJItihBccXPIqZf35TNixnnE9qbmGS
p4vRSemOJYSE5HYSWZwI7IC/a6yQLB7O03u9l57b+0v+4uhDSOLWbAN7FHGfJcFn
NiaLh8KBjv2meJK2KlodYVlE2J6vki4jHpsUlPmbBlKLdebLcUiW6grOcvrtjQBZ
MFgeb3QUPnHKcApId1Yow5i7KvirnEikGzu3eoNybKQeObRHDj1purBEgvhNoGL7
gBBAI00TeJl/3UwFy5+5O5kO8QOaOSC8j4yDoO4oC9H1+ml2zSeM1pbGqCN41MRn
WL7JicTZkviTww1EVjbYUPxd7lf11GbUhY807JSKuOlWskzoj4Cr7qAgfzwbV2ga
STsRglyPHa9XIeKL1K+cOMpbu8FOnHUUew1lqX+IdXQq9cGExtSrjzY+Lavx//3q
OU37A/Jk8nLrEU4XanB/qdI8vOcmZHJnGQkW513ydI2rI7s/HRgp49GG62G8HkNz
/dtSMIQIwt9oXVRZYH0PDrfVFXk+fYbCYQWeUcwdd+FcmnaGYEjKlhQ0mBpyOaxK
tSuJ18nDNsUuMicuJ7llwO0xftiH/mBRmnBJvR7jXvMfdG9u8TiWE5EJ2+hLXJQE
KIi9qkh//AKex4T9Mgp6AKabCXliYT0jUAPRbWIo0jZD+LFz+y+Ja1DFAG3t806m
ntdRxIF3v/8STl1JS6cKTX3OhZvAH2fp7HNZ21AR2RUjYJ9fdWZv0d8VlfMUomlY
sJEuiplpa1/Z+KyC2hdKvBJdO0vUnfBZEqwaOC6xvGQ6uz8ml6YRJ6ew43+T7VII
gngplNkhtwARcFPZKZ8VourW65zTpeNaziScRdG+R83xl0xKCsBmvrODHnQneZ0w
MxpQ1TwsuArbruBFmg43zCycThGdcTw3YIS0CK1su+o9gq5fNU5DANNcu+PzNJRT
oAe4bayJ3KnSX0dujLlwjsfN6HNUteMKbjd+c1T5quJOcKtOFGF4r5kszs8x30+Y
cWd/mDZSk6c9NmuN724d8jPcaujUg61tuTlQenVcbZz1YRbqov8Ff+bFJM8Rratz
cNUIc2dAIr8jivS7GsSUPtEbl9cpvoTQ2s7Y741IA6Hv/TJjcMuWVlh1lw1X+5MI
jYIpROAjs8SSx4ceylNlaLKVqe0DAjGV9lJeU18cp8lwfbvjmpjkWQS1OKVp1NOD
f0M2htv1r7YqwkPnIaG7qgpQVA/Co4AeekjfynX8+p6RvB1aHbZJbnFfwEPqv8A4
Bq/6R9/7D+sHdUEx3GnQ6dyEo+MWMEJeyIoVB88/wiCEqZStpJJ3zCi1eINYhl0G
BmDiO1wJd3U0xmAUTNqhEoLrJqNKz/JzZzLIw1Yh3nvPS1jUJqIQBFG1rPpSK5ze
B34p0Mq38bIwY8PUZMCWfJzK4cptKypqZBY9UuYUX6O1/0KjyMsudrjrh8NcJBzI
GssQn4xROWQ+YPmXGj5hDqfZJ9sAkItN6FEFGmTtECnb5PRBmpW6e8XKDs76fkSd
UDnj7ToX5S2MFGGmMtSKPLfBYxB0gOvi0MJpnYp9W4mszqSKZ6bGAQXCgoFEduj4
OPVbcsPEKqhh6rkuEQLHCfEGMtrVEkYTVY5YDuC2UxwkBsNK1LAI1aCK5JdbG7TN
+PZ0mk0hIlcNGQjQdMtLboE+rcYRyL9I3eRA/hmQ5QzF4kK50HFV9yukSbZnPelp
cv9rs0TkqK5QPXxapEvrEY0WIemmQy28Ysi7UEp9V68r1TVb/QqvZXfuycFj/NcY
bswHBH4fT0uw/mYnHEIiwghqxDCB6h11MpTqBjViBFova2GZgiAgLS7mJCPOz5Qx
ZFuMPi5BzYnAaaTQQt+xbQmlHwWuwgq7/4PfWBK8xIdZUa6gAe0o3KoP8SkJsmwh
yO438grW/j4NSmwmJgtsz0hWzrQ+K1w8tCmxCn2pGjRBjxWuCLqlPLcgoyknV8ER
kQSYHIKY2FmN3F+Di+c0+f1gDzfMrs2yHo1N3MNxc75RF7u5mo8yHAec+xOFCD3X
kRoFwuHZTo4jfLCFpmVF8U6B3aB18HacEpZ5o9gAtV00DwpfaIqn9CkW5v3rX6Ac
akVAHGB6xcoxSZATl6QrvQPnioHjcvQUuKFFFYp1y1/rI9SgRnjgWwkL8w9c9nz3
Ss9lXwbr0VAipCIzvsDShqtqEtdcpRuyAnNTKW+mcxMPSd8FqBWpItnD7oHnIqeI
2VWmduYkSJlasUxLqCZxqaK8kohmJsP6h8o/CjJ4pQ+/GY7GbMW3Angt0a5QqERb
punsmNHHkIAix0/3AZzn0m/ZsgZmWpLg9JCokjB9sQA2HPRsB+sf2Z2f/FVyeHXd
mjWYYrzb2W4c27dIEO6nkkMTjofwGcPESoTwNkeE23j1iBQMJTKlXHeeoUftPDqM
ueRh28I+qwIzntp4XYYSKKsHPpUPHz9kQNDhdb/+ZtYFOANYEeV2YaDJPbpQ9Ax/
sS49Y82EORKa7TOe9qRMWpmT7tvUhVWDk5sHme0t2Wl3uj8EIml94fj22PMwbjWg
Nshw7mhQSTaXPFCyuQCEGMF0Z95pULmCESizrIlzvZBDKlA9rXBl3+aoMBGHwupq
QIy6cH/uFEhKb35Pg4MJ/0Lv6XlVwQ4aZocKSh+m8RhKsdhgKw52TcjoOOZjXral
aDofBgD8/axAsO3BMPBbbfykrqVO/hoPp1KXhffnymL95sQHfMkHgX9Y+J+YNJwU
dpq3vV6g0NiRHvyadFGw0VuWmRe8rFmvtyr4fcXExTWYkOJH1I9EqOmOMXdueqBW
q7Eo0nR+0hIpCGeabzJlg8f/fVtK/lUJzPYkYeomY/hbAwhOY5rEbBBwZINaK24O
tZKdYg45awlAuBFjkjL+8FJDNcj25ZAlYfWxtZwV7WSIj2CxwYsRRRobBRhNbhvE
XXROkVSwjIjVG5eF6NLibL+TwjJvI3D3QW2T9v6YgJFBjuaBK8vmYZJKMVIkCc1D
I01RaRvEkcpFCXnVQetwiKJMKXX5Bkz8upkYNZ9kooRp3CGmAjuA8eeCH+CUuRme
l+b0B5Yj7Xtax0AJF5aofKX1UkMUULW0IA18tzh7DxVuEBIpSNhrL+r5HIGatyWX
PwKhnj8vDt7USSlW8nYrhj7btogPgo9BJI2aHrhYvTQueHiSV7vSvja9GL1Vr3pb
QvA6tCy3PznK0SJ1rNABtzQmXNLg6FGKvWG6Fk75wCwlFylPB4D++KYSlpqCXkF5
HAaNsKbqrgms/Y1lGPTaCdWjDfJzqndNTSfOSRoLHgVp+s6DoJ+YH8M0ntjz6P0p
PBulUXukhoP82MauMpObR4fPGs2i2BfYv7G6neg9uBcfmnUy4so2++KaNOsSGkbY
xr28XTXGnAUekKa/IMk1j/9GmkcB4ogRkMQ2IKptJvf+GjBRO+PAp+hpoORR/e/o
ECSAfcb3R/gUTDB/0QZBRjyQtMTGkiHKUP4HwnXt2fag9+XQh9lUPTPdc4VD6L/K
6BiMxfu8CVaglWz1akCOGMCWSe1vkw0498yAfuDdTNyFC0wUo7QIerpkAdrnMCkk
g+UdgzpT/OOzEXGKVZ23HjIZnnvmY9w1EUyfz8bPYK0ZFt6pCMJZN6geB+3cJhEF
+dJ9Yl+RlACrHzCFrIMUbQTEKvt9b68BGRxTT/7BrfbekMN/zj4kh9YqPs4IxqOy
03Pc+F5ea+zGN2EBzZDCq5x1QyygLuzOS4FooLY5zycwF2pkc6MXVWPjE/E92+Mb
DM48ipsyMJdZ9ET62BHi/2n9VkxN5iea+rg6URdwhqkxVe6+U07Y28GWic7lg+WH
2KtiYu9ekuTyv2Idm1LMScKXdUa63HD2r2oTsucObIwRNijtHtrqud6hnAHvRovH
W6hR9t/eBxgmTwu+O3zL0eu5JLb+Fysv5P00CkAi+bdXgl/pYV3/zDlUirFEbogu
xd+pHE055pGY5zMl24O8fPsdjpaSeJqKRkw2Is9ND0+mdQuQ+JNMFGCT61/TeB8g
0nkolPYgebH+BjKth969Y/Qzolr/Lu2YiQb1BEQygNgaTlHGNfc9UVP42n/K+gp3
hpAebKb5CCnHGRIFfkjf615J/nKLEYjbTMxpuQCc0MfTlqygjCm8BT9vEU6WbEME
JaWZi6kvYIwf0hBHdRiOAACRHemjsCJbn0+QpTROJ48HOkyxg2wFfQ18wV0JdtWZ
HzbDCYL4u6J1DyW1ROhObLXsMYW/ilG1HAtmJO522ffdEHFRMeyyTi4Q8FInzswX
S7cvjfT1LdP4IWHgbGxYoxktTnkBjS4ofPJaF1Hd8xz6OrK9DlVrrjxE39cf3iDA
QglEOMVxKnxvaPz9Kun2f3aoe7driuHP3aYRXh7T05yqjH25iMdP9hvQr+GFN3+q
Km4fuEOtzmak0r3epP2AhVgIXuilQszqRhHQmdc+pLUGjQl+3fA9cFLC4vu3q5GY
C9KDRccIVFCMHL0z41r+W2DVscNMODVM7FcqDYEQ+Fdpnk/ziKO2alWpxYRnV79v
wW37r3EQJQh88i8PJeeAcnCyYtNdEQ5gE3aEBgEApblMNkFbZIxU9G98XSosHCz5
EjS4ATOU8WR+3NBL96K148MTLlloIYOBA2dI+jMx8PL7q0jkrqjlgDMO1s+n5Ut0
BfZAVe1/z7g1MjmWuJ7uPCgGikWuxqTaDmDqOMRmoO5c5G0n7S8Byq7QEi6Al9cz
eMXTsFNOqXS1E4WuMr95AI3HwYqHLUOHSFnpcDOqONb2uOSbNC2wBTYWSNDTQnbK
IkNzSlFLGLjkgzInU5NOgfEdhk0OfcspY3QZeiRHnGmXIjS6Z11BIJmZBu1hPNuu
8q8yugwq3/ba+6El9XyzY6vW+xfD0vz9lI7jCAg+Lz3fTc7TQOWK1v9zvmWUjrmg
JSd6sXC7kvAIS1vqMu1eNuypJdwf4LmU5JEE4PXO8CU//tsClnhjS5/rvIG6c9YH
5ijqOm5kEoYDUWMFwmKRvuy0I0ITN9ZUb4lSkb1oetmLuD17pBaMnPGwnToZDtTo
qCPB6F3+nqz+cyyRid6kGwXNBdBt7UiEOGcQKIzrLsn5rIx1G2GeAWv3D1Ha2YOR
9Cr+0LhpouISEHGPdvjIbCVGBXo/WwPRfUu3UI6tl+0/hhZl8FbZq66/Sp/IVtrb
bF8XlHSStPOSkI/HF5VszRhbX8QagJwErVhIT6PzFlO2cz7lpeZHzcglzCeBAh/R
lSP5DJNmkqbp8vyzJjb3XLy+vLlFqaI0NUAOfGuC3lud08d678d6GDnWGJwIpAia
SSn8PIf0AqKjC0P/fwkCwuEJsWxx81j71Uohgq5npGBqef02nUH0LVFJRW0zW3HR
Vctcd5D1+hPLrffMGU+xRYk5pj+4/ywlJWvFVfo+euhaNIlT69zq140wf1XG8pdU
/Xa5/zdr+5y7cWdxXn6NGYdVI651N+j25SQnvLPQG9ywSsVXTqC4DI86M9j9baFa
lhdE6CRMBNM33roHPZpWUPaznDdsgYEPeU7HovHETB63O/29iACXT/9onP81Gy2w
rHElnuw8OR29097qiu7SzOVhhogsKAbtaPiX+Act2SasXihanOX/7eJXKk2hi8H0
o898lkA0PiEfwd0i4xSfRqLPEbBMrC6i7iBQkyXIff4jSYymRKgGzsgMt0sdqdDp
0CgOB6WM9OMkLgJ4EP1GNczb4UOcne+ncW2QYfYwnk8kn07mJJKnEOs9PKNDvSvZ
C2byC9clFPtXOW+OIeyx7pC6zPmBuIlNX4CVOLN2Ke0/rAN7iQCXe2TCx9xW9NHl
N6T20gUHxOGbCmIh0D8xHITsrf9viZsBHcuxzXmdJv4JxKF6Rm1NI1VVtNVLKzXx
c9tPLrsIGA7bpSyPmfDSj4vf5Mn1Cr3iXZIMfjiPxG8YGEJpK4apd4OpEDMg5K73
D2p8czgXngb8TwazdE9DBU74iA7QIRrXt1u3YCIrjCxl4VnMIX+3FDRghOVXrwg0
yIfLbYdhHtMI/tOjfTfNoqoE1sGWrCBBYmLZ6AB4NV7E9FUZAxBVB5RL20xWRs3F
hIlEdJibVDjsTi0gQAYf8VjPeT1B5ikYiW2V2+v3x/ItHEEBQUdjWOF0AOjYvd2o
cyh/fmdGYLvk5AG2SrhHN4DEoXCmu626YHtdAz9LbqqVxy7I5+F9fYm2lMXSQG5B
uz/Pc1z9OO3NJDi4Nlryl4OfTLQb9hJ2f6NXIEJqNp8/HwdegRmrfplfgqlHK7W1
FDGtN8eewe1kLotckodYOIuYsdu6a0E41Y5jsbMBCv6B4mDNyJ2vpRxirO5Cp1P9
NFYpBYElYYHK/Mv5ui/dskEaokNWAnvlrSCwo/PMEsNsv0BHJjVCW4enV2OajLR7
UlC1RrDQAmV27Bz7iJM/TrLdd43fS3tT4s3Ppa700ZB1iM6aSuxu13TeEXK8JvJI
BFgPPeg5+TrKwOaTF9hWlEVyfrSFo19Svy4A9UxYtU4m0XCSLC6WJU2Px2+HuMFm
P3HqbzYE1SyhbyuI6YIymeIVS0jDpLuoaTei0gc5VxhzUO1ZqBcYOOTynOUrQ30R
za7Wf8StItPwDxF6Vm9kLa7ef+QxakuJP7pZ3VMZZMi35zWdekEcFbnln6P9s9sq
vQ0pRWwgn0cB6IJV2Biozw2ypRQaA/DHmMpOk5yIWN4juEJnVt5AvWSCj68PKJT1
OsA9+yorR2mcGhsPrylSPy/nTsVxSd7r6bqDI+Va3mGQz0QuLH6Y7+Uk0oaUGd4Y
Aj6Jrz/AC7bEoILPkmXqZ/qsGo8IPLzV5bRy45EuPDfhCVqHoeZj1WUjAYeR6IXE
Oi/XStWOVcUDjK5hxYfvQUOretLzuHtZxYG/voZJOBVUR/m7beayfiu/BKEhIFfL
Hx6p+vpiOKuTobqGj5APzy1tXPnT6CEwWDJS0zcTGiTftZgWIab6Hde98xgJ03IY
Bwv5zPrWapaSrSB4Qqjxtue2CoUbjNH1MLcUMiS54I2W72LFhgyoYFwJUNTqkMvN
auONlNNzYNDpTligyvyIworFut443ULyAiba4Ap/PmUQbDTzZfATjloRYcBx09kq
e5p3CGqk5vhyf0qEJ2z62oKJq/WSRFN8WVkbXc0Z65yqVkeIOvNQNkVs98CGW/h/
r8dTalLEB+JZy5Z37nb1uTQNZEpuF8eDYU7WKzf7kEWgkzDjNIkedDxzDpuCysKo
IknIzug2KQwam4rPQgx4VWe4qjWIL4hIHdlJtCzScqimATpfTrITQJ8X0ex9hs6h
TIIe5I5d41P4AJ5AoDIGmChsxNVF8NIyfj7CFekgH4aes+pDPc6BTH7gIGIT2OM6
la82xMbMtS/E/RUDNd0JEcg8MUvf4bZIHZFShbydtxMmqB7zqGdVZcsN670br0Rt
sHpIvYnkNuE3b623nMvO37w1/ZwDej0ropGlImBCs5HwYv7dCi0qDQyoxLFfzJjt
IAoK6nmEYU26uedASV5xEuStkDWDaNSzx+SOU11spb8qFF1Bc9CIZu6XIX2GBxw7
G0iRWh4x7N2ErN8ooiVrTo6r64DPSaiNRg0WGU/DslhB7RGEl3xUSs5gd//BYHsO
W6sWZ52gqWmL6qjKWF+R/aBHEDqOD2EqFFGERfr2SAgK3JRGOmTOT7WW4/AQ9siY
P03h9CywzdUHCZf6a+TmWpx2MFD47Ue5Ihc9AuC8Bs7+NXyHFHJ4CULbxPYgaS8w
EptjMTJ7pT2voxIALJHnAwSYstk9/fhMTpxF8UA3Qf8GM5zDIFLgRisKTaAKrjKS
G/cKk9OLQmmfF0+t6iO8IiXKjSl96E+0nLH+S7yFRm8ysSTYT2hj2+m/o97DcmdN
PP50F9r9U7nEf2nyrPDuzhpuN3WNpPneaAykTcbUUCc5DfRAKZym1G9zepG7J45H
9U8diT7tMbFWLBQCvKnACCAp09p9SSA37kDdLN39tIoRjgjBjfM2fI9hjHkvE0tQ
MX+uPbvWEslbDDI70c/VsaEYVvA4DbCXMbXQBqpMmJVVQwFNDr6dEE2f8aK56tvb
S9ECIVPQXRZuuOP5X6/NUfYULHdNB3I8zd8zEau3bMIqwZiXkMBuoxWx3bnAUdGv
GoH6BApRj0haxepfrm5fuWBQy1Fh3k7/hT6THh61pjXFMPozAJeejo1Ic6gVAX4Q
BKjN+vhKR4RVDhuksRzR/QG2eXWYPsUBhQiLmmIZVsreRMcvp6yaKO1wm6IYlMlz
RmlMKvGYWshm9iYgttsug7WRwM22p7GtieYHdM0bNgXIyP0x4p48qCke7beR9SKm
Ck+jcQdOqG0LO/Kls6Ma67gNn0YHc9zbbUvfZ0LaBxA7Pe+6Z2LkX4+XcLCzrdLQ
jH5hNxYINuPRBVcwBKbHxGUCk9tNiY3WmwH51Oj4Ze5iogYikwmpSEakRuRmtbTL
Mjb4wP2BWgt4j04f8rztNyE9I8n8Jw6WfQR3rOO+yX3h+esCoCS5o1JrXlPula4M
FZMegfdx0KyIFRLE0KCvcsiha6W0uhaPwjWTyjSDjuiw2yDbA80GvZIfGr0FF8cH
IcgtDwTkygAmCaEYKXShw4fC1Lreau/ZUxXZRkzsuAY6vGu9ZTBRhCuTIn3hN17J
fGHAVW5IEDH6k+hvtULVBA+mvLprAVyKHzz9KJJmQTU32lASIKoTWaqyv2aScmdo
WHtSGM8Fbo8QKqFjMWT7F4YC9l8Fot26DOxFKYU0O2zPrQeZ6l1FjDI/k9BzKtyy
eWtjm2mSvO5BbvegfDzQc9j/CjCJwCj1e4PFeOdX0Am4p8Nfbzsw78v5xo+72bIM
IfpftQy8uTbdEtAXpELmpQwrl3Do5KzOMYKObL/v5zZ+rbtQAhGtkKJlp8ORCjCl
TVTJvrjXcaBgLE6xr4wDCI4rABfcgbOeHygLBL50+yPh8TWHFQTb03zEcxjJvanU
/z9+Wl/HgAsCEZiVJY6EBG4Po14ktvvsF6k1LnPYxAE8N7iKWQONWWz36c5ibJj2
28umeY/zrJurJOs0VNqHZDT5pz80w2HwrBdadfEJGCewY/pDQGwE/SBQzr74m78e
3FlWiw/o8zOthpMfohGGJ6I7XTJtfQlFjhPTemNUeVlKX2ZgZkhJFEpORqw8IgO6
Ms4O/hM+SyMjYevodXwHfCVjZCnwWV8j070cJhukp5cZT2mSUTN42MEBBrX0/pg9
JexZtxbvjxcOw+SKttyN+iX3V0h8LlZ9rVH6z0gb8LxcvDq5njrCIZX/w7E44LKU
mV0NIcVhHUEUBLDpR7/msI4qW7oqUrXUZhFqZweqinE3pyQUv8jp7HJb1mG7gqS1
+DHCZaatQ+u9z2LJBnxnmxnUBdLEfs2nyTSwzDbdtcmMWWKBLw1PBUHE4iUV2kki
AWS+BWLDn5Fg3socBlOf3cvrgmkcPR2pmndfXxpVC4k2rNU7DDjkCZSLcpxzZ/dA
U6NlNdsCaagQu4/gbDVela+8F8KaMyEeA/gze/o/rz9hlPvMmq7E9/4UM+skWTZS
nkk1RdxD+2qHfC9Dnxb7LFDTNMQ7/C4LXj3sPauBtIM6M/N3y3smbAGi1+Vh188G
dQXUGg/EcU+8xSClGgP9mlQPAonRHgWR4Qc3Ere1PJo6fmzY9LVFxpBB5zo2FR7s
4vuRYr+0TV8ON322MWLJZtXccLDWK5PTJ+aaYYvwZ1tn8GlkCKEqhplSTfZaIKfi
ybEHFbRcsaSgthYZskoDjpXzjO/av1HcQiLRXezRkR5TLf32RbC7I+w0be+lg6ct
/zPp6Lsa9H5VYxDRP67yo3YOIEjW1MAlWNVPicT9E6273w+nIhbLFs8B0sjIv4Eu
04fjchxQ7Jvxwa/KGxaEP3qrQjIwgiMYngREjxQGNwfxYdfYi+VNJArR2D42gywk
81+HepncjO174R4l5ScOzq89t0+uecRFi/d8IZlEPOyCvR1XgyKkHyi78CJsdxQI
EzLj9piYpry0LgmPEpZ081vgIbym1y7kYL6a4tFZsKSteAQCG7bqJGpUV13FoRk/
acyQp1a4Vz2v7F5ljeAK9YghAueMZdfl5vZLdOeh3Cp3XkKRNUM+jEuxSbyrlzqu
xUzWcSxs6VgWMV+s4QKHg73+oQ8/gStvxetDD/MppM7q6ltApswkhcKl6NLTZPbq
EOO2U92MUFQ20ewB355+GWEIueQ1w3lDmLKd7i+uT07bjKX7u3D6cNC57M6pK7Eb
dyYwnV6vBfzNow3vdG5qqvniS1HKKQ7hIigCo77kWq92YWZwO2kI2Dt/xwQCUsPS
tOWG/DBShERgliTLalkmKPU0livl9Xg8/lkoinxzZHA/e/hv6K/NFWdDtb+dZVK1
QCN1fFcOytk+AbrsL0AS9w5YxzmnocSZx0C/YKl74Vdq2BVeMfPu2V6MNt5kBSTM
/WjTM9R8CCTPGQikvBTs4Saa/xIFGUBeSHa/bN7dQUfPt5aqGNCnYIKjq7j4lcwv
wcNoxAMVgrxPmefD64m2AH1A3qMGwlQL1CS48T1NBtmRDJ9NWoqBZv+anUJ2tD4U
AkHUd1THWYCFWpQDDKAfbjHOYRkIGjQ+ckwekXN3YlolUU38L6cdkf6jJxfHninV
kGUz9UbUNhFNCRuMn1NsQtY26Cuc7eAUC10oSF9DWl1joJhOjfwdLVOP6eWdTAru
rQZ/Cv3wfKIsyjggPn5mX3Tu0L2uMgIZWbEpv9CIk4yS8oecUucs9NtTfvwIcr5u
y3HFj5E7IzviY0gUSE0hV6O3TCSNgnNR1y6m20shRgXP1D4oHMw5QZHllQYXiY7E
6lFa8yyYicS6JbjoRvtG0NnyvRsPdhJbhfFL4wOiVlam7yA1x9fPxf3bXnCIfdRn
CmOKGf6DnwvwTaurDWDPXn2pD8x+l1rERM++Lry+fvcpF3XrdWcvORqWEtBR1Yul
KNcjT/1w6nRxSv+rFjuk3DqYx93uiHVtBKvbM2F5MmC+yizMJZMqlNAAQ4HO6hKf
qA+3ZAXaw1u6D9/6wsHXDrjhMpHkUO0lY4LOEBpkMqKv+7JrDCx89z5e1z5AAfDN
VtwlnIf7WZ0Ss6HmOBYMZPLRfjx///jmQgcGq18dJnufBvKvpUzXGao6ABsAy68r
Qf5qVc70cRraGpU5aKXgUKlN5BUHJmKZrftc6XzbYkPSh/w2D6z8M4KXFuC3ATPj
I2i/YO/JcY/SlEXPtRsF6SwfZo8HpxqsYLwaVd/VHLZffNZi2GBJK1fzN48HteuO
dBH9qR+t+J2mqx6QWG05TDRDX/G6ophMyoMWoE8sqCLTZ0KMmXqCer4RoxSvnpGU
+JgYT4YN17ZxT+T28d066+L11c8jisH0SR1UEijGRqota2iMTuE2n27NVjbw/rEV
JAQy0avnTViAg/v0YAc0XgnlpNDIndxjH0zTuqjuobhuPAj0ZPsdXhhK8qgoH/BF
YNVoe9+a0z9ISVxUvJiva0fU/A1JhgkvW+xo8Q2ofXtYQRSjcpC2OcuYtmrllnmK
aISqZfLts8G8iWQ0folLwFS9XdlsDbfpGjKy+Q4AIOljFwA1YggcCWvaScOP7Zsh
ztPsDN/qM810f/xv2b2ivnkUbdQlgpsW8lhrtLobteDS/9MmjgY2KgOPD6RZJY9J
xyyETArf412MkKDeCyRwDx6FgSY3AcYuy3KV3SJdgaKLWDTSFtdmlTT2foc6Eb3u
2qEpP7s9R1xzbHMrsbDNG7Lj84iIZivTo12Gc+845jOSZJe7h2x2i0PDrUW8Dpe/
+x03Gnsw/lFqQPrwcu26/A+kVhKs2kHTo91IVz0fPagukrSwHnPFVjNsriw3dPWy
mTQL9Qk3e1bhsur9/StRYxyUzitCltDTITL1kmpGlUOt7WW49Kdu/xC/57FNR6hS
9x9KKISLsoa5isNNF60cq9CTcKRcv9vhrL/wmFBvYJ5DvdkxJdb98Iu15t7DXKmi
GuQr4NyofNG7rTJo1WpI2zifLF1PQhYRhHa9DKB/y+Zuyg+iRBxwi06FArjZ3QaS
S+Wr4cJ7JzOealccwdfO+fb3wFCdUWFPjkMezH3CQJFgqS3urMNm363YmP7FCCM6
/1qd1eoWgoDjVjBiEjy9UhNewO99MXaBDv3ycs1IW1rhy6EDzybrdQ33Md2nmha5
spd6ICorOxxMyu72Pupcao+upSX9iq9xgBagHFQZAz/IgA7HYHrFcXVDmUkG6lKq
YbeLH1/h9387b9Nu2qs37Yb3Akds8LXP5LjIpiVcVGUPPJl4tZzfnB4N5V/zzKpy
iGz5k12c/g09R/kkJ9eooolkmCJYCyn1PMvFKZ861GJO5GNNF94C8OY7YlSAIvWl
/CHGCTThNdiGYHJUFrrOBPonpejZjWe0UpNyifejmUSzZqP7WkuUiQ0E4YYEOfZe
rh4I2x3ctEwZ/ZGNtgA79dxd3RxvMEpAc+mh1ZJ5BV6G6KQ/5IHKdzefWJMBO6K/
+w6zliylE6KBSVcIrH4FU9e3LPdrMOOQqhZRjuauihP4w920lwZfCHFPRWbrOdi+
DlxX0FwQ+HizGgu4wbes3IFFazaF5+7OIsG3rzzeaq5SOmY0VXDU/8UUuSlBjyjq
LLG8umK/tu1voRXbMnaco7x3garC/SqIs3bpNfVzAe21Zo6cBtqMKi2hswZ5PYzv
foYjuROBIyADK9WE3a5ozAF6oLTCEFH1anfocQ47VrXVChchlzTd0XqsWlGlCKTl
/vmSh17I2rFTJaCHdUrXbl/ZYqB5LnE44MTW6pIKXCNXKecdFp0CjhL/MUS4IYUl
leqnqFxs6bST/wXaOSAWOUZCPyKBkWwRXejOMSsD97EeAu1kal3zRmwUR3Hi7NM8
xDJBsBQltECXxOczGYLABYtjbbNvL0y/JyhAsyYnlQAFpBhb3BmxDxBYxsp/YDai
QKc2kPm2eROq2Q16B2qc44WynC+Tm8rDG2LWuSqQhhI9Vrcf9DVuryKogDkDymlo
SJixrwRsscLyvIuMAhSwZdU/GvONyFwv3NN90xhbpzSOiclGIKa+6iASMc2pgQ5i
zKHTy4/JvjMS12RpwRzERIK5xkBgJQN4l1JyyPMntBwfiA1/zyIwtsoBRB32SpYf
5gF0qpuHjoSRTH09ergnczJfDQds7CPp2k8wc0PmKW/bqcL4QyaLcRyue6Jo86V8
g8r2Emx+zNbvwQnnw7PDSA6sp3MaHeRLBWdmlmlHGgCgxVGm3+sh/rU2Wc9/HR4F
4ywlxoV9UY0pGxKLQ9RFdbMbU/fUkhmZPb0u93W+ySSq8jU+TOvyeZ6vkkTfqcON
JH+3mwEZusMflWFt5khKPXvJQF5gjLVGQnWdus8IrEoBZF/Y46y7M1UqfqpczhZp
YMQyxOSbNz4vKv6Fie3UMgbX0RZmP1pl7jmAs/1h8h83a7dBdjZNw6+ce+qPSdMv
kXqUFr3LQ394p1exqA50phP7bpEcee3ccXdDq69VtLzkjVT3zrp27NtJnS8NXgQy
XBRtpxtamo6Njp50cgwrfR74KSuQAr9LoHznNekD15rP3A6o7hN23BR9fh6RaMNv
USBP7jbT5f/xp5g7fR40Uqx26OdcnADhisU2AitbBQYMCG+cUky4j7nGkwu0NZR2
BIEnMv4ocqnGIYNLTcqVIq3weYkooatWxRrnFGgUmvlG/Kt45+B3ST+uXj8mWYuN
N8ub2rED/AEPdEVOgUn9kACcRs9ov/tc33ZmFTkOWG1HHDuaXScTr2L6cYgGczia
iBBUpC6kN5tjg4Ckv4jFvkXngV3PEfTGQ60nLcdJ/WTmsciTfUHohNdImOCux8RA
9ai2E0+33XAQn0ZrlEiWEeehEZLE7b6oknLXc/6Zug1QcHVbKJSievzV6l85xEtT
Q0JuTc5GeQc8wJB8fZgdwyaaJlKpDxxRAIzLc/gXi13pDewAZxIAT21fsPCDDP6m
oObj9yaG/nwUQpy6HRq9KGq9QlXWGd1uYxobN2F90+L8xhf51bBUeARYwEHHVOUJ
1Jx1wOnRIa0InPWUAKKLFmzp0LMlK148D6g3LMCmiBAUMdyUj0FtkPFB72j/kJAk
XdHC4UbGOF7gr5LTagIjtIuzKG6vvCUQ+GT/f10IdsglPcBgUokhRqPG7cOvYsU9
T6gmUhQIh7TZRvdkErzbHH/rBIMKXjw2r71vs/XR0NMCmCRjCWu5YnlpRbee241Y
KVRw/g2oTdimbXLf0Vs+FBdsYWbo5fcjTjkZUbcLc9JpcRt9iKrq4lM4ZQszf+p/
w6lZtNHRLKnOzD6RnrxlXncZD+xC18BE6AmArRaUMlq1/KF/2dK3Gg39JAn+cN0Y
xG/k9B0YpZ9Nep8/O4oQvMMPFt6dE1YOoWKPK6zTytx3z9k7Wrkx4OADZblLmAOt
rMncuHuQhMcgVNqHT84HtnHtqcbrWAjfxMcrY2F7e2LYEAFl5qrkrtYpI+oWDCk4
LZLpZg6HzMibDx76T9ovEYJTYl5SelC250Q9iUFyazbbzws6PXFOPqhuqZEabPuq
7oGfV5AQAXSJFE8/jbu1oxvZ5SxUqhDu798nDGYw+gkxkYbbawfB1EGQyImtibir
x9qTbC/Rj0sVo2VHr6wDwD7ux7WLib/niFzqkhHnudqmQP5lpRrZ7x0tQPpwaMZt
pSTEcyj59nSz+pVtjYOmqFxJoAb908wmY9NaMFlhRfkNL66o/0UB55jZoJ4uTtv5
nqySKH/HC69r3wJzjeJmOyXioKSBCnpG3Ij9c1j068syDotpPy9DwgfxtYObHrOt
HTwoc0Kzu90Rm249B8a2Vx5CbVV/YzBZhFxS9TKTHl64vc2FhqPX6wkUYqtmG/am
0oinjCedEsROZ1x3HAlPjEbPhZPmDbFViH8cFa9VjsImxucLOEM5F1oLRXSeSJLq
E8Zs+0kx50l4V+6ahx9vqFQeaxUHgnukytJKDJx2pHdMMSh9pLva9Qc1xfD9+WvL
OdvzwXOoTAs+cGETEWni7p7qhj27uC3iV2c6i65PjEd7rscCztuEfsqPSLq0DzBi
qoio5+jsff/ZyTvHnQoswzder1HXHiWgCyf+iHg5AEA9+SbpkiiCbAjG/0ECcbR1
AFKqayv6VupTjQivD3sGi/6Soxi9J3twYjo1pYQozB1sQ1lQ6wLlf5XMaGuQA46D
bHC0mQUxCT9miUKF+gwPqUU3kFVWxnQ/RoQpc/em5mnJI036qqAFtVE/kygUyoxA
aK3K1Z4ZZ9YEfYVG4eMySSRLBcSpQo2Fvtt6DTkH9wcIpLE4goCWGtTl/102+zPn
2BKtH3UStLY8elu00L2vMCNe6nOTZGu6a5flfg6abpOPpvUYLj18dPw26F/uIZbs
j7L1WltHVL+tQx1hQBGRVnywrlNlHNcfXS2lVJlqrQ6NUu+m09u/oOPzF17rFj9e
IPbhCIHXyIyijejEidYwufT2sWwssfEJn04YftWIzqzciukRmV4m4Fk6X3wVTCUI
SjZro0YMzjMQ/bPfBEdU3vST/FVnqUvBbVFq2toMTvcsMttdJr8N6Tg7NTlwlQWY
nbaKnYhydCur4roT7XPIuN2imTY8JB36OX3+7DjwDtRo6aIHNKIntvFKdL0QHErK
y6W4RecZgEw8xCLI/P7KEE/VNPtB2lqOgyv6A77wuVkv87C5S9o7hcR4CsbNWXFZ
axZEazDo4nsEBHpZT1tMCyYUpDxcvFeOl4h+J5qMBU+PzuANLoOyJ+T76VxCXQqU
QNpSfDM8nmDg+Lfd3Vx5eRZDA11XimWEcJ2tRDwh4G+SudgtZtRwIUym0JE3qin9
j0weFGE59LJ3GZdZNvznzyG+ifEbfbTJaE7MuAE83pyWTWoDAqqZ0u04X4FYBbNv
OTdR0lPR9EGXGXE5mBotmfHoDZzKsTN3uTAUT5b+dk69ShVVitqdetNtKbSMI693
zNCncMW9nSTCZKHEnvMOGepZ41Eh8W8sgbZzC8W87q5tAiue3AJwGz2Jd2PPgv3j
nX1GJ7ennzMQjqnfcQljx4mhwO4pczOh159JclnlCbiZAb9wXVMFKNEHWjBzq3cW
oRcC5zo+4u5fpp2nnvtGltkXoXjPBNFyMTiFfue3rIdA6U5VLUQ21Ymb0TAj1KVt
vgaFhAKOLqaRhkUhyADjicAEBo9Gw7xe+mAxV3g1mCcgaT78JJN7K6Q3DhZNp+AT
vkJ7O3IkIhUe/dg8nfB1Dorud7Bq5Hgy1gxTJm/+FXPYw532DAK78+HvHL/Lh130
FpBP3G8s+WP3gQDCkrjpCFWRN5piBcyywI8WRyGs4m3iYXzkKVLvP/1uP9NPjvnf
gAnhVk/Gu9G9MxmOl8eBeoGni9v90n3usnVCdBs7N5j6xMmsg0wsfDas02VgWzpB
sSKnBlzmiSSnswVKi7vVdW40NAsw930P0Gv2U9G19MsqLC5K6h4bIYuG4baufqBo
b9ag0h9HRGLQ1osASb0eAeYKgHw2OJMSgblWhb5NWCKebBBHYFk+VKcgqelbtjvo
wjnjNnrn/ORwXERCdIWwjuMgAJYY17XjYjCxWoRN0TMIIv3ltjCYpJpCbJ4QjHzR
CVt2OE+5n1q+mIq7GwYIlLUqkmpKS4PSMw1WfwtDelZgZpGOEeBHLt0NoyQsZXaE
xD/a9SoOW6H99JFnHGxGd5aPaR6QkH3WMFLbrP+HeGkLcpqXi0j1VnSo3d+XIA6B
4ZXW7rM3T/ftuqgAneZVeUzXP58hQLyqr91AqvGihdAH5HzpQQf02qA82xWXltrY
Q2USTgu3OzQQF/lK+dyGKIZfg7eRQbRVg85jgGoo4A5YQW2e8yQ9m1ErVIsPBydh
qcVZGFSQVYvJSm2pRsfo9risoPYmWrG6BRhx8YZZ0fcDySNS9e/T9Eal/UTyo9Hv
Ef9uP6UPy8rRPJwjLsrziQDbD5nXyyMjnUTaJCI6jyjSgQZW5M8uycTQc5Xupbi6
ANdEVSskC5JPLlwtHyTLVHqGT8NbmQKCDLCDF0asHn7eeg0pIth1BSWzEt0rY6iK
TLqK/4KVhQ31MVipe5PE4DfSpzIQk4gjmCCiWzbh+7f3u+nE1cbYDDItsUGF1F1r
M6csCiAqEmJOXWEGFV7VyOt1O9b+aoz9ncQtlGUgDFMmSGIUgLsDIBInem3tbuFy
Y0A1luqpAMkS1P6WahDQvtauCZgkbSRJjq9Q3wzDK9X99gPq/2U74yRRgl1DjYMw
auWEplp4+OqfC0M9V5ykjP3Qbqz0+7RKEVWzBNFAqXcNQimtrc5tOk0Kts5Hq1mv
u1aI+/wvJR1p2msDyMGv7WoQwKcoWP0b9w1RANGEPDn6B0gbiVTIJiBADpI+dCHT
DTd28BntYHKiRMGSIozc4nuoY8zkZlzqDHgBoV3nZ7wpr85Fm5ZXYVH7QZOCq1kG
Z8DGheLAl7vpUuykGo3GXLeef6JwgeoIZTnXba+Y9g7HKwF/5H08pBc/t56lK2CW
31QXmL81l9fLMn5XCbO456dYjvSjpv08yzZBu8c/sv6gJsRSLl7ZCtDONdcqQeel
io8gD2n70XsOAWhChOm8GU2CyyU/PN+Qe0EwbuHbFuNsexAVt4JPvJtFagxx/ecZ
tJ5gmefUB7CAEN6JZmWQtTiVQOAEEaSed/KojcUyJhVof4yYiLdk041drf8SYeOz
HuEc8jcnLTKcfd5sCJh3OZ2iy9pyGZPvFtSiw5OUcHrosFjtY7/vYa7cJev4cyKX
msBRqiXqRt0TzOPMzLJr7hS323OiwAynoEoP+lmw/fD5Ko/iXu682FfYih6tHEja
ND+pYwcOOmcNvbArA8U5gqGXtj/wzWSdo2REXODj72mDR4r1ol5RlxDBmAVuIJIi
/AjRVjTr0sZsuZ0GMCxj7G8WgTBiFMT/KmgHmB9SUqEnAerbTtl6GWYIsq/H01az
wgm2IgPitCPHa+0Ch1Ve8zz6d+ULeQW7lS8rfBZt4ogSRoQ5PcQtk4rYrgAPUUU+
u2fQQG7TdJ9XP9esOcqogEmsljQVxOMKGeT6BNnWFB66RQ2Y6sh0VsleEijueSyo
KHAPgso5G8JXsBTcqmi71acwrY4JYhtJZeEw1pDusyNehY8j6aGpHTsu1Loectc7
Ha51GCEHAT9hynY8zFS/Z1gJVrttkqLjYYZI5R4z4qPzB7mC+4vxH9AjLxxfMQV9
xhgAXnmdDBab4v//nlGBiZqJdZ2esGqxVCRUySyLQR16lGsETK91oZi7JtfLD/JM
yLM/jcuGycQWvUwp+5fG2V6b9XLmpzHjNNWEvTdMQjCdWZt2I/T+RYbBMEsuDdtd
a0Kljx9L1tG5ByS33Qvpc5gX9F53mFDCCO4udAhfWi2zk1B0MArvVRZe2ht5WkGX
LdzmzBUZDTLw2vrEAa5Jq4CBXEZ+rrxGkkPPuOpOKIHhsrZnL6U1F1rDOWgGTsZO
Ir6ytSvmS/YrwhFCSLiMjlSo9Lcohw4P19e9QG6+z99XN8bQ3vprKpE0kxTYQgTO
1CW4R7B7jc0pmNwdQ1L5kAVWGsy1LvIkazPBRjY2bi9BDoqLcl3Vzj1cZZ2IR79H
2quL6bsyN5lr0SZjNqUjnN+5n6Flca/ieBqHFb0mSZogT96qvXvMrlcuVqyRaTZ0
3kwTF8WPrH9Lbp6Z7qXubL8afeXwyXSFFIfZHWjpMtfxpdLbValextcMw3G7+rRp
e3VqE2mrNrOHLbllPxIASSQqH3h4xuhj8erCZo8sSGUhMYx3lRSB0upLENsA4Ttv
8wBRogQhiHqeBMlhLUmR5X0ss4erJ6m5BB/Gg5uPdX14HxMNYhZwfqg765L6zkfl
JJBbMoLp7rePxH3KfrkKDmBJvSZLfCqHZ63fT5HS3ydmeupVfvETgQJuOtmfOsux
mKYceQB2rws7dTV8OMq0daNJJtu/UhOs/yBnul+jdkc4O07RoUA7Xxl0Bh9i+uI+
nW+xEtyurMcWuTap96r14xocYPCIXYfVhUQLOMhxSGrvqm/UY1q3kCq1pn4uks85
4mPOTmTxZcHWudJxl6FyZIewY5OTUIHE9wnivJdPTpxnsrD1AbNfzlF0UKQjiJiM
YMARF9lJMpILgtt9Ax+ZLHVK96QwucUU0sFDrRHjnZJIUfjO0ivVX/xr1RrkpgGk
qNLYbEaceVMAZ6v8RM/ftMjGZ94mVenMVU2Ux0nBHn85OuU6Lgibk4Z6G3OTUTvF
+/OOirecEwnBPYFzyV88IhT61KHf3dy8BSd0GqVaPnUfJqBoEMZSxOhS5dtfV5Gr
AXFosNuT2C9jK3BkmwpGsVAavooX2Bk+men0sdvZgQ/lqYcwwLnBlLCCl/vYvN/U
i62PzLlCs3Px9ct+W6/OJ6xwB7uAMjU+t6P9zM9Id/riSE9QcyaifqpQ6s/petP4
sG/9b8FCaIcI7u4iX6MagZdWvTlsv9n/LpcSAz1YG4kI0WXkT/rS5Lo13PRVvKXY
OuOpOw4ZUjCC7MwBxQnfMe7twz5X76JEeXDneD9h7eLqODY0yOC4WBYICEs8+zN4
o4A4XMJ4QHygA3ADIgh+my38XcDmpgppAwCNTkJh+MCtHH1SHp6/HsuJY8k4q3fC
L4a5PaqI3XU31vfJ5FhqMrnG/QrRV33jfZJj/Pmu9ODrRQIJ5ApWW/ygIEwx8SF/
YY5zkIevALycapDoWupWRAaQMd1gxJ9fM3oSfp0nMYOuyLdHwkSsmdmq/xNNZYtl
81Ws9hE8TJ5q4+e5XMmLRbcCRK6wbzfDJI9hDcwRtAki0bywlFZ/dgCjmr3GDWD/
sRDKlc1J91Nu8YgbvUbLxy+/NgliCTQwozEsT1yJtn+KXqhuZqZpBZnezkGBowh4
bLsVDaJkpYqR2PJshVkpYtIxKw8LOKZLXo2gL852Nt3vKeaZpBct/QRv/sQNyidT
Q+GbYdmokPL4zgtm2CktcCTrOPDpqYWRKGNcYEGz0o2jtQTjNsk+QoPex8RQ4bI0
gsGMaQI9DqPpXkotzKH3IU+FDaWY5sqSj3p6XjiBtNS0unI/wsK2myK0sLTdWkC1
bQHlk1BLIByNHzJzlp1BQlIwWUzP2z4Kq49CmzP4qBDL6QmT571Y2nCHFxZzTUjj
5RoFdkhiUy/YPBawrjt8+DMvuWgtfu6oOU7d7+nTUB0wklUeF7UQMxAimnDBMP2P
bDYKibSB/HxLqRud9R0JC3qMnmvVtlDglXE2M3HR3F+bKPAJSljnQAwnkJ3j1qQJ
3hWT5nWXKwms97NHZlPJVWM1mN5JYAkbOw5LiDigRiOuDUA0AMAMxjpx4gmQIWEU
pbaQH3dtk9iDcfRaF5Q1Wp8BkR5x/bTFgGKCj6zNKduBey0Fyyb1Gg9SuQh8XED3
1WGgZmDMnICet6srbH7vjY0TdDv5nkSG03uX15TYBre+4QLqyB+9jfUoA7P60Rdd
O6z9AR2zLSov17EKs9HfhSAERJhjZ+S+EzTg4BnqatWld5Bou7kuUKVHd0xWhHyj
b9kQt9OwmSqgiV9HOZxi0yzSo2FrJnr53Wlo1BEE5N/tDeaC/oJncjEntrrMo46e
Ov5eqYspTmjrEWHd22QFFZdf7+fHwDvmXrfRbPg8vOE8oiN6k3o0A/hJw95xfm4y
yKYo+sWL5puFjc6/9XmE5oFD0h3i7+YZDnqn1LqRon4tFEmMucgAJiUHdZfyiadj
JU2h0aKgNkiKFqyTB6BDI7d+pzvaMiMeT00z+E8pZaMq49yCsSMfIE3CZZHtBxFY
HFZ4BZ1HweFRWlOn5UKODLpte85764cMMY/6eIpJFVtkLwfVh7Kydnr6brfTFXEk
a1LRVJQcqGM/H5gsMi+On+4NYDP67xgpYU6Lm9Hnzm1bNcj9Pg7YQrMQeVM7ECgI
4+dmk4freRYkIcB1p5m1wbyrEh5H0SWvMgZ/g4dhvYWOhdcq69mBhwrI2VNyBZEE
+2aKKvSD15AUIJvh0Eur7h/UVZfkTqiDP4SFLEzo6P5g7WTIxpZbg/VG8tl/wcim
JYJejOI+z5CWzIbMPoUWbEdLUN26BeNqsM4DsqC6IvKOEThlzMu0xULuzKESjE58
qbWMt7p0WmUAe43PeGLFLltqOjuA93ZwVCB8wS6DILoT3z43Yp90SlnzCz7Afpou
UQmtr0Gd5tCDE6AT9e7gSkoL7xlw71fHFNmraXuqlH0dqEy71lbpAqWkiosA7aR1
fN1L1eGWec90mNFfTzfd/pHYz62jJkJ+6ETbsT4a6OU5WQYil1EO3iM7dAItbzH1
JHe8zvMMYJfKz1MhBi7BIQnGL4YvOODd5iJq+VHm/09R5FsSY8ZpDsRkmWRPc8EE
Sn1nta11JQw2jdD4N+ym8IS5VHMweSyyulcEr/mtIB+0CirdOteIHANgt3Rxvtq6
WgoQQsNEOOY6hBWccGefW/cCzB4pVWCB4sMePeDbHoahirvjw0U10x0zFacokdfN
PoGSpmmCfCMU8oft//smjH8R4nYWdzBhJij8nawdztIfnmfihDnMrP8Sx0LR1NnV
ZDDEala0/k8FBV/zZtLEKNOFR/Bq6ts6U/+gnGy0/2P0kuyg6ZRcHWLZaCtjRvQF
/7dZw2qv9brsxczFaU5y73jgOtkFniBPagMJpbuI2XVbBzQwOKremv5dyZdgHs4M
n3GD1Lj9CUm05X9KZTCU3xFrl2lLTuX617y/1UrxVkrZETAhrwiQmtg/8OZTls1D
OhMu9b7/LQVxbcpqKc0+y34iltzjAmKOe6RJlWI2klLNV1o8lba6fdV8rATtPIUi
Z501Kib/Aml06y0y9LaQoOe/V+oGnUI7DiuNkR7uAWPX/Du8Ww8FTfrBIDmMWxmM
3aR6KoeaOtbelFyJPbRHHoMRhvbO+qeu5MVRFKMEO/fQULxuJECC8FpeWWInQTZq
TUEaNvvBYkZ0FqHIo3nO7t5WzX0GX7JV7eEZEIBgZgUBrHctxTRpxiitN9060l4K
sVwqV9fKT3R6ZLDr0F7g8y0OPx9YE4/6WGcAB84cibxFPXZAyE7R2wBtIGntTHdh
Ut1492tJCEdyQnp8EDDK/L4thDfzpJC4RFWSUShCRrzb5Gqa+pks5EKxyFgG4pSK
7SPwP8p1jxHiWxVmnLa/eJGyCuDY4fYXRO2F3W6CHuVYWrqWWNgZaIWOOgoCc4gu
whiTO9rXsKOoOLo9e4AcrBeKXHvmwKoln+NesDTZNUGxvCqpvl3DFyjH/MNPfEgy
IJROBW9unoDmYNdWXHCQ9rf5N2k3lx+VXVK86gOXSeqg52v1f8qFTDH8rxyeFqQn
EPi2/6NzjGNKNmNLxQK8R2LHskvqAxJTA+FY9f8/HFUhfHqi500QWEZW+9RdAOAX
1UVZ7J+H3eHqdrChngmLOxBYxe9C6VlJ/8yjW7Y0ha76ywHihLgpRG4LCd1FFLLu
TrSVeXSgsjafiYYFBYsm7MCg0lqLCY3OZGrswTnvi0pG1uSCdGIjqiBEuxFcCE/B
+eGo0rkb0KkLpHqt4PjYHRjzmNXzwMRLd4fsknq7GdE3Mkmknj0coMfsCpN6IJn7
g79u4ijofhw6OUEzTFq8C4DwiugESJlZrw1QeZu11KdGho4lKX9uW6cSMU0kcqUZ
eFXxo21Pmyig6ITmpeei93O7hpufvBfqRUBC/Tky+nJ7t7lYY403ei68fCEEJWrf
ObWZd4wbdqttE54hSAC1lla+tGIar2qmrMTVNrbFc/KmpofgSHmWWK2EKqujjBUp
dA/a1dK8O8ifcyfMZWh5ktJxPRXXT1crcATyyNWtC1WzcXa3VBTo2HGrZ/uK+DVU
AJtsIks9d5dxS/KqlmjKNY+h5eMV7mgV5BeZcZryVL5Znlr4aboBeOf8DzUxOczq
BooT4N1d2fEHv+nKbuhgSS8rqwU93WJP/fZkaJgs5WQFQQE5ByVEq0lI9VtUvERl
6SEIT641akioQIFAbAjyHJk3A5XLuAxMH+U/ayZBu07MSZ8na3g2+I3c9Z5IuFsw
COsXJv13SUBxPaE2cYnUh2Hb0HesKTw39PZqiU23MvI=
`pragma protect end_protected
