// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:02:11 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
UVJmTOJK+83sjGmHvIg6GQGqMrV8qWoTYR8ONm+1gtY40aV4PSd7CUbuDLLfdnOt
f/cFZYIyV/dEMyINooF3ZLa2+6eEbaxrMMfXAkZZZusytY/xkMHNJa5ovWFhIuAw
V6Ku5TPpJuHy4U+pB2Aa8ZvVInN3GBPJGrrVFnCVmBA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7088)
XpKgRwWSQmbF136qMOTVzOY/vwjKRSfKU7tJNlVUQW5HuKI++ufRnh+6o6CcLDeK
6OnvFKEqinTOQo3UP9WiRase29pcKN1b5nm2fXigUmR8QeI4UYAQIbkW/9RRcnll
j5z1WRELRexuw/Zg8GptP2RutU46CofgwMTWWjyYvhq2nf9ATxr3n/irnNY6dIKu
hdTcrObN0Q24EdGds4++6D0jELTmnG/ttwN+mU2AAQxWY7OC/SZbnRxQiTFRaXwW
UquwydMV63hnvoK8AHjfV3LxsAfbnnTcQfwIuUdEz4GZ/oHMudDMMhDr2eHk08j6
gIICf+//79lyeecp7tgQLpd4hoTclqwIlNkrqThNG0YEQZXdZb7++JuFUwBEYNG7
RbN4argPoTy8CqiqIQI9J0y4xH0pe0LLWCBKugIEPkuovi19xDZ8RpsZxLAHG2ND
9jJroNu3a8a1sUhz1lSTZCJgQFtoXLbUq7DtHy80CpWxusSBsM6dwdbqpDT75NP8
xj4BMpmIweN3u2Ld1JDpFhw30lI7WmTg9f3moixTTboa6jBua7Blz+g+H2LWsz4t
h3ZVOqou50QIHy7bppRE1YYPcIQxzs5GwXfJNJVdwZwFPjwgnlLn7MDSf4hOO4p/
06ShFSltBTySTPOYfQ39zxlp3DZSyxPZXcfw+NDtxJQbcV81cMWWjvQB5R/nAoM3
Op7wFUgjGoQ1IwjUMrRkbvUgjMFuXFDGoQqrb60NiwMrAeWOR3f6NnY0h9dSt1lI
YeCIeyFo9r6l5QZYiJbRTlC0mIEMCu72l48fpEMxRLQj9iuOsomDXvWp1tliIDci
wOGJi+LYySFfhQtGnRfRfv0u4TWB8OnHlhKgbxiQIyGr/XDAOtGdRNGygZyjp19B
jFICz/1BjzVCpgyiMX/do1S3tOfXQnr7ffAn07exB5VCxP5lIPB5LAoKFK8xnueE
XCauJdroSarXJiLlRdF/MCc4jLb0VAFb7Yb+A6QqTMrGeKrT65CMi2/hkqAl8/Nj
9gknEa9vtB79Vl8Dbgzm4g0+RK7rgXd6DDwtF72w8hE4o0V7ofDqYCmrNqii+KeY
mxX1xPiePMhsr0P4QgzPrpYrscnxr0Mov8e+tz54ZEnBH3UhznCZrUcgcAW6Slfl
S1X4RC/9+AnqCd/Ok48AnRx6vyTpG+z0t5G0SlMeIFU0ieQCv26w/qr07/GmCyMt
yFc1TfBKAQ2y9y0YkCkXCys+L/Fr6Lj6TP1eKXxS0ajbaYYlq35DEvjU7M3II3M6
j3syfEmSYFB1MQ75AOgFqRxJvDXSwSIgpA6AxkAh9EMtmpdP4D1sU5VHchVGEXqU
XTtY1IlzcPGJTKuJBEVW5rbIcntRzprbV/EwlxleWoORq4234wed6iwBuCUOiFeO
BgWBj1dgEt6fAwOOjTniw1XezYbQvl13jZGXyqKHKtEmDqcliAPI3zIFv24hu6cf
zSe+DrE0ya2kCoRlREVewuO+C3eIWfWuEAGD9RuVfXva8AVxlWB9uI1XC+G619rj
265etlNIdx0Axt6dhx6THcpIoH4ORGtRfndzQOLcy+/T5DC+vqy5owsH23QUSRea
Xmj2J0Hco1OziahFgJOL/rEMqu60xrfcF9rUYcfQcqYCqo1SAYTRnY7ymBYWoxzF
Vkcw1jyLGFZ6vVE86r4NmNg3FCK9viYeWJbGE7P7a+M8U96UQZ+vaqMGyUaVRqxW
6Q7oP5Er95KT0fyiqbvFbEt74QxHHa36e3Z3PinyjKWIxRsh+3neri9ltXXdFDYY
BfR/V1KoCPbgGKkNc/8OkeuysE4UkWNt7752o2NvagPZl4vsxoo2PTMWpYG9qgzT
hV+g+GXwW+WAxxWJyl6XI9yrM68mYTjtp/+3QwfwpD6xynMABAeOvRV23F/JP+bs
i8xS4J3xzCskdWyT6qc0aDjnLlJTPQHqjWTqXNX2k0TFf3a4ksBBdElyC7hQXEXI
NB49kGVR3D21HcvMBSP/ju1yhFcghFhQuyGGEMPNeuJYVxE66s9Pd6jU1O7U4pj0
VidmgMiUtLP5RGLjbkPPx1ud2SC1U66kPbXmtktkdikGwVZhD+lZJdjaoKuY2W0v
5ndlJ7AVyeHSaLyMlOad/VdY5pOIeRijk1PqIsQHlYDmmStbiLXcO8hnESUXS+PK
2F4+c4ESjtORytRMJWSPSNWXEGLwGCvj9pR3hquloPwQ/49XISayjNQnWLXbiIVL
tdJVLOKha27ALkxd1tniAGRNsqkmIxVwg3H+/F4CNIVoGGN9hZXo2CjXXRs6X813
IvPe5rQ1ipNpc+cJXGKZhajdI2XwUXipblZYR35zAP1PecTY5IqAGAZ26hO+68ym
tWYm+SKXkQs2fUl5dh6B2KWppiibzu5OCzAZtyG4fNfBQpDoYHmloCDN5CFqOzov
LYpm3fTUXmxyM0Vti2psWsI4DkTwWnp1lso5FiUL2LUxP4ownE3T7298HZd+PHMq
ROuJtE+EiigY4+Cf7i9rlK2Kq0mkJD7Nbdiz4cxJqPuc9Ta9eil8KDJSlBsmBp8M
aKJaT2/Ivje/mykm4b8p827qinDpVcAaptDPhNZbPawjhfNX093EgeH7mIz38Avy
wxg00nWwLribU5bnhs/ib3OhArB3Pl/XRgYEo207SDiFRthiEkPaBB8yT72IiqxB
jzw2e1XT3jVHYC9hWbJid4aR9Aro18FzOTjpKzJiRag6+l6Gw8TFXjFMabGBZEaj
WtIAc7z/Jc7MzB9uaZEgbVyGZc0+VpgOp8ElwaKrGEIerMEc2rwplw3Gtu4aT7/W
XopYCCgTeUW2CqCtDZMchczvJFVB9i3Lb6W0v4BZaobGZ/OczPP++aLwotOgGocA
BMmBdXPWbC8umru9HW7xxsQPfs+opsJFxWUKeMaPXSGgzsGKT69QZsS/ra6GtqKT
cgjmZO4ACeYYHv/Mua6TMXxYYCSbn+0nqdTh+3vWc5xk9yeDbPBJOLUSwy4Upu85
2yzSmcVFXQkwkAV7JONrcBN8Wx0ZMj+Vhh6yb+bfC1VeKdGUg3yOIgC8iNxQ90Xa
sxd5BT6hy4SvJhHsqF0hdg/vP1ogjw9+lCBDZZIghTNZ6Z4FZYgRNJPK3hhK0KB4
r3pSyGUdAnml5ZsnRIjyopp05USqAcrB2jOOTLOlrpmH2HUu+3pqYZ75BpekwxS3
iuF8/ptZ+TIOldBWDLrng4jyNLZRnIgrG3y5rWWyjY4N2JKEa/NYC31i+9cioSXK
EB09Pc1g8UqP1xyB4QF4+QJdsjN6w9FEeW2wDE1FiI2f0hVkh3j7VBsFXFn4YKHt
POHsPqWhGwEMKO0S/UmjzT/qPMGKnHU4ELxabX1Td6OvtsTX7w79q14nP9Wlba/1
XY+05IzdJ85N7wYfLyZignvIoZ4kuanWDgmgFqybX9hRFyZwoQsPfMkTKpJcjnbR
KEo9ofipqX9Pa0BtYpc6CszfxK4Df9s6N7zvuSuDhmLB9H6PGKQFILEzPpTyE2cF
j4XOvbDd+gebkmgSY6JX9ABtCEWNHPEEeOP3x7JgVyWIKmCPRnqYoYRdj5fU0q3/
szZzMvHYEFWNt82S1SSXAypMOmRZtSBBl/KEsB+z8GHQwsM2WWZWw0oMh7tdroz9
k5XpC6n3XRyHgSYlTWHzRw1f3c4T62WZY8jv+Fy7RNb8adnSv/FoTL3cgiAy7OKu
jZsG/Ftc7ope/qQrTolO+XgOR4wzcCe4XoYsCuAT4aFelRT66TsaBmVZIqtv0uSn
Y+mRg53WU0QkFgx6BAK3ob4RUPyMd2hXnYIuGVhOAjyfsI0C5IK2wy+mtwszjL2G
vsrSjjzchREOb0oLqToEl3tcTJnwfON4rKWwVdZT8DwSaRZvhOetzYwmWM4ssa8P
OUiGWm6imu8am03CrGBoCUa6W1iWW5J7hY0Qumvk0Wg22R1qJxjiMY+rU+dZ5iQB
iXpfXFUxWJa5A+ieTw5F3TdV3L1C2we890Al0+SVcdjbSLADHYDWmoWf9Zc+Z6ka
Ikg43ToLm2H3R8qgn8KkvohQms6r1nICeKH3uIjTBPuFpJlvpEIWsvD2KMrH+5ET
dk06Kt23L9o3qPHrQml2wUmyNA6Jv9+1wyYCjOOCdmaHO9rh1L+aHQAC/2Ls7U8L
8LhxlSSnGETvC/4qcHOvQuygMu7Zh0KlHLfM1j1dxbB4T0BUquBDHeTpa8bIl5q7
49h0cc+tbziksVrXANU4a92ds5SWG5qpXH1746FRPPIFJ42xzlUoRf22cTGOqTwu
JjJQmeFJOR+uX/dpOT2nRXFQnGHJN2BGmgERkvFXvQNXxrSgiLik30B2PFHMUVWl
Opz9KKO4U5tWwPUF07Pl86oEXHLJKbbYvwRI7U3g42Nstb9dGHlzZIcYieFWCImP
g/hGpXGxqYB9L4furmnDbDd+G1wocgP2TPbxHjpfd0NPsD6UKDCeS1ZHzeQwPuOW
uGTt2gwax35KKEz6w6P+TQTCI1oFNGvnntpSu6gHna6SV+ms6GYDZEvACUFz1F43
i4yxqAM0k0lzhY3rlHUR5ywZYmGQbRGb+yJ/732Gp80hhOrJ/J0Ne3gFjIfmvGF9
9svJbx9Dgun+dW9IzXZDgXq2IFWd7n4gK781iOz4nF0rDHIN0SzeiDtKv0Fa5rfH
7KMpo5UlfKjc5g82RbVclz/Aj3yGT/DKCWYZ9ldUmpMhaW3XjwxtPjVhKDuXf1wO
J5MXYkv0Nnl/wpa0Tc/+9Hsk3elcBkpEGrLwtnAJ8BBqkC2A7HRKYg5SWAkLm1Bs
0wAcbXxBv9ACbMh3rNTRcXXPyGrLk7Bkbd0Ix/XhDrAu4197eFwVXflXeigO2MNO
VHIclVdc4gtY9ZfhYW2Isy+jSjIroBPVFoi3nxHeGnSQ4zy3vfrN007k7+ew22Mx
Txz6ZcIrPcLZeaFuPEU3XIwvHBt5BdvS4XsvplqotX2N3LhC47TKusrFBQ867l6x
ecRW4WKf2bqZB3n1NBQ3UC6XpKmA6MWwn4CVRFkW1jlju7qJ7vKXgwMS5TJPSgyD
t5YiuJhN7KeKj9x30EN/zCPeTMhSEGENZKPdL4yWUBbJTCzRBjNIq8TzArIWnXqU
KNot7ezkO1Gq1xlGvEb8puwWGWmXRufAqVndL3MpVBUL3/DYu6AlO88cJ8svP+3e
apEQJW1vv+laQcxShEGBpAi0bhaA9FVzPep3srdGfAJBeSS6oepvfCmQsqPU3MYQ
3ZmJly3NVcdPltkkwIMgUzxbi1ZKmuxL/AnwlhG+qRvTCdRwjkVhEMhCj7L3TIyg
Zc2R8iqWeSUyumkXWFv4A59fjjCF43IfURXVwKFNavfYI0cUMoyJb8BBpHzbVI48
8hh4MhJfOn0E6fQDw4I+0H02YpjT6w8udDdOwG2XB/cCFPn87z4yjQFaqkXgNz2M
7XqdOj5REsX2pSmoC6zmbciusjCeLpax7wmos1i/DMitMHFa206AbWJBWlCuik5B
QQqfXQufB2m4jTSdcFCoVYKHOQ72UDEpmmDLmGGisHvTLx7qMUgqGJawDZdJJKiO
RQwzvrTRpmy6fnbmNoQui4xLdfsViJChhUkH2Fqq0N7OOo60IetEc+SIohWQrM7j
hDE8P0iobot+maQskNkkS/VGJvdCasjMowmEFjS4TTrhgQgBQ3Yi9HT4HBtN8xPc
/ZLH1T3PzSXl8idElkkVYpLGnKS2I39O5+MiGBkU+e3V7EiHAbeVjg09ZtHY/FMK
LgPYC3FhldUXr7QxIyX7ZU58ikMOB2LHf17oSozQbKQuxgiqijiuTc9XGruiEWCx
iJbvtaTQzhBoFhkZf0rCODXWXj2DBATCfmKwgMIHjVJGWduDzAco0On1SFLv9uhl
7vIW9QdKaGJnzXMrUYFxboKZE67l7NTBu6cutZt8ntEfRnECq+qyLB4YuyQzpbvR
TnhxLuDaghuIbobC+XFpom2vzrcIx8u4n6L5xBI3QFQTy9TyuhzWGczxDlBj1+v2
gRAy+hFmRs58UXTJVbXT6/WvUXP6TAUPvudRu+IZ3WmgJjRuA6NMhUsP80Sg04ps
GIQvAnX/PP4xp2wAzVFn5S1UKRv40zWb09hXSiCextMn4kRDw5kgXeTGB1Wk1Q9A
7msszvSf6VLZEKlSiCjrQLXK7vYlr6vuYpthWrTZe7VA9qtPxTLnEReSX12MTij3
7scXB5is94qwppsqZOdoJtidUy4sCi2JTrh1k4nvqfQownNKX2Yhn6ZPid/VqtLH
jDLwyFOmpLb5Iw7sBs687PWZ4uIbBktV9uk3EzWUq795Z/k1AWgS65pBTqo3AoNt
KmPaYBv2ZnCvCy1LdureBTcmcZOFHg+EJ1p64yjw7KWo6xIdqxvDz3sdW/xiaH66
hH1pGKHOGKT+XHD8atTk68CC3/GarSb16nMLjtcIvpu9btGP5Jhk/gsPSdQ/clO8
yg4OLhvxHmUydB0SrBESgrJQoWyeVcixrcTGOQCVkgMMwkcRg3ixsw9MQXoa9b54
OIurSHflBfeNSCOyeocrMn+JrY6tK39lkF0FTl0Efev/X/mBKhYUtku+JW9VhJ9W
zFJZAGn41ioe+X/Ku7P6E/MmYayb0d7fNQLtWeaCG96oh15pdIp98a2ClPFLLEtN
DMS4tPi1p6O01iHEY/4fs+5Jl00/hxMBp63x6YItpx2HXTRXm2bwLzFOb64jLQjZ
xomRvQC3tXZQc73QGw9dOW098Zn9jI1CXCJVbJLb9Cg8+5qDUK1LAN/BBPnUeBy0
xbd8t5g1ZLZiOJvzTxyqO9whxyO3yyatDUf7qo0CZI/PWyu2Ot06YkvisZhvw4nO
PgFCw1NeYa+vI9+a0XgNGcszEM2cCYATM8wzIu3PMwy7iHPm6m4krO3GViv4/F77
0rViFnFmXS48pNoaHUo/GnKlnxVz0uOwZjP7OTd8afXgyx3jZogeO6AUg5byXtgk
ILHyoAm1kiHOkVW9vLwI4Xlo3+TwpzcEQFrVIOxi5FPbO2xzQ+GfzqPb8pACq6G8
5SVN58LR/dmjdb7b2T4H0856LMswe5IuR80eUCPZpZYEUWNfFSKp299NuuRjvRHg
ymx7rzhB1ptEMepAb5Setn9OnY3ush21fwmhjGXkwKwPx+nB5Z0JQTpCm6SjT6Zo
iUn6V9anNSdiDcgFHFIpxVw9XJl026tehQjGbs0y3PKa7btxOXZkOuCAdr5CcgRG
BSc09wBm8rmcz2sAnDc+9aQaoQNc6ZDYVKGXG9C/dmGUTsYa6dPaR5I018eZO+jZ
pYSFOO6/z+VU9uDUhbve59J0kIA17c6mswT3p22ZDGNKHBL5Fc2RRs4HyGzK+6VX
J+7yJwFSPgGXakVhSmo2v3cwKl88x5HgehFR51AEDXatHbidWKGgE8yTk2pQWo5F
tR7rPYW9Hzy1CAQerZxpG5MAGFZPo5zDtYVPpc/MOTCxnCDNl0lPEMNf5IxXzqEo
1FaVpHXxEtCgem2DsnhG4v8eBKYZL4wpFbwus32g7Y3idqZrVGgsfk7MuviINTGY
uX8XgmrhF5xLlCdsIp4aS5h7rVbrH/4VmJ79y8gfSuHcDs+d1hZiPFZtxciLBUG7
pTMD3YQl39YyDHQJboJh9CHQtXkoTy4BvIq9vEKt3T+EMsieju3dBawi/g7IWCMo
oLP8omM0WS3sh0nYpFgL+Lym9BxoHlANSXfDJ81Wong9EYKVv/CxSH4G+e9uJsnM
qs48uNNP2qYliBpelpVBAA/SfWKb6KHyfamhVKxlkcsIgQHJhJeB9ZTllZ5wB4id
7kR1EMMvhZzGlGkKAdc8u3JjnmQNAfBLiCYcV+8MlaQ3TM/GOcDdZDkNK/7KuBln
UCAg8xUpMVpQJVsP9MNfRBThLWJ2rRBaYOrWNgL9DxkA5YwA0e6RjsMNYl6MGbhD
psqXreno8Hzmsqaah68bHHL4KJd7zy9M0AxPSKaGdhAJ2IuqxGax6TD8Nz05h3P2
iu2iVvnImGSRvK28u+BlWd+fjClMTjF0wrnUP+MaNtuz6OBVewaEslOvZ6kprHRy
e9O8IGK1MR8YS66vAhzIixuNmMxx/IBQqPel3e/Dcx2DzYcv8ZgR6qvLdagBuRFz
JOj77HhhyINlpD2327jI1JWPKyzl3HdeV0qXDdWXgrMreEnoGBf1blwv+MjjTRd+
h34j/xXOVxGVcIeJLNusyN5KZzXdhdd0T4ggLMl7VeRnDwb8n94v6kWhtSJVsxpa
78eGpcWSete9VZn3q1Sjt+Se5hhlG0H/qsLG5YX/GMMAKTkVsoQhJoVCPbem6+JI
Iyt86b58HTpNgzxF1euar9jPZ73EJxFqkJENuqvq9iotVQMGIHikMcL0ggNC33bf
/5Sf/ms1jP1gl16HtUpNYxjL7zFtcYZHl5ymxRli4Y371HBgvVsS+lCnC9v1czWC
yRXJ5RSbrc8/Jlwq9E9sjeML1Yh3Eqn9ay/ZYFKRX/DO89OK90dmcZY7SR6nYXXV
pTHFH93C6E67lEuOZFEABqzTRXDrSLYwO2jraVgyHKC1ewI0ZUUXFc6vBlvX6Plb
gPSwIgUaxCXbsSLQFTpzIxthYslPRRfcQ0g+u9VHZ0eY6BdjYt2U2f2AreryeB7N
bOShufaRCNuVpBOBEjC8eql8iMhGgGIoV2K0bR14l3Onv154IXq5T4tiYGsLsoe8
cHh4yawLXBCaUbsb2RGXoaaLIUXdZGAuioy9TBVK9u85JsbCFrZSoYOqgHi4goMD
1CsyEQUwwQFnahrnBIjVIf8ffZjM21weExtdCP88FQmZfjTvxUjxxofMNvqqH2ei
/FyU9dbUsMJ1VkLeOOr9eDIclVI5GW9KISckC9cDnOX4tYmiCNoTSTINXh38KJxI
Ev4QMwAKQDXAIAadjdD2RVlUlaKBvrttA2DMu0fODSivDJXau1N60LDsXjnCEAW+
zQqbbSGFAb04eiJq3vErvXGR4sq9J8NpsbsbUFtwVWQ0oPp7uyhNm01uFm9wtmW/
Bwq/Y7FvJxOadskjhIBqr4mviCxxItsSC9hcP0hdx1G9/zXirFVdJtNYkYMY5kUq
MHj91IoiWzZTYg5+U22auuZiBuatDY51UjgT3L64hH7IHiRId5dzjQ5AB/mMn0tP
GC7lIVEGscBrLVERwE+NQDITr77c0tzuzAyitXp75cJAHLOhTg9sypEBoLy1Wqx9
u7E4hL/o+y1SnHhQkV8k/bd9XlPYZRwD9/GGY5gdyNDr+0YW/crLfc2JDRGmswJg
Mp1Tiz9sGFhYPSbMFn9WYix+nmfr8lAZjW9V18HL9ztcBOkVHLkJW8/EQTAGxrEU
t2dpYAt3OshBi+jBvlg215vc90CF8sw3Sdvd/X2hGQJeyZAjtNxYFpjvbXGGA380
qbODbYRtNMaN+FwQLvN6ZjKyC+zD7PKOykBWEMhySo0=
`pragma protect end_protected
