// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 13:57:47 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
bSYpNcJg+jPkoG2sxD30n8CEzQvlvxrSEjqX2f/DvyoVznC15GSEqTfF2X2SPzgG
ggC6QljT9LUwl96FM+FfqkmkE2SjAILJT56b4wkIgnruGlYBObA9imWzruAnzX5Z
IOfcdFICKnmccFF5KrnuscGaHvrw9jpnBlq0lvctiJU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 15696)
tpKDSgXAM1NX+21jjEfJsNwANOcBvzIvExYaw6MqysUza51rqmepXil+hoo5EYm/
ainK9cTxPnvccm0Y9IFy4Lm9Lt3gv3Aeo963CaQCN0X1fOeQbJt8CIbEayYWod9h
u5ymFNf2J4qmko7UI8WpCzFZuuSsB83a4Ort7+AdCCWy0w0A+D/4n7CSvvxfp53s
tfZ4depIDk+Gu9IDrhrf04ePntNpUSD56+bKnC9Yu839cob6LinVaUV4A857ReH+
FJYgkpw4ejtymg7dxoOT9W0VEfUWlUMBIm20n5TsBmlhMuepoNc3kxUpO/x4XVuT
N2omVoUODWDZ7VvLgDbWkOznCipQwkeZWR9GOigbrnTBksMiJFUSl9tTGf/e8fjo
4XnvLTSSntINdOfNuyFr8Y3v5JOm7MVPLZMdaplv8TBRXEc0CD9tWZGMms8qDKEY
bKCdbP12b+AcvdeqJ9SJ0Dcphi8KSoXhGKozR7rqvHlElW/xDEedEx1Q6zVcJ6RM
6CBQB7+2esg9njaCMY050elq5xPkOfGCUJEF+qJrefEehEHDycSwLy5NVfR0O7Ej
lPmkSvXngkN6H/5cmeaAikpDceTYoYldF0O0Id2DBjiVLj+KVHauRvJOo1D8AxOC
mXh6ICBfNGZKP01B5aAE9UqjSMRRz3GwO3Wy3L3X5Xy/65kBfQKbKH4jBJYQqJQp
RIRsha2Vs2c12APeg7cXeNx1XVPtRiFPjUlQYLeIIVScikK4sw27uOivZIEzvNId
M14FVEi5FnDZz2888TjfLpvrqmpM2rd/lIGUvY8oJCIhgzVZx8e4gE/O8knqOw8D
HJuKAT6+pElihgy8npjCBK7EYhp770j71dgElMlrjWTo5FlDuqiLo/izNJmuL69C
UHjJscVejyZVDp9z3TOUXVA9JpjDO1nw9KpSDHR3r0HDyxM0OBvIyaEXEbTEW2lu
aWx5qdbHrOFG1cCqMI66WYMSCQKUZR1b4YBURnrVmnYbNGIVXU1WFjitiwbo33Nj
zNXgCj3plwSNW0IdXp3jq9G80c14KsOEWMQAO+4BhkRkR5ilyR+mqLpKkfUPi5Wh
BXrOZbWXq6B7DIeXkVKTnKLgFVuhaEmooPCq1Fis8AqshUh425TUWvGcuujqM4xa
GYkQdbcmB1W9lurn3j4cBcYlRc+q41Nz9za13UywXvGeHRuLh3ShtYre+pAbS0s+
HXBa9ytM1a72X5zvLe7HDGugMm/eeuzHScKq3siDlD4tk9nBpT9EK08bfjsnOFW/
SpJ0a8T1MJz7wJKun/nIUKICcjtoCaZ82imPEe740tBANWt+TET+FmPHyd5/EBl8
JL+cMW1viRNItZPzdKFMrrwAOQV9fJlX7k9jZO9ghwN+en+Ay3zl+MnBBQrpFkq7
GMHqZypqVCCdzIg1saG+YknwHVbED3tiX7ObzDGYPmX1XuYYR9OErQl1hBNqP7LF
8Fuy+3LCbMlsTXiYJfmoszyr3Xm2zf/j3FS/XyfmLr3kdnRWWPeSu5rYmHrcsA8e
7wpO8HAxjxbSo8GErZdGa7cPToP93ZTHtB0fmjl+Gna6+LM/IYFVT+xDtxPm5yEU
EOhtTvsizX/dICgYhcc+04LzlAWtN2Opasr1C+qJjEe8YQMVs20PcGDX7D8IH8Tv
W+mElip6iP/hHyHBXlbZuIL9lsCZSnk47od8ktoa+zpac42f7sraiLE1A+B1lu1k
5MyCDdWxpQnPLL9P/9p3xhz/bTimKBkF4GWSGLfPFkGg01/Hz17cpIq2n1MKw83/
CqRwHHGe8OX+IxTF6crJ6qzn7x1VAKwy1FAqdyRyGd6APpmDSn/BAGNvbAVgrOE4
n63o01NoDvCM9th8WShpyHSwaDjfNapfjRcBkxzsJFIsslCi15hSB+GPPbcXhKyo
NWAE6Oej46OcGunLS6Xxi4Wlg3UvGLPaR0XqqeZndcSitQNvLVXu39Sn1yUtUmoQ
2cxYsjgrIYasR8tgIyySW6DIVkmHzkNwEENx8RuGNRpSHyg4prjuR+rq2GoJIDlW
aZAicUXWybp9BoaYuzSA6ZjXLsg0hpIUERkTnmX5iI4uJBfghDGQJXSpcowEYLmO
u3lGr/Dark/QAs32zyZiTclca7NHr79VmoqTxo2EZrOh6ycJQtLLEb0NOIJavfzO
mYxqMGBQBiy8/QXc893WUsfkCfDamVAZp0Jq41wGhpF4sRYCB5i0ERrhA6bs6QKI
fgZB2oLBva4Bk7+iATErW3UgtaNOFvgVwgPwCF/EsaGpkNVOu3HTsmDGzvi3H2TY
5pSurMIKNEkLJoMihiKWjC/fizetvXfBkoj183o1Mx/HSC5/gjKIGFWVfRCYNa8s
Z8orlm0Lt/otXdxZZhLfLUbkJWhlnRZjS4c6M0cS6pQ9vPFXQebd+bD6dr8UyGtZ
Y/6+DZ7px7+RSIm2KAs5MD/nY/yYuCid6A+aMYRDZkoiCRogMgh+ECPo5O8ikKy+
ZR/sHgx6fL1GSdQY/xqTYtqlJ6m51sE8ShCMqbwXx1vlnIVwdEIJ3WF378KISPsy
Z6mwCq8/LcegW/JO71E75ypSvgo0HUKxlCBL2v6ucw14RaS/Y8p7Nm7qBL5qyJbd
aYJaXSb3Gg6eFZKy5q/36QwPYqSaCCDjKsV3pCT/AmMomW74W87iZfLVh3wh17lK
4hYYhSIkLhC2b1VZo2jvEwUTr8WH3rvqF+3Wwj7a/Y7QItvVL+W8jXzXlliJgmtB
R/VetRT72Lx2UaiB043udo7yAVWQL61GRoLQQdpG4TI9UJ1A+i/5JC9lsWB4IAO1
PHLO9ZAqSHQTBNcVxN/9x1V4hynUuZw/ULiU1ILhuNy5Bu4sVwABK/jgs8+0GmNO
/GBvGQPUTiJ9S8FUyUIiDoASdzt+KaYb3jEN5d2CtiknW6TChEZfCcwIJOhZ9Bv/
Jyp9D1xKWWjSFlbQv99vxPBwjJH5ADPuCVqY7TzxRf03TBDtpW0LZzlTdvIhSdGn
bD9VkrDyVP+nHD9fwjUDakiFttSUhdwjE1mS9z6lJPUfGvQ5NCGorfa0nSlsJdZ/
JMP90GrZHYx/oeOtrg4UPQ/qbteQ1v3lHjv7Gd+Ssv87wuORcLP0+NXgZ22hgWyX
ZZHcjjgCKiYjMU92TcjN9xPa8X398Dqnx34M879p1LmyoVlMJA/jTrqr4UmvOOiC
MJLZv07bPQZCSOtb/bQgDCO7XRZ1255gwlM/2AfnbdN+4GF5PyukfLsYE6XA7Ofc
WpOTtDHUKqaVdMYmegjI5xnDjy5ecITYxpkck3oLgf+Lk/QnNDxi+x4u5mWF+iJw
sqznrZsV+0D2fH657ex3xyBv2puR1vrkL+tysD/4pzdE/TBOgY2e0SlbNNe2RBHK
UqC26V1HEGwSpEBsl17+hhj7rxa1LGu0Z/AoHB0qL6NlzKtOI8Fk0eWZ51kT6NcF
qsKOmu3+3x5ANyk1JPkLtoPBLMyCIPIPCubTOnLkihDKSoRlmLXapsNd4cG8uYo9
IDBiPokTgokaadqmW13eXqHaGhx8uyqraT1wGlwGzJ6KW8ydm9SvkZMhB1/2uz4J
2g79E07GyzqkQyM//P46489CCcgiyWX/4M/5E/4/ggXBstp2ccV0/UavHrNkevvx
Y8tOzT2G88hpzurZFJpDwVaVmyk+4Ii2kjbq7rU+vSBo56f2ILGvEb4qJGqo1j8o
JSa1WUmqNi/U1hN5xPiroA+2B4oPpjzIqvcTnx8kMhLqPm09CZUnPPoyRWPoMwcf
7c+hDkR0nfc8SBGvl7vuh6wUfiiFiQruhwOy0S5MH0j6dZS67aFA4rXvJdhwjivR
eDH106Zlh+r4af5az+wcaIai+4493UrbKtd0QU/AwH5FED1HIVTx2tZDIQFS0mlN
OnIUg1vQKxviiyUJRKnSr59wDx+C23vQ6Ei3UbVjN5CfeS5fi7yR/Sq730MIsJn2
2V5SXhdiPQQYkz+tKa7vHMtgRelrsl4zTV5HPDigUDkjwA87CDCpPIOFrki+xS5V
ZRmkxHld5Q4hdJu4hPYwaf50EMDWRVw0ex5NBiRX+gPr0meV27NVb2B7WltaGtN4
nIfWIOEnY5jNLdBAWbtrvyNx0EddKYrsI/uDqr9jCNSRflFLxXEVsVKkEXAjkHDu
0JS27OK30gBgmczEw+XiCb9OYWzBmSh3Jbx1Wvfa5/Gxg604m82UuNKCBgolLQ+I
Z4BkEE3LXn5ozlLJIbn0QWEwoC/sta6eQd6JiE1rIy6/gAY0ZmAL4fC85k9ZAKHj
wUMDVvgIxiUH+EhU3/4W0tZwMP5pZdW7ei2oW2xVzROH2o88wNC1RU03G7wadkec
te7k9sVTaVNJ7P6ZxP1AcYAbg1xpF5zmuxKAGex77ZeN7y1+Nb/IOl5xaNl88f64
zJByqHMwxxDnGdTqgtYZzKaDwO/XZyb/XOVaoMU6hlxLVjuVxjyVlsqpLi/u+HI2
qveXCBKh6mgGSbSaRLdW2LU2PdfZfdTPrSrsbvI3a/K0d7DXwLQ/oPiICaFQG4Z6
C4RCXoxPAVOJPBs/++DT516/riNF1DRTPMF4ImRn4Q0xqjaoED2t6kYHo6szx7wS
3HrryDYg6FHAS3etDh0mGZR0TzcESDcB7HrzLm0KY0DVR+aOT5D3zLMKU4LrKLw4
r8olvetu8x5PR7X+EJu3T8z88ny8UZaPaNkA1u2doCR9XOlBxUP865VIYbK61TqL
wSSTeBlRCvux5PVEyOXJ7e5zJr8XErc6EHAKe//8V1zRNfxp2+Vnj5OJynUM72az
Lf5KsvjUvUs+iR5t8o5P+5cMCUK+7hgr6ZjeH0H/otmwOZEyiBR8977Q4yuEyBDD
bnbq7rViWawR3k+32DXMTXmmJCD+aNfg+4zucKe5ymWMkGNI5tlpDecofpatiC0D
xKL2cnK5ok5x9YkbiFJJO2mU5hKIvkNSKrYn3CGa9l0Fs+rs5wvpdPv7nzM1WMAL
nrRlX6xOuPpcU6voHyzJwllLfsTdPZuc2+vP/ynU8MTjhLC523y1bOngNxLRCwzZ
9utwe5fya5MAIz5qmmqSK6jjLyD17+RzVKDaLa6tKSP7BWoHqpcdJ+995m6ultsS
mh4nTTxN6C2NQFrjfyNHALpWXaAwIl1joOj42na/Nm3k94gN1cKu3qmvBc1t6KxW
PZ+vD0UaSNflC54idFoaEavnteyLMtHMoXFkYXSDT4HBmZRR1GaEydrLYXf3xFJa
kE6EUC1lnVWCsk7Oag9Rm2Qr8J1GGvUZHrFE0xxZA/PneAP3RD6yg94gSKuP7mtM
XSpiZHW9Mn5CDfyX8AxImkflrmZxM4ACsKXVC/SgJO7PQEd1QWJoVMhxuptRvxrA
drhmMW+pSYMh+iFoJQAEBOD138tgIhTmzjzcmM6w7+wmt+nzBZR45N4ilRuJMuiV
Ou1184vVPMYYUwvN9YpEdce7MdB6qCKoe9qk6Zf4Uw3aKcRWCki+0VVRCsD2+wF1
VXRZEAeJHRYSyiwwiDwEXUqQlEbhvk33bji5Hh6uzZqwVgO/BAKrm+ittHwUUkQX
7NjUi4JuOS0KoZ9LzRoWkcd86YuV5jDGd6ckT1fbanc963lTgWnQx7nPYVFAz+U9
2JQmiFbeOBUT0MxJABMVP6YZ8NCSi/uV82PGbqykVXVeddQuugK6HnMk4Yp7dgzl
pLT9JZL5J6oLJ4Z/lrMzymY05HWEIoA2qphhKuGNyfz36FfeeEoZwfKEaQ8sfEQI
Hss28/vYLRAqHRJxn/WPhKXnJ70r7uKmMi1LI1IkcjRUV6p7G+JgfkdQN7picxoj
/61ud9X80Ghn4mx+0yQ8G1SQ/3DD3UebjjZW9stOQY99swve952aFiFsSrLOhNUL
h2pmTSPlKQCyOvu05F3xABye60cPndwbphMjITMTWiHaL7OTkGjXq1FluCfzH+RZ
tBloPpHnnDxfG1R+h5WVnjSVkK5tjWlu49/36rn8TJT7yQ+Qf5jLnmjHYz0wUZNU
wHYG36flciteW5hPAtkUkY6qAA8FJBOF0Z+3+hBidfEghqXxnMFEle3yyMQ3Qi7r
md9RPdKC0h2HGRo8umzpVBINKc22Zeyozsk2fe3qQlb/JOzojdLNoFmtbjRWXfiq
jmLem65hkqdP33WlDuIxglF7QejJxiDDDwW0nOR74xAYLwC2zlVc32ToefwRVP5G
HSTzqqXkohHjET0dOP7Yvnw6gJTIx5n9lCZMa27TxHrpteXcm1QQk0zJzG+Wr20b
BQiWh1BQHAuDDLY7wqs+v4O5skAgn/iBESvlqbxL7WH2SdW9lwO0yjU3BeQlAsb1
BJGPilX78fwUoSvNo4tFY0Qv94rrJa8kxPy9yzTF+dscN9U3+jTEAJA8Qh4AMSXR
qxuLN+8m495QYZeQLMPNHIUZL5vz9Ka+Vura4wYnhWQZssR9Zkx4KdazEvq5qwte
hj7b9ql3OXERbolD7TQ97KP0V85sbjU37++L2vPSx+ZM42hcOJzTbsIkanzW9Vgc
4H7Ob1MZb2bzstDMtmxCPRmm/bZ322ipm7UZ2WL2dFrG31Q/tw6qBsMg0S/1ao3Z
u7oXOxGDOgTzsG7W/dcnzVoc0O1qMofU1erOjTQ36HkIz0ajFpkxMn1WRSib9etm
BLei35z9fLHbgWO8WXTAv+NVKVtjHPMoV6/nPelUz16GB7hsQ9mmSC8QvX7akrgl
y1zSFzAjKlMcJFCLDqGrQ7zH2zzOnXBNHRdleU7thNSkVuecBmH1NDnZyj83kjbF
KMn6n/LfYG2miq2cCAIQ42lveGsSNgqI6cD9dLgvr061TzrgDR5N9P8562UV2tAU
Bbz9/fU6EnaNv5e/kwDjYm5dX851ECCaBAbUZnXAnqQyJ5ndiXfIFdUbgYddC1au
fH1R/d4VjqRx1Zn+MG1f5PvdvJiMeni+OU00wZSo93jZdp1JLfUmzJY3eG1Z6QMD
F7kR5Ph/pDkmRf4V5zj9/63cVP0aYlNRuSCv6Nmm2mEGDuFbug5GUqRjctk+cYQR
26uAHYya/M5rBBTy9I8DT9U5YjJhVqM8Bi1yww85LsDdFD3awaZXahUE+xFpjvLC
uvLu+xdJu8YkW0IvB5zSz+wZJ5ej8lKzvGPi+YQJ0DDq+qu57Yr1qqxF893mJzFr
Zc7FZogMJYM9Rd3JsRb+v/b/B7MCbU+B72OhnWgbybm6i5S5bk7ttPkPAA6A9PW2
EQMlggfWkmU5+xYgAsfgJdYdy1GkeD9xIRXL92uhLSzAHWdk6MZnag8flRYd+im0
+wM2soeIQcDCVJdQWtslo7uEhiM9ye6W/j1Wqk9NT3JwNmnq4Xgv2kvPtTQA1Nu4
QyU48K+EPuB7yF9mlLEOyK9dyJqERpQlW/HalETXY3wXnP2couxLrGPA0U+NCuhR
Fj9UAnwBuCP0Eb1C0TEdbHqpSQKzpPgvfHM0E6vTZjdDDQsGYx8R2zOa3RD5dneQ
+VshueHgG5za/ALL0uZo84qHAQ3Z05m3Xiv7IZvHPk8cX9e6o8cmeQZDJKshLwbX
P5+GxMoaKfuJWD/gNqJH5owgyrdtrMdRZbCV9ORjkJ5+cBSSZfHCTKQhCXNPMqHF
i/lfX1Qvznuly82jrHHlS3Zg6/rBFDQJfaZysdwH7NlXY+dBzh1eA9jzYCaztCfB
SZG9tU8VV8aKzPFiUSNs5Mz30hjKAfJBXrq+JMh1j/l9ZvP3NdCdmjAGn+zdu4pS
HhrRZ7zel8+ea+s3c4YltXSq9LO55XNkgL8Np02uJypE/wxQR+Ra/Ti+fKzO/Qn4
YwLZqJiw6BOOKReOrhxBYxFk5qu0SoQdU71yXz8hDMWi0sIw1Ut1NClt19hLbilg
PiB/UnQtV/d/cbALeSmRhub83by4L+nTGVgYPFLeKvPC0Vgp4mKTK1UFZnsDvXnw
9KHr3TzZlFiWGovbpd3Qwk2JwE6dDH1uRI0s/zSzdI1HgUbTWV5jT94SfOqEk16n
8YxUKqpPfrwiLXVryhJ0R5zqPjL9IPFhBXdeuFfgsPYDczSojSP7rIrSfHVsBCI/
EJ4HBd+bMtl7hEimI3Vhl6c6Px7+seISB7aTudI2si0HO0Lrg2sz2H5/ySsj1A2B
d87knHQpFInlAyMbigARJfGbf5C3iPIE7UIOuZmfqvL6rofhIkv8UbBJdJp2Y3S+
bw2i78z8r0+Cubi50038RT6svNCgNHBSJouDcKY3Zrovzsh0MpTzdGNRPJeIcWCs
z7Igd+UjK/+0TL30y4umcVCNpZ/to6nR70Z5H9FUJAo4SDtFH22t05WTgeESdESe
rOEGQmFydm6Ei3kvz7h+dV0n24AA6qTusI423zh/TuH/roAvhJosFVJIaxggCRSZ
pvM9jmXHR5DH8AMnBKkwGMWOXtxODx2hPzwqHzZ6m+b9LIrjJoGygKHSwCsS1FX6
q1pU+QIAZ8eOQslxkdNBarnsPKTXES6jLFXbLnJeQnsEHmCipNgYQvX6X4C4Ydl4
7scuhjh5tBqxSy8fY+roB2Hdl2fghOL02cESwXDk1QSc2M9xs79wc+NuHe+d82nm
nfz2gu5DZzjuj/M21UBHLvJxhAu5nDk/CHbqhxLGNn+lcNayettE/1DFaP5BRVzD
6m0kroIbqVeT4+N3GNVXfk0ekQrKTMTOMFiSptKwr4ArMPsCR8WpVezFtYTaBAlr
wNq7ApkxVakhxmf+ahHt5A/iReKpnIx13SbG02lk+e3PJJfe53zoVoTbmNuH6Gju
MHVzZNJjnefZqWezMIm92k4vxJveKoB3l+U01ZykNiFwl3ye3A1bEbr4bhu/VA25
Gdmv19za3ZqDdeSrTebxJLd7Hcb22j5NT3XZr61BEhj3JuHbmhSo/DJ6O448s8cX
fBlXYKCVe2Dh8Qqk6XPTsC3xvsomqtqw+Izoi9VCKidIGM+WUeSE1td7ZSBa7jKi
RZsP1Qpssb9vZBlYlGwiXHCBSp0ZDdourAm4bnXRCpMmum2R9yGXW7cPlzWyMMjG
+jlsGiB/ZyCcCKW0+cieiC5uYDYgFohYwoq0QryyXqRIZ9WBwmONZdligtQ0AzTh
SoOK+/PegMzEJovBxDtiE+89kHovkrixumHrRX9xnH9kUPROOpEcxnZaGvhS7fuI
ZPpaz6BtoM8UrXWf0RkXg6Fv1gKvVyXit3iLxIwZxUXDvdvZiGbC/w2rSwNAdXe2
lSTr/NxE/jRkZ62uvNWIpKlY4me/om6HOvV11jzB1NmxzpFjmKRZsECAsgX1tX7U
/YSj4Y0GCGABIH+qdc9e6lKGUg7PyI9afczxKSy/RD+modDigtyKtxmRx3B0kfSb
/gvpyp8ybyIbe2F8Jog7+fM4IeAkeJ32XengGzAtPVsNNdjym+8oGghQ4J2Dsbqp
LI+SQ+YfvJi/gbybQSyqt8De7C6EEC3IDxGgMnWYtRZyd+CaP7qzztq6UTvxiFDE
vgfNW69zN3vGOUzo0oydrQLSpAyhrOvpnLtneRwjOgyLOzxW9yf2SzurOCtgtw2w
Y+u+cobvpQYWsaNq23Y1LaaFB5ILgo8snAhfrbjvV29ameEthdgh+/vWkNYh8VxG
ORr1oCjcwYK3VzgPdzsk8yl4/lNDGjNhx0Tiy4CJtZEnMSADDlD2+bp0q1r7HWKq
qnXzAr9FrQDbDtqSgrVtyvfxr0eb0b2O1q8JxhDXOiOq5B9H66aUK30wnARrwhZZ
1J2+nWWHrslzoo80uesqhm8wg5imRCg9+ZO22ImRAOFZvWGEn91Hc8pZ+65tWhrq
21+qNmiVF+i7eIBim7pSl9dKincy7oaVhV9evraTdZGSRuf2N/ngG7kDWTKb3Hr7
CeDyF8uG+vmtGyvFY8qZYcZ5JK2XQLk8GbbZq6uKkFyi4dYrDpkXM0C+gTmwyR+o
okoSDSzkeZ6CtvcudRLBnkGbCRrk4ZKHC7hu+75ZWi8WyzHSVmBk97xiJrvoKbH2
U5hPgl6S9SV3LoTQ3eseofJDneXDBG7ieDkYcP5AJ2tz8rbYKDtXQd0QffMFi94T
bpgJLtNJhupTbuou4afmFvhU3g+h+f046OasIOeK5oA9qY+vBivmS/1fV/XkCxS3
zMzquT7BPWHqIQsNrRkX/8EJ/i9jVkycGCkIbr3VXWIFH7GxYF31dsJv5f0xfCDK
UPUZzwF8NESfL4IOAO2fBJIF9RTT6VYTGwTCErER+g8xo6b8LzwfS5Bz5AuPoDCa
PuW+TO7mva4zbpUQ1Hh6cJbsxM/7lkl07Ha89qpVXJiK1aZY9DmmPjw0ERH0eXxX
y/5P3zP7WknLc5DPot9PFxK4xWCnj/+zZCJvSH35LQZZZma6GeHLADpgR9r6+zcz
DEl1PLVUwKnYvzjN3gJk9gkVwEOvQttwFuVTNcaRMKc3UoCdBHLxpyzsKpCJxI1n
/1QaJ2OOqK4dn0eStrGZ92alI+IKSTYUfBiGfHT10UnqYm6T6WpKbhr6DMJHi6Zc
QHlkzIpKcvTU4+ybbwJYR1wnRxXkhjO/vxJwXVeHafHHt82xQjbke3i2AfcsUC37
XP1+B30Y9UX1EsQZgyXhTEHIWJUGVbMvxhgN26SDm8WY2IYUJh1mUW2NTL5y4KDM
xKXqVPXouJ1+4t6ga1sphTE2Urr9xHvbDsuLawVrxq3WLikH52k+UvMt4pBvppS5
xxwDuOlnLcxSTwK93RUfP+meHKOqLcL1ZpL5lEY8WMn4fq1xciNtflsZDud084Xd
xnkibYdF1mJxQpp9/XGI8KQ19rxdWqjvtlXHKC7D2nTunwQ8/36vvYRBF3ypQLvp
V2gGfxtkYcEuEbGNyTemRgSR1GrU1hqlE0OMCmVBRVeIPdgUyb0LOu2bZIzzvw2T
NOiS4c24SUT4ciP1x7FgURfG1qqdIQfNBC66wNo8UDFAD+Tn0Jg7TRsao5GeIXzO
3QLhyYfDiuojrCS0P0KhYe3HyRetWiYB4jfyezJNr7RC1j1jnQiNByV42FPdzJ3m
wfe6vsrBRAuPyj3nv4IzIRA+8A1w1+se/4iie77TLa+dZ3h1QzbSjQU2c2ZcvRiB
g9Yw556iyoVhnQrUWyXXzUeMkqlLbKH+rrQBy79Fi6ptiG1apMCFOR12bdMQiZIL
lRVWI1n6PT0jRVZycgLrXDSr/0rdhdpFN4ThFoPlv51az4joqEF8idLGnfAHJKfc
HnVoLUSe6IwPcafmXSOZ4WHZnVqxWIejgSn9i8cs5BhRfQ9G9OBnxIgxpPJuoX7M
Zti/ca4AH4yVKUhqN24d1Pn36zNYN2R3dDQmFvms12NyQSOdRXVbTvIPwlxVjZta
5peBaxBCNVC2KJDzgzroqrFDJ2KtJ9/nfhPSAvptufN+wl+xD05q6jwxj5+ew4BX
XFMuULqAtwZJC7tR9PkAQ76NsGNqk+czwM3zEriR/kWudEthszfGO+WZ0jquQ8vZ
BV6O8nPulc18U3e4eTmxFEvAPayXoIn+VygriDehvk/sb1RQG65gEOTNAutZPKNa
fvYm5CFx4SzvHQiJ4760qAdS6oPmt0ZWSBtJrkB8WfcBaKaCBkei0FmG2qv7BVS5
bCkQ4ojbfe3dQrLsFKcE21obuN2isjYsNa6UE+C0mV7kDF354SZejOS3e97vcgl3
ZAsPYPvEgcH+W7RHlddsJKoByCvj68kRo0WYYR19kSqPOK6euKBjaRZLgdrDamRp
aajtP1fPhtgIjyeYj3yyLYc+2LROZqxlufWfol/zn9acFQxnQpiyVjccUeOLJYOJ
366gLisn1Vzy5OlmpMHI2Fe4/n2+ZUuJ8XyWHa3JRKJyUtYY4/v6LV7NjYIaASBu
LF+8mf6aUkw0fzLWBPJHis9diAltDHixVU1C+twIoK7UIpCbrfee+jLB37zY8jNT
ft3MI/5/ov18vcZQnO0L0XRWDYEBZDJta4GwXry58UBuj3uu/jKR0hyI9I/5uwYT
2JMb0scbAtdkzILnihR3DCOIMUBJzf1y4/XVjTcN7Ba52QUYd74uhLDQlsntrkB8
KR5ZyexSn1RUmJBjkGB8Vp2KNm9Q4uNsABHfEZWFSDDTDiOncqaREpBFJzeQk/9k
9zqliQuZ20ZGiKs6Eig4dZ1VLK/sP4v5oOmOzjcomjjasbV0rXa4ssrCO8D8sO8/
geDXnox8oYRolipQgs1L1tbvUbiEQ2Qi+WBb/wvD+95ur7GJoKFyJUXG33rYEU0v
rmJ2pURJssbL8kaDk6/b7BCol4mpBW929JyB2+sdwU59wygVz+Q+nYH/9LzD0WiH
nktOA2NNf3IPy4bzvRPBGqhet6508oIMX2/RngEZwUFUbcY4PNsog5r5md09rjQN
i3eyUtvai4oMjtnFcTPyM1z3xONJQqCTX/FSWJAWHrPnSOTQXMgsx/Omtzd/n7aA
andGlewGE1lIOgnk9X+wHPCc3983CVCCvLHSAbRO3NJGfqQBVxklcpqVxo8RarPf
HkNBsFT/TwZe2RG3YiPRlTj57HWmqKSoT9jEnvePvMhGRoMoIzkQ01eeZWaS6n8D
tUc2cTA1ma26IXWS9rTdrrc7nYaaanGg099aMQg34dTEtn1vDM69t/QSWBimkZ8g
/8MWoX/gTF8o2CZ4ySXhymqd/LH8qgihW+JtbslPgb4jzz+SY4tnuFmhjRYJTaY/
coWC5rG7hfywbMk+mfEdpxuu2nLARIdgJrGakDgdRJUMdIzFUoTalcUQlW3h5Cz+
xUx801fbi+J+e+/GjLu6tgjj+jer+KIGGc62fIILZmOAkMCJN204uwWilqFZSfnY
dAc3tic3u4A9qkBvwxCOmOjdYHOBev5kiXd6mzI/95aTWlaBgb2Wfy3z7BZv+yo/
i68cVz0yUtoh4WBhymlDNIpjzdP1IJJt0zxAmV/4e+bGn0c99fLRNvGAaLkFh5A1
/LTum6ujCKWkqUcSiMuxmV91/OhRJM0VpnwtxqvX54uICw4Nn3TNOFv2YxE2sNw+
VaW1Xt1kfdvSySGmrBAg2NUHQzHgDxf9rODq7RDW6JHz2ZMacTegxhW86oxWevgn
ZWQlwVQq54eXavf9RcJz0CS1sXW5cf636+/HxAr8d3d3LgxR/XbrrtsTLKRlzzX+
WWRJqjMmOLPZhyCJqHaQhs8cPYcCCydaqJf0Wa+PF0q3Bum12Bl6o2wDeiLKZNHb
Hl126HMhPMFhzl6OV36+cOi9RHJg9VbzY3rcHYiouFjngxQHWiv5MI4aLl/necQR
gfGjEBKccgMl7zh2WMSqY4rPgZIjbyvlpFO7sMTpFoFYtsnUZ7hyjMOj6C8T8/V4
RzTqUwHfGNL1/ZDBQGjngm1oK2OEQdP+MgnCHxOfR27U03DXe1hWARuXd9ssv+FB
XvveedmB5qzbrbxQq34eznDKScaUXOG3PmgpeAgE8KXvuVyd71KuP7sqo+Yt2y62
fgpqbtElSimDj7/26KJLXZSX620o4Mo5ffO1M8zbfICdOJsPOFn2T95SWUsA3b7S
vRId5IPYpSp3kabSbt9rjpWTyLKR96Agsr4fiEhx/8AU5i/tVW8a5U8REYFvCtoo
fQAcBGJ+lCHrplCqfxm0cnErRePF+K/rhCZknNFSiUUcg75mNt074pNE0d6LLBix
DXeuqKF5TMIsbxyBoNYtlLPbI+ukcrGnBmzukBWvsIoJsOAeeWAKBacSSzV2nh+H
1zLITowQVSybdS/J9+Ud0hG/EOO6i9NtkDX4YFaFrRCAWBi1Ohl6Unv0te8FUBur
Aajf4wcutl5ZSBHAOvTnivp0uXWYMTJH+yycmtFa43NnA2OcfUzwAsKVDz6epY0r
6ywiSKgD9umYoox6woLPrJbPqjdZ0IMGWbx3v7/7l2nmwXE2myFR5GSbq7TzEQKi
j2utUo47xyv8hlfp0uivHDcw4L6rGyEGPdiTzwTgeELjNBH5RNnHjdcyzuItMLq1
ijOxNF+LJcX8cetX3H5nKh6+4ayrTUXByaAcWbjWk3DmBJ6jNqdhWwohpw4h7gwj
JsJWEk5diu/5VWNdo/PoFlqPlqqgLLYlFe9delyR4HHJ2MSItVw3D6s/w+3LVLpj
g2t93mhPE6y4+rah7mEb/cmUeaLL0+8M1Bgw2LlYBC71Wog0KtEaRDfgNL2PKl1L
Z7syJ5KG0q1RGffYhz6wbsFizBC0aWBYUQYHevTE/tCN3iEcSJGMNuPiCdEJWw0k
jWkaVcLNd7sZUyIncR3u8H88N6nY4DjiMYgOXWcm75LdOAlHMZmlrc1V/3KJeHRJ
k8ghs9u2X8bTw2lKo+1aT1+fYy7V6KgPlkMjEzCndwafdMzxpWCZOkDLDMAbSoub
MhEchbSc6v0QmwxB7UdWG8Tcb0phcbHrSAjouwDhFJFEARFPCp3/6kJ9EOmBMnQi
neNgd9iu6bYWtPGJ7DQS89rVpX7zckYKzTnB/blCIa2tEf1nWXR6Ze8x5mbAI8rU
9vcAowoCmEIy5rs3xv/PDRCj47s+hElDiDeU1T39UBfCny0oNr6r2CcSGeKr/7q8
GBkogc6jCrBYAAOXFhqWsOMDGbGIHegXmiIjwU8MDY5B2AnY/JgAEEjQflE4COeD
7ETzcQowxQjOhKEomoTDq+53fS3xR43r1y1ePYNZpcfE9omZzT4xdTqke2aBs0g+
OhpVgfnpLLmP842ZsPuRTZFB8w8C7DimGNKKlocN32CjxAX5sejqHVcxQw6SK9Iu
GuPso25IVSyYphxOGBc/JaSngBXQG7bWy+ITLu1dvShDsgKpsDPSnH4oCoyL/MLm
SJxFGMCXBFXjeSqtxN9pLASZpaWMBsz1ZVzmY5V61u1sWKu4DfdF1z8nnPlNLeTe
7mErrl/wkOZq1FEBEwdO5w1KUHvPkywKr5h5z4YNqUp8zhjsEKnDW+cMYR+NPvxp
7Z2XgVY+OCPm9UUXxUJq42N6CUGJOgVrk90uzy4r8nJ7fY6fzP732eOQ+hKqqtEa
UzgyVAwClMbNFMijptcwe0R/2sqbpkB6n3f2tqGdDGD4w3ZS0hpw/WBRpmQjd/ls
mwgFvgQAaWBjzrw+6Bj9g+zUXk9YQrOcL8gzRxRvVoHfO0R5t9mYmyLNZ4pubyDi
SSimMwvsNWDG8XhfsT4+xX1/+n6M3IsjR6HEjyp2em/A8pnKKI53VX7FKPv4pAGP
apqd03kuIex7I44O4DgxCcNMSpi8RyUXfHu/xM7SxLTKPciM7Bsb3T6glhNkVD5G
srIPIGzu3bN6+nzbiAj/UfR/57VD9pzeOtLkhQvEhU0L4JqPoYs34HhojaMef8wt
RCfy8TcJZEK4M9+l8bnzWGooYgv8jwJ/eYXh1doCtkqmQiCcYm6eHHbVIPdt4Mlb
mAjTwu57U+ql+dwqEJuMzuV1iLC0j8prBFw+z+He3k6I+wYWbKEQ46rx5HKutXTO
DnllkjwHfHOUMluDhcWh50bt+TIxaeke5ropLBlPmj5AEedh5an0JDxmWCgLT/se
r8tHCNy40DnUR4AgxRPN6MWLk0//VWAraQpDO+4pztAz1m+z4rQuReBfr5VOnIgO
uCSwJA9py3bB3OPYNpHn1geqfrXUcf9Lhp8LH0MBZvceW2rQqXPcQ38Em6QdNQlb
UHCbe7AsOwkfnY49OF1PmtqjNKmEQtA3vnRkQUOSQisI4ZR6bm2PggQ+8QVO5q38
xcMuNM7qUnJf82vhxN7l2diD2RmjNovCqEYia4MhKsckQ4ViwCJ39qQm9Aszutcf
HY2pIJDjlaRqLJ59I2eNSpyZTIx0h42O6ip2//4TRiYjVSuRsu9k1KuA0HX5Bz3+
eU4xt+trEtPftbiR8n5RhVBkPNSECh9DdtH5g2w+ScSTFf3+gw1P9Sbu1i9nfUf1
3CMAFc27OTC2B3Tbqhf3TCl5Z6WZZ9VBs3zZjUGDhJB1j4dIemmEGAhpk5LbXjLq
q//xy0qZEmEdkntX+rz17w4jEuxh5KQroZGDj4kAXqTeuG5foMGPD7IjZeVeeDpi
xuo/h05IwUtHHWwQrwYz55Mj31FGQn/E0+qYpLcZGTSwtujvSHUCz0ZfX+BKl3ec
XjVAhSPR3g0jSZkQLnu7XVkOLnfAGBIqN+TtpogSmkZVCFa/aAT37yDMjJZy08G0
yMzm5DH4LC+sOkGa5oWkXxESuNLn5JLfXkUrBuqt6+ZZwPfWfitPKLajtEt4abqx
TFQd8k3LF4viUw52YIr1nJs2JKRWCP9MZSO90oVM+H5iaOVx97XkvfdsDVUKdxJi
ED/e5jaX4w9fGieEsQqUiw1QRWfzNy5ceOkuXcZDuxJ9r5uJxYnZ+jQy6IjijK0Z
YVZePnMkIH5s30vAYzERMVGf42qMY7fcDzqJQQ4EP0iSXmSj9R9mMvvDj+wImIHU
u2J06EzXPdCVTGu2tz++AzW5hrt2HjYi/YscRrssddscEdHco/olheXN6xMwtq1d
H1yGbbCZa+7nS9+k/pHQweteEF8gsABvaNQcUD5yQwlMIb++rI8RNJl0zLmoK9x9
T+3hy672K6GKHGNBkZrsL0MW69f6ft0ZUjrH5uK2V9xTiIAyEKr6sA1iPJfLQO+N
659m5BrSQRYPwTo7ZsDqo8bMrMoqtRPYsWqkvo9dVNTQptONhle6YZfUiyDxpNLQ
fbSN/8PHZKqseNFyIXFc/Le6GEyXTY139CMrDfcVrRnxl65qCRuAOdJXGNuu9rv8
K6M2ZRfZiuJk5Y442HsaxDhQwsQhbaUEykHsFpziBBYufx8qoIXiFXDsN31eNXGx
I+se/hGd+yysMudv8eJRnikG1JUyg+uDtfKF7abz8jJbWwOXg/ux/Ki8h2qwaD30
yXPt+I4A5Yv0arLxm7MPC1wTJKiWB6dzJXfwujqFcYv+i+BafILaW73d1OD6JZko
FAH8iqGifmkFiOWFtAf1etV6wLIu/iVP2yXKzPPC8UG9oqT2YwYSN0cli6lo5xrA
WPf2Pp+ngHSoww1FyZ6DZMXl1p5rrMZzxajDOmHKWvk6DISKJ2bFApDeSN3408M4
+VUtR65v+O7yUrILQOdLCsCMYZSEsvFxFD4G3QtviwYm+xgvjh5Wty0A2HQKzzff
RhA/ASPrBKQFODj+2Ov4z0L7MZKpbKS9PrzVxIfQwxgxYQQTV7HE5auG8/vfTnWW
7U3nCrLrzNkAuyCfCZtGTt5pYsUwnY1RSwGB+gQW7Ift99RdWKhupXdV4hdm13XS
Eu4rQCVJI4zFbb5m0pbvs8JE9dTEISZJvQxzjiLBkaTzeW5qVmFj+7dE9EF3qNXX
gX5iVQ3SLpIdeL/uSmUVNudOaaT2Se2Bf7HBZ+XE1nBVoIKt6R/lvsymfNckpVK+
WRHFNN5YLqzZNHkjfgNJ4Nu+UqX2+M/9yWLZBwnQDgvbW9iUJSMZFm+hBIEddtVL
ewXi1icb9D1QrnogWmwWPjBEzPTzWNPtx8kQkGVzWjMMEvs36x+L/KZ+xHpEkMWU
As66Nzmi69+RxhL0o2Olit0pgKESi2C+rapnQeeFLMLXucGjYH/VlAXhizv0nkb6
zVVx+E4lCPECbb0nV752K53Eh9ndE2fQK5/YFujEvQI7Y4XpNIYhpqGgMtks5k2m
vUttiGAwS1L78Pxno30moYW7xaifly7+KjzCvlzdtyBsHS8pzYQ5iNk91Vd50/Bn
3Ur23NqBjuwBYe+BRlIO0QOQiQRUPpY/2QbsJN/zmU5M3VxTekro88cj1RsMTahY
rJVvV1pUc05Lxsc0RJ5TZmdqrqjqGj3l2aRn1JPD6Z8fuPTaOGxcB9QkL3bcKDw8
X4t0zcow03eav5bQVl6Ns3ohRiiO3Up0U0R/g59eCXi2JRKnNo20G+I6Lt6mb8DE
nFDLz8zoD94dMR9ENmDnxZnIDzWsql1HAkiy0x2ScM4Ej9eaLyxpP8W+7KtiW/V7
Qdupm3QYcZfehbilvcX3D3YZ34thHMHRGeNAIy11h24W2uzcr/JV+X+W0CybzHuM
ibBBFHLpfyE/QM5/p3OUJw4pdcfCsOsc7ZR4qj9AnWiyMPQ8j0azZZJSMc4QqZ+7
Gkj5s3QBxLQSCYC6xBqqkZa4ZAlBq8gmflaMJoSK6I+lCTWcKlJdu++eDoZFFnbT
KjkmCAjLzCtCcO68YOs4HxlWVMZ4XEr6CDXdNg2vqnPuMQijU10+fQhKw6L+Ikfk
LtqEPz480L/Pq/AptLntltpoSsJbL4vMoKKvIibInqNfFhnFu0pRR1OA0eq5qsDG
uJYKScxHbPqtJACt3KHJAJ6uhbqq8wrNoxoTxux+mvmL4zTCEv0MjE3fstlybEQ2
oArEc6KJB/00Fy18CnbIn2/2ML27ZUL6eCJclIyej9577GTZbi/5P4XRdHjeVopG
Lhk1C5mMJDViTR1TcQJi9ALiXfi8v6EVh6w+Hsq2Nm85p7u7gxhjmpy8qVxY5a/E
uv2fQT/Tsibcbnhl0CZ2Tvz18G/eRd2Zu3fhp3nKM0XMrButNrNn9szjZLFBxe+M
8eyjsfOCCpU9wRGlLaVmQ+UXi4TYyJVxI28/iiKKOMrhBZ3rleD4/vXrGMHu9zA2
MKZB+NG2GAPogIAw6hCpunkDca9iCfYyq/P5y1z1Jza/oL4vfbDzhdGBps4ttuKC
4ixlxncLHKYKC7q5y8XADEBqImeBIYBeKI6i0LdEOzu2zjmZ0ldczR5nwSVluKWB
hAl4P+grcPhj6ix8GgZJj3FjyIqEX0ymlRWE17arhsuELy5HN1RtRJokeQwC5e2R
LyD7bp5HTqSB27yvfgezkeGCJw4wj6UlRpsMQIwuWYJu9EqJA0MdUHycT+tPCCva
wZhfrekuKJMG7rOSL8TNvPlPZrfAlIJjIVSulsLPMpaTwwD/ERkvYK1mf8vwXEP/
7G8K+GK0cdKI994bt1pgm+nPPJVlJJ1gvtZTCBKmDwnJzSprR6suXFrYk4A8/wfd
sC8UrTxCefl8H/n8TV+PlFIvJwZuR5AtvZG+1FLIz7Mqwo2j4P8iG/a7QN3whyTp
t34ZEgXi6OdQf42owPTiJoWQ+2/tq51zYsmm9Bi4bNudfrzhQleVc4zHEWS3Bfvf
UztI5mJJuJcJKUJzLh1novzzo2W+3Mk1S+RbD7/lpGb3LXLPaKmsL60R181gTYOn
275i2ta/gHl0J3c3wxxe3TaQkHsn3SvQOyFIaB2aOSR+kE8evSNjLptEBBm83nZK
+2gyeP0VgEBOvPSPEvDNpAxL50EnkeVDVGOwmKoRjOyuxXJYx5ofiyI/lq0GIvHJ
RjLFS37wqENXAsb/jMUiEeZJPJzxmXifvloi3atPZpnHDFUFhcGP6/qpZq1d32XT
Uez7AiFmDjzRCVWG95P7cP/CZ5+O280B1pcT5LkjAtyWx2781GiGqZ68Y+yHkU4y
JZTpBDKkpJ3X9YNxdfwn5Y7473Pw6/ozFd+E6lyIkWdWtx41oD+muPkizexylNms
N0RRQN+/yCHKt6/ZzuGuVz0LTKN6lCb3CTZHGDcp1pt65yDVHpGqMYMuUkhM96gN
zSRSGV6dK+IIQh66Q0AqEoImH0P7uPe22XDV8oLCdf07cmbrYuJBuBnEyY+4Mt/h
YWdZ5zUTQfx38K2v3RvT3OTAXjkbmTPUJRU8qp3tyCzyvu8FtBzx30l89l77AdBA
bWWABMGIh6rWr7OqbDBak1CajwCgwRWUIVqWvpyGCahzzYyXM5EbPOXHBh6wCC2P
Hh6Jh7G1XdFKq28K/Xv3tUqPZacUlfSqazie5LMaKrVtyQg3l2/hQTYzopiUTG4Q
Mr+tCYreaNGO7YlUA2NXT81dsHqKP0BfpUgEWAdHeuhU23iSEefo3Zi9fdC2gENf
6cHAGqhAaJ3XpYDgUt7VxzvepqW+gf11RrOKfz00p4BookrIrakJGISSXlhnAi7f
F49qEepz8U8t5OiFP/h9lIMR7XODI+466qWreqgNXzKuHxG7W8+/rKBd33rETwWF
l8i7l5ObPfGdQTRsu0Ebq9RV75fNREjoCGkQoLE6EMRRf7ROpZ5EaRkVTJckmwB6
qc1N8LLS69GPrzvfja+BCB0fK6u94qj1HItEg2/7kj8wYTIwgdiMYfhtu4gOeQH5
lDH1BggcVF2Q8qPhIaDGN4eACgkcbvSBgyvTlSxw1+/VXkavSCPyao0drTmTE0rE
O67qZPnk4cY/wbWHTeZdB+mW5ehXaSvjOjrc+skZrIgWVfM1iLw+3NRH3duP97QP
PxwNYIVl5CAAkxsLfwKSLj5s2opkmCzq2pKLXXWFFY3zX/+x24s2BVxwRgCbIS1V
O7g6nKOqY43h1AkNARlRzuI7MKoyVxh+Yxd/U3snIqEuzs94t32kDKyVo7glgx2+
R4IfHbGNgOXZboHyqGUh00Vr6UurGntQ3yHlQumt9hUB1vWYidZjo/hY9zLpzf32
ryEP+v7Q3KKs2w3vJuNgO1z/7vCK9/1rXWUmwhBVtxNMYLrx27vYm/Fj9MbhyXzl
Ex0Qj6DYF0k5w4EKxvu5ku9e0vL3HaKZQSLaF0usFkV1TTfDCXCCCPt2K+VpABJ5
uuO9tXGkVCfBgJqb/8DAZu08j+C10SrkbikG6qVanjZ8RR3NtWzjpCtMyTD1rRK0
4m+HzBEvSfAkKIcyGeFsNVDUQO+AQkaF/qQ52e63L0GYvD0xryNVPLCken+/1fBy
RMdqistuGboIsFu8uFAE3Fz73Vs5TS36OTwxm1SS3B4oYmfU+jGK7YfLTaOb/PSh
IRzivvAtamwYaWyqutaAhbWjSfXfc24PilYWcCMdQHZ3ofXbXwoKalCzFpW3gW6S
gngkduVVsQ83nl4ucpKM0yp5PHozos6KsXbK4v2JHUjDeW/Q85NqcqIEwTOC86I1
R1pczHmyKLhpumThk+rk+kl7zOcMse2kz1XRhJNc1BHV+aN+hUVEMeUA3/OVZZax
`pragma protect end_protected
