// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 13:57:49 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
TRfd33uYWiNcexfOzplxwKyhXXn/7Vz7jmpPXudDNuXmJh3PiRIaI5g26JvGkO9B
3REZd/ywODfIqw1Bj33sbH2JrgrRayZGTWRecfaEHuyvDnABHGMTlIEd8l63ZCzc
a3UZ7seHen5d7RtkHWCTmS4W/u4rL/20wcP1K40BY+I=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 18368)
rYjw2+znnpe22vYi8pxYlQHVrgmZgQZ5cbFUInFxFLul2t8s0yXB/6HsHtEixqH/
OIF02g6KDWFgaIKb/k6Kl99OG5XQjxhhZd+bru2Ty8sO128RGChn8GRdGmsA/m/Z
JFIh+EfL11DYlx3M7VagG1xs38OmwtcWnY5bCLjlKlBVMjH+5SVnOpfRLFZehcHO
8uHVf/NcuPghnqXZi6NsYviENb3XAP/OHF8kcysRNKn3J3DnIT5qyi3wjaxs/9MH
aFu1moqV63RiCmBIkSr5XlCS9rcxBggxrV2d74Vx5TTwFtp8KvMVG8ycijOrvQks
PTblrpji2WLuSq+QHqNf0HHmztD2t50rZx50xAiWkgLlsf805+6IMZqMi80lwJvE
nnabQ8Oi/sFlU9Y4HYjzAYwkpTPffCJp06FoSFq7d5AqltXXhGib2jKdBfySqUkG
46JoiNMhS7kRCs8j6EXirMDQWZm7nV4pCigcKrdNCTTLCGA91YGbPPd8EZp7wgLK
gdjmdTh/uPoC2+THmPx6+7FUnNs5cp44MEW01WDocILN3qgmYUHjNFayJbCzVZr3
iXCuFIPg8YD9Hx0wK4K7tHkWqLBdL5/G1EaqYobURjxsMAnC1ftcHJ303KdZd8yd
7jtyTLsW3dBydEAL8mL98ncHqi0ffOq99SWovPuetr7bTrnYRR6iXFUmAw21CgMF
fpGOf/V7wncf6MZbDRZwP45CCy3BbGwx/pMmsoHsXi8F60cr++a7CsfMIJSG8rTe
4pn5XZnuFCxLWuJAlZhhGOLFljxYWDFQ/sjsrPeHrCWPHDxettwZ2wy1Xv3lLdGf
Od76hAfbHbNMwcniDJHLlNd7jDvpwYgWLRX/G7570zYUoQ9Ad/rA1sMKguBRVmE4
P+aUivH6YYRl+fbaOJxYvWFy6YENMksmpfJKv3Wsf5ZCmr0b9iXKAUj8/P4nlrRw
DoycNzD7qC2frIZjUUdTYNQYo1jDE902K8HbyXrBOY6TJnIra+vxuVahHplLHA8Y
cX21iuRVuZK0slnEu2zXncKofHXT5c8F0sVWQ0roprkDKwIjjcX0C/nm+deoXKTL
ob+HWTiBiUYE+hf6L8hiTPiq4plgAcTCVfufchnfYJQoo439jc5iSeZm7PSuDOtc
MtkC2Jy0Xo5ZSn2bk2ZCj3onAPL15D/RjSu4NTp/7G1f5RDarJfk5QNK4TtvC+r2
vhxAYS3NAncW4ARwd5w+RkEWvQN7LUfjaKAvliafcRcz/BQKo6Zc9wJd6qvt5f9G
ykCmXiQENCcribbNj1wDrIAR5XrTLthv8GH9CahPtht9AUlcx/fR6J+t5dWk4e/e
4mteDpfWwcIQOn6cHglkQjJRnCOkI15mRiWqRTgY4MeUCQrSxg/aLc0bUbi9WmE2
qAjw1usKqi9Abxn6XfzZS+87FaMWlp7BNRU4azGZtz20Hcdt+cBuzEZgSUwqC4pW
I4Be+la22N0xJ33L/2sT6ARMui79S837BTbQ28PVhEr28vkuP3PlEoAZ9B+FGiyp
9EPUEyViPM8m2LPDcfzYgsDIVJLF+lgj49FCRfgNLrtD9ZQCSCPzTAi5d99HQKWc
5TZNFoCQJdy8I1xQLQQVFbSOo8n4QeFh/tCPXpO6nEBwxH8SxD+/vc7EAcguWNgT
WXPw2rvjmIS6BGvGgpano8gEHk/9xEhwDRXNdJLfyub+vac/xp5rKTToSpubiw5P
/F6L01lPHoyZ2VYActR8xab4GHLjKS5mldjZlh/l5pRrV7Xl/H7p+2j5TCsEVAK4
77fjm9pLwrgfIp5lA+Ssjp52ffcd5b0BK0tmGB7NpblgnK59/drpZqroRTuObQ62
HgLLp7HYO0Jj6TILM2XSI/tDeE2DlgzmVI/MLgf/xGK7V27smom5pQQO1R1bS+0r
85yOqk6oeF/2nnYmaj6OHOO9c4Hgk2JYWvB8nOmdUkFr1teTU2DJo73Wp5ySHnbu
dtA9JhpP2iKvgrllbRZ2yhOkfHLyb8FS8KN+1wxaWByQ7e5Ejk4HgD8wk32SZuyo
PhQ3oj94p9WZMt0rAw+hgBOiizRWhAjANM7AVJfuHL0c3cninnnHg5GqBmO/uf0u
a8f8+CjKuTBAxEtJ8oOzgGYn54UgQr43WdQpSIgneRi0bqyHnKh67nXrDoNDYS6N
fbwUVQogRpEqvXj6AyNT7wk6M8fKPnZlCfFDQByZ2eIvtuimRUFMhdxo+eRxy9xQ
NRo1vCAGuu9liIbBOxFqJ2AEhkB+h0kOoVZp58pDifgqYxpXP26R5YcYK0keiAnV
FhfoUZcUfrX+1xpHHA4G0tGeLW8n+iioxSFU7X2GN3YD++g6ngsGctEGSW0LFZn+
Dcw4ZsmZcMKioBSt6ZrFr/WNWLh1YTBikXSHPcoCwFzGWcsngTQYohAs6hsM711Z
E1U0qiGPUkIWOwSTH4iVZIHBiHn7zSxc9BD53KsH7ODx+7WXBCEZRZxblmN4dJSF
8KdrL7b63S6uAz9lo7UhXdCgMC6WNOnW0teiKjxBRI5AYXRWIUtxcs1HcAK6IYkm
Dz/ISUEdarByPvYq70Koa0y/ZT1FOfS5jAsCqaMcq6cy7lK3pGbD5YqyFP/SlN6n
/46Xw0gAyS2x1f3qw4vN7lZmcxTcXAyVptHBKQon6z8xKM7XXg5EbulmxY6PwPC7
2euPRzIf4x6UVr7v4/UYSQhF6ZJhS7Yxe1r10EvtuT7hD2K/1AyF/bRmZ8VjMmIW
vD06AWYvoLF7zWV/Yu/JFbD1E/dQnAPf/S/qE2LBbc93nfv1BSzYEv/b0hOIabm6
0QPMIiSFHe/ipWpokvDTYk4yNYFp3jDllFVGbC1kK/65WtHyyMos/BQtXVHxSQpM
iNbpvsJZoS1UC8EvJ6LNEr4nxB7Z17R74i0iAyaeh81GWKUi/aMJu6u/3O/02N3t
WyqMrIKn+/bDulOW+tuoNBCATI8NKmmi7gUta9ZCA3dheZvkJ6Zk6hNpavcEsjJm
QDwcyl84VwcKj6NTHgToViwf1afe/ZRGs6neC2u6pbBrhvVPod24lTNr2m1usxq+
+hK7/Uh5bFLf8S1UmkD1yxWXJwbZPFIWkgiwQRDNy3IIQpDYLZrDHgOBEXp5c/JB
gS1GZVT2u/w1gP+1JFeyPyPwX2bsCT9J2ThS4LPYJBJIJ2qxGYfn8sYHQcFAcgop
TSmfk+utCmDJGJkPWxqf9stGgM5lpfhjULlgw6Mgztis77tgv0O8DSqi/DzGU6KE
zHcYCVpQgk2VfbYjHUbWOwBMwGm3BpqHE2TXvR0Maw3QmdYQWgB7qPNw8hWofdrv
GPAKKG0teNrAxzTR77C+noa707R4YReyyDcsv6ko+Wgw6IgnFxrhESxojsqHoT22
dZUetoQ79ZUbpDONW0vC/ZmpagAepvG95ZCJMNHuyX6oQah+Z/VJpr25y9ryg0LI
w3mINadSZIlfWuMSdi+1VjmggKoFxOy9Eu+rnSMW0Q2RsPtblLzcPFdSG58O8Pli
yUXpVvoXjjHOR0xLFdEY2BRns3RmtXSrrEJei3obQl5+BlmvGwXc8QMEAeMkW9JG
A9dkmV4vRXPywkN+dw/MmEctJoiALy9Edt4gXJQe+JXHKBOf514AgprVUQCoEd6U
1srDpQtKvLAjZlJaUA0Md+9eq6LGMvfsnIR+OG4E1XrwWEji2vulbgj5DYTcgBqr
KmGG+WRQ+3bgEFks29KyADtJTqU4u3DFzv4+85E3r7wc8tj1PpYuYZ46bvAViKD0
9PLF9z7UXANvApEuCrTs4XXmTwetdTVFaOJlncV1acqYEYuT7Tjl3qG7MCHDKVZz
XgEQgVLUe54+DstXy6Z8Wl7D6yR3NtcSQnSp6RXdmAd0b/nYXOwMWRsiQoWGl0aw
FF3GveAfupBDXtS59ikIQW+6MkpdQ+XWHIqfzx6pdIftjaKJZTo+r8zPRl1gx2rv
5cjISesi3Hbt1s+ooZc/BpjBnX/uQd5KFP2vvnrNmo8qpBEdQyAtzuigOl61n8fm
0MOFNGfCHJ4hsZnP9YyQUncOOe3BSGPgyUM8EQTgbRgr5rTH8KiNRSZwPjvLOPzU
HwmJ1FWXgt8FbhrM1D7M8ANmYFxwkHXtDb37bW9zYVkxAnbYCf9DPB3l8tf14fdw
29s3JwpWxq3me3ftDlwsMEHjHy0UKEaw3+R21CK5lpCPJAnqXfMUZbnGrexwiHoN
AHecs0oekBMmWLm+Y/tKbAiL8S7xtkdSx7GL392Ztvn+7tmfFcUMrizy7RnTIJ4G
yx+8NTbhY08ZPZ5u7ssSZQ5HbW4hQnKM8wvx7OTyr48A1TLmyisWUsANf4Nzfwa4
rmjA509o4PtQrlb5TAid7q6ydms/tV4cJAoTMXewhSVL6q+MlOtqS6eJk08Y5O3k
4SfjucGGMyDMFvIAD/RJ/nm2lPaRE33aAlLsAGu3Yvf2hxTDseGBarV1D2tPi2+G
aN72jNMmxZuto9d9I7uMLd8t+N3/HCU03vHWtk0gMWq7Uu464wbdPexPGI0kdkUx
/BSIZW9iyJw5peSnlBPDjvaACvdQrmtac3lXGVKPT3wodyn4opmW3X5YEKbvoOkz
rN6Gv8sOSztk30xzhOyLs/c200dLeInXt5+0aveFs5nESTVslJW+rwzgxw8LwMwR
uKSt/wlgGoebMMRVQictoBRdJBx9pXm2p5jgOUo/W732b0rbAunEIPxi41PKN6Kl
K0F3RKMCx4bOeTvvx5aZ/s+dDyYcTiC2l3hMQT8/FrnMSvEYoBXhIIKNG7PboGjz
0Xx7AlF6ifb/qR8Hg0BNXbEqFxFzy1cMwjfkaR/rz8jvlaa4ns6Zhykl/F8P0Iaj
86i7ucJpPr7bh5mp+C6P44w+OT/8XIdffK77wyCF+H86tKaxyU06Ry55BdlTy9St
N5Dwp0apyMl/BfJZOcHiYWYaGpqbYSpJnoMidHL3fQbYwLjnn/JxCRqjWVj+kdQg
wJzkv0/mulaai1i+g5aOvc5WwAICPMzE74MuDIZ3cvwwnzpbHspLbzNtOVjquH5e
9uoDzBtmvOB2pQGQliAcZmpj7UpoITY94H4J8JWdswMoc5xpHrPQL35jDG8ednox
vq7X5DvYiu8vXVk0Gw/Puf5d+TbNskjpt93306JI3wC01T8i5wZvnXI+caDuQr+O
NsToeXFHgMBS4A9nsk3tyEapZdsA/VJfvkL/4+lo839mvB53CDtnOF1FlgfY8UQV
8XQS0MRZO1j2WbiqL4R8GNMWE0KAQDcbiAVE67mWwR28/eed/eJjb5rGgBFxOg1Y
aJK2e4lv6guNXCke3YT0DdkJzr7AfJUlkx5PmSZKXkmnLwjsn1+2ZxlymR8aA4Iu
AXxTCMTBZB4W7YpoYuMQeNDPXr9jwZypQ+30Dsi+r5nHmSuNLBKZTohLfKsiTNk6
1T3PwD3qdaJYumXd4pK2TVfq0RNAqe5WNGXo1Pt/YDPrzHm6mRXc5QcrOtIki60X
Oj5VWN1q1jOpA5+Gj2XzGu5CSGY8STRqEKaIF02jajToTmOmVPBN8wypq3x5gmrM
W30+BXUxPonGRxCZUr1+22LEPyQ6f/lL0wqBEI0BVWk4ogTmlBMyH9KQfihjcI+l
zpglwtx6us+kpedT+XQCjlN/qDVhvDAS4K6i+d1/6phtR3bOqlf59wNJzRmVIVGp
WGuVYp1+bzhiT+nvF+h9pc869TYeUA3AOEu4dw6Agsg9Ba3O6WQDNnqH6i/JPnil
JydgLcPsMCe45Q4MpsvxU4uvpGEuwls+9siEBDsbjFQkYfFlIjZeDKMrxtGAKuYW
J56yxX8AS0vSCfjHxQEGkBgB/cVqxkNLZKzXqah9SyHxV35ZDGSITcfmlSAgr1rb
W0hF2pq5syFoN96DFSlzlbq6QPagTvZM8NSnYMEhyfrGIDzjo4fAiwwmLYDvZsUi
Pg+ugQohv8SZ0HrIFoEP/wjZX+1Ma3pRzTwrfPbjNWDK/nMLol6k//J8eZ/J6eoW
Y1PgCo2VazremuZTy7WZwlGhlfuOU1N1eOwLtZnJqrYMMqxFktePGYNhUGi4EYMc
Nf3Mb2k2fQl5CRhEfkwCi+YkxfQhTK/Q9hEUjHEJbaOVkFAt9c0C1Ywc4fuKe8x0
YFR/kmCKxTgmA0Xm/QOj3Z/5dmnkgkce2yNi0qcDa183i6FOXUOUclVLZ6mgZgem
FMfet2Ph3/WCPgcd8MPRiOkusGl2S8puNZxnQDx3NjIV0JRbGSYPUhR3wDFsAvQ1
SJEj3alK7UGRf4PFrDYStAxz6RglfyFi3hxO60UVtyCLapRap9GgNlgXgTkeMkhl
UNZpQ8qUIj3NrTs35IW6lEZqvYtZoEU8kNanJUU0FCJdYW6rigfb9968ZpYiFJQN
yd+Vt15Q4a+Oz+840dJgq14XCEztePWU3q8J3Ng0ekw3+o1+IrxS5d/mIFW8uTBe
uTOi9ICUDur+ZhgdPMlTh9575SjEnrBNmQwdnif1+nO2lA54kCK1r3sVYu+ia25G
9RbLiHBtcBiOLATfVl1yRBP5SC8M85d2VobqYyXyJ21IyhByNNNZOVhotqkbHgSk
BUHx0MKbPo4HoiCaBROrOxPHA9Bd4m+eZeAYP6MOvnqY0o638l4vd4/fqGg+m+Xc
fN54gTzsnjWkKH1MM4eZZc2ob9PwFMz9SD3IN5Fx8Rq/ZDDA6rx2WnJFQ0fLFzsf
63dIpJeYayo86NekttCXcodfuA3zTwhiXr8IKpbWHqDmJg3yNL5VNa8cSr+qEn5I
idQRXl1aPf60XyY5diqDXL8KeWmkcBSXCuaVzXrNAgCE6jqPq+UezZPFTRjl6fm4
S4P79Z32rQyU7FbQ9D21NFiNVovUCbsQYDWqcHj5sZ/PQqsrJ/0RNxEXWjxPfBg7
jRrHope2nAkV7/rbZpPJsuqEoQQwPwoAIok7VKZyD7EjKGG2f0uvXhcVbLEEOhlr
qmBkJXqdaMNsRenF3hqDdNVrWQvAkvXqWE7AjOA0rowS2KR/9BRA+SJaZVwhVzcd
u38HNhr1oCAugMWxCqeh2YHvKXDjOL2UNbxlAqSqLPz6SkjkQWTw+M7FPziF6naK
hd88OBv5HEJDitvo/ZRivNa/gDCJINBBGY7y1jjPsXeAUOo1wKjvexvFT4v1FOpS
za7oJ6DrIixDZ2Yh06iqII47kOfanb/xc627S01mc7G8M17GsazrrU3lmczEEPbZ
S3DFjNYQSuAun8KkxZE+WXJ9LhVddvKc2pO8t+M4+nep1ZM3UgVhFm/r8yqWuD7u
ZVSCDQH+cex7AvC8KiIbW25+oCF51+HTrNkOh0Q+DP7F69FJJXF5ym7mYCz5+fVu
iVsBQnwypeoSI5cA+VQYHx1Jg5dD6qZqJDxPeKn+afaO7ZtLY2LxMf1KEzQ7qHPI
XhiUXIS0AiQ/Y9VEPn+15oIZeX2teWJuvtJmWFsL0fAVNXJFckHQZgtszQEMUZc5
fQNIWHZOMdlAmKxqL/IQmlVcN6Dcs/eOo1B1tgXSPhwF/1AN7qOZzua+/qZI4kIt
GD8lsq8BPc5HJuz4oWWcB5Wr9Fut7jZLcjkIDs8xFZl6H1o+X46IXr9OqAufxjf7
Qr2USJ3MyDbepNjSsQCApXNdUvYMnIdaCVYe/2wru0a14TgpGXKsIqpvAaqiAVol
Nn5pHgW9jZ7WyDvhR0P7Nct61RL3Ba6QXmdZGHlXer61TI34wUuMuv9b6+r+4HA8
8N3ldb0rl+1ERGgvGDLzi7ChB4Cx9K5lZbRQCpsxS5aJZsVWJLnKarPELrfSNynf
8QFu88OwBQ+JN2oTKTDJ4NLiibpqOaHG2NhEGcuX42pKZN04xgyvL8y7dqWJxdFs
rkI862+6yCd2YQNo8eJZo7HCtgN9OXVZTL2w7hjslajbhPhp7BmfuTHdCgd+XITB
2ezskRMTOlwx3AAhLysxoyM/6B/0vDogypReh9NY3JvUB782vPRJ0JYh7gwDl9h+
SbGgCksRZeX8ZlIjbKCi6Ihzz7OPzFGK0KbpcKz+rdLstJFP9PhvginjTkEhB/8h
+wHrbKB81jY7qYrr3kOzOceuaGwM5drrMfk97+QFgu5PcOYxIYLcPKi3maVRDKcg
Uyv7ZWPFmzwP21e77uRKC/RjtnROc2zFNN4dC9EpBfUu9Ik4Qn33oO8nSnNJnPDR
th/PTE+qhJI3fqw8PjOmv3dAjadnKsXlXkcOU6QFjdvstCfaqVlIoYCeh0tFPpKA
s8ip6Epl6bD/4TDOulEjuow7ED096I+lKmKYoqJQJ5ivFgVYmxwbbvjbz+F6i2h8
J9GnlAH3XfZoIOWSqyAmvBkHzE9PqUUTZh+EOq2R19sMJt1HHz/SQyc8g+zmYuEq
RjjUWFXLVXv9twUzSeX+8K3cSdoibF7CtvCzYourFNkMwR4k3JKx6SoOK/KhSd9h
BhdVBIZSi8qqIdOeF6vTttcO8f+aWQLcE0vYK2eENDvJxedEk7N7n6zEoJuR0n5T
uTKczA9niSylSH5Jq8jXbXY0dtXUKOKfkgdOSj+2yKYB1//qyyPg2PkOE4kh/uRh
86pj4gAu6fDb3uEhDepsgffI2pWnRf+fGrqSUJ1FGL0mUHF23IREAMTo7pjUDHyh
MU+FMhi7pZ4AePcrbabhhqrHT8/pmWguU/vZzDK6+vjksk99GVyplobt4b7TEQCt
Mz5fV3phAp8JCR4wJ+UTFH9zZry2NiMU72xuRlFk5/BSOY43bIMCbdjyoW9ZjrHr
HRroMc2bGVRgIDn1T5Ae9V9jzG1eekxBw6iGBEJChyts7zwrU2yh/TBPlHfFqsZD
QEoN3s2KfyQvMmIDDCfiqKf+W6S5s40jq7kvBThZhF/HY8cDYSzAcEE2ZtgGHoIT
C7ga34X98h6bmF7l5tk4XoOqVNBDq1LDzGi2uA72xGz7ML7qpmKP9Jyc8VRMgJYp
hq6AzzPCpQTtwWRFFK4GvJtqcrWGILJ5+FDUfAtSJN5Hwiz8DTDh4llHMSMopjS+
SiV3iDJNIJlRFcq01x0Ub6vy3FRxPnrwJA1/3sHnN+/llsqn2IhxQACZe0rH91WX
pQ2gBykH0lhs93sH2l2UU7b7rZRXQFOK6BKvyoRGSrq1qF0tDG47XmPjV9gotQXh
O3p4FSYhaSfRdoeShIX7H2XKwKaSH3sHSjX0XrJDEDCy2bIe/tk5k5IUf3ZNTL15
hvyf5AKipA6myrUCLxwEcTDoye87tPJfp98MwP2MEQzZ/U0ecyi8wgDGVcI05ncs
pW/5idgY4C4xOKWHnTHluGE4r3MdqG8F/jIXIGVMNdajmedG8owR0EQNm22TgPLG
MyPFRi2SOQshGg8OT2xKdPn7nbl8gt55frN/BUcdY8oy9bB3Me3PLbs7yXuncOTj
h6AcG7HKlwr24FyVaJ7YXe/6mN8s/xzaXJc2WjxFbSlASldvyllQ8A6h+5Cblz1I
HCN5BGVztSSBlGWCdtXRX8R/jWF/f6qHRq6uWoB/nf5y3JwWC2iNQI444I8Jpa7f
ZxdQ/6PP9R8+T5QIGa2S2e5TVGUuaVLU9ICikhtV2y2MLoE7kZn3iPEtPjsdrhhS
RT7euaGG8K6HkfEJ/9VeEgH2YsA3RXgWJkV2E3ATva6fiKA/PZKDli6Gs86pS4mk
2Uk95ViRvZxyAGDxkNqeSqVZI4gG/iFEoUG5DfyB9GAxWdJ3bn6K2+O2ghwELggr
l+b43PW2i15tVPIg6khf1AIVv5Q1t9WBu5sALQ7Sq91QwuxNjgI8+4MzIqteG+Mk
6DgxrRSZqwAoQ0cQUEodBEtqX6wp9sjjT50/xgpQ/JrSwL4DPzBNYE4bAVs6WBzJ
gsxFSOMetYEHnrYTK875GGMHd1KShiuBB+dWjs6bhgegDoo7qU0zOFfNzB0AJWuD
a1sNuC0s/PPO55zgdNWM61CLfCbrP1qiigspX6XCfjiipE0YS61UgHbh9RuwL7cG
ivexsYGsTlgUDvwxegwRZqF6qR16a3lYpqm0TeJ6ns4I6zCcfsTGQ/xogvSnGXHl
G4boKez4eogrojRWWVSbCXGYbEdUWMjzdCjmW5/92BFVYsB9syV2wCbqrSIhW26F
DlYxNr/y78PwkP8YEOXyQhsdkJlbbai1XfhnpQcumk2evudUsRmxm/zeiSyRm5aE
dnId263xjgFnU17UJxsOdA5UX1hrvwi2rC7MmF8DBv1em+/URWE0+0347BhQeDuc
iZeWu6Jy9SvB2byjErNKTnXu7rCUmOnkSQwqkG7S1h4dUNbBZOuw5xDhspnR9glB
o23d+jPud02VUbpm9NbUpxFbZQ3T3/w4pyf5xwwupxC4uETXSiaywoWCeShlpSEA
0vG0i9OJ30NB2SnPAJSvHsYxtN3SpNxLw4MTGl9ciySO09VM8nlyrblUq9CyvL5x
rjohYADb/WoN/lKgRKGEdf739036LE9SFP6M9nl5ij9DT9Dt68LguFRDnUOB/pz8
QzzKRbJNGtXh+Tp2Ix4DVdvYIYALtZZquSkARr4QMFHNIz67m5DetUsxBUUHDEj4
W4adQQMEUXO19ZzUAgwPdSC3HmMgAA+70xjbS23SUq5lbxH9M0acCEm5Z1wdCaVd
Mk/TrtnHyuvtq+pDt7R1AXDhaH0gNC/FvavmEngLJzazFuvzvWgEWJgnphUdlz8F
UZc+fbBlLMKdXevsNdZ7iDPTIpa4sPx3Ur3MSEJTO6lupuT59n3iHRcDCeIiGtat
rFKe9VIYmTFPypunOkf8MBALUcgBnnMpVPG0xjIdNElIhaDo9/euGbFM8yyDvDxU
07uaFoi4xMxDU1e70snXG5Y/ZB/oKuRQHionD97XOFSNdis8LQ+dL2+cLfLpD+vG
BELlRmFdiwwdseFEhn8RvYEFVGpPDKqX7n/mG+8ceA+tkOm5LjSd8aphQBLgQ3J7
5IQ3MlGDFs3LzBY6dFVQSxNCwO8fGfd9kbRq7zWUvy7KFKBgleVQ0TRZ2dl72wle
vN4P+aTMoYV45hKJqa0NKCzFQ7LZ5YsuB8k5kQ+wxiyfFMk6bsEoZBGX8VBtYF+e
CCFSSGOvRSax1CYAU6LFkOHVXLgDMsJv5O1TarR6/gIyfYY77E9T8A28TqwjLHjR
yc338x0yhCeNcx8HYSQK1r7eC3mp7p7Oc8uIkVMQlyuCJmIVyftdJbg2/VOCb/Tm
WsAdbvPYvKGzEWkecP8wRh0Xjt9q8O9q6yQOak3GeWEoZJS5RYIeYa47c7CaXKJC
nH4koPPMtvRywjLDisfdYvTCtqxMIDyCTSFLZHq3zT1L9RBj9icOTnQ1EXg6Rdyx
zXONsx57KoTPDwDKyCpQdeIbxlqBR2IxfhY7D8r+Wx5kmBmbnixO5yMRyUakUboo
cZ5ifH5K1ErgpXo427BtMGxVL3LRTAm/roYy2Vvgy4nYgATa3e2COYd57GeT8BDn
fNTNdlYRUyNcyTPMBa3AVvJrkES5+KniHt1yZ+e1LwisdcZ7aQ9eVrFGqhifx+5n
vTVFc7okC0FndemJ9nyMar8SfScUDSs/1tywatXFJDdsqLL1pORkiVQTj2CEy/FJ
CHyqZXfGMMSI7/6fajoh+dMQ2bcTjVEpFXaGOebdyGQiR879pBv0Zdi4zLws1klm
yjJ0C1tsSpIl1p/7hd+9+RdV45AktWV8yzk5bkLxgt+//Rxb9NMalS8cup1G7AaJ
Z5H6lW+p/T2u87FyE/rjasok17bjlQb3zW7lFxrAbGPbPopWYtkKQHs5nLQ3/NNT
oczG0VscqBu3j6tI/4vQQyaGeRjxbkoPtL8vm43F6li6TxgPJifFAIshZl0OWQhg
RfgCsM2TCX9TujAyqYj9C/h69qV7runViXDG9X9fhXqh5ZHbjFYcS7PEEK0r1+Vk
VdEll/M4JsY5gwfLmvBysyQLfUvphhX+hWdJj3Xz3SIe4YdhH7mTSn9pgolBNJWT
Lu+njqKwObTESE0TCBL+8qS8gdDt7dIOayGSgocUKp2qxpxKWppZQ5/s92X6dXP7
hvCflDlOElCiDnuLZN21hhTHOFXq9I6sAJjmJ8glvvae6ac6SmNloS7yFul17LEb
LFYI99nVH4VbkesvK7cF/u5yX6Sd7HxRF3NFkCVtIRai+q7FBP9M74YSYjEUT3LY
RuRjMvy2mwGBwDrf3zcEld78+8/MQ4N2I2ejdfGgezSy7ltpTl9eGer+Keif8oml
IjdYV0eO1ZGW9dZt/e16pDoBr4RDaXNHYKShqBi4bnhF04twZY5hbN1RySGBlQy4
aZQ+30UzrMQVkofDWOweA0t3m8gCONKy1Py2JAL7K7CaL1x1+FMSHB7n+Rm94aP9
ucefyYiR5BLde8bq2DGUv69zZsck0P5ZSj4h8jVc1GInTDJddhuIAFR2SJVN2FB9
hjim3Y1NK7hTMHTNdHZei59a6Cw8k6k25fGN4Ynlx6DZJyKhuWoVII+uXuQJU6/d
/6vNSuqzGxPwuBMffqHKVkcclTKuFYNiWa+MQkRWyz4zLm15OH/vj8WNrgRlMZsx
BCz7D6mr59/ITJ2Ua0EzrpznVWyFukkNupmCfeg/GVe2PyOL16da4EvubvGrFUIB
pOxLzzHwl3Lx7iNrsaONyWrKXc6GFCpJpLOWoTzRSl7wzCDI/eNJnEm64H4uYzrm
hxBj6D9/9b7L6VAqGgEccn9ZUQ6I2VRQEdU9snMQCjNVnsz6V/jRn27m/HNVfd7i
xf9m0Sa99X29M/1t3W67FWKovW0g/3Mfu8uQPvy6QucA8XYyFOeLREuDFwzCdy4V
ZwXrj7GnhCS0AkAKWHRnmJV579OW2/sJguoZ5TsnsYlIS8QYJwBFolGRuZcQlqgi
LsJA1TP30u3VSXRc6mZQ/z7tx07O7HheR3PubYgXo9nCv279q4O1ohNOcD6ftNbE
DXroGtPdw8NIEGPCPLuFIckkJ5p7pcTGYrS7+3CplNOtNByMBoMEh4NWbJKcwPtu
ZWW3+fuk+f7WgPSF9gkGyd9KChN2mE0l31ibXZmh1ViI1Gl0dPc1DUipmXSdWje+
GDdhGLU63C2X8fZwIzz4ofPVZQyjFvp4wmoe+W2g8c/ts8BHjhMHnd7YqZ95Th0m
dI12HWabz2ZKKcbUJZPBuh/Hz+e9fo3ZMw23rVuE1wMyzNW0x0Q6VcD/DZ5EISq1
IfmAFGsbUc757JBcWvEy8GJ2zsmfWWhBrcqnIZhA0GQH/o490yfNEK5+dh6UHsUz
NLI70crDrXzdYpmqMnylVnOnMHifDNXAYoAPGX9qTqA92HPweDT4Fio+s+ywr123
FSM085eYz4d4IGwIKNviQa4lmvfzMfrhsHmnLXfCforNkTTlwykYgfC6/lRDBQgC
gEEFkNPDMNqF7kz9dveqVa0e7rn+uu7K0XaKlhBpEmddb/WMsgIhZo5BmmzSPIWa
p7d4BWfqtevfFHetTl1YLeN4bGmDwbmnHO5d8m/Iv3P1v7CTwja7T/cbFSG5oQKh
Cvjrsz4LoiZWJnuaIMopISE3cZlpG7aW1VudC1s0UD/JvbCWlTJ+0gDWGBNbepct
B14/rci/XL4XgxdIR0E73jZGh81/z6ws3zV6wd/guEkVNNIEf8eT9vTdP0mDYgTv
qea2YtANEtpxODHAw0v3alkz21Ok0lvkbYrRfnG8QGWMDcHuI30WaWNLomd1nGRc
mPRACUe1JCCvZNSw6WoXQKQWGc3Q1E1fj+FpfZ9E/NKJLz8rqkKoruN7sOV9ldHd
pXZMwIrGlGq8eaMOFROlpw9Hbqr1x0Sq0aYrmXTLfSbjxkBRhFMvyjgsmZXl5Cfj
6mXaOhqUrPI8lX3YZSoZUeDowFxK0zRiJR8HF90CBOM13pJwhTkBmMOcANfV+9/S
3JfPzNz1OdTOiGH8cUx/j3CidhxHH6LCdoaMadB4TgN4WYQ4BPo4IdWlZPLrvhJi
qdxk+gzSbUPlLEqdaV4q/Qg+EF8v1VOohIYtQ8RRmY/ECEQGOoSD2QBe5HyqdDIL
eCnZy2Vm40E1gmbMTzZ6k2RFb86WojV2qrHWukCJQMoEWum2Lt6kgHy0s7y3kZjH
qP8L2u/Gfh7KU+FDawxDZqyd4ZAeYE5tq2X/VJazJmiPnq7wOHmUv1g0QGi0GRGL
pZmf9Zf4sS3bS6q1H6pf0WVb4v99lNtRvOudy5UVejs8AQtUa/MCVTnQBN1R5VEC
8ojROCZIP+ujOMhIyHyKDhDz0JlrLXe51KI7I4VUC/lwE+hiO8r9Xz0cxr/2c1TD
gHhlyxj3Bpdq0u9Sn3JXmCmSpO9Yjgn/yqpI7WmypM8hyKgZ2TW+DNzP7TjUk3P3
RDTs/If2zDNSakjDcEqvJexE/s9hYYv1++yfv5ehklUjnU6VJhIfgUZXPhjGERHj
UIqINqqnPN0Pu50+L4l+ddgYxWBAuxGe6FS1eBs0XNIzvRGdcVBcVNQ420DPO6Cs
M2rLH9c6JCHfQE+FEnOcRpl75aLFyW8RyXAGk7NizPxOWnsr4zJnW9nqjm1GGUFf
3mGiG+Kp8JG989hBvBkqJugAphp/mLYPcl6j7Zp1gbBVf/DN9xeJ9Rcikq+bWy8u
ZFQInsb8CtlG2+OvsFeaLeh8mob8NBtR7DKSX2UNWQp71T6BytHBYbcRI7F/Ej/A
tnp6mZvrWjDCsnGhGjTKb1qCcri6cCSKA92pPtI1yJaTTeNZ2KPSziUmSDBlcvkW
b/W+QpzXIFxnSfCiSvznBXJC5vq5TjefVXf311J923kO4aRNvzf2N5gtd9wa+YzP
xqWh2SK2MYQbEHIMnRkKvHbINHiQePi0dPuJUYYHB+y3l1+kX04ca69gAEfpD8i5
lquiwm1UE+/Sfn7cZ8/5IHEhbymi2Fr6fr31PvKqMOZXhxZlQFR2xbcys2pYQN75
lEZ8T3AKZEl5lIebI2C4L3uM8wgcpOzq8y/owkUdGL7PipxYaCV2ag1xea6aThQV
eEO66oz1S96sg9JLCKZlGXBcImWyVqMZ4vdvMe/IhWk3H7+mYVpwEsr53uAKq7Mq
XjJc7/yS3idXRCSxPfoYCbx/bWb4luBmLTXfD0kkieurcVjdg9JQ2TtguzbsFnSr
HN4HgEwN1AoVyLpr26wpYevuiC2nCsv87rYq5ibQcTN3nsOzv9r+z/j/j6m1Z1GA
N+vi/zxDlLY1NSb3kL3qW+JNQxnT339/NSfMVgabgfLrgVpFCMx9OsmAfc8Yh/Ui
w9GJs4S3AnGaDfUpPzdM33gRnQnMAMEFT7QSOAqXtaPdSvz1m+HonbUL1Nhkx6Xe
sxJzLHjJdQ5LxhSWlAJWaSUMh4W6WSZPI70N4U/jdVWYC3g5e1jhdoiyyJGtszQR
gg8RrmSfuegu4SIWhYTh79+CmvO2JfOhT+/DfqRO/mH2IlutCpNEtGak7A7XLzgY
3XzcOCx7hgtMv3ql40qb264bcBsBWDJphMkdAbF6qe8PbqSye8HzwWL0nWKMsFWg
TXRMtUIM8S0FF+iZ8WSNs6wFX1P1dWdEqJvUI1Pik79I7mfq/Sd+QjgymsMFmNsb
feodRMoKDie3eze2eh4NBzgCgLJcjYSLNsopOcJIPLYfNrqkHBaenbhsakyF+Kkt
SIN2vwjUbbGmrNKi0brFcmW68LceLRbTwbVlpNXiquZgxyvfC79BnLxPnil4+s8t
xpJng0CwR3ki5kcSxu5GJ5NzSKxHlHPLasYjvfRmwhVItt2d6ExHLBnqgMczqcv8
EgIQwD6/mISh+U86XUwKFSmonmrotmhi7cNTyqenx5biJbhBO34puLJU2yjdwaQJ
LZBGGMTNJ6XzLy4wCFroLQLQViHckZ9FUhdBxG0xEwHRl975ercdNTVsqAt7ceBL
3aSPV2S2sKWpWhg1cocVm/niD9Dmyb/E+nUxkjm4PD/6OEtm9PBer4QrwcvpzG+w
SUyyoyfI8Nq8aHL3WMvdV0hDKOWZn+PTHDu/KsaFuUEPIrtvo9DJpou1HJhHroVk
BLbLypzawlU6S2dh0OlmHhDXIOfKia9lSyz8PXvACEJxOe9mdrTsyy6CF2yNx5yW
zp+m4o12LPfQwZ8H0o/DeH9tPu5CmPqdjklDaZCQzy1VbVzMgLdDeZVn7ySrLjb/
0hhGWjZ4+qCHDFPdPCv2VBAj0dw0KIZzcsVxgx5VDq8/vuaF46tgoeeEF7Ek57RL
aAop8prkR9e5ZP4zqw9A0ff9ROgibz5RrZPQdnhtxEvBPiycezSyIem7BpW9DG0w
uRzTyaMfRnjPSIzrceGKskCSS+M+p9NhtdwInmbCzAFximKKATna8f4if97i5UCC
zkWPqdCG8shbaFTiOwIzavFwFPhqJTYPydtNAn58O5LgWoXI3m18+1MVWjXx896g
csBsg17M9t4mncb2/a4N3y3AiC6YxapFSPT87wvUfnGE7FRTzJMRU2Em2g0gMIVO
BZRxxVyzithvXT1Xz+mYI2e1hOvh5rt9xjqxPDm6k5NNC4evguZqwReG6qJA7/+C
rvl+fSdSPP9ysN2HV4JSLFMsZuMncqpFjolQnkNJP0TQvLUBMtNvWv3szNQ132Gf
Y5Yy8E/PbltnnaU2lerduPff3gpNinjglpTNUNvNmlEkiIkofHyP2RO9s4nP7h+I
6uHsXGA95cy6YWJVPEH+NFlRla1y1LsuSpHQo+JL4UYLz4AMeN4Er6xErA/aSzKI
7tt426koords17+gLX8p5K7+AmWGhmxNkORWTy+xtzE7Tf83jd3hs1BKPyCkdxke
uFRsiFcGVnk17ySAV/fIs2ookYbgBFi71uiypJKkIhJxMTPlXwGvyRgyxC4L7Ken
Q69jop6p5mQp+d5IlrArA9oIGbbeLIGWapl0XsDu04c2SLSaeIYnPdyFjWoaCNwO
UZ+M+KAmzSV5HSzj1vxO0Yyii8SCeC7Oa7eBG1cIJlXQqmUZd5pjNPtXoE3yLkwW
Ki6aV7sqlyVEC+f86BVo8t3dhrA00D2Ekuf73TcHPz6zLIPmfNl0DKkRqVbYIt7h
guxKVOmVq9uVFQSOBThsBjKMcatj+xdL3MqjKIxi4/t2G9w7Ummyqn4dzvgurDFi
cY2+/PdskgFJ/tfQwWNAuZPgOIUvrkTtn0nAyCn6LifeHllW9TM/cDmNOU2Pxb9s
SosVWDEKlsOUMo9f+bocVX4JFmDisFNWF3RWaxfUdE6XEqSL4pylc7YYGP/MsRLD
XSA6OPdwKMig5tS+xhra27xYPOkcCQ51+UugVK42qzDZ3ESZCSUyJ5vOcZN7qGnt
g6GUH6vzD+xdqaWnp9cFMPg301R7/2J71U9tJ0yCNNsj5qUthh22Rn6mQ2yGC31R
Ma6btyWW4L6evQ9J0EtNu0/42+mQhQtKaXv5i+AJ8xOrK2SmG25ZVy7hwCBLD/S2
B0dXa1TN5a42ErPmLctQhnFyhDR56kn8lJwUnx6Az7DnK/ZjkXwLjaQYiXa4BOB9
zMqTjm8CfNMc9/HTNuNsWKMZtjh9yA6gMwor9uTX/WNJPuRfebwTj1uVKuXLjqMU
riatoYLDHUtaAweOdNs642JbvatXnEgyiXRoE2QgHGLAsi7VGDFqYQM1T2VGF6hC
TCOQshNLBShKvSRjomfHUv1ZBBJJ/VMuy+F2AWKeXmbQliuBDm1so9oj/+mGzL3R
ttIiu3Rb4pBOXvn/JVG+2ivBIRh+eX0FggQ2b4cMwCtPjIiHkIC4+GdD7o5BmQHs
e2FmzjZn+Rk4GKaL/KuzVgmrxaf+rv3uNnY3yO5p/g+XxQ1pB5/BActv0WwU98fS
qk/lxMY2NaVNAPva+MWd/IwqQw2YcXwf5LZofeloANpAfMKWj8QIe1Tn+AqLwlNx
ScDRasRf7jBiwhIPuvpf6EjtD5iCTlWp8rzpuvwCUoeSJqo4qJSVfBusiufTAfcR
jqxzPgW8SbI90BbuICqIHV/5fkBwgv9xh5MRwPlwxTbtPJJGop7ejHfZFqZHhSog
3IaCn0L78cfsVU0OEj9kd8lBQ5fOAbavZ1Gxo2MHF91Wd7m5b1bGLNlsRxuojvz5
TPKbumUEf2U14TtrjS+s7NLqpS+iir/IefXjNnWOKgw8rxowNQKhSqALiEYmTXpm
+rMZ1NWhBBwUT+0Mw0gMB+NA51YqI3uf7Jua85xZTHCQFdr0Z7vFMD+mnUdUqVk1
Z+63lwVRJR7ePk5zi+HNeFID8dQAG22edtITOCHb5UNC7iTWuvaaECCLi12kJIEG
vJB4oUo63KgaaMV+77sx+1pFqYGBRAQQv0q08ycXUmG3Sk9xA4dEzhRA4ewbu1cf
6OC1C0zC63HVjugcNLujvj7+etgtmMqxfec32DTbC5CBZBirzea1psjN2XMQg7l1
BavID9PpJ13TKvEIepA14VDlQupPTEsmg4BtlWHDs9COwUJSzFQ8htXwl/sGu0sT
qtCaE2QEjj+tZlMjoTrlUt/wzni/BjEhDVzyWdQb+TmG6PSK/tKtNqFinD/3D8fd
jXsh5nMworzXLA0x5/8pIz7xRNm56EDBKOHueSsBvhZBK/fFKhNsHLO6nStN/0jm
30Mkpl2v4ja45vgOYbLJWcoWbokiCgWKfM+OxIrjgogQ2IOe0i7uxfljIgHAVP4j
W7zcIqwgPkvA8mKwo+mlXtHRSuSO3hWD2Lg+/r4obDHQAIWRAmPuZQ7AKeMY+ZHN
38ovo4djF2f5VGphpUbqxnYmfozYAIrDswHcD8cKkPOmjcOq33GetDRlagK3PoZY
zJQGJW7TuDgnd5MrwlJ2DCQxPE078d60ltCVyYy9uYECHLeHijpfPdPX19O5Trii
F1JSmkrYAboDnlP6pzDBLz+ZmzL3stS3YSxVk2M4upahBry3cRoya+qaKqremnCU
nifxccM25CZU4R/foEJR7CH2HIErnuIsj6w2mqxeEpwYTTPr18L0DxCCZcib2N0u
4lGQzrfDprjFQsEjf64P4TIpEBNC1xAP5BDR+ErWil7jUWqW1TyjvEm3BoAVB1RR
olwawGEpRjWxOeTlichmEQg4HgtcLuQ4HBBDnPQg7oR3kVfa1aIZaUIfK9IlEF8d
PxAirAnnZKZWy2swEgYkeCSr27XuEXpTWLcdVX9ZtvrM1ZojNFZ4b4UHWuna9Gun
6/ftbUZEJ8bLz206+jQD0WJXr3+d8It2iEx9JdRrjhtPQbR/MTDcKY7xw1P/TrfM
jJGsZ0RIHNvAZ4FKl2cnQ7aL26AZuZIqxYkofA7SBo9jHcbQdsZJJlGzNHk1nBRf
KP+FF2vx132ufQ3kxmK7ghStJnzybNclXocZaomhwPsO7Zrd++jlrr1XgZiOTkqw
nd/6ZNzb7OVPzMQNCGeP7W4ypjijeVH6sM3ayGQC5tZZ8+1b55nBNW9tnYHWzDfp
yU5+L0bCB7/LQsUZH153CBe6vmZpZd6Pv4ng1wr57/krEVYO+XuBp7nvBEXMQwnJ
naTl2GRPAvIeDQ6AKKDKio65hq9slWQOMa5E2suPaT9W5lnZxhDoeNXjW+0XjTsn
zbqbLYSzWAKIYb7abAEg95tFlLWSQLG3SbEV4zzuky7ohSH+oqfPvXTucDi28xpj
zK034OaCiK4Pa8DKKGPUqCGZX5zl0U6E+h9SEwng79oMwu0lQheG1eaqM8gjaD6T
3GBQcijmdrdGcP6vjPjVczMSino1IwjfMYUO1CDQsH8+SGJUWzzEAiAOSZqBE0ID
VZelPd6tzxfnUbhD+lhYEGq9dGD4EifiO2pORAl4kwq5ww9W/sUC5Yen2jr1N6LC
focE1h3XRSJeAmqTFhsdLb+9IFeqAUGbyIIk6CIfGzH8omfO/hMAvezwDNDZbJHo
dJxJNuYDYAS0x1BR2kTlrvtOahM3hdN8LDFOK1+3982mTJ1JXA6ERs3mOxDftE/6
r2y4YVpC4MY9cHQFEBkwmPqKwJlWB9iOzp6qzP7s8p9FR2v9cenrk15yBiHXaaYk
EvQHHa9oQ4qwvczs9GxOdSSvegAPwh3JhMa94ZOLuT7F5vU0zFirNJ2GEmnByA7f
85KQjJ7A0eFZnFySRml7oNrCN5HGI2p78BWQRhOoI6uVJqJuol3Pj9AbiZ8LKdvL
rFVySG0f1tEHu7u0r60rRXc8TzusXGKQch/mg/94qWmeTx7F9tn39Ee+IanRPFf9
Q84nZng25gQYkLnCvu5nu3wz1bCRGa/2HcLBAqecm/ql95/HblSXsgQIzsVWvAA8
OtUsLdzSmrLzKoq2jcpf9rxxVShunPS2LTM9eG+CO8j6a4tNSicknJ7FRYwJ/vYh
lSAeckZIKsX/V5uYXZDQUij+fdNQzNcv9YNIXmakBiMLSOeQJRApLkltICyb3g4U
+7mHighoDX2qtzDFgpWeNmAgVVR9Wv3a5ghRlu6n9bBrbKu5iTZlR/Q9PQ5RqWrJ
mO/rq9Pke+AnsaFYIFkPYMLtaDi7U5D8gBZALGe5AaBySUt1XD5UWSviQxy8jP+p
s5jkm7pGczSSfp7/WjjyBF98iDEbMZauuq+luGJdnzAs05GJ9rD4CBkCV5v4WfJn
u/Fv7tBdESWUvpX4Q+Jp592HE/mRNsIxdkB0xt5LYE4TTcjEgEJADTswaKlGh1SW
+9vBIrv3Jt8YMFSQY+dJHD97KTT7h7CFp8Nfot/iHTB94qLT5L/mKwCSZphE55+y
++Sys3lEwwWkw2oIZYfN2GjNBMx79OwqiyuHfwFMcpjPyHmDpnOfv6ZKxQ8Uyd80
0k1OVMgrWLxWOdVFQBhpVJW1XanWeSERwcadH1buR668lnUASyKHg1QoCuLZ8AX9
GCVCkiB0/7cuNJv2nsbS8f0s0ezxHDjaGf97XyRoQugPP+prA6HRzf3Fb8kXzSw+
Bbsiw3bfWHNxALfjRgr0XP+IfhUaFVXsMrIevTUZkTbMbmXY8a3DFWAV5uz/NyjT
U8kP9vHZvEIIUAoECVVV14ECWrbvYsK0p8A6n/FTBUch4k4miBORBhUSzkL99+3w
6w7RIUtcC1cZbCBo0NEgXRIKgEr3jUwzv9LW4+JP4sQ5J0qPyiIegHdp6RoFRA22
0IZIxWrCMDDNWEUlHdUhdSngkVsi5tnOzEYYzZR/YnPuDVg3M/ZzjHXsAj5+a9w2
JpEGal3j0Ha5mVQSZFw3Jza9dbwCV9hMV0KcUlelglJPxZPdVo2BjohPyjdhUBFg
a0dHubZd+2rDxjuptxkZ/b3m8p6v3oH6frGEa0+3VJotlWaWas+Wx+Bnln5cFTRc
vMkeIAS2+1AfZBS1Uh8Tlt2OQu8PZ5MbQLndRe+8ohtv1FbeGc5tsZBrh6MdIuL2
ysyPB1JYYPvfeqzjilWEhcMYFWJVhA698rbJ3zdIdI3EW1Z0+Z3IJhoSo+breW9i
d3rYMuHj5dD+v7MbwBf68/p9wI4wRP9IxSX4lzUi/vdFigo3ge+Uj4ID6n0bGVOy
YCLoUYHBzgIJf521fqghK71KfvrOb7ktPceW7m2R91PPjoU1eDuk30Dk1DF7ot9o
aHWnG5eJwnM/RxH0OcdxxltF/eA9crws71Abrc74oUf8iHpYb/J98BqCLOCJZHIb
AD62MqEF/wSdbgkoz+b0eydbwY0gjHeM98jRnuVim2QXHqwGphr4QG4pxeCC3P3Q
HmQj7fqBy1O132M2BrBLaCOT1BmQw/UeE6WC9DMEmMI7pI42c1T8jGN2Ja+0F1Ck
jwTNUq48UkaeamwqAoo2vEGHJIG7oZ8ee+NATrG2Rkt2UNdAr8IXYCFitG8d07cq
6dJvhcqRVx6JnMzDryfune1qoJKk6IXAbM7ldRiGoowe5BkG6j76nQTciyjf/+9y
5vCKiVz9qsnbmRWaFcNP0QaJ/iJC3jyRyub43+isE5cu7cE2KPFYTRnNHqqtAypY
umfJTJKRu1nuGM+dNb/gKR7KYbClNW2ph0SYYbJStaPm2ylqNv9NpxXW51bcKvue
GJxpV0pFzzU17ygp3PTP+u93PA3++Q3AqnhZ65gdsx07WgYzDGTY8GL5dIjBdpy9
CinaKwAm4lmVanHj3jFCIK5Kzc+cURGFkvaw6a2z2+PD6zWn0RTrBahSykt5O6Xi
ucdAWJ5wmeztM3Kmvtr/9tm2wWsrhELyaFzOc0MuUOPYtzJW33set2K9rasl4Fj2
AxlVgajDF8FJaXmAnEYhPbhEJoXaOIdS0Kk8iVuaKgKv8+PxF+kj0QnMm6vd0373
mqEXXGOYxhohrduKsyeLS1w/PF3zmIDsQOtUVURuyybXteh5h48wPmH8Yp19eYUS
UJED9WlZWVSMR0i70EeqvfPM/Vyd3rdTUOSiR0f4IBh4+/dPRlKI1BuQpooX3T3j
vULN76gtj910vILHERSRLARcF0lq8c4vmvEf3dQdbOXfGVpTRjhzJQckX5p3mjkN
ifPRUAPn8ILKSg6kiomA+nhoW82yeDgVg9XtQ9PAOR7aJuS6Im3szRvO8gydHIYP
Ime+APKrBUi7SaL7/HokMzoSvY9KxyTd3V84vhnLZpUNPkOUsO5IScWFFXyRFNJN
L8C3iqwxboKAKGAkCr2rxk5CTBCJG4EvCZn5jn+Tc4ZYtS98wasMfnuU+LpzaWDi
G0g/fNTgofHOiPii3+u7rr/+H1YYN9SBOEU0XTsBxe9fPspfpJXENFRBMvsP1vGZ
xp5KOpRXTpeK/F2738uw3Yr5m1PoawoWkapwFgC6DSzIVIJPyEjidhbGtdhiC7XB
VlyVvi8aGLRtB5L0A3omUMgozOpUxO98nUMvisR40LoHqMFPZ+gUNcS4maj8aejf
ACT95uegBu0TqaWJ8W78/wn5I9tFaEe56ksVdNztWtuZCHtlKAm3wGyp7HbIV253
kQUc/0BsLbAE+O5OcYD7QZBQAdjGVdLcIqG0KkOQ1eebUTmo8dKQHat25UrPa9Pv
Fpte/alrIo3Z55mIAJLnqq/GMdfC4Lq9vN+6new3EFUGgs75Z+Uix+HVmNQHcKA7
gjaS4itqrNUAOL/eWUtbku7Z+T+jmc1vqPhSpfkDe6qgVdd5AGm/89fj5PZVp/C7
DZa5JPbWQBtv1FNiFjXz2srwDmHM6+noJcO9ccQmjOJFFkm4buLaPnKoYjhwzq2q
FB2AO9xz5hiw6T8YqK1tzULH+KEQ3D3RvqsgdrL+ilwGZUdd6TzWEBeB0UAfb8T6
mpCdluI3YTCKxrJgnTtGyKEkUStzSZAv/lvhmxhYgmgbWH96Ms6l5FWMemehGlb/
jaq8CWEjKWMl7OXhd7U0hnQ6WvXTb/i28RNkqKTjGDAFOrvyX3dmc4du7HSbTrvR
xCrEqfQLg4RzGuTngKX8W4m9z4cjA6rK4pSwL2Zp8qU3bELGSaxJTxW9r4gjbJZi
u6Tby0XM3Y4fLeqdWDxrlyDL260iVhpnOonOKR11aFN2ovJEwJlZKciQHwlNykEU
o8latFHxjMvzx9Dv7X3tVvUSDXYBjnCW6r94VEJM2Im1OTVZPa9Jnvqk/qH5+xzm
10EsgDB3i6NqSYgMfJcr5raIwQ5KgC/lO+XfownstT0ZNH7zKooCl1Ca5HstPt5u
JajjuEwmOg37dvpu/8o/bOxfmmZBJVSqDVQjZMtqGXkaztu51EKgD/LFY0fFz+Bf
Rd79Gw/ItilTpvNhprbl2cKo29wjiLlSHolSPNfyf3gpNtuCXUMAJZ5xnN25OSEV
1FWFlLSSSKgUYRHSC0R4ChK1uvIj5GI0Uvdtugh1iKfAZBGVhg44sAYdEfRcqeO/
XepI8jg5uBKq/IiT3B9Er5SWTm04Wvac362htZpMM4dC0Xads3Y+DICm1abAMjiv
y+rZsSFvr87tkGiQoGbJf61aIHF6itZuVsu1i5Hwdw7w/4djOTvgXgdu4zya9m8G
SW6MsxLUqP/ydNBvhbO2yhaGKUlFzqSGjVkIK6ftXq6Sn5MT4b5TnKGIClCLBDXI
C4TyagB1LqpRdAg4gE6WcUiagW3nDOhUoUs3nZ3cWif9grYMuMXWrDSa11CsKBqY
1TLLvVrp8+WsW8EYq48nPOHp+4+Qbk6FLKwGTpVFanJU7HJC97m0W/7Sxq2EUC10
TDmcOhM2EbaZeIASmrc6vBmosdwzjSpLZ++jI0/bmjFnGrcWPgd/C3KPp/WNFsSC
wTg5JIRJO0uNtTvsdfoJvxy8T4IL6SpY7wbPKuAR9dpr2/Ivj2VlL095Ec9rOdk4
W4SxDXL44RtRGnl7z6dTcY1L+aCW6Jpx3aoNm2JBsia/1USOXS16WXf0t72XO2nL
raTm5o6Yoz4f2QjWO1wOqI7lf1q0r7VfBSFv4RiagWucjL5sHqIPb1pVassQJU50
81C8x2U/mFD76aMFAoNnVjsa4jaBHRXD4K3pePWT6No2rXETkU2admCGKOQG/Y5m
Z4riqf/2FIWGBY4xOvG6yH+2owi0AIa3u74D5rhe4sQgniE5E7Lz7nq2FW+2HR5G
T8FXFVC4UitivcbFOkMUqUcdW/acRRxOu6og/WhgqZc=
`pragma protect end_protected
