// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:05:30 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
pl6tu2ZVDwmRAWykPokW4tozzUiQTuteWf2wUtbXalpmFLkX8yvFXpHRReyLmuZP
6dZX2Qyrg44aOVwotWcTTfnU9mvXdXdsdhpKzgezL7gYPvM3yggi6zJtn/jqBeFB
kmXwdfa62q+dauoJY2D0FuW1wA3Vtu7F/Xj2b2ha+ic=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5792)
IU+3BBKYhb1ILMNFF9CvscwjqLqg5s2iQDPbUhoSP2stSEPA4hUT4prL2nh3TbIB
rK73BRWcuJJKrByJTFnFVyfNflk59caqvIGnGUXMjeBq+xyZ629YmgLy2ChxrXFf
qZGl6V+ftz2eccugd/Nmk7cKWT/y3Z4EPkqJ+ch9rQC+lrCa3225ifMv6aWARbXF
Ve3krXOJvGHOV4eCwU8LYOhMKbEATOkxQVP/sHmsnsYkBypFXPqyRLw8Erymcx8E
ij5MbJS9h1UxUBUhfmMPoMUSrpUALFzf0fw04iMBPMglHM1LuDI26JoD5NAnRAnZ
gfXO9liJn93+v3WcW/vAnsVJEzI7dpnfqVsMnV1Z7UBpDBHKnFmRFyy21svVkdEe
jKUHXPLJqyLyjzlrs8o2bztwYgWxHXSp877ypyhdJX+29Hn0MoSL23CMYiz5J9/F
jfQ8w94kajbW8uPEwzscbnJT/LV7BC8aEQ7dKlb1ACeSYtWlLUiu7xY4njFEdr00
9nEhwEBhBc5bFUazpynGrisG8c2qtminwtKc2ObOpoBtiez+GUSMTxv1W+hctdNM
+1p/637y4tSOUF6GKDfbB8rNOKU64dF03xGEqN+exEAT2EICJNfg2ycVxMv2ab5v
0K27AHNW8xfS1OO9qkDV8i34W5ob4Ow144bGrpOu5BsXou3AemD8t3g91goEdbm6
meCt94HXRvhxHBBach7cLMfqnUOuCCtGfJgXa5jeKdLO1Pmve7iY1YISBNXnjsFd
b/k4J9E4o6LJE9st5T28cYmF/V73UX5n/ebFBOJz4Owap4iGl0btxOUGpt1ewJaB
CkuYEgy0hgcfJm2GPi2yLRN+DCEz191oe9e+kVU2aAGCWZ0VTCgAhvr7IYmUDR1h
lGQmpCcqEnhskqzXmfRxfXTi9xh3854r7fXfL5vwICpvMHi4r8E2uimkKnEmrrQQ
chyPyQ5dfpLUrVK5sqQDnK6EszGHTfSyIjG6OdzdRzueh/1X9QqOEZfsRLnldlis
QOafEtX50mX3bVgIIENJJJNWMh8gda9wmLGbLLjvw1Lxf7xD5WfPZkqRrt4lq3/w
ev4f9PGHb6u9f5R/J0NILtdMSBkC90a+phfkyKHdIk/xje7psK19lvUm7PPtYaoW
mslyEvsr0h10c3QBnj2UsufrE8AcZis3r/A3XqyIMGhRkE6Z5Qdpl1hFIW3MxyMm
Xjw2bUWwNeG3mADL4MZwkNHer2+keEG6r8ACCjxk5/r7Oj2C4hQThOUysYm5G74Q
gXhhr0c9fspzSgvZvwWhUgcLCNERYacry9KO+FeOk+zbAIzDD+/3ROiATObzKniW
XVKhHviJ/uWOztpE+7/V0ocFd7WtT56SwjQZWZMBovEYCN6VNM3dEJuIlGi0Int2
TyuUaYQxrgv2CzbOdSlbAn1rXA1XczBJ735hTiCvXVW3IGDKGDNqkKt5Hgsvue2k
kp4AAf+f/KwdLZ4xhOXfsxi8Dero6cWb8uVXfowVp52qv9YJgmnjQEvx7HeyiI2B
5TN2Y3WVALDlrCfG6n4mUyM48kJ7eL8HVokI/hY9GE0dvKlm5Dy4DZQECj+W4f57
doVxmLGoOm+Zo2a4lh91Q6gJ3tcUNhMyY7xYz5n5PIUoMEz7c+/Cb7peAGOlbnSk
6CaZHTOB+kKlfXVeiaRHOlfwR8OWnQ0D8w3kxJZALakmimdpvrhAKoGqChwwnCXn
VXI9sgr7ne0prIdK/CKqNbQGn4DFOmkcIaMsXHk3FjFP7NgbxAnBvy6Gg+xFhWEH
UL+8EOEI1sxni7jMyBWz/gWn/XiZbt5rWzpI32Yko19GgSWpiBYlUarIbaUD+n0M
4OSFN6awPwX/Z+bZmTu2mSHp7bF2LyvliFtBo7L1GZARd41Uq8le6N0HtbVfFuiJ
AyG610MynVvP1mEGoFgixtWvdtUgPYedCW1vC5/Z/OerhYomIiNGeKMWIKwPTgRS
jf83yx2IOkpJrfhpVa6GLDtGt0nHQjqll9kXj8Rllal4YvQHx2f9GJHJBhEaiSDa
IsFwIpsYhbLHFrzB8U+y6j7RGzVbjZSpJ1Wp6H0ogNw2ai+kCyK5ZWas5Mx+qPNN
GJmDPCn2Np+GtGrcxCWdBxBK6SSAwtIcmvVlcbp16qUBI3bu1c9EnBkXyLdRS0xu
g2KlOjA27NaAPuhkWx+GOH5m7W/MHMd1UVK/2/8JF7oEmn3eaniEL/S9II45OauF
3k+cEURp9gvXSK/OjVU1TFssTnB6+FYCpRQ4YAXHB6mD4fGsq0P9K55CJdGCzb1w
5Kysz8aKfiI3hpx5WxTPdKO/ZgNR26JMlneaGJlmBbENX9+QgdVQ6Idfmd7cchQs
4VRpYloOfryL5pspHmflaBb57USnVmdJgETSLFKbjW8NnZgv7T69t2S870FIp69n
C5A8c4memZ5cjLpzMk4toP+7A5MlrC2HCrqTJetv06mLhRfcs6JSgG3XdNElgfmG
brUy93J2/KIqK2K+NkXNqySwpbxgehrtUbUbwQXXiHumRQ6/ibh2hGRquzZ6Hneu
kfDPwQKQayQFE5f5N8X+pSesXrKcmlBxldNoD1BZlNhEhJRiWb5J5GY1anwIQFbc
2HyIhW3q1Rm8ObdAnZipAUZKVnSv7kMNoNk/wQ7+M5h0ta9Dp6AoJPUBJuLNDe9c
0FfpvC2SeVSzE+d7VwgAf8KkNyj+oMbF0fyetfepAhd9tb2PPoJXN5hoR9r+CfaE
UWJZjZr0gErySBzkipcDmF5usH2cBCEUkaENv3o5QnmSxj6wzRkaVrlS0DlPdvG8
hh5lS7TcD0FdCYpWc2OzRQbKqkdZSJeffnuJmGicJoj1PDntv2UAkjmMbp2tbOBv
8Ch9OF/1FO9zxBjyk7yQt3hyT1oMqLTC2u1jz9W8YxMfIpn6AbhJ3Cf7Mi2bK5El
pDVLW100pVIaA659FfO1E8fuU/DRcp/U+SEQg5tstytBWBTJ32a/2uJCoPREy7vK
ag314HgFcY8YaZiUvA3u8y9rvOvkSn3nac5jgmTEQsZP64YzoymknSYreJRy7g4N
ZleBXvFmTsICqHhEcd0Gvwh7N++J4D1SpR1xVbH4vH2G2n6PuqG4PES08vRpN/D2
uJT8JoLYTjEEEmwIiEtd7x4Wa824Iwb2SJFWGAIHj3wljBM7W7geChVEdejxK8Hr
P3wXOHfw59oKUuusA5XQg95u/jj7z63Jtc5ZeL6ultP3pOo1+XZizMX+QxSLDZ8y
LEG/YfKggJAmYJb7sYnssQkhVAxJCe6AvnOKNp78gzrfnTUYwGuOrob80IAhG685
8grN+yYZvysAaZyWmr5tJGAskEDipfHrnHE6nkwsiNI50ihslI6sT6HsOfYPVWmT
6Vu4JsEcUvOnwqQ6SVn2iITRBZRaJiIiUw5E1blxsmuk+OTiXdxfZqIubFxteyOw
D7Z2RW/NBwS21LyjK6bFqgiBJr/y8NnP9A/ZlJAy6ikIn8oKeWRw6/MqK97aPXxJ
KprlqHkC3ssxQtE5hfjWnII/+1Tl518TI7lTwdBU2Fkjxdzaoc00c24YagI5PjH7
2/WPmGkpenGPYsrKlQ6sSCqMDt+GxjvM7ATqNcu4QngKZRdkDMdXGWaPc0Vldzyw
aiH6neE+iG0zka6kzkYdzFv/jHtAVyAop66DbZIAAfJMnWmEmc8Uu3gsIYGcHrnp
gE97QwU7hJAd4JjzU3YZ8ZsDoPU/qdKLsBmv8s0BXsWa4iqbs0ixf2PDNvR2QAhq
hnFqHg89iXDpQPLbGqrf0i73CthtDpHoNFrdvBGq/wHfbAra6b9t9m7FQfM5ewD6
Nq7pcPOclpaIEG3pZTAi+4eL+dJn1J2EsA/Oy99lkJDHUW/XWuUSBCLcIGcb5q1t
6Qi/krewn2obXufgX8YnESVlFXNk1B9+OwpvaX/EBvXPQY7wKzvgoaK6C2Ytd67n
OPFk04HOHMtjV+S1dJTOx/4G9vfrLtJt8RBdp6BYl5Zs4EYsIxF3pAe4E5I7qN9i
Bp51U/jxh03IEsajZOCLPjXI3dPDbHr0bU5hbZhi92zhNtWAapHiB8BMDK4D0YkB
iL9McdGTi7230D/nHzYVPKgrQ233lRGW1plwYBxEQDg5FrFK8c9toYKWmJKMwsR2
DQevLlnVFo0CXpc8RP9AZoKCVPzgt2BKlulAUX0yrMqGFH/3/fJpm5AFaVoyYB0J
KlbmZn7SGUtV1mC0mx0WwN3S8GlJ2svbsr/9r5JvkBLAOWRoGHiT21Pu+xzoP7U1
mWFY86Gf4XKtB90MBDuNHnCFus42HWDesXCveEhOLmBVHsQiaCRIKaAdcU9o7j9D
YmXrRQ8twQSkYBheCjVkRJT4ZUfQ5/MEuTQGeQh3EO8K8P5nktXfhQYQR7rySRLq
Swi3Sd1+jXfXUlM/kWLKU96awuT0GodQv+P4/qDZ85LLMdfsmNlkBaPR06w/B0ZH
3tnmsliVS1rFiwwzvuErGOo3WPxwMk1yjdsmD/BHVTdT4CvbgTueIH72EGPkWGxE
4W41fX/EDbgy60DJPxs+1eezCWSUtJlleejfqlCoL8vEIpp/aIYnuP4iOmGvtwaD
GsN6iJawmTaFLja/pYGsVsECb/wbWTJxRJgfLRvYquA1OEcPr/KPE1mrXwcBhZ1D
QQpgjbWNWXpUeQgjKwsPVcpArqkYm7uBtdX9kvdoWkxgkPVhRfB7LstOmH6MoNWp
WC+THjFATxokzIIxI4hv/0G5VEsxYGIFlXOj/duxmppde5bDJAoVhSWDRw+KW2N4
ZNsVjRYI8CucNLdhIFVlMKDiLAXhacmvVActuHMiEwV6iDXp8/BzSQUviRaeYN6Z
9uBCic4PvqQ8ZnVbFoEX9EtyKNgWmMaMI+i1EIUH9i9kmiTYctxvYJWEiSfrttNL
TUABiDHOT5iqDX71J9XUBhXUrf8inJQRKBKPP8ZSuFGSfrtxrmnOM/T/O852Ck7S
FnE5M8CKBQAUStIOtHnqIA5jFlASZRb6X5x5n33U8oOBaoUmBvqdGyKcxiwKyY5s
TP/BO3gjJ5hHyKYSYG8Ix/Xk8hlxlT5N1MeAIR5Gnpwm6LjFwdVQ5scsP0fK1/2A
alDIWq9969qJ20L5OOtmdhi4NRw3dxwWEaKQWeazsf3RN7fr1D2FqBZhBCkYUPrT
YD054wS6SiB365fnuc1Ew9765IYNaTNcrVLua+RVwWFzIDjG+1k3ieGo9GnAWJ8Z
aQn//UFU6iqW/5MkBDSGwhC1M005RHPUaVu5pHAjDrUdKcfW0G3ahY9H/ZfGF6p7
Gn4xQMXV584B++G/EShDnENHYYQBEYZdmNamsLqlkUvtJBxMVWKpbCeq3zDHHueP
Aw05Qjn9aNxdQJxEBsVOybGZCglAN+nFGCf6J+MSUqoOSrvktYIiZdUL/wRXFYBd
b8ME3BFL3WxPGCEuVfMr3Pgd103fGvScxU7EV6iR3ty2RbBc2Zqm/1B1nfi2UliZ
PIASf+v+WsaKGUYUeRYZCgq5ZyWSmHn3VpproensFDMSL7TQLpBi5A2yCcbtgxjK
tpDLLOoUZ8FequOilpz7ZKnkAaW/6ccaZy5hdcSKboEgOCyrd1rTE8enDIIAJBT0
x72eEdmcc6WOzEE8QzxIfDBXgVtgYn3PlaP5PziwzAlHOFK4WWHQLBSrqJXe0tFn
jeCFax75dD4oLN5cm9B7BLOKJwl9wcLM24d6iPfkcXQe+moA14RTpWDhfu0VmUkC
VqPluAg21NnHFGDZv3F2lhT2YrZiSZVBSdbflx8HleQRQyVODcpIFoXgu3IAKoVh
op4m/b5CA1TxeNxyASNXs22Dv3bnxj4Z5bevgsb3va2DvT08080HEo9patlHarUU
NmOenUEXOtjVxejHB08bcEbn9ZYvwVcnJnmPRknWvHroUQrxz2PNhxFPc6Bq+qWJ
KbHwKb0COHUcOlaS9kZ5lEzSf3ahDASzBdKYE0zODm5PpV4BRoDkCcHpfq5kJgEl
sTnjSR02ZTYWt56iW0Yl13Px2XjNMURnKM2UJS6yfZExg9k+zP6RMlT+ISuiYm1m
nLMpNDxUE5o608A4pRTTP8BzoJNSWp6lWxH5+fQoqTm8YeY2tzZ3EdWSCIn08pIJ
rbrz8hm5p/XT32uiYJHW/wqzxR8/u8/tWPxvBHMMAc3s+FdOdIgbirTq6JpzAncR
jB/W/7S7xkNLZWGhyrCum2RPLde53TTU/Ku7JYPuNxZ5eINnhwnGUH/dg8UOZcl0
5HWMo7iVU9pDjkOyGthK/Q05z+j23+4DxXB96C/CvFUgVg9bp00dqPCMmG5a2dxY
fUb9AYKchfdYExST/3VFdY5qMPL9WT8dS7CboLnRWTFkyOfdWlYJzJfO/CF0YTFq
14RzugI4ATh7ALQIzPfjjT6szsrbaBIW+u44kGxR0b9xShhp+pXT4Ke2tltl3TVR
K5Te0fQkwgrp05/xdlj6NaSJdtCxiKAZqCkPpGtqyzMOSqe1nq5VQUWdJjOZAUST
TApbpu7WIVJxyOGkYaHcWZx7UkH+Ql5+jRjQEq53kMBNbMbDT7lVSFLvqNb/D0J/
LmBL5qMkg1QZYyg49eEpZfrwqzUC8Yl+GbVx0JWf55M+QYvddDW3rSkA4lfZeXe/
MMuDNixVHvY8qg4sv93LmTol3kQxrf3qLRRlHblQaoqRa4xlwo5aLn3fcUH6tIIk
YoxYnH6Y2guSo1tNr5Bn3+243I6HB3j82QC3OomdIadzZJPDPPXRoXIbcwz4Xkwm
U4ZSbkLI75MiWzZ/IrdBAvvoCn+eMGj7BuhbHGGuoL192NZO96latjNmA1rH2L3X
cLHGIxPu9okKTwyn9WNUHFB4Wx1LSiAq4MlyZLqeXfIhbAUGa8oA/lu1/j1zsj8l
OkPvnWonfQCVK4YxvKEXcqiTdyYNnOlzNPHbmxxX8g3vNOqmQKqoO9hKc1Umd+dK
Y3+hMLwx85CLZwSRxN736UeaHMWYX93ern0IYI8uM+oALw6fK9fWtzR46vsDjCKy
KXAzzkmaFnI7a+qR+m0z/HbDIrd41cIGBUC8/zZXOaTt9236NiPQH47Ow9w88MMZ
vKk4NAtpaXj41WV98boKH+b7LrHKrCzH/eFyHiq6hoi9JqCihH9cr6OQICN9TC41
3BDTZWqHRIXqZo5AvGDyJS77Ty9LFmAlcrCcIYJMp6GUIoTTO7QPoyF7f0NMLlAV
iKhAubv06/eFacxJjJsH8f0fZe6rTeYOgJKAaSIAFX04XLMb5QQlNfzqpoUEXfwC
Akmt5p6e6pJrlg94Esf2RwzDq3hIbrbijRDd0w+Ds03kGGWbfZCzU/mUOtQwMTs/
q3hIWx9vHZiSP/yFwCM969hEXgjffRtU0vc7DnN3OIkqmIA90BDmgzz4TfNB4Uiz
c7KMwlpDa+1D5zCnzQv36j7WQr0ZwRGY98+Z624P8EUjE1fK1V3pZhLBHzUaADrW
Er4W3Yj1LoMksTk2bcKgTtqw2DusJIw2CGQU6lB9QCjJQO6ueNkmocoDuY7S3Y+N
ZVfCV39H5RO3DLPeVYHbIGoOx3HagEl6r9hBTYv/A7Fhn7URZCteLLO+8mhARZiP
SbqIa3B166UK9UGXtSNLIg9qQR715HhWigFm+irXwObFA1ik6aTlGAmzIgyjuLLh
2m8hf4kG52STW0ibVUqN20tAE2bWGeTjn5+Y2xrfH/w=
`pragma protect end_protected
