// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:05:37 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Ln0BmBPXo/1p/CMs1AOOAi24t9i46Ff//j6RNnLUb+hqid/Z3UmTe0sp2k3MPBhA
Gq9L4bWN/YHRz08tkofq/lZGF/hhOHkQ7FhJXq05qO0Ly0KW0/me3FOiwguIZ7Yd
Nu6VvFq96w7Gvmzns0tmrR2TwJZ9zpBohAYWsR30R2E=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5728)
Umykilq1c2eKHVd2GdnjHGPKySZ8x+BLjcqFA+FIiODllTC1vv1HuiCYdAY0V6eS
3wXlwKaQt3Uk1amBc+r4vt7LI+/1wIXlLtQyPGibPSt+utUoUIqpGIUBWTc/+nib
HyA983eFjzp19ELhDdgM/j1QDb1nenp9a7krdnE4EljqSccDjZxjFToesSPA2cll
y4W6NvrCChEzSJ0yryigwIk++l2o+dSu7f8tyF6mVCCG/MqT1CQtoWz6JQqhmBlq
580KjpOUxo+zMMWhpb2AU0rmHC9PTEeqbp482mGP9zOAq1qmjcjREzrEwAhrcZC/
pmXYL1pmT0GJOdGlO+D1SeS7bnvSxPdIhmU3zLvDlwPWUw8zsiMslK9chxJTRRzd
+WXuHqpGI3Q1tLx1uVZ2+N1r9yARjS/BhBRPafhZcRemiG2eZICsZ8oD6NXWaisC
0e92zbPWdLMcBvj/wsxMSSdC6s+IHXUVB+jddA5AxIh3T/YNBgdc1rBh4FIb21g2
UgPSL3YKS0qSNTHE1dW627bF24hxR6ueeBoS3wCu4hGlWXZu9zCma6MvAp3ZJd8p
i/u8XjTQvpXMou/WIrMwwKcwl5xa6qaD06/UhZ2PCb1+GEVR5Ca/oPoCK76UCKTb
39M1gG7nJi7cwjYxhPy683HLzd9Oe+29SqgmXck+lugudoJySmOu2ELX44qX4bkX
srJFtbO4gd7BBrNy4sofG6KchQtnux96G7fdffU7WzRfN1+oj/juoMR0/+HGRpgn
/vAUTMl8ZqPtfrn3qyOZj6CLsXquedpJUtpraE5GH2wFrojcg0buAJPqdzuKXeb8
i+w4KKiOEFO2h7dDMyVIHFMF6J6IkQGjA73MYsLs5T+ivj+WoRTu+OmQuc0qsIrb
IpxEMb5r2JlmjKsVLt+9IV5qNZAcL1iQv1/Dpdf5YrTS1zmJVYbv3sIlHg9KSPKC
XwO6VpIeUXZz+FeqVqnhaj1tw15QBlDtYIJhgwCEemgTwLZ3LXC1LaT69/2hvT0T
QclzR5XQYfhgFDF2UeOND7nTdIVqKx1JgQqmDxkZBu5QF/PlrRbD8c6s9fIwrfrC
upoafRb51EA1HETYwSPMW/DUzUMQM38U10Z2gqk6qVNcdeArDz7+0rQGWWQCpQWJ
BgP1VoIVRrT+gFC8xnRNsaHUdgFTFvRatlHMrmaab0PA7ipnZVh5IXjTrpsLDCC6
CMZK3yPKZR0eE9Ijaxw0PY1HUkBBRLlEcx29p3vNKvQIAjRGrRkLU5hteTdol8lE
DK1PwXCO/CTTZRE0FaWVgYsCaVy8fX16/+3o3CPSsD6QMXN/HShUqVtPdreZXIZ2
wwOG3XsgfFEM0LCx5tci/nPcpgTk/6MKvFvb1wUHWcAPffyB985jsBxfJiTr0EJu
9kwSOBYiXoWk7E9T70uYLcuZCGpdBs/XD84NpY1oiP35LqfKFjGj8CrkxYNZVG3U
l77rpw4FKlMUPjMw3evlRTiUalgYoTdv3G0Fna9Ue1Ktp2bobyHRKH/hegfWAxKm
3bgcdklN9ng5parYUc1rr+g+4Z3jenb+eWTyKBfkOWXyHESDGJBh3bZwMUX2i8zP
mAdol6NkxOvy4haa16SpTuXwqJhfJHbRXZ5s3fcCrrSRarTLrWRP129i/cjrYI5T
CYt3HoimakPYBXmg5WBfujAcAoHSdJBR2Sxj3IvtOLXkTlekS8hUc041KtjI0nWw
/iZs1XAy/vC7iTYPQW1zH1jslLRd6QnSUm67iqXniN0acdSUE99KW6kYCFiyUTK6
IIxHMJ4C3QXvrTUzxu172lVVx5vqPqOr3as4ko2q/uB0emYrSwy4S70LxiZxh9Md
w8Ati8eeAkbf3ZaBZf2ftzfAwItZUZ+uIhtPs11Az1evODV5sn67f88ovfE9g7mz
bP9pkoeO8rjBv6AAqfWLBP05SAEPV6Qh6F5yvgI6TLvygN7kc7dBW4J3PuE0jUBx
CGP67wSqX1fUZTG/dGCxzRF76uQx4okXjD1nBnUV+pcODkQGnlvk1F00mCqOxbSu
hq7/utBdoTPFt2PHMwfLTF19kO5HBALcEg7QXnLGWQLyPj/T333ZnCc3kMmB7hZ0
22hsgyzvgXvFNWuVliFiMpn1GO/c8TsFYNahEAz0X9bSJTz2DzAElgdORGTfJxUu
CsPrf7/A3OrmXkJjfRgC617CJySKrAUfaZEqBJd8AxReHkoai4Hn/vn/obAscZlZ
5s/UIFyjeQr4gv4QZkmc5geZYZ4u7FVFgFnBlZr1b6bnIwHNLOIclvPL6ervrHgt
QW8K6rsoSPkvI2aSR7Bks9pkaSEt+m0nJupN4/uUQjEguPB00+Ag9HnTiVuI5IMn
Ld4aP4U9kfMK/DWUTckvd2KYgW6waIDhuo3SLDznF8w6Tnh4DSyD89jKMXb692JM
ulsaFndvVOZK7Pm6KJiwrgCycobi/8rpObBTmVlaASDrzfz1MPp1b7DywEQrOMGd
Ui8whSEPDtzYOrgbZ2Xot/chWNJiu+yrSF0JJX9+SXNWVyR1vS9FaUeBeYsSc0Ed
9jrYh1Wlh63YByuxmSNlK0W6nob4JcCVF3CKwjL3BrrbIywucOInVVywFj8F3z8c
QdbYBssu7LRbeC/zIOG9kJlAjo2gTrnr1xYEFWMMNKjMSfVBgcnHKCQGWPDujC5u
G0fuGcpcgSMLrSQqVCnAJToGvV6eXWeK5o49+UYsKfMoRG/3Obx1N1L5VEVg9v9m
SyGfh3BBS/pkn6Jky/4smxY8+oLtedXxMgaIOk+w33N+IsEJ89tpxA7VTEIx5uIj
JHFMKAos/TaksKcYAluV4gq6f8bBSIPBtZV0sk4aVt83UfwRwDwLPaxRlvhw7uIu
c0PXcgrixy99fwzmoAxSEzoU7bqxme3k5IHjZbjyEI1sg0hZtMMue9fuXX/nk3yq
0Wk1gZgkon+PyoFsjQ6CuOrOvrvalyGwpBEMwNL9XZIdN3cAovaq2HcYojyz0I7l
lQgTZi57oqFqWnCW7KJlBA7hJHpKC5UtSO8zwZKWCjrwaw3khpQMMN8tnxg8+fjo
0uy0noVGv1t7gIvQ68ZxqRTrm6STXM99eo5UhBfMd5FG8Msni+OaChraiOHRu6Yc
qI6dJk2qzuR4hIDBpYmKbBw6bKCinbrLK5/XUHQsEHEM0XonYA+xboSxsvoLxCUt
2GNLrocus6iJ0V5LQjmxJKPfL0eA+I8cfrEAlmPjYo1GxWZOe0kPNHRpIQC5MZG2
cWihGsZZWHHzTYdlIUUegCwluvA4joj1Y4f24f38WabNpsTyOJkPOKRhEErlP0z4
dMGqHwqO29KAX0L2K+KGHq0uzuGc9TtayShtPQvsehRI0FYY7jhMu/Y7uwXqwBnN
6W5ehu9i/HvfLnR5ieG6/7r0g4HVfRsh++h3aqz/a84QPeEE49Vtd65SKXGwlgTI
Oql826Dc8PHOe6mLTNs/Fg8KevlTioUhYCz9iphYP3N+NUETRwePhhp+d8jC8NpL
4DVeK1x466RtLjV55ekVSE4jFi8pQ9lqiztVLZ2VykEZ9G4VN+etgXoPiEl71dj7
mIdpV8dMLx7+TnREylclUUNU2yRemEWu2n9vUbFLI49cu+WVoyNtjh81Mdb03kfd
P26H7bul4SWwZi9IsamlMI3U0fPKJkssz8vOnATibme/knxplIzNFsu2GP4sYPJA
CgULvKBpykuHPEUiG6VHNl7P1cVIYK8lKLhGEhaSmtuSJsjTlpstW50VXPbVgUEs
mbM1ySS019gzZo6hgtLLullHPDtRl4Q6DGvlgRLXUVpIVJj915ErO7vtGxR6pjMa
VeF6CbgaKxy2sykRELCPLtzDMrDUJwCudpl5ZNzLvFVEbFKyUOdOTUrdDpgISVI8
W/KAH0OtXOtPqyoJm7Tnk1Vlt2zX9B1OdtRAfbJo6N+pN1Nb/4XgNcPEYRUPIS1y
rVI2POMTGQnNDt4VFcsZ0CF8no7dIignuA6EQ7DHaDSueMlNCIfVhQXQhyEZ+htJ
YbZsVmN97eIvf8/MW48A0Z70lvcpdSQbQKps0YAyfOpGnduqHTsX0agkAkr9foUj
4hV8KZaii+O5F5kNQfSGnmPNr7ieV2LRbKLjmLtG+eErvPhQXVMpZ0ofbBllM32T
tF6pcE7aBoVbumicxImmdCuhFiHYNcSxxx1wl3R4HeOHCWLUDLiiGRtijFblNi65
Il7ZaMTysl8DxCrjbIQybHnRP+o/thrHIZOh9M1hkVHBv+LHnKBSeAX6h67OQymU
ahDMcALwMceumKIXx76hnknn8OA2EeMLYPE0NrfT/4m8e+qgfULrU0ALE0kUIk2l
HWRR44Wdbj3YIV3bJ45LmXOk/M+VPo+UsT0SdgkdLiSjVuQINk2U6h1PZSqfMj6o
D763bXRU5cVbdds+U5pZRoGRxCd2egJOjP8box2MH3GIL/KQBxUAIHNZsO/u9kMO
F/77/0yYhT2cf8etrpvP5fp7rUki0DI37lv24bx7gDYTryTbXlI4DYQU5muZQKhn
BQtW6UGT8nUiJJkc4FCuE1GIDZH6Gxsr+kNQA/M0pMwHT0OoS5sVEoBKyQBW3YmX
Q3lhSiEkqkbx5mAFefIA8kT8D0IOp83M2acs+c4u5p49yKx3M3vmexmg3YYPRfGc
cfmDYJwagiBVhkRiOiTMKzsWVQ8ED+ur+If9miEAzOFkBwrgEzbhD7g6XDOqdT+i
8tBHjSTaiG2jgeCr2PHDDovH5w6026gOrikd52jD72RGc8V/tt3qSwZV8b08TqHR
EpZmXCuz5cYl/rPRPSeu/q8pepvdjZoxB0A4DqhWimZbAsuOy2Nnivz+feXW6WgI
2XkeHrF9xLGNcfODSKlf+LBM4m6cAQTjyfsi4aD3m5RvtovHGjuepGJW5EH8H+36
HkKVY7+rk36XroXZ/o7XHpLcvGBz8oBvT5j+tNpUoQ8Fg5baAEu436wsBb5I0kiB
wVkXGGPm+KwDEA0r7lGOWT0nn7Mfx4tG/ktbxhCJ5CjIsANmdiPWQpdPteRb1VYZ
Tajeu4+qnztF1JNNLG1oE57qbTRQHkQlaCEnJlteaJe5673Jjo5pIGJJPA5b7I1N
ZDqu8YDEFxNDxVrVk/MFeQRQH0sJGMSVhQXBVG9dL+YzwgVSKBT65z4y2+dAdq5b
bpsAVWvsP+06s8eJ2ztR8oebyXTpyei9dc2b+8x1IShKn4xktuySFr7w3INlSidF
/Z6KtzkRwxWbHmzepd5PpR+8Q0WeszJJ8zotfaUTb66wJwFxT00CHlkCLHf6c1iw
Anj8m1oi3jQt83a/AOwhn1NbEu/zs+K/kO67PYF6P90VCpEw/Qp/IuIuFdvwqfu4
t/kRdGGR1MirhB1vvXZICRfUPk2flhWdOAgmeXAhlUnWat4wqJMloTz99tIU9ekO
bCSxRXjPHcWJ84Hsc/GMRfKuQGjeP/I9ESeq3ZHg2FQml9tMjYsFzG7JO+s6RKkd
7d4nHArSdPEaNNo0qXh9iKk+U0g/v8m9VQEYB7vCtvhaeL9Vi9lmvENXLRS+hRUp
CgzD87W+lCNjm0rNSSBMqEExNF+vlG4mosn4uqhpii2Qmz70sdPNTWqYnk5AIsi3
PVBX7OCdg0T25VHhMAwSGlJyNtYdlmZWVhlQqnQNEUGYTEQfWC0Rwg2y59yxC7Hl
lEEn70RRPK8OksU8vNCbcWsi2Wfol9FMdQUlUK37WG1BLmWwzBhGzBF1sbK8wFy+
tM+7+lUPdEMJCQ/5+T42sMMspRQVI9hT9TMa4sxOXstk83Fw9eJZyKxJZv99qi9s
fzcmiUf8oc/II+mcZE7LbvZ+CkTM0DrXXGVOI7oW8j7lxXkSl3Zs7oXJtHhGq432
YgkSE+JENBrZTISwkxKffTWQCidQhGyqan8lFa0aHSPGqZO1F/ocSrpoz8RAalkK
oLlZQVyg3z4qYYIis0ZcaCuxchDgzfQtqqEJ17VcJKEQ227gdp9pqPCBCypA0S6q
6714wuaLHic4YuS9a3rmyfmp9eY2TYZklWgCc83HcL659zSh0Aw3ozfO0eLULqTg
RAMCFUIChPeHoiyhUQY46Ghy9Q3E2j0EKfTwZ2kMAMk5PwIEK0IyAWI0Z2rA5fkc
tM4rIfx0BEEVQhbaSiRFoM2lIOrJg2fm0J4B1OIHl8aoFwdjn/EztirXfi3HGcTI
4KC3AxJeCvfzS+tnGgFoY2uY2CZjutnEf/Z5WhHyL/y0WFktiCd+oYZJCLP3Xkg8
4okPEJ+g26+No7Ts2wuWrTLG0OD8aqyGfL0fcXuKzzI0L4zwhA//iq/nYEYqwUfB
4i6qpb1IHMsQCW9fU5W4TPrA9xS/dXccw2zukhUFKphEAhe7uzZse8b/WvYgzMsv
ASgC/kDdJAJHIJ46ilbahJ6Fx6EIhkvJhz6uWWaRlZeNhNa76UClzu4ZurnU1AKG
hPHrZIld60EfbcPq4aNZ2GrLwJR5h4MENlinG9dfntTzSfYWNVTf8NGNBCxy/T2S
tjLuY3TsJ6radnP6tx6oxMY3BbEoxfIKQ7l0kDfA9fxfX4wxQs94rKkpLRxkL7L/
Vcs0kiPXqxFyaH9gn3DNuQQURsOML6ajMftLaezkB1suMyVbGJFfJQwbXinUumbl
+s4MWCQKH211gPRJRTv6lQhFUmmoRS2VZe8t9WS6Sd5qTkv5jzR3wp0cH8Wm3+6M
AJdQNPQgDiDCKrDXRAQwz37Ft8cTCkHj1ZDEV3UqAUlHlpqt+CVkubk2enpZMB4z
8tWmE+7/5Y7H7DtIM4vbnjFzuYowauBPjMaj8etcQBhHotqD4vgPPW4nFspuTmo0
TKt0VGJ/Y+gAZEAkjiMq8th+gL1WVenYotMcTb9cT85l6ZW1JizwpM4e6Ru/hdrj
3W74sPOyJDc5S770rXTs8PiQlR08Q/LMtk7hVm2jFx/t7/Ihe1VXFvGAFZOGNHgA
369fCtHBSoDtFUp9GGEH4RT9mb0IikIrw527iH7Jvw+r5QHFtDFjYj/rokrgMM1N
8JpnMv3glW3SPEigjNEXAhUEySnASMXXKW13ZBvsljJjQ9aqVDr4gSmDVuCsIZts
aNhasnNC4vAdHdUQRDM5ungjOQSmrBfd+cVE0qGMQVKnt0Kbv4e5UaUVpRviGA8j
RQAAmN6Ke5HWmRcfL6oHJ4HCL7sJ+CxeFWilz0srqvvMAe3Zy7RMfg6Ge+mmUSPo
31tocb6ewtADtLW0LTUorzzFUUJFvZKOlYcKtUnQ76YJ1S6n0pH9Bh5tvpk0A6dK
hwPVCWQd1OcO4b6CWe0cT9CgyA8glJsY+6MUpDV66hMrWt6zQZNCcj+mJY1llVBS
WqgpE6u0GrerSE7fPNlsrOWMmvMNk1Smr4oA73bc3RP5Ks1NBRMvwgS/R1kfC6ob
aS5ZjDcEw9M9ckLEkWDVNbJt7jL3Ps326sFTqs/StYNYImC4KX69hY8uvYQ4/zbi
3ogiJcIxyTbRuzOpyuZxcw+663Euu551i86h7CnhxzdRO2fMDM1P41XClSFXlS0K
J3NWIf178xYThJH5xbNpokSKov0mOSg5MJXgkzzs6DITuerg1LkkEvMFzQMpbJ11
Q4rxeqgxetpyb4re5TFVOg==
`pragma protect end_protected
