// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:02:14 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
oluBlI8aT9uuf+YWqm192ybvtimydPGnfJ+Tpxu4s8JbL2azoo88swrQlN4d7UPE
fC8JCGGYy6X+0mbfj8zNU5rJB/e7xOcGe0cUubLQNkA74KOrUhQnVInnqD61ElAq
LmtLu+x32xBgbJuNYi3X2t4xKjt2yQz7dOWjO+/3Jj8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 135024)
KwOKSpvgQOUoGfLUCNYKB412zLG9KtKILW2V5DyO8//X81QEJbgY5p6JYVOAFBDx
9y0X5aoLuB4prv+pDqzlsY9yyPasucR0RKMdK9EYWGOBBY2BU8ZZozOXR/fQVgjD
YZ9HnUYzT9jUwefYHNkURiZjRCLLbKErHHdmWxQydsyvkj+wSq6OIamg2jE7KqLJ
sSVNRB1mcZb4nw8gUmHbsdQ+8+MylMTF1sRmifEPLXzQXpW7iJdV2YkqIvKfXlTG
BevqHCXxJaeo6asfQuDyQnA3LgBsT/zuipkIqu7pTFhjQ6wMb5yLHteoZPN+aILB
VyjqJOa9QKwcKU+BWLF6+OmjsFuOi5witUTPa6mK14QH+tfzCrYAaC+niTxbLLoU
FtKaUqwUZnUpUUonS6fb5at1i1z981SvydODQtqjLfGb70ZB69/RwJhl9m2veC/A
sfeMY9qiy2Y6ue5oP3J0S2dDcCkXG4BP/+zVFTC7DwVHP1S/CZKKHPjpZi8OiQ6v
rbXiMbplqdOk5QC515pgmPYJaLaSB+Q3TYvNDfvWW6/CquEUPnXCPNPEY38MKh5J
0WPhUAnQetJOFv5c9Zh4zmQOe3SgHTiB2QyBTD8gYZnZDGotU1MSGYgqrC8tOUU+
Keiwg1eGcoSTSnsV0e6QdbZmnMQ73FOs/Tkub+gdqXRdY7dD+338MHOBwB3fy1+2
P6DUU2mOpcCW2YNZavI5rYLLbcgxXt9S1LEhomcEjBlz5s9HuehylV9ZEJCjv/Mt
sglEKoeq1PqdFPYpPjmpvZ9OQzI8pbGiFjy1G/NirvJHnd1SuyjbXk+igQ/mJADR
lX/hr8A/PjXNtnVFgi5fu9ty2mwMK/BcXdSXwaaW54oXLNHs+icbwTSzyVxpqI/0
uQByPgrollW+1SKRNOcqYVmjtywipiDAZxTyW6sR8tJUYOFZx69VwfrfCZSXXqo0
UlBy9cm+DrW/LGpzbX95IH31EsnJARIH9ehVycHKFLCxnJaFFBimcfU0aTVx/jm9
seD7wEosQos2DhqozXJAw0T3Dqsby4mDG+u4D2oewAprTG1KjETjQQjvkls/iPX0
79umRo7Qmpfk/esj0068CDBNXqIh4oMwSLcdIm7I+FXf2/2uuSaxqyA2dy3NnpGY
99+ZOZ3mpC2u5eQ6OhKgBs8jNvTz0Ug0gEN3zPx1Yd9wwXlno/nUU6CxoDa4vO7X
GQDDs4wYrzmnekegpOetA0Wjm8CGz7+06NzH45MrRD1+qKTKSnWGbeU8hmCzYs1Q
cR7P7NWSSVObnBTBNdOKdTEXOm1YVuEXeKzJv1R8Kbh2+jIQUToRUmVV+ETazc62
9nzblBefOX/Oxk3DdcHup/2jksrweYUMA603aHmFjcbvadXon3wCzYm2M4/mt5BW
J7IInJkl00xqguza7k6qNNizKlyGblxcJCv0FGGI4wnHkORV95LUIrszrc9yvKeD
A5HLVvZUpU/yaJneQ+RVqu4kueFKdK5tU9qgbxdxyDhG2YMJUnEcJAmu1jlSti+B
EpNcOZaKwYncC03oP0UTxcN5voFVwkJhy0GZtOF8tU7E1imaATNDQDHKftyQnj4x
gC4Af5MeCbjD4Sziv1A9hhukW6q/TMfwjASB6PodHQERTNRVI/vdofMu8wghQPaS
n32QbleGs52zXoskuBiv6Mai8YSSqx6UHYOzRBS56JnQcjpJVyoMcLGhHA1EKGkF
yqy/aYd434kjn5tKKxDSLCx6g+Vc1ehaBOWnUnSBxFciktkU7dIOcPioVf8OaRup
RKjKyoQ5Yjhj40JgXwCNBjpszs+rZ3LshmcRCJGuyZQtrYwN/N3cdylFa3rHTYu9
Jw4xU3yY9BaLzIjUcn7jGk1v47Uc0aQX/4MCZnLU1UgPTA/QbYCTLat+bYUy0ZBi
9UKM5FsR61p6FOGFJX3eGSxMA0+cKSNBQW/O9bdCwnobTa7RABIFjVKabBP6RXIg
yRjk/ZUmUOEWs2c9EVQYpXlfRHQdDG+YftlqyR+J3Kgww7XDic+b2M/SLl/KtYFB
lM15C8xbp5tbi559Eh0g8Bq681PVqQESFiN+PEdXHqJitVEv7PSzH5y+V5Fgglwy
+cTrgCKGvyZZtpyBICVhIb9fIjaqYq5EoGthcS+YFJIfIlHN11BSZFlpF65445bw
9BIOKMVlp7LmDZc7MY7L6kEKpcF6cpxxNJ35ORCTTm6Q0neuzV7WOrZwt6U9phZ6
Kym46fybDfx59lSVnw/C13+EvgSRRQ8tvb2jdq5zsyu8eHmWENIyCXI4v/M63/kS
7V6T/YiO54ugm9IwUHDHi+J4QPSY/qBbSXd29WnM9UXiMPvT89QQGdsngIgg4nZB
T6YIFQofJB8EqLNtdmqXNtlZLA2kalcJhRQvnNpz8lE+T0SyBsCKUahpwk92o7yV
O+LLV5mhqdSOzhyat52yAf9buDRTfdAfdrUJoHdSqGkW6+tuKzNkurdMAEN/5Xcp
t7Gu8/vFap3OwUAsJvwlamc7Y17jqJAIaIkB2xVNOtpAh16De4bbk3KdWn9B/Sgh
Dw90r4tnaJ8PxObCbeg4FZ5L/GuL2zZzNsp0TSMMekU9Iv+L7LyexFJdByS7yVDQ
mYYwlpdYEf19MF9hpWn4XL4YblzmAWh54StxfIQ+wlJhO0dYJZJR1wS2sYbVTZ9/
fy8772GIjv2wOZx/xz16GUcXsW2O37/CYQNryKSUwCFEo/a5ylzqeuZDOzyqUlDM
9e9aB0yHwV0ufJS0ARLVskoj8h6QayYY+oJKGRlUGwc8PDPVW9hS2Wvqz+BV/3PS
cQlSISBX0gk597Xuxdvk9J7WV+wYbiJWEowZVnbbWZOSwTvIo7VEAcLcrlKwR4AM
fnAmuUeoitWrfL8BLS0Ze7siHyt7TC+wSlDGz3F6CQwGkmy/3alaU81rdroG9/si
LAnUoZDO1EX7YNqvBp2/RTEoUAq+JiyI0y19Mj8jP9AXuUF1McwWrQWwrfgf5o4G
CAezXdM6zluoce+ukPMMoRw/uiuiNiUVTKnVdwNX8aWgvcoAT89ZMHCvt22QVziI
rpP+fG7gYHfTxFnNpKDZ1VSbl1IR8ldsTxnJOx5JPGiwPvLjg7VCM4WsitxuV8yE
yHKj9UWJvYQKCg0JOd/jkil1d7fwROkvSt78HtDSmYEhhaBidCiyupyxBu0WIJRK
SnGGATBeFA2B8sCm3Cff4Padyw9ZTccBlTm41v7x30+Jmk5Cchn3QOkBzbais/ff
udVV1hqEnxorxCq44RNDEkqCKVS/gJqcoeFoYL73GilMDaUA9+rY+CuKqIRNm50f
zdwPg0fp0WfDRtJEU51dfw6G1un2Nk2g82P/vii91iGUFmLDNtencleF2OBBn/MJ
nDv7cpxfi4c6eMEFXyl2tYs0cXUHnTpOs6w+0GIUg8C3JM3OqQxoBG+7giXgqhaH
NNIZK0XQlLvNYAqmyM4jJlXJ12GnoaMsM+SPwbokjKQBP7uiEH8yhSVooHBvVAMt
j8X4XHnptj8HfsCZoi7KKjfYeFEXBogicmgQnB58B0Kmh5bT8VK22gI9H2dMIKlK
FGKSfzxn8IKrwsRFygoF5kauwsuJwfsnScn2bOnSPxUWMvQz7uWXljyvPrWmQ0dT
fR3VccNCv5ByQKKoAW4UITREfoiFaugwNsBykGFhIG/LQlZTxnnAvgMfefe3aoxu
Jf7yaz5G+SlYtQV14vzdqV/9+cvNIs5NG3QcWW98NVodJDQ0wr5MugoQoTV737Z+
KqzyXITZYWUfDnx18wTk3R3nNU3hUS/41dqD8RTzL7RSRigfTtke9wA7w29wmCZx
mq/NrNSg1qzoDrEx9Dq0WvSobgrHXSB3Sav0Q0Udk/qJSfRGLsT+2TIfC3kJDsMv
PmYz3H9wN0QQegyxUPpIULBVkOLoWSmo2ck5YGx7psRiZ+UzlbqBFtM4sM6K5BXQ
D5vdyAnk2EnO5lBqoUh8FUL6DAGiNyNDsXYoOR7x1Yd4R4MUeuAChUD79Tq6spXo
3csKZGUgG+YmiP3KeRG2cLUo2bNYTYoqiDJjvB/k+68eE22Wwmi/XsCfudOCeFf8
FlRzkgVnVpaGmUk6m3HRkyRpBqm5syN0CAzty5ENoa9e1MPJ5n/GGnbmoChD9LrD
udtOOrAWfJgUMitpVhv7CfonceLF2wIXt9hl05lNLHGPmB/CthOTnm+9L4AxNNBd
mxBFIdBw+3j1VXxwLcla8EGQeoSGd22ZZqUJ1iSVnfVa3Eit00NssYjmQUfAp+Z4
oDlVMEOItJRWR3CUGil+iZ5bUrSg49bkXSCms4z11RxeSsNp1EXg2ojYqGZpm9D3
5vMq8IqNJURxB1f4Laax9VPRHCzppyHia9NOmMuQnIPUFH0ZmOxSi/pb2XCKWLZ0
3lJzncQRxZ2qGtSWU9iU9R4gCSyfGK44WQ7393FH/ppQzHrXLDaen8zLsx0Uv9wE
wHtIewHWvHBH7aMoP8Nnal72NOHHf6c+zoMjgOH3LH6x8VcmBM68kqRzo2R3L1l9
dzG82Cdsgd1F1h4F4wJjYxzlN2noxb1TwEp1mr5exDpDidVMBfux0v7JOnCNknNb
fJ/sWe6qpFpkYOyfySUATpb03rD54qmyenWw+YqWtbCOudc4mE5FUQHDYQUeyNex
lZG6j3RojogQmr2KoF9Kym7Clxo+bp3TweAQEC6T3eibXxIYh8nFNQ3pLHpnQYTv
tR/sAkjCKDRv0bmjOkK0LkQHXbKN9NwZWMM8VwL+kZhYfsppvd3TA1nnZtDp+nJE
IPgI2ocpIDFL0DI7mnRKTJls7txZv/RUMrt02X8DqBCSfcpGyKDUGE9kptetgFgt
dBxUX0nmavAQCCzdehDPxJ8vPfvO2x6IPOG7Fzl9TOG6XgrVgM/8JG04gvuZoeDV
1ZfynwPfx66Z+RWGXbGSXQqRRMl50r8L7pGlOa115Z1GjdDFfPlAalHmNtNnDMlC
VQSH6Xh0wmQvwYI6ValfYZd8UP5DIhwvUt91I/e19jY75P828KQMZ4qUdALAXZlS
W/p+l+yIh35lntkRBv0lo3KWHRik67jfI6NxjVpq15UTn+PjSrKOUewzmLnKhXU0
QR/K7PVVhM9J1XUrxlgSIAsG6nNBL66Kamh0MJgddKFIuKtpHR2pWc6xhTiTZIy1
drBz/gFCf/Faka6ddkqJvNRcaL4qlBhgzKKAp/C+K3wT8euIPBYQJyct6pz9EYcT
jL7A+/IDAO3E0K2Uu1U+48vHTdLbk3iA17YoSdhw9Z2KDKV+mzkZAdUubj1BxmEF
p66ZT3CSbP/CssZwVe/+qB9HAO4ozNYPZvA7Bc6sjw1LNSO8Nw95E/VgGwJ2wKEt
rEQo4B01pFw5/pkyPpyAarGGTqCviEzR10BGI+9M+LnMn6TmlNFB2r4MJKXifug7
7SVJZ6R0pS2mei14LCVZQNH2rkhqsz7faLRLXeofQrqxvCwvIYXGcFYmpQxOJ43K
+5VI+JcQJxK9eT6I12ifYgRfJZineOTpHzCz82zW0/f12GRobu9MJ/mkm/9zZHZa
LOiEXk64pd3Y2I+7SI/f7l18zrltw00qay2bEg9qI1BjwnE6SOONDQlu120lyU4t
fdY11uhi6y0iukJO43LPbbGbyC3LjRpjveBCH4RETTpa7hd1ioGV4a3flmyoXJM1
sqLJe1YCuVaL0DeoGjAwa4qiox6FuzAicMiLi8MM6KgtPnRXmG/xVVJzt8eSWEPv
mEvZbFi8/zyKJ/oWmdSyRUdcWJPgY9EZT0Vo/pRnppLaCvDJvN0Wj/iO/lo+3eAO
ewEH3YfH6JfV0clJaQyoNADbq7aA1Ccdbwz6xE8N1c3Q9O5dYlwCmtRiWjb3IQF0
MOQ2qYTmmYuFjvAIPjy67sUaIaCEIQiSFjPKwta/4WB5Jk9Eh4KE5tIT54nHMs+h
eA0oeB7bu3MkhLMFk3eT0MFPOFRJnAwYAGZWSYGp1MJyawsPfP0UOkm1+y9vJl8r
m3BpiigGGR/PpOD8m1sL6/GA7VCFYA6lJjNhwN5C10ETDYR7oWRV6jxNPVFCDrIy
9+3K0SbrNEM8txVbMuJAWRC8kz0OUMXmBaoozDf60rOEKFRHyj5BhRs9z6dwd1m8
73Hive99KzEJhw40oEIJDi/CWgiLakm9wcfRq2iLW5d6cSJPaX35RXcENBjeEINu
YVtAxTabq15/LuK59a0kxZMmIouS3hJYQu2MmkuLys901En1eSF1ZlEcJujmilW+
Ry6GzDumq5sWrupvdE9z8XpRaCwXkTJze+jBws2CDjrOKtxwAD+uj0QFCid2CFRP
D1fFeBhBYHmb7dpVITOyiisU4u328cJ67OjpyIRHHu01ktV+fiKlLmKP/8u/O6rX
/orwGJAiCxq17pENtQtZ7CEJgRY1vNKIVo717KTCbv3RguoM6hNk4b4rNBiy81iZ
d+ozaORwfbBW2JNkisNlKTTE6kpySk6tblWp8+cFIXJoIVt3OciTJr6kY9lLk12/
nSLkx6AWNJRHHmPh6dsvMVBvAZMid0NXn+uCV45ydV4vGlqUPFv/Yt5aPKa1Tgvi
L5T2gwZGisge5lc5Eiwl8QYJP0ghebqx7Aj+hs5L/kRael7BU9jC1w2Tyiu6mjb8
RUgAHipzI99emULcCBWpjLZAaA80HzKlFh0QDJHHO8L00OeaQDPqeeIBH+KuB0Mv
peAnO/F+/OOpDmjKckYLMFBy2w0HcP2s6ebxF+ZqTot7ODy1m+ZnBfT+NmNLVYAf
tjfr7jYfO7i8HtIGSWCEa41z+ovV5RyHcQu1mrnVAi9MTg2beKsKfRHevTFA0lVo
SIAN0QCKwSMmgzTBwfUJiCDy1DUjgMTPRiaNT/eX36ullzKGH12ceb9FuR4nks5N
yyjIfDCViVfr6VvUTDLc8VsMC5Mpjc0THBxUE4r4z8W8JPZ0zim6yVmQjgt6xQ57
m+MXx/nMZVlOUY/hlX2s9YGUyzZVyeCzQHnVwA7MulDhIvc0ER3ih/TkIiiog7S6
b0ee+A6IozWxagEq7rEKQyM0d+TAjB3h0KB9cqvVSASSfJdDefuDm+zEnLAp/g28
dA7fxFZk81capL9Qr/wIGKHnWI8XqRGL8EWyJMj3Rkdj54Bmdk4CzPsxMQKQ1PNG
4Z9synG6nd6wqeZ8ZnIZUyy4szPvRCZ3mxJvUZGNLGt1KLItFR7uvW1t3JWwblGP
LOYfBbc6lIG4wE3GZo+4RND9IQIGbRFIncIv16vj4/9YU+juKIhEcODmtIQLsxSI
i8FOIzWsTQltXgkSA2jBLEiWRFFWIFbcr6aUs1/Y/oQoroMsgFEZxkIaUXRKqV/U
cyrm2VKGsi7T/G5rpb3ITDvCpzsj7em07MH1Hn/pRR4GnjDdhQwuEgd+6OLFDsnb
vHCzpb2uu9pWHUzuDAxHXkPrYCCWRFLb/TMRhOzTbT7oEW90PZd/iogKoYrdF+oi
EeXheTE4PzxocpuL+c71Ih6HUcDXMO4ZKHdo/RdmjLZVtIB0I3xndesf0Pr/F6sR
e3zGO+o7B24VetBD9rtSUT45lAYHKJl1pbO0Lh8Uk4Z0tEveFf8JTChaXOTIiv2q
NT0+GhY3/91LY93Vf/YLcSLv0EfLyGgAa1Kpucsn3ww+EQFr4wj2iDe3/d9UZO+Y
H46V7wRmzO3hXg8CggVgOzApQYQOgNYPDuY94VA9lzini3XoDxePVK+sPY4hKv6k
Dyf3lPkUV4qaFy2qjRDOLvRlRKNRli3DB45Lf8RZNgGtfS2qxL1waw8ROkZe+lVa
lcuQKKCXK2NcmRkGanba5IRcZsBVDOdirC+4TL9zu4UjqFXRVf2TTIuOv/ZwNu2K
RfyPRhuDBkhsyUo0JO2PpKLXAkQ0uQ4DiUWItQwLA20mYIdbrP1ao3ERYozjDOUJ
qfu5l2Ux35iGnRStlEKYBpUcZuYuh3UqR7qd+nUKStYuEpug8BPElFzdPViN13JH
DDYqL6ysFjSAz6spgrEFqmIJvpLfdBWxmSco7GwQIr8Tf72ewJo1pc+dJAqwaU3d
A36TJLrl13RlgnJ4UaWEUlS5w1EYJfdYDhT+SJb2dWowuAipekyGM22jUL7cXnMh
9CymXevi44Cp08yXTu7zVQRlWTaKGWMllU0N5rdKB0n04Y3v59xypjhOriZrtCHo
GMNmy+4hBbINik2LtgKvVVVD2JxHS8sVFNHY85KZGqfjRJDN3QGDipEErabxYbHb
sU1Q/ArAX9ji3+GnWfNt9LmvMDBMt1lALkPLdVJmjtbt/ml5HEqwKuuwX5mvx5OR
wrCZvRwU5Kh07S0OPEOB0OrAOvyC0uMk7CkyogZMNPUGR4i6t71FgtuKfyBqlusJ
1p1Oxa+TeKUmfwQpBYWFY3JOdNlNXIU50o+JJSTbTDFC9Xbyhz2DGwu82ELLQBJY
ZNuAFnMEg8DcsJwDzXE8wNvlfxuueK+WmriYJC065iZ3od3agzfO/XtR6N5whh0q
yOIOJ5Z7jX+QtL1bfJZkeuL8ZBK7vDihYeb0/jbiU9iBXUvslHPBt3qPOG3/6mVH
211UbE3sghDFnFtepljtWb7SAzz5Yggzi5XzXESS9krqiLFzDwdQtQCaFxRHC2/S
6ww1i2t6qT2yMkCL29tuS1Iw9usSGhNoJ53mpmHB2XJ8KFIkfTnx/8zuLl2q6P+a
V8Kasw44iJ1iIFKKhaztSfwd8OxxIoQmrYFNdKGbqDdrfGFBF3s6QGAFUDZou0OR
V2T3SIAVpvoiOdkAo81atDtZSuMzV7pbK0qSzXZhv5Qtjtf0LTHlhoxDX2w8xXK5
H9cli1R5JnA7KEkbpEXkxdn6x4NSumfxAQhFRIjqfLv3c6VN0chLiy8IRMuIdyEw
kFwVnXCGKm9J0jQXmdAH7PvT2/DwJwBXBZxEhftEQM0/kro3RInDtzwKhbmNLrDi
agsHO7szSKd9aX5yB+wQmln/r2nwcek14VIntP5ak0cAWQp3IfxuBXnY46FOqkqp
VsWSC4chJHpCdaV3qj+GAmhogujw4Lbi1YbUrJue5XbKt3lwgBsLv3gK4iEas73v
bQV5bNMmKKZaN0KQf8ViSJV87dFB2ezyCx9So0699OmeXf8wh1DwNXcZEdAg8Cjd
xi2OkPtAJrcqB9RjCK9fzBMVyJ6pyg7BePr27quOVfsy1O5+ZqlJhKrwVqIOBRBE
t3PKS2xZcHmY6qvCSPOl9SXgd7xc7iE8DrbZXiMZ/j/1wj4Qily39o3oJBX6hKUK
qdzqNqKylP93kiN65b04RZ5th+PFq1IZH+XaKijh1G1eOlBYNJVcSoG8CctaLMJo
PQB8kmiTreAB4qIi89jT5z/vwQbkwlrS/BQepfk/W9tTFUR9VIHx3S12rmozh6Di
/btz+o5SykRh0ar9uh5zosPUsKqs9Fe5qtSH7wHin0VAyucYlXBMRwl+jWOzpA9S
BCujo4wXk9HAJiifin4gHDhH3kMl2u23hHqEvaYeQ+O6wtLtLqFl0+c8AfPkxg3c
kmywx5vFG+jPB0ue0QSQeDjzNy5wDrj4fuuJkNzcPfhMpDzVkvIZio1rtV5NV0HW
RspGyXzisw+kBokB0d22s2PYqNvEOZmFbFtf5QNbp8JExaWneL1su5FpKoOynuaz
l0U9mQxHYN0dVD4GXBUUUbJUvay3eFjugRivhZs3rfRA5/8RDBI4HPJQ806yAEez
MrEOBLudrq50DoliZKtldK3uPCMCZIaUAmKJO4tB6cFEqne1IaAwxebOfkhlUoy1
eWFtwzLIWFOKejLQG//AkBeyIwGKmHdNJwO9Et8cxrJl43FpT/5IpCT6RjZIQtPK
v31953jalggu6f+c9yfbT2Hcn8+83KESCluJGLyR/QhdHtjzIPytsAAsroFehT+2
jdV5WUg99i7XoDbOqZYJYi36D3pTzbL8Bj6pXl9mEJDuCEJukEiJB773cuqnw1vm
MSaqGWY3qRl+G+DkUYDzJCbLsGTzXc5zfs7Ms1EKNDENkzF1V3lEXpcepGy3znsD
Tqhr1Qr3ZsLb3SM+z1/0KuXBhYMMWhngK+tnZ4EOzleKW7VXgQqM5cKHi8zd1/SK
AQJmNfwFWkV6rrjOMhZnfcv014Pxdta+Twp0W3i/SEvSF8BDj0CMSkFieNx+dMbc
r7/tE1rZaBoNfULlQhZiGoSmjD8g6SJG/pdIOr1b3mi1ak6ut02X8nxBTAYm8HkY
VKpiWuHBmVrHQJr5W54PKOdQpQxmCDu6vFVbIpCSDKO9DhF8WPgBB/i4+qjB+KsV
t8CJgr1OCTi1VzvZN7evXMb0QxGGAOjzrD5zUptmXOCG0lg675xKGdXrGgoUUHGT
kfT5M9dMwBBKeOqF0bZCMhJnIawwN9pNeBK4ysWuDuYbDHNaT0NrfJa1Y97mvoWo
xnmMxPNUWPWXjyWlGrp8p6OvyUt/iPm6b+4vC/ex58EUF0L43QrYZSXQi8pyjJ4z
0sAPAxVG2yjD36bxJhrG4G0nsNban26jElqhoBw8/HW9RoQ36vB4qXMPy75sJ8Di
So8fEb72yoGNbuCF2AeqbTkvP+zmvhbArQIHhh5mCrAXWRMWDNJJcNgH+RMcANiK
iI75Vh/4EWqDgky3HJTOnTv8lfm6uHDA5uktBnHJ1oaa17a+ykvA03UXXhaBh7Vq
asyMxJlClhxCVRWj5gfZDOvQlSkFsAE6e12dhew5epji6mChWVtiuQ2mP9vNMNnB
M6h0kHVV6e1zoponWsQC4jLWptKHjbc7GofdgSuly7p2V2Nh11V3A9qJ3K46FREG
JGpr+dYjSxnUHq/jNzR9CUiM9VcdhruhjdBSER2v/WJgz2TUwqYyGJVN8htYjlTy
wwULe84YySGPSBCoOXurnhit10Uc+0+moKc4cX7M0OUgQgFx/6N7KlI6V3ArdGH6
yeltqTVsX7X7XG94v0WaAbOUSIKR0FUn2NfHnzA+n7CiuNELfuBGP0IF6/dLDMom
DYlaM4mU/Fye0S+SAFrXUDFGasCJSOUtUhpSa3Mdn+/fZckeTZPRxv1cv6JhpPVL
jSzhV+eI3jTMGJV9DR93F7ZhP+V0w3Q0ZyP6f+y6RyG+G+Zd1DPD5krhgGKQj+VF
sWEzDa4SP0wuV4zYjYZrHM+qNFwIUya8YgPC52jx5aNzEVypdOJ74L1xUbSFCVqT
/l8sLhx+78tc/6JGWcsYp1771i+H7uqfW5zDtHApqUDJDHRIvTWxYEiHzCtBQCd9
LpMFXI598xzH8mi0kuL7rshI5OUGyfDRur+jYrIjNVDtYinYPPcw+4apkv6zfW/D
SITceT0IxBSj1hbXikm+jLa7MFg8U8k96hjmg4NFjnoioPozXAo6RgnugqsV5k1k
9rJwg5U/q5Q/B8Eu6LqxYdp1uWAVngyG7pyYrTZK9YM0K+sntrcfyK95dJksRiqI
8eKgeYLAdGDkNAO3EE+SG8OxttQmxZDdZ3LdnBqXd1Y45Jox6bQd+VbKDUIPZ163
eHVzIaUaqFzYtZUeTeR9sh7quyjlxbJfHVGVlbrAFezWSU+DV1kk0h0wIM6ML8CD
Ua7iXNFa+2c5NIA+JApk0KyZ2jSKvlIoLkStT3sBA6cCTlqxpmassG0r9RAPeo9r
aDJY9ZmhHfa0fcQ//1MsKg9UvJDqIDsc0b6YZ+A0v1FCuM0OEQvJFjdV2srx5lWU
6G6q8ZmaVNq0WGcVgOAfy4mVVf4O8Rvm8+/2JxVH6R2o3nbivbzVIuumqWyo0rQU
ZVxMzgABfv4gUvBTQ/HDDg7VZw9I3myhR64vboavx7Nxa6/02KQ8pCYs4CdcfLsl
F9KmM8VvZoinWTAF8yD6tphYx3JWzYR9CG+QVyAJWTlWt2rQ3eFArqaIaMXw6icr
59YqA7kEzpQQVw69HD9zTvGcRAKFyab65oCIg6UwAjk876vZyWcGHnKrUsNvjwv8
RWKMuokZOq92EftZzMhQV4Ai9n3gd0OKgxGTEkkoGU0uWUKMUGYw/M9WXogf4Y6N
XQTTbYg+SWndg/Mjqtw5uehxptcXXZZAERg7BJHRuLi3cV5F6NslqVY/lrCq61/C
L2ykSAdcwEAmODLQ60J5Pyjp3zJyfLXlpPC0FXbZNtxZSRQQUNY2ks2JOhLFgtnD
Si++nvBXie+2b+Ivg2jGs5nCGneZPx7dof9qlQb5hVfapOAFxB2S/oMEnIovtJU9
tiFhIWkswfE8kqeGnyj5XAbOIRIuMlaBtBGkufog3uX2xYkyfq0daK/Iyesc3LLi
iMRxtdcvSFDn2QcbChfuDZ1nhGwmjFY07W+ezAWqE3Wy09Wm6DiFFLqLzF5k2EvB
7z/omj9RBW8a0URUbouuA8DiKJpZonimCr1K8RP8U4AcHv0y3m3lJLZrc6QsOM9H
Tw1HQTlM0AwU3WvcL2P4KLjDkQpk1dvoPkHrRV1bnN4Yihcr+/7zV2dcCYx00qmo
5Va0mFoa5Gk2AYkvUzUESr5AaMuhpalqtRU+jsMtEkgfCzCmsbVW7CrqWPOAVCZ2
vXM6qz+b4GZPgBYb8ET7cPgaj3tT3EUfdUga4zZpqEp6GWqPeqz/0r7KqDQJ4l5d
R+w4pdmG0f5Q0z30xX36syCZayChOuwGFa/DDDSBfj8ctCecTy30fDobOPFt4uTH
2lEsTyJ9b3veIcHgxLoRpBJMIRXIHECjHPkYtlMl7XrwOBWDYu/wfeH/Onsy7QZI
2JoiZBLHK6ElNytmBjDxFrwUlqDbKHGqg3k8qDTxcupfu7iTFx69utrhs0ct49at
UXdfkYCwgfukb6PWR6stiuDqSsghn4ghysFNu9LKVCXlunZ3LFr4rhHZUsAjFEep
h0djLqmduRCdGjgBcLHN+dBQYqWyUwdACUs5yB3BQgbl8CVIbQlSCACqFvmv/CNC
K7qJ4iZRSaXL+ZPeBT2ZemT63mlUMCrgbb9jOOEs4bYnOi3wfMVOI55gs67jhlsa
yX/kqoKx+soJJd3921a3D8rpmm7UtAbDhC/o33JtrJlPlQHu4RdmqAvZw+mc5IcN
NyTwqd0IDZ3dJXQL/lC6bx9Yc5lSDMkhEFnr0hkEN0krYqpWOCyUCFqt/nmK5SF4
KZYUEINX/HNDMpopMPcex9JdndsfETEMtB4VZIIrWWCwhcQoVDjWznbwiEWhfDzn
iWmwwtWBvyRiFcmbtxUuaX5ECDL4EedlXN+ttazgFTp/c11su+bD7SYeIOGCo6bz
aOL+2SHOjvOIgj1BrZPvlt2unxjoOEshYHHXObW9qwIhtBFRw27QHFGBbyyn8eji
3TyN8IONxkR+RkxlyaIIf/WYw5lbM2wnhRn7xIdZU8eANzRxbMk88nRQsq6LlvDV
7rR9avFIAXyThBqAQevPd4V+ghwPTThwHcl2e7w3cXCa9q4Ek0FqFkcTmw9JLtmH
Xq0Z44DNm/JmDKqLOY+2HNU2hid2q2Q/Wil08lLNGJcOWVwpmC2DB8FZTNk4dygQ
+ytRvHlTwKqNDqqTdqsdLqv19r4bY5iQ84d15+g2oMWzMzDhKW0pgL1CSHJi1yu9
ZCcpBF0njlOljk9caBKNulVe3cT5YolQYQrG2eWD/AMQxzvD5Qyuye1zimAYgwUj
uOzPoB0ikKMZMD0kLNt0DShLUSbhHNfciYlwqkDWh9VJWMMQ07hlZZVKRHcHaemC
sp+niH6ZGPLreWPkx7X0WlkbjElLPxJgyK+cA1vQXVWIkeFWgiLs7vvuPP1FavL+
OhGsdBn7LTrzq+BTj0RMG01vpAQm9/Hy/GP1HTVLPj3mmysDWfdZ0gGf53Cie8h/
sJIzTvHjojUWz59vomWy0zQqaHmSZ6f09VYlPS5nxk+MTZ9m37AezeHx+YfFWKTj
GKkk0vMSDalIT/ZzTYwAwX94gualWrcilKcVrmmA87P03AaAfoqsLiAsYffgtpWP
NjjUtvZfxV5q2AIzUfQsIn0ZwSZc2KF0gzt9vEd+YkzmnxxbTrwt6RI8jixbqiUm
sqo+kMPNSt0lWftvmQqpCF2ACuJI29ebIx1qOLOziwlUvF5KsGHIBVRJO8+DBfYV
FFbAKvZYiTelZpvH985Wg7XWRdgy8QF/SLFPFKaQ93dA6QVXELhpbY0LUMIIpesw
RD+jsYgSUeFSsfrcIfMgPbtNRPLqhejrtn6GNjP739AZJsTnxB7NQsP326I4nyL6
CdiQ/r8BDmPTrGkrSrbxO1IWcU7G8Kn5TC1oeJ8evJl+bFRCe/nqiFWvyq/A25wF
OZIXdtibt1+/ckCz2xUbIQBYoN+m2ljpO0hVQE764OqWTAPQbvgfsbdyQpTxcpYs
NBMcrNbsCdRJHYxP29u8pySbtiL7vBCL/iZtXc1hkRIo8D7y7ymGe1UJ6CfV1YLn
qLk1GivshZNoLFtPntlvSTV+/OWxjvRpLsMDhMh2/zS+HQIPJolUpJ5lY943p5NA
eCein521Eynu51TPHKwiLyIHrmaUyrilRd3G0BAdkd5WkX6iW0DZWmUMLmNOprJS
/2UHResC9x7OrXrzceb1nKaKX6f22yt+6Sxn/ZAMZGO0/HfRPX8D40txXvi82/y5
aSpeOVFCKwtvvb9NSse2aHdwNJ/F75ztDtdiK8/th1oVKV1IXo+k5VGl0aKMFyTs
csAmpn0ZMf7nzloVAKLKnjZsiQnBuMngoiCgh0pqJth3JaV1LC96xrFNBIIcqL0+
9LS67YX8iLbdnVP0OQqchp5bMMi+2VafCWooZuatyg0ahLP0KuDCTGX8tY3o7Vln
meqyETY34Qmplr8ejUMT5PlKy9EMyv1tJI4iCb6kLr7pplySE324I/zIm9uB+dpu
o2stFc8lCCu0IUWrXIXTif44IMjae4YNcxvug6CVmhljVjDsq3NmbOk3dqw/JsJE
fAdak9mD6snnXLIaHXzG3w6lM3N89/8lno0zs15oRontJc399e2IA6pgTrNeSs25
hUgpYYo7NLl1EoGeqRYvY0im28ovtHSS4NBZ9cmLvzJSO+WXTD1id8fZeNtHnZP2
y/1spBYYSyWnhm5ZY/avDnnoKtdbW4W4VMguSrSdNfZphixFw6BJAtTd5FOTgKMY
bqzpzJ/W9UykOqsGh8ET/EE6ke9C6cwDejVo9Es0WYqfYsgoK9JOVCKmYIpGaG90
69mky12QC4LxB7D32lgtHkKJ+HTbqRB181VUz0hHFczH8HbH19GjcXnwUjSdgWSS
E6fJ/uH2hlU5BM3t+d1W8qLOvJ7IkEbHh6ihw/x4kpghN6NXFmq0mc7i4NKuIH/A
rv0gPkGUO1OjzHPEdVbs2xMCGjMdYl1YwRnARF5Bs/xGEa/eiUwGsvty+w31cW90
8xSKq/Ja0SECZjO3kiOqgotc3sdVGcVoRxgr/MZitUvmEiGmpOHC9uEpy9cqA9k2
VtUqEqZjtArb/jUUZQedqCLaxWZngKwANR1UsOp9Xgs9YCun7+Y4AjqOMJPCOTfd
FgAoG9JnO/1Qsb5eaLSvSSOFYOTCFocbthlka/HFT5APL1YE5VVzjfX56SBKxQYl
UMSiVLXnAxlvlZ9r2T1CMW23/IrPyfMJNciluW2N7MmXMnRYU0XO21LrIStD2hDA
iibAadpHMS0iSSyAoQRn18nKp8LPSm3Pnks9R1DUlq8pf2WebkukaL9yZuF8isfK
NGP69I8V/DJUg48xkQeER7DZ49Lukssml5xQZr+y83HgF/R1hXeQVm5dkkocI97l
W3TCaURJf7GWjFlcUR3iV7P1U84u/0FJqAiUYprLkIWEviEsBAZa3eFrn2n8RYZy
pU8qkF/s242KsVz6fLxdMnOrSW+3T15AI+1Cu48p+7q7liovVHSNxE/7364l7EgU
4ERXqT9XPJru2A5K9w4BVPSD/gf3a3f3q8rlOW8XQkIFAJoJOF/2DrwusOZWGe+e
ln57SGt7bn31MCIietPsd8anmPG3oJy8TIQ1U2NVXufG0Wq6r2ISkGpxffm008WT
BZiLVOV2zHdDO1S6OqVkwWW4g9PiWMvmZpyI6H8DmCPlba/nl7th0OkbgGepeWLr
od/RUEoXKnY6eXj8tZorHcML/z2Ik+rMWjI02cked+WdkFZLHRF1xFHVMDv9p3U/
HbOt8Ccfyd8dEiZfg4/CogNIXAhiOUZDricHCOc0Vwf/YXmkSTTVQB8Ge7PJm7dK
Zvvu7NgMUmyYvxt/j0GSEq6RCnfg1msKZ0awpBVZIq5iG4P/voD9kKr134rLI4ZT
Mp27x3U0L/XpZGlnuI6ooVjfKG6C6lqvJZ7oksw9i2DBenZSHL6DbcODEHmBCodj
ucV0B8NysyoUgFl9XCawwxFlBr1W4KF7m31NAidygun76mJ2yFiQ6dyd7DYQtLX+
jli9Di/qgXs1eu293b8QOppK1QigQ1chAoDyEa0/OLNyuk8ZS7elXEVUdknwAENs
xN0v0Vj8XosF0qjyg9Kdm1FpR18MhT09U/0cNwtuKXEdznrFPVUoUpnFaFjdWTxb
kF8Pfw4qF+KpFXlcvqe/68PdEX89bvl0A0jNYm5dsuHPEEpVDKqBc0fUs0t1et1h
OgsN0ZbERPWxBlmgtTJQlNpZNGmpGiOroB86J2rTHG11lsQUhuYEQOuKqlmDmWee
WaS5suwn488BEYL1AV3AkgkYS+IvU/Sh8UsojWjqV3Uf+qD+HvZAvGVTsJC1buus
VmAhm3OiadWyh4GYYKv639Wf1bUQv84aspFSwLp7PmSACDINjPLagCSJ4+s3YuoJ
KIQGdURSHXlbR1RlnSG0iQwBd+a7rGxgtp203F9bJK9o3R4ICFzPV8Ta2GGApVvc
D2aLrt6Zt1/KG4zb1CcfgFux2Ni6cUPX2CQd1105PmUJdebi3LStBG46AUXgpwQr
BhRYwO5KV+AEuUvBEEBi2hpk++fqP15IfYRSl2Z8eecDpXJnWCOGu27kjjgIWSvY
kx9O6gFmMgpq2WMbBb/JNDcsSxaleo9a1Ap/+rbqTBayFh+0sNgDhN30Dwc0Nik9
JufP16a0or2ycLE9C0wzmqSEiC5wRAXzTUrOwgL2nAqfB4SzFKoC85SAjCbVyyvz
/jJ6Jh8q/uc/l60xbYZ921Dpos87g5clzwTaa4Wp+7EX0NfWXW6oDhQle5smyU0R
vw8oc+WsoDkOaZ2boV1lILfUW+xPjCGhwKugrGpo1w10BpnJJZ1uNRBHALCMeaIc
nJzgk/RH5m6es0Rh8Ck0MtyMDjIA+0hicEOmaUbDyDlZYfB9T/h9nG0vYLQnjtsK
gHH5bi4edA+L1uRgp9du4bAWkWaY8x1iWIZrT3fBRs6AWbk6YIjrTjevrQbit90A
K6ZX+7CUB2OuAULTEJ+5LhCcXybQq7wjZwTpyCxsip91Dt8NjHkBfOgq5SMS8fzN
OKYj3tSPJsBrZ5lOoWUaHIez7FNFfYdvCRv1+7/DiwS0QfMpXqJ7dddRR44pOmSn
f6TS3i/Xh3HJsJCIIm0PKD5R7M50+Nf35rkSIkqkmoEluYIqN9ZJnpD/0eIRZ476
FlRec6b3kDjadcOz5BE2VudIKF+fvq1H5GRiqP6FAbJr9k9HOo+ihc8BRPu1tWC9
/qNaLD6iiT9Wjwi8XcMXlJK/ekcojgczewTw8wEBTcUZ1T9bPTJS27z5GPiQ7v++
7ZG0tFvqvrRa66QC75vLeQ8tnk47SZ/gkdOtnxwPYK8OYW1a3HyINTju0L0tPByD
jYu+AfeUYHa2kydvDbR7K8NQGqJ5kuGTJmFUupbB8Rf1g7+QrwQF43shcbmH8pCi
H9YPQbP5H7xGNQHDz1N4jaYg23VUYI8NUgWc9Xaw7sOCGDDyUbMYMIVTvQs1KQpX
2+nUrDIijXtLXlWZ9iiAvzBvGAVBmP/Ds3zpSzSkoHtn0rPzzMsPpgFAmNLiI2CX
n5PD78dMKX4cbtwK1/0JQ5+MrrRJShCWR0/8KPCnf0svjsJICx30yiyNKJHZSHrD
JDRqIV0C4mnarltgIhaY0rBy1O4Mp0omgk8831I2lOAM7l1uytc0q/4dtGOvRtBd
dRdH7FxPyDU1ia8VY9MeIMfCtktlZDKDhYLMQaH0A1Crp7fRVYLzi67ojfHSIsO/
LdyenU4mwHHrdtN7eZBg4F/oBdRAUKpiulVZsBNaZEh/NeAGgdGIeMVu/0Qhgu88
r53aEvjsQk645poz30owdkE/NWsciBG99YrDr9kDQRV9JdPcD+ibvgfM6jj7eMhn
0kAt+HImE2euj2Nz1sONev0uVjvmQ9IRcxVKvV7A1kMjFaJJxr/LYD0SfQZC7ZGc
7dba6Hm6ZvYfHUsHKUldlU3ENCruqPTMM1q9CaC9WdxHuVsxI9volTXWs558cJMJ
u50H45wwfkH/76dcVBnIHjYPYCsiB6g07yL5r+5qT4jSefuam4qjQHi2CuClB3Uo
HkXegzeHxAX497aloKslSe97M1zGLzwvWGd7qXpmFBO0j4/B//Z67udxfipB5A7p
4/ygC8RX3Hb/3UvUfihqRyIOXYiNAfaTQmwq4VHPvi7VjAaHIXPNE+T8m2lMVxVc
2wslmQNPzQNO4C0TVrb1XPkZm7ZjRtbW+3889Rzp14Im236Wv4Os03aRDOdMqmD7
iizgW/XoY9z2/uKBwMXFnBwRSnAKzAa4LI4TaYU275U0ub5gyskqY6gE5+hnp0Zq
wL3AAqidrvVXGLVS7PDb9LEiPKfn6M9Ci3rb6JLxEnezpMgqVyJeUcMC97TCsiWN
Zhs07BzVCZv1zMr/9xLa0HKqeHwYzTbpEz4n/KcP/lemPX6VrNkuNTfTZZAyxjCf
tSLjtt8We2iERqDLlAK7trhXVueqtHTfPrBgqm57dZcPJjgjEIZRO6g+V+jTZ+QY
GG0CNU6l6LqSkIsPOrD/rfwSOH9Bu0E7UYubOpRAci2pzdXvcw9mScDmV+OhGHhh
M5lvdQtgdnUFNIMetnuzsowrVfbTbJOZ/9roqL8Nlb7B1XVc0pVM6UyU04P4hqvh
O5e66wp+MF06Y0+Mvtkg2iAmx2ennArfPzD6wpWbrkOFLrMzaOkyeAiIHy1KqrLI
czT3w7KQ/BrdlGWCknmlGMQIz2NdpC5KocS5E8/TyrDzTiEmJBawlL8BWs7Q9bl1
Pxh2llaVqrMWV1ChqheR4E8eWyZl4aDMEuEbU8cnmlKl90yUrx3a0DiUqb655ItG
YmcnI799Herso1bO9+5FATWgXZyNEbBdr6+8G/aW6IA3oHLyIpFDzoZMY+fozi96
9fT4UTGdLk9+qIeCDMfUoKw1FsAyasZCTZyg4fHoMnTiM/31cT2g9aaz9DPtFys3
puAxHDdgTx5mL7LYHZzFGlnEHjxDiijA9OOkWzlEKS8ULV4KGOfd++O1ptnmz1eH
vuog/laVjE6X7Sy20w8HRgHt6yvoGeXauaA8ENYA5VD7nCVRWOgTk0JOGNK5mBHn
rjUWhXXhFfe4wV0nRJ6JSO2+I3yWK0vx4tOypGgV5ieetWUVsUTI0zS0boXkHDCo
q9B6SqBRqikLLB4fogBVuzNBT2AiC898kvHHLe5AAIYATWZvskXlqW48JivSS0an
FRQbIU4Tmkdum20AJWsd6Wtt2i5qlRgq2NOzA3i1xkLn3pMzn7vvHDS6ON+k5p10
LQLEgggBehLZ9kfrySbq3+cqXiVAYaQN2Ykacn7sZ4R9Tag+4Xs5NRrxGWv3Yeyh
E+w+la/jwoImhgxKCY+krHTc+KzBVwMESrlpNqzoF4GBS4bgtvJk5kqiVg1pBODn
vObTxI1gWIKr8FwGugp+4FdgSdPIlTpAPKOojm8fsS9PZ3N4Ng/2uJGIy6VjvyNp
GL3OAEsT6vVSB322okl/qgAmov5lWOcumE7L+wMFT79OkLWGbUiqvNrAKj6k+dod
34IfcVUKMdeMJIYvNY+Pxjmh7E607C/cr9Ws1sykt2yvrJ0n7I8TWwRk9WmQJ4/l
gh8yRt4nPHgXRTchHyngrxxYd62MS4tZNe9aXyKRkq/T/kSppShD+Dv8Za4Ib02Q
NQXzjBpPli+GkOnTo3mkdHO5b1v1LydQ1ZfcG2hW0LypZm+9tYoXHbcbdpV37tBB
DGR16ifUtrPgTpRbmuQO1pgPh8/DsQNbLg/rVNvHE4vJxc6Zco4eI1p7h8Z+wMeu
7RIJXL1MSxqNC7W81wDhF2H+PZPspSZnZfoMAp10weRDT84/oxK9ZJah0FeRHBCh
8z3DQvgZCn9hwgtLM0OBP2SBAfoA4MSTx15dBK2psxEATqXoao2vvPEBEPdLmAbh
zxfra89rv9U4L+NnZvK84diWFrhkBKlNz/DubFlIDTv65MUucsTsVPzM4VOZI8Oe
ndTywzX61LRWMVduVbpTL96rYtzonNR1uuCGHuH/UWCYlRYY/Jo3kf+BBbZGveHM
4GA9cRBYQ7DciwX6UJf0hCAFUThcYRzmlIfFPLXKVmpHTKvpKKuDNWdV+UTwtmuz
d0d200hRFnw/ZUBFyD7sIQwCH9cpPU+pVL6rcGK2jIJGiOFpv0zbx8cPm6mw8sd2
R43OX7JpCC8AYTt62XToCx3tVp8euTUf5UCgbb2rfkYS7togLIZSvAZLhvjsUpuI
V6TCE6qDb/4IZbdULAsgwR5YDzhiR5Xf/m9g0wD7bB83hwSO8gcrlQCsLXfGuk5L
NrEpIqm30mShYp7JQD53n4WftiPu1p4DW2saMVBay8/5Izacrn8Wl9WUW4MQssoJ
+3MI467kOfGDGsvH9RGkC5hyZqP/hOd8X9LEoraTdTkawmmXX+H1ALPDvAOy5QKi
9RVicKUQc3o+2yN+O1lOa0gSMCowykrsSrZt/UpI2UufThuzoCqbG1YmypDI7vA9
WHoILQPW7GjGtg6+pjyOXNii7d15oXe99m4uBRmCOAZT3y/SeZY5oO5UISLu4sLh
6fnt0+LOBBml/9zLV3NXhSrAGNpkhTsVy5KgmsCFxekfSjsD7H8Ufoe0jabgBUkX
usZ6dvNpQTiBi/kc/s8YXHihQq5zz4FgMMSl7f9D32TAM96yaYVNWWoe6pb9V8TG
gT5dI1o3Sx24w2CKQzlN7swKOkbU4IoHohMBNKOsI02dP6Gz3KDw+PhlD1AJgewB
7adVgF4J7s+LUHkEkv0zTG653O+l5o/3k9ddWjKVswQV1N0DJhOvfa7t6OWBKbs9
IM+s97WQGkOeJwiE3xuD7E3XSmqtyYoW0GNjHuvrJfvuxvqaKRXfynRWYxs3C3Sw
0qdVtEZnPTbiGe93RiZFaIAZQaiSuWyc+4I4zAtJobnVGBwYtRqrwE9FKHhMrd8r
3lqfbaZXQKF4rjVjWawyreP8AivKzy9mFMSasqmj1NpE6s1vP0WT4gEhqAh9ioNf
d1xPUgS0kTcp5wiAv6XpP2CI9LgSH/3IUwidbO9F0IyVvP5DQFd5SzdCi4dob2sf
KpOs4GpOh9hsFW69N8htmwVrEPQiM5ckITthBC1HF314FdJd9MEUn2Q9graBj7OS
JxBj3SnInp3d8sRxabwAOXwHEAq/VAvtPeQfHk46kFtzo63INoHHx8D7iuDb9HCt
FQcDtBfybimRJ2h1fLIY0dVUyKbgDqoeH6GotAX9Cqaeol/ASwOzn4GZXqIq+aJq
sSKMv+NjKTkGxsamUFy7iOvdsUmHYc7sdE6WlrJ4Rtn2EMwVfFCs3EZAB/2x3Kkx
ZPUgcQlGnWjMUQ7DkPp80nuQ5GKdZDKQ03pcjg2H/zbeqDa7m442erKQVBCXhykS
uwq11XdP/v5F7PXsoYZwJpsxrlQ6Ycb5Be3JzH2Wor+JUIp/MyvJIs8U1+Z3uhOI
urn6djQ1BWroCSgqQjcmwWShl/umYMIIcGvu4ZuPcCZMgAuofevq0hw4asFkrfHp
wJv2JaCEXpzo/Qqld7NoeTuCpC6yvO4y0wZWAnBbZG3bYsZ9E79JSxxhviH5blsy
Na8KLnsM0BkSLHCqcf4kYK09AjgmKqXNC1WPH/Jw25oDHCz0Hjnv6uecfQaYJC7b
aCkZl/uJuZn7Ap4E8p0Z0zHVbkKiv0fzoxGZuXk5dEGdipXofVrUpPhUPc+93ksv
GadkIwNMapnRZAJR2zxeu+x2wEzNBoWuwgRwaAdc+sqHFVxHjBHvQuYMZp1YGUZN
Sy+LQ53QKnH+DQtYdccPb5GnSlur01IL2njzzPt3C1AcyuXmF7o2U1oOZLNaLGyo
Tb2AqdWZ0BxwXRMzbOh2cYjl77CbrYZv0DvczgLQi4J9lJIQm71DSaoM9kCx83Rn
7h4xO3ORFzD8osx3emMV/lHE/a2avHCUPK3yH0l/y0vQ+bQce0o8qle/FMUz0W1c
BD9Bax6MR+SrBVC9NtlrhmcHwTDW+v5tTVvP589IVQONQGU0GGjRoLLxMYGQ5j2/
cJciflcIyo6hKll39+GgvOa/wrDqqPi2NVRDD+C5RZI9YZ1Wrv8130LhmwkhLjB5
b77W0wXsIshjt8BFMJr4PyTdgYG/qrhlDhUQxqIljg401zCYoYGdnd26oNgBbOpI
+rNZwnGv6fXaM/Yr3+aNEmH+L1JCU6Fo5INJNZKXwifV3GZG4n26dfRzoifTZIRV
rVQIof9aVDhAcZqXlJSyu/KWp1L4APE+68CIUAExeEMIq31CHGTc244LWbbr1QWE
gT1itqUOCIU67USI6k5RYjulFViG7DjR1nKzeSngMaxTIeDgjLtMoxoPdX1WpXm1
s21AqKmJEiKhQnFdDkJ6PSrhw07zhFZ3KcWhI9sHJaoKSUmvQJRFqe0YZwUDLnzf
d8USpQmz/2B6oBxDWkzFUuqsryqfH7HSZv9RvYuoElZCg1Vt7xZbFA8VuuJOvrgt
H0Yks+niFJlDK/c1uPIG94QsyTJJwsky4pidKkXIvAOlZyx1pGNkZNoT8yskZb1B
oejVB/TjRV/wRg+Rw+ZHaevU9UQKReKsKC0/gX3ulmdPbkLGxHZOAOjhri3ltRvS
to9ZSGE5XJAb7qoFex7WtKm9eJ3GeZdeoXU44JSInoBdKZI2KeRbqv2yDJmF13/x
gY1Gh96UrSc3wvjZmucgyMartsFWorSyISh8qdbr5xu0kJmoU6yq8h+TsmWCfF9s
1TKhT4RDLe/R9tiskwo9kBGz0tzH8qc4OXurgqQDmqUIraM6hLyAQHyc9ui8p/tt
SRAtOayOIUQCDjseYUrTSLTJt58agiefEK2JPoK+5t46VXBYw+VJXz3D3torPI+u
6G5pix31Qnph4zsxCFo+8bqGtsyER+I3vVLr/l1MDAyatwjk1yitBBcngp1NqpN2
oXGIIX19mKO0OLE6d7b9g2bvYWiCPoocN36oVn/GFuJzDbYG3tIZ5qv8Lcw1+FLA
ixRvqe4AmckeO2lbghVPdItc9B5DEeNA4z1mfsEYTM92TKJHPQ4Ezly3TcrHs0OX
JRixLGyJ4vIM76WoT8Yg8iyHtz+/C3WQnGC9yAUkw8buKg4eWlWIu4ncyMbSm3WN
LFaC2K60D056bxoa30I96uE6E/MI/UVAiVWhXYREtPc+YtdzAfm91KNYaVNwWIBS
KnASQSYPWbx6mnAGJL40wEU4JZSHjtBikB4+D5oFDEX8g3DXdfQ+tS1qLBSDUTNn
lvLCrDprPRCOo9mMXVmjzQ/nYqO50bfEfZWPqVGLG+QVv1zEsFbQvUmgdgejFL3D
EnVQ5bfZVl9OiA57zESE0jM+sCVrxpQWztVUz0XrpQTN1QyB2vIP1zFJrp41+NSQ
tLRfwVXqlZfxzRgwUD78x73N2RPGRXtjQfshfQP4nmdlstvysnQgSjgPBjf6GZph
XVU1yo8axCqSznwElVF5mp9zzuBB1Y4UQLVh9hj3DbBc/jRVMJN3Fa+Uc1Ykwh2A
S94rVhdz9uhI2sUNKIQlLWAyyVO/6gFwWT9Gg2dPgQa7F/c6btySCrD7PD6LY44j
GbLqDNF/YKejQijgc+iK/CMX826nAD7d0wE7E75FwG/5TIAgv80PfFDu+Lw/yAV/
yAR8JnXM8+PnLGdO0g9hwgJcPojWEQs5pWDxqNCoDfbVhomcQONxPy2rq1URVXQx
H8zjWvkTqiZLYzbp3PA4uucqNqVZiNSTwIaqLJ/YvORWbwNVpt04rA3cmues8nq3
3AqHvRd4tokwKmfQdN3OkKb+ONuiI/JShAU9OGp7EGk8uRYkLoK8jnst+t7bs24C
25MyqKBTRUfZyn9e1xLOWFI2IQRtppFApSFQCzfkQqB6DiHOn9+Io/v+db8iBgZw
d9eQFoVZ9FfjxphnYrIz/LePByVlQ1fVb+1dzwlSDGMsMQ6HfKexKFNKVkO5gCAS
VbS+yETAgPSpfwzmhNEFduvyOZZa3jnYfF7jgCgDAiKnhxvbMOcHmuqyb5MHSgae
s4qEf/VIdICAcamHkzyzAhU3kdtl0i6r/2ADhIkifN2h7kkvwTkCAETDFonWz/wW
GXDLs342BFPkqUYAKhwzyp2qy2q4IiDDUXteoJzf/IW8/xvMa9AWlJgyCYyZn1kO
jvyJv7/kEzszg0YjPUMRSzqGF7cs0wU/sw8KgsxTbaalJ7Wn9nrmJqjLOCSqhTGn
qgA54kopKgKnSdlgaV8AJaHLb2guafxaNm2OM5ZfqLCnJuo0rS/tKlN3UpNadKJ7
q1D1IZMqfn3C4aKf3w2aKDVU9wVvc7jQ2j4CGfYIkhnHgAlFQYmGQILTlsMfp58o
xeS821taInoQF8/TvNhczF2mF3ULBA+Eh5rXEmsdWC83vFi0omA/dCrEvJuBvtCV
m0e4/W9L7Fi6ufBo2zksNuA7bkyWndWOwOusutAQC+6/i4KK3OLNTQ3vvWJnx79q
hLYK3ia5MRLrPJ5DGQv2tCPDFVfFRDAdJOAcSD29EcvB4y6lBIxjNv7U7C6Vq+Sh
MP3aqGqeUt+q4zSpOVvsPCORWmAOT8dq4YHdhgsRPFzHCNFH1eMgb019M7TM7Etu
PylRZAyc7lR56UmInJuOrQsiKaQg7LE0GhEYrvZYPl9BESFhADBRDAVFW5jR5mkP
DAIGTRQ1fgAs0pLKole90V/Wi3WAWgGwUSqC7YvG1pMWReANe9sjSB0HioyQedc8
srXHlVx52yLFooZ8PGPwIvvbwMYso18ssfsuGNll6B47sy9z0Os2AobNZLrKHmwI
DqxtKYxV8a29783POe8DSgHeRWE3S9+47AEaT2CqnH9Y8+39YoqzI5haaPhWtqBG
cXOmisoF5xVu86sJSobs6x4eaXjQOwA29w1HHDR+GjSyfpkyxJSFBzhkfBYGGDwK
Xj8wlbG0HPZxflFEVtqqx17CASAfJw9UIpeCM0yDtPHY3YUCBoj8SOh64vD+E8h2
HfZ1EM5yixwSMMITxE+B7bQs/LcuX75vGJd8EOqv6jdIiZ0Ggo5+7L/dg/thmyos
QKc5Fb7GM6XftHZBQoP3FW6ZGPVD2C16y+NZzsNSEiJgweCLvB6N51LeCKT3bhn9
HtEeOGksurFpbYUN8SiyDkj+Lzzif5DcdFVWjLSfAD9M/6GngfucJJ9aiyDf8wcZ
/VQIh+lzdp/diizfgrn2HYdm6VCFq/O5FfhiPbZp7DGmNCPHVh7wYmQnzjWTsa1S
FXRpQ5yQUKwXQ2L2c2JNlx/ZvZAUPqKjycUnQmNuom6GY88h5KafZtg6xUQE564K
WBxOV59yC4NdihlWchfyPfUnC2o8gaB6uAk/sLUOqQROKVu6vyF8bWSyMhZ5ygNe
0mK0YVpg2+5PuHNgor8w6GTTtJ4GnSE0h6OUyxgjaf/1WP2avZu6b3PAtvvC7GmT
mdbyqNb/Xazvtnr41Tg+cP2ke9CBFst3YO/Bdx3dkRWUoU2fNRbKzST9m1V5Jc2m
yKjjHDAhTCvw/+oLwJcHmz2nXA+uxJoSVBe+JB6qVG0A5cML+sQNs7KS0g59fjTi
cdwz9PqOhvhRZJ3Ob3lenX2bj7PrsndKqRKyxDJQOscnn5UbS23J7/YUT5q2kMU6
3WJG390TdKjpQwkyV9liqLTHJZ/J1v6WakTLxSwlVIUKegruWcoDMeuC5sxEanFm
w96SYmeYjRJIbJreSjCHMmlgJgYqGpPUhydgxiAtA+hUtDFhqGWynP6+pcnzKzDI
rJI/9q5C8uuGG6CsV0bRQFWUbQjXCkyQEx14mngSPzgPgE1zmIjnrgPjyx0K/gxZ
C8B/WylDi3ViMHw7+KH6pbQVQXEoodAgNc+6TQRyLrBCciyQ6iPKEHbl+xjarD10
kXpk/AUfFabmgPythQM3d/2eUq+jEZFsy1+y5Pvd2srA257oXtSrxMP1zN/UvWYr
9CS51zmVFCm2I7nkybcgBlGB2WzNF7vaeLy0DCt7EzRyBVJBFHB02ClG4APztmrj
61Csw6Ei+1akDplpsl7ct7otETs6dFzcrFimtBe8oh4ideiUZFLlWmxjJGE7oTkX
eOrg8+YDPs2PTrmQr8a2RqxfQisNiuAA4TNWneKQ992iSLrJiyw/RCFvV2eZBGej
r1BM6w1lxmR+/IJXfLg4JEtYkqRohpKJHlgvu9cgE4AIPF+C6/0Y2y8s5Fykv2E/
WPgcxh4KnYX5tkfcM6Pr1FhadBM4orrNLGIQ/0q+BszB/zjmyQQ4crrE0EJaXq0K
xZbM5CHewVU/m0otde2Jp9koZLtPWHsVNOLb1M/ID+08pZxt38+ANoLnXtr5djA4
u9vYgjkyPdkqWYrUl6K7hihc83gEPmhXZ6tRjyWbhlXY+h6JBMqUwq8mUdIZM36A
Ry3r8ESaCzsmeDQWLeFbnX6Wv2TNEYiopdCZxZeizxu1ZFXf9fG7Fu77rP/6rKwL
7M++XuIlHwIKP4WysGEXkvYV8+g6jJ2y4lxIBpMC23NaO5ZYRLUZ7t/sWMYqU1Dk
ajeP2ifJHGXNSIfBrbXvi76LvWlE5FIcD4r0MrD4XpNUh7/hiKJufiMQYeP6MMKa
ah5sQe1WYdLFM0RHjX+CG2HHwl1bgRXT0iYdxfKAYXaIg4PV5WBYRnYKz9WY5Wew
hejS2lhwLcL6x+KPoJGyE0DX8uoxStalLEOTPtv3VSSKEbS6aaXzmDlyehJ4s4T1
pxx3Lyn8dVyDYLsitvSeLkKDqapdjNXI0RTTpQEreFPOTO7f2JjBjjFHVqA2QCMG
WALiFnKfTvyU7c5TAOmNmEpGwnlFE6xDG+UWkE9TK2flilirigdbBemh/M8d+Swl
t2plsMMdzWTEsZbd0GvAFXkiXdmGEvAftngIa0p5Xh/b6oSDmbmgFEqNWBtBzZlw
od2almLZjrF4/4qw4XZXU7yVrNZrmA7PzYioZJgNSeKT7vFRNGowsiL7iX1XJJdq
8uV/Q8406wh9f4ur3c240voBxlge3Wu2bgw4Dfg7SX4EAeFxmsA4uxwI5AaMYt6l
ZsDxh/dW7V4CQICsy4zjKkq+z1V+ljRu1D99ED9CdupEFLH+Fdonynw2wgMB7oFh
+8NgQrl4GWhVOB3KSm73GUW2yA9FJ2LoKpgeKKZqwSkloGx2IOApd5ld8pKLpq5x
alYC7HAQ/Z6WH3lWyD0iOXFfQee4xL+vKYof/X0Tu8y04ajIcDhzxgS18L7DWIeZ
dphJkl8eUPUkcVShkqgA3poep9NYmpA03iepDHOHyWVSJK73d8hOl75Dv5A24+3k
L0dWWMOxZ4idkO898wY9DUGQtQlg+bW38HrrUjTsZhXRw4J99vyCdPRuyoFGBagK
zGMn+367NvPmKZJTDIpdyFlhNO8WofwTbst9U9zABHlASnQxE1nHZPXjaLLMJOov
oOKW5KszL3wcA30Tst1qKoCJodCSiP2cFArZS1JQ2OiTF5LkCJUeuUe779JEP9p0
U4Fg9yP7V1AUDmnj9aERO7aNdv0l00YhGKESLI/y++eKb3NBZWbZLaBa+Wjolutg
eiBXDPJcGZalJcZTSnWNrQDWHCto/UKRvY8IQkuN7UWttE899IdYLByAQbJzuAU7
vmAHxfTRdwm/bULJW3Hdf2Xw1luIZ8TKPvYAju2nRwWp/vZdUdUO41c8fkiBFSjT
ChdY5qJD8zq0R8isktLLUGJyaM4Fnb7NmRn4+V9/+NVaNpSp9Wk/jv0afdPYGoHD
k0RM154HaEkXhyxXSlTVwTYjmkB7kPWnf4DIfedVsE0zhZn9yo5eAQeTERE+Bo0Y
EaMpxgTuOJl992agfYDLRRll+5a7h/F/qBTLJRwxIb1NBZ1du8Db+Hy7BsVukpMv
CFJ4eBEJBYTSoYtQ5gZ81RmzfVeUW/e/Y5LDmOwVLiYmePB2/eYc/9HkC4NA9XbD
nuxroVBjMGk+sQbaoy2DRLAcGjjMM8HiMsGviQPjTj/MwJWBUnjYQlZE6vxI8l60
Eyhx5TXJnmMvX7VchLAK/Q7k1oBvlzmEqjT7beFKoA9DTaDII1QdtDeulZU22M33
mErLKQhMT0rovnflo4T1fJWIOZpwU6xqmufsKzl/tJg9k2G2cDxe48JICkAGqpWO
WuEZlnBVzTTrNVJCiaV5B0f7LOWd27vmLepyp4/52Twg2XrtnLp1bl/7hlymYSky
y4fvXMJWQKTXPQ+XPzDGmf8sjKIisek08jhrgbIoyXoXHN6koGuuKOL7LP9xUNNh
ElWK47aPOH8sYSU8vIo21PuYYS3b5S8FPpFrNVIdx4CbRgKWANzgd+y5aXuiY2+0
UQWs0V14a5xkTCm9Xfr3kfmrEWEZ89HlETx/yL1Ua+jkMTuf5Ra0ZazZl1fb5ep8
lXFbjAXyfkyafiJFt1bpgQ/G+YtPkOLcqCsaN3LLqPgDo7vlhmqjaJ5TdkbxEfCS
UJoxOfOpgkIvA5NwDFiIaHkwZSO1wtfe6TkV9cJq8Zvj02yO00AFNlccE1u5rqVT
UkxIyjTvjEYEDXjM3bKhIapwFUr6SXvV2yXAZPA02eM0KMypFPR0QNEC1Fjs6KIx
Q76Adhr4uvwN9RBN++MuZbTAB0hfHfDFr25pDeSXSqVUs3LS451UN9Dxs1JTRZIY
zwl1PK+z26P9uzY8PezDldMMAngIF2GykN9/S3VpfsTvQBIujTlnDQaN0yRlwhC1
KwAdxGD5BEOvg/W7IdYa8/JazYdf/Baj5XYo1GzcXmoUodpn7D5+Cqwy0HnSa60s
VL2CCrOakY/fwr805gSvQpYJIBoGuzG+ErsvQqHFa1K7wJBvWPiDgXgkVrj6Ag0e
NBAWBNl0pMYePDVXh4zTQufK7wEKw9JveO9+b5U2KTnLfnDAZ7CT3RonSQpT2MQy
yvcRAiEuWtppHS5cUxUVE7QOHLQOWHsOggmZ8FIde6O+IxEiuSassUnN2PoU86Jf
1EbnRrGpFZ55/OEAA600r8XtA7aa5JQlbY+rZLC4VLC9puLuvAhRZG3WHStceAmO
ZqCfDDG53cJCXLpPnKO/PVoAklZytPGC7f6tQxEEthgOzdmfGfWiy2IrJueXn3er
quxxnf7JY24Qf6bxp8r1EkEo/NSaKFNIeYWFHTNUCnoIQJIJU6g0lrWINFHm+M4s
Qogk9UXjfrYvA4Quxl+ug05po++qyiXPbvheJD0iKx836WLPB6nVAXQcj8WSR9OS
dFwS49+Rxtecp4JKX70ozZA80kg2RLEWOIHpsqVmiREfbMy5uQkf7XeCkO4jtVIi
bteFpBmTZvRi+G8ZvCxuauZJFa6pU087cMLhAMBE9YSsi8ULMzF+s1SQjWf1xPtY
97BS4ZF8qS1h+RiqQTYUigVN+FXRXLBDJynIeb5VnRSSXRq8PZzMtEm+Ivgkeq2/
+lqFXweohNAaIKjEOGHA9yAOvb0o4U+AGAM7ZvQlOrLKeAo7BAjWls1RvlX1XAbu
madXYWstHAiGGV9nsuu/lxMjjfi2o6ZwbbY1aEcel4Vid4upAJPCiFCaDq3btCfU
Z9UmNWfyANT3gSXeWXHbRm92Nj1KEDR3w2tVrHMth4Zx4Zji2upO7MQJs00+Uigx
PJcP107aSDHC9LEWMUPzMrDIjievl5Ow2Eks7K4mK7prkoCpWs98y46C1V9KaPcP
SGsznI9k+NHbThTsy7fTIuI/VsmQVBjUc/oyuAyMOeBzzfxIoMeYodOhi6EBuYTn
Dd62WQ+A5g5RZC4xK1j1L91mR2d1QETX1Dr2luVWcvxz/LGiVNyzH04fCTbmvyaV
I3HXA0vVb4h0+XYFcJRpFucOI3nkHKPpyMl0GDX3N0XTIqlfbzRGorIR/x7Zu41D
9jlaWK2X0UkRGw24O7rzzspbQyEnRflQaGccXDjLSssEfID3dUMZiAxc11oZqauo
v38BxfX1qEEoCgM9vHuemfP1xOkuqC1h+84wDnKBnULAuNbq2S4+hqZM7kom7zXs
RIZV3QX3t66BaWnyQ6yqY13hQmOntn7DDgNmE2wjEgff+GuNMKZWg2xvyVxenJ55
CYOEZbuHmsJMA0VVT1+MQuNmc7jhkmGGkCeQ/Ym7atcOdG8DgDj5sfrltnGkl4EB
Z5lFXu3VzWMtaSrqVLZhOdvc+GgaI9Ab9o2ik9j5dsMHrrRCNcXxvzMTZawgxIqw
q21q4+rD/wxPueO4dP6b+h8+ESCHBJZMPiqWYm2ftkMx2MyrGDTRZRvdG6I2MboB
SmiAlygMl/p1WLbu/3dnbT7QO21ov5AfSuNU6xlpSIzqLGxKcAqk+oPmBr580k3h
Vk0LVeufhknC9xOmsVxCix2jsp+27SsuGPcHSUx2Z/UtfQmUwwhWLKedX5JCfN8Q
dUkWT13KQMzCdLg0Ve2jGmfRtlMwkLOWtJUsKe180azsSS/N5hj6CDDNffrjXd6o
vWFwnwAYlubnIOJWW9VWR4c5+uV9Pv31En2e2HfpLv+Y/PCOSLv8jWvdhlmMW+nk
+24orE06wE5dmO+ZH/rUXZ8MiVEz+DbuO5bzout/xVnAUtqrIGjRa/4oB3IMzsHM
k4ylioj07Y0+hgxxhYCOSKOKgAGTLGAA0YNuwDQrCnz90/35We2+3jP9rm6qsVjr
FZa5GN3QxBuOo5l83BxKpku5K9ay3LsnGJs1f27OpZYOJ0rIUEUJHXPGIavpy9C4
XX1eA5cnt3JyEUN0+4SCXJN1PrRTEsIaieoKOfO0uT9eZS08WuOu/ZVWsWwN8og0
rFlYob4FPhKFQt84azEZQGa/LeAc8l1mHa6oqDDzfDcxTVCjOUEz9MUeWxM4f0XP
CUqF53vYrwTrPZeLNCY4MSEKoFDLa3UmJKtCKXcWmrb5Oex5gKAX4XXMsqvQjC74
XwyCe05sKwMCv6wn+1BivLsZF6Zzcb1YCnYSIVYzlOBOx+7yCiuKcvm7Nh2jrT24
/nMLImYd5OzrMDR3Cidh6cc9rS79Q3iez6yBm9V0WNr0vDlMYRYutZdpxfdBP1nC
ydGpM4dCt+LgXE77JA3D4Csp9gh1tt3uID9MBzTqaUqlM7rLpLKacCDXpP/QnQ/X
RnXgEvgIh+CC6Ufv3yvIau9uEWHL+C0tpw0JURo6RcFiVaeKmbp+L3SYzwMi64LJ
OKb95TMpNVYN+5M/XMh6fkaQFYGiSIyhQ/Gtg/YKjVhbCvlZ+tUFme210WGKSkIX
3GDjceVRyFKVimzRUbxAYex1N5C7l6xn/AkoN5RLYz6yyQ+epZAUkFtNrCoAjCmj
waQ1c4hi8ANLDCS34wQgPXb55n0ZwmU1ZMYhAeHvye9zObo4KnesEuju32dtWRZ+
w5DBbstdLrMT3z/ck3lrv/IDgZt0+ueO1nxjp0g0rRRacQvTIOuDQ0z8Q2mrK90e
Vy7fZx9IPe8VwmyRiGmehsEvcYBKPttUqaEImiBOIKlG7ujA/fmxVzmnFVu2yxBp
MvB+kXM0TSm4XZVySkUnN99FbrRruhccPgZcFPBbRDiltLbqtfFu7cR5UB/4f0nS
nWocxyMfhx36bvafd6ESZLXZuddrInl4znwagWTbJenZyuYaqJX/3Y2QtQ9//lRj
G1fxWC6OLcf0Y1o1NoD4JeSbJmk3QAmG4gtIHNaIghqhwNPq9q7PQXYUO2PDRrKQ
Mer/C9hutkBOuUuEJnWfekf4M291lboT5pHi37Z2zROtiLPLFKQ15xAaUqdbnhd9
sUrNpKS10aPadHLuhDNJqj3iNDEZ1hK1PWaD4MUaIjO6mp2banMubQ6YLhfnxkHS
wGNoutnhSDjL6ckC9CqKOld1WKrKujUBabwvgBDOWa8wCScOjxeGjueMkZcFAsuT
QmDAZf8YjmutejYfrs3zPqGmZKtOhuUyXu/+JahiSRr3COgsdWVRSymrtrYWa68o
leG5COls56hc/6o0BAxJsacsjaO+/xA3fzlq4f2q8UuK8O+H9iFB4cdTuekkpUuh
Neaqc+i1mrPQxLpCl6lQMoIxgQAMNe+IHRe5p496MXqFCnS3zbmOxuLR24BE3kc9
qkh30v5sc7K3QSp4JdVBj8HWzTSSBXCLlNdRlBijFYm0VRQuVUsnR7wMi0jx8VIY
wTkUHcaaBFjOmXaTc14l5Kd3BAqMKMZ1pGQ1iK0sSDDGZfQChQZn7Wx7TJrcF11S
nkcJ+XNIBRtGc6tkkH2h1jstKr/zTQ6ESQ07DD9Wspq6tEyZlVwPm7qsALHHiXoo
tJYTxaBzn6tcbuj8DBgHdI/GR02fvn9Y0qbeI++J3Dj8oRccG0Appw6oXin6AADL
Aw6LpuGpr8+1UXkHcs2W/lmwYQlKw1kXaG0AXfYyGehVjEcGStDBsnkyqWYj1lDY
SKSrrCnh1KvdVb5IlERpxDgXiU6EsyWmhHt3+7w3r6B48ntLNQD3tqvnZtPseJNr
M8FM45bQqcSYjkjQFGOnBYjGsWaYAdgwGay3NIoYagcuL9LMy/puo/YXyTn3no7q
hC1ZaQcgnWzUCpsUu1dcOlVTjfcWUaqyXq2TwnsVVdflLFJ58HmtJBAfgyhJOerX
n1aFAS43qDd4YBqCgxugWiNTELOQaFvZrKBFprvQnlgh4R7jqDX2zXXQ1xnc701h
ujFlE3N4iKffIEAfseDmI0pJznO2UOAq3kp5lYL8Hg/chXJnPJRL2G5+pvWbDltE
g8RDLGYkBaGMkAY0vtUkI3MifjGAtwSKX0ybenSttElLjlV+YDGpGZ3iGhq8ePkv
ZMLb1Eoxa7ASCifbZA5RNR/1jh8LMxsfjCf3Ia1NU1e4U+Wxqta/tGqK0VCW3E2J
olKfAluM44IgTkKC4RfjPL5UggIl8XAxE8ef04RVA+4zXt0gFp3Ebrhh5QQp+ExO
k+l7uN3MH8sVwzyNiG11YK4TsnXaH15eOKKgIMLlS/s1h94pahgbtA6k1JOyRoqQ
BTIU+JiIQZWkzOKoFAbBWpdDyMfnOYXuft5kZ8h1dVZKI4/u8e3dksXxMz0m7BZ8
hrc5JeDhQz1cNQ7+sZ4P+z5DyOQHfPE+fNG/xA8PhqKvXFLqtznvY6IR+e4Mzt6s
Ya02a+QDGwFF+wOTZcSulKXcTaq0rC4ozmr6W2qKVnXJWvsONnJ9LzEU92mAqRzH
rsI0/9c3RD4crEpmRYqObCp8+NH81pjwOEn9HrUGSviW4VkONi0XX14ZVt/xoMhm
14hEspl38fBlvXkHLjKXCpnFvekHuVvNJqfCzEYtSoBF0vnoHM9nsPeUZG4USRSD
frGk51Qw6zu51lF8nYVqmU1jlrIX5ryavNwsW/qyLmF8LTXFCGoE1+OUFrOrtT30
p+s+exCS1Z6fx4RmE4Wbc6Qz3xQZNMKrJXm+57W7nFM8/YltIMrr81ydV115VIpF
ZyOusPerLB3Ky29SYRwEY+Ax1XVcUK5/pJ1WCnOoJSFa3qCvAiHCFU1HRNtyHdSv
WugJ3Za5ivFVfcIwgVs1dQTcu8ToYQkctYqWFNBPVTMPYFeBA1YSHx4BV4CaANjD
7qENS/TdVv4M6Mti/5EMlTOTOgBH2t0XvjdeA86bf2nB14lgZy6I5OYoYm1I00ZW
mB3/plzbu97XnWu/8tFGYrAK6sQzSUAW+SN9m4CW3sa5jkTLY4ZivijGftwqsP0x
0AxBreKK0TEWWzbUQGQiAXQvMCZfqIpGzJX/IY4RwK5RBCrh6EMs2JiACVOE3e7V
Z4ROgFXdwauhThN5Y293IzSjpaUrAvCf8791f4Hxk4+Qdy1fvBemqpAmt5mh2Qxb
tL4ZWndpOvp7qV7F9T5ON7yljZmB4xa6KTH2YQwsEjfkyTfR4PW4e6KQropr0B6E
0GrBymrp/2e+wIsSHDaquOqw69tdJ26RbpsJmbikY3t3dPcYJP69KgmY4p4j9DAF
9df1t8XM5le+8JkL8fwz3jQ5nMNCSxPH4l50QqdwRaYDGGFRhIz6WYqdBCeskHc9
zXvcbrkze6W005dNTH509vFljRn913eoz0EcqWnDOrXnvvqIiBbhmr0WgLrnitiw
zOBog2bhXjvz7SsIZakHnBZLu5EOLE2fmnp/q0O3oFBJSy6TQ0p4yRB6FeDuBp6j
tZlkVAKwlUxfJrTrGmdJ1pVYvVEBrBQHXSV3Mdx/uXo+y3gVTpAhS8xIg6nRCz1i
TXX7EpXQxX5ep3WxW1GuWvNklNRPAf9aRYn5l6O6HOBLDXO/FxAQW1KAgGm+5JGi
nZstFJshaMM69RmOtIkeIn/eao77/58kgf/yNBrSQQ2G/YDwHkenctILOSTl2cRN
tbsCgWRlLNtBEDTT7emf0jE1qNuFydkiC9rPOjwbSYbiVXmwbnDowELsJS4SHQIS
9fg4hP+/iDa2E3FjSLLUX19DXFSmgIt3CXpg0n64tPuArmy8r8apsY3nxV5GRyBu
b/fYOMoIDlHepskASRDd2YjAcGBxJqLd+TKEbJCPXHxYjUMebq52XUjPg4pKo7eS
r9u/s7jAqFJRN5X7Y0RCGPbFRxj7mj/60hIG2v+rhS557ZAbxuetSGEWTz+zYrde
FlUpCRlVprMPNJMYUvEJHpXsejTSfDHbGbLYIV6Muk8WL94I+fEyG1MUZ994GqSk
/yF2c6K5If4Zl141h3gVobXq4FI0VoqaZhxxQOueG04s+p+y2MSFd9S8AKwqqZbw
wv/s8IAijeZkBKYavsIE0IGRd22WMZjKeu2kPk19AatczVW1uMVfFh/cH+/THhrQ
k1xaWH7T9sLmgg1hIxI88/3aZ1+Rew8I8uwUFf/3grmR4VrH06jVHr1CwZCAFOHX
ingu/iBOIZgbUgZZaTsFcXTy0LuZCDMq856JHIERb4QOZY6araJsTowP5zDF9PfO
0wJsh6Iw6MbPVurVnPmfRJHl79CinXKMwQ/GAtivdMlpBgYKSCeN/hjp6W9yPZMU
OHwTlOdu1qNlPH3ozf2V4q5SezXbIaFNm0i6ckMSLKgRATruG8dLkaLNaKp9SE1j
HY0t/cK2MznF9TRPtef88iz4JmOYgsd9b1wphw75ZyqjuhKoL37StKAahrZbVuFn
IfNXss5xp3yf6Swsn91sJk3IsRkx4tMZOzz70zBJMunem4x9wm+Iv90k1g7qlRJ0
MW+QVrtfwL5PzFYrYC0CMzJdlAkjvhVaGxXywxYYizxIod4dZwD6/yVXHdVg+MBg
pIFuS88OeHGNhgBoIiPMnP/qbeAzIPLQBhmlonFAy2Xmds7mETnTzVXzNTjPj6J3
1k2H7ts3nJWC1NUbvue67XzZ0WPcYkmua/tjB9y/UDEuNMvm3I1XQL7oKytQ+JTw
O29xwly37GaaBB2mq4lxdAlPbjFbTrbI4TdDjfSf0PM4F9DHw1q69XgUukuD8cw0
+c0rHNnzpPcY+tkI+3PPiCSpu6GAluUPYJOjaGK3PsthlyNA4A7sNM0n9NI9Ipbt
V8Fys4TpJ/aDphAhm3Yl8A/jFRpLpSmx1stEGnNuxEZoeKMf7OpMf6nYMW+5u0WK
ZtoROc+DCHCg5FLOzAajp7OXtThiqj89IIPNiHNrlgfizmLeOlPrNLHsP9as9ErO
Lot1mruN0vO6ApAdeXFmThuI1Oh5oirlowWLUiJjHu/Ds2RDA+wQZUgcBmRLCFJw
ijSTwbY1D1q9uMtUQnFu8gTs8ccCEG2vXS8Nk1SADcggg14Vr6gC5PCcyGRf0nTO
Fzq30MEbmfPYlGAWSxwTjIlZfbZ6zkCYNGRpDXWu1lD1UuUEd/6bBsBdO/PthJ+7
EysSxFHuvzbnMgggS3ETLGo1ivhvNhhpZq9eqhTvbNCYe1aQGsXSap1n0VEnyRlZ
k5A7q/GLqJsirtkwt9Cide7Yz7BwxrwpGchVNh2sXMsRRjm1JAsvyszDgvN0MWg2
QbMpqqtYjHcJ/yBZH0G81Zmda5XUO5gmerI6gdxo3l155MnXOEA2V1QJNKlj4AWO
gMnxn/OVRw2Wo22tZ/shqbJVoQy3LIWaqOuv3tOf4jmrOAmFuDeYeIvIi+icTQMm
xijiPF/nanRIHl8GWJTgMbAGei8xrbzuu2qUKEbMmjNGi//a8YJrcDNwjfdlEKVT
LHwLpuQGS7RI4XnPDJfWVKNvvvZPCrP1wdW/IXwqwFgEb0UAXosVrM5SQJsgnsGt
LjdOJxoVQe/0emGIz9sdJWYug85brbSxVYHuXbJWgMi957vmzpKE0bJv6xx7Dur0
k/cwMV4jQz7bhpHDePO44O39BJqsTvxxKgJPwjp2J79KgfA5ohwIUyfbwoH8/Oud
gwR4Cr0fCHTMQChdc2cd6LhJ9CchC2hwzPkOpani++c0JC3JygCPvDIp12wLFyO5
zbcbhAh40mO+WDQhtdWJxKDA9+HEFBxonw1EyZBY1aiTqCVVOJYMNt7ajOMmuvUm
qzjPyawlFtAuN9oNYNPYBjNcjPHq9zWVvZkpWd2Evt4tbyBan0/NzEE70Hn4JdJb
4zJ1THaBkDO+CSlpFEg0WrqppSAS77hYY9CYW7HCv7UM7Umj4n8pyvAaOnPATriw
FypOMMAMR3r7F+ck192BKzS/cTCc8NWTjfkrFgsVI4W7dPxX1JN1nQ9uc6HGYCb+
qyjfig69QvOvOObA3ZE7N2w1bNLY7uAQ+eUED5TPA69LoBg0NX9ACGbvcjIF290G
nnMI8QoT1NGkeJE1BJFhGBEjN8Hc5rBQM7qUlm+iu2dOMlLxwMEg6e80BEccLTjf
jMYOuR/edTyrRA64utAReYDeTrJhSSabYtY1jJn3+8uXvMD7qA0hVXjvlpCJDklI
46jiCg3GLcswNqTdemDiy2SAPAlouTNzcH113rvUWtV+9XlxERcyv1NhL6af2A/g
MR62IKmPOAXl9HkTm5sVtWmy2wYxbh1/zO4BG0RgBuv5N8LXU5OefdLSagSuNERE
Un8myfS/VMV3tduhk8uNGTR6Kdenj51nTzOAf+mPWvVDMbyoUIApmV3awV7G+33v
RnwSiISM8Xog2XwCcsZ/Sol9wuLXRYfLuNuh28pVDKEqWILEUWUlTC8i9opgEwGb
i03uVFtklC/bcH33/Uo1LaYWxvGpzxsfrUFvAJcWpi09YaAhs+u3tZbPTvl+DQoS
CvRomt93CL/G42kerHV3UQ8s5xquIHtIlKWyesSx1sZLLvNq18L3yf1/hNxoiLkc
aCPDltPrXovRJNavf1/5ZsRwEGhbtTBNGkP0YjLbN82O53TVfDx6PQ+bJDE0T2Bw
bXX3koWEwkKbgve2i3w9e4O4kBSE8s0mDvduvq5jBVswjdkmbE+Sb/dItICFhc63
tYaW8gUTLQtrLWrBQvkSKKZnnQDJmhvViZSktozHF32Dyt/7EtA18rYwmscLAzV6
rpUl2qMTx6fV88P1RMrf/kLhPv279V/rwesRU2O+KGT2ajLJqkON1xzz8MReOmoW
iCTNrSArU5HciT4zkLHhP8CaEWky4UNVfoDnwUNpcuKTRixkfZJL8KCobhT5mnCj
Tv9rQv9uT6YBqTRsXRP+I/iNWXBwKeQPDBGFk/uwYj0xomAJrp3OJf2xeDF5b10g
QKjOkZha5fY6hhximxqKg3JFnBHWrlZLWHSoNm2967d9tSmWz1HhQAUdJVdAFqJi
FwqcDZdh6j2enATUbsfl7M2+I2zXjJGlXwzhPvIvfM77sAxwLn/L9nClbgOZdh53
O1oNcpAT2ugkrvb1MTtDw18w47pC9OQWqOSCAFHxPn7uDxr6f/KTD3TiWG3LKB7A
km6kDWXZ7UGc0JY6TAIVoEkkPJnSuL/X42VvUE074B6faKKXe07AcUI/KZZrIIgd
sLg8irKf07c/0OK3edW6haoR+zwWiAESpxHwVfmlGJY6W30uC5JEy8r15KDvw5Ak
kNYSy230LlLfnca+dct3GXXlg28pGMlqtYY0zCq+vrDlvthDCHCi2hzxbQHEoMgp
Gl6E/Mc/rUxcwlxoJVY52NKPcQ1pFfdw7AP4z/KbdseRUW4fFkX47uac+BEF7A9x
kLfhqm6YtsaMFrHus++CgJedthyJZZjsZJZIeu7vhSIJLFWiHPQDpkDTD/tuXcIT
WFAO/YVRJIPlhOBu0ifxm5qgkF7jSmsCRXskhgqZVVtnuHMh4sAN9MBXHN4iXyoh
dTDI6wEWnKbKBhV7ggMWg3fkWKmhtIfCa6cPyXdDDrnQrechirY/w+fEtlUzymWt
F4BYp3OUjgBpMeg+tGdFvxuVV5Wqrq1muITYgo+RgMv+/oaPWIoh54z/vZ4rB9Wq
tphidQm/rUpddkanZqZ1bB8Sq7pNkY0AL/9DIK1p/zhXq451/6HZrm385O9oJWmV
PV6+Pfh2NJGwmmaaakKVAbRGSZXeVOEYkZ+6JdzswY1u2vkblMcs4nEwqWlF9ys5
KvAO06YeX4KEno1SexacMVliNvPxltB6UY7cCCy5bI8tZ/q0gAfG9mU+pfo8cbz7
rbBRBbYEmz0leFrtMiCMy+NOzKZnmEKswg956AhjzBK5B6OaA0yANduRt6ZaBHpO
nNU5g6G28/wOtqTm2IWcmMMjt8iJ/OxFCECVGpWJ1iepkx/KyuTfJoFWKNSXFCAA
ScQ6RQX/r/QUjEZZvMkwBLMAENAKqwcmfah9/VPeq5MPc71pgDGDn4BBMxcr9FwO
NaoZ4li6SDtu1KIbLgmeJeOz8btXda3vr2BB+ofIZNZwBAwy3+P1/pqZPZ1SGlVY
hTiR0ClMRlQtKRStU0PAGlTCorOE1DN4H2o/utrXsyLTbBWhM50x5i8sF6vGGovM
4pQNbYpcy+eG7MHKgDUZoWvvACrfOob8ZXpga5GtlV2YmCVUxqLaSoOVGNGT/mzA
+GrHxU7e4BqBa7fH4fBb+PCOcJjQAs26VE6EIMkGiloHBA+v7V5qiOl6tZqxS1k2
eaU+hox9Vu1RQG/dree+N0eao0sqGEQc8c+zJTf3XDVnoqsNortgfc0WKyeBwEcR
C+lWyXVYNWzRuIdmNcGhpVFOPsQpMpsVfcn3nRVhiFWL5Ci5dUNEumPkVSd76H9d
XQXV1YZuMcEvWdvyaZcH4AgOwaRynKbfN+ARQWrGUSztjm9obp7ImEagnBGYxMYp
cqccB9VxwD3YOmgUPXkwqu2MG847UeNuGCumEdWsIcUzc7LEvAGM+eV+WghQ9uP0
cy3GEZhcav/MxRIBnXvux4HYSrL8vepOy8BKHqgLa0I3KOhbdIGRyuu32EOj/mbx
MWB4WA6w0XMF2qan3CrgDm5TrgRAaI7KiOxfbPu4KrqSqkPdMvnIrwhMpTuk/L/G
jhfH5Gh/DxdsFrk8Cdm8fzjSREPkM/ok0STbxbyRQT4R+HNqE2d/uLWg2qafP/Bh
2dOqyIcTrwAQxxyuTKD2lrC2jSCzbiQE6IJ+EyaG0y1hDimjS3VxPh0USqcl4v2A
XqcCkJ3+icLKtK39X8Yy+EVmIwHWWCX+1VAQf7qh9bPwUz2JWzkHcCjY0suLg3NA
y5rsi7uMDZOiTalXT8UIvC+voJNI8V04O/gl8RLvdshzs7NzFLFNpv0rv/ZWt8HL
WvDgDvMAzMXZDDRtVdCO6nO2SR9bKRRKPLSKJ2II/ix4aLEjTdT8vcojqvqDlozJ
rh+G4u049eFuk4LWjXuIxu1qGnX0miqVNNKgMuCMxWMfzv1gabBUf+ED5AlhuRqI
AO8mYNFr0u/f3M//wOCDn9PnmoGQRhyrGuC73b79jQL9f3ug7SumUazW/HX+dVVM
sGoa42qteKyokiK6kEUR5I+2ZEvwZ7eZx3e4fpR1JBaFRxZzZHI8CT842aQIhKPr
TLd+oBuumKa7vZAIlF1XtHFiNQCxcxeCXpIaaDi8uiAvzH/IhWNJajP0pHyfzdiv
R+pRi5y6X9AL+Qln3ZQagiSB/elGdrYgf4VLWi1Me9/3IJYuKkhWXkdB3lNnVOtH
yqHfbpKykm6wUxNwtiN6/E6gzt9SvW0y3LXMpcG6qamLfkXAqPySJmJkxDsDsvjZ
JQlTQQGhLLu+ILLv0uNz7vFc+4Ktx6BYcGe2CJSHmZQt1iypx1HTMrD+P/UIrfkY
UkvwtibXusbgKbKwJ/Iy2R7C6Hv+bye7iqbsmY1uKo4qFn+3ICq+WlkPX7YsHxT3
2LtOsQFKfS8lbZizhOqL2ZoOymsiV8jW/MMN4k4u4oDS0avoqV5Wj4NBWOzprrQf
rQkVjspuGGB8F20zpkWCBEbFO2LWBf+v45zBNSGmA3XkGz6RZS96T24TasXG+z8u
6RhrUxbo7m2mUtGYo38DyxN5nKkeCVZUoekoaunQcPDjx1VBMYYfKYzUUgQ/nlVc
5ogZS0HiE9eJ4ftQPd5ghF3kVvA6wYVvzXD6UUThgPBsAzawwgPC1Go3AqLOIKxo
tj49+eaHgvLD2cUGnROoGK0jGX31SWPeZbfqyw9s8Ky+Yq+L0xfgFDHmtpG7mGT8
6BrweUJ3LqwHfDvAiiPtuTCjpkrGqhOSS0KhZ8s1bdwk66/VyGTQVDke2xpUpEpG
ZLKfRA2grbCMtdrPdSJDQIhNpgfQTAs2BdOLjngxw1PWhwfbThGGDl7vmLIX5Xy8
8rNAfWzgJXrjBECq3OgyUGw7HGck0zDED3KvKhscGokg6ZF7NMO3/ElVa/wLGXnI
jphQ4z6STuUbw4hPikYvzMpSW4DEU/x/hBZHI93IfPDgLkiL/LmjbWFuCTvpnMk0
Plg+FD30VsUd2MHVlZ6kfSimJisw9CKKZb5V3ZxUJ2OKJ352RSgkDKPXEd0xj1E2
8cOeSJpSXjxox70LcI26x2dGi3kK8YfSHFCRlsG+KkxmrlmO8J+CVfWP/oQLRBDQ
uuDzIWBbZA0tCY2Lw4gC/69IFAMMgTK56nRYoKZJ974yOUL1ZmC6v18t3B3+Y1MU
WWMrgAGc38a7cMz5uQqSX02XJ2nUOQZHcohR3osmVepCDN0uij58PHXAqkCE3BPy
CB9I9VBfJsrBZdB07lfRuSAFsmEB3+wCYtFhRHoxgtbu/rB68aUjWh9WI5dEdlIq
XQWo/1oErpgXpBljOBydPFrjRfDLH5qew2n50Ww1LFfcDZsS2QpF3+K/00oS0aB6
pCM0K0zeq5lrup58WkBW4todDGxzGSiQ++bG0u1m6szfeDpB9H3BRCLdAuO+XbDD
LEe5xO15z7gRW1PSdyZGm/9lOnJsiMNqn+8dcGX1GktbEZsKsmOeXWX4cHo2w1dy
LqlN6/ivPFfat0jCezEboIbpUEvZGgp/cpYJP0e6fLUwo9yXQpErCcownyJkuL/9
O+1krvXfaBNdjxdazxY6YiK/+uDgQJg4B9Lo5keMtfgI8259s/S0hb5+loEUGsyl
c83BO/gAt0Xs/Ini/3AWhoVdPKfJfjBlzAvxE/93ms5SB3afrK+yWPH2fSjaDRT6
kyUVdjWAu1TnnsvWrM2lY1cUoc/F7ufCaq7I97f/SrUl56roq3HmBVNo4Ps3I5ml
vLuF/SC5rq4TOcR6xUHdQWWLuluozUEX3IUIAigzlXDm8bx8xAspHf3J3DRS3e/l
LTI5tiRtCYof1knEqEfYvJBxF/t5E+awCymVA1ZOOEAO0E2rrUAjLq9PrfwilQA8
mlQym/oUoXPkP0ri78D00JBFsqy5hPgQSfzS1Ta44XVTMQcsp/bjG0nkt0dooogE
iDK19mq1Wu0E5VKj/ODQU2TQ8oqz+YdGz/vKdkTgEiGIKH9TuzO56nExWjOszaxI
oKBEJB7NX+37NHIaiUp+AEdRJVduu1f2YQDRP+zGINoRRdlRRp7fGTSBwr1yqD3x
8HBSowq4jpMe27OeZp7x6K42O1sF6bqh71Hb7lsCKO5X1NiRORrVkxGKTjlhwLIP
RJ9Yg66DuaLavJqipWOg8kod6hKlAgpusIlkv9kOjJmVOqmn39r6w+LMmqxI4fEv
/SjTaWELYpAHnEQ5FFU2FSgH4oD8+deDZs+7u3dCXq1SWbpUKuRzUC/2T1cCTlHQ
DoIbJcb45yksMCRdBOPwgZj8yt6DYCJ6wXqSwyUy7Lw1X8SNjq0bU3Hv5Ii1qZo2
Hq2CB7nyaBzb8KPTgrEL4ptARz7kNWTmqjK3qrWYfdBFARtePyuJWHWBPmLHkatg
mRbkxYH8tLCbM1g9TLtO4DJxD1uGbFFb5RbmMYMeEOD6KhDJmjX/C0EJLRdM8NF1
YcViARlkJduDixFfoV1E6uptmWSyYPQxIQzst2tvRTa1gQ6LWrl1oPCLFFKym0xM
Lxuhz0P2qhXNf5pcv+QuwfSYQ1QljtGW37EeP8lTWNYKlkWeXgHITrl5XJou2W1b
CCTmnHgGMy612V4J35HNG3bA7zLJB19wyw3c5uferVg1O5Zed2UYmnNMkQcsb3oB
/IKeJhsRigTzcBq7HTKM5WAOAKzOeUVEZiSoPp8MSAowOF2tn8lwkF46bZXG4tTe
bqd1rFahfjaCYG76IhZOdxi2BJ6LckAcom2At4ONR9iULcdkN4JVq8jXkjqavm0L
OYzUznT0IorJcBFtMvEh777N0+LlQeo2HMwD6VjywspYIqA75ve5dx+jfb2EZbSe
T+2lGFOuBLmeFYgxyluzRVUp8zXQB6Kb8MD1m5774TDQpTegiKAknE44GIxufRnS
uYXItnZqE+oxRdYsC224Whzed3j85e2qq1gtCSBgtGvEM8AVBKSpXwjqOGw0BmJY
TQWz4BmnECKpUgdWHOcVX54Kjp63aHuhcevLpmIZh02ElhB2x5aLaJtrA6MnJeBw
U3IwykeeczndDJuKz4IsT1wasYvHijosa6Kh+dkG6AKDtgevkoWioUN9KMWJSzZ5
vYCwAjKbJIUsDZUmCF8XB0pyrtDYeaYw0wEnFKlPtXBECaIn6BTykE3NT3aodpaR
ELPxoMltbtb3ggDFrnOem9lsUbgCI/sj0HZCYd0EZO16GPKF8kc0Ul4ZjiYdXriu
Rvw8mek4yiYdCrOPb624sguds+Fa7iXrYtGIziJEHZ2k5EDHfBCykUctMPi7qJ96
huK/gDhxLHP5VmOU1RZEVleNjYxtUTLur1v+xOI6QUksym0mTeu8mkkYBz1wjQav
TgskuYTXCGPzaswKOsLW2rsBdAIdsYLIVosmcDhfrVvCKMD/mDh6/BKQiuivywcn
fSxuaMDcthI5sjcceHMyfkLjgGQL9mnC/5DkIXit6STSDJan11g0YIrsOGlbM/AK
J0WVnx0hSm24z7DdIVM3t81yAGIm1QwMHNqO3luSPWOyQmZ8aA5E7jAEFSmcylph
bkUhraaqrZW/1IQNf2R1ONL4VQeLJpLIlk1l7HMOYAryXLZhpDXhGs7STfpDAeos
9gUrEZudyZouj96koC262/VQrjaEu2AoRSAoitUEhfpFgosSaG8xXyYypPJabG9N
VuZ0sLOl+qgPHdpYomlsuYaX2BHdBUvArbvtdFQe05WF3S9SHQ3HCx/StUCn+mBL
qb2eudnNVZ+bwA3YglghdmtFGW/M60pfJWS21khNQeaLiAAUClA9kn3CTCFEX6wB
KUpwgNNPlZYFEGhEuPUHK2hRgZgGGHUBjCM/hTQuO59ptth/PrTKwy35x57Jf8rd
8iGsV3Pm1N7Vz3FF7P5WfCEs3cpfMTujRFbfnkiFd+k8BVkIpT07etgyfSQKX/Nt
E14U3pe+0zP8T4SMv9lSC3nWUsm5MQ617gWZfnPqQDVf74U5HNi1UHEdOD1gRH4D
rt0fIZVdF3LhANaq5wmurg8IbaZd3skOWdHCy2QGrEaB8kPvCA/3mrS2s/IDUqrz
n8M+5EmiAXyQAUaDWXpLp0O+Qnej99ikQqvc401nWLlDv5BU0esKgGwdbOxKWHsW
5IyHHnWOnGOkcOSirozqwpTNf4W165wlj0MnScZhgyhWTYDjuvmRZ1cV1GCahtUD
tE83dQv4FYnAGEuiFi2eIZrhbH+eMR/KDv5hc5MX5eBvRfAU9z15sX8v/iie7c9J
JfD8YuWOyUHrxNxc2vuPNjInWmUNoak5ullCQHy5rTy93eVt041JVbHEgrqnRI2L
D/eTKewOSkFDAkF0X2vM3J/67rEQUWjdUOSvZI9HUyt/ChGrU2fY/JFIZyNV0EEq
La7/zItypBbAoXiaMGANqlk6GXZyhaQSN0gFWVOM8IllnLXEhX/NJDyX6oz5yFh5
6ZmCbn/XzM3+24uwqylyyI4r8ZSgGPclfrtllRSwzZ6+LxFw+aTc2A/eTjpYZyLy
HOXz3vsi9ZAvaz+i4H11rl91/NLAQPYZswNknABMI+6V+vrCi4B6YyFeIQXBoPUh
VLxs0N1OvaD0XtXG6tA+jByVODCO1jWIN4w/xZ7ww6DbZqP4Gb8RKwHnnPNb2wis
eVgqNSwn7a4/5U9EeJno8AGG01UdjAAg87lkGcNqZhYQNELhMaEmjkJ7GVle8JQe
TrwSLH4BvFnVQwzcCD7eF3dznAzc7A5nPEJJF/69vYBpVt3r7kzqJJgI1WbBVeAx
mwixDmfmxeUZkHIhBtkMTfMRhlnKh5EoPA6jQrS3dc6wJQxQ4kVoWaBXeOtfDAmK
4ExUy2Otzmwr5Zf3HAedDMeEHM/7dwshiFRS0kOKuX6GnCcleGzjsM3qdK/otF0/
v3yNNqOexekfAq70Emrew60hKp10Hxro+psPz+LQ6C8svxfJNnufC4Yrtey96ick
jz4ErhcJqb95mObObJISV77QIJY+HZsgCpJw2NjL/7u9jBQxuI+O/iO043s4S+O1
YzfypUQs5UN0t9QfwZsMGcUXK30/zmRbSWhCorlzjuJ8IcKXD55TcCdp/aU/3L6y
JyvubIkTzx02Xa1YECDyL11BanrA6JXZufOJQDZxeSnHF2tf3Y+pV4+ZN7bEOVhE
QL9lBWM+zMZ6mkrd5GM1QCe1ARFapL7i/gR/fvvua+KXjoLnYDl0Q2xgKsfEdMLS
NYcg9lFZliU2s/Ji2oQegJRhxures2t77Z6qp9e/pyQZvFznmtg6RMUF9bQP66cF
0862pE94IZ1+8ro1BLmw73Hyqi/dTJX0slNkYmR4ly3+Jla9WTkM4plr3YXy1Sfx
H0aqxlpHIngq0lRcQuNeAKcH8YGgJVhyECgyDe/vYif0HyNncWSH02H/RGgFZaeZ
NoUtDnD31vrPOVroe5KT5ZsYu+4rsUVeziZjU+drDYPOBtE3h+HVz0OH2oj6E0P4
PbWn/9UWVJ+LOgNT5AYv+RHmTYDSZYizhZ33v0Deh83XLCRO9w2mWff5g13QMk6o
4//xF5f/ijQDDZDA6UV6LUaeo7PlTj4QNReS9KFw+xXbq3k16GS6O/lTYlIz7kdT
h32pRnxMxeoYuh/uPh4fpNlBJGKk9Ifpn5OIy+4TD51MHft6bS185oc/AAhh8KpO
zSXXstIjFIUTqEKeWgICynDqwAfEWhWB2Cbi5lMDYzlD/oq3vFuRgYrAMOs5yy2d
lpMezJxF5ID//Aw58i0W9M1benK6vHHr92YZs/QKBhKe8lQnMRYp6Xu5q90wOzLd
URleQGdN/WPUalKfuWR0t9PR4nI1sWt+A3esjYNI0ChpIihnSodkZ//RLDjOJ6KJ
qAuaAH1dz49lzFqcXMCNkYpLNwae1LTVTLM7JFDiV7ZCkKMhWEA1RHa27MG3+h46
lIyVdD5IjNBWWYMwP023nc8KqiBMHd92yW1vnyEubxfpyzehoqI1N2DJ7XXBXOly
fs1um904SOn1tT4v7y5LGvvRCD6TUuYUyX2OZqw0NNI+r+rgFbcyxmhTl4+FLdM5
KtO02esnJNjcnqXWuW/KmmWXAJZGBSC4cTJPJ5VC76YJZq/5TsM7dTqh5zDIOiaM
vqx49ySAcoJk+bAEgxh4l5M6TQXxKjIMKuyzx8osa7b6XGdegEaWgukM3u67Fk2G
4Ai20S7kFmLjYH4CjMqzWKdI5u8glRwGFFG7SKJP/MsO3gvK8ukr2TP7p/ttuTyY
HFkZOJ2XlI9vxzJ/RHEQ+S3J9D+AZoa5Suhg7mk+dH/szGw2CVVB2d2ASE0W5Blc
SLSoOsI05ouqvGPeTZe53APD8gvx0uEuUd1JsxESzIFuOVRaiJEMTtFSUuDD+Pq0
HzIVQQBOC9UzziSvqiLKSzZeTKFDYrOyvvqVB6R1nmu5vm5ehTQpCaviNtjsCgl2
fsVbVDVgxs0ykpw2yMABeTFBKyyruwBMvE4NB8K/xEy7GiYf9Rh8wYSudmWc73Cx
UHyqlS6CN+2Qo701cxOj2Z+LAoTEdrEZLPblAPsdHVS5uvl6BP5PeDU2vp5++Q39
2zLXOnPJQk5n4pNpFvyuZbnXVslQRPce2NKQPzoSXPvC8RxdxF/PWu5ygLfk6A56
BMaPXlwvcSuqlu/KUtuH0y9Ce+w7B7E0l+kGkVIFVPsu8KCLvf5kqX7VEUAfVqPT
BfGAGgsCSv2TS9+G1ccBOj5lK4+9ubTo5CW0fygIZ4Zgej9z/3kDU9gJP7U/WxF0
O2UsV7dgJBVFOGKulWhLIMCleXxzzWisNDDju5FAaAiGHGwxsrwtuTYya+UmPfQP
OE6z7qfby9oYpbwn+XcmE1KOLdUPBOnydxltQMnbcKVsgH54NMsoN76XYmwV81JB
Bu/BTbF8OgEhr8ZIyRl6bIB9/Fjqrv+P+XNyBt0n96N/j52itiddWyY2TEOZA540
WBqY3COGXJNAx5q0uO46uBvdg4KaqLpb6j56PYGsNWkiXyiZADiTzfcqQpzOuOtO
VQDQkrKqsQwA1KCBXm5Fwed45QaysXaFi4tbGxWIijxsyk5sAD7d9YGzmlYQnE5Q
utKh8VEJwbAfCpaJX4jMhtEfIRMdoFAk1y8lcS9jjE2Il/pxxDvlq6Vy+YaHd6i2
DncxzJ8M5H/256qk5Wr9GsWFoBJx1nT6lmL2KDgWjaQhi+yc4yJc/ZbVs+gSJbdZ
7TUQNLRekI8gj5uhzNnA1MPvbeiOwyT0SJDBJXYliNZG0Es/RptkpIMglBZrhDRI
B4Ja0abtAv3Wc69A/SV55jh5rbM3bRQNnRyz8H7wHJLXetZCHw7KV8Ki7VhlBR7M
BPl7+Gfl/NVff1BpW4I26KEUunB0pHYr0Wcw7u9LDlauMTUuXNLIi7Bw97hKSczn
5XoKBf/j9A5ZxzrJJVnbk+O4DAZx38iiNOZWnOLbkcij415M8f8NYu7JQTU3ilcE
7/U+wrcMmKWaPlqM9No9zAnToENFJPXNk9WEAxfpE7FoERM5M7U4rfpB9Jr5Xozx
U9WA9najCy/o+rsOkDSpov0PWm7QQ0BMoQgJefEa39Mk42iVeRPXzFZP4GSVH7Vn
SArKyDw5TN5ScDjNpJsbno3D0Rl9QQ2jNZZqXPIxuUus5zS76c6ifM82douphqA/
8r0qQr4OM93N/0kmqr0i56wRMYC3eJ3BCps6rTmQf3ZYStEphdAJq2Qd6Ju7a5kM
cBCZg43uH88h8EfSD9XySYWwcM4yEPBmSfVYidmUKwzPp7Y5Q36rasGdVkDHzXnK
yJvaSDSfujFRtehweX33InUfDXHmS0266tQaHrQU/DFYgTnU9Ssbc3oxYw48d5sc
B8qmGKKZvmNLZfcoCMSrjPtrGrjCHDt9/twXSk0IwwL6YhEDVbbIVWCk4XnuQEU9
Z1H4lLf/eRLgZL+Wi+6vEbRRgUkb450WHAr1+hNgZ+fKEr26fRuWEkb7L2I/zoEF
hsyRq/fgpNDsHRsVptXomtO6E3upfO9DskpHCoKJeXhXPRB6wZHTfvOrS5ozkmTR
vf1YyS7tz30rkXu5FwwLG2QS3TFRWNUdtXZQOBeGeZIuCuehzAx3NDFGHhuME0iC
O/ruWigmpA+x5r7s14N7TUnh1heEyg5nvjFbPhrc65QnbVemxRl+rr151XGCPz8P
jbdHJ3q7dQ86DY3/TMDWwEvh6X/jRU//e9S/eDCxHzD4urTP8ni8c8Ti09pW0bxC
wamKfm13c/sN95tUSo3X6a6V2XgoX0pS46zU6DEDZaFZvLDdBRYBtJmvMmgmzrc/
SYWU8tikPKmG1HuL4/qZ8YnPvJPwr+P16pt+nhS6fvpF3ZwYmK5qUhhP0RTo3Opm
puUg7LdgowCPkARoSQ4D0hXfyZGrkuoOJCW7k9/G0xe9+vXobh0E2d4ygo+5tOec
BK52c+OLcngOULUx6mvyzTZrOVuCCq1gDIQGC6gyx1EHNWVCYZec6jvRSmX8YqDg
zVwDmONCJP02C2jpJVtzA6mwobRw7LebwZM8jtvokarmGAkdR1eoH5FcANgM2+Xk
FoCaewVjwWQ/rs2zDGUORySWkSYBFMjFKkmJd3K0WSmB+ue2q3iFIcZPhw4UsbDJ
RS/DAjO4IPBdLQEOpY1FcgrwvOaFJTQxuM4RRV+EKyIUzWbAUZbEbt049/r6IfD9
hADHNHbCAPgwIYGa6MgqEIfbJC1FwUROe9+M44JXdN5v0JVc7dX0WYO04b4O/cjU
RMRnvYlusM2VxH7D+o7mXwumyJbFT8wJ1GbYVsvulcO98kFEx21tfEwWRVH3mMwD
fN9t1lesB8K2eC7hOUUg/K+Qrewk89SciKkgrSuFz/9euq++ZFlbih/geE9jOkus
KlhFm+ALMfPUcXRVXvY+/a+tENlqjGVNDbz/hGmZQoeWQTaisSHn2uXkZuRFpY1C
fYqR5mlEDpuABqH3kjwdarNkxdEC8QozbGSqlMO5RyiI/sPgcZeBzGyl7NOEQKE3
WmzHF9SxDO4JIo0hqSQUVvOTEaZ2t421JZprYJDotYAtYYN+BRhJujFsZ7veB8LC
P7GAupHzPro7OwcpPAqZyfPwbKPVh8n42NIc0kyyUOyiCwSot2FiezUDy99PuOTZ
TX4lX1maHdpmIPDInYNLfvBE955heX2mnO+PfUeHoFQLI5EUtAUTusFvNFtIrp3f
pldFyQfeWD59Qu1DKnQlQ9BbR2IbcB72pVlVTojaUcUos5RWoapJKisaW6C/Kz3h
joDZHQynMeemCeF+GXvKKrq0MF8SkRyE8szLIHzICPL8O9OxLmU1M128ENuxpPzR
X8s27VTjkJtM2O+t1AM7Ded/ZURE7zzjzOEcj6XmwgCnHroSoddainXxtxB5saoE
Uiyb/IGZkshxSarT0z0jsOsPzCpzJ/AJTkC6+aE7OGWVdZwhYJl7P0SygJpaZ7ps
22OqLGITYCemJ8KXnTiYInOkQElQ0J3/kmbMd+MIj4vYrz1m0QWcYmxZG64+MHcI
vmcZeog1kVowKs1aMZGb7XQBMIs/ygLTd1//SvAnswfMFC328kto/CvGleHSEnOs
dRUxAa7B6p2O9jDMhPX+BgTi/hr2NZAVAX5LkdKDEnkiz8N1iOny6VipAUL0hNgT
CMyJcLiCItwyQnst28dMCwJho5iXOhiMwoM1rKlwamPD+LCQT9qIdrnDSCb5vEyb
X7Y0X73LSYsVBuZ/7nKSjZWstF3ZkG9l/TinGL7/KcEh+VQmsb8NgBKN4LciDDoa
oAU+tBEsYSqLFlU2n/eoWWzam3bvfd5jTMR9VN0rAyIJprucUMV2OViDmCdXRKpn
yxliw/7Oy2MaQO/jVOmE6UtCHXWGeCioOJpJdAO37nBpP03MN9UA9wOgQeYlFBPk
/W2QW2klGUXcBZuv2SVCOMk931DR107v1MerIxGk6zbjqvID+ugTlt2YbMOKK9P6
kpHSX+S3LhkDUAiL6n7x3BtRbEvldnBKLcod/GApLYHnRb9zCGWVZAshDxEjIEQX
t6QZkLitRy2z9xSFINKc/6Dmt6an35xwigsaCNOHrc3j8D8Va40Ygg+kaBPsot34
IcL/ZDM56bmRQGiAaxZEk7e5tm2RACRHKF2mOnxWI9UtE+DAMx5VC/4NczsV9/xa
TrkXxrAlMNQtia52DUqJDzPlYnal4gegKh4jV+A4q0xMKzONzqclPUrzCR/l3QxA
ZrKcSQTCwO/4lI7viNZhQ+rJgeitXDDt0GRnJpqKFNppzrfvCVfxTuTlOSe0milf
3D6hy7b1i7Dez4+5QV1eRgAQ0CIZo2P4Wyfm/Geq1uiin7Z1XKN4lb8s58lhidKO
EyLPw+9h0qgrETuLR3AdNKWVXhoKHI/pGkCQ4ZApFPYK48imHL0GVONu3+cezexG
lbnC/WLN/YoXw3m30UE3ACUuHJc6JCWcbiyCfSLka2/o59mBva6A+RzXLJXmWuIl
gZvRJcaIViesD0jJA4eqQAMe5tY95upPOQOEzwaIbECrdLP0TH02Zr2cnoIlk85+
XZxS0DwcQtyiCk10BikYXU5Pr3Ac1GROPheivfRKRAoaeQ8K7MpCp6oIveKqklAX
OweVhSVfJv1gDvmlx6Su2LKioHgNBqgvAJvt0yWmwpgNiJP+v39TszYFG8D99loz
qq2X4yJBKu1zcoaCTnMzlm5qK1VMbf0BBKg+k6E5y0yP2xzWFvN4WSl081nQjXBF
TD+ki2r1dg+OEM2NHor18RG40380RTEMsueQF7NJK9YCkHScevfoFSh8lKnRdqj6
qYWZ4JL//vdLK+22C4jYwrvOgMVohuYReqlCoMvpwTQDeLLp5fchVrCBOEVqfl9Z
vkWEMmvsvz7nLcK1ZqkE1XGCKvDvvQeJXV/1d1qbhg83MRACBhqJ4vJ914Jbkke6
ktM9sFWzt7YaHSQod8z1+wI2nbBp5RtAjQT/BupF8KK84HRVkHbks2W1vZ/lb+NL
ZLodhdHRurZCRrzhxVIdTPvgimqoEOvximrC3ubTkMaVzAhgc40ihLfa6Q5Dui1Z
nRkkTBopgRqGrlevnWxHb48POXIAIDpLapcov1zZuGFU7cscrvt34uhz0wpBByCJ
+rXn5ES2xAx2Jo0vBNd4C3Sk1w5QdWUToCwZCpNiOgwj3ZA9PEADUW2IssWFJBbE
Qj4aSpJBzZafF4SQ+FXWY7v2FhyxLJbPm4cuSbM5sH/7zwjhwAzTCUyWicGtUIxE
c2GEDeq/t2u3cciIJYHiWijN1okKXBcg3/ZuZi2bw9i64YYCmubcGswE2x1KDrn6
DMdPjogU3bdKAf0LUuntSpt1aB/eJjz1TReojEvK6HJryzTM1AVcUtbYRTx5+rU3
MKj55XTGexQZrUPKuLQIvrgrmZszKWy9uHz5SZuOGUjOyOfWKf6dgH/1U88Ra494
dkoWYdo+1U3xPG/0220Y1M3WBtwILG1Q6fvtSrJyg3FF1x+TTfdHeVCMVPc8CXf7
RNhNMvZzBcfxe8s5/BJcl288l7VJX5DeXYJ8rjBH8eQqLtRNG/3jO50kpL+wgS/M
dU2+5eAhRV5kPZEnusbQTJ9UjHfqDa8+/mC810Db5KX9qoE3XhuPQ6dGTQJaTUTi
ak8EjAHKB/fMmO0haxJ1UPOYB4X/Xo/JsCMkcJrg8WzNa0I8mLBs/JEuzuYKF19N
29XdaemF9XmnvIEgyl6IYk5l7wd/HsLBg+tOs0XgJOai/CnQIX2fLRgRGhtmfSOW
a1BOic15TY5Xe/hHxzYK2/y1Tf8NVoaeS5LZVh/OyjOnladILWg8htq06GbslhAp
uXFdX9DMhEmkc08saU50pIFr2i1e70zj3YU7MVzjtWgjRB/ktTn5LCCQhGHy52h/
3KCaWNphEVgmRLAckIUMUP7P7HJVSL6/PUdft22ylaUmiyyVOZllvVm9C8AEyeMV
/tRbLP8YjUijI7gON47aqHo3OfaQMoYh06ZaQEwvZa9lgJSB9BOPt8eF+TSeL1QH
gh3rzvTJnV46zHJ3Opinnim1ZSK1ZDlQtS6VhRwpY3hrFM7EcOOn+9dUWgX95GQ5
wDEkwV/nfJ5dpMLf5KGZbXkkXSXSTAIbVII/0bc8I7zHbGUyshNpGLwOo8JroRGZ
/WyQN5xI8SfTWQOCxTL056ht/jcLhbOJsDp/1exM3GngEozRZt56DP+wsOmaUqx7
MAJR19COdta7eSq8jWbi6avcIR8K2yQD2G3dtUNJwtEsP2UIjlmgXCUnkNZkJVGL
9BlzFMrKfeMlRuFdVj4QBed515B6IRurVI+ehH77kikeb/EpeH0GXLePVfntg0Bp
f8NnaOOWfWICSlRKgeZ1GB04/XeRR03/BZJW48Sx3nyR+eBOGz/nhPPo0BmjA7Hx
V4A1dTkGThxVs0MQZnQQyXCJMpZoyOiXEtS/fY0y0+uToFVYQ5EfOsUwro7ccl7x
FKQ/jQ4aoSmHTNQi2LSq0zJzkrctLYJNcV5kVBgLTlXbGOXToE+AqKYtl075mKm4
r7szbHa3S9LsYdKTKRDe71Uy8nAi5cm0CBOnmMgl9WsdsurH5ZTO0fUe+h3SvNcE
DlxfT7aKir3JmRMCmC+bkY7fhv4fIehN+XlwtOvM2WxStHTNSlDNZLQtf5Wzg6Ek
cMx1VCb8/wpj3YSundioupDz6HWLmNi2lD8OMAv06OdO50IiSJeLDQrBs9o7Gslf
eryQ4AbMvduYteg0Cb5OMGL4w51Zhh0SLHqFWYYtTMgtXoOuqC8CaoxNuUD0hFs/
9DVPJGtuka9DIjt3GtyrGzRR7RlMfdB06MbbssFr/f6/gENV4qnGWQ6lBSsI6wS9
5ELUnWCjlv9wVJGjZePGGieKKO1IPs73SXbRKY5Zy7XwkRJko0JejY2zwbSBCR2e
RBFoUCQaMVfey99p68vEhcOy/CyHZskrygeGiBS3wHeC3cYCbPNM2x8hs8OeWaOV
xMplZJTORFM0v/Wa/L687pJt40sW+7bO7rqG+MHIqI8ra6SF+kI/eS1aIdbN1e9U
NiEYCrxIMdROLGSBFYI7LEP14MxGzx89LxsplsUUcpixYki8UzpApYIwFwMXedA+
upx2wGyz2kDDXslEHUu82DxHl9s27XJHYdsO0SC5+nga4PiEQMq2SgcWXASjM3Mg
lw9xbpFH13lcmavFGfUl6iai9KNxNm5mUxrBrPzgGGaiH1Xr5Au/K5IqDx9QQLif
P32nqG0Xy/W2GwYkpBfXUSZRKXqAPQpJa151ybDtSk0a+HD/JlTIW3vZ98nxpUpv
0pyrK4395kXARD+SY0PWKsYQ43mhVr/k9WXxG+UMDQKNezcCks3d7KRWBl8BIXYo
ulFXjlOpL5Qu0LkxKS5rFz8zzgvCL5EZdshyUleoSrjx1IuiFvOnFvMGqJLXc6Nv
zyjEhDWCRuguG7VZjUVjkxvs+5OUrx/dC7/HxvBLf6zOnM6XZwJxXr7QyW0VcJIC
KkwsT0xsk2mTuy+AcfyT5tZgDpQBpiO9maFIQj5f5Q/AY10MkmZt8HQfYMFaRbkh
U+PuiBeP5BGfZE+WNcRh/VB9h56Z34ClrK9GCj1GbW9azjLPPUaG1EAoSLuWkewo
s2wZEdH+U6Hjxf8ohQAJ0p29QZZn2uKWeVDDnaEvBvVLI1c849FHufIXkdAm3Bh5
7GyfGO0Crj0YyOjp9iyPLG0Ugl308EZumypyzED7uZuk2gR6fvYg1IaCSfd+7san
/XdTpXIEEOZQV/lFqAOiL7evigB2xKpHzQ/0t4hN0BCGOy0s7Exc52NJuQfrX2Bj
xsaHF1l33CuifpanQ2lLiw8rv7iZ6pwkwEprdPYVpjuPCBMpBVrmJT3Qj+RLxK0T
ZAyTJOFjF5iLH6B51A3Vu6+XmRvgETPMhQUcb8SWZw7fdOGe5m11/GqVNzjSGnkc
VTiOE53YBxbybPVc3v9tXkPuCamII6EJT+HRLx80GB5v+iqad+DC8d5nOsICA7Sr
qnoHOevpDppM6HdpaVJZRWLpwXqWA7uEMiPyrxG2qcL9L402hbPJIkJzKF+DAJOi
mPha6PeEVNV9L6qVbaPbt7NhBQQbCeJ99qXdpWF+Ai1H0NyiccETsF2UCipWIYXj
uYa4EA+/B9IiX346DNrFouWXnGUq7Mtlfsp6be1WvRMolgF8Qr54bddf7mYDBDFx
Z70k3WiZE+Y8rlt/UTx5OUW0E6F1gwUFJQfnw/tvINbAbdAMsrKQCX0HmVicIWDt
XpFvl/Yp4B/OxaBaPk0JzymqFh1ACtlfuOqAR9rzaqmej3RuVrc3fo0Xk2+rH9CT
PWFYUTio8nBlqJ3/HIk+igZhL4GWhEGAJdReSkfZOHRG8Pf4bl8H//uSew/sTRiR
r+ZOxtMQGHfB27zvjt+LLeAKzHCWa1MKAARmFrn/pdLUilpx+HagHZ79hODKrgLr
9EzlA7k77gAVKPiu5rWUEeXqjClmXaVcR0HkPWl20j59AnkJ+WRv5IKRJZj6x5ye
E2JMZxVC8z3toJ9QBP4bmKCwlsQsFyPUTmzy82onkxl6BEB6llsQiKnEkXnplTdu
qS/F+/8ZdfUQHx3msIvAtx7q8UtUJ+pOelhJSycFthyvkqXB02qc+jnx+Te7+vM+
CkNCyi9cvAGs+lmGXFqyO+A7lmpQVo5Q8APwyHzgz57AHUb+jV3VvkdhHqpsyTiF
EPP8i8PTw8L0YirVQzXADSGmvRwwNM3T8hhEobUn5Usknb64yU1c8RiqGroohe7v
KGwYrniif7tDsDIBVSxS0ep813T/LU4Q2T18fK9Ocfiqkq10pQuRZtq1vbTzNkLK
VacE1mJDcxosV6y+puLBl2o9dVNVUJvPsrAdPl0HM5aJTGxiXJ9XGNVrpJd4Z1rU
bD7t1oe/3spe7Zga/cfY1yY9R92O0f0K2bdZ9U9uonnV1qP0qGTMog8Q4YD3xDjW
zWE4vV/HN1/EGv54RU6+ZCu+ff8JusZKI+6kZGUx4n6VbT6zdEzvjNqjYVLzffJI
o715tq1XCpiD4K+OLMVDyY8vH/djUwA7ZlOKHGMDuxzZPx22w9r4fn2TuxYxibyt
tKrIGe1yeJCDeQphq9KR2fL30SHZNSaOu9IJpfbu26QbdDDjOnN4Oje9OSV+TTaX
WqrvN6d/xqBLiSWkUTJBi3Kvwxfh3hDnsg1hv/lfZfNH/b23oUSGBYnLuFMXqYqu
Kh4KGPY0ASOUX66wVZ54dZxJnqzFqc07K2MIUzY1eE/BKez6+h8YVX48fnfysg3P
nlo1YPcQoGoTU4ti+woM+DteEB954vDA2TduhwftTEVMsJuztYAXNlBWbgSR66So
kVm9f+8I/v4iKDSn8/CoSwHgpBr+QPq+N4IlmBp9RxqZU23b9zgGasu1vAI+f/iT
qC59t5pgIJ3KQt6jbpksx035EOOGN70Tn6f/tH+pq1kUjS2UkbiCJlYGIYCY75Et
MwKuOo6YQc2EPubQU+4gr0rQ+DQKXZOl0g+apRm0cHBxrklsMivbzxhIhFwmWwMA
an5uRJWgbj+ucVayGd3HvdiDGyA+CLeWEc9hyoEsoEPPcx3Ew1bK1K5yaVgdD0r8
Tr0g2I+F1Lndk6V8duRM+Ryt5ldG6l2NivudNjTcMzBBsMJxIJbJFQIP9/hq81vH
vvp85nbNOECpe+nO+MbPuHD0NXKS4AwKx5t3pgXtp+dzdZJ+GK1PZXSOSAxjiena
sMzUIK+3rtwoidA2SHZFnEniBBq7PYgo++oYy5Zn/wpu5HKfh0qzySXBZNspTfQh
sdi+PmWx3h4361VMgIMeP+71kJYHTEwfDRgrRpmCg6r5W8oxLsLJKCihhKHf2lnq
GdLpv4mZCqQf1zwoP4hsT8Fn0oVS9o8qwFWXoTQcKbO3IyNQrORPLJ9Xou6KaeTo
OHM8VF4MINEUs3X6DmMRFaUYda9dn/77YNjsuIA7lcOrAIyWemakQvcQiCV10RQm
d8WTFFCNYvLlhQti4Dpj+uSHOB+/QDk+aynR9+xzYjb4WvTDi2UGgUIagSGPTs4A
crs5VA0+IChJxk2lCZuHrxlB/v0wmutEaBVmrVKeNm33EhaHk4ETPAz/Wngro6WO
G6obIo/veQ5/9qKuXU77nmRoT2TFAmREHIxCxiS6QVnXfCKWEoIl8ZcbWpDwhy+g
WTHCZ1MPqy+i870nzFuWaEA1ao7X9oMqjuE6EFt6XomO9Zf9vCLOyxFg6dFSKosL
VKKALuZCHlXZQA524wF1oioktBf7vMIHxxmNPHtiCJpKfL4N9GYu6XKo+CM96g/d
/j8IJrus37BPuKOtQyzfugPPnSNsYNnIJfuBpu9qBb68A6R5vFEDf9PsL2hbEr0X
k6wSUWgQeXPcAjHNl5PA4EqwK14w6drl7SV/kbP3RoYYglrcY6Q/SxDJZdoqt1z4
H694D+i92bKPfJtOwxu2iGPPrDqvcFGJAiTkDjTGVVpAZCzo69Uj7RTm61KflaZR
gNpmDGad+txFG1w+iWzd9bE+PDOQTT8rrF7pbL7GLvdAh6hbwJp648n8RR16g3+y
74Oe1MuYpm9/kUKbI1FoFeYL74Qz/Wp5SMz82x4oAE9IYoWbr/UtGAWgQfKgja+0
V+o61td+qUqtV4Vd9MyBWcV99OmCBSwVLTP3aHTVLveKxmVBhZKvJ14/kntzv5Sf
55Mpz/Vqa+p2zsBgEZbgm+yv5qfXxD5qY1PlkTgIvvjkdsVy2cUVmnmVx9i6EQH3
V50wx7zpQxUhG+6/GPs2dJIOsShbQ49+aQNsmcUbXw5AiPjxkImwi2CUG917wOl1
NBwW+pRdLR+fWujujzNo2l1pdSjUznxtJ128bjXiGyYOvt9PNw9NItlBribwyMdt
cCSmcPn9/uw8p3qVPF/SSKuW6XhpQuDc6Kq5HEJs/LA2oFMTqiT+DRUvEVoThdbc
I8WDWRfRN9+6OaVEQZEjanHnwbIdtmUCLFlPdQ4P7xkJwQkr6EIcTiflS15Zl56/
8s8Nnt5sRjoRX3FlYc7WzoyEJW94bZJirn0pM9sgh8iLsJE+3BEdMz0bRComeuMv
Y7TsQTIK/9GvOOTXWb8hdZJlMBERB/QWWoaH8fy3/OR3iwdvM6Rmdd1pq6FWdqUy
SLFBIX6TyMAxVW1/H5jh/vi3yvSBNwgJpQIanyRJsBGJ+DQn/y566U3VJUq5J2Xm
zzQ4ZRzfNNyHBqE6AvBzIUgJyCsTj8ahJwqkZ0k46cgNIoMa0A2mqafU4piYS4dw
4fnrJqxw+jyBIm9LdePLe68dDXvqoMzLNQ0LyB7Pn+wa9wUjjRoHDswXiiJ024I7
Sy6l65eIl0AZOlGTuGU7d51gBVtHN/ZyF0YZ2rZ4oZaEVphHFUIbXWclJpD6hJCx
Yb5KkBUZnNIPfIe5f9e6JWrYAKD2qv5gakVWP7+KIBJvuVwL8nl92Ve+Iru2yzDl
lqOwmbvuCX12/IiXk3WS+dSadxXr19z+Bafy/AYEB/nxA8COV2LsySgj3N83LPPh
4nSFK0rWcGzGDrgLeyqyuYsa7cWUmt07ps7YOsZ1DnyLPNEcbw5w27UJUA0fXXs+
EhEVY5hXddu5JSuw04xYcnu6eItNMN1FDyA1L4gFt0XWprayrSFD3PONa1xAsLhR
Kuc0A3on0SI8QLPcZ8NEeklLBSNmFON5CXYSwsirtMrRJwo+NQUE98kknyQVS0dZ
ocpTAIDW0R3thG9pHNZnQWdYRK/ubMYinrkWvD6INrkWZlOoaiD+SLwiBRhi8ajR
lIDcXxkcR3MSlwXFCigLbRKV3IC417ZZLqe2OICvV/XEVBaNszaC5eXhlhdLHXem
wZLXO0YH4f1XFyoOmzyNWroUBzJwmaTpbZQ/dAU4S0uLXWctczqKgIHyA/E54Xe0
zSa8RX08bzb8jkBwAflHLQVRwZnSCOM4SqDvQkBTxS3N/+P+qn6d2tgZv47Y1st3
KXLq1JX6BnmjXe/Krqyc7Q3YVlt6G2/u4po5Df9uAkRE8Ymkjf9UoVASZATkUo09
4seH2BKyJ1wbjQWRyo+T1fBdpB48yyI9BoiuClLQtp2TW1QaoXXtcZDSlbfR/yCP
KqNJ5SEyfESjQZ36YI23mvFtwZvPiyMtZbvqVnMw8DCVo7LboUmh91R3ggsTvCmn
2Lyk/CW4kpQjmPtebVy+Bgpq5rCWsGQhxPVavlrbGTxZlAmpt5lyI0Nki0XxXnyR
FOMn5dHYpC2LAoZgGD1en1i25To8cZ9A2qWR77TQT833pgz6KC1L8j4IvMQk1UIn
1LIG9DfnBtf4xtaxhxToZ+LMszrNXff/4uiB6hIHcL+rOSvBFp7+KSPsGXBFVWM1
4a3ijb7e9/Lw5nezgSLBIhvYrfP42HfGzoZREKFiXkCzOrguVLgD2Hl0/iFuayN7
mJV8P50rBsjre4zg1WbS+lw4O6AuJOZNI/ytniIGn9UkLmVrGiIQ/L3FwIeS8ljb
KmsvFvn4ZaM2mVSlHmbKPuoDUJtk8msbdTZBIuS1fiKAK+DOvhJ5z3aRYrOIy2UH
pQGvQ2+J7alTSG8rifg2/4t7/DS4tShnjlpNIMbrgSXZgDFi7U7jz6S7yaMpiPo0
K/boj6135HqzPbs9g+0Vm8uwXNqmS8afdIveL8BQORvU/tnJ5o4NgTnB0wY3Zj/Z
Ty7cCEIuaRkqdmGCE6pMjbl0aaWqHiDBdHjgTpOnu8X9RbZ2nOdb1R/lIhyaq6m/
mwoCV7pRb+HHqc5mCP6VTKe01CjsC0qkEkTfmEu5kfuL6HUGPLvaLDNiO/sWKMCB
4IpIzqsydtKPyafYkaRp5UhdJeBOkYp78Gdg8n0N26jlqXGqQOjj41hNVgrSFjOA
5CFlANRvjRZqExVnrDjKxNzWCWOuDVis4xWYHF1tArWPBKfrqqnpz1d6xyoiBNde
kLEXF4VNDnEPZQ2iZ8zZsm34oybn4IMBWRUAX51oH1bP8kPywe3Jpj3B0I4hJFFo
7ZrGyTVrXPUfP/c5GZimkWckrk3I0PKIX6x7dhygg3GGFXY0LCZj11ce+iC/oHse
w8vqk8GoRCu035zZT3S/95rjvSrtyHffseOB5q9V3TSTWCXJsPQvrXL3Pxgfaey5
bXr+/Jccx65ZhNbo5y09Zzs7VJFu9O0IeW6Gl8jo906WxIqI4HHoN0HVTWJVH/XM
a0fEbFO39Lh8QRF+g2aZJc1aaKve4PxKaUe+mtag7TZLXf1OwOxQ81LIoRvPeR4n
Nre+7vso/WuPclAZJWqINv4cZzhrjyi8E/kx0apifhWsD0CDLlWMQWngM4t5st0R
37fslhAOUMBin/JROZb7lsOtazkEUVmFDK8VFOfpkCQg7mANyqwslYckNSynIuh3
NnissFnzSG2aFfLicn+lYAvw+yz2BZP64AjNCBJZuvXvukoame5vlMDTD/DCckcM
IAHt9oMTn0JQfetIctDysqRRto2OLI2v8l/F7YCJmwxH/hJHcOUbt3d07ZlemveP
EZctc144HKVYhUVRWiwJ56Iz5cKkiOigqD5FpruJ7P1DBdd0O3E4aXLSrb6GOCUp
TJoJ2TGhvPOLDlI/UrHzKub/l7TtnAOdGmKT6czPX3pw3EkuGrvPo+6mlQY/9X3f
UJA+jtA7IvSUkE5xYVmq8eN2KDVYHkigdE+35A+6rmJuBFQ55E6qnNH7aD8xpkeV
HSglOySVlm2rimC7dBM9TiBR/4+LuyGZhndsM0qu6olookmui1Kxm0ED1OIXMLEk
2UbpezSbwoubKQboh5/Aklc8+x8iy5PeRD8gsbc/WkZYYYl77KCnAjxcZL0ejLK2
Wgw3jwDuqqTMrjcI5o4zKar/Pz/B6LVSEUck6g70YYrvHGl/IEDZSOiOg0mk3nnb
I151qWFRxIr9ZMdVTpJjaINhrqjXV+fGdYrVfq21sTExeuphZt5QyRtvHpB6LUap
6kUnlffeLGFUsU1A1JvL5+pl38x3PPyFNjpg5T+nE/oppXnriaK7qhfVjXBMnxXV
x2MhDHD8oQhEjZtpiaGtXsgVn4OBHHsEts4pd7q4gDq3YfMvm8s/i3o4sB/XADNe
rvKrBaeqBG4v0XM+AF4MK0bh2zdoE4F+/YBhxjC2yG9h4iq4EifEnW6FCah24xFe
SLwNarFdzzWUH17C2dW05KBhk/p/FeHiDR5YNotAY/Z7u39xC1Um3uEw2oqrHpP/
B3vdUPFWy5H0xWPpwLruL2voYN6sASp1TY8t4cO0dzfdjVx0mQuqL2QBmO9w9XPE
n0PGnz7+kAg/3gPgcFMyPoTFdxaU7NGTGzLrILLxl73sX3u0RXbtIHlTfbu37BQZ
I9y1UkJLXyDUaWDAxeSNUrM9XVi4+lATKjK+8MOw2UY92a5QXKO+PbOPu3sxcgsI
Tj/atBeHqF3RrraKHdbY81cEuQ/EPj3p0DnvMauAE8efRdbmmq1j0ZXewixrXWSW
wUMyBvxfxe2M1XTPjssuH+0C55ognqrfft7RZi0fl3rHgkHkQemp0eoJ0WIJgHAX
vEOfWPV+EytoArrXxqbbBNtdz6IwPL4Tu2roTO58F6IuuzMSzHcQ/vwvm9/983yk
mYQ/LRIRCIA53x4R0C+k06eKXvxMRQFlEND4FlHnUQ0wb4QxGpK/WPaW+O/Y1KtV
dj1jf56XCyeSEH6tO6wIB8oaBgNFGjEON7Tsi5X0cqj8aKS36sMPFrPS4k0nlqtc
2JxC9QTSxA/iiTvutBnmrTOgN99An1y1X1QDdNe2Wt0FF9LFGh1lOrS601QM39Pr
2sESI+zTdTtUpFZ3mDknXurLrZxkUkHGjVk/zo4qxghoh8kfUwqjSY4GVbzYcqf0
+uL3pzkYJSHdAkxd61k8YMrBkqWCoD4W19ymt9OtFklpaCBpwlLxf9VGY3LMfKbW
H63HlSOxkeIArG8truDaq6Hdn/KZn7Cl9knJe5i/NwjUlh04eiTE1jU1xwNgxzOR
HQ84kbZtx/HeKGZXFUIdqibfNp/81dF4PqMDaC/gnBnqprV00PTZFTkvBxFS1nZA
GrGuTpaJM8VpYNT2bnqUNgb/3X9+J7gtsM64ywaQXfag46cxPxF3MzBnwHJHyIBq
Afe/ebuqByc6uypz9SbDQ5u/VnSggowc28hbUarZcgaAIN7oWWXYTZS315cEtSFM
qbjCpINozL6njFRgsQlR0l7iRGIAGivi13k2NDL2/xGT7dZ7OMc2aQChYS3IGapB
Hf8Mnu5B69KZsJmuj+E7nfe+2Xa5ajl64CIuu/zBVbZGAO05GaNhzYGc3Qbv6j6D
Lg+FBrIuw7xJ0GWFiuapvCmHrnaUFlApefLHJa4bDD5MVwBULjh/FYWMjLC77lpE
BcLBNBO+TdDUSvG+3wpYbjCE093T9OBsZfMgoZbWvh7/58l8gK4y1cd8Cn1HwpzC
enYUAmSBvuE82o57gThCDP0NEg/x+b/8OmuBUtzWOCZNoUpPOAAIxMvunDEawycs
Tmn5RWUvPdoOtekrd7UHkIrngu2EvUpY1uUedCgkdF6R7qDccbpZV1MnSV/uBrt7
6xAkDUdKteERy6A+BWj8l40dx3x/FrRa0Mx/InN6sPNUdHVvI5fO3Z7UWebVkvYw
E1H7wnHMW1+7kPRTVS29dsZUpGUPDwfKDMrpSogZpEMrV4PuKYVzf61ADAANWN4O
OkOsMjLBHDmpP2zI6ITMAe60x29JPa7hPKjoWgxF4ICTHHHHFQxESz5VWntsFGBH
LGiyDfObX+B8BiqBF+XHhLT7/Sb6hHS6oVCKpMH4epkLVzE4CvlHf6x09oQ/hS9T
8TX2omygpjk91m8/mU4u4fDzg16jyIFJWwqwH79Qbo2+MWfXbUtQKcEiQK4Ypq6z
Ul+7+dUuBTXGtReeVEhLu1hpXVBXN6UwV6Sh6suqWHU7gLedLNRSqWu36qmJluv1
nZ8eCORcfKz1C5b1wBuVuiRholYJ5An9538dDJZgLy0FKtwymDDb3iK0aruRQymT
6Vy6iR80OzSW5LndkgR2J0Md2syieWt+NiO/Fsb11rXWuA+Gt8VY20YAissw+Wl3
gZQiIB205QhKuQFfwzaqmfaBwBY70nsm0TB41EDPePIkjzJzsHpauqUusuG6vtFs
oN1vh0RLGmGEWNdgrw6haYycR2zmR2KE+8yRpkKgRRTr/KGnQxwfPXunt+cKkGSE
2bxdCUXwG8DMV4r1yd5BuptUqFsarNWx6GRYbAiU78hKHHJK+UstdQmHeWShx/4+
TZcEbbFSA8iG5CbT0t5zJsh8AEubu8CT+o8JGV0NEPsuCyV58Vhd/eaIFfRVa3XJ
hJBybc2W0/HTPb2By6yF3zzfsc1gbSCtnDOKVdD+xwBfsBML/tCVOAV0WJVeJcOM
APb7UtIkwuokhHczCi7oWKEjdcPx0dyre+5nvSSLgTq6NZjhtC1CUryV7uSQ2761
5z/GF5go6muKnu29eZ9A8BaARiyL23A31R9nLPVgUlRpUUeq5NGYmbUEXWZibGiz
6ynVDICNRSVezrwszmchQQb0byzxCfq8hcQ64ymV5KyMW1cUkrWLxjLi3LRaEdvJ
tGYfyTzz3N33If/cHcA+e6MYOGSkS4zvPsD1N2roHAXVjnA5wPbHajQjxleIVEUd
1ZAhdBlnKGtlOCiM2/902x+gCO8Bftga9P0v2iDDgDNh9GFYvtgB5x+jij+Qx7Wt
2xezfrHacUSIgKuygfrTIRxKgW8/NCC8OSJG2Sm31IslkvOc5mtjMeuj7bLEwK5Z
577eyce/k3e4O2hyh0JjXpbgwnSzmiUcFGvUB5Uv2DAaG2xGuQXmb1NVMZVl/OFe
Z9UciFvZtXQv9UUKrcrQs8d+dZ/RSsP6JAXAo7YQ3T07HHTFff1iEjUT5E1lYWCC
7gynZZZtjj8aIOG2RKzWKCSOmBaBulJUfkK7ou1uWleFInGCV0qaRIpoph3WZlhy
JcNryKM7G6LrYhDT3htPDQfThbA+x5XRkiFCcHbmvMj0ZnpMYgI/B/GIm9WcgWso
Sjtj9NDrST+avDw0vbL0Qkfh5AaLOiNnmBOtoIbwHQhLxwXK8eoR/xVGBq+fjCPC
+mJnhJcnbg/soMEJbv3FAATw2xnmEmLuknQNzSNg2aES+MwNcPt1vwFiRbtCwnpk
VDAsVrCZ4pMu4c7ek/4XFHDjTlhMhV/Ydxx40/S/7Dv+KBTcUYiKf7Q8HaYptFd0
e5+5yurahnmoIKy4anQoQLS9HDwYDv/9BAtuUFGHDsOQZovvWS9WHlYgmnn7qGio
a17vIr5OrOZgJYaDnSPo3b1tt98UR3TqhlLEFoXVaVgGIldNPrnBIXlEyf3Gyq+n
Lvm6p5O0MI+aM0JuMur1YIWd5waxI5eFGw5YP09uIrtg19QINFaB4fvH1x+KiJYa
xoE9mw52KsNmjqKnWw2hSdkpNXa2EKjYK6x1h3obmTjR7r4I/G+CvpwT5qNwiiRa
EhOOnhtLE33JObP2rAjtUTHCuoAGNDVqtXZKVp1f7ebXG3+JL8LC7106X/1vPkGk
6Q3BgW6hLpwAcVgFcBaHX/Y9nT2tZ4koAmorT4+5VRwh9U026kP7/aWJjnVJzoP3
gpN3uOKDBzXnoikOaC6RHhrEp05tj3kSXAhJ73DMbC7dz0i8PbHInp1ddVdlolnN
oN7Nn+tTfObQpuxn89a4jvVo4vGqt5jxgepkIHwH63sywWKuPTnbZ41kljaDSEkq
a9CqiRZlK7aaRoxht0VJ5ZLxhEoxPMUOVX1/I94Ippoi22B83GKRAVDEieXN/Inw
umTRIWvqIxKz8zUlznXL2UB4bjgU7GZa58a7gqQEZODULwzYMNXXjGQMkUEvwzGt
zTJqRzFEBZDrAkHoD51RknquCqMeF+l4oroZOZzyZPXVLoNjnZKnbmyBGaUmL/2G
MTz3QfW46bcvcdhJ/iKNFHbrZZA3hLpk4OlFlxKifXtwfdwfd4p+8flY3q46OI/E
kjm+eKZwEvaPbtUTCrCX0mpMyA3ET7V/O9AlEptR223AuYbP+RVhC4DRKZFsdt8E
tGl9vp779qmQvBCANRzrtsrwAhEHTJXOKVb7mZuq7Nga78Klax3uRpT0fWciXfs9
bC+zsBV5uyEsMlQW/ZxUFRT4DUfkSCNz6FyLpSHwnvYvaxRJ5sQc1MdFmFKKXNVI
JW/94YLy9GCwXFLdkwABTLnJoOhH39LCiYuiU1GDMqmeLjs5pfy1WysBeNHx1VfS
iwZLmZIUMc8QYweUFbeSviuRlfXCYwk1ZRs8lvUHCL5OOw2IeGrGvall5pSSUShu
Zc6VFLYZ1mzIssZMvOeBjZYk9YgqpOlRFByYBzLw/WDx4+kDTK22mxUTdxWQp53Q
mjBaPYumJ3gi1EOwBQ+O4NGfXvRO+hYgHKaeV6mTYfonkFCt6y1MIST4B2jsoSSH
KjeYx6fEjKPvcHAj96CbCMdGwfyr0+v9jsKUWdjFY2PbzmcygMPZ+aJ8PwORXSNL
eYFhh57qLFV0tlWf4/2+RDvqOLyCSzrpohBO7gbqfw1OwqVAaX6M2sUHatTqgtFz
lNBfLIbl/GvRvqPrC1VKt7W6WqzSyWbrEddrUFPqluA2hgfixjxXeehau+dd4TUL
RHC/Wsj/Qcn9gaXkK4gQxBiUstN+5HFTqtT9phFIpH5WEokwvBkvmlkZu4k+lc3T
ZjSZxZIcRn6gjhmoKNDbyUu9rfYI41Ku4EjPZBljlxCDVBkMmoB43uSCt346qQh0
BcP5xV71j0XqlJCLnr7+jIcz6umCMiDM/j5mPZxsOve72BKAvflVHjiPjQidh7/n
U6BgF8cvUy3BHaFeNdu9Ex3fMQjIJTxy7tYSPQez+9MRZnLiPdlB0n0873lUUyjN
AIM2XzRgFWjcmy/ZFh4ylZ8iR3lK8LlOF2OWKPfR0ljWYbMhVOETy9Y0netzResY
WC65FjhXxuWDrS02bFyMN4tfxsTzAQ00DDR36n8fSgvgQFR/fYR0y5GdqaJjwCrU
Pg46vB7dzopALXoo9DCy9VappgppCUqWNmdbNHrFMj7eAtVZgpd/3iYDBKCU9vUJ
8q7HAMe5RQYTyXvHnVry3bw3tyUJP+5AdYA6JeePVpnv7kq6DAU7mFkiDZmjz4bW
a7is1UuPEABVy0gyE4WSHCcNE2wr+au3qQa6I7xNk5DPTXPJ1kzx4cyjKGT25S7A
onL3N9tjvh6GoDEqKBAtmaHI6Q0tfyJ2W51UZE8hEEnOXr6cFMMUIDmu+9QVR7pc
fCdonOXTd0Wbtz/zAECORNCq0a2jiRU4wFibzAan+PTWaU+e6Uz/vgEc+jk4h3G+
Jiendb+uV49lmq21WOI0weFd8MHRbkPkOv+bjtakNLQdC2+CHyvHFtc0/wUqb0ib
pG6nlAy1AuiEbWSvLn9eroFb3fU6hsp0Wdu2YOrfo5P4T5inFto4dh40uAEFAQHv
07eKXM3BHWbUw1b7Pgpd0+1YTeZz+pfjU8INgu8UvOB+QHF1V3eQebs/Nxh0lI6Z
uFOZumOxrJZuxE57I8u1eAsl0Nl0Lo/6LXKqM2Sghh49aBwmR9HkcyGs+m6EV1XB
g38X7bBKh+5CjLUAgKdoR380c8uwxPU+8/c1iXqI8/MkpD21jOr6TyQarMzxy19a
A62ZJicra7cblBTGs4583Uj5UTQPqXvgdlfBFbl+bVqraD5kdW2LRa0/VuriLNzy
9f6SlSSy2q3ETB22hO0fv8cKReZkOKemznSnizhfLTNWY62qK7hPc83cRoPtAWeK
ENit9P7ybCs25SmCkYOFH9nBLmcVyNZindgTMaAFy3AoIeM8CKH4Cvd0DZW2PxT+
2f9cxCdDDelxQBbAaqoUmpGJOZdim+a1IAU+iZh20QhzHKpKTGazMzcqV3W3HiAf
r09l6N37qwx34uPsj/qk2ZiKqfloUjj7ozkAOWoecsDRFbBZj2DUF3IIZa/Oiyhy
9goYvMuh2zmGMtuxCS6O8/gwGWY4j2rDpCExpZcc0DMp5std/WJXkvpEhkz9tqlF
V2AcLApNnme8hB7AOJPaWDwb6W0m2r8ultCvXuwCylJyk+t5FlUd/yH87IlrS/5K
IgLvUsn2NDtYonsnONf6hgHqhczacjTp2okDJEV7JdhKDp7fhaN7c21X5VrPhxX4
hhFZpoTATlx/Otabpgi09dR8nqabkBJSWRo5xlFMNNPEPphta+WW8FTtS4co7ZFs
4JxT0AkUVgmbiFr2mAQyaA11HguvJYQ/G6y+JvO7IQTm/0tatIEUUwTRL4N91wGB
KcN2M2DsaRkU7WO0Pn/dhhdesRWaiDD8/JL+sCJDs0+0Cc2tBqwb2sXfee+/CQSR
/TJhMmvELMsf4XsoHkgiKXo+1c2H9vefkmyHaVnyXfp8DYiM7rAEM0Ewm9Aq1DWV
DgzDlLVkjd46Ix2Ei67b8DdM7W+Ms0wS5fgsIOubfIQroVPbFThhQhu6vpV6IDlm
z779lHEAricXf/j5HjTv7nOUgNENAfTkX6hRhQjTRMh5RQfYqiA/NB4/oKC3aXsX
hsKddDuHJw/gT0DCDFO24yJ+84HKuWg10xHBrOV+g3s0NRXPjEhPuAyqhDbCwtSl
YF6U15BLLhEGfaKffN+oiogxKOWT/6mj9leew+DZzLCOls7SaEoMh27KrJpjtho5
1YV5k5weQXSSMiY2Gh4I8QGTk4f6fyPV+ecQLjtI6hK/qer5wu8W/sdz+9sFbHlX
dUAtdLhzU3Dcaheew7m40juLoHqdrFH/CREIeeExJ3SD9u4HJsdMOe4ReG7tBxJG
mB+BDrZ4L+l51/MkY/vXzNhjD+JkQYKPqGskU5mZZrg77gGBdkdHte9ih1bb5vII
edE1lnH0GU1y68sk74Ttil2TvXVXA0QEOeH/nCTAlcMHD0Eo9lEH45UmKakoHiBe
AF7AzF4/6Y6td2Rv1Khqn5oiZW7AWLZ06YRK/9djCzw9TkwV3nl2KfSCvFVe/U+4
sfwG07kpHdsriTlxCphd56DR6Hg7AGHl9XTXW/i+aS7orWeMgGuGonU0YvmQUux2
8PDht+IQsKLwFaNYgasV30OS/5YfjqobZCrIpmwMm0e0P7eU2wqNtk9dawt31GiQ
wsd+fA7ue7JmIcyxA3lFadm8f1n2rozKI+Tu23ehybZGfMqStJqE9rH5VGJOdS96
0PrTCGyHsGQ/actX+nbWzrSX2GtjqkQfGhf+XvS31oFni8H2N0+2JJNozmNmZ4lO
4DkLtsMwn59gJDEeurECNQJvAZA9YQQ0pxcnSbtsyoaaL28siw4p+rNZZUzraFCm
Z4Dx03UKeJxnmiEXpy4HbrOBO8TjvFIrv3jVmEvW0Qji/YOCHzc1rDdcqnG/EnYt
ZQWC1y7h6kgtlzEcR1tYx4HjL2SUzpXEari5BYZ52ARAxUyUWC6t7xJGN3AdlU6k
r4zo/rp9FDLvHoU5E56HZd9RsM0L/76ycB3V4FKzxQTxsgjbZSOaRJNRASwH38PF
d9pFW5xEMK2C4dERFjjo5sAUJOXwkRqm6TaPa/gHtUgtEkJCaFmTgsepXSVMuw0u
IewBZFd5JXXDHtf9iXtbmFwznDmbBC6gcamxBC3LTnTdAEhK6M9PFNOhNeCtT8Jz
qP/Km4yUggtNeQrYfNIxEHhrn9h2NvKYMB222fSbRMXpaftuM5Z964VYrRTwcSPu
OgIGAGmNHrSjwNZ7XGkkWT7BO+JRII661EU5IZR0umo+Nz+gjwh5jseiSFR1QIFx
RW8XWGZNJFQSjDBcku+OsOYvTLLdhYoh/sC5QCUWfPw3Gb12/o+tqdXp/nmBJ17L
0ki5t+Jk9nCUIIfP7XN/wEPwGT3JA6b4dryTNe7RizI5hipzCgSjUE0LRG6CQnur
vZDBQJD6iDw1g4zDRikCNuHMJQG8YLirvY04z0yKmq8jpYFE0nNV3RCz/Utpsh5L
VcsaEQxL8tOanYT51XHvcT2p5KT+/8gza8xILXZB8ahc5QHWY10xS8YFJBEOM/gQ
3xqwIgZOfOoH+M7LKvQkH/SFGbkGFnXnHio8/dlaaH3J0UvO+rTfe1tPYQG5UV2R
NrWZHG5yops3eqmEXEG555quknIq+N6vMybwg029KlCvBzPLz+bs6TXHrwaLjr2i
oU2UMM4NNhtYFu3UGRkDhE8zNYBoclqvTO1fADYBSQ+e7TlJgXXDMZExxI5kX94l
DR9Diltbte4i2rE+8ysNGCNl0YZN3tzvrZmde1pUnPXRGgjnVAhQcNb9i3G94T8e
mOmy9B9MLYGpKziDn5YQFNKQwf4MA8p/gxb47YTvNGtF4evbO136BJHkM1y2IkJM
Eys3NOgCYWKRp8z00BgppB610Tu5JbJwo1Cug38Ot96bLjDg0wJScCBDK9DijefL
IptlOBzeDv0Zuw4h0eXq45toRswaWL+gDm+uTeYeOU4oFMWKdS0S1kcZB1C3Myvh
83JPp4t/vDiXQUgnET6zv0rTX+rYv77+k47R1sCQxpOzsg4qLeOg9pTxzJKlIrC5
6a38d7GzB12GhWlQLszLBOTsLJvZ1B4QbcJU8Teks6w69dDpshdR/bESauGRJto9
DnUZX0m/bjUY3uRjagixJQQm9C/upB8y1XLKNc5GS5yYcAVIzcHRYz4Q1lkZOMag
bWOPimEeM3jmHhylAVo+sFpgZduf7SmbCc5xNbFCgAVkjTStpQaDqPm3kbVSU+od
mjxjo84BTXkkIqA18HY8uZJtn8+U8MhsbS5gznaRH8L9Er8JBHkM8ecjDxIEmo98
rmGR7JdVHiPd/4tNuStGiRwv3wxVL3YM4eIsGQ051L8FfjSTL2FAMXwgNUllIQJO
XyzdDXalkmPwM/0saWKw0Nb5bKmdC4neql02QchmkZssZ80KDCRI61Pnrhf80UlM
2CKyj/g5/W7vVh/iW8GkGCqSDDBPzQ7WeMHYWuno2eX+cd08nJVwieWvL1eQQUFl
lPn/6SQLyrLOuaRMvoeMxxKVSkpHJRzFuFciepPaxDduiO5Xjcu6n6AtQIEvq1GH
vUZuMpHgDHfMYRIJf8MAtYioirqCt7aiaqTOdLXrbzokeIj49jfcre3UazkZkxle
tHsO+DNFrcd+8POp5hI14sOoWwlJ/A7/AnIOQC8Q62jEkHOGhUxpTpoSY2MBp9Tl
Gpvy8GT2w+tFZy7PT+9vB+9zv13mRLgw+PO62tUoya108AejzVkzQWhcqMHi54ga
oEoyahwe4Oz8UxesMv7icvLGUuhOv8P6Y+FUYqJ4iKcvzDN5Z4V5DjGUXcYXbUZt
rhXumqxdT5xtPeak1opLrcjBMDt67DDVSsxF1tDG56ANfNWKMWqcKsEvqOydfvyL
fD22JHQzju8qBxbg4LGS/cYUtO3PbXpnrwwqJeCC/Fd9zi+bMiqJCC8pCf0JlOdl
rtC/8IIMTHkdKWN8HTOpVZeGuQpgl5K/4zsiTjVSVndTGcZ6H0WYw0evucteIlM+
JhdII/2HV0u5S8nEBehwhYbOmajmy1dcExcR7J8zb2SZVm3J0OZylsxmrcIqAhjL
x9Hi6shYPgcIx8K+3kN/ff2MRdKf24AGVu4hkfsj5VaU1HWwvfg3udCzbVrLjL4b
ajVEsppVypN4xjg1IEKl1twD8ne+5A7BuMR7NH9/XtLqU2ZMhWrEiEuIEaTrxCao
WQN4USFjKlZ4XZbzDwduKcbyWJles/+7SlVQu5NqWYVR4Bfvb8tQfb2g4P7NwtpL
QlQUfk/S7I2m9gS+SWrds/zeBFYRx3RfF9FNKfUdX0xZwi4WcxGRU8kCqVCJRCNP
quIY0kOn8xsRLvvaQHMsDnPVYcY16qH74805cpvhRuil5IFhqW8XG61pHjAivQhz
f9t6WiFyWbM6k0B/L8jiHp0Tw3kgYBD16HPBbGGV7y2QVYk7MOcbGsaMqiDg/XqN
ktO4L3I84WlZVroMoRF71sOJfIueZXOJ4JOL6v7Y6Du8+H/YOdQ9JdGHRmebRx1p
ojW3zpl3IXVHwDaIQ23ICQHN7woODscWYotzGgpXBRbooSAyVa2Zxt/DiKJp3lFS
fxKVtad33QgT4kTzB8ll2IM0EEI5bGtJx615wW7P1X8uAieZS/RNYyRIbMLpTkEB
l9X42qQ/j7p8FToHVK5GMP3j3u2WbyZwz+wr3xCWqM8QVpZaNKBLM6cC7r93as2T
eAZps9K/lCORlfUi2+doKIAKi0ebezRx5EqQsCm27isQ9T3n8Psi6TytQ+txyS6/
0M5OGjKRGOQ/Mhabctd8z6JfysDW/wLBHqwcAczmVUf9E1g/1ott8Gl5WsTAVc91
IGRcHJYnOIv+9js681f9S0yogJacGnEaF04I+9+qQrbWYNk+xp6QDm1jcjy+b5uZ
6ju96S7rU+sYNFvzRjPHWVUtty5cllgfEf9dddLpf37iTB0NJgr1MZbWvsZvUlup
+3nhBqiG4uZAyJQON7nrImMcrMPhVRBFeANxHnZWraLF291VRkV7ik2UWJ3V9eiu
gjkUp03qMdCz0do80rQZjQxgddrOCTeDZIcq7t1AA6h4MpyMCuafsanN7nWRn1TB
tAKpPQihMR4OI/2v+/8rEP1yTd9J+paQfcVTdl0KYkIV5TId+Nv/2U/5b3WMT21R
C2TrPC471JfSQ8CtJLY0MmSVe0DaZidYSqT0s96Jv2ghfbkbEa1jCMiiAVvzYcBJ
AJ0AwvcESjDptxbnUdGMqRGvqm/STM55ZODQh9dJd+btdcq92IWOlh7dX4998nHD
Z1pTxyeGrFBxlbfZdVbPWLVRwTh04haH0hy2QIXPFkdi6kV6pJaX6b3I6hiuT82u
+p/EGhATfAcF+SqZ46fKjB6OEC8CBiVsQO9xwkh8dtDGgsKNSUwUZ4bJ6+lxOPuu
G2LnerUxkhMDl36YX9/nqOauFrpDXgwTWMYa2hOrdh7/P4PH3p2Cf++akQ0IKsZf
qMeV2sETxtfVykMXrTkcaMOg2tBW9I62vz4EPeHqWXq4KTbvcdT6aF9w4GVQOHhA
f6dS7+/uaYNHgjlHG3+DfZhbg1YvPGy0mo2YjyfYrv0FHrs3zwfQOKgORi4+Hv7l
njD1EabTef5RLEdFYLrcOCUuIouKNiailZFKLrmSy8idiq582ur1RyPb4mVFSgB2
2R2X3mFXoI9/o+0+GK8NsH21bbqG3i5JxBhR9Wdpb24wCjrdvFiqFNMzFO9ny6Gm
0rzg7DgFVvB4urvFS1J4GzJWeAem0qgi6qsuVh/biM+F7UuzYJ8EVkclyS/aLLAa
ZM7froJlj2UxuCIRFQl5zeQ55rlqZIH1jgnpt8AVEpMD2tN8jvgI6LFpqNB5sSL0
tm+bN1esEBZqx3kL4qXoDqeZL09TgBnKvJXsk6cpxwjNG1mT39l2Q3WH+FPPnuD1
RYSCOIAznXv1QIsRNrfyyXqDNd+L62FizlTICNMA8bUl9oi1341usCI8gPugAl53
STRNl0H/5+EW0ap+uoM1XnyqrFKDi3lIjFPSa+R3dqj/820InXpfX+20Frh8russ
K2LSMk1SW0b5snELs/Lm4dCe/U46R1eL14ld9zPRCD5+aXIiGPhWM293QKm8aXil
5Cw4QKhrAwGwO0ZNBe6esTQ+ksbwmnyrqy3St4ueHHEkGvAgg/0iLaAkd4FXPgi8
67u2q+5IVo/LQBoHrmf5SABP7IamHeuba+yZyTZuPkPAb4DOwawGyjM0AmTIwrWG
88P/6jITCqY09Ce2bwF0MQZDVtCxF5LMAoZTFDnN2hHjoBDpHfn+g7e296zhkAts
VGY8s458/1323HKj16Br5v/xdE47n43rfmdODmZId8r7TK01bCk48CtXCnB8yJ3r
fD56eatJSm/OxtGxO0QPHhdqIJRv/mRxvUWcUFbaSgSjkQmRkn2xDBo6ctqY+Fw4
kUHvyA5rpwFkxicJPgBOCfuvmvO+ymSI2ZU6w/cwSdtoNulX14pXHUe4z/Ljg6Vb
P6oEfhQbf8JWHdCFJB9wwGJERIZrRP3AaZ7p3xuS9t2fZ8eaCapqwBhfdCXv8rfL
Vra94O/JRdT7HGrquqbRXIj74BCtc8y/zzNYV7CU05P6lrcRscDhtL414updk9QI
VZJmAZfKemK0r26SJU26MA0Q8/i8Kh183fT966gmgUrz+wgZTocSDdfH+Sk2a0AG
ZNVEidNfrZqsoTNrMncNU6lD4xv6545eAklL4V60SAbcVWAIupmbylj0g7IPWILz
xyNuXQKAIW7LUlRSOHF2OPODgDwNI5Gv2f7ZPThOHrEhh/L9Szu7+Si6ygMIDTQV
nQthBJ4bsZy30YvflD6R+uQ9b2Dr9lo5/WWhLssW9Moep+rkoFHzo9N/D9eFCeqk
30vVkBz0jlexWHr6YAEiLufhY1hbkYs4OQe9BojEpp3vvEwucj8EfJcS6T0TdRZx
DSvhYGOpcI/6ho4RcdPlq0MmYj5YcMDlY3KEcsaXS40FaM+yblIiYgfe+y5b+KIq
hf48BArHR+nF8ocFm00kBiIcDVeyIHovfcf4D2X5xsGCpGjyRfwc8wrTYB31DJ/t
W/63ca/fQ80/zu7vmd67xvZdnbYz+nidxJOucO22NxXwlOY8Nhb1MStYHpganJjA
biXJWnHAfQ5dV8ryR+yD6AEzGMNaz5lRsnaNa3pQ9t+bPLyh5RngifLcP3iJ+Miq
AN7akPJF4dNyhSrZGbetpQkN+hRvoBcLCdqSjqSnvThzvXUuCGGUS4mJQ4uux+yh
WVX/vbQ8eWuBsrkTShWhK7y0KAZYUq2UzFt62ZRagnY+QnDty89rqfpEGl7BcrTQ
Rf9cFBRyHqQTc0GbdugWzA/ewxATOBH+OgtQDpmksJ6OE5nwLHcqZ9aJv7SalN2v
WA6r4O/ltBmDAjABpSVYpPiAM8igOXrf5i/FosTRvjtx2FRf9nD1ZteJQncXDOeg
A+6Hml1Vy7RwOxTLGDXlYHSv/lu8L0ujba6tQApvWYlSgR+zJeei31S+ZMMdaGjs
NKK4zwXSgC5Jlr5/dvfJLwdAvjIRwu5wyHFCkBfgYBNMotVGkPr6QIE79PsCyFQN
0JJod6EyqWiORHinHiObg1Cykvfdp8IyoAva4MoxFq1hqd62UNXrpRUd689QIhcE
tbFXX7XychbEa+4LhPrBILxSSvGEDbLwQ+zLz1KzMx6ZzWYpulknWRRmUuMDjCdV
J5Td2bEKV3szwPg1uH88nzPFX8pk8VeOBoNlz3vvl6C+lVWqgSRT7xw0SWYpZupm
vDybE9weZYXLJXYyfZFGTGNswDQJnMRxaj2ouufgya8kTJX1TTy94XSMgeHP6PD8
Gc3lpAj1FouEw/8P+P5dmUoaedP+dEy3fiMfOgcpBt+1XRZZx6ogr/o1aWxFywJY
aQ0wpt5pJ/glyAF2eGruWLbyZqC48erm3mA2ZChY2f6lKQRQlZ8Blcbmok276RjS
cWQDtLo3asGwOVIH7H6eRhEoI3tk7l8gIiIcoadI1YVKZUi3OPVS3/K55QHnGuFE
T867rDCjPdLyVPdWvrH0cQ5osunYnyRfSp6b9KnoE3VM1KDG8n1z7MIX634OjfpW
q14K1xoaFvLbmQ94Grv2rhY5tOhoLk6V+RsFbR4V+hlFYdIOT/nq33t5n18g4h0I
taWXod8Z5CA+7NhSKqV32/Vhlnk1eUmGn7ftrIRSJHhLAuVADrF4Pe13f6XNtxr9
sx3oFU5yiDnsqM57FY0p/vkv4W/ERw3E2E5qEqgx3eYMeIdho751p6n2ewRKIy6o
yGLqaVSRDgbuEhuNdQ4I4mHuFKla7LTxGcj+jX+iU4KYy/ah4X96Ret4mPEPI/CI
G4pq82naJ+0EXlsjAHP5zg5PpDzf/Q8SYMf/Llsl4Im68n86E6bbpXeWpy0QoDL4
JARb/wI0JnPQI52jiFrr8RA52AM9SuuwWrXsEKUXkofMB7/i2BXIfEdE1HDocw6r
itPBpVaD98ukvveRkYqGFJ07PHEMT2ZmGQ8cvnPohWhKGY8oxFD4f+C5VjU4RrXY
HFDx3oaNRXuukCwq4nqr1MhHCPwhkMhW9bFv5a1Oq9D6YWhievYCkCaKWYsXyM5n
wU84JM36aFxLlsMbfSTqodjwSqT78qoR37TXBtTtwHLy1u35Pn7KsdeiIkEMsEsn
KPalvA4YYbqIiQDGdq3V/QMIFvvK5QMARgM8HNNPBkQCZ56is5yqIv1L2Q9nvA0I
Ste/iruqzAibyQdsGdxtv55eUql8FkK3hVFmS86S43L/L4xz1AF18VWN+JcGUhmB
x/kFytZ0dL7L9FkOVfUHBEYZaMldPvoxr9iYM1TJISeav+ONG+dVb0BGmPHk8mkW
mfNR+Lt3DZoaVIzhnvEIFHE5MhXzqMoEydTkz8+Ftrez82qmAjRu2H7KBLwgEia6
4qFsvCFU/eSyAsN3pxd2mhaUQnuI7svVRr6AmtF9TMDAbHzhf9TamGGJnCz7W/V5
KCp+X9mkHtSaGoP69x9z4fFSKQBi02QRHcWfSYAXVTZn8mYzXlN6RCLTXFE6Vnli
fQRBEySvSFmpH+jK9eIyTnXM0tTcxVB3Rk+c93OykoVF5c766ltOlcbbCEgU1LF3
DGtqaukAuyXMo3mvpUo0RV9IXFYjiIcK/30uGFAbGDMty4e08GnxVq4BiKmSH4FW
wAJw5VRMbEoHFf0ZMQ82ZomhQdnDd9hK3baBWFozyXIZueLs46/yK3wPOUQ60qK/
G74qpMAnnRpBpd+NfknSgJAXY1sBhL2LkDmPAnBke+q203ieuuVkxMulih1idimQ
gfC+tqyThwDoHQy0wFERnr/NYIBssVFfqs4c6u90+JpSEtHXwP5zp8AgcUN3YuG/
+hxfXKtXIdKwxFYkh7GD3OEyNI6FjHvwkJP+Zf+NpdsBcG0RMYTt/5fQnjurFvHx
PcHcqTIdQISsboxuQ539YCCzdgmOU8NqvmRjj1IfZZpqtdl1i4RQ2dBO+8iBfvPf
wDec4A0WuIeen+8Yz/Q2xeIp42FroAu05BRD1vQDmQm8p0eIBotbLSGdnZoXLfJB
w5KjOMG0UOc54qzK94+XpoUNhE594yYNdhA2gHh7vArT8E7qcevz2R/uuQr64HnK
hgRLJ7ACe604ZwsrWlPoMJScR2WnlheqHBD1CwEmVd42/HhGLSfG9h4eOID5kp08
K832F6L91IDI2vYAwTup+74e0+/gHW8WepWlZaaHOg114gieHjGTO9EnO9OBaQXC
B/55uI0ZyH8MlvgawFonBhK3tSrAcfWygFsAOpnVkz9KfSfg0yDojsthKdpyvOs3
3krDy3VXGB027ScHPxXvt6WvOVs8qJSCH2PHo3UTWURQOL6e1fZHCi7f03LiQYTU
cnfNiCPO0KbwUlEElkwvO2PLoIMLq1QP5/IZ2klcSQCbcD+/f9XkEFVIgcT3b0yU
YsGNCVPcbzyrnobmT5roLO/vBuSWGncQE9vLfhmG6O1pZWcky74+mkuTfST+LNsi
KiSVTLyBlGCBbS1uwNh7p75Bvz2pK7gx6EWAjnjL44XV2xiqHEMJcjenmIg5qMc0
kQMy8E21AXK86Vbs/XVRhinmJaUWFc4I+c7rLPTLv1ZG/shhKqYMMLj6za1gxgax
JV6asZP4tXGp1LImlYP4dRh+u7Dm+kS3qhuJoAOmmGjGonALSW0NTY+yWaL4rHZa
V0Y/rJvQzAPACAjH1IZtGjCelzz2B+OSbmQ6PDF5ptQzIk38LhtobDVc7PzJoAVf
CMFCsa0tRmejg6rH8lc8PfeLG8pNfO9UJiBruUConUI2BO+F7vUX4p86096I4YSC
ojyCnIZ7epYgLIEj/EBoYHJb/XEvHQrK7wzPJ3JuOy/lvvcZuftzg1R5QryjCXtM
p/p9ScPVqBm83DYON86LWvXsqHMNutuht7VBFjv7Se8R7id0jyQMjp14+HDZzEK/
h2Og8ZWXRX5iZQLVnyY1yufVgtAQCCXGPaFUmdWBHaaW63E1aznG2wPT9RNSAJ0P
OER8Y6oXARG96jbvRGdK+72jKiUD6yYQ2L6+xUKe503Mx/Wy0OkCwPdRzdNeKdtF
+chCdYDQlYGLyyWL01gAYMz4b200fNqIB8T3nqjDvQW16JwC7xAapLVC3wUImmXp
hZ4dFnYyx03WuzKuXZV8/wAJvY2NuZiuTnL/lJ2TF+u5B2SzwSwQH+GlYrPeLUOr
AznWNk0k/7alw8PNCrsSqmQqngp2OyccoQhyy6BUI68wi7RRwgg/chBTfXVL6nGF
XM/wvGiJ9E2oboxhOjT/e3SXV+Y5IpjYr16sfGLAxJvUt7SJbwGCIL8HgNeo/1jW
DOQ5jWlctINwgxq/Qy+Tiahrsuf/i+LLmyt28f9MzYpDLKPHRrajo4OOLkz4L+Dj
253GuiLWCXQpMWAjEEkIjFuyDKdhHyvGLPNzhdluq2m6c+nIoVyW58/D+KDenp/7
lDwq0eNXoxKxiQGvgZKn4NnowSfht2ChWFYyDBj5/m9iFn9zcjU6ah0Ewd1XO8Li
Cx7ezimB4l6BmGdx4B3Q1KDZYDJWkkEIho1+Ww+1AAyKB2QU2jvOGZFO3TpNLHs7
RKop5+7tqInZcOgbGxxasyDEul/8uFLjlYryrlNqvR2dKD9lXBRnPJP5RFUOWNE/
1RSUswAT1siLkvFRoGuIQlmpZGCYM0TFRUzDL9wS2RUfWERObF2ndAp/cGcTauu9
m4NdIk8FPAmuVrr+aHYF8QgNv8p+uLI0o6jlJS+G6C9IQKK9nUVBg6XiIe+xk9Qh
m5o/O2ijyMKmqRjTBpPAK96VqbMs8cp8G2NIVWrJfaYdm7IgBWosLRXrhVlGkRbc
IqBoT0I3lAFklaZWyqVk8oCvhPrJMrH2exsLFrqLos86sQM4QqBATVRZobGXzVFD
mbVq5NqnZcBK3WjbYoT5S9Tei/4tKyx1haP7Rdu2sdEN5E0fDO4uCPHfpZ9ai550
Jt5VXnrOvFxKiaFQhydSLdXm2y+TNwW5282FyUNsMJTQ93MXNwk3D/EhRZkTadw0
wgo8IiGFJ3e5GWftAMc09g4vuh1mBNLGd7xGrI5OwhGqvbolY0HuRN9hVftMNlgk
95gZ6wo0mn55coHZHLj+LO/XiBeVht3ZICmp1umqJF72iWWqpX3zrxNWf5Hg4c9B
5TRjfb2rbj136esc30TDtqe8x/AJ2Duyb6PsHzCMkNZTAAtzIx01nnZL+LrjxU2G
S0ZCg8mppidPeekap07yJ/THFii9b3jYCG0DGaInhwUA9/YqUZdZ+sTKyPUQ/DO2
Vc46x61W0Pc7U2Xxux4+eNfIfG4jH3oTdihjgd2c2gp60RzCpewoY5iQby9iVcGN
oYRMkC60P/a467LMHCK3QD08Sx/U4MJtTKI4ZorlBRkHAjzMbSwqwbX+q0x6yKCx
BOVeilyOVMJ8LVh7yJEcKqsvN6PlQywM7CrpVOou3+6BwHzNzDfOlk356PM0bKAI
ARM5NMViQPNiY3z7o7ubLz60x8go+tzrCWTtoOj5U5N3Kq/ucmfPyFCeeb90n95K
jyRrE547/EFPJMqQS3rv441x1MozbIUo7OyafmloDJR91kXmRE8LpfI4mtevhsZ3
ZgVsk8nORwpO5HOU4Jldc+W8f2YGTqP1JQvTIPTYV4JEQdXu+CH4c5URmv/wvS0y
/kdaEeSp8BrxkBUNousnQ64nseplJe5TNXpDnvOjxjN+tnPPhb3FfrT3SFoVk1DD
s+2XScWkL6pKuVs/ubKEif+rrNuYg/USaaHPElIY/q3Tb07UfeoaYk2F7glyBQyP
z/Ja9BWy5ZVoqbNPZgcOidbUQwTrqJikgHIw+a1VmNuI+O0mqPz7xgIyZOsddQBl
Z7jywxLNHsFw9nqgPhCk4/060Ul63Gue4xZTcL+MipnJRuQXMGIFXCKTotNHD3JB
NW6hLqCEkBN4paKnrqRgD0i+rwdzALzF7asa5d1Z9j/Y03CAc4B2nn7KVHxFFDoC
Q1TAFRPO2YPQ6dX0Sf3U5bNFLrkZAkJxhqXJrVqudjnEL7SowSJsK6aewpB5yfN9
oSv2M9e3HDe3XJvicBrmnItzvDNpYt42sKsOEo5TYqnLpLHTwZYzSNKbwPzGVMFQ
J9KQ4tyD0TdtyWaZSVdWySHFhlJj92jrC4EQaGoLLLurwWibW9yvdKRTsBs2Dzdw
JSf+yvsDyODRZdpzATlLRYyp28zPh1xXB7//6rL1ZpfJxQe9jnVKztBHQX5CWayE
NE+V5zxHSFmLTEmiWmiaio/DQewKzKdRAsF9Cq0Nf/RcEdIuIxBob4dJXPVhdyY5
Ofwg6u0XiR+aXZim58jZ39v47QQfDay82HQaZrVAtePta/zHO/m9EANWFS6i/CYY
TtA9h3L/D3fLr/3cUzAU6BtOwFJ/PPhC/9QBMBPlnQhMthqsR/m1ToLKrK1b0c3v
4/e1nENoEXc2omtm1uXL3FDsMNMZL0BrmnKh7/ygWz/o+Tu7Wlv5cd59qBIIFCxc
p1b7KGpYKtHZx22yhbwCHNiP+99smETH9W/9gSqRJ8cjnTwfRLwQIeASjuhxqN9q
xl6/vKQw0CgTxjQZE9fP/V+WR1d3NEVRVbbAUyOSm1aLMv3gxPcuV8/XOSyZ0C+C
V61WFIQOCmY4sW1J+NJ+TiA50CRCWUaABtQCZOEw7m7vd252Y4BrWTpi11nrRhtu
m4Enuf+2EJwpoXL4OuouQ9zfy7wAoFn1HPsFXl5RXfgruy9vmlkusZpZf+Ca81ap
yNAWdqZMSkN3QD9hL7kNwm7o9Zw6Y3K+Cl3DuaBbTdqT+El0y/OmtutESresYy4l
d6mGKAlkVrle8Ye2f/NpSVVZXSBZVxmHGNijht4JQ6WP25GEPtIvu4ysomwTbqr1
Lf3JFMo1ZnuQvTQLSGcphgx+tgypFqZ+142fSEZ3EWi0qy6pLPY5hCi0p2wvdrg2
IOQdo+sDw6ntFNgjH7b/jsb/FUo7EcSGq1BDgVqRlQeIeHcLUB89Wc5MkhfKvYPX
vEzRtY7Z7NQqT8JIgdlQtnaJ4nx1dT/to9XNLuJ/eLTNqIycBL0ZZsGjJR9bS/4M
jr5+A4VCJSlq3/95LdATSJvAJ5T8sXjBW88ZCj7GRGx2FskQ76bjqh0ItQS6AUEN
kXg42SVHrfVADVYd7zbZSJN4A8dCVfphfGxDqxHCsUMj0BL/H2kRDUS0dYpeupjZ
srtCr/H0jVD9Qj0XAqDncWh1UshubO1zF+9gBrbk2fiAoByaJknkj7dBDSZZuP3s
XPcnQxjpQ4R0DuYTgufblG3NlXQie+gLoe0HjbokhSHficO60id4hyUEF6ubRtw5
2HsXzLZfFp0GpbVTOVbAffnOKsQaUTOc+zSApWWM4WxFe1+dxlhHN2WXj+W6Clt+
jG+TxpnukSzOoHVPbcT9Yq4Z+44c7R9WzOziSwjvYSVdcrq6FB+uX1XjMqwj2G0P
LfKhp1Ok+BlQuEzUaXrhmMzfL18j/i148CFR8BkX+btFMgvUronmiSRXZdZiFluO
BYPJOZuflexmM8esLT2tI7J3mA2B6nlC+ZlSuMezWiqwMFKxIuIPoqqxQw5a94lN
Rn7Zihfykyzj1aKnuAkTimji64+Qo9GowFGBDnFfpzSmk7DrcoeoL1fAUVJaqsnt
behnfEoloaKPL+XhlayfpAsJSb9CYHvtlsxtpZT6ahRdZNwEdKhivQfly0Zms1GM
5Ameo9tTmhYiyPFYFkjqiTjRtyYEZMccc2Y51Rntr4/mOlE3pHwC+3VhtjQIcr8o
dHFgrfAy5RL/XFtPd9lQcLANfshHGNrNenp5paxNo4WDl2FYZrpBF/HemB4H0MzA
cNdC6bYtCwGDXqq0xnT+/FMc+rwZgl37/vKvQaL26Wrw1VZckCv1jlF1u9bekejJ
ADAbpHvQhd9Xu0eR/2nnuj3D32b2rayEldXZAvCJLzRJKvIysAbN6gAMuEqpey91
0yHxgMwXABA2faRogdocsstM7EjofWPgdjZ5FMZggnQYaMo6ykJU6OfKy6Dn535L
xWFDMYgDkDv5bOMO4m6xnDJl8AfTaoCtfGlLD4ialb7b72TE3CjtH0eDwcEaMboC
PPzvJe9XEfurUY/XaNhEuB7iKSPmuzrIVUsZl7F+GU61aWvkq+2NJrAe0lvnNHvM
HVf/OX1X7CBE3VWpp6fxol1tuLWlnwuH5LVt32gQQRbSuTGO6ltCawXj5qQfGC4m
JojRp09OJWKgovNAO47FQR7Qo1NcENb4eCjOS+K2N3CACp2mc/EWg9ydMO8f60jj
yhS0DRKFukWpk5MnwPiJhnASyiNVkxTzfIKlnqWUd0ZmhNhPH6PIemrTUCNH/n6d
6UGqajpb0W2CdupvP+WGM6CGb0Jvz5i/xX1b1SBo7R7evCsU0/OokzbiAtFF52wV
9R4LtZBAP6mYL7Txa7yNZs0FPlG9+8rTap2G913NuCEAOWHylSbNl9BUiHx04pYJ
iZuXd4CRzV72CgRqtG8LCYalEsmdb5yjlNRPRx1IqNdupceENS+ShLwApq5jpqO1
bg10HouNHWLIfHBuusyxKoOrHBPXUOB8FPFuQgiQuWoZq8+KgH3aWQWyadjCp1XY
TKqF7JB/LsWui44FQzI4nAXdQDfxV7dACXRdkU09dH8p4Z8Q+AI7XAR8ErxiAOO/
xyVO+PNLSFahdfV3zUQK2SVrqfs9Xo+LGlxplH+QGveqLEGWKyDaJ6YN5Z2yJsWm
KvDsicQVbQ5xGnWfTAC7lnp4/p0sPOaRxvDxL1K+WIjgRIB0/4jkLNRA9nThROh0
HYRT8VqS6ynp1bpqgsc5/cEONvhRWDOhnz8Yl5Y2ekZ/xMF8wahRsJV3YsAJd9Vx
kGXMIXqHbAnVXV9glaASlSG6wlk35sb/SRoHAlUKlxNNh+lyzL6HBIUEKsPNUc4W
MR2vsw7KHtlo8utK0vZqFV7yUv5Vhfr13EUB0+bvN61Tm6aBQkn+rdqbMLPHanTj
FkJwOY6scudMp8G/syWFqj3GH9wX/fhQGe3JdZgkl6Mj10o8XOEPi+ilAAgR3/+p
ONNY9sFbIZJgagSlrpa4+QfOc7rlz++CAUjiEsSV4B9IAX1FCRAqRSBphIsQPTQL
XNyFA+pBozYVwyQzIzs54KpT59gym+Q6H2ReEddeuaCbfGjS3UyGps62/GoAVQjH
uF8q1HZaUVIpfkIVjA5SUgiL/mEnmeTW/gXUHJXfGHBsudW7jkXAIIE4Rf3u0kXD
/sGKKHbjx6LE7Xpl2nMjbHveAoGtsZ13qeqhLEGRf2+rMHfWrJIFyqPiU0fYx5Hp
Vzg2vjz61zO2ujXS5wfHPBipdrnRQJdyjdD9Myab03D8iuBk0nkIb+x2D+MO4olW
/fH7hm2eecvdWZtfIBumGe08ussHUr7GmmkZ4KBOSLcwetd7B3r5Tzp9D55frEzI
+mE0Vwz3THuv6NFs8Jl3yDCUlPxwId+PYLvrkJVDo4jCPoq+ZBqI3R2Tgue6+2gw
VoKg0pxm98LPP5gidR3JWBO3ZHNdEZomLdOvY9wqiBJ6Pqh7Ak9Mzd5DLrDWZPCz
il4waX/DZQnEoFL1mbZxILbOSpMOtvijfhn7cL0YWxWpl84RQLKW9DxeSzs8yy4g
CcU8M0eUjgSVwkMivpsg/SczrHwTyeMppWrhNLy1JjFVAyGw4xdXNUtJqREH1OpB
TJiklodFCfhDCdzd1/YxtzUCGm9+R30TFVC2EW4L5kyhd71eZz/WwzauozM1bges
teahmzqxSq0jNvRGqr3BXIeVX/lTp+tD3PU3U88wTwuPOblRYBldvF0cgbvW9gCh
lG3+jAqUwQDs2aUhCCeEoQsGCYLW4HQ9g6lBO7PGF1c5csf/zUXOnSDaXSMlA96A
88jk7FGDlUEZjH0iW14ipuUI+XzrXkSqA4fsqSSv4XTlmJdMTn+YdkRQMFrbIt+1
lanRJxf+YcM5THIf1Q7rMh8BTGHjcIwHw8JnAwW5vUYNN7jXghnTe9r8l32xLG6s
OikclSPc8fWDuPDz58mQCKSocbvOyKkN7aqOA8csKvufQ7s9XP3jOGOCOnC0L4K9
8YrPtZ2kcrgIsKEKVk5pzuRBZH/Ro9YpYJgkE+o+J8OG9OYqF2GPY8dm4SdsLCXO
U31ptRl14DJyBk5eD3XXtyvG7JlG27lKbRJcVgU2T+lVwzHisEfH324/+WseoNG6
kAc31h1YqCTbvVS72iIOCtoKjpboozmL9X3j1tCErhnF0zPAQP0/tdnNeScQ1lfY
aUeGMXeTujsQQIEdH+Y8Drhu7w5rBeeD1ytR7k4rEN1kaMewJR3o8j+6jD5UmXXf
BsuSMMv5uF1ud4sOGohiHmLoGzQOftiILqYbCWCkQs+WXp5lG2wazmg2PIsojpnS
m5Tnbt0qA3sS344qU9VlxJPUAxEl2O/Bwf7gwMia5Mpba7x1d/rM+/SRNH3otjed
kxsEHVgOKLAkBiISVMOEVGSfZ8ElSJcmG66kXAyGuH3vgClWxJCiCX9sAJuo/6EA
umUfiUmotCscFDsHKqtapG9HPF0JnCHxox7i84UocC6jMHjJHya9rXXMTFs5HkQe
f5SOTGSFa/0rhd0AJBRmgbsxRxxxgJ0sRfFq2u6k39RRdPa5UOTHq/uRRB1TNFLD
elq71WlaN8c2gvpczFHGLyLs5Dn1JauhhlT7N7Q/tEsEZ+rwViIujyU1eTS/azTH
5nsJ3Zy7bM9TXUj6+j3msXZcTkHkKV+354nWRSxwLHzATI8dZi+YPJAaew+gUEMr
1t9V1APjK0t6jI9fiS+GHmc66FDD9DhQSRdoWDA7rs2oieObsV8tNBR+WtbU5nxJ
kk03/NIjnji4uDP/lZDU7xRsqNswutOigStwtx962PUUESzfgqWfSru+DNwl7G9E
kk1VIVKCLaQDqO+O9yTE80pgDEXZgKSZj1OggzLpY3hHU2R3xjsFmtLjXM/h0THz
RQO+MVyZxYsDkq1VJ2lXON/nZ3lUBNQ0QueePZ9oCwN2kL2XlbKdgc6oFfGqz4P/
6g1TNT2sI7ykdYqUyqBPiQB9fsDs8plg4GLj4WL3yaXiG/f+wClVejjzoWquvPJq
9InCJ5wGx2pz0/dKAVssprMe8rr036CsesIEJJSZqKtz1PBTXsZmrbzsph0I2W2+
fd5tyxUTs8HBCAfh+QBkMsr2Z2WcOrQKJBis1LH63pN735/rsY2UFE2F1/UrQeYQ
5H/PdC9bQmrOeAOaRu/nrLg4ZXjCYNgQL4kyly+2SlsPyT1l2FHoegaYbHgkezjN
drQSFq1N+xQEuYFolTlOjDOu+KGPLURwVB55MO0X5y/yqplXzHppZLTzjvenjI/r
5r5cInwhMHChUs3naCTx9qCvO4IUAyxUVkF64rBAh+L9Wd7YLPLPVUcXtFbF+kHG
K73dGGGrG0A6z8xV4FFH92ap0/FRv/NaG0ecdXEaqOiDqFWiiVMSCY7nE1mxRVU3
7wYq68po7xOhsHNb0q+fkDD1HHpfOWKQ7941hqLUQPO1kUz+D/unb+6h24VU19OY
8FFD4tRtH6RQQHjPbQrPOu6/YLdG0RXR1pEP2LOmOS369WmNE/1B+ciD2sZnxnQs
2t8oXvu7mV3uLv2Zd7JXdKewrkk2JDH+Q7AoE6hlSlWO2Je70XBhIHiH+zc0hDLY
8kTFxyhWeSku8OY1DwjCUFqQLUhN+7ZqbVuQToPm8Ju3OfMht2rX4vdKqec3tcUc
JYIsASeUTCGjJ8s7r3F6wyxBHJrSOKQUr0foB6sLqHlY+7O/qrlcxMNLDuuPnPsI
pzOp/ha3OV9H2eLWdevbyG29v9eBoG/BczJMNAtcf1TjT/2q113c7ei0NeZGfy4Z
q7PBwhOrXfaEUR+wgpONkeMfc+PEexd9WYs6e0u45hxg+xSUYIEBh7WjqLrVd9Wj
kLXfuI4stDmHPpqIRTUWJgfj+ab3lGsuD87OfmflOyGnlXRmCoq0ZwEiXxEzwxDp
6G4sDNWeu9gyYxchF42HLdajcjs956fDsVXNWfrb39ucazJpsVZuvuquk4FzGtrO
bLawPgx+Xm/QJiebK3QagIDCMO1EDWiYpBqtSlruTRyXiA18UKxcEbDvxevNKpSl
AEWnfbFGST4AJMexla/FYDunSlwpdj+hIqwvp4u6IOP1EVxdfhgJRI7qic9O21nP
Y/gPvcVOpK1n7XrOHPY6ZfvuFbr2VviNMPTPYcYjBp8pahCKMvTdOBnIRRsEnuIC
YkE42YsJDeTeev9uwa+GtEjuwCWu3Y1lGW2Fb4AivA8MGkOf2fSZefcMRuemZQGg
xThcJvMterW515SfLyUHA1i/jeE0W/OCN3v1oxV0m4VKVEp1UmdWC7zToBp/8BM6
IAs1+y4Y4zQrKLGEaEfzLijhsc7KnzvrX8z2HHA8EWE40TtKsV0cS6nFqahDYkjd
5vz4WWUlkirAirHrKfKO/xpXSEEnnF8cNfipVXgj9kLrZaUEvV8tOETGQFgpFwNX
9txt3aTx1updee/HmlgR1Nh+0Vdjd7PfJKbMoeOo6qQ50tN3CyaszPJpsxana5bV
ThKJTBYRm1QSx3lNJpp8w7iZ3DaCEwWpZ3xs61fCVnHaa2OM8dg67V2Rafvw78Od
p6qisN6OHIN/CAxTUYpBaLYBYMIAA4y2vuLK1sK96i0sfmNUTJVhRgX1bI30C8a9
mS+S5VgyOH5B7HZ+rPDDv6K0N03qfi4RbQOQEYrwtSffAALSiIx+83srCmFfQfdv
GVeYWSIAehw2Vi7sAnkirDCa+R//0G+9h38yyWXJDPq+aB9zrMBNeb/jDPufJe0b
gBbO47tyGWALwKLqdHp7JowDgXuKP9RwKvO+vcnOdKQTW976RJyFQAfmzZWqw/xm
bnMehZ+ZwmdsAC3oach/DCWTuUylTwLS77g/KigpLCe9LsLZty29y6Ks04mrheGv
uF84DlH80OYVpkjpTtWHZhFZB2oQxD/5UpTVBjChgq8fw6FKM4bD2IMYgVV0iBsw
q31OAYC8yaquVAzBw6s18VUys0UkvE6rm3SbRYkMZIfMWKW56+dpl/wMZ56rjE7l
hVwwxEbhyfsjAhQq4aKJgUSeJ9K1b2ZpeteiX0nIX8ZFcfg7PIgAMBtWhJrLbnN/
PApGDceQN+mBHdH2T3yWsO4dO9BQkI7GWdifv96wOYBSbIuExsuiZIwuOR744hBl
Ll74QH6Q4aZV5uvw9FnXmcTNCe2oTu3/cy1t6zhfRtXC9zV6tPAVPSNmkKBuNyVn
FVh2gAVQgx/nltrt/Z9KAO2CInApesp4uFUH1bXnEThZHGX6ZWQwNKtv7Kfs+BZw
isdqv8Rz2Bnl5DvWq3w7CJcp4onvBckMPO09CCC9hZd10EolQY5T/uq5PmAUcEbK
ALgv1gkGziOFHadIZsyqgs5nnAP4qLfjMU3JXti/fz4rdl5GY+d3I1lBSJ2iUHw+
ye5bUTEvkilDayEW6aAyFmvr1hNlVCx2oSqEHvPmktcLmkDA47xWC7PL4VW7cmvH
XmTZE3IyP24WtA9QMxpbua9xYmFljR+W3C89kWVRLXFyn7XJKK/Oo86mEdfw8FVw
Bl3QGcREVJpgjaKn/iJoX2ETyiu9MUB+4VQPP7FfqC/fYGLPS66+AeV5DuRSUYBs
5HHYvY+c7ASZ2lvmvpXQW1uXHR7/TNwqjjbpL+8KKnp3MrfghUaKwfM0InSg+Yi/
4OmQVj/izlYZT27EjbSEnsBD9viHC1JLbFMiRRP0SKhvGZ/16rqVI6LT1uXbT1yn
uxWYRCFROpj/oOu8qFagy+8wAGtVz+mBP6qkOOLxzD08+elh/4cQ9iaT06Hj93tx
RDvFzL0y180dolcl9Hxwmx1/MFmkjDh+PBMQOeLg30qZePiS1y4YFC0e2RDu+zWR
LV3BGUkHGi2/v+ELCMUQcv2sTQHrU7ktVlf9nYIv9QCnYbDnt+ERK3sHJcr0btqc
Z4JYQ76myEVEgPZ/F849yqz6McbCQeHVxq0Iu7gVaUGN0sslsCXp5AJJ7rHVYyHR
SHHaeyJwKOkjqv3F54C91PmhS+XEgVne4xP6X1wAr9OU7Yv54eCBzQhLiKEV2g6Q
NhF7iJ4IscNKOfoFmyXeGF8dZGzHmJ8R0GNv9Xe43GZO8b/8pUZ98MDCXqaIp6OB
GtIElcZYPGRO0mP6WqNjtsAfHPR319wf8Rm/EDtED/bj+ZFskQph34szhEZUnwQn
PtNKJ6nWdPNcjcSRWgOzQPVYkXsNvHqfjqym8/arRvEPNifpu6M291DEIxeSLGRy
8cJcg1qIi4cHpVdrt8ohUoxlS+F8yKVlCaDgZIpIyrEr8gtXMRbou2G2uxP84msI
BvxvEocGwKwAoTGQ06gaSBYXKSn/XFF/ZIF6h3f7iV5V2gs3AB4vAiBYDewpG8b0
82ZBV/Sb6RXZUdm3kf9hZWXSddbuvHaaN7y86ePsFqy1j7jCSr6nJQHhngS/L2Jj
gnlp7ssfyDxC6TyGLjA1JTYFj2jsevu7mmwk/JFjSkpniVGDRkSW9kzDGLgCYz7j
iCY1FdMn+qaU9oPCx0wiNj1uNKWlm+Bt9P//VUB9kIO+w9VcrSLggB9pTGJDlc/C
lvzktLswL+5Otp5KtX+jS2GTWleddhGs4yrV1FGYgMnA5M4DS2hF1FtXocw0J91x
JNEVrivkfqyrskYKBSC8b53mhd2lpX4I8L/UfijymkCYESJqlVBitYvFkyROmYZ3
tQpvHHatxOcoh5vE4fe0N6l8E5B09ePTRJNEsBDxfTvkFNlFxsJYEgMcUFLlL1l4
Y+n2Ep90a+DwpxOzdS2og/DKsswlP/Ih4c9gI5DQTnvPt+tJs1e7imsDeFtpQHGO
inG/UTiGvgVmN8Qzo59Yt9IYQ6tHDDlrKxM2S7KkuEb9yFtk9snC92pOci/qISLJ
snrxC5XUK4FwHpTDudzM/lqxMZnl0mgL0TubvnbCj4GTiI9FDVU23z1MYVD6kmwC
jZMytlpcmy0CO8cZbFEpmqqYitoOdLl6B6qMH5qM3J7jwnxRWmFiQ0+Sy7IM6gEz
BuwnWoaBk3hhPQUAn35iZHOz4pGCO6GPDoXN+YOX1ppghVieHBPXazJ6N0I0Smp4
xM+UFyVfmHjQzooVPePuddUVC0j7KEau7yvDXjI5kjNmml/a+d3VU02y8fLXECKQ
PKydQNNtnFo6jXSQZ1beEn4en+hInbw30tdOlHsuFdLcd6tilso9obcRIo3SU86M
LIEPAg+6hxLiNoEg3pTmjKbRnCpsJWJD189CYky85Iss7vnieHQk970cL+AbfapB
q+7eHFR05lr73HdLdaLBpgYn5LcsNumFinW1iq5SQEBu9BoR6qMC/2ypDl5yP9vS
a9eHfHuzBBpDuJ/Cbv3JJKUUsLHv99YdIy5Zwi0V9rSSMWcb92v3oQoHkK9CC6CP
/U6ii9RsRDj54Q0lIMUFu2zouJJnNEFGMJD7urqRaE+n/6KdrniM9Sa27gP3uHdb
OYkRJ0tQxFw/ueVcs2QNbusWj98PLJHVq00duB1FAZGZ1dm+zEOMufKZHLF+4V4D
9qcy1a9wSDRFaqsui7/5VgNQ9kodni+MqAlXng8gELUNxbv9vYCfZpaHV70Az/xk
BLvB8u/CqzDQcyr68jGlT0B/oZXq+nwqMjDw8sYaybE9PtoieizWOPFvZvyHWjvL
mOs2chWKmk53YIX/zQW5vdIAS+KfAq4FQfij8kJjNjDfLJLCzs+3Yrkksqz2BoWS
GzpXVNkq2wFXUnPJqyeLpRm6pB05XvBRJctSBrhKSyJjSnFaWz6WWpAYF9ILoQVx
sF3CmrTa9tEXQEjuOWpKSV9drF8AxFsFglIbxwBq2+Do9/K3TXRnP7i6c80DGd0E
WfOXl9qOLRHnKzjHb/vWSdSKZhvLvhEKSra+i8d1Oy43654laGOd4NBFtWeyePTY
IjZKVRsdGBDFtChQVFU6sghJCvC1BIwSPz6tEAZpXkScEZx+UlvYAGkh4Ny5xAgB
NGqiN2Arsy/1gSng3gD9nYBOqmqjHq5PohI9oc17aOSyH4V2YnYIGDtRtmTOba4O
K9SyH5xF8dCzfs515DfgV9WmsVZVZCB8pVthrVnzxhmwgcJVIDDu+s8otD76ogWC
w4820kC0QgJ9lGvu4E10JXNUDd4I4F04TuVC7jLaATyZRMVW7SuqZl74IrQGG8Nm
hwhQAdvX4EORYwqPdtq4AJjtVTQW6pBJqQMMQmzieh8xOc3LAwrxVCbU5UF3SnaN
w6ZjqtHl31spQA7pCV6YWI345uTRYDVTenA4ow7z6W5jxhi3OgmSh9/VCP7h8TtW
kWl4OVkSZ6B/zJbo9CluarT8hAqqmakANeKEUDJ2GCAAKZNiMV7YXXr2jZnesv6F
2tDGucKUAnlpx+Gyw6LfFaX5zyT+Rlm+/P8mbGNFzFjsQIr9I90zesAYMmGsD0s4
GQUOT6WXFV+TB61jdloizxdMbWb1x0Yf9qn8GTqx+kMr8FLIiZrNsd1gX4oXpnpW
i/Un1x/qDmbTylCQDSCaeqUc4cMoDydNty5K1AcIU8UvjOWIh7RCB5oWKyq0HDZT
HHJS+1F71udyg03HXK3Klr5fxpdbn69Rjp9sI0aX6eFMU93IvM1/33Unoto+7vcE
Ffruh7qo+ckF4jkeYQ7sR6fvG+PJHtJfHfW1SZjezUn+stbI6NneRybGIOARKeTw
FozjvFbayeOslmF4swv6U4OJBb3GBPX7n8/yJVZ+myo8TzkUdvSLSv+2JPohXYoE
ebeNwq/Ski0rihBrqzTAYlxMs6wpKUZjgcJQp15cezJ0H7n6QXi1ozLKMHpLvvdJ
3Imx55qYD3mVjAeAGRme+fYjfIh7ALAcUqxjNa/DZ1HtFgzMp2rX86DHZ0t0KbwI
91lQ2papv9x8dphyAR+JoKLGTFe7EjgcFi2tK8ZTvZAyJPRMd25g26sBomVXVBku
VQ2f92LfNZHOcYN2Z5eE7gsGf/0/OFYz70Bl88rssX/BK9IDqyLqud0/7rTy61nW
dVJsMcSfTD8jCRx5yVivfLW59yhQvvpNE02P/Jn9NJvydY3G6xpYuL98y40PseTt
mmp7NnhKFy1oFtvuat/8BOdmMpcBST12SU8tXBp0G+Mjklb9tfTUUgMRHsh2+qrF
WLVhOyb0z8YqW4GzVR+Wiw9PALnmbDNag5+jpYz5JIIwIcuHas+PrQrxR9C+O7Hw
6ltfCH++rvnJ2vKjRM+d2MC4CWyfYtca1U+7F4BRi+Fqfdl6jr8c9m+h3aE91ksF
5BNuVBVtI47qrA+Kv34qYQUfKbIv08Rwom5tCMBiUfTHoNmtdedUHV7P+eSFCa8h
ySZ3frgSj46WZRXv7DOMGklTQ3O6OyoUP4miYePEgZOB6AmCXEqw8LhBth5+SeC0
Nh6biO0VJhY7Uy9Ij0DypN+WuOtDFZpeRh0S/iHZOpzjG1G4LYMzQT3B+++B1+xK
Se0b7YdSx2fBh0FZMPOrL/+UcJKz8Q/Pxrf0yxdgU0vpLbJ/BP/Z4sBTHaozX2XY
jR8jvOc4s8fpKVBaHTnvMCoIULpYYOh4o1snYVTXHwHUSFJdZsajPx1kBELR0P7q
SxmBJiHdoRTp6++YTUSrwmO+z3K0cjuSLOoRdJed6QpZxqgilarzG5umjvBUKhaT
4+UUjCmfUIA3RbA/q9FgUIywKB/sRdYNHXi84hGN7XS+FxfpUhFxcZNu6ij2jaWv
287BKmhZsQWXQ2Stm8XlMgkaByrmlKVcN7m1FPe6jgQNaUbNkOLYS4tyXhHI92Q6
quJVRMUKtVMUFt2njRScQrchX7ONb3gFTV1hk5SbvNKAggr7MBYMILjIijs7oKB6
4taCeYbDK13LWpFYnNMrOEmpo/F1fP2OSpZUpRg3FN8Lsja6myVsRo5DDv06qA95
9/GEcKV+4fMKWrq6RREzJ5pnQ9TzfjHR1K0x2asBe/E2LeByIAB3DS4KItjLuSQ/
pQsz9KVc5pjV7EfuF/Ts2bNpJ5B5PJXkTElRDligZGL5b+vz3MvRng0NRD/UssSI
HOdg+GnL3JPp7cYxOab/a12iAzYWdwj0KLL41/9KnnDbKwtRQULzyqe2r4MmaPYf
GgvrQxGZw/zkS1sv0ZV5kVT+RgtzdkE6vTELpRHzuNJN54UDxQXjeT2Rvn/qpwFo
XPkMekamXHiuCBpy9ACjep6sb68TUjjYM1VX9zdcHVBLh9+5FCiPC/YGTPF5ta+I
Hw4HCTB3zu9LdJR+oWY7CX0jBQEKrWsRowNpM7H0b0RuxLLGeP2diyyuSMaGmv73
GsyN/MIsH9/93fkIKpPL6KKeTbRoZr2LaDA8LOwNTuYA2qlVa59/WJljjo209yNs
FZfuJH8jFIU21JmY3ZeiXyt9Ci6/VIpzUj479rZ7nyu5brIm3IGI4ekmdiwyVK8o
tF8+ygneI6y2V+opeckEP1QHxOaTSn/yrgU/5Avdey9ADCPvdnGTUnKO1wwL3dU5
FgqLlItfSuY6dlDJVsFwDq7lJWXzyHlHEY4g+mtS/q4J433k+Ku08gaxMPOgmFPT
929zaus0Jtsyy0giRlXwoqmk/aNQ6WB3/GoYNOpoxCNrrQHpezAuWYwLlzEVYSLe
wBHb4cHa/RFMscVpY04eXfgTwmFXqJ1hfKS281iJxcxdz+9nSCVaJYUT3nBtbq3h
yqtKFmW6sES/kp1yvZcQXzz9MfzYFFKm82Av8hTWcmXyinmnkqw1dFy61KXfqs4a
phsagqW8ySZVtayb7D5uSzZWV44erBGEVM5hFWjVb1ALkwKo1voZoSoaJe4OZDlA
I2nAdqVWv1NjMlAffSb/aGirpBwFnNWjFeg8KvhSwTnH/MvvPrwxuT3Z7ESJSPGl
ImTW9r2jmo1IPLalwBXkD586tjhuf7PmJzA2A4yaKAcrjeFKlLly1aVadJnvJZCU
atK95EsH5p6wUZWNA0dHDxYhyvM0KFytPcZdKIDO57KafNo4YrbGJRQSlxhPRbhQ
xD//6h/B1/1hEnG8yECXR8j//cdaZ56biABFSdgf85AYibisengdTxUNvZzSoz0A
+AkE52VTKCJUcjqAYckn05AQN1hrRBCmXBlQOirykibIVqwA3rXnH7rDLROLTWn7
UUsUbtU7yGaKorLU3INz+tDn0kyLFUopyDlTcfUaTSmeI0UoQmvx0rrprKV84JEL
sKSw/YNXGWPQBgcOHOQGsZpEvEh4XjmGWGZdOuz6grnZvSVYd1/kKxqbD0++wyEE
rjKiO+VeG+LMMf0Av6vt8O+ji/GHhPfbZ1oErdcQ0dI/QU+rJKPy05G2peSOuDCj
3M8cQETXmvaeD+o1ArEDiOKCSjNN7x2xFPrLBak8JZ7Ob70xJpRxvSsarjvG18/J
H5V8uhkBFVOfQEkEu7jhJi+INxHAsJy6Chjsrlaw2q3/WMjdKYJaYzYGn+NUAb5o
OUC99L4dhbQxIwbgvn4U3uOHnM/WAITrYo/m32IzkhxT4TZvIPD7AFFOSw31v331
Df+FYNt8rpwiWwqfqxoWeDxFHH3zQUuZz7dmavkDg+/rKouTKnrl3XfsvEBONSS2
AfNjSZrFdpgSsDqDTL8cHQDrG0/0x/nfV2HxOkqWPGUmSAZvqDLfG4cTMKRMvJzK
APHlfyWunwD9moPl/s2yw9yZ4ywWXuPqxES46FE3JryoL/dREGPjWMmaDYjF6zXj
Shaee4Ofz8YWHnWhEnrBsQ1AmJ0H2csyucUF9CynvqDQWeI1kWCebaox0UkdMXon
DjT/yOsGTfHY9+jd+1A+EGj1ARtsEfXNlQirEpC/kIC8q9r/aK2h8vc7oR6LB3HX
rKaG/jsahjKjH0Czmj0RUVC0mbbsvdkKFDGfqkKUlOEc+iRVqk5hItK/xuaQHn4Q
rqXH49NghZ7PEnz5apWABlNsXPrUQbZZGxGQ2cAieriZCjTt750NfxQ5oLDRgTfk
xW72eMPsUUDM8PeSlNOChijbnWz31go16mjx8OPbOaL4rtbVlPXAQtlLQCliP38a
qVyRUkIVRmE4MFSY54WHfJhDKM3hgwvHwqvA+GmQKp7I13NeOkHX2ZEl6d3Rvgeu
qGqmIio3/Yhvn0kgBGnHnAovVMOxirbFBU5ZFgiQBAfSoDAiauQoRmmzeTYdEq4F
kK5aWvYgZPjv1t2Xfw9hih1Gq+LV0XbzgL3BtsZYG1Y+7Of1d/auaF1doxDUjeNO
G2OoZC6r8rPvUFoAWaPPVaFfH16E1u3cb2XvG88uNhPrIRBnDDKK/RLThv0TOXHh
PBl3NCZMBj3F/F8UvzdRsMHYZ1Nn+9zLzDcuTwb/Qnf27DN9CO1+MSw+rybZ1aqO
k5ExbMJHnDHu3WFPLDupNgPbpiSi3D+Kyr10MstXqmK5DW2ck1yXZMcTFqbeIhfW
nIOy7oSVxtiFqu/3ztkrt7BkMV1o/iBpn5ixGCmBdZmnmBEugBaS2Jm6I+lTKy40
Le5+1k0BI7Ai9NWMsXTojZsWu648wwriIKkExdf9Ty6lU0TiX/7IqC0RZApzxtER
7ILUA+1M7EdbJzhEYU2YiVBKyICzt4ta0AgZPkCeuugIlRzn8JSz9ISsK+/JjPnF
MuxyVhAjhw5ZOfOlPXBKJ2bZ/UxDlJEX3ao02zQNeVW0b942HIYyHbdUK5hJNd3q
whWovfClboBcX6wWkRS+OzhPluCIpq1g8EPlSCd17oc1SzMrPrQGtzJczG66TEln
KtoWURV724fGVHcq4HnGc019c28/aZVcI/AkoYbbYh8bTzfp/XYDxIKuvFFP41dm
DVvtaAn0wfsBHyDzFkpi5KZY9dl4S0dPKQW58FKJqfmcxAJ54aYOoO2iUfMsS3sT
DJ7t9eafz+WKQ5EusbZ1R8k0Q1ampueyBr+OjMi85koeDie346Tta/2G3IGDeqPC
djCF8kAVA2CIeDNRhqSLjC4J3pF6mzFYFOezQBPiL2sFea/o2B8g3KkDNL19vi33
jVuc4VLVmODp46VnsR5lnl9W4+yqBKNyquF/6ORLk1zQCU6BltTpogVqJhF4sFK5
TyTO5Ceqn8C+XTibMlAFVce5o0rnkIqr/QFQ+wDyoEmKZlbCQ7UgdDAmeRJzzbtL
GaHRwRtaM3h/fSDK6ZmFen1jT8sbfpxHjxXLsyZPgQJYTreDmY1KvylWXJR0ktYC
+Par0saKP17sHwnTvD4Mp4cmXmBYSgUPxIKn7TpmRJIeAs8LAprbtARacaMkP5Vw
98FKWYq/GpzMeZQIIKlMxTcE30DGjAke8NZtDW0CbRpLneKM/QJGv26qjc55RPYJ
Na254K0Ms+slI4HjJPsN4TZiwonDF5HhvyksFXxsB8IXP6ajGOrcspcp6aw4F6pf
thMpaUjGu7oEKRSESsu0JgPPeryyC5UxP2CpzTpxdYBE2RSYLvzAGXh1IjPVLshs
oa+KeEFyGxLnJB6frR6dtVduwltuPQuJtkrKnX7h4q0lDzAiEBwCOT4pQ4B6U0Ai
CDHzYR4+Ay5FjWpwmAVvjWQ+CjEufMbrauEM/SGkXy4m8hXs0PxG/zKVrNf4UhSM
Nen2H3cGroFtFq1SKAvWstCEC0Dq1JcMrUAUhCiyCwIBzMwUUVV7zxn47HTm+I+4
lRhYNfA+IWPpA+nopNz0NZoeU51kSEaT+++tkvHbmvqt43fiQxohiU829PMXAkbj
poOkQ66hjj1oAImCQ0gePwZWvpp3o8wdLMQI/Bwf55OqZFxBIkYuXvFras9eaqF4
SxVJM2EXlyXLpo8jPqOKjz8CFS1OgNAGtXaDUzHjqIi9C6f1XVrj1xUc+A3NIo1E
PnZD5GtogbFgSPi9WzzfZrSR/kHkWDpmUxkW9BURXBcPTyuETkxH3ZUisU/vZD9U
tqNpQ7yDPYW3gusKFoBpGcqb1/HOxLFWSITIEh8tzihHz2Nug5Qdj8qE+GOUFpkC
fQMkSmDVC/Q4oLYs197qYdOCzglFRi99Px2eccUbUPhxpMbw2Geb5nSkHX9dfKy2
Q3JNRBXziDVsDqHmkLA11vdzOLQkOF05vuseDk5ZmBij1Zoq8flxk4jk+ZDGVm2u
xO1y91F53uvcqTKoIMXqw4lCjq7c4Gw0dsviUQpKVlgVuR31KNkp5PYXZsP4bOCF
6SGDUdfsJNSMFdVPnsgYu0udKCSU/H6Wn8WaHnTFTyWchSVQgpHH3id/hAz/NpbG
MWgeUYwrwJ8uxPwDBjxB6HQMoptY80S88jjiHRvtojFNaz50SnC/f2f0vTcVCIgF
vgNUVgPp84eybQcdQmXcBKBvh2L/qU6XLr1+x7BjPR91wtg0GwSS0vx/oPRTscYQ
EKWYd0hUsirQTlGCp1MkwPGO1dh+s2XavIevVXGisLh8aOr1nqt5wTLLUBU/xouX
D+lBj/kvPGjjL25VMTLT7+J+TbI+XFpEWARHq1lOFAjNMRQFyLBokSC/s8345SmZ
pIx/X2b9OmWIuWJvIBB6ueKT/Ciuf8xLaBIRC65iOfQhfAkKM4wnb/MeU6kK99CR
tYKa8y+r38fl8BCJBIL8MvQ2JweUWk2uKQHNnYBcAt2Q2nUVMXC8lfi7nThvb4PP
nqmuF1xeQeKd2dvvpZdvf18XtfByh7ZYswoZuSiADMYiO1FL1uR0ZC2DSn0rWvJx
P8AXXYBvQDjEM6RA6CvFxXadta1K6LsCMpaMCOF09yQDlc4DPeWtvebIYYoQNvhn
kia991yEIfNtv4y25VB7gL/T/eY7tVaTqmptNgkxY5gfOExwgR3m1MpatFbKE/H2
rBllPFhXfKyIz8puzTy+9iFh6bF8zS0TWrhSH+yEabaO1dSHNZmQ/0eLM/nWR35E
Lkhd/6jQl3izz31xqEGAvL+KJu0U9EFSwo37acmdWhsdcMLgnoxRRFIeqnmL7uEX
f1aR+OQR5rNVLfTI2H+2cYbOy/bFzH9Df/NZ3KuaZ740799JBY3o5OWu6s/THBGA
ZqP4633MlJxfxqAnu11ND4IFU5O77E8Oxtd1onH+sIfN3mRmi8zGcsql5jNkLxHY
kZO9WjyOZavZ06jreBCLoLL3D9z0ACr0kePG0DPJFZxjR26pLXA8khXi2Mns5uvI
oJMKHw453H0kJcObbHxf7ckv2XEbrxJh4dHZt295xfqHoNt5UCx39D25CDp2oIub
D/QboIJckLEu3xQQt/sjS6i+ghEyQ+CdG/UyvzjoLFGM28ZGlEMgZj8FxN6B1dUQ
TV1T6rywpYJerXiLLF/W05rZ35gxGvNWYRiXGWkozwDtSu93ZXLnX3YUdHGt7OdI
hH0F18/t0pFMFS7Vx7NUaA7cUsBAho34PbhPzN3jxQTHDFhNO9W5y0D0irZXh8xX
JAliMF7grNeWnWXAGs0K7hm00Zty7ihYvWHXmavvmrRh9Dp3al+vCQXopxLXxxff
yPifn7iq1zuGaTZC8/9G9wdzst74iTegNXvihsdmcm9KwxXvPcsqWwuL7r/YhPTH
l7J3aXMrdG1ngVUivUstuyJXNDxHC2IwFjH82IBbAyXXiHHZN95l71dGFWGY8SJA
b4sRq5wqrlkJDiU5Xwzes0nbADZGT7btOz7GK8dQQZzPQWIGgBTDbPTv01h7RG6P
noJ9qX7LxpseJP2EhC5r76agmn++8z2EkMrAj/iIKMtDzxHztFn3bKzqy9kQKVDi
PnwlDT6ed1mKKxp5RGNOrbG+peoZzhTETB5vDegxDIigXzgDuIxmBjARK19OFp33
c6JWN8rb82uEGsOBOURIwOSTJJ3/x48CGUv3HjhAyrP33F3n3XVarNy1fub3gKUM
mQ1g83sdePpECvREnt8NPdgQo69V3Y3nud3UVCKVbm5Guo3zjZqffRBYQqy0wNhD
GJ71dWqAHkL9sR/gZqFTN9/U1Uuv1wNLad4PQoKAGn77Prgy9vZNqVF7TPgvrDTr
1KADG0vwjFqgk+wtoYJLfliDRgGXmF2kidMfHdFeAts8HwRhwshpjlY3vE0GOAGc
7IJTJUu9ouk4Ides3IjDThRBbHJW5I2sdRUdgBzE89af7rslfJEknWYsp67+pMzO
eXfFqWo4Tl6O9qHzIp1VOsUBNqSdV6U5BoWbP506x3ZeWy/5O0RO4BhWN6ZRMRdK
UBzD4cqgjjH2dGT5Q+GV3QBOA+X649GCycv8L9CxogBC/fC3oMhz/w6lBOCEH0T5
mkNXeU7yIkRCIp39qf9YFsUUBfU8Yz+0g+q0//OcC+tUdiqFamEUKGFpiIkgJUTz
r3zYU7dFTxOnI52YNy38ko6yX9vNCpgSb5FX/Es4R4bn+4tei/fSLPwt9cLGO11K
gQYG1zUqlSKSgPNM2CW3+6N2PorEsh4Cfv7ceRcESpYkauy7+EIMeK30NX0KZq7Q
7w0UVtvO1RRDrItwC2akrMW4ee3MGKtc7QAwBCfJ56cQDLXnQba/K8a3YSu3+Zu4
YO97RgiTrIVF6JiWr8i85jmh+dsaQdVOODnd3ORIoM+vqmdwFByflb9LCtMWGFWH
Udf1QwEokYR5Hh6AHvsFmeh49ahwus0ANBOyphFvr4EU9IzgvZuGDGXW1TYRUC+B
yrvztkh0cWRpd4vx277lhbz6gH/FgShVaqySMYfeGQPJBNsbNRG3oUkaVPaJHJhH
Puoul5nsjcwJ0sSFgZTBmAfFdY25KBLFkpN/mZh3XZ+70yIiM8+2feADVJoEVj1V
JGDp71erpRrk5va66m4C2yInET86AjAhHtNZSl0oyCIzHY+8QkbQ3w9rEVdnnnvg
XazEwv+C+wIhQnL4dG1vnwXRAddSMl2bLUjA5aI5XjEGvq4BIK8M6Y+d5ogzdgTQ
mD2S2e0/NDkaIWB2uYr+yztu8vqtMnPKoKhacmq+BwzseC8kjKVjTrkKaMpbZ2l3
LnJLLaD9F3fLHGI3gI5KmkSK+YUH+1U6dmYAZmuko3lozXMpuhqHtnD9W4gM5vpZ
9Wa/fFeAMx2dDTnKCv3IvIt13ZThyY/EAp6vejF2TOria/i9Bkrp0+WS14SXGfKc
5VPl9FMBbLSA6HF49BsONam6bCKKtkJxgFJuch/tB0Cy/yfGNffA172i6wqqSvlT
gucDTYe2Up/SpXR81pNF8/i793ffyusG1IU/JFvbJ5btbBn3EybqaFpxhgvibZCd
x1UU3P+77+D7ymKt8u0xMKECsJRo0j/emXIIFOVI+hvitIuklShtNcLGI39sEvGZ
wm/MpgqOyZcYiO84kAGyYR6rpWH0/xzVoJ/X6xuhQ0eS7zIzOZZrBuBeSFLDPP2M
SF3zQ0J0Q63McTfFqeoTaKSVhxV0znpliMS5hdjQDdRQaoDdVf9R4ksKNYUGHZAW
OSe0l81kGBhMJ3ksxWvbA3pKWXbVhujl0L1hqRd3h9AnjThHQWlYXfhrvcK3/Uy9
S10sMNOE+0EXf0A53t/yQKV4oUd+/WMxJ5njRb2XnHFxOvymjDWo7AGafC0BI76R
08AHG84nmpAqzL9eJJnnfQIDIHj1M/V2lKSsJInCrz/mflRRIuearOFwMG3eeJws
OYkLvuUJ1fXb9FAqDoi2MqDNd0FpDj7RUXVKYFD+mVqgMnb3WkGJEb93WMgQy4sf
/YEgFRrV74f1dfQpp0R70LizMKT/dp20HcbtV6Imz6EVZtWOq90texfO5qN53H2Z
zP87v0XsTEB6ZQ4/rnfMTT5P6nyjRWvg0vGNhySZFKbJLpMxlndYIIyv7GkZjL2p
tZF7ZAUUd1SCGVTYdsC7CQErM5VPLMi5r5vmQ4f/Vv9bPvPSEiaccY5EfTgscJ2r
BYGbbp61bhXWh17DF7ZIVWvOotZWsRfoCV2md4TTxIbSKuW2NJJpBX4X9RywBCeb
Ze/nQ+/WkhcdstXT4sg6JHcP4yyqrqrPUMvL9m7lNA1OEkNOzTfL5wUjZvKi3zy1
9sx5HHgByVkrzt4MguLi+bzEN3EXGyOmgTCRLVPof6EDNRajH/hiEK0VVVx+ZXuE
mKEIok2M73lRpFtxDlviMrxFXE5oPPedUuFMsKez5rg1FFBvUKPQaN1ZJCk+v7cE
kWRrBRa+eh19KT1HlaPsw6AImRVgT3w+Yb9dVKJkIMTSF+vrOu21IQ6vGM9SL2Ww
ujXWUQsqi56OcpYpkDZdkPi+JWBxD8CqWshPNxuNGTFjc0HeeuhnCX4GUAgHIBK5
v3dGgDZsr/hJw4Phhd+YOUmqCxzrub4zkX0upg3x7Oa5hgq0+aJafUrGG2CkUf5W
PJZYTCz75xUBJq8sa/CJ3UIDTJgqBqBXUUzedpQyZeM9q8LVRQvqNbTivabVpl7b
lzdt4HJ24gyKXjsxPAIjRHtFXbpbdiDv45K4lvZbWozQbZNLWVsgRB9w5EU2DD0s
3fsYz6EB1P7Wwptz2mkrNbqi8mudZXW7DkXH4RK3Gdn6xSvk6jd0dQiT6TanYxSw
87UfQGxF6xEvOVF9VrXnY8Tu/AimODAcsvAsgyZQIGeDXLSX8ITDQKxuSqy5fKCf
1MXCgVp/D+l7OBYzyvJioZRK61FpoxgQ8DWbl5yQs2DSXXX1lfr3jt7Xc+dpa/2/
ilhVpCqpSB6c7aKNg1A7qqHyBN6OBXdeUmo6WZG3+iUfWPg6YRJ74k5qfUQIEfTe
T0eQW5rpi8pmsU0UgpyeRgIG4n3f2QOXSQpsDoq172bXY6eXJiEb8qC/L5rttwnf
aPHTxXEyFsRzKFyxLZhPyiOOARyKNjlg5aKUwneMh5qdJI9lZ1sXb0RWVPsgRw+K
UtnxsxsGTzLo60ESXf0yA+zRAl53404U3S8K5njKcU6g6PfqS3zikYQNExpvHBCp
S1aivIF1oXCNQzRYFIHB/qL4ZuNNPSCw64kZz3qu+ZBf+XxXPcRkVyKPqsu4FdQ9
YucqZBLuTIuX8TCiUKvFCn/3dl6ePXI0aoHdABF1YupKJBi7UkHdYJM4/sPTQAGD
Qa1XhdItKmDXVuBCwcKIaLPtM3S9IakiQVCHUo6FUxdjh2Co8pBLCurJXc3fVPLw
WJ8J5p5pACBI7sedMrgWpli8M0TDlNb/urMcP4OVv4yrdIwoKG80jV/0KsNX03FI
TlpImcYX9pDzW/nrDGudYjAcM0JYRh2Sin2W/h4bBPZ+7a2Mn5jg/paCT0MJKG25
BFNq1ftv8KSq3Q/ODqZOcqBZn7Kk8CUolELnSfMcNAxfZvq3Nq7SEyfN4qWKfxbE
aGRY+rmtLxMSSc50d/ysRPrGVHLUoFlWSlEy1R9DLrOSHFeAh4y5o+ZCQMMHu6EN
qUo4vvGA+aNNQJByixIk5H1eCDpXyjytyUBYEV2LlFNXZtja68perUoWbAgqQuq0
B0nRH8iXGUy5mfnrFoucbIOlwpq9bTz8LqNszIR1MmCo29I1eefGOGerxaaZACxs
F4vGaALniptRnXktB8jrOE2t1l8H1LWcPhy16kNNnXjYbduR1RItx8z8ahy5ZaKB
d21EUSN4xPaEyYKoe1q8OOLLnz2/toSTwXd7jPiI8sEGC33l3iA8cqtuQHKbTGja
H7WMdnWYbcWjIwAL+kWD+l39XkZ1riAKgl6lEVJOmN0G3+zsFEgakr0G7O/TQYYh
lgLsCK+e6XHurZ2PhaBcxpGmoKPbV+DStLhnBkadk5bCNYLdoP9UbD67HOWALqr6
GwSgQ+73YSyPs+fkW9AaAonqq6eupoATfZfd+ApFn4ZtvozpavxlxmUgfFt2aQ/n
X5NgYgszLPuu933UT/oAMSsZ7YwIXFx6M6Ym0DcDPUo21Cs3i+06e26LnKBPcfMe
9wpsWckUjIfbNvOzOuJnXgSEbnzHR3LMR0lPj8rZ/VjFfxWIKVDbkfp9nCoWFqt9
6moqw+WW1udz1x5nZvXmOtSsr2WoLPgQNEBbmADezHICunnyeBJNyyDq6g1y8nyq
ArQHvu+4Ov6NOVpaA4hIouZ3f/2vUE+6zcdvNcmRU4p9x+peqacZbOQ/JNPXssy0
mlESB6xqmaHD7fLkpmIfVut7aQtxojDZmyTzOJJWVgRfhvCFThMK1ToY8wo8VFhe
inJQqofGhyEzlnjcp/keCpi6IxR1cF4u2PukFBjYgtU2e37YUbkZaAQ8oiktWVol
ptrRUG3GC71O+326iExWv9xH6nD+Ww5YOAnycmr0+algKU/XPfDI7PjgFcxqPDBx
hC+r4WE32vNP89Ds65H8e3e3flUxZlfmywx+q3Md7S1vZaSMJm2IzPb6QI9AV7R0
Xr+N7Qc2f6mpXo3ZNwtMOICyttAWlD4/7EZDUb0aJAtiDWjnaU6Hreht0z3hV8Yn
vDCbEKrURsm0zxamYzizRlTpogp89gtz+HSZu/lK1WW9eBNNve0O3B3z6c7o/x+P
kxYyWzxVU8pA6/mRi0pgHVftogZE2BRSf7Ih5E0vY7U2yD+hVpo63OufipW0BBwO
v/AgVOLDcRGqqqwlyGpMJV7wA1vDVzc36v54WBANZGSSD4IuFZZoSraEJsCkgREQ
eodItZTR1QSyUdf+h+0PBWCsGoIh8ngJrDiHL7pt2aIdvl6v9nJRQmqZ29RTOP1d
Vv7b0dJEOW3T5KoCLExVy9BrwnM6lGc3Bt6/3VY4ZzTE+PXh8c8wVKdJWua38+In
o5S6zqJPX5RkDkHWv2fEQY4Dt+rDE6qi6FEN62cwIi2CBcmJVSOpdrLLC4PErVFQ
zZDW5+OY8d6P+WzW4RqAHTW9YcVSDaxutm14pxrjJIAvy1LIi6liCYL/ERbnbCia
wdS5Yd/lXPrG6+IJwGUvpSASxWqZzAEctLMf2pS+YSURyl9PvRA44URKuvDD8U4e
fH3VFtYZz1tixBvkqc03aZZ7cCMafaGvrKd/dky7piNlQpGQY48Dpse1hXCOHJGH
kDpX7IzdMaakGIh6rmO0mnW3AkV4KSf+UNlV1hHHsqKlDjIewNy5U9hZH27FoEM9
BIFfrUIKiBcHcg1AyLqhbvT4UYpzferXoNNP0H2BnET1q49iirwevlZWzUlic4xG
aBSPfnD48EqOay1ok6mFN/cPxAJT0MHRqsZ4UanzhodOycgbhG5ltNM400rw5bz6
FeEWtFS/kCsXh4asldWZhR+sJkEyveOdoN8uDKieyNqlGHIGeye2/H9lvI5MmhKp
ahMaakRp/9UDq6WBjOn3DlREZL833jW8awVwetditeJlKZx8G80dOyXq7v+Z/DiB
FwYVy61YPk2pkwM3V6V1lDdCDXdLRIQvLAuO11NxdRc2ACw+oH3kJ8KeDpaJadt1
GxExw3AALhaHxcVL3y09PCWMq3VblIE91pIFp5bvL0W1zIlxxJctJ51riWNJouqv
I4D8btY1naY8vEE7gqyuFjh2rPthvI0okH7EgSPxbc+6eQn1b8XkOu14vG54bd5M
7HHMl65g16PMspSKX2kj50lR1TuBGKs8tzSjsKrIH4nI+dASd+z/TPgbf1X0Blee
IzYF1o/Uk+0IoMQJzj6rhL1/BmyDO40EBGJyvFGPxSBr+8HzoAMEqfVVToEvxk+e
UuTGrG3nC3pJg89dxHnvWptzwFedsaO32O04/9t3I0cm+fGAr9r1uy7tvuU2DT94
2IGgLnGV+bF4L8Ucga8X/reg2NwQ10GYbRH5FK0mdUP/ehP8GRxE0I8sFekq7cyL
ACKep4/m7YtJtvObekBLBlfO9wpUIP7mANUXZCwxg+y76aUf/EmUq4P9CfsiC400
MTMtdPOKiDS9pnMDkN4uszy96YmreYHH0l/JHsGFpjlA7DNgJdxUsm97rDuZcgON
rZ5eq8Oh3JR4mdOlUuYcJaWxlpmtzcIZ/Wm2GCR84vWqk97n0BGbD7YdqNTDpJna
arMq1tECYp9bOF2i+TF9szMrI0h/A4TZDI6n0649Uq85ElFA/0BSWjEpktFG+CIk
gOrVHhnzE1YVqMR2+K20xhlYJxCc9f/8mVCxx5d5i5ld9w1WuTdKInqzpZeVHtht
F1pyhlqTuKNPijyKgZGRCmDWTzqEbzogZ32xYPYlMrxlrTKgYtnlQhNgleM5rDf7
Jdh87YgvmzJmQ5Sw8nfTPC6kd+Z01n+EsYw5LLGP806E+UW04Tt/8kZiSJOxEByx
GW6xMwntm9Dac+rDw+Mrnq7s2fxjS5lVWbdrADj+XIec0pESJksKfdXO1ebAqgZ3
i3CcYFovLf8vcRQ5iCtQ05ya0WAqF/BjBPxqyKo0RGxL8bKbEAjuehj0lz19wcam
G0HpV1GdP5qIDBm/z+nhQA84nxMsEY2fxHOLEB3rZ9xsxzXdXnx9nH40uCyqaH5q
z/Gd19gEkx2Mav9VTXYHqxZ45tdcQZMb+l12HoOdZYaFQTrVGNQ89vxkiQ3B/yxC
Nrh9F3bEctrLtqqRBDrmgBgnpOtQ5bkHY5IpX1QFYIjvlkRbpS9CNm6Lv4gkn+sB
HdfDSl1oiQTXAxMA7D0CvLsMsDGoQIB/VnbFzLFclgcdlPNeDATAi6RTo+tAbs5U
yT1YdXzwzpE7b/KcUHi8gDC9H8XGBn/iopzP8+ZQYRx3NsuLXQ754ZWNAfkdwdky
JjVxiZRBKWH8JkcCLPD8erkQ7xVWDagStWQFX2P96t2gbYcDf2glvhHDJ2a1jGQO
h6mErfRFqqJOH4Z7oybBCTuopkjXKlryYKL8f0VwZOwPZk3geZGaK06LJn60ljbl
O4KFMzUwssarwxE4uzrKbkCKawvibw1kRFJAGq7Y75sT4spzpLC5fuPWxmmnZbgq
NvMbvM3D0oKsHLwcmRMFAMJQAZablQVvplGzCOhYMNJJW4HhuBQMdCzjIsAPOr/8
354aVDNoVz1oRqLz9NQwCpi+KVESbW2edltJvkHfBV4bPgpejqB2FFmmarpLeUnF
KSXL3XTcwHlR9UbQ8gAV9JY3sxJBdJC9dCUm3KX9UozbVPmY6sAUefY/Vv/XohDf
B95GE7ShXKY0hbZqN2mry8Pg+ysS+Zz1CJwAoLhyOhXrlIAq/RPoWCdK+HUb6c+R
UyafJCsknsCikmB9SAsdXF8HiMWaGs4e+n3fQbGkGesOAOzyXDigkfwUZ/Eq8mme
yb1/EbKWtaUmvVnIO7gCL7jekr2+wyuuUz1pLUTnmHB+fp+8p85S+G9SOM6D9xv6
nt0eDTCXdc88YyT2gaDH2bTjchDfQUvSpNOU1jkShf/jj2+IpLgBYEIN5bNkUfIn
TkZOCbhBVEceKImBvVmJM3JYmI6EXJ958GuUGkPy78FOZRluq2r7j36Jt0KhsqLr
0amWlPWtl6zxd2Rtx06pp+7EA3DR2w/31Yh+obNSwRiteA5ALrkMoqDJJnvCqsaC
c/PLRAgni5OuZBYnZERrSnvhqNwL5fm9xi9CKQcN6WethrIcP2PvHseX0qlfm/7D
W7Z2R2fJNgXlzRezKA2GOYM3q1gacOUhIptMGBybIj3RijBXv3Nw8BlzFmq1ekOX
uyL5TDHkanw/CmM0AYKBWcHYHUW5+jEH+pgwbmEig+4YP18dAV4V/wBjih3dRO3e
I0hQR7lLBpRHHDFkzOlBlAsf7K6wCI7FcRuUfYCSafpy6PATO1vRBY/G1gW+x+ao
GxkjZV+8Gf9MGEhapArX7rPH7CxhxyS92+mgHSrP9O7sGMF3nhkvhMGau2qeprJN
QGTqkxMOXSsxeg8dlKYYip3A1l/juQeHlpyaMccDiOktoZ18LwNA2IWDj46IhB2r
78+FyNai4VSxz5X8rM5AbKHJpj5ERjKHybHkXg+KZsYatpSS0nJwI8X17CFKFn+4
ZZiQDQ29j0vK6w986ojlc+b1jxCbbXqqnPOzPMTCvxZ9h7tyj4qpXS5EVnKSIyb+
Uf9Tmqm8IB6a/Mgsy6tUTVJ7GGyrEsOMoB+KcMd7QrWd+pFu6RGb8tal2H+Y5I9z
uahgT/p8v5I7UPjcDybKKJ6i+TDvvBlBalrxFO8BWJW+GYzMF2zUbvqe9q+scG8q
XGTKpFhEOofzK1VLWcYPIsC40f6wE+vLxLco9m/5FpmiqOlR7TxAz6Bb/JUIQEM1
gYUFmmq/KWyxPMn63ZW9SOC8wh/R+fkNML+typFenUfCcJJ/VcDRoN0UQDC/8/U4
P7Gw87Rpx5YwgsOfpaygieO2MBwhTpx/1S7GC2wfweQBCTrfcT0vve7dNBO05cHK
5sEwZq+1cqN5IAyaOl4GV9wFPOTWxAWp0bYUPiLcccGOBDISMg0db0JX5S8Uk2Y7
88QMdQFDIjfA/5GZB5V+q2FGDM9oRI3KQdw5blmFL0kACugATfDLcI/E7p7PX/mB
Y6I+75mi3BxMS7gKcHzv6eNeI3RZNSD/UYUtWlzcN4JQofEMoFwUcl6xkVt9MNLg
VNn12toxqiGowDUydGEd6StBxAzDjy6ZOFhF8G5gEf8PlWfmasptqhhbY8KfBJd4
APfmpisvPy1j5He8mr8g6sr/g4Ny3U2PUUJIAvcV/YzoIRe1UW6XPgBnkk61ClKC
0UdDxcxu18/XBiCPdKF2HBOzImJakPzL+5UQxRe6ElS5ueV3Ldwoz5iX7sYNIwtS
4xPeUc4sGUS5fN75cEii+oL55PyBEu7r+D+l/9pLF9sFaI+XusugTsl7KW7M5kPV
xmwbLnWo0e/srbLfdgg2+Xtzrc6Hh8w3wFr4fSbxDAc9An4jXOtRzU+gurrNd25K
ERlhhTRuVKIhVHeO0EYd1KIvSoEGwqMCZG84Yze5dJi0wXVSateLOI259ueEdbIm
ee84vPfFFvXcFgxIyRecHy8UKqH9q4Wz1rbMNT8+nIYOlv2C7s8Ktlm4JqABKi0C
1HdGj8BlW+Dl/FHLxxy7WEevBhoVKztRDwiUPzMd04yskXB2E5eg/NdG81De98tv
M0d2Zcbz2WiCbglzUJFSlbY9W9HHon50Dp42qr3AW1MusI+OJ+P4WX+uAwvJ7yZy
NG6cEvHsr3x/mHZbmYblqvnm9PUx26xlJNKl6kv0XSlWu/jJAr+S/9oiG7neFp8a
birTgaUJN0cJgvVNEVU/iFYXfH2NH/qezvaNuSQRIaiGZ6LqQHy9TqwaNIeuJ6Fs
BE/x6nrV7qoWNp/f3Q8u+mliTh5yqSrCEkWeSTtGnFwrHEjDtLVb8V9MBjF83OWf
CsvmNZSmN9tvaNtJ7rBSqE3sakbB+GQG5e2G8JDOkPZ10dF+fleinxs3XyVFjOEB
Hn2h1lm3GWt8Dka2k6D2xBbgedGImIDTLiDbXA/teaFp0fc3UCIyeUeXNUUyJfiL
RGJzicgK0kFnh3iClXE8Ts8RWFKHY5Wf2zWdtK3nZZK6Yvs6Di5SlCTGxBP3d8mh
Q3o5Bveylfpy/yTE/QVNVJdZO8DyPH7o+pHNnmZt/L0yToQJBuHGOYdzhdLsfoYw
Wtd6kFdbN/HXqEfFzhAMhxgwiRwjDRJ/7URWXVwcgxWVbKDRkrnTH6EM4RWnZIJH
e3ppIEo0z01tvAJkOQfcw7PahQNCeHKSarELd/iXmI6vjncQTgw0k/YT52aiyAIe
rVuMyVzki2fQ2Ev+VFTgITejBW9m+F/SUpMba5j9goN0o2J6TugXfbKr7vEPHLUN
rCa9JHPnk2vlHV/A4gOcAhjM0hgVcyJ7GDdTPStu+UtIk2cd3JqyERN3PTP8P0e0
MHebpNOMDeLq/hi+GP72X6up04Ge1DvJ3brgYGs4rD38kZWFahj/HC7gKSeOQni0
O+vJfeN4ZVQN7qUA0LRFOvdKSu29M6m9B6j7qGWhEKFq7wF/i1mhXLizn6bWkSwC
ifT7oHLveEAqNu/jAHsDJ0X3UPU+W9r0bx//ci4LNauzEapnrW07oKRjv2zTdrqb
dyuijLEP7KVIv7jwYylKHKH2OLKRca9KQPC6OOWCyz6LVEki78ocefsAGK18XY1f
eVviOAD3kJzGTaUDaoBNH6OUt7GIdPr/c8MkT1PUdIK60zmyQLRcOn6j+hWd+qBG
BM3nKZ5jxjR8KDkfKQSDNMefh2ApS1jWxccNUkmx8JIOyLOY8SCxhPm97HWv8oTm
CtXeUhzlVUBjykVepxHcqc2GRVWIDZdn8Wkbq6zAxcnfuB7HGevKDd2ICVWsG+hI
732eIDL7ZGuZqyAJMwaGWcsNVDdWpLdGXqHgg+/QtdHK08pexjU8j1U0c1JjJkyh
/nb/oiJ9lH9HCRNc2NN7RZV0EDy79lxpP5qlZei+QVO3p5F9Jge25Mlxej86p6Qf
Fmk0+axmyUKj4hRwWCv2UOJzN5gL/YwurLf3Ade8e2Mud5yuo11+gNJXDhGYR7p8
AXeiajTRJO+ggPj0VoLK+vqTQt9rIMyg1CkI5QzeeaBEuXEjdQHhOPhk7NDt5jH0
rdiJA9nefpeLHjDWHhnxIlRarx2kmUE3PPgv86VD7TCKIYR9HJslEIEM4W9RiuOi
XqEOUlszPzKI+gB9WoAfUOtl81Zq+myz9qeh0voycwSigBHfLZksjAZL2zzIyzjk
aNEPQWth1+3gfNT/a1rWhmQJeN8y7vQht+WucO8EqvAEbciTpTp8f/GJUVMEJj8q
xtDGU2lzBA/imWhFhuKzfv7nYLanfCwVkVQNV35G8NhMSG2jOYjlLXieBUxNtKl+
Jn3Iia4LBsj/Ujul02cq0Rxn9i0DuB+BS1o/UGD/GTfZb1OW3JAMdbj7NzkwaxRA
dqSZrXeoMR0wbNYq1hqynRfJ8ufrdgtBJnBbsqF8flGk5WcK5supYvHIL/E9bTKX
muOPdlEwehvOGPVPZe4Jf2KQhxb+Jh+AZOkfLP2Bcz8ljUu+qeWj+kHyx6OU4Ff0
1UK5/TRYNFhFrFiIeIUf22xAkEAJZvQGlZHeY0MmbEpI9Ril6awCijtwulANVdiu
c+lZaBSGej21U6KBCr4tb5kyj5hyoR+Wg/aOOG8386f8Cp94pj3LK2X6Ks3mHSZE
P6jBX0TsAIoRXRUKuOXlBfNM0mxALkGCdZbJzcWDOU4YcXDW/e3DJAl1wgwcmlNh
IIUKjVUk9WbuNWQJf876/mjNbvqdDm+NXq21pIA5mzmcqL9fncLpuMgp4YcW0o9S
aMDkFuxnoAVmve/cCQxdWeNNa2Zu+C/jvHJpOwJtdcROihBHFoybHZhCouX3d1w0
Csu0hqQA2PmmPG9qHzBDOMdo5IXAqWayOTyF9mZLp7tlG+VlPRaGFBA/Kx5dmWb5
yhjQadEanXY+iqzu1qh9vKU3wwVYgjGqhM/zX1LF5TdN61CxoY/K2lp2elqKelpJ
LDBVKkXdbEbec2KwY/Tc1Hfzh0cSiU1FT+OFHhEL6TbLE1AW61A5qPwSXIcoyEbD
67geX+A+ThTw7CY5luJ0So52yhLI+pq3k4QLyw0LiwCEnGNfXHk88UCIkLmFQePR
ldS41Ezm6FGdPjvPaT/RhjJfYH7SGPAw5Y6H8tkbSyEVuG3iGDc9Rn+jzgEl3Ta4
8LTH3VMuxdJ5dkkEP2yK9XjXuIeic5Z40O0c+JCdX0/jhm9Vef0AhdARTQMwJNHD
Y2N169Bo/Yfi2BpOEd5uag2MVIXhhW84Hg2x9+LYFhr8Sv9k6gegk2GbriRJCL05
96QwnF0S2Ua5IvMZse4DcGbdwJtHV112yl+0E5FwjsWSFD382Gusht3AI5aHpfMm
/25IA5oM4N7rPydg+GBe7BCeDt0awPLfmvUQOo+NxEVXC143uBzrEBGZMESAiUkb
Nf+zjkAIOaJ0SXxkHTa3bGhCHXvEkn88DTZZV9heSyvIQbvdshjKm3rVeTpV7nUU
R09JxscIWMmadJayllE8Xr/H/ktsrsqx5G+B8aaROfXW1gR6qbi4huBLDj3Ic5/K
qKPDg/8de9xO2H0Y0zIABdZlCLFUVibmuvpwTm1kC+2F5YkwmOe8NvnsyXVhof+H
1FOaR0XfnoZyxoxINbKd8ed7SntjHtO2Ofocfr5/Y7rxwUuAn2PIy1sZYGyQ+esx
j6W+z4IJWD7ldHwjbFWscDVjpDXcySlEa+XUIg8phqhR/h57grm9xpIZYw/zEz3x
lG+p/KoAhWwPvZKK/q9dNraax+EMhmIocutu+SnPp0ItNM44fjnOk7zkUif0CwmU
rAx5YE6fBD6z3D0SGojOfDuzWBF4hwjM2DzIVVcFbsJAJbvvmGNrvyWsWhVaUan3
giMP3xfSjdQlZdo6ore6ny0oTlD/2ZxvKn5wsu1zBDnpRHXI0fZP1pWdQfb2rUTf
oxKXD8oUQnvQdiPVyahBeCDrzyx7HskzymAhupqvBAW/htymhhBdUY142c64XjyW
TDFdfWVL0j0WXyQbRJN9zTWREf7z3HtF/Q3teYQhYf4opaCcU+xjNLzOVlVc4iXH
LprGCSmdONM7lKq3L5B7BJmDCIttHSBdEGCU+bKILWNUQwXzZoWYrmMafN/pRRHD
Vf60cr2KU18FWcSVqVjQxN+tqBapCwJlrCgwSUM5HSIwfOMeLh6X8AmQDMieIhSQ
zk5PwAcY/rxG/5JAHOhxkdUGiVZHFcSCK70uIb58MCtDc5lYVt9pJRJrQbouYT8X
iln8AL4dPT3oA78mHbgH0zQgfis+QF1BWI/FTNlXXuKzIqfnwjZj1XT2Uyubmkko
jZKub89aKuY5inymtCtUdwnvcGp6sF7Mp2+VEi6BjJM8Zeir+rH/Ojh4HRdiVBkv
HV1V9+kSCWdVy+8EL+iCX/20R5ti+JnWyNoWtEHPz4+LBuazmIdJ+Ve31n8p1iQE
EyEFaK3pienFFp3RXtl02hax149b/ETBCqjn7Cp4bEQXpwFNuR3WuE4exDV+JSkR
HLR7lWXQKIk3e/AqobtjZ0jSsPK4pTjFye6zbQN4btKfNbiUcb5xslPFQPj9iIsk
uz9j+2KDmS4xakoNnksboDx2vGJUFI9r0KOw8D6HTliB+IA+2NPSiwLXTlvJcXKi
mmHi1w60nJDlDahTB4XtR40nPX6sARuALEah1hPuS8CV38Bc5VvAj1JdoRCPTfln
Ypf+TN27r8gQiKLCDzwcnmATA5Jgd+7E6zIBAm3XyamaF723MrlfFH0bFTvEkjZX
PvS9xzkP8YRRQkNqwvBRDlL7B1E8SMlRmdymRV48ShGxqaqSHvvxqJ8Xcsw2qxme
PQ4YT+QMM8cj541sCVUqrKeLG7lQga1hsnf78jihrvxeyX4SdR49aNTNg8YpNm/Q
nNaFpcAuD3XCqxs7rPe7Y4x+/3ufAxhCdPZROed7jZS/tTiWfJMCuJAYyiIruwah
nyWpg+oi/QEJhVdI8axYAJ9YNVUZBzhdgFLNXPPU6tDgiDp9e2G8xRNM/Ihf1yAT
Xjh/0q6CmWhCBrqhON4Xut0dhrvbIswQB7alNpWY0PzAeQFusH7rQsuqdofkle/4
iGabStXF9tQoFjSeCd2PE64NL1fXZIizSJvK1GU+viIy1x7XC4ja+eLUZgbyTd/m
VHO0ZXxFT4Gn1grfnex5cpkjQyp5/iZGHcPOiiqKDvHQB2MejUeenitCYN+Zj9no
JIiLhFDZ9K4HUD1TWtyKTAX7KBw9TY2B63KiClCYFSpueuQPmIs1RWo9zP35/oVa
WrqSMjdyWW8xNedFcZ5IjhgPpUaZ3nreUALWFnlbfRd7OLl/3gtMCtiNYxX3babD
oOHG/XrkfGLCrf1fPM5PzhNWWraonJEcrfjdEqt2a+vFFCXZ7S1bWS7p2idVhp7p
Jo46Akhvy/H9QsuvSDOEcdjEXIq1CK2zlyNDpCiO0dWGJakihCQtqE1wlo4hrUZz
wtfLamvEVINHmWBNAaKiF0nUxZfNN42LIYwjQCHXHHzBbbjtvk3j1m5MOKPVxTiG
+vgwRlHeDdYcgSX51IV8ZkXUZlrYLw25wjFmymu17UIDJMw70xB+5LxzZ1cELxOd
wlWPt6h0n993Y23X46yhI6YkUIiEAtAxaV2es3boI7Wxa1+jstPzcNWGlU3LKYJj
XjTdT0e5wK4y95VsOzxkXX8G3yz8ObufuyDznDkdzgNUwdkVSzYlwZsngJJKS4aW
GaIhMOsQzmIeh8w6jZHC7hd6mo+RIWUQTNipP+5UlTMsOXLE0P+2fisnevj7bhGb
svCtwXqndrTZAsqUfcN2QlR36kApcVkbZQ0qsnqbJTb8eo2yvbu37d0neiqbbNb/
6Hw4L3BW9XHFhM1K8CN4eMCvxcZuDSDXaGCrsz4VWxaJT6W78nUdcAtEqnQ7x2Pe
SUiJw6R4ah6m7Sfarxx65sJbN3NDOCUhFP3Zg5XpE0jIk823StB4vqxqwxxKN+8u
uStkYG8ijUHpDa7IN+AOpvkC8vfRwm0v64JaZa2Q7BVulFAY5YJZ70MRCr+P/lh1
5g8bg331jMhWa160NdalCy0hDFw20eVqqV+pBKdAClVhbKrCO4Z+sbfhR2oC3uJo
O4wwuO3YZiyt7snk9wFyRDjUUclrDC0esRyGY2oEBsoLvX0PRmSG1sH6tBMpN2WS
eoPLL9lpym+muaZgesqxen3W8xeSrt1Rjzquq0Gkw91euiRemW73h0itF497eoBc
HTZtls2nTDm9pr/ccv4G0xQr1g1eR2F66peDkM6gHLcCwf9Ae4fno6cfj/7cEwTH
Qcmnb/XXle+RueUdvTFSN7qeRRVLgtGoDfaZW/scVGjjIft9EW7IZFjiBLlZKhId
WOeIjKBbxa1nqIj7xEfxNemnYcTlS/1Dy6FQUKlJbcvWOtCJMbMa7FvA+nvSPHl6
JRo7D/426n33WOJh11GXfC05f1MV720wgnA8HlXZ6FMS9B6CblFSUnc8f1N+ypy5
hKJmXsNreNZ2Xg8Y6kvikhNgEDCY8/TV752UzDL/XX8bC9h6i5/uTapLpLFdf0mA
7ikgSszqfg0jBfsfNS25xz34zsXxGDqdUgFXW8+Z4/tmke/5d7EVGLdeUHqtBBk3
Wt3AXa3gIJ0Mrohubz+jaZ7tcXBTfjK+KNeNZ3/ICeKVDd+4vinB39p3twtUVu3U
j0kkZTuiisumpM8FGK9GfvZESruoN3RoN/IEN9JlURvrF6Fk6F+7w+AM0gxULTJD
kZdYMiir2htndGSM17/ckgGe7Z+58JgCq/DzRNe4M6zj05GA5SzAl/4wl89aPUQG
XQoGdudBS02n9EmrIdIVJO2HaLFdVZUscehXPq0XRAR6UWCrstHtfd0m9XUokkaS
fYsUWB0MXSeEGO1Iiazpbcj4trDiFRPeQ9uIH0lZd55e0SkolB6y8kR8lNOfRVeq
dyzyxzhn6FZ6N0wQeB9Fsx+xey0jDLrNdN12CQfpwUn1vlEZmKcLkqDMdAF9mAh1
zzfc4LWrzDHEA7xznvvb/mSpjHWSx/0THWv3+lfYF+8zF4k9QlgGy+eCVtKHWhUn
qmMnyq0aZZt/bi36Q1qneB9C0Bx4LT98iZx8z1efCe24DjTAwij2lvxLCD0Sg++/
LmDvYHQWAM4jIZehzUarxuOXugGH94LVvEehsfSIoU5RxFNli60OPJ5/am7Jvn9K
FEkrEPKx92bx8HK4w6XEotReb9P5aZW8s7L//qtwrGv+3apcid61RSHEgimVRfJ4
w2wo4/026vQO0WNKMbSMZB0LlXkDcfUIUHIB3tD308owF4Zb1j0yu3RGpwFuXmjt
NVWX/YiP81OjS+Vt5EtU1DID7rIkcfua4/QAkI/GBKUSiqOlnHv3XsPyVBl9mH2t
pTf3U0BQFLeNLaSlsgNcPAS2WaFBP8AJzj2Iwr5pIj+KPiEOOdIEGcdYumVltsSA
i9cXQfi2v+qJMMtt80GblsMkrcoyNbshBhXWQviwej2nNOQN2wU/O97lJKMhwp+q
LdXhB6I2/RCvdCNW11AOXd121eFYETAQlLblePA1TzdpMkaDIQ72L3cHqIIOziPP
ykPA91UaRbtYzs+DYFToWO1N/bnB45sKxTcxqYg7o+2ScJ4p1AEPppWDbRudKsQu
qoLd0/MpgYIQKvUmq5mQBlHOtEvpLd3lQctCgc0468yUZ3EFk0SiJRXzn8fnVPJb
3FUqnCcvxr7xjU6H5c+MH2HGkwrE4rA6jgo3cV2XQTHUAY5cyhLMM9ZpDje/z2hG
YyQfgJwssxcpTNj3DqJayNp1oB0PuJ8wHxSYvau1r3jUuE5MQt8vWydFUaxrd+BB
ntFJhwI5b7OYv+O+wQK6WigNVZ6VYC1Av0R/aLqhBgMWQU4YZ0R2RvqV95psq8Dd
BOKHSI0Xs7OQN/KL7GwdYrtutQqWmok687yoQY6GZX4detQDWnxz9aZsfOaF7lfr
zQtjQuMk6MnK34Ser1df1BNWNWx2wAGScxMrVE+6gehUNarmnO8uAhUIXLXt3Yl2
DLnB+QnMdi3ofgYsdcqaUOle+Dz4a7Dw1+4ALK+5K9fQjQ11Wavz/9iEaWXQC1Vi
GOfc9hMqGf8H0NvzyU9w8o/soNXxbbLm3J3BdFN3B13LBva8kRGcnFcBPKuTqkz6
AUhOn9fijneKJZYfylYLeTiV5UAID/IJnDh0pok+ESOWM9XV4bKmDhA90uzh97JS
LHaaX9+snGShP5ndxJHCFO9p3yAQlVCeNrzs8v1/nM58/zVg8s2CAgyD11G9abTV
8BNdoBImGdVlYUcfXNxq+uX3DB9oSTEkZPtAnn5JL6eRQoFG/yMvW0LQSTjC5uyH
tG95zStsxybq8RicaD3tiS5PM8318V7xYswgtL5+5zrOY82A3izn5lkWnUNcdX/d
eQvpw+X3UPFyatGD8BE3Ku0ACgsW7Bo/UjLwaABcfDwkYiIpjteF8C/NdYYdVVML
Il/Owdc3/Ph1yeVhgRDw/oA3nZLqAY7bVVgv+tsuiQAI4os5zwI3XchoaAcgCzdO
0+rdRnhDQUkTy2rxoBj6GRZItA2Tumv39H5+gkxe0xakjE4fLgxuXxuNXqLViKnY
jq+yV1Wt3/xEHs07sOXSPkm9q99DbIyh9mCnOXH7oT3NMHFEPiv7YKcV7v0yQ+Lz
27g323cQPdh4fsfsOIzZ5LFN7zR5ZGGhlYtav5bPuy+EdzBzeheNpWkbgFEETobF
s4R07SM9LXko/zEJGbHyJ4ey5j2xFGoJ+enU/tp93Cc7NYWO7mQhlbvhZJV8aCEB
mvlPUQBqud9UoIaIR+ZcPV9j1HsjtzFQMw3aYL+DCC9B6dbyfU6WR0JiXrthwXOu
Y7KSxi5LQHaJIpOO69wBjYtiyI8d7u9iLML3xswrKNFot4Gy7U8kkOnG/IjF37qH
kQRn0OOtymG4tPeQQM5RSVrb5SOAomaGhZgkwbSJ5TenHfp3GZPSDj4cwc3RwD3C
rwbvOrOWfReTD9W3Df+GXVNG2yDexONfOTc+kw+K6j3fAro+UdgnN0elTebF5xJI
8TqzkIjfrnm7i5lRv97BltMZfhD4YwDjMB6qtLhcW5j2NM6x1vvgIDwu+vtxpLEw
T8+boE11BTzsZlkOjnt9Tnw6Em50xZQzXdwZPWR7UUTU5PKEWdbfBDLLmoyzsiUI
eNBWTRMeyd3PXbaJQqOo6EpB9ClqcLdZ0Q53fGtUw/LuwGbbAm2ego1E7geWqDUJ
bNyBF/gDCpmEjcerHY1GzQD0HSMdJlck/ShjBX3pQwaS657Ns4Q5BBb8jnHvAo2/
YeisfakF4p9rVCRjpTXPQGidSll0stna/KASDKq7MEX9BcEcvy8YgyGRTps6o/C2
esYy/v+VOL4iozt/4glNbzv6JgT/x7F0QXgW3qKmkHYKm1AUNTf/Xf5I0pDoNkyj
0Gie360atK9LLZp451IEbY2Afzqi7plEbTevGrdXHc63jjOorhwRE4uc8f/rkcfS
r+plHi0GodYKpHr87wqrx1jZ052ci/lG80eKQcRCV0Jy2ieXm5OsnQ0F9mLINklX
YOCRpxQ6VEPnjhDlAKOxa6PEghEe+iw3kd6xsH5QxAtdltcOEPWiB8l/D3WYBdhb
+6dZMjxKQFcLtypu8zwjauXhhyC9Dg6cSZ8m2vzMVHnCRRKOk/2/czuRld9dhLDG
QiylbDoEaecJq472QOkUN4tTRwYF8sm9xkI9PtJe2c8ZGUnEAk/Q/Z32qoEpNx9u
MQG7ziJ0Vsy0zblyxTPwpC05sRn4FpIEmbiR7Rxee1ckjKAZ+Yi20J0qOsLP7tMZ
p4QIKca7PBB7q5Vrt2Gf+zkHodTa+EUjOfE+p6PY5DV9ou43GS3lDSdeQIU7JAxo
UQBuJNaZ2v6WVAgCl8Hwly0FvH8qtFkfYaUstr+pT3H8fGEEX/IucYKzM2NAvWTL
KXg18SdluFFYTw02vK471SVkJS//3lZvISakt79yrs5i3RWbrp3J0pmODvdNK64l
Lj2ZuhHvb3ihQviPUsHBqX8KA56PBSvRTgrop7Gxql1nKHJOKWMmDvlwTHejEB1k
riFORcOQRf6xth7Gjx0N1dXRX519z3WTnEwvz6XzXYDjfqN0ft4+aXey+EfXAREF
6b+DGI3TSa4KVfoRX9dUg0FvojfzWiqGDRk9A4vUEJtfeoH/+8Ctglvhp46ZoA7U
VI40h0/9Jh50cnSZnwjRD/dfmheomjyI0ww6itUfEKYnb+w/TDGQPcbmUPciyjwB
3bUJy/dSe/pFLDm+upr1c3cyznwWyjlOm+cVkUoMEvga8fZesMV06F1TJZz2OSW7
m2dQ0gcec8L68EhB4f/Rnje9urXfdkziPnKkYamJ0hpw9kf9IAS73MnlKi4jtG4n
79krLwrfGmFlB1BhTjLjzgwJmpsl75AhlHffs808JzygEOC7BUEJe2bzormkodKN
Hc5enz/Kh016QFtS9XLQ+Q2T/g/Kl89RsSdWF+uAuZ2ff34/GHcuanrNmwm9kjHH
p9b24XpPFCZdsGpTGSIqPVf5G/UySV9p0HFfNVdbgEuM/6Pi1JSSLt5O0qfI4/++
EtOv1MkeSWrya7F0s4EtWzdyRHS+dFC5zDU7PAwYbodBaz7NT2/J1zxNkslrkwa7
r9FIxoWSpjpoJuahXF2Inh8RkfCFu2z/UfJJ3O/B8Xq/yrJeL6M2bAR8bN8FlIWy
f2gZSxP5J9n9VilZ5IGX+Ky8spz+WbOpK1rKAsy8dsdZ4CixvZrXAYnU/YzO2WCP
959IFkD67cavXElTEgKZ5geQ7poNQLYDz7RiVhjBTQ0IckS9ribcYO/Zr1e2+QzK
yW8ejnCDVPuLJSucTimI/aejcNHQrrLfIAnmvq9FclH2L0fs27wYSiNgMvLtCRsD
1fu3ewvld8wrt8pqr1s3wREmyPjAMSl6GPYOChi9mXCJwf7Jgq+M2K6VtEcClHTX
PuSdAHyeuo1/dezKr/J0fL6Qam7+b88krevovaysukd1zyVvXmh6seTMnPOLHh3u
jh3PjExhVpv1mXD9GwCWO4omOQPHKX1lUA8Vuo7pfeEmt9cOkpga84kxWgVmIHWj
KSJTM2VcwxAS8hy391WWsW/SZMNuKL4Wb46Pr3Z1lofs5FyyTAAyQz8T85wRvjK5
JJXPCX6h/xPKgCDFXyRTqyeE/mICD89kBuIpf4dx17/TWquObNrP0S7M+lPpnBOX
DNbtjnrhVeaA7Vh8hZU3wEOdmMbg3zTBmNut5L6CP9/jNFeN9JDGikdjH/syBdf3
C3fU1QJPw6meM/rmpzrts5vxvpnZ2H/5REgfG58p20Xh52cssFy3KbdPHbZwAgvf
nXRCwBRYARhOvTn3i3szI2S5s6t6U+m3MnTBoYSS5xSMi/re3V0w2Fa/LxUH0iue
r357TNb6alzOpph0kzVBM4/csxRMFcscGtk4OLQ4l8x5LQIY0rqHI220BeDMgpeN
LoBxcTxHsUINbHkMrFvgkE6RwMxuXex75fx6jlvjEeX8LsAWrdi6ipcDvUXTUD4N
hB50MEu2vuteS6/1BMn9BGL9s6mXq06s3Dgf/Yrs82ZxLBeGVCvIh82mqOLtPAbr
9ZIX/N/WYoM8rSfuQbF1/ZuhK+eWmaukSnvURmANmzWchyvyC2QrNpyICs7FmkKZ
zSjqPeCvpDbEl4scemX7KCAGkoyFZx5U9SFChRBtqoQEL+oGputZCq5D0IbvXdiX
Tj/+CzQZCm+5Cvjc3i/DAYTovfEBLByTQ/DL73n0mcc4AlLKIulgY/l2MW9K3BRc
NBeUka/gU/KTkPK1k0glNGH+krHONipicbkPPnh7mfVzAFTxFdmiT+x+gGOx1CWY
LXxb3MHQI6qCYX/6FWj8XU8nu+7J5k188zB1QCvTvT32nyG97OkYdpUlysjvAmJM
VeAMqW6V3M2VnJAHuzXn8Ws5m6wPTWjNXA2N7VuwpnxLM0saEL4cLyGAkeQcNuCq
1wJf2BYVibBOvyE5s0cyUmtRJO2AEEuDcORKBhFtvHp4GTrZk6sOtGZpmroyfRp8
TA8mzltHvN66V2NYhNtduCyebhrXH9PAj1xKCu3jkhrKQMjniPyL56owoeVBazZ2
d5p/HXpHFTwbw8/D6X56Ar1EcsRgypOV4q6OC+FB8IujRX31YaCt4cf6sJh6MPaz
fEAanXkriKEPdgT2v9bHveQVPzt5dWc/7gylwyfrWu1GajSOkA1YUSCAnN/gikam
qgDD6gVbluMFdtlRwZvHmPO+B0yt3Bvsvxbu1PZ9ZfIV6KXx9WkzgHpirv7PFrBa
3n3yT7ESgiq9Qz70sPbEeSy6l6uw0ug8zUG/2S5k/eYJs81KEltPQZWWcIH6aP/U
/b0AICWeS3ndM11y0Z701KRVTeHagpBEYKYJZUz7v05Lts/oVB4FBAWOJsvg1n19
NvG2HTJzEppxUVHInYk+9YYEPmV8Do8sqMc7PCnD3/JfhkfV8kXvAFEunb1jYt4A
VWNnimskH/NveF3RKjUbhWqURz9ktUSkf+UWmeo29uS6cXNf+04Lw6P3gYveauBR
eHL0txqnj0c9jUPRnLdW6Ys7d77M6zKD3Zctd/6FY32NjDnIKrqzLnK86nodlSoS
y3hj0UAvtf78v72yWpI2B+c5tr2FcH60eE9gzrf3o4FOZrPuyJO4tdFsUN81CHkv
Gic2IiUWSeWHV272Xs5UgegoZHoX6UPhHnaVLTejXuLxIZVFbDrQlkfhRZbQYzi4
fhH6J0uNcbdU/v8RhcngZbcv5SdiHk2i68my9+6A3e+wP9CHIhQ1klVm3K7CL21p
Ud/xUdLpjnbDtQh6BhhqtFeG69G64YLkjNOfj7gKW0W3Q+o3b3iBeZm9pA+fRxLE
Njss1hN66DwEBCmJkYdJDWNZyjP4zD05zsT4bOL6zLkfLa+BMZWV+Xif2JlAgwpj
RExcCi45yd9FdfE4+dI2IIrG6PRJulWURsQyFrkZoo+XDma2VE2zN/xWune3naCz
koQ2bVCFbbSeD1RE0bZGThyDCoKud4W3C4JgrZIeGijY/QshAQD4h8XkSfNeNF9O
02LwG0X8MyoprgH+SqMeoyg7wPC6etCPfSkqhIDuNwWaT1Blh1FDohTEAdh8vrEL
n/Nfjyk6ke+YbngphhIoFdRDqKUB2o4ow1G5xOGNhg8sqf4/2j9pHpuYzA3aCitW
Uu8VPB8y1B3pxAMy8G1xiSDzEKCp783xxd7HbvuaWaFLMRpHaqUNUAMurt7ufygs
KlA+IvOd1OoXO196vHY2qhf6YET0K/k0uAjfIxUrAbRpgUxoXGAVOl0K++4s2vrg
8P39l5jZtwL2HwkpKqPLbPIAeGRafg+GPGw8hVlpmlZh0ajivLw4wFNt+kwm0Gee
+cxr4fgCe9UAb36EsYCpkADk+k1636OeuGl2EDmH0EvUmnL9swOvMjJQrY/Vzs5j
rsh4/sAlGrGZB0f35AkX3/6EsyVLDw6z00fjuUKSTXc9AJkgOOkkj5jWSYoyIjf2
DkQPfW/1w0BPZv4O2tDSjEIG0eJIJ3PDX95NtOj+GSVWubc6/xXYLUMe2+2B8ftu
nJphG+DUkOtWMWytNC6+cQ9A5KFwrCoxtmwQx1aO1OO0CGFnAqatOkDY+Lv+oYPN
ynfinxcLIB30gpy6yWBtog+eDQknmKPsA831GbdYZlsVCR+iHNGB99lNT2YWX476
FZmafySoUro2pnBtIl2kJfzxkxtrorbtFMxb804L8mtzixyM8FAWOiSgiozlE9OI
5ZffVx05T8dTrMg6+RaSbij8FqsgM5ZZLgF1glKXf3uQXbKLmpqCWrp/YUeh0Bet
Q6AFLsKKFAcSUNdsHf8MbecIwAevtNqsiE9Tn8uh+//6YHqZTsXL5X9XBN9pP6iw
bWvPJk+O61FGmvKYCoO5nH+x3G4JDnaRFA2DDgLTUSBaa+TEFdiTZP9Qp3dDkq1C
pEtTXIoKXGyvLJp++AKBK+gzzvyLxNoNWVzGftHCPoWpIURL+GQ8GSPvl5jp7u/1
QorCY+stRUSwcZF88S6ktp3tmj4H+zcDjd3Itb/lQPYCNu13sMxgDJvmrTKKNQ1T
1CGrk7qboCy+lhvy/rmpH2fa9JPrfIvDrjX+U0oR8tqC/sCYF3knSSxIkpzvJ4zN
kLukWjMkJdAqkCxLhuXNZWUDMCJmTd6R4i70tf+0He2tuwq6aa629K7DWGZqBXl2
xGAhhKnwLcI12ND05/m0jMbtoDXPumZVWYo9qpVai3zlry3IF4B3UKCyjLDP9dtc
S+sv/G2wmCK7/UWjpmfnQLtcgWAIYFXkAJOJWaABhlPkj52juNR2blRmQy6iMZTC
yWVyw+M3OQEAZkaajuIZ1bjq0zWjp942oBXVQtVYwDnBm0zk2j5Abu1pCA/srPpF
l5DO8nTW6vsf+Y3W20kDl9ykMD3HqT4Ul9yAdlWa9sr//sYW0SIGvPXpaYW32HwH
g783gTIiDOgN1HiWWDVbIm2NpYSiBxCQodhtNtTH9doGtdJD+Ah/707Hik2Ehhns
WIcY+CLELB78nbcIGKrq89wFBo4E2kNgTO07ZqGrpLFfodfrB0OlmE+1l+rsFVgU
uT3iTcd0ho5aMpkJFlUTCLIahxtwZeb0I+DVU97snGeKQp4XtxeD4oDwV0HENneC
MuPhwe+Rv6zlr2mxfAAzFqBjx0wmnWd8T3K6XfzbotVfwh9cuEUwsZ7klQ/D9/uu
JNb1taqWdTEYz0Sa+aBkJwSTfOPqjKfoeeJJu7fYM+PY6CLTQhzFZdGJQv82udnf
9Krh0jScOHv0KUjXQe51pr1kZcUadkuZvhaE8ONIQp2GNusBxfeY2QvqAeT75Qhm
hH0aIIek2dD6kZJy25M0AH7z7s7dFwtmig1TfkR2aWfNMxwphoVMl+YMakkI3d5s
duz7h6A/hkl1Sgo3fCX2HJR1gh7VWgtXAt1GT5mlbLuAZljTvVXB38LA1y6oA36B
/p1WEC86UaNxKC7c4hzbWLC5Bip0hZl7uMBWDmQ/YdOPcPAXLF0TQ8Wl3aqGaPov
droqbFBMrPQ0WOqSun/shSRsUXPSLbkf5djopCYyp/O+HC+rP70+lWyClBziKtp9
XUNBzTsXRK+WgAR21T5hRmunavhWNsgI74NBQA4FuaYtjoKgUXDjym1/eOKzHc+7
zMOMEevOWBQjP8lsUAOtWSP+17gcD3BT1XNgeeytuhh4VAy2v755yo4OvqYkQrhH
J10loBZhfeh6AjqAHDF7+FbyP7FzCkzpWujOBq1E5NS0DPtlMaQpU6DUYd4qFUIJ
vUOIQ/GwbXN/zKj4eg7kcWqzBc780i7PD0UkRGgT7hCQcTHxH7lk2wbJFUboqn3X
DLTeFkQg1LXjg101YJCS/5EW1SJXP3iXF3NSHkTQbI4s3mQhMdYBmUbt3yOU8Yl/
1fmCksNEn51hzfNqOAdIah61ExlNWMVRp17GGKy+k+l/R0RVI59PiAMKDuiw+X1J
w0z3mRqfcvzXHvTJK8dkUjOgnrtxo2WPm+Ix9/UrNARnGtwhlrR8+8yqqK4232j4
tY00QdBaG/C9oZLe66gbQ+sAAjJwOoKbB2iNFMvlbKVVKF/+07inwIPgYyPiVTNV
w6KCRCoCNZBU/DpTn0JgKrjGz2OSkj4cUXZUZVU2EWReVaN/zSyRX6ttou+V7FgH
Ho3wBpMARv1YhfO8WKjkQD18vWJIibYkf2EQqvs1pJsmJryqivZZe6LMggJ4PBcn
UNeMH96L6iV2Jyijo5tiJo6qvW04y+MLejdHIztBm4npBqRvanMzh08Z1ZFcNkkE
JY+FS1ER1t8Z6r6SaDx5VGkezvMqexdyMC1A5fHFZ7/0+66axO8/sGAlxMtepnEX
yUjp/K9UyGAY8h3f0ZzmILQVdeZsBG0dk9gH3jl3jS+muxO0HSjHapJI3PpA2izL
aBrBK+tvE5KpqxfiB8W1kuUZFAcYNi8f41n7voVP/+ty8pVHK4TW43uFKL1LQain
ZoCiRwPHQpFvxyrrJq06an0n9qs1Xex/3aDveT/AWMf/Ye928lcGuS+ScaaoXwN8
6MpEDGCbKRvbOHMl1HCoCmPklbYotFN+ZUViuXOHFqohKmD7mwpyiBiQ/Sf41ifl
Pi83CovvEZsDC1cZdnQS8CD5gLD9iLJitnIl3YsaV0xvObOPYdkp+6/x5oDbD7Xc
Ld9s382a1jmIiiWouAFRTo3RMiRxgL1Cr2kESHVjO3yREasX3fLhCY6pwE8x/pRa
JEMIqBI/tgLgIYfbhCT5SQxPeQirGqpOX7LS3U6SbUs+v0gaTsuSNrydBCuhX0+6
dba6uVfqbYdhaRDSFuKV0HSYGW8wQQORy5nHh1SsG8vd7OojAErXjIkLQxTJPf0E
BE2TAckFKC8fftK1xlno55sriUbyfJFE939SxknItdODquRYgsTx8k53dzo6URnb
SO+2LJuZ1O6D+VXMbrSJhEvWHU0ytB3BN277l01mLChF/KugLhFEBF6jcfIMxek7
JKaSA9lsH26TNYcDqlnorcahjAGSWSYC3Q9wP86KTiSsi0ZFZyYNwKkfnblLQ4Pw
MK0tpH+tpXuTOuXNb+C/gv5siOXIkzmqozvI7/4bjzBdhweFqRtiRdlD/lEMm3l1
bxYHtwghiPKqXvws+woWf28V67gR6K1a3r1mBNMKQ7Sfk2p79dDvOyw8iJnVrT7L
Omx+FDwuhPlKDFWf+blDiiBbGBKN8n61+iz3EBz3xvtmtaPqdBpXvHJ4Y2HfXdrH
hm8501GnQC6soPhxFX2NG007PPQDy92QLlc5Paq3yr7pPFhbVIqgiBZBdpgyGXRT
g3UMEov11wG4JMC4OvBTP76piL/GuOFB01pypl+lkxmuWiBX45ijUvixoVZD5sUq
XKT2p383dJQstwQ57Tg2REtI9Kg+XbAJlmCApEOE5jRHPcdmGRoDNJXu2OlxIPTk
BjPeCJCDphYTpMFlt9fJxIj4S/lRLYM6cXzifoQjBzUIbZn2XcaUPNuvlrKF5iP/
GjAtJX1BEYzqRQ86X1ysb2tGH4pbuAb6dZ6U9pLIzLjkyBvvM1H1/ZUfOXsE+flD
qfXsQVtj1HEE8SH/T4ilN5MShcHUyQyHPBpBYdlTIhp3i/2Lyc5amGtinsyT91DM
5oSoJSOu9NqoHTyAfzJNMz4edXOLHd3qh2iX90Yh6kXAvopOT3gA4RNlJ+6ZGpiW
4B15RCel7szqjFsmqDCWWa++FyTJip/n3kSaiGZrpgcqvvQmygSG3F5zlgKE7v+x
uendedAWna+FCof4gQPBfwNPMmx1UgZ+iVsLy0SHugDE6upNf+8iahl4uUSCGjsm
PjHDSxK+zQN4zPfxjdfPmrWMhhksdA5I3ncKXVoH9bcXZGpY4wYuKR2saEC6Tvv4
4z5MhKQIxXmpH7ivLe0ij0Fi77J4dq9yCIH3GNPWYWZb4HfG+vzC7PhAmp8NRi8c
u+PrpS0E5VSLm93sFodmrRSumkBEWxWxAMJo6UbG1w5EW0Ijqee8Av3ts+BV7HFT
iHA4LNe8bkXauDCG5t32QZW6MvWNyO/yTStzjTRpQIgFpBdxkKRjIbleAeJjOn46
/j6knE/CqG5fKqs8xN1cKUBVmuX0XqsdQROYE1YQXmthPw5DxHppj69ohxewBC5T
YOtksc1ovoerVlOnZSFPtihS2Lxp+dR6kjUxVkis+PywyewHGhe+YBi1yww360Fb
hrIB7mxV8xwtjz5WL+rLxFg/4tA6cqJiArpb3vBgk8uWYA+YeVnl0y3fs4GXyiwD
gbcQ0i0COXJY0+l0uVrGAy67w0uCtJtYhJil5IW5U+C2Sf6KS5X1t+vmP1Vepsaj
vvPZ2MskWQcRpWI1YCIj5Gem8kkx/BbDHIlBG+RPddjNFcMTa7h5CfyuZq64YWkq
WTlOhiquWp8S43EmW+WGURxqXWKgE72q0e8pVhAlSNL9TQa8dyAoofXLc50rhRos
d053TAGwePxvkGAl55Inog+/k5lTTZyfeUQPPypOwm4n5IazzX4OEvSKZOMplZQb
btIL9OTD6MMiqKFFMRorMSUOw1xE9CA0JrIEzGlxm+VxAKgxRbicBObSCvtWIllg
+NsLrJAQDxkGUGQ9jUcXABJK07Z7CuHnsDg3dpE3bwJNPJs408ieM5Mf0IDy+fic
XH29lUA/gPPdhcoubka/0UXbAbALtTHtVxH7HFeZ1wyoqaAHtloTkYxuyDeJ/W/g
zIF2S+uzWnCqEgUHEDCILwiR+4VqY1lJhOc5YCg3REBVHxbNsROgHcYSUPd9og4U
xWwU83sp+xf7vYHhBamaINWWVlkwCLTIZLlL4vhQYDpbM8YcgWBH1qmsASDVcjvy
7jYg6qWHZpP6MFwhqZPhfVlVN1Z0YmYTAxW6quPT3NIX5bqPM/IFgfgVmNwFE9Ev
I22xg9iAJ+ujJ48EmSp1rBXhW/VMjNpGGxuzzZB1ERHdM1DdU1ripaIaqu9sb7vg
qsJMHk69EDAadKLgjGT84zyIOhA5E0MyHMsTLCGMeLtPDOUax5b65mV/LcYnnYWw
PIlxLmmzy/LF9cFYv0dQmiU8sSIMdSV+V487sOyGUZ2oVUM8CJdcrxV9CDoAOmhc
aq40t6uSFrkHes2E0+V/9XFGa6OrPYgoInOK6EZbp/4CjCuAgKMqT/X0h6+oGERO
wHf2QHch8FJrXBoJVemk01M0r5q8HOD1tgMj9BqCdYBM4cx6tcVw7pNyZYUklWTY
eBVNrzN6/KsJtGp6xJ6a7fNqHKZS+MR4+M3FY8AR83XnRTPlGJ36GJkfKplS2P9o
mvMyJgmvD/F9RHWM6l+5LTz/XKSoGgjflbM4o9uHNvdO+hfLUVJkboj1/bLYnaQ0
zQdVnupmCxGBb2YyjkXIwnZwUXc3c8or1njQUhNeNv3sbmlCzEP++61eQqGAH3u5
WpV3BT8EPA0jPl+aP5LvgAPDhdm0+APWxSXeQyA8uUkHLNADjElw0htnr6DApnsU
FgHofYgK1Zwt1hnZLv3bF7/gUqXPgURnM97BDTbB7GA+v4vJzi4zYUGlyGlnopur
8Jgpe3jX8mScumlE2seC2N2s8UCrmRAACfevMET/sJ9ZYxt/W4TQaiWhxzyVJy2o
KepLxjGbc1ziXs/419V/QEWXgslYLGOTi8mQ3n0aFM6vVdJQ4Wu5BLrfTwGPv4LC
E5cfu0ZuiCm99ETAa/KbaaXQUR4F9fK/p8eQncnDXV0SpEKA8J7e7lQ4McudWtgQ
i3TuVeBmBIZO302vBa3fECxNUJRWafu+E+X0DyQBsJwxfP2LsBZqKlTyJgiIfWUC
mipkMV817TpZdC9mU1TDLZbtk7LyEcKX5TsFEAoC3Drb2sA21b7d06mn5vzXuj5b
EITBcUoJ4Z4ISqPUIfLcHmPv/EF+tuwSMbP9J0LX8VpmEgd9DjiO7HXybHIXSmT3
uOG2YXp3OY7ztNzRMI9MiKLi+1TkX76Wm+eDnQnjU3VOADBaCeqK3GUis+5SksRV
LLL49o/TsFKHRUobNX1sOMNzIzoGKNCKNjl5cgHyBaKVN0s8nFyS9oJsDroilUiP
FRVPigliKWDTphDcHygeiDMbRLMYgrkJpljISc1KrMOZyCbxWxMtLiDDS3MxZ6++
iVv3daULSrqJhgzh3/KON9XC2d+16WBmKWX0hL3G20R+upCLuX4tXcuwwaVRdfyT
9/0WeqZxBjfmaVwbEr/L8vgaIplDr0H2Jer+o7d0z/SDDYiF9flso8CD8xkXirlm
mgTpIL/su6tHN7M3gTbuVc2eHn7rPodp9vNnL5Dsb2Jo/bm7oBx2BFAqDbSJbgtv
4sv/wgZWJIHdDocYrOt0UmzVAfD9o9pBTpRJGc4n33uEBGSwNorTSiEmTreBs+Po
NQ4i5/VDGAV8t4rRGsbk/2m/dmRNbY3yqj8IcO8mtx49Qv/53JnlrvP1GX6y9TXK
yhT/LWLIT7+psMcqVUX6jmUVvqA8CNtoBrZ8f8NdLY3BpIaL7pzXrKaHBy4Q7vHs
5zl3E1ZSxBarSJ0WScQmklXlqlQbpHUmmI3mUxlA1PAc2lDDfL+GQbNSt6ikI9Ht
ftksUBsb1uz/Zo42Ha22RqJFApE1ck3m9HiBGUj+DfHNRMeagnTXvkw3Ws+kbK7S
EnBdUn0q2b8Ms89cgRt9LWil2P2fRTdLkoK/BJQO8U2g7ULnOl1qq72SuasEzajj
6UaXFs37oFJ8hXJZDHzTm3GMzAAbns5c4qX7eDNFB8NgRyk+lI4LkzK4b9C6Xaoo
Ke04H/tvY1dd87Fw8d5lfcIBMNfj16ZbaVwoaXs9CQHr0FrV3ian6qPfUd7LYO0g
E0VfLBgvMHR5ePFNgyI6dRX+FS8DlDnti8Sk0GqK5V3xzlI2mMITRLsUz62lmz4T
3/hx52FUu57Rz8sIi61T74fUXoe0vNzvP82DsS2vzp3aKr0Dq+vv8DIFKBOn8IjW
YXj5ipzjQLW1yM+vuKcaPEvDoYjg7RdzMMviVf3B76oPUTLYIDNuMNyQ8LFxEaWl
vYPqnJ1N0NMRfAGrbM7vwg90q69hmiW7vys7jxILgtU3PLPAR28e7nCMUYdp5mq0
tS/FhgB1i8i5h3cHiOqfRKPsQpN1QP1X/NdWlz1CgwD5jUh/EpdsY4GUoy5PTHEA
7NXhh6S0xkj0NYm0t4oVuaxRHqQCXBULNSryCYGgc0XLootqVF8amEB5DDrv6+sF
MS57Wp9+gpQin+8jsjFh0xCnXE1/Y3W9s/vtcTdt9gzHp9978FJw0aLvGch1SVQt
ihA+JuZOS4AhgpVYZLQh1sQETKK/rLoINn7rf/1JFVltwtkAmH5g07FtMiK6jS+f
FC1LbIQuTwZ+CCxRGDKMUa2B/MBMLS232ow8l1EfIKJsvhabmQ498BHPbf5v3u1r
UqDq7Q70qcpNkZd4QVSDC9LgFMhRFYi/nFt9gD2vs2Z2bCrqYnsTQyz4h4DVuNGH
J932FX+G911fwgTq4B+O3Tps8yJhXwFG8jeBw+0LpIUE7L2u/URCwBC7mlTrnVCm
diPxug0f/HqwQAO0Mk7/DujJuex+sWj1qgXR45zFTOtMknYAvVltWUxJ7tkqOmEk
k+OvrEDWWmNg4GK4SEsSu2D60YX6UyvG0iDJNR43HuM3te/liODfY85YBB0iVk9l
xIUFwoZTw+D9TlbQPkgZ2XKmQmAo+5/svGz6V2D1wNkddJonEr8hgMO5338z4i4P
AyTE8FFwQgKTnWrzYl8Xm3+E4GEKBYk4WrcwngTIS4LON+SoRYbhmC0zghbY31Qv
6DxfcK5L/3enELJMkz8wAvzLpNZRDVTcdfYP7v67WtFz9KxBSeZaATYeNkj50B5T
s5KpR4sZP3jrvdJvyXYk6SMH+zXT1k8bVYFgW5h3ag2cH8AuteoIpl0SuxjEo1Ud
zscpLcJq3Hn6jj2b36KyXqPzHHJOskwg7ktU5VEFujSYgdoii9KRn4Jm9cDgJiWh
J13bZ9dX2QoroRmjcv2hb3xWCCdRNl7RD7DhrJ2csF2MRbR80mkXUvRgfid8o+rT
Xbg5AGTSjrL6KKnmGMsVCMb496rmfle4BNz3tdRTsAzzP2Oceu5DUWWFjyR5nT0e
K437Nm+YlTaQEd7v+Ear2KXYGDfFFqsiulmaBP1Hfy/esqc7MuM4d6XAjMZ2e//r
2ivRPZxrllnBctoi8nQ7C12hczhp3htMitwBQ9lnT90WL4sXXZpL+L/fkq8qkoK8
rKjaj2h08WtVcMlGOc4koSUYVTg4xAitaA3BOUs8MYOlcb1VuktUX91nRJbTWPNh
t53btccm22TeaL9Neoaq1WZBb9pc2TBiOE1P7JpZB79c6WqbvoFV3Ygv9zO+tSyE
muAPPueZcAqjubFh5p3tA8Q/bNtYiP1fXSUgZxjMhTd5HDHig4TsejPnhdT8IPH1
PjMGaVGRLP8VRZkrMUg8xMZPqJqb2j5px4r5YqVeBGwiNA9tncJRTBcFp/sbFxHb
UfIQ8UNcwQGXrXbxPK4HDP0lQs6s9Iv9YN9DZiuRW5csRhHv9ogubMYurIw4Qi1t
cHwpGSW4kJzw0Aotd1Kw2JJRE81otW70lVRnlSQPPiILB3LfNIvK5bZ8v9TQTd63
DNCuIXu6FlnFC9i0myLn2MJ79V2HwsbF38Nnv/2dVRkFrn/oB3QlKUl4cnoIpuB4
M23HuLyiaaE+/igFAGDU970sanUWwwe5QX6cyDRK0Q2biTUTGPMIjLArlaqfRtoN
CsrIcAUAzrQxUioOTGbUVKdRHekTFgbhM54XHNxdZv41S+5oUA+6xtZJGPzPwqjN
xrCmAA6hvHzmBFTby1zGo34g8AOStfAv4D2SwMZmidGKJqAHNGipM8VJdRN2m5ZJ
xxRmczNAVkBSndItCQp+C1Y8pWcfT7kuoz6j0HBN7/DdCHLXqpshxqv/4ndbtvpY
Iky4PCpOFKr+zYgTW8e3zmsSP04mcKXbZhLkazol/K38CUNY6SZ79AYCAFFX2wjL
6pGu/hVMOeYACshr6XxFnanUy5tSsHIb43bgteJkS1d5VCzvM44QlmiVP5Q6c089
9yroq9DWGX4oB9UlqRe83O/aDMRoin8Pg+sI01wA9K/cBx18CMFDi8QaSRIoOztY
ku+PxS0zwfJX3HR/DfckmYXNiXlUaUcAT0RZ5WWJ6A/o9viqOc5puTOjDiGhYTWa
no5ECK4PmysVx8JR3prh+ZyWqPM0nITJl5UDcSq4SLdL/aWW1gyqAj53Y5EXZlc8
egXlkMvhjIjG/U2rQAy1nvqcIOfVRUQkRB10C7lmzdlywuFrz7fxQXcVD1UoI7jS
voPegzRxGxExSF6oXfpq9RuBOJqbIxvMJFckm2jPAQu2OZmkP5ahnNvpLeiBQFaB
NKfcryUNoZGvC5fRVgqLwhTDVQBN+gb0WK3kQlw/UW+flLnwmVFdn+VZBLGqsxt5
ExFSH8xLi0u2Lebyrm7eG4ZX0qHf5rnayCRHTkEUhWFfd34ImFmNoX97uWnVdigw
hiOjckAjtW5LiXMzAG62+FgQeu5MTpjYXDBQhdsl5i3z9UFFaAt3Nn15hCeKBc+G
s1SwmJRJ5RF/IaZEpjminDnBM6o6/UeQEka4LXxpqTPxNkXhxl2MkarJlTBXh+Yv
1LVHdRxexcdaLt6yBZiGf/47KNONd+Xazp9J2VsWmDwsRgOXF3aftIiNbnGYkqkA
v6yWwiTKu9NLyvtfbvPhmqmXAopq69bgqd48SraTvL51E11SfsZgs0fTnP4wj5Kd
rUuMxOmutAE/YO69284h1HZMpgRcO84ttA/3WXPAXWcZmV4eqAcTfjDoTtns9Rn4
CzoyomEpAVrWqWJsQuX4+s5IN78P0ZPltXtZwy92Amv/Q2qSGBz7am/E8UyVk4iq
lCK4E0H/ME7aI70tqCxF2nWsWu9xB3WhGfgHvXak1FJitdCAP/LdUQcInhoft6yn
VCbXEzn0ezcv2WPFH3iR4Zc70EWPZ2Rvpb506lT/T5Tm5twuZ+jD9sCVT51D3wvA
KnIXPZRx+loPgrnfMuXq08uBDlbANxViLbfLbR2y6L9w48Y0YF2yBVciVC3qexht
r9C/I217X5N5yELSwqebxhe8rhoZUluHzGHnGOlYWjmS8KKL+kzPVNIwCIXiEx7b
s4DuWoFrZLaabFTQHY/bloRztcu8ktwivwYhSEhbsDoqxllPQxdc3rS6oK3k2Wvc
N8PwCXVh6Z57aLWgHdY02OtSkSsoBK30vEU5ifhyVl4zgF0dc0/TlYSt7LLVvn9F
6f3n5pyMsoxhjXvp80J7D0+Ne8oUv87Rr5m/99UPSvaI7ejh2DGwhRdf2xsYkGGS
l6n77z29gBnnMQuoSUUn9DO61f59QrzexOVPEgMK/F3yYf8acP3hlQqus9eWXVoO
5gRpZ+7CrVul1XDwfE6toBpQiRgISyiAzo52PPkfx4/zjkZDyjwpfUETSFPSDO1D
zoqVFOY+mlNXLkmWpvH9i4XLLp5ekpjxnSwdo8/6dYXDu57CAZ89ShE5ISjyJMl/
3krqmVlQ55ybQ8hicvafCuDXMI9D3cYbtSokzLqfaxzF1Tu47En1hg1xcXdsnNRe
rQ4OZ8lRyFNSv1VqVZQbMyQLOCCEclv37cl9Kzvr8UkxwovuOxPlyN+xNXng8/DD
K3FHmNT4TQ7DP0a+e4r8H4Iie+3MBJPYNudBjfz2jrwQefbDS5AYMAcFzT0dTDVE
F/vRAZ7Wv/NDhuYJ1WX9EVnUvqz5DLqSfRpmrTfpxWJCyav91yjAIGm/EX+wpBhN
X9QLTatl1T3Em5hJL5GZguSXcCLN/CDvupBh6oatn1y1qKS17OHizNcY6aEst5fd
fXgKcYtQGqFsj5ENb4qtzVE8bdqA1WxZf5ZIFgBdRt/jkIDj/UHuuA+B/bNC4ZZm
gDiz5ucG47YOzcu+iCiV6HAyLu50l8YbxWXHPQ6L7Dej/NXeVg2CN/w1xGUacC7H
LO1OJRl+M5r5QopsuaQPq1VkR6yVtH6/hB0ZucDhtdm+/h6jk21kgM7uLWm6f5eE
5h7LTWJEVLrT+PjhtBH3Ys0CSvTR6lHqcLd8ELCLhC3gIjeqrCIlhM2EFilJpShh
1YT5Qqez8iU+VzUhtwOBWQ/9UTFFWcaAV5Yct3fOp5B1lmB27/7sW1K7eH6c96ks
2UI1QR0hXA+KmhXIZF5BkdZZRe6fN9fMJrXn2YDq56tQH0KI4M+UVcE7OfeiJwAI
1QKd23fG45Bg4Yt6mNhKsmB05ZPKJSa6g1kMWnE7m6aXe+DSy7fU7biz5kQuvk9c
PXBtgobduTT7assD4VVvjUkHmT6uZc2aM99f8bOkDSET9Yc1VtFf++2yqWXKfYV0
lWoSdylki6A61Gq0epv7IC6zYUR4PwVHwBAT21125jeysF7vpSFEw5rZhlVZMnE0
UY6D2e8ahjjMmIjXtp2o0ifrkQZHxzUQ+3ZiSk3p1H0/mAIxzif7YhKVpIwJ7nfW
KYwd/mt6WPPfATphsksSH17RceDz5S6xb74yJlKPnKVFDh8SqLZGWspDSx/rTW/y
AXaIgtFIcE3IwPF+irRlvIYWVBtndL0k/rn7WI2JQ9r9nD6i2nQwMzMsvRIX7n69
EmjI1F+kAZ7aPWMoR0CNDD7sJ624NFLZFEAWy/59OEqyrympnaUn/HcNU87Dl6B2
vQz1PZsGTIP+wHV2QiUWSmq65syF2Ybg2q1JEoZPQ6Z6RGWg6V4eOyu2ntGJfNKG
ot7SH5eKAJuQ+HC2BHDZEdvVCftXid02ieRKdZf8KF5MsgdFYLJpxRfk0FXGeWLe
h7vuOUT4v8bHg8nDw+u6PImOpMiw3Dbo8OmnK1q57umnYovxvbCAZYSMpnhOIq+f
nOnM9k6M+F5XAM/E9UIhVr2m0oGAXTWqgsqVdpMsjeCPPhgLado43ZyZ6b4Bj1YN
8awSsTUW8QJhAF2HSlwtfbpDIcREiU2dJeThXTV4x5RTwbFCZjQ4Tjg/jHdvS6l1
Cvnw5XEw0Tw3onnCvqu2F1CcndxX9vxeUaBY7VVQMNNXR/seVF/4a4Zp0aDRNsvy
g0zq1jbH4c5L1u66FSTJHtqSnjXhLwrVZeuwD+fTVqX8j5PfosCJNwkLkWCG/sGp
EUUmMwqIYPu2hsCQcb9RecsN+emUPaN/LwtIG1edN1XPwJGzuJjDrMveDaNX+kU8
3VWcX497SwDNUJ/Yi+XiZT3FyezmJH02JVGwuHwYP1LrTsAgfXSwF3h4hcZirJjC
EQuHtcXH7NxZTUaoKkDFieCL9WXhYRwxf+jOwC9eHIpbJZLkrp8/Dyd+zYAb9UAs
T9Ipyw6+22IGctm2g/bi4DhkW9llRDv3IP3Dk0YwHLVb1pT9gZIRJmyOBXwWChi9
IcnsEL6jTEbt3+j0BJaBzqcvGCt/oJjFQGf52fffWIoJ2hBirViL0zIdzlHlcbKs
Jlyne6uIWGNHWC0sAuXVIEzFwafC0Fh+oDiMEGV0OPDLGnmD1hAxGYfMgYzcSh6k
CzA6qTFR9QxyWnR7UBbk3cUa27gkGvQ2g3Wgh9qLckl9Sz6s05olavrvDw2LQBQP
0aOuCm2qmOz5MD3qW0KvVRo/AGIEhVGhuUzBfJR21Qx7GrYTHCJvIdwudf9B5pkb
b5kDAF/tivBY5dESukwquAus5V1Y6tT+t8hTiPqQ7l/TfIK9Rkgc8SY5bq3aM/gq
JUYbimj7CQnb24AhFh3bDZAzuMneApJ3yO4nu65iPXKck/X68eL1l9xqHt8Q+Hnl
Vpqo8Sy31YIHGhjnYScaS3iEpcuIvgnDPk6WU/ENDtVR79EpfbppuC673Pvi6s+l
kUjUevDtEr/4B1AP9UdFgui/5rknlYTjxaNJFVWJh71K9VyYVWQiAC7pBjMyGO34
cXjlNYIYQETRoQNTsK9pHVTG3N2DqgNge52BEswKA2mF5Q91Z06dDD8U2ktKlXcW
Rq7K5YfLJHP5ebgCW4u/umZet5JmK1EG8xCAjfheu2pr4oBAjmFHJDaUYfHN2DNr
KMsnS0qg67g5iHABEqGj+MEbMt1xNBlN4tz4r0UbjxEz/dv0Uy/xbD7WNOvq1RdN
yG4CpVFNzhab5chsmKRNNlghcBmDnsuXkmI2ORNdb0Nx9seGrIW/s5HeM3El3O7n
C2avgRgWp2QY7WuZiyJCKljzDxLAgiSLLP/TLBZroDMaW9+u3kBReGMIM3Lj0/Ae
2qmq98ELiuXaVzlcUmgGSbcM2hLAIfvJxg8MdYW1Cz6Yxq1pZc23hi4KEeer8mmD
kYdZb7zlMMASXNoVdIynGyEaKELu5Z2mqt/A2My/rurbW9bKnrg+ul82M2Q1I4aO
3OEL4qdv25wmpmcS5vAds1EG5VXyiYXFiBiwzWRDrOYrTyrIyhCSjq3devnwzcOY
CVJ5y6cK6uy4KBbn0vhFn1csLtGtfRTHR3Rstn3aFTwOSc0f23dXMOlRiVJb3OA3
qJQZ5RSjKdUl9dfkR8Q27L4HtrpOb8//CdOQQSmUt1O7BsHeIgUWZ/DhqJjH0G6V
ZQfLdpffDGFkSMcXqP9ebhb2/KnDp4p+u53wuXk3+Lc6TSGbtFfvHYlz9YwVkIiQ
GI0cKrBwJKGbg7w+SjjNJANhWHk2zE25Q9fx3zDIbezJQCMmksR9SbLh91W9z5wU
E4ykRCvpQtcd8oc9zJqN4HHczKk26gRYbwcHGt4VvSiXQBeUcxMEVCeCZEiXQDWs
ZzcAbZ9Shev/xdyds0cmQlrKjuFZsQO5/Awe1EAvLqDZbaZ9O+vtmwA24LBeYH4x
DFtV6kvjknGfKYiiWRpN7IcBW6IivPnNmoq4391Wjp4y6rKb2I7EVJFQrBsiCuxQ
Heew/8dIZqmdgx4G6v4sbkkpirvvTNMVCoELeqiItEnSAetchz2FQ5WPPQyHekUO
wYjUD+EauGrgEzyUgmPX+PgVX07LvH852rvUYBtsBccv9boN9y5WKSqgSLuF3U/C
oABQbWAj82xwmTAUnui8G/vWRmwYpvpzq8+p7o94DOxaLD+Mt4TDNFUrh89wZWL8
r6bVg1TV6KgnpHBRxaXTnxVroBdaGYI5ekuqDlIiVcnf2as/V2SvnJ271XSjWaQi
EaIBjSegEr6Y/ean1Sr5elnepyA+CFEI8NIkt9M9qRsqEoaDmUyjZVnrxebIfhly
YWQvAvFtak4f8CfagcmCVtCns4Fp7Q7g5Yt7uj13ZRix0TZpYGo36djGhXsY+LSI
SQthXQPKEFu8Amw7/d7WOJL2XeXvtfWwIX03IwFVbnEBs4fcxPhD+oog23C8/kg3
/N/O5S/ttt6jcJsXh+EBJfvv2bX7qxR67FfbwBYQVFquEozJ7WDdCrJf16GUj2bm
hgoqRpG3H4Xm70zSIex+bXizVn046yiZ+QmIisQcUtWn72K3ODuyRadB4MiyYPXS
Atg8oSF2ROHmIMjd6bQsJ2F3G5RPT8zlGxfz0GsNy0Kq6bjuetTbFS0fdGIxM45J
0AiQ6B7Qzfll/bP8Zf9iXLG79murSEXhDqu2VhA+WSllCZ+t29tWzqQjfVHQy5mx
UjjYfmVqPfrjsRE/AvF+yFKuofntQhSJvAk0e16rPqgx21WGOa7cupcUVwRGZtTo
C20MH4d6+rb4PfzOFiMh3rNY4gpmaqcEtY538B4lKIOiwINAmUV4X7XA1ugL0Fmi
RE8QQyHVjwDWoMIHbGHBPXK4IHrpYJ3jPdA8Lsp9/qPRUFofEwD/zXqi8X76tTZz
LtugglABmE5+XMSm51tFoGZRP9BjEcr3HcG5f6+i0jmL7Ub1ATaqu2aFxW2sGe9f
tJSUPFJUx7U6Mx4ZB/bG6xWEFV/HgVJWiemQzFUzzGyWt0FX1/MhzD5DhasvByp/
epQvpUhiBGRUDpCngqYZYMW6cY47yYWbEX/qNWIlOy/+vtpgDLWJopETHyDRTE3O
7/UtKiYmuwkQbJp7bvL7OFvy2mdIfHDE6lhZq7VfKAnLzk2DG7EHi6IBCkUt45F8
R/L9NjKyYEIA0v2roHJI0meWto/4RBdC5Bb7yfPslXXN3qxDklOe7dyBhrgG0Axv
7gZkUDadDqMc/hMQWdRFMzxsvIsa21Lh/ZbfHFWs3BJgFCYSe/joNexkKnUuAsb/
P1Ea/YjCtMumBgFpCieXKMzhVYaWGHY478maSLziWoY9sDYD4QIfruNdlY8PbxS6
aJ2U9qRydkBb2xlzGBOCl/8PqWFvQwPGSnMmD9LfYuJ1iiRqoempy1Kuzh71zq4d
ChGeOM+inx9UjIuOkDzXgDsqbiAWaxSjqwLwWvfUkWOkFHbCSvp5L3zZ+kyyhkcW
jyl+K1r8yuS4o01boLg9DFn7F4tdqg50Lw/9n/IXfVOqEOy7BPWyKKJc3WgqlQXx
60xNvZMRApbrTxNvq/Pt0tacnnMJBRony2C5HGwBeBSFe2MPsbsiaEbGdkJKiu14
sIMQ4TiQyIXPg+vZmxVhND3j6szQ751F0sviVJ3x1LVzOPuUsfLKWCRIqya2G9nt
kMzm8qBNqxxa4Nc4ZZ33b9K0U/K0J3BUNKGjxNh7hFAP2EWvQElERRz3YcMTvfrE
v79LB92bD2lMDvvyMNe79QIos5rT6qTy1yIwjvI+0YBZnIfHr9i20vKYKBgUsdc+
zbHz3RUTuUqvEVg+6WHG1l+aqrWGbV/U3qWHWgsKkVJj5sL16rYcqrtB0T1RX37H
5EsAfC/e2UU1RtFV5MSM4Wvhu+ygOiPBxRYJ4vmCB3tXULdx8hmuI+XcyacwIVkH
x9rRdiWsm5BEsPmsAlrH39kx1o4+0u3gQzX+FrHYkNOkWC+7Auc9lsatOTxiJW7W
2WKsc4tQD5YSDlFONB9oiUt5nPOopcpnOWx1JGbBZ36Fwn/qxHtKSwAJAgJ7hMCF
uWaOlQn5GVvP2CJZoLn+9WydAUhmUCbVRDbc0+vZ5Q6BH8W1RYqZ4MctHAcyHVbj
D6oQDXT6sJD1I7cOwDErxiVuok0IBS87VWAWUjfMbkCnQC26GS4yRpNSnsOivwOs
cnOPOuEEME0/lQIuwMS2m/GXj7u8FJqCWmuYGyb9jJZMKoO7XUGstcsAKwqmZ+AP
/fauWDsm0Mhliu0/WfA7nogtHzkShM+7Na9ZabU5VjsNqU7Xwsm7Evsfvr1IPKwe
v3vfWNmrmdnxwnFE0DHr3+fMKZ0T54LAR+hvybzyr03GzePqvGZWLkpAisjBNuwP
A5UBICOp1AaRIPC73QKWne2YqvwK91/1CPPNhqqA9LVqXKSFc6iTdYJbp3I6Mph7
Vb8Jmwo63PHweg1F8Oz2d06LX9UCtt0cmySfvdoz9he/BoKpmo5QPptTpvWsbKZd
/Q7sEeOzSvg7JqgwVQcwQs+wJeZPHc4Bkt9GYiAx3O5Wtj1AB2POpgkdKCUmVIDb
X1STQLLTCG9bziwmBh8g4kmLehBC8Q1zPDa/xPFXSwpgdgyToXXdLWzSajPx6Lpj
Jl82GhSOwfWMz24Tnawfl7BGAs/m41ak5mReSh1DsFxdjE9CxcKLZQcrImcqb4Yu
QS7WBMw64MxhZmg7eKBxTzbHyf+NCIBPDK4tEXtWJTaa3wMzCmq0tTSnQQumx6eU
oF1rZ8BEUyTsnWSi5ybXMJHGFO8secWQZtb95uUn+xSnJvaYIaCL5/BW7ymTXEqN
T0QGG8wvrkTsEyEC3XDOQRMXTDDfmX/c0gPzLV4cfNVsivoqZ0Ii7UeO4fP92Wmf
PfF7k4e4KU0kw7eClO7PcKS5E5eXwUJ6fS2QqfXIi6HECR/pFsxsJLtc4Phuwa2O
aCkUG4/usMlSu1dLx7NDJiMhSVdF5KiHg0ZdEp5bFVdDfFeV9ZQcZZwZmHJ+W7qe
vy/zK1ApeVS9RFUuXs+RI7f54WczCuVxSVCvWqjLzgTuH5Rg3RtyRhNdRIOpOJ79
7rv1eTIp5bbh2FdgEcnInLyKFiWMI0wo8zDUkIbTgFgu+6AGFVqAB2dr8RTkAV/e
j2erQe7irKudiY6uoWoCqiw/lKrpPQUpLYym6Pqk9S3WtNjN901LBBQoEGqQ0zB2
y83gpP29N01arFr+qSqWBLqQEkxVkN3d4q4Z4LT0gD3dVuDtHX8mS0xCFbs4THLc
bAE35xveRBBCmAX0eR5Lwl9l2UbKqfh96AgprEoNtUY7oc1hfgh5UBSEngjW8IGq
EqyRSvMT1giDWV8KACIedOlmEWKstLT11tYUftW3z7TT1ewlAYWxkBt090/dP/UA
ObDZEFENPpEKOSUx35OF+QusZscC0RK6hAB0waNSOrDu9YkphmZFiNNMPqvtXrj0
xa3avKjU7UKph7MpRiI2QUQwc6S3MsY9USlW3WJh925Do5mJA0WntZAEpHGyza92
VI4kBBQUEUpl1Ue6Oaf9Yr/v/zDRmYtEgOVJwRW0S5hPFYvU+XIuoI20DzI3aMg/
RosM1mpnCOCpCHsshTDZiyPbXsJ2fPf+3rdNo9zNmuV04/sgpiTaM0pTQgiqNP1e
6An+1Ede2K9lB3g8pNLAGyj3EQsc2WvDuBoSyloow4UjG9G7WzvKTpFEi9RJA+7Q
M59qOgEezmBunZtj6ePPzPjJQ8eJyXmHniA9ljppMx7AD2tLXWrWy9/SEM5itbKk
lJE53JNX8w4fu60P7x5uZESt7zGvcRR4CtlRin7BACGvpqaFUsSjNzGxseUQHx3U
WvR4j36d1YY3p7NWcQy8IXFez2wI44rrCyVth2oarJS71J2CFdWexB8FS9lMChgZ
v6WGPyPc5oPXLra0NlcgwToZQXn/1djbrbnbPTHgqjISh5WuMnIa1WR6fBoYt6ma
RuuxQMmHFCorMSHcjepExqtNjTvsPkLbpd4pyN1Ps27vgOaN3DzbZbaRkttGC6aa
+QDYMjBtoLcL7wKHJp+XKfg3yiuGKUw0rr1RWa0vmU2C0JH09PF3HjBL3VUUHeYV
8r3N79vg4wdMsC3lielv8ENoStvVifPTty58t6x0z5Xr3iF0h2Nzp77C506UUQxE
C/vn8FWaCewYwr4X4RrajdDD8rnlcbCe5xMpAH4H/9ZMr/09fWceSEnmSSEJk/ZW
DBWmBh78ogNJuIQJL1LUscKD/3nS/1VJclgPOUC/stduZeQ2EZac+eNTMKmPr407
prg6Qs1JcT8QJSgtkMl9f70alqa01t5kxa4IDUowxoY5F3skLq/UO0enZG4oB35F
r/2kuHR5HC/hdsXfPR5X3gr8A1EmL4sC+msj+IRZV07kacEn/3U7n2wcJznbDW+d
7Ro5siBnptsevDDJNFsXGIU4WXU5FOfpZPhsp+qTvu0A9tC16BMmLeUMLCAudDW0
QpjM7YmX3z34ehgLHKIj6U1QJP3SbBV6DpLt/P8bTcB77mLB1AgV6pONx15inUIw
TApgTF6uX7WrC9AsNc7q8wHo6tFL2ghltQXa8Jaw1DYAPvrGLBrOLloZyo9Isy4d
gRz6wukHRx4HkZ3vbeBDr9eB2PyDxNNsDiUIe2V1jL6wsI+B3vvxxAdA6VstIGPl
woOgyK0w91oZ6UdUijUK53L1q+JE97QSAfa83GyLXPLxw30j+bW2ZdNjlBTAkyHu
uX4EDgA/WW3LJEQZLV0d0CJKMLJgu+nTcfIw8xrU6Ka8Pj+4Xx9yXcQU80our6TT
tlLxfiZNsmHB/r+6w1RENYDl4STEO/XtCMcnCPNatwV181OpEgD48sxcup/hwtHH
XhMFYeELmUAfjCSLAEwemZEPdOwSaREsN0nO9Yk9JoPhR9sEk87lQzZLo6iJ3DwK
IU+xobPnJcj8WNaXeOYDbq0rc0SlRT+uBccQmGf9MctMaFB4cqnmUuXN23Z/bnsW
yT8FU5+vcnnotLsMxySRG5Z3ZGh9MW99GcXWXPio6Xno89ktbqYUCkNHt3Xvwagp
2EAkYN49QxUqwF4pbfJi6w9ukbcw6uVNSKkEg665nrZPgE/9yaBhwRY1mi6EgV0j
qcIWjMVziwMyxnUI/6t/oxYV3OaaBcpHqMe1Doar0S4/nRPomieiDSCmDQDgnHzy
h9cMYVk15EkG4S6oa4D+ofeRuWGnFWNZZl3A7VmNNPD7Al/k77cCHTeOtBLXdrFy
MAVcLRL1vqto1bm6ZF37pDpPBnxi4xCRyhEOyfavQT2O2UVyjMiXhmH3lvDecogE
c3rKw+PJN/sD3Yyzice6aygerwrHNn0Cq7aTPKXIbBeZ94UKcoiKy5xrnbe7BLfT
tlciWsgOFvTfHHcM5ukkbyygX9i1z+Xss6FMwicONxSUX2A8mm+qdWzyUdpvdFdj
WiJttY9Yof9nZlO5RwSf94fQrdzy9FEi3Je7IaiciPb2OqpZ4vg/WEsfUa5ygoP1
sydaUO7+VxzYlRmxyJGBNmKeSitz/4a0dP70znHs5Y4KfbSgpVzjIOFiDCgMcORE
DcEnLCEWpc/ZOrxudA16NgLBqrLRZn3cdjkBDPNYj/TxZqPasojv4LrpGXpTXxGU
nUTkXpEVE1Xl6A1mH0Qbyiz3xJW+kKoqF5SrINqcVrc/1Pxfc+vatafQxO69sFi7
p49oYnslUNUESsqfdcl+c5Rv9J8Dajg2ngkbY1Yp/xhnLI3RR3flneAIQkvXlc0V
dtR+zcMPRQcqtGOY/tYUIJ3nvuJJTI7jg7HVHdJAPiR33CTRDBl4JUwvG36s1Q2Q
KY0DDxI2RRjvtnRvmYRw/0bCIx9SoUXbCxuxMtE5aTZGwEQ3aZEqqm5HI4O6oIuW
vTV9LLIBsR9Xo4/lejE/8HUcwGysRuvg+262li3lY723IlZfxsWR/sLpBU5mw2Hx
fN2kwkdsq0ruBf6QZj1tq36wDKD7UuSewEEz1ynPWt8ghchsz13xd1T10kLqlo/S
Wvmc3FxiB8fjsRT9uFXesK4MHkVN9Uo7Nbtfk3AX5MGF8Zq4BAVbRt0wYv6wLk1J
aLmHB0hg4A6r3eKwX+8l3F926YxdWuHFSGt2mxEzgTJZOl2kcDZGTV3ZRbeaRqXR
APmyudksbB7fRDN2GrijoDAqR6RPeFf9y+3tqbhxdkdfjo7Rm9uSnelTD/9an+wc
vvUDdqugFjB7EG2eFDdeJ63QkLsHJ0QfQqwVqBJ+rYpzpt73oymJwRS8X7Lwaf+f
n1+Ix4ZV8N5IYyDcBeUJ8iWv5XjfYXN92GKiANV+falLMGiLbxGWQ0lFhoD1WD7c
P6/rt+pwqBYZcpAlftfuVH0lwToBASQ+DFkRWwQQTA2q3l/YwdKcuYnRs5w9ioig
C0J6/9LqIvcCGRCsRY+t20dwshYeMK6coyEX2rOn9H8eW1tImYIM08B7mADjk6rW
oncdox0D89s+ZayUuT6L4PQ2YQ2VMFuxYRuuzPvVgjGMOhsN2X5dsQrdQSDx8slX
FAvX9QcWAsWhD9CzN13en0LpT+ElOwHYXczaZm+Vj02AJh2QY3x5Wc/JgNOmEEQf
ZK7sM6kSO4PkjZmkMhj1SgfffcmwtVsNM9Cswa6W4FH9/fnnl3g0vdEjCyhyF+lD
loMEPAWzO5sM6QqEMj7c6ds594mFuF+/meL2v4oZo8VBGFjW3wMZstHuS+lxoe7L
3tOxyOFsxmVuiNXZjDBKPAADNXQ+YnAY6gwKhi3wo2NnpfFo9FGTX2ySWBzjVMrf
xe7XoRp3X0o6akeE78PP4WmUrCxC6Xn6BW9NOxODCyPZD0qVzc20M++iv+Kwl1Gt
BmzzLWzzY/AXR0Hfsuuorp9gHQYwAyQXHXyx4OJHyPVQRodTIjj0UTGJOIFEK6rM
CGqeeRmmT2/qAeIQ4ecRQpPPtv1FNIk5jrV4E6suC8pZyNZ4c8kKxBXeODKRTkGL
v/n5oFDa0NulQIHT/Gr6D5zOw5fDWstM4rN6oBTFh4mjpLEkyw6qwzo1jpReK/6m
y40L5oGEji5rOpKlbd01hg5PHa+MXsGRE+gGjLT7nMP3KMF9IX/vvqMjlUlC3L9L
yaMRAJ3KJ7nvHeI1xBUKEixTxNmK0w5HgafGUbpIrXuBcsojxsnatm6r0KZXzIL2
BZWwUIXQrdVMY1zAcusR2/RNTYsKmwkYjyw751IYLDouMNgCvhLW09GOuSxqZXJG
8jxOlsAmu65CvRmPb2bKW3XkdciPa+he/zu5K/M9u1PEwbIPV81bBIuK6aBvYZtW
vBzUkun3V+qYa/Zd6djrETL2T7pzTEEqVqvgVGR6L5irHDaXUtOcjYhEC3Bk07G/
sj/E0SmjILZZ6jE77mig0dmsKdHut3neR8vxA149tIzose1mKyvfxfXbfVvLeyJ1
J8n5iWmFqYrOA2x8GHqh8N43U/OfO3jN/IvcfRGKqexCEHzUB6A3SjU9XVR2Qr76
Qlde9Hp18OOh5bqLkJ7OV7VDDdJQNViiHb36t1pDpwH9rH2BE6LISC6OS/94cnuC
2ItqtYCl4KQPyty88gOfPI3qjqrwC9VM0WA4wPuuroIzSEgMLrzvrJN37fvIOvm/
rubEmWI06dwHig/IaQsCPc3CKFHwI4uN4WoEdT6RAJ3+xPdesFSC4xRV+Q4d0QLS
4i22wss164gKw1CcbYCaFJN5wrJnDq/tD6dAFJuprlwk1OY7DKIesZBDhBMxjqD+
0TZViYV0fcK5YpRlaIhVIcua5KRHeaDJ3i9PrMZzUYuB5BBUMkJkbQ24ExVSRObw
NfsFU+utZ3Q1p+af/cnNqTB8nXGdmdPwFPeLdBdbEmqb6kdJcgSYmIDmPLfL5q/v
5YoJw86Dytzv2Q1EvMCnXlvAkfXisq9BEo6CDvj1e2KRzsj62YPLGF6VkTtsm/li
QH8i7jgJMkG8UBT9Ajpi0y69u4z8zGMN9NoeULC52GWwmKU7je6pZanSCLHflw20
ga4vT97r2/cUALI1iw44vHbXf5TvnWC8X+hPoODplNLONixdENJ2AiGk9pyXqsd/
/93vW+z+qTEKZ6GqKXU3GjrSHtMOlsdPDtCLOkzg6GjRxEYn6CiX7W1gD2BOWKC5
aLdscnflUDS1YTPDU5bW/DZ+DQ3DN3eJffPE7fd7fBeS+Hg6qsZFewSCkC73IBPg
TOGhNHnT4bfdmqK1FMcacsefbGp09K9XzL/+TNxhpIVj52n9mnq6u4qeuhfRz7+T
VU+BgBDy1Fj9i6SjdZ5inpywtqc5aREjXVeSpC1xpLj1WPnYHN+2AtBP3FbZHLTF
ObDawi6dEfZfL1KAlu2HcYDB+s31MgYwa6Qkh2U8IeY7yMHM1IgwykN9X8JnnFbB
JT7+iZK50VIH+YiKn28qC+P6dXpQvzH4JWMPxwn4JU48fvRE0KZRWA2cY5d0QxgF
v0VPa0pTPnbZXWveY3XzsMf6e3R83vNyYkh63XF8gLFTuS6mVoKyrGEa//nl5+fi
LNpffrHtpC6ZxozLMzhIkq/c5rHAIj5DWPKzlD1DXAUANvWE/Re7BnzFjKf6iYsr
jtlrXyf3yvOJjj9HyNdgfvvbuxgQkgLQ8kwF9Nd2ekr9bQ3rXFdkrQWYio2Xqnq6
JUwn3+8EArugt43gMCRlw02Pg1goFI8J/FzZAISHRlieA/hJC/f+KePogfbYNwtF
ndykH0RKBDIIw5BH+Ed/i4dmZLHHeSMZjoMv8qndwz30S+nYb4T2jgb7fkmaLO0f
Lo4MbdHHog49R2NQWqNzdRMH9YVu/GS9bv53LoeY6W+hd1/CGrbBvtmAuSBp+fpU
1ETYbVd28DleCfch+XVfdhNYH0fqbcdy6Za/CEcAkUk8ZdNhnpR7aSypGn+2E5ES
NzmRaa/UL0Vj8/AXvz+SpJPTGIddudEkjtiFrEwdi66noaHvGtWMNvQ7u0HDzxqp
obs5Jdy6o73wJUxl59rDftRaycDOu5ohe6izvshgkvk/oUIFRn8H7yUrKHZ4oJU6
W++vey50JjiCBpn4vgSUIDo+Oe32b9iRviy+YY7VUKguxS7TArQzYIVq2FPY9nL2
6G0+Uk8EuKpaVfsTBR57aDImqW4h/I1nw5rUmWk9EmU61GIZsX5zJB45EtZD+ACL
tg8j5+dKM9kWwPO17kaxssreWnwYSg7sXpnio+jTQ4Cf0aQqMKi3ovalGGPwUj9K
ytoL8tbjm5ItWaitiD3wLvHPsZqHXggvmyc4Hm4HfN+x8uGbybLkUXgr3dopJIPA
cLRdGBGoxE/AQU5BuFi53tW7aDcphra5Syf1KJA5sVTVw0DXZ140Pdc4JfOzdtiM
3I/WCujLusVnRwDRUG5Fu1VI3HYKB7JEqI8O559cGrzDLlaMEpRTyUohbSrgjvCk
7XYZcH33wa1gC1l/1hv0AQ1Z67ymAf63vYTQvDlrDGVK/tHKKmmGzzXs7vvdXkb0
2QZyErE/K/xsp76gUNHeOIDiNk2KaNuD/371SInNhIKpSpXUO2hyyBCJs2k9Hmn2
pda1AtLIPh5wUjMvJv5l9ZYVs6fLnjEePqXUYltdkAxrkwviFSMF8r2+tXkQfMi+
eIb2OP6ICxSWgLnQ3Hh/u6yrluJ8Ha3gz5Spi6UOdHlZWBVxhlUfag+W4QWgQmz7
0LOyvzuDQYhOGFqFgcCnxFbyn3naKLQ5KrpRFLj2jC5grhey/KOK5P2mIXIpHfVj
7vqvpGwGO8J6Zimv3L4I7YDioV0189UmHp57xbUrZvLnANsr3KPrsasCTZ29KdnQ
AEC+6DorlR+xADCTJyQ+fRserScQsNVPNkhzovD7OpCurtK2xNwTkhQYpuLcZsJy
hrk7IQntwAOPKJJielcw+giGlPNlSQgVaCKfFXZVpxramcnssBHzzC8bBNjfPP5I
Z+p9QiEpzOiCJoZneQY0ROKglX5vWMLbkp/d4ncdp6a7eAx1M+5ISDA49jKjDYMe
PBsQ4fw9WtqU9XEmtDOCDSy6ah/FcXGM7mZebEDAHQZsZgomTTc3Y9VGQo5IHTm+
wNlIk+0DHdimLeM0YRwORVtZGRNbp+MR+w7nIsl7dCqLHCSS6iVSnqYiwrfSyV9v
HRPpQh58WdNAuehgw/BXTi4Uew0LdGYM3dTMEIPVbT+sgV7nfBoLlK+X3FTConaz
7cT6gCI2UcXyUGSvTQynVTC6aRO+lNP0agGco+rTVDmXnyQXBdqlMgasKFOa9C1y
iaeN2uoEFbkJOq9rfWjQwH1GjmH6UTlDSrFtp59cW9zoxZXXP1WmwE2hflEEaA2D
VeBA70RCkKBpJpohfKeczKmZan7r4Y0k3j12Zo3Q7Al3t1tXsAv9/tw34rCvaEj4
61in0ibM/NnezQrkeMtnqqJOW43cFZk+aViv5AM8QPPhh/QB8n7d7ucogKNhb4wF
PvxFZSnNq2jTCnu/YyiMiBFz9gwbQtuN4a4Lo5iTA9d91CD79vYW2kWc033nyx+u
gygCiwtwM+VomJtFXKVhZZ3UCl/zjXQnIGfj46EgfpjDAhDpUzIPFXvxgTZHPso9
vgllXP/733bbc3w2ztWd1tIzUoCUc0VJqv4rYfkHXdTtxiFv3fCY0xQKbFDF3dQC
moO+TQn/d3+Pc9grwzGWWHq10qlKMZG8vJt7a7apX/7spvQflKLOl/DCjrv6t4Ke
BCTg82YjCQEtvzvB6GPRNJHxvDjbbCBTwEg+aSSej5YpX8a4jXVUmk0bCs3gQEFc
ayId3+HQy2U4i4rpbFWqA9S+ks7sb8CpQFGP8lgXqxZ10wg8Iu84N7Kx2bBp8v/V
4yjQtvC5aM1G+w9zP95A/d2itlCsu9/6ymutRjyDCGu434iETU3CvhxrIzQGmwqi
Z2HVW4iEUQiChlTfRuBW819nzrlbRzFtxa1WKyT1FLLlBdiEhfzHoQhDXyilfqTa
g+bloFFlRIptYq/A/uSEI2fSk7lsiHkBJeG84oVwnsWUJUBYF6018p6YPbhmaofK
tKvxNP3ToXo9CeHfv89ptq+t1zb/q42UZhU8GM5yh67X1Ucfkv7L84Zp5I1DnUCp
/QZAU/Xje0SKjVwh1ae4MUjza7Jy0/hIMxEc2iwJqvO2xgyPUl9Syg0Egj27CyCQ
DAX2tFjYDvmtZJzNyOCDcYEgPz7uTGw+baIwx0PSK/C1k6yEjYGnOAyp1d7VXYZZ
C4lmkswpkbo+OnPfPCHEfNvXlxuQISmcJlUdA4P6CVUFoibakjo14jMbxa7W713f
R++olkXWAdQ09PEflz3tNV1q2HzT0bvsZe03YV+miaIdBH4I6EtYcdVoiPaX4FQG
bszGRP3Kb8kvkrq+7/ot69/6zP3J0FB9hFNwpatyNv/fbCiwCXYiOjOBPGn2dIKx
2KRBvoZ3vDjQM4AWdpFIuEtOVWUIcPzKkvatTWLCL9XJvVJFWmthsQkP956FSCgD
f/4ef50E/H5egN+GJUUu6zeN1yRJ6V9LVrgS3euy0dKX7XCv+7MSQhQUGooHkm3s
KSJjgjnjJex9U46kjyClLijQX7vR5IQYSl4czyjo1GJBQVFumRdMJ0mnnb4HwWpd
dXtA6nugjTWN7ebsXqqovPO+sOM07VvcUFAIAVct1B7OSQRHLwQi+nEMzB9xFCx3
+1MWk7DebOrX54ulwgZ+A8gHjOhzJNkHQMlu9bJuQNgdto0bRVLDqTfB8x6Yu4cb
kZMXcB6ZtNd8YZzpYFI+ejL+jp//gZpIDqh3sMjEMLIU3l6LvuaZXHiyaaXRz93P
sPz03dykty5spBF9Di9eBWplXyPz8kHOMojO0Sd4YHRcH9/SQveuwHS3RP+HuQ0i
BqqGW2xFFIUt47we/XQPsHCOewNvGXrxnexgP8xJA9w1VOLhnQKiH93jcNv/mOB2
sDZn7EYK09cOV4wr6G32+V4u0hV/NlLTL2rM4/DQV4dmSEGXlrnf88AR0qrbfNsL
3apFEu7FreW2yHX953ulW+hW/JS2PDmTbpEGEnl+GU2qmsyUPDXIc2Ixn4rQr6ee
0O2LUggh6pcHFhAaCVzpmOpGLcE3Jv+smMSv+eYFqLDa6FW8mgZON5WuasikXrgL
eXlnzjChl4XWcu/XQ8jjKzF27/aFetWXR8DI/UTAANL7RaPWpFxY41vg+P+XHoVc
AZuoOUWLrJb7f9j4rLkciY8hWEkAZuEy+zhpl+ZRgAJKo0O2qzW1Q8NXV8+rYwVj
csyY2Mq8t3ED+8sUzMTYtdWpIOQy8ZwAXIhXKM2Nbw1PzC2LD4zPOh2iSogAqq+0
fRA6dkpi7jXoQpMv7wXmWBw2zGtMg4iQulzN/1LPdyefkAgg9AB+3WiPWxIjvfMM
TjubZfdn+7WoN360Du9Gane29asM0aTVj/ynjx0i/wEfjWuy0HhhCFgO7YSwhykA
t3tWjJK0xSkzmlH3Uj8YNsO4HOLNFEoq7Xb/7bgAZsDw11blP9fACE9p0cS99UID
ozoLeaMAU/kS+xEhO6pSwxumQM8nZUG/4ggWnsIdQ4sE/fibR7bM1NocBtnm86sX
tnaAoqqwDD1R0ZoHiSvv8dqoBjYIGgrBdNm/GYx/QFdkaWBI7zn1q1mkM5NGCXk+
Ta0RvpJyehFdnl1ofuPDh87sICWUR2+/A3Br/K2Z6BJ3CM7fVryAKhECYx7fOdPg
2agtZWzefwvJUCo1ctnKkIHeXu2cS/f/CPasaWqbXyl7PBrEvx3Ujg6ctqxGyKKR
tHchG9K36gLzEkuRk8dbi69bVuB2MhQEW1B2tNEr0wbxlFgwCxpHRRvab/PLwGTi
lgkoxYmVWfjBIGnIRmZ3xZYTrBaeLki7lsxiXzr7vv6+vRuchrBnWVoNprTXURRM
z2Zs4aGDx4V7ZSQ8XjA5Z9XgM/CMNurM5u87rxxb7kx53OGyj5DbFP7sypj6xLI3
EtFBT1FK5+CyMxBDH7C/n8R3Em2k3xF8+Y89yIRjKmY2XuRaHyhg7xLa9AIGNOr0
niM0jAkaa6g6OVin30uPiIGSq1D1/XBZ9t/cjl4G13OPO3zLrIIz4yT3RGJ89o/J
7s+P6TkYUVlz22zpIvrrM0PxhJTV4MZs1Fn4jY8AKpCkW4K4tGAiYLBGQ9apczlz
80HkjP4Ru28xXuEBlmkE7bCMOhvbikDdbWg2i7bmT4ElAiEUYM6LceSwbpehE62w
JOR2kCJs1mxW3HsbDTY96UFXQ4vDiW4uIWZhlu+z0I8PcHG3XtvsRSLSvCVdFF7B
b+N7TPZXj2kT20sQq/QrodPDZyjGdNnA6e999oK6hPe1TSTfM1AP7V3jEGblUtQ7
XHixEfhE0sMXFd3IXz1cxEq3kqszsCL2PK5cwkDL03tNu3kCGYjByyrNmgdd0akl
07Tl2ocxEcG1I/EQuha9koejgfd4UCdf1zaNYG9B/7WL8+yeHpKqwTEkKp8nha8v
sXI++n6UdxL0fPmE21ztuEYxQjYhU1yiPDf0hkE6jya1uo+TG8sEM2AL6Nx8/vW6
vz9FqgMNN/MypjiUXYyAb8vuVC8xuFof8dGlHSCNvmdp9VuN3g1daYSw5l/8QFRV
DQOYDreB3RV7fG/yqD9Nfqum+BYDIefaIVuNEgPgn23HKJb6gerrvhQnBp6xYwWn
A1D1CQmpviNxF1Ya4N/OeBf408HUY5vsDCRNz04BBpfajCS/qR/qyz4dl6V3He/R
/qIdOZxBwoeJWGywVrIc2oWJNJMKsiEz8i67rpGW48HDyOEeY0LuoD0na3PtmWOU
8fSlxO+ewX82CJ+u8W3GLdDN6JJGc7iZ26li//FaJketZhTPntwuUyyNTnJ9iOE4
xsTrRtVzLdemKotW9OyaGcUAd1G1rSkSPLVsxcGodBaljHyJHN++h/w5pmJwAi5C
3jJip7XavhDS7kseSJ22ftEc+kt2b7ohMX/HJDsGffuoX/Ww9QfldjZbtJpANt1D
58frFCVCV0DDcOmnODIQlR+GY8nQGgs1XOxTfT2lhjglmg02/ov4D4qlWBkrvhzP
WdaT+VHvwjhTnrrbX4S+EH4BMYK/0OurHEyQ0FBcEiQyxbGqWuJvab3qsom45TC8
MRv4qjET+CFPOGVdszj6zlD94xRuH0/7aHIY7AIxRRt4eZnl8yDd+xGZsdyL5cOi
H3/3jPRwDyFFIlQe80paPrx2nIJADAiyeNLt+nJE9oEC6CzGiwIVHRUelcIW196S
YD1wj48ksQA58N09CXnlUTgX+hmJQ6EQbp8dKRf/AooOtzERAFZd5DvXpT7i085H
55dpy2oGAqSpSJM2hY9gnNCX+UbA7IKtXRZ+PVTzH1jO6K3v7DB28J5YWHwV3cmS
g3KL3rvd+J0yT9bDzsXiGIUKwMAURNYMbI05AXVDYL9ApfyNUqunOnDZ07/7nAKW
rKQ/w+5yba8A/49+yw9kE+HZCWSRycTv/qgD/civUaAjZY3/SesFlUuKJ64yKrAr
238P4ApzxC7QgQaF4zzZ7HbTfCS0NewiCi3omYz97CYFmh64zBqK9d0Aa/tm1IBg
rr9eZ+cFg8n4tzMUIFNCfuaDBP7HN6q1M74Y0ERC8R6NAvgmo2pc0uCpH4GMLRXS
H6ONlaT8yMpvKegqxqshcYpGX9heziRCx/q2N9xtg3oZuiO+jXmNxo1rxkRMBQKb
83fwYBJF6qEgIkrPOVeFjhdXjPcAq82I+qPq9Avp0p/YV+X5YmaE355zOpAf7lX8
LKZyb1yYfIwn0wezGE9sJ8yLXv/r5DRc6FDrscyXL8rzLyhpVenSAuGE/uk4iOmF
x8bdEljdI7NIO4imyugd/OpoYiKzEZ5nT9neDSet/s4US3uQ74J/XEm4ax2nRBeq
BUiHTJhKaMQprVEdKj1R8dbdbWOoB+/+Sfw2fnEWm486ATkGkrHRN6/MQk6E5gbp
Y67mURucrV7pxz6rTQ3+61qnkOwE6AKd2C/azTNAdVw5TOqnB4WEHfSlhFMhMVaO
Tmdqla0+wGIE8UOyYv81/6MgyWnRY1ad3jHhyTtgZ7YNckFUNOFaYmb6FcZN06Pj
lIS+qyOXqcdiyoK5Ww095FnyP9TrpAhvcXlgxincTPj/lFnWULZN8J316HVp/ZyC
444tSJ/igqomha1EfAQxcCBQQP7YThLIB3OrIWJy8FaL2Z8IRQKalIsCnT5aUFTy
2+Olj9AJN+3t4MK5CIXoOeCrsYUTb/G2lJvHml7W49XqAQ/82sE9i9LARNi9I1Hw
3vI97PLWKvF6OyA2uCrMeG5E8sFBsWUZhjgNYGu43mz5WSl4U3TWiCbCjWl20mRa
EztkxnofDVQlmYhyn85OJKzQTKE8wcoDmTERKWhgOz/5SutOY8kBNtDZyQOuOYMZ
LZQyrfONRxcYJpCvQGV1c1f+Lzr/b8XUNZCdS4hBKYfAoNCnnNBkNGnsSUYyjYeQ
vdqz6cl5+nabL5/I4sXWccxT2mzgT0h024Rsn2pErgTbN7+l3jPPwi79v+/t5IO9
o+9MG1weF2aRBFl+tOEhiTzGfC4GcE9jupXD+UdoK1e/NV9Dya7NLpMe/hWIP8H8
8Mn9DL15SuZx6DHG54ivTyrGzF1sGqIhkASm23EiAXHVb39tMDvhqPG4HF2af2Du
F2vc8sAQ4vPeprwPak7crJEhkVR6Y1VWszyR2serN5vNpW1X2VcMgbA13wbkDiZc
PSJRSAeJJaer8pxlQXwHeTzc4Ho2XxLCSRsSichHVhXmCwEE/W4J8ZWwVUQEeMh5
/lINYo6Attt3dZhc6XjhSdHws7QuGHOTE86B/dWUau3ANOuO2Ug0pEclbPFx8+jT
cDvoBER1tJjn6exWd4UzKdF1KoFG1EtkwMjiNF80+WbqVCUKc6jSrLUoWvCq4dA5
3x9tyXvkFGEPFufZHWFW9eBmg7uFObO/sIFx77U+xdCNJvKgB2UH/E6aeRDjLs9L
3kgOHIB4aJX4WqurNFljRyHJv9z21ipi8N+TN3dPheBDRp7dLKsTqLhnuoGROYrc
alBAfACwnSX/oePz+3lpN917wkt1DhOFmDwWYnm7NcfB8AcD2Hj2bo72Mvig+BuP
Cp8w9LYzBQUuXxx1xXr3NzZZq8ildsnLP19l7q/31cqpg6ire9vrjznyYWK5iccI
2FWWSNu/vjJ+ScZaps0VObNMmBwANdjcgzULDWTUkNI1VnQDOfVS6gNfRmr7nqoO
eQPPNydWB9lx3mbUBk0SV991TgqJ7oI7MEvn91l/uo5NNqNTS2y31F/p9kdABfhS
J9JIjca6eptAQaMOhs+3DNJ6iu8ZI8Q/HvAbD6V/0Yy2UtznVeWGQ1DOeTMr44pX
1K3DVtfCJDh1OAt2Ti0Du2vLajuaMsA3VFzDvFlHg8v/uWIFwkwx0n0fhGYov7zW
bgNPtwsZr8WziBYgZmApvfLwJjUUdRfWURryqyuGjSBKGTpCuOZ2nV4Z6kUAQVsQ
EzDrL1Mi0NS4BgrIP9nQOCyJDipvJrj+ZENjggSgnoc9EyD6CzhP9QhhkZo+6foj
GQpE6eNPb3LcjcsfslVLc2YrwI7YwHedNb6VbC0MLtqcmuWrlBCYTjs4COPhXlRO
bK+PJdfzrPS0viTT/58FU/UbBpsNocN3VcjMxmifwmfU/ksObsJDBaKFf/N5BmyH
XCE2/uKImen/WR40z0mowNBFZc7fOojzoEnZ00QcEPgJ/2PZItsXMjBOnhh88l3p
CbQfwl8kFRQ2sZFpyw2SpQ1qRJAHjpbTo+u5RbnzPLmefw6+D4PXS9kCWAFlVisC
EB42m2rHZ5QGKjgcBMyjUTTRSlW3GgR3nBn4Gq/67gFBp2ZNhsF1pKDFWxuBRPkq
whTz/DnlJ7wuQlTagHkvGbAaxIWTCo+bTQSWMCGNKFweeUoQd0nZBhTz7zkWXtbD
7T8Po5Ll5BoS5iD5eGeIEM+lo8zV4/Ja8vK5tYeEvria3XRjbXgcuFql6UtDBqhl
+uy0KZQsyeufo2656pw5w2dejyxiKRpExKG9cL1O7/9vSEjycEtssioFROmTbU7K
iwAHgMl/zjgHOJ87eTNTA2M8ybxPBA1Auw1m8NWJFJ1D8YtU4sbsdKlTsdEWevKM
2YJwUGkeCDy50hOmffrrfw9Ap+WFtyRV30f/HY+iMESYbV8NknM8TT+sMkW9VS45
O1NSA8f1bdCl+AHh55XKlO24Pkx0IrEOgqFmPNYIVwAwj6IrQQny9TGbH7poQXiq
uQjLGfxdRZ4peGAaobAwR8qnvqKg6s5Sc2t9wjH8B4AuOVdsDW1vgqb//QNcWYUk
QSJKXTkop33kBdMM5zyJ7m6XkmFkigmsGGMud7sImkN/5DAg3p1SiNTs1xNP1dlm
9RzS01RjfGdGw4XDpDxJ8HBC/lsPFZKtPdNmuy2kHbqke7G9LcUGjF4Cnl3gRN0+
Et0jds+w1Me3l5RUh2GXipGJ5hjtak6dOCDjmA+wgD7GuGfbN/QKgme9GhWcazLG
bvexPzJBYcreLJVGCUpDpoQm01TpMtQSapwJeuFCqrUj6e+TCFLRqUS38xyJScun
mqX3N0RkCnrOjq4Hv+VBf9BlFWh30PNVuklcj5C/pEkv8TcauFAaKDWdWUHbpGx5
dtmAdK4QYlAScfwKjQtSuaslCox/1PblszQdqfM3jJ3AD1JNITU8E+RVFYdbngEu
aLqmPk2wEFiGmnoe5Fm4cOLNOJHlu3AX4Zud4Hi5FWI2ira9h5wugkpmINTYVFeo
YHd1v/zIQFTQg4GxoDkTQPRIkaD6eQLPU9qsMKemAGCzjncUVkQTzoo+BhN9XmCh
7qlhjXZkIlfTThsqXPjzp+3KsgxDeUf44RS9C9Aev7LzIO/iw0CrbijFLi3F2ImC
ZNAzs9ZdVuxMJG9ssedOAPqe2Cl1icK/mJpeqACuLBFQ/0NU6ruFL5Oh46TbhKCj
O3LVnzGWLum/YEr8sXZHsbVTmF4GvR4IW0yDunXWs4AkDu1zsQ3FREsRhyC1DPEp
4kfYXgt4pp1fAeN8A+bJeyss3fVKtRL4mvJF8tkn/qeOBeBhEwR42sKIFXeq9YXK
gwaVdO2wAnx6peiGmhgznFUo9TQHlRNOCk164M01D8gNVJeU8w64oRe9/P5WMxSh
6fCaYdD7BEfgbyZC+P70NQLPaX4O88Ta2qTwNkUhn+9n4VT3+ilZwf92T7PYkzdO
qGpY6Nsq6rTmPJfBRTB/YTJEb+MAjF4jdTVc8gfAUicLHD1s9jCSSDJepKptp9t7
3yX/j4tb1cEMW7xMcyQXC/NLDyKv3Se85NeVGCN65HVHzTCYApPj+LIgsiBCOM3/
qiP3n5pYfAwUczhuVB5aUSTxS7sgyQeU3kI9sjeF79YDdD+kZQsZ235bnsI5qo6T
LdCj+WTo67zN64jWBUs5ejRXdGn0vSIxaozitwBCTrAJ4plLIZVX9ofEUW9Atp/L
yoILUFQglu6GrM+ioaGrJQP0fEzt8kJAY3Cm+uBCMpLsCsUDWBIsyqr+Vp8X6VFb
YkRMAhzdM4BpaGFHPlPH2iSTbR8rdJ8AL3N0nM/MEqkCba/g68Eb8mP1wiDTlSJ5
GJfh6qXpsdN+tPZlPj4Im3cUhx6pTc0bOqzijJwy3gg7U3HxB5L44PUgtCnMAtR2
0E+IHzbIY5o5k75ki7Sxvo9BvBylG843OCdE1yALeERfQfv2CIVn6AeIcl7Oyhoy
651uh/qfzmlC3alJ/diUYwvTePn7kPF5MrdifBRX6qRkmyUJ3PHjvOot0KAUgLa2
W8IR+ppQ6ZAh7c82ibNXDap9upsqZYDfpjgc2Z7E7ZVHGJG6L3xiYeNU119A3B/Q
kHCv+/jn3TUrDW9NPuTpEkcxRfyFvlmgqw+lYclu94ihuTo0MJcH9YJvkZoyY0Q3
v9d2+I6Op4J8ypuSaPp3Wl2bUGpdA6UVO/fGWiFCXrwG+iWx+5mJ9wVFJzTit1f1
keGXKbrNcswkawecK/TSSuYHNKCcJj7Fv0pNzzH4r4iZBfjooDCRS45z0H5aYkDs
+MRNKj+y1UTvrwSOawUqZoohn1ZI2Kbdr38eMemWhb74LoYSFuVHax4nD4o6fPUq
Shau3TX/kl7A5bhyOFVXDNpoDrVolueZFvRR1rjdjT1tIG91Ua7iUEvVzwgwFBRy
1R4vRCIg98vmTw9ZrKcVfv35UtoaVK7xtLV44qQlB2hOEJaBeAH9CW8dWoFmzz+Y
H7VNO1bxWMo07VM97HGCgHqEDE0W50nGYKvHbgWxmDBO3ymouvfNZEdQ5kzvqzn4
EdRGwucOzKye5Qy0iBpD5MFPTfFWPJ4pA3aNuvK3TYXjWIO/bM7R6j8DE5txMC2p
rUzQ+4CKA2tjJo458PKjPbKOmocYPnp+TPC/Gdv93yG5JPrNH9fXdUjA0vaVDdic
wTmZjx8Jey4SIS+ty9TthwD7kOhAIW+rrGannzxGVek8leyM3HWJHKGdHptoW1PH
pZY+ck5LtG6FwtOiMZHE/hkt68rbwEPOeeXtFEotV58KiomEuOYMFJNcsnCvaHle
9BNF91oCEwLB8l6CkGELDG8+/bZM2pCZ7nR2CCivWVV8gY23oS8RJEk1/as/5q93
W9W2fSRwoAzFEdJyAZG8j2ac6NVzHPnHqGQIqC/FduqJe9M+vF960TznO6J7QKHI
7izwrz6BExQO3Xin2fqlXtfDcM8u+yonaz6JpUF4dmWwQ3yTss6j7We/o4pI8mLy
k5VSHGzZGsnY0s8L5vAj9Glyr47G/atyw68o8JZ/Ig327+9Iy9l7nyAgFqfz7M4E
ha8roR8hW7jzzWOOlTPYZ1T34BMoO5SG0zKZAHI1o3DJiyO/bjHezCFHZ7y3dYXr
MqCOcBhHyCMZk8fKZ3r78veF2gtEWpf/5wfGF1hXnHp0DBzZLXw/1YH8BOaMb5F+
XSSjsPkrMjALjG0IcHavXyCKlaqioAtNiM/edQR7Owh3rlHIVz87k1a4cpq2RA/N
Pn4ofuH/1l2dsRBfHFEBRx9k6eKcPmLkzzwYe8mMeKdmIAsd5sdhfdHIx9U1Oqn+
VQhG4EEBY4HERh8YBP4o4H7MkQjq9d0xeArwoItIm0tgUVNRC6W5501mAJ0oYUUQ
QJfglCrTXiG8YPEtAI+cvMzgfD1iAG4TBqFMHnfLqMIm1NYWBB/aAv5Ym3Mo7Vnc
45KODUJSDmwyTd15Q/dFQsT/zMElP1ZMMrOdvJgbxV3Y4erkh06sOqn9LQm56eAG
0ch4baNL9M+A8cX0LrHldeg7Ve2tt7+SCxUUl903UnUwKPyIRWxDlcsA2nDuP2cO
lONu5vfKvtcD87VOY+HU9Xyjlc1LhXAQ/94are5AwdsPS38rzqaseq4OaGXoyhgO
98vJUOzp0IOkfF5u1gAkeod34r9IjE2EUEWilsQzq9JQiIA8t1UiFeZZFTQmhsg+
b8UGRzPFamSQtugXvqZ5Pg1N/C4qYhD/swvIilpn/frAF/l0fXADlLBTR8S0UrTu
PxMD+mUcIzDP+1bw14uMbjrWaCe2o4E645xlPj0uSGIbflCUGAWOZpcCiAnrK/Sx
EdJIsNqmTA/H0w8jHcb0GM9OwAK+Rj8qEhFQ36soO6Yy76TZXEOgGmvkA7JoYbaW
Ij3caD//j/n+LMBvKe9X7QNfi/tZr/mqEeCUgWUpJbhC1J7VsSuCn4fr7axrajpr
0iCars21hhdJ9QVI0OVA6hqPf+RtXPboqN5EWHAEsLKoW0fEFqf/gnkwZ5jrUSfQ
KVSHSsC4Jr+R2Kh00iQjAjy8HFXeGxRd6HkiPBOJfg5AMkLHCJT6mPbNUSKuJ4ld
p9prCZT4AcZ4s50HbV4feN8HdEOFfHaoe1dgF7y7TxDovuECvazjXElel/7Mqf6h
sDM14Ow2ONO+/lYi4vjiZ2hWhOSG2QI8rCp6JF2d9GDpS0kGyg4TmHKBNYYpz5Dj
lgsDmgQ3xlK2yvq1ckRGm42WN8pilbGPmGeaq31IZsBGsf5aniK0zWRcxVMhp5/x
m7SA4PjkLMQ5c/yZhnFkeI6+YcAfyNMNkj+kDRxe0gD9C1O9paiG0SxlHOd3dIAL
ryFM4mWjFlGvohitSr+WsTbDGyCL1gCcDu+BTD6qJ2ndMYiClHV//iWUAACNkocS
Te8g0Te/E3Cej4VgzjK7viwCDVh+FP2uGJDkx0dlEpsJSuJvuMlO5IyZR5twyCIF
WbYhs6SeBxZS+B3r+m8AWZGCUdHx/imb60XyjZd0hdPrZbtUPvHqI9Sbs3iYmHry
3/z7Gaou5gfcAhKmeDDA4SS/re0uKZxBHy5qakSUC8YkwX2yBTxzC/+qbSCCjcry
Wney9lK0NV6ysKUrHbJhYwSYkRfd8uU65HEqSgeTdFyz3A+EWscDLu+qzLvDtZIU
MoLkMAt4Mj427hwGyKprn6tkmsBijQZIyNYAecEuYBkWDAL/qy/VXhWmo6BsUjzo
3AweK8Ef4HCPBwkL6Ii3Glc85ck/gSRC54p+gaFb0Qncq8+s8iCS5eWp6gvDp8eo
k8r/pFWCAizG9LRx+krUXl3bgmt1DgEqlTbpYzo8bMaJkiN0x39mbts0R91zN4FB
9VxLM5k48PfXEpwSXCwgN2l9AOTfGm1cm9/DwZu8pNgLqSbjXCCIdktIsGvAe7Ke
a9pA/tYdX3Ou+pI6SCThWVa4aVMvEq1EwhyqnEOwH4DcJWEiG0hHCDZKjbClr/fL
Uh7Xu52r9+BB30IfjAo+4sxz2UswETbv3mmFTpcptvOrQXQ2synDBHTXXHr1Ii74
JOxTXfw4vdNFiRpkxlWYcY5rTqtmc2TZEm6Rfd3AUguAu4KJkvaYCWXwWNclMcf3
39Ydbg8dVLnvQJLu4kaV6H3sTTAHNBFq1HhWFOiGvo6E8Cgzac1rL9/4JrICbnZW
1xk0VMtrUnN5TPzXlj7GWra/z3747SsTdGvr9UmFuEb8138eW1kPZtmgtxQdSpQc
HVyFctCwFS/RgnAmytZKe6P4iNXe0xXZYh2JbX4zRzV4HSQbyJXFVgdn9nJRPILS
g26nDiHTOOp7jVnjDp/ig22SvHutFQpOEfNNAJNHufNwFWk5S7E9Hc10H/rI8xth
o8mH0DWhfrk1R8BNffYEWLCOWrvLiYdqYkr8JPPaJJgEh9yxLn8iuZ5XL+laqV2O
lCrnFZvczA03RJwC669kLrRhf8YHI2qaGBBOkrU6sDD9H/E29+iahHMN5Gni5742
6V/RWthhDT7XHPABS17sUbry4rb66UcOkrqYmiy0vqAT3ViZj14C4FqLd0ezdGO4
uHCc0WSVRf9YN4pFAjDEWKGp8sVP7emRgx7tmtZ72blKcE6zrobNvf8Wuyo7t3TE
OsMceDjYv7xiQdkEyAYSIFsAXpPIcTFQioFAfkxPD3HNi1WZqCj2fTADGqVZOqD1
4n42KMZzpd/bniAUPKtW4sEjTzbT/SGX+YJDmGxNJj2UAdJ2S87WSgk/PKH7ogmI
MRkfvmynp+dbgnc0i0VC7WVZcbRgD77ZFrXNXGe8FsgQK0qbsi3OytNxlAFPD54C
FKsegT3Y+zaLSJ0TnLPbX/FWEgTVhWQ2btTd6F20j4gOJJN2H23nIFaXevkQnLlu
i6NGhbFlMEZ3dAQR8wyYkSkWVtYga6Ja2qy3PBVbLVPyCbqQiMkNd2KkkZImSafH
O1Ohi6rV0XlQSVl9W+/RgIDDccLGggJmUpfl/1greOeXBSqhtdA3QNEEe4adI4Eq
+yWWYEEif9kvFCxPNLGiQe+bvBNynHO0ZrxDmBfJQ6UAoSyLjDsYlpeqSWERbosG
xfK9fhiP9fUfyMCoXnJY2SwS0xpc5dioJNSimY3eBrCW2xShhv/4OIgTxSgc5Xto
A2pNp5RswB81MmYnFO3OadjmdxPSt6vz5+pKkjLCL0xvfEtCHJ+dWjNm0KCGNEr3
miIZ/oRrgpKB0yJBdwwLGuV2cLZmen8QndVxVbYhl12J1w0Mi+sH+DdaMVi+DM9S
O6veaV8PllIQAxR0o4qQiADHgKA0h4xmvnKG9ltodVnakAw/48QkF4CPg7ndzL9M
u2a3zPNVNmDr10iYMmhF+pSaarqOFV7jOc8Hwlb32U3JLcqK5gUvhboJ5E5ZeG3d
xH9y2h0UeW6rYynzBjVWXjo1uygVb1g6X/YK06+wutuQkhfa0WNXEn/o4rRuObuK
Uxy3wUO43mAc+yeU+eAfbLLNHe0OW5A3xoB/dYpbUe1HdxnFBBBFcX5ltYkc+PK+
+MjApLUH928idCBpZYvn3XUpEmoBvXsiE/Z4JzaDckhrd5yYjmjljf7IqG4wSbDa
DdF4OqD5nBOwVvzRbP097oTJnazF12FVyeLt7yRu74NvVX7Xy/4cOZ7yT7IZyxQG
MJjC6+lzyg50Kix2ANwqeVWutLIa/vPrN6z0scJ/+sZ+4V0GSzxPlug7z9rXbOye
Gkw0aoWSRBmFod+ul5/WAVclcByyVYuTsYwPVKWKpHysyE/CTz+fl8sCL6FjzyYo
bHlYsXGhpMbxr4S3Iy88f4sBZE6t8UF9cscxVWDr0ksHDwEiGwLfbJNtsl3oSCFa
C5jEjxhwxdw20T92pla34p0O/iOHOhsJwPhHta4QFCBAx1jkYSMnBzjQa4kvEPts
g47+KfnDYUoA57zHRYnpjXBSd2x5nqoLj21POUIn2nkpCd0Dv2LUo4tq8Z8G5JqF
8GZyX1u7Y9dIxoj35QZckRWyyRunMxkJEBrWvBqbp0OmlxL+dxfOaA7Lvi9d48NV
FAVANVlSqpqt8SR0TQxqr8TOVIJaAlKbV9/PqEUZRe2Z7BQMcRWByX3bU0XehK4j
49unUSaf574iAv8feyXRKLeXfWwp/qz6Glruw1bdUaKHmUFgv0VxlZe3hiwZp3aY
vNCKHTIKeqvZnitv21jqaOvm5FP/2lWy0ZU5rU3U4fiVdDTs5uCzScuSrCdcC/wR
m0D8iOEqLR2JH1lzuaoTI3ClAtY2Uu2RwNDxpkm5Ok3lpFLQ0XXDm8VNkqkqtp5K
115mSV5cJsP27DXALV3NhMmoVCbMdQvNRsD8pKH/J+JA+xNsJWdkD+w8rscsvjeG
5xaS5mpHV3Eojhw1s/zffz+6RImKEF8LcmtykVeIOKTZ0wlSM1B/7vooxlZCA0sM
JaUzcTZSBAn07/qA+e8KTtHS1+TRGZCiSvnojwSuI2oKpG365MOCcxDHvwwKiMaX
LwiZ0DweWOuYbsf29xcs0DuQRbB5QTidK4lqBLk+mWWBX/Ur0dfcBEDD/jbtW38E
yRAos45MyyV9/27ArHyGMryiTOwuhVNc8ppr5/DO4QK8z7jyNoUImybbICQIdXA0
RUuQeLxmLYYGnugZOi9NeA5gpgA3rsUbzTT+rZysF2I1U7+wHMqkUYovjxnZ7LsY
6SXZ7Gvo7VNmE+gZxqPJsnSKZArIa/egf0sKGWhUexjm0N3bKOzQMHXI88eVQgD4
zemcM8cx8NtOcwVe6yIw5w7mhQPedYufHRgf85GH0fM36UVjBFTcDlttbvEahh1G
a1E3CDs24jEtMLaIi+xa+g31lbSBv+G/gdGzZdQo8HGS4+pgA331sq/zf08XxRxW
o8UJ2WF9glUrgydqzyvM2eoTFTdwwsuv6lUGUdeQLFkBuFO0xBlaZKtIH6pPMxej
ZPcV9e/Wt+GHPy22o6jxn9b6llO1K3M8JCsEtCVxUkhc4td5piNjs/ekJmN34jl4
A71nInwFm973iIwbYEr4fqOrWv8YDLV8qse68zBbWPHADC+SV9xSrlCmwo40/v9V
Z3I+Z/0d7U30bUgob0XWchgFDh15NEFIUeHHL+RtL9AA9FwO5trvH2sdXtBu427D
60yCvjXe1J+SzroVTW08UCfcTDR43Pib2Pxkrxj9MAE5Hx5eHGNtPLBY28c9Qdgo
MmfWNojmyk5QaDRiok+XGR90hJsE5yOSY+x454MlF8MzgXv6p1bGj5IEbe4p0v9F
P4mRdqmNasUHia8E2XAPPJy6jCDwLqvyyrzHezp1LRKeAxeeVCCokXpEsPTMRtQn
H2jKo40CW33hbCrEoSss3RI+liFo9+himexT4BRpRarpxXTnirlFi2nNPL11I+Gj
ILOpoCPk5Set2KBesEwuAbz6M3Juu42wGQzIiQP7KxBNL82AHyZCjHRT2DfRsYOX
yJMmQiRr+m43AWDaJaR19M8YpSjfrYbEpeN2DcleLBMYRz+IRpY+d2ANOluYx7hG
yfSlM5tzHNh/VEbuGfEQXP5rOfA1atcFZ8eBKpAK+zIJdJQyExNzIfF0RZPex0VP
jqJLyzsCg3Db+xP4s2HkwkHQFN0ojZ3LzYPLQXS5F+VZB87St/rXoYzhDSAaaqnf
P9tmayL72ThxnAePI12MYgGc02KqPAEIYgVy5FGJ9ovGv5LbNLJ54SbM6zXN3Ckc
IubRKsjmeVkHiYmt4gB2WMqoFX3+g9hmM4kOdBxXMerROHJzyQmb5D6tLbIaElQN
LrYS9+YPNQAEIzo+DwrKz12U7N3KtaPNqLey0IIE/no8rP97pgg2iSRhzoL1jaGf
0l3/vtLpK019Zw2RoHyjV8SCc7Bb7iU+m+ve8rQxcqrRYhkwNNniE6rUw3MxGXKC
PxcdwEbyEXhVNh+g+Y0U8VI8xfZqSuvNKW1C44P6i59p0eErCRZ60pyxtEIM4N5j
vwhNzQYJ+CZMBQq+5IgtyJrP3PWskQFdaFDH+EAEWmeitRxzKYyIKhfODE9YcYEI
IiFuw/azDCfh78IW8lxLzV7nufO4DYe/jnQ5KI561sbNCRPE0HrxTDKial94Enva
ayGlRaHWwzBWbPwjLfYZB7IeWMZ5atJRyldJ9Brazd1XGEkRa5e1LkJf/lagYi4X
pHSICKq9lidBt2AQy+KHhRAXYnuH/cNwa+CpOPOp+4enB9BkjWZ7ZH6kMJsLRUfj
rYuwsyVYm+Kb84vusB/5Ne1WpSnLnYprgpDXSY5wG79Bp6cRMpleG0c8+lvJzSnK
rOh0iloo3G5ttNR0CsA/duPPol8AL3I5r5mTPPvzWsFPQ3iGqONp4ztDXfM3Rezs
GSvyEeSzQo43KS2Q8B7XVg2ta1m58vFBv2J0VXSbyGvCHk5oBQxBeC93Vz2UXvDN
d1Ju3Oo79dKnPmVlqDyuZooIpdGG/TIayLLWI+zmus1my0jOXDKw5t8kCNCCnkmK
KfOnu+dCRMFOKDO5VKx0s78l8yEqJo3Z6ukASGWDEHyyi33Q377JMez5TPfwIRd/
FplQUIx7bvo2dnoh9ETfIzf4nk+3WiB60jJJpWQIQoErDkX729MZhxp38te2I1gs
rY2lRO8jj/46IW4t3ynPtV0Iw2jKIZ5JDqZpJklYZmEgRlqo/YvXTm5Cp9AIfbCk
7VaSNoLqufY5Mu3DUP4DUatsWHczFooUpUK75tkJvD4es0m8X/lEUxHaPD9/fIH9
9K5vcKOMhgkjk2v9/wQVO4wwXzVedlWtIl++DqgapVYintrugFD2Ot35AkjhhrF4
kRYX1Ju0QNgpL33qmvWBl8feVSSRUQOE/DxiA6Om+7QXOIQHLKydQgJxb6KeH0eo
xtrSVBKyHNQUNiXU3qN2aRdn/gEqnTZGcMFjUMD/JH9ElPBSKh0ONVZPAUDw+Eas
QbYob2HzhXC70runKvqUV+kymnn59CeSN5JPSUzk2bSJYFL0cZEPx+C8PAC8o87Z
LiYBfG/0swhBahjl6bYNkA4iWm21i0IWttuj+Yb0vbI7T3mWijTeQOm72TcxFm3G
BWadrcLdsmqetXKcsyntA0euOV5g4AyWV+jnIgz0iafNE4DQXf0OJgN4uJLNroTo
n1lApx5rBKkv3NdSVTxw+UJUTwRFS/dkhK7NCsi+USqzcPTAdGXOSgR3duKnZI98
ewx1x4rnCgp1iqPB/e4w5ECqsbt/nItVwKIzjbAFu4aqiYSjF6qlDjeXMa88gNDq
tyHGw09OundARBA44LaOUxdS1sblmw19YNHXmLplDQVFYRFa+f3FrHYye9oDNJS2
c3cmpMwi7GuT4PZ2pf65oU/y/+fAVC1mo5na4JPZ0U0rNSnUFAj3c/QsjrNreE5z
CCM0vyS4Sw+dUiB14XTB4IsbbjxJxUZkH5H2y561zIi38RVDKQD+yR5tC0HszU5p
hUFgrz4R9MbToddhH7IbbrsnV2zkb128LKRxg7H2sheQQgwSL4/KVkicObUNPhB1
2Qw3Yw/yC2iku7WkW5DvCKpIDJPkIjlKmTzKejZvC2gwwyBqb6ppGvYE26Yj8zYu
8oz57Ib26v2kKDvo+DDhgJoupuC4VEi501Brh6ipmipxHi1FwOb3b8BZDUG6+Omk
X35Fd5Khgsm8CuAfworeO2bY3lDx3AOl/8L/Ebn6W9uje6TjtRX0aKMmecgwgIE/
0WJn7iHbtMOzqB89F3REz21jv15C8/i1CgXKQOMw50VhkSy1Yi/IL2KJnv9nmz5c
WqgZI178jsyDp6E1EzPbTIhNchnYyQnU/QbjcD293/HKkhrtyg6FIEOf3muKdynA
UhMPWF7PZoc72GSLkvmK+XDXbfEKYGQlfjn8l/uDBKTasSTfiWCnh2RcSfgW7am1
c4JtvN6DAWYB2lqCmOefyTomXAxrBOVZzB9849SmdW3AbMlpeMCuLKaU9pIlbPuj
0Ay4PYANpQJ/rUwMZJ2PFZi0cnXi1bPuUyNSlwk64IItS42TXlqNhJxM5DiEZOet
BtDb9uwWSKFpMQPBwMF+nAWF4fgm9StbhS0Ztr84pT2ZwxyBxktKE6AbvoZ34I23
/vwSWb3ov9wqifLorbwG8Ptgwn2nWmuHi2au07S481rWJR9YTZl0XD1qqzj+9cpD
EnKG1QFZpEL9NuofqxYdU3NJonkWA/Ft6Je2Im5or2qYVkBSJjD6MxcOlO11lin2
Cz9aMW0Npy5BkQD0zmwO75DDIrsxvJbhtl1iz2JuU7ev8iV83bzv5yxR4y5clHz+
vsXRxDuqk9pIwQ+yjI6AG8DLuIIPR2CGk9BgzHdvZAlLefmF5Ko6gLXTWtiMCaT7
cSDLNZLH0y1/G+cMCy4s+nNysbpO1BeFyW2FViwSxVa5K0p0//JWNAqyL8Df5p4U
U0qSYbqS8fh5CJ9QO2RWkuYjKs2r6aYVNYLf+Bnr33+2eD8fqUJFbj4T6hV9+l8p
vS3/k/QQZ+pHKLrizKu9goojq3n6TGYiJASimulolv16slLIsDzMgHU1Hrld17I7
Hr/pPrebIhPSnrdPJnKVmAMtiz7R60lrtpsgxKXjO55+tOYpt321dwjeufdglQTF
JXaZvsI2ZvTyHyU/SLsMctlMqsl17pH5kufd68rVumcnhFVCF6sO2zkkdu8qLgbA
6zixu2QeiksadWGflOUeta1JRD3LBbwu7ItxtWuZ/2VBdsJ51VeV6f+zZaakHUhA
pO4jLdUzPUc5olZ9unwtOiDfT9cL7m2C3ViT3chLGAbmwT09BvW9eojH8YNBEENF
M2h95VyUtxDl8Z9b39LMslyF7oNqslMOkJSe+BJ9Hej1R13O+Ty/5ZmnqSLCZ7Vt
/iSDmt4CLwrVSvodssWQOWNuq+YW/yWt0fTRGTkkIeTYNacaCaGU4kdyYElxYbHQ
WO6HYWhR1J1MAfCJ/qpWI6FoUmPL3sp+qnbdGTupt7KWyaTX3kjrZVgKXz7I5q2g
6oeZJEvp4dBJNthjJbeYGNTf98HqD/ZIxDLDGCrUgkQ6HrB6KfzQIaG/GsXcVioz
QkTF7aQOehqXEF5rGdmstZdWM+jPm2khTU/ayaFZWio+elJ23tn5CgsO56RaZWmg
nMCFEZ2QmQNGGXRmjMq1Sk1rd2akLFBvXpQjbU53WyuZ3YHRq6Pvff9TIbsIM9qZ
LLBdiIZAeSLkJ09QxK/car8MS5U9cW9U0VjTVKrIwVF181IbUdXxkorYcPjjGECU
bhGDallnmoO1xHVaL4T53nksW7TVnyZuseUI4zlb0mznEVj8DTS9NEE13c/cp2GI
rC5cnlVgfxUlat1R6milribSnDsoW1lwD6ei6rdXA3RbHAaQD4rqyPUDLvS+fzML
itq/tBXEFuzhyFfOgEiYAtM4V+esaBzFzKuJ5WLVk6UfX7OU7lTr6s1iL2C0wAF/
8ll2/qAfsdHcl4WFXx32CGzBdxCNkNHTcwYjBtOzOcOrf5/i3nCyvLV6P2uf4GZ2
txbGDIOLVOAUn8WvqDaGkJu8Uffyv+9yMQ0GjM5XzQ8Epwge7pNjxiU/aNTulkKh
SD7mAzOcRPAMmcq2WnYRGqR+EFX/sKoEivcaKv3ADCN9URK3C31m3A2G4tBgg42r
hew6fBcPFiWmA2QJbBhkAOetn4hSKIvroc/jwV0notjdxq6d+XPYwUP3ilP9UXrF
ng3iKrQXWUxLKra9lEX+E5SVVIoQ5U8lJ3JemApHVJqiVGeG34fcAzJJ3UJe0Kw1
mRGFQszz/dpdtbiSi+ctP9VwSQ9otffi3sxWFCasgV4pcaVGfP03nUHu0yCWAxY4
tv890pve9nHyBLlSru/UTeAfdcFCMqJMcDmNVbaKX3/excAMzg3qJIQxNtc1fgWj
cA5FKug73Ywm2jlaF3EMDYI3NfJnlYXTzWIu8CKdPSh7bQFNNop2UkOcFB488Gmy
zdCFMK60YeZnIv4pdtXzWOvEOuwfVdTv7UhOcKEP+yFZzUDfm5jiZfJIu4HPche0
NottRi+Po+vEyO++ivYWXonqLFCsvc4jNRiuzh04Sw7ipPjnva6qUe+sl4Hjgrs6
sLO7RQWhjtvPPxvvrpCkFWPkRb9y8cWgpwyxmmM/1OxhaF3eZcndPHiApTSyFKo6
NZSmKw/gEfa58fG4M0R7533Kd8JDAhuiOYRPeWDVLpRBxCCTq043YFwa8c0LtPQL
921nXnR5TEdCZGDb69j7cuIVHRiDq/bJJIZd+2s8BfAboefnnp1RXqp8Sog3x7XQ
11Lx5uV2EV44T64OPdQj3lDskwhgtvcpHvwbkhcHtnvtZMKNcO6Ui8xRokp7jjWt
OQ33AgyTsKF3ieF5wXZHssYI/sz7ynDjubWgTEOk8X2dtrnqygZOA+nC2YG952wq
zX0V5EkUQWz9xE63MohMIzFUHrr0vFwOAA7rrCg67svWWc1paVTK0ourS63G7uQQ
ed2Dtr0ihdVPZ6KaS7soiDK8L/83t1r0QmknYwb5tOY0bfbP7q6jr9exaNiAr3IC
u5fnGD9/yTqwOyH/HEa/1Qb38mKD17eWBkoOBQoUDgWMmE+8d/mYoHgbUhd4mq7q
OG0tUXTBp79C7pGmblf49VJm2kie/KK3JJIDSnNoF25TSzasTby/N9QHE02PDVap
E3jb/EhEFwj6Qobnz7UFyNQYkNYum81mTzmzpbX2Lo4BPPaIPqbcxELRJR0R1RXe
KBRxcekp+V2KQT3A7O7KtPNLM0NWd3ElHN1JzIjIgPWu8qfsmwNd372dmctWGyAI
NydLtYJvuS8HLQpCpI9ZB8EAkFYRKZLr+TRPLouvsKCBwU4guR+XsLAicw1LstNs
KrulFBGzeB/D7jkz7vcFUrOhQAhOJ5kVzHPOe6uTj4x30fdMnycsIAtyy17TIqJ+
8IEiUdrNMcbh84VvnDa92PLeH56MF3hFaZY9eDWQV2RH4mpWD1YHjTdzDN1d0OmQ
lrXVQ8vWCOGfeKuWUgZsOrb2o6qn5Cyxe0MOlpC75iaQB/2ihJH7Er2A2Y183+NI
VgpLhviB6QkuPAukZZ77BAUmbck6RGAoLGAqNf3V7ojXlaFH7YOhwxbuKcjo7Tim
QiluEOSi+7/NsVK4iYD6oWqZjyxby5OPs0+uDZS5NHtTaUDVXt/tWrfwpi0mSzX1
XeYRJ78qcXq9r5Y/R1W+afz/yufDi49pN2129NVWyIqQOIYiATH+nkKWv8Igpk6W
puLkYL6rFxsnfd+Ecb0C24U/JJ+qJp9YIaIcjWzN0RoMFHj5mybpqNqscNTVeHqL
3733U/zmqyarYy3KuH0PCAuWwqpOUHePW6fZIqCYGIIzSm21oSZLUy9BDxPbn7QI
fb9aMzLlKk0c9zO5eoCxP6pCI7i1SbbfrVROloGw5rnCU0ZY8nFL4F45B04jnypQ
1tutjvbEQlLPU45B6rlABxoZ79euIkfFzs59wUEXLSb+KTAc+NSQTfs97mw4Phdf
GQB5jtx7K7cUsc3A9en1C498UAJXgpQhhT++MZj8hslTr1Ydu6FkQpJ6BLY9WSH6
UFaKBQC917vz4Pr5YG0RKLefeIEmlVRPwt68oe9x+ovQnmIEvSabs/K+a+zr4KIn
rDB2iDvanwZ4/rB+aRHRKjGqLGMsQSzwBv9qcKSUQTyYSK7EwfBYI8+MY0lZccnC
FA1UxJkTj2nLMaJi2/N/lUvfsZLaOvw/zLSE6sogAv/AO6KK+evktC6BtLJDYNbv
iuwG5nM4gVp1+yp6Tx1Yw6x8Mkgl1HY32cGU7iubMOLCNcuzWJCa3+himDEMRUQt
TeykASouyww6dqmj6oXtr4XPDrNDWzfU5iijK1W5bcYHzF9us4LFDZrEtG2brStm
I4NnMqSjXAT69HjYJw2OU9gQEagpjug8SmnNAv/c9NlcAUst194fEnawdKtBDlP4
dnHcIjvZZZPfNvlefASCBZoyqCLqtrMYllfOkZoJi3B62Dzfjf9uwkccywExJk+g
nsC0H6qVOsy3jVW/JA5B87hwXP2oC1atVv3u4R9vfalYJHF6LQVDzeKONXmdD60w
pHsPUsdyCkPGUmSyzmqt7SF0QO91sxd2W0akWms+8KL7eCOfWizKhCWqfnCdHuWY
572PQhQ9kWBDYTYKjnH8xWg0j0oUe4awy7DUjox3/UQp4hDtStLcLHCLLMF9kCSG
WmuFhFVwRbXHb8PXWPEsoLJIQbXtlUPMSXewONFcn8jxunwYhzKhe5r3HMA7HJsz
4zzIM11kedOVArfLkBqW3GMQvTiRLD5MScxSt6DJeDAktyGq21ju2Fud37Oe9JQc
27EhoZVOZQHiWX0sUPrPYxpz67qG3ug0cFGITEA8Xbkqw2dMrpLB9CtCmgfu2fdB
yWfdoSj2axiu4ULu1tp5IUSk6VT32E4R2vidLaDQmhS35xwHV49mJxPAQFNI6uck
zYgpodablg853CgzikQMopcjkzgbdGYWDJykyZpOp+W8gZBjA60O/hrydmXo3QHE
tTyAm/F7M6NawfIiIk8JRoL8B5O6I+1oCfaO0LIrQFwDcltnREb0QRQuh79vkJp0
XFzzJcesAlHoX+mMohoeUjkvwXCoRAj6/RCwrOB2wILnzfMKsxk2PntZ4BmC2sF0
pPsik4Vpcm9Vvow3/85a3M5J0Z/DpRU93K9Vg/9L6JJzAACLHWcH8pkiosHxcwFc
GRlTa09+0G3ecHUaviD4tt8EVchm+G4E5xtno1s0qrNiN20zSvva0ZacI+Rl+aqc
sIea0YFWdbkUrrrQP5d3/MHzHMA91Qd/YmbBvwG1HAnZbhU68fkTyFLxS45GBmTd
f6ZJrKEfTr321t0NbGdrrvkxDHWO3FzYZn0jpNOfnUSFiXWF7T4bYofYvWSldiWf
xYZJdVQrnHdN+1W7YpbCFhb4lJAiCJzOKivlOhQpJKH/cxKmsMA1hmKrcw+JqfyE
awkiangbggzFMZ18nDj8cE9KN4EKQTISBmLvHUD0jv2672j3OOiNK8wB3JHyceZW
unc6E1GOVRUX63RxdJiD9NSB5DolUdPG6V0xVC7BgYHhririQYDwzn5NzsE0aD/L
Ej7F3Ne1ArqIPxd5FNExW16r9MPOA+bJgY7RphfhS2kOl/RTBt7T55n/pAoTubGY
MFJCzm9peAJJ9jBk5Mtx7odONDE3jpAK2YxhLr73U/hJFRhbNlgdeOFKmt1qDHmq
/Z5qNmmYhaHKGreRi9vhPeOv5u18U1aPxeUntzMnQj0pSlY4+ZL8DmUNdUIcfQEc
Xa/zf+KihxrfxTtARBSupBJa1fmYJPIvOPctN2xf1Rm553QaG8sgnPZgf7HdfqTH
BODcaNfGgDdjViMu12iE6DGsIkIHRdFKkJkqvVAOMJRNcHfvZslxaBgVsHlgISOb
f4lk+o8b7NdA3RtF8zR+wq+O7NoqcJcENsn0ZeiHPUYWQkgYrFgPQ/8UbgFsFgI8
AJH1y5so4jZjgr+SIjIZ3WMGmGHeAiRmWftZ2XFrG0/c4gJzGDbv+7PjmjsBk1li
OPAUmjN160mMyDFDJRJgwonoaL8XUypQmoFpUKiDx/K1t5DlmSojtVCaoaiMdly9
5K4aiZKcXA9tq/3V9Ik8WSwKN59wGCmKuyy+zFRdi3UymZcsWzN1SGmKAgozAZpo
yKenc/OKTIKsYJayPn3mVIw8RhaaeL31wsQbrZ9OcX8fgOrJ4vIZQXvoB7xBd65T
U12ln7/c20mGxEIQh34AUutp3QnWjxMN3E44jlER4QwWl5KZIk7U39i56HDX4B+B
Ga4t99NnG4TvZLYZTjIN6G+d3IEt58qrqV/Q1S6l9ulTmHYYJdH7vo9AMiELws+4
qNqgA9twjYH+kEVnP5hg3f1uq15mknzRyu4HUcFk/r3G9CWX/jTox9lQpnjmN4p0
9+d1S3pQ8knhRLEYKSQAl2xZugTwRyFnL2rErTkfdmPAB/CnE/JXfpK0dbvWXjXL
nNeCzZ9GFl7WRcSURT/DtWbKpoPVIFFmCxZ11uyPXzMHLTefRel+9VytI9X6IOdI
XMKQ+2Nat23tF9sLKBM8WzmBbcgGmaFRWU0b9E+fAwNwzpjYlPolNUpu9IINEgZU
1A4RTi+/wjE27RAm3lV0cFvU0EwsKMWkFW1VtFi50vrOi6FT7jr4VteCfniaN5+v
ZdFQTbmJ71uH/NUbcmA8gKTAHkFxcyOZYVeai8gLj5VS1OEW4+wbMPQrOEt2uKkd
eThRBrQ9bzTQdA3Lt0K9eg5EXUe3eXgIwUAj38Q6nGcdqSDNSKDeOJxrAwEd2XTl
66Th/nMPoDWrn1u61S8+8HY/xx0nZ8eSsDIDMuVp4btZnxTHDdVDuDh8M06Pw/ut
3h581Su1MkWElxUhltRNF0nE8gfz8KdlUv98kfRY3J6LYz1wXc0s68ig4ZxGqzrD
7QuHAcYsosVgHNCsNSN4HkvUgvuLoUvviGZkWColJNHHS7909MzcB93u3yHJW+k9
7YxXt03ttHok6aLyM7+L48oVzEE4AwrYTYi33S+WAN8xG9x3d/Cdzi8mfp4Lmyqo
tclzcK8C3VXAot8lG3IAmLM3saccc46Rkt2kVlIZbxPht2mg/eXuYzI1B2uj6MnM
8Li3SmPTkx8Qn5rmqPnx6jrarCpOEECZXgBI6yhYMDt7gK2jLfIyzKdIA7Wzvwi+
b8MtlxKymqjksSPjVO+2jNOmjtgm8OyrQ1QB3hz5AvMjiDU9Aw5YliuqXePadQBe
nANlVoMa/cnB1Z4SesQRISbynNAumB3ngkpiEdgx7/D8Tl+PEBvnlZH55/kmc8oH
vXTSA9m3/tvRJgZqCdhyVKLGK0uqnhm4ZCMbCYrDrQI5gXL9j2xIM4AX+6JzKxDo
vk5n4dUX97QCiImvTynFqar7wk/cevmy4BSfCs4VkMPbnikGSRZ/8xlNwqhvlkBm
3aT8Wjnm/edYs6X9Q2UWkapsAK3NNET/PsYEiljEiOggi0VjDKhKYap3lfEtco+V
ZmcVEyGRKIktMh/JrgMJ5a7Z8Z6Ys4vkM59MX0RKX3ZJUnxNe51TK5df2QUDAQEi
m7dWN9LEDm+/nkPZZMIDGS4f6eIW6o6OIjxGS5+e1L6spQYvKqsu0acmXv97EncM
aR0whsjHa9SaLnEGinG3lNHSGVRjlBc/NPSGMCdPOZewFbCPqAH/hC0Hno9l1jNE
+JTth/ejbJo0KOlJHty7Ucj2h2rGy5kqWSCocnIB9le1RuvrsxEIrmh53+dHjOgq
GchISoYOGj1C8PGh2MuNxBalny/rSEB4E3V7uzxx8ocnaLzBMKFxLvXiUimCQQxj
7sQzydqVLHb/AX+zXhrixp9HRyiaLYF4g37ON7dXnjdiKRUx/pqF8PA25j3wBzDy
tOs1n7Qt956fojqxbL+mKcSma8E+26bjQXQXBY4ubo2zBwNtCDjoiuQlVG94QV3r
yKjH0T3M033+EDkNKPyQUnLmsTVTe1P9fWxIhlDcCj/10F6R5nqXnOpaeYyv20rV
gbWcHMWfajSMyZV8dopzJMDHi3f+6gRcgjTafnxRrC3PUK0hXUGUF0RFs/sErrOb
1Vdt58em5w7bhtkefl5A0oCq81E87xApxeSd47xwZGY7FtwdxQaAm7n9CBmtOoej
o1/7RH1GACMep/J15euU6clHoPVxj47ebD2Kq5a5rHMp+pvurKEDbUulQbhokNQx
ybCJZAc8HY5yP2SIG/iyq+9AKpkObsrstsKP8hMlcdvoDoUa90VOKWnPUDG0QnlK
b9LLowao9UjkQAhTiFNQqKeHNxmEDOllVdAfmZTto9ZzXSPwngJinqG2v8YrzoJo
Iy6lS8WkTFDMSByUlh5R6rpFj1/ICNvZIDwcSA2sp20nFIafwKF0G2ndztBtd/4Z
NxXl0weDisSZjrBc34L2XjF3UUv4nEVfWUPlSm9zQJMcoGx0QSABHpL05+w/4CXf
N1KKY3rbikBels5u7yKG72bxlPmCefvG49l5vY+h9SRFgl0QloucSbHk7CPsmSdX
hFAW+tuMpo1a1kdIYA+Ey5m9wM7mYjXlLqgqGov8NdQiUuduMJBft/rNve3m3n64
7cr+hC0VfyfOjpiOAGRXYC16WNDtF4jb+pzLw8JXQdDYALnN3JCvO0i7RUOyMZeW
1/K1Omy1IRPUdHNnv52aL7bv7AzOdUFRrO6/1/jtqWnLetFhnaT9ILUBdPJREjZ0
eim17h3advlu/dq3udzq5/LI52ZH8HmSHmbSjSrSE3O/aKbyfAzMoqBRc3EoOHyP
MDF4wysnrtH0LrrZ8F67om8TUnvg6W3IcCkU5lZRVi/MP1FtpIw8+OhQowxNUgmF
CRjeCpmd4ENzs8lYl1Zd9AH+rtHza/udJCENPnQOcH4fvPvW91vE8xFeeVLcZXMu
gKUSDSLXtk6z7Ux5NevYr2kdtpXhJ2mLbV+aUa4YM9wOPDthqCQbow8cZ6NaZFLp
r1zoodQpTIE8Vm1vc0LI/ygc2sMRf3TkeEfQJ4tACV0ioibvC0CkVkFKnx7UxGeL
mgcn6UasNjGzYOOyjkckxk8Q1vN/vxmXp4ZyRlOalrC8Fcqg0AjWKT+KwC4cOSTF
HlDd0mINQ5AOTKDTbLEojHbtyqBgdcJAOT2XGKctmv79qE2yAMDfjD55ElOuRgiM
6Ih5O9RZLy5LWzSivDtrQfcP94uVbvOVvbF1sfv+pS4yPXpAWh6W6Pxi7OcgHQBr
a09SsUZRkLzlMuamYSZevhREADXT61GFqn55WrOlPbVxUlr6GW4vlN5Sy1f4cyPY
mT8qavEAcBAJxzE90dCYsSld8prI2v58dG+R7abQ8FDUfDpEwdRfGiEyLtbf+FqW
70yG0rArPfA4Gg0mU5XxnLBRhWaeUCXQHqm+OegncY1UptAmnyBUsK4q2GXQMKOd
2CJ5hwK+hUrf1bnZhTDQOcuk6Nd2BImXO4isQwnonb2rAxZOUjVawhG453QTalMS
B2uFgkjBDLpFD3VRnkqUpxEcGgE3uua2QM9Dehe6SwV5WL8c7oLZ1e42CZRHOg6E
1PmvikMMTfytkFa5xdQM40Ouet8C+mGigMH/UtWxQOEP7U/EZuQEYFsUhx+6Nmae
GK7jCLgnq78O6lc9a8ftYRXPYcnw3aGqm0OIf6dkIcyw3JJgNj2gDszNhCmd24Um
iig2Gj1li7sM5tm92bCiDiZixw33P9J05zZEevxWVNhDUDkAt6Z0jwCmSu9eBtot
5yLTTKgISe47lJKGaxssTc5FUHYWoIcou/SXi+5mmVWAQ2ud6Outu7Ho1X39cdR5
cMsNF2MxY/FXAyN7CCw98mgLytR+lqyLo9hizBKKi6/fhudDtNwwy+lMoY3vGU/r
K9k7PJlaaDNBK5PLBik546fcEKQOHWonEXXMQ8jgudeI3BgltwHG/TEhpJXB/M7Z
6tzxzIiY5sSJot/eWWwmOkfgJFUN5zl/uiWzE0W6FbOLf1NEpCFsU5nPf1nsKp2E
amQGfIe7TFGKEMFPPd0x7CyLDOUuv+TUq9E3D8qfotqbIf9IFTh+6MKasjFQ+m14
8SdKy1JJnpiZPJf1n3J2hwHCHheFWFz0Dr9tPeH1fQtNz7f0D8BvpjHipNQVXEHN
cdSHt0DO65TwxzGltlienvd0umrmsY7PrdI1j+NeuUTokKJmYRmpjjLIcpO9gYNt
8KhAZdvhvupL/j6mn7cl7wxQF1tr+HLLCf6KYTWoRKvwQ41oI+Dzq/mF3DwG8P2m
6zz2csYYRIT/0ZPLNfcD4+dNLK9Ed8eR/+uJCMmtEpblEabomqOCx+oxSltfD0fC
UfTnEiNB6pcjAqjml79Kaq+dY/as9bpHcROxz/7o6lv+NmwpBmtRc5+pdO8G4zOD
qVVxetLj1ZdwcVPdJsV8J9go4N81F9j6HUgGWYwQS6P6ps90NcjPlyXW1pAwke46
NRQtYM7DIwndyEO/KjtgVbFTo7xzafUuVSkCCNvS27pvbFoqcgI+AlSXqdAdj3X6
wSvI5OpmLBpkwIG6f6UlMD84CL9qtKaEvW7UXkvGY62mJfGLYlRcJ8kZt5VQuaLc
cxOwg8t/v5qpzBt2KehVWQkcxkHkQ3traOqZ+h37sEvV90PXz0dppTvghPuKGd+5
LkagNn+ZA9VBf08afSOlAUSmgXS8iL4zVwBOcWI+Zcx7cmS7Nbt5irJE7sJthb6n
MA/ywz3hbaq3VkPSBhLgIHpAbv1XyJZw9DRIufCJCXpjiSdOMhMtv/Kf1E4x7pBJ
+Gv4Ecg6k3erMb4+wLdxmEAusG+RhSLvxdp5r4Hz42JS6cw1q0ET04s7zNn4OrWN
teLaK79WDa9HPmfdE4hbrCbCnKOpCrMGZlJgz2FH324nZR7g+S72qm+60qTcZrqx
xQce35vT9IPjx08Nci2PVp3EGR5oRijbh3Jf9FjykCXrivNo5pe4nowL0JiVaTng
JPXVqXp/xyOlbNYxncHNr4BQEvA3LKW2104IyNQ1S9t3AfGtOVLU+fdD4xmZeB3t
gHSGdIejc7PpA2uRJP6e6wQeZQyeDa9RFW+AskQEsES0MXM0B1SOLU0O8dGBT1Kz
Nw3GBigiP18XZTApDdd81ywe9AnI6o5UcZvkGdLyHvFwEW42x4zmhigukkG4iZKN
O4l6R1/I1q2pohhSgYmB8iHpTsyVWvvaBybvAz0VL6uaD/5YSWik006j5Rc9wVFc
oF9DUpTRzSwKzVAPgAZZHTJdt6l6XdN2zmaMWjnWdTv0Ge3kvP9yq5M++j+sdgVt
5RfhkZRiu+7zicXZOFOK2xhAYGW0BfBggxZ2B34vvP2lN1UxdP58R+s5UcKv03eK
UzI2+TwR7HYP41pnuKKvziSQdo6nnQF1uw6BgpzPk+zU4Aab3ljLjj+jsXLLTPXc
aoUuyQGFP5h34mOvRMbdHLDoXmLipVydSAztEZ8A3dLMFDSyVgu16lNGkCSy6qXl
fy4oz6oPkE03Axb/aJPMHTfDp3gL65+CwIjVhcY8qo+aC6oBQXkx5JK1AoxTNZIz
rq5S4Tmq7JTNKpkOYbpLmQELEwlNAcY4HcNpYXzQFBjCUbZtYYxx+ObbZDJq+bQt
8EkKyyCVkwpvxnLxxiahyXHoZqEYo/xAYt5ordJxWbpWOuIa5NRXIYblTrwj7WH+
xC4Z/LHe+g3HkvGMd3bdh5XakjOVeetUBDPV/kNo9CbTF726lUj/MCY6+XPO55DH
vUx4raxuV7QzErWmLzPcA9urj2ErsOY5/67Zf8UTmQIlWsNsMNu/mf20sBrAImeD
g4SLFoSdoL/jDFYL/FdGCkk8vBV1KcVg8QlAkh254VVCrvs5xtxgq3FSoGQvZT1P
/UNgJetX1ckd+2rRyNftC+GMKZE0WgytoyihePJThiXJPrnh5jDFtj9RBlOQPvv/
QjdqjeopDdprcLlDjddq/nW/96TE8n9wnWNP0q6VsMNzQmbkOsWtqtSS5O8Dzlh6
KmNQUAS8qh8mlEehsdS3fUnJ1aL454PTizdufh/HC7Qsslt/U+kM9Bn3pvrigj3y
VfJ8EOLwW41suwpAYqtAlYqbZdNJW8IdBxSCQE5aQQjGp5OXx1sQGFfm9/fdZbyQ
DzHMatGoaEqxFd4FuX+/YcHHlw5jKYjGxFIIrx/WE/YspNn1vdAgLwbS2mjKBiKu
g0zaLAHWN1+cKCwM0wfuzDsx1d1LG4zTgOBKpmFw8yH4vM3Ouvnn9Z/f11G1oRoP
jNQxR5p/CRX0LLYQ7Q1HaMtP68E1blCCkBTkBO8B7m77rGN6VbESQqxoU6n2bxKm
3sCyjGeAmng10hFid5wwhpsUaZ37IX5Iy6j5R5pMpZC9zMbtgLBfx6kNGfg/fZ23
w73UdpKqEDMhrZz9u4vl4K+764nWhBD3NIhhhm4QgWu17LjXWFXwA7tziA/Q2oP1
7M/O/41j5LgRgaF76MTQIKCKKquIkBiDG8Mw+h56T7S7wOIl94s5dZVsqpj35Evj
5d7gg0s31zLhKKKb9EnEttUYbx6NLNaAy9+iy/4ljaR3I+X3A1Ai/JIXet1H99dI
j9gjCdwOCrXVG5d9DVrOUEwjblBd5/XSvuYfGCOk2qxwMeMt4g+8JM9dAS33lhGr
Mzp1tSYO7aN0KH4yi2d/QTcsgg1vCCJPRPdib30EtJFOVdJIaTg481ejRQ/sNTtz
cEpm9fx4dnUH7CgdEJssSUo9Qn2DMMialqISIe0crKHeD7sm0G9+SKxfY3Q8iqMe
1gxvx9VhIivj5Kp3eyStAbe2K0q3ZPNOZG/NJECH4ZmqQY46q4Uc9CrB9jta6Eoj
hTPBeA1D3XdCBp0FIbnzWHxqNWX7TxxcuiDRSkpCm/T4h1onYIwaoOYX8OQXvSzB
WNwdQaAz2q5Rez4OwlyqNgquAhA8LzXfQPniBKZ+2vT1i9X2ULs5VBMCmdKBslHP
sapbwivqXTszC/RhLqELMylOGIGSF1b93JOu30rFQzczj47Mhwdtpo1T9oxbpvnJ
pb5GMoh3vfVGwkd599ej1jjrn3wjfasNjMUSS8cikGRwJ+dbDUMa+j+rUQdd5aTc
jvefPwWwMbsVbY0WkI31xTgqq/4kZFVsA3axWeDvnVonYc3LDjPaEHnwz7KP4ogR
Xv8hq7nFaljVJGRls9pp/tDkvh4JWfeWNG45GhSXVEg6+suMpOmuIrOVPYALxpTY
r/wcRoma5h1g6vqGMrGADvIKFfp5AKXkcG+G868P1Cd9s1VTtsU0hGtEg5Il7+y6
2PNdw3wmBWlHTOTHhqurLbAjarZTsrfnvTJXyoDwU9E9eflcO7SMV7yN9xJAOxRc
cejKMwVb6rAtERABsnyd+4sx7PvygwBy03jaKXMLaHpc9FILX9HqZPe5LmrJ5yGM
qghodgjXZrXdem3VzwO/y9F7kVrw6RsTRs73RHDxMz3taXoDVDRMR4M2+lcQNgZe
EYk6D3x7l/MM16JTL/octouFSJHlIjInFGtrdkNrl1+yFt0a/OkAep85CTkd+aXE
qsaegE4l+tbyJgVvjdSbIkQAwxqVu5WYUSh/LczzoLpB2DuC312bSS5S1eVS8XsP
1sm9i/TiXtUj3SKi9xAsJqVCzVjGr/tsERBOppOaFElb+2I2wA/AlCrjdueDtGYl
Wo5ZAQ2OQZpcMrJMJ05PQH2gAAb1COiV3i/GVTxl33CVH5nXFzJAiwj8P2NLbhon
TPdxJ2/+3EYaG7/N5ekt6+7ptS2zUZrf2V8rFlg0733mfvb0poa6woV2Z6PTaMno
TgRo9xtVxolaPcvxqt7XRttVNFIZWMX6ybP9whE69DM4Lx2yEUC9u1b+z015Wpyp
eU4g7fJtCBkTp+oNSfj6+UOmLErSbGIYc/+52dn8lxB8OTeR/bzEXMf3pXUKd04y
aNzdncBrHFhsJrWXvcGsHbWCnlNxsSePUVYsZzwboMh9ruZxka7MeA41Wo1VL4lV
vff3yZdR2db8kE5aXv185kglOwO5TqmwIY5Mucg+nDQ3we+4tOl14TbQcvVbjln6
PxNd0eDtHzNGno0Q+Ui8yjpwRfnDlz60FB+JmEQtjCb6+TlVGRGudiPWmUUqbWZI
4ThwoM5gIDGYHBOwzQBjLChqkcVip11TXEWgeA0Oxhbdh+p97QchWacGeNQb7aXz
ceecTKrDZMnHfJqtJIMWzhjiyqAvDI/XPuX9Klk1v+HpbLneJM+pGReg5VgB7mjy
XRUT0lyFDKaNY+6GUyfS5swhsH4VMO1nhjYj6WBvoxnkGSNJdBjSv1zP0dHvuklb
LnaED4WonOd/oYhY+BUj0Hex+PRNBMqdLUdU71uEF6ov3GBy7xYqHWjfesPXisf+
UsdfLYkGukcBCO3BhSW7aWcia+KPCekHVUW29TONTu2k5nx0u4jalIZlRpPIqsBD
8pIwG2PCZc4SHblaeIZekBDJ4GZBCPr4zYa7v0TeG1Eo282ujIChMHVrgnrgdOiT
HyXYJNLrDpczt1uMWwOCWBfyKytS8Q83aBBioYdkGQtei0c/AkzG1o0VNeOS/4rB
4eqh/45gMF28rOFw3cDOUEWP947e60FjfqLrx6B08feNTvks+1JhikN9C377q3De
8/CjXENpsElbpvqCLX0q22Ypqx/KO1/0yrKzPif2uZvVL9sBeOw4U2bYrP+2ikue
tzMWKiMvxcB6lQYjafNsYHORTKeo4IRJIgzrzOimqlU75Vjdx5Q/8GaqXCme1nQ+
TmzFXwgLcP930Ywh52QIjBEUqqvoVOLGFwjdw/iZSgudI0AlAUFNHSGi3VEUSyy/
ce0VjjvHGJ8mDBpGnB0ho9oNE0ZwZ9Q+D2K7X48KYQ7TDZYtDu0s1qqM/lSFFvFR
GjyHRjB3IToKAiAbc1wigAEn0ctS+yaSVZYErDRnWSXxqFmg5zV3L8ojyH1YkCJi
EFLmKG1Ql1apULT/ahmm1bSgiV0mnNCThQDE4/mWACqY/xtGG1BOFX8N0h1J7fOk
4vHrwYFlqg0pQOE2By1Ox9hWDeg6deUtUPsXS58NTA5UuoKTMK1ePknwXza/tG9k
9tvo1DAUeSPCTN70/Vd6z/27RzwPNaXgr8z3KJ8ZD8TjV5Hvh8isByvVmFBNghrR
pky5pOnY7WaD543oB86VtgovmGlG3bAjSTdgF5uGj9HZfCe/YmpvYwgtCCinkVLD
KFCK59kTZ8UxodLBLel+sQVWRT23Qqu8FavbdwTqaCc2I50sZlf4r4/5KTNiE5Wv
kLbxyNU8W+kISmofE3u91a4B8Bj6ZcYCAe1BJ97PggD5NGNMfbeDSHsNZuG/D0Vj
U9Dc/qhRlCuuERAUWKANmttF6lvd+0hIRxub0P7AcSY+KdFUDWOZR/mt38WWtQKH
PsnJUiDZ9+3sF1Cm35z6KRM+vHxRA7QZWVt0ajH1vczNqKY4Clvutf82gavD4oWb
cW/oAbQ6CNiILCJnJZNZ8J9o5hNmJuxC7rbSbTyo2V0cg6o8m3LJXlhSFz5Pi7Fm
2hXlFBhzHPOcjl5k1HSrvsFfORThZ0Rd9zBWmETC5XOYl5crCBcTfhP8CRrljU9h
HxuWwCT4c91XboDTWkDYPgtNtc9FCqNUeMj8wJw9QRhTA88RctTfpixOl9WYBTJh
zdgA5xd31R0h90IxXQon8SpLHftU2LPgIBRJ5b4xlLcESn4xZ1TMAI0RgsyNJHkh
p7W6w6ZOprx1a9Q5U8M0eX6nwWQ9x4TX5/4Zf6JvGaTfzieV4mOOTCYB2vXYBlLM
C6iZ39Calmi86orDECQCImZ+4ICWrVCrWREIqD8eaxk7EzmVhAvib1tAComf3nOf
I5KgcDz3Jx1UU3nJHmsbYkT/l5Jz+tcbEBfpRs3u0LnygeW3QsorUEPw3LHG1j6+
u/VTM/egQxcIyLTU046q3Ska7B7YK2ivRCI6vJ8zFkvhVxysrYL5rBLhiuk4CCQJ
jZfGZlGaJzWtdhvuJ7LdF1a3FfcQTIVgtlqBYAall9jxrGJw2VeeY9n4hcJHEFR1
loCcQBd69BuMwPMQN+iUcZYcnPHz959AI1N0EExusqg3IJ2mgZkmX7nCIqOXO1yP
4huOzh+tRpRBHx+T4Ev0xEJ1gOSlMiqReXpiac+HO1nqWmrPa8Ej1cu4fgLVMgST
GIDfo4bVQav7jEUYQ7rJ2JFgkud4pOcS8ekBMu3pST/6IJ7jI6g6WtUn2RFwlrdw
cOLZ/qksP7tBIGvvMfjCevE2YqzDgW8wGGBIT55Z3gQT+9dsTKhWRXs/79qq9lMP
9ntVB2fBXSKN5tIgrhqtTX6k0IP8lPLrNr8VA2NbVlB3Jm2/+35dHy4y1i1ADLCr
5vpdZuhHM/LS9MRtawerRteMIvRomKx2q30qy4uTooyIE8R+s8gQq/6W25C8QVLw
yLuXDf2GlPBtuBwqDY+7k7kitR7noj8XdiH/0P5B7zZzyCnKB/gpQvi+87Wpa00t
2PyvGnvM9EBcQqYmyAlXZHLL+ib2WVKVW7s5Up44Z8ok0o3Qdie+UHdB1cBhCB1O
OZaLK5T2n+U2pGYy5/6GgOPfMr+TGP3udY/FqqK+mddjwJifMDMxr8xVOXbYV3Yv
mLHUWsTDCN//f/PTAoa5uP4FpzawLn9DMC6vqkFVXg6GMGOQJnoyORdPSWt+la8M
Pg4hqMScOHQMzn/s0utaMNdEbLSC+8VXaumpWY14QS23iqTSlendOAj6NmhjOu34
q9ld/VUzstTgRPbnKyvlQU6KfwMjNojFHH6wMhKAlyJkSnEISPx9vAttXT1Ee//h
w+B4eGdR1q0UdmosacNTBd57SR9tbzD7WseL4iKQciojtcS1oDrKQRWOJbpf32aW
Hb5bPNgNuOldGF9PUOT2kh1xqHdxt4M3IIy7TyMAnysNTA9Fia1xg0o39GxEIYqf
rM1N+B5cjb4OGm1dtE2V5gSpgKA8vEjH1S3mbW0k30VDKfKyBQCrcYUGgNVYCKcA
zxlehjqpTmTvQITi4c87geL5U5GqTdtOeu8GKIuW70VspR4x4V6YIbDVa36EZX7a
8TcXGvAGYP93R1JO23zF4BCC5TUWxHunuaTzxRJqzeMdUXtS+ootNg67Utwd/lU8
QlsIWty/UtiyTf5ZSSC4LM/3gKdYhYrp7D8lm307juOJxGw4f4rBzD1Epq1uxaT8
hB0OWWBl87OF+oMUo0yUtwnbEPgNJMzNm7AAn0jYPPLgZpVVn4ZggLxoFDC9vugl
fIHvpjd44feROxJhH/4FN4E2prUIewkwv5buoQWlYe/6P8RJ91euajLpb9sda7CY
gQV2wngMlVyRwoXqP+hkgoofcnL1Gy5eni7NeGJLlUKZQ9r2wjeMbKFMbOEeqo0T
8ZcnAzlK46LLcPN/5I1mq3X7C5jFT0/hJBEWVJo7xKd7rTjs6l9Wlm7o21gmGjbp
HV8XZACRQMkewPz5CcBG8DtlUnEZK6uujdCW7AhDS3g1jKdWPnZhixp4DDNOENjZ
krFUO+m4axqg/U8SCzuEV3JLT3vW4p6b49IFrU93L3aQuYKPmxIW3HHJA1191j58
o8gXnxy+3lrnvCqeZqDOSnuNROKGZe+Ecq4eEEI5QUAtLnGYXnkAs2cjgEPKseCU
eKaODHYLiFTvZJhAfFjILPTehFnreMEUVAVjQfq2++o/T/qwUKwI1RZzulRyadiS
5v5d1dPw5gu+FYZERakfobBG+oAI9KisF2AtVo7N85Z8GrJKjEz65UpwU606593h
zzorPWy325/GRG50UjYyaclGRq165uyQvzbPQ0+PY1yx6wqE41BmHyzHItLkAABr
EsozQgENOi5Cj1DwwB0Z6qaA5R1XKpkEO8aez08atnG0ls3juGk3elI1yP1STp9M
GSziPPX+Zb/8inkPp2sewlKzA0RROT22/peoH/uBvnWx87Lhj+E7ZHfF2zTRMD+/
1W/+gO2ZYqluB7Cf/NuVckHqDRYNXPRLwAgT4S3bclu2nk93uCEmgviiBpDeuOcf
JnsY/BZRUvT9oHLJSRdqGN+tIxO+cVQ/JAC1cnl0CDmqjFkDQJO5xlWrfv/tP0J0
+nIiDMxkbvGmzChwsLNprrtN6FL52tq5FDkIy4N1DuqSwov4fHFZS/wLRxqxnlww
VLhr++P2WV0cXl8w5vSGQKVy4me2SANDBi89VrFI1sfAMVERw4LV0c/iX/Z+C6HD
2uBXXauDeEWmIQkU+ZKoJw66HOnJ5lkhA7S+6U8RRXpSWM5Zv+34+63mzPCgxgR2
ioWno7uba/w58bVv2/YWbAluMl9fcuIqS/mR0FSZiAcAUJV/UzEsij4Elx7PhEjN
C9utoykQ4SdOchZzIYyM42tAxVYaP2lB+TAXKqnnQjBAofZUB5JZHuyIYzfJV+lP
DroYVUyAaRaukxPC3sbyFt7P/e3TxsWHiga8zaDfF2WCFzDxJ/KC6jaekWlv9g3a
HkXw/m92/qXs/VyPzzasX0KY+JcvprFW8fdPuKoNIBqF/Ed2xpZAoZ/g0Ur14rWz
IGzX2UcKUgJsrZJxCFEaU+86/XIRcvJRE22XJe2/Fq6go0Jmr6zW9TOVVf4wyIE5
2TMe5sVS0IaP4/ov4pIPFvrq7Ut8neTX03GDIAEu44J6EHXoJzaoCJaV4z5FPcqP
JaAsDQlN8EA4ri96Phpg6DWo1LMICOUmt4HPDFbYNAbC6UW2djhVSnxyJ8ojpsZr
Lme6GKRA03GQGsizv0C6Fn2uftZWjAhkctOUYnO2YQsoXgVoNk72XRDps4K7e7Tp
KVZXM+Zt57ds8PbaZgj61evB0jVefSoiruEmQgW9n4qClYut/eev/j9oh06xwygj
EerrtZRzic2kxLIFOeB9eGYiaJ9ozLnfqEuzUktywOEtexjZbdLm9k9zvRh5/sx+
gd69167f8dQWUIWtH0UYzNWFCcUt9rMDvL60AQnjq/aNUHwm7Qxa+GZI5Ci1hxLv
TzBw7r5hK64tMGDTlkoSvd2EA8Dl/REn25dlX3E/AbxeojFlHjRZl0b5B+hI7+2U
nxWQvZAFPiijlqpWuT9U+Gd4GkhEEoYTFQi0b3kTOtlLCo+TCOZoBNeQXg7LAHJS
o5lUNKnQrranmnOMZKjHXZwBooOs3TL0u8yDsAj3lk0c1ASKa35syZHktq5DOF/j
uf7M7Nn/XAGlmRTrSpn6df5YqxHi15BY6UQkfaHgIw3IwWSe0P+gm8lFN59bA4Oq
1PrN4+zDbfEiaiBacGCf3ti5woTUxwPDjx+YzHzMRYwCOaL0RLykkvhE+bmqJ1He
EaSmKDX++cXS4DoVYkhLYTkmPEKosMRAQoLSPU5bwv2KuLkgnEJNo6Y0QgFxmJ4Q
bXNnHb4l3lEXSzHHfJzUqkfJ8vvqqw0VPn/kBiyp+pzMKvMDsz7OAFWPUi8nudpk
f2DIZateFNdgf/sXdatNp0XQQTPdxSahsjcro6Z5vQXwJpzszuc4Ov8Ps1pl0PZt
d26OxPsu2wA7d43h2xaF4HFHL0e8dovPDaa1lgFrTEwCouO+n/jZj1zXIoeJ0f+h
4C/+syRT97OkTfAhEN9P94Ea28Vx5xE2bH+w0SJia5uDFgfsj5MfmRyjQ4ccee7N
tYoD2TxolRMkSEsA10BfL0xLPXkI7J1KuEGGmB4yjkK2ZjPYv2bLOWcwrOVTADRS
AZCdSHLd9IXrWkEEwEnQ7A3HHVYXmAPMI7PA2tjoQ2AYRLco+eo1yoXgaeQSOm4Y
AGpQG99DnamG8gOsKf+cZbN100tWFkpLqWgQSvEikIo+VuCB8VzN5eH7ZdNIdF21
ojdFStUNfCl+bPv1DNVPbc60HDassASOXKbF5/2xbJ+wGZjWSITo03sxeEu7zoZP
mz2Bm2fP9vnif0p4uxQcDTWqUrh7zTQwVbLB4XffW09wYy7FjnyOhJyApYuKlR1m
ssl8+OOok0XeMKxuhdsbxJVTjSSAyE1CYRByWZgwikrEpaBatSOAP6k9JH6Bltaw
+WKJGI5OKr+d893rdi38Hw3P8XMascva5UbOyqcK9f/U0x/gvoRHBiqPDfoQ9byr
RC6bY4U/7pwt2J5/eeRF3EBRpS/o2ANJzwcs/dWJU4yR5VXO4qvflQu+ENksWRFi
d2OuUzcep50K1aXQss+1HJydoIbaS2lXJXIF4tP9aRUHym+rEtIhjyVPMbhmlXbX
/ZMxZWA8Ib1gpCs5SeiNu7RQ9/440ZVTwAzD3zJNQQ9jBoyZanXjyjz9Zd/DgJVO
dUn1mFIj7/Xrk1yxmGwqcRP+mdoV/OQWQHGPqQu/eHV1+53KsjMGdQUmb9OWjrcb
EKAhVHvowfhCCJdjNIkK03cWpiCenaDHyh/NipozCqosvh117pRAMRE4PJ4AXiZG
21pe9Cz9dqpLOUNbtpuL0khIY7z1mIyyYa7WRZ3qosN53qX9wy+wnjRhf24tSG7e
pI/tJsf5zh80crWfi2qzUgTFS3Xz26CRYS3i4tdUPzfjl5Ptuk44Tvvyc4r8oRk+
Qvm6nP5wgsQpece5QZoxKNCX01UTj+VSavl0mr8Mbcw0NEbed9ugIkyiBV8dwzFP
aGCgCBglY0j5X+fl7HlBXOnSRrhpcpTzr3cnPcf+akt5oQGvZ++AhFPd0SHE1GGt
kuexVtTC70Riyu5yAWxnWLhYYE9LV0AqIq3thdh04AhR73v/I1KRScZdiCgW76m6
Mg/f2aRrIt1wRdQn9ULOHNExRFZ+sN+PXzo0bJP+whTJtmC1o2X0xbPglKHZDXQY
Ku6kb3iqswRj36BnXaa36Hm02YIaRUJtcm9s2Cz77s/Gy+zGqBxgbHTMpP6960c/
W1X7eHGlur8iLPjp6TNyy9oepQEtbFL3+Ce2h0O6HfZtBEhC6x9tS3Tou6HpUuBi
WFMG2UjuiavMmceVSpkkIQ/K6S9JaUqDsxO4tNiFIrpGNyHpkChSIV0SdRvUnDAp
3L7l7No08C83xUXEC7wREYMxwla/eCWccTx9vRepdFgjdNO5PLrBgW3O8Qw3KDe/
07em0kctIWQRIRrPSAy/XAvvA4qdCjQtI/9vl8za3myQwEKwYKuG+qMscmt4fUvI
T9PEd0NW9fSmcam0lNFvcvnzlq8tZ3CdyS82OpkDiSv2t19odsdGTSC7wjUw8tef
`pragma protect end_protected
