// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:05:44 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
YbpEeouv2yjik/ajr8gpC6fn6DRuKWmnvACa/DJ1ENnOOidb40obNZkfn7Z2PkjZ
t+uIN5h5VtIG5R2FicKsFIPzyp8Es29cNFOsHXKrS/UNLG0ETYr7GZAkJTbYDUt4
nhfYoXCpSMRRsyCQdj2txUrFC4Qggu9Yo3S7YEqePqI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 31664)
J8RqR7jvQov6AhfFta/s8lRW7mcnL8w8eaCVI99IHlRVr4uVKdzsKjyuHRPQFDar
tq/KqXs+dgg+5hSd4MX45+MDv5cbABxhhxSUuNSbsqEv6kMyqUjQGxe1p0Pth3tI
eyhd2EJn+rAFcSX2hcjr+W8Gxksrx/pqmlJyyjJrSJboEajK0zj6Xp8hRgFrTiQw
S/KU6s5b7nft3bb0yCfqe+PJNx50tihxBIgSx0lC31Tyo25yPhROgbCQJecPYVT8
k2zo33tHY8omFwx4KRxSGTWeZNMXqXJVheLZjQh+8F8Uc+gZh7lDnFiGLE5m1eDz
NHvFIttyFGm+7//BlCBvodSyqchaTufTT1zAhWRyEfczp6sZZ9O3Mri8Qwd/cBMy
UagncLtxwWrGEPRtaAdR7yt0BKrM0+jbmtyVTpBuSJlsw7eb/RpIDm/7l2+XKOUh
0FMO0udauiq+68s7RFicmbAqPasU2yiNuqVwRtTq/QDhNM/HoPoCXJETlY8oDHGS
24UpJIQ1nIOdYe306iBvhphsS9IpnxHs+WIPkHUACYF6cwvCd5kLDLiz6p7WI6lX
HwV/JptktBjOfX7kcKzpAV6m1iSlkpatC3FbDmtZyQX1KSMoKPuZeT3IU03WeLxl
rgDMuA+ZTZ2/TLADDuADa32Ng2oa9DrIK5iY4VWPZkmt2er5D1IEu39kSD7PjiDZ
9mF9Jj52mkJLtLo+t7pErJcvgc0Qay2QfGdHKslT4kIPXF8IFwmbuqR8LdW22Ijt
OwL/Hvy0/A+W9yK8rlxBUSn4YefbexGdmimJOBA3SMeCNo88AxRc/IW8LNgn+/j2
nfpD4qq3hbi0FlaEr3vodT1u8lBkxi7shajpvksCzXnXLAWzlMcCn2f3H8N/cjsX
ErBlxt0vuRPhctalN/A4y+RnpSs9y5HYoQaP+zwX6mFNknuhN81mgs1H2YMYlFM9
LGvrAaS9D2ir4c5ItqBKBKI9GwGoaO/TlMYoybINFBxy55xPLodnvJkoygcemA/j
TgPrhju1gF67r1rVA80kyABMk/ErGPSwQTseVu1du38olPvLxqLavA1vbRQ7ZB3E
tRZfg5Z1eKKmNjCFXEJJ0h7eZKDZbU9XgyTNQx8sfUIf2dJNqWTYPmnfA5mZ2I9W
eCWxNMCEkHOvVibv9+WFpzWo4Y83OyiFhv+4mp0KloMHlJywEhitUslCrN2Y0hjZ
sREXMg5vG/mLWAQjWiO+nBp/wcAi/2e9mRIawI5VBK4/MIN2jyM8oyGgpYfhi9pz
urRBylhNIdGSiUr/LmlzOz1GZv2izYBO5k+kqfh2EhuM3jkSj7keHViwhGefcaUa
YNpyMHAsW9q1QoAP3j9Azg1lzwFTZWFgEjuIHfDv7r3m9w6g+w4m3NtQshcdBSds
bo1GcJ8FnrJWEMxkO0/iPwCOZAUBUnJTw7wQyhXtikc4BPv8VVSSC0hvpKJlMRjS
rjhChwkR1bcHQKSPgIXeFQnfYgyDginSZ7Uxr3tR3bGZlNThl0wH4cMCagFCXJ2p
5otad4wOvdPSCF/08CaxEpyMx4yGvlv3za5Is9BTKoU7Fi9LEyJogHRjiLQSHGhp
Mr0ROE/9ZACvMK2a9Tvd79g/YjHMOZQbi9HtKGYNxQvaocnym2++u4S7WigPCQAQ
ERNexH3csgNffNtOSTw6KToGk/A2tXW+Ga7pn5HxP8yzCY3azBZYa8VNh6GW8iDI
WS9sLbUvqt7M1kHNSZxbjX6iCDv7qx7pbgEWKT2s4Ym/ytOTnX43mhvdUY9fG3s/
jUIE2ruNHpZ+HisEnLQ44Yovd9M0pAFEv0brPAR6z0jYT/XvPG+iGnSiBu6+kNnk
SkFf5dnucGc6bVSTwDizE08z+W/WfkqZeufK60GVZECsRccI2pDULc0I+38liLP4
mfCE70Dh4wYBS2+FUiBiTLQj9pdlq7T4GVUTS2NSnjQRyLvnFWlFW6+qQlRExLdV
VMrONasWkWXtgei+p6VutTTLmTVYwy21sBUxSpA8NH+iLlkkg2bSUiEjv+OgzE8J
kDe9/BKBBBFSuCAYo1ysb4JX91Yc0WhjmVyFCgZUx4e04HDl9zmwcoN8mTyMOgQZ
3uPc6oO5pN2MU9d9GsemBohSg7+vY1TQCeDRAPl9TzSmeXKzKvE4Vqq21vzkNRKs
rkOdA3Z31/2z+G28lDyH7VP5VHNTc5gTi48A+dH/y4FaD+EPS1DsqKGxNAWDW0sy
VMHZHaBYtu6M+CGB3dMMHwGx2byFqhhWgv5t/sPzt9i1wbaoTXru8W/ZPa7K4uO9
kBg20bCMVzhc35sAFvhgmqEH0iJOtxEgXZ61pHPXTWQpYCFOrgx088Y7kzYNymPO
cxGm+5V2V9wkDiRgBCfsl19HCZ81ECQzP98dq9dk5bi2OdMajck6us69TPR81D92
tHmdsz91mhVwzyuEycsn1DY66BMtUr0OoGLYtn4ro1YC67GX+biG/D0rK5ocoSQd
LjlP0PKTqGrjNWkfwaT8Q6GhmRCVhJ5th3KGqoSEZBY3Mu3dzg2GTdsQfht5DHBr
C2dbJovAog10VFrHMCh2xlo5KrLe4szxmSD/6g8QQVYpQ3B/YEzE+hjsHBNDx+5P
BK9GrpxA03mADEFMtsY8FE7lKBX0CCQqh+sfaGdm2yrhxvetT5WiRBM7OonTAlgR
wQjXf2pnhFWk+L3eI2lyoMBMmcclqX2ZW2/T3HmNlveNWkIMk/Fn2lvC/lsrmRfy
7Shl+Xb1lcWGmSe2ddQ5QMvjttw58VvC38upNEg11B8IAXLSaMXZyXZhpfROmtjI
U/uMuZgBxeOt3yYYoIl6hjkxIpxxkx5rzcsiBd8Kt7LDOIssIHlM17MTEw9PC6W8
nzNDDAgZz7AN+zFH1b/DVEofVhfyyUmHWDh6z4p4XBJYHRCchFuKnvpHyH8bF2m+
CQTTdiq6YztmBr1C5BLGHLKNDR7+7gGDKCQukmat3GQYYlg3A5SBN+l9TjfRkbih
ZfV+I7o3iqDo962+an0Htzul1PzueXFKhXLxudq/pfPuQdW0nS5RL3KvE0j8X7nD
pxlqvU3hNIbe1FpS1GgdLHEC8HZYz0+egUcntufZltgkmHQJTcRfbIxA+yem88oh
FY5rwps5mhTrpyezjPA06UTHZsx3cr9LltsL4Muxv92bsmXizZeh21jn3g1sAWIP
dEURlHAZWZlnIDMPIQXZirhtSehBSnKXgKTLSSYtuYKc0qHCamygXw22EzHoDOrG
NUfA/RdH6TGkbAVuetCppt6jGSBrjYZnFNjMnSiyezjypsdUB5nQ82tYAf9A/yUV
Xq8l9iWnR7URosJ0xdF17uu2q5cl2C6r5oG9wdonRbNGgEaOUPPMptHsr5BPlvwd
GVUADMc+ac5qof47B6pZKa0c3DJyQYvhsQy9BIviKsOsrsCppVzXykRc+Rid/HkF
w0CmjzayhG2YQ/UYWtDzmDzcfbbd8/i3bBZNlOKiUdb+ox6PLykdSbBejsVQHfxV
7naonfgscRm7hM2wXprqtcKcwgzevqfWl5MEDHNgDuHm+W65oNZKpJP9TzzT7MCs
SD7M+1Bs8EmgbGzPTrB49T9XsJ9Yh2eqPLqmn9kJN68EXWuqoPAgeLBhPERzhZnF
bt3mGVrPtWd7T/cdcASXSUL7A8to/w/5e0L6+RJqh2+iwRfqS9IjidfQ26wDZv3R
HNeO23YYH+yHA1xNLuzcvkNNLaYzi3zNGZ7zuWTRdgdiSfRTOiEF68wGx9CWNRWC
gNPobbN3j7iMEG35x4oBjUqljCxr6kBVZdA12ss1xENSHdN3h44lKZQG8U1XTlR7
EgTLM9nw5VOn+DpJeaGZgdFs2ZGZ1CTfzUEBjnJ/NhCP/bNQkb8l6C1QfMYcaCxL
2sCcAapP9YOYMITcUSu+lU7W/Iere4eaJN8A8xauFQxA1aOQmS74iaovAfZCLMWK
mu7nZ8JNfRXkX3tJF5LgGyeWe7DebqxXKP6MSSVu3RdTYWjpBm2UcH0tlMY7BlYo
NjY0VPlN8ChGPIVtSI6SSBXIFVftI1Bocv7lTaQN9XY+ShbrK6ncpsefplv0ONHE
nvyyOrcd0zNbFvC6TBslYctC1TQobQLpisW+i8S1I4VDFIWGzUMqyROQoA7kd1e4
VPJ58aekBHUlpV8Zce7A7+KcYac7eg5efO5ok81OluArMcy932CB2xeBHrP2xmaP
GbMb4UgWLMmlt1jH+h86DUhcfGYvD6j+gO6PKzWnCbPHb+iGsfjBhJGKh0JQAhBs
yT0zsqoTdwFXnzydTeRkj9okY+fEkHpLuFWkDTM0/KAWeGi59NXAeUfY+TMOpmsB
cDL+tzfY9OmBLkFkc/KOPfejP7ISgX7GKiaSTTxs6PTIYDqt6h6RAhoa9L2Eilt5
OO5hL1EUjOSWKrwULANBOPA36R93HPNVuS541NP/fR4/H9V6rAY0hPV72EsWbkis
YhSObf39TqKBEJB3svcZLHHZnOpvcJ0jrBrEzLV09STw7OCOSUK8f2QRYjIM86YF
z5byUSiUOdZeIihIeZdYDwaz7Jb+gbaXVLwYccchR2C/ANkzuVJMTEg1ChZrLhjt
gfbwJ2z8uF2xwzUZMIsDuZv8CEKzye5iaVM3OWXPYR9vV13VnWKf3v49Q3Bf2WR1
1Ogvfdkp42Qhr9vtiwtBumMSlimN8xZzg6OlASqupYnk8w+hozvR/78y5qb2sK+J
NeclRKgFmu2X0DVOksbNm3HyMrr4Bd74M6DHH1xIrloxVd25r7Twvrm4aotsPeqq
1+gpcT7W0yntbhru7EBHofaNstC8iePwmnd5z9tN4+7yN40wDhgNURcZlvjLs5iN
QtQ9zXQEVuJ7XIP1s8T+CD0RA9DfiH8uCtsTKWtKL/6mVxsWEzlRpxG47rdvVnW/
biGfT2VBcD8gvEvhXYR2j3ZHFPwYPWGUaFjU926gqxjIlVkaAxJQSUSGzLgAqmhL
9URHuIeUFMCWXpY4Gz/fEUT9dDjkWEO54rIBEzhfyLI6iy1GYkD14+aG/6SO7rCc
UGFBWQhf//yYcbLLecJOfvpBQjwdKweZhT+1+pHRIMzcjjvs5fDC4s2uIYVs9VOJ
+GPZE1R8CsJF85+sZf+YG7S0ObwGxOHyEbpVS69ixHYGfNy+ElLYH50jlVQHb3wp
sTCpj7L2KKB2pMNH5A5dQ3QHH5OoHgwQ6NEYsja0AixBCBzAj4P+lQZqbXR5BXW+
BhVtrSMEnsIIO6kqIJPYpGG40wIlB3fVbZFON5Gnf4tPvYLPlqke4xAu7CCZuPvq
oNIPFH7rJSQvssOO9Dl+UeyM7ZVxxas81uTQtZWD92HkfsExXo5yjql+mwdwuimG
ncX5Rz3GXmC6YJdzKCmLANNn18TKp3ig3XRCwjkcMNODi1fqU6P60qN7GAOWMwkg
DiDSFWQPclgKCUN8/z3KULkJuqWkP/Y2QH/jxnB8A6vcUclq738UUXxrvQZvnd8k
+KVlBT4T7a94P2QzxkL0o8yOuE4PIE40dDF9cMklGM/wLd0Pho2afPi0Ohtu8dps
COiHgcH5Kmde+VRSkP04/fTq3+aj7MzzhuSBkx1kvPUp06qgJiGNxRZxJ/MpRPCH
ZhRjSz3SVUP7YouHCUZsA51m/FFhXye2F9cqIFaZ0O1HozvAMcM4p2LSJh6hfdTI
ldJrT5QwxDK+P8NsGaAKnP862eB0e4eIrME1ALnchGE+FiP3cKyEz58+GcWSz3bV
A13TyD5Lpe3D9EW2/MWPbhfqDqLSuoi7dzxmb9UvD2HhkbUCC9WSpRsJ5fP1iJzU
f8/snIuj+jJOa9Kg0m6xbeZ3S6p1eh2TKhUD+N9prFCGniFjTVFGI2OtBF1TbYLv
BxWywSd2VKRvVS6ZjP81ySQc94g3UeUpRcNxL6NWt0cCXiu8jMKA8egn/vcXmoF+
+MhF70x9ZJPBXb3u7Di5zf9INBxbjCJguMWIVlNFDI0Ln5vIDrB9Vjvp+L/7LpFy
KJOm9cPGyAozYMcLgAyUdW2UGfaxx5aEydBNe2oSoDQbFnuMiuLO9j3ZUldiHA93
UHduUWo8avUQ8cVMlNtUfO3yNNiwSB+BZmTn5VNS8O+EU9FkydryozSH/kvrWTmF
mNcbl313AuaQA0WLSF31pDqbwKLKY3ND4CsPtV6QDkaK7c8ChyA4hU3Ixeaay8Dp
WkRy+LXZseCkA7H5jk3s/yaM7mhoaY0H4JxBMfNl1wEDyEpBKn93yMeJMtvuE5Fp
7dScA5Z5ToawSUILR+oAwKIaUoUndTuDUo8t7sgdcjJtUIXi+lXoKB+YMcjlqfKF
aAfuSkxi3LenSaAWFyThNq6zQbrBMvNGKr/yKTgL8c0PblwXTZrJqcUSlXrj6w6Z
bcTd8mki071Ve9Di/wraEx8kyQT7OZWP7vQ59FYWebQ9klNE4Fd3n82kk67EZVQr
OHir8pBBU9jwQi+aw3yOwyXmH6baugtHoRWXhSFqPc3P1bPJJaXZKTl9cI6PlIfS
EtRRFjXgqBwjwTPgcPSqyFRSKHX26ksdBbF0n2wqL8dOUNh4pOk9YraR9puJa4zX
nOls/6TCesnmRihzb7zAtq8WwuS72Kn56QVNCOoRj9mAW6+G1HJlyxmBMInXNUr3
IHHqKGE0F7wiwd/lH0O1bjg732f6fcRYosuwHwGm4Gl3qK1hqnpuRrC9xYRV1Ezq
emaiggClPO682fUCvkuNN67vU4nrgQNN5ZLQQzVyuS/KNFDud0eQCrSsfdhj/t9F
9CtFsqpPXecsgyUrCBoXew1LGX18hll+xogOukCtxeaVaO2EQv2oe9D5+tCJCE/D
ie94s5D7zg1p3hC0ssr8JH4iXZr51GVO15OFwbNoeI9tPci6Wf5H68lZI1MlfGxe
dOw6Zjlpgbnm7qdmBJuX5NWd5hylY5jA5cKb4kgtDEmWr68gtVao3Fdz5QZQU8pe
Eo2ejaNFLBTfl6wiBYOFlyS876koVw6xraztvMtDFcHpxpmKP+klIfkO+NS5xxd4
bYbXsYJbEBTbAO+/e/ZitlHgw/GdFor5H0LOuM9zUvaWJGOnNcXbjUeYT/yKwnXg
BIeEqnzubxJ+zpe3ok6kFteh75OxfqxnHz7JJ/mY1DnaXQ55fIW7koo63COZmXfQ
PWTxXBR8fXdy7H7mLlGzuYoNYxWY6JJ/h+AmMJdriWGFV+DFzgXCw4l/bNv/g900
o9FKuhqlNpP21fOaIcAADzZyh0l/IX8Kkdt7BajRkFjnsqoX41HSmWFG+Uh6CTq9
xkoL0F5EKWC9bkMCQczbOsbIt0WxPv1zllruvFRX4wst9/djLthlr6U8fZPOC3mS
SK6pE4Nc60NrDtUaAmcrbXySVmQOwGVH0NVxGtgQ6OsGVdXdFmvtjN4fl72QOIZP
uOK3gFHCP7lnMQt8I/6jT6eBUEdfKHYEy/JICzUWWB5QLiLWk2+QmSb9WkEzZ/9i
IdiYYumeJAGVGGHnaGaiHjHm5kmVq/n4Ph6FYQYhBM+8njbY+BTfV+OYdxhy5bJV
6a9IrYGzJ+LXYug+/iDvUbE/wc9w+lle/UL5msRZ+R3SgA8/kQBaCRzS+KCT8qww
GSBFz8GM9AUxiUwtpmswr94sZY3lBWtSn/GlNE3qeqnQhjUS/FkKR6kT+3Z0i3xI
egNqjggrLr8XSKBg0xK5bAEozPQcXBBr7L4oCClL1QUFa186iRdv4jhlcl/HS9G1
hdcAyY25Y3o1+P4TwwtS3ii+GqTYtg7BvrGJBR2dZXJqDq5a9j2M0YlUNkTyeWrs
cNUNCyCQBBcplMnDkJbz0a409jYe7xg/iz4aj4TDDrNOHqx4Z8jGPd9qz0U3If2Z
1wEPgNip8iedEmtLB5X+j90L9F/04QjVOVfr/341Rp/ysO5+O6zXIzsBNH5jMk/f
+qKAtYk2mQn1G2phsS6b77RKZkdV6315t/daFS/lCSFQMpa3arKImTuSbEjmPS/y
A+Bn7d7GrP5W4l3M7T8TOv0LOxiGzBURAhopsJejs7AdINHWT6KmBlcA08RTYf9N
JYe8X7RbtGjP09FNBQSVLToFVbBdfjXlFqGZQ0j7hKIpoOH8dLG5JEyrrNsFN2GN
lwT3JLF479PWD+82h3wIOuyEh7ru2RJdjaR2H+Ww+MmbqXR/5lQU4pDFjaIWQGdz
SknmbS7XjoMANxSUVeSNXXWCPsXpzN3aY7ZMdrNOH9JhmLJZCEwTkTP+IyviLLDL
9qqyb8H6GknH0Y0W1fVCFHlWP/JkYSuoRuMOs6qyW7voHMY/0f0CsokLdR+kM23T
N4oaslBZeP8LJXmN5q4VeV3ExmEzn93Tv+xF2JwAS/x0G9hapguOHrCT+aKs0ucj
SaxRiNv0Ri01RRxGpvg5PP0Dgv+tEKzgYGWdTBHyjFnrtSb5v9s5jXu0BlA22Qqm
2o4drQD9z4NoZXmr38U0iW2KiN+G9ImNZTpGWLEYZImg17SEpNGHsXre76YPCjOF
trm/Gg2CMKgDSUGVVtek4/vtRABAmUiM8bMv60w6TbVH2S2j0+r1vECZowhE5n9W
ORmXNI0FrMhT+JxeOQYhwXmc0x2B9ZEaRQ2FvvpNlKR73vunAiUplLm9S1uhr8fq
dnAKU1aqIPgICIeXyuHxCVKT24fnAo8ouQMRLKTALRPE0ytx7djL6sPFPT7MqNoa
egKOnCl2tpq+hY3waa6nQk+42+sV737QZG3o8LAoncFCmzsuO5DKdScONt/92MGj
M7Tfv2r/oD01tuZtEn4XvYeEVGniClBQPgIs66ZVwbWyzDi1Q+vcYY+jwseAWv+M
XI3Wbf76hjFHaoptxmlPiA6cHPU8ne5u9vXtqQy/PyJ/Ubu3CW90Be5yR1zctMqh
kJmfgWIwCXyz2/GRiiil2+uxFnMCI7j59xZxchEfEGb8UJHCEtzbdej00wnsfe9o
s/jkRoMYIQ6pFfk8HCdP20JrUUzT1tilXLhvR39fO+ZaDsi+puIXcXaftNJusW//
ZCkh02qGoULlHagQyfG61fuMLXV3fuW+I5XWWh8rQ1FUvhttsYp3dQosZIq/c+60
0YlRqpRNRzkdHOMjiMsBA7jmo99rS8zZzWW2mRilYw1mhsOE9pTQ8s/LJD4rlA6x
1aofs8X59SB/w29u2eyMkeWUddmGoU4d+bgEO8yOvAJ+jIBruXbtE8U22VrzVxlZ
evWmRUuTrwejgjHEHnQFrDcV/LYi8YRHz+wlZLlIk8qM2acHO5ZYJCEWeYi5PmwF
62VPsU7Qqgh9iY9bzHM+ohNTgGrFOR6eVHb0v79zkcukARQjtE5kfdnNycmtv02r
RmyAbfFhXjC1r93aDodijvCkE+P6um89Dr057Jt2bCtds/HVnYd3HqqE3/loIU+I
WGF9Wcf9Y7c6nLH990IpHfeuLc9vbB4Oy4eYy3GNE/AfYNQ43IgpBrpUKnsA3wxX
kX5ur8D7Yvb3nPekGIiRwmWTGKGqBZktk9orYoFWgtRc+iSvIMWlpEslSCnyHV/f
Ufjk60bTThXQu5gN6bMbR41GndE8u2q5tSybB2DEL6OIzRSnqwfQ1tgc4sCc0VGM
ZOFu+n+vOFxPJFdc8YiXyGo9vs8SIGPl2gyZwTfTRY193/uwdYdZdGZxXs3XV0ak
d0l2Jus8Uspp8Mm3RZdSz4OxNpd4Zy8//pbhJTmfOF+keiQ9MG8z2ISxZb0s60QZ
Tl6SskOFc5ij5h7rDjxhVeDY/5XWN3VYH4UWkJ+y231uySq1HvFTvnWbnem0oTFq
OqN0BBaZ/9UlsPXOIqrlIZmKxI/pUzxciVLdmJ90r8irn0oPwn0sppw/Er+XWZhk
wZLgiSYzepPtvDpJ+tx9Rx56BYPU1avQvRxhe5s/phNZVojrGNoHxE9T26+0Htfi
M65v1PyK2tlFDhteais1kLUnYjyznOwsIXRf6iiYepCN1SQQBV1uPTCc4CWrdF3i
c7wtuENbu+L9pDHtWCTtdIS2RN4aQvYqDMCWP3eiIEono80fCyCHqwBW6jc3he10
H5qinMPc+GjJum5CX1p8PkjX3g0gNuqszfwrXuB/7Zi1k+roTXhnP7+poScwONqk
o7qZLIiMBkW93mIGMEAS5vsr7nW6RJbp10mdvLPcToXDfcVVC+BTBMs2rohA3R02
ivpK2Gz2MfdOBmsNb+nxXRUoYd+BUGWKlqPpWnK8jDc1AXMCSzmFGfsFUByDEM85
VwxsyaWbXA2itfirndvOb7wlJbQ5ZfyDXgOMjuZs5BqVbkWoJBO75I50TOTWyIo+
m7gTH/PhhMmibrpKG24lM37YmpKLqTZ3b77lhv13FgO9YyIcIJ44sbjPRGE928gA
eWkcFCyS+O2+8XSDeMql7vB4Hz52ELjhEw/urSpiuvutBwYGZ243fl+A4lDtfamB
CgQ0FBefZUJGTJwjrdmCIIEeVfGhL2NGD8TItrkE5SeHKKZSLcbiu0UvXWRJqZXO
G47RpB8MnycDClvBPtLM/zJlzyB2D0UT1gJgQ0RQihI/kV5nMOSPmxkWqfUHkauf
lxno38gY0lluRxiv/GDO6RCgYCKQDLM3NSHjaPPm84YJC6EePsdkv00KtG+Qf3VP
9FAZSg7OnmLofL+5Kf0PxduA+6EpNAFRSQdpH8HP1ypPJjPsMokG60bx0OhgR/cJ
y6XFU8SNHFXNSMKUrqqHv5JDw5mhaIrFQ4rJ2GgHPp7WNi4wyj8rfWt1ijmUpNOW
LyWO855EDfra1JAiwqD5O2fW6vni6bO46QF1/ICUS9F4lVwtuT++/sB4c+cXDAD+
R5pTg7yNKrKGase+EXT2qsY0tAJxyVALEVeE0ENIx74RVVUSqWJgHojJPu36MHeG
T+TnULQm2VzPSRZccHU01CWcckF7JodpYo5n6/YC0OEJCa6Yn7wQC6H2X7aCFbRP
zHbQkGj/K3/+SL1XyoHwKAJmXBSuEiqptnQfXUdESyikJpZ5d/BfOFMymx6/AxtU
Z9d5KRl31Nk67zDJRhRGmaxfiOdVHdICh8MnsWuxy06QzScHcbT6XLURvMK3b2H1
gIASF8kwRYuitGWfTMunoe7udhMmP4MVuZYg9uIeklMTp0w2o3fkDUzXHPcT5TZ6
Za4h7K4L3Un9fjAHHf55P+Pk+dTZoc0lqxduM9LScj2Myi2uWlyAhYp6a/8d2xTH
fl2NxTprKLjiwGCoYNJTPm1cVarkzb/jmls7zyGCdkmMzebPyFwlgbbDKfW+wx+a
jM5FYt3qsDnZfbmMBr5MOOsrttydC8GKKjzKUka0VWlJRsHkJcdYa3RlYEZNTbM3
BtgLrZIvzzkOzOQSiyhTIItHuZttjsa0jgboupFWA8F5YruKJRroMdYjc5yy8ZNS
kErgHPRZ0ZuGueNhCF1AujSypu0xcew4mHKF9y1TKhe9Ty5lhOPbTlGYjJqBVGdc
J8Nvb+6AttLOXmEDvnmQgTm7EWwcETuE/Ijbl+2FX84a4OhH7VlsWr/f+rzlEol0
ASA/XWkwkN8W/oDu/l9dFhTL/LSrQ6hPidxeH8AQgKyyDvXWOBd5603xqgyhDY05
UaUFiWzotsHk4KPQskMdgoyXWbyUBrnkwBMXM2vjfoXYeCAgdLw166G3QJITX/vW
ro0XhAwn55YG/+6679/csJvkbgfsf2BRPDScG5GdAM+D6vZdAXzgPhLN/j4UK4Fs
DenokLS+20Vccg5xZfk6a0KUoZBZdDFM6MwLPfkatSqbEAG9srQWxn2xOphAxp9o
teFUlX+5VBnrZYpiNwQGZ84csXPVZx5TuBwDJdozjaqPDGgp9ZfAOOL+6qIsFD+7
wCwexYu/acb65xYX6dLzAjeylx9wKgsuwqrwK9OKgtbsoY+M2S+ZAYnAvkyJHUBr
rGGzC/idBWGcJueji+VleC7I/4MZA7jzv094KNY5A7iGmcVlgvn8LJJPFDytp8K1
P6m83O1TBuOXNukP0Ko2Tp3V45Bmt5wHefU0LDCzRRQs/1Be3enY+enWv23OHJJj
p4V5C+9yxRikUI5wkj5LD6MY3X1Hb5iTfSbVbphUh6osRWV/7AkVMJxnZ6GNcJ07
fVMpb7b+e9IvuWFjU757sYxXee0/6QoWBa019EdY9bs/RIB4VUgSQeBFYJKst3s+
lX8fcq4hBfm3+JxfwZPxjb2BHEhcQwjQgyTgrCQULVGCURZycL/X6llJguTE6IsA
W0j1wuab3AlkFe9KEtN4NqcDdwWCa6qAmX3qcmzth7e6LaBpP1GwMnRPxnLhjvF5
3D7NStfsJ7X1AzQ8KswPf+ARpyJi8T4iHoJD4lWcYLqTKLBPQPS+OO6pqhbM+Xg2
vJplgGTcuIdLx+nunY14bsQEggN0RAr544OO2KLVqjVRpmwiVBU5tCzDo5lsllLs
3uBdLBrmX4lG4LOv2MoKWjwn4XNsFT7zaG7W2r5TFturPDQc0ZjEboiqzfg+LdSW
Wr1S2hZPWl2D0+qkF6PvjGt/H9jHpWr/dOj3IbvCNxcJwDp7SKDpnsRXUDmn0ylc
QtNHy/EqOq5ORQb9WA7WoOn3RB6ZjIBn8ceK70WXt6X4tAJ6erjaPloDusGE79vy
tR3NYxewqsTNSqjygT6FrfFCaGcycTv0nrYhXlUtyJ/qRcbPIxPLgALCnTFQr6yd
ZJkokSsrhFb25LrDJCdi2a+QgVHpXb/9Bire4aH8npMr8+VwdnetXnsBqebwZbsy
N9m6G+/5943vvtyRGmUWQA9WOlPSCLRqslvYb52ZyHaWbFG/JHt5LC+MzFYVIWMy
MNuP99sK/Fn70m77cO1cOinOOlFn2+DQtnmLnC+OfhzX6zJkxZwDy3TGzq6gGEX7
xXU5AIixUwA28HJAUor/AXlEqsXR6Hl17BZwQCegjF4nmMN5Z7B2HHOkMbW/6kb0
vDXWvLB5lcNJmvQmResiKDyHls8nhpgcHznluv2QR9+Z8yZrmRE6/P3aBIUtj8f4
6ciWkiUgNhFlEnXR6+L9yiCiKJva0YqSHhDAqCXkk4tNo6awzF7QydEUDIYCb3H3
L3rNUAeFZ8f36urMEPPBPpx8OltQTvkccHPrGbuMJ8VVBFkdSVIZguvEWp9/D5kx
wwnb0NeTB6a4jnYwIJIC9T0ADrU4FNY55n2k9YkHuEuGiiuyiwaFp7BRxEUxGwln
AhS3ABcgPP5op9nJyP+6tQRMj4S0KhiPIWDrcuf/W/J/qqqoDAl5EKVsiPcEke5K
sjBQ/PegmJaFEqu+EohXcuOOkLDxsJDDRYa26A9260oScsSKUJTw9jtyeZ8mCH4y
5uS3t+sV8FaZ0T/tBE42RfSg9KYoVz33QqyXYKkfukmxgpmsziYcgeRUleb0rCqC
XHxo0RuAp/XlOz+pXu9tfYNwOPGfIDGU7GSJvhDrK/eRiKlSX3Ux0TLAIYsgAoi8
U9l2Lv/nP4SYcODEyjSAodGOzYQU4WHLLwwT5eIVDBmAk3UKrRm1fz8k41lCqVv1
BO6iGyNjnKu7ZyzaKKv2vEyYJ8Et/7xsbHv+g7ADbyFuE/TYSi5Ou5wSwi5Kdwnd
0l/E1b1+QJHs/PXu+Qm4h4x/7TdWC/U5oLFc8tUMCbn76OErLjmddpji7jnCNu3R
pK3BVNtt1GwHMgf8cqY5fm5MIK/gqgNG8MSbnVvLk3cIGiscvBKwqLvSd7o8idfl
BVQ64uZVDFeN+lvRJvxd9pWz0ZS/hAI0EPHQbbzOujFDZvDELSuMdN0mhNSLQbKc
3gKVV7PXWQ/8mbKaUkibFNZZAeWgVUfjEh1/NkaiFBhHVQBH4z/nWol69KnMpELC
W01Vrjxqxc6Tl8paYfzyhwZz2+mooUlXmHWm+akQMbOe6Nn4SMj6aUnuebVqbVg+
W25kSK76UtpxWQNqu8nut07hTjdzyIJF7c4RuEL6zwn276Mi2C9GHrq1MA2tjco7
ArREfswB1z2iDv/uejCc1jI2MdAILLXroCOMtOSWYWBfXhvsqnTAeTTAFRIzCm3Y
iJfNfjgt7vYa/fRt2PuFVPzSV+VG+TVcDcWBMdtFfH3+6FMWmU7CvdtaUkcN9MuM
YE4tTRjiv4U9zj8gY7X2sKptPISm1cMfg6U2ASr+T0fp/D6Nea9XeAf2TMeUSte6
rml8AOe22qMwRpRkwBOK/Iy8gWLLZqN4Bh/tbtw7TIBMzbviNoK/EQ9D+plb7g6U
VYJ5DUyraPIJwENFyY+fG0nGSkFZg48I7FXHa1Epo5F1tSikwa8/C5DhR+ufXEvn
i2ZZN4m23F4GhsNxjLSunMurkcr5fHoq7IWOnocn31u/fJa8argD9bEhmKLyZ6FH
vSiBXkul1qlgmYWt2W2f308zS9dgMorypSWT41jTQFxlNe/YHZ7a9RcGL+Gn1IZC
2Hj8gUoWaPNMWL42UfNN+jI0VHLJ4t8zSfq0njW/hjegltumKkPPzx5Bq0Pop5E+
J0IXyVi6vY7kQujHcGZkXXF1alIVr3tzkwDS29yfLNHhH7gL+h2cg4sAGscE0YH4
Jw227bySzCq0zG2B9jY6h7vilKsdKOQh+HwAqblzcqspuyX2YW9qTWMv2d5PCsUA
AwI4z8I8poZYMosStoXhmbeugUYdp5TZdTXN/kY23R1wUg24tcpvZir8SCyFSj4o
NqrX1onTFGy48zDJrJ934xtVvQqNVbmMkbZmtmVB+1AZPWClfTPOy6qL0eatMKQM
1y/Fi5gprhIn86OawCQEhKfwdBKzfBP3u4HGht6EXXnj2HpIRNBGVc3v/0uDlDEG
NepscpzKxosAybUvfWJwkjCSL8CzsZ5oTBAIjjd/tsjiT5Yr95lTQpD3woCvsjGd
XdSLZqkSwoBNmyLwWmLb3HVGfscS5M14oLtYKItZ0SyreWDS37nhljEoL8PvNT/Y
I0JIXjJLVHpB9ZirfXWSNcab9PaWEE/SCLrtH2OLczYdjbr+3KRIbxT6XgQ7FcSJ
C2lZxFCK4Ijka/6A5MX27gCoV9JDYT38e5T87WfVCa3E2UcGYsjBIa/FTeCj6EuV
b0hQ9ifxBMGzZjPjIGyKX46ideVVg3Brcts8taqBBKUFkhh1HyA5h3dHlEc26aUb
3mPkSGf6lS8WSBPfBCD2s4h3h7GG8+/Gh9Mr3IyOwMsIKXqUN6my2I7XLkW1S/Qz
Bm+RRe4Y7earPy/ViWkrS1L0Dnhlm/ai07oXDDSTu+bRIa/H+RbprlKUxNeIkwpW
LafCHZI1rpbXQaOMs6GJK5iJ+49HG4MMDJ3Lm5ZlehwnnT9d1nFV/WFpr2vyXOyj
Jlipc7J5MyN0B18lRuyRyI6DcireM1B3qkS09ahvU4+G6b6Hj8pHAUXsnn8LiAz5
PLgx5CgYtEwZhrbCzEBfU6KFp5AtJdYMbHIEKh5F6dI0N9PlnS1dN/hTOSwogwxe
gfgJ78kfsQzHBzEA0A1rBcSe1QuHkk5BtgApk2DuVtySkH6NUI03QnmIgskzl95j
QZodh5WRTMq+eWA/0O07AOmZ2CoT3XIdLrXDpV7QfE9nm86SEkKPp6GZAhEsb0/s
jJwNubk73ltx7y269PFbrAf1sZrZZrr+0Og7z9F1+S4u73vxGzlfhrtBuaJ7OW1L
EIvHIFmUYPXglvgyek8jf9gR1kaOiuLIHa8Sbp56VbsjibB9oarcwU7usiRRuYBi
bA49HkulffB3UxP0lvuV5ZklxGz+HOshmvmMU3+kg7drv7AVYkOO/76PQK6NB5mx
5bqF+38m4QZ4LBsDJacCFnwW7RPycKiABk/ZhmlRSrsXMUrHD8BW7DU3YlSNXR9D
AYaLjuHYHqhPgHZTuJCaqCcoF4H5ZtklhKdCJF64v2kGdY1T48DLXTX5oW+9ONiF
PVMwLJ6CmgEkm9WSVWENBdCzVF2lDnpyYPRzSSH41NV+xI8UfHg1JzQ9BKc3QVfm
DtVZKG5BsGb6/Y2l/yvu6gFTVRRBweA0UmCKTifUryq/E1erRhkMU3r98ZtlPHvz
8NMfCZXtFT6HIrgJZOuyeVkRaeNBULrlVDtT9SkKTUF5r8TjLGFd7b7UhtcYcTtO
NOa7iDaU9XjuE6Kidt0FVyfz5SZdcZdqsuxzTfK7A3qMWM8nyMkzC5qGUZt9T3WS
2jXP/FvDDiBk9YQ1hjdYinaTv1fwtMrOPgW3aHOr7cuc/QdcymB/atFYNdFO9O6I
G5tvk5IVcvVqfbuJJ5aJ2B7ltmhkXt3IsHpL+7edniPtNTBmLqjokj57D6Vx+CfU
LXnHKkaQQsuOMyw/nXzazFgXgreI68mbLl033LJukR4QAFKIqNYTUT0m+pXoK9FB
Oq0T/J5fqsUG/6LnrLQXUxuIlqJ3HSyX8N6u7ObK6ZTWbIRXffRyz5KaGSLkQp7U
InrtVJPWmfOl4oo0mcHJh75w1Cmv+hdIRrneOGV+ETUdbT+CFJc7WO7NwumKdsCn
81yJOBx4BPEnqTUb6aCUzZyTslm2i7GTscaNv6dnriB8UhSPUHHpr2eWKAQHWp8V
xNnxcjWVD7Tq29v6sEj2B3upblhakKUcqr7WRbIV+OCGOPmV/GEBvDHAcQ6/cKvz
wxS6WEXSF5cC7Msvt5q50zIBBvZ/8APwP0dfHN21DOYKGIRjM7jnav6Zqxikhj2X
NCR0cLOnQg2RTOJ7vryqpq88coFtGHEx9dHaQTfwUwL9vZAJ9rWkeGI/KFccV6h2
xXRWqIu+NDVpFJW5KHZFOvl04JIpMWviWFSOHXoi1LLJQupMBstAxNIKcfbGO2sD
98ybNfP2iCXxcSW0tXO1CkmbR9bmwNGBmRNkZudCAGAIudhqSNdE3QVNKrhKKmzI
QDlwIZyH14LoDrkKyFx6CxMXjKatKh3/lQNjs72J0hl3YrkJUFKvaT7NbYyhq8V7
3rsHwbWFU929YsRT+rtxP+4KduTFWuqvaMgLVCVF11RKDAk2+FtiThcZJdTI3s8Q
a7lHB6eCktNkbrY7asjWTvOXwSBwKQsLN/UVICU1mPiqPdhT7OFBuKaZSOL6HENf
uOtfKGrsLLAMlvZc+P8MytE5e+4SJm3l90gSqhktlRnp+TC3cxs+4YRO+GKjsw2U
Ysc5bzurvHz1YdLxQXEyQyfhxjD4dK5nhHE06ciDMg5fnjq5YAcx5HztNafqzsjA
PJYF+YY/eW4PNIut6V8+NiL4VvWVd+dJbarm5VFathegvrBNvJ2++rPkL8mx13XW
9UEUFizKktV7eGGNclE4gDCSv5H0OyXXeeQX+LWZn5WpXxpf+Vwu5P+shintx68B
+oG5bqNQ1C4MxsATi5liqx9qeV0N3EEna4V5wsBQB/lft+IziwfzIAEIE5Uhf4RB
Wo5IhCN4SjaRLC/uqlyD5xH/fTVz1HIXvP2gxZkHTqXoXWj+86Y15tlrXavYmLF+
140p86KgNBDuyO5zGoCJX38Z0PCCVhWY3wjyeW3LyBF++pqRvEeFQ4T5Tmor7Oqb
wN10F0gtTW63WhsvaqRpmert+ECuZGGaC8fQsJJSLU56idw3yjPnU2yQF1Qcl0i6
bYVPRuOG4mxIESto2FPIoc6zmYleUKiIf43QUqZSzCj4yVFqbuzroc2OlovE47rE
9BL3Jj9hD+SfgWm+CZbIbSQs3UFTETV36akQb/Rndbahl2+s9p+KuPnq/rybnGKz
fDx8uW+44DgIL2eGT49OK7Jok0wQnsgfRjZjh9ESM0J3hGRD4qM5W29nVl/01PiN
+6W5dCBO3L6XfHDB6Nh/NGLvne8TmiU9GohUZkNUUHPSnDkh05OqvCccNkFHpLxY
/ML16QSfbBreMldYT9/2enW7RLRbC7jJJ3qDeTvwQNL1qtDPUCsbXdECVUd8oQ3V
ExhTIrhZqGfzrSpzh+6VuMsyqO0wtM5dtZTK2V0v3wtdvLJIHtH8p2jbZKAenHTD
pA7lk/7NOzivK5o0Gertn+B4jA3I5MxNWPtRPqFJwe6lv+X9Wr1CFVH5Z8EsKZxq
3QzHIuqEo6svb7LRQNDLzpTv33Q8lwCqgC99RrFYjIAGv/DbS5DYnefj4Kb3aNGO
ENUoD1XPs7P6VWSwh6mjVllu4zQUGKA70BimMXgSkUDxvtbdgPkN5xFVy9srt09A
4L0ZzuPi0a+G2/cOGZjB9pmGs/mctUAy65wBboI8m5F9feKh6NsI8eu/F16SgdaW
7osjt/BiExOTLq0xoVXGmb68BP0pgqqQswQY2GPxk6l5sRRrGwEONprZordQvDC3
xA4aSXP+61iveHf8vS4VtWGdvrxRYkDjpxMHD65ayKc+c7z5qNqiI44zLP1QDH/i
7kl3JusZLckRLII/s44n/rE0/6qRwcqWhXz3LsG/bb/vJIdORVEoP+JxXTA16f6q
94i90JewLSQyYH62u10fWsSzlVfD/EO7v9px6S9LIkBkL94Ru8+xRT3px2vD7nU6
pNSbAT3HuvolHzEuOsLf98tEl/820B18ZY8/wiJC/TdUjOhJI8B/0f4lQ8jLMf1f
Gmdz6ZN1To68Z7/8HQMVQ/TgDILRrs8eBPm6qg0QcZE0+eMz4TatgieYkU8p0oA3
8VGubal/ktu3DPDe4qUGqthp6etvt4xe/0McNsxyZXOYsyK5jwpy6Q/SEeLJ+PRE
yrXnCwYn3scoHTyjrEN0bI80vGhXGyK2wjEZ+3EUxSMkyZ+McCDkuL4/3UEeD+Kf
AyWgjq2Utmjc2qZ1Pio3CE6tXElCSTT6lKv6weQKrG/Y+GC+8+hkE+SeTpyjdd35
incA+CBuWT3/20yL33Z0SIfiBm7vg0aTdAFCuDZwBO05/T6O8AsenSxMssqwtUFl
ZWMOcUkUPytefB2iHmRpd5FVl2oSwqu8bTw8XHkpbrXTq9PcNQwE4X5UdBL2GDMl
LhZDJTecjoO4uCNZz7V3I1GZYoQLUcPm12j/HEXJV/yDfgNLOYC/xMmzbCKlw3Uu
RFhdCOb5zbMMcSGi60gxnSdLyeRPXXx4oviBgVtKqKA09VskFOqW19qFPFgmgqHp
bs8SoUB/fjFWC9yIuZ4LCgVLdiVRUfCtsd3Jxj7YWhuUDM7GkHByy2dlTOtSWoWW
jYa8ivhQsAJePwnqduFA/SUaT5JIOuE/YYAjnvpfYbFEmOZxPgsy+7EY7UYXRWwO
4ZiG28P2kUuM8bBsybeNW7WgYLb4ONTPKCq8qyUD58s33hyqktAOB1Ot3FA0HIrW
U0H4Ke2uRRRvobTnDdI20awZEvJn0f7GMCXAx9L3PVkFXiwMuCofgrvYft8urLdo
AAs5n5iLlE07aRUTklLZGrhz9Jz72EsK1TSIM7cuxDudUbo3zRXzfJPVYI8JZO8l
IQxM/Uav8dUsew24yXnAmMdK0u23yj/wuy4Kka6TJ3i34Y+f1/Jiku+sjkRqbxsT
vgIkgj6sQsknc0WLysacUwnJb5r1wnvS3D/mo97gDqnztNGoaOeU9K19HwGPL+Je
BN4uTkAyE9QoPx8s24+Mg6S/Suj5UMEfbMoeE1ADrgm7OufqdAMhNb23OKuuXQBn
cDJcQhS8yC0sksoPOEveh2EqZDx6gewDMBm1QKiu7VL6cdmTdDNxg/UGbzmYajB3
YjY2a137gWdKgoCOUhTMC0g+NY/oAeHdRBEBA+X2m2+vWw11rid29Zc3yRXGAaGr
gXW/eMd4aicLIESsD068P6ulRQoNii/2tPRynghWH+qgGewg57Z2IYgkCi0/xan9
tExFqtfM7mibDuVfQOtraPAupJlWPmsdVPhv8VBdLigOehDU+vNkapuhYH3T2SjY
8hJFypm7v6FC4Se2sCZ/PNUFdF/f2aBNPIS8VHmi5EI91iwzSxGmbP6xaA08qMnV
ddc+UuDZrLgsmjmJkW36sXqXwPWXoxYBZQcvZMkGuUgMVE7vTnRUGl5XxgM72ha4
zTlj/xZAujsrE6Kt1Ii1iOm4En31VeHtuL7ekOuEKofY1OvNmzEcfruiSD88+kN/
Ev45EAbN255E6aQF/D7FwHN6P5VrtWc7xkm3EnN4/ko72LYiyxmWSgx2yv/OyWeJ
EAdXdGWNlMzY4Ttdti2VvazVNNyLHsHkFllEtnhmLJbvqoDV+4gTVeOmeyuWS6du
ZmDSnC9y52ZytToOb3ffeJ9ws0RdRbUnli5Vrq9lOeqIpxAajv9Bo/uhgaEiRgVH
4EsElq9uOwvaB02ge7JHG7OCkgQNp6G6W7aqAn/gjGejdSWVO4Vl2t9HTUi95UpK
UK+r6w5O6YFAjjs28IvsKeLy8A4sbBQl2BRDaBgnYqyjnIM2j7F7RthqM+3/6Zi6
j3iPgXijQ+h++Mj3b6IOFKS1fePGqZDrG+QNfxf18k3fppjkSPkYPKf3yTTOZ3xB
sCco9MtjxUImzBJ88ztNwaM1u+iH+VSuy4qvL8DdR2xcXj0xd4vsZzQOBfo4wJ65
uRynvWVn1CVhT0r/OEIljJDoaLIkozl9bHmfZNY9oaJ3BHR1rIW+Q0YnW+adg7NI
9VeC24DyfPzYQRm42s+iOFYeVnLMaTw9jc8eDJ72Y5tGMhPldfniK//i4U7QKu31
Z3ZZmn26ATO5ibi3pXdb6BRKFr5sbg36r+6REvI5rQ4lKexRGzlvOurbDEJFy242
bSHCrsvBS2p2W7NEMLSjd7Y14OmnkopCl7aZsdlOr+wZ/hWGPBcfGWDu+Hiy2e17
1ZGfS3ei8n/OkqaHxakvJ3Ng2Mg28XcYS/fJ4WG5fgBp1zwR04+8vxUUvbIag0EQ
zxX3N7VVv/gfoFzeKNobzGTvqdvRDzbJBv9Bzd/ElxsImmHAiP5Mq/T3d8dc8jh/
KKzYLCgHqDtiTNfguReY4nOCUBHr1pfwgABfBMOv4aM/es6rDF2Uqljw0NO58GyY
UtJNpAB3VRj5NNri96+d1pIEgEgTAL5SzQ3RpdcXlQ16wMzAPNlKY7c92IBiYe6i
5lCjsZiXf2aJHHNEqmV0L1QMr0vzm4cjhHxeqL9dlQYbWuDCBQhgndz0J9zSSo6X
NwJBIJEPyIwfob+FnSIfgatsLJLGefuSC+7fUv2aGejZ6oAkizNhUtBZ3SQF23J8
13qkhcaGbrto5lh4qrHTOfoehy3KbVSligwXGXZEab9Npu/tCdLKVhthtahD8HLI
zPi7bajVaqSZTm27wu5LNVKmGI9ac9KgRoLPpYWhsCbmf1KCpa0fWs+k1qX5NvO7
jP8HLb75d+oRcgkoOgu1AcUF3NhxAkALR/MUUOx1LgUPOR0LlLOTLGwzQXUb+sA1
yBW7CDAY6UIJTQ4ksNAUgfc+fMkScWEDnsmDpPywvL5WqO3iyD26xTHuZ1KF8v1p
LTvbxCGy34JpkGXef9Q3GqFbRtmOcpUFhMas3ETh3C8CWkjRhfFLRmiSKLhgS4V2
EnZZeGyCd4/paDX6T4bBJGYvY0ae6NZuuETI297p33FODU5UFL6+87HP3FQMY/No
HVLgRF57bNnLdmVurSgNz/8eF6CTY0cDoeLJM4om+84FhFFoCl0ciq34oFcMXAwT
WkjSTdeGqY52aGg4QyZFhWTRLg2J29YGIQtwCfMLZaP/Uf5yntVsP7e2VpqyXf1G
DU3jGNHIlOC5SK+CiFn9hqYSCvqxGm4nzaymezeDOdE1fBRM5+Nyq3VPawOC6a6g
lfgLC4QtT5rcRYTi5tJ1/hsfppO/fTEr734SRughZ+YXG40jSVByaS8rg8hniKv1
N0uo1VldtQAGcW22ozBgYTKh36iXNBrytvTSPjL++UFf6QsOQBNKMKBAzQuVeptq
f+lBjOMlHdav/7Iw5WKEoXorNPXcRKMuOe6Z8Uxw1Ecx98u3dw2gudlq1s0WOHsF
WQ8pZUHQNNV+s4zeStXpGIYeq8n7j8U/uElrmaujjBpuJNV2JFRSdSxgZfVsl5Vu
slwj+Y04x1dCggI4FkgiEUxqwIQfpC9qEpKZkmxSwx5lYgk0KQJKwGH3bcaAgYuU
HM7Rj6uCX9KKcQmXajKZoNuTeMNtYEfIE9rySqxpN4bMhlNzZfAk72DOByP+2WQG
WKTTInOictO7YnBKJryxsjswWx46haxIEKsbgTFQ/KTaVWB+//rD47OTlnEINle+
Y5HhQOENgfIY41I5aq6Y12ILBw6xN1wAWZ/PfkRAePJGnAQm1OTrF19b43d6uX0w
EbjEg5m/vGKiNEcYzJZUMw52Cm30DBe1ngyLbwjog1WSCgZiPTVQQ9EO5NlkooUP
KT8GkQ8IsTNo6vpng6CC5fTiQhC5J1stPFm8hyWKFACcMrlx+sdX3nwRfUA+yG5q
BUechAbMCMlEN2kwhjhaCujU4eGxhG4ztDuQdLXB4te/sOMZEG+RcurCw35Q+4dQ
tu6VRXn0ijPX3OR54qiRa4XXGNLs548Fsoc4jXTjVF/GhAjuAJs8fkdP+Ml4YSK1
5zJTz1iw66VnT30pflElFnCgqH7Yro85PhQbFeS6MIzL5qsp3zjjNnE/waz/3PxW
kNdrSAMywnR+kSZRWgp6G/wRIXiJUNDofSkAe6EL88Yt2/V5E4RXT2Ia2LymQ+C1
hVbqjR6VCUsv7qht2wl+pp37Ycqk69DghL0vq8AkffZtY8ERX1UfFrBKdBSglDKH
Fqhd6cFiBIL/1AdB0ZJ6Shwd9GFojziaG0u/E8+L/BGB3etQFvk5hyVZTJFpPhf6
Ij30uf0ITBbK+JcZHgdsvrfqd+tVecu/riBd0Uw3oyrDSceRJC7QF6WgcUAXDiu8
t8jXu3L2JfSLsuDvxj0N6TJhfWgPespo0WI2lhaR+Z8zI+rD9vWG6npSMfv5sgYy
vxxu3Ou67ppbwshza+y2y0pgOX0e9Y2nrpIgPNXkhM27e+pBxItTRtHrqColkFiq
9VW1qqai9ZIjnPOxbu/sZMAv9EDM57RmxAIOlGMMoNSa7clYoCyoujj5waj/aPPL
Y7xnWs+rrBXIHxR0i39d71Xn4ng9TESgLLVIRdJJVUhw3VzueJFCdGIIPI1oFPTV
/bs6qd9KINklSlSgvIQErnXlu7W+TYb7n3ZTTuCYOjMvMlTfxLQX6RFkiypbMV7R
KHdZpzvrPOalU64QjKxLJ1MPLDUsGKLVAj9MQdo80jS/34xi79h7al9dNqleQZdg
Zfu8IWRL2utlD86fSicu8mPQI/TVa2d8wF+w9r3fELpe3Yq8V2WQwXOmw6xEmKFV
gN8rXevUAs7CbhC0fyFdsuiPrRs15iVENByKCAEuHgnwHGMk6+LDE/LvPz5xZBzg
QMwxlgRz+jBvjDKjVTlUyqvAtkCo4o0vTPg90NoAmOVwM7DP5iAlW6gMngNikjz2
jnEbbhVIpvt9AjrQy8V+6bUE+VgGmZ7vPCU/ONzVgorNPZnw1aK+rCrnsQ/PBRMG
qqSocf04JOeDFGi9teVJs+QUqX9zGlRkWHC1EUGmnEHIhDq5FeHbMwdQoaYyMJfo
kl3dALZ8k3jdgPKLYGdEckx/lwRhH81NBnJbIhQZv7RFI293DHScbsVlXeDoy6+M
DbzyLtYgnwLKKOLKkGuB/IhbXKDmPCE1ANavB2LO4LENc8GAMnbxYSglHZ2fnj0a
sjlmk57ftHgCN4YSFpoXX1LlrqMuNLxc2pt25vO5UUSf5UGevLO8D73PqfgoVryF
VO9a4AS21F+6DNR5X1qN1myfELeXcsW8d/BeBpQgtWg6mLHufFU57WL6IWVyUyGt
Kw3OKl553e//fPv4RwCDPRSppx4kkBF3lsnlISh0Sx+BuxyWaVqdLKz2AYkI0rGC
IyspFf6yrS7Tkx40QzA0iZL7U7iVIcpxMf7a7pyAxgy9JnLxmqLtsW8eqHLzb5ky
q6WGRYVkmJLLJYyfQ9sVQUVTaYb0eeo3aKe8fdKeg1o6g/BmHo33T1iftNygWnuT
aFKOLkVbt8HfC1cqEUfW+r2AsqW3OlIj7fBtuS+W83JOHv9uuuAW+/sAWVUoPX9M
zznFNJhLVWlxJfsYXzaHK9bOWyUsmPxOSfKnnMcdwPzXWqzdvb6GdZf42Jrjyo1Q
Bi0pBaNJS6YS6IMhsaN5bJrSUqmFoVN1PdyR5NoQVlwGVGEHfQYBRcw0ZE+OLAAw
LiW2/UriULXdtGjlLTbYBbpu1Ucyc6ED7MySH2FhJtNx2UZ5xXG3fX/st6uD+JPk
A0bGs0/AnRJ2mCOwiU7yceiNE85+6ND9g2y6yVwuYffLdBDH58XASSg9rrgtU8QJ
YkJtmbgIRQh/i93waeYVXF2smt/kXcu+oeRNZT57eua9dvRHCo94SH2KJCJe4JuE
53tH87MWkhDX6FV37RRiExP/CTyyKeKlT7kUEyJnxxIJdReOULMq0PDbV67SnVNr
UPZvC910gpg/Q4sAh2lyZZuJVYBHKCzCxg8bh/TB9PX4dNjrO3I4qu6RwlcRncb4
Ei2XI/Sou7P7Vo73haZxNCkgG91vdh3Zk9n7e+8iFRFk7n1muBSkFq8Td2BWygJh
q6ijiXEr7TpjeKfcxq/ht93H3g7jdoFOS+maAvGm/gyUSLWSft+TTl85IdwLdZXS
9O2AIrYi6Yjmx6deQyhg6AEpr0enKiYUiMGA09fpdVB4e/OG3SUwivRh3JmaY2sO
Z0n/IqhuEtMH9p9g9FQo4WoYqbdC3pPdjgLB8PcFIRwBZr6h+kl7fVjZ3KqFkbcb
9goJIsf0Plb5Iq4abz5Cg3rEX0gVlUXzOeu3Zjguuug93re9Aqi+ixR7Awr0b6YN
0J1AteospbQr/3wGowTY6oeG2R3UhfkCQwN/Sc6fyH0tb/Q0j7oGe1v828tEQda3
NgqYjwgLDifBxcZKsohnD/aOv1wxwr74qY/6F6ZRBEUz6EAPwa4sRcF3P5/vxRYy
/ljA+dDJYUlmxbnoxQG+Si2qrgyiCXRE17DOfYUvx5lCLFvWWpXWeFtwUTYw8rV9
NPIV/P1Hvj1ynDN8lOLL0zVlAn2q39HpsVGCmiikoSMY3K56/6DIHPgbBVjznCa4
nedRjl8vqIIWvgYPGGbi8SieaKvXdlgPw5FnCo3hSvT5UeH2SVPQJ/WxbFTcdUHN
DlHjlRqG502U7P7hCULyl9dXfli+pxy4nO8ad20Vn2s0wJx1aDPqo9QXKY28lCyi
XtuYvbfVyTfuQKVGTL3Vj++iONrYn+N0QVPko+6zhAre9AO6zUkWSK34FsU6dx5Y
yEgNEqBsleNSjq1q0bGIWkrXcL7ox4Q4HmLGoduNDLJbej3sSNyB0HKPI5adzGUP
3ITyA3a7Hp3SrBvltRQGFh+kctsCmtM2XI1hGolIReOr/5YHeCVELrLeAWC7uTns
grwSiHR6Ey0mYjOyogj5iewK0W8t5K4t6CVIlOMg+ktVXjPy+zzrEGW9G+/pQ1dM
suzA0VTQMpuAoZYff+gv1vWSVrpZ8TCYd7MnQ99WCxQs0Z80n903y2/gmnoV8/eS
zj4QKMXFp/TEiwPJ/UxD/3d3zit/5mbgYFxxlOY6uojL03HWVTYl1fpJi/PK+EE7
r74HeIyuJnflfj9mYKD17lbwacHujpd/er1OxGKYSEKw0BHVS+XDJceqtMYG3wjW
cAsy09I5djtILMKDANoU4tY4l7fblU+QjODIA5ebJ9lYysSbBMDtKs/lOBT7+CYd
JDRvaIbmznTDNSYObcd7wwfIO/8EpVh4LITOEbeY13GFnwg3GcH4hpdXsKTVicKa
Nj0nB7IHhRegiGYky6gKOefJlqtFAKWWcf6scM4lqRfHQW9gJcHdxHkgCeCJHd8S
V5K2ZtzSTIOq3qzrQlv1Rqsxyi9/gcbXUuliQA6wip9X+WWgixWZ+a9Sws/T0GMi
tfT74lEOUTHcpkRMJ6GXuShcuILHXukAdKJJdQY1EZg8gVB8vRO1WVS82dJY61DQ
CDh/MvB4ohEBIMqhlNDiveZmHAzx27Xqj81f+9NMi14doKRUkltdF8vn+o8dEdjt
uQMR9QGbGZ+ztbKFXI+24pH1lA62MhKugolITwH2osuAh1K1FlZZcWZihbXHDeUi
WMolywvq4SAfgfXDCwmcNEPM28E0l7PlwXnhbIAjfgn7HVOS0ZwG5yno57qN0xlZ
87uCW/wtOzRceTN04P3KcphwuywYrzNTTvRgHN7FrPTtC9njTxl5CvrteHOu9fDv
pTaDdanbTELkkm+uL0ip6oC63QytiMmHcl2vrtVAFYA+AOELlw6xHc+w3jQM5wLI
gkUen69asAkeMB5Rf49bm+8rurytRDGRd6QvYP9PfRqGVeKeMa8H8M4oqwT6yot4
iBVHVMJW2crL4DSqKfB99he/Z26eyCNGhrlGmi/AkCevz3oL1kxc7DrXXjw5p8WP
DYTgnd3a8xuEtiuo2uoC4NKzzlGJUf83ktzauT4qN4OW1/yNl1Mbg78VTbThfYnE
bSU8ijV0eJpRmWhvatu3Rj3HjelWal/BeLt9l0P9aWNgnk15I6ExrgZlzFamPNYO
2NIx9qb6I7CeNKsfX1QmrxOD15ztyjT1S6Rk1toQ4w6LDnfRFjtvv1QDT14jN7GC
4kFYCcDaROa1tPLRMgDYg3+x80ZPDqGh9J6iYmWIuaUnrgVRvf35tiSMVMHBLfAW
eFfdxMildlvE3C97hqttRo8c0owgsM5XwhTj1xZkISeUGCBIQNG4Y/RLJxVk5iqa
3VJB6ePnEbgAh2mUASGBiTIbwtvu/U0cHBNqxAbCFwcD0deVqDd3KvDCHutXTVdP
HuLgIUlkJxhVug0Qt+5vEa6VACfwq6AL0IaWfWUL10jcJlj19m08O/xt0NrUWi0F
Ib3bDY4NaGCGRGjZGIO/1VWNIMBF+B4xTfAMmZWEqIWgI+emh67JKVOymN3vrp8h
vvBqXhuNHkf/zcYHrGAdUc7T3YQICmKq9BtQ70dUvL0533Y96hGnhtKoWIBTi941
0t/3DQH8/A0RuidFFP1vEGKoZXsjvXnO9KL/el/R/cGSrdgKNMddd1u940mQzrsh
qNz2M+o4b2bBTFyhYwTORxa4Si4Rc1s4k6lTJnx3A8emxnvy3ogRNuZSgtT34AIB
b4jd3f+/irMoJFmrHzlMFYsVhiOc6474RLRgrIQu1sMw3zSPDlq4vvJy6ZVog3FV
FD5jPskaSlnGpZqdQnfVQW53Iy3MITa2FENR2rF74Qt9+JoX0AgrTk62BaGT6O2/
sZwuQGVgY8vnBjDd5qFug/WuZtz4XzdRwSJMYV8lYbAEVrOIwGyShOKoY++qNKNe
ptUip0jgceZaixqoINb1m9iEMhm7AGdUMCfnnYCk1bjtrDFvhUnuingXjzvQTxNg
Ix754gkRzKJ+X9FAKahxJWQ+I1BgPX3fK2DGqaSE7X59K1HGz5ksG3FoeM3jhwgq
2UbHpBlTtFXNgyi07lFKS3K4DfB5ful1fA998DsWmm4/MZHfEg7gwRpfIi9YTVke
lR9ZVmVzuIiCdiWUY05BViTZ39v1YzjF0XJqJBASpvFw8Qj1VV5oZnUXrac/tyD6
MwTK1b6G3y/NSeUrbVR+Q54aeyK5Ar7yrAW4365QhUFEc29vUP6OKwOX35lNU1eA
z8Fb4cVT0/L7GL8X5Kua522wJLeUsy0furKSCmvQe4m1MFwjnBGCJYVVOw0k8Kkn
cYZP5DQ982RH7kvIMioFqIoEEB5g2Np6fEUeTx3a6LEc24Ajjkr9PcDfG0KLOfRd
BZMmah3RL71VrIiclR7Ts2o9Iu8UUxR/dIcmLnqDOmdB7tx+UDgr8QMyEf7DxTzy
17YdljLLk3WfPjU58Yc3AjdvkAOk6gSn1+enFpaOiTXcOxvLgKw4wbXG2IvnpBda
WPMH9GpwZ/H3SW5vHoWrVN4EoE9agvZIMfajJNKIWrDF6DR8nNE6/nSWvo1UgBgl
YTk3TNJBPIWMvOSHusyxiJNuw7H9lYXJEh6RWxm93n8TdTc+Hk2jcdu0W4P3ROvS
t2Juk5f4Mv7lsGt3iORtTkr4VGhTBMACc0HWE7TW/hraeRfprptVJT3gsEEzO0mx
5kg089fV0TmvM2uaVcGEE1rEr3sgcKI97D1V+pvxMMzn3F9g09/Dh8UG6T9RVfIU
OnmoqXPaeff/gipxEbYjSRBGl6FlEcFtdDt6Ea9zHMuGbOIS7HdXxanorqFK/9IB
Z2Ut51NnuuDOntvLgHtd48f2azpOR3qlA/i+DXa/IDq9JbSHda6Ia0rtlPUf6xTy
jm0OtlFnVyQ7wB2oSnrj4Tn+dkHSbVn2amHSksxAniM3eKSk5lgxTO2MWOcfChxV
tGDEyDTzp2Kpn57vxfn1NS9MaELw6cArL+NuMao+SamRMamEzTahKh578OINEJOs
o6yuiteUngLyjygHlcokdZWCeI5HFoLV45SiHBz8WJTvLLS+nUop+eBcjGWpsffN
9XQnG+J5qneD735miXaYlqJQAyUbm7CXNFsPrE2PfFQo0UPtWEOAOkbUOyjfQu//
oKcr9/MjZOmaOCfU7GQEu31KQsPhYJ6cJY7eUyTOOTmDPSwfFdZyIGnMsyGINPBU
irTgCdbierBz884SL43qbRoIf4JCRZQq3tNUvZMi+LCtChUP9QCPYHSUT53ja4Ai
91txG2Td1xnS2/k84UHRu0uUSibNApKrlj8qLgFrghm/1P6s0MFB9p58B70g9BGP
uWEJHgCJ44mtkOWMQHBO2rRpI9K/kcAxs/3PqNywQ3YkhwCO8++Lvsn9/NFuc59C
fXD7gJnK/3UzlHysSCtC0d/OTgcdvGfkoXVia15JT85Zrdy/06dmt42fun8GGpLq
FEQ+9116Mr7ZZt/MB4N+zOGesv7fb+nG4Sd4gL8xptE19DakzK95jMqxaASPZ5l6
I2QBp1bTXfAJPelCfiNKv/Qoi4P9P0KXBzKBWhb5G213UxV5tooRDX0Z/tRM314D
NuQ0+ZJOELmexnaJGXJO2jM2lZqo2bqTUHzMFcdWbHSDODFgSJAAWezJJKUm6GAw
Lj0pgyoi0AqcB7PkoUyhfkNxfiMTp0yBYGGXA8Srz23hIGPjBcaC3qRe4lIdrpHw
qsoAAi+ZnK+vWLw15mvDEddUFL4ROny+5GQDMw6USfg1vhA+0ABpFFxsWAQc5QhD
EuNyyMKV/YfD9e/lKJxj60bBHOKdrlC/2CDsCCyGg1GSjQqewYT+MB4Uc+U39lFM
tEZvdl7iZshf/9i2ZyeRdSjOgWpr6z70/LXfXn04I+A1jTab2kTVsHIbQhcDym+d
uMWpldZiHhRemUxyb1O5b5WxLvwMdbpIVNHZs2Qbx0YmErDH8wYSHrvhRNgQq99s
rw9vQWPrgniJwrR25hS64VWHpKNE5R42Jv+MsqC96SHK2EOiQVTQK4YdQ1q8j8Eb
knSTXRwwoxyGHFRVjpqlEp6N/x4GAgEcbF1hhrE03d/re/CCE5F5Ft/ht4Yhh1Ex
NEheF003SBc0rSzon/mIJGx0hb1/RM6LDkYRSWDHV2FsAaVyQ0oWavuuj4P5t7+6
HVW/Z3AiE+UFE38Jqyz+ZigRnmLH+Esmse7ej8bKkRICXRfogJJTSTjCi9PpiLv7
pempquGrR6kowLVyyhAMFU1c0eqPJehSkywfhwjM+uRdaw1qTRweDRdW1RhkkNU6
wSNBUMXX373ofDLL+YE2oWbGzGG7POn5d041mREEnj/j5yluGrbHEwG6IOxODCP3
NSvGsEEN+kamnq1by4CbZuvDXOSWg/iEGkEa9/hnudbHEhkX+Fc2wl0mxnb7IRjk
myapteHKP32VeO7EZAIZoH083kvIJgmIduE50sH41CUbqRG8QrwXl44/mCEBeSWC
pOYVY6GYBFb+qy7GL5ccKq5Fj9fBVr/3HCSCWPmI93L3LngiKfbcv3VgyDaV7P2+
QdoKDq4rL3jT2qU3DjIhjGTdX0NH7YQvvD1P/VK5s1u1tjXXb/n1Kvuy3P5xUaEv
11/L7gJBDvVBtddu3tgoA6UqS55emVOQOfXW4Dob7J7nWJ0iZ/UcqxUzMAOy4Nws
7yex2h9XdcWbcv056QrgxHaBo8UbuT6hkuow1mZO3lIkUX0bSoLGuiPUB4ZMguFr
BuXTlKoItqdjDpy0qy7OC/YdoPuBBvTGOhf2tPaztGvP3U0nNEDyGR+G2QxPq8SG
cJwzFSahwW2kfH2c3jHy+ueCbtdtw8q4R1Um8WEEGBgHwEquGxpiUw2G3AxnWvQN
yugMrYqSt2AELEis0qOqAFgkrYL2xFvnBfTSN8u7HWS6OP8KOYUwxXuSzKEt2uyg
SBKwsZZG+/4simsjTgm3E/qtRXpd3PuF6WXzu1Oy6EN8u2ojF46qO8F2mX+8Yp0g
qJiJ1rNGv6jYVGAr8UWG1oRDQdujA7WPowSNBwGI5r8UeHjcNqkpfJ+1jh1Mf+Ku
tQnc+NACB2OBAwJkDNpyo2l36rvd6pnJNUeWFMIwR7u+RUci20KqRdtibFl7ixIf
XxSVrZryMkNQ51r/kLLLrnul1DTo5mxl2exRTukwEaHZBvxzezVjlpPIJ8bcPNoY
7FI560Z0CIxH7JAXlhtG0BCwWw0CB6xeRf82Ey3Df7d+L7lLBAF1BLSTummGnUkX
mSUue5HBlckclxzESy2fKiDe2524Wvapwj3uJn/noz8fDD3S+o8oQAsOANxC13Ir
5+Hn4iuB2z0wrEXp96mG7eORL5a1cahj1yItHks8wb+KUCfNmU2qrj3VdXsDMWAA
DZPeeM31T/gT8RN1kP9O6fei6mn1bDd2aq2BG43pv4kKjVKOX+kx0PqwkxECrdes
Ms+oCh/Ny49s+kW8ualBcvrHRSLbc67Mb8tXwg2+L39iBqmW70HBslEuV/XikcBU
PAbrvpisLwzKTQa+iW1ang+YiIdWwzhkworHeZYlOOPlqvvDdMjdtdIyWQZJCEYc
SDKnJGkvDou32h+7h96kDkJ53NnZVE12Bp3PEujbB2er5Dbd4LvHVBnak/SOsD5f
4PgeObfAI66lCx0j+4amQaD3cS5vIjnpmzVW+EzMRGnRe6Q/iS1dGeBKsF28cTHO
+wbACShLPgdHJUlFyUvFgUAX3m/lEzGoS/Wh4qBKM7xjE3f08FEiV9Xt8ulQr/+7
cU5yIBSOUgoLln32Z+hJGtASkbo3WYo4j4Z9MskeV2cPc+pSncgKp4GFvGiz3lS6
ruzQGvgiC8j6rLCEKnPny9EyBYz4rY34T5Rv3nyu8SekAe17GIozsuK23whHtuJA
NXQoM5yg/5BZrztzdBg2NNn4d79oVF4ptijvP0VsksPVGJpyI7GNU7sqal8Qf+Gk
XFXZOxSprMhrp4H214ckpvoRzgMoCtsPgkWQnl9uX3b/0BbD1zrFdHdGaMUKN0Qh
b/An0DJ4o7EerEuTko0z8oy1jnKx/smT/DcLEfBgpt+HIgnMMLf6WxNbMOC7ulqV
eElMaEC0sph62G/a2JUlUjANXLwJMt5ZA/hvJXN0eevXyNSbhzDi7L5mA5kGJk12
68Wu110p4sfFoLLedql93d9nLJLX7LV02nI18nOUUpf8PAORyDWh3hK45mDUBfh9
uvCyZxLCHERVXsm/NyXUDDvUiGYM2OIuBoOcNkmUi4HVelXVih6J5ZRXeHDNaigK
I5xLhPnCWAKMiJm5betdxN5Wb4SQBMYlPT9Ot5CckTOG1OppZV0jgWoz+bxBBZCP
2YgdN2tMsY003Ml0SClXOrL9DhVMC3JZJdRK5PDzVfHiZZzA3QHvSz2g/E8mZqj6
w1jqRYAQY3ZS3uEFIijUUUdp7zKZBOXDkgi0dvED3eWbxXSb24ds10V7ZOb5zW0l
2+O+YeENyykfvRXje3MXEPZyBePAfqd0bYdQx1rQAG5SwFZggL2PA5p4WglgWt0m
obMOyW5nf7i23ZRDda3pvj2AcKLYbj0hBWEPaIT7FVXPfvo5fxNZflNz90VXjYDC
btxgesearVSb2UlAeTs4xcy0j6AXxAKXOxObBe/ckALGpXXatc0IvEW4rYp6yBLr
bAHTTmLY4k6gyGqrRulGSeYs+Iv+mmQdUBu/fsT1NXLsORe0nPbfzBiOgE1G76Q0
qmAoxWeshV5pPHc9OywS83RLOR6EO62/WMcPulhrVpel5dxbTy5dDHaTW/H/t4Kl
kTbZ+jNWcokOZVCbrktpmtiG/CoazhGiLFgldpqs6Yj4JG4HcZZDLnuTiCx9Mk6n
l3F2cZyQw2Qlz6kkwk/i5I8v0xqujijrjbXLrSMOtIXcNb+6et+LHGbAP5wt5qNr
uEiCPr9k8jRLQL4FFA8TMKfHvnC1pO+8yeS3D0vH+S5lQvOMQtLzHTA4jXr591TM
lbPgD6UhjxowMnWMIZAxIXcdXJEmXzgL0N79q5ZjluqasVDFqz//oC0ZSL9MRGL8
9dPifZ4yMXrAmZW2i3wv3znF5qM+onllsD2aXwOZZJCNJUz1a0HcKao7VdBQN7ia
cpliH1/9fCv+7rgLPtydOSDuRuhrquY23M4YJ6lxk2rRA8Gdl3OUd8jK92Nhnx0J
qpCR2Y6sCW1h22xeRCgQ5N5Q0ozGVnhSSLig7zx7fVKsZulpSeSt1q3wb/fifdI1
fWPlDX2YLuXa7/G5NHrM5GVBvN1lq49aubY7Ul4KNddtvGIwdnpYgrIEzXe6soTZ
0edyB6j6jAW5HpR9oFYBFiZC/xG1kQdFxrjOAiay20MBR0ZOkbfdpyD2X5l9qmB5
PP5V5n3Us5MmEglKB3pl2mBy9RLSYIhoY2vMSxorBCt8GlvMCOvQP/UyoUvue8in
1VthlRhH0lcsdqvVPG6anOKzBDxEg6gOye+Xvn3/UzaKfbZnZ/Sffx5ANGBw+ibQ
N2EYi2SiRLKS6shAqnVyzKcUjPg/UhhcgzX2OnmGuksRkZGfYsOxfOWVw9aV6S/B
st86d9oXCvXj3jo/z3c4ongo+yugPhetMIrwvhc3WKW+oXw8GAjrqx7xc42m1xzT
oQILrCsalVsnJYTPisVKGmeuBIWxHNwquEs34hoTEseIGAq7xXuUtBany4vJsgsh
zKJfIqUcGvSSKf0d4+tmK+Uc143gxlUPTv4A4feIORICh1AiY5F1DLAiqDxUoerH
grCkNREBbJccBKyG3zx+Om8fJ8ANmE3owM1m27oHLPMr2KsRE9RomUDpENNA4PsR
SbPDiWjjG2hzi4mCq++vk9ohj3NHJnQ6wrTH0onOl35LBAXHcNO+2/3BBLOyueVg
QW4lxbgf7s+swHOVIt+nwUtH+j3EKQIF3lo4FwMifScSBt6UCvHhy2FTVTI11+h1
gSXRBPYPXAduabT5YssEiAg9ekCotHvyL3NpVRrQfV471lEMtsBDcOuXZ7SdldjO
3H1FPPFtnlFGJtNkepnci3paNjXtRCNThnuEzKXmXEmmOCvyVvtYZSAyjqzu/nWP
tKd2HtZYQexT2t772z2H/VWy1eaFQ44UikaLMWm8X35lvJXwK+/AeGN/ZaAgYshQ
99W2AgqbD2cr39JejvNQpwvu3YaayYjQ4HAZDIwbgu9zTjgIFDGAZRtOTSGGvjV4
0hSI805WL4CUkmIfK0yOiPelG/RWjGav6yM7hOMnpLvIKDlO1m+zg4Ik/xx9raOI
5VCVPBAHoLf4I+MQQmJa/uTKXOq3cr3LZKucYzEODpz1rr5atOdv7rEf44uTx+sn
s5SCGGmt9pzW/UlTIMqsBmWBOQ58AvfpdB//Qn4g0DL8A7y7uIuIxRzfkXP/MQu2
X+HXri7sIjJeDImiEVgvBzMBGxZSX6KS+aMjKBBdqC1vihhHd0PFk10jxDjNa3Cf
UshmQV2b6BNNSFph5SjCgn6Dtcy98bCrk7uLSPvACDI2Y7hwRoivrzwQr7nW1cJA
dTrgwx4mv5VLkBco2hvTnjzwfks4UbsVgxWbW8HEqlI/DMf5ygE+GnPYsOcHKPuO
IF9U5XkODIIBhotVvTnUs/gy6xAW4aOJrqnmIw6C2EmKxK5mO4rHXM9ayfS4lqw2
EutoXzKxuV6Oc1xL3Rg4j3WXLn8X6ki72c10qowb8f0LemwGzOqao7KhQsY3eXq3
bI2QJoS8wSYdUeFbN+zZY983oBSETpFoCUhQmmY6ZsHGVrnMAEKQYBvU/CwyazuX
Qc/mc88uJGzLa8TQN2N1GYpn98MQVgiUPLMFcrBtgIHt7lKmBqSDjmWXGrqFyTW7
2t2CmB/brLUxMmpVkSTD77zygoipxBTmIXcYYhPU+U0I1NuB0IPzbaM1dG6Buc96
30Fq9tczthz4hmj+FvcAMP9Uw+Qd1D+oJ/5NRJgwACKEdisB4mNHnJpl3Es2myCH
tptXeOwKUOcWKoFIGF8hZauXdn6UCbzzuK9qgVVtsNg23m3BbWwKrqB6URborXAs
Jf91hEFqrdjDTzd1ROiC4nngez2teSgb6ZfV84yWDdjP/AZkANR73EmWEH+t4Vos
+R6hSGlDfQcqmSNGU5WXlYjgBjk3qNHwN6yvH3orJSzy4SLMbUJFSHKd3B6RijUS
8u3uNzOmMsgpWJYHKMXaGhwAxexj6xWTuf/76sQqQKOgjwA95HocpGIhAjiwQq/2
oxx8PPKkJKoKZNLHtYqR62hKVBrk5+YTpY112oLXyLSVTAp6Xtqjwf0eYbpr6ThO
59HFyC6Nr/vIV0SDbTUGXRJywTP+2Yzjs1E9xu3u1hJ00SVIqXpVxCxE/wnwbPep
xl26hdI3Qlf40rgKQaRPLvHHSoj2Q8swl9aSN6yQTZYXVHu429kNZ5LVoeslQnU3
WxToOlhZSQLGj9D86ZhBdVfT6Qmf78VT5JG2NuURj6qX9VlH5VJMPAkU99nAHrtL
k64lCzBS0F7n1kbBUYoUC6F/3SarNx+HV07iwku3wWfYPJPfgsrSuxCBSEGUZMtL
gZpcIgEjdMimUNPauK2yaaF9xdCY7YAmTQ1W7qK58avWn8jMw8zBhlyr1gpC2dQS
WU6pC3wjM4zy/wNU6RpCRUUNPSMas/f3mr4hM1Uua48n3ptGhibfoXmmHUZaUyvQ
qLFJjxs06wYEMKtgo1Flbd5MnlKzNvg2/6MuMWAxc1qttOLUHGAONqkgOP/3lN5v
Pos6HMGicR/PMLKbneYG954mVWnwn83Q2JiNqYvi0PghRsRImMCEhsFnRCvVjY7w
RITk08ePnKWHjhjr6JQyo4ghSrKL3w71b3m9V0OwrDd1REd63Dk71yuePOUESISN
Io9CPZiINEuluIKRnGAyB+VOGBYiPMpHpM2j7Kss8ZME83Ft0E/RVs4h3Ojk1Iu+
Z16Cp37+NzkkR4LWb4M/dBV0ZSHhQaPTvHeN1o8YTeA22U12B9sCzR3e3pOtroiR
o0oYib5ujia4HYH1TMKmSQXkolPLUzlbDrrPEWN/sBq1erWP/h5KoSg8k0l3/VRN
MTp5zt+ehAj3GdFzUtpq36pWYmiga/05+VyhSMCqyJtWUA9DZ2lwtgjgvv/1C8b0
EZpTFWniFGpPuROzPiTo3L9JsCtUhr/CbeLDP+jJEFZclfoyoSSZ4iyfBaJfsOzI
kbkIzRD2DofhIlxpW+aTAd0fUQnaPDhI9R/DmsabRABW2a/1Q4xLfi6UwyJY2L1N
tY7t4csZBi1Wp22cpiuIxFC67XBJu78OcjwoaDexJUBVxjsKz0n3Ib1UsWlPZ5Zy
nLSzk6/TiDBAWbNz3l9QmRIsdj9cdwslcp5egEOJQh00GqEul7t8w9FayXyJYnBg
1zunIPVEpNYhnoT+9KDoPcZVHAUtyRMPLlUfSX9V9rcy9oY+5Dx7pA1EuQ9Gu7t1
RUl4lye2Ikwo1/GEXm+assem5XFDVbUfj0B0RaXy9SeRklInIl1oMu7KpCrsLi1R
R9OQg2Y7qiimOXegz7jM8GiB0qS7pSGAJrQXhqPZ0HIR0dlxz12S0MSzmGIXxUW7
0TelZzrJ+HLVMCFh5KzUSOxBBZPSP24qqKOV4iC8TwrnrMdK8NWR21YhV94DGNZQ
1eBQKH41qT4gFyFaAMCaI96gG1e8JKvuFa9kdXJPfkoQd2bwY8rxPSDYDEEEb2Z2
zI3AAJtqBCCn+h4Krf8Sv3btBcTiFO3/ELssHASA5JaXzZp2q39ijdb1/PO4WUs8
ABLPNOuGgHjGJLqdQIjVSzDOFyb7dL/6w7552M5jb58d2Mi0N265Ti071osQ4nVZ
Uzgc1QKYQmZALY72Sfwnywlq1RJtqnYaBjfrfH7XlY/2GJA8v6Ex+LgmRhEkMHls
Q1izHSvdFnv8Il3bMhibZ1DvCaC+QZUEVsZGCParyrkBOHPMcsHo5WzL8RwIUjia
jC8UQZCm0cwdvb1dnt+qJixUvHQVQ031yDvy/AgwDFE90iyR7lYRufLcuSKdl8fC
J17I4eW18VbbBPJH/8zO64rbklB7vr+YdzV0/A8A3/g9oxZsW7RW/FO5xiTOqsDq
M+tvOHZyww/m4sXirTxeMfidb73bTasfEVmDo137LSELXInRYI/Q2tIQa+Hc1wbU
edABEwV7DV6OTJcVBv+PQLEZkOIpkRO3vHlaV+curoVhsE40E7y0YLLGGPlVEeoU
0gZIxGhcMVxgGlsalmgJUqgzD+NI8Xbqp4N9nOMFSY9ij7rxvlW13M4vOBws+sdw
4i+YaDR5sbvHk8WBwNnJ/5epK1hj54Gh+tPPO3R4Bs17/x5LZAvDULFZZ2X10JLb
hUWNixwV/gWJDN0TtNonXT0oGh4ePc4LgovwWZMMguFs4pSu4B0s74zVhH/T/ZlS
8hysTv4txXOEA7v4JTqVoOjPWXEpqfJg+BU2jOyIJh1FM/IvbQuMCpLHjW0nwtkZ
LShsAezke4TkRRCFGJWHylS8KufJWKvI/kmmu6NSlVi6FQ4IfcelrCkVqpLPRlej
HSlYYTl5UvFCG7gBE1QqUBN+0m2bgCtkP65VO1L10vv9cqX0tknVge/Q+/YQBkC/
9NhNqVcM4V7RBBbtQyGAj1sGEstn6dVVAO0mGkPNpoGczK3DM+44uy5l1AT49lDU
fNpWyS8NLNuUNW9awi9frsTm5Syzg6n6PnqMSG3su158DiJpxcy+Ge7vsPRgoKOL
DA8fjo5yqsFy83cYan4K6q+OgJd4y8IVMIKzphG1QyK3TMoU+2klCKLvXrsw2MYI
/nmGJyDkiuDnSB3fU6BXi1o4pjQ6+dWD5V8QAI1KhT3bJhR2fcdc+JR+DWM+zMWV
7XO+x1czJdWa5gbIK5QeTSTVJZfzQAKGuvqZFYZrKltE/tOpqtVlnFk49Ga+Sj2J
PMMSO8XkDJ+izbb+n50gRF2hn35IPQd2IsGuC/bLSnMsDH27irAhco3FK6Fu9IkU
4XwESvV1oiz/0lMMt78MDUcW1t59Hr2OosLvruA9SgnJcvmpq5cPKvjE/+VcLTB/
nKQ04Kwxy3Tbn5IUvUMfqbEHKMSWuBciMcslIt600PrZnChTtaR5YB2TJlUgT79C
Y4Cx4n0orQ1My9yvmS9PI8NEitkKd620nHs/QQvoPjnJ8A5lZRN/zBTZ+tvXlPD8
KtaFhPSSPXlSmC9wus27JW1QZTnpoadmccO6AQGCL5Ahwf92JAMj7QeuEQXp2SOW
GmvjraA77dKWdvfpcNm7XJhq+bUjcJ5yhz/40TJ12SiIY5Qwyn4rhTXF26/m/eSl
FWLi1mDCSel72kUC2rCu2hziHPtEyyn+IfQEE2M/tvWS3RVn33GQCjo0+JEPSjeO
gIHIwDapPLDa3QCT7dGdhuHDgxxArj0wXFjWWT6JChiA+hoY3TpQEcUbkeJBFDLV
m3xYrUX2da15bTY5Mb6o+9nX6z0clm5DeGQWAj2EsSg8wK/yDCYAfeLEOsKEcZEx
1RWI6I1Y5YpW2m3ihUw4Wt4Fgqw2SbZjyy6Yqop3tXTScdTGTnaWQwxDesbXNANS
NoyZZcJGnS/4oKa0YCYm6oE8aQqfflcW0IK+RgLg+v+AD8BYyPca+JEIKywaD2nv
Y8MC/aLN9xwCZIp6kwLzCfBAmUxhP+HTHvkr8FdRneqlF0jBxDaBAgStvqLlo0yk
Og82VK2veE2r6aT9P7SwDzD4bbxETwbPoA7CynA7+Y+/jWYues0Dkd0p1VqAaubH
aQBNxbOesQNdpadjTY3ncu7q39xeWSHUrgX2hYvc7/Pz3zMHiJJB3QY/33l41L7w
7BJzwSGzJExPWq9SV5G7IQhRv1tVSNGf06Ud+DtA8a4MIsfyAU6xjdYK8oqPglst
bzbcyEY0cbJkeyu174MgTpTKsdb7yHys58H5ywJbfuso27Ib/l4Xig8DUhZwqmkm
i9vtikNOcs5/zjavZvVsb48Ygfqei5q14pJwsGUm8e8UdBHyzL55Ix5yArMI078J
FQU2FIPyWqG+FUwrNtfDRjKbRFvMuMUUEiys+ftCKO4LXABnj69gqwuio/WlQs5v
22el7kIUnztxlqILl/Hq/kKjzZSn50z9TKrSxjLvyMrrN4hY/CzeGxBDvKxwx7uk
Yq13jPeLffc9ndVesUDIVO2z0TwU5CzaCPHsbI13tfLIEe8CT4jPOF2IPYvxzOGW
/sIhlsXNggn8cMCtb6o0eMvq990zB3JkCJYQ8EGqO2LwYHI3oOhfnUA52X0c10Bi
0SJVAyHYNE6MuqrcZjj1IiAbGSZ0vP4KBwQHpOULJrTfBiJl8nMfD/Pk/acBrgHY
z0gzidwPgQVtxXI8cuXEGZFnuu5BN8vO13kWdzFdNZkSDzcJI3bHw8syII2y3Ix7
gJt8N1matscAuqah0Lo7jI6gTZ/fJ3q6Mpu0ZLQrXktlFR5ecoHv7LFOkw5Mf1EK
t0NYd9Eq0T0A8Yewwz0k/OfJ/a9XtN8QWW5yhjxC7jEobOKR/TzJUvCZgvNdtIkC
9V2HwCmPAQmGnVX5Ttc7X83fiobsi/DzBQBlvgj6sXPUJj+Bjl3l1jJnrNRwzNB2
+doCjCZtxua5y7JNFtFHpbExOOvK2IrxUTfMEnmPZLy7denG8zpMl1g5w9GkzSrK
daFcAiuA6JYEb5Z3DTnl0BHI74w6kDvJclXxliV0heNuaVRupLtrAJ4gdeN3E/Ym
d9qaL1v3+5S0COxhkAYAWOvJGZO6dKEVWrH0cDc1Z9M4syacDrMJj/1rxTokjAO9
u7n2Re8fLHwoaDl7vJtiLndsKscgFnhAOQYkOAahBVZdr9ZXNO9nxlz5kcRg7aKa
avkOPcq64+Q8jBiv/Xdw8b/g1umDw6u09cHheDzXsQ9LxyqXKli8hqpNzZvySK6B
A3Q2jE2aLOf5gzqWwPl06THIFug377fuhKYdl46qAxRzq7UeZw6kS6JBbapHq+xc
YJQp1wQzNUEzbbs60quDxczw94QvAdgQpYmF2SkvpvWjhnAkFt/qymAN3VYuWrcF
9K9H72DSuNdSDG9BANOyQoLPaJM+ImjDNU80NXomsXbjmgEYDIszN8f3BA9j3j4E
EdPP0GZjSmFAdN0GdRenh6W4EJc9bTxBdszCumCf+hCQYZMkVsHDBovv0cS6xYN9
/Cy5KwLg4ZZyI0Uck3f1zRFOPL2C8FwX+ERBebmqXUOZQC+e898/O4ggG1htblZj
v50HRho72F5jRilFS+HxR06UoqdXYSLOPnUIyUREc/mhqYzgONqlepcpfGohRmkS
AknKW1OIOicwh2DA76csSrKzi4K202svLiy7dhbLSLYjViChJ5KUrpCKR2PkZ+4L
+CYok7BvOyFUuc8fBJp6ibGcCbT70wD5RAznOIi2S+x6wtBEB5a6qwTvsCk8Uix4
Kto/ZcV9KHX3P2QxZyRLK3bkXJkxjUFtKWYmLyfqvKXuWIj1PtqlTb2B1mZFdyVY
MdQkJNV0SldswcrXIEHWVb//Cb1UN/n70dAIazjIKHLXn7cKRlfo9ChYJSI6StU6
oO/mVorL+3a8X802nv22B8DgoZipmYrCSCZSY/+6c1NZ+mGGdVVWVq9wQ+8vTbVF
+2kcK52xQjqTsmM35t5Ks6yI9YZslq5CtwQv06CmyHIwO+O53NKfIAjWZUXz7x0c
Uc8uFMLAGVzgXPTcIRUHL1mrhfJcqoJuyWiO6eIW/OMtf2n25us9TefylcTyyefA
auXqWqCopp7hJIzXLVYGL8gpi6MCwSdYaGvdeqi2ydBTQWqhN5Pe09q5qg1Nc8/u
HxnOaiq7F/vIffMrhRdFgFKfnF+PDa6l9MH8A1Ajeb9HtSF+DnwEDf9JfdZOmWwo
YcnulRLCL9uvbQdOWq7UqtPJv3y+ql91iwPfeXJo04hsoWbnGoyjkBmPj24ElPX0
5GExgurlPsqd+HaZarqLfoeQ6MmuHjTFBAm2lPQbBT+tWEOYEJbuqCAiz10q4P9i
ycxAfxOmtKK9o8QloDdWHrqIRCpVneEuipj9jj0sEaXU1FzLCFoRbjgyas60XO1s
lGqA+F5IRyds3NK3nk6W9GMx4J1XFwKb4B/AXZsAHO7zMJRCFohkOv5nn9FGIxt1
Xdka+kVW4TEfykSLyxoh2xHctqGi5vrfW8NSiAHjKGnLE7T9Ha7frHL/qzb2yDQQ
Mf4/oytaemZW2MeOtyPiblzqXwpHxh465uzKe1nPn3xLB24pc+UDxS8StZHJv7qD
3ulmp4d46a7wWC114xyx89xNATUSfluZggtFF2c61lWbt9ulouH2l+xlvyvkJ/mo
mPwlkCJcOvb+f5lRXM+U8nGEsQyf+9E1uThfBjPlggemFWnd9/2n/4LvQ/VKwpiP
OZqD9PiVaxNwlcFfixrsYSb1h1J/FMA7oSN+WeqOEglYFtD+pkMtHsIPmyWmKp9+
GNyMZkM6+meX6WXDpAiMyvTjUNz7lrkAFpqWMEgG0hOOnZJtyoGcgHf8cgY+Dh+e
7uJ+WMSzmb/PljAn8EHWL8sfuRNcGN4s9FCGumD7ahuyKNF0U1N3RpPuEyTDXuQ3
r3bkmC2XojLgm8Wqa1Vght0mIO2iJhl7/lUdTmBfoUn6kr+4H5p1L24wya/GvHax
qsMKa2OhWlfEQ7RncqAbt7a9hmPNFLcwHTynS0CXkvEzxitL6JeusD+kR61Dty5H
lJecY0kczmW0wDrGa5etq+GvNDCeqyxNAeazwr/ODPi3PdgFmUjbz5NdIYH2OHMh
0+H1sXeZgg5qFKXW4maHOJk1CVprRTil/lPr8isNiJQAs7/cSYeDh2ShzFA8lbrJ
1cqgolJHnVUygiSMhV3ihEAW+xk7075+8QGD0kTFlkojbMH5wb8wTjW0o5KBr4Tw
fWo5SKsXVpkRVQfqN2BUF1YnwNz1XFbAuooeMS/LTCNUwoGTdLW5uoTKlJAh/Sc9
nrKU+a4Mh7C2pmHtdkRh/RwfVU0TLFr2+XM3nJ93ufHSwXSe4emizOmJNsidh1wq
jwnwishFxxj5M4OjnEE8az6eKk2KOJQKNd04sWFB0grYA91/XhVI1AZ8xef6GEdV
VVL8WYU5rQWWx4Ga1k8SQQFTRGSjqZBa5jIaRRPLXllDncarczdDWlmVgHca8mDL
Ce88MMskweyCqDlJHro0WbXytqj8NThrNlq4iuUm5+GhtCg5BkQOYCY1pUzGbjR0
RhZ2wJlfXu8F5JPJXw3cTNwg27zeyi8/aTVAFbjcb7NZDQXDat/Uhbln0SijUlOi
OT693r6LQHpfE/RzzHgU9igqI/KGmQ3sSpx/OULfl849dHJInMwriZw3XixUK8UK
DVZDXjpGYYf3mL25fmHbBeQQ6w9vgoeQlhgVxYw4zheXw7jg826VUgKOoOt4ka4T
gw5M6Xxb+w9C9+BSFI3o3yIi2FKoyfnt7wTpRuhYi4JTbbeIT52gEHesw7lLRFql
TfVxY70+R+upkpRKemxcZ0f3V0901T/wCaVGPV6pbmUVVbGRhzQMxH48UfqcMxtY
XEVOjQAGPnrRD66kESWNHyDRXm3U/W0NHQoOllNrIHf/n7caakG226LaZGRqyvfF
cXFG/PHEpo/iFvv7I+vpZe6oGjMT8U2NcUsCDhieX3S4BeBUSrXZwDL4OkzHMCLV
5gemro48D8NxdPcxLchNZvzhbiYEZgsF10q/XIAxx2TH1p63ew4S8xek5qoPkmWY
q3aA+1dY14zuaVnj+tzjfQ3lWEEZRV3NkIWTZKxJtmnP+tMZsyqM/o1W1nNXRUYK
NeN7WKeRRFUQoofD9GD9vORAU6UvqfW8FfWE8F83wTL1ggl65Rt1V8kfLI/ZGIqC
eaKxv2esGW5BiZ/xAZRQWDO4bUKuCEACfbC1MitzP/qMZTls3Etcvyw1gUuzsxzE
EZP2cvcjZqvCZlSZcHMXnT63G0Y3RMgGHKMQ/0h7PIk=
`pragma protect end_protected
