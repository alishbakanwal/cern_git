// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:05:29 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
NCQOJFcQohA5SaUgKuPR2G8sxpWbAqtkQQ4nUUZma1OHPh4iIToe1wlQ4AbhXuZR
xaO+i8joPTsETI4TF6oNIbfy5vFh5HFZKFbsyWapxPVf6dx/c2p8hY05yja+KmLh
k5ryWMEi0YSP4xdH4HAjzyK2su2fOj101/nr/fKnjD4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3072)
KHFD41WWcwEpgdG7GIU4i7k0Ty3G8wSKinP8//zYPNNTDI+ahPo2mGA1qREXd0Qh
0L8e7H6YvedoYQtvsvFoTjJ9+3oSf2Om7asTsMvkYZSiLAYS6mV3Ch4AJVDzdj1v
zw09Rv8dcUoN7tiLSaEHnzECnJlVJTe88mG6FTSzViCYbNCZolU9+t3C/5dW7Ex9
mh1vQMshFGD8x18C8U/KMDLRNl1GWRg2zw6T30JvScQdYzepbu+UV86nUsqdZJbR
gFNdLs3UhSA+GHOYi8wMVEWhwbepWWEh4v4Bt+13xO6X0mJXpGdcs+23DiUeOUDk
RZH4zaL7vb1WM5dV1d5yL3NolsumKghfSDVlcNYZZU562XofEJLzzwAIAJmCuZAD
JiGE0liat78LuHKaKbKwRs5CULqxiWRrDqqEq5ryDj1PXZu0EzRMRCmiX1xVdcW5
AC542klqZuF+8O2jRtLHJpqMUmksMsXO9ekcvsdv1OF1ALnOhhYEQiHyAbdELDm2
kV1vsEro9UWOmcUTmBRBsg4S3Zn8XFmFE7tI9A9BtsvSeFfNo5OpZU1YDEPomP6D
p4yfxeJTcpVF2/wPgrYETxe2WY97qjuh8mxMduP/qqIcDtwbye8C5uY8QCtXF0KF
HvF8e9zmn00Vj1ODsUjfX5uLC8IYxz4TK5dbB7IKWurRdB40iN3X/03+NzJ53hSM
PTE9cRknreof38gxg6hv/ov+8tmKkHYvkSj/3HJHUr4AnvYY3waHGrU+DjPq1RiS
FRsV/963mHMsuYfhKtgh5rjGJ7jCQUSxExdbVMG4wQL+eGuC56q8Xo/LB9gZbntJ
Xgv+XPz2TNTn347AcHG7bTLxKgB157rhRdGmhHwWc4kdKvlaWqVLqTZ3+MBRLwc6
vVMHU3EWVdyPlHY2Pl2TkFPz8IhxnU4ctZF0LAC6ffFVBgtAGUkVT8bjxuCMNUU+
cYld7rACFOzQGJzWHrZLjo56u+Vulzt5eTPqHSkvtmuc+QJv96OJQSOJeTLz1cFu
tCWtFIY5WZm5goVJQbSynqtH5/zQmGPh5GmeZkBdYy4Hk6LUgAu9/GLtqVvj4Zbq
L53ucY7gExBgHmVI9qEJxGMd16GwHF9ce48iouyoVmFtOdaKnRbMZ6AD7tEDDPUu
Nrk8+xc/Stb8XjkvC7r2zK5distkZX0WwCX+HJ2VdQW2zWrIfcvet53/qep5jOb5
zclwvtOqkDnMz1mVriLObeCJ4Z/Oz/OMHLQ1mP97V++LxG+oA3geoSVTacxk2ipJ
gQs+wjHulPLqmdEeauEHs6QzRU5Pb7ipHe7+4dLBvT04u9AKwIneOlnGn2ubeSoX
vN7Q5KFc54yOrT+U+9F47tXL1482sRobAK//s9KjnKugSQKVadHjRPINI+hq9qxQ
OPEJX4WsRBfoE5jLAdgNPMhr6tVMnITP94Q54+cTIxYbbkEA6BPsFfH0BsZhz6YQ
12fSvASR+EgbfxFtn9krb5ZXWDj9WZjRRUWVL1ypydpRYgy1EsaNDKtatNDW/FiC
jKz8aRnCwr3UMU3fT2+XnWO5BEMiMC7MVqy0VVkmmSdYASdba5yWZBcvVsdT5whX
RD8tPd+WzQeGZmHQ4KpvKGCndnI2hhjzDVyQrWPVId33ObEWv5Fu5xYuGkMHmybP
I2znwlyTQxxOqsrXReQcznQDhLH3C+AXUe2B3oX1WQn+rPm+R3SvIhyiGBwgNTRG
6KujDVPdNM7IbMbmgVWIbzIqOiP0RfxRtFUWa8wgByroz387PVi13VwqMh1sMysX
dHcPX6zdGmfWw3tO1gGeYinlXh+vo49s9s1/+DjPT3KbbvltEFSghAR9gRHImgNu
CITmqcZo9sYohkLyiXIBuegCQDQ7kGMxIjdfh3g/aVagzx73T8msadTLZwjTQi78
4St+X3GVMBFJy9aKTPuQcgSh8UIHUHCBWR8/+UM71c2NrZ/BBcnKfGM8m711Puw0
9isV35C4m5xXX3j8DA3sNmTo7Gia6i2s2Mf29L4tJozs0s5g2kN5Z7FoEAiSs5In
x0QqH8LSg5O7biqYQf2Yrz4kblq4BTcJnvYLWwMDSA3ZCmWXk9MHOGCT+UHjRJnl
yb3IBU+O0R9tnYX67Pcxohiu3Y7XNoeQUr38aZ1ROf5bR5yxYaLsNdgEbmDKvF4S
g9C3+0WTTKMuybburWZXqe+dYYje0gjPxwEvf09o+/duicCOunKQS/rDifWPXHfm
9sG62k1DfhGvuNu6XK2cYQ3y68a7SqhQMxTc1XXDs1vI8kOJZ+j1/ti41ipWsdJF
yiHXxWk/x3Ej6jZOx0Uq9QCOzeqgtfZjUIo+Y5Lnf6IGZNtKy5G40lyRK7aG6hJq
sbKUrg4YpblsJbdDqE/KiXS8leWh2kM2SqtqOY+2gfls4YdfNKHy+Vn8tTkLgEIo
1LLRge1asWCTm+PcZBDM0VVQ6G5MZ9dDYzLIHHCO4yf7pkpgVPHTbVzBy37hgGfu
7YsCKDvrhh9YTJoQP29gZai8Pd21yp37l/F/zPmW1wLybGnpAuW6j5mVKY4jA8HH
CtxpbFZ2VuvAZx2owB9JM6dz8xr10VolD6RZJ3gGewWAXrPU/b6mcsbOVK5kfJwW
YIlE9JfRuualIe7+BERaICMVqBTc4PyrzxEUDt197EcHEQe6maCgiV1YNl6WG8iB
XfaCGxRql/42jpBuLIHppBazwzDRSUIYXJQLzayEv36UTIEjahUjKHJJrwK46kx1
miuHCBs2CLQwoq+nX6HDlFkCHLuscvenVFmzt8zMYIlU7xH6k6jerQtZJKzk4wk8
4L/1X9eYOPiEz0ayXknK0dCbXS/ZmSZx/NnvgEMWiHY/szp7zSdBayZDUP0QlJP/
nwKxZhuJelQ+2+qZW5UHozAfMFjD0A5dKf2u2oAfzOjuzcmp1bFH2LH6TNcMv8pM
k7GZbz1dfevBpdK+jcLYoaUWiRN9mjrcanKWYmVyvs2pz7E92joFbHGyjVcYr7ZL
nrieQ8LVEmkHGMc4kwSjLhx9mluv6zuk0SazH7LHpur70F16iDJ9QrDhG+8SRSc/
A4pNdHUqgkqatni9wMgeWvmdnw4NTzM45OT/NtK8+YO8+cPzRhFOMYw0MN1WW5zs
Z07VB8vd3jcuYNRTOatI/gJUKoUEEWw6I8AlR7C+MX6ESFj7cYzW51KaERlvxRF0
EjM9aGABevJwC+7U3l1WZf6DtGwfHiy1e0P2ZofBnE94SlTEhmiaPtC6K4LRypr1
BXWjoCB2eEKi3CVuWBpNbhg0SoOCYxy4MVn7VgwzWA4aDhg6oChBfrvnMLkuTV+P
vnTxLypznXrWNFWYX+E5Tt06OF40imBcd3lf/UHzb5AmqB0ZRYz+1LAQqaaRpfjO
x+Kej5OWxR3wln8MTk1itR+njnGnbXJZPLHXbXNeuJC6yfRD9xyuxGxJCC7rXYCi
a26wm6FepIQ4mVonnEDDXM5QnxukpKaP/hh+avVKqIUBLbmSmO8ThX9H5Gab2FGq
R5QxnozDjuCf7SdwYCF4rh+zUSt4y58fj3zqeuSi5ROF7AWXMi+FXFyq3/hWBCQp
qgXpXLCllsiYbFCIvQbBTy0lIj551ayslElnPFGSH7BAojKM11+zcNuSDLD8jj91
184OZBJUA/GXjqW+FxTps1EkNghFFoTyRyhtT86kCPy2IaO0TWJihwOsAtHEAbGU
Jy6jMkI2bceRwtqjb2Tp9dkl0xLE67xoFQtW4NmI0r+Z57n2AbEMQblkWQpc4/n+
Wg23ShtWhcAsJyaWYET8Ve79+i5PQPZgyO3CUhE1dyXgpQl0VskeDpujqbAf+FHP
cHrCtHFRM1PeMCENqSA7PvOYuI2utRCB5FIn/kE0gNxnl/780AXm9wgeTUxGqYsN
BCmrqQw2NZb2kvdMxqlobFXWWy5Hg4yathA2ax9BHg06jyZm1WOr1ZCXmnJH4McZ
VXiQoolOvcpzE7ofrZWcIPPnRv8im39aqIWXpqqOQ3vyOLMbIhzlUxoUA1mxeDBe
7+wAMh35SQdkx/LaVkKAAIb0AWxukGxiUFBnyTL2xnRkVWrvZNXASx0k4H7Zju6Z
`pragma protect end_protected
