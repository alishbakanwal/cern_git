// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:05:39 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
mJbrhWkI01mKm8QJkp/RJ8DkDY86H6FHamYZRjkxSvvL/YpKmv2CVKtR7EW7xxZ5
nncj97tyf01UZsDMMYSVbIoWqVQRoSqC+NDs7u6mYdJZZ7raDem1iqYn+q5F6l3i
mxVGvVuF8wQH3qgFoYvy5VPNiYhl8Kf9DwJPpkBWhvU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5440)
zYrfWTWPuZjvfub2TiJJK/8zn1gqvNU1999WR7G1WiCIHD4kgqJL/sbz2xnMBEmX
2o2l9VksXvttfCCaTCh8xbOIMX+9foKMOGpT9/XU2t++R6UpNI4bE+AWRNwcIyld
+4ZL/2P87NyTnTKBmwV2fS0p+2TxZT4QTb4CuzMQ4b2lBjcNgjcYeVZt2+Pscbg9
AAGuLr2gXMTqbwRVm8a386448IDKJynkrp8az/nlWN+GYvYZCANxNrWVgC435Ohf
1xSkRnZ5fqoIKawI2QQ/6Ow1rWR8bGsLgZtypXZ/DZnBIwPsiiZGDFFuSz3aj4B8
oIFsdT4qs06gilEySFiVwdxM0BYMw0BLHKp4kBXoQpGjsxb65xz6amOyTcLDg58s
NFSHXIsA6O79nmeDUfhz+rsylcE1KG9WXfrkWcptnvhQiCQD2fw0cZFh1IDqAQs9
/sDpd3PghnSKjCO9o+SiRgtX2YW3hK8USSXpHpWnJc38gRMwM7PlcFeqeOHudZd8
M+imexBlmgLT3X/81IDk27qc+XXHm1PyKEoBQKkHHYj2YBTMyUyX4kn8ge2NzHO+
xDr6rKZ3uQ/HVOJgGT3UZ9dhxXoFzGtAElnA1HfIH03DdW8H7EWP+y2hYUgnEZyS
Cok0UmShK/f8LW+UuxTJF4D03tGYDjSc2GlESdWTt9dpkIA9OjjcZbRL/LHLxD0K
JvNi89sQmYNWyrl61Cq5c4Jfy4Ciaj7EBqikXiqtDGgRMyndpIKWiFYhiKOBPh8R
TJanfbPZ9t1cYSkeR4G9igWTtVxij11jZbYc9wHX6v2MxmlEnzmBDFz1FERJU53T
NQCRiTmQTHyYVp4l/r9S0Xt7F63S+i4NaS6Wk+wdAAgMbEkJwcHS4LukxWsYM8y+
mpKXJJGGidLm8trswviQaab2xdnRLRs18FjNut8/7JgXhKrx8KIpk3sI0luF4i49
w9ai2DK2pwFZHC3myRpf4vDBa2uZYnzPQLYuTxa3AQGzCY7ak/EOhxe2kl9h1xHa
dfEfPJZaB3yCKf5JMODxIFydDwxUDtgsPl+Pm/brbtCcXMT5BnaMx2tH7vYoB801
ecahX8N/D5qyfZLvJWZk4nI9J6AL9YIFqwMsx8h9rp+uYS559DxzAOokyxHkty7D
zG3tuRYh4Zn+whUp+egcgR3Xh9q7yxBixSMptR9pxU966hIIQfklcjWn8SnBF2uL
oqynGglF1FLeMaBG5OipcT9evlubEs8JdNsKEfCiLF3+ES8RjlqlejQRwZCXNAw6
baelO+VaIZmGOwOcP85Y9xT8AFyBogouZsWs5BcghGT10Ph9zz2leQ33wN+EVgCZ
YeZzfWxavs+xhL4XGujXCyC7DBG/gGUC1EzaSBCWh++kqPWAbKTGnGO+7KZcy+5+
2vm8TLkL2/2ahAGNEWoexbDmeqKK6aLKGI2HFtO41pntPo2s1zNs0F4rb4ct50Ut
VKXm+me5UBy6RFbJfCqh1bloINPrmAlAtmJ0OW0jGUvHUG1tTF5XqZGkP0AGzGRf
Smbwzt4DWWJZ0LihkgALtZjtl8mHjXJ1HwO5cehjAC0blFBEAxpeI2YnC8NKYauy
0rN7njtOJT09CNVjkWUQGkSkCLs06p1wW1iXB9AA35PveJFyi/Dslpy6h+lRUnCl
i81/+ldTSzpiAbeKivJEl1LHygbbC8gyS/KZzdRv+98qMv6NHmWWTKrjJt2ZSrO9
3BJtCU1rYiispc5PQyjT1qdZRRY0gjNa3nOJZm+JyLzKV7IUV7vifoCqcIqpdfzv
rWiH4coDKgzcafyB2xNNO53yMhKaqEkmuZmWakBX8GTJ40cOx/IPE52lGnexQ8Wj
Nrmj68GRR7ImNiOGYwahVcN6s99DAj+VEoqkHMPqgTiB029tERYDHZT9brVghQsN
Kv3FCZ8++cvbK7IZSIFgG5kmGjWtWJvtVhvjX20HWo4WR7QaIExY6TJ+mYJrcSBJ
LytMgaVPSo2YgeYJbCBPA4yZOVlCAFOjUbpbZIpuhlasWUbikmmvJ3YesU/ny46u
HmJVIh4chVTGVNlIb9lslbIibBYOfNngOJoRLkay+LK3umgIsM55y3OHIelB9kmL
c1W7fvB3u4fB1crbHF4oW67YKOM2OeZKEtRb0yKH4hMt50N/kxuNS/hLu0EI9tpV
JEMXQqFPt4t71vGrJRyvHoHEKmeGcJXCs5xacDwD9Bdu82alxHALOzfznZAHSqi9
WLufxkC2iqFI9yCj7kpTTtegxyRQCA6OYEP0b5O0W6Jak3tjlSAEdLR9PoYbka9p
CHQFXOcNhuAVA4LA+rXBTiTJjo6A+SCv/3lrgWZpG/rVbo0iQdpeCW4W6gKep88K
HnPW/5RdnQiTwYbmOIJvC+S2aqBS12FmdZ4La3TFTbZjApEaDMFrvr2CczShokR6
O1Y7Y8na5+NXfa+nZ42uIgivEh5rXbBfe7xUnWw9U/0y70q89EQjuh2QnJELx3R1
++j56uvG2uhe4eYbw9QVzAaQaz/RZjTQyj4x4BZAu9voFwGMqtKREErKJvvG23XN
2W5wEE6DzMteaX0Q0R6Cw1suvnBk4H6O5ABchihyzVNmFxe1Hbwl4mUVpGhYXR8K
yh7PxcLDVqL0gy6QJvVnLZL0ZoD4UzQ/X+g2Wg+69QCZn40ltBCZsAyPPrCNNOQQ
zNR3Xamhk/jtBlbAFLrKvmtiIAUs2XqeNQhyDMgDAsCbwGrDnFkr2qnwwfr7Qz+C
AEj2ATKO2BudlBVJKQeJ0it8IjXU3eqwvCU9dDnjvxyBzwOjZxWsXdMx6dGdTtAq
fVOQC0WANjGhpU2bevfHo+2HgLfwdYo5svD8C7LBUYLVI9meI+9iS46Te+uQi0KJ
vVViK9bgdxVIbZAO6HvpxM4rGairEXm429i/9+SVr9OILllBFzf1nXEvAwVSFGb0
k2StAqo4Dyi4HOwsHaTYfg9R26dLnWx3+CVeSN2r/GX2UwSU0VflRI6mVC3c4S75
LHz/Q+jJL2D9u5wvzjzIbtXI1Jz8dHgjANYppaONxf6jNG7zMTyYgrONV3WEdVgY
QRSpuPzdzOrAz55rjJAOH74bTSn2cVudNrhkHpZ4ac4VllRtwgcMeyw87oUR/x7+
x01aTWYD21+hZicRF/YNKE8BJmFxRZTeU5gPcKbl4h8QFOiH9REzX44e+AZzGliK
MMtGFlv9f619jYeCL6dF2Q9MB8rmQYkZdcDbnYmKpeu5CyIzRAhfXQcvPdvelFTj
+xm9zm1dqjGjRDK6jYv8OvH0NeXBFI/+BvAA+G3OmuquRJATtmSLBQLaMceFPSMs
BwUiu44GAvkyrsr/ZLkY2Bpiew1Ag7UZo/kiiJ1ygNY17VmzMYPz3XLcP5FLrhlU
2xGxhnOWJKH6yyY8uyCYfBhUpttzO83V1IVJwW0ybyR4OsYPnYJdNxbNMlEI12yX
USyacvkSzvaxEUhClas1ZH310DD/D7+RaVoFnDQDb9MsDpqBSQNH8LdaQS7Y2GUJ
fbIbwvTsVbzHNaLZX9MNu1G+lWbICcI6ZF+3Rznf3q7f0nLeLXFlznpCGz/N93eS
GmdjWTbfMqpUZ8WMc8SPd4nGN0DXt4p+EXPYAT97jM36kO4Wj/ViI+ZS+IZaJK82
GXKXahNbvx+Cg2mVwoXUKXzdvvzGoZz768Nq+lCjmXmu+g5wkrcsyDOaSAlBDTC1
Ghd7kCws2TSc48d6ZZHiM3OS/X2JKqbTnF2ouJbIVmFXEtYFJxucz+0rm2owK8z1
YPxvr6FYimRiND39TxB2n931Z/v5taOWNfgisI4434smUvzOHmdR6ucpPwqtD1uE
Wci0mJPrbDpshHQt1h99JAP3GBgnq4IJl7oTMizB6nqZBDJJPUMAw1edXCNfwrMB
nF2Xz0T222P5qtmyiSqCI6bfBhTGqSFIc+veemcPC1bzUU6SFNQ6IHiIPDD4mgnm
sgp5FvZQ4EVU2y0EzW/utoW/NO2CUYlUOf0svNWpw5axpGFaYuXHdF7zeZU9R/1g
eE3SPm7vJ1ogNr4mp+yGCM8gbVg+JrAuBQnW6bery3JjfZx8yTEoMNHI6hFj8Lll
T+mJ/xMSym6T1986GeCfNiXMgQWMv1/yGoA96Go2UdGFNC8fNmreFEUXNZX4gPT1
F3Tkz9N+Zh9wIR+K5pphCIoa8l5U26jofIsPtnQYTc8QbXxEtfcU/jV4aIBT558D
aQ0Ss9jsJ4PKPwExCyWVoNcZVIOYeLURt1xQmT1AxRkxz/IGmAAOj0iNQV06PRA7
IveIJRBOkL2aYiHyZAQXxNHE9vzzQUg8SPuRE9U0blBEuWJ57azCBpLkcBoay7uF
6QHGc9IncJUduRrTGI8BR818GDC3rtLBfPkMv+1oao686kemxQiujFG2U8r6yhVc
+QfKBMN9zPHcKPT9SkqPNLeYQg3tWD43PKIEFm6RU6w8sUIJB/VhrEkG21Z69OgW
jyegum/n6FQLwr9kVFDpqvVtPO5KySe8HWQxDtuAZkON27Cn7CQ6dGKs91LdJui3
SWR9XBIauc3rCAveZ9RrgQcwDL+d9Ju5lUyD5iGX6gzlQCD2jN+MyGQehG8xQIkX
1PrLWfjbWRhVjCnActdsstzlVpkCGqzfGTM99vF5110f6Hd1U7RRGCTdj/uPpbgj
WHcRuM5DgBa6gxmVQJ+qS+5X2Sz+1Q8CUujk0ZKy6SxKB3EOhqDxC5ov/MmtXM5j
mEslDKhk7IuZijvnA61qQ9OkIflWgkIAIU/wSCuzflaTX24bCe1TTTXX466lIDpc
/ZDbxiNBsfbmK45OB77sCQMixcqWzUbyaCMNMFnT2ldAkYTKvqyBnLCocH1TITA0
m9U0LQPZORnAK91zIhXRlMsrKV5HSUgzRPCNsp2gzWCSTropihGvT0xolVOdhGFC
ryAiOodyvS0XFjH/wD0uLYyVsB+IOnLXY5evlxl8n6iboTGtNiyZBt7Ws3sfwIXV
1GaPUq7QZeIf8hshvYT5zkncclj6OztBwqjor2MasNrFPzZpIhVty2SzI7LQQGKN
ebVty2jcQr9VzQ93W19HrXdMouvQRLbw8rRBvigNEDtXHMS5LoDabgzCWqbpLERn
YMm+O1eQ3oqQOKQxrhRF88DnwxPKBFAYNIPP8iYD4pznwsgBGsHesLnwMrks9iWv
yhdzKOJ0SffcqIaTLH3RS3VIzaSr1hLHZneDenPCYBLsyoYcrIuLV6dWHrOeQWlP
yLn9S0qhZDwjlRLDXKYveLUxlf5GTRc5Ylvob/uerCUdaYYXmjbzOKz3XwzOArmi
Mlko2zeyW4D4BsPT/kvvcmXMhYQPJGDPDVf8ZuYELGk+N9ej2EhkgdplwHxN7hKQ
Vp03RBViGzWlbJD9s+WQL2Zw1o8UMQjEp5RODhvnVGY/SCYKReVOnRfBJzJ/F2Cl
mABemAjAS/I1rFS18mrdn8vYMSoezXYDb6hYxXWdRo/xV2OanBka0hQpm9QHRR86
0YYILuLkV3hflFHCTjaTDQ+T4cg6H49DH5EJd+2228ucKR4sUoQTd++0jEcdX/9N
PlWmYoIxvtwoTdql/skR6O34R4GMpjVBPTdihW/JOPXPDwaQFwRGe6CCtnh7IHgs
ILue/vdJEuWSGiqC7XFMCOm7TkTGGJGbgPA0q5u1E49NZWGIW1uxzRZuITGiHq7B
iaLAv55RXm5D2JKVCQYMKPhtJ3L7wvXQhS+GP5FJmWYg7KcyD0L1wyFEyTt9as25
lO/5eVfCkmEYttt8mF1Q12bKqzuqgrm/RZr+MmBd9H0PKg8qL82OTpyKmCUdHDwR
yGaLhhvSmdTsCrxwaLUjYqtdt7ARNvL97EuJ5F2L/6O2T7bQnGEO9hS8g/WluTS8
V8RR2pWUzmQ7M0zPobOYMlHi+0pzQhjAcXI9rBsl3WCr1o3eSxS1K7hmlPfk6yyB
9/E7g7EeFMor5xjzA+GVSwo0GlsHtUiQCRtVggotcjYHACMqKjZAMZEeFdencB33
HkcfCQQnL6hixHrjpIf4KbQI2wjVoIH3tIgjH3EogW9f+dhv7eo7jzbDwu6kwHGP
Vkwwfn2w1ko+JNwkoEJdj3N3psLEEbtTxC9Oz9+06g5XanS+jU4lUtUilK1Pj2P1
VY6DoCUw1pLcxWSzEkVSi5GB250Pr/DKL8l09hUrLtFO+z+4NxM2CXN4SowVvDQe
KoPmk5Biv0JuqlsblVMBJ1r/AptoUXtOlkLbdOxIrBSXLiRnab/rmhKuR2O3CEsQ
XPRCnOOx/0prXbwdhq4yTsXlE8SkpNetOfrz+KPGrM2z0ZhJ8HWs3jf5FZC7b0nE
7vgCLbIs0XiJsERKqbj7Q9kgBVC2q+KIq7uGH072bhpZPX1vKtNOIGGspDisnEaP
8G4MfLUVnuuhGMwd93GRgAWPN9o6qbr68IjzKd6DWM/JXlCYAEGyxuYVrRXfXtU+
SLPZLJEmgKod8rMAbTibGw273U0mTQGafaTyJL5buFVfiRk5s8EVkqs0tvNPEmhc
KszFNAD0VKIJbFyhLhahQ9JG8fVNDyqfglmKRI5fNPQejIj9vJ/cGrbmGaaaiFAH
6Y6U3ajq54TC4j1/J52QUV9DsayDgKu1tsc1p00bC8j6Nj0zbqENUAGERZ0BrJgh
Rd8QGQNKvJx7mFCSUFSbC5vnvbEAs0AOXo7jiUNL/L0AqZ1seqybPnx0oMYhASJf
OkcdtVcgYNjRm+v6Ud5uZ8eZvrGUgs1y14sltGZK/D022oLV3vkpV/KvZ104TwF6
NeygkZE9l4TM9MrZn8gZzGW0+asb0PA4DQL1MbzTMnulPPknkSWcT1fZyqYU6fQf
VAMJPTwquMvvHBJAtTCgK9ciBj1B2C3qHmtZMmhreAGA3tSpTVUgcTQJTnw3ArJc
99jVhju/uUfbJvn+KAABWkpdNPTbAxPQWIvTWU7IbqUy4wph9T0nZXVQc2Xt9cer
0WO7X42jE+q0nMPyzh/JqM0R9LHglWzThe1DJUlp4S34KuESxJP5LDbxn7NW6gqR
6EpcH6QTdAwLJ2MaJ94z3X0bMf1wZaVl4PAmfYdSYTt7QECAgl3X+p8FdtTalCYX
uGSTN9eL54QjxMYvj3dISecBRPZmCCU+zPDVjBP/hQTgASdVQv+PSNxGIVB3DWAt
zxCLOE7YNhO47Cp6hh1GR71zh5J4g8Tc6PTYCzA+758N3vNMgrORMWgWIa1NgDBY
ZlR760xbl8jI6A803GSO+A==
`pragma protect end_protected
