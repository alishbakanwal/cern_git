// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 14:01:26 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Hruf9CzUW+bcszPc2njBecEETdyvq02eFBK0zWR0q3dNCDcV1FzGieArIWu80ZVT
ugyPswADCkDoozT1gAt/LDU8h1jfyquGuqfrDtjCGuvefKpNpoGv4agKYrUOrhPa
2FeQvTvFHcI1HmaaeAoPSPZD0LTiYievGh2Kd6HouqY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2838096)
kv1Cxm7FHm9hT1Uw1FiFLUsuwi96lAyg0KJx6o4+3LO0P0ZN7G4dka516CgjaCfz
uHhjC80k4CkgkuhDlLVTnE+VVPzmr2GYAXHbC98ZJ7FL2Wmd7yhAtCtblrg0tWq2
R1QZrt/C14KXpSeTk3rFhhRHM39nt1X/u0BoTabkOm7W867vICrxApqiQYpDkNnP
go+vK9UGB/WwJj5NAA95vbwb632W2jqtPCF6jffD4I5MyBnyLDUEfwvwXlJwIjDw
rftrV5M0mn3nuPNv20SUidKII67A1ZB7Dy7GmJ5ref2vkwanmP53bLcpegbka+kT
jnFxosdzmSaQfa/axrqSvxlLHamSJshk53eGlDY7BNWqfGwFFqc5QSEMuix4WxXM
C8fI+mV2TFqMHXpwyczXRmZISyEeOsXnjCMtu71+Q6f73nNNEkHo0/vrima+BKCO
ABm8SF9jkRhpjGkFH5LmQNx9zynckjiP4aMhpLrmpyeFsfqooyYcBWolfnaEvX31
xGsw6Yy8RYAuAhGQvp2M00rBCCrFgAPWMLhaohxQh3HdZrNcyaZGp50Pwzl52noF
YR1O1IhoxCYLCWWUrIFlDpn0Xnu34X2Y1IeGCyR5QZFyEigy8glfAPUveOSCkRer
U5M5YCBYRnFC/aKrrDWBAlc/8jB97UYmA8RPtNXfiC5w+GkTQ7xB9o0oSOhncFsM
0Yhd7MBpazO+x1VnzfvxjcvwfbbTSFfhjww2nqhFFIv643eBSVdaAUasCxEMi91H
gEiWvuscpkiGf75eGJDHhKQtuw2DICR6qP3jKOocFmsKyK//vyplijuFBsvv432V
7/yKX2Wvyn7SCCJZ+weVxLErI8Dq5k86xfIsGacl/hi687aHIzqigSJgahcuAg3l
9jXvxEbgFEHKhtUW+UFf/X9mFBQIKdeSJzsciFYmHV+YBV6a+huxdGZW1VW/+nyV
fz9xl7hUL8s5UNeOBTiatltpSgaKQqi462/JL5sRqWqDz8GQ7rSENLfUw8kdUi74
SvV2IgowOLi7pOADwb03IlN3qMv3xB4TwcUTX2Mvs1HtuDzWE/u1Gh0B3khHCnsd
03EVKTxsmX/9nhoT0jeY/iU26Yke+Rk/Qbixf88SxVPv9FlVKhpWD4KQkJwyB+ra
GdAF+eYp+hb88Uh1HVVTtJcL7QmBEloHn/SX2t8kxQ2Tu/kLPF1esPmGqtOT1hRQ
5L0xcVN4hmvgXRLnaPa7PC7keryc2DuOH4FFWEl4MTsPBcC4lPNv3VCOzzwI7KAq
2sQ1t09J+cVUHsA6M+HN4Z8IksrXybkWVQPZff8pnno0t/YV73DKJN0/eL6ivHwn
ZhugJB1IjFFNyGULPgr8MPuKqIFiLVQFKomGchPPo77ropNgUV34JK05/FlBAc1l
i3QbSYG0R9/ch/BojUoh/pPlUFep1xZ+Vj+i48rO+6ynA0v7oX0+Fizza4Cd8WVu
Q7m8aGKXuFe0t74Dib1F1EYsRySf6LktCHM+taWQFOjjXRXa/ykPinyPQ/rN3hBq
jBoNwXz8vzgvYedbcMbhus1nhcftx0zvqU1F0sRdGiw+f6zy9TA4VTS18w02E12g
BFSlS9C8QNV+EwMUyB71jCs3LpcpkjLoDCMt9v1nje7fM6DPpP9r2U4ba4ZQm51Q
T9WOnQ7M1E+I8rzG3d9m74RANO1pkI1vnbdAiZvIlOHtmjuDFiYLtnS13V6mPhQ4
eCHE1E4c/PgZxCN/5vkgC746bhfRFeC4tkvHYygytBkuAcRcZChZcWSkw0oMH53x
XhRn7zBBI8fa7nyCCq7Hud0vW+uGvgujDDLY00d3bOx0hxG6RwxE4aPTQbWZVWrk
SbyuwhCh+noaaxMdb2Yfyg98yIe02xptkr0ZBNrsrwkQEL+POJTj01SA1vWzYdZw
ACTtDHcDawDrgc9hWNehJWyQoVQV1Ptzv/zSISH2HjCLfUnQKcfZSCNil6vOSYUj
gMMd31yMpAyS3UZiMDYjsN8DJI80JRwmu+nmBlGsPumNDdU6QEeSe0swV2Es57mh
emga2yfrwVTZqJhFmls2ORiFUVncY/YRZmsBmVS2iT+AeI5ZrIVaPnv2wKg/rphc
fSurlbJ8OmFUQYZmDH8wVwGH3Nhf5hw6tTLWjb3uoJdfVCXe0bz6MWgpNWvmMfAQ
QSHoJXEYL0enZ8yxWLZrLGVfEx4EF2RdvTCfzGd/iRZzigIOFz5/gtRVp4t4hyFs
Mv4kwdchxfLPqbp6ATx0V9vU/X9aHoWFtJDnXe1BbY7asL0rkQkh8pWfNVrioXjl
QLaWZ0dVc5M8lYCFEjgqtubwb+z0oc0DfyVxrBU8cUU4O2g2VY4DkpBuU8ip7slN
ZsdemOcialqmwK0A5HT6btb8z5eIOX7G2Jqsqay+it0ixJfNBWt+jXNE7o5ixmOe
GwP7RZlwFf87UISqRP9VW0O3v4aMTbg/TyMz4Ho6w7y6oeRV1YYGgL+VQGS5XGMP
kHP6FXd/MfoGRXvBGLE3SM4OF/Lz7f2Y1W0C3ItNvva57OL6sA5utPIYVChXIihe
1TfJ0Bbm+OgLZKFvT5sqIge1MxsHCtyG2/pnbpruWmtoO9G4MvE3nidrGEl8FFGP
evvgPI4WjR9nR2Z5hniOt7oIz1EuGekjPSyNOuqhiqEWhICNOYaElLbSWHsC0ELK
qS2GIJU1097Vwc9IQ1yum+uWguw/LuJBMBHdqTANKq9upSkjF2FfJJSc4N8MdROr
DwnDdEAy9yHLewGZ+RASKPJaLDjXw6L9fi/VhkQFEiAI0Q5AnsPT4tkyVvuHJmRK
njKVUCRf5xw+9CC9RcHHo+geMIZ5kl5muyRvLO0Jm8OFMkjj49m4yrtV66a7Iidi
NgLywLoJC0DDzlTCjn5O36QOJJJtDJA28U0AIiGOTg7gQDuIaX3vdZzSiY+P8p+8
exwnIXGnsNvZatS9CgdoVvO0p7WzeRG6jcay29OmW4+UiCTMQ6OB7y6pj5LyXgCk
/Z/iTgt4g5YuSLN/FVwlh/glEzTBsurbUIPIouCBVg7z2CaMk0T2vEMGVgQWMsWi
dtG6v0Z+Y5hYx8Z7rWZ5yn8fAvt2Dft5esYYvyomityJJ5s7pZpstSaKNiiIqbUz
cDRP6CuuUQ4u6Ui4ofxV4kNcMb2XVP3z8UP0wx2D6Z4KUc6Dc+4yDZXTR4i5gwFW
ZzdF2tiejfCuWe5+gH0obbShzYLmbFS4jtbfaaEFTYzaOGRFEKMJDagSzRPCTrDX
vtSngpJh1ahhwAZSmvE3BaSNKKnf2gcpEiS8PiVHPPUANyIGRGOqPhHLbT4poROq
1tsDDiYP8vo45kRkQbRIq2TiWvDyb21VcWZmRU3U/h5SdcCF4ASA54yjn5nmFyva
z8wOidj6QVm7d/r7kAEnbFvH9MkR0ByhknET1ZjnUmusZcMnq10S/HVDWIYbTLOF
vmWAb1mITlbgfoXcLKRBZAJ/vj+KUo3nz8Uq53mWZPkQGEpKXWWi6qXiD4uAuLXk
Q9LNS8+TMAyQSMyq0POXFgRx0MYI926huZuVVMIZc1gNGVFw6gk3noSNAsIWXC6j
WgwaR8uSRSQUY0/jcxVH4nzNb6sM0+Rh9ZZ+UddmeYrqzVg4LImnRMBQcHVyXTqF
h0eHgRkt9W6w/WaR5gsIqIMrFnqYXMhPE+AcgleQfhCzkU8boSQT9W/sP4hJzqaR
y793A+ElrrDxAgiRrHmFw53KRDHOq+/PVcN52FbMKD1JYLOv/OKXgPNb5sMRd0xY
bT4tbk/HQH3zJ+n2SkQGhU5iIOO6pZqIkc8boeeYaOqAIhDeABUfyR74g4hJ8gb6
1v12++mrtRULLg4Lodw+XVGcH1kbJdDUzmlgxujdEp5Rykqt7zU6FkWIy8SWWvdE
sJ6hFGYjn72vKPK4xH995U38hMVKrA7+I3QfzkTCPNR8tX6a5c3HLTZ93eqG7STc
dVvEG36BoaQQWK4LGaue2Bt9EdJewU+CpZWUPZtM8GcGynNTbTKsBLKP2LAvCdlt
7Gup+TwSeWEJjvZLzFoD89JLIsCMVWkem2JtkZfVTNMKb/yKoTTi4NmsdnrMy/7U
20mET31C6E/T8Ref41V8zhIPHr7h/8dn7PR5ke4ZDlrcXEI0xS/K03+MgNtWhFsO
PfGwNYmOYogt2iCK9bedz7NGinxbud1dI4+820qP4h2wC1j25JYQS+kzKeLwE901
nVs4EVjq/rqzhHKVsSxoUcrnqmpkOXUP71U99kPYSiv2IhgXr1a+6xJFlrfXcBNE
OOi38Gevc29SFaKO6z2UyrQDOko7tB5cof2naW+AY4imdLEY478LcsFSSD/DgU/d
X2tpaVt3cKODZalTiWxpVbozsVzF9YpbaOJVmWm0U0w59Z3n/KnzIxbcPi7C2GkL
lqmyPtBAEFX5txt7HGc2rmGUBb4QKKm8IPP56EGZGBrjqz91mgyn1WlVboiMeMqM
w1wZQBBU1TJq6u4xkJxuIRIPSKp0BJKaYHPr53BFhfimEssUZvZpHAlI+2M4Owt+
ReXOE6TJQPB690SahVKoNVwoIbOQEBo6XHLO4Jr6bYLYyrA1prJiU7657o96dAaB
Q7fu4UtGj6E7UOelsn++z3FZqmW+eNwFP8lgWs7ePOcJ/ppD+NRuNVkEQ6zU/A09
iZkSn2elL42/5D0usJub/Z7sPLGuBRxi1t16gxOIqR0lcNGEMFwZJUgkW/KTCoVH
o/DMIxGwRw+l9Jq+Q1TbPDBAq/VT51MXTrqnpeWCgChGbNKsjE9u6M/SYfs5Hy/X
mwue/t9Isru9dNfqH/XyHPeE/qVYK5+cvrGAQrRdsZEyLX36g6c42NXt1uNvrwdR
ZJuVTvo0HZD98vISyIjlo+b+QCR1REr7j7hfTD3dZDfFgfL+t5gB70jvJp45qMP/
3wn4UPqkz9jtNKAC1QjAXAAPRjRyI8vCGwm0sE9kSZ1Op5QT5pq8s6JyduB8r4Cu
J9RwCwvWmpHxqKrUaDPPx2tVFdkEd8XhK1MT4oFOHjfxsBuwMKKnBPw95uMPkFgf
WaSleUDisvq7rmmmPy5vca+xhdC7WmwDHZUbH1ZE7Kcp7HddG2Njfe0D+tB27NQg
TfrnaH7KFmUlZ2Ng11JHJANtxAqdvZMA5aw6xNBv76QTSewad8Bn3stuY5WU0l7z
0979GgzODMcf4Qe45i7FW/zrvs8wKRVIdp0dgLaa7t66b4Kg9XczWnU+/+K1+nZZ
4NSFjp0a2BLs+iCsz8gxKGr9sC/uc3RPM9SebhCFpQByOWC7X5TfI9HSZPhHhAAr
M8qlazLeLcBuf5X13UaWGIDa9/uCcxKcB5Bz534kM9DFKe99V1k7VyLJQlo3ApGC
ZZ10MG37c3+dIjz6nQSt08LFKVfhaOH7eRTvtf/C5UxETPhlgUD6h0C4oZo0Q3+L
zeYy6Gwd7rdMyC0f5HrOgeqqSN4jiGjXplbo1HRkkqOuBV34MIUJCjVpD0JJ5+DP
Wfhl4efJpACFwj+ZRycTtFfYivcvSHs8pafIodRR4kFa6kcBp14dGajttDZW/ycI
oN5E8gkIf1sSpYMUFHhs/Xf/6sr0UWX2seIrYEDm/6rSE12ptp3yM9ZFi514oYnB
ZJXvRNHXigZ6ogg1gdGYA6OvBm2V/4j16NIslsbPvplRDEI862SbQKpueMW/BeKa
FUswMzpb9Pd3vNzl9Zk8PS1d/xcmMcDVr0i40N0ZgjeBIeikje8wx5V2dbyQuyKh
K2vBvfRFxSHBv7DQHjVhV/DK7jCgrYWhhTh9IRkzq0iRezbS2SZofdgMvVdoeHQ6
FwIk3lChqh2J8VSgs1vaQRgSAiS8aGvvC0gYkgolrMSPkCjls7p0Yj5EQf6tFfKe
MvBvBWCLFE9az75bErd/n+4j/Yd2Xjbh8ENQ0gcMf3piNzWU31wt3vlc0VjGkBKL
hKTR9tkZpdZWUj6vaA7D8ZYSpoBMAEvul0Ma6ZyaqNx+2JF1u7zeIer1mA56Zger
d5EDDr4PFt1XqLVBB6VxAjz1ZbmIhnllVmtkPHPnqB+ESMcok2lJK/oKNzczWXzQ
b6xnpdNT/J+SwCImxF8NdqCS6agzVNAaz5xbjMq09Yi8eKuF/b9PfAKDO5uebsHa
bt2C3Zsh/MLGApdT8ZdhcU6Jl9iOT5AWIk/O1Fcgai1Y/iS8pV3cEl346WH9eeEQ
juKnPeoI7laVQbBLTBPLzqy5ngjSe81HsuGIZbCNp1fZ6lC3hK55zKCM5amn4l6d
3bKq+D44l4V4/DowtmRQIQ8ZIeMBzCTr8yI4tEzkyRNBtZd8yO1n2OVWgSKCjT0f
yyxy7QyqSUJisaTINu8FLvEWq5V2GWnu7DTfqKgcbi0JZaoqYwMMwP0/BqQsIjHw
tzxW2/cW5K4is89v1lmbBVmnNp+Zgbp9RrgcWumR/pN7I7jie3U/N6u9vTA0bfsU
GnnNvwMQdaNZWQn2LFazlf38aEiiwQ0RKf5IKHL+wp4V0RPJQNnpN4PHxpnuTniq
2++1Ez2HTQ/7IKJE9pA3fyZKtBgFHG95Padiaiul6MWlch2yHOjUQwZ6bCLY2KRt
XHGhCH5Eu45aT5D6AhqeJSDMMNjfK5RX8PRXjMLrEVEe0FKWvkAb6cbXX6sf2CrC
s4YkWalozgCmpCWvL8Su9YmR01ncdrePbjAex4v3cCswh47kIesJBdVsv/YUCNJd
u/VAFAyuo9CDGcxjFh2EOj3zUkM0TCUlg5+8FuspWtU45cXaIiev8aKT0OUe4L/t
zxhxLwgmx7bz/JNO6BbciU3a3insyhUgfTA6Zivq7h7teUxMvJWcKQkt9mZEn4CK
1elrHaS6cZclgdftFUY5/qnVUQbrON1D+8uOXwt9e00Rh+UJnu7Ep7LqIKX0c6rP
u1KN6zkDAaWMaJkzZ0VhB2Jy+eWdrRAwc5/4gQ4McZno6cIQEs9tT9sppXh/vbNR
ip3lYmjlucpOb62YX8lsZohVS+1g8ooFrxQiAeK2neo/ULGP9wh7MCq6Eqiw2D9t
E0flEm+LXbIkt7c/AtpYdzqVowbAZ4jN/52uuClC14cOzT2gMazTXg8E1uurBty6
J8iEK74hNl/C64Sm+OvQrqNJmESW9pon/T9aPoWYDJ567ia1AOJ3V5caET/GR9WZ
SV/IC52U3gpTxi85G3zCeC2vj/26LujOR881rrUoUh/Gmcv81fwFLjjfKdaKlZ1C
ispjuvMVWeNFfvUVvUp+tLyATpHshwyvJ9fCxasBy4yuXGqfPXxYzdnDkZolxCJ7
PXZhQJ+e51p6XigvIBR+e8fg/jgZLzqw2DTRLSWbgW55cO0LVuKHNgb7dwfY3NS0
skSo/X+36LRnphGIFRJc5Jz56OAjHHrAZxwwl5iy3GWwPp1qSn/0PQd9TLnZ8hoN
m4+22rlc3slrt1P1xfmBKN2HhvTNJrt7vPM3VN2UiS83jo04BJ3ys7SxGOra7McI
13+0qFRNv/B4y/f8kO7IUz7rUFrrHABQbzbbQcvnSZPCO1iUqE0s2J0EKZ8V60TD
+nJy+9wIyXbRt+LJ9KB92SEWJN5rrOCLqY5eLh3eksUXYnLFAXC3Mb+rHqPHD0MU
bxu9/gvX8uYaEI+ewmem4sbRaialrSmgOFGlO5JKnElztszcAarKpfHIheHPjdYr
KfNq31ZBNMkAtN9ic15Y6mApQib0GuSp9Se18XpM7iQ5DD3jfF6tn4M1wOJMGNO2
3Pu2aRhhSv5VYtpyx/YVyVHB0ar6L/PxLjVk3OPtuA1mgpTxayqmtIEOLgTh5yCR
T5b9H5yoSKMt0D4aWaPAfD1W0KP81LmNS1nat+m8io2NYH3b24GLYYbjQtgbjf8W
wJqkYQRzOCxs5z/h72ejj1HGFALb5zGfi72mJSl4yGFcU4MpQd5R8qYa0ofGO6hq
l+A9Jn5BGMmOo3t7lQeFUNrZDtEBFeufsZ/arbJJq4g1P/UPFraUOa8JvP7G3/Yr
uE9UrNXnuTKADVNRx3Y1FSJ2q5Nx2S5Tej5RzzblLf3iWm3q2RcZ3O7AQ/IiVqp5
649lmcE3jQL25Aqq9Ax5r9kSGp0p8fc+R5NLGsFSqPx9WCF8oC6yYVRyjoK/TJTF
541RFyiR/a0CC45GKEBa/CIG4tKITkoIRR19ZJTVNtdNslvgRd4zqZjQ3++GGwS3
RQejH1zQYfKGXbICJd6mXaK/2tAIRwXFmVx6qc2WR3vCzNwFIgBOvMyu8B+r5ZM8
102VG5zCTG8UhwJC19WBtweASYcYzSBHDf98BynFYdzYp4302+HErxo8ej/U5Ptj
rpjCDklF0Kt4BiswSW7eBJNnVOw3xj6Kj3jZiMptBsNXg56E10aJtA7TzZyayig7
kWsjdWN1KObLQVahS3eg/8MpDVc43KN+/MzSiFX2j+NhA0Z/WKOwkxe+e/SsmeJq
HzDkNDBR8LRQ0rKQkWTIvA8dhoJjlyNie4K25JjutzFhleAPaXZl/v5n4VqMJlzA
VbCiPKL93Q/2WMS4s1+czBoJs/wEKuOC1pbbDmXLqC/ompMsMSmx1DCr0DvtFrfH
2YQS739WOPysZNIxw0F5rFND+WGL5FENx852RajyT+v73Drbvj0zzrnskhZpMZB4
Z96DVthg0n520ldV4vdMqUrbTe8SqcNY1P90MhaA5aCZYUK8iTw/xDxVzgxisY3D
53fW5OnQrvB2ZfPomDPEqpFy2N33LhUAsCyC1Bsmru044YB00LYil2OGSD2CV8MA
3BgVdToRmCHDD8x8u03vlTCt4qfX3j9ZslYABL0a44XJxCEEbtDK1FKUU/iHp9qB
eGxUyWT5ZRb12NL3REXmOsqLt1MdLKqhkOgd+o6ZOlv1x2MTl3a3440Z2CrVrqTK
8QTM3LD+S29yH8cOEivfQYSx5mlpQxnolDP4KeAhj3vCg42cjiLFqhxH7o3nLY+m
IQvGQWMQuAtUCLnwREfAoi1HeqIcMvT/hbJLFsWQ2UTk6E0LO8/wH8IzEK0RAXtr
5m4Pg48gp46hz5NySX3O8ka9H/RGNI5hCcRw4eI5Y3kRY3McWcnHWlpQQymV/91+
jnfZOSCO76zFUA6hjCHcsLE3gdnjch0ERAZrbeV7ErGpWwkirqrXER7suXHC3tDx
BaNjxruMPYION7JRLUo9r2gaxh7UwaL1aZ6blHl9joHOke1lNPvbBOzzWusYFasp
QsX/l3KJ0tf6rQF5BjMlRISnlwn3YDKb29088JaVJ4DT7JofD7g09jKq0EEbSlcm
+Pb7eQWDEfE3UOdZ8Mfb4WdHiY0l8RWdCeGnGm/Wnk81NOLXyp7Lq5w9nJDTTP7U
6nucth6sxSC2C8V37OM2bOTsfub9GE6O5ydjUUTYgAsgjWpwLiB3jusBoYqhzwfy
I4xoDW5dmu0PdpAmW1yO4BeUxfdXecacAz0On5A1qYHlJ5vKXWE7wCDvRpDsEC47
90+qnrzWvge7Kw46AWf4dCRyJA6tMpxCraVnEYWCemp0Z4srbjz+yXaOdUZcsFoV
NkCTT/DSPaFImh72nwmTuvNk2p2QdyC9v87VxKpbdZ875CObXE/aggljM0TaSkeg
KIegn8gfUeMZZCFDnfHN4MGbedxzdY372cCsj/rajypWMc7V2u2wmDvw0TcNvmfJ
hAdWtvHqjsv9sy/EbjjqMOSOD/e/XO4YBnD3FUlLQvYRtlBiggsz3p8S+/o09FDx
VzlSTLPb3eacSgLoeEUYTVeWcahgWaNKJFY6k+0/NMcGUtR2f0SwaiOOBtbGzTVm
tI7J0VdfTcNTM6CSgWI6rmofDCVeBfRLyl+9MAwrAWpXWodkOYK23uZfgXtKszEH
liVT0HQim7boqs0cwNELtWGTMsGtjW4Ft64nC38Oeo/9cCSi7CNHbuFQgS9wqseT
uPL6yxx9goXVZRRvZn435shVdIrqKuzSyFeV1Azn8XflryXRobYXQ5RAQG0rtsOh
NGXWpGv54zShfpKJb/EEbaNLV+LN2ujVu26pPz7Qbo2/bLNC9t0qyke2fRcpKAO3
+FphjU0e2YeyjtiQuZNyLMtYvJr6DxDFgWHM6pw00UeYZkVvkLUAyet7358tT4lp
Zzi+u4KbOcQjKtbmgs6dKF38aurvkiqjQVy1x8ZqqHkCbxosSUd32QW+r/VwgckC
uSGicMPtqaw1FbzVFPLs7xFGENYOgS107AOz+nYjS0pGCK2CnLNA/33NZ8X7n4rZ
fRN/MhpfblVNxbNfwyvebxV083INFl/vsNP57zObWsQXo857Ro5ErdSy2N5wQd+j
qk4IRNO9eSGpaLroC+5rCPKtDq+vaMLQZIX/lT00cLk7N+F8+OifVtjcBnRY3xhr
xCRMqN1C7Olzai4BNiMOYFIdw/edNDl4Zt/ohy49+d5cAUAHKVaX3vn684g3uN7/
s8Mg1UOECfHkk9Qji4CPrzEfg0lGK1hrJXpkuBMlXk7UVc2fAXpyXNpZKOFyqUIu
5j2USvX8fP3+XgrSXCDT0QFxBN61tcyW8s8byu8Bt7nWr0OBW8ohkuLEqh8lBhhL
mkMJVRYywWQHibL9qCxU2OFEfPNDrlcuml2/p3sqjfXCQDiDr2qWwH+bcBaYMALn
oQBrw52RpJm6fRpzqv23KJiiucwsu6Rtif2zZiDWnw6ELl6yyiLRztGcBy+QF2r8
BWEICVbZUSZwSKP3zfb/U5eaO9tsTbvkjzR2QOHiwlhusrn1YS8CDtC6vXPVBAgh
Mf3IaHE6ZYwSJoMxVVvL7M36zPXuwGjLd98/NGeHovXgNV2dPMffu+2T+/5clyui
zOUPxi1AAM02C2d5T9xJ/h3M5TI6+DPm6O9OYWObqJA2b4EdoF9R3GCrNT/KBUEI
4+RMwq1SGQSVbM/RcIy3tUjBM5yeChDObaCuAX6zBuGMBpFV2BtImmGtqztsvoaH
oso/abRK8+7ExTldkbp9TTMSW3oRL3YOxXnNfPgSm3yrtbZuXHx4odihEbxtytaF
hXpoaOJs8DQCfPj07+yGAti/cHg3dbZIxdZNCruu/Vf+BT2Z8laFUgsE5k1VIiCH
KWdsVqj1nE5VXMHD8LXRfkDlLIviim+5PsOjH12PL5sE9ltIiG8o6IhOuCosTnju
BXD10r/GQe3Gbse9+FLLkhJii/sQNJRhS6PTAf7hu3sA2j2e1YkK3jxPI8eCEoBx
MZHYZZQN2XQ4ALS/G/EGqyzdVqsvhN+tEsm3o27yx8wzYFFbFpRi1VtRg3bA9FJ3
Vp1ZwQWH9qaZfaadGWnhukG1uogZ9W+bbYN0NYO/WqZXGUBYIhRpoRWwln+F1Il3
7feRdmItZt8bCkKznUlsE+QxkGzmolj1xvYnAbJrna5f43U4Bzup8foyYMEyYWXL
FFBw+xDwEUQiFYRJeDu2zEUq22aMLMezEsArAIsAr5tr5m8kwTWN5txUXuL3joOL
jZPQqe4lIOZkz4SQD/a/rxbedw2hxn64/jsO6keQJNvs0iqXaYNAHjz9iDExBAA6
IOoG4Rn5CAVX+EPKl+NqheXnF5ae6g7nqQpKMLjBcs0++OALnTjgw0KjqzQKWC/D
5wYrWky/FNWo6EaoeVZ9Ql06zhRiBaHlBEK2WqGoCjy8o5SGuKDg28WxQr4+jCWg
Q+PyXCW5LqYg84F6F0DriNGyvDBzV+Jt3v0BK1I1lfr7r69p4T7CfmC2hBotuRDM
vuR9cQL1z4DULGxNM+KUrtGnIXY++c3sAEOTZz2jAnrJIUtTraV86+id8eHPq94q
SEeSD11dnAtOePp3OdGFAOYROyyUcai0Zp39JLryniHEd88cWTZCssQsbTH5ZlMG
0Exs1FcPmEyo/nWs56gIHgRyfSCbhnbgbWbcZpxf1EKj3HerQfzcXuYGBkTdvrvX
SJGsff0XKG5fb3JVjn8bE7Rx84THhrDnl00n6MgEhAq/CYME6L5wgOyi7pxFVS5C
Sw8qhjEATVHvncuDfrSNcg5ER5+YMUT0qdN5J9iAjA0TkxKf+r4xSJHkh7ixiQn+
u/mgG2y8VGNqMJMdVTkRcpo/17ltTA4oSNoSZOcc8nw5FEJ7QDrHxUNeH4hTNGTX
pc5RYx6ARGjuRGz/4zVUhRhPelx+x/IydL3dU5XBUMcWF7PFdaIz+MHdNqk3iF++
rDxhpLJe2AdZrYmIhWu1drwoeai8kY8H4HVD5R64n1ZBWISdcTVwVtnjSAWqev+0
xzrbItVBb8I/Ng7evSePVATrbwbt+zB+qG57C6INUh3qGSBn11x9De+qdXgY2+Ke
ybfLhc9W6ZRKeXh72NNHEea5983D3sE/VM4FA0mafuL9rnnTR6wMaSyhjFP0f0Zw
JGZceGDA+acA+4sUrRknE8AaqCaGQ87VKzC1vs5v2QOHydYR5QX/LnOerRkw8Od/
2pDPY3dXWRKpy3chiWWn8tFEwDWFzbQ13jikYyyXR3u1yl/9JcEWwiyEVJqDHKsm
vSpis1Z/hdvWpdzlOMTbVMtvELYrE70TWTqMpFUXyaHHrFpwRWzwtycUPNHdX+tk
aR7rICSaB4xUY8c6C6op/1e2dCStNOmwHEYTjutBkaNV3tgp0az/vUdfXh9951fi
lxvTv8WR/dvrJwCB+YaRdZWxbswixPdboTF0JmB2IV1LdM8tKVBwWMfMvvnu6xVC
sn5MXiLeafC3ZN9t0z8g2/7kSQb8/Uij7OrFJ4i4+s/vC2i2gFXhJj1EX5x1eM9D
wC/av81EsAT58K/m/zmxEVSKF6lhcKONTuM14vLtDZ7XsbJLLBABWQvFHi4b5TDW
UeWMur+AgnRal4YjJzwCAyLen33odSDooczFao9U6qQ5jtfKtAOh8/3Pz0HeGUQj
is8ivd89bLHEyNik+v+euyVi7otOlGbpnSIQ0PITnh1WZvbkCgPvq0FbbU/+RMCJ
tWQq5QuFm171208JWICG2EmC47ahH06McH61yi8wz/D4UjHUv1X7Wb52GsdiskbS
fQXmSG1YmHwToT3W7h3DC67e56KPUuSMn+bo6tGOqH5wMq4KYKN/H0KaLSw0DshC
rwQHBEzGTx7WUspP1D+whv3rvJwyyNUfwLogX3wDqf0pA8dTwGphdsV8sjjdd82s
KDIJU1cDJCZlugUEbfB7sqi6fLwJwS+GUr2PzO8nl9hEUwHsyIp62kIeGYD4lcux
U8/0Sm7pSp6sRv7VPYPylTKcirMwsrseIxuerKwRVIHh14Y/vIakC/ebJxrKgDsp
VRgTRAfWOdph1RJmjBg50xAFkZOKdw3Hyl778Xe3MarOwH2fkPKchV/IgluvhM6S
+jUrKVSTh+WD0CMYzNTlsL3L99IVgVBGnzCEdC5nQT2HI67H4ThHgTdlIwBp1gSr
GH+CyXyaJptkg6WTM+8GmjCZbb2yFZQjmZCnyu8OfvXB7DGbQVEYvlrotJ+o9ij6
GlGj58jWZ91Niow7sN1e0d8D3UzomQLBOO8hxlU+mR9mGgJYA/TJ0fBaNDBviWmD
Uk5rOKJbYQmued8Zuu6GpqdKFBT/VoHPn3yhsTWiQySQ8rywrPkyJouLP9HOqPnM
D1IDHDKkxomBORNSGgBXkUjzaQDPXe21FbZs1SpNl9kyhtJdJ8R4eJ0zkUXF8nMz
cCPzxX+OcVIhpknIH7ssFyKaYHTYTQ0V6tkZRONX7T+katc/u3PPmMk5XHuGGSc0
Nva15RCFCLy9Ko0DAYCImVkVF/A75RpSARME+qmNGq6Cksv1rBt+EYMlmjVoqJsT
/6yvkzLaEiEwRVOx3nNgUyfbe9VNpSFlzPce/qyDis4t2yrz3n1d41BhE8V+o92o
Bq7q67nJkGmKbpVkxij1dCOw3FIysjpmhrEvC0jMBN86Syx5fGytfI+gSTONIyjj
fSYAu+HGjCTd2D+1did3kHIspPeKuQ6eLw0traItMsqrXu6ZH9ltqVXA2ugX5oTz
R4wEoVBT5s8vhUv/n6RFLzJDmTZOivAdVM6J4Fza4ENF8rtx7PCCBzgqlrTcY9Qj
Q1ljnXgG77R+jR/QoHDlIj7217Jn2BWLyS0pYDgf9qF+2YJjwhKrs6UeqycaOLQY
5cjUs0E+2vNXSGz8vgPqQ3IFhHbvwpGONWFtaKdZuYKIwbVTqN7wmCdRIXdLijqX
9dPXRKtm0D5s2rE3QBQwfYGDI8ZLgdABFLJJFWlGbBNJVJ1bg3rew6vAynM+dsVI
No1T483vjH/TN6qZDwQxN4OKt8wGjGLx2Lp0PRWssoOPlRGN1pcGx/TvfYnZVfzl
tsPHvnOR9JE7kc0OSKLpsd72nnUVnsOpYy6VQFCOjxHxNllgW8ZJ1nNBR0QlxC5G
v+3bF5CFgIIX6z6+HHESw+0FqLu2P9YPY7q6maSk0c1ecSfbG/VJTUIBUXKzR5j0
JZ5wpE0Xil1pEfCUE9FvB9LsNmLwjqey/30Pi35WYEX1lAyJbg9TygjFEgXA40Q5
F0qmTthkY0xJm7NEKkUEZ/H32gpXq4MyW31HTsQQaJYZOeIhrrZ027LCAGWNeoXt
zLGK9zysbRqUfvS/9cRpeM4ePSjR11uIZvn/H4TEB7pE+tY3rq7yAcm4+vMFORJ7
RBoq+z2j0RB4fhUnITJWBPUTBVnUyZlD5vRf5FYtfk4hmwR0bw6CJBLe8+A30Bdi
fN33BUy73lbBzDPTjANDbx/vHO8ZMdTe2fLneP0yNWtxJB4tUOS8EsDmo6fV5WZg
7FJ1f930xTWIpoNi1D/03UJAAHXNDdbjkIBn6s2bkVXsz+D0BF3ST1RUKmCw6+CN
E4R2SufsDgtn6HMuFdkZJ6aj6hCACTwKKniw7pxL8xDb0D+Db9RumVA7CAx2+dMW
fvYw140PzIN20UC3f7kIW0DgqKgN2vnjDfDHlhcLQ/ufXpPQbYTeNdKnbFlh6l4l
0+L8N39Gl4W4+U815J75LwT3tXjh2lxkeFDOLXmmLkNav98fjbdPeUShJegyrDd2
JW90T9vnO5HDW/vnoCQCxTOllSYPckQlhoHSrDVYrZamnOp1+DgTk2uD1qHvD6rD
+iliYzQPEKZnKTc9e5K+g2Wp3N3q69hWWwaDcPiNViWF2Ie+feQBvrHO9h88taTv
+wWGRG1VjGR+Z1OGYgE6yHyooFkjl67M86k8iO1dxwMz2NkLIwP5DwUV2rEq9o1x
WlrkBDgQibqYd21R8tcdJvhmLNpEX9/fMYs5KkNGHZPtEQnuDd6YPPWlr34Jg0h9
QLsl/H0hsfeHUPb+7AaYFFO8ymIjrT5EzzlD3NOFnHUq0jvREKQZp7FgBMV/Mbjt
UR6PyfaYyXvUJsHKODA3iHJg0vzeFz+IiAaCQMCFwDL1Pr8q5XP6Y077oJNqadaw
GfIbDkLSuw8zG2LEkgottoUR9PpJRxO0emMNSxgbxYYUMnwTcQnyiaBKoVGqB3nl
P+6Jf67whGT8f/MF7HJS9WUwfMJQNSEMzZq/Gyv0FgwdGtGc+OsomYEv4QR27eJ0
9VXMQe1qPbyvOTDN/nyZGThChWuBB4a3nhkHYQViSyaTB4KagxS+Za5Oe/alXNhj
AGE2PiGBmIpRL6G/dFlJjtwxPNhzyjFGDSZICaK3BKYYIknX9GYQGlRMHsT5IHvK
GRpGh2z39zfni3nsmougBDhkNO2IhRqDPTavDlpYI0nvQfTwMlOHUbKgW247aBWX
/uW51XkgIwpPB1Ciparug4a3yM1gDc40b+n9bq2/Qh2lIEkhOATV/E5CqJ0DSJBw
tAiBpPMQoYpCaBk3aTb4v0vHpqw+ZnuN7P8UktpHDgWcKeBCdw5tB3a4UCrRPLGf
4wFN/K8i/4eGiGdXZhCHPRa1lCsYU3Dy25xo46MMlla1aBWFbUvklF+LQy5KVoqP
KPYsk7dhLZ6Vz5sPz2N91LUgZQNNvgSrTnKRPxH4/J9OWeli7s59+Fr8ZDeYM2C4
NOg50DD+dzRLp4eTz/Ph2u95YQ6VfEep8u5bvypVBQCv/05KScweOBbEfIO9xH1y
R+2dftKCKV7d8dWu/yTZCK1/H7k3WK6+1aRQD5qGVr91XGWpNPymZPGOE10xiHh9
I/GR4sEPbsfBPOofBV6pnnKakAGDHf63JgYznbhGoPvBrDREzCL9iV2H9kRIuHLG
n7oMU5UxJqwaMpQFYIlAAvk99zA5SaOrjEgPF627/GHOcuGqor/Lpg8iKuCE9bT3
US09PQDbsbFn33UTCWYlVKe1KZNivxNaAuJ2q5orn31+reXhFyyEUegZtjh4FybA
d3vMvqam8HgO8Xpf24/kJDQ1ekkEwrcvPlAvNTiA3H7sgmnwNNlzWTKFGdzWyjvl
Ncw7kBbPqrP7qPOF1gt2vBpSwOKBfqVflRJcncdiE8slb6aX4PZsQ032ksQLVkI5
WV4L0okdInt06siu2wwwVix/upJ3NUEUJVUc9669xAdmdlCFEq6fGievG8uqBLBR
VtY7xCNBeKTr4LKiUqkPJzEXtRP6pL/9evn62yWm7ovidtY2ygjTPDhF3ugWlv7O
9hV57/qjhBo5BaMfckQbasOL64krGeDTpuxSoOTGSkoFqwiU0VXPbuJD8IQyQ2nd
Gs1aw8HB6nHNiOJK6PuIVA71Nr3VC7MD/gjizc629M4kGMe/TBH0nde3iKB85pvd
z1Ij6fLqxxZIpYZNmIQNm8Qi5cEq898pihf3jG6yTuqDGjDOPqj74NA1KWbBuF2U
xH1JbdayVnYU4cGdGidXW5HwCPEXWWaVJFcjkExrfVWScBwrr6Cs5vZiE5Zm9df6
uJ/YYMCxNkJF4Z7uDUdtHaxmGqiayMJx3LU8lesk/rEiSD0/tP2lA+Nh9z8X+v6F
VgI23g+NWWojCSBKVlrMbRJCeahQO4auO47TTRAsfuXilw/eJZXhX6b8ShwqEfOv
tcHi7XE/lX8gEyaH04IUzQDpp+gcRXsXEOhjgxEQZdTCfy8plPAtckIPf8ZPWOiR
zfyhj12LKOPnoggpNimSc5dMDazgxrUw0qYDNQdIpKi8JHbhs2Ki4KyXUFvdeAWq
8/z+0XDOyZ5OgfM8Cptz3F6WS3KjO/10F06ooMhBRjyx6f07SGZ8LF04cNm0300/
WPYkUVmEMFkF2GDPHHfUkdCec5k8gKf0mQI6K3Dqu0ImRB61pM5p4Ed/3/y0nuV1
qzK9X1jq+76g3wSW050tDG6SDK4tlqob3JzFbTDIjQnOz3Ywge0oghBz18mrzLRW
Aad5c7/F3XLwbRjcJchxLE5983GwYz2bz09akvykM3yNUKc1CDdorYg5vb8eoMPz
4TNv9MThrSufTZXNGSCv+sHMVuYUD0QImojShridUqdBklMgDWUX6TTNQZy/qUn8
Wj7q9t3julFS3f5L3zwu6wOi6dIW3FcDYatObpSKQ2tFYQXVrvztRfF+tyNG3Lyh
jpeR7jLqcSBRCA/abhvpYuur9jULOgUMjiRO2aHfPu0Qgpen48rISKi8EeQSbR4j
Waaxo6KiNaU6vQ2Y287s7SCYnH+VpJU3VGr7SVkuuxeMIiBaWw8lOg56wcRsSjb/
LgQF6ns6e7b6/cFoRKGx+a9La/s0rd1VqJRo9lt/zizMqI+KRSlvm61nlyBbm8Xb
huEzAf8GgMufX7jw1dzKGqeyY+d3d0vvJZ14C8dmYE01pAedcmmO8OgUvC+91E67
EOqpjr6/KIS/qExESwWjJnqClgW1ws0Y6XScdE4DGE5fwkyUgSfLQ6RXDik/SbKy
rzI/dPW6WmSCpGPkie0VgjYNMRVUh/QGfQWczoZwlT6s6QoPoMAoKGWiW+kzzzfc
cXDIl3FO2SNjLO3PClVZxGLoNHnKgpgr62QeFPzfnsHs8NlFc8g+PZCKWpQuMlyy
2CACS+HbJCQEQr2yTcRoZ54rsUgqOHYT1Sf4FCWQ6T6jSMosdebe9uXxxW5shV5v
zDdrpzl/umKc4/snB2vSYz3tgrP3i0jVx4KBu1OP0ogmjapZLR9H0SZigNbjaoP4
Ou+OtPhaQuai8pHEnPutsYQIhw7PyAvgDc745QefO+a7f8ozfT/EdQiHfltgmGFr
BU+cREAFBIBjxWwSNPNQK0b2CZsKfwT3Zw+mQDmuZHvi6/3g2f7P2DbhUIQijOkH
926+G2tsVRhyM29CpmsIvHnAN7bEM0KrBxfs3w+FkJhg+UOW92+xbmnRSqh+eqNZ
W/8MA+m4J5SSmX66JKkcnsbRAZsvq/RvV040BT+eh+wFhshdZxHzXnCVAhkn6XaU
j7jgBLETJfYXcYE5Mb0Kuxi2LuMArRiLfFGbe8TfwACyRJ5Dv1V+lJ6DF+ZnTStX
2BR52LmvewD66qVFMcMHmSoKL7DECJT6jllgpA6fEtPt9LLiw700tK/KSQm+sXku
DfUwhEjl3qM9eI8qBc0VRqCekGJ0H6jvRfTVDThI+9TwW/ryKM7kiUzzb9IacTwR
G3/NXIEwbDTIh9BwlXrTvSfqb0FMDJLvJc2l2aaEr8o2AExVPCHEHT8hXqxHjOH6
O2V2W/P6F83lEuR8g/OKEBRyMdbhB6XiwX9AYh9ZW3YDMSzo35gyJriBneokSDNg
5td2C6DPirNAEMQwizNxnW1/c4jQn53BHTHEC6oj/WR5Pdxbp5zLUaUJDHwYQNO7
Gy86Xm16HC2VIFWt1gLv0MJI2cTmDNdhXnByUremxUeB1hn4aiCGQYZ2cwGh2tJI
5bHy8kV+0uuUPCrFxOE8ifccrNc97oXxDkHVRwlpuTh31/SPNcvPy4rFQmmPlP8s
fSNUJB3lQ5e0goQInWRQFyncEW1GgalEFipg82gq9yq2ec8Mktz0C5UpYPkJSDkB
ANktqM4LM+Ivfx2YV2/HZSPoyoTphPriHN5Js978uG4vawV17s5cMjCtE+EtOKJn
PpMQhMzZ7dGNSRdiMmXeibjiT/EmdgBm3/qch9lGzYv4gQXB4GpltcBBJERwePg/
D5/CrhRRVa5c9fI5WpE2KailX+LcSWUDja444GM0PUYUbhVB2SJZ2HAfAi6C95Ym
TB4Z0p7ObaO+Pq8YZq1+aIcDEEo214tbwlZoeCmP/2PFsMV7Lkcf09mTS75mglYa
hXEHVTzPly3rwFzKIUzp84vFO6UdcsDdQ5O/28pNESWWhmcHHl85uZ32ouNZXN7x
cTslSbwQe21/rGHDhUykaX0ps6b5fmgK+YtruagCz8HM3D7yj3u/4ZNSdR3WnMX0
Ds5WxkTcS02B7Y005rU84A+x1pW1yutq/SpI9hlBdpEP2o3tEHMutWQFYr0FLTsj
LqI2Yo+Pjbur9T3+h6ZKL/qPqTI2qQn6a0Qywtc8xHpkOsWs9abDD/9riETaAc8E
B/DLYMtQYJdApaCq3NJHsd0hd1wv8UtqE5ljxjadk6clRc3ueW8JelQhULFjcGOA
M48VHybRuJBb06ZsNkVxXkJk0i2eyZgQb7KPpL8zEEOPKyvXPf04XA5n89r/bWzW
rgUS0j0G6emj5tgK9GRXM35scPfM17ISgcrT2ap0dswFBvhUilr6JEC99GNJzfoD
jXh6YSJf3Yv0L/+A4v0qoGaynYfyOknOKIq1VY4O0qx12DhApVd8OPI5JiOPxs2a
pveQVcjDO4Z+suWlscloc2OTKYbXNlHz0FOhtfMzNP4Ok3ntH6HjLtdusH3f7AQo
SVgp+1km9ZQE/oDk/gsi+cERfKtqbFLkr/eFSBK6ScMldlSsjzct9rCWj37IBN/B
M6oKjG8xpyN7Z2yDow2eX4VIWSSJ/SNRniIhSMB0b5s11dZP+We/sSct06dtjTCi
FXphP4D2FgRZzLwlA/R4TIKxFq9gdhEZoBWklMRbqTsRmOtmjo+nXwPp86NTpBXB
o66Z1GrmsE7S2AsTVwUVMjI/10dihPmwx6zLbAbsRypXaaWQRUIUh5xEAwobZhaJ
8dRWO1qZKPEtxeWXOdmOI+1NOznImUHOxOImbKW3Msvu3U6IjPav9mJDPqHT0n4F
6biDY4xEuUZ8ykGl6Eh3eWr6awB5XOKceSGDkAdsbLZeW7I+pv563BXh3+Uc0m4y
OiMD1zDkFgs4AMvfYtoyj1XiOA2TwuSEJ2ZhRYKFyps1nge+VLwG2hPFD2HWygJA
C/N3g9D67jWRLzPHtpBlzGnx3ebHFGr09jlrPcFx290lYXChbFFUQWKJv3l0ZAV4
hn49DY+JZPUmwViy91K2BVWWN0xTnO+ULyYllmtmYOBx0t+2+YqNqRZd64Fz3SM4
ZrSAqkhu8bA2cW5jJE/N0+ZxVfKNrtvGxNT+Jwmoa96Uy+VBrwrhWB9LCeVlhq8/
eThuC+ov2TjnHN1N1SOTlK4X18895YKAJ2xHUeWihGnjal1c8NtoC67Up1E1TQxi
mJOddKUKckpsuOo5kLd1w42hiX+Mt8lSX+IqYzXs5aTyJ7sq5trUT1BF66412y+x
81mKDspCXQhvmscBqjMMTS8lZPwmMHesy1k+eoImzkYEs4k8d40cRYnNEra7moLy
bm28Dgc2DwZTP2WBzeEr7Hc1vRaI+cXl75SxJsRfCXEgiWmWr7eDEbBV4BjFYOwI
4Hh0vJfOhIiUiLX0OsyNprYnQ769Ruc1zqdYw/i5g4uYMXkNJvOn/yL/ISs+iMPn
YSNHjZie24k1V7gyz2P9Yuwy7cGH4FxZkLrSX4UnKM+XHX13snK3j6vXMD2vfb6j
dQhZWKiX/p9dh3kZY+53Ct389pssdiyI2K10w02JZ2v3bQJXVeTA2K8K3jI3hNz7
ZLY4m+YT1n6dtzFjg5SYHcscVCkNmym+zWShPkvpB2plbGAhhjOsb4oOFWS2ryg2
04qxFd3p2rWWiPE72tlM6Pcdv7DGvQRxCoY7nrde2i0xevqKuH7ELe/qR0uaxFK+
N/o6hMxcMP+b9BcjgOf+Ub6aPBa23ELPRpsYgwLnUKbbLVPvC/beHokmqU19kpRv
03/uvGIrpUwXkcmCwICGroNSwXlWKAEQvD5xo3ngH5FhJT/SuosAox0gEC2GFI9+
/kRUjUiH/TwaxLh0mgB4jA/pxPUkZnL0+kowusoK+BENaQct+CT8dwgJ0dXThyAO
aVJpxGwIxzPFwyrTjDVvrbZsKFRQWJLHC646bRBSL15KwjSZNkGg/CNeiB15CsYl
uzhuUzqkKAcno3qYP3Vd5lJc46ev2+2FXyK2UJ4Oiu70Wck5ghck0lkIS+fM/2K3
SFXX6Pv/EYe75wFrdiERaBuglC0Q4epND+AGsa4SdRnYK1tahiGNawR6iah47RdY
lMH3DPmyiPy1PtSuwVfFiXpdR1iei9ZOnQMVJtGcN5PVG7ngY10WMbSl53zz//xF
ChsfxVgOn8N/LpDC6yVk5mhT18kGsLB+AKyGx2SOu77iYk1Jb8hp1+vywH1yW4rZ
dc2i6e4iNtphqkVUdOICs0/k0qCbENU304jwOfj+90Ap5TmHQNNrKDLYgTp700s1
OxFLTZ19Sj5TssG7bmjBU0/e3jTiw7TE/HrJxPdRJvqZjl+dh0VbPUnxXBbO0+JL
cIvh4nVUnm22u9F3hzkW2ttY7g7+n24+GuZwDKKk2r+4wlSqeO5cbcX6WPHocLQO
OWllxVINOJJCvUMrLMYNECjL9qVeIO5Gh4vNOh/dnwp0dcIVr9EPNtWOmbfhjsbd
kMg47tMcaLT9LiH2I9IJbQT+4YhiOsryiyuqAuBAp4XF3JkgCrvKD0/Rk4+8iZeg
uD7g/wnW9cX1cDM+TpO04oOY4Dve0G2g2R3mvUvfMnzcHjkNr6EdkZpKtqB6/hQG
Befr7vCEs5cH80nCknf9siQ2T2NkCbIbMxE15zCcoFvkjLFPGDRCr2QE8iABZk+P
un3jPI1/lCFbJPkJMeWOAu2vW5e9P+Qe36ZWI4ivvtlyNLb/IQu0VcNhwAA95IuC
BzQNz2VbF4eYTirkP0ATajstX20wHq4ArfeN5mVJh8TBddzuZXa40YW2aSNid+rW
xVcB+pw+u1ozNgYQfU820oT1HvaCQeWy9rwzeiKrJFgQapXOJ1BJNSaQp366kI4S
1EqVJHgWqNf9rPeo4+s/yq9PWRGLbqfsFTrRrOm2D4VI3FTNweMp2vXaDZ4D1hxv
uTBgM/D0/UNkN9QklsPXshsmFMb5UYM49IYo3PvNqVIwicQ0ebjFxDBzB21LSafX
XvWctEonJs6wXpd255xAnPiEH7XiuFoIDhwli0K0z1ojoJiHkANd6A5xxvmZ1eFC
z4xW2qG5UP6ncB2LzO9t16vXEox7ldbue7X00CDXt+XovlWjUDfjZ78JoxcVZkXU
5C3Yk3AYRqeoIMfhKwSF9EOn8DOdAV+rLG99yzNCwJvWmF49U/hmNtYNaaGKXOj8
6shJ4P3L78JbvN4ZgCJHlY/Yr571T9Ke8Rw5z5KXeCtn1XTVXlJE4dbwSJpcohCp
vEd+TPgGeBcvsZiy7YrYV7d+PlCqO1NjcDkOf7dgCZnaPcrES1UyZxi95FhkKhN6
hIrXZZ/j0oAOtGlMG28FMWnbIFzgsR1gADbDT8bwgoEp2sRPO5csG4Rx9gAQs3SH
OPEJ0L22bEXekQqyozuwkVht2UZlktoxpzo+VYjdganreppBj+UjFQgFHBwLxGJL
26xxgiXzI4aeMEGjkWPDDvpJATeeUcOHkhwbX+CQPGwwRvtuC+qBp8UoBqEBBtZd
0+EpF8P+hQ42TbPM96FFQHvPJzS0AXYnPhYpn4piDT99/631dOCk0/NCtiD/kQUB
KkmZ1jS+oGEEmtzK5czZguAgi+DqtfXTAKNnaLlk8lGXpwCflX94Gx5X9thEPL/n
IQEseXGt0a5Pc1WhCUtmKuC9w9yqI+MgrIp0HA8Otv2hSon+6JZRDA8kWKIIhvq/
zCETfRqiFyBBs0DDGIbWQowTNhsUnKIZgYNOAPODtTz7qX2QrsffdIuKpq84nJKI
jm/elZXGmbP7XFFa3oZf5VSlMwpG2NmAMllCp7H9gwn/3JwgoT2eD7Ggi5cfzNQZ
i3t4VQv7yufOr6eDY/g4MGhXevCPebxJp1rxeML5QFm2+lrOAMq5mg3r035GNkkE
KiNFgEPBH2i0qAeMjAdezb0ugdfQXTQpR/fa4Wi8I+CYKwVFRiqZKaNNo0GnjJ03
CYSsdnlj881H2vlxDfCKjCKAu3K7lv3iB21V4t5INC4fA+qKR/X7VMxQO9WZ0the
DBSbgESZkxKkElaz3GqYL9m2m14qHlC7J9F5T/RJttrA3iBBeY/PwZkGpop645f3
uiczqFnz3CIRcqTH4aPG3dx9XOTC4bOEbK+k2JzKihc2REWxcXphVBoFzLa/RluT
qNP9HEM7YUQ/gOydXOcVVz28LV0HQB1R9AKvHFbk+0Rnlut2wkuKvcKv7v3mP9Fw
/dRyTuWn1jyNcomekmM1VkSfeSDlah0hAUaBWw2Jm/VstmmPD4EZWq+c7DXcvHDv
MnaSyHNlcrfctT6Ij/jsop3nyUBZRnewe5jRa2DKXKjsX5lB3IKhexSbV3q35JaY
MoChQ7GjDtq3InWkrF/6mssRl9q6ESuhcMswEQlYq5b+4TRUQdv86phI664mIn6V
lDaRDzfOYsjyuAzx6zRK0DLEeMJjxvlyz412PchIEREjlkgfW60G4+ZmBNaUeIYt
Ow4nJOyXPb5Yd4/M7DBnt1YSaorxOkPDNdY6obukjKLGItl1JAuSjmNBrxqeFQnZ
eLsnRUhCkz5SxTRM4Bu1Jtva4Qiw8QKW9Y+5yqpe7fxUgUfThu7Yg8OmTBf6cwmn
iYYE9UMLdAk0sNt62QHpsSHX4WEw9R+V0L85jwuFX8j66E5UVcoQedsjEZrJEnHI
tfJYfJmeQxa0QvZ45ZqJdNwHbweJQgV8ZeMRpHMGbGI2vbFIzgLkLcMDJRm4uIct
7u3lDLEsyKTvwNfnOkm0cZJi/l9/toYULmN+O11wZtxL0BVo/QJhBR+W66FJp2nF
jrmHW9AYqBpHMfO7ETuUbP3mbkZNKu3tnoDeo5M03QQvVztOlNWbCO6QzKO3gs/u
UBQZdExlU+6qVz14PqYGcwk+gdJt/2vV76Q2JEiOKcuxnIqhxINkQAWI39m1e+dJ
Q90tYMtwRo1y+nbfqkwBhYHFRg5ylVb5bUPb0nryrnSU5+GvuW5WNX/mXED7l56r
TOaYRMFPwIX9ENxXOKbexdm+80gznWDYJ+Qx/RvPp/i0SD9XAGmdXlZmmgDgKMhr
PrFzE3GPP4929dlo8wj+P/y0FN3/wzLk6if8PNyzgubJzZwpe1HxCsAH/m4mBnNP
JCBpkCUp5W/8rkkFOQE4BaXK/wUJBFud2hT2YxKuZ9dmphf93xIZrf1koOQ6sqTG
dsb/a7fbMmLWYHs1Rz1cZDDykr1xRKB9od1WoNmeo/c1PsR5Y41/bEMkgGcX55BQ
NUrN9CXWtcW/NpMn0ao1EvnYd6jgiheZOYRoXJHiqTZZC6W81xQMMeAamFssV2cO
yM5bxX6Mo1w5U8udocfgZw+xQh8GWd5n25AdGAS03qt3svH3pfSyrz8qvBE99LMP
RvFW9fQrTBWGZpajxmDRX4rvgu4aI42+F8DkueWrnC2KkpsIIyEYDJpnpduLJ74D
iz1gHiev483w/BrVZ1WKgne2X+lsTsLBbZmBjtt7HR84QDv0tJia5aCZpGhl/k+5
cbD7gjB9RATU3pFrJQHh9TF1Gwxb5U4pQ07qz9ztUBsy7RZ+jPTtPVOhSuAktnCX
TizuPPnep3SuDPp/Ebk3pxvYN10by7nQfmehHr8izLEhFiZL/hyzJLiMUkvy4tTn
aQjGmxYNHP1KYcODxBjBXmDYPa3w1700EyI2JHLrxId3oBhdsnR/0l/PqIZhuWRW
l8KQ4Mxy6iMGILB3lVrMaDIYCy5MYlNEWkhxLXYf6+hcBLEMSQfQLC22UXgmod3A
GbWOocXNASWsizX4AYtdHc9DM8deyBbeNXG12LJOd1Pln7hwQPFrQc2V+3JnPGUe
ipVWoZD1ZG5w1rgvO54jgM37zSnlEa4/AZvhcg9lREgjTqJyLynvYPw0IqFD29YK
l5psTsr+C1QAbvKKJe2vD7dJuxbrT/1siV0eX8AMK/gEdgCfWO38aa+z2yJFsBXn
zMcvR5NcdCmAOR7L2478Fin+dqX+bFVx+8ki4bLi7BIVHMevXO1iTsUUHtpjqE3t
zpY3ZVd9uJiEHeXgY5YNTedpexFM1Pmv2mjORW8ptJjDXKoBxJwCIGf9mkITOnLk
MjkDVL4ssNK1RT3Poe5b+a3eDtlTZ43kdjbfUZ2tO6njiGY1sE5qAKEpru2cFZ02
HIMGmPNY3kHqbDA3pcGZpa7S2Nkz/7tRrPnPsCOp7LpJnGfXUCZRzus/1Q21Q2d/
jQiU7FEN/tDhdiQI80eg+VvWMvvBiQmo9PQjyh6+4EkqFi0Ab5OvgNOhS3Bogemg
V0unKrK7q0zUIlH3xEJ6FflsZCz3UzZQgPvVfpAFK48MjZKCy53dFxkEOBpGGSQy
a24A+fM2GI+5xwJTNCD8lDPL0uDXhcWUQtzHxeq+6q/pX4K2fMKjmirNv1zCiCrU
2OvONDl1lpUqAUdyDHhmjx5GynzZSh+Dvyis2oQJJW4vBDCOpMa6jCr9ltawZqdL
2HkGCufF3CBFksicc2aFW5X9BEQdUkxUaogztEjXOaHHKLXi+lmfDFzZB3ocx8Dd
Wb5zq/2cQnRzUEFL29L53C3DH7z+Nldx+6LgZ5IfCIVSgr/Nv51VQHrrZmZaI3rO
unNvA2ffQNUoN9rhGbmEocg/lH9Q2YjiwhCZm6siGOt2vYncsXNkNtk6IY5/Fr1D
NJ3sOfa+rVzk3UIBp8qCjGSNXGUTuUOkOK9l5L6oyCwvc1Z6lFogvngQksc+9h/b
xclFb2yKXgUqi9+Sylsx/rWeI47X8j6+TOSIJJVeT3jheUams1qSk+DEsk63WCKk
7/p0PblwVEmQ9/s3YdWnHblH62VrpSp5vVXBN/yPgPbYc39ZANi6P4QV4akVSUve
ODyPAFBUUpShN4fgQMwkTJdfZioQ2RKuP7/SvSFVLjFvc80B7UJvgad4iu0r6Rx6
6SgxH9xPr0Zjlai1KeJs9wGl/0Jya/y/sRGaMTMfuYyw58zfFfKoq8fJGv4HsU6V
XstjpWg1xJqC+L4S41JQexOcH9BhPU0KvDJ1dgGkfhCj0NnElnVfiajED+7Vx0Ej
T75got0I3T476X6QGG4m0AkutdR89Xw4q1iE5nCE4DfocTovdrPjndpFEw285vyv
ALYBymN4yVGUkZ+7jFL7NHK0wzQnhNdx6YF9jwUiCJFZlhivWGpSBtIYu9pQmkt+
pdBw84/CXKzGKf0shW5Yr/JRyQtdnX/wtQoysMaVg/Lw/gpn57wVYuNaia3T0IUQ
sm7YO+tZkLge9Z5sNP1tV5Z3XexbhTssx8Wcn/MA8/QwqXvwgQP6b1xbNN/5+3hz
AqLO2TLvkAN+IORhz9VAIinYZhoId8MQmweenyhcoqv20OWeDwuE9Ll/VQUj5Ww2
DmYeACd+s67yoqkknvzaDpsKGK75k7PqPKGS+p2f/+MRImdvhmlmrSeO62qfjeyl
6cPhX3nDAgzdMtUHtK/pvBFX68y+6Od6maqYyxUdZ87UMs3VjsaqxleiNxzyQOYz
Qige6+3Xx4zGV8jJWmVVSFzQMuOdIax1fplms8Je8A9wESBAF/vEfLxWYzoEyrPl
fGzoO4gdX/F/vWY7dK+Os7Cf/YFwcP0PevAK+O8RjVFYV1/96JNwOqdV7x1HF8Rp
bdWk6Dm9WSMeYpLLWy6T+oujT5LJ4FSH6nt8y04yGAdmIVg4Tv63v1ePdSxuZq6k
Nbkot9HKSo4MoOI/xZzXCYcRUG/1dQN2BH5mQEZciyo5wbPMI8TZwCPBocfssg5u
zEsjm9mVYffggoFn4g37rssuz8ZmeCCEI1y4A6wERuDhaAa+4R9k9aqiqbWK96dS
sE8gmcjZqBHRPAn32UDTFFr8A1hlnlzvIw7HWCjRaxeK7CAbHiLpxz4LxqqaRdkE
vCNZX8S0w5yWsaOa0jkpGFhRkYcMpjHtCe1mPdOxOQtizFSD99AJWNDGb3ozD+9B
N3VXvULUFcdoHDYjHwAo+a5gQr0eNS2q5RQSp6SUB3WINg1nBGT3bLdRnWkJ+Qcn
M9DqMiLtP/fHtPkwhet2B56VAyrRD4zrOyZUmYU8rRXQgV2VDdC86TMQKxCb40xL
Rt7b22I9KmN4GcqepGIYJypSkwlI64ycjCQ7yVEJeZIz4XK9Mxo8+7bjAI0ORtci
MRldinq4LtpZJp6vhc5hdVcQD80TYelbquZgo9gEUrRw0ktYtT4NwXtZ/qc5/k0F
tqTA1RLpohjeqttd7mR9zh8pI6tSrEwjn6phowogiOclL5Np8ur0HBjp3nc9qDHr
7kmcNIqsBy48pS5XKHT/m/AnAWGnW75kTfOoqSZtbex1X43le3hloK7WIePakLf/
t5JKXel56ydwx3MKD2R25KIzeRIIzID1yEAS30x6LgWwS8jg9CLcqMko6Skl6DCb
ySw9h9ALnhR1PwJjTWmbTfx3AxnUmZU6K/ldsG8ZX/bWhdKy14sVXqcxAh9QIh75
wZ4oQc+y0f+dvDNeOMcJ88/PzsseJBzCH4HLXNAI4bl8rlhLNSEJcnkpXLQIG0St
jHbuRDGMW1nEAQXmZdoxUD8Hg/o0afVgre9W7261ihoYMKIrJoGUsbKCerXQmN4T
bTQRnX5y1k+QGZ8H+xqEehKugk44b1Bz5HxWhRcYbdNgYTbWXfzzeIvB8byF4xfw
mKBf0ovdrTXoSE/AIaOBQHasjKBmZYCECqNeWX/mxQ9tywh2zxDS/5j07hTC71qZ
0fzrVBctoQpLGYtVESSId0scgD94R5Z73xt13t/cCI8kJhvl/lgeSxPV/4d9F1sq
FEbowrej2ojtcTjNSt/Ob0deqma57C2S2vPHwgKB+GOg0Y78oTgFUcQoH772Luhr
JuTeZgHPPeb1EuriyNTiH2bumwOBnJJWMph4ukwW5hFYa/SabAxJYeeP3mNP9wk0
HED5C302rZD7b5uxt/ioMzvGeUbXhONjTkJwVdlXiuoblVUL4xm3IPk7qvd9S8hz
Jh3MPi6DUXvotzcq47h4y9WFtgB8RKIcVfpWKxgGncRhD+tSTeRtWKY5aOHquFWk
tXV9Bupd5Ntzcit1QHA9eBANiGGjf+Ev1QalJ/H1+D9kvRwTZUxn3zAx8wwYfujH
dMcI3CUUvdZRVwlnhKXGtQ02TI+ityVn/kBkVRorCJ4FkyGOCFQJsO6quOo+vpXn
Nv67trLr+iYeRUxdIIAP3vHwZ3WCrw81tRKrApohghzYzqrpz1tethLuPM91DNDG
bs4zWbPegM3ARubxIPR3EaDZXXDNFbNILsL8GNJ1ZCcI758yncMHpFQbbl1jesNt
fryf1SRaPmZNVePANluuZL2zAabH8v1A5AG2g2bdbimJjPQVQ0GHZj7txczfomyc
0k0GiHuRJv/gOwR5yZQeddozaCajfAcApdWEr4N1+KaZBsbnu+UTyJMUFV1t0ffh
Vp/77cYoIWf5vlty5G1ZNaYEUgzEHIHSgutK/hJzHAnnv15LjGxxvHFYkDMR9mfl
oETDXRNG5Q9c+ELlXsRBVp2vpCIrvSC/qvJGOJ9VjHPiPI5GnWhRWkFcsqV/MIU7
26uur+lB3VLSOjKkZSdxMpRNh8/tbW3k+d3hMmrRXMR5AxQZuWGPofGYqhHEtmVZ
v7A1vZ3xOiF+NmvXpiTmqOGTlYvFJ3xE1+G8kG2ptCySqishiDbipuG/s5Rih1xc
PyjtkHzXmzX8ZX6TzrYoKNzZQPfFcdsAyoLv9tn1N/b22ElGCkAYLvqR1s33BRT+
eFqNMfU5edY3Iq3XIVj+dJ1wa8QlyoaFPbLz9R4IG6RjBwSh0uKV24c8H3iYb860
Hj3o1zAZUUUttt7wtfVGTLJUm6thJGS3YTgOFbN+todAEVLxzZtjjdfCc0VXFmvH
pOpFiRIpBq++NUIILHQhpv1HZ78iQP7ADpTrJ77/6FD2/FBe3tM18wl5MrRW7Geu
EEMf+ZEkuV3QUim9ppwGMgCY+eyNsm0+Q9GTCTHzPyABSYFMTXiePY3fAOxAhWCG
MCzYftIrfx1C3s48NyT7kNmnKazdJ/PEUPOl5GfLDU87FEQu9GS3nRsvuidIaM29
zPtaUTPxhkGxcpaO2RZgq1C0dH6CGPXzTcY57PV/kS4qkWvgYV9DDdLlBaiVtY2V
UpjOV4AHFr/lOkyvO0Ko/h2a83OXwF4KbBusVMdSfyEgXz3CkqsUzXTMCEDryB1l
trH3YCbeH67MQOE6s+sJAFWxxIwo3f6Ubl9SuQX35gj5v4mJQr/LPSC+jY4mJTwe
ZUg3QTf9CwOZOsbedh3ACdlsvEx89Ea4+3EojEizI4p3gP9V9CUGfpcErjbQX94f
tN38Kst+pbumsnxcgYnCHEI5TREfAfLrQ/IN9SKaM3sG0ulwgNBYMnKvqlECycYI
DAdIVpYGzt+7Ndju/e2v8INzFT1pKTyb0emYXNB7xcra+J9bPi7H7QtBMaRHiAP9
dbY6x9tVuCTZrm2mmXgKi/7FvxhEfbmOuZYXy03QxS4aBh58pq5b91POSMGXZXD/
+jeeg4prbS9FhDKigJqD66joMx4tBaUqA2fHOI76QAc98igcSayouWLaUhNeFpa9
3k+xiFJByYXvlGRNOYRxNvBUEfNwZKmYJrMq0CLIh69irOAwiziO5JRqRIXQjjbY
RaQQ6hMm/Fs/f1AA/vfxZhYY4gvlmx5PiUSEhP5OpB1W2eIUAMk/EH1iH0l+e42K
RoOj7X5dI+vtMLH2DreudXjITN6fYqQF6v3CVw33X5zwZdGT/vpuT5Ovmq+owBdU
o15Cfi9tEveG0vosMqzPZ96T5PPy+0O9MjZieuhc1XtYq7RLBv12AmjpPV8a/oeA
XYLBbYnqoxDLNaBngCFX0ix2hujokjJglsCtAVaVC16Nmg1wNQdY2z0NgWOW4PJI
uuJndON9ulzmQsJdgTH3gFJlw3ywacqqJnhV3SZ4LI1YBBQgNq48Obxn74iEXjGc
YQVZORTkNQNpNN7z31rmlkma+2Sujiq6Q0uUu66jgMS6OIerSh+DlkXGdyCySa2q
j1yrCkU4ZzqP8GtEelGPyB8mXdebXdk0Fg1//EqgnXGADR4mMih1+Jg88BMnCzO5
FscujbhjjHtqR2jiRyAKwz0ljCsKW4PdaHpPrvOcmObGbid7gnzORsy96h5yxx1L
N6hLSXlB5rN1a3YZPDIK5QpmMfdgEYVBbJ231lPyKZUu9ICGV0288sWcXKZPiJap
CVlOXLc2tSzmN1sdn7wrC+9qGQYgbiKtJU+tmREShzGvo8SSCdTPggTbDcd88cFW
4RysNTurBpqbrdqXF159Ap804EtzXdr/WuosajKj7VYBTVrC2AoE+1iOuSw11UoK
hcRX9d8UnMN8qim1PDCVuIYkvKbuLn8db/GYqvUa7ObMj/Icxtm2kx5I813GW7Hh
55A5k6MOH9DxfsCvWXlwQmsvpW9hGP8P3DaV2urcnehPaxMJ4K2uPCythj3ay0n6
QfI7lWA/ETDLykmgswmPO6iH8aNf1efCw9gURH2Oy+Js7WJ4V8hNmEQjLSzPUUh5
In3ib1CZJVVicXv46928w7KjYC8EQjvhEHriGNCE0/q5WbmZsocOyZpjnXEnog5T
wbuABQW93YoFt3HFDHNtA549/bACH0zo6uzRdwjEv/B45cBjBOA0otTCk4YSKqxs
9AyjUlgeGo3oWGA3yOzTjs87M6V+eiqhGCYGWEA0dMpvblN36u/LTqqwE5yT4z8Y
0LcreBBx+yo/BPpG+TJNStAPMA4Go7+uMlAb6Ss3/wusw0ytOkzJYWsOjxrmOpS7
zEhULpRyFnkNf6U2nEFfLjZwYtUe/BzM37ybykrNblCzXQpyc9CaIrALMx0j4gBJ
+90sRHAWNz1GrPOC462zt77uIbbMsuIuFONhDBukVDNbJYBV+0FcJQqLb+CmyPdF
xDx3hnAFXyg1bl7W0HvXjBhHrxRkYsfCghD8cQBcW25p+7Z+qBT7/fzMxejoxt37
LJdwtXo61BbQGa5uMJ4zgjEsn8JETpqkkovGBj3X92Q+tBT9hSz7nSPGYPrjHgUY
P/WNFPneTngSDAFaqxqTJLDLSdNSLYgHQdybXBMPYUaPmUxccBCTgRUC8w9B2w6n
KIXYhE6tdtR7NIqBTVzrz5KmD1KAee5L3/RSbAWIRMW413pWtKXdRSDnhIf98e6I
jrXVy2fn99GTJzohH333usoztNLPweOrxgatDIfaHQgyFYQemgeHCHFyE6qh2EqR
ewI4EvbloH17Rh1OiA3RXR4zN7xCnb+42GdX1tIbIO80oYNv8lWoOiTDL9TX06CP
qYcke/FgRYeM6bw7O9m51vONjqDKupS8vUumdfnC9IpPnd66URKuRyKLO1miVU4B
CvJXVtiWwUzk3/0tkFCZDeL0NbnWIAGDlj09D7LEGBawzlZpz4iADBASNaZh/VEc
Pr/uHZSmgbOjkuR/fjlxdttjWxa3M+5AbflEYSWPJ+Chfpsn+76Y1atcf6hwUAyG
2XVpVFCnuJmAdpui1eNYV2ySRuCaIMsTIvvZCvlBWjuAZql4t9XsM8DvcZESrClG
qEZGxRoNVg7ZaRG9W5xiDjKH6v/A+foID5T3CgQiDLbwdsumNb4Nl8MwVmu72aBO
MxKRIO9Jo8b2I/7J/ZqDf70mijXeZEgCnrqbwVoxRdXNatQAZGW7F9U4Oekq1c2O
1N3QGF6tZtdVKDrAEXKqvddEHUdsg6SdE67wcStpSu3o6v6bf/knye/7tPkzwBfr
1U92qdGVYToC0icKvaUrBcYNusnIopWaXu/TaDqzK43G7/PFxKRj/hWrFWOEV8Lr
VADOqzmXXjKyrmENIRTGh31L4CuBUoP95SniZ5hsuy75gU2v0nOsudiBohcy7sMC
Yiy7KRdSJ1eFavfihGTZKmMAY3H7UWMrn6z3PyqVUUHyxrkJ4ech2LnZ3dR2TKDJ
aSEHoT+UPBkchDAQvPUhDIarm2PXpUa6BVZzXFbaRvbA4dEbkDP4JF7oVQHriaDP
C3zuBi3GHAmWHUxUbRXlQX1DoqwnX4OGgwkekGKqh+/QA7drVZ8/rSMwr80KfETh
K/lCmqGehdB4eFFDYkEAQicm77TKmUz+XvyjGl8DMGEf1bo3BAfPvgnMjJQJBtCs
WH6gcBmqLR9pCATBR3zfUVn4U49nzIwMN+xIt0NX4iP7IAi1bdxzEI+REzfToxyl
qDaU0COR+fJBS7lB7HZEHmC/O06tHuJAqsLxfX/R59RY08MnFyb+yhJ1Da7gmHVc
t9B+6/SfEb60rIRIt9fi7ppDJxn1QHusPi03wLrH7uH452JNmo/qpxaKDph0rtGs
Rb/dB3OXI8h63qCzAzG3XQes42+skhJG17uacSw4ftf6XXMNZCe+5lCGETBBQPUo
d600H1VAvb+C8L2G3OGtbFF2nd643Dp/3ssOx58hPJKd0Etlc2AOmnHvQDWKnMKk
+Zej+dGZlnXxSnvo4LfOeOdXRVCBExJDp1K23f3Ky9nL+0IXFlxcVHezabOe1wLN
7UJxN9kdQePAP51tJCp8J5yMqRgIJsDK7gZPX5e+lAer1Q4N4irNUJvm9fHx9Jf/
VRohJQk+CLsPBrEyVZNNqKoHvOgkGRJdsSMF1U3EnKigUcbJxZKVmGhZe+FRQJo6
QKIhiJQW/R82INLAfsAUrCg074o9wvB5BWvSbWYEaoaj+NfbkvJ/UCy0uiFZVFoR
5cc5ILC0J1SGytn8TcpiBafsIecyzO7VT1EOZljw5/P/o1qdS/osTywqXHS7w2uB
rPkkETBrgcFmwuJUScoBcZCylCTTs6KekGyU34fn2jyM7Y4BTKll2lbbHGHQHH08
qa3zr9a+HSHcwbCVew+q6Sd8AiLZKJ4JEa+KIbrFdYjsv7noiyt8san++CDTjl29
81XhbvpdaBdyC6RZZAzzn/ekemp+/5pwi1CTHqqsC+Yq5ZBfQIXKQS/PJ983QeoI
tBSG7+CgKt7MNPj7U6dR1/ln6W8ERSqukc4B2wMV47XqHLYmBHr28qc0mz20cvwp
LE0pCiEmrvtMKYv+JNLNoACCoVoalZ0rxWKBE6a+uQes4cZwgCgWYWAKAqZmPSpF
dXC3kKrbhlNI0q62ihhuod1fbt9C+ucJepakZnKFohwUv0LFjTtZmpM5lnAUT1EX
JVYajMjCO9Ell3oO+5fCPIIc2FGfq80Wp2yLoR3QuIj3VrQf/ND0XHIIPUXPsC49
fBGlGphAYPQJTAcH5dpCUkuY3h211TloL/evrGhyHqFMDOdbRP0UnnfA/Jp7il9v
F1G1Q1eB+9FG+U5R3QBCEaHEGdCTzp+iXBjhOrCxEb8Np41MbqMlzEx/y3qlHDwM
rcXq9MQXE51bJ2LdlUd6ILG+n+8lb/0YVmn9Z/7nHkuWMOBWoEaFFLz3zv2QrC9w
MizGdH76ryj7F+KTwHjHh/vjtQsz+4tyJJidWQbVoDFOvL0KGvgx7KQQdYJ1SwuF
b68NcRhfp2o5sDjT6RenB8zVEdz62KqAIj4gEUJWaIkjRy3pq+GiE6AK/QetHsWt
P+90u591ZiwQo4OKBnUsFnnbtMJb2v3/LrnDXfAvDnVmIo/1bsKIknDGOnkTT9va
9wW/3ABu+vKqtyFGiQ1cP72HE1kgfxGlkwV/WWaEKd+LbTna1Ji8abZ/p+0ZSPxk
bARtSeS/rgYnMpT9Lk55F7qeRERqM1YGrm45ilhbAlKlLCzNtD0LmUsCwdVA1AmI
mvBEtbiO+ncinV/duTiid4gT7aIsn2QA1goo5tMk5EkJdCgDpuH5GrETkTiai9de
1XCNsYPZgDTtr0jG71vQzRSHUsoPJ9gedS05XihK68if4d0gIcsL5ud6Iq7MA/lH
caRMJ2k7tG3olBNt3/P+/xwlZNb/mQR+ylzQTEqMpqJ4aPivcCvlKhdJBnvYk1r4
8homLEfj4Ch2Th1K4jKaKYYJMWimGqxmkmAmRtq6J2iJVwty6aJVFIAbYOwydl8+
fw1o1GHHDEz8kfMTJeRpGMS1sFY+bPgH7VcleBZb+azS6F9XXZkOT8jPYci7lcS4
x6hf3cEmcELavPJQ9+YOjkUX9idXO0VSEbXkSzg5sJXHtvgtY9ppYuotExuN7W2Q
eRMJgidEfR0YQ5JW6uU11CuaWeRPnC01w8Nfgg3gUHJLV3M6MflkLp+arGjt8dX2
CHeX4lg8sICkCGwzGCwA3R2l5DR3Yr4NMWSWGWjjXHYCFwHhhO/GCj8l5xVAfz+B
8EB4X7wGEw5z04rA31tkEXBltdJRHU0XyqAxJWME5r5TCnGXGV7kkCUGMSu2DmTI
SUIDOYSensbe05nzxyVTFf4vqBatzmSd7rRHMB+yaEiyk5IE2d3eqr1Wdhp+Ru3Q
tgXxJWRGAZsfHAkPuEb6OCSVwzhZJ7o07ghtTipEcYZ+jYO2Z8JMCgMrzXr07a49
P1I+GPszls+OsuLwbax+9FB016mfEGAF/PyUa3kMpMI0WoTZ2KC/gVWutUlOyCGw
CJiinvSWUrPMei91ckyVOn+KfZ8mkQM/22XHVSEUuz3ba7TlP8zM5NdtApK63spL
aa3rJumYT1kKxNDuZVXYMH9WLZtWtEqfMAYPmi4ry29laDu7EK38/wqpolzqEqy8
GaPXEEIT4ugc8EJLmxlZACwOpAJ4EMN4MOG5t2TOSdIjXSLGO7/fhGOizgBRhtav
t2BgEjlFuHELznagzh087KdsNgiMcTXZihjnZTJmjJvhGRUH9u1jN3Ep0BCfSBAx
6k2I1+QESoYA+dWaCjBvb3m7IXuLGylbolmGQlNM22qzywP21Kjr3p6lc+btKDRY
WVffwImm1OgLZx0KtdFXeKXt7KKQaYlByWZiO6rXva8tc86mhLZALtdPdZsPp/9k
AE64TqNO0mZP2TqbxST3VWH0OPL2slVHpuWTFDhkMnap14NhnnmAwDCqbBybHXmu
B+3aGGF4rkGF1kJ0oU3k9uSSgPuac2VHceyb98gXuDIIJ/RV+YLJM4BhCywjpuBf
FsjjqNLcf/iNGhNAuEgKrs4fWEXK0nUUOGjad7ghKXy0eVQ5p0vOHvTlS3Ca6Pnh
EAuep3Y7KFOOWSRXLMb0WKDZ9dM4rzI5P1snyIFl1SfHh/SImkSHGVJVRYn1kXWX
gXjdbHcWg+nqZ9DyMG/Cf+HQmFR72O+9mvRBMxs/LQmrx+q0F7MAJ6QcF60Qm0Nf
h+BYJTDaDfmNzq4w2qt7E6NX/Dojz8j4HIExGeZwp1kdgEKcTL5My1zXcA6/1xFX
AmbOPbWjX/dpHW3e9krxBusvmzjeW0hP0xuytih/8UfabyqBBO55pyJT6CyQFej7
8TnWdDwnXPEYfWw5r9cgCIvZKeMerf0v3zwPxsUzRwuURjHseh+514on3hvlnite
EZTTls/slNuwHRGQgzlIaQXZMmDU11yahkZZSgbURObywKxZPh9d40/j6EvxFVvs
5Zlzz2yUPaceM/j6ftZ4esY7LySGaqMhUfAQcRCgN20fCY1LkWl0gmbsvU7IjDPv
8qCCr/BahpC3gt+nBYdBEOTLiELM6K5FXqgIIzhaO++EwpwqEEf17xAX9vYP9AGu
1HiggMeyG2Izjk1uRNZTCcrqZa/PSh6KqqeLixIHMWJbrvlST6wPEv6SCTAgxZfq
to3513NxQGqT89EF1AgXtvbosvVW4MmDrmGuTdOR4B2o0kdyByxnOTmnwIu127L1
AD9/ABTl4A3ruz+MUCyadyDMJkpOo4HPYGwj8msHdCIS/KvwrYB7u6oTYyoyGi98
Co3UbCM1rcINAsqYoOJ92uXeFBh4CIhHPXzcj1O5I9bzv/p4n5AF0FxGqtfkubMM
WkMda89K1jGBEKSMVn2qMwokUAXQWtyajZnHwOk1ialseL1worW5Fj3orZGjh9ar
ejtviyCLag6jYNAlasnudK1JQGRYsBTxALKonDQJta8XnBcHBXUjYU8k7W0ICEE/
z7zHTi5KpOKJhDGhcv4cynYer5DfuDZWilroMPYpP09LV6xvJZcnAmTNsH1u1o/J
olDx7GbdKN207+aqghz8tsoMviW6/vg77TAt30EeEVlRH/0MLaZuKfh/gaQ7kHJk
Mg1RFHO0HVkmJ77QluMlgzkob90Vn7VmGZpOHipscldpqoMMK2dgNp/LCWaHqKtw
ZHOM3gvdJWd4VYQcw1I0MZSHCwejNn5LnrnVL8Fy9cyuQ+F91bksUFXYDD1wuxY1
E7FJ2C9MYjKqK19Y8sx2d2SjTCtbQYYqbCTYBSFsjdE3FN9cXeeUsIqabOVASw2L
APTnoqsNJdcv273gU2CMXTn6HEAl4i0wNnGa7UdgqDB52CEjsREx4qyacrm7rEze
oILxQFHys/r9Dn3Zf11pR4VwCkWPZyLyCUeR+S8Mrkd3WRhdnB7NYjz68aWW5/Ue
vOAHkpQXrU3HHkMttK5637SjtiDqp21VnXFx8iH5ypTMYYFSV6pBfzVNMf/0k0GE
OYq0CPHyJ0bQG4FDOBMfKUS2KPDKZOOP3W8/ToauZvJdepoTS33bZHIAgzknqr34
a19r+Au1C5pkFgcxboqrwq+VCrEdrXKdYQbihk9cI9NweEvkGAIdaAov97dQbyTL
uUvmrQD5e0bF5zpbfMBah6ZqmgkSx9wiNFtx3VE+Q8GHA3SAApagHWjJb3EQB7ea
/4oadmAWfKEsmyKcb4lWUlPqTpb/WmJcuhBl0YL1yHu3wW8/dVFIbZq+pNIcmQBg
z0Ab34m91K3cuKvJrTZjrX4p27Y70pkWDsWQ0eexhne1wT5t1dqJNa/ZNtTDY8xF
0BKaYhbdCPLKIU3IfwDt9aOlXnImu+GVFpjnska05CqSXwDATrH3dIKpfJDSi1ZK
9AFj5iExntzASw2nR4UKrvQVuOwMdBHk2K6e3cSRm/FuMMxeVeT4efhnbDCoFckl
VKqk/drXio4RMwOQnMWly9B3492lXfjs/nje5py7jHOgu8k4p2ECA1/2nVv4MwJK
7XsvRnK2hpLdLUNeoIMQsTp764pILMm0CvBBkk4bAW6ZmUbNDWBibhKDr6S89RGM
d19UvYJ6hfEq8hPdH0UrZyN8+OkdEOakaGG/DfTYSn22APcrAKqUHHrAkObPEwNp
VUDQXD2xEfAt2f4aKIuOWdlZsFzB3mYrk9zTXnpXO3RnorTMcTDhdXa8FC/hcmTn
kUqfsQKC9HHRDgeidLT745x0efIijj8Ng0DYiDmfYBpSTYpg2WCUrL8g6S/lSwNA
lhH6IDZsSpB2a3hkBZgrh78zVp7Mss6QvksJdskDynbmqrJbfzT8lb04CedEl47n
HBe1jwGUUAVi2la9wVzndHxvc6jvyUAK+19QOk0NnXUBJxXRGyXTW10bKSQ2F11l
GQaZT2JMoiE6L7XVJvxqOolcZrCPw6tLzPRamX18KNG8yQFn73oubuT66aedPXPu
t9bt5FpPn1dQ8ZH/GnUT7xsu+WrjwLHQR6MujVgHzArJEN89wg3sZiva8nOlQbN+
Ah24zH+Qi4QnVUx6hveXWPLX6vdL34zdt7onxVJKLivgESUyDsmt+S3vVLuJ3bI5
/2fIEG3SYmx7nSxgBExEFoijOU42XToPPq2eoWWO2LDJ3tFd67DBHHz57OsHeKI8
zGMmvXlzcZ0qahCG2TFDRaV+GhuPUWXqfWSoLAqNAUT4xlqd1KwDnlvRVAJ5NN2f
R0nQbu+kaH/L51b18Ydem2TGcET/WE01jL7BmhfaNBl06wuzO9q7ioLt7mKIZWfa
tOkkH+3rhJ4eDU+eOECKBaKtgn8oeTX8xSqj5t/CDF1LgfuETZgAkRU3B1NYK5ls
7z/Z7cqp2idOmpkzFmWy3NZFmhD2to7xVZw7/aiZFwCO2fJgWPtv/XyWFpT/33mK
X9JNzrVUL2vE63AeLdaE3LM8FU8QJcmbsKGKtfQgVCRKIC2DrTVkkk9gaBljaEBP
Q26i4E6D3mfk6xC6Ky8/Z8CvpkXp/gaYjdWOgV3L9IPBq7496vV7olssKkNPPEFA
X4ocZdE9px3UFI2SzOJi81tyl/PV5BTaD3Bj69T970fLZ+DmHlEToKjOXFq+9IH3
7J/KISZXKqlLgahQi7+5DneixsqgdTn0k92zSyG0HpAcXdOhePOB6AqMfapYYQrw
CU+UB6MZHSoQbbihFBnd9gg1CVzRXlQqLJFloRhw+qB+zZukFHt9U7kqLc4RyqQ4
sNlsxnIERqR9ZyRmMGNrUDqXqz5v8Wfsq4U1ZYWUkoducOv0MbxR8OravtC/UVOB
FpCheV71t+WWAcyC+TEZUb0/5cXR1lHVyPwWM6eb6iBgxO9lDjb84aH810gClAQZ
8lWeS5MNylZJd6tXioKsZkIQ+mZ8qMZn6NOWCKrE6f+sUIiOgfqn4YFhEti48qXZ
5TXa4G3+rJwn1vImZJnjDKJ/tHAi9Fm7KjKKdd3yvc3XwYEWgWi8wE1tp4KqHfOU
XH8WVK+bmtEMF7NqzHfVZvAlNnaE7Al6ySFQ7M/sOXv9o5Yh93j27r2DjNfduQOE
2XYg1uyWwz4NKupv8Af5RsArxZVzLkSIdtJJOgGvmbTmWVGBdO8u0q0b7SjbK9B2
6JmehO+WkHAB17VrfYwwVaNqxDyxhJZXmGPV/ewxgal2oO7zY0cTkgks1ChscAQM
wtqqokwsuoYSIFJgHsBQKyUjPojDDnebJoYsD/BcowaRw9PcXgYOD6pwLT1bOrC5
nOX8KJTpSVsazml3IMUi4ywxk5J7IZUVY/G+vivImNaeF8i8z6bOrjKEbEp+WoeF
xe8JXYdLSXavgiMCynaH0vbyO9l65ZHjNk9yRhy5/1xS6chLE6uj0y6vraS1/10s
fx/ZcUYkpY4N+yGxt/c9mtGbsDxG3jGr1HfbyhR580yjUU1BRK1PNwbDhVBiXV69
GQhAhwuhq+tNnPWNr0ZaGjgLm19xeREDHsYAAzNVBcjFRMIFy7NSwK910LDNQ2i4
BIQ5/TZcVs9PCswx5b6UeZ1ECRq07bBpI9evwa7IxucZxeGoP9K8mMBBWIER8eIE
+/jci4FaqAijh9ymKKer3sHS8NA/7ZAuRtQhPpevlvS22HLUFLz9h7vrRelVVMQz
ZmMELrxjOX6xdOIoio532TMC2y/BqXzQhD+ickcyyewIYIvKWUCwnUhsjzuqaLcd
UbiG1ayW02D2QiImORdJl0EKUQLE6sglciBSajbITItWPYAy5yf4kGb6VToexrqb
h/RwrB9mh8n85NREeRSRJjuKX9I9beQnK4RRSjQuXTUHPJ7+2FXMSNu273Kn4gUZ
vG+FciCz9G1U1vKpwcof4Eoo0kB6LvS5RDk8oP+7rjAxIYY2E79R2qXLLuR7Bcai
NtYtJEeiHvi9f1gtsxU7eWto6fd2iphxqcRfxOXidy1MbUuDMIPNIPNaHtvHUmu4
JQ7y/mLR3jRsst7+Qtcvs3yUvaSII2pcDs+ca4nICCbAv7bb0+zgRHRwUsXSIiOa
1VtgLY/5WkRn5PSSofV3TNP3UKfS82AN7Cc3azVQ2jS1WKsP7qPvernirL8ngwOg
1VKBdKF9qq9shchdfl9vA5KXagZKjtHFAyFpZtigE6tzSy6oDuP4nCKrfsO7P0hl
jbu5RC3NpIxKUZD58VDxV2lATtB7L2ILQEYtzWPMhnbbihUE4925gmYX6VbUXJm8
wf3J1lyp0Si2cmDpGD84Adxoq+9/uxuxKWdbHCz4dE/GNnX07HdLmu+QS8C4wAHp
A3hDpqF5jkLH+7nXEj+PxjfwOGsEtLeh+O3CMB06eKDn/D41xdrTSwKDeUmGMZ44
WXzQWC3DX/wxrDg/Ys0iVC6rE/10KMZZbVcn3ElvdEnbImA6a1s+oJTl2UQOC7Er
XCQk8MOb0RNgKO1Rj/KbCymWy7Esyjk6qH+92+yQOJt/w4+03LtrzbkoU13OkKni
unZJY7CFUVnDFIsUlfMdsUNfmgGeJlZNl6Xfk79Zofad+rhuqXgAqnClgQoyZeYr
Ji1eSvPIy2mI29TlHBDHwLVGShuUKJjm8VwqyyVkc4RJHHuJNktLnTjHouJevrO5
TtNm1K9HMcBXwzcmKDhZiUA7ULLJAAFJk8PGPG4O8Jga+ahKC5lWIRqjBQiOfB+z
Ig06uMNMnn3o2Ys4S/c6m3MXZgQSRwIN7FO3aEJi1Wyyj1kUV9CagzgRy0G0zfdq
guxav8B6WwvJ+uIQc8g94Rw3OQr8gZYxXL4FIDMeO7mXDNmIFTkrhDgr1kRRFKmS
ZL0WHfsodxeiqF5KI5aT1STZiLD8Pbnk3I+39JOv7XJN91DNPODebOpCt/CjRK20
KLmoCDBspO+JwHjcKbc1jsTPVS2U1mrti6XK44fdXvhWCfNQGyP5kD6df782IuvA
ztpXmJ7iCU4RCgAnOmMInMsccmViz7N3jRmQT5KhFHxYqfHczZ88eYvs25tRJv05
ce+Ay7ndaI7PAwINCYc8rYAA2ajxrCOoP5ueoHM3MgBNE4OxR7aGsAb3XLw27xJg
PXocyThUDJ8NkX902IeINfhX1OMWfg3sLX32Cr4nlqWA2lwKKGQ7JedKhWD9s67Y
upgG9I5gdcHAqxD28MKMQ2G1i1SQgbqRbWzpxLkGOarZGSA7py3yuSXMOy0yIjMq
8Fb8z+kyHJy/8MqyR9Wj2OhxSB7ljjXT8N0a4bxvPLzkYyhqVYaVaPSrRdVvNQed
+58PdN2LamsRTeDS/Kmf7ee1osUhftWgmf91Eu8xKWRtYFbanog9iKWv284qhSfG
5hgXl2dRNHD5PJ2C5cK1n/aVNXjPEdd5wGQhQBliIBwoQgVC6hD2suDY+RBLPPNY
inHgkKg9DUfxqfNngYOiCd916uW5PwtmbK3/LDEv7F5/GyKDWRksNKZnwoAhiEBg
7paUVNGzPMww/DsG8QEtjePWhqYOKvFlid5/PRuAyJDPvFlXlC9JIIu/9+FC6bnS
gl+NLdU16IVLSkPHdxYsmEJfKVxIQCrF7aI8Q0dW0hxCuYRsvmbrMks5fkoa/vSg
joVAuRG8Xeb4E1aT+/SBq7D0fdAHonfAfS7t56t2GDZBAovQR4yjS8maWv1xa9Kd
AzQeBvFGpGk5sPRO3ebaxl+37IigGJVZ6N1wwWIjL5Zyiyi6KTPUT9fN1WP9f+eX
zUP8+uaTx1iOqpgUKA7FnYDOHQiYE/3nrW/vBDhsmzAXC5kDYYMuO7U8akHenAr4
Kw9BXmBOxoFxZ87aKxj13p3Q+SZZxHlm4Ghk5nVY5JUe7s9+rXaqa8EtXsoi+fA7
zABAPzuV0krDun8aa1dX5taZkJPmm/xhB4kVvbkgYSd+F4S3DKNOfAy7/0uZUntf
AetQfq3V5xS6vqOaEPcf6CSuj7w19fvIqmGlsove98ld/DHzRGamSmvILcZ2zfk/
2eg7FQzE/3l/WClmk3ZMmDV9CrUMmaSFa7uaIHN9hiNVZUDS02aEElDOpjfMjnoE
gAqBdVdXTnzhO9+6SpBYijnqiQc1PgXgPnZDNGy1sCstJTsvrLLvcxvt/s6ZNYSL
AcAtTQcWNs5X2g742cQNPnMQLHSeonvoM3s8B5VU5JVM34TFQEbIodhyuiHcKSTz
+k+pAwoi53wDzoVTnLv5ktFVw/HNBg2sdps2podbJ2dFb30JYUBN+5u2IxViYZa+
B1rEMwV04wnPyp0fn0RPTAcM5hVbrZmokGIwR2Fp5/+GRHd+0CHfmSo7cy3VIbXk
oS/LFu9YHVY5RzkHYF+6qBFuzSXhEBo6IJvjVSqifkxDzf/6gbfZGA+REE7MJQyj
TOi/uAEwswJ4SNNTQxux9cKdeu/jhUEqBJ4H9QrocTtQRoyoGBx1DYIneFOv7a2R
8p5Q1BSaOCpF2xg/IrIW8oaWQCEBeXL9A20k6+swSXcczhHPSTqXE6CPnNdyw1cR
fuL/nd18qGW3bxfQ9GpEOT96o6Gt4CLEZKCR7h2PSfB0FsfhZFKeZVgDRbJDvgiL
AVUMlGCoRSB/TWFDOMEhJTx+mvT0lN4vxEZpNugk+DG4u+RApdKk0u7Hr59fhAP7
UTZiqrMld0pA10gSAHY0D5Ewvj2O9JsLlzc6PFj4YBADPIG3GEjoWHb6Q9Y39QBp
xwP3r1IjIsX+4r8l1zsHTMrttnUUEbsznHUyT1qkbnItgtA3lsooLnvfzLN/yeqm
n0cTXBgUnN9XzHsafwfNx1IR6eP+IehaH6pIPLOhOhQqrv92aGxuFeciITrBUgaD
zelfyQBzEPz/Yvxlxh+yT68ZLwrKg/a+HkNgKub6ezGZ0GduiAj+5iUPEN/jBIe1
5PlhCNFS1r0fhbzF15V1KnVui3TcmphZ0Ua8Aw1YGyUMDdNYeKmy7YG/Zsz+KNjm
6eVSvm6VSPmQReTL1c8aTHxVRLEDO7FnScOfkEDcryGj2A+ybJm/k7PJW5Avu2e/
HGSk3lqc08kKAhRM6CGZwY3MwfgT9N0vf8aRijL0CYjWo4e1Ibqrs/R89lEMbmf6
brzBon/V5hRRWN+30I0GE8oQaX69bLPbkwfd52ZtFIGfERuNNrsFMM+aNKfA5/AE
eXgwPRt/ra/gLTBXNKLx7Y8Hz+VRdHjVESd7yxNgUE7YXedneyf/ue6NPteYK94T
+j8ZuVw7E+VIcM2ur0x4l1q5uCAUA55WgCn69kMVc2Y/Waw5TWZ9+lYZSUoD+w3/
ZMzLQDORHijqW94L86OY7sWmqSqoEhqxMS6bpl5p0VCn5VXH9JnDo0VLJirY1+6g
xvBt2H4w+Z4mwJddkzziqvRz3kkadSIRWZZg9njGAvtBxFKXnmx3khyHVgJE1iJo
qerBhVOfJIkllJd77G3buT4nAGv2WqSjreDQyj6/V+i4/eD8cz1FHgl9FQ1p4XMk
hfWqV2q4fC9Fi/rtIUAYLq+zE8G+QhFQWFMuZ98EKiWTbBKuK4/NG5YP33wjHnbt
u+vsSp5O1DqYLjVEwLSQUi8KGclx0qKWZ1OLjwuxPdITbbWGgw1Ee9lXO2nd2Umk
foPpS5U87fEwFeCmTokaNOyc3U2+durVUnkrxPuseo9ykQz0ovyxgBu69XRHWx8O
I62PXsV63xESstTKHV7OfaC3khU3IYG/NmtqUz5FSVjNyZsgfjTQteDaGuOtk8w2
8AnvoP8lfrZkOJElbJ+JrkXSArKQaRtlLGuY1sFa6dfs6UZVWdT4SgaquTYgKPWu
SS6+S/WdRbUa7ATbtykO1qt+3kS9N2nESNBSH+SBUUm+ajgehSfjKj9SIhILUYab
UH1ZG83O9dtKOgGOqRt8Rkk9l3j/fM9PANZm9oR9w3WNHIJ1ZfbMW30il6JAiGiJ
bIYsIE7BMyvZuWRDkFbLQQLWNaX5nSd5ZZByt6um7OGuV6tNcFFL1RrH7wte+9Gj
8PG2gbjHNR2E+/BlfxB5VyuKQnyqPgC3LbAajNLwTgP//N90DtPQIZWsSuP+MbXB
zPtS3JhDVkXa3bOx9zp7pIJhmyEnXTgNWtN80TiO9qWrQNIy3XIfCCx44QEp1TJq
aE4Sw3FXWdAAgVam3xt1qLdFHpudtY8ZURXCaLZDzdW7Wn6Es8aYtoPO0z7WulwP
TVnn4aASuIkWUF8ImkYM24m7iAFCFdAE4sCuakEkoSU80dHavrPBWEuTIdOe7tOD
vaj58LOntqHY92rGur5gfcVKSUuHAcBepEgMTFT/yX8hBdCMjoa+qDDeAXuO++TD
eZoZnfYDVr4oKEV26HSNLeD/qsFnKE3QVLGeg2wo21AzQUcEp5Ztnywdoi7wITgd
r3dbEgmO6hRSFy2x5XSkTG4ATMNO0hvcS/BHIzS4kaCVWC/i7UofYagJuYzlaDPo
yVAbjn63XhqjJjClo76gqiwXDzTIsAYN9I0nC83XpOfkFFmUUEhHiXYD8m5Zl2q0
Oj1qnkPoFskF/Gh3ms2Fpum9CeaVQuYjDd3n/sTQ6fllZp0cHg63q0QPDpd5qsLg
ZbMYS1lUTQccpBPM9bzD04hHdGKwkPwOfcSS3uogmsWM99SR0mv7UmwjNfElJlkM
FHsp4Vge3e49eAqbkRkdyjP8gQZuyHicOWGvjwkb9gbNfXLbwmLagvt2WG2DTjy7
V97Ls7I5lXLnJkqnrNJ1vUYRJEnd/ABvPvGeXLGHDdxhQzy1vjsY0B0foOCIoOvf
FXxYStrjC9YzdCh6y51XsYyA1DbzgTMC7yrSgj6NLo9zO3G7nERByjG/q90lratt
6EWE3YhxaFvkCFDyZriTfVlJlDOEVWHiYhnE+Xct2CrHMBFJq918Sox2OrriWuWf
J7BsziEPDtCsYcQiXfsoO7I/yHxllLewNCoNeHKxmJ++tzQ2T2IIWwWO2VKSQiUX
7weJoeWi0Xg9TAOX1VQO8TnsnoxVVP3+8D5aqU6z63sOCTLfukUjkJN95fQ6XIUb
jlwqE9N5bhYkHcNbqDCcjzhOF81lgDoRcJFO5WjBhGmG6BYSS3UsedYytvPPF0T2
92fZuGSyGsli6LAN3/CyFs+o/uuhEKina7GP4GOSFX1ZudCwWv0o94jNpPw65YG/
UXPpaKBXiz06b4dhTq91VoPJ4E2utld1zylWlrPm1yaftHd2/TvkR5vToyvdsEdW
d2MHHGKc5NRWrK+LuLJAdNTHouzue++SgQwUrGMlk97uut78oxuMBWcE8pBLFoLw
3VHZoTFdePBBOD1rUgWoyi63J9cnYG6+nTuH66uwAPuBDNynNgrFGTfbbBcdykjI
IY8XTtV1BTfcnsioOoOlS8+1H94GljIwOO2L3dwTpVFZci2piTutZ2Ce8ed2renZ
ZeGsM/Ef9dFVfaIzBY30lBQKYCoBYHMLOQf7IXYJeEmAsaSVJKRKNyQFIGeu9ugb
7ZzzIj1TsYYY2WAbWSqjtn0I2RP5HWowy7etzDRdGBTH8oMWTZXw7G+5H6HMu1AE
r76kZ5E9cbg/HPa470WmUB0sHcZ00JRw+vjoRX4YW0bXGoa4c4mqM1qVW0bHnam7
JxRx+78mRzNDhyN12jlfiats7yM1pt6KUfXq9nLjZlN4FITeVAx4A2HPrLBmu9eb
UFim/SpUYVehG2hC7+VlOETSS7j/Ah0F2KzvLXhtupvcI9MH3fyzWCOAfJTTjwee
5kwLgil1e3VSMdraVcJaShAqeyhLM6akjL4Sd7FXaXB2mO/0Y7E6bz+G7lr0iO5p
2G7eI2sgR33fQkSW23GloQlp4HfiFRtfBnGrvUJPD4di3YatX2H4p4Us+Q3iYanQ
7QZOPsWTDpkXdxbz+ga9QI4sHs4GeR7BARxSiLpboQyDiHlSTbTWHKN+1Kiv88xw
lXY3S2I4TGi4j5m8YX2+mTpPV+NxI6URyAs36RHa0sXnQFl3+SvLyLRul+vsRu6+
SZsIGOq1ayK5S/WjZ3rT6r0vJBJwR2FZC7SchVZcjNT8rG5GqaWkd3+SNEOn0ZUN
tWve47JLNXF/lVDUkklimPmT/LaXUtbLHODI1rpe+3ac6zOEhZl4Ko+QtbpndqUx
tNfkPpBaQHBP58vmQjFYUSO1DV3auVH99wDqkQPORAcaried76GFEhgAEhZdF0ui
252hSqWIAk4qSflihCgZ7xWdx9D8xdzbe00cSRfBNaB60+gtkxd2ZyzmIcGkyHKg
fX8F4KLiFDq6azcF1iqXzYqdkULmxPe/tW8Q2Wo2WgivudhXoFuuQrjg7u8iY3ql
q4CfcM/2OI+vWkMUXDDx9urcRQl/7Eb6wpN3b1MX+e8IPhyB81aXCobO3S9X7nW7
D6pA4IM6UADpQBK7JOhPYpaAWPR1mXOM0tTZOzLCcJvpFTeI2RWO/x3pQNodhhtl
bImFvuOHDkS3Op3U3eJJ1PX+M12+48fbGCJDMtI5UZG4ItJdSOvZwCDSQ5oD7X2f
x0eCxADu3JkYbERfZDAyFXJcIdUNkeTPanEu5SyBWpcmeQCL523c/0dH4lzxThxA
4QCuLYSqK5eSXmpD3QqC9gUCN/pAsUJyra6JdBsukrW0Y0lIIp83Wc0/cg3xkJ0h
a7ZHV/Kw97sqahYs/21WLJs5BUNqQSBS5+1OP5LHh3A2vkSQcv/nV9STdLHESQNL
nGF+4kKy4s6KhB+7RDh0tTR/soTwhoADAIGNuRmfBp2BH1m9j+OQeqIHQaSLdnWO
r8RUW4RzsTTSAuzbE2jMi7OpYOO1KqO/VYPwHq1yUptzTtlb6PVsu71+7iTA9hk2
hWSoVLbor0DSnnDGr/pnfVlQANH4znbaixjv5enH/WGgIR1nBLTQOlDEVxYbqwnh
dvZjI71hUczzr4tGfSWAoirJrDN/N7qHjrbnymVNeubQEkH29koOXLwC0LOSRU/b
u7AEF1xvxRO+wPCU7/uLg+P2otaJ4J6oCfrR7atcKxPyyhJqwm7jwnVCVQ6Uq9Px
ESGwdRnGoWnCGBCl4fXBRdL3ICuSvuYqkW8jg6CGrwEX8NFcVzXS09LgF3M41T2t
JBiUqYHCedzmYPMF/XbKelP+u5mGS6PmvLl5FM47P9z77Sui/ecDSqFv/13xAwBb
rkxqlyEbkvzr8hXNFoVuncmcfCp1nVqx2eQUtrS0TgY7R+nDoYxMi/Pfj9ttCnw/
bosL5UDt8KGf7CVO2WzEDwAnPJP/ZxpCNJHUPm5fIjczN31rPLgeRehJ4vABZl1u
nwQBJzQfGDKVZFrsf2xAEN7zxAnZ0ilkRtwK1fvbgWem2rV42QJGXBrAeJuIMFis
Y4W7n/foupgtfh8rYYjZRq9jMBH0LJ/IcTn5NNl14XRIZFYhhowtyhZ19fAh4qVG
fu/9mWoX2TFxnb8dfqO/2tdYH8kbTgCP8934tt0W8GZxWantFaLH6XifzGsCbKdM
501t8eqsXssvn+FPTECyKvyfBJw+z13GrCSn15mAntLnJb5p4aBeQc8zFM9zZXXr
NezJtzyqK9qRFA087lg+x5pmLLr2oVPg9X1zqMLYoke9cWA/HGHQQfWn2kL+Uu5B
XJpbiUrnDQYZWRBiaFOzLp0fuLIixvcmwx+R4UsUmk0h87Gu3sAg+/q3tECw928j
VKwtLaYiVsEFg8aXUpm5lzBKZL0vW77NbqPvchPYokrOPhOCdbd7D3wU1sOkt6gx
pc0cjVdt3F91JTM91kBgr+gSIp/bMvSmm6sQA73gaviJk9dfSpPSxzEKzSCXR3CP
ZhSjlbwKqjTAFStKDyZ/hVK+YV7L+Le4rOx/EsXEBFRVhRDGTRaEYtqCNMxk+uGt
tvw+1CYQKjFHhHB+cU2bGj1/bmVGECCuuvy6NHKNq6AQjocCVTb7fW7fhbsVz2qL
/vvs1yLKbQc5PApDv5YZktIje4H1xhg3lJVOY16ddXAoUUSkjuOLcZSun5MUmAU+
ysCHijPd7uXL5YmIlpBELDmPphtnGeCInkYdKVXTQeiiO+wS07kIqZin86iAgAkM
OfMRBGQVI8kx3NZjVnsSrEF6MdHWyuXRuZl7/8V/2sCPasbSQAnHV7XIhrGTpcW/
GvJxAqaDcCZ9AtTjG3rQyYzeSOu3zZ9J1uGagMdtYUmp0y3LyUgfndMiiUXXlVri
v3GnQTNL7R+57BNeb2RVSLnTUBbgxrET/g5rvlzpr48Kr8rMloGcqExetYPw1Pv1
7W+AsbAVPRnTTadbhV7GnxljhACeT5APH0C/iA0u67Fj9gyZ661XS9av5H/j8bes
3/zU1yrLLtWoHsFwVKl1wDPGuRNrkbYvFM5DJrRrR8fCqfF+HZSfja6hiE2icKBD
Clq0S/CKFkTQp29i/R1vNd085plFotrFJFgLX/kRDa/G8bQO6VVQy3+amrlWGjca
6FNQ798ekBaOz2FstuQPKuVAL4AFGEnz9bg2nsO20kQrsMY4+wh0CLqvd6urk8H2
9EaMH0KO96AZyxn5P2DfabLMn9zwlKVTOSTw3SMh5iohc8F9Qi7wo14JUkr8Pgir
zfKwNHtUjl8EUWjfdchyGFVxhN6zxJwI0UbYIahBoXhT4P1UgmIAz7YkJF7yatpa
eIeyeM5VN/TuMmioIa1tBvjJeJL7gS41Wrqtcanx0+lwAIVcuwRjl5xPa2aloLqG
d3skCHkDew8vcFFlbm3L0yd/5SnZMb0iLuLS2MsPjEb2hWzPPDMGRZ7qfKKFjNFh
crRI7c4bVspBnRteHirAhlBkNr+uDzfGwkAN364kBXXKlU/ni31rV9r3oRO2cnSe
3ZWu572hwGJx4YQ58ZYR79KslnRz0l1EIrLKxu8Sv0z41zNPYIsM12tzdldFOuKd
gdsyNlnocFPo5HKKKa51r0T8SeX1j0ajGdojLkWUxyxIhM0mDp94c15qUpvn6Zwc
jerkCdtUm2qlp4mBlieIHR4qLpggtC8QHL1F3DKjej0fLKHS2A9SfO+//ZwAPTbt
CBg6V1kyanNrU2zevX8M3qv8++CtsD/J9ubETS4DouiOxUyyNNWkTkKTzCdHsc6v
dX/baU4k9jyKOIGsOxjIBzZsLRDQMNGxQUAUYXJAAPhVxN9VSRe6yVgUf0LUxLhg
UtpypXILLF7A0B5Y3CCBSEi3xmdLlcxt5f7ib5xh8gJF3rNNbpGGYl8EnvOVupSp
Njfow8TOn1K8ZBSvuwZwDY/AMk8pfxe8irbgyfAz1ZGzUXybMDDxRp1lrX4PCVeG
9zVaMhz0bU07PCyi3xohfhYNC6SUDkRsm/Vjb6eguzROcr9gbNMF8C5wFCJt+2NQ
gbyl4yJvVQNEzPejSN9g7X/1XFKXdIhx/WYoLYrxJMaVGB+06sfbOUeJVM43HRno
bnUpDx1dlw18obfgvVHHERf0lVsdgDS7HAnhzBWQUY/Y5e64A60ttmfx4m6F4LeC
MRiQoWYlwktQ1EXEI41RnE6cq2StTCh6D2r/08dsHegKxtV628eI2DFHj6eApGgL
LMRpS/Lj9euuAJgJJq50rugYz8/4USsYWnjfJmoVDBLpyCiVj4bAUwDvZVdk2Og6
Kim5fUEMfr05K7rpmYqHKbk/ngjnX9wDqfmjrWe1GAwWkgRVjl0ntI0mJWamghLQ
YA/JerbOoeXnkiy310Z6EBVT6LhgZUMILxTTCP8F/d7rXBEIY7Qf5VfH2Y8XdRU7
I1UZEmBof25oVq8oEGiZeR82NSQ3pLu2rCoOBAGoP9UJtDUGQxBd8ve856noLtLt
ZhE99VhOOk4C/A7HPD1MUkVbxcu8jnQ3X2nju31itqV0OtM11TcgRrsbRCRQNrOP
wNrXXWd0GJ6Dh/zpN3ErMhadDtcFeOPvjMHY9OU5nf2sujTMqWnZlzX1j3jKD8rT
IKjQbY7mw/KLHWS7tyxtfcStGYrsmRvd54pRA2TSZjAytftln7yiJceEsErAtrjk
lEf9nbyloqWM7icHn3Z2a8mvsu5I93u6QbSoshie2S664hImPnTAPwZM7hR5zye4
/mjhcHB7b3rdDu88WQ1uowrk5dLrDRkwbUkLG+HQ0XPDbKpRjc/eBM5U54Pu4+gb
NwOlXASn0OSCfeS+JMF54oezSEryd8RW8ejjgWtU1yZ2uOS9DagmrQ+9sbgJFdZr
kuI0kXJhhxl59U7n/cY35yu9Uzvb4k4oS0Bw6vYW5VKSUDKxTz8c/9mDY3BncCzI
FOK5QaPp5vvnG2CsXNqBQiUAy9iftc2Uf/NKR88uZe4Tte8wyrzGuw9drMNQh6u8
UWuBSdNHPRsOY9QHpHPO0n4byNrnyG5jBmv5+aZazt4F4OMxjhgGagErQ1eA4zgN
N8OHHRVMOAJZ+TrpxnebF9sygPCSLNMR5FQ7Q3S0n57y0RMWEzEQd1TmkjiwPN3X
ULfRQ1vKrsta/cH8WrAduizZxAbsxyrr+f53GnbtfvjXnGz5lcNsniTzr0Sob2T2
rbgg55Hn7Xp6PICSvLyYbfVanQMYzj7LkvLT+2DyOXazapv/pc9+kleBQ/AdntD4
q2Xj9W/2euh4zwBI71gtDBm+cW+UdoZRCJaCfOQ3KTBSVSNtlKA/SzGJI7KpU68E
WNxGvGjsUBNMBV1wtVHqWZC/AeUFcIou6uK4jCPL/FeU5lmmNa1lLLRjvXyT9bbm
Wc9ycJpwmWZkMwE7g1snabOIPWP/VqIq4dDxiEvsIn1QUcZGDuPbJjSkhOBSr2KW
H9YNu6OfarlsNN3M3TTz6famZMK1mAvfy2tIGkdaVR+V+xAM2fsMaColbutDFIOp
lxgzWya/71RGqVolWbh7bQKJIsaK85xZC9/tfsEWKVyn7ti9ANnsBy7AWks3fG2m
lVmFehL8tehsxGqgR4jNBP5+NyoepxA9qcqi/YfUXYMQGg8VQM8E6YBqVVGnLVrG
Gssf/p6Juncz9RPSt3Cfs0hW3T1fw9XBzsqA82E2sGPXP7JckqJhyhGwIY6khfin
mLNv87e11Mb6NyJCTnSjnERsBGHlaJJZvMeZJJ9OwV7+kk1S+RLeBBWnCVtfWTID
D4jUq6TOxLk1hr5pG0Z562S+/XoRsbS7OUFO4MiMGLIpEasFLONkJfOjRln1kXdu
LKMEo7z0ZXXJkF82otss24wMFSMFgZrEZ+QK8zBOOezvRaxv+b643SCSejCZdgMG
VZG/W4v9EkwWGyAOJdtrOeT6/iCEsQ8d+fTOdDs5ZwmgRLMCbjBDPSv6RgRU/+tA
6NTB+S7siuwE5JHQB5hV5vZwisascCN3CVI6NjgMtFAWxgosA30pfBowNDGqlH4+
1LzVREIqV0fL96cE8RIt233DlgnqMpVrH5Dt4T/bhMyjJ4ZXUupiyBo6APD+ZcuO
ngWnDYYMniLNLX9/v3wehXhJhF/9JH5xTW0YYROFP4Brnl+RXiI0EzO0rPb/gRVg
kIf0mn1pEqZmVzeW2jChOC8kXsrhGd3UoUvI1YmjJwAS9rGds49j1VEfg73RH+Wm
BCzebntD84EPYXbYgH50WbdI3uEgZ7e9rjuOrRKw9EiCbBYzyyEBp2skmwZJ4ovV
/Pyj7ZXdH5dLTAh6qjt3Lpk+hif7PdhxjTAOAagwhWFzBZI8q/kNVnYujWOjEXzg
j+KwDPn6dBsW58t1fv6/Qvo7SGEd18LYiER9UW6grOcrKRZXHxGcu8NrqRphJfKI
9t9jXS1v12srZbRkBtmZLB/kuGMt7ReUnrba59juuz41VQggNkbA8YqfRPgoA7zc
8TUon8rqTijxgi6TgUWfSaowaSetiu6bLlobrZyls7689TtpgL5p5BGlBkXdApv1
UkT2pCiUe6xnJvs2p4mKW7NkcJ9ZAami6PTm9a3J6Uu9/rS2rQEfXfqsdSQv+qgz
bBVPIEEzbheVaUZxlRHNSQANLDRDh6Ab4aJ24mqzIa/XrApBq3ZK/HsFvJthQdqv
NKux8mJdlDOyO3D2opIcaS/9+vFhoWx2MxXHSAZCHu1kuBWYHuA513Dpl+Ddj+Se
jbyGTeqi3m1K6qNaK6Rvn7WrHxq5lIYCwmNC7F2vyV01P0kzkPehUXW3BPZ3grH1
cTn2QUZLqMQ3Gqg6lPTcIAAJB/QT7616E4wtcFgcHhVfZpU2mysWlG6QOd5Vogl5
vKQWtZd8+pNZ0o2drRPQrjKbfqSZ4kOHFesEdbk5SWETtmLkWoQBcihk3SO08yFv
5f9Ns47UUx1Fp04BLR33fZ6WYaZGcrmBMaOqK3EIOfTx0xjixtjOKi/mCVXe7VJs
XELC8QTzXM1faCf0KuPCM6Jla880ZYGj1t3YALgBwCkyIsRm5JJ4w4pSRSEdEwO9
BcMilvunqYJu10bAhapO/OXE4Zt/KObu21u8hvp2U92O7DK3Yw6AOnoORTAD2mAF
YbgQNtKMZR9drvIGCz4kejglyF0jSoADPB32zixDTK3DEcglnvCMfLbI/8XCYrv6
vXCb/HyLqPsSbQsqN+EqJV3r2JVyOmKoQZdBGLemmkXLvHPZvMGdePcT+FLAt+Af
88ZPWnmNd5wgB6A8d371pZSctW5gSZJoCX31YE2KNFMgkkwjZpMho0mu+58SsUDI
6nQef9zaRxyqqPL9Nt6FPR4S+3/1XrjdJdJVlS5ljKGJ2qvZ5TfOZifopAwocI7Z
3CNMnSPL14RvlefsZkQqDlB+JGfKOaqC6sy/lseN8CBA8Nqff4SXEs+n1iOeq65J
20Bcd2ROlNopUhaDEhwkbVADQvJijoGst00EGAupdVWHxpusqoBcK3WCTh/UDY4E
RGdJ6aWaiOODWiLSaa9mXc36n8tESG41jErAkKNEVqCPN13tebRrgl8jItWf/lN+
N8FLNmoZdX4Xl3yllZ0K6vTJYwg+Fy2akYU2DKS4BWHfWFOF7h90cP444s8lETpy
6QYBud7UtEjYTwsbwbtkQwO6UiOprol43usgH7AIBN0vFlLQLQfrZn3uWbNMF8Fx
k+TfNpHNxZcI5UzC+YYE6AEdmVbfZglyB2MhCLUeF7k6iw8nIjnGq9u2IlIIrJWW
axN/Tocn3i3IWdOFlWNNn009G1LOvSWIJ8g7CdGS6/nUl1S7P/WPLMencca2znPP
oEiPwMc+xR1apA9Qegiskk4LxvwyLXMm1xeR64xkw9lsmWMT/7Wz5qlUwXZAUkpk
Jcu2YCrEyK+6qpniydcIgWXD4UhY+moGFhWct7rGSnF6MTmhuk6eF7nVT+vttgC7
8aVbGTuYlt49nsWxa64KlhHgHmnDT8ybSURl+1sfk6zozzejy2m3A5YT7HDYAwfL
RUokEXQ7RTYsQK1IIG9FxmnN2tRdtb4egE7SOlp48bn+w/iggjI0/sLI/ibFB68o
jzkolYoHn8m0lx1rDoWPdQ+4B4gO5N2WhhCSX6chZ22GFwKvPLTMVlvW2hVrf3Lb
cGrN6i4IC1NL334j7AR7fF8TuJAX4dD+9JX2+6Z+T1BTlZ9Tvx+orJs/3Sq6OZ8e
nq80gkbLdBiD0sjOUN3NtvUR7DwJFJk0M6SWSnUvch0wGRQU+2h63KCBfmMahkQU
9MRQSSzfPjXQxTjR+a4HjHqIJR1gUKc5L1BhSNHjHM5/xfplqySMu6aA+w4H6x5f
uMzWOr/kAO3mq1wGNhNIGMANpvtx0anhza2Awpnbfs9/6VSdm11ge3vonN7JBClr
cfflgXR4xPx5lxYllbR9xVJ7rmSoxu/dva40BvwEN7XR2TeBMdWurATIAOMA+4Jw
82G2lRdkAHK5QT0d0z4jzNrAYq0bru4AGVTnAlDE7VUO4995inf1uWNZB+QvgOYz
ifNQMHj0dDSVEGN2mToKUsaiGp6KXW2OFc8Qla754GhwEhIMUzYEUH+gPi1HNg2V
qy/cX0nRTVvHiBAtXVadbDlQIJcbDZH/lpssw9uZPRJBwBLXdqwQdB3r2VIIXvkK
RvnCvruI5wpB+18/5TMFn1ev/BwNNQxTkJIr7kHUURTzOtuf+Xjo+8A2CDUeTmNv
wdMLF4vpLGA4YrvO7s3d+wuwz9vJwZKUta390To4MRTmS0b7DkCCGovZsG61sNX+
UZz+9XzdVYon1tbsM+2AyB9srprrbzApHC1Wnw+l8voyRb/Bxx6b23UmbDx7L5Jh
/tB9/hfSsKwOwi8rfHTc7onrTtAu0sxxIuPF1IbSuKbdMWG8/itenV3WXCSi7Vcm
lvfaWFvFYV/f5AVxCxobnYsLVmazT2T0O7kauuAFc1AsY59vWeoALBuOcxStYAvv
iDtbHkv1lH03AHcIp98Mmu2TWBY6o68CG5RKx9VPA+ruG03BJOXVF6aOj5piGKy8
ZXCynrbadpTrA1BA+qMiUj+kzild1rP7DN6Q/BHTefj4+7wgMZg8LXCgixnB2oPN
zVZAABVX6SWGAUOkZVUR1T8ilFow0b70soh3/ZxTCsQjpMOUhKolCs5V+Pj+RwHf
pSZFKsCttCjKOzipetpStFM4RZkJuTL9nAk3ejAv5sp3Mh2xmXWI47osafG5HO4L
4Fzsk+RDgUheyP/0zvywNvVcmb996kxq0KF5xjoEekSval9ajbZq31Ad3vg/LbwX
N68a/CAgNL64oSvg2SSHs73GwToDy0w1TIWZEZzIicR9nAAa8MLBJDb78teDunWm
aTJ3DB7RobGSWi9wCrsvDHhRGNaiQm7mQACGDTwTW7v8rKNPfup6Qi/tqHUvwKPr
ZcbEpJgl6zZ/mPGVlAKHgNEahuMbKfkBTNLgZQdDOgg9jY5Z38lkX6zh/8tZqkmy
qvGXG6gtpnKbFbD7LzFueuh21tDrcAOZ3aXaQ5Wh4NfmUOegluQP7rc9qawIVGn+
NSUCnlJMEPEJcv+Xpxo/BthEdI6fNGbCgOLEp1BBl6ViZ69wxbtO6bDuAEbSF50E
rw3sEM6AEIFR0gbQBwAXUbLE/t6prGvG3eCBkidbt7PTd0LsvlHR7IkqOftHtGg6
wWtHkcmV2xgEz5a7ZbSwQsxPZcR96w4COA1hF0DSU56vMfh3vTYE46yTPM1/yolq
z2uU68rwOoH7VBKOukdt3Og48g13rK2IN4tWj3guVlq6FJtAouYSBqFFV3EE3p52
Wrrak6WzHLxfGRGovCQ2he1ChczzZdruBv3IFVGfxAmFH32g5WY9p4/Ev9NGExBm
jlvofB5QCxkFg+snu914MDjd5ABU/6dAqiLBpdYx79KZ8k+xvg4pofYSRMFrj4cZ
34cxdcNrp6CvRqvl7VPMWx5wpeMUV6qSltd4fq59QD5ULLRxrE+OPZHgrafGX/eh
ndTI3EJWdg5isj8iogMHk1JfPBw+d9U7RetBHVQtMwwoxOqkYdKYYSn0eKi7XcLm
XB9TC4HPccc2M/e54sPFq6ZeoeWyTP84JNG9E7c0rKdE/21VMcOERjA3y5VDuog5
E3PoT+C9tkJ0W2yj+kbWy/yVxMMvDCuQcgvnD0CQv1+2/MXY6cLcPEwQ8aCFhY5V
ME2MM2Rs8VhVxSwBRaT10XCCyBrhnsUT7vIIuq7Osa88nvakxa8Xi6yMshWK32eH
bl1xTHwGXCyvABu2pdrYCro+ilLvzfRYhUBM/ozD/uZ2AaZ4F17/IveqFHQGwzYp
LxrYl1C2Uiwpk1h2/A7ItQkYOgWgCp340YebZo1ZUQ0zjf53Oe6B4L5Gq2mxsldM
sqvKJW4V3zRVSUsaocsD/pgPNhH3I9AVqn2jGdxIAxxShQNRzTBH/PAoy8IenkMy
0Q5mTnSH6t+O0Iq+7GVNljLaYqqPev9nBUDBHuaC0TR0ioqGTBin3CMiBXVWr9mA
g9ZnF7gOe8a3I8/02jJHI2HazBIqW+5mxxzbKDVYx4jdHtBkOvK9ZGCY94Gldlw7
w3yuZObAEM9GJSbSwycVeo9K8xhDPqG6oAoJmktvlqdZIi3dIEyy7pjTVAjVlAcd
IpDHCR5kY0ejYa8ikwJamU95aGGjvHn8Eefxl5a4qUxsY/RVX4DCO2RADveL49MY
78egnHoJNwODDcO5IoHKkHm4DgGyUAk3WOSA/PuewvxE0p3Auq7q2NbGfvnH3Wxu
h4oorUdwLGUG2UpZEHQg83EeRI0SCqQnz9nSXyAyn2KVhCyiAGBh2qSzYIjaW4xa
Jpt8cB67JqXiDtLJOlgob+sdO5EOJ+wnssH/W5IwD8C+sxgJjYoc8K3Tc3lcb0kT
i7hL9nRJX9n9yXOH8twWy1ed4D/MJQOEatehks80wn21vGSJ7PpwujiG5AQUSh2M
msG9hhVOJ0Itndr/VV5PHtDbGvKXc3HxH0GXjSss8FawA1/tONsFGlpi9sIogGsQ
Sw4Xd3SVb7s5S5aKBcSHLAjF1GOjDS85hUsj3nSEUgzsCFp25y9+mvzFQ2jdNATU
2A3+FTBvoCzZ2oSGwkexSUB0eaFVslg8BP4Je78NuSze9s/0+aauUSVjBSK4pkfr
69ZF+i1yH/zqnvc8QrCBuXj8YkIJheJZaWUgsXprxK18pxS6ZYelhe1wKtyg9zCJ
CvKrPbDo2EJCIsYeVzafzMq1pZqa28hiftZgdogwT5ULt8el04CrLpcalAMn8wHe
Fp2mQB4vYgdUjB1wrUV7SuRbuV1JVmeBexheKrPmNcofqk0m8GqCgAjoIeWp1GsN
BRLD2rgqEq1bG4SXCjKyxOu0LQH0FH93BQTa0UF18u2CqtaxZfCU1WN3RJJY5Hji
v/Xd7YtnBcXuhL/iubVDWYtzWB6fShbFuqm6gikFBWlgMhau1yWEXclhCutHoJYP
QHRKlwycbPsLKWODjiuuceI6q3LOJVgu4fmg+r7RmeT8LNSS4xk+AS4kE/TxG/zr
LKhnGTc7Bs50qhvMYdZwd6GEyitW5I/agQZqAk+6RH62LyckkmQZ9BHS+xdj0xsF
0U9hEYq5a3P+rq6DngukcYRMIX3CxA5VbQoD561ry6ECNJt1zWSrX/DJidWA/MCh
l8x1/a787jA/ixPKmEnILGNzHwP/rPq8BCI4qWiXlHVsY7PcaoH8kkIms2Hvosfd
DzJvYP0fkMx+r1+voH3d60aXrKZ/xhZffxTFWs9CyQybKrmVx1lrrWyz4RlPYWsN
60G6cUbDrqIDAcvFoWcrhEk5eLRuO0yB4bw53t/d+a2Z04TjXp3ksTgxC5g6LCmT
2oI795vQG90Y8mtLU73NraPpAPz+N5Q3V1sfNchrniKGMeE8zW6CCfWWYjCE508P
gfGoqXZS/bWfk3oFhIdgte9TjPuVtoaZqFqePsf6Vzh85gpuHevxiD/J2G2WrzIs
NTSuZKyVyZNzskoeWvXB1geDKS/Qlsy29UMni72U5f0to4s8OHXhCmVJQb97gRPL
NtxMCOhvkmgetwRUozNUVFWciijfpY7E+CpYVw0WNIaFPkiBmIBaxiqM9AumcGPD
tANGnsB/ZjWqjwHUNSYqhu7rHmDygmd9uMbQzEMe/RwwtZEbO0KZyB1k5E5xEosH
x+fuwYrFyPINzSqUDjkX9eQr9b3waerbRCyoi2ctLNqUUcqNhVECPpN4m3z74sUi
lPkFQHwpaSVKzp58gdIGmnPu1W3gSblYtehupnpiDiXPCYQkXaIyehrbeWe6RvvU
hVRnXcdZ+X1dxXEI7oqK35Nl6d6fV6ExdZywY59yiVBSKC5DK/HYS7Yya9InfCWx
N1DsDEJWlsGbL7thsdtPEDAySP9LOx9n0g8d5+UvsIgYVvxUYn8R6tJcuZ5gWzOo
ryFXxpfc+GGygvcA0Be56ZKE3MkV1SmZkYpLh56WsJXfPFrjNeIY80sxoYWYWfS6
Gq4fFujPRKcTSY62bs/V5pP6i/dxQNsUb04mtMkCqN8nszdnqaOEA/zHHCMk2P1u
RAV9PT9L6zQr4OmxxPC9DlvLVXL/WxGFPP34NHk3cRnJW/pitfN9WKP5qVckD0yo
gTM2FohmFsjaHr4iY1dVYMHykYF0whQDoqu5gyg0BJhQ/IrAfuIUxfyGS9YVeaMt
d5j/mi/HUeHiykXW4c3kJHQTjwXHAVFHMup97igsG4UTueSH6O49xSDazdvn9izh
sTYuTX5VtnJEzQhmCvjS1ruO8mf4eSZcJ5MDioIDDymeaVP6ZhSElwNlG4qinnii
yBHBksZkRxBdmO8AVehaBwlTTDZWSOsRsueIBdtEDqKjdV8tu7W4gHOEb+tiSuy4
tadEgVRExHv51F2jnpkOIzi6l80PEEH8FR9Y+rqlRL6O3dkFPAl9otjRZ9KJGJC8
CIYcx44I0hgHMrIqeehlbhirJJ8C9qnSYqJt3JlUxVWOaBjDPHLea0oUH9tOLhIF
RV60QSOu/uioTfgu3vRhBlK6DkKEWEhyIYXNOvS27RSKWjqEibZkecVPnp0GY54y
aigKgOxmOZjLMo6Gtgjek49OLkOMJPmaqeec3pAxBHiYFGt4e0xzpxycdyovK9cq
Q0xF1Uv0lyb0506lu5P/2W8FBekyVVE1dsbMrupjvZjID9U7y+2swW7nAato0jb3
htMG/d/RwrPjHIceI3P7Vjs1hGV8LN64JZtJap4hk1WXHsn2L4sem883BRs4P+qj
SAWQQumidY0vLDKPogXF7EBfVfI1DDQDRk9LHwvIeByoBaO0eLQvdJnJT/iHIKH/
kZkxNt2sQODy5j3CMLx8wwQEc2A5nRhZdxTkfZNqIp1f3yVL/Br+YGaR9fx7Lghx
PnCGeTB/3kdCc8jWwwbl/ovhm7xX2dAUC+236D3arJGRBb7tw3PS7SGyu+1lj4fI
ICBS5hQyHzdCyZZZRAVFG/7ZFIeaOl24v+wmnxmBROlK6ZoJaEKnVYc+96xq7evr
7hRgsQq2MQzvejUh3zdOoqqxgdJFzrjVgJiPfnmM60Gi2AyjPkNTQ88UWJhRUT75
u37aOQRyNvlPT1J5Fsg7fR6tWxnPOUz3gVW8zZ1WHpjJ1nrhFqJCCATFeGv9/qvp
g5OfFp+4at/OmQIBJm+7KmN+tsIKrCnu4PkohCTH2qoETyRQahVhPm1RohhEJs0r
EZLEHOY16+nWH15EzsRoIhNrnyqG5TjRGq5l93Ekk3+4AtbcP3xorznhirgjQ4r9
Bfhs519xip/zhfG6vJ4S8BF3qGAvDzxc5Nn7mrYjcFrdwGZbKw3HNUCsHf6IgNDC
kyO43VzlrBd4u81f3QF8BCfImRDZRcTNWpEj6bWGvqtuu8fadz/zeAxjdyeIOktQ
SMduU4fq7faMpYTuh/9yN9Zhe9z7T8RswCF/8KGRbbCxfDQgJ8JFt5+bD7JdCLq6
oCOXQ+WgPEtoxm3OzG24kSY0uamnj8zOkU6aKorUPZE3gYhOiu8ux87R0Vfx5zNI
kgaRV3hlwOSBlLpSV/9BYku/FSQQXIz2VF5zFJRLCNypSSUeysX0GgnWglJ4GnNA
/I/M8jepgJteHR+Hr3QBRP/DuKZPhjeJT8cb6lMoDRjcoVT7BjwMWmDveWG8fcCW
jFJ929N6p5NAQi4++IfPA2Shan/Q+NqEQvTL35zdmk6UNQL7BaEmA4h9ebgBckAZ
CPl1MVTAOOaD3NoagyPNJaSBE0pMnv3ImRv3FrVTpzTvPInSqdFs9z1is0ycUgPu
omeDdzPpTINqIgj5WjgiN3Om/ES2gv95TH61SaqSV+qAfvV66G5V2rIFx38gwIRk
gix4OziPgvgGkXq1o/0GsmrrVHlg+ajtmBm+EVrOY98LVFNt0/MYyhkdGn8Q2akX
y6Ioz7vGHYWCks5TiuaSKYA2zPoQ7Vw7MCIVUBqotM7vss9AopGILSyINHZPeX8E
+T/L6vbkG3UpyGfRYqSIqn8UZi+4t3/iviflo/XUtuv/eIjlm5grTWzD69IWVIaW
WdCEvXve9nHSVY7M/GN0MqW+49IrFAXp6OI0d0kZxV+TjcX4bMIGJWdxsl1BEeij
qmp8MDEaXed2kvabENNRmuguJoPt8ywpePLnOt9kTIQAUej+3XeYkdCEIQJLd2t1
0IBnH1P8FwstGRGy5UKfQzmKGeRPhvZoyTnNUTTA8Vzqg5vVXyj36cBTcDaLvneH
Nv1K5Gqs1TFQJl1556N78ORLm9KrVTPqGbq17K8zaDXRxHhejZvuQx3cIa7WKWGE
Aj/qRySucax+dj4daXZ4c2HbeAznz2bhG1WeeXpoYY1gvL6wrlvsgz/vzp6+9weg
sTxCmnVbKtLOCTsxJo0HD2HF6qCyOEr5UEJosL09PZ8kCljla8t+AM7g97dI+zcu
0k1ZYE7xnFz6jbT/4o5lPe4sp/le53PmciLsyS0IIYKpKcZoCJwT03FA7Rn2jIO5
HckReLWRHHFgGiILH4VEkgvK3sPuuJpS2rqq5qkB8z5GX0yfR+NIHupPUZZBRbUN
0sQia56BQxGTNOzVepNVsIUp5jAh2B2WNN6vdmxfCSeyet0sILbdqMZ+7ptSHiqc
/9gSLjzfwteWsGT7iyd8cN0IHWb2zQ8VcxxNU+g5ujTjRcV7BVVaJnIIfG1pCmWD
lNKujqwYlF46AQuBqrkFBBAQRHFxil1I3aO0WvuuzdDUzYNjtmeVhztUumw/Q+cl
rHKhiK4IeifunprY0QX7TdEg002QHWUYVJH8SEK5l3dTrwawykgHToKtViJAqRJk
P+dkHty81GbJYNrQNIrUh4iNu0RMIUJ+yTYTrkwK4qztE4hINGN4H6ZlD/hxH6HX
esmxBSzR//tmsAeTULOjo5+g26WcVGRfxgYxyQjZl3s/QZ8B1jzCeOK1TTEzjJiz
TvDWAQPjl6lEmC9n4SO4uI1b95S0eB1qAWoj0VrxMI91hwQmafne08cIP3IP88kJ
5+eNn2filJghcvd0UROak5aMmbTi9h0y7lLDypAgtPqv8R8D0hQOCFst6pGy92T6
LjDN+bCpI1CRwju8CbOBflZME9d3rqtmpWnyFCkV5QKuAKMAlGKaXMeMRApqZRFW
y8Z6bLMW0mnLMZYUXU8MYo9v6ex7ipkY9Pj+vgudVmePaj1uGhBN32CrM5jKlAmi
y7XCv+a3JYuEw4yjud0b81NcYGKFnbgxu5uav5e7Bdf7knu3OJZvKqpxydQKQJF5
IQyhQ3BfZrbfp0w8Q80yCgpf2RKfJcSmF3Oda7p71Ua6atDU9op99KpXiXxXMHIz
TE4KmMKEy0C/XOXE+l13jkvZfVyKZ40+90R01FCG//62/GD/W0k9ynAXjsIyOp8X
PUSSHCEt5IsCQLrf1KcqBaIa2wzVaoRczf1MF4jO429wQKyZEWYLAFsTNwykGXe5
sE6b9YuKoKoQayIXWvNrpt16LVPpmOv5dFWWSyr0zmfNUjqevN7hrIw6dX0zdHSK
TOdGdFUekJ2cjsMaotpSHTDo2payaZSl0SIe6Ja2lMm5GPUDYOhdHX65qGXyoVm6
UluUkySg+/kdLXuXgEvTc213cPQoPHgu7rN9KpyxAVA5fjROjQRyCRinU8Ka+JQB
3YiTjVXQiXcxsVlMEiftN+YcQ72fWAjEZzrR1h4Lxsklg0YcUYPGDUryoCdNBiMq
1uV4ZPpp5pnJqVfILy28gDzItG60RiBUFF4ffZfU76wixExwYG9J6minB6Me4Kgs
GIcvkWYjN7NuhagrY6ah/6kANmYfX0b+DTrFCHyu1Jibm3/laAd+lhLXWCNJ1sGO
/p+l5GoSK/iqqRWxd3OT3bGU7sRCV5+iLcXmeCn6w0zV2zf941qkcjWvMS/uspyb
DxwjzcO5C9QxzO3dO0coN4z1wn15ApmCfUKv8adZyeOEVVvVq1ADcrH/TbC1QxT4
3HplnvvHG1d9yfRBwEBEjsKEKaV9BCdUAALpXv/+RM8zlrElnb9FZgGA5TvwZslC
4DEsZe7DEJYONLtaXR531h9aerXcy6D7DAJ9DG+84A0TJ075h6r20fsokEMzJE9n
nlm8lbuf5Me9NGX/nMK2PCHWUtq2klt7T+d3f5QxFx+KPbRzewePmigrMlaZtd83
uEVEfyJ2VtUGB4XZAfEZxupI27zL5sxNIQbP8CUtZXrl85LKtilGApcane6vS6V7
+7l+4OB7IlMeRp+T+yETWNz/7IUuwH4hRT2TDoGzVDkjIAy7FNpSIAUZ2rRDS71P
uOgtlJb4KSAJ/oLRGjsAzCR+B3T3EIBhUoUfFVZQgYRFhEHlvu87uClyjjX8GJSt
rV1VGvVBTAxBoioa2pAByl7hTqqFb1VGKyKEK6zNokUzUdPjbE5H44ENWjQda7tA
PKaIreQ+2yQC31/bg0AWqKJNb5tXd12gpOWQcFrkXT1fwbfog+UzvAsG6r9/cS2W
eYdeBApoHJ2nagXz1GdcXi6lsrDIeWJLANc15FgttJTnx2mTpb9+qQgJrvJa4UnK
k35mUXMnhjVhBMxIm+lh5YBnlnV6r1UtPC7+8I9myoX+A8sg/6trTEkGj24WAHGJ
C4SeEduGInaEvu7KIKE08SbCvXSyGdVErszEQhwbnF+YHtVfKcsRRIWDAPU9PMYL
LsFKSSx+g2HE+94qNEJ3me9p+g/V0z1H862s7pQ6dCWMxIIznIOEA5zFtgiUDMoZ
yw2rMHG3KPRNqlLLx27S34f6NBnTxuO9QLiKpr9n6dCZ7oOa8KJm2Zia1pkRULpk
JPG8kFQ6ZfW89xuQCS9nRfnccTqnyoVeZpj6hpzI6xPVAuiEs6WSoJD58tXHOcaj
VsE7HGhHR/Rahw8mCwIdTfitryQG5Jm7TYTNvMiIgqkybGWgNFa1nekgRcAlquH4
N8VDEehuQS6+9c9O6668g80EjoTEqSyJGBNBKlQNBVgqG4Ro1wMPp5eH9FmEU2Pv
T4B5maa/fcaqNxphucYbWR7jIcXhAbHLC5SiYWFfZlmYaX893U1ovpc6qUfIOoMs
4tppK6ceSOmplqMJHWgnb6MzbMBIzmOT22bLNHTGyvEfkkeRAtnD4tCUP3ls/9TF
9cMkWcSAbnCHw5IwDHiA70tQM5T99bgXJx3L/DXjXTv3nhmsxVpCBdDlMzOcEBaX
2cyZxwZszvrhb0xS53EEJGx41D90/dnm07vhG9qCEW4aiqrWguZMxZL0h7J/XW+V
+q5yEJB/DyBmCop+s7TtHKh93oiagLT1Gj+NQGbu0NV1glq/qexmCzQT5tiSOhbV
zaQceIPvKq8xTtEPIV/dMbnT6OlRFFhL5zORcwReSPSpWhypEVcoxJ+AWf1ZcAIs
95WUNTMuHZQi0HgYE7hgIBHZYZg7i80wxKxJ0lFgHbdtg0tNO8c/PGe/N95hgEvH
oPeyGJfV7tql1FPTIMA5G5MHBpybB+Ym9VPlBEZKwGkZZceSS8GkLaKxGc/awcCZ
oi3JM3OuXOE6E9QfJoSBYPPywTc4xUKo3ajJyLRtNtLh7M5LltBs0iJ4F9iUDyFV
F+szW1pQnAC7fCMHKeKpmW6u6HLnbdEqzMkccYPc483/D6gQxGl4eOVZxbKe4c26
XTSdeuier1zRX6JKvjZj2fen6VzW3UdSBzp7ujmfNXwzqKqeZIAwNn846D5+KYk5
Y8nYiujK5BQaJNTlSxTRU1gMdPM+MUe055ay4JQ4V7yufCVAQguIs8dZWF3a2YS5
xx8pL5ZdMlW8DKlNfNelmUNcA4ZuIQqyB05pVsuJHs+LVDZcngsbqgFG9grZ4BJ1
4Pt9O1bRyAQzKFlBwbvu8azFimfoahwEF28lGLTNb9KqgED15fe7j0ZVWry8L8YW
iJv3c6KdNbc2a2toSsNNOKWy5RCJYYgjGfyP5oCqxL3pX+1bgcyOpPILaElbVZrm
a/8PWNUEV3/wfj1LKCe/62NuIvQkiFPG8jdawLghBOSaGTit3eUvlbV5LgEPEfR0
E1WIBHYXYKejdwllk7SbVX9nDvFJUIWKg6qGjFrsdFrj5eRHqHQXR1I6eHUg+EBO
Bx75QAiJ0lfgHHRXxhTwbA5bf/18xU3NxCay7fz1XWPK8AX4zuPN48goIbpWdXAq
FWndJJfQdctS+JcGASplspyF62TWIdyD8pq5WRw3kvngqOzfTx8IdXb7v9JQHfZI
1bDCZmRx7wV7jhqXQ2cnZ9OvCEJ7Qu0LGUlLr2OSLbhNPAMOiYBZFkY9jzr6vgYu
x/ao4eTeF9UYUVDUjXfjmwTvzEQBBSf4IPYC8TnLtTGgNX8J1yBoy1PPTn0TbE2+
2diW5YKFPcAHgR78epdHojMtkELWtqjTr40iiU2WuJYbi81onekbs1DpCQWDR+uk
N0GCyxYfVoq2Z6vgMcqFxc+by/6bBghMV/+aLQrLcJNVIkvyCA/HCQQZR8mvtmJs
r+m6A/95uz1PN7vGtxvNwkKI2qUqQeguNPb1TsUXN6+xbYaMupMppkqv4B9vOAwz
xV2gnbWfEn7afF0HHA+RgYi1n0MKgex31KVnuBzbULsxq708JqJTCJtJRGb8AE43
6q3Qq7U8oYdQxQGiP/2g3iLvIk9U6usqqOKgFqArfSGyXseBUu2289Uyde0Urlau
lEBRemtytzceXBiLfuORo/Th1X4Xmz+coM4UmFj4ZmD8Z7z2zOzQ6VkJ6Qt7JFF1
Nxm6xbLV48oNeoi+t9lqjppWomlgsjg9ShdYKzeDrsBfktZtubJqG6xp6EwJh23q
Amc2V8VDxQVFUTn3jLVlNmojhb/mLRguqXCJAPvNcwZT1QD53RO2dWEyaGtPR6dz
5SAPAWhpE7/G2TOMYiM27AmsGTQoUN68H86H/9OBZzYReLJ8VvNuKDWXQZowDJtw
TXRInKu0kOZaj71XVduRZA4YOCH7l7s9d6yjZk78oDrZryKLsHipLLd42gDya4mu
jC+NG8gZfmqI/43wvBdK2eNHWWm2QhjgosAw27z2j1MJkUOFCgMvBtBiAf3Q1xHi
L093Jjx5oi2AbgyT5TAl+nIcgUefjyGujjI/MZJKfthqbftF7gewQbK7FsdnRBU5
co5Z/g9M8BqaV8cDk5PAfYDDkXxgBE0e+eJahlyMSXbqS+wm21bpfEAh5FAgEJE3
qpqnn4jpEf/L11JIRtoWSvo6fNf1BqQ7gCXfic+uAReSYz2Pr2/caBPXl9GRA7kM
LpDDqM8kV0QCbbDesigEh1oU51nuQd9oZOnkdXlQPwdpodWOycWAzs8uaUL7OhIv
3G0Mz6thDL91YEpe6e7sLI9x4HXYj6nOezyGEAYDBcHii1vYg5F15bGGAZHQMPQD
9GnIT1LaefSsjdKns9Q+dk7MlBFMn7Xa7BcplAjWvW3DLA0LZpCbVeTtI/ZljIll
SXGExz1BffsaeRplA3F+OZ+JbsnndMrWiTnY5Of+3YagBS66XVIxn8esnDA54fMN
/2Q2y7EoeNKX8ZPGbkbQRjuAMh0vYcF2vVzzx1r1rBykS+EJw1GGz9XKSxRQpZsB
TCVhPxXu+QocCCCPkZCSuRYHRzJJTDJh0nJSYru2boh4O9zYItYagtaOEKQV7deo
82OqqraW0uT1I81aUGsaPSptbKDuTLwz0jrywQZ4riS4CIe2HtDifk0R/P2EFrBp
a8+FodlKxDJcRNxuSYubpWP25tuy+YmV3m9rnEtUZ9Wv9iuXOFgMESRdl1/rXE7h
2nXTrRDgQEXGd7KXl7lc3BKNVVAApVMlE/t0Fpk4CD+U4aiVRIZ1wCMtG/ExVP+f
edsT+VeWbpqCt2GY6ph7q1MJbDbTq4piAz27voALn3Iu6oRSY0HY72kmSThPBmLe
dM7la4eHIsq9PC9tefJS4PuzdiB8DaZiXJ0Sj03voDwBKIizZETGUDmnK9mjeoGK
JF2IhiY6zF5shpzkeVEK+lnRCqEdmSf9+qnYmmWsYZSLgt/MtlJQF+l3fWJgqV1u
XnqrCsBaEm8lNSFJSCtkoxxFZetbStsxF9qxBWf55su8PgkYMksw54SlM11uAYHu
qpZkKL41NK+O5VeoXVuEsTyXX6f0hNAVOlMxn4uShLhH7KHN4MEaGhXq0mdJkPoZ
Fqaqz1CHH8cn7NoEluO4YEaTpFsm1W4nNUNr4Z2P5qL+Gv3RN3nj7SBdvXzPJU6T
neQMM2YwvuSiEkV51/WWhJF3KRbukmQRNnM/od08QjrV0iHSWwE4BpFbghKrwAcu
UUds1Q8NDNiIB03E0tre5ofMb37ubTtgOyEHCWWZ93hoMKkWDEMgLrHHAULK3xmR
Xc2KxOH62kVb8OQT3z5wwjsOgTlF5HW/eFYTE0vilcEssiFH92DHV0LDxmqi95tk
2ytq3gIFjrDThZQqDt3+THWeHC3g7Fq7jXnq2hCnwtF7cSLP8FkfRsygMxc1gGEJ
JPjW3JcigrMfrSQdJOKRebsCOua3YE9tHFylYpr2H6E/FyGmvd+nnypkVfRGxaKa
N5Srh1Fkxr/tIm1G8l/kMVRQ4otKNsTxaSe5gSadkEZ23mpMigRiZZ70H9m77Q6+
piL9gZyRqxR46ZQ88MIA+dh3NAPRy6R8+XC03vaEeqy2A8gm3JWA4ndMnM0aJg2E
A1/qrPXvollVzBjJLCMpF40vLNcZFn9b+0p/eoSg6CnwjQ8GTXmdEG3pzuysIcw2
PlkulsH/+g4ytDFFQkzMxjV//wSWqEzHxbBp+FR5I1Bc+xvFMOedfIDkqLSnaAT8
EnQEMUsX49pEA5FBs3V931R42mn+7YfpEONrvLQLYbY2jwSRGVQuv0JU+6D2JrIG
XETOsWM8XKsDwRxWAEjlrTWraJAmgn7i6Ks7T54Rgex2rOUgTuWWkMYB53yp31gF
tkVK4kiMRdV06B+KcFlriW0+41Od7Qehb6fV0F6jgdhUY71PpcAPym98lqP8tnZ5
rI4uvkpVOghsUpz8HcdU2sp64aGEfHJ2Hmmc24EykRBGZ9mdEkMKkHV1Sxmwecj2
yGKH5G7ltZ7wzAfDo/Z+PzObOPEiDFbq6RcWmFRN4ScJ/ap07CsYA28Gik7Kvzc+
a2oXPwo1Rwms8XRXbInfDrne58SQ+HJVkJKWWN288ah/FmyzyDFKfzDzpDMOiaAX
O75HEmp9znM6IJk1P/rzjeFY3pwASrzO4SX0uzJH59SNHs/f2ONkBiwiTwBKijoo
AbRaFkDjf6jinAzX6c9qbk5GK580CGIK9XDPISwZDyd261SxsWtKkr1lHNdB5TLJ
hzr1XwDTlkrQxR83or4bDE8GNMKtEs+hEGLoUnhqbTUcwic9IKzyK4YC/PrvUPPz
/QjXq96WkyCm/CqkgdaAe7HqxpZpd5jd9onFovZ+bES/abQQFj0etU/XI1KdM/jx
jzo/ttrA4mSRaJVXiIPTGLsL40qdkMYvVVTzMHjnq3IgDYQXIl0CzzBg9Owa4zb+
YKVECi0xOfeFGPgQXUPmzXCtNjrX4Yz6V36M5YY70sPXHuO8Yv4MJ0wX4QT9r1jA
CBbPQ2W9SaS5/inz0KG2y7Gxs1SneFe2cLUD/75cJU13OKVkJJ2bFVuXMUNJFfRV
LUOm442SWf3nTgcr6kDoV75RZylf9EYIuunB325Ft9oax2U+vj/LZQxU6rP3/r5X
tf2kgwOZWMEaal9iTEa6KoyUaFTYCHGSzk0I7hqsRunDf9WvO4hZhqX96RCaV30i
M5TR5dMqVeUCdqkipVyYV56ujikDB035/Buq3NyIByi3Xz1xZxq0feIlewBGYZO3
cWHMyE0rA04pKyQt7XG7M9QEP0rdcYVgCn/xQEgCdYb7aMENHLNJXgk8veuHkc2T
6VRrFp+2vBR54Jbfrah88JVZaR+JZ1Q6ESKmKwt3N+IEAyKiEzgsxiBuRcbPNEiG
6/Uk85u83GcSdXHVYBYxRygF4S/DFJM87DPInOfzAA3EWeFjm8Trm3msIA+m2OII
qRQRnVQ0GtQy5A6rAnGCLNeJXi6ofk2Ebh9vsGu5ts1EbpnPaBE3wbhFaZujR8UW
dIh+6L3R+oDPpIvO4hi02amFS90e4ElM+8AMBxXUMiWW6kXWecfcqd/J8AEAumkz
6HdhN6py9idkAg1KOFwjAIGrrFNnfRSxZD748Rg4jmf4SqD64coAfwA8iWYspG1V
B5RePdASsCxFPSE93usY+TNTIgwniU0+/mUUFwLhDtQ4bq8cBC1eMG0BQLxmyNYc
/jtR8QxFUljrZLb8PI0vQhHrlWTZCLRAUP0PTf30PGsZHtrJzwtAjegDvunZ9zuO
XnXx625wW6mFqJsgM1Tb6zjcyogftdP8ZgsY1Id8uFI5OkxjtRl+Mxg90Q03TALb
IaG3JJbeUJZ1c6F8lzn7mhV8xrdKbq60JiamJF1/C9CHs8jxSMdctir34vmRfhGS
s4puxl5K0EcyqcFyj04EoUfVIwaMuV+iOv7aZrpz3coYTUziKNH40P3nTO32cpMl
2LQ5w+6keSbslYh4+dHD/dVvFP9J+AUL97I1ssMY4MVDBHeTi+HS/hceNJW8E9w2
SmipKfA0wrrmL2xd8Jk6qd9D3NeJrKsanVawWazzSycfoOJ63aIZsZDUCNVIWFip
m6T/RU6dS4LbEAPOLILLu60MFecwaQ6/DV+4k6OzDRdk82o9hkgUOllgVyCn79oz
KSREvEa6jFSE4h2XJvgGvC/7qm4+XrJ6NOLbCKlosT+FzaY0VHOd05DKLOLcDipn
SNkgRQft2m1tYoEex5rfsVshEl5OcmYQlZ0pWquMJFMKhB6riFxeWMQXalaR1lHB
ef8coL0MSdMoTlq6iHp7Bb3KjM1Nkko7ci6xz7kWDJZxaR9DXnwxcd8EzzUuaqF4
oXPxdLFlE2WIE/jOGaatCQHBdFsMwyE4/uyHS3X8J9zYRF5vsEIx2e+LQI6XUTXd
j2AZfC43wkbDqNSHZFEZ6TkIvvYZ2PKiH0bbfmAvuPV9pmKR2VFVtYSbBvi87rMf
gSRRtcjEMQK8UBnxQSdwlHj/mtiEo87MrxUmXIG0B2OuT6lXGQf2sXM0W3zGEVc+
tQiFTRc+iRw2ioudatqFOx4qsaRaZqmMTau22totcUwvG7sGev1s6J0qgE4GngpY
G16mFVV2zjNnv2nk2mu5Uqr1U7kW9pKqpi++idRMHxbOzdckqeJicU4bzXJykV02
y2MUH/mb9CIRvtJgSkQoI2fO65qAX7DEnAN+v+doKVgxUjkGRO9v4HxL1wjoOhIQ
nU7X7W5jVyEO1TQrSCff8xLxWjmoLaFrXWYKGQA6ILAGgP1+BsAWAAfqhdwl1ZMp
JC5iX2AhJQ0sqjYWm8QqIgwJMz3IHNs9oYUmn1JSNZVlLD8XZ4OSubJgY7k81Ywk
9ElV5Qg3ufNTFfD3KAnwYhjSxJqNYfJWRRqGLwV4V4LIXmT2HF+eDEkQFzS2dZf9
OqVNuOlFo4a2EhtCmLxb6ViVHSf81Q3U8ZzN1z7CTDpwcVDki9fbjHWN2cu97isF
n8n843CzpOK2ZDWmOJXEOfQSi+MlHn2xV4Hf3bfB4XJlvbqv8CD7Yhiw+0IALd7t
uPKPh/rAibVNluac6nMlfS1OcLZvFWcqzvDFcbnM1ehOo1Z+SF9x3nu3eOXUY79D
gzalGeXvYOSX0Ik+Q1Npqc0tuz1h9+NygiCoTdzcxcBcKBgPzNmtdtsi1quuFy8x
Fb3frNtEHW0MQocgCuiRx8sPjTIlk6qYCuQ0l6RGahUa4zjh2wMkLXIQ/69c1jas
E6EqN1AvI9ddJ2nlmYZew/t8dMVNw1/KhIJczNm+WyoZWe1sD3sG3IF8z128LQzb
GV4GtqWA1Nn5Md/rirqgSMjfkiQ6qxscljQH0gfn6ETko5cHIR/ZFFBbR06Z1zdK
qJpKfigCHbkC7J2z4HEBDckVZELr/c8YOlcY1+4ZOQedegcEiPv2C5oWdbB69SKR
WNAzi6yxjMli/axfbrxhRF/rG446wgNyDe2unyaBy+BP9IpDPiTo0t7w+p3Gr9TE
xhVIxRxO9ZI/IONn8JbeCn946Agf75fVYWyE2+levva0t/Zzvy800q6JfP953Wpi
vy/Ln3XUVZF9020D5g9KRiiTPYhmMKWvl+EiNzZUiVGFV57BH5qDuXmdBqbWXAdZ
g5uPROazS7tJl0LYb9GS4f6jhuUxksZfcb2rHN3HWLYP5HJVUd4AlFt8ulQnbFlm
RC4LPOOH9SjJnqXikTuc1TgdSSBuEikjFBDMjWFvdTG9Gyql25cifHQw5dXpTMN/
IAf8tTAwsa3MgajnXHpG+Bwwgkg2VGcMUVFNZFwoiSbwPT5PY1aEAtX4GPaUVtfI
FyyIluaUmIlA/XtNz7ivEW7GFFImiOTHpCLrG9iQjTs+UWroNtwcGdp2XI3woRYN
zCgwfolPymuhLCORNB1saFRtDUEhFDqquyRiJd8qUuC4N71tXEZ1IkQf+oFm17d0
ATMCrSCtMl3qPmUA1OCShU0EijXv7PXW02uq3CSRoTKN9cSc8dsJXfHJNgxqLKVm
y/GisoOyZtiKh8w4bZ7XMY5/pwjrgC0p/rsiUfR+GJjTm5xGrZ3lN/fsTfVdG/Ch
tPVmXNb9I5r9Y/3bYMinzJO374h29c/ieEsT7hzFAaaLbexG+s+qA7YmeVCykNS0
V7d2tmZNjoyenECY+jE+Z458vh+R8WyjEdVDQNZPpJwLkNrY71dfu5dmb70AyhLX
Mjb3GtXvT0q9y6pdWggphmsUgAn8u32AwgOXAvJDtzC0iqRU52cI1oRX6dpRHkGd
IWkf0e5YMoKZ6LyFyIRcnVg3bxTK0JcKirI9f5nkpWa8+sVYJpDHLRNUfbN/Z6LC
XM1pldxv4J7KP8WO56fvQCfONISY6MY+jV4DWHE3ueDTk4nSa19avLFY0pa7Xq/Z
mEfg/Lmx43yBTKb3rqOFFdlH1txwmJZNxW3GALF/5DsD13+WmT0YelsX38PMrJiF
eM2xpYjUXPvpU73Pf+RzsGaTHXHoGM1Hy4uSqcdTcVyIGTP2rBHkiZfVLOjNfNHS
sY5xmp1i2FPFEBG6HiJop98btl+K0Px8OOAroaSTvbJa9Jm8UPgtdB1suBpEwIER
o4z/g6rGUFjCJ+rExuW2fbJ9PokrLenK2tJXDlwmeaC2mEEnuRUJ4xMmNu9tuLC7
6wpXBkqGkT7e+r5KqCe49uA19afl8UsNUrH+/5dsgIPFUIlV8ixWdeDW5F/iityG
uT06qF+96rGbCAVMlRDz4RCIgk7zNU/2Y+RXaurxnkRvm5q5QDELTlUQ/BGWUIfi
3L5gqXcUuvyds6UuwdJYQUsJPNke0kZWvvDAtWpeEzBkqUCKSL5elu1gjIwUNscH
Pzs81Jm9mEpKG0FwmpJJiwexvkpqgksy86a9S+B4JCnGZIInyfm/JyPn1IU1sC1i
V4z/j5cjtxeeFKeZfnQk1xXmlMFEuEgvb/a+1FUNrSpmi5Q+vUbbJ2I20VqYtUju
T3bt/iSsCGn8X8BBCWwoO5C7ueZSX2u8VZ5HZrQ0gaALT01CRoWMP8inhUhDWs2j
cmjFmmScgrwiYQl4zuFCYeK1ucclBVNmRRanzr4IhR9Vhg+Dq8vghh2ZyrYU1jxe
2QTNUayzWkW4kNihpUwIsizaZ0Yvl8WCaEZms4mniVICT2PkrZ+b+iLyrYRFOrwt
jHChZoytEaoGWwnILnuanFk11V6tAqW442WRN0GIGuvZ0OkSiqjBjsFawLG/dNsY
d5rC1SGyMluuaDZIbQu9vHjfnk9M+i2tQQRgispDB82fWcNzm3rjsAp9gamTjhW6
4bEkGGp1y0vjRWVAx5EataLjMN8PMdXO/uF1j+eWV8vrDk/OMm6tV7xMvJeWbLgf
j9JpzpejDOResi8iw8Uv9r7lcP+G/cmwJPois6e9pL4MpvanAShLdu1UAMQZ+zLy
umZZjlgWNnuK8wlxquLaifSfb8QKuIgBLiUNcJkeURQX2WtDnCuBQFIBhPTfJNIG
Iy7WKkDt4DdOKVB4ENbk002XZ+NBo8f6DV+aGCIRWomSDuIdVwZ1Er3xZE3acaFr
sP2X2NbZcAo3KcCOkMdpIuVBUBbXzb3kB2bOUWB4xWUD6DioE+6YXbRLlcgETGHa
z+/2VVbarD4cvjY+KmhIsrZtCdDwO2u2ao6OuPqmLLaBfaWDqYlVTZ5LvuF6/r3+
uG1/b+xb5ZIsYipTBseWCi6qALlbqVCkODAJ0BDw8zjWHzHIVcBRvJPeqRJNBnLl
YRLco4yHcT82Pz11J6x7rjoJND9DCNQYJsPm/TPCCYRCkyGUpoqtmT0UyZ6M0j5r
eEJUtHpAKyrmnQfZyjcD35760chjUBR9F4pijqOETswS7pvHgyZxZaFckBLQbKJC
BMN/6CGbnurlqUZg7+JRM1E7x21iZo696CVEjNbopUzY2S7i1dIDjJFq4O2Qmy80
2++U5Q9lotXjq6ovzzmqxY3G7Xj6GxDr+jgNP02HYbWFHpGwtX4IdMKNOTFjePM9
j6LENZ4EAhIGkGuprA9jukDW7p+u5VX0uQo1DOadszk38cnWTs8SC9M1GmOmA+bv
2Wx00ODpcRjUzTQ6r9/Lm77r7CAjbYbQajIAZOP1IrGsDbr0FGmMKqGwISimF0Rj
JFjfJXlC5X4e+UAAAM1q1X5kdvLZpK6jwQXytnEdqDyWCC3xkh8FRdPN8a57n7eQ
oH4yjeW1w+bZzSrJ5yPN5obdxiFJCN63qKuibf086l2IAJtmOAYz7HRGWfATEEeL
3iX+rcD7ET67u8Amg9+VY87kuJCG9JU1B3BJuixKy5Mput6n/okfJpzzth6SFgqg
dKOqFpAhg3dQO4LJK70kBhW8CFBD/10w6f4/BXmwAFIH1WgjrLA3m/+GIHotbr99
k53wrr/ngxtZB7O6zITWtsyQ0/1I+PiHmsQ0A3H8h/7BvYsBCV/5tzE4nx/huXTp
mxNcIcVVxzvF6tOzfPCMaP5dJguyMadd4Fd+ngivJDmq2MAYb1OnQ9xShkzT161X
O8jCMvIceF8rIDr0v05ju4ecQJmlgEwAitWETQZWzR2l3zi+BDGYAWcoNYCf67UF
1C6B6fEI9jUGm1ZqBv35cHNMb5mPstkTS/dyzdvkRwTwE6KFMMmeQkJMbKqEMoQb
MHQ0GqVMtq2l6DEwysXaS08nUZo+O+/P6LKYDwzREr9Ir/6uDfy/Uq9WH4AP9y2H
iextQJLHLs/ulrvfcr8OTf/j1r+L32wqiN9edf35h7zy/b+VKAVPup3NPqW+icHN
Z32mUi+PwYi9eY5NI7Vg9jteCCWAgWyvfcu9tz/ErZDvz4yyZ0XD2k5xK5uP+Gur
4miM3bEU0mTMW3F/9Y6iNxJNG9bJWml1cwd5PxdzP9G7P7OGcORiDNWkzyrlwONQ
vAnVJQMgWYdkqSJ3bVCVRGWSBBjPHwFKVH7BiKoammG7nVSDB4veuli7zrDM83Q9
yu5A7pzDWdHWSQL7ChnqvaseAAQAjWOkL9Cd1YVijYzAv/VrrtNINu7m3TXgl1YP
uuwtsGAW9tZhapayDt464z2S9+ebfP/8RCdQIA3OrzgsLaAy+xKicNmtRjLD4TtL
FgHFeac/FR8x6D9Mnm694jjiYGBserbJpBzHee6JcQBDJY1WLP+pULNMnZlw+/Gt
WAc7nP8fGKymAgaOuKzauQIer3IMOjAeb0quVM6hcWitM4aFL/NirBOxWE11T+a5
ijdWVsROXz1SIcwSaWrl4x8oIeo8oWI9zs4CQPLcI4bx56ApCtki8Wz8N4twH8WE
4KEMzrejOmoFsj5Pwy/OyxvTEnbnoNlg2an+jhQTJEJ1TgHz9a0oVuYY74o0KEtl
x/NJ6UgNYhKEQ8nrrPlcyI+gRU9n3wHmK+75VcV92W7y+vC/4O3UfWzBFSFq1HaY
mDZxARAmb1f7SUFEdCRSWSidMBtaU5VhVBzOO/p9wj9m1pzhuwJSylUBmwh+Ur0e
fuVAlkAV1oxBkzYtrwn7P5U6zhWX5H6VMDiHL/I3Xt0TgK5sEP1l101lnnbD5zkc
/ruVHRPBnzO3dx5V4GvYm799vgDvr+MlO/H6z3nYMJ9HqhQQqFBQ7nfkRRzcJWIL
XgdWexhALkNx6MOCMVZfupW9JixgwR5NwKFMugkNNyXLN9ic7YdPxrG8zOpYhMhV
t86Mzs14SumQZrQ7+hz4GKNa+gQADm/DshPwa86vl2ARtW02AlrO6rtGxL3w4+37
0UhnXRrriX5t35nMIt9XsYn3zVzZfvzoJKT+ldi8M7c6qYDOrZFqd13L5ty8xmEW
JVXTaNYBREHwlRhAREhaJT5EliA3OipnKEMCZvjC7h1yi7oIFvTQD7h5JDs2IFOe
eUqHRRzGxbXkbakuu33KyV+cdi3RqIyGqq62agcNxfIK2BIjMdDdSv3u1JglVEVf
dNp22QwAOl3U8w1P3vR41K9dJrzzOEfrU4hgt19N6vcNDF2jC8xFaYF7grt4v+Kg
QiTC9WCD3g3ZLw8MYbk8w0JrxeohtwLaIP0KK6v+JohM1jFFUshzKMjT7uq5cmGx
zXbjy1QrgMfJ5Zu+36hNuHVNdcq8uJWhyopzFrDy1Si5xjPt09+2Rx+A9kT/z2f4
Vakgw8E8NqVa+rPrYXl5QzK+xgdJyD2ICQEUxxMWptLLg6t2u9/pNi4zXhFeS/kE
l+s6U2HuB25n4KUMWtv9GBnShvqH1bXCCSbICy2WfkAOG2ByeHPnmKZ/HaSta8Yf
pypkHL7+2TtgyiYaogndPjjxdU6eWOBX9Q3VxVkzfGqy1d8Z7wgdUahF9jiA8qcA
5raYPX8UcKurxa8iSxr7CVb5RK1k/AE0jyWOnw4rLVVGJJxGDfmUfzt4s/9ac9Mp
Xnv3SlEyfHpiGDLaFvMPQJRpbhAgnJlW0VavlhcVENMq5uSWofv5q39UzElu//sN
o7pduoHizv33XKEEUmkxMUiwE4NMbtaC8V3EqWd3CtaNxjoP7ZBuWq0N4nKyY+39
FSokOz0m6aqgL/wTAGXwRMs4+QPqeRFcBgH6LR/YF4xqSllwHT3nnwjUcNGYQ2Pg
j3whLZY1aCP1nhS0KzllG3AAD+odJhBHsthCqkwhypApEaRqsyG3JG9dXRb6pomA
BpoHpGVKHHUbBbgH9UZUOMs74+Mn/OAZun71PyqXyIXu9h5zk4sWOQub7SU5dRK+
PBZp+Luve82O6t+0QCrjuOJJWYRTtrG/ij+t4sl8Sy6l/zUTC6Cs3/geUuyj6I3n
sRKKrtzX+mvsoAxOiNkmjTkyohFz8a2X9IZL/yzPput5+ED0ri9LbZwwq2h4ol+N
EMqrzSORxakkmE+ye6XlImk6xphQrcjxuPnHEd7O/FEDqkXxpC+MwDnlz9LZB+0d
YnbdwFlZWKgH25xjXjgTO6EYAW0sxks6pvn+N+Yehz99EbLRZWC9ExsjyVVuF6au
VrsOrpnIL3y/VRVAd7GCZpnSvYlAbS7dWbBND+arrEZllUVs2T3cQ6mTopxrejBr
6OzYSt7hyQmi1cBz5L0Uz/g5LqK/ejB4W//KfuKvAfAtfsgi8Fsy+UUWKK2pp3Rh
120b+6mHrpi/HK5dOjbrnhQ4Ntc0ZXyhAhIn/jQh3hJiCVQS8Y9y4UaPNaEdWoK5
c6t/HRpCuP0th3qIdy/Xph8XQsCfaTuF8XFtlybdos8ae9zwhfqaI/ZgjjKAcQJH
QxbUDxvmtBE1W4L+y28FkHY5UWDppL1NCweDZCOi0t81JxfRYWMscp12+LIUlTNj
b8c378NA9A7sW7uQMC2nlf3nuRH5NNUh05qajJrWGJwhh3JAEa2qbGUzwvlyvdU1
LcrxjJn6BiJSrShY+DORIz9tau0M71+2GOXxCs3jKO61EajkI9Cex7X4JRHJXGth
5KPlisyR76mvKjEwZmsjAx9vIZumay6KvdhQulpbSJSEJsrU5wQ3SN/q4hJ8VYZN
1Qe4PGY48t3OP7vh9z+0xczGsH6Ggao5SeV12xgQsjEv1GuWvvW+Wk8SgMjYtDD/
pEbG1FjNRbYLTDRjMljfwsyPqYHp2jharMYbjrOVyhxtr1qhm9DRzEhMunb80gYH
1Jxkb94oHcaNQnpWS7bb8SvhYMYjUsDDvoM5gick4WA6gv4X1YKhmXbLroifgau3
4ib8lcUEmckE0hUK9EnrnMrwA4p4c+Lm7zjZT67wHwnShJt9phCkv7csarrdisoh
vCTxLFFNrd26445Zl33noJj/4NqAqDHrapK1v/sfqOIMhKPAWt2n1N9Z7rhRPspe
p+GhDYsthiPkbqAr4FUaYYvfd1dUCL98XqErKCEcmVH0ygM/IoE8mBnq0D2hKOAe
KKHDaKIWZzo71IucOeuM/wCat2ykjZdaF8ab4KZkf1VxnqGRjIRzVF2EsFhdZnGT
mgY/J9wD9sNn7AvIQNwhYBiQlCCtPdZpz4RntVo4MMs71b7H4f6pv8aqtFvc5z6q
Qz394fWPQYTzcy1OaZD9UfHiWMk66yDBljjMsJpsZY+Uc9HDEmFKU+MKP3zQEvm2
8rVSxslgeSz4g4ulzFUKCVEmkf71BAYZfWOuo2VGzdKbfk7/SRRF9AYLNFz8+ZVF
CA9gVD1rokFPP5Z2asHOL5Nj7XXtokSbUZny3jXTAbrgbRrUjkDSZQneT5T0A6fm
fRBmbmbret5LBe9UNfxzSNv2IYUgw1qBB1+s1Vzzn5O5hmhWKsrYzTnDWnrbRYa6
MTEz8l58vV//Sm3mKcRepwhBnQYnyWBaJnUW44VGQkDmPhAYS1ERoecb4IwynnF8
kynvKz+AesjHn0wDqLUKg1MK4ey0F9oVf26fDXAeVEZ43WecjLaWFigLcYIbPLZW
nBt7PwEgaDg/vJtJfmxhuSRRmopiDETwCk4lKOly19YcKrxoZsCkxerv0NvEAtJA
WFf7ZtTYAiyOEtyQ+5H54EQJHuuHsLACfhIBkEo36FozHnh5u6p5dB7folfRTMzu
uMMJUM1qRnAXZWVpMIyt2e2Yca4RlsKiqZOe4tIKcDoV0I6q+v+0j/Hph7ynhskN
YGqRTZGws1uQcaP4Q6wNmTb+MM2UUCIsam5H44ebNHnMnkr7D9W7yUTxb5yL5XhQ
t6Y7dYyvm5jHXO20DUfRZ0j1U3zRW38fIQkV31Yql4yVAl0Zu3WC8NQUvamCWq0W
vUSNw77kjtHoedjzbzIPHlZzFDbjJbT9h36V3f6zfscmZS5ATp2EU7V5+QrEoQDZ
YTPJItD28u0gGfLE8odQpbmDFSn5ja4fY+srdK0D33dQKt9RcRr4ZmdrzUcHd6AU
82m5RHtvgsf4FWrFxqDgcVkN0wqKBpPXKc+VWc9wWFBZEwUkQsCNgBRPnhuj4SNQ
qvXlBAfPI5xOLKqsuya/XrzYdI/1OmDkjeVbddTDW7l4m8NxEoIygIMzCMDB0bkS
10Slu8b0tcBaOHlV0T454kAUfJAPAlQhorrTp2xJ5KNqJVlOfAzy9KkrH6nBqQVo
a5enzJUCItYLVIvAbrap0X+aXmo6xx94zP0cC9JLL6nrJD2oZwvUP2y49WgnDlqJ
FKrdhdAkEuXzt3MM1Yah8P5bZUIe4BwdNjVQiCaHGQ5tmxio5hrIhXGqOONxmwLT
iAG7UglHllDJH1088FYsBSG468/HnpVn6VwMnCNvjUhw6plL80eBmP/UW6RTaHP6
xVA/ITrlcv/CSByhUMjUAl3ZRDtEJOrlcVq9LhKiWU8f9CC4lUQMlPPWsJiNzbEF
RCgIj4cooJ7nCy9jTSFmp3g7Osj2SDqJjGOP+PuDsqPq+Tg6O6a2mXs0RWZqXRJP
GiwRgsvFZQMWMXcqgvRs9613LN2mzVoUZHvxd/xBe4q4rrEFmQGxhzwT3JThQ+7c
i5eat378iS0FyPBxPJ8BOxtOAbbPB5ao+VVF0v6DYiO+XY7Drkl0swv6PefjcSGM
FkldyUT9OO+b/cptO3sJGFyzf6FBEBXR52TKdeeiTUF7d004nczU/+D5XyiQ0Hnc
2/fa29phkiHGCQxnGpkBvULFmSsm6iVsuH2pOacAGmbfy8nNAySkbiLsnHlUGrxM
o0E2u8FoswFJ+j3IsIsOGmaRYqh/QbB8GmpweQDZhjkW6QOay52T8zkrbBK7dUSQ
TpkQNvFYOa+Ypgwhx3WfUFGFLoM7SFtu3FX10vcQbZiCaxDmmkS8h1DkIA38L/th
pZPRgdyLO4fWp4j8vPZii7LZLHsMgn5AjXatneen/0ZIIjnQeUOxy4Js1kUGCfvn
K7KIv8GQZ6L27K5o8BL2a0svRdGR5ZiNfC8/pq4NdffTUaetvwRPOue7KlKuqfg5
L47aafNEb+AmmZY9DaykwgUl21OhaUDQdjKQSKIkSVgDxN9OSmcLHL2i5Q+Q4KP6
7SteIty7RezHW9veVDexB7U8GvRtx2dmBcCkGv8TQ1fgfvfWiIWhgFHA4Eiw8Tm/
q/AMINBGOj8slwZQzY417w29qVGi4yN2sOcjptMZ+ZOtu+2gZtTVOhp3BimG5EPH
sATejZXBild8cT6FcJ9Phqf+nWFJQmNIOztLMte6LezMsyaVL2mr2vSc8w1rI+vv
Y/nJOsfxiSBVz50j2jO6na4lEzHZalD7zL0KuT+cjVwD9EFQLwS06iPj5rfcefRU
v28iRtPYFvPGpFexFFZZDu2grCaRrYfOpE1VO1Y3vDmJ75ff72pXeYv4/KzcGZY8
/U2iHMWYTEhvL1DTw0GuDU/WQKkyIzbWcc27f0ybm1pDDqIQ0ONpSf/9uWM9Xhk+
VWN0/pv1zIVtoeptwXFRiMxaHHA/F7wdzwpYCc+aH0xZfluZXGaoAeb25lUueilO
sCWQRSOCXUrGu4ekVt97iqvnHWabxC5TMdxVZgZR8ZBelbZC5+oaaTpTKq2OqJqn
TWDD14sgiC0wXjDu10XULtPcI8Ey04vONOIhw/FHHXtxCIqsT/N8NST8jJiP485k
I3gQz5AwniBRWzDPqNSKveST8TZFI22OZNvqJU0buLsiPMqDoIGe6b7zcjsMht+j
TCji/CewWwxqOEJRVJmm9oBN6W/i+50BAMXSdw5n7WaXGlV0G5eKMZSIs7nzHpbx
0mNg3GXjSxUYACASS+/K/q9sAT+DVEdzIn7Ila918cig/ydnVLoftGMjW09o7MpD
CT3F/ULwGmfDMeVTk0jTXA3bNYbwl/9sqcSDF+lR5E6IXDyjjlySu43YFC8xmlMP
mVNftODp1Qmue5m1Zk5Ln4CkcyN2E98AiSdFyXW0h4sb7wxS1hzl9gmQs0XZp+xw
kpJwHaSCbQ/Bshq+aAfSmEVeInYHJPsmmd+ssx8UHyPDr154zE3orGX5NaIZ5nut
TtgnmTUSI+jlA18ElR/bdql/IouUvyPF76HP4/TwicS25Dldboyo+dTlbdSwfLX9
QLCaH7AjklHen7xYj0uqg8G7S9PROuZblbNlxLcPu1Wv9n7ghb4Hv/KmK8mGCt0r
9GpaKJocmzY5qbcVvfLvUGPutJfdraeqv2xPnhlRJPKyRQ89lErpkrl16BcZY9gW
42T6AsdmFD5AQJvcrI/sc8cSzfMWLlxe+dov6TAHVQKCM7M7Ei1V4vvdwWQi1am4
G9bgwSXWyx5/dnrkVxbUgfcnoJ90i0H1TBWxZ9nNduBYW0yJEshtXcCXBL9A+yq9
9s75XQIjVtri7S6uifa+Bb0KluIufsytLbG5/kKmO/RHLBKYOWCK4AiwX9j8eQV8
of2gxCnIjzQO6ZGI9WEXtiTmh/7QEsLKmwrlGr1Nl+UaxhehXDW/52pUMN9SxkYS
Sm0DWs1nBO3UJT4RfIrRc4sPeEFUwAyigsxH4u7VzUOo/fqqTkWLyyI13IQS0r5N
QA6VU84LJ/NLkG5n4WnV/odsl0NyHHSrJNDVUblOY9UkEwc+mNqu6dSeY/fZRi5m
Q3HAA4HFQpSw01NQDJ89pKDU344QsySFF5efUdeB06xZc5Q6nLO6r9GBOQ0Z2khy
rHwHVrqfhl20PmSFvlgSayVdO46OPbMyrpIyJ/el6fqBMZ7TDcT4K6tbx0+mKZNV
VqF1A6Xz2xWsF3i79XnvrvDiD6qkAvJepZNoBpEF6U5LJEiAHMST+u/UD8YOzLYM
RsGRedmUgBgUdil0+/gTbTvFE5baII7x1Bd9vXCTyN80H92YsiEbk8+qel05/Tn8
35I2gZBlQfzISk8m+YljGvrRzRYU90hnAV7T0JCmDwPZKNGGoR3Gp9N5NIA1xajN
lYkp7MHy8f7722NH5uuAOFzDSC0DFK+CIiJE1FNObmhEUtuHUDFzKWwqxy5rIJ6I
2zoY1fJI0Y4650QeFz/xyNlwuW0n5/GdGvfiQ/g4yWgRje4NM4hWJVL/EHaxvC8m
iVTV5KNAKYDLwNFZDr35ila4RmmD0n6Ui9JiMhnRHimuxUFCxto2wcPb4ZVQ2l4w
Upo3Ul+LychxoSOK4tXoyCh8+5h+KS47jeSRAwtQLcVGI1TWjQbxRiq9W/dPSV5S
zdl/aj6X72s90Sxg8vxEtyEcH+XglP609W+hwAjUsuQprF3dZxVnpfNID1JThx3q
D08DeEMazCGOddc6u1qc19FavjwsaW8M6FeNeOCio4P6o+lqiVObPsK5s6EG+AC9
Ln7YtDRabp6+jYHYy931QJZAFHqJz3uczAz9UtNpfvR4srX0hYZpYzaSOGN+B2Et
zPe47NCZ5rjbINPOEpLb0aaJMZkAyxoFi/GUmBZER7QoPbKZs7QayRrZ86bE7T4U
pkuLcRyp3CvjLkEeNGlXyuk1dUVoaqUOqhg9ToF+vuBIKQKfyE99MmUA1kuvdatM
IB9bHnFSyzOQZL/FC2u2kpXgKJ4RnKJxxzRZJGWnv4JTvncUV3ncUtZkzVtG4UoQ
oaXXm4UqcRCfUxsR2RD9Ed1pGTs41eT1/vrxMayusYl5l+MI9HDLBPagkcMnyzT6
jTl6QsI/C0vF0y/10PWwwgc7DDTuB05z3bevT47e/1Kuhs1K2iQD/VzkY1EwtFwu
Prh4KHwW+S/N+Vf7Enfm+2VVK/T6RKbqdHUhX0I3L/qyp9E9a7SUpJU1tYDDtD7n
mHsO3V2poWGjNnDvZT1hi/6rJk3YGfnZ2qe2mDhbctMecuHn+oBL/A6ybfBHgIdR
u0GyLn6CUvrt9Ztgv2ROSXwpKnR6AhhPtobos+mquXbhWeY3St2ooCM8vjULddSR
5a3mJaj/7oGcSzg+YFnHjGDEcMbg/CgSjeKsKOXiTWChEHbvz2t8US1a0pYfkSIc
GUZ/30atbeV/Apt3v9SGyvwnH3Xyn7J+u3b7xtmTWfbRCwcu7RmVcL8RgBon2Nm0
9Zy607ftV9WP7ZU6Y+HpB50KxfEnWm/+8nT/EuNGFwaFPSfjpCBAOL11/x8tk1ot
hWzj9fMSoPR+h84pnYNfdm1ng0ugLCcNPKAH/cWM1WoWVeoKozhpwnCazpt1kS1O
8SV6tWnHhvKMYsk68M3+HFLf2hz7q2qotgwBeDkVrSU8HriTgEyBloL7mSyp8u1S
NvPuvtnNkPz+1WJeVaIxCXZ5TOq7+2dz9qLJj9KEfFu8amPBFvbh8UqWYwS8sr4g
izglB37rfilaUq5dE6b3lIhUHpRmQ4WLODssiI9DLILDI3+te0yVfcqPimKuxhHl
VspsCCohtIH0R+NeZzlzo12bspVndKtnrV+JIg7QTapz/Qd+Slb/Sbkh/5BiWq5n
NpoXyOZBiDh5Susjm9HozpNCx60HEPQ+GbdRaGeX1kzm7JnN1ivAMCZ1Onc0VbGV
NfaXSpLPpCQe0WLntUoM7sG+SInbhkcSCWW2+BAP2qVU0804OrESXrcm0V02aoVe
N0LWKoxnxwhEn3Kpu04z1tIlo9LcUtCtzZwOvsDyRLlSs7NcCDQXUpL9WIbNpXBu
tqFAA4OnpuFlkrOoyWn6+Fo7mlvYmKrCjzFnRIbLO0DYkjJGhf6RLS9Zk4az6iD4
fGvth4ExqWYyq90ff/6u4v0iCYU/KxWznObDXZCKO7r3YvRP6RMu/69HyPCbZpNX
rR9D3uYQh2488aaZBwe8T6Vg5BVQ4meTNG1X277JLSi6p3m4mbi80wp3eSRS9Vci
pOvZ00A1SYrSpMElxBijcCHRQAAU0M7cpTkn+OZn8QVCgsJB7a0w2Bcix4Z9h3gw
tvuKtPZHzFyV2goaypdPN6PkZrQdmwetZgsoqMoUsEIGteX0u562wV7NusRCQ7J0
Xn2KQ2B5TtBJqhyg8Guilda52VC3sRWl3M6PaX1M9n3CQwBdCU4RtrbJRiBVwrct
D9KlZOXW1LJz9B5srgDZ6flLsarJhfP99PrENh/h2sjUgXX3eVhzDS9bZiWkHr4A
EfVeVGsvUArwubjFACDgNU84naS12p+JntAI7AAc5XFKO3cvrVs9ibjW/cKCp+FF
R7rYfji8ugGJdTSXW4xUt3u++VNbR1ddxR0B6E7B76ruWghm7y/uv6lH5zxf4IKA
i7Sm8bfMXdueP3sU9RiICHJ788OH/pLOjCyY5oJPFUdBmjnO0G0ieH8SHmJHge8X
fXDgGxNnGePSuvy4DIHPoPG77xQAH4LTmr/qpgu8iIi/ujwqGQTZBlJ/PM0sJIIV
nlIrQK8vnLiEyR5Fpu4hBsB2DBMIDWMB+Bjn6uWc+zWaxebHchUQqKrz9Kgtwl07
NBSu1dPCV6vhMH+xHVmx2XM3OxHRBDIDxO4FzM0E5VkO/35xK7C5qKx+C0tLmp9+
yTbEwUyYQMrCbAL+hXjbKxgDqWksiymu8frzNMD228ODawlsyKUoCU/QeTvqPo0l
LhF+0nwSeK1OtOj3UXW5YPxUePIIGYghhNhpF4V7z+VZ+r3kJh8BRJkZsW0CC6e1
sErwcggFW7aDqKIGk9DE1+qA++RNGp40A9ceT1o6lv4WF//NkubTQqpABxlx6XPp
CNi2XXs2mIfxSvW0l0dI5dX2aHg8PiYTTni0Qd93h4Qy9gZnZ5UmzJD3DlxPQ791
e1K5MRmjF9zLNKT6foa/dM6miSlhJ7ovOflmgHnbNYsaynYU8krFtcdDtgLfRXkC
vRx97+wDhsQ/VGaHEXoqK7G3PcJxMOlWA13MgoFUOkFuqpvU4VPU3GyOV4pdZlJz
kgn6mb2yr95UHLp4fP2Qtu8TPKjCL9aHuDXt3NZOqpfxCGqLGgixJzTAysGTOXV+
UMH7cSXIOceBudvecr+d4Ov8VgKUyuyeVCxOBP2d5lz+ZAeIQYGV2hI9QVsTQDNe
Hi0mRlhOsH2ir07jqX5njaPlFZ8oCQYu1E3l5nvaobKbynXTVq2NkUoNOg4pISH7
gtF2JnwFVhneEC7n9udJySzF+vdnbZo2ANt9WFH1ZI4S9S8S/3p6DcVe2SUV82CY
VLl56p8QKKWRd9NF6fAkNti6HUIM8I3++Rz+28U0XMCjeqly54bqp2sbMqRsfT/R
PVsfYzIoLUJQ2V3rHQ2PesJtzmbDDIUELBq++1Cvi4vUq5ElFbhMrZCdOGKw5LVy
mKO0XyevLMIx9NvEI2F41v6OhCJ3tfk7yXcExzulAZrJR9jV9B9Mze9Rdhc5jX/V
xQSrBrivg/Xj0HCBspQs7XxeKbEiDBZ2ytlFsSMxLMHgOVY0GNQCjX/7ZivGwmds
uqbDRZ2p/bnJtq8ajYAgFH/ZihV9TI8uXAvGOsWujGub41LZ79EeGzanjDkH5/vT
jUQ64r+nTvc6enqqQn3OqBpGDT3hNozAtaH1A1TlHGrHWHyn/yhw4qTdfdWo8lCA
A/eg3OfN0A+EVOiW7P0oeDHukwvrQhryOZ/jmUD8EtkgkY2QbDDCgzBQbALLxKME
1zhkXKyxohWgFqlKFzjrginIWsaMyslv+CXZfXiHgZcMWjtY4v5FdPDtFOTFy0lk
RcucH2hBYZoFiLBkpVw4X99BKvuBxxgV/a/PJaFu/4dkz3qmgnl+i4wBw0eXyMSn
OXetOV5IvkPV/a2mKf/io47mqiS2yazDvSLRWbExdiQVEVyNBH8TzNO+NYJ2CjVY
acN424U38kqSvcoKGJwDVB9DqUQt04PHoeBkuxkJtYgKZ9xF/zD+D+HUWjG4HAix
3KmOKjXThDy0DT1J/cxIlNT1btlM6BpVOZrvkB6WAAKKFeSmxiT7Ef+gMb1jUlfX
zgxJYifyxEhijmBma5ND9wqFcYytDnbaU9BFqNM/3jrphvRIBcyDjPbq1JEvLe4A
ZK/VutJrPjanixz6HjHLoa3dd1ZuPSM8cp17ej3asbPkEzB7zKUncgptthIXQJjF
EcGcARvrUuk/HmEFmnCV+6/60Hxk2oJgNEuV0tbn7OMrhNGDzJNvNo+vE0Ut0DOC
4YCTLhdBqbHYlylHKLfBR08C1048HKIbGKHQtbXAsiZMqPn3TfdETRIjaIxEbP/M
o3pV/W2ABxW3EXpRKz9wlNl3ujex7DQSOWBpzcFabFGXSRTLJ5cYrSXuKHnFYXV8
Q6v4eqoEnhLlhmfVqyFP0l7HnEFwgvbhWXHDWnmzPhAM0Pm6bW2YtCKRwJF3+k8T
ZJ7nok0S8hJWyuixOhNXId2lSv45sD5y4rcyLP/UMOOmrHPxajayH1ACZ3KVttF9
BkMidS1Nzu42MONXRgJmXhaiABgp6blgUAZberyMZjgiPLLZUlcPlD/oj6ScLpSC
+w+uZemt4ibGylCQwnMRDlnzKznu0C3Y/Ae08U5J2cx3NZi82rgjZ89MYxmicgHW
5Kv6tRBxoOF+X3dsJ0YpnmPgO99mO8yPkKotsnq9keyXTZ3zKRFKeJh8NdKO7Wek
tIjgERU/zQVg2ySSAKNg2yPlJMyQ9KVzeBZEjppdl3t057EZI40M8OQHYZeGO/Nv
5dpMPirazmrtdrEIxPScVnLNJnUTh/DVV57phWsizo/CkzBr8TTyWjEKX1oBH2uM
1uQwURQE/gnme/nSHMsQv6eGU4UYj7wLrV/reu0/OECQUXSKJymurdfsWuOZPnk9
7Fdv4ORZLRFLyTrcYoQc8HSi7kxLB8CmCwmDU8D1m41bJtBOE5tiuLqKEJm9gKSP
VG2d/Wz7mhN5viAoPeHLPWBl3LcuzEO5aG0LSJQtcBkr5yWs7hU/J9N59NljaeSc
Mw9mrFacNyxVEgPcxC9pWLnbfW0yXmxzOqOEYegEtEvTJdzDzww9iVOw0IQCXaXV
et9KLssfesUUgdVtgo8RMu+nQ6ZVoyPq6eNDx/XyKuBwGvxhMgwbyUsH0pcCuT+3
wXEQM2uQCFexjDPwjhfP1QhewyqQzDlqD3kgEJwoMv0aE2yMHwmfsyZTLDIDwwog
hlFOND251+rrJ5dqJ4dYlpQ0JMKoU/Y59TCIGK2d7Qq0qQqKzNx35Jc7JOzvCH8X
2G9eMzgdWBniB8MeIUiQF/CTWAi9/lahUWS5dALow6DWJxGddSRdq0ptm4MvPgq5
j46qcvfpaNhdGC57CtjEMrw7mNi7sqev006uTq+eIOnfwvOGqTcBeRQL0ODZma2K
MLldIpnjRX1xD+ISEDJhTIgA+cO87PNCeCOl6Bfgtk5YqJsfPciNPBX32hBgo2K2
17wINELCene+T3fZwp8/cYSrGCtO+NQAzDY85I8vUPGgA0vZqWe/A9PjaHKxSWTp
y9Qaw9ka9oApqZcvhs8HunlaBCUbm0JkOsERj0OsSzyDUCvXFum4GzZtyQsfZGTR
b1BuDYu4wGZfNLTRHllS2Ffhj05QJkKhMjDaPFVNZbEqYAVMdSqOEq8Ws/MlVeH7
iYheO0ygi04kxBrFRZN3L7aSmD0Inlq2PBtl967gZpIkIyvNzOnQhL0BRKyGimcf
T3FafJRi6pDr/H9/y64aOtnH2erMpVO7wv1wnBcbFCQ8szVR1qpT01LgPmThJQsa
xdQSyA0iUCMC3lg7MaLuStTKg3qfef/vV7RfNuBSVc3vsO2T5554K7SwrmhJ9KkV
XUUmHGotY0FTJD3qOIwR+zkiplyLyJXmol5Noisre3q4h7+kPxxRGMBvMRQ9suxU
FcLsI96vXw/GpIL5zFa6gDT+KGAyLe9WvaEg+vmJ3LTXGakIfqLevahh4Aq3NaGP
AJN/oTEBvID255b7YdBlBv1/leN6Q3dQQJA16LIwwXX0ujPhIfqrtqr5ceY6gUk1
JQS+Afgle3B6Elkb8IkDz/fx7JvG7aEXYSGNIYC2Mx2N9d3VyB6L1HusHeb6FPiL
tD69hIvg+nNWHLg3nBla9sbLLuHxNNgOI80zFEoueUnqGBZLU8fRf8TlYpI15YKD
pTtjrUZqG/k7lqN27MoQ2OdML53289MRIrlE8ZPxQbdStM+1BmHBJxeG04dyCAHo
94i5Vu9MXzHSTQX2eKZZ+IGgvvXeDMKonVZXYeP0MRer3OtXbhM3jiKKyJ3x7LSL
KIEnmTjF4maw1wW9981vTPiZfKi0HJePD9SvXTy4GcBwB0ylwPll8V6gQlaI1UmY
Bnp6uIoGK1sWzQ8PTOYaUfp9dc7bo0bqXekYlYuuBTN1OeRVYPitfWkwdEY899gP
kTMsNNynES4s2jtiLJbNSl7Xw+dcI3kqeqj+N0+yO2UfXHZFW9rRFFckXzFBODZs
vjn8GjpCvGfCvlOHx+xUXo2pVnK5yTqNAXR57tqIxg2MhaIMu3mEXpzXoMGmCv8k
qMlwnkSeAGqWBGBwZWuj//oYP62/+W64cClWB29BBlj2Hj0h51NsXGhW/bnN/dJ4
stBB0IDds/dESaVMMRQ6mZzmAUFRO4YPO6Ic3gP1LNfszCxgaLCUMDpdK0RLUanA
dBNkYAaFBDgErQlrGGV/2/e491kdNGl6VkajQCIX357kaQhqQRWxyForiuCgo1Aq
GoVbshosow73UO+ObMd+KFMQ5GWfIiLwQ06dzSG6WPrcemlWjDkpx8NenkJ4rsv4
AeP4tI9Z+gSxjGzq4rhZ98a/VuCGUI/tq6XilagEy8jz1PXaE6/eQ4zJw6XOzRqB
+clsYOFTUjHhV/2xTl46HgdmHnRmFQGZ3eEh3mCANZ9cn/wOEvGCq/yUPX86hC/q
dRhZx1Oa+MM2DqwXsLwBO2+SBJmD5KBiXhVaQKWfNAXUvxM4ABpckYd4Mv/1zDCg
vd6a89eOzlQN1Ia3zfPU8pQkzKqwPFAff2Q9tyqVVdDN+t4nTm64vM6zG+0MyaKX
U7yk3w/Ja+ZxKD9N8nE8vMWkq9z1qzpYWdrKCat8arKj9OAwR7j4V86tdfa4kDRW
r8EFrdCdW7Uk1rSz3LkXTY9+Us2OIzp3T/SWMCAxKiBVxHhEdDjVSRVOXl+5Ng3h
1ICvh5ajxAEpXJJIeDh7mdTjghaoMsK4+toVgqAxYO1Lfg7hSzOo+n05nNtCpuHB
llk45XR3kOVcwei9RIkw5no/dhydpQIYXwp786uchSqHUJkIOqQVB2YZdO12VyKI
SJDdPBT+R65KbssgxxMvlG616F9aB0pXgOECmIxbM9N7kN2YeC4lpvUWN1pN0AMU
m/xhNiy9WBgHxJx0VdlgOG4Kl3eUSAZxnfuJVusieaG6a60a+YF9Mw73XSTv8yOa
jKtpytGUZWlBv0WjNMLnU4Ft7H9CYZzp5byDVnroxC7KZBUd7SPcqw4o7uHy4RB6
3+pedIoAmOMAt7OB7MBRw8SziFL7n0to/7AVNy/KoiyFDVLfQjtqFmmlBDnG3HTJ
W+g6afurvjt4fuLE0aGT/9ZFIBDBuc/Br86vSB+HnjdpUxMou9QY57W2PxOUjQvA
KaxOItZMCRJXy7jI6LpaA6NPw2z+6c/r7mBjIWzurlvGyhcEegS/K+f9/lBmnODB
GunHfgFnluptd3FbsbCnwgCHieVuHyTiggdIexAkLNtgZC+5ubGdvTc6+pObrLs5
8CZroxuo9xjJ+WPNgfj6JRgRwrVJWo99epxEL7ngcSsfF68sAWGkYB7M82PEfF+1
Cutg4lltYsY5OwyLBBH1nGUkTVueizUdvTdrXbpS7mR/zd0jdwk9qKGkNAYkv6l4
P+qIkee5u+YyStwbpYQdh8QjrkYMRRnCe7IWplJAWOIYJH7tzyIYLKvCaCVReS0l
llG3TuiPBkPndAhPJQGcDIAMzgneKd1VmcG3HsM3WR+s3X/rgTi5s96YD8xBUsFr
VbeQMHqWyTlcG7EQYm38oQjL6DM4VuvoyUrd5sVNdKBYqJVVn/f8o0Gat+yJ3xuM
oFe3whOGpVdzuTmkmxfH2rW/sj0VIiOmk6oJzY+cIaL4y3jL5Lhfp78JeIC6cY6N
54P4hYeDUxA9S25krsHpn1gH+7bYqvkn3QiS9g3FxSbUEdpG6IzgSUVUnjO4GCtf
J0tZ5VwzdURnMdTaMskIjEC4T9yEYkhncH8uvNJpYxgbXfMCaO80HOEUoyUh5uwe
d0e7jL9ivnbbODdSQSZMSsAPC1nUhgcypjQMqDLttG8TP6DJZi58a4U6dCs4MCSl
QUM7S2UQyhCxb2EfehJgezGzJtHI5EpTItFBRqUGzBR/saqU2zGnGICJvoNnnUvu
2RkOBIflo0PgYjzTsK8dfmdGQnP6a8qbdJJh4qKz0yJv9+A7lCEUp4JrRbDgWWUy
8JnIoUZw70rwI7ct5UVn2P5KKC9WEWPYwx3svB6tYV0+zbwVPUTFZmt/XZ4ap4gi
R19be0S0myCKP6YptYPJmhz7yY7tvDjaxvLwvOE/yKimDTD6lnZy/lY0jOzPXlWR
afe8eLreCOeMH9jjis19k9gUbqsWCIfKyrfyXysNX2WGUD0QdawW2gVS3qXupqfk
dYTzIy+rdApK9J3qMTnlEF/SCyua+rvgX5PNt9jivNVzys6BZ1MvffLptt9JKSnG
D95tqX/li8CNZQAYcp1Wq9ZZ0/2lB/wZs3mbA3LszDYrR0ylBNpeLt2jO3BikbNz
cvFMXhrk0Qgni0YSkwztGOfEsn3kRJnq77VUtpWcTwgdFlLGym10CSFcsKuhFxr4
CZwpMcwcYw4TlRyjBxCrPoeKbE/kEqycwP4nJ0EVahK/bCBszhQglHlWjIlyWlGw
y3syGoupp9F3Qp0w3Kwabm8Bf2p0LsTxuCrrsHMtxRq/1Q1I9TYOjThrjndUnahG
DIDmBLA9Tz62/u24i9/b1BnSJonKYWHpYyvBXSSUkO/mrF+e+LdA98B2kxJv0YWY
TFE5V7JO0OYUaZg8J+OMgcV/ODZm1rrCzak5/wb3PkHOi8+1ZnfdpP9tmnGqMsr2
J4DIg2kaOEsMGRMKylrv40UVbvwI1htPjYjhE9ZrQ200uGZhdivHzKHZGLDXhOzh
ocVUzLYIhjrc7fnQP38vlGisfok4LO9fhkCkTQUkntlSIRYgsSxjLsCyJ1p1sWzm
cZ39/75CT5ilLA06rkOWaNmoEeY0JDcGgmULk9xmojXlO8TQzSuV6sKpq8pNyD9S
jmZhmzKHMvzgaHCesA50YXXHtJ0CYVIdJank0aKo+oIv7sl4OEV3vs1/JZXjI77A
8OZ+H60uAjYh+qjhq43tGYdmMF9cWgMUjodxnFsWEto58OEtZl8+6No6XiqvFC8N
gg0UGCGdHmpSkI+2n+GA1BeMYpGo0c9InH88Zh1OOAxN1piHyp7u8MdSI0XvD3nW
b8Hfc7BjS0b7R+QpzJ4wh/nxI1//qa4hHvv95N7z48DiGX/hkh55t71F43jkMNc8
o1gCcwfx/vYgjA7Aa3ef9pz7zhxn8Jz1CNvQFiPecxlXjqD5bunH4BKW60CtB5xv
tBlUlkMX4BCqrrXeYa1ee+vvm5wNJmSlzzhKVDMf9bRoLyDifNOULpw/GKwnUFBQ
GR95Iy1yPQOIxIqgvRRgqCxxttCDX0Ta5kJnGjKIW/6Zp5CQuCIpW3/GOOnj5t90
PGDgvboa229R8TAsZrtzqMNqtuzdzi2bpCulcNlG00QJtAvMGpIlr3wcTBHbL6Z5
xZ7MIT3q7t4XYWH5yICFK2ADG6KXg73mWkp9ktB+P/yNRtxuEgyY3yj9yRnA3hvi
C/Oo1e+0qasKFnTYvGTx3S8V4B13pHCmnRY+nlE+mcLUuyABndf30SIb96TzmOqR
v0qLfWqOuistbZ4rS4b2Wr7NnDTrQNXqlHb/Xz14IYrWoyYPCQAcL344S8kYndoT
oL2ifhCwUfOE5ie7m89JX+7yC3vAn4xZHfFDTffR6BN/Kj2K5h7LhxAcXVMSrw/1
p9TIIEG7I83Bq40RrJ9SU4xI3+a87tCkr5aWfDxlTEYtqS2CeuAFhFSKSSSyJGaW
SBgdCmo/q1fAyvbaAmGIR9wgTDtFlLQWICljRcCZWic9wzVrZxHgfaR1Th7MJ4hE
1YcYUE4a4FEJlFSrSex+NC6nXW+31IeTucxsyDYP+6avzE6ea9t+cz2af+cIHt7H
2wJmaaZ90+KoBI6XiwANR+r+ETeJg+ZdumFvhnlMMgO0oEfUPG38DLBD95QMNcCQ
MKudPs5eRZRSo+IWeSmWNadFVKJvxAijeUjaVaxJAI1wDW5v26Lqo/Z/0HChDzrP
t6vWBrjhoZaCfYi9p2bfMRzQ5A79LSq/iuqwrD/4ZhpgYra//tULmhkwv4AOw8tR
1UfPp8ZMGVKRP0bZmsf5G92OdAj+uwgaTkqhrukL7WeYjN9Bois8Rmxct9NzHd3W
3ewuiI07LvMQ5D51DIGomEx2qtrV4kB2wWkfb4ndOlsUneRl02toARPuXcapz5UD
BRiCThG90J6VuqZWGXxzFDq6tcNUB3aU9TeMjuBRA4+nbuDodpcZ0l2RPdqp4N1w
daEeMApqM2nRizWe7juNWLJOfVmQG92e7MVOOVWP22pAULn9hZ3zjDxzp/cHmleB
hVC2Dcyg0A8WhQmrXI3UP3dvoO5/mJZeA0aytsJbXZb3NA0VmsNVt9k0YYza+W2L
r4cEl/dsfM+f+ct0n/XbIsieJ7kKFc/cmBoB7ut/ppsW9XRwJTNj/FdHMRmV3S5T
m+IBc7n5WzDiuZncjp9blbO5VjMOQ5xuI2tfQxUsiWAkrG7jizgQKz5cwBnzUFsF
mq6oRAccULzlqaacdfDPfhH+wahj5Zo0w0ZkLHnD1r0yBy54HID3OdQA9FvC5Q0I
zcBK25WApEUldqBca5gIkRPLQrp6fimaj1N410RjN2oLoJNmFBQ30VP7eZGC//GE
zygFi0uRP8Xen/tFMelMx+DWDMA3tCJx75oFR23U1zuF/EvvFDx6yAKYLWamTtG2
KYoxFNUVXAyfX7R278iaYVMywKFDzTL69IFaYXVWCAJlSXXovD2L83B03JR6O2Eh
RV9qQzWVoVuqXZ9dFrfBPJpZckKy4VC2JnvCVgEii79lJlxMTsCtYHByuWtYQllW
LlkPF1TtRCJEdTODuv3jzdQGWt8e/O7IJ21FTn8+wecjjZ9zSyXGJmwMWRbdPeuT
cJMEWMfeSia6DobkbdE0R3dyANRdZjBw86igw0dHWQNAqp1mbCeRknqjP5iVrbA/
8EgZwhOz99MsIeqbU9kghzDc4PTnZkCiVk1/3Lm2rfe7RY3AjAN1Fx1VY6etDiHR
Ri34d2uRxmRuvRJABu2RsOK3mXLkziDIv4hs4sBErRvz/OyjJsppAMclLGbe1r+b
UNAPn5H9Eyk9bo7W4OawE+CBv1h7IowK19soJqPIMaIaZlAz7p7X776sG1PqtaNU
vnyNjfezW8a3JlbXPGeFmHTfQrGPO79K60t5WnYjdTnsQDLI1HnL3JeXyde0hcl7
LkTYyxjN0vOJYuIB/B773aJYGvs8s9Wx39rKAW9XOc0Ej2gE/cZiNSkcha/hYupw
Lk15uaKIbPzs5hrpyJ52F+XzcAUUDhSVs38I7gLZhqlXw3QBEq08iPY/p4Sjy7vc
thTh4kCeIGf4f/YbNsQp0HgJ4jBZoIoyxjhABbd6A/NRb2fgPujKM2mSbFYeZFc3
4IhTDilJcSMwlx3liCnv+pCITGrhsZ3kFjP86vlUzvbMqa8PoA03E7REPnVX4NSk
YeY+RZnRnAVsDqJLlf1zDmY3DvDsF+aWnjOVPq9XwGtnz85/oL4qsokatAUF/fAD
DsOg/ZytUFppd/puSQgJintSPt4ylNN2VGzQOI66eeBAC2Fi/kB7ud3klXSoESkV
vImyuogxLUYFIKozwYK0vEEVLz0UNNBI4jo2HjW2mkoAoaJC4FXbbaeld5EdbZlL
rmbtodesrKpCzWtRL+uc6M5T/j1FiwFinlGgeWGsM/AThkqFkWvqhzuIOQyh9sZP
3HZQXh+DNhiaVt/Hn47vJh3UeolIWiIErSH1v5riivargaaDsYX2g25AzoX/zG+R
MOzMeP4mKl/k9mxby8MmVUDEwACWicVEmr+/KMhPxc5wSfNZLDCgS+zDSyl95lmr
EPujxINZhdBtDsPun8bi/knFDqVMhjAumCO5b8ys/fsPtUgSASYffARoN5hTO2PL
OAaUJg/jTg6zBvowtSW2NHxfxn0DPv3sKkeig4KKm1QeK3+Rizpf657PctlBl0ix
drXyUG12S8Rl+y0mVE9ao9oMsHqcf/ElYRGV881R5dsRjj9y9Cc08y06jQfeO7B0
hNhhuhBdEYYxRPpcfUwst2Edqh7veGvK9GVnXjIv1S3PfT/ONG7ESw7cG9CQidfs
OvnEedHz4Ma55WM5niDXdSoWHryDR0q/H8wQR/JZY3Opr+U7uKKPXBqCXJpIiKsc
wQA/0cwu8Nv/R3EQhvgFLT+jjp63OfND4G6K28K6jJvJ200HKBAjqusZ+udYcPD4
S78uyYRaKTEr3k9fhZc5xhbnxIw+CsCKvjgGbao4rPArHrn7i9i7hqQl4sntSY0O
1syOD9Kc0sKWpgqC+ekluFLuSSEEtjd1u205geLNEATp4lhfksUqynqxpjHNJPL1
4K2D2sYgxEzJWr6tQaOIBqS3+GOmE1d60aRo054Wp7OsL7+UHrXif6ccz5+8om8i
3cbZDRRSkEyGgmwTN+ytt7F321Fi7jUSXcA+J46M3FWAd7CZfCzFQQ0WJzfGQw0P
tG1rhp+ZrPfxmUIWm0KZgwQfXZvwfU8AHCLisHsosKKWw3RoQ3eedQeVLdg/0Z91
2mo8PHQoU7CKd3wjnxsOD87aooAzTcRFp5WvQdVOvkXRYJObIeOgqUM6dHLGRFdM
y3njwuMhm6NYYmf3PpsbTjw0SWMuXQo8tY1LC7XkLFbPbLBdVe6ty5PoSgI4bmW4
eRGbXxvs9Tkndyqp/Ke5P8uQLSRLDdRnrWafDze5QJLfmraMVMk8Rb+LOe9dKXPu
X27nzr/UEtNbQujcH6sTuIrM2Gq+xA1IAUhqHOqXEN++mThmWdv8L+PFFFUxwSoZ
MxHmTBDl1naBr2oAOwwB3Rjx+Jdr6tbWbyo8cIGAaraVCw4aMYrZgS11l27K1kCV
Qe/RIpdJEtKF3DdUR1rJX2PT1e5EJY+JdvKHv4gKCMupcsAJyVpfjCEKG95sO/d2
fAtwVbB+VUbi+h99cnip9JvCTaehT2Ke13bGLmmA/Awc+tJ4vlUGrrranCzltqo4
wq0vJc0207ypeMdSeXbjjtcQGJ3leXjvDNRvzKuZw7HFM6G46lYZN8XOdtZJuG3c
raCVp1CV0umRRCglS0KAWdVz0fJqBgrBR3i9lGcMpOXJ8Ko7Lw9/pF7fVDD4WfBU
zty4QbpQiit3y9prwBiz/vEes/DfqwqeoyO+Dg4L/UpJYp6bbN2cg7NFJ2jdHeEO
GUHzSpIAmUzmPhfewa0lzZPmnVn8PvvROsOYAEyJoHVCDV3zLyeI2hfhN4uS1Tur
UUump720lIVQjSHT3zTDeWfznqh4/z0ltKGEh20M+a2znNRlnzEil3ULnQlvmIqI
oGPvP0DAgMiyRtXdJ66DARpNu0is5J24xry5tBIIMuZMcllOYfclCjpcFIwwemAA
1j/rHhn4BZW224pCGf+kvYaKmK88x+Zt3y5hbisiGRO6V7AEd2w5w0bV/21b+tVr
8eCL/IS3r42pxq1JeFwLwKhav2YLkS/+jS9EqlO2cnVFNw/XJN918SXduxBtG2a4
0oktGy1IIIPDdFd3MHMkV+n/qE2yoCFX9Mvxxl61YRvYYOOQJxAXrSooM2y3n8hE
nojl5rcS22csUiwf0HnJrVepypAvdXzgcdyi4ccRQGOwKBRoe3cv4bglRiZJSuou
EpsaAo+kVaVHL5T4qnBQlt7orl9L1J94H70Saba45TVlK7zXmJSGuLGN3SGbgL9z
9HKc/u7AZPcoyhNu1KmMoepUKe5jJmYNsxN7feyr4Komgt7YSf7xYuF0R58iGiNg
HTiCkTfWteVHRzjC4D806h4EvwVkBzlhSWQ18usmoo75vVZrWIjTMrcvfMKBBEq1
q11vZaetmAovLzjXWCsTDuFU0syYkQg3uLyJS9T6M5DzmPebmBjSFR3NphOPDlAT
6b8U158T/gRw2hHyS1m/RX52WlKOtLtOB9T/kJPcyfem34jHWzXuKK1cuAYkjtiZ
c2qWcZgbu+aFhFC44xW4F4AB3bygQ0pj2/4P+u6FQd3fnZuclLc4FyKQISlNdbhD
wZdUpnkNonfVvV2OxPbbwEOLK5yvYc+R46Eqt9DHxffm2PiNRcEYMORcWKUnnXQp
5mjvWiuQjSV87PMavLia05VyiNTTnwlozTUmmv17k052jH1PvrAOfRT7BN02P7ne
sjM35VaaHEYphkjxOnoo6LhBdqgAPq2WMujhDGg/+4lYTgCSp/6IEiHKpMoawICq
IirOsq5yR156bhlxRipQv3wAI61+wCPgL5DoiOYHcdUl+4L9bbGTx6RrS8G6ANzZ
NZEy4xq4Ktrbj3W9p2CjkfwQTU9n3zdrelHB8ojIjz+m7UHV6OXzFy+7siXA7AKs
2dcjf0COcMjKXmFor+9EQSbPVyyZlFFyXswPzhmtueAD0GKuG+7if96f7C6G9rCn
JbmkqtfNqP5Z1pp720HZev2Z4eMZv+oY+Ar4GPWgt/kQks3SENZqujHxF9uqFYgz
LQDwI8Hb6aNLWQdo2VEcjURLwfSUf2UpjLJs1yLqPF2Ee0vGHIg3+SfWrAZFSzCY
toCbmDM6gSqY0rG3dkKmzOErHuOk+Z9Fv7mpwyrtBfDlyMZVi3q0gcxSWsxg9DF3
DAH6J4gPP9NcFB71tWRiwAk+RiGEJDueMe40IhkYivfCMWu2DYVrAyJjiVnL1vNS
TG8xBbqZm1OAYR6JnON803Mp+A2ZZYjblC2/rFD8d6dlb5oYY5+v7WUWIuxh5I0g
rpUXG2pxiJs0N+oeymomH+xJTSGbpuWpr0U5eOldgDi2IQEPkqP4R2vFnVWsa/Xn
ZWDJUse7tglPKjZxs9Qo4GC+Lm4GIfKI/wOE/q1AtqzD0L0sIAeiBJUAJ0oDZVrW
32cBQXALDRpJsWBrxFapVIYeBXPqrqGSyTRlx5kX+yfdcN2Ipp6bk9IFWLW0ljsa
nIgUpUUr7LdYByb3MUuMfgE9NfkQ+rv0tNugOJKKBbNkWp7POzFPqWbxkp8VU2ir
9gSPMvDWJpcKZqCLFdZEIdQj+qH8ysu9ZqqY/wiU3/TKf4GzZln7FHeD67dv1UXN
mmKjZ8atC37OzMVBpJOWXPbnz1QFvg/b2/4+RKpKy0L+naSKfMxJaB6BqixDPQhj
9iDgqr/wAyhKeQmOKfvbn4N40dOu5dlYYWMbd8t7OtgjvOSI2khNd4dEQ8eawQcn
uHsRaf23TEgI+gmVoClHiH7FAirUCwDHgM7n5aXEiDQT4gotT7fVIHPoomDZfHYK
+GJbG7fivOuCjGWjLwJDqJXGjKJB5J+zsW4geecvkXMmhxNWnAT3GY+4g+XObpFi
HGB2qMyMaTwqbtUq4VBjEoDRwoGRznIspMPyYNqMbpoxkSLqN4J9fR4FWbwN4IEK
MZEcv684c91cK21IzfazDUBAtQiNTBqc49Tsg4eUgmwg8ov3d1zRsTmQquP+mqdA
GA9+Rvh6kk/5rftzws1a3IvmhRp1vqpn/GsuodwnxViKw95CX1u8S3ZLIzbt2xV8
d4Cjzj1Pf6dlfYiawoDA7xSyBF0mzA1NFXSLUVOX/AT3UGJn5Vh42VlUTlAIY5BU
Q3RBNz2xeKdHfKwISoSZhm1c18T1Zh3v0pN/F8GuY9hwq7L0d3w10ftagz83jie1
qWOuhDOjlgUWZO/0HLoDjZT9cExsV/KSgAt7XquthyosyayvkH44rpjO8xkGPfho
9vaCa7etDN+Rk1Atl/dgK/YDRfrqaXEZv9WRk46OCSbrUDwSoe2ULdv16UA4Z6j1
ctLNsjgmBMZ21oYG/ZF4B5WC1yyI7I1bGRa17CQo7ATI4SlL+k2267vrPVAVFOF+
Rf5+JXeDQ/usuuSc/4J7yuNa2qF8wBVUbICKQYGatatRivDg8QzWX7GjrNhDFRyX
7OKRu2mVn4ZZnc/E2hEtJQ5PuKMfSjszd+4Sxlzm0b/7QyxyhsMNzCJevxqtaPnW
XR3YRCU/fWQNBjW4Wq/kmMWTPerp3olDkj6A8SDpXwTlxWCG9BK1IPYu5rdIwzCp
cgEmG16nii3kzr+23dY8qnlw/Q43EY4k8L7fTobJ8owMntjDqq3u8+U4RBrI4wQ0
eHbslkut3S8RR0pom9CZRoMe1yhDu1SdtvsA6Kp7doUljTqhgmUvxgTyaKsvj89x
MuTZ9y7zn8+UhbnnuNFFM6U2f2s0uH1RACbLQBM9Ox6wCNHgCQnjzefLcfIijLGI
T+h2Wku2GSpSftg6p34ZREWQuUD2YiOZv1UH7e8upmS1jrXZ8VKRDIulX7g4v+e9
cSJP+ml5yvq+zAgwjG9lEUZChpXrSFLRN3ajud72vFuDtVITatMTZ1+Lw3Bt9saq
D+Lc7DBW01dHf8UNKnVXf/eNrmVqbZMpoIpTvYbEjW0hcfl98k1Gj4JeBqdlR7e+
9JX1L/ZKl1cGH2/MvHWvGVJaHDfhVbHdXp6xNEbnhg/bvvrOnivcaUUz1yZkRU8+
0Lzsj0cvggEtfEuI5eE0H2SXodAca1OkrDcgWPumVVCsZSqeUBMAD8CzPgISA8Yu
6ctsxjFgYUvP6gnDfoSnPpQB7dYBE9pViRujJ2GJQddku8byw5XDcT8XkV4mz+RI
I4GxS1zWvZcyKA+s/G+zJUNMQF+HfxkPcBVNT1UTFpfow/g6kBywt4nWtjjMDayZ
9v3ZAARVkpQKFqHvswCijtfvp4uVDzmUXUgxmLxPJSMn2IB1T/ax9/5906fSsFG/
CCSruO+fR8ReSn6e05LXcRIKZA7oZMwQQzpPDMlKcy/1P9ox+ulEZGyaU833W0Zl
e6TqyIPtAQyu2UzzRm/ExeqO6mT19wFtoFIu9BS4nBqYxA0lYggDQY9i4u3ymzNK
b9A2ahas9IfE7oq1HBuf0/Pn/GjzP/5uZjEvQSSTInCv0rxYiwuWPjfLbQjbb+u5
jBjnQleBAC5PmeSeXhOgv9udd69qabWd298K3EAro3apret/EdWaAz2ocheCbCzH
QII+EKbnBEcGqwbaQ2i+SE5OVzfN9FtnMwGeOo1+nGQW8X4iovvNaZOHBVp0MAAs
DI8Yz51v/fl9IiYBj7ygKWGXp1Tsj0lAw/7m8RrYXPFdycI6i+sQg0hgTH8pK5oo
hik1jaYhaZ+YvXaW0xSugawM/ee9WADkJYkm1/htqOiSt36w2bcGPb5GIyMrm1mo
2TC7j64jt2t/I9zj7M7bJYkyxzOuhORmiS8qvllKzelJ6xMhvweT7fAD/FrKWYxt
6qmiO84RLPmfpmJRiYxXv16W37tD8UrYr6E0QUc27wmBZamhl83U2xKEqqViMXst
6ZLvpN4QCEitdHrNsQ9NMIEvblEBoiDYPN5btsmyzIQ04dCRSEfLizmafWjUCd41
m9BiOxDjw9Xxw+Od2B0Br2MSGscNEuyLsYx2l7J0xJH8GSb98ejjOm1GoMIP7SaX
KzeoeVqdk++TkDWITzk9sSqVWRwoz4+2bDuDLNzZCASq/Z/kp6RVPNEnpkUiwAHo
N4L+4UaUNvCNo3t5HnujhJRXTYXi2V2JU+8hK2b1Q2qB7nn8zPaf6MDFu7NLd51i
xjhZvbH6dxRzijZpV0KQjnOG32qdlOMN9CGStXtJi0SrMRIEFsiIyJG2Y0XQzwiO
hxKMApHnctMW8Q+dITgmjDVQUVU5YXX3p0yPgPKUKEaJhLRHQ4gOSzD4Oo6U1NUG
Qti4ay6mFLvPxWokToEVB7tqq4wOy7+JOBI9PCUwK6Hfh1z6/sNB5pl7wPY8N+Ag
MHt1e3PYy0AV8SlFmKVlOIGkfiXxdTgxKd1RhXS0Ct70eHnFqTpU637IHYP8Q/d4
a1EOSdOGG2jZcac5HC6ROTgxgYWexvsS9t8cHWdt9uqOb6n4SopZDjLegqYHMIIY
gC93x7g24OoWoZtSQt/pILP/2uUyJouWQjt5LOKU2JcSiIvVP6h4232NKe3ktQeV
12c5m7rZXOH9ATP+DsNRa1iz0EB+pF1sH3ZTdYgthnRk7zKE3zevOYrWaWRfEE55
ADUPKleskRFn+dzKumRrnRkbJV5JrLlQsdnggzDOU9MOZ9aHXbGoBNBr7Y6UKZ82
6CrSu6ZAbpXyQ0CKGWt+uCoKtamTIDV/UjLJUSfVWPnVNPJhuK9G3yjTNISZ5EAP
ay+ML+ZSMD5LD7jI2IGs5SjZra2RdXCVeiZoZLn1MozDluy06n2pQweWRohLJA8t
xGCWyIzIXTmmc4dREPXZn7UjAhqzFAxAdOOkr1/QGy0d5CGGa/+GarqFcl7teh4m
2w2Gjy/SB+M/z4CRmKr1aw1RwQ9p+7zXf+LosXLUe1pyrPyowKHt5OW/5EXHrdXC
7I9vn2hb2lw3r/3gRlv1jyxZPGOxnRgbkxFnO3U980OIDiAU0v8koOnsHUMsPpS7
efGpM+ARVIRpP7wxdA9LsVak6On4+/+P1Qb+bWO+1lndakj1wLXUgVvQj+A68ryV
4jREDbik3oN4d00+QVUAA/EFUFoa+2laNdLc0g1JSaNpq0aRQGZIU04mNzAe2GNU
XH+slCkuR2uzFu0evXeq4djQezsaNTIRYtj5lJ8RB90cfE/H8brBHGdBBU9hKbMm
1di4+Uvllj/MMsjejtpASGn/J6dLCld4jdib85g7LY140u5jUyAGxa4ZsKzLngwT
lbB+zNDyG4vJ5JEJfSihK9g/LVgANiAkiV/TfrOyapt2ZcaDplW55nAGkTRjx0KY
j1l/lhgH0KU6Piwto5oV5WiV8WoOVqPjuZoVyn1YiKa9PXRqhwTBvEvS8eisP3XR
lCiwxhDnwncD9ckcptgTRv9IOSwqaK5VMGatwyneCkb63A4eh9eDkXV0/CIvrHaI
p7Iu/tn3zBFy7MbXc0ed31KUaH2rt1kIcHTWOHJsUOfkNpjw2YiBkJnYuZX5P0+N
QWqmWmGbojKc7Gpl8JViUGyXxS84uLcPQifeJbUUuh5sg1Lk20ptbl7/rUfBVcXi
iXhrQ28s3XB+1PbaMJuVIGz3biDVYrsBsW9k/X3gQx8ohX8O+GeEIJDXlmgjOb+v
CiqcebziDR6rkHjDLCU3AqASLShQOIPl+wWlbMMqnz50qr55hNVFSBfp5zhAeD/Y
HpeACEQFbZvv1qaOUe/Y91pBncp46HECP2R63k+7QbA1YoctXrJivFbpv9qEpFmx
y7QH+40V0HNdOeTs/PyoYV+KZhKnLpWkzyN4CSFeDCeJP3Sy77MvtCbWTPzjov8J
E6BE+kgkKSb5suZgG0TM2JjJDABHuWIwLy0mX4oUe0ISFPmBeA7RLKOr8NUM4du1
pYx276wz2wjtB6/TwE339emvA8fLH73EIpw4WCnfv022/axQ9WU7k3i2F+5hCoN7
c6pdHI5dChqcaSHYUexg2k2Tb5WnfW5aS0pm7jg3hkOL3D4R7oHgG/Au5+9nxD/T
MYkPKx+Q5g+QJpYQRIqvQL1GXiH1tYTNGUO45FD+wfY9RbzHnCCvEG2j+RmEPmdp
4M1/pN2DRrgjHPPVVzITDkkkmHGmxLYqh+8EYZoxNpEEcr7rUOcWFhPaQ33kGwW3
bUeSSLBUOtUyNAd7sWBlg7CZMTWc/34fNiB3qEqTFXLmzVVjfQP94fdYAX1KNlUb
O8gLH4Oh/IhsKEUN93aF/W4wAF6qmXC/qoStDEsNMR8CQU7ngzMc/mmJgH5OAJdS
e4b5KNxEttWRs8qYQR0lO81VrViHXvfiwiufjgWW2WxJCo1pFhQVFz8BV7YnSKnv
rbIKDoJbFy4qmse3xoQW6a3rX8lUrAXx5PziuCLz5eQdsXUAj32BoHcmSCchpco1
9ys8Gjtq5ro/SmBCatiBXNw8JSk5Ep7VwopDK8ziplQ7Zfxsv5Ia9/QBvUurbfOD
JJ2bGPis7g18Fwxi5XtMu3bwBLybRle69Ly8fI+Yk+4deGDdm0SObMmnOFHHkw8X
LDPNbDN5+Tnx5kHzj6wch+6dGSvb2WYmvglVoonQFc1R3ueEp43MTXX9ro8+URC3
zYBXi3HrPrWOgDaGhd0WW/FPAJgeX9aW9WGq4td7DQ6QaRrWxpwWyqvPbzFenOnk
VuyTO3V3CjinfXQfG/O9es69pzf4yI8widb+BHCHs7oiuG/LhCI/JRa7Vv6r0yho
Ft/pS11t2QRMYP3iwVS9qz4S7ixVHM55mXQJrEDXUCki0UhA36Pe1fLXnr752xfs
ibKG05DyVtYrUkwcqJ+CKGR3Sdk28M2vPViuWj/HqZR/beEYg16xHEw6uIvg+fPN
yDr33VufiPa3F3T7a4vVxnS6Bp9yNGtR2ZmAEM1mbvMAIsB4C73xXIasKQobUtBX
ap94CcZOS/vPdoqpDlciq+aRMwTDj9UWjgaOMVJIvpOst1P1Lt8ATr6cTex7oXJM
jjkDuvbFqocnZl6QI//MOYeajqVSzuz69st4W/xf5JnYQG+x9NjjsRBHZwcGRDp2
84Jwbg1SSRefg16UHUxHznb5khDsb1q/BV4DY/YhX7TnC4UPXbAoUMZj9kYPF5ml
M7Vn2at1DE5DOnKmNtaOmU5xUh3Hd8CKl9iGmD08cPGDZxVVLl6tqAQ3DcW5GAAi
ED7eA5/Dm7ARHpXeydpT4a9ixpfUidiLOF5Derg9Fc2B9UeWmOSk3yu7GsCaHwyS
XfQk9zQ3h9g/wBuhVZ0VH1pzJgsSnoL4paYCrfJYwfbbEZQBn5TN9+FwfaCkNYL9
06WCOPzl2nL6PZCM3HeinmiOkxgdPhp9LeV3h2LYj3fu2XZ7U3t81aW9zKk3reMB
cNJVH8TfszcqGT+2P8p2xLxDgItkwuTb7fUyVTYIEfbM6Zw2vBXKmhTzx2ZNifRy
i8zpkvWSiWYr0I2E1CZhOA7lqzEwCekCJXNxllAd1tjPaJEm/NgYI5SpVUrOeuu7
fYiC3IuDS/FuoYR+x3K3rJiEGlCaqLIG5O6nnGVwK1dvB7/78zfolj7WuVQrs96h
TuaoyniLGQh10HV4ZzxeCYsef6pP5SEyEGbuLVPmTwXoPUWHxMv3lOrxix1MX75m
jiTzWrEtV0qw2P8oPz+4mm/iO3TsKjW4JqfrELShxZqAiIS6PmSnLAVkCp8RI8So
iIen8kjcGVJcjLFvh0m6dDPPGQ1WT+F0sTXDuBiOHBxzrR5yYS0OLS8mAIevCGcf
GG35qMArSeYlQrnx/3s/jJdvPcigi+G/liqUPjYXufYD4+4ymyFf1guGoMy/m6Df
DJeC7WGmlroAtbO1X8sahyy+bjrrOyzSONrDtfBMLCNqmWmwALGNaIrWhjy2516w
RHK30n6v9f3CpPEYfrmHj635ivmRW1G9FYd0uogc/HxONigs4VkDH4Ze3IoC8Kh7
QqExCaaqmJTqSeC70/1hqaziylBtZI5DatmEkR23RjWRrvyCiyidkT8M4eg0nc/v
kr5UA4D6bMCbwR5Wuyxn80Q/ay/E+dacM26wDWoIUzv7HUKIRIl0bxOJ93OPW97j
7RhGPTmQyG68Hi4ViJSfpmV7jhh/sB4Dk28h/vOG3WxqbvoVD/CPsuRUsXYiNLyD
YZLSNPC3YfQ30FL05qm9jBjbrBSPuCQonA2lEGUPeyXRhTaTTQEODsvB0iITgZoQ
u/plNPItj0EeFFCiBZR1c3dnvxyurmD5BbhFwEPXOvUAzcMiIJv9mOVJPEJf3ayC
qpRIbZwQ+dm4ar0zHsBMt4ZO1NWXKaj2pgaeFrtSet6xciIknsda6MkNjYLL2HhN
deuwKblYzZnFdIimsOEfjJCPWO1/0yA4KKfTCJuBaB6ieEOzEfX1DzTJnNiJyCYg
8BcmmRmRdU3QivIPSlkmPPewmYaXQjFybOJTQZfIJcvF1XKYp4yKmb/EO1xnkSRF
0rCj75245KFUnqkC1d9edobqNjtcN1fIE6PrlLrk4piDjU65+8D/fXBHM+7c0jXB
9U0jj9BqaDKsXke7vx1vrcm3sOrJwD3LspzUeWIOPQ6nhewuCdT9TVNfF4jDy0f8
IDSam8q3+nGGZ8nvinlmuL4HRANyjfGt2A1/9QV3TRBkLP0nWkOjITZJLagDJGHW
Tf5TcjAExczl1HB+pt/TWemug6WAFv8Nhde7PIgvWA3sPXPC3FLI8O5HubjXI4+h
/BJyVmtsIsEeC0JJlyngoiS2E40woe4COvi8IpAdz85so5PP5AiKks4mMrDdNfdc
gCIBuOei2QOR5MxF0u518Gnc/KWESh4zKeU132Hq/aEN6nJekszUYhcVDwJ9ZR0B
wrvpHAFaBcYuqAs9RnV1cm74puXMG3WwUFqgQvGnmGnJUOOewLSJHUO7y/5OhWqC
mQQpuom93hJCqmEkBINy66RImYuScnRrONjgHjGF4mh9V+skQs1mNgVXI/vxFo7y
5Ho4j3TmwN/t+rh3DS+qG0CT2FeNEHGIutw3Is1vOEcRMWi1jTDX34Xp+HVu6xjl
4gVRaQv9O5Q/QLIv49I1F6MtDNqjNoHsZgY/Oso9LmAc0z151VHAenQiueOk9HPL
SWr7r71Vt3eKrG/yt5yyS0uTr5++eaTqLYnbolcXZK40NXs+D8efCfSAetCun914
timKSga8AVlMLi378Pd5n+rCswPxVuGuL/ThyOfCEt30nwBITBq+IA+HJrw9FSwX
SdEwxLq5OsAyLPNKJ61b8Q6Yloa5zeZUweMhuVUIewFqGw7j5ifcQ09EKL4trFnE
1hFe9zMGce6f6cxsP6L5/f5krBPvwsvdN/OHoV+n8cvSq8BQtiKteOL/CAAADPYd
k2mVTI5kQLVxA6eaPlQXtVC4/JFcqAasOsDynITK6TtWTCK4yrK1A2JBtgsEtAUJ
rl4VY4L/+6t4rU6rpg/LmEW6loDlS/MjK/ais4uLMAzT6QVLVvd8rzla7l0taKI+
jaeeMYqtt3qXAa/Fv1bervez4qES5xkHJFSJTiIhC1tiutKEQMP2vIZBitybKsf6
+ASxc2puHytJiDKO6fReu+Em/reiD4eA00Im33KNFaySr2vr8qU77IA0prAntBrR
IDsaGh9HM78JK3hyVoIqTQfw3S+Md4hnYLElxlcQDtxiutWqbJJy/AxxHvq8zrY1
wuZZNJiB1dhR8QK/HUSaExTfhtzbq76lTKqXsgJB58T/pNWa0TVkZoocej3DKjaO
Y89vhFOhZNLHUknvPI+VvXARRjX5AFJDIpXf5KdO8IlCRhmMSsrZV4Dt3JjjQocM
mUqaN08sz727ZgbPnLVoGRJ0JL5A7/fThKiOS7IGWIFx6PtIK/j7cPmD0dzxSKJE
GPbIpF9u+Gfg90fferju5k+fshfUGQ1m8E070I7pmq2OhmKm/CI5AMmKKGZ7l2eg
zjc8ZsvgMvNVeiXgw9QD3et+wup+3lnYms+rEHqY+WicLmzNKwKPQT2Nnz7/G4LP
L+xbeVSOYm/MmWxVK7F2ZmolxswivEkYSfZOMQaxWSqT0U8/+1mDwUvZISlHOEeq
4Qbinw9D0RYrSxAZS9NAeV05yH7Aabgdt8j3u4RWkDphDs1s6dyzmkxYEwCb42s9
oiTKBZSQiN6V0F03zRtg7uLjU0ExyXcYkOdlvTk+Q5xg9SKvVyHL4GzvfuzmVzc9
tAZxFJRJziFKXJb/dPNhseie0iPqohSRyy/c40Jgw/jhSOByd5ReSICkWKBRdtIF
HZN+LcOes7QSHf9Okjg+72g6lVo8UW9Aasn9jX1Bn8Z/VKqTv6U3yfIvI7uPXsH2
qbZTqO7d3Q63ffb2WI3EvKERz8e/J1KaPySqInEl2/Uijibb0KDV+ScdvdbOFTWO
mrfNQIUjYqGCGk2QZ8Lj9c+vBRNjvWmcwE8RIO1KiQDehrYlgz2y3LfzuDVziROg
to03TYbkVc3N+i3/CEfC2hspJ5rPVtl/O1QrwIB2rjdhjJISYh2JiOzVasNNOSET
jGKHqVb0xQWP8yITu82bwSoCLFVAJZ1O0kkHnTLuK1XP/A3qmzqLPE57gNr2GcBm
paeJIX+rchRbnxHWyUWuOf8RoIKqec3jEIP+2Dq5I0kaqBU79cwvJbEcTOn+J9P2
e/BZr+OHuMGWiHN0TCn8FTWifAgAfwydQ6aNaFDCrQ1g6bFN8UrvELXPd1mGwrIi
HH2MLBhjk32En5DynMicxqEC1zwMn9escQvkIzOPhGTyLwjojfbwhgfvxo/iUOU1
sxcsvw7PqVIoETJySI8BdSfO9c/ZAMkSOGUfhuYVhQzX0SsOD0Opx07Xb2K/v/q4
hsMoEwSk10jWR/E6XhUA7cbhyjim6YxeRVpaZfplqL4Lfu7a0z5X9NbkWGrQjwze
6pF+YnkuFyBrk1afhWgfZkFmUZE0bOrYyj/Yaij9JYo4A+Juoa1CzKr3V/oLC7ND
6MTYm+5c3xZgqnzwVgorLcH8EAqVyjk9kK56ZvFzZXi1CfaOZ+l1sZ03PjBc7mMx
oE1iT2twqkiz3Clk9JiDJeWWCqtshfHZ7CZLK7lwLh+e9zk+t5gjofX2pMgcDXOC
wbXkUkLtrcAyFiXm0eX+31+2UM7kscdGxX5sq51O1er9E7rTPJs2NEeUeUjvmCH9
Ri5S8/c3M4hcRp9WyY0DRjsqnj35HXCJWaiotltPCdh1+xRBskKYVx9awTd9UEvB
wJ5hgmpsvw5JlAEPrZC4puDUuSBTx4ObpfaV2rWERLhXXfitrYpwC+Sb8myS9ezR
QdJV9WlGmha3kQVF2zKOpuFmV3BUwN3ZlRMiZH1qQY/HxnMSRWxCKmMOFtyogmtS
xOOWT8D+Q7Ep0J12X5BHV2Tkl2JMONYJz0+lHNFWzZcmpKaU9tODfKPuqUyHbRZ3
6fnhbmqoEGxpdPbs1wpNqkht2WN44LkfZtsVa44boxbn9/3JcnOY8Kr+7LPUCF0R
YXcctZMkXMcoj6awn6x8UPvp6cdspY5ovRwseYC4SGZ33lQtsxRTRmpoz+e+kqXd
R8IFdwSpUkExP2P6ut1JUk2Q6vkyHh38eIjksSWYt6xeWjHJt7ot6i7slOv269jk
SEnmwDmbl2TxHPd/8v9aFuZKcb/Fl830iS0sLAvibUsdebXKw1kEeWgEzH7eF+IK
UMpUpqfJ2qe773YC2+Fug6APPnUxEz+SUJyZ9k2vSjeVHat0bp9t79RhEqB+TyfM
cCUDOpha6M7HkHNhxwV/dFgUBJGHAaIEgzMXe7vnnRfSHkfdX1+kIVKFEDXE/er+
F3vM5KxW9YztYVUqnv8ZbbVI7zGC/dOi6W86MrenElJXvthO0PzUWG/ACp+oh9ti
QFdhlkyxsQufuObyaF532QQVZs3RuF0QgQ6ghvXELLKJyunkBkOBkdLGNAew/Jn4
7K1sHE6Gf2mm4P5cLZ4UlbP896YntwC1z9OEI3s5V2DfiCv1wiStXOGfdF9+c/x3
mpn4x4W/8gn8EE/LuMTEI/xannw9TApVWmaNKxtF71hh+7nCW9EwVhU1rYl0bHpe
sGy7c97U1EJjFaxbpC3pmRyXUQMrLp9wnO6AvjkjhyCiRGBulEoz7wJ92jYTtaMt
h62cREszFkDR4e+0LhV2Sm2oELzTeb8RtrsZiJnaM7pwuCW2PWexYlY/h7NFCdSa
DODEsoTWK5uiwji3zaLH6LfpZpp3Kuwg1yM8k6c6o/U4PtD4hWPTfnsNu7f6u9Lr
Q0PZZQDdwnvQETMz55uh9DckppQ+3jLat/J2ql22hLy6fRludTheb4p+c4TbkoiF
8EngVQphpSxjn2gliEkxzdrNgGjE2/kngv16Qz6k+4mjfKN8CMdzru8LPB1AO1Yc
r/DTujZ/DYAVMUaNlRVK5CV0xz4t2Z1zSkV/DXV62KOBdanzuEr8a5RqrjJWQU8T
oHmUh6bazt7Gyi4znLjkFL0nddzPM/TwXZGW1kA/tHs8EFulNybqOFPxjW64bsYp
tPxrh7Pb2qyPNjDIK6Tori7c/jvsKFeBETSb5EHc6uwR5Pu+YXZIZ9tEFpGlSGlc
kVp9r4F+NXTYuAUIBTqpKpN+YLhY1KTdGpwzfakRhV3SuaUi/u0E7A0n8JhTkJYn
+2RB4MuWOlE9uHU1lg+43mPreYduWIT76Pb2Skf15tQYhSCpw3Tu7DfEYy2UNvXF
2LqJmXWzlCZtdsxT2Mkf1cDMYnELoBqTjyJwfTjHGhiK1tKcJ4yWhtAfOwUeWwq4
TqmBhqZy3iV/tOOOOVgOFl1RcF7wvAKwyNtm4+ujzFn5AquF9dfCG3SGaWMlVJgL
NxFVUtRnUENmQTjFpWL7KSFhEIwFWWhdEjE1R/tNAepsyMioBrPLO5EnlkbB1kW4
KCQ2y1fyhfgO9fj2yz9yzfB8eUTwzB2moh3YPTobifqQ0UggQzTaCIRjAk/bgTA/
8+xH2lkSlFE0gjTvfywL71Bl4uQRD4u2SyvjHoQy7lo/C6gW/Np5y2bucyT60tGD
3cn4T67M7kGG+MkF4SgoHEmTDppJZuEue7bGEe4WAnlGKBFNlHQCSrIGfBwAnkzf
Yp54ckb20KOnHSeGvbYDww2EchWO9w7e7kP0BqCcmSvXKCEabT8rQvs3qlLSH/Su
/fSSxooh8dKpIcES89wVEVvAgaeXmqvzcx4QMUIZAnmBq6LGudoGkXmlm1JeUbcj
tMvD0mCq5KiUB/Uc5ng+jsPsKnwOIbhzivXcnepu1TaZfe58eRIAPcOJj2oEz6Lv
/tZVovJbw+7a/FuNfu7kNUeNMLILI4BYDZ+uE1xQONUKCC0LbYPRtOS+xZfJ+foW
cZTYB04L9jk4k0otyav7H3MwxZ/DNRvqe8PaGZRiV204edGnx2jxdtIHJutGAJMz
7Ku1BJ93dCSexOZeRHDHFipIzrYUDFd7rDF+0zl4k71qoeClVBup9GYA5nbJxf5o
S9ZJhRtDxvQo6RhMZBg2yjv9sX+FcFVdbH1z3XLKIrb0MBQuutE4GCx5HBRkdqKm
kfuX2MMXzqbCUzzT2aBFIadueQ2z0w9pXmLEPLwumq9exHSK2qixMojX9dJ29Vt0
gbpSn0eCsrLakGqx8dwA9R8vHVc3xBLSfupeTVNCNOKf+ibLpfDNe20+slopdo91
4lXveNgforJkyRv/kw5Q+GINLsaxHJ8IJWYtu4lQgvJsNesyr8YX+8ctOPZKyQts
D9y5P7RVyDH7UxYtwBcMUgy4bdNL5UTeRCk+M/TkTK+NS1DoaJWEQDi2xNYDn5WL
cxLsaYpkPdN0CKPhkJ9d2XMKRWCkgzny6VzDYGYHtsgrrVYRu5VTh3S4wLilsiw1
ITShZBDWgUfPBAe6vN7xlxVSzHHjjLbiHe7rBbOgFfGVLbHkyis41BeORyjrxbv/
eGJ9AQPsLGbCRT8HC9jzbSNDq1RzLMJ00ce9G08lV2BeHGgNAgO90yTduxWl8WED
oChcyFl9XBejKySoTgz3HsHuFTKRCTmDRvZSg00yZvrY1PkYLFLhuL2IPlDAryxx
p0/Os1GHWIDv1DlcM34lM9TQF4uCtj+gUGKf2gZ/x1qf+CVEZcGXp12SUCAtajIr
RgsMk+lJC/OgYrD0+JI9iSg9ABhkq4dlbE8keunuFzzpOeqhBVwOm5c9dEDwzAcX
ss4P5xyEHU3oGxKFgjvhC/3VviId5eaglQ2KTnkVOiDA+SAJ0t3RP3mpUZRSK56K
NVnPXZdg2u+WVvjVavhHgpX8rhYxYiPN5ykcDKkhg5ix+KrYRV48fu1WiRdrX1lL
NT17JcluruZCNyxMo8BabZJwzpHZ2NttdB7FWT2tsbXhXFLq1YhffO39b0GrxlFF
6c+IAN+MalNNPuFCKeJu0arnBMqdoc5muFDVfDCfdUZYaSsC/eTHr/MnffX8oA5z
+Wf/qTKlouRdA3ysPVc07uIFP+5CzpGKVPNwH3KPqkO+Wr2pe+v5DqMFF4vSVRak
O6mCu4+bBksJCWzyoyO4miXq0CgMVTqD6ERk4zh8RwZF1q49GJtjOxTgX6jKFLMW
LXLjrXgwPPqwwozVSPJpUy2iiGmR9nnXVhTuoDgUVcMiVzrSgnQyyRtvQUpUrx9H
MDjWNFNvd/AbuP1ly+Lm0eh1cETB0vcF7atEUlTVK5UPHggTf0xVPI2BOfwZNOcV
yguXP94eIout16NPgeQbkrZ6/nlia1Rc+QjnJ/YPXPkepBgrAVb2jlCsVzR52VBA
BdW5kbDVnLXtbayv/qBbGtZWRJ84lMtdzOyYomrJ8R1fiZ+LILCBOy8DgJ78VHTz
1dAZdiw9/pU84izI5fFm9D6ACNxdQnAV9XLkvZw/V9sesn4mQ1l9hgfRR1MPnIGw
bc518lXeRp2Mgnvrz5V+YxWfBckfvdP+MJKmEYT2dJNtghChqMrJImFHd9gotgnQ
BFnZoWi4L2CrUtx0XxrC2+0TtpuA7trd48DbEIeT0XD7wZgajUkw49AXZiy5535o
AvS0uNWax3MngbizoySFJTpPl6shDufqg5Ajxji75mV/0s5EtOoxt+i/4E3O9ryl
yDhgz251B52e8cAQLuAKN6SSbwMHOEmCpogmjKk4+D1i+Aujbj/Po8o5gZVd66xM
WXUeU8o2DBKoFkIG0YQGpv37Il2UtVX57Mb6YYQPB+FN8vVbxIH9J1/qzyup+D6Y
cPtPRmcZt9W91GP0Lgye2Q3c3Y0Nago5WxRC0pAnnCMVuztesahGo8veVV/rDWqg
8qlTg7UlsQ/kyNpy1O26qlzbO1STeYwLi+3tszaXZz8GxWHFtovQU1tOiaYwS8LV
PJUPY2b/x+YM5YL98kakF+MuCoErOmN12VOr3yQEXTbN9g2FWqezZykt9ODZ7vsz
GVFbdoSxP5o1HWro3GSw6OGQ8noi+uIQqZX9yKG6/Gr5k+9wMlF8ZGX/FhD87Ra9
Ak+DMCu8ZK12yCMbdoSJzKhVyV8r+y2zAdShHeYkChG2i/v8814BTSxZSM29ZKeZ
S2SzzTwInys2cjCbxNyLHmLa+sHO3GrPC8HvDbavOof578dNOmCzzjvKb/IMp5FH
pQb84q5eYhIm3U2QqXvxfwtG2Td///fNtZg/ZGxrU56YszEECpPjOn8ag9h21jrO
cp/FXPpTi6x3THlHv2CCnU9e5DVBEM8/LH5Zj0GQ7rSVElGD0b0ftCFmfq0dG8JI
5z9c33oflL4D2ZFjKoJ452oEu431GH43/ZUdVqUsaa67yR6luPGDzTjqPcjLFyoj
5gyjXCV1YIhwBInK5zVBRdPrhgkeErt8OleNow+uk4TVISq0ygeHlsw/DYV1xVkq
A6LzSv78B4BVHYu1l/jLXUdLCIfwt8EIrnQ4/I6w0aJVDHTUQGc9ZFQygW1bH/ma
4u1SiM4cBJGxWf5/iGPBLo3TYHb9lxLUjKzO7QfWwIiqUbwDLDFvxM8Y+KUe7dVc
hxJVzmJSVWME5EHhaZ7NatMqge1XfVgCpnAa/4BMA0MOaGqEXHDQneMvidfqCgbp
+IWWWPZNahdT3ZF+38+dGMLDPL29609F8kzqK6mIHkXz/sjwuR/baKXRjfrLpmHQ
m3xMlD8g21BP8lIk0vBr8Jh2vaAgP1q/9/vRY5v3cemQTrMS1ueMztmRqiuGAJY+
DfLtLY/F8t8ruNfr/RTuglvIo69OAcZLBB+gNzkT0sg20qVgZ/1pl0y9zGK8cCA/
Ogye144laK523/CldPEyICDUkyLzZ/8d3z4ySXZ6thhHtwGsdWmpA75rMPXyMoKE
ObgwXGqtb8/aPXYJJac14I4iSGF+A/MeAyT4K/kvFKf3VrWS0WPAGbPJ1lzjyMg2
fF+JIEePWRnKgmdzwOvTKi8nIhXCYWySYd269wtagiV5llb8LJ3vVc6bX1FLI5lo
A4FOt/Xwjk1i1tBQXm+C7Ws73fKmOJ7pzBdvgxtnsqTlMhIRZYUGPkGALpid9hU6
hC27MvDVf2BNJTYEg6ej4xQOx9qnmg+jC1c+AdMIOh1yY72oXcVZ0HkNOm+3hthB
b6+AwnD5lkXYjagQPxE9peH3yO4X/DRCmN1qZdA42LLOtY72H08XDF2N5N6cslaH
6fu25fNJdZucg/LKeo7Uj6atKonv2Kr28vk/mhWcR+dupsTGXcduummBuZLVtWDJ
VtJryte4AK9uyRmbp19BmeMx41OaaKFsEVwOfsS4wC/s6kbXZDT7KZ5T2yuW3FQh
CztDFz4n3VbAFba56RzX8fi7tdVU5ETyqgpNxg6tjfaibysTJ/0PEIQdjeG2ijLG
GFbnDLw3Kg5RJp14mGj+xOlKxRiFuB3bp/mBzSvlGPZZIalu2kNJdoW2Ko44p3WF
Mcxs1E4v0fYFLqZsvVgophTVjAZvPPr5kImtAi2hIpwqjT8ZWdWmHm5FtDQW80go
95eponPGbxEJ1QpHy3oE/1kExowZIjNi3MAQ3whSjDgle1z2UB7HIayzuK+LBJ7a
Pp9/Occ7oak9eD5AYylmzmQYjj4yG7gFG7Osgv40fA29sEbLtp8xF6/EqZNQiwzW
dV4rk6v9w/HXuE5pe+MxrHJbeYBNbPTJUf3UNF/YPHz6C+8T5zPMoUopbi3fGhtf
CiLcbTpN3vxcT2xBuZfwaD4sVTfqDbNyYixX/oOQg25PwzC05LIFtzSPsJ0zIVmo
TsceUMZzlRTttzLXwFClHKQQYhsxcsSU24QMd3DoS8RS++yP4A1nE/0zsSGnKAv4
y2+wQHeS52VOuwzSV80mgNwXDDhwiI9TIhXDXO4145GEq12CosIvBn37b9Ehqvkz
X6nZhbcw3UHHflwPyG6b1/O8y1uwQICLfgEPbkkm8SsyXJ5ZugHCKx1YwQr9tmHD
yZb6HYykyV2mC1UcBi22q3URjujTV8KFtYDbowMW9iTRU2DMC7Xt3JiBifHn9OCl
FSss4IcTJPAtCvXwE7avHcdAKN6C2/h89T+FhEadsLJy/3wPCfkmCO9APHjYeoMI
py1+D0wQ9rNyTJchaBvUwx+wM1dz9q4mijRD9GlGt+CKmpZYXmAuAErIEN0LSNjk
UPpvs3k/PGUU2xhUWDiGFGkmoiUPROTeVz1rCy7IEam8wN7ROusmJRobGn1QAa1Y
6ywXoa9fTYqr4jshs4A0MFCRRtClciG2/HCf1ULq7GFvcPCLcwY0nZvVZ/QHJ52Y
mHLb6LZnxUQlmgkZ3pP6QKkgHwNL1HG/PpC5Tw/XZY4gki1S1amw/l7i6JhCPUla
tNcFXq+s3FPYvsQ65POTJPfnKUql7CW5hhYcqV2GmxNUGiJRRo4xrzq4cM3J2obF
sKuaxM6lS2W6h3ykTKjz3Ww8zzY4T87O7+bjKepNv0qpXdvA1JFtrLzwame/UViw
3D5ZpQ73+LvuxcYsLIccj318jb7C1wP0O7r4gGbO87m3RLQAqlk/LWKYO9slW3wP
cAjjS4XMjeyuhHZySiOlIjNsio1gGo0gM5fvBcjGTx5kAnspjB/9CR0jXeq0eCXX
aFXB42qoB4wXNqxk8tzmGoZSOxuWUuXM9VHnDrD2djUbD2QN8IVTCsTgn+GBq7lF
QUlG/4TemOD/+F2fzUZWezJ8uVZ03g9PwFNDHjpNSNZYAPCNBPMOQDV3yCdvmEi3
wxyGPlzEdjKXOrsM00OL4aXMafOGVe2f9O4yaYiMKopc4KlEuXt8ldAhh1tlCtqR
fzaRYNq+PdqQs2ZPHkBrGlabp9q+5T86kX0Dr0i+jhrkSVDvTwhRj9ocn3oypl4/
SessCyRqHVzlpbAE/AHvXNC11MRkXskNt+K/zerckwIY9W3uzlhqbHJ1uRTqvmRm
oo9tC4NIVGR0oqIpq2BBzdYh+3rmmzx4k/kmJVmX1stq1DwmdjPhMrd4Rhtld0K8
q8KJsj3cVXqFuZTXNYeFoE28+Abr/1q8b+DLU4iMvK7r38nwkBvIigOh1SnGhvce
yQoAKygUF4MX3f0hIKELwNVKrf98atxndzkGSjJavUE7YHy4b92OXxeEqOFhoYAq
yYVhrxYpn1aEQEL6XMSG9P/3gGvV0q2XMkHzCJWEfblW1MbfE50GoPfa7UoqLakZ
bf+ZzNZo68I5hxqVf2J7yZqm2dLwQacPE/pCnxQ57QazO4zQV3TPMajSPcfyA9LO
sestk4MhOcbgITzBaRbNbg79GZk3InWrXtgJNGFoOHBIdg5PEux0v4DW4g8psKRX
xjaTe0a2LyV/smgfEl+Z6IMCEcvU7HKACj4orhiDsSYcuXEwNsy8PeYJPuloIRvi
u5+b5BvSI+wL+0rNR4oS2jbNRkHbeKp6UKwdgzcsfeO+pqqsrE4/UIoewm7ni23P
8Kqfu742tBA/zdJeuq2bqojuJLwrqJiLGNLl9pTl8CU7XvQTecoLX2eibQsixPJ3
KqrrbxT+ZXjCzbHHpmSByJbgE5TxnlYN+Lw77WXVEsaQPZ1XzpGa7BN+kdDvi/RO
GwJlecpbhUPphpMtwhFGuvvpzhL5arPxpU/VB4y/04mT4LeP/AsH7vTGx6+6RQlD
DgTE/H/SDGmMCSWiLlUJwgVcTM9bpatu7+LzYmiIODQ384ZzETmiZE/WvQLusG2M
41iv1PvGnguupncurJMkkf52sNWmTJirEVbCfGhtfur6+52IdCchwH0Rzsopi+/q
r6OsxNdfmeqFAwFe93GEn8HZ3spt8aFjuejFYeTw8977n0IyjGlQlwAgY2qpPE9Q
n/yp7yr5kdbd4kDDTRj80d4gNxbH60C5w5xrtq0EHImbIabMzVDSLE7BKrvy8ody
5LIfS9LWtdhEigc4ebmxAgod3Nd15kJWr/jP9KFyGU8XwLkDYKzjzCynltJUr4BT
HWDiw53yyc8HjWdZkTCYBRsXj93QFv8E3lQapEwq+koHU+D+f/521xzlKm2lp4fq
GfsaC3vwOso5weWftoynlPrOKWqDHl96xryC5j2n31/J7UhybDJHW58Ee0GYDRVS
LaQQ6Spp3sbY8P36BpF/CJ6ql8B7LA/7PUe+KHPd3aipQm9nxQMqOABTNZw8Rxmn
ru4AlGbXSDxmVuJBZWAdYucpoxvazwFR9DoY5fxg4Idt82RzhtHKW2YX9NOq7oTB
itjsb/2TfBinNbpPRrm7MicrVRq93dwPUnxTjtpBwH8d40ne1ZjrILyu/8htl9sJ
jFtjWsyBEIrFWtVQeiIcOSuR0s5L8UzgoO+rB+pNl0gWh4LgyvXmyiaWZ01XkPfb
iYcspKKFma0ZG1hfaKdzxWxJ00hg+LRGX18gclq7PZhwDfdfYUnhar0IbIxE2Z1N
TS1SnAfdVaQ2M/QH3GcyhZHqQlakxSoEwojYAMRkLSqR9mqsLI5NIB3LMkg4bD/Y
G6adqQJQbUJpsNszY5kNkE+MWf6myskIm0dk0ViJKS+htJZ/6nEhb6z457tjkVSU
B0MK4bn847B/KE0YE50h5J8hfOsRHw3/bNtFZppHlL2rRobCMa8tUTCa6XTnyeKs
g3tB+OrwKEh/yf76IROViFWueKeKZkITlB/k9/cSTGphBU02jYSqBCXkso5+nC1l
af0DhbLjrEjF/YW1zTVH3jRsSUsWuIDwGSMk1bRwhUHvrC92FeddOZIwAQFBagj1
jkDGA6QRLyTeMaGAuAVwMu+lQvVVISyRR3dVs9LN+CTptm+naP98ePOe/eMnkD6+
d/VlJGyy4M4vLBL39U2GpjhEQA37ANG8/C0/bvrO65sExevCpYSvvEXfGAyQ3qeV
EzqqBwrW3gejDBVLg4EMjzv1ckPs9KCP5cgNZ1idwatxH72Pknn4gUErdKbkfTKr
12VSPVAf3SJTgej1OZBQRyJNJNIyAebgi3y629vofGKbo3wT/4hkE8E+O0LujwtW
IytkzV4ZUj0EQPN19dDKJzhIk3ew4o+4C8wfcYksLrN1StuAJ0QyKjVX4GrlGlM8
0rQ9/L2nispB+WthjrWtbLPPk2BB/vRwFuN7XsS098Hp3BeUEKOVkZIug1qJxslc
aie7R6Xubm9Z0JLiab+WDQx2hwtQmvJs91grWdZPXsoKsVzUW3fK1TJTKHDgIb1Y
6aMxDMl1OGf2Y8jSG+YTPiHAq6X3GknKmZ8/PgvhNQNp9dMp2G4rpozFxhWTMzaX
+gFy5Pnsss/I00WpGR2/mflEAU5567DzpMViW70YuSC3XrTEfMlIRmXP0UA57tNS
uI3WtY78VX2jcLRwVkEgpKpRUhwPBp2TNIMzgCD310Xa3HKvpLxTHyUX/qO0xp8V
F/Tzyno4lEV9+5h6tiBpumrw3qHdYyNQ4RC3MRUMzwibGrYP0g0PDb4iTjI96bga
uzKujXVQDEYhIqXXq6/HAX/tXpUu4m0qOFvHUpe6MdVilLFTjoXRNKRXw5ix06TL
1CSXOW62HWSgJeqr6EkD7f+NkbAEerttCZibe9LZYTi2ftUWefqrEZTKrBq5wSll
jPajZ6ajfYTvO2Z2WMBSO1beeSTDEwalv1QDA2O9ZwKxr0oDD2g0lxd6WyQU7uEe
cWn8rftyB1WpT7Z4tQfTjsvnEGksA5AG/QsvK1bCVB4Riszn6Om8a9XYNTPvyCfu
cVGaSLy0tXXWA+mWo6lny8EZjbAKIeFZYnY1ktFUZVzlrsf2FmS53o+x9nZRG374
s0xaiJ2drU/S8n6qyf2A+EYjDFYgNZNDHAgEkUYYyefLXMbCSriqDpzztZw/GGBH
zqntZ2voCmIHY2ds0LSLsqJhEmqTN2d1b5/sVmYnjoH6ajChEdPVtW/kXgkojxJZ
m2RjiHib7MHakiey9H3UhgBli5KCNQPFEVWetqOExtal4MDr+81/cLtWYEkZywJD
C07wNjmeyQVRMtLpBGNu5UBzJAEsvQfYlAFLtAcYGoX4cQBu2IVkb8B+NrF5oGGP
sYUpLJomwUXa6koWIRSoxGFE6FIChDNm6/UGmiMZUWLs1lB9lzkUGmzpMKU+IYRO
ygkbh8G6fKKj0Jksqg3+wSN8yORyJJjEDn5TbaExx3XhY/2OdWqBxd/FImkwMRk4
+zcE2l8R8DFihza5kUX5tKOQRCGWXzB91sH+TogWfUkWP3Ojtd5K+z0bL3jaP6//
Dgxli7iEdF4nXJM36xtmWS7Poi4XQjYZKTSOUMzwrHIzhLOjXdQKNs2dZ8LDlUNI
xDmmUI9kncsrNlCQ3nlM2PsNJXO3qk22V1iLsvLpZ01SENcvLCLj6tjp2Zp4BjwA
PG6wMQcTecp+zwHwcRws8Fk9CiLxN9e8d0LQpzGPzngDmoFxDkSMiwdrHi+6pwo8
OGNAsujP1JhggFqjrvDe/F5uIgNZxOoUZMn0ApLJ8KDipSwe9ERyBNe0UVHlNmQW
JDkhSWLK4IEHcNgSl/JiSmwigIdubQ/nwzJC3rhmVJ92itiVZiUelx0NdKTWK6vB
3TkZb/H8yW0iRIlIa/6VetRKR2CrxMgFzfOBRnm9c4vzskFhhbVnxRIRFnnx+duc
hgQQGAWhhrfithxHs3QW9PNcQpH3fBArZhQLx/gHUFtlYtFCvBJ2P+6/wkI7UP5m
CWvDZC6/EXa1+7LJIRR4RMr+4vE18hZgM+W1we9MkoBdINZvfHEWl9dGPZ7yJiCv
PBVBgg4f3ermO9igY9Z3gt3ATYbxc4SMhQCve/tLayxltkm7IrFksjcL+z/UHOqt
XUgqajLCqomTRE1zBtvaTekxaw5gZJrGzw8cTjtxYx0VPGUfiwxjN0EUefeQObqE
l2LvzoFR13Fq6I9yfLsygZRPyudFlt25i6Qr2QqQdsP09umQI6Qdu1TxoHFnHHZC
Ou7076NdtWYkFgxOFBvWc9krhvY6mS6O9owyAgRuSC12jOyyZUsdNwroiPQTwuc1
6bAJF9fwu5/XMKNubF5kAagYJ1shTK4niV7HuoEoDqrl01iBjwgRU0rK8j0t35Jl
/KhmyGlhKxw6tpK478GQVB5sTRe/ytaMgekEB/PLgWJk907gxNIVZr3Nsvju08ht
G1uHJkipVgnwbNpY7P1kd0+ZXOXBSbxwhfInrDa2otkoImApqE7X33/13+ZFOU6J
uXadUI6K/O5aPwsdGTSm0uRXIyCcVkIh8sIpAc1y3rBW7b8572UEQHyZOmPgOzOF
H1e78wsr2vD36sK/vckA+VydkQf+jf8UWPysmiKJl3xcySgN1v7/uMHDurqGveK4
kkC/sXLXwZzXc+0AQyKQo3Ap0KXqOkxpJATWfbKGWljsfCXmj6cKZMNYBBB2kWDl
C1SqD1sdIlSFAgAUzefuipP7Dq3YksyTsw83MpdMjvuwUBg/A75uYGhFFsOBt5ma
5aTP+ECzalF46/iyjzLS5eC7dPhhkpp+XwQ1N9JvHsnbGhxG6Q7G826zdCl6qefZ
GnaM4QAgZdfjFvUbXpZtZk9jxtorTdPjKHrl5gauytDo3hVZxspOUHxfs7z3N9m5
9nPoPd8A486/o8BEmsJcSiZqsYlcxl+kc50ezndFb+3Ly4pszQceEgvZIK1zMAU/
jC1hVQ/0LA5e9E6RzxRamgrEksI6/p/LX6FF5U3/e3HpkMeJxIGM2PcDi74JUMf9
909JpHPBW/AzokbM33Ya0tEj4aKtuVZbctWNAL0lWpIP9/OpWfVBCknChWFvGKdd
Z91ShSIlX85uvBpi4rE1NGY8BXu4PK6n0YJTdblHKK5guQJlKXJ0wLHi8FjGfx4t
KQV4UI4yqEn6JbIn8zFF6JkBl3haT2DXUzcljPNaucevO1PV/XklOCziA+FHBkqj
zbuABAXOmkDdKlFM/etGGV4PIcVJHw9kGnHIN9ul9j/MVgm0vhbM2JMN4hsZCAYF
BlpM4c6hURsbE3IGgRjedVAdzZ4XAvH2PYIb2KPx6KwMIClOS+tVBnIfVjhw/q6e
So5N1797GUjCH8EeYVQmGBvWY5ZhgzofhGFkV0CJF2F0Kjz41SCitPwlH5Zd8IDH
39l8jmEb62FJGrXk20QVkkZSUY5F9ysUkGdkxx0l9/bbvuxf+2vtxRGZBAan+q7p
EyvbYoA7oO1mGTZNs98c0NUWDFyK2Xr8uDXxQTn9q+ydrtQymPgyxUqKZTe4QGOb
HgJFbT3Knx1W8/RfWpkRHmEnzJ0okZN10J2vB8aoDUpewN8glNglo/no5JzVh5wO
ihfJnzgEgPnx0+H8Nt3EM1+n9GPVUd49Jts3VWPWlVmSqQxDVCT9B8IA2osDdV7K
6/BJtIY9G1OcVzPb7oPByinE4ZV8IYCNoIWikAURklMcK5Bys6df5V8y8WmgNfCt
dbyliFw2rTLfXUsrHfhMUiWTviCaZyuEGJWi6mKQxIc7zbh47oX8yV/UmbHeEB3J
llAgJ+RXmmuXuiGcJKFbp4Ae/pzdVZ9kDnyso98+np2+NotRC3Hg2O6nJ3/OFdfY
QTKl94n5sKZggpMFvokQ52uXyytHP8fkaWk4FW/XzfvhdIQ6nuIr7DwLzKEmifcX
A21UxZm5EG4Nl8Aj9vwO9S7gkGJc+uVaU/NZKtY9bNt2yCjZfPkAnHUGpVt+QE1z
N1vsHyRAX1UBKd1RIEtRgKPEg0vbj7J6++hUu2htslLW56dT8m/IRY0sUxERJ3aP
oC/emf2vnFix9jVDR1iqaIJLIZgE0ZeKjhhdWoMFVJaZCJYPZnsMbh6ojDTa+CSj
E+85mma6/604Ey81OoVVHrcQnQwd76ZqNV+iKDzTHeT3oTdsyobZYF9eld/meEBl
QgFwhyPhyMJwAmWiUv3F47oCTczN2iWlU+xv02XXoJ/jQ89KwU6dbamr1WyDjCKN
ywPXTJH/40Jv/0g/X7WvtEXY6p4w39Err/cfFBMlHFVEJKzEM6uE5te5Pu7BnaUS
BySuJl4kX7lMEpc/ZndtHfsD101JwJmqyl1TSwxV7g/DF57+tXRbOwQh2LnZkGP1
KEjNJqKYQgEKCdRR3YBz9qdbIigaIDqFfkQhc6TY8/AzpoTFim02cqlyatT+V39t
S+5hytH8LCWdExG4wMYk/6e3Z1NIQMgIEtblaDjFdtILjaxtgrcCPGOXhaoGTFS9
spP799BOPfgM2eeiqPLXj3Q+bsEunDNM9nYhiEH8hzQaB6j0rIRCZLNbB+Yk9wzc
ke3LCQ7tp6fhXtoxKYobkZn2kIsKmj1OQlHZYR/4DqF97L1eeNceDUohKEdL73Th
ZqFt7ZHeOgdwSVvBJUsJC2ecG+c0KSssl6wn5rm490UWNDaTdwiHdvZqhFxE5tL6
FaQ2lHd2Uxt+bvSI2TQ+nrud1GK5rZCqtvW8NlGLsGwleBoGuf96/EpySD3beSmb
UKuiQpWfdqHDjajSe/lilU6cgCV2XQs2q2svSOwyroJUjzCqjSipXhhdCQRtrm90
FSjXD/QtXdNT+huH6nMgI4dtRjvnk2pgTrxThPfReRcitUns8d3Z5VkLYxnnfFMw
4HBAGAHcxP7kumIk8sdIoRMLQBqVl1Xgs8DOuUuj0xvLHDFE/tWZB6lYYEzJEFbz
O/auAX1Q0mRZzOOhae6Hu+Ii6PdN3kUrVQQR2aunHdHhUeMcQDMN3cZ+OHQsKzty
uNtyo5IH6VUU9f/0WhKjfDM1OID8LhG08g6HCvJw0Y+8GiJpEp2uWlBApRVNQdYZ
jY21M5Ht7DaqkTkJ3ZfcJzmKgYHGFyZzdjUzQHbceoR3ZJUyeqt6AkrKKGTPjV1k
nF21aHznUgZvudo919pNCS9jkJ0mwxDNLy+jedfYb/jwGVJeSBnpj2lECHWDDRdW
rDfm4WAY2EghqCwpnTwaVnwVPJt8pEF3F1ZooWgIwFun60DwxA9sIISb8Mtg67lX
oD5sNMR1vcdJwv2ifQzTuv9AMj8HkgSVSIrH2C5fLDY2fydxUNtwM/+iolqgEmGH
KxyjjkzAp51hC3f/5q3CpCDYesXmhQ2o/w66GSdaVX6DG9Cin2uu03SSfw3kn5YZ
67qvJnfVTbl3G3GmNpkMiBuJ//6N+OKSx6IS1oBH87lKcKbUG3uCr3Fl3d9ibJ+V
RSi8BfSWJuZRb2omO3Exle9Owxjlg6waHddIoIJaaaOc3YvZ8Zbis9F6MHxidpgn
KkfNyGwYqYvE0y/m3UdhDC80eVXGYuv03kE3Ff/uaYxv0N+sjA/0u7qIPe3eopZW
wBzaebwEiTATlyj/nEp++DrX+FD+8Py4wcO3T3B+L3WM2T8iRE4W1Gtm1ghLfVga
DokeoP4xT0L3O5jLcvtRyBoOJUrILi5mdWS/jPL0x/dOoGmTS3tSKKRRRemtXbqD
uX1BLkEeTqfOGHDD8vHo4vkEtsB8HqO3bNi4tcUzP2EgY9FSfKH3X0LfaBXNk8PM
ej5mR9gvdsYJfSmqewCMUCqdq3scmbRtNqzekIw5Ob3S8CTNysX8OcfTdUZsZPMP
hfsfxYHruj3CWQxXx76lWo0+bxbLawgW9jdUkWEZ6iR28KvaWCx6Ph/KSZs3fUPz
Ugd0WApLi2dYT4dUiJWiDhOzRRSCSL2hfFvkR6gz/jLdbHcaQtXUQTm5uTM3CTzz
cdaa/wvA9UeoAf1KYySayt+8MdDyrLqhyrWoonztUHIlG+3+ZI18OmcjaolhwwmK
5JPTPQFcnGM9eYnunzcypUzfsmkKSMH2p8JJgTI5KPgLDXpl1XtkNf/CxKa37lVw
hAQauE1T+iR9Eg4VIauJG+gw2VtMEhjtxhgB+XgRAoB3zKX931y8cS7NoqzBnQ2O
n5+z1kNNIPcD9zLr1tGoYDJ2ALlE71MrDuw8kQXaovd9f6Y647dcxSafPXFVivO9
lW2xlWMTlHJPRrvbWrrdL2wYgwzjPXcC96+GggRfBMDQCQam/D3IxDhxDJ6guBiE
9xhpM6o6okgHVwMMGQAO4VXhhsuDumXW5DMvbOZUh5I5lKqZu7l7iQ/UKIZ1XhBD
vrmj2ok5nVHBlcYcOCLSzz66AoujZLfE+jcxDfxHT4AArRX3Xx4VHX73joXbqI7E
bxI+i8h+bfOHCvDNjTCRl8ZkvLa4q9F0oQdeRsMpJaIZ4d4MWuRmVrQQHZAWHRjQ
f3t7wuY4XDXl+em9n0dJZ1xaAew69ybPSgyjMurtXii3Z3RMlhjClHP/WXUid2JT
cGVxbfP/rgyasXg1Tj5DKrdGeqcxZo6bjpu2vw24nsBAmwQNfZ1hzjx9WMQFMTTG
0tqApbrzSjZKmjfhDaPL7ZYfP19jVpxmvYMd9uy0V/b/ofruc59BeV5Qoepbkxfx
ii7nNzSXSjRzuVbffQ58CuloKmZh34lmqGor+xTaMugwU1OSE3axFwaCe7YDuIat
ZMCIXN+W46NC1NDdl0ezXlTlRhx+RXCPn8sNmcrX9e2HjVAjtI8AgBhkdv9ftZ91
OZG2aloyKS7ZKhGkmtA//2WO97JmxoQ25KZ7qLuZCDsZL7RwTGBa3ey1C70YoRbW
2Xqo6T0QyxSO/z+ia5t+/VtYNNtFFWMXIzgnPGaqleZdUAI/WGBxHKuY34ynZy35
So2SB4UlYqO39EPA0vqOvHmnpgrWBsfhitY7QyEZ3CAATym1FHaZmhzmDZrm6iwf
utSHK7LD24PPBPu3GZ9iJ7Lb7gyUsP+FLpCpTAT1F5fZLO8tcVgcjVB6iSGmphq8
HH/bzbY+PRYqlFOtN1KMvVlSlyxX9qTSXjO+AsUtQwoseKzkdfvbNvTWzSEDGvJ2
kX9i85/KuUWH3sRzVtxKNp7wdIT3RU7fZx3rkxizAVUQa6mUNxkV++nWKXDU/XR9
w4gSsoaFXaEEDzjBHE+klX/5BnnKVuqcURBLJlgiSOEDxoO9MWNZMSshxtSiH7Sy
QyyXLPsFhHO1lUDu7NB1H9WszkAtDskDGPcxJXuT+5GB6lpcjXc9cbWPI/Fonx//
YT53umBWxmNTBL1hIhCFi/CBB1DOTaIyjJIedQCMZHFWLHPU+JLI8H8B9FgoPFiv
1DvwinvuO5x8ropl3PYV7OaQqlnBrj3ePuRv94iNPrRN4VaI5W/v55iQ/FoLnPOH
0MoZ65Y0RqGCkVIoYv2pwm4dQT67/PeiYTEQwpZRcUUJxUYqwUYERz+vLzklmeZM
jRlaIZJep0JI+LcMGsuj85RbApS1onn7qKBqXGfwhK7HBpM7YFwTFNl1x0bi6Ycw
In/bhH3cS2dOb3l1k+rXOU7f3EFZHsUjiveXpos9XP75/ugpr6UXweh3WzyZwk+F
x0M51Onbw8gizptUoyiHmDNg6M1ZTWkxGYMmqXiAqwqvqoBRR4ntSMJ9CmGfDQ/a
iSM7So7t7yzclrEsOnE1Iu2vrTIVVj8DV6kD/P2hjZ0Omp3CSSo2g7H9vw46p9L+
22suJHPN+7yrbAI7CnDghpi5tImHiGcCapX85Q6iivbDgnvlecGiZLo+FjAV8tag
zwDTFsFLE3fhzvjo+ZMQ4Fc0SWxmB3TGd9p4BJI4xTyWDPD6Y9SQUI2F3t2Vu34a
b/fTm9JDXe+49A4gtL+iFpV0U/XUkitAWxBNrb6V1QZin7r9AW2cfmoCB0s1uX8w
vb+VgtSr5zuvzAt7BF+0evZ9Cm5OL9o0AMWHTNp58asGyiEGwNlnbr/WewcJn86P
G0x6LrMs9wtroQSBoSNDpVCLvn3KLe91RwQvDUxUFKVcZeD/K/1eVHLOwV6Y6/5t
oqm9ohAmWFqR53lerCz4wh32eD7wTxXw5zx69bQYN/UbRgLghGcRklVdapQgETfo
Z9t8+zqnegNNK2VTGx2qMJncKVQ9Opn6BHv64EMhknr6ltVHPP/XPySDzeyLsTyU
6WwaI1yoiGVJW2SaO0YkkUVdmIhjGQpnWpV52yi8U9eOWKr9Apoy88H2pi6fTZH5
aHbGlTlsQjsYyT8CIWJ9/MvnUQxc2BGi8OeL8FWKeXSJh3ENr1sAPlzC2i8LMVHR
+jNLpoTeKKhm+7kjMoY6cI/nKsyq9VuBJfDYqjJDJqd0O01yGptX8BrThVZTXqcG
9Amqw2xGxvdKBIXWvhcCghX8ZhNnpvxb+O/YCLsDxqRrIrl54PaSY1B3ZS164RUZ
UZ6gBGeZDGK5SCgihXRmvQCX+XJWxQu334kjKDNCg7OMfFcXuXi7TPReDOFOEozh
cc+xxyrvPFgbFNoJxQ3vRLmhGUusBuFzjp5iNPYt+FJ81zRdwxPS8t4Da3C38vwQ
t3ZmerUG/uoNF92UOeH+RDSbRV2goqkSYJJPxgMO5p+OETpCBfMLlYUyS5HKmOFI
6rDynP5ipwADubZkBItAZ9UYCuAaNFcPf+k3L6z69kCPV0tVYd1ttFwLJp+iL8Q6
swkojFhSC+e/nlkgIRkMRXNUtiDwyPTAzeQX5zfZBO3kW5zm9AVt/2sexVZfvryt
bYnIJ6l8/jaaxcBSgomFpzbaMWeKcY6FKDaD3JsXKdPBveGWscgGOF3/VrXX/Km3
U9H5rYy0S1M+EzJEeQDsCMOsAW4EkSzcs2iTQBMr5Aomq0xlfpClmkdZq6aFOB66
v96A9SHTsoB055CvMmD9Tn0S8dVdNHLwghQRKdZWgm0hU7mldPvGiaLSLLuFmo5F
nJiMWik4kaJLCKwxh0peXbwWbEyi+L138CPl/wxamPmiMmeBDvFhXu9b0cu954ep
Vynqeq0lr3FnFg7yn3oTxUcOlHKA2umhzoACWsVBlieL1q/dBbSGFwM1wr4+w8go
ASZQM6OeIiiAOZt/kCI6/2HMd+CcJGKIaV1lyaXbW1Q/mLXmTmMz9XHVWDyc0jgJ
7SCjiYkGTzJBiBcR57d2jUigysChnGp8/GqWAF3ru5f/z8F+wok8mFMyIr1Ku6nl
A2Au0Gr7kGqPzA8t33nZOMH3uiPq6qteEhZ7fQnXwOLlgIEZ8w17sFdNm6UvALtZ
KbvN+yKLHapGpZkecg+8X0SImVXyWRCpvcK2pTvxLMIWnB1mOa7RPVaDCfRVI+/0
NI0M/PudiFu9nueNIGbRCgM9Q7vMd/L77prPAkA/7YmgExSrY6igraHrJZ5tXyz6
X1gre40ido2dawTAIj2oNlBXSAhWGQwGrfq1uMI0Ae4OTXJ2r+9bMYudHuEz4FIU
nH9h1/UQeH36WoXmIgENiLpxkOOV36ouwLk9sJRIxdfqEYLrymuJXSkBbcwYorJE
m/9mWkosepr/7e2Ds+vYfWgz5AQEOMgE+D+MWx2gsNfsgSBPoIYujGIw7t19CHUb
zgXUip5pmXjrGnwaBaSM5YF0ZxCGuZOsIud9Ik18O2ViaP42cIQfAamGtDu70o6F
rtirTGDwIvPeH43wRLXF33djSdUEJJVgfnO+D0vG4cb770LWLLNnwSx8dVWqGoKj
4xOvMus1emqaPcolN9ESb1nxMHgLl8omj2lmqGRK/BcdeE8n9ByzhQ1eMMvY5/6Q
bZeArkrUv+bqW7BrwAKXZauKgTeMr5nxfLBP+w727vgmdhuCw9gjCLuD0dxiPY1g
m8AB4g3X2l0SXR7XNzv2c2cjcnERCkxBGE7emF+62y3QkA0GTz5RblTsJE5zQUfR
2nMOWNMdRlSne0L88/Qfi69ce2bIBCuGTyFyT2zmn266LC5Suf4szp71UCyJU3FH
3M+ye4WiH7W2+31/DQGpjkBanntxX11vKTGAy8PgFe5CGnitjbC3L5nRz91c/BPO
SHDWj48/ifFvmX27nT1NrT0Y/yowDF9c2G8tXrVfVW/X/kAHdnZ4dGcq7Y0h7NHe
600dvYyy1lZb1oktZUlYf0WA53GKupYwlYmxNFsc/vem4pVGvZVEaaa6+tk8fmLG
uD8xzC4c4ipX1upaUnVAyQZQEzaCx1nX3qJsfSSJ0NAiFL7+9GwnQ5vlJIJ2LXuf
dZZ5cKal1qdaHeAMfI0QlnGC5zZAXvFljowBx4/8dgTZesQPA8XzqX1XvnzrcGL9
0/VkctXh272e26ykfui89ixpVJIN4l/I/pusjO/ZZgA++Pa9Nxxs2SBIQFoZFryJ
5FV7y/bwXgMEBcpX8gs3ODjhBTGDnToq1xb8TmijAN46c20SSfJ3zo/czaoXqm0G
YVwFibbRNSXs0F7cP4WYoSVndsDY0y9KxN7sW7+RKx7Jfx1OeHdagqmNmWzBOjIW
nWwwrnY46pi32eQ8HwBt37xG3MKtv1ET+FTgxJKbqgGMRA/5GvNZn2FzYNkImmWp
bLryhVQjiv77NetvbAl0RHbp0n4xAiuI1zQsSSzhM2F6hePuRkq0K8ZDcjCMhIr/
LG/9WSWJnDWtQDdEyw2yI2z6CAHst+ac3LaZzppjrh9MZI1L3s6Ugw1uYLOvEuVx
RgY038IhOY4DMmWhruWB9F9/2Cgy1dhc8n3pNqIWdTqqvo6DgFhvbhDwTUARn23m
YVT8LGUkT4dHYYC6GK821SOvotQ8eCk+MJ0rC5QT8TXUzDfBrUsV1Za8w4Bh5uiQ
sF3Kgi6BYYjpd4y8qsSdQbDcXxNkoPR2Kh55TJarpDMdf767gcZJjR3t5Rhcvwuc
4IekTvIiK5o9+njAa5Pub0myDUD49CdChvRT1+S71KpqTj9VUB3UjV84wr07Jo/Z
26/Bt9C6njNPOExH1ThYs9TK0mtZlpagfW5yxigGyv61ewNOlYS1APsCZ7IFf1+9
6aURYIc3CxhoVuFVDtv/kOsOy8ALkR9+p7u0OStt3Yqjr3NDjKTPGN0p77YEvoCM
wY/wzXw+hBAHOXu+gjbAfpzphS38ZwQ9g/Hum1WdgjIAOOYfPiP1xWpTuF+H2rda
tOz9IBE0ikw8Bp0aM7rv5A475mdiTW/1EyaJ8woExJEVWGeXBQVDXPFj3QKg8222
nYkIUwYn8IOFyDXbw/sj+ddXzM0Clp60vyk8gpHq25eoXXsWd2t+D/Ku8RGxsINO
TVtwurVUiE/ln7pIu8RV0u6CufEaDhLC0inb3rf0RxpHeb2VkzZGnxCqIf3xCpWD
tkQA7PfQiPsoRknTaHzqbB6xC0YmeNZJ9XhjYNul+v9X6uC1ubIeM1ZdeCz0NCtd
ACX7rXLI1pKXDkL9adBvSpD5TCxfWVVrqsP8kSxfFZQUIbEDZGTmY4ha+P40Gs0q
Y5WMmdS3LpB/11v81JI6GJS36iggWSebT1EAjZzl/LJipfpSpC7y6idn5gMuoVpb
QR7FOhlic/DxrLH13JaQ12XksKDNc5Sq686FF4USjIyPXHCMtg5ITLDc5G8vSDSq
J7gTtN92DnNnoHNrMLVhejy7KzCqv7ZjDO76aqg8NWiN2jgkgyU5eV4LZsMsm8bu
HwANHJTo5+inlXfgQJorC2SLxv2JuwXp607WgV+kCnoxMw3Rcg10o72E54VgNvGI
zLZ9h71F9r7CwhrZNpxY0aZ9bjoC0u6f8t42J1l6BTJo7xKBZV73eyIsU9G8QNH4
BCrz0kl7iICjOnon/X6em+ot2s0yae2KUFxeBAaMLaPnaHdL/am04FPdn0vyJTNJ
1IkGIvMXFhS+ehn9G3Ba2YBH8P688mvzDRNfwJwFcqPy/nGTiPhZl3NQb3EkgYq1
JXg/lE90RgsP0bKjwOxRUuR3PzBZaXU5jDHlMJapTq+O0qDH63sRoaarI8wZHids
lSv+P5DifRea0rX8XjQu3dZDb1W0DxrPOVCUwaY8vuddsJKE3tobzPCnuNzd5rkp
OVa0UQ/vzOxS83jqsRwz2s0qNQtoXqC058pf8sXViCJOe89yQGlNVyRVJUUJxG4a
DJ8AwMv28dkSZ5srAr/tWWpwXe+t9wEhtBQObyrpv2zV8cXy13ciTbOleQuG+8mj
WPUIuMAfwkqYmpSj6tg9r+VdF871Cl+rtVN7sNjZWzXla6yj49lZJQs5AGISihd6
Im3CJVXFhFmveNaPTOdw6PafVZaeVrLFCOy3jRxhAwLHKUSCXKbtG1G+6/zVdE6Q
2M3MjkTkxdQVTZ8/t6u4e+yQ9DBFOWbmKxg7FHhl+RjCICz4oALvT6slfPvLJyRz
t23DdGlRTyRmLKfEw2Ln9dz98XjQYnZdYTvbfI02qn9UKhlynvqS7AVc61FI+3iq
RkEzg5yzsrU/jrRiNIun5pw4Z5MWIo4TNDGIXbtk+Op0ijUu3SwqCGA7dekWevzw
d1C4WyeLJAZcrC9HaGXW6M8exTkpUJQeUGOHzizpvZJbSMgWdC+1HeN5Zovgjt45
HrQiRDSQxsOh5wOqDCDQdxhxJo8yxkVv2XgsjKElJAJJyp3yycKlGQPTeNSqgyKs
XieYVM0r+Ki5CjvCixhZ9xAnjpt8AgOcR1K4KnA1euiMwMZn16RK0Zd0xYjS3n/2
Mqm20u2CC6Qms8XSVYB0iM/IbEQGImluuE+Z+QFdtxB1aNGCawp4AfgGUTSduqxM
xn5baJPfGjEBfuTVt0o5YrTp0OtU5DB0Mv+cKIJ+Ae6iZJDJrEZaCuIkmWXRJgeg
Cxc4Qo4nu5UYLf0CiK6fgjBycg7b3RIOIAU8liWucqmcPQMv9KjKAVeV41EYyfV1
LdS/FegmQeR0Ve9WUoQQVNvhmBr8k4902Vq7kQs9oSH1XnA/9NXekJTAxdT3iIq2
TpzRudEswNszS+WTuBKA01OZz/2bJfLt+1EzPnVriLc8eePPk6ZIDRHqTrA2qoOh
iTCseTB2MnMr8Opn83rH6M3exfWG21dgncxTwcQzT75gsGhkS3uTAtPaREqSMyZL
Hx2opvq4PgAoyJ2P0B/ETXNNATyPxabafsjf40zyhTTPQ3RHHLmG4/6HexO/GxDC
qKEeuaH2Ja8PyxblzJYMfIJo/tBAM1h8VjgrC6LsAZltE80xH4ERdYun0Eu+FfJC
xni/FFKfkrOAIVEwzToTh1FDH2UjhlzpWGM45mSjNuftRzUX0RoOxzAo6PXzOTcJ
b06rOQRFFb8IQj7BTlfarLWIjxq31A4sFotlOUW/ErE1/rpG607Ynvo/hhfJMayz
696Lj9SHxEtJnorIdWdzxh5IEeZ9Vrgf3z164wnRvXrhRj2sd78UYU6BlQH1OeHf
deqGMgMC7t8KSyeGSsJTL+evpZobwu2RbsXHnATH3KpbIZXEjfhvf0+DtJI08vwn
9NrWhNYCueUdDjTv1YyiaxvSVTYR8fOwJPtNgDHP5CC0PAKEuIqtCzTGqaGrm/Q7
eAjyWlgXZ5xaI1hMWoY+uMdSDsDRVmYy8sIY73O8uxMhtyz4mIsfBJeTq/lJsxsx
cptZZxolF3LjqJsI5XyiypsxlqvuLS+X/G1r6CEcfw16tAUhIK83srUdegPwXn2b
JSkgwWhcZzNjbuYPg2Uh4PH+rK2huChYcALtpycXIazCneavJqivmdzIFJnlC1Wx
DMQk6zuhjiSFE+wgAj4B/ym0KMzjWgSVz+FYk9VFxyvVBXUeZJqgK0BlJ0d1uhjh
as0+f8ERy/JKZq2Lu9J4R36S2rlJPrb0lU4pqwlXM6q1WJ52Lx0TOvr69+x/4OUS
evk+M9c5zRJtk8ctjCWLAg5XaLJkyMss1Yby1aaVOmfx8s6+Csof+AXYHWlTSzt1
+V+jPfbCMzQ9leNSZst8uvxHnShA++1dq0QEzrsvGmHHsq8PQP4MycNwrrol04QX
PnbaW1QwfI7hH6spqfqm9t0x46Ri/bXaI1HpRjE/JIgWX72QR3wHTzqN/7V1Ci9p
4l5cAKLHYfowsxDQ2FjwmEKGMR2RPgF4rXpEtROJMUHiPB+jr/x0KZLTY9gGekmm
yEYyrURroUkbGN0PJQ66/bqWze0I5uPlKKP/Qx2o/DZ6Stzq3/EwAyUOUu17jHXL
AM1GkAdEOvFfIU/ZP+KiBnmQr4q3qv+RcIsiRqmziUKsyKjDoYIZpnOhIBDaslZ1
wmHjFtfbCMeJ3lMIxinp/uMr3jQ8POOgLoNdEUF1KCCVoI4dy/3B+63QER4I1tXR
EvGG6J4ndFPDSGo8VZIkScNTxPA2T6ye1nvcK6FX6DM829wYlC6ZBkmY2swyoDcC
J4W6JHuaDC1wTzRot+wOOMy/jb743VqCWftKrv7DysFHbOJF9Og0Usv/0aXR1FXx
xaescNtNA6WJVwWT8txVHJtXoHCShP83Xq3sNBKvGjrF0EC4sawnqbMj1OYj4AFp
NPAkVogov8yUwoA8ghwJ2thPVT5ocKOqJ0eq5wxFq7mxZb9UCA9hL56sKiCyz/F4
/mRkRgi7NWYaN8rMEOKrECEMnYPFXfWLhviyw3r8ZRI11RNp5f6HH5PqQPklDGtC
gOD5cGu8SDHJMuFqWpu779oMbAx4wotLDB5qUIh/GokvA11Afw2UfphUptB7ULZi
/cZlWSYp3LH/elX40y5NzXmwfHZQ5odJHwHZTKZQy00VQwjJbStsqI6CT1pXvInT
7yKi7uMs3Wvrl7pL9DVGD6cMsjnL+5ElNA9oozbI0etnTHLP6KQQnuvyH5t+rUHa
yhlzuxcN/ssu1efM9ZotNxPd8rPv5dLTk8PZSBV8pRvLskRELLr3LS4oeuwKZpOM
fXP/ISsLEK7uxdyXNhLGsDOBAvJvCdtDM8j8lGjKM0IHnFneScpsJEEuiOaty4vF
RIFdIn90aJ5FRMxcW7crzjOUq7DZlNz6DPDOYZNbXqgXcCevodyyxttWFdv2nZsS
cGXkatcJf8l4uM70AxGJRoWG4vmeD/qqZ7ryM6VyF7mSlY34KDeXR8JU84vIwxcX
6z76mZP6z0HJzDzCVuK7nsFHfg+oTpDSCmzZrZEifyhgji6BJGjU6YBbagxElYVd
w+/67EJyNzd7EtqJU3trWDGcrgJ3QuCeQxHiu2zwkxRhIHMMaAhervJCma1vB0X9
3si9Sw7Xr+Cd3r0V5SSQEQqUcVkYh9k2N3i3uPjkQ86YTqb3kMM+ZhuBAEv5GXZ4
HlgTjIYpdLOI/47dPhG+psvTDzSlQqs9HiyUgbc6Q/mkRrvWhHjNpMD7QMFytRbW
UrokG7fH4sAc++PIZ89aqEvRkxtDmUwo/N6+CdleR9fYwneI7s50Kxapq8nTOMVI
kNRwaVECuolAXQfcw993YVdnyCNaNvnbRcrwCka7aFdl01XD1+ZGPvm6m3tWSJFB
nVMPF0KiPr5SkgyS/YInOPnnPLZE5dckcSzB6SLYGdd6hI4fqab6DEjMBxeTAhTs
hfrpWs9sKoYx7nevtSM513mGU7gBBJoQ5teeYB4cM8YaptpruEb7km8x1uQm2bAD
9QltAJefYDUw16C00NO2O/1tUuiiOEuNLEkNR6VlEirLOCLokhMWGhGeLo62GLSH
HFbzelF6O1+aOKB3QwuQr1z8DrY1DSnDun9OqqYN8WK7OMnTj6iB6MzTgJT008O2
/542FQz+1rmUXjEz2S0uz2LJDee+6zMW0+gloo7N98wgGnnNb9xqAzO7gzqNmagB
c5JdfHmSyURbkkg8sXOEp42di18fxuypgp2SLES+ASrV7IjOrQI/EMerEiyqxaRl
8QdVXBS97q8qbhmWxXxNV4jxO45qR0ZkBY6np/FpAe2fbwZ/7vQXcF6kL6w2f93g
BixTQTKTanqpjx01IcOPYTNOi7ekgTxCARsZmg3sz9kBWZJKLyjoV+y4vKLN+9IY
TIUC/1ZHwPkfOg+MkMRdwseaQEFejWIMy0YxBFUo0oav4ppGV2I+7kbh/PneZqEp
Q1BmejiY/6YUANnYuox0XVuPEmbYBgISWSb/LxG5atnCArSm5QR4gznuKtRDFeHO
KKU5qUe/IQJQDq+oK/nOdh67gaCQbZREbEqnX2ZBHirEkNMxM1+HLhTrMoEgi5Vh
TnfFUqsJkvSdivc4Cgxchb4Loym8TWmM6PAaclDZ1iuxkH+ClmiIJe6qDYF4Xrmy
t178OwPlRYJqc+HGrXQDCZy1xRcT1rhanUvpzt8YcQHlaMnRx30epCsjAi7YxZ69
F6ts5J7UrjwOnxqau4i43uCtUoR9QWZlak9UKhlZPTIt2lJ6C/OO+BC8OZJjDWtE
WDjQTGeQ7O5L6l4p4J0XOQ8bRswDh19AseNEdRnenDxXdMmWUOprO7hf6HKYxEhs
HeqQm9wTkM29qi1Wi1an71pWXSwKDOvdG8crGF9uijEABrthkQBAxF+5dEOkJ40t
Y4x069gc2+wxSZZlLJDB6oa8L6uKJQ6NIwwQMG54JCArdppTA+8OmFw9Tm5EgVMj
M4CYZAasQHC1M3alQb+fDe3D1MNK9XO0/+xSgk7koyT83H7NfO/bXG2/zdJ2Dzol
9gqrT6yp6y3JVlmQDN5EVv1LCqhRcmWAfSWUOwVwyNg/ZKWGRWGhmLFfTPv6oZm2
tq1tCgaeCb/hYreWEkQ+sPCxWs1Pus5PXY1OMIreipsD0niuje8+0cMNYZqufuh1
E9yuIO+UHyRmF1V3FeJyQ2MjEFBQ18laMFps/MbuAfYVmWS0VGRsBBXaDNMbkGNd
S3r6xHZ7UOc5QGeWYRa+8T1RxpLRLpEqCOLFF6jbHgstLKP5ccU4vbhCK3C9p2T5
47di2jmwr9ef1RQO+/oQrl7LpiBRC+gyCuq4oQqkDrJKvx7594iZknaF6Vg+5ZTa
mxOHdNkP2g9Z76uXZCGF8f5a6EmbQq27vVdiaq1hU1axVPIZXoBJKU7pzOHYOIsK
LGnTgcho0K5e7XqECMIatFh2BLfw/zCqcqWIVzriPOrdxIA3KybquNF+UZiCfpxO
TLbNYnvEyKXh665yxty4dCjVKz7COxQO94ooNihH5GrsdF7g/y462EqAtWDdvvZx
tHG8eNTi9zbgFM+dDOOslrHlAlQV9epK49YHsVKx7tnIMQs/fUjsKqJ8XzOE3UmB
mlCm27YfYxOVn2qDNHihmXBQ6w1F1fMlTaDQ1UTB8cU1qeE+a12mb4FiOzjrt/dp
aFEd/hRaW+7YnBv20+byNdlBpG+zXHg24Wv7Lnuf+hoDCQuLqKKjp0Ik3gNHzCBv
buyjmhci8nBhNN5ovfsVTBZvOFAygPpP7VgVqPdcvm2f5GNJcEBNQpD4Vn0voms0
IoMZ1/jJJnxPFrBps9ab+PNNA+uHW+QtgJ03hwSBiGOzT3wOuLWl1sNZsI9WoT03
Ne51+Makg/pY2LmbNZeBJZOLE6A+ENcYItG95RcDNA2r6ZCRkpNZlVy8akshdfTT
HaeC7UVfLF4uauwUzBUxPUNPAswUOs23QINvle+Y9HkeHcnwXlLrGUL72iKffGqe
lx6PxLa7JLXhzSLjL2ZHQOqaw6+yF5hKpRaR65+hRw79TkHrxmu0uCvqsnEjjAMO
779jsnhmyss3OsN7XXG1zYW1UYTz2cJhDy+fEYgF2jXc2knviw1cdnHZYG6kvJrZ
RrYgIqsxNms0/RQiW/oG9Z+4ingJFfQxSUI+0H9mQB6DkrInWJQitnPOjqSSsd/w
Ik3pt2NDt3A+lGtWCSpSy4wKQ+6nObKlNsAfk0zogoBya4X/c2rb8eD/JqZ5o7qL
BI1IP6xO0DPcQCcOFVdlF7F0gzZR5hnunx3zpE/bJxetMsDi7hh/QSDsl3xRYw+v
cCxc72RAd1lnanNU1AmC3+TUgTg6TPVRvImkkmGS3Rat8VHFkJxp2i2X+0ae49Gd
264fAsoy5gRKRAwuF9n1oOGTKBczrV2VgR3mGkb3CDwmXwJ5T1jnIdkmu0Yvp+7p
GhXkwIaRVN/rd1O9/5o1b/Ryll6af1OV6Kgw5b+Xmpcv/u28DhG1lVPdH0WOHr02
F3YOa/VVEFNtGyGhqeFuyiPAYTumD9xkoXDfyV4QF+UGs/ENYpU5Hfz4nxHPoLxT
3e4POBMZjswH9kipmgCXfioveInAVMJ/+MO8R5ov5SvABArIeJHjiMIFSdJREwSv
czDDGAZaKwvdO+qjAJBCp7VAjsbuzizBsyNN3HLMmFLW7/J2RbvdpECMOE1SJM99
9zdxGGlz8+EKrVGOg7PwICLT3J2i4hLlboQXrVeETLqxl52hcMxncGBGP9ZM5tXQ
NcxUYVxJhsjcf2bHAInUWVs1V66GREOcTnSzv7yhz6+jW8Iu0NxKGT54HUhlmt68
S5AS8/a/btaosmoZvxDSTWBoo8BEtY8R62nGtF4T5b1q1CevEPHTFT8pSFKLQ7uk
reJYdRIpSrN14BsmUouBqp7VDVmUlLIX0M5Z8uqfDaOjiYzDr9Ajl/ScAwJ6A4ya
fn7XMRYMbXMlIcYTwJW0IlEK156WebFTC4Sa559mElw/eubn93A+xSPWSnOOY869
lZqVpjgPgzPBl51zz7lAoWsnxu8aq8lbw+fUw6Ax4f1U8mZNn2wNUtsrosqzBFy3
WJfaS186VPOhI1TNnrDLpK9ToEaYQS9FuZdiu/BFk3KSoyYwFdvyWpC0APInHrNO
jyz5dwnS80v26JjIxbDBqdUEWpx7cVs3Unn6PtoXI95tQCbcF1cbkJa+ENUT3c1Y
9L5umOrP750Os2kKWEDzmOMw0YF/nWLrTILAbcjSyy3iUL6hcd4QuoQi5V+2Z71P
+7kW6HGB3i6N9BblRbBuPRPvnsfr6RiFXMz7bGlbAW1I5IeFbShckpzsbxqfC8cl
mNarPshGA289NlCpfAF476+n/aPW694Q4ma7qn728t0R2kk9P6EEk5ZUJkhwDzVt
YmmE4HKKr8jXYgRIpktd8ky+IN1HA8pZuigDO5SuiaU9P8jCBWsJJWcgzMW1iiMq
Xms5BTrPWWDV0XON5mXhfa71eaxVf5ehO9uW5DNc2K2dTOuEWrX9vNnp6IEIB6NO
gWWVDSJpJWfwUr4OonMx1dUfbGtR/wRcx0QJMKWZnbEbcavQuWJ3t/lJ6Ih9wkZ8
B22oYe3h0R0cYNzMvvCmbDnAEO/273MnPFgJ+fGS3AS65hS+u/2/JGOmoidoMlmb
LOmX0ZsEbqpQOhl3wbk94hcnh0bEk4/tPIxJy3DsQU2AOC4ieZifuVLLUoGVIyo0
dqoUxySQzU3ieylLMBUEwZrAY1qhlQ+kAfpxM74F+bvabD+9u9cwZGLrzwCc1qK2
zYyyoCHGx0/WYNcOscts6yvZD5hJt9ejMOlpywrLwPDw8iRIALHpDFZw1KEWDHUj
G5qYUHc7NSoG6XcT822jDDH4iveVLzuAcKcPJuYtaakcpBqxmF0sXBzuzYiQdADp
zJ221/Xg2SZJUGSHjw/IibEiVFt4USs6Oth3nuDgmUQ05/hSPjuBghIBtzGDxzKQ
PKCoH1mmD6uIyjo86DsRqbNqQdVubZ0UOTnnEy6sGjSBVGnKtSIwNj2v6Hinx6CV
2x3Q+/qKz7Quk6VUaxkZGIQF5QLL8akpheCnxfPWUVZrnQ3tbxZECz5+ioea0cKo
2rh+Xg7yu1OdT83SaqRyEuIgWPQeHCmZ0MbyyAMAldZcChcKLHA2nDX6LxJrxQrq
TuVJHjPzyCQaygGjuburB4nh4GBbZqQXs1M0EDEw5S+MrrAKqDalls44u3h9mnPR
I52AV+fuySXWpE3xc+e6XQAp3vs475XR5F/vqXD1stFAcpAIP41aYgCzV5lFNqoc
TtkT7f5Fy3pvywM2oiGxmb8lQvZle0epu8erXMmMsnfsNxv8R3N3XCRpNtuT+RgV
QBVtl216D3henbmHPRpnYbjzVLMBXfW7JV8tQt9uIuhA8M4j4cFD7oPlClHjfjdA
9Tw4oHhC71WiPpW+vPmvMCveo4KmWUoRSWxGUNbgrFRUULrM0RL4zZmrHvv+xwLc
0GEGtjgM8sTY7agzmiriBX4TN6yWKph+jLIrR04nsF4/k9RxkKz1qIoh/MHOevbC
eHKjbahq9dCM02xdCU3vjK4FzS1VwRNmiB9LEnnDjIQy+tdTWRwpzuu3Cpw3BN/w
FKZHO7HRI3zfdc7oTacxRDeeqWjBp/sSqm+KHvvu+Z77c3WleeL8j5+B+4Qz+O6p
ePw1YzvEWPWxry4Sk0lz8lwlgsoK3pHy+nOm53Eln87p89WZM1iDPbjtOTJ9wAsG
c3STRboS4y2nXEtBYnCoH88Qs3KiKX2qZqySq/ttW/Ab1169jSvPnNLUE4xm+Zj6
iMI9uacR+bO5UL1W5ouaT6YyTWlv7SufCLSdZ4BiCgBuJkqautXJCZNsq0i7pHcT
d1D9PvXqWy4FHDjcG1ULMmmRKbD0hb1vbiTlAAGw5Rf9kESuM+YCemUQW62lonQy
q+spTSPyQtKtyhDBTstDNBFF5TtChkR22UVrT9j3BmjrMqd0HvgKTYUbyqqZBhCH
gLBijBWPQnTNdr3mKqpELu7KEhg7Qgdz6cvq8aYrBoYQIYe/b1zAidya2fPLPcYw
TNftRV4MKA1azPY0pINVoL3AMeKuyX4S4LmOtQExA/RLIndgoJ2axUPqL6OhQS09
7/+nzDG8YCRfZEG0Gq6F/98M++/2O04LIy1RGr7Cvn3HyeUMGxnX8g/m4WfAhBOv
dgyT03WW6v2PIUIYA5/jzRircCCjQQfiKPYl/rMfKUARprVVHLbL17i71OZ1Owiz
7BqvXQWY84XGoNbZVXB53UoapAGSMA/Ab5PBvpzDlG+bBW+NHmUrBuql4mYGVUlp
8oKWYMse2I+ee0MfUqJHOQfzYPvc3S/MntVSvKx3/plr6E6bSiSQ6a76dJKVdHcm
jXNavEWSzEousuSfuDBGWC8W6TGlYS63wyBhRla8E2S0ss9fx28x4Se+6XK5rDla
m8GKf1mYDYE3fvbFV6TiGehCmKdAPoC55elPaKETVxPGxOBoyhEnaJQfoWsbuzc7
H0XqrqqAEeJ36QF5ZNEqApVxRBADRYx9nqhxuD5ddaLl9I3GXam92wsZRxMRgHFy
/7rlKwymklx0fHrWtDFgfQKInsTVXXD/ymsoBShkuCDu/4/HQxXnO6kvaMCrrb2f
0vPug5wKrT7imQ8R/TLlqS5KPTGoNd4AChSy/lidmDb8o75tQFFdhY/6QJRupkaC
1qkOysWr0mRSfB7FE5GnR4/51l9lsb7xoAH0VaGW7ZPJ5FOLPRofwy4Ee9Xl+u4N
TYpeNSB0HAobIbJVBckrbmgVEX6OS9uEUKCSkALuPzL/x4QYvsoabakHUO+pXuV1
1eaUu/cMrjWL0kEuuRN8MN+EeilHGorRJGbE9K1TGStUqhRRt5QfF7+AfeELYAvO
BOnVurjsga71EFZyUR618wNa62rCaNx73+pAAsAuFweM5D26Arazyko2KRrlLinS
fkm3Blf59WiBQMJYUMlWaEjKSiklrvT8DMIBjYtmLNu+zmnb3vm7LdYe9jrNxswK
MJG8GVttptsTNzzpRK2i5AoomNgCsmInXINireD/DIDezs03exaHdaqf7TxJwwW0
TQnhRccN+40StKg7oOn5f0h5z3mxO1MXIJaZZ0IacLQGL8nzMBHczy5GK4pCOvLo
5B7X4aRKyeGA7YUWNOZxz8UJcAlmTdgke1DXEGvMAQ/qH/jMqAIS/1eQ4QStNThG
B3UhwwRyhDBImT8x+9H0XL0MjoI4oKazPXjgcjM7gpyEUgfIAAuf1LR/560dzoGg
MQnHdXZziUBwKOuup4yhCjpU6pOy7G+71UFw4H5piOrg38MEfeZMTqvwNfIEnbe0
QAoLvbAomuSPvfWYMaiJJQNfBvKGJOGQWYMnqv6BQ5NuJxqp91gsrTjbo8vrqKwW
uBUIsEcl4o/2KnHTI4LBhGDzr+8gu7AxyIqH2df6O0t0ElUXSsOUJACdZlP+Vqus
4jeW5cHHAwWKQUmu+zT602FnUDE1p1dw7jejiVc8DiUFXVavVcUjWwst0h1C0kwR
iwBcngBwD1zNjd+fGFPB+9kuekh8OPVD5jF1u/lbWG70szkzQO5RwI6yKZgksT2a
stZFP/j7yKg8cbXritjy6BqK0GoV82PixwVsD3tli9DE2C8C+gutcNTQP6w/I0ep
uDmLvM6SznhuplLy6RH91/NiQ1ZWXD72ma5eMNcQYVVmL0bib4lv5T96tuM868Y0
+e/KEXxrNDZMsKpvLLXccjmlvxOCiLqjUn+ZsmiXb9vOJ62eTIyY8X7z1jOntdFh
ZBJaO+RO9G43cxALbaTgYhNt3JJGP4iYLY9rS8MtZKP6KmUvtiuaQOpsWNzEpF0/
+ygRR9vAkloQP2J6docRAUSka8SHY6s/rdbZ4YfbAiCIE6gKARNp70Z7cgsx6Ic1
uKumWVwY6Cwk9Eoa6IAteQjEQJI0htUD3Rhm28ZR5iTjskJ7OwFokJZOsk3kTnBp
WvhWm/M0J/KFO3vpF7EcP55FY+m45oMs96VI828NyLE3hAT8LjArLBRXma2RaLlS
8gDYlrRChmmr74RhMddWdgUC7N08mvnWztxhB8m5ttJk4XKUyOrrtt0FN7g7LOin
WaD0yuTtP8G432hem5jSVNdIne4y8SbdsevTtjMkhG0Sr/DY6Vsjm1/eg6pAhvPx
hLv2ihXZTgiqHJIHIKiJV0OfZS1tllRmXLDvjRdVi8RH8q2Yqy+ucXDW1jpktGOL
sxsTZj7PkBTW3Sows0YSoxMy61o/abQlEy78PCeRK8LGda2htYJZmsTCYLpK8Vcg
X0sFnzsRJc+u+KFLCEAOD3VYZkHgQPnInmqq1CxECcOhL/k1jOdk+GIheAEdnoAv
pqOimCTd7ar15Nyrkok4sgtIN0Sn0dy6pJoF/uTDk9LIXgxV5ffo6rnjqdCMauRO
2HCqKRnZhO1XxLRGnjYYWJNRuBdIFmjwy5WzQaWipI6cAFnCbBSDzTv1r7JW/WT2
kI8mJtb2AKaBSDJwO30fcL4d/lWgbT+XKBV56vrmXpUu5YLs6O/u6avnpQ25Q94q
l9LgPMx8CcTTsfb8qqFF3Hi8yUEt/gfPhg2qCuhktUa7NKRf4tu5Off785C0mU/A
HupoLHTp2AfYeCetX9JapctEa3Ryqvm5Ae18y+5pogJQPVopkQT7aQ0+GIz2W5t8
km7Bw/LLfwy25hPqGhM0pylAYgjw3kMjjFs8QeqR9UCkm6yRRebVVN68wyouL7VI
OsgFb5xZGLWVta5tr8nUKQpLT8jGPALqy+XR7+Wavv2Uim2dAO7Y8AitEIIsdXo9
RmFE1IVQTZgMtrM9Otb2SUTfgR1dDWbPveO4t2t8o24pv81Wjl/aaSnGgvM5P0Hq
/5s4frklP3XHIVWrrSjcsaEoQVvWtJe+TPd0vNWc9nu/IrNquk2fxkMCen6h+mcW
es3kYvH98pirWTIn7d+EXguMcjkgW38MtxsQSMiSdyE1fi9MTXE6LtQ23kU3CDvF
8zHdg54ae+PLQSZa/QBYdErxAmepem3zmaQsWrrQcKSOTDXV8SwHLr/bqxCIwejb
0/V9ILaLIXTFTdmbzfRz1F2botXMqLLJ8LaPbxaS2RSXUt8WRGQ1AqxWq0C4hZC+
J+zg7HiKC3W1HtDx9bnawxrzo+ZJtN3QmssowhgFYZG/mtqh+xT314utKS6pHNK5
mNiI3V5wS68tME6R8Xvb0ekYXq0HBNi0qcamCByb4TdKVcn/KIEEIUPqi0z4Iatb
JOgYjXXOQU4FsKvSF3C4+5nYBbhO0/RcrEGmRA00jkEC8sNA/tnTsqzj2FP5PjmD
J17C0dF2apbOVu05JOvHq/bIkFqBYOGbXxG+L0hm04ry/E1LCiCAcVByiWn8TEN4
8SBHebTrd3chJ+E6aS4tTAuyozigDkWHJKWxQof/Fi1BHAM6LB2KgRHxhc+iYiMr
+bsZR5m0A7EzNI4kuNM2/vfAVgByy28YWzfO2EWLs1pJdA0ArAkc74K5aknkKcmQ
txCh7cWomsSgNfk6KcqrQKGnAHAp4xroYE74QZqBZlFv+JgD0WBxnTNj1nFXX2Rg
tCtmoIG8dJis61LYohx5bF55Kcr/4/gMIgHLu1RCEeaqfO9A66bwiKAB8L9gDgEy
oxlzXkOenJ/V7eLxLLIMKCJSy1EyXhSGQr1XTwDV5uCPDIEvlp6vHatwQD6tayf+
EQ66WqZkIhYMIlwkCljhJGr15ufB+gLwahh6ywuBDuoKWcLbdifIBmEot+kOyoU9
AEVblpHmnyQB8HEI3qrlrZ8egaCA3jkYJ0WEhLPipIKH08Mt2cnVweIrXB4GpCJE
oMgv1G9nKhY7pUpcDpZ9CpqYRRWE1KoHq/qUg9qplxZOdtEmnlEC25rkLiaceiVO
P4hy/YHEV3LXhjBPQEFaAVnhVHSWN/D056JKQ8tLZcLavOlx22UeNg1Gbe1Dh7Tc
bA2aUAnmo9mD/B2d7gFHQLiQNnuKjmhrTpkrwwTIGkKXmztTfcwqRVoxZu381qS9
BtlxcI/4s9xEJUxAVK+fuon2I9eo0TeLgD+QnW2M1vnex4jiFR09P1qJ0suJnmJk
QYhVEAWf+SWAb735sWT3NIJLu9KgmbguRBRYYpLlrsy0FqPfEFROb/8X1s59bhwq
TGYJLdSf2va4I8HYTlh93YS2QHRZhX3Txyhkn8eP283nmpMKBZO7PHXXa/t2fJSU
Tz0xmVn78HyTdSn+OMzmzlsUX4ZRxJwQxzFpvro+xUev6MA8ohjQhiBao5Y3sW0F
Ho5k9CPBTcdfjsEeLkSdiwtcAsY5CHI/PTx31bkj5/9ULmCTscqYFXdUShUjpRcs
/UiOc0us0mSh4KvuLfsc3pKIxlKZuhlQ3qRvzvgSY2isql90cuqlxHrXb39ftYZB
WW08ZsNRsEGfk6otWaBlgvv1WMltF6kR4QOve3m/H+NsEXsov/qeS/fZvlDSSX2b
VM4d3dhP0/YmH2m5wpENBYgVOaTl+MVcPb14JgRVAl706VJclMFet6P96HVb9H5T
ncGVzimVw14PEnBwbia5LwJwXR8aKoin+qWAkLmKNXGKqvNXCv+4aIoLi8LalQHv
X5VspJbCMkw1YJnSpfSsnAaiU/mN+KQAirCXIUq8e4DQ8QERTyOhaS/t1lZUxoUX
NCWLQFfbnNgtbfnCEW+Jc18ymBk0vZzxV/AiCv2KRUCZtjuVWXmrkre6PLZq8bP+
2EortGj4JDxKJC1+CHITGn6NzdJgU84IcS7Sx+nudJzAmZ/iPDl8vk8bol86ANA6
FzP1XD/gUtyjazyQv5FBfIcqdBsk1wxacR95TGwOyAvd5pDGcbwZ4HnpPySHNzvU
E/dJKMrd4xNKA5bHpZrPGBYXMvV2/CmO6YpzH3k25KSl3XrgPd7B3UjnaiGzSLci
in1edEqBKVOt9ph4jale+UadT2ULZN30M5nJUG7fmUNx7worSllRy6tUVyH9Ryfb
rqcfxi+4Uv65EDqGe00epy8mfmwZ7yD7pjiiV7hnSaHurKTINu8m82bXWMRQdSHN
v4crb0m+JoQ0rIRU6Eg9EBbqFCtA4xxFHpV2zC0Wp/x8c5+UcvLxkXb21rSswxeU
WOOp6yFAa+nUm2i6+Zpza2I1ZX63Jl+MeFWCIz7kiSEBxa4UqCvGC/gNYwDCqas7
yg8oqrVVoKxVNWvFkBa10qBlc782+28eKCL9AgKyyQfXlJdRIvUN/wP+fTrO2/Mc
W5P+FBoLNwBsI4CSU8sXXkmboQTTeB080Ah4F7QvDqMUazF296fvv24/6B2vXDCE
d7pkY9ckpjvD9HXjg73HhBSjuyaCDyIadLqYyZN+7lELMeW2vdkRcvta5xJus4g7
QNERX3dR/sD8SlQ7uqYnBUOTUZ27AnmnprfNrvrWpaqYx2iZwXR9K6q5dXQLowQl
WlaCjvKVkxgL0nPW/BcC2fVnlWEozHOJpxeCJBeryITAEb24jvdAfkF7Jtf5znaX
Y/JEt4VRSDyZJKKMJevnpF/BD278EcoxqLLnZiJZoUX5VTlBC6nnRR/XD53eCfdo
3vpfMRH/uHNQCy+RXPihaUYMosjJs/Ghq7dxVmgbXKRBdj3URBtWbm/1NPwt71cL
oGQiBqW5sOAL/BlPWEc13KEIi0MRpqZVzaiVZlT2Q8/BRSakKpDgFrE8zssp7CN1
3dfzUkv8HYGvf/JI8N92gnOwwnouOPM0JMJIPctiRSuERCO4rgIvttVCrGANv0+U
Zg2IdgrleOSo5TL8o4GGffcU8/oeY3Ny9ejOMiT9bwMxCw17FsubeC9PPsywvq/j
Gs/KK2lUIXVDE6TyNqg45LK5399eeYqUA7p13YBExRS+vDl67EEX48QlIhF2geyW
qrbSOTiadYlpSelttY+u4aZUTKsFS58TQGeJbhti2rPeYa/TNgP+0iIyH9yDV9h1
bG/5hTFMxliXkCfHQ0/whHmfuBqUcF3VhG63NjwI72UKElFp6XxNmR/rAPEjCG+1
QoWWEu9h2VN8V0JFcuTwA9qlGbTtXViDCEpApHBMlYUeyXuqIz+m6iU427eZ8JL0
zPMM5eHHtN50/PDwbvLFLxR9R+8p15RwNhLbte2We7xL9lm3BM+KDolr4KdZToxl
MdCccdi91ucdTL+frqyK+NhNwf7rXJ7SHg/Pv9H5P+2E6kFRV/N9Q4Z1rlm6/5Dh
iIxVjBtPBPFKkmWU1AqoDhMu0O1muiB/AMgSZ0ddrkZDK4H212nztKSIoyRo9fcC
NFO4OYGvDcGvxPQBbh0IxS4dcBzmo6+B1mq1W83RDX+qRZAHoIkioMUxuTCDBtUL
z3WXkC712HDd1fWZAWSKMiW6X4/NuBVwe9Tp3sIsA+9gQufiRX6Bc8ihszo94AGE
uh8Apjz6eXfBUR2zFe5O7so0sFJGlrbI9FQGEBflTK4HPIgyDdcC3+cMOY21ujLV
T6ATFXKiXV9q9URGveNEQc7Ca1lDlMbMNf3JFQzjv5kFT1QwCpyEdfhSCopBdUwh
XoR5IuAPx+e0qN5IUL+jauPkVa/XGThn2JBxd1N8qahMSf5gvW1F0bvSlzVve+cW
gHJITiFMRuRdBDRl4lNI/jwGLNRqPK+ujvEnNn74wN1/jA9KSBwU74AhqIGQlpvy
XSzvTv+WMG2pSMRcbVtA6FsX4fxKe2mNi20nus/ZVPhPwJwZxZzWSOzPtKfGmRh9
bhcJCPqprmVSVaaZsSvcTFht3hCMgvgMNLJIvDTtWQgShVBWmr5IBdXDzOAPzNDZ
vvf7zjuX4Y5PmrkQNgbzTuYGJ/iwHBMlV9Hf5DJfHgh6ZgDyWwYPrppx8heH+1oH
J3SF+LQSaKnlewYE7JREzWfXW20cQUX3IAG2WTqTCHcIqXg8O+MmEA5jLACt1niF
bjUFqv3uKmeX4PHQlQmCDMijCkd1y0skLbPbmTxPneZXCj4qxPQW80o1yZxZinaR
7XWKVCFUkCS07bLy94ywQ0ZOU50d1G0d86An/WVm/vwmB0YBQFRmEOW87/rsIYbC
J/2lKHRzuv0X7lfVbXyHktIsEgggRCYZbDti3Ni4wZMWSfVpUp/fjHxmkj/8FFwx
4As53JhpmCQSa+NnrEBOh+W+fU9qDP15imkmIyh880KrKRwqVEoLjos0i7R323R0
WSXZ39ySMcp3INB6BdUAPLJAYTP93Mtu5K+t1o8pRXdl/JP/+1mOT9cSFS7J8F7S
+7rCUGeX3cu8SE7iOzOKjdk+Tg5yi3glfRPzWiLpNezax9R+EksAQYS8H/mJ1fSF
QP3lIy17dlTz1eOuezGtQF3AvWric4m73Z43/SKvJnQRho3d/049X5SbToPT/Pcd
66ydpNBHXUIDA4S0iXvh9luvqQxGAtoxkL/kyG3F4M5IHjxMPoymKdSsJ05CDgWk
LHapM1o1WpWW06gL0red4NEPMrIb8FO1WAdVZ9GrVILsnGd/BSUprYhsfX6+drPY
wKKkAwlvEf60lZ9UprrsWs6ZkFXxOpuJ+TPi+puYbvpqlv0cdx3S87lkMW4owXws
qnV/QrpU7IDJRSHp18LGdPSXo6rT+UzrBk6c1xWHjFBfO2fEttlHWjMZB57vwODF
5jzdzPU7w0jS0MjmPo2wWh8hFSrw2oyO87p0KvL0HImS0D46EW+ifOVrIG4D61mH
Ga3Gcvs4PWlSrKSVQ8XToyxAjfFFvmzDIooyRYmE8TwncUAL5kuNE2MHvsEs5vki
EbORZj1rTbDATntIB8syMFcjDQtdM1qLtXO2c7/u/qOFGplrKoLxPWQ1ntuluS98
owFKgaYLrYm/OT5nnnu8MqdjsRfX4yJ5+NbD47FApIM5lU5BqFXwCLViGppJ/p8x
yqiRb+rxVQna/2CsCvwZiymzmZotu9bkgPTgIgVdZZ9zeUBEZMMXXeP+BXO/gDbM
8gNmGxA7+ZixKanww7dw6xLWSX5LNPY+akxYTT8jRsMqIEESm3wwWyIVK4BYZHdC
FIg7ybAiEEF5nVscHEXe0IknJJJEUjvkURCAEuSX1K4etoRP9qRihme9dme2Nhjl
2cgPgDa9ogHWMvPinC4fElkM5BlKrDAk0tr69to9dM8Ipwmq/ilCGYS3ac6tAjOX
rMVcl5EKcduYYNjnwGJR2FzKKgF1uiyCbDNadYX2FfNywiYORY6s6ztWtOCftflQ
JJE9MK0IkYMEF+R2YOBFf5sYYYaKEvydPqfkLpPEt4hCTqN9FDbJEYDy9pTPfRiK
qoIITml3uuOla6Bp4Nc6mKsVN37p5fyi5ls6KgbBlvwyNaWhRBXbwNRiIyyNsrGT
8i5Kdk7B2i5OVavp+9mgpi0BpHS/dZOUhe4siipP0R0mQBHnD2DIr/SjfoFMdDZM
fof4SywTi00KRc6IvHouPgptgsgmuo5TgmRQXF9PDjM2Ss03jYJLBujpUKOGkG3z
Ui3FVkLCwdlEpi5A+ljUke1MTg18jl7zO5ylmrYJTCcEGLuyew3ngT69G2LyTURw
0MYpsFvWFESTH/H52IAgnozAcpMrC/9ySxHmjJoMcPw8Tn1o2n2zEj4SWu0u2iw1
zZd1I/zYZZytUtjLIqro1H4KgC01Iy89mfiW3T9ZnZvrj8tbGyN197fvrF8odQZp
FFWmvjRMyGh5GoRQImO/RaA59hrZypTvSSV88ernyuSqw5yIGVaSgssKnNZKV01R
x00vnc0SnSktBLkAmyVDQuD+az2XECLZe0uWiOuuDZ33Rw6M+jQJSBKYgElAqxxd
P4mqc4y3/uutSCO/UqoMLoTs5K8iZw3mWtnGT3DjQHlyIQCT9SHLL4O5qZJh14lB
DBKgyqTft8NwlAJKEjE051SvTenKaQFW3KXqG2vpKxqK4wPgknxXmUtIb7os2Xjg
s7MPbhAop0STU/dSM1139wxkXCWe3W2vbsYpN7gEcsEKNZxcvtJWLSUqPjsmQ5OA
P3W8TTp6f7WK3wJuW9zgemf4pjih2mrpV32WMCtm3J3lig6F8q+7MidGEeQ7Vhzc
M199ShdwMFlyS4McOoOMiu5qHywFvkglHqs0ay5NgF6/ih9mWMlwNPtBF+98BZe1
zpuZr7wpSHlEYBpJr4eP57iHUfe3AmU8SINEot4lR3fHMDUCY8qQ2AoLCsdEF/El
k4XU7PWUwOaYTAQj8SAGupUHMLRsTNKqu4kTVtKa+0FUkQ3s5xkNg2qbJ254G0hX
dD4CHIsiCl7A+SD7Jk3cW67hHfjgWoWTGqhoiisRSZ+WWI1dm9Hr1kPqQ7djUZU0
26XHaEx3t8psFjfrquWen5DBjmnqJIC3bESnLJ05uPwspi74QdecpiO8xa4BeHIb
sjINAFGfNDQxHBtx7tGQyXjX4VmsgfzfRq1Pxk13mjjqpMogs1pZXcruYww110o5
2nuNfN39UlnonXG3u2Hnws7kg7sO3FTIw+jYIJxboFJ0hADIaO0rX9Ym/hj4B2Xv
7jKTh5982WipvK2W+TEDZVSnsr/OE992Cbh4V8BHL2d7fYs0GfpLV6SBQfOVw71G
S/o/zcU5UYO/rkLCVj0VFELSolODrHE45HC2WXcIc6KHjXqvETiWy0vimNcTPv4J
sLpJZElB0L0AOZxq161fUKa3t8t8aKlQUYLOj1nZ2XQW9+BOE1VGDRMsHs9v/vqn
buuvSdMVbypDrcFfc8eBtGas68wgVKjJm7Uvp6tl2IZjpsk9xBzXk/axo8ZlxQgx
ox7+W3OOt3UVXfP0hywX0Y4ik3obaf9xtpybvNFzUviB/jAaXptTm8riBihlkNhT
FEYIngZ/4wD5ypBvFq0C2j71gougElklejHzOFxqHbqLIJ6Q1tdY+5vwsUh2Noi7
MgqUW3km5WmSafPuGeGElw/eoczbnTNsBM1GLUlu83+LzzOAEDbEhgheTD6UTqO4
cjI90YWRlTH3B1H2peUIctuG5Qwto1AHflBdrRN7kMupnmSxj21CcPYBrhhrt/8Y
qsOpBYHcjNwasl2K9c++AT4ZLOE/cL70j6yQbEkJZzeZ8XE+xKOZCef/e1i+EdU+
CANcVjATIJldmCsinlP4g5NNeHHh4e+ZMPpwz6IgeUBEwT+p4o7WJSmEKtxcJTea
7vDMj9Po9//IJy5E5j9zph8sBz3NkqJ0gDSBcRyRPctGpOMX4+bk2usfYDEmLJQo
MzWUlIhJStKeYtOZN8TfcBt8JSptAYx+QTsAK/rk1zW3X8EW+E960kHxld7CNNfL
V04Nz+IXc5MeeP8rijmPPai62Qs9csoUeedehByRMpIDB41q1j1rQn38G80Kjzl7
zNag4CbudX3MccGFiY8kgX1sWzTa+IBA5al28QPE7p303+7DLa5tFf1JlT8a9QSi
2sY2nO1nFeE35LXstGHAtOcG4ylUaq9kR9jfEVXrWQVdZbRp0WJE1GCNPXycVlrP
GJJhi1cZ4BtTYYqJiyN5W/FTmCpHOHEYetPHgGzIcV/o3hcgZxJgpUMmRqbWeNKk
fXeeU8lxwNNNrc7nc60Qu18CYq0rhefPBNRK9A3ulsSOq/d355cMv9GW28vjPX8b
ZTCquDhGzsWCoqd0Aeu6aFf2dYh/hT8aCgGF2AiVsaaYDrGaHURqwOZcqTpNjUxR
Y4tt9xcGv1zU79+LtbVZIQR/pcsS8zx7nEH6thvCO2GrmlCheLj1orx4L5sa+Zac
F1ZpM+ohWpeIZoGrLKp3hB+I5K2RMbEVQq30lZVdHdlnuqNeSyoWi/D0ojfrbrgU
EO93Po1nsDE2sgO8f0OEfFXwjTWmw8f4ywiVU0MpCPE+P93l/u5fTsJvC6GDgNHp
pr7cmJ8ni1yGi+I4WdYS+qQkgGc5PV1hlPbppDGRyGU9cb+IMVwDUdwtSdmFY4dA
4q663T8SCuOyWBg/96tDET0aqymaCXD1JmppCMWv6UX14gZTiZaLVgQ9aLzc3BHL
4mHdo+4CekaHMojfol5LzMsb57I+6A/H7kEY51FW/Ey5eU9BarVBzUMATXp/w+ui
qC+upYKAwcywsfBGrdCVXsyaSfTbKRJJV1QsP+dcDOixNd3jEAjer7zq69U6O4tV
um1cq2qOO22cmvMyKvrc43OGWOiTlJn95SekmRpDzlxwVh8lFSpTLcc9jmsqYvPM
UTMxc1YtAVa8TJRMA2995xpUcTWgd0be4Qyzl7SeeJVuq4XVMJkN4+GsSRyPR+Ne
pCezdqcbICU5PiFVm0nUGJLp/Ia64MTgIJ4FxMfCEPqWJA4bAYO1HKTuvktLbMNp
bzzmIVLogBIXq3+5j0LBDDjMVJty7U76iGZuX1aiHPx66kU0h/ukfqKg/DUmHtpn
3S6vSff2Bmh/OLLPPwqZKGZ/2DC4tx0/HP1RLYjeTAilaHe9sZ3vJGTI68macEdp
hTOsyFHdkGLani3gsjpLcuaLoIe0e8FhHi57Kruc4KIOgZyfGz2ArYnuca7pGKhI
h5qL/1gdHOrTPZ0CtoUeS7nHfWQu5QFLWPKkVUpIR9HlV3irjzjRr8g1WKo9v+7o
9a9x1tcBoNF9E0SAOjsIWjjRUqMJ3hbCjaNgK8UC8H2fdIW7+tn2g9spbd+78F7h
6mY15Nf1rUnGs+waviLum/ArrijyuJxq5t4wRzH9EzczUUGQrIhtooZ7T+itf/OQ
L8r7iCmOtneICdmFaOwhAEMcCYd23j0vLQ2EcRhi37FYglI8/59JrbLntXdQE99F
g0Ing6OzpCP6PgOohmQ7A2RRuK6/oVfN6e1sh9iHcOMagqzsWsxfFcPhED7B2mDB
qrGqj0FtHi3VpUPFzO2fVoN+YC7mWp7BPmEvJl1fXbB9HSAozlBLm4q85SZniOXf
mnRJjkygUWlMyfK3zcbb0v13+FhrstVG1NlDBJOz+YyzvW7ulm4rKYCj485Aqoi5
u7BlbzivyheIT1YTeAlOehgt6HoNobN8h7hdIFZa2VCp61e+UUAZKIVHoXkazVwc
ceqOLYC60m93IAJRhBk9UkT75YioGWmNyL8uehtw1uVI7XjvUlWa/Z5x5XNepNnB
JDNHMKBFtYICGdzU74bYQdmINHnRBMp3WjOFhGN32jHz4gCctB6PndfIx8mPv1kW
0zvCfecIFvF9S+kKhcmUDRRaeVJaX7EsDtfJ8zUl3Q62KHyQAOFyKlFdzlIY+EjY
0bvAUK5iTmeyz5r7CyxTVlJFsy6EY2OfGvH+eRy8/QpUFevd26Kj7TQ7PyYo6fzf
KylJA5opVURxJMXEWLmTQiaJDnHNrM5Okx+tBNwUd3c4HXj64A9DeJZUJzeSFGxy
A1I9J9vXKJ05Kb/sxO3sppcyG18kQWgy7UweG3rRBhMHUAr75IblT6dHkb2WvbYX
oVBP9pnZzvG050oXdhf+TpziPLAEvUFzOCKvPaRvfiDgARoD/mmU6cHKXYSyWduB
s1eyMQTqN6tOZ/16bXBc2RAh24jT/jq7tI7UvBu85U7+6BG8P5N+hFjtQu18bpHp
IuNpd7HqvNX9PJNQKcPG4WJEJkPTBE42g0otygudC3AsQxge9zw1wE8atIwM3EpP
TAbpes15bra82ur6DDdOjyWT7N+YYCexIVDKVeLCKchdkl2+o/OjXfFA1eQktVFL
ucZpfPltUos9X4fRStfRgB4GqTRlCfbzxEZ/Sij5vcQjWofdC/YvAtpqTdh4ARQb
zNF6UKoSvgcL0RsOMxc4uG6BBn1hGcSfPFrR/nX9o1uNyyd/nLsuq5V1NhnFT1mt
2PnTXk7o4OI+Ns6aUPjCPyBhujmQT1paOAiqDFXVgjQMlqPr26k00yDIMV1FYJoM
z+C8oroUP6bF/g6t9uNGL+P8hXhTjXez/aqIAyTy1vNG1XvtCscYWtaqDOy5G6Lp
oV8TIsjSoxnCIOMbCit+c6w8GEKS8oJXZHYUdMRztf15NezorYSpYJTV+z1/RKPm
GO+VgKAcTPw91OLwmZfxEAGnS11CtNC6BOeVOeNruLFBEfpyc34oYohPYerDjR3d
axJh7foNy4V0WpRUDmo5/y7pUYioyZrSH9GDefnh+DhafVmet3hW3Me+SKKDWKcV
Wje56quB3XyASLtb7sGCg4rYH+Of5+LwjknvynZwZO+FKJHZtkGn57lSf520DQ8t
67IVgxvc8aEN+zTQg43G+fzAWI51L8804omP9Q7FePMH0bNPQG1sMNtjd9IbbfGV
ujpMLjXVwq7qGdjsnmrB46LGtF/u1TmXraw92rL6SIHLMN7Q3cJ8iXYTb8K7Drfz
xW/vonV4asHA9MDCxvKXhcxQt6jUVOdisK7WfP8ScnwjFBV8ATtGRohErpLohdw4
jPQ8EcxgNofKstmaqAK4pMfqAAj1/Lj79E1vGJZgwbQ0OIbKd7WvTQrb7RWVOJk+
XNo147rVEJZhHUDkrcbUoJ/IMhoHl8KJVZdXhbneSkYAYykQTaE1j5RpuTa85C3S
oItQNcjnfbyRrbiLbrQPpiLOKX54lMOzKx87sYuOOgxmCd6QBv67tFxonF+y364h
sHzoqvgRaaxCvE16GLdalnUlkfrEWdu/75AV4ZxpgRwA2qOxjQEmkNckUdpmfhhE
Uc7nhaaivMVmB6M+uGUSPgV9SbmPNS8TMwcx0W3NoSvJaB8cbTZhddHo/uOM+2O0
xp+WdQ4aWg6kjzkz4Ojz/u4ezkPQKt5lUfoZTZq9O96ogX3N7uQkcpgioW6WGD1O
PYInvRgnpalayllK4XmMiB0m02xSrn3pIcpnc1CDKAjJT+j8nuMZI+9nfFivVjc9
Gst5g0ZQAlnkqdfMMwH8ifQ4QNJEYb6Jmrkq1Sz99JDwkZDBqterPhvpnKfXm9Ca
AhgTI5uae8/hM2JrmPW+Dry3bxoKdLjKsRkbvghL7HH+AHb9LlOvv11A821WxJq1
/iJXPIhJRgky7jBr5ZtSBang3DHFQjvVx9Ty08NA+LFUnmoPjuju0ty4vipEGKq6
scHBFdjNDMxji2BdtzFaS6ZDRMktakZF5efavxYnfWOHy7V26/+7RhgXBxaFXlmD
1GRjwWh6EqYQU01115opHcJEYbROhiJLN0UGcPvnJZf0xM8fUE5ogZrRVggNliOa
Zv97PHS+0WFeOBamAvjfK7jwMRcGnImRJWyoqBFRhrQTO2tcCl4zX6iLiOnM7CDa
Yy/YW2NQuG+OrkbTSrONCXcWACrTG4S2BG7WrIhArlGmPVxAO+MZ/q59T4fGfg7F
MsdowIG0FIbk2W6VSufMPbBSPVoHUIO5BujBHz4jqUixMQnpnuV9DJCBTqr+vi2w
n71CaXuxCkp0SbirxiWy7sakCB5tBO0dRWRvEhsiS/w2bD66DzjpS+Dg1clOuw8O
SBWTW+UeaW36ahZoQO3STgxZBgRCOFpIWgVB7UwGbffzh6lLBQnG4hJZtlf3IN2J
VR+jd4ehQkTgnAHAODtYbiy1sSCJUNRWb9gt9I7qm/YuMah2viwrx97Vd02gs5uQ
SXxgtJ8o211fgMiKSFDfWL2HbvC7UPLf/X/TS02FBOOQg1ax5LZbPpNdODz05wSv
h23BHVFCrJ+AE2IssrQP2p5ScPlMahXlbYTjR7o+S8y1tE7IL2N3oC0AUBkEV7FQ
42c/jv+HqSzDQRedW4vwwDJ7mztMhRaDmKEa/3BJuJJWgQVI+Jn9UD6MYaI3INsP
/F2PVf/X+5ImjEHBxof3j3WwlFNJvRycM5IB48Y2cVC7ZqIBysN5d4f4iEEUorLk
EdWlrK8IIz3pUnqkbjHn9oJUiX9BgbFqVXmDd9Ivp5hKDIKHJt8NKFKt6Zps/rYg
9q49aqG/uxLcYoo62Z0asRbj2WFFElOFhO+8YO+V/EdtRdj0GGsVgz9gNECxPsj7
zjIw2N05hAUUgB5qybl+2ZDSTIRLtliy/MT1F6tO+FaUS03zMTY5nr7Qv5wPM8+x
7wgY9batl5RewUlPzeh/eiMBp3TBvqH9VvlUYW9oqaiY0zp/t21wdim2AKBiVFqi
oRox+VKiXLqP5q2K44h3vhaCm1Qq2XsbXq9qGOwR3L5L/9yRx2XOWIWDTlptqC/q
23GE/cA8d91J/D6PJcKD07CEzAm3HzpQXXqc4N3Pgr22nEUcBWvEW5S/3hWONZHQ
yMJcLUGqKfemxUiZtJlbugbvX4Lv63rBjDXNBeJHlQ5+mmC8PWJjbqwYeRsTlVpf
5BCXTY/NN75IQLrGw3i18iVEIMVLr2QFnuRb+ua0I5ZMQ00qE/9sMnQj9nJGb6DS
nSM1pkY+9a7N7N7ZWSFceqBU4R8NY5C1BblXX0Hb3Je91rnutil6WRoEKiMzFVu+
F36Z1+DTLGItxn2mPbuxDKrz1AREYB3FpRaPeQx2nwg2fjUI7cSCYfNkIb6B7+PF
1Obh/TLtFoGXXBSZ8zoSkip/z5mGjVIy7IhP08xGYFOVDTayD98u++PWEqJN2Jg4
0LMkCBlObvdkNwfQIXJa21H75GqNSFpGMgcPzB7fqCD7C61u04E8YtiELazAzCJK
JmHen7iWvOGnYBdQmf02sXfi1dc9W+4r6D//A62yeXFxNPC4SnXfQnanoQojBPPk
Xb5XUpahu2CbkXklErNjUZHeusGaIsqK7kg1H7n9QFLv5XIzuUjF6USl8UJQuRc9
IN0pHviydgwELbP/oqAW2fOfLu1dLBWWExV5QEIio3+bnRnkHm+7q8n4i8WO7QXt
mgeiUbHzoSCHtCjrliB6jo5fGdkhq4tdMPOu5SVLFCvzhizOzxvSxomAqUE4cIRk
8IE506sCiRO1995pov1e2Rn5nMqvJHfasciXs+TQYu6Avd2kbL4irjeie9QUt0uS
ba9yQF+dPjz9gf77qCYo/8TaOwnJ0RPmBXVXVANhxqMvXNW1NyKSaetZTM3q5q8s
BjtgdMc1aiZ4mLArxb+R4/0zaGD+vAh7tcOUVd5gxchncBzZ76/jwVvvBJ1U1Otf
rBHVnQOeRzMASzoeuokvtmnBG/w9Km3MwmogXWiX68nqAM+nFW88mgFMX5ukDdBV
wZ/mDe3sFemxqzaG3LWDvS+Z01aVJiaHK0KVf5NssQA3K7xrp6lJsTyNsSgrQ1bp
4+TqOwWLOyPUcUQyEdar9yrXz3c1kvfZL4OECPOTByZL77eVEVUAhxV+HKpyXFhu
o04XwrYZJDManstIO0VYOiQeBEoZf65YP68CiChrK16y16HIYeyWqNKIcNxa9kiy
CpROcmmqT0s4q4Bbq5bmY66k0zRCwU9v/aBWmDKiPxctxwA1PY774PWmi36xCAJb
frXDfIFCjcFWW0mJ2Qo8KCpHr4FrAXRiV1If7huEQQZ9Q8tcV1uDahfr+yZDfyds
wCUeEtXgCo0XGWBuOL4bgEGd4/qX+yq4fAEQcy5YAxfGRd7jIve9vcohMkNzZftf
B+kY4Qdiy9SqUDHvG+AOn8pMYwdXyv46IFqmlQZI+n/+JkBKn8Jrlumyo/qmMoY9
daW63+T4LDXTL3yHATtHFbNcm7tfLneZ3kM9aLx8GVLAr8dTvqbYCoEYn/FPusMw
jixWBtIdKCz3DlLMmon8cVCVNTBBJt964jmN4m52YNRRtwpDWABrHTSurf3lvX3P
ZRN8GZNNjSCXnRWrSObH+aL8jLp+Tn29O5Ofwa9TL/b/T6+yyYXgCYaQ3q6GSUcR
q5Odo47kOjW2ds47qOv03KrFiTMQQMggh651Zn7mO59DEyWs+w80igiqnuX+nozi
n2VRabBVwcPZl8nlVdrkOP8eXYUWAgfUckB/wVMXs/K0g//GtJoUxMRGQkl6Q5wl
9hXxGBoZ4+NcgrtPOWTwI2tCH8kLUOdCurb+04MHDCF4rS2YmX9C80p1BKyw85LE
ktoLNOJQJx4EeIMdvOg188QbLi4kqJi1vpRf/QtdQXZdXHn4XUFPVFb2SwZ/fW26
Us4CzNSFCVFyrV4ouDSbSC/sci5y3RQ+XaoP6U0ipjZ5BoEvr8H/xXGySdCvsycD
nRmJL8hQNSqKfaVF0tZD4x4Xl/CNe2Er/sgUHrr3ePh/O2JaYRjI+cYXrjuj3B+l
aQIeO3RSljuqCrTTWdWOWDnNN6dWNM/5yxSh2GBWrUu6PWUb6GM79pSRPFVmIRIv
zUl3M6cMYHyueYKOR44HeXYXJ6n+hep7Ox7Azl/PbsPEqY6ImvhnwgL0HksuvhDi
0rUXaqK6BlxHy35WlRyqudXGGV2KE8lZjRiLrRW8CI1zHcIr46o/X0BTZcUSFiFL
B28iEWP1Vo/fjFlTO4NrzJNbS+MuLpMKBMIW09lyhjq+32Ws95Nkl62a1ROZIkNE
9RmXGrUV4MIfUatUhkkEH4HwiTdQ0iS67GUELi1lVWokMW1MChVjPYuRSkdrEe+0
CIc9OQq8lK+zo1Zsaq7TKE7QmrytdnqFarFwFMZMYSA3T9JWAfajdtUFq9N7Pxwo
xFKDvc8K/SGSmPJQ5cfxjSCGRY0Kr9+4kzyi43cGkdeZjFQwQ1QAPSPMI7IdZ7U1
TjdUVO525L8xzb3dI8Q8J1tD6nUh2SrLghpULFIO6bzWypXRyyDvdXqAfXoOc33x
cRmNKr3EbO1gm+PwHynPquwXcTECTH/1KToN5WBnKz9zg0h9E8ErsJT9DspxUB0j
NJFnRxr3gUTkYQBpSQt0cLjeh97iTWzlPRyPVzlk17dBb2DmmDi4bJonYhvVyO4B
2eg7BtmWVsHVN+RQMqNGaEDRegq3/a8vFd+TJpJeq21pqaSf42ZFlibYSPJ2iqyf
wskGl5LmPoUHy0zqtTXHzXsfuFagZc88WGZO3hLIMx/zwzlrdEGXN2mcmBH0QBh7
gaWKRpWWTj4KBM/gY3VujxwA23dyKAG4D9b3l9NT4+JS20WNdoFe0JUF8CY99aR1
OVlvl3baciBbmKfrDqJ+0YVVNO1qjtMV2rCkYwwf9odjJEI1iKXE0uWhURN1Xiot
F+Y+tJrW+hNVkSa10wzEVDBKU8c+aqz3dpg2aG+uT6qN54DSgA4e4dqvvACdBt9e
AakLAwMo7JEx6fh/VYSAShMCe3jpLNkUwI2KWqjfSB6FrRuWndpmQcQp2bqc4rO0
JEBvxB4VgVAnO1bWhMfgujtmVSs0U+emo0XW/YhtdPspq27wrfMGWOb6UY08xaVX
jGuG5qRo+TvnoOSAgee/G4dBF7FaiH/YsIwWUMwEoidUaP/COHH1yqgmyOAcCpx+
qjG4jVzmvx/uoJdLWHjFq7hbEJJgdvcQI5f/1cymueKKs2CR+/+YGkhM0zMGOV+A
Hqstm6o4Rt8uJIelrgN/6ykUs7An3MGlOY3YYRdoGYVjveEXJFdCEPbRmicoHp3u
OkiPPn/YzkWIyd0C056ShYNxUZPKvkmVQ0rWbXNOdHg7IoN42qTnMZlcPJOD0hb5
8hED8Gf95qRy8jVNfZ+ZovcNAf2O5DUGsAn2WAcEQGpEFFKM9I1Xvmr//mJrggun
1hb9tcHC5rL2c4lnRtGFPHQPi3i6LGp03ghQ2WpMvmNaV5CW3eA4mYp1v3gLo7eu
KAYKpkFHK5eTzKr2FHSeZuWY3mrpXzFnc74yI58Te7oJq7IQgYyzRBGy45gTzjbE
Kl+UB32U5UimsUuqLuAC/50ViIsQ98Zc6WDv67U4BFH1EvOm2tvDIh6DgIWiNR2O
+L8uOmnx1hQRFLAmG5ICI3XYkusuBaLdsl2XCJf4QZn0eXa6m4GcTjYZe7YsKImU
gy1WnooIBt4qf4Al1dTq8q6b7H0EKCzHQbmqD4GsKDxtl9fplqAepwqT+yZCtRnD
aCPc++ABGgGSiiMsZVSkKHCUhAkPMtYBLAT7PjgAyO69/jkju4IYXnnWiae6IdgR
cqwulgqI2HWpIexyV4GqW0+aUAMW0OW590bX56ny5LADMIRoKMqY1u5mSiTQsQYm
x+nn5LpeA8zxQWB7OsqcdUeSb2r+aq0K90eY0adKCNxII2ehj1e9VG20VW+31vGQ
KEsbiF7KfshpLhyx/Dxb5uMVwYymRK+BNxcXwMFbEO64XLicoYabGFFpEtGwPYqL
NYjsP9C6kKXEDULoaRPG6bjCwUw33hFVOyUDQQs0NolrCmB6uoLwLEI+jQpYpTzo
FqwRCMrIVYwXMMN4MAD2UdoMeFjAwClCg5GgWTTGjNbTQiWJleRGU1uctgLCUKv5
ziSkpD/5vlbx6s8M0/QC9tcWLq+FvJQZPwgh4OmNTdxLyQZ+HTMS0d3b+H4M+pdo
R/jM2Yc3KwQCbyHHLzueF4TCYJZZOjO+f/pMFuTCqosQs9tmL81pFYP9oHMQGVBQ
ZSsO9n2Aj10RZ8EQmrosyFBhyV2X+LUWLiKZV5sOZdsFC4D1YliIXb52rn1Jhw0Y
mqw9vsfBaXAvctJvowVxJcPPcTx0CFrErkRgBuwmh+DRG+hMgBhMrbwyPpEZfHWs
QgF3ioXsCuTqGfjbkeaDO73/H2GbrRr8k4RkKFWhKqYVe+Ine/9wHPsbWPfk2EQm
COdtQ+IY+Ha66SL1z3aDhvhtNJTgGszK9ZIMmhC9Bb4n0Y/zBFbJNKkwMIEJ06St
NvuyAC2PCBzxxrx8kOleVauI6dgxHxCO2SsSfvg+olu5+N8XppPy2luANW1e8faU
ymM5J7D+tZ+w56u2uxoyBu13ayjIvgORrwguBVl91EzLKCYHLlVXtuG5uy0AlO4a
DZ2DlnyPYcXadsV7XcmyBQtb026VrXSuVoMS3Kl0taEYUNUNV8Ou05dqdKCSJCzE
lB0f2JtTDJktlFinMaAZEhPXtXZl2st4NzS5fIwBTctvI89ZOXlhBvOT5qaJPxlW
ZypXNpeAy6iBPtCnjF+QYApVC6gWBSfeXq7JXXuq1BZxTMV1RGzZ0RzqoQlZymYb
lnpvxX3HkIOmi18qBBXIwCZ4bdW/QKl3DzKq9Uhs/p/emXez9Cz8v/XiI+E+PxF/
XEbrcz8W/mq0Sr2eg2iO/Jp6rakwUdG3WHJ+nAmx/SzcnvrhrYkbIhqBGDVmu2aV
hut8mRl6SUaqBnZwsOhwml+1yebAIApkQofYNBVtYcSrUCTSXqAkpQQwvqVuSKst
DZ4pGPxryBtYZiXHlffPpdAAaWvb28K7TFRvr10NnnlvxEHjn1sMZMNz9oUSJ7iz
2SqlMr8l48YirSnA4OukvrIlwF+rHWy5t4gRm1MrQv1IUL9oZaMXvjLpWyMoHuAn
pzXJqdbxUuJALf7GYhzdREdc4ZpIAwsFjJGm2TAaQGnZFuKNC6gQGXttUQKQ4KJ1
B0imgIf9KtJjwQbhTGO3mQlQL9pyU01SdLvOJToN+Zm22w9EgsuSNgJouMKXA3ZZ
6rOPgPkQcOGedBMf6tSWSSzXjnijXtD74XzMpVqe5x7vEXzoHxeVZ7edlxRZ2YFl
FPvq6FTgNUFxNyIuWkLWTZigACojnUmEANSjwqMcfrTnwepg51l8JQG5S4UWph1Y
sQ72GkGO/1m2coyaV0+R9PV81W9wFcd26P+TDcD/st98QEmhFDKHMMDrrmQ9BgHm
BC1EpqMP08Bd7MfM+gjGL9IUo8PzW2DdXHFeAEKZ0BR38q47Ep9BzpMe/tYw5uQR
gjscFG4cMuYzUn5Tbu3s25Xr/jt1XOd9qznPyaO44IV/KWqSW9Vwel2hDznzsZSt
WhAQcBHiYu1pjWpHqfNmvnZb52V9O0c3jxSwpkgTP2zxfN0pydlPuOleh1KQMFVf
HJAPgk165CTWvuUSYvWqute3JXmOHvHkQ8ueIMdKgKykbDUJQ5yi5du+KeSD0ihV
etDzKkVLJiK++rVANPMqPA36k+H/Uz9mElYDxlLMi7hk3H1qH/iNYs7VTsnReCMQ
ckcjRFHtJbUHRwA84Sk6/GR38OWG0MiBZ7gmuj1zYs5dfo6C3TzBuoSZjQpnfT0V
L+CwPgaqYTd2N8Ybqi2Gq0MT49kw6PUxfHYNPvKT0se0QLjrbeDV3ur461JRUsI/
attxMVs4eLc3/54JZHqKSRF12IyrWdxuU1aVAnNMkAJx4IOKpLGSBFWhttQtFJ15
1K97J3MC9aR9cm7nFivTBnD4tAyr7gaQNgIRDjTEMnCtQElDw6W1qSyYJqQc6Ie3
Y5c6dpSc0oSMv6KufRhLfMSwUKenKHggiQlmxDF6gYqsd7EJ0XCkI4MldGXGiPA/
A2SW7UNZsSzHjycMcNjt1nHLJnM6VvuLvXQY495pHqFFqWEvQUxXQhtBqw0oCVfT
DGYVFMHE8vfPD5GqHszXvhwaZi25GkyA6BTCMJKSWEhHoCXk+TIoOjWtvID56ksU
lmJaxWDRv8GQ1fy55mHtdlMnUCB6liPEQaKSHn8lkQ0w36sXdbASvRqcCi5GZ3BA
NT7KvtfqHim824/B1ypth9kI2FsxpidspqQpcwgW+jtsInyzTa8khSfquB2R1JOT
BXaEfC83FoNK5sPnTx0J/vP1YLWTfHjeE/krvSleNv3SzfFxcIc4zdO08i5zUBEh
Jp9HAYQBQRKvbBS0NhqIbEatRu1z2XFwvyqYfbAdqw7ZgrmMpZRKK+8dbILVYdPf
Btb29YLsXqEblHm/tG1MwokYzgfB2MNJ4kSRDxYmpRp+DXPaj7kOBX+J5U6aYw4l
x44BHB0oUWjPmWEtK5HN73vQwBcdD7xmaHLpTW/sXU3jjtcqw2SkMVeolyZR5Ke+
seTkSrLqcJkOApCO1pZl7oIdVUsneZpsalZ7NmR8G9sqfD0uxa8bELJHbapJ/YnP
4jS/no7N89cDWwVUPd4Lnet/tPmjBoeQwmvl3OediayC/nYr0WAwULsT5v8Etyc3
pMHHkceTwXG2PNl0tsUHUJzrcAFTuvAI5cTdX6Q0dC/rVEdw3r1y9a25BunYnYT/
cQgWgZOKum5PKyDfYcVds7oycitzjJRZrBsqNMVniXf2Mg3xlOkmumff/+sWytKC
mOuI2Ebp1P2/xNQu92gslVaFGSQKCiWt69HiWF5QBQxkAICksSdV/sRPsQrCg512
ysq23ZoX8RoeCMQ6+gf3tudQ6JFk2JxPsXL+V9FDbTcdoRRNig5OtfEyc30bsXMw
M0yR2SEIwDJlHOvG0TTBAVic2N4xaTxJWTF0OdfRmCeH0IzeYSoEuzXcAL6JkTnj
4+siHxjZmRsWrYmEuOnHw59kFaO7IqeRvNvEgbP6Y7/qm1GBEF/JCowYANccZ0Lc
3RXjA0OjtjdvwvNI1bq2zO9+fJ1pzYtA22w9Zskz8ULkgyuTuIUuRhlaf0FuLbG7
3yqZDK0Wlz9UdDd81vuKHp0u6zH6+PByC7wf4TitEPpSjNr4woC0Dqaszuj2xYsC
zfzvoN5qbX08gHI//qyEfKwezjk4xKEnQSdFTCxFiUoAPlOHzOh3XgSEZHFrT1Br
2WANGaSGxDeEnwiTwCB/j9PKC+4ohKP6UNW4BOWWQYSdBPr0xVRm4R4Mz0IC07Bm
UBxWoqZ+UYx5h19XLBysP90R3bfGAjq0vmerjFGyxCLwdz8po+gBIiWBzyGPCnAy
KRE7bmi7y3gfRQ92/tCgVIVRUe1PW/z4W5+zx29LTYV/DirsV9xljDXZlX7IqbgD
k8azSspCkrlZnAx3gavHrO2JYW14ry3We2eu7kn+h3LFb3JKT0BDPxozdVQ5o+VD
ItpHd8RaNPikSbb9mKt9oVEk4T4fiaX2IHbUc6dKT9Pbn1xgrWlrD4oSmrlpGB5r
GL/QziSV88GDhDM3vWcSmXiCxz3ywFZ9VyGTjNtD6a4M38ksO50uJ36F5z0GQk4a
UXkLLHkS+AFLlRts5dNtY8X3T15eTK9lSr41FjVf0DO9t3dO4EZdCrdpyvPCIK7W
cCETl2AZ7I6qnGu7UpMh/Cbr7h5ljFp3djtYX5EsBhz/l+ywiszEvDE75KMcPKdd
17g5S2KUjBBaThns0287jDVQvzyogidi4Ys/GsFp9+5yjGyvaCJvKG4o8crrZ/rf
oqdGR5Qws5If2w1ZWEPGWP/I+1UAWi4gH+bc0lLPnuTgS3cGsgmBC9+aSBuMs2fr
ZbgFytRtM2NDhqaJ7W53IeUeTL9GvdhtncUS8HHHml3t5jjUmKAzpsj4KVJ9plOK
i8UkBvVw7SQMEFg2TskbxeHJOJe8eN3jXNxtz49LHKzJ4TTB3lx+ARHdrOvUiwrV
7NfZxY21zAtERc9kY5bG4xhyudwxCFjzoDLLWFkl91hRGC6abQBTSWSpJwC3Crd2
rCa7qHvT7ysPTTxlGPo0ZrhFRGzux2nwEr6O3224gAEx4YgTX2M617fUCkdVp1xl
J+AoyBsxC39pBwHywNu7cbGxKWqEBXcygPAhpMjt6taIMW3AUrWdZPicJ+aEzz5V
14YR+NuWvnUPUN1MERw6HIunTBoW1l4/s7GoRbfhVBXV7mcetyNz/3if++d8hA03
VBQRpYckLFtgszGjFlUWxkDGvFAgRTKd7KCEI3kTzkYvseqlqE0ckp4z3AdjBJjQ
Eiax7flwYY0B30NkDX8VuHQDv2dZ+/VE5ATDe1Cevr8EQQBcyp3nH5RuI9uEbxnk
FHlcGvjP06FmeNJ1LnMEFN410YcsPCZcwATG25F9xr1h3MeX0ypaTHrfm9gOEqUA
REzu0zrSvuDRSDjAgCOR6XJ4N9uqDx4rgzubBGQPO+W6H0iCo2OcbqTDGW75cs9p
lDDunv5nB2ThgLW+Z9DQHbXDRhamO+hNrksaTw0wB+LbFLiOEg4l57JAQO+0JY9y
W1XduBZJ/Mf4MAE10xIcVxAAr2pOxI4tmLRQU8l0SZ0sk1eOTZ6tctKRcqiMjLEN
kUXxsNHRMhP9R2ZuOCI4dH69eebcL4wKpL64p1efdrvBLlT5Yd5eLNi+3AxLt/On
CQ9pUnJpCL9vvYXQbamQxemQA/VYx0gNZnMNOTpYPwVECVDOAE1ouJmcMURidoM4
i6yaOfhmQ7Sfyni+S+Vy5BWkjXcl4jLZDre2ljCzWCiUCyQa+NdMrMyMkeGU0zuJ
0eIikBrByh2cg1PqYYsWO15aSjQ2i+hWM//J6yjmkUCpOjEdcTurBSt/Nua4aACJ
wv5FB0vomrSOVeYf+mz40LQpl6qddaJKQ7DjekU4/0kdx4r8qDr7ucmUgUyOTDOB
oP45ZDMHFOfYq3R+EeKWw+UMBGxDLCHLnJ6gWTGu29M2ksxvb3abh0vIjPCOL8ll
Vbasqu63gYfJKIVy+JOmSCaE+Yge6VaNy9WFXrEAuhgCrDiquSiDcTz08V3chPsU
ah/IeZiGhz/5nUde8usm+Fx3TgknkR6rvlaI/1gFPoBjzJ5ykbuEfn7dMtcXgwGd
WBO2rEJaC0ucLbDNtMby7gm2kpn4nLZM1V3iwx04SIQbJKt9yNLaxJCi5aGDmcxd
06/UHYkiSc+rQ5cg6xu0CX5WFYlLEDUMYKgC9GpKDtejFk2lp0d1QHVhzvjGekbQ
mzeclzM4P+DNFEEVhoqyUSmVPkl5c4fkOsE7XhVCTjhIF7lzymk0dgz9fvxQyC5X
s6HYRwtm6E07RtpokVTlmVOcuX7dMYp1kiTqDuVKoanuEdBQxZy61FQu5x+RZ7UD
LFUU9b+XtWMgEp5zto1WAO4+Y0yIJsf9ECuQcDXcRAfSnHZFQkm8uUmy2ykpJGWL
yRk2VxEZh+6U0javECfKGROc1dAuiBeFTrp0jN8UXQIR5wAyIHCk6L/xL93+7XFU
BsRFTU+elPX02JAlHPOf8g/j5C8KaoXQklGjg+XgfBJlNzxru5RADO/LCOrTgNjh
BwfQyGMNRnLc7mFKtk/S7i2VeA4RmHffsdCTmoxHVmrhYo6RvI9/dT/Lp4XHu+AX
nvYSlsq3oZ1YaapAAsl3qb9QxA5J07xomPEVhgI6oikGzs/LTF6EgN8aMMx/Ryhx
hvpZoi7ai2eGKnY7fCMfTawr9ULGJxAX9qz/G0OLc6HYIqG/qdRbPuVsoePUIGHD
M6mJv75hoRPavg0frhjlExeAw1cjJ/FGf2UdzXDYGFp73oEBNSf6Q/PASeBfASDx
Gc8TWZkCEWXbS0bUt6iMTnB12x9puS45MD/qGzL0f6eqX7ehxmAEEIqexN3E++kM
UaBIHlUQJhDFdNNp8USIzfFQ+9cnY1Z03TZ58WD1Ee98rcMG29MPCr5A5za1/pIH
AX7m5+0mMV3hdyskP51I5yf864K5AkT7kvwrBhKOvC6jvLFrew9b0TtTnl4bLyJh
zh+6gw7pJQTCf3jdsXUpkg5S4w3krJPSFASrkTMIscZnyjzuyDVJnqnTI53BCuQj
Ntvh9zQGeF1bzQ1isaG6BMJu9OYwU+vpALA9/sU4SQyNODpKhgpMXO5qxvhm/XmA
yTSOcYjCb/PRB1zn1sjKPOr+tXBx8k2r7/rYtss2eiCV49LObb7gNZu4FULyKpfP
sSuXWt74eVsjto/uCEPHlMAyrVFyVN8ymCs3xmWuLNViyyDqSbYL1kNCgEv2AfSo
f1XLzjj/B33TozzUbXi2GWVE9XRpbjcGlTZ1v259r2uV+nK7j1bFB2NOLPz2lxBd
iRpqQwQ0Jryh8E0qvUgfTH64UkM9XFNRdWohsDCaa3kIA9OT94qUVBCSlzzEnl6G
HOoJe4DCHWVDjmIaIGrkx2UGntXCZ3yIqOSIgupe9uQf9qDm8uG52s3dg/4iGQLR
KVDs2ui2YABWicxfROEoWQPKq+ooDHxHJxvHwvpqxYoL6PcdBZMzIJhf39WMVPXd
/qn9LMM/s6/jqloZ/zXWWzUbV2FHiU1oEFJmMlB2tyukdevTo2QVIZTNHmzjLxH7
XijjgzsgslnaRHkhMaXCqVBy6qOX5ymTl4EnvO6yITGk1PH5+LrljkS0Cyga2/ZQ
CNYX4E+nRHrBAD8YreVreGbLQSslMk61Jto7XOe+fDu6/EBspLoeHLpk0y05jqJq
umlMvG1YXY22EWFDWntCAsN5E9lLOD6do1HOmDejRx1EFTyswGmr0y5dJyNhiL5q
KB2HVH4VmLXVDdumEcczyYUs/sW9cWeOHwy8VXOTK3cjjIvjM0pTEHhzCYJX6jlt
6wADaxkMROXj8Bfyt21hsxIhwAiaMCSN4nTjVAD4zsYxt1SK/qgdbjSGcTfAFfbo
IjdNOkczg/cMX7qjGSIdQDsAgMTME0T7sxPJo4xbQIpswfnxMs1V0HtKm33IpGOB
C29rO/T4yHjqyPd/g/ynMrhIaOCuMZiJUt88PTyfx9n6SCt+Y29L1zaDEEhZ9BEb
ZYijGya1rOBM+fQXowwdbVwEa7ubO1JwSVByHlVDrbv5JLr7Ltjc2i5a+Z9wpdwc
p2EWNjONK6IPlLgZsn/sgFbYboRGKMttkowUpNCpGDULTeiPN+w7+DkEL3jqEaWW
yleRWzcmpivxl4pbTvsoHYvQQHOeQTnMI/LetOHahxOqrZzxWbbJ7oG1H+BaLL8C
vyiRiVp7yEyDXYDwMDBU2ptJ2gEAJPdLhlpgwXd8p7WQK+vhmC/ZQ7LUqYwfMul8
jHnGdYu2fYuBkl7lxGPtLgy1mwg5DSLCADJd5kBDiVHqY/blPnXHhATLPSeDM1ch
9/N4cIvAJAnsRX+eWqTeysPn21R3NSomvrEBJ1JCixje24AFvdwLa3hhOLC+MQci
1aLMDDEFjpTAGva45vI20kBiQNKFvpC8oV9alRPrMF2Z0Gq5BNJgW3g3Sfh8jJE0
RHNlUQqrTbWKgBvY8XRkp/4LKqVdg4fWZttgDCEyn0oYpX1MPAOi72vW7KDLoqng
eSADApfeHiXTyDHL6Yv1LR0Uimg73K+X3R2Y0vIQXMsE6CZxCRyNk3W7VXhYCu94
Gv/9OXDr1btnU766Y9UlUBHqrGp4LCP39SlLlHAiF4bNvKm/sdUs1OyhOQDqcuwm
QVlubQn/KPZ12Dhaqj/01qLzCFi+cS5zcxWRAfNuWB52tJjlw/koyXKmiNmDLwyw
FxcXRk+zJNpG4vXC9Pq/2NzFD5AAjrVbsAM36nKbBmQUgnjXR6Z191dsC5zrA+7w
M4f3GDeBR9TeQW1/pXRIb3ZTvjjaSPUY29dBmrAkqHFu9q67qocEmf79aVKwrE8x
/TOh3GNy063FzdAoWrpvuLm0pe22yXwDerdKWH8Lk/vnBI4oDoVHdZo15Fqvl7Up
symriM7wZwDPcpGPUPgzausiGCuL6HEmm7FY6xu3DXqcjagw+ESCcC8QnPbcFFOE
kjHL7Rzb+1qAeyzCMKt7tj+4RoPXQxqq8bkeVQkn4V6yNiHdWGs07IXY2cJOLePM
Oe1t0BJM1lSicGrRuJM6VwhzXS5TT3OHtFZJsp8g4Bg3bjbIZ1esOPLhk+hKrADh
zddGkssZb+t2Q6nIKET+A1LHDXOaVcru8UUIIAfzvJVvT3QcwAPmGPG3uCAUTYbM
/37IiFo/sF+liZyi92q8ZMQUG2nYc09kCPALQqAowdGCpB/BB7qVoPUzWVrt77vN
t9t+eH0R2lXoJiiPAyMjqQMJ2CT50X34vk+Ehz1V6AnHsM2pN0FkUvFCcdKklU2N
zF3D0UHsyZs9TeLMjOIwoU9PVprEAn3hUyaVYnpKGzsMA1aRjhbMsedNm08timsF
PX8NzOer4v4usjO5dLsABI6J3xOZ0Aouu9KWhHbZQdhRIoBCELcRYxfDWI/X36Ly
QfdJ6GWCoLPkx1IEydwer0l8MS1kNfhZpFit73MAw6maP4Moy8yqk/vz0mCuq7VJ
0SLbUYjHV1tG3VQJOpqdcIqL8ZKv+4cT/nSFEXEQKg/K+SGtVHIKte+wt/xDxAHg
XgThFJnzbNSnF3LyhKYVrRwQ7Zs98SzPVqxG9Gfrzkf0WH8u6bGrmldeLIKAS8wY
yQOTSVt/ocB5FXIPwxZ9DLt/eYtAHjEuxC5EWtos9npMwLRdraIyL7xxDc2XS6Mo
+h6q46Ado4suzgerfCvQP7UXqzIxHmka5T9c0GZ5RdHG7f67iYKjU2XVzKMnRgQ6
QIRkggwj7B56qmAsP+cZArVuCdbyxABF+JgOSeN9PAZ4G484bAS2xAUN6863Xmxe
UpSRqsAM7mbnViumDHmtooCvss5iN0k8mZEtFihNOPaLXQWY4L13Psf7EIJT/ZvM
zBaAwXasyeUXZDzbVDLV7c/ti3v7Ff5gXB/e+g/pIjoitBCdaKyMC8EVlO/svRun
AiGI+EN8HYgySxtnmf144a31wSsuJLKdq/vrAXAQZtoAhXhdM3SVfsLlcdM00nf9
w2KnMtSWph8RBnnitSMe/qemTHtgyOrSvRzI3/rKTDw/REvYdDUTQbVakMqt/hkB
ra9Rx0N2dKx9gssI/SufeGsN4s8EOfz8PHWiQRRJj2U3oCMOGqf3wiHjO8PQoIVY
QYp+wzgLedqeWgNJPI4h6OggdfH51YQ4XNRg9e1OZJIp+DRyOXKS3TINOd/w7fm7
B/Dry3oolvqtiZuUwU+HLBESYNojWHGPDB6dHaytjSiqPMXZmADISZcCNY5K1QSJ
v34Xyyu0hcsNGNfyV47871cPMDbID29rRZEftb4Et/FTckoyseGLMVcvrEHz8Jqs
1geBEcI8EJlNxCG6FQGBKMps6wb/ZgdC0PmhPwcDRSAFd2az9XQ9S9MqXvenhJy1
t2DUIc2ZxGdFoIsDsBQZdPkPSuYiudiPLimU6IJP56LlWOM9thlrBLnT3ZZZIkuF
ztkmCD8jZIVQ34OA22f4Vg6U8Az2yzvMuTd+StWqfP7BMOObak64lZA7n5//iO3Q
nCEKGpQRhRipu8YHovibMoP0hwluEzmTMa+iQRB0HYSlkqEO1+ldLL//sf7VA8e+
cch7fUEVWMEkh56/C7hHrbqblOTN4UNUxRcSMp7f2YKz7FtBG5YOBJZUK86VpI7k
YSFU1TWdaXgq1bUmBBFRrdsJF0kF9ijAq5XKnxnc268cRHW1NUGXNcLqljEg7vmC
xNrofM8650Zi3Dxy1fftE37auHB+ojeN11GJdL0TUK1cKLxGxJVbSVQxjtBX1i2u
sJvWniN49Av3bqDlqzm95PN2mpQjbG/3C5hyA9oXCNwug06HUoPI4yGykLgpvBj+
wRpnLqaOOtRjvC4kbRCkjWRW64nYEGOQejsHfR3FuxZc9VweXXICkoWCmMyS6+zJ
j/Y4YaL75cscEmUxptvUKqoZlNZFQWDmQYLg6WsHEeJSMK+G0BK94KMLplTTdEO2
pwAGPitPAPO5EDa8wUe9K4MkoO+Q0acO28BYgGWQyLbakmYdTDZgRxoUMjOb3ifT
dEnqAP48Vszt7FuBVRjYW7IvdiO0axKAAwgjISW13JOWG3/x4wTwR0R88V1k0nRd
SBFoKlIHIg7qHu9Ji1AymhFm638V3edPqX/MbIy+s52QSnTb3CUVnYFCGilt3glI
RsR9Kx35XJ6t67KdjYwox4dJd4ROrb6mCok1xbFtge44l81RysdKbcGeQRgCQdL8
BWu27VYu5XTAWALgZsT7PoaNl7vo5TEpJBMhgBZ1lXDg1iNQ8d19UQSu+ct0aK3a
FvRA8nHrJSNViKAZhamnPk8RGZGBpUIdCEswPNXpcDSCo/LWjh4eqRf3kQfdsxXR
125M0eiXaH2j4TYIJX8u2AD34ts996X9WsuPd1wCZv+3rkzdd6BNhQVpKVOibcmp
8wVyEAnjoH+YbN8ciqK0tQZyEsFjCI5MjeEgbXSgvEB9+2F5IyZdPZkh5wgixEaW
z+hvUMOMQ3mrGdlPJEP/HG4ANRtThF5OZZvr4/TzBQBZ6VjTA7mgu6yzj237RGwt
QjCw331dJHpQuJSRKDwuhxjjnyjQHNpQIxok9uHkhl+Q1Duumr0JyMq1MHe7zoYz
nfRvk4KnDLrLhfI6Qg16FWfkPBepggWIY67aNO0l4VZy8cOoiSPbwSSUDO3sHgtK
J3DiewF6AwdwE8hVVN8SiKuKSbGmHnfPvYT3jpoUW7gmDJbB1rVOCE0LJe/BNSlG
MQdDfgl4k/bllvqxrzHrduN4DGsGweUTeOKTCKcOjjwaRtOgk0maqWel1NY9oPch
fDxoPwB3jiRjWqw6pJugxqQM6skyZgJ2M5WrLm7uARq4pZKUJlEaEZX5RE8Zaitb
CKB2izzTKgCUKuVF3vsCV/JTh4hIee1VLjNpCyiJxnMGTWG/bjMMniewuipqtykE
LsjAQOgLyNAWHtG+mqzpw5ssEkbNGdwuiv0IvJL9ZvemAqPjblpuUxrXMbXKt05m
CRwJEFoiMZq5NDHfaYOTWf576TbR/V63w8ovyOi81/b5Pgg3mN0ZNxdgnNocsJRD
G1D8zbktE5E0YV6HkPMEkSokcXG021Q7VndI2N5XI3kYrwRi0yGIKgLfqdaFopyG
8yClh1+13tWBiPO4Y5FEfcrz/3DgK6lXPZBt52gOWH0wAjIiJy94sHdxCI+aymB+
XA9MKqjE/dL684mTLaZ0n1MtCHocMRXhYOgHPuuDAbX/wbsp6SzmqZ4zBnhRtcDS
HUlUF6BZDt7FPk7GUPBig0rSmOA5TNLJIuImXYsffqRQBdC5cLeJW6xrCJuOiZhr
eLTtwokactyLD/harvX8gNzEL8kYA4iPyH8iAj22bsxPdizsVf4UHil7uaK/B08q
WM1BUdQ5QxvfZvEqHBDhDtd3NRMTrb4a2/mZL4mUWVxQJ/cZIUaal7O69mJicTCb
9mR+isP6uOQSfclnuumy6aXJTzGPbKXAT5r3KSGj0p/bQ72Y/5AWo0++wbl1PtdW
hRIRS4uS9/sA61ZAg6g6ech4u3MigQgkF0FB+grD/6F1uh0MUbB0z1Jml/oA/HNt
6ctBojO+ap9pBPyMTk2vgMeUOkv5PNR6reQjcwe0fYgz1kBsvaWn9sOKXn9ZcAE0
76KJHwdD1InP7ZG/+7H9Pmazkv9Wa5clNCCpctChsARoZJUsJODDNzwD5fNNaXiK
Rw56kS+vuMpfxI6oCA7j/tKI/dEc3u+5tUTh8xkQsByvbYSQH1nhxiiWWGg+glwR
aXNxDjuegLI7XVE4ukvDedbgZk7pILeqMJORK/fQIP0VrZ52vjaFkrHfLmOx4lX4
lfb6uRO7cWOyjrUw3z9ide6MwqN9R1DCDXdvkoFLlTCxkqtsHCB3y5gjVIwzsEzt
xyhkfrcQfarj8c1dg3307LOb+QY52n1sWjc+By9o17HiSVAJBCYfc7wmuB1symzW
Bw6g9UiGf6EH+Q6vXstiXeRZK3Sm3wIxfUvG0RlZleHQQXhySsYbfT+alrPhxhcH
9H1HygpB2eUBQp9p4ORx4heeKPY6vnPVj9FgmaGatxhdq0QSYm5Ihjrmb6Xj7/yq
fZbDnDSuHuVdTj2b6r/EEo5On6JK3LuM1pP4mFLjQtwn9agJowZIogA7tv17XJBN
BY5WVzpZVq85aBt4P1I1YQLvvHlTkxp02DjAIQIqxMebMScxybqIBIIZxuGj43zh
TKl2J6Ko/17TONrBmPRhjcZwIH8VuBzmsH6ATj1ecEEvYJTytLrNq4eGO6VXc4o5
fh6MVlxR7SzyZPlTaIvVjFvmD2Z8pPQBC8dQisNimQ1KpDiX9xBCDfMHymnVPQjz
+qAxh2Zw6FMYgzR8dCJ+1LkaaCe0fXlv2PYeHPZp0DmEPCgP6t85EGuqyqi6clFH
QaKz/Z/JQLETOMyKySbS4UJB0sGdcS+Xdm+Es5lw0HjF/PHyL2kg3Fy99wY4/FL0
gF9yMLkB5Gd/eJofeKJGvj99uMSzQJgzI5TyurbJMYcoSVaB/m/kZeTzikTWWS3r
BiNfLHD7FpChjyQb7UDccoX6q3iCAjihXywOwY3Bg/0a742tGpGTBp/LFAN6U3uq
jFfpF3D52KirpwHkLohgazs58RKe0LImmFdmtV9h5DdzEr1buGVU28sTZAPnH3ii
xZ1p2feiPTSdXnX6U8989YM5jeq1U7UW9rldvAPJYa1xpbbkLoqXLk3HFl0F5ZYP
xalRo4Hl125sIcrvib7YYEyCh6pbQ4+2SB8mc+qzk0yMae8ce863rxq5/4MkHA34
zYY7J5tEjVYD0agnYugHO1rWk03H8hw4FbE/ohKKtq/rKshm9vwcjVlDoFz3ofWm
SGSPmQbMqiZ23c1p4oe/Detm10cabT0kChJ8zhPVFOJGhtvR35E/qBfGu88KZIYj
AOB/aiOhcbyASEjdYHNIA3VAj6QuacXKIuXWDVqxNyVTn2wKx5hMJJe05pr/Lhgh
59JY8HX6ls/bSzZcb5fniarykw9o5/M7K9wqx2cAaObzkQ8Gw7Vj95CEiHXVK7q3
ephs5oNjji9MHtJOARcuLw6OHdPYoCf0XialhqbH8WJ0biQXgIzqXLgItapV4HP9
USlKcI99A2BQ+lnsYZzlUddl7G8FNvYlenbffiaMPiq9qzc12dGKpLh1IaOV2b9G
hTwjs/VidBUlM2dmbmufH97oOHS+A7EPGlgNttsTnAj2Z9f6vlbNxL5fQoHX7+6H
/uyUP0NXKn7i+fTs0eBo5OmTQdTKccIYqbaNRLOWgNqZHHmLHbKjzwfpklycLfiG
32gvB5YMxYXg83os6ELhvxOiGpc5O4isJIPjY1/MCnhsZuOW2nYSM7IRdqriyhV9
OsLbCr41/3XdDjM8vcwZQfqhP/YxK8PQ9WrhUGhmbQYmwQGgrTkQDG4SkkR7+MXI
Z04v3RkKMYrK+kqAcVgeu6zBdwu7kdZQIQC1c90qRj/SCgMIZ132d+QWNZDiTUZn
5y+rIMOkJ1fna8W5LAE3EEevHTqgiikEuJ4D/Y7Vz+Cjtgu9bZSJqii0NlYhWj27
FnEId3BdTJb/owk2eHAh6ahGRaYCy3gb8uIcAATU2hrFYemMxfDVyVGKliz1Iw3g
uqiXJbqQERlHaJWkW4lQ5Kj2eyoKthZ0aNWRrVehDJYZoCWu/iZZ5YDVyVxwXe3D
v2JsXNPR8IIhlKPrAQ3n8Yl1HcZBVBZlueAaIc0dO+2ug6NnglWyKs3XkIuYHfRn
aTWFuf4hncGl7vwt/5y7ziQyyN2JZiCebJslYT/DZ+seKZ8UL8RO+pTos0ZnpuWD
gLkWpTc8/jT8puLjCOit+LJP6DP/vP1Fvhj1pMxlBwQdaG/8f0L3D0x2g1OKvtDe
7Cx2aj8XDO95XBLm/LrgDh9ugAlY2EDSzAQ2mtXJIa1mGf9hAv0zCCoqTYKhqHBA
B4PY/VgIy29AhoDAy+KII6SqnO3QqbqtVeCtl24jKSxEAxChNzExrynkP7cb8gbT
x/cPCaPYvFP4EWTERw0xTdlirTCvFu7CctKXTFMT/BGnZ2UZ4Ycap9Xad3hLCC8R
RbacMRiAyzVtrzFBvRyNoQVpUU+hRe4dPzSGIzxinlgtWj5UJUVGeQOCvWI7RLZW
tIB073adhHpOPzOyBauBVGAgVGBq01jONmBz0IkUwha8/aMMCbFBPXs+zUTnJo2r
5knZiBtpXi/uc0j0Y1czTSImH2HWV6t98U4nwjIgAWw+Vg/vDuEboJM37opjJa71
DuTrQ0lwHG8e0n64R50vbqy3jCPSJtQneqPJ88JwNyRLu3iAgmXfqrcsxdgFn11u
Nqbqjoz/R3Bo+z5y3WmP13dzdEsVaKTDBOBhxyQz8m6AZL0IVBF0hfjfRiiafCS4
tKw1Q6AIMSrIKXLHUW2uD98hQO0ANXPJesfRHb/H8Lon3XTsekZn7kQm0C9+OSC3
vfM8B3MhUtVsFd0uRh9qJKNU2uzVymlh3NlavPJc0hGLXKSkzfobi11n36g6f9zI
/GESAM4tKQqACrB2IkS+QoWvhP0QK0uTSvcOkzJx5wwpgNPohxdmSl2GjUMz8T5N
YNFhk8s8wFF87pSpW1sQAMtz+nOlUb1A7bhwmgEhimlQ4FQkxXVRzueNlhZenuyY
1o7xsHRbpI4euc0734aRsiJwHC0KL/1ECQYQGxNU1YQTLxx40AaEWHTsQaOJhacH
FtgD5UkgM3CTKnk0LnTnRNZSuF8PUkUswJHXiWurLtEOhoY0JjNnut1qAlZBqove
F5brxiUO+Su0ruMEXGsUaqH261mQuK9/v6ZcmbHcFBnA6r1dm44CDyqmCgmPu6Ga
xEB1Q4jrtGgs3Qs/trQws1jSGCVgfkIdMGRPvbEInBqESFSPLJQzjy2gVsK0jy7r
ca0vyYIVpJXACyvIcMjVNcCtV6dSePqamdLsGstgBEuiUkGbhDD4ihECSsHtIfZH
Cwni/Q1XVXFIiQG5i/BHec1uEpDW+P0qsZ5FWpU6qZ7QFZXerxEbOLjwVPexZvRR
E6axup5ARR6OO5LFUTj3Neku98fWDE5Lr8LobCP0tVwJKD9Qh4IbrNftYyNFlxnq
MlWAc3FCjx5ENMmWe7b0xQcwrzQYGOFudsWRGjJJvk828aujRpMAc7JfVR0wPbvo
v+Fa5rIUqIiJnDsTNAuTzo5/EC3LUvGcuaLORx01NlhrBzLpSj3MRrnMT4ARQOcA
6UBCZkWJiPUSr+RVgyec148G+98OOvjB2xKKS2JfnOKhvRM9VWX9s1Yd6gEy3fbw
xxZ7teXJTNfea2nHLwNjs2umCpCiirNAYAPJ3fTsd83mw7PsPwlaJRXQFb/7+BT2
X3m/d5/thnOOfijybD6++JCDV7Arqh2KkveWIQ6iLbvC5nx/622x5BtIVpH5Op2k
Nlp8bnrMIm5LvZgRZzxi4TEBTwVMTNu8r3AMkUSDTQnRqBYluI20vjKBuIeHN4KB
5KrCGrwq/BhbB3fhqWNuobbMqcfyN64ApGRHYG3pfYCLCIY0zUnKxx2yAUwPKd4V
5F54LEJOUNFEmRsqRF4EHAAPTdBUGvMQLCRIa6GSoH0wDbT/w/Rt/nhbqNPCrm11
BcXRPkwB5eDRya5raCC6OHs9cdDVtLDG0g8JpGuR9wCHj+DJERzlaznwtWfNmKHq
BEWPg6rh1/vnep1u9oVowlvEhgxdIH7lRNv1UdsCKod7Yc4jZ+Y4U/ntgrYdNBCK
YlKtI2G08l90nGqg2XB+6geSv/uo4+gH5IN3283Ucayg+ddzsfyWo2ZC9cOM24qg
97P+67UnYcypvS+7XOQJcfeqz8Nla9WsYWCKLvLWRn1F8ou/AczX6Ag3Kp7tTLsi
mU/YNPW1VDPl8YTIdvOvBTjxYsaOm/F5FTHY/SlRT71XHUvGB3g6KnM0RGZDTn33
6tzas6+HDVVxS71dTyZJcsWpG+HwMuASeYEgVdb6Twp6rJle1yqJyQpQxcXYJnby
XuaG2i6bcqlMCXcrKa4ulRTfQUK3Y7XqutMixsSpY4E0K3k9sLTyz18uOmUE3FFc
w6n+rnrq10zjJ2SrEhhu9Ft160wEJcDLl4zqQConpyi5cx90rgc3oLydmNoycEpK
UXtj+v4D4Oz+gLZ7WIED9d/Pytgn4FJRkLqu8/fYelH+fPxl0wl5GNbADx/Q03Wl
5Epmlu1OZNmFMECQSNkUbwFBdaBIW5sQxKmLOqxSiLKdoVvP4IyTWX2r2es2CO/e
+/xh8PRcL4zku0QS6hySA27yqHxDAJOe1MoS9iZTxwJawA3wKF7TKvJ1xsXvFCFy
QEXD4O7GvmCa9knoedOtsUWGEXsRG/azAnxvz3iPVnM+eewDGiQlkNRj0Au1z4Xn
LDyq/eC7ehbPqohbNziHLn4EKh1+llD36ih0z/sWhkfsvA3Q4SKn9LrCh9s13yQn
nESqgqHaHZgf1eCApqz2+E9Kr5mJ4cYRDcvDGelN6FPgghTjf68ZNP68Q4oQsEBB
FRkpzCvHrXfa7Jt2jxamlovJTj7GaX4UtLDmUI+i0+1rcM1bOKllJYh3DSVFAesp
Do1bwPJu89P5IDhw7L8z/5krbMCVZcBur3MOjK6kRxRjlFm8fAmx8bBWhg8E+qgv
Lgrwe+ykv+nn29swhaAKCFB7LSmwH7uikONrBMjCN0IHcFhgYmhhAmqRnqfBQ5PH
bYR7oz405nURs8YOV0OM44eoPSihgy9XAS9SL7ciFsj0hHvbGkR0IGkRirP1BmfZ
AKxoX76C6uwHiub1YSIhXY+HOEqCWdvWe+y1tvcTd32fJ1aLIq7FFByavkZadBX6
KfbxOlwrbgCOX1pJlOoViofpFEtx0O3pNzKBv4AztLb6TH4bMT+hiBMx00Cp5IEI
fnJCAfWgKcNLZ23xVDQcPMUekopmN6C/1V+tuaBWCiNlzDuAIvzaIpe5mBrSRqFK
stqSiW0GeaJK77XoktdZOcAPkmlbhmNlSuoNUPzHZz1nJMcBI00LrIa+nou+/LR6
rmJZE0cEbFFPVmZoGck8uZ8CHDjcgPesEzEvqdrb7071Sk7hRQ6aE89azVfD1aJ0
AFNyThzcth1IwHtOtftoiqcRoWhWM6ox2EMDD08XsTydb303QKfVLYSfrHji5E59
ENzEMNl0tFNDebyYOhdlrjlfRSWcf0a5bj27En4bH8gXlz4cOACT29/vpDFe++Dr
gKVbCHy4UQavBlLfgAucHbrVj1PvH8TNj6iwifkpnCU0KLkh/leW6Zs4FVb40zqT
1RF6Fefsxx94bnrv1duD9A+NKGAa41mVS1VfKdAzO9ZRDbszUP5L/8ZUsMm2ggbG
Qf5C+04qQitBnxpifw0Lkd5Ex/GADDgi91mjjqPOgP1L+KnylAIrkJIxoXZAUJLT
Fzbj+k52CmnIT+qBZVuJ5kezLoMCc9eeWruexfx9tWlC9QOB4CWXvLaPH1LCU6g8
jgeW8AGbDXkZSjmqMgQAH09OdBMtAXshMCx/qJwSH1/sqUMDxcf2Ry8VwZ4T5jjL
s8WnzcozMeMZf798pUTxnw1T+ogeL7iCOy+wyOuLDTntcYWFRcQLTz5rs//BXAas
K2X9w85Tyd9JvNlSRy5S9wuf8GyPHKCze/KhYSLDbmRiQtd1EXXdSnjER1uxQinU
0LBqcJPwZuAYD5B7rabSlK4OLl7VKSXFdK1f0pWKBxzYIW5Ym2tdobYDRwLy1Sxg
urBHIdxZib1DDmh52GjRrVO0O2DOd5j2ue8ztgXylZl3yRk4PGztu4GJPixKrVvt
b3Bk5r8YbCcFxWvY2EarXDEXT0ovBLtRhkN3cdWqKRpDTFNQW2jF+xP5SBnTFKtJ
rodwXXbhTk1pxmAwivxRubmAXvqSNY79iqsgqIy861hJ5EANngDHy1YDODCOukR7
XDNEUMjZXxxQTyDcMLfUUeaXPQu/YI/6x3/GwcnkBo8cfw4l9Q/M2kCXizk7ybFI
J75c2mC/Cbd93tGTnUQ2HI6sU2U6OkF+QVSaqYWEStMLCqcL4T/qkfBUqIcFnfQE
ddjU26AewdOnMpEJxStOWg4xl/sGpLdj/fKcr4tmcEKImsHOCv3bMZIKiYABbPo3
SvLsrtvrrPJ3913/olKJR8yw423y8WJXSikqAsM3/tGlh4OycwKQO3q6uOo3cPx4
5Ec0SV66uUxdUCeq84g5ae87oCw+tDlG2azo+rGRjor5mFbL16iN4HbhC9hBqy6b
KeRfae8nw0qjeiozxK6U4lC3eeQwZ8pucOP/L1o5Z9QBVjAoYDfKj79TmwKl4O0F
37AH3zeTDkItVBvTckZ9VSJJcbbxXkzWFX6me0TCV27FFVYY+4PI5zx8WILPQENG
QHy9XJTh8Cb4/PpxrmAVH1EBc9n23KkESZRKXwiWiLnRhRcEzgSZH4jkWTR6m77H
oYayIBp2ETKYnc/ONRVneY+KwCgxHASHzC0mIww77+BnlvCIZ1T5WRtEdNckCw0X
4sLdWdmhhQLJmU+o9ZOWDvebo88J/oWdU7RMTvyClX5Kx6qYO+dfUD97/MSHTEwJ
efMQoxB10xY7+PN/ACXn5dwkr29l5lif0LNm95ZW/WX3yvlmDWzorj9o2xdHpLxQ
1KrvtAfigQ9MRqpsktliB5UQ1aJXZbeklkM4AMguK3sq9BpukTW+GihepC2FnAYC
KC0naqAFuUGf2MErYa8iCvLz2amZJmGKt79N8sZAHH3wLMlsFhnKDvVkCw1qgAU9
jHt41eThmMcP1grObE6CmCGJF5ll5UssAoYDkvAJJYLD4oKJhJUZk2ecVkmiSdTG
z0YVv1y6ZkNzNYajpdAiq6I0pMbhMsz1/8q0RxQp9CGbYu9kfcoQbfgZAm30Mo/C
ABw6C22i0sjnfJcXKYZ5EUEV8eFqUI62C8oHILdVng5vn0iIGi5zl86DfMhNpDLy
2+tOvCAMQy+VR41Gw/+9C52XTo72zydv9YaV9nz5v79ynGA2YMYRHVWtBtkjftkV
kZcRqh13NbkdM1d+yV5Fei98AtE53kWZpwoPBNlfNFhNBK6Hah/40kn1Qg8iUEhk
dHZkSW1Rj/YZpoJFpIyvutoMaXlD6A3ZFONfc+bf4g+SJcTvgkU7mhYwcBW0WLS5
yRvChyrt4mxA4hV0xNb0COfqd+dRz19VLtig45ssU7ny9fVDhb4MYMASiyAHsmC3
BQZD9KKUdiTDVBXZoUOU0XSt9ZEQWOmhQtijSiSdVMxkrvBNFythqyYN48XO4A8O
VpLqMLEeY2GMPVfmsJjZ23OSoIYKewS8Qd8nlLPXTm0GdBocCuxKRY2Ow0CAQd+3
nMYm7zuXii5mHNsR/gdSgQz6MIOM6n1uh/p0iuKx6xILXkDQqxKNcN19BX57l0fg
cGGe3duBKmjZOfdWn9y0CVtWC62xD2sowcIXmAYzG07OBIVnR0ShpHkxzdhsEh2o
FB/iFcKbU9LbHDwIIp+PmPW3Jk7jNvdaHHpsYtMwl5SiHrLeZeDqGEeTqdpmpOFc
lVyDrymatuUnnYYir2NeZKqIGlJTYkA767Lk32Jph9CRh7rXdi9QYnPSlE4DjMfn
orepd97lfwy6rj/jjcwKAhLkHjdYU8gLsjSZ59/LYTkGTaTYmEAtRPkkkQLBPFE2
OrBzR+T0vtJ6b4ygusd1zQkEs44MuCnw36At/bRqN2/3kRls4MNl2pMNkoub4o56
5pObphpnHdL9t3B/vseUbIDjFRLmUu2k7slIUDcMwpEZ6IAe20Ip8cryd0qsgiMG
tanj6Bhj9XaNXJp+LqepATYnYKJvCs5AdkgufzxBY0MCYP4+lev+QvneoleZjjPo
kONRVwKgxonDMLQ+kFSLWlKA7jIK1puKZ7eKnB6DHprkiJK0QVm43jdNXXN4ckJG
I1IRmdJPbBmQarus9NTqDzToP5Th129sDqIySqwN+3D4ECHPNY+dHIMton1vDmBo
Em2hdV7TsEyVViOudeiEc6VD+4itgetVtFhMa7yoFZVPELktwIs5dB8uqiCkNvjH
OeGaKcZTb7Av2ZBGCYVs0ve8+MGIZdasOjHMkfHmaYMYco0Er83gaCAGLDcB9g7+
xgYhha9Zu0ZoISarcusxWFGoLAfLCAJo5bFQ7dvcA+e3CohD6gwmCm60WAQwY38+
+3fbfleW49s6Mp8Z9IAZhaTt/MmxZX98kAjZsAReY2VnI0Ccd1lbSliUlYkx7Yxp
a3bLtw9dvkoFB3vnapiGOFG298hdpGJe+1oL6klpmodYZAdPMOEJpDddYFl6knGe
EMwjir1W1spFh/DDeI10AOwQXknyfHEFm/8IrhyoesZp3pbYuXSQ/O1K9gIP+OSU
WjuBaoEbGhQM2KGVVydjOZNHBDblm6tEj6IV79f4jAl2DumA0dnf/RG3jpvSAxCp
orqPQMvqoIKwhcW/9W5Xxi/i09tZTKlcsZUlqf3Kocec2+FL4nGTuXXk56C6DaIG
fwK3zxjUeTplPuPrVeXCJwGcsAG7jTDfMeBn8Plisw6MovkPsnhDqYQzVlkdGUz/
N8jMXDspe6aG1LbfyXnOH8Wu5SBBsMPYGlJeV5M1eJr0uhrmdDf/CCBqjqKZ1HEo
Ej/KVLUIVFlqGEvRfVXTexFk3oUTS96I2F5LJdk/mhakGSQFyqj5+x68AiZBwe5T
PBgODwl2aM1W6l7Jn8oFQWsDiMC2A22Cs2ohE4XfKdJ37XX9jRiy8EgMOpWw2ran
5iy+BqL/a7SLAcrm4axhFtga41vyqDjXR/1rxNCMN6a0tZKMlMQiA+PSJCXHbuqX
wJ91d8JeJW3JL+PM7rJqlNxcphxlm6weh2B+IQyTUvxbjxNSctcV7vFXnQ/uEa0x
XqKhEdEyQu/ZIvmHnUgCONaqMMacE+DzXo4AqPmhFi7b2q1KbeQ/QDJKEZrRf2QW
dPdoT+Ga07dmjYBvCL6+ULnJHItu0TI7D6vHmbAvZjV1d3PsTwyNQDcrPhFEGWE3
QeyQl0jxvvI8XCGiU8j5nOO3aaOybS5yyQN4bDTwKy2t/H+kGWzuwEP0CHcLC3fE
ODDN+umktFM3y/NPK8H56NQgXw9CFWIsr0MI2N7C16EnwENrTuZHankcCq+hchEO
PWSBZIW5W1TEmDsLrz/qxq2MCnzBNGnTK1sIWfPCojYRrN7bGoU16ikBjGKoTyBM
rydqJKdnaNVLUTshxXEpR7rUhPgpw63dKhsnAb5ZTrjxGtzMoJnOjTZ+8Z6dEEp7
0AyHuOhCTw3Xs+islhZUJyVVgIK/s6WA8HyDmOPVmcL9gtYgNmAGP9JFH4LUmdHP
Qvog6oNGJHIlMIVoNNsjQdBqAKCi1VMChz3NWMX0VNzywjChZwE07173h5EfEkC3
ZejNdZuNZ+edPR+ruWSIVPGoLI/bfpHoBu80UTNi7Quwecraktu5dSovI7bNheK3
3bXbmtHBYn27TM/1D7q+meePFvB6AzyBwSTT8oRAvZdxoIuJCiRFsdtGst08QLNT
CnHMffPkrsTuUyi9+Uh3UK93rI/3UZkFUZkrhAhMnO3tAd2ZARY8QI+6Vyx9TdfX
NYbrojIpH3FxptEwMJJr4qMjo2XQxOuTQ+ne7CVTEnyUvOWuqb71eAQeXhxJ+ciE
cmpya+iCZb6bEcbHdui0ldrAu4oE3XbT2sQvih9K2red6aMBDygpGp2OIHWa8ESB
JCgIIhI7B8qJJuHU39DqkRrJybQiXWivU6gWCr8DBvUmuTBQqYdmdSOkecwX1jit
GeUWG9gQHk00iNkPSix5MLxh/MgmY5i4kNrQglx/wpaXHXilqBGvsZJxXL1IrKLk
2r/P7E9p0pSxxmBati1SM7aaj0Z/j52wF6mHoMSomLs3GQfVyD8pUiJrnc7kSZxM
9FAP42bUsdQKUYrnZl/BipWWd93FHmiRcyimgbFopc0Nmr58V/uriX4Zeq9PWy4K
GISFqfMxxnkN1TBlF9TKimjlF7wIZYnczLRLsNkH12okliooz9fl3sCI7f15et6C
sA3BlyjU5ngioiwdcTYA1dd71iMTSDEIXEgRBO2IjqJ2GEbUuuCXVpFE+NLIEvsK
dgvSTpwpuUHlyWPoaFHPJRugkBp0khtIsHCVJwB9YN/GIP7ERTiBF124B+j8j4BX
/BJcrStrXa1kJEb+6AzjyKGJBSk64I9hZt6Hc0iyD3puD+D1mR9qp0VJ1qABctBw
ZKkr1/8hAul1Pfbcz+EVUe3DAjQooPef9xPYs5ZtC+Gb0oN5mv6QSltamncrFnaI
/G6bInHVtK0Syp9HbR+t0CUhsYiYkjFqYKg+xzqRs+4dUvNG3roXF2a57twr2HHG
1KauxWA8jBh9VycLLH3vI7tQbgvoVW9g0jpd+h/+ImrnXY5XPi/9h20WTwEuPssS
A1081TJjuqEbk/vZKIdZjzhC6GXP4MzULN/D8tj9iLeuKK/98Vftf2OOLw+6q/Tl
Gs/hmlns4dbM6LCMLwZbzwVRpP2rHJBbGbUPPjf77KB2XLm9pMSBboIlnu4A9wvS
Jy4rjPkxX88anlebeJITCxCmJFJhgw8xVViOPoAHtdcAqdD5ELnUTRUA3aivZDCu
7SMexUlCYC2oztxLA59IMoOiLPETXcfqQFyoA6HIzEILoX5kT4+ZqJ/S+ghsM1B6
yhHRyBDOUOBkyhdw6SMhKt3kMKNsljkxeQ32U7p+lEPqalbaTv7RtCLUjuBfB7Ot
Rcj8mDzm+7VYF0rkmYLCLSbPf3Zh/n1MXvOb5/QkXmbRAKDFzhXuTwbGCccoElrh
QfsCezANgnzUlBKE81+nBt41Q01wldRkOWYR3HDt8mMssH/HNdAuh0W8BNuH8STM
EbemgALmafVJ2wVTVQnR9LgnTo/oJkVpdablc4n+Sv6O4FEX3WXoVIAKwa1sIUwN
UvDK2rCr4qLj9/yst9cqOJbkR/xQ4uoZ+rWJQ1LdYnlLVmD0O0BQcrX7ex0271+P
VILni4CS3/9cjAopxolS2PJiaQDk+bXJHyLkMY/+8BLAjstmuVsrJybsKlbJXoxb
gOA0Y1IUoa8cqAXHkhiql9oAPMSUtHdxfRsbolvShoID2OzpOwvi5OUtkLTDWGlo
xz06PNUnlXRrpNJxf28GQIshm7FXKuvhXcWVI0B19jGE+U5wiE6S32uy9BTJxeAn
5o0MXr63QPbk7ASlfR/5GiyIJpeUE//hStH56DW+d6CfMrH1mw5gz8UUZ9z3cYYz
tWuJzwijYNNPi7aD1Lomd+U0XnCEKOtZyFOWqleIAhB8eIIhgATpsG+89WcTsPEL
ZEvkfFJN52cbf98VnBotz20DtztaagbjHSlRKQ3M947+clktUD3BlZ7RinbLe4of
SYPJgISz12n6N8tal3kGXQ5xs2QodMevYWzut0xZE7ZXwugi7AAMB7PLF22if6Aw
cApzo/Gp3+/Q04qwRFlZdi4muuQI7xwQvcyP4noPShwa5VXuFuFJ0VTXKK8ZFMKu
/j1cFsxVpzhWlwHNv1f70/tivr9RmnpRvEqSCNbaC7ErI0n5Z9/ops5ddq0il68f
PwGKWW0UoXcMEyhzHlCyjZH6I74qkHg7o0628h9f3tjd51VOJfr72DRF65bA+4l7
mrNkDvkGZJ0FLNEylQAhzTlXKR4f2NOtBmmiRLhZURi3DuI08Si9Ijf+7zc0pn8s
3uuQlQUl+d6HEDGcix81f/3sKmuZudDBEXLHdhjy346vN1GlhDYknLM3anXjKvV6
wbFpovRdR8xeJdnTww1Z9iATtMnUQB8V5vDI8y/sNddmlH5lUUrJArJcxsa6R7Vk
Y+G6Ms5No5yXRF+5xFE6g29zWk1LFC30wQ7yPsz8DlTG0xJub4lYwFZY2GMMMdcJ
3vIHVpor6kjiXMVWlLiOfuRXe5ahF/IHv2+XxE6bF0kYzHfbOrbpUd/7i03Vhjow
HwSKQAAa1hYuEaDg16XPBKHnDtIu+D7i/plqUUfeGWb53P1V4bS4L469lXsUBEQG
Rna/mfRAUt+S7BT94S6P/SEslYatOc6IDVqBKHHH8R71mD0F1cI2u3zAVsgm0e20
eRXCOiUjCPT3tBcYqQcUn/CcZKiGzLfl8FWgHH/wtOBBjdxugp12hUNbDwdFoSkR
RDQengRPHsRKlesvR3Qq6rBEHPHlL+0IGamZjolVM9rarpWkQvUkHpiPVIDIIL+8
FmPu0zOP+i4EHZjpbn+6uOgOLVYy+JKch4OWYXfD57Spj7O49FidOcr1ZxGGl7VE
A2HFQhdxNSndH90zydcOppeDp9b5xwgJkgovKcng56kzfoFdvalEOPJmDixrS8vi
stW81lEuqIt1Y4nh8ziDgWjyz0EwIcbssYguW58onKjTlcJUiLuHBYrBl3uoHs3a
B1b7LmxclJoVDGMOV1Q0WeixeZHZxuKbB+2Y9R/P10PiSSMqVJIUmJzaUw+aa5iR
w18qfxP69of8R8aIthCeLtMWUsZx/scUMVOkNAsb+y9qzmKA+39KQyo0uU/Bb8J8
gylvWgvYgTGPxkVpoW0ocJt8G3ftAMORNlBRrNLDiNYdQEtWOZldN/FEVkDXWC3M
gMeNggE2rYxMTDHZWtzUvalLT+8nDPwK8V9MIbFDJxcKn275NgljkMwV41r0bWxs
7q5gbCKl0RK1nRyHny/3g92KKhHk4pa2eIh1bG3EAJGaSd5FivdlYoTN+yCm5UIs
zG6Sbmik2W8AHwX3wNQ00rHgrGCeF+TozTNTp75QUdg9wWVoAGuvwVkIOMNWO41r
WJkXpQ9jCQbL0OnQGu36TI+Ytn0bOMokKBYXI2j/SoBCC31lQGqlOvRhy6uiKM95
uzJk1FYuoZ2AS4cB7eatC1Im34HsLbsLm02XarTUfsJ/RTaFETkYrc3iu67e959J
YdOqLzmVVOXY6uR/xtTbyqKSLdzRBfZmLNsVSZPIQAR8goOG97jg2MC3N92Z1RbM
8v83cMuxKaUV7a6EQK9sudt1w/pLkPXQXx4Gg3WMhKW3leDxzby/JfRiqHxkgzis
dNvafg3tgQ4qmL6GZzdWDfN7SuMR02DnuWFF9QETNya4rAxVfU1kzXYErlF8llcN
hi71JkKzeOORyHqwQL1MeEFFQNf4L0/J56fLvJBGsQSYd4nT7xr5a017Oi7xG40G
OV11TmtCDoKlHjTy/FtkG+PX5fKd/QXjHhKa/hjteOt8eD5apLgzSkaLBqihCYGt
2KoZYzTj0Cl0kNyXATHLeEjCrUq36DZq4LY0+sWQA7yD6Jo6xLfPuKBkDBFmwM9F
cNoB38SuagIPaH4edgIvWoOwMYSQ0BL37NKPqP0HSApV5Jmb8M7rkCN028feX1eG
2QA4tWqK+IV0807l5W+rA5Ua2ZQdlQ8WOpgroDs0v863Ix2AB6UHiILwwHPX8QcC
YQVoyYem063cCplRTPncKNZ3zVyqdpk3ilfbZLO/R8QXMRz8zrUIYg49LXyukK+D
wiC0g3KZUnO+Awxb7vrtCwS0xOM0YALbKh8E5Lvizrl01P/uVm80fXLWCglysmoM
9rRCdUsbUQqgNaq400hUIikVAUHcpTbNQW+rcSwqg//18b1jPCLVOEWceqE9NOmS
cGR+Y80xwcnOmEZB83Qsn08/wwBCWXnAbEpxjmWhq4S0PcwU4JC2ga2gCnCG9XoE
pAl0LTndbBTrcG3GJAYY/hmWhutlMyqayiGT4/31iyZzao4i10+a8asXRVmpjvbT
6BrBbLTZyVel/fFKNxgOwG8KP3uOqPj/Xbx4GCkIOhNUUNRKQepj+Vli5Xu/Mfz5
5CVJoGCj0mY2By61r39SqBOa/w+YjkbVrZfS4gFfwh/iSaQKfjtX4LI9Of5dDGio
A1jKqHrYXUqXZwDEpiiW2SQZr8ye4YJ8CasxNT2gQq5FMcWbT32QT2XfVLHBAYz6
HPF0XVSuHjAdetI+rcaCyd7L+k51Fh4WzwLsL/Ra96B8T7U0u5i6pUUv4sVAc/5X
gd5c7Y9Tx2WL2FrVz7X7jZ/hOVRcsn17ZDj+vrkxDX8TrPBC8nTzD+Bhg3gYhxYT
cCJ7dCMeMAKq49H1CQsc+QDf0tetKvMwrCuhO/PJMRrZVq8F0/7NVBjShgkIUh0Y
VlzaP0gbySLFOhvq6I76ywxfCoQv6tzH1O+MUPtGiwfM5hNaqJNqdpOdl3ArUam7
HLzy+AWHM2v90OZRwWu/eqBBUWGpP6z85I8U5YtEVI9pr4xTm384Z1dIW3bEjwbU
PC8kS4QutftRRm8EMkqhAPd2Ky7K78Lr/BY0W9x51yNngj0bCDWOA1XYfQSvelgl
Y2NcNqYYTA2xYLybQyuhWXKEqnE4/enmIgPn4d96dLcbr+GZktERlyz0W35dUb/L
1mg6ZVR9FIYNa8RTlgsuO0FxEEdM9KcyIXCRT2KhMXN6ioXaYEACW1OlBIP6Gfeg
+JcyZFkJGj7am3IdI0gpBULTTmXdxi7X+dVE8jKqgjbUY6tHiZD10hJsUxBf3mjH
pnCXOzNwQRIbo3A7fmdOkEFbzqfCyuA5QcJqeMJ7flAovEdcZYrh9f4eRQzb8qLE
VTaCIUEJ/vOb25BIWp3jMYxpjaUzjARDd/R8np9K+DL9DTfIntfZj6NjLar4HN8z
4lRDxxxTFgS9DF/QdRsfhIVxvuWKuIy5bYIzmkU5Pt81yiHOGweQLXe1075M0Rhg
j0pTgilz+dDbidascHIB6hKUpnNebmIjxOVWxwk6So8whuhr2+3Wr87Og7sZ8w4q
7vSDvw3z3vNZXYLIdCVse1rJEzqqZ2gL8THReC1hGEivBxxsUsjYCQ8kq1dsV2Ky
cs5FMRnWLpeWg6ugbn8NUKmEy6SUuBUrGG67GiPzleGbzg9SM7y0ALwM3x76b3Rm
XXDdO4RTtjGDhNroZTFJ8EbsbkII6oGsk+d6ms1pJbMlw3nogTEoEcwaC5Jy8+fM
NZLSXKqqKcw7JN4DCGQl22VN1uQ8AWdSz4jolg8l92Ig3lxLPdH0mB4B31vm2Rc3
aPlFXJHKl5mBb6HDWLZSE6mxGmt9Ut2G5AV08JHtWgRa+ZH4r/suU37Qpf5aHthP
eRovovGu9wkb/V1URsUTCuJIlJVypDeozmw1r/POq65c7e8aZ3hKRWNlidjnTeVd
HL5h309cmU2YdbOu5nXpqNLwqTHdazkKUyTtJ4Ac4ROGOzrHFnh+QlV9PPSaM9v8
WMUoOeNb349+jvQXvmHtWa4L2PQvYm5oO4QGTcSsHwYG/UKjoUQFUkfJ9R+mPEgx
amONSt7DlKQ5bwGoINYa/QnyMIq6rjYsN2ieHAFhfeIBiSkN2BxnUbMePTiJZmw4
3UreMh/QWxo2fA3VbrpbrIcASTfBpnIGMS9tsuZjSv1/2sGwsgHp62PprRu2QSsW
kAFMI8ZwTu1FO4v/ZGZ94ocCV8S+TGVJgHZTLm5xkCSt690oXD81498mgX8k9Ov1
Tu6/MKQxePFfZzOx50IDBekY3EJZ4hUcM4d+mpkHJUBWnv72vSrkL84/y4buRnMI
Q+F4LMr+wW/8iF5SpMlrpEMyrToBs5bXzI+Ff3cQxTzviRIuUS5085IqCUrUmRpL
k1WCPCzNR3J4wApE1v5eytQ0OyYPOd2eAVINxXjU9e5EkjsrGiZ84RcQxXKZjVD6
AsIag106h7UWNtb2sh+A7iD73K7KcBNaxQz49n/fGA7PthdXK2aesO2YrSXH9cM0
thU59Nr7c9js6E1kljXlDLPldRu7Doy9khXETPNye6NMPMzN+Yd7sfSNSQDH28Bx
qabCyslidiR7wLpnwEAHJ9/sHggVhKxkozB9lxRTz3OSDGH2J0UIXkgv9kiqcNhp
bZLUc68eXas7K+t764GhGsymKJe+nzKWs31wFK57F+p+9+zylufOEHch3ISA7GUA
3IUrwqpVcMFE0muIYJ0BXMuHQsDV/ACxjXsWvzm8F4ZYB5AeDMMB0uEiXOqpVd1E
FaoBeTVhMTfFJBtlzWepI12thiM6HZsRERIkJfMq4B2aVeOB57A4Q7HiVf+7C97n
iD/DkTEMjWjYEgVj2faFv/ebCpudgzvwNqHrZo1oVKmJK8FQl/3VxGpyG0wM4pZe
mS74NM9sYh90P1F3iRON/EWbSWmbtmvSs3wzmmFNX+xiJ3Fue/LtCXc6RK/Yex+f
zSefPim3PbOjUJm377JynOogvTLz1ntxgWmbSeCe7nWHuXQXtkMmg81EtEEdZ0X7
uHW6oopRAJjzePkYyYofOhb5lT+O0AVTGzCNlXqU4kBjslHsMvqo9OX1bNQm88fl
TTjn/tTN47X8cUrb8fykaXM0v24F2/R3Ex6FiGquL0sp5Ij8LYO5yO3z1kP8xSWY
L+IRJB7aCSRaF6dInzlK6o3Roou2zzyPkR4RCvQVyoCWl3nQkokb/t892zwi7OPp
y89uK4Xv9y5THlUuW7fL9DqJrGqrlNUtv+EEmNT6Mo6NlP5o+zb70Jx0JpODq9+i
YdpGke4ry/HFxtlIRZJ6aJ7O+mibCiSRhBe25LkEnccYxDgUiM9yJ/8wkLIMB4PD
P3DlVTaxRFJ7uZZOIYfMizghnyYC2GA2iX2FZrL1Mh8bHyljnoCsWIAT+UhVbxCs
9kNL30Jz1aDedTyIT5Z2yvzxBv8tYDxGP9pzqGvraauMHyt9oEg8+I1c+EwynULK
VZHVc+Pt5RapPM6k0PDHV4Zo8EziWSn++6216HnXMw/FgGyOBoEUFcx6lRIs9ElX
9FdML4TD7WNBySwoRnncu8oZlqEn+GB9M2glJF3kjK3daJ7cvCJ6Xnnr2aRG1BIP
/2737U1/9pLFgunC/R5YmjzT1GWQ50x7BNR9vad6WF38Hp9odaohqcg7+hX+dopR
KHeLqGYDw6cGeGQEceTCt9kBpxk/acEAuDqkCv9P6PibMNApr+q3USn2GR6WHUP3
xa9rqq8XsDZbNnACgF+0/ByCXOrPFkLaCMJMtaLVg4sZ0oRSF8xagPLswDPNSDaw
InZ6Xvepop3T5PHQTb/4tYPFpXlY3Sk7DOGddHbDOrsx5sEOWH5JoyeHi+J7lEP1
l0i987hVxBPlpmmfH9pcNlpQkqSZyEptnn71IOfm3IhXsVZB3V08yA9WCgZYEX5M
gtVHqoKHl3iCpkyTbyZ1kv/rcHGiiJfPLjyYbMDsnnmWY+rRwP6xE3TGD57KuWrp
7Kh9yC+vdQz2NQSUffzcTV0mnCkctw2fEszL1ErerxRFyUMJMg/9Vrh8RDa227aU
W5LUm497ZD+azWuad6rCDG+oooSE/Z2P/tz/sajOtJFhC8tC6LEPwwt+Oa8Lm/n+
RgiphBNEAV5ohBCjrHMmMx177Fy62In7gn8jHCW03GTfLeej5/d0w7RnuTwdygHj
wRwFgTcLqHVYgF3rkFvZ13gPeacVGbt5lEtoQ0SJFFLdsgYZ3Hj8ot5cx3TppsHb
e46OEoB1v0msycvL2vFLbLOW3giVmlJjR6NadXdPH0UE8PJwnsVDEX/0H0Q9udcG
zzLn+3G4w9fO3OK6csfF6+R+1ZCi77Hf8Vb6EE/CivW9F5VYjKPjKv5Dw6qVQe74
BHn/vQHVY0KMBZ1OhRkLcTjyUvGJx7F8QYwGdoEYrYfoSmwhcdFrFxCmCgqGWatb
Zpbww0JXRDeqTVCFiV++YyXlgL5IzF32s03uFytPxV5Wiq/MjmbduTvV+n5rrH/l
fQt+cvhhyVG3aelQ8bI/b4Lexi8sc2+tCmzkmSU139r6glvNKOjL85txyfqXspeS
wOI1Az2pxHQbKU+qu17dP88aAIc/1uQ4bDhEwoodZyJCKd8gdbDJXGVKxULHu5wh
C7fvCgrWh/xPZh21nd4LCjDdmXUisU3iNmQ4cTiu32RxpRBl5aAlaRe4dAIAg26W
/XBQ3m0NMLuq3gDPB1ZOqslk0pjgmgi9fo2UQNgBAbLPxZCN/9cLRwwwlphwNVw+
+x+l3eP9ly4E5eliHZ7YJOAHHH0l6Jszeu7tbosYq++6n7ZTnrbHaaVAx1ymCFPc
R3uLuQAysw2HNSZmK+fFR+aaxVd3xVXkgUILYqMHvQotjCDiBdUAdGd4vlv8MT5F
WFw6yBttiYmxBynIQ92FweRrJWWXYIwdn4JgsTlB2jL3E6+xFGl5dFVvIYNrARg7
+ZL3t0CLjwwW58MBD0H52XeR/jjKRdIuWsl/cvKaCA2Kl23pVmmFE4ohnc5jZKhx
tVYrJMaklEKgQTTeMITpWWnWyNNdXWctBN0UKCeoBj6PqykUM+dwb2qPxgVGBLW+
hzEvZDLd8gltZLkhMiEsDNG6+AWyih1xrQZqtjfK/Jg8lMCEicsS8L16NdGMaIpB
W1bcSUTuSJgA3/qpWebOwrJG8FpBaglqJx65GmMgY+gTTMCwwcG5daUaTi9VF5Zq
z5L0l0GpIkLcTNjwB0002pOX59VXEYzTDtzNmqrPCu9qhv3wf/jGN8j4nj44l969
z3tbl7uu8Bg+xWZCUeKAKKEewPozivLqE6bAA0i3F2d7ozRd1Mc3cvZHjT9Zm5vx
YHHBSu781KoZtB7O8fWe42AR4fDdg97wB8T+nMMLsENalybUt7AFxHifipfuzQwX
nGUOKKKA5sDuCfUE50NjBB7/Xb/0rlrXb3313Zd5Uso/XLi8hOB/HCWG0LP2hUJv
v6pK6HFJHix6tn6Z7HMEj/GfVh7wK8ZF7zZkklZGiRoJ3ROES74dmtG+Ov0UMe1r
66+WOhNrWX6Ja/m055jxJ/YSo15pYE6Sb7i5yWHR89n+GNUynUkVAnRjuUMr2bgA
KLo7ZD33ak1SShGCrIWSkzj94igzEV5+1IKRfGWiJ9cBH09X36ygTOhn+uwHIkgQ
bGNXzIStL+UtI4g7H5ee3IRMimV71DElqMx35XGeibpx4SJYrgXUrEo/dzEn7QvN
NOjqES9Pde7eCLUzFLMU/FIIwQ+sxxogv1de92KcSX2rlNGDuOijJ2qDFT7etaUA
a8Gu1u5cobjUfAmjWHoh/FMPlUBmM9CySiB97HQJQiYPteeuumovWlkExa0POcO8
1yFLSqy4zMH6AdMHKt1KLKQsLp7H0JQcZSrD+QH12qx1PtNIxyWXBVUlgBfXPDYg
PSEVUAbVaWyzFNl26kh7qT6k4C1NNDIt3nQzJZQZP2Xa3ZOSE/L/r1V/XVRcH1hh
+lSBjW5KC2/LDoV8+9gmv8ukHIGL+/mryj8FjRRjA9Gfx9rOyS6VD0eAAHiy2O3y
sJhmrGijM2z/LobkrSP3pQnAXPm5v36CvnmgPPBTU4GjftkqKWSv4nbPo2N3qtzq
0LcSxYH782FPYO3MmakYBcx+/+ujNGho16Yzuihyf5hzv96ILp3EGLnaSSd1NJa1
FYUTY9CS2Qfj4FGnUoI5S98HS0Aphm0jW0xEJ4ILbSHqkjQNf3E70BXh/qrpc9hd
/5te4AnCRZ8CKbWDonuIRq1yDMaFA13x9ChrMKJ7ZywaEliN9ZSqla0oxb/cHefm
z1dEWngtkDquoYF2kKbiHad+g8plmGTPPufG+Qhztia/3cmiAwZuGPPM7x0c5xpA
FA+PVCEfLlOUTA/QhGyqCqbRQ7trRcDYSg8GnawAyVnYn01Tyqmw8QZw6q2XxfpW
QpJP/V4hgKR+QX/dbC7GHD2Fl5RqHTTcHR81vLjiLWvZ0zDIpjk3C7PXdSGpzaNX
C69BxCTyB3sejYXrUKcSSH/lZxA4njz+KJvNLbhfGEMz0fhoGk50dsVSkTIwAF9J
gJfSUPzhoLr0U8Dc0WxT3CJbLlVS6bWBNSmjrjNQrjKlNpjDTxnq3u5VMjENk5PN
Fn0EZyn+Fldw6Y/i/uF3h6/fymgpBPm0l1LjmKFzNt7Wq2AkCu5Wqw7fQzWS7nn8
YanKbj/ZJ4ADeB99ZhvTmY84gpyEfWg4s5xcTCo1/PsHUh79wkHN/DpIVmknFh4U
NS/mph3esAi5sp7eFK1iN8vzsqqxLQ+PRRjmS0MN4LIrwy2WVq6lHNvjjIl48EZz
a6VWps04XAOKZdngKSzvpJqjPvYBZF0pzKrvahTaQDezcgAosaiZpOLXE1d9mCrx
fNb6IKQBoueyEIuAdCA5fovalfVv4uLIvcMoaAZNQeXo2RVuzEprIEvtT4faB0eC
/4n4tFsia0qM1o0W5vBXx/qfxfuqvyFzczN2ylYbLHnjPO8YCxWuKr//21JRdVwa
1q+4j1xryrK/zhrC0iln2Oo6oVqwyllR7pHHhztv52x4CXkYWIzd3FFvgtT8lJUk
1FjP8Gb87w+7TfCXNAOtUuRHmRDT7ylvLHFKVOlSabFUe/5JyOQ71wBogcH0Fylg
sZ9IdDe8umKk7vQRp6iQEJPdjmU72TLSm/4xqobslqsEZfu/8Bpw+hQpvxSjjixu
9fhs+toeKF/JbcaU3EAb1qG4Q79yo0sahL/3WTCuSaFp4dNHZjzCqV1SetVZOk8W
B5FWtU+f9eeDPS/wVLsPjVj+8DaDJvoTc4knj8a56qxLLf/GQWxU/i2Ce/P3nujh
uIly7ifARnvSNojtUpRn8fS89ZcqSUOB2504VXz0abMbnMmPpiJZv3K8WtofbJms
dhVi4beN3x9iSQGsuZsvnmEwQTs2e92VwSTetJL9/cz5kW7GEzWY8Cppyauke3wo
AaeL34Augq3m4b7ColmTDIx1XljXYcXJLyfOZoH6ffShsS80IXsBua1YC1Ds/Xh3
4JTD7JjdGG2mj8xJ3F6Ytk/lmaB4fqL41oVuu1r4OnxuFXNESo3zDo4i95RC84BM
Q0AY3r6PAS6Sk1Dc1Yuu8jWNP1G8Co2gvMPjYiqm8D1X738BDODI4Qbjz6qk/+OW
HqLKMZm5PtH6qlGaDcq4Zzh7EYaJataA9s9K9Wm3B03JRThsVCOYvyR0lQfMqf1y
ZADhvaddbJ/KgWiOrwo8mV7wX9o9h12EBC1OY4xD1MPnDuynnsqhy8euolbMzYZI
6qm7kI3vObE1aWdQfmdlQXbVgfKyeXmRqsbZjH+GeoGi9ul2MCDvoJ9xL4uyM7/i
BDhSWRDOcSV5Fu4IcRdX6XMtu/U35wAX6lgAbG+5HF4EMooEnexki1oRgz8OaXls
gf41U43yYC1QGQLe8fYAwhfp7pwOBg2+dGfJQ0Z2bLk9CcJNAF4pnz6bmctUb7uf
rAO+8GBiZdVcjnkYixYl1UiEImzMSQUR+D0gJLD5d7gOpmCR9nWnngzIcUQRWh90
lJmelsll16CAjniEb9lU/35m0YxRA5bnnajdk8ALby7/M1zkYgv+Ubi+yZPFy+xY
vC1FkuFEsdvfgUprVGwP9hu1ijucZxa5y0u5ALzlkahM6YtX2YKexYwZUk0mzONA
84b9iCL/EIeZqAINZBShlt/HgMfRTrB0SlEGjJPZpH10wjB4sGLpNXPCTSoFJtkJ
ECsGzTXYluSXz25Hv3QZ8ITMT9YGjNU6XvY3i8WMYU+BUHrGMzIlHopXVdvy84GN
V4iMhAjOC6L1aUcfqzGW1Jp8aRABYscSOGArNFbdNuiGdgAUlsJsZnOJiMLmQ+kr
FzK3J1R1Jv1IUVhhYOn11x/WXsY0t9PcYEw90+yC4mEwIAoh4vaSporFFBBedi5r
T1N3ptE1+S2a6zCPo7pdZJ7m12GkoGO7IsMPoXpKyR2suDob5n35GUYimf8pIY01
DkouYRKG7RkTeTJxN81agtCoME3NNe4ERW58g+KULXtJYH0PjgABK06c3YF2dFcx
7I13cWYQFahBUnpLQe6Ndj0OuEpURd4l8cBl1+Bv1nW5+trhm4XpezBsoigfGUTR
t1ndFOJ9QFHXakWAdCI6PtqZfL82PBJkyMQL/9uPdcMZdLQSYBziO31DFcYrHzhX
FGowXBIvByWgh9+LGmOkrQyw0OENVWdjq+lDWvJAxlYz+1T5EJLwKxBrCD+SzNld
J8sESCF278xYc04B9iuVIFcUbS7ft+8lk9u6c7wHWRd8Q3NI+ZjZAx448pqY2rB3
WEUzI5CInSdp4OUZIjl7Eeakbc1DtAnbH0t5ZaZdHDUv7iUSj6bLEjnLj9QSZR5I
dYJGAsSdQhoOZLWMn2lgjWSDlq4LagUNJZLyjzTGGHrkzHbwth1xx1lMskipohq/
vA0khpbuyOkf0YNVTOf6CT2nnTQLcOrWEcKpp1E6PAWZe1P4OX15he0FRmyHeceT
JojFAXaaRk9Y4wGSqPBEs8/zIOYacRdnqHn5B3kxvjzkIbSCvhfpq+z1P25mmIk/
V0edCptBXY7kHt8mfuF0vmaMlEJ6WipuCX9TsblxUC+Rdc/nweoymNKHtB/bsfd+
3LfwLlTyYacX3lekD7SraJYVpjDwnWlEXPHvYDLKsvtM6gRwrq3zc32YW6AS0yfk
PtC4DqQ6XDn+3WtssGloaVkTWM48higA8v/J5Ugege9BKB1V9X/cemzYcPHVsReu
0pLwojnEX6pwilvaDiuV11jNKAxweoOh2lgCCmWKjGAHmiWMikjBxXbdCw6WspE6
msgKi6J+ovSQiIa+A4r1MIyDuI/jaYLSN17rPOq4Rm0CI73IVPiWz9rzvg0JGEkH
1ChdlCbt7idsuWc3VLm2FfdE0lRdQkbabI7B80hyi1PV2P/jbGcu4UBKD0/rxe+v
a/qkqy9pinPulsJZJiv/P6N7PaPVu28RKe2aQXYw+LUQOdqCBH8ErVKnJfirUxZS
uLpYwjxgCELCyYfJLE7IEVaZUnxRNIk+y1S3yBV5WvlXLGmU03SV7gxqQGhu5bi8
0MC/YTXCdY0Z6FyCHyFxIAOLcu1vxXkdWkhaBOCx0fVUx8Wrsa+2jxv4liRWHv9s
fuUWyJDn3qEsKHjSioI3rYtOsy4Dt4s8k5qEZy/mPNdLMCysluA5oRTKJxdNKBGz
+PEfmg9wrZqqXEpedcj7k1V4e2w9/ktLd6FyueV/7nzkcg+06o5eX9RwLfefEKqy
c9cKoRA/pCwZZWgHNCNsqKiNw/agElpI1U0NwWj8TKNpOk35IoCU1r3mUno1gU+U
FrOudpboqHDAbpHlaYrPrCq9omPvHERA0dK9XctCXKTU/ITSmmqafOWoTY8MQQXM
pt3mAcMKsEy9VbaRj86P3kKRXdPa4P6pun/cqbstOc23PvKY8sxNfEJliNlz3Nmq
vx5cCWf41846AnsoJx8b0BWzrUtI+bExnksTxYFK+O6Bcr+AKaOPZJK8JR3SFjV1
umUAWGBEl1jisd1OCxl3SGdHiV0ClIXd9aEzERHqH+dN2dlEvuYMByP/dOYyFH/S
yd0zvlt/KYYcO3l1EyCr5u6rQQs7t2KZocbhRK9jmz9xMBp5eP7K+MksCskrvlML
foSPVfyBABiiZKNxv54pRJQz/SS2+rw3TJ79NpV4ZaJNoa+BhhtSE1BlKE/RnO6R
zQ/eSmFc87C6iqW+Ta+TM4v3bRMBZ3/bCZq313G/3rrbmSTjg2Yk61SMq9uMjlLi
xcZsJasZJpnC0S3WK4nd/f5AxJFffHF1k3TjOJYDI0rcaKxpqY2GsMX/2vaugcy3
UlIBnzjsBIobOIZZ7Wm8VzbiNN09NA/exgF2q5HYUNbW0cQcSEYsCrdd1p+lAtvF
W5luq0yktevekHqbPdEqcZDVRwzJaPgITB4g4zVq1UkAoKml8jVAQNrtVRIBHEII
dK9ttzqcl4ZDBcPa9EUphuFJCFYJLEHOUtr4tRGwVUACi8tOJ9TYjuposqdXcK4+
Y/YKbrFCbR2/7T6A8M13dXHBi4BVeDfFpOh/e1xQkoQtiAU0F7QGaDnK3LO3Yr7R
AzNnEdHUV+hFMpWFuXBH6RcgF9pXm0qKosWanEbmHBmnQjVNFZfU1m8UOaQNQmxg
cjtypp0f/etJ0QKR4/EjFypctTEBT8SeDwwU8rebw/8yk9hI+a3DNwI0XBVtHVad
WQk7iRaEmSFC6FUjIysYjkZ+h/Y/uEjN3qEthplUgwvNxKnGEATEWq9E7B2qyoJ6
bL21a2kxK9/YtocEycbJrQqNfNk6kfC/Fngqw4EPXVn9uuVrR4df5Alsce0/uT6/
Fm4p5e4JSYn6Lyjs3PZgbomBp3sF7k4dxeEelyToAH7rwSv1/YoP2QCYdUjvAVYy
MNA7iac6yo2oBTSaKDytJvTAWYzwV8EK7ckoZDTFP/39EoKAygS7upjunnbrEqfI
FxhdFCk6VGW//r/CydHpN8Safo3cIMbl3J64a3dBeW2se7Xh3ufFKtWmQRRkNr0g
sh8KjGq18Vz0ExwCp2TjZDBu2jeFcIMhcrFXe8zW2geFASLsq0/P0hT3sVvuHjjF
RHEt7zwWIkLpDR7D3l0KYd+Kx9zw3omTBWnzP3qYVi5RdGRI2eEzlL892uGNwn+v
gt2zEjq016f1RzLFCGfYZhYJe2vvFOIAwrzYNOZRb+pFip8KpeFSSclsAeqDY7p7
iediulXN4mIHOh3nybucQY8YUtanyYTmV4RHApYEihoRQbdwUvpaauI/18lz6iXa
uBLGM/91qSzvS2ZcYYSYL4Z4Zb/cfK+OVeJqcxqmhU8zYgZMJ1EV1jDMFWuqr5T1
BRL25sZPn+eJOsYlst47PC1U+U30GJN04jgKTQt3gr/YNYc+pLAqqZ8cTIve/j4M
4XZIC1G7sZOi/iMdiKqTmq98ZCTVAxckav5rD74eS2v8UXWHS7Uvx3lptSiW7bJw
r+zrrQOz1ep+o08GhM5A5jKZjyV4h2NmANgLpaw6g4qv0MUHNu9P4lirhNML0ABj
dF8VPbwo+EZhol1WjntCjWNaxCM0ybfS+RbBPmPrsM+RQ8v3aHPLVwRUgUTWMb7q
feSjQxlNkJ5gI65cQyxn5Sseq/pzdET6KVc20w0cIiq8gwYvtRypZdKNTERm8G3b
DcIjgWOZx3NrzZGE2WgwnChdGFnG95zkFU0Gm1aO/ne8sX2n1aIntEVvmn4LB6qE
DonV1J5w+qdUkK4WK0oOgftbVtpH2I3DDQ9TVDKJlEzABLY6PJvvNZuSFgc+eiH/
6Oe+hTBLJEhezI/cSD2y+r0FT0IVExH70SEMVInkFXV134cx9H4A1ljUVu/Z/yKQ
I3AmAR6DEGAG0GMthU3yFGQpSNY7tabDQA5X1EK+947K6lSqa7RKjbQNLjuyOH+Y
ywqwPf78xSTAxJr/KXI3mOoi4s1+0PIuD6pRkafvR3q7f7LknbjpKdDI+lUMbyTQ
/fGiYlzNi0D29mChHwrzz5Wmscn6dU9yG+wb6wt1TnWRqltMFRtuvOxJ3k9TGkgP
noPl3RE/7pwk3Q1OJgAAfRG9m+ixc+/sRi4HMuRk7Su6I/mzFYibB7qaLzV9crwB
ld95lgr5N7znvpWf6Sh6m8ewQg+ARCXuVyeDxqT2wuUpxo3+y4bpG9E/TJXYhunb
RZxNaKw3Ynho1P60l5giltwVIVhK+ozsQwl7tufO7chNKkTI0MEVOJBsBwIj8qE0
BnEYypsFpaZjF+txksA1GyXuyxic3wEFRj3Ymg5CwzjNwvRybWkyteJsihRPeE/5
y6c0ojcbK4i5WU13gK6FdfVH1oEIaAGo4Y8lfdkVEvDxGQFqWzzAGfvFBz0oaP3W
mC1VvH1seGTgmHF/EIM+hnv632iwkNM0Ly/8ilRYLsRG9ieDrus1RdPZEaJG24RB
t7MhQ50Vl60LL+AMlb0cGkXtPVoB9gkDrbO5M2bdgbm2puBTs0IBam3x8Aof0/zH
V06509230fiBp6mI/3K24lRYZSII8jGJCtQ4QZ1QgILz9dg8OM8Ia/f/hU/Kj/sy
/4KFWxmHOeDU86RDA6Hb4/Q3H/+LLevxGAtCXRk8kpq15TuL65BpwIuaCs6zUfB9
GLXVfU1clTQmqI/0XlLEKrFl/xg1KLiHe6oUMJHDDBzfbW1Ufa/kpdT05wTcv5i5
0GSng6NbCD14CZ1LOmHh8iUlJgua5DzE54j8nmLdsT1HZ+whqtwq02EMBqI5fg+X
8iuEx/xtvZAgRXyBf1TDYxPC31iDWdEFs/UIKzy2abT2L+4KbyuqRs8RWZycOzoy
1De0/8o73BuDsT2bA7gsBNXsX3PackmiuBJOQrXWCIdrDHH3X3E0K8Abt61NJlFH
iCa3bRnUlUcwSZsnr/5UgQ/ZD5Syzx/7K72sjZ+fPGxacTvhDo4eiJ5CxJY62eYs
WGWWhIEv6KcDRxUyGOEPFDdWFsBqfm/cjZXGoQ3BUu9cLb79Hkl509mNYiCIinlE
YuT1OaTHdxOfRpTB5iv7ZYN0VSHgzqelxtmJulOZYljcgw6dVq2acfLqK4pKYwCS
tb22P7b8XqKtjfkglRlicSE7b1uE1UY26a0EtsEFjNpl0Xnx2H8+QpcVpUfMfR2r
o+tiPCiFyy29FbpjCrXxH44QWsCaMUlsfwrYV2JS8+nwI0fh/koE81Czb1VD/hxX
cygRDkMF65KRW3T2+mynmEwvVS6zSWxP/hLBCltfRzj9l+E/YEw6ctEo/MvyPOjR
lY34038Bjag/eVr23FGg2lpeu05fmk1Bd06sjrgTAugiY1AXH0Xt+qITxUvS4rQO
PKwXuRNNCc0BvmlNMfl6CzPNc8zd4Yu0nlcpzk2A2h6DS3nkGergLSIUMZPKYgI7
gbtrpMkgOOicKZkJqN03q9mSRTewoJwmBG74yL/6J/Kr25uHPA7NQtAmrEUjIhna
ZGfEEpkG9Cz52LGO0PFs1P2lYediFfkpgBLhek83F1u3WTjeUJwm1H1DjFfXy1nm
TAdZUJONwtToyqWkSHVnRFvmnLLlPAq9hBxWDOflQhNlNi6Ie4gvIU9Xcl77Rwu1
n6mZo17DRrMhV62NYcm8pPuJjZxvnZfmOxUSa5kY5P7seWD5Cuyv7rT9Zar/7hDZ
bE06LGBlRI7CWLhQEB5ZMI+c7eIPt29KLzDO5YKrRTdKfdwdrSS+OT+VkuMIYjVx
JsT5q2mrLCkp+6nPUUkzNARxGqVWLTQPc7EELt8vLEOg2vVQoihzDTYjtKgwpqmx
/FOkQz96jiMRopySNLq92Sm55Hboi9gq+mfwB0lYLyDX+QPos4buitpYYdTpnqLw
Xfb19vXo8eN2rADdAtzFc2kwgqP09ZwKxkz6T/6Tenr7RAbUA3TCiWFiE0wbYT6g
2bc70Tgg3Kc/+pwTsT8LGfnUDy95AQ3ZHEHJBmISyTIvGN8K+/wssgifL7yLCsJw
SR1BOQ2TfLPKqU4uE+lovDKrnrWzxVc49AU1jd+p3E2cK9bNGiFGUsX4NgMSI6be
ifW9RdoTxoN+XpzwMedHWogBd9oK4BE01djCHXYlvgQ8sGPGfy0ym44K+irHjXVs
z3Y++S+rjG5lZJ/hieIsPOjVddy7fNKttzxkQ9XzNorG9zgFWmU4KuxAUrvzuckO
yLXhFA+0H2HnessVwoL5AThPzyU76JN/ZIi5aoYlD5usqHJcFb3LXGA1rOZQQeBD
nUptAS2WHTv/EhzFVVTzkbt67y44hw0cAzb8cnfhwkCZL1hfk+zXpcJOiPWZ6NsJ
/PKaOUO4ZM16PdHI4yhjnd93tMRAvRqlsEYtg7PpWjjj8SbsL7dul+dShTdvKubG
OYdeQcOSZEs+tqIfjjR6E6p1XSPIvXzqZrxI1FN6ODypu7Hj9XU52eT9cl1pP0mH
v054DXzLP3lh07A1DSusZ7QbXVoYZeFiveMVGRXgS7RPzF2cRO1OAiQzk2VQ0S3A
S3z0y5pBKNJciv2MYnv1a+5JAVax9dsygkE9oItR0OEK43Ee1cONzvLfpu+io1OB
pk90B7sJ7MTV+f5glg/Y4tzDwlD2GzRUwpZTvUEzAyKEHzeDCU721rw92J7mMFhv
L4JY+7iPhj3RFkEJmEdf8LPQ1V5cRQM6a/WzSyCz7U8nZIm9Nrznn83XEo0cRURd
NmirN6ayy3Q2x9icrscbAp18r0h4FcgdeC2agkUriNUjJf7DgtoONPNJ56QrVaeW
y2AMGj7G36OUupnxzVDsH8rymKmy26ZHPWRy6LdG0836FxnmvELjEirOK8/tPbHd
Tu3WGsF3p0mH6XuhbxuQejDyVVprYsbT0TmrWk1EjTcwA/sdE+3XyBwSjvPh5hzg
JbQx3TMa7NLbMe7qbPWSBA/RDStJDu2tGluassgfftykCpWtdIzkRd5/bpuCLciQ
NknMEnuZWy2lfQAE+CNbzx098tWG6tO+RYdEG0hi3EEwLA6kQ0WUB3fL3cT/1hwl
qkj9od9ThtysTXtdgh8iZCWBDDVAtqB6URjAM5xch8ZzgJ9SVrgR+Bdf19GVYzYw
NMdZ+jio/q6awVf1SFIWCPiluxmLrGXclsOh7Ia+ymnKif3JEyHO6wBL12c5mXSQ
jJ7stm3h9qlOZ/SOszuGSE8JSzuyLTDWEG6CmJncqWvBsrg2LEreyFimabNKZu8b
fMT6/Sb5dqvGfDYb8ilKIzlGw/1CARaa7onh/bv+l9MMkDjKE9JTeg0pPE6bleXk
mtp4bQWdXcvVIOG99QVH2lCUPMwq9LoPT+aYn04UN2zv7xugI+V4r2blzSDu7JEX
CWTDKyTiJqA1Rh46F4l3dGtyLXD6h8Ogd6gpCv9aelkhzwwO5pKb10fPWbf9Wpey
5q0r+Ioe6g1OOdZRGrvrMGzap6E+L2/hJhiBkLR1hbTsjNxoabTZr+luHGVP1Ov9
ZHFhdkKcpl+JC2+XgLBMHcXJwLUDJH+dUgk+0dejF3sWhvG0bAHzxq2fXuu5oNxW
uqeyID7nWFYRsDKxXNqY5eQ/hTnWVqd/ceDR/f/hTP2aLWoT7ye31tzVKptihkjZ
CFYETuC0lLXZyXTYVD3bX5Ecav53/PTSsAfCWoN5wGfyOmIFtOr61eWTVX1y+z70
bAozgsHVOb18UFJ6mePb6lbM540aEDsU4JGhMutSg4/TFeWozjSdcjYR85dscAcg
uuQYraLliVlHlzjTC4D/txQdpsWaSFwdpmgpnA0jY4hE4dFc2lCM+gyid5rjO30i
xfNBgYVLgR46dcdGCULpCK9v2aW01/kCyt8/M5QcxLhaEwDRkms5UhOy3SXPURqz
ogV+MkNxklXJEu+MYEG84nTU8+NehQ65hSHk0pGsWalE9je66ufsIxz5lnsSRe/W
7pdPNlJbUM6DvFxmUMIo8l+zxC+A7Mo4gI0qojDqOV6HVP0IYY0E1/ZXYyji7cMM
b+qdGsg4TYv7fqXwtBVVSCkKJvdtBj9vwrfl8ci0ItaHnRC9NcnJfFsSOEe8lyCd
+ppM6C6XZLtvSFvuPXpbfZkBV4D3IcvQObrqSXyJVJkoHsDy8ADe9n+Us1S+wIrn
6qhDz12NYGDacVh1g01QMyrSZC0z9TLT60QrHqWI/iGoCFy9LwaSIl4IDupstmEc
pumxd/5PB8kv5oJW2O3vUpjgprG+lezEDhmCeqbQTw+kzzOj/Ri+fNwcw71XNX1F
Wh0wmQ0YOYWMZI4i5+zIRgzoJoOnwvMyUZbHbX02mnMTR85S+162HrgX6D+Y3TUa
w/ZpGw1bEUM5g3UwcqKlAU0TEE76RSWpyXtBARmfrbNXgkhY/eTXKOBcjjYJE7m7
npuuy4lIDQtZoTskGwWMFQvhtghRbGBGCCFudunsL6p7cxy+k9SeXDJhMc1Cu23J
zbYS0pjs101eSIMixSsueqkBFLWyT+AGvnCr7ZUJR70sQ2Vu5o4oa+1oNwIYZKS2
YKLr6IY4tLhrCMf32PeEsTqMDNu9DxKf68ne8CKJVdBrum1Qphb6mPx/WNWSicvU
irlYg0c25kKUcCsjz7WYioqgG2tzfGlN7bjsgKF3a+zTtKoSNTFCGx8HStZh1PTb
j3N/jsj0hJ5xgoAg3kX5eSV+t0jxvnpW30HrTCJyL0ACH72vk+UpgiJ2ObZi1Q60
rPwm7Y+S0f8Xj16WVAHuOhs+bwGj1ynZmNMf23RFVK71oAkNEdbtnUpzg4K7J4uG
8/WhSBRVysqtxpwSMS7r/kesAUoTQ8TyXYd5uZp+XbHHnCymL6LouTQCfM5NoaCM
el7kTi+wB5yX4UMintdtIIZ6L1gBcfwaFOX5yTTaKPvd0RjYMaFDWaPqYCXFaci/
nt2NEV8nyNuSrheQN2DW5nXkGH16Kup7yTzsWTxfvw6ZM+t6+Iu6d2MuFVMWDI8X
NMEXPngBEZymcQKTUhlhr/y3fKcegh97bQ4yjjXCL2PDqZ3wZYPyN4EvY013y15O
YNXsSZnqosmyeLZIAaUjPpQhx+HMyP5t9y8mfu299Dk4uZi6yqoF9H9kIdksNW+l
5JjnSDFkJF8uvhDOGfPJ7qK5xKQRMTVKW40qmJ2aGHuEY0yNd8dgbFsVXmnpTZkE
Dj6U7ptm7rQ49MS8m6QUaKniwdKLY0VLb8KTb0Kiz2TZMs9GFhiHcUcfK19blTeg
edRxfKwKNrW2HUn4Zwt7WiwhIwDF9vdIaPHx+UfdF4PKgco+vyVa8uN+GFiZ2zRP
es7d3SvH94Dx985WDOLY6GyjAQRBl0/pOYCyRs8J2wqSAWz+984O8RSo8GIfKv5J
Fz1tKtIRS6yzHJO1Dyvio0jGRCnQuTbOaNnQCC/fihs58ArmlcPSkkMUkHSwIpus
YmNDFyBpLIcRtT3KIS7Qddbs2uIwtqTeEOGvY3jXBoZb5TZKmFLIPv+XJnmfd+VL
oGtFR978mSVtOwDxy1ocbn0LMNsJhJ7FxIDahhL2kVy54ir07p+VngCfGVOoOATC
i7go7nFPZihMUYlAGoGBSxfmG0qlXTU45E/Tt4tGnuOs+QTGGjcTk+k/MTqm9PLN
rfXTF8VGH9ooKf9Zb4K95kO+9/JP1Y4ds3xo4TlGeLhluvvjmpbhLUT056eN6XC8
sheoiQTJTfjnYU9JawlSgoTXlJOVF78t119/h+TpeO9EhiylnbjmlrpgJ+1szBAo
gJASq1FPKk1XvqgQwe+QYeUvpfUuuJblPib7sPx7BzDhoFLc6t7PTeHdA+KQmz4a
rN0gg5wSrURwEMmwkHftJ4ZyDrhI3Jih8rpIy+XHoW7DpAh80N1AgHD78cta7c1l
DC7/wZoj6sIMrgUbM7j63h+TiU4mwjDqCZZW1FAOrxr5PjxaDyeFNr5DS5JrFwVT
7QFJuWAY/ZrUwbLtN4msoi1ZkDv/4s2vZ9+/i7LCmMjYzcrwveyAsKWlPaAYyhMe
RcCLg8BBXID+lDHHUrtYp6+VJS1jjcVm5gtbloalyh+/+4Rh3nXgMw9lhUCMqR0W
onNBqidHRjNjmK2aKT6E12w9IUa1yBjdPFoK1mhiENghjW6A9xFvZu95tXzrQIKq
KqEm+D0f12MC3vGTbubWbXfBR2Ibrhw1ibLMVA4snIs0qyjPNT2e9eQLSlptaBG+
OVfGVobosCXUJgb6xD4hqPwHUde8spQStsDMGlOUtP6U374vSLZymWZGOpHHZgb8
Qh72QsWdCG7LWkBwrYF8if3g+hE2d8lYbkMZA0NPvo0v62JCLOfGGYAehikimPvl
nZumRdEDxzveSpGuYawbqVLqZQLRygLuod1tXkhdkS3+XxLxE+5OWd1NjBSnnj++
7+gAf40sxCe/GJgEHGoCvkHCkEV86kr8rt0XleGzTRtgtI3pVCB6uU3fMJGyQd2x
VT3zvxnwft511JqU6gwF2V90hg6ccKYVQEcwghAG2RU12L1OJA0qUEUQz/6LeVAP
DdLbDZ8W2i8hPy9prbDllRZ14yVwkh+oEh+0YDFalTMSR9ABwNoxq+KKuYd2zeFM
j/txsB3y/VEHW4slab8Dowb7sP+pq8lS4tMFLkrp1a+Dm9zwMc6+2VnwJMVY1bTz
jD5VmJuNO/nKQp2YWDlushmAtuxZtQbJlDJonnwWzrmQo9wrfB5BEZP3VLF36cjn
VwXQXrF9GytxpDq7vDSY8GQd9jKxdngMS7eA1M25jZk7uapBaaJTRK4swi63WVfs
L3XxK+ZBCcj6uQRrYAvovY/1fiyL2fz9h/BB+orLiuSqMbZsFaKYVR7Vnp88iAAO
uoF3XZyAylFdVX+Nv3rQsuYzYoJnA0dYVUg8t2O719x9GrOxTnmb4T0o15gAMOhz
jetz0hxl6eqDxCxTWwbwyKf9YepkJBEFsiDIMcz+je+5Riabbbd+RLprIY6xXVFM
8/yRYAUrveDHkvPzuhI14y4lruSsc1R53Cycxg/1xxmFw14RBi3OvY7pJgRNDHZk
2BLK62E+NRmK+/MWt4YZUV+gMXSfsegrhYC0oHUNCP9X8/PFr9NiyniG7iybz6xw
UQwlMpZxncYhzyITciOpfewcaPkgub//Awd/DxYhmXiLhT+tSrAFXWMdTWsLFq9r
ltfSR4jhx7/Q8BM+TPz/wbnJsrGtKc/tIgvKTTW/DHrzevkLznTHCBeXX5Mtc6OI
U6iqJ3VP8z4avUq/S1bmq6Vw5EWEtXw12F+c+P7kU76guMSvn3X/sXEhWdHfIGSO
4fEQtryABxfiA0kIHlax7kInfWMClZXMBXOanOCiBTxyPqP0YpiOcvoLf2I/DLm4
a/sZDS8Q/O1+Fc1v18GZrmw0BB/d9b/rMSNpHCWEGBGf57yhLYvEHCqW87gwaSWj
yBMmRxUXO1FBDLqTs8nMad3TgJnivW9bblDnZUI6mfsGE75RZFId79OWTLSQjuEF
c4EJVkRaMQvIX3MqnlCLFNUAAqdvtik7JZPHH8LnbQg9og/UoF3CNmjzkifzG4HF
6wLuQVQeb+xR0XS690bm07p4G6J92OSogONubvT3OD4zj2SzQ2Kf/BSO0vVeg0dE
HisGnEc62713L/nk1n3DIfejU9Lwcq9+WHz4oPFLxSP6nRCxaopaFAon+AW0yGtR
/DEM2iVZJoI9Yo1DpLhJUKzyPUt2t680NlQqIWStqZo7OmF2MCwEM2sQHoWXt1Zm
SRlXY7qXVbimAonc3AItZguVM/KlqXFDFKquUaw6Vfw8gkXBPgViO4Y49WcTvEoL
CuqcH66cnecCcbX9voT/JgoNVutD72qI0mpngIO4Z0K9a0cqUffl22hp9TOnPN9d
mz1LXIXlOR6P9pu3/PdVKOPiU2LdZn6vOZuWR3Ge/ZmVayYcwh7+liTFgyCoRahl
jrrCTpSYCinqlE+yE0f6YCsZeECV+r4Hd+pyffW4KEg2UsmAXFHQg401imRIPBaj
5zKDRj2Pkmavsh5LxA8CbjdCAyQJQT4HV+Yta/VJHbPLJ5KX0pUNzuVIv4BhjYNF
QUEx2aP+voY9yA7hK0JxIgH6Z3Bx4HhA4LEUVxlBfEQ9BGdDiUKmF7yU7Mi4yifW
Om2er+MWC0fCj7R3us4cQIZU7l+yxx9bMImrL6wUQNO5bK8NuoCPykk0uOOTk7Nj
i83cIoEdcQ/xbyS3cmBMDc1zgJKZAaV+sYoLq5m2FeFgWfAm6Lh0Ht+eYFG1e22l
AaQuc0/QEDGi22Ybtdsju22jq3XARVbNub76HBDEa0WKJu/BBKxprkXc1oYhnMmW
DQohcKuF8HlGqhGSiQ3y0/mt8rEjAktmfzwqX5BN81gWXXA6RFpLD5JaDFCklAOL
tdC93kwLG992KjpmJ0j0mhBUCBpVOQeGAF/ua/7JbrtgMwAVu4dqHzXYYBOwgCHA
FACJ3MP2ZeV5tiipLOu/4sn+82+0XRXsjC10h8OamoR1UdDYBQ9KXwSNvEP7KuYz
HHVeKSGvvNFisFLkknfnLFo2R0dk+u2XU701IURmrI4h0au+7KNdKSRlTq8NuHpb
u3GsEnCcDlhEuM0d25IMaMTTkv2AfTQRlBZXrMMEeoMwtXxDG/0iYximK/xhPgBu
UlomoF7WwENEX7JO+MOUjl76kM9enUhElcbZkxtXdh5s4aAD2to4FMfiqSD/kWtf
c3Gu1jCoRWsTf77/CN4ZLE5QKvPcL7yO1D1vLdvwjxJbYDWFr7WgUhzQ/B6kmKGN
W4MXj0AFCi0ymfLibVuZawvGUFfjefZgfYOvy15ctTUuqCa5gIPzo2KeGzVi/Fu9
R82If2jhVRKZ/4je2JbI2uYWNMc3U/XmYJFy5HSV+32dCpNkFP2GK6n7lhCAWjzV
DhBILRrTrBaQjPYmsBoaGlNsLONIggcHSFX6U/2mslZKSXChHpILRJv9i9PsFnNa
NkqovaUKJUZw4Ua/5GQgNaZB73rIPYN6nsTkdIvmYplg23pi8wHiAuY/eRVnTAWy
r+iEbMNKTcOcgyRAoaascLWJKGEeNsGobQ++majnJeBKXZWTGbpmFgc2NX4CsIBh
hU0LJ9HHZp/xZUrNHktNSdEM5DWIHu+qkjtSkrralOD7nLaWtwFQlH32ln4FhENY
vRlaD9dHEkpBHOGUPip0HbB0W9ONmJfV4p0II1C+Nm2Db48n1eXCCZ3TeNWOZTNh
/PsKPVHoO3WPsMO63r1UPgY5VsmrBXt9Ikl7Y5yAdMSPzLbNpXWi2XMY67mQKnUj
7cRHhoScEnqVbyRyf+W0oygXNrNfLijtTnXeqMP7Mz7jQxwUfD8t7G4LpNAkGggi
Z0Srryog5RY8xt8f9dWWkB2YzpWIuhqBQWlqsebu8fiCyzBMbmSlrA+ahKeBS1pW
DUMml6IaiQW8pr6CAeO0Jo2jOfIbFgTc1X4eyal50Xlq5XzNJft9qPUVssgMx52q
Zdp4kU5mT+IuQD/5FBpSutpfOc2w65JM6wfkv54LWxsCscbZcCleFFo9ccV4IGUE
/G1BfyHUQhKHVuG1bmlSiTsOkp0WitugjM0jkD1JsxiCcDqQ8QhyiDvnZqq18FIn
ehOaMlDH9a2+lpXiMZeWB7SjUa6SXV++FZ4jY0cJwAPKMFkAq8a8SC5/y0eGIyz+
eGScyG/POkq0Y/BbahhtOVBX5y+8QjH7ZZCUL2/RqDq9xmxiBjT3xuzwqXsYWpF/
bZJpTAE2LQrXNneTutxLrNWjal+FFd1ZOcGuyv5CK0XOBRQ9WRxHnkJpU0Bz70mt
Tqtin65AqNrrchlCLnY2RuGW4NtoCP6Vng0WLaNDus1sK9gtXV9r3eBb4pawPRrq
EhllZrXCfC7WjXRNFd4bORPxJeDJSgQou649wr7j5HXkE/hxmbL6b7UC/P3bEbyZ
lp3nnNEgtFmyW1shF4eCBJGMeBk8NmDFv4UWfBY1xDz8hxal2GlTi6Q+ICSZZPqz
1gH06kznZZvCFpdA9PZlYDlhY8vXXggIxc7LbV6PJxxS3y72bwkiKj+QWRzVDAHZ
X294cMBvFS2YF6YCRQ2OkEA4FinX/RUMGPEDm5gLrgktplBBTAYh5giKw+7TpNqw
3v7uLEwTMdusKqCfrQmjXJ/BGpe1XAozfbcx8ATNl276aqv5RXkEwkE6nkgzspt3
t3LccflMaELpRXtvATKMTrTQNtIdwdsMgu12ElGl5jJI+9JrjPYK5z3GYz3wxxNd
bNbZ6elZXt1Cbl4MpaxIqG1MHgqjJDXFV6Fpa8SNla4znVekypseeYF/5LVnJ5Wt
ToVoR4qMPDprnPITHe/7qLW5RccLD7O1BNHo+d5svdNLSq7Jz/WXBEdS87Mc3BRF
z34VGCfqFvHa+DBCNVNs7ottII0TAVUz50YfzTltSH/w8/zplq8Jxq7MzitrQMlL
+GkrToU8fgYz0Y+2Y6hN9bkduFt5QagOC5q08K4RFVgW+oVtR/yOQLueHfLx/22v
nhwzkP2IXSachaf4tF88b0oRNT4bSSUPDPlkbqfpP9R+yW2aj2B3DGS54J5vwiu5
TQaXUFx3OsmcgZj4CZGgKBeu8+gux9XL27owKVDajq23h8zqdtMbgTRYx0b7dhwr
ANF7PhXPceUnjVGrkvpL3t8ycfRwOfw/yuKJX73ccxoLoh097ua2OTXRPBs2q8mT
pXN5aY7x5eFgt4+WnyehmPLnLkxOWLKi+zQqSsT0hPysgTxM1JXl/Pi6DqyqHxrS
e87AzjBC3BtRrk6Od+GTVgmoTBcAPXSXqM1/ANA8xLjGvhGnBr6gmB6WA64n38Zm
t3aSz+tqXnWUNoQW/WlmGRdWilyp+owrdVlTq7IXbuiUgeriXCz6ssvJ6ZiASuJw
5Yxb6QprpaHeMkbvhQ31Egp32r7z2N7qWNmRAN9UA4eWQn9qZ1Nf7wIQ9B9qRlEo
Hf98aOZUcEUCwVt2EXCwsamIgDjUcixc0QgrdbRHY8QyAnTosOIlqcdTHlsJ4wNV
p8bbwFTjxcB5o80zbTV4W8l1MFMH84jllpWugtoFSsfp2zJkefCJfjc0ENZqBlom
JvEPRPwnjOBd+6MmQ0SnnHx3/jPNXQu7WfNe/Bz7VLgw2kIDNwfntHk1/ncUiDUl
qzqDGKZc59uZefDnrPUv1zqquZbDJ693oxdX9QYh9zKBtmbGApvT+jsMSKanjWjG
vjaS9k25+GwmbXOAdHfLonX08jV1vvBXurk+bRFpePBSu8tPOA1ZZG++VZ8HxkoY
+XIRUAs5zvXZvRXPhUgVQuQ3I9HWEHoXjr3/fSs9pZj5QzYsfKu2AqrwyHvoRDxh
lbeE+ARZs5LQKCFU/LQVURx3TcszjwYzluF7UufkGG/qdyECaxIKwQzJauduwBmJ
sQrkmpgQFtkSCDgoP7iBDi80zl4CgmoAucer8os+IJoAWZRBsFmndqwcfi71vzZw
wFkKPdS0plwIrFiHyyTJYGWqgLcJP0cfCICL2b8LYrYPXZL//UFKo69S6M+cqXjt
kWDLP+cNojl9tprEH77ojruCEuPnIBFdBw9Swp8SHwdcOcf9uUWLB2Q42o4U5Ov3
PSTgOcsiEt/J6GLCPE50TXy5CHmqNFqi5MAVP9RMI/ACM7gZ1HdOd0puktNJiGib
uobDMEJzExcaEDJBermW9svYX11ffXwGcIO2knaEmFUJO9yO5iQbyIfmg4tBFtfc
MszKah0ftZJHsjCXckU3Y8Fu2bEGjeHSDu+zJoVQab8Dm0ZgrV8LNC9Hof88hPGo
MFczD5fOM/VKe3tD3E5BWPteeK6jHK0NaMrzCrOFI3bIxHgJylt5PRCHU1YqQfhq
2W3A09E7j0tLyFUwvQuEtIfyUOJGLz98cyc+wbqLao4sQkH+Tkp5Q3ObhyKhdYJv
j6+wwi/7nw71yf8z1ag46KrGdyqACVfR8AT8dmITWjXUSDpEF/LZNjdcQfWH544b
XjftV5TMwP4YHF7woPOZsu731iZUdcirNWIVH1VB/BO0TWy3U4zK/mB1uMSV0GqB
UuiUBkWkNv2D2zHap8/tz/4BV1x4l18H7fVARp7bW0zI3FzBYMAr/2mfpZgThzF8
7bqFuUMsIsD+KbJruw/zhPPQD0jScpf0MDfr4szU2hT98vk7VGiqq7cR+NrAhd/6
RO6yj+NvyQm9djwWWtGYi8uG26wMjMl2t+mGgyHe+CQE16VRsCDRzVT49k+e9YlM
JdvM99S64TpurSL5d3OldExXs5eDiYRwlDx8Jc19i8n2RuQq20zOLlhJYGJ4ofd7
Yg6UdhqCHPtpp9mI2pF2JZ0NQ3vNB5FBjtr5pgEO1ItiWs7LE93RJqLMFi2fscsx
DGq/PQsXPZzbSDmn4urBxYmenogGgyHlmNUWKFDVX8UbwDiAe/kYrIfdKUpMcuJa
grQKauO/u0VOlfG7Z8joMrTm9CrmJELWQY+8trunfj/hgi51/eXp6cS5utFk/k6Y
cZUbV+debBNGzQZgwELr6V+m06Xuy1J66rWAXbmdcvivuhfsWx/fPcuRynwHMrqx
Xl6p8AkhD3wJs6jNnMiTcLxV8DS/F0myyb5+AJ/Hfym1lWC5NBcTrgUUy0C4gErX
pnjjg4JXPZpBmHQmzNfeSJ+9WsuEDMB1VK3ucPuoTqMRkgxKmkoA6gCmWeAwkwbq
eecHvpwrIiAXhLRfkk0wN2HOV+FKLcgJx+xXAR4UVX3ND5V05SSIdZ5137Eb2YCO
IWnNZluxvT11M4I04H8PVf9e9kZBsFHm0tWcwmW+IN5KKlxaDXuQPnk81jvQf2iP
qUElowwH3dI2h9gudiUveIHMRdStUBM0sVWpYFOOhO+FhnTU2LDJ85zjVMlgsYMz
y8haSYFza8NHNxGPCqcRaaD/aEABRjwTRHz9E0b2QwSZGZ+OakGic1G6e2tlZzao
yuW8fvGy345ZGGWPoq5GomftZGmVy3EnTA3v5QEkkkO9MRI+kKxN8+pKrpZXnA3D
nqhTbR+kCRFTHLUb4AIejKCueVoyze/zCbwoBFlmx7HBnE6Bl+VzuNeevCxTfUuD
JbQ7yJyHM6kojm2lHLTzKZ9TTMW0OECSvy3cWUfeGoclVtY0YyfUbUUsxw+uJ7Q2
fim8K1CKmRz8ilKUT8SUcl4OtJc303xRTINomyhkyYtqjAE5GH+T/MVfszugYUJi
vhuUIaYGMWQjXM4rTbo/eSF/AOVLJrbGTjdbjumzYdkQRgiu65gosK5GrY59XJwi
hdFEiZqp+MOUMNsHDd9q8NfBGPy6KnbYL6+kFnGslRPiuUg30d2+4eOf0EiLPUox
/m9NNLbavm0KIHUpRrp+wNE8fbMKi1/ZDi5KF1sdZHkFZkbQOQEmuH9VKpaFIxzT
oprFfyfqIEpNxXPL8RIPAUfF1mmoEfItxvzhw+nGgTiersIMO4U6i0OW/tB1U/yC
q+t5U1oWYpMrefhpPUuazFnjFwspkbUxYEjKakpx8EZ1Rwdb/RFPHCAhVqgYyuO/
CXWp1a+Qqe7CgIR5Iq5r5+eSOxKLUVcDxXi1q1MHeoUp/lwDNSqAgA3CLEGf8gge
5O8jSCmHVbNUlhM6eRTJ/YzpAoNO7C5AXH6TKgOpPlAtzAc6Y5i5yCEsi60ivbl5
6rua8QxjOWL5OMQlchcKjvWTE9UmUVlV2QhEcyYSDcP/4DhLtqEWKTwXwf/KJa2B
5uEsITPK+nKXI9S9so3WYwnYVemxpQfLSN0vFzJlU9aESYY0Z0XdSxpajY80nvgY
psoVhvEelXpMpzv58xuMoTiL3sOnQZ9XXA36Ej+llhrAyQN9jk2VFNccLu+zSZkP
xbQY2eOrktmTUZ+TlpyEV5mXeSa/Bi0Lq/0QTKgwaAi527x3GlNsxfODrNph1c5z
xDtAjqs164bJlWPxpDAreIncMujL+qQTUx4/sv6/oUL8ebnZXU5B/sMmofoRo4pl
2H3qkIGxlsyBbl3l9GK3VlFK1ZOTjQOj6Ko3gcEaBcIliyMn72KHQ3F6EYTi3fIF
JIZuwsp2nNXGXDms8aPE036Fbm7ZGpymIt208p5i4EdP5lGKj4R5cpzK3C8aLp5W
38c9Vdo3l7+TdcTFobndoQrSpN0arAOylz4g6gUGSHDPnec1AiOqXa4Ze6fYM4xF
ihJo/g5J119ByP5dUztlHZ1Vx9ApxcKsNfuAScZX5PcBwDfvfOReO+rME91BWFN/
EfILlbXUE3KdeKWl6mqXoufRtpWbIJaj48OXXW5m+KN2a/cuirJFW5tyzmqsBBVD
RcJyoPGdMm4/amf/It/GujBASpIo8ssA22bfRmuAS8ojufhcHsJhwQ/p/nquLzg6
2k3ehXPxiS7rCOa/jpz/GCsYKgJZZBP5FxTA6gZydIqjgP3PbV+5l0AxXjhWqVSB
B8/u5NHzeib0sHLpQsuIxmT0NoORklHqQ6irWL9LAU5esMaoxaCx5krRgT77M5iH
pvWfnBGIY0reF1vGs+FB7c7M+f5PFhorfFCa8Lmj6W2NdSYVNZOow/SkQsHEhbJe
EjfaFbUp+g68eNrY0t8G4ElkhWyXSjX+AYzmismb0JgxkvrId9SF9k/fwy06Fzo6
XMM9z6jfUxNvyOEc1WLLqZ0OIVFZlub3HGgd19ecFwsw8CPBG7CQKpTbDUCvVFja
E68h+3DV0AuRvP7a4atFD8+MKsMS95dB9vxZG6Ph1YnMls4XUwnqUvq7pcCPr1Wt
/elDU+miUgRTZunUMmVOSjXwM8oi9GbWj+TgfxT82jcq/SmJELME7H1LmV2Izpeb
DLUIABQOuIhOKp5ZQOKleNRer3OvrwVJ5zU/xCHG0X8oa0+1zaRNMZWU/EP/ca1A
P7cHoyF0S+zSBstsOVO7mf+RH+ytXLr0ipa0p4qtwU0lD9rJrQiZRuZyjiBaCTFy
l3U5Vc9z9KEN+oiiH08J88qs64DwFOXrICiLpIeahO5JtRLc85v2B7WFOXisNFL8
Qv8ceoQ+7Vk20EGdPZ4verRKitPTysa0Dyr/SeoRiUJ8w0LQCuNvQveBXKWSPaqJ
cwRvLrU6ufDJVPclxDuwM0NapKgQPFEATiW9iOxtZmxsLZqk6+0agbmzVuL9Rxb+
XE4J3Jw+J1cVPtTlszjTGcGrWyvex6/fzp298TPdAggLE+KjKZjqrBfXmQXJEqI3
8kC9HVpthWjirzP5LcTjqX5kIXnlYF/O0LapojnYFh0o+IR6NtnEVvnaEvpV2tz0
sxxhj6cEULOcqYAmDrs/Z8iO4JYu454b0xJHQalc+8VPxJ1FzYHPmeAHLtKxdlpp
gFziBS43MJpHyX68FeZc38/x+d+qmzLC/24YIBGEUXzWH2FTgAHSsDUms4s7bG/o
sKmIs+GJ7oGmnOS01b907u9lFogB/w00H4CofFhAcKQkwsjpN31sIRQ+NzwlNQSz
uSPCIEXqGmnvEcG15yZLw8qzJ0+x7NlocAce/0R+RlIGe8vrHiT4ZZQVoRDb7kh2
DsjteGyWg9bnWBxoAnxCKLPbqIaeolnvlGhrCTHJzWGByklnmSKykn8XGNJVnFw+
8GKkFxk77og2rmX+e0z6LsraqL65BR6IZuQwbbB7ZbZGlI+veavanfe6AJKC63bb
DHyCJCJRSWOmRVzxmP4ppqXJ4Fdb/fHJFeK6NoU6Cun/AlGcJvzwRsOZ8686v2Rz
QQiSIBx/dvhpOHTcsWohzMz0HUYLLyS0ANkHQ58bJizP9QqS9Jd/SiE5LnypMsaM
zwlxqfr3HcMIHmP3MOEnU1RO/bCnaDdtouwUNXrgRijBlvoguZYY46AdfZRvLj4y
2YcgbJSKSLGDnw5imBIhC2vdWIqN/+Kn5jQ3rX1QVptuOPhKOu1jHuLwbabN+3Gz
EZGAM0Ar+UCUCnbDYPAcV4UhVVM9pKOW9MpiEu/ahLNo+Xa2hdnz3RdrzrwlcZKG
XGbnZiXEaIyd4DhL6IDdtoF6uebFP9SrGj3XhiVg5Q7VXDm5g9mpIkqfY9dWyqZq
4VeN1eBmrbxu3HdZacybX318I+VBLMIimX5MFFiRxE/yUgHsWlaNumobNYZdGKGc
ObCgr6NhG3wuMp/BMMCy6L2k98Edv7sfT75oszhsTewkdNL+Yizh1PsLm+Sfw2Zu
keqrHYLi60RhJEF34lUOTkCQknZiHOaWxOfPeF6xHs5t5xN6V5qehcwuh+n75iSc
hIe6ULnXOmKEdwFpbZdlMDXe5DwI6WjASxzdiz7JO7BUTfPcVf8/XoSfYG92AcR6
9nPJVkkaYyjKLFdYqFw6GolEvCx/mdnf7ny2T5+zT60lnR9dQZo/EbEZTP7lNh6Z
dHmzWBuEZj3qEBGKGS55x2vA7hWYcrhief3UTYXL3H9fuJZkVEWDeDixyRoEoUfx
pY1Hiyx7B0eVVu+oyR6Uq5ferJlkm/cf3Y/mpMl7k1XpzFXJxh1ku2ffZQsJnNOW
ED+CpNhLIrJFc414E0xRnSLgDe4I/9fvCcmkCKrbM0k3ZWJV6lO6GMdWshrEjwWY
+/uj8xGHI2OYjnMnMAv6WEfrHjiU8LX/n4t4VMQ1y7xwHxMioHxMrvigW4JznZEG
XiVTfmdKcCEKWHhO3bI0NdrW/FCvQL32IUR2XLKcPLATUEZKm5+Txv6mlLwLBQNI
ACaG8+R7mqY9XIP/RG73/LXYNUEh9W20s9TdCB3Z/i+YbAcIkoSU2RjG3XlcL2Ep
/dmxbZ2SCJlU2MFFA5MOmZCI1/hoLEZyDccZVDywpYF98hYjWVl0lYCwdMq+SpZA
F5YRwE8VvigwA2Sw0286qq+67Deo1aRkhEI5faqQqrjiN9c/J8plDkJ6lnp8uVLA
1fHOtnT5HQY7lp/mK5qJ35DdKBcWt2r4jctKtOR48khOGWyQKOz7+0+xO6KrxRoi
u34G7ld9qQpaAdMkFukFrZDOfTOuM0GfnxBU+fP6t+M4nnwsDg4PdhObd6JpeU2f
W5c+fcTCL+ntErs1uKVJkNICRPADXIK7gniCObwcAK1DDSVduQIyLw3Qtv3NFa+5
uhrwrILyxHqa3SMKcoC57SCGY4qa4BJpVft3NxvxDmrxkaQabQzyLIlP5ViY0qGF
6Wpkvwm693Os50yC8CNXrj8I+T+w+zofUCe/viK2YP32bEZcVdUMyvYvRe8+XWBk
PqMmVp36gBzf5A1QdGvhNnfvu81idIFKcajZwu0pym2yT1LpbCe7ZWgKz5lYfKr5
L6QIFUO45HXZdK8RKs/zWoHa6faC9mrfJBaYsg1/Zp2xltVA2+3l5qiYIsB5SWg5
JdKiA+/FLmroRsgPsrT1b5TsasbwmAGZGVApAjnL/DaVMcn2vfClAWg+mvTDCXvl
ZxYpIriuIvYV9OAMs7XkbKYs+R0Dq2tZLUCZ66Bek0A/QTjkAMdMP87n8D6QsUQi
69epE/LFBV4wc8PlCkXiZkKq9kL7MLK1VcBaCVfrQrm8cs0q0ThazERYdROHcxZ4
OGu+8eZXTblZ4U3yDAG0lYZKcZXkBkclFWJTB7dbC343cPNa7EB/4XwDMEdT8l7W
G8CuShiNHyEwDYM9pSDfPKJ2zXtfrGhj2ka8X85RH7fnTxGBJzzBqoL95ADoxg62
eaA4nXzABN9aQyZrIugEckNJ33vXhdh2DD6fccGWm92wuU9S5rvrMFj3fvw4qI2q
vXVr0dq84klGyxBk0ijSlZjVJFbfaAb8vcGBJDMAzI7T5Der0+m5Cqd1MRBOwUIK
wANBj8gIoeLKHjEPpZlF80uOyX0org27yi3/bGpjnLodb84VwWolR7VRot2U5VHA
qhjUmJg1F3+W+R07rNa+7FweVMAOlhSJoMj9FXG0TlGhFaXXkh8I4ILTTC68wmDi
puN4FEd6lc2t7j+RWIXY9dk3+0Ac6XiTOsxXLqHUi2dpl1mcg6zQREw/j8TulIK6
53g9aL/aTfJDWB4gU3+3nIRCkDvcwEarOnVXsnxbIvuYDcxmrEQtBAP0p+pgxLri
Xu2s5n9XxpJCQ38uiC0AnkSTvGPX12k1eRX6MNxwIMUWgzzWWKqa9ZJKr87pOwDV
wJCTOzg5UmQnvO3dtKDUN6Dr7tUJ6MhOIPHjvzm140ai9//mNaoSxgtCX0Pzu0hb
pMOie7YWWxb1VzA6N4m54QKxSfQMZr8BigUjYPD97Z1MSsvKfANPYZ56ZqzN+W78
JObVyuF9EcKD0Xa+cbH9haqJxWircFk8dCPvC8CAiiE/tUrdygm7ioPM/HtfHqr+
uSmPUMNDwXxD4NDoPKMoP9UiCFBV+xtiZmn70aHUSbeuJf8NXFQ7UvnMoCyGqnyf
n5XRK1NCPpa30vxUazeUHn1/de1FtUsoCnfxO3C+I5HWP4Zq/986+RQlNz9J9Ly3
ifEqt2/rLaiduwE446FpBoOh4RjqGhQHzgEYqsp2gr2Yy9lUTWWvzid6nUUMgudS
Iqq0edwDdnlzkyJA/1XKG5xK2URDWQRizTN+ct+ZZLaiD9Gv3HWEKYChQVK4HM6t
50fl83/LmbxRuDQKCwMM8f7jc3GBV6noq6t9VPMElzp1rjdMfVpChE6g0TahDyzb
oPmLR5GHwxORnl9R9U9GDnF8hfHqZdJtM8LYm8x/JgrWqhawpvX4kOd3vfxoPzD5
T/2+n4RddIvfykKHFGAGMPMT8vZI1WA9AwPjASKSnnFxyyNEelbhQgdclwY1Q4kz
T9z8iEJpO0SOaBf+uRJNPobUfGrfIptxWDoiX47rbJviPi2M+3igM96hR/ynJ/s1
6xgu/0D7UIVxMaQB8L7QkN78wivdlifsrbvDTnFSwP93C1M9jZ+Edupd/wmrxLPA
1E+yEprG66Kn5dW9QcyNniKfGiAYPLCmQQjok81lUGxwebQZt2whs9kZAE42X2df
v6Ar094/ie7PTCJlwUPQHy+1wEj9/P4p5g6zBGp733UvzVPGw3jD2GwzIDCFamM6
asw7oTVcgca7cE7ROPIkIDmPQc9RqYx9GUDvuaPGXSA+mRL2rihlGpm1yujinSG6
z29DP1ayIi9HJlJD2b0ndE3laUyD5DiNG+BnCc9HCZpQdENaLJBiXja9iFisyspY
pvSoagCXjuQx5YlRr1gvS9KJop37eNmsPaWaY0isK5nznwK8eGIGRc7ZzAbUBOIJ
cnYNOk+1Sw1AOkUVIrPid7oh/UbiwQnoIlMnwIX0An7GDhLdGE++Ztj9OS5IBz6z
erkpMJZv7D1ie+o5lyF2+XJjuX8hR8b8xAk092bx5OoUzjFz5nHtOfaVnbmi841u
fiBrvEN3dMZebqa1AokHgkt2OgDa23WB9/9KlyqvmDSVOqURuFrOtdb7T3wsuOTU
8Ln2oZE390gj5w/0ibiZJxnAb3iRdKOceqpZSA5K3ibEbZDkPmtKtOCXBXL0ghFM
2mUccOkGhdzMxJWKBhWTJDkBJ3iuRVUVdf1UPs08sxG8Xs5OXHudN30DZphJ6Kds
DcL4VP/NFqLqStiDl5433jbSVnlZxooAY37ATP+do4sRdxk/MkpcnMfArYYQMr3W
2Xke22sBhIluugacOeYisIauxXRUTSD4aGt//Rxmbyw2e6aehEPgwwGOfGqrkOb+
vR7QTT/vKpcS7QkKNA0ap5NrxQ6Dz4jVnB/KyGSkHR6HLM9EXRqxSuXumbJ0Czez
tk9drIh4BCX7SgUjyH47fZw7RlllmjapNPpUxDKxwFcW3rYcT8B+tUJ+5jAz6biZ
HQ1Hz9aMJqPMtFr5l0wwW9uEtlTzcIDuO8XKujG8H13lLUkz1kJSAH5yJozWn4jA
ReMb5W0EwKxU38A7p5yxac48KwJtxN6w4Ae+AGVnFVMAOfVFuH8/8/V6gy/NFiVZ
TmmX037aTg6waYF4AI1ax8x5EupRM1N4sXxgioVKzOYxPURMTFgOEs0BXxJeh7/1
TnH+wO/noViEGrWkV8LxAiBB14pAnaxmg8XG8QQ5+a1/+hwN/T+WwuHLUQ8DJsdY
p0oKqc9CNo0An/qu2adpKDUDs+xbatQnAhMgayPGBO75ICds/f3N3s0tam2faKqn
jIvZNGOR3y6PGhaDKq7z/Ge7ajo2oevIbkLVo52Cz5xoX2DyLMGHnONPkNkOSw7J
iRoFpgfExH/BiOklo+7EGRIMKs/TXbnrj80XxQ9wbKQCv+5/vnnBAG00UScKISvh
J4EQToYUQmV/bOBwTqRq7AKiBYXiFy/ahbOu0fyIDqRXSVoIN5fr7L9SHDp/iKQG
5B/v9DrQMP4lXa9we5hDrOV+5aU8feNXEjlMkvVSZRDiZljC9d5znDD7l6DNKCa/
PYd46lhx04dLMweg5RJl3ARqhLSFIaXRJlUqrbrHorW8ndKoNKor/GEIACixZnYk
OhpEHgUFCIYiTSuIuXYLonpA3DjoGr7n5ChJVyDfh1SV5C+ugXGvLYskjJJe/ovD
59VZ9f798XCEqWsHIA9t/1Pws+Of/mXrfn3sk8hCUBk0b3Mh/HIZo/FQ8uGFpLMf
Ff0GI5K4io3GHv9AIId07obJAT8q+OsQcx9qPi8kq/tZ+yPcmUrCYFUFecgwjnlM
we1MQmeW6KPoaitunGDIQGHXjt0pNv0XieYmDiTgU1dvRv2fWKAHR/ZiVDvch82/
GQm9MgSfms8lpifJxcfG0PfhunuJo9NFgIq5x+YeDiPZv4J3Hhk7pTRPfefd/bpV
ihCV2c0165TN9cLjITEnwFAGegxPdTEYUSm5AOK4DpJ2XfcjSIofw828Z8eVp+bI
yynCYL45W0Njs0h3EVGLZQpPpqawzDPv4PexjzutF7z/SFfqO9qXHOTvXTqbOmQw
myDbLssIZnEE09lSEAypi8OHSEC/qZ5UuDBSlc6fxPNRccEBPxlzW/iWNHxlDKEA
E5cTh/Y9tMhbpfdx+XDGGSpIw5YD1cxnbucuhp7M0tbOQ2wz6XQY+bY6Ug6FNnJG
tZ7uYAxRVxmZAc0XWujDl71dKBlKK8PkQDIkNyunw3khBFpS0R0tjoEU3clx2wJv
qIxr2iKngOGz4lHYSnilU0qTaBIMACc2AuJloJvqpKqZCmeHQdiV30sAOlkzBkT0
2Dndd1g/ca3K/5wEQGEsxyuz2Fp9MeZn5DEBMJNKXZkeAYU5PT8j5e9RnNf8eUIM
ILM+0yrgqqYCnuKOwfZLJZ3LMsILzLfXS+VcYsNL8LF1AQ4z2EHBh+/i7q4W5PDl
aLd/4vn1GPb1Qqq8PScE7k6ko2vNyntb2Gbth9A0+g5HjclI3ACc9uwg6R2f/Lmc
iEEeA1u9lZ60wzCk0qfvqUcI1em3O4vYdYOkir5N96LKCUtjjr6HlC4WnFiGOovR
MtrXX05gdtW7OoSnx9OtWfgJkjKvXBCreKkS7vfCG6QaMfchXp2eYleVccTwpmUf
XFAD6cwRqqL4G1nGnEjey6Ti0V5BAFwnj7f0Zj604gskX76w1elZmW6RgHGc05IV
3kPQcwGa0JocfAK9CsUzPKQCYp88NbNB6n5ZaHnaKlUACIwe5q/7SzOXe7IQTZ1b
EfhAX41MdM0Q3+jUtHJrvHRR05Nt36sMj/w435TXDT+Idc3KIGwzRY4YcoJPKTt0
oS5dMMhJLChIw0ZRMsx1XZ9Mw1xw+7SRcPxaSZCoRvaCe8rxdkttNeHqxUEH8/Hj
1RZuCWH5VNT2JCSBaHAbipkykyLkqHzB3cj1+VuzpyfeuiqboENlS2Nlzk/339jR
MTSlXoxZLbdyDGbuWdiaCrHYSbSLsLEGDjhmbs+x0s6qm3zJ851oqVpwfxkVi0mH
v8dIhENg42ishLk+AHdKD6lJer79+BmNtbyY2/XL++vpIR9J2K+1E15prdjiN1Yu
wUrXdkZAzk8Qx4JgYHqd8QUVodG9oJc2lLn48s9qNoYgebd2P0V5VaBRQfNLu5Nv
FP4R/5Xmk3BzBKjTa8g191x2QoFI6OXnQDfDyI2CFK7xlphPBOYtZqWeueYm8lQ3
Nf/GmS/wQKcm5AKsvMOv58r0DVNncEp3xj0KjXvI1Sy5mq1HkOlFAd3EJGuRbfq+
g9dJcyJ6fPy7h0/D5ZObyyYFlLGtwBL9LewiPHgVu7FtyuMprICI3CBRKlYjbO73
HdNu/yXc8sHwYkJVmtbolbo/VtgPTTzbm8T5EcVtNpNHx0AAlJWrb5j0uNsilel8
G8/qMQyXUXAg+Axwq2qnJvOaKsQHIZrq8QtTLQK19nSGTdqz+C+AN1SPj2pIJZIc
T3/MUfKMY5ZFp3bhD3PCqoBsyKxEd62UvSTwDgmT9ChTGpy+X/Q/KSu+yUgDYZbp
v7QCbNSvx95Er9LygB2fuPeAogk+YkUI/WcdObOP2lthAEOyJwcnRod/dhg9YMpF
I/lvlfiI5P6ceykziKTUzzUKkLWBmIC4lu+KhQNAsOAxQPABM8elpKkEVAA/LaUK
A0JcKvTBtLWoii2d+tFuALZYEg/BzaI0K5jfxZsOg9b0J73r8daFuvXavH3gBKvQ
IcRW0mSQfoAcDfXD3Sb+MNo/IyO0n4MQktNmS+aj5nA513hSA7SiKONyhfM11Jr0
MQ/T9wZ8ZTyvA+XeBKv+5B5DX5lCyn9fBr2dckUg1O8iBqSCclwa7jeqaI6VNNmt
ho/OpLDjqPT58vFdPGnSubCD/e6CtEMKI6m+OJXuX5WpLBK0FxHAAYlguJqhlMvV
gj/NtXkRujcrkN8gV/W6xhSKq3NdBQ8LNG0QJS8y4spD4rNfm/9kQ3QVdHjqqa86
qQE2a9OZB+x5bc0Ez2NsLTXVKBKBQtHzD8mX32R1ifi9Te2DKTSk9XkxbWZ/3c5m
q7BK4ihZrUAgcZMdJVUo/DOYZLh5VXm/c/pgWLHh6se63UqM5NwbCW32TH/5umqq
iUeDVQVDxfqjm964OTNRhWw74o+Du/jCgY0WJp2yvFCi4pZ0VjHJ2vG3XWAJwLuE
lOwslUI2q/meqllbP3U5R3slyFuBmSlEhanT2g1lH1kQRQHfAm9CS7U91Oetksxh
DYHBJ9LNkntGMe5mgrGwObpavriRefyPjThXbmvBkReW8SUm3RXGcWKXu+O/pamK
fiUpNXUKbWj7qrGy1Z5DxJahJ6kwR40FgAs9zmKRjVn+Tb+0RTjsRm19Oqxc3ftP
tR2KvvUYu/oFuwrMmGHnOdHKVM7O2Kn3ia4VZYKb/k/ntf3sKKuDNCUr4KqbXXYD
iLxylrRswBvEK6OfQ6t0EbWBzlhghecVkBEQ0zS/s6XkwfWyARl8rmakVSksMEWR
qjQJ9J3Qsd7d/KaCqrXElsZ9WWKC+es3xB72U0iWtLQie+Rwaj37x8C1BY8uh/ZX
I7nIyL5WJti5lnYswknUOH3Od1KSCwIwOk4yd7YSHTsaOrclCpn6jxdUA0N9k+0A
AnyMgGMMHW1FVanMhNB8HiD6vs2rnlTQ7ALessI+Z6qE1XCGTZRhKwSSkXr9eyDV
BJjOa0VnWud5nl9rXp7YnkpZrjtYeK3yMGL0dTJTvkCAf2MP5FYYMOgvXk8E0Q+L
2NFuw0R8H7zAgN6z4XB3DnSng9KLDD0xFNmBWFR/SlKOLC5px8tEC1UQYeXRYXz8
QjA84N7ZPx/kTYA85aKSjadCdB8m4qGuhSy0CL7TZ/uYR4HgrL4NunlXS1Pems2p
BsXLPclP8PJfTjgO/rtZEE4mwV3ed3PDKB8ykoPjJM6PCxFW47poX08jbpRxpBEc
vV2CFRNg8ogmG1jjgiq5W5J0VwQ2AZN1NIjcOPWJsKaRVCw6/hGBIUoec4H536rn
UGZpUzf/JSMVK/jwoGWpWAFftcOjOmPZyIwQkTNE9Yo25sg3yg9YefUkBJgOcsHE
FGFEkT6i0Nv2cJ6ZDijc8mk318l6asvkY6ZehcB131ZnBd8TLn3HhA9+6T30rvdm
gDpSEgOqG/Ne1dvuEBSPGiOXTG+2CzgdKGxQ1xK18OwYBo48Xsu/SOxKJrUCNfuI
kJPwdlHywaMfPnTROst9ZvSTXOBYhu4wW32HKec7TcNf/zhZfe0bPcPDtmDAv47M
zApDqZwr8QvnRJaMv5NGMw9J7Xwuiu+Nj/9TD2da0QFKn1jFdlulN8piHLjT5/m2
hnlg2D1t17hq/vUuPJT/UpS+Ktcf576Pw0pjERss8A5Lf08R5NTQB3atE64jJ9ZN
EZmZ0Nw1SkrzTisUuzUlwxaxbKzXmYIfUsdnxzsBgi6AV3q5Xkdi4zEy0iQ16nTZ
vfZdHph/cYFJICgLfGPZPobES/5QaKVIGCAojKK/E+y+K9Izzrk6xQu45zjgeYOz
TrtC8Ky7pNa1XolDaAQcxt4MFpr+S4bHJt2chvinIYVKvyyB9o0fsEkq1WL9SvdH
FRuewu8K8DPEiji6Lnx28/b1ltSA8XgGVmsaTgCN9k49Z0reYvUtr7kUG/NsZF2K
LjFDSEbZvO0O3b4xHlakh0U5Q/0cY6V1dRTfEXHOyCIMvEwT1FC74sggzntm0dNh
iI3O6+I+U/VG1uhynUTve2tK1+u0PaRmvsKnLU1EvQlIIbHUjbXK8KoLaEZsWJhP
aP5DX+dQmkEKgN6+RABwKmKCymsCXRxULT0IW0L6pg65bz5u4de7jNoGrJeJNN1H
zGP+NKCy6WP+B3q1nuRYD4fPS5CHuD4qNYKvEIyQnb03c1btDbKepVYkPW6E4N4j
x/H0fVVX2k0lpbOPfZ20YYGtbdoMxGUUvLJpI0ez+dt+zH8X4T/dZdfw+Tmfl8OX
cpwFPm6IwaOfPB6C3XX+5nUx7qbnlihFIU2mYeLvNR632fQHLpxzr6VY5xUuD1fF
SIna+e8mknMR0jfvEgKnBcmBLiPIBec+CPR2i7JFoTjQjPPUDBWS4MtY/Vt4Cr7t
QmgFBoizKDp0nnbpKKN77sCF/CZ0l4T6BYoChlE0Hrtq7PYnqXDAhFmI4cZMv8cn
yCOqx/dy7tJS9qK2txz3/PymDVKZL2edsT6ic/R1gviuUL7ihaRyz+7FvSw0XoD2
JaPR935kiPGJoHHRef07UbAsBvkMpihEhXw3e4RZdZXQVNAP7NClwltArKTWa40W
Pdmi0nJfo6Uu2cs27Ek29V3QJFOz6FtQhSbATYnL6vQcFiWd0sP+aoVHwkRzwpbE
92xCtCwD4QSNzqa7aPcIitPrwHMTJv440C2P8fWMJHuCZkGB2rf7eQQXgVfLX/no
fbqgc5ZBzuMRUw2uHtzuMby+7ZKLKa+5eh45/XNVHVkPAx9VG8be9qh8R4QRykw9
QC0z3wdtAF1lmsOlnFdorBygI7xo+8SO4hloQIUbjO8jaVlsEMNYSN0994d2x1Ke
hemqWugOqVzd81n4+m1c3h2ljg4+ZbjcWqfNXQo6Itg7TQMA7bYI3uA28yZPjmai
yBRR5WV7TIGACFuPzK1kjoRbRJMADXhyzIOnOSjMYsxvmGy7/NTRBGN8S0AVcDKg
8rzJUeN/MUU6QPQvbVFMl5bW2LUZC6x8iNkgdYGBugC34NcE4dZzkXy75v9nbS/K
FYGURzegi4zdBkQ7WBZSJrpAhQy+vVOu7MW0oQqamDIRctThWvOkst33EF5lun3f
S6mKWz/YY0jQayibfiKpI8TSnW1MKg3zOtaKa2PRXhBzYnEdlmHtHe9+Cd+i7khB
2f62vxBYWPmuIR4+Zt9QiwAbHPQ+gWW+eG/4548+0k0kF1tCUm13OXvuHTZft0Zr
gu6qAJWRpzLLAe7CZVxD2CO2SrLNbja6ObLDOwRt1ebs5pBIGxOho7hK880L0A2Y
W9jkYW6e2hEHHzegXaPKimpcJDHfckROp5GoAnhXv1RdDWotGZoCuGqBY79l7dM1
We742JTCEv2RHSzDPOMrdM1jcZFo3yEQIP6QhebmyXTFfTo4St4Ooi4ENpgwmEZe
3iBBRq9cHBS5hKfDSy7l3dvO+5asbMSzI9NMdQwolOBzcaNKsArj89wWlEpBkmzC
Qzodk0KlQ7upOY8Gn+UcwLdHbMUhJtBqsrK9YDV1Qe7L4PYPu57YlrnF4lu1npfC
yG5pC3HLwkY4Irz7bVt6B8HpaJh+4XmzLLoqL25QyS2I9GrmI/d6jzmtaLoLCagY
bcUGKIMx8qUHQcGTC2MbY6wl60EMLPzKclV8ztIk+MWkLZxQVxNs+2dwehC+6TIy
Ql/TmQwFqU+b4gnEUemdl5tB1zb+Ar/eVll3coJ6tcpQ2gymuLmqSL+hwfa3qWvO
9FT/xoGfmsj6Jam5lz+m9PKHMfVV8cVKSe7cudX+QVjtRyRjG1QVsGqmjjhgf60r
I9IiNX3RYGkpSUCuuOhWyc04KF2qs6k6AW9HeEz7F5R6Ql4XF0ndCP5FzZ05d2lb
QKzEH/w0dKBvN1/QYqBvNkb5Tc6bCv1tj5ap/CS0lV68r8Rsj540TIC3mXro5YMO
lxvYZEVPaVONpQiia45TC2eCC7acw3l4Dyhu/fs4iYA6y3WAv/8KlxOuYSx/lRdS
db6xn8bTFnkTYx4sSeFAGr87IokEUUZ3l2yT/t4tPMDldg4tp+Z8j06JkgRJ1wAY
w0JkSuv0/lvSTitPboMnYwxPO+0IraDDaO//X+B7yEyGT5I/qyVBjonNvitdm5ad
hUjgP4qK7JuZ1+TPtfWpHnacxPfnKcK87uif7TfaGlfSkmLYE/CnAx3ItAb9h8dG
dIrpc9TznLt7NR6qqY6AlWJhP4oYWqzoAAMPOEBqp27oR+4xB3HKmtXDBDWNsau8
u1ck63dlCSWMneIkgnrcdrL8x2W1QQJZZ2yOkc9DAW2OahIbKjMT9rYHiE3ncAd8
ZajraF67jFKODWGHw730NGf/fG+uHf6x3smU8aHtpRl476dUAAGrzet8GkVxGXrS
0tjxLPQLWiQ5UrI7I6tTsGqQ/MUaTRvj76HHgoIbcaEd38Xl4QNBPJYihGkumBQz
dwHvPls2zoOnqqd32iFX2E9Nlhj5X7NZkvSKQdYgSeiwJ3/Mj4jXg9k/mdY5EsOD
KqOvV4rtLftjjKFJD9qEP+KszRF2Yb4/RcLO0lyd9AGmjeyx7nbUMk+uD6xxQ+As
ibnWTUKLHhKhzSY94bQYngMK9Jsrtx/C2ujvuspxFKJK+Rs8Np5NuDHBHJ+0eJ+O
M0apqbxmPBWzSm/XE/HgIOM69pXEp6wBVuCflLCds0UC0aHuIPjT3tkTpQBgyuik
H1KCni09THkeEIeYpSzIqhDmLwYGW5TbgVoCMBIp5rGX6JVDUqrxLnjQRWmtgzv8
KejpOhMtG4UVcI31Tjyao8CbvW4SzHYW1Z0ZiVl2gVwMQgwCofbZNdpNxx9oDemq
y/DlSapzQN1QwlrOygUtwuUXeXW/iix4NVc3wH5mlOHDZCVliT13AqIrNswQ5TZ2
nkOHKmW+L9O5gbk1gZyT+0fZWserkQ5r7OJpNh+iostwzEkI1yFvU05LHP/qzD5t
PJDbMeer/2tTtT3AToAX9ZS45lNi+vqctNtPQkjb5K1emblH688BRV18nvMjSEG5
oqA3MyAq50U7y485GSZzAamanpKDrWMacEeiJ0un+xM95S2ucG9PX8/911NvN2sC
/OwidTHidVWO+lyQxWXEAQP9c5gtYGUCgQtGFXW5vnEhhmDJD54TfbXuzfdamcH7
yHPcpdcvnTDPsGJXBIyLTmPeKL9pzo9Jv+JGzxyXPSt8tlK7r6UYxwR36PmJEJHY
OMte9pnTGGjopYd9lcGVz4q0yChhdug0SsDf7U/HcF5wXRic5FC07ipUoBsqYcFe
pqeRnJe3fxLLP4r6f7EtQVhOnnwDM2bqGe5feNz008DJhYLQ3OdP0aXTQJELZX9g
J2JZV9mWEbbI8xHXarfkANB8eJ7qxZFfPVEXqLe17t+2PhTjme7or1OuRdnaoUj0
BC8oNfKoJRds69uQUc8zrZckHyTRFJrWnDqggB+dlhK854LdB+Bu2Jf3g7McVqg4
9eo5XAxza9VUApsuFzo3kXs/gNyhWu210Tk3xKuD9yfXfVXM0CMCwIZLkmLPknQa
afT8F9Bnh5NEqQT1N2d70k3VbxJ8YQ0tI+iMyJdsip9ilH3lQsdDZd6HSkCi88de
3mg1iV+X5X4vxcBRjWyyijtflz05mFkuKhPEMdrfJ+1IokPm8aBrCId+6b5XqsV+
Ru/36k0ivLIzLa4JXjh6UBU5d4VqX+cKeZMiclojqOu20CQ2j9ei6l3KOD7wvzYg
EVSef9A3kMYy8hMmQiP7e2erDBDTiSz9YgesoBvtrtUJ+nNsxIi2Pt/mNrvVmHT/
hrQNhLXPpOavCixp6kvQjg/XOHzqOtrsbDlPZWiugs/RGhpZpWOs9X/YE6WLpE36
wPCQC55hEPKbF6dviZweDG5yNiyTNM6O82kAsaTj0MVeYG1cBvNjxLQb2Jm0VSNN
TGtufRU9wO9AfjcmEr8uNSYvIw5lzI0AGJccdk1l/JCA3l7JBmB9fbZt07LwkErf
+5j89JXTMBy5/ERL/OifhJ20Js7CjPbTP6GK3yL0h62Nb+eOq+V2ssr5r7TVrrEj
V90qNk8SO4uGknzmyzpsmd9YIKQ+igdxysSYahdwWcFKW9NzHFFGduCqepj6u6Kc
9g1v+qXBVrwIpVP7kwlgqN/kns9P8nsTBpQTb65YrKJR5e5WsSATeYYS+0ULeXWu
eqpGePDW7JYr82do3ofTfn1N7BoSaStVKAQR/NQrq7CzXLGbpzCYiu0gTyCo8K2H
gz+lQSJm68QWuzy23E+/uMFKl2uHN4JJJEQqH5yuvzaWWZwBpW+BmU2VTegcHM9S
VkwB6g5TNnDtKxEkLINFM3r3wGObOLXWZ6beNvVzOS+1wscLWh6dOhRO0Oz/nSsh
bRMSv+yi0RGA02GdExZ090IRFbkfvFMx+MFKwXR29vvgO1IWjyFAWcW8TSWQOjl/
PBGPvKvUaEaeEXuBeJmYn3xzJ3+zp8zx0CuKOPM8g2xaiU1T9S+39eFWTuMeKxt0
gRpJUovofuNcIs+yhThOrRvval7P/kycZ1mBOJEGD6zDS48eVBYB9KCir7IpYel1
lyTuHgow/LGdQUoWuz1y04x3GXQbeW++nHT1IZIOK125dvI1CoUiuhiOwO0IXpzc
YYWzbEfmLqU8+GcuI/ZoDoduHgi5GdEjFAY8z8IsCuCB4qQ4iSfd1vWjJUYiThEu
qPQDK+sqU5LjTuO+ymmT7FoKHCGYqJjPIIz7CkTOQwts5bpmgEcT/ENmApsJpx7w
kTUT6zKcmxnUsYbGzxxIAwnTGDG30Y5WNdMU9WD4OzyIjhaBa7iWQznY55H897gB
tCSTzvZF7IdQJ8RBBffAwiCUjjU/+RdpplP611a0+TmCGG8AjgLKF1FvOtcmATQa
l4DBycoErXc1iXvDeWE5V/nFVkCl2fviv7+ANhC453vo1XrM2jxgbd9d1PEaXTFo
OsVIIF5Xr+xvu3NE7HYaMpoWo1RrbWBVzZA+cFtBk8zoOtwF486EsC8zyVIer7zu
/KOs3i6mivKKjgYn0nLfqJOpk7apNkpsENsqB0uUGm5I5cFVosMo6wo4uEO1TBt+
A9soDcWFwkFBCGzftSqidp5AwQurelt0QDKJ9FPizNQ8NnAUB3J0yhBnkmSwlZhd
AKJ25mFk1ZFQSSS8dN+FqImhhRMACYdyRzuOuhLXcAGalfdicoaRhASXs+s/npFb
qOkjO2T5naISva/fLV8CVkTvfClLAkUzujgAxcC0DPj4yMCa6Qpvsilh8bKTmJjz
h9vOiMqYvLpI43Y0AZ6QKbhrmU7l8ObzEy7Qsx9sSIDny2BhxDeqUr+3MOIXzXNO
/Z5Hwxnwd7Bmi803zOnhzMmZwcCiG8aUES9oNv2buOR2TN9eCsZZFvDhuRnQCGsU
5B5u3FjX49LPJgrLiJAmTA1AdtFvpkOF04veWySBCk+I03i2f7iv3YglXsOmhjhA
MN0yej8Fbsy6Y9vtdfaNahwYyvnN4AjTSKbw4kghlLn6quyFQuN0HIAIqq5ogYah
p0w1OWGV2iePOMJnmkQ+nFAtXycUPm/dZbmskmF/R+gk7QmjrAGLhQqTwS3joc+8
6L0qy7bhMTi+/Nea6kztWSqnfwfzt5AbNSSuGSMpLvN9MLRT3Jc0lvSMGMmsMAB+
AUOeYRfMWQ7FWiylHoEhAHFb8UXOcDlarqlxga+i8GpIxdUYyuee+I5QGaqHs4OZ
hSE8neCruYg5PYsnDr4MC17t4TbPDAQVw0Nbrns9wF4vZnBo2F6Rme1LFHodAWkN
iO9PbcLrwEgicx65XgQWthW0jIoC3XOpNyI/Fp4UXlXRB6EJOlbbEGSBusWq/CBz
aDNi2YHFjvv3sM7SH+tGMahI+50UuTlE3RLjpuvPHXvZftO7ABrX8Chvacshfj/O
erQin00xSGVAJFI5w72KkVaQInIKstTTU0jF2Sf2i7dGw8I40rLkh185TinrSB4/
IyRc9j5plNFno1LttUWXZMqBbaUwf5ffVxrnVE3adOCpVlYbXmgZlwT5PldwmHcd
Gpr7rQuT8PBxDSRfg+cK42V1cDhqZhQG+7HAE3GLUcVBFUKJNLF3E27HxO9iz9DH
KiOVl29TIlAmMzIlSR59KvcyPAn/q93JiiOQqSPN5aue0l/vsFnhnDq8emjo7n1L
PnUql4d/9peZDaLG4iR5Y7jE4XE9j88iDQCKXEyMSzN3nzsdSjGGWmWq1WCx77oJ
gVjutMyAOXwXHy4BRer/Cnfkfmp2T+xq9cpka/n6L2EtAdW3/E52iRxTqSlqQlEe
sKBUcRJYzlLTCgWk3vl1Bge1N5GX64aIaKIhCLMY5DkJE2RLxRRBqvrd+ws3Gr1Q
MV4t/SnBQppmr2zRV9cq3g/u4EA/tQLSF0d5jy5EtzYpmgN1u9jTOj8N4Ih5PGak
AOOB+JO40emsJ+MuosqKXFTpvwqGNhQ9N2zgYnzGi59ECBzmZsAxSXqqKEp2fFzo
CdVZwebaYhmb+7QhzF9oYIDmdKyPYozesvSP64hnp6xcPHYsOhbUkWytaLSx18LQ
5IxV+ezH7UJi8h+HyQ6JctqmPgYHLOsjLFLXb4BxMyUIhx6TTrNHWv65iS59g/Ps
6CPSkQiUlxEnuJuOM1jPW2xNhvnco2qhBpvOz8EksZMGXnyv22jl+ERPPmnPoAO0
WC2y+MJ/OTITPxSgX21mVjcCk2Ql045obmNOIXZlwGTZCH6dXbaUKjN+B4tYORcV
sXGXCIY9iKKsiAmW2cweErUv65s3oKQDvThOECPu2j3e5NyG0p/zdL6ZW33CU3de
Q9JY5IVdJsNApoXPH6HrHcabgJRZExd7neFrUy2t5nrD0c4cfPWoBe9Qptp2FWUc
8E7SceDu5XJDlWh01DaJihuqFkuK4XneDsuFaVO0SmjiB/wuqM+Jbi6UmIKupKsk
I6qD1nViIzxoeEwUqWmm/7Zc5vh3gTmkJjMtHze1NDmOpakugL4B529o2afQbIwZ
Cs8umedAKOYNPYxPmUIf3sgF01i9SjWfYjWC7basf012snBe7XzY31AtkBB4wf4Q
8q/xEgJd7ZBsBr0SYYxmoUbbqC2tJeTNBN7LQb1JTVHpRhNdM2vPs5r2D/1i06L+
6BXGX/+BYP6lY0fvvOZIHP+GV4ygeHxFh6Teo6J2R3745phnAY9IOPWTOG46ihUH
edWoZhZp4qZwc6BCH7/N5oBahp813szrVyj3BwkD2xcNF7acggLMdaDtCmQkA3pG
h+e7LGvA3KzAutoZ7aLHGCVupv4WGhxQxNFbp/mJ6ANez91ooA8N96MjBL1+Q9O6
uWqqG1yZTGJfqIO+U2hguCKdQ0AMWCTLG04in6/Gz58Rl0C7apsO1R52O7lO3VA0
lkU6EvIDkckGqRkyfEK+ZEAJwxWXJbIED3K06JCXHEaXdKZvChdkad6QX9+sytTi
rBaBP0mrcZmK8IgSxk5KMRraPX76xeg0w4P4J8RAd4UuyFnWWQcXkrocqdWTWVgM
jYyY/bP20PxeHPABf0XFiiJfdpEpmlsZaN4WqYkHfcCVataazsTd6zRB/fGRHbPA
nYXwL5DKFS/6kwvVzh8D5wtxiXqA4ojMEHnQsNAZLydZjg2txedPn/hizvCJgZ+h
1RHgehz3ZHyLUYYeD/buicV/No4R5fl4ffM6S2+U57NhOKFrds0ILi2zbDreJDOK
SFZgVgeP0JuhoOifeOuF4+Z0MPtRC2CFCUI+AT/VLADwroTBW23jcqI9j9u9baqD
diVXf//YNpjdI4XKgsQgOh5F+w/vID233uhOP2FaKmeZ/19g7HoARbc6ZBKd1hzA
KWG/I1c5O47b4ls5HI+QTU50u/q4dXKpXZQ/FTJTLWUAN9LETwxa8FRoDdzP1Ng3
KYHXQLOFUe2vr8nYlmRZIqkVj/qEOfBMnFN4NAC5Hxbhhyp2QbsDCcQlbW/+cn3a
6MibwoE+gzXra+CQKIPnlVDwsH5A+tR2B0dUA9luZorOCGr7Px+KM+SL64cZgna6
thhX3a1M9EJY0ARdBjv6z3OB4mNcO8LC5dolYW1lwfAnTRLnqFjOQFuU8lru30qz
PSL5JuPzhnl2KVU/uoUS6YQuhlMmARblQ9LS27SMr0ZrBVA7yzk1+sc0HKnXQml2
ZZ28d8cv3Wq17ejSENk0asDjk06t/Q4XbEogkOYvPzh4dx8Klhw6OtIrjR9NsrWN
kvK82Lry4wbbr94tN6BhUB2JT9BJeOFYTcaF6notLSreM1KeHYBDWxXM6r2ScPkW
xnmmzih/8WPKiOGqMsCCWe/S/MCWCmw9t6+ciKzLpGcT/+/DKRsbe1alBrUe2VhR
pHvKz3bPIvzHuQcD04TwIVHLWegJ50ckL79dHNduh1pCJ/1ZCAzY1cqPIrJ81RVn
+ZQsJbHcl67nSw/rev5ptMpQKY4UH+IIDsZi5zxxLgYBZ6pVC0iJXRvPwAri3T5v
51Uvj8kiedA3D4TT72e9WQN6WZFIbudBNv+TkwNDdmi0ZaiTWeqHfKkaRqBc3JLq
RFkMzc0dt4PCHiBDSHL+i/8TyuqTxEk+0cdsFHETLnHuJFMGrpsC6xJQxBLupu9K
polhmsO4Cl1X8S++f5NRWmYKoBYskhKNIGxBYsiGn8BHEckjqWx6s4RDP4G1X1D/
rahG+yuChMy9N2vV7sOovY55BY5qv+hREAquR/6s00iibtlrCpzOwgidlskkKagx
XFeKcrbnqBu445lsJ4bf2q6/XEK+CGq8to6I+HHbQTdXUdFBeOAQgnfblsUPmUcB
WoSUpWsz3OpXVe+/CzAC3RrsXeqLVxgUxLLl+b7c/Z5XvMgQ1HC9ifQTMy2/fSMJ
OcV0lHPPTkhP2/gjrcvfT/PSSoCYsr3cBWgi1rJrTJGJEWyMkQHys4YXqDpo9SmJ
KYHpxK1eTZNIPxVT+0Kf+PRWFq5E1TfS8L3A0Z6ryCpeoF2qghbs8dU/ErLhg5a7
e3SDayWrWN0pxqipHFP8yDOmNdhv8APCZwjF4l51vawtnMaBfyc2JeYjGs71rKXg
5GurN396MQO86kN1wU2Ev+L1AFgbPZHnEJRUSeJrUTipmzEhvUWybOFlenJMoWhc
2N68wDZI+MmiVakXpzVrEUmglKPbZLhlPBKnztTgjv4R+9a73vaDotoVdRHvG9Pj
7IA447WiccfasWrMc5RsIqLYd+H9TDcCYhBZcpt8dndX+iBKa1IiI6a950t4syay
wLl2oVAySAI96wKgu8NJtL8ZaIGhwAd3Wcx2mjVam6n1HbdAcsmGxzgitoylUpWu
yKu09EsIqqNmSkHZTl3zRA5+qQjuMDdSNt+Cz1qxdmKUgvRBFgmijvwZcAL2nyIl
I4Bi1R6rWlAeUZBN/hFq22Qm+LtiydOHGP1NZ9t8KAS8GnBroG+JqQhMch2DEeic
VAlR9c8wT3Pq84NGAB7AZifhrpkiSGR52BXvQ0aetAVkTl7BY7grmuRNCUZbt8Gj
S+R9uyGlceSrN333VI1NEk7qbxs18N+F3aQF92bk72bHUyxV6Ns6EA/f+oCMnulv
pxIjreuy7r6HdGolwoKiZKJX9qPXdp799l8hNpEwv0N8zYBrYU7lJeKdt4rU8Mcy
zGky3dxl+YgMP9eKTUHOAGKDJExLHsch/z1wMp5ZukFSJz/RGtr9+MynSA1h0ipX
QkjtNR/PUwgoS/XMt+ERxQ9HD/LK05pQ8BgOMN9izb2ljxQf7B0mEs95yRYq1iNi
MErYFKxIwkUwLICeJa656I/NxTZO+JigJ1cDK1PL+LPeAeAJmFFeOjw/646SxLm2
7qUMtuM2WbIRGQw3VLy9xKW24EUCCwnwc90F73UMFKS139wD1qv4JY8Vq9YuoTLY
AkPLpkZv79I1bLTSMK0VyKgJbpR3PmKCWzJ0rAkIne0ddNUeDTU+P5Qb2H7+cbiR
GHtvUxW5t6Oxk4PXqaqE1+QfN4LjAP7JUoYc+iNoXFcVEAmLIc8xHWRdhZliBP7U
psQGaCuCijHrl/mmAgCYDQyFMe7ARd4n7dE497OxxaXAauijW18THBncPavfD9K2
bQqXQPJRfpVke8TB4gB4t9GZYD0hAuBmoMr2vMtQMOskc+mS3czje/j7WzzLQ0/1
PySOvOdqbo4r3VlMekV73qCf/edxdDmx91ko0a4uhQxJUkwEE3S4Dl7FHfNaXNMS
e2zhvZe43wyVmCt4ozUp1WvBQeTajmQkhKoZBK3Faek754ZLZUwVuWWBhYeDm3Uw
1LvKNusOL7gpBEmi4DgG4VfnduOwAidfe4SgeSOOeV9hDQS+ubNOOQjfrxaF6krr
siU9ghfcL1WvTy4aqVw+Tfvke3+tee/SE4diFBWoymrShaJSPYWBnFl83jD7gwI9
8FibjVdYZ50mpnK6C19lagiZJPYsQq84puy6wR0V+aU7DNE3NY+abesWxu/KeasQ
5S9nQE1cRpio7/EeARQN16YvjEwp26TEYqADl59skt26wL/W0SlNUaE8Ed4Ux6hM
veBmAzJQvd+5TaSmVH18Q50B/Z6BoAqqtE/ZBE8SA4vC1DMuUnbAFX3c3chatPhx
gAceIyxG5soHVlEPoqzfVDEkvDYZKy6hefrkXSV+y41/4pHL31s5TcOqAn8eStr1
G5L0XkDD5WA3jr3Rx+YXu2Ig2ipI2+0A8vxHeyhcWcbIUvD2UA2IhqglMbg9Rimg
2N6Pl1HpshYK3VMb3m0kw2/rbB7d3kRhrglYbrJUY4dJbe/jQA4zrQGkIec6Sqvw
ZH7qVc0zlQKjeifPpN82ckx4hJmQmu6sn4vHX/wM70MhQwjyhH7BmJj2lqNrTExP
fQiMffdLBJ/i3JqcvB76D/W5W8JVt5bgQew37yhHATzmVIrZ7CDoVIT0oaEtvOjX
MIT338l1m1JSK0YYyJloRQjhWfX9IM1P2Z+EsnYCtw7YPFQB1vUxKamSmTD7Xd9O
uwY9+JXqZG2G9StLTKCJVm4zypL8bS3wFdrQQFys2ZawirkiFuqooX8ui04OAPct
1k8jeDNHmPbVcmREYX3weKWoXEWL+8T0GggxzPlyCXFxmnss0AFIy4DGrlTFDVrY
uE2jfnKgQ085l0pD59dOwKMYAR9m506YuhFeK5MPlFjbmVJJ83RyLGEQ2IN0GfvH
ESdRLpaHEjVV9JjZOhUQGwlGsmkwZkO+UEAZ+de1SGllQIkiWsXicm2bB1+OEFhd
tYwcZF61B4KbVB8MrNaeCy7Y/EUaE9ihcFhAf/5EhBd0wIZeEB7QzVjRegbGOUty
1QhA2VSjgbTmRTBAeufigE8Pbm+wZG4hAnHOJNE4L0wd5Ntwyyu2SfMx9IVchggY
xDEK5g63iGMm8T2yAV/U5sO6a0a+HmhFDTatGvIrkdFN0tw5ke8xuipklXfNUy6q
H7Ut8KgyJSrsjjZ3dfHPfqrr7HVwSrD5xKp+flxWABuyrwOken8Ag7O4Ep6+oe65
InzyZJClu7onQynncgC9h8dRIx35kJx80pkNjaMT870tktUe90wYua99XMCl4G6w
ZWuBwdLMYwao1jWRliOxYFZPOZrljcKT2Z4x4ON3rCIYN0lK85nP9k4pUZFF0dPq
UwsvHAK7qiKybQVoE6914fg2LmGJRj7IIdzjb89NJX5ou/Fhoax5k2A/dGUz5T3B
wBIoKeicbT5jFe8ll5ie54jzo8uKCcyNwhmU2aC4ifjbH7nQJaK+cbxVpIClgO3J
bLIlsjElo1Lwcdn+iWt2ROKszy9Rt5Zy+E3Hg1rPGdZxvmi4RS3sdfb/gUvbOXUZ
HJnHB7Bl6ituILFSs0PiRx8lUFE57moJeKLpYI8PIF73cn4aN7AIoxXHi85Uch6P
QZRiCCO9nPhWLcurYtkfUyzstv7mQ2gEKE7D3uN/dOSNQEEIc34yOH8XcMmOFzY5
mSE6hHe2lfbHOJBm4mFYIs1I0EkbnyJowTPn0vsqKvTMMxV9fy4bW1tUx7DyCLJ9
go/sQE0g7zezhYVct8/DiiG48scXCf+AXRa1/udgsxT1shavjzlImbYs1lOil8Je
ftjlwZ8x4lzLGYQCOBmxqnxGZyam9Qgx16SLGr4cnZLSQBUPhtAJL+XEjAqKK7yi
VvzY7znvwBbCaOeGrNvirflAfjrgBetDrAqxLv6055AHJtdGh4NzLMaW9ukpgzQ2
P8agSeZ9CfR3ECWh+xdkoq+0a+c/UPy5/iJrsBrHnoRqLEh6nvsDqbFfYGO0Nq14
tHMXT3R6nrsNoCALoU7tzV6EH+UYNK/2wU1HE8pCoOtrdR+Qi0xotlkpKK/l/G48
J64MZCIhnbZULLl4utJts0h7eLhT9s/eLl5YIEaQ8j3n8w21fYoAor0hs3fN0er6
amCMsdHcOetIlB/jiQ1Ucv/hVR81qlJhT7AwhuZkTOGjM58i1fklQKr9B2192Kdc
7nLuQawqFO/lUfcD/WgPbN5+Tf53wVDz2aKD1BHCnKuxrwHD1XePDa2OKK4cu4IM
ekIAVibzIeZBwLBIPPTk9YzZk0gfXNtMfgRg2Dn1Z0JlvUWrVLLBUJLNHe8J9CuC
SgU7ojDueZmKC39FHvwP4CJYAEsCa8Ux5hMo/8kY5pAqlfEqH4+ytCmmGtF1FABQ
vwz2t0MlLZKAEiWNH2V93GobMWIfMtaTZ+B0tn/ejEDCKwecyM1AGqCDjNQ9gjmH
z7d7p9kbS+pzOR11ueGjG2ZS/lTUvKWwKfLr2UVYUxkUTJu4ZZ3tA6kuPAsi1CMd
lxmNGQIJaPWBfRxoEJZG/Ieg49LOyOU8woWx8HbC79Ckvt7IzpYiOs1DGid76oN6
sxeWw7nW2RUJis1LMHiuSqvlyyWD/R/cFngjlotyB8bNW36bEqYX+0qtJOms1yj/
U832k05pHrWUHw1aSnb/H+C5xIwWLWVMaUwo8/hAn4bzYIYXZSnHykFGuukxzgwt
GBkI6/r2Vw28Md03qjQCI8YlFz+/NsSfFbItHG746NIiFCE9H3OC++CiPP5efxZv
YMnM0yjLnWWinPBHVMDD+e2dQEDD/SP2eeJN7hAME8QDUYCuiI2Gxz/wkZav6k3z
5s1hH25eU/pkJBR7eMHIjJ+Qndf1sJjC/taTyvkjYMfKkGDjj3+X4OQ71H4rqgLl
t8hfB6V6Z0Vl8Evkse+MldwSimnvKo0TJOAE6gsARcdPgDWrjouQCOFVzA7Jkf7p
wjUSdAeNMMfUBcr1E1isJSMtIUtNp0TQR1jOREKTCFX10poWOcLLmx8dLj7/Lem3
DoiwA1pjXjoNAXIKzncZ4cFydjriU6V82FGWpo70sNrBS/2IFS4ecnUPr48kPEkP
N6Dk5wBXntK5I+cAW7nYeSDBhLJdenrqvGyneWHJaMxu8Es3hIV7q7JoH40rm6Uc
98d3KzXQ0vd4/v+I0+3wOGexC1iLkwPXOsRrFnS3bMbCGTofq/JMKf6Lclf6YvGt
cgxzl0dtT+wTJ7ruLDE9X+GefNmmNiFEbZAbpHSsw2d5hxFM2Fz45FRzlI28BElZ
ku+FbxOyRjrCXQo8d2vqtOjDT/y60NR6ZXBaLVtby+4lfYivKmETVN36QDNeg6yt
VcXNiX7/LoV+PoinF5rbQh/enBB5q3yXIVGNFEuk12dyGtElhj0HJcVLkt/LFHX0
gsSDR0gJ+y2Mm4feAHigL66ZsWJ0CET9tmNBJ43fDVZsuMBCmT2BRKxyZihcpESI
7VqGaPp74iNOTQyHgTQMMOIN8haAU4GZWBybPl7gQDpDRiS6vd1NJjGHEmWag1WA
s2sjeQBUwuLqfIJjm4PLHWP8RaScjMRFfW8uZoGywmMuEyg28wbHN8AM7smV7dd+
gBngEtLHzKjUkE2p6Y6euCE+PATlDWeOROmZsdxRc/BiLr9gigrQUkaF1b9LYwwN
KOdQE7VnAm4Y8XWr3kuOQFG0L4TvHGSD3Tt3zW1c4JM0zod58TOXOHPu5cOOWLre
W/f0VuCBoCkjJyyiugSqDgVens14chwbTL92HpBSW5pDcTvrTC/KTQo1CEqzPTnk
66bYKQGI2rnRDF5OYb0/YbaXryN0ImGqBLa7nlBP2mgvWCa79jfZikJ45v1riJyx
P2tZvGkXrCZeN/JQXzh7xQ9jA3UvVPXx7yo1RfkP4XqZzYW+0p/Y5o6Bmmvrf94D
Iea6gBmzH0eWolh7p0PhS8w/nN28V3YqXN2sQ2WBmY8OHVLRS45wXV3rtAn/CLbW
MHzFA6NPdTa0NRacfHTeIi2c+FVMoZ/q6vl7s1MW/FX1NylEH1CljMrx/zAdYfZB
yK///Jfe3P6kDiXB+i7S9AFd/m9DGhkyQKPgRvoU03L+vbFbEHj5vx9lcUAJNMs9
Wp0dH9n5HeX7zb0OBIcO4kbqmPPjs6GPBh11sfIFZXmK3IzanPlciupBAk+n/LEM
krycH1x1ZQUfIoXQztfcfKz/3PEyqXXj4hdD/872jZw+kG0JyHF/MTRKG8VwKhjN
ARG9p0MzT6/bcabrIomPohGldRGIiuMaBp7oMjtm6qAk6bFFKdjgTNTzm/rcx7In
Z/hp2t9mBtm1bFxwqFscdR1fwf9JQK3v//DIRwMwlJDJjC6BrDkapMVfn+OoZwAF
NtpvLTCHkZOkPOxvv52ht/yefQiArY76zp+KcdaoonCyCGk5cXY0hbjuo88TQuF3
Ri4IEu/7YuTWTDFCJ06GT7U8tT1DkSls5sisEMknZWe1Z9cZI22Ab1LYRB+7+UF0
5Nf9ro7sYNPSx6FWxLVVIbWqqSIcTvKWQtAgho1b1MPUch6LF+XlH3UorCh+Sx/U
xvr7r7hM7xXiQ+xvSYy83i8ukaxSP1PZyt4lpwiu3PvjgmocWuzelrzKE39+QF/v
+l/WEcZjuQoHAkbg6YhEC4jWxSuYOJzs66/hXHhKPjDxqR8RpO9GG4Enlt9WTu7m
3q/rihBwBXtUlSQIidb3vlBvR3yYz1RkwAv2BWGCMFkaoGybM/XFPQ7kfp+Pqd+S
HXHTLyjBw++E3ZvpvVXhbDSiER2eRtutQtcHK0LrTYFtcazDQUFXNr+2OjeYQXaK
Zuot0Unstap5NI8qa7ivg6FYksEy13nEii5D1361UfDOMntJuUbHNWCWVX13LwZ2
/Ky/gAhGCWHu9S4kcPqPuQBhnQCo4KRG9f51MFfj7IIaaPhCHZuaEBTBqYNqkAPW
wBSpxQreXU7rVo3SnKxi6eqj5s0ayu1G+eMyI3C0scorjNoJtlOXlCN8l+1jfzJb
ayuWIYXbihHwh4zvU2NLM+9JHZPQvr8VNg/etXnQvvFRUqCzQLVI0IxbmJOn1Jj2
d4/hUGmVzdnwTFpsuRBGSHpuG7vhrm0LJbfjqC2FjK/p7ttqphEj0iOj90K68UtW
Cip3Ro7+tjisb05zZytjUqDx4cjKK6dhanxdYeRFVVwLB3IE/XfPNfl1eUaj0az9
zzoaamxENxu06yCXWWRBCeteHGhh1fz+IDWhh7lY9FWr6H7ci/V43uIcmybWZHge
EjblhS/1poLDVGyJXsHXYlGJHHAxmmCbVyYF+hH+aO9nTdAM7+3AXGYrVuUAuIA6
BcoyTAXcvaZJjeSMAo6WUmJ0OZrsGXcLOC3Br8/phe6hRSCc8q0zdyiTj18u8vtH
6FonumKB4x7O0i74pZY1vt3CgSWRchjri4jSawiYxEXuxrmIL0diOhytkg6ep2Y7
lZCaIYk2ELcf30VFMYbT5EaBvK3KW1ZZo4X3hU65+9GAXP9XiLGC1uOGwnulvwZZ
jgFn4Mk8PkapAEYcVCW8e8PPnpPzTkArh3uSnSVQLqCXM3VVApK3dUJ8CLC+aJk2
i3aUYvv5KhKtXpnSzdYyNHGxA/z3E2f/YJKPuevDGojH2ETv3ex2UY/f/dxxmJkj
MucfrrogDwZ4MXAF4uDsoMjuqQbhc5aZPMul1LZG4nwm/JvNVRe26qx5mlPtW23V
KLfdtaFxigBzpAxzW7iP7W7TsCbNiziwY9DLvwKLu2A+JjLNlqsYTho9awtYogJ2
Z8IWq2OIoPJvYe0UPHVJy0CVjnNP1MeZ7DeqqyUhVfBfDCw5jRFIOfVRQzSJakfz
T1OcWjTIqxV33/n1358yvXYkXCAuo+NGE4lqBazV2TfzTTNvqXXP6qjrIcl/pWfa
ZEB0T5d4sta3gYHzux2ovizRspw4gUAzgR+L2fIsFfkZaEIDCQuuC+TzPtSgp6Ej
fPsNRqkk/liQ2iK9Yk/py3MOnmZ+J7tXVR6EApyJ3yQlkEz6qLc80U0GVRXohFXI
PU9fHED/nuOfdpfCcKgtRm4vy9GMnILB9ZZY9JXyk3p4l62A73A/JTapkavCNd9Q
U0SKd37BGGTAqcdj4gPXfn8G9SBxFAENb0rWRcHBpGZchSm0fZb1ogklw8yOER1E
ijmNqXrQz2sFYb2pedxYfQOCylH5ZSucJvBswIiphgZWkWaB/w/k4RjbGHXCtzyi
u3tLmL9qQTCaxMPkW4FXTeV+PCW+K8tpjadL4iiYSiAzHPnWE5vvg9joXtd/DIqy
xcsamm8WXUQgMwXbapbkMzKKD9LzcOTFUBUWbOS9Vqd1SLCD4vCAJrLjK+60Jwdb
8xwR1bZIG/iR7KZp9YA2Jg8gk+LTzO+WIs5D5XbQPpCynYGdxpuF9DW9H411os7K
grNWVsEa2bHbo3bBB3eSSIDHQOmyQgxV7BJzZTJRPFs/mfl+Z6zKwj3NQEgBmHo3
5rleJwy/fF37Bg/3pxchRT4BYhG7B7WcFARyo+00gHKrI3TWSSgurd4lhKMTyfI9
WNKUfhTnr6oJ+cEcxL2RqUHqnZ87j8I1pdRzyZ5voMrrVkR9tZ884C8iU0jz3RXk
hvOKKWCi7BpNdkN+cq8bTUNr9a6MHXvSY+QZ4yNRg6KnFwy4DIT1z7h9gO+3Rdy6
LajE9S6mDhF+ASC1eawSMsuZ20ElmK5GdUSAKPhoJEbfDhusd9H0aYtcPsyPj6bJ
+gm7P1wpRg95yXO0dyWYRcvKDFSZUefvk2R9LYS3XOAEuJ4Hw4hXfEwtO98HkiKt
SGFGieV5wUiDmrsXJ6fOu9po9iokm4tmLxNO7TY926Ppoks2Mav2zeagbcMZ9aaX
FVz29KKspg3rtmHi+1rLOnk2RPK0jDUylfakNdAXiZPQT/PhJpbbKoUkbsupDj9g
b+co44L55n482AUNj2TU/MwoCOkAM9CLudzjZaZFYzaGOkK9yPA7g0UUtyT8tkFA
RUQYEkxrii37Ig+N4DCbbyiFTY99Z5hdHunlhRKK8z/OJI5Wo5UnwatKhWARU6T9
t4jwrOhcmolXT3bMfvy17LdDYC00je7VsmHAxQ2jhLTn6E1IYpp4XeTUGU6LafIa
CqR+rpn11vzkb4DtiMsgml3Sr5JtYBhXoqaKFmocTh2jLlBaat/mYe3zneZ7trtj
zxxSp3SuSIIU5krYTmE0AWKM8qXid1cgic9NR5oI9VQalmbbfmx3kLZxLmNvOguY
qeOeg1XfrSJMlHte1YGUyMjn4IcVCpgI3tkmms+WJT0DZh0V1tJvJ6jVCS6/UA4W
6PX5yRmNerFKSwtG6PJVojytmqvYB9A41+1S/yAls/SKQ4zxD/5hddQJXdzen7eZ
sW5jVTii9Wa3sH99sFergHrj5Be3c6R4nT1bNgqqM7zlhdQIBZ7rhK7kWY7hEE9r
8d/1Cbh7ScmvQ7jAyaZ+prl1KuzfGycB3FU/N4+nArghChr5f8xgj0r+nIS3E5PL
0v1bf3nZkVq/zzwQ22mWbiQIL4hsNWR4BGpiJ9DvVI6jauowK1fcMDlIriJzF04H
SKjvq/CgTqgcvW1KKVt4aDLQA8O3AiFda05HqA/938KuWdlU2lWwcxIZSiHigcjj
ovZhKwZmBp07EBa+aMbuN+365mwZhqRZwcJ6n5/IhZAGtMqiJ1VI8AS8V44Gbqxf
87dj2ZsgQEhGRHSSE6WkdQyvg6esutlugqnkFpbOjLQZbLorfbaTPfdJf3mQeeIv
jymwTN2Eh/bNBOZXEgyY+5qZHXVnET3kDBYyBHvIziAF5Jh4Bg1gf54KTzUHNmHY
OpyotdswOFWLioy7Ms7K8MWBmTusb9FfH+nK+FXmSoxuIARJap2WMAldjqJ4D/D6
dok5rCmSVT+eIP9xVO3BGFAS6uCFRUeXua4nXU3jHq1otRw6KgVq6q7dlZGNmKKe
kGkn+kgfuS5l1L9DawNGvIrrzO0AaxXIjFT22lyXJz9suJlG+Lss+CuYFM58Nctq
eLczPj/af/sEwoSbLzW31zchIeFj3VSMcg/7JZso+r6M+etkGkGkk4nqHptWJ5Ea
QyZRxbXWCWSZy+GZmPkM4P23uPtOA5n+SmdCV0CVFuJ9t67HEURuRFTqgc0/ZFsK
C9Evy56BWhoUf42C9GX0Y+YE5/MJliZmdU6eqII+9OqzmsaCxP1WfO2KOlo1CDJd
g5a2YoZqahBhQG+1lFIq24UX/dd7FH6oqju/BR1RjMbbhXBYuNnF1kEeGLhbquUL
YA7k3l43dZotT4aiu4htyiXPhMIOlMpZOTDGDm4xI6NxLt6JuBqKGRHdmV7/vOcB
Cca3UhLV2i7F0FgvfJd2xlShn+3Pbwuvm1Coney19+0kJ9amXsjkUKulPPwwRLOi
LzwIuy+eqy4uPo8tJdbAHEDd5ITbQdDQiUL2Gcixm49ajcfQEuq8Bl/Hmi13CXaA
CO1U094ZjE9BE6zG0oW0WLtG1KMkmMNl1sn56jn5AuHrKbdgbFA0p4OVsP0qED1X
CC3He4Waa3KofAjlPTCAC0R2mMQtoyaQ6si9rMooa2upEj5D2jglTu07ZAcFOf2J
4j5jUpMRAmsNtHs1s8ZcWH2tBHf63xBFGEE1K8l4ulEO2e+BmKuTSB66Rz7iOQhH
YFeNoHUSvyxQwytDuxO7LOEUrwtkGZscd1P5Hpb1SlN/ZIRVqbbxKCmWHJsPMrri
wWBY4yz5VP6pqBqblHm52Su3N9d0JHpflgQ04TioVS1EtaIKurx2B1ohRcHYDN33
7QM4DF6QYaPQs95kZcWRUesRwGc5fV/4k5yClRz5FeesHg5KEtQ+PQA/1wmgqXhU
OaMB1bxCU7FeD+4scgKRni2vLFnY2FWbwSr6TUVxBcNmniIlc2AH7NjRZl5Ir1BB
98ZqpuFpItawc56ctbFzExZVkW1LgvkmwmAcn/cbOg1hsjW2EGSavmj4XsbjvB5b
b1F9gIPdvpDxOO+MyZz6VyrCcTfdi03h+QHVrGYDgzPp/uy7IdSC/Xcybp1syRF/
jdcuVcg8UUogGQNEZtqHa0ppPiczCeObHs5SEPCI9AKbvYjvYfy/1KgzkiVUzwzV
5EV4HypHcqgQGmpGKX7hwYIlW4jVpLfHrQJXLTYLCJr6Kur2ofN7l9kMmJANDSh+
WzkQPYd3Y20wUaExWfqQJhk5HwLOk2DA1b9U6dPS7oVSeRv4igedLIKGR/qRM8Fn
orM5+cHJJUG/iMFPZFyJ81GFlJPyayKYCsKzST3Kiz58E6KKV8lovETkQYtjAnRP
YfDF7np8SxJz+1/wVkZK1FAo2d/LogItmnM+FzAL0+RJBiJAgMAL86FAX4w2okVe
uFBgFVlmw8hPYLhluVCUOdr4VrcLVW9LHn0lEGFbnfZhBf7hxu49rD6+swWcxe9u
wf6PFeuGZHsQ03Uk4l6qsQZBaWG2I8V/QSWQreaoZogcJb+XMLDcefSSxTaQVc5m
btqWKepULSujdKzSJcnpAKyKKDSNJEE+jKYsMqs+u0THGRY0Vl4NkIg0XBAvgiNH
PpbgjRFBnOd8wcgyCZNIKhTXHWHH+J/w5+bstbz7F6+fv66CfeizvSz3Q1CaIKF5
lakSokUix+xEMupUO8+ND4/RoXNkJY+AT8KrpPiTeRrcZh3H+kzSydjTT8be951X
NC99qGEcZjNff5pwseuWbzixhSRmrmzUCF8m21SNGc8lrz43EzllhxsvMhFAyBEy
RqAXJXP//OW3LFN+bhG0YyhK57aFuql/krbWHOqH0JqGx5N7YGeGmxkpHP5+Zc2b
T/R+U+HpACg/PrQvInmxTRg+V//zNs9bZoWojodIg/AFvNk23BhpVasFBz03Ycaa
ja2n+pJlJ8G14xuPreSI4AwyfFH6yfUISJuSkJ63ZsnHUy3yKwQP7qn2eGr1d5RU
u2JoIBqDKNWGumbRy/SphSg+zbLYa49wF8W7l4imK2lPF8wut6BDVaiIJ3ZsmET8
DcC/LC0faPlRY0AafMl1hRYpglvPRx/mCQmCHvMoAKby+Z3tI1GIMbEhztot2bW+
JO5nKLfC33n9dQSvP/GZp7QvByLhVDYz2k7pFJMCZ4Ru3bUaTjxMjBJJsiACH3oX
bSs9G8IO7u2CIApYbd2MMnBDrNAxxrJpsq921RmiB2ByPWK28Ds2YVnH9H0hvCl5
69yZvL7PPvW+VWq38fGBpJhMNRG4+hZRde/9peWwHGCS6KU82jO54aDBtF9VGA2f
W8t4tp7PFhffiQUR6AiRjhain2bAhg2Q/TCBS3rqUxHxwkobPQgNmzPSXHnMR424
YHQ6pMN/9NG1GeijLO3+OmpIOlH5kJPf8B3JYi8To4LkNSO8g06jDiiLmMB9lxeS
88IUMAssD7qXyFjxi+90XmHjiZrd7QN6T3BNCrivfsI8QU2Gh09k8RugZmptXL+V
VK4waX29us/5qEWyjy4xViodACheRDpuYTRzxVcXMVvuS9P0LUWHNHrD+sbSMjM1
q0zGPx/kOg7FsuJxz/E4C5kOhvALCf8QzVXy+4afD/McaIk7hY33/q2pW3KOMOlv
lXZGVVWLxuIU+TjaYBOvfGV0FfoELUrdsqwssGhp8sAdFbcrPt9/rDtHUuaIORGK
epiPk1uZjNAQEYPAi0KA/39RuuS7Ok+mu1zeKfzcD+VQNjne5plrsov6Q0rBePrk
0/citJIbmTX34xLJqciwPus5WN2UFx1xY5FDKsbVZmC7/TBVGc499w0Q/dLivn4D
w3tPP+qsIbEUYzG8OljUQCSkCbE9Duylh5IJ0JNoGz2YMhBt5fdXwzmDet9+p3Vx
ijfknchBY4/EtSW5NwS6z5JF4vESp0sa/+OazN+hcrsasekRhUajKiwpa/IUBuhm
94blkP+II0t5e4N3lqUucOaoyJ2IHCRW8YP5gWd2Ptze3HmGFm5UtL4Lzk73QG6R
lWisWSrN41zIl1P8DuO5lDd1ediKHamY14OOCAiK2iAPHK9WWzkXAQa7rURczmoQ
ZugNU6MZsILddSjrAz82Iz8bQzpamppBUl9lpbGtqq1GgIlSYpJQScpgmM3wxKSA
6cq6xLB21A4RTWtPEEXbHtXqvn6oafk91apA/L8khVaQsRzhFO/p9SzKIPnjEkPA
J1JWp+n8+EgRMXodl4fQkUp/4LyeXQbE8bK8CNQwXU+MooksyKRiAJlE7EL1RULK
bkpFCAsVknN3bD0QaF/6WV5YPAdp319S/EDCiNCVGhgbe6mQmBEXJFbP5sX5ZdP5
EuNBGne8IVrwHucvMvIy/ghLuZuKmQHbaL/dcfI+2hIb55INK0uLIT5dVaJ2V4Dd
3Egp3al3uvI+QJXuPVS7I0G7Juw7LqeigBdYm3v8KdUgyLnQ+PJVIFzHNXy+swXI
EylNsQme4Z2nYwT0IaCmYaB7q52iMNhLIgLg2vuRfMnH4wqfDZAxrSoeKMAP0QKr
BX/X6syB6Ne48otCUT0bSXOpc1xtw6593grnr6gdmX3VE9X6c1UcEgET82CikP0l
Skab2KPeyFNtzW/nIMS8b0r4WGxhLEZkpGBYyqJsLoMxU2HdnkT4z7WHZ+HCPiym
+Ii3cPKaPiToq9emibk+Z9RuZvtH//V0RtJOqxokSYV8BvBpqSDg5UtfcfgwFtdP
wICZ5879v58UXCalfvPvqG/3F3YCkCw28eoFGyVZX70UzMmjFDr1NHyXmZJIJDqx
Yq50YJvaLtnITvKhKygcaPtajtHC8hgeQCfbZKXZqE1BeO83GWLHIiEGJ1x2inWK
4ArpZ9eI9rKcQFFHsXIhSA/Jr57YYQ3RbsKgwtYZFSkCo/nqsS2yW/WRpHB3xc0T
1IovHHBZ5v3u6KQRGx16HauldH6GusO6MIf+QaWsHWUpwTZ5lNfP+emK7Yffovxs
K55APFCijbTWrB4bSOXN/7abyLxMyuUosu+0w35mzQsXnLc5NOhnFH4SdMwSzTgh
ftHd0Nx6Llv+3g1zLN52XboHRxYm8AdCqD+ybxZlL+JZ7IwuPXgkyEDSpuJQBuFG
yMry/T+98TllDBqBuV/QGdwFT5To/DxGTzGpmaB/sof0yjc8BY2LB2Yo5ZNJ7YRR
37IGbx34MwGRzlZTq06ZW22qo1SsBxDw3t0wv9oX0EjBt/TiQKPqv7AxBmlGN7ax
WVq3j1NVqgPq2ITDkvQaaoz1467y4aMdFRApV/mAGRMOQz51j8RP/MLYMm4ZOv8E
c+F1ADipWicyJtHsAcUyqVlUEZrtlpyEI7gHPGm6r+3w4EU14G3cXh21/LNgHMUd
AartOukndElqPu6Txw64V3c+oCbw+jWAns+qOWqPH818xG9sZBskcSKnWHWNVV15
eCxABG+z4FLEIooAcGbIDHE9GtBW3YLeee9yBhHtojyKgdlQudGy8gdAVUNiXI0h
Q125Hu0mV8C4tolIb+SgG2bFzIrDenc5JaYB8wwVlkE7VPFpreP7ZghDq7a3Y9jn
uning9XP9+XiALrWwNtYBLOHQp07u1nB8ZrYAxW6sXaLldgZZ0ENM7TPCmlKGudE
yhK9V2kwcnP76Sj2cUGdeD5IVvP4UjaLf33dFvAcN+H6+BqN/Gz3GRVosXcX5ywO
T3U/YHwQI5aF0nU7qZw/dU8Vxb8xNePWyfax2aOm/mFItAOV1EmnfZxtw4DI+TDm
VNiKMgj1NgG5Dg017Cfgl1sA2musZRLM2Z+Tgr27dR+XFBasbOwWKV/8Q82Ts3nu
+3U5yr7PJ0pTRcsZnTuMb+sLp0ML46/ie0WwgEHUIeFANQPMeiX/voM9pbAL5kUP
Pl+Yn3Q8ve4zxXcpYlxYB8F8FNliz7kpqQLmI8sIA0nd7wa4RmFyc8Q+PyzQrc0h
nhTD0yBYUwoU/DHJ9Pn+5Sp1KZ33t2ga4+RW+bINCMJZsAD8CDoOQ8vLdbQdZv7D
k5SyAlP0fcAY7inE1+J+0a2fpLkOiPgSXfKXts1A7Jm69mZV7C2VVM2zPMbiL7Td
yvejJf41IjDlsqOBVx9s7xvNZcDKQl3/nj3SV9Z8IwxUxFRh0WyRVdvxKHF2B15P
xVsMnuhQQGM2/z84yFxg/Gz6XicBTMsg9oYRroyDyAjVnbS104IMUqdUwEZUpnFz
5fPsJ8SvnsXnIlgUAGE8TmJR5jdIa3Br+ucV8JZwvLq6NmLJ3BlmWIBcw1wkKh7/
7GMuMYk6BPQDwK/3yFzWaNFRW+nILJCIqtWikyjIGYdV2paOSuLsEQJkksnRmjqD
ZX9Nx/92YFTgkgB3O9c4Y0oTN0rp+2jKm4JjIEDJMpjXBj0SQWeihU7Q2znPqAss
ICElnAxk5xYb8wqol5cGVyiQ1daj5pNJr/I7VTEPSfgvOsiljv8cbEaB0R6+IDTz
uN/T0auCV9b7vNwKpmVO7KqLTdmwmn6pGwZAfQZgeEUkEmAwwKl1GFabFaovpNok
xG7g7wetIvs0v2bCqljoyOtQQdAWTw/Zcvpp+moXMnaVXwELLcEdUw/YcvPO+vSQ
tGgnsrCZwqEXaaKd8VQR5f3FWMZnRvVBJy6NrwgWZkW5Qf2WsrShVZhWACmi427Q
oMGvoBq+ghJ6D7ArEYgJ2/ZRYrWSzjOECw6DL4uDl73PutXP/zsjjFP3Jh9pIIzk
YnCodog9MtsqssXZESya8Gy7jq6K6vNGm6GxmCHoLfQ+ro1IGJJSZucEGUhQO0wd
0/S9Mn/Cow2T7OiuYHRZC2yIGgSRz4hB0bQY7fpb16YpXYJPutcwEy4DkYL8I7Bm
YCXwxBvtNrV2hOsTP9DNp+d+Mf5jPyynnGsHVPtFrk8GwhqS9d1LZRwVRf6CF1Jf
h/UsSXNXgN1fjZNO6Xgfpc+8QEgKIXMXQT0YnQrwiNjoUH4ibImhq+6jy2TjG9pY
MqVQWlUfl7MwUg9LtVKaLkljQG18NHa1e+eZhRCpD7KGgdAi2dOOmUmNS/KHwUu7
Jf7WTcKCvEj3hFVSKiapVoexoMGLTL3si2bEQFLKQtPm/KukhQ6pdcanLxvJ5sMs
a8g+4v6+yvBBwdPS9+/HRuHPXRx1ukcUjnJMJkRCDkZQr3wF7imQBbKvzQHroiyz
c4VD9yxsAilsCfHqxg5Zcwy8OOyKXrnhYZkqFZ3gHUWjl71NLVWI9R7sI8puw1ia
rCK5qk6IKnnY8FmPByZ2xSyD5HF3svTI/357GwDVn9fJ78IkKvkwWU16GBmbPrAa
mV546u7UsjpypFlcuqBL3hzNVW26JTsLrvw2BLXZkps35IhDyEX+doEV761pqFlH
tT08+GgpUev/sN2ymuo6cz805OhCJls9QIEOA6QhS8Fa9gGu4VzHH4NlzzMGZocg
N/1a02dHMtMTZjU2S0C6fyNOx0tHVxaOfcNEBcyNH0fhVzv4mGxOr0ugdIa2VTLp
8lreg/b2I8UV2sS4/hM9gQLnvzVH3IAg6s/5v5xh/qPK1EWH8pEch2DwbVQ6YA0P
F8MlIriROpD4C6thRIW/Zun9W+KBuMiIUcmYvpXfFKlmYva06Pmx0OKKPiFDJK47
EOhsbbFRbqWk1VYV8qCa5i5cVdMlEGuUBI74+Yki9xZhVDkbpUrBoUJGCIWIT0Hv
+OkJDuVfrzYhCrDyjPZe3TxFj3nsTa8el9BpEfW4rZThJcQD2Oa0c7zzzOEF68J+
7JBjPYZWr9bjVVuTubBP6UVBZiSKlGAlEKf/di3il2UtRLuAX/Aq82ciF2WNNCck
AEBEe7oPkYuCrxFC0Rgf2FV6jbVhlqvoj3xDq1A6a6gL7C+CIs1DAGJ45OHrZgqn
/GWOTBXjpETxpgX9kpUgEBnofAbA6GmS9IIfD9pN3F7u4A3BkZJtuvgPZav1QsVS
IvzK1dbvUJktrlpIb3/QdVUfJgh/DDY9JOUB81Hm0jyLv6CW9G0NjgpCf3SMdGvK
ikQRu5NSkAipvh2uycpvL0kP0hT34tDaHRAeXPgMUoeYPbetzIBX2rICSSCE9XFq
DydrDUhyLXE9dGpMy1eygDBssYCDve3XMxPWnLaOkgH5UgNifRT8fOBxIe5jlOQ0
E14bEYX7XzRGPrZe9BKmsXVCaNQt93gVvKNnT1yJ83NRlJTuA2whK3HRSLwkcemp
oAAtY6h1rLt99MYUXrT0N04/p1TapjIL4fXIstMWU+vCud+GSqZwBmZzH7EEikgQ
LZLfyk+ct0aH/+qVJ6EDXcKtqAFJnoH1LwbAW5tn1QwKkFeXa0d67tCEWdoZhTA+
UqtaA9ddFsrjOhNkBhoeOg2adTjXG4Q0TEdVXXXETBn3AUH2sf0zI+OQtM2oev9n
j46mECNtUJgqH86wVk2I5B/lYF9FAo+e9D2rqd5k6EaOn6faNXstedhOsIJWxKIc
mVSMwVzNh128kO2So6/aU3OnbC3Er0VY7ZRH2815/7PvVUfjMEVGRCHDtwesGC7a
T1Vhgs0vCadv4/VLDz5T2UZm63cjAmHFgyF0ednVWla6ZA5fVtC4VPnIREjrdpYv
lfT4IKdsaBdvVG38dBOyW+P48+VO4LQ2zTRvM4+nviEVAJljb+kJvfTe9mx9O7Or
uK2+30zeIrC5gzH83ZGwBHgznBZWKwxk8OWtoLn7K+ms/r4ViAz9Fwq4H+QcVzvv
7MoYmSKq6n5DRJCMGSC5g+16qoNzq4zmSZTSWdkhFw9kvOnaCAUtIZAIMoUCFTFu
o1a97DdWT4VeRcJgtGmnD3u9GmTwuiJgumm8/EQGE8NllXWXrjPmFQW36dsKI0lx
0JpRUBImVOsICap9lJpZkRTKenEgLbugOtMWbqijzUEwtwF3UrA2TWYc1SXaRi9w
jTU0smALNNY+vCbDvpWzAJEP+aSvWlekK4Z8xJqgdN3D4LGpU2dEa2uHgqdA4/n5
Xt/1tWXH+F5bMgqqz1N27l5AMUMaHdo1MVEisLS5OMUv5saEWchzA2XABq9GW624
VUTv9zLYXH0c38wmRjg9dHsuYuM8a3dxxlCPAr4nOjC5xON74rNftIZrd7fY+wg9
a3/XF9YJHpze31s10YYV8BO4dHPFr/CuMydFbQynXx5oaFNkE03lr+2KJ7Rrw8sR
oe5mbE90f0Hypqu0LTmfj7wh9zBaMgu64gmf9AnGn2Lwy/aGuOb6lDYH0HEna7n1
dBND9a0M/jtMzBgIbBkH/DnAmOHqqId3vKKlHC/TIKWM7A6lGWr3fz5jAtjO57NB
H6JGqTFhJiyn1uHPbzQx6IYVaAlwwA7r+fsn0CI6Ks+xZAtYfyTpqx2z3bYwh+yg
hO6kryNfQyOZNPf3YJu/oo8MJPjl0VXA+rvfh63x/d1PwhDe/BlTpt87iQI8JxsF
LOhPyEiuyV/Gv2YuGhMF3DqIeQlQtyeGjXPFMl7u6M0IIa+pcnykg5WuWn4Iap2H
rz4hiAE8+pKkLNjsDTWdf3bWgNPp6aaGKY4MkA63/vnPkyVGy0fLYFeU3xMYT3jg
U3QmMo/5UgzUf4U2cx/x+7MrqIYDukXXvEToat+CH44BVsvW9j/+8H+569+yAaAR
DgcQNLZaGu5W+7fzqOGxlzfoCPcKqvGZzClMML6D7W/6GmYQkubg0oYMscFXz9+6
UZLrJzzoCR1ubPauVOkZeGBGFvNaK6xDIOWBam115/cZQqIFHHfVGUS18CpmK0gt
nIbiGJZtKIdzj+K/uaF5vQPZD/0KnJWK4m8FUJnQlZNqMWY5oIiW1ZJz5PVZt6L7
3FM9S65WrJdx+6zeSvtLxGjm3sRFv8Z99WYbBRjKUsoGBPPcPoVzlbP9N4fVn81N
5aFsH+1PNp3yC5reoh72rrqTRYVnrXA93sRHVotthAw+8I4tEaeTlbw4FuTXUeE4
RzgxjbG+b4r+xGGrST6L/W4Qa1nJqZlDhw7w1X73HlarFiQtC3GsBSVTSLiC+P2y
27nWfYfp7+Ke4Gu9kEfbV+ASzb9XrDc1ce2MVuMN7hnH95m5dBwE8J+Jg6wg9Otn
17XeCz0EP3+tbYeKmoT6lF/87V0A2RU9IyGgYs0Tua3EbosD0Y15oB6xAht7CTLt
j3MDZlAl0TBGb/N1ENjvPdnKeaj2NBF3d884auKUKE3rlW1dMv8jRQ81x2hOLukr
pLS6Dm+RO411cFVBKVJUMU378aTrlwodH3XV4I/Fypa5dlQ7QuxlPzxmcKjYIAf7
bC/BnPAbl5OJude17UUifB2fcv76xy5+YmaxbUmDr75qMuKJc7vxFwtsl5Zl8fRN
sIMmxiaxKt7zOlXUAvFwBxc18foDOWmFQse0kT5d798IHsuo4EGRWcQQmEqhqoCF
3O6m+lsNHUzSQL8jH4wuSooMVnRXe+KG1u+QUKfbmj0HUVdMm6yxXjomNZ+RddCS
Nnuo9ptYEhTRA2V97+rvT+mXHm3uSJ8A/UxssZa2SjY0uB89Z8A2FBsgnm1TgJrN
JH0ljI9emBz/aXWVbgbueohZLYSLC4HyDbcJ5honB+mXvywyMCIEIMLLEIs9VKqB
H8DrmOfR+7L2DTLTJpghFZzlixno8NWjsOnyzwDILY5h6nzKFkPksj+z40RHpyC4
1OukSIVs11iVjWgO5/4BDGb5X+WSs7kvhK8hbcRHqoAkg6IcTttfEfCll+I7YE2c
UoN6ecdHH8agh5DTTRE4kBCO737/4FJVgXUnp07AJHGSHzWRZVWp6vDXksUkN0F4
t+jFu4xrFQL4OLWkBtZDQA0Dp/d9PESIScWiBphVaazU/18TXByr0WrF5MbS6gYE
V/rklGgDXYf058OeqFeh01AKiFDKSbqO22bXrnaA0ttgEXVSMPla7Jkqkh6zlLWE
vadfjySvDKDDaPK4zeHwwGhsOyeeT2hD9nGGX77sDQSwGBuu403VNP0jMCy9DUyU
k5IjF9C/UzswaawWV1lg5BtGvO0KmUSfGp/B72YFmJoUgH2V7loBEIEweCt85F0n
msLj5yg3Rm/G4Htr7jDa/IPZU46tGbgI6nntCsZkJkrFlxq6iylipXHofQwamMN8
oKKhpwbsLLuanAz6mw9PTMRFumhF2LhtGt0bewY9jE52aR42udJz1BjYaBeshceS
ERwBXnBin80IPhvWhOllbJowKzoq8GxIw0ivuckoMk/WuVt7d3+fHDKGytTf5zXs
mfjA/zYAVQEFPy6ua5twut+Ap3uynz4/vm4hgfL6PVW+fEKhyNT1XbQ7vkt+kOtr
JYK4+AxLtASK8vmwpzREPUibK66RBi5+FPRWPyvFPdW9iZzIbLIQDZMxo4gvxAAG
lgEZoTwozLO9BFSKXQzGf2E3v1mc8HY9OIkgPiIDHui3Lnz98Hyea2rdI+9yIEIP
ryZMph1q1JLW+nSvcOInG93gMEu3+KhD84K0ykzcy+albplH4ITyXr3b0M2gAhIe
pnOZ7pZsWpbyuUY7050wbK1oI8p0N7+7t0xEBGtNeGsbyc5HDEDRKQ2MQY5DM/QM
l1SxpuKrCzQ7gjdb0tm6WXRjfl4DIW9MkS9vltSYTtyo1HL7eCBfpPm6HOrIMSU7
BJlj+a6YZl/xFnJ1zGvN5i07hvFIEgmexU60oweaF+oii9vmEn4Nigvv3KBJL17Z
yGue3QX1FxKq7feUJRzNrcApRkADayi2p4WtPYKWnm0EvkD0AYWURYXQk/VYdHy4
e3ty8orp+41OgUnD8W+ongoIQaUeGQj1mIRVbv6+1AXpo5hc6yzhOc771y+HBkkz
5eJNlJC7P45PnWWpSt9uc/kniOXxXY/hk46+9va3ZIT7L+RaYPyr47QIWVx/mcqb
V/kHyQCj6c7ZYHwrhKDB0t9u5w/UFMelX5kGYJZpzam2gsrDpopShBBUNnGQVvfr
nQP2BNtKQudVGc1VRwQbpKic2+yzldjQUXDc/VDhwGF7GCABHjVAbLvdjV7+Rt1x
GBT1NXWalqLMtPpqrwo2tVVs/ZuEkKTQPA3076me+Hklwue5vKUSdxjkbb+MoNyq
rFUQ1y3JsEuJFPMn+CN0ro13r+PLH3d5WjIU877PMiXXMQjgINUw2NgBZXCvbQkW
4calBV9B8BhHXv59dMOEFx344HhQggNEfOI75HP6LkbCQJl/HZpCnzFFceBVMvEv
0J3IMJRLZpqKutQ+U4eeSYFgNErCRqmbfbKhRB5q+bieLaeY1wErl7+izvByUzNB
IhAD5LGqAX0PxpUjbFXef8i+2j+lNXFoBDDuoeX741t9d6PS8QnyjxNpWRmiXrUG
hvC/1Ot1sTKvAT/hDDvNpn/NOH6bayz4SbT1+adWTrXKo0J58lxn89T7WKpYmUnU
WrKYuK9AgwtAeFFhk2YVxtEB4dqogDqReQwRwJcm59QDvSKJLZXjdXB8i8KDh5q9
oqKO9I2SjJeJ/r7nisCn/k8/iIDGtP9B5/Un9if7RmH7Dvjjt0tlrnIR4AeZtZDO
He+j8L3LRKqU5IHsNXulMgTqLua2m5Sf1JBzeM1IEcleMxFGwZC5dgJ/9YE+SIsi
dYPGw/kRtS6bPQoTY2JuQxHK4ISYEbOMIShTxaDehlgYCzAsURirMWqJhdKgLQG8
F1t5HIjP2IMsX40GBsu6mkboFy6WNkj3p+dUrilh3+PmbGO7s1Ns7x6BDERSZOIh
Z1506KRH9lFLCwGsTbtYLU/OBwlPHjwOQiuHyj/+sV5l3H7o8tECoqZOvKLUden+
c+dDZ3ZwR4IcP1hgAegEAmj2jeLC6zQsO0gk7VMhEKWqQqsXOsokrLNX7UzPi0vh
pd7xEq4zfQBGTLlTZG0fvIXIStiNHEyhrgLFle6gk/jeoj+cjzfP0H4D7HoVBtH/
MLIDNfJs3hzi+UYO9fSnqryC3Snrh0ca2XowqwuiG3sztN2awTMRa2C8Sft36B7h
R/bOkcrYKx90SFet3hFGz+nQMAgrasfbR8rr8EerQ+eUnRTgSlNDr50aFFfqC5qK
VwWyQ8e/jyX8PvDLjkrIbXHaSNofwn/K4j1W1gUr1By3x3W7c6zqfHr4qTgxWmlR
vpibPI/D22ykakACtZh4cfCKP3HfpVSXpLTl/SzRqverN3eQxCe2WGP4azMq2GXl
FyObKw4rQ6TczkjQQ0uOtgLh1Xu8H9B/zLfW5x8FTMse8Uys89bHch77GU6bAj7H
EOH6xIMg7BAnHsQKq5p4faBlm3Y+BLMoO/nqoLX55WuwbhooEe7zhb0D5olGRg+t
1skGFkgwzDMxDx6MkCrYaERcQpJPev39ZKsQ2QJYX9PST7QEmGqxBAVbuol/T9Os
h7s/W171IDyUMw6mMUgjQiVd3iY+aZjgjhi787Y0ans/tKhLV3T4KW1HURB5eF6T
YUGsXOfBpCKIjVChsZWZSh/QHx2rFDUVFdyFpTfYfH1UCPGWY/sr8U9ZVd9UTCvI
4sXgILoNZbIHjF2CzRu9rfKxXheN/o1sB6m9wzByp4cejsRcS4Mny0RKMPCRNBK5
l5xrbkWLlfqsw1kQZ/9FuOdXc9HJ2t6WsOy2jnmJKgzoIz6ffk79ZSjYgsqP/WQn
wyOTcYzEpC9Xeea1PqfqJOlZJARGdYf3IEvq1SRPFvgARVIXeVq9pwS4wRIB0eiH
GyU9X14ChU834oCJQktX+PWS7JsVH8YX4l8tM/Ix2px7eO/O6M08E5yae9zoS7Ac
NWxoViF3FB4dJHntWWyO3qrDkRXjEmiWqUfcugUhS3CBP1/6hwfmu0twUp12/u4V
aMI0f6ALlfX4wEGm6Bo34DfFMU22ZN6LLq1rbgo8nxT5TWr14kalaKUVFdJQxkb9
Tm6YM65ausljH5QWG+iL/WYz3Bh8mvSHXmw/xA50KbFvxiAHuIZd6XcuOsb/qkid
5H0L/x1loFGAEyNx2hJ8EJT1T7cMa9gB8VJrDLxnl3AvEjky2FHgSHg55zTn4RtD
rmIZKQzpB+n2/nu2trMjSNK6M+no1St3/duYWY4waVofL4InO6OtzInDIT+xaRQ+
q5cVI5pIA9cW9LhHYme1TiCKZ/nC5BmoblwPgSQ0R4KxwuiSxO+BqdlpcGyDQi70
s+BZ8pj94trwse4auM52sUgnbjvn8H+1fpjxX1M2wwF9v47H7D23zRJhnu0iSpCu
8JgyR/gOvi0l4TZPXygFP83bc5mQ9lZdOYnlZ2zE7NtNNG6yBO7d5Oou4pW2Asz4
PnMnqv1WdPIdJsi3fp1heh336LRiDrhkhcg65key6YOh73yqnZNfjkizc6K6bsom
hiBw9hDZ75DG7TkV158BeUarWBtFYIiqBV0TDHvVhshK964dDjG1TUVzswPUD3yv
iWRog9oecqEgR3lnwTjEE9nBHLHMe8RRtRBObXVX2Kqg1C6YItoexXwLA8uFrLWK
zQtEzIBUFlqHYXUof2sPAMefjWvNE3kuygzoIjhV0DJiPGtJCzV+Wwv21Y6IrOr7
ZfWbLJWsOdh2uvuz6S75ijMDJoT1fz10kDbQzm5ZCoFrYCv0HSyrn1UDp/vNmdhU
baKdE0icEQ1tEcHs6g9NBPyd1CO9x8k8t11E7nhDOil00TioPqmhugUYoV62nC6p
POjdH7sQdP+UiSO3bP9VcndES0nX6eUmgTyJ9NRfVApx8DqwXwFE9fm/4MDwQgbE
CH7jGPyTp9CF/3bRcIx+CMpy4vcF2toC0ky08IUMLx74g8y8Uxi8ljvlHpdzd8P3
vtTM0g6GYlTlt4lOP+2CwikVm1AQxZorlnwgjtxoPgHQ4vQJuPN9cPKJWbmZiD3v
W86w8v9hDHZaw5AKZdg2jN0VY+joDFysWP4MXe0uvaKvn/eJWGjgotaSWa2twFxu
ag8CImejZVAj2Bq8mbCmhNaylrI8+nu6Pu1rCrJUtQ8ZjhKgn+RWPSvhPwu6M3+a
rMvPSmhjFjdgFeW90ASvLd2tjqRqx20fKCFJ8NpeyGPAaSTm8w7Hitxhdyrf7tqB
Eq6amzj9+yi23dD6KzFoHk9k7ekqF+lJ5JwOf2HuYZAzUU9vS4rOHibXa7o+4MFV
U7pxVhR3w4ydaLcI7ZdYq0bb2lww/21h/WkFEzmtqNB2YCxYj/lISYGVHWiqLW9n
/O54IfEURObBAcVAUGwdnj+PUrUMKqk1jaGf7jmaDFsj+69GnYuvG/nfJfyiG1fw
gHil0S4unbHF4tpnnYL4ZoG5uRvbK5TrckFk2nyn5N78qQpLlGQMfUrigDfWJLD+
TEUjp/NF9WJGefefGIx7IuiBsqdXQunF/D/StaamAzTXoVHiCH1zesAinEUGJ3+X
fY0v+hF0lfd4HXglGDRq3UtQGDi8KWlN7pKYZ8eK/3K+4fk4kuvDNaFCVS84PGIP
1ziOj59iCbzWrauSrkFWveg/wZCpZcrAMdcnrDIUJ6oC6f8t8r8g13PCWJysHQiZ
wMHUL0Ymcyzc8jVzzk/jOkFU1O9kcF1fOjUMD62HcCpQH1BvOpMhiNUbrAAaDEUu
KZgk5PJue6d49T41davX56aTCFhN+2NgIgj7h1OBAkktsPscrqbd9EqkoyyNKSxl
Oqx+5uBbA7XU6UV2nrzrtD8PmNsTG8q/1gEBnBS057EsnPMgRHie/TWIgOSrbiAN
4I0zTnE9Ec+ZZqjW6YQ5kPLfePbxnBzUKPN2OfD7SonIhdTBhebEK8qloU5k1eVr
CS+ccnplSCE2wVkYnV2VV0oY3XM8EaGJ4iNLC/rvS4aPD7Wu/sWKeZIBbSjhocZo
98xqgre6Z27Gn6tbje0kTIxGsoZ52jf1IrXZ/29wMg4WjWe9d6d4qm8IRDO/4Qb5
a99fZzTTysr8LneZ4k59YejDXPTsduBZP6leEL0KXjCYX9Sw1h3ImGUy76WyQps6
to/9QCAaNOKHyGRxN19LO5Ye36nTfcjH8Kf62Tj1uGcrnDhItiSQICU1ZL8BQM+w
Y08ejJmXQaekZTpYtnGadOpdM/qcAf1Y90sXr41nMrbdJxPlIYP5JVkOXxy9zLUq
Q8RzMBHvIPY0MOlTcXovY3kvTY7KymjXwhFfGFgBjPBY53rUBjYg0QOgfUX3Mhe/
IAhUZmPPhDlweQJID8U3lvGJuWrrDviYalAlXLLM06w5VNDXYVOhu6w+VYKHit+p
Nxm8agfvixh/fXOmKCQVCEErnnDSHYaQ3M1tDpw0bNeDFjtBzpYlSZ8r7Nz79hbu
QHG9lLwTyfkPgs24JotFnYnSxmUmQD2jpJ476LXvo2p5T0nX/0K+SP8l48ssTLp4
q8U8wzUcwjd/TiyBh2E9qm3qzplFhcqGk6rQ+8FvIjLW9rn0QfKCVGer1FHBYzoB
y2rTLKm9oWbmsFBsjRAo9zZAyxd0e3x8RS0+nnJujNQ+n6vUQSDhAmtPCHNVj8po
WOJPc1vhP2wrVkYOfOhvJ9+/yFEswvEzWElwYfV+NxMN/Eb+x2v/gP3A+1tPI8DB
5eYrzubQ+2PVkLTE1KGkCqTJQjB8HzOrKNdkgOQDNP8w1owbLfREwpmzNjSB2aAV
lYnW10gztr8KuPXyYLPuwJCr4e6ulieW//SzgAc8thROybxlgcREtLbjfiiJjP0K
mLMBBtW21+FsZeo7xHJQ28sROoGdprmWFZZXQCcQXCPls3T3BMeriayRcQETyTzR
SYkQblG/vBTPla+bWshkOqpusL2Tbu8eO0n6RIwg3bs8XiDe3uNbzsstms0/Y4+H
xySoziRuPlkclCRwbaXuZuHahCDGFtzoX42ItSg9abhtmsO38Wy21vIOFPZwDuBO
xLxfEL6np530LKp4dl/9T3xq2vqy2ZwyrPoYh7RQBamxAHCK/Na0xYZKbXmSDR+Z
J5zpHozQhRA1aFfGrlUESLMorT9nrt/NV1GxgtO0DDVUQGDRiixuYBqSBN0LXhNI
A3gmceoGyca2Aea08lAkxml1d376EYEShjobBqEBYliDjeW1hyzhJjLDpdxmOonK
kF2yFf1gikaf8xyTzxSSFnuUidv+kfVwUo+2tZk9LgvwDyPlwzY5MA+aCDg3ZM0y
VhpON+KP6RYLBHgNGQO72lq7anDg2KKCcfuE2sDol+s6GuHCspENn6ym9BXgZnJm
SQeOOUxo5I68U9OnPFmWzMk40SV7Tn5dHIjobMvOMxRBUIXzyYZKNUmjTsNVm7So
3VOWavYYH95oafNBI3VITfkWHgTUFiWl9+KrzRf2fo5zNMc8iALvQNfA/Qi7ZV6g
O2k5lCx26W3+xvR4FlsmSlrqXTBFQKMheGH2CAgTxOsF9F+DxYWphsa7dmPIuYf4
V2SZzJs0J94S0i3nF5NFP3mKK19TP4eFvtauuL3sAg+RanuVz5LlOYFBUPqO7tOX
HD0OSPh+ruwkU698sp3dAYgqw3N6f6rqmn555awV5+C6ZOheP4fTAM2Lygh+MLKt
Kv19VaG116mBgC/ek+jmSfn577h1j+9+wyjvXD1PfmH/k3ppup+GXi7wQwNxPR3/
uTCV70inSJbgzwHdj8FuUTRVt31FbzKDMC9sdroTh0c4eL7XX2B56a/8PadPnDSS
SOkbdOmuJmjXaVircnOicUonz0MPSseb6FqKhxJKLVGqteruNBj18wAX3j9FEMm4
cAiTrMYxLY2GodWlCSjgnTfulEnSgNOBkqqHRdykRfdeaaQNnCurT+1UGnwWBRDN
xw0zfh/wSElsK/oupUGzAeXpcgmakacGJbbhPSHTIq40rwaZklZ77mXqDt2TWazF
7jOvF5XVATPHUJBoTrCvTFdfaq+jvyzIfQzOd52eWhjQpoVgEptMG2zH1/6AEcDm
5tl5xqAeZrfixkFObKuDeZzwLR9P8rCVnCK2SvLllrnXlOns1CTPb3XmNl7y6OpV
rOcuB6vm6PMHM7GAKq365StM//jv4D9pN6/FcKIwaWjaRyu7m89CXmbnQ7IaZzRb
VEmhaFf8TzH3fa3z4/SQr1f3nVsOS/5fmzv9sUZtIF3upgvcPMPczxT895TGRUn9
w90WXDRKhNPTqWFee/tvGCcxQIJ5YndvtoPVk4k9NdVaNQAaVpSzwj3myqSihww5
I14Bq4yFGhi2cwtsmC1PCtzDU3SEQoIrK0jEw9C29YR2CTKpcDn21dmMI32Vzvaz
xoAVbYafw59YRRUqI02qceTjT1HNj0TbG6FWriCB0LlEUuMuApvMROsZeSPfrjG3
WyijUWd12nJDbqhcrD+TRfF8mpBTeDjgFgOQ1H6u5PUxONFYAoMHZ5GtTvJVQnwn
BtDfqYLOB2r5WySSRy7DplzKqBugt34B5gQ5u6I9FOdHafMgTEpSuAb0vvZ+v1xK
o4ha4B9KpNd9zG5mpm9nuS7G//PXdFYe4lD3ZjFv8f4YyOO45jId9xGpgNRSvedY
2bbj4cCqq5rav+ocE0FHQkU3EAgLoYsHrxkqlo/ZfxiDOm6LGNshWe4JWNFBH0Jq
gI2i0glP5yChYFMZDtIMNx6gMCV5SswRtKVqeVphYEZbe5EgK6W41DjF2MCDZA6g
HEiexEQpv3rPJ5YSFFsa1jeOkaEfdmCmd2BykJM/mC4C/QFuLKILwFJzReE+4IAq
dwmf9VqDA1k1uTYxi+GA4m0YFo5oPfGFBtRKE01MXmii5xOm0a2MWWP1KYcPAADr
7fsik/HTa0C2Yn0CGwXKu+2jjyw4Li2qayh40CaffSdE2yeTtQU5PdbqfnKXIHkc
uRJLUDexiiAmM+IFZQu2zUUkf6iA/G3h6L2aD2q+b02RavuhWmzn1TaosfBWdtNx
D3ssjwuljdHClasyJSNQ1yRJdHT7jTKWV/CJd6Py+YL30QVZYuCJEye/jqjkD3Tv
uk5NOFfVy20a36cwngdW23CUrI0eWiK4iRbo6bYEZiP1KU064Sq5gkRlDqG24xuT
nmWgfPExGPCmpkMX7KeR4MIKFV8YV6/7A5gyTByysJjc5ZLrrY9BbTBn5kRdvJM8
lr1aEIudnvkyIc0AhkBY/kLJ0aB6a7Od8xD6YAww/L/FdF7Hz/1yNx6ITDIvwLF9
QxVH4w9NgWr4XCwgevh6vwKMWZECpNdenf59THrV9koU25bEJffVG3+ukoedJAT1
cld5NLt7+QLgUsDX56mI/MPW1ymtB+oas4MVKJMxR+YPwVto2vG8hvyBlqwqaTTv
8ycVJ1ZeLeQmOVhjrUJz/Q7qmb2RYxLsvbxTzfbMLShCVJ6OaQGQdU1wqlXCppxw
LrSATS39kw2Xm6V/Vf3sYEKG/Fq8Qlh0x2re3EZaZbYmQ8bG3T1XhA7jZLyOYgxG
+UXJMs/AyZHTsOmo2zXkPrCTs1OjBwzeuVa6uuns2+JJSPJhOgvW2ZFz8e2z3iTE
dJ0RPeSQllI+Kh2gASCCvr8Hr5JiheSvUWTlRDfpQqm/aNQK0oTm9ZAzvKw9jBR3
ALadHM001ALKv0tiqTtRh5Nz3eojdBMnb6nMnFrHydtJM1YXC0kHW2shoMvuxGNo
oWWAz0/qKn+ujUFNPvwF9f+Z7sSZfMDmFvgJFdE62EU8Ke3uK4t9sp0rii5Cqo2z
Dz77GxU2Mi079yOS6qV3oJjjaYPmY4Yy4zz9v1O9l6ommKuG8SbjCH9hErq5dHY1
GN5ECxPZcxtXVMn4YKsn2yO9BhwnM4aJUcLA0W9qSC/JSyP4tgA89akgpEdjQAR6
7elJZ0MCFSUGN5cNe9AFJHFNsTcpL8k52a0etWt2H9uIx8aOd+m7yjpIBw6zqdhh
vbylNE/LnoBS/1bhJUufn299lB0jhxHPlKvqLQDwrRy9zd7Oc2MLHpqXMTNrKPz1
bv47kbzwsT6UCw5Kh5DXll41xKiCSvNZWEySjGEEelWpb/ES9V+huml928NViokD
2mY6WHgNwloK1M+KiBpV2htTJlAeDwgXthMwlLseOssYiOpbfTWZgp7x2z8Hkc0b
UilL2OS89mU7J5KlJXQo96T5fLyFe15ycuylYQdd3CYeMm7ketFOopeTSU9R/t6I
ic/bTamNgcwv0Jy86HQFrKn8+LN9TJxsu/y5qssFVllFAFsu7hUnsflOi6h4gBYo
aQwKAQ1NTHo1eH1uRLlWyv4uW/RTtaj19Xn21SOIL35XMfC5xDeoo6KyGSey4Zln
Rh9luoDNbOeQ+yx/FJoYC+N0Y4PyyuNSvnh14z6EsV1bfRr8ddmKOmpkc9R2ChWf
R8PgJ+TdPEkIHl/8pMH4Z68ondvC9+4DhfMtXFOndhu0z+vLJ8Is7o59FjUbm3+o
beHMzLLTJ+OQ/3Rn6DNl8piuQUGOk6HfQH4m01IbMy8G6wLer9+sKgWYRR+LF8Jk
LP3z3ioqWYHSYhvg4ZQO/8HcP1/sg1SJ4tNWgsisuMVO921dPDQX/l5KS6lr5eSq
veKjzClH9Q38MAM2WraI4MmPnCfUtkkXHL0sQ6kn94EoxXUPtdTiErDoQtsYLKCo
siG5r0dITWqGMzRGGYp0vUK/LQdYRPXOWlVOlIjDBJ+jjf1ECPg4rky3LJ5iDFu/
60GCl2XVBn1UdAykEUIYbb3yeq9oRDBHYhofD2WxA75riQTFZLbprGDxIrfSF8WE
SH6dA7BCxkE/icEcMpUa1SVpYN3SR9+rwbVUfYGzcc8rRSq/88NpACvtQAS4RLJL
PvMLuV0wXJ8jBLc6rj8Hhrfv7xRK4MXGzI7IsFRcUmCWx5EHDIgdH5i02fVfisIX
xDDan5ILjETayAR8/SNXc4MOIrfAHghsMeTq9CpGcUGxteVz9tv5q6S/oEhpHSJT
HckYv0mQu3+caLb2oSWnoBB4Nh35yTkwZsyUPb46YZF/bzfiUZEtxQ4wyT03P+Bp
kab21XB1SGSwyR+98fz5O6ieBB2hZySyJ54qgX9qZPva5OCWfHK/TK7qyFMnZgSF
3Rzi0/ddj6c9c58thCDHFT4vjdB3LPQM4O4dmq2WFAo3yOZM5LyMMfXd7UzPMM8U
zyrbelFDAPEOHI+W3s4hvWaru1FgcL0gZJFGtOjuVZoxH7BU3Vc4pcMlIGLAI9oj
6xAPt+mljYcy3BLR720sp+rD2o+eBuQGusQOBuYxtHnQhUy0Z931TOLLZPfyqvOK
XMsKMeNMV1o3ohvmANX/bCQdxMzf8lKF7pwwtLRJAv5SD4drR/yMA1UCyACiyDWG
FoWVgUzqhQlD/NhEPEqM/4VbWZDyt7sLQ5Uol6cwDVwPjJeJeD/tlAnDoGZNKnMO
E9w3ofKU++6dhGQ3Yt08qMawc884QIpCnFXkgkLHvDyjnaOPvLQB2oUn06voh8aw
WJwEaU5i4tWbaGFRS/SfWRKSHm2mbc1ODDrQWbzcakt3iwpY5AMcDFYJ6YAuekTC
EE46QDRFpCQ75r67BKtACOxedC/v1CSX43w1IVnnEmG95jx1+8KgE5SoA/ZkY1k5
zR82xXSOhNlfl8HQxmBC8OIJ7vcX2MkXoFIIgSlYedYiMKT5ZkdvURwMgJ/78RnA
IlPA8PTs3oQiF7pznQLUd7DnCZEzd6CuLNsUWvc77a0tzjWdKd1QjHjhxJwZtzjN
RSwcKJwjV0iPGJVjKKQlRuqk/1a08V8u2PQnuFBcNN77GScosG4teZD7ZrW3Du2h
Uc8tXIBM4tWle1Rvbti4zVY7/0yqm2P0Ld5fBAl5rV7yq668k/qGIHaUZ7LNw8jR
p/Lo8MaOVxipMZDwJ3pfdAZtwbbpxoxOhr7aUCWwgtNAyPYU1/nUSqkiM3ww5Xl7
EkK97Rrgk3Tl1NF9CAtEDeDMZgi+j8sQtXJmSPdRxK+FH9L8aIFOa2+qu3KHAR1F
rrDLcSdwQhUISXEcfDiGVV6MoMZuS7j00u1OQyQtipsNxKTBA74nV1SaTPs1E+xj
juyk7m7gGYDMXah6KPyUGql09oGs0mGBnhOfp8yngZ6HtD61wAKhjS2mT+9yjatu
C36kf7rgRi7FVDmRgAli5Wypdv+L0dhLAO3R2QTjhNbDiMlv3Uqi+01AZIL5I8jw
zFjQfgxUdhj+6zgXbCrVUcqDJ1MOG4dqoATLIZ21odBr8IQQhc7najBhQ21inBO+
772T1eZ0wps5MmhAQg6/vtJPDKMQdB0HYMnQb7zHkJGcSwCX+jDVg4v5FkiE3mhy
ThbdYRX2M5ExyOUQZLbqqfV4Ks2jAfMBarp+uQAJiYvDhjJnM6I6pJ2XpMq4wGi/
FWljV0Bjb0r4+yGbyd5gSjyB3OQkI/HOt3bBh9zEp078zRJQ+qfOl7ROy43dFKrs
Ug8JEwTwZXXnGtnBQJ4oFYelS7HdtbXeckvNtGavYjorYIazj6yi+g/KVL/wLIY3
U1PwxKoBHXPhRknvNtcCmC4z7Zj5Ys3+svkiIAXlpJqvkXk6k6fJOuQ6bns1a6oD
vLWhPcfTmIral5E3hGj6JlZzUHYYEEpH/ScGZAuUlX4sCe5Zd2x2W9tchQRMMJ/d
lMhmzPHkO0KKYRpeT82H48qS1/22s0bstyzpYOoyoMXHPwbNbDW5xO5uKPa4GZP/
3DyVDEnnoGk0FmOJP65oVnA7SKXNMnxQ+Ito5JU80o/84Tpnbhh4g6wpIVo56f1u
NGP9y7MZ/ElNM0OusJv8mSgPrlAAFhv/hbg9k2YPGioS5jOFG8oeWlDEvOprGgv+
+KRmUZPL1ixfOHVFs213pQ7zFxU+AQsoOqYPFiGEAIoCc/fKNs9yYgpgIF+F4Kxp
Xt2HqrCBYsIqzlVZshHVegpFMfj1uDDPRpuks2NP1fQ3nmWyWm8E7+n7F0aVBWkE
p17AC4nSVWHnARHKd3cbq36LNq7P3+PQDWkpcOR7wimEnA/r6BPQTSIRgtGtx/WR
ZN6AX2RPA9SmiMiFiFg+ek6hOxAyLB7eRLuNjbI+nK2StgRM0YM+BbzmbvVe0uES
9xc1ZoA5A60KYuN+udtmXobyQQtZ2dPUOHcWb4RYhfgVbq13PUQiZ8yzVLfZw+ti
WrAn9aJ/BTdNTGH7hRESC8j4LZUovfn19wxmaDW0soynsZipDUsLHnrrldWoVC04
cmKFybtGSCCBcqcbGGdAzfgBgn7k7kx3WlHji5mwQuT12evkvtrh7iLXFGWEg21N
ZwHBDP5EpOxoBGqcQi6kDPe7bcRrjsjHSR7Iv9daLOl/AgFDYKUpq7gNk9dl/Tbo
AJFKPHGW4RqtmrWlq3t6QUZtI48Ru7CrxCI28HdkrVxJ92WJN0CpKGtiupP8XBMs
IdlIf75LirEbj3RPSG3KvxGIx0SeEmtEQNbqYkaPEc1dfcISlkRfwlmnUgeEtKwi
P+DYh1YjUTkrACQmro36pDHU6XqEOdhfrGhsPgnJJSebXgz/4MrjpN0EkE5HY0gF
xjKqMvxd3CBVyInRfNWZWJVaCghd+Fl0a5u7Sj8YWz9rfeBTARQ+1AcFzWQdpMJM
654WRiSRwqfC+/WxQbZ2apYF9948DnyRpNUJOOk175n5M1rI9w17Rdk5f3mDw3B2
aB/WDqTsjmCEaIFmCPLhZW1biCK60Q/sU7cpm6QEKOqiGy0vWh7kN5opAFq4R3mx
n7nXIZhzXfuVMcoX3/WREn8cnTJ9DFArK/qyfnbVsyhNT9VmL9aPQ4d1JR7YKroe
M1Rh6r04JWD2ysGmXxc6UoMCPzFEvoY+r9ZAs4PFx1+WSASQLHvR9QkDJ816N7Jd
WU5u0wuouLoGEN0t3pTLHzziuUAVr6F803udhTh7pe4UzZODqrQ00BrNeUNPV6A1
cFEm69EzAdt2QCYwv/LhoravZ3OfKyOpToHKzh7dw/t3+bvSLF9fen7lxrsl2ni/
qQmzRxer28cQvDs4P2PnEQIalXmuKTtvPoFvadT4n17yzj+0V3Jdg4tGWlVtMLb7
Mw8/5AVC2Dwer/R7iZtzj6bEI8Ww8OZBgQS55NZLi2wi4Eu8ouNQWrg/Ru+UIKpS
K9mrJs4UxQRNmuP35CLG3nOjKqS2DKvXEmRD4kCN8cNA4x6CGFDiVyj/nft0N2AX
1gqJl1uWb3HSkI+VAWmu0TVZmM9PVQsU4c92DT4okm0znkVRjGN552kTg8a4oDjz
sSL3R07/f8aa1GLiRhzTUdpgkQBkwUCukP+kMsLq4j8OYuWFHl2BlDqsSv0tJWDk
FK1F57T6iQeNXHC/f2oeAB0x/J+A5oR/9UHIJ1DKObAHN4SUzhnmqWRpPPPqqOT4
DLMjYXLIJZgFsSMHUhAgZrBTnYtGBoGb2xyIxvQhDMMqEdIf/jf+H//PFRtJwGWA
24DKgUjbSAegTbllgVKaQL4hBIeeKFMfZ8qbSB+S7dI4kp14LCbMIPXUNFWvZsZ0
13ClE486HxVENoiY4qANGNRxKVrUN10H//AyEzZA1Zz9oHxIFYZIWXGdsr4noi1w
7lFadeBxlYwf33Fl2Wp/Fl2JUDe+62uH/CSGsAOEwtnqoBuTpsuEeHcHwZxjc1iJ
yxAyHPyvUHukBsEpG7Pv/OtMKi6qqvnxzNAARrJ+2Z4yrvmUYGT+qD6cFr15AqYN
UojExbawjW0kTWBjlNE7qPJu8zHkBtwVAZCXe9MiZLHPB002hJMAwZq1so7CuEvw
bCIA4yDrw353RlJbMehbKOUng4wRhY4vioXPWvi3oC8sSvZkE98FNBKDDMMBw699
SkMsDgr/AseAQHHHiqp5gRee8sz0wPPBomQpEGSC3xkwqCrtRpY/tVNyJQCcz3FG
uvpOBj8+JaBGlmbMFZ73izLtcUL7zSr9PcfWu/lVZpJm/A/fa1d6X1JU3w5lislm
mcMH5C+9PXJqWlYXlPcIMYnUAb7CWE2d0x90r0jLqx54ZNUJ3ltwskl4MaLCwHtV
YxgwlfYw8W2/jvxMndl7MiUHzopTFMXcQljDq/NcmCpuj9gQ60y1FXRruN0i+xb2
7a3f9NS0VDdScQc4RknatHy4m4yATL6vS5M6TRgCX1tH4Qahe80UBSVDIHhyHCwk
IdEh+PfKdKsBnwOU5uRXSXaqK3F6PNCM27aUYv26rRlnZe66MqDosaHKgck5wkdl
8N+wg+i5Gj4nHfe4dsmZtyMdUQt2CkTyb6z6GulGo2WS+52wtKJ1PrVQEghNh8ft
KRj/hY0P3NHqkqAAd38KC6pnSCAysuxrtk8b78Ky3ka3VLVLsW9Kjpe6Bqm7Ozjr
ztKtLlqIdi3HajYPsbD1/ncmQB4EYlVg9Mxr+wLyj9K1rTrZmgXpIHVd+/RZ53uu
gix6fXb+QJD3ieYFSo/t6JWkBNliic7xqsMFedIoglN0cg8TLV7+h9xBz0BBUa4c
6BVq3LgATBW5hpcYQR2j3OR7EHVT/8LAYElyPNEPlqo3MHy/sUirdeJJXuqBKtDp
DNETbu4KTAfgcmsJpBvbtC4hSZDK9Z/vJdW87XLdf5nbxZZN6aHHFYQOzMCsOBQP
G/HUzXjmfP5h14GADyfr/+CipVOdpzWKuCHop88PMjhUjLJeTlspDmh5tbPrkN+q
4Z8lC+OH8dNkahnKM9dVJV7sZJFqVbI+CTrLsgZtb0SVAr14usD4ZY8ffq/25XST
xQFnh4lbQ0y4AIEuIQPgXE/gmSl8OUOmA/ur73jFhdtfxd9DS5bUrd3CTvMCNX5K
99cHaChqCqapgN4yf0F8x4L5b92GXXBZCS8mKehLT/tmqdyG2SS/1tahZv0q7RpD
9PxV7mtEalUVDs+q+e1fTG6INzAS8Xpz/OahQVi/KehzdPVgeM8S522UEdUHUpW5
4XSKOHbLo+hDc1X1uoU63dkgGjzk6pSLUMYlbP3U46wmms6GemBVSqrBAAG7uFMG
ys9WOfmI5FxITBvjL5FAH3sUKTHvXYeyO+QzIiXb449cCjPOMrpkgT5U5HnOxiSM
NAeOp8yKHunQC1QteWdZwMYQfBnqNTeqDUiG1YGCH8IGLze8wzzxOVhGprvhTOxF
xI8GL4slmFYc99EODx3QDVHguIBKMw53JErEL3+19Jif+hTDNqs5RgBa85GR7wkE
5yqQ8zN4TmLqeCKDLq1aCX4zF2k7H1jVg8zOfOoat9UBbeZLyWfzlz/WSZUw0YdR
+I1PN0WBhUpSZfSNBCBovv2jOnSlIag5ivcCRnQaKVXjtJOOQhsYq9CN1C5qNlWj
8vo6wIgWo67lwZkj97yXeQP+kF9aJIeFT/2cGzIzvJZwFihLxa+yjlatvhml7LE6
htffSrE2zFPNiODmjkpRSPVVobmg2d9Yr5IyfkVyjyFP/NGa+3TcF8T1Tg7Fe8Z9
B7CAD2H4CqXS2K6jh7+El8w63x7w5ISNfUm3VVgrQCO9r/EHd6t17d70uN5OScmK
JYOevZtt+UZ9+YEzPdWV7whCIZ+04pGgt2TtHLILLEG7oYWREwMGfDsgf1B8e4E9
G8lBnXPAnL6iBa9d95Z9uKa92+/vtJu/TKRzTn7Nt0qetjlppRXLPkhw06a+nOiS
b0tILvrK/4TP9fksaKmoROq3SdMAXKkq4GnyrlmtIW8hjZU1m4zXxVP/s7Eo95Kb
Lk0qTlj1TT9pwx2OjaLTciT0o+q6yTH7w82QMTf9KE/Do231ToDrBKwtOA1diOxP
7ofCt8WIW2n3QenJUdGI9+dDqZdYpBaiTxfZ0WXkZ0mnxoEghcJm+ZU15vPLMYoQ
euML0x+1aHZ7US+95rWTdRF3RxrNpvL3KROFv7z/2YGrqbRt1Zwr8MHNiXQs03a2
phWPc2UXpTVn0xXKcuUImnafIzA9zO389+mPFv2MRVd+UwYnD3zevfbXV3NpLe7T
YaFFtZdrmhDgod5xcUBt1YkaD5dCjduCxEP0WQVKGXVmyJh+ti1aS0rWssp3RCfx
nVidjdlsNwXc3YsJmzHD9Z8BnF7fr2LYNQuPiFQyFDqrpMIJebUXAeO6/1MwPiwv
HgOWK3lTzyDjy0KzukElTpaFYQiunECF7TigXNSX4+Ee+cCOrfpmhVKDSETn9T2Z
hWcIMCdK5z/CUQhnAXcIE2gLwH9fOfU4TKRIhPFOxIjSNzjSLNmSmLUohYeqFJ5E
xbCbWoX507zB0+RLi6n2d0ji4TVtYvF6gZXQugLB4Nv/ni6zIUsQP0LTciCLhJJL
0LsNcNnue3586+TihPEAqq5iLxEVYQZcczkK7cuczEQOdR0MTha8vV94uAUz30b1
nXROmmrtbBrrNKXvu8wnR1Xo3A0eytKFIr1qQbj87aLV2vUupXm2/NxXem2kC87j
H0pEMDtW0yhJGzrOQueX0GQzcdTL+x9IQsie0JEfbbECoUCnYGADXOAI/YFmh7Ib
3EfRILDuZ1GEFTn+AmxNiz1PDL9fNcbeiHahCsTdpBnuA6inUNZKda6hBq441rss
D8UY41b9EA96ZN+gTpJEIAtU5po1evgR1zdDH6fXOLi8UEeM060t17GWTQ8YAEBq
spGtFfoqePSr51mui8QLJcvIGFzm1Intg2ExXE/ONmhksPW1LgywF3xPbmyfLJMF
FQA6miXdg0CQJn+ME0TdP/fxY1yiXvRLG/sUYeUoPywCUYzdM4TxzbwNr3BMVJdD
6h3K7434CzN3MOSFmh1W6OeYio6zx5E2S43qD7ENwqeNAzPIIby3xgjdhPXGinzP
uyZ3zTG/DQdth6nZP0GehWIKXMx96f4S7/TL0osy761zvfMtBNQIFhpnbVjH88to
DqOs4V7vfKC/yHA5k+5cnRd3nEiLMJ8Vb5LZxYgT0sAEkPjZ15TrPK4yg6h7H7ue
gp70fTA2VNjp1wPCcmtAZjPcBIWzKIGUzXQf3GPeVBV7BxZS9ySjvoSpu4TMhsEd
QOWY4+xJ6+0+y9onB1kOM365LwEOhLkRdo0ELcjvsTCJcPpKvz/a4uDAv1S8dfQl
Kdnlr5wB5xewy3Wk/CWuoO6BMg4BGOjpCnvQqDUc8zzM0De81fEPswsva+klj2Sm
B10l4bihVv0pdGdvLExy+BWvlzZOBq902X2DwmD3wlaNBF96aNKstKLWY7QpNilx
SHwg6JEH2ZlkAtoqawoF6eAQwiqYxFLZ46AbNjjPGPJX5OV7qf73PmDDvxqFAwUZ
DcMdi9eBR5Z8a+dFJvZhpobOTTKhGBA3JHEtsLpmhV2KcPMrdeClwvqSHvWas+UG
3t2pjFwJxR23JasEW5uUxm/A6RymtzW2R+pRhzdIYepXC9SenvT+4UCFy3FsmY/b
4s1eJJxm+dT7DZGdBqnp7hQbr0grTntoOdF0onm/TMrYf6H6TuibWJ6YCF3C9w/h
dXokDi5I2mntMxXEM9nSmnZgD0B+xQYkunoWTy7Q3s5zPxRslropFcLjj6DhUBJE
7mNNgDBIgxXrWKe8qhB6Biuysv8cQUudwBl82D0LGpLmc6toJ8IsbtQI0UUGsPGQ
InbL7i518VNvPoySFCYPExzsPNqsG8TPxfuv6a7nlye2JvDPwQM7hvoNEl4iSZql
I/74Qv+LwoRE+UljHV3VtQY8Wz2VECtXUvXaj4MqqbRUv38HLTfn2hcZkEEUv2xN
3rYOl8EZmOCMhKYZm2RI8v3rbHi4td8H3NyPklElDzkHd+5XtIdaaP19UXpclUbH
lHhy9b/pn4poF3LaAl3nKZT/4iMBHb3QU6dRw3eGVyDx/wKivl9gZmcA14RxeGU/
CXqtBWC6Wv1iGYQUVrSI790NCft3kYdB68lzfYE9ECeXQvM0wl7J3zZYrZFCll98
oxflVCZaq9dzoHnq5NLo4xg7lgseIbvItIDGiCxfZeVHHcs4RpBL7jomNcs2nb/v
Hwm3Uyc4bidogSmC9oLn8OksAwpY3ETXnmT1GKfEWxLgYMCS1I60pgz2eHtGhXGL
chA15yZuDHRJYyaaaAO4v2Da3nDG6cPVKHe0jhu2K6mwvh4q0n+Af7PAamJ7T5rz
2YKIPaBVSKDMFDysuP+02X9N5Wtn81wVQpWccD6MHekKd5ZZopxI8D6gAokMVu1J
jiIzX8p8NTF2Kqo7Wyhey4yH7+wxna/O1mXTxXxjM6rVPf9vEH75hWvfESbzJynk
Sv6AyD1njuCT6OXNVtMtPPwbw9UiYXqa+x1MGF6d0RybVKA5tXW/9CrS7vOnFsXz
rIWn21KbM7W7ng66kxJ7/GLQk/gKHmAThS9JA+F3jfS7+TaFnMVGfxRcSvpyhib+
EQvqnPJhoQf8O7fTbt5JO7TPpgqhVTuTH0Z9FbELtMQH26daNk3AP+gedrXIZYIQ
81I0GuvM1b9oPFyU3zYanhDqXlCNWUKKA7H/4UWb+r4kd1Wh+C/gxLPetQ8zCGlG
xNOK6E8LZb+F7Q/B5evjyLNWoy+3aylojW+mN4GY0IED/FNFCumZJwJLQkWWa3Bj
KQeU/yVOkrde61DnH/ltUhDQJwu7AsjUd1sFlG7OYuJ8j0/tFkcJSm9UauJixDga
lIcYHwRco1B0yUNA2139AYgj2zud1/BEAM7QYjua+ziMEYlnG8QMQC/uImW6PlRh
Aq35G1Sflso3CIlTFZJMoG53Ll/1HAgQtQU2QfV0hwNPqN5NcNf54N75u/UyeipC
qp0XD59x6mkT/uRM8Me2NFNkdeezIiRwfVE31zFovAjzQFtM0A8MDuTJdzEdZYb3
YA3IxfrnDPbtSyUq2UOzyTkcPsU5s+GHHPr2WKLxP9VgRInE0QILyNkMEf9D5phU
DVzYAROzXiLRv8wzpYyuVv4L2lgTZcsE8IDlWoSozazN7Mfm8WvHO7TS78s5uKtY
iESi8Clf9sVOQoXVnXZVLQ2cIUOzjSN8Vi/uMSy6uDNU0fDzGjuxIl6tQW8Cnm7g
9SHaPgP+HgLJjf9X9dF6DzLiDLVbOH6vfgMgZR6jtDhLuxHKsf4dJHUyHWUfSKMH
hsMnhy/L+3Nh0DrRPlT20sWeHYHMGO5k8erqWe7jSwNkZ1b0dOFNShEYEV3el5Vb
r79jDgdb3bJgN3Vr4oyMbY2HpnCQmKqfK8TwFHF6GsqTlOKzZ+nPuclXq8o5BbAo
3xpaQI1avgYJCa14+sbBRNcN7nv5q78hD47vlm++f9kXhzXtBkIiPv23N0T8u8a1
j6xCACmc5+yZENjojTs6LOA7hL0M/v5TKfe8o8thbTXhe2X58wzan09YFG6YOXDQ
dWEokdIs+A5SVC8+K1T1KLhOlG39JMWIkjz+Kx/tZmCACy6u2A8bWOSSEkiM+plw
iWgVYFuxoCF6IuuE8eEVyAkeuSbvG5Dj6Ir70swuO0T49cLHSZsCixYq0UK185UF
WnXNTa5CaPifghx7VEbqRoWXg3OMcGSO6s/HL3Y4Q17RTVbjl1aD/GGVslV+la/X
0rRwye/IsjUbRamcTxbUHss74ZV4XymsCztBQWUBTwDaVeYQ0xBT/V/p6xezDpoM
MqrZQNywO921j0xRZc/qhUdiL8O2T+R95ZPct8Uxs46EOVBhYB2YMxrYqMNNl+oE
v3jKhrhcqU3DJhgrBgNo8/AguVciP4dCnA5CvFL1VkBV36Mtn0UISbjSiMGHCwaa
YkeR1UR6tFMmnxb4WRLlamiP28sePbV/XmFKd8wG8e/6Lm+Ti6Rgg679AbhovWZq
pxZdWF7ExP06cIXuUT8r+ut9VbQoD2VSv0ixt2aE0fSAX9WshmdtR05m+PpQfzvO
laG1rFTjvpPb0QjFbn3Yn7N24kkMPmoUPJRxKbRFYOQTYrHsstrKrDPRwY/PFMEw
LjW3EYRlFhIYgb8aEZLq9DQT73mDvYt98rj2ZJeeBjhINCipfvvn5U7hNG2dDGi3
GMzjW9xTm+AOh3/3wXroeIxfpZy+ZeX2wn2ZEoZSgThQylb/zIYJr78DWHBCr4bB
dWDrl+auXPn4HeOsRgOf71vDOo0jNLRrqlz6ZviJBqZ2kRF4UEOfIm7R2PEtbBOr
W89NBeyfIyfFQhIjpjQm/hm/eNaMpaw+WBZeeL0DEyNHXvveRICOxzQbxSTdOBP1
UD4o+wUeV06JGq60SLpk2Uehi+KUy8rSG7HgldbWjCcCINWcRX9EFn2R6JkyT/Al
o8nJYU1dLJOn1BMz4zcDHwMas8HMWw2ZlSy8nBZEHu6mlOP6d3Pb5sFMiH1x2WLC
J45lGqJ0BIIkqMZpqZrq5/bw1mykx5oYmXwA+I7uuMbxRf9WNXUJgP60pxgoFOzk
TkHwQ8wBXQeZFXmk2H6a+i0CQAEWTKV7eEfM+HvCFiWl8wqQv1yw9acXA7pmtL20
PbID/MMb36TMtwf/qaB7steIBMZsMtqB71JdmAiLh/5pI9Rh7OINOdaBncT58rTr
HqE9o9uFWmvT1Qgyn7UoUsYULFtxGDPIIDolJ4B+hzUSryi0HtPfhOsuCO7ahQQ3
qdCq1G/7inJSnY8zotLzEeRs+GsEYbeANm+U15CFRDpnQZ8Fk/Xc4roOwxF5pfUr
RcoV9S0sRhtAmTA/IJ52grwZFXwvsIJuvNjNXqY8UgPZhM70dNMOVDLmAhApnkp4
VVsV+aSMu1yBe372gV31BymxPYRSWQzZoL91UWxs4DXghIVuqVFNN6V62jmvFiOo
ti+TahYU9v7HT1rAW9umGGQYi6H5IR8YRLd+JdRBjioYCDBVOZX98T7/5H3sni0v
y3NmS/cfdNGbXRDjNLnFyeUurfT077Jjk9evFS+NSGQIfJhYP/8iUh668Ihvop89
t5LPSLmC5jrQWJV6bQzoV8PnWogpLeM8H8NADdyh+bLTQNcV6yDdJtF33cvXFWBZ
X2rEjLiQ3BLEKH0kW480+BKhdfrur3ADSkvD5FaYPiV9Xc4AtFT12NpnYXh+myN5
6Pywu5mLuuYHhh3l/Fjw/7fryVRnik9NZz5J+dZTNWhZodiKM2i655KWjzSciAPu
K06n4XmvYFzqIeEgoGmhgHGsk0Sz2Q5Ty20aN1sHj8S0Dw85I89NX91aOxle8ADb
h46NzLRcT8ZF73XVRioQ7Dw3TtobOujB0SJi+buZmknQomhliwIYB9XXbKUffHls
XkMvEIRLv9voGZeAqvuAXXFdYI2jX7Ggo4aU01R05/pwJQFL8oFf92UEU6gw4IBv
jwnwpbaxpan/GV4TEih30+eYFv8sXoYiYXiuIGqC9GhknbtvpQEIPpYbwilh2dTv
tcBgmgTF5pDU2szaPdRa46kCb5iuaYnQ4jiM264z5Kx9UBf8a7WAlUCNAzeMN0S1
yBAcLhZIEPP7AdMpIgroDC9wvB4QIlKVyDRDKj4P+wWnlld8QM/MfvxSJMg3jhO2
JM0/al05J6C5Ik43aYIZM/8gCxOZdsilhXKwiDzlO+YEBl4jWRtY1ldt9hoA/XXV
gAYQ/CLrPA5deScNlofvumkTFH/Lb8zKNXeFjTxSr7eBdMltp0hgA5f0ZW49Pfxe
p+S98T1u4JCuNPu7eTzW+8X06M42v6l3pywyBVvPZ5KfnD7SvYJ19TfnTs2YJ56z
OljKD8DyqKojukcMl++sv6rrBVKQir1i1dFxxr1YYi35sEiQp93tVKCdVKWhjNQ3
okGksgeRbLxjZMnTcjm1ZBJzkWVL5P0TVpqka52VPuvnTFEIVGhTDY1pww9Pl/8k
UX5jG70lPTtcqOZay9BDrxZGvMK07IekOrWFNQ+vdWwyO0nPZifsLBfiB+K10cim
jVszvC6V0SMNFRp0/61BpRXkk6CKzd9iiwjt84N0mUW+b7JT+HlLiWRXCP0/BdRw
6icLhQ8DKuWxM/XE7bVQB3Gx8L6XymYBCwgofTpLf69QssCcMTULNY/hGExNIoo8
nk2TKMx1whfiV5o1/1xKwpZMtfUwFgofNdO1S++vZhsbCJwYB+vIKMCko2/lMYoM
+oUcLCvMFFDrtuesSjMuTRqEAlNIRAl8oAUOgrwxaLrvl59zncW5hoN1WxVXgNna
PWzBo0iAVDd1TyjIBGwlaFSBUFSvB1mh3ww4gGKdSLYe0fp9KwflrwC30sLZkKZz
g/DNcK792ildRwKigSQoPnKwZhVHSjnXET05FGA0fogc1fC0ZfKu49C1OBV0IEj1
sZQI26D4jYt6qO2N4h9yyibA1MkoX/AJVBy9vOEmIM3R3S65kI+4oxIeQFQhOD4V
64JT3OwloT9vg48g5EHJASBzo0hJgNZ5E6dQhh71l+tVgsq5JeJQrCG1IC8ZzuCo
ZGjKhAe8XlYE/57UJO7DcshZsowh8JmfRfqNeIbKIMxnJOI4BgHHG5h8BACA5nOs
R7CMIElT/pF1gSIp34Kos5VA0XrNCqFna9c2ehIwd69ZBxHn3YcmfLuOEN54IDZ2
etA3/s/dwaCFN53Q2OT4i13Z7PU66+X11l4aqwKv4hvRcJmcCFhDzf/6GEBLtoSn
+VYedSH9JbWlURf4zxTOLlqYaxisQFwnbauSJTG4hCylvdYquP0cFHvTcES5TzgB
fegdKNPidHMeAXA80yv/2s7gDH0SFrsQW4EYFG279CsOvRtoqrORnM2l/PBaUaWN
/pJbaDQ5xD1WXBx3weZf8Im9OHK0pa0zAuDr9/EF7Denv10PhPb6tPLFyG5A/nh/
UgXiipQrcL+KwxxSjNWXm1Ovy4+2OaM7mg7KAK3YsqPXzUtoBtnJpEBPGhb7ew3m
1J1y5ln18E6Iujxq66h2xKEPuTELmv7WafSjYbnc7TsMIP5VCMJgc+y+Gtb6zNxC
TuFyvGpBPe1/OValfnnrOFaG7LXcjp28TXLUOP4t9L9jPsnzqTyl4KdW4xI3tmkQ
+g6tYazTQ+PjqLHf9mW7RfdOvoCWnHZW4vjGWWwSe3OJSxdZDHb/Weof4MoTEjRf
ye4yxjGPBrbGEJRLudoG7fkltfIajjTLhKav+ptbckzFsG3F6jDaHv0CxV+H3L+N
MIUdlzRXNKXPeKAoCXgACLJGzxNF+oXFJhNbiPb7Xiq1RB5xnPfcYRxItUcjdYYk
HU6kX6uDRX/Uv1uc6jSylNXXsF+3+HWMq1FS/aN1vYfZQDyb61u/Mx00mLmVxJJE
AquuUAKuoA+tOXY1OkKUgs3Y055tkx63o5AnL3wgQV3qbfTxf4Wd+RczxjwF/u1q
q5MOMvdfh5RbbXH/VNwxzQqpAnXtuTdAMhAcXt1gxCJoDNyax4THAL0VDQimVkYi
DaIl5FBG10Sl78NQg2vZ7fA2jJ3LfFsgGZdoUFJ5a2P7m6SWoTuqc+pWdvoAUkdA
GnFp59dQgONOnFrlN1GplU92ddA+W+qlSHKBJiFPtg2gBiklWmPnITBruhQlypaJ
MeKoRZ2oU74EnWcQxXzQ/S9OWuFabNmvcBgzpQVbrHgFy6oenSM1StbcjCFxLkgX
+ON9WDoTrElD9MAiqQb1eC5XgMtL6qBn4KUaIyQb2R3lkfMqWZka8ny62QMH8qlJ
CSD8ZV3KgYFh1X1zb+witjDpjRk3WEqgBbmMmJ1LupAaFK53wU/pkUhyHPaUEiBs
EwomoFHiztSYN8/9cFhuf2qm9zhUaXa3avlj0NMIFqLJm4mTMPq9AlTqBcgwzcBu
eWPfLYOudor/4yCjbg3M1SQY7IRQONP0u8pIKoP7brWk5kVkT1RNfFjz6Hs17i6K
Q3DZc9X/LUQxYepEMMZ+ZFnoVym80at3V4QiA+eKmfBjn47qLs5Gw6CWrxdvM34D
N6e1KAoDz2K2Kx3k/F7KRoWYJM30AiPd2ji+YqVm9uPQRNzdynsB2bgwZE2S98vP
HGlxxJ7geFGSBGHGt6OSnyZepdcaWO2HTuuIJiVe3158f3kfM7zlIU0Y4nMyCFfj
//XpLbvrd1MyZ80DPpbZ4OcWXB6i98Cx9VSReLWnFCUZvkxJixl9dQUtSpxyRI6S
8PfukMdEM5F/peHoOYxD2p7BM9GcddDReki1IQJIku5Wx/ejf571+xxaBP808Mfz
WudSaW7W25e8NVQBybwfbBV4sz6JB85zfrXPJN04Jq2RlfGLRdGr357g58KkpCyL
rUk1vbN85YbwAD4r3tNCsijjZMcisOXnHEcIb1utVp4rkwYLxsYvz0t7vJurTyjt
Onh9WD3V2k41kSeXwo1nQO5yZIZ14QDab7WmLCB/r+5E5gxPOS1wc0WrriLYjulv
//0ML8bcRX/z6Hym+0NA/O6K/qy1VkNs7cSc2Qx6/+YQcmA1aS5/FXuaDEhdZZMl
IfEJSfspbPBspbS/pp/dBWNW+JLycDQU0KsCV8a81NwLDh2TjQ4wGhitMce9tUfH
bdt2HiZ9H7elu5luR+/Bc8XjlXMwHwhUw2QmGdXPHg0GSjrw5qtkyCQp0bHR9LIj
BT/jf3R2WPDxOPO4+XkTjfc4egbI3MOlo0RVW6LgXv2qB1N86OON+o5d23y/d45g
mq1JZS7OFTOKVNDRbDOT52tU2KkLeuov3B4+tCN00MzByBpVEVGEjxOE5N6BnHeB
5fcz2G0+shz7c68sHWG/WryDg4kSml+5/2FVfvULKcTEAgg11UvHRpi76TtxQPWn
8OQJhxy4tIdwVaSZkNuerKks9RwYYzD81CB4mcD0THq4s63KVZKYrHYf1cgMqBs4
awuOk8ktcDT0oYUY78My814b+3TFJYJUO7WMomKjoQG+ZxPXTw2PA6eA7ar+koGI
f0FjPhIKGrgEiVDahqwbjPIeu0IO4jo8yrTKzief5OWPON4aY+r4HRLhnD3bdPMV
kMOtdsdeUWScxdX/fmgIbvZ1u3Y5KjHZdYEqyoXtOw9hWFq7rkP9kMI+Y+frB+nf
7tAwBH4DGj2FgkYek3FDEObHSbDjZcFvK7YZ1gI7d48vs/kxvJ/gTQ7PD51N4FDe
aCJdoXtKAARaI7r/+PH7C2/dNa21l7f+tokw4O/mFPV0AL2Rk1mqNXACfN/SPUjf
Y1UMKLwxmXv8p0pLsoGFmTfnw2XemcI6Q/ZyBU6xzmqGLVVO1/4Xh91QZqIDGMHt
0DktqF83NfctqMEso4yXFKBsikNo/Mk8z8ocao5Mr17nK6Mpwj0ITzcQwTuxyXD/
LObqB0m6qTe9GoeCNH57YTWkmN78pv/hBrXYK2GzbEpJvqwtd5J/VKJ0N/qfPoIi
WP7ZtvreAG9epg5aXrIO3FF8O9bXT9zHaiyO3fOxYORcVkqi9r3wTXtpivZFWGf2
19RbaxiZzc7OU4PE8HYQTaTeaQnWmnpohWqurtgaGXFZliMqW4LEmL4oHCbrwEGL
Y64ljJqUuaR2a/D1UoG4FZRNcupj2h//FPDDLyuoHnhXPsJatCRYWNnxNITk10dG
HybeaFSBJWHTFKJ/pFeVtJXy10I2t+PNirV+9eYdPJ0m6zSZBhieJg0JTpdlHJ01
rx4y7Y+WmU8yrqzYEbghUF65wusKJGMl14kmiKhDOfwAcf7vQvwbK1gmZBG3pfZq
DNG9kfVpDIP0zrPbGtFsfNaXsUNpdAjPCSJJHbxA/AHU2RM0V+MWc/xM7hcJKnMB
T2/Ltv2Z9hdJ6IzRZNICO9M7KzkFqoKqVy2h7hUvMCzxheEo3D3xYk+AnWmYTWVJ
8zoQpFB50VhZ4haL419E1QHwRYX5NSi+5/C6EIYbEhtUMcsIZCg2Y5D3NCldfTh9
jqpDXjTTNRN9NiWCPBx1ZHYI22cUt702XVKwUp50cCtL3YbdZJR2cCKJSYpSgKSw
dNBrtM44SlHSCkf36yFQeuokRjk3NN3Z93isaoedBqi6VI5fPTXNIl4v3fSMAAuX
ODyxedC6//RjpEtcWDW/V1j5bQP6jzevld1+LhiO+xFd2FJBSUtlfHVg6P+DlMAU
1Ns2idnVo/mnDAVmKTti600Ot9lc+SLJ+ufEQQCCKWk+cEFUDmey8gNQkwOR5h4K
Zz6TGd18I9PEem80552UQS4p85FdU0sBcG8IWybYDklJaCcgp1GkbJUG5qy8D/RV
j6xhBsZmZnat5GM0mUAML4KB1c6QFA62c4fCeXUf3R+aDIdJusyjbJDUy1EmC8Ut
5BL7aqkF8CLR1HS8X7s0fEi9PIZHIbsAer9snoyRUmKAPudei4Lj7TA5Xr6r0rJ3
lG2AXzSmux/7hfagYNTwVmO3mz3Fg7lwQp8XPydCbDE8amfq2uWC7pb8fIq87Vm+
WYAhMPLeLUpot5BUmoFk1vWUP0/GehUFtHcYJGeXaGYzwc8wYb6UK2FT95+Mag23
xODs0PxdW62VHqC9s4GLiPGQ3rDsJWfOrjbV4u8cyGbTfU7wa6ldatnIQibIzYGi
I+Tn3Yb69f1Kll1TKirrGXds9wn+zFyw29Tcg3q/LXxx1Vpzlke3FCStYvQ2t2lu
GCkXqE3iFXju++tILw4dV1Mo0rD3InRsjWNmcHsTyfgpF+NCRRFTaYzFafhJ8fSy
W+J6uWr8he57cZRwhevtjKhsckwD8qeMlUOwHHmuLJOaV+LJSuWaEBlwP22tbIGw
DLfy4aqBkN2a+dMCq9bT7FKtmZA/d9I0zWQnVb/w1irRn86ThWIVTilpm9UKUEVV
jBU2CiMK2oS4EV1tkQv/p2CPQ9ohBAwGQktIPn2cfPKVEt1LhTaDGNvaHNR/TTxE
XrA4L1GuzQiPMIspAaWva7yvs8hAI0oiZQ0hRmmnB8g2l0nnfWyFlLf0BRKiv8UH
P8Wbt63GAsyubMkMwlIg1Nh4gbMfBkAAqBKHnPRNvaGhuWIbUcIZRTPv55WmktK9
mmxndmnrmCGP6zBe6XnfKYQzdJCS0kS39IpkCdDxuTx2YjKS6KW4+Utx3WRx5dFE
jbgXuLYOu5jd8wIgXHDgTJTgUaWSoTFb7fTuNanO/41KM3bk4BA6GZhl4uBzz+Uo
9t28J6Oy9o13SqQiRph+jJjum4ARhBeG8m9Qw/XxVkgBWTc6ZV0tetTkqHz7+cas
OrLqGNf6D+KleiXTLac5quiOBAcoVWLB31MyaiH4FOcFM9apMEbjlReEEgLVdvMe
Iif6I7HBdtq3KCeWXRhZApJGpvRqVy2vbof9K6aYM3PCX0T2QBMKWuBYGL80NQk6
SIiFISgWOm+eH6Y9yKBH2SzzKcfoNFwUeztQjOTeVGqO/9KNvYPR2h3C8f802TPb
yV3wAaRo7ESI3vQV2I+XwbCN2h1zuKCr4cUYVormZ4yg4/lQv23QyJ3kOPlyGYT/
vDeNtLJCtuDACEdO68RviUhI96MATSRDp/zIb0nb7gBtIn1y87eHFRrABS40JmOH
yjeI12WSBl9yBMaRFrmv9PiAUDr7HFHxvTU66czrlFEccfN2fIoHvpoXjnWFkVwd
J7jG6Ygu4HAggDRzrlxEorI5T57MopIVM68ZkRoVtOM/YVminNqWC8qd6eSRNHR9
4B9Mlvg3pA1E6QuKy1EHb5Z34/287uQeMcMoffRbmvb/0an0d7n26Mf8xAGJTYW5
8Yg5TjLb6f8NjXUelKVL9/JJ94WH3aqoB8imzYDp1xjtttIRRzjyVX90+0BfrZQo
wC7cT/DbEmY8d4jp1sZu7L9uQwjB9YfVgc9j3l286xXJdX4GUINY+mBcVP8hmlnV
Ud3wvBBijmRW6wxe7D6ErGvNNnF9HVWfLeDSo/RDm5I4AevN+wkeAhoPUd62C2gP
dFlZHSINV2U17vR3Kv3ZLPLHQciPVCN+H4ctT/CoZG1e1Slyv9J37RarIK/zrgPN
NkTyuqr2wbzmKaB0qvCRhk1doDYeAddT3hDbbfUT3F0+HQfYAjIX09CbGqzH70sf
IMbs6KUaKRsEqpEg+gj82PADq5iivIDg+QcxkSxu/eII3zXKq319Uuk/0Y/U71H8
xGhWwEIw3sUsIYv1s8yWjiUvSIy8bqX6rYRKk/urnlOLigfDM7b5sRucWOsCh4FT
2t82Aze9y17GE/Gtl6GeukcLMfw9m8H7ZBoe1GbzXLV4f6fqw1nfxTpJ6ZiNrOpO
Ho5F4/Hu0Qn+2OyS2d1d8YcByTqjx+9dLSuHY8ybQCVT5CPQUdx4R21hhN2ibzsb
6KhjRaxgMiO2S1Si8mIO6ikUvTNqw8Y0GZXhgiz2UdNqXZkbAFDiSQnDiAJnzNnc
TqYRmnKrZXRnLbCT8JpwhGkQlNdaOAbXpa/AtbuzgEfU6DerYhoyzUWde4OdIuLm
8V55ZAla6z6hWhm6Rg0LH1+J1R1zk1zBPCsMj6C/iwHkxFtih81ULP8mswL0OsRD
Ou0Qslwq2mLBDJq6f3DTpGfqevLFYgjFrBozlM4NEVxpCsKGB9NihSG9+FVnzzqf
GiiaVWLJGeoInf0eIxFiS15Zo7hQgqF+caUlPuE7bqQ0VOB82oCCf/fHrWKIVmE1
38SjJEH+GHeVGxIV1//T9hLZTkMEYlA2+ho49JGzHe0zITjx+4ImjBQkf2BxyF7Z
cV7/CnT7bflDv+ZQUUhBzhL1MyKs2a9CLtrsmHEs5QNzbcngVdHsVTu7HPKe2IY4
abcAy8eYmJXtyogjargZubEDc0Rzt2LGF0FK4GZP6yqdCJfu1mQDSOph2l5noveM
ECTHc0D5yA5R6+lri9kkGnidAH/+/2H7iTTSe2eabC5zmpZG2cnyV3+MwLxAxcl0
efNVtRJPnyyF+KouwfCiD35+9FLsblDB0Cwa812oywooHJcy6JmEBdztgi1yaueU
q5mvtlRlGjnd52gDYq+X8mKvjMEszheMottJor5P5rVSrA/cUNo1r257j+Bh5qO4
hpJ60a+il9IPKh0mS61mh6hlYmpQRhk6ijyfDRSve1B4JNhkqg7kw76AdQTB4bSD
yr15OhL3YiW8oGD3wobLrkWXCmOfGHMkCDmYjqbdJOJPIsy7rRRnGcv6rRJjgm0c
0CBAyA8/QseqSUohu/v29fP8ymebao9ep8KLztG1Q3QEpeFwB4eSDIy+rWOmLZJw
ICO98SJ7HNMTrPmRNS2v8aY4lbIGTS7w/eKHBLs/JT7qBDJ1oO4S80xTprmGONga
XZCxZ2oEHzBgoAO28E7aE5f0RdhpAZwl41naIztrQJhQ9J1WfWDVyu3UYdbBupNG
EIEZqYMhMcD7NcZYpsFImF8Wer5taEHAstts57PTKRNKp5niGQxPRF/z+1PU+yoD
80z81NhqVdLaOgz7onbzRWz5QjnY/4Pg7Lat9otbnopJ1/yFpYzrOoaFkdkZ6Rct
zEMAh922wMnNNgzgdVuRhXyEWhCPddk0BDttB/d2UfGhiclSZZ1W7n3g31U8svnU
EZunZlUpUX2kIv2uKCj9z/4G8d0+tJJP+2AKE9YmPQRSn8Ce6IqyytU5XOA3HSrt
uhwj1euqQO/evF3pWzvVEr8FlVJ7w1PmuT+UoCqxMFOR1YGngfmnBGPlt+H8fuXz
VAaCai+kfjncwa7nHglQThuikWg00bkNb6QMqIdnrAwgX4Qj0Gk7hXhAeI3ctA7L
0ggIN7l3Me3nv/Iff0rrst/iZZ9wsyYuCdw+r2ODI6R/qQzZAHz2MwjQycnUmNBt
iU7B6NEPags98x1g/MppQYi6W5op2pf1Fe2cQcqZoncDsLcqFoUV3ZaDBAW7Au5O
N6ABzETR1jE55uGfUSrzJIweu4W4x+wLv8IWXrows/uh1+O7nzQ6mN7j1No97XIA
jtnhZKuq4z2qYqVkzrxdT9eRnyUBg/jKmWkpdMdqIi6efMuQE9sMfQ8tw3JGFETR
+LRuU+Q2/+/cIVlNjFZf+2RFAiD7dhU+Xdm5dn9+WRvEYB6s+Gp1nlCQ5M8d/HHL
NhxrfaQndQsdvSpYiNxHXdzQl7QZYuSmFoWGHMcU617T99q1JUyjvECwCJCbfZQA
gvqM94QjECPRy9lXoC62vDBG6ub4wsb8q7lOwJj78E61y7GyuyoFwYrnvi6DGhkF
mQiP/9YOrnCrYWsVDQ0PXSvGU/vXGUD6W6U7OznwTgy5LdLsS3/RwppaqZeS2FXe
Rbvgbf+yq+wmWua2bWcDM2WOKKhbxNLNZaY1IvoSa5Fx8pPnmHm/kpVKpAykfqDf
oRjYzuKm6z82EnMIxQIRSSjNcfW8pdkaeKa9MF3yPwuy5JEfUhhWFlWSqMlOsmm5
RAK2cK/RScKeqlGuK4fT1x2T2LjYQfBdp82WXQsyGSBu6U8qLKF5bp5VYlSC8cEd
ipioZXMurpTjYJ2Pn5dmGrvH/NAQuIcaxhEvMoWnh++/SApbhzP/kGW98PMvy9wI
C9peD0/0Lmu5avWmawrVS22BThL2hyJdPSvDDkOG6dXZhOf2Ds47fpwnXE5puop1
sB5IgxijPN/9AS64rFauNdNuCywdpAV4GEVcGNC4vtHiXKT2H2JFK09vTeArdREZ
nrG01RI1fiEaMRY4ezkKuwxC+bRrQKzEv9LudWGFuyyA26g0iI5u5srxTXFlJvb9
o27bJ+tH6jA8H1egMB1uCfAOg05OGKNz9U0R3+wU5jQp2QbId9tyBISHALrtuBil
1mgXKRue5qU7Yuf1QCckJwQAJ79V01QVG+fpKsqeceVzCUAm9xDeL6zgJgIAd54C
WkrytKrmuixNczwq6d8c7N168IwI2aMREdwJvTNNhE1MIvfZG09nU5sSVHn82r/x
89g7CGShcgS11m6P1arnKJbYy9CnOxUGQGH683IQKTCVhyoLXAktSe09j7vWf/xV
im0w5/pJNy6rQZLw3b83+ptcmB1v/vdRqdelSPnc67zKUYfM6zEyboIFDvZacGS6
aeVOGSdZ2dWGHyQfe89EogxnKhHTLwd7JOOwch+U1BgZom4977DVEpqq/azYs8IK
tB8YzjRJz02fReyAkc4hyT+ewGMgeRxnxuPQbLlgkfoKQK9VhuPyubZpxPnsl2lU
Ind4bOuml9QcKD2f/dzjKvEx9GWiHp/MbQ1+My5CA+fKHYLOXYl8zVfVKzazvEcZ
RKkgKA+HJU/XZbAdD+im28UaREA3ZW9AWjUcRSowET4pQxQsSJ0RBmh4aixCAc13
BWT+IK2TY2mdQW9tYdPvvyHJ+RMfx6cJSdmNh2NtJHfPLSPOgjxfgUvEKuv5fY/9
BisC7nI4h/SBMixbxS0kO/9zUOSAux+uFWQMorjC+sac2oKAV3QeGB4KnGO0Klhu
m9YiKf6/Bvb1BEo248pp2NhuZVr+nzu1zhU5FKMSfzVVa8Rv/7ovJj1ziYsNFqPc
Ez9GSnyTjbIhh4gVEyWobA9XtL30qlE3h2yFPrIFmclMsZMrmYGl3EWe8TIjhW3/
Flbm8yMwmdRzKKJbh4BjZSvS87fV8hB8TvR5xlxXQTIPqUC2iB7HNCFunNl6r05/
mvwSp0HKRleeiWjzKrnwSnpi3pxIGcvqrxIg4fyh8GxlBnMM4EM9p7/2hEt0tgAv
CBdhQJpJQjzALjxtpH4bq70Qc2dA74rq9frX3I5x3p3ip5CG/8LkqRSFR0bwd4HQ
cW+d0hI3e+zueA2Y1fMYBOc1IV99NIKWDsyYnl3h12BSU2KL40KvM8oV0PVksbmX
9nmVvcx69z7He+y3FFpHRSBNJw1usgqyVVCg3MJCR0LOjCh6CwPEEV9sirfn6Ejg
mBGwztLy8vppiT8sVQ/kUTp0fi4UHJ7XAvDeWacCLzkLpieA1gtmHjGpopm8pZav
8qLaJ2KPkDNZzjfk0bmMZTyHhQJ24yqrdO9uU321oEhR0+OEerqpVE8SLxGfKH+B
5Mqq833W8dWlCZoVcq4lZXBcf3EvHmbW+AX4pFzHoP/qfLrzaVvWJHc8L8EqJu7Z
YVb/ha3K3iQdJIP1VQ0fFz6p7ZFxSonqdA0NKWg+ySnqQdNjI1YshcqOo9izrNAI
hw7yq0y+I0flB/ut9EIKCF5HkIFaQk0w8QyodshENeYBzJEJ8b9gIzOiTDDKKETK
eQo9vOmfg1ty0xyoGKIQ9PlLoWYhtogxQtH3jO5bcKpwMiPXJokmzzhuTRZpibSw
UY+tpHuoohxrh0KDOffmipTRmpZUQhMcsSDHBhu80rPRFRpCJrj63iofMDWDLViV
8P0HaOrR7UwWXyj6k8tzra53V5pXVhDFnAPLBoG+O2tiDX8BZxbqLxG7T70J5/jz
P9QhSXdP0XYG49asrzq97Gis9yFbKRgvJSaB9pG8PGLJMYsfbzP5trk0st/khbvk
M21mbiT77Jqr2kMIaP8HRenB3GbikqC2ejuMfT0rxh5g0QzOmKFdETw52cXFhSIW
U4ytAEWxIabMffrh6qh1lD8w6t2VwOriLNHfzKVfIpdh682/D87y808wkUFc8tZZ
scG/YfrQc/Ghc9z2oea0MrePg1RqzZAIne/hje1EftLweJCZk8hodyhsknGgI4LK
9ewv2OSXr095iRHeCj2N2p0SqHBfxrpBfkKAM2htYYe5TxyZfodGZbYc1YuwfVbl
ll5PFkW8w/lE8cwPMuzReBRjpF9tuylv07z0kSJ5+TI1/kOJNDsc8f2ojUifqhN+
lJeUQq7YaPdmJsl8n233mWk/XDx8BVEf8iWvDAzFUCmqQPsII/5Akmlp62iLkNCP
qh4yrlKzll9gW3xXF72k5gIEgtNWpsF/bHLcCQNVWKCMcUvtHMrq0c5zVA9Uq02R
vMFWn/GiHw+Xh0TiU9jz8oGsvzqUZkjIq+V3AjivsYKRGu6kd/WfCDDFkxQmN7eD
3lkgBDu1QfyXADdNmw+MILyElSYdhKFLjwSTQNX893ZuD7OyzM0hZeDZmJFvnI+V
tLySrdZ3qtOvWDo4JJox3pPiWoHakVsMlfkOnlBobmcpo6tFxERG5V2e6vwuFvV8
Y3MT9EUyLg4yCY1kF+grly5LkDpmWHh5W/9d1SEx1KswEFVkDPX97c6F8Y4Q1m5F
D3AXAvnUkSzx1PTXYG1FcSs8Irv9YvyuNZ5zXMxTdcsC7lV+X261etI+SEGM5x7f
8QouH5BsjoJL2h6LmRzsexmNddIWPkb91afND5jfpr5dLpzgGJx4+46pwm2VSsd5
AOAZ5qn+spuTNsHMBqxCbSMQblOYYtxtW066KHL3Twi5vtZgZtWTD1B/ofd+CNKz
jugABqF+4DnLBNggxqR23BVwPRygJCLG0awuYpdBAjEg3a6HpaAxyle4rEOAPegZ
wClJEtzGsZrXoIDlHhgMX4+VUF52PXvxaDdGu15EcmeWa1MHYSPOunMa1PVadde7
z8E0z8L9jWeBrl7GqPyfxBDHoRbhlFz+o5lUyZeV+i+MveMYJDjALvp71bkA3cTK
FQuhmTpVijZfXNAlpHIGATxd3r1RDXZHhqpDIdziHu+tjKm2ezfxpj1WIj9UtVBy
6x3+wkvJWI8pbuHssRCfaRhcOPp6KAnXo8rfTI4iktcS56o0Prf1xYthj2efA//b
vwrsDqEPcH8v83Xe5KIoInJTsg87gG53pTFBA3a1KzoY7c+R5zhJWYjqAC6T+Qsp
uXKJ0ElxOTtw3IdYObkrnIQvstfi7T3/FBSPS28crixrTWPChasY+RXKCVXuPZUU
mxt9p2f68SmU5R5XOU0YWG2mPQhqEXgwJxhUFS+2Id/cNNlHTDQpWI3PbW9GnhbH
OJIbEXizNOPOhaLslGJP7uBRAaKxnyFWLj5uIhXp+N2+ryQgZECEq/TqS11ua8tl
cyrnVgHhgf86prpeJ7GXSPGsLhgb/ucMARRBhUJRolrZoiHKjNxAd3U4ep9D8yYq
X0ZR/SdwDWDm/wBh7Dnoml2jHB+1V3frA56Uo8Z5jo378xVnOww1ZD94vIhu2+9M
3a4VeKy7lSmiZFx69vuXVM9ppWLKPbtDKqZcUZUOsaleHGSbg9+hG9VBuwqkGO20
vVqfS4NSYUv6/d0kxf3E2t+oSiZtBTcBTum0fKC6H6R74c1ViPmaFlsvJD2jraHt
p+9z4I6XgHfi07mlivd9El1CjtKSR6GBsJxQmzDVu3JvKE4/vbuF39861fJGAghv
7iGrH8o5YHTLRjT+JfZ4xfsKlHOwN8ZfOHHZqtxraP1jltrkCvAIXfnMBkflKX9q
u7vNkTeIjERArilUk9258LZh8d5zj7VlBhSfkRbWyrQ7vsAzsdziBKYX/NSqeS/k
Y16hxKw73avLO8TKYVJo/ILGdRrABGj+Xy3mQJ/GKWDZwLyBRHeb2HQDMbgLWENW
DMhiUQvg+nmakSCNIJ4MbEOJnDt3Z6sO/dVYwziOdOQcpW5qrFsqvBYSsyMZcXuj
Z3MqpXz8nc/pv5AA5S7XuyCZaRPCX8Iq/bGd3tABuu9KzA1OveHhsDmxqIeaPN1l
SObsjvM46lEv1+Dpun7Kuf/Xocvp7vulnXa+Q0agc9p/WBE8GV8AYPRg7iidIAN6
JnqO/ZwJLQUrtdcwJUiNUwHx1ERhEHjWpYGaqytFMVjksbrroVozMlXWtiK5OO13
RiOLEJzhq+5zdyEMMHT13kp8ckhuyjg9yQ/EJGZOX3Nzt1qf6IwAIDERWGw+N2RO
MTAZmFcBKxNRCoqxm4d07/8nEbKHhhzwA0JMxKQeFFdjJo31qlAJ3upruP2EKQZe
3+3/Q6AAJ16EkvJF7xK2RNUKxik8esQgSTs4/o3aMul1eNevhdd4F93JEc733QdM
S6l+H8YrggJ5yspZxyoyo5TuVDRITcPGWtkkhaduyEAnW1vy/86Mk3QmWZmibfNM
CBIgJNLLMA5rt/ZJY2MeYvuxNogITgAF/+iNiTRHdbwOADVfpCYG+QH6ue6Vrafe
Ds87QYmjKHb6BW2lLHgYKj3Gkfq667WHN3xo3is1P0/vf/SyH+deSD8KHSou6Hql
zdwc5gmqwhPAfzIHvADdLlo0aOsuSAIyPC3vWnv1vZcdET7L3UD/Xtk8wV6NDWiF
TTNCj6O0h3FZtPALzY+vCQr/Pc4Int2JtzgZiGHXdIbz2DG+EuG9MxVJoNl/X+ra
Ova6dcQhA80Zupl5SZ8pabSIk7djlqup93NOfmkob5nY/CpbFqAGBjJhcrkAulDN
Of7TTRFakkC1XNrKMmsgbsr6ZiJC0jT3hbOogDIVVv8oAhjkFYIirkKR/YrCBuA+
dXlf7pyCUAPA70b18LadVTqQJyCO1f6cdTcg4CGqdjoyDkfBPqYQ3UEqOit3MayM
ckfjJwHj74NKoS8m2dJLNJ597VIQIIZe/YFQA2734a8POvh7bdru+1gO8zUGT4AP
lvhKQCjitrgjKhFe9PG3eFVHEPK7+TOuKA3q79w6fye23IrRk/TSnDYIi9HJbafM
mhLiNLDpkIR24fFa4hfrf/CSTSt89UhSuqXMSTFulnRwBOhY0rjlpQcPnPGM+dXq
GBdSN9ubBH4UiQCrfgRXsh2kAR244asVYT40diDyF0E/oY1s+Yk+YY5bhURopFW1
FvROZgcubF2cgPYY1Ib7ue/0rnkcXepHy6YYDoU1GQiHpYdVHzHMM/TDr09CvjYP
155X5Xcd+iLygBeZSsh1tgbIreC5JZjbW0N9RrSl9yunggk3zKJ5inpxFMJkDk6A
xfHCGFgQFsx4G23aGsh15M4okMc0qt0QWSqfcet9nuPoQwpmKPtintF8EFe4KlZg
tYw/0r8U3CGsgtr59fdHS7E5k8aXxDWHCFVRlYVeNsTx+tSRkDzPtZeqeyO0YiXi
JS+Mic2gRRQgilwwHSELcPH5neuIKZ3/fHQTzjq2f+IjgeuMPxb5cHPSFvEnFzQP
n7Eo821+yzpfQPZuNpUArzSiM/DPup5rT23ry+4tpf0hPc62HNQbBL/nLFQfnnwR
hmbu36K7JbK7Vu2Qc9orK68kyPxMSQSyF8jFzopuL8ARC+dDRzJmIVRXm2cctN5R
+7HyWnVJXmU0AcLRKkVw1bz7Jvxk65PW5yjFBbe1vyQbdk2mW7MbZa+YKKnOy8dH
EHtDCzbXFu40Us3pW3Dw/k4nOMA/n8yRPxuXzRSlBcRMoWiru63cwza3eGtWD+I3
YXhKYiUCSA1ekBft/0HiFTz2ZnWRku4KSb1b//ruHtlDLrDKyyMzbZ0Z9lUD1cv5
M3XOfQwSz2tT//dwg5ZeM6Kjun7TZNB2YPy22EBEgH3My0dP0wkyOlKgyYycwVeT
J8k1Poud8rRoCI9GDtn0E4QZp8zFmPlhoOoRIhv4ayWxwVzSUm6/JqF0E/4AhzeW
89gUHGZu6d2csFmVJAsa2VALU/qpDUrjDNdS/ZhqIYcKkfORslS4p3H3uL8XVCka
A80hvuW7inQbhGyVIbigsYic6DRH4lRNZWxhSv/CCRJA22wqMU64TXOah2LohrMd
v82/vb5A++lyMuGGUkzoiTvkTvQm2s7L/cNyRVAYfZrtAjqSUXeDaHqYQyMMS7GT
yQoqSjxM8SGY1N/5M/gaMerwxMHl7YM6IbTgvetU/TFd71h0TM4L5J3EYb/xp1cY
TcFR1ihi5Q6MZegLjSkJeAXdOY2L4qpoFgIzvP8cMZg1hQxTIEO65ni7IQ0qRW85
He6Mh+qtp5yP0e0Dpltb+xBO77tx/DeL/AfK94XmCWu0vm9a/0PWZJ46Yadgedlf
YrhqQIBh606LHtbDGnzASiIVK1eiLQ4S++ZVVxLMTqwgX0/xjqCCiAQiem0rErND
ThI8TVkMW8Vx1ZNbhimxCJEcMRHnzRf0yIONJ5SWBidvnH0mHNlPDIgiyYeOgQGg
nPYtxacJlsl9m0PywbFt9upcTwfQ+qx4NhpoHCSkLjIF6WZYm2q23+sKKrOZD+10
KQns9jw9puTCSMLCks0ZEWEUb327bhtKyJm5oPdMM7Qq2fxcgO4qpEJ03nrjiZgN
w6I4vy5w6RILeW/7VLfpfqVpnWV01CIcXR1rjOOlDwG55dZELbTofoTJUNst7Vyx
0DrNC4D1yaHvHEOdV2QMdCQ5JRSDb5LP/VVqqT3J/fWNWvZig81MHI6+f2B6G30n
VxpWl1NcVjstbCdbzgaMnNIb88hrnUiVf5C2XeXwhbZpqsLtO+bpXQwlLXxQXqsL
Y33eKIF7kBW2VsSvvdOodhFCvteAWEAESxxc8dbz1YhykfHggix9pf8/TEs8HDvT
Xr1tr7MIiKteb4f/rEhqacyeu+eIRJNpiYUrybrSt5zPWspC1G40uBZgVKmXZnoY
Lf/belZlLTZxVub6+jifAWSQNq/096AYMvGSXPx4j94uu7BDJgc9BFo+Pujly0Bk
ohLIBl9RhCJez09i1MfoVQ6KCHB7OUk6WnnAgWC4FrOOHD9y5zO5wgD+Qjuf2Wzp
XFPO16Br+1vNWKtYEdvXtRfM9z4wEt/pmhS8LH+fMkHplIDIGrB4fhiwa2KVVX6z
iqSMRgPc6h2fT1Ym0UY9OqRvxj92//5qvUIG84dn2rr4EJ2dwPFLAjBjZCxsSxQP
3ueLcnGSnlQjfIOsN+eGHDKpET78fQnBinEjXvuXXCcmWNtsgJXrzMUXI770X2eK
NWw5S3ERd0OC/6U/spv0CLQ3qz6hrh/8zPlyc7RhgyCcz8IA+Ghg5Vi2McuSBAd4
oKNwY8drCwdx+zqRTV/0EearqXlxPtRjvFgUcyWnVinogiYJlpTcZtw/Wgl21Zgw
Jx9YJU5sRW1TYRKY7gJ6VcW9aRVur0CPXNRLXtiRFlQ0zjVp4butsi4EQFKzj/6X
R8jUZqQQWfv0yGbjlyUH1E8RxAfJt/NMF4Rm5mSRDhKPsm7A0qzM1wluU9e4f6UB
y7jKr7UGG7SoCzLSg9Ocv4o/BRbAmkCkafkBZ1SSUCqwsruWAG1mELve9PfNtupz
h7zSMqUb9vVQYGfsg35jAqzsJeiF+IlRUTglzfbGPPqJskXV0YNie7DKaf4xILL3
WnsMVr9xElfh+5DROozVkz3BokNIWN5Jui1rANXJIJeefwJCLBNONU8tsxTxQoOR
fJnWLBS+ggZ50IPwruyJlJc6al28CaMu4jSlTmxbmG307JGQn/vrelrdLiqCTVEW
S9tI0+yB9xy6HtcO6ajLLFs0hv/8e2vcXrQ9TBm+Doqd3OIr9tizDIovnhke7OPa
Z2mKrtwdG310AwveWOF8Dg8SHPWYczyT/9+iK8Hha/ZruvJi9j85ZTaCNfSE/Stc
NLHQm8uXBzGTVq8swsDdN9ux47+KDT4CL9/UBCpeeheCueLjpqt2KMsok1LLl9hI
zW0Jpkp5IuwYFdxsYSu+o2nvTscpyZCLyHYW6nAMfuNrQnG6A0b0oSSy0xchHL5q
gNSu9SULfGD7bRhQ/l+mVG/2hfk86zILRoLE7Z6xHbY/HWKjmBO7kC0sUvAk4lmC
AgzqvmeKYNgMlpkIwVehtGuSI2kd5qjwEAiRiq92l9PsfJ5EeeJ1Nc1SOq70Za+s
9f5L3CE8H5IZYH51FM7S1Dgw13RR/gKbGajMi8KO7K1TCyZJgAKsNXat70IUFs9u
UVOD8IgQLUGxPFLnLZbtlprdpEvghdz/sY6fk212YSf7lj78kapYdZTfT7EzVzSt
kSKekJ7beZoUaz796jlUgYOmBcHRegQK1haur27r/eM08skr3nDkxZe29QBay4SR
PJGxVF2IOG6rOV8CQFjDvF+Hz/FTsg46m/vleCCs3f+5Xs8hjzjx6h/MwbdikJYQ
kIGmRwnTb8IKkv0TAXmMBPgqM/v2Rct1FZJHd4BARNq0rYHo4NIAJNESM9kxH7oe
Pv0FcOouv5tWDx178hSEmNATVzP8uFcfSETGoDVSxzhm4/H7zSNJQqiT3DoGL9KA
g6Wdel0gYQ9V5vtdTUGSsxbJiHw5OUE4scwxV+crRJ5Q8s2iPKYGkVWm/k0iaNUK
fRu7YyPX697h2IxMOqsg4SHIsiFCCFgfPZim3NeliXYWBPaY5pcR/FJaI1qdGpOM
mBBh7KFvDaOE5tVuhkiC0m3LhfACkwMBYHOqGboCQwAFx9PWdeW4eU/9g4s/qOig
ngCV7yYF5uKNlB0e3EdvHT1PD+l7vAr9iZetE2DodyICg96FXPquFth9k7B1uDLI
hZFKjEo2AhrRFMQVHIxfoTaKXPDqA/lydAjEuD2RRFw9b/+PM+lNFtOQDap6Qjh/
k1fX4mHglTih2jUq+AN9fOd11NLvPGREOIUgX1UV0mNnYLXiT5y+5VvlJcSPnrI/
5FxioGGqyYZcW12uLbJDfTJgyRxeatkOzi8+RzjivrKT9trKbifMf5Rcr9XZXbEX
SGYhogNFRiA7NZNAZxaU3Cpnk0L9rvOMOtDLZu7gNpoisOlhLBpY8m71SP5hZ42R
l3BPNHe5glfxhp4hLuAt92u61+X3Nf0qTGjiK87BJz9nt4IdTGcrfcNZlt5BSUab
IXWpV4kboB5QyfX/0L8xv5R8OEFVDOtT8jwITE+HWYDY/or6PZRWhGsdEoSqmsti
QwYtNPjJCqWomjSfiHQbCnUkjWgSzFQGJigx6V7A23PLxVgUp/al4hlZNNrsUx8K
eW0BCFZwb16y9SVnZU5DgmODcde8yOUJfb8M8YxNKW7LV8fgjA+xR0JwY30dUd3D
NUbo+6ik3u+J+rnAS3/vazIHR8KDd3jMRmWKPelSk/g9ofP46yfqa8c7oI65qppf
Oo631GX7JUCn84fK6tFneFrACEZeVxRt5NPQ3WSuH77nT9oU5Xh55/W3/Chk1YeF
JpZfjn3JYpqCBgclGw8uvcEJF9jcHJnF7waidtK9GELkseS9cx9QT0Rj82BmuZR0
rqSU6Qy6LayVX+JcYkGSKb9AqUHkyrBPbmyGJjCWJUSLgcacSxGpy0RcFpqNElLH
oVY/CazXzQmv4fcQJzvz+q92Bje4RpVggO1MC4DUDu5v+3JPnAnrptVpbQX4pDmE
lVRl5wwMIu2qsbKT8SWQSZtT5H5rhARcdFxud2NRRPxLstKidQD5lBK9+qSt8kJc
hXVZZiaerSpVPgexQgkZu/orFmFs9/O9hYhroa6qeB3C1vKzRXZLRAaRKPAGfvO/
oKB0SZKVppMz6FxCSaEIk4n+nmjylObNRxUkZqT+RThcyFITGRpJbKzD/r3L63aj
HlhXOCsonCcW9n3oMw/sUpmjwnAu6v0ukSbjRQwq6tF46SYXnMtgu4Gaih5AwSo3
iRnwRBY10dZYl4B7CdmP0jucmzWJXp5lRtNkG/lEvp7YZI7OxWn1gSCmbL9GYsC/
vjdSEUHIhB1QZoXzZRBKngh6OiHGfQIh9XGysjWwbwgQdcmxlnt9cnbQvjsMNXKJ
j9azFw6q1f9e3+APY0jy7ngcJBIrbrShxzWB9NSb4OG8lP98Y3NBeaig5OKGirDl
ZzlF0GttENKdNlTDlwud+/F2jXa71vuVa/6kZ/9rzonACDaw+cfWqLRZxsMf28V8
MfhbWS/F/5qj9N3wzZxsOls9DegAnGuRVbS57rmxtm3d3Oq1tm+Cptr63Rscelxg
Q1qg+Wy5Y4GwavtT4rSl+BDcHe+avSJa3UJCtCD+rJgS64+aErKxJvgSg+EFFFvD
Fzmfbr4ZFcVTu9Yxv6k75xfqTUZZnRN/OtkowQXzRfekP/r5u3Ym9w1nGhZVpxGW
NBiUjg6gjkm+yelXpm3Ood4Hwh10Wb9EMfVjX9C35KUGf8+WOmMG+bFsTxB58Y3K
iEKPqrCUofeGz/kHedIfrwvjByaL9sSeDVwgZsOPS7PBV4kmuC4p6TD4zeV6qTY+
1JVfRh/dhL23H9/3emBeFiq4Py/NXhSkgOmiik3ivMhRprY1Eg6rwPJj//AfN+bw
nU6LdCxs8+eUow/Db00nbMPfRE1jeE1bf16A3ggpOT+wR6qYjIOJp3Uuqi7xabSD
Pkv6WDymABTHDp5zRs1792TO/rYkpw2F/S7iaeZ4UVGCoLzBQjSN9E1c/UEaNReU
X29JxV4pWWCD4K8mcTBzNLAg6X+vgH4aNF3jVWWKWZW3NGM1WvJzmpp/2DkKrpRz
7+iQbMQ5ZXcdJHTkNPKHgtcC87yA8a2tSRt18Ct31TNNIx+3pLeTUaFPuxcp+mEo
tB2/00/10BSo6ESOceSF0P7t6mtHr/h4fS67IOuedDMODNwGG3fgiWRSXkQsVfUH
HGRWtvJ0GidyBN+gHvslEA9qgHWzwGjpi/EcqsT6xe5TraEeojGjhqSxL0pSKWPr
Bs4Scow+fuQSDsna5fXaSLHbVGKB1DGKZhTJ7H2xJar+YBsiPOpnSMalb3eXx5tA
C/NKbF8eT24OxtfQhW4IvGjG5XmHq2Pd5gI81MfJxmbAMdG9M0NLUluOs6YFibbI
v2gaEU8EZ8E6zSCLZH/KYSUvWaqU9HK26Zl9yFVH7PvijBSbZcag/UKbfU1amHtk
mSiNEFlTgvCVHWBrmXJ0VRKJOi6VMdpTc19OHaG21qjQKnNU0eJhFW7N7Md/gXOV
OZeLo5h1gruONfWg5XYYmjJPseddXV5ugE2y2q/nyItttDGMsztb0r7U8eqHwHPB
1cpPmJjSanQJpWavw3i2xC8p7uXcT147xU5yLNhAZt3SLx0PnRJXB9UwPVTXksrl
tGPIRcXygjCos+uDsfdVQXpKV7nMeMyU4DPxOTxZjUiGEi8oWD6hXi6PahUwytP4
8lseDoT9wRuM90YYrVBiRFnIfmsVQK+cPaAzbI1/jRP8v2mNqu5pK6BgznVlA38p
eUXzOy10MX9JJUb6vWJOiWKfhadnqfTFhd5fcMpTvOdqxvshIhb9+uiaSJpV5yAH
tRS2yDUG1rZb4bk+D2I0jiUxEPbQHMreusk0T5ljxnENF4M9+epy8zP9hLeiNHQ3
D6n51UHJT9L4KkiOh0EbFgHXBsjyQs7gx70Wt1y0P730YLuDLGVTqUkfadVtltHV
tcxjhthm1Z8HDYZdDh1W3oqZvH74Lbq17R813K21VJ976e5Iid6dFIQN3h9Uo6Rr
oOyXcvKUOmlvOT8yWj/ERuIGWU3WxubqzrqFhsFuCseWIm2JrHkwZm5f2GnQNope
90pTZQWKkNV23fViqwZ92LibZlb0tw4ZuuthQKquR4YAnCTnf80/9Xbzv1RWKqFa
NSJUZ/xlc6tSCAIHPWEPTS5zE7a9DVAlbN9sbnqEhCAMpy/zT5+8svtW5aVXb4Dn
Gf7gsPBqOaNc6fP0bqr/GftttHgwgBmKWTDhhUPpj5meiFqGB9CyDI7Z7YH6BiH2
x6UZCBWuc3hf/th2xs3oAjDBiqrRyi0uRVNUnrVbvdlQU1iNLSHCfd2G/qE0y1/Q
C73liewI2MYzmmCHZqpQVFptyhITjTolaQ/ksavEe7ffxe/ZxsbeJfuSpKgp1JvL
0MspAqSb9RSrJ11st+eG777jxhEGgYpgiIbNvgC/Vhg3wDFCu2Z32nuib13PnaXk
nW4DRudEr2Jrzlt940S0+/KAZGZobcmjgLq9D3svgif+R7NORs8A5ehH1KiNwWHa
TkovyA6mPCicXtugQhKQ3tL0g8U1zoczHWyOqiqCTdrWubH7ncT9tD/+zsGMa++K
iU0ZdTh6ueac5fpUTxqYjOoEZh7eCMu8cZsCWVkyRyjA3PXQU1451pnOiD4mik6Q
ekTKqdps3Z0w7XF5KG/RpfxXSAVWcAEQSeuOel79AiSr6j8tF+h5jgjF+lB33n04
bR4GYQ9XYhcOQXImvlbHxq/B4DMX6vsKbytaXpuOb3EOdhvkAUSpfuHLnqAeDDu3
GkFyEX6+/VfhSjJRB9dZwQXq+6go6MsION8MZT6cujL8oXe52FRlEk1WOQsyF4wJ
PSV3GCcz7kKewppHoR0NVPiwr8digZA2bDn8G/futU+2ECfoITM9hqcfjQROA/Wx
N2y+WtRNun3EFg5RLO3erdglxzEuN0yKSnX8ZmJa7uEl+y/PMZW5XKlFvAtR6fKF
2nvu4Qkedz99uawba/v3NWbu7nZya3a2HGY4RqvECXeOEUyoDi99dWb2T/E6fdDU
/gKbFkfebozX4LaoKoE5+2+eAiu0W0ggockEu04ZZlu+IALxBPCUHQVcXyVWes27
Z99D7uESiEhco19KPwkqljndE6O8Pmd8MVBhMkIzO6nc8fVsOPvrO30HomKaVud1
ZRR9dfuwJx7IrvN4hX3oFOo0X5i+YkWGTLuAx3o7wHBzNwTlI5e1Y8fzcNk3gFO0
grHofgHpA1SNV3QQL7zqbcAwpdU9yuYzJ6cyDYY1xHxs4MK5SvTmaByCIjYSlIGd
LWv42UwyyOXP5LpBwx8ej5s5AFnawm8oJ2dAngxkvMfRHF9P4z1/umPOuCN5UTBS
i5Ynh5FY93BjQZlBj0t7Bz+Za9aaS0TfNxFYnHw/3vUIrT9A58UFId6KDKPLsD0j
Z6TYg3F5aMaujHP8OTBUeAlEKQVG/KVDsN1bxbg3PcgEVA4/BNEbfpf+u/a0+mdj
JUH8UtQUMyJkj5/cBnwais98P1gehmFArU2pduvFRaEyc5wJWs15CgtInsxs4zO2
hd+dgTOvcMu+f9kMCeXJ7x9PWQd1BpU3w381YBceayx4VI6ShVGlT4iRWdEZIeCw
TdfTPNyn96ldjZo7g053dTGUYjTMsg0LLrA6j4kiYeHxE842Zx3oKYTK7X+T+Dap
1cHmeHQvVP4pGePM6VChgKQRTpMKJr4mqusoJU06Gpxt/+NX0MEwqz6d/Hg2Ehp3
tFXX3rmDpJCSv2S3ejq8ZxDvyel8TYWuMY/iepC1fBbVwj1fxvmQ9oauC1h5Z4oS
xQwDJlZxGH849AFDhANfk3SOjo/MzVeVDCta7CfZE/3ntk1FIifnpx7T8wPxUE+N
z9Ja+NnDgxRv3zoYjP9i29lSbnKMu3MrAVkFFwL3lno+SOLTiL7pclLN/L6ucZyh
RnlTUnnRwVZhOdzbq2+qWHJCzj/veQCwPPEzCDcMWow5mJahoxzkg9qZPpecfYeA
P0oMJFe5uDEPWA7jnceARHf2cr9lm7L9nlr+/sZOLs6ZpE3ZWgRX8iyjHf8BNZgn
eTls0firWPGTW/kAYTV09WMnmeQ0mhuBqty05A9vhP2+f217pm1pdM5YuLqmU5SE
2X72GHdXJesOy3s9VAxfpuMoU46xHy3JkyWtZpLLkqFA+MDKLLCIERAm+L4tn5wt
W2TBwrqnYHInbULUPVofQP0UaxBX+5QqbM89Jz9v9PzVNqUu7PWI9s0kR3lF33Ly
QiO2AfqN67Fv9TUyJaT/tlOhYGDDOWMoUTv1kVOVj0xqWY12Jzrs+Ysym4KUT3Yb
hEAsojOXD0EtJkA5gpEWaNfKZBsMnfw9o2kb4Em9mUYEBiVs/Qn2GOnJNHo2iVzp
x8mZDdn4LI2096cjAXo1V7AcFKKzvI/PspXCE0MJQMs3p4xRBcoYGgciqwhRdQtR
vZdQYHtAKhfklSOWdTCT0Af/YwJpe33rTAiH4lSDG0rUK83cdLWby/ndO7sh+LSn
bLP8/sM6M5wobAmNQwvvnVC/CiyLyzxfhsha5X2Eg/vFMr6Yc5qwaAfnU9F1MBjO
18+x5c2dFT3FGEiUcSkBBYZgCaqGjF93letwE3KhhT6bHsqUC9wj+wJuOvsYH7ux
PWVCAVM9txrm1ECDG0w4/8/VhkmDJg/ddRPsvbhPN3NlXRHfbCBfWyLC8OONV0wZ
QD4CEPe+SNN+HN9DyVX1DjG6mJ8AzeUd60KshtleXWdPCqfro7JfxKW+hU6Q9lRd
WwyQmVZjZIN7nmpAP/gF+wO2R9CB/rx47OqChclAd0VngM+lmg3XS1apdq4cyoS0
5j4KPwmCqqcErKSlur8Rtb4K6A+io+nEi4pWS76m/gFqDSXrjP3/pFojGNJn6YCg
LgA6Nsh563pzEU53pEECc4dFcbthgL5Qd0SfKelEOwfLmJ2qjqDuo/yoSqZ2DexO
CpOlFog+Ik5YNyFx2wIhx2CrbG0hmRni8qS2PkoSewJyrm7YJ/BzTrzx1W88amqe
vDnvQMCRlYxykBE2pgmzuSvnlLgIJ5126jRue3wSnJCNOmX1/m0MyHZ3bhraAs3N
9tz5HSdoNW821IiEw1zJm5bgqYwjUIUCuJJBkvchqim/NjzqfvLG9yXf00chrdp/
SF2ySOPRmg7m+uIhCM7yfk/zVPDZ4VFEp69hQ78+8Y2aea0NOPT+YlIURr8kk8Bw
+vNxyHs9DflDOx3GGpyqSssnQJ5YTPIhczEeohTZhteP0v3EDz0dE9vkajLnwvGB
YANvxJXxCO8fPmoWxNcW3At+x2RCA8Zz3XgBGCp1pwUobWH8+wP7d2hrhwwLuGMs
DFSE+4/qwWhWhOZgeLN0o3z4s87dWpA9dU9d4pv/15sIgjHhOuJW6NofztnvdO1W
RNIjBE3nR69G0o9PJ9Sj9EMr+F4BNFjUsbMCfT1DOZbznZCyFkGThoLFWZIAUxBV
/oVyJMM9BDMXu1lwtsA1n9lVGjPWvSqGJpjzabzgZJT1VMk3ajw2gyS40WT11ilE
cEB0kB8l71YH0pMe25WRasps1izdAYU6Mk361B4evPthH2ZSQ1x1keTVsAcvwgkn
JftQr4ax78aOZoRCyLGrXmka4wk5NhXNVuet2VM/pCB+VdcpSG4wkV15whgUpPsw
kbJ3QOpJcjHHPjZKpeijh9wFUg1C9X3PD3lxwipM3u+CX6IpQJNpESJ+b2F2AS5z
Ea1e78tboCYHk6/tkNKqjg36++acfAobJgjhQxhPh5F87Y6SNMJzixG6YldJk8ez
aDF1TLtpNNrdUs8nPVvJqhAo5mCfZDnsA+rf4E7iLUAE6rMK+kvq+uhmkeReAaS7
o/o2GD0ozx6m2XKZ+I+jwKmYlfULLBMImDUJ/kwy0u6+jeP2M0dRa5DsH3s6XYpc
OTRFnr9Vjcn7JIgjOjrUYdldzGiFMAUPC7IWIZe1AIpY8w73a7VDMeg0XqcY3uQO
Re/7CbeQdPgNPjTX9sugVDo8yZ8lVV/0WG3hIneAlVzZ7iUaMqVcpDxgNummqLFF
ggEQn+GwXr8CMVZTwMJzxwWs0H+TGCDirrUxSmZefO30ffPWz/fBWr9dOwuHMq49
T28PEJLy0kdKWBkQf9klX995QLfekRVqCykX8DcwxSrdR2KCvquwqQrPNEAi4VNs
hjTmdWAhBUgqi3Ea9Twcs355bJR7kg3ip2tahEMcIRQAv1XqiWVZrWPaa2ghtQDg
i1C/Y+APXxPsIpl63dGcD4+ioT4DXChBXCv0uGA2vaTc8HqcbIhCwVbNoUUpp25C
GISOZOcOlvRfpz+f3gKMAMjqr8Gk5SRmX0znYqJuEp3ooOmTiqlgnex5e3LHucsg
q3I+Cxxmfh0ejbynF3AgU3EGEa6xgGVuEPXkhX3K6B+1cbWa1vqD75umXk7PAAbL
SIC3Pah99LJWkPVWV6S2Yji4DMZylnsRgyZLvGnac3LS6OEbcSwLvPBQb3DGuJOl
7rMVwy2BHZPy/l/2IQASD9pjdzdDYVFnCcpc2GWW1gLI6WC6leZGHKUqhO6t8CUq
FR46y7rrlZppR6ttoAYZJ2T8PKS+xTmP5zUrZxKnv+Ay6WrofnGWGD2ES49wsQHG
rrAJZ43gFGOc8KBC8W+7b0nPcFBvihh+1JXzIycsq8kGIwaB2KnnxJcF5jrCoaby
wKSUmW3S7e7SICqhjBRSpLb5/fSvAaUJ6wSE3AaqNA5/bCVFU04VsXxv7FJ6dzr/
5nEKS33RhppnNTlz4y76+Y7Qh2LKDtdpuVFqTEMvYC0mlLNPEjPl+xD1rN5dOG/F
q/68nLuK/UbeNwV8nLPIxN9DVt6u5KQQUA4i1jNjl0plHBGySNoq9jJu52YG7KzW
krFDJlUN5uf5GZjx0wPdS7QEK6jYB4ASdTVhqYUr59o2ToGtrdt2fgE5zkab2U1R
Q5PAhwdoFjYqL0gJ6AKO1MdGPQlxX5NMcUOwW2rMxIZ0FwnnDtqYzE4G/Zfjpai+
Zr5S0laFrtLpnmnlsmn9gNnOm+AhMLHFeuyhnJErh1WjlvOqcQ0qRyQz3vy9fTRo
x//RFhZw9RrSGdTRNEnMeN47ogv5ep0H7k9lJqruRGRSStK1X93/wEKC5h4/LMGl
6HfLQylSdbvkISV5zLngFBHxIqote8Yel4HL8NmxO9slSbKTLCxqyEFf6DFmJqGM
74gopbYv1rsqxi34qY6df7ETBRzwGbpSPSOZ3j7vHpXZNChG68z6JJtkNn6NJef4
+iA/3SutKbqpg7Bi7BLpVX7jz/ko/wINFgSkkL02udoDglQyAifKeaHU+Hg2GH0M
sUqNIoZnu0mGQr35/APHq2ljLr4VgC+4olNeeqdZ1yOLtl4sPUQRc1LnCIAzvmUH
ujirx/K7uTrwzgtEo5wLeL1EPdVGqIFx9a7TBqbs54OS6sf+Z5Xt/jaLp6dTW0TS
OjCFIi23ZnTrUjW7P12udJswEFPA0lnKymEWMfnuUpfWihVPKXBrcVcO8WRxwsiv
4GP0hg966KZvqOJcpJVCzreF22BJgTa47bH9fHMDexKRazGH4bKaT+pzAtKCCIho
S7AZI/MnrrF7rkI9AwstKE+Pe1YsdfpTnefL0PGdGNDsvE4Ov9lvdllZ/6GFQEpb
DZgNrL38mIn89pL1eZrJQnxsgNdIy3ZTLdCa1HTE9vvwKnlCrNhg5d8TD76jY2ta
Keo0i6IJh5CAOu98zuY7sOXWlPwSyqkYLrSaoN5ZOKVg5sdahfEseF4BP0wj2Tku
WHXJ1xljk8w+aQd4dlnuG5/zRbXTzKQffZprDYJMxQWXOXi7CvF/BkGBlyn8qxmd
24NycQPCTokp07JGOorx77o8TICSkyHxW3kbXFfGSjzfv6ODPwOHoDNpqFqPLRE/
VfwP9vUHsCYdBllFvuER/AWBobV17Dqod3jSb+5lfvM+wmn24Kanfj90GPn2ebC2
GuGwxPrkaFpDTX9FG0k/FNfNdHeDi3swDpgn+grZpUdkpIZ8tYmRRR/4cYN9I2j7
lFKoyjAm2JT++YQqe83RbosXg2uiSBiJa1oD5fpkWC4ZA3zQILh+YnsoGPkf1LVk
YKPmugM40WBOd4UjQuPwHWufVfl7QPNVV9QMhhzTMHAYF1JwFKBXKjt6vRNkJLKg
onms25fLRFR//nX3jkrBuowZDV5YWndsYhWK3bpcmYKUXeZ12w1F8RTM2MlqVQvE
cDo5n4D1Q637605m8MDjRrybQ1BOFjydG0aryxCSyWAh6jXeWrKUzIGXKe5qxgYB
XynNWjTdfevbSwPykD3jZVWJ07big+npnpkMYfX/b9B0k/R6VhDPO/yj7r1dyYS2
fMxU2/X7PtrLl8C2sowpk8KkTwag+wXzNHRVbXUyQ2DXihEBu0lpTBM7sQvX3w3Y
U8syVEDSqJ9s0x5WWtYaf4Wz80qTJyvoL3qszi2Z0IBPhCUl7vDjgKiHU64F647m
dbdFvnF9QCVE/qfpjlan4spEwgo6FxZVNcPhGaZMi2ST9GB5+8ht+Be5chOwvBzM
zI509VT0O5ywPbGRn2L4BMu0jz1ez7ZKBJu9dAgeNbtRyOjphqQo8BsBEpi/gONv
iRLS16Z265QrfeYc1btF6katw2Ab2wqgKoVadI+BX7FHZ5O8n3Vy0azeCE0YMw6p
Z1gut796sH2IESM0gw02QCOQXh3GvVVIwERFzaMxvadgD+V4UKeLu/3tML+884/0
3C8W4I5eXYnYkm8Lf4i+kx8NbSFZp4ESd3/FFSz2vxbWw+DImPngbuMy5ZoYSEtr
bFE++P8eUB6mC1ObLFhqtDXjqgix1cplSLyovGFRLb5g+SIQMDNnWChmns0TVPtS
WUlNvYlGoIH5xOcChb2iX9mcsNwC87icJTyccvGZjBxCNEWitGamW3UBis8rDnWo
zaVngL7qvBSlbntVEKMfv/R7Ty/r65PBTI9h6wrueTOmopHRt763OxwVpeZvgFsT
f5AN1lzraQjkn0XuRwEFXVf05EPh5A5rpZepGc0OsGjNbXy1e7K+Jcpp5BKzkAMQ
0vhP1D2Gbc1xY1FiEjaMKEnlQTdsXzZKhJcFHHL6t6F+yZ8t3NCESz3jE/3WTGxK
BwpWL3c/65sETFzcueMxvMKIC9V47RY/m9jTpEnetRL96V2z3KfgujIhHc08vpSp
+0wuWLLGr1Rdpn6hugx2JlxIWTsMK4D+qgVa0O5WMIJQHbHQpEjmSOOCBIpJj8OH
+vMEy7IV1RWi8FxK/E0yYJkeMGeN7FdjVUkTkH8pHllsJHUx85f7HSe/gNeuXR6w
7JA2YHNuUe5/kR/5Bnt5+rkmXzSx2DJpAqe3JJL9nIxX6j/BFuRT0X298cWahQ6j
NNBVx7PbBZ0L8fpBP2LsTvv0O2HVcS3UjDy2yjTShE0I5ziRt/Digcnrf3bWEsLv
7wlS2Xjwkoxd2HlEePEWPVBP9huKRm+TF27ZMroYl1kagy7ot/3+6mEuP03tw9fi
F0mxG/zPzotTcImcTh1ns81YM3FHfyE55CBwqK8sGGII2Ca8cprsiuHG0V8++vwp
8NKafq4OOzoRjlwkelkzXnTayAnT/6A6cU1A5WpOVWBZapGktiMVQJPwQZ0k1N7E
naEaMWceiUDfUMoCRIqBjfGMFaqCQfhTECyhUjuKv4xGqY7loBAwqgXychyFB01D
QUJpJuXO3xdrAsWzxsj+y3zFwn3lK59JTPzIYjZe+GpiB1L0K2usw/9GXLwgMwZU
MnpFR1gyiqIYU5++qGPW2VIk/l1kO6itOMmA4b18vLp0FrHNICLvcASOewweX4YD
++Ch7QOt+2vu8vceiiaPw/jwhBlSMCjK/Fh8F0tWvq3ZDcSkoHgFutE5VtILRjbB
Pb/EraqfUVws1QhvCvAJ2cKFbY0WpREZwZntr1wKPn6+eHBbplb8aYb49gYwee7o
WHjQS/wMMwRkwfb0RfYrTfqkrA1oSt5iwmTF3s+EJsxdt3wQXfvvjRjD3dAvEFv9
d0XMWxRy905t4loIinrjgdZ/JzEOV0/Tg+jdP9PpZwfDT6sZox773aiiD9cm9AVg
/mQOyRYQuWU8v7xM+ma1Y/PdXlVjzGHyfA37AlaLeh8svK8Cf/UzGBbCrLJsRp3q
U7atc4mYg7E8p/liYbX8sCWVa5aDDxi9FMemJsX3oHahvcO6MD/7l0YdD/eTEGK3
ZzfmmORg66rS3PccELGODJqgxGfJfsBGC77P0SwlIlk+4j2UHPAJUmzTcNlR9aAj
ZdfProBj68hovzgAOJMp0T+W4QM8yF5RYzIEWx+l8F87qk82BB+LTN1RvO3bgJcS
hWooTBWx6sAM6CJqf2FMwmCDar17/iJuabIn31soGveh2lUKJkJz1TDfxVL1yrdZ
mnp5JjMg39kc+XDPSYSEO0zxcNWARi1V89IleJyP4Pn6+NKcZ4W3/QPwvxQ7UpUp
zHIjUiQjyC+ljl5Y+DS6iPS2J8nd7mFte2UuXfxDdRbecFA3toOmiyfhrJyRcDOh
MJ+uDCnOtSE0OzogMAJ5wuLvjNe/A9BCTAISa10bJF+NBT/BuOeCns61jnLT9xmO
F6oFXWH0zR446MMWd4wxccuKnEyERg9EuiO8FaUOkpiH9LT8BganM4z7TEXfdblV
y6MNWnCVlhP4NAw17BaRLwpGHLFJDsgLmhFarDrG7bj2gRe7ReKw4AZ1poq/UUor
en1PxjN4wVfmuE2n3YYdimXTpnjRx1ovf4Zrd7MMNUVNt7k0C0GygJPhfLh43Lfm
VYLLGOk9ITkYcPYEFW8NXVIWM/W1MG3NFPHDVOxN+4nUpZsJIo5fYNfguOHITTAP
5nMI1vLVlXFny5j/WsZZQfgo4roRKPWqkFI+E/r5k/R+ocvEbi9NjlRgSYTrRNFk
xvKYHhaamxfpyIi20N/m6ulzIBS26undhjndj8r+9tfJF6aGrsBu+QFNSDnGM0i+
cdOi+vdVVayynt2soqoXSfORO6bn0vouEoAnW5GPDkq1D8RnzK+ZYP2nwiXqTiP0
GV43jarJBVtiQb2CXBvNKsiscBdPQLUQ+IynPX7m/itjWTcJgF2jCiNlA6WbTvkt
/2oGiP2NcOt0b79vr8mRXYZ1/PUNf4vk25QH2jSPFupfSOMZhT1QuJziYWk5r5/8
Gl7Xm/joZzvqqY596cXmDHY3cKLOyMb5ugvu6mPXRet8Rg5QW50stcLgsEF6BNNB
PqnxmDhoaCr9cqzTvMzNPA96NadBhBiKIus2YTmb8or0v5260LLwdVAQq7GqyBxy
ZUzF8NQsiezoSibSizNjP1a1FS1tiVKnekWRPoBLYVfQtGbkilV5IyJPgACd1Gu8
FT+xAJTswn9mnk86xsPSY3xvhPuFdc0P/6LdYFPpffH6GaQh+Uh1bnA8Oszxq7eT
VYx6JRreCGUnOBRLCxfpGJ2vlyyPFJ6HU4f2C3zSv9cBByU2aK7C1LAuyzrvTkvA
i7ADvD+L3ff8ZK8U3bscmN77JKNovHVsayr/wBNFmbNPAt9lHuW5sK11TXXMuBnh
iVJWfZ5idypjRF2OCXX6gssRCKgojGRnD7juBKxfoZmaTCmJpB9CLmFLIu/7Cxtl
4O9BuKgAzm6yi2ysWEX3J4qExycPTwJuw3h+tcKfgpq6K3HmmIWPvqbUWm9k8EPT
4Y8y5pbnnfUBfRsd2HMl8gjSK+M7Aj8wf3umQpawJJoq7C20w0ng+0DjTKQzDIcb
j3nU+nA++VVEXVWU3cp8+3S8/s79L86KIYIvXzhB2Vtu3CEH3moKksEpvPwGa8by
8lKXaGz21oduVuX6oxvJmb339eeoxEx3kLQ9s/v8btHSr6WI+C6008JKEzOXs/Lz
0j/clyiGce7e+5qB8lFWQDA7ain/8xCCoJsGZ/OCljhMsTRBEyVjruiApBYzYfFV
FI0Sw1FROE3LcIiGkr1fiELS9Phkf05g0GR+LUhYdB9maUM3Unbuwpl/Q+77ytSl
O2wl9nb17lZoPR67Jm1KURZuy28Jt3X2rSsYR3nKlESootVKzg/JCjTOJbMjh9Fy
f8bgps4PTEh6lsFu8q3K+xwfe/h7t9oJ9r3Vr+mtVjUxN72JxU5tC9N7b+bb2F/x
e93jgnZFaupdodQIrprKXIHhMeJEUafU7LuQoiOowgWLYx9krDWJXDBSh+n1NkFN
klQ3H5Eb9Q88FzIPNhKMc3ItuX1eDeqlc9G7Fg9cLTfqf/MpU5an4+plm0uIUVUc
UIboqnTyNPXdilfi4LH+ImbzfSkZJHKYuvk0blyqgeHyAqt3Ny7nEBZ6EEyCeMbi
yQJ4MHHLcJpEr0SI5fyYwOYPj5tReNyMs4nQQleqrYj552Ve8XXNFBMkY/uge/BN
vRSA8jLFPmu/0gQBeFxV4kMzkVNvZ6zxdrw1AqXtcLli7nUZIvhDpsF74Tim7Viu
Zzyo5JDhljEJ5upr/Ke3TtLkLzl1K0j0DZupySxbtYipxU7WTmcjCRnXfiFH1eZO
n5tp1bO4GGyiBOmp/UdpwI5lUaA2hlYBX3Lw50N9XjwBJnu3/LXoZ7nFZjlHsAFk
lxrs6Q9d5fvRLLuEdTiflkSzQOXkKT3aEVmsoCXBlVBHsw5+lJIH8ZZROyLBK4EF
6rll5xgDDoah3o4T338yNZU4idKzwo8gR1oK/wN4cKMgg3JUS2dxdyTXSTQUTkmU
JE5uEY1j9bOLo80XAgGkSpP1u4NZCIrAIldifOAbIZTpx1/4zvh0YWq/aUwhzl8i
ilysxnqCT+ICySVBCUEsr3xvM2wCigK6TXqF44l6/7WH8l6nTZc6tlkxjdfz6n9n
5+MkvdV+XAjkk1v+1JnEw+Qqw4jRdArgG4SfWcGO1x1zgH7usIyTw9gnNmfcDjeH
ts4OU8eW99huFKOZthBm1pb2bu1btihXo/W+vRAPLIwJTxxrF5kgAEyvBV7mfDRE
xWYJ34nyiTuFlxPkLYR/P53RczPumOljAmEE2rZNdJ5+H1fruLPCeNndsaLMmBDj
xtVVwv217r5f1ZHKKkUXIe+qk6tHq1P8mB3jTaIRDAbThhzgCzUUBtNmxxzN0002
8sK6TY8v//zlIJ2MnuCP9Xd7uG5WBQIFFS+pHrAFi+BXlOX/wyn4itSdEp1osa+X
WjGRC/A5UjgmY1Ir0gLiyTGKv2AsuuYT+lWlsBkbpXC8cO9UO7sO8ivg3oq/Acp9
RyAfN9uCUU8LKUc7BP3Ho0SeuVYdya0lML9taSHOAJmGij0SLmWiZ8cKyLRsqOZ5
nitvSH+Ev0U/Sg52I32X4NlU6qwmuSdopYKSVXgP0pG/VNav+pi+lOZ1Lzjk4RVg
vQCTkPenmPB4CYmlJ4P6q+7koxJvyJgjvU64FnH5JpInDoiAwnsbU8b/PLc7HUxY
xeY529IYGJS2Tk9bgM9qiw4nIpNv108bhkMKqN7mOd+OkwVP2m/LrEClE1Hb1woc
kjEZHJZ8qaNlJcNMfK31z/AjgqH0wRh0Dse/bnC6NWQLZ25Jvrd3MAARDYHAVfQ7
PKQ+DlECBK8kywmj0OOaZVER41q2bLEfy5CLngVe4CLYc8kaCtqydGddHCXgPq7X
PE0r1rS73yXaaooX/ves81b45EPxX5C0IgGok0Um7CXwha2FdTiz0vC2M2mwZJkW
C4ecU3iRE3tjdu+UlxaoN/E8xu3MoLUzJ4BZ71n70QhEildfxYFmoawpxT7GewkT
VBoD9Q1ENIYa9VCT9zLDMy3ogAxaoqFt5hDrBeiR/T/FRZYJ1aB3yM53BQyqsQVx
W96PV10/PFYpI/13LLtIc1epEdVvZ8jLN1j9B5Y+p+mHq6z0uVovWvla8QQt4eqI
EqgL2Fes8MAHgkyH1/JC49Azy3ysbe5CLQY0qEF+VQ6VdTH8M2Xnv7AsC1mM14fe
/xwmnHT0wH/4ThCYv855wlTjzq6zAlW61JOtRt7M+fVlFG/MSDo0wHmH4LHRheWk
MQuurIyGJ6OVzRpSb2J2skHnUQ9FRjcunl15nxtTUxDENUYYihcaXdZMa7hezaM5
8Jq9Bxc0Ms2wT/kEjLVAuUnR+wMYD/9FOgRaEqCcZ7WyCF1xm/1z5jodMYGa1U4y
JOmYEODFhZO6WxLqNFFxqv26N2quoyZw4SMUFCDI9gE+AE+o1x6kTuLztvwxfrpA
818ps5WSGTVNiPXp+LVDmUrkI72Sdh9SAYvUUS7Wd7UMfdQ1HpGfl0BHTyewdKfh
MSP37yi1e6vzUb9jfNZSeiFza0FRcznvu3DykH4ZpdAYPCy2RWbwzP4ioISpeNDI
JUqH39mRQ3D/Cz21+a1AWG1KbU2ZRBjvziaZIMV7C5i9JHKWbDYvySbvcAyuIshq
8UDT9WN95gdRbjDvUeLFyUnGScFN0OVuYV7wFLKdPuc8kLbR1uXJbOfTazYnUA7U
PD9BMKQ2htKwMh4P40AML694/RtPFxqCSrQGB4Wo0CD+L1PAj402kwGY7y2X+D59
z7rxKJ/L6q61ywvJIdS/R5X/UyGnvM/IiFxivC2HDrPrtwnb/RXD46JH8z35EyHF
yhDneTRHph34Yc//pu9dPd8g8ECL2BbbmvQgCvvEftMIM0JDKrpOoRFmdLf9vIha
7KTyWEkaTPcarMJ1Tr7/3B+jG/4BRGIj4k+Qyyuj293iQpHUBD6KupVe0t7F/Wt/
Pk0kbpEgJTrgksF8Uofq1xeqhgqZhz1uag/7fpDzPqAOQ/ekytZ4SBNkxmPeo3SL
1fHnKZKFiUw+8KdeBCps5Nz1PT1BkVJbLDEJp1zoYsVHc9bIiSky0i782Tcsq7PA
soNXDjjCebF7k2W50WPBONjw04xFbvFcS6WTL6HItAGh0XPIJ3OI80Z21Tjc3Nqk
rIiY3nZFs2AR455yDhq1U3c8yEjgkumHZOft3nUEdNtiECqEVzV8x+SliJ+sHksW
pwX3BAcMBGEUVZdYhxG7GPc/7z1y3JQKv9IJiNy+muzz6KQU7yETpYW7ZRNlkhAk
Ypx9MWny9c1hT+wE4y7XrIP6o5XYV+Ld6ikno8oimxXAjAuD/xAHLn+Xu4n+/XxO
3+h4FodxSK4Ez4byfW5vHG7k1TO7x3CSamNJPkyXmSPQe0UBhnkKOrOydGLZJju7
bp+J+gZdxcLkmmQK5DOAdeKlqAQAKILBr6Z6CyLl1p91VGLaLg10YF5RohQmGlrR
ZQzqUpt2P1Y1l82YaFMo2FnKPu2BRsn2lAKdWyyc/rOd5kC593AeaOke63IAGUKj
eTXZzvMRtdr1tMncHW1NBsYi98sLdSF8FjeQemk3RZMOVUUYXeEcpMLn1Wo13n9v
ShJyIq3k9RMZ1+Wa1oLU6BN/aaeFgUniRLjGPzu2D5Ji4v1UgxPJih1CSTr/8+/d
F0+b+HqDuzFirpDXCxVUrFedt0f448dSWCUCdACOhPLHUFN58HvRwa32Nz0VbLXU
UKGLUKpnIwkRL2RaCiNDC6Zq7s+l985lKu3xAMSKPdpFgGnYe7U7yEd72i2vFxPk
eoOwFrDd1a5jMzF17x7tltjrVw107svoCD8UJ6j/YQubbs3U44b0WFOuipZnR9Yh
u/6wk8u/hYa+anJ73BJcEKKf001v0JisQGIVUDbMdDe8t4D0WQIQOfpLzHlsujO7
XQ2Lw88h8fazMhkJjgys+ZkTpLs5kiUQbiAmjjQVO/2MuKb0VfLKHb9DEzhlNGYF
w7Kf6s2NnoKdPesc57lhQD7vyv2LAbxW1pyURUxfS1gZ7SMjOcP+TwI2MmegTId3
IVdGTwpuTcDEd3DtfWY69Mp6iyIbOkgGk9ZDg3vIb1bTSMposq8BVxjiRoWruphd
qT+sjxtax8BZToL/XBzmudHdOmpVT/4y4SnaOMLYtXKk7Tom9h4T8qK0cO/xYWjm
cGU//xPFgdSfzAC71UNC1hUMRAZ+OlSzwr+cliFfMI2iGcSPOAZ+XzQfIgjmXc7b
1Rrr2O//kColVyyV5vOJoxGzQ7sq8fNW5908uWI1/ygPSa9nJuUbo+0+2OzVy7D9
PzHlH0fU+nIt3ytxOmiCMYQGiG5eX520P+lu1D30zQYnfNYSk7x64iZl4SVQpTFm
zXw4ZqZFPX521bSvMxu3Y/YcIIFqty33dyT8N4iv83TI+axX8s4sm6jcnQ/6POpf
uyw5nIfpa1cLgGk9MwlHq4G7TwwKjoYDLLDk/wQoSUIy2XqaJlhvQuq1qL9Ncgkn
3IUxvVrgOphW+Ql3ZELdKKtotBJYOw2oX8r+EWHUMcfUQZ0xadTPKSLFo8g5MSDm
zgSC5u8DZ+OxekSQudflcmA4h+TNbjdEYo2nLTp23hIzHDRWla9V8RrGoExdC8Fl
LceRZyK0NIHh/JIom36G/9DBkOw5L2lo/+0lxqe1rQvpNAzwhaGmrpsDRrL0F7rv
LcpVWFFjDnkC1CJYsV3fm/gF6c6T+xr/GqY/H0RaF4K/ck3o/ch2xOafr1cn8Cni
A0YeGqnSgugk0yXVnxKq9IBolwxxjzPuwNcOXl1lSk6E0AqzZoOTUxMZgvoKFusC
uVoBpdAnODn6Ag4dbGlmv3adUc+WXhaUd3a1IWzGFmbrjUSm3XKU1NZedpVcLtQR
YpDQ4R6Bq50uKKt+xo79MDUGNj9Diei34Tx8jsiAXiFnijtgzINFefore7oAI+yD
Mem43ADR1Uas3EwpBMho81CswSzsxJS/oFSWeA+bPyv9o9CGvWlBfFYjWOK2ysIq
8lwDhR1sKp/hCQFDhcnJCHTRpsx1kvHSeQyEZcXBQCT/9/WmiReJGn21W2ZJyeJs
wD8gjIhRZkR2+t8+JRhDOMK87ompUfupyZtgEQoL/dSSGRoYbzfN0Q2vMRRaxUjY
kNgebxk9f4413fOXqO8C8FuyzVi1JdvXPyDVcqkU943D7C6bBzoeNKUW67PLmWfU
Gna1Tvesk2tOwE2gK+6XUQj6zM2hstT//dggFkuMkjsnPioOUjRyKuR3Qvhal8qd
VX3j3onRS0kuWh213QYUdoGMsK/y0EqCpzMFeYPAcqtwmvX3w24XObwoYz/118tl
MQ+dhzAdlwav1LL+cyk7Xg0bO15s6noJMEgCOkM6ssGwx1oGmuCLqIDs+cjGOdJU
pO4eH0eVtXIzt0mlQPDCOIvkcIiOs7iWN8Y8yfvx7Wdl8UzIj6i4aH3keE4Qa96Q
uNDLA4k56UiCOqunluCtjS2GJ0hqi5Lr7hFAqxrmFqmeRFOJ4k0cRHpQocdKLCe7
1fbvVgCTx1KpzvZ+3uputMzrdbN0JhK+RPyho25PcBwHnsb/6iuuBdSVJdnUrRm4
Dpz8gm564w/7gebWlunkkEeOwxULiQuOKFbNX8b64ZnUTQR+rE22AD6w/8MXg1aK
AV1Eue8bSA4jHhy8mucw5AVTPeDhis6aWKe35eALqpKj9Ymia3xnXm7b1qbFLs8f
RvyrzI+fEbLi4qME/LVMGUyIH5YbMfWMBHp9DJZPbPaj0itj8P6AbN/We7z5kjMr
/Z5ErOALysmEqz+9LwYfv5lQGgkeS0dbieoVh7u5mHuNHh3aWSb56QyoK0i63IjH
pIhWgk8n8+EWNYEszm54IPwNCFLPOgN1jqNBtO1WnegAqTfdq8CLCjmThnmqqx/8
CEhHZG2OwZGwGYcl6G+SHEY/dZyvA3RcJTLTt3xunzsFCuRiK8IO8ynTMs8gBQKo
2/NUFRAVieyVKddWENVvo+SlBA+SCqvId1spCW5JEbNIqT/AMb/nLmOaEoxfdDGk
2xXndPC7yGVWpaTA5x8RLY5uG+XRzb99MhjZScVL266QTZL8jZ0YwRNwxXdCD/cm
lqDXeGsJOYwZpttjqwImMT6wKWxGYNeglISGF32xJfm474tLSGPUpiD3oAVTLYMF
U7FCUex4iw/tNuCiG2NwDJ8Qlf8egCWopT3Ca6bMLd6+v6x4eut9ISow6DlP+b4T
7a/jVWJmedkeFndLcvqq7dk4dt9uZ3vq+/GL4El/Ehb8oCaobd6mXdSY+oUZWDq0
C87DZlls5OIGaGqLw7ZQqkzdrioVJyAvmZKX/NJ1JYfqunmpaZWsa6s8KNnQKU7Y
qTD/0QabzuMwSl1kXJ7ft+Rs7oKKHpV/ZdobO6tGf/QJ4Qx6IBrTvMo8guDA2xa5
CPXfe3k0FEA5LdGA6SW8qh63i0dk4jK/tXso+eBcYGM89H2ZCRK1taTLand4VDcg
q0sqzikYfM7+bMQLaJLkp2UJuWpADZUNjAVnvSxB5IzHy6Dqlb5KVXyb8IxzEdpV
/rtPU7dQf2TE+TemNSl5BKK37kQBJrDHh8WFTlb4i7TbaKdJ5mjFy1vKK193xIOK
YK+yBArb1y0ENaQXEUTgkFofLSx/51trBJQ68+vh3vPdx4YYcLEgpiW1a11Pou2e
Mat67Wnnn0qaGxg/vgtYiYVeos25AJCOSnMwKX5oXdk1OePeguAbp8/vz1vPMpeu
QKbm3JhpdyMkCIidcZBWPHAUy7HlEZioJHbl3PN9PhJrD9a9X8B3GEHxjmQ2D3nx
oYfgj22hqWH988p7SxPx/rNkjv6MfESU5nlAY0T8PAm5q/Uf/dGGQYzyJQ/IMopA
NaU9F+T48OpW7C5SzNgxJQxJiarm+qjqW9aQkQQymIt9lEBKR1gb9UwAMwIWDyKl
tAW+IagF9aVcbR6uiFpK9IKuqvrMlVPOHMwNvGwg+iZRgZWxnlYUouBgJUPoWQlT
dDEjPbCY4OOkxGytgEMC+wH50Aq9rwpctfkTx1uN8tFNu1U4XE4vjFCozY4luNvd
vp0Uz0ZR0emF16lt5IMi1oySRRyKXMdi4ib7frEY3HhS/vBEKDv7mvHHVzKnvJL4
u+nEoyscGTi2Qh8hCv09JmFfttdLaAiAMhlixDeCAlu/Ir2Znch1uVFGoFUaJbPl
omDKe/KgyQxioTEqESyxz9YcBCAV1mmZLBxbxakmw3mJGrLmZrOxbBWAIHIx58Zl
Zpg9zeuNFowJM864uVKzidpf4wSIXcZNDNWk8rRygDFYWlvH9Fycy9aLkZWfo4Jf
ZYT4j1Wkgwr1USrgJWxG0znn7xuLRvykeeU7kRuSEevr69JubPAvqi5OkHu3Od4N
83TQKguelPeqfQh7g1s1tmewmGJyyNT/0CEL+StFO586hYQ1a6QvynA42ljp2GR3
nF10Frla8daqa7n5VkCD65vwuP53KfQutbs+un6wS+FzxD7IX+sBY6nawWug7pfC
i8KQ4LLDx5ga5bSg0tLVV++hqV/R+8lsJFOv3DrhTErhFyWV6XzAnPacToRELD9J
aHiQJg0zOuVaK7YVyRMSiQS7XaLsIDL1U2nnJ/gBEEgK+XRs+PvFjBEY4mG2/ZkO
UuDNYFZVPeZPys0IeLrnzvOqA/SohwVOUx0cM0eACN3HWtHCGeEHTNxK4Sb9ihMI
+EOmwwSAZiWmIRb7ScssIPQfgOASnAZW4dsyFTvHXpsUuVnO2I1+n5t08Btg/78E
A1vjcbb8jug4DVqktaZRcYK8yZCaWIVEIb9ywKLPlBTzx2vdb7HBnVfeHzHis1Ma
qA+wwBF6DL5VG/1TwPghwyQmtMYpgMM+tyxr2tgIoYcS6nkG7aHwuyEdgygfn7Gq
FVCQbRoqoGbMwN0aCRti/6POYW8np9B5tWW1ZoZYdVzxXDAzuHEZ5K4YCdvv7QgN
4TnNVYR8Y2mBSPuVyu3ufjD86p/Dj7gRMfZQPZTZYZFCd04o6NNGkaq3Kh4wSUjC
PV+sCwNYF0cRN7KWlPbt5s+IKGPwArFPnEUpBH3/w9A11Woh7mBd7y3D4IfrglgE
QhmygJ9QEhQDuJk9ged3QVel2BJKo8SgLeh9yLbBnnULR2J1hPhdlWyS3P7282MX
3ojC/sUqBHqngYZIPGbCgrEDBFSEL9ExYV25/L2aOk8Icr9y9jqf9u9VTHpjrGr5
Hk9+ma2Y/GGCd+ezHoBziEkvo6gCDUCrtUY+PCR9wxg8iLELxlznP/CZQ3IhtF5N
A748xsy7m9JynlnKsH0JZPhrzTrkhje/hDMVppoxWjlNZ/Ho1hkqQPQDJHjPvDuK
ZiY5NQiz2fL0TkYineonDg7l3hdeoJmH0v3hHOgu7GMP1q09vJTmHiRY5Wc5Sdg4
q/iQrkfdiY57inlyC/Iy3cRDjxbfZUPWP434ADR4WcRfi8HLWSFQ60SUORQB3ZSc
Znj3JAC466QYamLXteq3gZnGtoDwif6/c9VQb2KaepFlZSs+5Oz9sEpQSS1a+BFr
wM9DN9p7mTKK/cUS9tEiku6jqIIqjBtG4ZnhMyHLFrsWphzCiV/1tM2dJmLdbxmD
F2+o1kA/FSaIH6/bec9rR5AZgmn/CInLZh2GgbEU4l8MVRxhaXoJe2DdDSINFPtX
XOsHsuTMY0RUTeLrVhqC0jrniJbf/dote17oQbsNfvUvZuhifttE6lMxdhkDvAcr
qnSxFHVdzt+vHLmR8RbcU879LtKEoH3UOXvPdgxN2ir0phCqa/ZgZM/2isG0BAJT
4qlPaSnCwK5CCLY61Q0mgdtc5aV5nrF31T1TM0FpvJQwU45r6OhUfXovU5KfIw+B
CUGlWRPgLeuUhK1hkNgbsPhId/XI3MuJPWIiRrg4OhqM+h63It3CklxVA5lVJj2h
IY3lLUBUlzi7P5a1p7XkyaGA6fKcMJaIASafPKaMcDuxmoWMhiBRZL050aLYLZ6l
SvLkmc6Zcg8HOkCI0JDAMn7NLgtG2Plx3svnyuZ37uKVK1B7XPCbsiEQ6waa7Sym
/uCvPdggpGEWS3s9MluC5riPjdbpCQk2aq8PfD50AZWxcS1HHdrSZNcS9LXdlSC8
LAtVSvAWz0m6XuK/6yu3lt2Y8ylSYUq6lBNkDIBkatvzxhIjf8xywomX+D/vHw7l
Ec+qdg5Z0au3SwEiecwfJ/V9IGFjhZwYILa0WfjlSiHNjISAAzjdVkoB44zwA2FR
ir4Bktws2Dtc+OIQni2N4F3JA0Uv8GaFncx19tx33Gdz8qcNTxWB3N2oe1m9a8+A
/ppdhh9XfsmqzDxazXkW/+goUTsqh2V3u+fopEji44KB43NQ95AcgyE59yeQHbFD
UICoVz4R6KGAHwP48Zqmbw8M+6gP6K6b/6g/pYtFLkRg3x9uePKOwcqdsGtzzxxU
YrzQn+SUrRtj9UsklvTdf+rCL3sXyLgunuHgzNI+c3CRmouNGyjovMmoohE2WCD1
Agmyy4rbxiuBOgiKYj2u81vnL5VZZFuqNJlStOu/EKHVCzhho9Xl1vBsi/Y95fQH
G/40KLuTFZYnLTOKJ0VPV+wmjep6+Avm+6jImrt9ds8tsE0x9aPoo2sNxsobAFC3
VV6P7LOpgCeiRWBaJG/dVl4hdWkuUz9qRqJRX0a+C6TddHUzclfShuOI+IecMZlu
hpPMoYir9gHGDgfYvbAD9XISEOikgnQHFU8RHTHLPbgWFAeHtNUyZluabCKpcxs0
hBYr1aRuhWmLidJ8wxvFggwlNeczcwWC/NznLtbsCg8e/JxS5VhPPCHav7OQEPff
tyE6g4B1XukSG4BicEMKMWkKDrZMjILuVLSM50VGHDiHmk+7exAoyIatWG9mV/96
idfY4nipO5SPeYPIksXO8H+X5kNbxCmxF5zleKvPg0jUYBTk1PZfaN8FREKcg5d9
qhLoUR/aW3ofBC5WzbIsR5WkaSW+lhMi7GWn/355vkLzuRg04gZRfCplWUDlufQB
Pn1kvUfamD6wohu22yG5WesQaG0MCTOHnCUam5gfLzfiwQlNiE6EsVzIBfeR8HaF
1MtIkThi8W/o+Tz+oDgHGfbQGSTTRzyZlqPHn4CIuts5rusfe6Dxi1UZdvKpINE0
9Xet3oAZbYk80NWL05IeggyTbvA4PaZmadnGNywrhZjzI9x9IUG9dORO2Bpb+p3r
JjWEI/3N8fuJa2vQn853B9V7lngEyeHxFpXJPK2tiVL64whqUqCO22nT8h4mbYEs
N9j8sYUGXkbK8U0h0Z9API6moFO+qTjnhat5njBU7eOG3jp3OGsmZ+nVOH0Jz2Rf
V6p3ljnCK8e7PnQ3eBIitpA5vtFXTLyh6nldOArJHYa61Lzdls9EnfrIZTj9JO3o
LqkIby76KBBdcwgriiuGh7rw/Mo6FOlCR2eb6I7YFTrenLXjEleMGJjE5uwajloS
Hr7puM3DTsY/B4IgVQ4Ix7IEsQ/iQAFM4JotdDTNWy6BD4vE6WxfMceo5fRNuxPB
sEaTsDLsPU0MLhE4anFp3lHkVfmkJP3voxpMUVUEsPNh+15CkEr5k57p8NzE6JOJ
EJazTGr7l3v10qpcEaIDHuS/9Z+tyhDyUTljiUme8XO5JC+ROZrDISnSMuvckjzx
kWMEiLNUcZplvDeBw59ITRRzq1SppIqq1WDSJo4O+zSQwx01Io4ZhSa0k/85idsr
9NA7sONJq/5KUA3vd5TPYPvZwkcX4ukpgpZbSbYa9bv7tQt33BYZwG6Gf+2dQokb
kZ6HpYXVeGUlXmYrDfvOrVfRe/qTu67oEpEF3u4VfPQZbZ0V1D9yIUVNS2q0paEo
s9CbC2Qy0bUT9haUGIbDTGivkG/1cyHwgpo9qTMyt0wnnaJ6h1yRQd1QKMEtaNBI
mv/IEx1PWrrSe3wUWzOMrbVJ8iX5sl8aeYe/qxfKsLJsAFXv8CFvANaTLK/ehn+n
PpKvCejsWFuHkhWPjHsx4+T4onyWmvC3TzTNbz+GbL29+xoblJ8GRWqmOMkhIEdx
PWibmH1NrrFyP4BXwYTL74MF+ZpGRRYr3wYSXiNvMv4oAYrSo90xiUZf2ckAut91
w5xqOATvFy1Rqw/eolTJjIKM5NRiDftBGyIrrFkdxD/1+mGbenLUKlQ/UK4n76zP
lS/gBfK1I1mJ8MI3wI9tB4Obpe2z7YTRJ9nINiG2QqSoCW/yi5pMDSRIzgK2kKC+
zFdgJ8LOuM3KQ9tfZvELyso/ZH4gIKuolKs6O3R6uG6o1oyGH3B9VOeJQsNPOBGW
PrfUXkbw2nYMOoihpQTqhZq+9i5JzWcfktvWJsMzbm3tuvifPQlpoA352P8xMAia
NDNGOBA19afqlobEWkT9jZKmFdT2sXvK1k/qtVXK1QCP+uD/g1HH2tXAvIqoPxYs
vvETGKxyi4q1K0TvQSDeyqIjFnXpj8XfXoXYGaSBLbZjbMzv1napFRfCmafKV2AK
kRWUYuFOchw9xD48NNoSv/25d03yRzg4qASNAEtjDL4H6YhAsbLl5Ne+/0FUrcoC
pRSNf45gWNwSDSEGsUdwOj4sjTNEF3R7TGyTlXdpYxIWY+G5RSSPHe+eDB8SHCLl
6FYxM9utiYHcQZMqFYFndq91wZrDLTsPtRXq8tWzvjKfUVp91jbKZu4YkK9e6UPx
yMmNkVKsb9mC/6xvHf4gnzaFC+6jLOiFuIoeFbCT959CFA3A7IrqOe7NiUap/0Vc
wKsjpWFse1IbtgQubFiGopFwtScEitsmElIccc4i2b3IGx6vD4yuJfb+5CVXY1PX
hKsJDCj3faImqfKrALhCVVbgoBE5RBZ9Ei1z1zwN3nWas/T7p3TLm7604qxQowwX
298/HoThQoWjH/0TYu+ia6AWwYaXTSViXm/oCxuMJIdDowdgl4E4SuvJSsbDQuO9
Wg2jODz4xhsQj6h5HZeKk7P1ORQ+fe3ErhEh9XysI6KH0n4QdtKhucZmxK2dKTTZ
m5KbKl4JwiOppw+wYzkcZnf3F2cu3l8VtULiOMjaznjFzlbckNLYlba7n2BMVa1h
h5OJs4TCVb1NkH68s+donN9YEN8xH0/VyPX5ZAkbklc5BHhjmMc6Tm35pSyC1OCi
NcVXGw4yJ8P8qW/WlYOpGm63l7ffiGxxPI7WtYP1ZkqH/83XCfwlnz0AmtpmpWpp
RQq/7f+VYxI9FtdZ0m8QlzaRRI1a8zNb0h6VbUAt+ymbivu6ouix51rz4WYYsspy
FkQlNZXLXGmyNi3omvq8d8EoOuB+0SemJJhbd+VZZ83x/i/vJfYk3u9dpBJ+oPGF
V397uOplr0Yktsh5XBbV9YhJRDCrkArLm9DDqfwU61qKQygER0NjueTna10fHdkL
dj8iQZhmiZbor+FRlmMynR/ZAJmAvv4H4XdqlwQaEzQth+DZC+RAkupQ35avMglY
eMrVd1qA2BsKjCl0vrWTuugB0tRHiXwPRZZASAxD3WZw6HOI2x7Q6exdnlAiNx/Z
/A5jvLTrRklr5Kry38nf6+51OeOxvTDmTsaOzeyY+rEX9QrcsgVDVqzkN6yiBEf0
lTuwU6+ZTSRnziXndZ8/Vi9i+BgMK3SivrYaRSeG5tsi3IKmqGt3gWkFTnWAEzEh
e9Yu2KkZRCLJUoBfpKp6bnj0+YKlJlBe2EMJOR+l+MrqUepDl1Wue8nTdpo9ypU7
cxgJeAoGtTgBSbl6f1LEdxvIGA/kvcaCwIMszSPrQJ1VGIUJkZi5vShT1jqX8qaT
ekZGf7BCvspyucWpitUFUqI/8tUbcnovPG4kg/nos4nDszLyvlH7wNqniJAJci29
D0CqqRbrYRLK7KaLv+IyfBxGUoak5NVctCfzdIkbEiXASMsAE0o5IzfsIgoGyHTr
mY0Qou1Ko8TKXKUOE7bBvzP/GyaYuxgIC/PaAK+MlxPfPAmnk5kpTLlO95Rsta9V
hbq+hb5R+ZGMr18fPB/zIbTlKk9tyLp99mHD+JEKmmXP0XicElQ5ZJrp/KmugK/c
zdPirmJbUaBhwnr1JlXwIlwkKqnMtCYfUGwzVZFlBvnbOVGuCB7zzOV78ZAtJnlI
ZyfKdr52ENkxPREYwoO3Ux0hlyFDwQhUdADj7ed2w18NGNCVsWAcbckQBiRUoIBW
gvOlyzhvl3E3ZScCu9BhauZo1lzX4N6wJjBDNo2y+K+BNSFZ+693RgUMjjhSJn29
9Di8qNHQjkZ9HjzMwpywIeTVyxjbHYsrVQZl1qgWE7Cd6IF1NW7VDQ48p1Ttqys4
SXVeNv4vN38Qa5ZDOkLkANiryuQTap59p6HRmyorb7xYTNlsgjCXlLIqe6UJD5UA
u3/VLnnX6rKg3n3mU0KaZdkw3WlEaIWZ93EE0QJZbsvZ5Y30YXGk9+Nbbv1uMqDq
CK0+k32hsNgNZFC3MoY2bU0LCq3AQP8wXZZJru0HgsHxp3IQSjJB82T0ose/qKir
kLWiz988OYRZqWqFVMbf0xsT48qWlMmTOdNeq5u0lNsVXAR4/MBrSbYauH/gEy4q
GTHy/AJEv6cECRPYFVYdBdo5iOked06pfrjjaQcpz2MhvFFXOlmdw0OsVwNKlaaj
4JbjrReh0qe5VIgpJZc2GuqvsQXxmFbqaQyFVXof+LlaZnX4aNBatv1LuiIVyW1R
tQlsmYN4aOLxVndK46o6tUQVmy+lcV4B2kZxOpfo2l71VFIwA3ThPDQiwkViD5un
0f+kKq3IvNeDdj5/635Mqx40EOQe22cwniVzJ6EUj5sqneAYDrOqPDo3yCPJtpUB
lG9jf7ncVQV2LASzsoD77Pm/oLyoylnkuqBmYTw9cBaOaIw0vkR2JyFyxDbyeLBM
3pqtK338k1aryQ23IqzR/rYMIAK7kPdn8DSBONHCYHkXhJZQyM65Avlq2hQfXwRv
4EapV4FNl3RC1ww8DfyZr+zaxi8TAP6W+q3j5jsyLQU43IGmWUJbZPHZwBmf7fDH
iild+04TdL5SXPSSCq0Qp8ZCeASPelaeep5/X09ZNn3XK6ecu8DR7PJwKHrHhDQQ
6IX2LpXn2Rs+usrFXvggdX6ynlqbob2aSzcOoZzaz7AT0SxNUIS3RWhzyYzOrNQo
wO+30sNnksA0cKFfaB87CawQ6nCEIJ37eYxuzYFFmmHPAAVAq2/541RoaQ8QpwRH
rfXQIP/BNtuL02u5gXTILbKcY3Bu0/RGz9ZqWCj45NOwF9Zmzt5xXZ0g8p7O4ku8
5TvBWOIX+IzJH6nTh7FnmhoRKAkVGJ9D5r5rK5Lq06waZN8CZT6tpjUA1Qn53e1j
cs124o7gTRDMAfnDTc9PVzthNgEGeppAyv3yYNXuO/jTvzxrF0ouw2fk4FTav8yj
rnNmPw763Do7EaKw8ajdRGSZd4JKAvKrpwRLr2vlAdkh6ZMF4fPHsy7apoCiemvO
+3jyxyJ/E/Sl0lKwwzdEpNDoFh6GgrCp89dau5MWvLDaRRjE8pihYP6bWNPVkyOX
Zjcbfg7IBZnqhKQG2vo6MVBhSL2u6ID2iuIHlEgdcNpDluKiaf0Hshhxmus7wHVV
/FaU2r8EIHq4rB3odJPToRRfUQtHLHrvjDAnLGL5F+nkIwR+08gUaVOpbLzgGfUp
nKcz6uJbJHIZLQeHwPKDQphMkQTE3HtqMf65lbGfpmsnNa+PDddnYqZ28fFtMbb8
D9BcOTYdsIDwwIIM8dk832Yly9XKwjwgEnKuJX7DmpsXEgBFa9mP8cTpUnInksyC
2mNU/huh7lLXb7vsAqcbwJGnpAEDZcy98ZvEKoOsLcyVnWW7K1Wv5VKYrAnSe/Nk
fERkeKu7982j43bYq5gLTNT0v2YPqHbHdTD7kiB/36SYBk8wvPzd8zJJ8ZckNZU6
umO3+4vT4hceysHejhZ09/TdbFb7cph/pClMBpdsKQGTh7qGHVsPVpF6ctaTty/K
f+UhfBAGbyqYt9u3j0AZ67doNJTxs0EFa+pEm73f6GGHz/HiUwu6ye7U4FZocSjc
Gh+5pPRtfFdi7jlNH34SFUwu7WCRtvQM8URaV67klpoBEgu5D7sYkGfEdlTrPN/3
fp4chBlDC29xUMaQ36xtdtQMALT/wZ/UeZC86f6HQdLrWCHwOkJHQYbufrhuHirh
Ijy06hLpy1zMBAp8veOs1ToyYE4T2cWTwpI2TiIeOXsCVYJGE59a3D94TZphHFhh
+o/ACL+p6dlH7mogUkY2suukBxeV14mF3RjiREY3IXTsL60xcAJ63YDEKGBD5GeQ
0Td+MTyX6mOTGbHVoI/EAO24+E4X3R5IXwcWXfSmHO0wTWsD8b72gXYXoOKQdKvh
g9PwEtyButh7H/IFcuAZm/wgsDD6HGjkKtuw+Gel/Vlcgr70UhlMsfoPjS29FxCm
OSc5+a2g7R4rnFS8dGp/M/b5TxsBTY589Qv7Cvd3i/MsHCC7T1vvjRhXoSD5LHhN
Mmty1xka6ZZ4PFw3i5QEI/iSB4coNMme49ytWndQg4i+ubHpLsfc6cpLv9Dp6viZ
OUf95sg2ZhixNeTpAWbkMtdvGoVygEacvAfMvI9Zb4pXFaT983kihluDiR2Cr/cL
Qlf65JQSR+9GWjMlICt6jB7QvD5QKAFXDvQVAgerpmFCd+c9UweqSofIMtoMNY2N
GScg8jJRssAqhUSxqnqRw+ON3MssTuxtt5LHeeJ3aioM43RQGPhxKlo/BBarM7IN
SCceqFc+j5W0PR5JuSZcF/N5vy9W2HJp+LWyqh4DhW77rlPBlhr0MuzfIxTGzqDP
mP3bXMwQz82gZ79uJovmmSsMPHTVE2nlSrwPL9dAgYWW0pDx9uI+G8GGlcqq/qNc
7/Dh1fa47d61tElpLF+ZT9CoynBanu9EDp3oRxuTzGZzkPSdlKD1VxljuorqOqK4
pVLjC1nKAhbIrWiBpydjNyaaQHsYKWVtPW8DB7YKbwKpDF7V9v3j622twmss8fuE
0bHKryL8vtKWZHqkXTet+yoUOYXJ7dzw7CMl3uEolGjDp6Dn419Ew/alntN+SbIZ
SbJP3o/tgaTa7z/yhJk1TQYyRofEXIhMbTnbcr4O2iORCmx2/M/TPnxv6ihjiATP
E8I06FNRHEy3icRqxIvOdqtWR70o1YOrJzhgurv3StZgey5J1AusBcN5LW5Bhc0F
qQRU/dypajECmx+J0eiIZIkER82qAPSDsQ+w9HtFmlov/rCzhv0lTXxKiNFgIcAG
ijB1ROPHmdl0N6O90P4vY5P20WcKyM442fu28o+zNyGy/5g6eZbdOPQek3dy8PaS
Hax773dRahn7NW3FchOn/nfQ7PYZRZIs3wLdYhxHx5XC5SHdqyML/6kezM42v8Qf
7C6VqAmVoBqWZJcTPc4jN5dSfBPRVyWP11b+xajfRitGInLmxcdKLrl8HJvMqMZu
CenspbEWUXVBYIr9sShTF/v/PvDwj9q+LuylP4WysETyOn4K8sXtC8yu4K0ppbZF
zbYn98i5Yi1XSmh/HaS1KwGTbhDOLj3RIUAsPsBVJhJSk+YbayqkvqfpLnGhqaaB
EKJhV5idM28BCK6ilPD/p1HWchbLani9bp2PZEWEhewYGKTUDQkp2pbmNVYA8MiJ
vgZOeyeUF1MwlZ1V1/c8gCQm2BfVbAtvBLSjscfJDGmDiXeI4k39uTTiD6eJ8mYy
VNlReqin2qqxw1mpWE5cMrtj0dr9+uv+3rr+JEyP5GzEnb2jzkStEHqavQyOr31j
X/KgOFJ8JHeVzxhcPt/yJLRBfyQCafq60IhV3um/YrGV9q+slHzmXGAtMtC7DbPj
cbjg0U2rnBRVwKeuPsguOn3f6jTyeGiNdaOvqwNQbBAV5nYf438fxnUJ3s+wMxrJ
EE2Wa3i516rwYjTO0+Kb+bRchgDsH58kYX/m5ip+bLOpif5Hb8WCfS0bGK/AOeCa
skRAHunWKL7l2Xbq/KFj6SubWyc0d3REjcE58MSlRE2F7QoO4Jm1UV4jj3mhxNAc
yzx85SvArRnmVC9yIg3Wa2pGOmGnSnNe6EBnZt1LURzHae0zsP2BsKU9psNX2JPl
EPS9UJg4aXdlIqNHXfRV1Q41kLZar/bEsYQtO0jiGmFfoJiyRYJynSteKahfRnpe
1jMNRMBG2F21O6sIk3hTBkp7d88looeFdsgPOOfTq+1gcDTzJIP0KNmHlsmGt65M
jH3I/NjRNXcFfZ+Bqt27M40s4IjIIV/2r6/NE2d1PRLXsYaVjGW1ZP8j91ZhHvwi
Oz5dVg77j9AWHuxQmusiMqA2zbvP3R/qKB9VmJxS6DsjESc6tVdGxOp9U35u8HOj
Xt3hlEBz8TVU1DM4S2Brkz/Gj+X4WjGKfnQfFlCC/Zu9jq2OIdkQphHoG5HktVCv
gVmMnuysAHfZ7pcGubeOAoMupuAk/+LgbL5oWvwOuozbiaiSN/TecDlLrroKcpFG
1Lb3gVcEQFYNG3IGIQsi1mXLVIlqH1hk/S0XQqAeU/QoRDg+/XtAC7DoSIFYYih6
7GYwN1s5Drq4pz35WTUlll8RYvsUfVBclain9KlHVoVPTzP8i9gK9xd7pAyXfErA
QXPKcWW93obahx1I1AtJW/e2nVUktVpW696XyJwvMYxZlIIVwyUXCuedDx+2YNw4
E/4tiTtaznQW/h0RXvbZ/PNPF0sSu1h3VP52NNnAC08KtKMzM62/qW+MRuWuy1gl
SvqXqAVPl+EwAUD5JlM/WWQvy2LGRCSw5FMvmDshxT7rqT0Tl7/UYYsQD6ypV8Mc
8PzrLVugEdFVWuFdFS/ifPcF0YUm5TMT76rLgLUu05P4csLR+9jnz5KKhyj7HGUc
6NXT5wsh5IgjlFILrgcbLE19BfiuIoFwlc12n51r9ApghFOzzcpJVNifsDGaxuLz
lGFa9R0GmQWGYsleCyki8udgHFjRa6kukAXccIHcKp2iVcjHUUuqFcm3F532gfSF
grwT9ky3LIRKTcAHSbsAMUh1ehls1+DeKdIJbiYNuWm0ZibpHfRJcTJ8O9ONvKPF
H8W+E/9kzUJArLWobiNVxNpTtKPVKaSrnRiN0SSGGy7PTGbV2gdC5xyd51uH6l2S
Te1opjnN4Q/y2f5ll+QB8mu8eI+9xLHA3jpF5cANIcCocWXAiJkjYsccbs+NKJSU
yT4VxqJcRzATHIo8uRKtEAc5Qo5vqtoWjqrBZ0Lj16219/VaOTL2LZGkXnlXgikg
MWXWyS7urxF+NwKbcKRxwSuXxf6I4Qc4T4WifiDPL00QW6qulndZlBDyuG8RpZZE
KRrim3KQ36/GXzAyCrowow02WgSEtCAHI5BfcD8BmPaIbUMRjOqjF0NIDH4QlQHW
cQ7sCc9M6CE0vc388TH5fKc5OOclubri9eeSz3hBfN3/yTL1JmJUIH9ORIqrbl+Q
cvmXVTd17cDqebVgObc3HLsNF4ATfJnnfJ7GQYX5hIEGe9uS4rIJjVMDZch4CuZU
X8HtElsnjOjVepT/N67OEsCchvMCz4TRQXcIKUuIOg1dn7s7aOvWBq9x74mlkDv9
MmKqZLbOysyJimCqMgQZbGenzcLp8+aLEfoicbjPeHgdKVNwL1zQN2WfdJaQjlhu
isRmxWo4ZYxINiS0x9lEpP9WVMBRxO3hCNAHfxe/YuYjXNR+8S8HXBB6kiN+oAO1
IyV9ibsis5cFkiKuCnrE6eeYimULzvPAkoQRGNsw85PTBhjfeh3pJSNeWVcmImTy
iE2ejqH/S3LW/QoHrIF+Cc8/plnRNvf3rfcUARxjqTxvq3ttItbW14hfCRGYfabD
1AtsOKkUnMnQ0MxFrWKuW04R04RULzeA4MPbCHIWbprZTgnhkBuFUKkNKjT27YlU
a9Jp17FFbGgV9GXt7OI8g19zji7Hw/v2BDLB47YXL/oxMGUR76gp6iZ3zOLdk2qW
EIA04c6/3kPOT6+0nCEDf1mnm+kRmdih/4ow3IDetTPMw2cEEAE4FCpX1saX/ewL
lulpQ96oiDshOA+jbJCncinYnqhrAhYz0kQqLH5kjGV0wtYKx4028TUlf/PC9O/P
+e3WVnB5dwKpEk2OVtT5/qKcEjkSEKtdHPIlw926/qPlRqkahHUuJCXCY+u6PI1a
sPiytGimIe6/EnANLJego7xe882Q4N5VbL5G9bfLOONLbdtX5uWGZHIiC7+tPoK2
+LcE65gO0q3shFENZ5kpuWB19XaOhzDpza9Mdv0C8z0hC3qLZ2jwQClLfVl+tPnI
8GFqWR/8ZZEUugs1NHrdMAwCtKGtmZ2krysajwus30FpLFFcLi1ZG3FPg1A0XcOi
cQM5GMlLXowU+BPfTNnBZOrh0cqYnoF9lz0vW47bv3K5/y6VRfFRtZkxEY3ETeoW
M/4iQ+eR6nUKrLrc6DDlmwSCeixaJGETrxzsfMTLKQ6WmItu+1RYskn/6EncTvDk
PHkzghvgCjzEOp26PG7kWifjUT2OOogAhnah1ocoGBqWJ5IpQNkPghcvGMVZou5E
nUh4X4xdB+bDkoQZ3aUhHDDSUc+hyFqqDnFWmZBgxmP81ZcZTQrcYX/nEJHGfYGj
QJG9gsGMp4LcNp3s470oSxZNBWyZAGFNhOCYaiy50xPMB5o2NO9IiHk+yKVMVABT
yLaFI9aNU/LQ07xpGWD6THYUHVkpoh1bsAMNcs2D/lAM3Aad6kUpBbv7wXVVaopr
SbFe8GyZE7AaIn0QEmm1gNekeqVwttYjFnJHfnev36+pB+1hh/a0H8+UU0mqnHel
De8GhwgNOiMEHFeddtTd9rvDplJAOSkMJ3qqP8MqmF69UlVRXfQqpEequ/wLncBy
jXUtMVEx74nSgfdr3fL8X/+3h9ROIj6Se9unMzm7Z0jEUA96cuO6L6YqfafmShHy
OLSD4nHnes+Hc/c8ltYsyryIIopNiTQZnTXZJhrXEppyw5h+XTiIMgMrvDmmmBCK
lzrdFuQ46k0pGgDYoc7ybS2z6k4zH3Bly0tOplzr0eaihbCUzkiCxXN6hrHEaWck
8IxUQ4qN7JjMIKwJFX6i1R65G0yzutC4LLEMb0oCd/Mr4uBwi9k0hBH3NnugfXXn
lyGz9bp9FoTmOjHHOm1QbRPvzgoInG1NcvsPRDyJLsd2UD2DvJTu5uzbtlWNqN5i
+HdgaALL+LfZmnQfkgHgKR2lefXfMlSbKlzOO8A18DHCne8TYwoEbTSUI+9En/xo
P6dJ18gIia2tfRZcLf6b/gLE96JyeOKdYvnKH7IfPP0qX2wGpwu289OmoUYWTm3T
6auVt7sXLaTQpFKm1INuZ6PRFtbFbVOkf0HyHlsLnSjHpRy1I9Wbi52O1+8yJvpE
xsZ2HqatnRa6vM34ej3P38inhjy1dFdWvTRAMyvlMhfJm+weaWHqJh3q6PGhuSuT
2kLX4EDxFyIXbXhunrF3WFF/7IlIfmoqlYWpkIhUni94LBH9UXilwun3Twfu/CTM
0f44/BsBBiOUNVCWIg9dAYODOPFV1i6W9cAo/0mJQwgXZeZ/klXBYL98pWx44Lz3
c2DRJm3SA5bgIiTalIzadUKulyNFEK2BuK1GjaYcGWZfnkQHxrk+99Z2dUklZC9I
ICF0TSvVkrHpATIAab4YjA40uGTDFUlYj80fzZgpAhYb+O40Rhsg5yhpnAg7FN2M
zZBfA1sfCI8an+dkfegQnsRRDC2xGSaCD5fmhoIa8JSE2j18ozh7hCi+Qpt7/wfC
KLPH1iopTPFqJzBFaoj4TsnVrYginOND7FfblgZejenwnLMlHAQY4JwCwfoeA5By
C/fACw7cO9vu8ryaeLreFPOBoIfrVDA3O0UknJHyAKofn5q2wpTblVBr/NYgkDST
8YoIMjeQ+OUPX7gVc8p9xDjMgEAa3M1ewrZsgYPZYa3Dr74qSZov4ywpyVLgnFes
eJ1tSCJ6K2NOouv60eFYToJjIa2TMVpTKNWpHrlnfgBCR9O1RXCt0cce04R6eP2s
vZCktY6qwRZW0SP6aB+IqbZAMHHGFOejM/BlErPm4KIjxbTJ4T/ay3+UVO1qo8UB
VZ94yj9cUQI6BPG4w9HUgQJkdFf72Dzpwr+xId28b54lFSLBXS0GN4N6uIqP8jL8
WPXptWo7nFYa07g4UdDBvB61qjBlPeEvLBSItlHzwEIlmodbX97TRe6G4z5v3G2p
7Xgnd7AhdAi2C6f+0FAxIHq3qXdGRwA72SJwTW65Va6KKPCVnlW+j2SAUWsHJjAH
bUWvJwOgY7NMaAKfS5ku7IQTNmnwJ4FbiYLh4duwG9FZ9/epdVvVLU/YlPx4ORc5
2wQrPCEZJ6T7Dsu509LKjGD6TbOORlgIQcucaPBCfA4Q5Bg5wt11/gD3VivSJqi2
VO6SotFuhg6YJV1+MlZ9d+4bJXBwTLE877zuK5rrCdjd7UV3oQF+2mvwJIPHAkpR
ydzZ3yO9El07q9Pl00Q4k0wAu7nvpHTIV+Cu52KAfCXc9lGtUTO4QMZUxplbaCHi
HOZIQEKw8aCwq/NqOYnFrXzltyykYm4vqKH99wsUb1bN9uvYCdqp4A5wdHiyCnxD
KzcW2xuuTm/hR24vHE/fukK8GEyexSUhsEjoXIsXyOBq1T8i/ny0LmW92IO2fqUR
7hYsuYRbX6NYWffJUxEbfx2Wi9nMXQ4UYMTUmNMU8LXMJ9xB+kU/lQsy2+5fGmcx
8QrX6pmrau7dYOjm44yhZ/KZsxG6hStexewKhh2nneJyCtg3srkqB7ib25Rh9Wb8
1fQ5maoouN4F2MgKghUuXRehIn3HsSV4k10tu8lamT2JFv1YeZOwEb5K1F1rI86e
g3uLz43LbKXWLMQmZNqEgSH7BDZzxTgqTj24iuPOiUB3GkZPqaK+OUaayhkmY81F
PfjSG8azeM6EcZhg81I5CzOx/lT0wgIKpK0HKjRvUUG6QBZ0JDoHEgvYt15KhFSa
iGl5oJjO5Wc/rmxMa7bC12ioziGRoDvBHBs+aI85mQyR1ghkP2e93ibRO+rernqd
R4T1kTLw82/UDDlZ9u2OmHMZr/6au9Q/9sX6Ms+DdKIzGa7/zMp2+2tTzRLKwnci
sjBchkq6AjodR2Y8Ia9oLaft4gKcrOaXDKA/Id6b7W4t962K4PhebW5+KY4QIRKO
8OyBBJZNb/8t8gvcmBuF3iZGWtr0+h6o3oeupqWccSZxmNyIF9whslBDdIJW6oDp
9b2ANxWZmADfthWCUul0a8W4aa9zVOCxeQVAFQafJavmxqkjhiKzhMOhjOumqg+V
Uyb0uGkySJvOdEVI1LWPOIN3nCCzs39IeeVp2HBvtnnMINzDa3HSYxicB3C3bSMv
I6V6OijDW879WztmMNxVG0kbmsHe+Xnog5YG227QiWvsiSu8H5nkRlhPVwAa4wNp
+dnMsaIhY+v2yxaWqbz0BmAXCdMPQq7NnkYK3eAfOh6EPQ8ukBietyR4RDPlmD+J
G23WqXuzAZSAx/j7oFujLr8tcVm1tISAEkJQ26aQ7XFUtp/R7aQ30+FPbizJEEJG
89Tj0AoYjes2l1dzh9LNJgZxlD+AQGxzpXhjlYU0SBhtTjQWV/ObUUPSMKyxGEEu
6lIJ/Ij1ausvVeEQj1MgFbPoZ1vIHb5YdOnA1qzszNneTXQIVAxoKhSCGxBrvXsh
KfBab7LHls4dC7MgI9xWGjVwSA+7pB25caHGlHbzXmnKtY85O8loqd98K6uicZtY
uz7ha1UriX8lyp+zO4pxvs4Fe0cx1nTmXpxrKy+GRDgWHi0RjJ77y7OQoM23RrTd
NXpGc8HuEEkJnhfzXSElf4qPCOISKHoWQ9eYntrxddRueTpNs5ZgvaIniG4zeh4Z
jM9cJe/8E8GjPkARz15ewokEpK2NqMhulAaw6/S0ASa+86Rjwy2gvqfwEZhI13+g
P9LqnT6UJCstfcBRao4ig2dzQqH0S7epgOUbmfs2Pr3RHQmXV75DYfmkZzjLflVF
WZUSzYuLXSsZtkMeHoaFpMHK3ET1ks6AO96ArMnWbHq8R57qkY/MmaXQ43imZ396
cqUqMfEYFFe+c81ID4KqvsgFnnWpanWcTQ+l4EV1sQqiNj7VDvnc+cc3SjKobcC8
El+gk3TjmHJI5Lv901cdlE2O3GySDzLwzQuz/1+CFvWYL1EsK8TtJ6Yrb+PYZetL
kmb/Lh4mU/U4BFgPqAa/UNAk0s42oikrjpzYpdCUJI4+wWwwuelAkcrrcpkyuRcp
eUAXtV/OQOYQu0wJZ8uaBhqFtpBG4uigGDj9dqS3tvBjzx+FNMTbubYlSgSawWMT
lDDQcUxtiNuhvf8eQwOEYyk4ckYNJcaa1Bzk08QsW9nRf2yVOit6W72cbPBCED9E
V6cWDe+NutHaYt+P+pnh+nkDXOxoysHEsQFbQgvesg1xC/T+a+SRT4ejlHDW+32n
BrMNJJEAOeazK5ep0X8F2iUGJEp3Hkz63ufmc8oPc5Vrpbl07mPi7B12Y5OXCD2x
MwZWU4MFjd2r8edyMz3Y1cmTtiUl2mk3YMbyzVySdJVmGaHtfYaumuCwEZ3SbFWY
2WVp4K2ljxDQMHuA7CWriwp0+h29TeINKYApZctwgxmw/+sPkEl6yyXDtmtYk6fv
u6Z2d4voPH8ZWnBuVuX4ZpgoUAqrMuD7PgM3qMnlUUUu0FaiyNUh0jQyo3sSelqZ
Kti1vavzd8bLuP5ERwwuhR7aOJfVQPmoxsAJJtNJdBtpCL1wrWfrIf0AkAVq9yb9
mTicFKMiWjCS6i5fLHNB9ETNcL9maeLytfahNDZoz8wA0g5CSjS9s681Akx0SUtI
tWcVBX+m2x56kmEaxOaj38lruJNM8LrNcqY/v0JGHtItithHVqtiS9RKNDdFsMfm
vF+SKrE8YGlz7+fwTI3q53np9A3cjNp+yZNQQ5AL/2Vr2Bf7NRLhwh9jY9UtuiF0
rqqZWqN9jnF4f9atsNjzOrIFsi+o38+fvuQYcNDZ4LbMhadUzGEyVLwQ+Aaoa0ZE
Ky/Gi3K8FpwhCvyQ2YELZPB+qxhjPaL+O9tZI42CbMKwzQWjgodGVNY9RghOBDMN
sAHuriQ9EcENvwuyA8SxH29JCXK3QmaLlLjRJlCxqM55Lkisiv1Z8JgWRnDcqrQo
CyWySCrg7RF/pXL6LLo7fzn1PiUjh4XEjdARvnnNdqcqzVZ4D4/2E1EoxX9bT/Jh
SDl1cmMhXYM7vFQGqUPcsbUjywrEnaGZFq13gI6XuE7Vig6lAOB7PStX6+U+IrD2
uHjLeu8Nxui/oY8J+8YmOn6rhwk47YdOU0byLOmJby3xwVsdbFKjy7lnMHLOTTVo
xe0WwOWLT0Z5JEaw35Wi2tReC5+99XyI549sGrvrJz4czjwIDv2gXgmmyG1NSnJe
wse9Fx5zeLAiL52bshcG/A2lyk+MgaGCeseoEj3rIh3NhoS1i19ueuw78/9sS8nP
3WurW6j3XH6dclie7QDTy5U2DZLA2ve4D31A6+g4RrVfCsdUZQKIeujAce1Zc3zw
lmmBivqe2+zEgbYM402KsrRtMIiE+HvElXfYuWs+G2AGTbfL5gzTi5/N9ZbFdq/y
yrHbUMFHwqFfTKcTPONLvGdqeJeOKC4Hr7M76q6rAQ5wuTBNkGZDQAccUE45AT/z
taEPGZ0Ipzy+7RX9I/Z0pjIic1jogvjyaLAV8rCr1r4+vxkdkFRsFML4YMmyZbbq
oniBSh2Ped96RzrMdVRWRO1hDfaekxi/U9ORUF65aeC60+tEUjr8vHZMLR4dKJNn
L/w6+7/OZKz3ToEJrLrkGfvCRR3VZf500d+0vJ9K0E732yD4uS+d5N9wEw/DngXr
D2xWk3g9z8e2NWm2DvVugdZnNAnOo5k7H3MB26+ZEw/fz2iy20JgWWnIJ1h3Z9LJ
F73lpHyKPvC7afZsVA+q2cG/4M8rsKls0w3dgT3dZVJSXCmskq7FRrG1amPGJ/6d
PLP4U/LhhmmgB3UsiD08QaO94u7xRPrJSUmZ1SGT27OLOWW6yROPgOslIGhFrlGL
O5Y9bAT4srcXHEfcnjDhcWvLegtAwIL4cY02wO2RZH9/vmAdO1A+IdX3FZ70Jk9P
412glRKT7r0w0XT4g2l/QE6N5g97wM3FS5kb0Sq/A8KcB9+rT28oBBkEL1AXVtWE
SO3gllkGLnMPpk+UfK8imWk0tmhB7gU+GSTvu4z6450J8OvTBNJkMBoYP21SgiTI
QDTfpQBDCGtjwAkPT0VV5JZ7E5Bt+WtS4H5bperKfNMZKkF7DD00IVwHfjfkuRgE
V8CIzbk2GQbNfRqIYLuYPQnjgIj4K7cKWIxBJUpk+C987JFPy0iQhPoOPy1sLecG
Hx29kxr7Ydd0C7F5rmcIVW4avvBwYNJZW9Y8ypPEpS2OjTE2Z04i/5WwIUD4twca
fb7+U4Eb2qIuXkkHR4ys3/PcvwSaC2IcJN5jZGmtCtJKC+ZvGaYX/7S/GoOpP460
tfbgTDm7TckqN4zNqnxwS8V0e1OS+QsZAd2k2eqyMoLwdibw/wG6duJwpsSzTy3F
QoDzNHGi/ogSNPJ3OAuGDGTI1Ma4OlX0peXlfREb1d5vdtrRzfeut10Xic0TRkZW
SCtq9+XQdqZhTScqFUMPVYQkuIyn07S8amHqYl6ZOix3PQ3vGSICFO15PjCtqugq
2J3X0NnR9nNLuUoSUXUP+/1DNaoCm4mSoEEYhUhk3BPsQmmrP1ChUGt6Q7ReeGIQ
Bef6tSWLF4qiAmP8zTy4VdQ5BcZgq/nDAwWaa4E1v6M/iHmQwiLA79XeBp1WT/gi
Fi4lIcegdoOKufYH/TIZdnvIrC/77Du0LJ15Jl3yFSDuj4chPhSnMd6Z4F2w2Ioz
3ue8MPiu5YcL6kvDQ58n/2kY+7x6kx6KPqS4GtVEONXHkllT5+bPbLT0mPuOSRV8
XCev9qpR2B4LpgpC+6qAGfTzes4NXKZXUHFIfJ0HWc8d7W5hT0C8jiapB9Rw+xs4
WLeIEebPHXq2+COQfncBSZMrwdMZdzezyQTNAT2Zk5RZ7JKEyZlBLhnvQzXR0YPk
6BxP/h+sxEt5SHtm7O9gXma6oBBzV5IC63TtzOmEqIAIVciDuRF61xyFdir4dMfR
82BQqeGYl/Q2h2Zn7rjgEFlnJdCnYUctgb9vXdNssPJWzTFBXuthw841FrL/niiy
3q7RQLx/9U6xaCDZ8aSj3LgHsUnj3yUoDXYTXlF0zCnttktV22iLWtnkUPpBv9h1
QA8QM6SEdFfJnwpZYLfnxVqb3pb34JRT8/dx/CoGaecBirLJNI7mQH0xEPzTgSG9
bafFMWFN4raPw7DgDEtACDqu27KMBHcYa1tHa7ic6ivD69Ne5td6I2LtFufh3aQp
d8FUCeLPbBoqsRBZQnfwj2MPnm+shmX5LsHp7IfbfGThS1DXAY3NBI+Y1Mh1qIY5
MmcfYhZPXZmeIt5scMcrc+3ZZsPkYfIGfGaldFdxw+c2XxeZegiETkJzPJ6kK4JV
yFOPl/pJi/igBCkM6ZL0gMZoSCiQVp9rGuCf+2D6wpxzrAyYSdlC3gn0JxIAE4TT
UCekAZMrGxMEv3/xb5UEy1/YyNQz+QjjMEsCbR+y4wxnpsWdeg4o+FMa8189owts
hGlpnRU9sRe4mYz7sOIjAmuUyCQ0/RZ0jjMvRPLr243lsQ15O/DUYkZhKEq9MsoM
LB2GLwpoDbYet68L3jB3qJH5NGI07DmKyxYtfK5viSzgCO5bWKqlOI2AXg0Rx5eS
M9/BkR8FoE5DJnYiJpb+SGijkafdBamgLN8HJMHrrzy+n2Py1gubYyJ1hto9Ybyo
pf764XBaZoGyxYGY+xiQ8W1m12VbMKeS/ynrDX0qempKUybPMYw1xCbb9oTcADO0
tVIhyUuqZ++R80G/RCX96oKulMgCwXhy87+pW+GXeH+rV+0sIY2IYrezZ2xUm08I
dTu5Vyw63qKWnOCca8AlwJxu/AngoeZnDu9k5IG3wRj++KmPLHHExNQ0BAlORNQV
SiIaR5HAgJvWIyLZmaVBPXJc1D3+TX5ZohOZuUM0o7ph31StpG+2kbognu6VRnv9
+PBtHpI4txemV1rkw0EaejufhXc7DnM7veLUXm5/+cTLaObHBsxaW6TaPNGyNuhi
6l1LVmJ10Xvq5zObwWLI4nzYNGcYpZvHuhIDBe6AId1vV3/DjrMtvgFuBqgCJEOc
sR4CgvDAynUpeHtU4awSD4F7R2PGXs2JT1+79/uvAoWIq8gF3yDQtH/7JdRk1jlk
umWNdtz4rcjL1txXheYmY4MoP6UyQaQ3k19XfbJoUK3UNmyi4FLVh5UEuV/hOg2F
P02cgJDGHAd/xdd0nmduX2L74qrm6KLCFOEmWqWyphnn2sk4DYrYMJNNhLfnicb/
LyywdGocus8G7Dz76bGglDzv4Fly/tDhISbI5srmuBL3L3ps5rKKD9t7eTPajf/P
jJq6cnU4IUPTJmTWezLzepb0LKfMyUY7u135tebscl09h2kf0TukmzhYq+dde+zk
tjHt5NgA5hqVsHBMKYmqM77jvsVNdH27BXV8N4avFyWAlMkSRtpdbUFHiwtGTCjk
AdsQFcgUybmTd3A2sXqtSWuuTQis5I8medha3R556lMzSN8biV4fcmv/p4ZcLx8v
6l0NiorosR4kZVoKXUeh4UssJO6NYCT8KvV3GympvmDtpNm16FVSut2rgyoTvn1u
ysmFri8B8FK5pdi4x71jgP5IN0B9gGE8VLDyc2N9Xu85gk07pDjibqYkByR9DFqc
JbbJ8W9Op7fQfvPK43ZC+qqpAayWp4AmBMlTVPydiNzknjvg1bA9qoDMJ/BisknE
HkdZihooLqsHOAD5WeRoU9m7BWrX9gZmE7Tf3cXcxmPhbUfUFtDuPzjANpGHZsBh
7Y8N3Ag8eamcvCUIuNXxICbDsa6FabRwysdWaNrrUp3vDBDoOexntZhfRlt1ry5d
s5SuaQjJSlVqZBilQCSbw/Ui458itvyH9dRG6tn77f/W3DinLV4jWNv3kqjjFtFa
mB48pyMyJp0jAT+NAqi8Vm2+EfOXh8kf8v1nKFVTjwVOM7/GSTsP2UOCOYcKnwzP
8Uigjyx027w4i2XO6X4bVu35XG5jy0qHBPpitfHe/v3850cjDcrTBeE7GZk/jKHO
sxf6KuYi6flhFxFQy8Do1n56KadUC21TuwJUt6XMquVNG1ZB0kNvMV/7aX8Ja7zM
yQeZgluengOY3C8EXnwfJkLK2kD5BtgMJDhdLePBQzj4P0eFbeU+ePQ0fsSCRkN9
zcqJKwTZLK1jbjF/YwI0R7/WS7j+jgBDRPjirHAO3PZhOWXgsUga/hLguKRja1S7
U/7oJeKNNuj8bhqGfExPe1wn+0gINw3LGe14dEvlLbuK2R6F6gQzRVICBaYWvLSe
sqsFiFyqvtqYcEEFkbyXnUR8hoS9JKKvxHubd1mHIcQ3a0eX9/SWhjxUZFTHjPzd
9KslDJUG6hYTBcRtpKGbDF68F7dxA2M7DXI7x0fPQkbpwPv7V24gnpDF0SiRvdD/
jQjPo89nAGNAnndoCRIMVzqcVHRg1v5mj9qq+18NM0RNIkTVi7y53CpnFJOqnzLH
6Ikk7qFgxForsHO1gooOW8czRCoK1Yi9/17if0RvGXQOL5i2ZYhoVDUvyR3Mua/J
AK1kO2V9/4TfCKk8xVKNUDUa9Wf3aKtPh7wybmRf4cPwjjjperIeHOvuYkgKHqez
Sv7VKgBkwCbHdNNFH7ysUuCv5S9JE/yJfpezmd75T7+Ax4aqWUrRbi7WFZh9ZYMb
dcZPbup0HiCMZ7Duc1sFs0qCANOA9gd5lV+Sryg4/bcS71PVZx3WsHGAS76smTl9
PfedW+36qwJ1Bqk/EmYRIIPhgVUCRi1ZK/6gbnk2WZmUnULrLZy9ObWSMNpcK9AJ
Tsr33+XExnP+JIRCSh02PL069i+YSmCFf19j4kNTqUrz4RaofFnjRmJ5D3jfpmLn
2k9+FO1JWOo4nPyxh9o9ozvdpz3z69tNEeI5ae7ImnsVVplPLgPgq3Omm7OM1sUi
DvbvLIAuNhQI9u4yZGunLgX/P1AysWp8uXNE+K7jTQIQxtQsLZA3btiyJar/AkvN
QGh2+syBEi/98cfK43cRPrNiNcJe5nmllHN1qJB3pmuIj3fX7RHL+LgwB+BAuraD
MoQfLuLpR085GzIA44IeMtjzTz96P+5yldiN6f2Jvlh+8NUKggUgIPHQojeR06QN
dcyQ6Pb8LSeWXdj50yX6BFy97EFZFyO4tK9SFFkToaCnmjyXyGmddqzwG4Pr1DML
+xtQjmgEv5uc1/ENL0VrNzpuneb0H7A4lU2Y7DIJSQL59qTFvixUR+dYuqopWjDZ
Of+UCJvyMj59FPr/VOLTnNWUqcwYATpPCKHFG4hw74HRQzSDJv8jts0PSLapI1J6
/rJJ6xMUPzmpTDRi1M5ABR+jANrgcb2T+43V4hmuh1ASajXsUGbmgpjHmq9Jfw1B
cRPDK7ELp/P+AtMJvq/FGaojU3wEOk1EuKoVGljC+hVSQAFODw+VN9HavmDyVWNh
X5iPDrVt9lfeb56ZOHsnWnyMOANqWHhUgCWOwe0hywARS7plD23evOSazm4nBdLW
ApmhCRJtVb31aDPJrG/zS0MwkXPoIaeBS6crUE75LH9jvdgZTcgVsZwRp1PGFkqa
1rTbc/pNPNypaxwi88B2IaUzTPf/w8L6kugpnnP1gkVaAroN91C/xJ4OPPQMNWtH
7niJwDrwJNqUyLUqlarbgK7RW/TtmDvk3DUn0wqUIEEuHsDC7hzsZSTJSSO4YpGz
Zbct9VXttKhPvlnlfkwk/zV9SFX30UeY/vrF3WKue6Jcsx0YfYg5txFNdLy/6teU
yuGoPEu8W+iHFZsSJtS2fEVZfjKczV8kiyvjJPZITS1dNCbxApP3Y2mm3tsEr47a
d8GkTHTKk8buUcMT1KrR6ZUwTC1xA6MYX9XA3x+7g7Tg+Hf33jocak90Tbj7cwWP
MxD/kd8c7dk/FzWV+wkZXREwvySAZmvHp9pf3R76W+tI8DJk56wb3xEakv4pS6Gq
v38m5ge5bu1iWFnA+ER09EdsVB4pFW29w8/sZ2YR1UMOu1zR1ZdFUNAxgNCsQVDQ
2/jQ2goecDAEFWHu7uyt9v8+/QbV7hFRGs1JBTRy+t+ny2qPEDo6xpt3TKJlIxoZ
y7KYX7VOF1bmjgHMKfeE2v/v5sjGuBihd0pMkZTp2hAl3DZJQP5cdXvzcokHvWF8
ITPjU1kHWWaOBlTdxeRGYqr/b699JL6CmSrKAQtJZ53U6K268SOU2bMkdRreH2rL
3lROIxNp/MuU5t4mr0ttxOJWwQyfS3yKIALwaasBPTLLw3gK0E0zD6rvjTNxddm3
jLnSbOfd3I1YXj8Xk1rOcMYOt7sgb5rnewuTSLPDXgqrdHDPNYHzLJaqDWqz/pUj
t6csodU/EfUE5KpnZdhAwiDgezWIT8+pyfPhC8VIYVt2a5k7vtYx5bGGKdNdrciK
G9DMSv9QIclgU6KnPV/XxP9iUWlk7owDrt0iN/4472qDnVxHkvNaPT/h5sqHhAbr
XGVwiVCNxYdfGHRKkC3Nt+CSJk4QJlANDzNtYWOJBcbT+UbQOo/JIuJ7nN1e3/l2
XeulSBogLqRAcqQikW7TwZqKy3nTuJHeXwXMlHRtw/H2WHroarpp5/nbbijKNpBU
N+pueLl16TdnAyh4j21GbBjEU4nVsiCP6Q7kCnt4+GR/34jhjTroyWDw/rHQpq20
AEW5zCaKoBp7U4OoFHABcbQ5a9Ue0ITB/cAVz04YVYCTlw7pJdcWOQsrYDarfoP/
ZVnIwWBxZAZE30X64XeGVqUUQlOJIJn+gTP6neiH+7weiWXjb8t79CjQRQ0x3XCU
4hqAU2ekS99NJNSp+q0EgHCbpj7KqtV1f/qcwyxPP9Fza3/GH4RKPyRiuV1PxZ/2
CLf9ceHkSqldYuENUZDPq0ahHzKew1ieiuKUhKC4P4J0aTs40txViw13aJzyJ+X8
pyHA+SatDeRFrCt1u2NKzbFFM+VrQfkuElH86ENe8OmMsnG7+bIeRsCqQ23BStR0
R3lzlG+x28U7g6hDx0qdSiBCEbMIIoQ/qfVaV+DzKH+NQJUmKDRyWXcVlxdDZgFT
cbAkZDaK82timuuE7tGrH0sjJef00NDT7oD/AjoRmi1QNzRevULhhZT8jrAsbM8m
Oce5IVY8Eqf+Y1b7PYhRlYf9vgqP3bkgcNkZIr1AyndpZNDJ8KesnkMe2PgsxTRy
sTJKtE0WqaBa49lTqfzKIFg7E8WK68CIGPenqlCKTywxlk0MaHFIQ1ylw+GxLcqS
FGuasYNH7RooaRMSYuiqrQoS7g6544ejkgRVMZ23cBniJkxiqGuAxFXv9RLkWCnQ
kUtM5eMFIBKZnabuwj2QIXWgJ/h6Fl1DHWVpM37sdj0tFT/8p8fFseMkuIb8h4Li
SOlGUlMSUp/oLFNL4Dsrf2FLrSI1qVold5GZmC7zlrKsqoRQj64rveuKOhTCBB6f
e7cmMU8l7X9IfSRvKnOd5r/zdFFY7nXgGdCxj1uSQHOt1pJ8jcb4FJr3+WzndUvx
fAi754g2Rpmc8VYL2AYif66BlQ2vUfvDCC/Q65NareT+UG5x70bLIvsVM70ZzfA7
VukigWOy90KZSlPbkL90yGesvAwGOzMjWc6KzF6050E1ZNAaDEbwVSA85g2e6jDR
ba54r+Gb976cY37ymYKckHZ6XBF8bcbVhzLl4FEANllp4+WftDJ6mNcRJAciwmTe
uaj6kr5O73dVnyPldmPJpwcUbsEroMLnZ6RgLAi7lZlxODMsbzfk9ZTBjGkmLQJV
GiySGrPuvcRCgGfCDonrAOWDtqdUdbQGJQnXxIQUURLbb4YOoDrL+R4P9W1AvnQ1
FM0FEnO8bLuDkzMpZ1AjJ7YoL8uPN91vBItzeczTm8VRD9hwcW3lFOCes3gLrN/d
5XAw1OJI6IppWJAT/cMXCDnvlL4GdVd+CD8r21gYlGYf0clRTne+glMCLorgvfNF
JUGc2CnsztTXhJddg2XCCBK2Rm4kbaYDqhi7xgTt+8wXJnkMxVHirWNz7EfFOp5O
IZtWmVbZynYvw4j7Moim9koV5ZG8fS7zP/SGBvPXCTdxtc0ygM+hDGXOBEHCKV9u
FO6IVH3SkM811tGpmULffpTS/EMhF/kNiFuf1Lyda10WIdPiOnC6lxvUJb6I4y8z
xPW5vsCIKtlOiG9Rrb36Gdhn4ROfbm3GBtiq3wmo6eaM0D4CvR3+JUA2Uq3feGnI
LpYspM71Ujh/XR4VYmM9IfuJpoeiIZ0ZpI146kOh11JRAQAsmgW2BxKO/57VZ1DB
vlI1edi3zRzQbs1sdHeu8sFk5pwM/Epg9JyKszVmROJeMG0UvfSLLhhOkLmWZEFR
dgFkagiVwPgnjxhEAtwzn3iIhviB3d0esiD31n9p+bizF7/xAABxrkaYLOKhYarr
IAdblP18NXdy0qD5rIyMuia/Ho8cfOuyhqx13UfMzSNP0moJ8T04sLd1iI82qNbI
V8OY55BD3XMkhbi+UpkaGY3WVWLmIvaCfig272mVVLrCm++1n34Q2GO4roOoQ/ns
h3onFe9LKF+OIDXTzqWD+OF9gBq7NgggipLoTCN2hOsy/24YMaB1kVFc6G2WlSQf
PLGARXiNSLkMrnka2CbbiA+RRg+ABv+0ELxVIVIl2Gcv/5uGAiuECbBXtNckJAqn
PqbfJChM3PmIttpmE4GhJxrd7Dbs5LsSNp9Vqez9zgWjOXLp9onD9BlQDp/AOdAd
zApJy7HzgEf0ZkISwrbVLxjLFrIvcDqVSMl424rXgyA+ylbMqBlTjx4Srs2zPQ39
jsgY7lBUW+3nuN+DN/pBQuTwCpDmBidAQH7Ek72nBSubnmnRjKtZGuQmvbXjqiCY
XwHQ8KTwBRVDuUPWH53GC195nTeduauoF1U6vTKScFOl2co7Hdf3jLhqzEGntDOV
SiQSlZ3AFEOZGAOM7ktKbH4LcxppAvJE8UnREegLb1criJUd+2Ws3hHhFmpbcKKv
dvb5cxIOreCAfNBj1QKDIc6dlfSOICHyH6bP3Sx6js4gnBautF9Op8egBJ5odWB5
yzQ+GT5iTdOP3Q5rp++SLOdLjHJBjFobmIrA0WXlf+sqEaWbAnyPQw7gnk20SOp2
c7FFySTr4OPY4Mo1i7TZnSgnvITvCsO8K66XRwJTz+IzJlqkXJht5cpFyGcrosU/
6/bHvP9h1k2peDZDFXlRd31ALVpGcg+Ab1r1ent+JdrOYRpDtzQ6aKoogrjvX5F2
f+Dd3jrJFPGGjAeg/6oUHTmnCohHsy4BKEqkk9VB4jUSyZ6v5qDz6Szuf/PlFxN4
AdwUqZYxAuoJbciVdWRmqSbgBCrkCqOu9apKUutGYEGKaRWO8NvIzj5XqjYQ3QaE
NOsjXKIj8aI0K4MBE4oH/16yuW2yN51FlTdoj3DYi3RUSYJo69Of6s0rn54tqCwR
dQaULc18hOz3liFlZ+RgL4MNb/Rpp+HlzNeictp6T6volG2kwbXxJ9MHsMlneHIH
U+0FxYfh2BPDltnh6WfnKu8asGFwFxC7GbuFPFz1sya5g/QSvYvNS3wRghjo0Ake
aRTVyh6bs5rp5dMxjklsihqY0KiEbLYUggy9+KPYaGn3cCQbQVdXrVDPNrYllCDQ
TQ4OW2DIx0c5SKDMuSMA9krWdxIdli2/oFK/fzNXp6eWpHEUWDsUPnDa1iddkXx5
DwUcdhNGLs7O7EuQhPVO2ez90SG+2QReHS19usl3106sSGZumlm8nhZYrbTIkvdt
6UTiBnDoWnLgCRTc9VOySxtuU50Gq6k46tPuYwTdn+KvBgv1lnFLfc1vwsPADbnm
Pkl/6YrBAAqTDRwQYQoCM2poATITMyQLl5fF1JY0BYjuPx/8ybB+2YWoUF8GdYd6
2JvNXXzvqvThJcAnRuxGaThtZ3WZcojPc/DepscORKuVajqrvjhL+Ep9RCV65pzc
4wklgWdZvz6k3wpEIBzkTLvmjtldnU2kbTm1ja8x2ABFdBEz9yv+AvUbvPN8cjh2
8C2QCVD/PFGVKuHdNo1PbuaEIfIp8Ysj7OrPhzd+o/KXYlFlGX00QdqWJ2fM3C6X
iWn1HrhCISInYCnR99m2xiJtZAVfDUw9Sc+G8tM9oNJREwl3/8E9NcSwxSa8kkV3
m4NoeB0eKv9gRGIRmNqoTJb+B9+FUhk+iTsMsti/SI6ox3sSKyjvKbwq+ZSDJ1oJ
OcpOF41E+lq15KfZcSjE3lObnsT39uj6ap8DDO8rAaJjS2xPEtWppEDLHFo/t99Q
Nr1LVQx+AYFc/IlA2qqBo4gWN2AnFsaOq+kS2RvVcXVX5Qu+OcQSszDnmawYkvBy
3mwuRmnl7lrzkF3o+nv/fh+fFqmto5fdPScQZBJlG4qej5dKq4IEcnUpqcBlFe8s
5paEkTNRT8wU1bTw+Pxk2+u+BuqM1yifkmBIBaeyv72bGeaonr5Pogw2eAbPjTeQ
ZWw3ryRz1meVDkXIa85XAJx17CHYtsaqRRvRCx6UJGzmSMBHx0oq7/PnajGc/6Md
GsUZqvYWJj2KXuB36i7C+OQOE2sZxGSvBD2vrNQxdKkDd+Nzegrb9zhtphkQh81/
WycA8LlX9N7wJGA5kQf75HXBGklFJ0QVe5HA79sYdKciQMToZGEOb9B3eXCe4wOy
7eAyBKiiiWCnkKd6KGC5CEyn6g7DsDFjmgij/7zziIqaEbweus8ZtyGfCgXzdWkM
rNLMBzrWitTjWgW7V6NEB/Xm53C5c27Y0OlcdeDOT6ePiQI6HWw8viO69TOXvNWG
HUEEygtaUe6FX0YK4jg0vCeTgJFQOG3qyOdkOU/hxpxiwvrvo5pqUrCxneUrfLsp
RsqllpH3M6KP4t+yHxXH1F3vwonxR0GWV3YQwFhMBb52sj2B6OXtDgyISRKg3Z8f
ULIjHTmD8W2XMhs+JvraiMlAyE09hjMmAvppb9uRUs0YBobzzrH6jMSGeB48iRqB
jZGhpWTHV44ScZ0ugrhVrG+0U1DvQv1vovpYlTJFpbnIgP9cpiZ8PcsksnYLnORn
TYZ1RZLpA2adBX6RtUiRrlvmOsk3xvEBu9D6eJCEaj35X4D5AxF60dJVj3bzMjWk
lhBikexiVYMbL/iraZdy0hksrjIKPoEKT5iYHxuMC7PlnjyMDTKWTF/FodS+93rP
lUftt11m9qiR74PTfxNJPDPDBKWHosEkKchP8QE2zdtfw55vnkyx/u/0OauAuZ2o
Za1X+54qxf3X89U5JQgNJAvcm8VxsfGYHfN/aDYpvng2z1iq4z7mCgr+FG2WHgJR
Zq15/oQhG32fByaJUp/gTy9TY6RJUDK55/NDREkPTqr38+YjYv/u8O6MEDtESqPp
Z2YAc9T/BRISgoYCtnxr0xj0ujFTBvtIs2oXYmrQT3L1uHCzNwcmEDN7o6ksYhzg
IGRR8Z8eu98rNOuWpuo+ySRYycloO42Mf0Gnx8wP4nN3dOCayKYlnRW/ftSj9/qN
Muh5ublPpbw42sCsR7JWyFzpWpGYZtdV/8YE2QxcXi5AvnZuIVeb7MpMXjQ78Z9c
19YUFDN8My5Ufrw1fyAFyGWgFMdcN4JPG3ugvrzEgCYWeds9lYUUg77efMt3clBK
Ve9WOtCytI7M1yGvJFKrujdt4pWnUTq2WA5sxU1zTBNgM7MPS38GHF6JBirqutjn
wsk/m/v1fUyAziTcw7nPy1rVLXudUoCpu5HYXqILU8zQmsKeltN5j1E17qSji9gF
4OrvJk4RCAfhVFdcJtIfPSIXTwN+23GOyalxKh3MJ2zVqAkSolx1hyPpjETI9jc1
GX+cxAzo0EEaO4P7Bztt+aXUUI8lsotM9moydllYwyczkb1vH/S2Sj1xWJhm69vH
NUgmEh+/QjfYK8wRC6zhTxnTAV+NSnNOlhPW3lNhRNwl7CO/lRFWWoN1tax2BrGk
5enQ2Zrd7BPI4JOacLWKDms2IJP0mdrXHljCqVcB23VpFd7j/6kBSvxczbdNTazX
09yFx+Qo1jXYEJ4ZIAOWS6Y2JxDf33K1DtqIdmgnKKfBoBgayWnNErDdjIAu45jz
s1hA4gBlSe6WfUMnVcQVkNRTAogg91Ll71CqlL/8+/fHzjwsn0kKeEd0N8yVf3ww
BGQwra9QCrq8P4IkuEiUPcvZJ9PK2TMXlWHIiRHCgaDDWvHUAZ0wTi6SW+tZ+NBF
08bXefdNusXXix6Wcqu8htob0I7XJPzGSHOiwrrdvYnxtkGsUGn1wWsd20xcUylO
P3iiz7Kosdf+BwdeWS6IC6Qx8W6QThvnOQXtL0qR9xqVMWO1FOAksAp7a4ZkioxJ
f/8Zp/56lLgz7WY54rYfGtCVdlQT7j67oAx/rfgfapVdpRTvQjolrcrptex5GAZ+
84yqIBTONl5FI/VBHYAjtSf9NoxTQRvA8zJUul2wtj9W0bb6ZQwFRVrDsaVmZGWw
qT16UGUUFbwG3rMVc8YgAaKGkW9evgKmmIz+bKOYMrmX/y8ouiT1zv7nlHh2WL4p
ubLBskiQx4iosBh+O/i894pbEUhS4XEsGEVkoOfrvRhknLVv7G7ukV9joVFmhOuu
4qdomVRYOue71OKYOWH4fYQkeuYlVc0Bf6Wg0n1w2K9hYZVlMG2FWh6Xgn2gGTez
hxi3nb0vpLny1cmoejbhmj6IJjs4gsRwl2k9ZPXl7dGNwKuT5zO2Elx5qqnNqsiS
NeWyQ1lAikijZ0LyIXQPWh5dZx9Eime3cmv6cOBG9+xczITxpp9MYCu0nLTxYSyC
Z0GfcugEnyWL4JECgBGijPyIlX72ugSoG2cNhePXaqOT7gyhSu/J7v5m0DogdlYz
hKXo1icdVsIAS5wl1gaAbmGWu46Pyc2OVLzF9UpElxI+fmhZqVzqGo+s9TFZMYga
TxOdNeA8UH+iVD1MnoT/QUaaznRMznJWyY44hpAgefiINcWdCZHrJVzm0xZZWugp
zVb7psfhX+ENmLfjDUWIqgSS+Tq6r2cwQkc/jTfzRElN/BMng6aW1VWccaPRS+4Z
9zyyu6av0VU5EJ1sRS/L3cm5vMOAYICzNVxt2V0Mn9sY+j+sPDHLzwf/Am/osVMr
3gGDrpjl5Ca3KFpTJw7/llDm664/IRSbiTwwWG0b0rU1WL1UmDT26cUjX5+n18km
NLkDlQcGlJXANjFto4n5GtiEQT7dTrmFfbqQfCvmjeVVupmtdKu15tI6SwgkC2HO
H4Nesg8gtyN0jq+F8rkKmfD2CwFrHpldk4F7q92qxkbGDkhFsvLXs0rVO9GAodxt
mfJ+XF5vFR/mgj3Bg99MBJUXOIOJwHT9OSvzWiVWBc3XqSO67bHpxrgnPd+coLLl
yvJQI8qrRz/mKWKmQBGsgBBG6y6HLsSt5wW5GLjgMcxCxngRFVEgIuC7HyZO0qVh
pE5YF8eua4JCp1ifJfU5Na71mBISY+//Zeupf9UTQQLIB9lTLM8PHTQFTMYmjjAV
TGzYHwdpZLvq6KXMRQAMIPMGfO4tQqHMUZ3DNF2kLiZ7ip5lDXXxgFigR4pN6OIT
QBm45gFdfI0t5W1Ys963uKRK7ie+u7RtAUM0vuE2OGhJK4ZU83THfNW5v0PImQnb
cu4TiMHV8ajFpRKmrOOAXg8TzsAy3izyvFsUwKAfUHR23ZOLjOJf+BL6qNnvOu9I
M9VUVOha3rkyYEn4VQUJQxOtg8lIRTsiry/pRlu67uO4cmjpBiSKxqBC5e8nY9xf
eMbhnizH/qPieKrA1SJEVMw1Y/2IPm6mgdoTod36UhfZPNTW/A/P4CmifdgPJ+0i
j/M3BVhdId/jLJciE050WYI2S4CYiS0qgNRPXOz81cnvZfDcU7L96GDK93qawVRV
Y5Du/eT+yZy8ZWEtuVkI9bFJOYEsxYlFxarZMyO9NqDlNLykAe47/rhJCjZtxemU
hiTugFKac+7LJdFsvM3GGJOf2StOcNuYRLGMjJV2//iz+VqPZBnFWSlK3hn1BUbi
iBeUedXNUiGJF+URF9STIPCl102xRsfOvQQaWnT2CGPWHD+EcjVnWHLHW8PS0xro
2KlI4yA8161pslKGtHU9J0aT8XNCr/+ItRkQh5s7m2q96tumint7NOk0xm3dLOZs
7M2j5H3EDFpQ+7GaTEj4Ck59ClieHCW3emY3LzQHZsXJ1HC7hOy2ojteTzBaTq7p
yjVdAnmG0+XkZOFBc2AJx5XP5WJWxVA2XaE59HWfoOnrRjvTPRKdL5cruobWe20t
0ukPeaex+TcWUh+8AwAut2PhG8FzvyldjCR9HH84C669cwiOdd9CqZ+NI1ezm/y6
pSwroLg7eia3hc0UbR+/VYCs3RuxaSSxGrf+OpwhS3VUv5FhAhlTullk8cCZibZL
gdpzdOlNQVPPJcqyxs+V489ZPT8aCEQGtmT338IO45+EeHmq2zd0loUtef+9TUJV
ZJ6qtUEV74cEm7tO2V2IqICDLi0VeoTEm90Iy31E1wNbhn1hHeQzYmPuNHsUAPm1
Z8GQwaf+m9Vn6NhHUdmk2ayDPFJF90UY/KE22JvBco182xWcxL7WMC9aiR1As46z
FvUiFuqdW6TbEIF4sD+3FI2igOAAKkGrzeEZFV49NiC36HT6v+eT4+5KeEklnKOY
z7xy6WK3VMwtCQoDVQs9Wz1OUUILJXdChJ47aoGuJnEFVY3RqpWbEMtdLYcVsgvd
QozNQo/wiFjO218jhWM45orOi+ATXkP+KERI+vnXo+Wl1Y1FxZGO1ibcjGwf6UAF
61oERlL0hevaoWpujcoBxpKOPct4HOh4oReJY3aAnOCrVznpxdPcF8D2f0dCXqQp
AW+XpdLQKSW6piLOGK7RBjlx2HAVwwWsMVvPjDFTO/TZdt/JwJ+nozTBYQpzfv7k
8Vb/Z3W0dPMCESU3gEoAWYQuDPaxpLmDr7TdsD+i6Zd6drDrxmXMue84YMym+WjK
0P1BycRWfYy92WImAogf4Pf+lNgtf39cVfWBvE8KJ50M2Fc7fEK54aPajaz5shj6
ViYIbxS3dIXTomG0RnfMb0JVSnwWCLi3p7CQNw5tL5YJdNGRBWB9NkLlFARXiLdh
5UWHWReFddYgpk4ERtPao7r11qHtcLteoEPe49vxj9RdWjpWrIaoVL2bi2YOuhCT
84dZRnJIYqBMsgAfq1c14M+kp9kgLQwLm+CCQNhKbxXe3Af5t59CG6xcKDmJE8QL
p4ClXpgelC0B2uHq4Zl3ROmjaIA9leE531ka4X5fM+FYgPJxtxhTrraJzVH02Lit
ASkRr8pcyKg3rYG1P0L67WvcqNmYZGD9ElUVueI86NkA4sifqj205qn81EJ8r9zs
tedcFUN2mv5DksEgJPpIVpAbeD3x8nYmqqBJjiHPyFwxWvlE61Hc76F9xfO+RokC
UZ0PGH0RoGLFP5KQOJgGmgKfBKj1NF7hi+HM2dKgqACvKNalrL3AGD0MyeU8DCo4
G1aUDpvgJ+mLKI1rFgUcJFge184Rw1nZIUEiAChtexPKZ/zTHWelpP9voJ+aTkfH
ISaMoDHbWv1RzXuZiuQOUYLc35qGExNrtujB39YhhFN3l9e5r9nmAYq63wXWlsyD
ANYjuoCxWQnHR2okqC8cQughQk8IYCBN3Y46WOaC/670Ck6a83wfVfYU1uergZml
j9UYjwuQR6C1/L+0NfMkeVRgBoTcvRMMw0G2Y5DjlqCu6nLiGnthFlg4tvpgyBLU
e+DSDaWimXU/sE9RMbvl/QeE4lacVJY60w+3bdCH7rZPvrZkddBDCBGU1CR1Q1VR
VfjiWDTaku32TeVSadW5jo69tTcr8TzrEA0NPc+TsfJByVmg6QUWBI9qzbVBzagV
SthI37z/8qUyjTL7KJmyxKnCte17+9RzyXRHUGgN9B2uYMQIqZEhqz1tvInSekn6
Sj2s76wGYsl4lUinIgldLBdsFmtNryodTBVsuGMxtGR4oM26m1xheGYtbdOGaTcT
oS1uLktbG01sLmNbgU+RPrY1YC/ymMCX7AQP/Lm/htj9cNWIG83W+SxH3NgDHoSM
G5CENlMEMBCuG+s0K8Sl5neMAVcifqv4IlrHlcmlVAH0OIQk1R+QCB28l62K3O77
4ccMs/lLoZnbBTNEaOe/JW6W+eHfvVNv5xS/pCQuao19DQ3D+xQtHMqZvKsRk1g/
NLgMDEqiMjQM3g95GoxmxEGs1CWikdemgtgt3Uh5WmvPaZELQcF2iK/QKg+p8JwU
iCFxuJ5nXZSliDYrYK4QGth9KJCkJnhZZGzM7oAxMBaKZQ9f5FornQ8KYMZDgdk9
jv2/XADJtqgAjTuWpsGoqIXEd2ON0gh3sZpd5zXJv9GgclHwo/ytpHFEOEOOhnQN
RXcg8xwJTex0ydnmYfxLgvOkI+LoI4JX9wU/SxHCK+IMPI9STIluC86I3GxPWg7P
QwzaSU05P5NFtAuk6W2QVFw7GExjNeICX0L7186CrT83xIo9Yw7uwq6YmqXCu76e
E501ugd/tVZ9Vls+J6WbU3wj6sFxrKId7ovsoXWJJHq5h58hmHAZ8AQ3UWSgH3hX
nEasVw+aGt2ouBfhf3+7GyySL37/2B9eFSOoV8etyzkkS8vUWljieWHDmvqAHZCj
ZFAOfUF12FTiuIcTsGm1xQ1eYvWIU/vmlTLJqr931eSeCv5D9q2efgE2TFZHu8gh
/wqwPcU8MYf8HBlEhxsJFT7E4rEWtWEnbWCW1q7HHjlH+bxcH9s9caAC3v/ucuEA
CAR7cI14LGvZMwkwYEIGphbkwAIB0JT31zVlu45QIAeJKRKjsBV7vEdOJcyDXi0g
PaHtvaUJvvbrsfZzq6NfFqRZ65Ku0tzOjY4tL51C5BTvfRtUbkZvE8sPy8IpbSgn
B7IbEnYxKl/5FRKmXUD1vLabVorAzbFz1Ed8eKkB5yorR0Xh8I2ADvdSaBLYGuFw
UM+kQc64DSxl9WMZsa+GwwexkAoWzRtmltb2g6HrLxeYWiaQZxhF7lgyrGVAQRKn
tPKpp0Wlw+gcQ5xpCax03jUVU+2mOA2E3QYGLuGBr6gWS6RzcDEE/U97pOqWax/F
/307e4P9Nltl5QsN3kDlvaArqRUmXzYR3KEWIBjAoDMy6wLF8nbN1pO2EuNQY33C
oix85Le3J00MbnwP/nZOC+rG0ROM8QT5Dl0GY06ijhP4YN2YIx/Ote865OK+fMns
nPYep8/Oiy6RZTHJ5sJwRsK//KzWV2J4OJctN+xDrE7O534VneNX7mt09S6qmPd+
zo7GVmmI4bJJgOQqAxCLywPvvUlg2+V3vbvk6mMLOd8B2pNrcm4q6TRITgLbZ+OH
08ySNKB0MNcELfiY/RtoOoo6eJ8zxGOy7bTpP3hFDWspcj4y7/1BpvtSNLP/ELxn
u2z451juThiak8sMoujChCF3cI5C1sUJkucqJzXs8K8X6RTsdXVMufT2HojMOkTI
f5Z14MO+eN6mazJ1mPDJaavjXupCAJTL+sNkpxwnK194vUwrkFOf5l1/+oSpVQio
P47fjJ1D16TJs4q18kOd6YB0Wx4gnLxo7JmDNNDmjGexWd28vhIRE9BiEoVegH/A
+OsS6wzyaFsBnOYHKOGtF1JXI5U4j/BM8eaTS390SI1DP2hEsYHacc79B3yy1c8j
kvWQMERZC3zNfpoFqznvDXICtLqf1MZtpNLHnEQfq4d0GEpwwLeOmxJddEwOqEMi
7+AELd5rz8BfzAq2dzvFSw1cfPS7VfBl3RLa8+6piFZx0QE2kqpwJtaLYUcNEz5g
i9hO6NHbdF1J3DP9sIevHELvKD/qhB3k3dPcbmiUclf2sy+/6SbRrvCQEKMw/7K5
kbIKHKYeCVTgeZEKMbsR3OkwRHatm9KPzlnzvtU0my26yCa4fkrXYxCy5OPR4qK1
SOfiQ52MeVSckg+WfyJkVBsUoffDwQFVYLGGLo+NeEKh0ygh0kbiJpFN+MH4Phxo
mA6GGvSufiCIiOuAXBB0nONzp6HMgEHa2hg4EVdSDhRAPnq/qnASZp8k8q7T4833
Pi+aTiBjOJMhfBFMrwIpy4i3NlYTa2JbP1vLfXuG23kFqQYsdouF3VKSEuOo96ZX
rCplrkMWpsLE8UbxQeWJ90c/mgObSQPxRVIDJM6U1wuy+E2jZMXROwiwz239XanM
4tBaotBLDZ/ph1QAkC9b6N3CmdQJSkkp/IJPeA9KaDapziA7CChhALzD7er59aDX
buSiUV+VmX0QoMFoYBXE4Zb0WJxa8FMGGx7hTCrghTYFzqFKBaJY5yUc58mfcflK
iC1NM6Uqn66xEe7C9WAUigw6aqVq3xB6xT9lnZwRwlIa0XgSTrB+eiZEgb88MYIW
EE3iwuWYV6imYb07YRSngEc3hzkmOnbYsPc77bwIRA5yp6eVykMVBmrxaqGHkvN4
8GfNv9m1SIUEMPg9kHWArs3e+guEiB7Yr1kbaWc7TYt2j6r4jDgx2BqWywmCa3iO
pHP+VRdoNMcGN5cHg0+UMFDehDJCyDUhuDDsaPMc9k3swMpsPddhMhCt7Yn/SJb0
Tqwz+WyRWh1IZ0R6UUJMDg29HD1CoggwSmDHGHiuU5zgXMiUY7k+gVzVAl+UaSyX
wpaqOoGUfRn7IskQomIiDKz1zRVSETFBCO6xSb3xZxrGquGW3toSc8MCMkMGuIG2
cNQ/jsw6Aqx1XnYOiHJNuSDKJZKqR7vx+2PYgLZ6k2IocvXnSok8lCexig9Vs8jT
m4yBdWGx3+8+yuP+3S8hiUEU4CpjGN/CC9Wlt+57mb8OxMT0NC95wPrV4jjL3ol/
RHmKIRWUVfB4mi57MORwCV1jxv0JgBN3TSZ21yJAQvPvnHHBZBUXZHDkB5KR2F5I
aklmp8QY5kNqGHkoAEPzKB19xNS7E58+cwNxTcjM+MNTOo2Qvp28F1vobEvv9Zn0
HgpujhCEC4GodyO47ooNMQqQLgMKvUaz9cG09tiTDHF9umeCtrJ3KfKTFKw8ItJ2
bO8ozE7map4hRmjG3C1iOUadqFc9DZWsDz4NwzVp2EgKumRbuU4mN8quP5qm0vI6
1X7dJtMb8HaVljXCeOgBDbtny05zB+ldbSwjzlel1V0RlK9VRiRmlJDJSqRKeQeE
nXidXhQc1+P6irExapFzTwttXCQpEtJE9yQD0OEYHd8CNIo/AvfO5T/VGSYuhiTV
n9nT2SgtcyMNSeGXfR7Y6W8qpxHW47dPf9guS2y/HybHSz5CWDVS7XsRZBgtLIFu
EZtDtVzqxjGb0yGeM+4tI3hPB4bXRUF+ccwbmkh2K7iEYBXHB+nCu0sQmAe8EjS6
IoDzix9WNKKIeq5dU91GWVO1XYtVHM4vJU0t9SsAHlQngKoQZx1E+U4+ANyBoHJe
ydrAQnVWfshoqJoqltIGOsF6Ik5rzSPpxD7tXyN9OcvhGrXF6gu6ZFWVy+WwaiU8
7wSFywnXpcsfFb2QFs26rqBZdJlkmmTxgBAm1qq3xNSi5ZDihJu+T4yeskqW2pxv
dEXPMFYIkgO5oNGFlGhHgr/bEzJEiQYetTOLyZvv2gb5HpczvIjfb8kNQaM32mfY
um8u16Wj56/8Z6Wq1E9CcNTWtBsj13hnzwe/JflGox4IOWoW0PoXVcrl2It6nK4m
6IL0GqXi+YhCajMEo8uOqa7jZ0TSNGWbVg2vS1vQY4d/XCyIhkuvPbJGmkfqST0Y
ihMNxkf8Wr0dSrTRgYP6acQt7rz/KeapYjJHF6/1ZZ8xm71cealin8Za4kMw0tD8
+KsB30ej8jXZ7Q89lMs0V76g9eEmyIt7WpLBkxF87BOjOuDLnEw1l/BBBwX+JUFn
uInpKUVtPpz7CUPFIuCPnIJ1WXdCqaseVPdBfrng2tWGzkE3jeRrQm13S0G2X1Z2
HMytKXPBRijM8stPHI/wVPrAkh2+MuvNdI9kXe3PrzxYt09bLHTxad67/Yzw6q6Z
Fo56QzdQZze28MVJMBEOqlrKL3+5iBp/GPzrHeGsBt39gFrB1t+dEn3xyIMcEc28
1LENj6tnY0VqtT3UmI0jy0snjoIzVJ64TXscMDu+XLhfWjrR6MwB7LiMbYfVOEtw
0kWYSz2atlWcl8dE7+ugFZ5iJNTZFqF2o+LWlncpGcAcS8EcE2NVfxTC1Bl7Hdvy
F6rY7aDXG3PIRY3AXEHaF7kTEH5uwiDhObRDYHlWWgIdiXhWcpb+Mih64TxUIGCh
998ExCgWYVhnlhwDsyTLVODnsYfbWxymUiOr/b+tzDiwKuj0G2kRjDNWdOBms2sY
U/NOlx0bZDfzFovk3wvp4y6kNt4J+97ZSewmWafo7g89XW44pw0M540mR7+69gPz
pfuqChnPh2mG6CKlKvwZ2KYdP7Do1yBU4dklKgKkIDaxv1mNGxw7bd5NQyOZ1+bO
wVOvt1Q2TJlnpNvksP4ktePf+J1YmxWt1giCGHpEeZRSAFg/Bszu2VzYhOiuEWDE
hYBmtqnB2I4sr9JgTNZpVthqsIlvRSL/DQTUZlsY+NpZXlPvGnCypvzikHB9jQUU
Wxyqv4ow0/yYlZiOmBNA65+a9bL7wwVwdoyDQR4cQHAKjrSYUaimEWWa+n99isXm
ZbsWD1PXOCH/q4PsABmcC49YbaumHAL/RAyDVv//To8pR6xAHazc+4zYT03BTpaG
q91Z7w90UVtpSpMUHCHZR/tDu292zTHI+4PzI5s4xJUwsFHYx9iZ7hgPmjxi57wa
+cgooO0kdU1PSlF13EhPCQxdvFpMykNRdK8TLsOC3+e8QpqzeDNq4+OMXOWLF1lB
S3IicgtVdSTxOzOTckAS7E0ZHr+C5mD0tH+4xDrPXHSxXhz5xWe727z4H7qiTqiE
zrrvzGn1b2pvCD5Myu452Mq/7EmQgJRYUDUVM2GzqpQSFD2Kkv9XGUclSBEuoJUt
zeVpK0l9M+yWiV15Hri32hdaVi9ruWOVgFCkxPCHw2eFrNU+c5OeqaavF5+IopL1
J5hA4DVZu6J15NrO0VUtkErn4BB3prQaEaKslPJvb+20SYIV1giCqIUovtPiUGfx
0ftgq9ttF7Ta12NviW1atkx4atWwIUzdIlrsF+GDnaPScqPOEGS6pqb9tGjx8vEf
jGNJ6EtIoNXgDKCeFYmsvMz0A8LsNfVuraCbs0pJAPyknbTz0wANY4E73r7202qb
mL69M1sM1LDNXZF9MrNG8/NnWsuCKMwXn+xmhPGtnaOPIAo+0glyGfiFyx0m8vKG
l9+91Jr9B7eXN8AynZ6x0C/XGIhQRWphurk1rlH6YTn2CwxQPZwFJiF5/lx03/Lx
inugbzayfOJTSsfHpOtXEMJ0e3Vo3kG9DC43OvqWM5Q0xu3AmGfk7lAtUPhwW/hA
dQ+NCy2y3Mhn9Kuzv0G02VNOLf1i1oyEGJsw6V0QoYEFEYQ6HEUbuDgm1gk8X+xL
oKIp+HFP+u2eboTPAjaW816udMItuQwysmGdcOpmS5OPHFLELHtwhBrLdgm3gs8H
+NPEmm3laMEge8v189yaA1HVvgluDvOZKQj5oWP1CXhtdwUPAmsYjEE7ldVz6sjF
Hq+g8InB5keN8666i5hJt9pBxmCzjRxzkGYk51l2nae+grmSw9eNNJE/rDkY2k7Y
Z4Frz7cc/fPLIQzS9KBTW1H3+FkyO59jBI88eMubTyLr77xxUyfck7RUV09AyPP3
mk/gY+lCILfuFXN5MrYmUgc36g6MI0/XRlvUzKBE5ZLnS9QAzmJHacRSLb6Y7gKc
vcmNT6pFQ+b1QexsCLO99PIAsqNA/OlOgBQP1uZF3IbNLvaL2QIixq+Vpp1pbiGt
FOeNVRW84ZA7RUoRAjJhMVgVlW+wHuYYzX3WhzC1qiLnlNZq3CkMRNRDVSF6m3xV
aFypSUUeoh/xZZ7QVHvA9RlkYedfakKGc4cPoUuP8RguQE3ZsLGa/MkbrY1Tq1Dx
dGbdPMbWUeYcM8seeynOd/JThBekWyZINmyxJPo+HjnJmFHjrhv5B0Lh255J/Kif
SrRHGYlFBHqHB793pKNEPvdiaUDnOuYeIPiW8gD5Rh6/Sto7JS4AAh05+LyY1HNG
MJ5Bf2Hb+Nlhm6Kkhl3cSNwzmZcyQU9/LyGlQ4F8pQpYStnTgu5TbtksRnXv4K/0
vffe+FR7MmYkc6DxZWVDYEYKiKyZ8zAiX8jrE/7unwOWrZdB/vCORzDI4k5ryVrc
a5bnJ39jV7vj0tM7/eGzXVMPcGXOZ+FL8xIDUDfJI/RvLOkIuAhlGq0c3c0CG/4b
z4oiWHheESVAW728HWBl3qhWaqdSkIGki6qVSTKAMUtux4zfejjbXM4F/FmaLk8G
w9g6/8oA013SLSvx6SXviwlG+YEKS1Ax4iYvz2SNGUKhSHy0DsP9oPQB3nvHTPWY
eR9jfCmGaZu+WGLcEcMljv5qwT6H04GyCGgq6HMyON5lA6JzqrU+qRtkBaGbWr6P
I4Dm0Vo6nOZiZVWl2E/dEQBJa6AzGzmCWMNVfylpwcwJApSLe1oRe5bCG5qASDhA
HdKQIw8+ytZ+2cZIJmk12UyGyqvExVyvMdR29289MMMrJVuT6kDh6lw0GNhL/xhO
BfpzzuKI1GsxvKBvU9l76/3QA6r4FHHXD6cvkld3MiGjkoez2AZYQgDZ2l3h7yFo
6JWbGp4z4C/w1DjkJKIG2CuFa3PbuGfxIkD/3+vjfq53yiWQ9G62wZECHHXiK8Xc
jzTaBNMoJDjMoaz2PuK+83t6lb/GRhEjrCGrxIskNDXr6SIOhML0QGvhZYNLxN7R
tpfMiILOn1/V5ngeqZZySDy+Hwq/Mhm7rRZXdHp5k4/CamcIapbCjoDE0YwvlBz0
P/WB8qAsAGsfZT8iF81CsFWPotdmS4wjPA1a9ZJ9CyLQwkSMhFIbUzBY7xr6hqb1
ezwKfZPYeMzaZo9x3ep2wrLF7zfwXej5qnHohve2xeZ7SI6xc+dB1MY+8HwXruBl
IwC0eebQARhrV8X9mbu4rqcbSt7a0AoZLwjix5zKsOJ3MofkMER8OLWwe04OwUbQ
Yk0WE5NNTw4Sh0VW4/fOP2bMFrxHNIMqm98E76ck3oji9rB0arw36qwaMcbW/2Dp
ZNvhFEvaPFAHHkVv1moLp7Cuu0l4Fv8Ndcb9my9Tz+uoD0gUDx33+POzLoReg69V
BrY3rFSGh+niEUzLVMgMtmK/TnYcw9StJmrpPN0762dz6mFXuWXGHObBUV5GCh+t
demUAXOsroPahpn2lYjenIpEhYhDjNAww2z9sPlFYhJm/xp8mOX4lnMWSDHDXo2F
9dtr5M74QPEiHK4ny9+hOYFuZqQsyJn0YbOVL7nU9mxAzg7/be7H29/ePz8JdUwj
dNfZK0q1K2yv0r2RIw8l2gwtrsS5ZGo7eg08HjK4lwrL4Cs/E0qw2lPBP45X7uvY
rHEp9hMgHZpV5BsNDW8mkAJptwRHB3iP7I5VyE1X7qDkKGQ3aba6iMY2EHEiq6Zn
wHtc3MnpZL8+RGxvMcd7tKtYdBwITzxCaARP4KA2RgryXB+QrDoMmda+JLBejVsH
kbI4xagGHlw4HDOheY/t2J2eVidD2Fa2ktfSXt4yhYY+Jz6faAzuyZJy5QC79qRu
ZqGo/aMe51UcjTabMhs7ulevj6jEwT1JP+gDZy4NKaKHWu7fCodLT3SoDrA0gniu
jje0VzQUP986HU8BWZaWya7jXW/BsvJbsWngoYy5PKRjVOPSGJgX0scJNrNR5VDA
NoaVk1XSqfbYp3/m9f5L9hzUwX/yvVNcHrv2KMtko58N3gmVrhZNs4g7MObfk6SX
ZGW8wQO4dCnkn/srRMrWKBuxgH4bGtfVX7C91tmO1CMboKK6mc8+p4k7l5koQdFl
BU6eg53VB9AXwTlvY7OlZmCI3Ft1TyesQAbXETkF31jI+EzDvGXNXRy+/uwckdrS
FodgS2gVbp4X+gxfv5DD8DVtJ1vIKOZ359CjbiIYZ/iEjlzOiX/OseGWCK0+GNMp
txAljn1rHTkvai42THMsJKtkt3j6EBmmw4YDAndq6zYnSdRGvTGenUFrH8AJvB9i
NwkLBTHwf4FABZ1pmygRtO0xuA8w5/usC9FH7MAMu+it2oEjXA2igdKrFyda/5BV
7SMxymu3fvgFn+wFuQB0Kn0BDaErScOkqhrz988aJkyxu+ZOBPOlGf+W2OV0mWQh
RQJAY+nPfDJHV1Eam1l6d6iSjJJDrlsIVqTLf+1ZQaCnviCDo6T1l0XYXiy4HXWZ
uDHvzQ7YqTm7G1TFxZZxA4VjuCXt7B/MUC6YBsLt/Xo57rUbFnf9w8PzIMhiALP9
7NiEWGrD3D14x1QEh8gQTKsUGqkSKftgvsvMUjNBI2FuI5Wx93FVQP7KY/NO6BRU
/vrnPQ4A05TVs5AWCslqtbr3rvI2VNU6hjpqlN4dos9OWTebJB95LMFDlDeeeN0e
JHT0CzOKKbgjPX7aWRQQ/JGOjUpYUjjsBr9gLTThrNjysF/UcB2GB/37LOfZjZj3
cpmfV6O3rcM1PW6MDVu2NKJK71NSJI578TgzijeE0MleEm/eO0IHgwSRLIVWKEs/
xQjuNey+32DI0QHsI4bVq2FC6p2SSirO0/07ixHIENN9Ujt2fPJBG1RhQG0iY9k4
fUI9edQGYXFkGVEoO6VGC20Yu4Mt09Y3ryxtK7Xv3nnedwwC8gdWNZ5eZ+SLsUKt
f8/ynQ7yZpZRU1Ot3NpafXqN/CuTMNixKw2WpM55a3AnI6Sh/zsHO0/evZv2CxKI
Qchk+QcG9FvXc2OSYwRy3H0cZxkIrNesoc8BzZKqNsD6jnsplWz0lHjUHBsHhkIB
w402VK2GfRpbpVDc/lHtUZA56PydtHLg82SeXwIvKxDnwCV8n/Qbo4nD9zuavlAq
Q5KgHI0LyMW6Vc/XsIqzUNXpw0IGxvQcGpM92FYTbDHrhKFFk5VlUG84tn4Y0ZC3
xlU33YaArG5WyVwFf09FGd2ZHxS5mx1BnqEPqzPGer+PzkQxpwL/LiM5w6bAfh6W
bO4MZdTLzK6AxvbWzNtw8lSbgsgr2RNkWK/YiTSpLg7Ew93agb2Zd9UgyPVC4kNJ
3qJ99hFyMbyhW4PUwaDSr0sh4rS2+DddzYVVyswDpFybG2HML5DLHF2hXc256/bY
oV5kOXveferRbH4dgKzpqueRt3R+NQV1MRl2xVPYH2p8XqekENc+RmGqJtOVbbG0
pGK+u8K4npQnB6FqTRut02rYJvpd6fXusrxU30TH7bi4jowWyIaYhVkm67BmETvm
xNQK5prPGRiG9BTCa2UVK5NIqXKBaygnu0SeMQIjykk8and3ja48zDTf/hhV4JmC
m2/tcFtt1f0W3/7JEZpXPWz6m0HdwHHeFD5pO560pKJPI2Ym3NpZBYe/qR5sdpeJ
htEh//d9y0otyDEriSvfS3YaYyM42fVEXiA6Cs6pxNnJvcLTBbbBXytAdzSwL2Qp
AokYOVkpYdyQsP+6FcviR5QsWj24Mh/PFaqpXt0u9p7vHG+HEpDFEzS0Fmt6QTTZ
X22GuFejUnYMxf5k2KX1tREmL7jZyc+vRzxAarzEjPEH+0GSrVNQ+1SwuAsUDWSI
t8rpVGQlBRMsW6Rxxr6v8LPlCxcUIbQmsk1czJoBBPmfstiJVzvAeYZ5v06+PK+P
VJ51Bn5gbMqCshsxf95SHm/nx3rBYddM4KqUwcPo3Lv2kiCAYzLkj6fe2PcAhbIp
/xuGLtJ2I9DY9aSPs0IIym7WpQQehCklazJqnCb6/YrmHmqc+WgXZJB22+jFnEsB
G4USZQ7y0LkKLwv/x7Itc56cIztx3cUPO42gEwuWaY+EF9MC9DjEEzWrwQxzWYrZ
Cq91yAXyaTEa5EYbH2Wv+BG/orH9aECN1tIRuhMCMPz3aHFFpy+rBBGZNmBlcpNx
NbAMkYHUv+6XUl2J8MJw4c9OUGuywpzcIDtOs7TssqiS5tRLpDArE2yTrOCer9TA
ICf4ddP7luq192n4U2k9BuE5daDPdvWh9iq/P6rH2Kk25DTzi/4uYWTSh2ZIQrV0
okN8eqcgAYL3TxPks+akUEcDPK9hdsj+fGo4vGl9rC9TFL8VzXB1vmTR9zAlfJh0
eP2VLuM5wSVJTxxPfcUw1tkqMoYeRQta5fmODhuuvfoWkyoRsul/l55q7599qB86
5FvwaUnX5dHFsHjH3pV+URkr7z58cbHb1CB8uhynZwBRtkKxLp854y5RbLYwbXXR
kxDrLeMJYmQKLGT6OeMTSmoCFcLmwelcrlS4MFza14l5gCJ2nAEcTSq2UT8EEf2K
KlY6XSrIL0kGwXpYwT5q6FeDw9kaKWfGY9rhNFx+rXj28aGLu5Fw8wYBydoc37X3
er8TJxCYBHcefQd50UdwsLa3pSQqCnX7klwNdBqo6GSYtLRtVJKaANQPDQHGRSz3
No7o/EY/6x74UVyYGqsPY/I0orxkmOnyjrMVelNKNQoUBpEKpQU085k/GjqFB9Ie
MKph3seZ4PImdokgsvuYLX/QjDQOL/SSI0ozbO73LXrVwh2frsK/xHwcH+RAHhlK
gfCdl6udnJ66oniXuCDzDLYMaPLXsmJizRRqhkIjWanmt+dWh1ljO1QT9Ckct5pp
pdvDap2zMacF6fcno7ZxIqiH8GRNicTMNM05MNDpA2w38gOk0JR3niUGvUdEjcjg
erxTbDmTbBFtl9jyBp0Qmp46eUX4PgoUHpJuStlXLBBYlU34VMSp4a191AiK2Zm0
PHeS+dybsOKIwDbv5seyxfQZAec1KXlIp72ApqRo2XLQdNMbSy78jL96wc5ue9D4
Y463iA/L/wDrGadfn7BMTu5bfkIuAPD7eBr77xxg+sNqayETUSrCF/o3hnTRE0DE
bBXGP/Jc6YG1NZZmqK/92diXp64YZsQHZJ3T6iRBc/B3k+CeMkRfZZua/hvP88Ms
JUHaljY1uApZ7wC4+FJ01Ehd+aNmQEoyN234eVA82yWqhtp0EX+7EmJZ7EGADCsE
BLYI46uvKYtEMrZt8r+Q6PAwF3iSiyzIxJk+x16vCc4f2Y+IeLzPsX53QppN4lwQ
u+k7u/WAzMsVKLds5Hs++OYkFjN/aqDRFQQ1gwI0oojGmX5gawr7YhXfwBhX50pg
5VsXGadbgl/LLpRASKNNsdE1cqltJJE+UVYAqo8/eBi1P8YjuRKx0s5UFFz/GWXs
KXS2yzen0v9NS6ZozFGF2ZawfTTPFgyrJAiHn6UpKYFWBJohDnqVIC2bQ/RBr5cL
+mm8bEkXJOpVQD9xeA1AJBGGERKcJSAWpCO0F513f8LS8skQJXbceg2hveag8pvf
+KosLvYlmbJem2L+YNsJNxhuiHnBuVK7qH7kLGiyFrIUPIQRG1wVwBptDCpF+y1N
8zfUbq2gGWNan1RRsscx3djmldpEo+owi0nrNvmAm3Gd6LZ9bA0uLTthV2LeBnfn
7XCHdxc7eV7QLOqIsrebFZZfA4IS6EaeCOZapLRbEM20eQsr3o3fPWTYDHM+MlAv
IQNE+DLcy0UcxPFLpOs2LmPXrvAl5JFYhVD6F5Dz6RdhFlb40VFclNkhAXtWCq+x
pdyWQHe0tG+o2z/Us5z24MNgdfVAz6V9UZ0P2KtAqsKAM4ZWJWQ+Se8dm5Zod7mB
LSZY4zoH8laPhGvxtujMv6ICoAI6/TAGTRYtK2qkX/M4xYjRDngrpG4dEiKvfaxE
uyx59lrnApSRh3ywMNI2nCB8/GBOYcqXZImMME7JvRELzza045UO7fe66ViyT5fK
6AiWoAGk+Xi2zGM8lXeLc7WenwBp6DnApXSoB/HnVFGTrDnNdhMcr5/XR2BTFIOE
2wSNxg221v7YnL/l4oDZiR80cQKXbO9XsX22CdLUvDDffrEWNBbh1kFxZES+bIG5
UUHXGsXirL0PEvKDegQZXbpwBm6VDchcrC1pgSIJcPhKaJQGIMJrBfAhUQCiPyrN
ldeFDPP+38NDk4JWyjuWtQvakJnXG866ulf/jIWNDBEEJprKLgjFlk7wop9S/Cpn
m2QgTYUry0oqWnBhvJKJic9TpByvWrx02o7xLRjJylsg1tovS+pp44fzHpkMbMxN
si8zp+D/oCD19bxLB1fAyqW53opCxMmLuhjLXgepj2Pet7wzdsVCb+/J5rdZ7Xby
wu2O/gVmmqIZgd6GP2c0GBzmapdgOlZt91F+OeepEBoL+M1Sslzx23D/+IwJN2yU
5pWgBFEam4O6B87Wv/Y9kenm2P4V9JBlUstIMJCMhy2hLtbjmsLNbpnTZqB6kYyd
ShO8e7X5JGy6aHpoCtaBd7zBj58ATwSWSuK5XhiR23YlHt+ov78KsuQnzuUxKBr4
DEorxyUwBFYthyXlRFQdWk+AcZgnp03WgQ543z7iRKDPhCvQPkyX11EN1T4tAtk/
DcWO0L0+W/Ew2vL0p4uSEtx3xIolgG3du6MhQINgZUaVYIIOVkWHfI9QEHO+Ne1A
c3t1NDETt6D9OZ9elOcGYbSSI1U6wtqzFdQxj3hR3DDsr2Wfkw1YyzSWXzc8E8hR
xaf4+8gOw6wG2o4/ReoDEpDZVdx+WIioK3Gt7BU+impHRjKoh926HofX92l1XJ/Z
AFksWUwFVaIczIy7hu3EWM3FkRZfjMMUOUFfsM++95laBLPO/+yGlcfCCzNO9d6b
T6V5xBYpiX9kc+EGH4tqJ8iWByUHRVsDwonDyDvVAa2rmrIcObilAd/Ehx45rSZk
Ao2l3HgF+xk1FxqOUik4NK7e1XvJLirEP3DQlgPgRjcf4qtaCXXHqC0VeKvgfdL/
CScbyHx2BVc92bYfuQYOe5NfMh/ySI1MOylPHOkFs40KQ5T++dvymP3WhZadYNQS
HHSPbY9KqZFubzxYjr/tOvoDzwYHzBGeTmV+FM3OYELpjdp905qrwco1r2loEhk0
0blojaQr0F3oZqhqH4/b9rW8KSAqgYO3GWQCb6Ydopm4NE4B9vtwjEhVN6j0QiGT
g0aLhbZDcWrSIzTzyKvCup7ykGLWCbYuAg6/2MICfoxbet0Z8YHyGTYFqGdrwvxX
llF/dv0h+PxPsswxGhB+hSJOoNoZJ///d5d4yfG/NnyagaATZeH69cPdfcpiOCL5
59rwIuTRn/mURKCpqwRDLuPUa6is/NYfWoThUE+Br6LQwhrmUxri48luxP+CgDV5
VP7dWpsUusUw4T7cppHiBkMBjSk8kfUphoorFLo2szFCjxNYARU2PiqSe2DD4Zil
5yc75EnTF5ZfAIwBTEQQ+UwYzJ0Z+rsQts0MLE1JCsBImSz3EvAUEk4CDaGkudQZ
qmnK3F1+Szmhvol13cVUwG+p7ar3BdgIzu/BZlbZ4Z+mC/9ZbOV4xN6prirlN35q
EX5SOAygApIoOs8h2XetJM3GvJI3eMjbdRBxjWdJQvO4YUrb8yzHyZK4deA98UEi
Y0AkcRPjHTFqig59Avw/4/0yIQZZOCwYJRDV2FosVflvcO59qyCEvpYazYVQyVMZ
IPk4CTobRuhX/UR/jrf5JcjgUTFT9vNL8SXghrBTMZW8oMFMOfArVFW+773Ia9R9
pTOJvnhQE14+YEoEDCNlPx8z6fnCvUSoApj990oMGrDbMrofHJGQY2TS3eHI3z31
K7Rwk9XjAiYsyOl5yDmF3OxOjN2C1eUk0jsqswneLM24LOJPN58PeV5sj5id0wQ4
0i95m3kzdTkh68awSw9ZHEjhuUTbFzZh7Fs5VtJtbvLh9FLUVTLlHUT52Yqbpud1
2nD0egiL5M/3luqaRFrZ+aiokF/mc1leVfEIpeS8VdIVkAhR+z9OnXed2PskQO3y
Y2lDH5m8a/uH7sdySNkOtq3Yb6kF4GqC8zwSSnv0o4O88yA+0JlTp0vAr70OkHo0
LBX8h0P02X8LDULB5ma8NlvgA1TKvnW4jSOKFqwoV56prj9LWZyeMf5+jD3Zah4S
tDLioxuD+UchJf/wc/sYN/ugk//Aj44qEQ5DXGILJx10NMZv3vY5GtJiDTNL5XMf
ql5rQ+oxPITmEppgamGLF1R24Wh2aIagsBdRyvlGTRIGl+0tYO14OdREWb0eJcnp
DW9mkgFuXWwIxRP76cpAoMZvNMxRZE94kNn8Si91ne5mXQ6/RksV9q9EChrwUmnB
eBDxDyJSEizbKEkZi0gQrFtfLo3rdqx2oCEoQ+29E1p29BbMYONQYHHzIXJQnAnn
M+XMKdY8p6KJgTlTYB7aJvnKB6PrRaSh3uOrebkPNSVJwlTErIaw99+1OIYfE1k0
0mTDmvmB+XS1BIJy3F8pgWHRe+mWi/O3kuG8UAkeDYDmaK2Gol+rzz3bbbBwCIsv
2FRZ0lmSr6wMWEu1fuf7ijFfdfYCx0Cx31VEfx0TTl+eKph9GKbRxRW3solMN5eP
jGm4dF965Uqn2XVFYkmFWO+UGHraZC9igRxVfHeOFaTj0oTJWUdozw6W52oCl96q
zFZkMbBNHZr6bJnCJTQBK9tXXHucFLntEUB8eNLbIdbHH9H0j9WuHqKTguqHlvlm
wRXBvRWWYIGEzdefiqCmJ3/JbBPXfxV7IAk74eHIjLyctg0whD4EJ+Iv/Cx5JfSt
AhIi/oPw0PboCPCvgNmw/UZQooqAjuBrhmE5MN7t7YZl/LZrI/yhxPE06Z9ynpAY
I+9pxmO3mfpx+sMlPoPaUvqVrNex0oa9jkMiCYrNEfPDbu4zav8SCrhbjkqNfjOr
+R6VOLpGlXMkUpRB96tlcMEK8fwMNrGb9YJ7VDxXQSj3taKHnQqm0jJrtdDr2n6u
+Z+vOGMBWC1EPntjJ2onBqS4Eg8s8YQ29eznSodbije0olb5KForOu700+7VHrhC
3A8njdMT3YDIxmnXSVrcV3IM6XlvOeWvXEEO4KpE45EXXNq2dFzNWSvWv8kmAw50
92XZ5u4tTI1HbiogxKDjcEA2fzLLKgiy/Fh+mULNMu78wA9vh1q87ff62hhiGxuQ
ejL5F33eN48kwhNTw8aQXt4nKhFrkY6J8S7FMYeezTeY8veXZABRXFJIO0J9R27R
4A/hrE+Bzpb9wjYNnehOgzzDBKMZfvxgPC5FC7HbvQwY4IvkYMENCzbNK8rOF1DU
RcVEzb8sDwG/OOrHK7D9tEo0iCKKOgrkBqO12KhEK99IIHAYPACcD1/W1QPZhuOC
BIz/36E2y9fLcDUE0ik0Y8JULLjHzgEV+HRTlP9rf0Imf43Km54pY+4wsFrAlUag
WbyWfEuzDUoRwlvxiQBsCtBsXQRO5ynZX9HV+Ugr2gUrMVI6fM+06GG90+vPVZAB
9onCR9FL3vNf46kdg3GsYMKLAcyPGb1u5Ux45s60j3JF5gf4cmGl9a0Jk/8vuFRQ
68OtzF2nsxhA6o/y5LuH4igjDJVdIUkP0LL/rUdPIhVO97hq72jmokIAi5wL26gc
mvooQUTbhWDieY+JEGaZ4ONNZL8h0d8OW4gcCTMIY3qRUq1BzL/ywlY+f74wMX7v
5jQgdWAdN9Oxr2s938LfxNQLwNW4huJSHti9wmpBePIDhe7/xBF32j0h2EE5j7zr
UFlLJRn3j1FJsIfooE6FrAXAs8LyELMiz4ESMZqpbAdJ6+wPq7VC7KD7DFmSXFaY
mLW2ycNiEJ8PjZGHS3hYiFxQraKXvYoRSFajPyeiNJseMl58IHXcqBqo14uXGfna
s8+1LmUL2+vKTTmGQ1nf4cbx2vJZWi0LmnBEU78BvKtGAcbZjHIqIxMv08Adq4ub
2y9wxe6AxhddNEPLpYpfOLim+XJzs31oIAZWDQOtacEEvw2qQ9jvS1bMWDvxz8q0
Gb4iamzPE9GqDU23U0COKF63UeNldrh3JmjAKxMcBXR9KuoaNqSDgRNdbKNywWs/
uAePr0a+E0729R3gDUEoJUG2veQwjuz2aKYmG/brNaORzO91pSYn6dO/bqlDFq3C
F1qo4d1/1z1CakOFiLYM/I9UAq63KtRzzTf2f0ItHO7zQaaJGt3YZsoeA7T3NvbX
LCQLSN1894gsRa5IdcXHDJmvJ6vXmRe/LauNunI5NL56jHSlJdHuX1eTjSqaDqc/
vpQ4Ufykw3SUDA+qsNT7GgY6ZkpmFtbH3TXjUtU2CjgLEKA9MDYo7U/8fhbbBx2i
RnI/zKZT52Ttu2VJMfmN2EeTsnsc14l74kxXCoXBmO7AlYJp1QXF+zPcWdK4RdYs
k8uXrUoVrmq8475UarakDNQE3dHDHhOO5bnSvXfT5bY67l5bl6yoqeweC81tJ5Fh
MtGe5fyK2PbLgU0VkFxWsFegjy7CzzN+k81y/wUkA60bk90+crxDQtDoCVjKS+Os
360yjqThf2IVwjeQwNdICg7n6xYMQvC/ipw3zr1xaHgCdXZ+4qcNoN1cNK6CKF1G
gA7hRtR53UOCSaKfAIb+jPoyePudjpebMgtKtvXLnwhAFC7aw642C5zGFkDmj7/o
I+u8Xq5JRNOZOws5BfCelbORx2UAAto3Mq2bU0u5S2Vt0yJIyC/gxs+MWo+qXy06
ckvBWUec8kVTrEE8lLLKCh8ZbZ784u3JfA+gmove4e5FUyTfzq1sFe1Tl3YGbP3m
msdwNMsp793v8dg+1hNuhr1A7hnGhuC5Y9jTtCNhu6sDTwW+gnQtBsmjM8OSLPWr
7iUUC0QXEHyDIx68hbSU+Vi6fBYcIL3CRzAaVIAqxCtuEScK727EkZ7OllZdQkqn
pZVyZ0aoWW36qwvWzdy6gQVDDHis2JyiEbWQy0ygOXjzYps1WSlEL42GIFnJ157a
wpAzTug/Lh9surxylaG2EVJl4Tt2JLKsMcvgzC9zl65TQpFzh5d1czCrR704KG2/
nkzGqP+AV1MXqMj42DF0CFWmG+dRxeADgVQDJfdTCFik71NUBnxmDEBLj9Tll64Y
Tov8AumFBs2Sx0Yocts9Fshg8GP/qyjmoVimRE0WEohml65ktR3ofdbJjeeGR3js
lY/c/yrbVPH/80OaLnjkab/rfzv6X6KSXkcK4t5oh9ievNzSjUAMSBtbmNpOBswi
FZHsBHvoxY9bOSc3yv2G0lzmlwO5Wg8P/1yfm6qhuhxEtsM26HYMZabiZtwHRjg9
0w4qyzJl58vnv1ep0wM1V+B3NXP9PM4N5UNnIiA4ywlUVokmf5IO68uW3/rxsDTd
Ndpzf7GUWyo++lgwWWiytsw54aBwhMo6bcB7DrpE2oUamOTrv9h2fWPhkX17isUm
vGdk40Ny7OoeDMa1Pi9Bn/2AK6+qtGblsZt6YAqOJYHvsAqNSlEQC26Jg7MEIrwI
Wdu/v2uVja3nCuWLWb3n9Wj7rfMjc8Y7+lWCzctUXWk9yQCFxcP6+w+EVs6PhOTd
zcI2C4Px2M3sexKUhaRe79qVdqH9ObDUX9217gm9fmUwb/tpwjhOF48NiMv5CkVs
eRYKh0btC1PMdYITd1BI+BfDPxZraGJvgDBWOD+w5Ab5zjW8YGUb2ZhCSlCxabA2
TD7XcdfrQsbcSY5Obp4CcK5fNjynHTrYO1eLtogfgPpxSh3G8xh3tCiUUAEIvE7s
IUyyMGWd1JfdtZf/w7gdAXGXWynZVC4UH3+A1GgxjFCZ0ALh+Du2Vw9r0X13DmBF
2oSWHJGAG2BLs0rp+4S7DVs6zi1baXFrBYmAotRczxC34ciodQ/4hGDjIWC3OA+/
VAgnT2tTbRxF8GDaurAV90Uk9z2DmB8OpQ2JMZ6Ez7FVUxsWK5C6BmtyZX2P3S3b
+AYuTnKbLzqHLtmK0u77z/EZVClrQgaQEbSd2KR3dOgy2gEC3rs635br+/E4ICeg
vpesQtNnR6V8Csglf2a3JDj7/3Y7SWX1jdH7C28tNn7N4ikM0Zp8J3BsfO88AKwv
RXlO5a/9jg0mBdGdEoV63Cc8XWeicPVEpdsqMalRqgHBNfbPM85TcUEem1ht2r50
JKVW9LHDAQLfODBpMwwESIArk3AVOfhqn9HuddxbAYR5YZ4yBsRRdEX+u7rDSei5
GJvkhMCZtFtOQiQDiMrS/YhWLmvC4K6gRwcZs0pZQPGYg7/wuJUie4AMtGkJ3ihk
pfqm6ogF+jLQ+2OXxdX3qsfNxY+KvarH0piDPq8yvqaYiJkwV6ILbpENrHaUWNKD
p/8hzLk40upnLSfmFJJ8mfr/pM937kDE11bPcKOTLU2GpYl+x3OJ71Crtqrberyi
g444l6FT4/LdS1amLzRVISIbYK7QGAxpRm/gY4hDnqQmQnPR/yAXapDopvAa1uZl
YQcFRrjPALxzDsYwszbZYK0qjGv62GqjW/S21tzVIu5NYcujJ7M5gaQRp4KdAx0o
XcVwjMryF6GG4MxjBhWHvV34Qxb52qi3ubHOWfbQg9QCbr2Z5zFd5mUSsUl935la
c9VxVo5l3F92l3hUewVHy7hvAq5a9aohYNYlMMAb1BZom8mU9eV9zmyASeKD3VZs
XZ4Oaung2yCrI+tN+8tjaG05rWEXYNNkBJh6ibXjkBSjtLh4CJXg2rJTn2OJsMvv
mAOpvB0TjNDPyhjcoyeZF1kDYCAR0gwleZ2ALWk2Za8ex8hcYeq9ldL//F8UymFB
NTylSf7E4SHf8VnC0+O2MX3xgMREAZxAsiARanjKZDkU4C2noMhGl9nONJL1arFh
eyYgzK8YL6+dVDpQEXGZhgxmKQQzAKkQUJSi6wV5+7GAW9gGjUpgtxe02VNJ18/Z
kTwZbTYI/m2o3II+C9q/aOjRnK3KwaHxxq/tHkT96tDzlPbe8tpNTB8wyRg3kndO
9pkCmTag2dxnO5HjX/X+GstSBQl+qbH+I0pL8jsSes9FXgE5nx83mFLW8cDysWEE
mIdEnrlVtW/H1t9FpQsBLJdQUV+31Bo3d8ljkwBhLk95VRr7k8c5AYdwzHKkuxYo
lH3h+CRaJrENY2naop1UjNO1R8+H3339j8cqeN5MkBU1g4GDlMV52VdH76HpjzGo
CJUCDUXRpiZXuv7Fvjt0CHdH7VP5qs6cCMDwUR7o0EivwXe0T8Ly2YpmfZI2Rx98
PFKMPtMU/R6dgW4AUJvGpUjBd+d7a+VemEOmCVFcH1NUewh4hcqne62Ab1PN/pUT
qmAmw5AHty/BLQayZ1mF1nkziTGa7XtLR9NP8V+JUgmYGKf00vIwI2QtLteA8gvI
qVPtm6OXnOTJXKZw6ikjXTbVkt4C+whfFkg+Z5lj5cj/wSMZbFQWg7cK18hsu7UK
qdycB76Y04riSMxpjRdhTWnXR2Il6f0Vz6hTwbKw1ZsIQc625HW59pL6XG/iSVcQ
uLBI7ahLUCm/p3eFJu2/1NRy04ylNEO1jDVkZ0QCbA2uGHUD1UWwQUw7V+vG84FD
RAB6cD4giWmDFZan00tP5BBrBFU9oQSLmxALn4/c/tBe63mNX9c3yVBTQAWuNkjB
M6iFfO2CDX9MWgt8/c6CZt0TVlt92cUtl4yUL3UwRPtzU5c6ic+/rWcuxfhH1oZW
a6a4n0HL7jhOUcPfIp9EGQ4IKMSGiTXRmfACN8ymft/MSGMzusq3CCn8qm8q3FPl
CS11/onSA/twy7xl25R24A3DwJBrcJ1PhZlnM1r+TyX30H9rdiA2jyGfcup8GeDI
q3PjwofPxhiifV6BuUi+piTZgovQGZId2PL125RjctpyNAzrNCQZEoSA1H2vpeIX
Aw7tuREb+IjMI4AnYYWvry/zyU2LKwbvebqcWkifLJ3lSnFJiLWD+4uiiItjZiKT
TmP0IBzpsDwFHU/eGG7n0Kg9+AFgW6YjQB3d6B0dU0QaMQL03Uj1fJ2+GGMToxDr
z8iyPdjRgxD1TtccNEBitdyUJX67zg66hk9qHTFwYVXE72uadiaMnAkLG0YbyM6j
yAMCXRTlT04+l8QTB2P08PUFJnMPaXR75U1z18B0mkY+yfiXYSPfvgm2BkE3W5uY
U+9vi4o5PxiPdcmF9AwaWxL67u/MnsmY0sn/0N28722sgnRPy2LCMBUoy8rQRe5T
EnygBgFeym8UNcqejoIBQw3V7Yh4JGPSDmUXr+rWcK8QnInvN590VEpPAgt5R03R
EXT7XAPI+2cAq8QEsbVP1RQWj3x7Qblu1AsHRxHzFfjkDZCLm0JgFaPpvv6UxBZZ
/YlIoEQBFQYvdRx8WkVCizRD1meyv5r4g93+sUulGHW9+g1TzmN/O8ElTb8b5nhi
cLOk0NF7DCwZX+qlvpD76J6iQW0voO0NS5MyxVdjAHYnX4/QrET5mITD0Ji6AWCb
pYWfK6jEJhWe4uHtg7WlddL1rCPOKorFwXoWSRJUmjldP4ii/UqyDyuXpqECDRS3
/J1s53IgLGIATKiiddUlkVTOFdZLWqHNvv9ZsliVpD3icuYLJJiih/T0wm0yuq+n
p9fdGVpBDys082VHbnkR4c5IIN/8xnu9J2ot8xFIMrRFq5LCao4lwygbv/ipMoIr
R3ca2QTbPdssbOtAdCxnSOoKoJzVJ9sMb1wxK3Bc2Reuz6yQLAdzq+IEHn//5LfM
e5HIv6KetpQRXg5ARpJLZgyAZKwKbBpTaL5NQ795hnkjRRbUr4nyC3e8r1KYtJot
fyRODBVIbs+MvjFKOEGFenaAFWQfEPoXBOaYoTOfrPEzPn1XrVDsUdN1XVErkP1n
Eo+zTh8JmzW0p4vH1Zo84N8JI7X8ZQ7hf6GtbR1JEg0ja/zJIcW/i14RGUJDW2/+
Jtqgsr/fBowN2e2DD8bm/ZjQpRMi2eAIYrpzNsO6rAfFgDuBcocr0d9ikPrF3F4p
ISanxi4Su+GJQsvvGCNkrQWUQLtSUb5/sJfvNC+DRZTqMfYFZVwmAv5ejtys/ahD
E8mb8xyGjgyAwFlxSgMXt3tY4vw/cL+i3jduuGz1BSPAn3KQSWk6odQkJbX2MabW
lFaqtGRSSwBubm48gptRNytlvnx1FKCvcw+QzqEEzW7vTZM7vIfX7LAVOc6dsfwe
jrcwFCfLQl7R21u/6C1AKoDAckLWq+h5EIMqR0n+3rskqCAS6HKwgtA/fMpsS/gF
hLgI0qRyfgvmPGt70iF7Sln6mgQ36ak3QREj/bKiMH8+2AZ1CWYCpKNSPhWvXxy8
iWzbTzVF9JNf7ahwEGy1+WT+IK7zlWey9SiC2ZaydipeSMY9kuQxhgtJ7pTCyYGE
vMU74exQiBxaFpKihbDn8VA8rs4kitdebauKdPGmq8JFH5LRAwJ9J4d46Hv4e/iF
qSqevggchGkekm86oDhIouFxRWSX93q/sN4VsyPhki5L3sV9gVipMFeqGwwplnQS
LEA4v8kF/DhowJhmxHAb6E63Wye058CeF7wDinhw6Dhzl3KEHmy67wx9McmNqIfe
MZnCa8kAaPkLP57ESL7r4fk7fxgK23fEhXQE5kG+HwmtQQsY6atKrvYtfZmmaf82
a+IBc3NQ9k87PAlM0GMz+sSQ6ux5Fpg0Lki7hIo2peMzjEfsHDeOg1fEmSMHv2Od
99WlOt6sfKsCkrtnYFxf86yJymaMksWULTqj+P2j/mVvDJYeB9nrj0JdNWC9140S
xiLy/11lP6Dfq+o4g3c39pQQdOaNwPE0bcCuLbuckzy0LuR0gT3PXZEzlDhEJInc
6KFKAVD2RBlDaJTo3F8r60UWb0SGNhd6RAr/fBdW3K2+89npgsAb7ID7jeT3gAFh
Ob/USLx8uWfFGy4umEhQ+BV/0QAEu/XXJrQf46wW0XtYEE2isQj06JkbWfV+mcPX
7DYw1PrK6SGVAOGTmh43mSEp6bdG6mL2WR11hpf4zVyD35JHjMsU6P39wDPAPTbB
uJje1h5ypBKnyKOQLB9d86lP9O9RX+dDI0thlLgCfP3bTTw8SBfO1t0DC0EWNs1P
mvgHY+eC8MhvYuV8kUO/pUprLwthPQZNSB7dPoN93o3ByRz4+98/ejJ0MJmcUstE
+2uA5InsbRdK8WEnEpBOTI7zbciklpsMmZb6Jqvm05AueaDA9ASjb5XMkNTlGM5k
ByhhVq0D80SafzFd45m4c+R3VMwlFUiWFCnHgdEzEPbk5V4ZzjNoLOCgI0hbkRYb
DGOEeixyqdafG2JDnz3kgIg1KUoJBPEPXO3XW2Qi5WGjFYtcm31mgHXHTgrAvJ9T
aUn0HPV44tKTI1Mk0L8fShDO9oLfBJi/joNwZxWfdJlw+R5vzRJXwtHzE/LJd8QY
BuB/A6LpZCS5IXVAF8XADPbHG9z2desfSLHxvGbtWx68a3Gb5vGjHO3tfa/uDjiZ
Te5GSbdbqYuynjhJmKzsG9oasTIZxjgJhEZTE4mmAohP0AzVkHYtyz/S6NaHQUH9
rockBjyknGPM2138/1bF7ZvT26JQl3RABdLgzA+WmzVMsApXolRkKmryUTZCy/Jd
kJKq+bmTTJ9Zo7dZClPuEn0scKCDVw9xg1w61DcQdym+cR3ITNFIUH+2ABt7z904
r4MQNYg60P10yL0uzHFOI/MgbqDhvodlja0wcpvjg9TU2B+bHFg7mG2LgCj6sg5b
Z8p2zrJcirBao4K8U+bDQUuNuJYyltiM0fC0AMjxz0zzAIeGq1KYqlEcAsrRq0Ah
ILqVTQq4nj7g7GX7ErFnALnlqB69sL4tjfRJ4yiRi1hLQspOGsGBmNd3t/IZ2GU4
feTQh1b/NuzAHDMKtqfX+QezFQP+pwXZRCTL/zqJxvd7wHB7yauMiJWvk4JrZA8J
XKa2NJBH+JPlpH09xhGtRB9EKD4iTC1N/Fim+goHDrfqpWi3FlEKaLJFLgLLh4KA
vyeJZRIk1T6BK2dtEvT5lJg39XqQMpMfEvHEg/OWLJW2qz7hWa064Lc/L356Ie2c
+uCt+lswH1EhbFSIIY0iIe/KGk9/a2DxcX7luwXRb6OGhTd4H90oL3KF+PmfHfJx
VvIROI7khtgtvB5asi1WQ4LFKYoc92RrcbirHB7G7nmoWCvIskUHtgBjkpm3+Ekn
bXjanXTs2j9lY64/z5LELOfjZxXY0oArXBAhOiG6imdri6/Kol/oGeqeqS6eA84M
I1yX8I86T7A2D1Z+aq44TA91ZgPrkD5fm87RIAPf44Ye4hL0erHBXxHWb7mR059U
wtnTYoOLL9QUyUEZrPkc4jq4yBoQ2m3ouyBpnskTkmhtm5a4KeQ6REDv2zHAcw4m
f3YCrKsawS+DYrVqVtnGYYSXZTSoHEybk68rayG39un709zhHO383s3XlxctbxIO
6MA24o0yGw6D3Y1l2AJ4qYZqFXSRyHnCRoc9tgZorj4Q5Q/bhhqfrNvAxcNDePRB
8IAtlDFAafh82u/CI2sKU4TBVXGZdK+BWf406psY6TC2Vi2lksgttBPR9Frp2XZy
fRrIMe65/RTFwwP4dzxxjKrvpd9tHbEQZT2ySCdAvpxnL2WdpbuZOf7n1JuHRHNQ
V2TcKI0BTNziYHsK7nru4E5sPTH4y7kL2KuHpkS7SfvYOrQ663TL25tNGmQd7xey
dW4SF7Hi3nrxNhA4MCggBWKJnmpYlKQW9RdDrzVLrH2UCkZ0511Jz0FY0L09M3p9
ApV5rtY2DXz2P/BhiHswJK/50JgT/FYCAmrOBZhg/6c5q2yhNbhykYLoWinQeeI0
ITJpNBE3+IsFGzwyBrhHLjMxSrAXEEJKrwyuGtjuIBwXR35Gz8nMq0hXvKGsnLvg
8EBWstu6PBf7XNqBaGlu8hMGlxfpFZMx4s+pZZ2nYqgW/h/aCCtJg/Lhj6BG+8Me
pfutrUpTMhMIci2v4hsLY5i8vS5ve9YxDMR+HJ4rHjHvFOeVBB6OmHyCPYBOvDRy
UcJQPGdnKmN8r1hWSDInx9HVE0/ZuOc0rOWBqnpSXYXBpX2mrweN1A99P1Csd3aY
CJJ/ArwbBGwhXnLOOHuGB+RWZYULGfsG8ELxFo9mdYXhov9b1ac06RgF+JqAFbwE
drn9SybnmZgV2rlknEY5jSijUbk1LNkNZyEZ9EEa0FT03ogmPYmX/qY/vLzJrWLr
JAimL5wDTl8nhDsGb6385cRyOrdL7iQqiNj+pKpmdCDOJ17Uh1wAWt/eYoMfhKei
TqYtNf7oiFPd5pxTcRvdQE391ugEirtCgizQA17+n80qBTHMoX0bI+aPUQmdiFxx
jUxBNzcg6w42LI10o8nFTDfrI2UlVomcI+yJdyCE/7cJ7pO1ME6SR2pJ50CYO3lU
r7knlwMn1sJU+bV7pbVQof7Tfni+tyklaDijdQskXhtANafI2YQAMYGn/1QKHy20
4P43n72VafaOCZmwRj2HuKB9PjQ2hKtk6JWayEHdVk5F3FpdStKDHU7qCqLlWLGA
COLBn3hN9e/rOY1t5AZ6nxitxQD3EdTsGuJHyYATb3wRCotmoktNn/I52gnXzN3A
WjpRbYKjXDuJSSB2qzzB7F6jxD9/JddDrI9GIQV4i5eR04CK3u9TS4uX3CCUvISy
5tsQ3XOoP0CXjo1xZZYmRM67XWnNn2ucx2Vurw0ou/0KG1AN6M3aY1OyMpne1NKr
k0ND7Qh2gRNAI39djMsyVEQh7P3oY8iRgDCURDO3pO07ffzJIZs78SS6My0yUT6r
5ENdptyrYOvTVLLTtrPJVuaErGo1LASjklUMDoNQN/979ZN3gAc5hZdWPsNq0y1/
JqeMgrreWvBjafETqdE9CkCSMEnC900AiExPV6Eey9kCLSgnwSRLC0uyt4z6XgMX
GAC46BhkHqoMs8sTH9yRbtgX8kr0kJaFfKdTpE/r8LnCJvc5zKY7jByEpgg10oEc
8l7fyErEsO0zc2W4OzWp5Dm30kJP/ZjOZd3E7HDqztNcCCgfVLjxMvbQ3gNLWEgk
xWaqiBRE+mosRx/zJzmelG2KHurgbU/w/jJHUVDhTTQQofWdwJvnlQh42j/gltp9
QTfnSBXQh/bd52vdqLfsXBRoEW4pIcf4dVJU/zr7FVfdBcj3RSo4sDoyv9df2Vqi
kXtVOg6fgMhf2Uo2YO9WJqY6NjuihUu3P/0E05B+OV113A9rszO1rlbvR64LQw/1
3DNaoU/8niWWGe6xhXBQqYF6Ky/DD1kM7MAUewWBWnsXeH4YXQSUtq5lTBvBzY2w
6v4kq0A0k2gJueQ0FW3YNor+6UwT2HYiuAmvGtVWZ0n+8FScu3ldaD0eESrFW0AO
f3gfevPdqnncsKvn6tBsd87V/4kGvsTnAAgGxTBxoGByJ9QslJPlzC0MdMAKdvZ/
r6Sn76EpQTpFMcIU3uRTVDQ9M1nX2u8NfYFbztsJvRVAmvNjwyeFTzjFKHIogC6x
7EiAJuj7S/PiCLof3VZzSU+hHUTMgayFxPLRIYyGuSFe8WYL6BXb6OE7AzC3PWgH
kMxsPAjhnvsK/ZRKjPvFXKnLNFoHJDNlymv1LXCubu0YQPQplv6Nz5O2+Hj0U3Dq
RbZw+Dt8LSQp9K2zUfrj4OzJn8rIWXl61lkv0tjTDJCswasSnA1GG9eGC9dQMlQs
udyvhlWjeRwgfXeU2kb6TP1X3IFknhBY8RbzPVY2YFhrp6K2rINa4q69udhj32Sj
bj1mjVOaNwn+glpw/XXg2ovoE7E3X2zk2BMGkr2ER+r11SiNVxxiKdFa4yT7VT3w
nIjQOqWMVcoq74LUxGhghq1CK16bLvInCez2Ez2fEIE1z2SHZ1sMm3KTULOvI58V
t2qzgc4i0IWbOQOdknY3ka3FhIjtjR4VKmrt+exx5vQYZkrqTjIu0ZjpCTnOwsVG
6DIbBHRxAAJwYkTCgHf6Oza0RWBW8LBxJt/yoxy9JpMqQJX4wi4yXUbssv1WEUNz
duftoGE94IQYSurgaF1XZ//x/hB/LZVYUY72dD5WKLTud+51xXcTj2o4Gq3+MjfH
WC6C9y1joNVwuvkYbjuFHfvOXPB2m9y6teKD1YD38WnIXHvkaat0A837qh1sfJ1q
lNuMO4gi3EQdOFawqS4r7ymuQyjICaFc0z334iGUYJBtROkV7RafNUcHyyHX2Eem
BnKs22+jRJoHL1STGjYAsY+8MEFleM0WWelZiU8X7odMCu38bLz1mpdSVzbNxds7
w8F/EC+LOw2/JHdHfFTzqOfq2urrRzmKc8weojRV0NIEob4R0rM6XOE7QZH2i6B1
VAZRPkHvTCJtw8p3Z4JfUwzrCLAeQRl37zbmmBhbG9EPHLTXoMdOzp8cF2LtFEwK
qrhX5HyeWvMk5pkcUzN2Dr0kTS6tkqIC3AwtMj43Y+/lEqU4QtVCapK5POdn7TFF
f94CwNyLlyDAdaPh1gR81CSDijXfkC5k3LjOeNZ/tP/iRFSxWy2rOxx8PTwH6kpW
+bnrc25sjtFQwaNa9R1ihpvt494YA9gXZPPZoeFCkymKBXM8zFFT7hEBQ1k60ghM
I+4GiC4H+09rPv88FjmNldzXC0GpUPSw6W0MzevdZgMwr+K1sGdKOwxkXqKmS1+E
+35he1SBjJZ/1fVCiDEiU+q5G7PplE3LIBKvqC4sgttwSCrfOeky9v8b5/rn8r0s
vQjmL+SxdRKBNH4bo0+YxaTtjstSviQGKiyB6WhzGSOnrootLIhlWHNcFFozeR4g
lckX0Z/GjW3qP27JlbTjLs5nJNv9WBroyXOj8bNixDp7qT5OM9v3g9Nwags6J1vL
rzagH2Fz2k7xTRimRfqqdlUYFpEu6nLsJR5q0Wc5iFCTYP6hLc6G7BI1F+5m+ebN
RLRE0Yrqfq0x7S1W8Rin+V3LE1qVNhhYpq7IXWwe4SPaWmzP68k5GJ5v75isHYBO
UEQouX3MPCXxIU4DPLUwjS/wwwgdUd9zxpKDN7CMB2B0TTSrm8tbeVWGW+rEi9nO
wyAn30g2QWzXAQzk7ksz5sKi8Mt0XNlsKjho4nqfNcnFlNBYhXDPSScHstAL+LhI
ErqdZcIgXsvUwfuEvRJwOWM3pAUmV+/X6cDDdEMcLetahRWc+9435cu9VQFT3CLs
6JaLR9RikU+dgnHMBex3OwqRa9zUIOsdVKgBpqAAp7biJaA5uyDfBsVQMptJPQUM
+76FXpK1+jqmVBAQuaGj3n0nDUelPA9Y9d5TFJMSjzEO671oUet+CoSQnj98rZXE
QvBLdR50VHaEJxpusczfKHyINpTzR/CaFBAEtjEpedlB1gGvfujEmBnXmySHXxuT
ZIDCxJQ64L5oYA/NSqDy6KOAXNJ4Xx4qdcuyweEzO6A1LkullDXaZ/HWiFaQqDEQ
7fvn1y5QsANEcfViser6pi59K0c0ECk344qtbOHAUUsBcHQ3jih2Uia1uM4cj3wv
kZPr1bvKcW85hKT36hKzQiW6Lj5LSWWkkzzvdrt77cxWr/5zUuJRgqkBg5XFxJfI
sxb1JZXA3WkTNJFzuDR0UF2rOX/UnUowBu+eWDYV/ZFBJeq4GKnpzlQT6q8Jpe6h
6+cWZrdg4yb77oBqiiFaXZ2dntKSCS8ahtot38Kqeea6/i7QPNmGkinGQp649w/p
ehOT0qYC69l9Zj2zcF1lFmlFRuMILaiwpN/1TS/5+KOklt/lo24QLsK/y1Xz4fyY
d4U5+0j/cPD1Q4XqTrmkgjWvjtBHH0QjDN4pQkU0C2ujgLII6PJ/nB+SUuX+Det2
GKOdH6YDeGd8A6dIhf8BVCBhn84GOASRZqfOhqChCLH0nyAP0dI/f6bccdAkgFmW
wzok7/KALpDaWqWoyK7HmVN+CC3+dSq/5roOmwxe2Q60ev8odCGyCdOt0ggh8lJS
8Ig4Vt8kWzz3o6m/BBArEVLta73NYfdqmT+JFJ4pUU9dVmiMhBF3U56h2YY9nKiS
F196vktg9pn/n7eq54ygLbZaRihZnCASkLFPFOg92lvV7sYYU0rUPUWb6YKhGQGc
viTEcA6p81Gjg9RG0+PEQshntTdwxWA7YtxHqYWEH1iORNuFx3Hg2O/Pq7ALbtWe
Q3vem/um9Pz5YwBIx2tE60DvT3MiiYD8ytR8ODulszvOIQcik876PHdOgK4cckFN
yvujdvnaKFfxaK5bIXOZ3pwDEKUoTjlpNwrTasFJ8s586qnkwYVNK0Al4fKHkIoL
YmujDfL/Cs34JbrxB00Y0xScW+BYU5cCm7qZLo9EjzrssPlbFXY9hDxp5nnnRS46
kEtZgtMUhUwcbwuB0YFjkgYsflp1e0k+fX2gPhSoZQyOZuIQnmxU5fO/TNFxZUGt
S64/a9J6Q5nQEp9zJJO5Bo8Fw7AaLEdo5QaxObN0NA9wYdRrnO2xhwOE0yvIhEA8
ykaYHT2g053wFYeIS0k990RX5+yv5sxqxC/7HElw0ngK+qIIoCNgT7sU0uV7A3+z
E3D5/N1h5aJL8c5EAiqyogevM4v6wwXzBKiVEE0j0/WFwaBmDx/qtvHMtfHmBMrk
GDLGhanB146kumYze/REQElXw8o5YSBLj+qP4LQ/v2ILqmARMM70SrwBeP1plB9S
+6u4/zAfYB6qZpJJKpMbs2RDdh+ZzFy4Vz/T8njwRxpsRBdMFJ6FDy1/Sb1WuaTM
HfopejQYWEsJnpHPpNENc4+UQEeXokeiGGAs6oivMMPzdGfLVVdY8CcxoJoviSOm
iiN9SLghKN23sYn+ySDU1ZPV5TKWJ+ZRxixXsC9+iPh646dt+xL0mCz1kmL65X9t
sc2jzO1Ne6BZA6ndPoi0sWjaaGdlNzLY+FbvMeiv+2DN1agCByz/Ea3UrbF6qAdu
8Ig/yCm4MunnUYJcOXC+hQ7Z+UFfMKGHrREpdR4Gtqueru73vOTq9SlRR4JlK9TL
Et/6UOAHEs88Jl8AU+6xojy/yQ/7wiG9D4Cq1ayPAwqlpBia0FVvljCxX42wOmSp
uHtdLKRbblA0Dte+VKkPQNESXmxN1KH2LK1bmKYW94Hz+z9lUXiku/YDLkRXcP/Z
bU4a4yx3kP7CvnG13sbEHeKVrmTiviku8tCRUqz4qKrbhLDyndH7B8MPlkTezrOs
k4d64C8iABt3yGVwVwPvEMVK0esA6vDwmmcew1guFvBaf/XnMCjDVn93tsNNJdRE
EVKf/q+sCTpVhdqk9GI2Wby1We7lIg31PFue+kqlhizYdbztVbyAqSHE+UJNdflm
V73FTxB38llgP5YDI3mARTVcGNBqbtWnO62fGcJteuifb3YN6s37dhYYJ347U/Wz
RWCeBkjdC+4YZmvPwWUIIdeabhiGDquuKHGZWCW9ew0U9P7g4J+4AMGOWczcQaTy
iJNJyQXHBpWsdWnbXcV81wQfvNDbKekeDBh1yZL83e3FRotQrk6EtKpeZgzmBWSj
oBGNnsBTPfmvl0CO5FE86jvFPGjULQJJZk+g9Hn8A8XJ6oWdjBo4asQzDuiJ/wU9
KIN/iS8S7Vlh3uEUpHjvBJSHF6i7ri6SJBJrQX4ibuG2XYS46yGrv84dULGFgRv7
XxrJRrB0TEKbb7B/i0YN1i442mCF9ZyBDEK7h3QZKYN2PNn8YleVS0jr72JQzh/P
7XlUErefYCnjFF7nCSYjp+PVhzVJR0PDKteMMo5M/qmJ89J7J3Mp6YcWAFl2hqB8
LcXoISVmEsyUC2v7Jw9NsqibusoRrfBTMpBg/5WtFD8DIBhGOdYGzARG031QaXYJ
KBzYjXNC0xNMXLuh7T9u3+lwqWUJ24ohxizewFPrpzoU3HSBuMOqsORnFNWcWhtQ
wsth47x9epKfmYBnYpYy+eei/9PZTfrtyIZAnCSOkC3Q3Zo83vkOgfZXr2W53nbt
0S9GJh1/baaARskEfb+VRjhgR1yqqJSg/XLxw2FB7K7A1CVRMhnakulZ3KEo9JP6
09hk2ys8llrnjx59CVKrmt+O8mdvR5IshNGjmTPJHlvDBx+PasQfoOBTTP80a1b0
x5NUSiZq1imiLieWhorpihVSfRGD7kVxCIb1rU3v/r15rVl22j7zvXv/6VMOfwXw
O5R+NL5OpZ7WIcRxsNjFZHtUYKQFPobuE7PAyErwE3gaVTIZmWNswiRRsUPzfbbF
TfiURm6RQRe/wMwZscFHpZvC8KRkY90oIc/R2CRjkLaGafoqVkaHADe6x5etDwH7
2tPyrFeqYuF6bzaRF+vp3x3oOBZSD8EzoVfcQu8WAOKPTmDgvKcxzP8IXrp031tZ
zowcLXIfAubPggmL9YkZLaPQvQ0A/IM9BAJ9PC9ra3ufX9fa991pis0wAPuOuOoK
M81IOdlGJz2FMYoC9yex+6QI0o8rOezCr7oovrlr/1lAFxVCnp0iaXmHQpI4SrAl
61o4BmVTlvr5KUbGQq9LDvKwJdLFNkBM0J1oLIoxWSvPlJ0XS3t/YVjY2298pdsg
fe+TZCDY4G+6pyoPV6tPB0Kl7fKrJvFTAHFNuR9UNqJwT3QsY3Pl07cxloNDtA1y
1TQYm2/oRbfAw5NK/nMqMkrRE9v25+SF/UjyJAlFyfKcv+NWLIOhgfzVFNcMhhLU
FvY3Q2O6491NP1jnlF//Ixh90iCE5EJVrxmeK/8zUR5TAvaEQ7EiocGWpHI0VIuP
FfWzLPsGSaTK7deXCHRzpU7HFm87CfHW+z+TgvRROsH9VNNRLtzQ0QgzD8ZRXh5i
xA2y1H494Jd6CfkaJluVuUwlC0t8YrNsZNhwS7CQNEgYu0XsHr4v8+33UthQIO4t
YHaN8qM1wcBSJM2WDMl0eeYL/MtUCmhVl4teUVn26cB2Cizht/qcksrQ+WP84+bb
eK6bUZQ0rnV4AvyDE7p3mFGcDiUGdsOEkvmTveyFy/h59Ceb6QREqSWNUv/FG8J9
31wuM1P9GrwBJ6Kg8ewKqkEsdrxKKaskwIwNocu/6dk0sFTMZhkDYslfpBM5CbGS
4khSXjM2x6mytEAr/I4rkLKG1SC+HfGgn2qSy4tKEUo+vKAX52c0HlUepmF/L6KE
jDk73SrSx4e59u2vn3VJylZXKphEMhPypwYBHFbGAFhHTfCEO8K2ivHourWMKAsp
65ZFwnnWmjEVcRnA6jhFk+E2l/1YthbEtwNZDnpK649s8ExqkWL/7bvY6xJP2hUz
ccddnb/SqmANKifajlC6rCEArv5v0VLxZbvaqxxgBDQic6MFecl+SBx1FMjwDakc
E2BGQ8XNWNlYlwqkDPiTAb+gWE25UckxPmhaQm1uyt3o7sbxF0Zq19SX3zo1MGQ+
80GIPoBqbDXpOTqu3omSexAa0rEvTdaGQC8r6VkWatdrSq8j2lAKh4UL2qMYRALW
eVn6EXZTjnVsIUMIEOeZwbGfEMxPLXinrqsRTSy27uhOMNYJTo1LoiH/6Dc1NF3W
HFTQOUeMOS8bfZ3xkKVqg1BSmb9pWZmROh+UCRbwBg2Ipe2nqDsSGl30MO7qS4Sk
iessTGRWxWiKyLjz2TRNS0/IoeVWB7YEBCTIbfAO3UhVMWQDhIWgxe52or9pED2Z
NXSi737N7CZr7bloOdL2zvah7gqRLzfTNgKOpLCREpqyMmHfbyexvw6r56mViDLY
TLog7OzYvkdW6JrOffLGxESL0qsM4GGigmGIfVXu0Oj4FWbMj5I9FLHQKq4toEz8
uJlWaJeYmC8yCLnFsdebfIAqWro7k5iIbDvuOxz1xxcgC0RQS+8S1aznDbZ/n7RE
N4hnJvg+SF5Gfdz5f+STtfYor7wkI0f9PccTRE8ClebaZudHjJxAHCSvpJU1ZsZP
Oj4IcN9QLP4fx/bQnna9oGpHsqBKRVz8QORH7x548Nutc2XfuZ+TO3PVq3/nLOsG
gt74yNuoReJMQob0gvZp3sNvdlM3WVbd8C2pVMUFAmeLhHr4ODP7W77i0q6lpttd
Q1wD102YhQJ5C//ZmfL9fg8YWOFhsmYPg+7MZDEvbck+p6VgXkIu6UNzoZQ5ArBf
CoMO2u545jhRGUZvMQ5HUPAeSTZ0LpgCjap8v/4qER2Iz3T0uLj/z4zYojtrguD3
zbJG2dFsNZeALR3qFLIddNBwxG5BhJKL5InWNq4xsrIhHqAPF5WSbjsJ94ShG1IQ
nGGhzOzt4th0g//Q5ry7nuNSjxjQCMxX+Y0H0mW6AvKQydTnmXlcroRSuL5eh3Dn
e6sAGpUPfvx9z6nZxEOHhKHKNlUtsRs+ngVMKxy/IF6e+vUgJYTqDWFom5Jfj2LI
qEyTZZFgbxKl/s+Kdbec1rHOWGS3DCl/Wn+1n5in9Xqlsim5P3Gh8YDigOkQAR5z
Xd8/I1TEgf7oBWgeZvV4bcmqSnS5x7M2gdKaXvg2XIcxKpTZa6edXHZCzf04svhz
AiHiveUt1ft04O/nJ2l+Zlrz/t6MeydJHsZvB9HFfBKlLHgO2iOg9Ml/mlfC6HJB
DvbDktTScOPbqT/7Z7e6dRQiRZM4BKC7xQaKfOeRybtRciI5VdfV28vhJBRZCPkk
XgE96M64jmejqPk8jdtM70qoXwUbO/s1w7mfnZRF+IlQcddS8VXGV76VREKk+HxJ
OjFaA8pQj4Fl3YTQH80+Up7nbfzC0WEpZdKBC7mQrWzgiPty/eHFIJWyjVTByOKI
UMqxkyFkuWN6syVUDYgCwSFKFxCoPSflbq+ggXWItsHORxfCaaHFm9GOcOuVRVxv
D07EODqDexRBfUDxOYfMrfqPd50JkdX6DqL++QPwYbwbtchyCcgd+Ya/fok8Nmig
Ho4CHhCvw34DUYp8k5xHnEjP8qUzByeWAcEsridezjqXcQJ5Y94i5oKUnCQ/gtfQ
tfHpfwwvY2hX8FaLwVLaIdTgQO+l2N8w6wYOPfIhvI+na8kyp2S63g2oymUuOjLC
DXSkDODe5gu+VdFDBQMZMIUImXbuBCOip53a4AjFWANj6a7amtfKRIw8RLMcnzsB
ahZ7ILHoKLANeU7DZQW7/ELK9gsLhhONI6cMPBLGNj4t/ofgFCRxTVwzMqnKzPXG
CHh0yovKhnEz6clz6bOJwWR8fxeCdsHy4ha6FoK3Sy91FK5oq981F3iilSfDMwrO
dbntcF6lPiBoDhGSpOvov/b1NN/Lpol/gZD3uKXibKUHzcJBjhwkbwb8F4kqrRDw
NtMKhK8xEKArpEwYZzgRawHRfEH/TqUePuY6RsZuNdCtbvNC0GDfCjZ699J4xd1Q
oodx8Fg/yN1DsacpnKHQK2ixDWWAM3yaoIx7CeDOH8I8M2HA4MvIg9JELVcr4ZaK
O6FFFcVCpGyUFaY6IGMeUdfVys+8URgw+sl+4owRwYQLUs4omiK7qTDqpgCzfe5a
t5pg12eLl2pTNkSaBhbIREisayXi9yljAAnjXH32e4ZOaVaee+T+xjw90qbRhK+5
5LIAYYyqTGRajsR7vX7p/pDmq8JlfI3lKj6Pek4+zbK6dnFd8cQatNhAFK/i2ykk
SkCUJvhydr0cekgsLPZK9kI6ywhGW2/U20MGl1ueF2nLH9poIuDUCf5BwRuookP/
9SFDS8LGYNJzxcB9HU4fOVq2t1WA3cCQcWz+CXEXz3D3bkiXizoccbQuzV9uPKcx
DxxCq1s/A84N1Jt5Og6nJBXIv1s5HGkfs1dThpmb6tH0Klc5WdMrg7tKpomMTbUO
iqUgwtQ+9+jD+iHp0ZpZsnHjXj1qok1vjeySzrhkWN4B7Cdy6f2mr1UVIRZmSCYx
vF87dyHJcOWeguM0+ZnqFz+JD3JhGkvmjfDXavEmtmuiA4O64BQyeQhwSeeC89cG
wAf2K7C5cg9q7qg0RUI4MBH1PDFC+Juw3c9srmdr59suluHk+xZ2jp9TbW8yLj2w
A9pvS35IwNsXYP1G9A0SRWATQ1M5AFQrkOV/oOnYHvMriZEK6qYWRVmf4AGY3zF1
/YiPXJC6U3rtIpnXVXuGr8nHDbm7TBt0i2yJJMrql/yatIJWEZXCWHk3IBMrpYmL
zAAqI0JII/ere1NZ2CtIJXEl6slnATkQwTEd67jvWgD6KZ7unFeQaXbs1QXbtrQU
VVZx52eOLbdIJe4zHuNCrFX4mU2GJ2WEXeLHOos3j/adKRYyxpJGOun+GK3G6fnt
WX1MuLuA2C3cyYgwy9rgNPCnteA/NCUvsPs7vEcRQcmA21uHsoyYua1endyQxhn0
cuHQ441k3mKNmSH/kxsPcmQyvUFW9HfdRTFQ4teE8nA+r9f/lhMjCJO2dKpDF3jm
oznsZzE1hAhZ6k8I6kxSEVmd84kKNp6rCSJkB8yS458Vd6GEKhtv1byTKCwsPLhX
FsQo6jK6fhgpOW0E98ZSmBKixPygKtgewTF2FB4FKmhfzb6az2IqnB3kg3h8+kxG
RtfE8Qc0aH1IZGKg1KperhKh4BVaVmAGp8jfHg3UINGcnhVZ1eGqS4nRbXL3d8gH
5/sza1O3xi0p+gjXbjl7sTnNlOpaczNDByOnC4jRfNNquBjvYruB0WXMoGTtj0+s
k3eZ0qgKTmQO6ZR/bfP2eoHK9s4Su6b7Kh7yb+7/CllyKb861a/OVx2bOP0nC7Mk
zuZXEOGEEON4uXebFDwfs8qtoULjePGRSsSFlsn8DlKEy76rnHm+k2Pfc5V1+Sva
V3xxhOcrBcCmDxNCLQUMeDGOVb9Y5PSFQe4KL7v3VGG1DrY2eJTD0b6XJUv1HLtu
WgB2YPn5xSVQbQH8CXlSCSq19IzGaiHcgLEkYOhUHuhKW+BnZ3j1nzKVPa3puIZP
8fxR3LivSi1XoFN33D4+mhyJkjPRQt+dndvhAGltvRKO6WVlGhfPRjYhXR+Pnueo
kS0heNKToKMgRyXxx03C6IHhML9hHwnbKZB9AvYVNCX10KdXmaULFSDeA79ygY5W
t7EArPiUfmO9YPX4QW7GqQWeLit25xsh39mkhGRIPWTULuZkyuBcjr0H+d49grCJ
KhAOn0rI9/wVX6AgzyxFYbLPU8XWQyqmLa25yW+WtPWjNlggca4qI4eGh5g0hM+G
ALYh06TXnccOdLuy3D51YQjbghtRNw/FSN8iFIk07DZoPaOzJoQSKeq+aBrO/uQZ
fpDFR15c+cqSnU+LvxbQ7SITBP8PGbIRqvh72FQ9ns4nDRObv9geIDDf7UyVKd1R
iAvm7d9L5PCItfwvAGg0uyzZJxJ2NLWaZkKQxERei68517mqFBPcz6OzyQd7spZ0
Hm4LehrUizvv8o0Rv8X8jT7hD0lWlmsV7CZEo6T1mVXVf+c+FUxvswLNLNGt5Z7P
L3+idMXnHQzCLigf6O9POAqZ1y0ffREwnOPd6qA3b3cdDF4b9tcXIefCHsZAxyC0
hGVTVEVs1YnfGIo4j5qznWhZgi9PwWkZv+RUUs1NeLOG4li8TyKgJuMY/BGpfeyt
u/nPijuF/4gLkB3JoenCnMR1XPvAXwK6JvCEOwvOCoWvtdz9AoAnrLgvbd2H1968
CKN4HliyXVV0ilcJbLCMYGjOyunGga8s/Yx7t4vaPgPaKqVgAxb2EdJ7ZX5RaU9P
ODMxH9R6aMXPSxEsap3qs8Pypx5qdcadeVtKMUzHRgiPUCbFbj3Vdk6O8Wvrbbxu
QoYG7RjcpJgYCJ+lZQUYMagQ+I49xDzemzG+okhfslR4lGEXTry5MUFSKBe9DNnv
xNRFijE8gGWK4DmOIHGZs38afpSM+rmCT+joj8Rw85MQbyakCJKyoviLXj5PLuWT
0kM94v0lIo1v5kwqSpxcSm2nvq1NEzk9CdWPhqaZTzVQxHIu3JOhPedHG/xdQOJi
jJnQeo55vVfPGi6CxO6KJ0HePORe1C17x1W/7JNQLAQq+AAH4SUm4NMIADz+JDx1
/DbSxtZqgOXx+dUA5euJGFMXfcSu1/8R/9cSGp7GCHId6f4XVx2zdQMQyq3NEKU5
dEJ2N2qz5Pdu3Q+fLIy2dX/wjNs122cQRNgl6Hykcbv6/lkuCiXlyx3d7a4JhNc2
CUENM/yxmgMxr6vP9ZwP+XhCuw0p4575+Ft/JdYR+uWa8uuhMCD/4kbb2rhhiAwX
zbFJfxNXHUxtMmVqpJl09r7A0cfkPT/FSY+AstOgTaCvvUcESBsbm6eCWfzYkHfC
RyIgQjDdE5plpeVYaJKs8vssMNm3anAGIZkurif3/Ccpr8rQInopEsDVCA7ZlOtV
zk9Q8hLNUsUFsrMzra6ghOZWYokWPJsuMaU6q7NFqFrSeNZ2FZ3P40qudKsjROQJ
Qz1B19XGnq5A8dc31iGON8HSsvWa+INmVQ8zBvQsPxqph7h2VqrKSXZZ/dmcQ2k2
QQSaLCahXD7fu0yTcEGZ+6VedYbnNgGT1Z8dMw2avFMyFgpI0Hci478UvjWwCswa
TYT3SRAyKa6Hi5TkNTwuZrLBIm9PqRtZR+8hLd1TTk1mNI/NIu9nEzxZCO345IQ3
7Le/nBrdH+3wpvSu+FH57EoxbpJnSwxGYS1HmcIpZHveoIlUlspNIkHItGgG1JPY
Mk5qonWLhVHkYQJAAEsOgG7VJ9cqbSyD+Xof41S5wgn+pdCrY+csRe+RR9TIPWYX
ivSP/F1DEKTXzOTYALpTmcDF0mplS5ChSvDGhL+RZrMikOnAAlTYElqbhqoO7yPu
KwxsqE+vYaLfhZImdizXS6MZBz3Xey5gRM2pwi/lExApk8scof878ed0YLloUKnq
Nv4EtudXsNiUV7+kJs4RNl+fLjqXOIQUWpJ03Hfl1lN7tGaZtB4rjE9NtiaaxNFR
UrnMpupO9FML2BXkfteXDVcevZ0o0qWhauJNfxCofBTmr099/6NXFzzH1A5RWDCy
Q7QDKd2U+TQhSp/P+T+DySPzthTHA8kxZlwhWJF/CQee5jO3vr1wunEMXefpaVyH
/A9Ps2S5kSLZqGclXmnJFWWW8RZmwauxx7I802qyF39tIyuZbbOhzxFNes/wrtbf
Po2va8WotL9Kh5dj4tsdBlAXYaryf9gjfGv2DZyZwHANzK9zzG6jlH2c83Ub9htV
VkLskEb7+uuLK2kzrjn+El5tOqrMnqCsMPsx5f4+9oxz/hCILwKrS3txjgMNqSl7
KOtqLH895h7YqvXVJ30m/RBMrkv1ppcw93O1we6O64PQG4+HYpKKb3bTZhBYli1t
DEk6h5z6ys5Yi95RDwSpMi1PWHTQJumNaKM5mYK5dZA3zb2qSKnFM/MSE+kCZmIU
GD+AwWisYkCvt2DmXYdTzpU5W8CfjlDhLt6SdxeQwZv+J6f1MRl4gBqJym6/qNzc
RuF/74aZNfwo4Op/Kw5plcUL0OHuV3tvD+eyZgTSgIlxSk3wBVENxfjPRyI/C7DS
0unoyt/nq+0c9wXb8uYZ3KDPbJGKPiwYydsmvBya4w7fmlB9Ns+ZQlfEfyd0VIvi
4BRk1NCI8BPz58B5VNu0KI7aSA3b+OUFbIN95YDgmWKfuQWLPwaPffV2hdTMxCkO
fM2kw4FZqNd3R1D5RZh6/ngJflL6Sl48yC5nXTt3VePIwMGkwXwzVOTJ3dAlUxS+
mvg2R1srfvbmIdof2zpK5yEBVG0wiG9bioHvilqWSBc2Z0CIXrLnHL5x8i5A6oO4
T/V8dllAMGkwq1WzPx6mYgjNhtFkHZEyr1fTOQpckvfK+PvYQDAeyVgo2NVDFL8q
YiQtgG7YYJZxSKEQM4QBszwxlMrE7kzFhx/2n3rrH8NI6zXK0GWP/DGrQTbBknmu
snYR4br7PV6GZfttlVdzuVPDeZnWRUUzkMD4o59lCiThx4NPkrGmkTcu8XuSQNtX
Dk0R8uMqcTq9Qj1b+QcFknZ+1NYLz8dXB7yJ5PW0KUj4sUXrnriDygOqm+sLFlt4
BrZQKUHoratPsuSPdKkBNX1VqEGlAl5MDS4RQgs1Iss+OVD/Vd4ZZPZlz2QhSJm5
uUIRnKVsGzLp2dJMHsm/Tn1BYX8zbj3KC7aJywlk02LwRlFW2OmejpEFK2XNCbAp
RNMTvATeTejSr3CGnuHJOVIP6r08v9tLmdpV0qprmcheGRLnZ4PyMtt98mfr27U/
XaAfCdtkKpdVkCUoMXz6yVKV8NTzdcLXRYzM9lh/n/nEb3yl4SKPDx2+FWl9ZYCx
RfZO8zNiB6EzuiuwYYn1PsKBdhA6NB+mmMjzD0pUN5roZsTIxSkCg3pIOfObgft0
6KQ9NGVQ0c+Qjs4e+yenDznd98DaGDVBmL7cnSRELBesRKjwal4Os2ZhVejNraIG
H/bqYGZRAARyR6m+MlWkeV4wzo+CvHeN3vkW0lxJMHmPg1Kj12PkhpxWUlzywx0Y
I4c+uL8PZxu+g+iTNTPogQp0F5jq/zCyj+hrhME0ED5EYb+k3oCYfOsLHphp+izY
lEYfb++s9aWvz6BkYwiQx3a4htg+gLgA5YN1OzPuP/yAGbXAgxb3gV56m2R79bhY
Xrel4irO00r+wNJWVlzw52JHs3fNjfegjCzL/KsjjJMCEoY8WDyj0thbnFlE8IUO
4e8ANhCivBFTrGD64+1xgK3nzDUwZH3yR0zmdQY/ejlr8G1IcsTxEY8GPZVnp9KL
ERAGAlcLB+HptzHnMxTaWqb7o4Xmx5EHphO8WP3v/ByiAs9+73QfEUsHVq7nqEg8
v0zhM8pe7os2vT91OP7KQnTShBSlz4VAO3O/M5DbCzwOooZBXPMEDixQJnrFM4Yn
6X6ms+hQ6AbBi5EgX4xb+gef5YvAFKUpeMruGsFnaG/kyywUDKvRYoJ+QufcTLaz
FMN/5/OvpyaGz8PABDv0H7pmzSc+4FHu3jzX3jPZsYxK1ZCnU9KDp2kvgumYmOEw
aKWZUShzSgS+BH061YN/VGG6VQtfe80VTcv1ltoRbDHlbXSsFDVIagB9UzZq69gO
VqktNCQxNwhNeWcmCmvjW46ZcaAZ+I4kbCjIwef4PmirZW62k/ITH5zOo1UVp5bd
skUdSWduZh5giZ6SRMqiODBFtxgNT2XoLjMI+/VVr8dolf/ll6r+nBtaZzL71rBT
pn5FG5IW2Fnppi7hGGlPKOI7LcRTRcLIOCQmd+Jnu09SCEWIiJGhFu0B58W3cczv
9aVopNPh/s3DZoGaspjqVQF8nUUhvnjeQkIrwNuWrCbnG9dLuLegKEnN1m213PkA
38HYKulkQDZQ6HYxGDkZPjL8nskThNfi46w/iDDC4o+hMF5+uLKYh+hk9ytp6o6B
6j43L1Gri+9zakHcq0p2/ZpTyjR1h9ggG7WLXbU2md2Z6jwyMPUBj5DoFXH3fEno
F9J5wxyyAc1H+ovpVIlib4UdToLMN7hDrZNOvoXhwywqxxWXxdLzeSBOJBr9U6zq
NghKDyNDlTLIRtCKma1UCiAZIANe5rP+7SNqDtQ+97ow7q5HVGv2pAmtjvty4JtA
uHZgkFln+2V4m9Uh9LMRtBRst+9+UOcExfgY977G/ogMrLw0eh/nz5f1miyzQjUt
JcyRIm+dKoQMa+79mJGZjbLBXhqfHrzYxeEsEgoDGCE7nv3XfYAWSB1keJZNR985
LxEKqwk77C5y+IBROSXt7oKMDfN3FASUJxhiFuGB4NC4rKMKkFRwVpor4zWWNXiS
7PnLfrFM0Glu1vox4a/dYUbaHhJP8N+QN/ClANDw8tnZLJlg+7XLBH0tiP9MY9nw
6LIZQzuyoKdSNHTwA0puZ38pSDhfH9xO8CCDZ1HzCIW3nzgqlTXT81T3KiAOYnhj
lawKKT3ae85w1Jipv7uQ9cbQbz2+9pxhGEQcPhFe921sGpp3MYkuo8CkQuJ9+d5O
mPeTxrCNbvEkj6sT3f+mm3WZXLV5CVcHWmx3Q6+RXf+4rUAB8qgHWgufxLohfIet
WTrn+vpi+ellytXMc16eTfL4b8BIQKP5pQlQ4fylexEJPhK0y/mI0zITUVC61BSr
F9OC7oxYyHwhdeRjz9gXdfVpH8W2RhPUCM1F6bwLl74Q5rUc8ow+TGH6QqkkWUTa
cOFWN7WcKWH4u/U6RHBNNr/Ot5+HFokXXu4ziKJhhCJHw246MaYo/12Jb9iSybor
ofT2UB+BiVccqiuAb9RoY0tDctvfkCrBUFDsagrw+hK0jOeHg3v+UVk5aQylSiBP
vAF3M977YgavxgOg52m/2F0O1YJUGn28SQWUHDFKf5zw/uXsb1nxvQ+hSTgZGJ19
4eAoQek8M84K9mCjt0O1sgUuJ7NjTbhmvBf1PHQTPCazToEeQd+nbgoyuX76QvOT
dB4XRiPeViZ/xuzvYAGdh39WT8Cj/jb/Gfg2rTWwrlViPYWmQXB5X6ZH0GiAIVy+
ovVrYvMY4hloPestwow9eGhPy70wOOZ7RemlQPH6aC3zeuQ61n2XiV5c6fc4U/3r
9q9+A9yxxBZkUYgTowGF5N3a0nbizswU7wwhG7gYjciNrwDXIweIzxFFDnc5IQdc
RAiupW1STX9UEA8FeFuIwr7B0m/B+UJZTuU1HN7OdRGr33cWFqFCQIQFdDlhik5q
3hqot9tbNmGZRbDyfALQ4xbBiqoQzsy6ZGoFyM890wZ8fkNvApea6+cGxmMReN3F
w5JOBvVgoZk8hTdtScGFmN5cOtzmG1kERLwMfrGCpIB9r/zT3Rhzgzh22mlG5RmW
vpMzTqhSs55GA2BA28UhaqjJutUUoiyjIA99RMaXTPlwcFrsJguEe4raKrp+NpL5
rHNvIXYdjlTpfzo2GJRaHZll+QROMF3NL+yiTxfTc3klHj0l+40o7hx+40BQCDI1
SEN0qSdyAb6Ics7SpvOEgjAVS7JRvl3Edx3L1ALpIdokbvWgrujvGfuv7Njwiazm
LiSthgg8srz/8zfh1EFSyEgWC7Z7tfrV5ZVbXzEJ61ZYjf/fAEpryiBC/KFH/v24
puaTa/FBkLvkIWW1vZT3gWO9H2iTuW/Gxmjir2oh9Pr/lie6IyMCBuSPev6593Ho
SD1ln1WZxWaJfYem2WpXnxm0MPPmpUA6lUtoNJShxW91Y5aPQPmaiRVJe+2dAFpm
BrdMyPVbs4oR236cKsBvsdzEoKqp33sUddBfgHkVdP8eNUC0k06zPXTwbuUvLBf6
otGC2PVgYiL8S2C3y3/M3ZX0noXyQa8zNkResv4w45Xsu0GcwBs9nHqgz8wTNcO5
WTTREPJBDtqn2+jHcXHbpTH3wEowf2DaE0buzpbehCi/XjYu6VbvLDvZCIwNf/n0
QpoegFbgUOIfjxhwXdY0SGA9iELp+7WZJFyl5TNCawxuOCYc9/UC+vu/eLzYnvfw
5wVIzTWve7whIZAJ8UFccXAtlX+p9r1qF2YzYkwrsCok5VpSAY6Ai93/4ZvdhwCD
FggzRMIfEk50UdEwbCi+vo5t+6O+QfOkg6WNT0aDSeqtXZmmXZinZKdtTpGLZJ1q
YCSjlhcniOkoIwri68iINZxTCd2P5+u2yzHejFE4NwatONt1GmEnHHAjVzKMjIQX
pu2xdHQD7H0+tZzRb2roeGlT8cAo8qbipWBXmwePdtuYi2luXvJbhCLraX66uBo+
oMJ+nwZdrWciHe24rLJA/SKKp6HoxHJbJKelwJZswIlCf7CSKD4Eh4hgesznSyVv
Oj3aAsPzfsbA1OGi+vSrrE1l6ZJAlx+rVKb/Xz44bhvXtBTRrhZohzNKatU/QMu3
YIX1GTBOZ0ZOyFbB4Fl74B5gw7XthbMUQNV2/wZMH62FhW6mczNZSW7UcSvB7oCN
OdRUuLlgSQBj45q6RScz1yRDtxozXfjcOc/uHdaFUiLKLV+OOzLEZcPxVa4v1heb
Sk7E64GSJ1qlls11ZDXLJqVO3Q88xTRj7dK9kS+cT8EYD1TMAhYUVoPs24DT4cSN
wASkoPiHE3rtf4QFG37IQywZ56InzFFslFJbp+QvhY0qIq67uD2Y3T2GrCHwkN9S
bD+8mWqptNvj7FsLX/6Knsgi0cFfZwOXlpRhCaly9vwhaMoaXI9IVfVE73bgulLa
z5DeMuIQO1dVpmEr0JhaCDYA7aX6QI8XPwusmnXX4YQNn13h7E4xY2MzJDJ9TyNL
TT3wID/fzlk1CO9ujpqN7Cq6oMYnI3BxikFw9pv31Qxq2bDZZ4SMsjwDEN5tyX3r
IGo6wTYWJyT2C6gGveWMdIZFOJdQN7fCPrXO/vvSyqXix1ZBG5SsKL1YvphiriY/
CmLO1ftaLFC5UmELhrQMXIqrRU4h5+AREwZgZu+0bnpRlZETWQshSDkWRFIjDGJH
3UBx8Ay4Z7/ybsCamU8FW8M79aHUdikIliUcxQmyXE+jLEOL35BATSAHCXqaRymA
ZKmMoq5wCr/U6xHCUWc9lAGf56GEpZAP7WFAvmOPMUfteSZrE2hGAGCQk+380O/y
jE3C1pKD3MDNTuu0KJGzBvz585JF1n69zkl6oVPJUQnUqAWG6ddzp7sIntQEYJ7U
gj7h4PQTHU8zgl7meN3orqiQjfY1sRVqWsoroVq9mOGSjlSUT0JdSAykrf9Flhct
EbqqF5OwiyyIHRsoBOjx+SwxdcdurpOzgiO01Cje8OY5NPf03P+cIGFcWN9frA4W
quIFbaKxtZxAkd2IrdXN4g9QfhibJUkv1q9NzGMrrvB6Bk14kNY+F97Lw4t0Ape/
pWVAiCpfWQpGzknVV7koivNYwblr7fQAseIiG7I166jhngFhjInS7Exs6HWVDxuv
thRGoe4gjU2LE6YyGIj3EYhWw4HZMZy1LoW87859tjLm4OSPa2lxcm4/zYgnnj7h
/pkp+z+Mjv1b8ZXsGX0UU5FtxyHBENE10Z1yga9rHBXtPbRXaBYsqwkqJrhxrjfM
prqPLfUb/1jtFVoEB2k/9UT/m1rB0mEQW4Hb3OiX1W2yu68ghv7GHxzsRwjUYdq4
QbKooJiSJM2X8B9pZ2Q7kOCuX7ZtPobjPxTpibqsJ7Cnu2nMDvx/lxhFYz3s9X3F
skuyGO5ehuXpoVR1XVvFDaWVAojVlWSiOn/ieVR2T/G6eIFNqiDAU7GjrTy+9ipK
uyAacIwGb/aeZWuxuwZjbLArU6FVIXzD+E5CypQ3ZT22cHmxG6aR3uQlBGAM8A/C
wfC6cL1zp0scqAlJlVSeqKk+JymjiL+jUw1YI9OR8upJ+6sW+HG+SrnP39YPldzi
oIF5CNQvjuAYw4ougOWTSlbTkmU0K6Uw49Jm3RVTu0vLAlsTOYIC6vZe76zan1W5
HnlfmqW8M6RU67lmOzIqxvgd+WQbb/mAr8A2rrkfF/A0YSsqIaj1hU0mI3UK356j
p3uIgsRp7EHBpqKW9FDPqh35LYkaOasCcCvu7o6TncE0jBFj+ZTFqwIthbPfcORs
nnCClGy8vPwAJKtvDecfz/GvuEEByxqtMA7zHx7ZrOUBDAGagTJB29XTONIA5sm4
bVpFfEw53HEiwE5YSH617KWmuyzAzlV0Xclc00x3wmz5svkOh6hjniTTp+UnYtX6
7Q0FGo3ucO1NxaGKZY+bysqhWtAn1NMXpnRvaItLEJPQYxpeg9E44tt3O2I18mAF
F6lbHxdNbEH2GxA8J3vNbc0TYo2ETd3WIGEg6KHQNdF5ast+lBnxrudIG4XisEnV
YQ0t8OWNzqJ2H23GLXiLfsewNhilpH/+Po2mywvlZc1nHIxLOVBSNwHd0faJ74+f
KAM2mjmxlFonTVKg8XXiBDCiB3UMDaqW2oAoRYDycltt7KPBXmWJftc0SHmWeuIm
qtTnW0SbxrxYQVUanjJFYDmauA2hFZxg769GsuyLsViGbO4huOHI7DARy+1z4HYL
Vrpajdg3F768uHWfLWM96iykcNzA4se8s4c7gF5vsoAiQBhrGmaGwflgIOSoKwcK
9ufih1cBmGcRQ6uVkbsIs25CKRRbMtAxkO5q3uXQjHpg+D2h9XAm4r/5Yh2mgNKK
W90scwqwiTg1otbKjdM5XJAEJuUGUtDj2FJQ7D1JhhXxJeL5Yreyxfk4q5TmdnyX
pPYBiO5d7yf9hTqaFDxt0tiJleL/HdrDWWfckIGl3ZNODSvFUPb5tmQmwi+AzCmm
rZwxHHEg5qA8v2Is/3dckVejJmYD9wgteiMLdm4IdrWfJLgjI/5hQxEHt2dz++K9
9lFNQtyFu61/J7sI3HZ4hJQPM9nEKQfHEzQq6KI5b396iNt0oXh2ObP/aELYyIHZ
ulPqBbbMja5m/xU2WyIKzgdI6UlYLjBAB/I1h/lOx4GDshPrAr72HHB4Bg4y9wZz
x635hwUKGUn1Ag6gbPanydLyEacrlNw0IeJujuR9tc73qyW1WGDetmwYmMxY97C1
no6f8cvU3NwYvc6KyKwwdL9Y45doNT2af87aQS9z4S0qgGJa0o/tLYabC5ayFLyv
Ef4LGUBC6FlrcIzneT5zL5CPlcLDVFHT/HMp31l1hXYl9fl7yVZuMgvxuzkX0o7e
67tcff8ldeFBfEZht8xFN0+G+onKbwbswPIjA6GJ4HChfdXFjqIWEVmhXQ3/WbkS
BnVuZiGai1VdPOIAEdKvbSeCKFEFHdjrSlLzB+W1nmHcF3FF3moOixAbYYA4EoUF
KryHrfyKMZisMXEohGZVgO6oywCIO9mw6ReURJcbJZ74YTCjP5p/bt+ypAc366Tp
XBm8C31bqZibyb86N0JAh70PeWLTUHij3iwkWjJy+yxx9u/JZQcEEVsZrFdAiJaX
9Kga/Pa6ko6iwAoUmxbDmyw9zSLKbwqdYyUw2KeYwmIjKcDs23Oby2Y+jgVRUsV0
Pn2EpARi+8PSuwSF03tmYZmpdc7mR79sMklR5iPZlzHnR44xjv+sDn0zKWxyfb5O
abLtTj4lcUH4TfkFtYdScEPu4NWdSpB1JsIcw0FK8KNcbH0UbCoI84gjyky0WwzO
ho1+lXVDpo+031XD0zhC+bYS7BvBjNZPU4rMHQ3G3ThkbOk/Bkv3OvF8RDUeY1Bj
j20tQpexFWgVd9XPF+5hHPvxfZDywbQxOgylE0OjWTnAQ7Ljz7i13aH+a93QMGeM
v0aTitE6N/WYtqDyH8f7r4E2wzl1fIG4tnu9S42BqQNgfEGUKBm7j5pkJoSPeNYR
0lAqwvGhLoLMLAYr5EYI2/WGCxinKZVWADWIAqSZH/ovuM2A6BnTiZ0WgG6S670u
TDubyQ9X1KN6lKpjKcuGaYxeLK1A07ZFJRfPYY8VmOgpvVn9nxdc+Lh9ag/BmPxn
XCtM27g4JUN+JA7O7M65SfiJLkRyfSyxHfslFsDkMkJVNkCN39aCEH9m8AN2X1T7
c5SnV660YeH8g/DmZwmQKnqKf7rGWRkzXyxPtWjZkuuxsESC5eyX3cIi22fBnHBz
D4u1xnK01mDgAaTVC7pjnqdVHWR2sbzqiZy6rb7zTYhKy3GDmaiurdG57WA1Gii/
NMEisPCA5KSSATKwr1SB2UlPcqJyzffroBkknT8t5/ayRc484vlupb5HHMA326mA
T/mywhmlsaTiNqlHvpPxyHeWiJxTn3JOfuho18nQyCY7Mp08lKgQtE4JkKPq/2Wd
f7q54zFs+UqiQ26R+FrcGlG4hAOmmX9m3FJJvaqTLw+eukRiLf/zGANdK81VH7Bk
Pu4v4gvHgvHFo/JdPlCsJVmhFwYo0QiCCVFpG82UKlRBEopC72j3ElyazcyHgxNm
lGnrhdOBzDshO1BVwWi+GRCKGp9oPCtTGOPljpNzv/R7f9ANwZkNBbFiOqwwbvgs
Q01877dGWIS1dbBrSnDtsGRoxEW90J0Fg1PO/apMbeKWda4rhuMq6BSTRRSFZ9zr
L25X/t4PmldNI55c3C7N8W4XHWLxkP2UvfVWWG3cCi5AEgJBK1ltW8hSAC9I6a4C
9jRjAmGly3KKol4T+jf1/fMsYEuWN5St0UGtWw/b+JBRfsSsaQ2NGAWdFzuyfvje
u92cAmJQnbl/byi/lYvRMtM90cHl46nxJAVxxcs8rLxPMC7/xFICjysr72v2NepW
x5KnFU/Go9BK3A8OHrWRdoHd161GLLSb4lOcUp24WbVojTZLkVWMOypeVNs/yV5k
GigJPW2Iie5s6E07cidiD+7tbWXKTadJ0xb3o/AM6p+t7TAYJk22UEzf4cjsUp5Q
KgJ3YprMUkAorfyBB3awaXbu5xbIOnri52E7Q+ltq04gqjQ8WbdyST+eEqfJENK8
Ep7w2AwDdINf8x1ipxX149b7iNl/whkCID1akZHgECEJdfEXj6wACPju/VXSpGag
u6LoSqxFj9Wpd47D92hwk4DseryH/deatGboOKKIZY7qZl2L0FtAZjyexGIW8Ybj
jlvieEupK6V/TPuoZlaatRAP5m/oJ7X1c1RKScsSEggvby1CsiNdn3BA7TWOSBXj
vaPn9+6myZIX4zEG7yJcrel4sGjazhqxz4ox2ltpD7F2yGF+vK7/bM1mVDML9hVm
+YxOBDkYL8ie0gK/AfJadauvFHKEzVskWWoNvbhfl+xxYyrx/fD299oTLqJqWYcr
y8A+BaEnB6zmGuqv0ZZc8Vx5k49PlvYUWmWvtsvbQ398g3XB7VHWCtnCUVC6y2M1
33MAiJoPbrTyySoObEiUjO3fXCFLmQGrGFP9UJGCNCleyUQOkEyMplldFgUXQ9+m
4D4PDM3mBykv3qU4YbZVsk1XyLg21qq7zSWsMzWIRaASAct3oaG1gyVN67+aqXjH
hr9w0UPdnsPaMVLi7ydvLHNhyVW+ZoOM2gBufOFbKYIEH+cF9W2CeCsQiwLJxNlk
VX1Snh5vnMuRMbS0t/Lg6qYtx90Pc3SZ0IgYHnNOjokI5Ads7udY1wCpTG8Av2GT
V0zFf2DjolIYWL2IM/jexsJD4E0PcNdHjIh1CYjxzTgdXTu5+VQTUCYzvrAltULg
c83k2EHe1WdOjy8U1SxMvH6jJsKv/Hj07BYOHA79gK97lXfykhQacPFh+X1hmHVf
Smf5gXw7V0ZZqlkLPDwj+MDhvaHRyCDnpgSOr9hzoH+YE1nxREkcdkzkrdx3KmiK
dS7ngxy7sKMmDnTQI8qyoC8vzjzjeXHFvBZ3FQ0Eo96W+yHOBaTI0Cv+3LP7Ure2
i+VfdkzMvnEGYmyorhtvfO4P5SSuaoP2CBJXquB7Ax1dj7UW8WvRWeW3VPoBHHa9
Ge3un2EFWL5ZKvDfpvUlItNgRrhG9ZetOr3gOkkn1duke7GoXk2ckrrKLkTo2zWA
Y8UkiyFLgJt7lpCSlA/U9ey97Pt5OPR5iBrrLKI+rGbvbIaBOMxOaCQbW06liUzM
w7yPK3W5IQui8tIi7giVJ0JG2IG3abyY4EDpBbZZe3+zfiqPOJkzua0j0tuCTlEG
fkcwwglqkcQOV3GYEXaJhKoVK90K4w7Yeq8X/yzEJBic8X8Sk2OgEg4rJp1YHU7Q
uj4jbJvziDcqjYA2fv+asyjcy5aR1IiNbyl3MKAh22dlfQ/XKNuwRevybnO9LCp6
bEOljwDW3cw5tUZXYKldfHTYXgcGGrxWhs7JrygfiH6YqDMGJE9stMpwP7LlhiLc
BwI9xTv/LZL4FNDVAh/XmZfI20Og94rQ7PK+KdSq5N1KPBcqZW/hWBbnhFiMf1lq
PmMR5izsESXgEk9GkOoiNJfm0qsEp+VpXgVJXFFY0DlCxYBX+ntM9L8qzGVHZFHo
m85OjSM84idYzOI9CgIgvdCkmKIWG0HnEX1vn4b97evJQb/o+FUdCREczsUcL8U5
32hLRMl4wdT0jKU3qywRtLep3cDXaLNm9aEUYqqNc32uALg6vpGP3kIruK4ffWCG
54d3lYXQmdl0+u3/Hd+r9xKerBYuLn4BhV/coIrjZbX4cXPNlxeJI67peQB7ll0K
H/Tc2sMlPzPpls2/4UwTPq3MDOgtYbTcRr8CWLd+0NHoaQd3oFi3CEUA+xmZh17a
q9gaRe8+i07VUmCxBINw391VTsOBJWc2BkFbZ2gP1bVPVaajM0Am3lgaS9+KwqEh
VL705nSJrN+rtG+QXVBLbn0SV5aRyPQyp2st8ITXI+IfHUBX+/0Vs5hCICga/JcF
RrJiH5Z6gc+65+LEOHW6wmOk/0O2U/fI0UNx1j+Htb59zmyLe6sgoD/ujFRndOgq
URM5pAy5QNunLDoaaSwCNPBvaN3EuU9zIhDhttKE+pQiN543E+iH86nC8bnpuDNH
mNuL3+//v0wqDDnR3fzeFJtg3L96+/W0zdJ5zyfqfIvtydDH+iMlSJ23ZfYefa9j
owM5OGtDGFIsYmSu7GAZoLpyHd2VVQzT1QLVpqe5N24xdb7nuZA7vtI/Qn1XA+IY
URg+Sq8qVs2DDVSJMsGO7zpWB2b3gZ9rfWUC/pdBjC3RpENwja6+jk36iEUkkbRH
Y9dH8kXnxQtYJJrrqB9wVU/I171eEEjccxD8S98Wwrrtm+2LyE2OlRSvqMqBCb62
JsQEjt6BaN4w6poIyfN6wx9jIUbqrYDwi1/DEF0FP7Vv6UIVrP8ESYQIB6Auou7g
BvMxPFYrM3gKU/PiOd/dyREfUDihNft0M4UfD45NrleXyDUxaqADYZkc4cPSPS0B
AwsaF3q+j+9gDRseK9xVPzhJrgZe0RNUZkmolKo01zya1kUDDNJn4Q1lpGbFjCdZ
5tmqxeFvPdH4NGbY764aotCqtKhmXwMQJtg/gKWOZYzmiTySxtwXXxJ4zNLGI6+q
UroKYbPKzN5rTBIkNBNBrG+sjTw3vKEXzDPpG0eyQVGKoA8ns7RzqIOmql/O6CrC
Oy0Mq9cuLe2X0C8N3q7Xtzrsy/ABpZGYf7zoY0866K8uqcNTXrBMqF1Ecovk9Z0b
JOABHzEyWACaEHJAsV0RPSSGvaRm9fikzhTo+4D75B4/w/Kat3tID7Vjo78WFeR3
gb40CUYJCftjU5DGHykaSPAiFlMuQHSIBH2WZ2RAcpFalqYVuZ6smoQB44seujlY
iMUp9Nn7yFdoB7/cAcptw4bbp7G9idSiDRiYd5HL/+Xk+HaJa4u8ugYOdWtJArEx
HuqKGLO7gx5a6g4khOf9viAlfoKs6jVo5tbdmOMGrH0dSkGHCozwkrQ1dv8fnbT0
77SOfqDgKqzB8GGKMtIissKGNvv/Jf10S7UelE1Di7SJ2PQ5aEbTKwb4XJy+n5Oh
jdTj06JKE2+0TcLG5mak6teNZhjHJZMexX7IRjAfY/YwHZDSxhQY+oAQWCq7xbA7
C+HECi443qBuwTE0YCyXFWoPYUSNv1H4ADwoSy7XDOfH3nuIDfzkIbFtpENpkFW0
asmaux1RXCEZU4WA9IWExBnzdIyHYBKMMAQkx9LBvwrFSxfTfGjjwvcUJgJRF/0A
1lDImO2Yl+TCWEBFkrcKvS3rIuKLEx2xGVGWfYvvYYoWyOHVwx0fIZPclMSYbf99
Jz3ubk2HxIBuIenhfUCTuSK7LqVVcPuf3V0S5Dqg3NtRED9Ds5JqInvgEthpT0Io
4oXU8p0B1wsP4SHan212u7FET04yQy4Uu3Ic2JXpqJ4ITMGAjay6zv/oW8XCUVEv
0lLTqa6sZFA9WojaA20I3VPaLvmws8386zoSSgUubpG60s3TOkQKivEPLyJlzXm2
I4C/JeZffUdfTre53n+TYVa245jpXZ38UPPjMzZVp8Z+VMnmlny7CU4rmDnnS7uK
bNwiYUOc60P38TXT035LJS8ekQPtJlQeOnk04OglNt+JnEjdMf0C1E8SzaQORmnE
qpvXTdtK8ACZwcgFNWEHs6VFWxJiXqDnm8DJSMexML2UYLvDvH0YdxH/wWzrgoHD
vqQYMkn7wvPrjD6yiQ8GaoZNlaVNw5/RTkh4okkMlzW5hizzu6qE6Gw0YZEQwZ4R
xtq6XmrMiReyh4hLSRNcrInvIiod3aP8CZL96esb9v73KlEe8fB/mXZB3CPYo4AL
SHc/bU1fbLqlw4GBUr2Jscm1POYXFbe7fPT/Y4Z2ZuOLbh0LRqsJn5FZ75xSFl1j
J6zWa2E+QlqQ/Cpb4Mvo8k2UkE9EyMrs2CP2fbpg+IviOF9AbEmu6n7nYj0SE88J
YmhePvz805IBDVsov7J79gvSLx6kt2ATJTXeVVgP2ubRT4vk57roYg47Byraichr
SvbWGm6htfDzfMJf/iULN4f4dx/jJDp7Ivniofyj5kTYnHbX7dJ4Ac1j/a2BFDXx
YM5Rff+JF1/8HBl3wJIaI2bpYe3LOIWEvsa1BH+52u0rP+pwMgZiR9AWpx/FGL1u
PHhE6V3dhitzvv0e3Th0Kc1+7xNaEggZxxU06g1xQOK2Bk4DQBBWlm6w9EQarVeX
ggCrEmPnloWTqGEsB9IZKHvwS7uXUACPwvJHLX4O1G/6WWFwWN3NWGvRp1OYA843
ICKBEWyoyhMoHzg4uzv1ffLOR7mI/zDA+ZXfezHwbkjD2mIZzfRiFbzGrgM2sWCX
okkQB62Uty2r0zzV8hvN8RfVYEoK7JonTRk+dMdKWk76fxEw9lNE1PwCNFoRkbLb
ipGQwtyyNqrp9k0p+o1vZj71HLQjzd7PLz8OHUlFH5FoTjmuf2LTl7iJy+gSiD9X
M4ONaGnq/rSmhgii23+AYv/OmlyTzTBAUbpqDA806+TM8L7y7maQ61fstJXG0bDv
XKWPxd77lk7IEORXGvpS0PkP7rhSI7MhKLhCA0hpMJQ7F/kQf2FlQN2XW+Uaqg39
GbDkAxGhDbR7V/iMsDTTGN/1o5Phput8to4wGFtKCcQPHgdMhshyXZWGqLlTF1vH
OKxDVaOfqruowlSW8Nl3scmz2wAite3eI9kzmVWbOfPejkLRbtnNV2YBcZvt2Yes
K8pkeBcnSNjnCSXvduicwZu9kTqzGd7UBv6kxQVElM/qB2YtPGKpru1HVgQ7FXy+
Rh1AorVe6TFUeG/NpKsi7MUoGAEKCWbYTx2sOV+/Hwr0Z4qrqplNBT6NFtZYxUA9
+gHOeDRyGR6pD/klioKudYoT3k9Rav2D+U6APX9l3/17HPXXJLHj8SIDoSIUqH97
huY68KeROB4LLp5Q6pAbsJrVHF06JSlDjm9oEnBABXEj9NQb39c4QTKXxhAdpb9t
HvCl+rXATxusUnfL9d+jgFvj/9LYjrM3CmIw7XHXiCbuYI7zX3pfXz1GoZJIj1jM
g5OYkaPqAHZM5BkrJSRzyRlz4CBVhUiCEIa1m5XMqdlm+J3R/8XJH9KjUCM6xEpB
Mr+NibYDGrOuNjWl4YPvJ6FdlaJak7Kq9WQcQNx1bD45vWmeOeAFzJ8Er91UPvkc
s7X+jxCI06oKayHHfoAClZHXKrd7wCAyWryoGppCUkvMgi+bvDUGV8GpL3+N04I7
nUZcjXijR1Q5pbbasQb01/9uGHYwGfyUJ7HlpM5o7191xaO3GSjZ8npVlS/XUaXI
UEysiJUkpXfYPc4b7OvCdfbEMYbZjnq+jnvVWSNh1WXzv3vF1v1mp4iHUHsStIHj
Av7fhEEsvnm3QB/b5X3x8TbY184QPT/UFkDMcvqPjhXZcFZKdd4Bx69i/wEt9Yxv
E6obeevgQ20gsgYSTHgeV7IpmnRs72iaTMNiBhQg+yalnrj0Wbydj078WYUQ47Wy
6a5i5OKcJBpP5PNzMQJD6yUmHv3EwdB2hsc1MHjG8y4qOMPvIdGT68fKJgdRzier
H4vaHFEVVQZz8xVGdIHUGumtqTxYh644/iyHOu2wo4Y8JShF7iE8/wgngI0pyues
8k9GLwzcgnZQqztN4waURleQsdhtc5i6+SP/U+NBUUVzZllmdUnTO5f5MmRI21EB
zAUNt7CMK8dScWA+G7et5VpNPYOgUAi9b1Hf8U5kSZJ7GXjNJYKMmSXJ3M+4bUaY
DO6XTlgrF2/5pX9Cw+Yt+UmY8XtbJ/hL7J383gIPwQlAYz+wW6yJDKE+mZ+YS8k6
m32Upk7WrUCeKqXfS6cBAuKBgmCW9OmSQITNUB55o3BZ3FUyzZt8To87+JQnggna
L7olFCNwImUaq32pp3WCcyeQVePjMcBEnWVTAMD5+RBDSCDVQXVQZCeLXrNVt9e1
/Rl5BOoKx0M/Es9h8/gwcXzjELORCsdCCZDs7k/7IjQqRIgXITw1DrI7e2GoDWI2
ZARacjrZuQcsXkYmPZlrvzvkygTgEEM/38NyHB1ZzkkM8g6xqia9Dkqjcg6dkezr
5gPkZtHiC75M+6IW9rDXT/qtQvFUk8sHHPMXHLAsWfsQH8SHb7uQyzzqHJRqEFl4
5gUAUjSOta237FnDj3r5iaKZRvQTYbNPVaftIXSuv1AyiaTl2IznHB/Iyoipe4Mk
3Cn0TmNCi8DBgq+oKeJeKbgwWrCqykJzxVxjUbZKsmMHVfPn0DJe1Yhij6sGkL/Z
6zPJvSwgw3gK0tl7mL1npQyHAgFI2FchCdakogGbi3Kd5KgyT7cIxmdtl1UAkEPh
yjlEjSCRupYMOrA8Gc/YFrMHKNGxiggYxY+zV6f4Mk28fG46XkvDXnLknXAkNloz
vgREu+mEvdjDh+D2H+z/BjfXlixXoucXwF1T2fZ7zK3YgYV5ElM8cFqJm05ce63s
SdA4f4RMLVcszE3ODbkx8TLVtMvYz6gTVQCIoTOlrWaBNP+y6mdLSiu+D2N+knnC
EkNKHoF3q5fdG+ACm44tuYtHvi+EM1Bm/jvvARwjLmKBJFxRl74tD0ACccvbfz/2
oA5POjrcx+bTmd5mvc1Wj4aJ3Q8iE13YxBAqrNVlQ78jgm6GKlhX0+ymdeM6DWX9
AlEoNmIgbCZgV5aBa7Q9EhXhLDQuH2Y/rq5KPNEtP4Zw2gwSr5MlZSL4yZIxxoOK
B1qJimjM0SwnqzjQ5SQQNaFu9CuhXPY3TOESomVUBckF4GW8sclevglO+PsKmuNV
EzCh4HBevjvtDRdzqsVWydpzK9TEQUZdOzz5NKZMF193wtaddK8GK6dm4rVStvx2
Cvi2xcujnV/S3xFyGD2rtYj3K9aNr8MFiB0Qy31IZJpJy8WBkzSuatIVjxcihk4M
NdBROaKBVN49oZgtSm14MhqfabCcwr2mgR61ELJUJ7nXGCo2IZvvJaslic/uGw3t
S12YuL3tl3YPTTQj9EKUOGeVwPSsX9Ehf2RSYt4Ag7g6xxYmJvnVPjsdIjtd6Lca
DJ3YUovrr5tYuYip+Xy7DGEH4MAl5iRqMjK/LBfuzIH8QndiS4Og73kVISG53gFG
RaoOyxthambbRcz1BC8V0Z2ZtBiIAOzsI9EPmcam/m/q5ia5uDpYLRbzTi5iX79H
M4ChNu97fooaUaC6fNzKPNOTmDVEUC0Dd4KMJyIzAdjeySofnNLunvxnfGsaELsI
7TQn933/dwfLQ6VfS6B+lU2TkQ+2rSHnOxDDmb2y2Lqil4bqKnV0om0jqPmRXB0I
jT+qczhOXO2d4aA+1pQ2KLvS2bM1MfMCIFjoOfVpav0jXc3JfhTSmU5U6iWNMC7k
hlvjz/3veZoiFL/WtQGcP0E8ZyjwmveYmVeOWrUI3lr1r5wXVMNjUoQBYxsMmIsN
fJCFxa+lUv+i0xS85eSs/XYRX3rU2H9/APOe/rAAT7US14bCwkJZ8g0upXpy/tuw
HlVJ0PLhn2hWvItn6gOfbqXs3HMGJnNF57YUgWTEZNtBcuLOkAY1K/xb4T3/Zg8d
TklY3GTkBZn6Ibnkv5sWHynBd0hBgvG9h+QH270kYk/P0zL7+JcoGbpRC6zdx6C5
hsYomF9NOgP0O2j+a52UqJuqIbiJ2aOOYE5dLx5JtAZE3XUEOI2m2Re/KT6CutvK
HaFtLCa5qbUwCIjNBgfvOvH9qF7X6NchFUIEqvZ9awYLxq6fXFJqo3MKUvhW4Tpw
lfLn88Nsyv/lVGDQUhLNReePabMyz96VcCULwIB+AM7w7inV/BhRfKx0yg+XkjGL
eGXwToeEUbI0tGjeF46sbF8znis0Lp+IM/E9iVYHn6EddjZgruaEOBa/vgcKFwGB
1WMuysTDauHDBHKZOUAdujmRzvgnJzMo/UidtaUvn2zQ7E340TfjfYP+K4PH5xXA
xlzmECy+un1bwFpEdunEbvd7IOTSEbN8VQziKproLLdKHyARs80xbjjTSTQehby8
KaVNFHJvMYiAyVaO2IUrn9NvO1zABQS80JDMlIfdz6xkpPcePULdY7dYjUgWd7Qw
exKnM6kA/6pWVNes1o/8A86nTac3463yHnpINCEZDTTB2X+l/fqImOOm4VeKqjwV
j66vPJCpgriPw84jw+xoEsL/0XeXhki6CAAnIOVy59GFm78DjRdJjSG1nXGg/7rg
wOycQxT61klvBa81cnWtkh2D+scggcIp3m+dBNMwUhuVbaH5Y9piazmt8UTB2Mt6
u7kunvcum2mFU0FPVZbK1UIARJzuhx+0NBMnpaF8Dtu0yogpB/Ke+IkPaex8WRUy
+PCQa2/YKUBCekWoBLW6dv5VRQ2iSHhA/4fb1HYKDd+Z/NhRVvVHwaU1gVphWBpS
odeAJ0QSFFf1uWtt+HW7B8WD8HXPP7XjD15mjMdBaMuMUlWRWLMiPKevD3CA5Xr9
9xubw9zrFKzx0BjzkWOAEVafwkFawHUASOQVUYDXq381WxsOd+Vhj2UhxNAfxc9C
fun/5bpCY7JVw1bezZdv0eNO4BilQsfxYm91M9aG/rYg/nUA5pkiEAOKQb+EQZJd
+grp4AAWO9S/3r82BQ9umKM/yShZHxa5DfPj1juNOvqKn6KYokyprGdafxavlhIo
8fWMyXKQFzkNCwkeSXUl2KD9GlwUDKyp9kbI4KKu1nP3FbcdeMSrlIbDwSOEhiqJ
2thf/D/8TCq6r4C+JLJWXBdXTFW/GNqekj2trMVKMDnNJ6dfJsI9L+9k66YizfeJ
tQweZagh4N9sogdhpE9DDF+hhzawDvIbwAuQ8Kuzvd4cVn2OYBhrEu2cA49TwrcW
xvWbFPllC9e3/yD1WN4OsRv2iOBXO69iKaY2ECOLgUpODl7FZVuNpyn0asJFof4G
XeZgyRnNAjl1mCilY5omxc8IwEdJ3mMFEKaW/4tB8TKma5Q1i/whpR0/rhQot7ho
DjJ5B0W+f4SlKVSQGxmPmrNY48AA7G3aurkUqDWiIikOzdDfyy26JU/WfJlXr7uQ
2K2uG7m5yEFUNh5Y6jaxbvGra7nr5JkacI8GizbL4vgDi1ClxoN3nHYeXuieNJd3
B+pehZs2cYnXCDVhhqgrVaFn5TBAtSJ6AIkO1HNbarbTCyYvwf9UsavyWI4scJEj
uIOMzvqtM/2N1fJ6oLV2dOle5onClJTWrd73AyjlUEaniE8BK/qWA3trjz8LxFlP
9JY13kQWezra+C41nhCbbLnPmu5oT8ICtbvJDJGyisAX5UYQ8WKsy7wRmEyDabYC
mZ//Tk4jkfPVTYY73P2UdQGERU48TWeaEyh7CI3AiRiIxKxp6dEos3jsSiQJ/vxj
OUDsCd7ZBVlBkuss73/n1DxKQHRm00Ll7trbuM070K6s9kFymBIQ3rrp4DkjbvaR
QqthBcdrPfwGsVOPt3/9EdK3VrMy+H5H/kV11J3PSEjKju7P2wW/7y3YWWTk192u
Y17Zsowzo0Ib0FvYUtMmkW3Y0dBlFuzlU1BiGTWVftQbCQX3/OpZBM3+qKP2HC5Q
7ayPwSOC5aa4O0FAQjgbadlt2Xb/GHPdNulAXYc8T5aqfiJ2ZbhQZ98mTUraSjal
jnYSNfXqQIzENmNsbKvfT5sDKINIl/REYe/ZmLHwmoAQJ9oSQsjagRBF1QvuR2Z0
aXdqtTH2pbJwhKeXwMViGwEh+tjX4KLlRfSDSIBuyCfnmnvQVWC7zYDxTM0f0C/4
r41Puyq/+pRo09+CxE683MoTniIvEuafGw2RNelc5+Otly50OURIem6ZMUqHV1KS
b+2Ckc1i4pNaaS90kbpkbgKd2wEfs0BsIR8uTaLnwNlLyc87ZKoVo1J4wFRSXvgn
KwzSx98V2oYdJX4JQM8u5PIbXPtuIe7L82ULrIN2plcQFCwa21K9kdazM3Lxhv98
VejfRhXb/q/9+Qv3kQ/rAKYtnBfnhrTf4LDfwYXbJczbQQEi8q/vP4zri2aL3sRp
Im/wDaSb6jVgMROp08D+UKjJosrdIvEg/pXAbhsK+K66EbayDPThJF2vGeVPbH3l
N1BUZdLqZyjAd4FcUSKStbBlML9g7EJZOzA1/M/nJGdO6+mia6KKvnQE1a62bLpG
AbxTzQ7B2WYww0DGQiSr0kOBsrD1Fpp8BZ5VSipVyXZK2ikBtE4GROZZNTxO1F6P
GpBpdvzTcEWYguOt0ZNqntYnIEfSNvQEr8iLnSW8RxfUcEV1rOTx/o/WqwwQNmgX
AOhcwO9cU9C1OPguigvocgvlQk52AFpK99cCDNSQNS/L9KM42wB0e/lGUzGbVxlo
4EY9qcfehI9PqQst6OOhbUT/mYeTRqvGzodKqqkw40TvRoPJg/Qcip2AZagadNl6
VBEI5d48rxiSmO2teiSFOdfodiz+Kb5ukpRqHrYewlJOT/GQDdxZSy7w5ct5YySd
bzLTddoHnUI7VpAoPVvByn9qIeqftUsgGzPmyau50WpAu4c8AkORn+dOLBCZTrn0
ZPPNVOxUwhnTg7ci9UKn08jAVvH+iZq8F9HIjBtvZQYZzvaZaQaia0hYAWp2K/Pz
4MYxTfhWDYTbha8q03XO2dKtKJb5JF4y8JXftxPoGXCzuzjp1f6ulGLST0HCJmp9
O1/8rwPCEBykf5Soq7T0ImOaSCba7VC6tDa1kkP+Ca2jnJNmKgNlTZXy4jnn5FaW
DB8tXp/vuitYDK9jOY6YmILVPWOcPmzzLS+QvjENnoQvs09FbK/IkDvW4/KvScbc
0U3o7pUvuKnyOf5SX2ru1xVXOKrxHkOdgWDKhWB4gAkcfLkJF5ZbwN6LSDO81k/z
2MO2PH3PnB10aC/LPTwo5vpn0tgk2oOqCfY62ls6xKGdfOJ5wfNyiJgSzTLc9bxP
fEtoVBcVdKGgZdcpSviIL1GXrhz6qtt0VB95kL2gBzNjdg/L6FZVy01Z+xuC4xXe
1dZ9aapuA0HpTdkMLmzAIXJJyfCa6R1Ly0A0c2CQIMr4nRMqwNNfUDP5IZYIYElM
LCkh9SHmnZGVHqRCciEtHrs3f7X1CP5k2c2Vs6mwSZieh9yJzTSv2705IUcE5FeL
XFFy0Us2TkvjKBFKzMfgNgiJJQkc0rknmXDgV/2ezNl8n6FN0jX0dIANaYYNQl9J
xHvoONptooIKYQNPct0/07d3Wklcc4gTcjm7V/FbJu27xmkvM96P1JX35xV/X6FI
mAG07SaKEu0OwsxtMrWfYi6+iK8KM5FGk4AhosGK5Nb4nmmEhwoiMjjZ3A0MupfU
hj5VMyUDUFc+oc4WNgFo/MpQ/R32tHEGFEy6Xjjzpf7JSIB5Zth0UH95TMISFG3N
B7sreOOI/HMHb0R92RzEsXpv21Sd1+XEGtBhUrt33CsiRLZUA0HJbWtX1Pj6iuRo
3RjOm3ngTTkLvKH3lGFzPMdKe9kJwrBqk2R8tVlQliVmGHYYIu9elww3VtKxJnNE
Tq/n9y+wbcs7yB1Hj6+hQ4olJuMcMUw67HSAP/nljoTtyllncyBHj63Qm6atDwTA
mLu15sWtbPeSDcLx1GT3T3V5OG3VCpjVXxjhzBunxBPZPRAYU5iWYGeTHspTxSon
3AcR1zV13yZeUQ+YeUSoQASZFUKs1OUkCLw1ktVO+oK4WbN774IHJM7LPTV26QHF
t0GT/dkgkfCPTZfJwOecPNlQafZrzWpsJbs/bM3CWNosseVsNX7XkaPti+lhKEbe
+bgVgP7cKcsTGn5xNR2936IZEfQdnw83k53vvfCJSTBcQASNpsnk8O51lQSqBRjO
GmoF1PbZBDYHQ6EYFC3sl7agojlZhtiD1BR54l1a3X+rcxawoQcwa044p3QxDAcX
vWG0Hy4WdujZFwiyrvqcmWf8OGxN/5qmf3IqcpZV4SV20n6uPttP3HN7FytBPfOv
xTKBSHJF6M9uXUGt8KtCoIO+qLL364xb6g1b5raayPWaO0EYNjAxgb1PwTUGTq6r
0J/FM6lPIYrq7ZMDM3JSkww6FtD+kZoPjhsqoslkmb+hJjwxP0dIrMOokwMS/M7K
tHJcYholoEHExyA8VeGtgrI6oM6aWeSYI+NxV0qKclrTe5ZPDc/zs04DAOcEFn/w
BCaL7T3pNtj2o8qefkiac9bAw0L+YcL6aJa8UwmJOWGFuEWazK831KVHnDRg40QO
XjoKUz5WkWhLqW7kQbVwA0OOURLf2a2saYfxNTHW22/EIQ2fyXHPWvSFpec6Oj3r
TjJ3XW43jFszIeDR3T2J9VHXeBN+kzQ3sSFz1jZ7SEvY9WoRJ156JH6SbO2Mwdai
IAPjtQIygwbZHCNoSlrlZ05zRwGh2h1Z5h96cm3vVt6bk8fPH5navKmn9DEOSQn6
3P9bk7crsXOnd0JFlBT9XSa8LgZdRq1FZnko9pReMCMqOWdG3nfwCYHvPVKyiDRd
Sx17SZfdVxiie+C/lFAVD33NJicCncBY/PFWa3NqPIXIRi5uvE/U6bkbbXMW32Km
qQyU4tWEMOdOuCEPM4jLMjdSdOGPc/w5zyQ0+DZpoJgXR6IP2wv2+ytlUvcR28fo
WfypjU6f/dD0hZ6MB64YzOyfvWEY2wTgeGPn/HpNPG49Bl+EaRE6IT9V7DcBVumx
yjmKkEua7qifQI6B/AIIeOy5GcfV6MMVhDA60xJrW2gcEKTymfZcHysIKXeJimxw
hGsnNrCsOx7rRC8YSRi5Pafds0NxUP8ho4n1Y1NTiLUSbwzk0vc/2PiC4IUYXkFK
Sm0KB/TFGBrcqaXIDrzSvwTBywub87AityeYrXXPdft2u0+N+OlN8nwtAKEEiHl1
W0m5s8f5w0Roa4nX50W6RR3Or7Mz0WO9A8yJ43dIKWagl8sjKoX0jfxUlruc3rGE
KZ0Np6p39AzCqciuyFoO56aiw+DgGVMqICad6kQQEld5B0FpY0v2mTzYOv9J3o/s
7u4E48G8dxNjjBDggz97KxDB3M/lGbFAnsWUX90c1qCLQfLrkkPriEzX0Jgorrjq
097zw24c3b65HxvPSrxjb3sE8KZeXDqACrxYj7lNrMyrCpNuAgcS+8utErcb27OC
5ck1cIy5ULXZuqrnQadOjQBONDSDowijAvoAZ93N/NIPGUwMppD+K+3JKyXqx4oT
TWxSzqIG2Y1RjBxP8P4miIveXZt8Ziq89DeoAKWfoRrDDmhGWrlgZkPl8xTsNg5i
wrvfMfRhV7TVxWwAQg2aNKOjknl0zY3RTOy7gIDJqMq0eU51QBKvRFuHMqcMeKjk
TuZSloeUugkXw8+A4HWtEYHYHATPYVYGWM+byxoQ3/CGkY3CR+mtey87LY8YSIN9
/aSAOay9RF5OmuQp1nUd6rpxk9uHYCaDxmyNAn9euRXBtQS/PZ4mK9YbFbIOUbcL
PLVnkTLrEcwZpkTtFes+HJ198Bq3LLneSQ33oSaGdzwoZ3H3hBmn76F8NSB3PDKz
RRGFbdsfnoSct3X/J+MkXLCPB1NRNJTM4henNcNwf2S7IP+MhW+S+nvrzOu18ca7
Um+utBnmMYA3IKAsbm6pghDGGJ2LhOoJejfBHkzAqnmatLu2AlF/tgDvYFq2W+9m
jjd3Nxqhqdv1CWepRAXE2dJGX3zRCgfZVrcuTm/MzrB528C08I90IAGELJs73GtP
maBgH6wkFhlt9K+fmbcVXhFyQ1z1WbXBfKGQXATKOYYcOJVpTplNzoUuuO3vAAHg
Ns+t96wIMLvEM/HJSKnek6A6fyus189rAArAFfKaqQy1c4rRuH6+LJkNh1gIHKVO
OnBvIEG+A+FgpIwJsB8rIhRRMy/+tcVZizvnOAtNq4EtGcsaRnsGOEVsHVKDC3FH
o929YAwd14nQVH1+6Gi9lhv/+nXN86eWDQWRBASZYJqa1fyLezqCiuONmci8/Ges
l0R3n2qVxKJgk4qaagyOvbdsGx16QHBbXqHyN4K9zYfeinz5ScY5+rCD3VrDbo5H
H/Nn2XUD0oA2sMWuloI9gB1lIAAvjWSBr1U89sBdBZoIc/BIWEHg0SNhKIgti7nL
Jziwulqu7b8oN8Xxaah7R57C4XZ7p3DOozsEWRcUP6uItQXBB8M6W4LbqRJGxO0m
PffzHMh/8058dMLx4QLzDnuVPgEPlGBOwHtbdoAzNBoMfMh7t9bSSmbMq445TZcj
fUcxK5OSY4UyoeKjtqBZsQAz6A6PgCtJJgBQIqEcMREVpIPRj7rxM2qKldKIxHSJ
mVUnnObNYhwIvtxE77CjWS5itfB7tRkTaCOAObQtxjGOnAMprUNeLSocXK3HsyRk
624hheyWTp5aJtok08233YpEKYqHuJNkEw2C4Aurt4u4JEzbCslUPN/Dmb2DbtiA
ndR+Hh1rQUZEpLV7hzZr3IfoGlA+b2CE2wo2bTacb8fnhfylCdHD0CCeGHKNHXDz
bZbwkZRVCvL1suUpZ22lhKY626A4RQWV1LDa8axQqk26Cxb4Uj/PyrGLzy9NthhV
y2b5E88Gq0EijxhQFQwPbzmV+SdiztDd0xQLa5c7hVPvxa6YxCNjSbG5O+uzTcTw
mWaV/iJq+qdW39NP9i6Jdr5gXLs5Hol+JBRhutOR6a2GjBIlXa1kVd+NQJ7DzxkW
tSp77BqVVCZFha121wjjdvkramZQYquS3u/+lAry7EZfCADQe2sPWYaskAglArUV
1OXmREDWS9TEh87sfwP6NLGVMas6ZJb/huRwccXKAFg9K6AN/NLezus/3HqNfNwS
oihNqi18LJqgTdxPUjG8uPaexGh+3J/E+QSv9A9dgLwJTNR7wlaBMuWTBx6iqa5R
kIXga+HUE3wXyBNGVowBliJKyM8qGBDhJjkA+PbItZKQUJcdPscDiDIuOfWVMMhs
U7OExP/4q8lMbVhCBm2F3Ljikf4GCWn14m5LNBJghMSX5aV9qNjSHoBttnJMUGA3
Z3NSBseAh5xbTJL+q3/jhgB5vGIuAVThV/wTggsE/Z216OJ7VZLnuy6u7PmcoSKs
mss8lvCCxapW/Q6K4mFEqypHSTdC45ilhtL5XnjVmDAx8jjT0l6qEvajDW27cwN6
dyxHJYdQ6n8goa68H2rgwdiFLd2hHnwZKoXdI5EFUsEHwvBdDelH3D8iJuFTFhu1
QmFYK3m8R59roh6U0SaovAk4q/hQMnjHbfUKVHyEm77T7F8wQGM40x3hvJiRlYrn
aXuXrBZHwfZ8ATNuCM6+0iWqRQLLMpDSYzHjFovSbY4gDMNUIpDd+kM3cOjM8wnk
rNCbFzUsd1qqW1aB30qHoS4WIPdr8nkeoXxgd2L7S3bySQ+Vdm4lAiBSvBjVpKkK
ASjspRDnZNm8aJJLITdAhm5bRn7xFa2/FaXsGzOV/2td5hAsryemgYyGBrU4yVnP
hbvk1HxB72MT4KmDl5uSoQ6Ohc2r4/YNRiYRusryD7MQP2FInQ1pLVxYmJhw1uO+
dGJQgFmA64waw+varnaKhiOfnfAROGfOB1ccJ1VbDYTxmq/J7QiPYRpwqmjNF5Ih
EkiFzQSgPWQ6zjgr4PrAB72rzXyj02svgzgbMwsqb7KXdu1i/GfApIObf2QcOt8a
w2fFarSbJP6fUTHtXnfDezX0oRq/Odzw/v7uvg/xszi6hpj/bgO2dx1gkcvzLCbm
rfVlvS91tGu/fd4iaAS+4WEMjggATYJv6lGziJGvKUn4NlYPDVzMkbvu7UK6Hin0
MfT6tKnOuXRr5WDmSnoJyThG1ATPGH8tKX89xI6R8wiTTQN8mY+/ZfrbsEx7AaFe
2Kg7tr+RVarNE7Rx3uJeFtejAxfl4vZinF/JntsTWiN68ey0mSGHrFLjEud2UvJL
eaej5ZLBnaow+7GSXCtw0U7Uhoog7n2S5kYvORmSP0Dz62NxThvG6KJbIGKGbIng
0MWrKb9lnT5KAtv2ojp3qP6Oz8ZwDT/jXXf5DpKdPVzMa9usXLrwLPPplTl6FGrD
ikKXIAkdGLa7J9hV7mutCC1uE3GH8uejFh6uHAE3Jz0OIDiiJw6wRhd1nZ2mjcLS
Yn8ZyHPjAwj/NXxGr9d7ntG0Z25o1N0xHzfPUZIm7MZeMMMM1hjH0S0l9C8iogyT
PLUJKPdUbh/kv7GGYbJ8VtUV0VGBlseX4ZEkqs8EF1f7sB29y2bHjLS0HgMHPdTw
k7kK1G62HRYGzmuhfEiZ4eBuGc3ivc4q/gXotn6KoNCP1uStZakZeGcxwk1CmErt
ATMfnch6f3iBvBPm6h8yfXJWg1f5iWkhO0n7GsD+Y3hU5hBjZSakpq8dTuSlI1w8
vYsO/otUGFIeQ8xLXS/9FS1uXLnIAr9a6G33h502bPWRBfvPzlRzyfRAbOZBEpd5
2J4w/a3bK5CCz+0kMwSXy3UDmCRq0K3Z/cdN9S0UowiRsJCNeuagoGvARB4PWD2C
v1gYQiakBAZFOZ6CmJBonhVk/BYW3euMIivGGuM2RLe6KyYMVC8pjTvjzgQcX7KS
c/PVls0tW+e/QubNyojURHG3DWUh328VTFyjU/9zGNEk/hCgydAZe/YrHghbfkO7
pBDTWriv/Uq0HSYFs4hk5h3NeVIhKMPq1aKS/4ZhegAuso2LQbVNqEgI7jizBH5+
QjtyhRGAmaosY4/KntDAcI6ConaFIFcWZWju5bkRWd0Wjd4ngD8L8E5PoCsQwWOg
tZB1+Wv43JMIxkCKc3sOril/kqPvuvLYoTKX2XdJVlgSpFXKlw5XwGpPP6UQG7+Y
uTHRxmg1i0R8KaTzDyGMRKFq2I1v11Yx4RCHlggXZq5So1NqdqMFxYL1pQ0l83pO
EMkuaibFgWJe31gfoVx6E8bgC2rOXA2woowG3PRbMIQUn+bt7RRwexqWAhHptUfX
ncUzipcH4gpe1IxkQ4xxgDO9t5cmlzz4fAaq79xuylf2bToS8DJHfr1HK4JDMhdw
NI06pz0O8jMAw7jO7kHaC98ARmz6sr+UUQRrb8bCnuoNoHK2kkfdCofrcpTVanoi
wbO9aR/vI2rjlv1Korts/kngB1s+YnmMAPqbrEmgcaov74LP0UJ2hnkrmm6pbi8m
txrzTYDfeRk2AC6tGz0c9lvl5gdD6ROzj1CB3ZQ8P5g6MLbr1LR4e771mcH1Zg3v
PDukeOIQ5pqBcRbcZhRTN2KKHa5D62KM3Crz8lKlwjKQEfx1zdeP4VXF5slgHI95
Jc7d+vV/C54mjAXDD0tSv3orYN019vtqRuJb2TIgvS6DIo5/EdL1sW/uKXgtTdX8
qcL5AEFk+gvpPP9ljLgphIITsv0CueoTECsNRRFPKnQEr3DLRXck6R9A1udobeAO
QU6KhkVIT+14MbZFZ1K6ovjA3lv9leFlQztTv7EioJ1iEiolHXdxKJfpls3CWiUO
xL8nREAc1bv78o8YE+9/79Ggwgb65UzTCEvGRSOgvfHHnwKpEuh7RT+HnQBd4aVa
IfPqwzFTXhUQE6wKUhI3ep5qiPn11779f7ToLG94q2xvFhhbttEB3KJRgm0b+DLU
MWYiA5cvVKZZb8H8ORyNZer0EzCrPHRQ6N/gfQehnUz9GsSe8GEwlAGOPm2gyqfI
5Y+F+31S7roefNwsvC+2JbPUMrJBpldYZ+1fyBcuRVgRHDefwa2AP6wVDeS+CAMM
gCTKHWnk2gTsVWSx2A/80ODIGJ1fQX+pLIV7gTHEDH3ybqvWpyRqlETDyW+/Nepg
djC4bOqUiPLIhBrlX9BQe4zufNvo9YVADXV6h1+XuvO97UG2AuPaaqYYA+jw4FgT
9cZlfx7aO1k5ajiJdaGUDo98q4eHWdoiaDoILT87rfYFcm2a+wg0BhGab2RKRzGP
cbYTfVE2OIeA5ddoTArRZjZ6iPCYCgrY/YBLpP8E198Nh3HW9RoB7blNPtwND8H/
kH7XlVyX51bBqHzbYDl1sa3A/jzGHN1dtK7/FYxQQSRO1kOUGGj6/uR5ecHv8vyG
+TQhkd24PdSIRU4w72NphnebWOBpyweMUUypb2/PlZJVLM3brUrgfa+iv7NYalNA
JfdYdGxadoxdWaP9G4e4TuUfDxppnT+X+JcICavGBsC8vq88zaVa4CNxc59viDR8
zLPqOb1CiR1BCmUe/8pUVmHC/CWN5WYtuXGEUiGVmAcwUnYKVYl6e4JodQzuD50c
2c8Cb9Ltijo4HCJDQkTMwLiAvQlubnDjSW+omst/GET7JLCZpmxK1lKj254jEN1F
aObuT/3+cvGqqm/sDEfroQreiuf2wcLXkJzdkndSGSiQpxMUbTt82UyqIk2ZDnu9
Y7eMOIr/5MueYrK9QHbLI4Gl3P/2EUIXP9yQmYGSF3zj4sz9i7C2mjbm+SXlEbI4
TkYEmKWVl+MHpqlAKJwtcExnIJ0ptHLaTcHNblBN2fEbylzu6i/VDIPl8Yc9XKTS
ama0MKqeSQfDht1uzUxovTBpOOHoX/a0t9y6fV9FeopuZj5T+ro91p5+8nn9qPeC
sihu9mVuv8RyNXPMhiAkCCuB+fM8IsFHR2JgEYUHT95Izzs3P+me839agPVv9YrZ
k/sHYVjcqonRC8RoTh+5XtNJ9KY29kSMVb3MWE9cuPa/8GkAyJyB+nW6kYSry+vy
bmDw0you33n0svbUfgihmYyeWXIL8GtKmRqyI1jHZRFVYXMv97TUiUJWFE3rz3ym
DGSxmSCZEnQMCr0MrZJ6VEE26rQ7RkK8s4PVjV2fBc2ao/Pizu5oUFBmV9A3nSsP
Oww0HybiWzV/D07zoX0JB4/xFIcS0ZLfEfBMMpn5ewbyzD/MnKyV2Rm9xYRvNVvC
QOxH6I4dBGpkehkXmhiQP8/MyKfXj8IPMSBrBqBLrsplH0G4ngEIxbavOykQYyQF
1fx6jxE0VB2/9uaHkgEBf+W5rP3xHrZmYt0tbfA4mR6Id2iiIFLrbt5BpmbFmtKw
Fo65njykNQcHznTzc7E0vZGunpi2yilPQAuo7c2F02yjUU83p3P1J5pEo/BCZYap
FbENJ6Dea3sLLL0hixlEi0VkicxBxsJ2BwUHPCuLg9ZCSBTgZ/cOl4PPhU8X/aOS
cTlZ8N/WEXhV+FKWfY6I9TIoKoeUMtH6qDA1I+8kjNm2W5yo64Txlpq+J4sG7vYi
JN/+lhZNb/TLW3heaDiNmibNvKZ4dcfvcBmhLGoEl9TwjwZa9wAk9ym7IlMXwRZB
dvR0x4NyCUY+IqQ8MlSkYfxdDcRnvsYc7hMl+pgjLUVXKS0Z/8ZX0jYxkcsm2VWN
m2H67Wi0SMmyvdb2FNNj6XRUgYr6U87vteBTrzsplEO/oSOG6FhvNgBhD7MRL4Fs
Efih5Pk5xV1GiQKwy3wMeh988qBR1eSfKqEVDbhMySIHXygS3lfp4hi5r1W+j+1P
QbWQZKUSEUsjIcD/YJ7WOKKJiC1je0O8NRGwp2NXblFAcuYOOf8azj959xtyi70c
9iZbrXpRi4OdxEORI+spdLmYbseJ5ZlJo1mMbOBReMTM6z99S1aS+NLgbhIq2RHh
ljaNZ0x7Fhw6XC4esKxxlp87R26rqOT9uY0r0WZH2sjTC3a53OW9jxOpHHDfCFX1
RgY1vlLK5qGOm8aVC6I9UhmSiEk9VGg9D3B4n9LXLhXEMdQHy/Wpd/49NTfkuLrJ
08A0zV5OaDaG3/ktNpS6tEBTBfIc/O73vD4KGX+3zZKmSSuTvJ1cAmeMyufWYtPY
86JtlksntBhxRfnVRlVWZnpDOIdoabA9ZcO21g6+VbMnQJEf22cux902In2+EREg
AykvAorw6Stzf+hxVyhEfwgYnUvSEElZmDdxcLbHjH9HkTC/SlOr70yxbFt0cjYo
c7sGcVR/5EcX54g5Ils5uW+gOXZhafWnmQ6fyUpbBqe9wChnsmizllUMJGu5uvpr
nK2fmcDTSwmR8d28WqwFOHLG4rQ19kYGc3awae0VAZVTpicJMjhiIojjyGWdAgRL
s4L5jyC8ORm2wB+inHhQtnEC9s4mAAc/0SYBmf4nJILC9eXSgnORNdyRucHTMXwU
Cpu3PFR+ejq19uODeriOWrl9a5td/FrV0W/b3zQxkiMAFT2KvLoUzFVL9KFsyize
tCo6+aNhBRNUlasyEfc056SqzxjVDQyo/lujEGiJaWM3gh0VXSGm0VdF9nhWt0uy
JR/wKaz8hs+Wm8Ct7ff933ySmsFVpSpc+OlVvKEqTifq8XkcfEPFvjNM4CD2ryDf
yUumT+fAYNrePI40lhSvvvK2joTDI+aFP5nfWLD5VPi8P2OLdZkrTFg49SKkHXVr
TUj5/VxMNCFJZoucv0cqcm8PUQHqx5cXhon03fwC6Kpw5cf8O1mfct4VAljyKlSr
CNa5Rn/vkMmUTf60F2VGKh7HaBtI2deUbZOPXGuJzydxL8QEAzmulF2SYoi7/B3j
5iCMU7zTnpxoU0IGcfw4+UHa1ZWnFT64BhWZNThmOYJfnBqvJSqNYNlKoMElNKSm
CmTr1hOBtn+W6qTRFgvAngzHafKz423CCd/+rHOHg2+G0/vUfisNK6lJyVkXU8xq
Z0DlEba2fJmywxlSbNluRwt1s93HoEE6c7Yp40/6uDUrpT2NnwTo45TSfn0MduZA
p/fPJpcq4q0m+IDP4332JRA1IUANJzjVfiFdJeFtf95B4fvqNZdo593OyLvyTw3H
bFsao0vDaFXrzxItOKsT1sTmM12LhYXEfwOcDoBaV7W99/nmyOGL7VIo87CoaVUr
ZtY1MGip0TOZ+oKKGFKbfbzX4LxBQgqraD+reFigDdvGc/oKQdwy8AaZpIvo8jNX
kOZD/fP3OEOvuQ1VPd1E7oDB69A4VaeFEs+EKiwDw0YNz/rz6Kf1y7rKvSI7Qt2n
X1N0zHLxCFlt5hIqt+YMegK6l7AQR17N4kMQxG3q1vuXEzrUx9qFHvm3iAEWK4OY
d1V2r+S+BlYc0J7npN/AVrq91V8eCW4gRGJYmFBMKfmQK02du9LYL0sjJUeXhZLb
yUnwLlIFyrAjUeB3odFZC9PENlQSlGVtGzSzQJlzyoG+2OZru3o4IaYb3jqoDKcd
VWSBGnJrMtyHCyyBx8bWxaMtPwyCQWRBdrNsyK5DIfvbyttB4FXWCMKzN3eQDZ9j
m2rOrZgG3NVfeCKrhIP2oMJLjYVxMOzjx0USBYDOBjFq4czjFVZM+5myGJx4mCTh
hsDDUMb/aDN+BaKxZL3OXppT3me2p869TERuxwF9+Z6J8k/RrZGzHT2ymPblvm4I
yF8MBaIJMUbZ+MQuPBWoS+VI2u6DggA1kws0o9mMHKOimyymFKd3QtWAO3koAZCX
4vcmzvFJt5yEpUGqB2qH0gyOyDnOuMyJzIemiSMgpw8Fa6mCrzLu+XlTMZ18slO+
JiL+6jk2xN4qqa/MHSJJVqx0JWaVXJOmVlUPpi3JKA+dOYHEXYhOC3oBAlXyhqAS
JJF4Addl2Fd8M0LJzn24ZiXOEa3l4rN5/cx/NBiZ6uJ72eFT/6w7hhFxjLn1VKnK
FwhOgTA3VNrbVgv2mVTGlgRm3flJQ/WXIdiVl5RuFajz2zZJfZyJiy+U9uv4bIqT
6aUKuPYEDHugl/D2okaLmN8/IjQSFzB3ZcsD3O5EuEkb+ngDv9CUsUCYr2h+ZYAb
V8SoMQhbPS/kLMmmNls/uCMMIhcQxwRLLsekQyJQc7gJzTNgEYBidm5DOao5rhji
4oApuWMRBlfvbC0IwbILK5+rGhTIwvZvSnfOuJMgpIz07/bPFdxP8TXYqMzrGqt0
Lep0ldDyd6ieb5vNvv/CgH6aCQvn0Y2bfJY0KxNv0FUPU+pnu3FtVieIEywSMomH
ImJRtZWnu/kKfIKYgqmxd18FfBruo36DC5UM9pF6ar1UDfY2dCL636lwQXzoMmva
CyeysSzLqnWmmlykdAZTZYTJKVhkK4U8nVe0So9vmSu1lWIVciw9gEXIBjLbhjmB
PqT/BCvt2Ll8K89NbJekULtgl9SjG6cgcvuxsMCyhzfDvNTQki43ivb/PYi1KVdo
AwUuKVU4CSAaezKimRclOhB+4UOtZnUyhT+EKrs+ZyJryLqVE3RyXwCGy5MVEIjG
aA+aNt+bXYiauUkJHkA5N9lHdOuJfsP/XkR34ZBe5Lsshiedbm1Rt7IxX0MGobsF
41tIdsfgLC85MnUUs5Z35BALkN74qSSVctqC/ah3oceDOJpVlEbUWr4PrjC8hB8W
WqT+Oa6w+ONs7Fy7G9nbkCdOiT9sXDoz41hQZ38s/Bjr9bKDKqC4vn82cjrdglAT
UYPxnJEbS5LDHvbztn8RgAiASEl0qpMCGaDwpuzSJVD+CWWcJmegIzTq5SiK+r2+
eWFtZO73cBdWXKwQvu/MZphZNhTrF5X+nkkFVAnB7XNllYUHg7IbdEyyrXwSg1gk
CqFY6u25Mcv5y+CEr2CTeg9f1TrvFngXO9y1ZbfxApFWLpz6g5o95q3Zq/6g41p0
rzLPlB9V6kjVTqimWWacShf3h5W0iAv121OqomOOMRZ8tEkvJMdoP0Dhwwb3gdiE
VRbJy6RX9Lgt2Xky+u3xqoL4tpVdGUj0c6LAYKuCol7sFhRMKh0yfueZsKgeAdMS
eog3LmeG/e6c3B3LEgCpZfWwnWC5OEw70M0njs5JrcTlJMxwgTKSYBqFq7rqbpRw
OZZ9W+IMUsKyh9nIPE0N1xArcrbbiVvPvNstAXZxtn2kalZN9rQE9Se9UCiVcxOS
jSMCrxnKh0oS8S1Icrt+IUblUqemGFXtnQboT2/AqSKaz0weG7ufQxs6uRldsT48
qRXfAks2NBw22gTpweR1ugL8uzqbWfL8P457D5IKVjj4sqY2jqTMTmd++07pYiVU
/jsf0fD+vFIjNMk8ZPRu+6ydwrBRnx+g8k5Ky62Udpir+yJjvctk6BXm7S6z0Gs7
4s6bvAKGKb15KRUuseatZlLqfcv0h+mF6BxLPtQYk45HbuGnw1wOaFUdOMba7WRc
OuCImyx4Wnckgn2Ba4VRgy2NLTI0zWLOESl8O1XcPllUXQJZ/y0ScB8Wafa83eh2
6R0QOfPqhhaao8YTnbp2TzFkvR0j+EGaOQPyEMrzAgCZPnxAXF73OHslw8WcImGQ
xlfLM91pNlQOKdBdQGhCQpR4qGXCzQ1qfgD6ob1eagd717uIw4lC0YeysoB6eDgn
comj4K0P9Unm4Hv6lg97hjE2g5jG5RbMt4FFDY9Oz1t9zWISEDNMgyKy7wfhWaH3
C3eHrMdVPGFo0xrtWoEUovEwudULTpx2lj28FlSnTgEcjCPzE+c4ZdQzc6/KCk7C
0T2hjdfWHRf1jsymmSHa/hV/DBDwQmvDUvcKLWcy3EnDs5hMHMvw3usZPAy+byoq
WfqkYQM73kx/ee04YRoBu+iReKNwHjip52zrpHLuX8QzewWKZ6RNhhSNkx0pShPu
1B8W6fycMZnwF1NwTiFA8MSL/iRUwJQOIIf7ViVe6ptrcZ7+OwphHMRKuIxsjSAk
eOSfnftW6GZ7Zmv7FsPbUUIq6fJyB8hNi3b9/D2RSsU1AJBTAYcIg1p/n4eIymyV
YOrMiGbQOfpuTbcq2GUTu/bihlcxH0CGbQ1Odx8TgMrD5szn4fqzxyBH0bHD3/MF
bjac6ST6bjDdxfQ56f3bZB/cc1dmcxmAxfA0RFwxgbuSCg2lc+ahqsQAKk+6ZveM
4QfZkM1FwrnqyO+DEzhf9PCIicWap/R6mXjbYlLdhtKP9rD+kNPnpJpOluojYw0K
dCP4+oX58sPmgvVkukFXwbk2xUQvqC3q1Aov82AYrBWcsJrWg2gul8uVBjIVi3eG
j29v8HcYvNnOWiIMHQPISkBw/IjMpaP/YzFVKfSsL4T6DsnXymbj3pWebdE/mQ7a
/7QbOzG7UCm+PyT9qZxCuEaqv50peH4n0epNaeyil5wwQqWBwN/sYrQPfsI6B4K7
2Yxk0sax2jKKvYKO5y8eQw4DE1633osXXAQYNHKlQLe4/mxmC8c5zXZlGXaMQCMs
g2n9ksKB+Zg+I6bo6TLfsa8TKD70E6AsSug/qJe8ANB2UDdPGQCeeiQ8bydagUrD
p597yTUcWcAssXU4h8FIxEGxjqx9i5FAJQftVnzC8psNXHEbhczxT8sviI2sNhMe
e06F465R5zrHQ8OTY8/HdVmRsajdcw7M96fmOv8ztEY9Fy9ThwIn/AbGatD84kup
iZfGzqSAIJbHEXLKgNbBofLP/gTwKTKZA2NVR0MKMLC6J7xhbULtDANsazy8xj4n
aq8YvWJ9tW93nKCZbWKBhVi7ryWVhpw8nbmf3cxvTAtdI2wf8tpKTknI7lkW50GH
Ewgl9q20LsAiVTAk5qX1bdrTYbcjrA3zSMObJQ3XSLWISNmqL1iF/6lovoXkyTP7
FnzYIKtc+iXYwD//uFSJVlZ6rfG0yBUnL0ZnRax69JD3EDHIQ+Q0Fq+C97p8SKu5
BfG9jQrXqAbykjU25tQNazC1JYmoVbXkzNGnZJRLyI9HkDjNYKgGoCr39mXw9NoA
1wUU3FUkZZAcLPPsVkCuo79QNynRULEGgeZIeYApbTjuXq2MWyj8torg/WdbSNcF
lF8//ZY0hNl0VCzkplkt+rmu54AhmtI2Z9CmV9OHGGOdfNb3YnQPmtjjwGGowuMH
X5Uo6OIEfNxRiVg4vZuCLEID9OTXqBaEQOesK57/vNzDMIZzI1gEfK0a1bDBBvev
zmFhh6E8JEXPhsALy3FwvfmmDhqwejm9/B/h/kZG6mH3w67p1FlwoJmD1yuweqQY
rc8Ig9f5ACWmVXtLP9/oFxm8zAKqTwIJHdXTSQROb41x79132oHSeT7xE+pZeHf6
Ah+//l0mSfpjuz9AMFm/T/acKTcmt47GplyB4wV5AvP9uTmJPzP4GXe/7JPLWgRh
ScljJaO/uh6Q5rZ3nx/hR0s5uaXFqdHAFW0ldy403375PSrd7vfCMojHllEXdiRH
T8xkV6eUQNMputSRRt06wEy6U1Ct+zRqVUX5ACfYAMAStjYukNVRXnRn2Mor8019
WZ6yuP0zHLNzBzrKBOJjtUJLAYvNeBlWgiSWFqZxVHC7XX4lPKAMg86LlxcC9K5r
+gK8Jpd3R4Rw6TdDBwWraqibsI2OL1xO7C5yCD8jTUmIV/EC6JYLm4Jf7ly8AIwA
/L+Bqek+gHpn5OwHlfFiz5dsu+anIv0MpTd33DBR+j8K7ksYqOLwvBi3FFSKoq2V
2hITA4g+YK2elhDbzQlNrQH9GRRUhfsS4/WcuEHXzMv7HMUe16C1jV3z4qCwtP/L
g4lOe/qHgmCBRJVsiUrKLIP9SXGV1MGJUhpgytjaebJmSodDOjwb8iUPqFMBodMt
dyneL7fN6n5RNPh3NLipYZ8FuDg/ebSZaCf4K5L+v+ecuYHPIRXh2TJdDFrIYYwN
PgzkKaG7U7sOp4eeR7gwWiKn/GgBuvyK0DMz/VSTFMiYJI4eXfZfazA0i8+JZUjV
Ql5YG/RAPyqi+fj0cegw3cnXvEMGB8m7uHdbJ5jnyC1zP0fOpthRP1tEwDN/LUmg
7SFONnNciDKnZha1QQxPArCUos4XyCAe6pIGWP3yUNGg9z/ptulPN1cRckswfg9l
VkP+FUiZNdRTH6bdRvMIk34sxMrf5GiLbkQCgA1U3t6qlkIJ5Y0MhsZz38bRGxgU
4Yk/MmoWR+EpqpTxDXIALdKBWFpBXBRczRmBiEAnoiAt2Wmp3I74a0U6rsx4XDeY
rO19l0E1owADPBHigDEAZXEK1Ejmjp/YEUkEfo8tINhjDP205sUtt0DUjeZEcHjH
MJkZxPOffhvv+jPWsmxCR7E6QRBq/SqwnVTL6Ig9+LqO40xTVE8wX5+BiIvuZwkQ
ewLZdchrDhjHxr/pBY4f9VD4WC/Pd92xXwYFc3uS9uMdHh/NnPDczeycQ3Sh+jKh
q8aDLRPlJDRfh3BQm6UtC6TlzHpqRRVG6MFE+TTyXE6q5mMUxHCbgewvB33ps+R9
u53HdZvmAC83M2Ckf7It/GPOTOpihRkrDYVGCnRcd+wc9KOBMFt2FJld+K5ke6HY
OZZ6KgAZ4CEYk83llQibRwnR2Ywztrs79Gh+RXKnUBIs2KHCMwtFfMd/TDqa2iPr
TLLpn7OXH2rfay7Lrhd/VcE2hab2QYxTsbVPoDIUhqZnZP510XBU4RIRTDpkFfrr
T5V8upYggVmrQogyLp0ogY9c1WUoA0JTSrpBhSK9PELoZfwlV52/ARkkLrDtYMdd
+0V2Co6Ga5M/1OV09globE9vsI61yXIWS5yWpDIRK/HgmOjWPEFM6AXXpjMEOY6H
0WmNdsMPfjriHZVOUvijlvC6AReEwoUEdIRqhPLZ9Aa1Xpaywh5eEFUhB+GV2nW5
GWSxl5F9JrbrCtR0nSw+cO+sqZFRC4feJrfqUkkOelG/P311K3F/ihNewnsN+MP7
T0WP9XzKOdi+CWvbB9Zbu9HhjO9pjknT0AG4aSsh0mXEdjVZELioNT0upu4Qi2XF
uGlCRL/nqM672w82SC/bakVb7tYQ7i/Leg+X8r58Cw2yp5M3QTKSLIpXjFlo8AvH
iS99H4INTR5Z+N1W8jrSu55HL7Ne2g59RqqkeUVi6AiYeJ4X16ya+Z8rg/vcd830
dqpQX5OE+2wQYn0rOsnPKCIPQ/lnLA5UEH01Bw+BkvHx1aGDhjUNfVzxLR0rcXsB
1l/Z++Wj3DhxzAyjUjBZNhKEEo+RqkFVUdIL9A63kP5Td+1l/EFvk7dbAmMse06h
OrCjcw3edyv555PWl4TPXSofnqUlvzCefJmpshXr/a5Z3sHswvuI/YAVj3p/1qqy
Q5IDjAmAbJxoWBvkws9gmUUBN9tVu89wALOPqJaYfKlL0pmPS2vLPvF2WCeX3M90
OTTm2yUpE91JD3/Ct0PXErKsxwLiceE+QTcM3GJKrO4cTk7gGpN6uXudlTRMVhr+
mQwev7xrv0LNW+WDob1+uVJuSpIMWdaNhxSw2Da0YRCcFT9njAUQiFW2E+SNVcTv
SZ7L/j044J/4k9CmI9iRWAMx/z0sDWrwpNqdnfrDc+leRn7+tbW/JLU/H1wqywlh
bjKYtLYPe/ni19efQyCKFT6OLjIBS6v5Advmw0i8T251TT86zRSwAOmNLlF9gEoh
SIr6CqWlPYvalK9/ri+sxlRX6NoO1tfKBawsOOxu04r0DO3XKT6VFL3fVUZDhZQS
wFDAurcccW0jBlO53fV9JhkatGW6bXhvQl4AqVFQEnZqxELQLWpI5QrGovd4nh6A
1JezsKBr2rejyGzWWUDJDhZZtpddAxFYtduo/1XXR8nZcQNMH53XEyGVJ988uABf
Dtl2pUegewVxA3teSwhsQtINjQdoQLPY20P32XEvGrnOiyiffhz3GWutvZF+6H1h
UjSnW7z8wQy7Bd1YXOlgm38dmNRJFRY3pg4cUT+Cx2M5xhf4RkO13A4kt+fjczCr
jmuFM966NdTDLNEJtyrkpP2KoAHMLmxi+CL2pdF6ZwJC452ft3b+Aqb1VWj5tzSs
C/W7tB+EEX6CEuoARj7fM/uJ2vMoTnBPa4/LAc5PBnb+RW6pfO99wMqB6X8nn4k/
qBQ9Z2X6IWxVYvOWa2ikNB6KVx2ovAopEj6xDupUjNqwv5me90vjy6e8lG5AwkBJ
pRHHwg7V36oMMwhb6q2VRbm67pb8rjDrK8ZetgIYfjLOMYnTzqTCdeufzPGEyB7k
hPzjf6yPmf4V2mhdm0UWPzKclYoRE4MLb0xzIXnE4rfg80qXQ0KC2KdjE+uiiQJI
qcbVAGXwuB6Ex//tVCjg8k8sMPs7TVyzfkLIfsH3TLrYPDfY4FTG1HNDZHYJUkum
SQaVcOCy3nMd3AO2jNypNLVTHSxmRDtd3PTDXlA5GDINKirMM8Q4D4S5PbAqSIIA
xHBrDyY5i02FML9d/QTqEBBQyIgmpXM0cKZ2mlwk4VrThgqEyb9QqgoXRI0uPcPr
1qaWKU27AEBHjuHjrT14G9DDLmt9gBhc2v9vpisCUQd7nFuDFYnYT52pIXBugCyP
T5SXPbH0ZFAv8Xi1GYT7xveci4wK0bR8gZbt6wIP8lTA80MXgxb0hViLONrC+zU4
8J+Mg+c3jOYiHCEQ3AgVOnzlUV3r94yrEq6WXraaF623FPJ2hIL0COt+kRN4dfkX
4Ch15aT/DMn85yby7l1Ywb0PM/3D1nDciqXACxXUVr/K47cECVObwRwdbCWmCsen
PiolgIB+gMPIxJZXMcrEE5VyXrsJaxAi4y/k4FrDZ/nekvuAD/AsSo+CvxhKUUs3
xtAQjA0QqQDRpu8yj5w6rVMH9ODPBu/njkiQ99wDarMWsTxMAUCTRFI1KcWOP550
Ibw/pKQlPUEn8bqr3a5PWceMilEmjr4ek+fISkYfb1C5hqrwzCub2RXrbz4GB0m8
5tG4MAkG5JM8CZXbmpY/RngPP5PN3buefeUCgnqKnbzyV8hPgFL0UEm6c8K5p7b7
UmWWSiEUuuaeThfHceqBOfoQSmLP9xgSzKMHFWcx74YAazraXJyV6Kg5VVPS4hz5
JJdpBYON3HHSlHM5i6L8gLzKbqFKdRTOHypTJeMxdwHNt6Ekd5n1DHGwGVb8Oj6B
RUCsiaGcRBrTM01oJPXZbwdt4Y4TIh2hUeMeb2tazVz7AFew4v+beb9I2lDcVjFv
FTr8fZCsme/DKloUj4LTd+4LNUM407u2ukkeHzoJYan/9FTISuGQBU7paZrY+9W4
FeSZTTitXKOy+gdsE8H8Ogwpiet9jL0DZ2wjJyTWb6IsO9viz17P6bJOPdgLL3XV
0xaPoMc56fFa1CbD+e/VLBmPCGGAoOdaeZLwaiNdfAjoEwQKKabqrGbkeuIErOML
HDFIn0STje4Wp8WML9V6zS0tMOpAm2zMuJUpXtSJF3584DH7vDLshRdvdrVyzY8a
7F2EFK3CoUhbLtQRzC8MpOFLcbORFDPj9tBlAfVYVnISVvViunRYZBxYaP39LfaN
pPys2BMpbek6eGk34rKS/r2oJmuBSqSZVaceLe5sBwg3KfCsjMjTq1YYPyXVoFaO
45IHkihRXNdqjrzDnYMPYxkviU6SrQiO5NUcL9iCWlnjTlEEBOm6m4qSk7ZLCMKe
1VxQ/N838MKkpik2NSOEZmcZrQudw+aLMv9Awm8o6qVl8N/h2WEyvb2LDmPxj1cw
irP2E2UmWamzu7PeDO+hEwWYNhhqgUnNkf6mutl+dg115NpaS2hOflmxfvNv0XAt
bfhk+ge2WkF6Dfy31S806v08s59Nq6mmI+SqYkfnJFKQz2sVa0ZYZ9A3ubakWOuc
kO7YHA/rFQ0Ofo0TvH2G2JK9zEyUq02lLvHNM5R0a9jCZQH71HSOhP9hQjzOPFBe
oyJurrRVW4vI3VqF7Aazv8JZP+f5d5L28BIjlKE4tkcaFxAdcaTZd5SerA0ZdCR5
w2cDN9GI0vFTrzP/gXJuq480HxECbukZQU3jmhQJPZa9aFhALtAqMchf1nWEtnoT
2Ep40060EMFCyoxGl89YNpQrQyTJ9TIQ110Wk5PsGWCW2gfOXUGUlws1U+fz6PJy
K515SsFutwPbDprp98FzmS0dvwJVZJ1KkB+2lmFK0MIeOSDMb8Djxix6JGBbMYA5
S4veIZQx7FpasjzOyr8Ru/adFprh7GMxdu0G/RkOW+kmrSMquZpir+h2TL9PEk0c
lM+78j1HpxDD8eSxtj8S489S6/Rn2PoR/mFnGoIBiZiNmks0pFgDnekTz0lyDfWp
Cdy5sIl3jJcmi/SWze8pBXOKvYXqqBb+UKtJnSn4n9hxaNyo4nU4JD8lY5T6d76M
EX48w+AJ5ZQmIarAUKgZzdXgjIaT0a+vmG30ImHxQ94jaPCEQKqsN5koqmU/C282
MxQ2u1gxtSTw0FqA7bBkJTZ4qkMA/In8rgtdYAsmii6c6VvPQroPFBB7KI8Poppl
4YQLtJDBunhIE/UF8bMAwoxXiSvGKNdyQnQXdfJPorf0bDLOPbr5inIqVSjl0HxZ
3WUDG9a7lzIhT/Lw0NZkK8fikKnSGSBnf965w3z8GEYZ7IWR+U6Ly0LSEsVBDmK4
pkueXP9ioarL+vl8xYSIZSDJlBqrXkTVzVZcMy2O/aqPgxZ6SbumIjW0AXBIV1ao
ViwyjefSCR7xC75EIBMvakMkV+tMj375FmMeshpN2Kx5G1TFpWHi9ax03ukYaHBt
/w3mbjYRGeWstJMdeaCGI8IgZhkfSbqEk4hsAEbjMXTB/G8P/fEK4ZiWQKq3ipv5
jBfQhjzJPKobYTQWW4lQSJb8K6RL+joo+QwZweS2CmvYUN8Xo1nt0rcTUH3Nz6DE
uVSYaiomxDZBEHYFAk6OnT5BaJz1oDzt188ZjwKXuguNnE9nYtgHzLK7Sieuf2j4
vfLgV8Q0M2rfFFw5sSwHuxh4yVt1vyyw36Uvf0Bnc7HmiIs0ZoQVfCwfe5RPy7tq
HuVosD17KU2amUmuUemxCZmjj2yIcQdu0BKJ3l6irMJJy8js7OaTxUECS7CVb2zk
olpS9OQq1+KJiEeIfm1g0ohDssBc/ZcXKm5zzAsgNhqGLYcQ6IZxhR4PjFP49tzs
IwwWhPYzyBEojPCusE4R4yk9IyG4heJTzrYrOPWkknCuihdgFxMsYzvWV10p5TAs
tABb1sR485V0vMy6j7hxdWS8wXw8GKypginzPRdDOcdF7WlEBrhOCqOwAghq+CNM
zNSPU/vBAbvUNW8qTpK+iLDphnJwtDYiFfMgZGXuWEQE8txxnpAJ4NI1qjzSw1MJ
aP7a+B1dUOFTBqUobTV+N20cRKm+GHNTrCyCK891itbfrr+ipxMRHdsgM/jZIPv6
HUKHFAbjLIUNEIvuEQeC8l6ERpj3H3G2l17RJA5peTdy6CH9ypPLJ3s56ppHVfjm
y5JVOxz10eHDX5o1k9yY2NR4F8uNnftcAb27fQJgtlq23G4VaZnlyIGlTYoIjnt1
XV1cADbsBP9VnqC+g9/cBxx+/XRAhGXzrNqqsK+lKgHsTHQyujOsypJ102jPqbD1
D3bLxI0Dea090kViHyS15moyOaDd5ao0rJHt8UvQ+QGMQID4v2QGIOW31+4JxeMY
9fyRocIqUk6O5nKDYzm33tRCGvhrQhIkjM+vObSHYqfVf730oDwp1tYXNQE/BHZn
eViX9vg8P3kFzI85kFznCmb6Xtagmgm0P5QX9q59e7R30IOQNCddicUCPYW+Auzx
zlpEkwFa1Thu+cFHbEFzvfolSQCwClzQ2PACq2BvSDWxzAHNO6FycnXha6OhSY5A
5kM9jRmbFOpxgecmXxKMAMWfqXZ5j1fKUY5r91dH1KxdnKjj3ecBVxEeNREp9rta
kQmqLdhhiCBzBAajp3YsEjA+kEe3kvCKMZUG9onSNZYiyVHC6iCGfOlJ+huE6h98
G8vLJCRc4YnhxYhRk9RkPoIr7Pxzb7X/CEcDARyAnIHQGq0GxtmLzoBBMvWQTNVp
EWKMDH7QjcYfyMCkfnUG6l5gS8wkr34BwGCFq2N3FfykEc6DIfHqiksO2YxEjEHx
HoEZQugrbTRoqTLPYh6Uiv5Vi4FdecF06yl/Fe03Sr5UL30tkR+WMit7XMK6f51Q
4Nf0jw0tfgXiZW0e8Sjslc9shH3uGPJ5UihtZ0KU7F8oDfwnBjw9XwJBxMes7SG4
AbVsC6NLoiDA795M0Gn96rAJOc1vbXNb+RY++1ytZg/mD4blsH3MtI3ZpX84wpOG
AoKsq0yy+uGXI3ekpfHC1O0P7sfV7VvCWuXM63Zo7fk5QsnQRINvKpJJ/XvT4JED
XXXbvma3Q/eA8qpMAEixaECz6Igu0PR75xCBiSSKTKV/JBsVyHlqe5g2aXmObdk/
g6ppo4Gk6IGefv+J7VWONRiS8l58hqUv4xDa/R74yWbHehcSYrCUoJ3M8eJPfhCr
gppKUCO0t2DuBHt1UmxABz/7MT+4oGSkUF9CFx/+4LHzq12wUm2cr2g9NhTRRfak
iKmHzxJw5nJBaRmU5fBjB7H4l8VUJPSlpujIGnfCjJNXG8l4qcBqmJ8i0rHVCpR3
TJDDfAbOjw8QEg1mMtrtet5FT4Etjju6Jla5XrRJbZbgFHb2GkVKiX5O26UAT3VW
FJXkDV0oOQ4xI2b+lUzQ0vG4a15N2+ew6iRH+2YcIBlrBw9FLN1w/XfE8/cHDDME
24DS32ZtY2DmT2ffdzyhNldPZ2OTBBMTssDwcJRsaQJAg12DQtWi3UMjT9SXodFQ
TNQth/M8Otju5resyqX9iE6OPz2vpxN/wRbFxAGSrHvVMH5XoWXX07tzgUre3NQK
ULZ5ZmM7V+feBVKTa0Ty5IfjzcXux9TNFOy4dlds4pfL1mHhxCGtcVqY7b2vLX40
FjQaaJXPmGgEHN9195XRrKZOeE1HhCqn+zVuiEHox0w0sm5CYQIr6F2GNLtXfMdC
bVPRS7PTf5ogTjerOXxoX+G9z0R9e9jGbPDYl62ELAUkJBcyVWb7Dx395Uj8EtLG
E3inH0M6fvCTqCbz7Dyn4f/pfJL1kwrbrx4/MekQdMXmHZ+CXJ8k/1nnu68wiP5+
kcK/ISl8u/88quh3zj1dgmbXDFggkjtmfHUGRXzmp584GsH6SxFbcRAakHFhjUlM
Iiend+YEJB5RBkp5JzhZd/gT0SZbRZnwP2ZMMa+MQ+mEMu6BicIbeiOJnlM3OfPt
w9mzBsLxqviTPpBs/gE0+8U1729j0ZDskF1kDfntmYAOHpccfFCrZyelyZSF0R6H
hrOH9+aOfMqZw2SKTVMv5paThH+spzgE3BuhLPFxg3ZpcMOzvzhmZ9ktt6VpVjA6
7ISVM0hhjdtgJK4ODl8V1waTWlkqdAjTlbCk00NmlO6lJgar3S22d/y/dF2vOqlS
QMETFZ3NfwZD2fLSgxbLNMLFA0LKFr8cH+bp5kCvvPk6nTqIHWa65t5K+k65p3GP
t7wnt6W6FMtEH/zbqXGaTRbIFYXL1qCoqRrF1boiDji8fszW2EZJvZZ83ktPXBUo
j8QAxGUeqPbv1zvEkvODT3p6C7wA21BeOKNSrSQOVvLp6sgjXDLO7ovjMYzf2IR1
ZLB6+q4Re7r8mHSIRIL+Ib9aCkL+p7A066XG5sIbOAn30e98LxLJd9ZqGa4bfozp
vchAoQF7Hn9jOUYLNdMmK9PqzPpLoJf45qWXcMJPKX94HdvlLwLQ6Tsnoo2VPRPF
HE5xMyaTwkoTgso9exmP2NrVwZmBF4/hM8g70nNLKPhBUQCnmHcZrNckPn2uZTFc
U4pwzgin9o86YJQ5E1QMmpcXPMEy4FZhKATx6ZFd0tlOfjoB7ePnmMMld6s6wh7h
gejngWOrXCTbqWP68ApsAeblIuv1exIOSv//Yr25+a/klUNCbp9ZYF4yR4U8l7ZB
CYojX9Ontmwre/Hb4cIP6sWlxUpIBoDgK5w8noCQG92E9W3zt6o0vPwzSLjfIT82
S/4DfFR7+COE59+FEImq65n2BsTgX3oVQ5Opo7sdlny+Zrb9DZo/b1B+l2FAvHek
4CYG1YD4ym2LWdu3NCq6KvgGH+H1gGmgvekXcySWwqv7CrL8jKG7wEvZgywfPMtE
2rAE+x6eDf2kCMmHpVo6qD8fPEzr0SyrtCqKtckj7JYde/3c1DHAsASe1blh8XH7
1WFR/NEg7YI7eDf0Hxu9Hm74x+lwWVS1wGZvxF8Ug6Yp2SB3GO3aeHFTOPNThpNz
S0j3EUFD4wb/pRa3AiLArXNZgcBucEZ5FgkhjZtstFuco9Eqdw1vtxrhERoRGKlL
5k5wxNshCxfX0VXgMnFlmDoSkHwO6omGa4mBMKqypFI77uWOSvQIXIiGDsq2b5iJ
6Nai2F23P9xhwNYi3Dy9jfj1/MOVOw9p0MK48BKGTot03JOToBrHAERzSLkvGddF
XPXLhziJwhsYhTybu+1CoKDdwfYDdurqI5VQCmAbbnQaD1Ghba/qoxcR93VMpbQ6
UIssQXjPQ7DH2AB8gsnxvOmtPYz/HRYy5ox2D64GdHBfimx6BMeiaCJd4FcvtGvX
+nOwdBUYa7CJ5HNXFyxxTnyNh/D05pdGLj58X6Zu9+rNtuo4ZYrqpdTcrqLPxq9i
zWK3+63KlRW1ws+3cLbY2jxCUIhE8IoTFah5JlZptIBRxRPqPVnauPRSa9g7gzdD
Rhnkn6IPz2W/NmYkGHVL/DpVrefCikaG/Yq9MhgR20LbwVvPIlj06GIYh9hrAv4W
pn2b/xWVK89wnoedzuT7HkzLt7kJg9brptaxGqddnTmVe7o3O6frWG4LF29vZ/oL
/rG+rxxKiyRuvoPue3lFsDSu/aTYOSFxQ71VQ3YudZtlpiGNoIdLv3oEjC+lCLrm
ma65ezZoLPNcWih4frTjFSeESbQiHuko5V53JRxEHGdY4NilqUrv9cb3m1Kx0f5J
Rg52OW2csnpxlKm14sBPP6u/vtrB9yXtLm9qTdVk/VBfGfunri96h1BYjOfubE0t
uICG5xR5QV5WRdyfiPsgMGIaHW+UBcsrV1dqRn/qy2joWHcgaIQQqeOkNJZit3bB
Qk6ZNzURYxKZvGBG41qt1tZLm69BOrzL0qP9rVFFPaKMZR8ZWK1QTdc6W0CnteGy
MDOVwfeiATi6MWPwSiKzY7vgl8Zb6zBWNH4uXP55eBwQ96nkG6OczoZXWmy0Hk4V
tsEFT+L9SMmMoS2qALXhaHCM6MX6GCNMFLH0obcmka387r4VF+xee7BwEsecNuzb
LxgaOeKa91/XEeMtvGCjongEk4PXxD28hmcolwHAEUJ/x8mJXN4ju7lGhHvLpwqG
9eO9fOsfkdUD1gpU3rrd3mxnkYbLGlSDupoybGFp5Jlc81IpqJuMZAiPn1zMS+v2
OFnAsbA4y53NwLt97xZheiGuqdGGGJqpoJXD6vtciJTRpVjpXlPgGtoolTJvXB3v
QQKPQ/7SCS13X3NKOiDWSpxusF5WmWFGvzHevwL6WpX1FVzcw90jSuJzAng8PcVt
neU/jgeFvQYS6InvzDrYe4EqxMZx8g4COJsU8JUOalYMp/Vz/z7NqOkW4HYF6CW2
0hvxhxPYwxWHUkYz8yIa1bnsZWD5ErQalOEzNV/GzvHmTP+6EVE4IYQkAuQZAZkn
t8kwS/+IKbDcYJ8zn+Z0qQ5vWcrkQa4MxiwIH+UjJY0nP9OfgsRa5wLTsrJLuhnK
wZWUUMOtZy1NGqQF/YaVLhJL9pShzFlIv+5OzEdjIQ3epP0HvP/HiEAU6VgpCt1m
2KDP0ErSO/1mbOTgAqMDpWFvcPjaVhcC1WVFGYZo1Ofm1iZQVAcEx2JP2s4kJEc9
PqVPZoBPozzADuvjtACM1kcukKDmNB3QqpopvyIonoM1hJr3rlFoGurlYEWWgDQf
MUJUUVsKd4ZUGR4et2a9rWR5gDaiCRtZCxQzP0pIFmv+XEJkrFwQLa31eR45/g1U
Qy9txsBf950wYgD+U0JKAbTFTmYK0PwdLegksUJewYRwU4pbzGB4NwVndRVz2EDU
uJlq7br3mgHwv671bqDreC+vRW39RfE8EuC2CSDqWrX2e2addAaSRGKY1drg2uuH
L4G386NWEN4y+tsFLc79fAE9rak0sFkvFE/2p4XmmF9A3t5u/wjkF4ovgLHfk+a9
DBw4BKslf8zU/s416Ipo4Bveh1YjEZYOc8qTKexbr+1TxlsuXjUfZ4OazpsknjXD
/4rdzefBCK0FHCzH2K5pfABEDekqDGhAb18MdGx0U5boR8ziU5sUbEKFa3FcA9+l
zqMjF/UHY+PO9TBz+Ccls5u7hF+9ID10xbO9zDLuJIzUv096mxyvjGUPdI4yxWog
90ceOmjPqmqLjub/vjda7AX/8p/vHBG1oYgZwXf7itLO648RPMUhPE9k0ItH3hK0
LEweqbrXwuYywjFwKqEvJ0wSVi9/RTeik3lyzKNA0IHK/haMvID0FdHuPL9IQJ94
P7IlD6sxF0hp8LyEHmWw/LyC0ldC+DJZUEMGybi/xI3NOOe6H8v2T4sjlzal7WDm
IkcMop58F9vH3Hbr5n1UfaHKn/6zJgPXj5dRwSdgu+B1vOZuKufIYHD/kpqSOSZZ
i2ikwWF0YPFcChm2zsB4R6Rz6C8d/XLkqUpBSxkaGuZ7QNDTfhg44elWBOGoo6AP
Ngvm5aYGzgIPVlQm8VHNP+VA72qOW2otq4Q7o7swQQDhvqir/O0Ahb7oLB+ZAoP3
HBRYmn0t9OXM5xIxlvpxnI3/Ggu2fpaT+D45N+3Z+f5Cucu+OQFTpUPU8mWM9MmR
Z76NFgJZcoFIJ5XFuZ1qc7BWdBQMB73HkCWtOEZnGizR09c76G0jiAIe9DtIx5Pf
wC/+r5qtsjWz9fp3xDeMchy40RsS4Ab4fEVtjdbu/DLXG3Y1PdE/BY/oCCC0cHMA
Zy+xENiwKq/AHhnTCt6reE0iUnNFt9sTHt2BjvbE2kCQgT4X8D6yRuv/mqVz0QRh
zCGrJWTMvqJEw1PXYFm0JA8AR5QuN0gpciKZZk9o0SAIYyrvci0kiQU9bK/p5Tdf
gL9a94X1UqSzQa4LlV4V/sXG3a6aOq/mvm88NEFpUdWUI+7WUVtuvRbJnlweg2Di
fWOed4F8hrQptEQDsK4uzqA7hlgAUqDjbogv/zEmW1J7J8gkTH5KQE9KkfFM6XT9
H3ND/KP2DRkeYEsNjf0WDCxfqTryji2N6HJhNlSwqN3IGVCZDMU2X+XVf+Ub8X1X
aiaY4OmUK5Cg9WenSPbgb0khzHXXkKBxeXxG6s1S7EO9a4ICy/5fezx3j1MxJku9
tPKw7LpuofjO/eQSOjrt8WzDArjRdPfuB2AYnwQsaC/Ox4gwRyeRExey8kCehdnE
RPZeQgO6SbjvOho2VMJrNGdTs38oJiWlgyhKiArGN1eu3XveSfYty/9Gdw9yP4n2
/slSMXwa4jMVKciXaVyz5B6e2/e5GRdfyF1GjBO/qG5KX2UUYZ2nSJ78EjsvQcSb
HLldlGlDNem0o4oan3MUCKQIRhD5r8vKQTw/IQ5qbs0456+/U3mXLqNTaqQzDRCb
M0Nlv5MG1GQAshRUmCS+RZqCqljWvMpCOzqQhtEK6ksN1mPMdS0zOauCRZDDT7S9
SqXZt7hM+XqGSnbLsWSDJPd3IUcI1BbTEM8nqd3zl5LlZQ8JWnBB6YsvFj8BXpLU
VTk0ofLSVdwZ6puNVViYvop+nyO5T6UUVQIu8AgGURo2sGvkeGrfRwb0/WYLw8qV
TkRUPLcFgyDbOpw2Ijv/QxML4723w+h4o+98pOrUNzLJ0uM+PrK0lcRFWi++FaBp
V5Jc9sKdXvdAD7xaJZEsyVXELDr+S9GOkz4DUp8emDGcdq/9t7+pHurzs/vrJ3UD
HWv2RGRs7Lp35e/3/1GhiV919LSm+lDgi/S1dtllOFsXkFpKlBMvS8ixq5d6//qO
rQgaNJJu6Kss4zyaKR5hkWlSLKoHwcsj37NMqugVp7N5lVNQORu1RZ82wdY1VU3z
E9+ji6wlx7Pg1nIJfT3GL0s0Ah1xtFcSxDhARnMQ6UKVNsajA1Trb5qcKR83uDVI
pCs8OCGjHacmeE1ubXAIVXltcX0QDjSPyqHAQOz9iOoUetU5U9pg0pLjpws6a/+5
MD2ffiXsGQx65gmE3jTyI2b0ipzRbpV+Nx+jdffeG/nOSkI/OWp4wNxyO3vnQueI
uCYfUepQXAy8Nud4FtrY0xRAna3DZvcQ4W+r1/I/wRL6j/W/DqS7VtP/SzQqMj0r
xDQ/+g521IhujRnih4H9u4Cjkk1vFO5KVDQZqqrvwA6GCq5PSIRkjsP3j9nbIsxY
rrHP18cdNXAL01JCb0GKnAsmhsBQDuI3P34oAf4IrJjs8hoJY5WaAxBUg0Lgj1Mi
fC6TJvYXyUotTAR8o7nCztsDX/DdlgRSVTs7HmsflGVtiFIg2f6czfXF7qIJShnO
/9fuDQH4KpywVwq7e38pr+yBJ/jPie7KnsHayEwFXmpg7dHTYkCuvF6AeVJjI1mu
ClPo+4iJ7D+D0a77Kv2USgcwAAGbpLQSloC0YQtl9CEl6GGO2Y3HBGSOorcgJgq3
G7O5Qo0P3lNZXSsSdkPa0zREpY/ewcLSJ1TGMKCDOjLROp+SPpBBSsFKLxO1NzFj
2H/RK/lnNVup+nXzCWAKwvEFzxXrZTMcIrDCTYS26d3Nm3VHknLcLc2R//EBjj/L
qr60Dzp1KHIBZdrYLn3ItMwXfFuN6Km3mDZbaaOj+H0qJfHjFNk5xxK3BYE5zO1R
7Amk5PVu5+zND2E66s2W4+O+BEe98VE0I+XWmXRR967OFm6AnSKXsWXpcEhNyDj0
r5tubqjQVw7ydICAlg3HQPBMP1HJT0nq+uiTkPAH5hg+qmrjdRHr/wcKVjROlQWe
W3Ds8HQNXvn/f89euQE3uTPS2J6r5GsKj5JqdGoz8aMb1tHRPO8l/pVAJawLoAPF
yiRixPzUb0UUWKpqk+Je6hQKIgWs0srNheOsWpAqLpeOwZR+8BxBMsCDhvWwLqEL
AEFIq93e7sgy0q+/Jf/Hm+WhM/x5MEtLKcNAsRa4keBIF2++UYqvtrutzDIVIGHF
XNVPLACsDKOUuB3yALMAHphO41uuX/va9FqeJVh9ZNV118ANpO/EimaNJ6Wby5A2
nXmQTXq8QsALYxJWfaIjVEz4rALiGFNLLTX0p+arK4hazMSO6ly7uDY+QW8r0qIm
KRbcyHfRfpdhTIgPXwY+pRzpQarFSdxXo0IqAIdZzyU7xJ8Csu9rzM0w6A3Il/P3
jMyuwvBhPJ0nzvFL3Jl/v7EzRpqirsozFLCSyEkScqPe/m5fJM80TVFTQCW/AOen
WAPLj3ubX03giaHsnkB94Leu8ovJkfetsZQvLqmHICPWN/vxmKKwktNNo09tZyBq
HMi2RirDRJMjQUtOb9E6ShC/8es9XqUrNRz+sa7m4oD33Q7xossLJRfFlQ3eUR2F
2NEQejb5LMb4FgHDWRPhMaGBWnDDCFi6IlM3ereY05jZr2N6lwM48mGZ0Q62yEX4
qTqgBlFMtyJxp/hsqoeXGieyOK/eSzx9Hd0QeFGKdgfSF5z1MuAmj4cxoaSO6RJ2
K+J+W0KOnsvrojpbkUEY4cgJWnjIdLWgUDlBmKRXlJfkxNcxsy/1QMUuRsrEn+gf
n4sAnqF46XrQPL8lT/1Bth0JBNneAeEUAeFgtTkq9i5qzu43WtyuabghhakKYBqZ
0HbLBCYb2JAFb6AQc6mfI67FOA/dEzzcr51TZlSOIWIfksy8rFv/aETGuS55iAts
X+l3QuTTEYe6ZRDGWOY1Bx5WWRrD+4TbpWkFTFDVoMgmdz91iUVZhLrvja8U6Uhy
6qmA2H7WVgQCCggmatRQekRaKgGSoJLiAmEz6OUVn8LeHCPqksRCGhpfnFYOWEoX
YJi6Y9Bg0arW8I/2ixyj2vrPs0AHiIaYnJhj2uyX7upXaD9CPZURDhxk2Lx6NNlU
cN2cNWTe8YLodvJWy7X1rJGDaQ+D8r1nIw6JM5jZWmZ3ngvLh3eKGMeJgNNu50ME
71W6pVJL7JyQZa/5FYZKLHYb3Z8dShnvGbD7v8hv5r6QiwgxBO/cHrT7UPgTq5of
Oykd7pO7pD4eQ29bK1PzHQiZkfzc+x5y/PoUKiXiPNKauK7bwGb5zduCMmJXpO7L
77TbuUmgAQ04OO1USOHOBvMsJ8zwZj3IE/MtnH0vA+6VXnwFcsedljguxmU9MXWo
kcrfmXOan0pe8NpEdxRcOlHzSknA0lAsXp/7KdCNtHTuwGejFQ7nfFCzbezPa54c
Q3y16dlev9TwIK/wPeUEuhldYGg5braSfm9tMlXvXw81iHNvjh9GQuLOY67QLvri
e2pBX+m05mNVpNZ/qvf3jVztltUkCoaZpw3jgvl2sCx+Dr3E47YMNLfniMz+XGre
D82Vj6QqzdXhknYbMr3S2S1sYnW9bfxP6rvZm2k1KUR/d4br/1IaYZJBgT95EZq9
6rb+ZsF2HMQOCT/VDM2zR0dXE47RElUREN6aJWGIGRrts2cgHhBaj/1lmqmu8iv6
Oe28C72ow561n65XWc66Z/caUuIME58y9my5xwqYYs68cr3sFhbwDxEobxgklvYz
E4Vqnop0CxqhHY3IdU7yCNcemOFIuMRKnh80csAuWc4KMQbThWTJ+yMUnH9G2U/s
qv9fe7m5/z9E0mEnWwGUfsM2pJ77SdnIdxHdPFth/cjsTw5xzmYv1n4mcEGKdBVl
3LEgXAdrwtrui5MZaqzZFefVwVJ2S66VXZlIYGRonAEuXzeNg582XDcj5jlyUzDw
02TM1Xt5wHLDzBhwGzO9/Fe3DEmFzmfsQYPXdmZfJ9BUynnetC+et9e6xDuLxT2G
0x/YMe39F+igM7FekaQn1JeeqVY9s7yHfCSa5e1NJQkleACBDDTrw8lHONnHYs13
Ubzdy4RADR0PsVBBXywJkSXdto//zARaVdrJzYm2HSbuHI5Lcqx4vjUatJ1wsG/t
UbfSEG1pkZSE05+vHKXKWg66kIlzzYuW+qgmu2ya0zYzyYyk+enCI4YrgGCgVcKG
qQPeTBec/YcPpG4fdM57boNueflLkAv4xH4WZJQtciTT814U8miITIVLijVbzmGS
UgLGtZHBpcRfK9eqaw1V3tEciwx1wErv93Ic31YGwNJGSjLw+7lMEjvhRehVUGFG
K+N7gtu9KWS6HeNLOWZEjjpzy5C5bdVQg5e6oCZBRY3XMVTVZH1m7pUnTLVYEL47
4tmTjXbcWXhGzgBnDzh2PKYLBl9jjdjOEqXrk9toc2tw7Snyd9b2I8mce4kGgkPN
ke+KIQYfKFcAiVkHbZrjFudoEC0x/OwbeFcV6+pVcxr8SpAqaVYSnlPa6QI9bXEe
6nNQGQ2Yctv4OY3thhgfrGkXc6sahxeL+Ao5cB7AuWvGjq2I0QA/shSrYmod7qLD
Act7QFj/6N49I8JWJn7kK/Cke8c0xrdJPxMRed+l67tpDuEYllnc+jwF3V+uqcQ7
TjdErV5qAXKVzDY1YDejd/zyov7W5CV2RA0oM+qKqKOgwK1LRV87L2wwLRpV9yZa
sNgnhW/cGZW2FtpyLn7qKvW8Kg09XOe+HhQ3/nhNVgLUr6YRwkHhTEakqs52JXOJ
unxOcZRxHhw8tIs8g6jVMZKRHv6mxd0hw7mMuIKA8nZ70I9ji79x6hgY8dhb3Ho2
zvAOsRxDhh1CmaHxKFnbpExZqVq5Movp1QLNf/lyOtQ907/VC22H6ERfjal6u47X
Fm0GH9vTe+nIojyQ0OddfPISphQ9AjuIh4/IkpVp8N3+0Io+wOzksD5jnPV4GGtP
QcVSW3zOkmWNXLjZtoTYw6gn1gaIEY9NliTY6K4yu83i/euCzhAp1nihfWwYqLL4
djySOdQKRZhrSxMLTCGCOcKNjZT6cTf8+V+OaqKlsE98J68IEB+0LWmQRVMmWP8u
gFAEv0vPPz8+wGsDi3lFqMhV+906DMdtt/1cTBN5yBggnfuOj/C8DTwvRHKUa9x9
L4WTnzFFyW4kfDMan5JwSfbzDirAmBWG/jJVb0BNhno5nezY5L8hrc6opgFUYYR2
rUq/t6QTqTgdhakuyj8+nA4taJTuIer2RUcBlNQCKcS34G/5xH8iUGOCj/AQTiRB
DzyVCi1dcDNqaypRAZs+ydfQ1RYgT4KqSY8k7Is8vaoHFrdBaXtIE1hXLXIVKU2L
tF4jE8J+EnqknD2MZDsDSYoctBzeb1C9EXpysGTvzBC9a+OlStuvUYB/Wn8+xHoz
GZMFIihaXi493m30Qjm4bP/Oxkv+Fp4acOpgaGswgKe4C0OraH5FJtqSMQXaIBXP
AOz0Jqe16iXRFRI7NFmMs+QFtdaImEL/B2ptFw6bWUBBXAGqpNRfLd5/unvLyC1l
+OFYPKd/Yt8oOMXghoCX8l0XKxBzFedDZLlnLv8CWdiImpTNfxFUpc2TLW+aitK7
7Ggi9pk/6ZpqNg+xfEGJ6pyy7O25yQzsmAFANaUuX22Y8TnHgkIFuFKSifQ2HswR
s+QrKOdFRr3oFEAwFj1Jg44+YRN15IB5sj5cv3vkdxjp412WrWRsAam+ATIBpkpW
T83vTVB9rnry0Z4mtUnRvNXJNEAxzhIwxdXjLBhFjFRpS0o48/5SlHoxsZ1XfF+7
P4JAnNmUIqB8HXTrHBLYCg/WvxusewJJMeGtacm2XClWrjtu6fBNKhyahD+txLlj
Ob/MzpoARH94psol+dmXjC5zz3rfxoEO+cEtg5OgGq6/KCdLu4AdSZt0jwxyQ9d2
ph+T93WxPSWnldNytm1qtoVgPCNm/BHZjMaChCP79YgM9k+V+V+I79ap7SQdFGf6
aGL6zw1itG0NXTlLqwAuX2pDkEkYT8EsKp7sirwPhxJHtZP3F7HrSpcerOZUQw88
mHGSN0l8GMFbho9jTHUDr4S902QBbCCVcKqIHDlNgj3OnarU5AqKHvduW+omquLK
spW73a4bjIkMNsUcQf2qc+075uWcKCAxN+oJAMoEnwP6PV2ECkiUDizfQXkTPhvZ
xI+g5zfTSVskNxC4k1FSvJYI0Ux3UuLG0cCL9IpeHRwNtvTuuXr83FppoJ0dFs3c
BQEOP8bEAZC3bxCO0u/LcBHtmm80tx3h8MVjCpeY9IKU7Z3TWuNaCC7K9Esaxopy
OkgvpmnYHOyMcALr5xJnX1HvM07K4lm6VXcGu9cfr99kPVKzEA+OZS0pblpp4g7Y
At5S3LFVg28/wM/+OPeyFhs6dcjtdqK9fzgkHxvnIMppP+C1BzQSc296m+1NoUtn
Gq9ovtJ5zOMBgMaQN0muiSAjsHavB5BXcwjiavrfqBspa/6k0aVq4/aXb5QMRknP
neVeOCCssFgFlJDAEefbf9hvhaoi93DHh4nUVdW/i5yYezfKbao9cKkkMkYzCqao
cXBSeikpQ65Ydnk+R9kxIcAXWL5Vpbv7EQjC6CFGuSLEGhvLxnpNjZ3ZAb+/pPoL
/ayeLMoztP7b6oEDaD6VzDJ3swqDma7pveP99lSeCH+jSWE0ajInpNEoCa5Egf3E
OJDvxj/w0VetIuT97j96PxPCBhPFYCyaB8+N7hL8q6vLe13z65mbcH0w5Nmc5F5D
8rw4Tf/A9JVPOBd9L79FG6RgmQwNydP5c2IK06NEIbPzz3Gc7PK58Nl8jY9JC/jd
HBHKSxnaqXLwMSxaMR3yrNEvZew7KxN5pJ7YCXHJ/Gz7N6TP247qreO+C6tfzYRv
eTa2TAOSW2KV3dgsn5Kmjmc5fhHsLrbrxufWQuHyi8QHBIBJV+2YKvOmHZwxy8kl
08gicdQeq22cwEze28OUU75yQHm/nykySwdF0HdObo9wy1yQaV+oz0YNQ+gAVfTe
dRHkpViqnWa8aVOgwOuM+IOz7eLHao+OwM05qCu9w7r93qp5Ybv0e1GfS9IJCFFv
0WF95nfBvSdaW0VTxx3sIfk/HOuBhVwbIlQPwmUnCYKyJ5DPffbZcgowZ8fStd7c
5tyZJC+IF3rj0CjD7H82OgBDNOXb2zMdxaUQ6oa0eAuB1Nt7DHUIt+AmTzPmQLAB
rjncHh7Pg855A9KvkWsjdZSwD3zQa9jN+Q+qOP5yGLjNPTv0ltwidyJOVBKSZdRq
LnsWP4CAOxsHbXdejG2+W4SEKbOKqRBUZqA1xfipbuUp077/c5FZ4AQfeOP7KFeK
Olb5QLDCP/mupi2SJJEUCDcNGB31vKynXe7utXf8w9RmbtQGtP/moCHsA9pAU1TP
tEnLKben5ntmKDNFjzK9Y0mXQuZNq6P3u26qBpuU6mLcJ8Y3MvoRGxV6FUhhvfk5
5rWJB9zW/n5sGP9munJQ/VuvLtw0dvNpDQxMq93b6Whe0E1nlx+mZzc/1vzTII2g
5R9A6B3XLumyk7OtqoBvVi2cCK/xLzMdBsOj1vXROFxrMHvkm2cpCYtvz1TEYiI9
Vvaqw7tUmN3rj++1x6iGY0CZtye4kToyqrob3X1GDjb8kZHlsDGN4rAArn/8ewnr
9QRVhB2pJfUFXhXqxjHAjQ8liUjz/+tV3LNqD5lm57+/5jJU4zbr/A+9skD1CV90
E09IpUYhG8b/gPK2stxYE3iwX4S8zYUph3zr6rJXJfAuTmbePzzXkyowwYFNiGzl
DcLIIcE4xNdfFvJ6WZ9PEvSoNBTppLxVLybQyBGodq7HfbFZjoTHQYJR8VpjAIwC
Oklzlhvr97KYTcEALI795eUIfZuUaxNxq8lPJ/tYideSXye/xJpR+emlESNjR2bn
+WK+SqnINPs3EYUtQ6XkRMAZxjMrPWSc+gvmVy46shATTuaAlqRq8YTh637LljV2
XErA9lnI0CL0l33jFcuwQ23FtiYvjX3x6m+TQcWpciNPtr8wzFagqOJfvH2pkvkp
qmHNXBr0Kn3NhkrEOI0QzWzB3B+/VQM7/ULPtx5nLT2y3jwPL3TvK31b4+JkWfNV
ZnBje7foOEFmX8GLMKX/m8TfId8TGuCxLhA64Ydd2uT7wTYhL5vBLE43tcTk+TyZ
fIC0JCp5POes+fNmOQq2RdyOuS1aJXoVqeUxET+0tU0xrLkmOASor2Ng0vYgJ8TW
KzNXWZpx3HVfB4sl75+gaFGfFZhdwW36d07+LGhawqm7MKykDSkxozZoyb9ZsdPp
O3FkdQdluEEnO5XathapdTkp9zIx4CRuzUG29xVJOA/1R1gYb/OewrDZESVOEDZq
mCldcvAw8w6CGnVeVeAxat978W7d0QVeWgW1p4hVTpmCl38b8afIjF3/fZHLzTdM
+WD2IDjIznlb/H06MbgHbOEbEfhS4uHQrjPnM5IQ96JSEDJ+OrcZQ1pNKXsBFcFw
CyZ2q1O2GZGnRrhYHY4/ZfVKBxQ1xej+v445tRGGOp0mPU8MjLVJEwPPJK+4nygY
OLIDVjtIWQnXAuUF60dyrcTsJsLBGe26HPZXOFX4+h/xdOnKBj6fykQUjMBSrkbG
S4UOfX5nr2RtWBCmXRat+8HVRhRSi/sglEVtSqKabBBC7Q8Ip59s5B483B2Sz2gL
wg8XzCHLACYUzTvPCpClgP9wODA1h65zeNZCzb37EotBznuILXuMubvl/y+irYvr
mq1lSfjHorAr+DKa6c5FNu4EsBvNM6OU9NlYP9tuhknPmvZ0FkYojLJ3gjtMvDzs
jxLOnMq8OpZLL234mKlcZeE3huNPdxQqS1Mde51Mg4WYbMUDA8FwOR8dSMPA+Lge
qVEUTu0MDZ5WvvlCQDgWlobeyDO+9Y3v017fDAbwYJrFVyx1ui3uwT18IwJkXOm7
mtYBlfxir6DyGO9yKXm4WTJZzsHNPJ9E0w43Vb37BnJ+fIp/gIaMmZoj2gZgDh9M
vP1rOh9AXJTFblW81FZ7wFQLuasBHno6HQT9rIK1Icy/fDB/p/H8mgXKCaAXH1Y9
FaLcdHfdJjCSABeQYisCFGZqPk+qVWliM55jA5HlflrB3cFiukEIC9tIX6tU947C
BxaYM9QS4jMoJ3X68aK9KokVbLoPzgSr+V6uj5/VBUgr4Ptcy7ZcrC1qjm0Hezp3
URJ1CaU1I6fj3eGbs7zmhjEbD+xkvmHq4Uju4XRNFB1Kh5RGsS1WOx7Sq2eDLAZn
wd+NJUm10NaD4bJTlVWrcLuCEBXKxjZSv6pltKxIXISAhqSY7wPrQNBTsaNjquhS
n0ZHiH/8XQ4QCx0SeZToFsK5mnBkvtc1mNmlB+lGyVClISgLjFKu0+CWipKdunrP
6lzKgFJAiWtkbowIVNoF/BzTnEzlXPRnQzhwfAPD9wxAfbI4xCf4aicVBOOzazuQ
4ZkxE3F8/YGIvmUiZzEcNxHP9zPflz7hyCeG/cMDOVzJSUeDxWy4JCb3OUYuTwk8
z0HsjzmotiVO9DHBdabYZyNBDh4ugLvk8JnWim1RyXm+byF7bQT/LTwxN/dapLnM
r4rie4vtg9S0kcneU3i2C/OVHzFMtOlzDw9TauBC268GHYGiTpXbQYPA/G+T5KVs
kZHRSN4Gv7OrJXtQpZf5mS3e/gUJPSUlyeLRGKX5VUYWuYv/o7KEBZL1gC/FECWl
laki/TsMBB+ARI7njrIQ2eLYD2zI5Bj04SdkW6rnDQfmklmLnUSZHZAWezC5nirz
abhjT7WN603b6/LyHbsuvPTxhj1xJ0/o/Nsgx9BmJtsU4PKyTyD3Az5Hhq2Bjyty
xk2GD5lHq7QPxGK5O1pxmhx6yN+pTGzFpCFiHcR6/JbkjQLBc9b4/FzwClVICkxR
pvgXd7dgLdGsBy270fgYydh5MszYAn+iNqZkHR4Gy3k89GAbt8uORN2dTRgmXF5n
gN5yV4uTu9ue5N5ZfcgZPQhRalk314PFOAXC5xwuW7OnN06TdmmxK8sfZ9YEsCwU
rpGJGx7rtPK9W8F+FAuiR/f6RrQhtxAnc0no2mhsGgCtV0SXJcFz5uiRywK0lp7n
UdmpDNWy6iUWyRr1BqgNYdw9d8ixUCvd7SH0iYf7Hf+p0WPfcVoKgcpV70EjqoK7
W70ZNpt5PcomjtkqW/dmHMs/1PO9B1LooxRugjBo6eNyRYtAr+acr9SeCDjaR16r
De3fYGgm++GUdw1DcXnI+lCZG4phROFYKIufriHUzEG+xiur8jkoR4kwQvc06Dc9
P9ppDwvqwzZtzjzYTan3iNiqePtlf6FTglxP1SCJM6x7ZUNIE4givzaF+IOhhaTz
F4OuDXFzLF1ejrSgtQ6I36YgzacPBWeyWKZ9BoRKAuGjIiBZFL5t2ya8k8zZfsu8
orFSVi6NRcFo/QrqMPps47FwomUzl36JDRVYJxjCMfWdIOOcECXlnU14zmyQcx9D
1qYGEGN5vU/VbcF4gXmg/kWRwto6HCqOoSyxNjdHNV875pSS7CllxyT9blmVrNrG
6q4XHnIsDl9/f1WmD8Tr8Uizhgk+P5vqgCcwr4jnfCoJli2j9VtnnPXfNUX+Q5vn
chp9xMSPEcHt0EbQY+pZwJnEZj1DKCnE2z+P9mXVLUVygmDV1bFuDT8dWAvo2IcG
cEELLqvSRtdygInSOmjJvZW3UF3xE1r+OMBQwN8Mn19UIzkrx3gPstZv3mAK23+S
8VhjF47CwrdMlxduKVe7NomuX/pW/JMCE3hjNEL9DS+4ej/S9co+0HaSk6mLLT+s
lQRuNjsqlGMaJI0WCWDgPM36ERKac/fp/98BqJebLIYpv1Yk10Bsq4NgFNvXNkFO
RlpMVPrt+vFRLbTpj/DMM+FtGCmVe3LRwC+k1AabQPwlXNIsQVeTMvj7qvmQpK4X
dhuhsS1Bi2V0pSY8cU+5/G1oV7Xhw8VQM6lDd+H/t8AOH/T2QSwLohdOo/ynUkFq
TJpTo4YLc0ox1EpxKy/8DLFBlReYASkqXJqIhnkUjT9fdD0WEoRBnb+L4V/OibFX
LT5H8D9/z+BhmbCEUkaHk0e2FdV0IUubw/b1ggaGECyGJfCV0dp/yFZ2746mFbGr
iqHP7YIOkS85QkQK/WCLPsgw4pAW+hoVMSoiaUJ7dUVNhr4tMmsIlZleVs7HSGTd
Fiz8/u3mm3oeCPbNa03dAiuPC5zao+BjJBMaoLZWHLovOd5KqRpBXObOdTq88YAV
0jAJSDYWCOYvzO2iADWbpCwoAfucAp7m6WBl4ocNxQ0H51nXlk81mzGIFu3Twx/m
sgQIgmax4R0NtVdqCSIV7MMs/aWFPTjgOyak4Ruv/C0+N5PSPxZmbkqzp1RdQv0v
+0ctOeqzeKxAhrkyq2c0qofK/Dh+xvTtvszoXGhg89sYNXuyG21xr1WN+SSj3Bea
m6qiGDyC+Z1nJ9m8odeRhYQCmIXBYyT0X5xnV3/vZMmfJ7M1AjI6ADNE8zQt8r5S
YKpXFVIm6Tusp3Ku6hTLjQjY0Dd9r+LA3biO1e/vr/5If18+3uwEI8K5HZlfsY7P
YwUtwLODKRyjU7M2fQNw49WqhXfftXAweQCsXkHURo76RoyaWM02rumc6s7n37GI
dRg/wnx3FwaSnUVSxssWeALA9zJoelNymsWHNFJZ7lGK7GBOMaDLXzsKSFpviYRg
I1OVyxWnVLwP/Ih69zGwW8HmiO/R2vpKSvVfPxDP1qhrGi6Pn5SnvMNExjXo2BIp
VD/44M1vxJV1rutHSfBnjjFLbE/h0eK9v2W0ewKz4xWIBxNV6tGIAI9XHLtP3bsM
2zAMxg21Af2Jn6xrZySQ1RHE+GWeAbJvWYJP/BgcX+GfTwkYipPX+p2RPTfx2Weo
wpw1iOLn9iBrfEVyZmjNUZ+4F0d2Dwbgs/HxRyEJtTg3e40XqvLaPG4Kn52+sDWA
KsTxhsiF2tt89iM8Tn2/TMms6EjSNRFWW33CBNgg3wkWI4/gSKLTUoHKs5h+qtjX
7V1aN5QwPdWVySMBNrknDWdfP2qCce5iYFxE4ZL2+rEl7RUz6VQUDgRNReUD6aXB
+5mW0UqV2gpyAqdSHBvGkKh47ffm7Nojv08XWj6JszINGoHamOLtKP3lyI8gvsnd
qntWkRAaNa3KQfhot0u7k0+QifIbfmDaF3cipCYvs+EiHr1674BndYwwUPOIdpph
ptO/RoIH4XggajVC0QsBAMLyWz0rhMBqZ1GcDKDps3Mj0LAP+q0MouR+WQy4L70Z
rcwIWFwZOuJxNzW80JK0pleY/F1qtTftxW3LTSxOWCJDT74eklA6rOzIvDd3AVui
bVB1pEM70feghVXmlBPlDt1nbhSRCqirTyJZAOr7aP1CxaDDEpyBMhjpCi1TtZts
M84uIXds1tf1hKNkC+89e7SFLa51Pmh2ftBRpe78fCIc3P0kSrBObxdoUrsrV4Tf
/jysxK0UmSrx7C6wPrwP4YhT/PrPX7I07lJr5aXOs1aR3Iwir35GQIuHJNKiR813
pdMYo977p9Vw+iQnxZk5FmzUeg+YjBKLrNy/xOdPP/IWM63WY1cFoXAjITi1Xisy
4hDBt8DYyL04ZFs3pG/iv6OETEVKlkpdgvY0hQS8rQY1Q8NuVJay2jqL5IiYLSoH
zNKGsIlP4OynH9qs1A0afhJJ9EZ5wYC0U8d1kkpMN72b7AdAugqw/uT6dAXpgMP2
vD3zIxTNaAO786TBrH42GoPUWfyLNhuBa2iFoTXTl/cLV/+jlNQC15G+YwvvvjxV
BweIvtG8CjkqXCMNzuMj0QHejY8qH93QZeOJm31p543i6Mg+BCy0knOQYi7jxF9o
gxhvLD4KAsDjG58BHbiKqACvLUqtyDk3AcK2p5jDnymovRTaLwSfCzHxNjgq4BWE
zrt8Lhiv8u7n+B2ofQAzzzRbg4fvWkPXn21iu4DrUb6UzlOHoFppigLc+Ep0ezbk
QDHCU8bVENguLgymFz+ItqYJ1wpOg4XR78G026csboXq2huEQL3W+Q7UlESDxru7
UODCRGT+sZ+wSNF1w/IMbqcseAl3HMiOWWGewkrYCfVUglVMpDMbtOnI40usG674
ZYdFqMWpaQuFA51lafJqmZVg5VZ2UWdILmgGaJ11Wxr9v5c6AK6hitO4Km8dFiDl
B900sjQ3jBmaiw2xCdl6+Dn+l1CLWqlCvUh10gPILNu7QO/QMJ7YRBhmA72lxxZd
icS4OjrWmYWylJOnjlKNTsnBm98Gasq8CWUIAIRyEkaCUZhx6gQ0oFLbaQzN6Vwd
Pd4VkMZqAIrXcHcfKXljTXr8ennLxN6qM2+uI5a47TvpSkb0KcRbvWdYWhJHWkZf
TVL9fbtAypiVUi8+XhQ13mhrv4UULhDWruNxjtvpBbiIBXu7SMDY6/M8ImK9uiVa
2IcBAFXLTydAPYMAG9jWCKfzdTIcKd0FGIgreuH1yUqzgQZe5Zy+BaDvnpbDMKbi
OhOpYouvstmNbmJX4TGstdaRCR8xWV/Tr30k6CeztqA50QOrHHobT6t5NO0xf/HM
T4qr6zpe7KPk/uJ5/fqUORN2eDKlO5Yl4sWu4qoZiu0dX5DjtVJay6LAB4R8SW5M
wLgnmRsGWBecLJ4gFlk5iZGZd/NkXmDyfnTLhnBGNsf1BHnpUAk2x0L37RWi2Jsw
XW2fXvSuncdfhVtoBftb0RUhPIqjTDzfPnAaLufHBzXKTMxXwgT+VeGrbgqdoX+k
a1INJ/l4VVLBFOg3ZhKkhDKs+HLbTDREN1avhr3pFksPvBnqu55S2AX5V5EB9C67
JXkGEVYUgLxZ90j2i5Udzy9TeWBq2bGBE6UPWfGBdnmoCV1KKw8uzrn0Wlo4PX73
v9H5dwUHJ/eTBAM0fCTPq+6mG1FAMJu/QEj+udKwEuybH3kl0INs6X7Ofy6JWVgw
NImYbz3QEkLQHatpc7rxINSCPAW6JPH82t57OVsWSB5itfnQoAStL1rChSBRNTS3
h8Up9sgDLDu/5fhm9OZ/WGzga+xjvqC0RPpd1fX4Y157OU/x89cD4g2miUVVRecu
DGYaG5txSg4+IHIGCRVf1CTqlE241THIzW9RvTWiZubmS41AhJCcJXmb5fk82sl3
6C3Z+L3Vq9FNqI4FU0zfoFzfGo8vMMSPiAcFuMP38ek5PkNLBYNjv4yRiXmuAtj/
97JUWzTIAyFxjy+azE5tU2Sk8wpXoTypRI+5paOfWHSJiXrGtAzmSh1SaePJK9Ng
TZWU8VVoFxB2dh7XWFxalfbW6Mmun/C4d3EUYMKoaPts5JEcFVbMgWB1ln/DMjEQ
+p8xdcl0Zd/H5hNoMEuy16R558vGZ7PYV5R+offr8D/TYzfIpFuiYcso7++E+Wmv
Smihj+GoQssj/rPzoOtCdu3jDqiuuh5gzo/w+z8jiPCKlitzcH7fWzIk2PTFamD8
eU/ADYsX3qfAAoEgNEEig3KqmypU1viRxdT1+JTkaeI44KqlvRbaQFZ+B74UTWqY
GMBqgvgk+Jz8PBbSLZQeG7BVgAv9FNELDsmrszCW0H03I/KOec1grCNq0SXhmxHN
L8bpI2/WeH0ukQbdi+3G+LLcLNf5AhTNjDyYIZLESS7a+M9YME7HlWHiapeTBHir
ePTXLnOcmaqC0lnCJp+X6huDmEv3fk6FvTlvDG5mQFqPw7dztW2Frj8iP0lrGn6v
dm2Mx0P3N6TGgH5lByjSuBAlTcRQa3JNk+JB/dtdo1mGy1UIaHSQ3diET9SATy0S
iB45/a+JV0setHSqXtLPaBnsrPF6LU7RQD/NazSON9syjJfc1IaYWArbAI4HHkXl
mPxDP41nKWgraVy4WaQpZ0c05RBzlPKAHM8ToccZSPseNIwChfZUui3c9lFLcuxf
U5r5Kzq7Hoy0E2gyhl97PDph+tSFVBpG9iMz2XtRGJyau4a2ljDH/O61V/6/wiSO
sS6+aoKtZvXYcNBgRCYCmO0sev4Ebe2jzh0I36PVWnH+mBVFHIszyBUr5Lc7zxhW
J99yf2N9R8sLeWrVcZcVW2oirQHhbLAU4OYrauTn/6vIsbSJjKJZF63BYzo620JU
blacxQNrUUCbKMDfN17Ylnb6tnzNUtUet8Uj3FEKrzmhEv8IKXegqaqNx6bSacif
t0q0BZ8v5YZ3fe5oB4vUcm+KXF/EeZKFgRugOir/Y2KN11HgNurMbxWuZpK53QTf
h0iwwSWAvpVYQdtOi/b8fppZEFp6eh6LJWW+nTLbFqRbuYSTge+myjZZVe3JO9co
GQiYqVhUDMcuDK8+95nvoXmfx6S/LtOxwzI2FiDfsDPLPKXBqmOd/Dbc3oxtTbdQ
cQEo0t8WOw41SnURG84qYbVzZyq/fmKxtygpLrYKmEmUaBYTmqW58EXAX5mrc0Jg
XW11qARepOq42h7g/DFNo6XNBpJY4RlcMQpVJK4PvGRa0u/7mbgWgyHAmyTPmtQu
/THApx8QbtV+8f/iA/tRuPMcHTODDBy6qVP2/eEo0dSDbNXlH7sadCH3psjsIrud
tGbbS9TllU8USYS0ioZJ/HBbesjYrcWzkjrdTjbghnOM/NIaVNSDC+IddJc8PKTT
Mza6Idpj6p1LEm9/Hv4ZxlJlg+1fnvCFQwNlilGflTjkS4rqVKLHx94tMP0hdfuW
PhjTxhVRnx39B+MYTZ15ytO+UioFn4VzjnKNrnuaHE3ChjfCooXVRceVdsNqCMU5
SnIvldWk5Uaw4pOfI1HdKWn0DoN6M8MmJPH+uvYrC5VRSfWgr0pJxUN22lQTs/jT
G0COyBfCS7SYRGlEuYPyQV2iOSA62Uk1rqSC961iILxK4oO15Fb0MVGhZVatsfZ8
6hSd23zXlIRoLFzb2laqVB85WrfTiTE44qIQ923MWnW75TBVgQAqm+F4Gqs6uSea
3Nx86B563jIyFp41COCaMWhFjjKlPb0LUlGtn2K85WQ+4Ly/abdmT+tmJQvYyoDm
A1vfrp9ie2n6l0RxR8tZchAAKrUF/0+KB3dEJdS6WASD8QUyZu70Lr+DsaFgT678
8zAc5rAz4AAUpDllDUTHx3t80ZzXoBhX1Hoibe2+spIshsMpSg0JLRKinKuh5CnK
1WRCOpEutvMq4pY2n30yGTdu4BB2UEccA6Y2LbYjqWHvwR1sFDTz9/8Wf4Yw4HU2
m3y0ZTgYfPaBfcKdS4nAhqjNsLTwtW7uJIFGqutALz2xw7bEEU+XlnPP0pVNw+79
rE4Z9JO9VewJQrQhzx/YWiBXZxWMyJU0TUnCN7B2knjfSX5noVm0qgROcUZC4yu6
ZzfMw4GH8qUMsMZCg1/+k8hUYAHuvcJ1QqRBLMY/b+gtSj0mA0vbFWw6uqn3RL8/
YfAtMxHF4NqabJxno2+6HLE0o7/3d2HGBqEs4gatsdpszzSc6sYPyXGzX3u3YkOJ
ohQZPkcjj35k+9aSZfSC3nnDYAJOMN6xAfA46HB+aKAxsvIZdMGUO8nihWd/cxVX
BrZtA2FWNB4NL1FItLGm3DK5pSc99L+JVMGieFzNu3DY8cKcqsNKc1h+AHSJmax+
YfAzJ+Rkv+JuMjSMq7LQlBdKWmED5t5qDUi6reKHbEVuhKAlZq3Okbd7lsU7mXrI
LBOEfWwcoIqqznoHRpTgcVe0v0hDehjYBHAUo8VZSSbPR1sN/kjlJjMfosgUnmsA
IgvU38LP8znwdugQb0QZiS3PTA2WN2zmQxNF+9RuYPPVlW8231BZqVVkTyQPCjpC
wKX3VZA+zNu/l2nalXvBjnZTk7ic/zgjN27jXMlOKGcOm8hltvdVUp7Q8bXkpnqQ
ancRCBGNIYzYSSxWU1fpj93RPvdrGFzUtUV9R9Q5Qs/3jj1CpemaSvxhlEUdbxE6
KEb78PWuNWeJxTGpmNXGKexN1nPB5qiW8dDHYnRcsLgR+7vTzK7+EilFSJXZpegk
MHPT/d5KKvNJdb6YDZ5UI9NprhSRW95NAGNh3tc9xO7rZgiRRKGf7b1uVWgZlQlS
Uk1FF+SZU6Puhs8S0tXDvIfSEZAPT/PKN6q6DDNcgOzYzBGH5wqzF8i8F9rCHkN1
x2mn6rIrgWoC11K0DqLMLO/QwIuc1dkd3qoxxFYCPp2TYqbfGYuX5XzQYtJj0Bsh
i9/1+9pTAcMFWGG8cMSrApIGcIm5Cs9e3+RP2NPex6laReFUbp78CrlGVnbTRkFY
NDzz7pxj74d7AKNvkii+xFDbP4Ic8DhTzsD4BJh/m5QReiyrFUsejWzvt9bYlMX8
Sdm1vZYODs8X/f2N43goM8r9PGgX6p+FsbLgpS8BfJ+PNp9j0pHB95OslkX+0Nke
tD0Z5G/EbEDWbOAKEYGFWBenqcuyoAZpDeeja/Reav1lEieH1RmVX2nTVPgV9xaY
mzpHV3klsEXu7qsCl6p6NSZAeQe7sgbYi+OsWIOs6rXDXoxYbxQIkR7fd9XDi5Go
B6VLI03UU7tc390paP/169DAzZYxuNpRl4bpcdCcxtfL9LrzkUPQbKi4sIdlrepD
w0PHElq8iX1ha/a0xroWw83ajnx9V7GVX6IKmLmVpTyciyl/kK35XkBWBAxeY0E6
+V8z1V/2IXgzETmCtX+vGhJ87eMhB+YvHv+q0ptgICBpuOU/Nr2ZZmcxNT0gXBFh
E9lbQDvBkGqyeIbq7yP4M8lMboTugiEKbyLM/zTymb3hYHbvaikouIxXtkwWGnFR
ui2x/ZomUyDQbmlA6EoIxYfJaP7gq7LW2imtL6/Qou04masjELAlml4V3UU37csf
dDzZ2rIfnOlIWwDWG68FNU07cDImgT01ST7UtaAh3swI2yqN1LtYmayg+MrvAOjX
QsdT4CD16mxpGXml/DVrw2PVjqpOjR9zqgn0eeWZW7BZG4ZfHdYaUkqpi54dhBj7
od6TIWmGtSVY5nydoJlwFjNritQDL1jsjEU3JP6zmFsaLd34Jle+Kcu+Y4CP1I6f
KpVp/NQN3H0k8P7G6UHncj1ciHN6jCgjCYppOLulOUdz/pIO2hE+/gkgzpRckyno
ra+AQMFbUd69Ry8m9FVKdmWkh/IXvtaLlsfO/hGLV1TRLvbOeLcXINPBSQ20z6jv
z6UAu+SL9GHSZfYXKLwdURefebrY1Dpi+aSSz90srIo2de+VSFGG5/JbQliiSLmD
ABssAHf90IP9vxgz7ijd8Jg4ZMgYBJF4A3cIiJ86JIn33/EOUD/d6Pwb99GjK3ZM
+KPp8dHg1X0Av0IQog4wIJ96gNC1jpXxnNeZiMB2+en5pAkdBwOA+JUNxHYhNLBW
2mmL5S7SmtQIKr19FT2Hvj3Q3drYJFck53zrUEDNf5YHgGEmTiWlANMiCbjntMVc
vGQCE1qsHl1sLo3wt3gYIIQ5Uat7GVow70LcqPVyJYHD/hleiApM4EnImTHDVoVh
ATCPf4x1yIOsAuO+mbY2EihkUqtMcoaK3HyHUeyveKyAhOSpfcrKrQDklX84TeBi
n/TRhKaqw0nbpkM4GfEu5sC/NDFB7P92o/2NmcXLTTaRB1rcymwvP9MPRDKrAMRm
WPvYp1/+7JCJmqMpY+mDqw52t+PK9qNN2GjCEf5jsLkzzjsLDZLJ+6P3Thkho7+V
bPk4VBv+1OBbpem1C2rZT3/l5h2T2o4745Td5hYXxwK1wbc7ui35KqPTzsP3aRCJ
x055g6rszHGu4ws+fz/BEWBEd1IhO1/N/bs4zHiAxhwrpylES7L/6JcSd/vj0IZs
Hc45CrS/D0NwjO9Hp4o73ZDTUooaWxYPjhwShAufiZO0KznTZsQCSI/Durroz20R
o3bOmEdoqsKtpH1pfLgSBQRnFLbX7NxkXo5rSTDDznG4Ikf9R30LDgS7XRcbapnM
P1YQJtSDFZ0DycF3CE5+8jV6NtLlb+dNwTMFnwkFZQnziH6jcuw/oFrp6bJhFqae
E2RdLXBzPHVKGdNS74lFEPCR7zuzzxFkd4XXdG6KxEaKuQxVfMPStkTE5yJqFClI
YmaVIvhuvx7Uqld3gC8kNRpGx6mrJA37KU6RUtDZQRhZKlZ2ooYy7vn25fwplRHu
wreUPZuoxyavLmvy0fYrylgu3QP5fA5HhDX5V0Ms1t/FPGDeoLVPxd50ba2qKSgm
S0mwZfytts/oVUL6E4KqHT3owQ9ZAva7ahMcaYPiBDkKi13fZGZ/XbjPHRHlQ1fA
X2QgkTMh6Kzr1cbRo7eqVhFf0pCCLcFOWUlJts6lYoJkFMmVvW35oibvLtZS04Gb
eurIUg7TnQ1nGCT5p1k9BSRpXdUBUGbPLuuHX2Q4SyxIgHryYVL+CDP8IY+s7uMn
bfS1tq4pqX56U+V2OoSub3Su+9Ngb/twyAERgBZchlQRpa+//DwiusX7L7VuUfpT
6HaSnabPmvhB3Uuei/uGotNtwo4Am6ga3Xf5zmyqgUcOlzDi8x9ZID8jb+apfZaU
npCZlXYQm1i4igRi9yWZOkBwLSd848YpeC43+z9I8TV5eisP6s6gEArUZH1DFzA9
JRCtWljbMtuAzY+su8DQnV6fYxMwXvzIXpf/6B3E5V+TEGm+f2jQqNCrwJf4JIq7
44orkiEXLszhzHJQGHiXseWyJq1Bnz/zRrx3TCnrN0hYVhw67Ra1Z7ZPahbdup4p
vqAMO5a0YyqjbBA8PGL+jo9jgovS3ot9tfd0XoGID868t1p5qN93/CUAoVQNzKgW
1ViSwYUwJ+YUZx9JIBj4mi7oKnoxKYR5qc39CSkZ2Vsmc88oslnXQ0mymxboTUXa
g+IKpiw8Mo3HAbpxtImXGi2cS1wNbrmSkTEBEWtS5TUV4QN7qRryQ3PsEfsw3KWh
7lHy5woxMjNsFxWI7RO4MpalJtP3sgMxIS04Mg0iRm0YB1QwzdC6MCHXWHYFyPzd
4AiEx3st72ClTA13ofSkCIHtR6YGScLpQ8vsBzgwO965aX5QB+Fh/gZmz69BZS4+
lE1pjGNTES6/PZ121uZxcbAn4+KmcrKiOFszHZQlz9NeKqWKNB9OLL81aeXsCwe8
efSRSb38vm5Sx4U50l2Ft7UoabSMweW7oaR1XFTdr925WMzw2TaTV04fZhqxUam3
YYdDXJoNNJ+UDWluBXnMHfR+Q2wMUlyq0PmcIf88hoXwxQcJ8FZY2WvIIKJurKbw
QChFLuVQWud3JrCnRZeDt+NFDUoXLOwiueOHMFfKXv5cwZqo2/M8I+6qjcyRVM2g
wMIKMGRepbCfyRH3qozeROxiF/f57cRn6da3QjwDBoQWXUQBUemsQuD0yi9dQGbQ
/tOffW9vHCyo1euZUdPUWCrQuvG46M8UxxhxcCnng9oQLWVXU7mQjdWjDe67Dkhg
LmeOqfY4OZugqspk3NQbnIC96P/pQCBG1HMdiv86LfAdO064WY66vUBMdQhWyBSl
AMt7hJdilMctbS1bM91EsEz5l1tqJix5YYbVcUnTDGjE60t/6tvNsY+5GuZ8WF43
x/likBHl5wx+qAdEqI5riX6J6rnS148SbxccpuUGF+8cPQoNJNiZP895m1n3mEkw
pqK4q6LAEsASXjkkhF4p5x4GRuI/EMqQx2D0c9kaz8weMF9CQHsbCNf6tM1qAc8C
Qg0YMYRprsI/XrcCAMjck3/LCyRMTXtLP5SV1tvPD2JHQf9P0QtHJktdjFHYDu7I
bnl4bURWF7MaH+l5s9SRFkwjwWMEf5IeMA9XFUAtlH6bStF5acXwRUH8KYaa16lt
JbN6UTxDQ/XCoRgAdue3Kz5q8V8oMpUJISj1GTrerIxPE2+D7BbBJaSKv70hpJhM
b8Xs3JdvqEJ8Nly2G61m0h+HspP80HGQKSpKB85spfBAc7WpnzO1CP6ehTYdgXA/
+sX3UBBaqnoHAJNfkhk6tPXCDzx4+/slgTzWpOOuVcXfz8+PRBCXhqkLdT1NLX7P
XhFs0NdU+bbeZf/zpe6Wb2PI/7d8RxkBEyAzNIXt+EuumjXH5dQoIG83J8ZbhNCT
AfwwayuSxwXfAAdYlwaV3y+COwzuUOU2BC6cIPFPJoq3dGBXlYhF1gFu6xuQbDf0
//BzB8VIuV74sC2es0CfAwzpP3HuGfB83PYMGw7O2Aep3LGpz0NY6XUasftSqk9N
aAxWaYQJUjBnHC1wlC/7dxfhnqelyU+Qtlh+POZk9hc8V0uvJc0rd+AsLclKVbpl
KtlinNjc9KJSNyRkHtp58NWhOlz+Vp1hNIGzpxAZl+dyc0Mnr/yR+JfuczZWmaKn
WJJc5U1X3CPdh/eYDISFILkXT8dZGQyq1o4rTw5co2O7+/ZAj5Dxjc06GdzMiZk0
tm+Jeba6sgrvcGKRI7tkcnC/b3ua1s8Sd5pUcvULt2QQEvGD0Hbrz3/kM0G09E2u
aovHfu+4IdXmhtQ14QlQ/tS/C+7zRFdBtMvNiwckjnArj6iT9Qine+K3CqjPKeIj
rSosMQj0kbFU3CKfWw1lP+0NILeuzD1ChsEOwxuPZrLY3O0cpamMkaE/K2q34nG7
qIqUSrU7R6dnm0wvcddNCwJauEWK/2CB46i8PfVAXwt5bIhtRu3T/Ow9Nxm1tGXs
BHHym4Y4twiCSXDitixzMgjw1gbo0H7xt2M0xqrlwCQysHtzgsjDaxZyQjGeIA4p
NfyU0POBU5jgJ3Kj8AO7gFr30ONgBjhRuVzOUZNWx/slTiQt/JMwQFWSouVs4MhZ
dYZ6krIfn0N+VjO4AtiQDVDRoCfFZ/Z/lYD9jbDVHxXWisqXatMBP6vyYfD4Yo0k
yQRU8tVsslUcIDHWZHMTD/asmjjIKUc5oVEhQH/TippLn8n8vtEyPTnxB6PAXuow
FY8kXgQIUEZVCYsFhzhj7Gqo1QkhYO7BHZVFynwJeulXEv7w2QBgGjWE2sFpwhjL
ezExF6oS8udIiR/nBXCFovux9UYGsKJ+QHXdbG9OE+hV9iigcq3XTHa3e5j2D8/t
2sEqaf/gfKLZ7AWpOU+mEX/2/mjkD6L/38nk5Cqbl5PvyXyHxCgkNDMIT1bGjfiZ
G868EDPrH7e8cLzoV9b9eDca9mt32RJKTmUbXxwW2ZTl9/loMXF/bCibFBvHgJip
Sg6e1Ww/zDx8HwL/v1flCBj92PArn4Mew3erJFH+ZRL+wXEZtF41/DSLy93pxT7W
/9MxAmLLt18A1x8kRuv73IlKo3p60jMIzSZkDvMXwhONC6WQvhxyJW/ucTR+u9jK
MWH4KwXcoc/fcmmP2S0MOX31OsMc7IfLw9f1Iuf2SVYavfI6mgTp+9Jm+uV0gsXk
PFLluuF3MGE2WG7+FV+zYWst5SQOGrOGyUMutXGsuAFs0jyohTJQUJJ5LJaJEQV/
04XLI6l+y8o/n4ybKWZ/iej4zwf8cHgaCTo4X9cG5aYAsuLff2pp+IG4CQW7es9h
rKwyM2024frF/o/Uqy2HzvED3D/s8zA1Cb2yZcDAUYxPqlidWI0pkwWyWDbuPgmf
RdeFxZw9IBHdGgSSGhBc+A3+4r6wHles/J8GMGlxHhQczjO1Bfz/Ft8tMjnfcQdL
CXpYW4lhEE7fgvxM0ftiZrbscqyEqH1O7QgQEuZW/WVb968g5JAHZdYdt6NH9LCs
I32bGAiBdNiO7HJPyHIPWot59Tac0L2Uc1Ny+5EmIeu0VQvMZURebv0gFmwgdhQH
TpgFanUcq+US9Yc2FJscWjEh/x1lNbdnnJchNOe3S7skV/5XaAz5nTa6FLYK2gME
sw6iiIUu/YzPrf1wK6UOK65XBnhOdYstLz++znEdcgksX5icfCOttfXFvzIOlpmQ
0o9l+tRVHv+nogXwV3VbM6chTmVX+2o31dthqwDQdDatmMVcX+SdK5NxzfGQ9fep
Ek1fIv/6zOxG3VKoSEGhrwLGtkrVZRLGsERdlWRl9VzQxjHmhaD2jcRILNUUDVCf
mRPyhmjJh2paQk+Km8CbMcur9w/HSbLV/vCMEuRy3yShy0Y2LduGDpBxDmv+wPK6
6/3kwrqa1mP/Cy3Fe1fn/N7LetGB8sP5pxOR2KxIoTtmrb7OS00YqyoIvA+g//5Z
VY7semsNQaN9RMsELBHLyf2zUBLUOzgL5UGFI6Z7hbEl15gHmfukddQnPdcCeIc/
VVNDjUNyC0azKfO6v+9MTIJS7BRsd1JWajQFOZC4SIN4DyNwwmnm08xRD5U+wfF1
xQq1Uv8Zx4vJ7yZo2I5LSC5kd21/r13K5zbhDE+TmyU144g5qR5p62K9jHoyrA/i
jMPecUqXTw+Eznau9jZ+McIFw2emcFop3S++Ti05JgxWyBC2csqzDVAEH7x7BpfS
dEhVD9GGL/YWMZFYlJZXMKE7dYVoFcu+fW/EERDr11mbCV7gFZdj6iRBcLKzz/1O
IVjehWWIQ8qT7neHPsv5oL2OUWZeMYkZoklhSyVapdEcbfZSu2gAk+4b9y+7yp2L
aFFKU1x/aj7MliaIN3X8B9LYpWcDIdjoSme/EGPKfUTra2WPUXPqsSSx4yDNShwq
r/e4N1YGQszz5q9YjRL4qFlznvA4fNmRfdp0N4C+QSP2ZlhDDrojjIGC/PetIB2p
SB/md6392gzDg2oCCzOV6RwY7r8Gori5OJww1nIpyPqfrsSdctPHfGAZdj2xM/US
cBTfWwemZJUi8qOx1C9zbuhtoZyWKpjDWXCYtkJKN7c7yZUD40T8/+KeXGvCPXYD
7ASMJQR6xiL/7YXWYgIbo4SXJ2ubCuA5xCPfi/8q9NUeaIEU0zcgIjfcnOZCMMFd
Qjv51evrGNLtEO/CB1OcehL5FSYDH3XJ5pLcIGcrKA/4FKuUSLpsCH/ITHCzK3S9
NX6doyg0REh68xbWe2LhBknLJPAjF84g3Dd1CiZUObS7pI0PQ6bRziu2oaKxZccL
oO0XSm2fmJ8EVMwsobOqugbUkaWQEk7Gaqbs//nTC6kDrprEmcPziN3kzJq29293
rmjnbXlnkCq4kOyBvgVbZ+rVcxmEmyoMi7KsE+ruIe9b8EL7bc81LtSuaQ0hDb4l
z3ewfKQXdbDyFq5dKSltONHt6f7G9jThOqOv/mYCWZFQQb7b70hrUmxEwcURDjhF
nTqeJpQSryvunB3uvcJT5uCRZpKQcd2NTrPhpQ14wgGKCa3eutK1VvUksriKgWBm
QkTw+C619kYfApJxElI1+AI6dPBmmmiFTP3jy3BMdTwL4Bu0q9TdR3rzGvmPZ/gD
WsJDnyUT3IQwuIAIX2Eq1Hr0CeogELjC6Uys5lXW8zsBcjMDxV5vtKunydDgp+Gz
LBYNt/Gl++hvzJpdSeEw5yYby24wFdMYkgvIuC6N7LPKlXT+RU37Nh8myDdg06r9
Se2VGxaqqi7abnrEdaW+dkWiyewrTbfQYBL4Np+gbTFuj6CkKG+jsTfA5KrjhW6V
9QqGQuCAzDo0rc3f2SBvn8ZH+O5rGwr6HuobztNO5fCb/f4/XlVJGYAXZZ5mQ0nM
VoX2EXxQXU1zmBNc7geYCZHpLptE6kgApzYsqaUBzlm20q6wyawr7WRorXVExyG2
iD9IuR3HsIwlE9iAGOxHBxvxtjrsQV5dcZzs3x8wN+G0N3J81kgyWxy9nCLM2vFz
eqAVKq+zwrA/luufir8FY15Lr/xpYWWp6yGZg/X3qP4bOi3a0ncK10evyuFsa2nG
t05YfocJkfrv9CwZg1858Deh7DmAsniGT/Qp/3a4cEfJWJKvXm/A6mk/x04GUZWC
Na1pn2reWOqD4sKEErmXVB0azYvBwKePyt2bkKxAVOV9y70efYBy1WftW+5Bp/bY
sJjf791GYrZJMIcfO9NiggNQkxF4WZ3cof707EUKcR6DhBpc9y/i/aqIXignZPgd
FRsnURX3eNEq8EUSqUcdDx7UyMFRv15cK2DsdeSidYUjl7mxsHbPdL2LRJMdfaYm
KoxxdFdYI85cETHKxUIaXPdQVhy4mS6B99/4houD5n2OofeoyetvgSmSanSxuc87
i9159KrR36wgpB/+EvYug7t4+65nVkjMaAsC/xFmLMdLK2BNMf8ZkOsSav6PYXrD
Uf0i/fSx7AEmOMFhBj519rsc97a0l+VU43PNAJkTJWsBkE//xBhXzTs5NWtb5UHu
Q8id6jHktpM7COWVmYvzjF8PBs2bC5UUAE9E+B5kTIA9LMoR09AzYIoXs4KEMpqQ
USulrNSdtsxTd3Fi18uoMGLzhSFk7bCrIiEVYUJKuXAw77D0ePohi9TkI57IMng9
d66l9h8QhDTGopOTTany7kOZyY1sfjKbYZkiH6f8JvE3+KyGxe5WY9ef2guEr8Wc
s79xxYGS+KFco6qMFBWvkakRs+gKEXGuzxp49MrywL9pM4T2tQeCgRlphxorED8N
NTipoAlLtnNstBOTCFLTRO5NQOBc7/+qwhkD500ywjTjfw1SCJO49PRXFMiH3rw2
w6/LgcTTEe1pwUxL76jTuQpPUWaANRaKbyZeQKcYlPJnfyC1c5rlYtPwTcVZfVaj
ihbcyWsokW9u+if1vrBr3DWKLrpXKC3IFook8F7YvhjwOaFqCscDIqHpRNt5IZ+v
ylI/vohsLqH09YGMOQ40nEnsN1jIGsTfB0VvYGM62fmFZvdbniEh0zDbmWVKWjWM
PXPAJdB2mEh5EY4MB+AcvDd5rMnJZYaJn8cTWj/6/nv8AIlp6r7PahL6oZGzuRS/
S/5RU067l3eESXJ4zl0SGx6V44TLma/1efVpLurJo2I4SCehNCn0wZwzgDzYFom2
dkS1NIyanwJ8H6d6tNOl7WyknUWhqGiXt1KKOcjeLtJMj+7vSDE5TFzfGuiyg/H4
miKRoKL5c514IlIIzGzR6C2RTWOIttjjcFelKJXW+YJ/fvNroZdJHA8WXP5iG/Zx
Vlu5DNK2PgYgyKRQfTEfdcuJBmisBiiKOlEJIbgwSrB0rCfsOsht78nR6dG4D5Fy
kyyc3OndW4bvKCoo7y8Tfhc+M1EDfbTjsTmJrw3KyHnODfveX7rx5IAkQqRPd55B
+C9mM9Jrl/olch3whbqsDahxIw23ueIAMmrQdRjZ6V/aWI+aqDo6tqixdqNIAHMv
ZJLiWTCDivytOgK2NZcjFd3XuxUvpij4pdZKH5DmRyv1xah2cvL015LNxzqefcUd
+a0BHzOArgA5qcPFBAEESryzjRMkdgVhN2/p2GmoOQOKG2tbgTmXTMTc8aqYNjDT
9xtviCZ8u9iehK7OKIcrfrz/WOa9ZgiBJJPVGjvMJt1noQao1Wn2eTu3GTkD05m1
88ANJH02+M/y0oTVESMtNjWzsRXE12d+Ey3LqrPmPP7OvI4KiBY+m62WLuslVZ+Q
y/t7HevlGTZHcG0TbCah3G6gSJ11SsTh7dg83eaDC95avXCZHFE5LLM++RXCk+/z
E+UkhAocT4tVL5Ugau+T1KP1OGqQ+cbXfsLDAsYjniEiePD1d4+Vm+D547Y/tsMZ
8OGZRu9ULhYVLjDfhCZwc8mTLd5BKQXCPbWj3KnY/BBQilp5uqVy3uXkuN3CCEy6
D7kFn3lKLPQj52as1AW0OAOc5dPqYQjhm/9tT1kFXy5aNT547SRUrjjjh7/UmT/o
77FKRfZsSxB/w3J/JZauMOXLb8t1QSFhupYoULtT7U5zPcJJiI6aAw9dCzRsUg8h
eewfUR0p98CLxApU9zAuktkJtIkELsiiPLtmQAilDpefTX+ZhQhzRl30OWhISoUE
E69TVRajT2+kuNmB/D9X7fd05VipRaiNQlaiOxWBMbJPrTBs+DFtUP+7ydrUoWW8
n1XU5EmDiFkaRztdo4hctU6j0U92P6PPpSKSiNsLa8ygQ5sz08XxeZnwlOGqSvXP
k8JzSDFktF3Iwr6p13YDS2i0vy3clhWDg+9eWWL9gkwDb0M2HctWWxQAiSj2U/LS
eb/y21vdxm+htUqJgknqRH7wbd4fjqli62cmx3wiMKAexD4eq0j3kUp0HY7m7wBJ
bn8HrEPfvxP+FExYKdz/TDBqdLnDFCQI6tFV3F2SbsY/syN8Kh7rvmGG7cmFOoNl
rGwiqJdLWHFh7Wbcl4LMV4Z4E0+EUYEvC6UXI8au4qChIgUMEn4R6e6f7kiwb4mp
sE8i079pnjB6komxmDbJuhr0CU2oakYm38Dp10mUAfuzfzEzRK/bqnuxzX5AyTCz
F3Ebs0DSq1fgBaQJKTBLbxc505O5zPf0b+5GcQyOGHJe6+AnGoGvW2Voti9eUvHY
q0WDT0czqF+HP+eIPkSIbgus58aAfD2oATSUszfkexQo6KTg9IRZ3aWBgcSBO5M1
ZlHYwWvVpd4n/vTUvRPWrJ8gbKyLAakdnXpCQrWvbLfVnTeB5CsSdynwyQ9bOmns
A2hFmQriEcqaJ0i95jnE/wGDrm+G45wTQAhQiJ9zV2As2eg5JU0WUwsW3eVLnk2o
l7OlY7mp0wDBtt5Jc4XUC+2p9O4VEOmKw+gAEhBQYRyMIpKUzPimdY12Q3IzEe1a
Ew+xaGAARSyzf4tkyygsPim8OzNTlA543X4k8s9oxUkfOGFvuL4Mocf4I88AZm1r
uLkPC1yQj8Ra/fiGBvQJqn/QiFuyrMCbrpQNhgmbokcMRP/F9bahMOwCIbfNrtT5
2S2Cruvs1dFHdwoHfHjz3WhCheE3geK7NmYznqrv4qrgB3/5wA9y2cV5MURBbRRb
2XoWfkw+F8ke4jVGl3yermY8+u8SxNYqlQ89WwkMWEL5rFoeAMuE+dygGiamTr15
v+/e/E5Ir5zm0rtpSgBbNnxfMk8dcwLCHw1x0XQ3Ec+7s6SIE0Emp/LqiEerAqHX
FzGFPj3d54zFVQgVs65y2rmD7KvRJedGYZ6G7wUuZjQMYWe2zhuWRy7l2cTiJvxo
uSzpB3G/1HdX/o8iq4UhWCCpYJ9SgVug03Mq4gmE5SIdRPVARJDbD1ySgrGyaOKi
QkveGd32isoE99t3zidq/n3Z6botSM0gg9zBNt0exSKkPlSItCby158zKngDi+tL
+/zmr0SBl+051BjWHMmeKB+o0/QGGiVEG3Uo0A+A+3LQCssfJQZ2b2a9EiKS1oLb
6umMVa2bi/a8yiczJfpNoQh6vpYl/4Ph7pGmFWRBuMIJSGXdCSh6drZ16fUVXH6L
ypvtSPsOPizg3OypS/bAhJx+NXDf0ISaccsqfsYwaur1AOSPgrdi6ku+r1lSHXkn
UHW4WQnQ7earuantc/DgoGnopAx3BSL3EOvNpVoIewjGE0dtkQUPmVoEk9vtv4R4
TjAlv/9nl8mmelEQhxdqUwUncIYAJrsiUlKEd16Z4X3vR8wk/OlCDeii4qs+0Uhu
ROLqV3YTbWclq2TkyrawR8Cdj9ZvWh0mMIHT+crP/r+JwD48zLZVLOfrHuSXEDxD
gd/1Yd8djoCHaWX2Gh3FGPvMBJZFBRUF6zI/90q9kKJIks+OG951ALai0b6wMBb2
nbYUvjQdEMNBN3QnYSzz28oUHVN68llpu60mp3nuyUFYf+8zttPiaPicLwoVFrfZ
SE1rZpT5LmOpj0BuVqpnBmjfQ2zO18hiIsPwdDzL85RW+XUJYeJUmPIA05ziyHV+
0oXHVWxalND5+OczbD+E+GfgsKqkth7DineFNO+JFxqSfiWqlZ1DfrWgqYU37WIK
TnCNdbi+yxlRnxcnkE3E9jgZDV7gxOQgSLNH0z8kWML/bgHvJ0LAPUzsPXWSOkjQ
Wlv+c+c5sQDJeWaBIw5eTIHkECyOl8IfwrHOQUPFyHldFfDjvbLAFbpc6q86dMVe
zFCDdOc5PFCc9aqIoHFgZkDhGAuge8PmndCV9zdG4XAeTr0tk4OrAQu5vjmQJG+G
J578ISPeXwvqhvkd5ldZvMQDt429aEZYgY7QY0e4IuqLC5Orc5rT6xUp6NfFAuwm
73EEsjX4ostPQGOPJ6c2Op1iaGvPgG6jJG3NlBBXe+KRnGU7KOBC+n3W03YPek+Z
OfHgtf4FptdthT6/JTuCib7gIzCKEFhF6rgxh/n2HfmVmIizXcLmiQQoHnExZIob
k2m+3Bz6jMq01CnBRi8GpJ/Zy2XCN6azW50ZLfXRBhPN+EU3LdHR/zQBWepNYFON
dAQTqk5WF9/myg0ObY/Fs/tTgCcR8doZDin1gwIiGj60JKFe/+jZ5mn3jFBMDd++
AQg3zXW73/FsBGBJpALpen+Suh7kz6PQ0D3OfdI6pfs/9LzRG3ag72sFg19U+4V2
atsgRRVyHU0yfwPfMbqxRnkJb7bW2IoSQApq1YBAQiqXeU8MdpDYgLigrsPSgHsj
SdHYb0Dfjh9VFv0ooO57ZdCXuQ7bdVkDZ1cqtqn+H36Bya8zcL5MtYW7onGq6QIZ
+xzUdhtJaS5BbQPOy9fW70eJQh2fJMgpHa5QisZEIz+fMIDDv5vi4QnOt55oW04B
jDcUUbfx2gFDlUvkFIRAeOksAn/zy3SCleKaUTRaFRbzybfNNno/img1mGiH2GDx
eW+DvZlQiCuLzQp9/V8ndy9B77Wffv02XtDbawTh7b8+ROTfJhxt+Vr7KKc5WSqr
mpPfFgoNX61zaaxK3BNQ6XdPaVG/JRMd1NBvHjIAjovVw3f7NgczG+9XySzJQzHY
3dIlU+5GSUzRRtYTnJxMmupfyLA2fQrkNGURDyWsp94FK1kk3Sls+PYfHjHQJFk4
vczIhAGkc7xwpGjExeBGcdsGE1TDHSdTbl2LXlgk0sNWgl7QsWMS9J59JIhvsvXL
SMXD9Tb/1WJ/ktsS5bR4vydH5ZfGKnx8u8gvucys9J0HwCe/WtufS89Hgl41upI/
SgHJ8SxVZzUeoIgvCeKE3erB/PBAUekz8fUdjpjBhqlpeDTQYg8ZAn7/Uvzt9mPh
Aa44a9IjXjg9+3mKwgGZ+8d+nAhTPuQU61cZp/Z8IWc5Jf6stlkSdGLEs5VhQWOv
WWQFHXEjMu7J/+bFmJsTUSaIdaKV7w5yEOVR4cZlUIIdI9rc3SLx/k5hhQjN0jMo
bZH4/U9IwH43T5KbFzmwW5Mr87iN5gKMQ4pyoFLSzig4v//iia2/1IGoIkhUgEHc
AOYrOeNIdaYSeiaptR+jVLABaLOFsuP6eAdJCrxyujyKk04mXb+sp+ojhZ0J3LKd
Pd+RkESTrVBjdVl/78620oUc/8GY4ndxQPIef0RtxoW3irVDppISnCDylW+cC87g
Z0vA8F3XumYG5HaRJ4uRy26Y2Sw7WZMGohm7kVRAoIlEJCAJl9jc9Y7LTcPTVI98
MFi8kiE9EshzwJ56DQc3PZD+cpvdOH9HZy6adbdnmXzDcMJ1Asj0LINo0ua+/m4+
j8l7wRn6q3m3bqTsrX9zupg2f3l+XVoNuiwniFnTj1yndLlvGsVo4j60wRyD0cjf
PNy9PJgGZoOeoJ9vYgyiLSYHd8Wp6dVcEee8w2Wnwh8cJgOlPNKSxbmDYGSq92fC
BTXnQuSzCYYULpOdGNgc+pET6v+hmfq5EX0/f10FV3OubCGAuFDmc9Jiv5QQhUVN
JMpqf8okVfzjt84XctAAMkFvvQk4AigMxti26napDy9I8MOZVPkHTBesPTGVoke4
C9QtVWq/hjLhfFDMMiPy2IV+6JWAQPmAqLNvRKyxmF/BjiLCHDEYZKDiG2mbcBf0
4f8wpgqsEisbhNp48qigAtcURlrQxBqdprguY7lMxSTJIEXofhplh2G87IJ8DDg2
2t2M/pyh7gFOmA3qtnuK8szKqkKolIl50W4QQr50Zu6spFaY76O+AFxwcctZZCsI
qFvMS303DeXCoA+celpqclI4YDeInaaM3Fez+kPSFSZKi34y/AyMeyX7WhW3fWWw
FaxrmztAEkQO3WLIlmf10JyJLZXlViMZ0yAZBVEg7n/x1mFOzoowad585pLAnEae
4VOQ/yh9CjRQlcSQ2X9wpACJC22kChiAx7+1bdEnfQxoWDDeM6ESkCkUrJPokbWM
OlVP6dnwi/C6Lvg02eDfcROY45hUdvfuD/abUEG5TyZwqlBGZmk1ZWizej7hXdjf
DLZi/IP2mytVexLXKEPPUa5xtVJMf8FRk8auucFXBffvfJSsYshyZAmrA01iEx2b
LA+Zs/d/wfSlBmS70WMScQjRUsEUc/uVBhfIPO/Cj6JAiCjMJqsQ1tOqb5xa+8dJ
MjV89/TENuW7AgzqB/+h4bkpVuQ63qr4Ewq/ABG6bV9tBZODWtUgkgueDuWhiXU8
4Ghu5+IietR0iZuMtj9/YC7GIEW2dQTsR9qGoqs5pmnmVACR8A9+pikW6DdDYWsY
n6X5alAl2wWcHlOTah2cZP688i36jPPoHALqoPXYSLyv5+2Se6b9dlYFodq7UcOi
qIzhlxG2LBAuNsFOb2sP1Ku09psvm54KETo5Sz8nEh39LXgKPVEUVB2CiH7OssID
ysqS3AUcj1+biehLeGIJsrxpfm10WKPxnveTpngLK86AUAPTkpRmMkDepxSTqsDS
bxDS8HCI4FpGoM8sgWGeJmqt9DQg2htzuxGuS6I2LqL7bJage6gB0DLOhjKt6Tu8
05FuvDYO36Q3Lu+zeFyh5fup/Uo++z1AIXJy7JZexlri9OWz3ko3QPXQL0HRgHCi
spa6/6J7zhWgRxL2AkpXByur+4OovAVW5ReE4y0mBzDicqE1cBmRm0VO1+1fvDKd
wbGr4TvsFLtaqwZv8V6UXUmmw2lFNytAxbLCk3XJ4FAtIGBkAko+k1CwXsCJ8CuD
QoN3wgSPy9tTcsiYdFl6c2V86fE3/3WxOeio6SrKPkuaOZ7jOlMmUzyIoCONkG9O
JAvFTcTHalBaha+ZBJ6ufh5y0L+Rux/n611Z6qal081KQPq1XRMvZGkRw77Ec4nn
4zqwvXLyx+fjImTeLbUyIW4u24djM9DP4Icyklz41mvBXlJG6a4+7OHkz70D+fEr
8ZjXoIT/y+gPOh3KxXoYQiqWb/BoZutuLQe7Wv5j3FAK9tO9jdr5QZSprUqkufie
eBQsWkDsmWL16dFn2mD2FJRDyfpvURZ0QcrZYm2xLkeoj0eJtr86fmDTCwhfUsxm
PNaEXWLPxj845Cz0CWV8PYMT7wFqH4u1ih2r79mxiJeB2d2nB8Endieq/2tQwDHm
tHUH5fqsBsKL272BCq+SO40iijgmvrKh9K/BAgxlzI+iQD1tGkywZ3i+aFXw0y8g
JpDpjvgu/LPe+ssB0IyfPbpE5oPSwNlo+MWaLEqCuYHEWNF4yAdzoRYGVHg+VqT2
aOLU9jocZg67yB3Wcv06MM/xGhwegQ9TqnQobvCLP/ZjfU4mYIC+Q1d72Ft257ui
HV1NILzO++EJCP2cNgymFkL8NOPI2DvKvYBzbh3uAqBugZljqGetfgavAut4G1G2
mJUYvVkjRQZRZ+6wluoBnsmGg/okTov2WU/fuvam9dVuI8MzK0iQqDmk2bn8Ogzj
FxB+0rmGt3jmYPIl/E+B/znUnK7bTkf5H+adg5A/R0/Vj/jMSTyt7CBuPr+aq2Ow
swbkgnEVAfUIoylwF7kYnGp8kPUiYjJTwFpHvUv1xKG5SPcO75wMHuec9LMa2D/V
nS9HykZdTn0qT/AGC/uCkRo+FiII+0YryXttwguQm4OvY3ZYi6snkexcCO8Vnjrk
3Dzr5VMS0SnFWAbiiKg8DeT0aDdL7YyfYNrURKDX89M1naAq2TuF0N4ejoVSk8eQ
UXHS1qwl9KfkQn+bdmdjoalzcVGFBP1vnplD1wzWmA/JzHsNKVbXp6w7fy2HAz+N
Q19wDx9SvhxujlfEaJ7JjLO17UpHZvCWyQ+LDEfTsQSu5jV4GZ/xNFlZzZU4Mxiu
jljRJzz0yvhqvCn3oJON946Prmf6CjxXxKmGoSoirkv0//0Mv0WuUowwkATGith7
gpmApteBjBC3rvqhK3bo8ejtfXTiF67oDBS2aqHM18qloUezkRw2kxbc/RkADuCG
WtX9Fox3X+oMzlD/ur5NLwwhhOE0PaptLlZ1EH1/CE8NhcaKKiKzQwnyxKYYrtI9
7s69A/jW2XXQJW56KL/XCtBOehqmtPtiJFBmuNCbHaFLq8MWZXLKgOuOx2OQy897
qaaufQ1sd13yM89klJ4etn45LQ0gEJM522nr6u9ZvaMa2VUOG5GajvOjGdiLErAz
YHxWxaDRAkXkjImORPFuZRGyaNM9pBy6n8SOkWXwHUPizeXd8/xo3sR78h0WIwBW
M3+Bfi6USc1RP8rMG0o8TjOZMMtGhQGb/BoqQ3iwEcq/YfuE4OYepTyYkmKPVZt/
yqUx/k5SmpFdVk0H5bUSkMjiBzyantMCD1RAsFu8IZjQ4k8ywmrTyQViEVjaQqtc
knRGQVwyq7KEoKUJ1BxbO6EAjAGwPRE8w8VPCheshGP/qrBaoFW+O2lOJBVy5Gms
mLVXJtfeJBVFByHz5oKu+rdFCHXuC2inQX9wa3/Q35q49YDPXzNLzoGpbhoky48K
c0KiEbKJP5tFyTFTO7NzPYjitW2/zLkmY/VCuaXcwi0etyIomQkAA+Dgt6wlAsgx
eudPHrFsf2dF0RbgdzTk96pYt+6uJEuLDjDUyBCcCC4qm94CsNb0ZO4nt+i9srzd
8eq5NYxCyvHsOxoesUyaoCVun8EO9MdoTw8oLG3BTVmxffK/nDbsL1iuyFt89sM5
ezAdrN4RW3lbSL0Df0hKi3H1VBWtKjzfb2ftUbD0cXoja9Ky9c+3WZPdr0n7RzGf
1fN7qVgByrohAEtnmJ7TQZW39sWHmSz8z9jEgFiJv0TsOeHK4QaFY5ivv0Bq5pfk
q8jPMGmkqFWDiuhxG58fXUcxgCJ7YNQ86aPuIPUdkB2KixbiMcR/xdEZ/fWeXlbr
6ESQmevgdUCDJ6BCgtDnIqdeR1+PsQKUSMtV8begAM++Wb8KzPfZO/AMjM0tJalJ
SqtM/Du1MJMvOb5eMrPGWEUHm68iyICPXL+PlPcX5SFcdrM7vspRuhus0QeZi6JB
0Yc2ezeYxQcCExEbOI2FHBnfL2vktL0LxF2R8PProFENyBHCMAeN5pN8FpeLxj5B
RwiVToD1E3GAvcCPG2Xkhjb4ZGETAFC6YZXCpRQ9hCR9cuMd5WZ4GvHbdvmGEMQx
1vQ6sYTFO0ZIs2/HF0w1r4RXRrreob8GX1AIJdctEgLJW9fZnUpJVBRwWa4N4cjG
yDNHl3EfyjuoLwmZ9uHS8fjayvPkW2EpZdDJS05szcTa9xv7o6ppEDFSoDe98d2W
ni4A/WVDfWSyBKw9SMNGRUdhorfOBXc7m4M2oPt0wAGKVzUZxan9nLWIxS4n17VB
8fPCQo+5odALOcXcE+H6Wxa+7fWzd0rGrMI2IfNAPtzSX3aPAoUfTX6OiqkJEQW/
hFl1bVZ6WJ+wcwTGM9NUVJoPTMNzoxOkzlfbNduyfqddphZbjMt8rtOr9Qno1ilO
AcEHLakj1O4VzXeo0GeuQkpdkP2deZJ935ouaEIyqaP13JxSdsZMJXy+oNkXnHBc
9q3EIrdcpkkqVJ5vg2Y1l3FCzML91aHE2/a4ZSmaV4qQRLQ+P1XhAL8p1h0WtZi+
3cu6jX4wc3J51wQNqb7wGGRV+mx+3LjE3ceNiuI4HGM3mMErmgX653tGW9d2slXz
Qvrc6FFMXHd4gaUTmGlZ3moSaS6fgKVoBMlMSo2+F/tJpvdresNkCNl0M8EMg0Az
ol70feIZGVtzD9onm6cf7U6TSUph4cmbqjSxJIMSO/RGnjWTKmjPsvkMMRb8cj/w
pFCQrbZEeg50W7l1R70lmdvn1e/9p+j0pt5jIibInIZKPhc+7hbnUZrNQSl8OfGS
qcQvsWH+eP4g1amBndi9lGngwp9ju87GuM8yIByzmCAtB+wWXcv4iyVMWT0IiFbk
QdRaZRwqEeJuaXH1nnUlQY/XtENOBMQGrc+w0FX86L8j5bKqtEnM4DpJkVzSnbhh
X0EXtQ0ybPh6VjLodDP2+kM10bPcUcYW0VY6e/6Dlmp5F91kv4utyDcnpKX3hMn9
htl3VHVh8tuEK/+AQ/fuCZdcQZAJNfkEBirXEVwZus1fLmrrvjCvzquugazzovId
6zbheyTfYjNRK8I/ngrfjO6CTOJSV0O78uQzfC9SKwBLafpvTEA29uo2vzU+wSZS
VujOWrYZSX1204A3Bg2nWwXmSEEStA+6Y6d/wuebjmgLg9dfZSrNYGnT174BfNQz
wXmKf1p2Opo7+JGmvrC7HkDNgQ/F8LMstziBVeo65fKuIC2hH9Y1X2PrveY1l20A
oY5Qss2DaJ7yWSOQJyhP9tNVgQxBxvaUxEQd+097bChU+rJX3XnvzXnDDWTIpOIq
juXAFzVlm3hbpQIHwcO3iS/pRUv/eqnqFglZri4JN+re50fZCs9yzk6D9Iid/9fF
qWXs4lKiufv/cuHvSuBiDN3hBKRb6V/ha2WXFu3bhOiarnQgNINvfJuM5QX1zClb
Gr9wkwtIJf6qisqMSRtzLws42+t5J+mEIwCVLxS9/cotKC4eUSjHhCwQGTE/dWs6
lMqGw4D32Wk/t7I4LLJByk7cqwJrNOYq8mFi31++XxbHHkjxqAjMGUSojxUSRC/7
qIxuSyGU/aw0E2n6bzfB1RyBqWtdG9bnxr/vltSRiUHVp4wNtE5GTmfYChqs9Qn6
xqPndyqUzxUbAO22xACW0hHdbiGortq/3RKjYr6x91HkVhmZYyi9pZOZHP+Da+6d
TRk2nlnFW7KcuSHbrP+tT8JWOn0U3krn26//NedKDVgtxo1ze/Tib/j04uve4g25
pdD1SJnnUXW/oIcVHyAbcStIlFTeJmCNAnHVqQ3KtBsSpvfTlfhgvMSSSmhO4rr+
KudivE7JiKHmMyIQopSl2YW3i6UWhSoA22CoHZ1OVnQMqE/DzTfZAfiYua+TLtTw
F4A8WyZIPBeTf4mUEpJKBdy5k94GUL4DWGg9OLruWjjFfZpq5IG2h++M8WeGru0n
GxTWXgouRQ70vPDQ/6qKhIiTek/Z8gkUBbiLGJ2Dmn606xS08UATKc0h5V9DQU1d
gDFJv8ctnkZy2EgAh6UlxLr96bZQmPxpdcdRQm6Bvi06EWo3Wkj5Bd3eQbB8aXPf
4J3jklkaqEWfdx0kaa44BUhkQWQMkRSH0EC9ttUohE9th+8CAxSgz1d7c04HaUKp
dD0smVZBc869sDer9S1LqPckuD6JDHAxGqqmO1MBJ821XNGKkgHFjY3WkYTIfcoM
forYIciPet51l/+PgYjCPhpCDaehVxNCnPpyrZiLKeOB4QE6N8XPV7w5Ang4oYZS
l9HSnK078baiJTeROdi1JyT+I9/J5xGOwYU+gwwvGhAPal0HA7ogk5Eguh9h/mNp
mM2uXTRbkb4BuqrnVujCE4U6ua9akNshuCvY2bpBJ6Lnil4W2DfEJStf0+pDHus7
6e0WBMXvN9DDm3U0YwGDYbNGLMCAVYl1VS/zb5UBnwT7ETr/F68Dau3hm/ko+jMK
GmVObdBBxxdGsNQkPdLU+jEnRQZfPq4sC4f9Ug83yYtJlrDSNfhjxuvxZ5HBBHam
vGGhhlN0VXLpeeVQCCvm8CoGS3IoaSQTAFfQMOwYezImwuXeMSlzOnMkMR7TGlRG
LNba6qNvw3YXxMhqYWSS3s1L7QGRzAIN/4+SB07mslaMRXeYL1pMHn+j4XeCEbH6
++gU2oNJRV1hRSyqmYtzzUFz543V0v4q8OH2LNYx5qJwuD/QP1n8FyP0oupSJG0k
vLk90mHvlfsBorH9c8vtexeKcTVO4URwwIeNRNYwqYMH2O1mfwVSGIBl4/kNu3Vf
0RMM+OLVBffnEG2mwf4PaJh9+6bftYGwmWSF2Oi70Cd74dZO0sc40hdntrO17UX4
eU3UZ2VFBdS1O4iJO2u50GYkLN/8zTgDKJNBN5gXmGdWbzuBX8H4OFSEJ4xMnXK3
j7DJXZSiDNOCIOMxHLxuuASrHZf1QPZWZPeczg5nj5BKGkd2OivftvVrrdsI8rPA
YZSHMWhoba+F0zSXKR+p2eLxMdfdtsgJWxjzM7yIUmbBEe2SE55w+PDmkJxEm9yy
Gv5yefxbmnstyyCndkI+jGWrmNd5IdrU+y3NjSlgrLPZuXpf+ewYEFkKWBOmHOMJ
TGnYECLAasN4pXnZWwhEKwCCeLn6l8vM4A2h2ESiZc7kaX/lZf4hXyxuEVMMEWOU
j9xywOfD0LXtx1WjNYOUwqhux/titibWgUUXZ3NcdryWIO4UF/bI0as3ScZV/gs3
ElWehP+UIuDv/Dpcs9Xu7iBLd0GCXHTQ84j67/qimtqOE8TRBRXT8n6aii/DAt0l
I6kFrCYBQa6YRdmv0dDXCyOJCAODfkivAdUd5CzWSshBlga/upk509W769ND1fFZ
+3xscJ65BfGadAJT54nGda1cg0N53Rc7qpFI7bXs5qEI7QFYjo3dcHRzYBTftgtg
kUS7snX/G0lOpSvlHU/GdrsgqIaxlfyN0d+bOIzXqX17iHXTi01bULPMbhJ6Wopa
hz0NydACyJYrNeBsiro9us9XSIWBp6kFMsGNREXcpIwsLzUEdxg001gAO0p8B3Fj
kSHNSuCiNNSf5XHiZBOGHQrWYxdHq9jSGOlqmqTIXsSNszBMx6GUo3cKfxLWbL0O
iGuqfBBWuTnhKkH3piNzo3U+d8L1U6NZmMuxPXh31gYjNxb+5OgHGXOOIbx6qtBD
p8yY2YO2+ANS/kjf7rtVecHeY5pJdByEcG2zXRNnmtQQDSm5N3WuwGUnWtklRYIT
Ry+9cMbMJhHBInX/gBNove5FrvYiiyW5ikyCqRjwWOQRuQQiFfUcVT/dl4VfxZ+v
yWeTQ4iYYwsYO8PnfFJy1V1diXgXyPMK+lA691Dhfa49FATLcoDoK+6Gw2wj6h8I
cf/EKeBpWKsIvt7ZXieE/SI9oDZtYFcYuhwU0FlXGCA2XF4VitIo7z6wbTQZ2lNQ
v5vs72tGJSy5FagEB/u99oMH/HXSxuswA/CeIwkoGWLEkCIX35ElWUxBx1Oin7Y9
F5kUbXWR0fokkiEoM19N94o2WMSk8yTXYcJ8BeS1xWBEnN97i1Brphp8dmdMGUeu
rJzzzYHEE4ypwDo/Zc1Eb5kFpZXLtxblqlhXFWf0Eefft1ltTZDWtSJvtMJ72BEu
FyxJxUmT1WKFAAuIonC6g3PVlykU+t5NdDKs9UPtKDYS3x/nEPjrPMUqiFVpnqzU
cyXbqlR1jAhNNhulraijNayey9R09d5UeXQv8f0grsPUlXRKHzJ3GBJxRJNM5uLo
W+CxOXC5HDTZIyCw6nDid7TbEykT8PJlsT62zZH5IWEq9M++BVYtaFaQXMCH9Djc
EX9ZxClkUTcavsmX4QtGeJr87d+VR56OA0eeKVg/bK1840FVBT3+N1X2P2RMx9EA
n+Z0XvWTsKdnyi1Qjemule+pDeEM7Rdmd2uoHeeOCvIiz0Ef2qC5oOqm/Ro+eKsb
ccS1u1LHXJ4DWfRKQRvfoCpMxzlPva+VxdRlHO4hdZsCcsOJyfhWhNTQWtAXRHGl
erspEnQvOgehXEop/cu0Cq//SPGtL6oBx17HeBLZvA8/twr/waAUNYx2o50LYA3e
s6341g8faDDag6unMaMsbH4d+JVP/WcyxeRFcdxH2Z8RUoy8j+hVVBzclAxkV9Ed
vC8PiHGZsjk10SEbhwX8PCMKfBf1N7Lk6a36JNl39MWRJrvrcBl+yOOt4dLEteP5
Ie1NrdoDANMuH7H79Sh+q3D34EP6iqyOBpG1NR1T+CxrSlsI37sWgXQCGKuNyDO6
AaQegtuC3rxTyPDrdy6VicAs4P4J/YCtfwx9SyQIkkpuwJY5Swppoa3DzYEb1A9w
A0bMQZFIs4khCDXJrMsCY1w0vhOC5BNhTHDQ5KWA75mdp+rQMkuHxUnA091BE7a7
83E1WSsQ+UMwy3bTHyPLly0FFm5dMVH6NHotu/8Pr6DGWRf2Oc6L9XbvAKxRR1HR
qvOX0ssdVJzPWe5HzqEk4tpnRs1KlaHKZH/+buYechvYDfY1gV48JXGZ6XAtvOgs
H3gYmu/cnyDr19cE+8pCbcqPE1ux/QgxQoAPgZvlo2LJeXhXOZV9qCqVNA3Zz3j9
kLKSBaJVAy8DE+x/iHPOwPo8d6dT4UZJ1qeSZb7rzjXvhy3ZChDIGFEceL1mjSUu
pDh2yDpAXXM/2Ce7BvoYQFZCpBPmE1FGMeQacEhf/Smq3XcccxXolCorXLmMdS3y
44w3esA8QCG4gS6LvFjBfqnWNyWDWifqDtkiHWfKAS8Vqz00jkug3qdeI3hz6hSj
Gcv7fQ5JEtaeo2ApjEDUoACkGIEaukwhSMfdQ40SyQdlI5WqjQfZ3oNdD5BCyNoT
fSwLkctEGItQqeEE1blFhcmlQVbZkC9R/YNC3oNuFTXrE5cw0VXHXK2q7VWPZiDJ
G0o2rcBeB/fyr9C2NIT8EAnkUHyAxT+XCb85O6ZM9xRd9ywRlg3M6zZSwr2pbGp1
fwgAWcNdoCJhb7yZeY2QjE+VU772lJ2Pcu4Twbx4U7EuCpGI9002gbstiCmcaR98
Rvb5xXxVqA0c7oNKrM9gUzhEkkwWQQ0olY7viMJmIUl6+UvYpgDBETfnJsBswNl5
FikVD+ND2D4uBGfKTA0tEfVGeL6/poyodpbqxTdoecAHRjE9arQlCrUQyRYRignQ
dd2+oAA/Ch7unZNEFZawS8BQ+5BQkHXawTm4u/MNmwHSz18vYtLJd1ks9gmOVP5w
mVYnAPdTz/lmluhBB7nqfdJWrKcQX4mRUdVczH1X4YLFwRqd5xp8UIEeDBpMkfPe
EhlgvscqcLAhCeUQn5C8pWEV8IX0G6Hn0r3GriwTw119Yzzcf0Bd8sVMHvDOJl4S
NLoawEt6AVM5yn891Daw8qEMMUgnEuE435HNUpeJLuuWg9qAwYjSUdoA+PxP3VDj
BrYvQoBVU2N15MOzMSGZu16JgpSXbMvQjWo55WjqiVqJUQImj+AJBqxrZlwKEwtY
/fUfxBGA0c0f5K8TKpBICyGHI1hP9OWy7gthULrRTQeRqMTt3hT4CyOkOwE3RZwZ
nz2rj4aW1FlJ7ncm+gxkNrEv0iWIdMKG4f6xMVKhX0TPCN1hN2M9hjqHcwO+uHq+
1iqVE0Ko1IiCT4um0qaHEjItIh9lbsbBuZrhLqR2zU3p5xCn3CwAD1ubV62ui12k
TTtpauGYezis5wiqjpreWnYChOCT7bs3EI8mcfmWcY23qwVHievpfnCqMVIjoVSJ
T5e5SnrJvntMRJZQtqvUDwfar5l7BJwOnw+7ToO0CoqSOXNx8/33+Rqg1/qa+JAo
WH/02+LPuM8tB467hcj4pLNGzI7uc/ZENHRzdEXTpp4PWcKyqTBeEUG4h5GO2qFK
lUwegqw3KoE+WWLg1TE6GOMEZkXecr08k7ip37sFWijUsc65qOjPru6He2tdST2N
vCdUiCbr74IUTzrVv04/mQlGM/vcimnofdbggugo8ABxGS6DgevYEsG6/Zu985s9
oOWktlKOnVoH2OTXr9Q3Qxt//049i/qhnwkwqvpATj9a8hYwmtQARcdYBe345f5H
4edrREU8SHkMtjYLZj4mmaeW3VWRQbK0HwSgjqbMdjvs/cP+uNoKNBjTOhlBn/uD
EjY+E8DHrA5HbMvnLNwSMdLt+MfpipJs/5VVcESvdH4KpO2hARKKdAyf7i2ozvEp
54vQSUgmTTuwbjadwbUGpz8qrgP+Lvcd5nzmdFW8NRCu9OMgAWckEpAcWf0+Q+e7
dP5RzbQhbQdLT3i6WZQoXgb545LLrKudHeEKhNOhAm1Nmlg6SEUpKtxkJG80N4Eg
90zx5EiE+SwEWGbTeDT7vJ8Yv8v4b7ok51JitjN3+5mkwgLaLZL4U4XUgmD3TwSN
TpqfURIWaCohkkn44thEzpDKx3q+KlQAH3jcEIcEWcPO0NdIx6AUvoAwX38TFNZV
KldIQZgyiUQj6atGIe77UKNJyVXRHCiO4WcSD2IECGxl4/nsBT/HK0cn2VxOgx9k
jQkroNjdyki6kp2HcvKfnnUtt+UC7hzV1WQ2PlGKjG7DcZrZTGs/Y3VcnE9hXHJi
gX4xz4FJB5rHVipa3obTovuWUvqB716BRWbG1l5HBAnoV41zxYc5opgEhIfbl88f
AIbMzHbAMBuJyURshQ7rmV+0tytlGP870WeblTSSLZxJprR5LTxJ7tms+L3dsAP7
DkLjaw8JZyZhO30VZEVNiSmPxnfjH2v0Yxzf2YDKIdfeAoEWNt9Z6+i1JHzYvDOA
TKt+/YnBTqT3JzIGLjREW0kacarRFWNAOdhYql8ZVvt+c+4xMQvANwEmZTJcHst+
eA7RRSk5Lu3tFMLqryoql+AGXRmyUtH5xzik+L914hWTdA+NijpNbj8Tow+y9y5J
5+H+pkZF7w2Sfgy0SHgkFyj0RgicZuT3ILRR63nIgZLcSeGogtBW2FxkfbQ7ropL
2WnmreSqTVY9UzSa9KRcjqbQqdDjQu+6CRCsYGauiXrFZqS32GrfASQ4q+Ye5Mpu
ljHKg+a8OTpS0CODTi+hOdp8E0PFUeFDGrAwaOtzI2Hwm9tB1yHiLELyYhH8sV8F
NppxNvKgalLeQTmq98dbXDNuCNyFla/e9TzcwHdO0Drm9tW93ww6n9HXMZ6twG7R
NPHupVDcLXAwxaio2xnWrnaUAo6M/mvGJQRjsQ7RAOcTL8akETwMNQDbDWZYTOMQ
N3p9+d8h3dtO/1NkUA/p40kkkde9M67udM5PSb5kPlPuE0pvU745AWBQbK5XUl5f
7W/AH6zHBqCQVLmybgqKk84Kp2CdKgWbwOeBtzK+GfsCPcLhlMxSuA2wB3DssipC
Wtdw3MYm2R0wO2h/VWgQnI6I74P6eWiWZaIqKwqsneHsZLmIGG+X3VzSEcPiGeRZ
dtsYN3zeNtXm4cZ6KU1dPOWTml2KycahINEw5y4hhkbMPTnofgLDGEswciuenkEd
K0b0XtqMBNTon6GIgoR+kpgCJv/vc26M7SgCZ0+yFbwxNWt8zxjEe9jAtVLDHVbT
oA04qQqFFBZoWGtLv9iNS69FLIvwFtzjnE4ButvIp1rf/DJkBLrNriI3/V1hchSz
vfOMi1jhWT20xRdt+0xjzZdrlk2ekFMmUm050IRQcvB/kzvOLtra8tqrWmEKi6Ni
vgu9Ictome3pTvM9EeFzup+SwU7D0CUA+VBmOIKf/U1V4rI7+zaPaBtQUGQZ7e+j
KtjWwSe6eujyeHo88im1Bbn8pIMn+S6ifTh9no+QG9IZ3TqdIzb7bXEE0OgvDQjX
48/ekEGmdyprJgd7t2kfS64JKzxuFiHUvUEsb3nvqjXqYhq+bBt6Younz9aMxSy/
HpXPnUmZ88nENBk0UmlsyvXRkDb0Ia+IzDcoJWAgsWnlyV+UUkeUj4ZCjmmBONkp
8pgVNgvW2u8/1HbrFXVuv25UckUMLYPeHAqJ94g01/JN7u0DjE+3VSHsfx44k9/g
8w1DjikD/l2gABgg0qyWKX7LJEvkaSzvvov8K0B/+05tnxDK/iirxT2Vm35YbOZ1
YW70MVjCtjU8r5tfo28m7NTyteVicrmBYUX8s5xHE4c/XwUUJf3ERzUl8eRK6lI7
VP6s57mht5WrI8t292l/0GgeNAapBiZzbdDRRkBCJ4LZvHw8qTjby46kmooLErJO
7OG5/c2Uybk0q9rwjqdVWb8yaIYRUsC/Wnpsybr7dEZb5EkBA39kBdUwOSM2oOlK
F/3loK4OLqs4s0J3h0Amc1sBSNlaxxqazflqSCERPByRTqKZwbdU/tLW5kduHpul
J7cs4/f+BdUHnfQ6FjReJB/gsJU3tb+w55i4x9OlRI4McowQylrF+KvR+Cx5QEls
QxKlCO59dDqHJPUAgwC04DNi4BvnP5wj3R6xinEambZDMCajQQMrIpQVMhwPk8rw
2jZsYGLrX7mczpRLvwbXUIA5DP5C/X34g+ilcQdPwx5QMymPH1AIbJco4eqy4o1X
HuQeywp7Jp/MMWnAAlF52qiLCbFCR07iah6tKAYz4ZyvXGh6PMJ3Avkf1LgcTwhr
/xEyFIfBVUod4C41wxUiEPKrZr+TaVyrvVVFQgACkbCPQaEllRmKYMLtSpCeKbaQ
md6xQumiTkkotHBVX8960fBjZvzmPWWG0FCJ1bUEx5mYZShCjRzimt1x5nyJM+3j
AK9QAOxaS/obAI4gBhw/LyFn3WzK6a3NqUYp7Bijj+BfnLEc3vykUmoVQkmW/dpY
ou322on41ucipSzcvoGLY2KNb7ZfJGCh5/MU3wds23PKkQHoJQ/8zufjxzWYw1J2
K+kcFxePrFDesFiY5XhRZGpCvaaepI1upfOyh++McVd02ieZzSccBIm1EJl4izDg
iWtcO6n3TFCAY4da1jxgDIiVcph/M+yOfhakjQwjDb436jeByJRdMAQQrDKIiTAH
HXZ+oGg0+/RiCj4Dfx4XHqEZSzfthsKZg5vFJgYMYeoWtFEokI+LXUsnPYco3NzT
f0+A7FoUgrBsgL7CVwurhiEOSLXFzeTIlynQ5oxVqkLZmoabBMlG6GGGEOf6TAKd
wShR8MH5+SoFo0/pw2dmSHIWI2YcLgw1AMNr7K6ueJ2zdOULftNyQpBRNhTgBjRh
47eATCUq3FunjPHw3dLjZbSd4itxX6ORszTWcpo3ieuPV/ap/L5xI3DOv4GCqofQ
u5Vw89YRjZPscoyKyl94861megye16avGrnhuCq2ko1RXGMVUBXSbsFUY7wySGsJ
Bwmc9MnRCePakBLDyWSZXkJIK7el1zsVHdPtOrGuOJw4y0BH1sSCesiT2mLczbe4
fqZ4+QyATw9v1jTZ+27ciI9jJ4QbYbmWYd39QHmk75nMpGvIC+bFuJryv1H7l+/X
fzSyHINJk8jjifyt5XVQsUBT60APhtYeCtMAWm0sSp1oXiMVu49erwPtptbfvrKO
l0+cdj8FRHZgzVsuwPqtjdxIhraU87N10Uqw5s6PsYJ0js0eyRsRvumweHPylcJm
9cWj3IGOJpYLzPlgaVli8WFILJwwHvBPhP2tS4nfEJhARQ2Rvg3n54vN6Zfythb8
fCfBmqvvN3/U2z2MPEh9+SyRVSwGofBiYm82pqFdl8WqoOVgDuJUuJUiAtnUVqsg
TElLrlvRQgdDMI9u1ChZOy2L8fFVf4rMDVa7kg4YbBqiJegDvxPdZcjjpBtiRb0U
6ZOlNw58r4axSOYFsGleAT1TmJnhXhncUfo9zupa/0xZ/javcDK8Q/x0qG8QyYmj
Tvog+ajYanj6ytOm8Ot/iF6vTrtIWo6c+hoZU5r6b1/wODqYv7wHhHlSMBf7psYF
9jLh6A7sFEejVlNyJd0i4aICKmIbGPcNQ/ODUsgyiFCujRAhKwNLQVWDoZyRpRrh
PCnX5vzIkHCsu60un6jK+j5IeEshh1dHReYxTe2E4bykHcy9/x4netN/4b21CRIb
NPTNAx7UHvDPRQnGJ7hla4w+8f42ff3qfl/gyTZrNpWRO4/Ksxq4jBemSZMKVIAM
kzVPdOeISnBAZn7SRnHcXni+uTvjhXJzAplU9EKnv7Mdsm76OyQWAncKB1U88S3k
8qiYPdFXUKUH9wUsxVQFSPJP3wwhuDGLbc1BBExndWNKF4xR+K6qySWJyUtZVhJ0
2I9p7Xfppgv7bPYO6v4S8XO3kX2JfROo48+YI/1KA2OWuQvyfZFIWr1to0K1FSZR
WEUDD/1gYITnmE6oJjDLmVjg2pS/urm/sc8Q5Bejn0gcqvFXRku2jSaslBbU6wD0
L6rX5WkJ+H1hUxA+vbUrE4+4NoVyqyWJfAWGnw0L0QcLzmA3hq/Jfa4s1qwowoaJ
WN6vd4y1R4ugjgwyqDu7NKkD4pHLOUYcg4V85MftxU0LfXDWxqK+buRcZtQbXkMJ
lx5dlwiAONvRlnYZd6Qcu5IOPMqNaOqityHngliq70nsyfpr1NHeFzfo6MfR2+bs
7C/uDWGk3xriZIIm2pfJmrnQb0Geapfh2GThZD/YBdxly+6v/wGXZW4Vf0q4XRlu
iMC3OUeJ3IcsdXDOL8otrOHTND7QJIjHUIk7OfQchoE6tiBAchWKByryzRrD6vRc
PhR+MKfF6b8sUBE83VbSXn5z0oEet0CC4Tjl4gd8Yk4G28uBV0OpKjqiI7o0YKR6
GRH21O8rPCzuWcwfDIekUhff7A788LvgSyD1jHxizuuFns4HiyKSujHGWTYOoVlt
hxGHPT831tqkda2FX0kGgUws3SV4mc7jj8clR10g6kzlFKakBP3Vw/KCwn8biaKU
kfBJIoOOK7OMhIMrB1imcGEdzroUUZzfvbGoH3KzYE0JH7NswpwHNA6mmKikYpiC
QlS9RSnXnahLi0q87buZprTn25G3kBMW9Yc7e7Y6IOWwMweZLuZT3sRF5yHLzxdv
oT5F7KIMYDPVkJupnpjzx/TFoeU8Ob4t2iFyqMaLvCmsqxxTmhSzdHbEaPzA+m4o
CXAe9U5htTHNtPIsYW0O2z1I5ZhVjFNJBLrq7vcq70x/SiWmc07V69dg9/XqGDG/
CTFfNI25VGl1hLwBOuh5zawy8H3aFCxotcQdgVsaTyrQmUcZhaqRE82QSoS2IR3d
IspYSZlmqV6Qw7LDFJtvzXGm78DwgFhNI0pVj+gyruR7vhnTXzOg/RI83CilRn7b
yzbXOiN0g9gHqx++YnS0+uX7j39JcOMFtkDrQgCekfyuX1saOD2HDoExxk2QH/Ey
xCBadz2yuc5c3rcKfAcZAsS68ternK9gEMmG6+LA9s4CxN4oTAp6zmffaxgMhQSQ
/TvjOD9vu/nZtiTvN+KYYNlPeo3nEAgAvnygBBgZW1ea+V3rPUpcGQyOANsxZogk
TEoIBVUKiH/RnAemd8ewVlOwMGCSn1WfztnFUAFLqZU10upCaY6YbAyk7NVx+jL9
sftu35/CqToSr16jgP95NSXIuoRDJDheWfNTdztcogwZoPpgmrkBDqOfTsfJX0JG
WCNr3B8vtee2K1VzeEvT3VSvP7vryhAsnr/g6F8D2e/nuKwEKycIepJGeL7p8T3c
VgEwUqR9LwmWZlL2+8KI6MhGTns4hcjfoi2EoRBCk+Z2Ncmq0IXTE38SAZL4VMd8
eleiAUlfSt1IagStEqlQnXKumBjvDwPnlwDAJfbMFr/oA0D5VoiTJPvoYnX2eedf
exeglVctjMbye43sLEMAgIoFj0icTVJVgafWWVsd4HaQizwKard0aocoVUDlfYVn
Gqofwh7qXwOS2N6J0O/vlq3Pld70hhc6Fbiz+wNSPAtRXNvBStY5cWvC81ugB875
+Ph2S7MAuv3pvYuoblkKnizIiMkIkRC19zgOTJu5CkEJZI3I76/YL9/7sGr+uFe2
yODf1rAtdroTzN2um4SbxIZizbgylQUH83mV00rkNf2O3gPkV4y+/EE0rLJD9KtU
kmchh7bbGD29V9HxypuEleHiN+oYziIrpUIrJA93i4pH9iBn0EJyudhDUab3SZOX
EXw8xkv5hfhIjl34QfkxWIkzeMZnW+tyaMkfAhLc5+yuE5jt6YHYO9whBRDF6L8i
heb+g+yCPDRkYSRsjyHDH7AJbJUqeuIrEeCTMgD3fM/w2JsCX4Zy7Pc/v6mBipNJ
yMqFn/FvfmBa+0v2X2/DmB936aK8Iyj82N/agbxE06QqCeB63gw9y7wtWeVpt/kh
VEkZEeToo33b0d+8DlJPWNy3J06r5FBeg9JFhNPJxDBWD+WzplUt0mOgsv+Hi4ph
9IlsUtBkcmTC2M9yRSbWMuPqfUGdbSxVbEUhwg/ReiaHbwlJRJ+q75Qo+3FJSNAk
LxGVMjitD8QF4kccUUoIyk2KZSTpCBmpFAfNviI750G/4bUlXgo+MoMh3qAfVOGN
quurVIZKmwjjeRUarT7vObVl8EI9kaLYLTpbioeLG1OufFyjGOLAHVszuKpeIspp
1C2LaEVu7uN5kMuY6ow/9t2+OKteO+PmLF8dohOjbk1hwlyUoilRNLU/a0w0u2Xn
4hw4gLpsfMy8RSKpsJvyhRS3dmcPJ+fEMmbL+vjgWaqJe/6Hhn//Mtm+VzVVfrgK
dyjUKIy0B7h3pINkd6F7yZfxC+UWETq5cFavjwTCf+veHAaoHNeCCb6kyP/UjoF7
X6mSiv9ElHJgScqgXGKqlhSn1OVzMDBJVWUld1Azr6DIDEmWocnPZIT23ZHygfVT
Dp2Wz+4cxShfOEd8sGwWsxIvyOWWEx39fVhL3hzVxCleM/FcGvVARPkTMbrgEAWH
A0EVAaYQkbIUT/f/qTHnXRIccdpnFgZqv99sX9shiLgBkO7MBblyc9oiz6TNZkb0
w0b0lhNNhHIWrH99rkmE1DlgipP4Zr0b/+rHogNp0Xz8C6+1e05RbImTMOs+oT6g
oRo0x84/KhIXzmcQg16fFhL0vLJUP2johm+EcTWcxoN+si16jBdPf9vRfs7Pqclb
qF5t2ReapZkFQ7VDwrlzFWUO+cElvhuOqnzPbG8tsfVlbzilNvezJ9vhfXcUnUSm
HieVmrCGk1AMNcBBS2mPh1Yj6f2T0XWOW2Z1UALZI3zFCs54LzhuT3B5QeRzeqLF
s7AjNwCvgR3AtYvWgvsY8qyLxjA/6Lbr8rzN/zA0syHpk2WXEcGcjnZyjmPYob9I
aKB7fUkeI+Bo1b6JiNcr+3En7ClZ3+PK14qZInungGYz8IzEjIV6j8TiDYahOkBV
2ApWZKCDahboW2ljnNfGxvTPN/BdIGJmWR4QvC4zE/qq52euO8W2q8Rk7PY8zqUS
sFFJ0m7AN3GsC6A3X+mao0ebNbSzXHOlPQ2VdFMtgAe6yP7Kb0pHzd6d+c0v+yB/
S/l0tB01TH9ct8vk7ZYTonLTylSNPh3ce29Tgtsv4DR/q+1SQxRwBvo7et7vPilY
91oZh1EW3pUMFZrjq/+FxFInzhQURZMehNQj4aHmucO/CnVZs3+A5fd+Udn1+Tzs
0cI95Qi0y/nsSJAD/N43aisszdXwbpjpij9uSMvvU55v1U1eeLeBYBrvVqg3WyaX
2KFTkBZLoK7Hz/k0GD//w1MwMRXBbFRmKZxKZXg0CUa6r+dGUM8ztSdn7L2WwfXE
zqjAuqsvPvBsYOthJ8brUNCrj7ASKG3oqiM/UTZDb3sow0lFflE1TNP/gPldBRTj
/lnPHySTcWDNQFUtMfpB0WbP/WlIPI4C9hCWPHSjf7jsI6Obnd+ohdW/mcrSx68p
Htxp4MeH1P0eHjtn3n5cjUr9mg1VJG0SbwtRipwiUSlllzoBJBh66YWMa5tMHGjv
0ddgeDKR+sHABImxATRBAv+gb1I0HlT4Ld2hoVlQefMJKh+To4ncVnr4l15DSpcm
mQ0I+GXsM22CjS8QEM7sXxcQMnm6Gbg2ZXOy46vNSXJ/VccZLvFrw1vgb50a208i
yil74qNLmt42dtChufseXa7LZo76OhVnG1ynQ0v1eEeXpsF07SihlwiDZZByTCK6
nXM2BWegjpkd9UriCZbm6WHmX6QL7gS1fhYwcQWyTPHN3gOCaWWElpTaCeIKJk1Z
bblyNkjww9Qh6hGl829k5crqSdkHuu8h93arjQ54Vj0jrJaJbr8SfSWyRr4crDGw
PvApmkmY84AgZ9oEYaKWbViqwEXV8ch2yh/reSNhGUudVGRY3fhbapqEdKYDot19
O/6Hpsr6xfNbke+TLVJaC5/o7qaJ7R8brym+mNouurVbr5zYVAtAWlIQJGsLUUDW
Xm5zE0jOoAf7aseLF079a2fIpGdcqZt2URwC3DFqEPFXcdTSqNNVxadSw22fIzDU
IO9Ije+RBWvC8TRug9HQdpop/oh0zLKJb77UZZ2q+CmQH4D9nWIwxG5VP2ve8MCY
5CvNLFxX8Ar0PRBy4XZyRV/g0Yid2kb4HY8cN2487YGt/2YKQUbbuhQH2E/OHxuC
0+aoPZCx98lhYeRDvSZd4lsTfG9Bd4H+iaJ0qtpTafISV0EEA+9onv9ThspjCrkU
Z8kb/hvBSn07bkbYB68i2otJjdU5eVtnIsMcqK6JN2JbZlmTzhYJzZq5llR8h4yb
/LdYTHEuK0D+1RkMCKTSkOIVizMIsP8HLNJ7mhBesZXkdeZUDZa2HahcrvIzi/pH
aw2xq91b0DGsNmCO3S1ae6fS6VNRjoXuIGTyuTjVSisBz9Do6sYKDDMCI7WITSYe
dE49gelqx+LfDI09Eymx5pIzCR1ipO8MI7UvIrRi0wO44gufBcZ5Lw5GKCSkUpWw
c4YwNVEr/GVjYkbJt/n1a7FPKeMgPjM3wq2kRq0AAqZmoOEQkgIeq5UgS9u2KOKz
z43oYt2vXQiEevGxRjMB4CXxOxtdz55ykh0FPP4PRXOIgrLB9cJLgnb2eWADPHiM
L/6TOSSdwcP6JWGiYLdNNXKfSIwPjY0HTFPlj07rzwCYeUAEoFXw5XFupoTNoQpn
xsYbM45fmOm7JCtcudyrHDNaFiug85a7k3BQJSnstASqR0USQFVoDIF1S1pRhbGg
c9lEWC4YzwRCez52pFJDIpbhPQGAnL1EVvYzrfZlvehSVVvq6VlWjjEMqJcOfflg
WtB3e6K4epIE/17RxM/kMc4OTKu2tlIFNhCVSVIsvqcFkwrZqXh+QlNXOwkBC6gF
MldaaDTStVKkA8uhiNMyBpuLKkHfYwkNy6dil9u+ZSIg0bGGMUBPCiQs/d+RYzbW
uAaNYQ+e83soMU+5+pm2Mf1fCCvcwFr2RT9k2dkXiAIHRelh+K0lm6Nt2WL0qW9j
DkFGnUrIHc+XPp5gTFCtDhkHama/uMB8K42ZD28kxUvCtsMuPRCTkPaSNIDF4Iw3
zCcNQnVqsRPXS/SAZXzPflFaC8M6Cg9VXHVHjQaozPJLW5uNz9jUCiiVbX8PnN5e
KxaIY44xT3/Q+jd+ZzaqFAL4QTVkAE/zBNN8M/kPHacCeRq32bm5T0eqx5MKMNc0
aIUp+ezwG69KPca3SOjSCO1gZSU2rQ0T516/rfZTIGAQwuJ8ilvs2oRT36QA/UOs
qUd8wZmbC2JQ9NTpWAEmgsyGg9lbsuO+tRI5OdsetLFc1HcVt/Xi2QId5HZF94+/
OXLcmdfNNnEQqjWiZWZdC5EPAJ67LALoNcXPxLy5Awrov6Dn0kUlTUvzuXjReKIX
QWLfPuCaGZBNTn63xV4uwIcnHZnJawUEvxkj3txCFQYLfQ/ogYTndOWGFP17NiMm
SSSwcf4BVN5EweqrrkfBKcQuU8scTm+laTNVO5H9bK7t93czqlvjYr0T9Zw8UEax
0BpN1e/Lx4dGOzuFIDArebx2GeNmm2kRtJVAt9MPfrHah4eQav0IA4JCuJdtooAl
yv5d6upN9kLBzTXsEAfXFaTAOv6DLxMKC9Y09B7ZXPYtYYZrjAJQzQjiFMxj2OhD
da3JfcGqyyBRZmQeNxIeGie7Ir9pkpZcWXbv+64DwIisIFb378vfUxAixk0MAsLj
vuxb/WPzqCOBLkw7uj+h7oAcLLPuXKlRKj2wltV3o6zNMnk8YGR/9xIdUmXGtEXd
GuNUHsF6gKdcWtSSp6cdQ70oPYIHnK2mEyy6FVXl2GbsQ6OmK/95Gj1OGvlPHnc0
gTbSXcZl2UBtsR6gR8kD76QVF59Kz5ZShL27WPYfm/O5nBK/DNxGZXfSShIhVIAy
vQoONy5iW5D4ljy2jfELUMUJtCh7NcjVChUxNt17nd5EDPncnkpWsceFtg/ZVJbX
Tz/gE028rGKaWEYLISwO4uAFoF7XDtJzUPeRBuMzuFYW+qoob4vdaAwWnho2Zfmm
wx7pXzN2ENkp9/C2gTHqKa8ST3wn2UPh/YxrOEOM8aEeIulgfOJ3cjbrRkcnr4ge
zNpa1GYWR+JCPI9l1U2VD2+hqxGFY2zRaqmRoJ3PJq9LQlXUFtUmmtkUN9a3rkTp
YjS4zhzrmdhAhzRuQz6o+7gBbhsFeDiYYRAGHI9HJAmvNWunrO2l16gvU8r2nNPU
G130M8UKz27DYEoloyKVFBjsuStF3GKCFtinwSCCUymIFlg1nOV/oEmUf+xkYzTX
5ET+yi0FPkDjvNi2+A/h/+GpIqTQrd0CfjSKSPzIiy3fJvdGFpTcpy9jsOv+Kjcg
+b3Fw6nomHY254ywJxvkmqZY4VbBaNEFxJC3vDaA53JJSHlzzzE9Pv+Al/aQdeCu
bfSwBfD+cpkys45A1J/kbuNMJUlzH8zm1vS3EfIeja+Cfc0sQpTo7hyIIzb1e3SH
3Jw25FDb0oH+77EwlTmINJ0FuoKEf1HPGIuws4bwQpzHUBwjUYbu90V/IT4ucTOc
jItAntQIIMlmxtbj7BYumsgnfh1TeoMGlU8BowMMZeD1VxP/mYxr0a0A4eKSjrEL
A5Zrnq8IonHyU7L1wieiiWLLdrJHweEqhky75or/PmuSdnqeW8uEnEu4Ut3Q/0iU
QfUX82HHcW8BHkDIeZ8Um771RUjNFr/IB4VIWx8M1QqKCG6ZOLiTtP8TKcLQfRcb
vvM1xWWmMY/qGIlmmSQrJ+TUC7dg3PMnsZXpBG9kwS/s08aG5ALNKI8ESz7h78gB
NKTGNM3HgtL12z+I8FNRGlkIDD/rMeyAWfi55rXl9CRcY7gLUN74NLf9H3+Jbvg/
/rpWACvEZtSaMXiBTekKUjEcr2l50KcQOAdBN2eK7wcYGo18TwJMMfBbZXLxNzxD
KvZ35s3UuiqvKgVUPy4NfbeUOrm9J1fqrng7WlPctUWRQG3CAbO/SiNtDM0EEj90
21ttVjwnaR8Ap6YzxlXHa2kZXeU8oW09uLRmJ4gswWEmiUWVpezQXus2FcOKqfin
HarKH+lp1Q0kQ46l7in9Pruly9O3r9VloB18am6OQo3GXQ8xtZ6qIaJfSlFDMLy9
Z1gi1fHEB9escsRR+sqMZYb3moI8uPvYJh0loCK3cqqnp3oEEY5rrEVWElz/7+QE
jtY8FpcWI6O0+UXIIATDQsLAqmDGSmX05IpqVWMb5pKwIo86258I96TpNhZikeDX
3paQ5Yp18DuIXOOMPPdI5PQGGTWK0IcfwgDtONDGEA1s7znMuL1SpT7X+1UXqMwv
vyWjC8JAaLBfkGAKO0Ea/OkgJxv7/ymfGpRMMXgUwidZatGpg514872ZgcUE6+gL
L0x4E212tXKA2t5M2cFdMvVPBN9+RT1AghfF1G38O5Aia9d0/VpoPDanE0ymCRYS
GsxTHFz2oSJ3i5FCP0hybhtSauq7sQ2RdiyZFutWzddEH94q7K2NOzCd4WXMVoIs
M+kYqfsYruTyYBPcV5BmHj+Lw3doZVRYOoWDt/s4IpYXUjIXbOt1ilguj+ufNUF3
3EH/aOMjTPy0hk24y7I1n/1UAKmA7XgODVrvcc8ht/o0y45DB945ecSJquzNOSL7
1VFHNvmQUWDhJHgfqTrH4UgkVRC2vPYJ5vBeSF4E6Vv3SH/p4ateldKXziyRO00a
zOmEGwXxOZ2pzl5H/3BqUApREF1I9gbHSGpEw0Mzfk5izqoPrEU09nBJv37H7lsk
OJ9fgi+n14YTq9ourz8PzT6CjJeefSASaOqm4cEXzDAge4umdtzIui1qqIJ1v8YP
54yhK9uzZoDDArMIIGHjOWZWU5dcN2B8LuWeWHbP+SMlEoXPd9o9osbuzdStLBkA
qA5d7G2EICMsThrg19rIVdOxxtcbyk5RD9fTxcRnreOeCgMWijPppbHOjmjxSVqP
oGz+gH36qRw1tVIkjtiKjKZWVossDnMwNWdEpITkMRs1ODkMmVEK/2HUztpBY1UZ
Mp4NxJR+VEqBwpUMCw4aezt7WHHQI6vKVl723P1GJprIJilcVKdobojQQX+0VJcs
AYEqi/FuTFpMLt7FrpDMOO1gFdcxtpaNEiFIu9LHGjskMYit0l/M1Cd0IaxXeNsZ
BHgvjoiMjyjmHNPCLRWdudJSk1KcJq9ZCoSY8k7ZFfV2dBKDk+bS80RN7wA+61rw
eQuHWbWzFf7yo5Rj9mhX6Z9zkjG2OFE+D1k9USMAgqqOwiPhrKSdlRwGXEs42oHc
XqW0adzBCSQt7jOxWtuIIeMsRvCXU3hLs8IEmWoKxmrSvmJy5fW+0O/KFdmlyJMi
7ovEH/pydyybzlneuRvhNh0VMWT9Pz1PHiyZp7EwAKl5OwaFowLUDNVeD6K7d/qf
cVXIk3Pu3F0vFmT/0lxQtkUfv6iu9xxylOFgqaZ54/0kofxfX3kRxsnTDSNdL4ZO
U0SS20laxWGVRDwixqcQcAah+Ymroxh18ZhFZ91mFVp/KP9YXsRTHwqPhIluuJVJ
kB8AfdzPN/7Ic0k52bpW56PHDXsv0ccrXtcGEG9cVzAkGcbTNVsn5VNRJxxVWfuB
MCTVHNOREASG3WFal+zmPtyrcOkKZQlINmoOzGRZSiYC9z1f2KUldTXaO0yQtNlX
p89zRDkV9PPfLMIAuO4cbjRCe7aUaVu4TyB3ow1VMVQGMMj0Mvw7k5YyDPQ/CNVT
RND5AzcSivq1LIebK6N1eTXkgaAtYS06MRldbj5vL/tLoRJ3kGPGkT4xPe8+mz4m
q3pn2ZOecJHW+5dR31+Yu1ZrxoNKY+D8uY+cb2kRmVQgdz2A+5qwhtvs6vLhKTb4
00mkhH37BMWk05qHYiKXJN3o69QPHFQxjj8iNhrEFiT1cqAIzuSli7n9yNaVFWUu
AsLgpnZMmpoVJ+TeUkOhDTGIwkUZPto7QeY/AZA8SQHAznAxACICXyMJ8qykRdtj
3LJ3p9/n/GL4TdQZtlXb+A/2ZxTcJpZUxfcHJkIw1u6tIM6oxaBpSlc03ZlHuBL/
gwAtRkahrsUH7pVOg5qQ4mHNeYEDmAjzOvsNIoCfDcuLxKLTADZiU0QempRLbfM/
bybgHsKlt5UhFiAi/28I2aLbAsfKPCb0+WkR9+0xgIxNxuEfTQuavkEcDX6excHV
l3JTfpmPApU4O3TMqDiij51KKCaaWkx8UVQKAZ8Lo303J+SR+nF88w020Xof0D/N
3Uqiu9IWMR24qWdXMRY62hfLDdk0UXYwpAgVimIMEcHd5OTcXJerG+5E3CHgNqCT
Unz1lY6juPJIxhmTVrJaOqSFQW6x4qeYNo+l8LyDisl3vv+ygeOfu+vz8L5nuyiF
8+qLOKjd6rL9EJZjUYeNOtMOtsgqxlKMAai8qLEJJuo180Zrpw7zCssgFW/JtgiT
cllid7hQPLOras8DGLqsKrWxqqz7RuX6ds1rnkFshdQMHFm6GauA4gdZv5uF1YD7
B2n1kXbBppLKf1mu6821YbnVBtrxiCa3exmYm4WkfTq9hQspTX/qa/rW3VQ07AmS
6dMrXEyUTCGkmKp7gYdP887munvahBctyN+h6YTpwvEkEJGEKyykleRTs8JKhYB9
7zZF1WRArMzro0JhqUAjZ0Pc0lM3RqChw8BR1QaqdNCG+PwK7fAPJiVdl6RsLUby
ExDugeP3t2ClCDAZ682oZ11JclOXIGuLYsBVZLIpjYYefLutttPNuTf/P8NF6hra
wGsv23bm0YvQwKFjNQbb+PPUCM2tRtGLQAbnB1A18FSRR90uy4RpZplg3X9eggfh
hvyPSoAMe4zPp74tMYEefG6eUOCI3wPfRXlhKevWmTuHZxWHpt4rzeDhwX5nQILm
qhQ1Fci4tMCLm6RtfJoQZ/r8IAmNVOhKwdv8rvqSzXN733yA9DDExaIZtxkcUP+a
HkgStHUHM+hfTVrSI91Lr3/paRxWfhHSOihipZabMd6a81khzwGhmt43HfozQ28Y
VzRDKTz8dRybVqx3QPS/zRtB4KIQ3cKMQmc75ZQMuk4nEEVPIh9iMXmPTo6GKE4t
UEMtjkS4es2NeJy7QRygsTjv5aOjU+x6TdybS6c4zaB+ARnn29XAtjZinljGc2EX
g61QCycMytiBtuEd4omzGuyPX6VaPmJ/A27kkR2yiRqlzbENsSVbjR0tNDa4gpuZ
snmcQMS/plZI1IJmETmYYKWAVfsARdqvY1b8IChAeLfNQNi0FDMQHGUyZVbflgey
R8gkC1kbHWgpTTv/GE94Groa4cwoc3y8dXe8GGtq3WWj9uM/gwfNzH63p9c67fir
Vr5r9gou5ev/r7+d04kkmwX3HHd41GjzVBmCQeKiuogMfePwvakuIsAbpbKlNhme
e/sYy1oJMZM3fzqQkT2txk3etn4E0dWmkUqLxMHOCLtDk8chlgeQ+Zp7Gg4N6xPG
BfY1Od0KgiTeezfig0VpHEQ5D33B9MS7TjMRKAj1jW9sSxSnUmilEYJ6NUFSo2lG
kZqR0fPw1Z9xSNPROPKjPRr5HwQUbp6lsd4mjdCa3IlaFO/vHNUZlBEhhRSHjAg3
ud+mjPqW5H3Qqedf18VJKugsB8guRxjBaMN761PT5GR5ZCCX8iddWPOdO0Km/TJ3
EOV2BFlt8p3UN+AQE9oSbctAxTQc40K8WrXEoJEpla/BhSiN6W+cgx7DC3tJBNdx
cTSHXS5ZVSFTnc+yBqIBJaNkztkUQ+/eRdIxhpywhBds0kwXczPGipKAzvi/FgX3
yHSV8zA6mjKA8suzk1zLgpAOO0jNPciQSIJ9I4fJH3ZmaFcMBod/iuGwVCpWS3y7
oX//s8r9XMEPM8OFaYbuWOlJBm+g1Pj8POY40GoJcgA3AjdD3iS0ZboNaoQHVrph
nFKqkbsNUWBvFqMBAeM/O7u4qkiUFR/gD8/5bLjCBezHagfOWyEeCH1v3KwP4vSV
lU/8Wbfkamk8K0Vr97+fIptIoa8gtE+3o+AmpSIv6oRlS5C4aWtM1VZ7/fdq0w8u
emiqGrfcK/z+qJLwIdUeiaI35kAats/aQklkA51nFSg6o4cxSMgNBTLPRa4qMk6r
CAXE51wrfr7jq7zJztur12ptDZXf/BNwsyTH6bPtC2uuDIohBfDBxW0PsdoDrwA6
JG96ZhBTImx5i6ntUTYe/FghaN8qt1CFKPap+OpJm3BzfyxTmQWEpKVvSAGzq3J+
7MWd0jdV4+JONImLJy20JAiuvWbrpV9xCStA6ZmAQo7cG1a3yrh/hmuL/oPauV5e
ZfcbEPNzDCONYmQYsCgNRewadiZpknXDWL3ogLLsnInkFdDZ6ZUm618aVuQARep7
D+QMwSJOoodd3vclaxH03XZOVE6aambBedmdZ2ycEHXWEbPKlgBFUcFBMXzA8JPb
+f41yrASIQo297nMg34F1UT2XR4u5KSPS3LwkJvW4/4VoaN7aKfW+7h4svogIPxK
CxSp606xJGyauIcSW4MYfg9HMDULJEfiY5fXJygorbG5hJlUccMOjRG5Zcm5jnxL
j+i/LaH1BMoSllAOwf9cPsxNCC3iAhEkqpD/WpnfJr5cvn1C9bugg40T0LQobql6
sUG+Xg0SghHGF3erMF0a/mLnKoDJfvhQnSX+X7+YGertyAmTczTX0z92G7/5QxeB
Tix5P51CvTzjOeRuUPQVCT6ghcjKd1BrvVuUpQ+oZxdo4AJ9O/lLkTK1XWgu7McY
KS542DR1MO+HaZ5en1xD9vAipl4R6x572mn9kCaWcIJdLKc50ao9AtvI1RFbziGx
X10ziOPWdWHXwi6x+FN/Fu7X4jy9ZX+2ZSrlx1CWzjtoLEcUbe90YQPorYVcjd2X
Tm3Wr48AWKQMM0NaMNu1Xfkvb8vwW5GkeAqzTpm9eiGA0cRKoUgcy6aLtKeoa51V
8OUXGsMfJaI20etbld/SKH8aTfHDvq0YhsvUWx5qP4B9gXCy6DF/RQbNEkHQPcq9
RlHiTKD9GHXt0hqUQpQe77Kph+B1rC1bBbUjCXPbgnstuqjtnB1swz8yx16pZSXC
zarqVki8hxD0XosdChfKX0jtKFu7Q4FPX0B3S1El5IB6UW4ojaDCDvPZiZCqVDmP
tp5oIBOpLOXBTvnkQfUCmBS4KpPmo5Vtzy1CPJmahZ8nyA6+5tiC+VJnIlPEBaCD
8qP2d0337vSdPHMS2H/R3+z2XHLCTITb93yvOJjvFZ0rVWs/akUq7esYp+q3DW66
AZXfbotzcgM9tM/JhanC5PF8tZfGNrTBAo5Yet1y+BG315fBZyqa5nGbJEyeRD/6
xTxnX0u0ellemnZHsZtvmXjp3eRjPG37WYxfiX9ZYfC5E6xFmwKlCyXPI+942DyQ
ngHknwiLbflCnyC/HQyW4TXIlKE/PLIsjaSWl7WQuoa36E8LOYLlMYxWCFeTGYbp
247JVMr1s6Ry2iIWakuO2+D32VQ44VfhIEHsw80JFR7ojXdBwCFz8+byCJVWo/5r
0sUNqF1d5xuHwBEJorkzj1GbEWLSy9VQEd1DwHsO0uCvQaeK+MdO9DQaJ2kiqcPK
laM8xKiYFbSVMoPp5ians8CyhoMb+2mtmtdslmUXdz2cFROtoYuIWyFGPsqTE3po
CRxZej3OZr3bG8tjfIC17PpJEvUuMXLGOXiim2s5PdVt25m9FGecWnMZYEwBcmrU
YMeqW79kgaZYPKN3iC3kJmHeZ+zYdiyGn2jHvOMle8c/SEY3mrX6MXk8sqe6KQ5s
aMlVZOvwI1CFCdnfIAecYD8PzmlmJ6oiKjfJ6Vjn4KlGdvTCHzlQvUwm/3co9V15
qEYa1QGvUqZ1MwhlTqbEtrIl6CcV02FRjPJTQ0I+gvRYOA3ZoxWOgtC6iv5CAW5s
2HNnyMyHhFWMshyjm+6wHfE9//Q4ln+j2LAxr0r1VWBkc3kNaCS3YSRhvI30jhfz
0L+KgkZHWHI7q0ZiPdpklsrxfeDTsFOVAPmaO+OIJTw11x3h3ypUJbyaO7e5v1V1
eHCHeiAt4ATTRZRFV4Sdpk8oB4RQ0bsD52iN4o+u7MmfR5NvgqrWON1f2/SD6wiX
U0U41u0ZlB3ynwjclSHOUsD09H92hcmvNdFSJ8erUkytrmEhnW0aCgOZkyrthGpE
1JTUDwa0ImLtV6QV+JyWlTMiLSbA0N82i/iQqV5bNxkpL7VAM5iqJm3FjqoxzzhF
bQ9WWUZWQGWgC5ZRO9fEwUSjvNtMhtjZ/kQx/3vBTXUy/MxzE/OJ2D8oGHZyU5Ys
H20JxCfJhdXX/y5uhMdFyHGlVpXasRFCCT9gRFl8o156uTzqFHWS7GWSIE56uKSX
KKuma4IzcBdgRrrsTbQn0Nm0TSYqy+BiJ3Dj67qJAXeIm80CwuxGdKjhx992M6EL
VxV+dDS3zbsnsNxgf4Xr9yUXF0pz9fkkZNUxAoxeGHkf4P8/1vlGs5waTOQWmhy9
ogoJ4Y58qm48njiTGC7gFEZppeESvAlp9QVjNyW4RKxviQohBqrMJoyCrPPt4mKr
1grpP16Mka5c9ihqKV81QHYG2pVibVEeT5sCmN4YQaZDUB9Ha/DuYYDGwSkPz9J6
25U9MEp/qfVCWaEZide/ifyGI/GEQSdKjk7bDHKzTJEPKpA+6uOMb8IJMa0Nnyf4
DcF+G7DexIm3ghomGQguJ5LwLxRq4bFzuEAD8gJDZoz3Vs/r9W8l3iAQCPy9/o1E
aZSrRTBtpTBm4iYtoGPnCpU7prv3rQmztdO+W1jyLmtFSHoR45T7mHbRmqa7zf+n
ylpHc8020W7jK1yFLmOyNW8C+How7iPL7WolR7gJCFpy65uzwGW/86m2cxD4lIw2
yiGLnzszHYjfrK1lSQYjJrmgNy0KXPkZ85e5D3nVvj3Q4lXCVJKcPnmNMVeE8bjf
yZ9L05A7pbC7RvidDZy3LTNf48JpFq0WZbgx01NFxmPY1dJvEvFBRgvFWl5sMoFG
/EynXtye1M9RFnfHFl4A3c+Xqxc0dkBxvoYdB0KKKFokcbC56qd/mCI4HE1oY4AH
sJSKxxDOzoVHcm3Mi4ZVgdTLCp/bxmunicaCe9BAtrUuf8rKlvrd/tOqF/rQVXv3
0h4DOKzm/6CUkmUqgfgLVVB5zSFCaxWYAzIWexd2YwzFgvekuttqH/vSL74cTmOc
UeIxEIrBoamNx/BTGa6NRy4EniHN1tOd61hBLB8jaseAAFitWLRNFKMHNZITIrfF
mojQkA/f61B0QicHVBgKofasCJyENYjgWBh2z2PuwtiLYaGjWyW9XVAFYAC2hca5
tjmYhmHkeX3lYci4mjQTZNd0+nJUnUquUH2h7ej99xgzPz9JSQxEnWyWZAh8OxNj
H9lr1F66HiU0T8rc8ArcvZFwiJoKVsaEZrLbYYI8AqWi4N8kCNBt/cvRSO0KUWj/
OFizIgyaVNJuNbvXldernCK7duWUcAZXBES8FQcGPW0ydFsPwyzDaw7ov8enAaIp
hFz/E+XIL9ZHQZmLno1Zrrt+o4tDS+BH1GLi55Ftz2K+FYgCIomHFSerFKD9trBG
8N6ZEkO4jIcAEaxGDfRBqmO7n/rnzeIfp9UMDysiqBsHhP1vQE0k27IoYivJwqOP
qKmdha0KIwsV+qNr4xfGcVzpfQtj20YQZ74JrFUr5l8PSlPAmtR8RMOvk+ccvTqW
RUdb7Vnc6hY4x/jpwN57urTX7ijh4rCEb86ltfoTVLRFsfn7Z4CoVgucHMmAm3vL
TA3qpn5x+BkH9ucJtUfHjtTnjMEV2zUHa4B+eEgk1EcnxxMgIYHi5jsP4ugJavWd
rslHlqpLIEVIjbKZEG0v9W9yef9OgrtpNO4R5wK71iSJtt6pHHys+ZlZqHqU33ey
PdE11KHcmcP6iaIp81HF/k9Sk+3P3Nyg1kQB1ys4HHdpWcfiqEVHAmJAzD2XT8BH
25NpABG5LTBVLnmtNs2Zri9PACr6hTJm9YGAylHQw5fo7s6542XDXZMhJOW7oOc8
QBOg6ChafYieTRYyP6ugYr4hhqiba3ibYOmGYe13X+WvuFeOFZmUEpjHSGWSOHac
luYA7wj03QJciq6d2qHX2WTTOWbvDt/kQm7AXCaS2Fw7WV39q1Nj0lIsAhoVyBH5
b99oFmLWUCz19052E9CAZ6i1UUG91nbq0UZadp1fv0fxVzaZx9F5lQdGD/h35Lcs
toXAnhLG4kkO4X3RY8M926xlhPknYhtk4oCFDMef7lqUIdaKTZxpyLhMN8McrJwJ
Fyeg5PS0ZIjGgqxD1/YWkr1JBBQxfGJlxe+OXe5uAhfdxEnC1jzqCo2ty3PMorg3
IN3YXEb5tvKluAcCPgwrIswd7wHR6B2fUEl3yIi8VQ0fx1PJmkLhK+MiThcDE1Uo
V4DZVnVTCH9D9wFef5Ro7jVbxbQ/7C1TSydJX7VLJ3vvoyp2YHiI58zhzr+ozbjF
IT1nm3TeY7tbX5pYLhXaSfIJksDGkeWKlHPv009nnbLko11w8WmXoGHnFEZVC9Jm
4154yDg+SFJ2mdjBh0vmUB19IEsxtf5ZgYxzJJHzkSJULow6ouIsBvX41r0HAlMf
geLMs9Z+va2jEMFx/eMfl1mduKpTtB7E9uoQ4qTwwA/sSEe7NYr51U+O8nL3T1Bh
8B7ojuFysYpZx+MXT4rPvLjy+1ewXkn3HUeZynxW63L2FTfznlK2yFCt66B4py/R
qByyK8R+SnRVZdQMwW5+Kiv6MUzAcMGb4tts7T3sG+qIM1vEZOliXVo+GqlnCb2A
L1iToxczgov4EtKHHwMa1wAkVBKn7dkhB4UyqHOq5I1RwEpsB+6vc85KiKNlt0mV
/VRfl35H/PPCITdRU63QyfAu6SJEurGn1Lmj+QDhspiZg2P+TAGLq9z6HO4byrqy
tYrUhVYLld6mgvzp0tcjGreoV+oPlPiZMsyIqQ2J9cVl/9uh3ynvFYSKLsWu/Rns
AgqYFbrK2O0Fk7aMju4iej2ZTtqYvSZEaHKheUY1AGB+IuMOV53urMIqLjilvung
04i3emYQ5+Nt1jJoZ7GxTnot9LeXbhLMFNhQiY6vVslVBRodo/ewTkGSA4RRIl2t
hhagedYXhNWOHZEMTwl5E0a5wTfA/p92Roo8G7lCQ0wJsFq2KZoc3Iy1IzgYeeCB
+WJ1Xdn52GcphMZFvWRO2HufbvRp4toICZnKiT84wACJIOFyrX1ADYelaNvIPe2w
IvMmqw+GouEdBY5v7rO7CWfGuj3Zc9+HDSjqk9YCbeF4UWBYThpPNo8C3AgXZinZ
X262lVzaNac50jhq4teGW/9hvhvCEy51MnXruQzhZovh4yt8CqoZ2BQeEGjWA0V2
d7wgmNNql0GkFC1ujsiF8iFZIHw/KZYvYIF+r+hBDmmynu4z9ucD0kVxJbvbUxhy
0AwWEdom8Nt2St2wntMOcDNDEptgmbk5cYpMn4NUAKh4CwkzQBDje8Tlluuk6fVL
ZSVUftGZg0rCBeyvW95Bq7oW/9jg5ECjO48E1z7ek4LB2YSBsLZHI6AuGaWGs59A
PPrZ5q6LvkdM8gkaNiU85rsjsOlWeHkTDZr611doQoaz9GrpoziF7yq3Cg/tcXrm
a/wnjqH5vNrXrLJ2Efyo5pd/+xKpZioyCXcdt3+2JP7pYZPdqG5xjg1Ash4wyE4V
qyyvKyjKV7SDqi+sv5UHnojATuGhFW4rfjZyUvS7K2B9dTD4ptGxo3eFrStBSqOe
HxYAQ8HRgpIGK2DpDRyrEA8L5wBYpbJFjPLQpqrxyD6srpuye2TYMK1DzHy0hMMl
f/qZRFEwuU6ppjKH8sJ5nUITvhJcOEBYMKceFv6nLZjxNYYlHoAuCISWZ9Rcb/ws
N5WmzsWcQEQNmNPyUEkebwBpHl5k14udjqDRyyg5qyVFwvXeTW1ToTSucuyBFcra
GPuO9/mOPpzgmn+bR8XOw0nj057Gsi0AJKZqNsoxpZ+Ch3CsvT6jneyVQx8qdl6H
cduBx9YZ0FvNJY6o9zh51xCdOXSePbntKqw069Pl6457n8XMpD584o3NIawwOY9h
mkX96faJZ/hCS5nGMqS8pa5LqoyzmhJcf5tD14Q8WqdBK67GqByMxcLgin30/KSk
KpVaaSZOgsaKY7VNnXfjbZ2I8w0x0Twc383ZtNA9yv+JPe18685QiTQcAZs/XO4o
LQbn/VXiJumwh5/J6P3jFR8G7O4Xq1aF54P2lOi6emU6Ro+PdSKK26collLs5Pgl
ZBlIhhLJ5btPz+g4M8bZpnCE1mRbu+guil1DonDAPzd8QG2ruDGHWREE6D8hgFAL
I8RPG2JkbdXrxCVFgQlXN+GnPQaRxCkF5NahZmE/d36DczG5+qiD2ScYIFqGxTcK
1NPObevQ4egpyJjIn0RNLhtaT0X81gcdGsHp8WrAJcqi0DayVdXpKC/AlOXLs3rm
sIH18ZbX4z1XlCmcUFVZK/yVjvKwowG65vA1hQXVKEmy+Vu4WZSWUgdIR4WNOTRg
K71awc1/LedbCH+iXDc78VxFY5UtJNY3t4t0Naa33PNVH3sN93aOSTATo56RnNDw
fWFgM0vqE2/9jPkPTDWqjMkH+AA03L3rf494X1Hl6RysfZC1FkOI6xzRfuJIGsU8
Mrcn6SGtI+ZdThEbkRWbXUTXf4+SOFLCiRNsgDo+n8cwpsSCHOYjnBdx36zVf1dp
D7QtXImw0yEuU9qL9qfHouJ5NYrOPePz3JvfRrce9/KH9UzjpBNgaq/12nO1yaE9
U9sYYMSLHr2Xf+t3VImHQdnoA1uJNK1KfOW4HN4ICwZm1PDpaVFFdLiSBgrMNfAO
XULbDPFGzILxWy83JmY8F+B2of9rDw2B7kNYSXv18WwoXNM0yuRFH0Z1660fnjzz
zAY3G4Vb1y1IHbReN37JjNZoswqxTBpUIg+8ZNdnlyxXYIBlnKLy/c9hp200qAjj
kQsmtjitW4QosqqsZuHoTHNo0p4PrMNdxZ5xfSlnnEztqFY2U/g1/xdWQgcSO2Hi
bKgKxlkjreJhRHqwUwwwiQlUcerm2KpfqiBtrQHLxou1uu5KvGII4leqihHcriZB
Tw/99HA2OD2EPyrE5Hv1K5dFsbieKIr9haxuHSUD0PKEkHonyW/jIKdd9rMhOftU
0BP/GDX19EBd/+LI6xVU7PAOk8A7qfP7A9HZ3eMxulBr55xjR9QsurOt4DvX0Y03
N5fKr6kGzmJG5itzDPMw9UY/kTSvyVrPg8m7CFVPLI2b+fN/NAmrviqrhkP601dz
8Oh6QNqt53DQE1/KdF/o2OZC7ZGuME/wScpvVeGs3BS7g3bm6bE2MSRkyHHF0MeE
KCmFTSdBv+PscDNg8+fZOqmQ0i2Yp/+d5wsbNkVian6fMGHG31OyLnGc1wR8b4cb
s5mHtn4nmpESRJ5lh+xDjanGhNvbClNUzh9okdxySnh7F8m9jmE6qjqVfZcSNcEC
KgbxeT+8tjYDgaEMERzUsmUyF8kJEEYEkC6S9sywoEzr3vqciri0UKr5Ws8qocFT
d92wGp/i/TdDXPhBSybhgvX+JQPA/XxHzfKOAYW2/GeTgYNU466wD0fsKeBBh+pu
vYdqSWkcCbPULkDr/liw764XyAsfocvsELE/H9MnNxQoU55qYRPWSqAfHYiu3cx2
uvmSE//yxbM9nozZ9XM9G939m/jNJ8PqPtIhRQ0SNF2JAf7syHMAygKw0Y6pr00F
QabGthcoqAhRlTUgMEepMJvDOcwAyKixi7PR9nD14jUgCUnaUPNzzinYVC8+yYEp
QhXny4GVw+FNxcXzkmrVRCQ3boYL6GvoC7Lnadl5rukQk4BBJsZVtxiIhe+87XGh
dmaUpnaeevAT0gMVRFwJCaPhSRAeujlHmcyqnnOviDUqC+LPyaNJDPR0Fx+7P5pU
Em3QxFZ0wczAgyHfYmJo5xePWHZWHTLNhLwoNiCbZgckom//J6VmCsXXhbZa1nWR
K2IDQe6BImh+tkuXm2QQSwjfv4LXAAWP7JjxEv2WNaKduOI1d/qsfkhmk9cxbbUb
sNLQpODTiqF6Z/SOscAubFpDfpKv6ekNohkdcX/5W6+PAALksSX1ak+9rlHHuDFf
Xir0yqv5bs5HANvPJ7nUzI8r9FplJVf4G5Q70n3Y4Zf5/FZgiEr3SeiGOurEgAmg
nKfz2xefYYuHdLak1HtvpDeLTHor6tibNS4qXt6KbaJVwfFw7OkUyYzZn514BtBD
nerNfmxI7SQwHOgh1BGUyAjFA+wvN/8KxzjL7KN1FW5yMAi6dRYyH1hIA4PqOvq4
uoWCQIHjU7AiqZfgRngbhe92FMsGGAYJmIRi7U2Fd15RMPe9brhC1cwvQRCBEtVH
Y79QtEbryvKR6n4LEn112T371MyLCyQxdu8RxCYY2vEAM2X62wnvWHxdDv8d6ZGQ
Ducyi04CS7nxw8L+h/BSSsmZZeaKXprH79lQuxqvPVhQlELJK+3C7qWjPqWFqc/p
d0Mig45S+gFSRIJXTCw+V2Dw73DpVw5QhkJzmAc2hjMTm8tEs2OaCnn8/AnFYQ1k
VgNjxJSQbb/Nw47ypexVqFcvbKexYiSGFfkzCdct6aS6ArVsT184yHH8BicRrKIZ
0u948UGikWuWl/AK3sjbIXFlPrny25oRdOQ3EfXYyPwp1TVB/Jzl64orP+/hfS1r
eigtViawVu2jdtSOXtmAF0tIlFJ5AjrN2Mk8mPZ5qGkR30Ex/ABGlTX6HeSNH3Ef
0M07TpwgruaztndGlxlt1fByyJ8cfgaxO9QnzWx+1B+lvIkl0eaQ9cTZmSNwzf9p
vuedFlR49jD1Z/O34HdYj6GCTaIctoXZBnhgdmKY3fYH7clF623ANljrhb9oqTZT
z3PeE1h4nHYnp6ZhEgOqy1aY4tiyH4gb6RNmPtzuXRizmdC6/GVS1M2DcKlE0VZo
IZU07ehP28RcaUNVweF72x+omG5N2eNKsDXoMNmMDsw0lYqkz+JBV/K7Y4kYr6ra
DVts6FJwWRFlpr+j9upL3yZi3xkYJIMhNiq9n/mii/xYzUB4tFwNvNYeneHPOvsy
iIiumKVoKFhmY0W7mT/WSHyCVVabNTc9vmHs5cZ1Fc6iNBlceHqyechavdqrExT1
m6kMJdNOo8AcqyesJILZeSEHMudSTRa70Md+ZFJZ7KJqLYN9EiRmlcPU8n3X/2EX
319ZHH6TnlP8YRyuPizjMH+e4qQhRwbnXApW8kkMedwU2gQbjUkHusKxDtlHd6bO
2lctAAIdplxKqicSmcDBFx6JMKBLvAWEmXpbFhsoG4JhHoNIaGk4PCVVbkCgW5lP
VkMI2SRfzGBs8Q6PgalU0PiXoNKWJCCnsS+gUP3f7Kacqmi2XA2agKjy2ddtF6SK
TopwtzQO+mQk64xdm9W76zdVYHYrX4QQhWNYMieSQKYIs/qHKXkWxXpUYmTh1Tkb
BOdDDL6BIXuN14BYJMPuN6GQN9T6SU5zIGk7VRa0uWB2RnKdq9O68j1CBIKH9SZ2
64KuU2eWjseNc2JrR6b99hjJZCbwUwxcymEYPv9vs/U6OPZQJfCI8CRSA1MEwwWI
wD+YbRmxcwE0avU54RplEbFjztnf9uJlxL/ANuhjHYQ9EwWcMd6Zd0QeGKTXKwH5
UUetCH36iJF5pD9chRa+ZaTIXe3zgqUzY5yNsHbsGO9i1oXavMK7bnHQ+t33capB
jogb9zHBF7WwE7QLs5PTOMm+vRliFNu6GYmGC/FFoujSjXfhoYMS9y8yr8bQXf09
HmWLiZJJ5z2Gt6ecilLa7wtwmr9QN2NM62kPjPdF0Byp+Pfbn0JgakJvHT3hN9a9
fDZN4HgKJ4IqrAbIFWVBmlwS9e2hkHKuBI5Wd0fw0NLBy8vDtMBIepm3d4st1Zm/
YSpxG6htAsdNC/taP79LAa8jSmnB5OVq76dufEXkIxNGDU0h9HhCTT/JMhTKHzEF
1bU1JrOU792Mfh5jA17H8v4wGHr8EnHRaHcNAF6IPKUjB10afQYzQBn1yKY34Anw
d+xtIqHR4JKHzFrbFDvhIpxQY1u+SutDvdpOV5fenU+QlPQrQOrSse59pJEK2Zhg
c9BtaQ0Q5P3n7jgpyzT+ikI6Ovtp2IwLqZ7hIVHg/k3PenekLEtOIJh4YZ7P1Qxx
InxNPLYFbQJDxLxsYbPjwUupwXr7FAvfPgO4hOqSEhfEchw0xGIH0VxUb3uWG1Eq
rwtouLRFj8+eTJ9ZcEBXxu0pH0cF5eFNOOszTcPayH/Akcd8pBA4VR7ZNkfYjCKe
5Lg052tHZMvM3LEG2oVC8r+Et2HvRgdocJG1ueHzC2GRzppuR9URAw7ifTlVxtsn
9UETk38w8tiZ1+me+XK4r8pjzEkCKx+Qu5JuqyTl0HOVzj+D5oD1a0S4tGtd9Qd8
zeKdx9xPSE0I82/iZ9lOWlZ/GxE/bDwRbavrXy6yMiKskO1uZKMp3NHcMuRakwXr
KdEKAdXoJ27NS8Gjuz8eHqpLnTYoeANStWEX6IoMmiV120HYFSltxd6wAZheStZJ
2bnRE6M7n9uZCCjyCql8IyCRRfP1UrZTi6LJx8Kws6kmZVxLXvIZFE0xFXF5+KI2
leTVvYS2wBwMwjm+PIfkHCm649XYEZ/Ri+DUsbCrxK5WG14SCcOARYGCuLKQmpR4
y2XRt5i50fYoaO3H/T7gIQz3LrPMFo6F0LowUdSHXLxGdirif0Zl3uCesTgsK0z8
dCVO5krTGFE5SepA5XYqaBiU4qpqJsh1B8RmFoNc/h6azN8TCL6kBNnf3a++DVsA
+G4nxIxtCLgMrGduc//feK5bCCUeze1drYH+4x65V/Y5atzDXfJElisUzlVnehTN
wXQUXHpuuNtX0m8710D5pm2D3AVoWmSab1vvwsSay28tXnIheBgCnU8i7BMV2e0h
JHQAJGQlipnLFyONU/rwm7U6TUwmjTlmvIsM4mNNNANdWGjvLLaG+0GmK91GWWGf
3Ypa8+GpRe1DOjmyGQXPCTZzXCH+AKuPFjNcBRFByqctChmP/wpa27F0jM2eseUg
YtV+YnGNJcAdz7/ELLDB6fBma0ufLMlfnFfLT82nIiHrGB1eIbw3LxDNm45b9AG4
ToVMzgjjicyp7NX0K7SJ7DqeFfa5jOtVWblCJL2S2s7Y7zuY8xTq8/W68MGnn63z
VpePjOARZYfnoa+E+f5/bGZEshgy8JpA76dSujhVzkdNoMRGY8Yojum5WXagtK3o
fijxNWHvfF1HIxMiIdSFYtTVvzN7hnIGKxUxQLQZt0eSj1Hf/jbts8OYHfpLiX1K
XzPFpB6pC5s4DRN2DfNuLw+kRG6Up+vVz+YiJQSTLwt7Z3ajmPiewhaV5yuFXycd
7SqlTVmBfZ1Wei5djBusCrEeS7HvnzsMoo8bqlJzDDibrad7HtdU/lFyNjl5a17E
7lK0MlayQJLZ5fdIB/i9BYykq1Pt8zs1IODG4ttMxlGaqyVDe33QLiAw/x1kNqf/
yRQflicLi4bwEtMpdjW2k3ctJcnUECpLscbS1nJBB9Ul0Lthb4Hidf/3mIhcuDrk
a+RVET+fjwC+IDddehxW7esA6aCHTbcS2LAZYV47hWEHrwTmIpcYfWNFFAt8Vydx
ZYLD55Uoq+PUKOuvCnmXgIZ2XPDdxrsjFoOHgAXP/usm1WhuJWXAoEtPpIyCCw11
1DXGwUdVte41ePdcPHLadFYB2eJ2yh+ZbPerMwAPiVC5JbC7paeI5E5VO2YBT6O7
Ees87V+EPRQoteMYPQPfXehiKxnPUXxctADBXk6yGPDkTy4/94Ea1kTeBZcwZ5MD
A1zC1RWfoSUHX+joykq0BMuPxvK5V8nxaeuS1mToXM58I0Oeli56bHzEtjhpVQr1
YLTcHqkX9R02D3C2sZbXWaQvfRpt6SAxcW+Fiq2cJjLflQadUu+OQfrJGKD6/lr3
yREO6TTyED6Sj2+f85QJs+/oVwiokhxnKVCJHSfaYsYwqSF/L3W7Dk9BLBk5uBkc
bmJwyq3y2rJ4G+5b+LQHL8MJqYOvqr/UPp49KmCScMm7G2aKVdxbvKLGBUIvYEYx
txdot9/BXqEQHXiSjH3ItW0Ng8wcQdoZiYSqKYpFPfx3RRzUD1N/XooHtEO7JOwQ
IxuwLxWZer2ZQeRQEja7SzNKN9EPl8ie/ILEgy2gw8jxqjsRR9uiwZSSO4ZHNtCO
cBmMlcs/KRPghqHBZD6Ms9ol7IVjetXagOKa8o8R+ifLYa6UteB5bbCs81qZSXVM
zxQdht4iVUztWed9JDanQXz3eX/+6fK3cVyGSLrI12Z7GTcu+5La7oNQGjRLi0z/
ZfcZG+evvrHe9RWMTl3Kv46OtOgR787OxD93TOe5gly42ys/vOs14Z8hlfXkHuJd
Fz3vknBukCyGrFRyhQFQ0NTwddoT5zoBXOs5jk++dwkcYvu/8s67GCgLrp8QjBD7
QCtdyPpOfQvxRIEsSuiGQGSfCaHvvAs0Fp1vDwhj+/ZqGsK3rnDkpupwakNNJfa8
I7VqVAb/iBaKWJekKkOD4GnKYetkcxa62SctD+tQ7l0RzbLDhswH4RzRYNInej6t
Zba1yisAu4wbzDicuzLpOhz87fBtgJ/k5IA5k0g0aoT3OHZusn8wjexloJcBVigG
1hpKy7w3QzvFriZXnicU+9SBDUrCmQevh3RCYOgb4kTeDKFX0SRUNCLLx2AscBxM
jGsIjUbdToYOzAePMyR8wjpwnbpeGgzwuPi2aTMND8aSdeDYvnS9XXci0Kdx49YA
AKyPEtaw40T3SyDRN7uwgMN6wKD2whCOVTcsqHSMtoa3RXFHroFJylbFCZd5CYry
MwHX5X2zz1/vBXF3ANSY8lntBCl5DDO3ap0Am9jQXEd0Bav1LO5ojd/T7XTV7kCd
+cJkyZJ+yQbxsZlz/CTKDbRTqkz43MeOqMgAKu/4Tmoj2D9NHlwMcEDfR91hMEeH
pZZeXQ22a1YzjJMkuZW/ibMHNTdQ3+EI74SVj4vBVwxVnaSH71LGO+bssRg1IiTT
vs1UNkBSfnn/5FxjaDScy/LGTmp0LP6Yj/+9ZGhgCNj/hkrEACxVjXDNFlmNshJs
yso/1FrvHiBs3bs0qN/Ci29GgZoRx5w8a16rO9FOiLUH1ZUejZcYGJvOobXcRuDp
RION1oC+MAiIg0XxWXJg4Zz57DQYbrhjuXJu8YZTJYViJuOJJPzF8xKgL5+Qh3uH
+zcTQrK9z+ElxpV9ZvunbnykztD9nc9l+tApjEuBIPXaxk/dNSZ7q8B1eWTWgTOf
1X1ymPNvG7qwuAnYxeJG/N+GIHGYljbUfzpcZanZGE+/pj0m39S5x4t6AkMRXv48
r61eKEa3yZGydoOxcOxszdL/tfUI69WcEmHcjMF4BBxf/Nte8C7Wj4ieDXOuBIFq
zvP51/5JhE5umixa11aRv6aWjDNROqFo51dtrjgHGebTL3SJh/fiUhzbMuxqk9RL
FfDz/uQosxlL+iyccAGZWa83iShGbfG8Iiqre0bzZgtG78StfjrlO//JdRpUDnWM
xdSg7VFl1L3qGBdnFJp6fYQrI560kB34l31EBc21gtBly/HVhsXg6SErHVAkk1eN
THGpMDazw/krB95p94dkcZ5m5+Pm71T3/iMCXFTLTASu6fMVRWxSl4OU6zyD8H3L
fQolNtO/SZq9PuYfL9VAvg/UGkEu04DTg45yVwMTJXPnei7HvcNAbjqVlsH4QtS2
tOGgWu/J9OAy/WGZ/odIrL0EqbTVKa+Rpljbo6SUsstAw+7X/nc9AHt34mHhzUdp
uBGchrREwQQKE6ZFpq6Lf6CDv9/5xvjewiTxMBYC4iu9fjqh/pZCzRBkBc5PfWyn
UyXRBuaPps5QNE+V3YHyx9qcK7BerRaD6eJvPL8XkZ46j5fT60wn5feGQm+XS/oI
4+avK5MVZCXz/k1lPhPDOGPAu0GPxN3tiYi/X8k4a2zwZUbFQzp/25MdC4slE3AB
bgVJE/gzzshAf840JsswFRHN14LCgjiOd+Hxhmd7Ku8BwPS4xPIWKdBHcEZ4WMzA
ztx4TYi+ni7LcESYhNjSm6Kim8rQn5WVapPb+lCjNpKxL7NmZ00KLiI9ZttbU6xm
xIVLGIhSFo/3MiVetxOVrZEpXyh4hjlbsC96kE46wu0iZG7iCenDIs8zvjZ8Ozmh
Yu+ohFkDfHonNZmJjP6gOdHpQVU5EvVFlgRVFbjZ9t+vYqhaGAGlKEUhgSNn5LzT
0Yw3e7sIIIrJ2sVzEC4QPOtyEMKi8b0cN9Z3fw2j2KK/scJ/dGfrCOkoaA56NzmP
tpCMMmDwR1rCQAfCvY0DPI8/8KAyex2IZjj8/pugTC3KB9TEr0AHGXlZrzv52TXl
FTqk9JfDTW55J5KOAhYGkbeVm7ICNNNbj+Dmpqb6ZBeNTQrjOtZfhKm987O7F3wJ
NDdoD8L0QWetT8M0sX285ma20U5nJRhddvPboeKi6/Cf6rKqMod6BBgyb8txn904
N9WpSqQmTL/VnSMDKrPQenhdn2XUgG7+ZNxfjKOBV6CI5RVdc5+aJx3blixtxyHE
q2vNBlErPlq/b9HQo1082xHC9ENMF8F0un0a39PJyfFTBJ7ysy4umHPx+rCffcks
iNoW+UXAcJmJpJ4NFsHss8svc2ZEBOKVwZ1m/IvnTRUyVtQ76su4nuFLy2PhM4by
0uQ9KYoEWGy8cgd0xNEfmjWR7aDjNnDYAX2mQ7YNzGYBJDxWAQSUtVWRYQ2WLkyp
Y0Bl3D8reV8y67v/DkuQgpZC2EkEVFpSDfIE4X4zQSVs5IF+Nh0AYTNAAwoYAHaV
fadD0Ki/MFQSO95BpUWGTzqMxYuA5+IpjOxQIDcYKK6gydtAk4zFd2kSqr0PsGiQ
Gr6unznCbE3S7sPg5hLoOFatppdY5691amH403DCoKzVOKTlc9Wl/VE8PbvKpaHo
Li21BvkZUTpL6t8llJt2ybRpfG5XLrcvgwQ3qZc+cT6ENwINLMJPbPpzyq05DuBG
tdxs1enpVvKvKVxUl1sbkieFuhIW9a4uRP9lhlRRgpCe6FPUpBskjb3Vwx3EQZpr
8KXnQt/Tygz5Jq4Pq7kI+zAw/XEzjAEe8wq0RciuHzB5O6ROV0/O6KC0OCtKAyYT
vylLfMj9KSZCXkPGxx+JAtfdD9xRI/GjctKOZym1WoNkpIPSWCTKLv4sJFW3QnWt
aJsjvFS9lz+ScyWhy2Dxu+vDbfk2ijNzFhk8AThnIClVAGFAXF3xcekREnruFMS0
UCrnWZJPFYdlhDbqWrTGWzXRW++3JdcH7PlL8h8AoLq9geLIKuZpFba52F3XvjQ5
NU25I2ruF4uh3rzyQXv9bHxBg+oRt6FbsGGrPRh81ouKSKoHuYUaUBpEDfwbviMO
BPNQjRkW+SHxnlITN2qXX++Zj50UTn24doipmp5cYJPxH19IsdYPnYn+ZstID6XR
0qeeXoS+taNqjP3YYdxqGTQjOIIS0TOyZqqXifsJtLSGioQZUVGx6xiHcrUhCsaI
LwoqHJJSLfGxNiBsME2q82qUIuUpY2otjdvV0wJfpeocRcW/++lNSF+prVs350Ju
zbwra5nVVLzQOoYUEG68smhsdbRryUJksh/0t0xVNF+7c136xqYmg1czGCNJdeWJ
aPBpEF/UUPOrB1neMN7fqteyPJYQg9Qn1JcdtjmhF0dj1H0pNReQOQbVSxUJ4rfV
9v9ZQ+Ruml3fb7FdBSwWxINC48kR/tyklqu0sM0BSQSOSuPAtHB7Ljv1RjD6pFIP
/aES3dB/daTwaexPlHjbkxlw2Ulnz6FH4PTbdp230AAQnRRLck0iMDrRKgWs9wT5
0jzEuWTzLvRwxuIEiox+YZWX6YuHCCRasvDP+YILGwWlKvPkyf6G1hYjuCmEy3/i
vBwldoMnDtiWUB64i34UXZEyfoDY0kIL/sApwtjy8WzVwQMjn+8WLMz+wWUaj1wI
SUV16+8D0bZOC5BldcOh3HepP2VFtFMx8NwH79LGhKyFeW4scHMPDjHDM8rDi7sU
x5gQ5fuEmDAgYUE9bXjbIydSvqwGfMiJLCqpTaxKMDKvi+EiJaHeyH/Ano+gUPmj
1zo8Joj3gU4QJodouf0egzLnLypl+85e9N+upEwf0qK4+NIc91ufrR4GYdaJxr3l
i9UKlToA1hrpWMtrzRwCmcidE0JkHQhWiQz84jP4s8Y5msq1iUkqcC8n7Zot7yQE
JiVT5p+HfJFDLTBTw7oDxhTbWIYSVhSfLRhUsXMcDb2/eog1DLKGd/YAv8PrPSP1
+LTk7W6GReJdsgzubY1U5B2eANR0Iee4uSryPBvJQxqH8t326UKTjBVKmu4SYFvY
WaUEcUObJIpciGXnMbMnPNtBk/FifYDp4yLAjJiC/tixGy/oG1hDo/bfO2EnjVH5
FEUsLc0smt5jsSVAVLZqPIEET/75R/dPKn19zF7ZqJf7E6/v5Efe2NMTNTtZnvUP
a2qD4FVKMswzp9eH3SHnAgagEztJpGL0yd+mQCs6qtFu4gQ3TD39krmotCSnu/rS
utDvAtEI906qPMYIH1tUmylpT/NhfxWF4Ctb1P1A7DjYsQZJzOKIJ3lldaMnmzxq
Cjavqafw7bqIwZYTGBtQnfm+K2YzloCuOEd1Mrx8OddczHM3ZfB6wRTV/7PmBciH
bpfBotQ6IH6S3q6Xeh9A+ppTYZLhF4RuMRb1veFL1rJekhhGsgk2RAOMG4/CCnHl
lzY0TSUL65W3WjgiftDqhn2L3reXDW271+4vvplhfeyrz3CFafN69fUzfR42GsHQ
CxhzoWnodvEKbZ3ovRcDV4QMSTifCApF/RlMjmGl1NOfmOk/ybUV2Byk2/n8IzyX
2l5zOHDTZEfjzk1+MgOLyZ3RCZPsiBUOKN88GKnPjfrucZ2pYK+yq3/fvzNl0J1k
um8dBJ+/EJybkl8qpQkVsEfTNtodAln/h1ApUdjhLzmAevmfMOnQ1OItLXuf+gIG
8TGm1yUPbgt2gLfHlhnsqkEMfSE/LfTCoyNEvUMhvryofqwLJybeIDlr102WEYTl
TgkBrBXm1Veg7aFoxmAi96g4ZOt9SYLCLuwsmDNxld+QBZBfm26oFkJMpO4EQZ2z
4/AHvWvD3fUfKqI94ln8DXyBDJa36f0DncsAETnkY0Z4VRdu9jkaoTGgiSK2f8fL
xTbd+GiNXwVH56DPwvRi/bdKPdQtQs17CVyu4GytHwJptinQ/LKjfiZFlJ9J5Ezv
mwxeDITAty1OPi0nRnj8FQoxFxYw/2EfxKvRSg+Z3WIwhRhg19Kssyrmg9kBTOw2
/mhqLB3GiRTK7StXGjo2cxRjr8CT5YY1VIcNeXaSSytyqlCrQ4Ha1IbW0DOIuar/
zADmVJE7Y9pLgBwrQ/LQxRJR8i+xBbhXxYsPY3w8/h8mJvEBE7jNMRb47V/iUc5h
dy9H2kEIavXs2Y1dTHS87K+jh8oXIEWv871c+HklmXtTU86N9e72a72ao3yak9VP
lR0zBTM+knRZG1bECATLGq4TYxpFzhkZ3MdlgIRoYD5aW6BbXYW3v3ZXpFcRTw27
0P1qyT1CqvfAMpm8ym7Z44/qiUd63AyyL/VjW8hYbaHTqZDBX3IiqB+Pnp+a0SPd
Boo0VbtYq3X5djsHWQOf11M3SpyFXlNSpfPDIhka+W6T4sc5BPF5o4zYSNZ+oz22
P9I0bcbBT13cUw4Zq2A5Givw2kErApmRcipyvM2IAfyxgXJP0KrWtIObPiD1NMKQ
yzPbLZQ1ahLyuXnNC9TMGvCBa9WWrMA3Q3wT4XN2b+GHF9VTPvptP28Yc6udmrvp
LCE0uOgbUwwUlyHUp7EBOEHGdlbFATznF8RnSHWx5en+VscTnkhT73gg4yHOe2vu
jbIbYJc1eW4BmbKGq9gWJOc6Qfb8sNuvJMNBJjLnrrKxhqNGEb7wow+e4JkUko3j
qAZ3Qp7A2K1NZ23SRHS4B626Qx2Yxnz5cOfRUAtRi8zrOck14s7U8HPm41eeMIRv
qqHmfU5o0G5LzSwurCiK1GewqdQKMsEjpIlDWul0zVZ+SFVbqzT3pfmRVnFWRLrf
/Hyi5gbikpeIv/Li+fnhC20TcTBjNF2HZHWEpM25vk2fntLy47wEMwPi+PmwcJIG
IV2n6H4ru9pWSV0VH64YByCb76BHDBjs3UD9SsQIYr2wr6XxBI1vfj49TGqzbjvN
en5j1nwtHVsmvsTJL8LfRqhvuTgMzy8cQ6oZtNCbWHL5L/KNS29z0tKwiQwWAXfv
UzgViMl4NXRcZuDlx12yxa+YLYWA2tt5oXWX/OG6J9YT7rn+ftk6RUjRj7Nb6wos
XBDlCia65MFFzl98CM2RFebMBRKpY74qQJo7fUkvaBz2mmgxKzCi9lEvBJJny9Pd
Lo/q6BRxvgSNVYNtROilYq0CJ5bCLLV2UnLNX14B6LroEGP6P+Js7FiAREAtlFl3
yv6TIlqEtbCXt5ZjH7bZ41E6C0So79XhL+FpFBBjzJPI8TIzS4lbUF+YglfuL9cO
PnolKGYj+2jL4BhZqFXiZcz/6KiFDzhH7ThIIMIXJdmlwHrpJq65KvHZEXLKAbIS
dWJDqM6YP/77pZpBtTKJQvXgDThXKH7LMimz4YIyFdxIHM48OCSuPEKkR8CUb0GD
rT27xhqWWV2Y9CrqGuQ3XeZ99tTaeEaDJmTMCw4y0+iR4iXkDmFQHogvxyXKDrGY
hUIl/P4KffxL8AyYeY4d6SNdsJFhzT58DE8W/doSOO4pY0yfZY6DfHqUNZEpQrw7
2ZGTU0OD03Gxnktv9Wh2q1ojQPAqegRcHg7UlscMjCVy8LskW1tMjeOjC0hw3vAs
ocn+GzWo/XJCU8yShkelZWnyjgMNer29WY3DbmXhpHfgUBH01idEjOcz5QVkXnUk
AIQ7s093G3jKIqa9Gsi10jN539kUGIQ9RJV6P/g8SH+d3DqVDyR/f+a3Rqy4WQAh
OnCDWzcgHaHzPEBdnrhRKcI53ogjhq0rNXDtbuJSa76P8FP+xnyEOYipFEnigcR7
qBqADxmZeYgFUkY2ZH3NqbwaShY1KUyJVzNCc9YWOavfSMbFXS/sxsawpjapjpGq
5I7NFKljIsh3V1zA0RAsxStLZdN9bhgO0+kETdu2aUMn/UIpdHTmoGfTEYJkHFuK
oG8AjCGxaMuFQtOfJ+5ZwdEzXI5Kd0uIZb1/FtNX8LDZJs+v7pNaPneuoUxzH8Dq
qkkUxV/bbHdxUecsIs/qtwOAb77xLp6He3l3Xc2Wnm8JW+xWGi+ohQlUaK7vH0YU
Rl8gCl023J++sAAXG3KWO6eR7gxnQXhJvZVElnFw/kT3hzyMr1zOEkAQqEbR2d3T
GFELBKPCuy+I/lMpO5ji/MR3YfWXcaomF94NblhqG7iQw6s5foU1sdU69j83cOgK
bMEterCxd+XSSTYodUoiT0Qrbo3q+AaLfcKBe1appf/qZR7FKAwO37ky6bWvIz+t
hS9+8+MhNipODWJ/tdGEwI2NFxLOg7mArheDDcwKxs/o+sci4qkqszkOwBE9d/1i
5l3RhUQN6bIrS0EkOEhxn3cQK0KMjLHmxdIeK+ZUt11P5AALXH5c43MDmrWuysyN
YVYmE1YRPURXUc42D+nrHXheNZglwAq+vU5UvZBnDv50tj26jmAGhiWNEsKSlGiK
kJeqIdeXg1avyppBbF8YF/8dNfIgJlyk228uwokkzTqbf4uV8qXbE/DWWJ0Ab0Dz
uI2uRS3qVZlkONIUCXflEdktrGhRsqae/yo7BJT4tB2r0dLsJuTSu5He4iKUlMAZ
i1+61sh9OND1ZznzlkkyechKyHcV+wvyGmLgsuzTGEHUpoezc8w3h8Dz2OKcLCWn
1/LRcqcxOuN2IFdaLBm1tPNFreyZGg+/9eFbCtVBv4IWZDPe839nQCvqk2kMixSB
2J22sSE1hZLv9R/xmvrP+Z7Nm9AB+psKTnIfF2CohVOV+NcIGRDVWgp86mVZ7y0z
JoT4aBT8hcFVq8XbZEu28yDj0GSN9TBSclDWqj6nPaO0IWzyHpZwKg7SVLLRfEyn
bFZx/3eO3DPN9Rn5Dje/FTQiDxT0Kc6k34uuiqYEVe+Tjk2eicGZqljSNc01r5z7
/bFpLUDEl3aMR0fYPPBJuNEN1QlHz0sE7sBP3rUsz78EJr/X7KLiINSKbRnduP2j
Pk9U+76YPZ2KTyjaf23vjPkB9fPGodNQWf0IlGALnozVVVVfgbrEjZizUXuswNNn
hXJeNi/hoI7fpoGO7Hc8KRbfuwv8+TDRRNroS0MysZGc9+rZEbLpbF8ysTONofm9
4cf+7gSxSL/ATYkA4ltItPcFKdqzfDULoi5Pcu2lB2spjvCHiztjm9OH46AJsqq6
7IipPeRUrRZjnESbu0oF6ZkmvwxcVC+DIAxq+1EEeff3ThVG0EgwMyAzeDikTli9
13zkN9JTp2eEU21C9Vm0FpRWyVjtRbdfeqLhKZXqvpSE4+ygUnRkXan+XOB9vdMb
CAy0rSHaiT8ZCMGVud6hDM/XlGeVnlhY7Y1DVdGHDtjORq1RRUbM9uSNd6jS5NoO
bKTv3gS6HK0dTlawtV6QulIwO5Gu1Phc2BXVk19ncfoOiFKT6vEn0H8rfGlSurA5
1dnL4+JbCUbCJerwQ0Asf2nvv9up9t4hlAbwRuN1IUqN/fdJfWZtZ+03FF/+r3bv
DI9FlTj8hGbRlimXaymX7Mv4ORDEjyozpdTPD1WYccH9LKzF8TzxtTQBuorsCY5W
ua+j8FcYc8zbUub2EHLr4fJQyTjet2mtxwsz8LiuUGM9lsljPosssHQRIrvfZCb5
Y+f4wZ0VyE5gg1DvmSbeu7XRw+YX/4f0E05JOYAV30Ezt1z2G8SzczYYgHODjnOG
2dgVOhvso5G2y1FJzXOQ+MWtEMhoo0LeMaVtgzTB2/LNzAN+Oul7UnEj/x86YWQk
vS57MuOExSdVUpGrCLr4dDKDNjdEHX/lP/BsSwcIFbietKjeY9yO13P0GxXSryyp
TGk/ff13qS3+2K/J5zlUsmsszmATRWimwUH1uhb0hMrHqlmQ8SIuXrMqcXbRQC2s
4qtIR72iXK+R4chwW1/VXrAGa2jOQBFE4+G1EzBvBNAXUyMjOvmUBAkZgdSoW2sv
SN12s07NTPR3SPZaF4N33l0NE60FoxTtIEikVh1S1lNt2qTIslA39MBzjdJO7qDt
TG5lWoZ1x7ESfVEakCBfsFmsoCRVFOkr07DQQF5hvQroYtswXG+fyDU2LKkRfjCq
fJKa3boGyTdm3t/39aCS7/Iw3yeDoAnN+TnKVK8C4jmb6eYMbvTsOPNCPCl9TNK6
lbzUMAkjkRyUWOww3B6NmKE8lHKQpb8wyHZWosnnLr3DR5t1VTcgp1Zwb6ZFYWei
Y1Dvwe7NlJLikH8kw2O6IxmfAkIqzXhVAISCFmnE9lqQKHQq6DX/cBFw/2zGedtV
L2EpI+D2ZyyzQXZ1qxkVRWtP6LmYdxH1n5IyuQuWID7n1FwtBU9dHY7eMjXwwA5a
DEpBIJOqXM1+m0+FOvtZoXCtBtkZHLSkpR/jepW7Ib+W33lwu25QU21KVFHaVD+M
p9xLA923St58Bo/Ou489mQcf0AR7n8h7DPQq2xXrYvJlhUdhwmDzUoB1MESpdvyc
Sk0YcjQFWFN2F4XMZRsdTfG8O7VZx0QcTrlBCq+buLuqvy8mrMpXIy9rgSxEFuME
WQ40rZ5jmoMMT934W9jT2bDZE67gkMk16E+88zK8Hvulu9eEJSCgBlJBgYRzKSeK
JJhoyT4G7pe/d5eZzyMMYLSd8zix6vb1BfaNgWqZViX2FIxoU6HoLt1o1mFUp+cc
7WrLnhrKwBu7c0qPw1o7o33yjAdOmyj5pvvO0pBndMK+0IQJ0JquQ7Q10tFGJqDZ
fyJq5mh4v0OZF3DsVCUf7wha9pSl7WKFlFBWj0MX/OJwdOBdb8MFDGpF0WiYu2za
WI57JQH8tS4U8v4ir8M+qPO8QsjOnm4grbwllsg+Ss556ukKIUCMGD4wa2/jQIkI
8qlePan3emx3/H+GyNagxkm5laDvCUUtLeCdOf1M58iTRxIYll5o7eAIQ/nevAn+
WsyaDD4jXI9cwNRRjyW2mSgENrNoRX+wWTPmgSyu6LF3SrljmP3oSCsKIIS2B8AU
IoborPl89p1v+4+G98vdK2/LVH9MiXdq8+mhnwr8YJKMM81wnFc3ZW/PE8EFB+SL
Y7HsmEBC42QDJMXGNhWjVzSKZk3JgjdrwHlEnPtH5E7coWwRa7b8mVWYF05Xl3Wg
MqFFuPHnWXZUCxURaM6K0R8ozHpxPC1W50q5JBvbaM4uLML/b4vQ4X/gmrcOkvwr
yO53bFzEMYd8E8HJBhNoe5xV5C6kW34MsCtNKimYwoiYqsch0/lLnUu7K+QGccF1
5S/b4xKldOZnCbqsqZZXTF/eqzUtX7OPWYuABAXlIiO/W/KkvbjvsVtI1xLPcvA6
AqqB7EoX0TLoUJQwtjy5B7bnY9f5UfaRynV11ED8IwUAAtGPoUA3xTvKCBnW8vYs
f84tPDml1inIo77v8B5LBZoDfTc97sxGYfipE129W2QZGYtabsb0wOB0WrxZzU1+
0XpVyzdSsDLQpAZn6d8ALZyqC2BNl0dRVaorFCjvMHt/5JU4R2FrIo6WbmkG5ukV
zvzJbGI3KQ+iBxGKNPGkY0PGYJSaCb+ggl6NBvLmlMfo/oq8nPufEmmTDSeOK8PG
fD116BanHayELwVD8XpVXEJ1YyLykYCbfg6K5UhT8+VZDhXTS04/p9x9jpPvWdRM
FofYazRIQWYnqPlK3B4X0vtcVj3dp0nS3XcOTeglO5mh62tE4ibfl6KWr7Bckhic
tVMR3Am5IS3C7sTVr+Csf/RIs2yWkOAHymC4B/KQSjmQYZTW06g98BDBvRreiM2l
ci9QnLIOi9LJtRm2mE97fD3UO1Fl9LY0dpIcyyrNwmzWTV4rndnLMpLOJI4ag4v7
3jYQkdn8p9DDHkNEK27Oid0UuxDEE0k6i3GAHxyp57uAThRUCyCgyDvXMq34vr/x
dGjqmVmms00/3m0Cq9lpJfLL1CpmkGf9/Dw0nry0yXVnMDwNTR97PO0sLsxTpzfA
/mh7Y2NyVJbS/vSuLFO5YF3IaSW3oRCiu8hRkV2wUymOnZolFROzLuaRZolWM9om
8fNmjigI+jyGQlzgiLoaxw33+V9n8SDRoxU6aV8ivfNDyA4Lnt1Sng+oHwbql2dU
oP/bV0KRQDK2hso5PTU1skjgfNkACkX3Rzn7RJhFxvEbXgfogZOKuRNeZB4DAaGR
hcq+Le4EDNzKJf13XK/bbaFducXJgbOFnng9CatkPUtpTV0P4tPUxuwgBpO+y4kD
2zQNyyPtidAQtrTM0JnlQ2SO4wDMVVGd+U+PGcKSuHQp3C6yZqbv2bF1dgAdEgzZ
nR67BOCUtKpmE4Qm+mTaqnWq22CmSt+qKBV9HOORSuFhGAPQw1dHXhzYsugz8MKc
OQDrT2/JxD6C3pSOmvqL+laSeKtsejpzYFgBHVRLno12Tsk3fcQicTMQwZDI+6Gr
k6dzy8jxYpDQbFto42+FrejNBAeriifov8cYga6PheahlKC0cxTRsVbJynU9ZHk/
xjwjsF4+jm79Fq0ZkpQWboQ+ePoLrcH/78m/nRM/wG9w3QD/GD4jE9YsM0EXg8Xi
gt2MRNYQyKXp36gUro1ycFmJXC+a6jWG5B2vu/VhQdp3ZvkjLMDgMuDvb2gqoLcV
RhpKZG22rQi/a3gxUnzrTj67A+wcOiSyOgtJKokPCFYMvibBeUKdEfiy7hHD8//W
v8vzEih8iy7ZJyE36VOaGjEoS+PONp0SKSwgdfSZJv04gTKBt0y/SEioCEnedJI0
zgHwwlg8zq7Ja0i5pD5D3e+/2ihP93JAyWoUYzExYBNZzN1gOyboGy3nN3ntcPuI
tednJRbG99RO+t1vGikXf3iiRDY+A2NFVo14bjbMcS8v3XSH+g5JpKzEI7Sd0itM
5NGC6nsVyiUcgS9zywMLxnjLhNHASTD6dMnp2fbwGebmFeDodlp2ppvkezKGN2JP
3lft9RePI3cTMwXwktVlduEkPMEaaT1UarIBQqvXE1EISckJgZSuyR0lfoQWs5NK
FCWMGOXBHXVuf6SB9IClsdVmF71GGApvQDM0gBdZpOFv0kep6FJqMXat7Y0hkl6T
seTS9X1AtZ+Vxpu/CXGb4kdQPRL9YJr5b1W5ubPyB8QgPpt31BcX9cciy5kkBSOY
BtHNrExHiOEMVGqJebC2ZbeFvTEvD7KiSTOG5plmbHCTiBAeLXFkuX0ULlkmaRvd
wpXunrUwzfnQ9z2z/MhtBJEZx5TYqwYeyDrUZ8li17AnrAhIS//BLAgf6pS4v6Bi
qaFhI4lIgjNWI0hRwheqJrK32ANLwph6XY8pyoct+gpquvWXffn6yxIS4kedEThE
DTlVPuslWKr/gquBfWeFEp4YKeEllBM6synjAxBbC+KTkLMYYowKO8p5E/i/pD9l
vl187hDiWHAhIV+KGLCV/4RyI3+E9I7lxto0XS+tvs1lcDA1ZsT6iMpBLYs/R3/o
7ZBPyT73HxDZlsb9vStkr+8t7wmVnyParUdr9ISugrvHqzV9qfn8qcaoxUgIkURN
qGxmKvfiM2A00sLTlbd/8xxm7O5tmYzfeGqkvVlTh7JIOBbpjhGMtSmfWr5iiP5e
fWZQXLZ8hQ/NMSgozm2pI6dA5RG7yetit3irJM3aDIICW8alW8h667WLXISShPud
0x1Y1evv7qNuID/mmtmcmq292MkUBEBNXuOXhpNKsa9UfhpJUdhg5U8IOlZpU4e+
pXWhhRwrZVHzGueOhVUXAhoqQqiuQrr8/8JZ46onGZ1729VES9yEHH7oRTELKcNa
DJ8PA+VRHkjryGeGdK0dGMxpDBaDQmBfLmdlo6Q+3Q1nEmpUhzZE5TR6QExo9hqq
a3ErfvEikItZZU0JjyEe0Xc2m/4kxFbSe7wmPQWvFBzB/RRBq5bda0qEMSF12WBF
ouTWoLqr+Pmb7ow3G+rcmHZHdE39/sz4V+Hf2zulLiUuV7l0LPFpgk8KVeZh5o+Y
E+uoRHQ+uDnSzT0MpHSiypzEeVFl21T8fPaeV81Am71cS3t7IRvpXvBs8lmvoJ9G
AhYBMnf356NwA3Ajz9eIgEwBgiJbV9uulrPAA6ggXkoP5gAEucQaOf9s5PQ7BEIC
fk3bFde2q6DOO5fxv239tTeuDPcNnmwsjUTsnI/cHh9qm0zHWIRauZZQfT+OsHv6
L72YaQM1w72MJ0MG7iHvCtP+mqmSIXyDaWnEXKFPDBw+KXzE92Kg7h47cialfy+Q
3Eu05Yb16KsUFmUYajVO3TbYf8V7Q2qX0ypUp0aS5DU83aSJo1fHRCrGFsYhoDEY
XfJpYFmd/83YDmFhIru4tTmnjBJMgt6ZCmSdCwPRAsNawMBY8Luxm348LW0ig1nN
yjLtIRoGuoQmU3o0XCRp7f1CxlC9MWr35MUU9Yj7ZRVUJAF1JF3bLED02UwkcYww
j/uFwgBRG3ruOa7BPQbk2srzfy+IHvtEISBwqYkG9RTLgb4Qat7zOn5bubOPumSE
W0QWyG3lxFPKAp7iEci+GBYONSRSDQghDFatzjVFh1R00QCFZS0VxTfHgqj26Uij
2nfMj/sBxb8+6RLNMJhM67OkTcMT5mUdudZYryACU5/v6ScQ5Yr68jV8QxrjLynY
+hCjZ5z9qVo6rk3XQIdBHnx58oLHThXarttkzoS39f8lPnTIWJ32TcIjs0P1Jlfi
L4XnAGfTvayX2Pmu+XANpN064ErWfSyHYoymgq/2mQdf7O4W0VZgQRpCiUBp8Tqu
5z6OI7j4LLP7i70lIduN+XtHYF19ielDjRd9eBJUUMqStWGiEP0t+6FCDdTFolsM
VYFIjiB0x8ecHI86Zwcq9nK7igpXAvq29M+EJude3+SvTJIEYEIk1QenbnXMm2yH
R3807Bgh/7TeRPY4sRsCYNpJqicvtXHC/xg75j4eS4x+RRarrBDwhF3/Tx2Oj3Ul
gyK2FZgrqi55TAIwLmBEqnmG0nvM/B3RzlSYepzAvUazn8O+XoDHvr9AAb5m9kBv
EBNwvk7FNdhhl1z+6E4N6g7VYW79Pl98CfbJLhcbxOkxr39NWa8W4rrdfPb0Puq5
qcGlAdZnNXfsZw4VUFBG9pB/TwvMwjiV7CgY7jPckUek69vg7y77BjLWLPrO7cKm
pKaGmgsUB+FUSxjmvNZdzrAV+KJMU1qJiMBXU7llwVMPpmvEZyEe5SADK+rTMrG+
3eISPXSUQPkRSzeinSgEXq0R97xFQdF7I0Mhkd3pjOV0NfNxT14Ql9tecx7hNVa8
jWbfDq75zHUeElgI+7+gu6BQSbrEh8R1rj4Ty0R03shNn+3o+Cl8UNzSQIgCm/qm
5qzy6SSuDC6EJN3nTgpW0V58ALdzqbzdzkS08L60lOalJyOabh/J7uqkVJd9OgyN
K16bpiCNXwN6QGViofCG7V4qYYqAG+nJHvsbI3jPtbOfRqrMxHWxd3mgtyNNriaO
zaG/h2KrzPBIOY2uJGh/a8rm++xsApyGiDSCxoSx8QU4yNSSbZXm3hXvDJCGmud9
Xtr5jPO5jmBD5tAx+gdDoMHrGpDmuR5l3ZmfXRjmz68bG3Sp6Ps2akhlvNSqHONv
j68ivAc+S043Fa2TRefGh6mgAXlZVNeqeffGlqjrzEQosOocY1pDk94Nv9+RfRFE
HTKc/1CsxWuzN6WJRVxaFG9yU+Hynho8APfLrcI+/uZIzwwh1ein2czD/NbfxSTr
/eQYJB1bI9HViINOdJAwRaLxko1OVzvrfGkQz3y6cDzomaN7rEdb8XrGtBJuhVAy
MgLEjGtavlo00HhvfCNMfw1L+jdvThPOKFrMh9G2G54bptWydHKZ2Buo2v88Tbkg
MYr+EjqiYYVPkYHi2GLzAl5OXpJBuLMADGgeFQMd43zSiYtCBRPVLhTcL1jL0niQ
YRhMPR6y8TL/OgPQnTEbUM4WeoQieiofO7AezcwBqKwYDRAAedcm3bIZdmZqjZZ8
K7/Ql15CEOGzqOhalFuqIbG1nu2lsn/Ydwll/5L46uUWAOFENubVIiYpBqoMb/oQ
vkdBO47En9XawMqF7EsPDKkJCBCwdByDbPtRbjKZhoIPVgAJL/2WO2Owd64xx9Ai
a2g64Ij5P7SKQQZL54JiebKkbw0NEv5WS51b9cB1sGjYZYwglPF9otE2cqSOw03p
EjIJB3MTgVINuGPfpLLdRF3CpjBHhPAD0Frxz7eEkn91erzmXWSjmLGZ9oyrH1fo
3bJCmamZZJtURZtIsU5Yd0CN7zNH95d+fRBr8dCn2RXndUDdXITrQ7PpRlbSb1/5
Dm7kQfccJaMqewVF/6g5yELj4mrmzIK63VB3Vf0eBYS7gmooWAHLcDW6gEIx2+jC
alMmO9J42VyzojcjxmoU4XNy/kPyn3FtIYUOVKO/WBq3QyRHniwBOCV1nJub9/7p
29XoPDYLY3xsl9mBGfdxzjdS/bXWpu87gBT/kcUn2e8HSyORy/gwnDN53BnQl9Lc
7g8PPqhM/oqQUIl7UL16aJ00I7J7GKzmLP2+qoofqObZcD+Ad+FI7rH49yCUd6cD
VlHv6rVOb0Fs7I21QsqYrHEa9/+JV1QhrwcD2bSbkWLvqNupW6u5xV3IC4uwLMaN
ZU7IA4fNw3vAy4+6X/srsoW1iZxyoG0UHKPbX2YsCDgjZKBayFxhYh5xCDtwwDE5
htFdfmrLLwvEoX63xciRfNlFAsSVl1zVCvXs6GtpqzJfEsVt0327ncK0vt9iIhiC
2/kjNESrMB8LPiXN69Io/PeqE+zUgfVexsvyelLUfbCEEbWqFa2hCfkRWMFPDteZ
9PIxHXXBbjBk5zS6bCqAdMrO1EqpjO3CxJgyvR64gYibm8zwLoxzhJ+jL7Vq36ql
1PXdCq/U3CyUQUMKg9EZbIRe3czu6gASx5P/X5MNfDOhsrvJTsZGf/HJODNg7x8T
WgJ/gkHTVoo1NHZFU1ml+XFTAqfLPGLtuHx3gSVb5wvge709PAabSdVGOasmDOBM
QG6RlGAUAloL/WPO9BGxYVVpRyBoylaLoYAY2qNjRQi2squw9Htkui6mF9YO24Od
1Ain5wazONg8mxAqwnsLryxyZv3cwt7wKMrUpu0JiTWiB1If4rllIFvCWTLot1MR
QXsbmGwUKIjHVEEC5kHY+kZwZm60pWFrYqvodkSn8uPzRbX2BJWOArAPw+4NP3as
lbbp/hSqZsqpFG7dnegRIjRjMPask9NK502tIxIuGoMbV0a7duOh4OQYD0LHk2Bi
Lgi+X71l5nCIAZ8WuvrLDjUgRDqv+9Yvi+g4h3s0JxId9rDbXJE3grmm7TjSOB8o
C3Hmiuamki06zePmxkIxRky3YlLJMSycLikQ2Y9zaWduiMr3zti+5kmx5FvaojaN
m60TwtqiiUuRobkfBSCJyv6a6DWD8AeUYyF2SAYJTtEpl6QwJNJuny0vVoK0NVVD
qPI3IC25i5FNKAhPjpIlzwNjUnRCuiGNbTevpk6KDbyGUqJtjevv+wrTO8BKsIiU
23CzutibJWlZl/GfUABXjcTmI6K0uBFyPOLgrGJ7Ty8sAuASkCQ9er2kJjdsjW1m
iaZBYU2lqTECXZWDynGGW8+UMuy0vYBrNhZE/ckhhr5G2UzcpfD+5WBirMw5I7o6
YnIzsKSjKWnVcDX2NXJx7HGlTsuWg4ZvUghSfZvsCdpC9ElvqZ/2JRjW6IwSoXhA
NQSBAjldBkG/JWEwvLeKJEi7l5i9M3LZkrNADF77j9+uQYRfWepNDWDK/aE5NFGv
awDIrpnVnr2ZPPxPRmiw3R/cWkZoKmqy/lsh0CGEFDQBPnLxWor1svdzZOBbklGg
YSDMNRL68exGxHp9jlg2cjfpz868omz1Ame7NuDnsf/qpoVTqAC7pgxXNVwHQjOh
zjbOexO8MzZM75fbtJQBZRN2MD2bZSh7Qb+PojxKmPkOu1D6dRR87Z1bBxjT2r2q
qejde3tfHfnYqzG2d0Yd7tz/IpTP59AHWisIeHrFJ5bEvyUzRp1dfM/JEyyjZlMW
KU4Gef3cYh4VrfbVQB98YF8fUvfcJocBvtTcPf2uxEYEsThqGD5YnVHVnEu2vlt/
JQTNJHcxfY2J8M78kW9M/IPC0IVTrQ13PPst/N9aaX1TcSKhclpxvWlk5IE+MlHU
YZ2zUfSripTmR67geRFNOiyJqAYdrtaZ4Lm+woFs/fAidyYhPKDj1FJv9CKcttqO
PZ5Z7OTJyTneJfbki7305B5G3pYIfvQr70BtEWbDHWsk4ma7jYMh69QeBXJ4ffNU
uLnJPkXRoPzLdNVQQ9NeUIMOy1YIyNeRZ8rtXFEphcV26QbG34+NEmCfjUp4gdYu
VgqxY2dhrbbpnXX/LpHsNiPnsqTbtF5zd5Yxw6Bq/8yG8MIO6DOP/KhrOsdMltbZ
JpQJAL5ryM2UUbSXhnvU0idb5dE9cGg6CafpCE4LPGPpPyhmo+Ii/lw84zZ9Psvh
Cfp3KHIYo+iNDX8CyE1x0Yya3C5/W+7VZPxxYWbQ+CAwERbFt0CAqq+3fFIx5d+8
X3QDGNhQLS2m/acpihy4FWlAHXAiXx0PzbwMEWJDom4OuOsApKwP6qGfUdjzFuAn
zH6telhNHM/iUJPImx99NY1pGebl6krELLflV2h/S2C1fHAWZ2ILmq25yigxTDAE
m6xqPc332wRFdl3FTbHru0pZu+8QAHp/CsOTZZJp5Gm9gHwAthX4ly7kMAHaFgo2
U4Y6IeFeNaYOiTxgtIsWOkkIxb6gm2SCcvUl7rTTWfVsoHf/egDHxBsHzebNVH9A
8LsDHg3Iokq9gjjhnec0gT+lrfs0k5JOsxAx0LN3LHsHdcxY8UF65gVIsE93mg3N
kiNTIsnB/Zm8B+7+E6UF+lnAKH6SvOwaDXSpY4wZ2WWACl/BPvqaB2CfKvyUuGda
jalEkELYiRpPmM62BzgMUAFhFLS8LtXIKFsHCxCd6ZGR5WnpkaMQ+WYryWLMB/+C
gvPi0wmCf1oTG1Ilq+w4AY6R168gMtcachfxKHsd2Fe2WPJ2DdORAZaToV56Zz13
lJnPQyDGzH5VMs5iV9T/0EZ95l+4mdhQxJM5x1XtXcte4hz/dw2trHwuGfLFAn/F
H9yN5GNz5s6nWyGrxjz9cdajhN+gW2hJWtxY20bCUAlhELBDW3pV76JYrQwYWP8G
gZu5NDBxYwj3hEW5wxukySb0YBGgCvuRkb8AansxjzhkLQei8+aQ/QhWm8cwdB0G
27dq/RG18UP2AznFKLKp0QQw7VfrqZzTawDnhk6Vp18VrZG6KR4e5+uZK1ooLmms
L2yYuuuD1/xglk001EDWLsWFUENr4Y1bOD742ob6v1SrpujVdKevNwp2q3WNAo89
6mSzw9A8dwRzVShn+PNFtFHHlUGbRmvDZ6NSBV6I5B+738k2ZegL88/XKs7ymK0y
mtlpfpHbth0acPAdm78h/EyHM7Y4U2yRU8yzx8QC5u1nNJlv8aqN7aPXdx4zJw42
ITSRo5P/yUbJc9pk1jhkr+SFaxADS3zYCQTXQb6CMpsr+t0mMdpw2Ygc6aFV9SaQ
kZNTG1yvCZMsiRUNGNKp47pyO8RM3//NZL/ForzWWsTn7Df983z7owLceRmFghvM
UBippdkbAbD5qyU3ieMYfIBWakry8VDq3zIeyFMPi22X+4AYwR24YXHYV64ZVA4d
cdYwU9mBHof7lKBNqhbh8VbERgqDBDGq6+J7PaQ4uDkoz/Q62+y69g1LU5cqojT7
Inzb9ZgAXOC+0Q1ti7cD82QZNrQmlaOBXX2Tqa+Qoj1RJzH7D2fWKNLpk2n9l8ib
g09rNgRpWnEPUikYs8krdZsgGU9FfD6X6TSpgMiDP6sQCamK55/UKi8tPidUylsQ
oizYN+TtT7pM++LqirjehLTJQCGxYUlECv9MBS0Wtp/0v4LoUR8v1yKUfVPsKWH3
I23+byDbe4ydO2Hv9fcLlcigAlSDnTv7FrihWbXKoZU6wExsmCyv44K1AR8Fu1MM
5LovDB1M9rFXk0+jjVweASPqGVhtrZ1LQSCYH0eXTpy19bOh5fdO/y5B70OhN4JC
tyieb8QgVBjCCg4FiyJ34vJJ8PW7ptFbz9zm7crLO+/8OUdBBsKL+/Iu/grIcfAb
6h/nFS0pURBC1PhAA79uKGpMp+HyH6I/o0cJBxQv8K2dVjy5bSbMqFLPcnhOrO/G
1HZqOBtpkk1P7zeQNhlaXmEXLXF+ymInrRKYDMWybwjDSPxhPmGGWdgwNnJwOLem
4S0l0J9IeoN9+8jVIRvfuD8pBBMNnOucge0zQS405LzWis3GGULgk0iUJcYPtJQX
NNjXiOxz5x3Yp/WEkIJzSZLiGBlAFfLaiTZQ+BGs1oJemsVa41BWvPxW/X8+wpGN
ClWQnJtfmsw+mtmNQoJbdD1/8LiFR3dBDKrqEFb3wF/jyuf7jMa3/PQF7VtDhDH+
0IuGRPXmxB79xkmkt6T3NVBYX916p68ixMrAqxxG8j9u/g+0N0RTgh2DCXZLK2Gr
8U0x+kXesHLGjxP4pC/fMkX5bS4fdFGz5k/gym001Kcwx6hy8gkxirLIFHSgTtGa
RjFSXyUlxznwEtZ9EHTL6oMgYhUVjgwU5mRMUVGINf+1WY+pESxlCAxjcJp2vuiF
s1x5/A5+l+XM3+o3esFX3axwGRZcfGpxZJiuY+LoTFVeEMAX2+APeRHCXcid2SUJ
JrtN4KOslJnDkBPGvuqGZt+NASqPN/J2cMYrdsSWnlAHM4cmXAMXXggr1CCTEpX1
XIPq69i15CsVXR2x4cs1to1sLETP2VpQ9mI26cgl8tIbAfSMlPUf6cB5yhEPkkwf
dcNVz+QwmYbQ/Aq3Ti3wdOg4IyjCKFcsrlHZAH4usokD2dCD5uQ8Ve6iOpEF89LV
9nJk/7Iem7YG42W+rqhQl+7T/+nCDF67wHbOz0TCJTVjjNtVkRBhryISVYYHjcJd
4R0VMiO8gl/KP4HvFpJFz+Y1W77bAN3TbB4+yrdLqfkh05K3O824Sq8VJk1Cnsrm
VK0uY7MmjPds/FmrdoN4m4CiOZ4NiXsMc3XqH2Er0wYUDZjuIJdEG/hiEPLshvdI
oFRk45Pe84igONdP5v6+lgukg7AHba2futw9w0BHqQDcTtKIugPjN5WIqWTEqlRN
GRsWzu7KFHBwlTbNMbUplbeZJWaBMf4Y8i+VmrN0QkH4r6zQ5cyMF/mwmNifjkaF
PcE+gM7F5W0D/NtUOMDqOgduKP44wejRzHsopOj0nMnsOoQa4TfADuagKyXWgyhC
Mib5HB9/kiYWg+vsSyJjv9q6AEzgcd0D4AuC30OAvWCKrLKDE1FPHVfnR3XUm9qQ
cIjEXij24QD2tbH2iZ2eP1uPFP2VJcWAQ+zqlwtlv/+A1llYfEeH5MYhQiYVovpt
mxvNoM5bOmVvMVQUEAMp/xu6la6QBA23EAJIh0YB7o4mhDiDL1UozVAY1pYLFlPu
wO4Hehhyf0WazD3aK2h8oFKytZGpSGYSOSl6dbpx9jgsLXgKKUpSAzn5WYUO/NTJ
N1F2iCOh4IgVk9U6bHw4ScOYdTLh0q9jAh9CsP71kvc3rPNQ2svE5Kfu0CRraHDT
SW8ARq/ubnxoZxcKHfqFCJOh0IDNOPhn931o1qiyCgJ9xzlMxmcMnUHalEwzZ/p/
B0X3K3G7wEjZgFFB4WnFWzCMa5ltgqmnzKED+r1hoISuQkUd1rxCwCdCzXrGBvh9
E2q4VAeviIdgLr4kDLyZsHNDAmYmogzKDL78yeMRcoCzsCstnIOkx6N8HLcQ9v34
SGXK8A/fyILkZnOE4twZHcBgs/HrEk/w2YWuY8Tlpbp04SmbhizxFSpzBKqihPbQ
WYRwo1HCeKsvyXur5BzwxsJSQeN7uAc/IvDvriwgs4ZBn1MqwU76ylacg+xILriY
at6OAjTJwpekDXr2MnvLwO5xKsRDNW6q34/HGctZ9gUt2y3yS3BPxvjGzFuCZGBU
qh8QrI0qf1MHq4Mn+T/0Jw38ewU6HS2BN8C92c1nb/ireWDn4FqZls+9U0BEZG+o
ubRaEv9YIYZf/B2+u3s1aOFzTpFHXp5j0D0AQuu4LxmEcAKk0DjX+nZF55F1otmU
iHnESXXkBkMu5QRxu6m/Hg/XO/XH06nRleW0PkqzjdS09VUjKZrKket/AbwPxnwm
pqlWcA8na5P6eYxkwPqjI24ElFW8/r9AXy8X/92wElKBYmEx3wAf58OrwEmD62YC
QFHR0nIcDRCzvKk0nvaCxnhh/kYINIUAhphhhDqvo8jbfLEMdVDmlkzpiGTdTspb
10WbclUFmOzGQlFKjZTFuAAHCoJGud0j+LQBO5k3RhfYTgyoq+AJZ0PBsPQHzmnK
ou/C+5hoymrXUp9HaIjslAad/ToLDF+cCXIT2AFSvk5GZHKFb4Nitxi+mRwjZc6W
Wx3ALSRWO7UdTsu81+bNOOuPRVmbhPoMyQ4HLnk+SFI9ZupF8NXb6XNcK3cBCbkk
KInOtC7VUIxLXgMQMUCoSmy3YXhQjDwMQwoeBKevM4Lfu4vDgyy1DMUzqN+xIrP7
GDHUGkpmfoSPjD/2VqCa9t03h1gEM05bnoYgtowxmZ71IzhtacnNlMIM6WVSMf83
eqS1DmVE/ExFQ1RtNWrSm/dQoUm4wFkmYmXUm8gJVJZ6YQ4W6eX/TtkOyH6Tfkv4
ZPwyhb5LuxnkPfYrvuCtWE/XzjlnFeawSCOrHo1wIPlTGxfJ7nw1r/nYB8lOzzNq
5PSPRpgvwQ42FUI2F4dLD4Rh9Ph0HwiQo2qZEhwAZMmGEv+Z2xo38bdR/Oe4Q4FK
5QPovHgRsdfmgq0aVpO701H4i5H1iNxTxkKOVDgKiMuxTxxcJDD0G5UWn9s9fPpO
52h2n4GOX8sH6KcGA+M4mo3Uqyjs1rKubLhiP6yuwxBaLn9WcdR8T/oO2QHPsTt1
Rq5o5F7kXucOkEk1qYAirTfQXdAio0jf2+TsI8HQ1oSD0GNJbirVgiibhW7OcZT4
3EezjnNxPHOS0JyeJMhgbe0higN4gcxFI1e40r7ZNFN6RvBOEI0nFsZVaYBqbN1c
1Xf6pFGftzoIA9Tj5P1DHBk8rSZOAVhdyuPNCtvaWkyvtsEssrQkEzDSCbJxcEiI
wQ8YoFJw+XQcJM4ru1BMryfsd1APm277FYOOSOxgcHoHZgJ6mIgrFL77tOqJ6tFi
O3drp3JaNkt8Ng0LtdWIdkQ2CPPpRX0vUV347eV8APiFsyr8dz7viUIXXTKJW12I
+nOM0UTj63bXs4dnlvptLqHMzxFaOcsRlH4awl1Nmg86yKmnUINfmbISObGXkh/r
Bx80NSy8gYZiWU1UO9Xyf6f3GhDLuIkW3WqHdTrENwRoQg/ODUI3MY+Xy7NrNncI
Bet79Jsby0uJy0W+RMxy+vXCsQwdFwslegeXt536aGjHOqfLaNEAs+29f0eO9/qh
eMJWRlCVAszIQWT1uyDvtpvlS/+HsGEpxuwyateT/bn4xECucU1iJzEBKNpCJpm+
hPEkmI+Pd/2aBmILbyiPsTEhnT+aQjEbjY7QBjyAfvMqrhlYj3OasLE9ELtxZ6+X
kAcobNOAmLwZR0O80aadelitVKH300RZWtz5rNT86tjohhD0jJqagqLYOd/uNXbp
4XyztQqsRgApbniJa0MrTVMgAaN56iYOTNujz+Gsmx6i68j7z8M0h/zaH0PbvkzK
CySIPKWj8lyyoBEXwpQGUC7+QeW5VOEI2i65VA/xeQfZ0Dn3/cdHlLUbsHbg4sx3
ouI6r9Lg2ChfcfHTUGZ/S28CQo/grvnO0dNQUkHkOnxCSPcQu3OOcof5LgfJBdxG
dSanExI6JDFDKyfZqdrSzdUo8IUt/EJNJqBmqfgZaR3ipj4gh4l8zf/+4+XnOVX4
c6Wvso4+WbQQMZLG350zYlESXXEgeBiYq3QXuXeFD+czvprsiqWT6YYP3cbw2a28
n1h/N0XjmSlboYsRDRDZUt0mWmTkMoznPWxFXzzkoJ4c1B/Oww6FeDHsO3sc0KTQ
sRTaCcZDqGm2YwQ/cCDn3ufH2kCn9FFxP1Hug4Qih+3zozWB3Gg3+HAOmf4joUDW
rFkG7Yd1VIKzkyuUMk0q2HlHP3hQeliSRKeAYQsOTJDjwvVxW9ZWEnNhSqdiLVaH
phfJAbOqh+qFyG8NnSMdPJzsAJxdMLWk1SDlIzj4o5XpUXw109ZbVP0MrezPQF3S
X96LS3fPeTGew3Y3OAlmOJSNN8US1ga5VaC64O9J0x3TVKsxkhRx/EUzGCSWcwZE
+uaHyX9Vs62Gwznj9P2IyODo8vECctOfKgmmvroB1luSyq0f3WwJyDtHOUwJLHCB
0tgB7CQbn7XxdiJVfHE0lHiHGeB6/wrkv+a4MGN/GPpnTcDrUtXijQwpKYwBLFIx
kQmGZaXRObVmpp5vix84YwAAph+UTR0iLeszFnZAPI5miraV3Y4c2Uv+p0lxi05z
4rDftWZXuHjBqFRr9ZCVb/uOYch75C/kSPSDfMaH4+PmhkcUAgROLLeSr1gGqLGH
tinzkHc+72pmy8LP9ui+7idPozX+qXEpPdbeQBVCS5OVF23SFU9x4AynNAzeg6WW
OZCXHhSF1lC3mXBPKxGTPEfITs672zhgoRF+Qoyc6Xc7nrZyfTKcz07b3oXxvoA9
/dZY1onTIDhGUAoxeerNRapWgOpauSd3JjWQ5IPnb1mJPRmooBSUyqQHf0jPsP4k
ElxFNVcjFfGhWRjuZRlfgLSG9/Ro1953f1SjU3GMrqbVfnkT85v7CpNL+8569mlg
GnvCfax0/FTmnGOLRvfChfnnMwHmCHOHeJH8TKK0GLv2wG2qRlHpedn4UMwn8gsT
wpSZOD9W+CRtdmiTjneMA5rPbR6EgLXDLUJ4Ruyit2WFUd3GmDKeKYYEbfeteq4o
QLtJx2hFpO1ACQ+dJrqSu7A2GK+K0DUCJaApNxOpvG1G/4phn4g7X/cJvdvA3a0Z
nzcWm9kP+H0jaucVxvKJDKaLOZLcZBxeOSBXNx2ucRaxSXJlKsM9sWvN7Meq6rxi
BB5XV6tIZUWdR7D4Co78ZMC0F7YQXn5FDN3+lOT+2avhqt26aGhoECOeG8KjtA5x
imLxHaiaCbFdscLkRumG+J8yuSK+U6qv8Ilehnss0pxKbNCphHEbLA27h5N98fAi
DT5FjViXZ4qWV2+XTykgr5BrQu77Q/+MIgIHXzR5gu+Q17TG5cIy/JTnyVJetzhl
2yioThJSdMDYTyMyebxA/qV7Lq1Ou1s77pEbZwmskFPUAhzY3J1EDFZRS5PdoD/0
/Hu+WVDW8btzMl31TidFJyX1uikrsu6fjAhPxS0dAic2XNCuR04Pnb6H4Esi22Rx
0OHMK+rXqx1lFQBes34IxAKdPlqPXizhljSCj9hsbYaZPzircBs8ESphMwtpPaLy
+HmG5EF9EN0tTw4wCpFfVlNWdDxc8lwMvjrVUi1P32Ve6hpQPhkB61UWGusZgUqS
ZPV048JN/m3qjY5GYLxuAxqOjwuQO64BGCOi5fZHWTiL9yi95LRB7TWVuXehqx3x
cp6tZJhVnrKg+k3aK3/RQbPNQb4NEr+/kNf2C+Ggf89lzalXqBgZhMPtJRj7XwZf
vMRoPEdSoegxTRvhGP6yFZTM2WIRNN40PtXUMWHCpSBgMdci73KeZj7gVD7P8Ybe
FOJfWNR4zjJW5S+bpP5FZ49KDoy1u88+4h7hBw7QQKFVf3/FuArOwev8eQcikYn/
AoU8nEFGrXBjKLrBG6tw+swzjo914xZKWPVXyYP74uMZnd9HTUVSd6zlm6RyGzDW
6745pdHIWnQdULCxLlUrUs05MCKB6ZSehWmu/FZjDvpgbZmEShJ/iJxAax2Zkcrk
47PYHWRjQGTwCxg83HSzIvlyPOBBLLGt8vkyKc3nsZ9kHxMEZBZ41QoYQEhyrw8N
81NB/hH7crFFHb3g9J9jj7sy/USgwC7YFAlhdFdu6aQSFhFBPDOoWdNR6iNMF14+
Xffcjh0cKGTpY3PmjtieQK6kJxQBD+U14di4lRehOt7O1nG05I9lQq3JENMkePmZ
UnTJsJJAH2vCnH607Nm7tEWX4pi4oCPgoZ7LcRSy0ZK2p/ij7dNS+d5nJP2Y30LD
ZjyaQmUNmthaqTuAx1fFmQYFGSlDgabPDc1ai2ZnyBdd+aOZ1gO/oiThd2wNqtX7
tcc7hXk0/1aa7txlP03lX4WTIHWv5p9KRMxWO/lZMu97x0qF1QKfpRzhumQd7k4z
pWWUMJKbHt+R2ViwhKoaCmZTyzi9R0D6T2ZZ8EgPdrR98miatMaQVDep4YMYprtv
yZ9612LCAK8ofonHWwaBzHy4TXgYJ0g6+VjTD0lfYH9K/aDbzaYXjAuOHLXDQlfL
GckwsTU0zCR00Ozzk9tRA3LGM/xuaE7ct+n9tnRjf/UlrDPUm27pWOu0D+RJkhBs
EVOnsnwQ1SPgJFnXtVOPwdhjuv+Z13c720FMlhsO1so1wzPchbcx90SS/7GVf5Zb
UIp1FsELXS/u6Ck54GkoMU7kUgp5uc+i/5LcXPT6A3CjQjh2H6gv5gdH1f5Qfz/v
cGljynBUjp8mClceAlxqiZnMZOgKipm1RfF+Ex73yvkGU0Sx3FWG3W1ruQnpbSZR
eGFgPa/+YEEZcZozQkF3YTcGopLjArjThGVeSACrhfChtCxBVjC3ldt2O4eCMbcJ
BPwpsMBI6XRPi5YUHd+3d5MmLqnwiJTN87tcNFjZ8rgZRY/bWs2HqIlTL4U4Pxp+
KsRdil/oE5tzJQmFZKboHoh3Uc53+/Rc845n49SSsG06St5he1En0z37r0HDQLR5
jun2D0tRN/OeUPujfkZR+nsG09JzByEFm4nlzhKwmsNiZ+EkNNoZuB92gv1v1xgP
xS4ScFTaMK25CUaFdAiZsfLIIOcygNy9XcZAJNeZMdeJ7qTXSwdcIYefAs2fmalg
Sb78czFE7gByGmybpeoFKJ7JI3Ns6sarRnPqAx9YjWr2wNsvnJV1nwxcPJa82nIF
Uw6EuS3s9dvqaYt70RJf1WVXRwAM7/lRAD59V/GYveqCP9dekAM4x6jAP1JA4pI4
tpfqn6gMP8KlOL0DYSM6KJKBW/DgZdjUH7C+EqPBQ/OdOJ8k2vHXRdseNM3C6tXc
fQ58jjVyG4Juqr/T78GGiarMC/wFu/RitVPzSOEMfx2C3QHKPp+L3XNGv2W5sR/V
60YWbGL+ERaWOIapyfihXZfQy6+5GA03L0e+7eTQuB5JmAZRBY269SYI5Gn3vdZj
xM3Sg7220sbi5G4r7WvXheKZX90nnHH0A+vXRyy/DN2G0Ck9yi6OkKIwNoCXRDr7
yhWSxRhlTcAurqxmm7oI0pnRC+u/E2WEfczIcZsSplIWnD9MPndZVU9IiBBmwTZ8
atpvX1cr67Z0M0CNCv20hcKq+xJn/u0uJJd25EkMfxI4eGtVKEKbNhuHMHpfu9E7
NknliHQuhWPR5MlipI9iCWH5z+98OjuVtMf4VInWShNSqeY7b+yp0k+nwcg3sKnh
NhlWNVczD+NzxyCVBMhaMS0W6wW9QWa2r/jpUKUznqrlVKCPQH9Kn5aybxa3NtW0
ywmkisnzXjCZ2jPM9p6lt08FhEHVJh1zLWGCHOOWBeQi4ngAR3jJyA1ct5kIdxYg
Z0v7ht1mUB3IbAXmDfQ7tunzkfREeJdz6KYaqJRnkS1f4Ih3T1ptPnwzT3HCmyWI
H620+0FoQUGdoTs3sDO0YC/XVU6uviWWEE4oshn+VvCIzukGtx1KVlLmrltPzTY1
R2usowPAd3Nc2O1dbhJjdTtQmuQaR3jHL4QgK7aNNk6noYUpx+De+UxqVRW9BYoe
bfpB3s+YC0eimVShEfr3430DtQ5ML0EGjwFngbDHjsRUn60Aw5Fl5Hph4mRuAlch
fTD9K3vQu5EIi45NW8d+79xF42NHLB8VwDb192m2D7Ybp1JlwVRJ2a2Y5SPamaNw
lKmAE6XtpSPwsUnjleDSfU0bRlbmWbgeiAXlXCsQGZzySnm9eXxryDiahedXCixr
Q2JVJ17bWDgeva/WWj7qphCanJ9dRvF/jv2NN6BaguVWdIcrOiO/S4yqXaY6TupH
Ow0Aq4HHEzt/lnFJLGScSLqIwkNGaqaain1XIaEGYfv5Y/TmtGUOQ0u0GlLqppAd
sBw96x/I8KBtaODx2rTVMm8o1PmqW0ogZ7vCioWehg8qAGgN/qapzg9FsWx4bY8d
mBxk5BBCmO5vq6Bl+K+VnTXstzeUWjA911FzWHu5GrqajwQzfdAcVCa0uD0jjruh
WAg1lHwWP8Y8x6JI2R6ZADOqZ/pRk5GqAidEdg95txAO+Ns+lmRUPJspHeoK2LwY
mlBT9tBN7cnPvNA4wOwWupFdTolr+pd7CKzM1pC1VmY7VFV7ZeWlOZgFcbdCBPZ8
7YShc1Z7XZcx6or0ZF4c7H2SMG0j6zlIHjpdCfdpXBpjQ1pijb1jjKhssAwrmgxE
nM9TBOmSWtcCfiGGRbg/tuBr7UCekDCksch7NqvksDjzjSE18adotucLHDT9Hsi7
fj4XBLzKTAiHtI6TeYdBSWgM/P01e7jGVsnMHJJeZZMDcrxsmN4ok/aXHVp2BHU9
X8Toyewq68aLhpNSuH1B1mSjuzS56JfubKLLL+E1H++M2WP3KWxMIN9aO0gIaVbz
suUdFvXbxXW95JC0UZ6Y3XWUwyfq+Acc4j9mccM20EUJWYpvVzyUbo1sjlVFpehA
kgDR4Q99q1p6TzoSY018EO1n0sLhMe5NhV02flNGaGsT6ZP8ipVtg0aPj/0fZ83z
MApSVpXyP0rMyhZjSl0Ya852KHBV0kLa1LqtF/YwbIB+W5yNvAnC7avhmmxGpAT9
22GW0XuqM5/csiHHZczC5XaumlbAnPdF7K3UJp1PoyJO7LLccDbfDLqAaw3hVpmE
KlPxVrtxTwBG7UOPATIeLlz4xVtth0nY9qp+KXKqUduM40crfpPAK5O40nuzIuiW
/kxch30l5a5IH3aYQ/Y0ikQt1Xwr9cNhT3Zm/dwmghWPZXoI2kHJx2/BNHgz/oGr
Tr+GMWdlkRWEl3ZoCtYFXHzKgPYcY0GREeolORLJaMkyw3E24FgTIhl5Q7SHpEe6
e/6/OJn/NGKYZz+08TdUROofy8QJe2pdaoSYG5ZdgcpukgpEQWdgi/LeMDT9j9H7
v+MYJyW7GST7r2sCbu/Auu7gwSIqAC80oDzBjgUF1MF8SEW/Q9mgM8KYrgUNKhRb
J06CWb9ot/Rw469wWRf9lAtVdxIl+hNn6VMTcE291DO91facIEn1mNA7hfk3o7W1
SEkeg0xqKa5m7fEA4nDoUTqydMdZjDRBuOmgeN1pdrV8KQ119M0rru78fUWv/wSd
2Yn4zpnQTZcAWyQkMuyzmT/5fxsjdcIPB8OvYZyxo4qgAD+sAUxOesBAK/JNDtJb
qqXfKN9V66Hl0TNJrSybI62qpjfZayhkvvgXCU9i1jwuWHw/kzhYvLxFicYh7f4V
um368OaVLRZJQTsXonMXJo9JMsWozVt9fuNyqDFsf6Xl/fdZpMh2+FIsLRoSgTWp
lkk1Q8o5sndLn57Tf8zom9SvAnXP2uZYnQNS47iC/zRIPXvqqnsUx4KVszWWy+b3
Pvop9RUyfULkFygFjjvj49STI65gnzSfhtrCpBbOYb74/+bSHO4efsBBf/PiqYhb
tA+InA4yUd5qmVBEDVj5ocDmbVHhDXx9QIqdjXNIU2QE7CTZ4XQsevOtPksiEp0Q
WkF7C9idXgiRbPk4VVe/x2UkEKduBUjAlgNs/HCKWj3Qjl5nZu2BBrLfl1ZCL/bP
764kyxXfA4lZZkWrgtPsX8BsIWTHh6TOQTb9zi+2jShwKnwGvZ3QC7x/9y2amcdX
zontQaybhRtIyMxCZWz5ofItNGNd7oK+I9LDtxlREclLkLwUUmgcsbPin32HH7y/
Om1mjXlQLjep4gGvLs3GgrbY33Y8d/ui7MfSFwZfZnbU+PT7BcNBR/76s0Y7gG/C
WIU1ZluBKFzm8jbEEkQBHg0gA1N1xOBU/thuM+rE3pi19XKb3U6wQOIgQU0znsNn
zZSZvvHrtogXEHGWkGoeiC3n+ItEdV89oJxsD36ud+0f6vyIVt6/Hr67awEQr/n0
wdelx8DuGsX3OcAhTk7pI87UTdkSAYiZ8XHLwhp8KrrDbofgvIKYZxBU+XtuJE+A
E7defnNR18tFtlFBzM5bl182Q4Td/e0ocwKanvdVk7Pd7U6u26/VPG5y7O3JUTEl
fRxSSnH45JCh1QlyWEF5770D7bOQ3YQE5gfG5ywK0uC407gd7MAhaEZ1tpdCwS/v
BL/jzkAFVAzMI5UDHtV4CjCNDY8o2AxG90MeklTaF8Qt1WI6JOQjr8yJVzCUK5X2
kvObtUgmNFU0mtJ8cgILF3IS+zzpJuZIgyH+vm3TeqyAoizFyyvA1RSWbYIXLO+A
pdGBZDBWJzJrm0qUwABfd1uQBj2G4sVO9qPMVCWZQilLtam5mZxxL26oEbFlc834
Oyp72YsBXhUrir6xdzieBdNO4t0q1HZO0lrVMDVn+A3h01ewEdW0tKoB8+fdLf4R
Oa5yjqTBtwamObuDH6z0d/5nXl49yNzXQ44GxdzJPNvNNCSBDoPNnD/k7bdaUILI
fz1NUH6XAQa+e2xofmKhQ3Hf+ZMUEeaEZvuOe6fho7lOOMMS6WXCSu3IjZ46N3GB
PfNr23r0yq+UISXQMzTxarvjSi3mLGUr8Kawo5bLtpiKfh7ZkUFum/uXtOXdt+l7
3or3iPJ3Z1wBRPgOfru0NPRFEfnsd+q9DVTCHx7vHS289f9miB1fcDTq6KtVbWXj
PMd6t+tPVE30zllKJ8RqD1+E3zB/ft4RB+eseS2/VPW+XqxygWVgFqPKFXLnOWsb
Jl0ySHVBvYQjNVvLEhGZR2mE5Xa7ebQ0keWeY2enmJRmGKHV3kaMgy2DtmO1Y+SW
9IqL6xmpBUfS2LozyhHu1NCSwQaiRad4OQs8jUAsTOcIkpRhk673NJeLBGEKdQjk
rcNA3w6asMiJrQPC3tlmK3Qt7tDUbyTql87FC9WTmID+wukXL2Cr0FqctEKydBmj
WF5+5XmAn24lvPgTKku1GrWuvak94tOYPmjUdx4p7YcWkvZLz6ojSBv8fp6DPaKS
wiKs7bKR6WKc0f3HU88MLqxGypxIAEIc+zbRCEs+lvlOqB+oKbVuCcVgpqI3OG7q
Y33s4EshOMFkhl9daz+ksf/ieyZ0K6WKaok+Xe/FM7H0ZM2BZh4CPHF8U/RI6fIv
LHiAsHcum0RpXgQ+ZFgZRlVVw7BI0LXv9v49o+fX4/4EoJoHAENaW8wnmrAVcCiz
66WeAATrT3GYaC0Hs+3PWlDeAzjBG2UWkHnVcoetn7qfQdGMcSsiCi/XsGeVZVHH
s425vk7lvZERWwD8F9CSzb+9ua/0oefZa7Y4RnwNEE2VttJOSXoGsWaYFNXFNu/d
Pr1ZytyeuqktGs1dBvLfwa9ZnIBpgeCrn5E6HY3KcAh1Y6/SLWuFabsHVXhCMq13
O7ARTlA0FiDzLGdeYyVKrsDlpBvsx1YWKGPCpugu5SeLIeMEr5Xh7usbkZCdqQKy
GDTRtSUYHDYr90kPc42Fcp8zUcv2SBegCcTCf6PngMhPXdgUMEuuDef5OZqFNTCJ
++XIRFlyenpG1m139W3GA/LQt1QCZ/ZoX4dTmtjYhgGmIFhbQXhShS0yFuczHUCu
PwXtwwygjbNAnaOqZ6/IP8FgFa2e32fTYbwgEX2FnSfQfhw+2qY1bczwvmyTRNX4
4vPszCaqEFqQbFd20Q9me9/cMN2ZbzShAULZibSl+hLKZQzoejDhCAYHnycje/Zg
3MJ0XpCOqqswQoWY4xUMOYY3ClnUSpo1DdZbkJvquuK5dWP5eAewVwGjEd9qqn0u
gNRbYFVxuh726yzwUY/nxFxXmHjkSI4EA9iNiojfl1lcDFpemxaWAtBO4VHAYt/U
FrI1ekzGB8uzzlWI5PkjxRY6skdqmGWk544lzmmsTmXfVBvhvDX0s05BwbtBVmCF
yiy4gKcoCubV00jd7TVzV1Px/dCbRBAqO3a/CiWfoG6wKd/Job85tpNEXQAxyB5J
HWiBNRDDWKSbkuO0zcbpxXiWrCqMgq+BqXi8QLHF9sd+I7mJKyF5C6EPXOjJFb6f
eoyloopkLxbdYF3Ahiy8xEj1rYnBm2cXt6hwbkWFrZyty1es8rgTeL5+40W5OE8v
lp00EGSL22wuQg1pxtv6WvpUdiqtLajCzW9/jEySUCobhX6LpIxZAzaCN/2fGKoa
6bnIjk6NvmoZ/4vN9YWPgMneeoR126DXY6AUmeOeAaoBPA0kXT+i0KnGuuvzd9eR
Ux+U30JDxGecv3i9EVNhVJa8LyDnhTbPeY6kZ5eleNX58gVdTHHLF6Ee1FXaRQ1O
lLFgXjvIm2Lr+2Kj4+Nd0YKM70/KnTUPQPYztDfAt6kKLjkAaC/MQdmh1mhOEj70
8GxofDpJ0MAWzitt03wAVgqs2gY7uV780F4Tskhf154zbgVQ2OcIJ8ae5Bkh+ANI
6z0tIVbgqRQqwLi8IVIppFYIrd0T+yQFtmYAp2Kndp9p/+LNhoHX7Ielp2WO6Qjn
CD6aQKP7m/8Tsm9K5R46gzAzmNU4C4ScqER1VZnK+CbKf/bqO6B/f6PXWIt5FLaj
3fWLNJVZzRCyf41iUsoSOtyOYKvzMn8/Ltj6eoaJTeeQ4qdNuKtasQrs1XDL1yEB
36fLpgq1qM8fJNT0ouQ8SJcrrVrKPS+d539OE7wWpAF2OdroiR7ZET6hyjRhdDcK
v2l6Ods+YzLVMuehvDUtSRJCEenUnIA1MFzj8nMc1/BqX5jz9VgFmJQHs17SKW2o
hiTnVbc3kSJ8tFTATmz6dO3O6RAkiEDiPsNpD+mBHDO2KKcvj4FmX+SsSsIYsanL
DbVJIOTSgQg+f9IyPK4OKlcSFZCitKL24KGg7mhidxcaVqh1NlUjbu37XaPVMKPp
ggaVmVu9MHs+wT5JPRKrbN8RNvhRJ0QcVB+aTGg5cJ6+NWHsaiq6hpurQQFnMrGQ
okGhd1ruCWoKq90Vi133HEAeU1gCANvZw9tRxkD/LRlxVaTZUpO7eKP15xJ+faTS
oF3B5h+GAu8fiLkhbHCUVqqI4oCwAVey4y8mFJnrqgqdbWfr//mRWJksSPWb8+nA
+QV+Sx0AGGl95XM7rZ2rvX+pa2MPwMTyixJslFOdq1XC4Y3oMWORSz1esXSdLXga
J6ANmF01xk+Sdw/xFPSOfkoPlLT8fH9vBGu4Up4rCyWviTkQD++Yliop/Wz4FkLI
6ekYT9M+T9g2Ornm7IOAHyr8qAwxNpHjAmGdECpM0tQQVus/9Is0xdbEW5wj450h
f/b1F8Ycj1K4j77H8M+IraEOX/PBW5kTSmMottFXwJvVx867qjDtqLmoHn1gtAkT
mlm2U9/PxNYHOLTmaukOLOx+H3Q0uQbPjwEux2PhdHFlNgNkzQeqF36f73alpGdS
jh2bARaxdZDaP9/fek6hALmeJlrXBRcJZXG+gX7wyFnpu3irFGM1Buizhn74/c/q
AN+rXJkMLBrhTcKwxwo3yaQgrAyjDcam222wD9rfOfF/HxkYtgRsDpq0gSLnW5rx
KlTxWX7cbeo/jq4GyFsIA7s3yQJ6xc1zEvks5cD6FggJtx0ILRGw9G3T1mgUI0qd
twPTWE0V991K/wVmS7/dfS7ZN3sEZpYVBJH3D8YtoDaiGxCrc66ORP5KQ8g6CBnp
z+e3z1BlX1y0vB14PmogbF4kq+7BU1ULrzGmfqD9L6XPEZ61iT+iCjIC96tHC33X
WYXC3E0gf3TwPj3FbxkGF2bgs0m5JBJeRG4g4b8m1K1/SiUprPkXJ8P+UlkUrv5x
bM/pNR60tKhg7akMTtfgbrJCltLBgkqCwhowW1FLMfr9xKYQUfD9q7mnVc3Z+KdH
vaM5UWSbufnVTyniFzk5IDgEEnPdY9V93bad03r9b3NZErM0rATdUgOccC2szT2j
qrZli2tWT+s7nsA5QPWQNPBoLlRkEb1UtY4A+ITMYZHO4TI9yAzk8mLtHuFpNi2/
mfFGuwUFyL9EFvdV/P4BWK10pcWVUsdXdn+t2jncOzKbenGS1HUIZgCDTn2oD6Ph
ynbFgS8H8le0vCJ1Q6aR2e7Z3keHRkeh4/P5kUWoB7SNnuu3TFscPminZqAyTk5k
qLakwV1px/Lt16GD7AZuHEFEZf28nRJlrzKAwZPTJo1m/Xa08CV2hRMoOMYfBaPN
6wxFxwhI2QFJ2fLPtsnVzhkK2xKPFeOJKBe09QZJWSX7IncKVUyaKKmcj7NLj/2k
mzLchs+haUfIoTqB6SASU6YH/2gnQmjTL7axvDdSL3vXS8J/9clN4tHDmLRKLMGB
iLZ088kYHOhMMPvIFSUs0oN+edf778N7XtiRvgFPVsV1oxHrCybaRu1SyevwUwhg
NaAP+5b3rQB/cjHeDQZLhqbmJfJNe57BmG05pEuzsBPeNF4IM+u4oLaq+9OLS8ei
T8drFE1n+Zq36Drk+Aogrd4uJ5GamMkdRzIt3GFtR56IGzkoES+WtiXn5bD7ANjU
uv9MVmWnGTQLo9ElusRMYZ7DqysPRTOxABN8TAZH9rlU9wT8ejPqCQ3fcbGAny4C
fbP3qBlc8ZweO7T7VsU5biuhgOr4tSoMomQnMT2iDwEW6k47jlDCgoJu8LeWaBg3
bQ0K3Qhb2id0+V3FASRXGZVIIKY7N3OcqCLZvXxd6K3RbxtWWR/g5Hk66lnqZ0Aa
1K74exTn16LJ/1oTaiY4aNjT5nOlxDfFPOMtTKsj7LJNUbxihWYkJ6ZUUqlxEK7y
K88hDI5v+Iq0xUF7qwi4EnLm2w5F0cxTQBr7P6aVe6WXVMeyClahECyEQonO3UKd
ipLdUalheCiGrSN+o0dGFIpptjDShOskHd4TGNsW5Nu/EHlNjIGM2+Rf1ncCa8cA
8Vlgvodj/ze1BKhu0vq/3P+5qKL4CHL+9xjavZBYnU2XYropMO3mKShFM732sWzN
loKX3ff/l00iZMCH6eOHlsSWhwe4TxM4uShBe7mqJJBMuEedYXXyCjSCS/Aelryh
LEPfOwvWtM4isHqBnrC6LLeTlkPSFAEYetVg4Wmtbkl8dNEJq2loa123oOJwhzg+
NCaD1m6fDpBelwIkNmNlHHfkW19KThIYOFlPR2U4r0onWoGHgPYCwqoOGYWKLFly
XbEH8pKwUMUqMVZOvcIoZ7+v/nG7QqwTiSVOW6zmUxaGimWApITc3HCrv8qRQKx3
EzK/W2yb4Q5vfnMzQtTLLJDv7Vp7vJ1IbC2AW/Q20ewR9nAzu6fehHaF6C9cQtHs
LFP/Z1eFwC6OPcfwaoiturYxuvvxA/1vdWlu55np0aEK/IV+TYzrJA5zovzFRPEB
FrkcYU839NgC3I/GKMh0Y5w6+oV4V5bEfYObcUTrI1ldFggBTBhEOIUbtr6meLs1
KR0yS+mNOhRp9a/Qu5HBfIm5yWeqokV+npEsTi/k5vjuStNncZ1JyWZZF1Lmmjqu
s5uT73OfJX8lndgxDrRFq9iIpTWKVb59w7yqNeH96Hh/ICj89d5jOXsXf47ZSfy3
ppbsiq/GYO2kY9Ii/8zcyTvAxEyDGRvZFkP2IebVu159pu4wmfRts4jLq+F14KlN
+dpOl75Ug5XpWpEEYlzCqTRA+QXOYnF1bnTBAxdUNlzk+6alP3lLdi8EsVtlgQdg
IBW3cwA+f1pOLUkF4Emaj/zhg15v2dzVuW0+o8jfkivZWY+tRoJ846JXYAI0TKqN
qC7c5n2r5b2uGj49w5fpez/YnoSREhbB7XjO43FLW3ySQ4NzNS76uqKy0P7x2fFA
1/Bg7ph5dQPuhNuaXxM9CyNHITia8LiQ2bQ8nGKW/vxxAYW+nPTjAFpduAjN9HhS
kxIlc75gMZNwFZ/PE2AnHTTlLWLVO3D90uZ7VxGb2xZtSYYDA9XCRo4ewCAxrIIc
dGMDMaPvzN6gtz/9cS6PR1NMcZld/rKH/4qxBFgaFInvWY1/MJoXu9EWqx+X8vQO
x5gs3N1AxQg1tIiLZ1fBa1Hdm+ARQi802FD4TXTg3SLHDo+AT3ccJgPWZhGY+xQJ
SiXYR6g1MJQ+lgu9oPfCSEGHVOUUOHg1Ci600bZHuck2RIkMIe9sIWWtplPSZ943
QSJdXdxl7COorGCvyTajxBw4vrn/T8AGeA6uz3C36WTyIjCut4z+wFENZSVEZsbw
vbTi2KMAy3khEcZa3MBemGz6/5y1a5wlzwt9TejSWUHnCnGsb7Qq4v5gS4uhpAHF
mAP+McrMCZz43Z0EK0eKBuRhh+hjcHf+2EQRZwWdxHqkRyLUPJho2N9bdck3Nu9l
Imw6HibxBZVxWPVhewa+o6ptQE9AbcsPXfXO/VreVhFlozHxdM+5BxYdJH27ySMW
slm8tjXXLuAxF68aYnxiWX3O7q0PBRS6YHBYq5TzVqzYTq3Ovnxsue8CmXsHMT2W
jBiojEGS4ScgxgNMcS3LL0PvrFWwwBGr8o1CIgzDiLhfh9CtZz43wN83UfCYo1Li
brWhJyA5XZzeunEMh+epJIYY57CkGn7FI9Lr0t/ZHIMtjRH9tmpKZkzCc2s5Gtoc
f3bQ6/Xq6BOQSbMHTnOBGEjIe5SVvO1ZjKGane69IDCLpZ79LZ3Ssx71Vr3fSL4l
WZuWOu+miLl6ZTL2skpvtWlXxtYDF333lmmpoZlm7Z4wOYU108Ag6WMGjtk8va+Y
qcEC6JBv5W8EUqrgocCqB21Spk/bi3injgvAoj31SePSYpRt/ARqbSdIGawQqz4U
huaHFZWdeksPwI5qSJyWyvx+vrlo0u2+Evck16WrssPhj43fSWmKoX6lFDlQpO+W
oE/qPpQvg5mjXc/Avt8cWQEMhSwvWr+eUsCOgmw3kI0sKn2HwIuaOfTvWapwXZwT
AqxH2pI6XJTHEKLGDcxEcETQevafej6aCPI8tutaveJVXwS4biGiEPu7oG/hK52D
NrLpuMs6z+qh7ul2DJDC5q/tEZZ3EiKYHHAc8rzkJMPtgrZNEzE5MIM9qnMwqN0K
Nlz3xo2xRPEt1u4tbYVB4kajo/qnrgxcdvRFMSQF71KcJmquxT5a1WZKIS4pusKX
a5D4IAzaRpTf4VQ29AA5h02bJlLc9LouqwFOqvy/xqEqeNr9TyctYbhYmUiWvx6E
harUkQWcrGhZXQoi/dq+4GL9eptTwDS6NTH8BMbyQW6zFbj23PRqE4SsYzlSbnOB
mPlTXAGbq97bTL7rhn7YYSG4O5ZMXVAw7jpj9vSZQ+QgQzkGvnagWi5jAHgXVr05
aJaF1+GID2Cs3ztmekXHs7vPJovPoFbctbpF6wy1muKcw4lKrsDPwWa+rBe8QOWi
PIVqA7+XHa912N48VtT7m0dAysWQVvtYPtKra2D03ywVNdaqbl0+OetGprXFxSqL
H/7syc7X7S+nUQW9duYUkN3QqAfymT4pztC6jeBDPEGArIKIfVPiDs6CrNuQzKEo
GvbRXmoCvFy5NZObM780hpQ6+cv83e4PoMGY7I1n5i5KTQ2HW93RRz4uZhZ+3tKu
ArFEv3w6YnJZUxLuaBS5ypqmuakrGIfmMsmksMIrXpifbEDC1PoTr8qNDD9KeZSM
jT95+Yw/TkI1VwLNd4G6dKtbCzk2ngfKaJNH/RhOp91+bJ148fDt7jxHNhx/DUO+
f3ffvt9XaGyCtiRgw4F/FXOCoudx56Gr9R3zKqzNYSrJYs1anGE5r+Hzb2CA6g23
E7fxkw+WxN+OFXI0HA8I7lBKkNeXSIA/DPlW0udXolVDfkjWtH9qOxTYBdzHe4kN
0Xlhgl89GvxGMzIrLV2yaDfYp6ilGRZ4T3qkLISi2vJo3Q4pQdksjjSHjpZLBPE8
pf7G7D2kEULtoICXMnJjzaIhbvBromaXlcukHWZmiky8KznSS7wG4o47Y9IvXall
RKVsH/MWacELWFlIGuUvp3ftB1EGVfGQNHyGOsmbE7anqW0JeRyN+7ybuN7rhF5q
jG7uPw/DaxV1AfZeLpNSw2UghixR7jrc1N/laiOlxWNJafYLDkIKNkpna/DE5IaE
W6j3AfPsBnyjoNBbDy5yT+9DuH89yxmQrMuvj90Jh+aKkeEGKYuSLbxSO3HJK9ob
Ho3eoBb34E8TDI4qq4mRyOpV2HuQwtwRZgsBTsMMvWRgEyDFbzDTxdTAPdSQD0ra
EnhSicWCmeFKMtP3qbrgpSxkqMqm0DR6YIia/CMQWLNlsFUCL8UwpO3d6CJUwhwn
VIhUbuT6xFTkmQTMf/6UuoAB1PFjnT42/xBrbrsAHVnF0MkucAupl4ORzizl8Hl5
Y9f+S4XMm2Q5eJ9RXUv1vYo83Jbnq3xkZFkLOjKiadzOEvlX4hcBZbDKT9gZlLlh
pcsMvWQ5zqKGSlzbcBHFyXHlFTxCnhUcrRiadl/m3RsHAGi5r70f3NnbN7BjQ3cX
PH6FQ/FcpPUrIsqYXwlSzF5ShLgLKmjlJtGF/iQ0pqkeeYDBD3l5OslrWJlIQgRc
HdbXRu34AXlDXnpakh50zKzdXy2uaFyccOmIDRog2o8YlOewQ8HN8tBHccUy4SQ3
6vRpC/XDlXYjvwBlEMDQ5NFE2YaSAFKqjeYPrMnEfZGT+Kt8Ata6vMCmz8I80IVx
hJjKPKJCI1N5j4FGYIW/kZTFxIukB3mglds8qe9teJgjF/hLTBeb2wHNQ5vTJ4nr
Zw9y/qy/UXB6mdGUFbxNtwX7xTM0Hqf8GDpXvhJS5CycvFE6CruGSy40CX9dm1bs
SuD0YlH8lVl78HSJvEnTOrFubMrLV/WI0ggLBwZc/qSIsTSQ7L+WtyNj9/Q7jppP
5MYr+Isi+Wbyb7s5yLsHAbg/cn986kr2NXqrRbOmhg3FyFN+I2fPLUy0CllMyXY8
c/5VYfUS7bha8jb6lRhM0gBQBcoOdpGytndL19Ujfo6oD0qifWoVAbrReOrU8g7W
FTk5TtuhQwt2K2cqQcbRJLrEGacaFDH9Q0qx+3eq9cPaWVZPK8tVKIYItm556yJ3
0OLVK1/sNCGOgt97DXAzEwjvEB1rnnAxmLHXBi1EPnjzy/qcuy7RdWKQL9Himvrj
zyLWhiTPR+uh0z0q/Vd69RKn7nxenExefiR+ozF0Fsnnc7VX1Cge0Oxn75XG5ymW
6jmWw/PfWEDcDTCQp9SDwZDUQ83JyCba0Te4XSvSLrzBrGrt6Nvg7PlfPLd6lVLB
8DbQgb7L6z5xDupmOOh9qOIyJc6L1Q4WwgbIZTqojJ7NXobD5jry0sCHe58Eyezs
GjCmBXr4iyjTZDRubRiPoMYMMMDIKlkvKeprzoyw5rwfHFDLZQpbYBubaaIcb4av
61B8OWGcTyOqeG9/MeJVFlp+KhieWAbnjv27qydySSZ1ASDjwFq+npxYCHGVH8zQ
6xiP1CfrH6iGp8wRr3EHLXdr9h+pLcfVMEeb+SedcbaM7WG6EmQy1R22Vhj2mRpg
EqDoplnDTyCjZ2q2i7xtMOV3ji5Vvc5itA5C8VcVYSr3Rr93JXcF/HeSyoUTSEyK
io4GuzAKtHeFFD0LIJiXfdYf6cgI9IuX6uySwmLdiD4Gw8xu5bKVM0YXI629+FzP
gZYJyjpgqZ7/oFLuBxdWOiT1d6ZiEnXitM4Z5bEEGaneQMDq2dp83eRspb9j7KRN
ZwD0ACrBxgRgYVYDerTfA2p1U+zhIHydugbEHn+XH6FfwWbYxPDTwQCUGe3dbPq9
XzqwNFoF0wDKSSGgNzy3B4m93NN5yWG57O3+c8R+rJ9M1/exYTP4Uun0Zp/ltbTz
RmZN93kXVWVCM7EpE0caLzV63Y4SUlgXj7aRme21ui0X0pYBoTSxx1sLW4lmbKqT
WwRT3vJb2jmdV7uDHQfsxs3FHQRT7YDmVavn4p2XlieZa8KcQ4mX7iWcJAfXg82j
Hb1XTmDgodbpKus48t81KRxZqGWr5MHW3Yxr6egVi3899XYDbHO3CGahm5lgbMzL
IwCcblIn2f8HjV2W9sfYqI1C0jZUDBmo2KQwmu4IRixrmCZDBr5T/80PqrVUL7yc
oGf8psou1cRQ3/2K72UIodlMnPfNsDautL8LTbv9EI64EHBoFMup4Me0IArTCiV5
xYAbR5NUHhsXWjkkAeTT+ev/XVpoTVe91CHi8Aft0QIlod1An2CU1YuF3cBBFSHG
7JDE9O5099CbmCRHwc15S5iQ8OwgyoNfXZ//Laq5vwkXp61wwe7CDZa3gSR/M2Go
tyq+JywJyvqsc+ehZBARCTxqIbiSqdMhr/NH9gLG92sSCc8Zz4BzGFFWtKXDM51K
BkJoq/0W44RCKfzAjQLj4OYy2ZP1nHhqeGzVhsGe/UcJF22Ra+swpdOmrUCd+90s
pn7W8wPNTb4phbFei1lqh2njR5Ul4708DMyZJRJ9Z4U8RQX+9mdD0o+YPNyezKv0
VquoP8xjzK0S+amVjNOlhpRZKGO3cERjKb3G9Si/GQjnf/6fNi6B9gZphTY0yY1Z
cHDEowqfHYDWKgujiOGCBgoQkKizaaOK6+bgG6ell9WZHXivBUBLCRdnNtOX33XZ
Nvpp40ZgzwCq7ADvyyFAwGSGp7eXo635DXqyR0cqft3AD9WBjRv97nMdDFFq6YPr
cPq1zUB1WJF0zwIXyjfdtMwbwPXCUTExTc7OaqSzTVwD92xzZM3zSmaKHZhddSon
ahksb9R0GIpl5DaCR5x2i9D8FmNCdtrYrrcUuU++S6K2FCYKl3ZEBtomg8OUWR3Z
Ofr508U08ghAxnE2KT9ojvqUK3+TeamiW+17ydxv8yG8XUPfkcicHqs9vZn56Nuk
i2iVmxSK993Prpaj5r2z3C0iGg+DPfdugV1ZgxpN2r+bxebuvxk6+ZyNafypJ+8x
Z3yYfAT4VlPGkiRaxkVvyHU2qKZYsDmQP8u9Y5c/Zihb9OUUFMEdP+s1vMtP2x6v
sG2MVGPyYtY1DqprRb++tWAB+aVPbuCtClqsGA4tgqXa4SfBxLw9sAcXxQvFEj3m
7UwKP7RB2Dsa7e7wMn7TPnzQtDZmgYAAeEy6WWjhAvbdQY3kKLtd3yNOF/pLgtWo
UVUHTw8wsi+Ve5xlJGbM//DU7YuDzasNeDAkFAPrPOGlevbB655rOuurm8j/dFf+
40Zykei/h/OuiJjHPJ+IfJzZX5N8vU6ZChIFyABMY/3eqGgXtCkCSxhQKOXVRN5Y
wsABJfFqBR3DwD86Sy/IdXXM5CvXpnIUVqxD+Bhbk5m1M1PbsMfoMI0B+oN7EhBy
CK82Blp8TQuKvXty73T2rxTqzCF1TY8dAxOxOtUMatFFXD7KbVzOk+nwaONURQ3u
zKdwzCLg5JjOgaH1EedwEMNVO+zIcuWzXgCRBxVO4kzipuBgLnGO5Pm9vyKU2CqO
hKRLg3Pwtgd5e3II+DDpydvPBvEO5jAt5LPM6AX/+HXp5gzEBr6p09fsk2GSNwhs
hDPsa/fyi177tO2CJ6F8gMINNrlVJkl+7XP+F/r6ArjRoPEBkCNbmBWW17GaYtvG
WQXmNNgKSBfY5G1rJdamekQ1Js9eywoAE4w/n9/WoW2ih5hRq7JclCuXfS+5avxr
S38msHVWR7R/Wz5YxCYE0YsjZTGPJ10O3OXmMGTYGMVWbnDRRnFi9oW/aDviajKm
WsS1GPv442XeOmMHOGP52TrZMTwN8EBCIES8BjcW1Mh1gx6Adqw8+Z5LM3XmNPSN
kP2Jmm1CiP5USZbsOiZTsSbB01RMXes5XGTQcBMVT7tg+WzvjfT6u5638E04epvp
NJq7iXXCeNkoPfMhT50WASoJnkq3hI3QBoYQlu9lGWZcApj1V5yRb1YY33L7fCe4
1HDaOVsVzqmakL80371UybgqsCIO+mhBiGEAdy3cItwvY3ExnrsEaXf8ty3OZi8J
feegouhrMWaGuxkUShvqF8CWE7hJeYDjl2RHtI1Gapq2sUVmDaCUPa/6DjY4IF46
tuStgWdwHDquj/xY1Ib7vGGaWvBp6nnNxYXlwRO5kSeUyw6B22Nf41iq7WCSsIPi
23Sq7VTaqziteRtT49NblZ8CTOVVHaBM5S5nfrSquePrD0Jywi9HGi/zkcDueqAl
BzasWtOejjgQAvD7qsa6f+4NIwpfR02/xnd/yhhimxlt72Ykg1SBTKZUMRhDYz7h
yRQSsWBt50fTT11FqZJl57zf/MbVZgJ5aFnTZEmpXsrQXPIQiXQsYFj4JwfkJekM
vyJjPRe74s5qABFqsNE8ssIoou7djUB94pqoWaPnnxhM9dD1U+fg8Ml9nz6UP5Pt
mf8eAfOpZbbWgAwv4B3VbyKFcx0hUbBfzHBvf3xymvnmdm/VbMR/qIGv2uBV1Qsx
8RgpKBPLaInr4TcX9AR6Nc9mSQejz3HM1zZ7EF/k8P13QsKehnTS+j8d6ZIZ2znZ
Q/vb46ncfnSGRyeJ7bxNQRN53kzpEpUB5Z/1dpz0qowTJH/qYm/VM3Dm4QNg9Q/M
BMOaiBsuxzc9uxczxGzRU2aWhD4sqMVU+NSyFqkjB4o4v77xZ+vDofD3Ap+60KUT
zM3D7U6bFtfwtiIgw2pcu+SXdYmROocqnMjBEB3DBzoYKG2Ptj9vG4Heia4zmjAJ
RVAjpzcGkGLcZxeL5ygRHFJbCnt/o/zEAph3qmoaYifvP8lWM0hKeALrvL+0dFJK
NLJahS+SxNuEy2C5KrNer1V4z0HRKOcjV+Z69ErXYlM9O8vE+XQQkMl+iDiqC+rl
8rAfIRjIQKalpsvXqQjW/9/ZgV9QOfh5tOa36bRbYyrH0g3m2DgC7zIXKWSjFgRB
SQJVoHrYzq6jRifw10+MS417acv4Drual46Py/MHStx+KA1jk6fpnIaFKnzv2yLL
OlSUle2JI4KTzJpVGBCKP6W8ekq/wQxp6X/+EvQRZ0M79JQw18jE41Yn2rmVih2J
DRRlFq6fPq0WBFfLqpMZQ74a9jILq1yjQ2GreQDXmjlb/P+5YXVccm5KDesEn6vz
mKNTvIZ+hplQxHq6tbUMIfyQFmzENnQ2sqqaBYB2P/FvlI+Tsl5sErq48KN/O8wY
bS+KaTgg5FYTCpoPN7H8HNdEv5dxmpruvRCXvagYanPOD0eZvY14IZOcfzjhUXwq
3FEn3zIQ9w3Caxo/xY09i1QTLlnUGXToaaFpPe7UiuwZQPfAcWW83zSQI8Ljw8Ox
5JkUgMpgCngbXNcmDenejZXncjSRc0Mmhom1Nj1uEWq+81GIJZKPyzvtgpTkz88y
bQeuEODKSU4jpWMBcoYKU028CT7n4OMPNOrNpvDUcUFeG2GtHax2D+bZ3M3Rfm5R
QlmjUbu3CvMpMQX2C06dFyNiIc6PChqLv7W3RKnfFrL59GlkV5E3/a/ljL1ixHAT
VwrF3TUJt8cY6WyTj9IbSmTLOmON7RgM+FMv8ykUPgFh4K32WfqHdA9+NA57tLEW
nWlI/VduasWO4J4BZR6u5a2E3pD/vUVZ5nPASi2tqxg/X1MzTSCMSqbtRiB73Ioq
BS3B1gpHg4XZo7kKoyTmO9/SeVnu7fgdLNJbZNH/BKT1IhW+Z/TexplKMOwZULu0
2uOAstFZD5MWNAO1G6ZKXmrHDqjgwo2ONYspqZijKJB4AnousRXlyOH523slXR6s
sl61CaoyjffUg89FxDtSiJ+4OcLyeD6MjshqRLFfMBZ5xjlDOd5wF5t1ZN/tWJTu
+yznoB4+Ve6YUn1HasSwEEM0/HLzFW0NVe/CaFCPJDGI2a/RdRwQN36If7iAQAlU
74a98y4i8m9LAmSfZW+kPDsVSYy+LJ1oCvfNcs5ZUvn9S5zmO7HjncNiF+naqtq1
Qau6lMF1lQVxT5PotugjsoyfD5NUK51VASAr79NFDkEGo3GsmTaqh9GwvpBTMh1J
RgoMWLU1uuYSB6atjcbTRxN6+NDiP/VPx7sGww+GvDkdt2Hx7lj1W2TndiLudq22
f5wrsMCc3J/B4UsStJtdycgn3nKoEkOOaaRKB4hgeenO5O2BAKn5zQJ7n4l0RkSD
G/gpznv+C0W+C1V+HGMR51dMpJWEp08j32Z7u5m92Jf+drG5cnPt8mdFbUmUUscN
KX96zaPZpWN4a9uaJuOHhm/IhHFh15DXc4gJOP/Y/Wh/3sy9qR8igToHVnEUJeUf
dijhgh8Bum9XSUMQDxp7l7FM3rodXgVJvI7OJ2OmhXWezi6IAxZ+R/Rdb32HxVgO
rYe1cXWsz4MjOxG1Ti9WVwNCtDM0wBg8gLwUsxYcrKXGePV7J/EIUExOrrDirMhE
alFRsWSZnodL46t6CfyhuM2j9hoSa/SrH0jICOHgarEziCXY9sAp1pq5OlIPC7Pd
SsM1/FWaf17NGrtL8vUPM+Cilik/CMOvrZtw3eiWtNR26nLgRF8Ezg4Q0mt/Ko1q
JxIkQQ0vA7HtWIxRLfPnpuStMgJ40f0HI4mHKeJcwIsZ2pgeIM8r0VDLHW304Db1
HNYtsrUaZgaT6RnF1LGv1adbdafOVCPnFQ/dUPdnrkePMwNUzLXzOawqDDczDCcm
e6wlFFyShjggnTeL8CbOotJfvtDtGRMLXJy7lfftvs8fGfm+lepAKde8CkjHwI9+
OdEIprgw48iVGD+F/unGApv7jB53mRLo4eq46rTXVNShH/RywtzKRe1JIpf1nCAY
3mXxA/khyuSSHPUWxmNuOBbih/ZSA9ROSYiSIOxhjC20TzdzJ86pPQws+Z9xH/Zr
zjrMTLgR2xWWewZxm1ea5MqlQfHmgB/a8Ckd71s2VuHG+6NKyE8k7ZHhFuJrbBME
0FvqtJdSeAX2g8WCWjQg+FYsXER4M/BC+N1zPUnMqOsZ5HQjl4X1aG+DUWxWmW/w
IEAJphI2JuLB8ny6aVGrH7LZLerpdXD7Vu+SqMVCkLopciIqX0KW5FDo9C6VSnTL
3x8YNELLr9O74jnot85Hah2CgJOxOhqa0evv2ZdT/RnRsyTEUrdksVClfobxWfL6
/RTR3mUikx0UjZ+9o1g/KS07BcPY/lkMS4uKoXVx9Q994aHA3yIF6sCh2HYY+xWh
1zzhvL1GVvI9csBcCmSM/pQt/yPjSmxiT+kygghe7jpZOYgyCL7jsxLm6BGR2TF2
M5vTdUMTucEQ26kpjuLM6tb+g9yyHT7lmODA4DDIsb8f4Xi8pLR1sCx9miQdtYAh
EzY+R694/sS+mBRZseAMm5eJiDO68qcWNYN94ATXiJAszqsFbhA4Ah2LI6PsPyGD
EFKA8WQTNw14+0eTlQGwtzMJs2T85RbeIyYfSQ5hL9zuIVm0736gadWHB5UyVm6L
roPtdS3W6H/kHHRmPrjtjDZkJ0qK2mcG2VReCOHwyFjo3ITxQeqUzNDBzAjS7l1U
Esln15My3jS9eG8AMdEEk7rn/Do5HsKCdyEAda185oGHn6lo9AdCiQ2ztW60Aadi
NJX+IGlptR48doBu9HylMcqLdDndQxMXTcbRTuN85YX8UFnz9/Ft9adDqxaA+3Vo
sXhlRDCP70LYM9+RIxTx2Udx9x/hCnGAmSUIRZEP2Dzg1cjvdZ3UC4OOCOFnqGjd
eJKt3kkcIhsyRqfCxC2hAmCf8S+KFs6XX7DEPyScwmcwlunzGF7s5ZVgtVjSL1T0
ivto/efI9viF2CAIpKaxR18fGmSyNi3Kj2UMdkj4rTW4Xw37A+rZxNPk7KStdRCO
/SCNuNQRwPpf2dXTkefSq1J/PlVMSaW6VCQ2JFpxZk+RU5XW+URoYbFi1P+AB3GE
lSLe14KeFkD1PdN7BT5+or5cIOXMDdpMv5tQtleYUkFSvNwgTWXSv7EyMS1ukJ/E
LezWOvugmdHx1WVwWFD6hC3QOQZ4vn0VhL07CYfDvz0O5JwuLcuuty/mNOoBDV5o
zKD+30xQFF21eHdS+iP5LzWMZmEAvYZv9p9yvxLIUwyD6IpqUE7e2NMm/zL7wg1E
EvTrvHSJdRZ//nakj1rSy4KxG1wKrA42XBgND3rnBM5dohiaRaK+Kzf5FKHe9BA4
LzUasoQzliNxEOGzONqmsl7lJ2H5jDKPsaiOSfZYj0fYfQRVv5ZAeUSTT/sc+hh7
XlajQgwbRVDuCpmhj6FHL/6TEOz4XktsPyF6olIc/a+Hp3oltssZKI9Y++p+1EXx
qnkq+CAv5jHatP1GPJuZ4f3eQNq3be90CEoFbcosavALFLFT68Ub9heGAnei6CKE
vlxzYKsX0QdTkVnHdyxRqAqk/0r33UFpblWWKy9RlcpCf3Q/GqW+arvTt+sZmYFt
TBCv5avo+dvaQjS0PGrJ9TQusEE/GPwgwskXIPVg8X0NgsbmVHvMbfoyB4xnLhpF
bOjzP8/Red6UoQ4XaweygqQZSW7TWdCWZmYiwlhFx1fNe2yKIIKlDA6/JQbzOpmF
pbGq94tPDJ+SayJt9dBQc6qZq7iI8xztR35jypk1gG/WNU41UpGONbsDFixsqVSA
JIXHeYOBgw6EQ2ftR/dy2IYJXOhPE/c8kJjI4jI8V5GhSXv4SN4/8QHt+g8Dixub
qn3YDfXjXCLsuMuDMl7Jh666SRGpWZOia3MnypZGT+wufieqjMLbbtSBg1lHmZZy
o98vsRdxCAFhY7E2+pX+rm8mL0I7UOfzo2z+SYyFpE/8rco9VAXCoyCrPJvXBLr2
qMDjkDh2o1Q8v0Ng3b6EJoSRsugkKXgPRXqyCwlFJx3FAHsyXNfgErCnn5lhUAdc
WBrODBgCBQzHN595Pk2g3TuCueabIiqNU+Of83uCXFP3mbS0qCBAgPDfzWjxndN3
eLin5eaKJg+ikP/9+QCSRv37poD8yrgXM+4GQbmayPoxVJ7fUwEOuNnidhbvs0fk
phkST954kP//1VyoXuwgBVmnucGVisFO4d3JAk7Tt+MO9VU9uKFDK+StF1lfUAC0
ljrPrdcMjKZMmW4bP8gw6c3wcQsSdHk0u3iZGGTBcBEFpbRXlrqb66BtLG8bGPAV
qOoNvp4nFZ3/QDF502TmUg8M+5eLJ6PLH0m1zJv3earSGURPZfaYr0BFFQgqQCDQ
HFOSPMIi8VTTvS4b1/tXfS3LrOq03iGF9brQAI9i9nuL3nng8oDkMaomNFoLdXuC
TFcTJaj5QpCCO3YkzvpD0RVcYXN2q3Pr9CWyF3VQKe+qXjfkSVN4Y5UN/Nrxl4P3
QGdpvbE4lKhQ1HnGf94S00ETQckkWa3WxPY0gwwjamcUieSZl4fV+G2Ab/4Q9M95
8Y9GsXmBihcFPaCK7WIWy+YJ+klLd0G8p30sbUA4tZb3VG33RQ3lxhtfjURAav2h
NrTFz9rCwnvxWydABVOur/Ue3d/+F3OZplNAdoDMlfGOHTYOPy5CsDGWJO+gl2p8
z2LCHojiqDsMJps9YhFGN3qhADfZVVDtS9XsbUo2Q0jcPddx63N5g1oAL5UH1nZm
p+4hHwTZQK34zQROT05yHEqhzRqtmyaTepG7QhPpQ+LiVvtY0xwMe9iPf+aEovNp
7O1jaxA7S+vD3zLYhwfpmV1Y5GDlgXPtEX5UgGDPPTQdYs7Qv6/GJXLytB1rlyyj
UG9ChYG5or+c/dh4t2by55KSuPNE0ficCXxgvtUi9/d6WTttmmqZSpHH0JsZpq0o
1eIN4BDFwp2+Uq9aqnNv/zYizMHZ4AVTyETtKq9OFZQ05adLi9x7nCfOrmVq+01g
v05NsMBd4pwehV1mZFFWOc+QfSd0D0P4sqqqvkilgHyjP0q8g5wSYbqMhRDWRsMM
gaVDceEW2J9KdT2vPff5ZIjN6wYCJZ6H9AGkE+9UuDFLW0fxkGl7yMQxGX+kf7nA
HwDo3rtI8lMWtkz0CAMBeuNGiDPwpyJY0gmR9NJWurCLFr9+utRk2F6mwhGgZlcn
rm0yJkAeiXDi5bw1Y1IEoSc3psz4dtiYUiKlK5nrFHSGwIzsSuu0az5t89pPLPP0
DDKIX/xowX0bGglGAJ4VRFtIzsnZU+KAVXBwMqZDt+G+Ual4mMQjQ29w4pB6CNeb
XlPTi87LOPAIRNuj1UACx1KAbFaCRSdMAnmRdQB83MBp/li5mhgR6pCHAT9VfP6c
dgoHXARJgOVH8fulTQhDmeKtkTplyP/ggk0gEVkVUwXtB3lNGyuMaNIHYZaqPWVu
TUA6WJSbhFAKuNKJRS3oLLwkcQcwCITCqIxjWlzW9PvGvcRreiUWKyPSK6FpQU/j
b/HBQSs/3OMwDN1H9WwsyvsJNaODv5q3M2Y4zZ7w0VZqqX1AeA6hVjsPEUG6lt7F
b09lFa9kr1s50Vb2lGlaplQ8MDv7U8rX24TX3Oht1Ewq8NwlRgQLetf8GXXA8YBh
jki8WFtd9N0hTbwh3gWz5ORlGqG5Gnd+eIPMiewYXPB/UFEoXE7uQaaQhBJSKgmg
VxG3Xuj8+j3fyc75C8ENDY+7UQjPZJQHaqtkWUm6jBwwwV7xBMd+b4qNkTCFKePU
hQ19mCspH15DXEuToTR4HWClEslbDRxOl4p8PhXGapHL0EFvhfGP4UUoS6HYpNOD
F/vB1g7/aRmapeALZDj1cLiMnJ1OnBElmVL1IlhsZCVcWuDkm6BWvWKdow427FqZ
4khe/JkxXi//xgR4nK+SEmQC3KYlKJo/4rnlhRBDO3i5w/HfxK55/tLAewXhjLgB
jvn4wULfoK0xedYlJP3lvcGhPkABZmeukvRyHqRC/U+yQ9URX1vcPckVkzQ5U+0X
HCfPFAEVAe9LPbufuxwohh3rj0yDLKw5R0wHfnIDaTMOysOc27bTr+WeEXTTfbJZ
5cK8S+iviz0j8Okt891sdqJQUJt/13561mD7ULeR0BPOayviSOPD2boxnyGJE6zH
uoQrSeBgVJ/DSWBXAIdMomyvHfzYvS8vCON3AQfBqyiP1mDdyFY9Z1xqF3vl8sCF
esEAvR7i7HWEQ0uToFTsv0QXhXFS3rppcP0vEagaYEXuIOGKgly3JlHbi5pIljFV
MyJGrv0+/Bc5C9cNYKrecHDe+xJz2c5EE3W4xZqyGeDtWs4S73fhpCj5qSz+gdoj
aJlRn7QOlRLwhgS6Ea4ojrXbSSnA71xekJ6S8EWBMz2HwyR7RIK/t3f6wufPI53+
BDUMIiMHSK8e1xzB3rGf7i25h/n1ThtK/l1td0L+GLEOD+ekYxQs5pxxRnKmvip9
I/NNubJzsYER7Xfu2iAxjQ9wn39Yx26lrRggElfoPzqICVLc58G+VvnXmegL2/vy
C/LcGdfwe/94VpEXC0XomzhqXtl4AmOTy5NK5T6AbJFaIPzgm9RI+btzf5r+ACd+
CevA/o0zzNulS6j9+GYiwsPoaNqswWA/XGvel0pipGe+/8tbfllakTEzNkN2EwBQ
PfbnMUfysBDGJutWKihEJNEeVL2LFT5nG4k5DQm/YiZJh5AsNIVnlwA2Jy1P56qj
ydGYLHBYD8WLxctKavqQgRjA5vO5f/GzW7198ZxEYdBnLSnITAdjXYAsDr/JmIg7
XN9JlIF7I2j+CoITtfVB1mVsASbOEWoDqaquR39e+IHIpqwMySz+3n1bX3WA08Ja
fm6yqAcQjsyRB2I6hYKGC3A1xpDnFc4RrRO1LDowW+fUbvlTFVORDo3/EAOrJgUb
nAvbaWG56Om8eW/fw7GjjohPL0UJ8SF7W99J7OSDiDS+kg4k8KfO3X/fgt2CzEl/
AkVCzWGZsIY03aMawXoFcSvhdbH2hyxHHQbhsR2V+dgsjlLbN6gad1DbXyOxUVW6
uQ++IdCf7cpH/e0jYPm0QWcbhVlJ4uKU0dAdAf6t7hBRuZNLlHEaZj1cvz29o2D3
R09uhCF0izqIT6hZaW8kCnECfbh5Qk7k29Vg0XXB0FEP6tA/y/NdXY0+GsLyg6YK
oI8AHCNCeiLi3sBE/O7jta2ydBI+kaV41pbUaA9+wabyd3RPjiPpeAgO78WVDEpr
GvkzBg/nxJvDjRQGI4+6iBCMrAAOlmFPvNu92Ny5qpM2++mENz4R5+du1dzk7Iso
ptYK6UqjTmOf8zCGApA1Fc7f3tjmEix2+QFw1hMIXs1Scy8IXB3Y3+LPzM/iYYCw
OTtNfHECHibjf5o+vBo7RA55ExsiRRoC+rQJ477zLxQyvmevrbMvsxVa6WCaFEEK
LV2M71+6b77PoR/E8nj1ZGwsr+eDDBzQaUqsmsYpGxuC3m7+SvXluqGHk40dZZbq
yRrraGrugNMkqZXzR/fZYiKUz/2B3JWpJTbwtMEdsPlps5AgRH0XsUd2JM1SVp3t
AR/1jah/ND9DRO6H6dIcHtg2xyv38wyJ3AnfHkkRyqYPY9bSvU3zBxdUajtP+p0g
t6fDH23+6OCiCJ6Tsb+h2rd4lY0SRDIVIgDh5rC5YlWeWB5vBUOUqd7LQO5XXDOz
/CY1c7fHrXH0vKShHE4Bn8hPQL9KsRskxM/HRU5g0H6MpsMTa2qAEZTDxP7zYoGk
bJT3jWuKooFQ13pGv9cJJ129+H0P7W/c4CMLMSw8TeshXki14rsp11lbqMREN7Ci
eQVJW+y53sfsRuS5p/9JXu1E+MWXX50ZmP+1TvgIC7anGrbtcH71slMJixbOeJ2s
fVu2w+xmAi2lTG2XuwftMtLtc75q9csNNMKVIT0uB4kmRPQHE2PiuRrmnj9GG87y
gH/9XWLZaIKWOmHqvU9XVIgoSKZnjxITsilClr2Bjx1RR/MplUigv7oiwX2yeoFK
lZHTXwAaYV1TKbOlePG4rhhiM4LK5q6o0HgLYc92KJE2+heaqZIHIx4GDiHsqzKH
KsmnADV0b4MoMAlP6kkXeAOa9M5Qgal1ul46BU/m2UaWlygazmq3XeDr/8m/9kcj
84PKkRtjm/9PCRYI2ZEcPYx0YsG5MsWa/fqlJms9o5Yq99RsbR26TIu64vGZaGr3
oxnf9iRspoBW1cPgVVUFS6A5/yRfpWNTa37YyrsUPFnpSs4V+rXSr9xraq6Xwd1Y
Zkjc4BwCwBIli0KqkNsEwNmcZWWqH5Y56lecglWtrXQ+TVS11ONTys4cQuayRc+r
yP1Dca0sZXFgpqBmuWKHPzWb39vTa9I1M2HMH4cI0K3dWarTNanUUxnMdKypQafb
gp/qJa6L1+CxSmYu/sj1jc7zRTOUJPje6DyNuSXTxhGBpJN2BLBe25ux84hb7UGL
rfx9DGgbN2jsZzPrYDbRcVlL5lgfFHUFAKDnYQrQYA+dAff3bxZtjgPmrfpI19ek
YdFpPp2QQvFpkhxl7LoMmmhZ7W7J+2VOOYUW3SQZ6BRw1FKcDLE/YprEAtbzLwHS
QKe48XRHRE/irCxgMXoC4p+XR2zua2bNBE07pNQP9/BX5gAnPFfxNhkhTG5eg6Av
F3Tg+pNJcARz/KOvfaC9Xo1fUJiyjKl7P7Y/Owrc6qitQ2SGI1uSA59frtvDPQ9j
/njis12TcgduxSRnx3S3DPjpfNLi+AobJA7yKh/x0ZvZa8UWNXi832UjmaNhdQCD
Uzc4isiB5yeEzi4su0AVTxtBySr60lrdr3VS4RLcEFjvK/A4F7+VD0nWaGV/eu/O
98/cng7JtsAnp/DgZIBa48cPrVlRL+TgIxEs05q56MohMuHrGmbBNe8Jykhowq80
zbXJVA3mzQ+93eRNIXkkESWXTw5ewyEt8p+MkxW0O2ShStagIHPaG7Vs0uqalZKs
wI6BH9JAWzUn5UojjtKwu1aDsHv2P2sv49+Dw5dCdOFImHcmwoZpRg1MSrSg16Ec
hHv9HoHBebRfbxw+/38FztFfyqKvovVa5UgJjN7xCdzHUEvJBScbaWe858ZSPTq1
5hro3rQ5FLbZHCo1DGfKXWkOVeOxNS/MYOYHLfVuHQpaUlN8GBNWCElXJcaiU/dy
dlYFz14hZh4/guyXrizr5R57/Tl0Ws4x3YWuvmY18WwkjmP/se+HQTcuFgKmfLek
0ggbxYIVEDxi/1/msduyeFoqJPpWxSzWhezj0lqE/nOJ4TR9TXh2rVUJ4QXqTJ5g
IF+lgJI19FSXjuPIMZF6MlWEPs8uo8KktDe6h3MbcjbpjZe8fTiUs6NlCRjIFYLm
oCKRgdMwLlYkAgsirjaGKEDslE7Bu3zWxfibiyCiTwVHDtA06aYs+CcsWqrqHChd
WBe62Blonis7kzgSclPHSqkfvIUKq02vxTZHURayEF0NpUM7j7zV6J8hPEekK095
GsVVll+2hH7UuZ7NFMl93nE4WsnLeqHwpJF0efvkID3OCTpVmaGx2f7MXjzkeb8h
ekIgrJD6JEPGo3fEoW18NdkW3kBvjTjH9uFzHVr6zJn5ulTUWYaxoJwrjPBjyDGx
lhRQifcoeA+34TIX4til0nGwqKwiAxPdH58c/P497gXPayPxQaRVrwUmYspCL5Rs
29/GgOMOrR36vax30qFly8cpgXIYS/F6Qkon1NnJjhJLQDnunFkzH7btN3TAFpTH
tIl0aW1OAVqPTWKL36SotdCAp74Nmjt9tnNPfaLvcLn0cLC+4e2mkbkyaCkDjVQK
I/sfHwsIDKunHWGnzw5ddVhxsGTwXfsJOOa7Xp3oZx2H4xLW49QK1R3Pcw/W06Wx
gw8XKrWLRMBN4+VD20YQ4roYOF3VsfxTqaRpiN1cuNEA45JIORTnmETX0XJYP2mT
lBdMHyj4uH/wU6Y34+9IxYMyUI4kDeunqtPg0cs46MgfG1lNZc9fSdBmXYCiGN9Y
WikTCvCbCBjqzMusvNFIe38KSBnrUveRwmKOgLU2na3eDFt11Ow+jiZwo5f9NajD
ihh+fhQdt6Q4PKoYZY5G5LyzNPi5LBBh/yJOoq2Urt4AR80VXx5wjOYxXtj7LNz7
AoP8v1J0WT5fJqfvVPcr7DhMPupJOmWJjNNc3kZ28mVFKQw5EJ8Ler7pmLIYJMh3
ZGjXcg8gPI3x9ObqtPjmkgJf7cFjxvFk1oVD4KyvditTeNh6LxAGE8ALxu5J79Ah
/zlbuZzmb9PywRHlPn+nzYl7LxrTu6DAes3RIgnxg0pdcqOAscSXYO4r1MfK1znC
F6Xg7AhHRNRxQDaT5AKuIJa2tzk1Txibrko5WspcTxBgkJg91W1h6WjjAzIDEtuz
yVIpHiDekp40pyCrL/kEwkVZ9c0vPfFVuIox+yXWxgTLintuTsrmgGPeJSNFf0D8
cDqTfQ99fJXAyeIi/Wy85d8haNXA8elDSiVinMZKEo8Lg9WgnPCA928EtOIvVhsJ
zAWJYGML3fnzE7UbD5Jl/6eUpjwPH/9Oh44ZPvy78tIlKWQBW9cZU22y9BThVgUK
fDsY60ysMzNyg2jHvtGn4/kI02L2ikofFC72F2/mb8qydY6XNIc0jNt4ni8Q7+iV
e5We93tNimbEvSqB+XeBaN2S7XQV0PplwEvPPUV3fWVwPqBPUewzZdRjI/ugoYwR
uIhT8mezwLeq2IkgeZM7pKEkHSG61AfkvMHpjooHp5ZKiY+UzWZ8fHTy1i7dwScz
FkZNIu+MWhwD8ehzYxQmnozPerNiyuYHFjDP8Y1u+murcCONbWLFdbRT86b/UpaS
YtQl5Y/4okKLWogY0ESsm9ITyFq2L4kthmST1VV6g6MyvXZoWErSMPP5YqlmIrhz
2+Td2suL4b3oTJ2ChWWkUUzCR8XsnYVsoY4ISGLeTKtBzqMpWgMusvYAaq8Wo+E7
L2e0ZX+5DW9xKWfU/5H23OYht7ZlTuM8TRgnSw4vnaS9ozp/G4wKhPEQmfWMiObF
+lFnwB92dmxcWlQBwWbIsVTU3LGHzPO9llYnxXPLP2KNu3n0oFXf/rp7o1zxdbDc
3fy+zPbwLSEj0VoZjRFCIUgqUVjraFI0n9o9Pd2GcoPAkpr5RCbDa9LXAfNo+vqk
bv3bOdT6Ts2zmD0ucRIxMOe+BuuAhjjiL0QicbBvxMtKfeblTU1LKkIl5dUTPZjq
gcfeqLvhiRWB2CvZFgkByAjAWEglRzReNH3uT5Ghal/dZOTsoUZT5a2fX1v7xgRH
dpr5bjubBg7DiBIlBsvImxTaxywWQva9aJFI0hwiJsZHK1QLR9i0v+o+HQoxRV/y
2icJCRBlK/HgLFvRObkb6sfDgfqIPhx2sWVnKJRX559xN14CMeLrHWuiTid+lQLl
TsgWV+sAPiNlJisuqz/nOTMkJzT2eoOO15n16oxPInbEDhPfOu9pE8sTNyjvMNsN
2oVbl8PzvguPYIVAyv2WZuMT1mRn6nF9PVqeQiL4JCkwt/eXSyvcsYn+R4sXtP4r
Ue2VAo/imI1b4s1iJOLAl2482pmsH6Lxd6FQg7BL46yAXyRUBp638GogxfClqiSZ
+1q1VHXxoXqK6/eXtkmILuP2E5GzEW42D8R6JBOHkFQcTVM54jiHmNNusyWsLss3
prLddxJVTqrGFzwu+UZneRgRMKoim2iBA7RWRkTF3DY97jL4WNWU9f7fYs+pUBHR
mmrrAmZ5diu/KyzKeuACJ+yLHS+M+6br9Tyngwz0jgddFCQQwjv7EIl50IF56zmA
O3TDR6fjx9MMhaV1R8Gfi7Mal8xiYQBdj08qAnzuA+w4qk8BuK2OPYQt8WYJIho9
iOkZkjfZF2omMkXMDw+z+H3wu5boTmMgaG30DyXelDU4BiHjC0xTccFwqKaJLyRh
J9g9bbgExxkpZz+8+kuqQXaHdnj/332dbXKtJnQ/keMyv7XhYA/BScBk8RWty+Gw
rZCScvZW+mo6FV5VSgixl5tnBI1tVOKRQ8nfpJbIdfr6cSwO+SrtvlSekm1ceo2A
0GhDE5QKsPxejeTNZWhPmF4plj7zogBsC0oAdAXNlzftHq+T6E/OC50Vo+O31gk+
t9Mk0DGTxJCfxNkIJ6jX878DAKwCKflYqPcpyyh2v1LmBOq53qcEPIoRx8pBHH7W
1BD+TC196GXgjCMqPFZCMz6u792HdrPBPOoY4Tsr/ZngKQDvKtSUPWkLLzv4YgNw
aChSgyQPEzQJ63bqsCs3zBfNqCt20RhjC+hOM3TcSD/yMuOj7ryKfyfym06/8UKO
eLPWcRJ04f77i12TlUx9chrok0XdMJP9YaDy8wLjWSzJtgmA3yW8mOuM/3As3X6q
sxJtxcxi9BHKs7AfrSS2KgTzy+M5gCseUlSE1VkCxEon/tmbB3mq0ROMAG+UVXOh
D2N2Vz8uudrPy+mZwCOTQMqj6YMGtcR2E8j+tvoHJK6s4DK2xFNHFmzUSi+CX5X5
fS48ZaxDy3Aey51CXx/vcu22h27AnYohwtdHKj2+D4UN5iMv6Sij8mT93OBitgl1
qRHDz2D9b3OrYmDJyJufVUpHZ7GEplnXnS6awr7Z6EByLX9mxOM92ttixPSS0e0g
ZFQXSJhCCky/BR8PUAue28UumR6kMm7GtZOd8i4VgFa1zeu5VBHLYHwJv9gMLTRp
hHM3BscjJm7YGgjxNuTTlsZCVK9Ph4aQZkeX5z6aeOA3BiDsI9QUmloPkkEk5eVN
sAccNIRgPv9/FCkDwBAgUiQ+WaitVi+K/ZEZ48UM8XWeAm7bXk+KX8cCNKgmic5N
i3sM2NCaYQQGoQ0dPrwnUhuKKMh6TrH8QZSAzVemboX3BshDDB1G9tMWnLsjze+I
lPhzP8IVlsmX4JHFd5GSfyuBhRgn4AJkBhxUjP7ZVGr64+GyLETMZP6GST2mAgyf
TU/z2LdEf4AblUhgfmVLOJqiFAR88oiEsq1+bBTzc5mLzJqR0yivsJJAUJNjPPSl
ky7wpeVnWlP2y7alapCgeLuO3WPNZbo+PfHr7EJcqw6mcCbdWqworwh09LHlzKWy
Y8yPiUnIxIuU4dPNFs0FZRDOcFb8ZxLXC7Uxs/hwfKNiuKZRA+lj5dmCEl+IXYv6
+DghWXzHGMHhvaFdfaihQhOozPTCx5bdbR+uHcydFhO2OgHHRC0ERwPe/SGwzNvh
doSLRlKFHvd5oEmVoLsn54wKsYIjxVoadHRPEPprKyhuwNhBQLLhiwa7fsXrw5MT
oJJb8Gbd+rqGPKihGIH+H8jFaDAn63NRxuVkCn9GYT5JbXPjyfFpiiN1zPSE5eTO
TAIg6IFADKI/ybWL5+n/QuYTD7nxOfkd5Rak+yCv7UlbOJWU4sY5MlShbnVL7rHi
Dr/8jcoiJL8g+UtVob+u4RYK9GeMuZFEk526qvmuF+YeGGt0BzYSUlz99drAhuJU
bvpLHFQotLJqUD6kkn7ee4GDfGYhI/Ji30UVcudbXWz5Iv3EcWQStaEOj9/iweKL
0axWiBx2u2B5B5ek0qhi/5sPP5+saELd2F0kMnGTEIfwOkoqpnPMM5OJojhs7NYl
RD5pK3Jze01fN632Z4bV3Fpf8ONfsGVatsRSxWCfun2m6lEExK01X1kxjJkZTXb5
KxJyb0mzyBHPGNudCni5Wj+hXGXbf3UpwRmuVlPIiMWMYb2D5y2K+0RoEZjsaGxF
rn6bxrnLEwV/a0j5WP5m+kMQ/uXwUFj3sT9Uh6ej548uPc4JPhXs3CiX9t7Y1mvz
bFdRNxcSFx4sC6BTvmxwZSS04aeoPv0xWWMLjCJsEUWNlUxVLstBiq3QR8vDSoEx
W2DSQAOtpWXUPp/Bw50cgiNibmhF6HoLGFIQtaVtKJlcM3eQoPSKJPpmkhNLT/WJ
l+9aJIqhtGBOU6uKqEVHhN24GVcGZBOC37uqHoqTfGO/hA5IDjvI/L4jT35wozGU
pZO/kocogzggBnFcUac6KvSfE1dcnyBt7anf9XK0JgmGTtHKL8ZlfmU5RoGFiBgc
CU22Btt2+eQs0iB0ALTNgPNeFpMtcrL1VSwZf3pek/EPbuPHRfZ5mR4cCAZJo2Vi
Yifox07YpTgf96U2zF9rs+OJnKe3sT2dsQa5084mhrej1p99ye8zXNbe6MzC7wFi
A0Hnnw6DsUKwm0RN3gf+XAemP57FC62Ojv4FaEm9taTapyBH/zUrF9hNWUnfvIxl
zpNKz8QwW2bYasdRW8sObuUvJIkCbtVbimePV1pvVFDY4KFZJ0FnoEmts9kFo4yX
nmWvOpLHzNNj6PeY2yhppo8ipeS7YNliabdMOaffw8gs7Jq0jutzxRm9u3km+EyN
4gM2K9jh0ZcPZkmTWv+dDtjtQWj/XXX7hAfhbcfNjBlKPsMakJX31DsjgrZOPCda
9+TL7Ji0AeudywhO0AU2lFqKG5JyUzQJQ2S5yU1WQE6xd7Td/JSeyYzBNoxtQ9je
KsENGj31DPdfXLfu11/jYfE0xwCJBdOU1EhbVlYnw4Fs+1PGUIrGq72pgZajDQmp
H71I2xEQJseCQPRwX4/KxpzIAyPWy3Cml7ruhCNstx0zadFFhdEhoo6jT1I10jYB
BVk+1CyT5AoqhenojIWXHeMSUc0Q6040iyW/GaQcIKenWvLpIKnr+H65CZczGlU3
2qu2WlcXSOBgTgTfkEacX/pTM/cvQeM9rSNUV1brzfDLBZ5toYCHmxsajDJNfxBj
TgMgSH+jrQzkd6GAC5kw8NCZdIhDKBGdwhBrjg2FdfyKuvRTCkBt2+TQXBNXdpib
J1cecaC/2LfVAkzUxq88uvWwTRv2/PMvfTUzZlSaOEb82RYEoymk2GOvv3TrQJAx
Gx/Q/WJKesJ7Vt69YIJJ3cNisbE0uSjfd6DDO3OC560w/pEkbmNSYRhSyHPD7/TK
yZaWlBy8laeVfcCIORLqMAd42EqrFhfkAqeqvIjkjI71qJRhslHkTzh3oKGn8RlA
gyIV4OMZ8v1NQAjBcyzdxWa+cY5ndfcF2bggPgN8xeSoAESQIuxiEz3dllJz0qnB
n4GP1h74AIlO60Z2ucPcmwjocqyEiZSgr9m2p3+7Vl/D/KWL4CqYBpd3zsNh7qSF
ME7o2r+Or7BVFkxJ3GMkXJqJl0M423lCDI1BL+oBUc/l+I9KcyuXsrB1c5lKF3Jo
pawSwquQlOd08pnq8M8gOX9u+JwJDa766naOEmGQkHBeetiFOuHxSk67ihkqx48m
2Cm6K6huQgOYTeAn+YvC1VPT+BaxHyJdWMYlJ6JhK8ZgIkQ/YfObYfZmgaEe9YHB
jsVsfxuORfiZnmPcyKJlO9PYWvRoqAuZLAHVi5VGk9iUgmmR8ZfkCmAgI7VgjBxF
X2uURRtt19afxPrAzTkj+egRZtFk6MgxvhsbGMGaS5/sLtXQXk1hMEnaPoRH2MO9
5bfn+oAXpVis4p+HFyKGUx/HAgTc77cfDCL19twRuzhq1V+mGrp1fbBMlNDycyvf
+OoRYmKZwnajhFu16qbSV0s3UZwaTnNSiGUYidnX+HabVMjRfVC/svL4DkhLPm+u
NkNweMgxLun2uuztuN1c01Pt7eAE0OAgnfbi7g8Kh/2gPsdAh07Ud5hLIodH6MeU
R3npt0rOqhCPliI07EBOmtKELPbI65OuewmDDjRt9CBJSVi/sNh/dMA7SJ08kuPL
28S8+j1Qrd+oNuOeiyuOwXzisyNLoOELiJmir3/3zKqzkNSXzb4pH51HfoiO/fjL
vqUXgs5g4nZTaYHblg4BeCwUWWsx0d9C4LRCfEJdY6fCsk2SOm09oKBvOSqu6w02
hc0PfgfdWt3Ml5OnM2GC7JFctCPgRuKrzTqe+CYrpx3BhDwCnn27XoiJJ63RJslp
ULq+QF/68zyv/eddOblRIg6ekCka4Qng2lWsocr1NB4nK3vLl73h9Zwa4aKU06di
+3r/lVt4MEWY+pmhuSihLraHBByCTWH/kFKFwoPMtl2WE8PxbNeBd28LbY766to9
iEPAJkA91ck1HDVX4nb+t/TnZLJGewVKYqmlun6Xebd7MGkY/nvQwOWP7Xsb3FTR
ziozQtlaU9TNCcOd5yT/xwpMHx38cERkD93xNHT8719PomOiAiYUHY9Uau57Q4N4
9Hf50Pc5LgwotupjBtnYK0XL+FYNXWzMPXZRJEvYTdJb1XP7Rrnrsg7UMyp7QyuI
3u8L3Nb9NX4XvpEbelhChcLxpLc5xm5pcmPDw+vcdrMEpzh2FKaio61tBTD5ZdAv
9upYfu1FFC3jprP3jCiQ1qPrbfPaXomqpYjGmK2D29jJaCi851BSzg93ov0Td6Yd
eGTi18pMH3dDYTpKldWd+kB9FDC+22aJVzjEHRKZximwO+bqWWwVQM8ICb9dAYhZ
AaGMKuT6uRWTAbEINCBUj9hts/3dK3H4lZkLTYZEVoBWTOVc+wQHgQfuZt0Kntco
VtTog/Aq1K4Ojs7ik/jhBvW8gCYi93zm5gSg/GieKcbg/XOXkd/nTaQvGG0PS/rj
JTBATAUbo3Ao5iNoboY9iAKXHE/m3rQSOyFbgXngXsKo8kh6vZXkcOWztv/rFzpO
8P/M+wV7NzFOG0QUyWPvTh8iXvsQUaZRmfd+pTkTovDohO9KumeUYHh80RSTwH9D
XUAYj8Zbi9CMEi3L/d+HYf5xNFnR1jU3W+qTgnbu//QeDShQHwzdm0taAjpu49w/
guuFI5b7D1v3eis4NYMCi7ZXIX8QjR0Ka/wE/120JCHyWnj1nTSEtVgXRTbeIxNs
VmA5HS4A6jfbeoiSGmLQXwXCflDFI72GTz/NI/w/i7gxy7uqlQMxh+Sx7rkhb6ND
8C0ziK8Yw6Ol+ca2+AtGJ+97gSjEMTy2bmvDACBXu8nl6Hpb3lAkzwgTq5Pn54As
vJseXF2+Q50Ro52Li7kgbQxm+7uakckeZkHpO0nnes3o4uZMkR/ztgpNtum1Mc2+
UrPBMrq6ojVTg+a5nx34C8aWc/PvVbQ++WF5tYRes7NRGklUil4+iGU4U4xTB6ai
wYWEEj8fwg8GaiYy9Gt6Txt4bm7g1jkNEc6U0dPQeNJpql41rww7XB3A0e0JFNbK
VXmwuWLkw3Lk3MIUR8zI2v01v/SzsoHY/jbx8kHRFvb3BErfcVizqExhNvnkW9nc
9/Q9e7o0YOqTU1c39PopXxoF5B6ZqwUIdUR/+UxRTfaVSKzZv+KGIN43g/0jMXCq
CYIw0rWjmojPFTSdEcTek9XGKuR1TaXl6aig1DMGFt+1yMmqY7SjBb8CiztCZh8T
b6NtEN5uxl2b695aLu2LNyLL2JE5CR+m3C7Aii8+6kupbcU3I0FTqqLZ9zMu6fwc
W/eiewtOF8Pms0oVKW8OZ2KQDnCklXRh2cd/z3lV6BhKeHei/hqCbynw5GfLu1CR
IOE2G3T4Bm2epWh6CFimY3sT5qKjMXiQxCpLCWJzy8Sso/z4KLZYXc9L3SBjMxVI
2fnqUUfiybIRAzMAJ2DYkR/Sk+4/5GJxcfSvOyqDPXAijG92PIMsvQKqpkYSbPHD
oL1xc3kGvX496oe+Gb9+chnZJeL7z0FdkzY4MXgIdDHI/0jbFHgbjh/M9lDaZJ+k
u3565KC869UDA+N/rxMoNULm6Psi+0wYWom3BM1wCadI8535JenqIXD7OB09Hzx9
TRRrA4Momtjh6PiOF2VOZEj+0c9k+QghpdBbKHNkqLZvKEICdqXBHALc7jXHA9ls
aIIZB+LOpiSERI9MS7yipNXjnaiirvMr+7X9QojANrkHPeTMfaHundyZNRr6Fu0X
GaB18zTwbWn+Inr5ixKvp1PwkR3jUGWZVhn61p7ZdYdu1EMjvAVSG4hJwEeHdyRY
qqINH/ybizxMwwx3DG+gJ9yYBFwoEK45oGxzWFQ8KAIEa0Bx5V5jUuyvUuFBbpaS
vk95NYPpWTCyd8PfSGlOJGQwlrP0eu/6HNW9xyE9C/EUaJmKyr0xN4Fl/MIaPTak
a+mLeAOKFtM/22Abacjc8dimw8/16g9drplNuvG3ky20YqfIzN844XuuyMEwtGFn
sSObZxln8VLQy6xg2PYgxiglgQmIM+qusF5G6ni8CmIrOEIuVJ2tTRgK23EtnPi0
NE25uVzYdifzGRJjwkkIL+TemqlP9w19rq9S6kHpQqAXSXRLpeFxuUIBkwz9tOto
AAZCtKjlXEc8sc+wIYl41TEyG6TN6sQAsVPHMoxz5EIoVx4xlhOvGwwQMymVamcN
rk4AH1BPFkWkxKHCYVGYp2HaTbs5qaew7NbkF+yJ0pPl2pS21yZNUZ8pnBzee2TX
7BTJ/hPX5znCuXQB1xYyfKTn/Vq281vqnTLK0J2DHNwkpBC1swI7cbeWdnvLnpLP
whzthN+HMo+WPQ+Y6/U0FpmX/BtwLXltAUfSF+WOv9UfqvX7jNoUIPejQqcRutN6
0GgmYLFrBqD1iW3cagM+A5vh8HUYFyfQO/bZjo9sOMI3M/XlXlavUIra2Gt/YRvc
zn9ATRj7QLJ4vrZhrq37zwULoXS+CjjRAf7tUQ/vyIlmz1irwouXI7z3UC+WmxQd
Acgf6kuUCRbJOChuNHK0jFYlGuIzEIsX2u4nY3lvA3aJyE5nKv36gX2INiIJ6Kk+
SMONT9k+leGAcG7MgEZZxm+SMwom+d4agQmsKosK78/YsjKmGgz6bOhSrDuOqUei
dLEXh/t5+UAP7/WCnFYb8ZctQ51WP2TdeuHH8FZQauflrzmCs9Ss8rQQ6Ndmjx+Q
5FqUCKt8q8vYV4KknrWTUV5iHFN1n2tCY9V0jkquq4PRxrS2K4i8TpT1HjOKXG3/
4wUP0H37tyhWcX4QY5oGo+fprp+klSR0xfQz82H/p8aUS7hbfgLCgsT+TDtgiLuR
MyBezRa9VsrLhsDgVS1m+JqTv0HINZ5aehTNGDb5xN4VhuCdj4KORICLfjUpeViq
I1hbX6cryPA/9uLC9F4bpIgx3OKSBtPdpmuufKVBLgyqz4j4dDmQEdli5+N7wli7
wCYPk0vNy3EQbfGdCCw3f8R6ZXmMMpdXFvGy7erDa8gRcfG220Zye+u6H2PW5O6S
kKxcCqXdBwVvLxV1WCXu0HImbjEM//1CZV3+LyjCV5ZuRZXZprtO4Dm2r1cOdO/6
Jj6qHg6QVNxke4TwqKuhtsLZbcioJc3LRsxXN2N094psh4xMrLBBN/aiLFnfPSW+
Lk9p36i1VtPm5/c0TRcP+5LRHkUBcZHKPoqjbKAHRH4gtmbRgXTxDsCGg0iKtsi+
3V0YZo6vE3RuqfxY+tTEbKxqNs92WY19u8+LiDttUkd4200IIV3BHzA8rPAmEg/o
MOVifxyslhnV7LO7lpwPzCDG+GY0XIaDENWEb63lCK5jafooAPw+Rl8ae7JfKSxx
6rMvdO6vwPCfCSB/WGtwaVj20SREbfXHfAcW+ra6CVN1QrjSgaGfi4ZMpHUQG/jt
q1Z7px5hb1mbzb76hFI/3r7mHvBCvjY3QEO5oSnC97mwR3aX26Lz0Ea2KavrtN3i
5/elkparNcuvqL4RnyhkFfRenKWSPNtThxcpe9oCDpRVxHNq6W56wxstbkbfWmWi
wb4y9g11uYjqLL7C51//+w+U291I3btkNEcqdrgS/ZZTxXmxZkvM4d0NLiUqGKc7
EU7HSa9CM9IRYmWDUdVI1lTZmQkWytr4NyjOWyoCALVac4bt8MTUW3xG8bUoMMvr
qWT30KVTggzfR7R8q0dNKL00EWOrE09b/UKrdIb8kXd+QKYigb9ojz+OhGyh4Ujw
QPBdynCvFgcMDKavNiAWBygqyw9K8AZS6xAjlmCO2yvqbhE0H0BW/dLsM7qkWbru
9vl1mQUv3ozk0FlhkFVGImGW7WlLJGx4hFua1db3nh4p0uERB85A41bZltYPB8RC
E9/U7Jm6uRSi/L/nEVNgnRJ/gS8pp9UmFnnTW03moeNfSGbKuTv6/3FaU8eqCVDm
HE4JwYOdqOrszs19auKh8+tAvLcZxPpe/zHmizfnrbPt2MNsyQ65PG9ZO6HBAEa7
vtdKSjBbpsHpl59/gDjfLWbNrwO/WhiyqE6Aj/XqxHzOrOwphbr3DpeMfDuStVpD
ETS5+g6vjQdGD+et6sWLnmi03HBu5HcElZ3DeAPez1GCSgTYWxmlRBdBDtIcAiPl
ZwAF3eprINu8LU5NaX/XK67AVsNOkXAgdat/UrLumT+mTW1ggoQJBrbHuJ+fkxRD
t5aux5aeAHhLFbdY70CiVQDEcudmSo9dkzY3ImpEj/Z9t4hrfYxoalOc9K+nTVOt
mYO0PGY0ioMNHkh/le6IZVPg/2eMD2+uDluYTcYSVTV/STNG7rKidKeq4TN8vJKQ
hfjBUyAWUcNVRWGeYaYWKavqQxSRLSD2sa04hrARtsfAT0StSIRyyQSEXbZ3AiQM
hdcFC4UOdvMj0P4UvWJmREVeZS1zeHzK/GPFyDsjBdz3rLOTFycwdEFVKYs5OGTm
gGaJOkE/sqKfnnTT7AMydi6YWU2IB04sXk/9iDg/Yfab+/qQsP65DdZ2sBHLnlUq
kH+lk0syffJa37AFsFTWlYJmylE/UxXM8VdXSou8DOukqTRDZn/g46k7b66AfWLY
wPEx1uW6zR6ZTVNWjln44kMR0nSk8i7DwZIChguzyumBNg3oWvulbYaY5KPB6A3z
B2kyvtjQaN2l7sY4lO/oH0VexJy/8Z030rUHZMVk6p2/t25S/FEGcH7juQ7RLpmH
Idi7G5hNX/yMeOg84QnWUV/FaYbcbfQGJf6fQZNzeEEdKefkyvAR/8NH4ACzJUA3
kxAfxWPWhSKvBYBctnxiBSSzfGyQ+HyGuRwM6PTYtVD6W/hj9QxuGYh2GPc4VMQg
LeLxfadnmPACC+5Il6RnzImfy17PJ9EMr8B7X9KefrmPE7gZxA+moWi/XkVdDf1Q
I/+DGGAGjQFebpSV16kkwqXkn86HITuQdfloRkbgCKa4/eroqizUVIl/QUkdFS6d
En6F/eVYUTsrbv8qdgItAiZvPJEnMqOQCA42+k06HKWv4Tj5oN8uzhd//NETwr1h
pG60RVs9/qEfN+SSLTOBiUdh70XauZnNVh90tY46JQ0cUNJt+gHqA77EQsZ2cMBH
7Xk4iASrw6OwHYZ0fgGFXoD4qSGXVpRzLqZ6qwEzCXbe/Po97HrjGg307n05c20r
fIIwHasnqHR6BF2WQRbcIpti5XOETTcvAknuksRKROVBXx84lIhpvaDfuwjcR0KJ
Vd6hoGIHPej/FT94KfxIrYL5qaktfbLlUJU5AF0QIEAewOEi/oVWyJ4BfVfqkvfn
LJ+fT6wNuf/HjKANQi5Kwc73hOqL1z+i3qntRtIzP/KSy6HexPPDtYhyAQhdpRfo
EaAg/K4dVYiaEvGk2lE4Ude7ZozTZLkG8dsqo5p/CFYBUYAjxFqVGGH71BUSOl2N
Q3/K6/SMDB0iq3qyoDFRM5HnVUt9v6JyFAdwyfkKRwiQFfaQk9g6mv+P7StDtriB
5Uq1TYhsuTY/Z3mTgjS5p2NTAuWb0qelntWnvIxBsZ2nMIEAiNLbjub5MTF5pLBv
7R5nNWdcDTe8xEkBa86/nFEI6xol046LMvnHmK28zo40Pk/RZqCz8V4lsB3FRrl9
flOCOaTRnsg4+ZgGHguNgGWsNlz+z/jy4iGd6mJW8SjQmtm5uR8OJntEv/Rxgr4V
qPEwViRVr7yyaEwibz5qlUCkuuj0RgIxbBOcbzNwjX1zk+VbVbWi78wPwlA3Y4IY
kiJ8SWTVaWF38YsgG7n9fHgJZ6CPsfaMc9T0d0WTIhkgwDKrBB/cW7+/uQ9hjMN/
F1Opa51iiS/Ly+H2kssoZYgo8p5HjsQJRcQ6jGQOA1CWBmbI2bMlfEIWRiG3Ehjr
T4ixFKZBZ9uQJrkUL4PAQCzkrMJ6Gq0oQZWofD0NYOUBaPLa7uuD+GxpIuH/sp3s
gA44ccEThI+jag1BSH0tPqx77y7FPS2z6Pziwqom9Yjh5SJyExxCAD4BPozzth7Y
q6puWDIkRY05maEiQ4+CggsIFBGAwE4Nomx3xJdQxNEjZh3U37njPs0E0O55ctbF
dyqCnWNVIA1OfGHkI6U5xKWoOwX2knqc2pIX/J2pzUFAXrccRMW8Zc4ccwBJnRI+
Ojpa7aFHm8RpbhWFteXUJsisnvzKCVIk1c1uOPKDks16SEADP3sOlnX4mWgLMwAf
jIgTKnzDYV3HMlyo0k9msXqYCQnF1ReLhzpMvfJunot0fSpaQzV5nGDM7tSQMoVA
VXM4k6LG6iFbKn4fTcy5+UArg7I3US2CuGU8U+45UkTd6u5s4v2XSL0MlWOEEz/J
V7yHBwB1IRjFhStZQRsQqwkGQD5TalhUBL5CQz3SVcNBvEbsV53+gGlxdIxtPUBx
Z02m5b0RTukltUHOgwd3HIzfW8t6ZmKDuONBLEH4hM3mU/nYM0SlQSoyorwqND+v
4OkW7j0IWwh4+jsFlkpMsI4Ly4PyhYBGvO/HA3t8e/CjZzelgVEUu8Yr3ULYuqfw
xjWHzKJVV/7DmDbpf5/HcEi9pSsmVKZyLa4aqg2rFAcE6R/NkQbSA4nwvZyPaU58
TV9eLX38+3XTnwNFJ5m6eAmeDr8I2s3r+JOSN0zBjsyJ6oE4OIrXjSN9IvfMbSNI
BPmsKPlwsRASRUxYlXDJj6fAWbbT7DE/QM7Bqvk0YNsw0idB+6sYo+CooxMgcOyr
SlHp6ixlRB2dB9OQZZdWcA+KkpfBjIeGJQm9kHgViXrJTZyEUsitu+ITYIYJWPIT
fmm3WvOIQQ7yOVtUqBo0+yhG+fhP2rqGxma/c4owQnSOPYpVnEdCqENElgmJLFJL
a1uvvs9taYKhPgYxdDj+1C29FzaY65UsobzS5+Y6UOQGUd3GbTFm/iYmhyRt/eqn
QHmCwj+tk6mG5Tl1OVd+6XzB3vF1aS5g7S3VejCuXsBNN2KXg6XuNTQsCyK/6B0n
NMEbzNavkZTi4z03ZZlMRlpU6W6MzRDD442hJoNgcS+gpc4JFx/W2lBIH4Y2G5Sn
tDv8dkxDe5wXiwZnnkRa3NxeDtp1yjWOvaM+ChCXp76PHaXb/M9fZ0R8b0h6XvAC
vBnechFwF8/k/Dw50jp/MwDmLNA8mVnbEUHcaIzBLzvtohrJUWRcZG3XOogpS6F5
JcW2Qkf8OIl8hDcxo5kybsb7yTNFvco1UZp7wTb+HArG+4rBc53uYr+ZOUXSFL6J
ejqALTRkuh0DyYw72fu5/hICz/3GoTZrdQHS/uBRX/ga6s6hWns3lXoU9BU8bBB5
J5iHOLBH7ucGm2LhkWO4ElPNzs+QN8KZcNVqOhnSbO0LAxhGRJhAuRx7/wNgUuNX
dY0DM7tf+Qd6XyzAelTWjdTkEZlatSpjSQ+OZwXdEhBlM7rEC1qpicXVfhezhTyf
rF0/BBiXay/q1P1/xDHquO3VQaqPOTpkk4ZuTitbgcU5ZRSaxBFU19s5HXLMdsgJ
E2zAlb4gF6G/X6zDetz6WbBPw2dMQ/MioMknL/jt5tGBE36fPIOwCA2+F6+RjaRA
bd3ghkOtRmJyJWR4eGMnv7xML9/z/5XN3hHiTTAwDrpNczTUDWvxIKicvijJlzcz
j40rJuo0xW51I92cGFtS8RQwamr+eexdxGqoHxgxus/oaHTaJ8gERCbOGhPM+wst
fN1aXvhYorgfPrW7HguSuX3NNkaXHUug+/5R51cEXHaAhGEqLOZRm/osP/iVINy/
Gv2WL8qFXMEin2D/4Q2yZBtLq8euulBP03SQQ7Ra9aDVTErbd6wTPwhdkqux9Nh1
gnz0cEUB5Fqkp977KJut042rG2VuiDRz3t1tYX7HUBbmUS8yXvR4edv/EVjAc1uH
sMnCZCiUd0bwS4AadiPKQv19u+9RiXUnZRXpaOFHFvqDjz1JBIonH3HTjLYx22/x
E4J6zupbk9YhhksrHY8Zz6fw7fJRiGqLhZfJBNK7D7/Le5Gas6/YsQhaPtvP17qI
Ld5VrNbtYVX/FzeCqTyi2563tLD9MwRqk6Wm0rXXlWZ3IB3ew4aufV69+RXeyI+F
mU0AHJO1MpHg8ffThWweAFgRCsv5BbgmYZ6c/CFHbOlkp1bd4P8GWEiUywodCJAC
weTv7hQmFgpSoaelzn2RaAUEVo36Q2fXaSpIL+W/YJ3DTMKSfhVwjfodck5E5g3M
IxJKqbCRVbxzqq0DdtGTcTASwQjrnaTjskz1s0/r/A7HHMCat3HMGXt6mITI3VsA
IunG/rmsK4YQ39zwBjNkgi9q+YeUxnCZ1NCkZ0uu3Cu/uDEAGt6/twPqIWRsmnOH
5VHto6xjft3Q3PgUPDnYod4De7UkqRQAslb09OBOq8TnZY1u3zNiciFsXP8WF3Ii
o3HSe7Udv62i0lMFHcvwu09VE8RdnTVs39Qn5T5pIFx0rKcdUH9TzPMlZnpWIx8n
0YqUDetFP9gMA9Z9+eJy/XatPX5TGRj7VUwF3bnDyGHaAp0juhMH+fcQYLCvtfWb
EQ5s+NlEJSnMZWDyN9sQnHNSp4JADVqkNwQdStTfoVWgclBu90RZ3eiAaLdeusBM
r+YlMqQoVA3a3kX1JU9eqW5NbF8er9V+TqEGeCd1+5mME/Q93Y0GFh8AF3OcefdU
NrOTIFmYc9qxp/eg9gmmbeNRdGbOQaHhSfjxaGZJtt0729Jgi8TE7cBbb1k0ujkI
ADDN5IzsL3EviQP3CaJiFQCFZivO3TvngDi+w9P466d/1mZzwb6TrCf6xU8dMo6f
7iVDod1pUZJwxxEpRC8r36K8V3sdmNNbR+0ZZjkertA4lHpDKc1M1MHe2PDBrVx8
6vnFvnvYO6JJ6LVH7b8N1B3YrnLdriRUkjbG0DGupRx4939YiiM+LD9T4fgcjbjg
fQDL4YMLY40bxTtdvczmTvXdTAe10WH0EmWUB7XgF+TpjuNW3vJkcyyEEPo+Gjq2
oUyRtOoJMQ9GK8MXInz9IZHKEl5Ik9KpgH6kFfmMZZwZcNQkptf7oHXqpzn31M55
Is6C8OpeKijLtTWxF7c9G+dVRMn9ZKnYoPeSUCUpxSMfa34RsvwV+7nkMZYnQuRu
nFaMu/VvJM1cHlZrGDFDdCEonh3lWAwSc2pQUZMOnGQlQO7wgruXsU6HORthu5BA
TMOQMWI9JDQPyI4wpyyAJ3Prf9TcC6+o9AMlnQdyCVSe7jXiIKy7/ewFC0f11tu5
f19WT3ue3AKyfpjqmgO+584GbZsXUexAp4q6yD7yK9KWiYOtZbL97fx0g2sJgcWm
XCVpgWyknc74sY6B+dY4agbv8bq2RNZZMl9dyszTs9J8d2Xy3JBUwhN7t3wsFOAM
5IcghlydH0QiQmOgwSP/88lTPwAQqCqeEU8f9M4PAi3CdFv9XjtLwMqPyG4GdifG
qdyzGLRqGPwm+DBUzT7r0MdSvX0g76V/qXixb5DF5KKpbYDtN0RS+yw3bIF/ynQw
liRguqvE23+5aMpjPimlvZ1zuwkM6YT/3ZJnhwoEHeuanip6S02dogGgLE+5+yg/
uB7tGKRplFCrgxRvgHMpX7Jc2YtyF8c5AHrSsznsemhgAUUckL6rb5CpATv3zA/v
4T+EE3sznOYUMJ+pI+3xEPQh/U1402wbziWyMrwKb24je59AysqmBX3QGGkGDXYj
AkjugP1Kffa5G/1vxQDFruovGmeSMJaAFkdn194tlzwQ1jgHaDdgsBw8f5AmYOJ9
Yi9ne4V23g9l4QyeCuD7rQqNwsPu0/xCHnyf3mimysBP+F3m+T4aiL1VL2mnicFs
kR0AyKo8vgdpIpmL2WXwDuzig5vMYkmSY5kN7RRHdpcxYO8aSNTingBiAKNrhkLK
a/jfpu7t1Ceru5+V+Kg5HugGFN/RpqAC7d9dduPnBR78rtSYEJBfxHz3BHu0SIeq
G7cJn5xzRu5pBaEg2bMEZN73fdQWRSLqDAorfPQl+0mVc71chX57vuLv2W+xwAZV
MinC8UM56He/fjFYbePYoPMXR7xSuYUoeSDXpCX6AOavFMvQcEj5IGX3HR6zjfbs
EGwXv6zBF7ikx+s5tAIctqnounBiUcjasOjVzPJv/5l1ZMI4054zRfleR/rLW271
YTosNoc2YFhSnf6Epf06IjTRQVkeRin4kOmfGjWnjgFbP21zju1NvzqOKLekGBLT
kAbSxVjS0Ko0N9sbWaOXT5L1LPTDvKzz9x7WqawWQf9/VYQZlBK19TCf7YWAyei3
AvNBk7phLllFwxCn+KA+VSDAV04pxaRreohijQtuTcpA03oQVZhRC5zWJqRuBY1N
9r3ROkD9tZSErH/fOREV0JVRfKLGsacmr2I44Mf5mz9dbLN+GYqQSGHeZ3xVslj3
JYmaAB78W5Ia7wuwX2RAdavtQjqFpF4uL+FOgXKwWUEqmM460LqPOvcq1hM5Vw2t
GhX0bpmIrP2CKpKBbZ5Ikc1sE4ymFaPZaxLlSXL8PkI7T3QSXCrvqb+G0ELYCuF9
l4RmIveeNOIHNQCXckwOilgZzZRKSKcCNCK05SggswFb3qSiFFXROV5kIkmCqXIP
WC9DBL20nbRAgIK6Dah2Q1koaGs7hIc3m9JzotC3b6U6TRaIzhdiHP98eEYI+9OK
Tfzn7ROonfXesppB6EGBuLL+t8IUN7k2FKki4qS91ftaSs/srgFiAdnWTqWYHwDD
a174/1QFJhl5TtCd+FMzw4z1/SdmNhzw0Vlgp/kZy/aLqWxWVmhHuOGeHWbS8Uh/
0I5y5jllknnXRXj466Rx5JWt77ac5Lk5EIZ+YgBOIfuhtHs/wYDjM9iDNOKZvCSP
fNFzWw6FK7m+Sm5v9V5BSE5Z0LDC/HGzj0puxLVgVHGl+Si2ymdVssPgcPZDoLLI
BS06YxY/X7jXDFf4PhTUi7J1mooxAon4AQ4+5Rnz5iZ85QrbsmJbp6hx01zZ2gnu
LiwhnMva5eRE3g0OUtjX9+dRVMSJH/NwkqB9tpRSgFvqwP9KhMf03/ZSi6c3zc7F
6oftguz8Ma9iH4IYieJNp1fQcLT0AzdBSwSAT6l/OSX9vizZ3GCfvOxQFr+oGO/b
ZtKyjcVBk/MtBG/63AXOmKbQVuqsCJroyT4cv9r8MnYwc0EcnLGakblUaBxVbFfU
pln1gWVZjN+BgO/+aua+lFC/hpKx66H5mL1pjARJBm0H4TwM8mtq6jN1ZEszvygV
CptOCcfHVqfUmKaW1T8aklOQDMjIn++cx9zdr0vKtSIA6neocx5Nddc8M5scWe70
nwltFJqCuI6gjyC8xOK4waFmaXl232Tww39J1NwVpbNG4ZKiOhRRr8npKVj/dGev
5SkIopxtNPkwrbOHi4Db3bwSQJbeGOJekJV1WphEJMB3VSADHpzHt9MWT7fQ0quZ
5nSo6LypRdC6J7KW/ifpgZoOl/8f6w9uk+jFINQhXf2bokTnzEjcvmDQ0etL/ipq
x59N1a2LDUDBFdhqFV4tzyQGjBl5tkFsqjS6mp49xpwgur78gJEgc1KX5QRMq28t
jAoYF1NEBKZW3Y0+P1eXZRTn3PN7F9FntAF4bKAOlkYRSdNQG374jdr4HC9d6Szr
iDco6Fk851vi+IlNc3ZxtWBKCLLaAvjskBPlF8YemSNEDHJrP0wW/iRDeusVUzRM
OLunI8GnGwIWBvaew1NBx2/zc9MWt2c2huvoyXa7PPRL6vYqljCp+BovFhoo8NKQ
aWI4cYe48hyHLRMMjq5ihFBoSG4uRjFM86BduvpPsTDVDQTyAgcYyACirLW39hYe
sORnaPdWgqEsdiIO6nye347iILiVnlVVZrVdoSWWxO4etnOO7bTO+zmonDtiNHLn
FAS0JG3aRtGC9zI7yv5KOA9m9pwSXKaFDovycHrd4QuLOu1MgsyK80pBlK5nhv+8
gm6shza51GW96UT/qliCUGOtFxF95D8RtjsvKquZ3L4yJIFFpmA88Tg1i9jLY/yE
1rRixRTgQE58k5ijhstQDxUExtuwG4FdaWUYi25P9HZLXOOYb4B8SD4mdzC63Yzw
LFrxpOlfqpb78Hwv8n7VbVTexU00+5bmL2qXMuUImcIzvkxFTwZhhiTXmW7cdld5
O1wKVUzfvHGGq3iZD22EGHjPyQyPEHVXiZ3wYSYJdQormWjsd2w78JP69R5yX9Zs
8jy5PHFsmaKgbofVlxTbJ1zsBQJPRWfoiN6EvhUX5cz79icHxK6gpZ4OE+54inKI
3HFvzT940M05CNVFDO04cN7pgNeb8vHoRmulbG3Cn8qJ8YfSjtL7FZSfQBlJVRY0
qwmj4gUfKT/itSViOWL7BpcROfT0G7rbuolNB2FvHH3UTDQf2qBKhFyKdL0HDhsY
XMd5Cd33ggIIdhB3usOQvXLqu3ZC/W87ZSES8CTXdF0TCSbmsv/BdTDyYxLof1GE
wMGtTD+3VH1NLx3/zLvL3fdcYxPwDEIjA2KLNIT7G2XsiQgSKhnUgf/i48TLxaN+
yO9YKmqwuCmpefEZ65oB3KEbDxOVt/r8gxvDxyjeEFjPqi9ZWbA1wNJLZUWuFHwW
iyaMv/g2SLbx3CleFp5qM14+6Oke8oAU07n/uPohpl5Rg+6XEZCZ9K63iEd0jA6y
++B8+/Rpz5IeI/CTCXqRk8K4THX4qj84RAz9X36VEUw9BZ7pTfIs/rKzC+qTVALG
4XqrrLU2DGU1SQMt8dmbKptJF55h09pwyBt24+Z7wDHRjB70ARSCRJelXx5Jqrv1
tKbt0FuMgjs/digh+m4B0y6Bc3rLUdi6qBuhaCQaKCPc5nLx3qHdmiXJYeqo2pVa
yJ+QftqnIcJ2StnKSCxmuzSJiZvB3tgkKTdCGy4PmyLcrCCLYNt06wxYYdX3QuIu
2noNUMWbJMmp23pKXADk1EQhaevIAL0n1n4fEaJLdZITNXlkNVVsw4mUV9E4cXPP
ArRWO6BrSxjBIA8suU8uKo0rIYp737XruuPg/9iIrnONPBGQhWXF8I6F5Jvc13wv
RLO3J0eHgDMaUAEJ1qqq3L7nOtFXQwYkhe+OHSRxE/K1m5oKOoVWhzAk/6SHUxX7
ARhgpcZefWjtuTDdUsQY62bfP0oernklMlRS8G5wSFjeXACNc7UvgjqP7hwAXkF0
ps1efLILpIOlcN0nvDdP9V7ghzxRllN4x2TYELOJLChhuWX1q3FOjvtLi+TxjND/
Qqf1+J1tWfk7g+5OrIidEIdYpUh0hjjjRCcic9l4TdEZmAhm5FmP0mhfmLbDpSJ5
JYnqlnz/qecUNGKc3TBqzEaSGU3BzWJa54CRi/n85v+orbjY8QJy7kAhITeXLqzf
h+ziE1BePRZzygBYXFqsijzJLP1RgZAST/5fsQyHTGdQi3Uj1v8OxDtX0N2M9BHK
G3d4lgmu09FbDb1JGUBzrdS7gnHUP0EjcllulaE7TrKidR4i3zsVZkUMlwYDxiTR
bfTO1hupDnNzYO24tRcoBwGVHqXlFh54rr+9WgCotyV8eG66mMoDxQnrepXEiUq/
Ci1omefNG+HXyXtegXQi9D0oFXm8AxcSd2tR5zw50+kKN0K8mnuo2ylouxlhIndX
KVmtNxzfIdHOO3ys5Re+FAYC3aRzMH0GLgGer4ccjdcjZo3fYgJgvDxGZM9e2Hri
BdnLL8cqdJUFsrHCvZHOb0NqBBpqIw67yWehJXGKQ4XXjFsRMZL5dLbIlLwHz212
Wqt+8SfXVLl6Aki7ybx0aGErsn2dlYHa83oiCddQVDneMlyRJoz6qc56UTmaang4
Tz4AP6HxGLGSvwxenSxW840MgPqVUbcTthgf+Fqw64bh1Tzy8orHTkCc9/Gx8a3K
k79RWd2bA2tpAkPfl9XlHUj5wy2Z8+zmVOZJZ3E7Q3nQu+QimPzdBTwEWRpAi49D
pWHELkzPR7bFevXwYZEkF3i6HXmk7o1NNgb8ohEs/43CYJhDm47dJc32Mg789xdg
UhVDK1leEAe+tt8B80Q3k6jWyohFaZsAaYfWWUpr9bpmcCW0u7warWaZm9je94N6
KpuQqQ2XqgczpMyJbLV/E4zsR+ADL9iukdXEynDzFzbV6bj/6D9mtCFFEWR5htxu
6G1kZNaEcPMmGIAX29hdGNEaU99EIITBFd93nUI4hv+WT4z7xY8MgA/KHPmjtPxZ
DQp1mA+Yai2bCn4Wr4d03/insWNDr48KMgteZVDhihvpxCD19WeN2jqQb7r7lrZu
RvqJIMm+WjlmCbX9dx1K2bz7sQn6PNPYkZSQ3QNe7XJc+VV9PVpFHS0D4RaCEbAh
1vlWnD91hL+2dD9ZeDhB8LJdIlX3mtOoKqtnfkoSB4Pt6PApGt74UqOYQAucUv9I
9EBdTTqUnRkKMIGtJGqGTiWmz8VupEPuj+FBTAeqrhQ75SbpY8mTe1KWuqhFHDmo
OPf7ro6nSHKynIXdtOShxTFOB2xBwrWZhqPnx7xKe01O1Gqwcm+OEWHNA8t3s9Sf
32wi/UoRpkJGuaKzOBooevBZ3tIScL4MHcdUB5dN6gPGl5BEiue8qocQ2b9juEhP
uCzFAHEqdtiNzY+K1487Vo6bnFPPvTJWJME0dmvlGCDNp0cFILaKBkCvFFG1+Lhm
+DcSlwIltXYFeM+UbkykDvV+76AIvC0sE0rvUGqQ+i0P1WqiOXisirItE5Fw5oaL
qw6ashig9cIGtTC7Xh9KFcOImQBeynve5yByeKb1ZkXdBF/t1cMvpeEPaJaZo3ze
mF6MFauEJdb6qGGbgVxEGQXeqcGMQo6Zg9VBn7ohyeVYduPgKKOqR2xz4xYqAjfH
h3wNhfhMfwBxQCIFH97A+3MUnsrFHQqBp5PEPmcxU63sBDU55RujbxwkBqRBfz/9
DKzj8cfwLYhuOSmyfOrR8/udp2UrEdvsGS60o+/TeOk/NsJJq4tp0AAkcbtRYQHh
29cA/sOds8jjolq8B9YqHVyhebiWAX/sSHMRcEbFurqT2O4zpdw3jvQHoEb4hMSV
lPC73Ii/4O0JZkRq6Mfi6xamZWJibe4c2WTnu6bMNxqm1iRuMg1x33ugu4Ldu/x0
VzAOJjWnlNB2GwtkzHPsgnPhcehynONpct2n5F6eGWJrijyXr0N1txrGX2N3QZXv
Va7yFe/a0FTsDcLws1zeiD6PCPXsPInlVJSexF8mxJ0JnR5bW1NHoc01kEoqRGOt
BfOceM24G2phuccaLgSW4Ns0oE4d5N5PgK4uVmZd30EtLmCVEw2coSLXR/lgYPuv
Kn/KoYdVhPUyshjfc+cD47zougf1bxYEz2I7YxXmv/h17FUIFqTEU1+KdaW/ytGs
NtfaiKTCzdBAkHLpxAkbml7OECEnOgA+NM/Lvhx9soPJUcTU91hgCav5I5uKXuog
YY5tX8YrsWs6u8LpA9+TSnPLIm/ZqkyhOHrK21Tz19A6rnzQn+TEzFQG2+Y3NuG8
ArX19zr2XZGkUf8Bcu0HUd9p7NMn0woyoYHZv4R1hjDtMdMGy8EWdrQi3U6hjIee
0yQPOzFXO0CJidgHtIa8W8gI86i5ub+IyxBHR8d8PaI3+YY+LV6hKNFJfjDJM8l0
qrOTXnq7oBhjamP3qrWOlz9IwpqjVdVRE6pMgKnAd51z8nPYzyLh4rFSsGa09cSM
FBeiQIyzYzIA4umdBqh35KW2QNgRy8rZIPaSFGAcSDLsEvOFIfpcyn2lHevlwxXn
bJmr34RBY5kIjhCnI+7ewafXAdLcqI0m5WOyQrCUoIQBBjVQCviRDSRWOdoVDhh8
z1Y/WxkMhw0BRYvhpXxVNonSzwCMvDIg9rQlYuVtmSb9ca5zXsXIIaWPSL1uT8aR
/vyBxD0J7/LdRGCakvLuJWriD6P2246xEHV1uN+XLG20ih5a6Wv9t6G8kFDtwcHH
J+rY9Y50eaSurALd3QvVYc6e0vOyXQUVTtFogeF6H13A8LtUueiwoBTvhd5nfiHQ
lBsaCJlIQBwvpMgF3TsOE0PNiDq4cNU2Jy4Rp2mpQVaJ4ODX+9PGieTy5raLYVkI
OOn/0pH5SYKu2nWy/BEks9iOiBs4YRKE0o2xw5trFrahd43KckX1//HXyyPixBxF
nfE444mU/Mq+p0YPOcnMOnY+UXp4S2XS+sIfsGNPXJI8TeeJYw3Ct9+jwZpVz7yD
2YLJ9IeYM1JNIbAB+yzFusdU+eiyS3tSpUCSWvqpVgsOGMYtxka1vJM7WCzFrMuN
6p8N5VFPOEMZaok/Gr5j56YIKcn7pQbRBxsBevfPxwAJ8YbUF6nJkmwOwddgKgVg
pZyf085pPf4gZHTUL8r+H+2geeNPiXkKjReVjFH+1CM16+GbWqnLu94LPS4HLK95
nOHj/oJ5O5hXeM8Vj3HbpRaQ/vdRfJifb6lO7r7Az5OhUd/jZaJuuoyRnSusgKYA
BfTN47hN9HqQKdtvldAKI8iRJHpN2Y8F45lTsGMWTv7gkGf14RHnXzXW7kF0mNdF
T1OI8QZqED84th7vaXVrtOx2FupbPwvRa7U3JulyYHdpK8mBEGM4HbnT+T3n5PK8
EwF7VvJCKjobh46AAQYMPjTJZlxmmshOdbWzLBEWf55uUPuDejzdnGrYAqAaI7rj
HHdKfs6VQhsn+q+Q73VbBakcYgrhJ7R9NQJHsb7i9AcbJ+lfAhkyPp4M/7kYgEXN
vtUVDf4phWjNtiiOEOyyUdDNt5LtMbQeeQ8ZpEWKPQWdjmXD0X1H7SNLHMlhLdy8
A0pYHEftcYaKTsg7Uveof+OHtYBunHu70Es3IS/DRxaNa9PAOBL0WvtUha7hVQbl
J8uqMqT0PfUYUjtS66ynv/zyF3+ZSyUuEw3iuZp1dI+qOhK9NV8F9CcXwFFaCmov
xeQaCd1pw8zkQy8XKqp+KXxTw/uHrocPA+A5FqZZX4XIaaeINr3hca4DkZDMK/Bp
Xkd7n/1PIzLFTrRfH3L4lbsueVcvbZy8qL+aGvY21okuJxurVvtD6xd7BCoOfmIo
7hKzVrAnQLtFGTGnbsSGewu5BdrZFimApkQ0vFB00/JQX+SIMp4BFDjUU+eQgyXx
quxPT09XmjqI0aRw3qPUflwNsBmC622SWQXPQLA91DP5Pi2oitzJe1gn/8a7+iNw
kg5NRPlNG24HeWyRqn0Q1yaSG0i0c6d2rCAN//mZ33sEAjPDPWP0zeqH4T2RJOJt
siV427zyur6caQ0u1h5K5C1X9MRvJNl884trE8c2I9t0rkAfdwn4MezKcGkmhh8x
peGj/9htIf7BmtA7nYSWqwH98/uZzHNEb8W4esHHJ2+wIvT8Ux3nJyIWrZ2PpMW/
6Vp6sULgWCGuykHTP+nw5SwCSi4wmvZ0G1jnDXBiBNNcpXnxFOzKEeDCCXp02qRJ
ebyL8ykYUweCg+PrAptGCZP5IUx5JXy2fMxdWTVSTvMldc6dvrGTupuQfmv3gn6q
YgQE+GfW2yWGWTwisVlXKg53kgtRIcmxFZaRZxtfUnQuWvQR5zrNe6jfzCQ5itBA
hUM1W2iLhPR0HZcHnT3RSU7t5F0VKRYM/RjmJuc+H5mEqIDyoDYd4pSn62LV3+78
ZP+unyKlB2TZXqmGML7Z2lfibdDNVttE0EpvC2O07ImCalu+nsDmZFqJlG4867jY
RJllmFOINJiQq1dFXUDE5rMdRfCyLJBySAlZxTK4WCDppP30eTrepHmo/+Y7cuEn
NBbL8RIKBX/C/C2RWmPSAA7/lEoUaqmi1ji4suTn+ZUuw8+ae3Xnyw9Ygxgnzimt
t6xjlbr3tNWYFKKmx/IDC/sVLvZRRnb2ngMgw6MVy8AYDx1LzftLGzvgaTq94FYE
oy4UugiY9y1OnNXbukfCimCMUw6askQhQAUEj1RcgQlx2QOHWCoogaO5ZJHfdHYd
+gs9RrWZn18bOVq8j8f0waCXEcIXYKofyRixyVnME1+lCRLu3tKN9b+xEN2P4mCw
A0MZHP65Xr0iJfLbaYit0T2reeI7Km+wb+QBXLt7oQNut3OWQHRMKTM+36nLdNkh
ANMcZX3Nd+Dc7Je1g5EnHUjv0d15BxN3/v+LNdyiT3JY4BNAyC41e6M4BbqZlmZi
INavesRq53l+19oE5P6mYRq2T7SZc9H1/HIUYRUXJKfWRbCPeO5X4TdwGlhzq1Lu
c7jSxrzh10dClqMbKMtxrxnPobVmRNMA63DpzDEZH2xMlhQOzjfxh0KKg0ZqH4Xb
a+qY6nxYiJSlJslgDIU2MP83ghxUiqabjwhZFRuZZMk+SEn4w2dGZfCs3cIunEqv
psD+pmyanwoI6x4XufuKVek0x0+Jm2aOySOBH/ol/A9Aoj5/N98q1SVMi7u+yZ0e
mLAVhfXHj4n64f8/BuDo5MQoOhk6OSqc2J1RaUXLEoKjqsG69mEo6wkzrZ+XnDnQ
XF630O7kCkOo++h1FbhyzWBWtowQGT2xjI2/Fgr8fTgQSPAvx0HuyE1VDjPEo6lZ
I3QdT1nYiApRvSR9CPW++XMEWd5YGMf21uwThlOr6HJpQ7Suo0vD2wWlhqS1ou/p
cg3lDu5h3+zPpFMk1Vs0lqmO/nK7P2MsPdomJ9gY/PqJpH2ILLZ94Fnew1phQk3O
EI0mvT3njI4unLUsrA8uiAQbIVe8edzF6cDHGUJyNxxWloKhtQpV+ySZiOmsPZzF
Y5SPUkr2DLD5oWgVQgN8rTAEJ/vfCxGNqJUjLI/EcJebwwVP4l9OICzVDvR7lISE
9J8T/GLH4SpXJp03fy2Hl47W9oxpd2oB6fj/GNE/pCnLgViVfXcuVlK4Ldon7p4u
d4UzEL81yVP096JLLKTGsaMVFsGbVGC0WO+AyYfWYVbywjD6K2Dwx4Rg/znHs09z
x/SNv+07xfBaJGnNg8KZdOUmj4O6vXW0Cch23q481/abyxZStxneO2n0g2jMOToP
NxPJ7dU2JJzFSfXWA1LR/A6EC1DxRHsgbrXZWUcF5D4aMr+C2kXf9QdOZyVFZjQy
YfNK0sMUSKwNWe2w1rRYKNa903XlcVHkQao3IqLw9GyxTmpe7e+9vR6vX9DcSntA
Cz3JNYPDswWSfx0NmarYKpGKhwiB23Kk9LmodadmNZtugTV6dheHQd5fbMEIBfz2
vnvxZUzknh3YeKIdeP1cRFJnNbtLMmiFw4F2T89x0l0yiFmMJitW6QXu/EQiio0q
E+9t9aoHfdGn/nPmdUoGZ1xLhlnYyvD+GOJArNZSLYT2TUPp6QBWk6iHfgmpryi1
35PDqzWXqOYfIzC7NQj7B54437TpG+dgT5u+LDFKpIU7q25mYVairJCqdHHOE53E
/Tw8TdIAIHYwlZbWODH+SOcMZ6mb6+dIaROwQdNRJmlsg1SMLgKQG1Ebko4RYYkk
kW69UJ454AlRF1yowaGVcdg2bvx2ywhFfNQbvxNE93q4RcPWTVXxa7nARIgzbeso
/5suDVXdeHdijl9Vpgdk/z/L5yAMtWkY1FkvGLM+Vyu/tPLA88l7A/g8/L7uETMc
O2EjfwHYFMveF3GwZ7b2Zhyc1wr2MtTHWFiiHtz9CVeq08egUKTwPbfqQ6mR+H70
uzJD3TWArUXXTWu6VYCrhYn5w1TRQV8H16pef0HxUlnHEVEQFeGsuG4b6nwbbivI
xWIjssZZ+L3h0PKQv/n6i0IRDG0Mgcb3oNwgGDXQ1RN8+ZVH3DNJNuhe7Udo00fL
7Dx2cwhxKqY8J6VnGVnK3aOHGkrKsqpoPoCdds+c+/HDNmsgIGShLHmngB+bNzlg
2h+RFxYrVjIAETvlMeDqW68NSyR3gTQslg5WyD3zZvN3TNtDnppgKi/cbvO+AE+L
MEadgkhLVrUMyH69thXg8krglTA/0qtH25vM4AL1tBzuHVWWMKH3KLQ67Qwcf2Qu
CpnywsOjtAR4ZmEbDH7Xdrfv0+L8bfpEzzMZVmhXW4oGXpy0sSnRVyFhMGlA8CFX
d1Immtx8uItJyfX2jfiqkws3NohbhYjBRrT01v4Dyi6HL8pQVKZGuB+yrry0acWZ
KWdYso8WqoRSVx2eg5EEvlGioZARi/aOl0Dq8avacOXxFWDV79sza9HhJkOSrVrv
X+q/47JgK5218c/kOJ543bn2gmNxPLy4YKmHCHURzpeV+22nvtdTJHZacoPyfCE5
q4L4Gi+GoPmKtBB+iTFX60DXyWRTaJf0LD+9lZOHAcJG8HsVPX4Jazk8uIrbjQrf
xynZrGDxV1cuOnq4jhjZ+/5Fqp8hB+ijtF9Dk0E6foe9ZBj5z5J6BrA5/dQvuXhC
LvU7J16TgLKr6sjPklH/0FtGCOANav9WeXKPqC2sKeMuufg0hzDL9/Zoa6XGqTz2
EzXGxDf3XfxkmRR/q9fra0dgqJ23ftoG7prTCyMREKuaagYujT/zP3ChGGol1TLZ
t+gSFXI5gb+NROCjt02u39065Aba+jy/Pva64GBx3x0WxRCcAD0uBti5O5x4eUrS
DtGkYp6XQ/d3ROg1za1P4FkyGZW1bbJ12yNPyt85PpZTg6ENJsx+72jYII3vUde2
kmhyqTk3ASWCfz2ycpx2pz7uxl40hglcKtXXNHZIsPUpiRWrtZeDMKY+nkUx/XIV
JrvXLfj0Kvhh3ZGx2bFu4z/ueW0AeRZzyOmzM0o5kd1QdaoXXj5jY4z9G7Mh7j4H
SZOSauqr7+qlLuBEctNMImlV4rJ4cqj6S1V7ZJf59FynF+CQk3XtQFtzzgX5y1tv
yTrue5nngdXEH4lknTfvcxk3TFJOl7VogoJg7g04LBKHtYWCqUJV91VG1Cpi8PxQ
SGt+EldHsMeGSuDCgDW7C/f5XgsSiM0SvVQyHQG0Z6GiP51QgEZi9Txg/JcAPAbZ
iIaTAarRQjxHApfkb04X9kfUMCNerYy7go6n1pCCdybdnpeDIH3mp2SluVCs0Okc
oecQf5qNdXsgU4SpIYT8tUbLJ4hBLXWlX2WqOSiE5r8zQ6DpAvVmcRFcV7HRY3bG
sKXsDvmDkN6p8Pnw6n9aeOyvRvWhWlNn21gJ5/c9Yvc27WvK1evTRohnRNpkhuyi
1UUhuviiU3WOvvvees7XxgFq6k0rUZoJzJu3z71QcFz0nQqE65SYxlAO51dqYq+D
xmqAq/eUoDQ0rDNotOMKeMN6X7xeOM4kJyliqk3HTr45d0KJQyxyHlKB/OYP0vYK
aLHBUJgKIgIUIbqDk7ks3Ledsbf6hsPuC63yvTMat659QBV6HaAK2lCh7o+yEOOO
d12VptFibd21bDZHS31rLHknQDdPkf2rNS1XuS14nknU7dm63lG+LSJe/kdD+JE0
MjnjLGxfbBPTlROopVyeNwDQyjHXMs6mhI2RsW3kk5qbhH1C46CPPg+omUvwp5L4
tyRDMWzMznmiSM+6huaL3+3Ein3xpBs10Z2VmutLak77mGgy61Ope5WfWyvNHmZX
TZRjDAFqOCEyzQ7AKRk6vy7d655Ffyn1wu5CTMr/f5hIxWc4jua7/Rjy1Iz4a3h+
9SZzZOviYRPrM9kusDZG/sko2cjwwRz4OUguGbBbLCUdKeBLV752lWI0eGK8bpR9
ZuNCNfdsvjnu78taEt+lHwwQsKJumGB3MyYrBYlGq7wYDBwPAgKoOda/Sp+l4Rg0
BtmLF0IBxztzy7+S+byXd7uO2CB7p0BuNw0f+c0zLgG4V4ijvoFcig18gfSIt0RY
Nj2CSFslhz941jMnI39Wr3LzYKAb0ZHD5h1cB6dGI5mHwibRcVK1k83oNO9CSQ4U
dFwzmjX0tHS/4YenH4ahrXe5UkugIWeILhanzpFI664eZuIeafo5szwsHIpi4Mnx
m9OiAsmGddCseZ/gScLfxGD28o2GrsMX0fyCyM4R0vZksQ/TtX327ujM/M44jjJT
kHM9LxMz+d9/PImkRz2O+PoJgADR3HkaQFtNE1FgiczSYWUquS8oYTyYrTv3Stb/
ULTkIlC/SkfIdUkhJtrwcgWqahIfJ2vNb7+WxraeJy5322DDqMZUI5Q/gjQzSihI
dvErxKjEvsDWwjftdf7IIoGZ6cR+vm8eskzowHJcNBLfuKRFy4myspH7MG30nRbe
CoFIeNwBkWtA656G9EvzIHunENNeNHo4xhdrRI2U2yLLXj+NQJfsFaa3Rmw75+aX
qFAY/MHn58Pf2PTEuUeAmH6YbwSH2tjrhEpwOPM3t57rsZ1BoHOF7wGtLofDXa8i
QMVoIc84rikAGffFV6G2H8wCzY99EIapVHFzx+jp7S9mrDlpTgICqjRlUkyqcBhJ
RcxJf3G0dTwBQtQLqfhlWXzGg3gQgXoW251sTpg3NbjJ/Y3eMyAN6r3hhNhjKH2Q
+CX4zmIi6E1YkjJgCsB/7+/Hl8sGDV9dK8HeF8tQxQ6dcMe3Is/3CIq/NuPzDG8G
3uH9GtzOP1LPxp5JxoQ87+2sXW8DFfmMLG+qLPwOhTC3fzlI+5b54J0XNeyKSQvR
+AT3Ch02ukDzNgX69g/nPvjCn6YokrozobtbHQbopyoocJbNTh3noYiT1Q8ygb/3
aUHTrqqtZ6xPTRxOq2hxyJiPgZKQiZCbP/vUBs31j0tZH6ZN0p3kgNkcdFTomq0Q
9bryk1hfdMSxioV/Y/n2jfQ3c9OSKd9cZMrZgiZIgFkzvI4FfSkYGdt5VgpPiTqH
lzR0eCvgs4bjx5HTbu4mcqhQER7T53H1/evjokjNt35nYvw05pgxmyw5NSEcKUW1
pFPdOe1AZp8frj3pO4s5IQNN2yoanLjuqc669k3Rw9MGSJfIRL00kaCMYsdtRHHP
YUQqdHsLwSHy0KCJXHK7owdXSEIy2j+TAzMKfJ2O9kBT2u4EesznEg1xyFz+Odj6
pYjluSbV/jYdPHlfTJf0BUSY+aR3F9HAaefiSFLaFHspLu8DHgzBeCA/Xk1lH6jg
lRGFIRe85NsPRkt6NrIJF6VibswXVjH2jVL0ZzXtGKiyG5GJ9IlZpPVrhUp6grj2
p5NVTTmGkInKMQZznWgHt00dimx5zeaK9u9p/RsTxiLsuHOV+/pZxFvnR/PaQWNK
LhBgw7ndDVrrO/Br3Yiz7dn3PNNP9XVbtAOi0KJffFKG9uvZVJsOIFiykbZ8X2sc
UKZ02imQj5a4MbRSYBMKz7ZRDvXI/ruQh1NM5ifw+3cHhMRyMmbNn9h1+Mtogh0B
uy+pfk4TBcnA3NBfFb4BP5zXTzoxgRZMpUxZ7TV/Y53oH6O7CtZzuC8qPrKJgK7X
vVn1JzSra7FQ9hIaC3gHxiXDqpFeLXgxR+o7Uc9isMmG1ih9IPBQd74p1FaFLbt1
LWdde+/+pdMK5Z9Osh2472OHNnscF1vhL0wUrrrWIJ+kCBhIQ1mX1T4K3pwIpAqA
269DiMVFVC8I7oPqIkatM78NI0HOf8QxkYy5IVDdx1FXqODquQD7/ghTVhTKKDFg
P6wgveHTU25EJy5dAF5QAo08kSRBORMyyZA+ZGKbI42I4Uqz3tWYja21QMoDDbZh
jAD0WdoN0ubMBXiGFy0bUhAotwdyv1X0fo2TCxEgqmg4kH2izT2p80cyaJkbaCfY
sVJoG9hLHDfpQk0lLnVA5NhNbzprT0fvwfH5IV3v3TiBhS4P4fWgPLVc9pUao3IJ
5bwwBpS9m5BJhIS2sLVZn1n8eAckF/y1qyYMieC5wQcUQkwDb+AOE0A72zMS1B2p
Wn5ZzhxzCBW1I2W7al+YoC+VPILeCfnoxd+DHcOBsWMWcG0wdLCiW8b6U9uw5eQD
5Dhq1gGP826B+GDpLDnq5TZKoaxa8PKmemUZ58OKAm4kf0NJwzocwH3Z3heCiXQa
SXKIcmPmQdUJnX2kb543UjsnPFvj8O2pR3oCFj4FXJnUCp3C8iL5CPeKkGsaURDi
FAIrTLh09iG6eZDuggM2uL7Y2iXIw7yVPXiRDsXqg15kpCYrBgWYIdfhfrM7XxMa
Coacq9fvTG158vwp0GIK+JypGnB3wsJVERmjDIh6RwjV2yQ2Gj2i4enq80QExMhZ
gtdVnm1Yn8fvZayyyInnSA5QThguCvjqJ4e8ssXhk+kvTtFB8MzAhRE156bXI/8Z
uB9MQm6XYJXg0RKMC1l8urjDTFyh8fY3d4UfDeT04DPSVvazFcT5FJwuM5dyx02r
2jo104q45N6+N50caC62Djnmhx9+/7I0M1brUMxVnbUz9mf0GZX+utStvscsguCn
qiWGIOWROAFjMjA+lxYyU84BkoEOrcUKbn0g1836DGlmIRgal8n8UR1vzmJlbjii
/YqZjutyAbmgWeNaOukGEviikRbpBQmf/46ZxIqWqqKmxOx+ymrmdoPT6FZjPSqH
8glFiypBPhZeBlqEk0EBFHnHIbd0IdDpdQjnz19uLWwTcf//bHEyvhnWi0pgh+z4
GAZij6rx33r8E7P2o0OPfIQBWrKi8cO7XSUk/iSf+9cJLRJOmmsTf76o9masFBik
7Hx8VbbNJWDkMAVAr8wAf4TdsVDMovdTe/IP1nSP7fPy6PV/tDTc0U/X1mWQmeiD
0dmQ4tq4iaWW8/9atpUWhndJYQ/MLmtG6K6W/KI74L3811JOMVDR2OHVEzAB2pc/
aBhdYngBTbEZ1D1GcsW2tEq+i2lgXk29UT+RQspEf4WFd4INIevYFb4alfCI62xC
4V88d1u8dKy577lnVJ2PWHnQcGGRiIgcxlGYFKwPSYSAD5DtWHaKV+/c1oRu2yik
DnW2HYK5ytomOqel/Fjk3Fvkg84+sbovuGpBeffwXqRF/K5ktorKBHYSGLOpPdx3
pXprUDtjNbSo/NQZousynXn7oLRlk+KlopDSd2PtY8caDF22ZuHIR7ZysmW1ALeF
EuBNB3ZqyuG3fc1r6/Z/oB+EeA54+1ILcfWid5KtQTmC4PsZPhnQfhGG7qfoko73
C67EwyGwBj3ZjzPACz27sZRbCQ8X+bWt3FjDG4twFI8OLsO6edppgHYDXFotyjGq
MukDbL7DlMQsZcwMwoUf7OOCIdC65lGFMSBQ82fym2fSP2Og9k5Np2CjW4hXw6Di
A7mpvTe55RHfxhPeTL1YfcP8ndAOSrV/taPY9tLSGmDsyt2y0rOpkFf1njuZmTqn
UuZJ0z/JYOtlLBzmNkqFvqKUBTJMBiif/eoqXekg9yEfj3iybLGbom/je+9ZpTus
rfSUf2tdYd5y9RFxFzBB1SNzhsOxrmHeSLIZYp7EpowT8NSJcCeZpREzq30bJnOT
ChS5LY5qZfz5ARi+KTyX1TAMjg8j/0ToHrvKHSu76dLXF6u/kOvBX1rwE3QEziFX
wVkhqMCAOklIZ8idbVRgiaSKGaHQUodl1GJqGLYu9GcuCobaJjxSnJ4Y3R8pWs8J
pjuz6zIS+z90ei5oLEuRNWKbr6q8hTLdrixKyStQh5d/j5e1e+d4Qb3ewnzhBLis
4vH8VXNz6xLicCg3rvhxGOadE/kP1EbxE5ZyHUppAMvjT6N/Zs+uOMaXJGfwRH4b
WvDiRzAuVNALOT2fOQRt3TQIdcU0br43tzSbzqRZ7J6myoaCHpWCMVf8OQJrOJ9M
gVXw/SZv+NEqdV4gxoqt/itFWAsn1YqgAUS7QN4UCJlo7t2wGLVfdoJuyCHO12J1
gJCX8cAOVwpyPFmVCdws4oC0m7+xpvg1U1KnLze/8/FghpPj+bWJj9lpjgfu62/A
k0GN0JusvwtKy09Dp15QaWUdTawOQaOUgwM+WWf4n7yDEOwmq9t1QbrIW21XRXpK
SG2RdoIp632Kf8Oq1tR0w4LHDqtfcMguJxC1MlOimL3vXRXpZ7stK3cnm4pNco6I
Ft04d3wl45O9Gp1YfYt19X41CictNozRG79sb3tCM8B3O31CAxr5zvKPVZy60ZTK
gBsZSz0dqeDLeejUZnzoV40vr6TgznQhZUBcS7Uw6g45H91AwFezA4Z9IcTl4Ifq
XtLMzCJ8kl5zwiNX/JHoSLDyYQB0R/yX/kHs1ch6PC1hZ0Fj+i5Zl+xFpEr4DdzW
LwDewazY96TC+s6AdjRb0StzMMw2HXxYsp0jqI0Ty7xFi9R7HA+Wiakm5Edr66+w
NWhsJVsbTfMn4sSwo3ucWvYzYcEVTYpN6xI+J0Qdbl5LNr1YsLqLBEYYZa/Qzx93
tcJlV97KhR6iIuoe4CeuKaxvBQom0cGC455v+ZOJMcAWZMsSg2fC+eHJYRFIkvFC
ZGE5FipROHkvWMPZ+hBOgna98DZBA35ls71/GH7JLwTDk7O5L2FVf0F6sm2hccQ7
xDhIdCo9zCp+TuCp7dSHG8MOMNXwitGF2Yn8Y3bVAsRPmEUwCYwBc7padIw62b+2
y9SMP4nnwThS6/Eeb+7+MQUAwaztFto5hgHgtGxIr5bnXjTIf5nud2eSN92ovLcY
ZM5DQfgN6DA78T541vdiIzoLnSgD4AneIWRvu0H35VAsYP8ZNMYPzfLQ843LBEF8
J6ljlDAG0QZ6F9/Ap5TnymRhzLIqB0O3yDDACXVnoWlNJBYA1LeV5Epyx3xG2pi/
HPEWZtpNdYKsY6MWFgfgqYReVqPtAM5OumFG6aZKQDy4RFN94XzuPm39ksTUIyCg
ZPXEVnFbFyJ8I1Au7EIhSAKkyUCAc0VpoCgmIeYs236ffqPmxWvuIhMnOlBdjmpB
4H+tjCncxzc4QXgfU+gkcyxUTquPE+wTKcmn6SPWKlXC7nxKqxr22CJ/wn8R9BfV
iT6qY1agP1YPFs9Hr2+yhSc+PQEM+QCStNWXm43YWv43JzKdB24p+EjE4RnBvhhf
XoX6AOOKZNA+wttRTmXgaTUYzEICsfDw6Zp1A1FKSp5oPHkqvT1gilibJS2SEiSo
Wk2EGCC2VYMa5fiM4/tW+Q1nnG2JMcEMN3Iw4OjCQQ+mOIudofAD+7BwStW/WK1h
n50eSHoiCbOAznt1/ZaTz1evFx8HIBSHfijGsy6GPuRz8Qf+/luJ/SNZWAYKCual
Bb+ncHflsnOg6ldCgovt0417poShfUDYi7rh6uasD1a62wiMZtDFkG+4mBKI3dnm
uWRUb0YamsZpV9WZoNKthmU6yYDPe40PvWjqFBWUi4gVER5n1RH6jo7iZ1rO9NcG
NzRcC7gM2qPgMnrf44K9LVRnficEUMCisC92m8rOKy3bwSAqlV2aHizt0i2ELYEd
dilg3rDCTUyCarlaP47HEh7kJpqrIOKx9GzHzGypFdCCOTZROCUBsjoVKjWqsyfa
8dTXEvtTJy2ey2AghZ91AR2lQWhtKsaFgzTMq8+NNlCAkljT4alhM9YErRfsYdhf
vJ8aljzalh0xkXIn/qTw1tJgIviqWMYlRwtz4ai+frhuW02xygaFOBTubw6tY8zZ
zLgbdyuGIjgYtmgp+4JMZevijdw2YLcKvKIRZAgByjzgGExl+tFu8lJKGV+E5Lji
mRAZYHzrfLnSL41UoX3hWg2gqnnLYnTQxYRYy4ciUPWP9ndsFhFII3lQ0sEWf0Hq
CTkUzueIiHQjB+7RR2CvVpLngfS1pS+nHprMCbRxT6lQzAJmt5yamv5fkpuSLAnA
wZOdYcNVR5w/tKUqIb0ojjHwJMGr/RYjVuE84RfPT/4AXgHFkxC9CxKUnieYolTH
w03g3XleBRpxa6/BiIg3oyk1l49jlAAyiqvzNIqB3gE46v+6obbuyTKuOIWgG95D
mwMqnPm3yRkSS3F9+QF1eNJ9Ykt8pPjTiFhSbHMJXXhnNRQykMfRyLzGa/JX7FRB
hA0ORqF4X6fhwLnva8pW4VTYo8xfgQyUH53HbWI2kkq+yaWqTPBBEshdsyJjfhyU
nHYAd49gICk/NpQnVRrXtrOl/ftAcp6SaTXjvVBg28sEMmoJjRbOW+SRK9cwM+Hm
lj+YZF8y8rkIt6z/GZi8ZlX4J/8t1irXNxiQyBC1kVxZcOEc0zHPV/bG8gRTlJPG
Jt5B5DuWBkXpHkcruQKlnqYPMh5loX0km/PdxL8KkXZudVSiRvVXVJeY4klp3Qes
nJTt5+YxVSo3LhDfAS2PcAovrI5byWNmhXBUYvgAtGs0JyeLTOoBJlAKIzr2JBpa
WbHAVV9MD1SRksjas+GdsDamZqEACiXIM9XJcB0eDnslIfEQJo8quhFSBF29HK7F
2vYkqN5yYeHu9Ri8DzjBbrepv1+8enZmOpo5RSLG22aHjk4Nn/QJqfiIZvVi9bzp
/zEexGDVS77phHZxakWXfBBAWYFK3GVFk0r+65VCEhlOdpm/P60szzVsONdKU5mh
2RXlcFYyWoOg8TkiRNyfIpHJnGgeiqd9tZnOK9b+k6/zVZko/FaQUMYjux6bK3PD
M1yasauxMZicMerH+7W0G3LfjO2VoOaTe4snbmMgn/7nn+JmKCYyfPrsA6cuEX07
BMdOTJzxRFXSKFXP8G82R91+LqBAgkWjVW2CCPb0U5kVbOGsPTkVt739GK3v7jje
W0m7PozPOcZP7+7FuM59Rg9T9w4s0Zihg+r/cwi9O9qYeP2r2NDaWYVIcpMjKplu
bREoYLfTYJOXQkYgg1+U9CZbNqtdMBSSYZ83JSeRoYwLl+Q54gCINdF1Rk/O/p7L
33j1JiCS8zB7SROSLbQ+fFY62oa8sSzC0AgeGmYondhxEOUnM9ZVJHQi5kcsSWMw
CPz/mnXgO7JWzhCso8pXOaquE7o72PUWULmP6ynnmmHeXPaYXtZ+67eIU5+6pwEB
AbzLIIFQKV220TuhvF2ofMmjm6vpWV2thFqEqaqfj7Jlh5HUZAisku3MSMItKPwv
aA8LbnLD+ysPYL1KDwEW3sXVy6TURaxqNOSeulalhQiE8hhTbOUDprS9BISMB3uI
jgQgaJP3dOe3buH8m9+H10+V4tPmX+9RmgS+QNbupIhXSq4MN5u4r2kJlc7q9SX/
XPf1LTKWxbmrKNCVmmyc4epJNenryFChvqit9OurvyZyGtO8zynYZzTW+lwiYkcP
sAgTldVQA3q1zbu+ql21/iRXIDrIwpZnJ2Hgo+rlLrJFFJ38HBftAxFZ6bk9JsJx
YDRAOp4nIR0ww/NKqL7Gr5/9f69X0rQEOoJc23xe4izuWiLny/Y6tjkJwJ+F7soL
SHjU+9raYNNPrdr+lUKj2STgFxBRyikNAaqn8eOv1W+KaIYRO0+4WQs3R4BzTa9c
uhfmD0/nYDAYFwXf8KGiimHjvxQH5d1jNoys594CeVZ2dZur+oQUKy1zTTb2WNo1
0+vf+gGNtplkeHEAVDq74loRNFLou7kcSat4sQoiOBSUcIwlKC/dT88mV9rRuBEf
q8GtvOQ2/6dDKk2c2xe3Oy0gVJoy7wzNpWUSx23lW9z9voUx7hzwlqESMzapdaGt
cnlaIUJpJw7O8ehv4K/DWnBgNZ2Kn5pAi4KY9haGsMGEPPXB/zxo0unQwAw0ewRM
nDyyoLXLS1qoRxfZNt1owp7iqtwJ6Oob5g6SyydP2+5Hfo/R96P4WOrgbqcxGHV+
5+exe7COhe8LZhzc2RvCaYxeUUnB3lUwX8s2doH+0ZUtrSX1qV7OnnRCBiLqToDI
DWNdkaleAPSzZV1bJnK5AHOJzEGG6PkkeiXALaco+DQMa2mvGBOheWoxOVnuerAM
uXgfq61h7hA/MS3ZGTh3QRUvQP3wfVnu+WA6kla84EUf2HUtI06+Sdz9v0Ppwz5V
OGsmBqeydDgSRHm7OdGo0k/4udxyaQwsH/puwjwbOfechSsANN39XBtt5CBDt2dT
dBQsoXp5f11aMWFuMjMu6RtioHm0RT2KkfFfbzzboIuI0DoJOS9ydT85w1zUoKiS
9FkyqLb4BFebTWAoKuNdWNWddflT4uN4N+HU6IaI2JDIULW3JL3kzQy8kntnBpNT
gp3FeVb8Mj58MFFQPaNQaTQlAF9M/NiyjWcdbD0NDVJqim7vggwkVBkB7Q1ebUdG
MGd7CdlhvafsZVKEVeeZgAqX8y0WlmFGAIaZrJ2zKJ4I9IXPPfu9KhnsaXM/diqJ
cOsMOB1bWF+TgU7wEmhapJXDsVAAFL2Ft2AGQw/Xy9TNGRAVud/wYMRehxus7paN
GaMv17RtvNH2szmJs0FVONLtT0/7Dk9iLEcp/Sr60B4/GtpUGiqbCPaJVyJd8Pty
VtL4guygANPiO/PHXhaPK0U/DbgUvXTrrYNjawfNl1yeRU/EdiPQ0fEWiUMtciyl
VfvGj7Mu0eUwWUgTJeXMQ0qjek7WPWPfYNp7qADYX2UxqmW/o8ipo4uKRlgMMuMS
GFcZ/DW5/okXpsKSJhGFocJ0CY2vcGDjqyz4QvVkXoAk1Rgck7EMFAAJHVLrPwGD
r0jQBS5hxmqsQrJboimhxIAJRFylzr2CMOkpZl5FXVeGx3DUE5H09Qr8VdjBWMFx
NzNCe2LkRZMVFHpkecAbT/PXIXyB4AcubUvf2FRXh6oT3275ZQdj+RUI/ts+Czlk
uQyEXBwEJsbU5fP0vma8E9hJ3doZecgU+jNihKU9KgclMBboyMbirRB/a8JIauzy
UmJ40qGoObiSPCB1FAUq6S0QBA2RHHPHOiXfBUjOL4cKILtphvjphgJITi8UTnSI
mmCy3X8Hs+wpcEZECNwr/7ZUzyuMnj6WsYXIe8yUXeREj6rvrTfES/L7YdRDkeMh
DrLg/gKKdI4IJ4DU+2I+MpW5BqJ5kqvq6bvu0IBzZcXJqtGw1PifsRoxQVK2t/V8
b8IO8bpjG7xd64s0zt4DpcqR7CfXvnJ07p56LOdOxnLsy2PQkdOS1ppV4Pg3WS6s
/T31zDbrk4xq+NFLxTjy+KYNKtW6H9/dOLCloIyPR8BmHMkmrNPEMPiKAh73uHNt
Gj/VZLP4oZ66lrKEH0DxL1aZBklUnMNetJGje4gqPJ55kjjuzXbpcSgf0bP9EVNW
SBv3OBXpx5Y2B/i51DDunlreMBXnH6x/MbtfQgLvZel3PhqXnZ6J1ch+jSFb/ZO2
XHFg/gmGVv8DqO3PCPketlRdCSffalCwCGpbqsYjCvCCmLqyXx/JeKC8eTW3zR7j
s6+JZn7Vxxyztpoa6417tJsvFKDKm1dTEDR1ZbpbyflGWkMCZD5xuLyNI5JPNgxg
RGainKFoinEQL1EFLAB+BuTHzl98EWGx1441an5Y0ckXfgtyQKNEY9O5zOLeLdPH
Alcwsp5q7Y3yEgR0rhtxoR65a6IaVHepvgl4CQqygeTALdsbkrpIKZ7bYoxnjy6A
CBfdjdXbbcEhCL59P0ZdP8rHsdtWAqWkEGIk5G6T3Z2EfldVhZ/TLPpa67DgVseL
La4HrxNf7ULmSyh0AAEC4TI1XihEKv5GTTUveAJ0+GPF9WL7rNe3Q3GNTdc49IRC
C+tt3iMOPCB0URNjnEzuRBgMSD0rzZgnTulsidPlARJMqCRzl8l6KnayH59YBRwh
E5FQOQWC7k1Q55Xi+fNdZbOh9LEE1qiDl5VbkihCdD1VIDg90LDkaRBqNPSwE6Yt
NTwO+S1maevZf3pz7WsKUrcJrRdWHvq7xsqFMjyKow7aWFfL4X5IHKKpHlJTMJoQ
PdAODO8pl4jog006GsVqVcJz6FAR1fET05VKiqIPFMvsBcPYb2Qaxtb9XImONnDb
Ie5FsDmqU6FU1OjyQdukqQy8+GojHUf/lsB4GMrsI7Tj+I/eFZf8J/eTUgljjRhS
IH1+Ae7WSTnBNYoyQcJ4d+kH2mKfedArPgnkIlpALaddxo7sDvsVxmVPtyJn/OCR
z1xhxyQAQ1OHqvWtYtvOn2FJbeaZI8U6+Miqq/M2jHU4xQpJ3BO3w20Ti6/7aN27
8reyxUSKcHxQTSjYHdta4WbpAkyfkU7oN+Ijgvy4t+owI5SpMhMKqRDNQ6lnbLIq
wL/ps2vdJD0Bi45d5ay9ltB1uD687zhiWK2OjxsBJaHJwjRyJLSiY3RPxM1QVJi6
rkrLQS9Il7M7Dmja44yxqCtunIC0ScmEIEp7rREw1GqWZBLn19glFVthA4dAfHdb
lWtaRP2lG7yWW8OqjA1shTDNLprkVLPhY7QG4pkpZVGLd0hX12F8H2/4303DH7DQ
FCPuGri6o9wsL4eGiGBBenwU7JJZr0IziJ0nLlVgtadofUx3qhrBl3Q048VgQ8zO
eSLVxtS8nCNklbSK8qHPfozR71g9ucqvAkgY/utNfil5YCSgufETJXaZxv/Sx0HK
Cw9GTYM2sxZx8h5thpyAl165WVn0+hbluFEyRO7z6ZjULOrUhErAMII8jpWl5l1q
eJZx/wJTMBgQ0oTDKbF1A9eYQjqzJ1BYekP+pS+ofa5rTtWGaVPEH4tKXjnNlDH7
2QbPc6ZdIt1sJDjRr7EU00p17ZdMMEJWSk37MtIUDhDR5DW0rWQ0BvGtVEkpezqT
P3vTZFDlGGT5jqwdq17utqNHW1x87+3egm8cnkH9sEi4jr5jyfiqmudLVX7fbimx
WjmbOIXViZS/iMUPggkXVdllWUxxsLrL1PuQTRI6P6+VuBFj/p0PRyB/GHYYgvIg
DuPLhcJ96uoxxjKrOVzwW/E6kueEcIu8QmqQJGJHE72fj4BNuTLYXlhpk5ib5uFb
X8ZfglV9uM6Hf+SpSDDZ2sxhMtE2SZC22TKSVFLU0cvVH7ZFld22qVEITaFL0LtN
kKTV+cgdU7RkbeQXW8Lu3Ke/ftSn2512iqWoBHKgrWRm4iAqMGsMtfx/zDt/XoGs
/d6a/pPbtNCLrgZPmGxJb7NgbKqen4g/idDmu0EZlamVCKnua7tgi9y31sLWQ8hV
DNA84LqHqz4b8MqKoXiLJKzt/TG0kcGuzbSmHmg+4oE90Zwu7kdLVV5+9oo7Tzui
61LvhijlvbdWCjRYOQkmDPBEjXhK9QlMGo2MRzSrkBW9Qny74HE4qcfcZOHhMR2R
diCuwAR+m+ZN7qWaFC69XRNS+JxtjWoYZl5wnRo6d4c6gcUd8h1SbRrB+rWopNrb
ZHdpSrtGQCANIYENpyARp0PumZhWXeFGCXsrvY8uBR1amekN6PBs11f8Q9YikJ/Q
0tNO5NYNj4ZryksU/8TBj6uBV9A2PdAzlfUnFrN7FPfgOo15zhK5RmSr9bd9BET6
9wRWkRjX2zZxRttPewdTURHo01jwMtmZT0er6d34sB0WjRMf6HSYBbDWKRUc1pXR
IpXUk3uoH229i7pQiEZ+Sj39amVtQOj6JlwB2gfijqkZJCJ8RP0mx8hk18gKG0Vz
Y7KVz48neFr+K5rwDlqxMeRZx0jLZrwBhD1cry3/68ODkCqEqZGNxtbNYB3+BBil
HRvgQuCFDJ8CFuIHV4AWRVZOi+KuZESDmA4t8rCPLUnNQzJw13OrIQyWr++k/hfh
Y8gQWbxX1lvKRU9U93oDT7Dy2Ryk6GxROwfL0klfRGX3Lqu/1xSS1sr9wgATfHjH
yZlFgqqKkDqWQ1qe2D4wT69zgRghIFU575csHhgEhIbqKDBlZZVAfNA/VT4RrtMW
sS4ZxmpMXJNViRAtj7Ulzn4eauGhd8g9SGa0cX9JMvs+TeME6+64ySPLigOwmDV8
DLeYbpECZQnB/rhoGSu2I51yQhF7J43M1BOJ8CSkOnBkMk7j1uRcmQO34B1Qb4mJ
HJb8NLXdlPyxZbvYOS+MnZUSNMQ9R2BEumGkXKqzbv7LRAfeeDGWmjVCcgDsowrz
GnHVD7+SiXXpXeL9JF/+NYK1ZEPZw0PncOmi5oeYPO/1PUEI2LfIlbul7KKUacdG
FOjmjTsocgvxdzXU6Y6rAH3W/mzU2UZNROQ4Q15sBY0dLWn089fwqLwBQw/V/T9x
wi+3L76nOYy8oMCqbUX5XnxmZlir/alUqTqJ9ERg1N6r/uHbSglBFn8g2ROKsa+x
C/Jq/dkTyGNJeqZ0C/SHfOIMEAqUIJzDWhJtU21h/mV5JEUJdsse4aAm+JdflIsb
v6izaErmouJQCOuTYqSgEmDuy06syr0JGPjb94EkoYYvk68l6SduVZnX9ObXpt6A
tFLP31e1Whax1+2uqrkOFsvBHMLhBfDKbBAnbwH6Wi1vjrXB7CBsan96iH1saxSw
PcSDzixCW00pqUY72g8Aykm5+3MOtVmqrWpbWcs5tmPZf6affEid8OlagqGdM5dL
X7qnA1VitSXqyjmzF7cG02k6bBsWmlCeieVjo6CmzH7SK0kc1wbcQEtgF132Yaw8
AMb19WcX32RTULR15l59ugPvvNKbt7ZMjbDMOP2KW5VV+WjAshOHi6gRi8puEeS6
GxIOSy3l8v3q4nlU7XaH91uZaQP55gViwzwzeeos6g9A9g2M9JtKlu4W5AwC047C
H66kuhygK/4nW0x6fF9QrzLmyBb0Gm2rFsBTLgFHdGnc5G2zDFWnz/5tZa15H4G4
QjTgS4sXeF1k59Y/9dTOwMaSF01bOroOXWE2m5q8BWI3HWDJLBszEJfaCjgB9OKF
FUcHEI1Jkb0Mh8/NvmXhoqThXVnQMgsv1StDi073JrUf18QS3JSD86bBQQtPt1yz
puApVKDUIE4sszJO7DMh3dFY+xTis/+r2wIhRzrf3wEdEpjoUkJncv9E+IUcvUdw
8A36shlF8EQotIMUFG+55BcIDwQ07badLKypnGMwx1l6kKpZhC8RUi+CDPLfpY3u
oaiwVz6hDF5N/BguOr+tM/iZHyJI97LSrxLxFbm49YL6e2D7AY/8DqxECcxu3FVT
VJ0UApr9QEphMH6qmqARhyBV3Ooj95zk+3KWfENpsGKHLTMuCL4DPbVivOH9Gf9x
jcFspC2yxAOX03iqA2yE912tHoVEBVGm18CL/ZSa1FhAM4qLJxjZpQVdihEACviY
eofKH6wizUeV1rBd28unx8q8M03UQXadOKHn7AHiuePTwA5Z5PMLjPtxNbiytYeP
utrj+e3KIf7XJbtNjAb4A6qbhtQFovrw7Dz2qlh39yn7xJcb5Lai3Hse3ht7SU6w
2VNUeKmFHOBO72z0SgGVmsEkm2xRc1bj0GwOnSu9BpiT4482d7PLZ36VEvKHpXog
cYYg+zSdbkKW3iXOyl+euEQ17gA8XGw0ortzTC4+wNIxfk75KS4Jra/hiWzY1ijV
i4mjmLdHN9UPCqCo39UGLqoaGqscwnyGz94/HPJhXFxt4+uXQCVtKpr262oYrxdG
rkQKLBZB4Bt/Frv8flaCXh+Q6f25MALhUsn/KsDQwNl1RnVLEWLKaIPh/hypd6As
r2lRnRO8wj4aMVKINiKnfFJiSeHQcdv0ZNnKfmT5UTK+2pTUkRbJUslWshYA8vWa
mXdrQbqHYbJFAJLSDhn7eGHAY7Ha6gjHcSDRg/pXXf2WLo43DrN6L1rmQ2yzxb4C
+pJHUcPwrR9cKuodxyw1dk/ogJyfH6gW8RlEUg5uxyNWfaB3gFAHipj9bITD4LO6
UBsLGq+4JynQjVxgZNpob05N0gfHv2t7NrBYzajpo3LhIVTR2ktAM/ClsGV/SeZc
cQSCMTOWd40mRLjzjtGzt/ID4pZ3qbTaAnpRZtiHFImb5NNcPlZS1jy9t7N7IPJY
QjhET+EkoDOiqCs0CSbAgxPCzDFC6sTXCaWpQqzNfUbG0XAeXitFWqAI5S/RsRV8
JQV/N1jqOZpQmKl02B3dFCEWaVWgVCGAozScptqPCEenST2rE+ffTLsvTxDk2Ctf
8t0o4yh21wl+OouR8YBoLkAeEE1nRXMZtLojEl/k4BYDjtPQRstOWLGShRW7KYW/
fdykr2iju1amOVsrS5MiBp8G8KItCitxMio9Xc1aVfAIrzp6T8+2K0o9GN7vp3/s
3CsWdi3v5wCgpfls0A3GWZimetUxIrm9B9j3ZytVjHrq8QccG2Sw9H1i3syyWw99
CD0tz2NY/5kc+glQESVNv/GabwCi3Ih3Nb/QtanJTwoHFKIAtMuh82i51efrVmJ7
upGD7vEqZuIJ/0PbdFUb7HoXs4y5PIHCiysnr+5zaj86auGl9g17Lh9+XjFl9oZn
p7TOLN86rMotkGW3j0qsQ9BBwyVd5uTgOKOV1f4iUTcWVhzViU2yr9Fw1oOwwrVU
ZGFviQYIIvE0Ce+wizeEcW80OX/0Cqltk5y+enWHExU+DqfSy8jwT8KohGkjBpSg
KunKWSZtrMR2LTdnme1WNtzi2szIt5bfwFVUL9cjynZ1rDcuMwQMzvEd8rVPqCM1
DAJpSu8x5zHT3ZxEJ4lFmCDXtmwR55qePC2RvLwts67D16QkqsfWM7tt2znb/fAD
taOx41Ild7YmRW5CNChbL2xoKkmLFaVW7q/m5Hc5vL5HA3sWxVa0C8JFufdtzxqW
xdOouH2pPV63tkLvjXMgb7WZVqFcl+MuOcD7hyDTQSI+/Qii7593KrQnntX0vAJL
fjRxRt13WI9VFY1L+yp38rRGciYBOdpRBfHw3uf6yQlsThUhoSrjsUEIoVx6nJ5s
OEa/MjLEKsthdaos8cC+pWOfu1vyMujTP+iQuQwZ2mrtEkdX4UzMXPK24JMFpWpe
W5OmHwjksP2WVXzjpIZtTjmxMHuKtBMcSPxXp7P6UBzqsiBh5UKcxGjnyB/8Lt65
sKd3XWScbI3vFB44VJAJj+nR9SPKs3QFuDIGuupyhPg/HyO6yTVHTSDDf0Slg3Jd
AbprPSu+dRE5xWHeHFNRhCh6PHOVQYc5tWhdl+OAj/TqpBxXaQADb0gKSMlJEvoL
er4W873lOr7mtJ7584ao/Ghp6bYPsM5mmvXPK6/hpJ0hI31Id78y2JMkgNIq9Dv3
RofK7QUu4pBJNhgT0W60ljEffvevEO1KMKM/p6Kf6zAYlg+6JAp2Zzcrl595QpCN
S2HZt7VtrcnN1ST8G7n04BG3X+yb/p+kXSfaDFwwK/NIH7BRB/TdkyAEEuV1W3h1
6ggl7swwRgdiDX2vXku0e6NnYxdSXeUl2drdGK6WltcvlpP9GhUKHHvfyCqbQHLe
2FxxcfgPT4rHVIZFQ4hSsh+TO0HGjytOuLfRDGEraOk2/POWIebolTe57BeXfei0
2XjMneGYEZA4i92FaFlAEwM9kbdj2wZK4nCacg32z7OnpxFo5sKpZq3a534i+Ofh
3/OAbh+LM/SzO5Z+wbUe00MGHD26D8AuHdWdPz0VDQ8pyCUzEgBEI+G/GEBz9NmQ
auSSrpS2sh4rt7dmAzXYxRphPSzB3MObByTrkmr20sepOWLv64ta41OFj/6pJGH3
T2w39OJAlDXg5oy6pwxkcPso8iMNicdl9RpWfVT2gJfV53QvLO8zN+2wQsPdAmJR
D/YpsE9500W0MWL/59nMP/2Ha04jMrWloWExIITAJatNSX8GOYdBvGsg5yjwL3a+
xs90jOMlCucEym47TjdEz9eFxtB63ePWhk69mz4L+uX8olxzTofrHVXzbEJzgfj1
SjbVx5HbaLAJ9jpSTLARoxdUz3HlzMmv7j8ps9tDBZ2i/fnL47JfP0+Lz8WsgVld
mUnP3QFxuBsZD1lRew/6oLhUJelVBLggeviTadZFt2WeKAXCiSSlx7dZLz8ghFCJ
Eic1CWug2w5UYRbknbSXeOLivFFDdsHINiyIP+vIcRaHUqbR9nJxfWQqtHXxWvsS
rt594OBsfxik6UrUNerrjcIeruJZlOeUOoNGExK++Og6txCQTaCISstV8N/KIAYd
IN0wKqpNrQPfqWkDaKhcYiG9TKOMNmuPaKhdCYmdM3FT9ZxMYqrP3vHtlFUeDdYa
bneO0CM7zTfI1wwoNS8gakq4RGoCmHAIQsBMV2SQ5RR9eBD41Kn/ypTwvBcHAkFk
R9SFjswDhn6dtq2c0LbD2b0U2eDg48G7sYG6TgukrecUJ4sO354HKDwYaYn2r+cO
GvMrfGjWMF2R1zPTF9I+CfneLqDWX+NzOLdF+vv2jkBdKN3yklU/D2/rM2rbL4qT
7PYIJLWh9eGjnTXcZAIFD7jvALI6JcwKPK9rv4nYe4GRsgwQMIiIJdzbaTwjuRI2
luH5tUrbkGzowjhOKIK1lcQpU/JIwntpvXjRJ4+UHeGMCyVzETiUOsAhZXQ+SrXJ
VyGNnIWt7gcKMAJEQg2dWTWFLjwD0Py70cAWQJnXmfdX7M42gHbV/2l+JzMepaoI
QQ8xNZ5LWQ8YkDfb+aBfHSRHUtzCmV8+6l4akhZEONufwOJCeK1Az55X1yFWfgGY
Da/R6xd+VAc4NdiJ/r93TFR6kmexr/41tAfsUIJhsZjQuAOUv/xnXNLH12Qf51ch
Wmg4hSjaplexpm2AUkJaF/sL+ntNCSFL5UTE656Q5zTzR6BUJ8CEJcyq8fzUzEoO
mHnxLwpiflVu60P9mUQ5MhVe9smqHcpW2sb0OQ8xZHk0bXaFpKkVkw9d4U9esANY
J/0ycC6okF+5PfMljXEda8XAeo8Tns/FvI6PA7j9GV4eFkfFFvFTaxfy+UxAKkcv
X38YQQQ+3j7R/EJCNQKrJiBOhbria3csfdaCBEI9+bmRrcjz7ntkxAGtm9ZpYlzu
ipBdQu6u/IHzJgZM8R5Mz/3S/094HRhxnudDJLa4NHCvbDVeV/Pb08cEU9Uj5kLo
87u/Dq7WyybPWND7UpIbAI7CGV8kTXWrcuU3HjtA/zc80Kha2OUhuiSdwx0UPVDD
rEAcbg7l8jc+10WA1JMOk6dJ+WrkSkMmfjCUf+MupBsraHaQZ0BY5RSQ/dhpEIFQ
ZZfISxkjg35CRPwVktP2eY7tvOJw7XK5Fh7KJaVXGoOugT68Lbmf6nu29L+jTrJj
HSgVrHL9vuNJj9aLDpE5NQCkQZR7/YAKT3KLFdM0DJUdPK8fF6e9hyPw6TuHbW3l
qiiA6GK5erIi7PLXnAFy41h0NWpWKRZuQTn+3qhJxTPRC4swUifO2ndBPhFjnNv2
C5/c3zhRTuwbMiCPzL+imIYrX5YybiyZrV5zfAVYawOma/4ENWw+lpLilZVu27HN
sZyzWPf7rTE3gaxAW4GeLUC9Wi8scMe1v6M9yvWFtAiW1IAs3AR18KyKKMjj400o
ckJo0IYQdc6micmE5Vi0KJuGkYORzyZrBRbi5HVQcJ+HyZDbcrJS3rk/2Z16+fJF
SzaoSroM87zbHC4Kq9CkSZw68UbokvPzs3p0WpW1YhW7HQR97gPb7qN0XlC4AyyZ
uJKQknWFfROQR5SALNT6S/FH3oD/7H+jyLjhAaj7MwKwDEwytC5Nw3ZD5asJ68Bg
Ne/OUAZPparGc42ZoAdD39im255Misb0vX2RUUdEjwwllCfb2r9324MWqyS9s7ZV
Nzb0gJWUIitv7Qko7kT0DPPoCqe0xub3DftYNKiWNOx6uxgyA5XuEjP9LhX6jqTo
zjMPwzeFp7mekBoJHLbx33B9u1MxhYOxF/14zXziL3aCOoC/ZKeXC4WMaAeY57bI
95J0uor1jO5vPeco7JtAIJRRTos6QaFT4tv4+klrM+CJD4DZKQBxW1bhNmFpj7iW
1eGXV3QNJsDIek+vibWEaYfYiv6vlHgEkK7RZtS1+/7XP50qFMXZirij6Zj+NMiq
IX3BqwSiVq2oArvNLxcCFkbDaMv+RFd6EphD9MBdlj8wfkPbT/sdLz8x2J3dfZIV
Xqlb9+qUxR85Q7Y0BYXdP9c6CE1ac1ujt+6zGfc1QihQPjlQRDakaOtrUbFt/yvt
wXYoNQYn020FTzdyo9k8qc21OT4ST8oQ0sCDQxQdt9ifYQbb4gjjq3LUy5xtHCCq
eNekQGsww1kGxQmjIBArznXnjDHV9ILBqTRWkp4lnaw4Cj73cgcmisvzt3eFMaBi
A0zwKfDyUFsIKDAvAuaOAozZ+NBuLA312x6661AeE0s2cr8haJyOSEyQ7K6hO7ag
odeFeSr0FuAcKqtiL4M2oEM1ASlspi9JP+0ncH8B+qNKQf/za9WnjxG0oZMb/H7m
RVGBCwBA8SpXEjkt3CRF2ZXO25ACbRJ+DINPN9OUUjwLHyP0DRwno+JgBz+dE4gu
b2et+m5nbMYp36HjmkpQ2nb8BNJbKEQNLbl8mV5I0/htTOFmlIqDlOU7GGb+Fpmp
p3dbpI2sASsREponuiPqi0zuRW2/bf0lRdQWS03AX82f3IaaW8g+9Wnb8ihYW4FV
j9Ad11fbNs39CvMR0BIWIhrnQESi0zLOMlwGoSsU/snRN3N9kcI6uXc8Y6gmsXHR
8oM7IRDydSezFpDYi6srdszx4YF8dgmrPPC/VFW2ar4YGaCaS7U3aAKPPOJPGWKm
CDQMDuh1SEA7/1PyFaBlf6He9B5tqLPVZVFqS8SEuggN/MMCSzlF1A5wJ72Y8++i
rsotqyK1ej33vyQDeqyEIWiF1xn8K/eqqdcrUmjxrla/UTRli0eHULzJcBr/bGSa
Ejm4wU5LEqOIYO8fTewqadezWeniC5WxQx+sWbA1RaVV1p11Lk6xRDQK2KPfqKWj
lVxuoaWUrt3wfGOTCrC6cfzZsigH+Er7mxovLu9c674VjAYa7EQWiHJ7xMuLwNsb
mo3isugI3rKoG0u258S65JSa69ZBucqCCne13AAoXW1DefijS1WDyMrk80A7IZEH
R06ScB0TfmM/8BMf96uM13ZsQYonSxsBIJo1kK3B7yTikfhBvIR6/Mrh44C7KsAs
bHBRhBOJMj94bkSKozwtbi0FGxtANSMEBo0JgQJbsdnQc0OlO7TUtYH/GxXDUYeJ
tTN9w4jEtEU5eG2+tO1Ho8bevFvwPW/AGZmQnlZ/DJqqxMdS0stRNKXoRzv+ppZq
mf91d8gAYZNui4SSF7S97+5cKpKtiC8PHJBhIKyG8RfflJEe0T2P8M6JdnEx9DuW
Mo8cugLKv+7hI/LS7gJqh8oQvMTkjRDLG+QsKC964s/336YR7awT6yXPFsvsxH24
K5XzxGB/fnKXDIioIJvBrN4OvO11cmz//b5QXcz5KOpwnmYMj8VoRahT0iE2uSuG
Jk0SezDKvnXZYA0MAAU6u1Yn84cUwbgPXDN6w3lXEvoL6XRFHEbspOnC1pIUqc0U
hvW+2R0lBQLtp4lEOY5K3Bit+jj4hirEcpEUUNX8kAcR7zS3XXjhCHsk4V2XLxgx
h7HmCKuQE3gOtJiqiYDuzOdC16QmEzdIu+aZxumQpXJ3pgsvmlxcqkPh+4aALBZg
BPNN/39lYph6EHpzwiF6BN4Pa9GYggMYeu1nZqyTNUr0RGzHBINhL27YS78BUczI
Cvi5h7RAIDJsFYJPyjPfK4D4OYuqhAi5iCZu4Bc2Qfp++uxTaAAvXQ4afko4IuEy
7PRj7lOvZuAHuvQeYMACir9t3D1t4aGsvNvUy5niXDr7Iga2GO6UleinYXQDr8b+
4mgl5/DwnwyXwkx2Ld5bc4ySU1w/4Pxe7SQYk5t+IdYG3sa1A1ZjjaoXriD08TfT
ccJE6DjqcPYw7ZT0I3xCj09+1+5CbzP56ctq7tn/8v5GHOfc4IlmXFHrJ1jYp5Zd
j5eIYO5DY5ZJ/HsCRpMLC7cSRKY8UCCA5xGSmhIO4VknJbOECbnpLkElmFMMBTuK
167HcLE9av5QxU3gkTr9NMhN6rgMK4lta/pDug9JVVPye4v1Hh0D/IDaZHPfpK+h
oJg2WeEPR2AjH7+dAY7sMxxRDSUY2vGav4NmPMd0IAe9c5Fq2Hjw2yQcdKQ4GwWu
ZwDqCv3SbiapPfaC66IB/SIUk/8C2uycrNIA82YckLuSWgOCixy/lGPiEt5w8sQJ
sDR6jV9u+s0i3hCIDA6BaG6qUbgCk3MqByWsys+n1Avh+NLavO3/SezeEzED4Ftg
c5prkHtuC1mqyjIBL1mtK0X6sXqUVYEJwdsIbDqeayNc/IIzJFkDzZWI0HstNJWe
TkYafxVzy5ZakzPGNomoxHOZxLUCaVWqfM/Y41yPGconKtyAr/dTpFNpzDn5M0l0
XM8Hy1T14yeonugi7sgQl04xh/brW+QBWJ3AFj6A710pLG+U/AANPaRUba59FRec
96kzyvCXAYt/vLGDqq+ZzODjKzc5i1o6/+x19j4wkArS8kze7GlRyWHabGPl9kdh
UfRNq6akDB8sPo4bWHGtCItr81J7D5w8u8NQZZBMpgpe8CjdWzZe5dfv8dRcupKO
9sz2cDaGNrMSJRFI9eGUDAZktFIbL9ZVLUDV4gRw+WI/6gMUbTvadCIRxaSVIZp8
9kexYlFA4yd9ibRMeoC8hcF3C6AtoOtSIebwYLDLYNwSiUcND7ImFplMIktomApW
u+e+s1wg5RuJd2szfbmiqt6ooaAltgs4D8SoA+bzKwqFZvoZ5YYgjykl0owg6/EX
h1W5k36LksByn6m0OnSVnT3A1p09g7BQKALc1WL6N0iS2N5psgBPgSMY3DgGrw+u
+HKk818L9NjfeIYx/QfWME/yyH49pr4k1wnqTO/nVuRjrXM4WRGkV+VHqPTTzEu1
w/9IuFr9xDb0tTqX+CiMgQr+d9uX3p+MnwsBIBG6nBEyBzTd/RYegRY+qjADVEOy
Vr1sjY+2TbfbC9ZPRv1EPuDNUB9lKW1mtszTO1E/Kd9SypvD23PylyeY9C9RuPdD
tF6deMVYovkJIGrXpGvdsFgLUJ14LrV1Wk6tQVVtMNEhNWSCGVw0SwYlPrFc6Kj2
vB933QgJCLbtZzZDBm42CvruTYJMPbp5zS7OWTv2zru8QlJv1Piqqd6flW6BVpfs
xu5ZGWcsuLRHZIoUGtpkT0dr1KIPliM0LE9HiUX6jXR1Vx4jAJ0NMM25h7Q+uZrc
1+0eo3Derrul7jrjANX/JdaXaJCdTwsIFQVVwWi38j/SIVNkAinu8Gu9SIguPpn+
X4tRp3aA3pvckkscPNeZBhZs7pgPYKoCy3HCRTj1R1P3MDlom+pZV4BJklFzh/At
ldpQNnhoEePHtf/kz55qzmT4rGlNwY5LonERNGRSkJiyrvlJsB1UKrF09pM9CbNl
qM/acZH89bUcrbyxoW0HGEqgNvOVN1neRFPi0FoSH21MrO5g/a3cIlEHHygHHcnP
Et9vR/ATAcyKnivsFngVOnfPT0+eeIeuUWLK5Ne1IyFN8MfNGpxTJ2JS0qZrn+yL
O6fV1RipdguG6pkzCbW82bu2ADCCxaI5U+3MtpQn9z30+GWNMsmy6AqZjYFLTApn
FFhrXVGfGNpMylrNfR3yg6XTIRL9L6qhtVA9daLi9sttCU9zstCEsWYIrKb+qSYd
DK5VZiqtVpBIAe1BS+baRHxJFn7DEpXA/NEFw+Yd9qCFUGdOk6bpnvjsdZUI6UeZ
5Geyy2eVs2w+78hucXyphp+ffIkSPO320gS6w/HgB78zVjog0RU9Csrv3M+eG+um
gAAg8KPs/98U3criOEgP+FvYTuZ28h5hqwTbDAKok1jmUys6JPxruA3QXKQzKD01
EMJhTWF64vnwbaPfEPMwZ95i5TAxxm/Vpw7CgrmqzNPnk3fZxHDjBqbYJNQCO6JO
o6x8/CyAnyI71ayIQQpQC/fWlAbfz9++/W3JfQT/JvcDwGmSsgISFP02GQNiMXUG
SMF8l/fZZnoSj+DiI2giCrMHAL48GQ6axNxu5/Sna3pBxKG5eQyp6UV6MoYtQxyU
Rhz8gizrkSCt7qa/fRkTzi5xAehOw0uu4mYiqr4mcnI+l7WalJwusL9Yz8gGnoXB
bz8Wj8M6QQUKh4/i2EKiMTxibtY79ZZFaDi/ALVBcRl13CNMTAdEeTECTBIiva5c
GEJdRa4FRuNHGOdXs0TCGrz53xT2ulGs529eORbM+P+a+l3yExKX7htHLbanzj8I
4rCgw621riEPHNRX/yEuVyWmXTiRXO4QU+DaawCPd2ouOlAq1lsB+yQJwtX1kRSO
SLuUCcP5+0VM4WDCKQ0OMe5Ir/hO+d/uRpd330BUVv/TtBRh5YX/OnOGoSndyXLS
QOWSCc/+x0Nbw/C6Ey2m+ZbSFIhEU+D+U/fBn82VlVs+XNL5DD1yrh+nZ3r198ol
1ghcZlRVIOtWbPjuBP4IuZ0DVHif+cxMXa90s3Cz6wTmm7idV0GkkhJKRdzbVu7z
oF76HZsfCcLrKZUZgFrGnGDLZBtJtXF9sVIhGGEoFMl1BYYxgkcKltCNmOM6JDJR
vg0nzY+Tkd2Ovd1YR997y0pbGRBsjz5JzJvbKOUtGMVY5QgDd3UHOFwONke0q2C9
4hQGKP71sjBXsCdVB0flK7V/r/6jF04Fo7o3MXuKPmPoIJnKBGTnSdQwtm1SlVyl
XJB1xvJ/OhMEirXtr+V/IumZ2wH9Got8EYL7xRfeHA4mCXrplBy3taspuh/HLaEh
g3Uvg4b3lGYIBKOFHNb6NxH2lgBrqhbBvrmoTc51E5CTKBq+T/IVXQjGqwq2kUaR
PJG+jysFsAlgbXa4NwDJsgofQbty46WOH6b0G8rZipCU9PzCNn6Zjov1F13XYJzN
nv+BnCGZJwy1PEzWzvRD1uoU9h2vp4jYbPsnMCsyj/Yq3w2Kg8Ko2vZVsdpEr+7v
4HL+z+EZUSUjRX8uSVAtSIn+U8Dr1QyzLQwVxlCWOC/Cmj4Z+yQOaCzazKCuwxuq
DB7gOy41qyu20HYRFhmgI6dihqQ64xgtT08v0CZZUviMW+SXyDvcDTIpPPU+/bRZ
9+XpaXBbl+RO4qxSuMPWxaN+28PQG3rOEt7KVUnj2lQ9gSbzkbEilPhiGUQfCfqu
QpSWjgMsDU8tShYA3RPd/yJidHwBYojp02yeoWc9uiq0RI34N7DG0jFBnwvdB7aJ
DF4oW9rtCXmvCAJ2DroLupwfbx5CmNVJkuQ4kdf22cja7a7cPIjxKu0FkDJJBFzU
S1R7d6W3ayjofBjhbMP948FxiwOGeOjxYN9risVr0cIwzN5VW4JxnMhLWCI+ajuU
TtL9VxVKkTVAZXVZZQsxQC9BqeT0l8ywrzamd4ybtNMrMCETFqocTsdEQtqN0Lxj
lR/eXeTMRF78H9folbBKzmDaNtwGaP95ZspT3EyJDg0UZfdSr5DHkl6DBVJjykbU
HXHIg3hiQ9OvcrCjwNoM6wV0Lz7vQdVk83KEBYA4N44ZNp6UoPnOWJnBsjEpCBEd
8ftftuGF/gYsuou4kRYGfK6IPCZhlE2kPPw0BkpATylkfnz4hZx+sQbUw7Z8FXVP
z7vNQc/UJlDAuz0vGOxem1ZnUxGomivItiM3dObjrfhGbtILsydc9cL/JKBF4h7l
fXVaq9H1MXFP9SHfUZATxKPp3RluZc4fZ6W+1SQz0Vg8CMwmKIxo1GsdpDadcln8
jC5BDczUbqkTPx/jHbyzqRk1KJH2z6dLjnFs4SioKxKXTM30tsJt0nfOckTs3us1
iKbINgRCtlwSzZFptru/+p2y2Rsripr6VB0Gw/YsMeyTRXk1/KH9VHnXhamAjFtT
jsB0ylY9BWRRIq4mSdpkdxjeMv7i+vue15cSgYs3RhmyTVrJnEPvq20SjhZc3SnV
irKF5ugOWQjUIcrpmwxK6TObEoqKikBwsEbXOVkXv/F7VvVshvz2T4l3SYkuMs9O
VXeS3oTVEEm35XLZKDE+vUJ0FD/h1CBWKOMSOjibnK2NfH7//2sqrZTbva6wzfQM
gU6Dgob0Xh6b8SqbhRnYi8zFmKGhVPGi0K5OuqVcNyjd27yXs2C7lP9LdvkCwDVV
OHW+7tNmxwJSzCWi5YJngzDqflwUqq4DO+TM15GtxnBfgPeVxWyK7TvOulVGh4F9
/w/VAB23vgPmKNC3ULNSsby18IcZNuc1iXv6c+QrkHbnWe83JElFFAvK3tXPObXi
tHhI1OjYTDrBjk+qtrKeItItEBJt5O8GkkXcqgoSxmTM0B04Y/5SDZBMANZCvzJY
4plZtteOASzjiulKTCbfKxfKQShEO+0yketNgPMBSu2aB/bm69L1TKkEU2/Lsj2u
l7s2PU3SBHhE5jUp4S4u4VjLSSpYQacve9Z5vTJ3bmzfZJpGEDO1+GyxhnELmcfP
aFVtEFpYopfAYIHirsbq94Afw65IKw1jH9FAjUnOCec94pFy1C/t2/EFbiGj2F4B
lY99hUDMqhtgoRCBpCqa79rWAnAXUhibvWrkoWe4COdGGXlsZoIxWg7SEd8vdCsh
ktQ7XY2xg6ReFK7BTb5bhKSegF7I+wp3GQ3xtyRrVVDhGcnz11KMtaaXJiGEny+0
AhOJVUK1leLW3jefyvp4+CJEQ2Il69PtNeNCpclhKYNdCXSWUrzsFTxTGBqJGyFR
7jj80VgP3pF9i+NawNsKBe5GKa+Xo2sa9FFmOhqNe35fIq8CNTA/K7RBHV/fWacH
tQSDCTSODMmVlEpbRtgMMQeWxqqaqH5+Hpx2LCZeNpFddhFpbK0HkfX/as8PRTvq
PsqUn6I3oJ0l0TXxwH0nC8IfIp0bAvQ7f5URS5ovubKMbRoELZQPKGhiXRHXatUE
b8/2QMOIwPjMKqqzhV7AjIm+2GaqvPpbEJkfPEBzEOZ96nfX4hvkVmcQwdh76h9t
55v0ORi5vvxYK23nH1sxt1uJH2GHZ+OEb/0MSouZUkhXeKA4j5551xmFm5cL6fwz
bYDeXk/MLQMs13auV7Xx5jCjmVelqDjsEfMQoLZzDCrsBOVxklOpot68+lYFhcZY
hbqBGB2Ll1lFFJhdshtfVmqPkQavxFLzOAXRB+7Sws1mxGgK+X7avo+x7UeaTrFx
V3UL9Mj15Ym+9iDL7el6hZRV89I/Im4qRBI0jr0mb4en4uYH1ftST/LRE2lzpbXp
PLFoa+s7JShsaPHKRPFqjQjJ6zxTzhJZb+y1AsbDEqM/Jt59VSFJXcHvABC4syEN
MF7xFB8EGvPpD9Mq6iijQJCnefB469K1oWrumen6tRnMEteBEHN6svNMSgA4cSWJ
CDAvCiAJ1578uL8QVXGM4jnwAqLjcJB6KWDl/6mRr1d/prr9PxpR7IseJVxFtK71
HUvdw5G1u+EaHA6sfg7yUdo/e8OnyQgnUwWmssvQp6sxSY+9sS4wlT3UE8u3a5vc
5soh4EZyxt8BWvqFTazQHDdJZoqFc+0hceiaE//SKGKTaBJomy8P8Rq0py+AgTM8
xs/2BeMK8e+meKwTMVMpbSe9mp0cC5i/jz9nOq0Pzd0KZUdPusQ2HjS2VyT2RmDt
lumXwDADZ2KwfMPgNyfUSr4X+1uBHVjb5NW8nTUQkhCf4J70IN29DSO+FNSOcmp3
RaJ73UWNY2vUehT9zVaC1DAZWvZ65md7a7FvX0+SGceVoVkV/jFYI8QmSok1GyyP
CHe27tY8bd0dp0xwhZUBwmIK5MS23bKxOxlzc21XqMH6Ohge6GuuI9GXbB5DC+eW
xEFW10jR4mTT/8polYO0uqc1azvZ2y1saMbLFgLoC6DovxCURUpjMmC1snD/1U+f
CKzKUflNcuWn3dNGSsjRm39Zl/hoizWO8tKkDgXenj/d6merIVaU+mVPhScObXnR
wIDzilb2Ag4Ow1qRoaVzhqqZ/532crPzz8qFR7V0p1Vl+HBrqj2KWZ860Rlu7I2U
G885ZlXzHl9PVuUW3RurxKnnrwUWsQH9ZWpdTAoMlHP2v61xvE5aoZiQHp4dCmJH
cKP0CX2GM0zg0hGCSpI91W6fpvaVxtteIvPQxWCwNRofJk2NGsISMRvTREI2cqH6
Ao3Hmh6pRi0z0fYJjubF8oB5AgrR1PI7XJCheU9lNs6QqEnxKCSWFUmrg2FmYU+k
digf9E7YJaqPr8up2WUtFCxOQ8G7YeE+nS1QMxT/Rje6Vbq9bi7OUioU+wElhzHY
qNzpB8sMhZRRIJ/GNXr06QvA7ocxYCzb73lGKrE413JOcsuVqMQAjLt3GomucRyx
0LXlmFGQho61FkV4SvFpOuk0WGQMNaFPqzcf8RbDAepgry0CawiRmOM81Hp7fcp/
xpYW9UCggN0WaRGV4MAK5wAl2pwITXLzx7Kh9rhvNOS0GFkk4pssz3Yu53xGvehs
E32qNBSdGlImNIPZJZyZwthGzA1Y6MDXBcHMvAHyxhjAaX2z7KqpLCBq9csmh9wy
oXAg5XGV14Jw76aPP0yXFfERY43Bn3gIbMva1q2R1suBTp7xv7O/aQ1lUzcHRq5Q
m9kbQjuGV6fwk3QiNnYNa1o+G8kzqA5T6xTmg4n7EOZWCPgtOgnysRrJYKFaq9Lo
nzZ3hsiFBt1aQA/mtaBtxKlZ1gtS5OvD2B/35m0sCOXtWTPbZBp9PXrNBDyB2KCY
Dbtu54/Ru4ERsrcxSCnxF/NJrhgOAsLDYKnbGYxXRHx0DgDKSI6CFLMBfCNymzBW
XtZkLbj5hG8hxRe0X6tqIieZYu0ZO4RaxMp1i8obwlx2ODKUavQwlBk2ZbqlKF9c
/pxtEpJL4BnaJ88HTV4txD7uOSzbzw38jRFEi6sMT5SuNvmtl/W5nTcgxYr/Egha
egh3oG2gh/+qEN8jEmtTFQ6QQuunPfm3TNstk3f4Ud91p0hNXMAB4L4qnVOLMIFu
Ch3xzv8cqgCxwCqPSAXWxMpn974jx9Zs+5qtTw2G6n1lXvNLQ4Z+TpgYH+wlsB67
QHAmDclMq7Rp1lXPrl3MwnqGQ+/4BWuI4DL8NxwW1IocRv+v3qW7yHFc6COMCMc3
kIPxba+Xuqtw48qK65setecPj6orZn8wQWF6DkUR7rXCtyM9IZCz8lOICYiFHpEj
EMzHbNay7zbtUSn1yo0+ItoZAaDq3ToqvPGQl/2x5NMCxpGxofPS4Dbz8Nz9XjI6
QbfRxTn7AX7wYNEGRXwG6HXCMNLI139xoT90OL1P88Iuwh193m/QDxFt4BmkotjF
pDAcwq6rc7mCEf500ojyxvoTODG0de6P9Cp1J6EWu9CUdzYvX4afk5ZrQDQOxtEc
Xl2MBl5/qmcJnM42o64vCCimKQoTwO6IZLOrE68zbRYNnizEVUbDNOpzCryomuOH
klYVtoBT4fE4xKYj7DcWWN+XD2GxxQ7c7YVPVE1G+/RLANAXVfKOr5aW6zanXLBL
XttdaLf/+dYbbdgKTdiU4WDxzzTuoNow7K6DwfwK+2BfuCWGXYzqvk0yr+oo7OiX
Y9nZcTrIPsIxqBdPGRrjIpWAl5QVGiGAvj0qQTHdqsf5j81iIzNjKQAS/dYJfJDV
vLs/PJo549t23DKqH5VA5AA/wrIiz7ofIWfCA6gjVcqLqgrhs6WeCzL/Kz2p35e8
CzuIvrNTDUREaksiERBaIubu8EyHhUK9QhSH4E1WSn+desSTh3fVBFxEhP2DvI8j
yQbXjJScs11K0tQ+IJYgAVm2WN5L75K5nObnBYxycrvfw4W2iCFXknNDY6E3BN1E
IBLgWbNsQMIlx0F8uEMC9qRwcXS3oMfRUjHWxda5rBYL7TGybML7xPCMfJndw23W
PY1Mj003xTugwSQUvS1R5x4MENL/OU1KlmoJfBaMyZ++6lQR38VJAaqZsuvU5bX2
vhRI7syg2vCeoTjCga3b3d7eep8l2W//ASZlzbX/LsC9RaBTL4Tln7v0qkBWcuZ6
wzHbh1jY53lDrTpTsjYDeMEMnRhcarNb1OLtiWJNCy1KkisjkphyaJ0+rj929f8e
uANaXAZ4hIDS8KWosWoTr3gVBd+K7omvjjmxrjmH8o88bgP4yjbMN5QVUo/tsubb
ez2ckwo6Z9Kuznr9veZi8w2QXVbrHe/6hFsdsjpnazPFP1xAa7uXo3g97NOBILY8
KQryU0mM2Z8lU5Z6yWtInZV2WF25o5mM9vjCdA+/SL9vIujjuCFXsSFCI5mpuM3a
b51Q8zEU5ubenmO4XfL6FhkscM26u0EEWL5f867fVdkdw02NPpY5lqpaMS3s5VqQ
qCR9QbThUQw31P6wT+lrCYva0A709rCHuYjwVS6KSU3KYobMHT5VFN6pJyJ+Na0j
5nO3B+V1pkWitxSPj5gcJpgEdqTyAxLsalmAGmjKTtEqemsZsoyd5wCvOrWyCi8M
BrJTlgd/T2b+vuOvTlyeUweZTgJxDWSLSmvni8qFqzr20MDhFDR+OAaVoON5k0AR
9zSyUDZH7F2towleLJUY9GJHvv5/hul3nmtY0ZFjaa4Df6b04mD2koI54vcuoWO5
JCozzyGM6zjLTJccCgQFNmb/2H61EevjMZnVPQ1wp+G1Rrs4pyQA2GhdIKJs99HF
LK1qIyBLvDfBT01y7CVmXg77WmJOlNbkJDNJTSxjxUxM0M47IImbdhcy8P4ic4ak
zsTdvCDet3NCaSFC2osLPu5TlOjYEd+S/4/TLBb8dTZ9N0qetFUNdrHiQdnsNyu2
FMtHYmcsUTZKhZd4RenOKMc9OR3iEqA8cq3RysaLBXZFivR60bf5ELjh769/WWGu
NJncO13LpDjZ8a+HtsWJgA8COAkuc0J8kvkcMztjKv6AdPe/KEE1ytFKy4iZo1IJ
uijPUE3TrYeEJvC18/+UOG9pagenN2nwmCtaot/NIgXvOdQQC32QQl1Xvsel32TU
jq11+mIAIW/OJxkfApBYH9OCMd0dFeJD/dQNuHxp0P8GeB0cQWa5pOdaC+2BiHut
5KhafdaSUfrsW4c5VOVAi9yEp8Tsgo7vCai68xBsBUbTCiDxaJRo1k2EsIN4KEOh
yuioFvIYVDh85vJhKJuew/X5khgCWRmGbYj9CkZfGR0fBNs7hJQC+yX3lrqBrqku
WNJdx4x8fgKUG4WO45RHXRM37ZC9LSInDYmZiktX6yDcaUKbk1Nm04epiESWNDNy
czMQFoFW9KDaB0YSMef4dy4Qm+FNSbrqfwjB25AvZzWzRyBb0Lh1S3Pr9BwsMvMP
NH3mMGJ79Yl1u9VIPWHtGL4BAJSw302utg9vfgfEXrQg0r5dtWI2qAC5V6eNvVX4
1vc2vwC6Wkn9vGzWKWEKfgz3O3sofHCMQ97vvM6Kwxw6Wzrba1JM1nlNaVCVHEpC
2uPChglWTQY52hXoRA4cmGQlyMpkYWT56Mw00Km9vKYfR+vCIXRxrybl1m3cDmAQ
D6J0FVGiU4W6piegbL0hayeb3MwyB/4fcu2xq6+KV2oJD1yq6/f4K9wacCxE9kH/
ZikhRGc5B1GaVGzSJtkyXmAT38HyPfNsVQyQ/kU3sV50zriWmZSGhvRt73gQ5NhA
x2oiJOEjv8ePKYdisL4qvpmkWEK65MF1/0EIpsufKYbhHEQKkpoYeZn+4WEOF8GR
Rfv9MNyOuSNzyWX12GysHwKBntZXXg0rYV44blX3zcAw936LumLzclcKEwmvepQ9
Klz2qf981+0Bf/7NQw0kdkZn4hFrm4/ksyqfLAbEeeJ1M7eZlx9kOlIPCywF1PJM
U0LzDQeWI9VCttz1rUqBCOmhcHZMa52PXbZ72cUByK4adWbkFTcjWD8qYzRCbxpT
eQSNIKnGUp369b9TDHtcd+wVwCFKDJzKL3zMm0CLBqVST2UxhBORn7nRVhFkLtCt
r6U0bRIXq8457jcRQ7yesWa5GOGc+gioa61ypb5+IA39rcUTx1AU/YhS99GPar0N
i9NYo9Y2hpGVH1dNzByhRHcq9iQwpLWTETgFvMGfxLr6fKCA25uRMT+jboxiLAMQ
jdFHT7FconmcOgQixhTzc8zb7i3oMpg08n+bBCqzsZgwpx3Rt+TPoRy/PKlnwzDz
li+7RhUPgLxNKGRA06HhOX6vwCLQv8veyXGRYneKeAtoQqRkMWvkyXQ3uqXIoT8v
U1uy1wRKOnMRdmLF46DpugxKmxzu3VZ5qExHPCDaMgGEqjzl1uKtcHQvHaskwMwA
CYwXVsEHf/y/i5j66Ll6yi06QwDqvNqbAYigtkQmsE3doAfDHmDLtAxLHbYfjvGP
qxADoXL6tedIrvhVJXVZi2qanQBh1kzzgpoaY0a2BIoiV50GKhapnvoV+A1a6pxU
ijmW5EMxtcsTcWEEknqkTZd6BzCMZIT/HwaE+I9d6AeIU53rTjg3kVxgMqrECChN
b8jf3lSd12oDQ4upAUaCIz/06pbNI9Jo5E4PuhIDZEIOXnZ4lUxzGrA3tDJFTles
ldfwZQAqRH3x8bv7ueFnzHrT9vqDioA+S0oH7a8XAXNhKZZKYFFa5tfQ9Fr/BCPR
Pfue+mieQvXy7WUhpIkt4tvu/1ubK4C9nRsz/q3RIImyBhjxaXBI+6Gdl7P04HGz
y9IqO1JWSi07STWxnuKzL7DP6dEXbAQz0SpMPWiG7nyG5cD2gh+BJRfHafM+DFLm
avzVar8UrQTe0gUgjCf60bSn3Q/Q5xiVOnZvlmVx1ng6kEd2jVk4Obv1KNeMaWRt
FYieS3FCR5gmpdycOujjaFGza1T/lb16tayetH+qhe8iC1uY5ugL2fFAVCebhyRf
feowiK0OzTgqb10b/dnIhxtCDZNhTEkXzU3Up7in0Y7HgTBEX9wTADY5fxSMARdy
ATI8fWWq8gE4uZDnyQtJZCd0uRWysylMCvpzO2lD5u0T1AnUmx5jqEYmmMMZgLxc
9lMd6VVxSccWpqQV9LRnGCeqOisFTRinmEa/28g4F6oPkRHX+fLNcQAVqazVolCb
wrZSNT5KC+c+cxMzX7MOBiWk5boqcsw83hJo/F0/OITAlLe4e5AhCsbQ71EYhoF4
ECvv4GFZ15M5GctLz6jnpVhAIQCEvOqibeRqug2bMp7vvGuOlx9SZKk7XPqMV+HJ
87rjvFTYN/r/Jvl0qWWP7X9nKFi1kQHwBFtouyuzhGq0aSOSgO1KPGqEoD7MmygU
8PHv9O3VG2CB4lK/7cyL35MTr4r5SkpEn7sDpCHPS3WqNX6ZM/9jNGkSKX/zxX/1
z22gy+EoknO2BVUb/CVJSKFhmSm6vUuiWXDw/JmHHC1123m51mBf9fuvci92Pqqm
8TM9IslWleuZ7evKzPR68UsWuhAT/Atn33Vu9O37p727Gv1kLzO8jL5HB9uxNLdU
GvtjYxReDUIZ4HCB3QaFN3hn3nl8TPKU7SH33Ol+u5IHKhoU/cEKAkVs/OrkyzBq
RoTRIBubxRDCwVpYg4YFPBv4kPtb68PgQwKXhOCnRN7L+Zt8e9AjmFJONTVZdhSz
agjofQaEdv2BPuvboyCPJr6C3ZuvlaMEip30NhT6u2nw60t6a/sHlKo2tT7NwvhI
Ws0XvAPKJRu/e5JYZujZxfM8EuOq0+wspQeAjC/Zp7QSqUrX7GgQaTBdcDqh9qn5
KwL0NnNZvlw+vpIVvhPKuj7oUYHKOrrezDz00Ncz1/9QochKLaLscX1Jhh+0TONz
fTyoYCFWjp6gC7BMZMzV2cS0WbWLoF4zuh4O2zHsDEOFWfVWjXLWomLPLvdXgXRd
XqxSdB851IQUB7XNvSTN+F1Vc2f1B10pC3HDPM/LRAI28jrHeUDPnp5gnc/kFdXe
bDLUe99QC/8n4OcOBexLKI1kUXcJi4YGqWJTojnTZVzt2COxQmLyUYg11kUlT/Wh
R9rjBcrftblE1VP++IezZ3kVJPOf8NdrW+LWse33UVpNfNU5ZPZNoJqJwOz4hx2M
WJ3bIRCg33flDTDAsYRZJ7j9jq+SPZxXyVfYI6q0QYDrxVM7oTrAzNvBdW0mcA2n
qw915/0/AJuhs9j9Ee6gg+wzoYvdulk5bTyHmtjRliqOVMjVD0FLglO71RhDcEn/
FI8qSw/cG8algdXgL1spWoULPlkcfoi9DijNGwszoMisM3YtNSywnwXqHPOaoYFz
8rltdj0jyWJqsFT2YLjpJJEt6JqqmsS0ZLlZqlEPo3jhFBru4hAc4EK04Jly1yRJ
g6L1r2YH2obNwxNc/MBTNdaj+pWuHZ6G91hiQb1K8BQMV1mm8jLEWX+9Sr0E21Fk
5pShVheOzchrlsOt01/c3OYFEW+ltBDpttIBEKVysIIpkXqxZNLjKp4VUeJgpBDL
cwLwxaZD2bsGWJswdpSp/JS1C5mpbJB5Nompquhph04eFL8H8fHBAmDDf6q8fMEA
4KnNa0gO+4saVvYcHcsfeXClSRhBOBY2JgvItu6aBVHM3FA1QeL1JGTOeQEXLoaf
7cWPVH7P3GQ08yUtG0Hhi7I0ve6vwoOHklHKM/Q6sWrmZKgUnaO8ypZljFMeOPE6
GNIsSux9+wx+quqGsIhbQDBWgyKxPTW29kwujSZ4CKSEDflLFCHtFeTgfeN1hAbh
bG0H+addq1I/y0kisIFIahlx4oIT3JtYKTqPYW/sPnXzURe1EJgL9tQFlqmV/r12
EPRP9TS+PF72duIVQGFExZ9eRBQ+TNF2uqhkx2x0NSS1S/gcMtDNOXKujyj6vjEJ
YPXDrPDuoB4cEzHz472yQBFr+04xRlF0Of4ta/I/V2Fm0y8sA8zK0Q6cZeZ76FOJ
wul7k7JL572TzZcB2oynIG2k7ehXCUe1hhAoSVUi7QXDUBjzPVuUi1reM7T0K0jS
HoCzCxSPtylbt0Bq+WLi0ZlvH1lYyxadKW3X3XhiXQp1x7+enfk0S2TLKe6WmNui
aH8x4uZPQHojg5HIGW/BSTfRICoUFoT22cj8eous2nMvrGA6r+sKA3ZNHE0iMjLf
QuZy6LcgPrCmXjC+9nMe62xdHzbzNpjz0ZxiPdcyvmzYEF2mIu1TCohspcEAm5+T
8zUp6gXStnrMDs+WTy2hEyJFARWX1AcgTS0EPobnarKl6CaxGje7MrE47CtqxpPW
Gqm4F76Ke8/vBynmIrXm0CSFY5rl+QSSN+YmHiTloEtbQFRt22rH8mELKpQe8V7q
5kN0Lk1z6YaTwN79CX0PBAAiwnW2RRlahHPxY+2dM0+vosR7Q5OWulWLIHtSwmOs
XRu4k+jwtqcVMS7IqpI/y+KxsTLP8khuHGvi3mlJtnVYxp/fO5Tb9Ze/skZg63bX
pu1QcIweMnHNJvhrpXVUa2PeXcPJLEPwbDfxGcOz1NtVfgMeg5cNmuoBMJhekcBH
Jgh3zyd3HkLxC4umDbhx1IaJZRqRKjqnANRHc8z+Sv9Lm6Jnsf+8P+kb4tGrvz95
H6t1b2KQWh9io5RnM+wCN/YUvDHazulR+pjrZw7VCC0woTq3jJ/1IsxFRfcdgwaF
GF/weRd5DrdmT0KTsIoyz4W7w3m7lWPAVFG7cWtj5RwndFsyvi/A0AGPMGjTqIFf
IeUqIQ7IJ7VqadoG9isdGzHa3foZsEkGnr+b5zLXhchs86zMHKQyzQQ7qycTeMBB
1cAlbG8L+C27DCWA3TYK6Yf2JexzJjbjGcebGFshpuJOZbnmcYKwZjdcflqH2aGl
dMqPc7kkWdid5o69PzKXDUASWzz+4ffb3zvnkOQCpywdi2B4XXIxdCSEulcZPhgO
Ra7F+nDGhdLdttKEHcAp2Bjb2BzA18rLIZwCqkUCOG7+XQ1sgPqCu+VgkS8AJweC
oSB4pDGCvsAEQPLskmUtQkahdZFy9Va/mTtBs5g+KUDe7Cq9EmUjZ5kXjlzUE4o7
o+sX4ozMYh65q3FYdmg59vPdmbBxrExTEv0nO7pEQOPqRppNyawY2nObNlpAj5Qp
9cUNPP4i00wP9MQTelzX3WQCCKoODOyptseGfaNlGDKbZ6R1TtFoSeAEjxpnL8Ig
4EyJdQa9Pv2iABPI5Z+xOiUfZklHrOShc2cSQqxz8MAezveCA5mPfYJasONtrwtW
pSP1M00e2c1cWpNFM7rDn31aeN3zpqR76LsaRQNTk4qeg8VL9htGac1OZxQJvpCC
ZkWEbfkg6K4m/VsRhiI5Z77sy/YeNX3C8hKXS6BsV/RIfnBIWpOXvimA2px3GOvv
YdsCzgdThhskO3/DAHLLGFKACR+O9SrIv4MaBRDm/6Nt5Xt2VLqkHkEFsjGz8/Nc
NIlYkrpX/sDwytx3Z5fVHb/FYqoNAzAEP7s+seQNXQpG5E6sygdYNvt3Y59DLnL/
2La8Yeo3pQbbFSpBPR6L/Zr5jkPtTpRcAZazjEF/dAWFXrgdZMhI5zwg5TfqYdHw
eJTWFE6nbaey/URcNAdXQre0p4A9ylGB3EAUZwHpzTCdnrljzDJ90Jo6focjbIfI
kUMLdwFi7BbU6DZG8AN/4X6ouwKjkhh4gNyJyHCMODldgBJCbdsq0wDitTGhKyt3
kf8x8X3eOxEx7Tuax7LeNVMvMDJa5LjMB66k6nHiqfc/TXB3oQN+m5Vc9aKXVAES
3352bosnffB+bJ13XPFGPnR34on+zm6nix6Npa+6WsdtyWtTbkPji0V9Ll/WaNE+
WHwvcjHaTokNkwnCXNGI4NWmU4oXuTDMJVutDKwv6Z48A2MgvXFN7lAImiMeYEls
0xfGAkjuD4lvYBlRP+o1b2nZF5N7dmvDV5jJ08OM6lH5E1NsE/msUfAbe1WZpuaB
qE194qrKRHrreY8HXs3b8hq4nblwUeE+IJNSn3GXDatBnsoCagd9pibIKn0NP4/B
ovKx0bmMQ4hxTWV4Lv8/gf4eYyM8jHOd5V0EtcU9RDSMz9yHc1elYlgbDkVPFRnH
wvsZI/RIHSd7Gpd/WnUAowubhE+Z04isqOMT0t38Z8yNPeV9I6CpoQULLOaP0e0E
6wGhjBjW1w/xQoKaxy/ZYMs/sQax/F/HwoESq6DxUi38MnrBwpfTUlXH57+FXadH
5IyDFad8e1FmoTR2/XoG0rBEqSjaJqtjMEmN1bWTmZnDD7EMiMXuPlIwuM1CT6L7
dzThOs0AcYC/XkLhPHVZIImGV8k4xsFnX7NPSqNAeSmJYEh0qUwjcT/Bo2GB08qc
ukX638FPg1rCS45R6XeqaL0n9irDcUaewmoixlrejGQDut2cyi+AwXgs6Yprln3I
zr1yIrDq7iNP5SR4SeDoCm3NEGHxEvzvaW+1k1RueBsEDXM84T5MFb5lCKQzH9bz
pMHUAXZ3qkzhjYPFH3TBlF1uhgaslTyrsXZRCO6nXt+3LL2ClWLx374JpB7XFiwe
DMocrseszbhPxlc0XrTN/LXbIvSIAUbNPsulNvxsQalvCc9Lancp8ljTvEEDY1xP
i2JkSxiOAEmDgAeUcIosEm7ayd7HMxOAdbYnYfwZgD+A4pvT09Pp5sPNib/PNauD
bvWWT+fnOz2OEge3JXeXC+lQwxCFdgdQhpjpZXjJzCnhu/C/KcquuMyUQhB+FN7x
KuJqyeNY2R4K96Z2l2nQEGORkV04DdRhrTtQq6fjdA/8/JbxVhjzNrTIlR78KBHg
C4xaNSw4PrdKaCrYX9x+y2GZeVsAqfMC1WHYeQmc+MAy9KBQumfAhuIKaawnhdv3
U/4syY1PL2ylNwg2dv9E8PE4ccEBDh8+fiUJVzhJdpDPbbRqSN9R007aUQL9DKp1
ef1Anp35GagZJN2/gch3MTCSQVehb7n/BR5x/F+w+clbzTGnKj10yRPIgNg51SFp
p3mLACB7o6nQMAx5qB4Jnjy/grSNA6aucLkGECoMh5rpZ6lzLkbwCmvtO1xp+pqK
PXc1Cp5Va5BZbRCt/YI4Zqle4i7maW/LlM/Qm2u7eY26grLcB3m4e3r4vhDoDZvm
Y9WmHPJxeTwkfbrNb/RvvJ9bw45xj1h/OHqP6tL1AzEy0Qae0WTyKkuaQY2D+mBy
j4Eph0V+2DaRJcoN7jR3+Wpc8FepZ6uRALXLh8YKg8MNsBiLdKBZx6o5xBd0kXE6
KXCx8Wq2atHUlYqb0JObPIFdP+ehj4Iezh6iqCBjv3sXj4MKfx1Gvc+o1D08yOq3
MODQ/9e+X1WnmBItNXNtAXJLJzjhZgRjjZNRBTvYY3W3x61GJSFMWoETu1EQDrev
9nucUIPArjtvw/525TX6ZajndjXiMewDepNE5E+7ASsZpSwlyGEEOOphnuEbiZa1
s53EniB6VCWU+AhOgU1JE4npwQEsYbpQwN5lWnvHEBV0mObeSbl+cniR/yHagczv
gPCXhYNnD6k7f58x/Tkw2DlKzoorenx4mO3giwr/tIq+4WXzryM2NHOh7HqKq+fH
U86li0UrsHx+naUBljNLf+1OA+TB9tlOMUHh7WWbXLiI8VkZ9H5xSs9cy+S/dv4/
ui9W3ese2MSRwIlKRZKEDHsaqnezA5rUoaSPvE/k55+XHCV6rkS0F8RYxNKGlnbY
RxxdMfiHVPnjUw80YA/Hpa/YHLMImTs5npddgDbIHN6T9gTvgxKitVEY0OzfP/K6
AyN7EAjodh50qJRCOvdlM9xfnTRp2DEARHl4Fvy8RTZitalyFY84xQNF2au8xISL
EFlshcaRzyDxhmBJ3g8Bu2E9O8kwLlG1hA8233nBYRsMN/HvBH9QJj8/6pcAWfBQ
FNFOTXldpVG/YWTLDaeuQCeXAbAhp4VJ9kJ1V8ySaa9nVdmlVb3k/he2d2YHMypw
MNDuH8OZrKhynPTPPznfpfQH9t8ugRpD+yeE8JpZ7yofbE2FWTZinbnHEG54wZwW
a3BZirICiEBLFGnxa5GR6MfdtCWWar6STcMFxPUMmUi+JY43Ea2RIXHIx+LR9M9K
SyWEWyEPbHclASaUzu0WGzFZufCi3m1HuCV8BLGkFiR0V+xEUAlUUCHHaT16EmC4
KMsZy4i22XPgRNy8E8ZncPHi40zc+xgFqlY1VuQELvuHfKcHcmIGc2u/HzzOb5Dr
P8v8Qu9m/EUJky1rr92qE1PRTxuakzRcatyfGWUulqPDpLKjzdQUaTGXieCyiQ/u
1tVex5DD8e8H7GUYc3uQzhwWN7cfOJ7HRmWh8HZ7ACHSMSmQ20SoRtMPHjgKAhSS
9Uu0jN6lhtbtPwzY3pR5ANXNOzQackxtN5wAJf3ADIoAzHrwEzPytPh2ij9WCSta
AwIvykA1V3mbSL4+BjDp7sevdWo/x78QOtpi3qs0EhzJwFWXlBQOu2dq/2m1oFeq
IEHhgZU5Vxjua7sQFicC7W+brgSH/NoMDTqLXbNLeAxZ+IyGqX4OjOFhHxslLJAf
Bg40bgFBWQAul2kwm62Ta8Kor81liCLLqO9qV2b5BEYoUNK60neWP1yILUBtX4IZ
b5CgNBtCi2She2aEKa5hmGaxN/9/1j55fQz/iuwNW0HziGiwOOMTrTi9StGqxdc5
0QZuifw+z2FPSxspxp27aaNcDoFEzLQaFDjac92ZKSpVOBPwYKkm/rt66WHa7o1J
TqTd8kC+XqRGpq/alX8eygsj1+vU7+GU0dDYeUpLEV9rn0hWoJx2P+4osnSmkwU9
rrFkgzBq9XEeauXFbG0THYWgVkAGXYXExNGNpQ+ZckjQXtZ4OdY4395F3FtUan1b
JUSiskSQnq73fnOmQeT9zMCaWc1bYsWf5NjOSfAhJZGWpyQi/AXgI8rhuZe/a45g
QiYehxBQl0gaRMuN3pjbdkYFl91L8DrMtqSeNziBkU4aKfQOIGHxfpf8O+AXD8tD
bhXFymNwZS7UdIY80Z4h5F/mWNnPRFalodeylU9NyHjWzBL5rZt8j3dVHyNXLSVy
h2TF/Xj280gyNeI2Gsl3bdgBzifiFKq6Mu2FpjW9rgx5DgUXxBYWtbSul2D2oIq9
kHA+zCXcjgQjXpFzKGJGyN2nTUIUnbGfQqVgGsOhCvfGqJaLYEYEioreE4EqKl1M
9IGTK+yJh/3tUUfwa+vJOIAh555mRQZovyfUFDakNfKBIpjnkfYTTbUcpyc0diH9
Xjh3S5/0y4NVtGQTIBgE1DbW6sAM2bgmB8d+7NO+f+0i8k4KNr36FIeWiNf9LUJl
kG5Lj0deogw/tNe21esGBmmtCpIpU+QKEKpktMWy9WRyCuskXkTUDBJunBCoGiad
6fFn5X9Qtxyj5a498fceSXrcqSUg2SiX87lOSiDBmS8ymxz0zTKH4d1WR3alJW8q
/i31pLXVRwSjWD/ZzTn1HVe/F9jLKrOLldQAfkt/hkLN23yZ2eqzWEwqxOoXHVZy
L/uzm1JkVhVitI+A73I+SO6jSPOwAeO+g8by1nUiJHDHq1K3wTRiZPoo7Y9QMf2J
kevmL5/uk/SWlUG5JnwKVh1wFiNkQIZFAUNlSm/DsyVp5xUSCxQc8NhK7xFMrqQX
7Cxs6PT9GPrhn0n7OfEauZCZMU0A6vIwcgb3TnbL7xbfY9QA25mzxpZWqlwdKYqK
LSzXUlBmUwxpKxSXifIzsO2Q8Btvly/CS3qm6Xt2l2xy+xs3yoazsYslQ8zknzJT
JktUXHstvCl0eoZ0Frz7Vj/6esyOIdqyG0GLeJNDGltFH9SMnnJ6mGuJ5b0T1PNt
LsnrXGH1jsFxaK1vndW1xSyH3K3rODN2V1bOL1Jr1Xz1iz9HkM8Fms53lj4yKhdC
FqHGOuHMsF7QvMvY+VUGv3HZTmOvvVx8Nie/ibUkGerL0Y4inE2BLA98TKGLWJkE
HoBYap8ZaS3OJd2JpqBrTxrxSb9fcwCQDPTKLaS6nk9kJ+WPIUJZ51wtmIQKj3YF
wkbXJoQMyeoxkv2b33NS/fni9t5QfV1QxpfNb+t7b2f5gieENhs2mlugTqWj5Bsv
xa8G+C8DL1tcrQbLZsWzQB1yDZ3SVN0oTO7gF68wcao2VX0vtIgiScbjCaATPziR
MvKX+ci4tbyj33hIt3O2z/WiIfBUOfFUbeNJhvKK1+HeDRwp0sz/0qZBhnLPTILs
xQfTmfKkvAm2sCwkTa4+PSTrlT4IijlcchEmz/6OwdFfHG9JCz2qLPBFwo4QQR1W
NDuYh+PfObbF79+E0GMUMNezS3sP1/YuemKxG7p+kRt50iOkHXghlAeIYEJPCNEO
1kgTaVZ/Uh98yFo/N0zM2eQoAfrb3m/r+TQpzpPVoox2p2Z5yXiRvpO3wLStJmRv
m6+EeKni5lXyf6eYrCVMKJK9et/ZbZOakFLdZomBjT6qUx54zRv3Q4PPFK93wqBh
Bd41uPkHzD3YPf0A9DRV/Zh1TMROLhAeOKSfn6xKDNI8+1irIUdaV/aHX1cV1s/7
KZ5Z5zvGrFIZYitBS2ZVS0ytuVMQa7iS8QDfM7M1x9oTrRGtqDVn4FVUzrIDlUZA
t/nLvZ/dGHheTIKSpex+yQrRwjMBm+MhvPf5BgjFFhzRINQcKowymXFo9DPPhNcN
YIPbEF2fSwlC25mBEsyO0whJ0z+hTDAI6O0+SfEt5I36vLIk3tlElcYkqFFOuGae
D7X+Uif+v6oTBfTdLOn7gfag1SedtGMSMd+6qtsv8ZJ8/JXlcALq4EsmMrJNk9EP
sAXm583mFhLvpX2XmPgxcLTAqw4iRQBsTfzSRmNO8Z732jnniOfhDQUpGM+OMH6k
4zC0XjiAOptauGMuEPXXCozC8eVWe4hlj0/m3gKlKIAWTlL0CH61hziOb1+mt9On
JHMpa7P4SWnvXLDze7JzG4YL0cKzRFDvw4G4F6Cn3gkFLj5SBxex4h2iZYnMxUfK
bdkGKaCOh8wWs34oOFe+uR8StvdNvmQKqji5sSqKuwV+gLqJkR61s7fB/+S1raZW
GxpkCdB4aj7dRwR5Wnw1vwrqjN81tCrluu7VYt9z1pk6v8rE5nl05TQ034/dKFdv
c7YEB/S/aE/NrwopGR3yJeaGn0Zj4wSEeOzPhbXeBMTB5Y6ivFuQiee5ZJEQUviV
vE9LOUivF+6vG3yNMxLpZu1Lwh/884lPR7eYGBPfk0Fx36fAW06oBNWKOLcevwSs
EmeQlnqzi8SHpXETn3a7V9R4/vKhMGR44gOW8m6YUVKOUIfOxlOzTOJdKNlBzwBv
LikR9JFKB+5Fuww4z342ZhVSZje+pAAEyvuxroqvuESBnheLo2V8A/aZdTJR094k
l3VWi1MjNy9V4Yc7KdR6ANAEbtGhRRathldsN+ma4LjCwkqPIMsRpNq8gq7tS36X
R5vFbLDuuvMa1vg4I0Za70zaFl0hUqDC2R7eB5GHEb8ZQ8dnOeQCTYUhQIc+dI6t
Sqes2xgVaTATxWZa78WoeiVzHPm5jESaCUueoURVpz2tgjNuXb0TjvpO1yqjchll
+5yCN+dfUOWyuC8H5MxiUNb6Gk4GIaoTIzcOBl9G4CXLxShxXqVSTUMdficV9ezU
SkidqED+dpzSpC3z5Kx+IItwObeKA0lRCiDEk/Q+x4IhrNaXxwuQsgezalk1GuaC
bCkJbTT1ITyHQD8FXKlrvI2dnFj452E1mK9HEX6UpZs9KC7qCb6LY8qQuRzFm7tV
AvqSJNT407fVy1IdjW63b1CRkhpSG7BE9kuHUBieGp2Y7tQ5CEwIbMi/WuvwHzSf
S7xx3nEALL6poWY7f0kxuYnJk8K8PvBWbD7shFIgd3dSSrQfJhhcoi6zwt55VCdQ
8aB03NXrd6NZ3yMXY/VYveevRUnQuN/9teR9L9CpXyvkfVMHf3QCYCeGoRLb5oqB
DTZprXtqjpE5reWhVEbc73JBqokNmIyz3ETp5ifzKCMj2kMEU/OD1HnMulqtA+Wp
RHkMPHxJdAGVnaZtDiLlH7mY76lyBRWdz5MTzicb4bqLs447ISxr4lA58Ldd2U9O
GkPf5UZDxAaDv8xAS1rY9x4JGwrbG5TcHYKtpSgEc/KVO+Vb8uwNPjHGy8ZP7Iam
1XaLADr2hpyk0olad2THcXVvI+w4wHMru/5WYKp1x6fZ0i+bj8QX0VYabDC/MGt2
HSFyUbni2BaJ6x7xdGb+iLFx0l9BVBJFPYrScSdwMc+5a5a3VGicUlgszAhXHXkE
n7Ou/QDqmLj2mPMtbUrUYaKh5ZnPN9YRc7/DOIuaB4udLULGQRcrP5+PDbFgpypv
7jviJMJxKS/KH6x2ttm5+BcfkC7v8rLbA5esKA3J3UpQkqGRYEdgLXlnwSeMN0qs
4oO7TaLlrWc2iefVpN6Tdga83I7Xe4GMVkIwcl4bL2YfrqqF6N601Dfft2GZSnDt
FUnePJW9TmuU6q5+kj7+Je3/e+xhvjwDys57TYlDY8BLN3RAZ86tIVKM1uDD9gaK
NhK5MJfCVG4l/E4ml7PayOt52aiZl0CLnXWE2shR24a7M1ZnCHz7RTRm2AuFmuKk
sRYLZH6oVDYNsSPta5fdvn8FV6QHjCDWdRqZlidJnFVRjRysODCMD+p35jWbu8Ia
3Twq7cPqlxDV69dZvaDttxt4GaBDc9wxadmuV2qnUEZJ8trSJxyJK6rpsc1fuXp3
FUGRK2F60ABZvRoVdlP33RHZht7NOGTUJTQcVP7hkOg5ssnYbKIPknJgYmbTxcj8
8HMwgpN7Htm2f01PLtKDAoQdzynECLcjuYPUeizatbs9+MvrAuCce2CSDKbAyRHf
t5F53IA0l8stVEsYYY2Hjgox22OFOxiUAWjb7rE+6UNfSy80ipHtwegmiXMO7L3g
wOwGb2WqiwZT0lFr7F9QKYB1EsDBf0hsifymTTQbGRRrczFll9BQ0x2czY2IGvFl
PI26CpDESLTb2f91HbOosP1wX0n5a4B3mY6am6PZMqLsmSJUFGIw4Bo49vcQ0fhE
mNuCaCSA8/a4Q+rwROH5ln8trrZeRBwUiYVD0aCiPW1ZJRm2mILXnXW3yw9qrhY/
WZDM6viFWp9Fmv7CWEvbNc+DM/rPmjd7EWFOnxaXehZsMJrXBfokedD17fJIbUmL
coiT5vjamJaFxe4cyddBizwuRTx4ZkBt8aL2nBbBMEkIy72qRsZRixDO3ivfQEj3
cRoy9yD8cBwwt1a6ast0cH0oeaIwYsfCV+z5/4dBLfN8t7GWTMUtzQ4yUPZ046Ut
GlJQOwBSiF5pJhJD1kdyEDkg3S5whcCaeMqWTkOzR+183kgHbk5f59XnaFxvwUrp
EOy06FHIjqzTPDm06YolDPg7yDVkt4htEvSNWuM0T/pXyH2EI6dnOQEnK/vArWTO
7t7cKdH17VjYUGJxWEAWeQfsJWP1DX9jRxKHnqeV8z022X/OTTRQkNXaoyxDfKtV
6OCRjDzHIJQO0o3GYOCbjJl+ZI0lz6BVmEAiEAGVSxBH+DGFUMnmtJ2R98GNP8TR
Bgsuo4sOdMtRmlYFaeekXFacKCu45tq/9MaGW0VO8uSuOZPRg4GVE7lBNYjQXDQ/
HL9N9W92GjCUcqNluyEuJP/5ijYA4TnO6601vrJ+mNqFcGGnrN1FOpmG1mCN2kcw
94ynB93343G1VP/MY4RNDL0BlluatWlGEUCpyZVZuDGtSKHskmag92DD5wpqQcow
78lyinc2UCqAptNXyTdpaHUX/RZZr+E36kzXcTu29pHh5r5MmBSL6P6v2xC9bONB
qgr8EcheUcQ04b7Vb8Fb8eydNfPhzji1Nlxj3Ie5VZX2VUHYELGWyHT4P8V7xgOO
xigGOPdiryvVC7zOTzbAi3AF7cHjWWZ1foOvY3kAbCn1X34GHDmRGTTCQTP6kAi+
Sj4CyHLByYOvsVilKIp8a9FeZGc1UkOs+tvjPl0D6DMSOyUNGWmBXFyo/DtnpUTL
1Y0Qm7Hek33lHHK4nJqV0YbBE7W/gIlXTQEKfKr3CyIZhouphQ6sQObxw8+/ombx
s00Llswwn1p7XHPx6vAN1HxFf7nac3Gf5/Vk10XKrKldtKnFvAsp4NQNlCKtyQuB
/xeJ2VAiA9rIclMbd2YxJaSQwp0ol0rTX4HxWn/BJtpPEYE1Y6C3jIETcljkBsFN
KgySIy9PQjEnezRE+8VOv/EZd7hhJVJzF9LfGDOm8+dGVmT5RJCjBsO6LnrQ//Ey
SUqd9A3UvDvSE1KRG06bXWmKbAW6WeK+EpZMtekCUYpYgbZ+E1a7RWbl9T7vfnqz
UKLmjFyg0rlT0YcAg2rlAN9V9QZ3WWIVxIp6tvtmBZieN34JXlDtx6fsf4wB2TWG
++GFzdXqVJraHJbq4Za2pO67vwRJw3eMP0bRQCm0Yv4Kf0yPLp4zd0nFWnhgWsrF
LsLFf7MSHKWBNc8xzqKGCABJDdGccajrwRo7pbHJlGSaf2GvEmBfCcBBatOKqcbi
cUtwJcLjIFqwcWUenxsBI/SBUhYW0K2gpfo7KRUDWDC9CUboD2FEuIGrfX1W4VZc
93Fuy9fWIOi9cSu0BLPDP16weNdEcIZ4zosBZlul1dyDI7cauk8zwqcS+cmapAOc
zGMouAGZOI/zbCPiLtJhkS5kjppescuHddawp6odQAfsJ2Y2kttbPVfbmnePvrGX
16ui07nkAIEesvn3ac90TwTqLOkF6A4WaTcVSYcayh9hwesoLDz1U42G4YyQ7gyP
jM6FbcmkNTpt77rJNZn/O+jTv57oeTQ1Kd0uAjkrBJ5NccwdifDhvVPjGM151Ie0
LRRPocsZKjnw1hjKdtwNA2niHYN4jtT8yHjn7CMO7PDGV9vAZNB34voZU7lDRbFa
JMd9AmIAktHcHfQyBwW4auXr1+j4Yik5Le+6E2HjozCVrLoUKuT8zGIwmf4WGML0
A+CAQL9eKo63ZCTVWAQMEgdUeXpm1wH0wjFb7mh71VWzEOPvso2DJZFeWs2HP0nQ
oLJtloen3TI+n4GI7VYKzwh1lulgyFKcAgVrVPaHoi8AiruI8R3TFVst5ep7HgJH
iVRFZKuxJB5W+tvt4F7P9xEzh1IiNlFOepV1JvH6OkSkIsE3flR3nzQe1A0m6HZS
QFaIm4LTWVMIhliTWds71LIoCNr7FgOmfQPZG///sYjEQJxPXiOEjPKz0dIFs2Cy
Yp7dU9RIbW26dnoVn8/LSSTstaE3hm+lUT682yIkx8RW1HMfFpG5YriofGsspllE
XfYC79fzQfkycmvhN6PQhHWLDXJRKfdvMTpYeOU+aCAXYvpanDyKloDYEtbgsY4Z
099Or+Ih2x7GlXKlIszCC1CSMSzvK14zTmtftjfiCnFKP017kJNjj+kYr9cx/CXe
MRPCjfr0HXkg9gWIzSHvg6Y1TTMXq+QLoNv5XUiftYEonUw4CHgDp5shrn8MGloX
WMDrtwSNVa7v57Gnvh8/hYiPwRYrb6JWdize4XYf6DpM2/oSKw7WjB0nAvbQ1GIQ
h6jTNxNLFX00h9DEhxxGekrqna1xeYNS1q318IgVpe6rqmM5rbG+3GQBH99+SSJI
GfhXfItRKj8Cm2LnCY0wWcBHT0+kEmWtk8Fj/oKqGiGXPq6Q+yRrFdv9V2ScP+WT
+0HKqnc71Hje4z5Cq1p2QbJZpQEcxD/qkTxcnnriQqbfCCKzUu6zEzBvykkhzCbB
BObmVqYIR+rjRA7vZeyOsGfcR05cxVKjO/2yL6lCgwEvQfIIqwAIzDiNq5p9ndHb
MGf4ewHqJNiBNaNkqvwJHeI0OrOkQYyD5+Xx6hFsGMXzbNyPo7/Onf1c+7p+/fDW
iSjjnNy7/ZS3M24ZKy90rRVzhV/ZMyrgcsaI+n1cuXOzl47RVX5dI/XSRG4P37UX
IzcZG15NssMRj+CQEfdXK+mpbdTZ33ikLMwQrioD7iH9lDbHWkYYCwDdRa6b/Itn
ACCF9bMVYcmYX7Ev+eWy9CsqxDh+9chKIFPfUr2YzbJcCZDyQIF0U/76RoI75Jnr
jUCMBdPAUyOXpviBShvigybylmEAkZJR+ShOavfY+Z7EWWXUBueaLipJN7WX7tWY
sqIVgBzGbG5o/U5cr6vkOlvIQK3dOwSYCzmm63On/S1t8bo0dpxFfYHs9v8Z+PEP
5sQ1ozK7rAsbjQyKhEBQHqbftRa8OVzlULIsnMYslO1x4z/MtMHJJTqf1zpyuBrx
DOdQ8SnNfHaovwVcyqK9NgHyAHOZL2O9Yw3XS3GcQdgWZjlELEIcg0jpp63/+khK
DiCNpwJRbVu8XNE1BLFObV/zEH0LhWBpbk430HxpIFa87qA6x7QTVI46Qwxh9Tcg
p85TNz9B6BWDbPtogopzikooLDPaveW3whdn9jffIBzCCsApX9HBwuUC1k7/aqEU
W8k5t30SKZRkqhm7N/qx2icX+zJLTJ+Rx6V2WCV9aCKysBYTRSTHL7Av88NLNXR7
tIbMcdN3GP/P2oQ4w1l2E6lT8QVu3ehDXVHkV2/z1O+07Ij8BOhVuey7F+B4Wevl
f4Wp59rqz9zzxFzXzERyQTAPNizcTDK3xhCihL26EmPBNq67yDuSI4P65tJNaUmQ
FSuFL9Eo1ana2xCdCfJhCI/n2MkfJTCqelv2U5VnmFfM9tt778s8WDuwWODEPADR
3dxQFI2/+O7tLldyoQVcM5kWehUdfqLoXrgwdP1megkGiUn558bvO0KTzR7ubb0t
MncWMQRWGh9BeLucjZBVFz2AKdc1nxeyh2R7De3ovFZWGM0Q/9vtZc/f+YiXpEi8
nTYl7jlzzwTprtNJBFHkUeEYLwGOCxIcwlOWA15gJK4z5uEp+3x20YqFxYBfsgky
+4/bNvpg4WfLnB0+X1eaxSQzkCIiPppK/+mbc5suYf5MX1bi/dI4vnmuGzU2zVWV
8kKp/AmsvXiXzNUMdZCTFQRbxGMVM3QzlNfWLeVw3dBXjTBH6vkoLZshz3IEV1BP
OmpK+HrVpMsbZ4GHa1fZ+Bi4c+6OnDyQocmyUnTTH19TvJZzoFaUE1z3Mh5TmEp+
otphScG0dALUoJtT+XGpnQFqmJEt84EWEt6VPptQbuVRRtsrTXPQBNgGJEddYE1N
G8VtQgAHJzBQuTjmQ4vNIkyeLsRG+ByUqDBovgSJ3qG3XtSiNSIBiihz2wqqHYIP
oVdoCU+xQPmjW//JZ0/xgqa8gWeRCFtpBYw1vuD3QmTgn5mW29Svqjbu5thlHFWH
TKJe4JMaDT3vyMy3VhsBsqae4uaKnT4JwS67DUk61XM2zo9Y5Kdq1+cjGeLhdl4L
l7+x2zbl8jqar9sVkNoVbGgACjLw2AZ9QrrPgvibcJLvnNFFWSyIMmrYYsYphmIF
nkIfUhjCt3KrT602GTrqddOMFQU/9uMjP1alN/UefPLOKhScBoxVspg34iNlmvGa
SXbAQWFjzRAP6e5wh4OMKdMYPb+HF7bRxz8M2wB3sYN6eIWf1kD0mYuzs3J/DTX5
nbd3qvnaYp2sj+b7KE3n+QU2hGAjLz4MpvCoElK46yFFTG4BrJczOtiS8v52MYia
XtbiSKvaqqh7nNzV42zuLgInu7vX1J0v7z5iKLzSUcbuTtDe0AcA7oobKEDBCKq7
S8InqM6Q6PGKg4hYo6RIMfevvRT6utBFcRiwO9di0GScM/RLT/hu62TJD1gL0soU
jHGrrHFqqeyY2mATv0I9FCDErVYeoSiWOOl+bHyY0mYD9eqCi4cAGgJhmo+dNBIh
EaP60sGEsCbtkNMPecDQpulh4T3qkBSBq+e/HRX24RMNQCnWOSYnr7OyHICcqsYw
Ep3oG/rrhh6rKUGjiN5jRIypN3lyM59xTVvJZsWdODaXLo8Ubu7ashilDkLzX6tX
U53mEIu7wuWuZRfuOYn2INApV5nmPFL/29qYf3QpgxL3zux5P0GAiUeYT/fdReso
lfHRGXucrMYZmIdvnhdd5cNPnTFUUE63sKoyhAYSjK6ydOHpZ8JCuClmKPK4Obby
nVATTBLgdNpiBWwIw6Xd4Br0Wuc5uibgqGM2BroAmcs2RMXXJjkUybE12giCXf2V
o/yFGyrQ/dKF9pE+/pSiw7gyJs7H0sKlITBRKGfFqflQs3yBSIAEyNFOUpxVnzQf
c7TI+6WVfY1i3hZL5IUaOmGtHvqUAMOmFKqsyzUlA/G36AFgv86PclQSleikwNEv
p/7HzSb5qS0hh+CqRSDTzQEX2qHNrF8VyDu251hqXFN8sCRsjx/PFHLYRqJa6Dzb
lZ4rpl6yKpJt2Rbs+5X0Y5khMQgS1PH2XJ29+Kg3VD3IcWddK1zx+nuVtYgqlDZS
Ccv7vNZEieReH/3O6OGuGeq2DZbB9mrXtEOFLsqwgx2Yqe4fk7LmP8i7p0WiB6IW
o8uZ0K2q272HrUl+ZUi/ab/GP08Ld0JD7Jzhh01HsGR0qbUv4yhykRSrK7JPZB9y
gGSkuhvwDmQOZ+9YXSsyMA5gKxSILMH6QD/7f7skb7Zf4UGTBZz2EGziCJq/035h
1vpoxIb0L0BFPVUKvUi3h/yMBg0BAomfQfXraeIqQQf7aDD/6xk9nMMUkkTb+qwv
GixmOa5ceuAHHhFMKp8sXMXIZnhR+j0UijrLXE9mfrbHEB4KIRrjAEP+YZnMPFXN
5NZFFutgRbaiZZFLP8xShmSC/LcIaBX6X5ze0L8CQ0PHpLLNIxpuATOk6Jrpynsa
YVHfSJPbMMsrVDLutV90Q5xA1H0KwfthPHXo4NPp0AVsBAjcRv88HiMupsYN4mGY
iH9YDRZV8vYULZMdosEpwle4BXW88SsRgaMOnFO1g/if71EQ/MFMHZn16jS9UdHC
DAdD9Z/z8lSuj7eYPgGxgBkbi2Wh/aj+Hvq0TXGtFjAFaB1jfilUEhJbyO+TH1br
LSxVuURoPYwiGA1LkOIfg9OF19m+IBNoHKveUdUlzOY6yDC45OESxwJUPcWeMWTP
jiayENHV/XDVZ1MIlkNb2F8S4aFXODvAy8vf8Fk4xrCykKCG1xgDW30KKncAHiuV
XZFgHoyU0e4sqacTLo9IWfsy3vK+k48OsYSwxB6d31YDkSRXxlvVPvz79r1uJnaC
RRnHlPbV+dy5/diYOj/37YPlsBspoPoOVt9EBp07Pw6zjWwNJUogGRJUnBmmFpZ5
VsdgTmzBNzotsShXAmiAi98f1TwPPj1MQDvVOkHGjgN0bGx3xluAK8gyW2OIhh1/
3My89sGF+a+yr10WI5uh2MzeJk1li+mauKqpE0/P7Atv5n0LLsXr3QCG/IrOBy/0
fNqqiBTtDyaeyIV32vsEn/xrUqbMbykOKoHZB/LoTnakh6dBnkS4li2KYHZB+LzZ
p7fDjfOgG01XFh6rj93Ao4mxyi88jY1QpoSxYMp7P0NKJPKfsTXKB2ZpRlxu+wKG
bPNVcHMnFRlHNnIMjFXxpb7Sek4FirH5ZqfblTdNOkKw1BvwAke4liqWDkTD+c0D
JmIws27VeGykygdc6pMzUFzOFlNXFaIBC4JGySadJFI3lYNY1EXBrT9xvOa+6kPR
PSP3lJtSbBmekCdyBQUP7ouyGlr5Os2azvEr+76LqlOaPHUQfRaxjlBYRODdn/nG
jsFog5pcStlek41/OyUKyM//5MYqPjqg1DSioAwtWrTWiXocOxvEzMyvObAQCES4
vNAJIFVAcYclG82ZPnbkSg/0TpS/1eTv0pxRXWoraFa14gVqYjY5tqCnQS23/0FX
AX0NWp70qycIxoeXxUo7MSAsayqBt14090nR5SdmFHLGDR+DsRmJaFLYar8ZHN2g
aZbLKAVe4WtxWFGwbF1Uh8xPuy51PtzK+z6KAo/jhrRyBKt2y9qWculCY4dE7Cbi
DEL7YIidzVy9U+3KxYcifkuhe9+5Xzo3VpGTf6FVAdARiBtO1tgxCwWsSfft3WG+
ApuWbLSSPaYhJ5bAewjUX28NfV/VFT4QgkEvDYaxqdRkQpLiHLdbg+TtOIX4euxX
Lk1lb4SB7FvgpMCxKi0AiEhc8SgsJ5veB5qMXNobbW7gJ831svZ4z6hJ+hx2phHV
UlGT64y5jnfooWuZlXi9dDZh7IQFVj1qCVYFLdXpy+DVgBa/sityO+4tNYKoTwR3
okFtSL1BCXEVjBZjFcNhQZoB4rI1mNiKanV2igRufVDg6mxlEAi0R0ZRFu8aKPAJ
eoqh+5cRXtcsifsw9zr88Xhz7H0eS467UvrEFBhjbFlHwNZjhecJ8GtfqqSynOhA
TkiCE78b+MCYofidhFRvLWNx2EnA7HGtpqzioO9JsMG0G9p1fHU1EbGam5oHiCMa
4EE/b1mngE4WepOzrHeQa+sRwxulhl9/DPMBNQMXB1Lz87ZEYjU9ByHlXDIngvzE
43EAi4CvStcyZDpKJOjx8sXjJnP9I23Yd6TpVky1DzyZXWirU5aS0L7Pe/IXjaoT
Qy4fOuIlgjg8UYZuuwie0LNIKKjl4/CiGX03uqfR1eYEr0eBUfrL6ZAVvRj9nN5l
367W+tdWTUnz2Xwc9kA9i3zJD/zHHpedJCKVxeDN3WfGkUJY+GlieDHh5CxSFfdy
IWLNFqzfoNG0cDLrmz0F8aJgTsJ5+Pb+q5XZ5svLdn3MoPFa6mZqyHDP4KCQ+mkC
LcVJU7P8rIYaS/sUjyYBlqQ1IN6n1g3z3nPYP16E0vltv/JUFlETt7Xmuxbvz2P5
NjwiJZKa/ZpxqmKx1+UmOzb7B9Qne1qkEyDN+NPt/WixHntMWkTR8GH2eDNXmrsv
Q3wAkBu4FVeMCl0ZQGd7WQU7DL+yU46usgO9/jFfOa+43T2iFCVBQjwii6b7o1H2
ou6bdif068Y1Nm0lmWNbmxNbeQDuiLDqbr82o3Jz5IwYjWx8a2IlhyS0nnJYWl+9
6imI4JaVxkTW+AxiNbqhAGIA2N/rAxdYadgLT8Fz4rj6+MBxqLSrc59q3uhL7e/r
ctfIxkRo1Y33UGtuhDGrzWqyRs7iyilClifkpcqKHyW7LB3xo2Cz5NE2O7FHdx8i
fOedBxT+Mv8cj0qJAtTHeBbOz5/0wrdNZrSZJJaehXln5afvwmw+wGwIktajgUIz
SvF8475/W5n+b18ZMV3li6xasmo8sB7pXUJXc31q3QOYs+HJNhK3DLaKCrBFsbCl
Wq1ULsK+/JPobVIQZ4sRInnWalU3XUtIPGWzgFshrLairpnzc6kAPHRjaFiW0LcJ
CXJlEWQbzdoCqnXzmv2ZJ5zJrOFbnLUttBWx4nfzbRTdDD1r6zn7LFJhECQu1ydn
yuTO0uhLGJTPpepsNImnzu0TfRv/p2ya474CkXntrpWVOrCsvPAa6oMkRB182p0e
ediWXQazTvUUisBCBh1QfdY7kzJvNY5QIQegJff7hMK2bVuhDwFNB9X1sfdULFCA
YWSrjmNIi58S1CTxybNCrxHt2Slwi25+99fu2BMio1CFkGxkz4LkGez44fJOOCx+
ec9dbqQHDxZJ4agK/P5xSL/VozTge0rL8v6hKGTXuTK1qM++Edl0asg9getutRuc
BpgoqEE0lw2ezoGBGF+W/nQYrbr1FriVX3VXjbciwN2rsweQsZ7TOUt95S5eUHY0
rqEwWBkJHxOttztRpc5gllnMf1W1MQH2Poq84aFZ4ZYCU9xIm+0RB4M9on9w5kcu
z5mA2e0XoWgwtssmxfdLh2EJdOYWgsdIz81QqgK8dZYyRQEnARaLdY0ACblwBngw
qgV8AiO/4dRhT1czXyy0cxyGv3eYYFi+4xK8AdeNkbBcSIlJEQUtgnWO7CL4C0vf
MdM/6gLl0sVsl1A7ZnJ5cNP1TVuilNAz0kNr3RloJbAx/rKnlDGZq0LQ+YWzsFPY
K7hquRctf/zVktqLhqnQjTChL4xrQEl+/6pvSmHjl7KPwCBKXgQ+EYiNzIUedfyw
YdC9EuSLHYJ2YkAE8VC1CWsS4WUOfJBEtbIGatLwf0O/rviuL/lFx7YXgot0yje+
PJPqgYse98ngRtNONjqL0Ecxe7DjYJn5vzAu2dAERn8l73eNvVm6jmsLod3ps1pF
LN8WT5ckZNK8lRxTq5995ju+Uaq5IbtzB3gLl3bumEt6NSQZCEZnDlKmeE0a9KPO
iCGIQwNXqhhOxXVAUmrjwWD5fAlYaRrYdQohtsURObbzss9sqKUFsZQ2HTJb1Y3J
jAg1osGFZQj0X1J87KpX4eAjfU6CAKD/GKpc7YSE9f+T2/jqqX25GBnN1eS/Tkw6
aEGb5vsAWbgqvd1xXpbVlz0fKFvz9MPLRK8WklpMIaDF3y8nfgjrq4hfFmPPg43B
AiwU8XOlWqQKIP2RYh09MybzDBNebpmWlyDStM1riuAwEWFt1tMMZOWmit8DQJDV
FLrgHPyRcxS4ljDw1jNOGiQsjlKZGywMg5jnbW1VtCvtoqKy3Goa5+OsyfBcjssV
wssEQFpy66u5zvlUScwzs+TntaiTAo283hSiJBOPjnsqy4OVl8mNiuPi3Ugogtjt
8oDGg2R1SeK7eYlKy4IQcrXVIkyxjps/bn7kj6dMArxTYNOq3mL8LA0DarLe2CVH
EQfxf2O4ypH+Bm9Ykcs8G4OGggDIf3b+Ui69vb/7rAMqXMlILmKNBT0Mfl84nPXV
l8GXBcRbj078t/4JTOqDDPoLKgkGMZXkeAI1XCsVVQQwU2gPTs22V7VustB+Ndan
ZdxJrfba/+jURtfH4i2tZRp4HkzxFtMgN+AQvNBu6iE9oWqHKWWPKHMyysDhWaho
iWProT3cHmdksyis2Zm902ZUx/FC4l+On6akPTqYC/Qx7CchjI9PmJA4Ak6Mfbt5
Q145mV1YhnKls8QGuV5jvrNWln6FRhe/WnpiAILFgzYCbg+xy8t4iW+bNq2UlA7b
D9Jx5mcvDkqRy/pryTAa1qm7ZZRUiUZz0N/kSH68M/wnCOo+Sk3H/QLgrcuJ/0r/
xtJuyv/sfCIOmpKtml6hApA3aY8m6+E7qLQp49mLtcSMiv10T9rR5kCVqp/MUAXx
OqoX/4XTuadaaEwBYjMWDpa+0/ktKUPzzlFaoMHe7nfLz+m7+Dpj+IUnwTW9L1Ra
iWxhWFdAP584yOrd6A5ioJWysWY7p127v6+D4sogw52ynaOJX9SauOeAu3ScM5Zr
pd/LOPhpVOfZcgN3YGxBORKkTx4OCY80i1pdRfwPLkA/IekWOjmKfZ6RV2cMinKY
lrV3h7uM0K39e9e9hDg2MVDdrdcsgU7jwMtSmBgiSjAOdCOzU2UaXlCMn/GiANYY
E5e/Rum9UMScBlT57QIa8ZBgMPB4O6eM5AxLdTcI6B0Hcuwux705Lh4zMYbzbVew
7oGKN4G7t+GqaKVXOeu8/x0PiGS/cKub1G6tl3Ki55Z8dWLWI2emu0B5llODFFx9
c4i4AnxWrNLzISEvcgOVh34O/yAnT/YqjuiPtV3tbVjwVzyfdhkgGOANQ+co6ezL
s4SuBPceGNgYKJ3cjFwdv3vms03xkm6Hnig8gee7TiJFzi7W6O97Jr6uZi9F4I9v
oTP3ZWdfqPrqhYQUYlHA4FCFSnqRRZNZ7hms1znwOtXAXVLvPAuCtESMscBazk/2
AARe79Jc1AJMLYfvMm0Lw3/unzKE9WJRcNUIgJGyFePHNFDgAo2Rdwt6A5kKB7+O
r9BSSyT03Xi0i/EM+6+zqobVVX9uPLuw+v5Cjk8XTD4KCD8Oknat4jWAY5Nsy3kJ
UzjBIubE6SEL0qhXTm19YwAw2jAQI5DkmH1WkqtRy0KpCpV9vFAgUtq7SbzJik/H
NsDp/Ja2gdwY1AKK4643MjbFEItgEITyJU14pxWWvAT0E1RlHI3XPhSCg2Ai2fo5
HeeIC5jpwo17Z/xKGhKuHfJjQY5Do57PSmuuxHwEFwoFksZgwvYj31mzfhy20vQ1
WYOsVY9lGWV9R/xG4Tp5yw66corXcuGBy9v2m/CoYZKeuDba/0wt8Ev5xnvqsyvD
cMcJM26y+Ubt/I0xGre2b64owlR/HkXgZj0D9vP0i3rbso6NyXo5OG+15CSappqC
/lLhceYNnY4CnVRfI2oemUGYDch6a+Udki7ofmtj17XZRMS1eB7F4mXtRSrFFPbj
tGgJdUR0XE5goTwzAU1AsSaeX3uI1ZZVqp8tVFHygRyzgy3OkVVrcZicxOz4th7H
xYHxHGk7zheiv6UXYI5f+BxtzUHnw6cobzE3GnXt3EjN6/qpSwGixRgh6NUlRgag
SyS4h6PQhPbVG8qJfe3DGPdMjPZtMgCa5Q7I5JDwNREx2gONLXySdpYGc0mqXzV3
SK7Cod3P/MAt8kwE675aaollGomanClJf3Tr8oYRV8nso9Ig8DGjmgqIsB6ZodfU
l7mh05QiIS3BejAxNn6Dpcgrppgyy6uDWM+0jEMtW+brr+s129dd5T6CysF1Tz11
W/tPvWgNzgQkMWmHcjeQf7XwDIKzt5eO9TWQJ7JENh6dkZn5rYrCfgq+eqC9gIZI
Xu14/eCXnFEVlgoG1get2EJAbgpaYIDu9Wn8mw0g0RktZlJz2tRCQHmCxrVs16d7
qSbq3Ao4MTfT0nI6JSBwm0+erfGyEx5qETUyt3wIYVNxr7TObs6phpSsXcer5iEa
ErJ+F6YLh8OmPf7f4JFgkWdw2s9vho1Z7fvg+Wna33MWESbhpxWuEJxCjkyDI9Hy
2/wNQ+XQ9EDoc/t6b6nb3IULB7jp2JB/QHtQHPe5hnk4Iotx8Opr2dBP2pYOWoyS
5ahdx6bmOo5pJRWntmtpwDeSSpxvFNBHV6LiPd5xZt0MQSiDE0pIfRdpGcbs3v9E
u19Pd9K18Lf7BdXAORIG7er9lcG1jj1PtFENC6EZROJdbSIsKwTFlTJBn9+Jof1B
Ee21qq3CdJPSEpLa+LlpezcmzutrjjQ4hEqKESTnWmiSItniB54K6iNLK4AdT83x
C1ZPKF2RRglfuZyQN3vjjnJNiHMD8dXJWkdIwkb18dh6wmxnqy4KTR15heoPfg5K
UCY/6LUi/O0a14Qjs6f1sv2sJClN5yA410c6XkwdCwN+LCKtB0fkxbdixW0+ZJ1C
/O+42OLF1GzSh1M9C2U5LS5vrpM1HczzASRn9FTaQj+PCMX+sMiZNLga57lxAGs2
rRwiRKP3HGdbTJP16GqEDw/pWSlvgJ5InsnUygA8Vyq9H3RmQpoWxHdpmZmwK5Y3
fWMKG0E/L+URq9cVaWaJEyoR5yno/WnXTe/W+btUBmvYnO0djSTNB+jNHLHtnf0n
1Y40jhw0yyXlGVC6sZAj8R9CO47PqJCRO9MUOAXbuLZdr4lXa24MoSOU2V7vB939
qYpvFZwzDaIWmawu2fQb2xAJHLuE8tXh3/NdPqgdW9qu2PcSVyr+XHqewUZ1hQGi
bOcpcz8+AULJpQVrY6JolHeIe0/8g3hXMQXzEg7zUXlawHjnv8CK2HwOFpTB/o3Z
hPX2xdQLwgLM8VdqxsJQaSy4EL8mPKU+OD69YrdXMS/K4+2hPXs9EEO8SYzNZvjD
6sUzNejSaCXXUnb1Q5ncwBEPfrQwAdXcdciNJp0yRIal2+sDvZMvrEFcFRCWQ+CM
caGyFAHYIVdQHi0u7F5DzsJ54LNjyWbJfxZ7hMc0tRUHOMCjcITJiNJbE/26Ajzn
c4WsUk14eCoUgVmRdfiDEeNif0A9EWcG1w1JNFDv2zKWkq6V19Vs+DGSHW/fIU5C
nEv+CsiaOTiXtt4T4vXADLE3zw3COXc2IoAIlZSvI5TIZegEve/nDW8mY/NnxSnT
rg4RO5HiXiot9e9Q9G8FNXVS+y3bkcZKw0wjY6OwWudylTeH7LzWyATbE+BbhPkH
rBAaahh2uUzhATUFk4Msz61LqKw4NPtxBTYqkacLHzsdS/QXgJ3ZvweEo7EKc7zE
hqf1cw/N1wm10u4+oL/f0Y4Wu/wlwoojmkrWE+uw0TgHHpehHIlT0uQ+zLCuS3vf
c3RsH13ZVrJdTaYC5NjV+7DysRTO+Y6A3HJ+h7e+DRYBpWfN8oSx8ZgFAL7GFYYY
PEycwzhrIkf4s+f/vxRDVuVFx8myHBMhHNtLXU7SlxRTcI9elVTTOhZtZ+EVKaLd
qO/MDx1brVh9tJdBj8o7kg5RtDpqWuDj8t0jZMM0f+rkVjEziRFH3vV4PA7G1xIl
zwRHStpkQc37Z9SrPtjV3xXEudMuzw1Y8FDubnlCqup/MgPmIDitQHOtqxf1mBhr
yKnXvxCG5XazQ5EjPGaByL86BAcg0UySmzGuEWMSav84nEqlrr0ixuLqFMnovpNS
uRtIiOM6u20xOUe1cP0RaUZnKZowR4RwCXzEG7/YcJWZjQw5YGXWYE+30lPnqWrR
jDcOwKBAADi3HpDTnwKWdAJHrgOg0hxADV4ez+vuBDYJF73SbdDHD7Vp/jJiC43H
R09x06VA1y6hG3eHfcvXOvBvxGozgotKBzAxNanzJehRgDsGpD1nLTQO7UuGkbPt
4lpUTPKdiR4z3jbqql7uzAWeQZ+9fnOM18fODl3bxfloNQyanS/H1B0/7JHZ28tH
Vkvfgp6qLNts35h7TsOOHhENLoOju5u57u+lT5fYnkKEp6vGfRHy1yrQz+f+R/cE
+lDZ6zXuyulnBDZX6nRj2opWnYjPue/AFAo/Wt9cdcz5PZxKmPiP6Zp97/qhWWZ0
g13HanDXy3sjctL3bM4zSlUlG4M6o/ZGuxS6imQ8i6ze9+nnGQZJ8Ym2q/n5mCiA
OJLdWqsP+iYfKrXcoJr0eu4POdc4kPBNhIJIpHhmM+3x36yQ+zFBDmmrqlCcJolh
xjCDC31ZHljY+ugftCX9zD8QmEcboFUGwKrXfYPCpiAAuAX7YD4F8KPHmwr8d2Qk
QnfQrhxIcHmxWa+ibp8uVqRg+p50vpAE7aRteKBbNILdmoPcl5Ia/4hi4rVwpu4Z
xn5neNmYcDdkuyqFH7UuqZg7w2U92qdnBea209bz0dJ3mQOEa54V+Ta0kXcnE2Ng
GbC3CiArQhUpkAkl/Hs9rqLC7Qfni5zFln+rh180Ns3NQ4YKk3tAtdpg3bgWql57
kid+sElXWUy/oY59mMpEyaOR7XNVSSKj3JoI3IOUwyGVTPixBAgD1339Z4H6G1Ha
K6CJaTN7HnVQiqKujgkaiJtHVC49BCoQJgEKYEyb6StbuqIg+j+sNOdZnjaQxWNT
cMeSdgxZob/fEIKNGPpyn0x2J3qQ385ZP+3ZpjA24A6xeGhtsSD30pTjtVLubQZ+
6Jb0URpkNgCcbI9bsIxccxe4tQCXPwySaYrFkN//E5bObtMKaMF5eovj5xMFjvll
wnzWNCaiQMWZDkDAHtOGNcSkVmUMdecl8bxv9TgAnBFLKoehH76vCTBMx4nBSMTq
XS3IogunH02VX5BYahhP6hSfuQzTOk7Vq9IqLlU2EWB1YZz9LdT2ErfcDe8k92oH
ErapPfl5zqWN25Hwy1Tenq2oA1vlHEJ0Wje7p+eMhpdNYc7JyJLzAg42K7Wtvzya
30Fje48zPCXzLSLWYRxehJ+kbjZfE4u45YvzmoUhbHHUFDQHab6451/JEC4uQI3V
/Midb6Pxcs0aOa8f2i/GvR4+azbszjTeoYGw2FyX7zHgmOyK5/a/ltzNTdbhU/X0
8N6uQgXEMjUXT3bTSKEFOFPnSWYZABxZ7BN7Uple869PpauvEecdSWi+L8hOIfYh
UzOUXoaiyvexNMhrYBzmjyCm5KMNegUwoRkRODps1HjC6PHgd+5tRmwZYaGIXqvb
Ml0rX08KFkr8h5RCNMYfiU4f3FdZqHheGnL+FT980WPCfo70+hxy9/CBXyazSjC3
evaDKoRlHCPB0MQkcQCAsH60g+qKX+A92+8vFp5BVKTuh8q1pAAX6huPl+fW8I8q
vgNo3wuohSfJMZUg+XOdmQZur/ZnX3hhIEF+FU+qKaius7WgaLh7sSlWurQ0BCDH
i4jrsmY/Nkj/8t/oSQkGE7g1klzYb6gbpKOzDuGYbKO+fKPgZFStizElzW31kwiV
3KnzUSyZXW8FIXdYtJc1bCSFit59kT6HHlKenNs52gaF0HrPWfY9cgIEh7qVfuBD
lL3RmhuZLWHKb4K1Jk03iyY6cy7p8KUV0SrP8QR3x3Q6HZ1cDy1ftP9V27Tk8GqI
aFzZzj77tnMQIW0oZSVFcQvSHTvD25kxDEN3G6PjH57jKIfVHVuNcv9KfNJnlnxn
oAFjTwKKxqKUtfg+RR6zjGg7XPoahaiPWvAla75GEAomMxGpu365/0a592eL5jLZ
ZpAGDfWiTiXig8cKnn2QqJhjn/4cbYprU1S7zTkq986P2ZsspRqdQNDDw6NO5xid
VPWWMMi2nvmjuwlbUr/wxxZZlxVtcM2g3nvA1zBPRkrjs+4cCruWZOMBbvJeBBCl
0XQXoGCMdBX2p+Rngb8jjFHW2HeD79+KltF0z+wbYSiT4DU8rkSMqZqb2l0zmw9k
q7nc8tP/OG44+BcDcaHqxxYJXw5i+16ZuptLx0RHyM8bKE5xaTwNiDErz+zO3Idu
KIlwxg8+tdjzj2mwThhXHGH41SCIp2r81eGsJOkyhNrNHXALFu3sDROtCXNoGYFt
h5ijsBG1J8iPX7ChHLV3npyjEsc+4qpZewy3dkeoXiFJl0sJReDb70qHSbFA3WJF
AudwxIe9C5+8pXEp/MZpt5DQVxpIEWkGg9q6p5vdDOwKFLFTBNuOQ6NzD3ZMLalb
cxXb2nqp4w6uRcwoFof/u2Z3s87bnllfAAXI6cSX4uY5/JPudsfF7LM+YR6hsab5
IymZqshtKxQwv8DByYXIKeNFS0xsc9zpqbZLPELvbMZ7foMUZR/pwO/VURsW5k2W
ucLjF2X36CGHdeypU2s7NSCtRSyGfRWf0aZOclzPdRk9xZNrz1kjgMPjlsaFErq0
2pHxPBic+/4lVGqZiOPPHLZ10POiAalApZ2gCOnOdm5MxpWhSu+1+mgut+9Rc9cB
W8A4JHlb/GgRBetfM2fiyDLQCW+HUCVXJ4rCWfbUPu8xiHtJDEVURByqW7R2rJ80
YLx67FKZe/13IiNFEJKlFsTox3oYgVFNmH7eGsta/qiB+3oo8aBgdS+pdiLt3OL6
Q098gUrYKjJh7Do9oLOwSaJx0JDMAW1H9FGDt5JcGMLwP3c9+TsH8YfoHBxO1wZT
0yM8Mklvq1tJ9fEWO2ab+6TllJR0QxCU45SeQBi5KPRR/UsI0yAUxZHGGQiFUZ45
jOs8cIJ3sykQJ5bD4O4BcJYPg0Dq8s+6r/vgtjNA4t9rpf01ICJoEAksJWinvZ8n
El+8nGHxiQnYm7cJ34e0LcjTH2LdliSgqxE08tDiMrWJ+y6wdqykDOB9S7v6qiid
T33yTLpv+PnbOSbCaelNR9daXlJryaYJxEs39biQm/rrJOWpkkXE6sbG16rnEFWr
rOI2LJxq1upJtyTxSNhQBOBqed4HGfifq7kQHJLhjqqqH4dQbhedF3aqANCnKUdE
9HKdNEaXlnFHxouD9Ty2SR1pDzhbSosCNN4wUaBVtSbxtb0AMamSNEkjy+TCT6L5
oZagPucbOhQNb/HIhhMPTt9/tJ2xDOd3ErR9Wgc4ZokKIt7Ni7KhMmjVxRUpQDIg
BM3HMPFSOj0pDXAEP1LZhANACTsDU4tyGr9/sUMiMPf3Oure0PYxeWPrucPyTuFy
YuCraHiyiJNmZgKjixbHJt0Y1osmShe6hz0Z9+GLk11he4a81Esp3YVRlziGb//Y
jVGJWyNaJMw/CLRMJVsnsGz1QwzU2ofsWIRw6B7d81d/IrbRO+rRJTSpo5JoXcxI
ZFm8R8tO+nNmY9HaY1da1OABpG2u2IlBW7mJBNJ2RWamJHwKvXn0RKJ4QPoNAOkq
exAyLjRO2PgbfttLhwprksa0RPB9l8xKiM+DwKsbCi8Ajt0iCld4M8MtNC+tMJd+
c/bP6SmWwftQeMpjCjFdd/rMEsPfphNuGCKdd1FUbUAUBdGuu6Fqza72NoewOdeV
d2dxd7OIjfX5KHKuF2OCMDKbDDNW4JHF0mscixpvj6FADRZaJvqXd+8yCeQ3z512
58Q8oPJrGxR/aX8nFPLlBFFozpRHgm87ykRp5y0ph2YXrt3i4NoK0aAl7SxGRzdp
EY0NLsQlLBiWlVuYYMoKCOMQTu2gHeSaRJeFsQG+GHmLWXuStT+9JFTbxIPUFILA
3JE+LBCm++oh440BzZiKR97/gEKcR7aOliho8k7NcByukPj2pvhsd4mEe6jySjVo
5xthvXRR+YrGKfJfbSl+Ox4RrilgkmJZ7JMecAi2AVn9ijmD7KpK7/be5f5aKrQM
eNc+0DBu70sL2jSCSSIhhPMldoZT8V7JWZHx3U+3melyI3vsyy/1sbG6xM6M7i1f
sKDxfHe2MwwBw0bOZTqX69uMI3E5ubrp/IHtC3Fhs7Vio+lEZPlVdPA1TOueASWU
gV5JjWZ5F/aaYvXM6tTtssTulPl3+nx4ypqOgctOIUmfYyvYHgIHCEoXXTAX1teF
PhxMTuB7XnIY/VxwLnONhbXQhqFGls8EV6K0A0DkF1OEcvjk+gYKecAxJImy7oSV
O1lXRWfsxiMDFRlg6JhvfiJmV2gHkzs0ruRZ4x/suPROwmc7w9gPIe3DbwN6tXPU
A7/1DuIlPEh89vakveO7uBX+D0vzCvdPbms3Xi2qdWS9Ycv6y1iOwLZJYVOG4g/p
H4rUm8yOhsoxkpGVEVRqT7MdTgbmqIYFidkApA9rwlTtfS4UV070/pleT2zQZWZ/
+bxiAMKL4SJMibppRx+CB1BXFrYJAf3ctlNBopg003trGeYcU/8WTBELINwKDuve
KVqunVbi2o7wPqmJujdcCyAR3yvavv0YI75y2vyYh3cXIegrn9QJzaXzJuj1b/2X
bjpwVUToXhp+yM1GXMcE0SQ44KcxLCObPO83GWSlylCbowNUoToFrtrjGzmRpXnm
UtdJ9voY9W1TKls8gE2PwyoQa/Dj9ItMrGYa38CQWV9uOqWL3DE8xxhOngdG1xv0
65j76anjrkMl7rhGlB5GVOABWvGox0NDH+HqWAz+Ti5eBm+uO6oqld1moa+FPPkt
IaMf9oPZ120xfTYUxTGlILpXhrDjjuw+kiG0ZhxxOhXoVzKSx0FTQfW6wu5Xyu2I
gmeFsFE2Y2uenP8BJUn1Kyrckrw604KcyKkW5Fle5YmGopMgEzPpQSnI5YBl6UlW
07O9R03Ck+rZY3/2yNlIgstz81anPx6/EhezbFNVHqNen3w9oRWhot+/sN2wN/Sk
MhRZC2Bb70ClpGBWJ7jZjaVOYz/fZ7Yv1AEXfReQOAiQfBigm51USmNvdxUeWwJi
P41X8vHvwOrFAPU7kGZEUfm+6khIJVlUMNKLm9THRS6Kh3fq8JL1fZvyaYGJBaqL
5rzdkX4pSqUOeVzYHSRQr1DCcJRsIo+ulXgD6dhpWcqkHUcXd5MtlgNLF1f3GwSY
E7y9Lc6zldZGTOObvLBlifh1qDGm/n/FVxlObHCt6IfIMCSngf0iV+oSjLCrFvKo
fKiTNRCDQyCUwYv270VMYmk4+9bgK6/r5ZxxY94B0zHRlFtC1Yf0aaMR7Bxqm5q7
JI8yAJzqEy1RqIidIcsb59vl14Fq41Da2CsZYFfP8c2EGq6COS2yP68nkW8277e9
29D5BrAVuuMylXFV8oVEf3cNaq+iHJXbetuYhIyBqcI1On7WNCOMTPvOvONnKwVw
vPCdVeLLsl3mmCm7VKU8PPAPH8mkP7Ur3jvWvNQhGogXppK1cX0o7HYKD7YXjRci
3MALsanXVVzLU0VPEZLVLWlnZ0KqFVRvqNQfB6+cAM9GIDVdt16k95WD+InIz5Fo
DvtmFhGYJ6fZuSgLx31UHlsA1s/1Ih0t5GSJCmAj3eYqt8GA+YitiE+DtSF6WQit
bPfQHR1lZPa5ea1KF+yTSO0kTiDIE1X7wi4ofKFRWNZI9cGKQ1fMJ54b4xvdJPJ1
YycCTwnXna/IFlx/GlshMG8N15YVj7qyhQkqoaVAwV9Dj14vujTqA8DUdLrSXnMO
CVR5u3IK8OiOVeqi53+NV0xbtD85ohlspj4GhPVIKyoiFSgNU7agVeFKNjoV8ovD
tH2BdLuZgEKES08SylSTcy6GxDyKdPBv2DFJ3DzTBuFYJkF/Ytgp5JKGk37gaQiC
V5pPwBjjgLycMzcpZyUp3NusnJKzyWoYUN6wSxxehyRYI5rioPej+6oHQ5P0OSQG
borZ2w7r9DnAnxbwE4BKxWAJi/RoXcpGOF2hRBzrs/tzBFg7NojgRcT+S68lSyJB
ht7+2Aodu1jthRLfMpj3Gk/OAbah9TgxhIdLVn0APVzG/edwN8W3O5SyvavBJmXG
90T9PdbFSSHWVWpLty1YANTlqQfrfY9H3Y81dhx3Yy0qnRa4cndLliAMwmQt63aL
l2Cc8R8Rcz9JYow2pT8P6yB1wXiUf1+qlNSt3ExJ8klTnln+DJIDiqQUvAkxShGI
uiTT8sKhMCl8RBBAJL6pfIubiwudGYaSpEV8YJTvNClYJVtswxo/QapTyE+yas2t
I5HXqGls/QzwxnFcUq7cfEFFWpL0ywR8SntjoFuAND/UKwdhHVxaxoKCGWFpIBvH
gFxBtLnjsb26qFjhURbUijgQ4gIaiFQWRnxk1kz+xTcd6aslzu5zdnsf90fgP8qy
F6HdBizYdUYPmBsgiUqX0tjsb86mrsR1wtekh8uS8LsYoEvlgywwr9fA/i+PoKkf
m/SXXgzO3WVYszWxdatJ8upF0WeO/zNgua/qInbcx7bcYR4RxVQQVxRPaph3e//c
wm5ObeZ6ZUo8evKXIJ4nSxcrqloNYsGWX5iaXFE5fDnXvwsoW/qVhCizqdwZG/NY
jqZHJvPvpLRZ45rc0gI4wKdWA1cj/wM2y8HDbq8S4hYvm+wNqbFjSNZJgL8Nz9Qs
DJxXSe6wkvETIWk68VdciIVtDzGELDP2Gb4HwDgsvCT5vEBGCY5uoiPkMsrBvQ05
yK4IYJIZsukVQaqHE7MTgRD6F5Fpmby/kz8S234kp1gL76IqUn/wbARvkuPJGLHt
uPGXggKNlU9ekMt/L5dRcNW9ZTDYZTnKwGHBX3Y6vpcRYzJNoFD92K2/3TLN05uJ
Ltup248Lv33JmmoHKN+fTmVOKW8vEBMpqe7X0KZ/qC91OnRqD52UPYkAmK37iZNt
Uf6xHl31HHl0dYO1lDPPPU/c3u0R0zUo7KNfYI7xs8iE1WuqfHFFxqMEBVYOvIW6
6MpaAdY/G3LGrhaIBJwp/Rz9SvpCCGNucGkjh604+ynWZWU5RDM/jn9VZhZKgBS7
UmbgSir9XcnLY/2Vn78muTCimYJV6C9v5SJSeU6o7i5259GFbwI9Miytj90Q5YVd
OvqFRy5PjrDb4I1M0d7H5+T+L60RoeOxXeJL/k//XGPqEPAbvL5K3W5o7pSgYPby
esz2PJCMHpMERmzsw6WKcfX3ePOL0xA+2CX4ZE09xn3yFc24WhIKIeCDqIzwlv1C
b6w8MZ5apXn1KTX2woyjsgPIIHeqdVr2UCqZ66Bk7DMVMVrhCPpeNVT8hn3p40rR
uoiete+3DqobD8kkoN4Tv3aQmhiFXH4SUpzL56JlgMgBuyJtPMMZAKHGUlwfkFOA
RfShJ81LgtUsdV6i4tFGqD5uKJ7E78LOcsXvxLU/kfMcqb61A45t5Jkcfe2MJ8O6
kviQ2rtDQQi20OhAzCP9xA01rHxRpc60K/7vOpVCeyo4y5bSRDxBi2AXahEtOg+Z
Mn6PrwFeAYYIhcwyMfBJgU4okeRQFygcZyGEXnQolgzhfCup1PNlJNybtKCUgUK+
dAp5lAvZLKdak2vs4Des/kzedEq+lCmfg9i5JB1rbZzvybnoazqQ18oynV/lu/zW
Ruh23ZhWInPe0DACxlt8HoKo1qzK0TWZpm7vsvCiqiCoB1Ie7QT7wOc/zd8s4OGo
4zQbK3mmuecP4TRAyWSpIl2s1vAZhiqIxFUg5wuDe7Ua3iYXAFZLq2lVHmrR4JOH
rXNEGtib7hchTpJlQh3gVLNxWWwJnBG7s9vlcxYQTSNP9/fW4HM3bW+4fy/jpteP
MS+4wOMhUONKt22miNRrx4ZAZmaLhgaWCPHLqkmR0EAJfgqwTaV6ugWKLv0LbG+E
zIx1vMZQc9X5K0tc9rYV6i9jFchLJlDXemUyrqGW07q2LWj8W9F7A6rQlOKWkB7Y
PGXnzgu76Lx7i7BICsWOyrm2HyP7DQOb6xeRyebrfTK6JZLFTuZ+VIG8rewDFn23
QrHIbfj3PIC/JXT9b07ImKhD/nBducQld31yzBMxjZ3u+4QgbP0gn9k1Sk6DGdYc
p471LPpPWZelRw/tqgVj78tvn47PWnrCCXLa1zf8KXb6ZGw0pspK9QXB0/EhbxsF
ULTvgXHBeQkNMoEzDD1GPWKnrWsx+Hll9qTfmvu7Tjf4NPGwluwJ00jnSHeFLp7q
m7/91H7SxBoqS5sebUuzswVYf8I2QXvivTLpqML4QF7PWzjNtNxb9q5U7T6zH2N1
wJL5WMxtfgyatYqoUWsR1oBwaMs9xGR68/TR0ua6lk29wzZx1mh2rS59rZGFWF7F
UvcjXCVOERQVF44H+fjIuQdTBAqGmHMTnoXTVgnWgRCPUEETY6mtTTVHb2F6icAV
eXv7hnvvAgzmnGC4jYz/rlgJmVx9IRUDArQqcdiGGqIaWal51GCNtjB0EVWNaswp
MeVxY9dCJRhkS78UlTIhnDid2g6ySNDouN+OUjuigf/WKSoqqDc+NEvJnP0dCANU
eCP4PRlWE62xjuTs8Qc6jht+xniS6aznlMxGPx0gx7bSREYuIaS9ye8B8JiugEpR
HnTw9SurKuMgYUDwAiIMGPfA38Gc93TCAxP5DA0znjGUVZQ2+9I73hCf1/5tJXxC
a5QeIZr5ODcEuZEfRwi250rEoa0xFcQ+wDzu1idsD6Z1t1qoheustnY5pY4gHdb0
uq8lKz7aP7SAiwwR/FOttAMKy3WnSQcc/U698NcFXdPGP9v0vLglb6rXEbxQyRY5
nWz3JpvAhxWHw7gqTnFpR4TUsPInte7h3Q5aKPw6e0034BZsY9KAZOdp+XeiHyxF
YfyU78iwIVAumo0APRq0Yd5ttNbSN8NHrE28SVu8A9vmxQi3/rZFFxMeFI2DLwen
JcTjKUJE7hCL3MFeHnLUNNRmR5x1B/91bq3IJ+W8zZN9gfJfpq0XUKMgG5e+h9ls
Qeg6QWsUOb+6gB+XHYHXo9AtoltL/mzB25vOhnVxetgPb1jNHS0I9EVCZ7mqdlpA
bSHMvMz3q2P7mpDsjP1Zy5XX552fZ69KKBY/uMUesGWM0iqvzw2DYoPv0VHM9t3T
AH5AK/by5nbPjeGkEheofs1x9hFarcKk+fLRSdwIJGC+Ns1LUfsOO7YbWNHdB97t
7oONc0631Gxc99JpNxitL/wEeaWGt/CXRyZgyWZbFQHHTjLryzsMlxiXL5j2GfTX
7P2tnUK7hwsmgmrxoeeNaIIKpKqVvlqliokYpH/HWlnc0Wrr6b3PrBHQI1lAnLh+
nHUAnLTxWYjcCm2dGEnD6DT9cn/cpw4bXwffo2juDbZZM+ehvoP+Wnwyl99LG1cK
JPMYuIkK+A8Mcyl0ulKwyYkfR7UIxaSWU+LfQmHYq+cil77Q7tSC6wE64ch3cESF
EQaNHJRF9kQ4e3MT6iAkwH85zThf2YqSF1wzKhH85a9D0gOvKGVp+fNU2BsUOMy7
5Z0O/U0J/POnJM3ylVzvSKbRXr7H9RpHWmecqr34aXMuGIVkL1X2fe+TLx+pMZwz
JcGf9yHB51gCKRZax9AHrHyrQHoj2hbLcUgKmGK0BhY56NEHSDavfGsFdvgcoNMe
74YukcKCpNFxulb1fz4q/8fTwWli1D5aEvauCj8qYCyDG1BL7C8CTp6eK55KRikr
d9sDcO6NFNxJ5AqDnH78w8BAaPEEkmJPnANg7wAVeWogX6phsRKd86pE83GXenPx
N1LX4zlqFR5W5i+zjmdvzzAboTpigkLG7ZsyJEkgrVC0oarmfwQABfVU7oHWRFaX
1d9vP4zXSbg/rxejX8AaYF3r1P7F8Myddc8wW3WFVLNHj5bCEjBj03IvImJf06dY
0ZYMMm6wGAzaRzV3pWqKHbW7EV2+kqzfuIuo2BKANKJqvBFbgsuHquvUinm9Qykv
Y2x6jp2uTnsgBqIvF2QpQ4SiI1opMwplwjpeN6sgNA2S4acN+SdJaaqYslm6PBbF
1BRrgjYR9pUMhxXD32U5biQW4e+xSIHHdDOI5vv4XMI12cFbug9/zGcb1ng0VgR6
dR7ohD2J/US9Wj6cpS59qmimAdVWyPdZrg19VMZ+hh9j6pnLYJaw5t5ILYlPIeoe
E1Ap+EooWWik+9EBjDHWq1g9c/AMsqVIe93VaemSaeXSJJw+tYU0W+1EttqnSbgN
PKZctZ8EcU/yWSfIPt5NwdYp80LlEyHFsgQz/uAPMDc2HFIWyBKmfXdbm5AfVRAZ
8AwkgkDWsuHyU8Z5f2JbTRHwevARd6ANsnXwa9aqSw1NGzTCnxPiRIMcUa6SfoOX
+9pXmIKSnRP6ZvE3lnn763FAIKs0RwCVa8Cu5hdNbzeaMt8Lz+9IFBXwAvIxtUOY
4yX38X3j1Xc3tjGUEs+S1IAlA8jFRkNGhWDWCN1h/MPxktfBJ261JBVLZOF+Wu7p
pyyJIbZ0vxrDfn4uOl0ryOKzs+TaYYP/jOnmHYtFTLLNeFK/Wy6hjAe70UkGWHB2
UEXVdk8TQGJOVLHqd/yxghrKBqUjLBQjBnCqU255LbIRAWmyzyta6qQC0XBm4++n
LAtnIv1IAqPJrWL56HXBcVOSh8EqtQ1Baj1spQ1rd/miDsLKmlbRrnN4Io9I5E99
rMMmuCzmTbaVLfcqkGqZewSHcB2Grqe2xMWyMQch3xXLwsorZNX9tcwzXDmC2O6/
IivqvZbM6nUafDwLZhZk7ihvA0T9EyDDRLzZILsIfT0WMh94JuhlV2fTqXPBl1tn
FrC8rR4VVkTc/uq8nplevMroWRXiXdxiwlpiwJiuxwxf4vZDVnhb09WCm6ZFNtLo
/aT7E5uQDIjvXhalnD916a/VN3U3ntGLcRdcT0Jr144qHLhPCNNxFOWLwbGcfRrt
LIGPd3XS2foO6qpbd4kzURE+ChdVNKDvrp264VmOkFHE3Sohp/+EC8Zmrm+Bd4xw
rAznUph3BJi9SCIsiFFUMDhbb9SHvJ8/v0le8vfRRDTylsYd8frssTJfyferMVaj
rllOWkbWIpfdmzptp6J9eLHbNJTgJaOp/YClFRRZwbrB/YIJQtB4uRo9BmosHct+
kqlk7a9rKDLRm5SE4fRu2oDXjk47/x/p7NUKmoG70tMu2zRI/wFD5/3oNlXHm01f
KTQpEs97lGSVdSOQceRincBhn5b6YeW5UYUYT1VwBfSkgXKuxAXOTp5xIAmCbhNI
4hxIhrSDLapx3XDHy4yGDKs6UYXZu2R1A7iaHde0f7CT9YPJq5j5YthPjTjdCjaJ
KhQsOmSXs0x5BYxjJynPKIuDKJEBvXH5xLdRamw1YrI6AUn3wj6xCGWXsngaTfly
Ab4XTALh8tyNWJ0xyVNKRSAxTx0wc4lbtPcMh7IMOLT4PRLa0UlLJ5LOd0v3UC8q
YIflS3hUOYSxvus9hxFOsSxDNuEwSaZ89CfyP/QyORUUS9Y43lAwRDItwJEZ21pi
mTyfqkgU73mx28s/2lVTtMHMdxD9gavxAREvKSea7+8yUCbjv2ryJcQQtH3TkvKS
uBOXfkKFDy9kyj9T1wfOSNGm0FDmwei0BaIvE60ArhXeZ/n/rDZW8VVl420Bt3s8
cNBeZZCnJwCGfRHcv7UlX5s62fJw2v6ZcVFbsW4KGHjwXdMfI8lbCRORe+RZWcHc
XxeMh/MyA4U+ZOsUYDhA7GMj1TUezzsgKVD2UM/Dn359mFuDClJ7voVbtQs2wkHZ
5G+1CyQMwXq+5ixH49gW1SeepoCxGbwy3SHiGK5FZd53Uul9uxnGgdiFkGTpz9s8
X1/2TnMW2l4wvWwBu/ILxG2214TYbcUiyGkRHV5irMN0JuEw5Tqxj66gHXJk5l9P
U7MvjZWSxp7XBebWxraV14ROLs6MwIsdUhf7kIS7ENeGJad++IvFQupZu3lfmKzD
bzPMsfBjBFR71s53+xjFV7WrsK+A1AO1l+wRCP0dNfUDoUMMWMDsIRNeaGRApOWK
DocmQvWStL3jUpcDttqOTbH/J19XBpr3ORi4p3iElRfE8twrp1952u9B0plkdS7l
1dmqpJ0/wJbdTzZCQ7uV4MN3cXO8XuLzpGVXIy+E0A3+9Ia8q+il4yK+NqsrJCg6
FpRl1Hp6aLpRMxw+JjJdq0+WELrZTjdRPAy7NM5946tp2+X3xblol9aGbNP/63mU
cmPeeMMpkq6LaA0NVqEQyqHOiKEFh2q7yIkQH8rP/8Wgs+46Xmb3nyEoTvn+FVKX
eVq1pNAW3QQk7O1jXIiCHJoLPsXrIa+iKOJc1zGwgBl9hLTxCocc1kaQ69CAWu05
MLjVQ8WgRmcUNjmbKw+Wa6nsaR4vFqxAOP/I3NoLcFfq4nsMsFhcu3n1M8zAQmDT
0jedKIfd++t4bOQ8El3X9rOQQA1Ol4PiEtwAyOXPaUdD0BK6IBIBV4hqANLalD3q
xqrS2qUpcurHCf+TgityfMsEMfQyGJGxPT+OfbN1Nf7LY7u4qUFWGYX8kM48mV6e
x/eJ5hB/dFxeuiwW4JCijD5HTDF+ewdEb+aYVXBUQyU/yr/oq1KkllwtPTv6E5RL
IkH9gFX4L1rGSRRo1WLvp/NH7HmuiZBPMevr1Mm6hwuz2GUSCDDz0B+b9u1wzaPj
chA8XH6xV9y72dpg/hD/pD0aOy1Hp3IFaaNhEiR+x10FJjtDYkLLpVIwYwGy72rF
SWh32IXUia0PLAfQXl7u8vSnbZlpad2WBvFW9k6WTdA4chOWZ4mlgoDbfczWWjgn
2+1f/u0a80I5uxQIuc29vauirLVCyXuHsciV0gB3FWV5iE++e7X32OzPKEFjc5Es
I8mGhPjWLfv6vGYJuuMeNwV0+mnUuUVFx4YE6Y7kD2QPbQWJzHpBtF0EkyHp0lEj
zx/OxhJ7z5/DpRNuTLpUqkErCNSHyunRvI0rh9JxkzyHtCAVPUv2dIf1XxpLEFVE
tYceLxYhcB0p9cbR+o2xJEvtDPOAHC+/FTEZs4/9utGGKFJzwBVwRUmCFqKvDG0/
DdRJzKlmGlLsB7swLGUsVd7b3kFpZtJOdpkd3Jvp4BrsttFmCh7acJriIC+35iK6
d6OasRjlc5jABc9pvJo49cqRmdYh6yXq7sRnM4dtLhf7UBdHKoazS2RRTC8qhViO
8YHw0CHmND2MjDp9v5nIeDJxAF62acG6zYJ75qZEfKyKbVFIKvFINonLE1SJG/es
X/Zi6clufZc/8n4Zti5zxKf+KajsSXAlI6ea9hCGtY6RJf/gY8F/OydDDa8hbHXw
dWprN3hm0VabEEcHqIj29bf4NxWxYt8EcVUzsiAHgY6wA39U2is7XWfsWPMZgruz
F6FhhP9CB6ekpw29C896iy4GvwIjpozyDCE02ewvEv67yNJ50Z42nPsD+sF77bx0
+WXaPPB5siKtouJAFfdPaujoL/MrIJIGD74YgtGT0zOXn614vPN0vp31ta7zwYQE
2w+yrJBP0UaPX3YtAhBDRNCXYrbP2VL88UTR09iD+BGxJL9UPW2k6jiTwTfxvJmm
27KDhg+s/QHhxLtMbq3ja2muh4aTzEaDm6qFDU7UnXQ92SR8/oq2N3uq8r0EFZMK
oA72RXJCvTr9FVHs/Y1vzfhqKfpYYtrWY4QuXE3FER3R0uXRAG8mKuzeNLY739Dp
3GE6xLuI200p4pVOMawghVopOqqvVXvxVp0kIdnm/xbtK/tErKH06U70FvToVnC6
sWYLlRpVvn8AdGHu/R7vrSKs9NuMPSoR2rKpd5MIX/DScA1fszlgDP1pTVmK+VAE
pPGvfrXEXbfgRVI3KQiTdwOePXOaTCcgIoRlnY3haqrMyYne4L10wSPseUkgG0/f
i+77CbTMSzprbFLKit4t+qAIs6eCZO9XXa3Dytk3wRHdDL1ZHQJv1TaxBfQydOCv
kiF2Eo5M1BvuvUVSuDgEKQw+moaIaMiN1Ubo3isnJzmt3XDUp6Axuvo8hiTfOInR
fGCuNzuX9wsqESVUAgmUzrir8jcgRtK30adeRnM7kcNs6IHoW3RBICOhCzHoZ4EO
Qnn2Bd+CIbvOV499V7EXehegRkUB96LNs+UmVTGoFnoja3D0Ck+RC3SGuzXu76Bh
lZKUtMDJ36OZCL6E5YoXXT8Nuv5HjHVegthWkFOb/TeMjTxvjZC0T2BQuk+UqIdV
LhCzW6HMdPkHILmBgB8T118v4gCTbsqN+2NWhZeRVS8DpYXY7JkxS/Hg75oqlq2Z
SZM9z18x4/q/2oniD5QtkE+1Z9NtMIxOcUoK8HAGMTm1mrv+V2ku/3ENFoctKIQ5
qALTaD9+8B21SCPjqJG9NZ/L4/ia86R1BwIKaE6poMG+okCNZpoFZ27U2GrTEszP
9U+J6lAwHFrw38b5nXTchXvw2PJR4RP56bk/sdMPAzWqdD955maXV7Ue+IAoBqpO
ALAOcAXFHpr3LL+3sH8WtjIng6+lA0D/0fbjD7KKE+Ut7xUOUFnYO5H9L+RzzeVn
SPDkg06Amp6SGZqzsWGhWFqpEbsXH3f1fD88OxVFvBieAQGeoK8XsTLhtRkFAGqf
MhNWM71/p2QMDVqnzKbd8TimKVGRstnoRRditzMyK8aZecO6qCnbLo8b3AO5Ha0U
/ORMT1nhWw04FlresmwDF+Oxdcq4YyybgICmlaABKqN49sEymV6BxR5JGlrMKaw9
bE7jrKh3Y2MWNx6kaLcKUlc8OUs9FgQ+V0IqKJ+lXmkW5m8QyZC53zitr3NBzJhJ
HJuWsl1QisZQ0x4a9oFQYOiUgdvvYF4DqfMDjWZjIT9gJ9XtsAd2Ujj0DFmW/NF7
oUbl5+crLu8HyAremo6zRdoefsU27y62jJ0WwJ5khrbZ1ildfn6x9d9P4KqeRJul
kKLMzbE9B/HIzdKIJ5CO/+FLzj1/oyiJFCF7o9AusaSzm90N+Kq26B2hLMWE1YDn
srft35tggVmOtUwO82IWXkEIgZs/olIGVpSH5DJLdinXsMmmcrICYoFlEkWMJxny
07wRfIbn+inGp1V5FQF2tMonWRZMyc50/FZjdkgXo4XcHZijqvDxswEpg68pgHsi
y6A28CYmG0lsPwK4ZwhvFwYAn4RfragAQfG9Y9Cz3JllRDsDd7RaMO7EoOZF+amK
4gChSa5/LFvbC3PxgeyP3yeFKX5lXytYGy+RKX/hNp+x4s68KYMdqGTROF05+NSr
9npoPdRcfV+hf/1+gg6ALtoDwJV+WBLhSE/3ehNKBrZEPy0WdsEv7AkU9RGgDOGa
oaaQHVWDUZqGPCkCZDiH2BOq4L4rfEgglKFVuRFT8on42oJJSyeX6N3hMuEb0bew
2EL5q669I9US4MoFDw9uMsJHekQdcaO787yQZvgEmLcmcM8f2rG1RNNp0f9WJR/h
GW7gXZbNdeLv6KSiU0x8jbhSaNeQdUdzIlzZgYYbplzjkSo65ACbGJV4opEta8xM
XZ/IxC0+LT99mIORBSz8gmOlP+8XLPdyR0Sa51TtvjoKj49wh4jRksEvlhnYrbU8
AjxSIZkWoUg1tpKX5Ncypk/Hx0gCyiikn38Wn52TtJ6RpoEUbpvV1DAZj8esXB9K
2uTkewezCwv9PUgbVoVjV4FoKbsMmTONEY34c5P9Js1BBrNSqsgLeGudhvYGiXpy
f20m++f+7ppdjJcuk/Lm0P3ZS5lhitQXB+Ic+330j0vD5/+fYHhjDmAEWe8I8Z/J
yaESTSJv6y+kcbVFb12guV4c9m8G2an5yzge9F5NgQa8ewzCIiYAfCPST/fpb01U
GPSZuNdseaR970RI5LvitIzRk5N2J5LAV1eXFZ55g0E6nf9Qg/esV1OHnoB+y52K
FDTOZzUZEEX0j8Y7a0Z/1EhF2OnkthUtXMcU67/BnVnQxbhVjkDr9HWnKQC2jRF8
EyOo+ygl+Zg62CiFpKsEJqAqtCSzqo1/X7ulpK7mPuQSEuUfQ4agdetpjZNqzyQO
ChdCIysnuqZfKQXFFyyjXTbXN0yQntRhE3QVg/Y0xzF3MdghtUMqW4J7SIjziZVg
Zcs2REefyDK+puwRb152lSO1fwoAQdR4XVg0ewfOFJu+0FZet/OOEFaoFSCbpJaM
GgoOeG5YLeZa/pYFqI62ymyWWCc972/n7HCnxNYvMxIP0M0KEPepeADEULpAjBkG
3diJ2qe6+UJ5UQXmzpZHnFtn8Q1bRSfSt/sAKXQirjIPWxcbPVrngeu5N7AfHS5/
MR1pH7arFijBvLTAcH8lF7Y84ypxAhQbgfXgXBiRDgOteJgiXKEibJR+JeCSOmKc
lNQhWcZc4eY2JWbMATKZlu7dqCGpdD3UhxCFMZyiADDt7lHn95hMH6y0oJfr6pUi
7BcLT3KoVk1WdhWMNtK4lRRL4x6vBfgDsH348yAeeIavAUZlrYe5IsJVCdu/FF06
FYdNyfH7EzBrRLg2Olpirw2341RSDKKS8eMaZEOGt3nxY4iTjNhwbiLOhSgM8V6p
8cvP4GYVHItOUM8j0XFwXUC9dRkUMm0BpUkQZhwof9u9NcIeWm/EloROVZaQ25nv
XCyRltcjN2kU5a+PbNyYWPnHpHMtY5ByFZPbdJD2PLc3QDuzDaSfL91uFRy7+EMO
8wsvW6Z7n+lnMcCKF/jLDZtd/EeMdnx6gGFAoNTXcINUXQghJoZBkYfRa2LSE0kS
ihlqf9uCjyulv1IZfwbnFZEctL4oxynqJPEJssnntLmRwiRKe6xjCUCaJCoHahCK
mwAT8w5kOUCKC3vzq+eNubXeYH0b2t0InAg7PcfDlamNwcknkknl7E5OW6ftjN0K
Vopun2JqlQl6ag5OGeP3uwifWKZq6CP7phvjBkO0KHemEb+l7tQCuDCttj7rCcwK
ZhUyjwbuG3/efbN4Aybsbp9VN6zYeqEHgG8GTgBXEgtWLy6Aaj3IpVfWJTXDgqJG
pRz76JRy43+ZwaN9t3seZ1ku7bCPiFIrYhp9hl5dnBaj7yPWu7/BqMfP3UZjUco+
1aAKYTTKSXR0JWX3gyUrQ7+tVwdGLhK0bENneI5p/pFbiAnTBOFkR5zte38HUPHQ
/Jk3tQ3hIjPArl9dZBNn7lyjqiye3AGQZn9moozU3MEPssEhHg0Yo9hjYEp3fC1p
nAVsLrjnzvQ9iCGClqXintHElGQtxEGknk7y/hRxkZMGGqXJV1xpa89GzBrUq+BU
PHyK2Uv997/NwQlyKnTxO4RkzHuuZHTV6TzujTL93wu1qXpfDZbRN7cKgLIymyGE
AVqagsiesdOGVw//T6DXZi9c0PODj63eIYWjuC1aSyrPLQzeq5MkFIIOFI7YQim3
3rAe5I4095Ut+0IcU6a/2fPkMmsvQ2rgnbjM2UH8JCI2l9iwzw+j7/F1CoDEUCia
s/bjB8Q4rOXNdrEldStfQRYtXfYY7MLmysWiPBS9HyjcoWvIsCVeWiilQWNUYxAj
6n+GBUGA1MzcDSUlzC7YDh4doEC8KVQfXThR8jxiyxwt0+xyCb9yL8nsc2/ImaSg
yX8OOaMRGBWGZ1c/0BbA4vQZKTltXAjX0EJOSCCPMQrwQYaIkl3bEQjHV+khyEaW
5cqofuSkPvhGQ4SvdzGQasYxYZC5fHBajx4OxxZ4Pi3ad1GDtvudPh1rG+cFZ6UP
DDmH5sRk6I7OzTUkOb71CuK1iY77hNFNhXIW7m8EBTniuX94AKWxNhPSBRDIak/U
gSI4kc3ej2iehy9yv/cYJC3nwg721HtuiPPqihcqrSjyDFC1iOjOsN8OE/97+ZQc
e9KAGnxzKXdnmLb6VZyP5phPM317yWRCfEVRG69bYu5ycwESTRWesaeaxqG7U4fQ
/cgk1V9BTEFIMa1G75bdIr/NvLdFU33btbTiJ1QS9BQ0JelSf+uoW81stMKjnF4w
Qu8e+vI2JITeMjo3NqYaQkFIW1MB4x5TaE7B1EVq/l6XCkpnhbPUaQRyWcgcI1uY
jPiPk9rwL/8d1ev5M7foDOju5/l5F92CJ3U2zw6FXK9TQG1/bfhPnAsvXAfLm/er
2Fgr4OtuEnGIxbBAU543FkW4iE60QLH7+X+Yp83DAaW7KuSAcxkjdvSqhZOpXNIJ
ctKZxCWu4KUVzH49rklZCr3Qdp5YWyyyppbo1Iqow6tjrj32S8jPlGZUBLu++3WK
UvnRqZwkeCHDfCLZ7+yZx1/ybH9HrN3ufcBAgUR4xlKoiFReXfF0SDWm5wgR9Mxh
8q8zD1H+GEvzmWlYNKtJ3oQUcYpbB5f6IlgSQNCKEVs6pc3tTp7ZqEOI+M0U7RXP
JusjmjlJxWZCqQHbzj1dPn3vGc4krEmlEMSU3Oh20iq3EAVeSazgq4NEI86A+u2U
8NekkqreFosMYUH921PfdHkI51QDf20pvU3MCOzNnciel5Fl6LrdTPPTxNn5rGQZ
cYAsSKFo5TiPoHX/Im3QNoxfFAe+khrbPmGr1PSKYpFXHeV2k1RQaRl+wxUSzm4i
30YRyLU3CVOV4uymiVO8ptXpB6S4NSkPi5MscHJDCO/n8GeSK0I5vAwDfF0/EFZN
DJ5sZd0T2SEp/tuQVCrHBghlRG2uROqCeR4zoRvc12jICw5tYQX+PPwUzV1W61To
BHN6j3j1HaUxKlKgApJtgDa8KRWHil1yXRmhoJ6ZQ9+Tq4mFVRf7hu5Oa1Hkwgyn
bZkkPuahsO06EPSVKwHBvrhBvwPsoDgxnn6LPzEqZkW5/uWu233HldONf9u8T5nz
/guClUGTQYVSQ5zugvXXXwD1jv9hy7jfKFz3FUUfmbx/6Eiu7pY6BbOzLs+qLdrq
tcorHysD5axRTT5hg10oaFIjSw+t/dPPAjM01zkocN8XC4tUxyyw5l4jOHWJrSu+
CjUmdjbc4wiZiFxgC7nMUVqxY2NAL8wUu3k+r0SBZwDrRr/gqOgP8qvlvBaAt8T3
124WW5crdlGY9NzTjpCnXhbSIxJI82wQ2HyKuB59efdDPxuBLtnfGDOdjkcp12yr
uDbUIT2lX/iErE081psWfJeNwEWIZ9j60QWzHB8pF1p1g8uJlBWdDBI39S+SMddI
09aU2JoWPqPtmJjzguDZrAbZq1+9bGa7PtqHUPxXdfXQKg9plPrVM19n7NHuPsag
NqNhHeAIZKGLiA7wTpl+HMet7xwn68gXn6RE4TaltgiGUUGb7lKEw9to3OpteCqE
9PJHNt68HV8PFrovfBAify7dN73xlDZyouAE9uuo3O5jQDIXpfr7G47S5u5oZBoH
cM8ONZBYQ2jDxIzxGlD660am5l5pk9IG7BGEe9MnrUMhDczq9MnWOqnva++p8yf/
CCnc6HQEXS1vrho2h6qNoeaUCYcy/lXTI4bdqh5JGoGiJR4mZXCPjX4qoq/3C1n+
MHeAmTW7ueliuiuBOFkKFysR0jBKSqYU2fvBx2w3zeoTp9ZoYVcgyRVNcSzJyXn6
jtvFS4YUrHApBLDKpKeSilJ3BqK6VlU4JG3sI40Xonc7wzkah+mnMesJCfNa1eBT
gMhEBGdLKDyBdnjDTSVJZVDHT7yxZVOpD70rN1+g+PQ5njAmMqHgel9WEK/IeBPr
vNTpR58nAVkLNzQb6Urp2SxGGTECMDEWwurIycDk2KMP+u3uErmUNqjUbfvpXwZw
N0uhWrH5BsRLKTxK+Ftf2GIwL1bmVXvZBSyM1+rCfvYYxeLXPSArKUho5NHvpI+o
qY73cLALQwg0cUOFyrZDHtUyB7Qjrga3sv3oMPs2aar+C0ME4K9YgKbQZuuANjCP
sWhQOPWHWZWAQo2SM8FT2uVS7VSdCh52B1I6U629Syq9sOFhHrqKb1iF/sP5Z8fC
kt2ty3AW9WTdxPYx2M9b51097U/N6GcgbpYKhwVo2UNGA0Goy74VUX3JGRY6RhO9
JYgFvMzumHYsTcXaluNLSJ0N9sAZcemdlZs51aCvuBL2GblPcilKawcbqh+sz8L/
np0QaaolGP+g0ZYhArRE/GEBbUbX5T4byyHXx1rNrfQ9/MOlSI2aDi1Y3LUcJxcT
uR5elOFsd5DRYYEai5JVddKFN08I/arWCG8iDk0juaNtZbfT+13ccyb9bPsJpa4p
6QjDtxzBIu79Ac+1hFne8sI2b6utSb7s46qqXtcdcC0G9nrMoYLEDFey8/iX3PhW
ax+XL1HxJqllXjv5MzWo6b1cKAyXqRciVrjXMe6JbQKC+CqfrzQ7U6rcN5KJydbv
XQwQuLfttL5Hl4OwDW3j1NBx5y+4E8IMZ/RtMhAUOLQwj1UMG4ZS/4x88/BEWrKy
8BcgDp9LRwh5C6GYAN6T4dv4ZmAcVpT4HgVHdbGI538XRO2bkjaVESZsO3CB5yZD
c20il1RIPI8DJ+q6MROokHbo1H559C4KDZyDZTmRtzPz7+/i5L88+p2E3C6LI/7y
GEtI32xh5TFTJQQrTmEnspF/eteFkhlhzEgFmluHF5pygwXpJR9Sof0sdvsorQw3
fAa3ptIw+BM21LPq93/AJfcHFJHon1pabyZ0ZDv7zhj9AqkMTpxc+x1RTRXnoZWy
Kd9CTuoeyMVGURHG21uYOZvqQ5LKlC0Q6hbBg8d1+LegtZLCyZEmjn9CPHlE34I7
LqYhiUQayp8pNmBIalBz+FqqkfWSM4c+41gt2nY25u9GvNOfQGf3Xk3YgHL1e2kB
q2YR5RJ0Kl2MMJzeegu4S1J5qS6VZnY2lUgjyvBap5HjloIPJnvhtWxuYfAWNfCH
XjoC4Gd/EDrmcQghEWQheUYt1BUj/G7eQ6jQZFxGRaSknFBbrApbQprX9neTU3wg
BwHa5TT/5be1VHS/K47I5Iv4nia8IIeMXhObY776QG6PW+mxAiWvGwE5CQr//06s
2xgqrF46Yxamm1maWkho88qGnt482pG0clUet71hMfm++h2vohOBodO4feHbZSp0
BEXnjhOanl7bmpXatHAd2a/mOvRbcLh3MRX4+MmTEVygyPifsvK7dQx7VD6qrGSd
Vb7F0efOKn7ImwN7+f2VA1zBoWzf3JHVz1PKB/GzLw6Pq3abFtJXt1LSnadLxuiT
3OpBNGVVY+tx3MMRNx1ATSGdzpIGr/0BA4SUQ4Z4QbLM0t3r253JEcdk/rQkbtKb
r1+ILntU7RghCYdYfFORlpohRzA0T74UEKEpEzSuiFiouR7StdsUk12s8qIVbkiD
EisDKbo7Zk2iNB5vjsiZ6od8yBSrQdwEYLQFyOyhzSGZoVvt9054e10Pd1RlZQlW
w508zFZIz/HtsfHAwvfQA7x7C6qBr0JwOU6IiyiVub+DEfMvkC67m4BQgiKm4NPb
RCTKV3agAn7R9/g5yPSk2E/cwmHaUc7+IwT77nW6vhwff3MQGUsPLTtp05vASnBH
r++DDfAimLbrA/Fvq6k4rdY+Ni9DiFdPVns0PATSTlIVRWL+qxsOuWYTX3slizMm
Qs/Dg+ADLUuxdXWHDU8ifFv0y6n9czwu25U2IYuAq9XExDTNgOUvXZX7caLVZ/80
5PIKuLlz4k9Vozpo9BvDXjtlPLZg7Uv5fXArkA4c7BYclC2mX3nUe7bQkveRuUYQ
uQQS+eEkDDRIu4aSOQnMPiPzfVM8R6UvoQgBMedTkX5XKDRuTO92aSGiYAAL7E7G
Ohse9B5Z1h7i3olVYGWSaz3cQX8Dx2QKTFy9G29wuwOW2O496hPgnhs+Trw/O6wM
cu9V2UJFgUhnl7dLDJ3mQxLdfME5awIySF92uni8Qek3fzvUaWt1t+yVZX2clw/U
E8yUmlWSUM5zwjxsduSMe9OAbNQDGB6/AnbC8WxFiMj+ZyT5pqdGWTGzaKAWAFj8
0FNGXIB03lHvlgoDnffK53HeMjW56bQUO9aaFbB2lCwjnI21Zzn+mUtsjyOQ8VPX
sbYWTYMT9LWBKAFTZjlDpmSw2P/NlzpEwlPaM6HlbXqnnnVPh6Gp9eOAAvkdmgQx
GoaKGBmEc0QsYT+cXQIBCt4apolWTVMtnH9kIyyeUJwlaq/O7sKi3yvSW/Gd1UHO
EVXLn1akIUT9l9d29Yq/izU/X7pKkISUmRT2H6WVqotzx2ecr8cSMfIHDQiAfTRO
0urVnWQgW2bqsKi7L9DwaVCTfML/sVz5BE1C5p+1kg2WJBKy/fsmIPEMft2nRgsH
CRNqj4JNAGIdTgovo9Tcii5EBAo+/vhfqssFARl1fBPTuu8voj3ihcpmg6G6Ujeb
nTODY4hzNkLpwduawBxd3xA3qzUdYHK806tnGW+s7bntcu4Gfzbh5gK2slIdA7th
Q5MYZwHlSL8JHwkNVK9d7f5RsRCfSo/BMbShRdpOjZq0pi7NmB2kzU9A1SZkpXbW
xJxaFmMkrtSuKtl5Zv/U8qnHmgZ+aZ+I23JllTVgmj20UWSt62FfIiwi+zxroHpb
TaaQSNZ2vS2fJP3rEjH8hanzQIRskzqHKh251hmBWaBcfbiPuxUEb2j9SRjtBYkT
5S+9g9Fqjb1ODxeRWsbuhMovuX3QO5fISecJh91Z1qXz2NnofEr7tv+L50zON4TL
j7WQY9QwgMG5Uq0Tzn6ENmM19rlAEQZcxGZ+zIEnC6kQyLh8GYuMi5pnuf1T28R6
GgIR9gGDFga2n3Nb6PiFxQSKjHDU/UXddhRYS+KnDFhK+JRIwtK2N7RDzt480nNr
QRGwx4J9XkGn9MfojxIxhdNsW65M4PajzRG/pYtsJjJLViH7Tk7OudyNSw6yK6jy
IyfspJr75+B7ZjYU8wMxYRLMBJGnBgRmDxihMNhz5/VndKCkptjJ5g1XNTH1Man0
2n/7pcCBE29vkra//jiq/k04fd+9moET6bwcSxcvZVOOh2TWf5x5m6AbcpIfib+Y
IzZ2OXGg/XtLsu9fu6+qvJ7zLQh0WykGbOb/OHjrjBlVmNaiNIw7Y1xq8Ezb1afv
SzutA4v4HnJjCL0zwmAajJ8/xIe3s+NtgfPEuyY6Vs7ydNEgghehz/c1vlnwUGNK
BYa8jsdktJ0QVY+nn0IS+ShXlbnZD3aaXCufDK6z6Xf6YciyTKznWLawKsuS8qdw
NM+kRXp2Vqj7TdVNrf9E7oD4YNvgKBCs7hyOnwHLY9w/78ZYJphDrgjCoZBrr8MY
hyHaZUo9hXEmbFvPYoHMHuTH/rg0f1oYRH0KLgYihvbZQ614IHN/Pk5n4CCotrUd
hzbOmPvbzgtqwV+5bgY+lx7rf03xhHDPuZKt6TfqSG7/wiLWNAkz0hw0AexR8LFi
hbgHDeC51MeEy1B2UGChOmS59MdmRtatmK1fUNx1pzoG1vPgPTLygSlLv3tu97Hj
R0eUVrLsoJaENQ+0xBRvFE0uevry77FZu6FlJs6hhNvmzrn0O+H3pW4hv6MXzyKb
h275nSJXGC7IEGqnRKH84a0Qoz0rrl+iD6g1HN/x0F5iUxrVeEOBSe8zAuEMHpK0
6YX/M6FnYyKsl2Z2erpf7X07NlCelBUDjUy+hPj4IpdBY4Tjj+Gmt2K0utS+xcdB
oeaSARDgEIGDlYt5//PIFmzv9ymqhs8X/Hj1zQ1YLWmOfrslCyJI3dTD9EiNfpbs
vL6ULoUDm6NLXM8ASuPesQ5adnEYIu7CMcI+Frolnn6JU8A6bWpX5PY0Ge2TfIlF
q8xAfvKrdZAKNDD/Bu6wu4dT7LNttvZzlKu+3jK4XxI8CVKIiAjg0lByv6T3InbS
I493qZzv4JhFY/eoreg4oHb1Ryfp9ZpOS+fgA17JvSKWGwnonopwon/2HlSDMIaM
YZQZJYLHVJmki9fImgdgEivZPQPM+E9tBujjAUmZUIjAMM1r3QNOZ31EIs6VMJan
CZrQ0nC9XmRdB6hFt8fL/nF9L3vSW5dXVoMRh5yrPqHAOf2iuH9TafYIcl2sUbzT
aNSJfu/3N/BmliVmcSmjTE+8yF9ux65CdsA8WjNmsEjaomx6pAD1oemR7ghzIrdt
JZ7jXbqTVin27nG/Yjy7Zcfz/80kFEfcbx0n9Vj1vCjNtcnXJ9fyFrbEAGSnH6sr
5bN+35jOVg08laOE6BzL03IWBD/nWac5JObx35K9zZ3wNofj49BpWru/IW0zvZX4
539prPVwF2Tjrgx6y47L465VocXrVoYPZ2hPGjLXiHA2hQlH5uHaV7++FscDuGeO
DuhIqV8qMsma1EgULQZ95O9z65gu55XPj4RO7FrLtY40K3nK7rE1sJajVTkYiCtM
rf81GHjk/QpFi+SRke/xJQWpqKdHb/kjHqNUOG77ccB+kwgUAz1LkaX0lSsGkO8f
RKBAWdn+HQuXeiKxrvfaiiHj/kGM++1u/0SfQlE3xeZHwlMB1tTAioR7sCOSjX1s
SOV3/phA5V8HHtKvMnX/iS/HXccwKyd6tvYoDsw0G8kpIOU9Mi+Ro2mGUpCYy5lD
Qh9jyVmhauzFo/c2VPGDKOHto5T/DfHjPBRZb0xmpYUZLbIHXHhxpOaxp7iE14sP
AyAqSnxa+2sYXvBaA41SqxUOEFBF1uDBBUnh6nXWVRV7wnUPi7/OHfU7Elpo0mSd
kyMmGF7HedKf9r+7caQEnDKT801jZctyp1LzVnXD1i8XkMDbJYWRAxa9FIy8UnSA
4kaeLhyPidsrdD8xJfkPclAdvgFSTo3sXkc+azHwhQi4uftvJX01BRW5dM7Ge3+K
21NS4SVzwOq/ToNA8VYs0VTiGxSuFUCLJd/VL72fbC0A2Lya4wKol3E/+ImzkrnJ
6gKqixAHfsqr36cz2RDr4FLVaZX/3rzXp2qWnqeWEUjBKoHwlBj5WWFKNVx+QPkZ
3wwDaBwf6L9g9gjF1tNfcJZF4hkJKFstUYvu7HqDkjA6dqwOsb2WsOtW+KPoBv22
p1DrlE3O2BfryFkvsgo1nYUDsCF0EKk9b0DgW+EH6aJEcq7uQBmR/yNWmvps8ydW
Zkxo2a+yxdJASYzFcYO2/cvESmkjlxCQO0+2RoLMXJdnYqSJO/t3pncpIypkpFnL
VMOWiYijFkMZQGHEZvXPKyoDJRfFGGX4j56Np+z9Q63lO1W0vfB/WEUPTC/DnDge
ec71hSP4DeQLOYuwvwE1cAkZdFbBCepY+ROToE86sGhH5XJMUSvlqTclbNglal4i
V2R6NNgxFOV5i054l3AS8ePmp2nYWJpMvyBszVT8Se+KiDcdZwUqQDcRmXfk+3A7
+eEnRzm2sRf7rb5OaYOlXWBuKxm38179azIhEdo4R7Ng4KkGaZGSPmJyauO22U0o
z9W4hb8JWKnTSMtKLpNBtkJjYlEWc15hgFcqwLTzeRNpnN+Ym4QWfsJuII8Zw94h
cBE2SlnL8CaFe4VqV6yhaSR+CA0ClDs38Yu7WQe9kJBIYrBuu/PBqVlt623nMZHk
kbJ6MyGJK2JI8PWLa/rOp6y060pUgh4oEaKAsWwMDdwg2P6WA2fPT1EtlgAZ8Aj+
by+U2K5tG2z0ITT3L2Qp19GHtJJ96b2UjtYCIUbaCFJKmaxoMMsQO3SejMqtG10B
HLyF/NkorVOMP9Vutu2VqhSiA7qD+9rc9QdOdouXNYYGHKzmoZhNaAy+zxlj500v
MQ1cZ2aSkuC9zhi+Mr2Oz1lCota1gF4YUI49ra4iF/b77khkXXwrhv2qF5/s96Ok
V/dNwbCbxhc9djXTECKfKVOqYJ+hmyt8h+cyJ5n4Mn+niFIpNXGgez24rKaK61JA
NtfNA74asByyMXXbGSg7axArhfDgi48mUNHdjUkVDLu5/i0Et+kKjrCGh6tLhP37
ybXjO4YwuwUJc/DdqnuQPt6GZQjdp+T8yr4TB/ZeE9D/N/W9lVvvVX88lWsjNn0/
UDflCiJtU8oXmHs6JgLJnpopkG8wK2rorsjDiKCEzRPYPqDhJLo2qu/rWl7MSFWD
dKFy9izcmZ97Yemg7jWnJD4qiGsxzMhsnEMcjCaVix/8TaVA89qziwutS7WGY08G
3EkBTDJpMvX3Xoac2G0Qy/VpXHwNggWUY2Gkuf4DkHQY1p7FRmBOlDD0HaVAaECN
uPNznJzJB4qF/jsQShAfaVQVNjo/rC52ji+eSnXrvOLU0yMapMpPhDfCwoMD9pYY
brTMdJ4M+pv64B9GHVarzcHBWNVTxQY+gru18uCgkOSNHx8+Ml8nFa5ELp2G31rX
s0r2R6qeSSOZ7v4N9Qyv9pw3IQvSTN1MHrgrjkjo8lGXwo0GTZWcZ9BNC2HPdDbT
N/caIdEc9ugoAeFnrOWfnviPFlDPBnhc6en8qT2bdJSyyki7pLS8S+B+K7iY7vCm
R+w/+ZJBNHtAoGY0hNPL2S3BEyAd/YC84i06/7C1TuVhSCqkAazw49DsRZwILjvu
dGhrPWe57qm/XuoQpHqnRC2z76aRiwrNfwK5zDKkEDRTasRF8TrA5RWCptKK76Ps
Jf4milN8skw672ly0YgIRcqSlvVka2mLTBiqjB1O1KqYxC12CLpk9UElB4NA9xGe
eV1ZDrvKB/6vcXJ/Vlpah6rkHzMmYNHqvGT+p+sQw9pGcbsf5FO2AFPOqm9fpxop
+4i9rDH8v+nhKmMmMrC3lormmmnHGPwPfofyPODCrPtsVLFsWM62MwtLz1SgNTnj
xCgZ1Aky/0kIioTFutWi0dExnBLC+7opoAmAbChbGAgdKYdZdF2yQtUfiAeaNscD
cavvb8+0SL2x+cPtN6W53RfSqScNAAo6BPgQuxB2Yk/V+T39QvfLOFFf8lRILWXu
uIWkwvUt9LSoP0NmhkJkfz1rUpb26j5hI67CY6TZgkC7Xg+oMz454NirdTIV93sA
+Ou/pIFchdWIqQCBNIy6tj6YEv+uaugpc44nhVptFwU6aW+rLKVo7PYhtQhsEtXY
8gpR5P5pLTZLUTSFUUoO8zZKBH7D/NxHR3Z7k+7ag+IEzWaObM6AvqICCjZN1G0c
jtE1yDFF1y0KScyagGeNV9e/I0QCe+zf3F+KFWU69BHJaT96Z02JMS/merN+KDDv
cjVxp20V2TAolvi1+rQTcTILr936qNp+SiOvIXpdThUYsaL7XoP4s2pYIGVqvcWW
RwlGuFctiJl3IkHPuqm/WLhpoqHl3UcGxqPhvv+4iDqb1J5vehdx/CjYFkcZIyH2
FnyqeN+WsY3XXtOiQ8flX07Q+KnEYNtqg2uO6YQ3YrTLw1zOhQ0AXddDyiH+BwV/
aKjIafvBTVE9z1sdgbjpioHrK2ZeB4W+TL0pL/nI8FiD+G1j25YcRAUDgMjKaTNG
VnevP0Gmy+2C2qI0PNMC0POZgEZ6wiePy9A+COLN++fSoqfj1I6t5djrBv+2LIAD
n7u0Di/WbB6GCYFFB9/Ha8ATVmBJeqH3Bn/Vkd0o7+3TD7vukZ2axdYmVWgBC81L
xhc4pVS0WaIcotPz+nF68l/7D6A9Q6abJLvYBxd46edNpQK1DQ+Q5xA0b8TYdT+0
K3DQanyJ8XzUGX42D757/XP5M+ckSlYtH4/wxOjLkZ5NMwixMGoWDNTv/RtMPpQc
qdE+QwoQ0tHYGKY7vSAcPL/JDskCwTAQdc9IOGsTwIq15LSg+90Bn/0hxfGDQwS4
oukwWxnO6X2unl565No+TkggDDBG+X97oM2uEP8bGSzDlLEWfcKa7+ilXhhqdDuX
wVrJOl2d2pQ5qZH1lNjFo1IG8UElbCtb/5wRRHGIxrI4qO4TQZ7o71pNVfYbH5eT
ngTO5aPDYpF/Stm30u5NMESuSgk0z7v7F8kMGoFYMRa7/P3By2WR3qTgZzkcg5a4
7KGX6F5JiAE4iGWv1qoslWkg1E5uLqU1wwbbSr9liq+d1xD2HGT0GPjlGY2g2fWL
I0Df/vVVXDEEFdZuZADpJSlsAAoZagBoTvC0YTkJo8dj5TNf+sQ/jzZBp0Iku+tB
7MMhUoJBRtHmMYxYHlDlTshiSpsR8lcQQKRIBzmLTue7tN2Edcqh4X10nqSIQKMX
liPp5wxwsRKuiR8I1pr3LBXKPLpRgaLsaIVhLbsZ0fEWOAK2anMA5olZiVNrV0xU
5z3qxD3IXoLnuuJsS6RM9TnFly8C02Qhd1hUTRRypLB23jkMed/5xdVGMDNq2rx7
ZbfxzyRpDiKlvePWgHraheKyAYhLuhxM8iY07T7MfA1vlx0yMjY3tqnExZ6CppBY
ErwpQIpk43azM2p/yXvCVWqeKMWFjRG+gGpqnl8Ssg0JudGyWh6tBSPDLgtQrI8z
YkBCRM5C1BYRQ+kgeiQdCOfYakU1azZsbOaP//wZqmjT8eSj+v0Mb9G57PX5DbQk
7PIDALlqQmNNmTQmIMtHPbPJMVTEa6u/XekS51j4jkpiLUiTdVN8Wz9vE5+wOf/L
djDoeod0fJagB7jf/JZFF06UnNFlpxOJ5/7/2K79Xse2rAvORpV0DPcZYsZKIRM+
4/dUzI/mOdUyybKnYDP15RJo9clbV1Cl22HdQQlXM84DnxYOrgx7C76ypTr63WAf
t1a3WyQyhrXtTl3FD3GO7OVi+hx5xPqtIdoxpkIQYb28JnIqjMjMKnSD0okDPgyc
PAWSyKsRpANAR+/LXq5N/JIahnA9oIqleZjsVMh4VqX98nyvuD7TDrbt+WP2gm05
EX63E7hmNUhIQgaASqzOuPj3sVDEfUJGfmyqNTOHELUke75208QlTG62zK5hxpYn
qBwwl6TBbcMtiaE+HUR4tnHHOmdLMEQAEMAUH2u4p022aOlmHa5lm0p4CDXCgNJj
Wtu6IOy/zDFTVLEInD6Mrgy2/yfEL1D2ifTtPKlnSSB1SyKQd245kmJ/plgfvi3d
7Q6sO0r+cmZg/CkncZjGX/IOI+7ZSrVukqjFHmWJSUsaoipFbWSmIOzAPxbIBEhZ
XDRkfASmlISz/FbQ+PsNVQTV6tdWa0gWDfomAYHwAaOq/2VcLcOUDIneTkopvJ0/
N7h2S8Hp1KNUdWTfzEnvr+g61huO8GIb/xIn9tHw5Qrm1N5C1qRLwPZVop0jJ6rY
QlyLkMeml1lePc/qqe2CwSrXcDaSUvtAphzQSSAEfOKKugMfkMJcDuWPhwUK46R3
pwSnlbFV7UzAI528fhTtnVP1oBVkpETVvSKEifCFMAUbiYd6grOJruX1j7w4pHrn
Iq27uuTjWa3VvIGJbMWwCRZQ+6LO9X9+trea6R7wn2mCUO6GFW4hegde8tpBUE80
GnD4VptSGrDgC68BEg3sV0Wuix02aMkfyAAvol5qwmeBMbG9nuQUlfxPdM8nyZTx
HztN+ijoA0aadXKqT3GMl+Rba3LXY+syaQ1Xzd9AjiQAqk87nIUEqssvldtGiGY/
p3+IKJXzuqQJViLFcMlKYwRBxvree+ITeRB63g6rGzW31rhMMUB85zoA4Ibj5gES
znr3q0TU0tJt17yH+97sIO8opgHZvi42OyNyYhB1ngLZ/foCkV9+seWkZlvA9PN3
gYIZz/yKMATw0rbC2bzCx+emEW4DrWYUAez5lVq970Wd+KtSkV8fm/JfA1WjkzhL
ZLRUcIG8wi/U+7gVqc2YKe8MjJgx1/QBHqvaRtQQnlPYOTF1rIyxTyiTmXS6Zlb9
gUn5SNn5gER8Y1b1qXNcq+3mqbE8IF840CfcC0rIkot26eTPWJhDNlqXr42HpxUw
ibR1i2who1si94L3/5QZnh51VAbovlIV2ttamOJzlxCPaIXwSHLHB3rdhjHdYfIZ
I1+91LU2FvwgePRZhiUcIASdHrC5F+McVp0zSmxEXQ5ZL5l72/1GPYgJlEccKmwj
sbWbacwBmh+7XgA4loZNsiAZlFIeKJlwki27Vr0HXF3LJ971TledS3PqF+SNnQwv
djOBP3mGJOPTM+TO1QDpZTTkx4iA7yp+gJ65Wd/eXgqvVHtY2noOElM9jtxlGcFd
KL/ozeSpcndJA5KNcO7GtQkzvNedHxMGZuFDqN0JB4OEgGmAPeS0zwzQF/FZFygP
Vk83J/y808XL+kosBJ7SrmJw5Pw8s/jhEPaFY0E35S/tqbuOd8oDxFuMCz91YC86
RT5CNSJ/yU465XM0WPi+RTdfWr+FzczsHBaNuAorLW1kh62VtYruA+jLbkc2B8yI
VOV3BwAKyC66DeCPH9a7kXW8ygVlIMPC2rfWLzSxhafAOTVOFqg3IM9aASbNbely
HPqH5YNMGWQQm6GcCTMUI4qtFMr1FMwQEljPlMtdDXTFbk4Amlf4aA6RHvFlarJP
cxdz0RGTu4n/Rt/MZsSYfK4MEPllqMERRIMJuR9FfmVunj52WWqS9uTA8RY6Q0we
1XbBD408fic5eyFPsdaFHFt85aMnJno1EIhvDisNq842Hy/nFSm5Ypb/Qjb0CNB2
YoScJvKOZPwb8yDiqqkGCKlQoHeL2/yL4pZOzpabTZtjwVMIMrN3uMzJMmquzN4R
AGFJwtOi4OAjToDEDuKePY97s++tcdwLyNyGq1xO//Jm9pYhU0ATeKyKaZ9jEwYw
yGr8rkFXqeJcEwp8t+GzeEOC5HrFES+N7SH2vHuJ7VwC11T/ryTPw1vPAAuIc76V
Q58IqAe/25Unjn6DuYKJoK3OV4arljEAKZNWtHuCOU0yelf2xmC92ZULzr/NRPNv
f8/MykZsctttyZPwoA2Neulzz4A/Gjo+T7+s5FqaBUNV2ZdCpP2tBbI44XqINudE
5XlUdPpHHzq4pSamU/nT8Y0U7wIdI/I310AN/Qd5RRuySw5et08BQYA0ZJfr6hAS
MxN1WYLQMGpLbwRK5oCb2t26Ph2016/2NLnutddsElt1zk9kz4d+KsMtzkgm3fMk
WZ0yW62dAE+KrsJpK5JxKnpV5WTLKMJVu2pmciihxqfQ81zLYGx1mAb1Rzr7MDsE
UatISjEXaZ81dpg0hAq9wGMs9L0y94FlUddu0vdeqxXGlfU4G/clmT6IPX+bmkGv
wq/9UZYCsf3pAXbGAyV9rZhljJ7Mhq3Ok0QuvArn5b0Xoi5NYAjeA30kpIf2cK7m
gTGuR80jba4nYB8B8U0+2rKb3CO/evL0NNZvsB71CKT3HTVeaZZdhSbLa3WzmYTu
t2683SwDVk51GcqzKcqg8KkK8p5/WEp/yHu73PEv98RVURD8RX2fNx9oYedX5rsB
JOdPxt8Q78cNzj8NzNlVssP2grnc7Dsyd3Pky1ekBYAIZFtt34y1ok+JXnN1Kfnu
suEOdEQFMFECAmeZ54y9ZKW9+jdzdu0e+SUxbe3UZSYHO4MHhJvz8Pc/uJuwKm+F
vXz7tEawF2meMvYL4hzB/02qxrNz5Juoja9VQ6FTvgLCrM92YI5BzN5OThLl458f
0PkZO5nrIvOBqbzE4DfNuuyoV7gk65EFEP45680RlxGI96vAlWL7xvO5dzrxhDi+
KIv4Kz1Jd7M7q4w+/4h2UvHa89hiOc9p6x07gY6pEb96/p7SHuW8gcVdQUIycphY
/RxwyNMf+dgMT23cZkry+x0tBZF2tykGlpyS91R3YHF5MWpMpEWgQH0pJvdVgiv/
tqcGWSRYQfhs7CYXUIFN2EaHMzHygbuUKGi/lZXjOmwG7EtZitGXyAprPEtEdzQE
0jVKN6Osn4rLdC1Z33EvYcsf7yzJFBbiyPvMnwk7yhGMixBL6n4V31SyZxopTaLs
J+vlMrNf4in+QowKJrjknxpY4xiC5hMGXPANXsoycTxkDklVE9MEQc7zT8ZmpEAL
JU66RfiLFQQgEiOtP8eq0WzsS0TORNRpu5mC3H7DrFGClciztMSgW72CU2XIwTwG
rKwEE89eYFKd/MGypw+ddz12fdeD2ot/jD9KHpvFb6oxNLp8yqkiic5ZOwLr3Htg
BKNj8Yzke4nuOj9np3SHLeOSh9WVWvToYA53yuWFftTIc3Riy5QpCoTvJMS8ps3V
J/3RBTkiab6xy7qxve/qJ08SSRloUJoFce7OejIzOIp4UcfNCDujusH5VvtKFNWA
n+8yP9lxufggN8x0oHAa5T0GTRfRCKS33wDa3sH0U5bLBTMvvhVG11CvdfnemrtC
TVAYBOWro3MYvNscfbRnE/9i0daxBL7duA7JKsHEmwej4fOHbP6UPRb7a5z03TLd
OpMfP7d15nZ7Y7+xg9L0o8aTve4cOdZj9+UzrJIl4SYVAMbXXmyyHSE8o7VIAEKj
YjICARvDRqezeY8UjoSKlGVhVnt4IySZJJBicRhV+K5vt85FZy3pQ5SLyyYOFzof
l1DNR41ztj3yllqcJTRvpVWkPSCZI2AKkWX/lggeUHbDI1K44Lb1Sz30tOdEp3dP
nRCngIDvvHzSTk+sBWIgE8I/HXapd+1ExYq5m8uJtmvGEHtS7Uc79rJ/N0JmyEjO
T8geaR8+2KsEehjqZ9ryO1YoCylmRRcx2nABD5xDeK7tucGoee1NTM9vDfkus1iS
O/SQKGXBtb4UVKxNqGDdhII79DDoEoQzh7ZvmvHwUyrkxadhmL0oPq/93f+gcQ9B
rGUHgW7bU+YQRRcz1P/pDhS21fVcKiPFlUUHAfVZoFSodWApxuht+vgOvQV0FB11
H03MJnaVwtVT/Kg1Zqp0xTvQLSU+lr0189tkaK4sApwwh++NfVXE0HItsxzqgIfi
7IgaMal6Wsy182rc0E2uxUeiiASP7qt9lKikPpfOjLkyMv9MkGMWhukoa5YxQ6QM
K2YF9JJIBHJ8YZ8hGg9tv3mgNc6eRr0neI4ROKEG8eBCfm81qZQKqLoihQem/Fph
qTquovy50kQBOEa5xFnTQDULLtngXAde35TmN+lxo8lCzoFfYE7vqWVUty5vUq16
7TechCwS2wLAa6514V597vSW4AdEW1UJgyVDjCeGwJvdyKwYXet9gy/4RofA1iYE
X3sV2bB4hBQ5zEPqWJKXcG4fvbW4CIksUNMUMy6mhGKJpPWzrasqftKAP7gS6ja7
nQ1obNnoRTAQUwf+Pk/DYpxMc7XEYw4nV7jMddMYB660XDGjV3rNEvTF5ew6wpgo
e31Ucty/RdZrfapL1Ct7cTKVPg2ZesdqpxAXjw5KRKHcE3wTrp9OX83xqsV2/Pta
ygASGTjPZp5lYqD21dV8HXD+l93Nf+lavGmHqYh+gaym9W3Avg5RTnGmGuxqoGKG
kXxVBjr2C9YP04v+XU49SkOeKRqtO0eZy3IpkgZQ/jG2b85W1kHiFJzXxuTMABrB
I5F/zVjVGvR+bDUMeexReApJXib+GTuAvkVErpgj5b+JSeCpPCxsgQ4dOhEZc26p
LMWowbAFhfkWZBZxFcEZAjVTLcFf4N7F5GG+BkUICG0Cl/HarNVhN4PxWBIIqs1o
/cJSHwtA00EkX4EEx6AXUcaqoOcBoOhqRbdj/DYjL9RSDAVcl5S8Bw34cJlFGL7v
GjDOUss5ioSfZsLSmfs5XpUEwAClovOK8PVB4cQGxkjNAJXzrCug+ddTAbHQXkie
BcIEBmarTtZAeByFREfPF5z2k2D4j1bNPxHavjFnAcRWyxMlWxlgoMiyV3LfQQY8
YvcxSZCxJJ8Im4oVjbvk4KfrXsNUSFGE+2hys9fIpizcXvI5/Fs1WPB7jkYTE1vP
XPfJP5AeZ5F/FK4xIUHL3HvZYgUBJnB2HYKAIT3eAQjahDLWZgfn9NImq+4UE1ji
QxDi87S8AE8XjOqP7nnutuVewgiTI3NQ6cZirrY3QQoP4XWPREdzgH9Aet99xxzY
B6EsJaccgCimpV/mOj5noHEEinz+pcgEKJp7F1Ef7cBCwsTz76KQEyhUieLx9Kwy
JxTzpertQmvG4Bze1CdL52SvcuCsBvtzA2s9+2AUflxsDm0picJQ+v9U9n3ziSDv
EerGeTw0grJ/CkpRO+u232MlbVNcWOWq/f0E8KjXeq+eVY29+wwL6HaCT1u/MYCA
pjI4Ikpae5eXq7QzUGrBfU16ZOM+8cz/Wbru/cZICJO7vOaejhcxx5BPVak0SbIt
RgVr8/QDECSyYv7dUIQTiaZ2t76rUgdwF5EG4Z2HOXMkQ4tWeKRXkwXFXG8t3Dup
lumM04d+NMd67v7qmMrAA2QcdahwQVOq7Yuc4nPC3WvsS9ChOEKS1tKU+v4dq0T/
Oxxwe675GRnPB6hLBe9Pml5lOS9BHotE8S3MhxyNotRhKzueiWuSoWlhCBcqFqP/
BlpHdmdA8/Ms+7p71/2ru2zDxswcP9xP7Wm4WFKQjCJEXld45+bFG2Mr7QPqo6tM
enRTrAr4iEloaMTVJL3cx9L6V7HBsptYne/ROFFUN9DBGMDeEaqq/ZBNSkdrhiSo
Ae+DyiH9c2ar5mqddwXjF51HiVPnSuZshi7a6bXPFZ7+nsh86BuLJeq2+xRHT+ml
aOO/QWfclRlcJy5/Q7AEz9X6GFc9ZWKHBsVtaNZ9PZlLB1mvhGbsZNJ9ZWQyUMNt
DQqrUY0mFtyWguEWDmZi/hgpdbpnVOKutaNJrd7w9BqEDAAFUKKVaunbUbk6A+7S
dEiNP8ldi2GiZjOyb8qXf3nCpvQQi1RQrCZqPVB1vgoMIQldMn1w7BaD+69fxIza
xYfzc4JYU43yffpHXYyDTspm/w9Afm5ZqSv9vuC/y3Iemj8LiEipH6vfMpm/PrqC
JLPODQR9miR3dLJva7YtUm+JaAENoa8UAKkKf6bQJhnCzkCLULTme1RyhRPDA5+X
lQ/7qeNlZsEubiFt/ntuLDSOBka/i81r9tPVRgicPZvuUppo6+6i5lSdYQr9L2hf
LzqdzwMCV6L6yGVXopTgAX6/LWO6dyBoifUKt3mM8pJzvw7lloW+EfswrpZcqNf5
BPyyGAqjCLWr2hpWAq6MNH0viboGvWKbWG8yEztvExs9+h/3PQim/12VmpCTRgYh
5CW6QNYoKVSaIjvVDWAQpG091NsIUH2oiZTDaT6NvMQdgn65e93IzZD9QkiMDRQr
Bjzxf25PI9Oo0hfmghrD1Pt7qZKK1P4NepIXNtNUnwESF+1z8Ow7oQlWmC8GqRkN
WmsFrlyln6pQJ9/Pof24b/yu0O1W///nKoUThr+JUTRJssoVlskPMinDFodeFmUn
TKMzoRB90ECfV62TEfHu5RMFoduuIN+qWsVuYbq+E51TcWJQMF7Qt+A0u4UBOWgj
yU2s5JaqPHhZKnH6LFPwzw3fOPKOx1NX4V9XEh1kpJmkleE2/9Q33rcJ05gw5YQu
u8FvA7k6dMKwXeLmg9eGu0eNR6MMFNt1pfVAzwZwH3I58nlEKbVgtJG7h6B8imF0
W4z64zDBxAA7N4k5K9OkabdhCNzj07s9ZWNtFQhmkcRyu0TQ80iJJi9erD37KwqE
B98o95dpHLXoQkmeulqv3d+TfdL6VvKMYO3424ofBkWm98U2RvAbj3BvuXQ0BaSb
0qyuV6rX8bwOW53cm9RmdX7Wxv9+4ANMPIzJ6KNu06EyDLKCwWe3riRr292RE2qr
BehVhfPDrQi0iGtj7XHkQh3cVk2Pjc9jsNGwxlPyg44HE75ucWndf/1+TPsGq76a
fUxvuqlyMmTgR5sB3f8bHXCjqS+PJhC/uAffftvCEMJ7qXgX51G3j9zrsaPnp24F
8Z3aAOddYjGtySSbv5cWElpXIQxN69nhDQOvjvZDlyNKYO34lNnSws4DJhtciHT4
yi0GsRYVTh4ml+F8fdEsJ+GNkkVE3czn97THPz40t4aom8DJ8GZ70IePfA90xtXc
y2awFAg2LVqoBhbhCKGJUyE6kdqOruoFRwtxMkYNRNH3T9/4NFMyEezp3s1vSkO0
JvOWpWJO7GhE7wX5N356iZBzvLzoJDXkaRgvjIEbqKAM705GS7QAfOmyM2S7ndlZ
OTcKox/CYhsqbXXldB0F+vEbugCtUejaaiUosaQLrzL1uzCSN4UOPsU2y/lN9/ny
CxldZNfI4NJ3EY8bMtnEk771JNm8MY7z/dhOF/TaTqhj3EjtvSzvKoD+q+8MPeC/
5lB689+y4K/K3me/ktGLKufYtjm9ue9KlqHOEZin4fnD2vlr4umIz+q5xlA0oqhb
6yx/2SjVIz32du4Ye0ZxfNgiS/T56hZL3bRYiqL3yOdVZpN4D1NIAbHJs3Gj2341
YVTxUF8/gMaGAJx0PXTFyD49YnymTA1e/ScwynjK06b1fsTg/b8jSp12XfEnjB/p
cCPb0mQ5VGQMFHT5SKuK0eY4nx+zMtjjQPfNfOGHWW1Hmixng5ApVNuC9apS69JZ
Gm6pQ9eYaSsZ011bWLVZu6zDf+WkmopYqKLOn6ytjmAoN3rqlNCaeYA4+Rlrhaaa
sq/4kuzXu/ze0nUESkngtzHPCPCDOao38jQZ48Q6Vyh+6KQAjInDpeg+wND3BnN0
d5GogwTKJrj6+a5hhG2N459+7xyBDz1pU+LCtucbzRH+n/C/Hm2UM9g7THMlxpL5
/nJgDJevu+7zWewzeEjMJJcLXfvN3ARI59hMfU1SEZfHklf2WP8QhzXtyGMcDZNN
l2APQHqgq9QYxRGEzUOSFIVbLrm3Y+2oLOUz5MVYYtGstb+F24vwbPOsXreqinfy
OSfeRInA8K0gy3rap5ScEsfEGCyCJERRihVeOhD+vTmXP5rkcXZ/YOMVNURiU8Yr
ueK68Al9Yj0JD8a4r1mv8AhbBeWFJSy1RZsK+s4fhyuIBdUYlcbS6rMS4EG0KTDK
HUrrSgK3Zs65IXdxvBzNYC1pgmZfi/RM8aCSLP3OoSx+iFPLgp8hkvW5v6DXdcn7
7Wv1SodyWcVreR3ET83PMh+Mipc8M8vmUq3LL73LcJAUyHzVm4hf0Z3AJWyFEWex
WT1HmQDKpFbPKRa41OXshPVQxT4hDRxrhrsLTv9gmqvCTmANPJ7D9mtY8g58Vg6k
Usm5FwWY82+c/Yt8/kkt6117arZ72jw51tgeljy75UzGgc/XbdLWIuuyoJ7SUZN9
Si0pwf5Ex8VItNpfbXiS0/EhYfWMzFp2zwpWalBm6AAPo4mwnJvRV+KxSWQjj6HT
KVSuBjmunNPm03tIfUyDJuALL2mbyGPJhTQbAkCiU2Vs3owxwhqpB0oF2E7K7T3d
2P5gWC4Z07EIrwWy5gHVPSJfcAR76TuDF5blhMw3rD2P5lNOoRyDdD+YyqG66G9L
8xNDi9tcbIRqWaIUrQRM+vDnn3jop2oKTEF0RSuqbs7MksMclkfwCC2xrEDblog/
beqYrjFixOql2aj0auw1T7RubynRIeIpY1N28Nz0ZKcGjWdPaLN/WznTlc0TXkt0
nKpZiWeZ/f7JBKAHoaFqnm1bjVi/qHrRltDRQhHy+kSNgzd+UsszdiD07/vsR+Ct
PupSdgWOT1TH8g/RdBOhMAMZMyLDjEZEPAKQByekpmMzKVzhskztRHQ3nOM7OYrN
y/vjg8PzwR7xYRy7mCVRvnEuknidKNUMULUdiePwhHpMWonTrRfBV1PRVp9rThbI
hlAk75st3hDpSZ2w0hy4uCCI5iZSVUbQGFCgf9Cds1vtJ/cNApuM9kbSTI21Fx5u
YjV1i4nwsWlg3I++y0RhigkVLxZhJF7PaqfR0pZXEZYttZ3aAiy1fPvph8jehOzv
v5OLwl2jhTtFlfeLzaJxf7MxsJVZwVOi3KdF7ro1VpxDd0UgofmEkXWHO2WcqMWw
+29UGHgL1+uaZAwizzN7v9MA6nvs4/4pM+lKX5bnY7H5osrBHMC8ADWmNDV5TQqY
tj78fGrTeWJiz/zoiuNoqYw+FwdGOWV+IIdhNucneORkaDXVibY/ldR2rCJfGqcu
w/ZhnUYSNrCkFkCvLfKMcFowWkDaAPCcY5X52mA15e8RxcRhNJKFyb30g8TEdDzP
6tqCvtde3YrjfyyuZejjcS7Demhri4hQkSMQ4q/Lc2qlFZhS4lMPBTE7mvjvoTYl
MqJ6gVJjU0g2AS84Gj968+Syh8IbU5JP+JV48sqaHciJcIu+eq73gH6Mj/8rnq33
MIy1TLyHG9QApzPJq4z0zYMtBDvQrtVs/UXAk2BjzuQVwiooHJh+2WmRq8rGfJc+
jQYssOWsreiQg76TdN/2gUst/64l13gJOueMLxusbVAtr50Hx/33YpEhTL9eLbGZ
kDvjaJ3loKI8WZ/8ddNrIGKjpUJpwjWOMhNGIhkgZjvvGgnyu4Zn69GrWYLHT3Ot
O/EZwYvOmSVVQLmcorn1B4thoSW+CuGDYRZx7EQRqkgwRN/LYtEopz4uu31YJdrN
IdJct3L1jlm7YcB6bHIHvzUUYH2UX8vqJ1lV9ETSCZbW6iLXZNACghv15ycWxxt8
4D2ccWbzMYcJTrsW0N0Jhs3dBL6ITy7PM30mfW0ARt5YCFIg1KEVUOcNxIpnfHdC
Qqyse73qTSL/fK12owUjqxGi2kA/atzLrywoT2TJZ7EjElNb0j4/kNrK4nM49L5M
HE3DV42q9K7ITmpWclnLXBit0QHaVgeWV0hy1TYqyMaFJ3pxxubkXyou0WR1v20g
8+dBeNxOui3S/dEMBul0n6DtUQvpoY5/zU71QsEYAWH9S0v8wxYKFpbUyfaSUZdO
7R4B8xiCu+YUfzxxrZS218gbE8kv/4TtqTh2pnZDoqmSOpgv7XXdBERVZL+WJEfZ
K1tGiefP8P64q3TC2S0GAQtrmoS4JG7pedRBvM8QLiPhNnbGwk9cu/LomrErx4sa
TIhediZ4HMm+y7tsqsqT6NK+viFoj6ZHpug1EL9epBRjM11WOCDKojdFI6Ag9+Tk
5Fbjle7GvnP4ndG9JkJxKkPJiaTlauD0hkU6UwqGTMyLjC6nwA+JyEWXDcUMIbJy
xRcMLn39IujhTTg8oJ7wxLu9T2m6YzN6pdg6yii41dZQlGXEbvFmODUnTyyrclnt
ho36SeJPkYWUxZDJVjGZ5CHuuUbr28Jb74lGXS0ndzY7aMNCk25bcnm999BrmJ7J
A2wJqQNIht24SxzLLPXlNzn2r+5CxpK+LMPtngP/dIOmoTJVld8LFYmxJzq87LoV
Ye86JXr9n0Y/8zpwFPfATr11JodCXYIk8/XStIDZWfu61I88MJ2Odc1z9EPtVvGy
e19WsO4yXSVEonada6vtb7Y+ZnicQ0Nn/aOUP6DDrvGCigGMOnpbmefeylaEaOYl
SZ0ika8G6oVm6wmYKx/FW+35BQcLGyqJZhIQLrzVtogqGF8e28XNnQESsuYJERgL
swtSLpnGHkBL2i+rNC7nYiPELQqrrlPoPBSjHl53WOpjt/6tHkDG32y9gJMOmOG9
7x5Th0kcNIBJxRBmOFVWLqf1a1QYRSLRfvL3mbvMNRaNqSP3JKdTuPCJ918g2v4W
PqTqCPzW7FVxLUEIMooWY47LxImTa76Hf+DIcXpJ7KMMIAhsuaO1nZ6Xv8vjsIVg
3sawS6ISx9mCROyzqsGNf28YHUwpqbuhpdmhCmLgUopi3Uhqi7K8ZdoDzWh3bDhP
mjMkrfFf7myvzBHGxuGoaOUhX5kbXWvppi0wHe3m4BT9kv091B+/jBIcDuuK49rf
k8BiMsFs+TUZapVUnCAIrPyzqP6iDzT/KQgMLex4F5yWlg4keizYxLLfHR7p8Ou2
f+2TepVCeEUyQsHJD1udzdwGffxaqfPOvSCItFCyXoOGlc8GaWv3HCCUSWT+yUWQ
1DW2IBTYK8mv2x6k5HwEvFW02NRoDDIQTKXCeX9VVDwsbnsQ5SEZrkDO0BaDY/Z+
FDi0MZLgfYD7tFoyzIvvDRSFzHID/qmZoI1b1Srm2DbDwPqRCUgm1kcZThCh9R15
zzeHAemmLqxIQI+qqpQ2lMiajJKqJGL4kZwTjiHRAwJEfw/2Ow/lc+g78pHRlS0h
fjJXnp9005KPN5YYhXJh33K0NByujoTlL+6mnAcf2u1T1whbhSWaCdS1AEhfLlyg
KglqnC+z3nfMDOBvi3MjWYZtfMtov3lVYOa5Rbtg9B0V7fX5nqUFfYCFwwf8/w20
+EduFOF7aoNVgGN7dtYAEnFSnhrZ2Zq3gs6qojBmSQsJMYP5o+mN/a7M6yuteISt
sKcEiW5lxDbrX7FaGO602TFPVHp05QnHepdpVy8NGuVQHzlpW6vrprIHj0e7F/FV
QnoQ25HUyk9Teagu2F0A2Iadz2pwZl5ifr0sUMeKuvmj3Xqfml/eBDSP1Hj1IFuZ
yxweaEJHxMWCjxhETLu3i1tHvTkMocVH6jtoZVHcfEb435pXZ361M9FnVwvYJjJj
9pyfnRlWVi1Ts5smxqmRFb1SGblXl0pxZpBno1oV0KfqqPphhTg4ddcZ079LZPZ/
4etdH0G1283/jz4mwwei2imugnAMt98HDd1X6OhKE7DhjC9UMem3PEEyhuoIKnRz
4u3xMFMHQVLgnyQ1EffPhrZn/fFZPnoTW5uZtaMDpEk46hv4Eaznd01Az28croPb
L3V7vnPsB5sWzN4enA/1AwoHmyhCayBNXqgqzUgnU8YiRFiUuUcJ5mGTCKamBuSA
9aSNBfnS/Qc4OAlwoxtAP+nGncqh+AsjbsBCi3vGEEq7fe5kJKwHJ8kgoMAmwpxF
VbkQx1swBpieB1K6Ay9/ggXg3CPd1gwzk+KPpaANSJ8j14p+xb1FVfw1oUsWGsj9
PSsbG2Cg0ozc/IEp9UWrPSb+UCkcHqH9vDMwL1PTtXjkEJRuwjaIvKaMpTH9aFMw
KARg52dNK83cCUJ43slyTAnTvRC2PS0+i2YRylscLgn4/43Wb1MlJObkqpiIfTiO
gqbbDEHBwe8NgRXAkpDuEalFR0WKGHRq4edcH3Ytaur8t/jeBEVBu3Gz903x5z12
iWwkeXSOSASV882dgBLZrUA4ecMDARmCn4Urs81pDGC/ayaeHbAAMOhJbjbnBJ92
yQSy6ZRQv/v/j2jWKs0aSP9FXVTSspHsj4crtJO6PyCf1klGRl56LN/0YCbUoWGu
17zEsGLeiMst1caCda4K3Y1FQTcO5QYRWCb1PgYANxas4UJpVKpvFnA8+EKnkoHQ
3F0u1zWfa2zEA40ZLu/locZtMzqClS6jw5V9aSUC8YOYYOX052Mz3/fOWKFiMOGb
aUDLnDu/r/92HlHbyw2AypzYTrnExAN/5Qj0cBSHjujWbey+zYoI/PbNHH/1zAW8
p957iij9MddZOlXUM3ruwoQAeyvCYzYJLJHyIko+y96aWpypp1X72R42IO5EHtQZ
MFhs2/TLaojqQPUBaWXBfTfr9o7c6xlWJXPlJ6G/HZuGtidOurx640w2/pEDvfby
tybQF3LoHE+fStiyQqvawo7bishU0IyvcQctHwYc7++pn6kXastcv0S2XBNEAtza
JCDIfsO2YgonfQqyVHdhzoxCQRopL6Gbhwy6C7FviUxyrWWmD3pe+JfDuOUbfUfs
BeJy3mctw2JQ6DOcNOlmNEGqS6BH2wKpTgPvpk6W9lIK1X6y8BvSVFHn6iNub/Oo
0vYPBdOvO2B7lFyS1eDgeZSPQFFuN0U6obhUpuIjkTRxWUDvu2iP+Bd51oOJ/mXL
worADKUmy0Vraq6p0hZqbZOz4MmK9jfyKWEuhg09J9fWzhh/6WxZKI4OhpP9ruOx
R2+tZWoyjSbgYbDZLxUORyByGxz+GiEMMc+NBxFH4y6wa8ORRVf76moGd6LJ8Htd
tLEoHlAGhKDA8laa33Dsw3ZcK029/JObX8cixzbWtB3ut2tq/ZjhkwQ6aTxUGyEt
NPbBqnmR7Cw5YqxwyI6FRN3CUkSK6M3hUQ2XJKcUtxvWIHGtlSsn7/h7B3VfwesK
H7xmoXeuNSvBJ3pkSaHe5OeAKOk9XqdBtUxuKe9mouLdUZxKkah7IXJyw0HMco3x
FcmmG7mxnhAxnIvPhR6yO/S9wh3zFAl/QgNB/h0QPw7heLzKWgGYmzTX8v6w8O3P
1X0NQZ+JxZSAEgtI4zg2C3i1n0yJOYqxEv4h40139dbC3VuVVHjYW2L1ZM8C0/q7
6w/f/LDmfAsTzPRoHYwvNnc2ysgaC0HqgirYM5rK+khWyrEpsm1opaIGBgCs37MA
/sK/cs51Cs1Mr5oQbeyVt5s9QeBKnBWWrH3MOfq0LgjPAZMsmJ7ObczD8VVNP4T3
Yl/iSWXS8BYwP9B5K4SFdh454kvQ9YLo2KYL90DNabqflMmLW862xJdAIyngmeCy
ZkRTCbBw7vntQTjgML+VXWUgFmbmdAtlEviBtl5+6TSBtSukykwJsgeEW8JjUiRn
Lp4zEMcKr3PAAv6v8roC+hDX3dcXS92fKOFkgrYWsF6CB1Lmb7Ja3ogG0PyFzKWB
tJr9VBRvEHQpWV3Ltd5V0zya+NRysJp/jbPIO04wBwpQww8cu4Uvfmf0fYRxRNQI
HvxKb0+mkw+aCILrHjaoMCgJcOtOd9Ke3C0qSAwfdGGMI9IoGT9vlyh111p4Ta4F
4MwuNQkSXr6M3dtMRIGhAj8r9qItdJD21CfO+T7MEsvSsyWjIz4hSPoy9d9hf2US
zoR4FZDbKssfAbNb4PJuyJS3J7EAZYiC3QZk4ESn5utp5sK8trCxvXZrMNfJ/bqk
YJCDTIDixtGCS148Te8Cq3RySqLQcFosEbHZuJdxi3VYhr2Pv8gMTW1lKJnETQB8
WVR7a6s3+Kvx1ioT0HJ444j4rkBBbv9JyLg2h+C0nx5VW8RFd3aPQ1ewkm9K3Jnx
sNX8NYDDGk65tLf5X5aZPmHY9JIX1+NVpx9oztfWmp5ZIpXhUfXLAuVc1AIeaP7E
yabiKdQrY9sPQJOf8Q3IBNTgXTbLPG8DbrQRS8ccF31HUb1v8LgvFERuiapyRYI/
OVqm8IXHC2PvuKsEWvVsjYuvsfUtRWLdZcvc8a9B8uwoAxFKfvhXcr8Rt5rRTod2
SBxRLpUxEu87uRFZDLrlIbL5EZWP5+pZsqbciUt+vVxxPXE+jpRABqiO3z2sU7kx
xGKD/u2mRmvV9PT9wMa4A07QGEpItgzT7BtwOryl+WUtVqVo4m1owfAGV1vwty7B
VZ5QJLjMw9JakL5KBBypb60jS7F4AdM+41ckx0C9tuM7u2SyJtQDJYmecGiIlgwF
/h0goj9KXn+crMNOeY+XpMseTBSdl6NxXFgGyWw/z3zBbd1/sj0+UK+CCLTG6Wzp
BbJA0vD2FKWbAyVHUBqtpBpVZt7h2j5MshvaiQQ3NHbrbNItGF//fi7Cf/WjhBPR
3fVLJ86Jmir/oiIbCFDelAlq0WTIHrkFgzarYjyHemHsOB0mCEsx58VvzCV65xoX
9uEcMvPdH0eLcp0nmOYA9eeqbiuxTuI/U5k2TqcJh30iIR+fJFDU/64LrkMrmdKb
BpVCDc+eDIXt6UhTGowitOBWHkd91nWslBEqBztQX91Wqb7FbYCHhoCqV89Nh+Ul
FK+qkF9CSLwSSTemWonvhjS7sBKa1VYAjjcb1A4CzOI7/4Wze5njiqEVHjAqi73n
fQdrxwWo8c2sr2R/k6ChfbVe3xijqcHc3QliJK3H0VHI7vXPH5x252lDQQ7nEO4M
1tM/OIIBaFLsp/luusvSuT+1R8KgZnYkaxEp+HlSKbF13JxJURhccBvyPrI2bi19
1B+XUOs7dLpHiO1obLFlWewOLY2lVaGBG7Et/LB8Xv3NFB1h7RNFHWT7sc2WlSlK
PIGsKjjfRKlbfjuilj5yEZBvcGXWKubfZ8kQgxlw1u3SCbfOE+fG78pkXoQ8+C7M
0TqYgh7q3pdJ8i3+To4nUwvhTiBgrGp/RpN+aM0YbfvJJiC/e5YOx77C6bTSPv0G
NFmkSz/UaHpIfWSOHGWmpnKxix2JN7n/3F3y09vE5tS5XPNFH+2xBjvyLS8maT3V
OJgxAhtcNPzjaIw7zGTMLlCWyXYHrBWk5cbku+CyyjIzbBslPqYvqYK401gc1W7O
NqkY39CM4UiUZfKxRVq0t2GvXf6x5sG3oXD9FK1M0pfrrhVrvY3p2HEv+1eFMMMj
kyhq67JDvoCF1wOzWznHCeFJ02VseRrfXg5q1r17GphrlLIXijee9R5IAbnYrLJM
A2E/I8BidAcqnJgYtCYZJ4bh6dtmpy0U/3RVEA8edaTmuZDk4ixO0264Wv90Txf9
FYTpTSTJW5VIjG0pjXlTEkcAVJmiQAFOQbDCw+T7mzAUKX+BS24pfplAcp21hUEi
hWU9NL0C/ZQ4BV65YKhLUWWLyoEgXitdZXWmNqXAtE/48DztpJ8y8V1LlFhMHSHQ
vN1Axeeq6702/9FV5gnd7SN5O6lI0s9H/ZgEgC0a/tT1FKYRqhvKVgbLmOv+NVkw
aMfkZYCL44iA5CLTV6kJSOoN4wZwV93WaFnxAlwQvC3H/z/qVsiy2osLzvoS3n5w
2LKyN6FjbtoL3PWWzTnto8fy9u8uOTHvE7VNpP9q1D+H5VHvcXNDRCFjfQtxoNy3
9IvdYN1R93pBzY5U6T8AGfJB2Wpr9LCg+DGL7+VCQYQcr/nCHKSDFVag3vYfOlji
HT7DmFdyBzWk1LZkYSVAJQtNlCX0FN+5YRS/9KKGlBVFiXe8z7pr3jFoDlDzSrF4
3exZ//AdR2HLz4QKlYodTtK0N/tjIinO2exd6XLvKAe559FnV49SfyswwaBrvOCe
LEZPT9JsMvOnhw01THDSFOETHh+1wwjM7nFqBv//7vjoMJZCbPUZn3zTf+ur5DTM
x5iIPrRsB53h0B/waMXIB8wxd2OIW++Pt5xCpMQA55Egx9GmKQOeZpmEceXSbInq
U3V8NYGNS6RO0mfFjUiuGyL3RdCdis4k6BWlKPhlSaUY+/Yl6ADYZqT3kqxnS15O
CkPzNSjveJQqGxUxHBOTMn/vcaZEbY18u54Il8ohwpZ6AIkIDvjtoduk5dNmPRDH
WM88Pu7GKQNpID2VZOaCcPHgyhenn3qZl5ygkevAsDW8xzY+LMELWEgjyeKikO6q
gfjuGrWA4wpm7b58pAk2efaTkcu+rxa7t/t4DLpqkgcboO8ndtPX/ZyZn9ggwSDQ
3Rc9Mv6a1yfTuWlWXdhzrokYU3jUGfqJAlf23HwoIC7ZuZv8oZ63SghIVAyqL4oQ
niMhnlz/WykvT2Fncn7OnBcMvPMAg93rD42Qjs+lPJDfK2DaPfxSReY32wH30xtp
WE1U+Dw0CaiW9uMAo0pTl0T3/HZ/DlGru87dPCtlVXt+NKCvr9pG3wm7MDHYXJLc
CbHvgqDKI3fB1M2aj4SYia/f3+LL23NOwh1ZehCAF0+Y02KVdkeTvBRngI8M3EXB
1xV6Z+2kt5/Qe6H4uXPG6bbXkmHJkGnZKE0aUNH5rNidjjjM7urIQUrC3d3/fu3F
0Z7fI96TsIIDuEEJC3ULS5JsC1636/Sw6WwR30fzvYe7LnBbo3IeqAMHEAmBKMBM
qlZTmLGjDDytQAYGG30LI3E/7fM31kmwthOpatJaQPoZClmV6j8/jVlGN610MPhC
qRR5ppQEcq507DIAebzT8BHIZYsfwaT9Lt9CcflZR8185vjQvUdRMauRD33Z4AXD
8Ir+tGtow8f0lmmuhGrFeVZ50EHh7NfthKibQFVd7OMJ/yRtSwZR4k64vx1glUo4
HOS1Ulc6Bgxc8jeEW6DG+rXQlsRtNnMPDuO6Biae46m7n4+6VD5W1Z1hOMITBKaP
zJ/DPdGdIOm+zuPuxyY57+bnZbNXPvOcSYHr94XwXi4op2MdMAJ2O7bgoEBhPspR
oiGcdfrAh+A9o1uATP1VCCivqsNiA195kWLSqJADoVMaVILu3DIg36v5tY32CtmB
gAjJaOAayU7EwqXxWti2P/J6ED4XnjcDIZpQ6m4x9SWpoLZlOduFefQuQH4hdg8k
8BPOLpmmW7lSMYq+DekdK4Lb5y5wf5rZzLAQHBgxbzOQK6lv6N7ipfEKVD0toVJi
ZSsACczz0pvE9w9dIbbR9KHGtLofZVJ9v5hvLkolfwmr4KCP3cE0F9mELOYM2f19
494XbM7fFB3SDimeMZQ4BYmA10laqrtNcY2shdD1zpuYLe9JHzjh6TwMyuyVT8Ae
K2lR92WM6Ms+SmkbhFWAfbWazLIALIrm1A+iqEjCnjpdUUVb4xTd+Cl9wb9uebaw
Cg/zp40MRBfKWg5iBJPFGmfwVgb+ABCGWNa/Tob3gfCzXgYB0OkYQHdrWngJuDp4
umW9oCNMwOJKvJc5KQvZtIqy1dRcg5AR/N+tKkTEexq9NpTIlTSxNoHhrErBIiRD
Jh7sle/OPJG58B9FTKcexqsLdaHSRsPg1eL2t2w8EZa5imm48+ck7bRitbvXbUVQ
IoF8kKMPjNw3shexlXzUqBkMLhklLHxB6sVOsk3CX1ltxUExMwwVylI1uOnlmdVD
eI++FB5zxpHBhPzAtqOBKySm9dSHkqyJ+IDoEPeFoxJdCEWXOb9EbrKLcEPQbXgO
IN7LSB06VukjhmKTSFxKVdj24IIPy+FDvsXLfTsm16Juvzlb19K+WP3CuhUpi0z2
DD4R0RclvbrPbt4n2BzUrvsJ8OS6HotuW4FbbtRC7T45s5RI0kKMFe9LBxxCdIHl
nDE835YZT8nT3zJSK0Me9H8wOY9immSEelxbex2/AOGGZ58+rhMsrjWFnxkV/0Ya
3JHM4OZFIGe3YTFvPGagzoqaPIj8F8RhMGxmAYabCHPdAhJBiZULS7swFy27uRiK
YEqwDsgm+fukzbvEgi4Bea9ZPIYqipp52auRYF1ykF9gGf9zvXFDkl4tgBFAoZft
+KBF/CWwIdfqmwGVDIhbcfwWXNQsL6g1oBznB8GCB420K8lBVTwco2SuOOCKrRox
g7/py0ZFzVJyAe62vl6fJVL2vaa/1clQtza70MLmeadf3vc97OeHzb+lb4xBqOud
jhvbZdwUSi4FfrKhWqTMB9TAbTvpbmBwqfaabdCoSYJjpoiGABSmCHHrrstlttCb
q65Y0AhotUGsGV6FqxnK0Lcb4mDgawHTQmzUq098d7sS8hClYRPYgzFZzYw6ZRV0
fRWQcnyfJZ8GES+M/UnjG404LIoEspwJrYC3YET3Ji4UdGBluFTdODbUaPeqs8mv
8fkBgnuu1FJLG8F67ssuCjsdntekq5gB0sW/62UwT0r5shdZJCVE00bPSZ3GltJW
TKcBiGhJjUNjkTEK+KTlfhow2/MCHW5Ae+Dj+3D4OFWEv9/Y+IF7d6vVvzXwzoom
ETsjbxmOvpJOt4u+gYClCAEvzf9DY+EAHrsJH8OEEMzltSeYSoLiG1XBQtZRJTAy
HMPo3aRXZGIj/qxVvtsECASL13tmA701q13vYj2UZzDPHKx2HZsiCarnKLYOneva
jXiBvbspdit4LUGcDLcbh1zqOyCYFlTecZ9/XUrWrPeRDFL8H1m5RvK09ZclGKMz
VtErzkk6p5KYSpsgzM+5YDFUjYOkx1Rhl5U+h3z4aE0Ia7Ppwo+QYijsgZZr4QV6
bZQynf/R65Fud5t+TL0CEt9PYupsEaA4sBMyqRN21jqRIFFY63uIZcagAs+DN/O6
NMovxrPQPDvbG1XDq8uaQhTRvrBq/OhYgQqPNhew+HA5gDSsqJfwJW92IrcK9TaI
7GZjbYFZyte8P9yZRCtUlv0SeQPh+Hs5rxO4K/pZih710g3Vjy41632AvynqKxop
9ZqZ7JzFefs8yS6Y9yxAfPTcMyC5ABdEEyOISjK19wZASdn9FN4tzHgclwQnpwjI
akHq4whJ6npeTmc0PHkSLaBqrIPVuyvWa39oZpVnKkxBNbe762vQAJwI/1bQ2YjR
rtN5z+HZf7l0MwROlp6pyG7glrnWRXJ+uX1fi5ww8TRtOflhuECST9x9NRBOWW22
8qI9o7xns7/H2b1gDO+spAZFGdNK9cYx8HipQRwhFfQRTGk+J8DmYbppTSmTaTik
ISSFyPmhLxoRQIvy8aYOyvn8NChlJjcJjtpb1KoOqnpxr98Dg98PXcG533HH6dp3
F8/lmmQ+EfgaMgnjN5LshvsOWzIdmsLHf8hz/jWCJZq1ttcgywK6zWWqILoeEz+U
afcyWf5d12KFVN55O4QV4iaXbYQkJjpiwCcn8Xa/SrHBVJKnBw5dV0XwGHEbUd2T
QSo9LzO4ceYmnT2/JgcqMIwkfYphVzi7xVE2GK0wnSN2JRCBgiZFNQOslYZMLsIX
Zmm12IRzwJhLKzg1CO6vRWu4oz+ht3ctdEn0ZBM4tQfHLMYsOUMmnhjKCmZj5Zqx
VMqCpDZr8kHlyJdp2hGuud9DGL49CZ1Uwiq27ZOAoKDR/xBHK6/jiJI4NP/IyedD
nvWhLuR3x+Dzr6LC4dNjxg6B2SZrDI0FrzgzFbCXEF4Fz+SeMQ6Wtnsvwq7PHr+h
wqSO4/2aZnLtZM/FqJIncipvO7OPx7RUO6TEObqp9ceLCKxoyONynAblMO1LfOJc
hp9QNOa1OAYYK7MCrdnKTp2m6tteubEUjbjbvkjX/Gf1TtJUsuc6Iv7aXXko78/n
Shxl1xuyek5uamfk8f9PDA9nYLrsFXSyi/lham0sGC3ditvno5jHIie8ucBd+aEx
rmTUfRot9fpeamzYGfxDRQEYTEUSy2ifP1YTD3waUnIInT+xaLdW4d0lxnCGrC9k
UBFYJbqJzq9nTpGgavMNmvNjpJFOBGg8LoL2xBfW0lo5IjOPgIGjj2Is73RzXZzb
OFAgHMseo/kNmf0L/w0NDK1/BUCnrdsboSbbSAOGKrSZdkLF2Pwhp2U3lEW3f7IF
c2mOYJmNnALaY52LbLuhUAomV3Wr6WupqwCu9JnbQt8NfBx8sNPHkOT1cUbZvkTs
/FNBe79Mqi/NHH67upqKEHSllVU9+fKXzbZSDEtB0HtuXFMY61hMSQjiQfs2p+6N
Ao+35BGbI7Id6MLJLvqVvQ4r++RLWiepO6DCSrR4n25CqeGWw7vx96jMAbgSFln6
dLLH3E4mkTBxE0NyhfoBVoP/FLbLOvhOWQ1DC2nLTG4kGwHgvZ3CtFRs5nAwj8dU
wbAfaPFaayT9PM6RcDLhcWO+j/oiNJo8c0Cr96gity330jbatwVkIKc0S0fzGx6j
UVADv3FC+yDQKfq+BcVyzgdb9nFgX/FLhducDuhW/I9X8uMfml6PKsvLQ2/cD3kI
/3E+GnF8faStUTFNP7Lhf5yLp9bEp52mzoLtKzCqxkDcQypWqybFmcvQf4QwgO2q
mZX5AMRU0HhMK3rxK9yyLHtD7iIyZk5sN9qqAnxKhme2C0Ut4IgGBT3fAvRtgg6x
gvCy/66assvWk5mzRjrAU0AOkHzE9ZdpXb95j3JBLjnURYVGJ6f8iC/+QCQbzBy4
5HYB9SfcoriS5qGhLml2nyrRqdPfMSBmepiYJktADFJMvAAGvs/GQMtnGUCphzW7
l9MmmkBmf/sejRy6FOwWY3ORuI57PMAUItmYwkZK0wcUewjv0OhKX2lhKkMWXySO
ceaoInlhA+Ky+ciBi1DtcJkD45l9hAcu0HsZ6qKNkfIwJgjM+o0BxhDE8VohRK/X
PnyB3/nS3qMBYRkP/OpAB74q+5HOIVTWe20hJE9U0A7eqNY0O8tsr7098xXh3uLq
/MbNn2HmRqHomxZLq+6jDcvkSmA4+GYhMpPEoC6rSdsnHfXsdmbclfhsZZufuxU7
Hy3bv8+PUQvw+hvpDezhrtdRfMbFKglT6H3lGyIYnKQM85A9sxAoyUCZ+YSU6O2g
MHM067ia8HFNkR5em8mZKPLvthUQD+P8RG8oRbB0MAmFO6ww0mLnCjPz0Ek0D65e
kjd2JMtNLd3TweJeUNesj+pOTAbm0ibMx3W7qtZLXh1Qx7jLynRDIL0twHHIQM8q
wIRMgvdlkC7K92uosKIYnJXqheyDrBqcJfddUvNMEd0AX7Jm2KU0aVsDUxft7Ei+
Rotk+kRf6Y1JL4YVOCVxlnr42mdqEYsRXvxxDP2bjcz81v/N5g8p3pif/me8aV1Q
5ZC8ZekljYqPrryNYeaAXn88PYtAqQnRmx0fPIwVquJ2zxh+PYf2MPEfmn1PC65w
t7vnAvGCZWKgCpAmZ6HynmNuUuhJoX+oZnOh468yNxK9Y03zpNPCHGZ3UhCI4FGg
R4WmZtqlawZSYwK1I+5mOKCcVlNILIxKv1l/TLPda8llxTjIWwVJIAelWDXjXTnU
HWjZQxTb9xYOmtm8MWIgn8ptfJ7Dn9RaaBiHoTCizVGYF4isMwPKOlzXjMEvoulE
p6TZ69MG9kdg8PHCwcJnmUsnNYYG878hVG2TaoZ+KcDDFJmC3CkpCWy8F469pvpr
CaSRNWinYZwwJjja1ISjQ5tenQPBFHijZ81YPwnCqrrDUTB1FiQmWJvclZlc6V50
uYj0069b3Zb3HYm4DOPESBK5oYvnZ2kITqP8BWHv5HSjnf1ghViCOW+kJb9gZ4LM
9WRrRH9FsU2KPycmAqx+rpSeQ8rDym0nwVKMbfP8BPKihH8UnTfI7X7Ar2LuNum6
ukIj1aG8Tz32BdQJC4lMTPQDyvj/vs12u4kznbSqawAw1SjgcD62clePkgHOnfTk
qKWOrP40UgwbuNllZDkjf9llE7ExS0oEghPaFf2hmES93XGfyUFm5wyqKSzpRl9G
TdN9rPBxg/5ER6UbE3jSr7ZdAQNUfukgf//0TlTnc+i+N9YYy4/0D9f8px2yCzCQ
3sm6WrpFMl6GAnnjBAdeqA/kxa1fDTP8QDX4WXH4GIm1jTpNAcJ9czMN5d4FxbRq
Eh683bOG0Zuf/Z2S8VCxW81b9RhQ3bPzOUenXxUkU8fyr9KQocNaSASw6AeVR878
yjy/rG1EmUs0dffO/FlwxT+/1bQg19t7l+PCUx0ytlEZs9A1zVe4jn7ljOngI/CG
U+rRUo9G5aRqjNdGYV3kOgL0QAaXtUdWI7AUa3d+Hc0mdGtgYpF1E+mufznutgm6
yqP68RXdpIMQwp7P43UYor4uxWkwWKDi7ilIcnD8320vwgl1k0n8+H8hHI04ULPY
6ugguUDO6a3BRB0GA1ZTwlMqj8YsisWFeJsaBhalbnrOzagR4RUXf+yfV4MeeN4g
qMh6g5jK1pD2b73uA62RFTvAdNCipBXh+SIf3Xc797O1syFdYfiZe8TsqPB9vL2O
hGJtc48POcSEXOeWw7nf5MuBO6GasK40BOIm2aHoRT/oxhn8bKaIlMLXfxcC5AyN
ug2I7tL4YsugKoZrd4nNBUzlnQ9gjiohcBaymIP5jJB/R+wPY68Qwqre6Ij9KpsT
4SwyuPewXPvgHxmJlMGAdN33Tu7XMEJMzFDQYrEBLofiq0OKohI+r0kSehbINGYP
9kHXeEVlPmWAH1cHJX5sVFo/5HWr8LNge+OUG/As5U4pIVOt3GWZGlofye8y6dSw
J3je1sHYCYpaF+ftqgMG+sDiu/SrtGHTVWqsh4MyIAkme4ctU+2B9AYM9tWqctM/
oQxYc8su3RcNOpvA2ixT9aJDyNh08H7j/55kdME8/em8iXgQvWMLAcFD/amnYld1
S4ZjT4/xC+E4ahK77pcvuO+b43uNbcId/48xfFMxwp2NVYhB616Csxxg3hGcjY+p
HS1evMcUl2I6Ibs5sNMeU3HrhBJN2cyMMfiIXUMyI9y97m+p6f7OTvcFf8wy1PB0
0bPxok9ZT0wMWNTZM0T/F7hHUomfTQm/PP1OzCDx70x5nZ281i4qxVS2KvPdjZv5
7nsRCKOvYYRVHkg5yDlvdUcbcEcN+KtfpZQ/lhwXRNvNdmqUNHdoKJRH6eDmN+hI
yTGsv6aWfhgSECJttCyP7Fo6mYOi/jbxEZp8kgftdcdzZoiUQ7Z7CeHAlVl1Nyz5
bWW1HDrcHVfNSeNoq0kq02C3PEcWdCQYzq23n4024jC0PcL48VRrbb2/vOPuyAiA
FI/allY29Ycog+Fz/ST7zv4FLp1808LkgD7iDrrrj0h2gAKijYcvnpvuEz+dzY3Q
KZCisxvBQQpTD7QVnhlwsNvzHgTbkYEztn3pmJkygJmosiWlTEY4hSamLZft4h1x
/V+1crY3RFZW7b7g5WFxjL5tchAZeyQntops0QHo1MmAFME3n5SvkyOImNiUG2jB
4GxFzQfJuENK8qr87Xu62ZuarTTd8l/nAtgV8YNuud0uwozDseLkwLijow950abm
paabatVHuoasUwnNRAs1m8n0W57GQikCazIy2+kXZ6w0d9BtigjtuupsXTr5e++l
Axual6a/ZPZYaWcF+YsbsJkBnhWyu4ydUMKfbHN/u2DXP8FORM1DmsQqg4yjtXIx
V/ok8d7CRarI5BuNg0p9pW7KXWhy/bS+6jeH0fCypaCKtokosIciXGWwLFHROpUr
RPO+zWE0zaKNjSKpab+oRyiCVHgGNMvGeSoxp1w52/tEJ9GOZ30XFxim/f5M6onW
IC6uZ+gWfyQ9x2CT/Z/mgYp1secI8DbpjPSPdhwCyDpFPjZtDOkVys/XORimWNTe
eeZxFQLXora0Q92tpBNwXLAL4hDRwTWBM7zkq0OfRINmImbXS9D5kTbVR2n8SmKa
aYffb3B0Spc2lrAu8Un9j7ro60DBgI9NROJJ0uRngcZN2Xgnwu3NmqqYqZtKOOlh
AuqeL3LXiwlRgoWUa8+t0qaSfik373olEjuAlOEAgc48+akdheP2pL2fFkRXvu27
41DaOZsD2N2Id/Hoe+1zGcuhPOdT/+1Qk7ToW7a6ZRcXr4/RYzwtOPrDIc1RzmTm
UrulmU1ZBPnSiJFLdMmUHsZyzycTnkgw+hINQYbSGUWHW1get1XHK9WB7xG/i62+
gvUTw1zM0QGzmPQNiljUJ3cJA4lwSJT2CB2MrGL5jXYsfS+w2oHfmW9sy9qbnNLK
b0C1cTLmtCfHvs+Sc2qt0pqjpUZOofS+YrT0ZNWGzHluukmacUhH4s8esdvvOQ/I
N+exPcSAY1Sv9ngvXU+7CZuyLbl4ggWdW9BZZ5BSVdwT3MfKbrq7UtWSNVkkZxsH
GgREiIAfI+dwZY7N/GzbW+6PXZd2uccOSKolkuBT3iyzFmfaTDtPquH0PQ6TniRc
GY0jIk3bXyGk4W90RZ5G2mQqxsxKAtfRhwo90UBHE6fmer6SH4KS4KGG9Fbg1jWw
GGvWx9DwS5M3YWWNNbJq2TRWtZ8OjCATaCopiMMOl34lXCswSbm4YkkE+W3Rf69d
tKR41BEsYx0N29m9y3yZeRUpAemk86VlslGPzVkZZWdiW0kjTnOp7IdAgFi2+vm4
J88cAnAIAQyq9B5jK9ECVju+N3g1qaDEad60GSSFmXnFZE2AuhuHLbSZ/n9f6UCY
iKPN7QxOKeDuME7dzqKCmBdSPksYN52s/Wz0iHEiG/3q0iCLdoY1/nRAh5icIeCL
Rz9e0QPz/kNWj2zVwMNuSRo17K3gqucLaXkiF/MCSOc8xxG1ehAxRRydE/s5gU2z
Pnc0nJhIkL05kp6Bi+Y7D8KYaZPeBuFcEUoYqBmUUZJoBMQSTBuWDWVrsYFZhbfi
H/x7jykCDXh+eChqUTzAkCZ1Mfp1/oWtEiFhEvmHDGLjje2HJ1kLHFv+xqGYEW42
pEMIq8xuwM8MT5Ju61Glm2gQGeUZvyj+vKmaM01/pA69VPo83IQ2E1FMuGiVWs82
0XHdJwKIVk+KLHnkgyazBKJo3is1FxkRkrIFNyFgYaJCsMdAivWSb41S+yJDtJwx
XRCZjylgiRDC31H5xr2ZTf2pgKHcmZ9hq9VIIMyQClHMAqNmh78P0Bn+AoO9kQyF
vbngx/hUdGatov5bgaTIT7ABaKnXmc7n6EHP5aIiDBprN9J5NJbbLYsk2DbCxsgu
C4OpdnKE1JWsf5VoXQ08w/ALEKEMNaiSIr2yhtVRYFn23paP3JhOdvidoAjwSPcu
PdBIM6ll0MhGE6uwtvjkhksvtvXLcNBZed2e0C87QTktvtTiBFwNLefYuuknmfEp
ap45qMKxQBhpdWmpGmTBHhxteDDJRsZbyIUObYY3ALQv+H7ZKLHUpIl+Ase6xodc
HqE4IN9ddSaDnga/jqylB/Guu8bXzZ9vZRIWyMkKxxgvDt68uqX5U8ts+0jt4t9l
HggR4oZeDClr64A/1e4TF31Ub3U/1x48R2gY+u2KGmRTMI/U1lK+bPm9lXFLUPZj
z65duqIxCZOU5aKHGlfrghN4f7qW3LyR6ckZTIEuaLfiuNMraavUBMJ1oW74yS7h
AdzA2sMmUYMq1Fcm/ejTedno83zKyM5qCu0CKVBT0706yfoJNSUi73NXwCubInUi
qraycx1IZEt3IRZE0zmDIV2USJSGF5y6QdBU29qBGz0JK9zdbiSsMkELfTpMplyE
T7dxuiZXPyUMqbPBhuINeTSKt4jxITBQHzfYrp/JdXk7fggcKiJKbDrEsIYu4jjr
o0w6ilcxFNMpnSAX8CHj4Lq0s/qiX3WbEib+20Zqko9t34HZZcGs1agCjFcKdRbO
RkcOuqLQjDQhybgfXJTUDAa/7rLKe65QBGSSv8/3hnFuQQv/HacXdPtnjbZFTY36
ol5foLuAjjWdl7T3PylBYSt9fg6PktrVU9+s0vfQIk35BRt/6nEeXr1HxM/cUpki
rhrkm0RrlT1qs2FXdtHQOfU3Of7JME6ZOZySitiPNwFfupSrcGEy8fWGaEraNV/e
vV10ER5RE7P0Zpx3h3F55zv6RDg4imKIO8hTNJwiO+HBitKpbNHcus6wliRvoMoi
VSI/9oNTSVBtEyjTEN4LFMT7mCSQ8FI1dCTWBhemVwwYnKU7ukTuPyvFBib8xPUH
kCgvVnFSaTAteyZUz/H6Ng4amHmo73mQEUGWATcFhsTVtU7rZM2AS+eQDqPU7AD0
GCyxyp9M0NS4cSFt2L807tFYLD7KhPGuX5neH5maGWg+MYVHHvXLMLpQ/Qlc10JE
4qNv2e8Ctp+er9QJirhm8BvI8O88QcwJ/veKGzT/24KgspInGes7jvl3aGLLoWTQ
ljy4qr/nH6DHeCGTjfifVZRMoYLxpXWPG2GXq5NXRGV2nfStidqxHr3d7J+IabY6
kDUL6qQZ5mmDgmz1JC7K3IHknEWFuUqXWiGH35PhuxXtUrt3QzoQ93NklSp7R7sP
qHMIJ3SoP+55+3ah5U/FsQf8ro7AQ59H+duFmtMLWnLitwz/xduLvaXKP0492y7Y
LKSAZX7lETE0k39ODSw1nSLEdDoiuBSDtzJNeohNQdzNjXqplUUDmavrMsTRmONt
R2zXKqo+a6amTbBxp2XOEOhyHrtFPYqOAqOKcJlJOSY1QujZO66nwBBbQYfWfIdV
PUB2cM164TDb7afUzQk/iWR8dq8g9+tY55EDU2U6flymOk73s+iwyekAFSx5BNgN
DfFbGs4OqJTy+4/fyKMUs+yfwpOfP0FdLNOO/schqrlA5Hit1AgBnlxzl4hJn5yv
Zn1mHpF8jYJN8PXG1Hmko7hWMdnWstL6YY+EjfPWk1lEqADViBLmkdrqDhJ2Upvq
9NpUZZjg0Fnur3mnMhYb1dUiZ88c4mMXyrbRg+naF+JqrPG1s6YmrO0FgAEgCScE
aLZ8ymbnD+5lfCJNSaODJAkvT5OBBkoDmBAJH1dEDHh2nzVGQsoYV1wNd9z2rfbP
0R5R82AXgkxyuOeQcQgvzd1521H5xbQBa13i5BK5DBM4drsGUOCh0fHiSeIhpTbP
tuutFfXAhKoU/nDZjL0rmQO+IdzSgSqQ+h/YukwXZTuFg3wyrvqx7icSM64ktCOC
CE34qa0+SEnZw41ppFhUn3or7BoxqBz9dokrfq1a17hWv+D9enrZLfhNGTFybR9S
NSuZKg0WovfVFm1PMol5eOxvt3s1xqviEQceY3v73xD8/MelzSJhB/pkxi7OV159
sDmcvu8RtWI89R1s5W4jyzmY60CoeJBiesOkT89srEjGk07Aacuu3f/R+ZAv8eRt
pSq7q7sYdhSMt+3eJI3smNFPJF0ryeDIAo8YOia7JeOqI/vBWvqb5PHLyBA+dKoK
eBMjndvsSRtBA7KeT9evXsRQcCHh4atMxRdyjSbAw+2f4HcLE8lN/Mou5pKZH7X9
Kl79EZAga6IkqPXUt8l8sL0tzFHTfaFbGwomJ3mGlJaEI9o7HQnjXVbmtFb2MRmI
L5nHPQQIj9I0TdBDmTbjdCodgjeW2/z4TzCgIsa1PCMSI6GhnnRgRIk9+bznynMB
/r3X9is3lQd12fHK0FiVeY+l2/820uurhHa/EcsgJQG509x68FV8rDdYH/2BNxpC
4ruFX1TY3Y7FPE7fzH8uNM5G7lAKx/fpGxaNsrkOgjfcte8OJ2oojyotN3H5RuZ7
R6bYED9DbxzNwy8/0Y3SIyX1d5Zm81lb8QS9kd4oooJmiPdB/5tau/Y/njISYUTk
ifVtbM07oEVS2mwEDIH0AmsmvRf8sROAOm4XI908ZvaiUmZ5Hb7j1+08g7k3b5Yl
qk8YcAMjxmQjwJDXIU9r1P9HIxz6w9lnQBYZqsbIMIj+78p/WNS91m5h24BJUlnd
hHk6Y60BbWp/QiQGK8s/QlMj3RP8RLiDKoHdIIT4D+K5Gc3Gb8xA8MZZ+1NFAOFp
Kt/CHB7zExaXFqIXcHgqPJIGDoLYhNhZ41NSqZhtGf6x8jz+cq3G36HJDAY+X7pS
EEi+1DHQ+zpQT9V3gXUpItJsrf8czwaXiencE07WhQkR5hfpOTGYgImgtvINGhI6
RB5+4Q9r5IyJ+QI620Fi9IONumCqqThjRHvNJXqKhmaHzvnFF/mkymHJ67phtQ/8
YS+IWYPSwXJIqZ5kynZ1mPOOj1WUn7ns4TbAMbL30Ac9wKtlaEBLPWlHuZ+uUs2A
Oy4mI1NZYUhWEb739uuFr2K5suRFIs+VebTgdd3EsjRe9c4OAywf/+IdUpqj7bL0
tJPVFzcGYPe68H1Rr6bvX87fobu8ujHEjmdqC/jVW1cRwIrUysSkpfQ9VxaeVI3o
aEV654Fzqoe3oiDRmEBuTjFLPnKedReM29YnW2/CjOPF+GaWFAy9vv/N9cCTIPpw
jxao4v15ngB0VMLeKo2RPjExgw/K1xZyOmOaRP2aGO00wxt223HMXimyrOqnn97E
NR+fH6gwEVj0w14/BerxTyP/QQhkG9235vbsoqiQncOdXhiJN2NqGyBWC5P3VR0v
atVikpQL7rDgDtn0mLzqf63yRhaEo63cP2PwesaXnEgnP9zmd+bbNPZuwXkGOMcc
sScq4f1I50no7EOCYAlnpHU0RGXS/0w6atasz9Uob8AOX8WN8edhbBWmoJX7B7UD
WDfWtbONLk83x/fFNZBeLDLSfexnwnIKUq9PlRP1Ej+vxpjBzpK+UQ5L2YOKU147
cHvaNDXVyrLktnAwidddpPumxz2QiKzKhYL9WHK5TXuLCUfF4rnt8aij2XpuoDl8
jWGwhWf2t1thlG/EAr5uolgoiW4UCLL9wMHphS6zw6c6l4LPb3YSIvhKZBGr2iuD
9dfOLjcDIZElp6LLIY5dp5WABYYqbmviTauUjYfGHpz2GIiBJoHCzZtQQ1fbI1BP
suNm3ejhwi+05kjnbOpKfXfhJHg9tQ8SIJbFIGy8UvnpXQB7l1+mab5vJZZIZ0DT
i8YmswHBfgQeFv+UTEtLt2hCcrswJaSrBJGNWL0+lkyE78lAWfGMLLoAcXPkMIRR
hTf7VPtBDu+gJ3J2n3HHk4vlC4m87pPcjZDhzn+yXVXzK42Dahc7SeYErzoak/Rd
FzQqBYBTJlVzFdjqwW03d7Y3Tkv8ge8NnISrn+owGNgLC3Ux6kKlUuf1ub8g24Vi
t77OhPmKZKPu07fpHRId3itMn8oVKLgl1J18gfQ4Q8qJQDQMUD14HtexkIfjbpdd
h55ORknfIIGD8wgqzx5/ERPF/2v/hnSN0isDmk2qEQYu9e0RIqFJF+g8dMN+FzcX
nfflMEXgMCoFPl3sqytbPQbQfS0eDULDJedPMr+T9XX2oum4txpkPsnP9gAnw8kF
qobUAXva7Vl70VPzXLHay9jH3xY/uJfsyn5eL5+6K06BHKtDoGdloiOdY2KClmu7
DXFRCP12UPof7p4Ykr53JmiH9V6476eXw4Kcg8wUJ715HpOgQCtOA7QEGMxuhPJb
khkE1OPA2ypKcjr8tE0xGG/mQ1PEC6snDSeGqJOGbcpte+Ko2335Ggr7XoXsy8N8
/07BpHSB/xJd9QTLGs6vq9bpYLId8JrjGEkdRzqU5eH+pA1n7RY/83s5d8dptMG3
mLOYHxuJtvLXgU6y90aa5PmFD48/ahn0dtMLzQaiYDxEI5Y29Qowe9rJE/YRvJUM
jdCt9LXO/mzUG1EyK0WxwZ0lgetbtUTrEsXYMrTAy3MP5JPze0zUr9VZMOe84gK2
/KwNSlKU0V8WlB00N4reaGkzzazlPLIxPS8RB24s33dG5F6KlFNXG67/RNXhLND2
64EuezZ6KmmB93qlhjyxYzC+ZJCUE4RovkHsH2ACqmWTLwy+hESDJwZIT3FItBwr
sNlJJZeY4g8EV/T8PCdzsPd/IMhItei/q9v85V93diFF2UBTgZmUZJYu3wcn8yWD
4YVpe7tDHRKSNZABcGbCSLlBfi5jM7sEIXmhzgFN22daHZWe7T352jdGgXYn/mWQ
Cqkc/gcq7ZbeLCRyssvAx4yYyPU+UEy/GqsZz9M++2TfcOEvZhNRvfjqJZBojnoj
yhIfrOA8wzfl6ommRXse7j3gjEloChJJ5r7P4E5vZCJD4H19tebnfL4V+1j9H3Cw
YWy6cs/H3yLIDzrqo15HFucG2njckchATYZdbKQS4gKA52tEGyaUy9O09lyjnyLP
pAgjGzhZqB7EHo52fRFRl1KIUtqmnUlO6atxbri3gPXEt8/ko9zkhB1CTdYWfAZr
NTXGyh4ucCe8lO2GFxxDAbE+LZAduVL9qNEa36xDQq8jjpTqodsOwCXwGIKAMXgE
Z0vNfkWzBDjTjc0lKBnnGgtcqNUoS/PTqIq4ScXGgpiiYvw4WW8XUo/mQuAbnJQL
6D8gHEWIV6VwEPKURj4zCYkidzjaA5NqsC/vN2KpjwjLF0461xHJsNp9AKpxmY37
uoKBGgnUGUhYUAhbI+kI79mJJkwyI6PkTVpBC8+HUYJt9LShg9hrO2auw0BQljZE
5VmzcKDpRYOkpOIBzQXSfvB1DN1CPWevhEN7JE63stoVIXFOIINW2BAgQ4JOPfKc
5mZ+/0JFc6KRabkGZpY8UBJhf3/hcr/ZjnEN6kMFIvm6T/aQFaew/MWVF0cjV7qK
Kt8TCFBwd4epUGIoZuC06Y9ww8N1/h5QXMd2mmogzj3ZWhC89bplrXHT4KPIVIlI
1gYnHhq8g11Y9zlCPu3TQfAWnwO5wi+SemXYTmOkAr/YngLxwEZV0L0MCn78Prlm
tnfCfivKFOxpsvKbueztAEs6vGY0T010aY9YDOkywD8tgg/OyrW9m1B+9Xc59/KP
VLM8KySVjeLbZ7BlMaGOa/FdwTlBaL3+U8+NpaNu6Fjyc3JjBeB1SGpUbgp4yAdB
FBQZ+mDSL7xAl608kr00Ds3m/TZmUh8A/2Ip14WAn0COQ8Zk52k5xAVlVtL1/CD3
DSjQH5pUynhgTXqBfAGgO9gjur5pWzM8SCKqqriMWXtY5AGoGaRCC5gEnY3sKpxy
rPEt6EdP5GE4/XuniNEk3pvMYX/Beh7+ntTwaUpP/ZaOznYLcZAwN0H8vSYHcDaJ
/cIZUQ29uWD1TTNp7chRO9R6VyuNfAqX05DGJlAtksr+8sLKVOBQlILuL/wJFebs
sfVAdfFhEAmMjgsGqht76y5DIx7M1QPaEfE/yB8uMslowm/hspxC5d1m1Pp/2XoX
xl2cS8I0BLBuSkBl5TWqtRvB/GKxMuGB6za5Psp0ffLcfdPuLLoWUKazrwMFn9kK
oQKQUhKX14j+jVgB4Pc20SFGIkNBr7wPCacV6Y6okqobWn2avbOn+blm7bAkcy5Z
Yf4wudoXAtPAwdCRaNfuuoCJN6Qg5/3RkbGhZkZaiHvy7gAhsaJC/g98W3B9Yd+4
5LNh49lMS0STdE+jrtgNLAKF8isv4GaqNIUxBtZRH2I4rBd2kiLd+VYdhksQK9BI
Vp1nR9oW7QBvSnCF+5lxiQdc2uyZ0oEIyeNNzaguzDSF+frViUYCOMNdKN+I5C0T
3bYu1eXPPp611e/TpYR1swW7wK0vXqVTiHVcJfMOdOvxhoCe04Hte4TawbYJRlIx
BewUWAfIQqdMeoJGx6ZWNZ4m/TIgev06NI/kS7PStlSaLWPMHrcGJ7uPdfc4uFLe
6HmBjs4Q2l9yxDa+8aQaK71uTTfNAOsV/0RzyXMansC7ObEpBpFAUR2k6dPTceNJ
tGfzRnsDUPHYDor4JK4Wm9NsnzDp+Pab3p6rEqvg1g7stsKSidJrkzDcfqD72eF2
lrKTu3CcgjLuNtu4/HA6W6X3v5VtbCGJT51NglvAFr8jstLguylJMPRJ0xaZRQd8
UIbP1MJrbGvLAH7c0qcf8KPrJN2pDX4YN1/koHPVdQK5XJOC3sU4YlhAuY2b8A7D
x9wGp/q1TJNXTv54XSW2FngrloJU4PWeM2eQC5bArnBg+4V4DTVzwuHe+SxyQzQM
1oKlPvkTbLAYqrAe6RbzfNz+uWNz5IaG0SlnwIbqOPzPfPU0pBJTRr8l3QNhLqzF
T8zknmZK8Wgb0WUiohlphZ/X1tioYiyNiKdyJSceM3CPXmBrJHC8xAYLQZpICh0w
J24TMjNW8RNvUeAl4qpdm2xamjAw2h0XpSd+Kr5RtvT2A1EHeWUAGPlU03WoewW7
NSrG4/czz1CVNY6Xb5aU8gl1nR08vDMaRO9icz9A/3n1U+0jDafvcCp9dCTGkTuW
BwP5TzOHTwSlPi7GT5IfwjqrAIgftsVbViGXN5xiKoDqu5492xK1w3bCpslzxglU
t8xWfebUViQgfpnh0dXt6UV+VSWsOBMGJOrOifaW/ZvWlcytCjUPNNPiO3SQIyWs
flsGIToKGoFF+LuNTiPyvdZz9yq3XYKpq0/u71jeq7OQAuY/IBVDlPUqxqnZ1QK/
fq/8ev0++U2GUrwNq5Qnt51+PodeJVNKw8s2SxA/5geK9IpOKokLeNdfaS2CdFcX
yDoz7l+kQodoAmSSWAf7Hg7tfVuKfSAxT+vR3GrAklkQ0HGLNYEqvkc/qTWQRawf
6WLXPHlRtR0kjt3OGqjHtoLaj0uyXWoZD+AumaYmSVvqF+eq2UbwDem49HD/TBZu
skpDHlhNuNFSydAs/otBB55EhCK83y6cyZtNkbXabV3CobFWjBZuZZfHCkHCYlcn
SGMcRMZZwVt2bMvJ3Y5P9qdqMoN72o/xhJ+Zyg05uRyj9aRvz6R0bwTBA10bwbzD
oQHJEDiKLmUh8IAC0aVAhLrANoBJwi/3KqLcjKHw+uCK7CRfvt8o46k+3WhfWWmW
GIGAZNsDDXPzJFGKYusxbXgk/h8lbbiSUMhyZQ6i8KTpZ9pgzwyKBA1hLLAfBKMa
6t97xn1rSHFJiUMwG9IOXMd1s6yBekOlctjkVhkH6HjQ2GxSJq2Br9Pk8gW1YYIV
kNElsC1k7cVPtr0a/KnlMJm7aTtCZ1PmOECc6FrVujbtrQ27uydKACesXRcJN8Wy
4h1dgZlAJt+KkOGtsKLmzm1knZKKsTQAjOIcaF/O+1zqqqnOmhY6dWzgJ78rMQSI
H7wqe9rUzH99b4eQok5fRhFMbfQ56+Vn48hdxY+f9lNbQzHh8qPhJmUvcfJtwboo
VOvQPpbL5mjY4BTvhp0XKsMTDO01X8cfAAfIcoA72CDMdqmm3JQHRerimeqlM8PZ
D5ykpljT28+AZOl+bAU9QrAxtTZfYpweyy1HXJmAZmazGVgRKdBV3XXovI6YcSPw
wb9K/impSLRz7id7KAmveSt0NzlKt/axk6NiuLxarBkVicH2CjfuTf4ZrzZwT4+c
z6RV1CZpGyTBM1uiLWbWQgacscP/rn/uiDpTqCVD9pudZqbut4n/8IedPExzxhwG
SOOCN5bzYkBPAbZ7qHbr16He0sUF7sLk0V8VVGpCAHl333q5H1CCEZTmxHkp258X
KgEujSGT5wMl9EBbpwgV/PKHVrCvWGlBluH8WuS+EV807mrwH4YNVlZYivLR5t32
xUp6chWwonAgwY/haT6HGN5bwK8fq9jxT0u3gNpSVgVpw0KAUcJrxaUf8lWNQKEg
7fgWYL1npiuxMHkS8IR0tvkfAnxeCcxT4hgHeVfSnfMpGuVx7nNK/9wWv4419hPu
6WLpgWcJPQ+UUVvyy/nOODLfNmFcx9oiMDbVd+ETDf3dvT7TR8b7SMJDACfDoxSL
FjEBbNaeUmKIda7Li4K45YtRit8catg5kCQAASsKgbNUibA5ZqCDMMFv8hM3yo4U
njUrI7BKBdvy4yaedw5nZmY7x4L3vTKwHv7cxo/fQfIxIvIYj0ILYd+4Qbks7obk
9aCAv4eWXmsscP+X08o6zv2JwOsTrK7cNBlrTcWxU1ul56EG4Yf+5kNP7UxfO2pY
k1IdqR2k940rNHP3eb7OHiRx3LOg+bZHeOYiuz/OhmWlBcNRukA4oE9N4Gf/ZW6i
Hkg+H0abusZPdzopvQa1tlSpH5B93u4jWpYaV5+Xsw4lY1fI9UsC8/j1gCq2Eg4q
tvn+3Y39hN2ZvUkKCMm6QbIBVJv9hbKGFBCrV/zno4xLxKWDhYvofkR887w87ASX
+xAnwJDxHiWIDBnswq/jcLSKSdY/NxMN7Sntp3xA1/V1TFzgoZdSkYxv39Ue6JjE
r7d/eSZ1u3QkZ4TOo/Ru5N7rm1NDHjYXKO5rxKLJdY/XsxLGRAbSPpiHqEAao8wj
DPHQFxx8aVEs9vwnEQc0EPSDODUGDq7lXRm+ahF4E6IhL9GokTLIBqipB3CcKfmg
vAoxaSU/bOwRLCHYLBdWDgfs8R1k50dmoL8ST2jnNIfnpNqa52StR6JkjDWm4jMD
AUG08tnozOph4Cl8r6GZeJuO0QnlQTMaNKJtGDAHsLNQ3/fC9W2cg7nyaik5EYxG
6tOdLndd0LCJ9q085mXWJB4vcRfcYpI6wsxkUOuCukltJ3q747f4qmPXzaW2XrBA
ySmdIqqvTi0RQ1DmisnDJBp5V0lYf1fyV5oxCaTzh2wmaW2jwRgh7H8lGdfgz/4c
Cg+urtJesa8Nx0DxBkrg6uhzAbi1C2rUjOiJfHOFcbWEeWWdNVjUp2qHEVGVVjiB
lguuYkmacsyBv8RO0HXyxScmYBda5m+jikyMQp/ASzEw8DDb43uZdt7l+Ic3MQ0r
Uee4aVgllF19mbVIZYmIV5+N/7PeeLxtkZ+e7F7LFvXsO+TfYY6Y0W1Y7ICPYdOH
CV8e5rnWm3pMXJdO0URBbl1UEEyAL7XUnLsfTI8TJmIgmO+n40SznU0GY5dnkhty
fxyi6FCVDWd8xzyA1+CZbun65CjCN7rArIZBtgHveoonbOS6Yvyp0FK6Bjuzhh6A
rVOMUO/pKMp+IX3ZsNkYG620AMA88uYjeJXPbsDQg+Z6rp7O7JH+Hm6X/QFADysy
Q49ophL5lAEE2qtJaCiQkfoLAK5PC78s1beU/BnnN652NltfLZE49zucASkNoTu0
NwRcELR6pM/SXlChQ/xbg6NIOiVbNu0lIzbBT+Qafjg5Um5Kgl6jY0sYKjX2j+23
U707zjqb9t4tPqNOGybeX/WgYbGo0zgSVKDugR/d2uuFVEgl2uOkI46zH+GBmtBq
R6JJ8GrQx2o2llAznA0dyCpR8EOHdNfT1xPfvgsrEhHSAp2Gj9hhmpxOF4eRhLbb
/qrreIb+4a1POuNW/pJNs6D1n0JuCcEXOiDFrOXFJbEotAvrzno/UxTLWlNcy4Mq
5YWZLe3xyAD2GBIQGssxbDqZZOLOjmrZtlH2rVirUophuVq+wQzWkk6OGx8x7Bmv
f6o6QLzNlaAaLEhj4TQJkZs48+MJkje0FW3IGg3dqL+Ucd/pVvQHo01KgF8eorlv
jws14ziiKw9k4qHBG0hgNtZyH62yO3e80sRbXO+AxCa/4ZzOKYkCI3Jp/URbHvK9
xjLYsQjmmS5M7laDfFvCOhkAdvmBNeMBiwzSnhzsBNFXjX8h7LOKT0lLlUV3SeWP
uj7uKNE2uFRW0yyr088G+zY7tOSRL68mucUrnShPukV7Sl7vU1v46X/4gb0hAJ6a
357aCPI0fQEixtKM8IonyXMM7ILmV+teo7P7LmKPJNlovsT2zhs6nPuUKcW3c1Wc
tnmbMXpcqV9sEessttBuOzfUVBI+x74Cvg9QZwLSjDSSliIOgnpPuKthqiimEOx0
p9V0V+GylhgWwBeoB1bBRAlg3F9gsojxjCGuJZSNjyBTQ3d7tqObcxB/s9A9MYR1
6nsWjAp5z2WkDtgtraTJguZcGxp/8xWEczOHdI07y+6C4uF2vmvM8MZuad4rXa0A
8GrrtZ4GxX+dBYeVWFP1oUKX7cT8mutZLBrhEM8Es9alN7ZG84IkeUquAPFJvPZK
hw5WCRuM3YyC6R06b2y7bexV+NR9E+UG6hrWdZru7YD5pWN1lTp1DFO1I/Q1lpns
U1nFLj1k/otVAAa2uB7cz23YqEe2u7d9LzciUpJvosK7c75mTXvZRK8Iy9ooB5hF
VxssAtyhoYhv0Q3CYSs6g2CMY1AWYC+IBGmlgYAGOIuB+nKqKVma9uP88QZKQAaG
X4xZU32lewqMMzYdrPSvsKx8UoPqss1DTBurEVggXFM5rYZAnLUdZIwneOxQud/Z
jHsWWu2X1x01q2fSj6LcwYK/iQIjCbc0viefUj6mXgWPFiKfK8IEVjZ8b45F5VGc
up0arOA/hbiE14gpuZY5R/CJW/0DYEDcyt9AOIhWvHJL+J93aSz0gjwHuTr7q9bx
wYMrM5sezyKB1S/6WeLXE9Rg8WQHRX6s8Z08xUVqRgxdXozMv9eN204dwZEpWGON
fgmrX30VTCsshrLSR/VBVlK4trn99C2G0170mBQV8GYPXbS/WhVQ6DkHDbNkq2eJ
CbxQ6pdWvSdkjzK47LbDpClxvamXuDF3F0+e9CL6+0Z9uVgs7DelKqweajJ6Af1f
dYdrS53cC/zjtpeStk9ky7yGY0qKzyvpTlFNO59RkRk1ol6WyIZgE7pgtDKIpzpm
Iwxy7b9ZGszNdOJb28lcDDXWDPfiTrvazO7CguTFz1FnEUUbqrqnW2If2fsPaV+i
TRORpvwWUd9GNHGH+drVbyztVv19R2ubzydAoIcUei/8xuEAVWBYh/r6yl/rZkiU
DhARkuSH9mp+IYNhaoWeD5Il1Tjc+WXwkk1jZZgrr6i2ZhwigDWb6cmsw+o1yfC7
BzbXUOdej2hUS/+pQzB0cFn+GQyDF5repJ+/5JpdsD/r/PNIPD1xEQhvM8sEMgNV
kD3/9KojT3NQ1ahHZvl72JkfVcCs+Q2OHg7RxG/dvFHK9tPKEhEn0MQBWZjh6Ncj
vWY4hqhd+A7XNalshfPL7iXlnNsnqsX1bgFrU+QxvLIVr1GI7uI2agH/NSvhh8GC
7ZAzrjkbWChJrSRAGgp7jD6eHqn+8zoMw2OzVTyUyRRoLIBz1G9tCYOcqg/esfm3
P2A/mAiOE7BSyVHE8cfnX92Og6L5hc5gqXRtPf6h1CSX3wwymHthjf+9pfTRVkWp
53rH07RNjIKmrsW+wBmX4WzoxEAdKFTuef4yiZOFtJL7bcLzOeKwhZ74PQ3uFHCy
pL9d29GbxjfonI3nRHDgRQnA5eB7M9v1u6o6XzCKdNj0K36iaZFdUCLxO5J6SYmL
gdZMcCTpF/9yQ+cgT0GquhgQY/TxO+8RKXJZ1RbcQ/AZTEXmpnwzAyLkOh6SDb/Q
nlgguiDhAnrXPvlaWAlZg8Xlciuax+xL+hxJbYTh/Ly9w+ZQhAGhLVVwUrHUFLTk
2HWwi1DUaqaj813Ivc5VsMZsam49OOQgeKk70x/e9Q+JYTSNYDJKosrDxwx0p7YO
CBWdBC8Dm+BnY0fS1qE4gXqd5xfBjS+eazH6kSxAHZlLA2ybUs18nZkWSxrQpK+N
okGIgfHq/svNGILvlpPWqqsXC3VVhGjECTPqOxoKfq9Fu+fkE1DuI+pjVNKRfrio
0RX+o77aGncb7D/OaeIxmW2/QyZ8RB7Ssa7efPIqkQgLD2IGsMkevm45JiV2FQNp
L+CFtz/DyJjYEJZmp7DND1baksOVXAaw19Fb1AdAvWnGEDhSvfcuqMspmDSOMtO7
sQw7VSU0PkMEygCJbNSK4U6i5z6gFfqGSxI/T8622jDClyYTYG+60q/7TA3cOgGh
TeXR3sRZlVQnVWMycGXPjmQK9PeBItRw3ailmpO72Rzrc+0o/C7SDSSOpZHp0P6m
ivA+rjdmAXO4my+SQhFD4TNb8GXTcpUSpg9gfNvUZ6Si4ZfKrIRqTZ5N/ELIFJEg
3GSYDGWKdvgnlVbhGooItioID9RC4LpokNr3IdhWSYNHeZ+/6RCLXZPhyVhhW5pj
ZsmqOJ9+WkUd5Aqw/3Y5nG2GIHwQqb8WFq3a6csCRklDi3vqBBpqTU939mocDxeu
mm1DfXDK3gUSwB82a8y6fm88z36pCskvsUTnIo1qJnlRuJlerqGAaQgHVPWYnD03
F2tenmWM+xIVWENlKk3ewmKdJaMP6nUu2ZWd6ykjnW0wj1VJ6Kz4XR4oJR8UZ37N
Q3+4nIRUi0ifG4FFUzFwGNzyf172a2MGuaZDHwXxkQ00nIjlhg2oVeMOwP+UpM7K
0gKrx9aQjJhEDtrcwiOFZlVG5TE9AvtYbOlfjJNS5UciUZRvjqCJi0Z7QKOnmsLK
b0sqFO7Qii03bDrKU/BffoToa67LNhlthBMODEFaH8ybYd1NUYMrJcy843bO5Cr/
kDrzI9YYhotqfXX1dQTv/sHRqV7FIiEHEEZRojFa8PeUyELO+BOmpLduX5L/Li+R
o1DSWWgHJB+lAQKKWs6TymApVbPVpPs1rQ3aZ+X2IjHcK8aDzw+1Qsuyz2KAJZdR
0LF2XOgYzimOplN5YkjkauLGYq8cEAvpJqjG3sFN0LtKrD1GwCPVpo8dZ44qLKfc
lVkOLmDu29lIh8Img4gB+XcwpXCxuWrk5+1ebH3sdmYtLr+KnmBqeFHwWbPfdC24
e3JJaWxiKNRiCOnO5jE+6ftxEHvAonq4JIBkPIuXXVQJlvCTlOcgHTb9bH6cYck1
G/cA6eLfI3a54IOX1PR5+Ml9xotELfkv0GZxONTExfiMaGImiYkwNu5wSU3SxHhm
QPXI3POMNQ1QSSkxbAtJoO3E5Xqc+RBITayFCUhP8DB7vQ70NMbWKo+5tpsLJwzM
IXmrAQ0LbSGFJShfS+cSaIGn7NONiczWgW7SyT1dow71sHzGNxFX8iR25MFxy+mW
RAvkjjH1adQhWE1GOBtrleo5GTmsDD4cdI/SYD7JNoTBurYlzdEuYuUalS0LuAtB
4hS60Y1op1MGd2s8oZ9U6m25MpscWIpkIM8cPtjkL5Mx/LePAcIO+UeO6v7PW1nc
rrUIyyVBUKkXey9q51Eo6yZLFQw/76evU1goJlzWp1FlKYscUrOZ7/KjxwCQpfu8
s/2kz0fUi0iIIoMu0uBg//3+sd2+n3vO9lnq5pjiYj1PA9tILvtDa6AYRZPRyy7I
rctUAjOPdam+I0gvRRNH7JN2F3Pl+ZZdnAdvUfmb9cCnE4sf0LEd0c24SLKxaAqg
Yh6YyksewAU8PqsOuP1zEx0DiCGM3XOiCwPbOVi8PG9rZpPsdIzFa/Q4SrGJ6Yte
S0zesfYRn2RMGHl3m+H4DwHotj7sDa3t/WFFYiU+DjLhk1++XWxHgp74PFt+75Lu
8ohexYo1R0Cy2IfX1JFKWLT4ezkcICfqygl9AoLNAWsN7QeY6L+8R4t6pT/A511X
58HosjqnKpUXSbasnMDLCNrtLFM6a8rz3cOhyTHte25Uv/AuEg1IGg0YFdefKspc
Z6ulGaDQ9lhU+ij5NSTmcR1mW/DWLk6OFMC3Ef7h2yBIl9FQkYSy1Ugh0yCpJNrP
Yfd8y4PYvWg5dCFA6EixkLS5h75mQ+lpVtPtscfyyWqpBTrAGpzgzk/cjnOKlAyn
YV1sLenVOLzB2H+y5igHDGPf3tZMC4dpMbz3Qrlx6jcqiMaiJGTAs645LyUs6f1H
wz2JAWyvyV3P1oViSHPsZtyxauTVJMFl9LBx/xHBQ22g/DfIjFnwrqf7BiEHcc7S
3OPDJm8dMRB2sFTtIs7BmT/qjeDkVEGx7BonhBuLWfx9N0vPNdr+aDA6bPovDtGc
nHu7K78FvFjfENnag1oXEi4GFljwutLL+0AChjWV+WP0fAAZipbXZNHHFxRHphDT
Cp0hCBHg8gOdtUR1E+R1NIc4oIK+IMbuCxobmjXbHy5aLVye2FNK+5mXdvV+WQE3
x/gX0IBl8/Qd21ckmPbogpL+p0uyG8eQnbrK5zBk44sfap5qVAtgJf+05Q8/OhFm
6h28hzPUSe3xz6rx3E9goYOp8aRsgkhnhhgOebihfnFRVeXSQ06Ihn59K5MvZeRJ
E9C4L5INpNp3XTZzwqTGdfMsCTSRtKghd4HG8K4OAP2TvNxLngAGxzortVolOx8T
FwcCE5uz7g/+Ojyo6y4EVVR50Dsg8kFZF5wNUdILYJ0pwSOp8HKraFWDiG6QokqO
kVe8U/Xqz5symBUpFUwAdCRJ0bYEX4+XJAh49uet0F//GoR1jL8LECcYT87m00c1
/7fSZLYTxGZ8fYsP4NG0vcRYKgdYnlSy/aI3zijcTDxZCVNWWPrG7Abl0NQ6hOND
D61zSrlOFpExYGN+rTQUosgJKY8yjTcme8SCDCkBqdxau55nSi4Ge8hzm9cAyGpd
EnWJ8hYp7Es44dZT79ENFytE/XgcosA+D9MFnG3QGVO1R3aTBdj9FAnA9dfp9sTW
CLPgl5xTi+ce5lj/A2W6qlL0bvfcNqJE5hiM43VK8+PqCS1pM4MYWA6RFqSluq5U
zD37hybi19yq6vYZiqp7RLZr1IOdKY/6jizzA9K8i0b2Hj7VQni1PSznKH9shpMZ
E6ixq7CCvf91B0DQiJv3BgJxbnuiOaXOMiju0g0z0GOh+mESQVIhrCWbmwUP46x8
syZ/rTO0//sH7GyMH0ZAMuW6vrE/7uY/5Rlesp5YPE+wJMYD+9gl6SYfVN6gpYvH
f6Xc56nAvTxIn0anF/GMcLQcf6BfozMH3XBzKIgOEoIk49svJqds+4d8QdigaXr1
mRx8M3SOyG03D/bwr57blF3Z3S8Q5iDG7han93dI2yXh1lAT4UVQlnzrisfWhkWT
Fp0XRvs0enOBKYibuf6nQIfxgRNjRTvcs67LisJE62ym7w5uspw4xCKnuJg7CZfX
/Bsi2ZzJu8Q95MeLPyF9pberuyuJq9KcgkSOPDuk3d3n9wlHUZfA90fCQD8zmigU
cuO534ZzTWH8P1KQgFbakz7P/EM6pfVaBG/9GrLGHaQ4Cs+ZauXqvHCGLmqjLs4O
ou8VV765EhBjHyj4NP4dnIBuWRIlyKgAEfJRue+VF9GOa0H3adbO9UJOIDTvWTUJ
+DUeFtVvCJF66XTYJNQ/i62zw1y38584wuOJT8MvWfq89uuWJf/H+tk5A7iZ7ooR
hIwnz8D3NArTb6Ig0JtRqgQE3TTK1Qt1ApWMwahfdXTMyv2mvphze1PPyVmBbLDR
tYsS45cKuo4s8J2/J+vmYKvJg9ju7t1qbenosZ/7+fQ7Wwyg6V7iFZgQzViGe3kV
GS4oYHYT0nD/nTd1puEvy5Km2cmls5nIK/p9cUIjE54W/81zUdLkCSnPyyr29QLt
Ig/3fKF+ErRtkENNQvYmScsfnzXLRL0il/8cOcHkzV4+WYa/FH6w/Yig/BDjyU7Z
tfKur7bZteUPYoXGtJNq/sUYFr2p96FuyLI1pBMQs6p231CqeXcZga9Dfg7kWu+Z
uo+73cLzWh/S4trqCNwRenKz1P8QbYCqsjQQyzgKS138HzghrEMdPHapgWQnw3RC
oM53YuTT27u4/uJTg1uEanKnMCy4E3qWIFrg2firWGEy67NXg/fqMxJ2MbFkofrD
R7HeBLIqrxkETSuyGzf36Tplp7BAglLpJaItVTyYlHFFfdOP5f2wbgYUqNHjqfKX
kEdi10+r74frBh2vclaV1k45ge9P9v3Qrs4RRTOw/+iGJjH55DggzeGF4o2CLXBw
t5757g9MiVnI0Q7566L4L06h7fbysZuBmNpS9MNyDPeyg/jOKeYXiopLuS9xbECe
Y2Dt0LsE/bR5lubCMscQYjddiwtyuArBa6zRzntiC8YAs/njpyy9RWxhGasQAf+5
q+93h2eXOqscv35OQdOqaQa6CtzDO/HZf6rZ7v0FIsp7SSnw6gKT5YkNQvt9Rx4e
8c3LRGoqgT3V632bW/vwcaa7D4ZivNQxuofgIWyltGVEqELSoTGBiqGc6YWSGA7y
76+JQfJLBLKuEpLg8l3IUVp8ukt79kEraVWbR2KjRwfceJ690uHeF4BR4exVjMdq
KHFaMtp8pS8rF/4nRu15+UUL5aEaem23Hqa5gmlUS4lzLI3L7IB3/G8yzjs3Icmx
LBIHx3LN4q7AjiIe9OvpDRBzv1C0V9wbNaN6zCxY2GfgiKAa4kOOVGcsn4JDUrmn
n2+UstT8fp926I3/3rbIY04/stIFdLOeaLa0vpfuDUb7SykCgVb7TxpFMrvmJ3Fe
U0Ugyyn1fuGrwbW3F8DrA7LNaKR0U6gmnrI1abnH+rDxKZuQ2w+l3qN0y2/RaLeZ
+uAyc6Umul/CSe2hIM4I4HpgLL8J8Ll4x+SpO5glp1kQvWaO3j6R6HQys6gMc7/q
JE5NojeZ8FRS7JYm5gMl1nAcaZG6kHqfp+mKgO6s7OHYqs6d2wjawsGOspes891C
xRxUb271Qvy4lcTJi4QOLU/ERWA32H2LCdcUUQ8L3bWzA/0H4hiL4zwVtZJiVzk+
O5rf/HaHWaLM85n7vYZ2vAbvLdy0eHXG34iJBaOqEamxIgn2V1JHsmITV42R0c+r
F/eZhmReK7l1i+uK8tNkrkw3CoHTR+ylI0fHCRDZbkEkgGNw2HkDpWqugSqiKVIz
MOjndC9YCrKTmdZlKTsHaUYqkbwpsM9P+RgAuii1T3OjtzVC/+Fl2/Ji1yx0Mssr
JVgj7+ENwAmRfQrdF/r7NAFmjSXQLngISOqg5NkJtpYQMOT+OGdlsoUkOdqvMQpL
hiabPbRMxf3AzOblTxLuLUlx9toyyKr/z3JdyR7NS6+js7Rke3Rk8c3nskVibCNa
FqQZ6z+j62s2ovrwD0oURXqJPnAbAC6WPRF8IzlMvbLuPRwgyWqJskpJHGNZo4Wz
nQbv7HgZJt+SG9Ls8wj1pjMUCxlfB/LFgcDZCAKssb7vt720ziWcMchtJ6rcm3MH
vl6mpZyW0sedmMfB/7asrywhiDIW2+HOLRsGcx0OfjwDv0aH7rtVOFFdMVkuF3Li
ME5L70JvVn5D2rikWkXRheDW1qmt6v2WYDyIhAwt8ostUKn9x4aYOX/MvCNrHA2Y
oXA6c0BZFc5UVLBxixFAMXyV5hhkVeXp6+19r8kfi8AJa6V+ymPO/grGR6uIxj7L
59xwU63mB2yXt4N99pr9UiQZ7HEt+j/vWsMFa6ECTNR2gxz2wFCf3/s9mAduArRe
8F77aLJRnlUxc8az6Xs9levyr9Wm3iLd2tTyRdtujIBJjlpTOul9BFozQMN0dCWg
G9xTCekfVy7jz0VQq0kLnywnupXakcQ6dKhqSSrfV4JD4sxPiXdhooQQZ6t/ZsbZ
4mdKyLUsC1oFaCO4rAJlW4D1zcT70DDRZIbMrsX50sBp+LzyoGivQuYdh1s14Po6
5q3ObGtIQMnC+P/8MYY+HogoeDltfdS2FpFOGAV7mRLxbqeJyfTt5zV7WF7gZfkG
h5vA41P+QRETOD2s+5hNP+DgtXLot5d5zvFUS7aIM7iL0BC0jjsFu1JOI84vG6np
4Zbf4+BFWlbZhIJ8Cszv3mY74NaT/Fv7/IWUeiZTzzYt2rbYf9bWTfuARC/CzgqM
UBis4JoZBMlnx7OfAsclB7njqJMWCkS0z7kPQcJTX6GMAhXvCqWRp9Nui8fLmmCk
mCHJxfv+OAOA43eeaDgR5Df46xWre8V3omurWGb6GnzhThdJtpCP37GIJxSfVeGc
Oz3fuZDH90WKSc849gIJMcMnWXcG2uwq+6bt3Nf3jI1B/JG2uJ+Z3BvSjbrpgLbF
DogpcT8KB/iojd7e0bel0P5R0boMedtcwdTj5lZuQZc8ppEB2Tw9/MiOJ+hCZaJ0
QYZM1H1wbUVabsPPB8/FOQnfdQbr7CzRPJpPqGzoh5Ep00nFcUrhbrWb5E1LK6Mn
QwWylCeN1WrzEaiIrEB43KlLY5OnkX0EMV+zJphyMpph/+VO2m3DbvuiOFbVJK98
q+sIbY899KS99wX2azfB1smGNwgfbVIIEr/VNzDS9bBOMIRmhOi+kQ8vGkHsZl82
nbTOM0c9Nki4rtDd8Fa3+kcloHPb0+BqBMl081MJM1+EDEXUMHFZ0wbDvZU+MI32
g/waOpEEiRt84jF+lG8IqAwpGySNOtw7TpPWETCXiPPZgUWg/07w2COXS6JlsbR/
N5yeSlbSDZGm+RkVTr9ZYUVMao8wrZo7MEGQJWKs4p3eJqbdmFtiH68mcz0KncLj
o9QUi2QJH6ZzhcGXDv9hkjAZV2NRHs5kGyD8b1g77Sp7jYC8vNlQiafTPWFAuf8X
FvFs2DbezmcdtSUTorYs1U4Vdo9yiHi2c5/PHSi6OvHMu9wtcN74TAqfueChfL9L
do2EOajdvPZvCaQ140Y4e6pCd5ONsPi+tEs4/8XV810VPnRftunHKR/GO29YKEO/
Eie65FjQKWDeGY0Z1he+8PT6OlZRZGGa2rSH3ObrC6sGBfP7JH4NJoUYSBORobcX
FpJGSDj6jIATZFgPfLSJshvVr+AT0rnVh1Vbtx1bqVAgSJU0xdQx+E6O5JCcdGjU
E4b/mV4BpvchOtC0I69pZK3qX8nJIQsB9K936Pyc9gaRIxuxeMHwuzSxDdYAZh2X
xXpHy5JLJFO+uwhYMyjVmaWJtDjJqQbaMUqJ5MBuC0LWLytsgykG4sCXAzWMflCL
gNW49rI7oeu+EbG+lhRXYiH0rCbGqgPHUCGQHMDCpDy2KHMFwcO04xOIL3ohUI8l
6z+/KcPkIbN8EGMKxtOhLxg01FHFN0fsci0AOtz4jcFXM39JRIJk5xtOu424q8En
YmgZ03HW2qIfW6c/hUB3AKSeXVu5GEMnvBh8Z5PkQwoY/76Gw6aXZNJyRxB88yMu
vpMBQkpnhuVGNbHOB0fPJ7WwJFEPbEJXFBdX45mK7+XANafbXQPVvFM3K8KO1Ynl
CnPrU9A5krGVZQ+YnU1HhECh4PnjuF0oD1iCN6wBsZfTpHcym2+YIJ0dMQyrRthS
mFBZGa0xHYn8hPzC6D5lPY8XDFX9rlxByHxzvolHjnRnxJMz4RMxcdoIPJPgdTm3
RQXbxYruTYzdycQ3eQf1Cz6DvZJaxtyQ2pXgHoFSGOhPWh3vFPpP99AIyTU+4qnG
7KyYl608I8/PXiSXMc9/efw16dl2FccGhyVjdl3EzNGbu109DF7xCE4LP0ktWmiK
togudfExwsaue0x5lnzb1eypzBKzUnX34OXxalfoCaE3+Uc3B0SHkgdYM1hg94AZ
J4yFEIlSCMwpn5AKhN6WjwgsWs0b6rh4AxmM8L9LQMVHN8R4TQY4UTh7jqPbqjhj
oKnh+t3OcD6x/0duVaLNnvXjzWlScVHW60LcQ4CZgfhXYmSjXpobJSgWMXCkCyXR
zST8/yO5tvCn/bz21cJoPPxipMsZjocKCDF3+ahXXF8ElUSkZ44kBXvyEevwJd8i
vEs+p7WRFpkbqsmtsDnkUrBIFPVkl0BCpWH4KQA8IgjD+c0K+wtlfHfpu3CjOwS/
Zdouom5m/yHK/JL3Rv4NUFmDOxJpRU8xofTcjl2WKDJfC8lPwJR1r5W5edSQKJgs
HU+ZNAXuZDd7GThIOHoT9ZUemjTY/CEH2XEzq8swW4u5y/WHMR5+nvb5zB4Pi1xr
fHDXmi12dJVkgJYDMPsUT5I2dTGf46tIXk8kBW2emIVeaaiairKh55CtpztUZSHh
px+B6EGVoS3FZdAFVj1uEDY1wHc5QA0kcuAWsbsvzyxufjLidd2e/mRJj5tFvD/y
Ch3tJ3DH5cV9boIRUpP0Ux+LDwvJV9SrZNSm+IET1V+H2BftlW99rdDTUPkYE5j0
nKhjTuv0e13LOZP7GQJC0gt70GV03YuAexJ40qdSQqAw5m+fAJ9NQd4PkIvcQ08w
L/PBLB5MlqhKbTiELfLUG61IV3nsnJSCYn0V9W7RWshS6FdYGs3RVnbRKGEvqGtF
K9MxR94kA2d9gqAnWWj4neSDDaFqVCcPbU7/N87iKDwMy4q8pmQMvMekkfONrc4p
rwQAXRPH8EI57LM1XpWZN66O9p84prJ8MqWuZHg7s4JhwGUwQY1Vp+JWQdFWXZ5s
+vmMtjYDYSYAWWCUxzoC+1ZvqYfAryObm9kkCpExSwntS2d6j8u7iLRovOnLl/Cz
mwUkKRboGEstUHaUX5GqU6io8URxAVdyizaW4lVbIHnhm3fPS/nxm/fPg1apWgNE
zg044OhunQE4udrK84KOFmchX8bM9Hz6byGOXjbNRMGzFdHupI2AnFBhcLOZTIsU
o/tA3DKpD4m2HSwXSnlt4A30cL7nRh4QhCU1zyYV2LatO0x/PaTpYLOuJvxe26Ii
wbCHXX/f0/EHDgEg0L49ci684Qzh9oTljPiSHiHzT1ya1oxyD46SRowqCvAh+t5J
/dM4YzPLFD2TIju/w6auU6jYdJhgZKBT6H5uWkPgJOKpP+Gkud4kC5jUVfbAmJg7
eUoKvbzuIIGyJAps5Xo6hLQ6E3JFMZPDemSlIVxdOnldHnGuKZ3IR//8hWV3zp83
y+YYGPOFDMTQrzZbNuAoKGdvIVghs8xuAhHvdGCS7v3tYiDPyLPt6dji+WsuV0Q+
ChOl9kHvTALlgZItWloL6D8yfBmfv2FqJxU1s5KlyRL40j3H0S6Lmhv0m9BwmA2O
3fxA1UkTZEvO5bKcIIx0vpJ2UW1SkrCO19tQVt8IdpLbIud0m6yY2GJIQe0OPsCc
FJdrEi8O6KekHIpzMXF/AT434jZTwIuaaTQc58bhw/7nW2QD+TTcFp87rwHTt8xf
xucEwjhUJvArxVVC58l96/Y0w9cS0elS8uSQYQBKxfV5x+6OJM7wGdO6aAwYUTXc
fmDuR3clWu0jFzM4oOSnb4FEO3aHbKogp/X5TrCuAuW+U952sOLjauLYwf2HFPg8
YjRziOGy33yhXl8UqHi0/D8Jq9Fh/F0SS5fvsMlMH0GCbS3Tqd0KkyXqmPKLZ7A1
vHa6r1oCaL9hHKELBwVLgV/hse7vwVRIvG628okqjg4MXURNUQn1kPDf/cxWEhGD
DBJHfz8ODRwZ5sCXFauqk3In8KdGnqBrbTQNWOwvEilzMe8cyYnU6kWg3d03hChh
pHv/CrPjkBRlEhatOGuIWFAGG2FQdJZ/sGVZZeR7DvOsCAFKDpiNPU2bo8M1Dfkv
5stHhJaHe0CkbUGA1zR4JA3n1e2rswv+9kM+LS2RSFCLfRRmO71ipP80cxoHRjlu
0YhSWXExroqMSMFDCkfBBY2W0vqS/5RUNhGS0UFJ/NBitCOiTVza4eyN0ZQ5g+yQ
al0wmyNcoj2bEnIPIArbHKN79/0Ig5QiXwMhzJSYex7/2sjuQvk4g5gtSmQAoHr8
+VPVuhJUizURuII3ityS9tVNNpT6b9gii6myN9tjC5Y2aQUUdk4iT3gbUO3Q733M
gBVb2oRMI+kts5PxntwjLHlRCDk5CB9pFm1QuNA99oSMFRW7nYg14uQ2UcnLdHG5
8xqVd6jn/RdJABEGqpUlj3RjZ6eyTZf8mTEOs9vp/QKLcPlD9P8db7ukcKDHTa2l
NA+A2qY73a2TYX3XA6zdr9Km0d7wu6iT9KtgcJuVIee4cocJUDycs9glkH92vckn
Jv4SUS/ZUvyTwPNrTQvAbla1lskLFPvgVaoGWhe3ArKYgC8Nhez2H8yajtDi0yaK
2UQZHpyjSALyh+7Rwgaf+0Oh9X0ZXbw2FOJDAtmNOcaYBJlYUjqeAECZ4Bg1e869
eQWYF9i2EGH+w3o4/Ltr/9Aw8mSXGZuzJe2CZ2HLAb4nyxQ6dYPbavS6MGtfy+5U
6eOTkZGPkbmy0T6Y6G91T71Xmqt8TxBLRs2DvAzBBXLT3QNAGzjONaBiuB+Q7+yJ
NzGfn47BRsLDA9UPx343rX4lhQ6rcmvjHGQXykxU8qcQCZVLF0fNGgVUD6tVys3e
Tfz4Kwd40qnzyHI6+lk1nTsTaYhkrE4fUBdAv4jK84r+zrUuYSD/tjjbjfRJ6VGC
VvswQDy95sza99NIdMO5FMlIBIXML1Z1X7ZsxA56xq2G1GdgpbO2Z0Ha+jA6ZWEf
CxYDdAgjmrRQeVpsQBILsr9n2g5oraA/QYZ2qANsSpTTZ82OGo1JJCK9WK4UmOUh
ZWtM9vSUiPFsrfpvdne4hzgdgoCrb07+IU8gP3NZOjsotxFhUdQ/SZuhOkOH0JUB
UuvKygS8cTiHdeLoTED859GxuCMnnbmWTTC+grjzQaKCYEESTS/0DIoSge/Nygs6
eduOcRSnUNBdq+VAo3ILrAmhe5efN3UQkAR+n1giPJfkxgDvwN+AFF5TmpgeILBa
UONgClIgvi7BLnh/9+WfAS8qVhBqmTSinggfQ4uUDUSejv4lVTvk6mAXnedCY7za
Hwhs8H/1wBIevkkTCszCdje4i/XTXh8Bnnom+rbBiWBV34p+fOIsl2EMcUPRkVTf
l9vovgazFsOsg8I99xG7EHOnDuPDzcW1SsVP8dYVoCgM4MSQGgx5zc+xhGS8CI/6
XKGNX0LXgNLF3kmgKoMnCT1gKD5Fu2P8oUNzHHctj3OJVOwbNJc4HaX4eMyvkJ/L
+v89Fdrc6BHp+MasMH6ZdqXa9BcXXmEa/aaS3n92cmrxTm3cbA8Fj2FNl8Z3OmSV
PJcCOB2FVCJgDyIyVcqD2eTGUMAjuF9zwIUDOAIcRRFfhNlSsRjPLinbxolVGBBc
5hFAfL/ExV2zvzcJs+uh6GqaWrkutV7ul1PCwIPuH4TkYXttUJjIDOd3rCh9R2Z2
PmYvRM18pd/ZNHTrsJaaT3qZpcUv8+W5oUFuqxw9aNO43ElUdwvmuI7vxTJL7l++
EXrDnt4gaXiPMX4J/POagp+L6Sr17tXhPrA3sELkgcuxxOyrlbNNKWhtylxBd75D
Rr7GtczzNGHv6npFHegnRRGSF6s4vLnpcj0A0dM36EYuBkBbT76m3pP2r6qHG4pM
YYt3UTIb9WJVO+7nnUqDlu9L3EJxgfRHoeWgoIr7bnNlK5lkfQfViA6U3I76ZEem
vh4zBTjjIYZtf8N5rchzDte3o/eK599dvngPr4GSauyjxYp+j3OcSymd34PwM4S+
zxjbQAH2pLV8MXR0HtNHY04YnjJrPBXD5b2Ncw7L1qIkryMRBiX3uMUimEr9WkFd
KOL8Qc061yqfyLEpvN3cWpkG8Dg1Qi9wXh7EAiKjsgRTCSE1iB0ZlUmsjzQqv+YL
ELAQh+l8TJnKhr7+SP1Ep4r04db1BQZwjF3AQnTupcqPxFLKJ3Y3nhK2BK2/aBE3
5UTzV2UoztsZB9PJCHdZEkfm0o2mf/Q1E3qzzKs2FuAKorDV7SJuoJuZaVB05IEE
0yYfXQy7hQJB2dthJwYmavF9B7l/a3Ijpf3JjkHPOqOcwF5PePZ0zj3TploHrQtI
IdRbpSr49e5t8P3Af/kQVQ7yb1DpBQXFkyu8XGceHxfWtFO9004TdfJINsTBktZy
uzTfgFmlTPNPZf05BidA5/On9kMB5fLG2OLIhlwzNjw0rTcJX6XUCysovGDiDTP8
MVrtprX4JKlxBXFKgT+kiENAvp71DW99a0LKUQRJozhUCYcGT6ZrgjGCjcWuZ2DN
jyDQI4A3f151OXxnjx/G2i9+fx4ykBYiP8nJ9eYzy1GyThNxnKwNwTg/L/L6Fz3S
WiXQewgpJXmn7fKqBggbL2V5VZ4MahQ7+g/K6FwIh8eNqX1eDXr8Uz84BdtaG7s+
xtwWRxU/9b8lLWOYXUJl7iPhkBnKn45/+X+9gHxML+KysC6FQfO3+aFzuGi/U9E0
Dcm0g7V12ik8EuUNDBg36KTm7gcNVgtRJFojYczQOCVGiUKwu41UyGZkquj5UJ+S
zNBLyA/bZg4nzLfF4SxWKos3mxqpyr1w3QtC1Q4OexA81eavzoPpeWY/6mjZU6Vs
YSJs8/QcK0BnJqKlAlklV9jGGF0DsI8YxxuOVdvdbXPIyERGSmmRxQacCTfB1uE4
q/CsjtWOm8QC/90bi/exHLwpSdCtVXJ0HriCDgx+L11KvmELW08c2IClZh/Me6+N
nZvr47kiNo0S/t8VGegk0Iqj+JnaQfxQuNbBZqZmj+IpUWkPsLq2KVyq+k1jZ2Ul
T6vUUiO6fa9nHlIGIfTQ+5aM1C/33/KYbADvVo+Sllp/GargKNT7b4UTsX4Qvfv8
Ozgv+kZYTjT4x6hD3LuSiiQlT9lPSSgHDIs3ZfynVII8yMQbO92FbiRzn7Ms2xry
oIItsTu8vKdHsxxg9WWTm0FYs+kc7JUDE4kN5yAvRj9ROcdm1+kieHDuByCcKVkL
/AOyvqc7ZjEA3lCEos75dY86pb/MlaqvVbpmUwZlrR+K8FJklRgyGlYEqaUjnooD
/OLupKYKCNl0pkSSy+OJymhI/ZqgdMB4sksyCHs3R9llPIj9tJ5TrbCCH7e2aRrM
uQtcsBbfWTpLsRgbHFl7JbxaiPQTRGRiGvj6deHyGKTDEMq7HIANWcFFzhuk9Niz
RFQhvu+xufxhxPwN4iyuz/d001fgbCpnUPFzxQCY1M1lffo8C4zv6CWEPDQkh9SJ
VgAEhB7Leifud1w9YNskBzuKGHjeBaCcJUrkengKoJvQRPdNJ2jvy0Q7TtlmdZD8
feyvgpRf+GNad8B2TkfWSXoanUMns5q4YVVbYlP3ga/W3EPM8tZIC3NsNeMvxbVH
Q/Gqz5NhhIi0jNTrT0Eh1D0ryYqXlfHUjnanMc6f9pgpUB2nhI3CPGol6p76jcha
EPnRLdZ0nqroroapO4nTBUYR4WdmocQS/rk4GjfSGW5H6WuGVNpl+Tv8Kxlj5z3+
yGsQnki5cO5Q2UqS09UJhJ+tFWQ0ak4lPQura9+Z8CqSg5E4XKhHOWUE2jknXhRM
hCikOxzAnDp+sETQxlAchXM52O+iNOY4Gsf6msaUFh7CLoQDAlYNBRMBmy45ssD9
pr4w452Pc4Tij3LAHcT/M3XE5ZjCDaWJ6PfQY08Ee8bCFwp4U04dDaqsDm2rSx8q
tqCAGEgxJp+bTSyPy+E+HUpvY5ZrnKiMeZJdfbtOTH8i2NgnPA6wPTKBZgCudGYa
o2SP7BG7Udc+EEAsk47pzrs/4OeuY/KMlgWGA2gDfyrECWrmfWkwdPDK6LKuIO9t
h8LoWKZXHvBNnDf/gW98KN74kP3yz1rcfwA3kcMgOOC4u+Y77wyvWINzmoILqEx5
/e16yDsKfhtTP4mXfZtTunxd8j1pL7V2pdY7I8lLs6gM5vp3qG3dJbNMH171tq8L
Y3rwo6WBnGJCDd6OhAC4XtRdQ45jqzv227D6iIzQ0NaXZTMZ/QaZn9QPGZbAk0Pq
0cfsTTgpXlMxMFgWqcGqEnw9P3+n+z8YHtv2gUpHmyh0XhhQCsVwDJGJxKvipajf
xEn4KdL5xUVbqsTLzYtQcMqn9y9IgOSD2qQyRsnU0ocQwzA4SvbZ1a2A+QfY7NVj
0jRyWKXAV7k/CqH1O6TrJ7lm2JLWzmCORz0n7z3MHyuPV27gK4MxNiVkYihefiT0
yx1KdWrVHT8Hi0UKAgva4/Xub+Y2yD2StBQGds45PBgg1BkNEalVYN7WJW5qfQJ+
mfWqx0BXoqqu3Y2w/XHfxZ68ATxFuecT0RIKDUG1G+sOraABtyx/7dojOCsRVTWf
a+kwfQL+ctC5XAXF/vcHiLIAsNIDmM3MGShT1WmnjsIEEGoNtpxxGyXq8dfhgStn
1k4ujTLnQxKqc/MV00FBwBsC4HxmYGRlghcVgnFbDZ+oD50QEKlgu4AvooT9HZBg
x+3UFFvgIyqmkWVlik0TDJqcFVCsF7FwrhXPxbxeu/lqvdwxLeYhyuyERstJJ3Ui
IlwCzpXDeA2P0C475eBEHeyG9XKE9hvXsIPwHwwqW4PM25ZZ/xQf11OnlJkHOqra
WMXXZCrV4+tTH4LZwrDaOxrVoGPcmJmnRhYjMrBBVB5LADgzxWY35GY6Mp/K5cHe
iWEL3Nszskl/cwjbKVxxp1eD/+djo+7z0QusstDjqP0x20G38Cba38T4+YZ/3Cmg
GKlKbaa+JnCdPkY0Oak1yWbCO/z5igmhH+cA9iUh1ySrm8zsAI2qy32SFqsBTSwB
qDmEyzIYQp5f4A1k8LoOB1xthYD9viT9ZYppaS3qmmqpiKOoY0CqWZvykUCY0HGZ
QIMoRqm6KinPqW3qHrgxIMDiSZ3DplnZRq3b2zhjhAdNiD5zJsa5j59acGH0+S3v
GOoV8F6c8WlKG8n80NVIEx+4YQ6w6Tz966UDrDwbQzLMAnh16TqpY4QLZwDTiGcP
feF6DsISLhyancc4fvaB3ui3+mMciekNNB0duWruvzTTMeroUT7npdzDlyBbnZet
2dTdamKV1HbDP2aBHkqQMPowrCrqpsCyYIH7X9HrxMfUP4XZ8FggODaik3Nes4Km
h7sIppwkYssZhOW4gm01aVIjr291oljE8PAl4d9aY4fI7X1w0UtCs3+CTexFVvGa
3lMa7e+yDU24LH4cP9GI4AKCc+DRAdoj5bkSUypWcagOVUdj/gqQL0xX3ywITMzN
NQPXSxkDF033EHxbduT45B37G3O+hsTilyw79h6RrRJDUqN22BKT9PSkezW2pS9B
LuRSFbJ44Zi5kq5EnnqqdkD9vaFa28+dng9nwqFIRfNlJYlqLGwc+FDuKrDi0tqc
E9IzXA7/zeP7RyAWNg/eKvVRAGbtpkUpF5q45fxYeuzD+JMRbaqlMcqFEbDDB0ii
wntk68X7ZsjNhJ25DSuelfp4CD+JYQfQP2LzObnNFb9rK1S5gfwWGrh+Yo0dg77c
DOsMLXElBtuenPsIB86afat+uyxyC1EBkWUw8t81c0gncL6crAgdL5a3Jpa/P6Wh
3CLFnvhpi3oCz2KKkE6XCDQ/XxmFLbFnf+PSdRQWDPAcwOY1Pki5HR5TY7WWAUTT
hQ0zfrJbv3G7XQdXYPHaUtZnBi1YFlBrf6yXvUqsUvVzHOB8IvnRUDZfBz91dVOj
Qez30E7vhQKqHucpJfOfwt2MhqDpiQ2XkMWS1utPt3vZypjwcMir48o5Kk0Zskyu
IWq+sxt3NRsvnyxtXTUBPilL2j4E+V2uR9CpDnsB4SIgNdlxJt7Oe+6Ej8fyE4gT
muo18vfGDEuiVTfPtsYMRfg+ewfSwBm6hkokW3diOkkLk4zF4P2hLqFt2wyAwmJD
XGN+ViLUfnxFE3Wx74Su1VXWosDtcJInrzPTKhrzmkVimGR3Xb+LC2gcd+2DvrM7
kyisUSiZ5jZw6yerDp+ejEzMNwkEjzs2i1iMBYQTUbn8VeEkp7Sp6b3IXTDen+bO
MCtb10zeWXF9TMongmaRkYo1b7R8g2BmYnyA8e4+rIOblNBa0IGB7om1ZeD/MFuq
rBrmK3WEyguLcB4m249KNqRVCm4CT8HSO9SeUEVoAFzMQyhPk3PdLHLx7Zrp9gOo
MgraZuT2oCuDEyzG/TaEHpcCPYMySVHlqexsOlPmaMcZO1v9C6M5gORgTLOTLyIc
DrcYlS9ak8TVB49OdvmcE5aBnoKVy5vBurAAAQMho7jaFNladkWC3zl01ebUNteh
ZQCQL97CgmHCVlv+9F6I7Dwi3YztcBigEmQAfJN5pC+0mG5TWUL8PqTsH8Pi6Ieu
iGWrk78iP7AN0VENSKc4yDcOA+heImxAMOdSCBwyYGIsaYR9lLtDKi7IdMWOzSlP
1dL8ej9SFT7DwYQyC60u4uV9Ab7Fi9+S8HxjwMue08cwtnHd3qIpuOyMHuS6VpOw
Jn8271ND0AuoB2DhDzLyIAloIfjCUZgJHz/0pwySvN/po10TLBPmoW91WJuZ60lB
ehrVwVPSpwSpZXxHFCgOCjSWWrmja12YDBvVyI3Lu7v74DbfKX91FBbb5Ps+l61d
L6gBXMaLit+uBjr2mOZZV0Sk3s4VU3/HDAOFMRC52Oa+iNViexy231g1YQ+de1bp
wUmKGZg9V5F8YJ+uFpC//ZjKcP/OTTJNhqY+CIT57LWQJdLm7sGGRlpflYmhTdJS
NoeXcZ0VWvgcmJRNW6+BXNUsDr1nZJ7Ji+peyYsP4IkwF42XNRCtKXU0AfU3RKd7
xm11UtobYS2d+GLBUFFKiSC4BHJCQaSmrtIy0P7r7gO9F6d4wvQqmDmi6tEy8LTk
JPn6rdWBbqvrZ/dQ/g4fTgOCCv/DLuuP8gdw6hV9Qhh1qQ0jOM0jlGm0rGQHkif3
nBr90QZP6QtX4i95OHPHwJt8ZM8NGvvPAvj7TctiIVvjfaEZBn+2N9OXDomZT+zF
BOo8b82/BT2OTceoKjlX/OHCHlivxJuuS5NSm+zDyw8W2Xgffao++qseZG8PI0WW
kyppIyVceK+qx0zQKONuCNLxx32j0ajKf4FokoHurSi9a6k+UNAl+wumMsVcd/Ug
eXXVoIxraUpftTCUonRLCJP31Xsg3LYKOhIGPkX1d4EjzENy+vNTVQFC4p7aGCYy
GdTKY63XhxqctKO53FfieO1t97TmWnOGqUbqaMbRmASVhZ+b/w7OdrMT5jr4vsIr
RxYcHgxAswA/QfWPpv+4ITqTEoqi3Df21LQSMwqIy4CalyDIIVBt0TYf1wIWCDi6
ytsmqFUOpZm4DJe1no03jZyyDGs4F61aIb4NtRsy9l1fgNUsFjWFHyypc1RCdXc/
dUAbuXlGMVGJK2KRH3DlICR85wY3YHaHGPdK9n2aw81qbjaq3gv8M6KCm3CGjPuA
diYYyE7dbY0vXWq/BA4Jtu5RU28EPXBfUxmjiDqTp8j0HeX168I3Gji4973lt9/s
pf28G2Akkyt4nNVyksu9d6eF7/fmyIwGc8Q3tLNSlSXzET8P8rxqPyJHzcI4Tox0
Xk/BbZaxG2niCXjqfeBHLpdaK4zF58Rd+76TRJFV63VRxbSU4FHrYvDW/6wE3hxV
U/IU0RZEhqYUWXYpezINkGrm1big7sMW9EJS7dHJFBeUTrv3AIO3TM033X7GZxtj
y5blHXNgiXiUDhYqhCpSmzBPqXIW9SzkWBuxkMMBg7DI8wd92NVJkhYb8DvKJnyJ
i5cbVX4iuKxoJDM0v/EG/UcDQqh7NBChPOS5AYbTWDFeJdt20G4O61usKRIYHLvm
0KwhgKdyQj0qNLxNIba4Y70QSxawYTv9fQdSn1iqzom48KjY3O/P6Hfbw0BAq99c
YcZ6zaHJTVxbgXmQTEbF+wGaskHrdF6nOHcIGnjXTKH/3n1yY3FkZOVsa8/7xjII
AyCgrT3jys5nALVqk0Bubor1KDUMi5jfVLD1jpfKjhDQecL28q5p7CyjjyqpsyDw
rrfHrs5Wqbp+aoFnnGUzldjKX7R15pWS2PJ7N2R/ZAoDC8TXfB2y7Iyco2gdy1nP
J83E/hkSu0U3rymWQnE4W5EYag3jCa/Dmho5Zm+patpO6hrggt+Teram96GV3zIA
1qZYJwbJ6FRnvWHKNZ5bbE5MQUq5EYu/bT19o8lEP7RcLP+uv8xyDm8gBf2JZaWA
d3xv8HkMnPqGuvBK+msbCvEX9IDda2/nD6mVbvwrf/cyDzQv43wEWJBbwsEz6N3R
TTa9BN8ob/ep4sPQGelOKYl7qDedDpX2UtppZ8JjN/W5tSzkI1mlLj24yvy/bGFW
ZAcu3i8XAP772IAYU4dZ8R86xYwjhvtZAAjmkCOGNzYytTW5uoK4YnOh6zFPjyEy
0I8dCIw271O0j6xVCvXLA5TGQOEELjQyD75SSG9lD4tFwA4kRbzn5TwuDFVro/Zd
nHroNAJMHTajazMrrT4Fhj70r6K7/P/YKKaK7ZZTSirHkEgsx0bgwTBWtqE6jP4M
wh3M4Q0r+XYAbkReb1BDvR5721Q2FaPJ9nQ5nlpuAqJ0GrvDPP+hxU2RnhVaSaHQ
q4iwm8i6THPk4zftZbkQBu867GpRDbbEy0NNX5alWMUkVrktdqBHhpnIRS0BE3OF
MYLMtAXp5aVkwZ/KHBOloqie/jO2xuarDbACWdhicSWadQbHkw1PYOByJXrMOAU0
C1Axg45HpUxcf3MI1qBxvXusg5eWFjqkhLDU04pLQdYrkc04MSXuR6NY3aaAH6Te
sNV3ngqcE+zr+HYVrVOxytRVynrOVYWrMTv9iIqUehcChO8MGJZ8L8niKr3z31Ne
MQFDA73aBlpTT6g2ZixNuwztL1y6Fvk2NABeWLi/oWbjNS8DSnHIBshDy+f1yjDW
MOtPjZt/yaEhZnqCG46SCmCMAv54KuPvnnAyGw5cZ+KJCgZAOhA5ddeXahym4mlO
7J4lWboCxHNEFhkWW4A/B2+rmpnrXS2By6zOo6KcKErRDJHjgfv56X3QBj1CLnBY
IvgcttbKRhByQ/b43yK1r/iO3+PVz5qtSG7q2hVBZxVoNzcQGHfObS6vo29nUyN7
rTEIvVmoKlF6iGoJJ6hRbmkajRFFDCKsUh81/n8f4AGbAf1QR8YMqao/sc6J1zeF
H5UQkZSINXqwSJX1XiWQ0uAN3N+LNlqEeGDFOkU3P4GFch58eCsBR2T8wampTZc8
mbNfCxtjnx+sCO+WZUFguPOsnuj3MIjA6gtT+VmfMfwezIKMfr503MUqOesqcSEY
ShRSA51ymb3nYVf+DqYGhuUTsKG5wrPORhK1TIy4Zo6uAhrfxtwOICm7bB4GaFQ+
bNUOASQO1JFg8Vq7peykRph1ClrwWMA/MguHoaVSi9M0WmSyDJ0y7UjRbKZf2MUK
A4xdruhkrQCnu4CJIt0zAKKtOeV5sa+OzL4TjtznNCkRoGeVTPFMXgMlYa+iTo6N
I7rZZnygMYDoFgR4Bl+tPmt8UBa/hXlcY85JdIXqoCL9ivHjq3Krzi3yis1pSOSE
qYmZTHdpqpK8inc2KkR2vbcTqkDo1TxDrBuGI9UwlORV5wu1b0FIHScgwn6HdjUr
aNSdaFWudsPPVa97+pT+n24QOQYzYDKYlXnm+P+XTocftUpBh55GBBzfUS9yiGrP
2j5UUN8hdv+Pce24kiNg20qWtcfLknJ+NQv1/CIP/XDnqJ6PNHHz+hekyyzcpHuW
ziYCXWY3xR9qLh0YlGIukyK6I4pRjlvZAb4+Z71yrchqls8bxsTtkx7P5WTxfiIe
TUm9++bN0ib2o7a7nI1n5j/Gk6eq8muEj8HbIWo6hj2vGC0TnclfOqdyB3LdPFZ1
4BsEev0x5fSEkvScgyaxylwhfZo8HY6kZ33IjGOwve8efGKsugXWyVQJqo8W5Cz9
NhHVkeqzn/PbwzhnyMVITLwMuM6Wb96xhqP0CXGOyb13J14XyAkQXYKXKLnjGCEx
REU/5KD8o0E7AwXgVMnry0c0ORORSavJFNg7+2yXA5d45dt7PbL7CciBdS/1QJRq
AfNL+lNyJqijFux2XqO7DtQzgiSx4JmE7MBFIXRNkAlT7FO3Hzip2hZQQhRR0Q0l
vZAUflUW40Yfvrz6ZdZ9ZKOCkAFgfpaJHjvXF7FJMqs6xtNsHfDilnMC0H7oUpLt
MhslJYLTWy928UFJDnVFpEyYu85GRMa6CgwfCLr37V0rQV+8LOHNc7VD8iO+Vqyc
ukxKQ3Vktu2GPHcdMUzZDRFtFswfmSCfkOByE8KSVtHPDdwTbGpkDh3MR9F0bWaO
zcVkMqxLxiO8Hl/ENpyYCe64bgHgR3Z3XTtXcBF8u/ol9LCVzaX3Ykq8PcZMQyOz
gn53Ax3tKwi6yqQ5JK/JjzXkdysDNjNneNdKEwJ7Kj8w+ylc2Gz9UEuV/C8LjIZ6
Bntuz1w2C2XOxhZf+3IekHIP7IyIwO3/EMxcNDSHnnZEKdg7NrGyfP/cW5yDeoms
YIMtVJ4XxO84UqcL/MjWkxMvJYoDsBGB48PTcDilC2dyqUkFMeXZ/gj/PzkBSGrk
dhh7lpqnoaeObc8bN93q4SryKNpF4G9gN8RijyNKcAjiJkbdlj/MMLoTXs9Semxx
A+aXmxhFuTj5VqWrZqa1alcVzjwHbYXpdwssfUIUFdSoF+5yD40nMy4JG8OiJSeR
1uQRV4WafwgIRW9sBEcVdz3H4pcaytIu13LmFvADPz+3uIPc9id+sWWSYJTmXSnO
bi5RwAej+cG19MjXOlug31eCgH8BbpS9NtgFGZ8ZnqnQmZY+A+vtg+FHmqB0QXhm
wfn4G4+Cgpbz+7JpbTyHsAqmw9rixuo2eRjyBcW7CAvJSCIn9/ckG/LPJS32X5kY
gip8L+sA8pICYwcOvOEtb2D426UNHoiHIX1qBpQU7mvTBBL9In1ewnUUqWhSdWRY
JV7aYsZwHaxIursM9rGk6LjMfMWl329VLCHJa7GUz4ft7G5oqTAqeE4i3jdq3obn
qmKoVAnNxhsZiY2meAwwQcCBfkZuZhbIaRLiD50UvXmQoDBkTEFLtNFfFw2RcsWh
OW2wQRf62ahdIO8Nh/5soxhk7si8y5U5Obbzm2Xpn9YBCQU6OVHnMP3atEA7mA1y
M4E5YOTaYohWaZ7AlK3gN7ldtIEHXgf1r5rtGR/Vd+nSZbLHnb6m92SjnZDTWNed
hVjIlqeBwLpeNVV2pNwHjW/jGzN4RkLDJgJpLrs43i9pAOYctHnpfLFJSyoVxjk/
Qqdj5mHM0WZvjGbt36Nsjgf00ivbc2/w90/OjQLm59sC2ZuitG1bjxSVmpVB8K7S
QOG4gzSSM85LoMNTZiKVj2lwtoBlDde0WgJTNDXoJy0SJbwg45Ztzpmx3aGOByxp
c1ub7yjjuxAxCvZu7krsmm5iPsTF7h2kfdoi5VpuAtrPIlo0sfY91h9uI79tXzM6
AvGlTnCUGPGC0q6DsjwL+SC5JDEPOHLlN7NsIRQrgq8iFzH2d7DMEsnXCAjZQPFR
z4myU7OPDDzyaw9nHoXGVd1FxfE+37edaeAhCi7UaXDUwE1u0B9dcyXbF/AzwYej
4IP/Va7gAdmh5ooz/Hy3EbQSL884SUTLGWVIelMmmaK7Iv2iqdgED1Yvk6TdFwcy
CDdTlYVC1PZheFvh1UQVLe0qz8rE7LfQuQnMzpyWxepI3F0sLIZpirw+tmPRFVgl
iCkDhasC1Z69YKmlhEY2JE8bF51gbauUNiQlxfagyuLPCEoq75iEB2L1Siaig0UG
p3Q98RxabpD00Dr5Xq1GxHPhiJIUnWLXu/YjnIP039pVtl47t1IzaY9wVfAdZSLB
3Nx4gGzGc7ZuvwQeTahRCqeufUfZm170yse6DigbrouktvYpwL4lmwJmjEhyGmFh
zV2SPOaVFwm9bcxuvbJ6LUf+3jBUiz+lz6BHhLAjdX4OhMy89IdfLcyCv9TIkVHA
UzRUKOjcujyQdeahxx00tMmUz2QZoZlLDmAR3A8mqwJXta5FzW8ctd4vBtO7x+r/
JDqkRGClG8DDSOYr4kGFEKvCKjb8NGi8eqP94d+N2q3QNJxT95nvYfModmLTivqr
3/0NTQGx/ZmY7CXcVOyQjvbrlmkhT8CdDieuEE5SRGAIwyHaeGPFQcBe8oZnE92M
OXVtpNpEtOfrlsMR10MxkLRDeZgE9o5spTPx8sDeGQrxymv9S52daBEKlR7gXfy9
I0+OPAZ7mwn2Yg+iGY1+8d7nQr4tHtaBsYDk24Ak7pAb8uYzEbwo9eFja+7UdrRP
Azoj1mlIRDIlUYmwAqI02NY8kLZlVNSTEgqszIDgt/5RZY8k1CAhXHfIHLg7fB3i
Cgb+Gfg+F6Nqj92Gl4ZjBOHZYP+8n0xL40rQbUV+Zhggu3q6iQu7BM4UPh0g+e6H
kZe6PCHHioul3CpSAZuzr6XtfLqHD/bOpAl1ixnb6aNPuBopCFd7qh6CLUdUpHHn
QepNfISJ3my7xCEwqIJMYaf1w5e70Fa0uz5t91P4a+EteOyXEJzG+lxPq7YDYJlu
/oLs3424OpZBgC30MKHQTH5SgyMMysotWtYNlRa30lLmLeRSXvoiMu5DzE/UHCjW
OkJHwylu+ZtiY9w8enjoV/GfGOP07urBVKysvIoDBvCjUqS4oFO4Z1RaPfqnLT5y
EhZt3puFoHdDgHJr5twczMfokiJLl0ze/zFfw/NUD7yr2dsdUUkfqO8y7BqcJhQs
atHhU4hTxx5FvgElURXJEtWJAlzMhVp/LiD5ciF5Y12H2djOvLj/ZYn6FxR/5bzK
Xuo5qbQ2eePuVG++WZCF4PAot7nDuuuGoFp+bV31AIGm3eLmJI2jWvz0dWHM9b29
cG5+g5WftJN99C53+fI93NNRHPd6lh4onCaRdq2CQFldTlQqbSmTAAxMtuQoXv19
bVOjZGnBvPOxxK17F3iIK3fnkPFJgwrfCjUHt1MhvnPVpZywbTKRS5xamBPzVJQf
w9Ckyhq8QY7vKD/s9vxjv6bqm7BSU18PxSHFr7u+z/MWwCYAR8ZKXwYMbOzSETxV
BfI8B8OtyqKXdXNgwD+whmt+KXhQ+zzMkkrNNz/mi1hrh970IYJzX7jYdY8VZ/w7
LTE32lT0Ofcn+l7otQjZMyOc6hRERcYTkq2QR1ZAIhPr3AnGlfLrweQT57Yj1NJP
qfnplkmn7d9u8bq78TzSE/UT16xPA5352OnaunPTGP7aiGsu4ToBDghtTvVK7qwj
9j6bYAYTmOJR5Zw6hK+sKfa+22WNrDRJ8OG4wntfAXKcMtcsBJtaVpJS7cCqKZ8K
ZbttYhQqUWkb+JjRY1Yl3l7n+/Mixams2qFKpk4QaLl9vdbBy+WxxEY115fbA90q
l38ZYcSQFS0MlHcylWs5IZsMmpKGUjKlO0kUFyMIbyeECGYKp042MNngh7ZcU/4w
OR2iBjlV8oCo2KyBeb8EdBWu+w6RZnUHYlytAToa/Dtpz6Jl1B1LM/p2gM03olwh
z+DquZlVeeabmSSfX9oFMocloMphedScH0wLsnEBe2Mn2XMuVoVLY5YlfkajyCv4
qSPzF2ggxt1aENdlsb4Dgl2OmuSop5QhdZ4pOaJO0aDxNhpZVVxYKx3c1FoJhwbw
dfkR9oLMSFy+NnEpo4L/EzhrDCL5usKXwqUy4FUL25y1CVd5PKy+DhF9ToCuxZ0b
lzAbmzB6zdQ6IdDptb71JZ8p9mCi3G/uP1Yvz5E6282aUv7kp7vqw5DgLIkqU2Tu
2jnxdgNdI2ltc6nT5DKoSr4ye93HqF0V3kzomgnK1ybi/yG0EgXmdVxIL6bJ3zht
umo5bM2HH4CGzO3EDgo15Mhaggo7FcVi3ZuVcq3MxL8hDRWfYvPtH4bXtm9wqI9I
vphXTJjbbfBqcUGRpgNWeb8y7SNaUBUT79gKRdEziQJzodVnWUJROBufdmoHIjTB
ldDVxQV1fzOVVOisMq/dy9vVPaJGpN9uu1vn9hvF1D4g+3KuFZitubyfGaK8PWVb
20CjWNYxuR0EWvt/xoMEbxeidlOmiFOd3mIITFeIbK3sDgMZZa+YgrQRTaWSqOsY
e7vdgJsQlvsZRI/y912RsXCirt3iLUMtUMOoizkz+kidCxs1r7GWtngDQUhCftUQ
5LGGFznCmlZX7gcashJOciYH3k5aXnbliWpC6jLWlwpGPNXhK/6NwjgncD3mDv/W
pUIe5knWPnPAg4e7DSekd0iT66UU7abYjCsztq+Gbf4I9GlWGEmffUZh5IXOBJik
8KsAhTfPuYBldovBjrOxGRBl/r6IKPeI5rJFFdAwG5fqP+mhTd1xyZ+RBZBjCt+L
MhlJJf9pIMN2UXfAmwjNJmPscf+cPp33EA2m9eOwkaGJGNGGr2qR8HLSz4aAnieg
5jdhZDI1LSU3IYR7upMB0J6c022cwr9QyBE/L3xe7W0ckupSxGVEH9rb4B3rA58l
hp1CE/JbtaM9P+IfGEzOPVqDwQz9PWpNGsts685Xu4KKXvZikm/3kgdHZDIr3uD1
BuLaerWPMM7yr4sZnjqeoYET3leAfx+/0x22CNEipNbyvxs+YO1t5IWzkD9IodpE
r1DN5mKg3Wx8OEzkygBsedjvgOa4sH925gb6+SR27brCYCUOqk3A3+ivvKF5Dl2z
ek+Chmep2W38I1O1SHX/xpF4WTtdHc1HqZy8wo4scM+4s1gJGGbbOrT67pLjdDI1
bckMLznRCZLJE/DcfV3j69pEb8q/blw/SfF1WPsR962H4Cvvr3CNbuVwBeu/cvpT
VFDZM0DIsQZykzzDRNYZgBF72/SvQspZrkE6DBXRD+YsBcINHytsHM/LBZ6l9lpO
d6ezUd+r3WZtgThyyWXTRapJlSLGY+2ck5l3CB6sCIvX8W1VAnWb51tOnZra5A5t
jvEADl1xuu/wUIz34PrCntqoLhxl5wgBLOGqkU5I0D5oODcSRtuOCOYpVoTr3R8X
WB2RpW+eBRXIg0O86exoCB7SQdRTcPGjfJ65RXmthfHVlyOf1FFnzRrFb2BYw6ci
cf0wb8OqbhE1CsK4MnbCVmijRU/LiR7byaMF/LeQq9CNFShlpy8lDhO3Y+/qicw7
RiPhBh6gvEdEie4fR/XYKvbDMzq2BAMVZmLUwAncYDTHyf67YcOiu4rqLATBtZxK
DAMZZMBuwSx+iX70fZWZbbecaJ6dehxq5hdIv/rYqI8MmnPdC/YNdBUxoh9GPzc1
Carl41A1GQCQyTPNDXcfjRPDDWJgMc7cfhlKLcJIY+khYFsX0S4bQ9yz9XFtEl5H
PpPVMHaCleZSnkDWU0tRTNLdXv3rA/V35G81uQhoTXEADZ5Wx11orWSk7is05dwX
+024BqvOrAJrjFrJdMzqZMPF2zuB5dVJe36oGnFqMifVmxGA9iFmxXgsKSrFZPO+
SH/cv0uhHnoo/Tg2Otnef21xvZE1LZncDm8uX+EiPtXrfpZVGkjD3Zc/bPFCBkZk
TNPNz3yc6QQOs/TyJD7zKMSw8G3auxiYRKT/DDTksNgRkRRJZdpiccz55XZ2VFlV
4VhTTCECXHIMiLk9LJ8DQtpQh7zmWOpSIAYDmpzm9VatIjH4IVxz2wxfz8lhVjnl
dg46e2mouYIQUZXrYXYIHKs+gZtGxKJqF5vgFAu1hCGK35xLS9aM59JnxYc2CAgh
tOZ+LJ7bOIs+UgNdRMIq2eJXT4xkUEmByZcuIf4a+Lg3i8NAqPJJQYusvEgdrL4x
1yr4pEVlW3nFhRWzZoCE+KKlbk4idYbgMFdO5R/mA9O6rALyn0vmWqel+edJVBQC
fpCIOkZ5ibk9YgiuKVH1NssLQdBxA2oijC54aJ2B4L3V1iGgvIeSj6E5u5DkNqDt
q2qvyAa/Epw33lw48Kp16ASlFE0u4PDsAh1EwHe56N8le7XGlGfrCrDyb/8FQfXE
ZVbsqcb//sXwi2EVncSd8Rudj48WpxfRmGG5+E9WAndwdUzC51epkfKCjxuE28r/
fc4jvD+OHk2V90IJUeW4Yn/B5ZBUG0gQUxRcztnLu81UmHHzRmXg6K5h01EnjOdy
1nSCPQoNKWWQgKZ3yJZwkxDwPfw6qVrloj4k75LBfdDlPlzGiU29S4qyxjo5trI0
GizIdo3mhP3GuB7SKTOQnJvK7f5JRr5JfI0/yEPuX86D5+BH2nOuuYyxhhe1T0PN
dQcfZPpRfdgZ+gifBOq8O274sq1W04CdZgK/fxxOvYUqlAhWg0sUQTOtyLr8JWk0
6TPFogvXCebvW69yC+5OfQ0DPM3Xk9bEC44i5LSRl+6KT1u6M0juZGrKolha0qyV
mVxR66G7M7BAkMLSoH15eOf+rkaCvy+Ap7w5StMFMGXs2OvshRLqz2sH8yS8Ggef
8XZYKSDBQbpMp2H/xv2JHmjAC6hjjvMIs7aODtbOxupKOEvbsWXYXPwzaljiwqNI
Qd0ehwEtFYUBI0Qqu4yIi9CobyfyKLqfex5Iijho+F4EowXBstSz93R42E2sK7yK
PEmMKfwEWZRBwEFEigoDCXoZgwRSXXKMVVgcYaIEIqtoOEj/ytFPXBMINFU26jAJ
mVpvctrQIglECvzPtRRkVsPoCaRjOXgLlzrrMa0VkP2DTqOK+R7zuVhhdftKSty1
68vkH+pP9j8YIjTfcY5t5UxdVid4fs4sFnRUzPa5u29WevlV6Jn8Ubu3/pblG9wp
28xFGJHw5KbyA7Db7MDDKyuFMXPHQ1Bu8zRc5KLQO8/fqIdAzo+cJ9CbgYWBDDDI
RuAI5P1QGd42cqjWNB/RREt1BUcS+OdEgLjWMPqpGYoc9ryt8Gpxe/2MqvSsg7yF
/8mqs4PlH0yNnpLgDm79/HSQlriW4wYs/YSznzx9+bWmLFoDiAh903rq7BBY68WS
QgosSe1t3g2vE6EkyvpBXAiVILlGEv6XuPnR3bEy3WkT0ZfpX6ToCtYW798gpQRP
5OL5lVBv62qyceJ+3lb5xTg03OwAc6WJSKPRTp3qH72Y/451I//DFwCxnJH6RShT
XvwuwoGEmCkrvmSPG/SXbEq9iTYLtu2G1PxLHmTaDshZLZFcXbqByKI/X6XaddfR
Mx17hqb5ASxwZP5QkyuT6u7RP1uCJS7Gn614AMgKKa826m+Pq95JuSv5AsEXT4DR
j67S1A492lEfWgM33RKFc+vD4HI8/5559R30N6N/nFARrub7jKSHtXMe6z6Chf5n
JbnURkagTgV+aYzVg/6jcfYAvpaIUWkzWmL9dBKrkkx+ynMBm5U9SzWjI5DxrTxY
k+aiuOhcC1NhAUy8x/iw/XFvTtNp3HlAiera5C+3qPT6mCjCZ2Qmj5k2HSZiXeA6
pNlk9S7Vc24uNe5h91EX62E78JG9QehJUFriv/TioBxtlDbB4at0E76bB6D78ugY
QUw95pPeY8m5dZAWe574pFGGICkfKF3kmQ/7SudyLDgz1G2g+UpFQE02YW0/Hg+3
gt23cvL+BVwiDZQJooNfr2pOfv2Y2N5hvM4s8j/oQOL12fpJsEnNs+bTFxs5dHJG
Svnpc4v5KZ9+TtDaH87LSfQhJ/szMKETPBZ3G33ZJtS7TuRAZzIc52fE6adgJgWl
4m1xUwTheohBRLWU4E7sLZGwy/wQc6NkS/jVZ9LQFNHCxfUW1DqgWSwa/BPaOZpr
5/UHDNV6uc79aYJzw4wg/LCm287lcoE7SqiOSzWqTpuMRK3ypQwPPJs7DruZGEVY
zQFaeyeR98QuHvaHTVaWNJDBZC7gOw7oCtbj0WrgOF/trSwvwjaMxsGfRIjASgS8
9Xnb4IoPCcpgRGakw9S9ojBKMhMe06fyRdHOedZr+dNTAi+2hG4rBmIjLnOUiHVP
7i8dn5VdsSooVwcNwXrwWAjyTEvYOVmDwaq0XBIMNgd5vivnOAri93cb2obFXmoQ
dUkbm0tkFFGes/ucNg6xruMyEGsmC0xiNAXQ8Ef6chOg/4p+JMvjBnxsRFGGgOe8
mqzUnUhzs6iHuebiYqC3snnIfjvgiDZtRjUdZ3LruSmGxoycwOYQiGBA8AcCSTZy
vfrXv5aAig9fld6CJTCFdLM5G+dfUe1IE3eYrX5qCpsFGQWyU/MSKiYXnt60Xd52
wIW0Fyz6ng+Tu15bcOZ/gm0pG8ajveCzl0nEq+agb3RaUZjm5ieWShpoVq2xRGy+
aaC339LyQiUxwCxgCKsh8jBOXGkyvFTqJnhpo7dMfbO3OPYSIDCOIhkhuCwyCYQy
Sw/p6PE8yI3Yv8QwZgO/3mRyjLL1wqU4s8j9OVpnkS5tGvO4UD8PYXbTxoyJEHWZ
iexbd8lowaE1DSe3nMh3QCu6k9MN7P17d0x65Fw7H74Vzcla4eNn/sxlk4rYWMdX
lny/aBSYa36Iq+YabVPB5Wn9dySPvkz1EeY4hCe27BRc2nVuKZZL9r8MNko46MlS
dhtKGSIuO08orDhXNwMnK+86Vo8mrRg2XXfAfGPeK6282WDSJrJdOyjCRqvddlzD
pVaBh3S9OV/hhBHpWvhkj69Nf3/RWhVZAm648r8yY2CthTTBrvSDLp09EPh3PsUY
0lxQmmN9V/vkB8q6qPn8CB+/sBRjT4Q4WvUkkDc6Oehn+sFVJ16j1q96BiLjmDOI
uo/ySajQlQieouVCsOppQPZjDUxXOluYu9w+sugypB1ByIP2of7OxRADPYK9hnWB
IfSCmWrdlbL5ivkXNIvV8mfCGcgBocsmaGsjGVYGBVo3JMOn4P7dHhuKS/dRaO4f
Eulz69TCe0dryjM0vFLqwDaJwHYotS0MgjwAXI1qwa3LbUGrSZNxpNQYJJmQUodi
sADEpklFe3eiybthU9ToR2IdZ8VuGYoZra7yjf13B/82NR7k5R4Tz/e4Ye19tggG
k3Z9AYOaWLCb9Nb91D70IG1Y8bO6COItXUCDqCdcC05hboHi42buvh3dqmlOYXIg
RRcp7tYd8u7pit7iukTw+CwUhn19Q4zcqNPhzxh48M9A0Un14UOgFqNOP2Skc3fS
zVPT2m6VrAj2bSmuI2ee2acmPRWgDzI7vwTrAaqyXJunfrtJdTfbA1M2jQCHBUG9
FrZKSY1q/kQvRA84F6hWdWoaJRduFzhh3Awvn+VUNSRK3O5Ggg7FLvFBGFxMgP6a
mJ0A27u+/Tkou0FPXTByVk03q/2aj3ptsksXa+/tL+klGK38P96H2HvHHDvtnrN5
VlPwMUozuT+cqCv3l9/DEg+ikpLTaBRr3lh3uQZU/zYDeaWu8JqGgpii0JL5g/fp
oNFyWHlelo9AaS0XCFf5+a9jBGXqkgc6XX1dai+nVwKiBOXkVD42nOUcG6JR/dXJ
BoCDARyR1c3PxeYFGjb65WeZ9mVRc0GaXyDic1LCYXBNzYNPFFZPRn5TfR2f30um
WFhsUbgjnDY1nQbtghZbG+IwKg5NGL9qzYj2YtDDhEA07PXASZ0s2m8Ewx0+uMLg
Yko/GW8p5DzZSwvsSnySESmn9qGb5UnV14fswI84Ut+LS3eF1Y2imnPoTSEeHlyv
mu4DYHyhLGq0/boDxUc9NMVgMq13+DcvI4hvvpD2n7lD/F5JjBjw6HGzGMwh7qR3
r7xuXoY7Pg8tN70/fbIfEqrepVPJN6y1SX8RhkwxsiFsVPu1KviluEV1FANSA6nu
EYAEluBamgpdo8xLAHxiYxdl2lMMXFmZ6B/k5arQqUUmpxVTQOsy3jdiuR9cUHZU
1CkdZ9SYnq4ICo0ahVn49f5UGvPjGwRabgmmiW8sFl/3X7UL4hKL5j5YkNVdLrO3
rf6WSan8sRHqvAB6E4MP7PoSzqCgvLbhrQaSBU0XKY6VyIjaxy7DUucq25Idxkr0
YBcwYbWJfRfEgJmh3rMB2zsext31tgdpy3HQjkFr7VheMjO1+baROmhqkzHw8Kd8
37edO4hI2XVjH06oSLj/iomlygfqAq+kDDdKqwewZJbwKpHFDoh1TtxOw/sjb8W2
rqma82xiaPPcabRzKs24l0amP09BYqBNXFx0JGz3kFWhNXaM33Z97T0g7a7GDJa1
aneWoU9xc/+jkB/0eo6ENpw/ueVC/VKmNbG4eA1doL8P1stbSZ66I+WzcchcalRf
Y1gnLr2yr67UslLRx5TQpyRc2Vs6nXi+FBcC0CQrIjF2SsHb6sm6RtOZWuaKj20b
Pk2/ZGf6U2J3oPVSZuAfnC+MQVc6l9WBwUa6sySKFTzlvD65RJmibQl1g7bkUej3
l80nbUkTIFgHAQ/W16B7qbVog/12sP8N+sJowoCsAKtnUGAGlyuZbgFXPntEZWMf
6SykPjKvMk59KmYCXSdR+T9kp4P+Qdb+U2h5pp3b/C9SSERTruVgtyJICGrRNJJY
m2BcKsZOf3Sm7KrM+dRKVlnim8Nnxrm/KeVDyJRkrY4ZF7agQMJQusRFgMEc9UoF
YuL19IRuL4Fel2+J3Dl1kY8Q2PeW69Ff3A3IdtGoy11/32cAExrQwtIR94uGWeRi
fDNxv02aSpxKUZY4uFyiInIua18CuJDPylBwkt6hyy0pOIzHvCRZLTlGL/hQ2Wgp
GhYxKVyQdfn8N5oid0FZxw5XYa+YoHFaP6GkZOBLeJfHzKOGIdWTJXqenV70nqPU
fFB9cmRPZ10I0jd4MvHtxf9Fz8wyKF+2ErQZ+XLagoXCzBI4I0djDnsIauvKuZWQ
4YJfs7sNn4cfadR1QUSRH8p3xxGN/3XFZ+S1EXJokMNaxjkYZJhoy0GGuteeeR+f
+N5RkypaLJ8qnvSI9VzvZzkacxlxhQPc8LZ13zEb8NAiYCibftxChKo29MU2gPOm
dPrrPPkSbtv9vrj59tFtShgKNtE4ZdUeYM1p8R0d61jZBByeE5P8e2KB1/q24z7J
duAxY5yu/zY7JZgXyq0brg9Ai+HTkVfG8TBVCyI/vYsMGwDMpcPIB4Q8ByU2ofIi
Vx3QVF0xiteNYI45SteerYvThOPMahvUF8qi8V1kxyH2TjnBtdsOQ5AT0Ho7h1Nv
a2h5vgBn1MkBnxe2cJRS8U46yJSMcnlPeTCvM2MXxq2yi2OtNFg791Jw5vRbnKpq
VYtrmrwbEZtzdcCiAfzrVMve0hHGaH4gMN9aIwi3ZAlWOV59oTqozU7Hh6M+qTgU
D/wvdTNGtcLpoHFGiheL76san+nyrfJ/nNj5dyCchPRcY2nOqZ+u6TkzV6KRmB2o
Fvm9RuQfY9a1Hz78zrb7HptiMqwULRlyNscwoWaAjg4W7tWCD5q8Vcnjjk0VG04w
KGEzBKDl6sfixROeg9rsc/Niih5zEAZZTQ0hQO1bEzhz+G1ylX2xb3W4qdTJBqsr
9jStXfN73yIviay7ZcB2JGw27EEHoeaMvSmwWh6W+JjpbRhPgjuR2kjM9Ka2WIoE
b3ymkr1OfSPeKWea+DMD6ms8h29QVIy7otdV1YCcW/OCPuUuHsfWv+orWe3N8XB3
v5NWU3nzyKO/LL0vcCGfTZzmzbUGeES8t1O3bSLLrJhlf8wJseLbxQsoGieW/FKX
et0qc8lH9wNIkZZAMz5DT3iIGHtUyJy4+90ctMcGJLrHrnQB8Bi+ppWingRRtY2I
8yslGqVAx4KcaGnv29vgp5xK+MTkAWxVyXYtTMQ/Dt2DYOJOs42zPTN1mVVtxDfD
Asu+82O5pLyM8OxNrDAF83pb/p9i5Kg+Js/+t0UmFH3lgiBIraaPBbeYmmnlBAad
umTURWEXsfjMUwGXWHKPZiTQxeJH9MZMHZY0YNOvluI5pDkhcPJpDYNH/348ks4w
Q+386T9RAHKu5HIZ2pUxwhRlNCnXh+L29V1eCuAPZ0Qtx05SFYglfl158JkQyNE2
/PtLEX+0UPyVVmW4MmrTitZYj6hqGgmzPd2vwHx/HWjsIyiCz6j51HXpw7j+reWY
l5qwmSupzi6xAoU7pIHFJQ5eYap57A64FB0+qv4v/UM6SHsODKGj68mopwVSF+lb
AZ5wm+GJS4iXUUlxnyxjZomvkK/yEz+U581dDFj2/NWdnlpF+/YXyKYPJhlGq8KQ
AG7R6BJOYuoci13k1FSxBIUTg2a/tfBwAR8LTpyWOl47BwrDsboQ2hkVlvsEDJk/
mUoxKs0urzPepsJv9hHsVzj5PPrpW2q0US/geFAMHc2NMfBwHyaHpX6edzFFInDt
igIwPe997grMtFzh6b8zIqDBBf+v9nR6aqi8NXZz5droC6T7JfdPsFSEEcrlUEZv
oodtXlsFewXgdRjrEygHLXEQZnAFZ1PJa1KHgd3zGlMMe5NwnsOtWHNfKQ2dt1Gu
25yE6VkjOApM5yLeiCv5ikZvGh4MNWpYmKTxUOLb0yU/x1S7MtWLZjUW76qxfws5
0q4t6ZQRAVms/GXTV4xiy977qUfFmLBYRu4dNRhOVHnM4bit0TQBxyvPiHjYKr/v
wHxz0gmulC35sylrfCc/vlnf+1RrzmG1EZ0Z7xWlYfZdqPP5ggWpeDw+sOIv7f2/
XVB/zrHb4YCeX17OBiNa+P4P+0g7X3LxQuDpUhuyFpAPPQq2u3yWL4B9Ib1Ckgv5
3c0pAxlaH8HN/zppkpnOy/PdPugo000m/sGylCJo2cB/7bg8Uhr9QUqfHH1nnCri
eAs3Adeafhth58CSNF0DW5QjuxOygEsAZGZy/i+L57qmZtPAmqFv72Nw5TTmRl39
UX/LalHSpm6NdkQFp+3zBIS12Qu1ind5D78ytnm8wTKKJ3AiiMEu2H9/JZ2GhiQA
TSxJeBQhtAWmG9PaO51h10JuM94VM5r0zZF8M9d2v1Ai4EmUiqIZyY7uL2dM7gla
yZN/lHCU7aujmV+AOpRbooz+WLW0YzzBAGe5CCefTrIJLom3g5Z3QIg5deLIsAHW
d4XCWudzqomoDfvB130Kc8NaayIAu5x6uA3+0LTGXRqEOVoJW0Xn7C9dpnXoLdAv
vymUroHtwynv9c/pKmfBOBuOjXXRP6hxJsieOpWcGBBn5XpSmg/RymJNhd0nsXyd
7dQkh3sak0wUQuRKZlMnZvm9P5aUDB1BNUY6cQ5h3t/xK2Hv5ZFl70CLaqDhubRs
9IssiHe1OqxBZfEf+IuZ4GMcJpXiiKCln/M2h604QhCsmeGkkVoSCRyjNZv7vfWM
uhR03mBwX1gRhsq7IXPu325jTQw02ML8Z2HNUbKF/6QKOQ3sxRcfpsRDLFEq8Nxe
2nsMq/3Ggexo1QccXUrh4cUWZgYGfYeYVKbNFd94hW/4H8qELS4M4CzN15jM9C1u
Ig46Zo/iT2Zz209IYCp22az7HRKRMCCnHWjhCFMRgRmfN+djkiqAdZjoErW2PcXe
YqUHLm0rs06FFEDXUHd3KvyUb59aqd2Ozf8n7lK/tZihx2l3nwQPmaj2gUT9jOz/
oEuNAW6EqakXV45lH7fpbGN0PsGzqW2BlfXycMHWPFfEzE7lwWk5I803A9xbQfSV
En3QFwghxAsDXdjBr+RfcxZSUkn3/r04E2HeGRKX5rsvAuRjDtQwtzor+I6G+4pV
pcTLu34tjqZfzY+61jKy35MR6nHn6RDu5nsfgTvl8mP7L9THG84wVlwEBj7zICkM
a32J5wO5HL8VOlA3/4srdOXjIYoO2giqyUal8G3HbpQrAfPz++DD83sf1XgVOz1j
Nex8tMkBJyoqSbn7el2Fq2KOH/MdTJ1vnLZ16zCF0e6qfztF1whgaDUYlW/WJgLw
qsAvtelgM5Dxw/2DgZlVSj5+bWmRX+ar4Kvvmxvq54PhZ9j5dczDY7ge7BPPmUw4
DWiC6XpN+JsuFY/QLVTd0U+FDI1B93Ixy0/o6j4ZZ5GJVGzaxLFAop+R8Gu6nppn
p7arRhms0as5dXUSxP7i77azpzyuLkKssb394N+hd54tUXWGUOOOTS05l8crKzCe
TJY0D07SaBOghbxLvNHgBIJ/asols2w/Cec2mJZEQdzwCid2cZ8YaSxs9C4q8BGV
EROCW2KqTUXsSs4aClsbLBWtSj1Or0+6tAmUitiqzVydCXu4yZclFJm4+jZSYryx
BN/ved+ZW2Ty15wahDhA8fOKM36bqPvuweGZ48QZ59TVk7f0tNZPgxYiAa4qWGXV
9wx1u89yjeJQ3tKyKdyVP0+7cJF6blDPVl7e2dFWgk24NF+jpHLaK9OiIqYYnaE7
o8/ifJZ1p0qT9sPqVWt5lyCWojONRL/ZykRLuWBLcK6mb50h16RJj0XAcfcoE9uj
jbz5yzTXcjBLmQkwIINEUBfF68SDxdRSHMsbojjzKkb7JrTHQtlLAHP7F46Eej0N
tZUrgrmOTPUZAC6/Z2U3ucLVMDQoGQGkvKTyWkeqZ6QGDUla1Au3xhQXvqho/16J
/dH/fMBzh3jkC/0PDn06arn5GD86ejjQC+CnwEPa+f6ukqKoDS+ZqbfiGtn5wDoD
oOZzxvImsZKCgcSbXRYfAibs8Hp9lpX3TS7kaoHtT/tCWRWr+s/rINt5y7l6K5N0
bz1QL9FMUzTF/9u3FFeAuqoKdFRCVJ5HjCZ9o4AC/G+M73N7PdnkjduXr4tC+7JQ
nZbH585Gqp5hTC8+jiKuSsJcj3GPonQ4VZVgs3jSb7O9idriTZ/8F2cisXaS+gQk
NUDGkENLvDpsupiiVV65heUhnKM4AH3ZiByAksMWyBC9rBN0cvFyFnvIwdCA7I3H
RRTKnHkJgr8zL8Cck8jciZTwYktfHSx6hXviICpy2hb1mKPHXUXKgIf7Vx1IYekZ
8TQN53tHZJIF9WJ9JYJ1B3uU47JX1BCPMW767t/bnQA5qk5kCdu+RJfBQqobzNXW
fb/esMohjNOLOR86gd17z4YKYuFfXRVXrzzSJUIw33GPVE05Nh0t9Vk26YlUr+E8
mcm6Uc6U5hCJiDZ4nra/nEkV6ejxkLBcTy1oQetwgoinMnW+N1ur6Fss5SvetDmN
vJRiKE3UxNH/9qRI5tlnZ7dOH3O6xgz9Grj3PrjKoF6XxFUQj+s7Ow50XUrLDHN/
7l7PUty+4n0waqdT7pO2pAn75cU7VkXLi8v2pVuNDAQVj2MBZsBvCFQmoaXxV0iN
leJ9pH0sTCa0xp5ztEoea/JD+tYQqkodMDQ2iwOrhsO/enbNLP8fqmuR4yQIblJU
JFE78T7QOs7+V5HoE+210ZGe2IeGwgNOcap9EVfJuLwjKXXvfZ9VaYqTIGeLRTEf
C1DE+sbf60dwj7Xih15/aOQpSxDTK5zpiRL+aF0a0rfDDE2bdQDsHICVoeId/irJ
zxeZosg/V3Q1F0zrLL7f9uW5v6s4SlDU5yK9Dno+AbeDsWBy38ggPIaeh5goiT4k
i/0k29KS6tF6R95lSw38jK6hlItmJszbhcrGdp4v1hy5stZYRWAehn7m2Jj/jX/X
HgCPg2IpgK5cDR7qBlzQeCHd1+zaeM14JIUma0W2eCSMsSYgwgqo2A0ruU7Y8Nl2
QfRRimklJmNxzpBBVcyAILTB4C1AHpcFjTxz1bi9FH8wRQJ5DiQni4vBdztQu+8n
DZimCeMhvactuKS4W+g/N8+C4a7CLujF0aLqMPW/ewMyy54yffUOSYIkSHFhtKeU
SXJB4SYnR+CFoKfPY3ZVOvndcA4mLjwFLSMY/mcLjd2kBXs3mfGJopFKr7rDLaJu
nnculm9Rz80+dqGOFTWCkEz7Gk35bD3pppPanQitiwYR8SBFBhDo3ef3IrUCgxjG
umuuKoCI6PgGOHn1ikN3weyRkEQvrx/9vk4TISjNF2gRUbNxstvbktMy7JZq4GxH
KQQ6tm/xi/tZs+gKlKyuGfs5qSZdi7VPHHPCPb4KW6nnTr5QSzw80NEq6Ag/o+qR
b1gFrz73pFXFAi3Jf9APPbUaoIY71NlG/KmBoknbk5jxXFx+GLMna4203rJqD/fg
pMUb75RYGt4CYGUVyYDS0yZ7hJvuOa6bMvdfI7CLw48VB3hWZ9eCPJZPKGf1Jtp5
e09wZgC9EC3xO5irkcztaEngfpd9Utw4DITkwOcVzhjoK/ZMiFo1AqQlMeCcPgbq
A1LAJ5N1VSpw+En7XHpvBTkE3zXdmjl0ZF5Rc0GEIm7P6H/ejLjzHARSmD4nmmDw
9FulqrVR2DbuY0BfzKcanxmo4GR+vVfojXABsst4AqNir6ujDw4WAJaW3kJdXj3f
x22kXT6NhLL84EIDGvR7fUulFfwTDiOqK5PRB5zIpU/ih5ifVv5TpQRkq1ZCl1Ij
LAkJhOO6iOSIfOtw3lUhfVzbdFgvVyJVKiOfbFgDHtYOYHbXlbnOrb0BcCHyGCYy
K/6F8SSfRImAqajkjx0DQ8Ocxn49QiulTxKZQnm15E0dp5YrtHiKGZLV0G4Vb95C
JfmnCjsUHmtJG/gbCEBPs5xmNME4ztyeZtojiJrBd23hvZqD7q6d1Y0g4rhqHxWm
kq/CkAJh0rm3iIepjygr3M3Q3w5+sAX6uD+ycz/LDiDrCxNxk2Xb6C7lRANHlDUy
Nz3XE/IfsWKTYnow+rzkVvXweR6zsbiIo1YvB6YuZhFckzYOGlaBLoh5QS3+TLEn
RMTy42iE9U4bYtQKWAJS1bE24WyZo4XirDqPPz1wTD3hbXVyvBbUPkpUYW0z5Xui
8oqR3lhxEW+HYYkXdNY1qGqPjwJkv9sDBHc/uF0qjXgDj4j1g9BdwZqnH0pBMYfu
dyfFPwanE06Rpf0HLD4QsajNmkktZ/e+47lRzseYdmtDQY3jYRjx1cHqGiLW3rz1
DuT4RlhH/Aod7kyuPRPk/RKj+TIMBYs2p6Qre9YQX6HI1RnZoZZVHsb3Oc/caKxw
Z+E4HF4gnO2pbvFvC2wIW360lIO3Icordq1lhBI5j/51BnflwxCo6EkK1i9wjXNk
RuLLk9JHr/0Vxc9HzM9/9XVUIlDE/5CQIFMs70mo2NHU7uoTYCNqhyZP7av7tO10
0xWzTq6YTtsniJ6dnyIN9P+iPgcdULQw7qtbkFcFwohejHNwPHfV+OP2IOIXgiyk
O8YEPcqbVmVfpp3uDTNMHZV3bGm0apmJC3QEvS8jb8AZGC/Kic3h4d0kUfZ9pvYD
3EwvTLAiUCHpbWFiYTufXf77AFwRY0MMp7Ulv91XC+K2BBIBcuoEvcNnAwcKFSua
rEHlw0wKdF8F2/qZyxXVyv3ZsyWcylki5yRrjzueS9bzEimNLmIdmlNDI7zQ5m/C
sWvci6QZXkvrZSyliQSfdiRxfOZnUPZZt1g4r1MizQtRGhxzxVJ0R7FmYZi1FDoj
MRPpJGN5BFUcNL1eCiFszQzdw7FbRU5dauv+g0oAeOEvCUeXtceMY/zz7GNpV93R
WXMCQJL4bb/doXLaccVfVJPjUSAnGdyPsclEhQPkgMQHBLXi17CQBkMERVp+2okp
lroeo1aUZ68KnM0+OZH57K4YAuJ5Tvf05wI3fsxLS3Q5booJUR3EMZ5Bev6FRlRP
Kgk6L1BGYCEi2RtWXS5mpJ1t5TuwfbNy/HdkoZRNduSJy6OW1HHWM8+LscsaVHbZ
m8DE9kp04kggBQAN5l1umANpO9CDNr1+LKLIZoofKgT5PguNEqtgyaqvHy203zH3
HIdQpI/3URimhwdSCg2dBtDlTgZ4Z09GjvLK+psFqq9PzN2s7/TjzZlcHEt3eE+i
ACS42jtAbB14s/a5oxCSEYldo/HRa+vGdWXoaMOP6u3gCRZ46RF79iny9TTygDk3
S2ir5sQP9MNH9atTGL0Hg+jVwonxsE/YdlwKNwqhmkd4pHC+mtjRO+I3ewvxTVNu
ta5vLn2gIuO6UEnmTi5sSU4u0WEj63W8KtwatAOxcm8zk6S8DudoHjjhdwIqPx45
o+63vY9qz+ehlhw1JFaoypyshB98r4JP1zr+gExsZETk516rB8Sfxa9JxXAXYrUM
AGSQC6hN8v8OwmGcp0YoN7tBvq7LPnrI9y5sQ/CDrV0Km8WFVubHlYO98xhKp4aY
56Ux4r8m0fyn21aArkM8xCMtBqeZ2h7SUAAuo6vuoEDPyy96FSuAdFb9QqJfJ8kK
FD7BP9gOAKuaXG4nkXuAOa+9Bnx8eWyG8DHx1ZbCx3tZyJ3nB1aYKfJDzDyZP83m
QmRU1qm0eFSVTkiloQSPQk1sWjRewF71b0ogzzYRmxVID/jNdijJiBwzWOYGcnXt
IxTCltS19qWxjUHGQPbUdSsqons8xQS0i8M6u0ff3q5ajr2LZcsSL1cjEWfusORc
9nKnTjiRf+NJKmAc0WuNJBcmeBMS2HMrYzoWUK2Ix0DIIYy+pl7HVbyqaCiGNGP2
XFLTQAd8phimESEgBJHvXqPJviItzkps8kWP2NSD32KKsRWiAr0duM8tmPfdHcxB
bWubWn9JvCxDovqGoqLny+Wzfitn0gWoPMwjRgCF4IFyyEHElSNnksXJuvX7wEz2
uM5pOIFR6EUbWRk7vnmiP2XZ0Zr+TUa7lgvrq1RzQ0WdI/a398jXyZnY3XN3lj3z
jVKai1gpmS9cnHrJ/ao/IrJ6IKgXdAS7j39iKdDyACLQaLP0uaIpbetz6jzVM5gA
VYeDrM909Z0cJwXKEkWsYnrxf1o9akSRShgskaxxT6/Vq9F+RQpWsApN7BP7SWIc
5VYDGrV23vfJCF1xudGneQEqoVL5vo/YiDpEH/1B3SdhZfR/Ow88abp5HJb6eZJk
lUgVuojggVEsnjqPT9WOiD29+6/BiYbj0u1YcXeN7kTCUZ7ncLPkgGjSovT+CZgo
p8V3WwBhNXGu7jw+wrdzqz2FDHV5/NYX/+kBFoZ68c21ca5OSXQdfR5GClOmbgW1
x4/BnaxM0Rqx9fG1GFJoVbwK3+OrY2qufBBxLhfpZZyJ11yVz9DHZyIrtUTLCk32
fMLJwcvd2EnDl2ykRHSoRLMlnHEd0KP0WNLUkMx4/3HBFovwoMcIt+oxcc7yDE0d
m+AqL6tiFyNlq3ORFxGJ5T5ue2zEICf/fDb+M4wRCMRgkX0f4IOiXY60kccmD+2s
YqDAE7QKWVr0KRXlbDNM1mQSOKfgxTqfcVVq8NS4XL2M8sKCdcrRIc5d4PRULj6/
NahgIM/IYbB6rX15VCyZMbLr9DRojk9TTHZUnsNdfDtvrWNQDTfrwocTql+FSFb8
DpbTYSQ8xqCAgP9Ph1rz/8LDrNMnuLdrMNdkiuXIoJzRSYszHBLzWJwRk6VpV5bK
bP5wzcCF0TTvW4OUykh70fne5BERxJfOvc1ASFZZqp6FCAJCVjdWAE7742Do/wRz
RWIRQyO3S1R3TYaYERHzWO7dcFZIa1Zk/795rm7BTJz7xXSqGLfitzfSFQ8j3knv
+O230tv5XTNL0bLEgXBelbd+f5AIGzYuo4HmJaA6Hawke8UdE7PJ8TiAVkeuEr1Y
KQ1pcEFhOh7feOuVsUF3OqsDr7G82cayRwsL6+IEYzrJq5XMxZsQIdDMr9k7EWiv
g+b4gM8oPdRLrNz+4yPxQ/cpDk5ozzUGcByH2H0wYzuTgXf2+PgcwsrYHz32bJhT
gZxu1gejTKO/rB7ICYpGSWxXTGK6qnrh2NKzFynQLDXUv2T69gkL+ASKaAeq/e3V
NcTmEkb7Xba4PP4lBqNaO/2iBBh8r9G0z6RfJzS7PjFA/mwA486ce/GBX/i6wAgd
hz53wUt9Tt9MKs0i+ttlwfveQEIF60o/AWw6ibN8MvtbH+iGaAF9uGKkvGx+QOiX
xE7RTPe5homdwRg7UJPNHVNvRQ7NxqzvjqORfnvhKr8hHN3LSNtiCmQNQ+9u9j8m
DmTY2CZMd9H+t0IXCoqfABeAqN128hc3ggYEP7dh0MymETk73Zw3un25TwTQXcfX
xw7v40JGfp7hzLxNk97oyV/0sF+ED4H/M496C/9ig2VdYjoDV94CPgnaOtFIdUvj
5QJMD9Of+oCDVAvOwDZcPNN31cQA2UxgTsTFp3MpOgG32Qy1EqO3Ql8pU71g2Sin
DHqoBijvxnlzmzQE/IEBmDU7Nk1C5uYGfqW9QuZMHhYgfpmgEPCJOmEZ3sSsLxeB
8TXOBLYWwlgSVxacVtV+xHYkW2jU7lc7Y5A57i6Re3z4dIzEs9ko6s089gjNl7TV
CKNw+AwLWxuwXVFWqU5c3l6spbXkqMpwu7fFFHq/DW33CESqJevNTB93/0mXT/HM
NP7xNdraqnsMBZH7AZfk4sMWCqw++QpYEDM4jbMZGpm307xnpGhxoFeRv6aHn7DD
dN/p4wyoFBx38KWcPMWoYPqE7eJOa0wwDSQKwzSv1F/12t+sZLSbOoh1i7+D3P1/
zwUXCf5Gf08MsayQgortQC+I4k0V3h65I4Z+7opGFEoLBsUnKNNXK+fzv6XGpT8s
msLzOdmz8+Af355XmGROSG0rCzu42zWYe4yxvKCvDtknP7sBk2m5h5nHYk5uvJ7p
KNXzHoZXaD+LMKazw6LaVRBkmcr3TowGiYOcjKNNcKNQ75S1wmFeooEQ/3uIvybR
HufPeGnXtOdRu3h35kKr21rsdCK9Pmgg4HviHdxYFwVwE4ScQulUYdzn/6dZNb49
ML33C4NlRJCXE/IGMVHxAwm2FYPRDNweE8EU1qwUoMup3r+OKpQNILJVYQsS4+yt
5NoMMBp8bCjMHzEZ3HU6NlyOaYQgR+SG45fUozKoczm8jhZTcBNiv7VkfHO7TPyR
uAynYHZ4P3ILv7J4gVSasjOCQW3uw40b3DIt4sw9PXuGET296DJEAk8qvRVKVItt
IsTNWUQWDVhmU7bHFbQkHF2Yp+sfjCuy6z71dPlZ6I7bchameOS4uDv4cQ02KZZp
u9IyMCFseB3rysPhdwhei2f8QRi8Bgp13Uq1TORpA6hpQZF7NpTsE7n1O1ijIdEV
4WazDJvHGA183z2YZ3kKalqU1KwAS94uHaDMTjmhbov3Q9kO10uSsNjjp4mfoOsu
u0SReuos4oUR7qt+X3HvlZd/lZ1LGuHu93luYJ7rT8rVOJpm4NNpLbdRLwdC5yCE
18TEUKZGj7SnlALpGmbKNl2Pq63rMqLVkd7DMrjNu+5t4TXCRy3NhHSer+MTPwYo
VPD4c3lMkBzFlBgr7z/1Z5poLuoQaGdvainnXlG7pvTy0Qo9wSX77t9rWCD8mg+g
87wtpERpVd2iVI3Tk8CYG3HgBc8JZdD2We0YTKGYqXBE17g2UQU19bPomAW1TWYj
OYtDRXZyozYpmq4JR4I2wqmV+6MI6vYXseN31IbIVu/o2uL6o9jzj7TeYtsjMujQ
jXRcSIzC/g3VQrbxlH7OyBlsg38fN9PizJQitOqlQy+Y7pUbI38WWZhXHd2RrxvD
tlk6qOftzXKD2z+rnTsr3mHV7/BmcjY4ERRtwOIpJP8Gg0EhKiwFxl6jqmVAWYuY
skngN9elRpG3eVOifH3dagUFcJTXcSNC8aetYjVviXAe1XETn4gdwP1aX/2qn1Ps
N8ZfiJm7O9jVCMX0aeZvkhBw6on0u4RCwozJixflASPxzVBugkPh+3Qk+eitH1hv
BnIuQfahezu7F/3y+ZXdIBKBnKjpMijFUgUgJLL08f+PudbtWozCUZWmwu6j9df6
U8onxjHeS7MV1acm9gFFMCwPUzoQTGyofnbwE+ppr18OEjo1cheN6t0VyH/x0I0d
Am0aGiyItdYttahS4ZtrXQID8Md94+At79lhb+O6qBDJo1AWg7JIES1GvGDjXw/9
J3VnBKxLWz86WCGqDURNOw+vuG856LqfgODtwpWuytQoP262XhbvC9PgzcTlFEKG
C2XIUZP2O2JJrzCXk9mJjIaQaNrBS1MWNX4tGU71AVKKrDD6LI/9+76tXKioMvNv
oRKR6IojRjqGWeaneSnTKaYauiLVdevItcCRjvqbFijTZVLaMlooxDtgN51xrSrF
1usJAxbZbiQs4+NG/vWOPWMQD80YJd3mxUtl5oB1jgQH6ZGTmKfq9IM04JJRpsdX
Ruu3/85sjBNhsPhy6RM733pwE2DwLteTF5l2+RL2gMETEb2utLzbTP+MQoTP5Fij
1TE0aKkI61OTrWWee9mV/MkkRm5Rsh6eg0BmmOj2FI00vjd+1Qn0vuz/0SMSgMZL
TvaqAp7KpVc/QJzfqmrgXhcpTjFem7ONvOFfcYazedTrvjqE0A6NwAElkTnYqkuE
0gGao3glxGh9cbTtZ5eN0EN6FyC0GJnA6+EaMg1ylmnhps72iDIWUgCgVufaq1Kx
EFe/iqqEyMoN+oAiu0D6JA19KGViFGDzvuWL7pbfyq/IzUtD0MquZltkesbRskCu
43xl1n+ij3RkqKwiLE4sFxNAo6dZlNFfn9ZEdOXgeOOAuEevOYD+gmF2PLw/LV5j
m0adTF9R2ck4FTS8R3M+ke5XEpHDbR8Yso4xyGPaDuGnL4OgFUH53YwqanP4Phdk
YcDUvwa0fxGqq7J5ADHDbTfqoZ8uBw2xakkYafuQsNu7I6RWkAo4tchZFE8S2ejr
NtZ3zIsM2OzHJ/O/3m4n4L4Tho1ppb2Qpnsvp4MlYwS3RVUsVm/22wFcC4VlMT6L
QHHljS42YlU8x2rT/C8MDtn9v2WH9UorEMCsk2L+LpQx/QwFR3TBrNQth4lYyKR+
umu8Guubel8JxwgelrsnL8JbBfuvkxkSdiF1k2sKXDkJl3ZNr/QGh4f7r+1AqSFK
N0WnfyY2H9umjFaDnlr4NzkhJC36+S3cVb6GeP13rNUaEuCnWs+WdauCYv0qa4pG
GtH7nk0GpY7r7fKnIrQeRlax4rwWp81ZPOJfqB3/TQkJf480fI/Z3fBn+e+NkGgH
zjQW9Y0BrBfcIrvLwdLo7NdRdlO6a+dNz9S7BptKklvqs4kgryjSTJpGE0RHNypn
h/O0NApRP8crR8DPMY/BUBs0T1Cf0nSuFzqtvbGl8/6UB4sQcJjEAOgOsbklDTuY
aalXNyWC+Y5bl9cQ4+dZnK1cLqEWgEa6ngmQNNGWrgaB1tZzK+6U5ykaD8knv+1k
I92sHGfECJxNdD0MTgzwKdpUBW1GJnQYLPDECyErMvWiYW7z17LbL0ddQRvR/wHy
CAMsHn9114NeqDpRBIXimrLCZn4ltL7u1aO8Lnx6pYw4zORJGvlEkBONBsaRpx4C
gKo3ElYKxBUtOtOpnfzsLOyNiNTDKrtK4pJBEMBNLes9L350BPVZw/vaFI+2b8lA
tgwP9Eqldv7s0C04NoyIfY2t0bNe/IGwPlwZnU+SjsuOx6Wyi0zWhNjVG9qwKiJ6
1hd9oE0r7YT0gjf440H48D4pjZQelNPpHFO0eBfVYgv8inzyX/0N8YKe+KaQsQkq
fRNrGBnXGfY4EGPFkxO9/UWQWLf/MxHtrcHV/H3ExASpSrbNkL8U5ldvmbjPy5Pc
TsCEBQbGsQVSfMvkcQvvriX1xhP3P1rXoW7Jk8Z4wgAuXPXMXMnHxZIqZv0IfzyS
+yjsA02UgqsUUkgxoUTq6jXnEKBEYtYoVTv3fh/SGA/hcl+Q7j+noJx4PCBFK4xP
pH2r4++Gl2mqlHBOniaE0Mvt8W/VdjOtwmvVUD9VP5TZGchb5rWfQ7EthpuvlKwV
bwByF3xBBJ6DkhQ1LK//txEqz3k1asrN1Tx1PuVVZ6WbhN+Nym62Wtpdm9itRdfM
VNVeL7oKQF+BwIwL90SaD6IsBoiA8wMep18u0YzHGcA9BRuDWAQgfAqj0nX6A+J5
Ne1OJzlPwITSOauA8F5gC1LgAUKG9/vwlRNstYUW1P9qv6QOuTFssm6MiLf3Uzsq
6Qkrq1vEoHWhhvBq2dSa4/CXYUzY7x/QeKQRhVDjHE6Rn3g1WydbWGalYHVQj3KE
/BfJ8WSsmp7x6UTtOpxxUEcoiy8qjCS8Lrc8VN664fVAz7dMWZ6E2JRFZ6ypsbmH
sUkGqVmoZHpRNU8mFe1WQ5Bsb4g4y9p7vCKMGwB3eRUuurKFqdEtTUKGlL9SUBNz
j7/tKp+UWVpwy16QGycUkDF9mYRsIgRVP47iywW6FDmSjWFNG+IFfIASv1IiDnaE
Y9njKJxuWvGgY+l8FrVmvjClbN59Y7/we2COqQ3mXpsmNxtpa2gtOi+I+FNNoBeE
+K1duC79sq4/q6CoZfu1lPAx5YuxMkhQs1Wcg3MZ0D0TCAswh9V3G5q0z9hSuPRd
OHC7O8J3D/5T/Q4vbOjIeAuGMeYyB/J0yCW3LNrR8UTf/QDE0lWMrecVkLqbhgW7
HWc7kHxfTamONHqEYZRDEkYzWO3XWYyKfSDd3ZcKryJT/0IIcM8VRoKIJo8On8y7
pKCLZJFpa/cu2sP+3mVLN7IYE5bUr9s9dQWrzLsbuFW6O/OxUiEYzA57bIO+YW20
mgMSqVWMjXNmqNCoWw8kFP1qFJq3rIecAtZH7pXlxrNdR4so3ZHQMuo313APG3J9
Af5iUAO0cIYssQATa5q8C8wz81qX0PL+R21z9D/n4Rpd7T3EwFisI7jeB1kXsLZ0
x3YeAbgmjzn/y6wh3BiAkS7Fw2YJBoDUQcX92phlY0+Tak+hbRElnezmFJg4/Pib
N71YEqNhdGkLzyptU9p++BLele3BY60LSKjT9Pd5GbtlxZrzKPJTAQyO3ohNMixi
ySahcOL5sKTLGV25iEND6Gob2loVF2AJdrakI54ZEPIH6w7Tl9JOVUSI0IBmjLAN
/BnyRcWI+m/XfATlqPbqcjDlzjCVuGQxcGgMsevFPZZasFPVqMABGn7g6QFV2qHF
0L6nVhGBIfGX7KlYDBN0U7idJk2TiaXQbncLg5x7uaFG+g09Ts8cYjBOfSKJmM3m
33MkLh1/Hdwz9MfPWFKGBLdz2o278JOpIhXXf8WhuNrjekIYvDXgk5HblgRUbRLS
OYlNKsJ7j84tk0UvJXONCSl5kawPuQ/9tqnHwyiV+y5zJlIbsK4bcujLMeQpfi3Z
slN6aAwU5LrJFb2pDte7CqkqlWscyUQCHo1rPZTNFN5qkVej/fiyPqbrcONfFfga
pJDfhFCC0t44gkLLSUHQMRZRW2w0Pp/NRKtdVK5yo3vfYTReD8GOuRIp0jbAGNTR
14alYPLJud2kqTmozJpq3aYSx7BCDi/vTLVe7yI7V8PcajjGK+M6sjBZN5on+PJy
tKC953wb0cS3dSMGqWSaZtINY+FOyph21YsTub4lzw+dkezOX830UTgB4clGUJtN
Qt9ws2oNK6c1d32XCwoTi+LAPI9PJptzR2nUd/s4gsXk5ovh2izacwm0cqyPRdyc
6SNUi9DF9PXnBxMYKoYy/TcGpqTXA4oozuDTfDSYy54wzWKdFPc8piVhE+Juwywq
xEDbSnlTcrw2EbqnfElLy6k1RldxbVszh27uKFeU0UIw0SAQXYOGRuf3pm8mYmbn
f/X5bSROH4gHGZ2se8Ticiv20pxS2Cvaz06SSsw3AjBog6bM0FymO2BcCXK01LGX
+OOBxDiIHDtIDBaUwUJcVM14UiWygcpujegREobP9Iv6TBOe2gX2ny0plY/E+dKf
Zz9Ij5563JHV18ffC4EiqIvbd2lWqZEClZhVp7jVcdA0oAkRss/XUZWucXC7BUAm
vdy860W02y/cxG8c6ZH1AfCHm+FejXZH8wvfJ5yKQlqISyw/zfdi9LEEIFquAIgW
yVgqWE6Hi7EpQXqVfL/HLjED9PAh2Ca6ICvB6T1ZwstQDr19ba5dkMlWiZkGyi5r
2ae19hiD0hea4Cug7/aq4kbG3SC7nOvMLWkdSV+8kz1gcBz7nFsBDDwexxYot+aE
GPINbhmArQbDRUhRPlI7aorisbicDO8QyY8jq34KcGlzC9rZJxe7PRHQflUP2LzG
xO5ME4FlanfuloN1c41AXkcIhW6XE/lRpx6hckuuMdHBeppsAsfU5AOOw7sN82CZ
c41hmctSFmcMC0pToviUUPoRdn1EU8Gjj3RYFUB2BQ1cFQJqNYiPi2XTGTUvic/+
IfbI2FKUuFNzE2sMisfDKZGbCfBnI5+mtudxJgozrG5dBiHewIpeW5GixCKsUW2a
Pcv+H3uxUiPsq2IoVGbaMa6LX1TS7G1Kcl2rQguz2gNzMiWYYizOMOf4krniUBcn
+rYaF8x5nJue1B1fRZRJj+rnn5wSUY4OIXTDufiHvbl8TeCzRw9CSujrpDD0nCAp
cl4Dy4WueeO4pdedWV6LdFifwBGrK5dF1nYCydYt1v1TzYwMm9HE/RDtJx3amPUr
0eDLbDAsx+KoGinjNHv9ArbtZ+bO8et1GFxQyXWMoyhT90/cOqi+3oWG6HRzAfSu
OCA8kJuxbLo/+J+i4dktkc+QffKRL52XXqApFIwqjucmhoqHaQMJmyKGM9SGW36o
oWsc7C+9jvlp1fWF5KCh6NMuJQco7xqiRd23iuy7b5TbOTn6K1E8tGFh/8V5OG5x
cer1frj3fVhw4FWBF0hHiN2U58cXMxxSIHj1j6HOMyaS5JjuA13Ts1GYPCcv21wv
hu4ZTkeBNiF1cs3nURlbplajaVmOeM1ZInbsv8niDhB3r2ere2xwHRQKyycFOvlx
SJ3eGIJRNzCFnYIYkdZKOigAoQmOZK5QHkF8iBc0TvBoYc7bLqkAW+GQdjR6nLr7
g0+5gjmXeECGPSkhzlsI56UjxDB9geXDOucA0d3yczmCD2dXwGAPwuprLObzIuBP
i2UMYnYmHMUP3EFIZRH37DIHkdyySiAEVke8vshTakktCdJ7uTPl8I9gnQHGL5Ov
pGFM3Y/cFoYg4pCXnq7x3JSSPlUnKLf1h7/vx+0py9j7ZmAyKqizyNrbAoMkpFCm
3PUx+6IJOAlByKH3D1tuhhp70GUqvThav0u5Mf0Ec/lNNHsPdQzPVV+fTUkole/O
9npHBKeNuugjXuzXS7ZNLNc5RoHK5XZuzL/5foneqkityL6gILLIWUavNdH5YWkD
+IVQYKb6jTNv7fPbKDAI8Jkn3loFC2ZPKNkvK8T1W3u05xlWqg241uvr4BsjK55h
0Hv2dyTwIGBemXQdatnVlibMPKApqyLqFsVRSMbaFNreaPFQCWOORfYiOdHMzBgu
RHkF1AlBWN/GUOCWi1MruhOM8xaYNfn68mzQQqlKdtxwyKKl9Z5MAT8sBNrzqate
vhL7MjkCxoUWW074RIvXlskfOIEqE7w74H9qHt9tqAhCMm2K3MOhE2qtQtXNEYGf
1dc1wlqFcw0ri9zSuBxAYuUEzmD0nJb0x8BcEt4nocB41EtA4J8v7jJR0AnU3fbw
jsL+tLFwJBTCn7NVLRJ//82OV1jnPBJMDCA9TC4Q6AGQYwMSepefFsEGKrJRmiDP
oX0k+ahmqazdv11ayisPceEKMdPFbbc5koeEHkt1O1DU+aNw50dSa5rqboS8B3Uj
qlUszUtS52JDiM4CPD9Iov2JabsQB+BiUiDQ0XWG2uVN3AjZc8aLB0rCRJXFhrDR
8BEnxSx/qHku7kSyrNn3G14AFosuvdmx0Bg5dpIp4uVI0ToE3YVOOkdzs6UUS4Rz
lWmvrL8ZHQ0uofzXl6eKJReTQ4jGaNmLoUMQlIxOhrP0JpNuJgwKSUovraHsq+U2
y9hGKNwn8K6ScqvLHTBlQAsZAczVpAeCo3/D+lxk15hVIIRrkrwgyUf3V/EwVD1s
xlDBMLiJLokItflyqPOKbT3BFMEzQrbj+SEOOzy1tOeoRsqNYLCqHVmB5gfVbASb
WmW5IFDD7WKYNXKCb6iJoxDYPjmbksR6ZigQ4j8s3Qby4Nh30RgWyDojyjRmxq5q
jI06gpeXjAo4OH9kzAsrlzdLeHZEvTnwoKsyt0Cu4Zv24eAbML5u7xIQyE6syqLY
bfiVUo+QK6Ti807gJX7T0YVk4xZ6GOT+EbrVToLzozR+Ci7aKCJn4Mf1UfWYGfwk
vYeAx4/heuYGfVrbBppprPQ9sRynCnxR91AD7EO1tFa+a2GA3qCotMuAo1XUk0rP
ks5QEJDKbZ34k0EvSBK3Mn/lmAElNwy47iIwpDdvEcYu7PP5/EHRlPRWNZKiWINU
MYx6DjnKr7hRQ5rZTDIiEDD7nmy/ccaz9E3/vbnFSElI76t6z2u3YKs2sHKq/73l
Wq7QXXzWnIN+wsrNaoe7GnariqbkdYasvnDNtGuEar8jelZXrmtdMmvNnhm2gpaz
tEBgifqms7ZrwHqPvWOQodib/nmI0o95sVajUUk5abojuHqCH0w2XEw1shjZSOas
Nft2/nq2BWnCGbXlPndRez3HisbcAa0Wba24pSt40TtmvGnwVzG6zmZWN9PeMT20
WVLsCoWL3MP95tO1bVnP5JPYQIbqo+4/s2F6XBczy8Mgl25YVaoojtQZbjd1z9q2
ap+KJucxDd630ZIMZ9eBIwh189KkVhiRMVqEMMffLy3lEdN2XvyyzvCjtf+FsNeH
M+dlHnlKhoe7RjJjFO8fygTle9VTx4rBBigk/kpDsnfIIlDuuXeQFCC1XzXWYngH
qZWmOOhpw36L6fYxNlaA6wYhNVMuOouaocllkGkStMB5M8QbW1p7ujqb7etOVXb1
jmky7N4nXe/3z2juFV1Ec6Lxk/ObrVLWKdLx1CBbrAIiASsouErD3k7rWJeKGHfd
hOktMCk+fpEYGw9V/XHryljTrYwbH/Upyn4sAbsIJkTvzlhP3kGsmirjZzgRoDas
kZZJrzAJF0pSwR0NbYu8e6szv+EmJJi1pqHzWbYrQY/WPhegKziXpeE97PLli7pi
BKrN4Jy/P5frJkVKUC8X0aXLfRGNTsV0ybYhE7hXMputLw5j7UyZE8Ti/TAhFWIO
CTkm5Of5Fnlj5X0I/EiF5WReI8lsNAeISzbwxfydmKyWM1pkFcErf3tyQlUdwTXw
t01+D7aiGr4CNlMfDZOsAUzrzcA2cJLET37sG3rDfd82OCIfKWDjcayJiddhSSSx
++KKgLQmuylEvgWldQ086XARLe+hOjECudnjZSkMpTvLEZQajEXcpz+xeN/mVGJu
RIZAYYw8AoVBNuFznIcyvbDZzqj1aBiLF4gI1bMbo2X8P33cSo+SbEcZUmIqLRj7
6XFZP5/NjBC2aeKen77Yx79gAz/rCldSmsnoPjFFeRxoKa8GW9bLo67tmHm6gboi
M6XiKXyAPTvWafN0kc/QPW9urjrKvDlBLqnFAtyMVTKbI+ebgRV+12uSHlslf1WQ
bVcfEOM7WGbP4YW/8lVtFf1zEBh2CTJkzRfJu2clkaMgEE1WhEGmuXKmPb0ai2AT
sLaBBcj0kKDxvfh6UmrUKuNvr4yF0ko6cxEHEj938/+SHqYOFeqeEMmfvvkrfit0
EhY7/qENIHAKLUcqy60R8F08cY7dTL0f2c84zdY8V8Uq+DUvC70Fk2f0/yOAelvY
VggDuvnd+JYNaT7pI7jYfxip783KcyRnFmz4gT0jtli4INQp1eFsZ+YHI096ezAI
TmIy5e7fYtPfPo0JvECzIVgZkmXPbet1FRxR/pZhEPR1QlzSdNwkTGrZMx+VHKqN
L1BfFfltuibc6WRkH7yPxqU9p9WAldJ5WZtn+MHnVZLOUqtJFb4cOIrdzoO/msVm
iysOVk3e1I7E3phkXZxgP2MSgSsftabVLvmfQ809LSw03RbetHBr/hQrsJWkT2xl
b110x2XRsKkymX1bBxtdiriuU2oaQXngc7fRAWUCytk1eB+sLCZ+X+Uf1WAWjLxw
33FAAQOmuFU0or/CByqbWKtRA+Mz7NNmoCxja3h8XNldBrsKrt7EAcVRxrhW5gOM
Iinw4Fu3ASR3mGUcyN6LdftzYjpiP1P8S5O+bT6Rwus3EuWRADR2alNA9mgZxpQP
z/VeTjgBzAcLSUY9HjJUl4y9niv1wYBUKJs6xIEVK96WeghxobGEEOxgwBK3kS29
K6j5I4s5ZG4yPN87L9ZxJjATLZON06+b22TzL0Iyaxhy6XCsAeqwgAjtUudxHvO/
jJx9FDTzPssgRdb9DWtq12+Xb911ccELsnTB6c2wbu643gCy2V3BsiEiEb+ES3Ho
HV4wv2huCuiiiA3AIJK5XZYWIoZzPY296hyS4iXvYYBapeg/9gUYY9PdwTHbIPtF
0k2sRlAyGNEPTUp5tX29oRIyCQaUqnzHoUSR/LuW7syWpgrNucMBDaj0+BR/2LEA
y74d4a1MAZMQ4y4QV/Qa8wJSTQJVBfmJUIVusyAzYR9jaWUEc6ZmFKpasL5qcTG9
AZvDurR8HVEPcJXx/hLE3EqTta3vebFVKY8Ex6MV/YR+E52y6DzSm09cdKzjdSu5
pNnn6bH3SPMeXzltBTNjXksKi9sQ7+YBn7u5pplKut7rLIX1Gey+NeQa4zC7u7Ah
y8PcD48sDfEGVYowTCb6g171u9gZ8Y2b77+XinigPrbGvjZ4Vin+hi6q313+v/8X
Zac+TTGu2EAxLVZP4g4rPYXkf4EVlZjMeCgcn15UtCFQOgp/muykUBG52NjVWXIA
2IS1k5+CphtMC/lE661jz1wk0RiFof8Ei6Vo3Tmm5kDCSZwX+vDDSu1WKJaCbCv7
juP+5ILFLLdxERyFw7bktbBE/exowhjOBVpoC9hpdTiu/eRlySy9Iv4GINYBK0G4
6tape8EQjCmAcVDPuL9GIB43j9iSI1EWMbLND/ifAfAS+32LQWnryGarmx5Jzugv
gnk4jdWI9HEcCUIQy7cVSUT9M1BxUPqjddMye2UbkGFELT/gsNFODxhNSH4OjgiF
TS4pzumRl8ffrgDCyTmXqLMrfyJW2mVQhO2HU0i6aaYEb/5zv/6WOaIs2P5obFRX
Ny6PUu1q38CNclNIartNOi+JSZ2O0zSagAQl4fl7kJOajVqjH8tPj/gtn2e4ZYNe
cwFuPikpRm7lJgaQtSmV/oTVSeoATbCluHwdrSFVWreUeuWj4/xQtNINd8qMuXr8
AC33KYmt7zdUBCHlAX5PzoLDZsPjBcDjVTZFv5Qbfv9Y8rX62uvTpX6EzuwpSkM6
fyRwskYXyrBXp7e/HeJx8YPdDw5J/J5tDgM0WAvW3jlE1oXCj8mOwEoozWnU+A4g
aSK04Gwz0ZkbESy+VjtidIyoZEEySD14OfWs7b/QG4RXskHylg7qadpp1p8Arb6y
s8X8CJlNOc017jFVwEi0aNHyeBI8UtDxWMWDiZHz0EZhjeXpJHLWjSmZKsTfJ+rV
C51wd7tv7rmp/+6ac8iu09DfpdZpBbzoeamrLDQWgIW08I2r6fTRZEr45ouY9gRS
whYI5bh8+H6+eBvmwB0h4FLtH5njiAC8HJ4JMHAGit8eBPhI805TmGGvAHqEhHYU
mEI8TqzJKJWuF/IIQsOV5+VK7xE9RLmu5y3dJ+yGws4wJmJe3QdyKuCACoGZ9Z4X
/93tr1dPEFbXouICNWr8q0uccQL/l/xraOVq1mTF03sVDBINB0evQLe/C1wXyOa5
t9G+bbPb2Qmci3nURkZRAbZTmw6i7qTLZklmxsGAL1Zx4RclrqU6Qt4/ZokjVz/8
CkMdLf+QI48sm28qObKYbLKbUo/yTqT+VzBUU5DY1QiHcsL3abQhBjARZPUE6fyA
BvislQuSHwC6rSRpoBBvYyNOPPqtEUQSi8rwkKcMOiRatOOT+a1N3Y+clKSQggNh
ez7Ud+xfFQaNe5qBIe4JsMMtSTFVObhB8eaHlM1sgTg4u+0PpexKtQfZk4UPPeXD
hF1h7gBfG6dXjC4GSJueQXOLDVXGAJ+s0SXHjQcgeBoIiRPmpQwIP6EJGPT2MrRF
HI4ENE+To3v08L0ROH4UUk3Q8nAyZNRvt4X/nGZ3qfu0HTR69M+TU28HYp0K1wio
M5Bup7oSyW64c36XCPhBtUTUETHg12mI5bh9KO1ZbjeMB1DaCEabVPf7YT01oswj
1rBEhR3kw9GjMCyVIZGmNl56ew5C9Sy/jutdeVtq7E54qihOPNxz+V+CSU7lWNWn
/y5C7PLJbaEvSWdopc0KQm0Xha/vI8+bkXnndb5tSzFARPX5u04k1V72hwIeU0al
Ts8/rvC5qZh+cnbhkzta2Ce+yXvJ6ah0N/DEc5+6H466P18y9maMWwXRnUwf8+S7
z4/xmNV/qwssP2qFR9U/vUYJTr6yyOptrR2Nwj8+C5+TBnrSEWfFbZ507/fMuWWH
8K5c6uFzo2dwjKe2HAOftw20S1r56q52KaW2tp5Ilmx3DGaFPSc3onyrAAqkgDNf
TNV7JvIVMjvKMLj1SCyzpzm89jm8FrQR5H9XolxutVGHDxPzi8Y6kXyTiX41RfIo
Kq/H3WoVZiA4+gRWjPfkYrSoIu9VQG3KyeCVQCF215wkDXrxpDhvoFwIXCt8QCSW
NqnD/9F6sUD5kV49vxf+S+EK5lVfQTnU1GDRGBTS951rdszK3/dtLAXhn6Txqgv7
yENmDlMMP/g19HBUTvYFQQwUzHiP9zi3CY2IF9CUF/vw5+ZA7dxntS/fip2G9fWo
Pi0bSsN4NaMq38IC7Wfi2iRjrPN4pnvpQdoJh7f48rjjHkeWR4zuJfO+yNojjVLM
dK6qs8sK/ozi6PdwBLva7KTMHVArKOS136kK4lVMaD/OylOCKh/+bDdn6bVJ71+1
qYSNsC6Y0yUAtquJeIRWEmhejGuqJy/mbpyRVXcK72CmgSvDggvS2Zu74G+Weuie
Livi4ql3xuIoJJbxB8OFQSM1dB2+a713GLZ4q7+nqGcaFX8xsGDgduXeWEGkT/lX
zov+/8US5KYOgmidqLF5G7bmwE0n3Wz36cJAWymcDvTpcOy7+S6PPfODYaLzfAun
56KEGcOr3Vq9J4ch6iG5D+ceCuxlym1cEKiBLv7aObvZV6UxCQXPnfe95zHNk6Qr
lPz9x7JtxoCp1MD8Def5HlRvqogxdT4tW/F6umiMGrxNor0a7Fv5XHRO9vBVMiFq
aLl1FVOyyeDegNH1+g+E8SK5zQI8Aa6QeX3Zysps6Letiftn4jCJwArA783P6sFx
rmW5H/yEN4iGwgDN//GjegEzEOduMCACSoK/TbMfbnJdPeKFkEHN0NzRu0+LtHFq
jCEGxCsw4DWUCGXZWjmFIreGJvzUgzZoCLGh0R+bmPemz+bpXxYOwgXq8qNlD/+d
hvw97IvUs26Jk/7XCfKAFnuM2KpOi3yvxdd+2axYGjtrDYG8u1tg0vzE1i9dwtfv
f4pcnWt4XGkNFKXIRcNwFol606GrYma34469qOZfQJgafmZ3TzUlnPBVF5Egb81G
jImgcuJwCQc6kNozMbYC0Eb7WI5NawZUCRKEhXzlvucSRvvGDetFsaw6dTXzoUjI
tnmrRcHbBRXse/kCPBlIJtjKi1jKrwGgF6iwzBZGE7uDP+4tJ2PXABRfF+jGIpIp
7TIkxjtQ/Z/a2rs0DyTWf41sQiufRfG/4LBLAE112+6jnk1p8k7TmJ0sJf7fbrL1
1LvU21HFAXUSm7Ra0ZJLbaE/s93vza95SiRRCYc2ub0EB/31UfHHrXw0BNBtYLwY
uXSDTi5cxyDBnN6gJfW2+WpRcMWlf/rVqbpRPyPTUavZT9WodNkfZVo82+WkmkWi
JuVAIc3EaJ8dGsH/41S7gSV0n5lAZZplnOmM3AgQ4LlxMbCVqie/IfYDv+fHxOAI
0ea/tkPIA00/r/c39edx9HSHKaRgoNVqBhX+ZWbQFyoMnH6UOg4U6QAOxi2IdAnW
9H7SK6y1ecDBmVqGgvf4YqT4q5WCqvfWhhEAtg8lNKb0xshMgT8J9rQbHsk/5GxJ
6y4JYcBOYpiLyLuQTQ6d8OHppxAODZz3bS3yVjPtCuAFotLdv1t9i+fcrZXYRC+v
Bowal4wCsWudMlpNYebX9Xk9S/QgmfRJMyogUwHL5JslDRlMOYiBkHCuVyLkHlWy
9CkS5lxM+Cx/H0JGsxvdtWkxQApwwhfIq/RqT4k1vsUBPtmhYDH6+gIgDsux7JfS
w5vma1TmchvHokD0Zg4g8SCAeBDZBSfji2eN6TODi2iJNHx/YYjsOyeYtqbe3G1e
7ysDoHXeyX2Ooz2XuzUCEicecoxnmfdSRxYVlqF441o2BPZ+5op9ysFxtpBG4IiB
w1khq17690NepWMXW477jW3CBW24UMfEpTMrGD96yQprRGDzjVY8hdst+22nW/qV
JBlBhBV1PAFlcCR6RwAO+WkNO589HPLmy8qqbbmzkETJJT+2GzyoYAiJ5RS0aQYr
bdsXtkQ+vUbDkqqNeELKABakgnOh8BCdezKy6c7J/dzHyRD1jT/za4PtQVtdwZBC
Mdr1H09ad14/pOmDDv5wxXzlwffQNqrTpJyZRCRYcgRqVxLHahDZ3tEcsJHAlYtg
k00EZFW7Hjab+766E3gMR7GDSi3IK39wiTelIggkq5owjfN0ImPGrfNVtHH3ozgH
RCZ9W4mqp9hM1uGAiVGHvwuY7vvyAF4dfPPji38jJ374bmqYRYcgxODL3ue8v+b1
bCmRmRdLZyIuHTsfnHIE9cUl3S2K8yGTRRdch8b+IJN/dat0BMSXfOcLOMfB+Ss7
g8PDcuEpEbSOUPEKXrGnWK2zJ4mP0Jy4bqVyhW+6LLGUkLzn2HpVanYhbPqKteT/
jWXFitlMA5wgSKAQuvW8z9sLj99enxFx37yxKzVZkzyBDZ+yWc9Y6VctD9BsBvnH
CAnzgukjf15LtT2uA67MGUeA5cvgIBMDPvdxYqLO3GzEvR2zf5Qsh2RjHygKkarH
zO21Xt1asndaqWKWsz5CHp4xYhR8qo6GUsMjp+YpGfUU0+abBcCXOMwaLIHUkhO9
zBf9i4FdEyTZOAqRye/JOV1Akcwvt/yPngLX8KjC9qmWDYTOh2GpUjR0Iwk2of5k
EYmeq0gSTgTq6zmk+dOSbx0GrFsY99JA+E6VyE9VSHFKY8aAoyYVsRS0B4Yl1DY9
L2F5UevU1eCS8F7bm3N7SJGBQIXkP5T7UMwTZGqyes6lgZRZbu/8beUyXXKNof+P
3TtOCZ+VpnmEcTCwUxDNjKUp1krsTyS/StcoviyEy0n+whgoppHVXfpSBpz1BqYG
4k1kCt5+myCDvkV1lNu9UngU+TB2uWJL6spCYoy86pIdrMumiRBtldyDac+v98lw
u3P47WWKbaG6yYy9///dH+G0pw9y9hzyNDO+uoGUetP1tqrwrtLlev75TwIamwr/
4c0QOGYlnXYaKsQJjhLopbQnDk53cFp9k5hK3QUGsPFDj0nzJIwLyzJ+NSokaQ8W
5/hB+Cu35wiov1/VUyFi7K3mURiJocez7U9x0EyPyXlJZ59RHYRpY40zCFtKhIbM
zYjIwV5tK1Pcqzi+ok449V+F3zsZIOpc9+pCsEhPr/VItaKOLro/nJa6avq0lvxL
wqkLEdWSbQx0cuGYGJ6b/4UoVjDq9orUbdD6+TaeNo+FerlzBz4M+E5JabK6HIFM
UhmObiHgaHq25Yd3JJjBAObyCKDDRyIYk22xbVdL9Uvncl5QePfUSF3u/VkOk0kj
SkskXFp+UtdanIm1LyZa2j79mEKOIKaqJySWmA02i5UhsFAsFR2or2IcPP0yOTb8
YkiLJlWOdnokL1jkSd7OKX4MvIcgXuAJi1xR6o6QdGHZAeywhOu3eOxw7cIAQ+/h
byT23rsL+vVHAnRmJuljo4wC4BkDPTilRbhL7+UcwlkqtLyiVvdwnzTpl9fgDwCx
gqm2abchNbH3ystd+Wg+MMQduIcKfD+OhBk+dth8RsV20foJ5pXDKjFjaOmM9IWy
mFw2oYQtZCEfILXA59V7hX92g1NrMOs9s+GkHj4PXy6fEuRa9w2Ys3WXSphQKz3x
ClARaFng0EnKP9F2fPrIZVeeynmUKPyi+kK5EJfZKuw5+BJJNJGZf3uF1s4u8VrT
j629RpbTv9kYetoORbQpA7HBxwSK57D+6CgHfAnZcqOStmIx7HFqK6yItVHq8mSq
2sTBLLXKc45TgHug4kDzvBQyVjyTHDEfMPv67Y/k3UmTlqgo+9ThR/7iTmxxgski
NfPwJuTDCvUiXtH/Q7UGiXT6DmW71tx+XMjiHBrK1Bq6JBr7RdS6MrXnG6I8jYGH
Jgqd3RYFgEG4n9WlmexYf5jVRD51FJDjhRS9ldATQEO3lotbDR1axY/WG/a7fE7i
JI/i8eep/EV9A+Sq6uGDbeIejgKGNtEcrPFFIrx0I5mXTmCcfRVJtSXXfkv1FPUI
h+NpNHn24dUuiKfEHvpwybS+N8NLRkyagoLqdcggD6AgPX206JCZJ8HF9Z8faeMo
Fk82S5X6lczxHqT+AtXoo3R6a+XbCDVtY1QEnB8jIK2DaBNeo8PWiAUcVj+h5mvC
G2NfKeZY3QMuT2Or1LIFeaUgzV31gVQaO0odflKzD4QkikDUh5WFlxPaFVBVOtTC
OQ3FNde66+JF9Ge8SVlRth5K3Ixg2rptCSn9fRncbqXMjQn6UWlkPeO7R20GAxsf
MXUtxIq2HrBwN1/KWEn57nxxeAIhZrrxuInb+MsG0bbFOA7dAqOHcHNk7dq7Oxe3
oisr+4Qt287ohCCvvFjpMESCogg6MVMKtwnG79X0nj/0L07q+LRDmUKn8RJ78VDP
XkXgozKf4rRNUBG4NFvqJDE7hvJuJKMgqPZfEKOFWI2lxG4lDEu7zVQn/mebD+r8
Ah6Np0BBjpU7n9vVmZN0HBCpUs4esK8CJrLvnxGd8CnGBN4hTnrS7UHuMTqjog2a
gHJuG3nS/PMFsmokAFEz87zIXCPuL/ZT9lxazoavjgG1n7prBFmgnegADlN5SU0y
K59n1edh3XAc43q/6bnbsB/5YMUoELsz7aJHMeClIQAFNshbDpGd8vnqzXjSDfHE
dc3bpqv29m8deowfWR2n72Rk2AuzlbQJvjTNpAN855nmJJbSqVsoK9bi2jFvQo24
X8PMG/kq/Z4oDCaNcWThGn5uYniguvQOXbQnOHPDWHeve38JjyzjcM2YEVGnHV2R
3vxZivaEEb1lckaMOyp8tdC2s7rM0kadUNGGBbWXxoXR8VPIzerNvEta+pBGe6cg
ZORK9N9P6XRWcVRW+bi1q4X8VSK6ZfHnnmhUPyzltnKvAJM1hFtTpUXsaFvr+QUp
4RKOtbk1yCj6jF4cQhhktB8DSwWq4nHMT87HhjYuJFvLSCE4zlo0CE2BRxNrQbYD
MfgZ2hggnijQ6ij0dubzWgcxsbCPCzc68vzPutRX/EfQCkHzp4E5uBqm/fOpwYXO
bOL5BloVidoIbMUr71xKmc0I0XuCz5nwgiF2ILPnrVG20ujRRuk7jb+ly0+Lq7pO
AdIEIUNZou8zZc7BUqsjBi1gO6TdBBGkBzUAmID5JWgngdaQ0ITsTnOCoJke2IWJ
DBCBfC7o1oUsD2H3CV3W3yORxfgaGzhRpe5y2BelkDXViEhMLsO8plS6of8AvZSm
vvM1dBAnIi1Oau+YFCuHp3nldx2WKuvF5fbAIqrZ7SCYhReXuVlKT5jwlhHrQj9z
42NwWRG/hZ6l0R14DIzBct/aoLiOYn1ywlrwDNhCuBN+0y7oydRBiIbs8nR040KB
fcmah9HS4+PCmcjTh1m7BYyQ35doBjzlWwKk4JF6IOvNYPw3ku2HWx66Vc2E1f1b
g98po+6U1GIFhOQ9Eo/Vo8Io+vkLVrRZa/uwYRJXaq3fW9xDlBy1Z0NkNKFDuUUe
SqA8KfPT0taLnFImTBhTW3u9K3znGeqsrcDhbcHUN6/lAJ8Cwgv+3dPbIchEaapb
0Nj5sYBCb4Qe7VFmMFGyN/FRNztpEOtdGSdNOI4prL8J8HOjRHv0TDt/oGQA5gFg
0B1J0coTSdSQ6vM3c0NVcVnnscbLbvm5xUltkTyRDFZYVxwcugvHLrMi9+ernsmw
PhT+vQuezoo2B8u58yXWKNCIiuQgvT40vZFntPPqDKXBc1HLaYsHOLiBbTXqKAs8
3k0U2w8SZ4/j6N4kklNGQ/oCSy5SKD3ZGGW225xETbzs5tB9A62zxjAR4deXJVEY
iawOM5MkfPyeUsFr3sp3tqGy1IGhh4BAgA1pDFzg9rD0oJXk/xmsb976ASrGzEVB
P8WSJRxN+gXfvB2Ab4A94Fm8fKQR6HjWV4h02sySIl0x0N5q8dBNuPJUcHwvPqsZ
vyh6zia98pe68L8zIRGrCX/mHT4F7TOFHJycVdZcbCZysmvxfE0KerMeoQa/b//8
6R+7F/Tf2aG5w9xde9S6IV0D6xEuIA/etL2obEbtsz7XsCRc/5AtqvBePVQ70/HK
p0SzcV4CqCWnMBmGddI9b17pkEx3kCfAcVMb3Bvbb98G20/1NoDOyootcIGDi5Ji
ZW+iny6plgr0gq5t+oyLuWaYlZeWPuy5SN19/phTTzdnPxZ+kOa9OAVdOjrrb0ZP
WFl1r3OvEUa79ADMTCxkV43H8oXucFMfteHyjeFdZQVa4YuzehuXehHm/4PmF4U0
uvg+/5USzCUPOQcu4xhXRrB+4X0dYCDdwrzYpZyQjkq1toXLqTmIrQ87Jmuq3c6T
sCqEWPp3G52fAINz1rPeX6VcWZErzHsnGciAuGW5hDQldxF2KHpf+tsTo1C44lIF
sQa+OuE138L8ukZrZ+F0GxKs20dwneGjehlsZHCXAQI14ou1gKqxmbemZB7Fbojd
oNLpCh5FbjjpfZBkyku3/cOhUzQ9YvVq8mWtyBzzZEXTZe72I9vIFpWgrDv5jQfD
WZyB5V2L7b6vEve++o1AQnYaJHgvfMDXg9FU1cFPUUWHplm5xi2PBkXyi5K6eP9i
4RgJ4stDHW2jUixA/GLsA1W9bWdNRcxprrr5sWP4DkTuiDw06H6dosmMlG0BgSya
dq3dSNNtZ0mu/bvMpxoEk+cd67URT6A5ZUYgdONtt0ujCDIkCmkbF4CAS0aI9ZDl
vjz5dF5jdKAWEHA67xcwYjqyeBCr9k9obKiqjgdN2fqlRDzZDRDW3+VAxJeKuZJ6
V+air8MRQgvfBlUnb3aybTO5rHEnlYa8ewrkCiHfZ9+PtH1pAQYWp1+dAz7n6uBT
m00WAyDcH/pa8Xxg4wi1qmoRqUjeHGqQhoXWGsXzeDdG7QWrqUiUMgFsdlR+TfmL
x3wz9HG2tpYzcJAbICdN4gb1LwRYNKovqQGO0ncid0Jb+PqexFTG/AP54P1LljV1
T0qqWaHsU5DEoUW9raUYcJxU87hmHx5SuV9HUXIM7IPW0taLzSV3WxeiuAJy3IM2
VGDH2RaKxG8OFTZRfPiWz57hilTGy77+V+RyLZq7gHIzDGTggGBKKm6hE4fMJJ85
ihXy0Z0bnbgWsSFNEt87fT+gFoKPFuIxrbzzTRZozsaxNLNJUmFEGja/VVmHbsWG
j87YtvPnd+GEfyg3MQNpHuf5fdyUjNP5HJKlKHHl1QxtHSPFTs/7XEBgxusyGaFi
QWiRkJl2N/7nSAQdBQxyETW9dVUcFu6ePkaQF8VjjGZR/b3hNv9Rz7ylzaYmHGdb
l65MmLXqW9scXQZOgoTFNPRNZt9U082zF19nzM5o6m5JI3Vl0Uicqa4EAILkiyaD
GF1UCquGhjcnnbqySRZhf1SYtQEM5/+ey+b17hhZXOZ/s28cm9qFPPehQOUjYm7d
3ji4o7wtMN51solPV05L8ayD06+TzzzhEj5l6qTIGggbISmp+s5zoQTpk3PtCnH2
xQIPyAAYLT4CUby1BUCsnMaWR7lKS7q7BHNpaV/fS8TOS62YidgWcnKPWhWntXda
jfU5nL7p9YxkzeuaALb2/pr9NGa1+7ZzbUXlA50V3UCNdY51ZSebcJ4ODJ6KA5O/
WRGAYyHaWVUmK5Uo6k4O8EMz8hsoV/0i45styrfdQ4KdPO62OTovnhKW1QAvxsMK
5UKenfte/Y69I0NmZvYqS8zfulvHV4pidl15RaBsKkPO5nB09L91zmU8qOHphr8u
/iVMKmMAofPaALJcu/OdvDW2k64Cop6LuRyG3heBDmxl0erXEs7a1Fp8r741WzcV
9lkHeKKjXhQ2L3RHfxkahj1iXZrFktBvmtvWcF80eeUUyeSH2OZJ3mUFk333e2Et
yLGijA9yNe3tvVxZwkymIh8lpeUW2KT9qxY675PJZeRopXmqIj+24AmbZvJdQhFO
fN2Xyr89QOcE+f3BpXy6vHZ+r0V/khq9THFUKZj5WQaXMSTcBNkK3E6T7i6ldlB3
qQjiURsSvw02WUl8r4hwkQZnkKUpB03jeU2o0MkIfBnui4ZAGkBxfNhXPnEoSvtW
DNjjFFmyGwXlRphGdgxZhaRV/m5HmjKR0122cM9UWMC6+5gchWkIlvT2EbbekcNz
8cZBsB28R4aVRrvi40wJ19omTb+ZDwqSC6rgXPSzxsB3OD9dR8CTvQgniQ9u6/8P
TE8sqChNp557igK/L2DA3QZwX+tiwoZh/ul/ufgMl/NcILkbXCO5pq9yzS2ryFwk
FxJAu7REVONpl6q11so713D3aFXD4dyreUpoOJ04Tm42yGycvOw79dRJykZyItQs
DAiAQrtmdyOaUc1bDe2PXTeomwOKtb9IPgi3jqrt/aC6lndapHYJ0SVqgJz8gmUm
of7jPbsOVP+5DA95bWPzt6zTH4YEasgiyKwY2citFkLSlRkOdL0LJmnwyII4zsm/
SXUzb7MQhujCZ2qnlXw+VxduZpasAN/YJmFTrxo7kgOjDvGYxLBxxuDybsMW0bCa
+tGjH+HXyqRc7+Fadw3VNupRkjJUQr8iqgx8w1uM8oK6eL3qs922/c8NpABSzopN
W/osNiepsm+zmiBbcyOXIGa+HLhI9/XjqR6501V/kLAwfK4zJIadXhxYg5cy3MxA
c/HMny+e70hA3MW9CecS0YQAB0ghNYIewwdhJxdjDN1kViJmhSllNtYsAqlfXL6a
oOc2ogS53r+wZBK+NbmelVjScvRRXd0JZP5ADgJwXk4ik5GkIRCwXQ0z72xVdS4x
rCfD9zr1uht76zqXFjWIGT1Zvmho8IRssbUb3519L5ks9CM8a+wZjJ4j91vFvwZp
X/1tYvfs+Exc0phpI60DmDr6maDzbmPHjVHo5k2DQBcyr48/g5j4O25i5TLifJGh
R4vZuvu994T64s7XszqtUQW6kXQczitL+ioga1GF6bbGzV6aj8TjQNNGOMhn5VSG
6CxyCrbtuXVZGY/lexIOgp1Xhdoeutx40eUeGFf9ErVp5FGKsTz+ri4YsZc/13dl
RahQsyI5DILUBbOKsDyhbDGDvtryYWTizm77Pc7ceHFtXaohz7VZ4dukhQPLfXv+
xj3rq35QseVe+++xpjHyqE3jTfKoqHHskO+DFxtyGWqHthAakOCWkU4oVgqWTRf9
TySAv4UxowaQT/x356A5ig3zEh8npX82JHGSzs/kh5g/kidaPt1+pcCatg/dQUt2
Dvm3phBKeZJkTb+mMSZe2Kat84R4bwtf5Gh2thwUdnHnb6B3CjYeQ/RBCdDP3OdM
CxYB816UKjUGSWCMUYPnNOHAvjGgfyMGMoRO3F0zslRX/4466aA7KYclGIrFZx52
lnsNRWwjlGbUIrcRWfm7GrSBTDt6xUM5D4loSB/d76pndreeN4OfSaFSwFeLHkAw
86m9MYqua3G7cU2/xT7ycP79zN0pW2++uYzavP3+e5HEbhPewMbZUkMDV3fNSFRz
5mvzzxywXwM74ioBRHzIqt6QIyOQh4PhfczBgOzZZvRPjZMA/lhlfGh7sHAex18+
fBh5F3Bk21qz9hbtR9hvLvwCiLYOUchl4EmZL3F8lTYn1mh6bszPrgh9Wo0Ay4/T
Y9RlnJ3eyp0ozwTnZvpXxHEGdfbaKusueRL9lphn0gTJzHM7mzvyIKr/qREghBQw
2BwMuxAXTfdGwbzyO24W0hNUxeEkkrjimCltrWysOaN92axrsvbv4SqLPD95Zgx4
eR/ZAFlUQ2MvNJOY7IcxHs551OYNyD216gcYnbBLIVlIOXHRMaLAqt49yd1+nERK
0IpUmtWs3ShBtIyFJxp36lFwhbr7njIH6U6Ru+Ctd9FvfNhJdEDJQ981AxAStgZC
cpqDnM54HbhmfGlm5a6WxxRFsvlhToVBSi4bg30QN4upy5EjnGM+6iCeOMKh+0T/
OaLs3GvSI9pfFPm5vwzJ8Tyhkcfz1rqQjhpZI7W9ab6Ubf1Vw1HLm9d11dUDjsla
lLet53pN0hDfcyz0TvqbttjXEjLtrnbm4GauokKAFcjQ1d15f+dybUTfq2RINqQ5
/E3Booatbc/1Rh+H2lg+BbmfPcXYxoyzFmbuexky8hkXCrbzP2waQExDHgEknHop
VHHZf3T047KmabpRfs0oQO04tEx78j7e43whYaPRnNDqvjBeOCxCOF7rqsuifvdg
wLD1H6pbZQBMCBgzHVVhF1gPBel0B+LBCLb8xxmg2Vce0EU3Ribh/ILIZ1i/BFSO
CM6QErxXR+s4v3U/VrohfBegTmYINpXLBqYaqoiwDkhnaHCaObrIm/XfvfdcKF+z
8JFVrIuwxb6vmRtJJn5w10hZ4j+LjiVbss5xog7EkeGruYw9E99K77CDk9GUEUl3
MbqjYdZg3bmGedIJNsHhGSbw0MY+bHeFT5n4V60reSQR3K2GISS/NRogwhIp8lU5
6z1O7OaHDVblPLk/3CK5sJfUQ1PfF9Hgl/8E8ujUKQo1DXUe/6DaeD15HOw+OuOR
JbHhE9i9o72vP/eX+b8P0NqsN2Tp6lYXYgt4KtuJM8OLkuv8Y8ciRsZikM9Hxx69
PYzwnOPKeCWgkPLHurSVdMw+ikY477rorRbz3Z6zVSuwVMh+UWEnNwKVrY/I91Bp
ZDAJpnv2aa4reK4Ej2zgRF+Lwy/uSKo+iufDasyTrK7GfuyOtU7EvaZLEjjLFwhz
vtggo9E27N6gosgIGHrbJ3PolI+CzkAAJtFohQ5BxtW3dPd7tC9Pi95387zsvgg2
Rl06Iig5SJvdYc7Tv9Ku1yWeLFrb2TMXaLYwv2i8bJeH282bD+CVpYN0sijc7mM8
ddKSafmR96AbQve2QOvJfhKHL7a8llsLN6DPdBQW8QKaFwvrwzKa6k9fGFTfi8yp
WBd3Il6Eo0t4C/igE+IY8RjOnwYIUuXKSptnJOcGzwT8SztRUG8xl1ecWoXUGCo0
UeM2yXb7ZmThPoPOYT5rFZJqbNzSDEO6xpm22OEDDQz97rliTF58nXqxZUbQcuPM
IqGsfFRxCUTb4D0Xr9TIQOmKniI5W1pXkpwV9nZ4Cu0EUn6RbAhFPOm8CvE0MenW
5p5gL0QbBGwT6PIIkQSLvkGUHyY9oUnMyGZuuqJ+tIjZ9vuD28o/Bj+c3aiHzHTu
258/Bt22kVo5KhJ9unAecOGJKha0yBATgo/Czi2K7hWDyxBCHY1zOz4pAJYXVR7P
lo3DwrN6XGgEupTun1AfyoLxQPqCfPWSsHPLbtn4OA72zUxToubNZ2s83CHdqv/y
7D8OU38PctLgqkXPv0d6YBjAFhzOpgW8TRYmHrJ1FRALQL4igs9xOw9mW+ExzgwP
qyA1ADY8vHywc2DxG27YGvQk6WEBWAUAXAlWxgxfgdyADxdHDP5QlIGE2Wnyo0wP
HTCzx/qNyQtZ4kSd+0DGcfEcCrEd4TuXtmuzVFqsxTjBoT2/GeGEYdbPZU9cQyDX
3IisaM8nURRT59UqTKM71M+0+TbJjSlzddcCMq1pRhT0z0RD8LiZCscGM6kUNqUX
n7nOfReoPc0gOPY56mB6TwD+NIhLomwa/OorzQBMbbqv7nnXPmlIswcrRSJqVRid
ljnBuQJTu6PRy8ZLfv+Yeu5hezVWBnLCKhSeDcRBj5cS0vCtsxveNgV+/mt68weG
mT7AIgumxsuzpo7DHo+QVs1BaW7lzmpaVBM4k92Y+1aXYACc7AXM8QEYdSENxM35
Er75LngMe/CE/SpBuOwobOnFOgd/hh2qMw0kQl6gjWsoXTNRAy6B/JbGj9vDp5+O
rQ7cfAEMWYAJsQsOTBWBi/0IZPgH2xVvToh76k86hHy9brPZbdQ5cVqs8AwNkPkL
SVhvU58xpHN46PhzTNeosNsz4s/zSr04mbqacSSvqt4Rpf82Zmj/I/pYwo48njiQ
a7GDqReaixVzSY07cMX92dJnnmR5uk+fy8LrxmPfiyxzuwSKTJL56RfenLGeCFC1
nvaPyowGtN3AF7rWazG2lN64c4C3incCkiOitTAX6V+qSZQopcC5DJXJ0FLvgswF
aj5gQ31R/gCYX4NAcJHbT1HlyB8fpjYiOGi0xiAXT76kOEGkshBQXKhD+XpYwRHF
SrQtMk6cIUOfJMPEdE1CsoZ5Zl5AYu02JGuz4UimjC1W3RQ7BsC9oG0eumOomHMH
UKXZ/Fvj7BqokxLZGieGh+159/FiYwN8Trn78e8bO44LIKoJvIUkjShhGBWLHTvR
X9+2WhW5WYVXCxxCRmJGmFdjKBwCgt4ChocKcOmvZ82jiNim1NMZ5tR3cpHVyHTl
xwA1HUPy4kAAcu+aTG9vWJ1FFXVP4WtG3JruLOLWRqvX1djpd8NJWRethyRR4D6A
zqh/6opCWXewb1uRi1thD+rCcxdKYINMaZj9O2A2AO0HY/osQt8xOaqmdnxUa3ym
RV3XjpwtoUj9ecLDWQPAJD964HnlAc84OkxTcqMRTDaI1R2xkWvDOzpe01sGsiG3
hx8NUK8XnJz6ZV08/aSkdg6ETYYsp3ZxYCrVmaPwfl8WWgBzheqxjzHRZGvOcnuA
S16hypYm5XAHcZ2hyEDzO7ic7kwCOFF6EYY9WkNRBzes2jZXL4LG8tDBiqFV6niO
aKb9d3C+0+tNKoRBN0qX10mPrxhu5PsM6ObQrgDmQD1Oc+CmoJAbs151fZZSJsLX
MJ3GTVx15ftpRDKm2CGE6TN23V0oRg57CTsSyXPV/loK8sMLnXymHobDyvrDW9f4
6AWJR3JQYmf/s/0YSbvXf2FK6xomyJV2MSfphCHUmh96wCH7O6Lm2iANX0ydr6Bn
C5mU5Tc8hpLgwv5vNaO4PLNHaT7dzg6xwnAdILoJwEQMTYN9mXG7hmmHwJzHFv9S
gAlO4WLjtXJIFviQshDVrK+e37YySwYj3aGvyrMCt/ecofvS/Z3hQjom+TI1Ym5l
W7yzn9PTf1O7oa0lAMgWQ+MmADn2C6AnGSSaiD59qmIJpc+J9GcDDuww/nsv2ixE
75NKxzDQI23mkEDg5ovbOtNFQDFUfSDl7elk5DBv6Tn7y8UQZ8et4OzPb9oTy8MQ
9jAQ/Rjt4FxxufHyK3iEdpqVDqO+VLLAna6B2dEfxbKsQ6IV2WBbLnXzQEcoD3r6
ZZZiKjz+I3cPil4bfICFdFzPrih15L25vEzUYQUylarBJZBLXGa1Jc587qUwZ4m+
tSuBLFAqzOspRnknKVEbKW36za72f3+DxjlvldHZ1thXqrVCKWIw8cFijEFNjLWA
po49nSoM9/L1gNJkr5Pf9dlG6OVsc/Lc9VGZas27VACgYfAY162wdGNqXd+VpHOQ
mG/uMiv6MUvWvMFr215BEZCPK2yhh3Pq8i1BMnhl7XYQXl5CtfL949pWYEeDnQug
wjsDI7/SOT9xZFi4uGFMURHBQqHHZCse4bTBi4j9tWtF/dXE66uU2Z5Vi/dciSOy
2iyeDUBB9F75IkMmgTM/ZE9kLuSglB6fxiBGArppusDrMbXbb2aEkjlaj3iZ1rjh
gJ/f7hCLd3zVw/9gXYymxcDGar0n5x6NIDPIiJSaZmWiFaMFfecGAD6LNhxxZiEQ
weywDhh4JfVQHbRwsUnBdbUT9kimb65FKGFApzdDJnqWYozFxs60Q2KXMqesQxFa
ZJpj/vVUAnSB4nuaOTVx0lre4R9+WfAfbcSYNTZldoHVgoeONDJUvkUf5lI9O3Pa
SHRbdCapMgMFPapWryJ5ptmWBC3HWd2TUdHF/zDxq2kW2fTn6HtxkEBiSqEp7hvH
o5uqxGF7apejGNZm3HKPtY4ORk1PPD+evYSER0cZtOUnTK+ivJw313hHfjwo3hII
PuGRDSo5oFdsZl5xkcXvG+RwdPCDzPEu0hEzWJtTFlTUW2V9Ui6TsAgAPe3qJDes
mDsg7dcQ8pG4tKaJuS6E4SIs7msthUyNE9j/gmn6bFCHEboNx5WYzTA+mQLJvmKX
BCzPY3I3RkB0rc/q3LtLaBPkTQHdXvNxKLOwY/pIpvZ4QEI1u4zzvXFVkxbqQDZ4
N3KHZCQFnxNJtFcv64of4RgXfoOOAJzyIuFYXz+he9+kjTPtr0OmWlDQ8rtfzqXw
Hpr9+lpO3RUSaWdIDVIY/iwNSlBtD20Q6RvRVvPxAc00NasdXgv1fDYZJdhpL+/B
+4vowtKz2mm6on9zRdtIzjGheXOn7apXqn9yvMHdaM8jLwAQpvYvawHBUD+h83RP
HMeTbDMqf2YLhzGHJkjhyO93VqklUz3dDERG0CWLg1YF5ykpG25sEqWIxuh9fpQJ
IXsyMamf++6wSy/DVO+o+4XPTERTow7w3L86G/jNRQK/DKp7EnnVmiyx0V6eRQj3
/xbipMxev5pfCfgy57iCvGETTV/C84+TlmO2234CEx7btF15WEMu2y52aoDGyMTC
Fz19BsxfAMSNcX4usOaOcLzfkKEqJY19yINp1GH61py4qBII93V8NJNpcXNV03cb
bwJSsbgT52elKChVA8+gMKaczA/u6eUCDXB1YvDDii/FjJkQW5/7omVhWkWdBq32
nh4MwkHLahxuazqlVQtv8HaP/q1ofJGl91V3Pcck2qHsU08vPn7ei9FSTyX4CdmH
hvjAqUah1/oMAvjaprgdAhwWEQtempeH+Z44HF9wwbiwHvY+V1Z5UPqw6JaTizZE
m4uMTFtfM5ws+SlaiHX3cHZSgsGhkUkeeCaVpLBNN32jMLiBrzFCABu1Hp1GAtIB
+nLUSugIEGGQ2PvurvJ7Rwg3w748GUG8QhxooOZD8F1otCukwCapb5ysc303BgH6
Y/VutkAn5yLYlL8Li6Pq3oVXuxLJSyliDnad+wBM2P9E5OgDJOvruG0ZnWLjVMl3
Ns3wmG5ahICF33+t7DcWfmJDYBqALSIje/8keVuSXnMxaJ1rTu2qd2h04KeRUGoJ
ayX8A/FZnsnNao38tt5lTnCDVvOWgGkDO6P+InNJTnQGcXOH/F9QJs5A0eI4h5OQ
GzkGWh4bTAVDpIkvZBFXNudD+sSWek9GyVdOjQFKT9lb+0kN5thK1fwG5xyN1Ygf
1xDt2i+QtjzrqfbTVft+T7/Hf8ghJhK7/Gn8oJQCbhj3NAASjxj3zJNLQPucO5cD
gBNyn84HUAhV6nNW0lzKr6nl1UdDIED1/qhNBlL3oz4t4DwKONzMrjeF6OQujN4T
PJOBWb+DhXeBIN8hEUppVKlXx8bW5SBd6VoLRVk0SRJaxmO96gopu0ffwGtVI6aQ
8+DRznYNjASPFneshwD2Dcc92v+LCCv2uHZEr3Rx7o3PNpeHrNyevQrEEv6gByyQ
l9gPl/xMjhWzNL/1HQJwnqZB4bfZQe7XLzFbmMhvjF22+tHhtYyjRYAVVf3AEclz
Y4L7nWtErORWi5H6wxaodMl26idL80rghs4OTQMfhyiiQLZT4WQlLg1s8Aj+r1xW
n9wZxymS+HnfHc0wbqN59nR9Mq26/RrThl+SC0PsLbM2BAK9w+UtOHDhRhlPejuZ
mEsPd5R9Z7tCCjgRHiVTBsTFhU2VSx2L3I/ngpR6SONm0NPgyJjEaeQYWJ/JPNfg
zOukf49ICU33CJ8/wYYXAVs2jJkqV+I/dhKfJmI5hzNhqrL2YfxCQpjvmLkrUqPu
6tZ1yPBaHCwKUGcBgzZsoHVvMHkDZYaFbljPEwc5RqFcoErz/Uk1hkn4LIJ6C7/q
/E4LVtzSZsmieE0xZ9KZRpiZGCgQmaueZyoAgA+NYACTzwIYUJIQ4LH6RzzGcED2
34lXa/6nZ/geOlXsrvK5FnfGJvfb0iZ4M4/qP1JMAcrxXnFQTI24vY3Jsfa+VMv9
Q6ANDMnUNi249lv6cu8fXkwi7lyw+/xUawCl7FDVi2AN54FoREOG7mEK0QA20ix2
V4L2oLdrLMvS15cL50GFNXC/FKsTqj3Y/mlVGNI5n4KmYxiJm0d9XPkjylkIW0nx
AEKV3rDyWw9+3DlD2zTrd7H0sSBI1vXteggQucXFdVhUcYtMXRXCBa0qhP5zz4w7
H8t448v1fPlJ7atG/UZ3ONjPi6wgmFVD/QNDCETN7sK3VgoHTWNhXCkEwpdXBJ/t
YPca9gEegqocVIqYw5m2uvwHLqyK5yvlSEaEcvt42K9NJWlrhuUEVhbLRIekB19Q
xqGugIleQrrXqracX/H/RmuTb55ML+Y53KUpfpoYpjYtlyjVowgFb115pEoTNDAT
z6cgsK5QiMdBTjNF2nZUfw/BMYl16+GvWVY/LzO4dTV/ONEplWzQ7ztnSKeLtgYj
P815zifArrk3tGIsT/wL7hAuiBID0X+I3hNF51mVs3zDT0rXIn1Ya5CXR689sMWL
JTi/T4nc6t3H2FmbyWHwIkkJ3ETv8pMZSw8FMcZ94NE8fwJi96lKXSTxoJxMUj3S
QLsqF7znHXqCnjluobKlcp2Jgl5NhzpkxuR/zeOGaflxRgI8ni6dnup7spb8n52v
3hW510dX/c3MuAMkFC6WZbAGGZ1potAFMVcJz9Yo/H+/3ZJC6OKirY4ppwnaefmf
m/abgokRKo4iG2ClcZrokEEjI5n0M5RUscW77GJoSfSX2AcRgOa2pNo3+RZUV3aM
+bGw4U30PFU5eZuaU9sPbt4SS9+RWzJNdmGC6Ykn1oB4y4mLzXzAt79jvudZzLw4
yJ109N17asXmssRvTas1p7mRoIMZwuIT13CBdGSLLCumBPeNtnLEebBzAoucvkk8
TZHuf+SkEOwfEOCOpIGraQodV70Hbj2pp/FI4ifdp4dygxOzxajNDXeNF70bqJoQ
pOnxh3EJqnp5j7z1JGXKDcavD2V5a2pN1ieNyQ5yGhckZX7kKluBxgCELRv63TiN
BjsO07q653s6CzSQTRRyUvh+6KbOV+FAmMlteRT6oeZYeEl9SDE6XZECCobVobI3
EXRyIw5NhL3ih4LX8W8F5TyoDHgPm1ttAEbQ6lByTs/InEbRDFdufr4DVWlUVtz0
/qnOj5yAlRUTEUVKBeO3R2ht5uchS6I5ccSEW9yo44vb2U9zZWmvHo83DUv+o6N8
wPCMUp4/TpNIzSacSe+nXHugS1bQt7EJjsWHkQ/WQBcGpKuEFxNHZQEnDmjzE5yo
DJRqxbRlwA5ot7dpGEEG4JPhfQHFYrL+d5ovCopDxgJWfFuKsLS6eHfA8wC3obZK
52PULT2VXObtXzF1TMNBgqHpHPNZf2DDz7EOCnQKuZvP+puRkxg/T5rL8j33ujvI
GvmCZGg1sDR0EpWa0y29x3GGKnaQ7h6nrGBWDwpNB6i9kXOe8WrGaKf80gWpQTgI
1mkc4I4MpD5t+GYmSHpEKW4vVegWJX4XT1i4Lse0JmeK719OKKPJfMbtsvRXYZuO
LLaA4d2t+kJlsfAyUFEkxELndFg70jij90Vf4Ac+6WyAJioGnM1Of3KoFJEcd+MN
E7hE6S8Q5sYfTwnCJntksTIKFmk9Rpy1rUWbmLAJ0gMEalONrG5cMqZRnetpBU6r
j3jngBfQYXihmrLCWOxEDIgJtwZkkgEuISX9JV8igAvaJhTgDxeke9n0vvouiF0L
IhusYVsZ95dzqaXtTZz3iNqQJAvj2uIFwOwOEelKaokVA36fktQTZyKN2OiQs2Mq
iSIi/zNxhA3FgUIRkOWZZuyE2+UsUxlSLyWpBbgmsUAJyJI37VqnpGrn+bAsgDpV
A6EA3kt7577J/uScERUw+zxghtYcEC1E0thidGgZOrhxtEn4fRIc7PEYtUkj3cHd
1OKIk6b6RAPOsIBbsCpLsVXEF1TuUavfWAQJvVc3Jb1ZVmtmVt3jsh0XkqM9GK7z
ynsjNqaMeGvzT7j245X5MriNl1/Q4cgp8wazid+/33MbAkUOwkkAgPavT7cISwf8
x7xAmsFxtR55kZ1UtZ+TeldQcOF0iGBa0Pp1MUZCCWcRRGx3HEDUupIe3Dqxcz50
lGM5Evvk18xpww7OMGFGbG85ol+BxqDPzOQpIZFg6eX2P6Z0/iHXHwPiNj22gzGe
2DtXl5zx5MlTnwVAJI95B9CI+yHJZF3UnxVXxf+xmcY2FwQ4FvI/KuS+TNj+dYwK
Q0JEgyGkLSBENfhJYC3Jzx71kNhrqk+3VfUvxoYyZ6SSBYnZwI9w9u2diMfPlCCG
quzn8mTnPeJZ3EAHIIn7lAzeHc7AxjCP2kLuUxob8F2Rx7Q3YkL9K+CJb2fFp7wB
c/9lGR2Lguq7TjnO3dKIglJR9tMSuD0zGAiGBM+VFObBLJPorwiqFjTh4eiWPrwY
EPbnhC3Zbqhm2Mvt/8ZYrpwhljNIS2iU0UF1RhmbNskwtAR/LapBpGd44FS/IPGI
TpIXkX3CaEi7g627qY/E8XRRz0xI1nHiRjhrHxNdU2Y9PUSW5kYYIdEtOqPC0Nx/
zB2UHPXvS671VSpwSgY3jGEdqRGDc45P6XWmdYW4Whd+3+hmouf3V1NlSmqiqdSK
LAt0C2Lv8ROA34K9VOEn5cNip4uVxnU7CaUf4JH2UqFOCGqkDEaWFgVKYmUmbZQ0
gb6AdEaPOvDj88oeu3scYIP85KF0eggzH/RY7QK5tqH81kIJE/uZa+JggRzxiL/h
EPWbbrC6LdUhkwGB7feUX4dYCtLBqQhKLXw4pSnHRVQJCHaA1ZcXk7UOsO1PG9wW
mmgRBXXHT7GlOMOwwYPu+NGqkYrAALfuj+woVfs1HVmjapW+cMeJT+nCxbt9c87e
zjAb7bVA70xB1hi0nV9diUtw7I/pmzM9fUzRobzc7fkWIHAHlgEGnNFCAtO3LlNh
lgDdsO4+XvLjNfYMYD0r+6/Of9Oc/FnYyTdRkNNqbKyqv/ELX7hgPKU6MLfYk4jj
zn4JsRX97KuUx2CbbK8HixAR5QJIbmmf/52SSsD7/JPgtmgzgA8FwLOPMvd+fif3
r5IwM5b53BaX35OfphcTTDSFe6l1Oec7edSaonFsyUtoO4RIMmBZbLGUxMnFgSNv
rSsuDYekaVuVDgGwG+mksP6IHBrpW0kq4SnwgPrZeE2vrWkXOBzsXzmdYbekn2jk
6kcTHDjTBgfn1agRf/pZtAf4/uG73tAXDUzqHOgyR9164/7B54BJvGkCMcYkLHWi
P6gl+KedNHPyu4McJIeSGHFYPGSj3xGhjb/IdZwvyomLJMdVayHnHlccly64NPgR
86UvMigPruvrBaQ/AAtevAr31ZZCRcBiIrQSFmLZNVIV0nOfkEzytn8MF1eopMX/
kPy3z4E+W7PG+y7A5dPgLne86sw3+2FHG+tujbfRnju+LNZ8PDKoz3Pfai5Nkly7
ZVX72sfiP/WH7AjgdH1ifPbhq/F6xTx9a/dJ0A6ycNxeE81tHjS0eAbGVRgC1d4t
up/ToVblD23N39poo8c+KCORs/NYtylA6nzBqTAVCDqOeNSSvoMLRnf1SV7SoWcA
7po5bPsAQlUCXUMuDEYkBUhEiG6qv7VFSaPP2nGuhVhcF0Q57bNILsNujK+y8YeY
jqikhTuS2xKhSMntUgQgRohrTvNuFiGIDSDmBt+xZeuPyrZSIzegnHjXpW/RtSgU
G83dA7taqbwh6MMQdF8pneu8aTn1GAcwGTqBkqSeTjEx7Y4FVGhk/KQ6GK4ZLlcY
YeSp6yxrkEkoRXju3B1TT+tErhE42UOXhGiWdmy9hTuKcfNBiPNMlPNuZxY/cSav
s5PTlRNTwCwbR82Cuqd5RvfM5+0DB2qljuzyo1dbDN2ah8MCoPTFWZYTPV+C3vMX
3Cp4HuRftbT+JiV2HcP7BWt4H7fscuwCzsfn0IJNAzpC1Dcqd7rH+t0P2wt/Fz18
cIddFbzEaOZ4DO2w22b3e7bu4CSTKFSNebOOwt4bJei0Jx3DYV98D2mOzdYQNa9l
9/PpFpjMngnrvtLQ7iyvW/zJHTGOQCuqCGT/VEQcQGzujK2TanxKG9aOCR85BWAX
d24sYbGriHxRnrrREtX7+0ptwJB2kzVVqw326KJam0bwxFOYVEqFpHdGjbunv986
pDzC3TMTjOYOue3b3QnANOXMSddRBopqqwMwEpi7GWAdaBMEHQmTBMXcHjd9kUkH
BpNT8ablvVe9+Mg9lO1mJVD2rWogqYLOZ8g7KqMYwEjTOwf7nG9Efc1j49zzj/1i
cLei8cZPFBoVgEwToK7fgriyGknlJFic9ewkCRd2CyPLud0HonxAJSyRwXXc4mcA
7wDjxoIEyhvZu/yluuP0MPQO1vCC2a13K4j1Db591keVD8E+wQNOUATiwefpq0QT
Zl9xL0Vpt3SQZS+K9094MOJNqAii6xtQy1/GSQWrI3K6Y7Ya1+p16HHNFpXN2W77
Hm8SYY8hALX426tEEnpSeHlmPZ9pE1s881lLXSpSlcipWzeXVqHRQP9sPptWCDDT
iRpm6gnTJzcG7SFo4alWxxcOKvstVNg2OAI1w1pgaxs8PXTL6fcMKgrMr8bi5XLP
FnvSDLCoW0Fi6G92imAwkgA6udZQhrR700lKc3IPzOOmXSl5HlKf1wYeoyNX7w/z
EwQt41KFfVsR74xaUtlW2YOA3pMUfqApat4pbk1qVLkB5cFQ0Kb5cPe2auU1Jypb
luyVHK+iJnFXvW/IWuSpfFS7vwFectnFunsYSZM/Ow5227SHPaWHYGyjsC/mnbqv
eyCCUg581iSFRRHDk6wx3kQkW82IC+WbnedEtcs02EiCZVkBMsRjdPoh8kFfeinh
OTtdrr52OqRpfXibBH91gwDvpXZMyJ5qD+CriHswEtC9OibjLfJXbDwNaNUe5jku
vVRM3MZ6LL7mMBtmueDfiYuzSgNvMTBXcsEEL0YduzPFgvqalZbe3hZTQjqOl/aE
TJ2zLRpKP8K1wuYf2HRLv6j8TEiKwJBNOU43UaWDOWdlyNaCA6IRa82uYf5jANQM
9KXd9O9+ESzaFtJWuR9Eo5U6bwDcOfXkEemGY/EimfixBMDMiKJXaJWWVcMQlbGt
baDkqFWjtOVTPxuR9yWc//lMfsKpeVM+KX9Cw77A1V8LU5lNHLnRorasSmn1XeJ3
c5y6qodK8X3o9iQMLIyBgierO8Ml/1lecdhiNRCoLzebkur5icsGldKDyxH5DiXQ
544UgKDf65mZH5MBod+SMH4MB4Rx1V5NLdnmhlhIvbw3WpPpt5F6RCQ1Lr/LOcdY
PpFy17/shV27rPaHf6n83gMAxoofD5VbKxvTrkswef3nJ9DJItoDgbiVm9szC95g
+L0gsy61ER6tRcvhNzVszDKHt4fFHGtLR4H6EsPA+/qPk+bjM1NWwEh2TnCfUAvL
kex58Cm02YReMpq7RXOV/l11yK/Jx/jr0ombDddxVhUPj6DrcUzBSiESrTd733ud
Z4e0cIyNlCJBXKIMWpv96Fq9mlXKmnqVWv3BtyzgmIIY3d8lHTAYEwN7UFxSFg3M
rPeku2fEzv7/t3Dpqo/wVAlsIhm1X0NT0bFHt02PHBL35Q45vZZu1oQnQtkNi8i3
KJ4PlQhY/gg7yN/zHXWxzpLRtwKYvL2Vq0HH3LXXUB+iLYx7x4MOX+FwHNahgyi7
vatninsXZj3uZc/JBDknQJLdeKsIwEcsz1fKk6CUsVYQ0xel+fQgxtAqFtqZ2vga
w4ZdW83AEZPjouPjj7MMoq462kykNfPRiR0M8kIni5TS8ELfhfATlehlN6zqHXIF
Hwd1E2IPaAfjkNHBCgcvPnhku77LESbqj3jZbLMcgyfP4/OTiJDuzJaUl2LeuHhG
CbF5h7FSKBEcREQ4iqVimaC89yY5ENPf6y91QiyK69RvOo9PMoIHGM2Giz3D44Rh
zqQ7NwKUR/pgZVq7GZDNousUnkEe7RYgyt0Gmpz12zS43VaGeNHkaiX0lp91230s
yHqNtnjNAdAqkNqqThaRW5VJOoTaf5IrRtZJ36wk6yRxr91UIMrXzSND4V1NY96R
iobJ7NUok+PyIMLETqcvdXik6yXsF+T/TBFqm9hmC/essjTKlDxX/7lKJi3gXgrX
y0GzuQnf28RGqCzYAuilRQp4gDijIQw+EKuppzxw06BWM0TUXORNIfY/P0NC8MTq
keQEIjtZ7wnW3+/pebOTD0rwoHxkC9+jkT48HzV/T3m9DlDxIw2xhs+Ay2b5/9Zr
KT3uNB1geGB5glxVarQUX5f/oXAg4+IccgOjDTcDh1EV11pEm0qbUOI6M1sAGgcO
l5IoGqG5vdeoJmb9PXP+mO5Hev6v6RIw79smFUT6FLjxJKBwsY+yIQw56nSjeYMW
oQZgq2+/xf+rq20Gmzp94o3Pb/ka8CGB+d1lQ/A8H2nBHS0Fq+XfCbGNcJfWEjBX
35Qy/fhnLO6Vn1jC65dCIY0bk6jMkTbXFBmToFbZjk/L1h1q3H6bJTWCPBTOF9hy
KgxCPi41ZYRqBnTD2ctCZwoa4ZbLe86XD6NcoOrDdQngve+tAJfiOIjxOMU5pEUr
rpG/UIBcks2gjxH9rNPON+p2lA0ui3G642HJS11lU5rTC4bI1OPXIs1OSA/NBgB4
MeUt2FiEeeytbbyIHINc9PO2P886xi5nYnffP1zN52KUnKx3ayRjV7dZOWpunpip
2nZp+F1vyLdHSsRVZ0H2nig2RQNM4MOvtPbASFoRgFujaOGSBUyC3Q+uxOVz3FSM
oejffxeugcynqbIrUg+b0pCEj1iOiTFa4ALhwayX/A3l10Iq1N9Bl8yImeN26+e8
f/ZKJTYivmhLyzlIJ6r9uxIxOoz83cO/h3TuBHMsdZ2R5drPE5FOrOzURGZXFc3Y
fQKpj/RutyMmV1hWfDD45BA4/TtUjjm5pRUY2o8ZMRvmiEPAdKgD9Y/4NP5IatRi
vTT0Q5Wnawg3/olUzYY9GRc/qhVYtoMMCOpRetMBVx3Orl9i/ZmAzJFhnol34Ksa
WhdekS9+lhGCt4ZqWpwmYkPol02jfAQ4bGnbVsgUqDA0GNAu6Xfuq4NgA2Z7mOdt
n8FqcSD9PDjrmdUTVU9JWyDbAQVXwNroGDF4kLMaWcSylCucxD5yw8S+TaA4NFfk
4fnO1erHruIHy15onYjZzwqMTnWlR4ZmdN/Gu3r10I0rIBqBb2QIRxPRzwuM+xNK
Ydouayqat7W2Tqrnh+c9yELusiSVkAWxoG71ryRIjhj1nZnspbJGfkBYtAB81Qb7
KE2PQhCBtylAw/5/zpi0655UkZwey4YkIiDrT+2++9YkK0bCdIRRQg1NzAFpGB+/
I9jgqWmTPwJYeUmsBNa3CXu8QvtbVxq8mb7YQv1DEqWC+MrP+TXlyTUpxdS3x5js
9i1JbaIGd88t7T9r30az9RqRUOfKRR+JUqn+AnpBhjyhb7GlqBPJdIl0GVK2lPW6
REnp/7CLQlz/KyES6a4YkCwQnmtsHBK1DcAkEXy438NuMP5fH3zqMHGjkKRIHPjY
f5fiWK7R6eNNcO9wnkqrl+WwWHiXvACve/DF+4O7zbQRvoGPNiAfX9mI9jBfB9g0
RHKWEcy2rhnxGUciKP6BiakxC+CPIXx5lKloLWAGtx/cujemI0AbDn2VC+QrsSop
KwqmOfruhc3kF7C+/OISYwWOgHTWc53in5uU9OzJ8/TL4WszEhV2gLzjbvuW4EdZ
Vst3FZfB7bzBUJmVEG6GhkJxHyD7QYc8NpNl3ZSyeKE81hzMK/XFRgWbMJve+w8h
Fbpg9eQYukRkf5Vvla03T+2GaCZuxSKlhyeCTfmOYspmprplOZtUMsZSfE2isW3z
lNrISiK3qv1+cX10PicB7gNhRDF6LeqBXCY8aioSotbgAzWQxG54c+QDgjNUfIPm
wkOicOLDm9opJn+gIiKGz3r1hZDHYdZIhtHRs7kgMzE748D1TEaXg/khVqUcH1sx
2c09y52dA/vfwtTj0oWyMvd9BT8OARoFpQGy9N2hwdj8n/0iFgADuyByHFJlQy13
bThGDHnpsf2IegvpN8O+3XqWXpg4UL8TlO5dO0/iuZNmi5biuS2ct6qtoCbsk6Lp
MlyOuvH8x1TjhqidgxX5qx4HFLJQO+Evu389f+YzRppr6Mq9rfJMZPfTMBHt4blz
RbBeBlEOaJdFeSDvuYdpYkmbVGt2xa2Q+ShEbOw5X8QsoMKKqYypFNaXx6g+phl+
Ckc+FTryJglYGu55eiZxVocHhvOB9U3lzCEWtArvzcfhGpRdw3+ixwIScDDALE4b
4o/rWsKDebaY4IywmqqBQMjNEUPRn0pOB+aNjJm8lIt/oL5I2vrconV1lQ/oSYUo
MTQza1A1F7RGGKPNdOo+a4fPhUkMkRwOBTm2esrtODz+O8kzh/tyy+iHFnarLKnZ
ytfwZKbreMhNxDSxsGGpWgVt8LXUtbdIVnzDpZ32yrF2G4ujFZuT9EBT+FrBEac3
zEKyByv5afwICqhv1MLuktZ/VaKTTyXDyYaNrYDNZBDQOLPP4NJEDjPu3Y2G5nXl
wWDW5VE30xSibQ7yAfsUmssAperbNLyuEEN53ECdA7UHC66KcbgGSdImOqnzf5kC
Iw/CsRpKzHi/KNZOCUrdZdUMPjmWedaGQte/7KOKk6QyhbPVsRo6gQ6MAW9mWA1o
AjjvYdSq3mEB1/vC6N7ceCwSCGpH9H9hJE/9jlDRjVCngZ3gfGnbOaL8mWuMhmzd
tbTqqXnw5BeTzttABHf+Vkg3JOpBrOQIXZtyNScogdzMGemseb2GLbvv1xNWoEaw
ombGqTfBv4FRRRvYpM8ZhjAfxrZUppzF1uNV9zps0HqC3VDwK3h9G6LGGs4gwGpf
p6fqfzEkfGXxVACedPVECr2TqRGf7pXgCy5FonFj/Suyit5yC43MMkXjHvMI+cOv
f4Bd3iUSk6H4URGMOv/rABokXIZPmxAKav24SOGQFOyCwLn94OJKZ3gjuk9+LM2M
pPHuq3hum37Mekq7kNf9VfYtOZEDvGzGk0+ZsjfPRN7igMPR0QwbvVrQDJNTsEoE
HKtrX5xX/8RMMYIKmozQaraMFaA+Qyx26HfQFlFJYaTNkQjRofsMbMFx/kYaWXhC
8fpSDWWnB36yWGt8DiNWNdIRB8nNK4adPoVOfEISHX2WKJpGr++IG4ymlmFHnzw6
B0KeT4H3u0u+xhlpRa+El1BHvT4JH5Y6AEbtLpSpwYxSMBVReDx3tfhOi9hm4nxD
bwRKb3UDsaDIPCVX0tty4k1+PfOp4XGwnN7IaPNU5ti+CqAZXd9x064aawSTZZsy
5lpyqs4SVh/TT8u+LdE4aAPQ0gY+LoAO71ng7cPczMLyPgrXOFqEhuNzX8phAXkR
hpxq2Et8/4Xn5UVUGD4ZaLWPTslD7oplyPvHl/tujUfB14yzDt+xTm4YnCj6/NnT
uVgaWlF1JpvodJAhnl36oSoymxKEm+NfyvYg1GuasThDSaEBfyTkXve0sV4f4qKS
bf2hvAvkp+HGxz3F7396FqVxMMa/96IEkEPhpRPLFyy9TDERufGljmRlr1Ljf7UD
ZzuydTkzTW0+nhJlX/Dn2lHuISGKa6TsPduhlioPNnZY6+InF6lOUl+/CDt+eih7
x7FjHhH+JBiYddQ+zTHyIUwRfcK5zH0C+DeY9HyCzG5g3SSX9z4V8ERy+TEhvDEK
sUCKqCukx+/evAeP1FBznTTQfK6KE6x5Z+aWVgJXmrmho+6ZIo7fHSUJWJyxVm9v
bRljGViOu66yMOnOXLBhGDz7rmZs8BBxeJ2F5zjHZAiDqSjHCHaorqw9CqF5GrN5
/xrYURXapX09cSwaEedHMbjctqUmN1oRo5ZRZU8Ak2pHBl3Mw2apLH8eDRhrAF9T
2xDaWoCrisj4AjkK6P1jDaYhdHCb494ruyA1esdrvUParhiEeIzhs9LqEekiIM00
My2dwYKPGLlXdOsFI9syaZKnYaOfiD19BJJd3t3MlzegQp90AxYxwd7xpL/Ujqn9
nVrfKBgvMttjCXM+mofOzhl6Z0JvRrDPGTQvPBlLVJTHfE4vHnkhOeuwh741tJQo
Ev8xypPAWOL8QX0hTjmn/H2/ixBs9lOCYNgrMebKour9WYKIOxUjzlCDOoYeJjRL
nuLxZKtstY+SfxseRXerlxRBjoZa8A/QIUTpEEm9br0ogJeKYpRIe2LHATmHzZWU
DQUHNqhytcKULj3VVSNFqot11ewDOchr9a/ilKY/4WdasPcwf0RrtKW6vsIyw4yp
Nyu/Sv/OBFWPmEOKZSpoU6rHqJJe2CFMgYEubkPUsTFAuFDL5Bvom/eC8sftcqLp
1Y7nh4ke2HPgK8rEGDP+zONtrnWAZpHpATV0dQIPxlwDq0IVdG7UqVlqbrQv8R30
6ZaeyH7mM3KJmxQwovSShtiYG+jgSu+dWUkU5eCqHghi+Pe58aZdcm0ZPvyAcQCV
/lwF2A7JlJbHs+z3DdTUlXP9/L1DZPdQXnbONnq8AcMsafpE1tBOf+ZF+3NWVK31
JKmpfmHxMP8JZ3jqvqA+cBV8YpgUJVCPHVbwzJTA1WqjAF7+lKBEw+gYabaL1dGO
NSipJ8D+ax2+0ggfuyDClRmdEq+3lNbeVtgReUiAtPLs3Fl/NvgdbbkqxdjHI/Pp
ghuWyNVCHeSw2HUJTiY88bFq2uxw7bUzqeu3paQqYChwfQ1nORmxIISWRWZ9hIdu
rfLQ0SdJEBVLsbiUOTDhEGt6IZFAhtN1OlXj2qlIq8wCNXTkUxUOE/s2kIkIaZ7S
rtyEqpc1jTCkOpQb3zZ+6dqIEbeByIWPmSxslmOONdhSYJCpD4Nlqu5CFTwIMeXD
ZA1xwZbeogjNtQFoRy9lSucmwrvSK30JLLVypu3TSMret9Bsd6C/+Z36WCd9C8Im
kzrkQJ3dtcsJO2Sjrdi7ZcVCK70ekWnlBuTYZwRJ7IlG8giDLxnMRZkzpe36v4Du
rufZMNA5BpWo836bjnzn3takh0A+bT4GT7Xrq4mIsrlbLfWBuWzD2QdLnkDQ9nDh
RY5A26YYMEtk6MiN6DQ559QIuu3mwxhxEe14KjAlPUo/SIFzH6Zw0/TmSEffY6Zm
SPiAcfIvvt13C0qP7dfHVPV5WxcaDdDPAanc7eHrxIaYfF6lRjMMt9GRHbuOBESK
hx19Y9EQe9cCVtXEYWvyV7Bl/S9L/qz04KG9t+hPnlNdO9o9qJ9L+yu5Y2Xo7j2z
To0+S30HW3GwctGoWWn7dN85EyoBaISuxgXetQOsIl++L7DFW2CoYCh+PHUAjOUL
U4E8zT+4iEnN2nO9fTAo7jo6dPtsxWR5OYSWUZVNzSEmgo9xBi/NMGcVVnLDKn0c
C5wC1NfrHwHnaaT9jMKHxkRCFS7QrOxBvNliFA79yPgJbcPTd1//Be03pPiE/U24
bX7KRPgrPkdKMytZN4Ccpfmh9X5vehKmN1q2W/E/2moZEoyDRrIkLdA2Ln9VKPSs
geMIdkgxQhXVzMcHxfr0ZKu1Dmc2DAqy3ytw0hmbLmyFybZDjWsXzNM6b3uAjcM+
Rqdjng6AdEZt5mkwYRxgA4ZUziklpAQWp8NhuuxVjEIUqzZYf7GUQ5mI+NMKsGBc
1p9kIpGLn4Fv4OI9jZg78A1fMjvqZnxKvyov+EckppqGi+CnPUHBFAzaSFJGekbh
wwB5bu9hp/4DYpx5b89OR2HI8J8+AeB86XxtIeaduBTk9aBAalasM9RvGexMbJOG
pgK+auE8ecANxQeQVXq6MWoqZBB30dMchjvimDSFuXi3JLDqUluk8n6iYqcln8WH
+4I4UKIYekKdO4E/hKjY33NK5k/T+NVwuJKxD6vP8KBPqhOFZ7VWaupKv/r5WzrM
deBg8mkbsqVMk9eNSm/QMRCxYWtBoqSAFkl8JjfaLYADhXG83G3+Hs4RDzBxQKLi
HASosAeyitN1h7PHEDrB4iafrivp68wRKSoeHUl0zzM/qzuD2GuEeIO6i7rYqIWv
mFcbPfK56igeFonOPRtPx5D9hjBHRnYeTPUAMM9SL3TIIFOyk0IoCiOBXeAdX3lX
Gt0ZPc0yMRkvRwl89nrgdLEEO6NYD1MBxPOhhnPXXs+JN/U/SNXO6epY4StAQtRe
EMfd/qPbqQm7R9m6Db7yFBTPgO4v7eHbP4osGpJGjoDj52wPAjOrf2eObenYXx+d
t/5wz8rwk8qEnfB3zJDOW2+fnFGaYJWlnzFlYQll/fA0TKGfrVVXXlLb6/QzP3Ol
o2Dyut2VKKTA+9+HId1XAICVKzWO+6iHXuwin9n/L+shlbUj2A6c344C91bOVJd6
Y9VagRL3O4r3eL33go7Urm3rVZfEV9cV/5MTiGDMC5ek8t/MR0SRNxYoxKlYf3Ow
iFfVKBLwHOrdvUEpIpzMAKhrSpgd35tMa4Nf/suidAFWLw5EyQgw1g8S1JWKfQ4O
gn8GojVRBU8s5drbn09W30934h/oOqLJfRyUtbfu99gozx7QQZF3Z3A76WW9z48G
cuQ1hi0LkFNN7kuOB+2VVPjHpFLbHwmTgpOxtgtuUp+FkQXiYoX3T9kD1niwh/bK
6GIHRV36rYK60JRxKDs3m8CzLjEZuWDC9/eGibBmPrSxtuB28WDUUWTIUUfHyNB1
mSnfmrwaJNYJQW/SMrPMs9kkKUeYVf6BEgdYUTFkpepdJf/tV1ExuFeUHzYJ+NHR
BxOKBS643Ff7bfce+Uz2qU+aHxyCaZm2WNWGCcc6TIbnP/PohZkMC4J0tctf9gWv
SwKRGnaCtEei+IJVOVte2Ik88wsi+3mIXdb/82ntMrvdpQOI0uDsatIjKITND/Sn
ZjCFMcOZDhALAu7hhtUE/tupYbWt+kG4iTM7IW20Don4BZFOWiERdXzky3sr7lrl
ST1hvODletBJgBbnPJI7JwhPIiD8fF5XarypnDNx5fI/4mxdyNecw9qZQpHzVPGY
mjp56xI9B0rz9QDSq/5wRyZRvZ3a+l8AtXwPpmrHnR3j5mHx0HeaJslWv0CqpjyJ
IaPUu0Da5Jg+DRgAmQ9mapYg2Li/ItHgccwSrFNrhisPCa7/1Z44deXI5wh66kfR
BsizvEXtFiyF/9RRHlF/r1fl2nlE1XQ66AKXbaV4jbO/45AjhyhOklfCtXRmZsEp
7IFg6cajY5cNYujgXc78ZGG8AGZhwpqO9HPR0uHkDGI6TPuih6r5YXAognIbjmop
nuHCZCCfwrgFocgMc1zUHO8T+3TE/NIDM96HYAQpAPl5GgEFCdi01cwkSvLdK2kz
wFXXfr6CQ9BWTZpHxvTv4tpbN3k5S8j3ahU7a3VZddyzDGUZiInK+9vODNILp0aU
Amfx8rErllJq/iwE+NgpxNhqH2weVl4JMgV751XoDWHIMYTqq1UczWFL4zyb5Ugg
xIZe3yXSFWJa4qp+0RhubgIVFFbrTUXoZGOhbOU9pfNJqH16MhVezbAoAVQkosl4
SE1ZLzkoRtpz7L2dBKpJXcH5OcgcCNxqqogXZgpUC6WsfBc2px91oYh/VQUd6Wh0
o/WVVJjxRaCTjcwp88EYuDAxn2S9p1MCS8RzxoI6388HdKXzLi77473M8p+Eq3/h
SWHtaRBqIgntP6VYCzOHxPyR0/VecS2ZcMZM3FTuicGPAiVMStIolK/ebzHB/S67
t2jSHymj205YKq+ik/A8DdFRPmcE7CjQnXNz8K+dvrSQ/ASoESq3D3taz4EP9DOG
ahHZ+2fhuxahhd4D46jdRvNn/gLvH4qU7Vs9IBaq/cLu/x3TMC8rDu/NjWmI2BE/
xOsckiB/ZtPZvL77k9c/bx7S9Ue9Nw7KzjCC6IyU6QUqoPBvTHQ0/hQON63PboaE
D2PItGqj/G//+CxV4c+Ocs7c6D0GR3lwbLqhsvD/1edCBD3UbBWIL8+jkbyS+Y40
2GJEfKUVXI9HEQBQeLcXgvovhkIjabnUKB6kow5o7jBgDn2cM0c8vIc95iA7YMsl
jWvcxA6eTw1O0aT7s55vkuBHC+MYlh//FbW0rxQar1j9tTxdX7P/UrdrPrJGpph5
/1/Cx3c1N3PiJENgGqklvUHDJbwY+ufVfb57vNJr/nommck1IxsT+5li4r1AZ5SL
vzoIbReN1dhEtk2i9YWw1+TcUEq95UY0b1EeyLeA5AMcuFR7VDo61GPQej1G9WKt
l1nKnHL90j2fVkLQfdIlTCDbgI9paGb+MsFrQ212l6DDH/9FrXjjzuDwPzap1KT4
VDWzSX0Iv3anK4D7mcCMrhCUNbqK/FBjCJGIQyEJ+Zz4zTb+ZW9M2oHwKlPD8rI8
2Rru2QUZxEr+cJaMKAvn3G9gTjr0QJbt1wDLWcBFGwOUZwH9fY5QGjrsmHy+x4Fl
BQJeEFOZzt6TW3lKHI4ircDoCus6W8VpJoGtW8X1pP345fSj+ott2dOVwjPl4QEL
idHKSo+jEEaiMRAfy42hSKyrrTDX2seM0pPMOBPX7J4azrdZFDF4EO4slSCWmAdz
krMefZZFwYGiTuHgalkdA6RrNyrWfHsCL4ncoFKo91ptxI13r9xAPE7lEo8HsFGN
IDxRH9ZCO2XmOox1njCoWyL0j7lUKngWDD48bQsQ74A94PrZcdJ45k3rOYn+etr/
/QjhBXVeYeBdA5Rwz3qH09iaCmpBQPBIbMqA6ZB+sF3SWcYnM9911ie0EjNDW5kw
JEvrSkqL6z7DrtkmAkEIQoEDdkBsCjMugE5aXE5yfec5c1jlmSjYD4rFDkrnTVOo
tZ6HPQBonCrF3spf1+ObD17H6no/l6305VLHzGhK1pPHBYFclt3qUYoPXavrrhlD
o7e2RZj770KAqsIm7ZQvTf2V9JFs8JBLBjXzNqMI/z8yf9ghZn4lCr9SO8agd0NJ
JU0RCeZXWZYyXQLk+wUXgvsDcrINfynJQ4KkUKpzMFCJVEncNcwMe0Cq0zFoF4LZ
Dxmhhg+YWSGxoGYfrwFR8DtIu3Pzt353M/fO3YYuFKJ+8gelZq/T+9a7Gj8USFss
2KMDQbUldg9Ixqto6ryCxWnEF4NvS15M2e3OMBZpYJS3ypK9ra6uM8jzGbcPTq2e
FfYlAKFFdpi1CaB4Bp2w83GAKnJi1In3kCMjdtGTHVv832v0Nt29cgWWts0jsWef
vvoFMIIupE+DGY/MsDYqLFXqO0wznRm8HuCdE5f4T9iFzH0P+SSGSXIxWcH8/09K
aa3bWvh6rNCkXpQIATHrYjsHvZpm4V2fcyKyiFlOH+dayLpOS5upKYiLFh2dbMLL
wnzEZFoAe9wXH2LKmXoN1iknlKh8uJWj5Rn9UCU3/2OhbwBSo1+9rF+/36PBMHWB
d09Wm98MNCtOLtNe1nsiebj6xNju0pZcWN5KZQKA58lOGMFCP+3F74OKwt6sCE5D
LoRmvtHMyOrKCsAbq3Ovbz/P3Mn1V/n70bb+q/qAtbwRO9LXJs4WcLqGRbgr/P/P
N5ieiFu8I1eKO2gdzJwW3VTwQNpzE9bcKhm60sjBHv2MvVVNjFLxJv6+i1GPQdSi
Un72JxzG/s4DxCaERm11MC5NX2VfVasEto8tnvVMRlWCFwrNPh5n/ZMcp+7LWaqQ
4kFwij7iq8+pxNVChH0/NTIH/6NMn/wOgbfvGoYqpQ/dF7szaFBX8rM0c6xAXV6J
ReByGtnvnKmju5bY7rHKJKneaouHQd4ySDDM2GFPVktrt15O69egjIQKevGNmrf/
I0yZxhjuBYxJdOhIp50qWGgRyXZmymsl/vSEK6Sz7q19nfbcbpuelqU7Fk7IxnTW
Shs1WbFBi3MWGiVeP3tX3hiZ+IHWEdrNCrjswHa4zwQZtJddqr0xgjJSkWYur991
2N+5tcdxRwD3i1B6VoAl1y/GEREVmiVrLYhqInSQ1Dd2z4OTPi0atqY9zYTWiZNT
AaYTxRP8l45oG34UVRTwal81I69DkGS3wkHFyGPjGjDpiwgoVmeA88hTMrrBGeaU
2GM2e/ehb9aUAz3U1iWKQ64QqRmZB+YpWwPN7/5jZt0yrOzIrl8Si6fLhrRrmORO
agU0vSk13Sim7308EMn87iGb2jBfaTX2G57wd55IO54xpIguCsYo6rPwSHfctZ0I
kAtA0QxphbjXQTRoRXZhNPoPV6wlB1yQDi9oTW1gJxLtNjBMMC7Qxepis9UsSrDv
CYLhQFfAQ8o+1r9500ljoIyQAi5JtPVl1rsd8zSrOlQIgfQp9c+xo9X3ygzMs1Gm
RSFiObbovbmbne9K3Woaua45A4MGX8U7T3I62M7Lpp1vpPYvU+qjVFq5/Ej2VJog
oKlrDr0a9aB8MeFQnx2yeaBDcMbVZohfF4kv4suo1inL1jy67EIeLtXDkXUlLhpY
qIhZ8osVh9M2QQ4dmXZt5qfw1IIhhA0Ij5oXDXFdHghxkFbC/IDqb9Lz53ZGsm4C
W3FdJoNUrdIpkRETGhuFU/hG2VIUAPu6ejP3ipy47leBcsXBk1CZAMtmhlJFu5Rx
EOj5w8FSb6UdVSlRajBmicm98gaI81Eg3uHj4+TBG7k0m+WdMOyzTCz/U5obJbH/
y57A0RVqjk43NIAqicCd1HosRROowyaO6HGRPLaFFv3tAgdUzMFXxw5hQd1/uM5E
qiTxPYY1r9U20Ot9RzIg+jPHoBbMWYlAilfZZqYrcL8BLhG5SN3cDEpjXxxDRvO9
ajAMsVey6joDaVK3rnDdzyPM4f3PD5aZ6587C7AncP0toTjj7qsXH9qmvIAhzF5L
EIW9snB/F0ebqd3l49vPXoigMRyaiJy1s3jVqXjCRTF9PKlJta3DTxPPQcqWTaxV
dEJfSjH00vAYGBgxltta9hSFh9gkJeTcbBlt97P2pe3FSXfvvdO4JaYA5uZ+cxYF
AAncZxKW5uNpL0Qdoj3sevwe95knp3cWK18sQhx0zdFaBz+8kDembLBnaoj1ZNxt
reXegVAZNJQ5feAzrgdX4mOUoKimdtk0099e2JH7A4+oV89Kq+4CMjNRd4iFuoKn
/gN2gHQx+lzlPjZbvbdD4GHtFlb/DeuFa3QLViLbmDT8DKrGAQQRfqUmxEj/gbVJ
DL1/3IS+Ab4EegKbzlX4DmAaZrZWH0CX+SU/zT6YUfvixoZwCZktqCVsPm9ZuuLv
9jcR5l2sv5iBRYnG2bFsAXZhi8zOZ6Ce+psYhFRUxQhaNAO22ZzEN21fPZA3FCLL
DS+1FVBKkJn9bsqJdksPiMgQZLf404rloQQ77MFOpKnEZ/LIYYwMtuIXC+s3AICj
3wvOz76ilpAsjyJo6JsJHzD+o/VYFghlW7Dp2ipCswSVFP8jby2wTUzgwcJ7wVYI
23nq22KR6Af7AJP+8sVmEDv0fLmnqr7fUtSpuTrND9r3VGmEyqlp4BhYD5aZkch8
6+pwdAugRaOBI/5OuMuMxtnpYz7+35AH8nBq1OcTgiFx5TB2ZHxgUIn0ncfLWBA+
uLd9akaoE90nLde3L8nBVJv/2Zsp7XTPb6WOA5Ny0H9VyirlRT8sPgv8DGxA+uGY
1SXgGiUIzmRQKeat+NbAe2DVL+DaqZSrOCSNqIsSL4VdTsDvJ3q0kfTxNL/BThOo
XjsQqCex4ggPWDJfD/CeP+sp8dg85Qm/wfEeLEYNnC+/yENmnFPUF4/kwdWdD5dm
F4YBoMbTeAmA8wEKAfinhQhD19ZbtcPdlVXa3ElGsnAbP934SV1z4i5tZ6ByAiDg
o4YjjuOEiFSy265dHhjUIMiN/fCABD3aTfA6kxaxFprY+qUvxTnW3R9AKVdy0C1d
yL144xcRTq8uN4A+seG4TgWOVPVZuFRH681tACsQA51OSsoS4xkeVie4C1kqemT4
HGVW/9kJaOv3qdPl7qg9Tghu140fbNtHvya0YmgZ+HWzsYmPuyzXPLhcFx3L/dq4
gg2UI7NzDm8Rzy0SaoREsuVicQ8kusa9AVGRF2R8CjoHoNv2aAKycT3d34rmKOIf
z2Js688Ypgk3kOpthTOTb11s1wrD3HRdcZcQrHXiA7CkFDbhwhaZbPIi/MWe/cE5
Gdw4b0VejGarcsWNNlg6ojfdRncpD5oy4Mh5n94A9jtTHOmLar9/T2STPhDwZsRE
BCJ+i3xvvg+WTRbHphgKZRcpIs/pM7x/m9vXhaz/w2Gr4fQ/CiddV9qNPPfCmPgH
z7KrrLtbF18YMpWutr6tTHFyPiWpH29PxkSJX9AYD5MJ1Ld/N4+fhsR45FUDQTBe
Y881OBQcso0Us6vpPaAnECCjyo5Uigfx0LAPP/fmWRvNz9lcDwZ7nxDyDZkX922Q
af9TYKNbLxcz9gDctFIeFN1UWaJM05Hs9UZjnm5t38+5d2fdOFdL+ScE4Ctfydxl
S+qqzPIYVK9ze3SKN5H7oxh3XE80IUXgfWvECsf8ihmA1NxjFRQ0HV3FdPTeAqHK
4aa6ow6Om9tgZ86LYeEKG7U9A29IEN0vkaX+e9RkfqKOYNfpJw4RhxGgYCm0Ss0z
W3eCEAMZRQnsFnCt5034NS+FGZLwkTfKCiyyqXpDjLTo455snJoPoofaGbcc0E15
ifYoFQG1urlSaXj0QlpaQd8p8fVdzk+/VBrd+ObiEbY7C3punMNqIA2pLtz1rwLE
CJnhntMPOb0mMU21nFbjc091dPvd6CBaj7QiaeFhBipnQy2vysPM3wJOg63fu0Yl
ffhXpQwqdM2yE4xdL0tS/gdUG0UJ++DxBlZCLhnkjh8nxyo5/2IvQ3n4fE70sCW7
+M2qO9VAi37xUCFoZxZACauMEDDZmetXMQcm/MGMI4mV201cyanj8prgrCPLE8UZ
hGAoW0xLLqeMAK/7k+3M3YqLago/jEM6ZJM+0gwRsYBtsE+1o/rTAHGzDrG6/PCl
Yj95jkqRMsRGuhIJ/GHF+MoGTDw9PYeEvhTpg3i1CU73Xfi6zbmWegJ7Lbd2Q4LT
jJC+uwu7t0OK7ehffMcPn8vVpFHYFE/lRqtgX6At4tIVzaGw5grkUyYNsq97QK58
7Wi8V6A04j97P7AmI68MMNbhNbhpinRoCTYH+he00gcTE4BIs51BFBwIbSYQHedt
jcFcso8ImH9tZSRLV1BCNJJ3zBchqQho+wUy/mnb7RymNEizifA54a8DOcuCAOIZ
m/1iBKymA02dieTtbfbQpmHILmMMOC3DgJQ3d955Px1/UDKPidQiyv8MOb9XlJPm
j6QrXKfBItY2WTOJaeR6QM5By8vUBp5I2hcZkze+wPwmlktzDevu5XpPKgaEdqfE
WwBp5LbBR4+uK6lCDwZ1MFkK6cGgirpamJ7+ApDcScgodIyEDTZJSCjyvERgbUGT
gvjClH/lzhcy0IHe3P7gCv7P9co+lPyDakdhpzQNmn9PTg/W9gH++GGnFBJJyIBS
L9OPm6rwnZSJSpPbw4rybTuCky2UxucRLKnl0tucPFHqIEM8O3ApKUksVw3u/7Ff
GR/kc0neILrMOuZzI58qtZ7vdLlv1r27v+eZc9JfOIMIcxmum3shwiHUM9Psuf5X
2rxpVDzvKotjaYJGkRejDi2pDQ+Ry+WzzZJKCrdtgvxHlNkbcW5psx3hwiyu6bMA
h85I3IUdibsHsFdJqN2PhJOwhzWejz8+XPSU72xnjR6IweHi0NFv7Jep+p1hVSO8
yDX//IsbXBvwPV8SEpn+/DZzJSfPmgdwi888averIpPRuQAZ5dKSQ1t1+mcVXZek
viUA1xCBidHxepAHaQmSOwwsvVdpexIM+lGH1LH32zn2fehv2TMv2leeovsb2aYc
fcDbFGaWCvgcLTTTExlRB5coxFx7bnoH6hoRew6A79I22kwjWCMeU7KraPBA1g5K
Y7UXTg69MKR486CKeFRAQzPlDP/S/q88lAAzIfa4A7TdmZ1siEXVauEJAQdo0TQi
K3gzBA4P4RmD2v1VEfRnEDjGLKwq/FavKq6/sjaoa/N6n6aCOtDBiwRNUPnn/z8Z
I/242K8TwQCYaOIcNlmVdKXEkg22UNq0suPY4FiIb7IruogsUUIybSO2Ao0ATLpU
3s1isf9m6YORmYXYqFP9SkDjZ6Tgp/w5DVCLdvMRprm0oKuvrhGfTNyvZeBbpjBo
7kAsvs5/obnJ0WfJ/EIZ4d16Lsnh0yCywqsA1dHXWj9RgwWjZP27wQzFh8qwjAJe
2mQKW75XyfVfqMee4U7UMZVXnrgfFhchEF6YlnONOmIVIRfd8kL4RAiU27+2IbnO
DfcabP2/FzKmZVXV3PyTjtt+pD7PF8xwkJkYXyoiLjwjmmmi0NqDv0MYMBeKoHRC
VXdkoqpBJ1qvOypG5tuR3eJ6gQCviLjlDuLjC/V/cby4aQRWZu0yIXMTDpAKWFNs
NU1A6bmKzwsEXArSh8R7oq8iQk+1NceysPJgqKWXJFThkKgRk+2QByaJ7q+d/3ZN
TWjxCBCmHhPFSL7W6ylt5sI5caWVcAgN1pCAsrK3HbtBPQa7wkuOc8b7aVT0WuSa
TA7o8id7MEwluctHyKNMeU3TzmknvHx1uTU7ky7vW647PkKZGD9/ZLGd7gEUBmJU
u8RBnRgrQpzqCEMDqSTKJbM9C6LL3sTxkCqA2tTz3YVA8zYGNFANBI/RKMm8rq2n
MGWgOwZFZkx+pZUu22wiqSznd9nQrYnw02GJn/PaLMzfLlb8dIGe3/PL+cmZuokn
9ZULMAytMZr4aKb/btAI44sLPtbFuzxoPhQP0UMQJaSybpuHIMKKk5/xkxrpGK29
t3r3fPm1U3oLI6+FnOkkNWiqKoNQ2wSVvZyQMfxoZStAfKYmRRI5if/+eTH1Oc6x
Z37lXeOz131cQuEnjC52ranECnUBcx8gdXwdc76xPqq41QoMdRSbAAxO7GdHoNm7
5zmdMbqI2yzwshiLyhPBAmLqtCgfoh4NKftH2FPkvHEr5EffgE41Q0TlthReKVgp
vdj6DkohobojMR0JGgBlJcliqGXLGuZ0o+w8BvG4bryUMahg1MquESiXxcZ+PT7A
yn3pIplzAeXI0E3IShbh0y/MpXWjE7dPhhyudx6fAb3Z0qz8fMoRyopbiPw4VaKU
g+/oi3Q8JiXSA5b+D7w9Gp2DJIjzgUmiknGdwGMIXIk+xVsGV/4YpUHrcULmC5wL
QIATRIWvRB5RkRBKua3jrY3jAmLeZ6IWWDqzNZOBT4tjWOt/pUcDYpmMMSyX/lEG
axnxi/jdhENxR2efx4EFNiqhj2T/C7s9Mt6Blmu/Ogbxvvxl4TxDtLve106KGG2y
r8bdMEhKR5jrGlNd3+t5lBjZNuHpVHwxG/5StRgjkcR5Lb135VQgBUms+oQ8YhN9
ZhKZ+1gGYL+gzflcc8OqYY/Lg4kw/C/pcONoBbxBHFqtGOLo4l4/rzDI1tFYZVYV
Ky5bSYUHADQqMz1FBOyKbJkGSUY/mRBZna5faCmMyR7BCOeCR8oSM0wtrVMJvDSy
IXxSEoJNzg2hVjs764C6ZUT6O44edPBARRiJgsKaNPttyqbzjjff9zslt9Akc3NA
KZsnD+x7DuqcULDZMmj/3s9lsZA5cXkIKNocX0AAk1/a8hIhcDTohQEXOaHA6wha
jeLTTBZOpfpUhDhlvJO5XMAMSGcEZY3+9eujO5jBNM5kGgmrI9z+GOyhHKrvNYpp
ZDJXR91A4JSFhwKJwYSraE8YxyWnHsSg0+oKdAVMQX7mh0tQNSa2Bzot8veuHGD2
uv/U3nucKuV7O92mBCzBQxV9c4+jseR5ptaUbmRx1xlXfN+nkGnAeud1QVB91jme
J48JeXs8OHWfgWJLfCF185IQzNBYT11GC35tF68+bQY4RS5cHxfMFDNjhLodyPNR
EpQbdh4W/LU/3uVrXcX9QxlWQ+C9OUnqL+QYCgDBCQFbpNZSPN90Hw3wd0k10ezq
mj94ehEgrFznnp6P0LFzWvz40HxdEgR4LtDSfx3Lv9qqZKCeBf4vbORMPZrpyE6a
3cZtbmaDtFkqS2paT2NKR+bdnMrzukKNuU1AZ+Z3TPoIJgrAjjB+uvv9LbLyUth2
O/kJpFU7lqRSD1ziMuI5sQd2/SBT4QHZOA9yC7upqYf+9eyucHlDI5gV5xu6BJHA
HMVE/5w41GukDEszdQU0LZKHu6+QpLvooSPmXzusaOQoZ1YOI6BVf6YKNm9FoHU4
VwRLJ036rL2SxwB5qi0Lnmh5UwSkbskUl5crRSxh5+0IKGrHb5ZenprArSF/+rmn
EMz7Nq4LlujDtrYqZqTV9t+T7Yxi/F48Ed+R/CTJaZGByMXQhmwW2JF26dhr+Pvu
1JTxLuvUGm+O8nFXLYI6rITe51nnMaot3RTeaJoxin8+nLiz/1XXu1VbZssvr58Z
+SSZ6YXOYXrGcl3yGxCcE5K0hu4QdxuJsn/K9MDRt0EjdAjak5KoPuGp8xk+VDxW
2rs4zZweru9kQRMwHVQqyFv8tWMiNxlCEOaliEjH27ShkD8lXBsBU3MXASGaVDZ5
cJ0rROtA2dIOui35kxZoEPF2ezndOQWfgzW0pGm3KQc+o1hTqyg54a5CpL+M50k5
32HynXA8ZJ4EI+toMi97tzKm0uBQfgkabPYtN8tBqzRYIhKHr+xyqjs0VoeaglHR
nLQFkYwvIHFzVhSojSaSLRBvUkm44QNMAuuAB8L7gNbij49Yk+5hmXPUrpaSTqss
LeVq9XvJuqqpJCPyWsYPNp+5f1Zcy+4JpRQe3iI1z7WyjlSCZQol3fP3T1bvLpCh
IUp+fYKBWVb4TKr1yjLUZ/RMS+6ral3cXciqqCTmFM21w08GTLmfjmAeSu8wfXQ2
ihXyVypZXuNkQfe52yAWowXlZSSZahUYIJ6oZenuLYbIldnamW3bfEYbXPwamzK9
TollKg35loprsf836Y7BjFhLSLsTR+WwI2dMCAjjfFJlDWTv1z5O7Ri9B3oLkLPO
rsJqEPuMS5GH7adMp/tIs39Mf3zKYYZg3luv7Wnp/fvqdrrXhhKw7xX/kDxS9Uj0
uWAlAUyBEI++4u4JdxDK7qUeoGdZJRIhfHJvDVVxUzxKjYEPPePOGIvO+vMexr4X
9gyCF1dXP/VHM3ldwzPemvchyFKdl7b3V1l7ga7Bcmzf9yRtSOZchzC0HhBJz3Vi
KF4cGnvYrOAee//yZ+G7i6gZlxv6DjsVNdYFE/Aqxs1e20Es2lSq3IsHyspVYSwI
BLoxl+M56fQ24UfD0DDrFeTLP947tW+QGmvRKcl4c5TQOVBW9u6+rOusL7iwp44w
objnFmoNtUp8t3okj9nNn/9NVYLoVH8zljSsqtUUiA3tB6LdD04DsZl47GmnW8m2
dJofE9eQ2R3LlfE3f+b7FaUe45mzDIJgidbn8H4DvsohOenclCXiF5VRcVtkfR0Y
vJJauEhXxhHqUyOUb5L3uf6rOVqs7reblhqprZ7nY5pZXxyNOEQUFTonk4g1iy90
f3WT/mEtvmjMa1Qt64XZtRNlkcUqvPuW+qrYJL64xsSv9iGQ28TE55Lk8p5ODH0z
szaOz7UY4W7bkhmD5ylvjdUsQb0CzUOjuP3qkvDNs/0qMLriH7kSUP5jLZoRn2FO
Pki6eIKzlDP8SistS8uYJcT2pCL5yTFktz8TMjH2k3VqudPp4KOxOzZZn1TK1/Uf
Sher/dLFVWEu1PqpKWpKe7qfM+CFJid1HrbOlGyyhm5xRI+Slkg0Ja0NtHXU1u6l
GGfVpuoqkXquN6K6CRYc3tSnEa2tATynCKjBa24Ywh+PQz04lLkKKBOAR589nz4u
W8gXIgsN9kevUZ7E2/JMuxHplLcD8/gbPXObEl3mveSVk/96OBiOClrdMJR8U7Gc
L2+sNBXnatT1gxtYWW3NLDZkmiW0GS9152e5fkIoqqJVpeWgExalitah31lHJU4h
D/RDXTxwqOrInp2++Ho+rRVHhMsnsRSDWVjli49zy2fpN9+xcM35l6B5QIq4MXjT
JfS0CHdBUxsObY0Vx+ZCQTUnv5bMIPVt0oQGuxL9SZCrYzdMTNpfa21tQk82pPy3
r1dfNms+uDN8D0tAfzPU/vHHYqPsztcZVVqYvEoNqnQRIKyrmDiejr/dikjrD6HM
DnvDLTX3dWLbPgPZYALw3aLeWy4C8a7Ryft82F57OyZnb5q38PFLris5WqJ21bxV
HNxw78zUPm5VzsWDpWuT3EM2PvLIrXEjurD08S6lC1eaZfpF+AOYIrQojFjTkUU0
eYK3g3/RhoO8LBzpeUzXMvNZkezDF4dl5OD4E9z5fAF8qWwO9bhA7SxOAUEtgKEC
tLS5AIhxm6PmJWKV1iShHrehJqSBdGXHVpOPRrYtB09djDwuZuS+FejfPJVxNFES
6/x/6t7Kw67+4+RJft28aXN89V6aat8qzf/VUCAPR/UPGAUXbg9ZCjKa1Xyapq/k
WApJ4IP5peeNy4o4vs2yj8OCoB++4iSvF+T6me9arnHLErk2rSIoEtJRPh4uJ3Nm
fPIhNaAx1BnIK5gRB1FcS0d6HA8R0eq42ts9eLHK4nHdhy6cWYAopjlyMKgxdiRD
i8/PhIUTzz8IkWvZwhOzpfRonrGsdgKrcLOiD9IM3Za1dJqrfqfXSjqM74eza33y
JKfJMeQam+43oFpYM00Psf62LiQ/MKxRaJLVBUHStWKuKE9IzaPt2mAAz+/zWM9b
gL8OkUevkbKeG70tT8iCiVde+tz9cY8lnOtCfmWNBuC1Ww9XI6dpMowuffAAZMd/
5dt2cNqurGCmKWaL1jd/ay8cSATLX7apzDBivU1+/c1sF7XDj73EIi3VupjjCBQs
U4ZRsdcJi+plb0elzqylrmG7cCsReQA2EpxoPpOrhd3YfGOuJNncsKPSTstjb9Bo
32XWx6WJz7/Svky9lWXjS/xRID284f243jZ19ovZCZFsAaxhSAqdYi8lfvZLvI9h
DnRRainr0ynAz1XhFl2nGcIXj9ANhlzCALxtKeLC1C0XIuNYyj8eVEoQ9FYecpkO
OT1QDh7COGji9sF5MWHRNHfSytuB5ytE4WswlBTACKPeZIrNZNMBgmipw71aUxwC
HDr61f4L2yCLk5V8ytA1gh3h4GOWPzHzh6OOR8Hmc7kISJJM83Jev3zFX/U/jjLe
FwJHHWkxOKDXcZgo+6c6NTBB8hfY9h9VCYpuMSC79udWXrjCrGP8sdHq38C7Qupr
/iuXtb0K6G8ChNtL5a2l++fYxFURM8d5wy0vNgksfTDzMz2v63pCweg7uc1B1gai
2l6PFqSVJfPKSGs259hL+OR2ITrMBA8I1kH/+ZcqohU9x/cluIhYIRtXqW0vzTZy
4oQljVY9+DNoSThF2dqEgwot3ZFnGpBGNFzdBfmCtxEB5tJ/uzedx70g80nWpxkJ
3h2aa7gBoNhtrZB5CP9xl8GNEG4VW8qRTr/iPv6aryl5DbMhkSKaD8S+W/x8HjoJ
/CuczrYegxbBMl2JzoS0Idiai3400GyOmgPhmU0GjXIXg7HjzUBU2Lx29Tj5g1ut
8f74XGBDzonLUAgBy7hBpa1IiyZ1iTxlOn+5scweFuePOWMhIwUfCE8dDh+3iUda
z4chf+YjSZF3v5P26iBLTV0xwo4EzRwk+9zLyqu9iUDnYEUPIBCxkKoPX1P9iQ8H
8ShwbsVF/ONtUGEWHye+bnu05UufoXI1lR0HnOOWiSKfF7omyeUUDZzWd5KV9nbn
TO060w8EcSw2fNQChwIrnjoFvUfkZQCzQ7/lZQcfOpltWfRMuiooA8t7FH2jwazB
hMoVS8gVVpAfWEIOxIlLr0czlA4bysHfTgsjYc19MjgNAcZIIAFbh4khrwGI/lFC
aagP0C5NyA5sj9+jxJQEKtt9ZU9//qTvl741GbZiUWn96KAXCQ/+g38HSDVHdE26
1Sm/2T+6Gc+v4GWzGzNCKO/4cqFA16938Sjk+d8L8/u3x/26omTEgbvPt4l/48qn
0BcuOKCRPWSzz5eUKapu342o0oKUxCThLq9+1lydOZqaD/sjVBQtF0H3T0d791Y2
75vVP63Vfaj7eRKM3Lgx54usReal7LXN11Kk9eNW9AkCUEBAtZmS1aeJflWbWH1I
eGEOWwAuSIBJlfKJSaakbxuBcKlSj4jVtBRceNTUa+TUcvVammgns5eoREng4zNf
SWKofwnoAiKOEkkfEIAM+7xdW98J33aXNVPk1sMIp+XKnL/WeXVjVbHg4h3XMJLD
RdP2p45w1FFiCqzv4H+xBHTMwqEozZMAum/+DCR5e8HfbC77TBW8Mzg0z6DmXMS8
bV7IXeegqAs/b00fxOyCNSHizTg4lAbOuajEaayTxZK7eIIU3BA0Zp2IYzvlsTtB
RQ+bHCFTZKx3Oub9Ilb7j6GyHvYqlLyV756+NL/KyMNkMryK0b3SFUyUCu7CuJUg
+RiHpKzPOlZ2hgxLAuSefXgCepwfecBRRfXSMh5nbrEb1MUSllg7lQOnaZGQIf/5
iy6Rq7IBKX5LFXvozfuKQ/k5o3FfHObqwopthvlLhCTiVgdIBWm8iVKkmA2ra5p4
/n4APYZE/liflR7Te4FmCn7zyiz+KQ/awQCEuaYFJFoViE/qExwOWHjtM9GMojFl
4KeOnNooI3FR1gqaYleS/ubrMRvV7Z2Z6gRoB9gOKrV/T0n4AwiDJxEy8/nbw2+c
HAyKZX+u5kE0gc6I6QaTYa5PkhExh0EFe8UD1xfIX0qpAjH+a28gi8ik/bxvCwmm
TwTCchaB6nEZgKiRWG7UGRcPIhHBHGfIig1E+3/KhXVDlZnu7bYDqUqrYUha6uBR
OX5utBgIJNe6FuwGrlXqDiXVtj/oXZBgSBom+19t/5RwPP/2IjcLRi7B9illC/C4
BR9j50ThhbfXPDGHIcS0PS5YURTI1TPs55rrTLOVqwRhrMupZBtIu9HqmLZ0iW1A
fcuCSWT5vdB6BCoAMi6DmdvVa9yvUpf2uX1397FETI7poU6xj10/ZDcUXCoRq0AI
RjpEgErz3xc+EvI8/ipV88kZWJABzxa2JEzCGODlZPL/xgcZlbNkeP1hF4Az9oMJ
zrPHCruO+cuh1RfaxxA9piqxjGQVXh0NB7lW9y6VcBIGVeHXG2Jy8NxmYs7v7NcH
bmBxGpMQSY9j0pyq3/w//LBhCRLclxagBN09quusqesvGAqxqGunwXjkGz44g1bI
d4RWosW046mi7DHyRyrDWuDbsiTF8PQvgyNr5dFDxgtNLIRENLgZCYRi3xl4ZRm9
Vd/480ZPiXCQ1NVnTNb8UNpe5ImjF/sK+/yVFuECf1UdeLCsVyL8doYfWbqv0m+m
TFf3ymawZ3ThYDZ6UOJ2iXc5CLUksgBXjjZrOIA/CBy3sPSckpR7rYSsI3cKWx+W
6at3YGCk+3WoLkYErwflhngfyZ8R4iQ4ihy207NeSJHJRNLqSNymUFr52cwYGqZe
yUGql7cUO4XwioVtMoMcv99U9d8gs59UTBLFXm9ZdHK+Jn+tVcynKoKesrhoGqdV
47tlSBz4GD4eA+hZEbnGKOmP7YVUYC8DI34qjC/thkkxbwGwMDVaIJjK6P+rqp9x
AwAPpKTV4yXXRHLMV9cor2opMgUb58aVfSMEYUqJvrV6g7v2YFWuN89Io4IHADP3
8zfQb6bgsDkl8DxVoxhCwu42ojT7Fw5zQXd4PS+A52JpT+z4oaO+VEyLYUQwzwM6
vKt825xAoLamiZ+NeA5mpztNpNwYYOgFf2GlnxwrFaSEKSogdQKZSr0/moha0hCX
mvBsjIwSc+ckWYr0i9cI9bvjpJX7QJN8IMaBIGNoHqtqzAARlrm9fNwfd3C6g3aN
AQ9B9i+I15Fw+xOjpTSzTXURvnSb7gVCoFgvFk0oT7SimJDxIfj+WKEKHG4/kFZg
Pq8oznxCLdFYEVYy0QxgaGzPKRtCfVViK/Fx/VEWKa3r4+SfXwRoldUpCCXWCMt4
Lt3dBQPlIvMTt21nbQf8L7Q5CdBY1kmSL4QWiSGdKfkL95C17RHUyKu78+cz/C3q
Gy5Z83DsYgpmAAC/iK8F/IDKj0l6Xur8Xp6PnSm4D0Jf5chhh2KElCNbBDNe4KNt
epJ0dnIsN1Z4pkRiILLCba4cNXJg8Xx/5Xk1vFKGi7BklbWK+JAZLIspBRBGv+8x
JWb0EvIYyPLEktCMGqiz6IQ38ukB1Fwt6D0jbHieToOcyWtEh9CUXqxfluwc4V2p
zkuRbEJZcZJR153ewtFDFbbwhuKPTr/HDVLf9OL6VePPKP+h0gLPD8G3pK69Dmp9
jbfbTRYYI9wf3h0tECqQ8AVrRI/k47P6n7sTC2Oj1hpSWPSeSQ2VFvh2HMsWDmWN
CDXKE2BynFapyPxC2AaJ/vnNbup1Onxngv7Le1VE78e/C4I1Cb9uxpps6RZKhJqE
ARt6marcfzrZCsRkul2rZI1EiULngNmRvJfIenByedCmkGzi4T9xO16Q/flScbtP
IkwtsoZ5bFSzrOEry9bh8Ycwh9qRnJoO0iSNLrJp6+AkqE+usbCCLcrW1XT2vuG9
thFwy/6yxLElAAHnJYVyMjuq7acf8uFVzYHe7tH1Qy7OJ72PXHbTYb1SWFNAyqVr
y8Xke2XhyF66CvRCMw3sV2jjWanwm81B1D9h98eto261cjlZAi/gZzLEHc4wuhQQ
ixWfNKTqK/qAKk0coViNetvIL5b20smaZBJ599OMvZbCKODMuTOiKRdojVagIoO5
BolZMlcSlDSRptSSLkSh2Dx0LgfG2tOhW2zYk1fKDL1rOK/YDOqHXDcwR3sB2GGg
EuNvwJwW+f47EDY3c2F9nHDjSknw7VReSrYuSVob+FdO5UCUJON1scUk31yt1R7k
/k/7zzP2VNTcKYlgf1bvg/34R8ZSRCC4mGKDl8MzP6ncXACph+C4Yq6s8VrwvCBj
/54Pukd2Y98W2B6dHRwcbi4wY13BqwhL4sOv1xtNRua0hOe1AIaPX3HShEWPUIWe
Kl3u3XJSgjceErmQSjCmbLy9kCI0pGDYYj7zlX2EqgZ697SmY6p/x1U5XwFWN64Q
VulFQmDHn+VL8Cv6aEWq+L8f6PU81ogbnD+79vDCwtD8ZS1tesqVptLJILn+PA+i
o8wg6hmpgzLfnP2aRkrzwz5rEIChyZuNp9qPuEpudGUep0bDi3kb+5Wp+B2+Z+Ab
ZtNr26qfbWnhmSeRHkC03jU2B52nmPjV7j0D3Zs07kpa15FTejVzRmwlUrheyC/3
VRLujoUk+p14pHHtFl03tRrhY9PmrKT5dTruuBtGrcRSuZCQ/MSHZDD+l88WnrMS
XMxWSIf9kLBs7hOFFPVvAmBAFjqcMGRod5aw+XVaeytTPffsI99V5X8YPjNbpz9P
InxkGcHyOwy2nBgI2TUNXCl6a38c6JwFBwuCJaSPrlDQAyZ9cBhtuypnauYhA+r5
VaQ93zg8TxUgDLCg1G6LWE7pvOPaUenzENlbYuYD/UeWTtfz4jvDOHUk4/jTGKyb
foD1+z2LnHA/7NuHHctcgFdX46rutYfxxhvnqRg+x/uHzsiVvEhNZMPhYPGpvwy3
VEmGoIgVcQOscp5SP3p/rZkF+kDs/ecko6LNtOEhy4CwKDZQTz2k9eLBUhmY9Ot7
r18HA4F+rdlkmT1EVUjG/w2RWJflS5JaES09Cx0fEsxxUanV/gEUbj30E9oL45jv
ShNTVDkC3CWqFoTfX3lEhd1LTW9dj5IIiBOV2+YCCMI5jBwHsT5HLxrRpwBXfviz
+HsunQvGqzH1XMUhQZknQn0KPmTUi412s0DHwGzWZCgLBcLjVdM/4Ipl12kcHskL
w3shU0xIBEeupnIkY7qW3nBrhjI8TgVFyNAlBmfle1QbjXLZCO0yN/qKPAVM7Al+
7RK79Pb5DGlfElBbiHvN2EKQU8V2tClN0vIrRwHR2oXXveA7mTd6p7PB9mWveLX2
f52eJ67RAHiEDt+r5ZxnOXAbb/UOgVDzPpGU4kQgQvRlnzgwv8562QF1bfa7WtKK
mhfzgH6vxb9i/ynfaZTZLgJ9X0ks77g2QfXK8QWmegugvEsrOJJmQIL8lAyH/fAJ
ZK8L3ULHVBcT5qvm0OQEy38AnPjJYqTsWb/hFvQTbLzYoBfxox8xlwH+gOa4iP7X
ASfjakoOEcHGLLNKqmeVzH3aO41JHUCYqemo9i/hhppU8Zxp49FiaVlsuc4d/t/Q
OjZMhDVTW1puiaadQGFyOD/BPQX4P/LD+Pa12u4uw6x6joMZQ6M9kbgFx2Cfn0IA
8ksI+PNu/jaTeU58nGjJGI+pI0GvBUHkCNFJ55Cf2A3lWoKkvPgcyv3yfnswcfIv
89PHSLzbWCAJ1wNjL31sylVmE2Hh+QR8k7IOkkz0bOazeS6rWW43I9IDYFDN3WZQ
v3keAf/RH9R7xZXtinPv+kBMIW3Q+62o6f2chu1maZQ4lFK9NJ8T6unKwlAL4vPO
d56+qqC2+2/mPLlCGb8EexXIdU/z1gVSNID1vcwVMf2az12Bf5F5Jag182nEPcge
CzxjTzjw3Kc+EDWye200UG0SWDv3uouB5Rm/ZfKd62NhS6CQk7F/b3fuFogzpkhf
N6ts9+WeCdNj7M/BRQ8ZMm7NHHTvXISI6TXoDLcDhnJHlbsVGJB8HnyWzdrtJVR1
m5gbXnjoxfEAdI9Lt/WZUEGZNB0gWDP1vyhXy8/PULzmM4TwdeNW0uSSJI0NsBj3
3hkXE/A6kU/nsyuWxLSCdGsZjfwHa2lhDD16s52/6OXRvLy14L8RN2ehYjPybkak
i4nBrfKXaOuMjuQoHX+T8gRupEgdombrYqzeLvrTMWUqUmqzocNiwzHp4pB2kqWL
9CXx/bHRNO4c6hz7v3SwG4it2P4JK0uxYMOtM4deuwMoN7Klx5btwnyUTmLdK8sv
ILh8N2CpyWdqUZGEmSmArMrpAk/O7aLYn55qS/ALfNGEbPY4bolx9b/kGkKWKB7+
k8xVNp4io5JWzrsf7XViFiqzj5odpZuRMihCZkythZU2JjfeHClp9f7bVQD7/pfT
bbPWcpTW6bAvHW/dVd0e/Y+C4ft+XOwGfyHdKoChl7kEc+DnQ/yHyLvdYZtC0H42
GLEFYonM1JaN0iyxPeO7MPM7gfZ1k1t+aEXjcD4VucKLkWOr0i6DvKIHukYElWPW
niqM8rizz34gMFVaSXi/D9+Xw3sagyqpXtQeHLCmvoz8jYBD30qwpCihLpIYuKb9
bl9gXeKS34jowaYItJgeWNPrSVDwPHnbWHALWrTBLQsOA4/P4ektKsX1in44QKM/
sdrv8InlczYfKf3OF/Bth7qUDhrBP+CKDmmVqpY/Ic2d6PrXR4dWQDnE+5c8/0N1
86U1uxgF4jZdra2ojUitui+b0pjbm8zIoOcThsAQVoQmqwRRNMR2H12kfNbrlT3/
7Mb0doKt6DJcvyNNqHuGXy5uYRPvxR4dfBdQz+hYbgB6gPSSzvBSjEN/7SIgt2tW
ArUJ8UcklLVueDz6qXjeMCValEUIvSqFh4qb+GF3MLA2Vu4PEQq/OlU4Y27zzNrO
JWE+/+RS6HqKqP/g3dkoY4uPwPtVwGd29CH24ZCVxRB+m/snE8cBD3yrf3GcviZr
gjtKezgk8CSNT9y22Rum73CrTzR0PBBQsJ3Q720Btzv+SamC7X0ksCivGcMVTXXx
4fM/9vJb5Jjyuq7ZIY/BwtEF/QMx17QjTRoMQHWe7a2aUNofuJGv+LmDzvvgWywG
H7YBTjwMGymirbnOheSNO4FRacVv/0MmVrEevfjD9IDjCZ9t9lP8TPHni7Uzsghj
sAOqOqPhTyEJlYERyWOR+raGAW8GK+jr7SYa7Od9Sg49wa1Z1/NUvnPHveTwhfXf
NpdFD1+ebJ4vPCSXrKGUHr8i68zX4LqK/zeFbatMcLgag7rNVgZurOQt9mNS233+
m8QcUGO9yraosZXkyoZ6gWB8NtSX/q1wTOOzUj7HFl8PNzvtFyQqDH3+UHMC3Pj5
fZrszLsUYhrnnST5nHF5RQWdygWnIi0cOxWOND/BBu7mshnpwz0QNSl1HNmHHO0u
HCf521raxkqh+t9+qMFOCDXZGog7AHeYYz2dNhQ5vPT/dzju9HSzNPJXS3wNiU+y
GwSuJnZULFjJWAmlqB4KCV7mlGMF9qlC894s5JFjY1EEOXOSJ8NiEygd3LwWJiF5
chlvuXwDps5dl367P4+V7WFIupfl1gquKZMd6/Tfnqmnt8wFkDtc0uMQLrLSmZPD
KZilT7kZa2H752+wGlV7NNQuHkk/cUrJpR0zr1yBcQ3sVYxkCc1KB2nW1pwzesde
3lOXndkCCvTWR+WK8fAklrtz62W72t7RY+EZWkjwiT4MBi+/tBKdriwQw29Se1Jm
RrbNT93nnPzucz1I/cGMFaOXmpPVjMggCaFYG5tw1xLWnp+ytnhn21EVGot8WE7b
pZSVqr6tiDN0vmKeOYUAwdbppAQnSFlagJ9ir0Sxi3IrVapK9GLzZmuKwuvwuXcZ
IThg3qUAzTrODazmQbow7Um7LYhw0MT6ZsU4UmZEzrWc2tRURlAc8B4bzSJ9nB13
bG3u4hmZCaQoFt7lwc8xf7nOTU5F27kfw8rPR+8u2rEim2XZZH/KH6XO50T6prck
kcbCuqqHSiME1g+0t1mkfhYxC3IK4t9wqY4/ddFVauRzvXnUOatxbDWam9O4e3G9
v0VKQDnAZTuO4vG+Wr3A07Bl6fdG0f8vnsmjnuzcOLmIcVbNcg8n4RY113xck7U5
IWhL06aISrdFCOlzg9YJ0LvXZ1VLRKK8/acnxXPmfA9aPcVqzE5025HZOJb7a+Xb
TE16ZKmAnjjij4gnd99ve3rnP2FUAus+rV78pB+A3Y2OdarO5pWLVB2upWDptNUc
0U4+taz15a2CafX/Q//VEOy5vCO3v3zUuEWEInWlTrjl8R/AvBBipEm70ecOPFFN
CfKGgCKE0Hh54aFSBXSNeTJ7a/ZUbbAmpyhvlJ+ENTrnt6/58OwGPfqcdMVau91k
EIoL8QF79EYFrkpWo0ydJfG+fiKQhDbtKFTK5WgmwGWaXPIMCO0nOY7dcI4dvhH9
Pun9vgbhsUEHgapSNlj4AIeNbgBZLYJZqYbnzDzaR6suF0r1N4e9pJgofL0r1DJ9
tT7G9W3c//kIgwYEqUvZcljnZwYAPUMzari5cxkkTDjRkj5cZ3GZsJvE+DuHZpXa
VxePWGA7UuB49071/sg6AxTyXyQICp+pGfjaG2mJr68Jh3YBANwP7nsq+BNuE5MA
6dFlfgNKJRcByFXhjkxRudzLRejFuzx1cjsDpKlpivwT15mez63NjSQuyt57WUQu
RTq+9MvAvgqckgDtFjVTnbWegI/VgQcpewd35atl53/ldgb9BYvNE/RhK+oN28vW
/woQaSxd3Uu5OtRuQY1dfzxXBQzK4xI0VLQIYIlIuKyeHR31AFYcqGAN5yuA2M9s
oZ8A4YesR4KAVambOz6VOXMdYfxnqmF1fmF+9G9hguA87ORbLBk24kfbTJGfr4J3
Z8B1hwtOukj7OTmNPzJznXz36LaaMnLBd3Zi1z+LT3Bdu1n7q7QyyD9K0jb8HdwN
wPX4SFN6B/DJGoLXS48i6oz+iOsSGq+/J9Ihm3lzxqCEQ83V4k7TScKFZDExm+zV
WRaOBWN/e7NUWchNua2ARXFA7C3+lJXXzcR4xaLaieUf/tg1XSvYwAVuncgIZi9T
4SykrSb8o3xeaX3g3qybSKBbC7V5GO0dplV0j37EbZo2k+phrjzre7WyXuVOS3oH
Jte/vpDaQie0qeSNlLNNJP5aIBWHSQCE+mOZNkYR6h8NTm1x3ZpOPjmujFntAL0w
QC1EX1coyX//Sg1rSMVBN/kkHDWYC0pm8zVVbRePBsxapRgrW9MJdqFBWLFYnTnK
VjNT2cUtS5iCm9wJrFABxHxmGfTzP/3vCmQtWRTy7VLA4tarxrEnnu78A8GCbhCB
FzkFL3YEL3yB00YlLqS2nzEOMeiC5GW9kKxvL7J0tjZcCicjEoK2ufXDORkHbFxR
fO9WWy3a9gFR24SV0Mu2KQohzpO69OeruSe2zpuh/t7/FHrxTp1jk7LvkMd/n9jR
QVPZHqt7+C6/OPSqBWy4WZrJ7NbuvNKYF7oFPNocgL+MG9IaPtk5zuhysip7mL6B
2/DKmEq9NrmIhT1s+KMahV+MyZG7nKhdupxEjiW1Qpc0dwkYf+iD8EGyxcbLbqDO
KKyWLBT1GAHAFx9VsVPGqOZYzCW5Hol4Y3WQiNV6YEYxbQ47V9BKPt/EnyAP9WAo
tUt+66GWVMFY/BN7xPEnlsIC+ubMhYIusEoKgudi2SBRLORfAGBR0fG3D9j5ZFJs
ylb2URCyeoRwfo3eCt5MCLoAH+jHvJ0wCs0k4Hoqap3zf6KaOcDupvuad5v4rH8S
uO4dnjtD6iDZjq7BvnSdZvePJszkr3uJD7ZNmZb41WddwPpi+lKf6XezXXEFCaSz
hMuNn3nlZvpd7JHaW5/u5Z9Qk36YuP5ch8lmsefCzdSuLu/EfPw3rAXDpTrZb8c2
k6V8J/UCC4nmDorf9Z2uB44ZS5GL49s8wU28Yv1/lfuyML0dbOKPSY380OR6PEJi
CFK9b+VkbHcaoV4VigpJ1gQg0rhBSaJIcFbqXe3GBNdkyZlyKPAP22E8z6STdC9A
41iea3ckykGOuMOXt85scxZIYt9DMBt8q49EmLg4yCxoBB7bIyv0WHXKSP8TONvf
JXJorIMPHQfsIRtjI9JFDF+Kh6MVMX+oncfkjGJsfNzyfyR9CyD1T3IMgzcYtSUp
pQJXvODXcZdcxZIn2c4+xGdGFCuDuB59kUo9kQQnjcxz+pd3JXjRUqHGrKAAoxEc
n1RYo6orty3n5VDK+DlDWF42HJ+G8OG2zUgBh4WKcwmhOi6pCfqiL4ZixloR9boq
17D5XpynRrEHskWJEHT23/3xKDExrLm8D4qJypFNnl8D7+G4bCeneonwl9o8+xAo
JhUKSbqlLtKrxsLuQob0XYSLRSSrQDBuinHNeNxfqP6Gl8bUhl3Por8e7JreGeli
QLWYA3h5iqLGkYLzzBTtyWyVDPSHz/MCPU4nDQzOT2jvj47g+vJqE8Ms2iPdJ2QE
FXCpYw/bIUsgcoCTiSUUfLAOvalNYpbFp2w4i3IcoGlVvaaGxBjGmDKY71/wVuN7
H2DFUHwuWkI3U4+iJ7/iZ076NaxJE18GMmPvv/GE2/6MtbbYZrN6LOieYC9PRoFi
WQLB+vEkgKZ6PycGeoeQQcHFclnJXkDV7oMrrZjhXvaSS8Ki5mIlcNtlTIo3pZCs
z1t6+YNXRsV/bKTrDmS4ozLWe7AvKNZrK0unwF/U1SI2a1a3zSugHddBdpGS2XKX
EhoM4IZF93PluR4Uco7A+fr10v9VTlrq66BwZDQtfdgLemtYsrpk4KrvwJ5tid65
loTk/HYjiGUi/HF5mN6WFocg1U/142gPQNDppQP77cith+vIXKgBI5zUffv/8yyb
GVaxOwZ1TDRI3reUOzAHX9V7HzY6XQWRfOUgqe6/ASYD2nirqNJminUfL/pkp4Qm
Tk/bfLvD2frESwjAuouxWuPrObqnS59bv+3UuJVNF/PglZtkQxAHB9oarJv5gwKj
lc5rfjCnaq8QnWwA3PIvtL3zu8bcl9w2joQ852qyk7l898egsJflYDz/e1KgEYIg
LmKyJBSGKxUVhujqUG55iXfBD4Ld2g0HMPSvYOwILig7uXMFQh3e1HCf798zGK+Z
PZQRpoecL07B6gfT3P5eqqIjqQeQ38gacU+BuloaIlr/IJULebRflkF6LkpuBBnf
SpKfXlOFM4EwhgbydrKC8VV4D9o8siiOgkz2V6xBrXUqAiGrX2psQJcViqCc5uLM
hYOz8NE2bNYUsS9jd7gEZON1QGALq6942l3KR9223zWIN+axg3VF2m/NYIJHAZ+w
U8Ja6n5Mk7UVnMDVuZz6KZ9sVXNasSttak5rjMMAT5MVUYBCVDl3CDmgRVKfQm7P
XXeayMUHxwkTLSMAXi9UgtapZOCCQJCvTJwaXdVf0H/Q916cjiCD01R/BBYy7T3m
kxhQ2kZcQxYNTBCi3FSswFTdUnBRnQyhtGeeT0W7zjL8DR+Dnci8NFo5rxD9L2an
X7rH+XZ7GZlKJjiDH9Y+MdsBjRv3+wh3QS87AMNwWXAcPLVYRDmchR/9/pbisedX
3wHzOBunI7cF+fmMT9n239LKgHmr6JYGnUymX1n2ZZ9U1V253zsVYySwz30sdKu7
LSvEAFXXtY4Xdtx22h4jchJeUISes4L0jqyAiuT7lRAN0xEGQ9RLbUZ1UGAATDVj
n4MIUUEbrFpCUibqjanSWZlemV1ZxybmIsRAYuJn2ExdpSWlwi+EAQFcXNtbSzc7
/OHLxo1GZbN0Y6SoI2GdiuVFuO/LX1zcaPdoA47MArNBazhbeTAZQqJMglw62XUN
V20pu35EguTlkUVsxbwUMEL71b6jdx5paYrotb8vz9zfI8jYVQLfnvQM+b18L7dH
Qe+Ot5UDnIK9vZrossa+RuC18rUiwkC4/NRBYUPLTsgnFmJ/iu7DdNC0Unu9RPwr
HuzfeHnEinRkRRCzHAlmJf1EQ3PRgnscNMpxIauyRmVum9CC2Ew5uxyYvQyyJitf
j9WkwS+F+I5K3sIrrL8etr3jjSCZb7Lo9PU0s5RTx95LbL7H4WHk8al40/UBVV0d
dbnN2B4j+C15ryqjgkeeJYU3axYqooc7Hz38I+/SxpBPbB2NA6esEvWXvqr4zKTl
jgBPMRr8JWHzp9r/3XGLi8OV2twzwv/uuLB+0BgvyUPlUqz2/F2rEyye7O40Cqz2
DS7Uv9hhrCjLLXebRsVdgJclLfWZDv0gFsnkxcN/VIyfb2Wo3CDY7YRk31P81Zbi
Ok2n1o8M2lnvuR2o5q8+83hv/jK+hH5LA9dxUFf+NSd+c0zo2Zpfs7tzH0m8DuEF
Dh2r3Bf23c90T4Fdp3/9RYnc1ZfLbNN/I7YptWP2qjfDEpY4Uk47olYehVCUxDDX
v11YYhegif34QoFVHEJKRCDIZFj91fjUFE651OAiNBTuxapmPRntYuEYx27uXtDT
G+LoB+bOcpIB7oJgg/ZJS0yH+F6rTHPJ9V5Lrl4Ie5gfsdVFKGT641c4QeeQIHSH
4kjaq4MrvMejRONEiYwWPLBJjx65lAowvSF9ljxhdCTgBFiB5qdsbsItThRJ77EE
peZxt5mfyuG/WGZ+b2E3Ys4IKNFu6Rp8LG5k5bG/yReFjb5s556geuY8MTgVSy9S
RAmg2EDwMNsEYwN1TAHyj7XG5+0EOxb2a6m7GxgP7qyOO0ByxJpsF6sr3XliQ+2R
ZxfAAD1UYuw5zaZms5gnDEd9LIFIzxdsBDenD/zZYGWGje0+0u0HOHZpZ5mhdNPU
Rb1sNevfwO6x2AXIM3FTHkZnow9m4umKZR70FWMbNafWpI8xE4lqcjjfLx2sepsp
j+iWsSflmH+dbcRd6RRefRucMuqUyqTCnugDIb86gG7nQV1GzqqR04+niCOwT+gz
SGEc8NSdnTb0ZwWC9Ma4GMrE8ntz9biT28nqlI+s/qF1mkq3Yno1l3iV6EE1sVAa
izV71IACSRfEaY/iuOhWAaplADxttA5vEbLP+zldlKJkYGHS9rkbghUUMpJgFNOm
RXj6InANgpZtfea3py7m2sf+1QdMyLigaEI6xjemLvz1UMVksTxgpOMQtbAVc9nO
veY+lWfYmXGnyYqp7WakKA074u6GqMPdS+Y4F+lnKNmIr+/FQgLpndnOvtcF7Rbh
YRco/Hi1gxiKz912hPWaVgf0/3E33N6EScJn7ZvHO1+qEilBKyeiNHIC12rkX7Bb
62sJSLxSC2kLTBqo6kDp5DO4xkFTyY80E/c9Wfwo/QKyOvCL9WbHy+ynvNQwPDuc
jhQoDkjU22Uk2a1yiUoe7QYNlcpRKLLgu6BZO0MnYKFP5NzqPmqRCae6QaHJB8gp
h8XI8GpAckoT4vCIiZPKhQ9nClBajLufDWLXjxm28VCSQoLax4hQUNBDbpb5oRDU
GEWSrdisgok9Stgp/LqkXRIZF3jSeiGiKzzQOjxOgA2FK8HaF81agwgOGVwb3jT7
TEp036vXpgd4HzxYSLILcVFS/PLcKHg5JN1Elhh+76dgeAVQ1mwHHtwTPTw8WjSx
0H1BC7FnhyI+RsDvVB7YgeaOP4beIhmXP1J0Ofsvitx07RPu8bi2lPzVOsblcOh3
bcvArBqDQjM51LYCBTAIJTN0M/9usE6ppfD5QUIdg6h+2XRQiGOcrkvxHE1Fdh7W
gCLM2uW2u8cyQNFnxBKsDtMv4DIQsLrTeMsxt72IKVG/or1OyFHg626nArkQCw2D
UYHCPWwWLYOgHRnPXx7hbrViqSahFCr4euvu+Rv9xlRArNsZutzzvnfaOSVqhqV/
d0Rcnh14e56JpM++IJSpcSp4d4RwqoDKFeXPO5T/9bhiatc58zvN9Nz6OrwbCHwl
biU8PhkKERz2xVGTVs4wUQZclrTr8aJDoiX8wmngWTtbWqFj6vTp+k8fNSENRH/p
5QeYbzYaEOt5HSAsQpEeUtQuQFNIdR2AZrAKFb6c6qpWttmNQThK/7BB8dd7Y7xv
ZZ65u2gr4qrvua2AeTaqcztTLZc0sBsAfqweIDs0z20G2TQ3zs4dfL/gx8useuEu
A977kumqK0NlOuR2m9xd2k71mEkuL1eChoyR7IzisJjBb+0NLj7Vg9Rt6x3z6/lX
YHyhN50UH4iN/YsEOsui/fEMCC8M+ZpwKzSVxl3dmKgn2DyYmrJAEQYAkvoJtDiA
cM3IBEw48QIIdgEKjczElBpDTMiWzR9ZdxEhNqbg7Ruq3fhRhkD6QKmV4yase49j
L6Sy2KjakNLoVqZWnxnIeBLTDGsYdo/eF6fGDUSUY0ikqHZ4sXMoMyJKJLyGkdr6
pj7BjbTZQMmpASFa6CayttAv/n8mLW63ms+MwERzRdBlp9/GFz0kIQPJZLsQFmtW
LVqFS6d0rbE5UUaEMWOunx31DLJPyaeVxNCqeABpaMXHfdEYtKWPgD/5ZUtY7CwT
RuipMv6ScGSt789tLzeNrInc7aiqdc4xyzjA2mNABe32ADs63UiU5PeLRam/nheR
CgBJDRj9V2AlNrZgWCL8HlQQnk0ZuTHUuP5HRBVrUmhkCvRqhukEpGTHuU0gXd5b
73plag+3cbre4eXhPFUgRjJZmLfZwzbyKpOi8Btzf3YTn6EwbrP0jr61bIKQGE1M
1rl9rCEXB5p40zibOqF9m8fADSX7Qjc+IlrvQh24YfIXIsYX+2kEE7hoRbV2SiYu
ivzr/2W3OZf94r7w3bLJYYC6eVsVEd+cmDCOIE1Cvy/4yG0vrklIhh/H2HtErtla
U1CfhrrKI4X5Pf7j0u+HDowqcVw4b8UrtpdVEefFSFjIKUmtsGvz8aIyDbJdVEqp
Z9/Kt23kQtmRE+c5V2sTyAYS4H32o1GlaMQjHzTulCwdMiCA2aTpxmmkkg5ipBAI
uOH2DLLlRaala3IK7fjKnY7Q9a3nFJ9fp5uUlrnA+wKrCGyXOaWjyrdjifh1vfCE
A8tLTZKkRMxqzBV8X0MAEG+e/A7v1v+QLxSfEh+4FmpvDcpOgcgzi88qVO3RwgEY
bPjxf1EE6QzkgmAQGcCva+EFSuwVoxHKWUxIfDFJXAdlXzU8jBVbOomPIXKH6mgV
80n94gD//HdksIsVNZvYTYCMf85cVU3TRN1fpbxGXQO5BaUBgi2t0N53gjWIctyu
mfxp7TCBEC5CWxwtWyZJY2yvT44EbpkwnSMJXYfdMvgieAIA8J8FY0JSWWVEh9cG
WbR71+EQZhO9LcWUlCgWzNe4O9t9Q4CRc69Qe3Vax2nG3mdMOY4X43VC+WJBllP+
ZA/+6hPtKj/LBPULXExlUY4varl6i07mgA9H+ti1UONHtvPxwjDnfAi2D3kCp5Vg
MGUwv4ncGbh6sHituDHzQX6iq6Dwa45gKZayMvUhLKheHu6kzozBk3SSDJNVMurm
r2VhowIR6dsSUdOYHRsPHVTjrmQXL4Q5ILBBT/PlKGtYWutBi9uZT2e8RrjLFGF+
rPev5KAuUKzxRtCBGdhGigl0jsYcm1C7LyYWp5SMLpSzsfuNLzgZQl0e1AabN5Cl
FjTMt6zsof6q3RHicPw1bK5UgofodGzm6mRRi6aD58h83e0ARvYU/uizz1lKSOLr
mHngnFqnBnb8h77nqKd6XR4eyYmTH1b52CjOtKFVXgSc6A3FINC5MWEIKhOF9ebO
pk+eWV+vKsdTQ4VeVJhuApvunDtdB75AukwTRlzRz7jgfuNKfxxVbchQHTLJZXN9
DR5pkXwQ0e7z2/F22C4SJex/3/NQdkHOtfgWU/nhmmACbWR57p6UF++HBDAxzj5n
5/Cl0QcK7DQ39pdygH7NkHRwxbXycuRpR9DTQw+5l9UFgPgWukLrk83qhndh4eXl
FnU6wRffeRvdNuQM4oShrOVjE8w0m9Rj+e8ka5BFeoQCagvWhPBGfwnw9NUMgrBX
5aO0wP1qCOyDBEhejBfopP14x7s0EtL4UeYin1IO6wpqLIDa5znyp0+wQY++ofIg
Wk2GIQ1GWnOdTyv8+UQ6U2nTCPeP38GmDQgCKbwT5ZUAENb+1OFiCa7PlCfps5ft
PpyBP+ccBZDFJG5on+M7D6lEGGiezmdeI1m57FXbBt1D3UGEGTw+zPHUw5uEbNQv
1y145+4MIbcf2j5/ovGx3jVMobFQU7At1FRmbdhSbCtOA7BQGih3dHD0LzQS68Wr
4VfpfQYVTCWrMK9CDm5xE5vPiFPvKntmonqhVTwgx4bBBCjkDR/cP1QBooAbuJOG
nLNqe5GQGS3u18sHytE7qLJw46Cx+bUYuLjfLtpinTgt5vveS/iQpOgB7lsvrmaD
8Y18vSi7sjs1kA3bncPs8NU+16kDqu5jzyGZDZpXBmT6muaqnaOxNqtV0bwMI1q1
y1/4Z0ZRV82yclqvHZP+OQbUsR8ohHCln+WDPE+RQbcbhzAbaTnAuzFZe2pHFyy0
pgk6LOgyLmxpiS4FfJ6UYb744tItLYff8pnmuJsMq/wJADOuWEf6RGq4FUK1MmDn
/N728I90XXAp/xwq3xJ9Ps/fpcrdsal4mdIhS14qIKt935djl9HrrXzrAqKkNirC
P5iyBf90GZi7OOghuttiPyEQpu5pEYNzsJEJMtHzL1wjsvWAiCX0ktvF30t4Be72
u24UVWrX7q0tQf15AhRHDcnnG6VG3t+JAEUyITD1F/R6ITv6zg80pbslvqlJGBQW
AKW50YWhX+bXnvUeJCJuWiSSFBHCrCmzrhGeG1HhyirictrclbzvQeLGA2dZ076S
wfoQLa+bgI17uOFqkUa/nBUiqrcmyeNMRpYdYw03tKu/KUg41QcGZ9htcX5kIinN
YPKZm0Eat3AE5FaIFnOCNXqiwgSc1VipD7CBupLXYzc9h7eLGlDcr9VYIUUvofnR
v+527w7vOW5fD9epvcEVgbZlU7/O+Jxo1MM2TDQjOZ+kh2HfntTALqmYJctjuoys
l5ilJ57jXU6CHqriaeGOj5GpanJF1d2OsEthJGocQnCVSfnkNlnmWVeEhpRKBtsa
vbP4pfJerhIw75lt5wJqXWOBOADUAjGVPbzVi9V6eXQRB8qCZ6HPYgW2dclymZHJ
dpR+yHHNnM/UL7tuz2pwCbheXKcyMmOjmUrxxpva2nEmUvVQKVYt7lrJhwZ9wmIt
BggAvKJIigc3zh/CHmy+JRUD1qIfGtafwNrRuv+t+JiCSgCAXYynGcpt8dH+gTcK
FxV+j6TVUpHP2hqyLt8V2NN+A0aWJmHMaKaaWcgwvyAZ4ck9+AlDERYU9tzazbLs
f84BWQ9eimXptAOUy/r/QuZpCgtlU7jlpoCLt7JRF3Si8m1iHygE5SF083YYAuHZ
k18u3bEHS07SeehEmZ8VHOLuKF+14dvCAVWAuSFewhCsWpDajp1DQwAogCc4/EwG
A+7havxSGr7ci+2+KaB8BENCZLSL4w/xO6//WyVRjYHjMYF7dE20VwmbBWwKxpZ6
EAcIVC5xwz2WwctH1pxJxG7VhYdIBGfDGszn6ntRgoUtsOZaX93Zd2XUGTq6NeGM
Zo4gH/3j7tW0pLjq+RQxH6tahfYkoKCi/dPmf9LcKgCwym8qnTB93ikbwMrpQ1Kl
MOCgiMfaPAvNe8bFTD9I/YQzYqnY6ckuL88wDA5CF+GEhZ+/moeVHtMAcz7Vioml
jNjg84F4QnxoSrRApmdXLCLCVOFI6qwQpzTKh9crZDrjcHO6BevA2BTpDVBd7ajj
GPioVmw7R6FXDHHL3TeqYvXIUaK4/d72xMmhg0Ou+9fMeyThJs75k+Gw7L/9tzod
HuKyn47Bv0xekQ1yP8s6Mf/KmUrdX9qKfSvJfTHdfLbzPqHc/g0HZbxLwA15xz0M
GqPF70vfIyh9FkUecoYZrzld3uUZwd6FDC+AT0hKJrcI2CoZBZtvk+JvnyPSu2WF
VuVwfBAlQcZIHuWMFsPtgL8q5Uxg30BTJv9KN6zBCvH+BS4EmDVLovN8OLfAnVHC
qdKTL07HUQJAW866O/+iu7R59wQ5Kqt4hTyJpCN4wFwMCN8DpldL5yY5AyQ3jmZ1
N4BINsLYCETcYac8zD1jUFT/BIDPQn8HG1mwbPr1MfFQYeCKTJzuKf1frHoSrT+g
onBfpbhMfDg/EGsxk5b9VSuNPTBdBJDkGpGdQpHfGuObJerzhBRYmVgrw2svEh+l
YthePS8KN7IZWVou4rZNboJFB3bXzCpaOe4c/+18oBxb44IE8WxFA/4eyGx2RK+S
1hjntG0UA65wYyHwuhFATv1KOFxyO9sKR7bbYsU9DA2j92E2yiIxU8Fk+8VUxhKw
TuFjSr6oQDbC7NYW9yVbYLwfKb30ilUejuvMl8ZpCrlineVrXkK3A6WS5mhbgfoi
ugIWHGGR0MPEWmYhDC/JFyBHUThp7rK5ySrZLRJNMTOQYMd8qBz+l4Sv9y0a4tla
KnDAtTw+U1Ge+xTZVSRn4ZQ9psIHg/PFOGfIuZ5XzrpFVPqBmuzKjE11Xds0G5j3
wxLwdaEW/w7LSvbJrfAdpo5zg3ZYxuhVAZzUsNbv9JVgus8c8qq7s7QU2uYKDdvN
/BJ3YxqSYKLatuimRTlOvp+9jeWev4RzbHQTWeJpUOfUAI6H5r+aLsZ2iqwlANaP
lyS96nHf+Ix82I1eAKVbojkjdPzuxbG6sla7WVFFLNqSLZQAB/Q0OEPgUsx3AMJN
hkmgQ/n5ynKNEFr0NpQAa3dyQHA2ZXLVQ7dsBqvLAAovdF4AX8inp7Q5Xro58O5c
BaNHgjGxN8pdEiqPvGJaVB6I5U9KMiHwbnIUyoZf+GbYMSFs7glnkTsGhllNvSub
5+89F+XcvmuR9rL2CDPJHMYLs0wKXXosTrukkA6XfL/NewPhWI4IJIXm6IHNMbRH
BwH61zHSdDr6OLu4/BGJc2YQxMCR/EyvM00skPkUHcqTTAeyjEQPyMQw4BuHZJTQ
Nfc5WoffHr8dbL2y3Q/btece7y7KsNK7LNWlP42vebdJqOlgAr/iIQ6bHUFjonim
XgV1IfgdcqNLyC1dtgd8cLj+R7l7BouC6fBRv72d4lGDZ1EJB3aPELq5DbIsn8GK
E6x3SJv9/7PnegtfqmyPdHg1oxQG0efz8qYJkjv72WsTT7LL1WUjD3EI8scy15pV
M70uhyOFsrzOhOmb9jK92au1zUXLfoBKg0QnYShRMe8dNhiJnUI8Z8+VMy1n7kBm
Ip1NQjYJUppEU7LBtpSaYm71GdQXowiPCKbRssFeTfORx5y4s/Vy4igj9TuaK0mg
+xPaWZB4vN5aOWbcohM84ibNUKOc5viAPH4ekx9l6MXM0vZLDR5i+K2FHPKyVxIK
Q3jkb1N7HELHJOrMqRHkaAMtIoDXeFMPZ8QgnZkjiFOyBSnI7g/Ze0yzBmU/ERh1
kLsEVZcLYHGFA4kJAz18mMzdtphp+5U+AK56EwGGLckLPhE2lT6RsCW0XcZpOZ22
b5ql8uRcBZPgzBO8kE/Sv6Kx2Sh50yMcn4nl6KcM2qiFfcu5RemrRroLULKw9iwm
ESb4aYr31qWWxYPY1wsdMB+esg9WgY6Q79oTHE6Pn+xEV485WIgKQEplz8YKa5hE
NIdT9vNq06pUT8zWKbkheXdsQOC3yuZbHYwZwEs5CG+BGws/0diKALk9GnhO7FXF
Bqs5i5j3PIJOz6eJZ7UOx0GGRaXvTDdJgVELSqtklBXXB/uhy7H1lPrOa6dW3+66
6Kik7s7L98YS5D7HwZpLDOGk/2SpOt3KfbZy0d3pLwjFQqnS3J6JV1Upa+FLL+EY
nPx0p2M1ANia5HQZ9syYVNOs+UZTf13FYh+/sbMXM2YteIFBlADZBAYQ/z3151xU
leBVN42RD4FFYGri/Q5VHD4SWQlm3MVS+OV/ahZ+7vq46ozn6Jj+BhLqcQ1b78fi
N/1eAvvkFzy300B+ZjQb7bsf7zQTy17AfN/0wbWlBQMBeqgV4Z9VdT1ouf6mNRKK
jtpinUrzM+JbZq/uiN8wlkswW8jm0z+fXuAMXWMUdkzpYjmeTHSZD4jhfCM8QRsX
O6E34Dj+ZxrnRdJ1iLnEqeP/QVySztsReWLEsuziYyDx1RQ5RNERO7XGUZy7ekO2
lkfP8xrOkRCH/jcZSy5+Yg0SlG28qUG6SywjKdqnaWM3GwjbCzH3CGknWaiBdyfJ
9K+7mK9FJ9W1XKj8OhjyGMmE0ta81huNrKs5cpuJrzsVLy7bjvMUoyrpUlDEUU1J
viZOA5sioDecI71tciwYaq94OV5KDBGc2K5fYWCzrVQZ61bxtP8E+NqATyeF0BeJ
C2An1qx11ZkqIAV7XLpUt1r/hsJ3N3hKiiVAKBfgpuCBCVkloaqj2wxZ7N/yNtm/
z/5tBfnVbOIgpDrU39tdIBsKNuc1aAtAQFXvJbjSg6Zb7wpSXVbtTAIcc+CRXPFQ
R747KabUDAjmx0MaDMy6+O7D1bZYKHuYrJXVwx2mLb239e6qFV4h6khwDutfmWbp
VYVA9va1P6owDYKcRryB7smidKQwS7BE+HFYXRwOSyo8dPHoN1K7/RzBuYvaOPAf
TpVckYF/0Zvy6bdRPCjOMQF3c/+dKBHVLe0iCc/1YLnlbH8BqxxnYuPbXPoevKxc
ti6tGS/gNUVTCQUloRQ+cQfjKnL0T2Oye1mWUJQ3xS/e4URXxG7ShM6dARLxFd21
VncRgJRbCX4zckuOW07Juf0ixZnLmbqKoyUEO5rsEf9rhn4HcgPtCQCD3qFjG22F
UXHfwbQQmgDL767GxLIQZhvKZw3RngPnhkzO4cSymz/qcSN9f50TrFZx6xxQjCtL
W4iXVP06uIP+PSwH5VYC2WC/1vvtZ8UKVNYy4joeKSrYB5ytaMiEMurLTr2tzNjb
e0C/dmrGswFtb7Ux10u9bvjlDP4jvdRmT3yQB/18vLzMvXlx/74m/xEr3Ngwr+AL
DucF7hoEggzgJaQTUgUvmebTBf8KGt+QHk+SsakVtmfoC8UErLJMzr5hmmEu/kpJ
Gkgznvy/2zDqFibi8u8cEWAXmYMwfXPW7TP2hZiHh+W42CgEqtJ7qaVg1h2VKfhp
yjLENox/DnKrf/oQRZ69BfmeR+PzJL8pQ9nGJ8twO2O549GRo/REudOYtNHZQDQ7
P8k4+O7bQKFDA0bNaPWNGgg6g7MR4lA5kYaGjF7i0uU912YGJaOZtgyGd2ZQ1J+t
xtIOuFbOCMDD7ZkM3ONYLszF7NBhHgVfO/5e8icSSf24ETQvMXPLmBThsbDHbOxD
vBiZifBBfEh9i0pzExho7IB7FAK9ptPA0p6rENWf95LMyquOEnlhdnAXJdOwX109
PeHCCMEgIfhLTZNGPUH8qlHbDGF7qMx0DVzT+MPtiMeuAk9mweX6ch+N4dljMtOU
jbv/cQqZZWvj2JAyF4GcXERoREcF1RxTi5ynEHmDKjzty9Kq9fOzwAE6fN+Zjd9P
/A962OOAMLAxS9xRuTisPH1rtVVzXu6UDtq6kILbgvdcKaKzPGfpIGKLMtcSRk7g
nbWSbip2ZERHPwAhW+wjpdEt0JhsVl9qRsjZ+dDYBIlwJ5L/MlJ7K8NdsOO/BkJG
mXeADUsj5Y15NFShwPNs41fbzS1wCjQcSasug+XTajTKI5ZXnhnHszlFbxiZ/Mc6
qi9nnPuxjJ/2Ydvb+ITIB2UhkySlJ16/wHojtLBdA3YqhcwrnCdoPVw0ttcJ8Opj
fwJDLF476+HlFtEVIlzA800Ea/Kr6Ssg4JFi6F2gQDMkKCGID3ZDnjI56dVvQBaG
dQbwS42BAEHnZTiycUGvdv9fZhV1+3jrWhvlmxNT5p0z/NbecXzMxdOyAOzneQ7+
QVyK1N0wUgJIoFm6dxuFM44Jbzvz3jMAIFC8bSLD1unZ3IrT5SUslhIHhtmVYYr6
E5eLZd9fLTdLJTyYCavZIVG7/Dl0nXywfgeXAUXym2gbWBayD4NnGzaCliiSYq7d
8KOy4DXESFPmMXdN8d3MQosk5CS/bAd51NcGSrZh5jTmmQfp68ZzNWPbJcdFBMrP
kolNfM6O6K4aWxSnmokT/Mq+FFosmW3JaA+bpih/Ra4vIfzdiPD7hJo1WcuNK9lz
a3YEmg9tDj4CFbEhQISd3G+qwCMoCEfrtLvcYu2fIjEhmb/gmK4QSNPw2k5RIpbm
Le4/vzUKIbjs7bzSZZT/wDvMHSx39nQItpJCl+bFcJOMMf3v8CdtuypolsMBP0WM
OD6qMLc1hvR2fHUWo1oIECjroKjewrzYBheCbWisK7OFPUcdhEXG9o5oYy6RVauc
odfDrH8nyO10rEJX02TfZTW8AgHv4wmGGgIMFAtBimqPtGvdSywX/psE2VGHzyl1
ZvRd1nWaE0h9spTn/xzEFa0KYVAevYOlxk9ffUQ+etRlinJ3YTxWKKLr3p+MTL0X
MhS3+iOwuddU08I9d/7l7FIMLUbEK8TPWDBjXW6tduI2vwKlxydmgi1GfzMIjmZX
VF0voWUBdOrwb6ixMVNwpCxLOElVJGmhZFxdvFGIW5yf/+AX5E2IOYvRFf1AjaRw
ZMh96KyBvnRFWkywicu3rG1Uw1vHST+aF24T5y44m8CEhJ6WRVe3yDOSaOR1DrYi
dSPyA1P10oSkk9VgpAElTJr5Ul/l6Jo04SmNlnJZLzSm9tVuw5gp0tG/vplfx++q
rKA1a/fBJvN2qbta2ZBMMnkgv1v7Bm7vDTOb9Kb5NJc6ilv34O/yve6SpHEpCb/q
gRwjhxB34JoHPbMrC/9fKTze8LePo2yetmmLfNd3zTSjhK6jVJOqM2vpJrsj2SYf
4C4FIeRym0YZpStc7QeEM+JufzaApbGmat3wiOYlYUDxwZqBdV+XKRjgK16kbcA+
56lsX3aZmm5NAazNaCX3szLnpD3dxCuOXQH7lkUYBC/A3VSygNQ/InVw4DRTqMUt
pJ662gnSv6ZXGMpvCtZlTYax9rYFWUJRvxaDnWpwAVt/fvpgSRDKTRLMd9xcvvlr
YKqegTUWX+Z7QiYO9E3lBZS9IKV0ofaLkiHBeBLJg5EfFuBf0uPH07IZF6yht5bx
9Jz10vIScZoM+ueescu+TLlJsBf2JX8ThXD43qHzAbyTyXhd256DtFb/EjdEfqeI
x6n9aYdUbcZ/3q+jeNsOjwqYr/q6otJTJicCQERjhWHeeVkZSDbajShHItTfNG8H
ESi051wc/jmVw4m9LzG4wxTxKSQsSHM6CSiyKAkf8lU0GFOmi9r6g6fZYFTo87vm
agjl+XtWUJ4m4/9FDR03De73vC7FJHikDevaJnfOeNSN/uTOtUoQ4VFmgIiTuVLZ
3oXJ7juWaeUC8jv98wJmFoUE/8kuoNiLIV+CxdPXa+8j8xpA1hM3tb5MPPfFE1yJ
DRJ3NNDgXI3iqHc5L6gFx8fFPQ1RN9SGDVPgxG67ZvA1yBffkr6CKRTIFVreOg1J
YWyI5ndMI3Wp+U67jLiDq4nTg6wxhppLlSj4F4GoWPpk+ghp9OZ9dNUd9tftxGfs
a4lpbRrju9TjIexr/h6MCiPGzEbBtoCiEsqPj27y0UV7SmHp+Hf9TGXFcsJ7TwDH
uHHonocUqW20q5J3tOGGvJs//U0nhsPgjJoN2NjmnnOqKHZxCV0Q83Nm3g18XtxL
QJgAwgBKL47hp0mr8lOL9l0A00//GtnGxql+VXblWqkwarA4v7K8x68ZDah16z2J
vRISvaVHfWQrRUSaeTfHaE0LFDXqibzW+KBAA8E7dlUeHfOc7s2ARfCscTQxg0GP
jT2raTTDHtKeXLTS3zDHfjRL6gSM1TUOu9Z5p8QWNAehhnHi8mzEpryOnEThKB52
/H+s7dlmtMkwMN46HWz03Pz8XfPE0MMtwmIcUVFoupBlhQp2wqvBMh8tVpoVg3Cq
dSSX+SldPLIArqnofmntK8qkPu0PVO+kiHpJ3HlHAW30mzdKZuAjvwuMvxgQa2U4
/VmigGP6wwsyFx32s60usbdLY4tXfQrjenn8+E2Q2TY4lujxdhQwrWUouQqzxH80
WPUzOlzBdtAwpK9LlZJX4bsuMtnNMiXN08wl2OGgI4HTdKzxsrnLqbQ6WpImzYtZ
iDEJJbGPvzS62citcffb1rbR88pVa/alQk22l9Qwl9sMnwL8AwALEA3WA+EZgneM
NkBs6d/FNE2x5xrNc5V8/5beR3hH4DOf1xc7z4DH7V9EVU74sRX/+/5scFNE7/XG
FDwNYNrf/K5+eMYkF5YVJMfR3kUvLKeNU5hvqRorjYCgv0WHWSb9hM3HoY15hrYn
WdwOnwKM/KvEoTbs5gb73GG85ALcKzkg2YMdlOSLvmPzAZefdgaNO0Od2dQ0Hx5M
ruuXX4Gx+4ik2Lcg7BgVCY/BdNtW563hv9njSaFxnPz9MHpfwCHZ0jPZFi03uvM7
ewbGGP0nsyYJjAV7lAsq40nJNo4ciyEeynCcPHlWhf7SbIqbohGU9vxDcA9gQ7Lf
6gjQVlpYEe7WGB6hEd+9gcowk44V1PqEg6Jq/zVytZuMgjdyc+elqqx97ujwLqfW
qydYVHFTGM2vcU/W+EZmOfUU9N5jWWIJUK1qUqiOectpoUZ4SmaWPqYh1TYan3Fr
3cDq4y/BwP1Mv0rA+ZP95nagytj+KlZB5UXqlk14HBdJO62dNedFnJhCwOp5aIR2
KfFWixRESIAdWDpyqT3q16gMffLNRTtOYbRjDYYyLI3SMzvMY+yP3ep7qKSK1+5H
iP6bCLfUC0ngC3SLo4+rgnkBmzxzgRVTjrspueaf4xrVIfQSRfv0R9sm6tHMNcIL
+cQFzi2EBBdn9yYiE+NZjm2vFP+eknOM116tLjWHEt67A4NfbX/8BjhoYuJMrNNT
ZoiTX9jB6WCTI547gWBeBYJ7eSWRLzWAHRrNGnpAzfaVZx9SthUYarIsWIg8zqIT
fzelxMaAoZXzU8znbJnTsLLl/XtLoQCN2IaYTYZ7k59In018z+4RX0+2Tu8ZZYL0
vEp5ZabuVe65eC4YUo136g5QIrSDlAUiu1GUk+i7q1cxbfz3KVvF6BDgO7pEi+Gv
3837OSkG3SmtSqOXHr8gR/L0/EweBZKHlX1BAzd1lAf23mscrVISmnYYKus4W3vF
9JmmKEt0aUSzM0Njjn4Rc3q/4r2D49wpaTlre6hezpb16cXdj4LagcpJogvOYc1C
bhxhjVrmXnb9iGaiwMlbVkSeFNSGDhnl0x4AdueoHqydrixArEdn7AsBHiy8e1xo
Fx65I5qDIPDhnKC1N83spihMn1JEWPtNfv2HOQruMCbGXulr4er5P5F+mj98iEBK
4nRl92wI1dhdlGZJ0K+rGMvx5OcYchkWB+PmyODTWdHd0e4OvLL4fC8qj99ntDQq
fgWlsWC8X0ZDkgPLshyNVtsDUF9CeUcEUd5Q3V78pXGV3tpqS9sqOYdohP7NLKeD
24r1QldtpjloNYPQxAKivTd8iNmCtVX0VuVQsYACCE4O/9WPI5JVAs2rbv5WCNLE
eFrUWl70iA3ZERk0PK7QSLH9BLCfhBXx3oLtzDYkXDfp7aXXLv6Xco3T7poO9cna
UwRFLsxHBesFfC56q9HdAbm+CKRGNlske4PMmVeZdC6LjculbNFuD+xu4JcBVgJj
dhpbpNqNgjQB8DQLbV6mu81d0y263JwaJLHE8+KLI1259q7n0490KJ6eTh3EEFa0
1ADu+NaKTEMHq7TCgSHrPP5ycpAfEGAW1P29NEYEWMMIS1Vj0031C1y90Nk8KRJX
ZuYQIer/PpQ7f+Q6+/WM9YE3mzuXdZXJduiBcf0GOx1ZgOz38/6uKvO/kcsPiZHh
bhcC3h23jKCzrVoELrX4nNR7sHG3jVHEN5+xHns99vD30uJF3RIBaK2wj+4xD0Zt
MPZGnBt9oNYUfKMPmrHXPqe3fTS7OMd0XflvXr2L4pnzvPktOGOTB8t6la5bSbpN
ZTTZc1cKmHmLXkyX5m2bqG2w3N/YV6DXOrTFlr0laf1FRhhkV2IxjO9o6KuQ0RPl
+kq9p6qFmEc5GAL9brS7T/Xfgzr6Jx0e3gOBryvnnPbwmOAPG0cM5rq13QNE0Vv3
M3DwyP+/3/UnVYleuv9g3uiosFABjMoGqjZWIzRaVj2m03z5tzveLdCJLt2u9Vji
773o4w1+VKCy8ImGLtQNylVFw3slKWXBpRk4LwopiXWPqsvrVpDCaYYe+QJwUqzh
kFomw1Tu/amBTZ4gZDBy/QUE8ZkxaCY5gWea5LH/nAYmE9DEwhXmmXUTw4AQpT+9
++dcMPdkneleNodKsmK4mH5JR3aoUg4/kZ3n1aTlz8FWKHMnRUg0OmFA+IzHkBgp
0BobDBu+KekQHuG/9lodGg4wtPqzCSfUNIrIX8ZuhZ/bulpFQqqGKn1+INvGEc8A
Ctha6Zn37+SBI5+85CQDNDyM/2ABicDDPvLNaNcxx6lkQUCOEJSK78lVa0gQ51Ot
feDyRHhaqB0xvnlR1WRLA5OwOiadIssPbYs8QSTLuYlDlJOs020siF9p2a72AdnR
fM61xpjHTBbuXRUee5UuZ1+UNVZihCNyIAM9stlAWYnYnQ3sgKZMx1yYDY/dfZ/Y
bMiw0zMYPDJFPJOf+mM0kXDZd8kBphVNtYJyuG1QD2yIykaZcpePmBxd4ZCsnnJc
iOPR3Rx/6G32hqh2pLpnHxR6XIqiG9/umyOmetAdP5Ki7veuGM+RcGwozZRkt1Zo
fLqrgma4+xNISCCUvV6OP/sDsmgn5yFKy6gMK7If2fhbs2zS53F/mSihsJPZkYV7
cQAILJAJvDximYiqJSVMY6IlVx1IE+gVuml19JDAggSuRhlQL/wchWKPTD4cZbkf
16M9kPOA0wxgQBBIUIPsdR3+wzkEWA8+ZAdkmP8vWgvUfCTND7GWlFOlY7YAiNF4
ASe2wNsb7egiijlVkobNu2rwKrPnvJRriPlPmO3BfH3hpybIug0K6rMVnMPShMVq
r5yEsSGuGjzXth4saCEKkkWEvzL4PjtzY40sXfWztTpLZty5DXM7qoO85tM1Rk23
FpKonrqNJ4SNKq3AMXkql6D+HunKE3da2Skngl0FtxyowLeECqNsSpuqb9Cq499M
dsJD1fjRXLSnh7MIpUFevncGHwtFNUZCrg80tSyxi7G/LQjHvwJtydfAYSmlG4i1
88ADTkv7c0IKY4TQG/VFZcqNMH2UUNxm1suy0wKhRZAhBjfFbE8ccWJPHxRsb8hN
GCBZ+PHeapfckK4dDlIw0wCvd83GqVE0WgtjdCQ7EgjoehdiN9AuyM7GjbI9c089
VVyZzoJjFBi+Udlh+FjcndkhvgIiIY7BGZURdB2vTXhgBPsCTblCTU5lhEOTMdc4
Tbu3MHNQ+eAkrRW+4+waANHOeFzjkOiA5ZEuWcWrlfd4pjgb4wYTFEv4CytCvboM
gks/lsQQ0FbFcmc50AXzBDtuc0JuoWIiGpM5sdxYNurq3rGW2Sa/MGQASUIfSmPr
zF95JCwNZppN5uUwSeoH2lnXyAOLbEyMSglzc7VpktSp0N99VYpKOT9Aerd1KaTe
Tr2Y3FVyxJCh+vKfVbax4HPhvhRP9yAm/Sl/hQFhzpH4Jm9Xg8NfwZmDoen5Kp5b
aE56dA5JaBnERtOEInDfHf1HhgstIQcRZzjH3FAdBUMryHcyYlAl5YQUbTAzeexQ
vUkGh7jgFHDzbvfaNEf6pPSP5XVWS2436odocJyKbi4DEaEof+HREAHYUy+OoCQR
fL0I2LKt2TpejVD/nygp+GmNdG5QAZXO/w7UTa+DJZ6sWWQvOhOCXRs5Qj2KJxXs
Sr3bd+4HboZt48hwp4Xj2YzDoN71sYCx/57ut6olc3xOqFpN5vVpmU4Nx7ErkaDU
ezRP4qzEE9PHsY8tLYdqwsFhMjKJVxqbG04nvdPOXLIEshi4g+6CgaeTrAQe6YTF
8vdU2OOMeF30ia5p0EMqNMc70rL4GVHF1uD7skxH9DEoTqVGUnozpDMr6jcU9WR3
Onsx0jxBcgRkg+JDx14k4PwSaoiphetBe/vHbhpfDv21mdLuTdoZCAEvPzYt+nVU
KEwZ2o6QMh8aajjzpED3E76VwnjGAEt76Z4kYu/8hPJa6g27vHN0lKxXTEOmih7i
Pptv0Xo+bz6pqFp7IlbXXr4tAK6XwSUO6xiBS/tw9ZnlPxCpNA7xVjjp+frASjUQ
GIjEhSVhg0YScmu5A1I/QMpEd1/lxqCcoPqGJxw2acgjId4GLfL0F3o5AMesZy3d
O06ywRdsb6OC5UJHZyaD9qMeZ+iBsKrqY+OgslxOQMccvMTfsPyLzkWL2y7ycUHF
RvRQ4WPQLWWIZYLy9zPlUB/YnMD/k218dSXntYjVDq/+kk0k5KPTjCoQsVe265EU
UQALsGAw7P0s6V9VX7Lo0Fre7QT3Qe06TialyROdzynDlx2ZAiRBlQiZmqcRAckJ
YqOwEFDxUR5MqLHOoUkXvQpVxkGILcPdGWyBaPrY6m5641HvXfPqx23wkA9Rq8cP
79G8QqWJ8z+Vx68K8xPjsUbZ21HAK8/RPvt04yWKuYFR7AR668p6rsDNWN/OHSB1
GUrvEZ1+H9GWeImlCZQBAArIYTYxJVgqMAgdsg6Fpa4FiAkNFUdVRNzXXJFin0mI
r+9nR4GElSUCJvBbF0gSw/f4Fg47qkwjMF/mqoe6SvOtPqqKHsxZqegrG0HYpzCL
KMKMnRiXBsTnZApNEPa0wSyD1kaHr+clYyHKkUoA6XyhRcjcImMoWSN2HZKRbm4Y
Dw/Nz1z39dQXNCrzDjXmgFUibZRd6HZahjYT7XGfq1X/IattAIoTxSENPecL4/v/
c74Prt0QMuXkkq8Sg+q1eLdcUyXGCSFcgpglvlWYpCHUOiPCOWckbGsL5ea83jtX
BtOM3UP2XFQ0f5GLqYjW6Mh7nhE+biaO85p3rf1al87BuwBNLpM1Htf9IyRlDIQn
7G8PfReDGxYDaGotrDk7NS/xm4QUDsSoa5L5ADGK5N1TBqNWp/qGmd8E9Uc0mYXN
q1kSXA1e4tcrN9CUFOWL7bBEEqqjHw8GHf6tZ8ZblrIl3lYESGechFRxHgKoAGjB
Twd2GvjaxFz/nD6WGdNoXEzREiI8+zM2jSPNqw8+mWO8YvLfcDMssWwWljJg3Hbe
f977zN6+t0sxSKIn1DLc0zqgHAdPuLDeGJVqOIhKNj1TS0JklraYC2N1Snw/eK71
/JgrfuQN/k32jwxRNB+lKrjM/E6hxet94l2DxiisMzo/sK9Gbz4XQ9vTrkYt/RZJ
wR8GwSDW4u7xQ4ghUGI7DVHZkr3UlHkw9Ey8ZkEwpwxRZtCRWRsscJ6Xgjz6tDYk
KWmsvcpzo6GzZ9pcInUCkAfxmrbIYPS5LDILiTw3CQ8cDWoiB0xsJcPrFc/tFbkd
pKWaZo4JF2bNwwu+GxBS1bKZ7LDObHtgopbS5m8P0nDvRT/0aSQ15o8ObDkw0X2O
Ft0MiShW0zaRit4VU+4HJXOjeVCacrv5Pez3hKVBgzZTlqCx9tsoGz35LwaGZOo5
DvEPQzkVF0enrOiSX4DL/LCHzXa8MrTBs2k6QeDAfBkQCJqAHwXV9suVzUWigX1j
y08vlCNGIbfZfmTQPfRBoJiXzNBdQKTH6bvQGhmiRS9+0W16/uBm2BI7iMNURF4I
po/ISfjIvVb7Uof41vqyEabJdMW0BGH/QOumtavDFXqSjwbrBeb/hwNfkKuAs/vH
pBSNj7sQU6qXmcWh+o+DjfxAfvC2gVC9RZbkThq1GZawIbwe872bHWDYJzhf+zXC
MN2ESLj7SCiJhedFvqOPPmFoFf6hMqsiWSzvn7G046lPieW0XjgMDvR6ELpMtJ8p
F/tgIejqdEkAaTmKQB6hgsBpSio1TdHeswOehm779fWgITSVN4wxYnFxpxe8bmAL
byAPzMNUOOgMN4r+I2v8yNRth883LJ0p44LpKaFrVpTlKnfBVJ/ng8OW7I6+iiIs
AiegjUBh00TeaoQriEklwZjPQqyiLif32855PP3/0IwKSJGJk3lxYQ4aw4KHmKK3
sWZHymwajBfw5JFG1kgyJbjBj6p/92EhYlw8rYXOBomk00rKYxP/XP+R7vAQpa/1
8qNizt5u0KUOD+S4AzobNJLcvyw09LIfFPm79YFpkFr95nu9+++cosqnNG2EOSMF
VqvTlE5ndxNYn14YmaFRji9nvTUqOYcxGz8UaGvuCk51ATB6cpLRPMD+x7GErG0r
eHUir2PY05u91u0xNHk77unadUUNNZfWaPI72pBzQH7vHMMJ1qN6TScJmCMjGB7o
7ax5Xt5wVOsyg5LjJh/0H8xwBv/BQU/HEQBPTKSwKmqUnBlFAPWqAnuh+8n8ZfNb
5l2nlv+PbmGotncYgxO1bhFSeCDgYpDxhbJ1r2yexUzMN4myyMSznj3ucxo+dq1c
EBL2lhiHdqmRfhaJV/2pEuDeDy2EcE3CAcFg3nqmhgOdYU1owpbmk8YZKlJ8lz76
7ZZpxHjVZOnBTbDQ3h2IG6gJfEoiXk5s7SYnLZlvVFGRI050VUNkaxxOHE2CLr3c
QTLiN7WzsmSFBgHF8ml/NwUaN0BTMLuCEfvxSBPm4H3KPEcrJ32Cp3lFNBPp1CTY
Eqt4sIuZUAUbFylSwi/mLEHTtknjpLMlNBUVWKH1YzY5h0V9ZgdMXHQBXUS8XdKs
i2VizpuLM8IBMvdC7CuzN5uYQ7ZtrbNR4vaZV2CJ1IlxYRK6ynsRD1mWIkx1NZYk
DZ8lgSl0xohPnF9Zul+sUVjpiM75Paos+dBzbGVEtD76BqV9ojtVla2b1sEwJGjM
LrP2S0TQhIOWNz1icM5/0azAeeDqCHBLnr5PT6zBA00hZAqzYJbyBriDerxbrBDm
IqjRnUQTFdyJHITvem+O95732VrbRTVgLWR4TQzls616XJu7WiZXZhwPY6rdwCx0
MbUSOIzV+5SeXHmTo0gKUYqygk+o83SWNt/ShGzGC+8MCc3pJV8tpiggQmjT42n3
iF3wtG4wg1VnxgPeMjvTET1wvpaMJSf0dh21+LmDwgiyO6xv53INjQ5EntCXoZhg
VwZ1bcL1M40W+REO9YMPdNRAfUVUiflzeGokrSDqtJyNlKFNa7CmytleGGbJGnP3
P9Mv6MsbJAIrSCJ2e3eG1bO4epgzHm8zHMaK811eWAFEbcNQgZ3tqncOetKEICEt
s8jrQh9hoMfXEFoWqvuYPhUwIiGQbJ84UBnOthDx9fMsgyZbtPIUNc9f1kxwmmby
3oJQ3CV2jlbeayvG718BPYobRpY+5tnfZQA8A0UxvNLVGAnD+kKJOS0gEzyrpMEu
d0CXPpBC/ntMeYcrhaLPSWaLhu1VFm17AZ65e51PcRHF2L9FnXCzM406Co8uEPuG
RZB3pb4GGcrGyFz8DweOUfY1ddyaEXMzpeivUt87NB74vsd0MaZ+bAEtY56MpuUZ
+BDKWBghW8b/0r6QI5eeIOo/lXYo7N63k+dRLCfDfE3OyNP6nBcGc9Mo4UGqh9Ux
8i+gkBSQouP+xfnloXBlQX+bUfI9BowgQ5NFMC8vqa6YhYL65LomKaWNXN5H387C
dgsbFXhW4sEMPFbnqu2Pnkxa7NWNtUN9aYVY9mj+O1PEeES2wj3SYn7PHOxgWGUQ
YZAt3nfho5DORjY318DJrG6qiBVglJBaRWtZwrcjujZZvTyG5oBvr5z8Ho3LsmTe
DtA8P4JT/K9BM5jx29AwLEH6FMGj9Jlcxbvh27gm4VUWG2q27LVGTBmyQHClMIsw
b9NahAIFFnEElR4mwfEa3H8F8LR7n1PJdneAFnfLyuUMl96iIij7I6Dw8rzF87w7
g2TX+KGDU3UHd/Qop3hsVOxok4WHrTMXFEYBga6lGiQjFqsvPPazKCCH88EFUfaz
wI9iOIVwER8XLy3X84YlBkzm20iIzeqe1NG5Xytf8/STdPVU8U5tEl0s7VIBX+HM
kv7rLUJ4vglMVF3MmBsl1a40H2hYYNA9PaSSthh3FggLL6WrLNoWLvbDmn7RC1yt
dXuuSJWqXy1/5q2OzjtS/PCf2aHpWvzbPgEf0nn5w0neFj89e9ZL0pU4iFLCvBJi
DecbpFKkLD3e4Ivl1gPpxUiUKBicfzdgqnE3Tu2KAv/sCsur3ZgYfSNghztK1Uz4
80Pi31QLZgYqK4rSm/CLYWL0IK8RpoddhX8dNR8lpjhplPAy5NmI+c5wTvOzdUNL
OJo2GFrnf8Iz8wXLR4wXMs6hDrG5fPDVRZRBLXcJ18VetMkGB/XyCi6WhMuY6mZw
IuV8SxCHPCUyP0P0FyimUgLnSgS7pC4mKfgXnT4gtcyGOpJ8bASIas2NFWS2xKEh
k5Mn+k5Sm5jJDXnISzADaN8x5KkH31AvTbAb7lUItnAQ4QRmCCWqqff4XHZcPg7a
cFl3WGVRDnoqXIJHu/muBxQgt6GSuknv7Ies6pNNVvTi9TM3ddzRd7HbbsrgjKpJ
OtVqy6/0ILRg3bgAnld01wokajSi4YUolca1n+1HrSNhwBJLzohQZU03+1RK9w5F
sG4gao8BuL0zw5QAwS1OsfIQ+wzYL7K9EOhqAW4F/oyvDtr8RzjGq+ZjwHfbSu6e
hGE0fcCgF03xcJT1RAaSJFQimJdByrYFFtuBtlwddX7USb6oQoxpBu4iR/bzZPTS
3PqgfDwD2lIxpf/1V3nVUx0q9sDybvAvJGFzs+jKhOJPTGWySrDLZN6GCZUpG50I
fMJT8jYRUYoOOrQQhjmEnFYpXwBH09CIlCollO+VkFcQCiFsGb2/REoncRwsfhxn
CQS7YskesYRy8m5m9tj+tFJ7YXMVjn8VAYVtpt0LcE06D/z7Wt6ErcbjsBybatIY
J++cl/FA/NfPpnWWRFz/QNOWSOKiqxXwylnaQ/RJQ/sDgSWMjMUGy+fpVkLCan8c
0jBehX0/B/IStuzN3ZjWRTgP6B3RQAlt12Ix9iLXS0G/i2gJLlSbYamMto+8Oswz
azzIsHYD4Eo6GGW2s8uddLyEkjX3KC4sx5FE/707QNLgoLWMgKwgCkcs8ZoefkgO
rqbE1bUC4tDMcOTVVpAz6rwxy5/BiB7e3Jf+bCeLAshqLhvFI3GjCaV0l1QJoaOv
xmV8/afnQmwS8/q7RhyacZu4dBJCSNYpo2JY1h83B2JC8xPiXXWuKyFZ9dtcdMAl
0cCqdU49Y+zjoirT7Vvvb4wZogd8F3O8Tmyp10xyC3JBG3qDhPkIEhP4Wdbm4sOa
V+E5SOTi66k/Ho3/9BZRSjqMvPT7NInhDoaw+rdmxJxG84O5z+1PPYDM47DwsPhw
n8EjUrftNE02LqD4WzkpcE2Ugx50wqLrCbqzJU2U73bLYRZXaBxX+1TxNuD6P/I8
waESHpffdnNBKzyDfDUhNrqa9691y41Qzsr4S4yZIStzPMp5JnD3sgpGiXLUhhwu
Vtd5QG0alHe0Op6i8iX4B/JyeQQzZuTtlsFEHxaxXAnaYJUjKqTg9F2ilZBSRHfG
7gTMWSw/X+JCwtSt7lIiADkqQQ+hNfa++iLaw9N5Oq24jfkeQ5sO3I2iVJ8eaW1j
L9+ykG9mgt168iteG9xR2vFt5wnbfKyKYFPzlkCSBhIHSzRLwTmQp+kIili9N4EN
RvDkcCA3FgQnj2cVphgYtxuw3wEJczN5mzbKlrbGxYJ+N0gVWoQqKzUkqDX4pZRn
X78THzx4Dbv2AsjIqCO3OHqKLpUNc8I0p8yUlet/anYBSPo07IwI5vxlWyU2Am3j
coFHCv+XaKqKp+GPKRJhTBTmWCw86boss2jDbjbt6QfGNE5YmlDOKFMYz9NEJd8U
11Inf+QFZWjqQxNHfISqOAyRb5v+QXTWbw7UcIA6Q0uo9AWPRNmPOjA1SUFd+7fs
OkMhjFt/MxNLMRWziLgsAkXrcP1tTwEJyr7KtSmfLFlNmvQYnabaR2k+ZeLfuKqN
+WPhYKkJG1KS1QLGLCM43B3XmR1vrRFUA5gRr/BXAtjOI5xBLOP37fmvTEUYe3Tl
NilTTYwrIPH/uaZsR8OvQrTjX8YIk4p9ckMoDaQbWY3ONoixdx4olIVB5jL0vree
Aez0S9QyNeVMtWL6r75j26mL5hJ1EclkC8axbsXsXiqSN4A0q8HdDN74mRSOSnjp
4TRI02oqVpJ8TCycsrEy5GW5hFJv+Vg2mrkGnpBmjqqGT0VombL+/4XCAu1EatWc
8cu696sNzZQ2XA0VpfUaUcLHOAL4c0sajg/Ow+cD6Zb1DlW4+UGAF1wdGQrtJO7L
Xe3y2l4Qw8xTB2MLE3LAK+f0mqaGlWWjbabOcKBsd+90Ir2RofnFmlMorlturfg7
oEz3l37s+YT1lRy0rW3ub3fTPqAEB1xjoasy25NkM777KdhboYX370W9pACRXVYc
KbD7chyFXKJbvVxGwhAPwsofFydipM0nEPC3/+pi8z4cH5GiJ4M3acunG4u+s5Mm
c/3PNCn3cc6VvIi9mEluwnf+dwkaXSwMgrul8IAieSkp/wHtylSuPeLVmfJkXZ3u
S4B+fnFyTSKUvw7X96p86qHPqiRqfRw4xOs1rigt7dumr1k6bAuImEr2wP3dQyaq
33LPKICbrLi4mRmJ9cHNLUpUYsoU/KZc8EmeWivKcYDElcYDwC7gwWn8Db9rTg36
XPktgEDgH8R8k+QNlspX0tuE4UYQ5afrUld4YzyrVuFdg0CB7puEzjKb7B5ekewn
Loc4Uqk9emNSJrQCu1sLgITRtkM5UAcqUP91zOYyYlZQTzuyumgRdhZdMHSklGmX
zBQdFbCrswiKnP1Ba4PvHtzCWWeVFdYHq9yjtanmBkyHCGZ7tWNgU9EdNZZj4JbK
u9Dj4lKZZvnvyVhOmfvbGYIx0K842NTdBBkFehFxhHU18Edqtv3qdrf3Oj7QpSuv
P6m9VX4dl0x9QmSvpUsgYAb+L0CXi4db4Hk5HhlcD51tE087bEqQwcBRhnURkagV
Zcai2EOCDmddY/KEUDmG8ZPxDKV03Phai1LK5OWyC+bxnjxsrRUf+d4WV6JyS4u4
FzSFKHJ3Vqptnx2rF3P025waIOot3dFxkhOtcAmJ9/LadW0jI4o+zpf0fEGKdaAk
4OnIFCcJtJoRgOfmmKzEnBfo7n+On03V+vkeZ8wAb7IBR/5QEdJVYpzTx66Ruidn
rpV/uuTWdfQeXnw6RaIa0TvT3RrIsWLjamMvYER6xxA8PcarfSRnYjsXpXoczXm9
pXHWIE1EXyueu7i+/EI9QPGM5xRK7yutDRtyTFGG3JSax1YeYExbZ71PlGb9bte3
FDMaNcReHbRsaX1dMzojCVI2L5DeQDQZO8tJlZyOCUl/vTsU/PxvxQiQGVQGM/Rr
LXbZ9jq8bUjgLvjjy7D7UOr9ZjMO92wdt9UJ5BREdXOj8pfrcToL83miohXiiOC0
DW8YJRuZlZMpbY3EcLEWI64jTmSwJxAAYimMCznf/stVGFd6DPfCHlITxd9LfA0y
MpxRo2aQwsnK2v1JlLFyUbdZZcK3s+o3gNxGVeO9y1A/+yq9Vs313/PFmJvvQXU3
pfN0X27L1VjiXgINokX1FULEuAwOQvxr4H1m97iuGDo1lsWTdSRtcVzdvFPr3S1y
BknMfLa1EZRmPXMHsNuj+kP9eEuPr1ZzLDBMLIcNWuZi35+rx2jpTUIQmHJ9ejfS
kz3RxFaGJ2wv/uqu132KnOzgYp1dlEeJqgfnMZriVpp477t4ds6yZFfvwYDnhAf7
cVXGTQyp8l+LOY8mvkP00Hq1N9R6aYD6K9brbtSF91MPng+DKndNiYk4Xm03BVOR
KGy6Np9H/mqm90N0yjNeOY6PP3ESiWdo6pOs6qsPDna9VkborLthYmSL7R3/Uy/e
B/Gmvlxb6+xnH4GXcqxVif6IJhjpW69aJv7qCFi1xocwiVIKnj+myzbGhHO0MmsE
miZ7YvEBksYr+0aKEHA6OKwyzXMHPR5Oo99AyKuDCuAzBHf3YANOLvsvnlFl99tW
pwl3RGe+RfznMaqJPG+KRBoimuly/BvjQtLQ4KkrKJsFYYW2NwSEBsVPtiJx5Ths
BZ9AqBwqvJyRZeGIUSfJvProOokuxzpylT4eCfJ3l8GfhkkQYjQcDe91DiDW9K0o
U4Gs50TNAxKZkZdVoCnxzcGfbGgFVDUGxBpAh6Dypki0J94O+11k0IW5sx8jSo0Z
CjJgYol60oGgoL6gAsbtHeRynLLzCkvYP0MebzVbjyxp3aHfyb/StJOIzc5bJXN9
XBS8G4eTbsyna6Hm3Ki940nzHpl7Dy1jZ+DOwv+vFSGMZozSrLiUMq+6rZGXfEO0
RYJFEVNXseKEwXoFuf/nbThzBvgL9q8d+SdmUeEA0RIZyX3DB7Y9PQ7QRjZgtGY2
cwyx8D+wG9i6feVPafrGmadwn/Hp2AAfZL3acB6ZDqYpw+5QRYmHO7j1yQkZU4Nz
hX5AWcvBG1QwBikWI3ENJfh4G8u7HuW8mcQd31l0y7SeRQys713ehSoELxyoRpdH
diHCy6fvcxLVgnvbjQiFwrulUYw3zMJi1U9+vDuEYh6zV8GRgrD3y2Y9QsqfD5IX
P9M/viF9CRk/cSWlmRdfinZGnaBzjKTNv88Zd10tjSaESioHiPIJBQTRhsbnLaBE
BJg3fCxwoWpipULuMlocR+H/xcIhWRx9qnMly6PDqzu2dujw7tknqexariXFA3St
9y1u1V5Ht5joMzdldJvqyXzhy9WE/Mtw5f4hLhZyXqP36qwyJHD5UVwB7lzTOsm5
jhx9JgRNI2gChfhxfTCFfYJhRtGD5agm+bSVE+xOoWrDWR7ExLBzycwPhUo7gfYu
t/OvpK+Gb1OF54+YLeqLXZcJpC6yb8Z/dkI7RDN+f5gtetxAcVCx0tmA5gbGV4fP
hgT9fAPrJoWPtqwBQ2KtVw+d1Kse7vytlRD9WqyExVLtxabdkQTbEUTBWDMRrvzL
foAMK0hioRioi7TdGOnD0+oG6gc+9E2c8znh5iaSSVDdmjsMFqxrlVGcFCC4yY51
fOkM8C56h6SsABbG03DwIpomcamNSfkzUyjVmceuXE4BO23S2LmMAzqlls5jgV8f
sVfO89XnTUcMiq8Hy6jRnhcujJf0PWMoBEUnQ4kL1bwIVdkN0iYSpDEbAwjY7rNz
eKqNnjxJOnSP8vEFfYfacn+vs33mMRsTSFuYY0tCtY9Ed1AkM+iWvBOz/xTVj7Jh
kpk3LNMuh+wURmOrWEKcPIb6x/rPop1LmD7tPA0tWZkSRX65dNkxXVg8rwUtWPp4
HeM3LeQyF1mN4SH3cZtPdm9873V5tBDle/+Ddjv7CIr0kkrTJylFjnsaLMe/39cM
WNVcSiqpmmXQtbarr4nDnTBPTVflB+1WPhXyT8Ea4hGCNmd1hnKhlWnCio+rJZGI
oI1e0f98R/HnNa2CsIB7LVukopnwAH8vQxXi2pjd3ISIVWq6xyOYvAEwu2Y+ofsT
FuM263cq1WhtHwlIDv6pU+4Gz1VfJSfDYI6ShedwLggCalZY1yQrfWeRvyi400Hj
l0+dOsZYD+iETeNZmLe9NLmmX+0KK+P6TriioxI2BrS0Cf9Uel15sgpuJ1ZEs/p/
mmED7QlMHHuj170/LhXlz+cx+tdgmHwp7QGxjIHz6oqTr0ig6vejEEv3D4FGOwAQ
m7j04s+1jW8CeOzV1Cxs3wkUqv38kp0RK5CVV8QozGCEaLTOK5yUL+4KQWtHppa0
LP+ouQwOSAAUVsEe1MhPZdtQ6HMp3OADsUI7cFET7H/Q+hJABnPvVjUOBgGJ4FIK
GOXWgejPh/YwJ40cD/ce04UHz79XDiZpZMGY4Mul1oy+TFl83OXwzMwFuQVRc4ER
tCxeyJnLthvUFCZtqXnWWkGtu5ZhVA3fnZSkH7hyQxJjR5V9Ndpdxi0QLWThalQz
3s9PC4sbD0Ynq6imbW6JUaZdyv5d4SPOiXnDOK3dUC8Q8Oohx+yYswzkQMXRnEsu
rXB9gCOUc7FKb3s2XU6P96DJJzYvQu9bZ6Bp18HjsgmkcZHOKbkPYl/WoszHo45c
6XmHdLHj5uNta3dfn+vFPI/ttOCMhuIpBwtM5kudE8i8oVIC+XjVa16wVIYNfIG9
Oc0htu3LdEWmY2ikcUVGSBt7b6uH/p35OSKbehIF1642dKnjIaN7SCEYwHx9yC5q
ak1y+EiriuP4QwRu+Y+9v5KHdIhwnZRP0j45dHvFaAUV6GwA3qGGsxE3GGkBRdG6
9JKv4JHNe77Aqy9SL4UDhXbwcp2b0Sw6mLsMtoE6bXOTOgkJDW5z0wf8f3tqCTqd
tpHu497U7zPnzBDzif0LY2EfsvRRdbdyactJ6ewiG9b3FfvZMwx9CG/icAliT/ox
+mZ+pgquA0yvR2x3KLRvSaogMRkzJbYjKhJdotSD5NF8hls3D/+v98DjfFJ4UhmY
DOyTITo8gIe4UeWOk8YyKlcWOh3Pyaeed2CE1J6RoCwmCFkbyFHPNqXHMSKw3AoJ
rdq7Y6vdrDxcFLYWhzvwNCgQbVYZbPkAcJGVVbiw811l8YXtAzU4Df8b/K6pHFay
bOKskH5605a/mJL7+nwpGghoxzsZqZXpOPsU2bqs2inXMC6VTfTCOwgMp8s4meOM
DuVxI2vsxGE7X4Hi5ccMqY/54xISvLDNVV4X37F+iLxyWe0+qYxOScoFgJc/0rww
r/XnmvyJ65Hr/rFJpihMLokeCBXEyXDWaivaQUQQF/5NdsWZ0oSCToBj5292qN/P
YhU8B1y3wSROFzHT1jweubl5qnu+83l/04NUXdCpCP6+NBsAWFDBqtmqYzlAIVf5
ggM2ZhSbc3ecD6Ojre34oN17o2xxsOiCh2LtB0r2Jdun1W+VcgHYCnFYiTtHBtBi
ocDNc5gTy8cybOqfwhM+ol0v/c98sc+++xIBA0UWjFs1TZZpB27ahc0fFUJ0wXrk
8FYp7yTGCrid4rkSqNYwKzq1iOLT2NrJ5XHoVE1GUgaOLu1VgBP0+ABG/3KRrkTR
3VKeVPCY9eKpccV8kg2YQ6SfG3s5vWYIOqedRYkp1bmXmooCtREHQK5Qg/UZLn8i
RZb8zq0PRhbqqG6tejAmOVnRJucl4JdPoNp3WUieTW8Byp0f4MlJqGSISFNReptC
z3zW0B+hlFrjichfPtVdGIU1TOA29mzOo/iCKa0xaGi0tVQ1FvnqddW5yt1g8Ze/
XEEM28y/Rz9Q+nytMRCAFjIn82Wzr2YCxNQChzD8Kx47B81GnhIbafFC4iqW8xMh
Avr4/xPSlaDmh7yFukwxfdcY769KoyLfIXK3NaCjUmhPUJk9tOP2VoBFzvpQ/Wcz
jn7MUssyfdp/0fHvc4fr7BAu3kYKtu0G9xkCqdMSy1aMOkV9bV2i9s8Fpakg0/lY
W2GgbRgJE+fjbHVaZRPtgYH7X3e7oo+aEn0bnOi8fOBbN0evIRpR0Lmw76+nDz0t
QKMqs9gYwpUA+Ew9lLDHTV+Y5gfXqgoLpQdMb8dBWu5EbR5CSttsvJ0bd0njPbmQ
lA4eP4of/UgVH18qV2ThUCl82VAl+x5/us5DC+v9v8hC+6l72NjnIl8ZJVg9DTIA
ilSsrJFGn2VuyBfbwqwVaQ5K12zGeySf3SYG/6VByKCpGnSef3xi+FzwHZj/B2bl
VyFfjF6BWiVBG6bb1cOaSJ2UVqu2Fjqn2IjTTNEbtgW/rwV3VqW0oqcgiXg3mvBy
N3BeTqUILhXHsrs6SuC4kwPOddrB0qXBYdZ22JDBUbPQ7xCFU9xhSapTLr8+xJF2
B0XXSrfXNjqvuovJAp3tZIrS8+M4njMPKrEJYfGcSUTYzReb1Isj4/2Elao7lqnz
d+KpZidX1YWA6mS0f65ChwLQDm5esiPPBhJxH/jiyDw47Z3RAPOOrDL0SQmOHeuO
R1GmhJsEdG3PVStb7GXA5Bm6mivGMKfyhwxdwk1HMHN7Bb3XSvZiIF9Bt5UCX2B0
M7jB27wDP+Rw48QCsYbabP/kFyVcwaf8w2ezKGUa/oT3mIrSCW3Z9T8u3RQ+1M/s
n+Ni0PUXtjeChbYKM4bzkluvi68awhS7Zt/TOK3FoETb50xnMHVpQ4IF5MNCzm+S
OAB4mUAFwSW9N1+CKHEvya/g3Wf413gjVZzFxoxzKMDtUt/R7nIrrE2eV9l/uIYD
acMaKbg5umBSPl2XtGXHEdAIfInbFt/jpmJLX4TuCbNsNonEIb7kPkT31LO56Rjz
ftIjNGGWAyd0jf5QjEE6vDzTzzmmooBOPCgz015jwziqwHY5BP25qqfizndglF3w
rIaZE7mNR4T5kyXIt2M/kSR8oRpUBm/wpXVEmwML7mkewvSpqqkz6NUCXpM8PJOz
DxYCz3LhI5CU9Vl1je0AkPMf/Rd2jTYzQn9DvsykJ34p8JEglaqFdEDEcbM0yQWF
cUfxX1im9MG3vuTysurQdTQ/3lAzt9p9+CDpUAq5mFgw2BQ83Z4k3BtZ6Nulfl4f
3Tj9X5r8vE180QHcaDcxDdEfUlJGOzhGdTYL5p4lermCHZHOttiB1I6SopUkTG3y
0dGkc4WMMu7uh+TI4+9wOkK/j1fFpgqWd3lukpGiCmn1lV6od2RMSSXKIbiIj68w
lor/vP84E3ij3i7T4cC3V0k/b4j31dMhck+Rx2EwqxPk6sw2/Bv3+jwFE06QApND
slJnAONYlUnT1YWK/ANrc5CN6YaQxLe9D8a1KwEbunrnrFa2Dnkht3lUApihowr3
i5dGBgY/GaydKLckVz9RSkC5kSceXeRy1x8zO/X1qq1ogOLiwm01vFrNA7NogQk2
K6MLWp/t4PiDrYVdY+qRSJO3D4rHy4Cqqa3+v9vVsf5K50v01HXQKc1e9q/QoWzL
YHVdilXTMwS+WZo4stoStB4U04ovWWj88QbAuAClhbyoWPdIDuAw0700XYV2NSph
2qn6MVeqyr4s37v2KTuOSxgc69eyHhJYQ3Rv9zpNbiAgLCLQrIJSYYUrIj8M/bMx
uVsMm3fhrbau4SO2kaAC+oZLm5/i8CaxsBYeY9NGByjpkoCI/KfyZVl7ExTJYItb
bZq3FaYuNlYHDWr/UN+sHuVsHQot/lgsE1jgkOwMWAU0Og8Ss6+miArJayqMxbUW
gjVMTEphrZ1y/yvchQ/fJPvbg2NMvOHwuYP5FjZmsUJaVDh+pUIllEUpmPQP4puV
TvlvlyqKstYJYBXW+R54xomJDFLIVvjXg1BTn4XRUCIlZsDllnv5rQp5fD8Su4q7
7utD/BmvAPhilznVMFVO9mBQByCg9LgelLKzm/Uf87CS8gLEr9SWjrdXsaMNYvWB
/ZK1NMdLrlXY81ure6NdRHQx5c5QPHNIvCmOtCIrhLtSc8Sq83rl/qwRXHZ4QCOg
uVGeVh3FYT53Qkq6+UgKewjm25DDf/sq7gxAbuE0UQ86bOJh43i/plfqSztmVVLR
4X9V+Ntp7pC/KEdLa+O7+rurudCJQ9+cvNMy83/cJxFbVExfZp3Ja2GoRRvO2M8g
lVOmcKDFe2U95BQfiJrntgbR0A8JaykzgQQWflUJa9CGqiZt9EcBesw9k1yTgxXB
ePBFBxPbi/3t2wclqh4yoi0ep4yaBqVa8iPiJntJYlZHWGTaPeb9bD54lew5OxT0
XywAzq0in45zPXK2TDvO2+LVjGBpZRWBQuM6ojhOlTdqEaiOf6NDHEqvj/o8EOit
NtkY/g8gT9G4nN0ptrUo03r2gnCPMiTe2pDghrhBmUhEb9ACOZog3Xerp69AiqiN
uXkqS1ROcnRuEvWUy8bqNSCk8PWi2E6fRsP9ZFYzM3MKB2TLpJdn/rqFFUOqmsx2
VNcFoJ70Uxut08EgfbHV7TJNLVywIcTBxkbhoMLstjol9Kt9kRW+HxIo5jK/uktx
ACK49/zL99ti8OiQBlH53DSZ94sS7QFzaO5dSplB4m/B9QHzRsVpPNhYJraZKHTa
3HuZR1gQ6dQV2au1t1MaT0jpGTdxsRP5Fr3yPB/GEclEqgVgIMTuG3QNH+foW+zx
nXPiZvqCg5CPWKsVnBk5do2XKSc8A1ZuhTWa+wC77O9ggAqCXPkJatfq2bU70tSc
J7kchVJA+1QtucnJGTVyqsQEfeYVoJWAsgdrT3m0AV4xmMtPDPEDYvlLSJADNnHo
PTaptiaJqNXSHtFhdQhl9oD+RsPrzMw5ao6YHSDSYv2HtNlN5MVK61LQk0oybbyM
frDaOpianM1ZbNQOjOgZ8OPFFWy85rpz4WoKmqTsRaHl6xlb0H37LTqESt5Pq8pc
2YgGydxpa6QYt1e++nlAYegaOIEAFd4yNkdAQvX3WJJEQf7G2r4DNPa6Uv1e0r/V
ablvGA0y0irmzlHMDMOkEPu33ngTd1HB19cO7yGqq9cUaHkL0uDzw0GlCD9Tvqre
uMPdcWQp4h7qHY6YeAsv4dYxNgJjP33ub2+uEup0Hrv2VyBsfKbzpTHEdxXMqVbM
huTuw4MchccLJxW90tSfWAg1M2bYWUzEM1rcFjcbo6Pho8/G7GzVuMHAqUClmfuT
ynlv1ZDr9UQC0lvNlRf7nf82bwKsw+8ROOdHXWKbyh5prpsS9BtB7K+kzc68Lkqw
9csSNOshDDdwj8CS1CKYhcXUna5Lp4tzAn53zD0p24h0FwhEP9vKypJvgxT3YHJ1
Z5v5Fk4K1fb4+fQ5XVll7iNkM8k5tEyGtOpT6hS9hVyZbbPX5+Gks4ENmIJ8eYmJ
ctfbJs/BSUJMDCkQMLyD33z2uu0sqn8/g2J5WU+s7iBX8EVdKegKwT60AbnZZaZK
GM/tFDlwd5PTncLUOsgZSgobo1Oqu0QTbyf4qGdZfJ5eoyU9QUg9mQrLPEyAEPRl
mBPRTWHaRftoRgp17YduGHOiB3eET5i6NaxF+RnQw7KYlbe/atoEUn4tq3xvcvfC
ZrT2YYoDoRgylq8Wv38/Vf3L991MRWhZRPdTUhH+h/Jc53X54IHkkYyZxHThigWv
sOEXjDBuGck/I6KHw8L3rIhQiIDOkJMREzFcGnxBoXCfPfAolMqKTn0IUAFhjBiY
GhiYj8w8ioLh/uT2gULrxY5PvCsRX1rPaQZ9r+csZvfk2HCw34lfeb9wp/8BCGck
428rBXn9/T9vJ7Dw/nSy6QDr/h39C4mqtImlOSaWFGqEuQ0ko9i+1riCZ2pfexpw
8sciWvD4qaqbVdUUp5EU90fvK9AjUvml387xnPNkUZkZzW1Buhr4rIgt3Bi28Flt
M6tujjM9TyGc5+ZAPTm956IU8WoXjlNN8t5lS0VrdmReQJ+p20CWHQxODpkOLMHm
iSdG12Jca32WXD5HfjhEYseg2KI/McUwPePPYrf1gTNUAT3eeO+CDYrmb6i/UsAK
6aLoZ0okncP1g77igVbT9LAr/BNIq8joME9ukiJwNYUt3EB9ufwb2PyyOJtWL7cD
n1mhHIbd/y/sAAZ5DlMbA47glJQgqaJ8qS8KY8pUjmhlJhUI8CbvsTPjil6aF1nz
wivR8YA6qbAIbhVPbfiv1/Y2nfaBtW8M6d0Mc2N6A9K3VQIgmZ5SDBB/3eem0uTl
EWykcYXZBbEYr+rYbsv0qkRd2Nn/4nPmVZF9Z99hVxlsxHG4vjhcYNoEDQXcmZtj
50DtqSwC7kGolJXMPIP6b9FpSxDa6Qpsg5+qe8wE/aJGKXzgNNFmE9ydB5czJi+q
hiN/uIZlA0rvFZHvjn/mxrc70eDiGhfRlDberD+goV2/M3S5h2PF/txs9ZmkmzEl
VUsc3BfrEUu7qEAP6yrVVoncMOcNofpOuYpB+RzGxQtpdpfyc40/d/w8yyrcm8ny
AprOH0GVEZl0fyoS6OCblwoWKCkFtevVJtinEJXaZI4pS1aFlkY+yuvfC64t/bIy
2V2BJq5uohHRni3sFiIdxOsWxjmPIGhaz7CnK83STCfebnXdegfFe9zK3pNSGMdG
v26m8RqSdzv4wmU3IjcuZZaq8Cf7oLF16z7R6GejuQy3sfdPHq+VkSlXa0o/0dP/
NhukTWXKnXgbOp1hWOvyIxocef2w9O7rjDR6hyTVXr2UpnYALzdr3mh7xClCtyrX
f9DlwgT9pbgwHnt6aQzpB/LubBOPMUcfNs/87snkQAlnuGfJ4anuaKPuxh07760B
yArRTFqFRfyjaMQulFeZLgXi5Eq9pXcq6w3o3R2qguWoMZ1ZO5oVPEPlga5OThaf
HN4jWKh7keVwil4HdVwIcoWG6bYMvSOhUTWVstP3ITqspUALvgH5J2tfUX7jpgJR
6ftDytpwd94KtrhvHO7TBfzyjReHuG4J7m1LFbri0FnIv/GAWyvnZruwCt0lVdX7
qCl/CqDVcJ/+qZhnwTiJirS2Q8VFIFEYqE2xKemtfYCT8Nvs7NFILDxKzuzk3I5/
IDrCKNnQCebJpu8Q7mtRrkHDtbd5pljpGd2Am4fhstah2+DsQVTZPna4f0Q6Mh8T
uotvgZZfJBjyhAdmfDeIXLh8LV/0RBRGQIdqatHIdP02ewSqL7X2RiPolvMSj6W6
cq6cWBPptDdedk1CYin+gSRPcMy8eI0TX7EtWoFXn9l476xmzfnjhzIX12VWYnMj
wPXgxbd94r6U1KdUxJ1MT/zt194eJWjkuaDfjqkoEFmoEZggXOCGd5ZWBVKUXzVg
xu8NpmM7koraaXfZEAw6UThYI0fKxc6SaVvXC9/1q561RRTJwD5INsaFIJUWQxRQ
aJrhulfliyI61mlv+Xl0mi2Diptodgteb6lavaGbSeOTG/XFi7WhftVdFgg8Ug06
+pyOtvfATQZa0ZerpgdPrcBk5K83oRH5m8o9h65I94NHeVBL3W34pTOrj2XJbxAF
EbRu9unJazw3tbatMmBTDaMvwRtP4vnC/QkSqJ1ywS3HC6j3Jebq4BNR9Z5wQPK0
Qy1QkCAsLwmGUiZWgHwn9gk8jVih5wEqUoC4Jmh0HaB87xSNkd+fhGBKw+069MDf
vCU7fbKq5TwtHTK9wW1lbMws2dOQUYM/L+WGcxVAOuOOKPC0O3iw6YY63Bykrc7Z
A5CAFk7GHyYs6HrW16Kflz1JnZKbJssd66Ecy01pSIo36blT3/FvwrZL71t2wVEw
tx3mUqL3XAA24SSoLeYQ0ycK6O/bpiz8uEcrub3ajUtRc808GJ22XrNOaj5vCIRE
+k33Qb201Vjm/hKkcCJBls3tLC0FIzzSk2O+sdmL9rhK6+P8xt8XH7IUPo6xR/Zy
n23GALgdFzLhQp3emb1K2r8wf64tRMn7oCB6YC4f71GNxk7G9qB1tjk5e+xLk0OK
ufJrGhEV4vVFya9CZLRNrK3Fk2E0na93rpQjAZI6AyUVMzDAeyrX9GAwPh/RLwq8
W6pcm3kSba5Wi1TkwwoKYoMDBd6DlEC6reMv8tjiBBB4va3j0IuaMQJFgOiK9j81
iuCFyfUyfEWmZygDfL8tV2qCQZaCdqURKdrpALmrJcZJyDs9xTgBAbI+e6Rd/anf
nen6nukJQOkv3g1orr7NCWAayhGDm7P4hYk4aajCMe/iIRl4tmoBH33+Wg9btc3o
+1Mt5zehuOHDONZHAmCWHJROXALK9KA3dv5ozjAXZs0tg/jKxNWMRDysEPOhzrER
T/wWIxkIDlp/2sKORYL/vrxtXhuxuJa016murbuzBv+j6KyAxF7ZNuDkuvan/fWA
e/TnmvuHov8uvQ9Q0iagXyegqx+YL9Jm2qMyn6lp0//DIXiYpsYd9ra+/SnxtLaL
hXsOGnmB65BzTzqpWngzVP+OaNrgheex4a9WeWLSSWYKZabdPI+DHBig699q+sCx
EysfzXVPHzwO8WlMlMbD5jgDJ0EdBcNc5aZ3wUsTZRiBIS4iNpbNlrx+ItzeHawV
4qRulmlrj0jhLhe0OwpNm9rAc3YiXlH3tSSikgvsl+Tmfzz5QizaXXr62i/3HGnP
Rx7Kp47KHhUrIIVWQEmk3fzbb1rdC6TIgFxqosAP+Cg60gLeGJjMbL7XOH6upcUt
sJ0PRwoR+iCuKS/9rx64Lb9gLZjLkXkJdFJFYrifF1fJBqM5ICAyKy3eH6qv/kbf
p5EFX05+FX3AQDXiT5of87N3wdvS8OjHvQVUtrkjLKvPVs4lzpVDTwvjSJFSl8iv
zutWwRkUQ91Ud4y5IA+L9btsQYyU+aGb0glNnS6Of1I+f5wPwP9ipEj9oJJDNOF6
XyFRBd8rhfV/TJYqmWwlsCslJ+c5eas9femaXvhNaZ6yilHHjpMfGodMqpAY1FRn
x6DeZ/zDN+/6z8RAqgN7YdrH+H976PJhg/l/Kqx1mr1EKeaNCBT+GIc/L1TiqdHZ
zKoTXHjepk59yCYPh9n5g2u0sHpPasp700kZy3Y4CLXK8ejzhlXkZVjpMhuv37kS
wvuT9ZyESyijufRaSmCbsBKALoETeDf3N/fDNo6j7KnOylLrNxmJgdfx94ey7cNr
+q7TgBoV+LqEnIGQezQhVc3hmtd3FSxBwgNBlNRSotNUr1L3CwYPFsDRa9YQTVg4
fYHcgKBMh1QCInNiqi17Ubq9cJQTh7g+L87EgsLeB5bvIj0jHKJcRyuKHKVLRSC8
uvT33J79c4QUGdel1NR/aWmiN2/P+oXT3lUIGn+8gnFNVVvbXfGQ4+6hih5RRuoa
kBWeUIz16Xub6Q9Ts3OqBqwzcZJUwDSOQ7skP7uKlMhmHTrhASIm8ABk/wcdeGNA
GcFrGFRRb6pv7mdm4ycwk4iDlOmqCzBOZrDOQ31cuRBZThC+vd5yX/PezfXqUwQo
0eJgEP1P+YwI5+zQRXaCSc3r+ylgUAzemFVxZkKRjFfltSk2+Zo6m8xa8DSFe1+h
jLtNDV1tn7bD3XZatsB3LM8nDzlGDHlpBEomjKm3AtpuPbdyK6prMzkKyrwo5Klb
Z52FtjIXH6q0K04eNg18ByqEhng612KHXr3DubUaXqPkLpJ3S8pOc4NiufwPNxCU
ey2fCsqagskLJhVkNDmpcQHz0oegvZoI914m66zr7fifVVr+SAXV0w6zvpDDF3h7
YVGU1wV5sXW7Z4/ZYMyfQ8DZ6emQRdFMc+2ZFdgusqUBcrVYAn3ub2VipkO17XtE
SAroMVAa1Ofeu9Ae0M6RZ8Bu0Mepi4PGib2M5YpCox9KuL2DtvbIHF6GtdNFuthv
n5msxtI08CUHBNvurOh45kFQNV7pmINigr12JfC8JxQ7dzxW+YgS6BA73Q3/eBqs
wgghbrpyNkTSCkCDG9eqCw7G9Q4VngTmv1zy/VLXQCbIIqBWoo2nYW0J1ldBG9n+
KOGSpONZlNhAXinb9rQ0AVF5gDt/cBmgk86Vw46IaqK5IPFuHUoYCrtTdG6oI1r5
NJySBW/4EOTGYozfT3cP63pyxKzxQ9VpnK1bvyTTfJw6lcg78lTVjq4jxC1y/WDA
rXsitQFVhE5GydjdkG6NWJwKdiUEepuMnOQxWoR1zzRMs4wSMKIa8OG5NgPuD5Qu
Ybk0oGYk6LRrlTbHfbwNug5VmDqs2tVkOV6SFThqN2QSffVdKbeb4UHYCSR+cOZt
FJrgBmLM4sab2yGx9qDC/XjCHLrBdZo4zn2MemNWXAuNWHajAe/yZQDqT4oT9DqK
yNDoGUvWoRoxbdLAFUNT08pcbdT9rAszCQbDXf5LIhiroFONl0u47XuzGpjkeoR0
/vgpe74iJ1iGY5A7YiCrL+SlIZcco7QMH3cdtPMVdGbq5uwUXbn+wgbVhvBX/Cku
DmojUHwhho6Q3GwqCBjz6kLhssJUYtYz35ayQ2rr3CplSCKVOYmxJeRS8x3AGs4j
hChle3F+lHIZ7TlB/7hMTWTb8wuQ/fEPbxdXqjKX/2zbeoOKwmYuR3egBOMSQpD2
s4PWp2vdWL9gFaagJ9pHi7crd3UWQZvN37zs8kGqclX9XUz1lsSIHqck+QOv3reU
h8jIPqZ6e9glPjar/aMRQjB4+t8WOUnBcsziBo7oVrLT0f74HGOnZzcodyDc2DEs
yAOVJyBPYdMrMNIMeRjmim4CtZRMd0w/WU8zQZ+54rUHsIZsyXK4l3d+tNDSalng
LjZ3VxbKegMzwmxKGGt2KwJ1sj58YBUFpATB+taYOrrsPV0RMscpc4q+dc6XM2nU
m1ishFIrtuAV/lDQXf4Tq8zN2E7jSnMSX63BVAzwW/avb2x5GJVeag6SyGh3bUyL
t+DW6FVI6rEkDZYZem+b6ptbRfd0mz2BjAVxbfQirZK98J8T5axP0684hab8tbEg
hPSqnwk1Cdrv8zya/0MreRlU/wxunNgOYKMKrvo67MWxnmgkx7D4ME/2uyb+l5x5
fCEe+mfWPa9mJkPjw0ibsP7fB4I438w67S/nisxsMY6FK7w13nSCfq0I5DR1qcOw
EnCxpwEMRu38s5Cy8f/0EHws6yAdKqyK9+eCP8zf22qv+OgXbG4q/4KM7WdPKk/r
3nZbG2hOlF6VJumlCCO8P8c7+FJuF4sv7Q8nERtmePdp0g5U2oOV+m/hARa6fNAC
ulWJpC2H8DEK+BstvP+AcWIrJcAZIN8I7mXXfNPe7vYDUSNLzEUC0pd8CS04V+JD
LOAgz2U7/khTjWw+3n4yOlG9LLvqtFChe6D9ZApsZyg3j6ITWD828eCHNXXxETXn
Cuu7v9M4G9jw2xYooZ0dabZH/h6lykU9RaBv73QY9ghiEmAEnG+EHkqemzk4xUKY
xMet80RmqClplVPjxvwi3kb22LtDCkvc5+IwrpV7Zz5TVU41UPm4/PecaJxSKR1w
E7q/J8UL1OOyIe7Iq9cBA2UmCpeZtk7fwY3KrVz6QEtf0xHlSSsNWythsNW4oXhC
BYxIUkcvdU+gGE8J7rhKXQZgvWYK+8xOgf1OIQqagy9CvVB9GUoBi3OcQoJO9Ene
2vCAVOnU+f1uq3+Jr0ZqoadFOegzuzmW2dURmHpVaFdS1F7iJmZCgJ75UVRw1GzX
okPuxlsad9RstQu8HVD8v0ErE6xgfX6dCCwrYuKmGJpAyBgCa+6BznYOSjImWIk1
1Cw9mqrY2G2/1S+9vqHrOuZRZcj2Ef0LglkN2EOIuZY2SBYChoZWpRCogkgEjcT+
P7LZpvPMw1DZ8jPjIVN8jvxPNhD5q6JbDObaGyDwaF2YbCGh4+wZwh25B3vh0JJ7
hohz0G2RRhAAuXPyU9gNANO/6o6f6R8Jjdpd5W3ixOyg/u/2Jszqq14I9A9prVNQ
3+mXP1wrPPj3bSGlrs/YwpwqrSusJajTXHMNzzSUci06pWWwyRCPynT3vSZl+qIi
QnRH9LwVbNoXdtpBD7a5sQEEAGVrA/SneaFZRJPzO4tg3w96stE74LkB0TDkJyb2
J1nY9vXPT7w73UYqkG/YpbVwafJBzY1IKr4SNpEwaosIngop9bbuLsalSJbL2ug5
zOT3V5M5edoAeEREtSDeP8As60GJ1duOGH7PZQJgt45VqgObpka9m2PWQy2Plge4
qpGi15rRpRe5aq6DDunLNd2dlPY1dUiwJpag/vawrIL5qUcURAr0AoG6+LJ/C4yt
8Tkj1mRUQ0rnKTtGBC5CiKQ7WvX3qlVC3LqLUK7o5JrB/BtRexN5eq8jWdkYho5c
PI08XH15ZArnxO1IFXLp8WDJ8EbPHW0LJJNIl2WuhLrRiJoChxMt6SuKmdF8YTaJ
B5fNy+ox88/WlD27MDPPWstVOeGraRWNrF6lm1z2SQihxJLYsFKrUIgBIUfwPJbD
+zt2XKjqq32Jwhzj+9epeZxSARiIyVCG9eWh1KpgqKqeHehLMnyFi3SSJ3oVPUfM
BiTxgcN3mQHWUYd5Q/n0tKVeSsLK/vqcykZ/Adqub+giGRDwoIejSzO5kF+CCiC4
5NCSvoZDLEJroF5p+tYY2Xak5z2E+rdNKDAlmvpXH7OE3m9Mw4twTokXeqVtElkL
Yt3FugMTB9nMzdjW6AI4ooYLlS3Sa0OWFuR4oKliFmCGiKfEXl9ujx8qpyJlx97W
I286wd5zeRwC8/YgnXifUfrs7x63rVqshJgl0Xu3DjpAqFD8Fun3cX6+yK7hF5Cp
iyqlFwK8tWQj4OcV9QRgU76G++AUravP7Ouq1YFoxQupD3w3+TNNChLF+M+/M3Dn
zGNHuv9AR23s7X3blhi4cHveq/V+SjnHU3If1ASI46jC8bPaEawdKclsSzTckJ09
QTSQPGuhGW+Dm/08jlEacnvha3ZfKH9Bb16a+rxWD7xXDLvr+asHC5z+wzYQD5LF
/JKe415BKXZQ4asVui/QymZ/wH+eD/1dr0miP+kTX+RTILRJ3VVO/iIh7X/tRMKW
x+8ouVgx3CPIqtd5vdpVAwQy/AOW0jebDWsbtP92LFHNmR3pknanQZNmnI6rZ42g
j0MCMFoywzTyN9+qxCfWqZEGYa6DQ7U5jfybS3r+8GzOXeT0qOjCTg1vopdoZp2L
cl+UgjVFx3tHTiR6LzlEtCaFFmwXxC96E4+gNGUSuEDSlwoaQoA21h20juK2T7tf
TmSsCfQu1fOEeYPGgr5eaZFlzhDW6u5zasLGSGEi721YBfbROEIWBDpfSgnvd9me
CHUEH9wgTEVAkin7rVmWoi+hSa4daZX1cTuR7rAf0AzqTUJGioCq3Qz5OuwK+Mgc
en7iadkemETnTEs6SnW2kIuSDl/janZ7uiHjmOwLqB4asGm9QUkCZqVi7DVMqcjs
/N5k6kVgGe5/pgnmglrWrapLz3+dqa6rWgrKKlweM86UHSxs3uWD2dW/yhKi/dYk
A29wxa/rokdNspVdJqeTqLrDNteEPbYbcD9YmlAur5kkP22jnCgc7gPOMKUx2gNO
Ze5L94rJLM84a8sHNWV2r5mvjXjMo9LzvHBHNPSnzB+5Epqbs3q1KvEEjWEbaSQz
+oVyI7WgpNCfwJ83i+wyLQGEfZozt8XFS43ApWMCP+16YBgH7nmb+0bAZggwgSH7
YKfNQsaWjmXISGrPK7QqjkfnAKRV7clRrnRzL4uWzuo1fmSR5TMIe1FaxAvfS5fj
JyaCBZ7DGeMaTNqf8A6utOO21WepSiioYouA/neMjckpjk8QdBgTKQ5Ff9k+FwJR
mi+AhvAqtVFSgRdr17AINpLS63F45Pfw+7KEki3GaiulE0jVHXbwsTJqzwqdyeo/
tJUbRM4SIX34JEyHBgD29W4p+7yo+23fcda2XAr0VriFFKNzKla61w4ki1E/CgQL
L8ZpS3Ru1K74kfxX+EAsQFXzDlW9gjLRxqSEE8bDnmVm8FRFs7L8ole41R99FmXI
jVei9XP5CDVRH9+aXlyKUt4Den/fDpF4u45Jo8LCw85Q26Gl+cb72x3CofXOX+mc
K5Mjpy+6lSF3ta/OesrGNNN+qTqvpEXgBeyvRzaPyArgWmpKGauqAwprP7JKqtuO
2Mpcp2y0nzDUMSJt1eDGXg47AXaGFkWdn1PCZmmaiqDR8LcgpCS8ARZf2XJJ54HZ
IF4BM4G3SV03rfYzsE2qDmHX3kxAQnzslC1Ys+0c99OX1DLEntzqwzQt0QprwY3S
E+r3/ETAgc9G2ifeLSIZQijWQACqsQ8nVgikCLKhEgqj2wdSfSqzV6UsZLobaFWv
iRG7WKxLDIDPX6EPR85ZTiR8Qccn6qDIkrfXc6Wlbm2Ihy5nHOia8i79dbjRmXE6
AZhSQYCYGrJ20y5zFNV9hj7VF+kh95SOz9IIAjxVYX07H3AmsJEKQVKA6YtgfQMM
fO+Oq5dndDW8yfHxqtU5FF4mGnH69ghBgLinziKpOaAV25axW8Bz8/0HzwJjbwoT
Llw9opzwgAt3piBDYsZjz2WM6l4BVuUJQD1XhX6CfbEHVyAXj+iIzhqH9ogJxGt5
iH+RKr7tlFH/KjhmB8kKpNvF8Ko2LvxLE/YBSc5gENNK+XJ1m114cTpghZHC8ttl
/JQYjY65q7afQJSv3uxXxmXHylO0y0LYv0Gp6wUu3cwesKkUABQnEF6rm/bUSnDs
oVNwxqeKuOHziVaHqQZbnZCMkYRqvwmnZ6X3kLrl6SNJ4gunA1YbKCMqs1MUF1or
JQNahC7eyU1ksN63Lqbf5QUgFOROhv45yDvfsyGNV6lkvUt3hDdfc0S7mGUOtHS0
x7VIJmqS9e7rAQr1lvXv9DNfywhrJX0yhdKxssY5DMNPkQg7Jsx2Dc83g2/vjiYv
D9gj6bBsMNgNxIKrwfO4SlcoMKF45K8eMrWRN7Rbn5N1H6Xl3l23HDqB24oAgdGf
ss3gdTyBXXk0HWv0FVh4VvT43hVKHisYbcfXyG9F+mCF6dlQ9V3E/SoyVEaVPYIS
j92NQGPGQdSkCEU4L94Lz3pL6sz3pA2/SkX5Hues3cOGPBlFoeO3QfEYvVSUd1ad
kiM+jOBqnM56UYzmrU8k9jPqtyDQL8GqBG1fNXQbyFnzp44aa+/aAri8d3FJj57d
EZ5AN0Ax7ZoL+gBxZznoqEhg+49iJB/38/9oGmpKDUWCfgaEYw29nRRM0REWRTKX
kgGWjBNdIWlw7x5WFuZ2fGRN4Mbozz/1fIt4Euro/XQm/hALqHFJljut6eDZkk8N
3yhl8yVYYF7FHCBOEOkgsTckQG86vbKUc4m0Y4CRNUng9vNH+UqM3NdxiejSnmen
AUDeyouvO0gpPBataE+8EaZNwE3CJhafzjUNuJCfxH+T9QTMadLprfXmh19TWsl/
60C7fs2Tj20/v1NASMh/k+rtqwRyW2Buu+vSegwsNW1CASIVPIj8fsfjewXIhXO6
KVytqyNsHHwPnayCe0AOt9V3Lw92NEZsQ7sMzps6WgtxBeH2Y1yiSI0DO8Tk860N
bBBll+LYSC+Pp/0yjp/5MUkD2uAhqylLZOKrcg1LHnW79Oe9LHztS1BsW7mMg7o/
qTYQBBivgWhm+AfpAlxml3agQo/UhSd5sU+S+kflFsYQn5HJbpgVv5hkwKpuBhor
+ImuTedLjYWPmw4sYouIPHqJGLBLlJO1LDZoRGzxBom01Ek2a232LXueOEIN0TJe
ERNaQIFnVpwt2/f83UjAoT3CL2T/L8iE+shB67gj9Udwtkgx+OHEtRlPM95yFRQI
KXT6e3MSVWipxz53JcwW7+zIEjPJjfWPWQ2DLiWG6PUYlonaf9jn96p4w/moUoFE
chRhLRpXPGfCxEp8hiuSpQTmUpW1IrHXcJurgEdTiZR2Uhg5hJVRvxj3jSThzBVC
xn3R9Rd9vcJko+D5X6DTRCxdey62D8ilW45Lexu3AK6NIUr6r3F+gC5um5ydElia
FzEQMt8aV+DO/6VIs8SFtBHX1fHOjRbkEPMNJ4KAh6+a035w7T+cg6WRHtAoD5YQ
Oe4LWZirsK7BJxyNuniHF4OACfhj+xUE9+QodRKvYhGssJRBQpLza45kGIcWtXvU
oL1w75KikUGhBO42GxavvyCBEu4W4X858OvK48/YpPw02bIEjBLU/VxzxCXlqVtw
uizR2SZ91YzEU6IRswmly2rP5wghCPwv2kipmVL9THoLZgA4p/W2JuYu0P0a3e9/
h0DwFlofP3GmPDIZhdyxF4qB2PCIkbOS8nIb2XRAoVqFOg4TW7t1VLXJscUlH3xO
CJrWnqV37A5g68A6f/HpIlxCKcDPnmCidU082M9xhMHx4ua/zbFtYx0CmVBewvKB
+3E82pKLrC8MZiOsAjJXLIpHxn+pbDxYCYxI2zZIqRr5JifENiiKyV+rKiVvpKXY
1PhBzwp86zIedZqgSpT244PkVuwszL9cpXOaiPEWbFwXl8s7XVSUtYDM/kV+GDs/
jzqmOhN9oSnz0SFUrKfCPioLUu55oas9phu5Uuv8ifm2NemisrnutJaaz0u/TTsK
GAz2JX44Hf+kLBxpXCz8O7dJI9jHMeE1LA+kQDEstX8z3h0k0GVngcD0lUvRCpUV
luh+PyYb7TCmaAf7yRWqqmsDnBtWHGMBqzVsPTZprH41Hj/hPDnUj9eqOGKpyJ6S
CjCCzLfcK+QfwhOFPgZWk1AxNPna5XUjziGfRQ05jJI5v01F2umtjqafLqfxMFdn
AEe+iBiIyjw5F2gM+APJ2qFkB5Chca9Tev1namRvPgcjztOHvtJNiXI9rdZnijKF
6NeDjuiwWaIUQrQfjiGNsi3zO9y3ulOq2f1AHcdR0nzIOLejXRgIXA5DJTQ4a7T8
Uneh0LO6stkmZJ+9jsq1bWF5YZDhsuF9BHcCVyvv7cC+GOz74oFIa5ek5ooswuTB
cxAT2yCA7HOFqq55X5xCyrOhT/KiiSZdTu7yMkjGsAsf21sR508Fi8yBqPtxCsNs
Fl2EgP+AYk8+kh/NluHiu84ca8C9kw2osGKixmyWk+BNfduCfEOx4khB833L032S
opngmL0UwUQ5txiEjwvU/qujZ1zY2O8T83zxjhYTddyFomX7wlxb4bH5R1u7frSA
HpZGxbGdyTi00q1IMDiASe2Dl/+nPTRASgR7u0ItOXnKacki24z83ErRRMavGhCd
PJFcTqNTVs+lGP4aEVcJ7mqETeLydOLPpgJx1QZz28RxEYu+6agJuzWLtOAO+vbZ
XUyXKZuoNIIB49of5aiBKO9CkbE868k1Fq3QUDf2/HTo+ElBFLAJHVZTVejwhGTI
0unxyCKAhoZL8MncEO5zJ241Uzktv2YdQ9yMkULNPQ7Tacg2Xi7izHt7QD6e7uMq
mqSCpDAtj2icyxkb58+W2pX96Vk9EJiB6XhPCrJagag6mpAl9PYGdCgLJyx7L9k1
NiJ95aNi5B8fOkYsmUAWu6di1Ys6+Wb1N/ORNsU7SFYTT4zmqnoQ/WzUMXJm8cuc
1aw3rOXU0m2f5A0Soa3n/8NiDtneV66qksovzn9yAJOfneYszGFFZw8hudE8N7Ge
Paa4ruY4DqoeuU3c2PNI4b6OAbB55dKk2xiyZxD0KIUM7nDqR5fQ/1KT1Jy7TY8S
iaV9Qh61fKWcERprSFDsPal5DIhQiifQpVAjXnrW8R1CwsJJw/qsA5W+f2FHZpNm
vqKOArE5XIx5Zd3AXtdV7ggOmVCdpsR4ZxkLnyatLoZEaFXFQeMRKA+n/wYMjshg
Fjds4fdmPrX2lJX3ruZ20k+XUF5gRth9wmGFcpIZGrMpQnzwrvevgfuE++FZ9G5q
g1AVsMUYGPCBRejUZFZPaNv3M2EkSTFbQcC9R80AxeXF7NGtvW8I8EZcB1vPBVy9
Ts1grP9liBvmnn9BdoIVW+O9VEfNjnjVaH4ZzBiNVLi+YK4qAqS1nSU81a7lkCpK
5IQq2U8wyFTqb1fT/ukwi4wYaHnsh/ll5VJLJg3suBKodbMXSR3v16cmO8aQyMIf
Z1k9V80QwIjTb03h7svgn6Ybc+vXvqoep4FBdQyz12Q9Ul5zLXBmKHoiTN6HNuar
YGMy0PQwIRl4qfzWHOXEKaXwlyY5wN8SlcIFY9eDerFTxggymeoASbMCZr+0d58X
FcZwMd37PsZzeoeGt4dmjeOF5hruEz9rrOwSbyVJqBEnGlPGzFaO7ylKZ58vyH1l
cvUodrPePWAzP6615r4/qw4aXuIog7NLXY8mD8aGJg0HOxIViTsHkO2j0xqIwvv+
CsOIZ9J0b99oeayxhdN+fywhINZpZchwjOUWteu7Kwxfgm6JZfZW6PkjrfjRnjzm
honWBx61N6S0Eeeoup91aPg5JapWuicNoxmJ/Lr88Qqn5Suf2NhQiujCUh9x3LEg
je8bW1qA3lWCOTQBrCZ9+DkxWOA+Ov7uyInCx2YT8OIzW/pZXhLM9eG6GzoGbSIt
8JUikBcPWTxdJbgyfCsVxH0C+WT3r3HxdzfjPn1xHIuPVVhtKzzRRF2Cx0YPMZ3Z
imeggmp48VQIHZNxlKZL2wfO7VaFnPJ01h92I05B9thR4e3KlV5xcE/+Jyd4elsH
4GczfY3os4xXGA5q0SI95EemSgQVHrE7j42cZrc7O2N6mETQxFGJuHQB2yNHk1J0
fJFafz5Muz1NT/jDlEZSkzO+m+X1mtUJHA4g0fsUgqfZCCwR+3VSjtOmP7lDvTpE
fvtaucmUKwGbVDneQ5Ig0g3YCBblKQqfVB4yJ4kf4yRTicfK5bz1/EZC/YSS7P9B
SwNDXUEJ4p7ZpjyCQndBUaAUpR1rNVMBDZScCmboQFSO96/j6dABcVcdmeONAtcW
O71P69wahkwqW8H77518c7vkQsaBFbKwOcApKNmmcU+QoP33R8PZDZi6JqcV/heS
wlU3l9sKsU3uh8lVz+ZsuoM3wXG+cOGlKVdekDTRmrrF7UciudAZ3R3HTCC+ijXH
bHgtt9ilSMRI9MJflPhDMfm7xToAvHKk5biShGCJtVnubN2369kA6oLIvteSdMkH
t5AIZMtZuTJpwxxpOy8CWsKxOBqMdeqDyCZXVkYlJDJQjehM/3O7ZydW/6f5Clji
ywQ0cp5qzuKKxvuRTboMRhh5ZFuvJKH+5cyuAYkqjW7MUg5A1IaydIfTjXATVlbg
Z0Hb/+U5NGQcHG6gGJGEYSVRaAGjtGPNy5uXzrxNJDvEfy+CJIwySTplMEaEWv6G
x1xKDCXNLM1gRwr8FIGFt0A/44KgTkZ5PDJGyL7a1hXoGieaXyGZULsccEP791vU
xuo3RZQ4ijnKwVqxap207X9jpqYTsHtcXxhKZZLGURFb+ovCGZIU6C0rKrfqNbj1
8OIIIHm4nhM3qFIjYkGoywQEwFiL2YEUGJGP9ZP9btu32rtD1/FOMnNiEOdiwtxh
defu9xZdDhkdrQkOGt3z5UuWwFxyzKRTO54oEbhZXahL7xN2g3CdRPnpujpkgpjo
TfcFZdV++13rfnQ/+fCBi+jvViPANqq1g0Hqs2xaKBObEYOuvZqSHoxOQgoAuRUm
sT5tMPy5ETFLC7ce8F9xRkvImrUGq0xDAIJphUyHz0n4P7pHV3/u79UQP2Yaqvp3
bVqHvpa0+yB3hBAfqsshC+D5H407kXoEOv9CnfsCKTO+jZLXPD/KG0B6UO4I2Upx
ycALWm4pqX2F17l8FMQV9XC8Joh5sxQBweWyvjaWxSEEWRuzqbpe1Vc8TjM8B1C7
KJs7+EA9S0Uxv23eFiKGbA03KhlQZnZCcdHQYdoAjTdFgmz61+j7pIj1ug1eIApd
RY4c9DNtg1HIWtrRvhXBLNw1UAZX6LA/P+b30cPBgXceePK8tO+GGGcfMOFbK8FA
/IPktruE3iOkJ7Xtamxpxzq6yJMPYyEgOhEria+sRb2e6wLAhLnzPvkluoDd7goQ
0HROTagvtI3kna6BRycgBOW72Axmit8rMWIOfSv683DXWC4m5Z04A/p0jOQzm+zL
Q3SDYmd3fDYhz7pDkzJj8Dj2MzWzTj6oYFnpbqD8DBGhoyPs02sxRlXcvmp+n2gs
2CndrmltWGqwfRKnydQ1MufpkiS/05c9GB6K5TMNz89O1nWvDi6NH9FMcSCew8cq
Qo9XgZAkS7Vh1DYKfTQYVGammzHNrtzk7faqqkKup7a8PGtq/nR3Y/nVQurgVqmz
f9cNgxiXva2resIwgZTRj8FoJMrlbMD3FIdvqUTGClSs+fJrGQ3narWnCK46yEjd
KKCNbI4e9/xCfGt60A40WTUuuhsbfeoHwa2evsg8ljTCQYVdiJBvvxTaQMIvlPhZ
+h1q7+5dFR1pTwo0E7rvUZU8F1Yc4mEK6kOCCLGCZNcgt7EHMLdO70MYENz4oiGQ
VS9jSww/joPHZLFtTEHh3wcX9eWg/upoS6GHEBG0yML6n17QQUY2oh0TK1HHWF9r
/lUCR+US+7g5duNabSdJJHTShf9xJ9s+qop/ly50N6ftSE58YMwFqG6Ax+grmDFy
qKPk4xRAVguUHg4MN8YWXS9X2LJ26ZOL89fPDvBAf2n+LHhoiKAQYdTgksVrEgxe
md2DGH6ze2wkPIVLvcOYmqkKUE8Ap4hPJH8v4Cff1HhYyLuyx8b+fW94ceUDZ9Aa
T1IU0H7Bw3oawm+TAJfeJ+/yRSim+FKwC3idRX7yrbC0rC8apBLjebE682QW8Lqi
lOm4enLLNeTacpNdwAd2TW1vaZ7Bzoy6JcH2a45CNsXUL2yDux74G1F0IXSbKJG0
mChS4SvyfjAU4J9kPJEc7PDHT/yad/BhOQhN8qlCqDWaqYuFhO7dtYfJnPOFgW8+
vZamKEsJE6cUZVjB8BmykkKMy3/vmLvyrD7dYNu3nn7gbtu3GpdhtnO/cDiCwKIX
QrFOssSpYWI86Ko8x43F/4UCmslZ0X+0psjWY/db2TR9zset3FzODZQyQ8BS7ko4
lckDOFK9pOCt6m1yls+ILaqzlOiBr7sF2ocXhRDNTm1dn7t3afmoo1LivhkM0zk8
j4/meAab4rI6P2S0KJLR0OdDCNuCSM8mgB1IHb+sENplO/G0tqCGd+o+8gfYgkTT
3m249Hebx+57e/6qM+XXM2TgZzvPXi/vqz5XV2lA3MqTRaT05479HMRYqr4g4UAb
82DW1m5FnsLRAjKeEO6ZR+rPxZN0PGFyOzIVXbq9o9EvHBxxn3bc97vCJecV0gM/
yxei3vll1yTuTgcdak1NPqkaCyXO0DkHd0BCtE1M3vINjGmo2Zt9CTWXpVYudsU3
Yfw5y9z02LLzE6KkN6qd33HlX2h2tpg0p3YfpKogGnzYXE15YKZ03QyjHh4fUEIh
OtrdxQuQZ0gGy+cm2WcdcFuHXDVLEKfI9cNcNQwp3L8JVQYi8EEBdz97d5WgOFsZ
fHqASRUCkd4aUYdS55nvealkgErW+p/rGni3pxEcmDC/AbIC/3RAe8dlGLVU0scv
a76++strZIkgwtW8Y76BysdjVT1pflQKKoTQNmBssNOmqlR0NUiFuhQsK0IrElct
mpgPqUP0V7sUfdCJM1XOHQHOsIoXZDY2Jp8MaeMaLOXMsNh6vZ9zWBu3MYBD+Q4C
ogyKwqMG8q1nlWpGmyMJ8k4vIeHiuKFFz/eEFsfDNNsP7ds460CkTI7gD5QKT4+j
fjRGOQBjjukeeANHSmNkNAaN8T66Uu0VhstHq+/c7dQhZozENrNuEBcceg82gyF2
wL2hJsd9+lHAnDNHrtd2JGVsIXSE5fxb3lNqn/egeSZcweDr8Ov0Vn8CAyydErEW
bKm78k0teoSB93zK+fO8WAx8/T5arKXRqJzz7ThEB2gKhf+yYKR/BvW1j1ZOrTfS
7JfS1/9R5nbiZK5aDLSNGK7iugQowBAD+CVQqnlvHSVOX00AXFLQ4f6pKaohbWJ1
x2fOFlPuEhGjbvxA6vX1VPAi7iimSd5CcG65PxUr7Wi+UpcKuhqSdUcth5Wwcilb
vGBNLk/E8tL73WB2wdcFxIs95Se/lheo3JF0vdN8kHET7u9vdTvKzfHF2WgGpx3i
jCob1q8LmUgVRhQX851ysRgLDIWa8AumEfkM8AFk6opYuaXVlk6bKGwq968QKklO
WgxtOwImGgbp1azJt35UOS1rYFjVw+Ao+blpwOwZIBdbgca++TIumq/n98gg+26o
IvjFmKWHGXQN+97Ofyr2nt8JuBatvFAIzxWJ7LYxOoQh1qzlsveieTlpG71shp7W
rohM18Us2fB5qxrOxmoSLaLnpgyuBDKSC+rdjs+qDFK+VcLjTjCVQNX9Zvf0YOI6
jpXR0Y9M0b+znozof+40UtsULkhYflv1l89pitgEfeghfIPPdwgFv6VWvY/WkaQS
xK5E+kciglt9MqkI9SzTkzYh0nASUxARGpwvLVSIp82kRQXaVq57ElNlSdmeNIbT
sMg0uYJwGP4Atp0K1hRVNbwp+fsYrx4VhEbC396GLtK264057j1BscFc9sX8twmk
UPjULmQ61ShvxplvX6exdqNfNhCUp0GF8b+ZVZ71J1BmYTRTGFm3y1wA0OpfHlQ7
fXqpxoqVRpcmD27bNFQnK5FTHoMyn35gOc4exXePfR7cR/WtZ9+11Ce15ymWMCBx
h14WrfS8pxsg8Rfr2sNLD79uiODUbnCMqUuPRrMbxLvnq1Buwq9dLen8ToSOI6o8
QWpLv1jL8RaN0QmNutcmpgunfBgqT0eRJnFhj75Ct6fZ9jd/3POq+BEwicUfrbhP
2RxABtx58zXr/uL4USV8QAfgIjK11mzxZo3d26s6RJVbXmvnpKwNYnp/N4/bxoPM
iJ3Uo1Ek+l639Mj4Yurhm0XmavIYOMEaXJ2gSF+AgCNKhAJXOC1C76E22ivCLVcE
ng1FatZTxD5OyXgqBrWvtOjT8ChpysF+xizp3Px7xmLqRVY7YrgGm8huy/j1/+te
QXsgjtNeWSaFDkZ1uRdbFUIen+wvOPMTt4BiYbbfTy5kTBS+yHJNeqyduuGwwTm2
kdK0qLCyFXvaAKV3PTZCdGP2C/Tv2EOh1giplD9QKxfILkUdaMsdsyIR5LgLwdYJ
NKCNARKCo1PdolAFrEdQppsbuJEgiXcBJpjec8iIUjskEEavm+4WVGIMkSgUePSp
l+BrH3TFiOImM9XwUE1QJoka0Fciak2lujdvQsVBYjTer9uGW7RuNOZdzF5XL9wj
9ExVVwieABlIsyYUfPflL0vHDcUcpsCJ3QfiWZYu0JFhUPvgQA4+Sq4PqXFcEXrV
oBkxFo7ydFttyxYNUgpOkd1PSsBV6rNFmHJIy+I7nX73cYkWZnRbUEGh5tNRCzK3
a285MJW4/Vod6HeLuMI1kT3GMcnLxgu/ga+dl8QdsgsBKkADnw0w9Oumfy+aUVtz
l7B7z4ms3hK0qECTIhu11Px9+++P26FBI3srp670xynNrCcT+zdiSM7q84P+u2PQ
lS5JNxC7ExAiU6Ythzs8VZYLdZrvVefxw0G3Z513QlSTnnU9MYQ+cgCzHivoa0VI
41UVF6feEm5EAPOAmWY7tHBg1sI9SH7FkI7YIT+ITncL/wOvnR+afLmonO3RnMzb
Pm1mvTlM+8c59P82JPuzfAY4LN2uGclXQLzW3baBc0nkP6B2f1hi8I/vpZC/UFSR
s6oeVC0+H6zkDD1MfWm1z9cTWj9rqKV0XiRZVzqka63pZi21Z7ZR3OwuslKdCZbN
tG8hpnHzvP3vRk3pbpkmJNIxF8S50S8NyQ40fQPB/9tDWSpxkDgWgEOqTWSijt1P
rqaSjWJgZQLI3EnfsJGKmlL0UiJ9TsT7mnKSyPwieWP5fs9JEj/KlI0XD4b+NVCb
VGtOoTNfc0dus7mhaNZteDaOEnysBv6XFT0buf555t7ArIS2NJPSMRSPhp5V3ZoE
O/Ae5SLMTMkFyoJIaEpHPta1tGuDkT3c40fbfCbNgoC162oA6TW91LDCdNJOK+9D
a+l5eJzSDMbgNANQU4HbNPw987VQZSm9XbRwlYUmccGvy/RJKjCjBIyFCK7+Aj5p
yxj6qF7+++jiswLFo7OLjsiUTccs0OfEyx87gEz/849vc50NXHfMuvj2ZSq+6Lhj
1cyNg5oldv6U94Qtoi1Q9c+esEh2JvZq00XKRyP++pp/YmiJMEzzku8F7O0us6kl
/X7c7dsucFC0bRliexrd9YQzQFqOl6vXScDo+yy58Xo/y5xipxCkzIBe70r9uLCz
g4rq2lFTSawwyKdMz9skMszV5ImUdwiA+AIryKGsNw2vR0Zx6Yax++pgpXSGAL2U
uoC+emIrPuUIV8Z9dAcIqv5hRefwVIdIAqdzehMOiKInYL5fWndifyvCiilYg/4O
KKpVjPxo2ajD684pGhlOGQIismVDBmiIcNONNQqX8bldCRl9iKW8DRF69o/dwhOB
1TZiu9vARtn7F30GtWZnk0Zv7flltq1R8P4M+buvVEgci47tShbu8H1rW6+YtVVr
UkiumpUozNiDyL36j/Yty5+w4zG3ANjcRnMuBsNDC+TS8+8OQP8OdlmJxiPhzuTl
T2C6t2ywVMWPlFMn8yr4TKH5ZiCvZc7BXtxWOg8+xLxCEtqjVes+BB10zU81mvCP
bku+33B6KLjTWuWZNybhceY8dFj//4bjXF8Xu9KdsT2FKxHsf/folyh2syzDPLdf
7wW7v8cDABzSlmV21XIBGtlnaEQs5iZaEeInE+xIKqg1QQyNAiWWJAC08+mkjy8T
jgTbieayYHN33T/bzs+wH8+yZeAKqgzbWUZZuBOIW3wDYzGtgV/ZEFmg6quGBgaI
A44dbdAqQ8VAwgMTRjUuO0nRfnF/mBsdyVQT6gAzhp3RsK9qxHfVgsADo7PoQwVA
YmEgYuIZSUvi4fLi0jJhaYQfnX2WdmZV8Zm4JCHEcP5Z2r5THEZ4nBxvU6sBR815
WbTiBlgxNtynssidEJwqO1kyCKXUvP+YbcvUkt0nkTFpLKHdNb+1g9SQPP/s6sTx
faXQ0nSfLivNwy8lUwngZlQf+06Bq8trFObkIhC2GWQ5hRA7ZGsEkY3vTzGzCfPI
wVKXbbLBQkNylVvu3GX14NJr9HGOGxVTTer7j8iB0jF0gVV+NrJA6VWCOouylX1k
XnXQGfHkBSUDA3VrM7zLKR6s/f275D4p49OnrBkMzO5HOBQjvcNYW03oy/hXnA4X
IQVWwAo+b1KBCzgCCxHDRI09fijYPoOvnIRNFmGAFwe7MbzuersihBmLiabnGlwB
7I8V7j/BSnjBxlmpfTYu+1OQjAGjdWZYXDiBE034BmZ4yuVGFnH/PVZLhaLg5Lb7
ZNFf6isZNKxAw3BRf4mwoOk8FnmKn2w6NW4VSjBaTX5Pn2rOTtzVVSMMtN2MNmUr
csVPsal1yWDEEMkdKVW/Bx4Jwft9rPX1cCXnaPGGsOIQXh0655n6Ec1kJnkwNU5g
2zLiRJpTvJElUGr8uEmT2EBxXJLTYrV01ikuUjpR005dmYAxEBNxu9g1MWR5STjI
io9+SeMm9acHDf+SMMtoVYpONO/VCtU1Mt6KcPJlUzwFg7UXhH+a71VfNP8b3KlB
oD15X7Kb+Y4i8TtL+jxEJdpe0ToqQagIow4gpmci24TJBogQVihSXa8mXGUQDTWN
U4O+YVYV+02Gs96ypEd0sXOqKL0enIPpbAz7jVVYt2PEjHSnRU2y6ykxtF0QBIsh
q+5aDR9ZXpVQR5NHqUDQGp2oa3YsWWnE5OeA3GwYeaISgWg0ilQk6LK5iD0l64np
xosqlNIRxV26nLDxwmWprHn8q7SBUvKlV9dOxMfxzVUWxlxgC/Ni1iJXMA+5EOOu
55ZFJBd+suhFKxnN/i+lPufjAORDpAbALsUu5xDzineqvAnTQc+SoshDjcDbj7Nz
p5ggDwp93aprffSRrtfTd2u0OjKNB0K7vSiZAK7VWAA5rOBphck/pbe+Hc/KajyX
i4C/O08/pwb7xYDT+F1wBDMYj51esaI3dM43JFdkO+YLxPB9r46bW3qRcPM/EH5G
4oAyVPJk3tIojCEfVTlZFh/KhiNFIQCeHxpKxc4feugM4jZWct2p9lHuPHCHe/Ns
wez30f4nwhZ+Ney12twnTfvGG8BXT5y1zoKEa1ZP8j76MF7dZzlGC7oD44TfjOaj
8XeRpG7jKMAE36LHJRH9qhNUxCwcfvfXyQHCN78wvqBMl/KwxZl6v5Pw24VgopRL
AVYpp5id2/HJU9jKNTt8y/ee9kk23f34tSzTZD3H8iBowzm9LgHVnMxj0k1MdZbN
Nq6GkctbkVDlES8Q/+N3/WxdpY2NEVt0GYdjQ2ViHpSYDi1KHjrWtUpcAJUD6uh8
/I3KA8VGG6+j241Cn/p4r2+v5sVh6MpGOF72Pvgiw8t/PriTXEYP3GihWoaP+Y56
r/T4fs8EplCXl1Of60UtXK5s4eJJkr720D/BgBcG4BotW3zcNh3RylOQn6DbG3yD
S5Vr5isiOokP50PE4gYbX9EvS+KMVweHvrbDlPa2wzOMn6m354hfUnRXOii84Znw
3X3mnY7SiFiZMVueZNSwpRLyB+oUgkdl9Xe5WrKDetDU/RI0VZx94MK9iTYvZDQ7
AfjDU+lwBCIL2I3+vuveMPO07LeSo53LsYvE381BYGo6ZK8zOnTjhJP4nfgnDC4/
9OJC4zoO5rhTrig+990yQDHAgYT7z8pk6C2wlGi380c58AW5ilXetJJ4Y0S/bxAn
FdvQNQ20wnAApYnXgfTttITaCQtUC0vNBHAxDR7MjHjQjOk9KU+oCX1EGUKHepfc
5imtOn0U0n+kgNzOwxaOjCGvyP+Hz+BD2Ft0c4VvqQgiT3o9UCY3bNczKlC9b0+r
h2eoE/8e+nqcRfso900pTkdX5C31khHXJ/+Bd3sOkNcu4vKUZ2ZRLsqH5BUBnfkS
xdsqO1JA5kaL4+MkTzyqkQ4Ly62YD+a92OXE1qo38iaDR4UABrD3j5hAhgAfuD97
3xzMviKGKp3+d42SwkyNJs+A6xSf2uk8pfGX7ZchqsKJYt9W4Ezdo6XFPqS56ha4
ctmXdxZnBT8TtxuzeiJhuethwRpc8NZpKaAFWolqYPgh0m6uvD1XtefFbchnrKEj
W3vSloSADk3hE+sXzE2isIQ8ErbHXjD+i1cZV+e+5WZnl6XvRu491tnFV+mrfZW6
ET32ccAz7vnAWj0SdVLTuZuY1mPG2VNG9TZJHOM/dBmr2Bzu7wU5U5yDfvRyNhtA
Ba7pkb0RcwG7LqRouPfJmBJQjenkRfgUijP6nnHpxNQBeOdofcigneMJ0qmkJdob
gtC++ReCDB9ntYkXBe+Z+lwTURqOo6n4tFJMY8Fc5SmPcqGsb285nsUOPkh2LzJU
XxeRbZqpZ0FzzyCF8tLxkxl+jd0/HxBHczDH0BySzx1vGhE0nUgHTtU/aTzts7tC
azBUwmQ4iPf6haZ54HAzDDYjMWSpMpPmLmQxPU1mNSbdaVFlL1mZiiee9RqPPRDy
uvkztOTqecSFnkCv+BaM9pPQk9o4AredK/5NmWcweh7+kl6zTQn8vY/oCBUNrHxk
JTQ3nqW3cMmVTisSH3GISGqgW65p0t8hxLz5UagNr2ht7u7ZkOYpVjUvjPFZPu5Z
OsYen8Qdx+F8pZ2g8mVQLluQOBNo0EEh1eScvede+/Kr2BNnLvqBDdkK3FXOMyVH
sPMvd9/wHGF6+5+WRZ4nQ6W08dx2vn0CbUDgU1fjqZose9b0q9fhqSEWsZYF3U+R
MoFNithQNB5zHESZb4dqhev5s3bbcUqTTvVN0EcqiwPSnnBzisS+xYJ4as9JTd7j
euuKBUJeDLWDBeclKwboFqdPTbTmgevyM7d0f1BmjhWNRymDy+Dv9/M1JEvXC2Fc
/srUHPkDNQz1Bprw04Mr22z9pd6czhtj5ReVOaC/zCwX9kWPZeUaQ21dAijnU0vY
/wYAnRj709paai8vRJMoOtUEg+zhV24qzTGhDS1xBs+fHagzpU/UwPzPVlpDEIV/
GLFRBoeEy5s2t+33IrB290BY5EAx8vEKHF3zvzyB5qquHzmXdXqg0PyDfyOOTbiA
Temv8W7LyC0OmGPO3Y4pINl/s/LFTyrPWQDAk3a8n+pSdpa41eNqRiirpiQim7Sn
5SFpC87JtFAd2lT/KZyG0GoVtxB/NQ54z55quDbVsckrWTerzvpO1mZwWpO/uSDf
mcDhapXcRJVsHXAaVeEhEdq2Ecm0SQ8v8tq5BamLwwh9PP2H8m/v9tPZoDcx6kW/
4rOXrbBW16pn2RIdneQDFpN6mW4j2SGDKPgWpDdGxrfi/+BIyjgQMO06oLvbIVb8
iijJ19cXg7tgeN5QcNU2DG4wMt9JkDwTVbIAIVBkoO5/3ctB3fV4je/d054bsi83
XB0uoKRiHSETdajulefb0mdj8kGkgEoh6fDGy0iTN6+viLpjYiIvDGb9i+GViL5Z
JnGdc968XukJdyhaJmtmGypoQLAJkTgPiDPYk2uac7txbF4tOf2jV4fAejAzIN05
snlKmeNtQXCAAAyg9y3ZTis+0IdgD6feUtLGHklqJOW2/fYAutWnDBBfiyxsA2Yv
W3RB79Gf8sco7iXUHH8gw8oFSB1+dClY++Z4g2k6DP5PbaV4pVsgfxterohOlXNn
3edG/LnAGTThR36zEeN8mnxjOOFoz/+wW/GGdyWuRAFGugOxTmon9pCUInSiwi1q
4EaMJiDDUMKty+xrz74AzDQp6IvrhPl7CFBt4IhrKjpLcNIx2fUxlaxQ+JVF4kUz
iq5M2PMJcAXGpkGGD0d6Syz5V/Fhk43sZhVpp3pnrFPCl4wUs2dOsR28cn8MbjbX
RZYg5FCddL8IofjJVVidAuNz7J42f5JE51f3QQ7VoorwBPhyukMvdUKxaTrZlaet
7dAv/8w6Zvbl13VcoDwOvi/imYiPr9XaU62J9L+eyAazk3bkdO9hv2DiY4/Pln+z
XnIS4XfVrshIQI9do131QK5v0qBHTv59hk5hW3PHpHlWE+SSX7/4WfClXwBz6Y87
JvNB56cY6BY6wrYvKRjagDrxMXYbO5jLuQjuHSt4BvBHRt3vSRblCaVygY1iJGBG
RHbdWf+X5z4ygduBxfXhB4NfphrzdsdMPeFOXVop1FA3C5I00+pD5quVBR+oe4La
MfJfj+QnOpbpbhS8LGeJPFI/QZXx+ArlGtrAqfanqMde2SvuLdKCwnfkCOieGOii
4o+FeX/ci2xfPyXoW8ujHNjQaV+aA/IZ7Eil5GEuhuiUscAB9PQHDsEARmgegKOK
Ngi7htnHI6iB3MpTtXqwNmcCauUc1gqi1MnP1V5L7yELtYPTJd/npAvNAHWOnlXm
UGEpLHIg559ipzkkUWEvsTe8S+clpT9evR/OtjI4m9j08DGqWvPMMr5y1Erp0uoU
wcqE79Peim+fSLvYPocEQV0Kw8tkT91rhxfmZWPGhD1yR+3KoMffYuz/Thcd7cPD
x4mVNQYgSq3P8kkRdDKT1qlLK6GhLoCEcUuKRdm8DItZj2sxiavumJgY4GMjmteU
tmPvdKlAD/BDaCCWRT6M1h4RoKqAfdQsypUO5Sjv6JWKRVjvRLeGq6tk9nu797M4
x3giQW3b9mJNujnbvmD//6A72pMPvPGoj8oJutXgvq9K56RG/OnOKSOPDljtVgbB
yOtAD8GU3b1Gf13rMp5Zm0zv5P6VH6WPeB4frbKsp30wiuuJetHqpfL2+2Vfufum
VbKbuF9tp4EFKB+gMw+GnMEl0sM/QHd3t4XZtiyuJQCAjGvuS0zftwdqzWIQC2MH
YAV5wzweZOesWdyB2ZhUQ4Z5N7nnqOCMZanTX7cQVzKJuKXj6UZ2zj1U1lt7IPS/
lIT3V5wot6h/5MXXXhQo+4RWAlAVSM6PL3RKYaJbREW+EbjJu7/HM2tQRorrISTv
gPlRFBQuGnaFQGk2uVk2aPg8TSSKwfY8wQL1JjFX5U5SHaQkDACxl/8jTcHJDOQZ
O6EHzLb4R5fPo2q5vsn7FHz+/lQ6DLz5eOfXrM2H6fHo5MkJ5yRnGNA5pm84JHNY
cPY0AOYnMn1LTq7GpkzokyqHnD5waUhZWI+hDO1ZQkedYLaGnPOPW7dyh66cEaax
7Fmciqp84IV+0y5QYkYPSnbihKZ3Tn/ZdGRd8Km10S3jyglhz7cprOl53SP5lxH5
otpuqH63feyNL+lAEH81CyI1THdAg+VQye/Soc69S4ulYscxFi2mr9v/K79Jk+C2
LnzNiTu56NNHN8yXM791dUUZwITzHM2IlVKWoUIXUbfl3iD0EODR+Ik/ikb2oIe9
oF5QPqsNSW6d6higUqBjKtTrwTkKSEddiJ8BgCWLu6G0wxFqLCbP/3xk/ooxdFFq
mUf2kFEyOFCuSMD8BAhBLMyMn6d2rKL6Yq9cmL1M25/LMGMg4/wKqutLdKcn/UkZ
BIbps3602GnxRslMquA7k5wbUJiB34uINbQWm6ZqeFoD9GBrK9spxp90ysxZdOoQ
1oNGYZ5zJg9e9BWNIF3Io0xmq9Iuc+SVzlfulWvtCVjhxr+2VtzTAScTwPgOv3Y5
R+klcIyg8q2NjCzfuT4mvrJGd1GH9oTJyGq/8xWl3Y/eQD1TiQWmzpETt2Bi5Joo
ncH6XfWGk36RLp7fmVFTzZGAvDOueX/BxjtkXwpmJtTEoV466E4o7KaZCNp9fmw2
PZgDjuztE1Mdzn1eoaX2ZSHRKC0bdf1iVrgmtrMzyq3YsaKj7YTDzMamp3JtdX0T
7V+b36OISBxpXe9N4N0APx30d4SFP80fsHc0n/nepy30gqDhsQYNx6yhpj2pnD30
spdMM6Vgg44HW6H4qdO+R8jINfgqr39CQ21IMSdfZ88pz1F05FJ675n6gEhWaOJl
1RDt3rJrXbfDAPhpHMbF/6LmYlUVY5Joq6DYhz+QPTD+CdDv4CMDOJVgq75PCMzn
dX4vR9wBuzlGz3BWS0epmWr20r0Ts8y1m6d+JpHzdbInE5McAj4aZH1pbTTEz/h5
W8zk7cla4tsmxIT16VSCusdAzYMkwqDaJVn5tnzqTeiETFBj6sjW8fYvxlY2962S
3DEzbW8Ecj17iXoL6BtL8degDnYNx3D3Qt0rXHKhcv6ReuDpqHbiNz4U5/zaNqCA
+7YIH0cPN1NbG7CFwa+wHTtxQ0BoXkffwBc/cWu1t9F+uZQZZaRoUEonv+C+8bKB
nXAW244gJRG1glc1js8cn6eI5u0EKnwTdpkT2392FWo0Wx24Ge5o4SLEFVB4K1Lu
UW+FHTzaVsbYwWpO/qKwp2Ekyqny2nHTuLiirMK4dSAeG29BUp3BhnJlSBVadcOd
n84zZV8VDJvqWoYRia24dRNwZ5F4tKJNrXhnaRWDKjNXEzIk+SSfzvb8HqWAK2kz
ZXuJlA6kOw5S99ydxYDCs3NxahUwsr8zU1orjSvthoa8Hfs8GR2b3hOwHMlQLZSp
Wc/brHBcK/qWmWpXHU7NJ//Ps08SwviQFjAFKXuAZ9T6khNTM4rJ5GwQbNcyZfsM
mlVqQzfysfeAHzesIf1zgr7cSvMeQNQzeApFRkEfUdsJEpt79R6iYyDgSzU9ee2N
+yl1fCGlpMMVN3vt+jq3ActJd7SOvO/HY7lbxQoU+RB+u7oF+t7ilb7MfrjST8uY
FHM2ZeV3LwppKQOaatmQPd+T8uwxWp3ql3onVut0xHCOrf11whRwb0DGHkydFYmr
Cg+eGJ89TwXUmfp76zi9brTPgu15fUkIBrYfzac5WGoh1GfRDvG7WrbjBX8WA745
2BSCwUW5dnROHJ0BH4CTYJGdcEUoHD2k6xirdmBzY/G7vJ5fl2nBcPKHlp8tiYL3
u8EFIcr8G6pltcYwRKQKU+1ebll2UA9ZoeIQxmbC2nOo9b00SOTQDTsn47kxOlyn
Eud6BZLeIM9WuSqOayF/93umFivtH3cwkmvz8w/d8UmaIO+arEm0gL28lOcaFKag
1pIbeT8LZncCX9gQzbtUHKmHr7TUEr/UokLU6RbtQdBUXKbKq4ur69DU9Mb0BVbr
ZBVl7HMQcvANluQjh72H5sLn4P5kQWejhsywh/FcPUbD/R9FY9u4dzSiVZJ1mlme
FQqtC473PF0gY9QrOPzZH/gBlKO0CesKJZkwIHIUW2DybDVkwsjs4qegCN8t4A3K
j9551ng+ghg6E/a9koJNGZdz2pQ0BKzgekWsYfcDN9ioO83HDAeFq1VKDTSX0xls
ZEdEc2akcXh5fi7Ju+opXDgnw1/HFjCcZoShJgoYyAwmR1A0O5BfhUdv/5CXm88T
o3dPLFSQKWDoq0JNrCuSHI9dSgPjmoNOQIiRRhQkYhL1FuccovxDIiIUyyT8y0v8
1Vw8di308C5k2tBUnq3KhKfSKWYWFQurgObbdDCrPITxxKzddgS/G4yqqp74FFx9
kYlPAaHfAcm6iB8pqX9GJqkLHyH4f7Fa+pVk+9HLg8o+CDU2ZqY0e+wclB9K8KnD
sMVT6Cr8WR90CrPHQaGHnjtd4xgSP9UPd+jMXvt0GfZGRmapBKQ2Q7e576MhWw6E
8NtJmBquNCNFjBSiwBUhYCttLw6lGhasziEclcNS4DXJrKtXFi7ayLF0HzfB2WAa
H3G1pbUK9hGPznEj7Qcx81SR0LMdL2Ek50Nq3+zMriEpMPmcVMOQgVdDp4aCiSfj
PwptNumShE+66g+82rCRerFLBlYNIr63A5xOQmo4qaeEOmNuM4JSLQiUgH/0Cun8
RtgiIGDe6ix9DxSZpHdwXH80UOz3UDVqQPHMBpBryOv7CXCcpLG5ydVNnZg9PJHy
MFVxKx7I5m5/O9lA7lEkgDipXKsxNIGkqnmRnFOD0+A64xEXvzj0NNWXdWbsaFf1
g4knRpziFPfbrZjOThzTEExVKu5jLDZkjQjQZqIlSgc3ez1sHXi/08zCjJT1V+PC
rnT92yt42MZu/b0ER9gDVx1FH9+BtpO5fa66GRff04unqrnI6aAlIZpv65STHvVU
x/RECzaYIvE73/81U3fNi87i+syOYM+a8rGxfgEkXgSmgBi7l5KZumN1HgLZv+1N
NLKH/YT/w781lvBAWW9CakfT6imssJT6lKRqIL3mJGVE4jU+qlvfhs9iSucUtIiM
pVtUEyOTsn23EAXqfwHXbDC/GBkuj59Oan081wgoVmRtXe7VvCpPy7uZ2WIpRuzr
F92ocCyJesWo7B4e2aFCIgn1Knw+WR8MZjvKwVSg9mV3j3KmMBsBTeNB08vfOGNQ
WXSXtTXQbDFejfZtV05EAweh5vPcmveGAkYBWOB14fb7XXvnxlwT2QMJLAcC6yOi
dK7I4zQcgF7nLaBNWjujddSlqqQjjiQilViuGRwg4y+fETuwp+r6gXYHq49B+CsY
cM5M7tih+geosWCnhUZJumGmr4jfPB5hVd86HgYXfFdqcfIr9pgaPxFf3sFwZSQ2
tve/gH/UUfsz+MGw4yUScDRre/CS/C3ZvW0cvXZnBqVNpuCkmU44fFE2ClGUkfKr
/+k0CpztChsjx0iyzvGCzgv8XsO4opy9QIzSMuFWWRrtfCLMPavegkmWkJ23/viE
V8QAePIS9jDeooO/Ax3/+AgLeGJfqrlFdbsyJhl2cL81cGqyfpieztMIY32niOXV
TF2mZAElOy/k//JlDn6ZHRogq/zDFIhbnb+9wbDYLp0zznT9rnPZuIDAbOrO75Rp
UaJnlscu5RiAlbmbI9cL3BTUzDIN/yIXGYHKgTRHRZPg6m7GWe4m/O/qIQiqOPIw
nZSeGs0PjEfp7e78dSNHEAv5smYCaJ1eI9gbgWr0aoEdwiqc1Ib+x2Q+RLUreDfu
GbZa4n/OY+Kxe85i1NmxthsQIOLZHvx6lbQjZoiD8+o6Og2OCVMvp2teVck0rhB3
wg9/nFE/lHrthIVy/kw7q7JggggmH1Jf3hkhOHY6KU96llkiW6BKJS9SjPTi0Nbf
uzGmMIbjGR0h+3jJ90+roiZCWsjMb8y4vYLCZeCD4a6cB2pvkggPfcRXbKGoqG4/
tdjxZn7SC1SH2o+D29743K4QNSffSjEKh1OhCWePhdLQ+hR00u5KLYb9WFJ8kJI9
oMuqQ8GAgA4xCUwUCGqsGpjSBktFe483Mf99ybQLKHwyvTLyICiNT+TYAwcjxZ6t
qr37d35zZ+oJVt3m+BI5/JiVCOuzRK0DINrxpuviEAPDRhjpd5NRV3avm1b98GEw
nurtryavLH4dP9gMHDku1a63HwJ/hfwRgUpAKH7mwulmpMgloNKC0HWpXG9ndKqy
dOfoWKETZto/sEZ1vTsJxljo6Cokj2qDXcotlNtjat0+dIzJOegSy9Fx5Pm4IRjd
idYKq4LZ082Cd5400y6i9WXa0xrz1KQTwEWebg7n/mkCoUjsN1TuABQQc1cjT2hW
jZQ19ecbMVPn9/5YULw3JqMhgDF6HeOwXqSRxxelwJH7Ah1MPhqJ6a+fog9OJ53X
JkSnNMDfeVmLv0LpB6OKbM0eCibNBBrqs9aHG6e1hmLL6ASg0mIh8MGOG+C/nxPI
x85lRJo3NHPqFAY91hbZnrKy623H1/7Qg69biT3g/4qiKszGJaOZIo+zxy9cnDKY
37nL5R+BXjQ6iGynD9mIKYjvEw91t9apMFDQ2UD+osyGh9WwOgL94cwqgCXN3728
3shz8fUuwiiOWfHUZ5QkfQtrBIOg0PmQia/MlvGyfKy+x0hbN6Y6GDjSmAO79USx
qevysZEzSxNQGGTVnwykeqDH/duyXLLXDf9SVe50aWwoKE/WbWKQipWk7qZwfEKM
WoB7KDe1zgGP7ANAFubZD0sVMgcHb9JOBQh5f/fUJxCvFCXAcEdFE2GxUAECDEg7
uOqtLw/HWRGbhjwZ7Y+iUBP3e2qEwaU2Po0HV3DX2foDMXZV+BQ0Qs3XPScS3Fkd
bBi9XTufXhGitR/Bj5BNjW6K417eMduTWq+Ug7DiRRRDzTuLuU8IuOF+zaqC6QyM
QanOyhakS8Eo9RMitQF/IJVMZpwUiTJEG+ZcwJH6M5/xODSWJvzWA/elOpHUQPkg
oU1NAuZzZlJ5nUrpxmJh+0taRmWZmPgYbPJYnRzNTyizPc+8IW3I2s2lUrRbKGPN
mV07FpgYGFCsr3OAnEqr5uSBj+ETRXT8gqaJiecnwhTNpuWqnJc2UvE+hCBpuTUK
N8pO6umLuNHTDGKABsaBVgn/E/dR7EGuDQspsH/+MAskda6JJ+vYzszFUC+cKWEs
5HMsk3FkieRpReF0S9OqK5u24uoFjUriuB5IGJ9Pd1yvi5sm7yYD44i1SCkfYX+R
fofX/6QUW+E7Zvf8vYuHxVRy6MLKaoj0iyiZ+R0McSomLUMXViYD0lng51Kfqh7Q
6kZkVU5bADQN3gf/tG8YOyEYwS0IBSSffbmzj+UBgi1bX6yoUPhlHdfCozbzAvzg
wPU9mwFzDAgtdlAhljXxLS9eaCYpkxJtG5mbET6BqHot1AIsXN83rHHdUZJlYMd3
0/R8/ScwKHQMvvCn6jVtCP9wwUrBNCdApCYMpJQc19uK/C3ZnDHOvwe6xtdCB7/x
nRQFog4COxIZzVNUvWLriqVrXspQbcZByJ8xuseLIgXfevfKMFwc+fgorPE0rXEl
q7BA7GDT8MHMzc5V5miLrC/avUGqjACKc7VVHKl5CFf1eQqwC10tjGDhDzC/JXtR
Wn25Ng7fnj+bVhf+8/kjGmnFQUQyI3FEyoaoua8NTDu0drAZSPZ9rH5ELWezcYB5
FTwROUnX0i2BfhhWRZc0eXPwHbLqfV/X85C3tNOFb/Ys+lnLaRnAFLlJFUzJFSOU
R1NdOaiUDwlsh3LjD3TD63G2Br7ugWB3kyZfcpA61A52nK27TfZEZxcBflqsuUcf
iLaRi6AvbjmD3atBF4YFP+2R5IoeUkOtXzBMLvvHAn3qySpiIrAT2mvprAC+uanP
V+eBHCSCfaBlJOqDGxW5j5fzZxSXIVBIDgmZWYUoBHxOf3FENTngRudkzbvmzWlX
MogksmkCVBEvpU80vU6fNnmFWSmjcOUwCDXK97IGgv1nvpnq2PqxDCPCo9rw5ilq
JobaY9P/spwrWtbmzAlFYO5d1/ifkxelStSRu+XY4U1taviP0T/kBGikvANBWKfr
R72BMxtgj8Z6p6nOq/EuNSzug2eNRDCbtmHVtQ3ndMeRqZc9+PcTT+lErEdoZl0s
LsPLyvCLxvT+ibC712hNH66Can+fAucriAeLSUAy/NHdrk4Q3SQdonsMUICK9uot
XSwlWWE7fW+KFl5ba8+NIQthWJFwmTSRDHo91vXr5UGaZTuOnsJn5/8juaQ1u3ty
6qCdsYcIsiT1vvpun5vGNTnLfPOdGGT/ue5oaCGvGCfjzt02P6WY/4VoQk40pQ5j
alR5U8VRdQ6bfJUfGoZz5RowsvnJsS5awzgUCKydOvlYxtXzRk/05wOAQ7Qp2Iww
8mmcbq3Kjik/l2EwFLeE3ou0J+5ta9RgMvs5x19ibNhWj5nMBA+oDw3V6sLobch0
7g+p0CfDtlfMuuwC3vjN024Ar8H/GZghnIyPxpIjrnCF2mOvi5TZeLEAWYLGwTuQ
6UJ12p2W5uYv9i0fF8hDb1yLkGgZpO5iQUiZr+JhoJNZ/HL4bjgUYsU3qKYFqfYj
Q/NQLmh1KJw13mbidNxum4h1H3xg9WVuPciiPmJoJtwX/A8s3bLihJTMjibqVFI/
oTUkB1kkFWdH3BNidqYPiLCGeJUbtQBJlg+fROkDNQ0cNdD2mOoyE0ZDVCqJhJ+K
dT9H02fMtOIIVcUc26cPYRvOq5TiCAsQumkraMSm2Vcifdc17dQQeCwnfwKVYVM7
VsleCpA9gKq1NNscP+CpXA5AmFk8G+PGQ74cjc7m7b8hKCn9rPQC5FUtwz9j1Gpp
0INhoQ/swGp0707Kl8NrbK7zfFNlIo5fM1YDxJHyqfCLCd9Ftk9GU2zgBDEyDY4L
BWJ2TQbL+fB3Qq78+fzxQpflBr9fJ51czPexwun6gss1h/mE9ZxLFIAxpyGafAr2
WFVugoyS47QESD7UtfmEJIE9PzwpBXfJWrUJx4TBHaP1hMymuQKhCSvEtJAfKjPZ
32FvprDcXHqaMuBVi3YfTq3Gi1IgbR7YOZBZCF5ktDB91JW4YdQdPvgFfIvGRdiZ
t03mV3jVzg8AONp5ErOCaXwnzhLs8kWw4cw2kAG4MPKgQi7+q7sL6b9Lc8SlXqfA
SDb9LNpRqmoWyg8OwqJRGwbmEce6Nlbd6WaN/oNYegWCDe1aOM6JoNmEX3WuJrXL
7ein+hQZn+kN34vJl0pNHlal8bG4uYeVRcTFi6Z7JohJs2apaPK7vjvZymQavQUP
oF2cTXpkp4rsOFO6kJx86LSIL05VMH1W8AEagC0IyuWMTcD6PR8fAWDyjKceHFKf
Z3lSuLh1z2uWJ3NPrIgBNmw1bl6te0hfuZeqmy9FUPS/BEuqgjZfDMAcbM98yQht
uPVAhhKJhEAK59hcrdLHpTDy2qgzhKfTZ9jJa/wzUyU6DfL97DqjPabrjL91So6R
J9dtGsU+YQs+heTK/k4AaHWzeUEms4ksWTdPCteHF8yGo0JYS86Lr562YwkBz9mQ
SczoNeo2oQ6z33tybqzcmzXtvOkp1G7VnXfETfU8jF/JhBEBhMuJMggOanD+WBfk
A2T1ALwF1wCzFYE5F0WRzj8R+pECA5HEtHCOQ15VdFR3egkzHgwqt5nXlIAG6Qmh
VZ22QNhJXFYr2jSRV6on6kQcr74TIK6A9LM4l3xzk7WoQbxp9ullvTxU1qR7wL8k
APE4gwE+uQx4m0GDB62oGL/VJQI8e22uciqQUZgvoPB1MR2iVY7hsTOvmrQgxD7r
OWY/oBW+Hw131dCGegY/Ety80K8AkeTZKD/tS2yKiOnsthrros2IMHC8GeFosI5y
6qg8oBCQXswC7C7/awL/w7Lmz4IJa6B1vmN+xlDKNSGe8mduI51Fz7GTUuznttBg
uimgSXsb67b2s4oGgz5RahTjLnrCcPfci8DmFakvFS9c7jyE2Wtfn0UCMaOFwMnz
J0PJlffBZfmfCS5kM2RwWw9t7OZ6G149ZV/3J1UkHauIW5SOKwdWhXan5iFEncav
mL63NakXTu5Aoz+jzhCnha1AWjVJxZgEnhaedeIclkKJHlDc+cS+j2ri0PDB+A/y
rhuo7fzBQWUKpmH8gY2s978qdF50yjg/wOEm39DqbDknaXi14EV49IihzO4rgVxt
Gh88hzMRiLLyD5HQZ49yKUecJVvWgTXHerfbJz4wjpjVXvrUysMiCAqgaBKkidNL
cFh7YIxx4NFzsF2kWptHITIAetMsAXIbaaCLami7OditGK4LNFJPHJsr0rwnDWML
lLv0KyGlU8Jg/xT0hBB+h0+4E7Gl0byJhnk6olyNzkqKhP0avKHLe64spTlB5KuW
IbacI1HT9wTSGrI7vg1A4EZ9n6E5D6WaCcb+uc/9KGlVCB5JZX4LLfigG0XT2HJx
ruUJvQ/asCpWWuk2RsbMiYIk4OLnYVia6HMrzf7CNLLU1a8i2EsmodXthkyMNdsY
x6LPn6HWdsuzNcAH/YU2Ou97KKRdWh8putBaAGIvXO6VVU5J2g8uUcwrNW+SIEM4
duhU0HhBnt66tis0JJ5SHZ7Nf2y9CEDbVDEskaEu0As82m+yMioGLLQa/KnXU95b
95/Uc9BCirS6nGj83kQsJVRPIAqCifZq3PhS7Q6NNRWSdZapOMUgqXZvPF2sh8CQ
e3awX68Xnu2v6NvbvJ7mRMmvK+hd7Xwe8p752F+hepqVABbwD/R7bKauKFwzNiaG
sykk2VKBx8/3QKTs6tUKFYVZLUSaxqCNcn+KLwuT8l9EQkomsphmPDVOYyj1SO3E
DM0yr+RA6z5Ord7XCww3qMW/clNC+Z2NpmaW9C6BWH30U9z1jJypdVvoZyXTE4tm
xYGWfIuJlWOwSxhjsHVr+WoSSsU253iWOmrAZ2bfCmG/K/eroGGxw6dPY/1+VqDX
/8pbusmZEt+ODBHoalx2j4VuxNRHfut5lkkZc4yjx3kmvM4xk+t5V/Xld8iMQ/EV
vqfvofZ0uJPBkeoCv5Td7iOBivDCyH6dWe8Xwps3a9Lqqn9gTvYR7DgqrnF4/biJ
GM5Jrvx03rozTW9MP49G+cm5h5dwS+Hc784yji1pxiw98eCjhTqj4DxNYx21C93j
aZ34idDOss9WXD2QzXD3Q88+DTd2UKUiBxd6UnwKuZ2brw3Hcanz4JHCApbAAdig
WDuAuvmXQugl1WT+wSO6C90j1fpk4PlaT1hG+fSGzczQgu8TJN+s3JGznPU3FN0I
UNbnSgBlJyIj6drYrOsFjkteDGc3Zh8GX7+T87ycvcgsIYhrwHFaIzA9pg0MpXSG
2iDhu3PcE9Avi3Eubgf3eseK9vKCHlKHm2eroFW0HmItz7bVPmyEcmefL9tZM8cB
sqYTu1KbVHxyJdu5LCNaqBrfOcXzTaHUCJMsRrDOKMPo0ExwFte+aMjnSCytPQfQ
xhqPh6SSSg0DwkNODrKpn4zQDIV2BvJLnf2XYoy2di3D5oj274lRWJp9s+Gp/Yw0
jgl5NX0yFDmThvhGSMr3D39SVym9vLC7HpY1Q3bNmdi7sbCgH7ftKlC4Y6h6jbfL
1ktig/CdwDIOexX5BFwuh7PrI3G/Y4NZHBi5ySOVKy4SiMuXHPfDmqnea+Kp6PCf
gYAVw7dx4RJpWqZYuzymQcFOQlarR9PWxDqB+vgebFRYM8nHbgxHu6s8ZfiIi/RH
D0j6qxwHo4lx4IBcIt9G97TKqWdtZ3Qyk/oc1P2ChEaccBkqL0h24z+wt7787y0e
UNXxM9eHELwnSdvofxsYAJ5ZfVHRZmh1ztgeSdJvFN4K1vnHHEg7lSx+vQVU1W4m
dJAwC5xmM0cRUIcUuOjcgSeKj0a4azDFdA9Lgne2BQS89A/UMXBPjD8kAPoUEYOF
rMNkjr1J1mO439t9fMcOLDjemDqOaeaIUEq58757Ac39oLJe2kQa4V31FrAhdDwV
n1xteqtrAv8hQV3aXtwoEN5ZmAiV1XEdHFLlUh03iyLkuu4SDAo/lxvQGTp7KBRJ
7wVhg9jEvwxV6esz5Wgp+3oh2w/kayb4oat5sMQBd0YMMKw/gKiztTbFqz1v1HUh
oq/f408W7F50yToIt0Z69VZJARtH8f2I3xdIewooSwBH15q0KJmXRfAqu9N+0ZI7
+PCU9nU9m+JEyd+Iwtv6v8Hy3AVTXDeHvhLwcJ3cfdjPayPhPtn9wdJPmLGt40Pa
znOzUwBZnoI/JDcG3bIC0JC5Aixj/I/BlU+0jwSq7nXydvkh8Pko2hmaQqi84KeL
rKFIqDBee+Unb9vkSWRQ1Y4Po8qBMAEUsTMFJrPfgnRfJG8y4l7rF3+TDfFNwz4X
6Un10FvjaijcyAyCi2cg/JsWN3EmJdo2hpmUh3Qk0tqXjmwGvZ/7831wiBDMRUVG
FOty2IM05TE7b63axIdnUA4b3DZgfb8nSanl1Zf48CvY3MtNi72qztMjeQQR3zgp
rOL61uy76NDUows7ZUIbHzcqLjyBxPZ5d4/dD4OUEJFCLG/2r2MPzwX3BX7d51PK
alP5K4761dFk+Zm18d+EwIppdlHwqYrq3a9duyrU+mpppyPB5LCvl2m/N4liD0e/
b5DcVTh1wG5sRvo1JJc155JZSf6zFfz7fZGNQW/2WgzSODV1oJOMCCneE5UHB52x
cQRldz6DFmYICVz6rBeo2xElWdpsJnJgOJHnuDimmDVXLwCPfsnCzMHdMC0DJykK
cJj7/dTfMR6CHKovIjyaizZfc8OjzZMXoybjdN3c7mX1lj5LWIt91HiuJL4N4Ig9
6qTmT8zYA6VMscsacc3z3HAptzDKZ3T7lx64e4EI3I49qSR4PPI8gHVj16wx4mMN
WIovjHCJXLXozmF/fsJ+Z6p8+4iA6rsQJHwJErrb5+8Z0cfdEYdJtzK5h+YvHepi
n2T2kW9WXyPa6Uazc5hLjTcQn7Jznhb8Sq5KUkci5DCcdkHigzcorwM2caKFLMiE
9ywWqwsL78C2Ro3Fd7tmIoPQ041KLmcijeETwEfNleU7v8QAFsO+1OB/dV289V0L
NglbABib+NZ8uUD57cSAHWzyjiLn6737s3uAeklB8+E9OGm8tbZcehvZ++L3fqWd
/+QtzqDq4tT4kPnuYmLKmuJ/7OPNp6RNslUtqVMAabUfn5lW/rudwD2PETMnf9qu
eF7LxIZ2NN6JpqVSe1En+rKtz7+vGc6UuEywgNEakhvzDEdbUr3yt/dfmTi3j5PH
3NZzKSaPJencIh55oUwzYBv3sfY6I4Tjtl6N/JcntB/PgewZmRNPJxDQOo2c9T0l
pxdXXYP+FEPawE7f73Gmxt47ZZXpiQjskk2rmgUN01HILi4IIrqqnlxPZ/m1zHzR
iRZhnbQpzXEDTgsZiQ4xA1vDcFdBxlVjjXDirI08AYRq5winzO5/AaIiUD6Dqxpw
EC7FhZkmd37J2ZPdk/CJvPDvC+i2E6ouygRB3YyHIMQJyMx7dp4bqXdaxbVb+OqW
mAb5d3FPd5weQyjkAkH+8Y05uxQgdmsQskZrK4+AjtQpTyfeReloquMvdv2BkvNW
y88gLrefH1KCs9cm1WlmfVuLrgIXwqJ6Fg5jpPWTn6m1pSTHuidzBkbrAnbuB3PG
gDNHF307dulbJharyMDUGCwrF/aXcPUYELFA+KlbemZbpWVdRhgGIIyk/H/TXhYe
5E/upkOkDSDQp+RijCHsO3PRJ+232k04BuU0nzSA5wltPXByNE4C/GRoRJAK2NZe
XHJdh/Yr6CWXLqCFlee/KF4CGXS+AdiI8XYJA+jyembc3upxW/JFvldZ3rg3M+SS
ymHaBIlkzj5NooQEs9kI/iYtGQdpfXobTzCDSbvsB3yht9qxjWZ8NU3KTiktfq6n
3C1SknuoVMRj4BqiRCyNC9Cpuj6op6uV8k9M6pom78fMNFdCfdkfaCTJIDDqb7be
wXj5E9tbZLQW+yo/Z2uGHM1duHGq6PGCq9hBDPjsRQCJTGYLFvLB1IwkE/8dATuK
O9dNVoH0zZuPE00zfZpFHYenNJGLzwSxv1dK5M3uI8BGx938QHv6xR3rA6vhH2Dj
QMjIC2Mruof5097/p9Jpc861BzOwe1yZu47p4XFh8fzJr/h43YNg7NWJJEz5zeX+
xF9++2AWL5/aO+00U1JIlLep3yTWMit8Md5hMhzkvWt7e+LzvbSYxMRux9JgKhuP
TaI2scybiq4HtSqBGGs2pwCceCO3/HMQuXo44o9AyCIjCPR3Nu3FTQ+sXQLZC5lW
KD0wv/rlN73F73lo1c6F3ox/HKBcK9xOSp2EPC7mvEu4ALt3FLvGCwO13n7sQ4HN
Ezo6mHp66OGidaSgxv5h2ZcSv9JcsDN346Zt92eIO6ZvBsv5LYl2EjhxybqSkAjs
FrAjAMs1c2WHHgfMRFqQv7AtXnHTiQKvdOPp29tkNIDFxChlFkEH7iVZEhyi02Xy
OmQJUsMluGip0TDulq4G6sKRra/C5xpP4/s71jKuuXx2uh+jcJtOT9fg6CwPiO4B
JFFmPGc7eLz0irBvS1iNnUl4wGBl4rhIuQ/59Ku9vo25Sk2Osa2uEwbqe5q09QY1
7fWTyD6mDOpWim5XaPV7G+/4jBcVNsfHHiomSiS6oTg/NGXspLJ/Bd7EtyCEt4dk
MlzYtLnHZ/v88GNS6j67UAZjXV6UtFR7wjtKi0RGuCXGOcLyJGYd9qotMgZJubQZ
+44xvXhbRpUsQ/5WBlezNcHEk/UqwoUzC9yeBcKzZRot4WhTckzpsfhRQ2J16JfZ
yVyg+W0dQbTbwCJpsy0K0mrLcMFwLRzyalDM1eNhy3uxzVfnCha4o/i22dR/vjh9
suyHjkwE0bHqA8k8mK//9dJ/ThrMy1vN2V/9QHOfMNNHtTA+rsIG8osuXQzwYZ0t
QCGTOWquDG6tuJ8r0QbZjJoQiOilXPhWdqBY2dFWVmz2r3uJAWN4sBF/fC6xW0he
k0oukQUKkzYRotTyQHomCQ1yolIVm8wW/p0P6xCCsJMUGdbzaHK5sQo0LEA2nahV
lPR3LygzlcBAXYCwK4Nn/vtHML2tDoMkuNwJqS++3c8llbQ3jb6DH/zI4So5sVGQ
YbW3jMQNO85cvWvLCZcjnx+2GlU7GOFoehL3aILMVsOAdi14pkk1P4TUzNqkxmzw
b4EQEMz+858D//Zwr1J5ZgujHVT8k6P5ZpeniG+4PfOMu8N1c53oRNjCyHB7KxC2
bOGgav42c9rlMf+htF9P6PwC7gMHE7kMzAdbpfPBD7lwB7+qcawu5T0RNw9n31xK
xhXcIjq1qPmegIyEzo4vPUUV295OfVrrvNkYR4VX2UXU4hcSuoa3bIko0V1flHzG
L6VUl24oMn+El5fJv6JHUOofAvx1/w+Opbd9oVK+/wVHBrO/keM4kStdKhe32WRP
nwNcVHzhfJYDSz4F40D923jy2FrOpBHPGds6XGoeIDn2IvkR6d+VFqrEhTervY5r
Y2exBnYePFRIO2Ks5G+xkk4ePt1Ef4fMOUVS5Xs/RixObVYJHZ4S0RnkwLDxCY9y
ujddqcxoUHYzl6E5JluZ2L+2/eaRhC5E0QRZVm+vWPWEai5hIp50cO95YEtZ8DXG
mpUerqPIavrnOm7MHZxVPlCTNflsoiN1eYnGv2WnpfVBuf93slMlGOdgP7Fcg3gf
BDhcJOYUKXHQpIOS0S9JGZ35iTR0pTRrHku8qggjApwQkFq2m6yvzyE9P1nlyBF1
MgxGgj89s7T30orGmcTmPLxAUM8vCBRzvq1NbjRFqyIFUe4E107gGSdfTIMtvKYt
uImh+g8iC8PZAhRsopGPYhWpqTRrhPNWesHYoUEFUmebP+dfZW/CDV8Pdv09fwF8
HE3aodYWtDZWrVnqjKwGFcl0OqKyTddxDzUIXQAZbazZ1CG5eLcimrou+dQ+fN7R
YTmfOkezkJ1zUEV5hE0PxzpQF/lpjXvqezOmQSiJPozNOaG/uw1LHwe9zuHJT9Yu
5AlM2v04RZITGyg8RCP6wvMAdCNcwBzWnuDXhxc9Tzjgb3YpSVOCa/MfCY10OzCr
/JVp9EY5pwHmG3bhoiFeB2Kl8Qt+2EHTo85j4Pg2uzr/IdkFRF0typQt3ABWAI4I
EWjB8keVrEqXEstalV+O2pQYjXX6q5YLyNDzgGUWyp9031b3Q7blFnm46f8BS1at
HecP94J8pxGFRGZxzGwH6UXLRFyUAfBUNHC0WMtJvmWpzQuAYgE1uA1Lmt4meUcR
JmWdw6xgvKXYwgAhqsBESWSJlwVM5tJoBpCzUeDybiFUF8gutbSEKr6XJp3GfGHl
hrgoj5OLqOm6PW8f0GItvCV5EppJIsYUi1ohJ9Wlt00qfWWoSSqr7uVyX89WCMM6
5scTRha4esRA5HxLgJAP5KJXVQ1mEZjiBdqixUisNb+d/Y+kPYSZTCb67O1yCRZ2
96WOxDegks8r+1JcWXwAU3Ong8HcxBNORg8JjkK0/sdELbZAOZtvf5du/zgzH1dc
S7sGFrOhO8dW2a71iH/WMMU2PSBtRqjzZJENKA0pLP93tBOcWdM29KUjjR73f5xB
i6wSo3LAN4NK/qxjzZvM7kf2vOXg/IF2EzMqDRdH3GPW3RMZzZBWZMDdza6vPl5a
07Tz+z/+2L8kgjWoziPRuYMRp2cF48KjkY+8FUxocoZgWyNCDs9ZzBGOQupU19VR
6VOxSSPisJZamQB8PUg8fmJ1jNzmt6QpsesyzXS1LckDts34RYAnt53q+ZYKrEeU
2ldVSZZdcPy4yiC6T4K1/Ltd45HIfNblpCTL1c+fUPLCqv1zfrJo08/fpiJmdINg
ac0wj5HW0oaJxzDBNg21irGr1gi0AbGRGRHMkiCylsEIWMLTU0Mvp428tKRVtA6b
i2ltHcj2Rknd90ncXgfW3URPALze14i8NM79sEyFEEos+Q5sOkGanwxaPm7Nsrlx
REbbFcxXhRaSi7F7DcosLTOnzCt665fDyUBl34g3Jr9Fo1guGCVXW8KpUhJy2ibg
yUnTlvuKkL0J8p8msgc1SRAvJDgRbCjIDLrxQe3yH5Xu7uK2l2I/vmB21t3P9dOQ
6W9kn4Aw00wTduKa1xXI3DkoadtNa6fGcTD9PGTrxoyKuYaehhM0L0eaazRraQGG
6Bpue6k9/CVJRla/Sdb+cejeKJ340h1fqdi2bbCf0FbUiLQmWshvqIPGzI9WBmzZ
/OrCHwnRQv1QNp8w3a40MylGygfRwefbdKC/WlmPxkRczo6AynbU75jjOOZoXngX
3D9wCTOhUrmb4tFddi/us6y0zPxxto5ObS82H8uiW4haLWgaiK8VwqzTYefkl6zc
MY/N4wM6X0FJvLuaFDYtHXwe1YS80JuQrfi97QS6LycSGu7e7Ds4euQfvutD6mJi
SHj/Q74SiLC5a27dryzbUrWb7h+0V/2p6pB6rztd7BRquXKn0e7qlHoWw07SHTrL
qoxIYtM/Q346ZXrt1dFurnqPwbcB5T659T5X3xFptSXRBCyjpi+zpeQrA8kAq3GI
fbDEgiJjJh8h1lPdbuCFH4mUrbR0XWBkSihF7ZdULU0LjRG3JcBylW/h+Q70Di4A
OORg0ec7innTJLXDGPi9ip5F46uypngj7AzuE9YKs4qKxWnTngxizq/ZTNl6LIWI
bvzJ2yrzwYpsnGCTlFGBgNkThImMTtchbPYfS6ZcQiiLDEdDQYe9G8VrXSS1lFKb
pgAjyrcyzspsm3ncVS/rO50+mngbzRwz7jRQOg1V3iTnTidJmx21o6uG/PQCYjWt
5fLDLl7vvxf2H1f9/H6CRrlA+J9LgjFgASqfHYQvIqpXl5UPVtzqsY8tQC6+Lc7j
FDA6iSJ2ms5t8RGA0RfHC5i16owghBvt4u9CqImp5vpcbCPSTK7qp8eL03/+Dz6i
teOmjZV2E4llRNC8MLMkw3M6Iilnpj8wHq+wm9h5TFKJfwmKekjBQWG6rrbpusLK
Zzbz8dglGbXwhQei1dmzHh/VIhFUAexK4K0xKbFkWvL2r5LPNz1L/udJ7cZYWjxN
nfjweMMO3cxi+Hx3myhqjZtbkoRmo+ju2MAZ4yufc6+iAIOhNSpoNOExAgNc1rrx
8ewLz7fqJmCabVfkt0vL4/E5hAUN0NjT3m9kUC0+YibyhtB5+8vceSqKTeKQIoH3
VlVZgnBiUE/pVSLHOlr+R5lgOWjP0mvJr8BYyxXVDUO2LVnB1ewvU4gVhYFbHYIA
4M4SSRXCk5ef7hSksB3rekbGuu8GGya16fmDwtrEFE7YuwgsqifCkrv2Nz0prhC6
XE4n6SCFWcXmgYcuzPjVD/xRlwGjORYBUmCbq1iKaPAh8XgnVCPQZJR6igBN8v/b
LK/sX2kOQ8Fyy2L4IF7ccnO66YGtdyjWbUqDM4pwhVFMFi42X/i522i9CzoY4Cq6
dW/43ObiN9MgR2BpNTRaSA6C48aHSk1kMVlTUdpO153aDqSTFjWbss81EGqbSakV
RRfCYZ3T9jdEPqG5Oc7XC2lfKoQPWJUSrPRNNjY0BkhpcSvwwxYzFAA+kBVmHw3T
tzaT2xMTK6XNe0gNQ9RFUa/ty4QnyRrCFNyMaS9xS83GS0PRSTL5bxAkAsYDVPiM
ocZr3y9116Rvaqop4aeFuGxRvp8Byqcc48bGJRU4y0/th8ZMzth+aoAQY0qSC2K+
mDU7AFI1wXxXgY4PZEa1DwHOQOJfk/5K5BpjjPuj/PsJfZNnwji+chNxa4QtP6B4
wXxqbTBjqMfns0yinayjmArw6xjRHA+dRDzM3UVEC0j0rIvJvg5Ex80+H86SgL78
oKTxB1RbYgZ92yNjEdDIbytS6l7qZ/qd5NMTYLlKQD6HCFiguOHm50Y3xdWvVGgh
dwYi2I8OuZYEO8RVM9ad4AIBDaOEJhTaBrjB5oqYKSkLRsqxP7ZRMBdhek9Gr78b
LJlY2jNFqnVZlXbxBUzN/pFkSU/8bozRbqtnUYK1kX+L4e6fFi57jDS1LCZK2+c5
/GfX9vp3TANLPeqrKJA9gVqiG+EsuDnBQynkYx+Z7Mpu9uPMB3kdVK0byxhDeBM/
lAEomUs8i5Ym5lHdWHyOkmj4Xu5giw/ikV633alZK6D9xLcKptZROq+N1lD2ZZ4e
yLubw3du8TVa30j2zIAXnStP1y5qOxc+HeMd3A5Ls7kUkYaZEeDem4oYkjh9Q1UO
SMD8B9s6CG3R5IdLaAjfQQkxA9pBflmV419EhZvKdALl3TjtgI8kqz6TR8Zt8/0I
YmNPS0qmOYMQ+k3BgWq1Rlyz4OLsVycHgi+HAiTYs9HGl3q4/WjqEapUvUxELiAj
iNQDK+cw4mc17E5L2RBpDSahdiOnMeWnHA9MNvwToMXm+3DQudECMuwwkUPmWKOh
qV8dqYfwsNx+xdI8OzdlMJq5eir3pEVMWj1pleALmCq8/OQwD5VPw7RgyhpbyANI
ahimns5tdFCDc57FpyrOKM5egGco6HaljDwOPDNJKcLc7IYWn13MXty3lIuPyiL9
dRVpyV+RJFRQeegJBZv/VQ2O54MRsOPfp28g/F+kkKsKhLJWcOty0tAV2YscnE6J
tC2SVZXI3Cq6bpVBP2E/CeHtaESQz1wzwzp3JCnQppeajNtH+CXPe7Qq8OPLp+pN
vsLyY17m2Bsm4m0+HbJzFjT/xyhhzLhK1sNst6IVtWDwtMk3ZAF3VaRd9SoFNAjQ
J/71w5nx/6YNyATcdFlK5bJWjoZ8Sm2+v91c3q5URdxmYTl6aVZg0BLEBsj4n39y
1/1/AXH1UR93vFumAv6capmDKN/yHgJaDBWlm+YnGoctKh5qdFOjA8HdP9PfHpB3
Ie3VGwItaueEZwav7D5ejkRBSw+F+ki83dtA6jZZpv9/D61eciHSPA38i7UwEomu
mKiR/doTY9j7KduwUJcGL28CPoK+RzTR+nbsi4rMlJncyJU2vt98OGqV2vs9YHfg
ora1S2kgO5h/UnV92rEvxl59OOKWwrnH4qGtOpU837SevUfCQJgWbLtYKoO3PX4M
aYNFgwaYtY79oMzPhxtu0yOd6eLAKBpQPYwaVC4s6ukCvzO6db9xFn+PwI3bx+fA
ojIP62cqMVzerZkAzeXo6cMvTSfqOusxYrM3MA0SXSrf1Ixeh+ZovpEjHo9k4AYj
CHhV5pDO93vRalSJofafoBHjXFJHInu5HIUmSHvBLRvW6SNlCOPHXe8Y0FDTg8n2
phHVAkOJQQehRttlodNMYdEDxYxcnifAFzmVd2OXaoLEMiwP2D6vMq2CEMsxn1Pm
zpsJ45eV6O6DeZvt8155bMPvPEk6HhQMGM9vzhlT+80/3Kc/0a0QB1dfnqV6UHx5
mUJY4z3IszXT3j61Qkru9XtJtcDfARe86kzaHbdi52hq60HxWkat/5EWv4KEl/u2
xiOOXuHlLMEm6fgOJRj6R+VoonKaqax1850AdUalNBEKHUo1ytXzQTGLQcKevQLZ
KT/WkftXnLIPKayQtsW/n8gAEfk/xkpmyYjBYFJSDq8ovO+xNJBiXdm80LPh+zGs
15I+AJuWj8KCkwqFiA6lCz9wzLvQTzDV5MdIwXaH68XxzCcGPYgdo2QcC0xKvL7R
ICKE7U5U1HvDQ1xn9KwkJHBS85c9KR1HWxn8NQ4EzwbmndQibXIYfUG5bun8HVcx
ORdD8LPToDWZB1Fi1bBIwpPe2iLC3uA57cFV+PY/jJlRBLN704DAaNypDDeVoWw1
JdvsMxhsYadmTxrgdPKgd2LVW5ID6KHkQAypAe0Fa7Hpmvo0SMS7jyrUpZ2KhQzx
JJ59+ncm83wrqduBYbEpk889vZmDrMpl29U2mbIl6aeFdXe/zvqgHmA3zkiQf8o+
KVczfPlwfrAuF8n8Y7AGHuaEkPVkHxsxNJk1OeVVQBhxR97CeukWuEfbO3rwMqJo
x69xhgyXpQnwLWrIME8NKjHrtqJwP1js2GwhRda0W3XmnQRnyx1e5VMegIlo9SmQ
80TusddmWkXw6hU2PN3wdfEVE8gg65wguQp7a10VuZE8Asc+Mz1X8X1oT8FeHmm/
474KTFS2L9HhKVdDqpItEWQWMZ5A6jCVTpxhsG+WAf17whRnJNcpeq1I1xUm4Rpg
JfdTgYBgKdnYwvnMALpWj+AYcLTnJ0ZusYh0oZ5MGQECX3niGr3kCkOPg8E81S3O
qHsCjvOwH9YyPYvoO+HTTWDi5zZT8Zs5VDOeUBOiocb+bFiCptpctv5Fyt3Gazgb
Gz9b2PTIgMAE74MVijciEyVjJuwWp6o6QShlrONali2xbN+a0+z0V2W/uabi97sL
MRc0Fqphn9PsTXZCVYwryJwSKgwBrV1uq1O7bYEiJDGhPgBDBSLwhoGLKI3vl91D
0wp20onEUPFr7dNDW+E0Pt2wLavhrut3HRwxb1wdw4j6wnpEFx8O+4nb+6e4bCQ3
n3PXTugecKpcsAMGK9/BGXsSi9WH8cs3VvRUN4L7CBcnbvLYXFKdXDkI9oCoTrRT
qMr/+hr4FQHzDWnU5izXB2JQCNwtCKmVN91bLPvLnlGvqVw+KZxu+mWjGIwqGJ+b
JXxmwB9cSVAZWvKQ2cWIdfPAdTPHQS8dooLh9VFZ9ssG2yr6mIJvOIwmsDIsTcig
CoijhADtyNGhLuMjJsd+xeooQHAUd8He2z7lbrq2ud264gzpFUkKcYG9YThsiBd8
7zgVf0MkyyRI1ooX4X1pADtoplW27ZWsx6O2zuPHnMQ86BLy6HQ+m5HmVIzCbg1R
vD1J7FR6LS3pCvaiPsI3kPCLy4oZq8Cr4sEaSJ8TELAjLjsA1/HSvOuoazL9b4zm
9UDwTUX7aTB2BU5+IpfiJf7m2PKBkckHQLjWdYYFzHsB3l5MqQ8KGlKe6oElmqSw
U0e6ZV7AVjEI9uug4m9iJd0RcmWIS8qs2oNlVbTYggBPaz+bTztyk/PvJ58INFvT
9XwfY/8dRRAKVbY1cQscjoYpq9rw+bXQD1GJWm93GTdWbtArEGTCZKne85ANalqZ
2xh62cNXc36WIkqvcYadZXJgjjYUO5SxUolp8QddpehZsuLrnTc9TnA99z87FnbZ
LEQz4833s7oTsPxzzQbyCVzd5AgRU+9nHaIGXeS41pQx8d3plA5yfUlA9WqSxstr
P8XY+CyBSN7hu61C3uCXkOLAByze5a6sveD9dFZNPyd2FE0QG2LidLpmiC7+jqcw
yeSiuNMs+onRysAodLIEDWZr+CpzehnyvKOUX21O2T7is0lbwKKBo0DaoDembJ1U
x9JL5OPwFRyydJNSLRsKOPDbBEGqDmox1dttSkjfnnZkZ9zwpigXsrJK9i9eEd8/
w8PnBd3dwOQqD0tCUjnCc8E20J6mv6ED3FoQhAzb+EI7d5GMD/YACKTnwRyM2VjV
T2Qiv5qLjGT8y6jN0yms7Qy1I+pSCQExjxFQc67bOSzdnGyDd48B+jvrHOHegx3a
b09cZMhDOjpsSbwhPl9MjTWrIBcP8GDWq9e5u4ScXk6kvbFk33eKd+Zma1dRPf8J
G6qoe9ivFPaR9EXriVkTzIEZDbbS/VKeINX/kkUuV36kAZ/Gc8XwfjJeyrV4PgiM
6XAs8HyAfbfVzFpPmd80u1vQ9zXngXyK1nPpa2nPap/bCFydwCy/LaX/WJLAV+iS
rVaJPankSmX3q5Kni1BFvN73I7PXCBfIMiRtGdPVo7xyPAQpF0yb6nRU1oae0Ik4
93jIvh804Ygl6nrexyyAD67T3j7/OqWoPc+JiW2ts6D9YnSjJVF9BfrtinJTrjtu
5kwuL4gmZaAi7r1QxtoIG/b1L2nTw+MiAjhNWyh99/1jMXmOAnCZgxbbm9doVs+7
JtJeHkgEacVVgE20vnZD0ZRdQK6HsITkSdIMcqs9VF1eZ+nGEGi7CqREfJN5tct5
kx7JdLGzE/TwG/14Vk3oPPzpi2ChqwR1XHeQkSl9Jyuk2KD2qao1BmTShd4d2iEc
s9bQKOK0hG1BpgkQpRtVaIAnf7RSe+8TyXJ4XPOsu7GRQuzj8Yngg1W+UzTA/i5W
H7t++TXIw1UGIshQ/FKEqnyk4h4xxQDO+1ftB69AGxZliOc9kVM6xk/g0L1oNG0d
e9I6SavPP1x3CGot78Igq0Nnqj5/fRG+JpDsUT5c/PNuXvQfSag5szrK/JN0qqAV
XezizpyfYpTJfN5gxe9ZaGJeYkpnn16yed5YmcVuNKhZ1ljPOQh0s1ctpeqABwFn
JkB9HIMp6/8/Ralnl1ARjSK+8yUTohvP59Q9psWZpEJcgOaqoFLRNRC7JPWAmlF+
kXQLYtHqjqeGqN3ai0YabzrwUAkgsDyAwHEuBtM1i/CS1wdUxnuB+cV3u5cnAX1t
F8IXiCwjJbgumstf/NWdL+st0/CNOBW6zyWfnBGHXIolwRV8c0WwpKfYCKQWqRkt
8XpUtQ+8kb/Mbcoasx7VA4JxGIF1i0UMywQqzEIxtIZsAALo+zG/c8wHL66uqT9i
msiANVnap/MuXMdM5EQ/TlOzVBozCjvl9wJOSBblNALB4+TNzqB/eLq5QVsf0fuK
l+20FSqdeIPeKmoD51RrM1iyX2s5SiqFHJDiO8uSC4ZBHfs1hrOFiY1hzso1A+dr
5QQ/8vGtI7rt7pAx72Y/r6AG9DbJepZ/MbiNPymkB1n1x3gS51gsyGJeWdI/u+Ih
wPItujDY3j+5CYK6QzOed/Sm8EGgBfc5dkIs+JFwKwX44MXrmvSHtCFNXKheyUHe
RsnwJikOgT1BsTF8RZ9lPXilJl5QXOuElwSMXKV1Mbd6SmynVVMrb83FsNGmY/lr
qm/NzFRJTQ/e+p0lFTurKny5l15FuwX6oDl1W4qbCaRGpZPXNRMFd3gWLAy77GN/
dbaPYsAZUo1oC3iiqTRZoE7fnkHMDyvs6beO+D2aSFdDUGSr3IhfDg8RUyYcsANY
XKzVPa2BgLzyJYIvdn4bmSsjLcXTFANognjUF7b76uS+PlFUBiFrLKU9CLcDTjZ8
wYOMxCND7Iudd539dXRiCVOM8WBZJZ87A7MJfK2AobOj75SCqiZnCG1bMTWdS/t9
WPGOtFQUPqZekz1WnoA6DIORYN9wNDLOwVdUodDV3Sb2QC+rNXENWHuBQpGoLJST
JKW74GOSWsN7NzQ40Q5YW6AtyZxrmHD3Avx+xNsJqgeSFBKv0cj9Dls/ejyaMzml
JtOQxbQBba4v8ShrEkrGFf0xeY1Za873RHMLU18/vEeEZa2e3BEuGKCK35vYaHza
n+s+64otPoMWovGBEfwNtspV8qRrLSVBEhWxwYzzkE5xQYG9mn+AExKkwiLkxx7U
Ov7MmRWPob6FXoLDTp9OeT/D21gMCS1a6+Xogxp6e/PEaJFlZv+htiTXRwngFfzC
h6htHz3XT4e/C0KWXRQzqnkjLjWjXQEMAP8EzKUFENnlMSb5QrTx88CyVpPnop9p
FX6YaA5QXjzGd4yM0hkF2lObqskcNl/dgsL+5LDVBq6QNsteWhrw84U3oLNeTzwT
mWeDCAAb0QIZAP8sEvPSgeFuVVIxvdr7Y1mFho9sX9YGpCh5msZI7paeAMU8qObD
CryC2LElS7fjkA2XTPCIELvydZC6wc98zyirsuny1FapzxK/z0CWOJ0fo5kShV2P
+VNxH8APXvaGCUuVGMa3NU9EtRSt0b9kKE1TaBIsnz3J5b4EB2Fc9zuB8iO2zaeU
yaNUjCiaxGkAAsNCEZFxcS5YPFAwPrydaXuM3bvT2hMAxmuNFabHIXX1oIrG2fIA
R9w4L8vWIGHkHlp6CFLFCOA4FMWFN6dn93XVlNcWpcfYWShM47aP3KNQKaNcooC5
KZWESgcQPUUU9zpP12kwjYbXtz6WKjA7+ioC+t7b/CmRD06MQC0VyIJLR4RNOTeS
RA+uTOs8fwnrabuvUA/lvyXJDGMcKBIBxcMvXc5hsB9yBtpvPoPdac8tVhw92pRU
VD7XuYXOqzTTPs1vxprij2Q7Te1ekM4Es5qtpaqaHSbri8uUxyjQ87wV4l9TaIe5
k7psz8AHaA4UvZ7Jw3r4joN+IAdaga4e5NMzT79AUZQ29HwlyzYNfhZ2QmGFlROZ
R+kLl0bK1I+z++P2SkN+9T0//OI6CWbspyAJmxd3tQzcCgGHBoVMKnmR6509mWL9
KV88gLNS2gSZTH5DgwQjAwZEz0F9P39K6Sfuninij1Z0+kF7uW+4jbHXHF437Dd7
ij/9gyWLlqvTYavDVooto3A/V6lgVbu/CIvGAMobDRLRQJK6iSiM02GLdr+AiuHT
M3jWbGI/hwJobWUeIIiie2/WDLqNHxJPwl5SMmvB6MINIz87fuH9N6r5hSecAFyy
Jv8nzMf/8j0wowVoVz5Xu2U7ZSvNrw82m48/h5gko8/fc29BYXdxizLqLVhMxj9C
U4yxhyjGB5pBG4x66+M5/CQY4VwVPGzs7i5g5urr2EJumNePDOfjjii6rqB3yCXz
xTWI2MdNtWplJG6Yvs+AZE2ooEe0ghp+d8z2JKtP+4PHUOyhjhYhqHkGDPdhnG5Y
GOpzlnR5oQuwZizVdHgN1LAbf4kETd5augpMNhyHL+Hx7pXH2ErONA2GV0qsdy8J
GT1Irw5yytXfJ/CMDfd7X0vZjZYiCwVMGY8kLl+o40rcgOzbdE56FU4aMyN1vSg9
7mLEKRc2k8BG8TFKHB78tu6Oc4Mtfx19bViOFxSZ/rWGt5hC/ywA+gkpKrXtIBJV
A5yVfit54UoftphrJRYK0klKyphnYNs4sw8kLBSUHnZp94pgckgBACO75KrVxHaZ
Uq+4XZ4KWhrKYSOhwAySoS1kkbTq9QU35oICLfkB3tpKcoR0J33G3oKEyslqJlf3
u2HMH0I43Z+lWg8muWMhpdwlY4r8XjNwclSFdMCZBbr14bXZtMrQg54GLqF0e/RE
u5Th5aOjg0tbqrdVYeKdHZ4FeNcJWHFQozo9qwWmzQMNRamUJxtVzA5gaU4R9DPw
LySzHOuHRqxrMNE/J/9atDC2a4eF640Bp/uRiTv4T80fnmumXqWrb+dvOs1AZXgk
Bl25TGZibKkRhPgFd6/kvZ1Yb2y0upFPNbvTsrmYbpUYmdbu5gB0JNDuyYBva8Ic
cX3gkfq01kFuQcYpNu0f7EPpSm3f5tV9sZ36gpwti23krMwQsG6fBW8PvQftjn32
tFmS7LDcDMs62mH3ywG/+dETKU32XXsfOoZA9HjXSYYkxHq+Up+rlFzGieNACk5s
E1lMD05sHGqPabuHT1QmwqDgmEKztGSrtaW0yKyfczGkarGbE302Vfwb8mhDQmoS
tvSPNSWvLhbhhvHoo6/T4sR+4Dp5nHc2oBqgN/u0IKa8ZKYDL0MeUSa0r1VNj/Op
//vm0T99bZHWESn7GWWnjso1SKcV9FlVhH0ZIUJqMvyhuOZacH9JRCVFjMp+Y+97
bBTuZtQXXQOILLYNfQ3S23+yxg72oSOBfHW1ARLj33Phls6z1zSMMZ8uwdrw3inF
JtyRL+BBLfORgjNFwYNSGSzN6ELO/X2QvHs5ESrJsZlLUmp2LfBT8xs5fSTrRKzR
TeO7AVSu0QWX3GC7I9vpGksBiOm9tlo/4cPqiIVNk+FK4tcLitmfVJsUbVIxkekn
W6rafgzXIQavNNFfy5dpmWr1VQeG/s8J6DZjLX+fVIanpBhlQ7GWptW7KtQbbrC7
asYW+D/rgsFtmUog30o/GWsqQzfhGamDhQdfZyGz9w7tL2I45JvEL3E6+KdRje/y
+D1CIqeUXCgbH/aQEkunIEsODez3pI3+ee5K+dWJbvI3CMMFp4bZ1pVn1QRN5G8V
yxVNJlU4nNng+RPlrKRk1AlKLLzodkAv37zRdrpIIcdKuuTqG0f7wf6Rv4kmny2C
9asGODFuE7q2rPAhj2fIgeTl2HgYFWkBFWnYH/9UX/QN6CVyqsRCndeEqVH52mhO
8K/KmCW0FoV5lWCglSOfZSMxtvJq/NIQGFTcw9XA+IBhHVg1/n9RQnOq6JmDhupc
GSZk4f55eW9HSoxsegM++p/71lMCkOX7vadQfOTfrxFgDVC7W8sbB/mwKoKJ8U4C
wXvxj63IvXe2D1oPR3bFXzKTHkTSYHJrPkGdZHnMQ5GDNZkexOoJRBnMPvWQveZD
ppfVMw//51738roS0cnlJWsklYGnNOS4thVSu8CMwpl//SMn3oMqUZGPuaWDVn9I
Aj9BmE73Cc6KWztWTD9VBNPD1XiBDNjFnHCYLrJJRbPiMJdqakC3A7aim2AzjmVl
20VMSFHAGnuK8zg2PSVTL9Xxti0AQ1AuGBt1Z9giEUvl8yXakX2dlRNu+gVRCbEw
kYJYlU1VbntQBMYyThPRNbcpg3VXt7ypXz30hnTCNMt/Dsx+cI/ByK0w1EOP4FL1
MdiPRoXmvbxlG/yQoif8hYY8hskZQ1QA72lUtoVaisv+VGhbzRMXfj61ogB4EaI8
KHsiLg1FAWPxbkFF3cLRWriZD/2JZ+daWaECnrSyrITVxaL5cSNUlq3lYrjP4J3H
ns8zglklgHo7aWZXeFeTUT/YFL5yQ8mSW7msgAIsUtq48rltZgiDP8LUSbnTLyT+
3sCzkfuC1yuA2Ej+cnkfnxhygDB5Ays5iZ8QVzn1dTAiuHVwEojS3EA5Wel8tzjA
Tuv1SJ2l9PrRX+8ngJ2MUq+T+N2+rT4EWEdafmyG3XhjzicryyznND5W46tvyyyF
rkk9O+3KYgeY6NH/SEcSXB8n30O1D1bDp051zSdP9FJj+mgSAVrXKUKPcj1f3kel
pkqG4005NxKlGYeuSQ3448ln8YA1zmDPaVTAsxk5CVqjZeFch77EJkyTJtzmGn4V
xSIJrgkO4FyIUpBIwskAregDOA+Ag8P7ersGFOwQxY6zl0OVFU+6CVVrlEqAlVhz
URSNmc25iqKmD5d4Fz5xBnWCEDBZo3goHCLeqAZkYqZQFxqITqQiYTrTeRV+h4LG
hI4BzwBspwCqK+5Sj+VStl2zGvjJSb8PWbQy4F4n/eE/TSbTR0VYP0IgR2Xccb9f
MdMQO6ikK6iv994QbVqJ4r/PLzUghcyw2Mq2Tr9ylyf0Bpdh2OCEiPynPLd0iSU6
YK3Nm1vhfl9OG0DHz0XKEcV7avQtmJ8vCFAHwi8ALo7/dNIZAbGgd1f87sajL3Bl
9JuVLxfU6/8yyKlPuhcYSmRui4CUGThbCiHU7zu4nMNS1NeutzYzUpEFyOOh8Yau
iaROzkXFCpwbA6UByZMKeq2xkvk38XepitodFwaFrwhDbeaTksYFrOrKeUfxDBo/
qhMl9NxjcvWMzfqxW/hSsbhCJ9j6/xBWwODSm0hziy/O8RNoKw4onDh3O5OE9fvt
W5jlxk2K6chanFeUxvT4nDtImXpcaZKmI4dYN6xqpTrqZOrRH+Aa/qJ54ZHJJWnA
QVxRDnBA/6NE1T2gf9PCgDtu3m5msp1Rn8T1jKaFZcQzEsGehZBgi5K0ZjSage+x
s4T4W9DVIMtPL17nWwIwz5V3pDeuGkRhY0r7gBg/4mdBHXjQmyFON3tBhqnTT5HJ
LYNu7v3f0U6VACDRSAkd0VYDJTeA8W6s1nAF4McvEefWNeOPKOSzZDJ0U1NBHAAy
J110g5DnceIOzEVoi2OlalVF69ac19GIJDjtElGya9q+z+24p6yeMGFl4gGI8bTz
/Sy9AdUJafpVuPOZPWCS/mqNhXbppoMP8N4wsQ49o/b3AuTJzN6TVehzZmrgvKHT
QtwnefBuyR1kPt1R8diTUn4LXNkdyMnd99Z7KUXo20pm6MtVanIJ3tU6gINsPmUm
M10l3aSvbN/zuQNDN2z9Fi+vkwylidXcJjczc4KLN/XOJiROE7wX0/DZmk5scbuB
PVRTy0jwibcpFck53FIcT15CrJs10icM/7u6V5KZp2fZnqBktDoHBU2TZfU+n+kV
FKp3ojNfhpjUZMCNuKwwjmLdbCH7XOz6fOiUvmqMZ6zUXmeOfIMMNmVSWAUca7Ko
eVHbVfHs2gTkUghvKo/hMotZg3LFxwVzemtlh4OLUZvuWxr77BfAvgUkKvPcdf4H
ToQeM0dbViTqBAXCiHuZ91J3i6RN6DMlMemnaUB0BcB3aMXG0Dypfr/wQgdo6W/p
/pG276N1SRbkboqXDfVoTNYyLF/tgZXrGAoIur3E8yurJXQYA7utTrkV5VH/UUK2
zUapJ/VDPkb4CNfJRNx05FR+tZuDiS+Byv3hJu28GtCgR5blWl8GnD98lzfK8S/O
pAiOZfPT3cbFG2wkxOIJ06dZE2tlDT7OxtmGUu7wzgfg7KmcD+68U/icPsaBgt8x
muZlIUt7LJo2JVRZ6+6yqUq72dT1w4wKQndO/eXZnrT/cbo2gUQIH0dwn/hXDTao
e8ozFdZ+sXQsi5rBJ9gtt1ViBci8lNkXaJAiqi5ngZLzIISUzDlT9tEBO7v8IRsj
GmtHymrrAibwUmmiwZ37zM1eBdQhb1SXuW9GkfzPrN1UwTXEMw9nWL3TLVHr9j8X
3fm26vFQNmfpeKoneP/OlQHWP+npOdtgTPoHWJR75NQnyeozd/3aM/qkF8VkIZF5
GAZaU+YdGwQNS1xgZJUu/ZC7Rr5LJkybRgPHy26LdDWhCic7OCRyNi5tvz4r2TTg
mCiC3mUe+OJU62CbOQ4dvP7sXNjJzIm63ymCS18TRtwz8Ar+m7OzF7Nsip5Yrsv6
Up7hwVeg5DcDkq3MgOLG/PKrv1lPDKXP2u+iXAhjqTXWUv64kPTagBsXaqKvaAGb
W6I3kfGYkdvKUqSqTexnP5t/WcLR+SL0D6KpFBoJHHzc5OQkObe1Nn3IdnFcDYBf
aBPcVOAMZRmLppXUyn3/2QIgSSba6+wQNchvxY9WWwCcpVmiWkGYVOg1ECalK51m
rLZ9DUIcS0EEYb7Ni7FsBA6OqqVwEiSnQfmceHyFJPpWaSFnN289I0FTKKOniPs1
U1fF4L9q5ljejQ6Udz1HuEftIA3U83L/nLes/Gnf6natllcmSCmGpgU1R9deGMtl
8MVauBYWwjZQxG/O0wTuriHiY3wBp39UJxc5gp6U3aqG4R6l1sOzth6nlzfwvMqz
ZCoDTBcGvid/oLALY6W8LTU+agP3g1ObcDu0ILSEHiehepLAmBHyjg77YiRpnVYa
fIhqH4TpCeGTmA0FOBvYVLYNLN+LYW/HABw74v8/BVThIj2Qw5oUYeCZPZxTZdHR
NnCq4pAdUR1jp9gq8gzrm/HmD/KB2kSD9F79q/42KQpLLUL6Uc5+tZXs9D7Q2KjK
GJlc3Tz65sdITaFQgPTLmPQNCrqe60e140AhNMrX0lFbLRrKWf+PkUCRBlIqlLCY
oh3KtUpR+VqrONa+cB0mpmRIMmSX2d7E0qji8xxl3RteTlG+WlsfPLc2Pe1vflpM
VN8RXJi7B8ZdInpd9ez73I2D1Xnf69lAbc7ZjwDHirqaa3X3YG5k1dhQDJhQ6M8p
3hiSEH9/PgGDk/od/USv1I+ptaQr0O/MFMexY96kwR156cfowrMF7eea+o6XuZKR
+VJvz9fOBpM8oWV44dZpVWQKoeQt+zb7ap1bKvLffn9jFNDUvxC/soipWyZQVW2K
5BXE6+3XRQcv4IyNsoJ3WRLIUs+MWFYsjbvm1Q+0gmWFpw1WMVHST0aA3TI5pBVT
C70Uk6T3cqz6SM2RLBa1O26q2PZTtUHmz6Tbt1Lq2gl6MfHT8hGEf7RdB2ZDN24y
kTpuvXk1mi/wdKJMgc4n8nwnkhQW/3XHmGfq96gnSgFqzk023Vcj2s9Ng8Tygj9Z
c7ffVIRwFxBeSnmC3ESdJxqIEtMCsswaCUX/52vrel5+Z6BZMKBhYZ7GLL3w/GLh
nMmtHvswyWe6C+wE65OV3QlfVOeaPOfi3elWFTT252b02W+ljWxDmv9T++147TrK
8T5qEVmV4pXsKpAAJ6qsMtmyzi63ILCrmHBdW9wB4cHheqx6ZQeCQWmXjRpBx1e6
bOi+2ZbUpYqnoIxJy/s+1kreJfV3G8Yz4C8/8jk/7+RAPjKp6FygZMUPoxJ53LsP
Yk75h4nGshA5NpPRzCLXgenP7S/lCOyu+iO0KSZqYMyr8HP+IWHCnwUq2ACTeoLb
NCakLxe1NzgwqvTqmIDWbQrgQ/NXExRL4oONgheO8/mBF4J8FKcTK4oZa2R7/h+G
iwtzouFabnRn71ksenAUhRzhs3ayBnKuexmiwqV6rKyioHguEBkadxWUiodDFy5W
dSaAz9Wt9vOBhPX4dnBCqOf/fJXoW+o4ZD+mCKkFKiS3ECQSIOsV5N1EFcOttpHi
9tJWRnRb2I7IAqqcdN/VUw7MK8BHqHUmQPzMMANy/xeJFZTLdA5JgvIHb7o965MJ
WcmNHXv7SY0Pai/XYF0PZbkHM8s1uCm7dSoS/e8n155o4IKc7TQGhPg1zrwhJqIo
/kN1mYXjGOriW5r2JQ12xN/7TWqxnN/Dfc9uBNIYCAO+KKgetDEoBHuqfpG6462l
t5aSNLJHSsdhTL9xajdCNNcFK6psvFKleeTNevFJoafeKIe9MJrpbGz7213kgJwD
r9W3vM4IQVROhYDo/fsvxXEg/AtveXguOKmcrKFq1YQZjLJsHuxTtFVM13vP9Z/y
9eOeoK4GeYDq2fU2l4MJx19IC5sTdvkXb6rc8YfvuPH54qFOf97BH6zcsuZkeIBo
TybJETczsTlmT+HcNYu6DsBadZThLsS+giqaFF1fdKECxYzLB3FlQBpy5AX8hNsc
5rBClat6eTH2IdhmCWIgrFZiN62yra5Cn0CxqI/gL7xntkn5RBBvQk/96QBXeRrh
9ysI11nPY8FRDeOE1gZnuFHa39OI7UteEkx3Zs87GfPRWOpRI2TnZL5uhdtEJsEZ
6Nu0vwwoxAPH8908WBWDVGVzkLpkIGxhVHDMv1f03YnKPjpE3pbtAMvgu3inKWhI
SjdaT2SE+ZUiUNdC6DUQDf4m1KA0QDT+JtQkS3iUvPQy257AaEqNAEppB1oVUri2
7aUvHY0K7qEBd4uOObWA1V2LRIcsQ15IBdCGupzluG9LPHJD2oyRUHVfAcewfTX2
30v/QACzaFHjFBN8gFP9hi36auK1VddslREd48dSzElrewZaIX8P9EdE8Mo1UFSj
m4CxYjLujdS0tcjZ4nKbV/eYDz01sxiijFc7avfytA3EzicHwKmdBKoNQuEb+c9g
V8HzwBy+zoFPWdQPdFyokThLAxQ65all+PLHTOMvnpIujNkVYoItKHbGLHSgVyGd
K2+f2SyPnQ+/QL3xrrcWblJPFpwSzfnm83hwlDDAGoDVz3OLq4cVrou6Dk8qgcLf
XwDq6UvrvAKJs1kZ3Mk2GZX6X5+DmKlOhtY4s5LuyJRF9ArK3XoZbe0R9cy9jGlP
+EZSbs51vQNkOsCJK/U5pv5i/4FfXf3hLfQsp/qJZ4R/Uu0srplSjOg0J+3xoKoX
iWesG+hC98FieijW8OdR7o6XRjZIurnh2GQjur28C97MzYp5r+3o55B7c65lfISN
RUqSacHOzKVL4qp43byn+X6ArphHqCokZFk/bXOnF5xa+jdVAJDlKx3WxNLbWQIz
P15fX6MBkYYRoomfVla91Vd4j5YJKGEuL1pfR+ae0JFl9+gigfHZPsV6ssPjP+nu
sNKxyYLplDelkiPjcalij1Lkvxrck5sFjCa9ulKswJhR/pkaHyvIgYcSrqIlrgGf
kU1GbCx8SEKNRiaXtSKjCKfVboYlBR/gh7K/FkQyrTu2ucnJ/xwuL9CSrCAz6QhD
d8HlgsWYt2v3f1+jM4r7cint38IqHJJ/QQ61Dza12UVqxeO7Ou66lLh99gTzt/OG
KbLTYzjz5+3cV23peQGGOeBL9BW62eOwly3fqCgaOps/xOXmCx0ANHfggeQsZ3r/
GA2gK9weuS4TY3c8QxJgSbvi4m6oebAMVWa2iMNs0USQ20C7emfMcrcmcmV3TejF
raihSU/tW1iTqWnFhgFkB1vUtNp3HRcLKf8b4tN5aPToaXVv5lc6jrbfvFivdK1t
6VKd/u2ej5Hs1ryQ4CyKMXlxX/vGD34WZHqT3sQWVLNybToFB06DHvUB0Ekdh1L8
WCCy/OW/gAqt8E2+DjQ5v+HVTKn5aicGGPOLV8Lfzwf0uqkVw1wjyOXRNGBR4sU/
3Bcqu5VvitN17zbRdXOQp7SHJFb6ivSzA1W/8MWqZcEq6EFOOkNKgYx6YdU61nwb
ThhvX2Xb8H7aXXMXdNyE9nA3RFs0zaqoC3eNnUaznYmym3embqv0qOD5+Gii3edr
tzmrR6HAnfof1birOWUBfOD8UYNRgym8yXanEkz5U6Z1+vRLxhLhysomTraUfF9E
WqlNiIuJjyn4/SRCpSzm/HIZ+ygDf9hJWmKPTNSUucJRg7QLN08UbzWC1WMe5bQh
dw7ydm/3XygFp7m1cGzGKqySThX4bbNJkEgwQH3bNcww3iPOS9cGIq7048WDJmv6
LWYUu1aDCV9+rSz21wMcqSnLLXiY82iUaR/NqfDCNkK5uqcSzdZcg9K1CKniwXTb
5zIcAF6Yy+Pai68wrwEg+Rx3Q2/wJov13NeNFVr8aF5CdMkoF0DW7GrCIk1wpWd0
CKpruyrIEds9oSvglAFzfg02Q1d4SjEfH9/n0S0ihoA3srATj+m6RTbBxhfNJcQ+
VMmDFQ+82pFLXCWtF6ZCbuBfnGmps5QkU1Cn+K/TEOZzHJoywsFGsj0ec/DA3J3a
3EsDpySyQUMnblOTYgbJ4C/1edO5uayeeoZAvzyXq5l8OWMJwDAsFA/flOgAtwI1
iLOlAem4QNx9x40+lChxCQIlEjZ4pGpGsOK39JoG8IaxuBPdn0OZ3gY+qoLlpCuG
kzlutfc+u0B6fppCbHE4MibXe9QfsXD+JDvSZEt+sPkQ/9bggM+jx9Sjah+8kcus
rMljeC2vPVLvOdwe9g0h6nnY4lILeT6x5wlr3pb1TD1yEDnlKXqLWetWxH3Z0M6D
jFRc+rvPy6znTQyPS2OF2pNInEAz9Xw3VG4v2wI/r5FKgJenYaY1Pz0rZQZR3siS
+qSJBe0qcHuoxK37KdwKk7H1eGlOHRqiwZTmwV3HSnQikAPuDdJx7GFrYnQosHrw
6S96GmlK1RrfkhVFh3eQdTRyrdrVOa5Uks8pmQv5GTAoi0/foFxY25r6bmH0DyQx
ymh2oHWv3QxRc2h7sp1pqysUTpUZ2xy/0AYC2BIv/DJWBmwkp6zGj7uZRXa4OAet
+6XLd3XXy+pCd2fQeY8ropsRq7n3zBglgxgCi0wky6oR5Nh+A1YSN4gcYV+w+B+n
hnQG3LbvdWTAQRIpiKSqz5QwAvT1tv4z/50oWIrXhs+6iwUggSB7ayl6rQYBhJ4z
i0/8TPWuRvOPJiFRKUgcjTwCferkxk9vX+POTB6RzDfadhgQdunNighKGByVKi4L
KYg23zLDShKLu/7SllO1dOL6kaM2EMYr4ME4Q80UmprCCbLEop3nonWfJyCHJGM/
e6ZJh4UNgGJAzlGKAdKd5tx54/uSXBv//TkMI+yFiTThO+SXsrlPw1O1ba3sgO+Q
ppj1T1Cco56b7tcipRoOMrr3IwZwKJ1bsuJoY1egcRug6rD8ILDQfZ2qti95gMvg
jXzYWFiGZgq9G/r5SwZPSYqv5K40KgewvriX7INb7VDy96/YIvseX/sHbynpd4w3
SrB37plq+6E+LGTyJxNKPXJy7npidGnCnHIo0tiUcbipVWi2alY/J3/85sty3BBr
U8SINsk43kt3D4BRKJklQbR1oSQzqhm2iXc8iG8emYxieASLWVYYyhXo+SbjAwnJ
V50WcC1yGYYngAOahO/JscwFgid8NXiwqmiBEYq4JAqoqxulGKYd01T7oFVtcUj/
O2fKMUtgar/JJAMKbKt2pRkYfc0oPXC1o3MT4WW2bdnPArolsUWZlv9m46H79Pnd
fYNdmzYFP3Mg0thBSZAk7hhmAPrz5q80nKmJXocNLgxQS8NEuZmn2cGufHWvC9tU
6XgvKPL6x6Qw9tzyECDzOkXABJUiAN8m2GwmFczHyKIQo5Vm43e4x3AQNZHJn+wH
SSvCc7WktAtRlGAp/qxdWSC5tciEcWlN328ZOufmBMNPb+LYJOclXIcrPDNCupFO
IotcrjTt3OYfHZBmKFRGkGy2BcMWAoH7Kj6RR5FGSA9I3JGuHNq2gJNMGmiRSk0q
AQ0CTcH3NJLanJ+88McTm9umUXPds6Md+rCrBubx6jqW652YwbL+iSqtZxPYGR7k
iIjmjGZjg58MfwlknW8UZIympzA31F7Q8Ld5mABicTXSySEljan6K+uv7kN38LGf
0ag5C0r/JPEMW0GZJCXhsy73cfh08HYluyQqGAIp50V0yT4blZkgYhgHzuTKTPJO
PjuWgxHy1707/LSSE3O58lsnYbLeFCWr3UzLdxhYzKafGHghOV59MTw1EwM7UsaE
0NWCT7NabFmrpjF8Ed4RKvNFVpQw6CMuzhelXIOLA5h192CqQpPYS+3L3k7AEHL4
NawaOWqydNosNMG/RMQamsiyv2TbaG98cG+DjpavLfuxGq4kKdFaxwIzRDDaGJ4t
orAKUw/ZHI6JceKI3SZFXNrpnq6Z8pXMOYaphBqIDys9LAvwq11oJobxou997OS8
/mqtDVDY1acMpNqFsROwinKjZVsYt1ubeBC72gtSq4FgTbG040RwR87pZjWeFuOq
wcKjDH1v5AOwuGsaOU0eUbGV6Ui0cq5iThu4MDo29y6N1TbpfTXgMTm7u29Lf7bi
1T7tknhokqWl4rkf+TvEV3d6cNTKUgTFBG14YuiDlaWIk7l4fnCzVaosmuV3rIdg
Bb86Zx2Xn9qdDy4kLxr7nDW1i1x967rpKFCAF4ML+y3ujAC6jXccpwU8D8SOUF0Y
5ZGNf4zcGxpnaQDXYeZ2L81gv8RGF3GkbY5zPFoArJbYMf77s7tFhy8H/CWNsTDx
DzVbq2Uxmw+bCfNCW/Jh+EF52ho4H060IfxwprmZ4MwJQaZIy3Mm1qx+43QxHehG
lVE+jsc33ThfXlezkwbbrXkWpyZRcQep/BPnVIfsQv2ApNU/QYkyPf1zEBck4vZ8
8BqiLYuTV+PHnnD17NbTqWDZ6pX9EcicPKqBLaRHeNark6Zq42e6jCwajwSlwjXw
aMJd9dvzJzxis7vI6icUrowvPITw4lYxtYG6+VXz2c69ZCsI9DHgLAE6NC0h0YSq
NzxZFZs8VSmX1qfow/654dsMqpUQryLBHNiHVYNC4rTz649rN8ncyZ2ZntrKgmu4
5Aqk+xoqOPjnjG6QwwhXnK3YujPp3CwmYUuHaEvXgd4ub7iw4QtOFadxgPBeWRx+
SuQFa3I6gPGcd36Jxm/rf89S6CUbW3EIJNX5Z1TmkBP3mzuiyV/95wV4T+T3fbjy
LA1WkyZh7nWDn2nn1psJVHeDAOwoxtDb7i0TVz3XsgWz7+iPn1HBEUKqZlQlOmg7
62fWRQCIh50QguVaYjehG+Kgz1LxAS81vhkDxDewsp2fBT49NgyzgCLiSXZ7lJTL
cUa0ulMcUAeQbk1rQFlvHGHtIlrIOu/xPKgjuL3tuscx9I2qxCbGV2cRrsrx1E8s
OMK0i9wZNXxYvO2Xe4iUoIsjsU85VYpbhtFa4K9mKKKohtSQo6K4ml0wi8VL5T49
sIZXcvHN8otvtGKMZOL4gw4ilbUlREPyZDWZnbzkN08OtbQLvlyU+pOTQKrQxWAh
bG6A5+kxt+3SWRMseovBOp0JZNRBpI15S6XQwfk31OGcE0obuqUiv0ffeT+k4d5I
ZhFAM+/IJfO+91n2LQUZ9DVQsiTtxP5ca2UOewFuJLRI3NdRehr5vHbP4cHizADc
mBK6QSFw1zwFpI4/5xlxjuUJdMfm70y17YLNoSflcEHSP6U8GPqBEGeMvSAou02A
bgSiv9ZtpYhUu8m89q7fQoyB0Mkha97FD6hpu1PZTIxpl6QJCVWMfuoU/N0NS3/B
Ncm2qM6U+dYkyfj1qxA0/JZqIv8m5OOelLqiJfLcpgxJZ5gxGZ3lcc/+FDEz86WD
L7oKqeC6TFJVymjmQacZBi62mYVkOpyZEIKQsZVhxdyCY70Ezu8GNY2a5AU7Mj0U
rOxWP0uziprEo5kekSrdu3qu9tITOHYeNqEs3amNxLf9n1tWQMdrnrtkHRALGPYc
8w1iVoZKgUhEkGUfZ3svdSpr2BijuopYoCXLKc6rBwXhQKJ+i37X7IODbTAHcZ2f
X9g35rrSKlx40yOmNoGMP/TLm0UeHUyi2Ck53DVh8ewY1iEerXubuPiQkzfFneUJ
OEoPXL4KdGPcPuHzOR6rslIlIORotncCslQY8B0FZ6/LU7YekY8FwrzXpPdt+GjD
IteCpp7oiEJoixS3a3f7E8T4nwhB1H5RPc5Gb2aXUzdMAfFyKgOKczJ6l6q0yRHd
ohIO5F0Ba4nadByphWOH0KKiTtg/9k21OpZ+rTdhx5Eks4cAGMpgXqmogk5yGArA
dAqAvzL2y5jPqYQ+O27Uv1gV37uaet595/wWAv/5XjC6zcsVyEzNbWnvbTHzw/QG
tRwE098WMuuqmVZBo8jkcF2Ej17dbHtgKb4OdoZnCvEUUb0kuVzuiAhStjFuyU9/
SgrzBNULLajeWW+FPemCgGY+YtgtT+m0uccB8HqtDiRewGsV93KmamD3EUmX9pAA
/6bLBdLaPsXCnIwXNJpzNBGJbaNjpHZWu2MHvgHBJ9m2iE+meD4Q/4E3cgNfLKDw
u1YbtfMUL78SN5IEA9VoasQ8Q9Oja6uVRSjqk+NxuhRJeFdRNpPSZjZSNxbyjjbV
s0ymtbBExuApw0/eOh5YkZroM+5L3Adco4QldPXyJf2jCb3E9jJj06okfOhJWRud
6odqxkBL+4ADkKy6rdRTZqMSFTekeFYv7Lag1JgK9qCjhE6EpvcpMDIccYpC4WGv
WAjSCFSY0H7wQF+Nl+qo2JnCOROpO78Gv/4/zZ/+5rPcsa021iD2++k1s2JHJhIq
EC5TC3gwYRJtvL6GfTboKLc8IVTNEE3sItPObLRUwIOBM+UJF0a6Qcx1WhUwxPed
MvQUdiTZ6vjbyOT3up27MBDQrPv4RZk9oadgwuiYBeseWoLH8OkVy0s8AQeBxCxY
WXFn9gSPFHiLKKLjW3BwtpMgrOAWGqnOAf3qJJn6TPMvAjiC5o6prsohaEB52eaj
4rBcZCUYqApDV8++HBHaahb164TdgUg/YSxDnEHUUdE1tmWGsUJrfztLSPVRZM38
z+VSbvwzVpfsUnaRkdpy8fmDEr9/YB7PaZJVv/LssxPVxXUdF4ocQuQM71kCYo7/
4F6ROugjZ6GQjEENQmdF09mlCu0DaoK6CTEKP9qdDa0U3uXUwbmwhwwOiGMp0Zlf
gPjZCrtj1A/IJgi5vCoIJI3SFSU21RqfvKomARW2mhNS9mpgqjoQo/XFxKfWoLAz
8ADwsDTpBm6WTS2qC5TQXpzGSOJ0g/5imlXV5UHyZGZaArWNteYKr772DqdAMx/T
ILTVayJHcKUluzBs2PqWJNMS8oCkL/og/E5Papl8rxU9lpreVbw4nPINsni1Igut
ZL5Svk9BMdyTBxzbb9p9epM//LUxT6DVIPzFc5xrXCz0TII2jRw3vjjStO4xd+Ux
c/EeYII/yLjWhu7PP/g0up3BF4u9Wd71+twRwncvd5bzZEJelLoiOY9iXV4Vaqh0
KbQiHE/JWf8/C1nJ2BYjVeS0quLYo0r+GveVyjpaFWmo2AzwRksRUBaKFTuhXUG1
RiK2+3bxm4MEZBhd7U/a+OEj4aqPmIwc2RP12D/YJC1iefnhvhur8xNN9V/TUJd+
tynFu/zGPJua7+QY90MgIvYadOyYO494KD9vWmZRVE96rRgWoZiEgQJPUHvY5pUy
AIPCFMXv9+IywzpyPmIAV9SuesJLUVT9WgZCYFenYx5uMXp3NRFk5ObrpgPhGcOI
kxUoVvTcVECYF9FTzClc9gzg39NwAdIyMkFxVdV1IPhOTD9wkD9o0t0Xpl522QEK
v83Z05b+6YMGPdfZNsw3Ixo2vs2Jni+YLqgaal45y+q37Ha0wM4V3B1vZR2nx1pP
CxivecBQGpcGzIdYohGCdcnQuI0LJcKMf8r+QRaQ/7MBXawPbXPII0XNQSAZ2uJS
7UE5aFp8VEgMdU7biW4ehsZlTlEx+g59QJcVCCiyUB6peq9XjWatmjx3VtqK1hQC
3jFZ+ztp7gBlfyEi3MmalAiS4AgYHjAoPlI7J0YWMP2o2Ud2q4nCwuwgZj2jFMbJ
JGkL1g93qj7hYkROCfHb8Oca2wkyM/FSctYrFDXh0mAoX36PNwK+xsZ3mEOWkJiN
wnC3O5Gj9vfZpD4ldjlDuIXxEszSI/PzOWg2SntFFgws1/vNq9XxVl9K75SKXI3J
TdbvCt1QlX9RVH8Jo6+VICxMWn9AlgvQ9AlLAO5J6RHpU1HFSlosAstG2h+qip2R
oNPOMq1F0uv3Agw2ZFNyPs/PIEr4Q/kv9dBT/Yf8aBPuiwI+kWvX3m2rWvy44GEU
Ph7tg87RG6fwFLcOFn1UsLUFP+umFENcIZzcJurU3T92tieg+An3ruKH8fIbkPaO
C3wjJgOl6WHdRq69yPsW6tUKrgp/46YwODQ3NcaOeqo+scgRVji4LyBsCozhzSMe
Lnbv6598fCbvJtYejplN/Oh4zSKzgHqzzAmHW5mj1KZcBvc3TG8RVSXHffEy3a0O
9p454mXuBfRHmf8FeJyE7Z73aETaAgF2TWzBtLz4wy6rsx0WEpIIFEMQffwQstCB
UrZJ4KGQuGFKCgOHB0BBxmXK+gAwyKqWmlVEEGTxEPTX3SMMNHGnq6fazaYV0PcK
kvJ+N/OJBtzZan6ZzYJkUtdKRqpHjFWYSmm1gztlNMkYltMQXG/o3KwbapCrg+fV
hMi9UEfDxDcLUIjtXgzKUs8cZavl1oOLmQvUFa0Biga3sDJNR3WQFEBxENbnS+Mi
E0jJQXEhkWmGCBhSH7RsxIgdb6EEVU5Yh9f04M6AAfraDYguFqV7EO1muC2DPeFH
CFu+igSydQl2+dJBP+zP72OEbQfP47WvgPawCDqfwoPa7irB5fh1EOeOEaEXTyJi
Yqcul25nRcqW9TlfFIUHDkBQ0plmharOiJrxc9eRVB12emNaAFcXLZddZi+GZTT2
5SNwnq79brbxpN4UmNiftDJNk8jbRTudKtF/sWXSweGxgaaGloZjYTeS9iNnIq1c
wpe7xyvFpEaKjWb9Pu6so4bUTXNZmOgn3FhqeDUV8sfOUJ7vSlYPXgC1eBqSA5a1
uXKYxtohvk3uevkvahLawjECk2DmWGLRIEZKi0xAKqMXnrMx6QDwb/qjx2pZB4c5
4/4yKhivsalbvoDVzdoqxIBfLppKr8hDO3p1SP7kn3wVgSymx0wKqA2vjYPEPkSO
0dRFv5P5W7kQymRjekFciRxFs7PJnhrYL2yHIKkKpdhAMhQ/Eff8TEfUptgHVrIL
o2mEoFiR0v34UHsSfwhMF7X5Z+SmFxsJXHThPmGuWixhcbz6XKYF1EmE6QaAraXb
w75ZStYuXl7/R/cVvAKaotO2NJSgGvtFR0MC9A8uB8DVRcGYJMXw9UFFfkNUyETs
vysTh6aQSJDpQ+4rWLgoQWPDYWTv5w14vttDmuLW+SoI2MF/G8vpkiNRrhrlabu3
7iYusR/QkJiNDpfr+Op3MNtEeQI5mPWStqSFWRxYQ/Q2HS5lughJCu1zhZBifvoX
rEKT6/O9z+6qqSVZsKNT8JZBZYBf3UlKRjXRc/1sukzBl0iMtElnvvOak5kaOPtf
iOGYzW4lCy72VYl5it3XLkvNrp4AzUjJelxLzuNNKcmh14m7sod0Rx/WHHjF8nZI
I/fXtnCBqfJZVywCL3O2fTOJnPoBnacl0Rc156jVrWh+FRuzT8IdVvAbdIzK9HhC
Tm0UH4w0Xd2rczPnaCOuHsSlC+Isr8HmXMnTG87lmM+tG/6xpdfFLjk2xEJThi1O
MkldJY8pjNRb7qQfuoP59LuEG/mOT0HYjOFDaLSC2LjvYSMJyCEcWU17A+i0nNJB
nQeIY96ktoYfbgcjESQ+nXyN9dnpMll7NrcLBEVpJT1z13JwEqXM5Ro6tJbRg487
tofgp1hfoS/n+NHNjituWyJl4lQvtQG6mpSqTR6L5jHQZLnJS8pFUBnhkY9i6AEQ
3G7sbjGLsFjgncwt+Ta50phhrw6wOobUrb/MtImAXJhGOCxaa/PrYPz6piuX8Z5b
ERAAvJZavu1azKkYUBliQh4qURnk4d4I4r7bIGlatynyYF7mg5e1tG6h244OCCQ1
8+BTZIsKtteJA441rnui+8qPW9+yVoVAn2RTTTXO+HPuasFLevUWgXBxB9seDtC5
gx71V+Zn/Kos+LRY3tLV+6h85JWrRS9lNjJhV4yGZewGHYDZR5rwhUiBQehqCyi1
Jq0QrIp+uOrR3PnCXWb9mNRkGlhq3VcYoVpSQnklpVrhDcTY6Jk38ZFF1ymtEL3h
HgFq4YgLPw2bURZAf2FPdK1VsLvGNHd6ZnvOE7+HQ3yoo+AlHQPR8b/Seoh6KGkK
TrwT+qJBlEj/6DSgyFCZwvcAsUKXcRhINQqBd4chB2UldsAgA9JyPR1a2yLk/5pQ
jHBmkcB0vmbKoTDSQlCnwspC4xnJjLMQuWSDf/YlVKckdSPlOrD6pxGPad4vfC4S
C38n420tEd1kMAUlyD04JQx0/ZR7dkp18Em+ILiue+9wlOh170H6z5rYMTjzntY9
F5eHm19WeyKuiWBXjDmNIVk+fHoVn2N4JJZgvBih2RdGpq7MLptfK4IBn3b9cDot
BS2QL9whFyrfIEVQ+GtZR34s3+gFKphMuRf1PiUQneVKlZizQb4Pt/fu2PKNLBie
/VuotLzBF8Q/vkFiwuPqExJhYUorFlD9ZOJM43fX46yBwPzudFZHR5eLlbUnayFz
e+EfRQ+/2mw+pyK7mvd9UlV/n7fOZeUrzNtJnjr3lz89Es3U6XkIPtsauoP5O9qH
uWImXs+oJnLXP16/XqFb/2WC/t3Ft2ZcCDiIPtB+wmhsnz7VUwjVaAYK1EM45clE
oB1kwVxQA8cbMwGO0Rfs7qS2cpnURM+lRefMz6Ox5Pqmu0u9xYjFczipy3ndnpwE
47XQLuq/F2Froo42FtHuFk/1ZxTa0m1Frb6x3ikIO11IEXi7CPbeP3fVPcZUZfFW
me3ne7eY8f+Bsy2rKxtPJn82qOzr1Kx+OmEeNwZeV812p+KIdehyPHFL8NxU8Odl
NPYf8qa6goUVPNM6XJQQcffNpeIYkTSx5rshSuNkAG8Ltyxhu15HUZDQJpk6+UQM
VNefcbs5Hh7i4/1LTM3yhRauDI+Hn3J/TNUQKn6W6zrzvbWrcw3d3pqZRp2U/Ll7
RF4RcwIdXxSyLzf/aYUqdACX9/sFtTTEnzIbTqWyDwI75E2+m5/1vFA9lCYrjq7D
Jp1GZarPry+g+b0PJ5KdqJ/qX7fWjmzyNYKeFF/zE5+H8GBqW2HCKGp9jRticHjU
72z/c+pIaNRCv7iUeN9D1sIsHBChCADeNDFr8+OBavWH1i9Z5dfvjHHUMPxKElnp
r7Y9I8mnrCKRGVsGkMUx/ufD3xRATPuxnitcZ/aP1l6hiPOyE53jtMTKLK1AZJGo
2uV0fJLlgUunucBuVLMm9U4De6YRcZcpKazZ6speK3pVWJgh/6bzp8bRrrYNS7ZY
iDq/bRiWGvrF4WY5Rt7s64+EFcgIo7MsAfxgp9E4A1yfINr77gOD2RlM5341/tS7
jiGFDngCJ37wVD1QQnKyl3jLT1IcrN9KeD6xVhW2cMR8LIutiBBZW5OOzOrMLYy3
hosxTKKdMcn6QcOYLWCSnHYZl9Kixz/m7jTTBdBNzeWt/npeaqmqiQrbItmxZXav
Xs+7iTy6WyoL9prVamJiMr9++MCNah26Flfotx+5CIGyll71MhsmixAULyiLwSFh
21jORaYOF+q65EjgQ46GWjLTvFVY1y+IxfAdXPwZAC/5LSf6cAd/sOs0aUCj6tVT
c4oC3TOJOZmMBlq6GVYrF6j4ry/L2suV3Q1GPcpFGHrLKFTdNgSR0AGUpneCyC6S
+8gFDCOxG0apLFu4RxywIq0MX30JQGCtNUziR5G+bDk5lsgv9H02NHFw27qr3BGU
m+jCT7PK8CsGGiJ6LYtW7vyMNT1Ws/K0UQDDlGwyS6ne/Cc3EucySf9cWS/cDhu4
a54f2feooiIXA5sMjBKj0Q5PhVEKPXR2x5udm4Mb5J8wdMQYeFP1rk2OPCuNEdyb
4VI47Uagggom0EamAV+yvSBXWK7wFQttBB8Y+GHsUCLYoE0wQ0KGUc0L5SwWBPJi
3N9ScbYqM9Ryqqx9klBVeRxQYpA6vm+3qyEaakMV6Y/TRtTprzuM8OrvhMsYb3hD
T31Mk/bWSaxNh+0v5ttuXAtGto9HGRzXDSAGekkQZQcXhFC84IXSqVxG/2VzA0bL
v4YI1TbcgpYER0YoqVpaPwVMO7Ni8NlYKbxqKN39rkvFr4MBxfakKB1qkXOBA/Xq
HG8cedM4BlBe5Pakbgcm8VBWEnFY5vHCU4C2N2pK3qJJtDd3AIeTcF1tg3H7krwh
PSJ3K+30NAQ4xVKkx4NWM2yoYxcjXbZpL8jaXDeuN4Bj3j3cv5Z7Y3kDJyI7q5Nk
QBwCrw/BuH1hYVrPrEWp3Db2Sxh0hgbcLVaILT8QDUI5v64ZPKElOZG2D02Qa4Wp
40+FSKuO8MSvh6Ki2oP903aTJjNjlj3T3uEuxxAnWQTOcdwzyD9Mybj5azd9x9m4
nnaDnUcHiTwObEoDsXwBybmaJrrvNSRTSLi/3JUYKMLR+ZypnYNcqS1HLSlr+TAx
Lf3Fx0LSICQDVM8pQeQWhzmBxoOVJginVe1RAK40//SfeVYiekGBkdn7oZ5ZA4H5
S3mIDg2MDOKNHQcl4Zk1KJtMGM2lOFvEYBufLZ943eS/XHJENjch/a1cYCFc5a6i
Qf2RaUoVNcC5qUSSuqn+7Q3ehdBEf/xJeNmyb/UDemowq7bgiu8qXrjlBXHhDXes
N2aH8s2yi0uaiyA6Ih++TsLcAlveDUg64WI9+5yOpAkaVsU7dwaX70U6KnEa7lcg
4lwnZbQu9op0K5+fzpUR+HOiCapYMfXoFqao0Doruw9Obu+Fs+iiyK7ETCGVkhdp
tpDYtoHWCvx0knN0ItZirvZoycu2TWBSzmfvBvo3TbpB+h3KhhzVI4b1IyCUNQV0
/KQC3D7qq8UXXuwv2yvR8a8Y6pUccJLegdGCr6CGRYUDwC59zww5xgy6vGryg0Mx
1sFCgfgsDvGiZzLT9RD+8xH1yuLLrpRDWvY1NDUkKakQtMdybqPBrdQSBecGs6Nc
qmY5VlpHUAkQO94GBtJUhIvzzOHGM64R9EUyZrqBCI20FTV0vue/BLMFuxQqmlyi
Z9v0FXVCiWtWoC42DO3GUwFFDDWd9piqpmopYKUbsnu5i9xAcEIlr943WCru0Tq7
cjHRgQ/gljJzD8GKJXBRMn3tH/7q80MHX8qrlAw3k+Nre5BMMrIUAmvTRImyI5zJ
6JGtxYkfLZDRvpbGdlVGty2oCFQVOuRevfKZuztLSyfFyd4A+zc7pWS7s8sq7dZo
tuTZR2JvNSdis+79u59Q+tsC1ALib2BprfktuZQPTYwVmrZmNKHKtzvc9MCN5BCH
b7IKKq6bqR8u5VSOMh4EAEeYgfc187W0YIK8+YXOBHua+/vc1f14ywr2nEoy+089
jp0EtB4fjoL51Mpalshci8XbPI0rLaYWS9JdrqGw4rrfSQ4m5s3xaH5R31b08h0h
ViEzMntNGp7/pi47yYUeZmFDNypw+QUKkq0ZaSeGIGjp2HqMLZ1ppTSJoSU+AxUl
LNqxj8wD6s455hP+JAGBJ8Cu7ZRqQFkQIe+8HBZpN9n828uGNEiwy38oyfUSu6gV
gNm4OiqBIJPn1svxQYIVe8Tj7s5oTNleBMz2YyZxKoU1aAiZHtyO4Rr/J73M9t8l
HIuvUwfzAgXAE5mpvoya0jSzSnTP8zr8cKw2tFUEKmf04R6SwHSJeOBLv5s+Yjbc
uG51cIzk00LaW7BqmkIo3Sah8N+5IalGbKKEEXPeC4n5oLw3tqRj4S9XrTjJSGeF
2Lyy2MsB3ERcGJ/P8+R7byYSErn0hxnNRTpRjWcfRSfM4Ftk6MBxhbbzSoMnmEcQ
WoZdyeHxxYlVt26vw//uRpGmnYFoKnvYwmLT3tTLaUbtUlvEhWz+FblxDllDHUVf
tSRZG3815mF4zUb3J6lI6UEFVruKRxPoz+nIJqT/62n3rM8P1pzbmFLmuJTidgLW
BYR5eO/Id3AM+iBw2Vq6UdFA5iO1pvHOE6Aw9+8kyrk6GxVXjbbIT0HbCAJyqVV1
rHFjJKyS6ULpYfx8sXIwlKJSo/wphM5EKnhlC2QhQpoP73ZXxtp9ww3wKhbodTsQ
8R1e0h4xochmyfDG8azIDPYRWOs690sBX/qTGeaTFQRfRVY2NlHRjMYLaNb4EfSI
JOwQ2J80oyj5sLDVkH/oYpqRlP0l+ZSs/zPRoWYEeVLJqMvimopOoXFWIUCnDVuR
qtKa3Sx6l4b60xNjPBjDCcclZ36AC+gYAVeUeRikUyX119WFzb5XuXUtJgxz+tQB
ddV3L0iAk/hsruzjEI0SGBfPnnj0nMm+c8+gUx/dLoCrKwGDeYP6sR6Oqy8xrODj
3uzvdxxykWlXgvEUHy+FIiQdVtnmDo4auhsVE1FlHbGX0qpu2wX4wte6Qv4rVEI+
zLY2zaBZ9JB5eVZtXhdjElwPR08/1ROQFeaRz8HPX8Hlb/MwLckZmWUSkFQ2+Za9
Ga2Nxfa/40cMsU70nr/6CuQVPGpS++ktNg8IMFXy++XVtLWphRFPmpYS/0QDZTZ1
7HyA3yYe8k+rZuyw5mUJYjYyqDXvaJOF8cKvC3gEvFYX2Dah89EU1DJR43jCHznO
EEJPDGQ+WXCVGf5owxqWycpVPpeSNbFZUfGrjf+7OGqvcvXAfvIsU0m8AZYWPFjU
5qt2BcjP5DFvSAA8fftdppsNhg5j0dB0b6unHFUwvsAu4zoo07qHaCNb52qyKOl6
IGR6oWZ2wSCwp2CWzJ/N2DXFG+/uC4hvjjKycgk+/QqgpFBacwdrgsA7Xl78hzwq
94nUewJA9VS7jXDt6ao+savI4ID6z02kEfa46+Bl1C2QXR9t3lpthPy4VC1Ym6Gq
oiVKYXCm20k7UFNQfcqJ9c3wPgFIl3LtDybWOY8XRFk1i1Tu1FzipXHQOMhNc3se
ukyfVjJ/y1o6tMVCHQkzX36pzQ1jRd8zMfUhtc8CHKrV6oKvAks6Criu58Z9ngH5
funsRksrNsnPUerVv6GQ+lvxeQxWOXc2b4QRSHnhEmWuNFY53NjNZ8eFwlQCxESd
R0pEjxk38JTn2taz+NdWPP7DVbiQZT3hHY6B9WHFKYhiD4eWNmFUG9vYsUgKZie8
FLtnC2sznebzGd2AnztJ/B3DhTKSa/Xpz6fNDwSFyIsEHkbcdMMxYxVrEM7tt+Me
TyIN062d+CyKOpTF/CUsWrcmtvKTr2CrHWXsA65Gw1a9sNHgGXE4XCdhi/daqiZc
voICI8GKQi8f8LHF5lszRCpJLFM+sJklBvsVXHSauFNGaAaDUsTmLWu4iXTFDZ+c
9ETKAB7Z+nmLhH32zBgFaldBR4/lC907ziU4yiaESPerZysU5hoENdKo9JZ6dHq+
lOvyAJbmxJC108hcv310nUagItHc5LI3feXvn5dL/KJLVaXIPuaIdxJgfP1DEDWm
dduNsi3JSdBPSZHEPyluKikN/B3SwDDz/Y8Wqv7YyJwtZ1y1DtqLUCfR4ym3HEvt
3rbWpFwmy3VBWhzFaif0VDakYueFPlRGZ2DiK+3EMjPYJA1dmKyjvoTWiYaoJwtu
MiMSI1CiHD86Dhfhf1m+ZdFngrhxm3iDjPJeIzsal+87jiVtwJif8n5S5xmCOI/r
2MXgNl942+uXiQKZnNAe4xc2axPzunf+4LtC3ahVVTqojyy9halQ6WcpTJXY8INK
6rCvL9xYwIgcICLfkvE1xHuoJK/FGhJ71O9b7MLheo3ug3y9tbqO98fQOoVftRKw
bW7oglrsDb1f/4H+lF9ay9WzuHXwT4CcDNLNZFEZwTNljsEMjzhomddQjkbYppaM
7B20yqSkKqQllqmfoDoFZjf/4oJ7pMN5DdCUTrFI5uqtjbdPGcEpTqej/DlAgbXa
oYL8IPVd+Pts32ilVIzIvHn30UlvHT8ImC8fIRScSNFZU3Bhsh5Uv+kdhr1FTh7I
+c0eK32KpjHVX+MN0CKwHI6xedyoeOKBMLY5W+BsT4bGMs3j0g+dy9H1XC2Bhrmq
fjibL+0VJfBiS2oBvh+HTMN9KVKwU8UWtj1hx4nj+AaZA/Wia0Ew9q7dR69DEjxe
vt0nwONrovP6FDXoVdw+gIHtJlWNqYTt+OW0AYxoZfxWFucWY0RsAS5+6ioAZODv
oRaAb7p/JRoXFqrvfV1wPe+tBozTBQnr2at3f5uQEIUI4htMFkr3pu1YPLheC1QJ
alA9plxmFDDOzFo7eIaVUpxWhspuXMAN0MsP+sQpPnxPIVjNdhiNFYpzXruuxVN9
W3cGiFNlwwkNwL34ImB4NEQQEpCpyXzhPPNc9E9HLc0CMIKhWFazGhTordHcDk2F
ocT1VkZx7xsLH1ZDVFpfkv0xsZFl6kcp+PE4bleAzVEObBBeV80+B9CWKWuVwiJX
dYVVn34aF7K3wRHpASY9QB9P9AdGNxG8T6gkktH49jFEdva6PjkdAGggW9tAeiEJ
nb1svySXdUJFFsrmlI+9CzDwgSqAgCawduECEF/jcFn71iOcuOprZNprViqhFZ51
4JSNk3+MJFHOIy53t/SjxDDpoRJ+u8EuHviBGfuTMu4+NR/9ZJWPxkPi8nm3PwLK
PCOVuhLo1++2YnyllIyWdyoCFxH0+Ml3uM9tXkpMoiw/6a+t7t4XNBDP1ok1LclX
mdnoeVhpoR4pOOcZZF72DPNJALRNmkEzAjUmW+PUjw3eHREnWFIkSnIU3VjhznuN
wyrrVgLGMHZEroW3YDGA9PUwhAnOsaarxVMX4Yg9yH3U0L32hnuOoXErwNKr7Gaj
LAJt6KIZKx4uDY6MA3cfI5D8lV3A3cc9znSNcywGdlfSciBlV0VCXeIQQBmcNOMx
pzRgz22bRMdBFUqTuflOZnbN2b8E1rMWhqeMm5hz8PmjJVxmuLl9cuTmx0DRynRI
0HNriACGjKQODGuiUJZb64INZVkydVC5oyEA4skWdsvH5EkA5mylUSmR6w/Zgd6C
5zn1SxIpet02WqrJAceqXLq6jz8gQUgK6TCEVAVRQUIEqJN12bgeQp/jlqTCeSO5
ym/2RYehuoOHTQdTkrbROAoyAHLQetwbhzimS3ymBVnRtC+fPCUah7FYOkFaLr1j
Yl8qLFv7OTbs6QQA7h0bvB+SXf/RvgVA80H7YjTDsg7jddjoCo4JTU/vdrlADzx7
VDdHQacDheczfOglKwYA58MFKmFuDOZoGC8rW3qA5vqu16p2qb/o6aLAjqCH+fjX
ooTr/yZqxjlgPHWaIcTOmCXKrGwaEQ0z0aa8jdI5nmNmsXYJpnrsrpQ6RNYfbXHQ
rMCJ3xFHLB7OhBoh6yb7gXBs7DdZF0cTHLKoLziMSgHzrxGcPZJsUepmUMmLs3xK
lUscTfMenxOecuSQD8vbirYeFEp9EIPxdxR2I6OUo1DR0WeUzYe39ffYrLG6DiHv
V3BqGY2nIegZd8bUla/U45bapLy54jMZE2lszbi/iuYH0+3wrI5FhURjHP3y2j0y
Y+az2KFjJHK9WduT5wu7Fe279o9jiDoqg8lWzm8D2OMprWuuLMKEa6CTgrBx1fIZ
6QXVYghGBHtb1XaMtnQVyAwr6nRY1wXa1WJ4ubx30eX2oRs6zovY3X8/Kf33FSlP
a2R8XmV+RWjJqmfJE2OUxrZwoj7kREFVw4U3jAbBh2Bq/aF/aInQUtVTUOJzv8Gk
YbSb6vldSwDNn6snMkkJZ9VJ+9sqJPL/ddBitIUt/ewhhHBn83oGvRKTKnIWz/Gz
Q8Nvejuy4NSe+UV3gD60IdsYajTymFc1CTTJiWC4/hf/lJtx3SPaWSdf5lpMzkOI
wHaQV2Pce4WQaaay7Fl3R7XeoapEhPXCWre1AHhPCACXItPf6IYB5bSf+Gy8er4t
fmKb7y56XqNz/g6I6rRjuM04VFTaY27MWLdcwKBsGD2sHzv/ytFZO7axLK/hrRNY
LolpX8EdlZmN3tpHeyVzFi0jsNc30zaF/89qvRhrUkSNGCisSRROl22yM8/he6M5
adsNRKAZwZpMW1Fypgto2k52roZyeovkc6wAbt6WC3KUIYuGax44hZGV3ZbwRv6R
eySIr6Y2iePrdcv7JiO1mj/IQBVY0w8BI+SP/w23/NwzaJWxaMxoVR+f82iglNrI
ZIvOMRMLJIEJhfSeD/52lnF04IzUHhnjmfxj3m2rEWODJgp32dRl6oSp7/lRS+qr
vVNaLCXTmzM5GtfhECHFPXMHfxQHDGWkJHX1iSetzGVX7gH3Q7kOtv4rjH1LRgQp
B1PQNFHwsp2o2Xx4FitlJL781dHvHSud81U3cUEXvXBnsGBgCY1BZjMJ6yvPPv0M
nJ6ah1waeIG3HK4ZUECkPx3TZJn4gMbTsnqV6S6XKspZS6ph2mGx91pEVztH120G
LvRTp9OI/O3K8RYLuCDoU69xcujChAq0aeBL2lPnrM4YvfZ2w7dACdEY4pEO8af5
IUuFpPOU0DZzulU8aHm/qZLfhZsJb+TnM5Cpp5maku0frU0Tci0ZLtWhojvvWSjx
bLCTFxEEyiv/j7NpY7YmgvZWPO18zBbvInebyb/E6l5PPpwfHctQ/nCf6iGmSMxv
8HMuHcwccLdDy4nuLVz6GtDBqWFUBQKAkKHrZfG88+fVHg8kDSFerGYgGV0MMmsj
NCtY+e4fc/fXGFTtDPFUYBdbBzIFeUgCiI7JU73HsmcrtVwDPpLkA4C4aEZAETmJ
r96J4eI5SaF88UwI4WI7t//FGJ/KhowraHfqZNovTtB4pvnKk7i8nDERj0Dm0tMq
Tn+Iqa3Wei9xkyx4nKjwjku070iy42gp/Ci3RD6S291u7UcSOFx3DASb4XZrzTyI
O3ab0jXzdvEr2BgUgHFG4H5HBP+52/3zrk0zXCixDdGEdex8TtKkYfMwYZeaZtk8
1RMvkK0C8ad61vBHUksi0+74Nt1wFVgYfsFkktatp7J5iJ2qdUCu7+pJLwYlUfNx
QzO2fM1bsRKyEHfLeP+AqgERZUxGHBy5UTaIAqZfHpDZFJC9Cvn1efVhhHlQJo6P
pqSJAtAJ4hsWy6lTwMXrxiDb7SokEB6A1Yt7FOIB0Dq+I1kkAB87vGzxUSCnleKe
KHLCZMA0IpHhq7q+LQ7LfznKM34TMvIizrv2garFt8V4WLzn3MeECm+6W/eHeOMf
1AQcPT+zfvifJuSnKupRNdpv6vgeUaCxfEvrJcFDAhj3XpZlOfzj/7X03OGMU0qA
yvmi91WeQDyUVQZfOyMMQcig96Ez3qoKOEB4c2g0GjX6c9V7PJXBRDUugu+JXfMn
oLRtjRmfbxwETqqvfmOuUFqSISsYHYtr9Ei+0qChv5uoahSlKwu6nTuz7Vth7rhQ
lZi25RIVqIZcpmI+MYL9anAjQjrz88LOd6+m3lZBDfLdDJIhJ6CcqqVO8zcDpvfJ
woCq43JSvu+oV8AjtcN7iVRpHWqMeenhLG/CG4VkYxVn43yX700B+qEFSq9jHCXa
LAi61zgp267pSgcheyBmY9kKgzsCz5XKd9TQeehn+ZABHIPNualqMp4Z57eKosBD
rICukO52i3u2hnAvdWN+F7fCCOxH5nx1TCgd3Qhwv7+AP12NlvwenA9xd4wy5nkC
FZEW5VcAtkeLCttZINVFfFjJs8o4J+a3PN/38PZ+W2AHVPVwxMtl1pknxaIJvVQA
8MsK18pmqTlExe8TPflUhQAZdYkAL/tI3MbAzgLUFxNBF26NO748ZQmjPBveGt+E
8R95hEZjNnaSGpAu2xTXu0pIaGD+0LxuuZYgqjMCxxS3mlF69yPq67I5NJ3BUnLj
DpvFnuP/ZvkQrCUy8S0ir8ZJxeqPj7Sq0evXR/xdWe0BzArfoy1Wn1rN69ksCjY8
C1vCH+shMagiEu3qS11+cYU9brMViUmCN7BVOpTA9tVsO9GlPeDm0F++5bi7P8Et
8lrfJV7oLfFjzMGvoetoz0WeWj2ArFqpdE7bKBW8tv4Bl+AcwSl5pQD7C0C4JNPF
FF6Zv9nnBQRrEPkEPCAWqICIHa7PmtQ2bc/z+s2CGtUAbbGMVzLiwkMg8RKVUMpv
snal4Ev+qOUSZw+UDi3K9ukwHtvQQOKYcLJ+P7DH9IY9Rt8RwY1TAJGoAFZpnL1w
wuWozSqilQ/n9iVDheTMlF37nWIcqV8cbBaERaAqQhYsqV7PYuhH29S4WD8ILD5T
/zK7geppqSK6/SGBaxV14KBCLZUV64NMr24sWzvKwbuTbdrlYyHK9XLtrVdXg/59
hWMNMvCPT5qIOV8EtnXZit6sKDnDkkqMZ8wVcjmzB1Q/6psgmin94DJhfwO9AGQ/
tTnjHXjD4og4c0Rhv0m0fpNVq7wkBg3t0iQgz6Re5xTQHWWY1Cvvcz1UlQ6MiGzb
H/IuGrBUylmnHJ6rhu+KYwU71fMyWn4PVxGwM/h9XBook6GAKZ1D+oJFq7KoXSOQ
AzYObwGPhbasqXRKj82HXcm86og27mqxMlyKXiu8LKD+EIJMHD3XgIRDec/EsKVN
9z9SvMP6FZMgu9gHxp7vTKfGnBHj5U3p3bZ6LnGrd2QGaoOmPzSShRK0klj/sW8o
9DZEK4t9naw6QhR8hvPZIKEEql/9L4oY49BFuIdaUcbLs5CyCV3g6nOG6DyTThEV
BfDsfzFDOt5BArvRsn7q8DZFnoUTCKlrdglpug8nZpCEAoACuBiZGNalGhrF8F5U
qn+u0Ghq0fsjxexITI4sFMrf6o7bFYANwoeYMBuVQSoV72YdJCe/0pZunEj0NlqR
WHuwWXkDkYw/774qsSXy4XfffVzyP0zSMDiYdlAst+4un9kCPd8KUCdcxYL4HY/6
gByWZxvjAn1pWxfCd7m9tumuJYSG/kJwqoaoD9ljhV1SE50mijfjDlnLZ3ILttpd
WB9nwoINnXfByFH8/z4UPx6iJ8/ejGjT/vC70tFExzLKKjIMgs8PZCI5mSk5V7jx
IoHbFoGv2bOonaGb1Mo+EqvI00+CGbL6ExJ8pUzt1NLYd+7dPjszsMyGPmnUoT9+
tMEhIWvGnp9Mfn10o3TeBU3/kIaTB4gnn3tEfr4TXE4+3vW7g733sZrbANLDHRnn
gingOIwiKlnbQjL7tj3QybajoHRfTPoCUZnaSjLc2OmcO1YNZ11X+hMzk1iCxK7A
dek1CI9IJdSjIJq5b7RGwgmRndo1pLih08Cjw90wIvcW+YzUozIIkVTAFR6Ktsrf
CkMFNwT3FDyHVcKqqn5FjUkN9JP69i2H7uHP0G8ZzVnAtEHdU+RJh9imtR+ByTjw
bv0Rh3ZgVE/cvwvOliMPup+3c3/6pJgUd89Y0Gw6gZLPtGMDr8X8mDxMQqMhCTe7
8CcQ9ABsA1a08weToqjkzr6mdPya286jxeRRxcGvIhy5/qq1WziYVFFFjKV4C9I4
L58+kSZPmbs8mnXFd9WamUTSYSdw6TQ86YXfXrq1kxTCD7GzMT861MSxJ2iAA9Zj
aW49ulm4tDns5G93K0Rfw0DQXvMo/dASHhC8i9GKEnBRr3dRHU0/ncELElvO/QBg
6nS+fdpykKROMBiKAqk4X6OfB5yCXMjEiV3uYh7xsfLDirtgPMmC5PLo34ksvgbl
jXGK+T2SuVXeKKv6lhAlcZt2dvYNXgV6WNGtw3599sWwmG4xDIi2GJMdc6Tcnj6G
YC+CFBs8J/HF98vjrXsp/jWyGqCmpvSYljzxszxLjL/ejYr7einIrUKucoErX9Ei
bKMTBGp4rOlBfuDFv32Wvm4uoqpIC4b2mbGebtjdqEn/ntsBYK+15gYd8RdcNquK
ssz5pIy3PAXFa4SmP7q8iiogmq4KGcII7qTDQ9gzURw1UeJsO79TuwgUyam8TJGQ
WBg/Sj0CZdG3Lv7sn68xrnBZg3OE+Vg5B7QR3B2u0jval4h/0KsYRLVeTKCoDNOu
Wc85SGWPxJP5UOx69axNvd/cTtGdVW6BIgdyfy+qYEclurdwomdZxUaBbfuhCXnE
BnHZmeKG4IzCLwLjtiIFq2JrU9plx0Adm7QBZUwB0gKo7W7qAHhzulq4n1HQQu4r
UnGbO4CNXcYnhIabmluaWBQzsUNb/Drlq2F08+qLDLeRuOmSnV7oVhQwxRYKnwSH
w1YczNTgGakM4ShgmxW7SfEmTU43KLKfnyPPQWJmTJCt1WAJy0LIkis1ofTskHzB
gA8Z11f+IiiYmaDV+34Nqk2WfTZNrOCFZPynTffzOA0/RBM+fP9r9PqAEjKgqWVC
8ImSaR5JCdg3gCv2zOjxTw7JSF/Zi/WY0h6Fa6b0Y3UcMbuxOdzTsHcuBW+Z6oS+
dR3Q6FDgyY+wufI9NdnnqauZW94L+QJUJIEbrKCxMV0iRJOAuuq7AvKE58j3ONcJ
Q0GNZmxPOSebOUXcc9psDF0uR2VhanCnKSxdndHA0n8CCQyt1ROcGvFp2WOCwGIk
BTKvqpToW3fT4LU4MpR+oqoTVJc1B9JGgTr5BShLeCZMfCLZZdiCL2y2UNcPiUXu
acxGH2xfcLWY8lxupnO27SDVMdB5C+8UN2sgU2iifmZ9L9sB3B65G4/xLDdcMbk2
m0SySd3uxsS1g3gDcnU5M5lIEKU//38dvcC0+rIkxQbl4pngr31uN0crZwKXNROb
ZNkKbiFZodT/bAPjlEMRNbmgcPu9igzwJzx0nfisMA9sOpprkEz9LAJOMDv1OY62
435loIeh5nwzVkUfGHdldJDwJ8MvXqAiofdx/Ux1+Ez/vO8lChkxkRZdagfy6EFB
8S5R71xImWMHgGFNK7KYpQObyz70bSOBMH4ZM+eNhWqng288B3Ume2SNBTx7bGpd
gCXMrZt+nFpWtTAaZIcsCVy6UDgh+ZmB0bmI1/3MFfaJZ3MiXCzIMVGHggVpFdh4
H9ieqzuC5YhWhf2w+kHeUVuSIQD3SCSpcTvYm018iH9fO5zxk6IHqNK50fVtPlVw
kmlIYAuUnH78YtgKw5AB690/j7+T22aroabozAGZR3xf3EB7WjLMG9E5mrr41C3D
pD8h/B6likbJvEhO5dtQMH7ZXyX+OfW3JUVwF8Y0lUka8l6v/Gzc2GTc43rNLwA/
GOWUvzOS5lvtb8CHtosaU/uLY8EVKOokMzWu6GfFAJKkZkANfcqrlNyf6T7JYLic
lmo6vtZnqL4MxPzywBPK6TehWtIX3qqmdU4G6rzUiFo+O18UsRoxHIivZVALPl5r
8tThoEVgcTrqE5AsvDzzuQaCwtfUKM5DsgdXSRiSjhpZsO1XWwDxwnoCP/ZXDxZa
7phvkt7IClkTv5jMCeh6F0jvRafeAaZL56KmdUpX23+mkIBwHJcFhirLH6OsJ5cm
peC2SHqqr/+PWRQ7GjBxcresiREik0zdYpNKUqsJzoh/bhRSDLBXKAihf+2/gIkF
MvZBPa6AC+nWjKf8Qs4+tQ04MAgmySTDVDy5931cHLvDVO6LCb/w6p4TC6puPw8E
4TJ5IhLFq7DNamjKMeVbHcKs1BKapzGKgPmcTrzZZYnsNQCw01VCqZ2uEyFPdNM4
XYDNqLqafiyNXOaQwr3gecPSX/nlt8AZqwiLzu564SX2vhCsGSKjB/A+f9oJ08BO
oO1zSK3VmGWV0RqFOBJpOuvedksZyYPtbyIvTd929ZtNZyncd4VdlTKIzWICKFIX
FLHC4OlYs4ScDAr+iVn//7BQyRRzgJXzhaRtKpPjcUcfL6ioDzMmWli1YkZk9GLi
5lIaw9V+pS0UBQZvNbHpdeQ2ozzxJ9wWBQ9Ck1Qz/2knAIunSSh/LUQJvNAOxN4N
r+BuJNlinF9cJPYzV1UWXu0pS8obtTV4hYoZa32z3cZ8cOGwIlnRV1cmxPmlOsZm
0PVGoF7afCHIW1dUqRrdQUD3R9OYkI5ptcqdWlMbus51vUaeX7BXXYP9GJ+0eRZ7
/p6KvfLhxDmqXFwy47gO4o4uoAyvYIa7A3KznDyIO52aZNXA6sulFKrk6XV7KLSl
O5JZEnSyIxb3fP00XX7DTD/HMLAujmf5N7tf8kWOxlX2+gZsZDviiWm+V6eBwQWD
+qHbgw998R4wwnOMW03Q0sRDJ8pmg4Z+XF3+2VGRWxCIJC2Zsjxbdf71z/6VP4kj
lSyxaRdZgNgZ0mU1DbznW4IcKO4f5N3sI1C8k1SW17grtj/eRFv9pSPJNyPKkkZs
NzyPx2FKsU/ZIbxXcsEiGXn6sEfMWo0es6brb9GPqEfIIfUAtO2gPgHu146h/fSX
k6UywlO0w5nytapC6HhYLz1WuSEnmVCWHHDG1Pg4Fj7wn/teWggAztigeKrh60Os
LpBM5tZCKbe9a+C/hJzLUiMrFTJe8ELrfOoTdRSrKOFkL3lW5sy7rlmx0SLI+fkt
g+CYHEPdXvnRD7sQ0YoX5iZ+Ba6a9plxe35OzMQF/yjabOi7XUTZDxTsyQtTxda1
517xzddQ4TpKRHNjT7InGUVp09R8N2wBOrN5RYh1xK5QNs3Ji8ZuMaxV1MIBMv0Q
xmPF4BrKsspQrHd0neeEsBQtcQ+I+K+NkLXu0o7+MSvk7WTbiU14kIW7qpsCKwos
hTiIkL1Hx6SPTDD4C08zYLTXDTaw7pNinAHpRunHOkih+ZsmJ1n4TQKex7w9X9Pn
xff1A5bacsJs9WLAWpVl3gHxJfEE4bld6rJ4uJcwZho8qVqrpODvgk9quzTkSgWZ
R67ElLbE8lv9uFnI+yiPqKe1iiASnXq/O6cQ4DUr9DoATPq6xd4B5ifDPRM6eCW3
xIdk5sFUfcN0NBOBHFB1qHqmT2su6OnoeoUQ0bZDiddTeBdPkrAatXqiwJ6fhJVN
Jrvj4jBzSifh+7skc5GlnkCEsuXY/JomM9Lg8fEqxNwsHKu+UOYDKQOjnh0s8bMU
DrlCvuV59c2HdnNJf0I3X1lgpAVRv/J3kH7uCEaYLy2XtgoUYd4CcsE7GtqQb7Gb
a9XG6fOxS0PSpzEXQsZ/8qTbgeCpGog4ONPIOILad/8zV9HiJ6dcGLKeQDCG62lK
hvLaqBmXjMwvya+bgwWEdvm0aowU0fXLR9UQekaW86IPzpI8NrHIgwFXW5jHYiJC
QAclb1xc3kc8kEtppYjgA0ytPnb25hW1w60VDUnaCLjjphQcG+epcKlx9K1mhHaR
J8Bz1KDqTfsXGrl5IrPKlSW38AUzl48hpoqUsOAt10Ckrsb3oE7dn7215PEsCRmN
T2LwvxzhAtMkb6yL/veh0qlsSPqxeLR2PBZRZOl0haVQBQgNAVxiu2zoMTeIDxDt
D/Twua2LZGYR6B+sFRCRgba91o0kqodtNveOhgcQaA/y8kjk1Ik0cIME5pi/qInq
Fk3sOCw6h2agtfRDvaLq9X5Q6/sXI2S+xsDE3VmuEFsTxKxxXB79/9ib6+/7Vc/f
QebLwUyTGWSwwP95BiO/Nf2q0YYmMjR4cx2P8+kMFSDV/ZIKssZtTCHa2uS6jFV6
9vvsmZfBJ7WM5BCdMyejtiAQzJ/aPzxrHclJH4o1RbMN27oBVKz5sPjB4KrjOC5G
mzHJ1dg5Vs356I4j47X/zv72xgW5din4Eao+oQwXErnxjoqpSWtCE+/Bz1v5p7GS
cwqB2+W98kL2DOKvu1fIsi84CghSLYHdvwDT0Kwp3i8wV97yIFJmV6MVhlbz2ybC
MBGz2MeCjYVgciXu0hcZ8fhsQp5Was9p1mkeI9pdEBRpJlQclVw0EiJs9FAWiWPY
K52B+B6mTQQPu3/U+5gJaAudQKM5c1hM+9A6im/GqcCIo5ducU/Bc7iCbxZ6TaQ3
wWjTdAyu4CXzn+SJekRDoF/fNYYwV6ahd9URT3htC0BP95zWupItijyx/8EaoULV
bLP5vmB5bKbQDgQQCTiNeiCVdp5NC/DURorPSDcAr8xuz2u4ZvdQsSh4fNjfyEx0
rZK0b4Avs6X4EDOYmUw6gCh2T4Qu2awumre2d/9EIurP5t6Gv423ceZrfY2rrEoM
GlBn33LAuYMXH6YhW+87a7zZ3I4Z5p5gi9CJKVN2UF98Am0FLZyIFcY7z8SSC/Lq
lwWhglYe66oMMijkMopoiQQzDUqLINgbMDtOjObEt7/rYDteI3pkKud8AArfYWDh
Ryk24NnFWFjl6Gj1YO6AEyQb24B5Iw7q8Vy+eRh+GI2DUVdPL/Qm1dV0S0DVvAje
gUJuHp4ALEcAPNibIz7Okd8wJNPsgR77fBAr/7qICh1wNQ4DIRCCwcJyBo8ZFg9Q
UR+omuOQ1QnjpBc/SVUoh2TMuFm+nBfNz/i+AiKoAUgwYKcH7Z1WAiaefLtQNwEb
Bif3eb2sZsS/MhXu7UW+7C+NFaslbEzc6x5oZqj8tTN6qo0Oh9oajSHzsqtqVKVo
8+XSoCccThcpQMjJv440xqFPrR/vCNgqVA06+Bl4DOTtuZ1DA+5VRKf2qR3DfXmK
sOymvrn4KyRzcplohkqT1MF9y9dfHuiZHFg642Z6YiSDcsq5D/6g6LfGn3fX43WB
jgSoPYcXpoFfuTeRQ0+b2ZvsMlA+EOOvvbCqcNeZpC4aX3GLoK+tuSzyTBJUmMbr
3406yLiPH3hWKqjaMYc5emugv2oJPWYn7sB562u67kiD4Z6JyuIutq7p817xUpr7
HHYlW2AKkU7qq3QVx1m3Ccd5oN13KZ0BaRwAkB/5T/hSGrf8l++W2fVOIlTP8DVe
7VKtGubtIl66HyG4gr4NLsiS45k9mRj1FTv6qrtFhE1htazeonqsxmkT1OTKNYYt
7aKqbRCYwPFHpKi/9+L1JGcF0q9wT61rFN0JCdOXgdKul5184Glus0WatLpPX0FX
sFy9ijXALOs1ooIoOip7NOf29U0ZfoNtAqREF3oLoKe+H7l0EXSB3TFPTbJM5Rgl
IHguR4+A4JKGSPzJ0819n8DH99NS5g/R7OsPsUv+Oz2wQEa0xaasRihfTNeI6rd8
tPhAJYWfaaf2SWKSco9QPLqdwKYsC53+p30WN+7E2jmavfqy0VrbErz+wl0W8flK
pT21DCsBSeywdODExhBW0hKPPF6BuANjnyKQEsIzUsjNm143Nhp5AdtAJ50mebH0
JXU0ksvqVO1rEZeZMwzMHjETKeWVatzJo55JfOKHNVk9OlXfw/nQ6/mffxVLmRvJ
IchYK7U79SqDHz/Lf8DCQ1CHvdK0Uo7DKHNyQeQVxQH43NbayLa7uh/Xnex4xNhX
zc+QLY3kHDtFZQPxD+SB79jaBOedBmkx7h8Z5M1kSRV1BLpiqPH5r49dhSS8BAXc
6GdyoMIEQCzxGI0/BtnlWMxt0ep3HnJjac0gqUvgGORr2f3dB2l92ExdeIUrKFxN
ZP3LBdC8RReOakcbMxDWSlJqzdtMojdvsc364MIT/OqSx2mq+x4AQIBGuLHCNUQY
ve9yXpiyGoUKwdmJzRimudK7ELtiupZ2Yg/9rlzzOmEot3RjzR9x+aTKi2AbyurD
yCrb+/J0m3qHj7yY9wfNChtyobtez03usiUFlBvJwLAr/rRHHY1sgrOYEZf1zdIr
P0rl4TKfLIT9zTRzrW9IIyALMwTuXB6OAL3SEgdubVq6NcqQ6KMcq6cyVSUUaaGT
fJ1dK1qBFUtIUK0HAouOad1Cy3sJ8kVDt/npBm+4VHe0N+UmGkYcINJYcuTvjVnm
DM/Rd6YASY3x4ujl80p1fW7X6vfBzboRR37rQt87j0+qih/6s17c2ON6DaYECD57
94d7IgKXPrSgCbeHSHiCe35/j6RyKDpMY7F1ZscCs1BHya5XhWZuVM1xBxxUfAvK
00LPzj604wfp7+YLLYSUOkV3Wa7GYCoXVmWltJh6h6y8juTWGkmbr3bGwhCJYkeo
n7ebDa4tybs+FJUQy06JgHzTdtZ2rkwykBLVIVM2hWW7xNGQPD7Egcwq0mD9LZtU
gpXeoFf7+oUUz1DfsUSeO2iI7YSDbT5dIvj1AaMbVJzvhIaeJWCx+GGiY1ZWdXLu
n4XXqj2F72p23J4S4uVTG+4eYSQvMwa/0ezcT87+TjuB1HSWJRaoKbE+Xk/m2sXn
dK/XbAlB9Ie90igOIDKo1kSoKqpNJC9dB0w6/ObeWa8f1qBUEqaE0KTn7DNByfeT
PVGWZHNnUcNgVIsCyjTXDDe6v62syxWQiSggtCmHbEy2z2FCcjPe6ZIYUnN9NCww
HG3KEWDV6iakXJENEoo3S/XG6beo70XUbw02+6SGX8FMdamXOQ5CYvyPvsmOyyvS
6rdjhTdrVA4nAcZMqqpTYJMrvs8dlMcZDxpXK5KN9wSRSr7WxNBRMNLyfA3Zu0Yy
aW/zAy42Q6Mm8v+/ET7jdRrRS73AP78o2JqB4RsuztdueYhakqBeoSos3SRFeDzl
87ZqJFAL2EIOOsinQWpJvdaUOO4EPxeASxyh1KKJJchyXVO52XD41kQliF9zjb6A
sxydCr7+2CdNMw1OMeTtLCRYlDzu+UUkT8v5ewPAs75Lzs45e3w54MYW0ojwTkV5
LWEWkJUxbfz+u6IlczrCu7WRzmkR2fDZUyb8Ty93ffKMKhaawrvVxps0y832P/G3
jkQ8YFmWwsClA8LuxyWgIeA+PBhrHfmqajDOKbneXAf7fJOh8KwMpw6NzbkjCFZ7
i187xEOGaxAvU3bqgd1MUx1fyMUHcqOW19U1Z8lIjJ4eDCGDaIHMQL9MmtL9SVpP
Nx/99keUYsL3W+G48No30wNEhWrqwL+3Y43CfVMDzlhNDO0jxydWLJdCDjyrq2T8
r4nahYxu4ibIyc5tZKP07KaBmrV4diN0Z67W2jKZWGInKMWIuwfOO+BGfOapI1rA
5mig/kA7/W5Slo94gP4bS8RaTs9pa+qGEpH4jzSkUtYStzqABZBaSBnn1YtQVxaN
ZEs9+cFhsBW8CSY83p+fl5nzzNUmlTGna3RMEKXBp+GJ7uun/lYH7cTfHsbaorrQ
pQRGuHgHFZTntA8htwp62lQCw+adtnZE+W08QonS6VGvI55r5rkoZyxtw6DsLe5f
j6q6THrCbTmN7OxzSzQ7UmsmUHnOgpzDe4aW29Q7C9v3dK9/H1jQJzNO4HQXfYf8
gBRrMwSScKhDP+qsVcoqpj6OOfNI/njE7m1FA5ivevqEvCr3Qrm9VaSNy7x3S5ql
Ylebi9/0TrByyARDlGv+jURWfP59r5gNxIWKUjdn7Iy1JfI7xqsyaH44+645vBek
bqE01vqDID5JLzXeNMadB9tmQ/DGIhrxsB4QF9E7h2+SWrJivqiUBz783yivIkyq
8z3w6uc/tKgq5aq4xf1rZ0XuxSItLcKlFucFqkGcrQnOzESUKRgMYiyhmHPvt15U
KD/X1PuMJH3sviRfyVIyNbZ9ATE0vTSLY4moYXrEU/OQDPOvCHkFhB8kEaOMGTLu
ro/hudOWoMm1EWm1+eOZ5icgR7DUHXgSxPOjWBbUjkm9YppQaRyimPqSEGoR+3BX
sbDEoBDAoIzg+DzW2rgkDz9ozgyvNjWXNgnFSvyTPBgaMfsfumnQD5YnSy47bjeU
RGnkVweEn0wl5rzJ7LeYCYc8oAeETcvkngOZ0goMx8Z1Jp+ThXSPmgIlbjZI7hhE
AxyAY4lJLlHb3x62If8LXkt2qAiDrwWQSqeInPqY+6z9m8cXBzUHw17x7axl/zJD
aPSNn2t6ezlmhhENFoQMUPQOMzuoxo190bjaXmvVXNA9TeqFsB3F2TxjiFGLNyeO
dMcRndXVIea9gE9JyDPeg5Z2kvXhbDTbCnzkc6G3SMwdZm6Nrateykw/MC0M+UjO
A2AvxOXEhaZwjxeGCYxdZ61JzoY6pl6X8SBjP9sbDmsHuCswZPnywzQe6oU8YtD1
nV76CYDQH7rZPO9xqCwLKWZm1AnF+NvRWA/PUC3w5PNRlax0SA4sEp1BlD8jizDR
ag1a5r65qJAg1Tie8axJ3RO8RjHMu8hWviqOhbac3nZOrYH7/GxHNxwWu1iz6s7C
Syt2nHu6PZ0V+KtosnPpJNA8v6nVNAAlejzqd6ajqJoMK0Yo0wfiS+JYHP7VGAcQ
bkLq4b35tOf458pa+HPChCOG/L0a6cex07WCe+6T/n9VF6+xWWpKzRafc8TC2qYZ
xuwNn6bIQXdyVm4g1QUV0sMa4ADOmQke0AcWrAo2qvQeIRpRQ/QHaHBTyc2igYeo
BU8MPA9ZpaD8/zP70TYi6XJHGt+A9imatX8LERj4+YGuj8D/6xbge4Q6j6ckZ+T1
AcUJk9I9vcy4c3Q/gOVedYd/liCd0tkB0005uBeEcOV1DLWidYq0xzd7+ahzaja/
xdS5GdOJRlVSPYAK+TJV+CAeZgVMNHKUvb4RHc0HeCliQvW64HOQBj7k8U7yS9HL
jbd68enkfYfhQ20fuwub4XuhvKE+81j2U6nBZpwCuq3DjlWPRFi071W2D9Yr+sA5
yG5rGT3Pv99L8ojsf0/+zwBNlmvyWPy04h/JZtUi90GzpL2bPH+ErJQxGIIxA4v1
7mE47ThobCwNeS/G1as8bal1Ijs1+FtSMa9fGME0NOD3y74MkxJ702QMN/Ol6jGe
jVTtuRnhp1BQ9qCqbqk/zSR3JTZzEPZJsnSCm1WqjSFXN9ph3zcOCHJQwqNpdvBz
Qkgfb6y7bTSwrMWA/xKZAmvonvkdVuTOXm5CGAvePMZzMd0+qISIonXwd4mHz7T4
DmPE/jY2ftW/a2uJrLhdNlnHWIO6t/ibaJ/J2n8EjRCglxLwY9YyZxw0tMQspZim
KOdLNfoOC4pbzOKzLYxqS0mH1WJ0yyANCF45GZcVOKKzXtB55yH2h2hJ30B8VWgZ
1poXBfoO/0ngXubG5HvmeMtNPpLa72RF9AGQc6dAs7KWtxBuRzJh2xWb282ze4xa
124Kfsb6JY0KWlKbRI1H9MQw3xmSBnpVzpZjKzdnAZIafY2buqAobJQGIwqA2kbc
y3TvoN9Ol71JlTwU55EcRbLt0kqZw/8+P+17cNccpyKKmO9NEpy+4e/wiz6jxI4F
vdhZZwJaGKspf4yxkkDDNs6C2UY/tb77Y/lRnHl4OLYh/p0hiSFoyIRXBXxF39gA
KMVDNpRZTwLOAmRxx8dB/ctmH0k8lbP88mP3/2lo0xoCdVJaGqz+yuDBGREHGUyV
x1ufFYXXPoHDmk/yyTIiOab3yAuaqzEqj+9bznVY3ZEZcGprZGxImi5KddcIDhQK
0A4LxrIzmiSyfqpsrCwjHHur5AY4udhd81ZQWJYuiHWEtLwRmfVbbQ+lk370iOf8
BFXZ5KEkjcBmMT+He1DLGYTz6tSYhiC8WaIlh1D14iAhFYQYrqkCpm80eWMfSzsK
WtA9NMZel0lb8x5fqSJeeNMQVS4i5QhOwA/Icy0JEnj6Y1Fsz+5uCv3D8AK0TOfr
1I40rpUsyRIotoebBxtPomF9YjOWhqUk8Yli3wGZzTrw5pNZLIPWiY30Qx6Nrh+1
i6sqUwhEavrNxPJobbvAaAFW4XMTeUmE3wWUZFIPJm4Gnsu+NfLi9WOxZLpwiNsF
ksKeJtVWpg0NvA83LyR1foKWYIBo0Skyi9B4DY7wq/eTako6a2JlVXVAALqJvWNV
fSNlQgodwHQcYILKzJEaUv4HPJkB6/C1zPPSrgqM+1W9J/mFt17tnE0sYoiHYBLq
piV/izuaeLGAIfPcMDtm013FPkme1tTRhHiDFVc05vo0Bn7DyMjsMRnQJji15Dex
ruhqET/pTcoJpJcS9XfrNZR7M9C6HcZxj/unxlkaOaPMM/gFpCG4ot+SvU509J4g
KCU9jMXbJnW7SbO2JVh7XDEie/qmbsWfQn8OZ7cxCTmWRQO0W+L2gs4T3qV2C7Yd
tBXUuOZoxo0HuF5NqR2bTaGWXkuCILb2CAeMYmatLg0kIwN6c/o497GDAGTZTpiq
3vBzBnGWSIsMeyZx7bl4W0BWiYoRSJ8fL1nDWyj/BHRh0aWi7LelwW0ZFWqNWmjL
hEOVpQoDVhbLkgZl6zTnr2MZTb2sZ2OVgjpb1ZnM5LQhhVutm4cZ3vzrVENUkVYt
kSNQaXLceh/ne1lE8z4ZtXVSuKntGqjGuUqcZTGcOfy75HTQnklgTsOpuHnMO9ru
aHAg2ZcsPota8c/z/DEv/84S00XuNijqDyQqxxvw+Tg0kAfotJSJYLfRMcWrj6tG
QvS4VSjo/swd90Lm9wR6m4jApcpEfKAxbAHOlF8/5vWWYp53ojkyHCZtW81oVhnl
sadvlz7P7V5n2Ot6aiEt7B5rVtRY/+7dRafTk7uP+Rbx2obj5zpNDdpVW9eUfK24
0FHWoiRhTEWZ7IFCwaajdg9gV7pqZKFuQvmiC/uA7Bnwa1QdtI3x86LKDlWoWPTq
4XYVagMI5djjZedZuPJKt60oKp1nVd/up4BjiI7OlLnEz8g35Ixh20XJgRvCApjY
3OLh+Egx+wABW8XtlBgs9hLl6wHwAWsY+A9/25dLCmRAU8uyVzayulCKvdvs7/oN
yuH2+8iFLtDs8hIzLHYcLoT+gW41JyoamhJzufE4zhdm3P9jS1fuuBlRwAkU4084
n9gP7PLJqtit2e3hKNPri3ZI97sYW2lqWSelwNZ6mn1zvEPl466C/mY1CbMnPkL6
Zg5BmsrVwSXsR4quNdesQsFrFKbCRm1AJOU5JxkagXZkiQoZW5CH8Y/9ZwvWiiyU
271BrPMSf2nWvULM3dDG0xg4MHOrLBxWXBcu06r3IyxvMQ5H1WrLAQtgRo3o5s3G
yV87fJEAMwSLkboC0d3zfo3DJ+93QIaX7p+XavKLxgS1T8DboQlNP86ehvn50J/Q
qc/hhkgsjHkzowYXS4VwtLWgXb4rFufc1BGE7/Om4BPhKEcYy+qLb7lj2xNcgiWJ
TkPihiKXFZEelcvygQzOH3x87oDuXHGdug6IWReDpjjPlMMsOlJl9/Soh39YNSpO
Pvul/I3bqDsVPH3C19JVF/HESDZ/b/4aBh608y7WyjzdGrgvn2L+wPkFkN5ssqIj
9gV0GEcTip2gZJa5kkUXudcepwzUvJWyPbZOTqOhznzSDtyovr43g6AjwwWYJ957
8v75Vr3iMipnK/pM/F+JiH0X1wAotBZZJzLWScFpLC7nbYP2Ld440kZxUZ/8VEcy
lCj8MS9dULUAb5lWmLeuDg0sFbUndokgrhVGxxa/E/svYeVXc4FvopTsWCZCVNfv
dfu3+u6cavVSuBqX22rRH9RkRaBAr6R/upuPwjE0DQwWVYFpurxHKa3p49zhhrg6
2E1AGsJWI87PQ88UiAtRwjcBRiGY9Rg9ptvD8nfXRmwEDo6hM24d+jb8jEKXfVi+
HBPiJ2i3u8jyuFESpXv+tV+B9sC9VnWOSJ/UlV6VS2XPlAXz8Xajsrr0c/IfOkrr
wSBr2DvK2tF1OTAstQF1ndQ7PioOgTx7jirFFBXX5Rm3zKyiF4lpnTDaLyF6BSy9
8DYuhbSukIQv2QovnJ/rZuxPNbomR39RpqK9tb9f0FcWHR1Qn+cJWhXxfVPAzFMM
2aTLa0J9iCxOgE2IOLAtupbjAMyoB3OC0C9dzrEPr/U4njW0A1rpPVZf47ayDBLE
wz6Hsrcmhs4tSvZwJyu5LX8H8fAIN4BJfHU/CXOgiNaK1rY+h2gRfF3BLW3bcJAk
cEO8CyruypFrOc9PHk+BfQZFzDzykADxygU0jQbGZ/CE3K6YEUsYr8QvRbqhl5Lj
FXii47mIqeWU33oiVe6FqFeHSQfXmbVy2YDRq+vspsBIpAE6tsxfJECbwYQnCW+P
vLgeBjqXHFHWKsxqvZ1th/ZHb6/BIky++4I9yslAVXpK3qsFTtxSkiy5GM1/013b
T3gaq+BxPMwv/G6K9a3V8htrc+iRnV0/WtDN/xJfJcD26SNlyS8RGJUmbke9XoPx
OhGNcz1TgTvlK7XxIVFCixPk/BmQgz8WLKppeZox8/G9sUOmtDe8Bk7xCN6HSjHz
ib15iewdkUOPd3h3cEK4qeX38j+yJ4nSo1fimnqLOwlidNMFDTMXivPBaBZLYHNP
4clzKoqV6c6Y3iKwn2ZKhdZ828AOvUANgQmxpffBf4L/lsOJuqjxyVIOtXxingLx
X8fvqPWN8PvMMw/Y7idm3UeVk5jLnQxOP+rPS/r1VCG3FLF3i1MrHkGmfT00Wyo6
WIaz44OV4meYHyR7iweyjc0UyoUF20+kOjlnOtfFWXlDQdHpHa2Hdnkiw53wE5ED
DZ9ASd1wsMOCzOsBuShksw92ag4SAuzFBkeHvcaCSWbCkoW3UT2h7CIIk6QCtdKB
7+G9L5gqk40j4+VzJMMUtFmuFu8SnqEVVWnwiJzzKe+oYCZHmwg4OYYy7raLLaLn
6sbeM+A3r7EgfJtiP4Et0UmdmBY18JzMLy/5asX76cPMyMFneyzjCCBaNqCoyRAN
F5ZripiqQVNhtvS8GKmw+IqruhrddWJnxYfjMm7wM6Dsm5nW8zZqjzvKnVTmTxqW
Skg2KwUoUPVrv4uW9DRwP8GlF0KLN4MvAnjF3wOliVQi+QALe5eaLRKRYtNh3Wku
+Hmr3o6Z+jJb3+S1G3riYZPsPm7DX0TlDlKAU+2U6IrDzgYp/v0LFm8jv4e7Dmpz
WsmcC26y92fay0kRViYhK9R+dLWjzig0IeDuo3SnwVgHg3N8iaAMnG4X+cmT5/Fv
pVMciGDi3NJc90DC+4f5b6mrI5ncejeBU7vpPhsVJKFdM3l5ELd4Vd2JDZak5OuI
IinCUqlyEtg5f5lH4CK1y9jJqs/l9y7WI2K9l8LYzdgvn0P4QkO3VY5fjhk4oS0Z
4vlVM0mlKVyM0bH5yyNq6YRJfWe5g4gNDycZLtxUD3wpAcPOMv0kYItZwNnnsE1w
sW6wx81utN6GIjQKWUrusjqHVtBRjvTeP/HR3Yt18mP1K9qWolrYc9fb7LUbDCXu
ztHBpbh9coZ0HTF9RYFxlzNvbeW/GCrvFH0bIKSJ+c7RQtyCRXpLMboUlX92eVbo
0dvYT3DW+KbnjRAMm7LaS4Tui8JKzX02AjlGJFz6ySH24nCr0PGpnEvBgX13eUUM
zlxY9oP65TXmr2SKdRWJXtHsovFGoijb87+pPfUAhFWZHmmOTsRZvVbzzrg1+dkS
gLlNAPPbwo45yCSg6CEn5RLkH5JD5YlOmSwpaowUBWRsezWyaO54UuNWI7xOoln2
ldCGycFexK2zZ0iI7BLmMSZxCynCYg4ntQZ/SU1JJksDJRuSMo2JTGBQ7BrxZpd3
h1AvnfOXmEVLWaOaKqySfuWY4g5olUbbgLtkiy13s+dXeugM7GMwxtPgw/U7f2rw
IUGL1ro46nkVS8e5QrBMbzl5FkB6dUbXOp6Uic3nbvaBdWsr8E8267OySjrWmrBm
GcW+JVqdbE2nKV1Vi2eCO5eQjnNleIMb/ln7idIqQSWVk4Ff+KMD2sOGn8OC3KzI
DCmepKriVHSPT6eHUAmTPk9KFjhXMgzXPHyJIxyzfQaRQksxvAYKnoBv82g318NK
GQnv/jh6htgj3y4Ii2JJ4MKbKvejfLhmBqzWBEPsfzErt0ADwpDW3Kw+HNC9EZSq
S17szz1ccYG2GJ6aWuTFRdmhRBIfcwDbzHSSnpBxZCVSnW8pZziJparPeJjkhc/B
oc9uwfGstqjJaRrONA6YS+raPoYAISoRC40uyRNwg3wBA5zLRoJSK9W4mbwK5uK5
1DKxcs+y6o4wf3AKwnWjbaOKx9OVgOGyXafalzS+fEd4gmfywlvm92M5Cjg+xgwa
4RqHd9sEJ+EPJsG6TL+ZcBofF6FtDa+7rQ6pkzCuay32yCnvbjabSmxbRrFnQgAa
lY4FPHxZj69jJRP4n6PxRASR9PgNIGoopBjtuN1ZqcR9IY3rmitV32wXmisaa4Zu
MywBhFKD3AuJwYy9xTfAWDBHFYDc0eel7l0v5OFX0FoXyvnBd7gJ6pHh5CeWOWxT
9B/Ta6eVD4NGosy/brAezLbHF1pOMRR4QSyVaZbGMBNfeuCcoFDjaJ/dhtXRaOxb
2NhzdLvBWGAICgApOsI5KdwyRkpn3gr9NhAC1n6E8udaJijg9+SY4vPt3oiUq6kf
IfJRC5QvhzGPk5D6el9JQESQG53mcOxokivz3ttX+/W65er7akKEPCEUiYoofkyT
fnkXtdiJYyrz9moQcz08KJngrIouLIeZ9u3V1glw0GBie9ssrpnc+3gXREBJiLWE
kE/X4itqHhEd9HQeWwcyNfSsuD/wOsisCZGH/6kyLID3+HOYT+Q9sMQVBtEH+dZx
i47XyjAI8PqTBcPyTyEdLjeeoC4Ap/k96upkg9NmjW2Z8T0emLZUOHind0H0Fj5R
4tA8Fi49mkrXUUIZKZMV+9+TFw4WYkRAsjVA63Fz9vJV5ydLrXYPv7hJ8ALzGk7U
Q8VaKs1It+sgUiRiqdF4oKWBCKCAL0Bnr8j0vI1+Uv3hbGt4qt2kSdsINj5ZV8ff
bhd9PSb9WH+YRtakC+M5LbL4aimQgd9zER2fjfWrhVvNyFuocpBGrgivrLuuLdSg
fczSFhGKh5AAiAQFD05fg7S6RHhwiq1oFHFCEa4uqva+MfH9S8uZIl1+LaSzAl9r
NC3Rc4nSmePYSawSQpb846pRZxXMW6x35XI9XlO/FRXXQIfDVE4496ch9++CTrdc
Ur+rtKIxkDUPKGooT4l7FH1zKivSu4zHf1WxO7QLK8zfVQmcQHGayGj2Tgp6RBYg
+x2HIlDZeIp1Z4+Vy74RFymVX/AM0ox2sA53OAd37h1n1WcAMtJIphcCGKJfZbhE
X82JCEasEogxLnOYiQupmQMrlwa522avGTCXm1dgCx5hQx8ekMTiB+PbVhE7vndM
DzCWDkSCc/dsIRvfdSFLymwsmIw3ZA07HV2tQeNfXghVcHj5LNiJLdF2t6sHt9/X
V18uT/qBFtyGJpGKOi0cqRa/kMQK5uAGors3u10yMjlSxDmBJMniIn4a5Kxks/mM
g6RMUyteXvkvSLNn0x2DRFrL049abAFJx3mWiYhKHVEooERLDWfRpDyIw5KYQ36W
+5EPJ0StBR3nCCRMoA2X4ZzUOlkuE2v7xngyBJX0yru5anYzz1JTeOkBLhM3XZsx
UPwkzj/fc/NAHBKwumaVmy66qGlflKdjF060IDYanUYzhg5hSPx1VIce58EK05XB
SxF/mlHjStZKc7jwYIhhosY9+W5bnsEUdwjYstKk4qqReV28BDe2WpnEQiUS7XFK
/kV0GG9n21MIe0znimRSvytQ6s2jH/JPNoFeOvdzW17BqaqdXo1I1vgtChvYZqxT
BWuft8TsyMdYYnl03t3t9MozCV36Ew75Rr6nTAfI8iLO2MljDOA8Cfpbf8bW6axO
qUaYI/PIBlwUQMZFqXAiRny/dljlyEinhhbbCYod3SsvSmmnQFaNCmQq8geQnnI8
3alFP5IbevJuF5C2tMco7fwcVjcuMRfboUA9mkG4dih4YN0FEQQTtvNEbuywmtHI
8GnEWQHlPsjxLl68wln0uMv+CRq8YHq1qprv+ch4s8Kp67coYNKFzbiWfLWXv2F5
hC8EzvMSSVUSOsFa+mqiWIu3569sJ0mjtm9EC0Q/l1Rk7vRHhaCahbriZNAgwYa/
D4cmulqfZa5RViGcJaURFxZee6CzmJXJ9eyKsdaU6novtNIFdqC5pAeTBAbFqI/J
WIcQGnARGWgr8DmCHvRIB/w1M52S/tcWmYt52Z8k53wnzUIWa4UV0arQ0B0cbylw
LuMGyoRZtfSm5K1YkBNYICiDZDBLMLRSHRltzYvS4qFDdqm9RUx/gnUY1An81wRh
3gmmgawOA3GTf7cizpPB8hQ3sZyUIhZFB2NAEo++mxfeyyAhQuOY4MHqTfyxhMJd
1prTZxtNJs9F6QOg6VgdOEtdwGLOMOM9VZFplXzFsalS4sUUGsaBvOMxYuntx0v8
rC03gmRJCh+T/yPzn/6VVDh8KsVUurn5spOX58YhUhHnbHHdMP/S2W6fm91Hb2d1
DeIFlqi/6+j1618SRfqMpqNwVZffTa3UuHlRBiJ4aaXp5cIuxJRJ17lcNQ9k2dKJ
PMuL02wBwAoxfYwGCERfnm3sWqQm1Jhcu7LILXbzOsFoc1piVpaR6xtmEbTXh5S/
q31fG5Rmnp0F3+r2ev9sG9kF9wJTen+juRukuNXuzTHjh9oAfmMcpP4EpqrZA4DW
pA0F6ZArCIej6I/lkriCn2eIoJiYB2jqvzzfm3NlZdy4IslBafVpxO00qRTVi3qu
TgsN1IBzJh0u/+lz7FT4NPr9pUEc3Zb5mz4hf99bO57X7iGllWwEEW4iNbWL8dcE
swRs1O2/aHsLmrl+eUF3wG38E89wQzHAyFQuLPTChXUL+jUs1aF1yIb2LIy8Nduj
a+dnyK2QuDmPGaGQpvVc7QrOxMaNf9kfsnp731rqyZsWPKIY2dglB6u7Ax7aazmJ
zx6rJ9/Jyrv43xVABktD3kuThSRbXuMxKWeEJfGtp1pWdl7rqVoWLmKjKj/rvmN2
UYc9MqPf2lV9R5z1hNVhaARTSWCF0nm1f2ncNBAmZz2jIcfnxkVc27PzGuKjoqfX
S3+qK6U8gysc5GhwvkvKPn27wHacoC/ez7q4zvx3o4tyPUFb+qdUX21lpg2Cpkvm
daEALus8vnOqe/FKxp1VIpkx3wMXn5HLZnOp25hm37A19OTXxWyxWDDs018cIq+z
S3YNO0KcUxvlrzkfrWc/Bo5BAX1+WPvffc99Ua7ixVzUCRSDplSiEJBF9ar40ac7
xzxII+of7z4VcJeGo2KxRV2SuWdnxB80w4LM6cAmUsnBk/U0mpT5KyRP/HaDbM/M
DieySEt2uin3ClNCdDgL3VXabPCEeetiLi/vgkmcJu7+moDXmOEVXKeGlupwR6W1
Iid7FQm71UYViHWGgAgHDHWhR8mEbaKhk9YqvEcfIyH+IpO1315psmwkMvBdAB+4
2CvniX+BZ0rJc8KXRixC2aOeiUU1+0DIHgu4eK5pIuzBlNs2LlRPws0pZTgXSdJ+
6blPnOfQj89SURy7jjHBDX+l7VbELtmYnZH592BysKrqitOpVFCP4BrvYiFqY3vk
htRNk1vVzZWPIT6zv7mscumClbv0VAw1qtPe1jWsP4l1nkhjGI4TGyNFUrv/0OKD
VECtsQD/3c+cSCbHsu9D1RG6YJUSsQSoClW5DPWUjsXShTIS3LPf8OocPxQBr9VN
acbopCphGol/pKmbH3kqA0gYwoA41rrwr18yAJTYfU/7coeSpXMange4I6BjqfLN
f9Wt9uo5i6Z9s0ktbfW5lIKeuBkEX1yNcUM9M4qr3Afzr6MBxLfw3J9Lu02svdBx
fEXvuA8EKv4+giAVFtnlbu7bLZcih7NLOctzDRo3o1fDG1i5GfE2wOGg6+BHMT1C
pOv535RsajeHpfsv2V1fudVY5OSABDwZQbCGe77JnCbqE5m09auWdfzeExzz/Q1/
MvZBtbqcjbgAmKvc6IzZ65dBM0aP03CkyOEgS7HiOSFCT9O4pEaOef/1+wj3bxca
K5OBG0SIss6V8GR575s+CBRfzJ1FkzUES+Bw4Rr5QpTwS20KaO8bIgfOwz2WRd9B
IrPMQI38p+BuBqLfaLqGFP8Gt3K1lHMQiDnCoob73odxQPyiPzj2vuuPAEkKPQZA
VFodugr3cMO5VJENOZmhMvJF/+zb9SsIBssMT9Br3owJhw5BFnRyH2WtE0L0v8SF
pMk9xInJBA1rrxr/LwTCF+lyjARP8jeQ6n8Oq6LTZ2CmlyZ0gt1v1PIfFkS/4z6g
wvb4pAcmUiDGb9AmFVxl3BZBWH/EOF0amcvG+x7N15vZn+SKBcut4t6/+aTYyIj7
+K4103MZpI1O0lG2cB+pCh4sNat8YZK5s2qD1apQcjd6InNLy0p1ME/w9JZ2G5B/
ubv1RcUSB0Zuk3lAz9YOwJtK/i1k8stAwvP0vJ9siuYiXx3cjcqA7DZ0/Fr+9dKw
bnTUrKJ8stYpJ/o+bDx9/sBe/v5YwV4+Vj0EhNL6KjSjK9tuQP7MLhfPDUZN/bPz
T5b6A8ZYMgekNSxdALOjm1sn4j1RTeNBYGFV37hd6p9LX7jSF7hrHXi8jTll2nID
HSKjlcmcIKulT2s9Jn87DlIyXZFWJAMFgJyfnINJ5+K2UMvnucdwuhlS3ShIVYCq
fEKYs+0lzC5RGiOAQ90c35ZseaSvauDjJxeCndXn5GKcQZ3Mq+51QOmU2lrCs+9H
2i3lxWoRxfp2GFZrxIuFpHwv66MrN2JawmCDt2tvPLRBUQLbZC7OhBQIDFhGw0q4
fvH/RSms2lt6JFYYtm7+uJTWLmuOFmfWdQekgA/cqTRKBN2toV21t7xnbvDeXu4O
Hma2nCrnwKVyzOj+bM/uLWpUqoZd2/4qf4CDZY2xfRSEsAVqaMYEQQelhnyqDQq6
cr+136YM8JgG7/rCJjD1rXlAako1Sx1OsH1NiBiuUOR/aa/2uiEXWUDh5q71BKM6
jstDuucDXIEFm3qMgZxsGgyDELkEIj68TXPLudabEy38FzptByo1p8Kx4LwdCUBb
fwToFnNcSgRlwQlNS0MTPpTDL59oGLIw5vGEPbbW9sNb2JEKqDmWvAKD0CrhmOoi
q3kCQG3zz+f9OLiiZDBmEfH6SjT83sYn6NSFU04uH5iZ3KJ1uUcNPhwWuOjyvsyR
sYhZ2CevUy5ywVV/FqzU6L+D6iTT7O7fcbKywir7o5JL4DLD8T6vAZIRfjQ7O7wb
+147cANyPt2FM1VF8jpDPIotIOaoWzhqPIxKIVzuzQhS5Yh5njXnih5oQWSZzhBq
cVDfc9yixDxXrdM4Cy5v6QPfGyghsj4oS3yDYDFDSGEMBkWzOm8fW4Q5jZZZLk7p
iWXJQwyFn6jjHUpp4Q8dcDxl3ZwyYr8dC11QePtBrT/wMuQRJTPp2kiB1M9RNJ0S
SlvBrCgO0Mw8M1RyoIHdoUOhvfml5/7//e0piG/etaRCLRqtAR8FSAMenF/iio9K
mVUxsl5FT1bET2GgTMmo/mCpImDlx4LKd5uvYIQVD7grV48kBh+R6KJq3vaC43Xk
2b1gZHGKWXjRim1lVXrvim/OegSCBV+jhrvoCbty5LjVAnbBToW9M10JR11Sw3m1
Cf6oNv3O8DmQkC66qOLWc8PYVBOduupgMnMEA5NeaJiTZmZW0B9qXbjj0SaMwrSP
qNV/CWOYtG7zqG1aERtCqwxqE8EbDyyLjr3Ssriujkhu3lcch3/mI/fNFwhyb142
LxJuHPPq8jTBds5+UdL+QVtnP4q1tYRiRZbU2dLFKwvtyDYJvIOy7T8AtejP69E9
2joVtz3ZVB9NoE6xHuI0YQkeY0TfKh311M/QiDKnCH8l9dELq88hsdaaD21WH81i
61N95x5t38hpg5SXPKXZaUjH7QOzYtWpnpkRPx80GRA3fiqkdN2dY5cD7ZGawWvd
69Y4P4OCDgeCNWJhqkFoiTBFv98/qyKuJeT2Ek0Kk61DTG4i4kdVKiq9GsYVfPX2
tgwzaFc787J5RTgY1W8ymMSPa90M/x3/+d8xAp5kIbp3tbOS/mY5+JbIvmSkwumS
Huf4ubLf5P24oMR2zfBSVPmMjG9zo7gzMRM8y4Yzou3AXojR1EMENLzgrmivC3ap
X7wX29jKEHmZU8rObgXAfJ3azDjcSBWYO7tFWmtbk1829T75eY8dTqkKBg7UGHpW
oXLH39vBZwdKeNoviTWf+qnUfTK80O2FNSCC7Yddffqg6fV/S39xgXdtqzBe00c/
q6Y7Mj1ZdtV8aKqawopl9a/TBJZ56+a3O1GxwF8cfwKuENvELYjXwlElhknZRlcK
lmrxI6ghx/VmYsWZnpOjxmNzYbyxbQLcCVS8y/iIheN2R1Hjmv5nGZWxiZ6eKRPf
64r5ImlAVqoqR7twAiAGc5BCX3TRYSaIWERHUZ1bYAQeq7Rq4cAop32Ur/3vEvnr
zym0yUWQ1S0NZjrMsGLvcr69+zLpZVfPmjSCRqHyaTs/MRbqxK0H5hqhXrUrwYvv
RRAgeBUcVl0FxW8rt3riwbrwjdkdQmqONak5ettsYF+chjed6NVkDPGBYlmc55OX
BGg8d2V6k5BAwG2lYCzfZqR4h7DFcVKORn0cC82HFyO9/C/JAMFles9QncOURe7K
eEOss1CuxXW4VQV6yFTpPqtveLon23muqiHNNfT/9Gg9FRrocTLdKgsw5SUmydS1
rCBME8cNPfj4t1D6ll8nMRCPkb4SZLEWfafsjPn7I1hl2WKJcXULtTk8w+pmlXtr
aHxlgmWoGHZYGoKFWzN82g92deAz7Xmt1zH2jJ6d05bunGSQ/qhUz360LYrFSPcx
H3L3D8Y9KpocdqKZjttQvxSYo8E6CCSDgR9gRKk8NWo6mPRx07NTjtclirhM5V98
sEQIXom/hYclF8749sphe+fguMZsWEjGf4FQDPq1p+y5nuQIqw3jLElA5j5kmo3a
5v2C1A4dCaoDCpT/Un8VjdaxDZ3l1E79dud52Z2O1JXlY4/2qq/2GH58rxh3DBm1
I392bCuhqgVKeFreqGoQwU2RmFCwv7QWlcCMvg5wXdy4/AXGscBmtO1PIjzN+Ptx
4LREfrV6pXw2yfXXUO9ZGqHsvfakLKySQ3LNqdxx3E4iBbPhErV9wYC/PB8mC6sF
kYdtz+YyGBSwbemXpCrVwpZZKBDOSJmJA7nLy/kfZ6W31kQeOvspt7t12aKYIoBc
D06y5gn/+JzTPiMuVVKEHdWkJ5DmPIzJk7a4juU1sqCCEspz3nLZuWxM82wynkOK
Q7DEEus6m2oLMikDn/CFgyh/cR3vZsUBqC8CnRvjkE6VcPCHk9wQKsXdwdf3LHvU
YVivi3VxFAKbZge5ogjzxa8omHUn36DJeKU1dzinP2CQ/VAqQ8XPBvn6Xq3R0QU+
baN3HJUQtX4hc9y1t6qF1IWvgM4WZeDbvr6KMFUlAfXQdiA7N6JcMgG13ZFjW5Wz
fRbhelqFPxPjpuKMjCR+06rH7WRupMAxkgGVYvZ81nuDDoLIj63cyGf6lNnTwBgV
+IuQu3pTfQBjCaEJ77BBUBocC5UTclUokoEZcnUs/y4UUuAI1k22/Ht7t2woTEQh
r/m5qasmZpnoYcu/Dh45JKCfTZHhh+HDgLB05+0lEKCiR332MnIzLoMGcVfh/PFy
vimn5566Ad0sj4cQPLXeTgnPNaH1P0XY+E8c786WRXAfbx90dGIdmnlKB/T4SAYo
rAqp368MQxhZ3QW61pwNp0QcqvY+vUDLIvEkmQOaqexVBIy5RGCwGeKsxK3hH9/M
pHpqC/k72t269aGG99Bk4AfpdWqcxkXJc2rcUX1W4NG47wyqgTFvPyD9LCj7YR3o
/LtE9LsLJRMN6FJ5eJFz5zTG2F6N+anFFj8d60dyg6dzDzl6wjdqmqiBf2DOZ+ba
Zbkotf5txCWUJRjUTL/+cO4yAgrgo8Q0WH8vFh0tVjW9jTzDR/1HyojwlNaYG3rZ
jv2n2h90fx6UxIIAg6mt8e9TwOXyLfA2XlaESe3pzbax3Rb3RvGt2LUtnc64z/Q0
RYkMiuRRZvPmpwHjQKtJ8fJwHZ/p0R/ZDMR/Mih7ZPycujSD4H3DzHWJwXUVwEGM
QxTna49IkRPc8N4aFCXXbX8+RI+pNKMwX/ktaIG+zzkscK7eDFWr7F8ln0xCbDi+
nOtaBeTBoGbIGtGMHpuKJbDyYp/W4XK7CgKOiyg//DOL5Y7C3dQDj4HLQrUbQNt5
eyqyd+uojHcJEnpsQcCPBQa2u6Prl8/vjLJbcTLluKQRMizEHjgcMR2yzmvkU01Y
q6C0G9f1lE98stkZszaLIigK9Ty8g1lPJqZ9ogxXvDOb8sQdTavK6dlywsnQyJe/
nRR2cIWF5Jn7S4Jep6//O3OG7QN5gYWflQkOL2f6d5ypD/Its62xbJ1aPprjdsxg
ZimPkJjCmIDd/mOUF1kTKGdT0MdUHDL7u6wKf7hG502rOvfvrP3rPxRdKK2fHzKb
WDizaW8dLpB3+IyGQzBAt6vF921EsVERQB2UulENAr1glImuCQnfjnPtT0Ft8vnz
5l4VVy7eN/t+g7PWrBAzBdD01DLHXqlqgQJJqYslEbsVUcicLqjLh8kCQo9xbjE4
0ynECnWMjsLEsVqS5Fs32OVRpRsmsuWUspmh9ZyFJHjd5dKt/g4pG5OrQmbtjZLo
7yeuFSyHnnfa2z7M2+3cQV1f8/cL5xFO49XW2VN7ZjeOzPXlYBTe+zPUT0SUFt0r
bTRFoVH0nIstZx3kAQTjlPiOZfIh7EkkreQwGtIPvuI4en9hQtG9kmy05KE4voYy
p5WUbREaMiW7vARZhMgrcw9q84X7PKB0t1Od63/vIaeKfzD7/hLI1o5KqaXeBp/c
9uwbIbeMka2OBj9TN4q5VoGPmhWH479wOwGjhXWL7RGUq/0oyfXdobJGqLVS6L7b
SGgpZywlHbMUfHXTXGRCU5OhfuQs60U79BZNCwT+aXhFPNHYWW8k4e1XVTF/cxrn
VzJzpA3wwqSXed/kaiNjd1gTT0gPtQ53sl0kPvAX0fIv0H+AEsZJAItE+7sOmRsq
UP43+gSAMUhH2TNbs4kNye3/QKIAsZrSjWRfUBfAGNzaTPAbEfcr7oJ6bcrRnKgs
gm0KfIekqjnHfkMzDj8BsKDX29vez73Dz1QvmyfZPP/Mnjbo9k5sSHbHvQnilc7z
+xgkttAT2VAV48wviMJtms+APC2j67fN5/56v6aak6fVNWJmI2zZQRF75J/8Fjj7
jy/SDldiU35JfI5UHVuvygiF0L3CXOSjMHlhIc9DEr7YmKTa96JWe0B6JVTC0hRf
0oGje+/DGglgxl+nwn2+Tl4bSsyJov/0FQtVg91emQG4BM5MlPCtHTOZ1AJNt+XH
aExmnu0+PoeKeSUN0e7LSFSL9PlhuWj0ri8+qZDUWB4QtCuq8UfiTM7ePQSNDy/e
9rCTMLCVRo6AMUslAFJDWtHVFO3RKiEBPSzLV0EGPZ8fvU22/G91U5YwsHElGPjI
JlWR3BWPxEniW6hNSbwLwTdmVbGudD7uNXU9/4EGQUeJI4iR7FCzLFeRFwMmKLgz
ZUHSU4eKxYZVh4UqoxOdnmyjmUzM2kEcsEc/I4kekvnZK4v/bQBiHS4g8sbL7pHR
rMJ3GMWklJX5eG3i9Y6x8pKETSUTvrhrGxvb14Xa+ps+af7zm6tcUdcIQNNO5ia7
amR1QrNkq3TvDAkQJIn4LIOyLL+tc/u7ebel7BVsV8kxEXGx2zs9fiVsipzWv29M
GzdTCm9OX0qFkmy7oQUifi4x36KHmkjJYpcv7j6o6zRJ+sDsFBDiFmi79LCLM6uN
osyOZdBzG/lA5uFVk4oEPvTzSmc0B3V7r2+S9tmlpFNHR0nHe3S4zH7Idfwq8G8j
n5VmCBlWQUFVe2vuDPNt8VXVfG/LZbwnh2f6g5GLpnPBoMzyrW6R7sSSVZnKddOr
G6ER5kbx2w39e7nEnBIsgPmNou88EUaGDpSg3UetM+kF7IClUVRXKqM8TyXfG34a
v5piK5EHDKj17J5fYT9kF1cLvTn89dxoQxEkzx3LZS9YkTubuByLxxCfUKUVhozS
NR5T6UqOKIaBlLH63Bu2a9Gh/+zQR3a8Tu+9imVf/Ti3YkpOHfj9yO9vKjs3sOAv
f/nTryqZKkRdXo4mgS/L5ZXxxOBk1H3oIhNBupNkjWNU+7LoDY3uL87UTQ9pBft8
rCKzMZUb97S0mM2tG85TK68fvFK2Uw3ZNHrrcXazUDqlLO1AJxUQ6uJNNq55zkSu
QCwaRwnWfrfmAYYXBbHiVFTunwWtfFNi1NqNRr5UN+ocGHKNkuFJebkqqNe50R02
u3y3BUJcE7boX2ct39UspJDFd3FeYf5SyLt8RNkWgz2OKCtP4zPa/AwuGYtGv7Sg
IYb6quG+3Egva2gktPBP2txV5cj7ah50S6SaTbRi1QgORWZB+lmpkwVm0TB8oNCw
vhPIbkDxRgK7pXFN19TpjDUgDnA/UqYekvgwdsmbTLtAe9DCI0woMIQEPC7bOfRr
HEGshXH3LxE4MGFDNZGtB6u0n4JP/uWEUba/V1WWvzMXbNv+/grkev+b/jQeoLe8
bAHrQuOVJIvm1jOE+fEY1OC5kkPHWkjvbPHdu9/ausZ/UOzLQLwvHP5Nu9i+yZgb
Mdt/pHQCE0Bzn7Komb+k55nrvKh8DdREhaHe0LV4Wlbe3FrVTOAIdTjTzCv0T2qC
z+2F0JPzUWIIW2he7kiUWDNkGO0t++7DwGyVGzJOQBE1Xyl4/xNR6GRLHoKisbDg
dlS/FQpQ+msAcIZNu9tZaJAUPUJJErahV7BUOr3WCicnKn/tabnhoUKvMr35SVEK
b98Fsg0VmEcqizu1cOu/vS0Lq9ZKK51mYLzXIoNX1M9jDzbwNQYP8H05KvyKeObk
fQ/0CllI7ZdepiGrd9yzKHpZBpkES/3zPacTZ8pG+ZHG5QdYjGb0lXbeU/lgae6C
gVLh/Ngm4MaVOglvp4i/Uj2Nc83A0Dn7ji4EJ7vkjk+ZVivhFXDyLFuqnVFuqzq+
tmhH20CAd+uQWnyQfuXUisD9Z+tdZrLxDY9dxHHoJIOXhMseeB4bFg7m32ZA7WJE
8uJilvWGrNoNyKkXssLQk9ZmGZxUCEUfK2E3Jp2lcRKkrlrkVXe2yAZQuLI13IM1
9Vl7/8h97MW9qGirwrlrGSP/52AYuPZbVJ76OjPloOqSDsTlUb7Q6mhoXZZHFl1b
YerOVEtsmvbzd6nrqoNk/yrzQamgIx0i/SyT8XYmrXsgA8QYKE63uBARJ7TcdZrP
tuxsK10fN4tpqBZH1nttzj2J7aFJ+NIzPHCFQ3hNUXsK/vnq1p4RpSOMvhBxl3Tr
LnQKyDLegrOTX0ZgO3OzGN7Vp9oVJSeTNp+v9xkcVizBPinoLpqcmGcirFxbrtXO
Nl12g9pKeUQYLwTMu0+SUkzTydEG4xDm4vATItRRPaV5nN19oR6x60LX2/WYuHdE
PLXXag8KGo2vDSXG56ryBqm+7+pYvC787nd/9S4O0gB1OO4LTvya/rZ0AL+Ey9wK
hjzOW1IiQZKjGEV929Jq898HTDBDefF5qEyHHQg5pjNoapDi7VvYVARYzqEqiiFO
OA6c7C9lxIP3nYZUZrxLeTNKumNVBkbcGjdGozTJNkrQzvOvjJh9BHY0PgGgl4uo
UgB1M0Zp/Ww0OyVigdquGEDiHhGWagdXsGYy4sQWyZd1S/LB96AjgGQF5XCtja/Z
XcQyPcHeoJwXEXsIVqdXiUesJnS+q2tU3eUYHXtxaXXqJojtvLebvq9cLxWy922x
8f22Oshc+x4GL//ziIzPoorEXq0KrvBf1HoJI8artJhKs4Mz0vFGtarN8+kgaT3N
GZL3mQbZpXjwL97+y8hBz5E8LC1B/05PqA8GLTKPpOHVjK8BtnI92HD0Nu1e/V3Z
k7gCMtTNlrn//VrEavM2suCuTooFSrfdWEDcm9+8VZgfMS0IDCMvJE8MMebaRfn5
EGajWfhmncfZ1wgTeeD+DQJyu/7gasBA7SBFMZ8zBYUFnWu/kIgVbTGL5maN9oxT
mWiSuog1KhzDWT/l6DW6+Al2CU/rxPqTe7iY3q1R8ifuRPEa86QxzuPjb2Siam3I
2o64bMdzFXk3tWYqClz+xEA62jbf3f8xmTFbQ7ZOBUcvZzCwUxGNO603RXPj6SEA
UcmzwgQfotMxnAmDLnofLeeibGKvEn5VSl2Tme+920M+v6pEoZg+umE7sJgHFr2R
kr/OAVhejaijo5yIhdl0WVw8/zUMRWDVhvkYGFWZLxGILg3FKofS3kzrFSizX6PQ
i9eK8LGLjKyskgDpy6EHeVyiC7ct7Uy2EN0bMuKbl+oMHdlL6s6uRURtPVI6I/iY
ptx6XfZ/2v4NMdHEa1fHlfIluqz98fdmO+oEj9WdRIJ9fJEPB0HM1CgFxZGW2Dr2
4RC2pWKbyxVWAApTfHv89csFv9sRlaln33XvuMs150ga2fuQ/gnR2PvBDHB8gh2c
jdMf0HaOAMACC/LSnBvlzga7icW6u3yg03qyIvtdBTdd72HSVuyTW2pD22ttrRIC
NN1iDpk+f41nQNCPaKcRF3Zxgjsid/wW3GYDhsZ6HcvqA+QmdJ+P4KyCjrIroIbm
CwPw9Jq2YwIRdvCCuImlZFKFhcDj1cZJb7mqAIViIcq0qB3GH6zbad8qqEuj5jzN
gpcolg6LDgB3I1NjAjsWfWcVSoNw0/HVLUlLCsaapjxmqHUFJ+R0EHwTAVJjsfBh
kR7AUmX5cqET4QeI9GFG69R+ZQDO/7gbNoOEcZ8x1oiQJl+GzdF/7K8IbzUN45cK
B9kvQmvmQgFP6IgwspV6fJlVUPGNAsuPBzlmlgp+JSHfUj/NRihp33yjUJeMIL7u
Z8M/WOWggUc4TyFVjAtqAAbp9kDdqRsIx199K1gkgR52JgzaKtndJs7XcldbSHVY
dWBebz0yjXAuvGp3Lo8cti48kc065LOCzzQ/uF6B8VsWbSBkPAZRpws4Gs+YI7zm
wgy7ocp+iU24RomG6RmPiz62IdkMoXz8ZK0mbT5BjxzqKgACDUyB0I1O0oQpMmuf
FmxkC3rVm7yUR6W8F+mKS9JNNH2dp4+mpIAYycR5WsEn7HltWpAKAZGrRPBWwrJ2
5Runq36dnaUzir9RtikaRuebO2DimCRuia1Ac0MnE3HY6d9WwlYQ7lcmJnWJfoBZ
zG8LEia6N2WcTwCCQnKDwKYYM1YywlMVoHmw9ebg4vjIzTt63wYHsniHeKZ0vRMk
jCWfhyA1+Rri8j36NWp1+g1DgfDToYzM/Lz9ySh45ItSVW7+XpAtFIVgUT2+E8GE
yKRJMBIF9ihzcpbye7XsX/5NSJVyhJOzutACQZ6Aweqh273usauR0ZFuVSGZIAdA
4K+Pap/TjgL4uwn3vU4Nl+IKTVci864sPack79jmCnWZBcNjxHuQ5qon+TlG4aF0
Ra+qlBtb7SUa5/JHL1RAIOkpGxf6SXkn4sjxAm7clJpU8FmHz97PAWVEMJU0+Itw
7VhzpGTJN4L1Ly0ijtQ/K72xX0z1oxraMcjwgWsRdlJryg9pXHOPRW1yWgjT+PEJ
TQS6KKB3j57UGda+IwXzt/km0QhCbb9IsLBA2KPWP11gtBY1x2jWnVYroK5iz2JM
9OzxYbp57LK50wubPHEwZdp8hlyVdG5taWZhyo/mYA9VtT9F+aih/7C7CQtxNY8t
/fdEJaU5p9K9CecS+5ZFo1Z9CzwK80a/eeD8kUup05Ec/NMNg2fhWrl5DNSeZpuM
clni7yokA1OhWJNREETERE6CbvHBAwVJ0F3rh0v5CUAYr9mdyd0iEXb+m3+smOOq
AdZrPJFbxLN4C61GwqCM1DqbBrz0P5DZWfnQc1GlFOxn+T2Kv6l8NsTuJMXMYZmv
8dnHTVNHdHLY1KGzchdlJvmvMd3WfQV8oFXb4/2wisVITgcLLGlVIB8VskgAP2zZ
88Yo/SxSlsgVwD9u8HgtXnPsmfMDYA4alOqFEYTdZW0OklSPehyJ5PVkZm3tSoz7
o4Xz0JFLPBqgfakiajAm1kFcuiNMSlFCGKHqN8t3YTs9WXIBJN1bIpMTAlrj+SxX
DFQTGebUzAQ0D9V+HqGFdakze0Iv2ScCtmc0P9Ru/LPfzT0c08nFeC0G4IIXxWRn
t3y/D1tw8rKUmXN/mt9VZv1MMVQIQuCmzevslZ4/veWQvL1/2Vy523UvoriQJGha
vH47RiMRPo4b4WZhI2riq+d38/DQBPVTuFR363rK6iTkpMCCNYECK03SNeXqBvjN
E6Onb6gLctCdjKuQ79eP6O/v/V7twZzznYBJ4CRntuaO+UXbzOFET+vtYsS9dpKl
5/jawabKTSqx4bxOAhdu44PZuufFGewbGYst5Pa0Y5QZKkPPZAm26tcRnfEsyJ5c
STiPFNhlzeAoi8GvbF83fwhi3jeXfaAG1snSGVPhqdEIs9DhO2OnKQCFiF0HnXIc
uZomx7hn7U046HCycMripeZsgeJgAp0ZXl0U0qD1oDTRbvH9mgYSOx/uEqE4gPtz
mgi9h9z+3IptyAo7brUA2OiEy18M4/iaar4AkIE94dkUOUdrF50reXRYcOVCZuke
7A6qT8ZG6t/gIqEArQDJZGIFHy5VosxOSURi0ixJfWBbnmWpZsMOK47cNfox5rIp
snnG9Xq1Wfax8AxG1XKY8V0C03AudmC77cn6WsKlFT2ne2SpYpXbK6byJUMEz+SU
9Y7u+iRWBqEn0rVA5enrcX4683HcNOSw3nXodW7vNWQ+u67rAWv6R0/OrYSdxAfg
iCpI8FBm+jPaMuInKfuA+FcCE6uWO7sPMIls0jEI1uz//S5uV8FnK21SLC6LBokJ
EAGaTgbGNmQ/KhGURgNMzzCzdI6eQx1Z7f4fUtpldfhvh6AZo1WoMUDn2aIwzvf6
MFWCWTSdhA4iEQCvHu5fgCbz6nivNt6radPF7BTSyfkCsRiGsN7eaUGot2n48jK6
AM1zx2tPaTK+/aVQmpkXW6rhVW5znI7lKRuHnek1yuGk3YYbD+e4iIwOb4hxMK1J
Tdgf1NtW9G7a4+NT7B2mHPgbaePOXIx9TU/TIhqLR5IjYMRaT+Pp+FdEJJaKl+z6
lckMbXCPiWvB1w2FJ7bFL+0Ix6NlwB6WlA+bPT977PRmXQtiRQtsaw2YR+rvzGcM
dbpJ9ZAzbk0ir4PZN2tSjLn6rgVdvVj5+a31WFy27XlJg2/dwplFal1kBOid6jBt
2xc6Vq52T3tFhue2V9LNaUU3Drq+RhuWv8L0zeiywylhDJJlpwQWY8lvZZUdqRcJ
4ryMBmZTW0h50xTimO2W7Ckd+JmuY2LrwI3C8NmFfJZ6pJ4HVp0gbsfFjEa+gz7N
q0DNwUFB10MiOAtMm0ppCHrak3oQSeZrlP9iZ1aR5pcr9nxSwGu040X2lAMFofpu
4srL4PpdhJmJI7t3HAJrZRCjU8K0S3nK1CUCdza/IcGFtEMBGLUKGpKz7BBHHihn
TFEk7FWOLLVtY3n1Fswl4Sf0Hz5r/CLg9UPd2Cl2ojF9QoysSZ1RU0bg5SqEI2As
1zPfwuQAVFC7zqz0+ZKef3VoZCn8ED2bl9VjUxx5LPe+yn0ldSmPERV9PUDij3rt
tpTXnmwH4IUEIoOlypwGoyXPsrIwaksv3HKL2Vnp6TD75oGd3jgLWNhVcOUqS1GG
ZF2KdA5I3O9G9kSrjUWJDn6wJm+g0Dz4Y8xgNMw+xw++KzmeU0GiPWcNatngqWkF
LE7QLbH913Wo7Fm+llVy7INrHFLBERBMG2bAFYVOdDlpYiMcklwwWvI3lAyrP26m
5Gwzl3QO/enAcebt6nnG7KNlUYmcBq20XmvBJ/Dc2TOkbgSCNi1Jx91xdaz7ySJu
Y5hKuEa9icahKy1eQsPBlGSwZYIgqaDcEKkgYTltin61qNcN+eza33vc+wZAxJPE
8tYzAaYnn5KzpYZpe0xDzSTe6pgPM58P3WWhYFrkfaBU9dDw97Xv6dKA1cILzPur
SopWSyfX34olhqoq6j8KBimlfClbuKYbSpJjgalRwULJhPVv1/EPwwXzGd8t84AO
iWbHC51cZ5IFTSn1WKF/6nutlLk565HbPPAgHNT1s7jIvuK3Vi1/PkwH2c+y3XTN
ThJkJ4/o7ApL5Fl+evQ9SFNDTwcJaoFuwdrsNDRNAiqRjCg+i+kTY4GS4cSVkm76
OKIpugBuuatMQagdFO6b9R2YOtNPxfrND/RQq5v6PycUxI68cVQxojkVkgtOCWoY
m7xcYhahRuLd/BToIiX0bRXkH+7XsXaTxePe6KnBjEac+rd3KGDRzy3hutjaa9Dz
PXX54+UcziO+qXVPPZOUD/DF73XSPm0259yLdE87kYwZNJFB9IfguEaJBi0s7l07
MYeCUqrYb2Z05immXOru4mrreJ0VbmFZao5UL5e0DDqPMIBoMLqYo5SCgmC6W/gZ
SYD/2Y/6ReYGmR+Ylm//gUimJ4JuEi6iep8nkBuwVKxYlnjb54Hr7RwPVdBSGuf8
QKSxTPDSjyloWzkoNoTE/Z+OGidyNiPIFkTx7eJe3EuVB07IM0ym9eMeZ2QKToLK
fEBmaxELqoTSuoof2V5AGFBVOz6SdHH7GUcDK9lB/DhAp9sI4fq/QGR08CPc7yAB
RmUI87LgQf0fpnTm+3i9ncs+h+3PYkT3/jA4NEt7fc8b3pByyWou/oWtt2V/0rKg
WGa2LnOjKRlR2b8JcXUjDSzo58/eT25O6e5eGUjPE6xFgzNo2Gh3GQbBVkyWV1w4
TR23G9nUjSWnLOEWxWxrGgqAAYWq4BaWg09WY2OWXeRi9cicMfCG9EWj0uShJ+Gu
rONi2+ed2A2+AvW65/MACeDyz6Fh8XuSJL6d/T2Xot0IP1Fv4NcECsW8OAmNBdlj
LVFgUyfCx1hLifDAp/8nJ65ItI1mL1jCmkNFzVRGLFDu4WYRL2NvkbgT/lPSE/M/
s+Hl3/1wxL5JXMjpSFWMF15KUi/SqyDDFFfSttB8cgqC7JGEHCCf54DanCil9+k3
qG1TbVViSTQuEentD9eQ9L3kAZn7iIgPbWQzCLwW0T784fdBi03AlwqgXYOakjBV
yFevImjkKGwMqozVH+df5I0N0TstbO8JREPyY3s6qmz27BE8z59TdiicS02RifQx
ScBdLgeuC6wXj39eyujshZf4oSLQUARB6qEIPk8fpED0MMwLekpzKhH30EUSQbcp
Q6I7QzM/X9TpCTY5GAKWFAiKcsN3JeiD6WE9x/4oRivkhWHs9At3HYv1kL5JTZBA
0nDMfahrpbGFSxJAUQ4H4NGK8tT/8pVC/BCiPnRZKpqtKuqmRHLCv1XEzcuCqROM
sum0+c8dxwMeqtTKP2CJxQeKWcmMJe1JWV0bUqg05Z9k+zxbn0B/rRSGFAUoThfT
vPFmwqhuG7cbO1Z/EKmZo1l/ckRIjb3fBats4i6eJQI6hKDtn113UBSbBjfSvczv
4yfBD+oKzLfE+9uGh3n7dURXRGpfBaTlNGsMKGgGO7wtl1HFs2SI6/tU3rpi9XJt
Gbej/Nd5sXFii6JomNu6ITkEOBVAk88Ywr8dpvRWczVe9pCNgxO/PBbmi1dNkjwD
kjhIgXRDSo5XVWHhVLetsmkSxnFdBtbvDTN7grU+IVOOszofIDlRzMn8nK8SWC5+
DhNkn1Q4xfMTgkJsLhJK9GqsijngQdHJO8pKnzXFs1AX4KSXYavPs0C14gyPQoGz
8rkn2Ubs4/oIj6sRYgpdGUx+b81GpUwAoxHplvhsyodrdniXPXk1IteByiQ6IQUC
spysEamtWbFZbhF5vOvgUZDYM5NYxQeGLtt+AnsyhIbCEpbKLYT5KsUYx+xW97Vz
CgbjUfCwi2IXaArqyWM09eChVkS4G9UGpVYewtrl2dCYkX58vnbPtQWAqBtm/RmD
P8kuV1uweRy51z5LL82sS9ruB47gx9ZG8nX3acs23x6kvPtEIvfSeNNTkKWwEr3a
c1UGVHHn4C5QcX5lsuYlS7w9RQqKLCzgHMYZUfV/KC9GFqLUH6Dnu8ltGIKNbUfO
shgR3B3HSHepy4pF58wUls1fGo0a01bMlEXz5xZgoj+MR+O70RJAeVwp2hsHBeEA
0zAVSu/9PmHV419t4JDaehA+gUR/7wtzv/rNLu6F/wJGDRuMvK2+DiOO3XfPTeHK
SFxHnRYhfsjk/ZBLdWsAOWvWCG1rESG5FxkaJiXcO+QbviKOXo+0Qf1S2j02yx4v
gw8vulXwhn6XtUmRZRYnFw2YGEq4ixf03LOv+AFSpS0fDtygdPOMNava+7P9DvjD
OebIE6iooIysel6clSQ4Vm+i8Vbg0aQ+LUv9fLDZ8JiLn0s4dGHlVStAkMtT3LHr
NkxxZ2DlkdapPysyFdzV45POmDBLiscTKxUnWdiUEdhfBCiDcrdAaP64vgx+S8B9
ruzw5mcaezUMdtnXqFs5od1fXO0lY2s0O5JWTbrlBS5WSAt5VywyowAP84KdWPOi
YWonfDJ1oG6qK7v0yD3ZoRvgf1FWGcHP9Uj3nEJC8sNU9seDzhjKtLNGQ/nxzLGV
ly3OO7iV39fmPb+q29o1sFv8q9wzaM+omYfGfJ+TcfWW25qMEBwjBPt6vVPU6ECv
FMDm22W7CZzGgUpIu+swH/8BfgYcQPpt/KJvipCzdiNTmsw/unKZfbdXXyEllC55
ynRds0JND8SgJRsuvfDWi3B+R7QocUr61XZ6SAY5GilW6HbDJ7bXUqVkqH8/HJTo
ZFwfYbzSw4cueqbHJKfHycyQyYkfilRM4BDEYKoOouieTLo0YapqNwwoqU1CnWgr
JGx6Pf5d8OTXA64QrBSflsPHc1h6DZ98p6wlmFXpbv4w/wcFn4XcowthVp7GwjSO
cRKTyb9LQ8MW6VJg2VAM3t7EAk7cg7lCPQywOhFpJCJrslsm9WH33j6wwkvFiW0N
N+07B/+XZW7VWz7G6xqtICVUuFkFnQ9CS3L8ym9LCFDRoNal38ho+W1zKFrPI4ZU
/QlEpQBZ38krdFGFn4PqUIZDE09s0mADHXuEwWjqTTt8wanjy2MdRiui1yhCVRcN
v7cC+ozJt8q/k8UHo6QugZWFh0xx+c/McYouhe3Og/RsDo8R52H/KPZTU+Z+j3gp
S3XYwYTvl8TJPIiEbQLw7li2iablDszNhHipeQxTJ1BbmfzoMXXNQBbhDmvqZabr
MXRcQfCRQ8rl+cOtNxMYrdggxeV+ts6v1YatNmwKfpu6uhsnvLovsu78K8ccnYNt
YzK+uFkh3LL9XvYNC5SA+AVGt8oGk0B20PyF0AUbcKgorCSHYsTyfGoCT50pqVtH
2vZb8NBBZukIbAl5RcIbrGK623dYyF/NsyKcAzB/QCqtZZrGcu/L631G79sQI4Qs
wFAy61ph3PWuJkHTiLhqqh1/mlLfzn/OC5+MYJuctqhLj5vFAXV4glliY0yxh3er
W1Jy0pxYEQUABhLB1JnhtmY92nuMLEfzBWp8knjGAmBfIrunSAKOd8EVGOnleDbG
tokLdMuqkJzZvJlDiraV/Bqc2pXvmjoh68ZrhxPG4bHD8pbnO4DwiS8YSQvyGwGY
gE1eVK0bfBf01LhrWsqrniRc5CJ2Y7b43eaU2RbvoZ5Gd8gJCIRd5iZWxuBHdQDi
y7ijsttdqalkzPrjW5VdsDPqFaMuoQMJmCmPbQfJ8fkJvphfI8RkkO9qRmFOLTVx
bpt1eNurKaGZVF8BUx0Jx2Wiq4WElIYLObSNu+4PRrF/p0E+HWtcQsPP2HqmVU5g
azMjadkeXPtdpOIzLZKttM2jik3gaugWYPWAmWfwPRcCJsIPton+8cmQP+nW8lQI
vkMFpQhzGX+eb2mIyJW5ARn1hW9ajLMl7MsPOspEOasU9qxjADto4T/h1b5Dq1Hh
LM6nB6eGxAdphBaNFxrG+bueBMX6DlSXITjHDTPVkSqDdIq/SIe4DN/Zona50B+8
9B2oJEqvFepZOzpt8O7lysCvo/+CD+cO9DrO58eNdkAYs0FyuQk2478NcbgCUyLI
KgRIDHqHKwUATPoA3Mo0UVWL33MwPDKoR60xr5EJb7qxZb5gryynWkVazOzWcGaU
paNy8eKvT9U+LvyemX7wW8Ji2WESDOCKycjNCafRxg0Wc5tl4GMrBERu3m0HlxbA
BU9IL95w/CXFFQ9rZyv9WRCuPcPaR9vn5lKIYp+6r4pPferA7T0SmhzEfnYg2BF2
QigFbFXfA1DH+QK0oPRlERQ5AkyfvC6of5IuLkGfzn2Uid2YNeLguwc9yNS5sYfd
BmabWk6Hg/DbK+TEeOSD6N5Mi7Rdp/XuArcZTomAZxrCX3JENT7pi0A4eqPKU3nn
SVVgeOfM6Sa2VM+jfrw/mcxKXaK34tZn1cCd8dlCJeNMzH4j4/qtmvrsfuQE+QIe
6QPDbdpTafmHZ1uDFs6dz4cqkiZ8Pe7GDutKFuJIdVey4crGRslF64OluVCmgu0q
jL3FmBoEzBQSiW+7k91iJLUnEGC/Bf7YcWvX3OaqxKQxrHw75SFDkiuHSbZvxnkH
qIVfPM7VYfmBKWZmwYu/gT8ReumI/Wu0EGoHGlwC12JEG85JiPXT1/oO/FHOsFKY
H8nmv0jU05PweK3N0dRFDsQi7ZJfwaUPchbd50HMTPHV38QdIgLWSEWMgO8soN7a
AFRleCzwxNWbLJkUsIbjzWNhbV7uUI3queYsva+XgFnSrFOTk9/b4ttbbYqaFN0d
dH66JKo4IriIwYjTIZv3wBUEoQwE4A/PE0EC/AGZA0Hm4EwWIbzxUH2KVIu1eInf
+3CN3MwkiYfacA3HR7AOR1P1Nyy7Gj2j8Jgn4XL2aTsWhSwkva5TCyC0JoR0DhCr
49DisCl+n6PItWLHUQgaTGWBzkV6NEv4o4b5JzSN+BFVocjBo8pd0DKAGduyyInw
FMJTCqoBtfd9Dt4IK69kZh+6dtLtpmhejMYlDsgswFlB+0NiVqAf27vFdUMqMkKV
UvVP4AZuXgpTxxra8WDt8kFcaFfONyf3qE8fyzNEsAA4KLJGljPBs6A7B93grFCh
hLf5zxHvTXmq11Pi66CiGPU8XXcv6dH4rvmDG9HS4Lp3p/xAhv2F1cQKaDO3LvXF
6wMyoq6eFsyARbG5JdYi6SB9zHUvpUGu9SZhg3dd0UKPw/FCsjKVpGUMFRKQ9B23
xNgy3/hwBzkfoDFBMjAoOj4hUa0L2K4x4l8aJ1B6uuMQRHJ6Fs1Lm7bGDgie2mN7
jh9T29S4DbZy5h3W8yg0DuN/LzxGrh2aV5go7Ts0z0LYq7GZQJC0Df+D5kkWzdGb
i6tTnII/kC4g5lffPGqX7yRj1C1bS6aiYXRe/dLHOSqg8hENApYXX4LiXNzN4csZ
IzPnc+ancKjv7cXeKr0V+KQ1egPj1giWzfT7zeNgujmshOawNRiKD4fH29uidL/M
JAK4/gwsVQtvQeD9hBitg3zx3uYgplPnf3q/KDUW/SE8UVCPkVn5BNpY9tEBJypA
923xASbkLcR79Lh3CdsmmSVWr9T6JejCzfxacZkPN9ij+rAXsF+WLbTa6zpOmUvC
4yPl5AX+jgb+VmHbtAFv+y24MSVhjrEsfBc0tUrQ6r4tUOFryvXq0BJe1JtWU8Ds
6fy5uzkCa5Bp1PWT5qumpNAzLgcYiign4eZ0OHo+NvP7MLu8lyZ9FxmQ+5qBhnTK
ODzjNh8eHgt1tjOhFeVyPXcUJr+H6d6dS4EBFlHEoOclKgo6q5CXVmkOJKUQ1Ddv
DudMHrrBhn3ImymN+SUppmjolSymB7qu2GacxLs2gekX930BtIJFxRJefbwxKmlY
JAIRmrLjSYXXzbYLa+vf+ePmXJ1iqcz3S+bC6vXRXK3fbWbb7pA7xM6fsnIGFpXX
cw5kndCGZI3wVH1zbrG68LP3SusGSjVXTr7tK4i52j3VJIH1rCcNxi63Ql/xbq+V
SFVQBFNAR6B1v3iKp98B4bkZuCa5+8U4vIJWtVFXyCgiIs8sx7drUtpAjECWK/mJ
InRGqa96IwnRnhNudmvVfKZ1Am+Ghj3BDyQsmr5lfhtgLRE5bWA8iQ3LqDOgXRon
XsojEMEiBekqcIHiaX7B/68EheyZN1as7tVR1W7Tz1bqHw5wTHo6eu9KrmfOUQI5
Ij109gQMOn2dQWbw4i0UULQYZd2DoRgXmQGkWUmN6MNAF/rhamfCvgwZ7O55bsyC
K0jBQoU37cwgPZDvcA35WQR1gF8LI+oVTrO21poGKUd5F5UatVqGmBCxR5aoWRFL
A+0MedMQF3rdeJiQ3eqlpVei1ELrZ9r1Hoz7DvFH6oIo9xIpg4HfVP8y+6FEn4E9
gvTi6XJ9jRPFuvu7EKb3w9xekmZbRDxLQ8u5283uDvieQxIMHvDF1kJgZt1y024L
43XwpKEfKZshYGEWBNdr50rOgMIDHqmrfsuBDVuT+tW0UXTSqWLcUKX7ptAPrmiA
D1DTexKodvTX6dL/8f3zUSSkktdG1jjqz047F7WAmpYRYEJDQOf7MEI9QcdALSiA
OZcOsxNMtxLNMFrKeRt2rnvDiKuVigWlp/f9mU7fPLIam/y73iWqMWe/gR+u2IrT
ZM7U8YjLcGIvO7pB7ToAx09/xbGcEh66ajkkmdkcOeVUaEjvY6DI7ScQga3V+3/w
eZ3lruwY8NVrfjN9ZhXmoixwfQnj4CKtl00EFsBaIo6I5mmlYPpVbAIYj5gLdQnu
GzbXZAw6vpuQP45Gc1xnUVbNZdV40F6KSufCclyn60QVZ7fD52fpiVwvi2mTnY0Q
mbXUh8t95lv5+quo+nvGyDSz3FecHUpzYRJ9b5yCc1M1vJoOS5wZDYHcR/atUVnA
t6hA4vawn2y5oUvVGqcJu+CofPnPF90yapible9M1lAJ5SlDmSX4aecvpluL9Zml
LtAZMijLzqR8BG82Rs+grVV36lgbyrnJCOcYWgI0l4mxcHcMuKZSK6q05PazUQtR
mSX2EvUeaLamUiCBXqN33E9wrSHZc80ih8kospQkvxJxTk8N4/LRyBGOKlW2+NY0
pPuRcZdNW+JnNcImP57juRNdI2JOGhfynhKv3rJR7T8erMc8fCrn9f25DXBI0k9u
rVtc8tixAWn/QNMOTaoLytlWEJXf7O/TQsckQ/gCGCyT4goQ6ZRZhT5i63w9OLUO
lzSYN42uQDQXEfj3SS47BdN8kLIlQ8h01NG6FjlCbVO3qSy+qjiQloIUqdQvBnrD
POFjlmmikSDM0HKTKqWoWnRJTz7OccUJn5itIzhcKn6O+OVsOptKsg6354gH9dqr
y5Rf0YC9RVpgM43JwtD4Loj7nnc/zT/sFeVNc+bgV3Tg/kgEgNOd/a4BJKNDRj1S
/wQm0/VQe8c3bchbaxGQ/CJLkOgaECnO5KH6wVNSJ3E1N6jW6fAojPmV1oTXzxaV
oRELffVuAYeVi8FzS8eh11aVJNbEIFqRJ5tNPvoO/p8eRDJBmYjiEZ9SsG9GtIui
xO0flEW6Bau5U4OfTaqW4sAPcJZHAR8HqzhqP1UqsfTGiZQAB+MMiW/C0tZD9kGE
agbU6gbhBAt4VEntbB/5axotcE1vtYQw9Ku4kc1T//63M0C5jZmhea6HzCsIp7x5
w07c9cW+/lQeMhpmryM3jIwkr8JFlQg6giFeP3kIvIZz5KURFwhXxjvJIS2oAE9D
IVK1rzwFVRHVdQmofEf2x4XC4dMdhJupJNgcWo6YzJVWohBwCVBl/7Ne/7VnjS1N
loEzOZDn9ABpa6tIezeHbAL5GlSFDPXBYqGhUhqQyRfugTQ2cyPZECgiifvLeOXy
ct5X7DIxQ80cF/5vs3r4fZaJmQSKQsY5q5kxomksf8VwRpZT4xM7s+wmKQjr9eZ8
3k2R65KTDBQ6y3UphsC3ISpIs4IpuZY48cULEF+vyB0MancXII5JgGohqFPW6B1T
5Y7g3qs16UuoNo/r9m81cLh7Bv5ipqZq1CNZq8cFB9UC3GGdyCLQaJr4DPtTvDRZ
WtgiS++bXZkdhJTIValQ7rEz1ZJRQiJn5onrakZyYh1KwvQ1Ky+m86h4M+ljaE3Z
8kFzEo1cBmjatgdGm+paH7bdu3aSR8Sl/P87EgF8b4RhZjmwtQriwkrxgAQGBnDx
BXcv2MTf3ZfnuuW0UC8RlZkXjufClu/Pp28INs1/hxLG3GGNwexKbD4n3IF0Y1XY
+h2SYsF3qwX0nMYoKCK7AH9JOBmcw42GnmFaE/6t9b3VtaaGociSLSjP2zOFG2jg
1CYX2Z8L6vntt91QJEztWkUn5Gmj0G7cMuyFcmFe50F2WFG5epBmvE8oaZGpxjn6
F7nfVscPyCYo8HpFWq+e3BTYM2KlEwJh9FyuqDPgdmxuD2xGjp5YM1mEnvWgV5BD
A08FKzqVSGiWjE5n72QHiFHN/4B1MYqC1qd/NaeDNHpMuXYmZHDlryGv2GR+Q+zs
VJBxjNOjlqlJGR/pyid9RQpyennsishAVazlIAq9eVG6aSv1JMPx3WZCGYSUdMkH
94NQDX+pSk6iLj1oe9v7DtcYPFeMa7DrY5ZsCYDWYrYzeDG3j2xA06SVqfxGE02S
F5ETOJcpP9fcpQElq33Cv9NraQyea7+8TOYoVTVAmIitGLXp/QUK9gse+qDb0Ves
vsvTlH1MnL2xtX6rr+gwpyX2yBbYf4PH/6Lebp0jq3sy/8Cn9h8b22b2GPGMjH7/
CMqUHQCxqwfv9WKC1v0DCQP2ZP+l//im301Ko/R1qFOxKKMafKhUyV7Nr/sAfhE0
vE1Uwm06Xp6SqAa8ZqWpUGPsQhbeT3ccafFyF4DH8q3nJH+shLeJed1pIXe30XoM
inU9ZU4n8MWG0mcPFjJOd9CMLJeooyc04d86VIJfCj0xmV7sgUjG1zP2B/fVwVzC
sjc37hwXYeWWzafxKWiTuQbnl4PKepABlaW+amAQ3QNCv0rY27ar6UelRxOET9IL
+hvhXRby1fFCIf/LHqw49xpy/kKWI9nUXUHSDSpgLZm8BdMo5THSxSqhbUvxMVo5
TbQfJYrwQLTzdHImeYYPGM+YN0Wz81SSMhzpVnQOsRL8ReHrelyrJ/d6+l2FNcPK
GOZMVohGcAUiR5Lqr/bU7HULb9gg92zkQKzBCE/oL2yPLkDeZRk0HwlXfaLW3Vq6
j/zD0GYA0NpENIasBsfu5A66tGJ/sLwtul5bPCfaEijYQVb2IliOZCPQmo+aZ8wM
pXDnWhlNOyNYMvFP6iqHxyztyZzZb20Zx+p3ipwt9Sn4/w3O1G2o5vtcbPJwvPtJ
hxfzFkos0dGR8/i0zGemY2OglNQ/jT7pN7aew77yCJLpu+AHErLQ3XVl3bju4uQX
HiFyGrx9GLRxSWjQGejVzAkO67AGcWq8YVz52qJl7v3r6SOHObPKva7/2pn85HF/
0oc7nx44A/WOTmtKN75BIfBTYp89UZSi5hlqh7RGh3g6hQnZXgRCClZute2zhUQr
LVZ+oLlmD8zljtHpaighVauvXbb67/R7QIz6+hIRRXU4Ms+hYC+saRYFypAK7S/E
qd8aZHW5bxX8bXbydYuK6lVZ/zxCdS0FWA3b/Zwxezbld2tUAcy5+o86+ACi+ZxH
cpJDzpEGFgp0LaETCvS60URZa765PCZi8yB9LnuEAeV9RztAaTqTIflx99Hbqt5L
KKHK5cd5fqKfMIRceospB7Zoip0d5yYGD9hzgFC0lNX7S7QCysRvgysWuIagRMNz
BSI2APwe32CNSgKe5lTY8fLHf+ouIbRqr7deYosj/p1ymtXkExgDNnuDj3Ju16JF
qPz7EqhJDbHE/EaKqZUMdlJfQGutEegCMsNrQDtQjuWnI9UBqAThYtRnq3NJpdYV
qdHxeNbgf66rjl7+SJaUDd0CUO/TgcQGFCu51u+/alPTwgGgZFZGi1Jv0jDcDFTN
NxGIE+jhmyX/2ncU/6qwxB+HnUj3XTfeq/PBeu94jDuRwcPaHYet/xy7b2ngim1D
ABrt6jw3Zmgbn7dHxsVQxxx8aoAODWonzIf63kk+YJ3rEtAB3XvE1daW/DGmKoOk
PIYX8T7v0P/4qXOSvXXDLk01WugRmtS/IAEJKj6Se0FXmOw9nXIeHxFV5Qt4oCta
VDPJ0hJBhkwDji8ejKHVGLjH0jQgiCeOlFIx3i5F6TSXAVeLys7hye9Cys4X16dl
sYr/cz2Au4jXhf9eORk5AlUHX5PXrPdVVS878cHxbL5PZTNy6SD16nl+CpVEuqlf
Xj69WF9Dctx22o52cShWS2j9tpsew7OAn9ZNJbC9IcIS096x8ikjWLkXUJh4DT75
9wvrtT2ZqX4xJn0luxRwC2+6Lu1pdn6rSs2RQK3c0jbNqQSLMeZqwCjnrDXEY8P0
Ev7h3eWBj78xWj6uEFDNId8X0gWhXJaXZnow0IHjxRSJPU8xLZj38jE7AOsRzXKk
LX7Dz4hC/xk9VqKJqztra0h+6nRLBc1ooA2ejzl8C+n++A/be6aHgOHKjRoEhyJx
OqVH0KFXvX0hfEvkiDZTFsqx3mQwOXgjhhuNhuRjSKbHPQFOX/gPbE3BBTewiQLV
TqC4TuYZ28kFAH5kNgeHY7ZNRHpev94uSxC88wjl35cLr0v21jhS9cH6JeLWQ42X
VM4tIs1THlLBmXXoDQ5qUgdzEpFdF8jTDpLtjSEJH+CMmmCCWOUM3J3YDJxF2urK
pGPSqoYJFH+M05lzYS7ug46wHJOg6Zowgb95RDpqf37RkkFmpX4K7jyin++MjxpL
/om6pRKspJw1/Q72NET+IsMIfnGNU+B2ALxG1GtoaVlxjtL61gAGx8czzLP6xveZ
QY/J0zkRMJ4z8bR8CYp5E9BielA4EHeauoPpjoOhXWx7+M6hp6X1pFK5m8lp8m0t
rfFSIMwn8qtpVUPIdJknyGunWAvuXWENJOfG5uLtOXro3UyiQpM8cMb9TNpIhK8H
9FeDXb8o3R9YmuV1RAupymgitu3vyMCYRWB/5QM/RaETETkUqbCqaC+ifYrEgg1J
dSm/Uz+A9TFKjObCy8o+iLjGfLMswlR71E+IpGrpGFEd22jFvcutOtW3OrHYqj/X
rcOuLoL5CQFolqdzoXUj4kK8T15Pdwouf+hG/L7XWVy3htR++DgtkKEXBYr2mLY7
k+ga62TlBTD+lDKzj82qZgNh9t+qKNsIVNx7V4qXLtz+ZXxduvHVMm7alZ9Ce7wN
OmSFwsIzmCcrUgwAdIUGs6hkjheCu5XpAJKYTin843JmGC3PMdSkjuyfWY1dciW5
Rd0g6kyU3HBQ/9gz3vZKK+RXeFQLcLTgBv3RNHG4ZOyKZPLX056noh6nHXC+BIz/
KyQxPDSon7e8VV0zDnIndGZx2zgPHvOb1/6DCpTsy9WK8wJByc/Q+oDWTD45v+Oe
HojbavKYXwttKq2zG9Xz4MPjExjwiRGyGmY4ynxDLoKJeQFkNicxot49ityGM6Q6
1vHAx0Ds9qhljGFrew4nixsmpkHlgR3RfJnZxMpv6HPd4EZ7wh67OMBgD306regN
YDGe4hH2ls8S+gN5pcTHhoLSP52pTmlom7mfStZBcXZZnLJLf6TkNLpyCIdHOFti
ic70epZOkSuUGqv5oV2TyLRKn9vPak61Ep9NuBvVcyUgVOtL9gRK5Jq4yySjluHV
BX0A3JiOA7+xUB++VgqTbHSn8q4O39GwYkg0z0HDJHys6jo0h6CiKcUgkreAjWCe
W5xUimbWE0UqpKd/Br9CzYQaGfHADgZK0r7ZfHGVM/37VTqo2jdofYpGYfuYi1E0
ZXY8LCPV/tuhohQmoBu8APp6ul3uCW5GIin53/sBh1kxylNWDA75qEOSqPcp1Ha7
fEoeO0lJKXn7Z06RnmXs3Pw/Di4UhSg7b+aEaioo0lAOMmYoYew0ye58DOHK/Nna
7cHDAYUBUBTKixTRkNgdKH6FNwq28DRGpuplB5nYP1oLdHO7TCWw3FBssIbCgDRz
07TknrDDtvvc4MCko4LfQBfH5imgWfYdxL7g9aFcbyTnLkPJpEcTSDPLhhC/Zxo6
o9uf3krLSVb0CsK+2N6dunFIcX7bl42gOIChWlql5sb32zQAFKwwjAce1VrTtU+X
um/xQzIgb0S2sXTEDVa7ASPAVo3ELmbr7Ij+WW27x/IyrkEbo8pmuiWATfwMEFhx
7O0XfOVmfAlicjhgWKz++YI3p01/vM6hJkZf9EsMoe1Ki2ZOhvGigcbkn6dfLq5/
L9XN0z9a3lvdqIq0npuaBUNm/nBVpoN3MJ0jWAdrWqQqn6EjQ2630I96JuGxwwXA
43wUGFL+4RepyYK5aCCnp43pO6IvgBEvyqHqXo0h+o46pwTFIYvUFwARIZ4P539r
fktU2/5lKC1bLUfJGA7HHQqoLVG73PPE928QGSv+V5sW9voEvSDAMjYxvGy5f8TP
kB282UrkqxIk2Tc7fENQq+3ge+/9mjVBaYy0SDgrYlmUf+PUZ1d4ZNDUZ0+UWbAa
DvHvZRRjk2YXK7wmtx+P15m+Tu0D51iZjTnfblK/zeUP35u2kBDFHzVlIAKgrT8f
uTdybC3oYkVaP6JHbcAdkoJLda6UnPn+EXHUwUP8GZfUalU24S0HrANYCgMUBGVP
3krZpIHuZtmodQtxWZemgNQe/YP7u6Ag6eTFtG8bkzzQzO2Mj75Q0nmy6PVve2XL
E3gRioy9FRdV0xgFpbNGcQiIDFQaZr82gqh12FoFbLbuN6i9f4xkq0ZXHdeuzjlH
lSA4sCcNcZX1ITNsw5TtulYWPHDVmZBhY4xwy9ySWo3A8FehTwdqtY0Y66+Xnoj4
1LqMxAgmRdf2E+H1w7YCJlZqp0rGzytwNv5dHV2WJsrEPzxWluuD4/OCLK/UNdra
wWK3YkUlnYSicCbYpAUnDxEk92KIVSkQk0/ISJeyRkbEhyXx4KXFZJng/Sw8nKjx
PIBJ16Z8TwYfAYTiT/LDnOKZT1RRrdb+cm3HXp4tl1F3QT5UJXLgMAa89l21t/UN
JPCD+Zo8EFgsswa+9uk9mXAZNTwdtg7KMLJKNvdPRuF9Fli/mr2B/iWjVX1ShQik
78jN0fSFnE8FkcmrmjozsDUjAtpzb8xlWJHaWUlTJM2KSa96fa1I8w2qxnec4NbP
Hp8OKjq7k1MEyEnoW1ZDhK0Pihe+JgrGpdiSkWlTmduDuP4NGH+y+IsANEFDTjlI
/Wf3W2HbuKJ9uwG+PZ9qg4IJx8KZQxgMSnoweyiAe2G6/H16clJLfO8XbXL5J3zc
TNXFdh9Nz9NZYva2BSL2gPZFE31YJyblVCqWsP/ARTpzIGGqRze177DA1ky6RyKA
g2ryCWUX1yZSvD3nukYVRrVHzYBAuYdYclRB/9DWWrbIDodHT94M7aExzXEj2Gbl
bzoxhIFRT9GFTOJvd8PodySsnFK54aj47iD9/08dg5nZdKtZ30LYfkUGhzAz1mGu
kshYNQ+kTlBX3vxjiqbyyKghm1d8AouD0veHspmnK76vaVYHvdOohttWZJhV/EVA
6xWxcAwKC0kicAU7EulXQG87/C9ppUDrV2+sqBoHoe/QwCq3KL7br2sXiNgrkrB5
yCsWBxAJ2NpAhnQbLi0MJj5ceUEf4bHRQJEPDDrxkQSo8ihz+MlIflpJR17P4EV3
N0tlPSJPOkZIj20E6pCbEKkIKCIqlpgFrBVAAWA0Dbd12N/DBp7A6IuGZhY/TlJm
YousL6e8Z6I0cebR6DsRgm8JJjIkZzlrSLKI3ofctWRg4A9ClGTbzlA8UYTNNack
tKaUijlfRgHZnIsYAieGdTgiAfJuNOeF3+Pl90maa99O5IX/EyVtqaaGnsLHZiIX
u2OumAkDFVcBZtuz4CKe8gR459bKCyk64bA9iSaz7LqGE94RZgkBX56stVtyDQHG
Qq24QNJ4vWf0LnFRzBxm6lDBo5/sW3cIqd36DA58Z2XRHdubq1d2NHJbjeVdYLIt
RtbYReimNSI6Ec4plePi9T3cyh1eyK+d1NJc7ivlCorWrJCs5/29SrEA8vUW3q/j
Zbx5TbIXB39bUjYI8ds+qD+wWY5c9WyiYzqdA1AqMXbBz3tTDpqyfm/QNdkk4nak
cJ+TWHdPl6YjPAoYoJu+jElASTjzPFenET/WM1rqFQ2c1b2Jm2pOKZd9GPOsOuDO
RvUomyBBQ8ewN5bKPziHfQLE7YSlDrYTEVLm0SovjRqQrfEdF9NVJm+O6xOszXFB
j2D0ehtJ0lcArUkJnGExtuNzkvjPMVG1aSYjGDlBWpK8YYhQ1LkAqEBqcxjfvj87
atobGJjWf+1Fe3KsGoZrquIyHkSqP2IlK1x1/bJQ2LLpm71INQ6EqgikS7oKFWy/
9z0nLSbcC0LB5Cg+xfXmKlPtjqR/FRhnC9h4RH5a52DW5IJvQtu5XOTJR7ulceLe
ToH9X23FnG7UrVvnR90ecbkSTx2PE+dKUp3/CKVVNPJ8Eask61sK7v9j12mMikuW
GQA1euksTAunrrnIm0tXjVCAcPNK86LdIdxSElb9e4mGqcR0OdnJbXQoVSeg4gZN
kEowL3KGVC2oISMeoXzPB1moJstprdFa1/VQWJFcDDzJoK+KO1lxa/5jaIdyfNW0
I3B/bqEoOaRPSOs09N8tOqfk4zoe+ugZbJBpD0E+PaUml++T8TwWqZx0qVtQixR6
FaP+MSW+db9Bu01wZWz5sNRu3zls2mBkoRdcFVl+yECbeVsv0Dc6L5uKlSbFpLDS
i7PonS0ZQ7mne7i8Oy1YDX1AOHIDG4ce8wNqpN/6ucQ20svz9HgPyMVrXYFhXr8G
n9Q5zhg5fuIRy/mDAi/3cuajHpJmboR2TBPuCloHbTWKVubXke+qbSxzmQrenfZ+
hjPaQ61aa048kwjuzWz43/kTK0I0h4seV25ge+izkTA2s5klf41gqcdQ3Li7ZdZF
V5VfIF+72L5owxussZIU9Yl8E0iEqJItCshxiWpxea6Z7mwTeX7hFfC4bbXm8eNk
i6GwM1CaBNJUggJVY+SItf85259MjJwBizvTGRLJybeyL4jj8g3hUtZGl+8KcL6M
TiCbyb4NgcOsKOKf7PSkLMJnWLHiCDnZIvdHXf1TvE+8/2jGKBiEVt1DFn/tudPZ
LWVk7FDap78wJ7Ei6dUrMDHZBN+mVC8al8O1SZgk4wRMQzGE/wuJ2mihAMiShtpr
s6tL3+LCZKe4WxFWeyKVKqa/1FZrC3rrX8e0odJ+El60xkfBYiZWekg2Xjc7zlHe
Vh7Gu7ladunbcYYq9DKLdNsunKlKxTor3BjcxrWDfjNo8dqu9xFS70u8Ruknz5Wd
nYXG5Q8B8TpxShTR8eqO5WyfuRo4Kdfce8SygfLJy7tMA8t0bXs0XKlYjL2mDD3D
4NtfBVFyX8AclV4SLCZmFbTzFtWiW9akMCPsOjxGz4vhU1rtoJRQ4fAOirUkCmrC
32GeuP/6f3zn3ec6DQDQmFgx5ia4sXFxucUPb42Gipc6V6VyJRXDFgb5WeYEt1aT
+AWKzZ1dUkQ8Azr2QAFZ6qx2BBpUIR3Pzj/7G/EJnwhUoQvjLRTcC6cJ7g65ZSdV
wVs1mNR7GZGSUD+3RXRvnQ1uj9OaMMvhNTZrG8dwE6BCpBeeiQD855bm3c2Ej5K+
8Ed5PoIl/FFRQ8DGe+/S+M1MTa8eUAjA1taUFeZ/qHZNFh2H+TlMXkCZUmDDr/Nm
p3jt6Ctx5xZhf1u0CXt7UZ1o/Rj1T1LnfqWhK3tvrtmSF7TEBEyIW3xz/1rXfCyy
vRtechjN2Jlj4S/gGwQpxmvLUPaYZwpF/jH7ndCt0EIgV5s9glqpyEWdjX61UlQk
CcQqgmvzujbXEiw5jCzh8hqLMs+LjTf2Nit2py/RhZglvMM4tJTjXy2miTOU2gXy
IfJ/lHX5WuvZixTLFOEgKY9oAqLU9K35X0bBCuSpV/cPb3Yi9XyyQcXTcbvOlOfb
Oe6hGdE3utS0u6yt0B8B6cFyF7dEgWs4OiOQCHMui7mNEjAlWQ++nGShdIf3DpT3
nSzhbxMDknFbtI/0LqogjfXeuGd2b1G9etmgU03Tl07GWWbLSQY3jVGPRxt6h7A7
Z6WWtywFBzoAyHWIFD+NTLoaUHp1KmhVAVVl2uCk0RCPYJvdfDgpGj9P2Mvmuknu
XsKNH9W0TZ6ggcH0awo2AV+YOXWH8kgp1upIJ5bylr5+goIK0VaRiPP0dW4X7nCu
z7vQHHVomPXTLuqJbA9Le3Z3DEkdIB8zBO3LX+7X9RekbzkG4fWydcWWBN8nAGuN
zw4VuzIGa8smGwwGeZHOJY9DWj1WY5fQnCVW3wLtrruRW2OI1k6NEYSIwyyqMzhJ
UOBSiuvKAPHbn0wANcf40o/vt8MBFREdNOqzeaQKdf2fRHnjTWcH+Oi/P+wmQATX
n5Ya5+DnP+twX3UfpwQvie/x+ZprV+g1xBW2GhZtadaSMBiA4nbF9u/oj2sJzcWR
B8Qicd/r2W8L4M4xTKNeK2CFhmcWXyj4EAindxOq0USMRiAe3UglnWIxYov+JHrn
Q/85RSZ13DInaVmF7/fz9m40ZkWheO3BcAd4jCZwrisHJB8CLA6Ua0N3arQ5QXu7
pftJVWwJT17h+xc7IZw6gnI4cpIu3c6r67LWh1ehHPjD0NXo0JG407lAZtI7PMMC
1FNXZKtjUXdilJ0Op5HYsfV488VeVQy5gyHkf/XYyiMK7Z2V+6qztN7z03rbDyQC
eshI1kJHVN4G16lU4If8Fve+bFQVfdivriUO51ReuRXDt+fLpUToXf2hcd2Urf0G
4c3kwfw8f85cOhKMrrHAqEGioAwcaaKYRF//Ixs+I28XpxqCXmGpiqvKM8Juj2S8
wliYDwQbjGl5JZPE5wF+FLOQmgQJGd4Q8p6+OXiKrftdvDZCuw0w7/J2I3hqt8LG
i1/KLgv5UZgrt6cz8COx7eHNxiL9BM/FB6SzSnsoipIuvBa9CBrM34kWJIaFukT9
YCchjknlDyohwwJsNBv/lXlvddJ4p/Iaf9ZbMaAJ+Tnfy79T0cl0B3+Vh2fPUlQH
yW2qWvF1LMFMj+V/viH6C/HCMXh/nJPceCxfwFNSIz52ZjJ6RCztdgbJxTREjlW3
xk997eqHfAU46KmhLpUcIicWjVti05YXR6V0bVJLfeBy1eHR3J3w8b8JnwVVLCZT
7m2T0WEOs34RtfI9fMIdpCNEr3Hy5PXvD++qi6Y62k1zwNOVx8l9H+fjj+kk1L5g
Jz8t1CGfdiyP4fg43QaBSrsnFYb5kBnjzKUATRZFwJXNx4VWae6+D3M4yBjjE+zA
m+W1UgVph3mq82jMFFiFIvpM/8MMaAW7oGmilN3J1P+CjmK1MHmF9xAmJPQVfZlI
PEm/f82F+8qc8XOgOYmdrK/NPCJxF8YxTqCaMoOAGNU4tFYT5A6hx4bvXkiBDCV/
wFpxN6Z4T2WBx5Ukj/YeLVDuDkizIgYbLvuKD0syyRtT2CFjtgRRe6nKKwkaDrsH
6ipmzAVANmNXgvTm5Hx7q3MrXWfIiJfVSZHUJVriCDSMnD6RRcakUSgfVshbWqEd
dHcGM0DwTtTPlWMZC4QXxykY1sbgfIIjDdmge/S42KbFiOcH+p8w3VMAzF+I1Fqt
GKJPyfPwgLfeteG07qcl3LEjZN2dSqSKzz8SfIgVtcAzzhlGFuyyZB2mKll0jVgd
uhz5BLwBYHi8CXomLZRC+FFOrBQsD0OrA4TiWI3C82D40Vh+cxope4nLUhSS1lxC
UPZOS3XxKepZqaVOS00RkWYDLD6QMBKhjokLoNokgA1Xw9l18p+1zVWDTRxigg75
dP/axgvI9Q+wNAyDcPhAfQtSGTQ8vXAFzwtNgtyUUG/92jIwmRPwsfZj9n1CLayB
88uzglue4V7UX8vFUwAyn6atOvU8m9NpMj92O1eOI41aJPYpe7WLamwYy+jYN/jF
ngBmczOI2b/o9Qw3ZXK5MzUl9zkRnGGspwFJjgiDQlLdU8b5/iEN6WDXxnaOv8Yg
sz1nyrdeP28+n9/DwhiveJlutQMFOYnLtd8VCsdZPu8lPBR1f/hY2+j1nwDjBepG
2FDgH4ru2KsU+PM9qI1fU2zUSHHr4Z3DnB+7P6iE9RUEF6b+rMp9wq5/GYQ2z8T0
dpMTqM+F9tDO+j2Rr0uyzYVseQtp1Rzy+59Cx03p6Xp+zfTZYllEmKwkHoZU4vUb
zjNRS8zVsEFLUwexfAatNUwhFdVvYf61avIaTN+IGQQ0U+qRfYH46hltujm9NcvX
1GDqCjzQ0h/YBEI/VykkZRnHMRiyfVF7eO53Vl3xdSA7XDMQiWobYXaAjGVMHWR8
bcxZopxp1MTphjMYu1HHU7uI6cO91MuTG1XrM0dRKaAQlMh9c5bm+D4poGE6LnPd
SJNHbi5nRdkWJFlIOT6x62b09Q8rqUd4cvOvGYCSZjlPRVJgd4FSUKewMT94iN1D
4i/TSUt8aKO9Fy8aq6dgHfL8qrLBhs87dl3ciJmuJpwGiH1VepzDm6BGzuYt62qB
rMHYSeqNODrm8e48/fCz4i8RDZOeBgor/CEy8dryh4GD/pMny03VppkiWVRQs8R2
8Zltcu/Bs5R3Q3NeqcmlJwpxkRpGqmQuB8xgMBHNBXvbLlhYIKPyAedI6nT1Cp0W
huUJQTSNx8XyKfAaB2vGcj6/WSNplQpcQ2S4nOTWpkhfL1cca4idBYrE1ZiUrazu
OaLk6uHDiJINjEVvbrABI5zGaxOZDlECY6YfsUNV7mEHVHDfERD9rKt4iyp9jCB8
GODEJV6QtWH+Cld4glrxsbiQ0xawK2SKFB5MEbckE/yBKkVnR1L3JczuUoIL5gv2
CiLyUU8eOjLTlAZmbfuBBgv6oTQ8gxUgKD7T0c140sSwAGL1gbjErW5CYTjoi4x0
j0pDBOtXEGQYlxh4Rgf49UO1BeOnHyJTrsxYQ882m7UAuh7IxZhhxRztKuE3LodR
Vj7A560Cgx2QOutph0u+qhwTJnjEZvJ4BoJ9kWy/l8kxI4nHw5oS9noRYNO+3yr3
Yz0AIv1Trz7Z+W9hJdmmVkwZlHpseR7UPIIqQdz9xkRA4cCpwqNztkTAMSj18LI0
qboUP5GOZDr6FB78RFbl5bA68cbeYU7RZKMiuL/XpakGfV0g1b2oY384oNdxO+Oe
7f5nKljnaVs1EKP4cSvVjSa9w0wqFa6qscgPJkY+B8bKx8WVXO0JXUFzGah0nD8M
45SJgMq2lbkg/IIkgP5LD3SVE498C6SpkP+ktJdRQT24ymRb/bm9g5tQ2DC6R7CS
xKEcvYojbnSyRYo/c61A/LXBBEMHqlZWc5LbKKbvVrqv90ZFyb5EbYvKnSvzLAqW
c6uxUs9mY9fQQABZ/2/YjtKhTeuYl6oivxTjNDCS1xd4tIhkh9/gDoi7rlbbSkgj
/EWka2VbStJsmNUIx4/wGiMBWHzmLl774nISh/mAQiWWotEVYatIIwqAFn3M1N9Q
I9JnPrEjELMiTQriE4RJErsQSYgXS0n4CEJq72jR7dB3Bigey5uISBcBhwg0ZsH9
015DuP/IPPPhWL0xRxsdpn9hjkZRAbOgcv8ugsK+N4SloaNLOgeFnPJNXl6gnLw/
LUeAAoSpg3j5dXYb0HUjweZ5xWxS4OJBml/73alE9zl9y36bsWtyxbTj264dVZ5M
oLgY0GaPscU9UdXd31nB7ZGMSCuiqe98t6Yacz6YYM24sbr244pK2N3Z/UdbSW3Y
xuQDujUaJFlReDwTzR72ddJjnGeElHEvexlBTDx8mx0Dp54k/+VR85ikkPh5OL5T
of7G7k3bitpY53ckIR0ivg5HJiKkf6ckq5j1xkB/76TLXuMUCh1i33NNiar6qT0N
RpXiLMHFt2kxHF2jGg6KHXDlsJhe0g8/XSd9/NCVeQecjzASa7heoc3xAtw72uSw
lNO9TeEQqpALSQFMNAJyq7jwfY9YyHg+HROuI56RgzklvbWYY/VDpqw4gF2oxeoO
xnPMmd4yWI1MIbcRI0HD44zzvh8O9xJ0UZKC/d1eblRi5Jlxsq/kAJd/kyC5SQcW
mBR2AKJrWUOqWkzRPwzplI+adlinP/EaOJqyBJLiBIuUS/RLcMR/BNeaCb3lfcTv
Q17DZU4shqQwoSh9BL4imk6EXlewYR66svzeu+NeEZyRlZQLixl537vbrkguHJzU
5ufawSwacSG8qDpXD7OradGTdRCTGi7eHC+Ps8cH1QsheGOxVa7fGH8OPZy4El26
ltjY3QKwTA5V8J1LXBIAV4pA47u0ztdZ6k2usn+qUsDDTmawz4+nLsH6TfcmNzm1
RcLHQzyaCm/Uh0Epd3tNpR91Vp+msh8r8XQ/xoaOD9hxgahreqwUMhIi/z6b1jTw
WxYzp7vLtBsdkVPB3yEsByzVuQAlelF6LN/I6CiDi3iX1U+dUfIvpapelpM4av2z
X+gGffNBZcMBdixpqfCN8hmUZEMl+iv0okaC5can2n1e/F1Sc8Qyvedt58MtzCOB
2ZQ+GcUisXbdrJZHEmNaNQ08LuWoTaiMnlzAHP3VwvTY4bKHPr3oKyvYBv2PLGn8
oP/7Dc9ab36XaIEW6zuk1DDj57l9Mhp1rM5wcEp1icI/WzOkYOhzyo8TdmokyNaN
Gmsu5aLdtMw0tmcDGrxos8kLEo6b7TvPKWhCkxiToXqugq/vhA40RcrL6cnN3nX0
UaWPsOK9nk1lyhwUeubdCKxCNajqeyb0+aO2ELp6YccheC3nAK1gN/1DvjLCBMvl
+ULO/+Rfz7GfyLH1/UlZHg0ogRwXL7myyJEIwWRovAqkhF4bilE3j/IM/CsF1JNn
ZOLNI2V/S6rle3BUcI2oYg/DKef9S4JeiQr9J0NcnRlY4NEBgGERiKPEuvhwNq2i
brAO9ob8aRIJonjYWlRl1ZXxseCYeR9Povg2mxa2xCJzszyGnyWxKN3O7PyVwR7b
hYtn90UnrAbiKxaDNM6wiJ7LQl2QyKGZtETpQJNbmtaMZkLSVeBCy+D/bmtjESiQ
oL0K11qpiU/FAtzfPBFn0l9MB+GYxpXv9Zq51nyfRDn+J9MX4N6HMLlJNo04AYzg
RakkPRO2I5WOv9p8DZdCiqtRQZyPlEOIFjtQSSlKUQNa9+BnxZdoNjXAvIRU5Fhu
3uhnTIPebzIARiN17jCe/dk7+Lh+yRzo+Fvwx6ZuL1xQ/NlemTZvra56ErYXX2nf
8HQ4THCE+YKrlV8KXa7N46IeUW3BEH/iMNo3QBDClUu+08HonoQEBl9dMIXU5yvw
5P0BWFLtdebbbjtjVEsT3z4lYTsnI6kAC1onTcmUbUWAxQMam4AGk01Wq83Wq0Kx
0xDeAy7WyYLxBnuMyRmTri7cnqsdqrE84H9bahGTIVGSKu45VjrEhfxPbadk8Pz5
osi7ml7yOVHWk8I4KYRPx3LKbsXZ1mhu+469GbVFqHE/szs2Q5FjI/Hff5+6+TZA
87JJuO1ughlcwgNXmrbcp89AsQKz1DuSYMrGQa0nimc5H4K5Yk3Q2jWOIY23mybJ
Ba94AkG7eNKKpzJhb8LHGr5ZcjdBMq+B15rbz9PYheHbDgJtz9A668dGketLVLCX
wSXPe6TXg2CDhO9aTfDq/SyAlvb6ewaMhQ5mU6+nAAEAISjSlAEkNf4XriBn/CLn
UhZrgTHxT2RHNl2dXtXKhfPy/VIln0z9hRcbVrOjrMFkOTZOOuN+kYGcviJK1E+f
IR7F3MmsymXdtLHW7v4f2f1rI/s3XehqyS+xFMrbDvyRJyYOEavkjNW00406Hey/
2biDhID3IchR7Dwyh7q+L+dgnirSL2AP/X57UZ/NeZ1kJk+tdySUYFNoVX45ao7r
9QovXu/szXSxwXXfDDddYpfqiewoSgG/kK9bgiR9T2ZgZ6cl2yGnznwTEYKO++Ww
e65rUYTpaMqJAtSE0RcLhbeNnoSb3oeKy3VXABfH2o7Nb57qCFHqBXtVBReEHtzk
28cdz6YQcRxCp+kZk/KnhCXGWd03mRiKq0KZBAurdtT8DEJ/MpZCJIyRgKnGe8ji
qDbn9SEfVj7qnUr8E2tqXvMdxs76u1JphzLhnWu+1HQpbF5kakL84teAcf84ntYl
GPffi5uuqgCW4FDOQLkwmYWpueR+F7J3P1eb1ySEit48iDtxGSL4B6jJHcx4CmKY
T/w7lgwNwAhRW3yvOQXB1NDxuCFANIgMq99Hvc1r1vH/mFsb8oPzVzB4AALhXTEa
Av/6AJGEO4YN/+ZU8qM7oqHCeDGFc7tcwaz9V3r8JlaNToBR1tNxRj2qJfbcRYaP
GAFYML+Z4uvrHwgf9czX8m8nUtAqwIEgjLr/D4LyxMO/Rn/DLDKKNOQjy6PVMnqO
1qDHDrBVJ0NR0vCwULaAxZ2vub6RYDaVemFT/v+4C2f1aj0EGxSCuiFjGmrkbLrS
di7Q3wYWx6qtsUBSxyL4OuGGeJVC0zBBVz5fI3nKWubUixJDwWPk/Z6iE2Hc8y0x
RLkoNZcI5hMIMbKYkrL6ScHUr45pHu1Qa49xk1tAeJJPWZ8blPzMzFmteldg2OHM
UQWfzFsb8AcNjtvvJ1YFPTLXWtolVwC68YhlfB9v5OQhrL1RddXGsFh4XjeLSGiy
jdaEZfiG9ndxvLTgxbMIcTRI+TzOm6CWxLYr4wi13/jdSZcVdx5dVr+v+POdaO0I
IZVIUUkXsgdifs0BZyyTajNbfMY1fnMGjX6qCX/vUjdYEWCckZW2p4mElfNcjNGn
YrBzOBWetoFyNK3MjW7OVkIVqJWkHZHTbcjoR1Y4oln1c6QBS70vvXHjJ+TsXYvh
/TfhNOLjZB1IpoYdUlk0s9EEfniscDWeZ7cjT3tqtycd98OVpOS3F1fcJnsTeer2
UDRancYZ/grXCldhj0wSLH07/awikOyLL8tjfsmX7ASmWHu+ojA/g3KtFr+jvSHS
jUGiAo3pDd65vG3rY0A3Xm28bBSJyBTFR0gxglQoZiRjtkER/PeOg8ZOsZ/VsXAt
TC1wpUlSdRbJfnb7vN8kHemvU5JmUs4GVXUtgfGc9JjPdJ7c0DJEYAn+QgbAnBPg
YRLhBAFYDGwxJb9KYd7FEmqV8WswUrpBaIISXj52VKAUfWJOHRUDyCkbM9HSs4SA
j8iCk9b67YoZjSGvGKxmTXetNuaOGtzzm4vD2Hs5cgaX5Wnb3MQK098l8P+lq1Zs
EmX9W2uOe4lFMS7bfFXBUUxkd7jr4EKQRwAgrM/zFokdKclK131XDyE29/6bYMLb
hLTEq69fDCDou4o+JVUUKD+Sm+yOjijnEtco3KWgghmc4f2kKQ4d08DjUyRkiN8j
7oBxtJfUdkG8dmDqGC9+CREQ7krdF5b8ln39ViX3nyVlodbvil1/4b3cDl5L5ZvV
LR7acMWOWmQcmNh1d1vdulHAmwRv3sjGM7hwHwqDH76yiKo2UTLojljwYgu3J+Cp
C0MSxj75IO/GvZPZJc+g74Z7E2BUxD9Gqc/qBAaxkr9I46+XtLevxY0P3yajykTf
1HNEIz9ani8UV42czjjQsOAw1elPfPQQUSuAkaVyo3yvU7jOBc0hpP15VD3ZpAPz
L+79R/w4fwpOmAJdF51aIuvEFmcAH/ZplcUF6T58F0b5wqheZdDK+bYZatnm0U/b
xJ0ZmRoOdR2QhDKuvNxwVbMt2L56EviA22nDyv8bxXTAr20zBTOEvMvdujhH+Fns
6+2elSFQI+1nt1rdAWCi3un6GWF1EJLuLiLwiKp4THAwY431aGyXPSxOlirK81mz
0LRZYizjSUEISmUXymFzKG1PWfY/Y0JvqJWMPgmM/AcvRvUKhGONQf6rlxwMizgB
pLaNxv3evwfxh/dAQMXmvIyaWQrCon1G3dLMZzVdnFfyY1c7nO9tB+/D4cUtyjJP
zQ3hyFt9Zo7HYWTBaeGILST/zORQBTdijIwqOVbQsGBkRZcIQzaRcZjgzUAgMo5H
fU80PZ1Jmgp3KAGaFqrWJF1SmDI6EmF9vhMe2SLETZ8y8OCTsW2QnwgKKecO4ftN
18kpKosu3wna7CSzahUYVFncmD7xCkFAD3WPEHShAjGk3kwOR3m2Z5Wt2c/N1uh9
yluinvPYuL4c3c0Wi4rgyR+8vsCIT3I+hEhw7LQghGf2iIifZWottl3tLkqy3Zu0
cOSdMVQJdjbh48ehDtQhL4N73TEKfB7/p87NyzzubGsfXIfR5/wnvGvsXojhHrh3
W579FjVpxPr6JnKwgGzxaYrOFMQ8DvVaWPZ4YWtLek40MTF+aglf9zEvd+iGk13w
B6iaXBwxg09oet3uWpMth7awjtTvUf9Tpapypk/qft89sWFAxQ3rrPkmuVOGejxk
D0LSzQbLURnadKaAlRNun54ef8BfWbAZSPtBTJxLVXoG03GNhK78t65XaydG6p9u
g9CECYHgurAEO1PGTNWM49p8ZfQfm6T71tyeYpZtg6XLzmpxDs/ZjcL/UQ48fSOV
qW6Mbo2t3IF7N1ThdtYIN3uNPxeSoGUPSPHHpXGTfsAK48qozHYutSREz+vTPkh+
+GKvkH4M6hzl1VWPFn7IMYmcz4lM9EOVjoVpvi5JqUv3QfXV3Anc3adIZ8CvygmL
Vm6NMPiAuNYdovxz+e4MUBZ4P7CqZQNJlAIwjkBsBpyepwjq3GMfFb788RKBm3z6
SOnE0xAB8ggNp+p9731rI1aYMRJgD0+/mqkBOe3jYY8kLbaCE01e5GTeAsoHEydQ
qt3x6p3u75QKt95DaIB+9Nn+3CXz7iHdafl2QJcfIPyGH/6nf/Ynn6fZ6sLyfSjs
q1EYpuxaMy8CnqcyvKb/T8YE85CIqbCAEpraQ7XUSFHJ34TUonKyZsS/d8Cb5FYX
2pRw+fYFwZSdgj4l6rDJtmXECPgjaFoxk/TudKHd60xmQPfgJK/WM53zisJYPqQK
VqmHcaIXDcDgtCPmB6jQPgKYfvU6PzdFw0xo9+cwo4CAZAII3shYIuikS19K9Bh8
Z/xO6r3A8Dx4Qt2TP48njq8SZJ7FQDDJP7apCHav0vWwcr5KIRTsIDTbZ9ok0Vf9
exfoyTI71Jb2CZc1gAKf0g13o6NHEw6jG23VTWHADgm9AjnOG1bc5DCT75mgkt1c
nrd+Ld3shNl6Ccc01yXQ8r/ThokZW1MQUfJUheQCh52BI+2qEJL1qeMAPft4WMhl
L/gkvRlNeikOn37T55HkPSbmHNO8Q+1E22LtKTZQ9kh67IxmQKOt3as9DkHojcPi
P0+aMQcz7ojufEniLiwUjvWi/tBgswYTRW3+n9myv7SZhLO6H5euJ1uGj2FjG9Ek
phXu27hD8vSZErKKhp3Z2g092QQcXNUe33WERpHqEdEpWukzyTmqsgBIwLoRVZbK
JD98rvAGCxSiKudtiH+mJ66PQgS+aUiJUnvU8QkuVOjrRNvNS2cTDCWwCFvda11s
+VCrrvtwx2dgf4ZRiRyFj0fWole7d7y9cME4gTji1GwbuxjdxYGkHhFz5XBFHL0h
Ob3XOKWB07v9w0/1UDixW2Xj43q+VEkvWD6Bcvp6e9MStrv/O/IJ4NZ//V2ZjHMh
/TJV/3gcRIhAMwkx8BdYMl0BUMwCFjzuI8viuSMEri6a75yZyxwH3FB8QIyBFdLT
DL+l18y+ra1L2NOb9SCtnS27j4lDu+F+UM0W2HMY2PXfdm+Vxe4UY6sVO8vuuuTb
sd//9oUeDj1Pvj8pOWB48G6tPR+RNYGMzAy/Be9OIieYPmQ/S+LxDlrpsUT/C4f5
x9uwfFgK8AooknFks/crc3qvpHukP9DZOmVyYk72d2JuAdSs25JIwZC8Dus2FD82
aAKy5SruiXSPUQL+mAjw9ReM2fDSHKro3YeoMe4bUPcaUSVZY1u7oTcPmrJcBtq4
/DsrRZVo/i6MfXVJarilfpy1atpoVUwb0WIwyUG7qZNQ5o4DdaY6kp4mULK0vk+L
/nsRtUNm+yVpOJG31UW2DrPajvSlu4X0WN/93J/73Q8mhfoLQ+aC1JqdGQ5SHeFY
sr3TGQk7089EZ26bKm0jhmRT4SN+gFdm1/CkFe/08hXEsfB1ELRMv0t5Zg/a0o2O
b2dyRD2NVEpEfRjfSCD7pXO0Tbmh1CExeabfXWX2HFEghLDPJNz5/O+bMyHjxv4T
v/pgwbzhEv5j+WWb1s11l66afTPt61/V0AJpxFhMy5GHHn/l4h3n7G4PUIJZjbog
PagOnuItkVFNNIwdXPEcjvj38lTt3rAUYWirhhj05KHDfHIx1PAKRiZg7/HRYCdd
rvd7VS/ZGPMMngN5LZmkp3IaW9vmnTAc9Jb+m8h5SDjT5pFpgtvDmKJE1PSXQmYt
411q/u4oI7bxR9m/RmvuQhzhZVRry51ZyE5Jfs3vairo5KCy/TjEE7mNKWltjJ3t
cKN3RjgRjVuSr8rD2X+Z/dSKMOMutwB/kf44dbIJGzUPOpjfIr2WjcGRjRWOZylP
JPgBk2Ex/TKM2994jtA+0buY9vSXIXMdfrAUwwhPYADCrW8gQe9H+2bbzxGA3E3U
BlDhUNMF9WHP/JFA2ZpLqMomqWpNGg7p6Gi99d5dg7qRxsLe+y0PK91PXBddh4iY
dsn9rliGzEikP/hZft5q2bV2+TMkhJS0rFnakBQuRdm1Db9NaZ7c/Cab1zeM2SBi
TIqNM3FwccRP10GbsL8VHL0jt8pQeeJgpWieM+pN64pDSCC23P/9pvfSvSf36qVf
Wh/zjQ4qkqYBcfrIGgsIZqzs3eUqUORW/pgddhAuz4X7qGZUGWPf5wo5mSDM3xkN
TqXUM02Q0vPdjNetmiOJgQDvK5npc1X9s17rmytjvQ4ZFPtMJ3uMnvZhr9HCGFyb
Uafc3RcvdkCyaWOuEokAWI9+g8U0KVgEu994TlQCJPYMAjMRZkA3J0Urg3AlyIku
9FleZnQ8YQTnEbRAEwrT3UFabjcz4eaZiOyc6uTVj6ptaTOcBRmQIecVL10CZ+fo
6vaKv1an+WZsTf93MivUOxn1JR/tjpdgkPp32Hc1M2+s0rf7CjfaPrYWk5iK4cHN
Ss+g/ffSdHDHR8ovcOyT0FRqrz0+RGcOj0McpShhyUZBw4+uyuX9mRUyfZVBCkxA
CpWOo/T4m/+ErAYP8hcvUauRhTRQb0l8jJJqmdQHOV7ypzvfNMt/tE3koP5w1eix
8nFjjykE2rHVZrRGzK1jkolx+tvTyKmiNlTn7mSR+jeekcVOIeEnEl2LUIY6vAXf
CBO0sKR1hDbPs9/0jIINKV6yqFVKP50KCLVQIkgdImqhsQIx7Vc54husBVvAeGdd
ghHau+kYLufftKNN2Yi20GkH04XgRkGjhsI4uIR/y7PMM2tw8NNtaywV24Io7dUo
70kEAGLqlfprOhbTJnVlWokACK6ustEPmvpkxVDcRSaJ4Bz89esh23hGFnq8wTbN
RP9P5K/NrE47vij8A39NXw1LFzvpXyMyatzaUKzBHHNplfsJIBab2VxyzKvPetDQ
t5w3uU7JyL3mrBymzQDRUVd7BnhLHrE4PBGUhIJXVZYCfTHTWz+E4bYH04PTTft7
+aRUvNTOHqFNkwk1C9+KR5fZCZKNasH6Ifny9sKLNdGnXCEJ5PSUJPIEW1C/E91K
1jRuYR5XGoWHozRMDSSFNpUM6lqNvCg3d19SyMZ345kugiZDkOYZIhH9LmNRYbRw
s/cSoKkepgOzbypvbUSz1u3yE15awhI2Gm2k112pXOJjx+yyUOwykDy4yyaYfoNn
8W1RRQFkVD2D7FNGD9nVNEa0JDnZqLT+VOxnkjnQU/YGjpHe4e0o3mS6qRalr3+j
+GF8jaH8+E+5pG9NOy0vQL1dhvmdaorKR6NnUBKyaaoK4GDsYRlRLhDEYkCk5bLz
xsB6zplXJIjXJ4+gbfPYtOXkOvrAWxoOmGZuZPWMI/Yak7EhHz750UOr+sIz+53G
4hgtS9UFbXCUsRQrEniWBb0k2G+K1RCMMBor5aHmbaKf4GA6hp2cm832IqgLofCZ
kslFpU6ufurrAJasfuTWIntoBarZcDxxDJSwNNw2RqojhIhSwOEnBGEQorpzJ2bm
5392JS+HGZQSkpSvRJ1CZGBzVMZLRhlqdUenTJ3li5AoDB1whZ7IwlkuNVdJ3rzn
m27oLtEfPTJvT56myl6ch1AivalelYk9velwIhZQhgbYygyyyqIrGn/FDuAqVo6i
q+5S8dvMUoYTVu6IWAUS9gFociwWyhjJsc7GUND7Wd7QYPKbK/7usBTL9EpW3YsM
eoHJtngVkxu3RIgkfPixFWBANgNczEUDtC+LS5MHI7r/CP+6FT4/QrUjDxCmDrYt
r7+z84odoXbbRUlhBId6AqehtJGugNVlZdrfUOTE5PgLfahLhS5u/aA2FgLFuTcr
lWEi8AaGVYtmFY68PUPFOTvRMSXK57FKRPft9wSnjwM5OVYxeIXfkXJ5kNGUT5HK
rzjKb7RWkQbJ/izMi5iCgatfII+ryowRriu2GO+IcqVHr/OKkQeefTYo/Ty5K5uW
jALB1gchxuA6bZo4pCW7RcUbhELmJwPKKGF3zZ2TFMivonF5LCYqcQie1Gp18w9y
h5GIHn/2AUqLjc9QTwbi0GgE8FzJ9TwL5s5w3IyWWsxpLEMjqTBnCPMyGMrm0Tkk
98dpJa3xjuXuXkrQfh2IMZxmZblJ+vjVVgJfLCFGb68J6tCvTybqPZ9cRzRLlE7N
17tte80j2wezhGLxP2qgxaEvpQdQ2+ZiQAXs7KSuAJQ67lP+sjyDFN87HeiQmO+M
mvz2JsndE5ska1Ik3avgU0Y+rLaVBF+dGn6QgsHWYUw+Z7o7bRWrqFX520jOf3he
sd1sja7V7nS23i602yum1467NWBFvdKL2Y+8REx+fWsSDLUpE6d6QNCfq/w8DBBC
1r+EqDIb0Nohh+eJQSQDOh3tMVD8ZADnKZMfa8aZ2fb6jan7HgnxjDzN1tEer32i
8SnrPzreEubLuj8omGcDeluXxxRT0ZiaqnOwAaNA6tD8d1F/QlLA5uJZTRZpGq4W
JzPq1nSeLaBvYAalWgX3xw1gDAyNPQCxualkqzWoccL1PwXW1VdvIS74FHe/NR78
Cep42BxeN/E/eJo4GG5ECrRMGnYUURtlMlp0ZvVmSEdZJFMKrg+1xp2OqZcBeKhk
9e5i7DhB/tmmJxFjiU6EDEMAoeOLlwxHxoDOWL6jOYhaeESHo9G7oIei3E3N9q1D
alQdDctObVnJEQuZwv/v5LepGOktA3nSoTEwuSqlzsJoG/Zvmhc00jrgjKdMvcGG
+d1RCJ64HXhvH85VmfiTVkAbn0E1urhMZXg6A3IV5P5OgxRyBwuGh9v8flzDCS1Y
pijXLd5WLkl3qdmUI5wsYnSOMtOqiqcUt1Wsmbc2OyV2++Zb2G3w3RsZTJyaWTpe
XEx+YZ5fuiTvSfHxthdhD46upOgl28N9nPaSX4RJP9xYIcaoefnDPDlY7febEI+K
YJfq9jv6tQetiseF7gjOpV+UaHfo2UvxxI+IiQady5uGp3IN2YB0j7Gr/89ycsrd
vK5fvxrr8A+SVpL27guUtl1as0F58QmCxvgXrnKqyvUvVCUuxFmk4yBKWuvtW9gO
/bc5Wt6uBgyrJGDXipGYKkiWHMGiVxyWuLIbdxMITiglM7+didY/2jpR9uq7qcgy
Svx7ANGMaUreR+CgLZObkMy5drOXXBd/F89HGccVMJP0vUht5zuygauRubnM4Vtt
yGTKMSQVMFz0D8DgOxAFYc2qLDvQBjF9iClsDB6DESgvFH/xLJaZVeH2hxhInmAh
xgOo7NZTHd8r1WiFyf84qXW48KfCaQ8w3aV69+xI+tOXCVqLTE7aS/2AR0mDe7/e
j4QNgBhFjASesTefUF92wkS7ZxjfeNH+8oI02+YIfX2GkNT4t3w1FVYJipE8qIJe
2HWh3GKclas286BsEZmbqZ3vyNXIt7kdVNHBRozy7jWV4ElB23x4Cv2o2jHGHeLe
RLv62bgWf6PS6YIeLwyBm/JyiTb5Jhi0mBOaqqgDEiV8o7XPo6EyKXia/Xw8j0jw
JhdJpECcmvnaMD4zEv4UiqW7MwTEF96Oe+BbuozTnanmCjwYP96+XrdDzWzMbBES
DJdIPvs+nYLb1KhpFd/kQc5GSfXtLynkztpK+Hf/PI6u0Ryw/43TX2342Bbztpns
5cQ/0N8x9n/39K19L1xQ5y58mAixttgv9jcYqxO7opNAimbQgJglRrhexl04npuf
y0ql0/ULRmS0+2lDA4k4KxzxrIUK8oprzPz7Pu+B8K6SZwnUPmZG6KH8l7psxPsO
E+s+SFIqnuqndLtFQhy64cFyP46f3b+vbchQlGX2PoG3g7i6BphgauR0n/IIc1Xu
8moo38sGY5bSX9fgFzNp7PJrGCTgxaQAK/vBTnHGbR4+WklAdWx7+Q9scGhcVxNQ
EBjhYSwH+1b1v4VrmImie8OUE7JuSW/As7Bf+tF7xf/SvP8PraPVIdZzIOvezSS+
eqnwVW2W8nrYHgdZMeod2Z6wahb9s/7dFuV9q2nZGEQFY9/NW4+GlU/v8erJKxnY
lRGtsDqb6x65+gg0ngYkV1IaH0u+gfrYAHjm43aolVVhi4wsCS7bg+iTO+u9wD3n
12LFAXPlN2bPUBB3gSEOafuXiyph6RKyEt6m+CXbNdVljn82NeMm/E4RqYR3aCti
S2UHvRO8269QNDVpSbFYGIo8umasydhxHRbL1ua7LV1qnNbTB7EFjpsbpw6fYYBa
ByUPWEhQ1jPjaOR8JMBEe3HrxVzWG5ddI6PZdwq351TkXOAIwmfVvQFwl32h/3wm
zt+0DMVwnqtzZLAYHWESxSWzbyLUYWl5G4+SJ+mJdLZv1jxHBHaBGS0N+s61tR9f
Hdn/e9cDcbk3ZPs2wFb2YryfFkVRRxDBZWJZO+917jmBy6Pi6TxacILdEJRekOpv
jlejrJCh1JmosQ1x/H7k7ndEc2mczsaiLG0sew9uReBHgCNfyUIbkrIDXytS5GYw
+i/fSxpvXUcUt++nbJg+3EIZkk2uQ6TFFquNsBwaMcxIApYdqwIZdLAWxepVLX29
M79VQwws0P38ypO56O9Tb9kKwnaRb5yffgIDUMdrYhFdRUS56SalXT54Rth96xXM
L2ZaS+YHK7F5yopCn7S0WhiM6D3Gzd3qLiThw+TY5WJCnzWbMF7Jj5mlY7vgR/YJ
HABhzR3OtjMBJ4DRWUKlkq/9CfwKB2D3VezClVOiAttM/lnrLj1sexPRvHfwwhg7
i9Bxyfoyq9ZKDGfQAn7jmV8mGscaikALwcaofFWPiOd3YDRIGMA39MjLpUaKiPH6
PMIhQZZifxMZDu6E1VF8Ex60LCDGaOupkNsy296DcLOcCXw006IBcRD7XaAS0P4Z
VNjEBbDiykRqRtrVp1hy5TNqUPGW25uQiMJprWYsLEAZeVy7YZIADGNMQdoqRQWa
k9sVyz5DARyryAaK3k7QXWfhlVY26OsbVCb3DPEnCMwUYki2UwMncKW0WiV5Dk5x
SZmUFsuoI8qrhqayaooa0PzfiQ9L0eIPUK7ObW6QTQ8juQkbs6r6LwQLWJpp++KO
F+qi0DaPX/uk+0lkwpDv0V5aJ47rXu4xdNWa1jma2cpczX2wYNVRZrsg8sy6Q1fq
oGun8ZfnIRD8TEwxsnGLzrNSy3dLd5BFXtC5uE/Ckj6WfO25tWdqqGxLzxVS3PG3
g8a6PTAwzwM7RzlhLFQFvGhSH3iZBcybPNygA4cgZr6gGxeyfxoW7PX7k40+q/cF
YaUnb8XYdd3fSYKyF7Z1KrmSoB1YHqDi4Yjd0mYLOH30EMK4YeaHSN5ewhIo2X7d
YQJmct2WbEgH77L1wcyGuW7fij88Z2yTj3b49BnUJODw8ID2YcwRnNFsXvORPHgL
2TNrXSFlyYzmmgfVUIFs4SmHUz/uCuPfEP5CwXfWOkA4Zz02F55kiVStHg/VQ92u
1yFFDJJWurHpi5tFuapPy6JuCEDAR4k5Y5fJBqMiWuY+Wgbs2hEgvufk8Mqihxfg
Rfd9djUV04SIZDB23w6/oqsSPj0H/uE6uc45w+8lGVybcEvhYsrIeOL1Ees8utzU
FeCUeGeXhMEfSE4i5HYWU4iEwYsEeDvGA6BFrxT9d9pIjJO+cn+xa7cOydHIN3P5
Mex+H8ODl9hOIrsoAGn+ORP/gbE0lzHyRN/Y320wArQatggqzfaGjigc5TdBBvqr
yVGjaFDi0WeZtsl2ceE/Uk7T1gLD8lZIIEtCDlacI2IPUqTxc1rTg2A6EIKTTSiD
tqxXGdFGCMlu/BeevHqemHEKxBOAJAsyeckmXueZnEONAuykVLMgnqkOhVFbtzNN
QIv1FKrHBeRgdx7ePYjzMB/1ekl9+PM9zNxYtZ4nNdlLzrfXmoMUqJNNhHkdTgTR
JO41DGvexMmZYKVrVwFwSDy4En+PwbtjLd3m12sflMx8Y/s6vGSr+gKRhWxwcBXS
zZSFJWUsIt5h7+8trhhCayO5naOrORF+lg0w2+g/nwbutty+ttt+oX9QKvY+yNju
w6Y0W3FiVViPWbHvUA0nROsfnrkzfIJEuzmJYR4sVqC7c1TnMuobZ5xzDcw7Dq9P
TWIdtdVrZkOS3aqaEVN2KGGMIBo7USmdswVqw2BmxQ3GsdxVMk4uMV7IfoAbfh3b
zq2dkBgxA1Vua+pvry7W2vzLLMcTuU1n4J8hdYXzl2FdGY3Bekjjq0YxDZ0hytpm
jqLIlRmPOdi7Z7yVjdmyulhhGqnsSmlV35Db96Ko5buzXIv907vOeY3tNSO6u0Or
8IJurRdFu2T1mEBnIVh+i41bTzxlasVbqjcCuT13+ne8ALO2vxln0OXKvPjTmFFq
eE4Dh8cySW8ohmmrMAoyTxgrCza5/+W4o2mF4eWz7Rc/4SfPYEG0Y+3TyIFAbRW6
atZRnhLu4Zz/nL7ologil1z7/6pEKvzFUMwXKirwMxHLr7UBsn+NAGT+AB6mlmzY
tZZcrr7Rwczi19PS86itJKiNai0SrNhXonN+rwPESv7poQivkzqmRxIlcdm8T5Vn
+FD2E8aFKqfGAt2r+SAuXFuog6xDalipzN3ZiuHw2NgMOCuXtfgWpNQUwAui9tFj
aXr8o4y/bEeEf1Lz8GYVSv6aNiW07pvhUnCiOECwZOUwCGG4Hx2G2iqX+Mi4XaZt
UjNZ7fDvSrPaeouE+o0OV9RGzQ7SSMT6zcqFXr68xzRJ9bzIWMN33vivH/wOYEAA
eU+FCFVdxD/VJAto7lftRKh9OyVz5B+n3N066BHK4SYRS/88sGUT3b43KzKg9R0m
y99dUYsTlxVWrTjYPijIWeFShNwxHFFQ9jprpJkw3gaDDqC21hjvFGyHPWfCFsNU
a/zHAcHN7I9zUwhRbId3stJkBlism4KaNqNtQxtpux1tFmx+vj6aogMoyQnpxrVQ
i89waf7bVh/p+l+I+frgbnKKg6ZQ3jDTsOMJsvZo4DXJBSDtRPIyEyNokLkadz14
sf6u5voO7nQNb5kexI2LKTtjo9Bkp0X94Ya6+9350um7TB+iyjoLqcPu5bqZW78s
cpfHG/ccM6LKAbcBzPt8Ddkog6f7iXtCWq3gJ6ofy0RYo6A5dui7akdXnINwLnKr
EG1BzscsYCJie5DBAdUp3vst+BDJxdrKjw241xgkeR43x1/gx1v0XHfjMwV34A7A
Y+Nt2w63ap5D641nFKIozos+B/Z66eVlo1KhPJMbJHuVUSbLCWqpTlkgoYKGTwP+
pSyfeiQU1MeT0xP6x9xN9lbki5KrGIBdN72be2yYzv4XPgN9fHbKlPl3NoSePZnL
I0+9hE443H9nWAlBIAK2u66i9JB0m0t6KPFXC5ZywA/aCpBDj7LspAIVH8b4Wa8m
2oUlF/hyF638v/oG2UXL1Xe4UUNPXlR3kAyWpwfJ/z6tB4BtrbVt6uyaWBL3SQnr
lYuZ5r4OZ5NbAvv9u7Kkj8AXiVi9UZxyYaaxQfkEu0r30A6uEdW+bMRBh9UjuZQF
hgVD0ksA3DgMUytuvClYHKMjRQyP1+jPspqVoAfzyGAQpttFM40GDGrC3JxGD8Z/
jF/LTBAsEQbmmPCi2zJvRraHDabvdPXhRisa55cB4mfVyCdyE7ByG2toLhPars2M
akymi/b5afp4PDt+HsoQ63CV9/kxLYmsIF2Y2Gu+K0cTyp1dPA2i8RIGPi4EYZRV
uX6ybyCnX4uBbazorDuwV2PcD13RVApEkbDVznFlEOy81D5gdb1LwyDB/0/ylWOt
nBi2oK+lihLuac5I2xHFYLYPHev/gS0afvu+nLPnuoNxE1OEtc1DNuY61H4L3Tx0
6wB6qBbQuYbZ5nN4sB1DeNMhHWDlphxlhJ7VkI36OWj/ouuQiHuXWzZmHMIRtHLC
YVN0c6n9iMFZX56vvlIwbru1IirhuenQXKCR3uGl5COqbPGWHD5HxsBX+KmQZDrV
d5nZTIyKAvFrdRL8RvYCmdvbXKZH8rMGYTsRy9Knn+kN4P0oYgMk18iTDSILXGpu
9Wfy7MLp+KKkgomAE67gYTmkGlb7XJxLDw4Je/koSwCMXGjbuyAzFp92V06SVmfx
8PTR4/d7asOUwcz+XvGGMwm/ztH4g3aLsOrp2aC3rRhz6qGt/L55cODmBhzpfanB
ggYbFUWLt7CXEucEseN3xHgEuRMigCVRuuZ80/vgN9JXgJua76P1emnIJmqisw6m
F09+hHY92LN0T849xZxsHszJuviAPJPnIN12Hqcrq3szcCvdRjPRhcJNKrcPSVhN
iI/314hf7RQ3rtbF+bbCt+5XnJixQ0HbaLuQGxepCXRmvzyIVFlHA5hzu3BlLGV4
CsI25pUfsbMx6EdPcyiQZ6U9FygtfftjL5CenQSLKfYC5RUx6Y5/iUlyzUgpiVyw
3VSNLwQ5PuqskEFr4EMGcBpPo2be6Jp8uW4GTVAqkbAFVhh+PJhcFqUORLPScEOT
DmjACy8oggrdu8tfFVzKNtNvSl6Xo0WpBHHF9ef85JjhjpixIyHvFjnDJf/ZH1lf
RxcGGM1r0BH9+i4Hy0J69DZ7A9FtYpz/7Zgu+ZzwwDSaZ5JJBXBibVy0765XUZ0h
Ru76qfpiYx5olKDBGCACbGv75MHKPOFXUHN6Cum9IPm2ii6yYPULJw7SkQBPD44x
HJSaQ008RvUS6diLxuFPAA//7Y4dyZ0Wi5vnyZig9T7RSUoPbXZIJiEX4pF6Z2nf
ipsGHeC5+n9XbRQBc4GJOrgsdYE5uXPRtZ1TH04M4JGJ2Gm2JJdVFHQkEaVFUmLH
5knQHsrutbYt+Y7q8rEqwvz7wJ8s/F6M9KvQCXD2vw7oqN4qAvA7KQ4mp4YSSf8z
WmzAQSKuJyuzOkwzx4UJUzVQYNxSRspRbMhg5vbIlvBpldPjr/e478OEB1eZ3bI0
hR86q8oGXONoNSFw94gOTkue1wbhK5zMOSJm3hPQvcdgQCBreC/+gWMyOC2z3OyU
Zu8+TIAyiC+sl3/0SD4II+Klqp3eoaL0Lqe4IBqpBjAzhFB0hcS5x2ATf68DVOgs
zf4r1W/4suPDqVtroiGv06u/KD5ZHIVVMNcwomaIEA7qmrKNYFOAXBzuAcfwPXW8
+8iq6mpLBY50/6ZRpfNSoSLOIgDRMFhYAu0DcbWR7QZaGgGNju15S+hE4eYHhfs0
ybrpHahkJ6ywF+WXZhjdW4CZmFAP7rjLwUeW5cA5U3N9iMMw+Nm5psmlBEOdtqMJ
RPZGoXcNKt0wqX3QwFSEpXKA9sPFhR00ceI8yWqIg9hNz+0LCCPDzOJ88llGyv3y
PSM59QgZHRRTTC2fa7PaXI0ILg4TtZFiRk/TkyLLBVHfBEok1jiyC2hrXsXPvy6w
dKLyBS5PpBffheea7zNB1wV5b5gsTSkdT5YhFHHxIJPhz8kjDxuK9TiVbrUdVePM
8T+9waNbH9UGzE+VPY/7XmNkgTrSErlzB3xsFQYkiOMf9R0NrwShe/7cNskPDOXZ
mdmIVvuaGOw5NJSHdpmpfA9ev++gfz8zFQhHHCeyvl6H6LWkMAQkaeEsPJyZEBpG
dzOJ3eY/n+16EFua/8r5sFO1+wHfpcy4TgXZKUoWGDASe/i2nq/hfqc4eK/FvasO
0vAU5ehfr+KRh0bhIflqA3o3DHKJ2Mi6BWPGV4EV5lbOms01KPZVpUmJOOInRPda
F/J2SPJL7LcRhGtGlJaBIGCKNC/QS5fdWP7XCNovVwMK/sVm3KboFMg9QR25HKqm
qcpo6U4UrsA/bG0auWx8CAu5Vfnl6u17HgBm42ZRnIRuQZzSi9Z3eGFgeEwAKB0q
mBg9wT3Yio46rCu1MysHMYE+29lJQcWwXPRslv1Q1URn13G2dcbaF5CEJfSH6Lq1
XR5LMSI0RdjI7h/A85bm9ldSKbhTJai0yJlqMPFsUO2AZAng/7+9ZXkEU49FnDnX
XtuyZPFHEN/ZcPMyU8ds//Ij4lj4DhZ50QuasQmRGq9DcIk9sB9WPEnL7LIgG/7W
xg8Dd0CgnhWhM9l+vuoxG6igFUAOYhFN5NjnrLTwyc3e80nNc2d/yHSo9OzsjadM
6NZQXjdA/PvV6UirWufY2vANA4pE48WJYc9eCgLmaO1EDa6bdR9ojfFHMdyD+1Ah
RsMQftdvBqoVGMJUgCHk57PLRrtu2sAmXj5SLgUJRxWiZzDnl8sOk+VSw7Rzjyl/
NEUEt5USGWRQmKuV+SFFIYRM8NNEcg4mB3QODZWDcagY0QKRVex3/leOk52U2kU7
Hm7JIDBTbmERfS5CHdVu/ADcPUQXkbeiH0SegqaTscUJDZAq66GS7afQALQVU8VW
DXPWYiJzEDFUloeOKlG0rCZGIBSvn4swbqqAgw6qNPb79/QuPkkZOa7Sebsxoyq3
yxLRNmrYHZYUBaiA3kr3L/+nRP5FC+d82u+jYncF5jYv4TnKWpxBHW6DJbZmMD+D
MLKRCeCo/DhiItHhXlKgpFeCo4KyApcfdZ11grw80aVcjAdrOGr7iu4jM0HDYlQX
md6XC3koRSDKYwurRXH2eh+Po1jwGA9O4tZN6YefVZ2fUpKnFov0M8cxLJIad04j
z5F0f8F07uP4k7xOvSryqLDQvVZ0bZkT379+SU4qrJ1ae7k8TXMjFNtkUjCd5Osb
U8Hz7Exlr0ucpoOGw8+x+oZw/HFmvv8yzhhdoro22K/iHKBmmJwLw7QMsOETsGLu
fUFhJTtkKkDURhmnUKsvkFzDlgLdihYUPqjzl3+3gp1kVAsJr2bplOApsVvUTHZ5
0X+7/LTncUVME7t7SsDwRCVUyt1xmauGQw4PUqolQ2V9cEt7/L7v+kXvXaTi9M9n
J+xNfuhuL3sn4thZJ6CWg9CYGLeBlu2U82nHCcwAjKi+G2vL9xT0zD+to37GWXLU
jtJzxIuukoZX21LETVwLVuSjJ+G2705QDUSEWY5XnUIvWWpGLBE3omp8jHIZdSi9
NFm0jcQ/uY9vOEEuVs+5sbMXDqHOBhS7WBOVBMKjaBYTR9Mb97FeDEQ+PCQHzT/R
L2xnbPcjRhFq37GL33ow0zmalaceF2ShUhqA0UcdL+lMEYgB7BQfhfStirFiQ9Kd
MZ29CyqkNq1PDALjOtjC1FitQvVA4548rLX6o+22alaCXPlf4zGmBPyaQvg4zsqC
VColCCd1hAEusK5i6nbp+EeVBMeYAA4Y8V8iZPfc/DnqosPbPSRsTxdXdelnVC1P
5uC1dp0JvR5peNHhQzPNGenCmiBrSAzSU4O/P4tPp7HrK6gQli60LprGzUl9e5dw
CtG5Y3IbdgcZNVfDsTiOBtd9Ggzp9O/t78vVc0hr7smQmr83nYunFPQcZLu/eC8T
iPLTcpcG0K5duokdw8FixZ+3ZdE019YRT4G0/ShayNrfoxcVWF5t6DObYJJkPE0M
vrRe8LxnssGD/3x2M82amOyZc3dh6MbgLoYiiR24XeyaKH1gQhSp8a+f77IQvB1h
7LaF/t10bCexWP7+PsYiCLA6lb4rDXU34qIPVXGmpabRYuOWw6NWCoTzd4snNOiS
Q6HpsSo+SSbQSJ35QZ3EC7LypEEbODfr56zPju8ywN+pv2dF4d2vCSCNU+RMOLJJ
i0mpYwkmI8kB+ZFuW5ScQ2n56Spzt+w9kAnOrDslGJbs1M+a6ExC9lihlTKXQTRl
P1CvRGxVqwThL229qWBIXvtROue2K9tIe0XuGcrpCKmlrPXf5ea6NtiImPk+9mYk
9F6BcISpj3iajtj6LrYRB3smiOCIiQ5+E17TzX1iqzpL0XiN+4qpq5HmDNAyRs9D
6fm5oM1ifTGCEadH7bo+IB/TuADRMNjmXgsDu6fx1BYZIOgbchTKcBTjf/BwZ/UF
ojAnWd6WUUU19RV9EhasfPzBlQ6fGmgWRGvQdsbrOyoj3NVbUKSu0P53V05jBxg9
4BJQ+omIj67P3G6iwW5LY29miej3aSSZU8wOHEeufrarSftuBf+KNTLeqvgPsPqy
jfls7xDznFJD6oUOu/bnLrdre6YYqpU/x4qjur3yYKQIx57jd7AoIAaJJQXuv30L
oQqu+MMa/knd8zC3CXH94dbPH+i6HbW4wtoHOW3Buers6S7mR9tTorRa0LEkW4iA
PQicl6Ox6rujzBR9H0xbjyNRm9y3+oisc/vxgiaA7w1In+JdYfK+/NAuxodwKw6m
+DLeqYSJWInTvPUYTnwTKc2MARk9y1pApCxDo2czW7fXzcvpRt2ZSV+2UhnuxhyI
Bm5Uq+7IezcCEk6nM6UJHyYUoeY8Vb0T/LRGCXBjyGWzBjPd3Xk2JKLHBqfUC9FP
v5VUEyJf11Lytl5dx7opNUbgis1vO+3E+kTrZfueDkg1kUxVR5mDKsaZnIblgUFK
pqOZ5FimUBjO+3W1qcBGTXKON3Fmk9QGdyZxWEVSeJGcapbJ9ilTjzgBTLku3/wO
hTVZgdDw6ZTw0MSx5Qf2QtXMdTpdHUhEIo8n5NDNEAPtbkVRWF6vB2J8vW7mo4MI
9YimpXYZNdyIzj8sxJfihag1ZMPav5a+hA/jax6IajcF5CRmVTLfm95paQbvvakc
zqoS38c6TP4f2+8yx+hGKR7k12iNbBJP8GmPBZwlLtlg+DviDtYTMwwNOsfUL8BW
D2mp2IWgiDrIf76vARViwOrvk9htC22R7e2MxuL65y85AmhJpuJeuOY3xyzt8lXu
Eyp3uH2EIrjIkA9nAnTfWSswbRohCEC3WRyDISwPbeGruGY+wuF06geNgcFbURMN
5XLtSsyLN2AsdYPcOEjZHE3XK0lKp3hpYIYqspXq3Ys5sUk3hiBlQc1guchlnekP
aYl4Na2nrd614XWYZ5TuwgGeT3xitKryrzi7H/GdNj+5RpSlb2m0frKV4WG2NqYX
NOKi1/RTRJAxGfLrnmGtAejNhudrJN96Eu6KpKFNwlEmIf1cvV0qwup6Aq1fiIfF
pZBuiiyXzk7e0IA7UaBco3m96PUTGGJRbRGFLUjpxpgH8djMD7HzCwVO5Cu/Shs4
WMjac5/eracoOu+haf9SqPOyM6M3I9jInF4an13ExzNkpxrBXuSudipzsMA0MHZV
esd4btrl1Rp17tapdN7Uorn/1YrjlHlOt/CJX3xDW3TV0uAH07V1+O3Nk+xBnH8B
XYFvNTq6oDxlP/frF4v+2Hv086Qa7/3W61Qx2LZ2NGNAh5v8KWwsTEo4h23eBTI+
b+42KRlQZf0M+FjQwSWqZfddoTO9ClNrY+4IK1FV2Nb3Yge+AX+GARgQvXui/VlO
WkQhEK8l4i0u1SIIS1e76I7VfiKl+a0VjH0TLMqKtEqYyDUSvcooZoa38TITuGE7
vbpv8K5R3zEDdqvYXgbfU6+qQN2rCL20AdYSNjLh73lGrl5cWdCxXI6pSCyJsIyC
VvvmnSRAUiV0Hl1KzkgnX/3cEkEHjiLIwoGjgIJlnQxGo2mnwv/+0ADeiI50pfBF
NBrdxD5vF11CZwWFvHaDWGc+0VwCD1QDss78i4WHBmbmTbhUMJwvf/FYXUVW8Iev
T0bBVVwlMSIeazCWlCheyPxZSXvJr2nSOjF6cRhps4Eh1F88eCffEpJ2lqSJIjIO
Q9/oGu6F49dUZ5omFLWd5q2WK+HsfoOAARrCcbM6+h6smZJ4iZ6GqigQWhUQ7fRp
nZRx7kHrsdRrbBKN3mBLc/3fYiwKx/itkeLD0P69cXM9euglAk9MqZt3kGdHSaDb
qzrQX892eteHoiC1I0qOfN0en/yqeInHLmBgAVXf3eg+FbbD5GZEE0ACGrxR7105
tmLsW2xVQrV54vWi1QSePCFewU3y6RQzmtrC/A3aX1/hjqUD6qm2ZF213dtdWEMl
1dHxc71xj9GTrlrYXp7eFpEzs93BUSJ9zxP2Ays/WVcQDnrMMsD/URmjCohSqwiO
VhQ8ptQZ6mTWcUyKrrLNcXdzHV0k5MPwLtTbPJ7OIE+vbcP050K3ePEpxpsfiRt1
M5XwbA+S4J/lEOkwm6rWLPNI1nVibaGQ4XZE9n1V3ill1AckzwKm34F7ZY205UqL
TTE3iCkjw1wOG5NsWwfEm0qTMf/OJqd76MAOD6ZkMBalfBWn+x9LcOCRaEHdhX3X
wg1yEWI/8VTeACVj1zWIynZzgwq8w5YozZk9BS2yBe9vK2vxd2qbvH4kq2K9kjXH
2yon26qgsnK0g5Sea9cYdzI5xOfUMsUqmwVTvgkB7SC0jVI0H4UQnrPIq2h/jTwW
Tr0XXQsNewmZ88+ZXP9S6y9y1yDQke4v7hOx3ZbYnjnGFu+sQbASIpBqIYkMkEZB
Z62GKIqEq6aDiuaQxh3FJn32mcJB94HAJ19Xu6TF4qz9QF+juHQXpvOIkhwRwCqq
QRgNHiZS08t/7S5NOoDrvh9CKu9mqm/W/w4S1OiB8Fdh9cOW8V96b+bXUK61Zkxp
FmNgqVFpSZ1xo3OR2lO+jbVnRwOKnJY7Jx/gsTEnHwUoB1ov6g7cOyckQs0knvHm
DGaMimUYj5TPGlvi2laiHGIfWHWOCgErvIG33lmqqlRW6G9H0McZ8hPTo89huScI
x38v/RVsHWUD6p5spmcF0CDJqK5rNjllgT4eCqa+s76uBxmhEMbUBBIaqQwlDdWB
AaqPJ19IT58E1KUziUWnfqojvwT6mG5mQ/5bFBMj65LZuwQWQWOTePM8aN88s49f
d52fYF7VZSSYr0OIZkAQS4K1iOjwyKEkIwAa7Ozc1/8G7hn2FcpLY8Zt4DHt5o8x
2uC+ETAudfwkF3jL2vpnOM1W9XvDqEdFg+ldv4KiXE90gRiuSgAVJPXmdeJJljIA
XVcJbsJcoMTOoJSCfteKPesVotd/q5gu4mG//v5iX1TAShw7i01CY+GDJlGywlC+
jQ8Hz30JCRfhop0jWWNp4G/cyeT/Hy4ThdLU2WtpsUR7ZsZD7kBetWzeWSrtJsVi
R7LvvBSBsNbTgWt5n24NN0R5igLG1MCpksj9gdTie14x1mqKeK4rKR5kNVvkToNF
breh6bK40P+DMSNmjNX4tD0kUJb511yFVDIn5xMCr2pTTsmJMaSR2gV3T48HBZQh
3UEH0c1rA4/CLVG8mWGTh4IbBFn15gLqXGRgevSDwNVxEPHShV5N/O4Q7eT09+vZ
vi0pivlTE2gOZGtS5WmP09PGTqpj2wRoEh18Cp0fGEoaxbIV5jVnMHPvyGP8bYRh
aTmbCQ/89vDBi6vi48p3ZLdPavDVcB4Mhx4u2F7YvNp9j0z38coJcK7widK+E5rb
0OVJRF9KzMkeZPy5Rn/uKt5jFAskGOZKq+ODRZ9rkYoHA3FXTBV7cQGZtgHgOIrs
MtEIXw37EFP+qN897xBizlFlBe3vmWM6p6E9bBcNBdf+f1HWNXz4voTV4K7uIHQ1
+pJck5ym9eTl0bfFZrU6RzwegHMOjmyeA0wWoG3TJFyB5CkkknImN2B9zM9WoPsn
jVFGtVGjIwgCPnDUQoNq+xmc0+3OnqxsoJslFrzhxXCQDau2FO+fUftVL81wGDSy
sEyoWYOEca9mLmbUeQ1U2/BrXjPlrc47Xyi0zxdpECZCEWWu1IthtXAZQ9gab1r8
6+KqQLBfGOdLOhfGAMy7qar1gPJfXnoP3XN9XgpmtzBnXKxGiHcwsZyy/Nej/0hL
WQVZmsUYf9zvUhRE4Z/0bnaGsJr6GQrGFqQsahqsA18cC8VkzERrfi1C7r75tlS/
xZmFAtyweytVCsaUmFmpMYS7Bm495YE9K69pJM3cGyXqwCYH+owJIuyHtlUVF8yT
ybPsxTil7FUZhSMKcYnN6sDKAaKUMcnh7MvMr3yI3Gy55GlVIpzZoIg9NzqWL7hc
VZFczrwApHbIO2bPMJhAsjtSKY3kxBDynsgYCbmcN2/w3hzScRAe4WD9yDeo1RGk
rSznDmtECSktzr5nSJYK2XBfKqI9W4r6RDMvxFYJBa9fAv5P0EAFWdcd3WtCWix1
XWzxXBDtOgyaOtgwUTr73vPUHOm5LNph8QFzYmNSK5DFRIpuHK1sXy2al9vlCYOT
U6KIFi3UUME5ACxVYbQtQf1XccWte91vqmNiuicMTL4lrgq1OsHE3uSS/HDwHPXg
vKxMOW16XeOnsTp7ABXMq3uA5+wTBlIimmvkBSJVSE8lchnFe1+5UaUym5J4Gjwz
0EyLS1S1q8ndqGLEnjpo8LFuWyGqLUFEIBfdm+vbLSQ53O+8r1naK3cUtHF9D70M
XkGbgF3ruuOEx1ui7m8WbkwwG61/IS3lcofaT9cdF8tEvcH+O26Wu36QCcwJ/KbF
Zaj9abE4ibbEMgbeiwsafS6ePtpToQJeh9fQuu43c5h8aUb0po9E0VnVMGn+dOWR
oG58gOI5i5lFYYbkojSRTQCk2WyA4hKfNceGRukUwsUctJaDQ4HIQHrQrBV5pmqX
oqpdig5GkUSIpTLWw6Dcvpgy2wyjFWNaS1nzfCBx8ouX+W6/NKnLxwqzXV/Tb6I0
PzhOGiJ8lZ7ADjxVOnVWrTaAMQUVjrwBmKmzG0NgcbrwgKT1zBKMCT6GCKBnWBMH
jpEflS5Bc35q4JXQcF2aKi7ml2Ya66y54Dr/aTWccUUBJOQh1mtsFy23/6gjgYHS
ERga7QpMAhJ28mx2S5DK1SgpfgcwLO6mUsdhuJrAXzdFi3qZtYc1X9LPM5K933Nw
ij6Y76M1KpqDXUkItX1YNhHYtpAVMTFxdZp8AelfqlmM5W/RDzqQCAx9MhVwYS0o
Vh3If/A1iehRgjfPq+029btZn+KhqNsr1+wJPDDs/GEjcNAZeb58o0z/AdKSjj95
YCz3SrYO+MxCIOuHFKjJ5QMi6FTGTG/aquBU8f1WhoKVejmTbj4ZsWXgnlp8Fdnl
qPk3+GfLP7isd1sq/f334xS3AhliZuJVAVc5nWsh7A7+shk8prIuHJfjx8HU32NJ
VJq96oUiJ16fYvYR0rqTiET3TavEnuq/SR7FA79erNynenPwoBorbyIFutKs9YAu
AZcaSvtX7hDzAg5hAwAnHo4mLe5ntKSt/nXH5w2OKCnSB3zvVGhckkguk6983rhO
oSH415FxdzClPDRLIq0oZdVDZo9TwIHIcZ0psn9pKjFVMz94ZmwluZFlxp6+X2NL
WTbDw4AGyXxZPEJOlblqcfWQ8jTVD2A2c2zbt/V/YBk+2FtUOJdxOzGJzXCGHalH
K2aMHgtIChPRxadrHpazCD17YpcVk7aCD77pOvs7SWVD+iKmNLvjlGHMJ+hVZ3Du
TERi98zJ0ycAzYd6KsHKvQrLjrX34KEOjKWREtzFHvH+PpvI+I+v5dCHyaais59V
kEdBWRNlg3hfbEVHLZ6vuSGRfVAwXhxjUk4ijzq1UUstLdclNwlCu8yw4t9VCW11
/br7p84h05Dzgvv23tKpSw/TPKXNsc+l3MVh/cc8kw8nkJPm7OGrpB+wOqlVRI70
MqZgIuyRC3Gdqc/3/CF1M/usPAi357VzI5UqoCYg2RvI1REjLKSiM72bAq6O9sQc
0HBwRokDveVdfNyqDUoYXBywqUTqN9ZlBjY8Rs98XXJZ+lGnp3rzPQtS3NKwlgWA
4d8lGW04GaEi4ylVk3OPmFU9JFZr94tpxWfZoIoDH5lRFaMAtbM+SXIKKiJfuU6J
NquamorXcgIR2leq/zeSerEOEvOTLDbVOK9TFpS7ojZKR7Aysapsc+3oWcrgPave
6Fnrl5nPxBXhmidBOM/3NcBNZohytgFk32iAS9+R/HGgHH/Uwi+2XfVv4jzyt8Z1
WY0mgCdQbro1Z1ONKgZuoVBT0JxKdo2bQ1iiBBxN8afH80YO/eyChz6U4hq7iswq
2KPCEQ79se+BGRGWQEG+pFagg6w2a/TuJLbB5y0jMvhmwPG/8gMNdIrzfvMRq+oV
bNsp1Jd52qgNGrzG1yPtS1krdnOOgvOByE8hLioUgyR2xeEfZONYTn+BULBgrcZ2
e79z+DwcJSFz4m6Rc6A2SIPCLHnPgnBEp4J+Uf9JDCQnMFWm7ZbBcEwaWmoNkC4O
MattyXIo6+JplfeFTLoj4/lS13XL5Tmgm4YwKoK1lI4nsiAmb9XiyV2X8sinXCq0
SUxuzaaME2y1jp/bXryUvxvOZcpFJ1y8kYHmHdnskpygH4UnayzBViSZtEOsh9YU
qG4EIGid3EfH11KL0FqLiPsD+w/i7zUpbLdhX/sUBEe29Gtvp8P/HpxbD28Bx64k
LCRjGrQpziNf/B7jbWTA/YgAWNMG8C5mzjezmHsII7tPFLWqy6/mSqeN63VV2geY
0Ms+DcHPv8p0Q9DV7UmOg5U1exD4yDkhGBACoO3fu0IyngmBzEfRaNtva7a93QZz
F3jF9Tk9aOLGibFs4XSjhA/bzKb276LUI+I1qwkjwwLtV3hgOPT4Y0Jg7LS+3m3z
2XxolkY/Hl2EgAhhDjpcLjwCkOtOECK/ttzWoN6b9ACWT2whx9oyowpdfiNhUXWd
l8Cbt8XVAau/4Gbw2Zhi7vg/adO/3oPjLh7RWIYZkN1p2qS06hfn20OwDgkQxX+g
cdQMHd3MDGMYgXxMdUoztd5VtSaHHPU91YaW6S30X7gIjC0HVLUEksn7FkyXnxWw
ArPz5mQxlazO1qMNKyCAuL/EOE0PB00jPs2xkNMz2k0b6lHwnQGOu/1/s4fnM27b
KZ7cmYY1MT5AHdVHt+f2oN/iZBc6bAzPs7BwQLCGrp14W5EH2+YfMYBHlVkub/Qk
mair33/77j884UY0A8/kcq2XO+V/L5ojOevynTOxRbpAx802IJ7R2VtLmPe+yVzr
7GlHD0XBqhrjRyfTsnHTqnYrH/6aR/QvaIbEbtynwyqXzdHDQGY0jDcb7B/4QJ/H
SDQN6SVGUbYoEwX4Z57mcgagUd3EZnl2B4wyWbCY9vvdZL+UbAaqi4ErSti6hkDI
Vm+B5iEx6lTqPJ5LHt6BnnArCMBS2uXepMUvsTkL+/Ry72yN4WRMo1tRiaX8vIh4
jXS3jNwNijqlEBUgYxcJLlkcTS/mxBsxNRB3nf9lQecgu7dhXJ2pH42jc8y03bpg
pYu5AgPy+F6gXwCdXb4y4TUsU3zk/rnJotqj/ODiHNysPGhcmjY7/LHU5735DehU
GTrs3QCuR8WNOromJVYUfTGBgumPH2OtUZDvGS/nVX/BDOwp+ot6CuSzUXNk7G/W
5+v9xtbQTKPpZDCvTLn3a1dstmdzuxrZM/ZRExiIk5sKTnAjKuq3aW14igmVD5N7
4oRRsD1+kKAYDnk16brpnigoVZtbO+LM8zZ3ypMNTd93TgFbD2kxmDFDhZDyiTzL
SzlPYebx5Ca4LlQaiq5t91BqPUE1svTxuu5FMMz+9x+6CRyOoe2pNF1T+ZWjaPTF
RcP5RCWBHJ1XuEwUwWyEteYxwA30dqCgjESgX7aEAQyIufyqhItRzMw0K2+fVY6F
/MTrIGdEqTKVSG6gn0eSFHjMWdKalDHeJ7VRDaN3b2myjAU18mYQTvvXFbT7JKGd
QPnbw7DX+nm0UDTp+ZScJ/7KnO8NYmQ/O+Uf0xeJMTa+D5OqVzVrkb3cV8Mm3ONF
gnpVWuJajCoeNe+eYFL8Y+us1y7JCEYtIesBU0apuDx88EpNzfQs7Rl7sNfUBeOs
VwL+siC9kCZh1vzG10KptmCwsjGD4pQ78jQ2W/0Ms5wKTlPgcgGXDW90Xh379PZL
O0ythkbHNMhmpMAJv5dJAz+XUXR6X9ckPp/L0E4wrNMZhA7CK3oEGmgo0AOxFXtb
6hpotXKBJQNkmtr8i/rXDm1EYHLEufnCWKlHldUJf4MAR+2SUOI7tVAuYbEESpZQ
AvXNfC6ytrwfo3Hd5BQ9XatkNYA/1hC8eRHNK5Ydnc8dvIi3qT4glxftURxTqjkl
RWgbIkqw5DwG878u9PCMopXvVMODbZt/NecB4RxWmQrr9KU3r5DOblCFxQR6WBMP
ufTwVPCG7lXduKrUHogwBQP2ktht+4VwiYb3ykhq7ytYm7J7rjNpjNFjxP2m/Mue
mpYgqETnRxQ1n0ejYqvvsnz6TSgKx4e7DoA+0uKa3TfIMyT8OcwZxuAJjHGFOW+L
Uw/zdTzhNQ2ndx6Bky8FriBGQUm+w+Rfn8CQ6Pt3a8TKbpHpxNCf0b0WXVe3ID9W
EvSb1VzppEApJpvkVpobxGym5obsRhrVfC+Ct0D0k0jdA0xA2ZghnT4kkAT4a5LL
UxpOzYlUHbYOOv1JXv2jGN5osQSrOW3ibAg/6Ih3yr/tjDvH893iyjATnh/dRA0v
eX+r45I3wG35zf9cwb8hMViZ+DzgJxh4xU9dVLVdG3QBZ872ByDXZa9teibiFS5Y
mvlKsdk7+4lQ0YKwXbZwZQNeHjLXMu2ZO6fWMW95FYmENEIGS14d+JRVTgnEJsbX
ir7pNuvJgSiVuxpXhgr9rbBukJOoqpNJ+DWjQSAzMONkBOMn2xTd6j4rplmL+EnZ
LVQ4h7Zm9PTfVqaqq1NuTKjHYjwFaY5FkAtf6d08DTrcAbgaexMujGSaiFjvWDKV
+oYM4eM30QJud+EwJHGjqjcwRHj1TuggphxtgRN92g7f1h2nIfhw0qC0/hZtI4dY
aQNBDEcufIv4gvw6q0au0ZAiwGVZYBfTg36YsEB6L8S58gEC7LrLBZp2KK1xL3MX
lTf1Pr9sGGhFcFmGjf0uq7m9ny/1ll+9/ujtw8v8+ddPtUGRE/PtuNUrpmYrfpoX
5gJ63SAIt1ZryqmaRzZ2DfgPolVPugNpkJWmKuhcq/jZNzWEiwQgQYNexS1sSQoJ
uS2/Nn5WfPLKpKG/0Im81XiP1g5uZ4LswpdK2P29FidtCvelaHn6QDV5wnXCH2hT
bQBDszBqAnH/QM8awIshcg8yMpwk/fVZckYFwqrtpcJu0aoIaOG7l4qfOIsAan+p
IohYFi14G2cHIqMZkwwca1yhilDAF47sAIIa3PIIk9N+QwVNNKILMXsxS48TjY4S
iQ11PY3H9Lg6kLtGwxS26r4qv7xBjR+3wa2H1F+AB8m0aXq5zgZRyUA7BU4os57M
8wcEgk9TfvOaAnZwOR5aYllb11bq0kKdaGHUEahaZEuzxdS6Xfz2ANL7PgPqjizU
jLN7sVgJj4d7RygGzvpAoTvzBv/o+k8DAO20GZ8AIGCtryOrdstt2Ix0qwEnXKQ+
MRGTqx8V5dwn88ti5Nf7AywR4SeEuqGSMsgiEFJOEWmI8PURzKG8EcYbIO9xD0Hn
L/uI7LjjQjkYUwfsdhDd4HHm3Xw/zIbGeompmWpHpr01cTz4Asaooes7VYhGxVD2
7zktBtUa4y9Xm0N3Z4TGVPRwvVk7+B9DRAnq1TV80q5ElZrK1V1PO2jWGiVQWzdf
TFI5BgrKTBaB4EOATQDg7OHxy3AMPN78qznPna54RsTMOGn3efHBg2cCnN1wiooF
fQKWbM6+aQHTTog0qSCTYkVzQHagUZoK2gWlos+RHsF8nVaTY6gNefRWiV120GP7
H6cXN600mHocLr/qNZTKtkpeJqTcpynPJ33R1GpOOCpIUdehwqzYFYVuW5BTDUSW
Xm1AhRHjhH78l8nXQkBU3VA5J8yyn0coXJjv7UZxMAqJf6Lg6TC6GIX5spcBYWR6
CMu1f5Cy+lVyAAaG+sJP6aEzwIWYH5imZCN1ZcaFN09A4OPScNUGZtaLokdRlD8k
qcP1gz0dbB/6332P90DzUXtgxsljOWth0zua5UF/eV0vkAWKKdCwsj5C3kIrGEx+
ehk+ev2QYwNFD6fz4/D9iUn5ZRb8VYJvX+Sm/vQ4AkSII7wrwTN9JMDf7Qv1A7EQ
yYZNLO5Y7Y53eMj1+zvLAxqIFRzjtH53HPH+p5QEFT87GlmmSiDRYyDWpJgFnTKT
YDX4sXihLb5Ll2TObDXlVRYndIRNDm3d1FZxcrGsN3JOfhhSYBnE9vCpboL73uuX
SbJ2OagrCDU7p+jcdwaxEw2DNIPEznTczagFPDXHe8xKHlih3wdoke+e1Pt7hyCo
tIuavUfmMsQq/hw/+1dgc7D4xdnTFYk2OycOq7pkR1NbFFA2ykj+o4CFx30EuDHC
Hp0n2bp9uB1FQWDDY+yZKmwjD2eMmFfXFlhHKNcUmgdOaKVhwMKi4oKhgdS4i5Jr
k5E+Nqr16eU6IEAv9vYto7VtEhz/ODb6sofp0WjFQI1mIJhNn634aq/aoMg+nBxk
PSHDfXxuihdw6Nzcqb+g5g/LakKZmsWkMd0oX7dpuxHyVg6e0MTeJoX9s+IMHn4l
FWMzFLqtz2EJ4R0HHDh+ffT5EuXJkVDeV0LB5DCsSjlb52eCNyQOa4wTBayZ4gZ0
qIPE5VAdZ0zVV7bA9VlSaCY4HZsNJTcjnKNPnOtdu+ynm7nDrpjiSBjYNu+3uGdq
xHNk0lB92acV/uSTRlqQ3x1osx8S27h9FNq5yWi/XsRFUaopH9TcuEhqmW6zTrXx
m879hg7SQjplJT+vB7wse+uUm7TlrjOXbQDrygolGv2qpT7TXt/Caytx66UXaNuN
kBQcOz7Z1/1CP7rLm7VRItfPK3iU4mIpuKXTBmAqy2+W0wNqY09VFq/jRmP9q8am
0ht/w9YpvgPySKFxBMVDTv0Qtgz9wjDWR/L94phI1Le5vbt2KjtNiE/PjfGumU48
4lheg57gzuZpKXDzLWTO0zZl7Bhq/f9b9OxrvinpwEoGzn8ZHXqB+7PWks/tLJqH
KZlNinbmpNeUGLszBxIrzZ5WY0fu4yyc1OLMxZ0VTRW6mgkTBYWhIdCwF3KSYCf/
k8VRy0ddC72QzmRcrKG1haygadPGUQKNSO+k5bFmlaOOMdpWrj0xOJJZw4iorpph
sx4KhD5nZBvded7U0Wa0DIzKYk1bYkSMvsqW1fFILwraMJQU/rTGHVPs2RebS2D5
pzoVmbySGp2vDAiOavgLY3BlcH7t5I4Djtve1oAxVDhZQsJMxKk4MlQcc22Uhk/d
tU+1SpbNFyb+nD8V9n9K8nB+0ZmpA0/9SdJv44936ecsRVcnoD4Qe2MXmVezrAN9
ETeSx08pT/0tjoclQBFq/qgDJOFaq84rpBJ896d8gz4RAx91HFDl+kAJ/IfD6/0O
533wZpV5GLrIlC/csqH2mmHeOnsLKMYK4JgUFtV3IHZb9Jd9XM3rNfZAhu2bvqdw
I1ZWseZo5ntGkJ0fw0kI3e4izw3nNO/VRMK61Ijb5fsuSSuex+Jt9P2hxRnxLOl7
daBAu9TyurTNnczOxXwGUcjRxAMm6nq/h5NHGbTf4zzQ1le/MqgmaASr4mQSZ5mv
9DZyTLqnFIVWSAhR53TxGIOuI0IgO0a1XkiphVINi8P1Vcxl4s1n3nXz5WxIwW8u
ZVqxvxhQdD74Weov8D981yUzS7rA5Tq58k+xXKLp4A5d95NOAEoZow4ZmnxovNEB
kp0Brpzx16ibJTYfe66ToqpV/t80PA8gdE+CJW7V2oh8KWIoTpCbwaIktlp66BbP
79/fTbJpzqmXEPzKQ2LCZ43WRixDLG5mzeFCSdY2z7DquhRkq/njtF5RhL1a1vxJ
wv3Dqz+RSaJuMV1JArsaNYa/orCuLsxTIy9bdM8D3Y1WKnO1rX+ErR/+W296GuTJ
UO1GWPvoEpETSJY1f0sgRieEtQ3DccQ5im3t9UmePO95TeVu96jLo1TUuzr21pO4
DDXv8bY9O/gD685HKofDVTNE4l7LemIqu90EwltFnmiwsPvZysyUVcY3zS1gGJsE
aOR96S6OXp0ymUwtSNWKwXMN0mscqmWU8tRlXJq8Hmj364ZLkUNobwY6kGRtvsjT
D9MwXd1MMyEUgNd9JVCyjDgx2wK1r8gjcg1a6qZKcRIS4sVY5zVN3vekccqowvpU
rhZIsWhmyk1VXWZeAhJjvoCG3UjNjKlf2o/XxGhfvuYORNCkcNihkHi4hjn73vch
OvMWQN55lInvxmMTLkkhnpCVW6wINxYT+BsgfWehKBcodAYWf+OI1dxSAgxozX8O
SAdzDJh7pip7JviMPF+5kT+RWA5vYpUolYg232cg5/YsOcz/LBXk08d9k/mQ2iYq
Sysls8Ilsi6SNVSPpLnTIYhyyExctdflmou9RI9e3KAf9PFkVA8gpKWOlvluVShy
BoOJrO4WgLp6/Mh9ijz7rUuPj4nN5jE2Sg1R5cTspLqhJQl9dPa8IPHL9MJWAb2o
Yhl6ve8CFTqmL8fpQSi/BL6/Z9WM+NkQjehxwT/A1eEjneVlr3n7dB9KnWgu1bZ9
wXUr72FJeU0v9PSKGxNJtwpzjneObFkZL1OihWNJAWvqNfG8SuJQjcy+MV+RlYDK
BQhlJDrh2nMxru3rMYzCzRcjxVVQFUWT4khBBuCg98UaBTo3ggDlNpZfi2aFbdYY
HL3/XjMs2Q75rVPrrIC3wADvW0KXaEori+6zmTIWQbOKy+iPKMFpMTX3tydgkppF
I8rsQR0yU24n+XZVBMY+ABF13lcZ1wui9pGdA6kHkFQRkE99yCcZrW9hx7w1jI/2
mpTbpmTP/fauOdkh3LX0wGaM3EMSX7wyk/ySXIb4c/As6mmb4MZDC14x4wt4qdcC
KaMe4UgHQU/MpHhsIvpDQuwVCjHiPFfBeCfWn2nQh6K7mAaLpHK6EVyd2KWiVKek
soWpDfgVUuVAE/Sq3nfgJVcIsFfjIveFj5UrJlfeTXzynm958/6Zy9hTDIbXRkHm
tmHtSb8DIQIwHMhtPBFH9ImBGT57ZDvHWZPtj99dH9G/voXDdACY/ktIz8FGKS2I
pcarpL5X+8uB+ZuDcxE/vDl+o4rgnPW0phobC0+iRAu6BQMfQl4yszrnOkeUJNpY
/Lo3B62W/uNQW4Ih8qdqSm2bNm0zgL6WIJm/hhelD9Ul6S1vSLLSLFZzGp9Extaw
ChZTlkZhVHnRxdmc/6ZvO1Ft+I7pTShlqkOtnoJOuvxoOecErwdG0vkMuXiSCYp+
fSPU695Qa+w8eqp44dugw+R0/g+rjO9ZhMOaAiyC5Tlf+QCYxEKWs4tE/l5Mkfet
Tq5rK5XZ7Eqi/xoyt3JmohUuV9kchfwt1jk3WuRlBDXcvT8YOxilxx6RwlqNnaNt
wpJC6guDULBK2Tod75ZVdegHoqqyKF6+zGNCKOQis20R48NgeunmkBfjfdqCePqS
5HPr1T+aVCzkXGl54gz300MftrHyDIh9v+BMoiBUn8F/DpfAZiSU/2w+4GsaM+UN
dsc9YpEH/0uPqCXeu2QyTcKUuJqWcfhoM410eiOHpj9BJ2dP6nL4596RItEFqF/q
oaO2xiXv2FWVvwzPP7BtWw9kcdaRbTaLI+5LXZKSWC6JrumYSpBPTB0TGHQyDceD
KHegsv9GIHhf5NAxgiAISAWr/b3fbd/GPlybS+CVNfQUL5grIdAV+mn9TclPh/G/
6zi4KlDWohTw78Ruv/xHjNI/9A94oXYg0P+XJenBcKnMup9ieBYzgEMswHYpUL+P
EigAZcoi+0gCAdRXNR3PF3PLgzjTyk3D2YPymFd7vF89nb3I/IyDCfTuJ167F27l
1KkVX+cYcDcq/4INwFZuOzhvKOIShAsX0EovICKBMMjMzOUh2ETvp/zqJHG1ts3j
ImRaJ6oK9KrL3DSV5tRwf5BcZlvIkL2zd+m33REhEkKCozL5slUFFwVKjweGEl0n
Rs96X9KZXYknMyho5ZBYQrR9IGyvGVJ6UKtwK59E0ZrfKDt4ff3RqU+EGVqSr5lU
kIeyzequafMMM/Uvw5OHS6bNQ1N3+iVfrOxptNmkUYWjy//QUpzhzFBpevIpp3Pe
eUqXBXVCAHy0q+9HMuvfsfgOrKGYZOOfu1io0YWavEgFBPrKAbiHgTY7ELhcvVeo
sSEm0J/a7rk9A/mBWoPouCjKejaR1aVxFieY1QX+pFgkTfoDWJb50pwWHcsz9v18
oY7RK+yhBn/7YjwnjxCXIOSELHNZnuy/dr/H7HFtJqAzOJ31QsjlRJLavZTQwfwa
Kt19Bv1aOzqT/mpWiqGGbFvtIvjDnbuV/349AbTFQHvwVYkDRcEWmv3STMiUw94O
kLqFKZvCKb07KD3qc83xe+UgvBLgSlq42R2PI8zI7CoHskt6O4jfZKF+gka6kNDP
HjKq4WLMt04oAKfN6P3+1UIJvUmPXTV6kpUccZKmf+TpMRZxfji405YSMTeKcSY6
odllm5rJYmOrDmvzJqr9sJyczmcgKyL78FTSVWBdsdBPo0Y/V95EK01KzEgPNgAB
4f/LQiL6lF1Dufh0gcjxk7Mhhyt7Zrg7iRrUJHMmfg1EBUJVzynpPjFZGe195VRl
jZUX9P5zY13UICv1Vy/QsOG8XahDPAu9WH2atniY4K5urutEkXBPyKZC5BYfusLX
r4YECS5DJqDqxGTj9P9Cl8NycD4tX0De8ABQd7IMw9K3no2GZq4AwjEQ3hUV6NQg
f38xLK0Jwyht1qXwlda95TO3aX147ykK/Fo5wdrpf2Zh7Sc1GA8rmlIKgHmsxY+0
Gae84ibCtkAhPsz1LmeQIclAyY8BX3Ei2BvTZShdInlMOQoZPePfBXkdIYgp7jfg
2EZh9WZ0M1XSMJpx6PdWAH56VXvmp0QbDGsyDdBDZDblxUstMTJyfQ47zMK7PVCB
cr5sVN3AqQVShR0eHv++0xKWekZYlLeF8VpgcRnv0NMoHHK9R/2VfZyus1naKqcV
C3DP57IW1iB4jb1mDYrips/ikNCGluw0EcSgLEpqTQbVMSHMHMLrviPkcXQhMn++
Rfsz0YHnVP02HPcQirt5BE1cwahRn5KBrZb4PnVrG5WC+4ovjJq1Cuwl3Nx6D5tE
AtmB8NFPOj5bMFlOojOZ4PFlRYAxb39IQ6bBU32cxoINfCMlhO0v3j+6Gu6JJ5IT
7oQzFPimTUmAGX9C73lh8zUAijgkfpYQJKdEBGjgM2zXripJMcn6wbkH3BMzv1Ru
N9QkSdqpIniqfM1YPQzQ/U96HpCXLsiO492Nm2EzxFIaX6yAnH/fFCuKSGmXr7mx
EeNNfDhGVNGIN87Bo8z9/ikBcWGQoRCbNgKXS9O/4QjlKf5f+y1kLE8dbwWnMv7/
1MnBxG0AmUrurP+/gOR8juZ3KvZKZ7mpob8wmTlBdLuh4wkwCtHvoSR+9tjTflG9
T7cUJt7bcxerZKWGhKd++RwlTezo/G/EUlW/heATxI2nRJbbfty7BXjESJbC10It
c6rpIc2gzgnjrc5vM+/tz5Ta0AZR7kawhl88uqtKeRpID0tLbqRzgI14z2F8vdlJ
+Vc+6GtHPNKpTxaqP0U8wYgLyyIiqxW8v7NkgXfbl/E2bDZGqNkfJXv/5NVJmkjg
rn1WgyaNcQGVDP8+zyS2FHUvZZUjGtkUdQadWLFij5eFSUQcqf2CBgaCZkcWiXqc
cZ3JWjF6xu3oZZlmgtPmgeakVEVIZz32CDY2tLobg41a1OOq0udcKVTN16JM5VPG
vlgUotNh3ggdn6VGN5wbLe1O0VadT89chscIcGx9mQXRafXOQ0z3flnEZ5e3yNiC
mqq12v4Q6FwRugwQVedtsukvASzrZi9bOZUdefdsLD56b/+JHW4Nn0A2LxaK7Xc1
dfJCBTTCKoB3qy/IzgDpbvlW5dx23HoQ/Di99OpR18Nimd8xtoRoD9u7On+VLDXj
OcWXBX9prZSuykAxWehe908mgjg2/S8sa5T6blnUlVWY0uIIUQRdIVvCjvkNmDO7
lLMkjyjAJd5QdD40Z5L+vp2cVZwwFYThmYdQdtCONaBjcbJp6ZKFIktMEM4BU3h0
1QuExBJfMGdDdxdjPFlgJlHsT7WGRaIjBE6x+eYmnz4Xejep8ELlL9c0VYvB+1vA
W253tLbAbbvGVFxPCZ9c35ZWkNULDNyOQx3ZUdU2gXWPjBv6dTFgdA3UW5s5FsJX
cHTGOKW7OYcQKW4qDvWvVT8FYpL+7fbqeAr66wMDaerPT5UObS2okwEzKTaqTXaC
Rd6PLoMBLtryTl4D+1a5R5K7I6AZt2MHfCH+wXh/sGkS0WVIfXmmD7aEVYBQ3MYM
J/CE3SuH2Vp+F7WVtiS27PGVcj941Zm9XJiQsCQ2SXw8mAnZRbkKHcwpaDbXsFrT
GJr2jit00Og5pVQF0B1nmNJQj9a+Ns3cMM3JWegNBTtAXTH7ZCNiJfZVmU7a8uIO
eyVEgbcjEDywqadzYtVraa5/fjYkYQW4ZCCymbjr2Bv+vLFXVMTnWl6cVvti8C0Q
+OJ7llppKrK76woMe/Tiiaao3JfVShRNGcAQN5DIpa0KRyYpwe26l6YxIwmcVYaX
k3W+5RAxkLVFSfwtKZ2Gtue/WA9tUmfeBWQ0EpVNOZ9I+uUmbXvS+6gKm2lfUKLG
2BVio+XJPWNQ6Fy65nt3UKpblWrfrhu0p6j2R3w+Is22LmtiEI1CdwkhJ/71JhK9
Xw9bYM3DH1ag4T0TAlgbgsHTn3GRszoj4eZCcLeUf/1UwkzUBYPVybaMZ2+K6a3W
BEafuky/74iYU1MbQWcKWgY8TkytQNSJU8H9/kpxR/E+bOfJnqqDQCUOhPyhaRqm
shTNQ480XyrA8utTdnDJCXoreGmSCquhdOtSqy77c9PEn3dtm9Sd/VjRFCnII8WR
v7kqFBRXuJUFkUXCqisLZ82fJ6zzfKaFyVG27NhmLd4b+CuxHab0AdExXx/fDyQs
xws5os/bYHfkc4yXhknlUhdIvHCDWuvkRpCGnXHMYLwUA2ue6FFkMY1Y3E02Bicc
HBI1n3nad9cNmt61OIEZp69U/WV1xebqPqEFDVYwLcII/AmRuZEkfYwuFsW3SXSQ
3HM5w7Eg3p0Ic/mzpSEs/KUmRhYKGq8a3T+x1rTIVY+3E79W2se/YXZCYUdDS15D
c1KBEecwOn/FqjREoJ/86b//Zb/IPcYAUoFVPhSlxul8ONBfN/ru5OX4N0C/rVN7
8Bg5eYxzsKWIioyjelYScA7nnWUEmvljMAiIjjq8uUbCgpcLkwbBYh7AHhMBSaWz
X6DGigqVWTNi9NZiZ4yX+ZPcY4+zpNKMyBqBVS1qkMTIwdl4m7CmB5VhoggChPZM
n2mZGb0S8tXTkFyV/G9vynlem+M4KwK4FTi504jlWI/bGnCqFFr/SkZD6UFWtS83
JQGM1wUmsgu+3OMcMWX85SnpUUkQKfk3qvRupxba9WrOMUZP0B+o5GNbEcQVVBfF
AbUy0q474emEBUm3DAJ0CDhZJrVtXXn9UsI2WMD8G6oYjWZ1pifX9juhDfcRwNM9
gZ4+nMz307gbcVU+44elW40aZK0yGXYojdhTNtFD9DyheAuEQjPKojCucQMmRgT8
vd7BVBzAdD1ODdqQATCzwU/Fq0y090tWTMa1naUhZ4wkJzzhXxYiSTvPKJadkE9y
2TeqiO32kqRlIO4q/smGDnnFqdZmXQgZx7QyRmpktOxgn3yNhW8O8PKzbFTDwrqN
4wNxgf7y6d1JJC4SB/gEj12ZUrMnIQEGzLi6hlNmUEJbu25PSkpwETecFYar4uKJ
MCTCD9Q+/WOsrW12ps9Al5JCp0s4EsgLtEOU4FfJGF6yKCyXWYbM0DvGAy/0gIwC
DqIbJPre2UZrPxGytZB4iB0rZf0BiY9c0g/A40zBUfUoYVJmmaY08OuzKJLkR1uY
8AvrLoaFXPdUYzvSFXNSBWAEAShO/Lps0hzK/ba1vL1L1+KcU1tzgKjhzxtcxYnQ
Vo8l5o1JFlQPSVhL0gd9/xSFxY77TY55Eu/21/yVJgyqWZVGPpG64aaNi6uEkWOE
j9XizELVdowWhahfDIh4mBPh8lkVoJBn9C7JVAcmj62kGnyrKmFHZgzn3VWWKgYB
oI/ISOyTMjR6kJDoSXDLBNHys7Nq6oxtN/AtuYwdUu97wbR6Kox8wIVqQcLvlEhP
1is3vkZpkBBBOlldjXiLDekNp2psGY99pRyLUURwKRixmdJc4YdZ+ZjlL9DGwnNW
3RsYWVR2o5oruHvhnnij/AkoCmY6fXezU/LcekeMJ2Ho9hDaPvIRel+HC9H0+fYQ
JdS87ximI3jscHMF5U+w4q0QTduRU9LRS26ol4vudfWN+G5Bl3SlRUnW9yN/znEw
VutwhWUgi9u1magtOSU8/+nZwv/bQWHG1oTdWq566R0xl9yDTxuSNYpsM+IMdJy0
vFg080FS5ffketZb2biQhM59/BqmZkGBOMWss5UcFyAmPhKt3ZWWePhMYRqkeTmS
KQStSDMlg0nJTORRJHhkw+BCdWMDwmWQ+ydDFy7qP6fD21kXGqh6a1umHUpbI5/j
0nIIRckvEs1D4G+m60XLbfkGYr10K8nWMe78KCydffNPDaGlZffOj3aVv1f/QhpN
wcGny+ZUCetn1dzJ+GEQgyxDj2RBUpJvbQiLUK2ZSq7ARAYTokgoV/PoUzq/f9rj
YXFP9SSy3bEkxFCAhi3WqAf66zZYwdg8REWSQYyrC/pwZrHb5Ql5KW4tSmZRO496
1XK1Zvml1RsN3xOPknjVjE/rGXJcq7ST9SvMKEEPw2/wFNCjgt7aj41qKtwtOqHX
rMwUYjnXvEwaX6wol/6MlRmuYgqQxbkqF9XkpFsMHHBScGNkcrevjK9gyaMjj+kw
Ca9WDFYP+25hsu7lwsgujNQOS+Y/BZVL9Lo7rByeeAnbCCGPnO1EN1sWCvN8ri1i
la7X7krbhQADxbJJep5OdBAJPi5HiePExJuINJ5eVba9qG5izZAHQNd4C0aJbxiy
HLVTReRK99mL+/cD3tI6Nwzo05sAZ7LEKWqUYomqV7uAQ9jpxIwXcMzR955Muqt7
eYCGUz469Y7ORp31KhnK+1nBfKfCOY9I8YsMjlxtfVihi3+bh9Gty+obfEeZoh4R
X+fl+HmcaU+07zKQYorhcalcb3N9CBvfAEt8swMa4nphag2FSdC/QZ/i1O0YlcfO
6Enpo9P6/Wj5PEuJIz5u2KsDFN4/DdGLj7zmjUoYho1EoI4BFllHEpCBPgv9IZ2K
YC5UCF5MSgoIWJTvrDO3ziQD6S1EQZ6j3H6XAamPPkf/HWbRCaoToDV7UOBOOYhB
xguxYttT1WM199Mu9s4Xx7qi0b/Z941hjkpHYi47giOdBL7ZfySue8kcAyea+I/u
8NrfMtvtDzA+Tpkq9FSkvl1ChkjBxrAtEZopVEF5tiB92FRLJMFzoyi4Py3thI5v
ekp+oQ6BY/Ukbzk8UxUhN7MJJgVnZwjlbfVH/CGrjqiaPW7b4U99Nf5wLus4IzxZ
cv2tQKpJSvhl0N8QqI63OWabujCnX+Z6e9fu3rDNnNQ9Jds1Ver84s5K2yvlVteI
mVmKPwQ6w2/EAS5jm8J2cR7OPlSML6GlWPZB/LjQcdvSJXDE4LDbX5GHgKadwvOG
emPS6ai0RK3TVkNXyjYvWItB5lqVIpYq6qcIwJnZ/RcxY98BRXWc1uKfUovRVpZp
yuTOw9V0kcFs7284V3EXHY/4Q3rM1twdteHC4cMNc2iJTMYjHpP29DPzloiQbbfh
VX25fJ+AcEOgvBNzPro6y2m2chCYRUdGNtD/oDLUGzp4bK0cuasE/OxuU8YdvPGf
01+yKrup0U5/9G3+GtlBLJWUYrzQ2qv4SOxWQsrGGtZ3r9IxhnVNfv7/fDbKhRrz
q+aJYRAc3f8B6eUQOzaD5NW63oiLQCHgs5VIXeGfzoXPV26+ht54tbjCQg+0fztt
9JBuMIJhsBPdfyxvj7yaSdjy1FAYLhwAHxuYsAkfdihhifRHV/MQPBtbij/kj0GA
Y9gykhANxxdnl8IiWKpmaA0eiyr8Fg3S4KDO9v2vBPkE97SRJSDo0tMJaa7AltSV
OhHDKCNbaRe2XuEtGOXde/6r4CEs5R0eTT/PeWjbQHuTmAzhImQ2ruXiuRl2rWME
1cPeHG8ardePvd2uov96d3C0FYH3Je973M9C9xdQQRP7tDCtAD9Zx3dgDINhKwYv
iIE0MXWhB3O7OEvy773xgPq7RFLO4xq/YYA+HpiezcEY9hg0nT6xrry8ILtEpJfW
O1DOx6nhmi7GwEHKSgIq9GodvOMF8A25t4XKjiwmSxTNG9TrCgLqbYSkeJ/ayGWj
+zfxJHNAH7Cz7BAPKsHBwPbb0dPLXF14797w5HLIUhRf8R4YH+Ay6Vgg6e/CoOn+
FfNPPcqZy5CmF5EcxDrKFDe0+b77EIfRH5epv4BmoifrLyNWQEkWXco1dDCcInoE
BpqDBWGaVQBKOxz77OyobIoRfGWZ46XqLOlWp78ePNb6yle/UVbrBk2cgEyuHIXe
Pt6U9V3A4cwbtxANdXMUjb+OzuCIzvqE33xm2RrAfpbmVT8cpHioV0lTDLrmzn0R
fC2uKylR1pbblwShXNmKFSA6Q4EM0u7utjaSzM3f9AIOIoJxRK2kUMK33OpQLtUc
J70IScyCamvuava4tM/hnwS1zZpQiBFnJGMTeWyuOf9Mf3ay34YJZ+ZOZJa8Hhce
PRB4RD0wZSDXcKTWQ19Vs1pUjEsHqpRXf/BMVyLhDNB9kgR/jXY5jfapOepxQJ/y
YT01nVwURbpE2atJMCWlkcg1I241JZBm+tUMlkKkQ1AxisigZQJ9vzMlnWO5IC6H
ujv/4v8EYib9vYPdtOoBo2x9AUlNM/j/AnP+CD0RIyaMLgbMEfM23aMo3ufbdfZV
7Id3/67GcFYT4DS0OUgvqSMCy02xcymfgb0iUHpopFETqikhrVrfl281WkBaVf3y
0sjdVcl0L5qoQVdVhdL1wIVyYCRf19EJT6up2BhxfJX9DEKFGVfstMgv9GH1FdnM
GGoTsiW+zah6vAsXGrAuyEpna5tu72Kiu9R7NvyOuPCD1FMCXvpa0vqGr0bMPZJV
8X/RslB/rX02m2h8MzYibrU79sKHGePh7wdsENf5auVWX+LpL6mgAXAS7Hk1BF4A
6StHKURNPNFy2KtIfl//ntqoEMYpJvBMa0MOzqLUK17+b7AQq2Y787Xu+u6GLj6/
el68jXJiv1mxPc+wscgu6ca49Ku7njDUHAfKZ6Bo4Zzz7xuxJWgJYtl/O0LsX3wR
v+N143hNDG7HOPaP8awqHDwlGHBC3D5tu6y9SXAWTrR6CSou024ZHuypqBAuQQuA
aU48/AoMSI0/GUqewHZnrdvA3LzmIkecZ0YufSqGoduUekjUn/XJHgPdSpqManN9
iTqvon49vzYdWZk3klmO/bv5vM/GArvq/tVrzpTFuomYTZj1h4f+Ofs81WqjKcwp
HZ+GvcrUsZD0h36MqkVDPYT7AN4da1FeiiGlmTBbUSy1BStfKmjie23eddZ4dfp+
U0l7GS2VY5DisalngrqOCzNZOTkrrm1biKco47o26YmIR4DAR6e7W0SJUP8sne9t
gd4mXVlKF7JM0fRDgEXWL0Xo6rFV/oGlG4x193pFahXfPTO+DEDW03nByw1waJYd
S4en8EB01R3314kmuWY0+ibZa9G1HCTIrtp/Orc+R+JovbI9I99RS+UkF+VBbsCQ
aikAujP2MQ7aYtyITatglQX4IjzX+5iv6a/7cr8qCwaTDMvt7PlP0+5W5QEx25KR
+P+xnGoLrCnGC1HyBQAadYvZ0LXeTHp8gsAH/Yv1LiThoMegz5Wq+JhhigbT9CGg
LSSDs01kAtDMWDUA7krmGR5dqCize7fy28ZZ35WfmhBZaTEtPFUD6Mif4Lfz2Ep/
So4tPNlZA5rpQJ1LYurafjGy1xXw8BgPfO5/wXPnmzBROOJQ04rllKW7ru6Cr19a
m1GZNcm3N0KmRquPpufAs5l1dnfHQw+jMa7Pg7Xt7vxSQ2R50GiVHv394ZIQgWD3
ikv64gpVJWAcFo5iTtLa9LQiK0y3ZLM/MuMXbnBxYd+YbiSM015GIB69Aael9F9R
+Hrj4/Up/vOFweQN37qXgJyJ5D/rJVft31FUhMVKusWTDejFLWoJyhiqcdf/JoV8
qSSCnZpnb3NQgcrELjTe5sXdb34BjABQ/1DqA6TqDX12j+vAaFltu6BWUMsH5Xa3
Abl0sC0nqjRmooVmsXP1Z4oUKW+rOZFQ6cfL2uGAnAco4Db8A0WgxWzcCLQPayBx
t4Qpvc6TO8GicY3e8FAS3d123oBIV/W+O1V6gZcoa+Keap/qP86sAegyW12sxlnR
rpJVoi3fKlIrcVfIBR0NBsOPxYyU5FRmAshhQ+eMWvKbOx6fB2eHRDsg2jeZmN2l
V3N64R0kIV6vUktG3fN5aztEj8zBGrOA2j25e5E/Omt0dUo/XStavgZpXGyk65VF
3D3OyVpp2iXPIu/+Nm0ySIcifzJNJK7WaHB3gqG7BC2L0jOKYusOqmCy2Pe2t7Rq
JjrGeChuTSXaOhdELJZ863P+yaqO0aOBlETXgBbOWnbw829Kxw8C+rxwM/sRH2ca
viY/+VcZcYmpnjTxiC+GExxPpWh/7/pHyuYE14HEopf5Q7peMl96EUpv6ERwNiuJ
mgtzYZcz3UonhoVer5Htf5Pv16DJHCT191I0m8FEOASxI8U1P8OdhTKliadFK4Zi
wypBv2d+0xUM1fvi/64DkZ0jS64v2TVo2drkB9j9n68/KWRFQwbAunvlsPTRCkqi
2Zi898WE1vYLz2cDLVYvZbI1LX51PFMXCe/k6q0GrcsXW4pfg7yW/qydU+HO1u7j
J02U4Hw1Yl+dtKBZof68Gdrt9q9vNjmHohuYg4+jG64DVGbQPeVxFQkUj3IRkCY+
mOZd4yqSi5mkEigFqjPjug9mdvoDZqSfexpjCVkF+22bPUin10dHkrlRpop/4M40
jA/svXr9KROptO0VWkT5QOdM+/r61JqdpdzsTQY4T4OUB8gSgGRbNhmTtnllK4y8
tl59FByTZH1RUxNMK5zf8yVO1uiPBYkUz3yalaXnKkJLawhV/TiyfbhMU69N8QAq
yyAyqRpaCC2kua87eLAI7r0seQhWEOiezXPC2lluUoul/c9wpgPl8Ifl5tUlbyT/
iO2mF6KSZOJyheN6ITtPM+pTlB5C9RiVZPOie4VVbE9wgTWUKGdT3bCC7FS0v/kG
zVVSswTXK/opTKVUpzpgUkC7XFbEJDDqfQQFHyvA3jtYifEsjCzH3EMiYU1Ax4bW
i5nxETqhqSbcxW88ushVcOFTqO7EStEQoalBv7Pvo38okPsu/qWA2ndOtmn1Dwwz
ezIC/OD0TWqUApRb90229QF8WxFXv7ky2eWlMY84iei7V6R5cWp8YV+5lBjM6v3R
/qhcbneQSyQjCwf2hBV2h5ySqpoYnZZThA7Qjsh5pxFtVNLloxKUEGr/l0m02P+v
8449Mc5rOJJBvNhbHnPEqGUyo8gxz64oqXp3O5OonUyQFPZ5EN5meSPOR+7+xfyE
dsOnkQhU4/AkXQp+DNfSh0pCsSKYu9Bd/+CBeZ/aGG/BFfek8L67V2L8BndXDqRD
49Hg5Qp/+sMzIAnzyuFxELWi2Sgqk3sxBUldcmUb/qyopusZUVDUM7wHckUAcffr
X9U2Xw3ytqYj5/ac7uEKxiiX05izlUDfHBfx7l26F0dVo6Fz0IVcu7aF8Er0h0U/
x6tonprPtnkBNvHQEUSk39yUb09TkPSZHygJyaWdLB6nFVQOjCEUQHCEN0jil9Ig
mAMexbkQ2/wllUpaZHRzxVAy8U3zdRnc7F0UrFskR4MXgPixtHRe4WVC6CVryxSK
ODEZZS0EiSI8ZuqV9yHUvLDfhcT/wVAPePEJb+0aN7Zx3g1PqKwWlcl4xZaxG9Gn
zEpCQ3tpvUa0xrqZI5NXqSQKraVKlNGE3rpaWUy7jh6vTJEK5nfqcwkWv4/8+oEU
efOGoYRUu+fwsAYfvmZG4ECPIpgI4ImHIIESWhVva0FHtY5DCdRC3R7Wr1MPO2PM
XIKnrQF86OeEMPp/7mpCn3iWeU3/CPL87CV8N01SOQg21fywMt32Hr5YuAk+TrqM
qPr4+8SehgpAiO4tx1RHwp/ijCI0nPq6sdSww8odipy7c68z9SR+lZ+ztEyrRyv7
aDnXV407G67CgYTOVT8oI/F6sjaJYU58h+wdsGRt1pf68uRl6lw8AxPb8BL3CB/h
iqf/s4zxQUfzaBYkZA8wGyGlvKT84dXqSVq51lZCuN9y+LnXKksY4Zl4kaP5T02L
JXvUP1OqtgvbzAI4Ji39gJlBafnseXalb9UeOj78K9jlHBetnBF7Brljv9CeKKJp
hInDOYJjCPQYxM6tgdj3ZoN1dZlVBa5YTjrSJj/1FepsBxeH+IoHvXL7+NRGsf2o
PGTXtgQi0lZKjE0TGcdV2FicqRFzNKepO22H625HwPCTrlFHht435Iaq/sVDb+I5
lfoGvaM9l1s0LfxZwi0whq7q0M4CuqxJEnC47OHLOUSp7nforaVihblFxd4Otfcl
m1o1L72Iuqz2keks9inP1EcFb/VLWV0RaXPYGOrAEqb8oaAekYlDE3Fg1J1StMjI
yD6O0ENaSjOvy/m+qw+E7quDWYcfbLoUpqAOraysCQHnFgJqn0DwpzYy9T+GS5pk
560m0wYEih+qk7pbfIcD/vx5VJa7f2QZOXigoOU/vPDNuTX7BhegXB4AaTK/rSXe
pC7wWWBQ9lEHuA0z0vN3rcuVDWvX3Z9sGlezFd+mhb591wj+EYjydK28AC0TACMc
9QnHZNnlUFQuTxdZPzvp3cwqjxcpKeze5grr6adQOurykDuNXXsBGFcX5ziPALFE
z/cleJQakV4plYh3xHhJhkK6A2A0Pr9UY76vD8DgCqgxu+XHUmhtPxtPq16U4Jb+
Vsya4gQPgLe2FdbVMxIUlVbcLx4MNLEC+/rk2Kp2maFQ7mGuKy44V5dX30lGcmZy
PL16HSADvKXRNyHVY7n1QFsFO+Ec8Y8AEXF2EPSksHC3xPpVUd2aLoMREHUN7Efc
2dUfuk4C1EX6psllcnPDU1GzRbJpOmTTbZP0X5NSQZehVCE8bMn1SQRuHpFO8wDm
4l73pXs9qe2zSKwxUx74u/oAEgYV7YaI+D1yEQUiXVnkWmEi0Rveg7rcWthbOatj
fzMtrNH5RuYYzSLWVqJpdB5y8ZunG9xtWQ1MNtNt/IVFgaq4bOeOG9D+P1RX2e8O
vYb3YGboxPWMaSeO7cTWBleBc1C63kgPozgZaP/JulKDUQbX7gRWW/E0qaM1gklc
OcGOVuINib5gR4OxMexFD2bxMJtt3aNAldwl+TKc1jshpKsbIiD2fa0bOI+cjk/+
wvQ9VMemn36/zGISCGAFt7plMeqv1q2MMhYlkkNVPGUuMD2WBT9AnYorweFnDYTE
Sh7kNzSCZ0Yhh+Vzewvs3RhwQQqtg++hcUTLU1BO9MNJSrBj/HBdn+SqeOSgBZDz
KMY6I1q+IrltJVlT6zPaqKs/wdsW7eCOueOSLBUTMDTOSO1zFC2LTB9lGA5tSvQd
95HpUfek9yTsPG7UM5g2g99X4cAmnQkoMBT9e51wvhOPhZQc09whQ5vUneEO7+Ft
h/5419Phg+8kw2g2eIq91jmPR8olFySBz3TfZrA+47O97OwGSnKQmpQ2gM8KCSJg
nC2ZeFBkG1TRxghCD3Mhc69SD643rDE7Lr0pANJ4DZ6zjglXik6ukgC40b6iPHSk
UshWAgj7ojN2vWewVJhiiPljo7PwkbvH8YzQMwFM8xTXM8NWsCASDI7dX2Jw5+A/
6BPEP3+WufyxRIW3xGy6DTacn4y6RqnBxrtaN0PLm6scpGA7VfNsytq0NGjQidNd
DXIT9GJqz+MbzJOZ373pO2TyMYelYoTNeRHZG+LIfragvslRKQHvdPbWUam32FV9
hM1odN9SqZXcjuZfAV0kLExVgEj9LfNIr0yVznJHemD+55HqvatiODtsAOGQpypy
qDzZJI+xKuil1QVIleEqiZhSilHBA7OPi49PzPvEcdClEM5KsOs1mkrYBvxaHTSt
vAuouXYkqGr/5Z1BMV8hjNEhmuvHwJIpZDmXVBb2otCMpHGhv8E6IZ+1278KjcTo
qnkSmF5v3+9DQ8FRg17lU5IlP1FVNz3SIMRyJvE8WDEc/d8midBhjN3pLseuXq4I
KdJpaUbZMA9GwZ2hSLf/hDQNv6LSMDzd/tGDp1ynKpexGazYaUc2gul/OBG3HVaA
OVOsw355W6d072AO4Tfn9cOsSvmDUiphxntBLq501uaaQkTUMOAvz2we6npT1lBY
EN1OFx4rfR3gqxVQ03rmdcdrIMSoOlTny8pTTmHYirrAQmrhVx7F/ZANgAtKHN51
8ncY68zUUfkbmLnxDIbekEPJIhmIsEx6D4n7w7NotTWa6SlCA7ffm7OZI9cb6XWj
uJ73Jx1J4aD8y6C8X/CTFsksRk5Jbf9kh9b6vm2WaWB5+N9pZ7ANgs7PKdZjdg+Q
OcUK8eUrKDFGL0c58MhWdD1IdXYdDG5JNkoApcVWOjCIwJfWee6A93pK4AmKLOhg
lH6Et47pbu2gARj4yK9IwvGO0L405zQpBizMyJN/bQU19uZHza0fVJ8bXRy9K83x
mNiuDuM8dEZS3hnWZEfEcPBUWaN9nwORCnnFKb6ImlHRCLGUXRZQ6yJOTG6+oTZ5
SBht7wR4ohMJwgBKh37x334pgIEXEoLuqvnfXYw+BmAAxDoAc81FuYqnsNpCeTZj
JFyyb1XgXNmGowNYFuw+DCwHCiPFY/hlNW5iNwLTCzGr2oT12FQ03/Y0Tnepkl45
MWvk3kLnru3vC9bUDWX8v4+hI/G3IDE8pmJEq4BYFq9k5DX+GFCRkBQPoKzyVMHs
CTbBJoynjnNWfcSboYQOM5Iv1865bXr5uISjOf5AlKYwix8GZ/ch8xSTrzrG07yo
FKQkt1RiZCa4MAeRneKcW5rj4QCF/p3NLmEnN9LWNRPK7WUpujf1I3eASltX2a3I
SQoxYdCcTYnV6+utIrnfrMKI0ZIKn+mqjp6z/g8N40Qf06+lKlHSpfLBe+FJZ1Mw
LgNSEG/2S+grf9SgSautZfw5VJ8Gth1UXFVj3AdTlP1CtYg/jqGTiI2FunMuknrz
g+zjc+7YOYcwZVVwwmNZA4KvbIbspYufD4vzBihxRy+074CE3pv7Ag4ywfUlalPM
1jC+IjNEoZIIIRwfn5kuJaxPEcoz7cCQLaLZ/XtL2y0Nr3SgEulYMRVqHUiYbWbt
dLTt0SRtLCEivvtxWN8CQybuWv2egHPssZm53/CN2fXLtniJUkwKPP/YqTqkrACU
oLaxqFya5VWjfV5Oyqg3J6aBngmdV1835W6ZYJ+H3IwPxoJqhu38opLj9QyLJiNH
rv6GpQimOJsD9eXFiXPpu1j/MpgrJU8nvme1eMDEwrm4ZhLQRy/sT3M09hBcAbdh
RnQw1bawXHGRFY353tIxG3Nd+2+Q9aDn1aA8aY5YmCyFDB97oeQo/SiSuy1UVDur
MR5b2rSDhgFX4VRm00Rs0bn/iES+gMXZvCX2ZtMYP9L+ktYfYiBqJ+IvDjx6zCGi
bXVpV0OpEmSPZ4qyWa7wtvbZsessEzA14uHC67ndtzRGBPZZ6nVUbutShweLxFCC
A0z1ffuQ2HU5nBvYU2f5FvpgHrvWatku0PinxvuqZ1i+lQu7S7RYuW2SgRa6Lf/X
QvG2auDnaC8ufM0bWjhJRRvVSbui+XO75wmCafWOqQ2KTfXsur9S2ct+1Wn3bKqK
Xv04sjh66ZurZkwsy1ldiz+OgnzSG7gYVkHRKcT8cuLtbV0gUlGIgSxb+lXq0EGV
4I4IvNyEU7r4vFXkxTZ7Ebxf+lwqOf4jzzn+bsc6QiPFFB/zFF9re0HN5xIBC3nn
q1S2RiZVe6SRl8JyXK99DjCXu+FvibxJgi+GxrAQoCki41l9jbN0O2FRA67y5qOx
qt3yajaFTkRZB0n2O8E5eJQuNzBZLfgGkjx9i53gx/wa+UErIGDjc85Hz40cCRzf
JXwC9N0J4weue65jCq684XgLbd9TbR9ZpIJJ9wXWgkVZ/z13WsIwVDibwJRdrah5
9zWFRej3poLX13dSnJJNteAEFNaStTGA/zaWSkcQu98QqYmioqyjr0BdKpZjnACj
EeH3nFYTJJaIIjnAEJbKIOiiyn66xjWzjjCCRccUzhF2rN4ygGw35CbCKOs7Niit
umJVMKw27s/HnVfZurr6298bz2Uh0W7vAQqsi7tHwX70BTr7N2KD5zMHxUYwOifc
rLpegB78uf2j1Dyrj5U42X1oFq6jpn2UPOvVdah5riT6VzzUHCWVK9AjX8X6rYRf
NhzeQqIOaCpGKFxwI5aLZQOzMeEaIu1wysqiUZhnrvrNoOMINh3ZaWLyJUpe3X6u
xDZZHWGFLAEM01JgveRty5RIp6LGlpC6lyFxlyT4wTCInsL61+CtWhK+70xfXQYj
VEk8U8aefmdmkPHIoUE0oRJx4J3pl4eL7rFicKgY8QGKkdXlHsq4CCHol1N9SG+7
jCS3RY6Cb5BPPKg5O9S8DB+Usv/UYz4PrmX6RbS5ZZZPFalVeKW4yGVKi/9mo6xK
eCRVtvVlJhGms0lZFbIdf2VqvLH9zHPCHaWzn/d5IuNDzwtrLWsL2+mgVw+0W3TV
6/DafBP+qCvXrjOCt05eJndiV7xJpvLtxT3eMyvqSP1x/55hJgew3r2i66BzbawD
Nl51tjsPREnzUz6k06uuZTKPEmYNvPvkB0kkTmReYGIbpeRWZbXRca3mzIIyNULn
Ej7EyDxtkTg4mU6Ecj+SvS5rMC08+7Q5i7CMjIisb53ZMWa44BXGwgEPMqnOBUUX
udBpTC1zHqI66UZIS+eyMDP8wLKTpIh8g1iu3xYQcT66qcygiish0ugQkf1K0Vv6
fttPVQB1/f0aKXlx5F4qUbcT1bPPML0UbLeD0CeKTJbhGNNZ0y3BqfE2Ml5UY2+q
jLfL1ZaDC7hB6G0yiYxQiVeJMh8B/s2Rr9LrK7SibzU0eOBXpVg3/5BEnd5M4n5l
KTGV1BvnMyrDX8AGjubm4X0mRuxpq/A1FQM6gkslyJoJMz5VvlAn3dTjuJkpiugi
St3SL6MnSl7ghYVWMlA3hZaqx3e5nZ8VOpxIfqun6ND/PLynoeEJJ8nwIM2CHJuE
RzrgIxSAgYSJFyx8u88EYGk7HIePUQtpHf/PDk8EGHmhHSDB6rCAx7rv2A0PtjMy
bcoAcmuwR7vQgoo+XZHgbAY//edyMpWkm4N08MMU/E2q7B+Ug5AHL96SQiPsxIfj
sKNugaHAAFIohLS8T/F2NztwY1GbEthlWJCgpMDKoea8SCiu2qPnlbA0ydF3WW7O
a3CCrspQ+aBxt97j0/pAaoCBlZaYF/NI0ukc22G4w2FtChs+1i4NJh1n5jflAiBH
qRM7L2tskeH4GM9lmSjBdX/2//rJY1UdrFHEHo2Reupm3hR1t6zeZC9EdGjGelJ3
aH2DZ3wMSv7eDpvhIuy97OOG2FcXSAwVLljowLRnEv6ti4BRQCOk4oeIfZfMX+9d
dznK/dMXhv1UBm1Qwq2ROPiboqRnaBCNp4bqVRB/6RQW/cwWcbS14Ip8GxeepybG
W+hkky34xcD11lSeN+9iaazJ2aW/XfrzFDdaPPtw/+zaK2CNpufCmBtVTr1Uv3B/
3Q2xtJ1uAFPMK4WHsFD7XxyCVJgUJqtRtaG4jx6cEa7fySEw/WVevJG6iJcvB7E0
KR28QJGy57OCujuQwT96Z6sNSYGhqTU9NtFoKdr8U8Ivw2zWBWfqKCZp0MfLcyU9
N4ksliR2RjAxIGxTmQohq8/oSZrCSX7dZ2VaATO9QQt+jmxczUJIW9n8qaiBv4u+
7u1qEidU29VBKqme4/KkT8Ajc+f7Z1XXB17DqBJoVmg9U3QZiQIrG1XgiY6EfOh0
ANRAcnHYrC6g3n2n3WvxVCJpODWQ8sJvsZWCSk47WhpFDtJ1Yl1JgBX8zXwkUZXZ
TZwb/psnerQeum+koZ7b2dgvUceVEwsxv08v7TZv81FDIqRmYo3PEb9bJOCmFVNu
iXAVyVRWBfFmthLbh1RepJ7HrYSGlOJM4UajmijsLL7QlKAUHb8mXjSmRqXeMcbq
5eO66bQ5cOiwszdZ59adWwmhCIEjJUqD4xkWDG0CzktN/8NJ6D6JkksVzXKFRCvp
KUdCNWd1GStT2ErtXjkuLahBKynI5unUmtwLPbhvc7DpK5/+H9cJOmv1MNZJDB+L
DpsTohafRfuZF1G9mLt9BBzYjCziHYxmhuArM1xTXc46AVxGSdSJgyEY9MYVmAqV
VrctCDxMokYHdmDBhgaW7QI34S9xm5YiLP/rIhsGaZ0VbPy91y5CzwmPyX/G3Y7b
H7Y36W6V9yARcbKlyqJ58xML7/AVC7ZJLN7yOnxPDgnV0JevId5VYAXFGTheSe5U
/Cjpj7YU8mK/A0HCAVqYiAn3Wq9WrqiHTkiZ64FNl4DGl6qYq/7Xf0cY66DuPoHV
A5LR02hNzH/+JASqqfKKOFNcEy6qgE5te3KOKKdw4uY5FjQ/yZrtCjBqVb+zw8fb
D49ldlpzGWBsuFMaPNuHK45gXD55dABlnSPhrRfTjYdMbXIfD4uWG4ZTHqsRbxzk
DIGofCC5wTMObJQWkLQZIakVBtCQPUGVMx5DTur83mwQ9QyVtYXogYu9h3Hw9k1g
p5l9mMGR/BN3dRPtNBR+cEUNNolBryK4Qsix7ROL2eBVYDMn49+K78aydEqr0uWT
bC7lUMOQ/lf7mtdbGBBJKW6wWI/mDSl/ROhltpodEJxfoPuww1dmk+Df1gtWSdQS
kRoO5chaGB8p4zqjuX2qHdMaftIYIuH7hOwWtyFzmIupazSh3jKS0w8xKE/U7Ch5
duRO/QI2CZaRdfWDLcCjalRINPueSTm/LOj/0SEcZlqYBqZ/WYnUNFVFw1mHKbYR
67GBNJCsOqWoTjQuE7WD99PPyHFTrdK0safp/nAi5h8pIM+WLCH2Fzps+3tQvoeo
362EuzpjWuKDge8VwuUGABfWb445s+X9tTJtUfdlcOXpsxSGovom5EuPgTg5wAR6
6Dj/kMtD+wtLRQDRVMhFdw1MG+gRdsb296IslZwzsdgpDDRpPce72doofmcaD3cO
ffrFD0ezgOJk3kjLHlK/OhM1bqT6gHoP3whSytEOEm08KFBCAOEbkwUxv6Xxz0/9
dtWn9AKEcgmZsifPWK2OiQ/mJv8PimE4lD6EsEpWjIFjqlfwcNB18r9trllLB/Hd
BQz4Xw/vMZ6YDKvbM4cmMMMRgiyASPTtlwa2RVBc40CN/tyOjI9UXnPrT7NqYrB9
jq9EKd8jZSGWC3tHe8Nx9YDsZvxrpZji6QrG9pmFq4chgNL8lexofNWB330uWxd3
ppS/aLTW1QIg2NJL3m5nQJd3Gyr2oliQ/+1aA9HDErGSiNhYVtcht6m8/feS0Zma
uu0ZT4G5wwnJEjVo6Wtrqe1dHHM2kSrpwiU/vw9QW5ttc9j7auzBfLM6HWRXV5Q0
FFmtOlhG5gVVmHvF5n9/TtKuD720MuJfblLimaU/+H4R37mxB9V2Q9Iu67Khsoet
S+3VnNwtjSGFdvgcFgYTUUyFXqagCcqayz4dVFh+pNBol39jplAj6fez10rV8UhE
6+gUbJFrqvSy4n4eB6TXt4zHwLLAvJQMGh2/VhtbdDzk55KpN88tKV84en5fcKGa
bMaQQq40i/NXHgGtK4Iy/cQIzll39zG+3rcsvsJXKH8PBt4pXeUeZWthjVbYWXC0
n1HCdJSFaTlcNIrvFGCGVqKwg+D4MRJA80YFDLjN/u5GaKzhWauKUCPoMkljBc+P
7roPrzI/c6baJDmx/nvDpeu1x64EG4D2gFwvW3k8agEwkyhjgUlsdp5IMpq0omD5
QSE4XwCtu73imKiYBCG+bHEFsHiaSIZQ4+OYKuoKUQSyfqiLhQNoRd7U0ZqVESEK
PBzeTTU92WBDKj37iJ6XTxjQYcqsXZkVdPTZcJFds4eUz7zThaknOiv2QHzubnuh
+6UeX3i0oeY39GZiTQ0jWiXmdLrgsdAjzWE2ya90H/m8YdkLI3/RL6XSRg4qR3ry
ascux6+YRjJLzKFcl9HmEcgnr+YW0r6EEbfmhPFqd3ZwM2qWSKEtuHMviPYk9E+q
CUVMbsX8k2SYU/Jm5H4cehv3HV0I6KVwmihrbClZcigqvicZnmM6GDKvhwIS+u4X
0ZCkix51Lwb/V199HACYD26bGJW2VbBA+DTWiV7iXaGeakvOtdGQAhrui1M/o3Mj
Vvnc5gwX4RMrjrC3oczSXBqNaNJXqBIreyYmnwCfg8ll2iFMTXsC9Sc+JwIkbwde
mX603WG+SXGMjL5baBiM8oDgIOdCYACmNgqVQJM+n024oh2K2PPvuMi8E7OPZIjY
IkmNyI2+q1Ltf3I6NsEK2Mgf3Mn/1VKr8AWaRR7m+55OUyRz+6S5L11w/KmzjxUy
SIpAnepg5JUThbBm+n1JwobV0vgnwvqKz4uhOp38w/zgtOx5WPE2rNTzmyhhLLeo
AAt3NQOfU3HQ2wIp7dp/0gK26JECFSwHMEr89sUh2MA6GQIOmpgJEs4LG7EEzJ9c
Gwttf0nplINKKXFi6kIAEqbYkFBgnIFl5OiaOqkW9BDB5AonegJhyhvfwn7k78ir
ZSS25ZlgfP86tyQH0p4oazNESVZHMLkPdhjXDqhRUrb9YDiuiGOG6tSZyt2oYNKi
/8fhozjaaSeYSnpzw37yDfGgji/XKMXycX6o2pjYRx9kPth5caxCoPHn+C2tTnHT
rac6xhxD0RM/3AIBFLV1+zq+lioAbfFv1aTWhtsJP+QcmSjX0nqKHkPkCALxdyXd
Hsw3zzpoRUlvCi2ODEP6B/GSZYmULgFqJsX+gxMsTfWaD85U+h3JySOoWuvdpVbG
N0S3enQoiRhBTPiLA30g1dY0yfEzOHFkPG0mBJ4JaixbRrAscyExAKp7XpGLYnNY
9GvCkHDosVB3bdgs3ZgD7/6Efdw0FpOitJOgWQWvcolkAuPPBp9cDidPbblGrGHW
UN+vtTDBAaY0ipFTIjPFu2is5rwCUUMNx8uareSP41rVZf4mviyY2MHAEH2sEXsf
KeR3TEL/oNxEVjet5PlqdCPqH6Z9DcLqi8NfUq62e+wR+h0nLdIEn4nQ9Ur+u0+Z
7yYFUE4O3o86y3aXrpPrHo61u6CqrJMdl5kxPdt5MY8OxKFPALynSujwd0JTsljy
KBiKZo5byf4lyB2XuByJyNCB86l37xEB6WeEJPqqUZdlkLpB0GYBBJArT6TEPdSL
mrPqP/ovC6OpTTt+V4Aewbx3Jhbk53FCEr8SiCbXiBTPYOUiCyU0ddHfU6tQjs87
DbWwNz9+WX+wWicqVQADIz0ZsFxWl6Fich5Vr+OVFZUNJk3/VpEQtYKq25eGVIUT
Zov02kPCNGVcbyVWrSG8rAihv3JiiTxDxsSefBcgZDjMDGvPM6jdvGj0zsdI+/pj
xB+vsSvxUX5rKtDcEuc82nw6huvG1u6QvoMmCItVRDwvdxkMNWCkkbuxDfyQbSqj
VbT/EK/Km2cQa1tu2KpHzwgYXrwfkLan8hytqab2Xt5uvP8WC0BooT4C15OwNmpD
tIoMwyvCOSsi0hqiw2rx1EqEOLYtYolmWo9ta5825d2bhSvtAxO0PWWUYypeQrsa
r4xMPwuv/Q9GZxkz9G14k+THlb9JOni7vqNs3SGX+6g9XXXYL4Cu/qstd8QQt9SA
vLB4f+0whrQXQKWtFLwlM799LAO+wFNOcxTXuukaTdoucmH4PpGZZ0aBSg176Yrr
VYQyx/WLFIEjctCN00rn7+ETAGTGpZD+aa2ayUnZRXvmxKE5eU5QfoY5C/rTkU9v
WSeShB3g2gUvpxS8WF1tsP4Zr91KE4Kh+bEIoIKHYNGEERqrLBFf6WQoVGUjo0cV
5/M1f9nFgRh8bPddIuzJFTILFzWE+UbDDyPhGfhE3s4qFaRVh993Fve/vl5nH8x1
NhvIV/fkJXzJcoUnus1pzWPOwekuVT0YNUKyKiafGqNOzcvMAnlLRz1SaBNya4ix
s8snvs5wksxsp5VRpQdwiGp6NDe69IvnQQ93MU5dpVA15NZnTc4TrmEg3+bDsInH
Yu6SRRz3YUPbRxEWztDzCHinTdNgKw5MJgVVstNELRGezBatkCruK44tXrJ/BaRP
luc2UDJdLJJFX7WqMPvUahTLn2QwZqL8jLkH6gi122ieI/LES/cSvEpvl4TLIzoU
iRfXAe3qrHBsVBbV/g9lEzWIY32hqbWI9ErCiKz21MUXtSauCh/xERMGw+O3T82C
QzxtDxEXv3bSljXqSatyZlXx1wyopxG3zjowCZzExSHcn9JT1DCtczuU2AFeRsSk
uz/MoWMlqm05Q1wrlVRhGj3XKdz8UdmbAdzyaNERohZ2gJmOYwuGh2A2VV0tNwq5
PsNxrwnOrGgv57d6SpxQYrt7TGj7pBncWTIAGLvFXPeTWctC22/dYJIUvKaA49fO
ErNSXbS4n9X4Xov6u6SkbEZavm1R2HedxQW51g8afKk9CKoeQbtQcW6mlwURXMoq
4E9LWwKLFoieFa2tVf3dmnaiRvBc7+U/aJmXCd314bWo6YdvJOxOIGX8nNb6k+Q9
X+x7HRqikGSKHT8KzPAj4iRPlLenC14xf7iVseFFwC9YS4GzTTPWzLyB5Dh+zuX9
6AswcdgCl9ZbWOSKMgf0D6Bs/jX0IcKdmHG+tXgX61GriRqvkZ/eszyLV7NJZKIM
LQqo+w3KXQ1hLT9OQfEZHeY94VTM/dFnuQazmUeIERzyH9iYgIiGWL9GJQm3+Hvz
8Gh3cYAPZFH7pExguRhF+KW01XTDrCx6rqP4DyxEom28wgUhoLLm80ojhOT37ccy
U8HJXYC9gYFlEvdaUGt0IiUfGh3Gi5RS3oKFAgKeL3gehf2jbFlYQfQB6p+3vuaw
vbeTeS0r2UmRaPcFwkDuRVMnkddilA3CQwKVdzWje/oswJV8lO2Ja2V2ZRjhANUn
rEtK+MfFHxquCfM72QIZlNSQsCs5qhfFcikI2YH5nUB/Xacyas0IKnIdWVspd4tw
MVHAbUbHiz9MJM1+EaWkhnyMJ5DpplyNZ3YYpPN6X9pYNZIpwFeP1YD1JApdtQ7G
Cb7ksSObGJYL/NnzkjcC/eEsH2o7vWwVf9rZfHU25cDE8xTU66vWcEUsfeuLjC2u
kJ88AX7ngkM4unF/KJaWcvuIIdTxY0mgv6HvBlWKvKB60z1kYA93sFsjyakUARd5
EFXh1WjVNalqOVB+qKOaDjS8yTVQc63tJlbf0Q4bo13sCe2llupBWXjQKaOg9103
AuMsDyg/akD0LNn055zFj0jfFZ5dfoNY4IRPwAug3bRtGMPGu8enJ6U0kvQEssS4
gJf+GmozNHP13T5i8e77u1d4pp3jhwkYiX/3Z5/h0jNj7+3dZoDigXg/0KICH1W0
4gh08aK7zIPQvPe/xOaso03e8Y490ndv0gw8pdEN0T0ACEtF+ZF3WmdmOTmnkcsz
SkPMsmrUi8L3uV0PlTM4pIvmYGmwz9yfVDrnA+LKYWilwhDI+X+SoKjSha6AXrqw
uIwSwvxo32CoqA/E294vyUToog+0dvNAJA4m5gOKLmV48NTpsiT1t6s4MXLzCt0m
uOkOgul0VToEX2213D8c7SZS89qr7Xymv1nxDrZk0NSxJ+fw/ElJjIQJ+IA4eBRq
i6xNOva9kwEDUHD5kZk1jjEShkmrCsw6+vBgj0auypdZI7clNp+vh6CYW4lU/DjK
RYTDoXnFwTp+PPYRM34eHZM6Vj+SZrn23KEn9ipT6uMSwqQMjrWGE4j/QbxjC4vX
xFrPmU3vUGegQ1+hXWPrApkXkr+y62G06fzy2tPz9rrgvkx5b9ISI5e445wFsNyv
qWY9b7z5IFfSKmIpQF8H4H2lgZSojTeyFsc3QBnGLHJ4OwxSuzbN6p6IwuN8A7yr
8bbOW9fF1XCo0SoMlpzWlHWIW/rXV31Vuvo9QhDuNlrYtPJ3MB84lUDPXZo+rvf0
9dOPVCpCdjFoH2FVH3D1yuA5xoyzXp27Gib5przevy7Fkggt7eS/3uXRKM5mmT2S
7WE0zLT3Acn5kABN9AOPuDk/ixwCx6JganMMCutLnACI3d6mYtpybUi1Qv3z8EVE
wVKx4bVsW6hB/dbU5QsQyBcayookVT4ZkbiXhoHPR/k4Z8Kx5IAI40M9stZMNcFy
fo9O+xSZTtCKetlgoJyJ7r7x5+bzBt042GBTxXw93zaGTOF19mMjDeqhTy0oU7no
RHXCkRo06N1DzfWCsqvEtnSXdIHJpv84o4oJlzZqADPL1xBqxzxotqkgfNPchSAC
jOsBAcQ4A9h+48DC1nUtd7wo4wglcysGgghxFExh/LtY2MbMmVIOMyvXc17rACIB
Tqe+8eCyenIB56uOIxwelClDH4kwgnGyocvga85cRKZ0Zt4MXajyb6NTxVc/aPBf
TV7HzjYfUzVXANfRvAtnOEphmc8irDXVq9U2aAGBrxci2/YOri10+rLm9R/XsPkj
vB+oCkmHbIGy/tct10YvP5d1RFJ5vzPFawM9wRgyH75ULvxT1PnnZVZNgP2iS5Yp
Jn4RTtdoGhymd52UJ9C5UkaFteRdkCXfaz5nsAz5Jr/b3AO/kEEkKCncwR4g823e
cPSegg0XogU9ve1X665XAATnE2J0pbGBcDIh44IVt0CWoi4qxhU+8FKJKkig0Q/t
3R8jDrCkuqxPmz7IVpvi3dOvuvDARsUwzO38vKEtE8Etmez/txylI8zNfIkrIe9h
9fEgIa7viQx+UYaO2iWqr+F7PJvPQKtB3wDncyqD6mE8kIjG8oWpCWKejgPgYjUN
2hiRNtrpnO4xd7p7kszJlyPlBfosZSZPVKDW8Vm+PAj59MuXUVXCUlw2oKfifs70
cfO/tCAOLZVqBLcOeX66tX/zRLNfjz14GHZB+hnGC/hysO6KAbozckX113VtNRgX
BsnDCLEyBCNJiC0R+Dm8JmMnRgkWNEGtySfUMHewjjQ/9su8k/Qfoxex/aRFhJp6
UtmS61hQaJ0AiREItIhiJ8qGj7r1E2cBJxxYaIG4vjup+08elG9wtI6t5hli/rxE
VHmXUsyfDN25/xilMXftR3zdvrLMtbJurUvwVdHe08v0xW24rOIqW6UeyWLkX9Hv
psUYQJGgjhDbJqzx+qnC/OM6hOGAAX6WzRHJ3ncnNsdbG+d6Te5/qZgLEYeD560a
tdsVmm5HPQMmnYXOQlny/COXtnPfIo2Degvew/AmJR4X7NbBtHEpIL6n7BVTNmah
PTtFNlY1huFSSSXhQyXyr4iDY28+woioDzViemgUYWvPjWhIlddhzfdDcvIr155a
otI65LxciXXVzH7Tm1ufm2CoahvG22HVC9hSKYDLaFfcFpGjgnhibm6I3g7nZhAp
OrO+CTiH75pXEmctjDdJW/a+aJaLnpxLQqXVfi+M6Objdz+y9dWCHEV7/aPau7gO
QRRg/YWtQlfXVZP3KFd0vNWDLJphfZnypFNINYeTM9kQI+edG9ZnpU/dJdUXAttA
6h8zQfiAhUiymp+Mhjae+hBSbFABoDmQC5d5J2bPlIIvWxk2WOvPBjcVMRRejK5b
eT2h8EdKQbavmsoEEuCfDGDkwPhW2X8iTmUA/Ir04GK0os64eDej+w1I/LHl+B64
VXT5bUWp7qRqyFfbHzUXCfYSalcBcD1/If+3SlN7RK7i3NzVMyCs/7ZGbuMNUNVD
wGplQ8HD5vhcf+z3DAKCGs1p7JT/34Wz/TVPBd6w6Vlv5HhER8G7I4Cb8bdvFPzg
AJ+HchLeYNBSIn79VY2J3prjptDGia/ebEjyJcbAhl+t2mbkV42Zqdt3Ds12gEPd
CoBICP06zE+xak5LRLS5QPtcXDzVPu82svK2BaJpV3v1gJXPTcDk5n5JgedDfQFA
nRYfScfJXHC3pT9BPx5inGNBK9mDt6msgoZ5XN4yxQaD+OC6lVcpJ5FXvmZ/CkjL
H/+VwTCGcYdYMQrX7xGwN5e1O/0SfHFA+FPC9SckwPAl7ld2woDY5+uCwfs7fGrJ
0900tTX9YoQbPh+RX6E3yibbBYaGLUFfx2uLRnGi25HfdfwEVTH8QLX2Hs7tcy4x
0yLzvn9+7D3Mdif4iF8ASkg6cvCEegUcpxErfiYt0/fLPk50XJU0IOC1BkkkmsFy
qpfF24tmYVNpoJvKagyyspoo8fooE+umNJUtb3+7B+caWsQCuHzZ621GDdYfx268
Wqrj0tMW/UGGBilWFo2RFKsQZhCmxOMGWoeNPTSiaRnrA/BY8elN4Mww3bxtRx4B
gNf2WWjtB9fpNcQ5MPTTaC+dcyCkAk8BtOQ2BNM/k7CkmMu2TpT4G/AuJ+Ls/i4N
fw+vfKKG5pNBFgDvvQVd4oK3soFRhGbmv3agM7YtAF5n/75CLAfBw4nDBJDTrB4v
0N7Nlqr9+zGl4iXUxzkhcgXDhV8G2VFyYGys1eD0PYaAE1+j6qs85yFtFhQNphDX
62+QVVMyNbwX8qv6BPFZmYKsmTmWBeT56qjq0GGQgnW1p7QVbME2X4aUTGuQ62vl
Gn+FdMAAP3ps96pXODI9SAoyeh1xCIpMbfzoP2tNhh5S0Dg8MZh7txJ92zqqzzHY
78I8ePafB0nB71dzPH0VPW6K/kFbtD46dU5axpuonUZDBjwPSOKLDXaxmlgARqdj
C9nNrFflNlcIh3UkUbKOjZ1DoXiqX/p2UBQEo2UiUv9oPPK0WiEghHxYoYwbvv2N
2rxSmjm5lluTLKtk0BzV/KG/pdV9xC8pClD3RE01cYDKwSBrKFSuMOsiX/OTp3I0
IiII5XuWYhWLhZIsAxhlw+Q6m2JDtkl85Ihb3srKlUiOAoxEjfFucadpJfGvHuK7
HyDuP4hUITnwczyw03VtSXkN1L1VmwN7fTcTAKpmRQQT0iWO6jY1Rojw3YsaNoVP
5EV185hwKQRDCHz1Ts44xPMAEvfp3++sYfDJITCNosSDQsnr4wHcdyXoDaJW8SJ9
XkIANGDtI+l2Z3KPMgHn8C/mBlltKygLW6JWdXuw9+PhPXyZmjc0DlOJ4jHGVxyU
NIMftZQH4I7p1swxHzYuZ+wkj6zblHjQye+MCjTsGGu/xkkSELxrWa0q+nE8gM3T
jCQNt06ex72b57qWl+KCzNDkci8b8u523Ms1otNLD1t02B+kkcoNLQSOdmTFkc48
eZyEs26jdcn99gVUY9kAvsiyN6eeZjrp4wDOyML+guCFPowbsjG52t31pOdI/47t
p0E2XyRwhWR+zc0F74Q81MkkGowm0A2Cl0DXwiwcrBd+GTmxelZ1haJa/mXUj+Xr
Wu8d9p4V6w4ZLdXY94DtJwYtgafxZbqT/Sl6UHlKOvRZl5FgZU2JJHxin4nnDjbX
JwCV3Dz88E7xXukUn3HNbtnYkpIsyAwYG3kRE2kTV3ofmy1twD8wnNWx08+3c02k
6R7VasIAOH9pswBY5dXFI+OB0pFax3WXb/ZDZ5y5pX5WDXWNMl3RICpT66mg+WSV
fajAdPqPtDf7/ZHGesx5WHILAJrf7LfH4EZKQX13NBItwuvqkWijSJ9boBWrdZH8
wo9JggRLo2zwy2AezbBhc0UkVOhOuonP/AXT58H3UU622ReO5oe/zUJ2XJ/oU8NB
kkplye0lGZ77IzikmqADXRcNtkZsbKAbNOx5ZMaId0iUPSsf269pRFaaa/o6S2qi
xrB5DC1b8rBM++aO7krhyoW1W/DkrtvBH3yZf++x985V6k8cKGHx+MuFwoubxghw
IsuuzoAiIQBfel1GlvDRY3APfzVEpr2jWgOoPyVViqKPIXaPCx6LATe5v+63dNb/
zzYHnqup7gTpgEy1s/uM1BjiTc6HpcW9HjESxec74oK9L96iWwhG7kBgwZ8wMg4k
oFd3TgJe5x/4z6APchdycK23l7DgcQL9GR5H5d1xbII8Gdzyg1sWv++xxadI+cXD
px/BLIBKTOYUnJmzsL0/F33JMLIEsHet0opRrGMsa0i6hpqSKSHAe++9KyL1mcC/
wG59+Sl5BuvfovNqDaL+XfYbqetB+IPoO/oa/f2SQJe5iNFXt+5QQbNa4hmt1f1p
BVwHrWuVn0mFgRho+1RiVqkjzTO6QNUzrBtYC2f5v/r1h/TAmQYOEUuk7ylVhjTF
0MVn6O9jBrZYKwk+gqV8Kp1xruFysIVBM4qi1JZhlpyxJqJGOObDouiDuhCg1G4C
M+XJbmD83WbOb8b/unqlXSjihMqHTSO5IgXHzLOJm3etyMNeBgyY+bY/ymzzqdvr
6Ga5WCt5JHBgnaON1/dA4yxB5TvdYLVUuVeb5kaQZfP/49v3eWsfV125LFuK8vZq
88cYD1a6hjfQOPFm4GgNGrJCDtVMmHsMwN5Rp8xBA6RjwtWChVPJee56NfaH+fLT
FX7bBQT54xI6wkoMbYCshX6gLZAGfAjI2ZbpngKoLWez6b87RMRnJx2XhyMBfJ11
MRO9zZWmrB8DPILDefOxIzPeJenkuy9wx6bB075TJVx3y2+mTneX2WcZu+z1m5Xs
X5moYlo/jFvS/WMlDx8WU5rtzmPD9wmQ6422GbZGsh9PrH5Xv8RqADUQ+peBlzHG
Qt/eT4wC7oIvdnPVAH25B0EKYqDvg6WHPcZ7aumorytJc4bZaUvIr2lHimQ/1pWN
Xw6Y5I6D6T4zLn/5hTNmjj7x9gXdp2MFLCQhDDMIMa6Sj15N0d5bLHy4GS7aPWiJ
xXIWORywfCFTBR1Uz2fgxxteQIUAjr9j9+UhXaMVBhVnJ98+KIr/iDnbcWp9JgKa
GDPNwz4TfpPccfvQ4Ucjq268zZxcfZmvfGJ70XQMxy4DfsuwH3MVc9BnkQCRvv93
qiOHMv+dQTXQV+2267OHQec0EeGt4SQZs+azEPdMGf/7zTzsXfG8Q7gfd5xXsGEn
QtNz7Tj7mrbg9SyO5Cfuy0sZl7Hac4SFGIHHWICeA+Ukup4qnAChBKgInWe3rUEx
O7S4hsmr6qq9TGh9z01xJfO/UUiULFhxMrGoYVrY2899s+zVyDvPkwzmVVfUBil+
LnoI5cXlwJunPenqVH8DCnwSiZX1Y3EtNNXrbue9CyCblOSUveo3r+M6FOHoenoR
01TLvWshwfnTO1Z+O8V57nolUdpczxI/IWtZnNcF81MiPLp/JAjjFN0koNMZBdY5
+0h806gZ5Zous8ibSZ5tWXn7x/HG9Rwl7Keun7B6RJTmHkQIxayrZaYnd3rD3QXL
NUF4lZcPl5kuoKWgpTXk8jOAbFxUtRwuDCsawiAQo56N6bOVzvZcIuSR0STNxxuT
EoD1IJgoAD9+F5YkFZfVEducLCDOF5YTRHJzQgAiy+VF4OR+jiKq06ZoJpR7lvkW
Ef2Z76zrXqeum3hmbU6/1ooOfnG+mfVGi76IQnX41HBl4gs9m7qMwROS9+0z65mQ
OjYxYb7sHnTinzQP1v+DgQ8xGtJN2tZbnJiyVzr6rs0oex+fmfDA+VtuPZ8gpOoI
sGmmuvWj9yL5bMos+5VN61mT/rF+k8c3sf4UTGUL2ZoUY0zX3duqStabsE2EK0nx
/bVpU61Q9mdnjPzoDnzdukZYbCweJ5/PX3c0auOm/thkITG2w68mVQljOfH7OH05
szJcWogL4JIdcbjXSVqihzLRy/LL6ih4m3QRXQZjsSRlG5G+XZxvemfVxY4PWRGt
+eT8NfIyfSaGzsHqutnDXUN/EtwJZlSoyUGy2Xr1Om8C1oXiyWsWnbpMwyseHPgU
3ytZakAtQmZYYyE3TktbnqRvs2u1KA5VWQMRP0hcwTjkj8lR+Z+mVIFoGMPImUL6
dIyyvc8NH/Bxm4dwibCDI9a8ixkDG2GxPJtxooDjaiJcY6wXg6NgQgYSzsTA3lLJ
cMg0u0QR8dr3vBLFsVcTlfgRYUy/M4+FpXrSB3IebIo6Xya1kSLvKzSknpMQSM7L
cYCKY+eDBtwkz3Z1hijufgZQkfeoyj5marPI0CDWqolqneUcW8tdKGt9tqyo3pKV
DVcH3rcxUmUsFgE0rBp8s/l1NERf2oKFq7ivIolPRjWacKa2Eumpky8bHtKeBhmH
26oexad6hyOF9+y1ghNauUEvS/p42WFoyzGDnZhl9LmWZe96tSBtnfhHu9AxvY87
/Tki6idVJ2HaDua37i4JdzsOxKiQKhBkJIYeqIJ1qO0zkLusDtoYxWsVWyYuixQf
Yod21qvUOntOJBNxSY4WXW3Dl5O1moqw54P6NX8T8uBAAo7Sf9Ku6GGVTpX1V4eS
6X76bIMRzxPHQeYwpDMyM/22N1o+kexmlSHqOEel1UiouT9gpimkm0JQGupE8LS3
nh+adUurqMIN0SWVrrXEbNhDsFU+GOHYz4anPpNn3HUQqrFvYGJK3SgPl+yVWn/G
BMjToR31bzPabs2zhMsw1JcXzniY3NZCai89fyl0v4IH/xC/RDhJmGIx6NIdgurv
0RaqCP4CTYF9RejgZUE1Du5vcZB/23vCj48+hPxUeZGSHlFXKdnzmXaX9lFrfnO8
bM8FNyU9ZopRkvMzkgLNi2Hju0z57282oSpM9XD79oK+/4obBNSYsETxJyJFEwNp
phwFD/3zh+n+eHN4u0dlKdzW/oqsUpscSmkdRLK/n6XtN1uXffkiSCAAfNpbTg4H
Uk7llmI247CUOVzRKg8fZvWm8MuEp++M658zg9tpg1pAEviWQ1uKK4YWOTNioMoY
TNWr9mFacEb182wCtttgbSmZJQmNMzQgZQdl2uaCmeAXRkZiIzDkPEn0q5cLBNFo
vJZT0ruZGtyEDm2EMQFLlgAxXiSNlO58mibYsTSxXnBVGg+pvuKu2yu7nYCap+Nt
IdFsr9kwZCylzAsWzRZLlpEofjBEuqFWc5+9yEQUCPTevRuRW/vsegNjPOd1Me/I
nVyE/EHHchOM3i2j1+X+sbVgDZDsPN0L+irkMyKHdbtqIDF09/Uya6sOAxlXaHPr
ZQsyfhJ2it78/zcYwo2eSnAC6/v+Dn2GBf8Y1WLrBs04ICeHi9R60XjlR3F1VlWh
lUvKowiQn8YSXxTJtrzxMLLfqWLopBtMuqW91DSaVO0Ew44c32pp/1P50lzTqu3b
JH5iGOLMQUwcPKLJBxnd2d15klPntuHVPHzqWYzUA5BNUyYRiYcQoaX6a+Izoj/G
XMMPkHr7PJ5OWTHylNUS3rFvadJpHxx5XRHIYSFYo97kEx5WxG6XiPxo5z8cQcNF
vGCj8MTn7xgP7B7w5Q1+1qaVJFlFhUdUzLqHR6GLc7uFdrl+g1FkndKw7DRaJBeh
SLnhSRz4GW650NHt2uqWu/ZuGLS7tunCe69Z3J02uP6/Vw/j/A83e8oxGdvUSrzG
GbC+H1yMMzQm4rthQAvSlEuntJcVQQuKjPFaTcPnbjlYGcZSfHseg4BCQKyj9GOM
YmxLMGKVHCaigQ4QG4p5848bBS2SDFdAUvb2DuxKjFxWFlxENWZQlFyzWVe3K7rZ
V8M2CD3NUlgZcpzKHsJvzm+PDMiOqZ8GDM/Ns21Pw9DriaT50GQjYf8rojd913AJ
GZaaH+maDj2x8oUnq6NCur40azygqQv6QGtRDeFIfgXYhnEEv9x0DepH0BWVE3pA
8wDShYKfKyqgr4Tb5pIsasVlkMVICB1cxot7MWwFUFldZridQNvpINgPzrxbBgyP
tMyxQ4WnY9nnsVGrm9PXDNT9t/vfKZG1vXyukJ6BLcdbAJmd+Z40Hdg2k2t826pF
WZz5AsBS7Q2c9anv8yk7kk1ojo3eDSi1P237L10i2UbJ8Bn+c567norHtxtlL9Pi
+hyYJC4wmzc2WrNMT5QUeMdKTyZbJHWsMiBjjwuLePP1ZTcCGifa+391Jm2Qgpkr
4bIiHOh5FeKl04GVT/mnRRfwdfuAjLkR6fHd9YBw2UCn7C7S49U2gL/VD9B74VpT
ePOj/1gB4yG+mbKg1wBmI89dsy8mafU+JYdpsCwYfYQ8Mz7odXb8RjIYVBpUjl9F
AOV+M1/XwW/9ApbPh3neJfi9TYD4bnbXxd/nAzwstT4+muFVlIKiIVj7IENy1fE0
SZYgdCmmomOewIwU1jTotXNl76p4Zy66dpVOEzgq+EVXX4qb8mYWQDr9l0hF9c2l
cGw3wjy04IcgQ0Un8aDSxuyUw3mrrU4WUqNGkPxTuXV6oPqcpIXGeekE2tx7WLiN
WKG91BpEtv/FmbybMtuoYui/jvtvywb/9W/78f+SV/yHGBjkcN0sHggw8BBYD6MS
9AI11TNI7JJse0gjKghEsyVI2iLn8HJVhqkRIm6OA014dvZxWE9Wo6G2cYj7US3u
je1ZPaenMLZs9WdVWmZazqPaUJKBATkbGF4OAw1b64X2/+sYxVbOV5lfSapFAVW8
2ZRtNBjR57pDmh3GRhsEpyY7F10+AQYrkWAfCRt44TRbCtxSAAOE0WtDYi2IJ3J+
k9gf3tCEvg8iim9soTog3DltXhiAhWQ08kYLTYdfduWwCrQEBxOuMTiCdosQnUm2
PVFgdkIaQ0EezSQyB3tmzkWeDj7UmH61NdOiEhfmnkjo5tAy+iJmbiwka0buiaQh
nQfza1O2ngyxmV8NQQJZM06xgwoAAR0nrqknhxNhljKkxr7mYta5SUaNdKcxB5Go
gzMZdINg7m/P64jq0PBJTqHHWC56MPg1mxT2Fe02GcOZTetpBsQLXxuoI4iV64IC
U7RE/Yu9gq24kiEjZXfxxSKTtKuKpxLFndRV56PgFU6YxDPcJYg3HBBeIFtjenfW
fzx/okW32Bg9uoXyxiB4guTuyneBsy9qXS+woyUcivlk7YZh+QFSIDV3daWWRELH
91ytoFMY8FW5aeb3L/0CVKhYm8kot7lZNC9BLBT3J4jzEmtsrzrzec5v8yuBnbZQ
kBFGO7aXfVLG/hB0K43RrQxPdzJsxzr9i14f8gn9pAuAbWe9nytPy0NiRpRAPdB8
0eUeAjlrHBX+cXA7Hpomkg2YxJAhbxlYxWumAfKoVg8mObWtX4c0vhtObzV9aIgK
3/qv2Qk2Q+/Mh3xgpvDjYjVlMOR+Xsagp2/I3vqK82GHUzXws+ZIizffmymy0+lw
yWbw4p9eTxfHIwkkk6T1AG42lqJUinnYvXS38nRK14ulGRkdM6VbzIz+wV9j8euK
M53EGc+5mvag/itCDpspZdugAmryky7RXb4LllSF7EkWAxmNBZTKLPVBqBMc7mWL
MtSe7OmT4ziIAGU9W76OG7HOgRSBpAgB2vGbwCZ/NBvXH7qRbrxOOVFSumM1/tY0
4AtUEsHbqkPnGcX9gB0pRxk7EyRBPYBELQyRVFQjt2cOAJOeskX0bZzeVyc+ZNVB
BSO8AwwwmHOJbbONt3Kbyf/haLv9GbdInV4ihnltrKUIAWT8X5xz57X5e/7A4Llm
PqBs9NNrpJbHz0ZeKW+6ZgOdcWUuEJ1nF6wAGR7650AC7Tm8m0TZMc5ACPWz4J7E
RU7/d5rp8Q8W8aAGBK9WRpdMxDxah5zPM1h0M0sB0Mwu6GmaFRqfhqvi3vsA/oLY
ZbN8OeuBt7LR7n2PJ78C5Gx3pw/Jquh89iabsa68yiRn65YABmZp5CjSkqGfo5EV
OmvjRzcfW0JTD44fM3fDl5m/W3gEQfT+gsrivSK1GTtFXXLz68PFj2b6ol4SyN+7
zxrIkAtmJLG9862HtEWFvoEXhvGnM3A2a9slhiO2+W5ab6ErbRh/0JOlPyifxdB+
tatXUY0N0K6GFHlayn5m+qebSt+RRFb08sTkHJ2y5fG8Trf1aUEIZXckwazCMxLr
vg5y5n58OO/t2ptEi60GF4V2A0rmkRaM++EOvuhBrYiEwMDPbgoBIegaZ/JAYh0s
t/vfvyBWV5j3tx78wwGDK4HDv8th9dcJcQuhoccr99XuAanFfPSuKriBjhzTbiAI
FQO4FVmFL9IS2u0KSkuTrxkZdZ5GwtiWyv4IkZagpFEZ+m0X3GKqN+gnZJmPXHIT
STNdaX5lWqbjDYP+q9Uv6FWvAzmEiNBgmttDXG3OCvrnUSAo6pc4EJVbGmDsLa7b
QUJehOuOSF1xx0yU/1Y2GSqxPjTucsFk+DlShqp4L/4XQ5sX0g6LVaRHJLRDiSQI
43dz4lBx0N6hWVjP/9P+ozkR9N97vAqm35c/1tlOSpIXhfgfnjoLlxjdycApkbfQ
opp2OB6uDRPrg6QYI3K6mPwy0CcpfRbwFdKQlVO7CnlG3tqgCLAj/fBNBKsAnbHD
sX5mHTSX64WQC1PvaCEPjogfgYCyEa08BKGgTtiYp53QvjrLz6pGmC3w7y8pptug
+7CCOYmqsgpw+qpVL/y+6M3CXT2FdPjZsA4Tt4ZaDmVME2s8ur0P5sMhIupRYcDN
3baYEoQsMyLH5y49ED8URk7HiL3+cg+Vi6pn00nEg5MOqWS7dOk1+iyFl6G4ncyd
PVvULsSoiMVA2ARE6rvb+DZVz2EGxZs3QHwRbXyiFtYn24yuN5+tAqZQVG6r3Bns
4kQ9ZMI752T2D+10CPrQUe9vgMSXtSkMCOm41Z2FW6jb3lX471SrflcWvkYCaj+D
GA1vMaux347WYsZ9Ad1gbbQujRqD4hrn6Rz3IEtFr7puDvgJxsoGlKEu9gO4/Brg
/aGE0d8ZqSqGa2fK8sc94KcGJ1HObqqAvu1Dp1DfeewSnimxQaLkLqzBwr+wpxJg
tB8BN/L8Q2F9UvEsmmGHjmdFDxeSy9sr20DSipNMm6f50oFDPiE1mUUa4f1qHqAd
AakR5LqLyAagyxBOFw9FwxxpCx1/T/QpFNRteu6H1s6k0nqG1LPLpFIgEDd4NSn+
RHF5+izbxAhDOnx0B6Bs51+ZWU64clX90k4/INxQTDuDcp9saohcYsq3B+h2aP6G
S9lupPyz8mNJOwzT3d4KnPTaDh982plFS5D3m/1RcHQkIqD6h09TQxiltL2nf2qA
RTj7Sg/Dd6QC7xMePF3YCxS2FhOjZPi2w1EPdm0Mc2t6LlVqq3MXCIzCKCozM+8L
8yVib6B6N6tgCqUFz6NA99ZccGXUc/wxRTVFUsN/BFawHmYzKmLR4qYU5NDUrTow
IKrtVGALQwMzNBmxTUDllmk/gWSua0e/2soEDXGvgUXMf0IJdHoIo53WfiP7TaTa
Wk4DveKK7gYOI9A3D5zq1jNHq/oxpJ3IlFbVru47lLk477YHl+K2vx1Cwyy2lqni
Jm9TYGd0iUYLbSrH0dl8xGfGIUFVL0G3BJisKseQ8f4taohdfDDy9G6RLuEBOUkD
InZYr8PJRwA+8Y4T9JwX63VynxsMVyOh/w/tfHXCLQGmiz6kOaOMLPXUn83Q2biy
eZO/ub/Tclol9M8GyjGuBaFJicz22yVLu8djfrfwZzCDCT3PVwQ27OGrdTNpvJAM
e10lfErUrw4tsClHhNeFhJ9LeNM2B1TiEjfbSWwbF3dZCZ66u+fm3AX0herT/dT+
g2gIjb+nwQFh8qRvDqx1Q2wwGr2pkIPD21F8iAtC/vA0L1XRt+WoXplA2HZGVJUo
a9UvRwKBcYwqukBAiTUpnrONfZqQHXORZgiDRrtfzZgeoS01ZHU2bt+lI/mCP7aR
lWiKMWdXd7KQCh8zKATVGDWDokQR5FcVNnbEX8skaiX3Aro1l6jOF79TS1fNVUdI
5uLwewDk7Mdn2IkFFeB0LoD46tv3ulZ7xgs44O2sw6c7Fo4rjVcR65OFgIAuhIf1
lk94qlJFA21Ux6hjwe9qid5OB8RzSjiGpWYwL3Z9+v5163M3AW9IGgE4fuwK3o6y
TIsb0YkpGQReEBiE35pW2tXcZ7W79WZqMmgyQZItUSFi3HjIu+Erq8Z2PgowpTDf
apaxlx9k74IKyh3JPDzHKmsdsEIqpobaAYs82pOOTyZcSBhG6o1LXRy5qHvRIzAP
viXQgZN8G4KS2WL66CuO3J/lAIi1UHgb1ls5gdgI8sAsrdb1qlFqdxz7eLWmZywW
4o/l1NKTNn20iL3BXJ0JiNZe6dwSzxWy1lebf0Rdul9EcAPT3yuBsoCYFxQ5ZJwQ
2dwCXS/cio6SxvX2NFr5oJrEcUFHEIcX0LIuiglJstEatrKtBR1AwQgfo825pWAZ
NIkBF0P3N/p9UlqA4zIZHrLJtE0rXCCRga7XZwU/UaTkGWEbKQ/wuA6KVx5VISIs
bo4iPuCsv/IH1dqLmXkz/Mwf7qLPu/1pgbtcAw0hgDgEqKLaROYyg9lIFDxqplDG
F9dLMtiSJ7UOeyMCwAGVFp0/3CqCJ42n2iNHZlWSb4vjljZbP9YzqUS/9J0ypNvK
QA8Z2g8kd2k9kV3j8IJLre6/LuFYJJeAbWcXRByDfwt8F5O6J9W0Plfph8hCPsKB
7Zfjrpq9Wd3LWp7E2+F3MZ5K+9Oj1Y+1IfpUl5HXcHhQk+JeDUy5Uuv9UwWeryEQ
L2pN7+WSpE91GjNxj4ADSBCDGDDYtNqAaORpeIjM5ClHdDQ3Vj7oeids0TrE3GFP
yvNLOlESvujIdm43sc7uqSkPtYtKJ5BZW4EWng0wRyZqz9vGIpHjPlHW822qzdik
KbrkYbdVXhs0kCQU0+QH1RlHD+kXw2XjlUVIQ/WIcZCK2imj7tTPk2l9CWNTIf0u
ZKzMfEfSOb7+yJO1fQuN/FqeTCrBVx73mKFECcMZwZUq4CgPF/d3l1OcsufhiNo8
uVD+b3rFjtnFgtpR2ZKHvMTaoxZ4JthGpZaY4o7OfAfGXMMJLR/Ivq5Qd71r4sNA
kogqeatd+YHXEH9Mkhsfp8v8O84YwS7TqIrK/YP7Y82qiWf7VFO79ja6pylw7LZp
qSn7vN+Y5bn9XaiLetff2XTuO6/+w2164jBlkiZkNtsE63sFU/UuIUDbhoRetmHn
xGyTYVMYGBi+QnNtZ/nqDn9uqsahcSCLKvdPTGxTtX+JctYxzO7451/michwe2vH
o3TE57xg3Ej2P7K+GF0CnDnr6z/+jnMD3M3UOHTDrg7T/nnGWhk9anoVVFdcK+Wz
pBHqkeIxLo6wnQ0sWDnLBBjbgGMqzt4gNrE6IPE6qYUjtIcjubh2IgjU7D9oxaSl
chc3qajiig30qythzMWp8Dw7UlhUiPJh4lrGb6t/CBtLhp6XQaCd25Xg5JAIESDv
uYk4KZkq/eVccCEBCR500PyHR9HpaOGnK5JeT6T4C6wNOcabjjsoIoVjY5qadCsx
g0GYtJ1bPcKmwifZIMeYcCQVX6waRjUPxnYenSiW3QwFlo5Qeonq/We4b0X6hXg+
BLjEXK+M3c2NnmSNNniDqhbr2a2SzS5cB50H+qFg2fh+xxkoz7CEKUs5VEeTAmMg
GVmLTKXIfjt8McZrDsm5Z0r/t/7fKgtrz3mGi65uAi7FUhyOUDLta7c1Bw8XhBHF
Aoqr09W9i12mbtPqRFTNy+fRZuoztRqJu5setWP112dOHWv0a3rPmeeboCpMTE7o
0NnQRujVWfX5I/cGdHirXNFAOZmZ+NJmhsw9MfLQGLhd2cuBjp9TSKliQUEOe7hP
Ju5hyPfEnW8s24CGMn6H425AQNZ8t9iAV9ULXIQFDvGLP8lh0X7Hk16QL9VxlCeG
/EV0kFYhz/dIVejsL4kCf1f9dGTOpgDscoxD2UtL4AhOjxQ2sGEsw/7Zacvh/lPS
Jei94PiQngSnyqRubfDFK1jiraT+zAp7YeCUcxsp1Wut193EtZY7BcVTY6YhYMxp
wU+ip+mT59c9iIib9hP7CCYP4yqKTA7Oy+JRxtWt0tRpQ2N0vgvwnmzx64M5waei
cWKGzPtorNyPR/i8e6/fi1OBVcsWlPImlzANz9EhiTVRw8d+ZVMTuK4VvJvl/jjM
1/z7NWuEzcNxmKnrF0c3mO34o98YjmNF6WlYvS514rTTNi6UKLHSpj+UnLiCQcVy
rOQfjgNR9GLx3hSCes6pqCZsGOdBwUNtIUrGBoX00CEi1qdO5qFnQuD/MEZs4MdJ
5WVHubeCQJTRedZWPY49Em9yOwz/4Rp4zdMkHMUMd9g5NY0JvRXd+rnu1qUCjzGl
uZVN66sd4luhq1lFU3qPuK84rMrPlcXpPHf3JMfkW4+Pm6wcvDiPtkUw5+/81Jk5
9yQSpaLBZ+x1fcXUiNbqSTopx0bWvwzW4/1BJ2GhVjUamPcPXdDs69bgGW55qBdW
GNr2ot30157KfFe9mzy/MvQJMfYVyEMkRenKK/dkuHBml4OKKKeT+mb/ig8qBNKT
YtDQoia5REdYvs8Agjjd5PzaDiQ+7Ui1nj8OWcPzYT9AhxYJ7bS8eenSzMfjceLo
v1QG8M+gbgtSrpc72ZfDX1F/HmnTuiZhQpSwi0slt7485esLx2ogWGqEVjqY77SI
oW9YRlZhfElP8TirHGN6rlsUj1usRi10Hd1+ATdyFdWAvUtxkdySgVeWb7TA/rek
zMl+RW0HIKwbTN9rBFfmb4Zl2gd5m7+VHeZm8LDcEyJDjIbOlCTTTc4yjeOrc3Al
WeNkpPUj8IG8qB+4Eqoj8x7aNWFh0yC6AQZIRMSnfg47reLEZ0hTnm4h7Pat1MSY
O+b9JdXtn5+PrWs5DbwEhyU2INPCAykvZ1yi+tvMoayULRR6oQ+RKctqP/a9ot9B
LoK62vJvqQq1pBc72pKdqNouE5ftdMuF9yLmEv159+XrEkj0fL7oplk2Yz/OoO5U
u4/wTniZQymGl1rSWTmPrk9955okviqae5LKoD3zylFWOGd8sMpUBJ3wJVyJx87K
LWWpKpgVRLhF1dhXfdagshl64yOGxDWPP8f91r+p41DWHybUUoKz+O04rJi2EtZj
+bBRgBXCm2ZN80YhYiN2Hkjfx6ktBhN0Uo2DlvcQL8VCFKW8QYthEYBHRp4Kz1YB
biv2mAJj8odFXMGQOftoc5X++uZGj50CV/16sDgPwjhvP32/3m6Vw3Lc0ddHDzyl
fASeprrKXSHVx/EPcu7c4lIQNQG4ryvX8mocFerwdlckBG0sbyjqj8eKIA09h4WP
f7JZ1+cwvOY317R8YtqQy8vOxAOvJXbKsPI+dwK9NwLjCdLGh49tyKk8rF4vNAVT
wrjFugRWCf65ffieyNWL8YGQqDep1KPjL7Upz/Zp6KlzmgJzr1P2wWUbLIZg8u99
80K75rUrM7wDfJDeKk7Qkh4Oexa/D8gT513MQNh1mloKQP6iKoXht5U8T8xMBvZ0
dYjf8584D6XSJ6Dmoe1Z14qpJULeMsBXrv7Wcg6cpQDDpnKOs58fPAr7NB4XjAoc
0T7aseLjd7U787IGBu3/wgsmKSLwOkpJ3jE8Rm4WXivwd+djzIeP3EoPb0jD2OgF
+erEa7BMHPs/UOqE+Yt3P7dbn7jWOx5x7Byh7I6b4qEZI/7W4VISushrDsmRVY4s
nhvGsKgkdihUE6WM7q+Hk5RCYkchj0wULav/zKbnvevW2MH0EPUxnCsNPEPynzR3
brZDk2d6iag5SLAd/FUDUbN/sSmuSroXOV1uBHAWSCY8ruqOFEple/PnB9tLScFv
qIH4BVYfUXJ1wX95h+v7ElU2TXZrgcR55pZB9mVsAjoHU/EphZz1Tmqhfn2yjMJb
mqbh68J6CtxngHdej6rKDXfNJK/xdJIcidsxUsAYTr0s6tsP3Gm3tJz78xpqKIFL
jh45nxRshU2n42fEQTOKii4UtuLkJeCZifgSeffzSxZzDd+Fn/zVNWTe6HNtdBSt
TxXPxHcpumsoQnvm58ory1/rKDcG7EgnUXHUZSbwDiGJBPL/EqaSaABLTX431g6+
bpjzLl65IE4MDAWVYHpmDt4WNrndw4mYqdRyLanciRs9/S7QDtfJIB/UNLpVrhxq
U9I6fJtEsve5B8TBaeq6E77i+1vzhvk3BSnttWFtZZyrMdKg1hhkOqKVBagykXmU
m0Ok9Ux1Jp+hH6wcRaX/IxScs+7hJApnA6YXigYFITuqgYNmzsbl7ORWoOq+cNz+
nMJUeKWYG47F8elSK5PRI1zMOZ6XQHy4QZwUOuOAw5DP3XgiOPz3Ka67r+rnMSIS
QxShJeEgKEi1jRMNGkfveZzJTYYpClyH/cC4rSxA5C3BZkkNN7M1Sz68Hbcwfel7
bsh3CARVIFcPTeuGLgxCvNuKCoIvE69BrvmDgS4K1zKcodst6BmirkAoUx381YXP
BUcqVpRR5/75Yp0FE7cx+Cwny6PH35+fUNg9OiJUF2s3UEcC6dhp5DakcNgdg2ey
Iybj2RGYRGk7IBlIain0KYktSJVo5GqzssoSKvwRvsbj3KeEizyrEJbMTQd9KH2c
2jfFzAHy7xLz0iXvHxjZpsZOlEyWBaCfNjQC8ACk5bY+V+tzVwC2D+IuQ24bw2pD
DcoDtGqvM9Knm/z6K1oglJN8AjidVjV6ZlL77WzD7x6ca9M5tAr1aI1d8mBLRdkU
0whbu3I/OWdZTQkc+kmisl9xuiak4pTLtABlrszsnMZF+moBC26pOhWbBH7QicVR
zkROkwYwCp/crA4gLbU7nTqp/FSNK9aYEjBS5LRfreJxaRptgfmY6tJDDrdCd3nL
9vf7qKaiXDgPyvOnSjxUSshIQ/swGShiBLnD41yY56EFcYu8agBzCJat+Tagy3Sr
Cf/79ka8X9wJ0NeABJIr1Hco7zftbLUnWTN3nyOU38jNwZLmkKnr42WRL0tevCyt
Gl4AEG4tFB/nWdFJMr5QZjowtv7KD3ettAMeeud5UqwPgX+m5FcnQEQeDcx8EHRK
M23NeEuMwPAC+EYyy1cRaRFBeppYW0bAX5GF/nbTjxE7jkL/o3h5/xdtnR5x0VVQ
Qwxe2tWE+rHoA0ArE/MNu4eionvL4NSIODdo7FTudDu7uigjTHSmL5OnR4eJFYuy
tEHaodD393LUgRWneG5/rqaaxLap47bLi9B87n/iWvKjtGpNUru6M42INGhwpTko
9TeoAeYduVov5uRoJ1Nqr0tQ8Sib4I6unrSHaezkJYj5vahhVvaYGGJaicb9M26H
4iqaJ25MDz7RidW9tbnK5Hy3iYnG3mqHvbhH2jkCBsNTcUDU2RaaS74wu7TquYo4
DCqpqnQp1pIP1Ckrvbq9rmT4QMV8qOKsvsadXwrRbN4y/qZpn5jJBaxM93gkdk+u
CXud4js5ehi5dplpawaDhF0fimyn/S59Ch2mE+xVArIFe9nOGDkSnV2ouLN3GObF
Am35v82nnCHWkjQ0OhY3zpw6f99B8N79rVnd3KOnYpGyUQ8jJU57yW9xDt2AVSss
Qp7r/3JzvWNCJpu4qs2FjGdaaRZ0QdT09UP/+5yDExHnSJczHwOdhmwpi2aoxk9j
8ZFXQeTS4ubAkiYUU3+78nT6Ev17I6mSC7/d5OJP1jJnhxRs5JbVKo+QGwl5Cwk2
VAjeFYePkCFGmA6PJlp3oyOB8XYtRlkwnzg6jWSTFs1QF9r89jhKhSF9v0f5rlhh
Gej51htyCQPhBA+wkCfHviRGs5Ky3TuJow4bD+ENn4VtbZ9diM6ib3dTZi/6zrun
5JqhcioJDS/r85AoLsOYn3A7/TeZqdk45KhosxPYwdLegzFo8L1JwKKsJ2kTYEC+
cTKMHrwfLWFl7gN0fu1ZTNjfEPO51SEPEMLcEZ8CpOf3rXdUMmrst23CX2K4WKkT
HDGEYpQVCs5QkRWbjRlju63zsT05w3ukwb1DNPW1HJSkx+Ynu5GiuSIDzt8f458w
efXI6EGYEeBzdov+aNbR2Uw9MXduV4RGSm/j+8H1Oevupt1NhPa3WBgnaAyE1/Wu
48HKgFzWCCXQUOmE6bUQLt5mmBUNUW7pcXYWBqsGn30gUUDO0ej8oRamQTdWPNvM
MesKabw5pHhk7JtjNPwndiP2xCse6WlbwZErlo0Y9w+48yNMmhvl3AK+UX9Ws7Ln
3ldBibMJuccZV18PLLsGoESmpTqXlIVbNafIOLCzyCZmCX4rd35WemmjQWxQ62c3
Hofr3r7HZQRS7CdxKNrs2r4rZChT5GttMPrqo41llTnuZcTFudnQFxP+t76E/t8t
yxdLsm86Du4aSfIvZVcSFLVUpaltJDq+eS1WFui3dq+4n45OM+oGq9QskjrP5Hz+
/mqnNvfrbBrrjfzXlLMuvisOzfQqpS5FkCJYtW86wFFMuHn9UZnPHEZDaZSjbaJn
eq1XTimVrwQiXZNwrdAvfjHhqtt4dxi2V8IHFApttbD0GxKvokJLCirEO+Mga5gZ
z5t376qSlY+JtXFPeF3M2KDa34Ao88t3TuPiFGmbTwoNyrigYNmjhsYYrWxde8PF
dc9kpwdNYo9UXPQoaWLO1S9S1sXl9Crx1cumpM8Qvz/0dOyKWocn76K6KKP+/avB
U6jWiyTfwQfvTdx/1c4uoQtCgOzi5UgdpSpZ1ehmIKNwqqM9Pr1eWjZIVS3gNRpo
TShuRrSxdtI9drHVpgR5Bk855eMIP3k0o/eR1aBhWSWBmPIejpzGtsO71a0luchy
ZfXN1scpo8HHAeZ1PCPbtVI5aOWEw/+3UVJQAOeLQgi47vgoNQlt6uWv7oOva/ov
8Q8P387e63p/hfVW2nZbKzcy2uUOrcrSoikTdqKL9ItVYmaI8i7awC0/dI0eQtbi
m35pkD2jgvSG0BcBXYt9XjXigo6Ijfr0/l0rZ6CNrmmjMSUNEWBxQXmVrrd2e/3d
+RMzE8WKYEICp3A/KF2RyXUIVjZIejvcZsxfOQxkZz731bFE/J6uAsWYDvW5RmD1
ean+9fQVkCmhD9fb72EdT52+qpqItvzx07L74yRNoNxWp1XeCSeYsSim0its2MTB
FCrRqqAeA8jCDI7rZGAEmmKfx5ldDJ9SvHMWU6AQjs3fnEVV2eCMjQISK31PC+tq
yfolyddh2RbeW58/rouWAWp4ricWCYQwXHE25Prod/1mi9kC2QKTv4gPzEYCSehD
rpzghGni5bOk4eHQJGcHoX7qwoKusn6Kf916NYTxzn2sM1pCaPxghUTbXg1Pe0nu
OGGhIfiQRPfs+Khrt7xD/AA4MeOSZ6kcbG/QIKzs8aSG+QKfEMGkHUa6cPgYRu+9
04CanL155bBNfVx/Z63utpic+zUhhrX05TGoHSC/Ff9YvwdtBRNhTiBbsQvk70hs
9G+7cllb+OYy/S1ZQmfa3GOBpby+Jtw5JG2zRnQN631tmYP/v7KTMWTKhVu0yovt
3cBLue018O3ajh5aselWUWczZxDTlLHl82UatYUYfUiQWVfrVdpdXaU98r/UU/Ys
6kWMVjzs4U7ek0BRiUM3+6bJMEAJxvGaUdhOAjpcDfw/7aOgOlduEMXuvkk6sVr8
ew/4oZYdKt2Rz9cWddFlZDxmC7NzdxrGN+c3fKBSqS179JiU/GWlAe7idpZca7CW
MySnxoq3PWE0BpOwxD194wnBOQt9EnnotxpiUzdpfoWDE0yUnGmjugFAEbsn1zyf
SpOcfSHaH5ye2vkgdQhjAQFQ4p1cATxC3h580tNm4/rmBj91LwaicTBkHNmY7OUB
hms3DAT9W834lEgSqy/PpIlh9GCWWHkE/fz8E3vrev0wkbQrVJTybNEwCtPikMuy
I4Q3OcPbSnbUCWdAc8o6AQAg76+Wz94tu5iVBo6xHTaFyzr0pXEOrdqIbmLwjHcl
Jh7Yw+6SfFz0jf24wbsIZZWLf2j0HURRxb336AfZmCrRv+WBy46SlW62oxRVFsfe
0gh0xXNqOgt+GK+9yEOt/PEQqamxrKTq6x1KlNQfyjS2x1hvxzYMcFHg2a8x9WWH
V4gUUxqGdS4apLXgcDujDQ6C6SD0L4v0vOPNkzvoFPobOT/gZ/aiK7F1WBzN7dUO
XU0DsE3eS2c4h9WLNj2NoIMMt/MqUYIEHwXRo9wDe76zPJHW9xZybSprw6+XD1pB
CTsPr2GHu2uBXWSuOKFGjr5rrX7VribVvdjVxeCoZBuz7844z2++eTH/lLIyt0u7
arUJgFDJRrIp53keEUq/BX240fhHbwewrykBUiRg3kDaSiKiiFP3jK82eKaF9CF1
YKnE2rdYo+cdFn8/tMYJZpdCE2Gw/NZXF5qYVYBOtQsnuqYsQmwaIfjfabvmgGzP
DDgkQVM61Lajt8Os7MvAZoD+C+LHqQfIJSVRYM/EC+EPJ4Quoc2adbJsKmKCTo/f
+22Jol9Kw0l/E2Bh9ctf487r5lWncW0DquzPc19Qfnq9wTO5DGC3XjjfWGRo3dvo
5ISWUNorlHI+b7bc8/3FcRhY42DxAX5A8OLfun7i7FbDxZeSSDfagFkEEt6WT5+N
8foEOeJV3oLaAnNYYHnTYBwyZUm497x8ksPswOqVXS9sn5WMuD2xx+gY+fGMgVW0
WiUBFU1UANe0Y212abCprXfaSMrpyb3NwBNoAWQIIrRB5m8SqdehICB5WHea3gqw
57xtoDzzYCd1soOqOxYDre4Z4LCH0pdnNyzFl2hsMhAl87oV///pPsKD7MKiVrjW
pbcbxeVrFomokN2XQjVr+6mKazPxY9WkDfouwedHpHHkl6ppMAYaCYpxVHVyVRn0
rxvoYOaAkmG1MD8g+70F7YBQh7Ho9M1NfAYfg2mGnw8b5CXgaWGN4pkKR0YP4xMu
0jg3xGuI2oCs41x2jVND3qhvID89wO8cgaAOTQY1X4J8/OsLS90Pfip3zbEV+Pce
Bt0YGXZ5QUA6s9/TKexI8mFcE96AHbjqhNH5D/d7UeuP/wrMD8gigeuN/SedGcpG
GDx3wEZFZzy1Gld7okXCy6cE+aFyzWgtwBaGz0yCHxxVXnyog0ej7/R5xImr5veF
Iutnh5FMCrP89C81I7IKGNPeK72QWTjqh7ocRdwE5tF1sH/8mUoT4INCL/Bbcwx9
79ttW84RO61X8PMX0Bmu16DkdcR3rjr7BOit+1CG7LKa3gSZ3KK9SUcs+hGraQqs
s0YMCXCbRiXYIDtnJupDSTnUgKIzSx1JgRAW01GbvRx8twG/SAdTzJnKW3hFSV++
x4XmE4GUAv8c7DA1SAi8Yls3ueI0vdSfSzVy5aPM75PNrk2G4PhtQaYoHCM0EYGr
Jlth+g6/EQndFLWqkfUfO7pp5xP2QHQzFxVubod7f4ioQOFzORxV/I9MiyA67PHX
0XTIMGDbpTGufLNnKiXLL3RylqaQNyI0CK53e+QSjVoQd6HnBg4TZjOVpExNfsjt
7XPsfbZHOmUOUryx7BLRBPDQT2fUaGm177kYIGs3P69xT52rf0VkUMvERfhCxEwD
Dirf4Vz5zGbT/UMnzYy8Gvyk22/uWh06fJmUPhjg81wzmLb3Wbj9eelznRbm6YKZ
UIUpTTEDPrs0qyPNkzVy0vmMl7trtUVHefa2m5Ld61s8kgfEu9wfEPmFngkjLMs0
2AcIb91bnelsREQiQbijlfgyTP3QHFxF9htYstdo1IcgqWZN3+OKw19yRuH1s5BT
6avJqvD8VmuIsmzyEPJxjJOVurxTiOE7+DKdO1gUIwHc4LdXozZpmvFC/jJgtyw5
7JEWIZwzl4hqkmVGV6py7rRE+aaWnIgieWE4Gmbot9HdyZyjbw4Ncq/H2JjG1BKU
fuxnjlCs/l0TNB9vZK3TJfewIHGxVylzJCNb7jPxeChz2VNNNMexuyEQABPGwQKf
IHHZDKcSEBZYrkqXCI4ZcI/1F9mQ+p5PusycybPSzOQEfGX7fi/8O77WDVR2di/p
f0n8H+giAiW7/x65F2wizJlMnHIVsFaS0tSUW7zjGKM7FBi+YoWLqTbPCphcENUw
hPbgA9XIo+2P7zbXcxOmsBigALdfmwkwFTJdVyEGWhrqpXm5LDZukFIrXmNFzcwr
oX+A5lQyWCbXZHGnKt6HhEKQ3HFenGrjZXL7YddKiUnWrWlnqRv88Xm8E7S4sLxg
rr2bDIy5hkcnj/oW+6ib0cQ9QroQ/wp6Mtq7tALCTyELRagr54JltOL5sj2H6DgQ
Nvowgiu4ooCOp4I7/YVDBQRRTSx1SiPNCXcAGELL50eyahFIqI4+U2Ih34GZv/5n
jsfeR6KJfe8vysn+C+LOAzOQm6Oek3YlBCaW8emNPi7RJlOXciPKBsD8MYVgicMX
vxdq/FrCgS+PAjugt7/itNwXS8aWJTtEogbEehev0vWnXSrkyaQnINn7YDz3uk/9
LtjQggOKxi7lB0DGA3szU74RZQXGhqhEOVdEv4wOtQOEST/+oqaefM2cz8q9ZPrR
kkW/kxAOogQpKdZfVSJnjjnkCmEFCa4P1pxHF5M1MbrTKvBM6l+B94JXhbd2FFCp
TpzbxZwCPq5Ax3UBuhYPJGTjXthKsuqjIOturEAhztAFO63XQz1Ixc+WafJNL3Nx
SJvSviEJP5AE+r+Yb0LDWR9fpwdmMvD0eIiStufThJ0fgZRXIyMSUeFBScdKAwgJ
QeHP10obYg0hCLz4Aj5cdPaletee51bXzPrPXczMGoSx256RS7Dubg5kGUU3o+FC
XtxbWgg0R5nAhkGP6KD21MDWS7mcPbR53xi5iIFYIXo5gSnyHIQuoJeYT5KxIz3H
hOcR7wbewHNORj7FywZWI5hYtIhvuI6PmPvzbrJBG0AoUKhrc+VHST/yUrJhcn+u
/hKMQQajbG7orQjcxmZis3d31Gg1701yKTUP/lMXlZJcrhsjmPO73qxFJjb+R5So
+Ex78+OroJbFqs42L12yXvIgr5lkZxcpTCWXFykpJAYiifWxXwXuNDvJ4Cy1Uugh
lt0eC4G6gyqpSvMe+g0J3FfrAritHOFPmY+mqcio/lyq/BOaHLz1E3u93aOXalE2
+12iRDSEGjPq3H39DJTXD2pqG5jeRZTZt3qB0zJ2ubUfMZjHrgk7bpw+JNi2/ZLV
3jfLOan8JQodX6QfwYOvUITSu4jc886ifj1RTh71J/RI04zBQz5RotXt7g5FMcIX
knWsDbNhNtkIx9cHMXHF/EIClpSBwl9v6Wqj4QqKorHtMqm6RxNIFQkcD7MklRtH
DYxY1mVk5mNMPIf6nv+ICIBHjR6sq3XI1IuFdQ6mbf9KUCWweneXCGWY0Azq2y3g
FL+5f3oB7oGVQyoRc7MP3Fk82wb75dT3u5pWkPAKbpSNGMEc/aZen97XiahtZ/qi
5CoYZwXogH3tqra3QdwWNvay8hs0ok+jAt8MDMuDRid/VXqb1DMleJegR47VUC1y
8vdI1xVUbNkOaXYz1wgIUL2Ui29UHYRvTuatz/veoEJivh4kUOklYRKlTJ/LogXn
bmITT4tyFCLPFFQouvaZYNTRr+m4gOrhp1xctexb91CljAH/lLDhBL8ncKO+Iz7p
RZbtZhY4tZyUiBcc0TpdmUwDE7Toq4II3PL+jHfBnLhcSj/qc7nStDEIgYinsEuo
n7oWrd0GObUR+b8aeOn7FdHSzsgl0ukMDxaC/FwHBgCwQuhNK+Oi4pAQMouG0ipy
iQ/C9leCZOtiHUxPXjXV+GkI8RksvzwrQQnl0Sjy4rE+F2U0tXH3Os0BuoLhsilj
ZEw7alZqIzg1A8ZXOzgC2HYhE4cjeisRG4uGiOkSjx7LzR+m/H84ijPeCpSLk7eI
11sygzvw1E+mr3mXOhvRcdE/HdkbkzAWriCFQoZCewUMQovS7dPtA97b5wrFhRyi
LtiHhCkWum5kwnxkSwe847ir6c53S2beyD7EDsbpEhEn9sCWgqiZ0llGMVI8nv+C
MdbvpnAJdG+h0hbb0M9Y8NFvj/0U0f47lh2mlz5zs8lCFG/wgrEQ9/wqmTiwa/fG
Dj/AthAgC5jZuBEjI06KaElWbr/oUSyH+SmK/SPGMKLUaH5h/AORJ0ReSwrf876V
ymvpb45NTOih1+ljDheodVGFAXn/w+IVqnkIhac/mSjJBT3IAN0SubybiDmXPl3i
8oSYNLutrqq3bz4UlVOMOoapqhm6/bem5ZFqik972SkgZ0JZpwJfUvBaNRyq+t9/
ASI1pbK1fK3wRmS2g0Pls3RYYCGc/rpU3MLGh1UeE/lsr+EXSyZGOkmqkJE2MeJ4
/m5DTnLepwGb0/APf6Gx7utR79Iu3QQgnD3L2TEUqklk6pllRDIcqH5AfBG4a43h
nfLYhvKsPrMTZE2nXTEpavBFg9VMh9LzwfJLlBmXyZPJ1hyiQHXZ4kheMPKB+yGc
eYpecl3NIW82Du5UMHoIvvTVlAvZMUwIOc4WCSeqKDFPf1KOA2wdAdyPfBJy2O0R
3lubDqSOv8Mmx8Tbeq0b84ngepB8IPxlmJKQyDsf9SfI0qch/8xNCtuhC+yzcT0o
MoI6+Bwuuv0P43zb1amyOi4A+L84iZoPGVCJWjAxVOl4hZii0m70K998z6ZHWTpW
lSJGjoKap3uCu2ZDrVnTgg04xBSavT3zDZKTSKlcwcObMUMduDkSIHkFMFNAqJIb
e/r+88SMbRgXOepf+cBnDFEATd0EMVMwlhl802vYag1SBrWPNtNXnauDspDnfY6X
+997mbltEc2XVza04EYN8R0C9y6ogCYSwHyhYCnVd5Dm0ztsD/FSC7EbA3YfvGRS
qqB1AIQNMst9psMPlkXcSOtTEBFfZ0MPIKkyf5zOb2ELdKCSr9cAVORcbuV8d6p8
C/Uxj6OUuBcjeXhPpWWKiU0pQeGAFCMmeerVHdL/oNO0qkV+FqiL1w16pZP8BMbe
Kh2zKC5r0X48sdocWgml8eANBHMIcQ8DdG3PVl172bmu1N6SgkU6IBYRTltUV4Ee
Q3k/WD1tQl/JGG8ionQWIjIkzDgwOQtcPSgvSMWuG6yI03uhTdh+qj6yDzIomf9W
EXQFRW9tVt2LDcSgnRcb+DRwQrbKoW8sSuejvWn7cJZbDAIvF9UCY4lZc4mUvwo5
kE8XftNqUPMH8G7UcITkYTjLJU5PHNR1DfEchgi5VZ+P2phDB/ZlYUjEkbuLsZe3
rDvPhTjSYbmofpQRASp6JZBVcvd5SrAOeji2IOpwFaF4PV0+jKkkeLkfioeYLLd0
xDSwwOrk6qjx8CkFdMSoTZnjkEIcZMjeN7HswaJWGDFQrUBSkwMuHv2kP0N6+Oy1
r4CI4zZzaGybPV+so70PdtJKWzQduWkT1f8O/KUA7oaYCjLiUONn/k86F9sl00s/
FnHBVapi+O833itDXx/uYcmUT73uJDElkZdCv/EIBN1SROlD7akjs3rd/22xuKqC
1OAli5B8dn9GzA2UTCSCSn2MwoO2PI5SW4spB1ZlJISO8NUVA3EFty75HgTL++yP
ySgNJY6mxFQ4GUcAUpHPQXfYwmBdVE1HRBnoRwFmVPwdei3NnAiIsG5cLlEREcP5
O3ygjFjquSdDOIWAUXYLW6/EkONT8r+jRWln2iZxHPJ30+27aYqv6r+sdUye7I8k
+ZhhCVh/K8V0QsD9Svc7zbDvCiHlE63askgFg++s1FQU30Bj2pVT/vE3vHWH/8MC
1Dq8ZnF2e0NfW6TFzd4KMRp3LuREmf9fkWfenQJ9SeIq860skhLE61iBSb7FZFM6
kuO/QpKODQzxOvr4kLSHha62yEXaGDGskYEKFFaxp98ddGyAO/fYSd1TxYJlcm1T
Qhn0CQQlGsckSRWhKV2uPunEb2tfbwqYLLQ71C8Iaqoq1WYFcAmT7sjqrrX7Lq35
uUHRad74YNh7mapCgDYt+5plnj9N/B0v7lNtT3n9OeTwP3RvyhDaNcXar25KJhYj
QwZdq/Jyy0uuuv6xdWPhUvFwJgBF8zUfQzZ8zhVXGveKbe4UQN5QiX+pvBUevmws
+G8+UE+zlnuZDDSrD2BmfGDeYxN6Hs9OaDuNkew8cd1l+1kBLZYy27dtG09axe0/
HFlIqeAmkglhIQJ9EbSytQgzBTOHyNKxAyp8sb72NIIXRDusSdeqVQ+SvE/29IEM
ouQUzOMrvcTR0K2fp+fCU1eUYgHipELIsV3lb5DtxGbhsDKPpix0SpdYV35jCA7W
uSDRRZ50zPMAagff5dxJc0sYsj92A59LRl01dCHbBHtwJ87o5WA5Gcl27hXSROJa
q07KGIVv16TgRPsBlYv7ZeCfM+vvady3RT7k0WTvm7D7pKaud5izbBPxorWCY6D7
NDSw9lWFppupTWjoLUwaQD1KKOqYu0I4KCKrtTxenbhB7PDNwQZXZGAQ4UM2kiON
sGPa/7Bdovl9Jm0i1pzQdna48NVuwxq2cZ+GkMJQt9jMHIlNechOTcV2CHxtOe+0
Gm2HRPQmmXRDK/RYfGHKnw4pSpmStjEx/JhJQikfG9EAQX5IuJhdqoHUbYJLTjjs
3KlsIEuGjoytbXuLfzrICCWFRG5o6mFnvBrIfq3RezmX/EX1Zt4ErLQZJGI70BU5
6Bo3wlGwlyOzf3VIjZfImVj0Igu5LNzu22gTjR7/q5KVv9FIy9tKfAH03clwZhew
ynk2nkveqRr+ylkirHWnMT9Jx1dYBSDAjCL9WNiQW9DFoQuY/VC3wxQCuT55q95r
zPT+e9JNPrexeU5tTDAepF7SFFxhYOEFp5Ff9+qm634nSjP+FN2Z4Tt/TJiQkxBV
OUU1c7xfAyamB3FONlpRS3iaewbRoB2ZKAGyFvdlbszxyPo/dUOwJ9PMWEv6eugq
K7TVmj9Og9wtcLUUTI4A6+ssamXhapxGbPgA6chQBfvbce+ewoZME19bJ0lt+OYv
EYul7BzRrLYJdWzfVD5/OVQ4vMI+7wVU+UBYlZh9O9J7tg0LojkEl4JX7yOJMhZU
7zpUyzZP/yKPcI3V4Pbz9oSrGPzVs2TsjqzthGmZlsqvi1LsMlW2+uZqxitIV/Pt
AIFZDb2Z/uRX2nDaGFKQsg72Bf5iKAJLLoYRRMAwzwLrtmB89RFUuUS61HYYMsSM
f5UY07KMlUXhKOAdTzzXDlTo09QPTt4VJBHVTuINnFHLTB2h5hKFkUKtuCQmB8qX
cyIaNb80+cyUaXpvOTNpY2HswqYWYfdjrktfg1XOExBXAQzoCDv/Rz0tf5u2nQZr
OiJmfuafurjtPq0G7ArEg+z/6XARFv16VXnkkzBGfdmE+ns5GRPxohw0inbPlrnS
kRgKQZ/WwaStiOZkdrZ3/5ZpvahU7CRO8Q1bq6fubaxNktQHtk7Y+KBCFQ97Kf2l
bkaP32Xd2SEYpml0SGqaUo5D7BVAnVMg7qVHCM1tEalkaGRudu5/ObuBCiNxmv6w
5s7ZTygiEusd7zC9lPWL96wD2e+rY52Gc+G3F92vux5ySzry2fpo9RTHQunO+Vtr
QhxZ8x0rRb6KEqFse/ZTuMoKhPKcQLlaMczfvKsaO+d4v3k415dAFLleWJyIcJLY
Yx/9Y5GRxHyPZKx4nAQHKoKi10HcK9dASsKiIvz4McfUWdWHjfinGjYPaAGouEHh
aQTfEKnV11poU6L9cYzFE6b3RvpryqpSqlJoZWd4UJsvy8oe3lYAG7+yXdE2JI5u
Dud2FBnhN9w41SE/NFjotf6UyNGnnGNx/Z1IH6xYEPU2KQl3yEeYKanPqxwgheiI
0ZUFKrMdNRuAsOj+de85BslZWZbOj84B21FDYjVxelxEslTH7wlWxlGMDeQjTqG4
OqNZ0E2mPsxACxXNot2UERQ6ZJ+dm/9/reDq9UuwZx97saTp1s6lG5/p9QUyZClZ
2/fmd3+ahU/8ncWkXyZDVgzwk39X82AbjQKPzRaNobec/XasCBNPPgn881DI5OGB
P6EtK/wwe7bgAPjSdPIdByqWthZNNQet25rWI9YWlZEOxfexzEcQsQ4mJYvMdN0C
2w8yVK8TjnU2qXgCX0wtRy+rxdu2EGLQVYNe8fwDnJwB5pcfO8XjfqOwR/MRJizY
pMU1EmtI/2tZD35VHx63tSjzpWeYRnC5LY1cNXGydJZQr02D4ZxiqNy/Fgsnht3a
whipX2BxJkKroDAJ9T/I5AdM9nyvf8wzgSPEP85si1rEteZk5EyMQNYYtPFWXynU
fVgRB5Txm0Uf0nmzBuuKLQuGiMopjK9TSL6hq16oz+l7w1+qdFoCx874KiVn3U51
NqY+MMbnVF4e9/gFihSzVVQ+rkPHZvN5Wz2riZujn8f692dW8tS5uE01m/+8H7Y0
H6yuhwMwvKLnG22Fv9MDZEhBrHNHIgnrqx4W5luQA/nthFpjo96o0GpcNXVWxVr0
qC976L2c2ZO+AgsSNg+fEpWBzJ/fgSgi94uBEmEHQDqSvDfeyig6KGd0vKZkCj5C
ybkmL61qr6K8Vcdtz7HXTmMJZcYZMxy7Cc+KAqyAQ3uj0G05JtnA2XJSUE1E8PxS
rG7MM3PZZ8OQ/tJb+EJm/xv4Hip01t0Amk5um/1nRsWcCVmbZ4RE9nDmLj0AHJ4P
lxIZ12FqCS4cskodUqXUB84o3PBF6Yu7ybfohlvZjBm1X+uNlg/lIMzqqL7oSbkm
9NcZxuQVFjSjxHR1WEgjjed9hP8pRVKLUoAN1go7aelKqY0J7lLLY4y+0oz40LRA
ln+YiSZTF/FIXG7MO9QFQYCttSspzZPeycAfuInOfgWsyrglIlxM84ZatyaawKfH
CowhUPl9bt4P8c6L0p1T8tLv1Ah0HfXM2TVf87w5jfLyxcan5ZYLaI6fF4fgYaGe
fq7EfWEyiCkyNTuxkVqpAFTS3hG5Hpgl+wJxD7TPAgvt5+lL8AVcjNEFUy1GmNNa
HZUEAAID/LlbA8l7mgRtauHh4kn5pu9s9tchC7g9ZmAeOkphH29nWemDg+6hgWn+
5Kw0Q3ulWaMWlZj5rojTtllaX08pmjak2+RHy2uiqHaZP2yIEC8wLqkTOWBmfOC0
pvQBJxqm9x4VaJsPN/jAE7mT+vnG0df8MGNcNuE5ndR9U8+a7eBiPzE9MJYyFIP3
Q3ir4vv/GiYA6WySI9i/mbU4W85ztzY/2a03UawEejy2BfdlnpU42xLxzXYPwQLR
Huvvue0aqKR/HlORlGPogKtQ5FlTgts6j7B1fvVKpfsWbw2c5vy9jtDkAffAnWBg
u3IPXtl4Fw8ZlccyasSjRW/e5M7pwNzrDDvw+3Ni//j28fZuFqLv3DJy1HakYN5G
AfFrifefpUzkJy/kuhbGe3KdbFxUl/uRP6JrSIk8+o3NoCagiMez6QPwoiFGDzDd
3S7XL5oGudf6GJwtBb/N3BMMPyG23oKnaCCE3WGlXF853atJzGcjSdtg/JlZBDC5
rc773EVaWsXPhJpNOiq+OMLcjtcaLGrK6Wow9wGje/BxBtl5BR06pUdHiwKv19N1
KtMZ/XW1l//3A6R0zMAWka+NL9jbFd8QZtd6l8oMcKjaeZRpF4PWYwvstkokTN5q
QzxYkNk3GKtKNNygTgJT6lVNb3xfxyb1UwfIZmlhCELxHJ9ymP9UJ5e7+5fNC5C4
JjTgx+GpnSM110c6j+L7b2tp9Ipi8Ho9LF+w1xFr3aByNm8GZWkZdODUhqcpI7lm
lBJwreHzh18iKxTrJO+Li4mQ/jQIYrBbOZqj/w8DfE+LXqZ0+bgY83p6uJYxe5Pp
46JcwlRs4jBeBTaK8X4Mp3WY/kFJ8GrrwUxc/ADBaGdlKeVea2LVN4ZMPW2geVAX
5YDy86h9qw1MvwmsGN4AsIl5wze8vJqeLTyLOkU5Cbkq/KivHPjxLGLy/m1oVmcf
l5ZRjYdP3u0zNb/n/CWMU68KQhtbMbrIIRWLMKIIHf0zoTXS/CMN8jg7QC+qcN8m
7teN6xhM1XBeJrysPNyRMj5mzzwDLKe2uW3EncvGOe4oLiP07JvKToOO6xaJdNfy
zWJG0hMQr55CDVHlmdilCFaFgE6b89ev0YiSvD361nC/dexQEMg1ZVjmxBze1QR5
TiY8tyu7nQjAcV2ctRwvOnCS+Q8cZNIKCGsic9cZ8Y70QFBrgvZFqk0oDoKdWmR8
3Dhb/Bpnw7YKC3xQDZka/nNEOBqzpFsD4HMN+lJFIiwt70h0vNfA4hWRGBBP2z75
pQKlFGARQQ2F2/Q/qmMgtgTiNYtrpDthbWJe3Ov+nNmXHI/EV3VgnuwsLA7OtunU
1L0STxapAX7iFK+1Yq1I/5wEaBFyzL2cP1I+/Y/uvC6AzqXca28Dqz8rzdukw66q
0SdAxkN0tSD7SUHKq2BnJ8iYJOZ5/Us+wndNhsa31BBwCDvZqB4BrGxtrWwkglMS
fDCclSXAL50YsVDEVEWNFQuPqnk1DhEQNC/AJvmmm9jW52d7ssuAV9sPCH7lQLAo
I23b4k81eLVXslXwKsVaWzd2HLoCDcM/WrGZtw2Pc8oftuugGQNXkMh3EDwSNVjh
uHazi7htyOirEuGb3vfUx3ELBoHIqaojhBO8UV1N2uCnlD8ddz/LuY76ErnphLSW
6IrV1yg4SFVsWNwGg3415K94YdFSpq7GkSaQ6Hziri9BAGK7hvxPZe2Fq83JA5aT
PuTbHwpaLiRNYVx2QQPmKHGQkpNxJWoCdJliLCWFZNcQSH+SL+OKSy6Y3H4ISlpL
hI8EGE5OqtoSi4xZzn0jcr9wYS7FWsz46IgKRDKKN2Idn1cUruUNLyrBLxbkPzTX
G9bLlb1tWnf/gWsSCn9lwPZTM4Yw5B2ZPBMA2jkEiNh1jW0dDJsbJ6U5cisIjW5r
PFh0p4KMzMoLMjVqdjFBhCUT2PZjKvTiA0mvc5Vz07DRA9o0JClN+5Zyr6e63nPf
b4zUA4RTRF6wBXxDTz9mdVzE4LYDcrvTFKqYBFfm+j6rox7OLZA21BrOct1dcMFb
Tggn8VOZmxpQYTNiVCUiUrOJM8dKP//fEdEQ3BdaTyIRuNK8rbh5X38b66u39niM
XVPHKrJD07idPr7CF9FMHQVAOkAg4cva07ah9LNuSV5nY+iAwt/j4cGXKY8jNb5x
zu9/Lz49E3b+O/rxR0YTHd+ZkBHNim7fAIL5k0nMrrFgYAaNeozQBPQNbPSsZ1QH
JU4fcYKNnnYyer07LN6TgEMsu2fDgpQnVHSF3QSSJ1PMWbonye8HQdM0p3pgpSET
jBUa+MKzmJcvL9DuhSrc+YBLg7pzDNu639NN7Kg6bqi8KcnnD1Z//CDoaO19DweZ
LO7LQvPs1AUaXzknb4ICRmdGkEIWvzOO89wqIMwkq0f8SQz14vgqdox6DTBVj6sG
GjZYAf7lLVMOgP8bhE3a8n4Q48VnjTXB5iUrD/59S1MKipfY6EHUgR9Q7YiMvT1x
RCqTggEvOsTvZimnzG3wQXLqBFHqwUnH3N27gXO/je0WuE3wexXnm80BZNDda18w
4Ow9ioYyxBeazB1Lhx/IvTKQi97+NiCQb9F3NIVMBnHULOvnRpHRqFHeIPlRecFR
ri9qyNaa18JMCPkuer26vTGoC/Ix1AwLFwpC76dc33m6/wOgws7iPccmlxnyOGlR
mmoS27R1cukj5eolZHb5sHrBCpAyfWFR2MUDN2pnIMgTCr5HXvqv/XNFg7Gr0/OI
kIWlep+3uW7fzGaKMvL5vqgN5+02CdJtIU9egygp89VaaSGI2gZQZbisrOIhnF/L
YpsdLFDtfI7ugZ7qnB23NrOaetLaH/JIU37DMHHGCNkNtvWJHBaj7sqnvb0WjopI
zLc31LP25VG7+l5CmIxw8FoexaQOsgI+VAV+Z1YOjBd8HU4C/3+M2ytt/7YnGV1B
a+IrpZ4Ig01BAlBuG/ofEDJt8vXNPfouYk9Xp+OQ8tSYVldnGWehs3HdWY18u3jR
ozhEd/TFvdPyIW9Q49yFtz7Axu9pWinz7SMeJDUwSogNPpASLyGMbvbBxgy/dR4f
2QVfT77UgM/X/M+TCqaLixa6XXL3cAULTWHgqnMiBZ6Q0LoSYYd+jvrDs1oBYYI8
7g65P0Y/DU6pPnzHmIOa//CLenY2OZmH3ItA1YgYecahRk6bIAcBh5V/ldyvyqTH
YacCASN5G5ptgFXConOf2pfDhkaUmsJoKww7vpruFReJQegTk5YJUNb/28r5yB8V
Z2WBGVS2H1QxwxJ+cr9wXWxfwp+7kMm73qN8tOUBMwoguQ/kgJoz7xKV4SJWpmf3
R7xYmvrrYJxCBnpC/cGjf+LrYZznKSgguJyF7p5VgI+4S1yfwy9ZxakPTUm9954q
HSjR7/p6dAe/5zXso5nRREQ0dXcyOKrKykh9Z7jYSWA5Q3XJXC5olh6xByLWhonV
3GalS2HnmhCOko79m/THc0K0rhJXexlWNu6oK9lkKjY4xKeoZY3NfVPruQUFohV0
Go22M+QJEw504ZdAutewiSPOVcg3aN/eLSqxW/kJP31lIGUxB4W5VZNr/7ykJwFI
23n/cgJ3JLIC1KcAqKafOMI8W+RQL+4V/WiF7uRfPi5junejnhoCvwVYLnc+/zKX
yIqPKTTrKHjErbnFJZzxzpmW2FQEaij6+vstjWYMpsKsa7Whhc8fM5X4cn0kqAhM
/37FlVHqOzZ5h68THxd+S0QH6cdbezw3C5ZeUwSH1BqlZqSoFz7G2lXMlPmiWPY2
rAdDeGeXDzgqeRyCnEhC21CynxcNkJMg+Kv3DREO1xRcSSheiUOifgsIuJIbFN1W
XJkKMBn7emHNyCtiwJu+292JOgwQpEcnOUUnOC8Fnly/5WOY4aMB3y0ZS22WqxY6
yfl5N8RmGjkM27CJtdlWobrzx3BADTcEcA37aaMyAtdKiKrZo8mrNqI3kuQA3Qw/
Tpsp8QMjuvsEQqDD+4HZi9TA1TLE0vrgSJBmla73BSoq8wZFs7C8xppgALNbxgtM
XFv/XkaOb0HD/fHoz/uJpJ0nv8zQ+aBzU7uj9s5v5oEIQHhEJZSo9Eh+SgmorHMR
eXomGRfQfY5wGW3hBXf+S5/vBGGit40OR7JEANMBDQwJMSZJYiuktTWajhJ6X+39
Bvc1SqszpaAVgxZIuNEJ82gJ53vZINfLeEVpUnMk7WHWab5r8do4ryUE1Fydag6t
P1lPYWuISu0DtzxlNzQuOeESACu62YQdv+AIk3EA+U+EPbPCWFMsUNNysAXa9wSG
HcrJgfC8CcjTA2lVa1R5KG1Ut+m3ehfe3OhO3aWyZbHIiQOLhNCg1NnlW/vFW/aq
rl/jwUxRJ6UrTxCZlwLT8PjSwGw0wViKlSJaOGNZvDChPvYwsPOYMN/NnhUwFIbL
chIZEmYqEjoYm64g/c/VVvCT2m6Ql+XiOdvaPy3YqluL1IN+llsQuJV8UDLOESEh
twmQ2cBp0pGWGKZ4K4KeNrc4zWEntlaJVXuJgr54ufmbgh5uoulEXV1Nk/q+mFhs
6JFsYx6rFN6x7HVZkNgPf9eSWYyKacyPTMZAGXvklYBXxi4d3aGOvCO/TxXQHUAZ
2dnURhC+6iet6C+Cl92J113oMHWZLShjC99yuGHqqjm2uX3YBbX0tEelHy9C70S+
Zjj9Z1Vj5M8l3zm4nPZShE7X1S96cj7UfxlAnbxfKYWk3WSnBRh/YU61EUd/bLMD
8t+hLUQ2xYXtMRyWqN3Lye4vzo7FwabTNkQKsgx7qbaQW53PwZ1neYKBBc9W7sGp
6uK5u457xOlB+7H7JMJ6Mt80RhEntxNslbMbGrMACEiB6x2FinkSlGi+ZrsYyA1W
cVd3P10kb+c0jb9KZ4cix0HL+bm4J470QksGgReAwkyZtnznBuwTD5c5FqNU9NFu
Rb5ZztyqPnJC5NXqG/yZev6LrFyl1DvU/pWR/rGElE33kf6mffrFdPyc1cN0OBi1
K/C8qKXsCyuRg0FVk3wRy2gZsR69WFaFknkTU7heXlEICISCnu9BkJwucBRp7Kek
x4V/hIhgNmwhdIFmcgUjyQjEh8vgUAlRodLeL47STfvVRQlverzsF/N8UEX/lfYJ
ugZVMYDBEavBGk7KQ1DW3Ppo/wtSxS527wW9nA4cSIByQ4w2z/h7+t6YUGYfO+xF
8ZtKiT7bdqUNTeBJlxkNLR5f9njgaBu8aq7IngZRBLwMh3hCKq2uIrMDQYizi8xU
jd1fnoWWwIZLSDUiNEAfnRzzT8s5rV3jfe9VHXatucqza14qQvLPldoWt1l7NYF4
xSo7fhvmTok2ar7yMdIb0vFO/eCSDRUhagLW7AAUswpxrS/XFt17Xzqcl+izvUwh
kHPa4GB42YPoJ5q6D3yPy3GtMX+e2qKh2ztx2GwwuSE3rh9lEjy2wc1OXy+T6A2P
RdB+YoMgLZ6gCgKsxW0ss9uXPJ85E2NlBvdvkHnyg6R9k11hcbXb3rxlUagSKZI/
R17enNCMBSIH5fFbHA6r7Ffs71O7exnd/IchWILo04DSvhQiX9OY3syNVdumTn59
5a2zHgTYzlGGVSLYIwLKLZLQakJkDVVmArFiU/B80+yBWeEzgeXxtSfsGU2sIdUV
9G+JsIqQFWjkCGztAROsbRoqQHucLUE3WCQZkbn2rRXnZsYncc/afEhu6ENg9MXy
Dol8pCVsqbEYEN83zgKB9fN6wr5m2iv53fCpX06cgW7raFae3Q5nPOm7g06stYmT
PmO4r+XJKkOhi+cVzwRgh8OPr0GgCKnXeKLrBftTY1bVi4VY+MFwdCW/Mma5MrLz
MUG3KtDs1EzUFxQvu67wCW5PGWuYbPpu0Jln/38EESQoDN1qBpUCt+XzotRqASVg
Pn8rohKlzcx3or7dzXs8g6TEXOe10++RXmxhlccTKHMAv+Krknw8fYNrWEJqyOTG
N9XLFClByCA5kP/RG2cFZQvjJSXqGZSeVwDbZun1lJI/BiIFCqw5bnnxDbEkMQVo
ZFOK8FZAhKT+LUUAHeSZWWY4hal956vlUWPwqHMGQ4acWuyxGebEVDIrAIzlmWz/
TaFdZ9uUXXJs9hY/x9W7gRx1x3zNYDjY/F/xq5i36SlqJAT+u2ocbIuqwIvr92bE
SNCjZBLTDI2/Dff1pNuZROEMVxg0MsGwwQU/xck4am2O5hp49rzzb4xPTNP9hEK9
/SCOk8TAgSGOZhD8KA9dL51wPVF70+9S0MuOJOPXPN020QCHf3/S+oJWuHDxqbl0
jOfrLJaCyMBfDfa+qSsXftLjprPjpOaQy3or/otUTdaHvcIgIIXgZl1uDnsc6vqG
kCxJszG5m/rxfuNtrUrr7UwUcysWKfwU+GI9ISb9WgqZI/Hqg0tVeeO4ET9o8JV1
Mdn3bZs8JcFiOSNApG3tl7JMBnVk39k4SdL8SYBUhYzFtEsXuNrmFIYcpjZt1RQZ
SdQW6fsiMGkgHVbdk2zfghStsSoHVKlsBok5co8waZbJDdc8l1RG1C8U9fM48E7i
/EYzHcF0E5ttrpjcXWmnp7aBo24YWtAupNp3U1AXp2IG4uR9g8dpjyFIbWMY6OAR
q6MUMwjEUAj9cJIRK9dZqfSe/buSAA03OrfWswSVmCDGB99T729yYI9obZC2d024
BSRC353Gvg8Xmj2N/iePnNXQX1zwPXcpy8ZOVft37KJ7m7l0fHE2JtlNoO95jyZj
He/E9Vvc/nNOsw5Ap69NrhLSqO7d/2gxtSpyZHgIxsvO5zMtwQ5elHxIYYKMumBd
+9wqr93PCbSHxwiHpqwJ2Fcbecau/LFAW0HRO3+hK//SEbnHlR5BxHFf+7OVb654
pcGFbnX4zoqZ6cRyl1Dbl5mNsnLnPY0z4VbbMgnwlpplm/ozwhjKuk2vVkSsuQb7
Frc+guNg0IDaLPF1y8uLX4rWD5L5vKktVwmOMBSr22G0NAJ47q7UH7weYwU7beQl
YAjKFGDys24QultjnCeKPwrT0n9ZlysP236T/6ccfx7D/uoKIOo/XUg3skT4UftW
vIHYbP9J4zowzKKf8EUbmSG+jfof3bfiAzua9TEuPWvv/DQleRCGt7V1YZOAWhED
UPKaMwUG0whhSMkyN7YaIrkkFuyYZlhrRKyc76O1hv78yeQr55re1d633JBnHCkP
dioPAGtCDYybtwc+lr21/IXRLdC2JbrCe3bRmFABRrz+LADZhrOEki4K5QJeNBAk
4JwrTbv1JdaWFy3NxXlbH+RQNSe0fXDO1EPYpVBp53bG5OnFP9hWgoW77zuyY1C0
hsnGvW3uJQ1PQ3bGUzAU0KdE9g2TwwFQAenNxr5CS74ml/fEDsNJGRg/awHUohHU
MRkKUgZl/UOtqwqk72AHngCcARy186hm/9vpi0zCjvi/YBm65ZylfGMzC5umaWhN
W2ArGtoAw1Jbbz4bDY2krPNBJX/YSoWJDvX5II4o1ClpBVKZ3lJkF8leopXVnUNG
dFWnZs1qUfqvr+01fEdFPFrHz9m14uY4E2u0fSAfTTfVC5pkYfCYnsOL9WnSMYol
BH68tiGENEZz42bTwYSq+MqBhoedKlwBeGzxyycJuzUozxmppNzakXZ0jN5Jfg4k
NvU9sBNXDYrEJXpZ4hDW1Ljmc8BFwN/nVBzsV1mY8vwBwByrrIzNPigkqnq3SptW
vp16HLGMfjy5TlOQAdWAvGPFaQ2IIOtmYsYHpw68ubDlg4D9y9BuvYNRnDmGCzai
nUZIqi3ag6JBE6gnaNvo8gXCXrlkmdW7hQJ/m4fF+kYyA4RPHEU+dCcBYQw+n9jG
dJNKS6BWv1uOc6YZAV0o8M6XV891C9RtTV2AtB6nrD21ryvQSybTE4UmL9gGZVdH
yvyUn/zoEgBYwpH8Wz2HsMxG++uZDwlEx5VdTlOhhWdu/ZmXO1xrDFUbhNvMCObo
GTIEOSiSmDDaEFbt1eHRJ4ZFVFvahkmZwMfkhX9xRiGTTKSK6VlK5jhjC1V/lit8
gwkh3yHKfxLAbi1gIAYXzsc7Px81u21R+BI8A9h9SM4jW6/Hq3cPkNTri/cZ21wv
w8tZpm6RPlcHjn/eMXUT4gCXkKImzwoSlpw3PRLe0r7E7pD/F6EqP6YPHCrfkf26
nG4xATDZ1zlYKMvjy9ccVWu3fVYltIn/cmM7aM5li0h8MDM4hHHie9oJ8FC7C5Br
7LbIrEeI3ivV1iDMZSACR1X7CJH3RS2JB5MnwfO4Kzej7GYaMxiDH8PtYZ//lah6
AImRW8JJKyLElcZIFFaCIugx2ZxFZG/BaCRDNpuBomcins2q9IW/03inu/zlCME/
0ULay4cYIf43sV3cNpDAdpYda0wZSsJLUmTW1nH1lUwQABfEPYwl4zvXXqctTYnL
5G0lQVqpumxpFoTzn0beQj/IhF97ZVHtXKh6ATHVUJQQjZyCB4ItM+WN/klA2J7k
jt9/jPWL7KtFelasBf00/JPaNBEtfXYwGXEx0gaYTigYM5OTuxBkcP0RXkvMJv84
fBqUYnW2z3gWET1K3kkfVgRCQzvD2aLa+AXgQKuWg93PsOrMTdXnTExGn4A7yFWA
UrvkFc3DlolIlEggv+5NuP0O+wEoKF6NbPf9OrFFXVB21mNEa6HsYNLSmGnyhkB1
LXAk1m2SqcSuyareT3OPIGRubqX8X5d2YomyL8lI5xObdLPo2/QkVfNxAcq94Sj/
J0bM1kxdtt/DqKVxCn1YXaK+YsG8AxG2CjTvqGkI8HfEviYGdD+XJgPi7oOqLQCq
jghu4Y2Kfpe2dQLgDURctGoTygrMZ2slFzo7CdZpa3IeixzR8xVZuE/THqlnZxkZ
v4iLhBx/zHKh+lUfxQcYzOCg2SsSmKW6S8k1taUP/mZwGLJTDsPvNjq26LmVpi8H
nt2+HY7Li7nte7aAX5WunD8TtY3EtQ/9chAoHJLUq+1pH3Ds6ybxDSOrCCrc6pfb
E88V6egO5+XFeR7SPOvrvexNwlwbTA40qkOM/5LlHa/zBtkBvuslF+t8zjW/sryt
ruGlzuKirdXmH8rpKYPxEaROyxJemi4/+Y+m/CBjG57jZqeD4jRGfg9maWp/+zjF
W7lqNz6YCb8wSiGnOotejOB7emTWuT0JvRRlZSuqrnU7pZPq+z2J2VwP4rtKQLTw
PgWs9Bi8qMMqay8eT32vbQ5u24FYsUT4KyhuDsFVAE4/dgefUVdMunXiSWfmvMPq
6AXi8U5no9R0dbASXjgM8OtM53uiTkqhkkoSPkRgAvN44pzEG/w+lOgrv4C2P01T
pyrZUMpGwKcjjdN8311WeMhNyY5RAHJZ2aqYt99tblwKLDhbp5Tj7sdX8jFg+qbq
zAnw96lIKeegmpA1c1wN5buK4FHPwOH2iR7xlEyL4v8xouG+l1YQL3v/wBVuGMco
mP6tiitD7tV2R7l5RAjtZNEj/RwaNFDejPPaiUlfg3fgGi/VQ99SYut3K4UI9iGf
7AjNCXoVGl2asGQuBsAWyfdKS5Tmb14ezRuP65BIKhj6Us/qXqNV82LwvsAvCkpf
seCxR2EE/CMExL4u2V2Fphq8lMhjBejZMkACPRI0u1FE47d4jG0lsVJXd+hTbDJz
4OJj733sXqHT2xO1OaiRmkIEs3ip6Sd3t2OuOBnC1uGfYqdOIzU5WY3cu5+lfadm
NxMceI+DQWNpGkah+uaYdrLQiKpGuCjMNcaKo2QBPzqIY9llbMwEPo+M1eIgeF6v
a+EWetB50eNTYuNUyARyVykcuh2m9MmA38WiDjsCaJf7se/a+Cy2I4byxfBw+r9G
WJpSguMVcKrgy6fA56zOEL8UznnYIKhBoz41HVPYYBghx/mynNuFlLJdeIN6OTea
+/i6dc44eysx0rFCEU8cGNsiiUpIUYasWsqyKkOgJ3s4dO6IyUR3jMuIK03VohxC
FHcO9RGdc9ZRFVTMQ5AFW4jitKPYSTRqbGNHvVB8n/DCRxWH1Mg2cl5Ygb/44c62
AT3hfBEEL27daiG67zM04wuM00JnTipGaxs57qJFkADPzJQcC6urdq6tkhShkfz0
0HZymeWorkJiKVt6gM+9MSJmKD9VmGR0jsVgV9w3v0AG1KYu5bVDv+73o/X5Eaps
n4ifNS066Bs3Be3dmHT6DOIUUno/bZbTV1yp+E8uJ56e/3ZNFfE6JbTiZZTyH8C3
+Ou5QUj9/gfUJdvI12Yl2Xef1kk07PF58y/ooK/XNzpCE9TUlzSv1J1PCf98etIp
H51JZSHpSAiKz4GyUoi1o/W5ia+cA4XRXmHxTYMTymMSxKd1apIaytyuP1OldKj9
5l9ohk6iFSZyrmlqiYldx2S31fJWNCATLscMxBXaalQoCbaHtQN97D7xIWhaszDj
VxtGhR1+taaZqv5D0vSbvh0FUvzgJghfrYId/4dvEyJSADcnbJNNRw3QbwKqKopt
VhV69K77omdM3W8xagtMOTyupCeWODGQnttuz8NXxHb/7k1Hkw/J8F7LCMHRxe8g
XoUOQzAo5BJteL3tBLbwbYqLCSmklVP3sVfSJkvrTBznEaRpyZY+pEpQZ1oK/dkX
8eFMvPddOjTktscB5jfQZHEI507WZVQeQqpQelBE1l14uGk3paiar7KRzv2bB7h+
zH6QyLKFXxakBB9RvWb57qjqBwXGGTROjrFoaqFdPR74x5oLeIgMWSv/2ZUebxfH
UJB9tF9blSA3QTrTScD0aIkPzOKfP0gGgXT4ADPIRwwAy9P9D/HXuDf+1/1Oxhgj
7r/9BrCjx7IXWwPeYPvYpkHKxyVibgtp6ijCZis3tnu/yB3MDq7koOxyzv99/BC4
WDpjZNXxh5gxZEliFRIBEs4O5R2UlB1shWKsuteHBtOR8kpbw+KR14fH/s/6HeaQ
jlk2OY0PvKLRbszRs3dr0w3yCPOTsQM/Z5wHyfjLX7oMHd3SC1WUIbeDFZFlI58Q
tK+Ac+K8NWMIJzyJh3SMilNY7xHB2GqHtMClDLKjCeBvCoZPMLiBUu+Hgwv7IU+t
xhiOG9FDL2PiQ1tDM0vcbiNm1dJMAc/kkaXtUOt8GJsZP4mkMysd8sAeMz/m3xxH
/0VClOrqcEA+yGzmCLnm3RRFQILNbVmj5euaaqo104Fx75ls5rwQi72pVakgesEy
4GDjRNdY4Ni3Akr5ofqFWBmEWSeW3npsf+oz0rjSQt7mMlq/zgfYBywwRhv5PZFf
Y3du3Rq7dsg31F/xP8cLry89/ZRveUXLOoQZDOIu2H6VgfvDrUICvYVWx6hunqoH
eRXY1Jm9jQTC43gjYxqmv7RgM4tuu/6e1TzpDL696Xvy82xOJJLHmHUyKCEWVfce
n8kVmFzSZek6Tnj6QKT4dzhC5DbBxNx3P0JB7h1vwEbs11Ow33Yxpw5Rv/EHst/u
Zp2Uy1yH27OSeoq4K4nm+xVVKwkPsJHXuLzy6TbrHxMbEaMRUk71WE2Q/hr2lOgX
lJhFiRBhf2yghpFgrmRBchsV564WcTIkQgllbGgvcNP3RcLhBqViGgcxlEySsyQG
NsEBXvO9GLgRvFLoDf3njgvDZqcxlDDRasmwJayGezh4FCmTkNIAzsxw3gpWVGtk
4cyEhsVLCqoo5pt7wPFOAeriGByuyIywv7EWFqLxTyg98Kz93ntA57J/I6QY4+J3
ifSpIBqUdqJUwg5EkmbM73t4RsAJ4lwV7WyQNQyFlk93cUs8xd9CeLLFn8XPv2iw
Jw0VwFRPybVd7BPW0Ra6bxVd2aCcU+BKQg1dzo7CXiOj81ydAphQpfPjaspEFtM8
85aQgClMFXtc6BIAlpjsxGas+w/0UnEycVG2q80C9h40baJGdG7JQMKrjeBlCNxK
PZA6RXMW9Qk7wIUofWmYU8UDKdNa5SHom6Iswu+HCA2KNXXqly11nGNtSiJ8++LN
umlp/hVv//et+xiW+fHz9jn1GWcbjJ4aKJRJ/7QGcVZEIL000Z5XiDJohnw5O9Es
AYRzdt8vC6Ov25yXGRVho/xmPrFMunDf+ZAzi8A5j85vqWwiZTnCkBWq2KRWAx2+
wBuH5KJVMp7J/s8ePBla1Lv3MMr3R9bmWMYeOP369ukwbiWm96kEma6o/wybPHiV
DqVRiPOgQYoi6Rj3gTGTt9PVkXvcmd4LiZvufFFbpB9wNq3/ixaX30+t84cgKR2n
CHKwO1zoT5+eUS+QlI6HQAa4ADbvGHPWJkKewMIJeG23fmDSYE8YaGL8YG7t79so
SoQQoLV3NT1LvLAfc+SDHPH0ctbaYE14cr91Aia6EV4xc9iUTk9YUa0A/2wcDuaX
McKroWGBetTmOHFA/fAs50HORFriPIFW/Jnsq+YnLMAk1F2ti90Y78y7VkIjOemb
Kmalj9La0WgUM2QMNSQA/NKQEXqKJVhaWcte6wXB/+hLiFVG44QAVEOEszLMgyQ0
mFyZ251si17XxpUA/uvZ8jUCChPYvpxY2UCu0NeziE6hr8pX97EFplSFwADWR0v1
eypID0/LvtA1/nlqE7LDkFEQcTIOT27aQpq39i6I4CzInZSskm/rMEKLYCkD+p8k
6S6zHHNoiAty9Rqm4745GdVzRdTb5Z4qRGmaztg1QysZgt6JdIu0qxGO7qW3nx25
gU4nbl/+rIuP0jAq+rPDd9PfkXGAvUWMhMCYVNlLab/5Pa+RXVhWzJ8or/7I8Vf3
GSi0fzVRIeICq879NlZG0kmLUZoXVa83muDOPICbois+pn0XYTN/Wad2hqV9UweH
ZNMIKS9Pm5W9du4N+u+MfmpEgpC6KQDBlkz+DwAylxN31sGv3AuB5f7EDBtgDR8P
sHMObVDTQuLutS60KEgfb+Qd308EixLkRl4whfQIV/yH2sp9kDCvQRiaFjJdg6F2
fF/Q3x35/ttn37RI0dQEDqkVrU8intM3Qp8B3J84Vm04+MPIdtwR+dqHi2HNe9Uo
Yi9H03+M1itBQYaeAYoaqAUVyZFP5WUAPMqLIE+UTiiwDZM6q7xjZABbfUmITQiv
QGLjtobY0bq25D8FdtpPIMuLRcVE25yNMyd3hNbCt74MT9iG3IONf44N+tWfFwvt
bvcX2rjatn0OjGTmAsV68KXn23qYLPZKkSmtUaafNYtiMgXBqp/sKMwDr+HT9o/Y
HGwozRchE4EEGv+Xq1OFUa8O/tVClk2gF/yWXlRoVPViDBaHTSy9j98DdMleXFSM
jYp10nKdydrotgajFDANW4tRxfKR8eAnEWXxirNtPPvq4kcs4AyKB3aOniPAEziu
2PiP4g+tsY4Jkj+EoOJt8ur0Tv8bcpPOnQ5VDNkGsAnxFGphV1qKVtbrlMzbMKMn
QX1gnaQQMjluGqclbMFIDLeyXXJ8qAFuZu91za2cmgawr+fqPlZ5fOb6iUGCNYLR
RMB9cBkCrhkttkP0c5rEXIhej7bayJmkuEczbI3+sse0tegF8wERjKFtxPPlHg4k
fBEAZ1tUVA8b0ElDAApNaXCARwZshX1GeeRF5RbhZkTJfezW75lFdwLOmsd24UUe
yAyzgmL2ldC+gSYufPiamoINz80evjRK16i5FdLGNIPXRQHLf8sov/Dv12FpzvVG
qfjNbdScgCLtw21rC1Dx1qIiochD3Los5NfRuve+iwc1Y8F91NcHI3RqcFNEuwX7
z5wXp50oM1/m7b7t1xuYpKY98Ll4neVAmAXfS8B1eZB0B7WUuSAo9aYUnQadf3kH
WRkrNVrahvWlDPa1AZWtbctBspKKlKpKw+Gl00/Iyx28CGkpQCN79eMCNbcCEMir
cUyiNaMYoORjvAFmlMpJewrf5As67DAqiwVfhwdDjnDLte85qh5X4WDA0lqMLMSV
W3cdf3tK/cxHjMlvpDGY8NsdESfckGmhc4ULzwwdUfsoLouKcWcAiv+2M8+L/K+N
5vTFNam/+NiKkEynPUYomhujwAdarqrKChw5Y50N7rxBcNu5ndvBwFsM2uUJb5ii
Dh90mrk1GoGbzsriIEHxlbdBEhwMYOcycazvYVSug+Hhucakns8ZTkCNFDug8d8C
E4opOn6tBc4yTIDtrT3/E+rGxHjB1wCuEUDha6kHldNIh2rNVk9++xPtPLbsjmpT
JYykjNXn2c76Gmd8HgyNc9c/v/JpC7XtXEns7t2jMX0x9TdR3oRWShsMFw8CSh6y
754DxjTZ6GopIExWNWaW4ynNxe2X4IhleP5k9RJlLv/vVfsl8skMGxhP5WZSpu3j
RbjgEo3KOTX/Oq0THKcKwaPGoEpoKXl5nB1XiVNcQ6wYO/77UXKwkcEWkFDzeJiA
Vb6KGUY+IEzC3yjGHZ9lIneVRnZoeuSr7+lVkcmYFoNoRmpnh+qcGFgthxOqzvGs
nPDvgFPaXOD+ysVY8zhGgMPQjogb6OzwA7bI+44IeV46gWOOr9G8ASs1mKsSFcjE
Gku/uRu7G+FXTP+3Bpr0X9ETTw4xsr2+8G89pPfeEnJujlvUYFSfUPVW0IWn51eY
oNEij+gwk9zTGLPZEmmxCUh4HRzFaRzWuo5s7iySMFNyTOHT3t1Vl9pQxIDdc0zV
1Dg6o0oEauM9QYHcjoag0Bb9o8PBNmF3AcdbAjYVHftVsdxqGjRsklatOIylW/Cl
U2S7onh4Az2Hpki3vU1kE1RyouVCJfAISMk1EEwJGWHJd3OQvOiPjuH6OEleEgtq
9+SLsL4psfRxxWyErOZdZPxNeHtX/ZYgknFDAHmAFG9qWl4S9n32F9JHg7d+Yquj
CBqIu9gUS20EXfy2yHzemGjyMmF/tqAg8YFuujcKnR0f1mwHjTnBsi5I9r8E24pD
JwswtEuxV36KX6sKmgnKGbgaFCS+n7/PqZn5+4e66qzFPJ3LkW0lb/5PAcX0dcuU
0O2sX6xo8102YkLU/8zTGP09qrMuB+TriR354IFNQZnjoxR7YBwj4RwN/V2R4p3S
o6aOGjZ/b0GM87Wr/jObUgjA9NAOuA6dPJElrfwCMDnLz0OvbmLb+cyx/gNSvYXv
hQTTOUKTUM56nmDN+VgX5S/iuRbqb9jWZLs9OLq2mxGT3As3C4h995tOn6A6u+/T
yd+zpF6vLxMgN/JPlH9l6DebZPMxwRrRuJXSJOqaHoxyqJX8I5O9WoECyxJPb0cr
HHCr4QMi0kDIPm22kPRs3DvolGGf9q6IQwzhsCBZPNsxTwNSeuvcjBKqBmo2Hw4T
nsPgaFe1qxIJ2/oI5aeCxJyFiGBFrn7P9/5YhJ/ofr8tfr3R0WHQ94r2KiLJYwKx
8a+SoEXvevfiWEkg8Sfws91HPFdQ0VXp47sQSAoS2ue0XdbfhJN8wV8BhlkwG88M
ULpuIolWORr0qm9BwKrBb9MzI+wWxc38zfMDEbl2z/pzMyIPE+Xvi6oRBDjpA7sk
lLtl7bx9KyC+Lrl6RnP2GvZesGlXIQLqdPoxY8nqesDSB+gf+wi4xuSyPDUDt9Pa
txaD11zsRu6V4UW5KVOhDoPD5uVROy4tWVgWXwoCCLOO7pPhIbNI9pm7ftyhA0Si
Cc1llwTP6Q+vWKP7wuwqACjVtH9fdBzsDAC5nLvWrjRm4rgl0t/8KtKstaTTEZ2/
gQJR9hKpUL1lb0Z0KICF7orCZsUJ+sIZXyqKxVewrTVH+Cm3qLMnbafNSsWF4pHT
LddW4buQWQZ1XLQ4i+HQJU0qqKDkUKWP8+ZA1hHcANAPZx38qVKnHSfcuwP5PjW8
12pOIMJX3XC09stNvBiQiRxiwPntgKqXK2U7ICeunVYZKA0l9UPjkzhCCpQmmOPK
fnH2O/KQmmUYp1vAebrsO/x/MmE7Q0U3JKW2CE0U/PU30gq2SKAxWNISAjiDLhf9
++tW0I6o2uuBJW/kjtXKgwjyXIDO6Ks0f1xcWC6TQHglPeAVM62GkQHKG8xYDemQ
w4gv+aM4zfzDffFwcoJ5SimoLEYXcvU9WjOIZDZP+LUADHTAZhtENTcoVd4iNXsz
Zxv13OCybr3QRYyemAXz0+QS2KQh9Fwr7I4mNO93RcdsUw/niWxtf9R/Cr3MF/JY
CNUC6WUIZxeuQS23ssr74d9krVxc5ED7hcyrrIfshq9qDEL/UBR2/wA0WiKecFpL
VnoWFqW/4YRETDFy5MKS2o0bapJArlYMt07UPbTbNNRzUvPiF0aQ4/UWf5MBSFy7
6/BERBG40EFdcLJ5Xl1z7rtNBtpGYM7zcn2X8baG3rM+6ml2YH0gqCHwQRhP6z+U
8ejLuFqVttARi+UcSDt2HxSw+Whruq1TzIVjxmk0lDVbraMZWdxudY/et430eOWK
OCLsu6JZvu219AsrMPNQkrmMbYpxh4KxybfqdyP0dNxbLDF0it5ku0sig9FRdnYZ
nitZeA7oywS54QXKFwIpBo8Yz56nBYqrEpX+A44OjGe5WXFBKNtR2F7Ql7gzRHS4
RHaPM+w1JVU1Am7BhAVVYBJcslW2iH+lnxtTL+qbEgcRvITLBeQE7pw3yERhK1f6
Vkfof7srB7/3xVS2U3099QenDTXF5WmJ81Eji9Siy/srv5lAcA4Xjko6LWWiR033
7Lfd9ecz4+SLDd51M82JBnHVQlh31tVmyL5DrWBgljYW/H+OfWoAoy7dm0y4c8im
KWjWbwq1+eEXZFiUycWx/fG1hciemQiK6huiTbCHFz8wcisrr48QbXBP0HFuEXYe
HyyrFcHbnbrhw4HJ1U+qChRcfYLKQb6xyJq/AVwMfd9eWuTBw9YHsDf5D0FGlKG3
WjvGdHQ2MnpRiSWlaUWpUAKgTAbqdvqtKzE35ekcjoRETCzxc8Fyopp1kwE9sda7
H/TsDPM77eh9NBTQNtYLJlurv3rJbTI+3CjFNvnVcD+pf0MQ3uUuiKC3fz4i+etp
ybSmM1uzq6gfKebYxtGlvBewgOYMbjALktQkqnrJfi2f0iYfOk33NjcKWe8Xs9Hi
XVT/xXi3ZSvnjcm30xLFtmbnMZ1C2LNH+uhfnZXUmzkaeA6hHRqAv84b+5w1jlq+
/wUksDLii8ZjeshYVxMHO44rpliCUdMnntVPJdHxwuE3cBEkm6y6J1WEAOWDLz4l
LDYD8G1qaG3/2tAp8Dhgovf2W5jvQFRxkrXSfeIHniAaVGIRKKfw/UklbWHtRLpn
Bpr1y6vU1DRUykEgPcaJ0Cb74pm7tZoV4htYcNUbhLUlEjXlZ4d/ErYeUxYX73Na
XSur0679bT95FixihFeZe6IvYTfVfVxd3I337w79VL1mE0iwW4Amdx5//IZjM2Sx
Y0sf0AkeD9vfN4cebh+tKxbF9IVm5QiucfPWT86RrRNO5j8Okly9aeQdLhNQ4y9E
rU548cBImI/o8PjSSCtDAVCEgYMW3tfN6oazGL5ilcVxYMHkSgDxley8DqunTYRL
UcrRUab6fyKUwuqRU55AyUMEZAcBCih3KLX0VTwZAELbwoewlwUl6r2ksZt6xi7Q
q7twXuhYMgesPjn3Orf0O2wM2DPr54DOCzSeRsy8/YTd7Ax6ZrNXjIqzIFbyEauH
9g2roECtizggSNLcZeGsJLac6V23vLxjZJUfn6DdyzdbBU4HQG+b+JEXR5Hkmo7W
xO+/jZQC0gkbebnO50F1WUQYbHcHhQr6wK0uNBijGlFts4Xa1MxsMS1oNDDmjdo+
E4x+RkkuTWk34YYgwABHqjvswFij5zeDEaNM36b+PymA1/Nll3b8bdY0zR03p7Pw
EPpyaCXEHMgmv0oGCh3QNlDdwFkJJN02vAaOcugYlUVZhb2kp9dKTuhF+8nOa2/x
H+m/SvjZsjL1AAjfJ+Hsl3YdtQ7Go+glkb2A9xLAbTj7dtYOMeKnG403MQGHQVd1
Apko2j1NQYuK0VNYYTIX1oPDSyLKm+4Km4mbzJbUVpoYiVFMVoMRtjc1z/fp3TNi
z62Ep6utHOwEZODLEFR0iMpwoIxjXSdtRXeqQ9cR+N9IQN5KzRF0AuwoWNkWcUdZ
45p3LN200l1Yk8YluOPYtyJglRgavp9WDXzlLDAySEu78hUbuOJi5Qgkqo9dRdBV
i07ZblBypkONwbsrTzBJFh/0u1AuhpGVJpHvy7pC8ASsobi/O5NWVSV6rcR6x6H0
vCHhc2RY6evRaZ2gh0f0eYk7KMz7KDphJpnZyiChRw12HlsVXiX6PzU6T0F6RWyC
MckAT21uxS7Ibkzj3RIKyCRyKo71+Q02NBfRRN0StnBKFmOxgRcMy5I+swICv11i
Lch8f5ybDfejkFfvcAGYBS0v7asjQsR7SC6vTEKDjyaWJDlSOyfaY2GyYwVXuNE5
tnFncTfY0bXU0e+GO0uxGPw+80T5Ok3GqHdlOr+tLGSxXhHrkRUGagRJbsEA4nJD
IpgeP1jcgd4pLwKvGiAoudacLPHsMwbjbeepGjpl1ACB7azwBU/74iDjPrxhjKvW
88pmJHE6OMoiWlKJKqQRWF28b89pgivrymZ5etg2YcYjDj4mgAbCaTRwyvaFu/yE
kGdkchZYHcKl+XLbcdHzuOFME/UnK4tzvSQul0dYvzGoZAbBZ89UIjL1+4HNj9oz
GtJvJiRH8Tw1M7pcO6SnXE+lHuf1evxVPQICvOjCVYCHRyvkepJn0+aQZsxj03WB
fNpOijLkZrd/VsO3rnJ6huw/xX33yf8FNMlrwVgD5uQMniCMNkwEFRHiBbQDE/TF
CGgG+qiXkpznz0ieNAunwsmxN4WG8XoPZ3YG08G8iPX7KncZEiVrJ3DFLcnICgnn
E9jwdEna3JhHV78+Qz7EgNbVgaaoYlMB34iTVMeXbvNKIyn2exeZy2A/aRoDKxDn
p5EvbL58oYlyX0clJM9AFq5Xp55ux265IvF/HnyEqio4+CzzlLotZqExoF6ngLcR
mOtuOnBboF/BNEM0FVnCxP0P56UAziXyV1jfoGzRMylFXGhH1XiV0bpWl/pM1TtR
Roxlqqym0gvzSN7HL9OH8AwSOm3NhscufA4vzUhIF89R4eUIJFM2D/76CoC/TUjS
HtlywBXhFTYXzH4WxsZ00UEZbiQs4vTz5M+gfQkk0yCH+sC9ulVtNUyYvrbYq3O4
80CXRsbo1HPEXY7DNxMjnHwEbXqU+CPNMPdmmFthczIEUGxCAR0NNe+10hk58RzR
NWf0+pV5N+UrbiXPQnF58z1LyM9zOzd7hyUsPkJC7LFIfga4bOuDiABQUs7eTGkc
kFrFsVA9qWdzaXeLHuhZ5rQshuIEdwvPQFKz3WYoUIw2H8b9xb0HkFqo5E+WjIG1
KiOy/is0JVVbde/fwBOS0yCMaCaj1MNKzZ3Tggye9Z0hzW+xQF3g4jWpMqU9tU2Y
6DWyq2OyXg2Eiv6hugUx/oo6e74fPDsDeVMvQ7p4lZD8pB0ZRVPrfEKyuXL6oKfZ
YNYwB3Yxj1dvDOHig4zPjGRnjQGlUsWgOW3PmqqlDMVcgwvtI1bFFotWkv074zLo
9UM6VJNlGjRpbENpzqRUzkAWzID7xkSqsKkqy5mifchY/WBTWml66fJVsCBrOQbA
1iKhCruPtTHDXPoku3xgfNR5EVRPtRN73nkgImZZbpmts5tYni1a0hO5VNoxvoWr
55/f6yeyv70IS5ZYSpSzJ+EjvAs3//1Qgx0FrYGzpE0vC1ZVf5nsXlmb+UgfEoD4
NcjtqZJ3vvPdcONh6ZYyYooKWhDifzhfbcUIaUqYXsspGCI8pGIGK8zb7emFWcNe
kTTT2WZVssJabaW6gPF6J42Y/Cpb5oZGkZwiVWcYxsiTr4g/VmJylr+tS8vM/T1Y
m3VANluLOs3zJSsKZVONE+ayTRy1Bs3Lk+8qzkL7yAJJ8Z+XexcDTvY59meEIfkJ
paSz8fn/4lCnRDm3Xcljl+s8TuduVOb4+PLU4eUFkJj+eBAXNXpiQi1/MeQsBLEw
/XHeb0QJnNPT57LfAvDk77AJcaicB+jnDNS/tH0XF+T2xfm2YZGtbsWH5ldJDTKP
cJB3yOIxVdn32GGh18lm/wU9FCBcCAn1BhBYcq9CRMK2eOSkH6Z0TH6tsgm8s5av
LNsv+wTWVXGYz4rAS3rWnBai7alROVNk3wdLdrt9YhqVczH/Rk5GFKv1CyfvjStj
+BJ25pSLoy526ZckAhWENHYqS3NRNq7RMOyYjhntvr7MniVHi0Hu0+R7y4yJZdV7
rYOyoKya4+mSX+K12WcAKq0n4eNubJKC21DkZOTYIEIhIVajG5YSRVmuC9M3CjH1
NnTh+twiMcxh2Qb7mz27mhcWMkBwR2/jEgXRZAXGM6ud/zj8yEYw2h8deodr6Znl
X0jLNiMswGr8KYvR1ZJj5QAJLVaxN+eHdDQAzrOoTW8zZtx2PhLPowxJiulR6yvl
czrkw2GJNIe3oMv5lzT75RhMMV8g0c8PuKbIOAVW3svYs5yjQ5uCf2Rt0Y4E8s31
xsePZpukGNagLkow7reGcBSGstzlwgL0+3dqO8yEP0Y3uWQ3T11daxdFfiFMwPr0
It0TzrVEiaIh6tW+trHfow2PVhwFZCcCREQi+Ci3CIGXBPpfJp796g+5ljLY/QGd
J8WHywA2ssHlIAsoARy4NW/ylM2FMbr1S1Osr1VrN1oyRQkYqlkHGAktXlzKgZ6c
/b7vxT4YEaTydRSS6JxF2GIsBrtcAQKnRIgEzwQxm2FFCuXTvBC5RjM9OIawrPQr
dKvOnl+09/lBpAaRE4jfztjDrj30/4tvnlaUvsgwWhHAxK2CEEJPWuhtQCUJAjaW
e0TqKZ2AE2ASeYxY6SxfkpjKOFxPF8ZkOop0HMp8PWGrzEnpcC0me+JXCCrKiTmD
usSiS/ieD9O/qNq38OmhZwirfC2Aw/G/sb6+5qseOCJe0EETtEbAv0YVdnOmavZL
/itJ6GTfGTBNEYh1/myEUPE9sxsqJGhct1qm0PhEOdMP3+fXJtjO/I8QfE+es1im
s7gBQXIc7QnZXVrWXVNkMdmweaQirHgwZ3Ay22M8/DqSrR2RZzzVY/NaG1c6j7Yj
9Ra6cLLdCPxwMUV6owLK7Gft8iPfLgkm0PTisg0cms7TGFYgr17nytCfdg3bHniy
vj3+7zLF6Nhd+Hoiv/MPKYGeFzLkOwjCg1PDAWMVvc9hwO3uCKoGtUUKJlkCa1jL
erRDsVGVnvj2txAMH3573MjP34MlFGMebyxo92YOlinzCkhHpBssxXqWwYiNr26w
gKch1HVOJsR2M7xnhgd/K9yRvhgKFYpCopxWZcgJOYTlTAgZ8pHBWsV7NHKUPJ9B
JPuMVnQuYYPeJTt/ZlwtinxTCkvMkXawux3AaCITbHB10Mg25QfT/UJxRrSXGRi5
7YdCeV7zBHUcTfq4GOwGG4r2wBFMEmYOZ5mz839OkBY0Zp06GZMlDEoUz0KoIlGx
RTRz5Jeu+aSwa33lNdB40GOM39fVpdbhuVdG86GwvCidzp/KhLmQp331LSYtgxWY
1eZlVdTMSacs8lbRvG8t2acSGljturOKlJqENC04+0dW9jKPxkQSlisf1rb+54yH
KzOdplaQLV1qAsMNSwzLCkA2s93+2A2uVhtlxVKQnemuOZHxBXORO6Ru1/isvbis
fARHaVM1pFceaMlBGP5/99azOX3Im0t21VsjFwyMo3a6xl/NDC9rX0gsoiFNLipy
uAXJmNEMo37a+2GKiLsWpvnoCoyTZrlrUyF68CqobrdUyIIt1FTEHUiSzeM2VLdm
Ys+aRO3snDuFv+52lO0iDAdEB25tYaLdbJh9TXdwZmfs/UnSsi7Bf5kfst5F9uaw
KP2+5JxrmbxE5LBOR0sz6x1eCVckvD3chYk/b880KG32yMVU3etw2LaNl/2DGMLM
B1ULCKduitQcQGCHt7qtdMRWM6kIX1nTQ8VJsX+bwhJ/1b3VlgAI3ha7gnSv747i
sNNdrZrGFpbK9Wt6KiNLeAjMaROVdWDUPcN9/0yowlsuYOsRgwibUeMxF5xp7LkA
vaFdgaN22q4meg+dh8hv6XOPT+238ymBi0MUk1qHw++fgdqBgQEDHDUV6ILzknAe
dH+khdhR51VA/HxDygYpIiYEXkZz2oLiCDKJwfGBOz+fdNofDxSF/3q/rC3lBUwA
JoEwLL8d7lOU++SkWi3WZXY15FJ6jnNus7cQdsg3nmgaCXwsRQgwSWtrkB3jCphS
JrJ7ge47Fjbirb0UNrnC3Q0gT0FWVemrN3OHRSH8opYuGJF7X1NgsGACOquTIai9
jeX4+0VipC00eU2ZxwR4ftBo4p6P8ka1O0GjiR4qiF0M8rMiiTpf1epyZd0TeEp0
PQQm0HzdbRTrA3cG34Kg2SXfana9BF+cAV0/IXp+CCMtdOoftkTNL1C5twkW99cN
9pu1xT7OuHR4Pa61K1OOt3oDONMpSWbkanAngOyIivLW5SNaPGUKegxVQ8n4PP9Q
XLgbPPIWst7cc6f4pcck3gEuiCFpnlguOfu0PJKw8/1x4aKyQwodRUzMiALv3tBI
QPd1BmczIEhflGAEV90qkRFO469sv5ynKKYtLjsTwi38fwlexfHBkhvWP0NzaWg9
hzkK/5iHSH6owbwHVAFFEiYGS6ImEcaNUB4TD2bK1IOg8PP5rtWZiocm8ymjJh6R
OiYcXhoh7vPvln/fgF85XstQ9d/RczON/r7IROpeWfWFXOG/nhvebH1yzDqIqRl7
SPkyMLIMd6WLzfkPxDwJpuPb8JKYiDgfCbJK5ZKiSxYXItUCbfBOwPDGh6imn2hU
Dpdb5lJ66q3DXDB5rfRaJ85SlAEkL8Wotv7oZbccjYiu0SBEorXE5hm5YAWaTQLt
3NU2e1mRYcT0P+wMJmPhVMHlC8clrpnAun3U0Q7e8xIaQG+ir6AWFAAWkeItPBhm
dCDXxy0A1VmK3FyApkYFbEFZaSBsHty8IGWV7Y7zXCLVjkoa1yeir3hh4gY1w61t
WUShOgTUfOSavPrcLSdoCGEUOR0b5kSE7CjBc0KCCcFH35MgDRpbJny4iYKHbDPl
4DmUnzxu6dHZeWW5pqc63iAD5rZIkgrX8J4ex/4DaoyWdt+g/sARSghD216PJiPh
JFyeltTYnXRjeKxh1MRDboPv7JBvIQZwPtvX3fUYzagqJETcKrhRlc1JMOt/H2si
25+gCtH4vcIPHl8lE4GQqee+BjeHy9g5pB+YTecIsrMJlnIqzsWIYgJY40eJrv6h
uWC7jiT3HXI6UDYC+umtLCtMk9O95IaCNSxNI34xzmn1IlOPzZrIAcQcSO25Mtux
4mnW7IF6PfqVtMjYCPe9pJdeKODSydRqTRYk2gnzKdhEPEoVbxDJaezgJnc6EhHW
VPxK7zEO8a8m1WYvkwCVfDnR8Mf8meIH3Rfx9702dklUupaUfnSJH/51jKcUjE+y
YHf2h04Zrgklb3dqILday1md10r56BiTQlWUW9I+FnXciYiGC0P7N0QMOYTPba+u
ae9Z2laq94DIzMyoOMrbO2Bo2XqqFJ97YdSij5anfDMxDMN9w6+CvOsg43TdMlRt
o7nKz+mgILpmLq0fsG/3ItCsZOzmRrPUnGocKkrhB1SjOFiIn7wb2ofiI3RD53kZ
iq2wa9sW2E31VzFNhoRo3rwmbTY+ydv7IznRHHcWGkEOH5E+NXV53uruCPI6sii+
tgQbmTs9WKL2OGY3g1GG9BzoB8zt/JFUCUIGz+PPpuYHwjM65eCoBwVhVUXB1P4v
vUn3dfw5qZoS1+iMYTC7vcHLMG/BGoDvCf8Mk9F43QtUD5gi0xTo4oP2POyfDNkG
Yo+WDYu+KHPeMY7uYJwQsfGH34WRRAWui1JrDjqYs1nz9aouwSpT1lzbfT7x4RfC
w4Cvtpx0wY1VCeQg4J8hIXx+4CJQaD7NYC1cLYPR5GyrUbynn0wFkQ8CSyGygO3l
JLxayUzQhonXxzt6d5xn+k4m8LBRvzb8UZD7cQETgJKPRuusdbzjZEXuuTRPuJuX
PgspPjyejeewXt/tX0FKH7/W+XsyZA5gHboAWV2KeYIPYInDmKxFfhQpwb/Nvb4+
Fv+yWrmYGyvdwYhQpn+I0EOYmXlKcjN/sKSVgiKgMu3DcGPFAntiY/nIJD3YyYv5
HT/xQbSEmuBSEff6Ag1L7dB7Na3wC25i0QcfBDPVj6gdZolmMGmn5dD5CLY/3rnf
Ogps8XrfVay/g9rq/TJwmqpwiThMzZSplG2ACffwGGeyb408/1CYGUPRtXsc9Ldw
fxaH6R14RNNfgzr24kY63tIos3haU4MXmPI3uQNMzb5cu0xdAh9ApSLBaQiwJJU4
qa0yCvL3sPAIruFD9tCrb0H38nW07AvplmRRSIb3gxCEdAD8PChfcpRPpCw06f86
YXbDKBmZOONZy++unfP3qar3jGZ583suJQhKRrAWzEVU5bvBmQv3FXn+k4qlAhXb
IxmkCQeWSjT2rwlO+FChicPtiN2f0TJlumr+D7Ik2UdHvOvKaoCbwI43beMVf2U1
2AkD/VTs672SfjJDlLc5dNLyt6HaWLiSZ5Y4t47FWlgjYj6F9x0/vqMTHDXXYJTx
x4wQm/s6mvjsbA1HRxUBZrjVVo1pZvSzpzre7LAJjmwWWFllQPOi7dhLYnFEqisN
5CESpXj1bjjA+n6q8LiZbC4o/CoN5sZBx98sdL4xApAganBZcyQbFZQ+n8/Ip3ce
5PZHZgJSf4NIATuvCvnYLStpWwFtUScdLASvKsT0kGKS5VabF8Oo7c0qHGYVcnRF
11SG24lqz/tLsWTxfdi+86JTJ50z+YR2cYXQhsZjzfoizgLMBPrxNCqJWZG690YT
D4slskQ53F2JyjvXfNS0Y1yXV4obZKlRfUgudtAIP+6so40i51yagczP3GCOJrj6
9S4Wzz74hAlbjhZ5O7rAt8e9BTKHXiVodJNiIx6HtK93xZ6GvjGwbTA2kDlaPXiH
aKVcNKpMLN/VVGZbuH7RG7b4pf39q3rirahZ4ZZcJRGVnEBeFa7lc+rB3CigHaxn
3OdgKX3GL1cCFtFICazbOtj6tEzI2uqAzkf52l7pdpLTj6CQSgyvUx7TLfW/WNJ4
XdvvNZCuFfD8qsUz/ti8LMJnE8fEZSiS9Cjl8i+IIkrFeeuLKLSK5MZepX/y1WSO
AYZJ+YB61tuQSWbLsYMnJI5F3iGKNkzSIkeO22LryZAL6A1SRQDrvndzm6hLC2Rj
xP0q9KLA4G+DhQuUA3A8jOYaD86VirLq3XHMbtE1Vxz29Nfn7EN+BVWIz/q0HcFX
WuBYPCJowuwjc0SzETno+jxHOqi7FEfFKp1M0z9QnKTqYWwVWsmOfOqj0TArtb/A
JyH5dqWXWb2RqWZgI6JH0ayOl98k7p+zzbtUfMOSrHPt5y5EYwjk7sIkkqwxT2K7
IB1litXbInGFQkjME/a70AoIiypPXBFHf2U/X1B98U2Bm8U5JR2NF8j/FE80P9g+
6wiAOu3whqJ38VAHstgoNy7t6bNBRQ/qkbnfvQYKUAUNaRORLip/Oo2fxLY4wPvZ
g37g/vT1UW4dfiAy2PKgq86lGhDH/AJErPVHsRphcTbpy2Ahv52gwrAtDqzoR01e
GAZlHT7ZMglfbuq+WFprWoS5jJDvcfA2vS/9pEtk8pyxy7C6VLn7hU6ZQlCN8SJK
HUuTP7587A8LwYUP1mS+duHKZ4R/aJ+5BzUZ0jhZI2uiCz5VLwcmTAzZP01eLALI
cuBL9QvF0sfy2qygEOV0aEEmDYEW/vU/tUHE3x0tINgHPhgHPfLbCWUC3jePsjJ/
ejFTKLOM089U41XbbcNEsz4dNJiMWGAZJ9CAbLsG2lxF4Ow5dyTSA1moC4bw2DX9
ijvqVNFsYJvx2TzdYmq4Q92qo4qeW6PmSxB2cCl/hPmSUfXnHfeYdXe8KSxaYRfX
EHyMDnRVbAW/FqVdSedoIOQ0XAkshQJD7S0Z9X9F4ce882kLdDGb7w29FxELhvbe
F6n2FP2ccS65wAEG3M1dvzGigTaBApAP0CUlFish2fETpQGd8An1NPi/Jidv6n3j
gy6WtYKcyzxkEddWB3p/abn6bh34lm1JvA0oO3KxgLWyouUA0BxGM/1n4j168azm
Kp6T2EQcm6jOougHN1xPCHcaelO6OkS4H2GTz4vKAgKOHmlkBTGOlAFfmE7VibEt
9C8pOfNF6ESJ2LYR2mcDUAP3IbtiqXmVMcgLenxaMltrGHwjPd79J8vFSCAAM+G+
BFxL9a9bRl2/XK20egcJVky9a0umE1YRaFW8kIyRen++XFPcQ1cn2TnYInfZQXdT
ylPzaGSnDsKqxLeIyghTvJvegRV2Un8kseNjCxYsZV2IVaXXfIuoWQhKF2KTVFuW
WTiwsiFV5iqtpKws0b/qKTp0um1wQz9MR812jGpaBu7ifkM21wtuYmM4zxucg7OF
dA1f6r5e16KojDBGBq1n/F9ElwyDNshX1vxnXyJJCxFnt1ppTNyZ3MwwyFapsKYU
EXTgx4Mo3OjUfngux3WGBJeLlt0KUpH09zLPLCSThMTKhJ/Eqc80V2OQc7RTkgli
g5vGE1ZHC5po6YHLpznM0BIRHbHLc9V9aUE2myMoURPCh+GvGVDKD6iEPa0zaKuN
F9mYR3IXWMrfgeo6enzOUIFX52IXayjjEA8GnOzWUkCfkMYEwVKrAjirxd28Maan
TSD4+SuL6JlTJwafpRxYFzjEWitwDvkbHHAeHR5w2lN6chwHf5gfvD9AB3vBLg72
PdeJAP4GTNgYEqA7vOmT0ei9MvTcNxIVIEFwVMhPnNJg3G9THBAWLSDdQg5O6Q4D
PbRjV8HwpYC+7eWrTXfQlEaKkJDOWpWZXYgj3BPLgfMtt5zt0sTsm5J5E0NVBk/N
Vdl+I8907qNF0qlAzFqa3BDdopsDEDoAyGdDuFZyeO/x6O7e8lcukc04UQXw6V3W
KGOWS80gDsgBugUwAOMShIZfFz5rwMRCgU/uif54cvv2BMhODAkGI3cjZbnwLvQl
MNH+dfJcQCgMy7uLe5ShodEXCdJprl3rPNZr4qHwsfC5U8Wuit+588A1CkrGVf7i
6jXQUWLi2w7rs0LDUqE1r8/wLAMpTSGPPi84Ky9S5XYLaeB8KLf6z54Qy9zrxSGF
uBJJe+ba3BW/fwtMD5FlkldnruJEiJtoC3/R98s06sf3C4/QvqMDWwK3ZQebivu1
7hXaECCnqpLs+Wv1uaHYACJNxMfU05RnbI0laZb9bJLwrunpR/K/TuNkJGjM6lgv
xz8tKo/CC+iuiPBKJ5QeIaH6W3pWjJl0fa4s+BTinCAIAJrO+O8M0ky31dnujYAo
876Kzmlzy4wl1iBg8pe8CvJWU2yJshXnzGADxJ/sdHyq/IQRUTWXdtGQvoyzXdXH
Ci7R1QulOkY7FLLeS4zn2xwA+vMIuop7o1vBqT++q5ws4KVWRg0i+UvN6sgKKpi2
9i53lGuQ5S5s/oVsjXUj1dk4c/LtDf52eHw8YqSc+fPBhsXNoARl8QWAeiheHX1r
e1Ulrew3LyH8VXW1/iVpRV+AYDMI8OXUtLchzFybDhVxYDeZ/hb1oBQBKOyzsbRH
Tc3R9p6mNfq+GHjI3Vic7a5CPJA2jDx6Q/oxCIxFYi0yhUh5vNOWzSBEduDqmpcj
syajlodJY9svbrNd3HlayqutyZg9RxczdBkRYGM3XbCCksBunw8nWyaG7NLefg/v
iLVWIcsro9KEs61iFMHFRCP8xHq0D1o6Xaa7MKL+a4zk8vGLqwxxudAV102rIUvg
L9rR5NhEJO1MtNAEzvCgEg/ZDuwLDpyhByGWkl07hvra2gRMb2DgK4NCGJnITqvb
AN6oyd7NcdYHZCts5Y2GBzX7qmBvlagcPJYIvAahpx6gXZktaeJJnYApzRzaA3eD
IncxbVPxEAYmefGdHk9BB/eeOa13/xY/UfN6V55cZQMVR0tryWeG5CVT/vsBPA7J
rpFNyh1uT5DWl+7d0UNCk4yh/tSdVc1AOrauxW8uYvJHmB04v5S9+TCPCnHR9NeB
TaVeuYLgfCspXRbLX0ADpvCoXPqYCqWzosGxzeZZ++hyhq8KjMBlKEja7YSWcp62
HIjki56FUmi0fuyajvqarXqh4LwC5IXHdL/8T39Xpo32dC5AKQli3ZpoWqdpwZFS
i4ZjzUnAVLQIykRBQvldOEybElbqWVsM4hSYI0QGTGGw49IY0d2gLqoo61g+Kfic
gwiswuMENmr911LFHRYJY54nUyu1sc170k/VzCiv97i9UrIOEygsWGNwnIkdgGGE
/oZob8b5leBfsfjIcFCYmA4AfLgYCnarqL4zl14U3Wc2s/+/O+eHV06EHYt1ERu4
fmQ357ghT5QHMA9dPPTSr/VIboJAmpGLM/uEbs3UgYZHCFjYM+wCs7RkGdAeM5pT
xGxDDF+AHWikahfuUlXV109/0hTDldxeTP/V3MJkQudCyqNUDIvuDE10UBxXp54o
UkvcvtCtBe8Xv09MpCNRaM234YkC2eRMx/l6WsGdw/TXPR6xAki3JASOqsuYKBG2
5A0PndwKvBl9lyA9zH7PkhGsyEt24LjjapjFmdlukAU4s/nLvLl309bUlRINSa/o
+KSFEF3siUUEDo6BAUh5MpaNhBuTrueAx2osGCfO6JBNJCVdYp1N11/uYTDvcdyJ
DE8Wd8xQkL83pPMKNGi9eJ8z0uT2OWLwOYIHcpNXtiVwQgpAymjD/XC98367FkLn
Pw00Lu4pxq+9CMSGL8hdFH/0BsuhhhOmH/cstY2YRm9Jc4xJ8DCcySInBf8FPRvy
OwAmHyT5w+5gnz9wZDX8EFofVeABX4Zz/f6/n64QjzcF5GP6tuc2/eKgnNSsaySP
jUiTlNzKlmqG76KasWnOrxjiDSawyO+H852PXhGHzdBfJyDc0TIVYNPRwXECxTle
pXowXsxgndMt7/qkIgw+016gqqhvE9je7xkRVwd/IctuTZ7meMRlWIUortLPJWDY
xK+AOHwvTGFqYbEVOI24UvZI3MEhrrJWLMuH7/NprAdLjiRZXaCAck5lxmYIfZWi
NqMaGDxakgJjLn9wpZCAExBUaqFfdLCa2joOfNivUeTL6ZWZh/uKOufVcLCbKdwt
as3cJua1xlYQpb/t0Hw1yCJNYUwMGqyB3TiIvlZzRmlbC3ZjU19tzb6pO4eW2QkE
ty/0ZE/taSJL0Rx+fr3189qbHXz+Z701dul+VWnFVcZCUiOlE5pemjUIOxg+B2pB
j5AaImTMzGVZHCFsj6NYM/XCsCPM6WvbWFpmZdp9lsF/yLb6K5BKhTkNVRAPkky+
augdcJVcLzpkijxemTt51fji5V8j21wcE86Ar/aVGZjkGKISkSdH60s/G1fnKeRD
H+Os5NtdW9PpFJ6EPxcbXF1DPeIehIA1ruUg3Qa0TRenw445mK1QxyJ8H235j++M
SkZFgp/mrpZMLqLjTcmxJUqBqT137feAgjgpiTxQ/5UROiciE7abF1nBfPRQIkYv
jB4W+Dy/7aVVfjYY2Hi5BDGxBddIDzklAdJ/N9ueHFn5JgmnwVmgZ9MgkMyqd1lh
Ze4tO9cSlWLlvMUCthANt8iChPYV6XsqpM8K545g5Sg1uw7+zO/zoAwVcjrfnxIL
4LJQLuqrDZAX9GvrkNhGH3fRCghQUDV4kNzxM12Nbvw2FZJt05RebALgQ5l7W9aH
k0jnBMj/N9i3glOYw8zNkvcrxlgvGwtXFD3CPGq8sv+2CIpjYmzSo7oD4fzJHtjw
0sxeGqT/5xFBJGKt3oWgY2QgSY4KNOlYOdFPzVho63gOq/xn3ksPqH/LObDvqFyw
R/WARqwljkG55nu2eVgwQcgjD1AzcuL7J/ZcWIm7trrAs0YhMC4+zPxzbQRxBaMm
YCPPyyWNu/VwybPDk4FFFvL1lMQFhPMJ/5826gD1ymnUzaw2AhJ+7SsYyY6uM1LD
+UOT47yfZ/T3+S7eHceUAE0sLdIdlIt7L3+SIUIU85UzJOaZJfehdQXSf3jQAU6z
J/h803Wufj8Sf5tuvagIkswLnhRxzzc+d8KMiqq5riCLDR0Yc+2x5VnkCCqQ5sy5
B6bAbUbg+GJSXeYkrEU5wC0SewcxJONsRpRRhTg6pqodYY38jJhnv+9Z5zwp64D4
MMzawBjZZL8PdOe1W/gZ0XX1RXfcUx7AelWozIREj6UE5ZX3g+gNMNn5tG71l0s1
xJh+ck+W+vdA1gydsw8Xbywh71d0kb/OdTTSCjVmAvtALR6Yq+wVf1Mh685HC/jg
YWqEM9aidAxK8Xis8OxcbJABUIo5aDq2kM/wnLcaJ2QCaFzxFDbNc+TOEeXohnyv
PTwdS8WHaJL29hWTPFVSRVWZixLrsCxH25q52JRd0M7unEn7Pu5zJHz3noTlM70m
bzs0Pfme3MRSENIM2V3MaAPf1tpMsz81FxBjY+p3DbmaI3tVfC94CSTMRU141Eqi
c4Iy88w+laDjotUL/dM8HXtmg4yfzxYwUJEatWCUPAu2dFxCIvi0V0rCjgtKIydG
5S4I9jch3NJkgy1qMqU5Ae2bbWv0a6nJ0huArpZMmS2I4N05dCjm4h9PopcdIF2m
2883eMAh8CPf4nf8BqU17/rUecSJLtTHTALP7sB/GD7voXrvEH+kbMuwDUtzqxqp
pNR/tVuE0VS9kj+BjcBWtHQk50aqngaRdnuX67LJ5mFesOk4+y3liUHAxObv3Q8+
lPpvhMyLpodmYBY2fuHDyntUQtxDPmmIE5JkN+25+lEH1d+OerkwOX8qvdsXVEka
eZkz8QHst4V3yA9XsN1LkEzW+Xn1oFecAUGmZtS/fbi3dGxZBMT4f5WjvhStO0gZ
lVWvBVDDDuRYJdDCjURMKUdGMXqdBVxGtl9JouD5QfYT5jb3wBz73T7wmF2MyLqq
blJGPC8ukNm2ZfeAIF3/2zAb2FitoQ8up7035f5tgDVFoh5Gi4mc75izFV8JBlAa
zCRYPF210E6A12zj/yp9IBbMLlqtNJKp3IKSsV8yImLchHVy5DpNY9eODSsW3n4T
adLfXbKZCIaAy/lPf14fk6F8upe9+uf5Kq+XzeTnheLbmQmndBqxaD8mP0ZkVmN4
8RHlfUMiImVp/Twpv8YRiAZAatCMlYK41wkx7HmYmuhPzafxqxXef06hNUeqQZ1R
qEQoHwdPLvi5w8qcUJ1Aca6OpDkAuUMyeVpOZfnzYEZTU8XwFYWlbbcDL7AuPcgQ
LRs4m7qU2ft3L8mNHAlwvx0xK2X+rvVzIHsr0fz/fhuD1Spk86cPkH1Je5vOX6Rj
+KDka1VQYfmFjriuGO/ZJZv5uV0zCEBiOEuhWf+8znz5o+NaHERnLRUfAylIhfQH
Vd3oHB3uxsT35+YLT6QkQMj8KICYjkcCtC/XSowVa40S9bXMhtI5Zz4OWZ+vvklv
QVzfywshgsiqTwWUyTidd/dAMDhfCcenvpcBejR9J6wXENRBQnrHm/b+6Dc4U0+A
onxdZMaV730cj3gIMFZXA6z/uKEYYESiemMtBBUvUrN3vhFfQH8amJko14gVVpme
hJJ4eH9cnB1Kh0HfoE8K+XpKZwQ4Dbni36uofUts2dlT8pqzCKSQ2N8Vc5W3EhNE
DfISFZ3JIoqgOEBNCGYA0Uh9+iPcee9Ea0vN+K2jn6ZVMehgovizonfTrctII3zb
OWy4GKpoteom92lJf0C3og5NC2zSoJdP0DuP2yv11xTiQnGGpZKPdjA9Mp3gbsmH
iSafoDThyFwkVyZVvCZ1juqyEj2mX28Be8E++bOnG/COH60c71naxfd3dvSR8DA0
uM9ES2CLhqjMk6qVjAOvsx04A6tM2Zs54tC5JaaJsn3xv4/mybt8G/BgFO9WDASG
eNYUIyBnlr/7jpkG1hfGAyHf5of2v3OPpfa3yeTR3KIi4ezuTsY3fp90IWBsvELI
w7cYxrufPk5a25Rd8aDYoEAOUhNzfwrk4WKK/JE2Qy/hqOxEvChv9ePlSASW4nPA
bXdGWaaiafHVS28K1DaC18FfaAAPm885lwvDWSHfhjv/TQVO9ACRUGg5j5i9kjGT
xvn3+TeaPjzH6uT+R+tr0siPgWWhBqPuMPMpIZijUjW7Orc+C/m84SxVzcbc+JJp
OehC5Ld+gceH8vgWwa4DZSZa69xnJsjdzbKWWK0TGGb/Tnn0dk9GjGqxj4Sq9GO8
uWQqeRXO2vWXe18Te6s8mrbVeB+MvspVBvjWmsh+k18UxJ3RNEF4oalaKe2cxrdJ
VymHqAawLfiu387GlUd2okBtJ8EQMtjPB0+4uXOZF7fRpeJ0HkLqe6ObCkr/g2u3
AocJnyMJ/V8exWaj/gbXndY+V5s0A2fawOs8RG8iz47ejpca0O9dJO8ybWZuxezu
6DtWVrntfK8IHtNhW85C8UkklLU76cOW0gOFhQzPX4M8Xc+9OjulRMxU/o5tiKz0
6VxpgUkHDL034bOsJ6AQgJX0ZI1KTv5vOfweHZ0l0WAdzCHiV/YKdWNp47Fbu8lY
9wjlLXM4PoQR7Z91D7/flDiM+0xKlS4SB/VuFQ+hynJw8jPXmdUXlcS8aKWCO0Xr
r51gnSGzxoeqfCB+nldcLGWELG3/DvaRBY7ssmz+cerE582CsZa+1tGhq8aOS0uJ
jsDf2AqY1erHPiviVhS9z6YXOqUT6dSXGwIzbD+nKY8Ut5YFDtj+UnteJdlc7M3K
ytM61QPdT5Zbij0jxS/Xn/yS9+oi0YleH4ZjNcK+fpm7/qYJX7x4USf0phnRYOeq
nDpllVetDp/mm3Feb9jalorZKhwjV/X2FWMGIa7GxpKkW0G819HspBAiM0ykDFnq
Ghh3YmlFHnY6QBcNCSiIiBNYV5Bi4hYq5i9BQ/X07z/pESWc37x/xthaJ9Q347vN
30QIHVBHfrKCV+sNNCqnBsbbuHH+uLZmbI9l39t67bAHw9V5BezIxftid0lKNi8l
RldDxHYdQPl+iWb3IoAoYy8RTJeJATtf8+Nwey3Oki1fu2Wzt/Lc86W8hx8srRtp
pTah/cUqr0cMlUoSI0Yjhu5L1pdAvDLXELZwzCqHVOfFUJaL5JM59egIgeEhApMZ
jy8Rg6yqIBCBavTuK5hXIYH01bnQhAwuu8A9H/0zWIARCWT8whfzVAim9J+hDsyW
Br7EEG2qumG9vG9S3TXUSRCFrtL9x79XVGZ6CJ+zJGY1E18had0NTcX7u4UEIUQ/
XtaZzaeJZ6my2ZYLm3rgc9DNiCTdCF4orZqIU7rj2Zwm3S3+Dcn/h7xE0uzkSoVk
4QZGC2F1zyF+3tBZcMwPYSCYZ6eNLWTJkJYWRHgBsvw/ZWRJ+np+RmO8HYlH3RYu
txmODpyKWicaLaI/XSjtxK5S4tmZib5ZRtYZ5pjEEyg5XIYcT4l6t2VVvRwbjN/e
6d1lBg/4ORwvx/8xEnojkxUbLgkVFpwSTXmRxlu15d6KZpw+6dnkcmfrs8Iw+KGu
pxiSElxyisDCT14j71rlyIaMAyO3uZAthJcCR0MXfrhUmJdW6KHDfbyerkiyBzkU
bLjfUGR1I1S2yWvDnlXFRdEDo6bzVwaA33bqkHSFaqshWTDBKkAW8y/lfDcBDNxG
CZyf/SONBh5GjjjTuhRnT+9gdYMCpDjLj/WJYQn2TzvC2eAMdzUWJEe+VSgcbThT
/c2EvNUIh7/U3pOXU8IJ86XtiQ2s5nEyUJgkwR6oF0YIGi/BFEsdW0TqC58n5awy
TbfB0K1vk0eNayIgkyNgk4mn0pRXKAWuC/yDKB1A+nHg1vnOYA8KHG4Z2t2DGbmE
RNXvOgM+xR8lsplTqWE7+bwsSnxOpqzxfAUhcXfrB70vLEL6p5DdfXiGYWLfMz8Z
R51I7UkwEBjTva3vu0XdRJm8AU3FC6LNnr1sgcmLDOrVD6mjteB2wByjX1lCgPgD
6W+PciLIJPVVCJpPmi3Y8W7WV+kIbFa62rQD1cSbhwm94uSA8uaZGPNPZbCQwANr
LuyTtePdQZzIMkvepGQ6idQfg+VnZIeL75g984yn1HcAgf+BXWmjVsm44WlIlY5r
657dJK/G2cmqDsShW6zKmdKcx5gB2aRhhGu4qffg+nje7ZO14f86HR/zrFnqWL66
JStvuuQs0HdHvUVXGLrwz8uPNB1RwgCr4kghd9EIB32HBUhjCjy8KJlH3Bqu9vGL
O+fstNvEMWDvNhrpWgXleMAGCE9E6o/x3UaNAThcIVd4r/EbQbS428yt0agKrtew
KMp6JcSlQstHsO+jgBE8pMlKzjbpG8dhZSRGmKckql+Ez4S6Va+gf+de4qpELguG
ym3wfRwhqNJ0VGDlxu5+RdYyKG7zWLT24P8lkU5Z47JFyD/pDRSCtNXwteu5VYMa
BeTzPltroUI6risbTgEBVwfmj5nUuLKW7kijihOsPJOEf4sC+qwI4f/EhygqLV5B
IbDyxpEeazDaoanPvJB/Q/uptyOnx6AmMEuhdfQ1dfUPp4GNHHHx7vq5eYtRSXYU
Ogpf82GS87kIok7sHifamAGGPMchugMNhQVcbqcDbquq6HaKTk49lIefijL2GaGo
hxvoZcte5ENfq/L9gJou9o1fF5uzs/Dflr2epMNZZTXGjFWj9qGZJeSOpJ3VPObR
ncYd8BL5HOVi0k3BV6ZzIYlbabh5P+IPnmidlSZl+KLDcFiQ1cLN9TFayfpCDyLz
aKpzHbEM1SNZwIXp512RMqAIIxn2Jg0dIDrILP6X8wlNY5taewWSUuaQktEYnNya
iWs+92VSYvhKoAebEjFNiSXWR7obkTIQwrroLGF8ead9V9ppg0wTputhNTNKMIoT
73cc6ajyTKj0aPyVzBkAcTgbdw+IunMTo4Q6uFH1djEnGNVNkqp8PL5slj5fsZwl
Piy+q5cyNuJJt0CznwVNrt/x6DX7920uabOJP2GSO1Wdg+clmit4uzFXo+Iq5lZK
dwcM5NhNz5cyYNow0iNxP6YM9Hf0sTBwtQL32KI8iee4jutObOXgHnlwgfcwFRWJ
1w+6kxAOvJFqztmEeBr+8Bs7h8d5yNk5r7wzrtL49+SXuj9H1YxfQXXqiGgeuS6l
l9E/e0QywJWIJzDqoGT+6R4aqWo1WboK1dJKTA1DPKk1M0SlH+4qtltJ2E0Kt0Pl
QhDCIWdGzYZE9SY+4yYVtHbGef2DjXPeo/XklYD0Byf7KQKEkHs0hnhdsvDL3155
5/Ur1gFYc/ZHSsj3zrTGNtjJp0V7jBU0lwWiQTe+OT7moX6gHhdD+GfK4IykWp4s
6LRbv5idQcmYDnJEsKElWWcJ70HQTr3AJWWChhkhsLezJQ9UaCfdr3LRoGGUgNBf
dJkoKo53+pirKp1bHsB5Z0tRYARWFDALaaCUb+5Wv15GACHN+vTqJ1soB/DP69FT
151vaz9hMZk1fBw6QvAl2+BTWJsPR/ZJxWs+78Bo5bNl0JvH5hHih3dxM57hiQ1x
r5rsLVUTafGuF2yzfvceBZywHQtvAw6ME7bG/0A1KOHLWKCxRcKmJJ4MXqCrEHgG
4DGAMkgCqlJVfOVBBqNlJfgDtGHyHFwGBQ7NJ3cW48/td8vgstUy5dXb9DANlIie
9KDEIiqtTgJADAt5jQ3LkInR+MgXipqlWyXEzvZttThp5bXxIMp0zwVGyvc8c5Cq
AFutiJ/wLBmD6aA7qMGb+676nHZCxflXQczK+qzqjV3cSSQB2dV/7/5xbkjVDAQ5
zNZyE4uh4epzCH7VAk2lomaUGbrKPJMXJtS6c2CFb288HdEo0nZBYzfzi5+Ljo2q
i7SDhdR6RJGxEizHKrYIcXRB9r810RHFEFrvdSAPNSa6siLKNSHRKh2al4GqSLot
zGxzZ9YkQwEg1JFWsYEAFkPQzlERR40Mz468A4cw/16DdiAEXynZM1RO+7MRMTBe
fHpnjhxQnlwpTGnF01wang5b8+Sb+A9eXuzGaXLivGx7oo2hhxVpqs3heaYBI+uX
xzOX9izXKfEv2M6kaGGTDai7e/VKNHNQPRMBBPsMR43Qm63RBVBR99/Wbeptl8Z2
5y4IvMRXcD9zHdzRmpVw7pBRiZ/iXBRdGk6UuZyWo1qc4AZf+CGFJwsRV3njCEVu
dJScHJSXA0nOA4nOQmsYYETSEQR5aWI26TSGumcZ0dI0l4tkm3oB+TlDK18r/SAi
ZwDxr26+HrdSbmvKssE4jPQdkB+jcFaVv4pBBl99Bd96V00nKbQX80ff8c46EFek
34Hw6P3IpVQjQQamKV5NMilfX7hLqj6xAF0wWB5pQc5/Z7AMGwNeviiTXXXccLYe
7HQLXm5/8wPZFsJ1S5Sy3UEb0hseqj7Nv7ppkmCoGopVfmCJaRMhYPgHLL+CQYEQ
ocqo25V8X/oLWlXM2RUxXng+HxTDjhfw80rcSjz1AkKvw0Ms2iS+5f6fv6vRPulc
TQscuDoFT8Adjy/9H33ORyFB3joYfeE2PieRchBd4S//j2syCENEBoQZuW7NMlCU
O30/Nj9dknXHfVemDOYvtTaWlqunVQAjfeMDJkNahkoUesMTs7ma8MPfBB86x0fX
XXJF++MOetscjhXIINTquahlLFMJ5mup/hxdnGoyIyODv9ZobMQDva1vWO0u02H6
5pYdvrugNa7+7zNNy68DKPp+uTubfRwaVGRfzvRlLo3Fv2BEbLsQvBpN4zVZBGcm
yNhBSqriEIRP1yT07YgPbLIxvYBHXMxzmNhL72HLJpwaIIZtxYo7mw/koYAgMkzW
uW15hDt5JK4g6AguQQJUw6fEgwckIjxPdBfaTRz3J+PeLF1xzLOjFzR8Y3czwMqq
qJ8xLdyUKM4wnWO78bIvhedEt0K4kDN0AeVFMdQyJ/VDueyOzxl5zJMRGtpia4DP
x5yE9H13TDYvemXuucvzlBzUfMWNL9eRCG2hKUEFbFok2oq8eYKMiw7WUlZSrO5X
QL271hgcrTkNxmMtF2J5xk4TxLMW0qulus4ovQO4XwnKdnOKor2tuJziHgM49WhU
iWTuvAqRp07ZmF6U4rpVfcBYJu1rBTyJQZ6AYcldicuEKptiGUqcvcSYTij8KCEF
WOnyalg29ZzXxHlXxb1rhYKriJDUIb+/SeNM7OfTlVr5LPsTlZ9jzPI5XNZtIo+T
hwIWYr+luZT+AvxstOjzFtvYN8mEpFR+BxG9yhUx7p54kZeg85vszUSiq44C5n7V
4lWAUBYo3MSCcb9NLBH8GlbUeUB0OUiSdGna0RREtXoROsoK50+CGwBFjzcghrNn
SSmGwU7vU7UgwvNAKriUvwSiBJW4tqTQRHWIvhiiUPYRcIlvD7wXd7yvw9lT788W
5Vo/2kxwvJSOlCFr2qw9Ned24nT+kuI/6Vtzz/GbSeAoGh7oYtxGaaQU4ldQ84d1
4NKuqiYjqMHW7tEwHfBYPwo/jYvm38hVE5RuxBPodOCtkxh6e+V2Wpy8tsTsDscq
baQAg+OpkftA77rRR+Ltz1l4MYz5s5Ai1w/fokuRgIRSvIfCsctJSeU8ewUnneTO
k2Xig1nTIRmKNjwYIIe7/O5jWQGfION0zN70vW5t2LZShz54wVd0WduyXvtbdq21
yKUzNnoittQVVIv95nLf2XNdpL42syg+UUzUXhUx0jkdkXbbYVdF7uD1NCkz+O9a
etXkIxiyva6m/03Y/BrFSBfwlbWZBjxy9XPYZSipHwyBXs142R6BA+Zv4ZXRZ+HD
1IX7+jsSRYAIxX3FS/goH1Ce0svqeuuMs4cbRahgcE1gS+jyDZm802dh+PXk1cgg
Hja8A9A1IvfF+nZCT9Cm03i2B/g44Bdtoj4M6dfLfIQdTTzFSihXSh9NhjUwunZF
UjxnDb5bTJS1aA8rxibMEE52p+UyRWg3MQCzmUcrA+Cr8x5MBUj+/2z4S/kvk2G1
smEFBKtc8w5uAyBsRxq5kNl+lugvpRJxsYE2BvXVdX0YPR21Syn6eN6m5xhAuu6Q
6J9xaZcxTjUTjnLSb6BxpNBoYKcNDGcJDvQOcgXLmpL1E/AMHL0vaJOyLTyPVdku
hIpbMt6FN8xng1HbAh6TL893JuDVBhowW1Gb1O75lxbgHu3JnjxR+DAWWIiI0MY5
t19aTgXYYBkFqdtG+OaHdm+3VLzJ+GXygzNspaKVPHUl+yPY7EQTt1bLbBmPsPWP
WPbzIdIhdudT0MX+AOG8vZAOlpxy6bNZZg4nCZIQ4SMBPAqJiJTV2gboMNAqM27D
paNZumpxJI42jtGbXnDQmtsH0zlHAOyEddRTVSsoPUFR6eC8YjHcdQTQ9vMj4Tp9
4i8dpeFQ7ufw6XBeAXap+XTVsMBJtfdZgKJhENj22UwsT5jBdRO7sUKlHnbrFE+o
44QccU7I3SbP65luGtA5kkdRWUMd909B8Kz88lCX8almomBnB2jlDhn6ZQFZicb1
6GBoxK7Q2PcQ3c/YsmCDBICnJx6zj/FPz/6B3eBPcofmqgDxPvHMxs9rzHXg6imZ
Gg8P1T+hhaHeDJyVBjjfdGkePNzmkqr4L9Pv/GaMPB62lSRyoQ3oUfRKST+neeqq
knctpG8LGy8c3HmE5Rzyb6z2bLYta6OhcuElc1nQ0ZcNXT6mC+TqrTAywOKEWrAi
SL1yCfiEvmjWsAvpnJ0oN6tZyd7EEJaSwZXW6hQTdyD4dCs8n+e22i6TrNRrbLjH
RPwHuj6wx5+o0FQrKlBpGOiMGMw2Dz9FPe3xmKLFm7ltonWW1dC37qeN2AOQmAjN
69x53PVNuwntSuL6gel4/G1SYlcl9ajG1w4XEI0N8LUi/it6GLbG7WfNfUtzkgXu
ZguTEP2U8YadFRd1le9sBRKgcT/dBlvBaNkQ526PlyLhdcCL9LG652Okq5WTGDOy
oPpr91LUgh+x/jfeP6W4fpShRwRtlhXpIsEnvARS3Zq55HlRSfI0WYWcLoLJvhuh
xgvx61ewqTVKiid/Q/9f7i9BrB0hYg7ebVVYXDwcNSuHqeQgta1t6pr+0MzutbOE
F9zdCAVwNJSfHGq/hEnbZK+B8/MexMNiM9j9OvC3418juE2cyZqnFR1TwU4DQn20
a04SsNbJor9rpgBcARhSu5Eay5oSDiJH67TwOGcQvXuC6D88qCC4voDpt4imRP6N
bTEXKz/UTt8WdOuQGHPoXywaiWP5APH3ZdXrbVIpxGHlZoJN9N5D0mYtF0Zr4KY+
Z1zylQNppHEdaarS5RmUmyPVTavaWOeSmB5GqGoUn8sUhFS6JyRw2Mn25v/3fDJH
T+6VQVE9LsNkdhAGIFQYio9CvOTcDKRY18yF5UFVv7hs2HHnGnE/SRJp7VqzBJBa
SrYpSgMOw5igoYnWo9I+CsxfMxSuzoicRlGfS1duiLgenUtLLQ7wCgfylRBl5PkQ
nUr35VsdohZHgEWyDuQW4/fPdIJkobZujDDuQz/uqcpiwQEuWYmtwL/FzyeyV5BI
0FDRKqsxbglAm+QWKc3rpyZNusiz0vra6Ioe1JJmysMFVgtCn3FFvy7kzaMo226C
QviDN+DZw7ESzaYjAp6Rb+M1wtE9g29XPwLR+fxscSNgqHrOxxEx+auW22IdpVWf
NWkjiaHHErlm6g0D+gY44DPAE0a7QCqarlE3/GYewTZr6Xk+vMCkINsOI6lc58H1
YAhbPqGGGb0X6pYjs5ls8HYRVLFA7DE4+emJ7DvOC76zqcPS3nlV/+wJhgQvme46
brM6HLCVv3syp/po5WtAu4pAlehPBAYlBIfxZEHFiftNJYn5CNOJ+Rd6jqPHLBLO
s3Mw39uYUonr0FfFMFB4uPdt0+xoCvdnvYPcNUssN+G5zZCX81DeCqglVa8VJscU
T9qOXQVuQoalvb8YX1tEkZFrui3TQqDJ0hXwtUAVOk/r+05nMSlQANer2SZNbm+M
l966Y1sSpRZBAHTIT+WOAqVkb5qXVKVLjm7JRUj9AKFyr4Sj+DRt6mntBCG3itwD
KOO60Xm9vHTbAMV73LAHVk8Cz6Awmk3iUKTd200K0VFLqRtU0Q71QvUIPKrplTho
ABwGKz5OnqR8wFyjox7IbSPPPnF4Im43xSEm4/rGuVi4FkdytYH6VNPFBxnsb7C/
DxgrSJw2L0dlo/ikPBfkWXveu6ZachPVHe/YgvLhv76w39dMdCPU0hZsVz1zilC1
IZReVdavbR1pwZiXB8rVPKN+ws+Yv1bSIJg1u9CBXvAfM6IbtC3zcmvDLlkwFYDR
buzc/023KsdFAR6H2o/UyCDASLWsx8aBD8vHnyAT99ywxNUFHLieC98LhTa/Pktg
yScp33cKRfWCTPA4DVuHJHVOkm7He8yioREk4lElmlMOYb/Q1xxQIYQiuKk/jDKg
bM8fhY7BFqQAyo1aYV0ZvG2zkvXCzBrw0yv+33YbSDa+LiZItPrZ3zJqPkxyXO/p
/A4z7wynH90dZ4ARniPmERFD55WaqDJLIs4IP46TqvouwdUqoeo1BsYQUTqwGmY0
/RlsPKg3zNH+4NSHYOYqS/9KbMzA9gn3SfVbKRJFUViirK1Wj9XBD5242XIB0YxM
qJqIEjuDQB+7YtDgDU4JmKstDbSaJ6S0QghoejsfTcNWqmGxIhR/9RpbmpY1ygZd
3Cct0klfn2UkxXECQctTfjyWhE2MLE7yzdFFDh+VdkHEsf7OOiTdS8OBbJgLJope
y0VaRvko4bf/FKpx14bSO27wZPn795t9uP3uHaMmGcMPJyIZjXw931had9qiHu0F
CHMh5pYSgcHVj8lllhfA8KBtmd7YuKB0bCbdCGYorZd3a2fUbKJORYRWE6V5NgpW
WZVvT/5t2OkJr0E2DZ8mOmOZLRqau/m+xUrDkOZUraEwn31hoBYLJw0UpuDYobJg
zCxzTzteUhXhsYMeU+F8+edyg5WplSRPfSB1/igqh6ENn1SjiJVFxNX2+YBld/F6
u6RGG8fcRktcAo0Sh0vOn4faXK/+mCckskUr6k50Gg8Ni76x5kU7elEgeKDGeSNr
S0YXm5EZyqZWyH9j/iewlCP2tI7hi8NgjN35a6/1Ek8+hVjAcl60HUt8B8TcYI+b
TVNLvzkdbUV0G1PdXrFGcRrepACI6yCJoo/5RQNBWNop7OgCMNZK1ImZ9qRrYMcX
SORHMT3ZXg2lBe2b/3wmgRDHXv1IlZWRqr6DzYGTNJStztjjvSYPvMWgst+vqF7b
lmRqBFhMcC85UgrTNhaCMZtgTnp7SJN5zz1rFEioFHEuvoAXleuaFQDMB46nbMIG
zoRuqhZfQ5rBVfPRfb8aQ7baTg9XD5aOIJbnxCyJ4sApyz2sNU+kshdJH069jqFt
LvYOUuUAHkXjoABLeCfbvQge/ZZ+45awYxgM5Zu84CquBzcE7XYGWcuTtpleYx9G
wkxo/hhOp3LGvgtfvjn5I5AGggASUH2gbS5XBxT7Cjvn80Rpswj37dK04gYrlSo5
uHOi/FhTuThvGlpR8c2DUGn05owMPYSKuM/VToQt5uMMA59QYmMnw+BtC0pSk2Mq
y8UkU+76VO2GNvnQp6CVHVcEGrvfVKFN6G/SttolPzKKXGk0etCnIa37kk0SVuj4
lWWOv6lZTaQ+9xXXy1Cr8EO5rP5A1JF/OfzpQKwrNzVlBIG8vKWon3L/2+QwXAFN
gkocNkQ8vXsqmXzlNqDyjBJ89IjdJD8/Q08MHNk+x5graDGHepqRPvzbXV5YBXMF
VPVwCDlqEfzSgaFj6KhYZuZKMZDpkkixRn3W+pjiZYzKvBQcXhNpddmD3UN2CFv2
bgQ5yE1/XBgv7EagkxjbVsSsjvHLxvdCKCPOOy/KRUeTnr1bz0bXD6qB0Jp7URnv
qrbO7CbZ4B5D1GFlbQ42FeP4STbEAMR0R5nLx4TC8t9SG6kXtsBE8iP9fZzJVSFl
ZX4krZKbMVBfsXlBvE0FK98R51V6AAVjV1pGi0ST699/rmTk+3jCsFNRVstOwybe
4GMAouYru+Hpzdn4bZe69icDDieVlE+s4wx2v3xtA1+7q2dXkYWzcF2cTzwIpcQ0
M+maG81fZEPnYzpdkeBq1JuH4cmGN02gqJX9ou2r+mLIngXkjgVEsuJkKjohFiAb
paMJFiG2FM3Zk0xh4h/ocaMOHOMk7o+mAwTmaMxJneZHJWCQdVAyjwqxoCn++xat
wEbHzp6FGezWZCJzx6keGGUWvv7t7LBbo+bO25Ms5tD0Ov2eUIekl7Zob23EtrZe
o50ws7gfZb/jgWM2/95jz9tKRpMQzmu0AT1WhcvGQR2snd5JGAb0K/B2WIjoGsTN
7gxZCNiBOLlJdTa9ZpgY7zy9hKLU7jS4p4NJZvhjNglFTV/OuiwLymYMa8TTlIVm
HHzOgpkyqx/pbGHjWf7FMDMAQnZvrCHtVxdree1JOcNhnqSIVwJylsbwhIixJokd
PWpE5BtdJ3uHxl41KYGrbVbaoq3BdQQB8JKhwtjqJ6UioL8TxwETsNu2X/uo5YD8
vC3Gkdoz8ZArowkfnrQ9Lax5pf1TSA0SQZ4N+cmUXXelN4NlplWbX/c1DPaP7wkJ
odrs7JCSWUYVRX28elGN+/Zwvvvv1kKpNnyQZiOvvfbO631xdlVTJWvyz9hjJ52y
BPHO6JTBnoZoJZ1UKKQ6wgYlK2D2SAaOotmwklaQd5VHH96cIsZ15GV3Gmw0QRse
UdTd5H72yaHSl+CWfd64rC23Ac36IPpZRN/vt+UhiCrEj7YBAK9LXssqST7jngbd
FQDOR1USMkdOIvoeF0awatxWUn4994JYCySx4mAtmh3pXvBC85wkJQyI5wEzR6fS
AXGaHS92fTYmG7YtnR+dzAXW0weJ2YKzJg9AbsROMQ5QX9fg1164LcjGern/GYKx
lRTigMa/tkaRN+7C3EXUGcVcCGzo8TD80oAI8md5/W2g6XpePRbJerV2LUEC96Tv
23mcrSXR3uS3hI1v2XTPHpUhH1Dcrs8muZlPyc+fLibVBM+H3UkpiXDXV3AdC5HU
J8Ks1fVjM2Yy+DQyk5mMg3nBriWa1ZbVIDqjPXrS6esZ8AngpALy7WXqmcUgB/yQ
sQnZXeJoPPocDliO39u3HOj6ZcFwIGUHpGsc34GmztR81H9vgM02nVfIZI1kxA4D
3zH8wAEB7bgbw8tpz4fapYc2G3/FNeEYoDJVBzJ0DOUKeTWv78NT5f831oGBpktV
cMJtA5y8os4JgjU+IsVbg5/O+R6Cx/hRE3775idr6pXYES4Zafsk9o3FlmoxxhJd
mJjLmzWfvkaYPCNM/i95O8ELVHlVlGIR7dl+xBGLbJxSrbKB+PQ23WZMD7yiMcxH
qSAzM7DSrEIaQXATTdor8c4duDn/RHadQzvEAn++9Hn1Zd2ONpK8l0kqhuQMpS8B
O/6289Q/0w4TuAle+SmjqWvV9mdKxvR5oMJ07iD9CavzOHJsKzi2OkFnit4oQYOZ
189rP+0ldwa0m3WkoxH5jvL9AWQPhGQ2w9B3bzvMqU01DWP9b9ZUaHcAQzU5PaWf
VKoCCF40INE9VIHXoj2H21qSRAESfLnGEv50A033oYjzDdWXtTCjSdwawc+W05my
p8QvL/8u7FWLa2gbHD2gs3RdCjp+ZrE5D8KSfQsHs4dvY4Bx+rws0bLHMNHvlzI9
VaZ2mHWFwdu2sH5zXqU5bri1HKWaHpHaTgP8N+zTWOOO1qS+k3snnwMn7k/1CKOd
Q/dsewMsn+tBuej74D96bD0QfZQbAbcGFUfpuAdXcILhONjHBgKNXZdbIQn4XAp5
rpKHVpdZnyTRfIuHWhh1KBWyfo8hJY428KILQX2zqBVfUE5WImeXnsS9i4HlYAbY
D8YqkzeMsoe92906Ztf37HlMvsWIcCAKwu67C7L0pLahZZleAlwCVo7t+D61tJ3H
Hvss0taKFtMt3cCxY4o4jk8dJk7GFMBbzQHv3jrVi9JwXOjF8w4v1ROC3fflG8e3
6VRDNH2DcsVkkYlJLImVGs4B78J/xf8TWh9a7J2+w2oB//LnSfjE6sYlgh8pLwn0
RrE2RPfuKeuf8aSETk9BTK7VnGwmKsgdK44r6dBm1iyACZWWHttRxAlG1fSOMACT
SH3FNZkh3Bh6VI58jb9hjHmH6j+3Nz6G0u1jOGs6wZKUW3staRtjYOeDzIAqT2qg
bDfyatan/V6MClPxLpZgqgmKEsaEOFhnRwV57+KyPYWYlwZc4007byTgrWZWIRoX
+x75rK0asinj0sk3uKrT3k8PZuf1F5Xq20Lh9yl8ZhT6KOvV++QhN5awqOHaEZYj
8FQrA/bSPaVB1CDvSITtWDwA0jT8MTNTfK1gQjpxkLpGAeG+5B2alL3X4en52DFr
Ux/BSqfLhUCj1HADMe/lqERtDBGGg2G1ip+n3nkeHh5+hf0OqIP/Q3k3122Z4d4q
t6ut5Fsm7opw1iwzBFOQijZPZGybel03UO6w95aYRDerX5/83w0lXku15TGYpQL3
HQjldzNUfA8+lGrg+0f7U8Cd/LVUbQMmugn3kOJjSAdKHlav2QGThoY5J1pgJ0Gj
/0+NkzVJaitXTrgm7Xv2feL/3O7DdKwsILSSNJXlNrfH7t6DjaookFGiwviXLKzA
2VXbO3P+Yj16ZalM6Labi4I1ho0/Z4IT427SORGHU+4INlamAZkIdA5BQhwnBdGP
LFzQnTBzCem3vJ6XACmenFm4SNQyO3dprv+oo+2WCoA3PfFwRkEAzuJ7MR5sjHp1
91gLiZzvt8d0gWOZBW/SNdsfU/1stKzWSzOXsVxkFgexnCZslTitlVVq+NI3wg/Z
JiEKLLxj6uY31f2i0ijqMN8UD3VHXYkF2+1F5i4PYDKhDqecRsPViVGFz/ZAVPkL
qqT9TryOyFoUDSVastSU3M1wR3Ats2WzL7VJeXQXhCXYcpViQ/O1NKen0BHiCykY
j13vtK9YC2ub4jeqsLuzlWFeO7mYCpwYFAsTv7FjgC60MIJulfMh+4dK8gRXmR2/
ZoRn5k2qU5nNEdu/VY+OulN34BfEFC7GZIjazEDuGF4l8cIhwEdXmUxF84uLE/pC
A4pquWbj1+APZr8KEHsjE4bBmmbKIHoKvH4oW9I8OBLxbO+4b2FtPjk8GwAxTJhK
SOeR00PVLUVddjLOTtCOEzcM7TAmJj0GDYQf3GLr8b4P/97o1isJPTBOQ7Z23AK4
NeI/lmy0K+jPNncB+uwZOlwqb9Jo47aNIETXnOKB4arMQ7qktIY3bKm97onTuCIt
QRdx4p7T/uQ0T9B7tY43/OP8jIH1lenISmBMhDdYe4RkKi+PpHxPi6Belj9n4iSi
Q2gRQwtJYl71L0KSTJnI9yTe3l/PFKiHTSHj6iIbVgXNd2BcM4xImWGZUkx5pKUr
8Fh5Weit++cd3smSNSmSZ3eRUb7OgEkPuq2VPEx5uMk3w2gtkoWK79AERv+AYRYb
bAMsQvEz4iy8694eGoAZc/wksIqyNjyYQaD/IzcLeR9UBp7EzC69Hic8RU7O+Dok
h//zXK4Zyvf0yqvAEIX8Wye7ylhl1QrLdfqhGEiwk1QpnSmA3LeG6FcAeyLy2m4K
/FLEsEZdiDcIIojNWi8FP93XUC+dhdJmVgLxCiR7Ki1LF5RvDQ5AyVbic/JS0gPR
bujGq4wo7D65y6TjgtT6BfM+oGmoiz/mvwba4ojiAqcK3mrbUbKIz5YNzJToM2zO
Q20y6bX+bOBeqv7AH33pezH0e/zYZN4bq3p6rvK/i/f4F4rgQUwbLAYl56gUzDsN
cxz95/IF1h6LHcWhSQs/DaCRhdi064f3E/imqHFyCPWX1ejSDhkONP3A7YQBJmh3
LGYXx3IcgeLiJd8FZ7TKtRb2KfANp5Zsa41+JsZFM49MrTS2ycJzJIeAr2fGPR6n
aqQ1nkkqJOq4fJ1RM5ZYMYLS6z+YcEcsHB2LWrRUzHYcO+3P4P6wewkD29DW8egK
2N1iOgwekNHxDYS4eA8Zdw4jevk7ICnIa9Hm0dadZn4prF8k8JiKfsq9PAoHAFW9
BVKg4V3/AR9GQr1GkWwO7e3sW/BUEFb8NFoqB1sGD0ZUIb8yJ6wlsRUuwv9A1ZZP
YSFjpLSFDLPMKWq6gCyhDw9SaGluK0oEo214UkVPBxw4raOHW4yFP9jDcgtan8PJ
sm3Wh9IX/eU8D/casExchNBO/63stySWKvHcd/u459v3boMoV2grCTxeeQAsOVD4
5ZVi30O1h/eBgsxAomsk3qWO8hcqgwuIogfmlJ47QiMvjjDV1RJadlOQfPZx6Kl1
XkdwZ2dt60uBKMLWgNdA549ABERF56ZHOd90Ua8MbZiC66cEqccinkfpTYu50RsC
U26ARVOB13jJnRfitg6xJpbW09Skl4ZIGIDDOFK/wYavMhYceTBSu3p+biaiqKSx
PI0d/BUwjSNA8yIV1RINSbvRTx3ZhowwmKPl/UGLdm1wVU7rKy8erdHHZP5DVIqI
ltGPF/uoEkYoyPxZtiFLZS7Ehztw0+lPgfK3ZT9v2F64xDCKoqJfpeVCNiMspmA6
LVAgSlJq2REKsH4MKmygca+2Ee8H6IFhFyD64FybGOtJo+XGJEjYWSd+5Jgi2K5H
PzJaxfaVrkvFnp4UNpbRFz0QuIvUP8Gfp0mFO1ZJCw6QlQigxLAybW7Yuw/XtyPc
6MIu9iPnCo0yOPTThAGm/iGqi3naIlTN/SAIlR2fQPWUQBqirBieuEA7HhzATSXj
4p48kNzG0riWWyc6xQJ9NCLrDUlSKVIWUXCDnB+yRtSCmHOyY0/X/pQGg1J5Nzzg
69u03wiBKpEzAF5EUUag8zmRNin2cw8nNWCcW7/qd7mSlthuN0TTCA3/S9vXSFN0
8tNrqiejZpKky2eTzy/VMy8ed8S97gJfvnOGCDOnnDiReQLv0G8hN+HweOGaEkh8
O1ZMCfUtAW9MrcO2vzJJcUW2+QvV+ao6wfyr0hD0EizSjrdvbrGtH8YxSt6tmVmd
Eu77pgrFP7O8EBYHNtDsCOi6QO5TrqqbRyesBErpsjtVmQgK1C4QbpQjnkwXepCS
RxoMC2yhrOtLFT3z9U3AONwN+6iW9qKrldK3+agixpEDOmy3kUxgDP1ZT6yBCnlQ
NuFIBCF+wbHQ63RRBJ+HTUwiP3ua15d30S4OdDtA2Xt/yxOLxkMkPSzrtq0ZEc2y
CScCepk3kiCkN3y88ApQOCo4CFzNzlHGi3UsigHwhuNBHELRGfnMUkk1Ul1ApSvg
NMAWsSbdFJbf5cSkA/Hlt79NvqsBsoRYujki9GGW5Hoj1HsNamDBGfN43bSrozvr
jZSbNZ+MOC5r3rYt1W0wz4Q38+roYk+yGcW4U75xt3iRqOYvRXyY20B3AXtwxkPG
YeBZ26oDo7C24Ex8UnX4LeAqEb7mvtZOHHVDFxBWvgHlXFUwAy+IKrE645++RT/1
e1AZCOGMmA5HGqWqr3deN/Hy1n5YraVzkleOXer4shpjC9lEb8K0vcfFneoYwkmZ
Cp/aYPZXutD61Lb2/fkoeCRWVXisPe2rN9CbIyWdmBHABOTpxA24joGeXdJGV8Um
dSQlO4ZyscQNLBS76rMkhQFdGTf3lc06teM0QNFU0zJdzYAy/7eW/UTXJoyFTMqm
MSl9JZkuUSLaPZjPjgCK1IpqKA2caKRwOvdDpf9RILeXkv199ynfj8uL4lLOmYry
wwqEA4PMK3goyR8GXVqWRpQInrwlMlwuW3rBzgb9xi6EpG/58UrG5LxczHS9ee6U
8dbu58IazzmgAVTn64ag9pN/A92cViJLh+dofG03q68rNIbI4ZXHTCMlvVfKhnw6
HbPNOX1n5hSF1eAy3faQ4t61KwNqBPa9beuYc9atB7Ab3YW7KuGtZSy/Hzz+Ot74
Sr31Q5U+5i+efqRA6O62ZFXheBbCBYgmeKlVbiWOlbdyKhkhiLAIP9spxOYfQixG
fnySPfHQgSYHoIHjS8spqx61AYpCBeLpgKR4o9lrOn3dVc/JnybG1Z9YfwQAwhAa
M+eWc3a+Jk19VO5sxNQikS7v7HpZFsEXF76ZLYLmhkZoX+4MVSwCoUFnW/v1j/l7
XmGpckNVNTUIEbuS3T+k1aW+qgpKZfBDLQpf7UG03GVFhweWu943E5e2TWNTs/9i
BV2E7TW5ot6m0MbloLcoDJYY0msNusTx5CZXAVdCKjJzYAwt4qo2yJ2oI6LyNhu4
ePum29v19GT4/Mep2qxomdUYyhNXme2svrARxJoUatJjxKfx7UzGPhGcVXfzvCga
/m8S8HCpNnSw/MzfJhRv7WlTF8faG+gZYLYPdRtz4F8hM30DKSY2Fm2KIQva+F9c
/RMD9eKkkSMxUBkemix09LIDvdHbJO7tiqgqNUkK3hjPXxnlwYZ4AFO8w+y5evbx
mY4h2/SWLixrXrE8FDaLqHsU83nOKwFxtdHjd+UddQsMBPKvqItScw+GY8fIEUaP
xEGRFszJ0YnI7grTuaFV3NrfT8isKwVWpMEPa6xI1U1SB3MOFasT3qEGHgQlDlo/
RsVSU1gbMhOUoUuYQzX/XHrOHE2akbiGWpPbGOwjiAsJVEaZdh26WsbGtSQLIHvp
LPpWSulBqASCAHdLF8tw1JTCEZ4em54w7A6hhM78gJIojW7+s+bY8iMfzqu050Vc
dlrZ/bxQr7SDB6Lm2HfmjL1zX0OZd1DYFYZfKfqpS/yJvN1kFo6hrA8mHBGANqWY
uGmVFwgyjeOb82xkiDfNsRTp/PFvih/83U8kXcAHCYUW5WVgvvbsv4Rapzy0L1pQ
ZFhOGbJSQn/2alcDilvzLKoy19Uf8sNCj2OhFD1eMLmUGxkkXRYD7wi7yPuBjQTu
+xUXCTatLz/ZQ3CyJQrr3aBWiarqIGjasa0ZPXM60bMYK8fwD0kq8MlD6oLAg6uB
dvTm6eqKXhsMURBqSuHcSk3Kfhej6HRjZzxnuj2gCZf2C70pMiQIJFTpLWqjvO6g
Vk9dRZipX0wlTfvIv/oZt+b4meYDMUIPwxu/vhw4+9PZeJhi2pDABUWPAEMVRl+a
WsAPifCwuni5HtV2oYLkxxDBC4N1SkeNRJeFhaxT8LrSEfKgxj19CZGIpT4RWZ8J
+T3kGAUmGeee5fa8RwTEzxiVGpaifk7nAFWdDMIRJ1tVvb02aBz1aq6ZsgtlwMP0
JjHAZRvpX7GkbNAPiojFcE5BkU+XjyPoz778p6r0C19DSj4fX2jzBhakYvEeYqSO
uepPzgtL+H1fJU0IOwU+eVxC/XqGq7rIGPNwhOaS/zpEA8RW07w7wRBERpbMj7cr
1hPRFanjJA0tK9Y3p1GQCkszgMX0sIh/X20uNp9IJMLP5LRWZ7Aea9JENIaQmB4A
3STFgNMjyqiQSpr0rv3i4ydbTGOyhfDTmuQp7HbEUH1M3/mapud3NqQrhjNshz0y
t3B1d43cogoA6UtpccDHFsKM/mpqDbKa+KdYe6fN9cesdP9pSROulgDOxmHOcbcV
GFd1dbnXhkDYEf/BMa8LWV/+6AVllrrx9gYqLzOQdmXjgyTOpBMZrkWOccFQTSXJ
o2CU0WwrT95yQnZWMKGO7eMi9ZtwB746KVeYY2Tspmx5YSfTkxrQP27gKDi+uHBA
aQNgagouRx4hToUv9JqKCPH0FFr78lMiu8PCHD7iafypzRazegNyX3UggDoIdwLi
GpxHBRBFPDnv33+o8HU3/PaxNQSChTDWfvVj37cylumajCtayI+Ic8SSuwd0FQaQ
o0RMIN18P4hWk3RxMXcXB9y2ygJV7R3wslSAxr6FuKgoRsMMLp4nO+K9Ey6lDQpk
7KXVejacx4tJ2gXcFvlfBqj057My7iPyExMAj8//c4GV3cJt3Vl+sUvzDZ6NmcL8
z8i0iUEsBSovHM77N/pke60UOLkEX40KVBmPFKLgo+2mb/P0gb4mSE+QqTkpXxl2
fj9BwkxUnDIbcRLXnxOl17/IzBss4liGfVxFxGRy5ih79ZeKwTKyqmilwAt37Z07
IJUGNXCv9I2y0UfV1eMc8jQ2TcQ6GDZmk0MjeIb4w0OBeR0+K5KUb8vU/5KVNB4M
LrDU1grbD7XJhegvxfqAPjMFwBa6biVLbSNItRzfxPtCYXgmP0Ca9ByDpnm1gpXi
5nX2BiVNS9K/qgyIiiT/nlBQAEmDQvZ2L1Kvsq88wHC14iCBUIRGdLTZp4tLC13f
k1Shg16BVnyw/f9DV04zkPVNG7HsTjkXOCq3cAlDaPApsobK3AKRiZm9OSpwqoFL
lezi+hzZ3YEZdqiI0HtavwAuHGJaS35oqWtfh6+SFy2u+IKxDn4aKYCdd9ph+FiT
GPC2dEUO4CvBsIeJaF66bLmQajo97F4xBmG7jDXndz5tFBDRPiOPKZ2p9vW9Kj5O
2YwzFNhabm2J+eK7arGJZmAUE4VlMqSTXroJzu1/TUxL2Qvuz4SeseoO6vcZVAPX
nMDbbNxtKwFHV7juC8SIGGEZMsSqXPsCpSHQeEej+RMoDXQY5+T8xe9W1OMsVGiA
qw5wSu6DDpj1FnP8lwVa/uUF/b9kNh2pwIqU909bOO24fo9x6WVbRApTfL7MNDxy
Wpnpc+DI7J8gr2ilmuF3Tndqm7qPT+Wxx1ububQu2EpV7zTvWG9jG3UF92jYCqiO
IOCEJt/2S2Xw2RMvRqcIpwDrTInWdAynKUlnvJAEsMOlMslTU3WHlevdCHiFQ1Tf
xRAlvTSNi4pcIm1+Xi7vXSmMeOY4MTW1lVO2QeQsKeHln2CnlLYsyFsUe4pNwIk0
j9gTSmFWl7+YhJlavDfyZMbjV1FTpSAg2M201tc+AaBHLfjKgWfypTkaDYVH1U0w
x+zAl/DXVt6l8Yuk/qd77KcBrA6BnBRMm0gMQENvSnhpIps3RpoTSnKTXXN8GqMq
K2zT23oQw3tfqiUMtgvwhwRU7uEaip+PR+GBY2aDaoThnWoDuFEgRpRvZENJ2+4A
hlXzgsQN0kO9zBRGVQFEdUg1rTOfc/Cp7NH63FDi6TQTWQiXEsmE/dH8j+kRUVoh
RMZbNVN6Khmy/XByNPdzVQ25WOPiSqeuQUL/D6nFdVLH8AkI3saw7Hqa/j6LmG4R
EVlN7q1DUhwpJZnfL+Q59VC0ALalxBTqlKDPKauQRCCiAzQPpScxx8lF+hnGNXNY
JqLWqP59ifN3bcw+fdNEmBVuEuYeBZPwFJs89CeFt9RJPmQ95VxgTtYinQ0//QgH
Zk0bFij88dpjcXr5yVucjQ+v1IfVnfyzbH9TYAbQENpdtzW/odnsmcZBpAdELvTi
eQQQe/TzlgNsW5QIGT7gnx9sDBRVHZqYs7kkqL5wbk66OBTlulR+awicMWoj5t+S
HVLb5rwNVL5mJlDla22NO8zDuABRA08NftWoS8nBIliorJ1bQMO9v18fc66pgE7e
qNkAeguO8yPrcyn0mY3v1QQ3Lzo9J0yewwthYwsD89E+/JSfgstM931bEFciXBMV
qoBk0436j2EpD/mD/3J7Zsc4JqWvyakgq+CgylGqBs0tlzsd/MBQ5HCj5HTuBvTw
YttPDE4VS7ii2GERjUhCxPiISUzZ/jFF3/2yiZBl1/sW8brrWF4HdCd46h7dPH/H
yxmoebV6NxmMjnH85LELb1ysNaMNDBExPW2TZDgjJQo0RXYyUYN3YRHdtTCOMlbu
ZIRUPU5zvjp0/tXpe7cgVPvnBb6WDztUvzVTTeRPnZFAqBNazq+650dKRQGaUtOA
EeeiMjIR+g19SXiuxZgGRz1nF4i7n7DoPrzrqQnh++i0LYJ9olgO7c7pMDANPqgO
MYK7Kek6ojTlpKWYQ5UEXOwsZmTdox9VuIDRfe66JpUNLf8i1vGwMeKbyfd8FU9f
OBpNnEWM8YaoZFeM4t9CKmjQQS/tmFXiYBF4G1TVeMvSVX9ej5mm4DIOMa67Dv4a
G+J6wYKVYD3E7tH8hP3b/NXqSMiNdTniqTGY3kiym2G9Wgrcz9oNoFt466DEA7cg
NQ4I2t9B5wIrLhK9Zglrdnlv9EFDufJITU6WmDYBDhdT3g6SX1Z94P3lCLWYcPcC
oV+/VmclyB8bj2xe9jUZc6LuPq5bZArf0x+EVIRstHiKXWbwY7GS30H63Jx2QyzD
CgiKEk4mbUapt6oOv59fratl91sOCMcDrwqrWPv4s5vTMwQHXGgIiGFw11OcWdcj
VazD9C086qsNJReuAf8My3Iw7nR3sn/1ePsX4Pm6Fz8Eo01vUxDkKpVboRdk1wfq
lRTp9zdWDgb5/M1Rno01xKI+j4m/zT/Q8rfyHi6e5l3RBfCzQG6Ic0iHjCoHGBOL
LxoZbNokLqtm5LulPiNuDi7Z4IRs00yzLsIb4Y2ohjZoO8Ic3lCNWKGYzdgh9BhQ
2+JbRR8NC4n4EC9UKp3iJ2XOYcLKj9EMeCSlBTi/zDmgGnHswKDWNukV2WN20GSu
DdtEoZChxd6gviBGbu4YTVUtAkEbhpMskJvcD36dH3Fk4iA2P8n1oRiVKOWyJYvI
aJlWMgc/P9PqAMACMfuH9SrwSlIfgUVhrkG/LLAnvVXhplDGPJLkyQrAb893Q+od
RVh1OTwWR03X5MMp1RjHuyyaM4OjQXJMKuxyATZ443EAbEwxLBWrLI6l4KWRdZkZ
gN8ZfcvHnuhhH1kPvWqavxtPCtgjK8G6CBeB9meBA06s8Vy+8ebKEM+GMdiCLlsi
26dq0FQcQrhRlQUK0gOKnozkPGE83AirQaAww6Lh0F5f3gXJVs71YhjgUB9eHHvv
G+3qRyhlPSpYf0+bDrXU/EXY5Q+czGGcdbL+JehpKivkhrcQPDVIBdgHmXBgipn3
8fJh1v+DxNf8PRBb6OfBc734vwW5URREs+wJE5/lnHqvgrXNRNrakDTNBjwqFJZa
va2s2eIvJzl+4D5gjAcDIH6yqScz07/yI3VAfra2psCfLmCC/mO8Q610PCyIiN/X
CADL1M9TdyIGXuOSY6EOxGubDDR+kOblq4GWItj4nuGBoZdSY4nLMeIah+XL0/YN
GZfbSWPFYe3pqCRB2b3R8Q76PtS34KzpDRKrVqTvN33ryCy3ok557Q+OdIEt16rF
9z90zGWJEswAKSj/FDHi3cYI/0v7K7D/qjGEy9hHtJOBGF/+2YvY2/kOrx4Xk2Zq
qXERHABmxi0vPArKeyM/aXAQbE0zVyssMVktPuG/tbG8WGdVkjEyVat3qmFpGJZn
3GGdZl/qsOncktWOY6XWIfsuupfBJHdanGqaOH1/FtRiHtYCY6PDpAA1nde2XhCx
vDpkHNIX76jr3ZNva21CeTmmfpbNIgN7KkxVsTTmzkDE+V1qP4Ve59NRpW32HHd7
JK6sVBTR6Z1sbgcMywbfrNm8c/sUyXTCfqiQZefKDyCmNlSRfdkc4Y0Xs9Lg76Wu
3xHxdGHPqX4HfqSP9uVDnA7SHRKq77PF08uv4wdYK8EuffNFl/iO4Ndc3Bw/9EoL
H2198GSXQpf62XeIUxa2A+kW6ZynS4TJWO+5jMjyt+pKLAFCPRKcD2coAC40SHOU
4qZmYTPCH8is043BgP/WJFsXV2biecLUNGjZ9869QdOZ570lZO2TQWwU11AWUMkA
J4/kb1JFRtWCrMVL0SHFmDIeyHY9NUHVBAfiifOteaGLzPbq5dzjl+uwFz3WmoQZ
NUJB2103+N8BmaW6+yHN8eweHArdgoG7uLvSyisq+Vw0Nz70SHNua5ucX/Y4gEHF
rBgrNHAxLuZjKgg1bk0R0exWITQuYwMp2RstM6OYhAaQL/pckdckYvmzowakumSx
6tFuU5JH9mbm/qniOueK3cFOea00FoPe/WSiLMKZS6IlOdxmBKJvq+Nq1dkqZIwF
nylbGHPFal2lWPGexsxX8ksDQZpPANxFGK8LU+DZk6lSpAn1ijLrO/i2FxvgDsND
ib4Uqz4bA2QEgfe8+h7XYc0grGrUU+1fLJQ1hS8N3gDWk8hzFwtSdnlzEikNa0JZ
wwEM3zmEFtGH99ck9P4M0CoAPNpStdHYVuZLttiKOikxSQG9tb2ZXy8H555VW3gc
Ceeq4CJSvw+1BYX6oSFldIDrSUTkAn0eKlOuyRPbfQtOQaKjl0+EjcQbwvkzp+2v
1mc6Ov98BgDF3lpJuqUpyf0OLicwPOPvir6aT6nxpzO0A862HpkEzcyKQ99pEfrh
NhEAG7vH1vzuPu7hWEbIRGwXC7D/q75cJbEx8LdF8WuFkeyu+MBao7jNX3YXu7rX
9C0MttXMyrfyW+MSrSl6nIWdgnUpfZeqzUxj6oBNULVIHMFM04AbIXs0JxVlPJBu
41Tj6f0YAVBjJHA9zs+26jk9obvTz9aJ+ZOUT4BW5l+N+3mnmxARs6vKxNEtknX9
b20jR8dxzF+Q70goFhOpa6gtfNhB0mMofE6/gto976IfIjyvUKTlNme/HFbI+OWw
kzqp0/6kiV/iZZiPcxe8nbvaodeHXUaHyFjfefQH+pV+fnHbJ1Cy8vUxiGS8W+Vd
xt6FnDXfsromEWiAkhaEfBg/VCB/i/ZGxJHcaEmVEOEzQIUp8g1eJne6A/5Oe3XF
IvB/yKF/mCdRsYrEq2wpNfvZX37S9ZNAfbQLSzexEiiU25HTf42FXNvN9QRsknR+
NkYnN+IPjjCjDMKmFItfENlmOLYsMcAgEvR9I88iKoVjklwG8iLEvS0iuWrjc4xB
jPbKdzNR7rSkJblvMVpasW2asZIDJl6YHuSItw4hjH9QZbITYS5Gr2YlMFCfMUXe
QBpLW0E4Eh5WPBwW4uXzcPR01f/iQIkTBi2VNnfa1oTArqe03/U/Emli+BIEWAYg
aQweF8TDafC8xk3xL7p7gm6T0LuGwFD+1t1/+d3IvcGpEGLX1qQ1QJhCCcsrFzLx
YUgdPEo1TV/AGrglfI5wOeE2AraqYNyxreoc1h5Y3cuvqVJLJTTZxQrgj+3pMifR
xgfTpPZRkdHz8whxhXbYAR+CWFIZ2iT9M68ANwiyf644di1p4FdI7ngliGYfv/Xn
WGKJW7yMHKQX+Y/mytgOdI2Gx6K8ZHGxTkIi/R5Fg0TvRsySLjxo3mAEOcKNq9Mz
8wv7lq1CwW7Z2EzwKux1VwibXuSxqllDft8NOOR33zdosZZEmXDPQJN8ntzMt7zU
+rqXY3z6712yePJ8SG40Jn87z91XfaKzwei+NsEXEqM99oVf26hVbkc+XRMZo1ur
CB+UkqENv7LKYmy7vuKY2hMcTv8N874FWmVvITBALkqG89+/aajMLU8q6Xn9DIOv
r4gC7/uSlxaHFEmLV2ZSdBB5mnWVVy/SjwmdBCSaijlN8cC58ZjQfUuXDMJxVpsq
pE5oZU6j2u9rbfFEzGtOHL3mIXhddtG016pGiHlqBc+KTM81alT6VNA2gakREo7C
G0NDttmrvhP35XMVq2sA7hnNUKaOSis9ykEItjloSUOkwR+bicgSz7j93CgqGu0z
qRDxdOQiMZmzPs3Fiw3AaB8wF+3gIKUYoHLnmggOokjxTDo7biGkdspyiZ0y2jL4
kzQ0OXN0u71KJclJlW/axPyTFJ+00kczx7sVa4+GwsoL6Cm+Mzscp9W6RddT1Zvt
CmTu8yKTrArcANAl7DMuUSUE5OagiCJzSHyHvq40/OxSapfI1LBMmv/I6Zv6P2/K
vniKLE7ieiETvTcYFbGws2Dbg7sEFOUpbDS0mDY+swmBM7a76dMgGhH/zk4jjmAa
bbJhmNh8h4Mtol2xtm/7Gd5COeyeRy1QWHyd7afiXc7YbW62lzqTi0i+9mGc3zd4
0QpinW4Ai1+k77myLrJwUAwBskffSgnM+hfgbuDa1nhrIpmBzx2vY/uc/guhXt7P
IgaK/aWbi8WT/vbErZITcOS0NJc+e6XCmEwdjVE+mlutoWBm411g1n3L6QuWAg6R
VKYaDlcqHp8j/6gQ6M4wbnfNDQCjGCyzf5MBZoou1pzPewQ6+xSQblJwefD7UZe1
sp8MKaJ55b0ayf3wtpfNqGY2m1+Ur+HuzgRABgR42xxnaArQXsRdL/r6AxfoTjr3
RZEIbqaP5IND7xZrTfJg2r6SFE+TftvMp30XCCAfLcfPPdAiFQdyXrAh+PK0GiF6
FvJNWY0wP5o/TAgAqW6bFQkpzan8iItC2nBribe5iEHYeysmrA+eshMCeIIARAdN
ZlcakEZFXY2bJJld2G11G51BJwRICfDcjNup9i2xHgjEA27nQVI0xNVYS0YoEKCw
pEP43jRrIFkrCpfAp8FqX/vl3laKIX5HAYE7eGxme7iu1viPyfJqHC+0MgCM/0Z/
sejNhzoDmzTe6vkt7Hq+mgT35PzH4o+J16+UGgsk8XbblMaHGl6iBfCg0zxiIYoc
b9HpSH7BG4++UYNz/qqBbcw6e5sOaDr78ebgW7lbkK32icsmxeEiHU7J+ausnTGO
EocvNfZPk936PG7XQcblVTZ0UkMdxieDxo3aZm5sUcsc9oN3YLWxjJoZaxoVGw8k
cY3aSscH488o/2Xc2EkAXpW93KjapnMw/tMhfozyO3H9JKAr4Is3DyKIUJdqB6Cj
7TWSeoSWgHtGSOWMVQ1crDzr2HVyQcJJhnUj4zAG41jMC7CXmMM2DokbdteSBniH
IlkklpVpyfYyH0L8uLAf85BRicgapxilbSQcU2g5A4WrC0SejGPh03NN2/94Pn+1
GQWzGCG8lwPpOszFkNMC5JpbO7kEP2oBFXuMkv4O6ZQrryF0fHH5nFdrWN5nNI3h
/TzcTCWM6HTCKZ9aLkULMXSE0pUVoPM+sf5KXBouejOXOA6emAtqZWEg8x1HvGLg
OvHdB5xUgOJaSNYHN9lCFwYrpwyATDHZTW3vvESpk7Ce+ZtiL3qIyvaKy7qZtbv9
oLVMt68lo4UGJJrU8XlTf7vziZtDaBtUgPsc9i89jIx1ag7NdfOuhWIJV5QOT4Rq
slsqvfK/biiorblbPyvUZpIx+OfjnkWVX63noMz+obuRo4bbekK1SUTgkhrdcGV1
wmHeIi3vgAjBe+Vucj6SW9Rv4ushcinWA9hLI40vI3JtlMYYoLv53fXIW7so2YCR
XCkeKhEuIhXJ76uXkOcHM81em7aX+bRiivqFAHhi3ayRvFpA+JFTaT/l5PqWNH4k
m8UxAoeVmuRh+0G50ux1ZFCn6PWw2kt25r+s7SwvzcnqBqcNyZ+Mh0Fs2gmN9O2x
S+5I0FepSmoDk3cAc3XA0e5YOvK3IOleJEt6oesW8L3VJPY74p5l08E6xIKdQgfQ
N/MIyzG7ahK7t6Dh1prLfNDk/xCJGLeoT5QBdIWp9m9PU7u7Rxs2OdiHLyVYYhfx
3L89IcoKh542hFhC/6AlvnyCXcq2sRO0GfoRhsMlJ3SQu9Txp6lKlVbtmmswFPSe
k9opNjQGYeJOvw0/+ntYYnicmg7LdSFLoqNKldUuigzAEO3nsIqHVTC5l/g8KP9a
r0Q5aPgrOPAGa1F/7hdW7xac0MN8162okgdBgokai4mYoGTDtLx2LT4YTvb2U3eo
JILSapLLdMJrevPhuVSurMM/TrU3EHTysYdygPdZuPog9+a7AyBEqaBznJpNEfIp
l/UjEgtIpGsKKqciPyKewGvruuY82KwrA4jS8f1MnFCpdB6RWebKOtdWAPoxeWUh
KJtu+v8QXnTz6/XRkwqMLEvDTlP8T47yj5C8oLt3lAYcy71C2NuiRBfnSVHAPkRw
x75/zUFkve4oykEeMui/EP9DZE4WoeVjbF+xT21JwZPyjIx1YblkmfzKfnob1ZL+
aKLFr4cnuXt9PZjclhjkKkv54xlWeEegKM6eW36KhDkB2D5ZXXX4Hp4i7AkaUsq8
04wIUGO48Cr3V3wDu1GhmRFov8Ojb4+PvNqD6htkOjOee3k9jgzALydlo7xPdGMF
l2LgcBh3Ga2tgmZyEWxzwdIfU6/ex15lzhOPPjW+HLS229gvMOIAtp1JBlb8ZbRs
GeZwn/BIx5rXFzfRaY28kGBUF+ra8Fa0bCBP3znknBYRIDTJir/7XHsbOg9cQ5Lt
69trSTL3V5IR+RpgVuLTfmXY1FtpWIuOHH4mDQb4tCf/R3E5g4KRG3iXCj3u2yUP
p0FCetg4+BeXcGztuvHFae10DV3/7m9c8CFWsYoB66ZJ6VCdjfyHHsWNxMpfMsG0
iP13w/ilXtib5h/G4/k7q66UgcvvCC7jfN1Br7Bi+yOFvLUnosXOVqHMQv4MVs7A
jm7WJB03iekW4p44M1gK7qI+v20Uv/1LInY+0xdDnJ0W4RDaFELSAmGUUqmLnoy7
MDXeNyKkijsKLYjhC3TxV09q39mxNmraD/KWTo+KvGEvhRRYg6WxGhQriIMLAndC
xA91D78xVm0aKHPDBAxF83i3ehUQyTNERSzyYG5iyatDj9eSJFPd3mwcOC5zuNLI
XKJrm5J+dXkc/oHvK6RK9lDzLaD80e3TmylskQf3mUlzMY0KrioXSI1rWK4R4E4s
EYnUFIuzrCvk4b9H/qCmQbuKdRroDc4u1AYN0I5UQzeqSk0qywd0E8x1ofrfiFet
qeUa35dgiwfnHqxmkSkCKc2i8oqR4Ph+eTlI7AQxdr6mwBeQU340wduXNd9+GikB
+fLuZ6VSCNfap6QGOEXQEVQ7RyzjVLvfdEGMEthXRBmnzCpVTkMRSWg9xFDH5SjI
JPrRxYvSewvW9uAU3TR/0sdJ+0wXc7WsYxgXJMsgTYijCYN9oApOtXp6b4F4unx4
k7ZrfRkydTVnnzhHkP6rCIZxdZ78wKROyTpei6SPKo6nmPkm9PFfLC7J5Dgi/PVt
9MXvy231/XfPz0b4Le6jxcdy8dwVE5D/JluNATuPuPXaHDd59D7N0FCn/AFbqRxu
qJG1XBXfHLx1DOK4lUpxiwooi9lEDi49P3PQKMr0PRxo33/Tzx66XKZJQeBV+IUn
NgERQ9StUl9fFXsbdxvcQR6FHaYqngGvAXF5GC2Xk+PEkcqaYo0nv+zP29cw38Ob
NkD3XeP4hKUJhTv9WnR+PUA15FTQfTICep6XgzQ6b38e8SA53hg+qr6uKQ/bcyr8
UCqMBqgs/kDAn010Z7mwgV+O64et7QRee5LH4zwDxA659Qd869yy24B5B8iLY88K
2ylq4K8c0A1YThui3ARU5vXpqBb+70t3+aLGYfFQ6FZDt6fL3BGYQjEVgn+26E79
kQ6r4FxIwKOUcXTXbUbb9mxLqfLMZS2kqdD/lWy3rKlC3sWPSDTCVdymrZExXA59
fxZGUa9LKn2VEvxrLSfspGHaMzq20Vu7vX2pYSkGkE72GK6cT42QoWTaBiPMduXs
OeAFEP+n4pQyLSeUIw2hi3ROMK9dkORg9xJkxkbU/EUfxpALTodlJ0wMSs35uKpc
hRkFFPGU3M5UU/UN8N4nr9/tA3D1X5p7cRYAPDhbi7jVl0tTIUvRqtMcOwVkO87R
V4PuF0gxlS6hnQEQFIP/nzQ3Zfd2kjFIskezFfiQ+tSpDsIADy25ViPYgcBar9qw
h1DyR08OsLviUGtocchsLUNMBgwviN2o/uP/nuTfVFH9ZLkSVa4oRDSBomuxiqNR
5fEjh9CZs0BbGVhkonT7EBcNsjmwmgJGm7F1eVunxJ2K10Bc0lwGH+PbVVYCklhh
fkBvMjPwCcql5dYII2gIdnES5bSPgs62uqoVcA/HCoGPYq3GvUx25Lx0zD8oiEgf
p93jcdwgO8Z/54oLk12OKbzuxfMUY/Fv848SFQ/fEyIEJkQYWKSJ6lxuVTf+EERC
x7P4x8AkP79W3j5HIoLzbDQQZEkNMT/nGMroFCrT7RnU0b6q0euW7fx1Hp7E1jj6
Df0bVYlJMD51BJJDrtKWRFjgTJmIWNRamcC+DX60CCWrwhLF0NjZfXtsgRM30Ocy
ASX2txzifNVJnOaE4kJonti6rVtkold/8MPmI/TcZKIuYunEjuthlHRLoQUadN9u
ZTNS4XUw8G8z9Wq2RK1SNdTbRlN8b3Zv05vbI5Bl5pyjJkR9myWUL7ebj2jo0fm7
HsYG8H15BOHAXCQyf5gGc/dQFCAd2LJZlGx8LasmRMwX0Ig6gyWQlgNg39jt1USt
Om45Y6vRrQP/z86NyLdB4t4hnVb/jz7Xb8PCDZtvaJ8Qz7o6Op1/6BBBu7BCIQ2o
1WDazPIb1GdUZXgIjIuqrKiqyZ6ayTeuVKSGOfblEcPdhcaCAwr8TOZW6ARp0gfp
FuSZaQxsxtrHPTcHJFfbpP6R6CaF3EYBSuqbXag1hDLSfbcIHopfNCGfA0FbPYV9
zlEFCkqbADtrrLJtOtHsQuWLhZNqr4J0HoDn5v6RuSBNHifbdvRo/aUdR0QPsIgi
p3QbW7AOCQ2gE2G0QGzctxoawtCcVlSqpMxQAoYNkkUugUEqAASJqIWY6uLYBNA7
dmHTVvyQ4gd0kIAKzM3oAsNFLmFoiBbSKC3fQGmjb12MMpeO3/aevqPzPctsjWcG
VrQ6VPkqIm95vLG9cZlHjECYhNIAmvR26AAMWQnMNGwt/ssyTjIfvrjXU20e4aXR
dE5Dod18Qx9K24l53eMXqnLUGZEUF4lQWfgCaIu9SGcl+qxS3WKuhH7jP9nQ4K2l
Lqi8TMMBC+XhNbdmIyKqJRebG5rJmFw9itXjNms2Ew/zwa7e2NIUP6YvpgkRwqib
op047KlXzfwn2yf2GjTUb522nSRjBYP85LEY9JjPCsEp4o84zHJ9GrAsEAyt1plT
hFexA8wrRHUgPvR673lDf+QuWrV/CJ25Wd+UBg23QOMR+kDjDHn9/pFw2CCpzqH7
MVqTdSIocEfJzdNLE9s6lme5UWvFlnJoyfzLO7gE3lXXkvfYjlextLUwazzoaNKF
6h6h01V3u6yQQpTlnKdZurOoNjf8AxrcBYxqdjITgSviC4dDhYbgw7S2NmmIwJO3
ObXqsQFlh4genHw7rofzjAvHXUKkFd6kcUsO9snHDM+E23S6Zr5n4t8fbVpLm/D8
IGHaPA0sQYOPVOW/C1fKzPuENYljP0MEgumKrvskWw7ad6z1l9GuizSeiOZpCXZM
Fr/LTV4n+xrnKMqK49oSt6hMzoLzWHHvz17VWnY2hore+pRnd+RVXb5VTr6z7lHk
cYC5UJBuyiwG1HcEjjHUTy3qfEd7RbrDt1Th2y+Sz775Vd7OUcGr93FSAKiCMCb9
qy2cEqR0EP4rkodichotLUe7SPgc12dOax/4ubwnFsx4nd2sHESGLXWc8y6b3wPE
YGOBF49KAGXPejQ9SYzq6CqczGyZkrtZlxALmgZHC7M6wkaHjIe+E0eOTJZbFKCl
j4pJUr7Q5Gpu+jcdeSGihTwav/kI4Ao6sQ66hJ3HYGcTWCD88oZ4uviiWLX9X6Va
Q9/SRtuQuHT2IpA+YFs6A0ExBgkqLN47GMcwOvdKyo+wM6h9zu7iV2juXL+QLB11
5GIynZGCUmFMVlS1h0dMGLKp0rbhR2OWMRuu/KdSPON+iSp0TfofTuBpWaz46uoh
EBTz4HJ0ntf5UeN1wkeDlckfgjClLxmkf7ad1D+5iew99z0eazo+/2XRNOxto3Sd
5blJSfeJCOO1rK7mL1RQflMXMqCTUyoV1ZARtQIBknVaDAMHuYq1KfXq2gYToQHw
P/x4Zm2aX58btrEsyihr6BPDoOb58P0vd9bH13JDHqULDvnAvOoh/i7fA8yygqir
8SGDIVM/y4CzLv9iAxGQ8TNfUalC2RGX+PQml4LHxWJ9Ep+0FS4SINH+hOslFnfw
Yrh6ufYNqzlB7TR6mEJf7ONC/6atts7bzWXXx+jwtveZnaLm810+1mFdmKPAPLl6
vFu58kwdie90uS3hJl3nctoDP5kKxEjJUMt8UIsbx99b3uzIREAHGJpXW4Xas//z
5YIkqksFTErgI9BHNHsKxCDsYXhncjpkkbaJoL3zHyj3SsfTkdCMqNCuO/0Or0fb
C3xyT1iJ/81OOlJ/NA261cNWJKFFlevKPrwtwR5WXIbdAdPVLWIpeXnlIM6VL86f
5+9k2mBWQJpJ7rP2BSCLIBQSlAn3rlXjW8TrayNWT3AURF/2Nrrm7itvIx9T6pVP
8GwPAnT1gdgpbUiuJuJ2sshAjPQMPeHlt9pRlaoNQwEMfkna9GuIpySmjcWh7Inn
wlruhjRKOWq99A8SIT+az42ee/CQuPx2A4CBy649m7qeEydSHph4NtTIx+AIZ0VP
ZZxQvwwXxiaYvn4/Oxgy3niaR1/G3NUR54FPBnruuuXVDWioRVygv/xPZiGSyZX9
FEEUn86hcAPCqPalnuSMArVm9IR4dzb3Lsf22gHOglRu3NkkXf7baRCSwLeaV4sY
1ySPdmfpYPm7YT6wyixMswV25ZeBUak26VeDmBWTYCaB8fChvWgT0wzoHBXuaIf5
yMNUaCt0ceOHd603or/vkYXwRPDJvlUVpA0kXh46zFJtt3d8mgpZ4wA/wWQEzMhO
V5bfk9IcyUkbJWz4YebZKqdyFYtiOLwuEz6n7C+FejykqxqX+K24L2x+YlQZzfzi
iKoHywR9xRYOcVH8mDwXmCQjXTRjiZ87l87ozisbxvemve7QNNSJDvxmLiJJwG/o
Vs616wndCzm/HqdazgDDDsxfI+a4KJBNZq0a2Mp0X38Uhv17WGdaQLn/Oj+vYFRy
j3RKXxGNgc+M7LmYkxZHVLBtTWDPS3Ca+IVX22zg/PDf6ofR1DHkJUMqB+j7hNd3
LNczOjkc5KxOw9NNpF6PY09pfIahSmDKFJ4XSuCmVeLXHfTH9xhEub85Heq65FLO
ybVxrnpNqO0YwdKEyO78eeNN0J7/syLWuD0H/mS+ABtgezwbdI4E1H2SGMLM4+PC
My7VP/+ta7rSGbIxqG/6K+uv0LgSWxWcpMadWjjne9dawoFChx//erWQBQ/B7cQe
iUQi5SxFuzJRh+RCOHkKC8yKM3q1ajFxWxFwAxx2yi/Eh3WGcGoiIBYL+RamFkhv
iKye3RXOvVAOVyXDGvV5NP64fTAgEJcx3DeZKWnmNWrK3NJLjsgasH5bU2PmVPDp
JV/j1knuAqzZZSne7RkmbX1u5XAKV1kHVw7NoPJKKhv/Gue1fdZdD4hZKmiTxhzl
idkIzcOCgPOjN2O0+28aIP+U3MwtnrNvnfXJ+iHH3DCkYm5Y+sj4qyvz+d5QTAmx
sx/9Bq4NevpaixZytuHyDuuSXEjnegTqGV4fn4Gb2t1DzVPBiaG0REXLYhnsAENd
6uEZipw2HM/ssSbieQ648IXRHKTJhOZRC7ESDvaDE7l3YCaP0Bp0sQeycOkA1HNc
Ursu82Mz91/cwhGeDKOOJ15BlcTMFLRY07aMsXpxBw5vHcVkgA3r5hOArjO+BNWy
yDNCf867ad5SgEr+WjbNfmWNfhG4oobUkWGKsm2fBcinCiZhJG9zcZmltr8G6dEN
PjL8sA4kEdFXFW97h1ml8CiJ4sZ0AOhE99UNB9KkL6fqYkbw+gN7bIEAZV+MBk4K
ZiqF4sQaBDVeaU2/MW4xYeDt3xtZsLQrIubx1UBUI66hBR97FvfOHM9+bVVON+UG
8/Qfqq7uRfoZCkaHu2CP+6Tel12owcZZ6VJoPeXHM5qxpm+4V71aHPlwu6RSmsbM
LMMm/BXYjrr2AHTLVpmdq4yb3nrHJRw04uvBegNUl0OhnHfOofGl2y8luI447CmT
Quv6uvdv+RtziGEdss3YPePQutqP5iJvI7ycgmqVHfVtIxUqz45e6fm+jlFIcwj6
8FSl1cVp4DhJ3C9GhmjTNr1UjlfMuWRgobNz7PGn0bxxl1QuPW4oXfEolCyC/rE7
6zboW4LcG/CiHEHkD+86F1CgalaAxoVk9JmhGSpXjjaHx0sK90Dq0jtuDlAibB5q
/NqC+qYwOa0FqduK8nDDfFjRWB1Wqs99bE2up3wLh3cSKccb14+uveE3yOYfvIMG
zB3yyCNOtXfOStYswjHwSbTvQYWe82EFncxV/2FXl0MzZefsdFoQ+vSDPsgi76mz
sr35JbH70X1o9V5ATGcwfBIaocjKg7/JO0TNM1z0Xv/yHel9+MnOGLN5BIEe27uB
T0uxHQYolr2V/kSKuOLwy3KrMtX91Suq5hWoFYRH7oDdtoxNYtmVXTIhloHOEX8G
lu9CGDa4cKHUQnL1Sw5kyw4iQJBrTIIUd9wgpMrSBX3AJ8Nx4AjBhE3y0Aw0h2vf
cm2f8szqk5DzGiU9Ums5kBRLS20wCHUaLdoOQ5PAGuwoNW8q46Z02Xetu8YEbBVQ
rREmAry9Uqdu8piIan5mUYKD39bDvnW1uvDUmsFxqKQcIaxGg/UwdAqDM6Sv3KxC
jBCvlvEsg/UN3kEUSaH7Eg82Lf+kA0FmACIiSr38ljvl6z+BfzD5YhaZHFTiUR+i
jZH6qwZQu+iMHbUE7EHggY6LcC95Emo4n7IjT3eLpx7SF+N6zwGkBqJZIf0zCqVn
5ZqVqnEOVupNfp9djnjoIPWF0C8h62CgHwed1Es+vkl+DOnrp53U/BYzFDh+UtP3
ZCaqo6rRiUFVpRDQ6ZwAHeQidm+4X3lMjGmGju5AeuBFCOAJ6/gLHYnnS/Em+Tgk
Ie9fC0073VrIrRtHng+thg3wLfSUmlNIfUbXh5WjErQfdzfmKdO4PtlKheaR5V+F
azMzQ7JWzRYwQWssWap0MbHOm9n8L0MXnqJJu7AV/xwjmOMhoMlzcQGXF8+vSxUb
ezl9NoyYee8l3e0t5cyborWbsA/2HAaMDKvXxVOQXXBAoREIej4/npgdaMzfZpJg
UemWwgIsKehZhwJgryZS/VRIb5PIYkZ/nC4H5f378qzIbu7r1rUj9xYpdXuc6P1E
q2G3X+hrgv8D//CJxtRTukcC6Z5rqYrrF8xxR04DAjEiBv//Nh69gZQ6lxWWwbX4
U9Ut26CQpvAxnww3ixnN2GzlawoWlXhA5ZU11toSDPImmcmDD3HGPQKeVwjFFz2g
cBTSxtx2gUEOHYl4L0xvyTY27/tCQT80NedHMtRLQ0cjnAb+nmObb+rCPiTAxlSd
Jg4jdJ4r2d9wPHLg2pMhO1hF+Hu1LKurEk+A9uy/gH9ThDJg0veWyCX8wcpq7+gr
xspIInhvL2zBr2gQWeDtAtVGhC2dE7leyMHknhTVxBx+QRiPXo6rBU2gdzyDt882
zQXICtN0weAJBx0g61roENDuUIgFP2vGKro/fzHnomn+TpkFahCuWd8c2rO9+dzz
2hDRmbPB4dWyM3Q+YT/DlBGhnWqALc2QdbpM4oMhSsvyCMzxUu/dXAxwA9HBDXLO
aMOQs4KmOLd5DX2Q65hS7Z66qgtAX69l10qCjeztxVOzXt5/UhBpsEyJdTP/3wPf
ti/Dv8R7xh9shKhzXkGnZcnaZd1MHDqNx2PAgidy4ZnObZtMuAxnniit62qybHo0
O58CALbSENRYBL9FpchsmVGvkxfkw6/nV06fqd+y0OuuE927bnhKrR+YQIobxIUw
WGXCIcLZPcgtlCZJVBHu/V8SOIWv7hKfY3Ksdz1lBAzL4yTfsh4oALk4/qzR0Nsi
iz+97vTmNQppwiD676tuFECeL4K2c/9z5eNKzhze5PX2GyYS0GB7K3BA/yr40dSx
RyAtIeivBtXWK1a+g8fDjIvTnik+7OUOH+lTTsSJMU5JQmmNKhBdbb3C9hQ9NCmW
hpPwk0+OEoIt/4fcc+OWfpdrtraryUNVuKWZq+4pUhqMOok69A5lF8bz5CgAWv7V
vqsxHDncJAKuWCcuLV5p66ZaSrbIjcAkK5OrDU1czXRkYdbOBiDIEgncILCctMk2
rvf+H/rA59F46Y8TbsSgo99z1Cm74Aso1c9DpSqG9BzSkjtIqZW8L8sey2lXoOIx
9x/laghwFkVhit17gr0QQz9XwtCYM4AztLqreA3GSDzhJOb2cQMZBcEKu9CKKc72
v0wHKDXf4Wa3D1cb0LU6bHmlc86SRLsmLji6Zpbv65/R5zF5UJIatj30LRofPenk
EKg9+LqS2ABolGCONHKmR3DCQrZSPZQHyWEhXuLbmnTX7PQR6wK+Y2W3nyI3EiUf
RY/lnA/Hlf7YN1U6M97/7eAUZOyeLzYQ3PxuH8Nw9gV1tszu023xh6Il5pBDIw+V
m6EtjSiJzGNuWf1TLFs3O4Sy6XRiVEhqYrqfreEWr1wZii+v4OOFkytKfn3P1lmW
MRMM7l6SDG+z30elM0/rbLwuG4DoBuC2WNd/abED1yqm4XDNAtCcNx6OH4Ll4iLO
OXF2d0ItUj6wlKu5r3NnfqOrq+Mu7wjfm8dtpLgWJsZuLEij+gb3uVBZWAS+Bf9g
QC8qoTAeV5yEhCj9HQtN9HRgYUPnUFzovJKzd+MbwbRbibe9tCEpA39/Bx3qGJyt
DPeq80eBJ/Qm095tRRrHfSvB/TrOcSqtq78rPFgo2h7KzRtYy9N8n34gD4p0XNjf
TTdk4DsqL5FJARUigEmsiJKOEWnRgMddI/6973MWRrzxT5c9wQaWerH0iUmJTggv
yFc6MdZtpL2t2fR8mW8P/kbPGyGvvlv479TEqvsBqdbTzbhrcf+MCUf1ejvJMINR
ZCjW8k6HIrGn5iyUW0kGgPNVHao/oH2Do3t8Ex+/4USpxiouXjgTErJBxKT92arU
c06giLo1aq124efF1OLkhLZRGws1cSI1gUThj1p90120tX0+u5M/brPuZ8GMs1PP
LvP8Aje1oOL55t0U0BatEdigulKvGJZDIS7gJ8PGZrVqFll9fizGqUjO1EsaNaby
7y2wYCOpuX2cjOvqoXY1e2uIZkmMf5yRPCz6zeoAkPworko8FPrvtz07roqhD+oB
zXwpM8y8FNHT46L7vY5HdW2UhWgLCGJQJ8AdaJF80Y6JUdVaYDjFgtDqMY9MzO+n
hLeXV6bd9ItQJ35EwMjG7LzflCcVjYsniMyVRIoq5ClbzaLNo55Y0HvwCjTV8OR3
M8y31h74chZOIyGzQ9z0EZ2DXkqykzHZJ1ofIRNpiHHGzW62k7iB81KPGQHfY94T
WRAxdlFw7yRbrFpH4dAo7i8qwEexooeMv02taLvFoqwLWP3ZBbgigoRXiZ8MTDkB
4Iu0UcUv1RViXM+y8B/LP4e0UIprerYsSyZwpRNFOS6j4ha8QLaRZDvfL+0bfBqr
JBY98yiqrVTZr6DJzxOb3N9Nxr8WGyhgGwRB8qyK/6n9Sg/YH5/Yp5WNMbJG56k0
TnGz3mdgcmArOwjm9dsl/Lh03hARsAJfQx0puyicOr3+idouF+bshVsWGW2HV1ax
AMB1LJeB8eVz4q4FXg467IbyUqJ4vpBKkKhwJ7IdjbBkN8UkydT4uh8WmpMURw72
IyUq27ga35VWOnMDqNHNByICeUDd+qnLbFGvCPXt+lgfX+AzOl3M4GJt9vw/eo0o
bRi68fWUrTgjMCf1hYbrG56GvmsZB1TZuJfqWntx0mCOID+Mlq0SPzHLWpGeOELg
y9XyXK6BssZdTmXcbX6TA5zc7o9+8k464hgH22CeKuLK3bDD5DgOKQlTP2VsG98O
3Fc3GiFRQtOpPRpi06WApTFkQo77XShHHR1WLd/4O2kgGvZSeeLxPlCAE43WIwep
LPHEvICmvd8PNT9eF/f7OqHrnYo35qwIANI+fdZz5QCCsxDCfAXXnB76eO1pT0QG
jsj6lpdzLpIoSGE01QmprA3SR8ormdNgtY4dJz1AJp78OI0hf+A3mZ/++LX7289Q
VghkpGJ6YWaXmjJ9dU+higE1KS20jqzOsxXB8IrDZmU/VdVzOdrU8pav4cfMwjLR
cxAJL38EgXUMoKyxy50xQvOEdbOmEFuRjYbXNRHsqDs4scS2sFj/wQ2TAWW8Z58i
wXTIKun00/ZAxK/k8vWP2STA+geYkn7RQcwKsUfn+x8l7MlIA1Zk4+MC9IngBbzO
odED3FyLsNXXNYT01iW72xDDC43LPCWeRl+uDlEshYYpQmLs9VkBGuAxEajFHewY
3MJY+n6/s0HFDpuWjCKaM/glElTYM1j4S0rd6k23A9kJAdnQBJsepdKBsK2XpBYr
k3AxPDVOw51kc0E92mcDMDDhs//1j9P4G/ZESFO+VbK/Q41pl8tsBkjpE7IM969s
N/+0eyo7RRjERL8Jhyw0m+O67EwQzjtNqN2Q2GAo8zoa4/6XIwF3/6L+SswxUznM
/o4vxrpb9ZsnamQKO5bzE5KEHlfrIZ/PYzQ74Cltin/Svzgo3uOCVKgrxiSnS7jz
cHlEArkdHHczcTqJ1DhC8ZIAp9h8bX9K7Yv54r5KTRDOAURDCA9DIVSbuoLYkflw
iFuwWxhb69Tu3tdZ9P6BJ6FvLNuac/qZbzHxldfUgDbyYn4CEh4FJYUv2Joi4uPm
AOTp8m6JYdlDqZgLpI9Vo4nMIukB1z/GBl+ZXgkufv7uGfPmGG6l0iete5ScOyTR
3UGucD73+6imCpuVScVBKj7Z8mhRx/dPxwlYYZIN/kO5xjUrXNtB00TgwpeN6ReD
nn/32eefbHWdtFSkhw/Dg0ijs3A0vetccFbTDucOVYw4EOBpy14m4uZvLw1IIdWa
1oaG1QktVROTSFkFfMPY1/eoapQCvZDKkN5dsJo2F1Kiaf+1rY9r90wkuQdbydnu
o/YsfZKXBhk4zYrN1sFp9hfSWimGpb9sMxl1lVtit4Kg+yqQD8ItiO1XeKx9EKz+
KF3Bpu7Mci+liLsftywThvRFEv4xLwm5v3/VtS3Qn2XoGaw+ERZo+V+tGtqa+GiR
5P1rmwOezSt+Wcg2EoPxpFweJz0Nxutdf/7bD1Bb2HS8hDDvqsefOquLX+Kr2GkB
CetDXQR9eWUWiEjhp2zhNi9srJBWHh504zz0L0IRhGYs8YiHb9HnOrUPaMS8+/3G
KGrDcchC4G5hj1Codg/eSyjUovaFpbNcXJV2B/95sX76r9sd63MxEYs5TycXe5sN
Q/YQLT/6DOZ+wjIleLzrR1Gq22AXJLTYi1m6DaVJ9cheqy09CPI8Y7PasgewtTDt
9vKIzZ3vRJ41UYe95LD1DMqNO55lFa29aAGKt3EOcw4dp712rkNqTlVbTRhUdzFB
sODvFxfh54VG7IYj9O+g4CoNsUe/wSjRJbo8Lr9051PJoYWBzCvm8P9ZRu4U+jYr
5t0mVhca8VAH6923nOZPwRuPsiaydWMTX+qlApSRhgkqCkLG+I0YWbYq/yuXYpZn
htNc1UWxPBaStumsw+REAKPYKfwph68xfxC2uluKO9C5B+hgxRdtOuTO9D2u0/HQ
9B2p2PWzqnaPOZDhS/XdNG+cs2YB3dNlhRi3PpvGRX6iZn5sbPUhuP6uFg1TIuni
Ho66BxtbcXoNUZFx0xPOdSsQA1PgNo+6kmJG2/1Gy2wo/THziY8ymf/qwTbDubtE
kvy9FSr5u8OGAIur7CwixK5BhYFx1ScyW71KeA75uvUUUQqYaLpqwvL72eOdTPf5
QjcR3xXQISGYpIxJx79GL0gkwUd81Gca7AkpP+7ScXYnyE1QvZdBT9NuSGhWy9od
ifZuX/mKfgW7iaQrhUlji3EjfRM4qEJu9lkMhU/0AVTsEyvKv/dSx0BmrwDehdKr
q0fDkYrQ/PVH27pTQbGjzWsOcM6T3DT51X45T6VggYgOILKOfarIaELYFuR2o7Td
KWXhHtqA+Vo0UxWKkSkG5wpzP4nkB3tRX0HGea4KFtaTXGHZLw/wls/s7FSt3PPG
0hnmmjoroqNeEiE8WfMpcd9tZXwORzPKd5YdXI9jtBiu2APA44Za7L3ki2FsXexm
YQInuN+gAZXmJDv/liuwx/eKbMtQos96WfU+utv6aM6W6XF4ybaRzGx6dK/QHxkS
2c1QY+S/UJ2E6TllzTuNBviaZ9jkG/n6nqgY7uOMUG3yTB1Gr/l0qPu2kPCjnyO1
+1oo8HzntnoZWOGbOF1bpUAQCIxUsExXlQemE0Xjz6E7cLh2vC0845ctbwVdEPcK
kLN/HmHwZE5WbUCBk2Sovq+vTbowBiBSZMBeIDvjM0g0sC2oQcGA7vytNlJ/DPZ9
LgASj3qp/Wotq2PfyAqne2UxokRQ7zSVIqUBwMIXviHTC9pNUQNfbRAGoXvBlarq
qT428WsH/zo8ya0d3ffboQxY98kF2Bf2/o8yDoBKkthX8p6LUj8T7DE5FRQ103Ts
USGMe93X9Ami7gUs19wl0gODI0L3xL0nkDehf67t1CII1qqEYQUcGtmTbnhxBd9r
9WLG7+UGlyi+G1z7QB+zu37A2MGyEPTMaEkfVFv/ZrhlhrfV7S1TELEXesMsXHAt
W3QXUkKL+Mt2EX8HIzdjR2M6M/+M2bc8IrHMAGzhqGS0h9/hjRAKTAu1Wvmw77Bf
UNm8f99euYADXVTvEbOArMzRBPJPOXtG/LoFfhJvj+2uQpM4EBdNNKd16rryQ8vE
y0YHP3vnGT4XJ+VPvArDqwwM7gSkpEk2Jaydtwv5w2IAj63Kne49qx9GWo9fd46d
TXNsAGCpfcTl+BmfX021sGajSWgNtDjGtK4WyTX9LM/27j3e+V0ce/2l+BqXmZuW
acgutMtGoTydpfAL2P2L4mLZolSv2TTbebV01OMIsxMKO74amVz4UDq5DHu/F4wD
7fdXARaALIZioj6QJlJf9QfKLE19MdlIQL1s/ovqkwyKieUwc+aUZMtb4wP+5XWt
769T7DwEeR4tWDGjor6jRbsk1DZFv1kBtFHN2eS2LaJ5clHzEbBCWixO6bYB25FR
JD49TIx8XGCSDHSmWIvN8qKlVX2TpAwsKd/EXTTYReSznfo0cljRxV/Z+oc+nuth
43xtszvmZnlNaMsbP2XSkB2toPZYIl/5HWO7K/waepv9yNc9j5hEUI8z6E2AhBri
0bSvTslJsvGFZVK74Dg9nITQ3jjAAJSlNAvb7iy/JCR43UqM1a3/JDjSXheUSYsB
RmL5lKHQQhyZt8y8DJvViW8btVkJO74EkpUYWuuXAzZZHWcCKJYKmW9ILoyS9hOL
5OaOcV/rMlbxEritFxhJXdCVR/f2Ug/1G2O/25okFtV++9Wbj3hS8PEnRMgW4xcQ
HQ3TJriEk+1Jbx+dVJrdtc7XnCtynDdARA3a2SMo3CEJpNh/CfDeVrUpotpzb/bv
Qe1aTBIxYXGKs1NPRdhqpG5NHqOEG/HD509jGsRMKWbucDfBHoHrDn8HVfpt5Jnj
1LRUe69iF0PNCZvSj+8F1v91N8AZdyI8BO1vzqG/Bs4KoRG4rkCTEjXRNbfxT4lG
bcoaA2T0sw+ZM0hAde81AngneGDXXqabMlrIltS+TRGasqt8P6V69hucrdi8zKOb
7+NKIRGYnOTKGkbuA3viH0hFCtUSoDk5uK7xdz+ERK32qp30gX96TnNP7efCnPag
VIjm3hhHJf8aqu5F/eV1E25+9viM7/J/tbOlsLjwZCgeo846oeCRr5Py1PS5d8om
kUg1+ANiwcePnQPG9IYiqC/6hj7nIowJOar2GVxFYTHfSCNc7VB6uTR86a5qn6yv
iyEuOoZM41P/4283NizEwx6I2bM44EqDdNcwvvP10mB2dWGM/B9Q05TRMVpLweWd
4FTOp7pFFxEFhyVzNw+nN2XGAalFvRDt3fvVU5RXa9me+hs5yZcMOBSMM0DHgd+C
K9eug/U7085OJYQgH/Selb4EbdItlQ0QjnpbYTE4DHBNjO/CzRup0VeTfEo7Jp1+
uqg3AmAL5aJJvAEK1p3siYrS2ER5mqWb8comQ7YdHb8eQvtmw20SaGP4/fb7x5/J
Grdp0Mas4q5kCKXla62vr6PxnS1xnf+xPHy4sCq9hMypju+L5U098tM9zeWdOkol
/9IP9etqxYvtm19MpIo2AyY3+Y7NpkQDoP0MlZRGCvuD/wrNVaPEaXopAvRp9eVJ
hWnEwT1NgNgxPWn3uCcMmPeM5rUuSwiz8mSkF2o3u5oPufCMXeo6u2cRCO0K/pEa
Yicwk4IPWX7dhOJRQnLoxQIeh7uxD6bY0BCKSHwMo+Yoj3/t5R4Y/6C48Y0lJsep
7E5rvOx6RuTVB7Xk7s4Fw1rb4netG6aq3FIFkBCiuFbv4PfVKneJEL1/v1PsqovT
s/LTuD6auk5qOGiQY8dIDHd5wDvODboQS+RK3oCsAnECKkb9lKyV4oyAFH1bG7mp
EDaWYQtm7j1iM0dxkHEa3s1p9jOX79/czNK5cuoifdOkBky5oluvNHVbaytuKOLe
n6WlJMYnCXHK8nHR0qBKIC7m5kzoclLQ3WuWL4jjP4TKy0BpykpLzCHnKYI+H4Hp
VmoDnTZR2YW04Q5pil5h/AOl/nWrXeff0xSGs1gnHqcEfuk2WNEaVtqjIXk46tWY
JW8xxoy2h3KR+4Qg1Gr/POsCLJ9r9vAnbsEdF11XvITKbwe4NW8ipjEKWmfL9qGJ
sZTJbmUiWZyBRStZr0bTMHuZ5R8TXfLed755ghh86VIYDTGDdyxQBq9+JTXUNA1u
v0J103zM7HRS68Du7e/ue07m5DuKIsleL67flx8RVAgxPwEvgom0/chk3JlxVY+k
pnQQo/E74cfuOY8BQbIL3wBkjMZm3cGjO3QyDbnoanhJLPGYisZCMC1rNog21cRq
IImHT9ImMqDfwjLCvB9H1CcwgeegIan3GJHgLvCz7pjfnDY4RS6n6lNr47ydQ/6e
CzOwxcMTaHdkSXy2r9NpKtyTa2sTzQJKfGnqGEi1weQ7tvQLUGAv19X1IN3kMoSd
9N6PNt2hZjyNgl6Y5ENW82F8ibVmd0619h4+vsBFciWPTAWyv296JP8ERROLxPRC
+2cQ0V1aBwkPqg8BGFCeJ2kWCDS3eUOto16WaupxjTZTko2GEKPkTi6GoC7A/B4b
xJRZJTwDSBMgpQmEQkhBPQjsZkR0cguCuW2sYMnwNBtaakciJBnIMki3OoKse6nm
4rQmpXZP2HWaSKV7oliTVWLglU1t0p/zmmbkDTFgnvxLtVIfFQjHYN4RUp1A1cqb
4ZDuF7DJFi+w5w8tKlYd++wbOLGV9d6tC8ccgyLTsTJ6t7quXYLx8hFrVCkaGg7W
XUi83k+teHffnu0AlnTz+UMqKTN/yE5+zQIyGYUMgmVt21RTmOguZAZXCPHB+WlQ
z8ZlosKCPZuZKiU4IoXBENd6yHbIZLSJC4CV+gl9IpPKcnaaUikjcsjjATzgdOam
b0XFcd+WKlgCwCnocrLe895HT/yFKaxWS/sbAUeEIzkFntKEzCI+JEu7rA68sl7j
ARC1lHexDzD2d1dXo568h8juQj2lI5getPgs65d/pIYpR6tpyXVGOfDlcq81qsDH
uzRD//M+Mg882knBvnLmS/Gd5DC/oafzXHmYxICluxSi1KySw/cFQqAgz/a96fzk
cNKgfpq3yUhBMMP0hyulhWn6JitGAum24oB4t7ix6IhosGh91ApyHnVhGrXTgNLl
1ZLTIte42ry0SOnKQ/euK4MX73wSPn3+el/MSDdGj4IdS7LSTclGG24wkHxR3fws
6PxYDTI9xG6AMt0m7T8a2R53vOeJko7EJBLQSsUgdqeCZOfHpXWFXZpC8PTk37/O
iE4odrAkzo0AfH92Z1AqQAa+EY+yw5hWHVO9Ixz58VX63q3TUt7zEFJKTnMuhi6Q
Bl6m64dsN0PZhvV/2uI4c1IIukXuprqOcsXVMYHrxZhFo2bulzXzIpP1phiDlHna
dXGtQVahYBVXtlLK41FblanFdcItKaJbjwJ5kaJQGHw7gPxmVSc67ICoW+AerIs2
cQCD143AO2eNPelkc6Zs9wyrAw5IQZwhwXofpbv42W6UyhEX6IrercL0I6fiGfrZ
cDOC2OfHdM95cp9yKZdLuJ7bWowb/CkedCncLqlVJPGyLy6FG6JInwRKGcbewUrN
gJqU6jnmaNBmyHx41armppTmkcXzEa0nKd6AE7/cgJ04J0YXpQqY8qYU5Yjdtqzz
66TvN41e4wPdDohPSAgEdedeO8I5lX5YQmzWjsOJWHblc5p5ge50EiyAfkDMt1mZ
b3Pj4Y27nibvJyt3Iqlu5MyOlgfLaKiBBECxIMB9eB499l9caiivMLy+iWbe3DTa
1V3VOOearFgsRJVimSEw1DDNatoO3hstKzwma99f3b/+/5zyf8DOWkoS2RjhIh7s
f0ofdPTOdFC0VFMwe4fqfubAg9s9gLOy45nJRJVJyBNRlMq+9Ca2BkjNzSnLetaj
i7QgNCWjw1oOGegWTsDYKZ/bmIwHs4Mcg2+B+c2OYL4QgQOn9t9ULQb3mukBzT+I
8+z8hGxxI02Q5B8plO1Kp0YIkUAbBH4XlAOkzYeHLtqgbYmKqWyGoGu+Dd2qRJgp
m6teihGzbPIrwN4HG8t/atHkPWbAkgUffVHl9WNakJReAS5AFNHMzv65nTmBfBLv
3/0zRDT7vzHV9q2zCeeruOD83AuNvoU4NW+VNs9MMYQQHPqveKp6fyTabfRgavyV
d+XSyrPOlfpGIIEfNZpuI8z04TUr0gzRt+VVb9HeUdEcaOPZKwHBY38zDM4CAWUO
xwXjFOvMkzldb6SNjZd7EqLHPv8lJMMZ1+I+NVN5SJpgnQ58mIg6wQBh37aYwWWI
3MgzvUlKLPGexWxkw9gVDC8es4avuI+dK0waXTt/cAdzumkD0QQQ3FcV/kTLQTxy
oF/JoaV7NlpUHc7tKX7Mui/+D2s3uEFJlP7pHR3SCbiUauhK1tGGqrZGBuC2H/A6
4FqRXqCFIJWvzymstdFMavdoo2uM6w+wGesqELRjDic6sGSn9TZNQWSZ8jg3XLdO
guNLstP4ytDPDpacesafQntf9BnNwfhZdN/J8N0AmTjh4gUGm4ux7KXVcLTeCab+
aqFrqQjlVinOUYNDPFi4Sz61Bidorb0sz72JeYdGPVVWDotP/WPBAQkZhiOcPx85
ThDtQk2lb4yhHuZwE/7H37ayuzw1xX5n3rA6OEHd9fvvo1T4YTCJGd00cucUNRmJ
lGMp4K4H5K9TgLh3rj8VRs50POVzfqid6+WqpyBFyRxYNJDbT16uIDnYqYXAT1VJ
mFTZSoXsFTFS41mCbWRhJQdkx/CPjW0hSCQYOsyPGAql4G1r9CKvp4fOik2fO+O9
UOi62uRtGo9oVnnbdw/MYPD1pNn4D3OC2U9fJt1wCN20bSSvz/aHHflv5iVvnmMW
H51o3kNgZE5nOM73AuDRuptiFcHMjT8JRa+1HvdNgHDrSjTVNGyRZohUAl8oj9fD
/bnCvZvDQGY9lR8sCTUX+G3DbCVy0xlMqy9BvYwhIe0MBbiy4tkki7WXtGdjVvvf
Ls8DSzq1eeJ0L2X8l3Wd3GgeWgzEA7NPG+1Z78lG37ZMkeuFtTigIaLXSjVlR+7I
Ew9XZ+ZJwXlgX8mslwiaNoscWPDtR4oU9H+G+P+9tF2KyAjVEtUYA3NT0Lzff+zB
c24fOhBV2gjUICMbcrYcpkQR4luLM6yZD6DiWCU3Qb3Qa1GBNKasCBaFSrPMEKBn
TE3d8cstkylgBwc1WcfJcjcU7qyraQWXepWFs0f2hPOETECENg/pZ3S5sppWeU8m
8T6aYwDxQTDvbyB+pisBvfknDWHUpW/OsKi57fXNDzemSGDuZgavLC0/pg6RIxcZ
No0BDCxzlUg6PpA64W33exW+rBScVTuBc7ACHhfpZP3jU5nQNbFFKcyfYZiaf2Fh
aHpuqNzLKh+lglsuMh6EVEMIfc1rDJMsSLNIHE54H9uLdMRXnGMAXgogIcK5ynBI
+AbKOlbm1F2eLVI/PdKWqqODTr5PwCVFoDYZ8nrEjHU89OZVz1AQPapqrANy2DX9
dfigaThqWwY9eafxmUUdDTGvnBjtq2v9xgN1BuDoNFBa58axhmF1s7y2+aBnrUgO
rtIbhypIHOCl3cEsMXNAafe9FkafuAl1z0f0jbav+RhF2ZuKnvBdDNKAyO5+bRmY
2z51HmEfSrhRBgxIlQtT43NF4IkO4XRvcLzz8dwM3MEdNpJokB79GVvR0jsB8Jes
VbS+R3v0bFV+TETQATytDoUJMt+/Vv4rj6wBpbIPL/dCilxwTTWi5KjoQz7Lgiyr
W19n0jxKNznTAJjZjbRkcmWytUnOWP2nWf2bbxFM832ThrmK7cS4nVV9g3iQRozQ
bq7anbnRoze7jJexm5GGX8F/YfvN60+iC9tpiBPFJ/J+vP2xFLSVZp+BsK4UlLkW
hKZ0MxTf8ojbw3zn4EnzZsNj+XTmPZhgFhJn6ANqcYQw71sz8xe8/O3Nkm6m8SyG
i2mRLHITaHGXQQdkcNQ6Pqn9dswnGDSEG/5Iiz9T93s8Yx1C9Ns8x/zT0LwIfRo5
D2AmwZvhRDqcCTt56RXv5s5v+C6g+N+oRSHTZl6h5V9HIdyVN/58JcV+hkxjodzT
Y3vN9osjg59/xwuxLBpeUDVuTVzshRpgFQIbkoDMPM7HJP7uuEkBkrEFvWa25K16
rnea2RBgXmwkNr2qsbljjBpDrfNb+CQZyXm8qy/lTQadDt/1Vi2SBsiKCK8j9UzS
KMdyjNVFGGTbrrNMWxooyi+5pQXsSYkb39zyQCAnME3xZ7NjoVjGzbtPHMIFI61k
OIBA8QupOAxc6982EzgLRHwhOuH1v2LQ8qNy2DbGPLcdhBMRGLzw81R2Zu7/MSUx
j4iJUExrnPYspmmBRaFOw6cNmxGRhSVprr4QL7fYX3rR36DNLKW/5ePO7JKQAoDi
ZYSr/WhPtm0MFzuL979zineGOpx+KRW3Glc44xzQTdullGCIFR7Md25MmC6WlA9I
p4MjRMh+wTPthYpX3POZsq0YzPEj+Q1HYN8Kc4PRbaOJBlwXlMicKJKXDET+Goet
bb+fifzeW0J3umaEvF4vi97hrm59zOiJv0ESw4vwYApvroxkIwBQNLWGlSVOsjbx
MgR5P210xBy+SRiyiIyPtR7yJDdvv375JdfZ8COyTG1ngg0d1lr0SCv3qU4GhmRZ
LVAtmEFPvTlXQBTLhkU2v8MAnrjVrSfLZ5xP60bSdZXp0zZuto9gD0amy6dQfwOq
+HnFAOu6H8lf/llLAml7ucbM0do0PVPRsMdCseiDw3jQ8V7PXbjFaBaMhFmyUQj/
aARZ9iq0aVqoA41hkARMXGOrhGNIYIRTb6MJiL1CzvvuL5bebIZKXBykYZcPH0nF
U0i9wSsby3HgAUBztPSkL5fYN/mUCuo2M59Fp6L+s5T0IrX2wiL20Mrz7v+gE3xW
GF2SRUwhrkoGdN5G6ZLPkGJw4Rbinwrxjw6UODzyECsavg8jVvZvSW7Ca0v3Idvl
NyCPPCmIs1BZe73rV1AFyIrdvdGNBxMOq8Ji/Ko/0MuxBDpMoepDmaLQSENtKDde
hJW0oY7K1BYPV5sTPv1sYJ32j25BopO0O15asHjJZquCO6pAdHUfhIjTtfhFStfO
+dkfyY4Lkd4hawhnNoqszZAbGTWEuXub6dZknViy9lwPRIm/mV4sjxIWPHRDmRpi
UccoB3R4f+vbyEWjxUUSN9dQMl93Rid6S9jiwu6MPlc3Kc5tpMxJrhIV6clc0NxN
iyDrzFJr6S1JaT71wtfcHtFq7rf+dxS8dPXcNegUL5vzGwgRNEe27OJjXflND2wW
8GlXpINV5tC84CW8/PLnEltHOwOty96J/pk+Me4eysDSsnVtyxTh0UTrHfCvxlsS
jvjsAeYOjfoaV2BO3HD99x9aPn1X//pGx3OZdO9VSXfOU7CXRis1IYK4TJcAWfHA
gE1feHiy81ZZwFmyfgN0vj3A90HUcB6Fe+F+aPupsjWRFZAJ4VjzvFmAV8zUYa9I
SS6pXOax+nz9ATfiAwHugXxS38F2GUUhn+DlHEykERWetmFWwtE7HDYGuCULpobv
+SU5Ci5YnW+JT690Sbog1ORIohlqD6BL3XKVSm2RmNBxH8qoH5eMDrp+97y6PfN4
3lsvTyMXMc+/lJCL5VNHVvM8H2zfvb99RPvAfpWVuko5056X+JG0/S4cT4vqW2iP
0gTpMuZcQsflnSoVHbqb/36HaAQu8bxxYGczZl5nb8pj5olxmK3EgNALS4nzfRUV
82FSv3cjL/B7wc8lJh744sBdit4YPJ9Nl2WcpufdJectqANYRiSy372PjjcYVH/G
yHP2OgRlk7dbHWMf4hlu8RvPX9jqRnopQdApMH3fYR+ppbKt+8GfRCHciEreNY54
ZZd5ScJ2ak3nMz6EEwNefAlIxQxbjqvucFR8N7yKZxkzHRWTG6ZywaUTU6k+ycsC
JtTHYko75FmIEogfojlal59HucM72+4USJAK9kJQVdV2l/PdSlI+kK/+v6xhxSkl
o6S9GE59/fONIOlZp6eoT3iy/JNw28f1RvL9DvSwN0POsAJnV22dCjARjssZXqQm
2vkJSh9mIWNpV4KpPf28DbvJFEXKBiNvqt4kDrlYn3SOKaIWLsrLwFK5+fcTuTB/
r9qNNyOTNlfranasm+uc6gIE3AkCRl3xgYlcKBvF0WVTW0bZrcdaQixqhTZd0ASX
AEC6zQljmqakbqxSt3SqPT+L67YS+KEQFo/O/1uynUCGPldtCSgKDMT5jXc1sLwg
VWjObReMQNd1vZTphysjuVF0QDzhXLdo1wnLfCEbNHdfJKMEmljMsiJCKITtVXaF
Jxvzd05R78D+iB37Mblvx84YpcHQmoZ84ju8To4abJZ7Ow/ecpVT5+/6Oyr0uAi5
qK6CL1AebgC+FS3YjqjV5EAAZTGCOMyiIN6+EnQ1D3j5mEzx65OQYVBfPYBQvxOv
x3tRIKLcFOJ9D3u8TH6786oLg6IldQiWvaTZsQPwQjc/Y8ke3vfQHrbsCD0SXD8E
JopAPgTRCiB85ncwsmTN7ZUxIFc5fT4rv8WcC0vn4uuAjvVFoSQNhhQHYvmtBH5M
GNesw3bVSiCoUvE9pctlHNBtwHEv3QJzwAsWpyTFEI6BprQPR6BqOJA/U2C8UxqU
PnPPK3rqIwEIYQTUbjQZR2jEU95gK0ozInHdz1iFNOVJx0zviGN1fciqfDwOv9yI
Aopu7kLovJuucP/PXh7jUNMU/UKTdk86oJXvyFmr1fxkqzCJ4eApKq2jcqgvqNIN
pKr7WT5L36dUmJZZ8PZfsJ+d81ifCfYwVKAHQGi6KdfCpxm1Q8FgCZTGirIHLk2q
dTuQNv5TpuHaThmr6eGJYnU5EXyJS/51wNz27RuKESh58gR2MSEYXqRbsKUDVDzd
fo6/uwRKlFWFs0B2/WwV0QTeqJoCAn4M4z3WB8p+/boD0PzT4iQk43kJ1YKoOHmo
YjDjqfptxwSxIUrIK89hWoTpsRdwE+57hHDEKvcEblAcuHafKjV4Hy0EiXF5RkbQ
mEoiGcNtUqfWDH8EiP6N3aCsilK94j0+lmlcuDysaQZ8/6pJJ6cwBdCHlERVQLix
0N4tpgQLOedX8fyAAytLeXBIljm7ZXHzoQTWq6ymbKM5KXLL5NAwSNIwP0XPm3eZ
J/jCz4MqSqcMdPjeQJA25MRKa0COk83kIIzLmfvuiCZk5Snj1+d4jeJUSkno+9J8
2vsXATo8pjdrPVjsQ53zzhWuEPp25DC0wWp8LguqxZNH4+VrLZtsUvRK+MH9g4V8
7zohtljwKLhl8Z/lpnaJjmSWsJDHmHNs4xBsfpKf5Tglve/kdqskI7mLJRV6b8D1
IZrHK6bs0OQ3tmBXTCBtMYywm9ITYgr6VS/g9V7LbSFEOvwF2YtGpDKsE2cT3t45
pFoLcnrXotnjAoLGjCGJ+DSyVG5Y1JJeYgAy+qtF5cR2VLAfqaEeEfTRSqWy/qX8
bMr/rn0byfQqau0FKpQgBuayRRcu/m2mg7yfIlWbW2i07UsNlA0/mouGQGwz5nSC
70ENpVdiBsVy2WVd5tQNsVy6E5yqdItq+hWy4U7sepiQqdYYARIUucw4+TMMd2Ds
s+WvExg9AFlIkWsK5x5S8XACeNrIJoGdFgI6/u3s+p1IiR2vPcpEa9BNIqSTMSrX
I0ZKMpMu+QjDb8UUsUA1/e+0GaSBF2ICcmhJdT8cq+IiIYPmNO0VB5DQPAwa4+e+
Hhmh20CbtCXBDixQZJ0i8x30waqBmRXepcHXVwxpw5WzvRYWgb2AghEVbOq7Pp6n
KSwm5QE/tNytBYStgbZCR6oL1lT5NaYxpWwD5oU0NxBHpQp15o8f1Vn/CtfCPtgY
hdn2bxQvpTq+ZZ0Tti4QCUyGhRfPPhAt4aj85H1DyFCZNLWqYquPSpYJJvHK/gv6
ac8fgfJGTgoLHvACLRNEULBjKnDC2WTNbD7dToH9C1pBf0SNkBXODhkzGXmKeFdY
tbLtYCKZNsfQFVUVDbM7eYrKeGbnquQph6nK7/WIQK77HUOMBdAvuG7MVIIi3v0d
f6U4P4UfjvW1F8qOKA5Y3bpvKV7dZ+o5ioABHUO++Q7boJ3JOgnIhMi3O4HTGExg
jvspDZA7araNS04l23+gXHJi9bRbW1BK8BBtRvPktVEOnS1N/KvO2wmYFerGsopJ
eR/ko8h/l2jwgjuxADm1Nr4bFy/Yl1aXziHA6v8hbnzQnEDgG3jOfqeVGrunk/sC
81zHLBHWn/eOdg8Vpt4+AtBJ5tiLSm+7UYjqPNPLHJ4iCMTAvB8Sxr97pbHJRW8J
rAZSqA/4vXkk9XMIO7afvQWvq0vHeKHWM9BklfIyPVstNq25lWji8yCXXqJyunrr
xzy5d9ZbOOD5gWy2EFCYxqMcYmUdOLc+eZIqFq9dRjmQB80V83T/yNfg9Hbci+L9
ziLnrmB0ai8mC9Q9V1FsZiO/ENjystU0Kh8Kc+Vkxd3A1+POATl9i8u8zWfaJERH
Bypwuweesym2ntkN9HteBmmbPYZ4JmnUCMzj9dILGiIgZY94Oh6P3aCqobMqxUGQ
8LVoM3WWh5IaLOylae7y4VGU4Q1W9fZLguy7BEH7r9/10g70qevmHNOye7tgbIrW
3sWnxJqnDXAu047Bb8/d9zG6hSW/Sxk67uPFOsmvd0zdp/o2BClFdF2KbHRnr9uP
G/lxF81XrUWBn4gR3XOgBaYxHZK9cdzl4xl7M94NjERefCALZd86205PdBGfXuv5
gl3Kk0C0DfVMbTZUA2cnBQSqPLWSvvT7ZcfDoEBoojbk/LxflZajyhhX4pfrZRV8
ey6CKKa/on8uMThR1LR+o0pufdlm1wcxF0D3iaXuaeRN2kSRb4n2W/KMIbU108i7
KgVIuOs1X2XYPoHTTN0wBfDj/nm2xdIbygU+8PClciPAe6I88NwGl7CjCgQNQcYQ
mdUgyjrJvdDevAHvCoPpiB3eyUZi5ONFb5Bb3WVBSbqHOV4a8mZjEImXhIT8qHBK
XNnbt7csntnzaARm+Yn0crGFNA9n69Smkjl0VfbwCHMyml2JK7wEpbk16nOFVc/L
xu6t6cj8EWJuyfzlRCx5oqyHdL/IRDyLhbKIWA5oIk2/SCIKPLxhHtBS8mm9pq4t
MoU1M88g0CcizE0iXHaPpYKUbXj/wgnKh03aepdW6bSbehy73qwbaBFcBKVi8s0D
G/04okBbAsNM6/BY9Q4H8Nz7exZJfKUTJLHvx7Oq+TUKCF1ZO0+tThasKbgxUtin
wrnEh8VSLjxiuXEHYoXIMMhA2QCKRxX3PuoQDnsrjcH19hyIgqeQst1yE1RHbvc1
zuF1CbYpqU7ACjZZAgVmSDDSMBZ5mPYsYZ2sNmYHnuo/pDHuQFtiEEgxzzS/1Jcm
mzNolBGzxwB4aifUO3RZcLhvd3zIQOpL6LRnno2UURvlpHkOp1vA8bnJlzhVJMop
+dLzjdcCEwjRDqLWIuV1FAq7UYjcSx702UlN1rBWRv0U/L6WV+S85WigTDj5RnmK
p6BS1OO5pTGu+qc6u4SX/d/zY2k8kMD88j8sUh3/B7ZA6IcozBudmraCVCLsGQ14
LEqzzm5uYrKq5VLl6wOWKpdzY42UJyFvQ+VjyQtYIPGr1GcmPZkO8IP2ihtSqCM+
v+SSLY6BeVscV+VNUmQ2yz7vNOT2vZ0fLmmCpOh21Q//vVlnaa56WVdgVn/IaKZC
3uS9Kn3rhmt+m+983Vch/AA3UQe7PmFGlZlDjitbmhKAc4jcH7cW5otxDngfPNA4
dQUuIxAoFVRrlXoiZYzUPmpDADrFxfF5uutAPCYj4yKOFstUehPiWqBwYcXmZxOg
khtlWX8zwqdjvkf0hEN8hWSfAB8nzvwJWkgKHAneDBTAK+JpMvcAOWIG5zE6/pXE
M0p412LOiWM1UkWDCJA2qNOhTlXv0xGb+tMkxPsdcxsKPfmtwsStbCdcM/NUbf7s
IQrw3cN367F0IIYttjyL0nRHvkg7qSuwJoGbWT0pZnovj4shGYYhlEQqpC2BAy4Q
ETyFHTJX9XV2L2hdOET+SqPks183/8y87d7kyDIuOWPlKRwOENHO5XIO9oVtUgn6
qmlPa4j5dq+0i0nHes7IpcfWmDvjMRqZacAOmH2a5J/5Hv/4xwcz6HRTXx25qSQX
TgBUdaBLcGoxgTNqZ/t1+2OiEYe8mfFPMGe5VStU+8zDb4duajGA3QSuz20EAfxH
oPnG0zPOs+z/EVru2xhXZ449yjQgu0v7/dym/WI351R40oLY/pphuTE3KJ5j+8Aj
4i0r6b0dgVQmG8MAz8lkH5Vkb4JVbCg9iizp+7C838iz3O8JUYTYG7gUiiSG63+p
IntJAwZC3lgTfxo2sj8Pv2jFtW8UF+YamhBIo6DQOMnSc4+QjoGGAkHKJ8DzSzhX
wjLNMHb8JYYMEQAY7u9VhLXNwW3I8a/rU89ke48dV+GPCm9bxGiY3h5li5C2v+az
Owb0sF8OjkjstTveQdK1UZVmihKTnXRMsaCygVpB/gh5SpMclUq06o2tjbPW6ZyT
ePbaJrTYuuQFtTOleFOqw2anP19jZYEAwRGUeapWTXiei2BKS04G97g3KtIboMIo
NiX7UflZyXB7xAGUHgF04wf9GL2sYNMR5I1ggFff0XR/pXRMgLK6Cay0LWjxZ1QG
dcjZKxcBBJUN/4hf2sadG8ZPyyU8Ykx9Cn+ChPCQp16CvaHKXOzgCN7cEpinwSj+
fQcuVFjSZD+QPLWxjLsFYVRCFhNNDW4IYZ3gaMjzURXxapaoDSWCQpeBcEpSSNBY
780y98OjWly0TfMN3wHPca6U8Dhn3I3lzjdnbnO/aCz/oOIdcFrwzGCNm7ntke/3
nWToucKMjchcFjxPpRJJTvuP/q0VBD0qjACZi5WoFCgkyUvNrGxosahJmmY+yjKx
aEM70R1j5n/FR1wfgGFRFiR1PH6RRvex5pFBYDp4ArGOb2240rlIFUpDxVvqgs8p
WUgeUSZCUTU26CYe4I62AABry0302L6I3QmGt5ONdOr+EuZaGWQ7q3IJUv7F9sPN
rixUQyO9auYezzBrBsWYqUJRTAXWQ4uK5Dv4pK9HhGE/pCEHgqp3r2EgoufSCHOq
3taPFkSktxXBIv+ptpBFpMLIEJsvIuwOB6jdYosfZ65YG0l9BkyHZI+V++CK2PXd
/qv4BfRWOco0sSdRFk39iAdOLAm5gH2UrDi2ngqxA3eXIXG7kHokzVJ2IgmK1+6k
/A2s5+rP4p3p6w3hJ6M4vqoTH867JNVXL1vkVrf3Q04Et6iDGNgEJbHjsXTECgMd
M1PX7Q4AF5/ygtFWoL3PTDFFchXDgUxmrHhY6ZvGtt8Dh9v02hY6f6bB8HRMZ/xc
boZDVTFK1etIZmuHYa8T/zz/ZuM/o49DW3ZOr4ekmnN4HyFVNq63DbYOFCe24oY3
FKsogYkLZsNcra7r8mxRCoLv+irVEPv9+fUHWVxnmVk1Xvey9XB8wF1yT1pYaRhR
GxwU3gsvGcUBB+aHfJvGos/Rou++hhaFQr4MTdrMbUWeXESIdb/8THwXDDzpxmFS
CSUzKOhESmhyeXJy+ySMiCuw1XdUyGgGEdxj7IJTG7FhraB5lH6JvcBMwM0ppFSt
M4OzJedbIT7PAfClLYQwMEGNm7+rc3I/53js1rg4QZ/YpiELtoYgsCxirp5AN3h1
Qzg0KglrgxZLEGPd6iyOzldNgv1UHdOPX7NWFvWikfE/rBsqjYuyszGpJnKiBDZ2
hVCdHQ7H4tP16TlnvtRuXvc3xS4jllkMn2PUk3z9uPMbmWNwYlpDJYYvblPkrCSp
InfYo6hvJ4IPsZbbN3Ap3XAF0rIF0VOeK9ah85TRzDSeAiPooMt4+2ofFHtmZtHZ
A1mx6ibQ4KD42ASR+Vy+YlZidzz6HeVVG5Q+dXyfwXZyxUb+yxRlI9S9GqvPGOR8
HoBB3Fmm5mJaok4w0Plzx+M+iNaP0dwK4183/YFZUYgQKs4PkTTD5/Xaaen87MDJ
5hgMa+ee3EenFsiHnGTYOY4Rlfwursm3qjdaz5RFUltLvqmuzwFzHaOf3bQ8/2yj
yN7OHUKiUZu013ttOLQkJVxJqjZ8eMNNbKzEQDRZgb771ntWUjAz3SLReOGZnamS
R2H/ozupF2Lq1AZdcvtgfegJ+hcYs0QNJvz2mi66tPK8gFC/ER9S9kkHAMdHBG2W
ROjpdDiLIsbjj3oMUuN9Hxmbx7D3mt28D6P7rM0q2VW+XSXUn2Cx/dVl8S+hbkzs
9Zl/MHFNM535tD65G0n5Cq5zB7cdz1MT7wJT+FNGjXipw25CGAl+2jhvEx9r6rRh
hRJNPgk6hbyh5AVOpgidAPNNvPO1RgyyVLRPwzRDax1Hchmu+wseMJpa5sjbtElR
whJ/y95h3cb+jzRc7eYbKW9yG98yKQ+Vx4qQ/eD39VOdaE1Pff59JgFvewiEuDYp
rdWmnTHaOdcxvEOGtjZV1CgLgQjZ59Q1aPPYjT9zDWdiHWOKB7cu0edcvf25zdSF
LUzMPaYvgsUP4gE+5CFIuWu9j/or5IlW4qqURXWjYlHXG99RL5H3Y7lHX3MmnAKX
rWseoKUJt0u7DmNxtaeKHMJdkj+Hv6XZI3h2JZ7M/BqztLgHGazgcauN91xZDPHM
tCaa+FqynF5ffdbi5b/EJsTDzynlR1TKWglJlMCRAe/+AI+HcCYoq421qDnHiZmO
haRTuhf4Qs7ITw/Bm6tXLGacCFMrVQJiSKRiq322JtEuYAgUyLS1Rr2G1eJnnIUk
+46sqZqiQGJuvgk2M7QzLDDXSxJyJVGERptTxhtJvjqAsSMkgi37YTwK4d7exHOb
GYNp2qcBYqWHr3JMls06L9DcF4COKvvHy5yYWyhrVB/lVU9JXphq3sIlLQWz4KU/
R7YAZgb2UKeysa90jm6TRD48zP0Y/VYi5TwbvQMY64elwIn7LL5ZljGXZ2keaRog
23s4W/7yE3R9H0CX0F8qMLqU7R7zew22vKu15rNMsh+xNsfc4h/A0ht9axhf3vqC
xU6pQvTru6JJI64M5JibTjq6wFse5jig/B9rTvxbAW97ODf3qzO7c5OETEpdtrt1
BiwACCFhTHFSCQ1Owb2GZQG9vlMgKrl3hkKy0WahAlnn4wLBUQPRBPqd7XX0gfa9
BRSSeFS2O7qcY03Z9z1hW+Zzyqlko6ljWGFLxeXS5GpBqmzevdja+1g/Mw37aw9Z
Y0MdpLEsSqbgctLDhLm2ds+KvveQIBjoQE3XMP+14MJgM48GQmQ4gR0FWMVlpEsP
0nw3zxko4HXsBdYhjssj0W6iGTyElIQQw5TJKbBlnYW7zmqnmPvC3o4aBe4z+PcF
dKjOUvNz3MeUM9cn17NaALrrUs0LlYlsP53sms4tooHAPL81UxQpsMlDeQUvlnhq
RYdhbrx1eTm+x0Ecw/BH1RKNHXOQVFFV2lXLREbPewdUNzkqIcgDPZlHdwtBvSWf
+girjthOw5HiVHCBNKVLMO9wCRAtDBdEp+4hrdgyeQYgZdAlvw64ZzVmI5M57gw4
qxo+IOwEjNNPwJBoNWFxu3JRE3C9PW1HcDqbPWW5o1wOzLil4JJ7inPNJ8YIZUXT
atnwOdi2IeoHXaqi/bnI0ZfDg7N9oHzJlFzstKkhEbboderKi8zZZTyG9stpnU2I
OrJm+KEFlJFvzUl645z0a4+eniU2kZDWVWUOrCbEtqmQUq3Y/wm58oElJyUvY0KF
ggdqyEV4faEp3KDEDeamKY6C8C50cXGraYWJH4rW8zDa2hoFYDv4FAPgZAHKgppg
3gO/U6yv6Fko1bDnwzRbnTIxmaHNqCuGllZwCDJzz95qW6KGce1RzkZ0RRuWN/+n
Isvcwq86kKrf9LbGVRzVgjaY23oTu2F0GWthrrz9AdPmt78dXR5DIxftKKVrc7cj
a3qKPVb6OrO80CNjhR4hiUw6i+sa0AdUlvCtiCHXPd1c91NGhYLJWwwF/qxK9H4/
brVOPTk+NwrJflBw56l9U6MZtffaGkycOqdaSSWrvShHqr9M/kH0c7wlZsIEIIBZ
uxjW3iaVd5AxRpTnfxPKu6IQx9HxtWrZ3EHTHRXnGiQQuX/TMb3hffGrN/FbZOYK
usDBTWyS8RpoYm76i7dsumi+jN74WCjLbgPMEfRYAgNjtF0Fyk8E5ncbM9Y07KV8
B8QbiJ2ehjtQFxgWZO70C3hE+ZABMNNqzn+QFm3hhsuVd8ltcWVZsb0U3Qn9p4UH
/c2xya247CQg6rMBEFdUTDtjjxs+w89Fps040x+iiZemputhxgo+DibjGj8aBqUe
YT8Zr1XFKn6sxtGXsq7nWmVBVdvgs84H49rFIgDWNrahj+rnGWfABC/WTOfcKkxI
/XG53TT8c7V6irMZqLieBPX/XIlg+QKGyVX7MleiS/5Y6A8eswTR3aBw/xBQzDP8
zQNwfGnq7zIDAYXY3wLpuyd9u6MG2ZWIooN+r9u5krKyD0EO7K5ziPKcI+Z0eHu/
ytXEpXC8MoEOFHZ1BhCEwhYt8IcESZrbIq0E1rB0q/CeX9jWzLSVju7w03ivQX4i
uXy8dwDgbKUKNtyk/cKOaFn+30Gy2J8vyNRPchb7g0cPeJipunb8iPPVv9QdEPBW
y/lWShop9VUACfY+kT+n6/CRliOH4SA3UrN8op8hJuWc3w0mILCaOIbK0IWaa0c5
Eiybngs1O6L35p4mV3Ji6I4O1i++U7h+oU/XJDReyaYpK6x6/ThHGOV8tdO4qOTy
79Pv1wfWwcOW4guwg9O3ec38+ZQZiydIWo5Ddbkb2zVm+2pvLY1eslTwJeM8coXH
ElpAiqsXXLQHxFPMMTmrz8CQJ3Gs1sCquwbPri1ey/V/6QjYCFbsWeZVpXq7mvqP
iXJW3nC5acWNI1thSjuv/weEL9nivDInTWIf21MYcb4udtMBfdHjvhVU5tqH+KYG
u1daLipPnOODyih5EwTYussD5z1OGHhVVN6u6GVJOxmDgPV6MaWTWQci6tDJJ4kf
KI2RB6WSeIHu7SjtXJrWQ7eBCB+NXrhRbOMZdHd/jfWVVNAiEqBS9X6W38vSYkmo
Zqmt5zPxchlWEQ6bL0KcvKoxlFBFFah06XYJgbqQOI1TXolJ3QblwpbKjYm2ht71
bnt3I0CrsSL30mFxIBnl7trbBVZi5EdT1vbnPgx46d1UUoOy/sJ1s+DpkpJ/ILjX
y+hshJixA8I8VX9pES2b3RtCcSQlISmevV6uA83o+v1ncYI5rWOBMFc8HoNphD/K
kNm5tEd+k5NnOg3YUy+FcshXL4vWkZfNdlpfn9yuOfdjsHA4AXtvBi0a0rgVMAUk
pSpjplnxYgKY8/zN3GafsF3yR5Agn7TBCXc+KLHs14b84I5uB2zPHzg8pOlCAs8R
09P2H6c1DY3P3+24WjXZSWJeEkAhMOBlkVE+fNhruQVXCmzZ1IO668ir5IgzgPhP
aRxPZy1WqT+EaWXS7/etSJCByboihYXEL6+rBrJWyDEOuIm0JN7JePuMSZW1V8fS
vVK0C94FozuxZ0WQzIzbkEN6vZG6btg73jGvd16txPIm8ChhCazTf/wO0jRgYQ1G
iizEWASvqMX6ddyVpgClnjAsNIpP6lUfgfKmHER7WuBi6uJkyhBkuPbjuDttSa4Z
AIBC9gjPc0XrY8FP6L2UquRIbjF08503XuFPT5psZRAsdAM4L3FSm6+OtPWF+T0n
4LChb+HVmfuJ2lZdBxNu8hpKbx4gGr3pAzuqRz/QIvaP/5E3toS3KQM9dBn+uV5h
qyVjhyXZHWh/4gW44GkUqz2HEQzuaHCCyR7OjKgIiTzVh13us0+HrqI4D4hdDvkR
mW/i4PYuMTe1TYARoLsihfKf1L6pS36RiyaHXJ6jlUD85rkmLKJfmPzL7fEfNLPz
oVGgdfW+svFporkJ+rPvTGcVI8y0jGw2jvDAAsspryzDYtPPzORFhoTalxQcwLFl
ZO7QyzesQrZ8M9uHB1qfCO4DUtXnJEO2N4YLLl1p+q6nfLAvKEvTPELyqwTR8v4c
IZ0hcuaysCtzpJK1iz1L2gI8TpxypG3JqZq2IP5QkjN0ZejnPNpLUD1M61pC6eJM
+JsMnXUEFebT6neZQP2nPcNNGSfe6VccvDDwPt/rzeFHCPfn4mJ+fvoqxKfW/ma7
auJ98wvIYXc4RAtjJ/vNC3a2O8AiNHfXmVFmYvyWHiThnQz2V1zW1DmWvHV+Kcks
vdjv9dHMkx51rr2Z37k28EZ6vwLSKsRox6t14hhju9ceAHZLpH3aXYEab6Sd3q8q
bmvE6PV9YlG6GxF1Pkc3l6Y80x2E112453+0tS9XBuSxaO5W7D4cwnbwTPvkQnbB
suezMW7q3HqJ1K06cojXeQWFnnCxHiAvewN/hRNM6gNqgpnJBz6d0gpBJkF0aYJy
PjHNgCOY79rEZwHNcwzh3x50dFsueCAmsHhfGas37RgIRzFZgvbOC7boRb15kx/c
Uz1cLZjDY1VprvgGe3xuxWzQ6UKYiuBNLqY9lx3ILc4akyp3g8fBO4/Fjsq8VTqv
nbrnZWWODiJni1CGKBU59NHoQ4w3TdHvIRZEuSCIEQEh6MgqQOKwCmomJKKpLxrz
e2rV4W6ihzIdJg+wooL0qls8BtUOQz+sYIO+sZQxw1QR3u1ckWJfiC/9Eq91IZv+
dCFlJw01DP7YAMB3BWgIW1ov5PLaDiDS3tDpFEU6QlGJzwEApwXHf0lfPa+QI5iZ
RAC5vU5JTu5A/fID9JxYlds+meexBAcDDlO741j27SlGXm5d/Ej2duj/77RUlE1s
8L0q/k7glBJNJ4kp2dWju2EERfS+VOOV1T/wnheYOGOpX4nkdrZhzqFm9M6YWQtd
d+PyXj3tsgul2qdH3QdSnISSDzQ7I9UBhXLkpHlRqCEUp6TZ+vagL0eXllv74s4o
3wAPRLFMhc06oRWrhcOs7uaW6BMlu3Obhl0PFUiSRv0RZqRezjx4h/iRBa1k35vQ
xZDU8YlqWtlsyS1absoZiYpYg34EFaGzlgTYE38zz522h1YcOC4R6QCEzp7IdSdB
j3cew8L5ZDe+rv7AzxEQ8qxC1vnRB1oZwRDOwR+Ps34fpR/OoRmlo/EsdGxuVyRr
YFoI4ui3vRfjU5uTusER8HspYI8mKjhk/bf64WUPxAibjJwMksOKTHQDYrBBkmMD
6x6bEWXThjy6Tl4vWE/84jCkqdScAUCykCKR07VqA4VoC6WTSZIQGCLzXAJFrTn0
Ol179xDqC4TjW0F8OQcB2FkRFqRUhJqqSya8qvH9yaq61k9ogsgREgQqVNqMwt5/
lT3iBGTfsYd7ejqtqbKW8LvtmSWtJT9xXJ0ld72KW2tP6P4sbolu5/73ZtKfhFV3
y8w16R7+JzbF0UdN6IVFd83H0/pFWMcojYAN16FJpxBfrQ46Kp7fiYW40VK7kp4B
I7zB6kvKy6XSsoAcjr/mD0iwlja73Zgsi8D1LNOJ3v6VyvZJCrqRypiVSK3L/+iZ
Uvtn6lSXIlrfw6VPVXaGKHBICxL4Yp3T7mDxynXqQBuZzGF3sq2dqbUCmEGCe7lW
frdnq0Ce98IszcphrY9IM53TzwMMRBeU88ukJ/Jbk3gT6iCEDt1CxHcnRWjqzdYH
9z+Cum9FL5FPx1Rmk1WZ4Em00K9M/vrSKB7MP4yq5bKrxYzmstyk0oaltZG/74rC
oNB53ewWMWJ6tUhJ42vGSRY0nQ7mFyhQEaaAlOXos4lsb2k66yVNGyzE/f82eTRu
Wkov3j6nSTTK4Wt4O+RvhQgL3Rk2U+cqZWCfs0gzJ50vEawbF3QxiMnUIDYmzQMU
2+SKSwWtGsJqdSVMdr7fXJxQIc0p8RYKCEi7pYoDA5uNwTDbTtxGcJydv1e9S6CZ
4gn1reeEg1VZ2uUx9/MamxGmGmhapc8iunuk2Tgd4obrqXS3TDIfQvYpmAMsDqSo
TzC+WL2fhV6iuKr5E0Y7+L3voLkbczCt1hJYPqSqMqSp9E1U1pPoz4wVxFVJeFhZ
/DYwewjjQyxAT/Br3bJ6TPM7DWry1QpZPLmhKScYGL5hG3CIzR0+eFCOveXJ1nTn
J3lAoJSWynkeg3Dzpdf2mRAr1niFyOcF1599DsigztpU9tUGxdCRMfihuqz4Af16
puQWg75uZQv9fBkvqlGpfFiaa7KWfjDckrzTBuQesCDXBbhADTbJav378QEl3PgW
kHPLvS1tyAUm3yexdZxChBaFmDpaQFc2ZeZ/r+lRplY8WtWtdvuqBS3KPTwhpM4v
KlJRoBnm2hXOpCqFbMBrDZtewC/TAAYlLnmGbVLKmW4MzfgMqwcp+hNhbDBgDv94
+yOVEsxuTb59nZBb0yLHvR9v2Z3fbE5tQc+ivknCkqSDNw/JagxC06DuCBj3dNlC
BmzkXlnTySXtUym5kwn3e1B07r+OfSceq4ghks8bbjOvkb6p02KNFk3E4SizFzxU
vXhq1k5pw4aPYtVFJdnw0bWIo+5/+LPozx8S/r/aGPDrKQbHlfPVS+rYGVRxgkcn
DtT+0V0/pWuKCyspCZQgTLZ2VTfWUR8Vm0kCF8SVkOsYAbmjjScO1vxex3dHvZ51
X1A2+twqXsYQmkJ8u4DZAGIwrvJBw0odP6GjLq0iG5HcUys29c7tJLn+mze8TKTZ
FJ0k3WqWy1h5beZcDq8biKBpZALu+Nd3rx1OlJ4BTQkwqLsq7wQO0NkUsvQ15+uV
xBuaHXYl3CT2b/ntejZayvuYMeOYfYswJDefEzCYXFleH+WA6RQhjRclzvfejhPf
QbDO0FfE4O+0VKPw+rSvpQSe2+hiH9vIP2SeVwPao1xBeedy/Vg3KrZB2iHjMkeo
zBQTdbDMyn1DeLqoElqxFlXMDQrTdhNypmDxvtrmK7Rsi0wV2ikea0Fd9g4j4gmD
CW+gClsgwN6sj4jE1wFYEm2RL0QS9644DZBHdXJBVUqJ6BQL79XiJnVFcdYEOX6M
InQzrielvULvUVTy2vBZYhIRSy4J5pCPf9rgQRDyVp5aKjXZek0xtB5uK+a+Dq5N
GZj3Zd1QUw98EBaXvYEVWrSwUhhCjp1cegvmrwc43OsgvsoulSa7qWgYLH2d/AZ/
Wa+wuSizvsisT475bspJiLrY1wvYuH5Jmn1RX/X2QOJT4UmCy+1VUQJuJqgXQD0Z
4Kgqdpp2tT3Z0PB6m/25vCaPrGTYEzRdwC0+oTZlA6/2nMMFmAcXmDdw9ytqWrn2
UBqEZy2Zsjz5w85L+XXtZVOeGzFPIvVn9ZSqTO+1fwZ52COOzDJiyC3foTkChdq3
TAN9j9vhFc4IYaoU4e0B2nciN0ulzYAgHl08T7CBgdJ7br00/T1SgGvaSWmhGelz
Y8WxAcjMvVCJzBrAYrkHB5NWm+ghjSTsKseg1jo4Op/oW6OHhHZeeqJu3F1Aa7qh
7QNIrqJfpyTL499qRzuxf156+wyNv/d9+Pk/Obj1OYREr8iScNxbhe++tpSDo2nd
whLbZdvGxksIu/EkbEQF2u0K1Pi2WANQjc3IpVoNGUKiQViJMZ7IpRsh6czwZtfh
viIpSUx+Vd3cogCP1Fld6hC97fr8Y2qfY9nMdJf34HtiOC3psfGbIPOmreU78R5q
rhin2SKi4uN5iy56btwpvOFCHYtZBsgTPXQjqktnvca59qIee2213siizRosy+5k
QXNaef0EROFxNEaqT5T0cgdjAY5oWrUBi5RjgZDb+8BOXCtd9HgtvOsb8eSmOiCT
cv0W7uJreCfk2h0p7o50QSzRtrZYM7FsX3BuJrRzKRWvVPwhrA1J74X8lF4aZv4p
jEuIiRNs8mkv9o/d+M7hOsNz0JJYGgdY0BzWOdLfDUz8O8veXWZGsqDzWGa5wX5E
8cozE5Gyio46XYDsAB5nB54I6hQ01HEMOY9P/3LQdRE8bDmJOBT/NCSln8njhMRs
uvP/EiVA8I2MDoYFjwt+pRM6I+JhOCT5W0y8OvJDC5qY56vh7I2aHFovFY3CsYGR
x6l+NLdOHrZDk5L2EjBvqHKhUIFIhnbCdjJBtPxRU6Y7mfaku/2OqyjFFNWqllIp
BvgN3M46s+Eh+NRwU71rKsAc3+Gv/Sc76A/GhqQSq8fhUODtCvJkFww4zuuGyAW/
zK7oqlTMxz4VkkejxCa7/5FKFLFjUxLabNsqv7yl1gkUR0PE51K98Yaf5vlrYp/n
oQWyJHxir0lqnzD4PTycdIWMlgwUaKcfrSPlckJEE0duEBnuhjb5jpCwysWz6/3h
u3t3rIpNpjMPn/AxHnhqsNxG0Lj9ndi/srgSyj+1tlSQW+p1g/fvlxWVqpqGyzCB
LacyhUwjUJM5eVBe11nXf2BnU+pJ1uZ/P4VshtD19zhLHKyj7Eaq+toO6FVvWdl2
fpySc3CJD0ZeIA+awEBG9dgXuv3wNDwjHZVIaeSUyz+nSukSiwEuhG5WzjbO8+iw
TMldRGc3QYe9/aD7KBDWspQX9lFc6eEdda56hC8/kn0NUbGMLCNzwLfc530RsJAh
Tki1thJ84vl8UHh9GgsIMQ17r++rziOw+Zr33qyOU7exiiSRup1f3Ap/Cvsu/jX3
ZDb2g0t3p5LEfXMLjl1HqsSnOgITchNed7wWegOGyHA3rf/lVIoDxBT6uKFZhIM1
81urF/frWQD+u/tyYooXOlHbXXgJnODesg6hvmmz10+WvZjb1N+9xUtzrJs1n2F0
70SF8wyQ0aJL/4xTQ42YSf3jSBOG2O5GspOrbIgLPaHQhxLJm6FcQflcBSI9dAp5
zuxJSV6e5TXfKFrvR2crponyjiL1L3pJkc6L/hsOPma4j0HuDheWk8VLch4oUxeQ
gV+apl31w8LfW0hMZHQcjbbCAJY9ts1P+O3W7+Cwz58fnucedH6axdgYJebaNltb
OOYi8bYcRkT6oVDI/RkZuvoX5ipUBUUg90GhDkTN/xAtkY/Jh4BEBH3TM0g9nKex
aH1xPbF9rqBIJiC+3YwOWWt9bUFeySeFd8z+phHY9M4arqwUVpr1uEjJHyvS45CG
GbpDNBiZeUgUAJ/Ol7hbQADSdAw5nEGV0Tdgxg/DdcuURpsHQIYYSm9J8jrhbfUt
AD6Cetep8Jyr7PpP1dRrpfyFA+/ewTT7LX+x1B+PpjoxNrc3yMUbpum9VQ2h5om3
mfIdYkV5WgrvKu72vMeN026riTHlE1mOGVah+FbEkSMk4xoGo6aP/mLJQPFwOCtQ
6bVj/6IWe6MwkJSDzVlcl7r2CrUKaYtg0WTd0C8rqWdwsj+3HN9rEKD78Oh66Wym
yjopPWomJXyfyhScJ+Qwc2LKgYsIUOE1qTCstgbAR49f+4iSLqJGggr/OIggd6uJ
exgIkuMkUSJyTeZ0TTqVVVvGSoplEqsciE/gdmERP3pMnLY44e87Y0WveR9cbc83
Ep83Z+AxQa+S2Npx2Pw5jlDpmwmYjMu+YvT1YgkrQwUYtJsHZQgBGx9zF3KgxmKl
8MpAT+zkVWFfyqoQ/DMxbbbMRKidMcMbPTKiLDsxbfiGNZ0SnUDdTWGsnFDELcIf
w40Ym8JrqzpVXNca3R5qrha7dLaoBn+GMKrb7o+Rmmo1EgFNCxH+zD5fSjlw9xzE
wx04RQGK+CWLD0V/y3QODjmeTAkJv1NWf8x9f2B3tSHkkAvH+NHW9wsvlNqk35kg
BbtN01ci+5zQL3FWuAPwWCde6iexPLBtlCgCuZJlJVC+Y4EZZcqdEBEAHrNfXwNF
cCmE7Ep47P5j4wfkRSJ6ewLw0FpWftOmD6bvhLut58sty+BZMNZrhIjrLPtfMDm4
67FixE/CQ8PBYooSpcZ9FehIn7KrOxet7zTi70xnd8g2M04A2P1zjU6CqMf3qioM
u9ssg4I3t/Fhdckn67WQq2gSn5gyN09Mx/JF7/LxzeGdtSWR/kex+vNH1RnDZYhH
a5A3E4pcELZnWyQtnSzOAHP3n2GjgeC+jIfdRqVcLRSnFobrRGABWeLwoCwhsq1L
hFtzTx3vc/dFVs+Gf/Q6U98RFMSa/0vkudX6OUuM74A+pW6O9aaC1H5opA0Kg4nS
b+xqrBR0gpVoCtnLK2SX2iamQidJuMlZQo7b86mUSHW2hpJcPRvH0M3kN+aR2oVD
amZ8q3MG+anip0smDu3jLDddnZCttWhjcfME5K13G0W4hjZ0npo7wNVWBlJFCn84
xkt5AEHJ6CO1A2TflujbvozwXl2f/ZaSrEot/TwG7ZexksTiOP87OT4s+1S7dJCU
22/HweyGSuyJwATtn/BBOiuJSL4DyXFg0dF+7q4mwkpYZ7LJSWzIKxE0rTvEaB2P
dcYhDVE7ywbftLhzDe3m0bmSn00U4zeQT5ZORZof6Tde789PityCW/NmVPqbO2Qs
pg7/M+JW4k8SwgXsHjSyRNCP9YS5E92GJ8oHiAB3XmHJoLNGlCfQhUIp0xPa/w6N
BXoh72LpjI1qElh+ppKB/xbj2kSPpmFSveKM8yUJN6Ydi3o4uaGgqV9WiozMxHGV
a8jR6ove4TzUHQVVdjFnG0/xi2XsQ1QAvKC7nYHwgERYIUCsRinVFahCgtCxjLkO
xHdAlDOIMhKo3HLdil2DKf678W9YBj65xUK8iZNlbKoKtoxlmHgXmobWfU9JUcNV
3k4kxCmAStauh1TI5wrLmBPKPgbPC7nY/pEMX6P4mQiLqTVndqsVXL60qBMNxjPN
H8sOgpDWjxtpKg0R4NZNSKaACGgz2hujuvZp3VodYc42or81m5bXx4X6kyIIJ9xw
QQhK/PGFDGhiVIQgoJYDfsU/80oeHhiIQs8fqC/k3JidPzbIDddCmAB0oX4FAb2b
Lgw1jD/pj2tWCqk9Pg/bKeZ9undrO+xNM3LaI6kBOpOfc58crMW5G4SQNbvfKHxt
SvMKEKNzi7F31p5XGvmJ4Dc9Dtb63Akqbpd/+ysGpTbp5vw+rv1dKRdqlwyZpc0R
0IAgOToWIL0vUQJaq/x+xbhlq+ckeIqyrIuyWgH62elIfcQsU1nxbMHQveV7D0xe
aH5td+7TzS5lm+GzAeO2g7QYa8SHKNdMw2VeFqr4lm0cxBSWUDf+VB6b+vzVG56X
Dq39Fj1a8/cmLC2HM8uGFWm3wVVQGo+tODwaXIu/RofO9DfmSGPW2YSKVwWAmjyY
B7a1ROx8I0Q1if/qt4nuZUDMIkbthJoKS3V+wp06WureiHyhLpMWBDQ9W433jCB8
DoEj8Q8hKxChYq+/fcs/IDBL4KViLaHZ/xu+9dG3siqIl3nLsbfuydYUtWE/tMS+
dGYbux2Q7Kg4U7AKsTNcklAlruFR/uL7ylTGUmyxrDTVTncIEwtUf3dEktidoVGV
QSE9CYx4DfmcEagv7NyWI2JWb2iIafctudpAIT64XfamyldigiJtBP4whONVaQV3
dizzZY1odbsrUeCO7S4G3yviU96Mf4tzzTza5YQ/p2jvQQA7sTisvrvvq5K2XmUE
kTK+hzUElOy4KoKjqDKL+NoNuONL+jbL9kLgqtAYomjVK44g0QDkOZjLShasK+nt
HtNF4JvtKhRn4sP+A+PqUHi5RbO1ICgYt3EajuGTjjKujmvheUMFWWXMhNYQRtmV
lC/KFoyKli3Aca/fAsS6xgTNRbfXk7l4TXtidxjcELwAFkUzIydYRxNbMRalFshR
EhwdpW9w6CNhA/wjgeV50xdLy4w41jLySdmYYPGImU5ngBDWsi8TaFZhY082S7+7
R6jig+jWQKSrAirviMi4X54HKh0gQgoSd2ZOmmr1TOqoWHG5N4eBN6AYmeO6y59n
nH4LCueGVJtLOF3Z1rJXu1tvube4RO6+kXYzT/DHhev47ipVEkNrhSDUsp+vT4Nf
E2T5VLSiICNnzfi+rFx5FnNhGfIw8u5ezDPJrqsQpSGQHoDbS68FCrPD57vRPHv3
563Oiq2hI+0xTC4DCkCTrpa2Pv+YUzFIA5YZzLrBuweMsni8+h0UBvexQzhuCnhg
+dk8nC4GVDCRHGjOgjUjzNdKXV3x6s/FAxrCbMFxULBMVGuCuU4Y3BrvItmRuDoJ
oM0izQpC/svQsUp1E3W4GeRnUzvQzRQGKXMNsZqtOLk+brIThVJbuoXeD3xNwYOy
xVEDqOK5BeOhbPyrFvelPPy2Byx45NXLTm34Jn81vz6As0CrF9dUwxc6AoizrizQ
zytuTe57gxvGgtO7QQ1WkcI/ehYGJeS5Uz22Y9shLadIfJqE7GnWZUAYQTstf6Og
6ZbhC5jrEOhmtMUNfs+BgjkZSc6DMFDMidnTsFUaW2w+GDpjEstSJhUBC43Mi7AZ
pCtG2Z63c8Q2WhSRLMC/EeUdvg052VGby4IykY7JgPcVCnPwZOAi3dvHJUytmK3f
oLROcrOXXCdqzpFDVbOvwsOxVd0TmkUuYzHvTwF21Co9IalmcCQDvOzNAwOT2Qht
AnrQ0GTylk0Gcg5ZyFD1e0coSPQm/4yhFQQT/Xq11UN7EewJRDoZthkVQpF6KMQr
ysxqTvkk5cGL5kgLoSxYmb3gKwnr2xmEx2WzIbT9L+R3pOMZhyTRADnht8b54xoV
Rl+59Nriyq69L9ToNHnZ7g6LQM70t0RLpNhd/3dOzMWfJQM51LvaNKTsKS7gC5hQ
jvGfnTa0lkVCuL5n6Gd97UNe8pMqzlu61NCQHcYJSOEiJfwm0wlQiwhAPhe/h3Tu
MFr+BdplFRX9R5OY1xstpDaRms99JZDdQ0tHcUD+l4Xt+Z9rjFZ/VSLR12RD3c2B
gYWgY4e9hpQOpLOcofShN5z3faz8KorOrdKwz5aleLtLVt8HM1BmYiIwdjQhm15W
PI6bn6J6m5VhZjUPNHf6JuFjWd6Xhrrz6dpV21coEMls5WShftbJ96UmV4C9gl20
WgaMYcUCjb+FIeDW1dSwaRTF4RjA4VH00sKA023Cp8C+bQ18b5QQ6+lR9o5bosnJ
hqE1fXOIprTai7XMC3vcbbPHesjiVlxzMvswctld3d8S5sjkCLrnIyOPF3Y+pHbN
Ko1OdYfNnzsNuAo3pmwHVj54XlN3Cd4j64UeujdocOzZ5xgZ2/XN6o0RyVHosSlT
0K+HAThZxH3qZg/QoVbsEgwew7vsWN2OIG1ajKxFP7uN2XZfCEtQ9VPF0iDfj57F
XosNYGcZ7TcS5kYo+yYYDqee2lydTzLvm3BsU6qR6f6A2SKeNedEs/TtcboZsZ1h
KHTs4CRxyHBZDgSURbI4oiqovi7l63Bqj4Nz/bfyBjsPfCLgCCZfJLrhTZF4Mu63
OxZzhkvRfAVPRDk4HQn1YDxTy9dwm9BLNCGWsXAl4iTJ7RGn5A4K3qTwnSykRAKe
SwSw2rdYOvrBc26C4x78SlpTCl/5EFIqrb7apCWakvJyb8mkxeF/jIOaj8jI2emG
nVyvYnFLQdPLF0YWrfQDbapZKbkzuaLcp5ZhaG/mtLryOm1IhjT0mqy+TiAi6IG7
BoXUzmXuvMUMo0wyXAXmZcQLQ4Rh3ueRMY/4xuGQyHBA/uXDaYIHBvC1IZv6y5XG
4+UHO43XlPTeUZHhnBvmaTc+dd+FmEvMV05diox+oFBEyiL0hadZVqQR8q2dz6tB
SUQ7RkZmnxAUVML6I3/qT6tj16GD65fNw1Ioz/2RUrni2Yhr68c2yFb10vsXvYqh
5L5gQwLgxoSdDylRNWtkbVWJNjDHgCqU5jviuY/Ic0hdFOzmelWL1Qz3Q88EqQ+y
EUFdPgsjsLWNDEna3278MsTLhoUJ8Gv7p2jQYj7dIssyse4JjFKx9/hgSGaAJIzr
T9Y1iG/6fses5NoDAY+YCfv7icxWqtDrQ0ASLQw5GgVpGdB3z0pRlF9GDOxAh4sl
SPHaI8rEGubfFhOevXs7F2fTJj9ZI4W/k6T7HBl2jhjYTXtEAIpQxBY1DFga1hs+
PASVZ3QYEC0E35up6qjI3/hoRp0H4t8qpfN5wsNUl/GdEXZQKcmBbo0CQbFDtrFC
2MQQYsywiJ85GxYU4l/zvT9MzynreB5kp8N5OOaVlHVLSCCdfiAAN8gaMnxtZzDx
LiXbywYedPHknsxy7pWvuZO2NXOsBb4F5KXwoTaX06CB28R4ij+3Vsoj1g7VwKTH
vtfjQM6+2U4hFiwskDpjxKxmYlmf8AjZO4vhtykVt+sAerPLUSl+uSZupgm/0+mE
bU3nibfSuWYlLYfpxOyY+ttZSZA7Kmn27z53bQKH6yw1VF4DWWV4SQ42Aq6aV8RM
ebnvtL+gaXY35Lbu9LZKNxAengKJsit4mvb8usjpBsLLNr/Qglqf8PTZDJ1e/cLr
hPI/ZZ4+Dml5BWZ7eYmIRGYVy5qwqXkys46AGSEOItP1+Lap47/a/LNYQ/3sMIgw
81kZpwAKpw/fN9p2cXePhh45S2jcct7BUV5zJJdceO13LRE7KMWDWkxDozoRbE72
uSsxJFMKWTd56OUGBPQuLFsqytHdSB7i+a+oppR7Tb6AY0TovL6sT75lyXnInO3H
u93jkkCqYrU3syKUElmJzTqzBHV5LWjCiwzVtN/C1uANgTdeQJlmqcj1oNv9tHjt
BwLLYb2QVK1fwikm3DuNVFh8zQIJnBFFBrzKAOBBV3+i79c7dbK5qbbkqIVL3hFW
o8/X43LotSD5r+QhA+J4aF5MG5S4/pxodhNDBdf65MQJhHQofT7NCOCWQ3H19eFc
BUjcyDjF/ZWWVktlA7R0fVpB8itnqLsBI7ZsbSuQLPXo2V62m8xg9SDrFWD4RKuq
LM6+Neja4mYu7z04LgIeWxUHEU/S47+USeeJxlyO8P/50B1+EsFZiCAY3cRXU9K1
LZZOOC942RoOIwdXNQDc3XEhPohEM3X9UvnxJhXRQk4zdHOUw1pTuumMCXx8Khu7
oolOmLLbjro/JefAfaqn9cMIPvjv5q1V5EtslDS1WhCriibJG/y32Ic+hg/6XVj3
y8z5iPDDJUspJgLK69yreF+L54TLOUgkUi+IeANuio8UNUM18wPRc3dqVMfLWPQu
IOpa1crYeBSqfxz3KLO7otHcddjCOol/Aas6ea6XvCs+ZlNQYiPU+tIvbCHIeWrv
w274PQ3MQXJlCuGAyN3Pp4Yukk6b5uOms8YgLLuKrZufwC4MdUO653UB+quZlcX0
r8UexjLFMVHMLqeaF6I0xBmt9bKwsP0LKQXx9Mf7afJrzqfZOP1SJK4VyibuHieT
skXJRB3PRm6FvCfItvuB6Pj4cFEuag9zJSyeqCryp7ekh7EIpARaB4gRk9YzGfXd
fZMwa66GCGUf+B8QSvM03uRFyoy9bZtMRrPrts2ZQZao01mvI5cfUCIfYbc9AzCs
JMJMNrIw3WV2LFoLMTf3CkbngTzR2S+MzsdrdNlWRoVpJwEdunrAjqCQL3JlCjFY
cSCZ/nwN7mNdM/uIop8Blpj8pF861z8Klab+uHBdR5Z9SyukdjRhEkEfskWAEp5W
0U7CCy8EahSxGLG4WGTZDoCmFH53hYEwu8VoiGrMPqSbzf2Kr5zd0bO1ZTbh3hkc
+pt9UOQU/cwX1ZCttplZul7NabaR/rveqF1XFZYUzLURCntzlNI2SDTXZv/3xjZg
fBC95sOoifeIWowEgN7PJ8Ls5IipNrXGEYAqpnbvPphB3vyLAvVA7VfHpI2hPQue
hQMh8JIJsJKetc4+6s/M2l18RxV8kUqK6z2ywha2Qputggwh+us55gWlxRHmFTG+
BFAs+LYNN+D2M4Rtr/Lm4hnf/uemYZxkLutF06WZHCNzdqvnwl5GuxXlFmsejM30
kGFUd+ukDVH2z2aQcg934QbRNBy2klnFB2+x6W6uUgpJNJ6ze8gTog0tQ6teZlkH
GLlPRLXsZlbveMGqDqW/ca/2LoEI7ZXV4RXmsZxx+LltouitjMaDxsdoZUlqC+GT
hzZ8q2exUvgdr8uEPqwuv2vhziRgmn6s96YrBWugLPrDO8y8B8j/EfwjlV9MfGXK
zPElppPFd1XtpFP+96KQAX9rRNCsIl0piwupN66D+/WPmmVukHWs3VavvOlaBMbN
qbaKdxKj/vKxotcjbykTfnfVTU6XKCHs6OvAJt5WEUmmii3yEOAUf5U0W97lkl9l
LcoC8AKPOIWVmjsLjD298KL/xKiiMWZXQIAhLDwkYXhobRuPFGNVg1/zvJm8YrzL
F6gQ49UF8C3Wh+r6Nz6g25Td/dvppy0oQMDlhgSz/el3fY4ZpEuq4i8OMNslF0Bl
YHk7LkX2x6iUyYg8dhyTpZOJvdPB/JBwbDLTdPPyzUoF2E7wFak81eEfi/RNRZE7
iV9ShkTZfexvw0Tls6QPwVbzIjcth0JQksk1KnNuVNMQXgz6WZxPCdMlJzLFzADH
PI9ZhVqOSieBMoqjbk8cw83Tlw4XOrySJgOOUfdY6yPR4It/hG/Rr2jNUEv1pC0L
FmW/Cx9t+23FsjwL0XnC2scf75iqB7wXuxvTfb3l+0LCGqdJ73qIuu/9K7iBvzvx
7a07h7M3R5ZZnnCJ1Wwg3gT0742Ub5dANrOhKB2HWs9j/t++eMb7xMvKEIu7WlR7
larlF2YOfVyyKXedXFhJBaecoMDzqxDs2Sd7p/Stzq9kcqk/ozyDYiWBseeprwVz
MoPS7GKE3TgUazAy74/fogelrpqzEe6d9Epdxbexx3bxnul0lnOoCt4rEM4j1Ev1
rzlVMqjSCrBz6p4KvkwJ2Digmx2qXFkFCzSzrf9iDHVo3QS2Vz9JWrZa1ujJw2+f
vfPRO17NRA10/M8xP5f5/sKHOhUiYKpM8WkkC1KRPDK2VqR7XodPxIjxVHsq8A49
EIvoeXOFlemhHjyfIdZw+16JT/2az9yb9wtWXQ1oZtniIWCEsMSlN7AdeXsx+8lx
trFv6Z+Dihq1q62Yt6QrOw99OqvQKfSyVFzWjgxkU3juAnprHAqyukQU8ByHil3I
h0I4SXtHnLn7Ln3PEsiGEgZqiW6csoVC0ix7NkUG7EflbRUBa10lglxDz7+AU2vA
LFc43qBHizRi8nWxASLXRZNaRh6Wd3bSwAEiEOiZfe0Eu4hTTDiiPO2QvgIeohlo
rHoRqFEcdJwN964/IOeJNSpiI69fojHrUwlgH/JaG8N3uLERkpKXcs74hXZm5uMG
GM7sbHGnP93ofI1E6D73KAD83gm6ZSRcuWkKdx6VK00XkmEa1tIubmMZvM58UUih
SedLKvvep117pNrcM4cZgNsfUfBAv1CvNwOL6nGTHFLXgBfxigDif3BwAa/5jwPr
tUqDuAQNEonXOa+FGJiZHhxmkk5FY/a8D3e/+/P7LFoUvm9e6Q0vnwDdVhJ/cnQU
GFaVJs05C00CPdgswxvR5XpAdf2QXZ7+JSpumhPLdu2e703CSqjijUUWY3fWmyis
bwjJWWXyq6rGOt1cxKYjIShSpHk4m6kz6vqGMdA7BXDUmAyjdz+xyKyQ6+kh+0O2
EckhHQ9UZ7iQpDhP2VUHurkc5Q7wjcjsDW/dsntu7bR7yYRL+QCgORwlDiw8xoHv
qGN830eKUNca87twXFQ0L23g+GyK/LMYsFSgir8HdI5NyAQZ1ClzgiN9kIttJLtm
3b6mMEmbLksZNWx/e3bqea0e6+AXiXwltTdN28xK/FGuz9OVhRIZLb7aDqR8sOWG
tc4mGdo5njVu6dUbyvBVsyPjLeiGDe6cDpKHpmiX5CuOodZDqsVQ/avdWjFNrQ3V
bTWfGEaWcbk5rxz8KRtqv3yynD3xNjJlHHlmO5BWdYYvLpOMrb4RLGHE4GM+GToh
lDgDg1ABHzDGgTFBrx8zrkRWwW0FXiSYhvKIx9PWyDipOA0FzZIveN4UaJyoW18+
qPO7PFmd1HQBZ16jWH6/fkaFKwhYcj9oVF7wa4/WAQQRrUPSiIa0KavB60ZWZQIk
lHOV/stPIP3u38zzY/AVtlpGUQbcyV0i1a/zhd7UAss1scxP4i9y7Pq7/a6XDxdD
3G+X09uNLb1p+7W+ZXtHAOcnnwFLjmCBKpgldL1QpYDtXIlnCWIkGwdTYnMyczdM
o/C89j6amS3Vy6jU6xn4hofxD0lkWJ3MNZ3CBlcNR4beutCpFPVQL0E+zTba1I5p
K+XHYtgp5xOFyEWkOGR+XB39c5j4lnRP8FGs0MMu7yDM0FIwfHVgkOr4WTWl4m7z
mmPSJs5Hn+akixilOrSJnaq5xTLfZCe6ujlGY+v2jDMgVBP5OK1rnNn8g+/PLy38
jVsL9TQzZPKNP8D4BFN6eJcIKa5JO+RR6icmOG2Fsm03h0mBmnY3i9tsDfjdzUyZ
Ss4ZNYC6vhEu99PusqCSK5z49H0OuQYzR0u4VFkp/7rnpaca6aPaFTfNWEQBcnjy
IsPRqArnUc5BXBw9yCGryWYlPVChwHr1UYdj2VUOEL+3OQXlSqKr69CXeMCk126N
wCp2rbfb5YgPd4hRY2IvJZqrgWXDdTXwrMzgxKqBVHiiw0Fdly02NM+04Wk4wyln
FYr3XmTm5pdz8n1YOV7zXWLGxARGEzajDL4CJ0iRP9qroBN2E6AT5toCqT5Jwsai
/3iZXCouK9fUBBbPESJiNQKaQQXWwkWz0Y1pMR8frX1q8aUB5X8fFQ6o6gxMi5Dr
pJ/X6p/Q/0RUb6CLmT7AcozypxhU5Zw0QnTKKju+jFt6+Y3WONYJfZJW+Z7suGYx
QCn7LX5kl0WwdbxXc4sTilGm5Vxxup8FMTDPqLYFQhPUwHaolZxGuBqETgAyJC4i
0/pk88fFKWNhcNo2Cm5dzriu186mgScksL1kPdp0Ff0IqroTQznOfwvvLudYEgfX
zwW4lYNKZxjEqBWzG6rtR9MsHts9HTIPla9HpXMyu45VeA0UTHlnEbjQBxqT5Svd
tGdL4C3YCmwJed6xWezB0AnB1Hku6l/bkuTqi4tGIHWiNweBuYkiOX0Nigi+zWHH
g0IwJF4sYN3IUpXWtIljnb3FH1OYKpG7h1t5weIeD/pzETm7OJXwFft9uko3xfuk
8ujRuBAb29n4YIzgCwhX2vks2NHAc4StW5M6VKxHa7WA+1/k2mfbmNbNHkSO2nT7
9HDHPCLxbHIJjGxQpJhheq3R6hnqHKObwgTUgBoGu0ES+TO5DDYHSqMak5aU2WPW
Youev3x1lfM1QN+Fu2lS+Dl31oZB2f+1DbHWexSP60FboTg9BDGLNflMGAN/Dhy0
wWooagDxgCux970UetWSwzx4/+o//Wt4lSlAYjCxnvHhPc33ubhvoo443sDLeUgA
P47RxE6hnu/1ChCzq+e5KpA+eFbqNRomzDD7Y3X8MQMH4HPpQVJlo5+HAjc0kGzV
ASKyNz3F9hM83hrvYkJaK33KGVz/J2sKtSIGMWRK9/MWsgoqVCh8pvXVgnqC5Gt4
CJslo/hfh5oILX3sqUDVSREZtzxXlMFls2Ocsb/TZ840WBBfKLxHfGd2aotyTlWK
yuCtH5/7cUZ6MnwlEx32vSSo2fxUNQn6gUELJg17HljjdzsDx9u3bKqxSuFCQ25d
ScReAknh6ycV4vEwZ4qdWQzP7K/xu4Obbaw9XVJovA8k8h94wShKuA+l8QBpBxzk
ODNiItSaHjxhTAooKd6ZACO9kfm44S2s/x1OkOHtYg1H+MIfVsPE7WJ9AyTPQ2nE
Xx4w5QvhBQpy4ZmLiwUxrPJeALbNK75JOcBav9tizO7cyKENLNqO2vJ4FX1blRH7
yds9EP/kATfuHk37dqpLHrb6rv0vpx6fbgrwltIJMf+CqMXURx+JrZFnVgq7UKdX
Cl76SmaAtfjt8ZxZ7pdh5dNBP0lN7UEBapAhxN7LUmKvygGwi4aIpp1f9D46Bzmz
8qVQyhOi8i4tnVJIZXMphrPn5ZLxtMJPZduFJCYSuxjAYU3rnniGcvbbtIiXdS/G
fTS2w+3c3g4RFCf/9amIwjKgqJxZZwU6BSxMOdkhwOukAc7gqYwoQWK/CTFKpi5z
Av/bd44n8P+2RJ67hHMpGNvRKjj9BRBPynJEpHkiU7FkrIH1Bv0iym73655OUGI1
TUSSMyG/7O7WWgW0F7xAf2tlGxNAY7kcCtm3JQ0t2fXc4kQfEKipCTLgDOrc1Rcr
0I3G8USBHk2nVQnJ0eJigfmjvG+UJhpuC50e/7VRlGsLItUVw6cMPoXbZUF/SN3x
r9Qux0TT7Vel86xVRHFl6S+hzYyE94Pt5fLFcblmj9OBjG395yt4YxmfcQoGpoY7
401QIVcUBc8sv9fL87mtjuCVIBUS0EwAkP/eVeDU+LUChgtI4PuPJeJypIgp98r+
aesjFom67jlDSN5LTnXvjlvnz5K6xUObc25u8hsud5VC9TbpqEdYV5HIEFAKztva
qY8EFhbJsxIa1Rp7En7tLogRwZO6kCm8PVyQPLpnMMjShaRAkpD1J1qFYBaTmKVt
uqoo5E8F9JQJgcb+h7E94zKoEv8LlJ4AVo1IjoJhD3cngN2L2bE+jGe5l/xWvce7
27pMQbN1emdWC4j7UHEuLD8ntvTSpsVw6oFtrcw6lepGmk9yn767xFF/N5gTjw+v
07QpTkOOAVLnLml4R6m/wMBUCmdDbWGzWdRs+8DRUAua1pUscXL2wADenjMPiyJi
2CF7XURfItTDJmH9jU+uWry6NJgGAIrZbq0jcfSeTl/T29rpkaUf24grmjCzcb09
Di6Aj7i+HUYRmoZBFnHuuwSVcOfFU/OGIjaWXoA4OPFQ2VdIwhyKKduxqTh2xaVa
NG73nAt5/+e7ZNo5lT0RUK4jdvwWM2w9MDbmQpHXVRwtE+Jxl2HcEbUwNDtLUF20
aECGFkkNAkk+oFwntW+Hy7+L1LJigF58tRl3QHsLdOCgdJAro5V5CbgEg4CuCeZB
y/W44LGxf1NFbPiJ3BSbNR6wrQaV5LuUemii8s728K1l4TeZOUxeVor/xYxw7mur
/fhbgCItAckKdCyw4FdmrZRsUwWit/KvSPSnfihD5wGe28ekIDS/XCZiCIEWtoAa
7tZSSfzAaotI9MMnn0yoLLimfAOQaGc+vNzICqr3AynwHyJzcN60sbj/oBCVrroY
T86A8pNS4sMhax0r65a9Txa38T3IjXSPmIV6tcq+2wCtkrxn94eXRS5nq3LACrZD
nI50sSUf+EW6H5n+UmdJb5q22IJPwoku2WQwxPNWpUWDFvY6xR95+uVwmk6Um3oh
GoxhNSmKztpiEzjzoaTnwdEe6GTjacZRCktKOt4chlT3PFBBO4hxOkqEu4r90/hY
UBh6uI6h2oDDwX2oiD9fCjGGFF4Ig/wLYJKElgItCR0QCkMLdLILbglYP8tLvFZy
+VbxDAK+YUOAiX+4agAMDWDFaqwtduZ3bqvTOoW7DdocZmo/KgahdHs4v8pVWob1
JmuoBtm/SplS5kRAUiLDb7KzZYpwQ1s4DEbo1RCYi08K2Pq+JTc4BCbEvFzRcFeS
Bm7tekVmlxRkMyqPDsV0bVnfC3DZylbWip27rNdpbRrhrC3HiEMwIa38jnYTuveH
J6BIm+08EEprX9Rf9G8IJKSYjTafpyVvvD/+Lw5OJh+Wn2+Dbg6ywd7IFGHRWUyy
1qZlf1MB9W/RZHV8S23CnnF+1TqjLzDg10PtMD3nNOBEp4Jx0kTUOtvLfHCgwJme
RrLm7JXwAMzDlkTZan4t4IA1Tgm3GXhfMFRniIo2DCFr3DSy+yAp4LB7AsW7n2De
k+qQuhMUETlEw/PpyM7an++jRchgHTVuWu1yS6077y/6Jl4BRGMQiKZIk6duBUk1
jlFoPXhFzzaohQC7aSVV0cU+BqVCfyUXEf9Ir1xLSpGzfHvdN46zTj5liXlP+Osf
f+GbfFyTuP0fQV/o6gFOcgY2oO2ubgiqwzrnL8x3rA7WreMk6BRKGjumMKK3Tlda
IYzY44+7eTCz+6sax110kNfY2JPwq/BlecWeZWYc3ZJkfu2TPJ4O3fy6vyNRbXQy
71jjVcFgrWZ7JOd1PaLgDNEpJ7bZlcaj7UCCi7qNZa6+FOTs07AiXPLPeSgaxBNv
jyi5Vd7r/SizRw/PNFGbTsXpM28Bowf2BLjzuZVk2P9lffKTnW2jf3rm/Gl7isLG
yX0pTjqqG9UICxQQXhK6yVouBfh3sxWffV2BJBTHhetunZ+GciN1rzcyEO0Lu3fu
sHmP2cUHa7aNXZS3q468Ve4XmRVVF2S7ubhtVHoY288eX+ks+zoJvU5666KBVcKv
Csqf+bVA8cyuQ0Vb0+wqUyTJcUaVZp0TvAhGXG2bWR5Wrtay9w0Hd5EavBtS20rj
MIb8pq/0Ov1dJvuwSJwMyVko83QyWDD6vQhKqCFVFB3gEymMv6ja4srLM5PdR8T2
3XH14iRvEgSGplVUE5slHm2leOtoY0Y+UvJWsaahpiJ5nhiaN/ykAx4W1lXiScuT
A+w3glJ2qZbZPvdv4NBoQi/kzZBEfGrCh9xcj85vDjQcZsXJszoTUveJr80LRCW7
jmDSusIAoKNj9XlV2X8isbTA5Zjfho9hId34FDeT0SOQUeGZSikWoV1eE0CT6zeZ
RBDBJ4pl/AuypIrav/zXVdwqU+5O5DWJgpxirmtKmkOwMF6DDzMJIF5RqTRZS5dc
8aU0nbhmWHt+EbBgTC+sYYU39yzh48xNETt1rFTmM4P5jEnPAcc99bdPsMj4tGjz
BWdnFhM7EHf96n3rs7zG5B9x5TNi103jtzK4MJ4SSRRjUoSzePjEVqoiQy+fwF3v
AE4e/cVRYOQIOgmlWUM1EtQQ3maqy+bpY0LQmV0ousb70iTh/xxn7CdyKFFgYV9X
FvI2caNYCNgGFCi5kOPsk5ZUgFWPVipuPqOCjW7lrVgxImSEI9iobH188xZBuMUW
3qWrxQgLuGpQJaRDflph2HkfGbtUFEujhT9pSl+0xVvhlaqJn4YskFwyZdg3hR2/
eUK4k256IGdnaWzdDGg9pu3kRXEsO/zRL/bXid4pZYgKWuivJoO7UbwgM0usC4OB
r2SactyDgvxhvTtXWFDZjmGuMAUVOcQcpbpw+bvsv0xE41KohVrQ6jjBE9vDv+UL
2+7mLFFLkWbgW4uhuZiFIDwWtZN6UOvtrn1D0+CgJBsUGYWvYcF1q4fhhmTfp5os
HBLcG+GljsmAT1/tUtEk6L8jnVrJSxLYS60k45xhMRENuT5/2CdPTCg2rpQKuTgw
ARjkBxDoBb8+ZX6o2zkCHdnj03QpvQft3B+IwflYpDPXgbY9nPeMPhM5pB8ZDKR+
fRH6B6PF/yawwBvHy+WwLxH7ZPAYFaR0xzSKKpG3ZImnNIrgzefc/zh/tVxJnH0r
2DW35zByUhwSQv1FSJvZ7qqrlnM8I9oAzS/PTflDsKPJ6p+B5uhepl5PWbtNSLXc
2EJYcpXLsqMjzyR22OqlHCAb3dqp82gu6ACYjYZvZSCooWdKtsP6DncO+230h1Ws
DrMfskFt2biDOeKnelC8hspixM7/0wCUHrJwRDqIWqXTag8GDvxq1Ayy2QXBc5ag
nMvYcCV6WOZU+MBvb11ayVnUAFfJC7Csz8rMuoJWio7+52cU6o9gtUKQ7hTUhqpf
qZK4tO7A8bPmGnnfPS6tiLMFTvKDC2Ns3glNRPkVqVVgXLLUumZEz4YGJClAyhBn
9fcbJsRGrhy+ihzpnDVhSnspkhBEBq5erUXRvt9wSk5GcuqrlfMiV4QfuWYwb8DS
BJ/EzqcnUiaXkjyNoDGcqV0yssI089dQb8W+U4zvbBXgnpbYBClV+5qi8jy9wEAd
ItOV0qqxIRef+xA1SKFTDWYzp4p9w4YgQtPaVRj7mapM/KgYth2arrEkUaeVjvnG
t8cqd2h9RRppB0MeFOu1HtUA8xQuAN23S0LGeQPey7rEQ04MauUfDCqVCgKvK1d9
R5X4q9AmS9cZ9LCMtkT5wiGjqAplrDLMVKCrvlQPYprA+OxQuYv+ojru+moAuIsB
E2pz7JokEmPD1J8wIwdzHvkR4zSpHULcdAUmv3kAWDUsbiLRWakXRbWQdK/y0tva
maohVeZTbO/rGw6Mgiipmp4NocA+c3SBURyj44uSvQn6BfywqTouqFtsdAMF3IGl
26cR9kJLmdFyN7z7jkZ+qq6o/Da2EEImyN+qFZ8//8VutpYVu515dpGDwnH+YYME
DT2uozSSXv3ThF+s0gMlHQML/3QbXZWlpPThThdLNN1PZTGgLSNgrbmKXARnXgZa
gTqB6ZNKC+ZbfyzIC+Na1VjEPwu8DYu+9mvs6lqP0Yx7VLy780EdY0XzqGajroff
BrPrWchHxfom7R3lzcpUL7tkwIxYqOuJtSLMZNw6oxrky0CBNR6GlIgbbqKgLChK
xasqr7Apz+znPXaq9h8m61ulo7yXyX+TBFaM0GAp5g4VsWu9qTFT4FZHx6tpuo20
/sz/L37gG66IfVax7+Z2xR8h9e56hjlpghZsDdMcEzjazhlu3QV89PZzN81MEGt+
O7jzD/twVKs7X5FLt4uOVCQrvljIzUu8mz1KLyi8FSLgAcg/IUYPkKOHAAWvb+/u
42wrSDbTpU2H4Knv5unBIKnddAQtRelGKiL6Nf9I2hHRdRDqfw7kJGB7Iue0XCEX
v0MKdV2UBZYrD+366iHvp4Bc+jGy8u0yjQBvdXbZmuJrXY5teowsK4Q9HGkgddLc
AmkbelmGO5+hPgWhEAkg/gB2X0RdaNvnQi+ziW1Ohn2fQahPxTT+1RtLLQyUWvdy
XXeMPKM2jCCl/NuyBh0koCW1+dcc9dwoHrqYybcIwuERjItbhzmtqjJ+wdgmy/Sf
RZvH/xd9qdTI2q32E3nwgw2CVe+sxv840GprRd8crizaGPKpbVBXfwqUnbLDO78d
oWoBxmXbMMo1GgT6vePlITxMBsw5OQfAM65PwvfhMVMuUwKeV/zqGldc/QjJmTN3
1I2R1F5juqGmjY1ufq3mSLu6pNnaOIfFyjalQCIIQggG4EF2t4qeppgqd9A6N4Pm
Qkrz11T2nKDGSTNQn0noVJ++lXhrsPGWexpXa2O7ThJ9f/S6zCHVmn+f+vOWoFup
PSBuOJiOgfb1vk6BTk/qQoMymJI+nifg+3/n/uj15PTnaJPOy6z9VUM2dsxS2CvN
qtpJ/gICOuYRvwfx6Wk1SdPjrwSRgG6tfbnMxw+wzMMVPBOpK4nZmWERhoT8f4WH
0urzTQg3FhFOye6N4JBGXbZRcexh+NYxe5tvPMkaHl0Ivv3zc024h9aM3K+8Z0rS
F4DOEV0VycGu2L3NZNXu2jB7KT2Ik2UoYXK/kJMPgM0TA0VhqBkE4ppV3fOvzPI7
UHsBq1BIJR51rpMhdf9hyQKFcHN59ySCseBzPhD6CMBrxZtuxnQQyz1TCjPljF+8
yeLLUAjJ0KJXz/k5I5Z83yHWpDpqqabphepEmiVXBPQjyH8HleRmOjW5x9MsWgT+
bDTxCuZPj4TTzSCEpPISpz5lpmijjURqKpftGOiKWrRtvscpqVCHs+2wueIFtP+0
YBPvc5UEkZYqvHqfR2dwLuFzd4RWJwe5bh1khRM8xvW1G1rdaAZI6/bukR6UV2w8
xMjOORbSLBDoL1Vu2aM/k5CSm9qM8QiW4lFk2TpVOGOyQtt2VgSjD0ROPAf+rznc
HOEEiGJK5xTY+7l4JSWccEWLFbsDzupwzDev3q5Ui1R/DCG92tTCXnIS2EtevoaF
BVRsbLsIYdv+nC9oSdPufofNd99pkZSz0vGGGY2a6H25B3ZPLIj45iH27hxDLRS9
bVgm7LRrtQ34CV+Vs0MdOWRXfIedp9ZBn76mkW50MoVDrpCzdiBN81LMu6Htlnso
Z5wfonU1+gUB9rXY6GsgvB+rNYgCz8bw+3G8QI9hT6I8BGXRYvuUoD3dKUYnzz1f
X30LNfIaQ1z4fz72F9J6srjmTs1pFC1gVoT1x1lxswNjdEVmVMODrPqzL4l0h6jC
bKELWqBul6AV0OXatMwzahGTMKNgC+PXftUoss2NHlnlj68Skqro0m0cCMqkae0S
KgSl9ywPr+m7e/BhKz+2hDWf14wndkBpXT+8D0o2XK30oS/UDSA6E4BjRDRUrXr4
9yvtG0fYwI1EgUcXUmV6h7irU5essU0O2ZBpN2WyAOt7VnwJu++0CTuZ7ZWpPNxl
HJzTxcR25boeuGsoTDfsLQfZdB9g/gAfVGdfZa18lYn41/yoYCY2Yk1jqRxxsw6c
IZI+CzfwUCVNt91IKtZQRPR6axBUT1/iEQXOsXAB1XdzIrfOTwzNKHL8M0YF5BWO
nzpk/zDJSAscVS9EG8Yr8zq8MIWJPhbo+s4GgjyZlsiUKS0CkXr+N8rybK//Kvw1
XvIVb/qaj8xlOnBw6O7iBM6yJC585PAtBiKlkTzM0gJPHQ++U2pDVDZ/M6mLD0iC
5g2tyx6rVuHc40gM3dJP58J+8o8u45hoHhW5ZzcwznTyzvfPaHY872EG5hiYC1Qj
87ZqkPAK1PLc66cE60HOQj+ykLKOGRX1djnWs3S3TqKBaOMm+Qq0CAi0c0RcF9bC
fABQj69UJTQA13QBNBDUwq7t7+K3/Jyk6qqqafD38vplGXHjJKIfb4mmWIdUKiY+
Qb+qsz8EmdH8mH/XG+5w46sofAUh3TbS1mBYIICHAHYtEPaQ42zPP4w8fpXh/VSL
uAsGo3xkUCwQ9p0fa2yTYaDGPfBxSEKyWVpuMrj5w+kAXMgYrKuNV6dYfZYC3RdD
6qDDbpyZ7iNUydAi0hgzSIQWpnAVbqP3iOewnKENMoc2fauP1oltKxXkylz0TUxd
/yYd1JxYSgZx9oRz1YVcsShCcwrQhuvv/+NA+OM9uuCcVnp67UMPeYgX5vE0PBJk
MydAuvVyMj1jrjKJzbnUSuBB1YUu3HNhzcEjapY7ZC2fz2v1AjBLHmVTuykUwlM/
JtblNZdU3j96OoJSvecGUjYj8ZaBYXXxUAFsOKLDaB37Lquhj4K3YrIuWeSj43u/
rNlOkuA21bjn4OXOxFqfn/+/4kw44rVarQpk1/BTcJkLYQDWe5Tucoc+Tug00n/+
ryhYMHHBl2tQyAofKcD73NnNqymFvEgQ2VJR4PUq/2mKLTYip+oZTF3coPnd2rlS
n5UCkrAmhLlj6i4UjeFwWBDcEltWJbpfT5h5gIB/eFKm9wG44HI9fEKHsGdC0oP9
vL4y6ngSw/nLmuSakIWVFKPw4z8MH51AGqlj02bWClzgmpox72aeuAihT81v3dSB
li2mFwQtOxrKk4YJTWCaegV/FHHy+9y0Ji5NBdoZrE1z9iKyopKTK0kVVxKuHwIv
ZhSH4aga4ZqJGn0zynSKuRzArZkgEy6p26omH9ilH1Bg4w6042uO3jFriubUF77/
uzXycf8BtmIm5pTQwCUI+SE0Dv3K39G3qbcoJQmho+eQqJPdYQASCDt1H28gII4o
f8/zP2QBbdui3U3URhtCNr1qTws8K2e+Hl5BIEUw8An7TmyktuuGT/CT72TrVQoX
UjyYRVgpuysHLw26W5+Yk5gAQHhqLWAUrQ5e3RNFPO4yBFFBdoATXZpM6Flpv/iI
jrqRPHmNmpVFIuJ2vca9YjgRDPxTOM2rIw8V+jmY6y2Rj9gTUSfySHIJk88UMUwm
bKiwT/ByNuz4MdpVWmenByrJe6cubh8LCzgxMIDfmP51K8PVMrmZg7dwBSMbJBj9
ZMIR/HR8F7x3qr2J2PFeNo0o9yxcVr4frPkAX2PqKhnaG67PF8J+yMea4sD0kMVc
cWHsQgK6GshCqAhs+VL6fJ/K2feKPNP/hnaunZR2rLGH+YuGeyHEmPNHZLyzEWgS
lPs1ztoeAIphWdUXGnt9V4nvwETC5BGB9TeNXh3jVB8lTZu4pHZ5YGjk6zRjdmvE
1ykvLrIKraa3PshB3nm6NPDUcKUVdXHHJeuw6ycbWvraSroHnUmTtW0kRHWEj94k
CCxTvCbanjO9EOCvjn0+TCEVkgb5iLIFyCoBUUUbZgsAMCmgxFxLeZOrLr3UXy2T
eGobQ+gPPnWfrA0XUe8uZcQoEhiIJojfAJI5/FdXyAVzo865mgpwoqDHlLcEjUjq
SN5SH3FU/S48llHImnuLJxsqcOw/UpBF4eUDclWukrR8jESgUqhV4DfMEPKqDkPx
sIKQPN2B8xCtvUCUFJ+xS9AY2E9XNfPXi1leuboimbzisjEGt/aqNvEvJAx7fq7Y
JmgBUZfpH7dZfEAIppo1ZWIqcNKS8BYqPRI/7nqbQHM1eWOKg9nsFT2XXObdBPPo
94T6YCWzJkQ58WBFNc8mTEdHVrwH1YKjvBV+D5ea0viZnPKrG0CK2eSDiDo53Syh
Av9mRi6IbEwtxOwc8l3+Ym2qbl6Ag8idYM9/tRaOAIFN6rTuhmv36ifmYJY5l4Mo
kzSk+KOXJHxQyfrD2b402KWmiZrbwMo1EopW6i4Lj379o1Th2d/atUnk7pw9Gl6h
jyXXkJLT+SQowcfx8nMAOw1PvsVOz+/P31PR4klSDKty5GRwsAElWCVq8VVQRiiq
C/KyyK9GPalR6JGG6bvbg2fqbUdkqOIs/f29hGvDvByVPpLKcx3ut+nouO0JzrLh
o7HJWLnpE4aUNphrob3ryChnSPhezhslj1bLcsV/gEAup7MF1En8Kpc5PGJFu6ws
wFGplvC2gs49rXuXDgbM5M6zPO+Th1ad6g2hFUfg7BWKp6b4OYe1gy7PuXGuW4Bu
xh4uwCvSJuYEgIL2xzkQArG4K5NjOLF6PYWgXM5jHThk3o5U5oNbnZ8FokvQYPZK
hudg4ajJKrd9QPqNqNoMsxH76Tbnggvo4Aur/HQJXWAUc8b3Ej5T3QGu1neLHJEh
xUMBj/HgujY0dxrQnSHx2sE8F+y+WtcidK762jSnG8oJJKy4bp2rDQkvCSUhd7q2
DA07kFQaW0cg74B/anqAdMu6ZLUJDVbfBLH+1WiCcjaFKQ8ZDnx0PvVNznADbPnD
v1qGk/M5UoA1GbxvO02AliOejpsnO5DwuuXBl3eyBTi3RsK1M1Mjl+A31mb4NnlR
csSbI+Dh4aoxCHMp/+Qws+eLmYx2mh1gQiB3Z94Od3bQyfp45tKZ1stBu5xxh2Hs
BF9YA/nBTiIeYDKhxp23iHws+Nm324l3R6fYVF5zJ8jZJqcapInG5julwD6VLMta
RpwDTCmdq43R8ZUwzA33pZL4vwbuxpPleIbh8aVq7+OkNCPNa8tCe6RvT2ddw7D8
z3wmyQPjjz2BdUiI98+LfQbURQV2x/u/NwhtpvBzhnmhBnuuIjyBBvjq+vv9Nu3S
ier3xDW8fqrqYDx/NWLdJQU/lG8phQT77VcCSd0766wuJA7uKT1AkJOBDM+pKSEL
krPYmxEPhf0sp9mhz2I6aDtvZwPoNHIZqrcPOG/4zSHyaihIaTi7b6uo19QovE4G
ZnxQsO8rtFARf9yupFXcY30avbjWZXqm0ZBfy/VkOGyqr1wxhl5AVa4CevF6nlqr
OPZkTQMw4ZIifsJh+AFyO3EnjVH+vWrT4qf4B9kAQggXoEY41sFNpAx750tvJcBM
ocCm/sa5HG09WqFp3KDkZ4t3yNqlzYEXeGIOZLCVHd0EJUNmm/gbTGo/t+y5AQHO
0e9QQYheE1ljpML8eRo4Kx/VsIyyqGJxlU10UvBRUeB9mfu4VHbVKQpg5ylVTOYf
edF0sz1dGBr6H21juMxPMYWzztqnkT7Q0DtJJFOGeBlp0YwfOxkufhBoftGKQLTS
+cwwNpODAvJNroFTKFuSXZLdoRpoEbuBlOwWIMvOJAtVVVFicnN3DEsmYEioETZe
H6K4xNr66EMULF1WtOeQmpE4SiZlSKi7g5P1nd+k0m0jWeRdOZ8m2Lm0VbqeDrMh
UaM4ti9mm/eta7whq0vK5lXLqSO0VniT7alWrfBf47deWnd324qrbbbpXQV0k5tB
XJFhF9rSasRHSGPq4UBz0ZpciBQbVldso9iF//eRzN/+jtj8cS8ZAkFKOMmz9SQ6
6GCoqVZ3ftYD+vfqw+YEouqrP3Oq+MSQb/KX0onG1ydO1Wk9xRnC0bPLfFvqMVqK
Oe8a55dQC1vVzUfwFgn95Bu1Fz+1+9xB7CwVQBwE5lBsxchJqrtqo807AVNaQ3QA
TjAnc56qUIPZNvcetejl9nilfQ7TzOSWniNKwsybuj5KCuOcYNG9XSdU7yZ9g/aS
TbLhK4lIxM2RahCsc0zHzvRuisxL+HB3+9FiDHhBkqKUjH035r0qS8uDO+I0CMe7
1IWH1gcqRf8bHBCziEXxh180GGPt6l5n7CnXJ4kxI5+yOcy9v9VHggVbQo/W0llF
/SycXLJ6ECr24Rm1w7bir8kKNAEiOn00uZ2ab7/5YuiMO+Ouj8/VCGUa2bZvRX5J
jz/7u9BsCppBuPa5obUD92w5fli32xrmdCy+r5YRdwdv1kmfMpJUQYAnY2/7W2a6
5TUfP7L5/ga1trafJlNwuGofDkfimfXh72zi43IB/+3WLznz3B/7npv3vlpatYN9
833bnvCt2Lq3xXCkBop6rVIHTH6L/i80mSYPRDSQht0AxYJrQsY5FhtC+39zhRYg
0a2FVsWODRmHpi3IK6hAuUJVIHrJzX7d3m+SApvi0YoQKUqwDctpZ7ZzAe+yy1V7
qe0LwhCw/YxdczDf9TLpnb1ASXrmgV8uBRv82oatLrwykKs6XWOKAEeQY5ypDtNN
h/hC1vDhccOYn/tJW291bsgCUVLaZ946kZSiSouwapSdGOvVYK5Wj467/uHFf4vj
+XZD0cccubKmBhUQEuO0CZgZXbJIpKiHT7i1HB5hBpPbGBMcmnevE5b6c0JeW83i
ELUQubGaK7/XtHS9sJZQTLgeQeBJRdY65Jaap3MqRWH7cA0YDlaQtMeWZ13BIxp8
2hZ8ho97ebGZxnsvUQgiMrhHiH1X/1pEqAYpBrlQbtIgWUS0QUKtNo/uYoVDZFme
6OfF/SKRL+CBjDFcY91cNSSroir1gbzX3iQkEZvmP6epmOZGbfCOg/oAh7NpA43U
N3E3z6BWubBND2w95ur0d/ANzLVt2E5uZRARJexviaGTrmj5tbss7AL9WwvkAX1E
QLVnKseNFrL7Xe+ERf1RT67v4OdS2iZaFUzOo+yt1n5GJewL9TF7qbh80x3P7EG6
aGUHZyS0fwOt7leaCgfXKitTj8sIKgrf78GGRCpVIz8xa2ZTcETwKdI5YllwEmdm
VuByPy6U2LKfym8lZb7o2lXe8VOoB2uGShadOqbPQ4Do6mtsVtjUUjbg85A4iPUz
y6um6DNBpBRaJj0N83v97OEY/LczixH1BPi4ju3UNUdSCc5HgUOsOTlctr3rpG/4
cYzkbv3w8YCqEp4izpJSCzzuk90qlPWEHtogRxzZF3LUEvp7rX4SZxzON03cWk+u
E7ZKpcV+osH6S1Ce10EFPhk4uf+SpUzOJOgVDjEKx1LQaUCIL3dUjpJeTaKY/Ncv
iMuSJSylOSxrY6z9eaHuoCTpgIMpbGYzZeXY9b6bP21jn80bTFI7nppp7VZcqp+2
FJoRostL549Msfxh1IXAncOiBCt3vHvNWKGpkZ64lWf/KKTjeADwbTM2P4W8PB/B
Qv0ujWmhymNHge8iQtX6WkGrNOHzKo92HBJ82UPjqP1bBTmbGGIhhLSGEPxGUQbd
TSWamUFCHyIEJFbCXOvfYwYeBQS/OT1Xjt27U7CypNqm5Y1kBW9/kTiUUx6u3nZm
/QpEYkOLpVpiVyWkat142cy2XJszDtcffIgsADFktQebeAwvbvg4mRvrIz8Ix6Zk
NYQVY+LrMcTuTSQaw0JDN3PW68L5kjX03VOIIc5fxjdNTq56wLa7bYqGX7RK2f58
kJAU7yb/d//OLOb668PCFfHxV0APLYNfSznScMQ3pYtFhqbm6gw8KfvVPgLNd9mG
N/arpUG6w6IwhsrtYc5MYeK6DV3fuqb1PJi7U/RiP8KexiGbgfGMsXju4gFlxCky
ZlWbXFJzizrFauVNAo1c+tk4sCk3GnEs+FFunjR5X64f4qVzWzes54GQqaRg3RGb
Ua4d+AScVrYwbeOoeSK3ZO1Kq94uLMrxaJDOv3Och1pPcZUWjansuHVoFFKBLHfo
BmtwwwHDE4DPgbPe9v2D7ASfXL13V7W1wgC399qP88b1SxujdtUf1oo7335j7XUG
CxhDcJkeSEkle67eqBEoDONxjsmYQlWX0lwsXofzlghaFNyksN4vRa94Gx5AdbxO
/gUSRA8rIVsusNPEh7fQPRzZ6SfEMGZcbIt9DIpEG5suCQpocVLm0FKeorK6SDfo
4wYNval4BnXPFWUaqjIQmfPaASZFqfXO+L1wdo1UKLIn3uYq0H8wTSn16K+r+5Y5
v/qG7NHpP8SmuAEq1jGoROtbfNShXZfDIhVfEy0x8n0QPwNQsFBacg56mIHdmk3l
A48cG9qeelZ5jQgi+JgvjEPZVapwdDLQPdmn7/4Pgu+23s9cu9AxZ7KAPcT64QKg
Y+F6gRgfFnSpyCzXXUI7fxhONvqBTkGAmWY5cB0e7XcFecb+ftZajOL43E/fwdgd
nywYG6Efd2PtoPqDAWBgrvm70VLKXK2fekzE94I5GBEyeO5bD3sBz1KXeVlVANa1
SX7c7mNGlnSMyurwprItKZFC6KtQZsqzPN3aJillKHJU12F3g8tuBbQ3PmrIQDLn
pv3GhKvFFMlgL1wBzVryLsgOolf/QJRGWUENG5oZ9VtWxas6X349NqWPcUUI15K1
REXWsZppRoZdMNV95pIjbaZhb8PyTIZzSnF+L+TGX2C/yZD8lBfcoxQ6cYiNXHyi
X5P2ID4nh7IwtWSt8Y0uvNWO2jmbx7+OR8unM5QOGMf1S39uPz84Rcu0Jqxt67T2
UylznFRNXwcTQ+7He+C+wXLLxxQfoFIpAJ22Xj75dG21oJd7yWnPLJzvoKlU9hHu
WM8QzKIoqTo4QKQ5rwBvA6dvMxszc6VTNwwupsvceETp0yc4b6pNxy+TAkBdoVne
CyqrMbhEPPdQpkJtLz8T6hcFKZjabQuzbhndLatVRTDShPwOvej563RaTW8MNWUF
1Rhzm1/EG4S1coxGpcchQ4QU5/W87LoXJR4+De7vDQg6JUO26t+BmBtdzI9ZTUPs
T+enc4auMv8lkHsOGRghR+X9rwYTUJyIXcgx/XEXXMuTaNvdyoE9hAKN+bPIGyie
1gabHrSc/sPqa+Fi9ItqvZrrv/tsCtzm//49WmhgKcuwaMRVj1bvRrh0nB/CmyYP
wOhrc52fnqNmqKXWYFhaGcsmoE2XATkPll+3fRUldA3UBayuz6EJcc3D8zrHUSDi
ANU2RSL/+BgohRkS/nE6JVLMLsdMs0UmJpWmazXgyK0pYBeDosWQQQbHVoqEpVe2
Sf53PplQE4LT992kaWE1Xf7TXO5GzV17yYOQSFhJia8wSvcX65Z4YELIRxadZtkm
XTYOB+vWlkQBJ4FBaddyAHGHg4LwSjO22rPld3wbD1Hw7A0l+AL2HcMDv28rOwtw
8s8tM1OVQjGnisvnkRSMAhPkv3BMhz63tLWZcOfwYCfM4EYNJhlsmeJcFY0fKWXg
4CIdIiQ6KXslE7uOeVL6+hWl27zJDGgVUyWrCx3NA+xjHDcb42mTIdJ0a8F+6/Qa
kqrIhnyIaOd17jZe/gp0MFTzQQhwKQ+QcoXu20nO00+6MsBQMn7j4N9BwyP48lrG
Sux8p51o/R4H6PM+WdFgUwU4HLpBsBsI8pTDcmIwOLrkX3lT7IuhEkiKKlU4wkzO
RxzrhFz5TciVuLHr1j3ElNDu/8KJT0HFA96txYkBmTIgMU5sN3P/YRjTjN6pHDWm
sO+aFOCJd8WqvqjbSIX64FKOtEqOuoDDrC4ZJFXdQIrGIiI1DwBHDaQtrAFD7Myc
2NY3dhWptK30Ai7jh2k8RIXKsC4JeNp+tkXn4X0lYUsHymhi6vuLcUiJ5b7/tFz0
tv6LD7poDHE2Hm80xnnwPm9r8TFhdZ16JcgQi0ZS84k7BYuMLtl215jPIH1XPI9c
Nq/JufteXHoJD1aWxArKUObYQUx/+b2k2ZGJwNFgbAlN95wstM5nseDvBL34+UFN
VxoXyhhr7euFE7FtcyvaZYUAMejNH4Bspgu3rH4LPFmdryTQ1zep79pKVN2KDCIm
oJrGLWZGhlpwGtczRi7YOSSHKYceeCoiranAXrp9mI8H/HdKwdXfdxvcReeylF8e
4zow/Gcny1sYhsXzXKe6bQ3VP2oUpPRUtsZ/bW8D+FKKOl5923qQFTYTeVJA90+S
Wtp0UzSjsAJsImpA2ut/W6IiaXRN02t/dSiRd+Sq2697wOKgou4uKTMo72sYf2rb
juYa6miQhsc2mJw472q8sEN5vV9r4X0iXmgAgJQs+AejJvwVdC7DGvn/Qw6QUl0g
oxxNE0975AHkWAUMJ1juyuFW/f8sIuwC3cccRNTPnN7KhlyT5r1UacWUOzb+3fNu
0N5yRwdP00/NFLfuiWOxbn9qGwHdtz6nIW06ubrf7YnPRq4IjIcULqp7p8U3in3q
FYKFWVx66Lq8HvcGFbcCV6dWxw9I23hVB0kobdrVw6TgxXfRVYEjfOdlWhM5lnkn
HQSeYSRtaHmXsBWnXpFZUAkwddhx36VEiBlIRuszd5R5IuTXjFvARGnqnxr3xPzH
Wk9WBjsFzvDYbp/nJlMplQdA8Dt82cFRbLMgxcl1m1Du0EHqa7eiYKH5DYe0Jl9+
v4MiwuyiohnTBmteQVS4+atVHgZbKdwryr/KpuqcHKQdsNkwTehMvLwaVqWgV8/N
yhUd/gxJ9K6JMYtFaiVldjs4eU9QaeC40Af2INAGnY4ZHCiFyD9jqv1lMKysZYTK
qST2TU+6AgPU9lY5KHn5r+eU1pvUbRLTU/IBYRjVCKhykWj0xh/2qcPlJgO1W5OZ
UgT1ko9/oZRsJjXmT9RBDQ4hPFCyj8LLuZp6RkTHnSEGLOA4IuePT8zN9eDDwNe1
5uCrTxw6CYhEEdTme88UEKgG9K4i+OMUfxYP/5bOdp8/4tl3fBtniIfisw8sOm47
y9ip62EfuU0e+fJdrexCMxOEtQsoJdKcOiyPOPyX9DC5dgHlI5x8Q78Cs7rtxK4i
gnYMud2dOjK+YHGsr5Kf8th89yeraz1CXeosakgXDtwQEvuS/Wa/kzy8OxG+GpTn
GE30Bd5zHoG9BlbmAZ90p0Pv/YQ6yKaneWBX97MxSHq2fthKz2VxEzr6cfd58x+1
ZgFkans8GAeowDjxu5+fgdcq/4tBEb4EzP+2VwrNiDXJSHR4AA18EqqprJfm0PMq
sEeN+YWH6c71fN2O52cWBtZWIaoiHxqUqsG3CKU/dpPTzJjNCD/Tlk4OWKAoV9ag
uxccpowYku23/FsYRvlhwooT8Dq2qSSuoW4ES7O9U6iOFt8l5OhO9IhgatlNci7i
FN3m/43GaXicLcC+Nn8yH/NNpGkfFUkTFl5fENwsz5tFNVY4r9LE/hZnHLJgjOEX
aS1aUsr0RbQVPB8KtFRDqvKi9sQWHUdpI+RjSUF4v1fFkavvJtTLZc64tBl2a0xE
eu02q7XHDQv1cyYwCXs/bPplh5reQJTml7dunzzRgb7kBIJTw4UEXc4eER7XLZLw
JX3f6lGon2tkdhpMZJBMNZFXVzr2becpdMmrGJvuXAm/lHvH1v5CRt2i1EQz7exu
NDFpEuHjHcBkTFiFi3LtYQbI3i1IsBXJD4Gk+alMNd6TqxJxzvnQT4Lf/s7/NAZN
aIspkBCm428HShieRCvAFERh9L5C3jbO3Ce1EegkRDpHYbgoFEeuMpCeOfubJ8dL
1E9Po+P7vR1LxKM3Q7/uS0ahcwb2ytGlWSolTx/mYgSNFBeS96XfOz9le8Br2pCG
G2e8YH6SCYOul8RtiH2/5p8yYHXApI/C9TI8mtU+AoGaqZqmsy4PJBWq2chmOd6U
aGas+JNyuT4mp6W59Cq9zAJ2ne4CfuoRkgocfs6ha5aKUR6w4rfsPgLpoCkHuEjR
MqZWmIFCitxHScQ+nHj76oSIyG/ypX18jl6m8dyUbZTycj3kOCqmxIoPus8Rte4V
bFKRFCCQwgycmTIEYGlmQmzljbTihFi9d17B+2zV67fL0cSJ3J83EFpeo2cWOfmV
2CZC9bgrG8rXRLu+u+eWQTQbaaYzKKPmhrIMzl+0sysSuFwVe0txBaU5aiABakgA
JJ+JNC+OuV1iUEW6q127hGzm9FrUje9mYdJffq1XO1MJTMzqPNwbwA2TSeMpyRP9
jb07NBO6cs8mcnxqt0qJziP3Er7C/D4lNKKkKbuOb9VtrHZdDsbNP3UkmYZdzONB
JMXnVuMzZBopv4wZmhJqZzkvZI+ZSPNkF+4mMGdRzM9QYDm5jQaahgsTvDuxkA0m
ZpBP/7r6vBhNQvIkHjIGaoH5ZOKDJzyiB6MrPiwK5LewoFppDcOA8zqukvJLKa5W
REsSKBjCSvvtPV8aZpHMQaCzYb1ORwIrbMudKjQh9Ahm9SYimsedrpoNABqEJyW1
T12yZ0p9raEMUoaahl/gKNSEWYYFNRmFgS7x11qYPtsFHBGnxq/+MhIO7+1AMduP
v5XRc5C3yV4F8opTFLhnFIKaAQ+evWsRXXLMZ/j6b2bX2GRnTf84kjsWV/Q1WOKg
ksimgwazb+CLSeKfAlOgWrGO9L00DafZ1ZpmozR9nTTG/4FfNhVOc/oJIfJB3ftD
7fmg0aTE2gnGHhr0fKHEfyIajR+gCGuqCaQKhlMFDb6HuAyBD3SrKGQ2/bou++RS
bZx7QxaAp9sP9PqphnXUwIXA6Y+94o42ZdHiklXGKbxaeDilLg6owf/+oXBH9Vu4
icLda82003EhFEcT0mVcFXTwGySRYCa5rdrzU5Iy5NRLCuSAT1sgH8JCsPZ/WZfx
85M1VsxFtT/IAMxa6sRNoGO7C2D+HYFyC0eUnZUendOnLqR1XrZDspSRvA048gYr
MHpgaj0KOhEXJjDLGcJAnnkACwaVgqjNZZ9naJb+dZRjFv/WrZof3jc58hMPgl6j
rBvoJ90pr52C8S1KCa9XEvEx88ugI2dbR+wvP1B2A8X+AogxEpg/4KAwFWWUdwJu
/GwcxpwMbJ3b1jr7nj4fmuDSfBUvc86DzA+i4n3eB4gqDuKSUiJJro9tktoWPoQD
B94EXxTNDomMpBpa+h5+ITv1t7ogHjIq/9aop1HBtoUc8V5+S/DiJ9IrH2duRzn4
oc/vZOI86DwnGhI8bkKmVBH61y8SAUoNSoOGhYNW2RVa+566lDwPqAWhXk7mLGwX
RWZFaBXaPQP3KTWrQfuM/Ma8T39+n3CVM0G5MDXljuMHdUX+3cPnkVqShJqbLubI
3r+g/acWoWPXAntwQUDgwU5+Geei4A1PfPFSlt/hQKNdp0fhYpQLt6aDQvlf0CVC
GuUlkY0uAqyL+u1/fzSnm48pvz+InwA+U2nRk8rWrqLbQvon3cXRfPA0Gv53RdWw
hIqsfDBtkp5xh0uS4p4Iet2d3BIo0+svOgUkASKX7/1PoMERnBb4IQQtG2Os1c2P
IM0QK5cnUNUVIKjZeb3ddwQGLUPuNSl9Tm5PmJxpfqxLW1mUAtwu1m3Kk07ll7Zs
TBJ9QYbyxnzp5fDMEZKPASabhy0QJ2ZR7h12No2Gt7o5Nk8AM2Rxc8mr2ve8ngPA
9x6ZnYFvBD5SBEcqHdSMJxdGZ1joUmaF8vwxJ4rPIBdy8uWLd8V16zsld2XTFPn6
TO3tQEc/wC4wsaqZcEGYfVMhd8lPIyb539QJgNurcFhlaiYa6HfQgHCoZjeKGRxx
EEssEvgIX4dBeyZbMPk+21baU1TFqiYyV4M2atPmoFuux94KPPMvPDhzT4mOt2Hw
3yNMzNLx2JK+XYgVTRtZthEYF/ixySVOb23Rr5owzBOvk5ns3Lkc9zR4EvFJEySt
rE8wPQSPRMyms13h0kV0lXlG95/j+vJKyd8ifizYp9Jq/ymYe5L3ZCXOk9NAulok
3HFfO2O7bZGDBmafIsZfrf/g0FvnsVkoiQhTkW4Dg0YUwiKYnGLqwVNa2fWf0jzY
9wipm1YFV0Q1raY9XZ7roAdV5V1m08kpnKgkZ5F1GZv2FqvbptfZZuIZ1YFQl/WA
BBiSnjUH3lxfkBdPekQxhpUTYVo2isL7MkCa1wpdA6+eIatO5MnDWCDj9IRU1GAj
4wISvTjg8Iy02L96WSFUd9vFQ9SMn+09xoAfDYmOwBeOTWKGgGesbA2qXCNESiY7
//ksJkyNy81bLMotjllispy+M6BU1i9A8EoP8YXZvXu0hVMYazS9JfbmjaxX94AY
RF7UU9vaWK46yCRpXtlhKYC1qMosMgn91rpCKB4NfNm+Tmzf+ia6TGfiwgQ+WtjU
x3Dhu43MqvTTqxW0pW09LiGZCYypSX6nA7IHVMjUMiUm+7y392yo9M595C3DuaNx
a6+5GO0HD1zIRC04a2f1sepJs3fZEAHniHc43wjvYBr+uLHIsiIGtxwUMDdzlKAO
qGKvulWQXjeE2mrsJhJA30mbFxgcgnuMpZpexqIVYDEXPA/K08u2PcCled4c+FZ5
9klr4K4ygJyhu92btl1wC2pTVnl9G3is/fXEsV1p3tQU+tIbLI0epZl2bFTwUd1H
JXFJWhZ41y9aV46l40HEC7I+IOfCw4fEQLS4LN8rwyNVeNW/IhYx3GvGBcE/kqTy
lKCg9L0ydi76nKAI3PI/P6D+MrojrqpaIP1fxwF/BRutnNSiZ32KR6Xp4V+/7Hp2
ohjkAehE4dPyDYZr+W1AynaVw6uep7PZanXBacjpGsvkcLu3SwmhBkny6FNc7K6p
F6HxXBOC75CLiSjCGx2xqOh4QznBrbriPRs6jAkIgYkgOBhOWrjPARnOYClFi7ey
c0p/fjD+r3SQHL2ZDLH20bJPm3po2VTAs66ThlF65V9jgBxH0oMqpruefOz4ZHco
K8JJSrNUsTus2CMaxfyNmAOCCN9lH0qc1J57FUos9iksSXAnBW25IDpwLc09GVqV
g/jJy7TMSV7Lp912KISfQdeC7tL4QViE9fgkMH0F+w6WocwdsL9P739w0uW0M+c9
R0EjBiaWFyMz1HTRWf+SCy7950WINKMhafNKhWKguhBVkCoLIn6EWKf04uap9f+f
RvryoJ0HR9LOmwgCv0aDe7/0ZLz4tAfhFRkdzb+3w28sYKtkB9Nl473cNG3lPMMT
/gOMYvTFwh1s+g9h+1XchcHhAdkMopGnuH9kmimKoaYhb7j8SSX/op2SLqhZFhCz
tZDyG9TPHeTF/jiXl2P4OTQ28NJbvDlxiYsyUn8ynORf0nxn/g/wHjfN6GKehU5f
7OI7dc4oqYXExhzMTEQEXxybAdwbnXpZbSBCxINsqwPN8HeuvGQ9bqtD4lAiG4XR
2sAF6FhpEgq1sjJtDDc/NgRRB9dPocg0tqEtg3xIAoS86hWPshW214hHNTR4ApPN
ZzRPwyBhhxZv2yL7Yr+BGQnaW31mRdRGd1xd/PDGQBtYcgbLok5xRq06Y/DG2yyp
m7zAs2uD2J/uLR0OLt3eP8+Uhn4wLA1vOauY/riPcwV5eLToGQCcD9Qedsspfsly
B32JVY1E5bungNDYPaBbl9Qaj6pXtcLx0JgZiIsGsQ9A07XropordDCIqRPcdxDI
JYsZ5Xo3p8PzEaCmfOggEwUQRQ6OZMgQzgtLSC5bp3KECUcCDjUZKvB+P2nudEW0
mHMNnrOdmlETYXLggxLz7DeV1NDU5GRLGdDc6+tUHW3JIQMQLWsA1XF7v5qbvwJF
1rACLjjbeIQjMXqzkZXfCaMzlnQPYmpfdJ43+D1o9mckZGHwUTSE4ZNyTXkPsu4a
h+2BqIEgKaaurNBph313GkZKTk1fUfr6Be19lGV5UILNQk7iwQkzxGlKRaKLhTCN
drr8DrPAjq+6YgGjSANn1X9Ay888NvPcZOmZXHnwOTik7R4mGmMlOg730FHu3II2
t8f1jOtyf52S+kgd//w7irq07InSV8EYr72KKy96UoSXqFEXzYADq2wl2saYxDNu
xFFnMaeN30BK0flfyabrj0EUsLINb4Mfv1BWH68YiYP7TLT22XLnffvcdSzqUZOK
vedGU3hvI1LuIolbzv6RY6FVlX3vkcyGIuZlq6yAAj0Z3hPLo5uad/HGOFVJzD7b
fY3KwaOtUIJAYvLoxED1Z1uIntJfSncK44DTsgfUxFvIxoSPqse0Jv/qCQmmGx5c
g+b3mrlpv2wLxp7arSz6KffWg1ob0ALm4otbVKPa0x/K9sD89ZJVY2j9E9kwY5fv
qByiG3Qr2OZUCYgD/y+HEM+zGJMYEOpv4Vp/PrLtLBRmDR+UqVGkmrkU8ryKYZHB
guCColhibeC480p05YUOafyrJu6OSkJk3mjcqCNFwnHpmsGcyrfYdT05AMZVDE8g
8O1CFRpRx3tdcBpIy54YdvqThs2m2L/jTp/BXS4U+WuLal3LiXqPQj04bkG7v4/k
5RijvVsLqo07tmoi4SNRYDxrQSkl/3yL4KuTSI4uevS7az1WhQiFCtbN4AVybJBq
iYf226RyInyBRdE0wIkm+nkGiyksMzv+0meiJ6bM+zbkG7P/AlUD2ru730IiYMXj
G14YbHNeClamIIq2hRDU5RrbEuN4r10F0LIT0sdegnqIa261m38f/Rthcfj1Tdi/
rx/y3DkJJJoQBJ4PIAVwTvW4Atv8fufZDebzb8nKqiVFOK6204u+TZpw2bgXhu0W
TlUgwRLCMol8qu8lYqqQpAEpcu+eqUIsyKqO9HhMTUJEksiE/wQcEaMP4R9O5wb4
dcXSaX6G1O3LBBQ3OFrfzBLE7Qumz2Im7/LS/meBwFHq/z9AcgjMiZ1OZxZyX7L4
rGgvCOIjuCVyEm32e3jR4xft2DTqPgP//yAQjJ29ivsQ4kV1j9czgXTH6JmD8i5c
Xun52BR/87OmT0JHPzeGRBntTf+PYLXqFk5f02i/Cl/2W8UW0oWVN4TV9ztskJ4P
5oqr8EZB3foWr37+85ecYlkjrOg0ERPOPVu9hm9s25oQWK7mAMJYNJKbDJApf/JX
mf1upxMNu661iagmQjZXllBJZzIhLhe7G+TrOG7brvLKSlCBGKwzktQZi72BnYIo
kFaHOD2kMEUfJ70eX9ffxu1fss1ZSAcD5fcBZdvI9gpy9rmf2eGe5e1CFt4iGqfr
LQpNmuyAsfsZUFKLc82ydL9M9/AU+BTHp4ZGo0sj3aiT68kEiUpIOXB314NQyeeZ
rA48Wa9UeZvn0xmNcXRCl/2OB2DCuwBb5uwX1lV3wMslFlIYOsNVVsMYbt3086ws
q5XpSWm916ZcZ5HLeqAvGkxKF0WMfQlbeS7KncVemg/B0nEHFZkBB/5eViWgY89b
XtUimA7JNq7avfWwXMw9zAx+T9y6fs6LIUf3Ryp1n0S33H/EwMvM9bS6VLemO2w2
oQ4CvD5oqv29ZueO5hTsP12wkmOUWLRq/4Tto8GxRrELSYZLL9vdoE454yHLpgJR
1QOJvnLUFf5sviArMlSzkKk8kWQhv8oZ+PquQOvKRsQrnngnBNaxEir8zaJyMs6F
JcH2fRkDTCSPqcvCtdKwJ7kesYgO+o2r3YCuCa1isMEJ+2rtiwjNlJn5I22SqpHg
rFQay4/fsSRIy6xvsXrLyNWMRd26/hv0KeGMy3mZkQ2MhkzSHdHd7n9ZKw2+bsWB
yhFQWBiErqTvelM109OFRtG41zgmhH6LDcqxAcoDoJqUn1GbroJSIoj/SmLegRkn
FI7t8bSiIanu50AGzhV2pBg8yzQw+I8WoqukqPIBPufM1cVSoOBJ9m0X1MW9V9iM
D7+7g9X4vS5/sVPptGG2dNPxUwAw3Mt+aqAD1jxAt18ZTJcmd3JjukgwN9GgI2uN
xn5ag2JIVnNQXdgHyyZ6pFXcolP277Qed/vrzxFBo176Xw4MhASiIPnfgZrEUOMd
WlZcrwFzrZygNN1OjeHfkY44INFXpJCnBa/ObpW/CMSzPYV79ecxw4KdaFlhKfel
NO5n2gmSpbAmWrzdupASWzlKPRn3ORY0U4wQGTijxOsMmVwx38OfDJMwX72PrOMf
sWAxD6I3N2CmPdpBX55euCM46K7wZ2+2yqdjJ+xQ9zMk19kSCoYl6jjhVrUCyJmz
aQArF2/rGocHWudrMIexNIJwZ/M8nPu6MB+Ca1hXlVtZlwo4wmxSpl8JCjmj3KxV
hUeVt6tM6/h0Ky3j/gyyy02Y5KyI6oDP8f22jv4jZw2Zzbd3v+CADaWlYdTEeT5R
h7Y0QG8XkRQ95+QSZaG9TPXe0P1rWEtM9H3D8PPPwIBClX0ty+mQ1GpOOPjeB+fB
vALmLj7VHwYAZm8u2nRdBV/c+T/pCi08MM6Vn45m1tCqrC1okF5+2/zAvpUQdK9a
gFmSRu1PxNGG3fAxAtPNoPOfuq+meaYieEa97zAx7+PdJrQPbekgJubG60z7cmFw
cf5oOyADkhJETE6l6IxZqYHfdk9lJaAmRVqk3c3Nd9xE7g9cB22nnk51AjE/bsXo
xxl5B6M5IMaYe7ihSwXNJJAVV4jScB/Dl9fet6MB2DO2lu7uJUQdUUUT+2seQZv2
uZzhhtKlvCjhrM/TnRXhl8HqQ7c6kxmkmGKdspVSfa0ixe0Gm5Xr9eSAZ/bM88UE
QqmLt0jxMPt55NIHjOJF5JX3+w5rPKMX3GTud16XQ1xBJyQiVjjreOShBbdD7HsP
ckj6XracLFu7qh+RWneLuzuUg4KypBtfPpLZRpC0NlYFk7MVkt5ozc68z6EyapEs
FfnG541PRtB+1VE2hiVt2NYWZSe5a1/KxbrCip7MZicMLxwoElleUbWAyt9TnumL
xjJ3H/+DULsMxbBSrEuRfkTqpXfEpX0bFiVnSNhNdhjnsvjxpwfC7aZXvYYaqUiq
WQNaeHvgZDHgL5soSB9QKHi3pBxFVrJk9jCKGLcq2skorj8M+A0WpzpYnQ2OpBJ7
oAWuBRU/GsSZKeUqfOZYMLmjaj3MXzEP99iBLwu0JRCtaccZdUdt058f0XK2xmYg
0u2ZI0FkIw7xQtRlnaDI/HxCL2fbcZOQSUoNcUOu6AhdPsG3S3h/j+wmYLKqF4Qi
+FslmA1O9+uH4QhDOuKwqiq4uVgyER3vSBZq9lEWOWDAafk6NZdnHBRt9kEAsdD8
5Yqv0J6SqEbuep1fi64K9j+0KuEDdFPV7vcsIdrZdyoiUpI32DzCdMjl1DJvkZu2
7muyC1THUxSkB/DyfhDtiUkUGgkboORDxI4pvgCw4ctD3SDSD5SzwvZcrgY1JF+z
AInfuRKLMp3lzggxvJHUrSVO2hcL6GjIZ/3jMDgl7kdVu1gkny2VUFK4YZpKG7cA
2bd/Xz1hA8PeMkSx2wNfn4nTtyXFpuSsMHvceIcvCCj2ZH2kUSG2yCSggAf1GFIn
oV5Iv9ECkP/LLDCnr0XOmIahqg/YBHZj2yRhm4BSJQpCz6LGi+Mui1PKZ98mjG43
hs7UTuj10joNPMC/mXLt14V6CRH4SbaYAdrjKI07xhpQ8nOcKw1+e3R+25Vu5v3a
uawUnTHntP5uIg8h2MjOt6LCB8Ztd8vEVw9eNt6E2NEBjv2gcRC8qf4qAAHK6PuR
0/PLhOx5gAua7P9lJz3Qcp6XKKcyQcuZvQXgjS5bZkknQDBHdZu/pviPD1g3UjS0
IG+ElMxUWJwkSLj+LqKnT/ZagoLuyHghJwjeqAoc+FUsRZpYfXPQIir0IwvLTT/q
EAEPhJkjzovxczU1V40SYATsDiT9WamCaXzNC3I+PGlRuQEog/0Mb4nW7ggE6901
BfACZX6fBn5zoLic1FX24912U9HO9/azF2g9kDYaKabu4XHWNJdPct+j8xxUfTci
yIAW68nxRi1Imo22/EKsYjVbviiTfCGqlpF5a/yMYUK13fJHgJeeQrA3AN2KYebP
rooelRPAuqDDIkI4WJxHSjcHYeNOXqlI8Ni1xoWnBrdjsHA6UrTZtDoLqkt5nD67
P7l6U5z5bpAaS3YYFy+olg73HlMqWIiBGtTRPISiXxMQ+Gc9nLAewvIwbno2+SWd
nIaCGuKmcbrPVmajviAhTaZHDlJDhFzF3FEU8v8mEkcnyXDNN+FEOAdNzOBbzhYn
LFMg3iQPrbrl6HlKsmloSL87Vjk6j+Y3KVOTghzxwkem0bYp2iTZpSQNm3CvekN1
rEz+srAyUPWCtkZfjjOpT15KbuBtlZ1UJ3xLbWcUbpCKsWxoGptnMqHa2RJ/WThs
PSsIBixCRM/F94/DB+eQ18dG7UF0CahUZW5q4EM1CI1j3/qossalH6aGKaQQzPGx
kkjT6F9sHTTvnC7nAAL07vEmqTVtdt8SIpOJnLvEhjFQgj8MKyf+yqdy2B6ccu7L
hroc7Gf7n7zoOi8zW1BJata0YghTXB2TTqqsSk7OPRVTna6GhduYcBrG0ejDxtHL
ArLQcce4eJw6FMfvMWWfiC0KlmZgTbS1z9nQ/+IIZ+49YKDqpmSPiWycfFlJbSyb
9eSf0FNkaZ37mQ9RUaS/fuJDuwXfdP4ixgvczU2X6182lj5mtPrgq4qaXgGxoMzU
oIzgYsYMyZg6nuf+k6lMUQ2bomWe6DT4jymjsjRdgNxZH0rRGQaB5izqpUhyYNB5
bFHpSSb6/PYFa5zmsPy0OVIFzTFklMFoPWtRxuAHHxbzWLebLeo2zqjnyeL2IAgh
s6upQE+4U9uiLhdizGfuRc/rxBcRDlhJMll2+q7JCGv+12fJQz9TLToHDiWHR0hs
bw01eDyHOicCk7WKYx/U6nBXka2JNklf+xuXOnOSuYQcysX05A6z8db3qn7OnlnA
CkGfNF7NOTXtoQ/G5mB2WIcD8yYU/2Ddf54xgk8J7pdbIxfmagHPUjs5+iylt9MW
eSa7t50UThD5GcGLT4crNgceglLpuUfQ0eOCzL8rGLXyUQa53LuyFnLXf6S8k8Lm
Hw89gBza5DnOs5D+oFkBJh/wkzk0WQ5pPsXXOLNoPeqacklCrWpLWzuj1PavpViW
nuKMfboPuZI2lijh6W7OtxqE1xi3RK4XSUAGo4BEPXFrZncagBSquhN7aNwmmG6D
hFpihxfLzRNNX+ybEOkTcV8fh0rhFaSL9TvMjnX0jwcxqIugVF2bwMIHCIxPv/kV
h+9kzKNkM99Wv7CO16/7rXE8RHgD6dHJ+GtY3sGa4Ipvnjv8ZFT/foIXX+4oGrP2
SZf4urErpjeGKNiOx5pqPTuG5dzfjps1IUjkqYV3WofQz+vrtXzS32+4CMlEJ3qk
Txpibw5ty+BFKfu35oLIwogEHfOulDw8VVz+etHctF3ccaCIB1XrFu4R2xUDdRyM
/hRWxnUBUWAkzQz8BbNAGGWAmrNxy/vrNPGX4k4mnbNvcEMBAkluydQXEdh6Naw7
VWtvbmipEp/SarGvtN2t4VVNnNtNqMCCzw/gi2KkV+CpVvnOQOSmdLhRH4EUNRvE
aOvGzhWLrYUy38qiYCy4lGDHnyOt1dqvgO6eGc3xOmmMNSULVXrht8r3Hj/FsKXj
znEt87lMV7Lz0lN+ykfyo57Oncquq0Aeus05MfAlw690juPjRwblpvZQVvl2BlJs
s7JMkQRUuV6tCiQCzUkAGdfnSkakd8fnPe3CvbSGRI6ySLW7TnxbU0PqxPGtw8j8
K4DStJRh7EW9pJWTz2LFuYm3ua246fgT5ZFfjaapFawwKEM5rq+zIv2EJ0zD9tjm
NOzYqJLawtqIK1S3b65V3ANxzpmKFmJH2rQhwYijO/7ON3HmLUxxbgmJeUNNJBml
oknbr+8p5uFt5oOC7ao25GiNmU6nY+h2s0DulxheykFrXQFhJh94oAqTxVzngYng
UXTA51Kodz+rKDwpb9JmfeDGOKA/4VzpUWR11eBVzjuvznalQeIKZEtTXChfG1ZN
bHnFqRN5fsKkPlRe9O6ye04idnHBVX7T+ERB5KkrF/pciQas4TqUQKXddl9FV5YT
MjJEXrqABJr2RC3xUPhmgPoMSbFreaC50st2Gmj5mATssyZM8CQXfLnjms5cGSDd
gb5dOU2HD3ZVtYgowOaenQfb5TeiaL0Dt3Je50h+nLYsE/nn7MFPvvHhZ2Y3aYTX
3fxI6HpE8EATWeO8DQXufWLz5fXxyVDz7D94zI1lB0ShJDjhNTzQQqufBDggUZ33
VaaAdItAkte6G4I4G/abiRDoThjcGk/KJ9xZE14a1pIFc8r7BeYxYBDkYnaFkpDM
ZlR3avh8dOkmnUqcMF1w3ir29hD2C69X+BwSMPi44NZWKvEr/GthFoLm9bCxTB/8
ABGG+s2efst+92WPz6VoYlHZuLE2MMNgksdczTuFp6/HFYHma2e7rS1ILGa4u6ss
rDcRoL3aX/GaNniE4EUuym/cyoqXmrnEr7dTPv2UE3NdC7M//sbj71p2VVlKi+er
MKYCFMFmibyRlxPtBBlgakBMt+qgdrBqyzLQWutDcTDljdNZbkCUTN/LUMc5/kvR
5pBsKkq5XBC1q/I9xBg9zkvRRar+6OIoYo0HO/NB+dO3Q5IaXDLBVSw1T1jJUPR4
ZHZUgxSMzV5DTr2dbzrUEMS5bjaz5O/cVaVNGQAyOUoupQquS3+ocagh6hqUj2IA
C/A5LBmJ9ys799Y70YgWMgOb6kkQV+uoEKHIL2jdWHLuLK7pyu2Igul0WP1V/NlM
82CMc2UWUEqI+QFcDDfsZKsXyLi48E/djpE18tGBq4DXYHcCKSaezdeZ3k4hejEN
FJDRknOIMv5nC4QOBjMR42QGzYEAHIqiYYdhnFegdO6ArZniZqvTWMQgVYyyj6Fv
z3CwEPSSwqDShK/sszc/Gd80R6er4y0rpF/UazPHVRcxUr9sdW0A0RQ6SF+Fbwxg
dXohljDuKK8AhD8tMckVz6iKpJzMtPXXS5dQTOCOIvFGdjXs6d9/fx9yKDwjXfUZ
nwPMw+35KM8ZeUvtO/Tj1XgWfp6RKA3RMNjpMsMQy3utUCPWVYGkjpi0vENOH4ug
bPgqcl1Lqqxjxr4rgWf4EM8MO7ilStFQjmDCOWx86wC1rWeoOwI2Jxs8o5T6WeC0
0T0X3qJfZ5Op1tJ1Q4dhQCWnQ8kDwoMFESwOLy/VgAM2QfpOjrsORFUjSQnL07Sc
7nZN6fAlVoXUi9kA3MM7iGSrka/2hS+IGCjWq6tp4diQ+HtJDfwH1yz1Vho/OsC8
gBXlyNmRkiB04UkBuWKAOhuQUAjoHLBsB5uOmLqUMI/OeawohNWZYrxixxEoC4p/
nnZsVCE3OZpxwaCwGvt0bEwSnUXH387i9YGxAursbsgFFr7+KE+Ja4TJnv/stiOl
g5Z/Dij4m486CAsUVFPQuwGF2fK7yaphOUe8z5LuffrUeTiH4qSfzTB4pJIhiiN7
0Kjuw/dVZ59Kl+/vckMw06XObQF3b/Ct7Bh9wOsTND8hHeIb7lhp+VqrwyON5iTL
EhxfjzDsYZsGZC2g14inoVQwqryY0xJAJaUbSbAl/hbBcBHp22XZB02bGo1E0UEJ
9/iPS9k0fqHKRBqxajA38+kx3Goibhix8AvIoIXUVQ5KVV0yQMQZcIeEWkBHGIBG
fksIG7czpmUxgwrNE8QvI1KYIiFhMleRL56VYk+S9Xp16bAphVlp7qzTHB4SlY+J
TVpf3o8uhY+pf+fLKFXP2Ovs/tWHw2DslYee4+VtgpQwuD23priKhAJO7cjfRwG2
edCLgPrZmefg3UE1H479Wj8cJQxrTt9c+9FKh0MASGmwLnMIN/OTXEBZa4GWPNkn
Qr+KUQ5/j9f74REQqDIgPFAOqPODZLxsJ3DhwSIwZQFi1VYkvchsMskrprNZinVc
HMu/t65mY5+WqstznCykuPRv3B+9Smipwnulco6wiO8lC4UsViEYa7gFu7XvHxaO
ImlffI+00fqjJMVtT41b0pBaQFmz3Pgn1EYmK2Vsfcwa9rlkWxuA51yPJi1kC9iu
WGhYMli2NxshLZEG3s6Td27O0WW/r3JTGrXnvDxd306Sr5xPha8jI08ZXMV1Fsb0
rRdo4aYxKyeiqAndkBPg16y9HsTijz4Xs5UhK6QBFlCcBCPcDpw+tAc5uiREOkI/
m6h4gmOSuYmgirNZyBPqgQFIeqGegT4bu4yIEEph0BdmWvp1UhcO6OqImQKeHVHh
AchZ5BtYZ4v767pp4ftPOJ2qXnE03PKgolNdgdVq4xkPEP2T5iBEy5k/UD8oMZIF
5XyBWGtW8mVO0pFXWLEzJ+ipLtBOhiE9bSnEtO2Iwp1K4k2F/GrIl9BOF88znXCk
X6d7k0uFD7OdOaqk5eawEy4TnuJUFDdzWsu2JdLSpw/hprPLVDAcHfmjqfV4WiFj
9xl0yOPt3drOSjibJQYhWe9LLgaM9tTOxzY1CZMBFsSLafaD+L8O9RVRcGq0amuh
D8ivxO0ZbYoph2b1P02DCcQ3at6XAe6mGDG1SUEk2zRwChjKIjBx0tx33IOc0YKi
V3mZ2c7hh/v1zadLNV3mHTJOh09x29b/l6Gc06Yqsjwz8cxR/E1Q4U+jF4urnUfo
5wH75HFsi3ZcZ+KDT0//AECwVTwTtuDRCdc4XtIjmvFCLeMnUO8WqqoS2WNGi1LD
K0RNh6XMdjlJqHk41cnf7XKx3kyW8TccQ1fWThCiV/T/ChjtxqMAPByblfcLYnlg
22jVk3IAe5nbFe1fV8tbATGePGuACDmv+7Xd9laCNGc+Aw7i5G7BGyS9LBRjyikp
+j2GnbN31UYqxxt9WEtKKx2MyYCkmdI1+m/I0SV+5iQ2us0sxbmJ5caAs9ZvHO+a
rNRCStn1qfpnO83zy+kGTTNC27NU+B/V93HI79wJr8p52+cJhvrb+WkoITu2oH/v
TdzXuJ70xvL5NNKCXk69XgSV38Ge+eWc3K0z2eHY3o1vMJ+sAPHJWPWvV11xrlVy
YhDeiPXs8B7TjN+ZuI0wgtbMVscXAMHqk6eJYMSrKTZIlvcrr+YU/sX7Hiikj1ia
Bisb8ZHh03eu9GZPRjf4ulzkNiOj+6vkn8MVCN4jfM9JBnFa6OYXB8Vays8m3oE3
qAxd5a+X57M9wKsyDW9ZHPmjsfPIFB9a90H5qac2TW4f/yU5vPge12F4b0L+lORn
1icP8rEvT+MFEw76nz5w4igwY9Ycq6xOhS3SD82+0fv5C1Bon3SqnXrt2wnXAwWI
15MIUPNMWA9mNztlK7VaubWnPQs7eAhGPn/9k29/LuPqw+5dlbyyYvcF6oyQvmTZ
R8qV1/Fycl+B2efd3Z3UOVMsO29HiJZO1/9DwKo8B/9LJ9Cds/Xjzzffp8eee6lw
vteRPMAW+uH0/aaEmzM4ndd9zEaZ1hf6zvs9clvEC8zPfIabG/ruKxw62/zZs+d7
ogRLLYxsISWYO/j1DNCMCD+x4fGSw5F749ATkOjZM54mlStiT8Vq9kl3w7Tvi0fQ
7yONr3dPGd5vqd/lPwTK+5HTDjoag+0k3amsoivAv7GI2dh9KaBpTqEIK03f47fn
s+YmVMUHWImbeqxZmO+ekn2Jbl2Iaqr1/TjEx59r9dIiUSlmGQzLAvgOxcsMuuvW
53bjvUyoEyoM7u7qI09SRGHyyaqAIoDzjRE913Irzt994X5+T2xM+8o8I+zKdChH
yN1NdW5A9Trlyg3uD1dKwpnmrLNKKg4ONe02y13oFmLk2ixER64lBlonXBPvW9bg
THWeydzru/82SLs08i6YNlDNUEwrpfWFuW0gsK+9szhbXG61kIZudozGH9WCs9F9
vDI7B9Md3PCaLzpmYM3zvf4p5aUB8TVRitj7s5tFXQFGbGMFA9TfMt3g1JctWX7D
6oSl8QQ9PbSLshgPO5c6wB+LnULOz4cWgZOkqIClgYXGG5O5YYa2IKR3/TRMa9qK
VLhR8AXkeF6gzFtiVPZZQmtyeu/JjuNmZClw++FHbjf7/QHOFqnyqTpbEQO1Mi1r
rPFSNL9gWYe/e2dPHGhWLvrZZuNs1m+xPnSp+NbjXT5K2nrV35IeyRB8Dc12ZrXx
acUd4xmfRaJwUFsPDXfTTx6s/LkvWGne0TCR+OWSsH/vRpQ3bh3r6robVFoJWeaM
86qzfcEzYOgdp+RGF0eKxwSAka1Woi0qlx+gDMvArwX5j/RwLgTWSGZjlLQcj+K7
k0gpVN21iWJNS2eSnVjrLJw3hpnHEPaOC2sMEbjKK2lF0KyTtZQJxhtXhB3AR5sz
HmcjCV/GicPiTnDsaYu/tgHKpmiCNUXiN/tH7YfxHdjVkiWs2yIiNeKrH+rnK7GU
TJ+Wp/NBg4SC3PH79YVR2c5Iw+g2Uz9vJHKcLSfRATEgJhY5jUKRAt5rJvRbl3e2
GWJzqDwPOBKrWITyuvfbz2uNfurNWAHCIbbaSNR6k1sBMDWzz3aO7tRjQ6XfvV+m
rTtcRRaBxZa0ebOoLaDywMwU5s+N8eDMyNLvKkVt06YjQp+CVUfgKWVAb80/tAsD
Wvix1I/9k/AUBEBLM4EKx7r+An/Zifz+YMkUaF7JC2mIQQs077j9BggMNQJ7bqEp
eqPqAbGTSXVBOjbRpjLHTOnLjYoBpwxLZ41zkcV+ZSkC2efunHe6gkg+eYAZ+zfk
2L9XJa/DIdQbBNYiFg7vIXcukahCBuOaKEgIFuuHgcf9+DIX5XvK6yTTVotGVa8/
mBxuekIvVmT8J/3QCxHsDwwQMEzkffgscJj6hL4Z5KI+ekGOxTQGbQzVPYfaH4zu
aw9Hoy5rT+RTiBHIBNjhoht9i63EtN/7o2JkDtLcYSLaOIp+fyHP4R6H/ZDuyZeX
H2w2ez3lNj3lHSbQVMpiLbE9/4iifVO7ZWCIShcD3J5kIITtsOOMBl7q2j9qzPZG
1J5REBzkhV6+C+zjddF7t/AR+fMU6O4bT50mMM7PoNSIdo75QHn9MFbRJ2y8ATHw
iCSqiWftec49zsJ4bmoRaWbl/9bvyyNr6oQDSQulBjukBdHXQe0eqtoGKSZJT26H
UCLnZdos+EFQVe1jgt935UaTmlsOL5h68y33+lriqJ7Jl2wcV8cIONle65iGxVYl
Wrk5uoyJgkhTZlLdXMu3ExMhndqlyXiCSRFtcm0k1jw+fY3wALebAAFgpfG7BKwC
qfHGtgI1L2He8pb2hRttuOPYtYGm9juomcS4SkkPjB53/m59a4uK/tkYVY+ABFFC
l7gUaCTQDigL8l4H8Q5FgrVBkIS+bzuGuCmwl7Xy1Ij2utkHr4vuQJff7jubvFOb
SHbJmXn5y6F77tJzCBwX1P88p+RT7ek3Uq1HYQ0guunZwAnMeWz5q5vwiOLGkMtv
d6Gh8c9vajCsKitCwDKQ9yQlrnKJnPf7PgXzfufaSdJw3Jd30y0gd6VAdZB6Gj2i
m8oL1bSORJ/WVQ8RxItc3X/c2er95/IlT7E1LHCBUymjpp0265oym2xR6PNJ40L2
y2guQTPIjIk2juyq4Y+JMkknU3+otr2Cc6hsMmlb6pjb0ptOrD9covgel7SqX6Cf
/wMgnrljsdaaIUTrtGH/2BBx9fs8dC67b58EkVHFk3ckB4ON89zlR8/MS3FgSElW
vQfKIyimZFHREPQ4MqVLA4Whq6BlUylKe+p8B+OWVUsDDDnGNYe1Vl3sara2atGH
yUCMO74rkVr/ofQWzw//ttltEpfdYcuWUUPqz99kT+Fc/uQcC/9rCq3EvGhsFuNs
YEX0wEMzWciqROVp0ludARGt8jmyWi8cbQMPBV+QEJPpyvBb3AYAcsirNGHaKBBk
uSOrEkOrGorAYn5jMk7g5Fy5Vv8rAVXCWTu1xAoBNkVjZ/b46DKm6ExPIlzA+twz
MR4IJAbcoKoveMDV9W64SS7gVcXejX5CzQH/r17Z5XMXoYOWfBwcX5ZrVN2qA7Eu
8FZ6EX+Z4eYJ7pXcxFNehjHjsgWBd4A6fy9IIXyTt8gUj+WJ3r5jGGRg+J51Qn67
6H0Vx5DD7weVxKINKKcg+lfG04uMb3L6y57SOBkfgDWOvGwXg8aCwmZq/B/zlYWw
pRLiWu6vE0jgvucmWrMFdekP6kqdHYHObqLotaWeKa5bFalnJGwE97PKLgBeemko
t3W2HZbMzCgD6yeZoNnjTRpaCfONyrpx9eMI6hWkVka995ao6jIP4RwGw1kttMAf
UEhadtcJXtrPEMASjd1k/GKqRMsi8niWsZNfK607pwk8g3EUrpSGSAXj64CknOy7
gFatbiK4gsi3Wa1HzT3XwWNn/u/dy+7hlE7rnC9FZeokM6BxxsaPFacRNl1qrAne
SeJ9RHb14b73xFB8xq8fdDsIHtDsZUciPQBaw1KtR0meflO11doE4l0Fc2OFbcoY
mgl3LtFpC5XY49+03oSDJqIb1q2ESUmbFfdRziP6EZLkynQnZDtZx1tldPIyD02s
dA0XN2Q1qv5DQML7bDyOTqmMm0GLgY48jUKJwCm02FwkSqsicvqjxawdElUq+z9c
fjhVCkKUN99nxLIuHzP5aqs1Dm+Q9024B7DplzE5RZWc6cm1mCGf2f4MF1d8xJxx
zb8c9vgWiuL7WuHIvtTQf6Qbo0hTsGle+dvO0Go2dg1H/ZwAHsqbRCLiznj8mlwL
Tked7Lckm+zhKUcUZQPO19FawK2X6g1dl99HG5Xn3mbv0nbYnmQIY2S7XKb2PgFN
fB25ihgYua+va9CI33Rg/5vLGznAvrmoA6RTucsd5VR4ZRA7Oe1ohpUnR40TiLjR
lFLXrC6L8amGw0bF5RIRLRSsbAaNnAo/hKjWr93VYaDRegh8Lx7UdaPJDQmv8kHl
pg/a1KDJwMFUiuHPvVYY3P/ERsafXRzWX/+noPqumtxJTbfNZ8Of0ftEy9JcS2GY
nW9iK572b03roWgZyrRPty4na8dPMCKEyt+H54LvBjdQ5wXiCFmyXQiPGVLGAB1r
YitsWIwPQDQBgpGOzTl/+KO0RPidR6w4GCJliaqgS+XVvj8fnDEr30uA6JLBBYvk
GZvgOFH5yErGIWiB1sNS0hGn5O2uolsWKB4vV7HZjKhP3yn7IXr1VKYBBuzN/gpX
1NM+uxHdn07S1CwuXqISsbV689hyA/rugyRvWutpKBIJiCPwhXLUqjp3yXoWpMDw
BBtHjj2tYbKBLT80v1vfQoaavUooxJxgYbo9HEf8WJijXa/p3q6Cm5Xe2MCyW0g8
o6b7ui3CnUMx7uA0sqmK0jlLfI7N+meq+PPQyAk0tCWN1ybD7NlD79lOkHGSAosy
qk/zNTncq9VfnOvxG7LhAlgNE1jVx1yof5VcV530hA1Orw3ed17aqRLo4dB+w4W8
DZ3uvRTsRXciWfpXTKrcPwghByMryj9uBFbkKB4GCoWx+8pQmlMD3x7Vb/UhesFL
HwJGPzXrpMopAHG47yB5dfVKikSSK3G1z8h2S9Zki19TMrisjbBpy4kGs4fWB9OZ
jF0a0++4QoacjRNOBX+bLShSgQJMc5Jw2BKI1wusylcsRDknb/gy1UBfO4LL1WSk
aRLaybh1I5/ai/EvPPwPRZ/PBILe202tFuX9mqbebNbeCtwXGevf1vKILP4kfHg3
dMEHjTr/3xVeXfbLCn4vg60HSbhoZ0cJa3V6/2Abqx3M0cSyq8/+izp24coaG4OM
gh+GDAYSzVxg6NDzVfoWvj3/jX91qpVJxk4kKfSXsOCMb04S6IOm4YSb6dts4cx6
UeNg79nnThi1mtQluqg2EBxZVlEu+5slQ7+BBYpCOZZ6rbn3PzxhMuFSci2T6nw7
wAbEnpqWshQo8Z6+J6rS6JPT45vHzQdAdc6h05UoUQD6vHhw8iLFBVkGc+Djqdx+
gSM4ZTmWKdfTFnlELpHqdTNlNiCpsEY/BNKie0dVyi0G15a43nmiAp8MxKzAV8ha
/sdvbZOsXR2vKqPCS/cKSf9S7TqY9DCUm7StjrpgCTHTE4fIumYpBa7csEt/u/rG
mugLyOS8E9yxnqwHWJOeG1Clg+picRl338hRPb/H/xUOahumFTIjiypiwZpSKZ6t
XTDFsp4SL5H+jCMfLuoZHBlq/5NV0T2LIiimREse3TYMyxSvQ12mlNsWQTDWuQZf
SRQWFvFulT6e0q/DR3QtenuL6o9KL7mYeNu9fhp4p7pcMPGiHFcBqyc1f7k3RPXx
c2B6aBKqplqTWJHoRwwsvhMAf85xzfb7/ZvY2E3F3nH2wi3J/yQaGWx+oKPXHzHq
cdAQOsuKoTkiPsNv1uMovk1Swvkp2rF0+utbR6k7kO2RDYmniatHdlpZMFHNj/dG
n4OdehfAnkvwKIEQslFWCRUUsyiGR7wRdsz/xSAKoJYUnrrfQSVFzWDcK1GQhB8J
iBks38gY1WtANP5kMbkCha4vx4pyszMr8oeEBIEoAWbjgPdy25lK+WnOHFN56Vtp
BAGCIexDNmOK60V6iwrqeTnJIsGK+czcAR7VsegDcBP2sCp8lmWM5qv2IezPClLc
Br6Wh+/Joj8hQefJIJYlF5VDzLY6iVH7EpkQ5jxoWk7f+5fSMkHVzNvfOJCLzOrU
PKxypSIjA4aI0UG27drQOZ9suFCl3FfCTGgnfPDFA3pPQ5l5LVKwpFvVdG1zpnxV
OUiV7QaYqxyb/zJGmVurdy+7LlUkXbPaFOUUUnda7F5eHDEr9a+JbbEzRTbRVIJ6
ratltFrxwfTGKNPrlB4ASkH86zoWSiGSukLgNBsWHKiniodvpmet4GK6rgYl3uGQ
XQy25cLwSosPDo54o8ZFfl31gcXA2KxOqDFKUmqXy1Z8vg+/RF/0RLj5TjWAX3kn
FH05ldDkxg72i9cwZ1gBUoQKXJDwvCTJwCHJR+A44kxpnqkxjYXKiwvKzlKg8ROK
K1VbGclmneBpF0hH02IQLajO7VkMz0xrX8+f0BchQ1o7youxp0tai0arJgwKbxgb
JIftujTcvrK9IvuKJxPT5Y/2XMKoT5wBmLhWZnGeigBJlSmR29eSeLZ+71Qj0Rwb
GAguKPO6cQdggC+LdaOVPcLPgKNu9ImWZ7Tdhxj8x4r/P8b96GyN1z+OoMGmHuWy
Ln/OqDESqTZqZAuIofT53PioiTcDUYkVD67Czon21y0GAh8K3BEBlQ6sO7ITb8Cf
H6QyiIx0NljZTbXTlsnB66yl8V7wiLiwTCBdDnYcg4Chn+64GSugU2ESGAHHgLDd
Ep6r4nHoWC9luPF9IPilG7KGj40nVwDabXy1Yh71tqTflgG9OxWyC5NtU4rm/hco
JQ+DAo2tlJ6MdDNKFYh4dVlsNkIu1g3oOE5S3WvfowG09nfSarAnQljw6QmbmDwy
bjHLkKWrhcob73CCxn6MEHiU7NkE9yr1btIYLzibK8dN2MOCVHOju/38QCHYr/ME
n4QKIrK5nOv0kT5hxcp4XEwh4779EuIFiAqQxJApKKv1tkW55meBz+y4fhK7661V
bu7KbPd/5FktJYfGa5qXmtb+ppLj46QbTtAcEpGhtMvJyVk5P+SCsdRdxCgZzPJ9
lnkyOASYmqu68/fqnZraROD7jM630J1KTx9iof9lblMMttxMdTRdoMZuoEH5h6ve
PObP/sWQlBlhj1FiIgmeCe/IVSeWI6ccXwXvWEtXLW6l6xkawt86Jrtdl9ankHrC
8LcEX4V28uYlV4cw1i65LHA5uXDD/sHqBMPNWTEicqQexjuSPUcgyeQQ4UJw22+4
9JyYE/E0OY/4dlEmfBU1OvrsUOFs48YhIMsBKok5ceM3MBDTyzvWvmW3xXl1eKtU
A4hJk16OnBvq7vY+FGoAMRYerFjSDMi4BA+k/1HzG0I3zBiy/t1lBjiH2ETIPpp0
BYtw7Ho7+PhgJkH7xOG2PFt/6UD2FMOdccLg7GJfgGRzrK+nH0ijYNnKMN2yWAoz
8t2AikpwHJ+A2OTflR82hId7z0AgU74/KzWfxjVSsMWL+lCMYJmeLi040zgGyNPs
oTBiVTIXJWUy4nGSIc01OOEnUHKh7fx9wkqTIWjttghZxEUswzP5kUInPHNeDCca
qcx1/a63sEbfiRfEPflRxjjLov3pJYZZ2Ybt0TLYlKj9nPS54vFZh+tTBCFMIaxW
H3dm8s50XB+RaNHu0qUA8kIovaxxg3mXe8GbayetDcUWzYxHx02tI6sCUFpdgrqG
8fgYuLIvz4vaLaJLjgkppSnvAOATQ8In5rg/suLin6qi977Id6e8ZZm/VUIKv3LJ
e7gH/guKbeZUK/5Upxp6W/Xc5efqrCCr3q3vE9yApdoH7JJR4ebhsxYr7UiYbo58
rBTs3QTuLCNe1GIGKOoyANv6vzV1Z6kHx1L/uI8qIy9DVA9uGpPVrtmOL+ajVGvu
ZoQyq9rKf1MM0npDv5WEsB1qPNaJMWf8GO7At6cFox28zNyiUKgg44Dm05gqW+lw
iHXY9znbs8xiiVX0w8kpbeSZ5/SUNTVlCJiSDarpz0XVZBeU3BZA3naNVpEnvYoR
+1fIUvug2gJuSTMi7W6jxOo4RDm5JdqZr6feuvrh1tH36NJ7pFollme3yIDxRzGC
LqjW74pcYGoUOh03wxJSZYHV+rfSG6oThrRx3aosRLuHkeki8tgTRHMTeJO9lvxc
mvO23TO/eMnJBi2OoB+GWQF/2AxBl7pJvI02TzkxyDIXIrtjLjUDPI120X5xTemK
UJsgyCiXkL+IkOTnWNpmX33bu5imyNULuR/WdcDKrL95z9SOZM37VbHvuu+Ix3gd
qQ6V6ZGsDYc+L3VMixHpaJXEsHd5LHb85vw+/YZf4ZN3ZIE8LijFXBpDCXIKxj8B
tLkxVTh25XsxjUCovbmsLkqPZMOz4/KvPlrhcfMjMktiumqln7zRW4l6A9u2wrqS
i7IOEfOrDubNuDPfGGOVdNJYnrlXqepeF+QWccFQy7cdY19xl41PnfPhKrXZeGpH
GzkY6Q+NA6KcuhM0yDaqjA/zmBMNT7BH7yz2a6XJKN2+52TLyICXjWqcFiBCSTre
Po/wfAwDoSzt6N7gQCPiiLUkJb+w1qxrvdwSNZh+3TOJj7RsRN/Jj65eoRiexCbm
Mob61ZCiS3NCH7bE/hSRL805fzDwvsTT9qQUT+kVSSPK1d5ARMV2J+oGbBeOce6+
6FHkuBkdrud/EkPyKokh5hNLayiz/ODvdHg2A7gRXdRO1K+NapWv0QKPHmOihEtR
AK5VCgFXtRuCv82sVFveLZ45KMzlgC/7rTdIwd8Rm20NMUktrj7/MF8+VLtBMHPQ
cMcyaQ/8ubKNqTZu5dX5fjWieu+n56ZXS7vkD/dRh9tKe0Ovg3S9AeryHIEx3LoN
O2P8waQHuyYUSQGgDLmlvlCdloPLpboEONVjbtERbd4GmzRSjpWV7OJdLmfmTAsH
SG8AKkQsuIorVh/Q3yMZ33tv1Vg0cGtWVGK6EVVhpce09o/gwUV8NE4GSsG0BhFx
mwqk5bq2VPJ4psJFc0YpyK6Yhg6a1HaTlsIMnsG1vVxczJMD267D/HLopv4Gkz3c
ll3jAvAyMUo7f+b2izm1Kj9O42IlRR/dyisGkfyF6JPfkjQxPg5uiR6xrNjxXNNN
Ka87q6WYGDR6xhEDlKIi+uelfdfGLXRUZc5x0T8t4RHve/1ffruv9gb+ChVnAVvu
1kwlTgxm2GC0D4BLZQANMEdyZhpdPAULRDDCa8tVt0O4FQOX4CDT3jt1RCA1I85M
mUOll80Q7ZS/u9XY5RdliGxX+CX9whlZRTQtbRWwO9qu5FdrifBzmZSU9LUEgg5F
/Lxy7G1GT3PgCLxI1KYEfzMLsp1iTQ7MaXbv53URxUZoSsLT1vVGshIFWHDXrBUE
VN+BD8toujm2xyEOD7BBtQl3t3R683ajKlqEjs7fK80bh52X+TDxH2VX0smzSSBT
uAZMOqpE2cl3oxZfmmNsFE+azPyFkBYbvx9LycfG2TEeiIYzPv6Xap8H4P+mkqbW
/Isu7ybmly6MkGDZ5RTqH4TqcHDqbr8y/umI1EGkoYQmQLK90+RtK/DlXzs9N+GU
ywZTEKahGavxSvYvdADn5hEu6jbrkGEgjSKKbCuNs8QcQ9JnuI99INQuA+YB1fS5
/gy6O0KERy45u38mRK6oXxn+NIT7KdYROgUPpqXVd8SsU4JD9PNMiQLcRHvZgVhx
72mUlcKsp3BH2JpL3xc82WQ/wBLI6k1YVVlq7P0EHPJX9Kn+G3+Ss8yH/xmZhrfJ
KOUNfALkaHf4nmenr4mMxON1tznYTH5YAUa3RvB+JdFhucXrTy7sJyNvlQ4mTgIU
pT4Uw8rh9x6z8q461vVtqEIkapMRPSeM6P8NR7M0UymlBAAkYOuTLp2sXL82641c
B7W2xs2y5iUtsXDQTJBI83F2SpfCGKIdhlBcT0KCU6pDleM8XFL3WqA9xugGt9BR
FY2G3XbYeuMWNQkJZqwGQd+XLS7g9XO3hNDNRZqfTfa+FPPdMRItKSBHH6cqVRwK
c87bN34g8pJfalK+Mv3CT0Nf3mw1uZbCQxi6TXzs+bn14JTecW1no1tGHmqB+qR3
CCVXAHcAPWvevfjELaWCzBFLXhfVbt5AUf7SxsblsTTlZAAXPaFWNYM3ER7NeefF
dAwqHxxOwFClJYSkBmw0/4VWSbhpLn3ou2z3aRiGp1/I2d0CGGZRwnzUTs3bNWg4
Se4EpfFVzFudJ4qwXjS7c+4RpfbzR6F/wc3K0G/98tSqwc/2crUe8OXsz/EgxzIa
kZTGC9pF3TojRG7vyoCggXcDx3yNLaTP/oQXjc+4v+7Nu7mQmluTFli+IQ3ELcnR
qAgvTrSmvi28qgw3N/UI/0m+XV0jSYLNnZUKBQSz2Cq6mL0FAL94PXmYmsrjGrYv
N3pK/U0KwSiebdBGelowOYupp2awIgGscDV4KD5jjSG0R9WQJDWv50F2EnLDLb8F
1U43s5dROgFCdIP9FG9oThEgexgCUeZ/Yn+F+A8ZuXV2zJhD8F4YPlfIz+gihrUR
XpAcBrv/7g7gUw7YDbRvNjKG4U/+WReIacYvwN7ZNuRPOPwItX/+Xn+i3pk4IX+E
LzHhB8yjfnoft3zgctyx+dsURrGNOK2sva0uXvy4To99vTRZwp0tHhhftd9GVYR4
7T2TJi3vYs9l8mprmfiZmg9p8/ro/cqotL2jzzWu7H4OdG56Kcq0iW1tbbOPoDhL
moYQjBq8apeob2a5OPI7mC/PAwWnFPWcORYbvHAZN4+H3xnf7R2IGfR5Q0GkXIhU
NciIzLbIskGTACMdU+OGNlBLu3vooEbH7xQwsDtnna9ej9MiY/w4i3HIQ89b/yKa
gR2Ba3oCsZ+MDsJWznsP3K7cU3ohIfWfoXSS6+Dlr5qgXwarijMMC/lMNO/SA0d1
qC8zs1eIf7pCd503M/+teKlDzlBBr1TNWBZV+kQL8eLEpQOkBFkrcDwEUU56cX+Y
ckr7SkM9X52DmePIKOnttstAiV5vYsjALfXoHIqelGgtaiyg3/MKDvVkM0QU5DI6
kDGTokFbCnpT82DnlDpzZYBdExDw/ci52PJalVvN78sbQrVF5R0hSdph9DKLkd4u
OhLoE9+Jq4goojiiQkinFElIAIRq9GsFBTVkl0XA72HXV8DODCDYERQ0rTqPjn+I
eCpZwGjcZL3bWSSEwl9Jt4yW3epRthlE6igxb4xfrMpaf7Ls5uzhwRmTyZXKGQzk
LZosEkgvFSgryE3Sj5Kfy1gpnB2BzQGIzquOszuZUIhnmrKSGh77qvpa7RS2FS5M
K0wtn4q1cFqHF8zdnXiIpArIQnMtG3r3hoSrEZW11+WZn4nR+/153b38RKSEqg0Z
vYb9yJqNiQ4o0c7oEGpHWmbQAIasxYKlAnFPV7olzUQMRtPerBVb2m/jRiaajYSx
mdfes0XxrQYC/40rcD4WgTTXnlzCJQ2GaXAio6bJ4fKNxcQc8pLpqKCvI+AdqQlW
eresYtIuOkp8NmATLuX/K6OJLe8OwcDlJd6/KrGn538/OhQmxOqqx9juSgkdbux7
zcbzOvb777Hsh7ExCt4R/6vAWLXYoBqivsIA/d4PAkcWZq0FHIbcF0tZ0FM5T/P0
TUe0lPcbEQl+cZ935+FwlU0KadVY4buyxQ09A1CVAEcChdZCBnX6qFAmKM0jOwYh
HJ9GQYRhSLV+v5xupbkBWB23ncgox53Kq3cWeqZjR0AXDiUlm4eXGFfb0jOeFdGT
EQUUGZNAA07FS+SbMSpSc4OdiNbkDG5KWe7yAJegckML0jO8S/UdQz9WD/hnfSgT
EOxXLLqNINPJy+3XQnuDgkNwTO1OQ4HPlDB6swk3nSiHIf5RIj6x1+XKx12MWzyW
4iyVT1MwA6iV9zfBw9vMzHM0yr0QEzO+bWwwmpDS1horsLZj+I2qsAl4p6nqOWJn
LvBew2mkMaKxd7UHI6pB9PWhhUmit14FEDTnEZqL8j5W0Oolav8APNkG5r+cxtRo
R9/OcLZntD14XZj+6ScbpSELq0F7DB4mJMqlm9EvfeB5dWt4iQLjNN4HEDKe24QA
lXBJlGk1dNpk4/F44uCMEWQ2pou07zQCgiZoirXHALJk62Q+MSgaMEDDOAGE1cju
BBSGBIqJwoN7pakmrRzgKwSp6LISPTPdVJocfbNLKaxZU7HzRrzMCbu6Aevv9V6h
4TUfGpOD0upbRLRi7FyuzXQMXY1kYeHgQ/5LBmB/jMFwcs821XR5ZznXzosMpS9N
eAGZCzGAj4z2TmHb3Id1IpZNdH4zBDkQRRiDjbbDlJMFNX36Sdx5choVQgQNoUpj
XU7n7YXnWYj+TDT0HI4WuTy4cMaLoHmQLkxwSu/OqmeaRDEqhLkpF3xb3GeHl0CV
sZfZa47+H/1bRhXh3RiRbs1pguFJ2qmgekrKAADmgENCFe3dNfZ010ivCQHPnpQF
1vlZO3Zi2u7+qmymukVPp7jPLJ7huApjWrVKlPNZVoMwKVLwbbU4q5Xqk2HpZyUp
BmnL+JIy9LWg9gsErDQSQqeWcjmi7If6TApVt21/XB7NlWi/eY1VLEOirbLRJ0J3
UWf/IOlJfCvvaxzfCPrluQODdvhxpgkGpErNev8KAt1/INuctePx08zvWZDyk8TU
44jDxpljF5au1HwROCj2WNQVPsQtYF3RcdrOtUGsGh5MrKt6eSj4miGo32AIunOA
rnd11kKc7XDcUbCqcxmfxImHsaunzRS/mUIUImfKToqlcXviv1Ea9yB+BTEl/v40
UHrbrxbsemC/vP/gu723qvd6CeLqJeBlke+KDl4QgnvmtHDacgGXC4wcbMFxxlXg
AvockDNNH4TiCMHmDz8cT5+A07wuKk9cCwKDKvdOzCJs/az4+o74ty32ZExUdnY+
sdrjcZ4NdadGVhAxkWunCCms0bjsCn1ImgbFxjv7wCeKRwYLmssAHzXtTltdkGoC
jkksId6xRC0s8+QeRd/Ndgqg+hASW4A7R2mKE0GaWTf0CgyREHVk93lbZq9bI85K
vl02CWKuOvM1IFdVmfr3FkaRVYliPBN2k3fWEHJBY/rnLv7vV9jI8loXnZGUHCuM
+MD0fEtY0kI+3NoJXtaV5+JUoTBq/afZV3YTeY4R2DZfKq6Ui3aQMSM6MS5owaAt
hTt+jH4BkT417wyPNa2+zjJQ6paHSaKz6cVr4Xv1oExo3BuTtUm530lX0PhE12yD
fCZLjcm6J3hs+qeefhMPz6AEK1froMf+SZwm6LVsG253a2Z2bzfIa1Mb55qH/+Ef
yxr0RFz5hr6HQkp3yiLUOTO/nC7ilLEfER4PbDG7GlY3n8VKMXL5ajbtpXPZwXmK
nw/R/sa5UiOhae9c8xYNJN9kuIJjyif+oNEwy97KBpSkZ/shcMiuNYZfhWKtgxA/
1kA7a4GdH0IfxU9BxP1EgQfqlAPGsdFq8vC+p58rPv18s+Tv4neTxoN0+tQtQ8N6
/jtsvUVJVe4lF2FFLc3RqOgv13SbDnLrbvhOr6FEZyJbYfb6qdfLVqZXFN7/W/Ih
PphNzPjkQ0rXIp+py5ppTZArHlwbnomcCsZfNH4Sb+nd5EMa35Ab87HZK//iskig
yXS3rA8S8P00TGjafBatxblkhKYZqNZjYssJWMepwAVbFRUji0uE7ITGD8zxpU9W
xLg3XtjmvXUJ87FlHvQgjqyi6ejN0nszBR7alTn9WpSdZKrPMmOCTWD4nPCATEkP
ZO+dfHC2k4ZamI8t+FpTRmI3QfzEalMulkL0IYuSaq/KTSSKiattq6UkJU6BRP1C
JZ+0RYXWhIdewyQ/08H3YU7DTPVoYrvjckzNqS5vA68vhK2VYO1WlINoeS7aHkdm
nRIlqTcAfW7q1hg8RJXfxXvzDXuRnIFjxMXpCYJrx1btlpsKmfuf6IRGbnn0Ze8u
FWFvEt2uSqu4bnNzxOiIAWYpR2aS1xnAE9gpgAKNdwx9csWeo0Lzqs6CpbIioc/W
ViN2OEa9PjpHRFLAH6RHFkr/qKjQ8SfTNH7KEbX1Ng3QgdVYAvchVr66N1Fczvaw
s5r0br0r2ezd81emHKDa8/nTLAxqHkLiDnwNWK4k2AaUTLXtgCHR8j+WNjZCfNWK
AXB/5mnoxC8O6TY/lwegWWaILQTe/XRb2nUOSbAEr8rphoRJV3vEnir4TZP0ma2F
xfpCNnyQ2gp3zsu6tgnYk7fZ1VCOVGpacKQS9GnfFeyYoToeqHMxafu7w7zLAYSU
69dl872uPYmAc6vPSQYXhtYzj4EsISNFX3ZSGMjPQr7aModvLoovllNytI2Qe9Ql
twEYkPoHjt+xkijsqmcCMjozk5lqeLXJ+zWGsvreck+YQ3YTGIhfOsvW6gRkjbca
gH/rd0xKqrqRkQdFgcfPzry/idiEb8f5mMe3TY7Qq/dZpHr7zq1m5sdHwfujf3/i
IXrGI3ecS6TztLaLzQVcphO92W7OdM0KRDOt/N0A7Fqc126J52pQChArtUm/NLdx
mXzH914z3ApQsja+0MO7m6uqGyRnHMacFDqA7JmQkBQB3BlfjY4Tkq/OnF649h5p
MzYq/RyI9TU8+T0tX0xTTVOkS/FWKPBYpdwzRzEuz+SVws1Jh+VsBOc8lizLHXMV
U13dfC5BfRhiWelNkAVkRH8RSOyBDYqdcT24OGIggeu4pVy1XMGcHACyDPcphnwv
H/UZZIe6XXYZzsPye2XG9ATBmjui5x9BJ9FVXACA2CXMRgTl7spzRhlkUQZtDJhB
jkgT+yR2pizQxYaRm8KjUx1r8gqP1FEjz99CIb6ll7m3ifyjpE632rELhVyZgoXG
LmEwV3bSX4YkNmkDzrvsPpwWAjP5x4hJtRPBb81Hi3mcwguu8kx3PpilopntpSLx
gFgTLF2CNapLA3KtMkhCUvoD4GAxhw338gUWLgsjcOjbyGdxp1Pv0WWGasvojKJH
Y+v0TI/+rWUbKQ+HjNNFXua1/Br5zg/n776OxsO4AGGVZJIbAwiwXV+Wq39DuTDG
Q9UapEBZuhvWIEhbyE8370e57PD3qzs2DAmi55p+VvEHB8KAbRYadWlWZM0hy91r
HKZGZ2BvUC01Uyw0VavS3VLbd1Qt3CUu7/gjHMYAGmt5m5LJeFqqmMv8pI7+BsuQ
mWJADElms7VfVEP/lb4Jpg4mu17Keh4tHuNZkqRQUrzwL9YwhAn5Hx9GI7vKMWL9
75zhAshR5RBI1zx3oQ2WrFRC2+r1RTUM8W3c7o8/p2E854w00Ko8FICM32UZZEQc
1tPxRvGKEslqHeHAt4YzJrUEwO0WxcjV0QJrzjQG7RK/1J2Cjj9/NCntWGbaZNiJ
UxBHV6/2kL2/y8qwITApV+as61N19QhSC7F1r74lq4HKkhxo9aylIEpZMqkwUdBa
ij8tzVEVAJEtKbRuX67RHs2YinIZGjR/q3Vjzz9gp+eXg8PL1LaWkSnfWWNpCMIv
9rjLmaK4xP8XBzGwxQ/L3fKeM558HNFkUH3Gcnxtr87YTWxBhXrsNTz9Wzemns5H
ny9ADBoe8dY+VOaCOClLQh7SMLLiKCGETFOF/5WpmbAiSRT2R3nhxBg58I27x1NW
zRaTbSf9km94PT9DWBXixuA6vRHMapwmPMRxQFPotrjBzuOHxU192mmuPma/G/Xg
RiwUdMA60lwssQRr639RtfiHvvE50x1UQRNRHBi/WBJ23boYCp3cocNCg1GGBSiG
sJVHL4ldptKEx4RE1+ePr+fSLKkqMSQVqwGi1dTxjdU3FUe17+QsNsM4LUWEATE2
a/sKVOVH1dEk9lELJsamHyEfyRO4QZRCdiBVuGNnKcwlgj3C86Q7kMaX37HvEE+r
bFi/7zTUT9CH/sqha2H6iUPaHmSZjGl03hKphu6smrdMmXHwXdosDQl3Q09wEhvs
kVGw0OuJsGDteTHzTt3fzf1vtLk5Yr8wNh0IW9X0MT3ij1vH4x/mCKciDoUIPSL3
66Ru2ljCTOL5HTTpei1vAGF1EZHyx4onwz7ea0GfOcdTkg5FaQuJYPhAL07/CZEW
3FG12vrSvI+xhXEgkF4RzK7clmqrTEG3zKkDsx0Gul3FrQaqrghorWxRM6ApsS+p
lavP0+3Dv3Ye11H7EXBDClJ82TuL642M9xcqk5HTmCu28scvZCQoqLKvFnwfIOKr
yAl+Ilms4JTLCBl9KsFHNNnEajKZjAUcuEAePOoDx4GILZkMN9XnlHsvOrX9ftuf
za+hfmfsh2YtMPv/4ewzJzmiMdiFk3yQWtJBRSMvi8c3O6fDZx/LhTB+FxoJ64UB
u2WbKmdzHJhFUooD5gvQtKyJpqSWr2gfKgPTN8qDQifzz4uNqCb7VZ0YiLPZAwR5
ys+5ADK3JEoj3Do6NRdmNsLOs+qekE5wrpIc/F/qp/IwuFUknSYyTX8iZLTNkuHo
OdqaCCfq2yqHg+UKKfflxgLHKD4KmsrbZAyBl6v721t0VE/V4uKzZetcjGrDJeKw
DtlWFdXr6m7vwJeq1bxtyamtNj159BwVEHwluBDnGZ27v3kEiwVaGRiqTKQ6asUK
D8cRjRwJXmL/cvShWvB/g5wWpKlk67jWmAJn0GoGSDoZkdENyGo2+O3L0i8iJevJ
BBnpT3JOmWZu43m6VGzjMpgmWJqeJJS/l8RH4n4HMLaxZ0rqZzeD1ZM53X9BRRrc
KZ+fhXVJJAaSdHcdk/MM1KbfgcXNckvG2AvqatJtXw95kB5MDrySexfb6h0tebST
I4hc/VyDwBYayAa9IjetYDfHTm1NieefnLuZkmwtcukBgqs90PkVYJUvrbCRM8DG
zIXJUQZzaxrEGDFYSrOOz9EDH6U2Kv4HsbQRsiQ3do8N3+u1j7c6mco/NUctv8DC
CUzFM3fwxk5FnH1S1BaxSWcwd23kYgMC62lHrxXy08PRhHplSBKHQHGEUYm8Jv0F
WboMbDsYdog/D3NVCrKVQt0hKcqHXEw5dIZ1ZseoOaYJGmpZrvHYuXyMFH1Lt2ce
CxG38s2ZzmLXtFZbm/+xCKqT2aDMcXW73dxSpoqUcI2+Q8gyamZWzxMRIZOUFZt5
V4qLUpqHk7bYaysHu61gZQI+BbxZyfXSUTpmoWhmAVFMG/eMs7/WX7swIygR8Pcv
TIbAf30EjeJNQ7itK5zUOsCfKC5By+tKTKznOyX4JMNuIVNO+2jj6TB7dPbr4D/o
Luk4/A0LGpr1tm4cjguHo7B7uceNbTHHNVIasCdawwU7tfjp8Y4MYUrWClB1T6DI
tQW9GQj1sTMc9K+L4mEyZAwqTxsQPrqTrV/IycbIexyOV1ernpW695UIPYe38lJc
w/V9ofJLsscD0reVlgq0GGPjsvktw1ghljDCU1cxPhwl0H1pNNi9pLbl4v2ocnMr
7hm3p2DA4azJABprqUi7pNjBZkfBX10luH8xz+W1BXWJNcUrW90BDKCtYk51xAft
YocfYX38uA1ME6tLd9pcT1lRnyGjR6y1ohHuJ2s8aGJv2MM4mUPLWRhPUN436dhA
pOC2E8dVJ85MgENcKTm+WUWPjShgOpA4nkXpaQU9PamivhORUvZhKKC0jVjVLPja
2YbuLHvSgZhFNCgfBih7zrf/VHNF9CWCFDREm5qUow/70ttqHjaYMlw8iUnK2Us5
9dPDDzeafC69vssipx+3XMr3zIZfTqgZHyWTylyZnGbfhZWXbak6SZdyxxBK9WhK
eU/wiDB8ye7nPRtkZSNQkOHbnFxfh0UHQSesechsp0QFkZEXSSb5T03fW2O3CpYW
jVq1Ja5LiZUUox3gH78jbMs3PxKOdL6svhxK6e+JlegEClHQuriBwhCp3imvKw6z
+rnHjTuKvNydkx5pcZCLmmmMvqlVQKaD/pC5XC7Co3HjoqtKH+XqnnKnvf0QeRRe
vq580Xms8V/mNkDOMvLzRFxbq/Wk0UgvA3Eqk2vG9+ZQT/2aLvHpoN5LiTCLRxd2
jaTMc7gxsBib0YHTjdSSrVGbsSrNE4ztn3UEJKz8kUchhPL2NARok3bxNb1leC2X
xiT3pCvTptyKP+p8LWznn//HBgPelNPOvrY7VTgAx14K2RbFX/H0A08MDoSarneZ
+mM2lqzyiPClrsgVAql9d1RnlibVBdJDipz6+R1vR0bpP8M5xB7eGFGg0WrQvJEY
qGlyUV+Kt/IrhyW4HJfZol9qMVtVK6jXuEXs/7lO+btgkMKYDNFcYvhfVgbSMm8v
JnkoNchGo4j0cFfPnU8ZFbHcqv+kilDh6V+6yJpWCnoe3+LYeRWiRXPpQ840flKs
tXSzJYGX9DabL7JbvVHc+xGxRypY4Umo7TRIYQI9Fp03baFQMwLa1of1SGYF9gLb
wy9BPjmrDotyeP4P2eNB41jrTrk3WZIag+1mX8FUJk0TV7QOFJ7bU3V2VIVsyAFM
7yUtwVl+um7cuXXFU9VNK7+gQUvbKifiy2Kq8Rp7Mx66en2rn5xFyyu2bgJpkj6G
j3tpZaTZSsI9RQYbAkcYGHysBUZz/G/yJROcqWl19sxkm848iBLXq4bGa4t2PChk
it04u4syjrc6wQxfQCbUJ9znpxXjW4TN0s2aoPOEtcQGVvb1Zd4oojN3VgWFvTKC
RyNlsd33vlARHHg18fQSzlsjwrgZGi3yoBWq34aQcis/WYJ4wbgujY8z9jmr0Gyn
qqqsjKjDso27H6HDz3ZexDSSIdyCkzD/iTNNXPo3l4ehgpwfPYbpfAB0lRux3H6w
IkvPhpuuPDM0UQ2yNGH0mB4AUuLHIch0z8wP+GzeW8cVDE4yjxTsG7x+sWZlcJoC
esfrOvjjrcAWVdjOMq6/WBngrb+TcPqZq4CdH0bMI0W3kxdORALKQKN5S1vlRTrY
xc7ol2u+9ERQMxoK5R0wW4KexiNSYLBCoGTiBcSsuG0M24aiBDHCDfCVQWr4Itu+
PzFPyGWUudC4oP8DXhZYBJsfhIGpQIpeAPAwL4ewM1kVHY6yX8KSHFEDydUa8ZHy
Us53E6Rk2usW2Cegk/VzP2zhTedt+efNlaLBMdOFKaybFjE82IWYXzB+AOF/Fsb7
z6wTFYtiwepbGWKVw+qSzvT2u3a9kmLiaLdaBFyGCP7Qc7dtuALPLi4V2fePyvAN
qPJLp7kf09NcaHTncjFEC68Hh1Xc8aJ7JyEXMMdMHc3aKWPDNakD3zlYx9lRRH2t
13u2zBXPGJlmxJjCdLjD2gCsxtUWSk1mIzgGFMtAfIr/dUOjD7X65gkZGgZ4NVX0
R18sYJpMddCXLHAoTLOZixmnTw+fd+X1x+zvxTOXZGxTP3C6/+2MqUsI5dU2KIKW
HFhDzwfkz9PVs9cAAVbtrXP8v56XfA21VHVC5tfUYSy5GA8qMUO6fn0UG5TH5PNv
52TIuoLbqQ0/sTAGNwgTUOSguUKSMGKlr1Su8bMGTC/rJACQ32KAOx+oRmY32Lh+
sZysUlkbP7bzWdcu5uMQXQEiblX7+RX0pvVAYEaivFbDoPLzgyyFDFZVpsEm6UUT
HawluBMNOjyDwGqd6DdceBvSqH5rHn1PbfDtdj6SNzgZ/BL4GSF+s/XOB7den6dQ
zFO8lsgoJ5rrpolzfiSIC0Ca/EyqEnrG7cgZl4A0xtimnGldH4EPGImkpijOBvWD
fxcPTlDcCMJrV167IvsfR9NikUjvUcWnUGVW1MBX1tyULz8LJKNvkb7FbzK3zX18
83iFZQaFhKO5DrypMbPMDxPTR4mYdbbxwmWZH6mk1+qLtT7PABtYjsRYPOBmPCRx
L5bP0A1ubJRXfLZ/T6eHVfRna/BZOpC7pxdqdehBB0wffTjozuj1YXEopYSPa9ey
g5+6mgHbNQw2zt8hO30QbEpIZxmW+db2t2QuXebQPhu4Zvc5PVAjkYXKRw8Kf8zZ
6dOpoWuBkF046vikIseqSbG9vpK18Ux1Tw05il5moowIehSztimT589yRU654YiH
qzP104qvg+DRNAZdS7pyW/YMUmUrkPSgooRKy7ep5WpCF0ryXDA3IIRkNLc3eMRQ
r2+d64/YzhZD7dG1bpg6GM2BIZCtOf82fgrHoO/Rb6/QnUgJ13c0Bz3hxpPOc0Yd
Hke3ikIp9bGJUlxqkG5XPm1F/yDpACELtm02HBtc4UpN2ELDW4rfNzQ/Qj+5VrgA
4myaE4Mx3WEK3Ano+Tt8WqFaouf2FYMXaE1XI4LyJG0z3nhrhTFhHUJ0NzCRvd6J
KZ+gk9XdqLVgkqG93d6KZOhp4YV7iaKsgvhC5QjVS4dr4RK0cW2cHRgLgy8ig1Ft
eIeKrjjJO5LOWW4jdfXB1OeYRAJk+io/X9XMJ35qYLZE/O9C61TWM5uUE5xZgp96
+Yj0MNezBA5MbMOC6OXgbwNuRSYMhOeYpQejfuUDL1p9ttSX4hpc6neKN57llxaI
EHTxZgU7CcZYXdESdg+ZnP8UrGeBpKD42SgzYjgXlQHw3z34deKvQ+pVHCbS0I7j
j/P4c3khp9PPqkw/tsdTbElRORYpIr/AWD7vrNsows1UZiSv7tqZSZQa2nyQ296j
PeEq5YvLQuo7c87RwaU95CFIMh/RJlbLcrwxjNiLX92ZQrw0i6/Uv4CR87mH8wYT
H4z5E5xjqHCLa0R8s7X0Ax/rNCwOb/FrAbmAcLTzK2ztlhzcfvfXcCIos7EOYV9S
ddHa/2oSJwYFOfDOKit3BH22XeQ8UAqc2ZaWE8gG0kH+UgYaQi5xCvczqEvfH8hv
aU++U7ZB+ovTiPVcA1whTtyhKPZt/2CYuLbc744hSUUMH9PENZvdkGw5+1CkQ53q
u8DSGSXRQDnAHCfZQBjWHJDRZ6xhuow6RHknL3UDptDrfNtZGZqEc7GtDag/vdmK
5cM9i6f5uoqAyf5JGaJwzcxP9RYe4OkxKpbG0i64rfA9vP88c9Vxet9DQ7WhNw9S
wtKanJqScYdiRdrBrDiL5qpUEMVR7pXTPzwHP8dUnjPrPW0OSiigjmvjTudFTLqE
6RQhLkpLyE5BFv3nQb18+8TIuVcSg+FKxufuGUokqXiEYz8HomoSClkHt+HbYI4r
2/pnvZC6Jk50RBdAHctaCvWLl1N6KygnpvLmAhlTtG6zHs+T00ayz8LBKG0Fg4Hu
2fgEJ8caRO1sbO+JC9bPqwqn+02WElSp4Ekolnzp2ELJEf7l5fcp4Kes6nDpdGxg
JsJol/z7MIqDrDss3hUzRskYcceiXhPd7d3GR5hEJxpHg3YYMWEYo2ZWwn3G2MS6
60/Xm/KTb6CFQihk+HrTiHRuguMPANQCeSSKFW+7rjEy5ASIdKUXMV5wsaA+oJ5S
cvvKw4n2bmYU8psbXy1hBtlja6MkOBCLF09Ug+MtTvkFc3AZ+gM5MYgpA6PC4bTt
k+VPyQrRH0koUtF2O2Wk2DMJ0Y+n+aVJ0aTTbq0j2ekQ5lSAgNR+Sj67FrBb9sSa
Fvx5AooIqGo+tv8DCzh7gbb9bMKCTrvPDwigXRgNHnrOtZiNJ7Qyi/j0xUmed37g
W/ZUqfe+/c+fsc0ATxU35+OffACD6Qc1CNJcQUtupSAqZa9jANvbvcM9BS8YxKym
9CfPXgomNtaVnHSyb7cuCPQisoTThmZ4zurR8jRQFdFQVm1To8RoFHB99ce2c1UQ
u4vlQz8LnnGisnGtXLPnaqWyqjf6CSbEZBc9K2jqP3T8RtQ0CdnKrL89WoJd0JFL
uomzlCPs/UzuZndUvpzQlEFURyZr7zZowMcZ0J6KNfAi6Updl+wYve1Cn4y+nHJf
UPv4JwkTN3dGVPFCrEVaTsBSSBpxGSmc2UhAbET4mw78kpNHB5skx6sA5Qrqq2ty
mS7NsK2H8+SaSi1ILvyjkXB4vC4eWH+Kwwm9QHb3rf/un8snqSSX174huI2KfNkk
qGebWl2acPSqlfmQSZ3ty1s+owI8YwXy1YcDG9WifpG/w//UAXXLgBSuVJ/Y2yo+
b1CxgRwnWx0/Ux6+GETlVGXdqFfpvGQb0zugTFMPMPS6n5n3t1E1aB24dv5W8Nv5
z6GK0Nh3W3pG36ApMhbh0tUPv5ALfC/grsw9n9ii48LNbGhC6cGDQmUaN09s/36D
LcQeIf6OxRnWPG+quNDVX5wd5Et5G6Z2iGqP5sSUPXaQhXvIeIW8dlAmaaeS7msF
0Kd1tec+f/XeLdu9CHv999K/44JFnkHPCA7c79T0yW5x0M0XNXf+HKX/Gj2QCKB7
OuarLDsnC3hY7kECd5023txtymcyZN7P+QTnKQfL0dh6V13fJvGm7aWA2aLKP11U
wsTN9lerUPe/H1CA2TXu940rXoy6AtXtbzJyJfFSGvDWOsv/LoNtlY+ZcBeSpnjQ
U+m2f/5qwVaxdGdX81uoByujvj1+JrYMbjVwQEG18h2wiBppr6s/jmIn8VHXBcEs
626h4P2Vw0+M67OimO6xXSYz7YBFwJK6fKZFujtmUPtsunsmAYujwXzH5gXX8enE
mArf+o+nWPFiz96Tq+UQcyT85+1a8CgbZTUCK9Fg/VzOhzp/ZZnGJcDtuXfxAdXg
pISrqssBx/EAyRgJoBJ5Dv1Igu82yBGOFLfMeVKhRWxopg53Z40xXy2ngPVqzXAg
6qan2HZWrmziLdlSkoPMiv3Kl4p+k2TQgIYKwo5KoAI1sbRlgcJKyg3eZ/MUDOFZ
RBY8fgIVbnnChjyUBGkn617AeDIT0DpUNa2+ZH+jQlEafh5pw6xkQqCn522nHOio
fF3YwN9qVcTYp78byRv5h7GAYDdgDKYeY/eYRPcWMZiFO3Lam+jb/fXxZ5q2lrgS
RV4KY4LQc/QkfXxrcEqbghG+bQ6ChdWWrEhiLuRHvHZNt5YJpumR9n7vPsOAydve
RmSkvGpVg27Uqkca0rpyFJydHFkm7D6kGRzi5U1C5sb8lOcnmAfTYqy+1fMNRkX3
dDi2nebbTyapES79fjCfiyPqJ/9w92Px0Fv+MAs9cFfkfmSysMQswkOEL4TLOy2Q
5IJU7ja66u4SvMh1j42TuuMguyyFZwtt2+OeO+kGD5Erg3FKwv1oUF6LdZL8PvoR
EWyhyorU7e5XCyQr5pLLe1h/HicW7Jg/pZg2Z/MNn2g0j+JKiCHRCIFwU0YELL4D
SHl9D+vHvv2Dbvu1GjGTmsaurDPZK4Xiv02ySX2G37yyu1hjyaPBcRPkUkNfyv+8
Hz8uChTWbomYfii9BEKVYByZkZjyp8VfbS3+kw19tSmuxlHtAkUYuM3+x6872czo
X4s18CVyerOHxIcgmn57ALYDVRySVlvOFzh8M7Px7M3FVnc7ONukkEuTvnpUkbgI
IIQeYfw3I71+3Q6vFBs9cKXNtG9woq3H5uOXXvfFkcFVC0xJhWbhon3NACk+MoSb
ze0aiJiT7jTc/v+EDyonj5X4jwYZJVFie6ZVaXK+8A220XNcA2PBCXcrJ3qcmgx4
/OiiFb3rYvP6tgP3M7DBiUxHUcXQgM9ijkE5QPESMvSmuh72kgDFAxQltrLbmwPV
8cf8jXbviuugWJKg9nYEU1CqMxp76JJuWDbJsGId6/w50imf8XySZDrQvN846tjS
fyRvabppsLa1/uptNemIQ81jGm6UrSlwTWYGkZDWBiY3Z4F5gOUOXl8k+dQtcW9p
qxQHhcXDtu4/LZnz2L9NhrsL5W4kYhW0X+fDI4XkSe3Cxcn3d8BNiHA7jvR+Wkks
yMAcjhkUPkqE1kmCQEYIR38KK629gqhvr6PBMOAziiemTy51KmD6tKmRwhn4GuxC
afbhXgM0GNJZNMEb5NTNKtDnaaUwJpw+lVBhVcX3Qj8Rkvtq5n51paalNuzfR0bk
7WNMiBnSReZRklBKvWSQylAwtgNcWwKBvWhCaeW6Yp0Nl6OoAvRdICepQBGzhGVV
TWT7SqNA5huCosb8WNTcwoTL2hcerQMKD5JZ1brO1rz73wUCr2PnPZJQzdny06hv
2SF1Vief1LoyqK2Afsdpn3bvC4OBu8guGFC1G/m1HjC+HjKYXy7HxDZ0sMjQaO7h
bYygYydBu9YkB7FzFVuoiik4H6hSqFle2aPQJM7wUi0hh6d8l8mlxXaREz4Kg3S5
OWVlT8etbpp22q+P8LfShG56+M6AuYwq8ajH4xnpSq5f0yjYu92Iq5v50hRanm9W
DCdSRVnH4D4624HyW69nqr7Q9THiJsGeKSg8meZBI3GjriyfG36ZRPZZv1PjOKo1
hoWmZX6kpNGZhXdFvH5U8FZnsf9Nm8j6ucmm530pwMLzKEcTYKbWtoUicsEGJ6H0
9Qz+bnDqJX8ZTqe/pBXbs0gCY9bJieEfKFuWUcOrV8vzFFCGQAroFII7TfZcAOJY
c6C8OjMweh4O6w7hlE8ruIWK45ezNgex+vAtCDPtE1oM17/8P9vu6svpzLAWKCn1
H+rrSlj3ZPJYHiseu/8xfNbzkz8XDVSVpilAE0ZN+kbFbAoe/pv4UaQ+4v+k16nN
i7gvNTd87xjrA4ICQ+ZV0l+ujE8EHMhQfsSC8Ho7qb8MQMAAwVho+0BehRUGWAxf
0v0+4xEC5ySjwjsiLt/fNN/sPKAlMLXvD96cuH+kZCQKNLhYiyYt6nWZS4zKNg8D
A58DBqoGByW5aZ1LNwqq83Si1j/bEzIMjM3OQYf9zqZd1MH6J9zOQPKFZIF/vQEx
lBD4fpF8Qyi+p2bwPwQa3jVCSHxceXpHIOwNXk9/1kf5xiAu9rYz09lh3VMIbmjg
Hzetz3cpi6bJOeKUi3ytPYs/R9oA0rMC3w5MZckR8VRb92vrBu6WPaedyoLdnkcn
XkB7+g/fOrIH9eK67d9wtMXeJ8zhRr37FkjbuJcSSu03h9FqbQCNox30qJQwwd5V
UMj4Khwc0Vki8MMK+qcNnXggKTpmWyVSHNWzCr6Xjs/YV8OLjOjW4VupJgYpP87L
vlhWac/b1tWsaDbFcaLVAAD9eFCnH/3nF+4X0dm/oBOAaEzCs3ubDLPS/+71s3Rc
I95xVS3U941ZDUb0fzNkyzYchD0NP18LepuYOwo9/xmAhQoimrLCoCO8PnE5LRN5
l72onTdjbE5QD4Ui4O88Y9Xlelvy2wMHSd/q6E1g04Zn2I6d/wTI+8PXNU5BVS9X
kgbwtR24+uBG4AbL21ADtN69cZTICmw6IvOKjmQexEGNg+HiQX6S4wFbjMC7m9LV
2SxqMNEYJYvhk3GsJOYGgGprqNMh9lgCgvZiu5mBLNl6mHK5ZkvJiZmFrlFcI4SE
gL8FbNuPoxqjYkmXULG90lHldXgUAX0bmN+sPrzAKSn9AemTozn2jwvsrHNgVtXa
Le1PvVJcjQ7Tt8CrC3nqFbXCyMviUy2++DVr7lTtrXvLYV2XwjYEdyo5UpaBqOnu
k0lkgL7AbXCg4v9nWYSu+57KtQfnn9QPjEdqKckpxHic3+5eD//mBpFRzz7SpO6l
lhwcHbK8tclBc6ZSEjj1BLQ7O22qVIr/4Zr1rc40L3RJgeDMxwh0Vxhbk7iuHXth
OzBxvFEuvtwGWcs27qQCrZMbrrwGWGE8IQgmVIb2NJwjRKLOwzkHjZCN4pI1r2WV
MWAY4ntgggpHitOd2Cv7CDG5d2VEO/DWjLKusjuwdJ7pJ1oQYyMUDirqJW4ZIxFC
qS875lmM4tSwKAOBKHOX2ojg8oZrKpQOxPBEGDRZ20GognSHAyjvxGE7uRfhkC7j
ghMSe+HUN3P2SI2St5Lm+yyRiFLqnKNzDeFynJvliV4BR/faWYu1wLqTtkJ+Mg+1
Wc4xzWIciatfBoQCSs9f8WTWVBiJjelFR3WsyaiiVtweraLC4vnozJ9Ckcothnrf
mwPlmc7vP8ZSAgbgnohums4N3gpgY3kKwk1ilVmdwgAmzEHScuAF/8yWKc91J3hw
yqD3xoeNTypnuTGuk589KpPqZxzWNb4zNiovnc6idzC4kQfdj0eMZMNOjwsHojfM
MQKUr0X1M3p0oJIvlw0Zl9ANBqWDO5vdEy34O6zCsuGCfBWGUNgqxhiHz+GrMHbR
0NzpMIIy2GbTb+TK/Af76Kz8pcD6ovA/VEX4Lp0W4vkx0ShsI3IxJJnBWlYZxS+8
gSl091E8eYCWcNkMcRHA8h7ReBX3ZMS4xsdUq8kkGE++bLzN18E1Y3rV1b+U7nql
qJrZbHc/ydgKq0GJRV+RjoeNfr5KC0c2xbyIoewtRHT9dvjBntNSNjKjW1wgeozC
Xa1iOplBXqlg+W5YiKlpzoUrE3gGwtk2dHpVy3PsFjkLvkkHRNQjzmC0+nInfBdp
cR+F8YlsFxPpYUg9ufnSj8PSaT8J3q7qsR+mDMAVHVjGCjj+os5DKnHOAY9wLY2y
yv+JsCkUodgtiEft8YGo/F52FTetUw2HcNKWjrg0nnuxmqR/m0vEz8iOy8yNkmkA
hy0tHd5uddMkbujrr1BYZ5SLA3MtHFqBR/gtZEcDPf5XGHxdcf9lUubVYbI7mcmx
AmiGVJjVDLfaHMbMsYZ5p1HmO/d8E6j8ZkEmOTdH1WYXTLMx9eyxq4fadfnmP5k7
4PlK0XAYFPHhE03HDh6nrxCeJHp4V4zBY1fkhP1WU1c5D61UFHcwAAJn3P222eNW
GzqappjbKCoiBuHbNzZnSFbZBy1xyC2B2UubWoLXhfMOpokMf0DT1oS7P+P79Txs
0KAda2XJisZA7FnNLO2hYdRJNkNrzQUuxjh4n8dYvqSU5RUEl2/L361h9MdnjhNU
hQ/jdIDltCbaS89wCDBGvp94AP9fQgbtDi0sF++Y5L2dWp+oqW9UUpqTIXcrvpCB
7YAx5uhm6trQf7g36mNGLG6k5QYt5Lsz1GaElxVvaBsGhFcVFJa54gjhhz2sPTiE
827N846llFFvcODljU+XC54frKXy0H1CP7epOQkCckWnAmmnYmS38/KNG1A4ADHr
uw3iit05oDxOwBlpuR/ub72rZZ/A/JtTCp5oySWE7A4gvPms/QacifMF8WC8+BGY
qYWI4VtXHgsujQPH8nEX8ha3kx/QV6Xb9PHTN//cgstg2wKhR9hP6akI0NrsGNan
9EFvVG6KzmCoVkO8T7gSbqYHxSw0nQLkLPeinNz45gkkib1dX8QDXAIsoBJoPs2g
WSn59uUz23qPwpRyK6RMuqZx7b5gC7afXFTpfXUbTrtxXhRNoJo2lqbbLyfENUXl
slJj8ubMoeJhK1H5Yx8bTd/XlbEyiblTrH3eA37Z2hmpWtxC+Hw7Fr39fXM6hdA+
gkvjR7COvKu81KkZy05a1nRkdb3vK5hy45xp9KXwFyDONemmDe1fge0twJW+dHpL
UyRfqRPUraO0cWHHYZKW1nHRD/lLmRQe6LnwllHX9qz2Z7rASmW88lYft5HsF01y
IfLOTgFoRUNPNisFaZrUGLLvyPRqC2T7Rm7OcKHtq8oJH+Vjl5gsLF/l7Iv+4Sv3
OHgxj+STT+eG+gSCa8bZ/rCV+3sa1UPdJAOmkFLu5TI6N5+vdCaABrArUcO2bHVO
Wy9fHpwk7pmmEsSB2tg9dwo7Sw7xQl6RR2J76LUy26DhRvhrtQgwoRTjRM1Bys63
BSo0gI3wpTaaWoceogEzWI8BOdNV7FMvXlTeBWGhvluA1Wbr/wiWUQRdhQjumgk8
95GPDpnsTu8JlxJRV4053CAQeRjXWvplhULwzQadZTHdOFuQUsaCrMYw2MZ4WW7W
shvnKe5J4j/aqWuEA+YyQ7sbRjQdQaJKAcT1hHcMRThla4Qm8utAXX27FvZT18sx
hdTlD221mH6J9FFGLdbCK7v+ePIuUhUMKZ9E7s3kv1FQhISPuC3JB2l0csvRYse9
FBwI/Hgb2wBlClI8NbCtS7e3o7xlh+XCqVbKDhQ4Dg+74A/346B+QBS0m7utJXdp
TKRpzxz+CiL+IkhipCbbcb3Tv2trSauP21wLBs8nKBMZvurSllWR8o/haBZ89Ss5
zaBNV01K2VUSuzmk1yuD4vXp66ew8qTW2q2BLe9bGPLFPIgQuvVjIekC4GzuiRoH
8+GkYO75/kRVbJbDf8YaSgWoncOtOLo4BfEE6y/r/wcdr5YonAiv0VA+nhh025Sk
/S6xxydrbqJ9cuO9OgyPX84t+MpUkS1geQVuC6biK9O4Sl9wMbquyn/NlEOkPlor
sTYiUeY5KmGyz8/5YaHPardLI/Lz8yKpOivOzz8iEZqDZVOqdeb4KLHd112mYHE8
6IvIh1+Vv38QCiDOSmcSWFEJodfQe5UYoX1srOo3L/dgfrGOhy1egKZeoHLFqg+s
F6qEL/8QstUVykPDnPf1bhaRZT0yvdJh20QrK5s8ViARdFvD/DCy4iaD20iDveNP
85zjAI7EzCTDe4DFPBUEPfjU5ZP/Wa1yjLBRg0ig9V9z7+p/l8ecicGtTVOk9R7Q
uMo5y30uP1rFWU+6qk1T0BHXoOFYTDXVqk9rfMWTurSy0CnQxaPsaThBhdQLp1NM
iNgEa9RY0HFOu3sNngIhZYoJIN8t325COD23A8sx3JCLBawLLBouHUcfEDHkdbft
6CQL9rVkOVO9rHv2QacEiPBCHjMv/RU5p7heWjMutSRbYVyBRIJXuhdcAFsX+8iK
B+jVOjh+ultSzpDvpp4sisxWvPfeed+swBPOp5XuRTIsNlr36Yn4ia+sp/0qMWtr
Olvey4C5BgW8YMO0UjZrdpCOnDepGrfcl9KKKW2lK3CI9olC0GO3S7Ch8rJ27D/W
g+sNZ8OGvlvUDLAaRUEsxPAh/A66B0awc2MeGnm3fM0ObCzAbl6qF/GNu3yiBpiJ
9niPFNXA60l8SJUlP4St1WK+yX3lvgNTklO7GC8zvwL1mEnNrb+YdRGhUtucocKt
GLZbNSzSNJE75wcGUCGduGgYNOmUqgiJEAOk60dq9nFv+PNTpKQ6dm3xShwIICAw
InAO6yCRJJoU+lFcwF+V1PPEtAayUtqsKZPdNvqHA3uFVrDCl7Ld0RrrzcssOaEo
VR9QyzE8beiTFzdnX6uhDx47cAzsbT8japr+R9qEQbF5FsdRWBpl57zeVJHapJ9n
LVhQ7lV6eMqbwEIa2RFmZjb9Xxnfqoi0y4EaAE1jyOgwe/17HO2sDQRlo4FlWc/w
TLfZkB85/t/qL3SKcVuNmRPgNfmP5WD3YuZvjElZf1mnbVlpowQ2OhAbVKamQW9w
CuboxlqtFutN+GgdUOCtFBVRNAzReMElLPnc2ETQE6lCsFyO7NOZX0eepZzXL322
DwSNlhovRG7pZQ4WDsazJPUd7NSeEHzBCKdpqE7LbycG9TT2fpS5PIKPDckCtO4S
DT5u/Fjmf8UDs43QjxpoNuy+syi8GZxmEEhKy0FDPakd2VCYLgdVkBe3/TiEovVq
HGMr7zDMvYHCVwBzwWFPhAmETpw663JXJparvRUw0YcBQ3OJZmi/RMo5J2iGpULq
xu0YIeILGRtCdLGM1EEiHNjQaFwkh8Vpt90mjDtjmIPTNrSJRUfH7w41zu9yy0W4
izFXyHdFDxcq1941PZxqtKQZZ/m6o+jMRc5t7pw0JKKJC/KVgWhgt26GQgHlCvu4
BbmkxpuOO8+qSv+UbNQk7GnbRLhLmtTGybN/owxCTljSN5pWBXrJ76QUMNaB7l/C
JRXREnXs7HrXTq6R5pEnXV62Bpg4GD+wJzFCqU5cj0hF26WMxlD3ivVXa7eBDb74
5S0vF6w8ql4GVav19LbfM1OCSFUu3lpUlLahMLIofC6V7wEpEhinltqotoP8h5sA
c+zxJCWg5XSeDdBT+9X8WmH8/wnLsd2Aloc/OicUlA6HLUMXAXZmIx/chz7kdGo+
RVruA516wc49XRv+laSROILGYK56LBOtswNCLYoFd87bA7JlWK2ALfQZDXz/XHfB
OXc4aL2/yVIUG2IaoWcsjFmWlJFBXly4UEnzULmwOBIQS5bRdALeM7CcXgKd3TMe
5TiBBbbMPV9wf3JG+82jWB9/A5Vx0wWSXpkEHi4uq+/BNGD584xauQrl4rjyvRU8
rKgWT1rwn5AQaZba3iH9dWAgIYd4f6nI8HEcVfvER5vG9CDpxTENNDdAo8bQckrD
Y3NhKW0KsNYWH1dbUAjbclYDtNDfyhysDUPf9toGmcI74aYcoX+CAhPo3wDlr/au
V8bPixLp7g3kELGfFoWTUPWKBe9aFdh5yilRM/a0j7lqN1wLJYiInPCnBY+JAmkG
koV/GLQ6i3CwlSA3EdBbM0/1NaL0sCyofTCtunHQwbSJWmC7GcX4nnErboYPcaLB
9JhBYFcAqHACngRwI2cmdYGf8kxUj4ubIjTuSFbBydS8F5wAG87HE3DU6YmBdlFl
HguMfYb+zVpN/rkvDSOv7QlpE/zzskGKxzQMVf+w56JmPwOu766aOsMwdBwhjUeZ
Zp2F9hd1rN9FN+prxBwLawCh2NLAZ/aKSvbLt0A0y8FIHWU2nIUF5neIinmFo3nr
tMDSnGblEFwQhmPgWGvaizLp4owSxbha4TNzGksxhMO9XttYDCiu3wjlvJeXTEIB
uDBu+7wi8Oc3j9dzesVW+i/tLwo2gAWaP9BHBTmgYqvfU0JOpShN0lTRJ8T7vwMD
o7t9uGdZKSsWNIrMNmzU09dm+Z9Y+wYcAT2LvIMhwImyMsVfUIoi3v8t9E3UjggM
4ngTVVn7gAeC1I7cE6K8gBlaJkGegcv4B7Zp7DtcjkNLvDUFzCqqSbTRKnB6q/7N
GP1iQNlWpUhPdhNvqmfm529p8MbgthjG18QG2yu7enWQSbt8s0akpcoJeZyH1EYa
gJrdO9hU55UQEG5fk8snxbs/xwX3nVJD/DCDoaenyg1wraw3pQpDxcQeYHdgqtH5
Sc7r9Ll0sBhh9fpoa+F2iO6MF4Ue+DdMM5piz28X1FfQnfoE6f7dM07ReOihOSIY
I/vbbeD5xZP+wgF+W0FNO9SExsDlt+Wryvx+6IhMtGm7uIAvWVH2TZcGQXdcgtj/
9u8PZBrNx+97FDilLo3lGvZKF3HNag9riP4LZgszmx7IlUziCOR37bAlMt95/wR1
s4d6OqK/6+V20icB7alMCaFRyU0d9qMSHrAO9lMLnl6Ixlz0KcCBXiw9snBOnuVn
7ryod/2RmyUFBB6LgJ4HeXdEiHmIT75KGZcbdlnz4JpGewF+EsIehORJVyemdrbA
CAKts/lZ/y+KGmt4VVLK9D46yd2kq0uDgDlyNewka+ty/2MzYBb8A/aafO+A1VxW
TPB59tsogY6iqm0D/u53JB2Bv0TTrUQzPvYDWH1uG4VyMmZmqXSrxqgM6wLtt/Na
c/kjOjBuIJVMFk0M1oZtQXGNc0hkDipPo+i7C7piWmaBqciSvo8FZJEc89GJT3pn
zY93RXfNIWQZB47xrrAImQ0kawyWwQkYQ0BWHzwvyjR6dYwgMGq/PeXFfibM/p/4
MF0i/laeqcaXWsF9n67vyiMXO2RN8FJ+F0BgdEhTHm/Xfo3t6f09Rt/42PnvQ+YC
N7oE68tFoAP94ThCJTnRApcfis5nxKVgwsv8sj7eZ7k8z6eVMN5AZWdqxvi6Plsz
CpTyihQSwiJUlD69Ic4rx6onQm4BHJoqKAE43qOJVeEyCy/FdIX8Z1OXkZPfDYbI
TodPKuNL5fsgU0ZiYPNatwXQTfGp9cRfjTD41Qp3TY4thbSHPNcG9M7J+/hlwb8N
qjUaj08XRec8yMJx2pUin/PhzDmZOr5/8FTYtMXiYnm8IrFK9c3f+XgObx8HfRBp
uxy+2eikM3bVTISFn0PJ+rw4AgH16boO2zOFCV+GfC76lIjdq/D3bgAR/GA7qoMz
E2cimbaHR5XEBKFCMlKlrw/BNIShroq5P4ADg4CHV2n6P20TRCTwsxk7RMQ634Ud
3V9xXoP9fzbsnlYQ90QnRiDQRtctGvTng6ECG+08xpcMQw9lYssvIujLyudOcjOt
0A4+5xbw5vON3fFqnMox3ddXDqkCTwX0g5cHN9m3eszN3g400/4RuUI/QtNle2Uq
lNGelgqAxrbWKnOu9kyVWd9ZWua8KZLlz1qwkBA0mHmFU73ayl6dV22DttJ3ZyoL
3vkbp+Itonyu4pWWjkg0CsQXi4e//NnVjirXIbqOahBL6lRUlDDO9H6uPVNfISRL
eu9/ZTGuhI+NJKmqXS5AfHkr18Vm+qGnWvU76L/17u/9tOVbOY1Lo6T8MSfi1jWm
gzOdx1dJP6eN8RrQpTgDQZZX08XYZkwS/90/vutx9n1dcJa3lWLkrhsPZU07IH97
zyok2Jdvoh0v6T6C+qXM0tcicelMgCUhLMQ5M89hnNlcEu6O16JEv+NIG0MuVjM4
ij87dfJ0BD7y7WX57tNoewaUmo60+wqmaQBloBHO8hdrGHiafLKvNv0B4P9bbYty
lLHYnk0bDMudyikgPqUyF+PXHJGWui+juVVJ71DtHgtvofpH0jn8IlcssKYqrUsP
v1Y6DGEBY4G6nlGvenZXU7KQhO/yJrPdldzedsiFf6mFVkBQcZHAqpg+NUcp0PYH
e7MrSOZKvbrkVO/3/lisC8s/1hKkoTlovgniKNMK4W/WyfPeviYexdAZCrZK76qX
iXiyeiBN986I60/Ko6QNXA6RencMt/sRKd32DWBYvQ2dFLJWyTFfri4gR9xL/qSO
Ity96PF9mxGR/HaHLtegIa3bhn0Jen2MUdn1ww2enc639V9Grm1dlHoyV/cCqOaW
2wHD9vtInPuPHm9sDSijxnEYWhYlqZmZXeBJqr1TSK+mVGk6HpTRCY6GojHyXPn0
OUEM6hxk3AvgMH/xNIQSb7qolh97O1lEOXJLkqi/baVxzjLfhgxkg1xf+ZRw1iXl
cM5Tv5KslApcXp8C1b0J3I0RdWoPegO33qb8O5e8wdFG04PH9hJlPQ4NsgI9HzJk
75hbWhkuGKLExDRwhNd4MVyRlNMdFlVHezB7uRTtHbrV44N78nFJTeqVEbMl0B47
Xd8y3Nszv+guNIXJosmNAxIGh6nbroTUo8ciXXljrMRRbsWQ6lreLPxY3e/sCDga
2JPSAHZihHzY3k4qZ24Fq9SC0vVgOFeqMu9pkKksEequn21rZgJBfkx+h8XAcxxx
dEAXJQ/RZvqaRdah95Y2mszoRDst3W8+Hl/iwlIYIklqplRWKYQusJsdhrduergB
GYEZZP0DZ9lDye1w7ueH5enZFpOeIewU4EIiDZC8Gvdu5i+tIDfKnzMK5A4EKb6e
o1itdXvhdJdy7R+97NAx6R/6Y+vF1EOzskEgyyUnjqWVHLfI6KhoCzMOVvy6MBNv
dLqjJzfI3VFxPHRzPTHtIzk/apuGNUEi8Ax6LCKqrmh9eOK5iQqD1bCyZ7frNem+
U33x9pB9KkNptisWd7mUN2GOAkN/X5KnYPf1pjpERd+lIQgczrYRuPiY2mdPpEAG
WAt47r+gGolhq8p987KZcZt8ng2bSt/tFKAp0I9a9vglvsyCxMVCjwbNX4+JuTVE
L9+Dys+WbZURyGwcUZ5atRi111+jVpeo85lX6bwkrrDOsdF6y3rbq3un1I7+CNvG
3EZk0OfdDr4JuYFVR77qa74vVJ9ye6FKdEHNdp6ciLmX9EZFcO4VlhsiaW0ZxAh7
inU4B5BVGrZTJ6CBdBZWMll8XlltZIOyJHoVBbpK1WjFXS0muznjGVrLA82S6ZSg
akYa1+lVZQS55g/93TZuppNajVgBgJ5fg2Z71Z9Jbe/yA2WA5qjRBF/cSVd0ccU9
LZcU2mPUcW9OgwBk1V1V1KSeE5jM3ByclYv3HBmcqYHhr3mjXzD3kazf79NfFRcT
g3PwM+KPziI+ue1T3Xtfxk1unUsDy9oxW0Wq2u8GDM263FWTjzcK1CPCHixJ8p1h
b294Hryk1bRWtxSIxqLGpHZiSK1C0r0GuR2vxA/Mu78RjYltfDzy3NAh4kJIBfl7
IRpgszALNss0akAQRTwgQJ5HPwHLyYgcrZ5LD0GJHUpGpvcfEkwKUj7HdUn8QTD7
sA1Kwg1xJ3gCVn+ud2jaxqcpyYSfQmvE0uTrgqgo2yiX08R3vF2WO+j9BGS1ceCo
8Zsex4tF0snfLOS1VhYvLK1RWZwPGmbdTyHDtMfr8Y8WQ4C/bb8Ypxk+RjNdZUhB
C1Ab0soRsaojsBkRya7pB3MUN/JhPqU4NCTkKXN1qIpycEu7qttRefTu3y2t5oTO
j30oyZQGU8skAK222HElaN2mRZkfLGErhumyj0hdhbhGNIvLOVrnj73Qi/HX+fdu
5KNBXfcTJMAJvtezQuzP7qsNhlY3HsST8ZjCTWddWHZuM6VZa/T/x+D03GmCTpIh
AEtq/5b3pw1OnWANNkMmm6QbdfAAHX4YlFjdBTBnNFMt9PlxESWHf0w6wiuhyMQa
7jo1aAasHFJjLWfydYO4zJ6SXiT1wAwSN7gOmAid+wqL/eYcMg0VjQ2YrbLqzpId
1DkpHPrd4v/wLi8nQFu1rL8cLz1kuNeSnZEWC9xs6MrYkozhXOzdxnVlFeVxG/mw
RK+JatynCCJynvSKyWIwUVqLih4sy0vDX7zpVH/HzVtkjq6EkcsFOsT9XmEhkZvB
D1h0rwawRUAztZC18blR8gNlFpjIiX42r4l9V128WcmbdSottl/bqPue5jaovjOv
UnpwpyQ6PKrViNmMGtNqI2l2vyP/+8uFq4OqyZJmF7gA8Ggb6az+1eWZjuNvUPBO
B5wYdIEbU3Ej5Ru9Dfqtxs8lhoDFidyT0Qn3J65ZRsklQQh8g7GocnAGgS3NHFhK
xwJUQTZvMNhjz2438YJQk+SqxsO/OONHKGj7//3y1UcIRBo37vpIgQHoFg2xi2kt
/Z5P/39Ibc0d+VTjSPVDk71PGmqeb2DtMYE93CY1znr2VqCSqCPzca/BuWYtYwbU
9ScUKVnCN9iRZWUodc5JksnltQEa6MSB2YUP5CU564ZrekZdtKNAQ7SpOhtaIKfD
kqhKjUiMoo5xvSMf/W5tcv5IgWrAqgTNGMWPTQTbEC02AUSRGsfDt52lPq8BBFG+
SGqUUTao+RpHy4J6qF53wyHoXy0U2A8gnQh+T2KU+j5SUsEfq5KWhzwtyIV5yjRp
sT28F0A8KeW4H75DHo5wmLlrwloJpWdlZns/BJroK0lK55JJlfJVsmXGpFczuv8o
HIfqyWMDf+E6SyxSnt9hrT+LpRq9eur2vzcHIuYfPNMFJGBTi69hnvxayrl0NPit
P0rUGiHrRTyS03aINN3ry7UOrM+zHRQwOnW+CtdVm+kbtsL8vNhcMm5m0/fD9xbU
H7VXzmuvJ4bp/zH5Sj2tS+1NhFXuQQ9ZsCV4a2fzpCAmmKqpleoqPyMgmdZYcW+p
hYr1gRdtSzv5nQg65bH0/dWcC5n+I3AH6s44D+WGiuWvL+RYloCeQYbZ/a24kzLw
ZXP6wxbFc9O1xWR7nZvxZbGlIEOTaPALUdUg3JvZBo9YBE9BxLWTHueg9g6zyVLj
OkjQCiH2efExwPFQbNd1DoPFoSR3g7AkJDFk8EUEDZrSzQ/wPVfCW+IPBzd45irH
KQ1gX+E0eKAJwR+iq2mfebWi0S23q/mD7J9woe2+xkswVb92FV+r37Sf1rD2w42+
LL2lqJPtA2R36T1SEEEahYbxigLh/JcfqgR5nmhClhVa/VdjWuLe1EE4k2c+cuZG
0IFvuu9bIiwYnK6k0Q49SkrwJ8STtQp9srviruzghlSrVgH6G3v+9nvtHPQWOjDn
lo6xgghWEM9GTP6+5UyjTkpvGRgdKfXorzroaZJMm2nH+HmB11F88b6F+q1nXuWD
Y+wY0RJWX/rACwlV9ddEbLtgCSg4rIzglvigY1UVlhwcuxkofNk9hmbsMD6wWCh4
X82p+mDWUPzaGs5mvyxFrY+mvGkce6xmwMC38WIG0dNhqG2llYXWuCvY+p4Ef0YJ
82oEAMQ5WEOYStXt4tC6HuhjXqC5Ehb/9TN/1KlbhfE6GC/5EJveC3+gKFfi6QSC
eIPHCGTNBJzoAMqmYdWQk9xqHJO9Q5TG6pgiHMuqD4KeX/v398XsFvNhfg9WKMPn
aBojCmwbQtYu7xj0a22yzf5aechwOh8YLbCkQbppyUTWVAbRaQKmhQf24PIPRQc8
NcBmWtczjGyEmIL/dpXtkkJVkJZ2GcEmf222HyMOLl4WVxDnON1BMvuq5BlJHtKd
dDXgW0fWqaAGp8Y1hoYuiu4ZeFldznT7Drh/AQetuaoNELS7AYx2VOFNv/jZhsRc
mAoEL2RiY5V9kdh+t/noDpiUbFoRlHWO4bUGP6S/4RSkhdjOao/bc1eCBAC/LtL3
jojVeM4yZ7GAmm56MbDuzOJBWVzS0Cd4bFzXzMWOXsHWq2HNwrfKVmHJvATC1ocP
FgSUe0etxIt9JkiYLKgCZRqXQN4+1H3eJI1Unf39jDfMQyk6m5y+L40oQxicH8fT
mPaYoZXCcHWZWasgK+4Dbj6KoGCcmtDIOOYOZe5ak9shGu22XfcjvuN+YQ6Hx9Zl
rc/t8nysej2zuUvpALWzcLIbqdfK6rUdyEae9H2dG6czuhN40FeRP+135i18Iwin
deLaCBi2odH1QJ49k/BtZORwBkoRrln0+wPB7iJ12LcdpYeieyq8j3yNjv/QCGWR
diwEDwJ3IIxTWgPjCEB2WSyazkWfWAKLF6t+eUdFurswYVK0kDU7Kh4A6x/wtpe1
dG4/QMjEJUALGHcXg5Ba4Unz+Ss6nKn7i+nQw9qt1nz7t3ne8EWaqsg4+dVUc3II
WTdpM4pZY5y0ophGdFj5c1OHoCFWNpRuQHt0MrC/qhBKfJGG3+/E6bA8omtTQG3J
e2kwo9TCWDOEtIf3oH8uqL9GT+U5c455b1pkkE1q6oCpG7B3rQ+PuBv7wyNnaemX
JatGYcmAmRRi2/Crqla86pG+bgAz+MeNFJhpkq0fh3TZ2jmi9GwzmsYC5qqx0pc7
z4YSjNywj3i9mFwiQU9hCk7y+ECsyjeTDqhJyal/7a8PvyywoNIgEt6EqsSah81K
xdSWTGgohpDyYYln0NWkdrpVI691kyXP4E215PFpDWNZisehBDuAwmLC/sSk6acn
dK452EXV/y0K9NKaLkdCw0RlqHOCJ/93vvemQSiZs/tXgzEYAg630MYQDJdkzmIC
er+BMh+aYOpe1EUG/s/aHOSdIQE6sQ8tgUXkJ6g9zWnIDk+cJ1zyW53gyrGur+ch
Ilki6KHpXYVa+2IJRPIU6ymEvmhVkGvh2lrbiYoS6/nsfFBpLd/E1k3VvXVSGNTM
fORkj8jsdbSJ5f/Nz5WxaB2Fu/wuam9fRRrJrb8hd434TlK55lxTY0I8Ytn0mHFw
qTRCzrR0zxUvwqgKxNLsGSlSXOROuJLGXTiTQ/YK45xUsUlph8M6CMKqG4yZCEt+
NtOp9DdwKx3N5Io5dJPXTcWuwN+fhvrNrXKZ2q4J8HNvExZ2f6qIJ24FPY00tvVH
bbKxqe+nsJlIDso9qqkMlO3gx3TBOOtPeZcDtN319SHep4LEnYlYiY2dKBc/PfWf
nuObvlxVQytDbp81R+EgKlbVB6rx97iPGcCjUZTrX2ihdwomBSqW3MnfgY6iSdhI
TAogAP/IGMzofwz46ElLaG2KvFoBxrUA/yDVRox1ptayBv/8p0HJRL4DaeMA1S1c
0s0vF9vg4hAjknl5PHFwroAWGOZ987tl47/azWYt2Rg5HOQ8y1MrEcz1bh3OBg3A
JZ5hx4SMXHgjSj2CBDDJXPhMsU9JbZzwR8hOlBzpsWj/VTrFAY3q6u+5sPX2nbVP
WWgARW7Vn+DUDKL2vSAvFWA1HgsBI9T0lQ/MR4jUuF+alffp14mhJpk+XGEHqXM+
iLe9U3xAEkWM8w5BZH7ws60gv6RVViXUKrM7TvuTwF/cnUPpXeXlvsJ0FT1t3r4a
4dqdJ/+Z4YqTU3I0yzmJqu+mG2g5gkStKS6YsYGYDhuAp17qAaS/gra+s0RetVmR
iWB8cnnGcrBH46JT5WGb1RiNhSHNiDgtXG4dqqQZJdxux0dmwizT6ld5OipCSnrb
BrLkWRq+y2Cjgac85OB66R0FjNE4SX2QJX0J2xgUVpx4wUmXrHkq5jWWqF+DL9wz
373YbcGrC6FNx7YpAOK2Qksud6EbGLKvM/SXAJUZVEBsC/lvL2fsY4hL+dlIb1Ck
DG0HjKrRtENev+gwF+PRgn4h2ZtpjBNeOcIPJTT2aFTs4VRh1w53m0n3ZYXgejj1
/qpz1gkCDqNwoLJCFvQ/si3UADlSxqhFQgbbBvPdAaifIQqepu9XuXNsjV7CUDXE
cTGDWBpp+C0wZVUW5mZhBYIuullLGCN9mvOFIYVolza70ynK4ST9WSHxDecMoW+6
SoKJJudhXiiD9gCNRXxj3VQLZBmyT5eFgUpkD+sQ2JIdzvXGJWSJPNnKSfJaNpDC
FhW7a9q5Q3FVfHLC1cq30+JQE08jV4TE/B4o82PPCTZ0x8wKsuwYMw1LYVyHTi1x
vCbZBtBCvTlAA6YjZxhLnT7SnTKBu7G3iAiZwQIUDG8GSi563k2yrsO1jZzsIn36
KA+AMdMAoUTsHGtuojCUimPusS1IuAOckKv1+XxiaEbJK0ECpxYe3mAG9UXPQbPL
S91ZBSgonXlMdq33AR/II9G/5Oz+WvI7Mzr/uko9eEjub05Ux5tgS4ir4OrZxGcF
0XAO5m34qxUVVV/n4GnfQhXWKdFHO74aKLggBzbIBom0BehffSWuwOMiBNl17FEd
96EAdJDiNaOG5EsLOsxRwze43KP5lKx7ch51cfiL6ubxIX8vuW/zD6eicntFUHhP
vkPaxdFxtCsoiIKvyVQHu7jXE2VbaiNbkW0hwB7XrW46a5fZ356r1JCIDSe91X61
7NrUQkZ5twbTYvaBkrsCCO6udImiW43QucHrjlLIoLa4zwoTEcDNMJjDyjtOxChl
1PZNwKx6zXscGvNCO97KwtbzAUVnAuKKAcfwVBYnQKnaEUQBqXeZrCRBSHbaS5XR
rJrZGhrf3iPQmh/ybh0F1cYGwQ6bZWXm2s/U3GzauV5pwuaNh7GQFfdh1wRfQNu2
ZkT/g3JnmhW0qnwfNzqAelhs9C1eikUZIwz5HIQ15/7F++B/AdTwmiZ1k+5oS2Lz
eYtPXg5mOeVglqqVhmzTCbZjUqlbAWy03XpmXb6wDX8nQV4teaUGCnk416qmQwLv
rt5U4uXGU+HCI1OyptX/ETCIHzaV+KY559nj01O/j8/QLeZojdYvmBDCR3/8BJnH
H3YO9n0ic43yqsFa5XHMeRj6V9hKS/KHHRO2Q/OwkC34h2gf/yDqRIxJ6zxxieAy
OTTItT0GJL0LAaUg3EUPjXAr0JZh6awDg1jZ0bjPITwM/pLZFLCtBu04tlbVhoUR
4zLbuvDjMKdW6IBQEWfMj7LN5nPgkoSWL8z7xVpiVn7Lv/qI+73mNB1r5Nd4h8/k
XhSEizbgNy5XU/OyQMXP827NyNJ9j1P/sDXuEvtR1O8yRjhw7+B6qfZb7h6y1pkG
dNwog7nSv42+g7Q95lgzAcnqC9hv2xl+DoNYSbcadDTtildXO2VjmO6c35dti80w
KXd/sT+b0GHADNuCIOkkQlFw3O+un57kEQgY6cKAbs/4o/Rw2ir0Yahh1i4wFKrA
LNURuomwbfoAEGPW1Purzw3w/So5xOeo2yFQokw8V0FJIIO0iJttICmPogk4oR/d
GlvpiWuy+SaOEi7r7eoyc6oyjqH74dNcJAnPPUN3w52WzjuWC37LtvGaMk3Qp4Gb
sMkJIgBgs/i/c8vz/turVsxI+iVRaMkfLQWcOUrr2ahBz5d3niFhhbULlMgUxS1Z
HoRzdGH06XHefiRLhVxi9Wytw8n3ko6udogspYyrlNUQMEwR/6Fw+Wz7eUkZPX3G
UJyIVN/3g6eslTuEuIyVUM8euJm/1nxfEEhfInqCOs9RVJzZuXquBG2C0qseq9Mg
t2nenJV+Oy5P3+RetP6xt/lNgq2AFYDeFeSsfSuTZJeeueUU4d+BZ9ThGIRghUjT
VeoN98Wv0NdPGhnPn/qcoBnSnA0ZU3/3FErQWwap4YkbVrW7c2C40jY0W5nbQGgr
Px0jPQKt1Fcp+C/RIluljD7wYofYK5d/ngssi6dDDZCOnQ9nyuoi1u+ZZs/ZdCKj
BfRakMOnL3YAkaWZf2w94TGRmt59ngKQ3ciEN9P29th/C3chQPsQ99yfvJHVA63z
3S68Ir9VCDVgy1hABwk+eNAEf3XsvjZgl1amYD+w9XyAQjD2CSKVKlNo2fYNhUFN
cksR7hSBQCiLN2ZEEFuMVAEFlsVkOvErnz+SVVMYCg8b4zENRXCgpODZNzvfuiV+
M3hZs1u35MYpIiN6QkYawx42YROdPjeMpYNS9vc1x85JeOhy2jTbYcGuLRHLwatH
XGYT532EUOT5fjsjTwSWtVBZSFpuHY4FQKx4qAX1VosVjTZO+QiaMPn2a8mUZA79
HXZOjeFAc9vSN31DkaNZRuZEPNsOKwNrq7XLYCwBDoVCffTxp3cnajBtY2qRuwjn
6Jig2UqnxNbyiWcm8Fn9jFq5ADwZhVGFYMkS2lbN1QV/eb7dNQcrP+4j4b6rKOUc
x1j7IkldPFfk80YdzxDCMZpxw4VsgreORWgr1u1RGzHzmrIy9KNj2Imq3N0YGT36
6W70ZYYqBGJHFVxwGqLzQeUwf3yMDAmMjLmMvXFGs9VZDwPNESjrA6jlm87zwiCy
ab1QLZYPClsEaHkXies2dXt95S6CLDzNSKL6/tQtK/5BOTRAhdTHe0ia7CfemrFd
ho19Qf/XEvL/k1PBrrjXHi3SFi0bR/A91Dr0ejUZopmvVr2woakC2M6kqFx1UBJO
oeR10cWh/BrGB5/4jb4PdjJYM4H6yKO+eeij3X2of/j1sfMS9qfUyudDTjQbW3qf
MpywVQuOzJJwT0I7CKR1hwJmU6N06cEQmRpiL9NAwodseuPlJ6glFFLZc0Yrw2q3
sxVe+S60o5fIdBECBV1JpUDXsBGzIvSVBhhXvqov9bJfS2Bb4F1UPmjPtOVajm9i
ucL70uDqopiXdmqqrNA6aCr/4heECCfPO5V2PKC82gxASu9QCuPVXO+6muD07kta
+q+xgn5mwhOy8ZcGPc1M71ElnVaCF0FXyhKEkf90S5MPYLBa7UBZQU+cAuiwsoTQ
tzYW2bLnNEc3Nt9hpvldwOOcj3nW+7tJRZyF1XI4ZWV0JYSitXrC1sld7LrJEDiX
Ywq/9hN4zQxGnNdMvmyPYz9tOptkJzSNSsZs71iHHiD3iCta7aFrQIIL860b9XAI
/5aAdPc3KYwMqdSV4LuNuUAvV+fIsTL7PeRVztmlgfjWP5QYySTcHCk3I7sTqwje
I+nI2kgt9qoEjFTM3SNumE2A25ebgIh5MVBsTFAU5nVLRNaAJGIUzh+vr4M2FxZh
7XRcEUU/4MSajwiyKzwTIq6iRr1BlTS65LnjKOPcZ1qpng020F9/ce7Cwx5R0tzo
2OUwIcNiXC4wpjM2ghQu3aLgBAMmYOTeDdasPdB+jwio63pzAJ7t4g1B1WbIeuIx
APuGr4It5odtAL7VXXXtknfj+qHXrETY6dA1ZZxSywfCrURwTw6ScksW4FTmHlV1
1ZAkcD99GtS05KQqHBaQkq9t1OaW937ke03+6MZwfP3703a8eRzB2ihJKqa+Tw5H
NUTmhWGUxSpyA/XC1rebdyzLyc4ZqnXpM3avTzR8WZIV+MZ1zn3D/3G3zDu7o6fg
qpTLm84KcRFe7jwhC+D1dGHHKLYc1Fhm+KCcxLZBMF+aeScoTZJmXKzGtIVkEnn8
xnAHC/IaJtxlbjhvIpk3KSaxZx9fJXbtImG+cEecDMaO2YBYl9cSx+h6LoqwXy7Y
XrSfBwsh8oPc6QjsmufFG6INP6l8siB7ETYVLugRNWeuJs5jXRWVLGbvEGuGcpus
i2ylzpxwvRP0OHa3j9GOf/Xh7/ixOf9v0IEpTvTShTdR/PrlMld8IboRjdJu6YQe
gSbajhYIAfz75ixMcCns0LX7sHcCIEOsAzkAgIsBBEbb+XUDesCqv8kz7Vxkw7P+
NE2wJHkpblMIvLp6ZVkbU9Fh7UkG51Rhn0gYzOjuCRuuAuyts0aMQD6lrC7BqLCt
uF6hc/EhwcsGSK6Ud4dM4ceosarE9IMoO1AHwm3zIfC+NXqMgNBYLX3eoIwM+AsL
kPDfDcdhiEzwzR1q33EAqLtgxlP9pML3hhSChGax8djFCD3a0SBstvzn7uD/+oX5
6wrw59ZhxAmYaAF/tkJMluwgfXyTLEebUwC/8LVdeEnVjZ5miN7D+/89QD/uK/4N
+DUsd9dV93V/93ebBAyeMZLZD+IHX16XFnSTPy3PjWCUe1bpsgupL/W5JyuOFwsh
UubQmrHf5FtkpD8ob03+aXozV/sWN3pkFh2qNU8mUJZbLvbL+4dzY81LHpykyhnH
MgKpwqv8hLQrW9J21/Xq/LarANs/OV3N6+eOtnPa4JuG1dK47bCJlboJCao/SBN0
S8d+5MGmhqGo0YGlkEQFR5qwvFGn4YnyN3nK7bBnbxNeL9RXkpnJUn1WuydPGnLk
AGyHigFJ8XeF17978+WpFbL8zH+7QC7WkPNEl3UlSl2MvsLxs8D3wK0oDdbq+cOq
3uUam+rxhP2Vm7Al6RCaqBRx+aF6z5rg2aGAAjpoWloAM2vTV+1a5FH3nmwdKBuO
dmcMoaOlAcvJToNSWyhrJt29056nskoBGN6o9kQ1OhU0dfvjnAl1t9aDQkU3Wf4g
KeWNF/ok4OhsOQ/OPo0DF/2CSgSaQY925vsvzzKjtVKjBZgjGreKErG6rDcDCHeH
B1UtGP9NKXGSn79puDO/RpCglb5eA61mj4R0jSRjXOwdvszR4VaXVQe2eFZOw6Cw
TfBCaDdfNSXZmpKAdYzdfPYDpxtDHvvxebf1pJszxqWvtHKzYKhC96Vn21YXyM7s
MMjHHAbWuAC7l+gpCJzsyD7bPK7DV7fBMCee1rpn/qUiwmuVQ8MsdCxcsvaHFSTE
klCZsLz7eWMpInBwh4Puau0Zj9ovURRBZavi38UCV1VFiBYqEStz+jl8HbhtUCmI
HmDJ2nLe4R6t3PIssmUKcvnwclMWjK/M43N9B7ajrly7EV0UoH5eQrS2ab9vZ82Y
VTxyCWxLcvGDpZ/lcN1sekyn/HseHd76L6T+QvoE6+oS4ZcP5HfRIcZvC8PzQU7/
DRgJV99vi1a5hWQRGZO/OtNRcLB4T6aQhqCkF3TsIka1lQvd8X7gcwk4pxFbKzKj
vea+i5cVNrPtH52shhFtzZDux/81v/BglqoSF4wHys+ndUPHkDXLDtIHsLP6F6Ez
f44HMpOdqFskVQYMj8UjkonPEuMd9iAILEw9S0klo2rqIS2QblE4bZV4lIFD4iDk
2ZevnIcyHrLwat/YE1UUkCnipEneihRv3eq73eG575xA+nIN4NfZYLFj/6sGCDZj
rP60/j6+8dWkOTRkEgDi0NzpM/CBy9OGWcuixhDyk6KtwiUKKQZra9PCXd8MDUVh
LBs8NcEoqXrrxwmHyMbNHNvV1smAz/qIdpiO7tVs0+jQZ9BIOUuQWd/D9knKf9Xq
IWW2MvxN+8p8VMYpLJnRH9r3eGlROJ1YYV8T4P0rjnVZWr363eQuTV66yPBsIxxM
D0GeTGuWdkrZij16JgN9zvMFJnWt2P5JYU/02FVJSz4TBKusSNPHvngtoeOSWUt8
y0D2FbyY4QPvM100S/YAZYbkfSdXa9QQt0bK3AwnKNXh7WVwxm+dL/IBQYuGoQSN
MBg6u5wvMz0/fcu0d/fUqw/c3b2oVyacCxKgTvC8G2wQo0aKqqxo9LvpbsLD8ExI
s5/0zMSFp5woV3ship8AT8I6nFTI6xF/W4wuP3zJcuCI/pjua/3TEDbbKaPUcukz
pZfx+tvx1n8fCMqq7fs/N/R9PfxIJh/Q9U80BW8C5EGANjX3Kz0ahj5NJH+wZ7Lb
Bfu7X+j2nLwOwUyvVIKZqQsLC4dApZZUThBYtV12ZaC5wv6Y26mzct8Hy8Ucdk+P
iSa7XznXRE9ZGAFivM9BMFQuySD4HfKtwUqgR8sUkrF1TSm/D+nzyBsJpy80xBrr
u25WoAWDSeHk5vqFpPBdTNqMcFpv35UjpB/0W2HxXzZ2LU33C7FYuKJajdbQ1H7A
QMtoLWnHAC7taVzOFbPBgGcaGNyNFUqC09D2ZHrrpHo0vSgiwN8MDgHg1JQw31dQ
Q6eQaYzVoY11AiONHLjEICFe394hfz6x5VJHQOarN0T7YPyJ2Ftj3DsoT+46izF+
EXwGTcV5rvyW19q39N684ZMftL8ReB3If8EbqheA762mtDhx8Yg68w9k/XLBIYWl
o8NELCzQVs76KS/pJ2r2aFdmtEHsUomA8liVI/Mentz/7PX+FT0EWSAonNERTOR9
efPdLFetU+nSA93TbvObESLU9injKWTK4uhvvZR5sV8LXAdxX5UjUF0anqQ9E3MX
GR4H+UaINNcjzJkl/qKiNQCAWy8hM3iumul2gi6sxOu8ovDsV1miS8WAZ3vLzEdp
X5bXRzIEj8p+F0l8UTpvuijBp77DSWcTZmiV3d2UP9j+UJ5CIkeNT7prwetov1UL
rPlB9pblXyYnigka0xe6/fQOFt2HXxoT1pWpbvMr9Bow/aUb0MYgpqoXgSVB5VzR
AvkJcc3mvjV5Y7tfSuaetVEKzqW58/rtHb4gbN29OlnKU1m54/bOSUZfg9vaOUW6
MCgoQrgvG410YBcq7qwShGm+f6lnIwLXC5ptSJUdVWmHmjvXIi1cAvP9DqXN+8Zl
v6s+7ewQI5fLRSfTZYalA7DJ9hCcPdSir1vvWZ8HFmsmkPwo52gY01FQwjGYXPRy
JnD4h8pyGiv4kaXIfsYWVxWMM0uf0TdfhoCOW+h5mbRoZj4Fy4FiDu06Qy0NVu65
YPHVMb1cWZ8pyVMSa+qSqCiuqJoUmH002meAL2iKuWQ7c4ne0kPM4m9xYP1GD6qG
ekTzeVnad0HLzMIKfvo3lOwXdBghw9o4V/cyQ7XeCEaqM19WtIs5JZFwxG1KZT4j
lZJv5OVcwJlf0zFwY8XFaSG3GY4C0FKbs2E1mzWHzKUqgE++F/f4cBnHNw3VK4ds
a5HznaX89IbuFPMVAxCVrLpPc5SkXb5EXTImRbKuIx1zlAtFxJYpVQsChJ5bOo7P
1spr+1Z6apQ47WBaEJK6v4JB2SIYzH6CaV4A6dABxeibW+4PCnPRSZiJbahEev6c
gd7SnMtYMIFkif4Wri55YR8R3rqSFmb7gO1arQfVj2WrxfvloqEoOZzmpLw/nkN2
mEZRloIwy6xnnr0ymbnd8gLdKERHZB7SN2z85pKq7Qhq71RarGPjiG3URMcjIQxS
ZwfLpGSUBomgKY5r5G4SQ2mEZaaW06FIv59N0tpb8gXHUN+GeJ1RaSPTyWI+TTK5
I7n1EHWERXnJVBcbWkts59Oai4N4Qr6Q20EM2ktpVzAVk5nMHLW1F3EGzKYIR16q
b3+P31DCvMvmJmjZYaXPA9nb4UBH89tuY1kEwqsJap7OUWkggFuqdQ+7jFMUAwXr
tUS0Hh9jYa24JHY4tORLCLRjnsvj1xYEXC7YdtZrupMnUTAYD90WWeHmNTbXetd2
cHmEkh7K7P3LJkTluaS7Qyw409L1BFX7CWAhyar7mp7U9GJgJN/baHnaAN7duRXF
3SnUdqgUyKsWZadC+vaogieohYYeOOgkR+wirsfjd3h1woRQDqw0alf2h96BDq2b
t8Fhq+MtcQeksEk9l2yqg+WwnOAydNZTiLfGZ8u5dTyzemqOUc9lYBzaYxPvSRe4
Nbp+zBzyfgiigtJCD9R73hKcMseLvF8o0LCnHBMZI20Gbkt0X8qGQz7WiAGuotj1
ygFVUkdbMAKns6ghLD1m1xk0I4Q4iBwssDlOAT39SMnbJ+xKj5f4b1SZ3Us/uFRI
B2ZAcyUuIRk0sSuSd8ORRwE9xjiEnPdW7ypvVeWRiiMr6F+OhVazBp1ba4Ar+LFl
NQxXQcZXXx3kO0NiBMvBW1A64YbDqfQFDcQM84b18XqIMsWloHD1WK0s/8zz8xe1
HLDzxUIQZ1eoWlJNANtK1wRUQpNwIwmbsLaSmaqNUA4GGSjMSxsfayakU6jVirRG
0kCixY8rK8oMca8n9aRGmvMVEPic3qqghl+DgDMMQF86xMWzw1dUsDIS5wl5n9Q3
JsOXfch1RZPFf97oVSgErbMjEefhUJ9dwLSNHQNG1vWF9yNA652JvP9Wrf4U2Btg
sPsZEqzJ3u55InjK0XF0Wq5toS5N/puHR3EkEkP9oyta7weTwarFUX4ggrH7hQcf
5dnAgIB1yY1mNoKUPG6OALJyUXMLgd7OH/20tWHX4qeCHi+zN0l6ECGWP7PBWbip
OPik8md8IwG/ZWo8H8S4X9TykEqVh3ij0cKPY9X5HVT3J6r2GkzlwfUbf494OnsO
VS9gjLQo7xqRo43wNw2pMHiEYpGhZac0vAkrNUnb5sdHBinxmb/1sBPsp24XFmdw
s42pD9w0wybFj6Er06oZe10LPa2mMCbtG24JFehTtx82ga5L8RfTTyqvirlFzS+N
EHQBsZZxaQc+nODoNN7Ciy9aqIB/qdn1sHw/hiNx6CT1fCS5thi1kC8/GWXlpcUV
sIVv2R6qZSJp/FHK9Pv1EZG+zmFaZiS/T/jN083I0JaB6gb4dharzi+qmK+jnh+W
1mhL+xemvya0mFKrv+1eNdEPl4h5ce8v0PJFmGUVEeQxou8ttRiS+22bJImMwO+C
yQWp+bj2SfUW2osWR7H++bPsG32d+/N1JtLrNyHfLNk7ODbJuE6hqHlWfqQ3Yo0b
GwiN86L0JcnbxuR0tS3RCuWPd5zULCIzyJJrInxcPY7BDeZF48QuXsPXSE5C+nXs
uhrLE98AJftUY07sPWtAqmz3Q+yXBpGjo7kk1KFE73ivtM8OT05Lh0jzJ1B6UtMK
66ISYMUxk7+QpPPm4EBnLZ9p+fa8e3Zay+UBjV0P57ndulruqIIrodFfPPzo/FNT
JxhFCl+ziEFJIf6L9ndxUoyP4E+fImlQ5PTK8/fyrvUVyULcMN+VSMYWjzOmFKRU
zpi2PiawpC1Mtyc5s+lPhidS3wXKbLMv/FzdNhALq4LvG2l0Zq+o7L6HYkatFBJQ
3UJqujahdLBsRJ/ZTAnrLkyXBqZCm+VviSwqTL8n4BMyU7CcnxCb/sTzn3CLAHfH
91BMt1H2rGtosMhBX2H1nQ+5mgdAzaXk3RMFfQxQIuQwLK9Jm/XS6UzHv64uOueM
BKL6SXaeEwL44i+8XolbIZYjiqSl5b55KEgx325/7mRIw41o5Q/9gQiG3clgz8sO
unLN3zI1J07XjqHwGMP6gt469hfTrlALVetyZnOfN8qrisMB3WAYuDRE0Zag3sUI
cBXRwGUZ5BUawircvQmK7o592vbN2gotV5smbMCjFdDl9wW3LH3qfMZB5RkWTpmB
ljns9IyfzjqVvK8SBZeOoNl7o++WkkFYhjPgvTWblXllgN8TkZi7XJ1qJzPxgnhr
OO8M+H+gdbQrZuWYCkEkanJYaRcVFX8DfE3OloCZ/3WMy8C6hNyQ6HHU3LKkWKdK
gD5a0fE39XJYhAt2wiK8qHu51gQBYVRhj5A8WpXP7QG0+0W5XVDldXnQVpLgMzfW
kUNMjAPf9h3uxbjrxCU8zrC9ByLb10xXuw+aTZ17LyPW8qXx1JtDW2XmI4wIKdZV
KF36BaVsyvIXCF+bgGycxqbU7m0u2bgJJu9GjdDWbrmn9jWhZucnS0rOaXAX1WuE
EaVc3s+2crNuX/OAmzhwvbSXJy7ANls+Kzd/4nApvMLe0gjII+lU0WWNsKR/VUmY
PplOFTZU53SGv4h3k1nhDCXLxYKorQJo63GWKuGePAloPYXVorPWcHvnVdsRBUbS
UuG+iXTRmXup0EuUcPWuNYiK+ShgYWHH8Y5jO7CrDj34G1NQG2tycrCNHrURsRFH
OAO+hl4JPkxGmae4ctXd7w+duBw2fYMULSneeRUXp55ZeenkXNyZYtWACaD4YGe0
k7C8RIro6VNvL/Tz2hz5CLuTkDvAxnER5hzaLJyXQHo2M3s9z1iXZmFklQUfwn/e
A2t8YxdhAELM+lzJTY0owG/yFmohvctKcdT4lLcswhddaD2jL4UQ/E3j96MsAfwK
Jib7Kk4Y1CRANzG+HrPIms/lnoST9L8wcwJipWFxmdEO81UtgN2MJ9EdUb2DzP7k
n2OL93IoPZ8myNiWa4qJHukZNWFqJRV4hSUWnxotiqZ0+zWVMBEFWNhvCwb89jlF
jqp74EmhMRyBvpLWZHUuwY+rnGyz/Ot0ssr4SFXHDN1TMH7QIPrSp4IgB1X6Cht2
EKamOYasIK3Qvb3qCQ7YcgsDx6AU+u7bJM3d/fvNkh3T2gUoOyw8S5KoyhiPdpV/
ynJeiTdJju54VsSMfzp3RI+I7hzDD6u4qfgLSSygnHNWVtbYpSeg2OyMammMObiX
HUD66koazJxtdoXzQjJmRWlhKzKdgBIn9/NmOw/4Ih5y1ZjguVIKHqXclE9HWNYn
gykSOyUWeqojovweR+ypPTdUC3QO+O4PA9KRiPqhOypk9OKofjjnyrd4sAc/AJQs
o7ThjCOGymATlqI9t8PvzMacJYVS8GFuf9hUOb+CdbuKbiCZjxEZVK7lRUlcn5Yd
fXxl8MHGLHBxktX/FKquEajkREJxLRKYST2Njd1laYCX+RvfHAbLUkoLbyQ40mcw
gYvq8DjkSRnxp2GoynbdzjsT2PUFOTlJJrl9Wl99aMdicz4hqw27t7I+UhNO/DhQ
SN4SrVnaSTSoeY/RTkHX5XUw6eU0192GGm7K6J3M26Mt2dGcIFzC0FYaQ57W3qii
gl5m4tBzQl4JOIq6qhEj0MKeYv1aT9rHntkij8beUI7E1uLzqXpPiAYpOeq7pf+M
M1U5wUZEMttWn6KELxSJi2RrWi783rFla9FItZ0jggKLGgmzQIJyhQXIjmZkmO8g
IWWM9+UvZfRF8Q3g/KbSuh7QH1NWqTtcJKxh/CN4aEejMZZn4JzXk9S5rw7Wnq4Y
iWfbZMkAOM1TsyuELO+xr44jM/ESi2cJoT5EXz5pRyMo0QuMOJmfeL6gXy0WuzKs
HLEIU99Elc0xTvEdp69g5ThVLRbj7ZgCANoU8FB2+wunysfJMgrx1EdaO/2XHPqC
VO15RDqWZGvfKYlu1I0tlR9W6sIKnQl/MSFqsrpmkvsCJpywwsF/lSBZKZNjbQZC
LvQkz/PrAXtMYGC7YWaL088pj++m8BoOQ9O2ief5rRJeuAvUHcrwzRBzJVn62KEg
lO60t0letBaM15VVN3qvy8B/Ev3XJqmkh/8QrY4vqHU4V+9acHmeT9j7ia2PCTCa
lsfaWFBldMNP5E4XvISqFNQiyzqJ/wOp0lgS6AjSPq6ENei5gcfgK+X/9MGeYSX+
xPCieKbAgRAK0Frzf2e4zd9fOy0Di0P0DRMlc4XhjVJ52eEE4ogreVKULi0/Dcll
g8Djx4pd5LDGfr5wBr3rfjUz5ob//dCgD7HA/v2AbMVnLgTW73M1aswdpsBi4nuc
PlVzADg7tgkGD1wrlnYRAqCESjy+SHbj5YUlCAflo6mOdN3Az7BqC0hxG23KkRO3
bLdiud4SAJtoxIGExWJhJuRxsTQtbOfUfsh7KqXQiP1Br/lPUmof82sK2bq6GsH8
xzV5MmvmHD02tYEFUjpc57W/1kLcUn6ZoPHu8W86ZLsiUFnIP5eVBgSYpjfrRTCZ
V6c9eQ/cyPrsnLcvgnf60dnkYdlxN7cwkuL2jg5NngK/SxKgzA7m374yPMCkDj7E
X/Am2pBgBldF4QLAFu3qw56JMK8vB3ZDYgUbi4a06MUYZsgGtak+EXaB4h1GC0IX
SehnutoTOEjtGDZJlxc6g6eu5pLly1nK5c0mIq91IFC/OWxFx/O/ndkjyPzL1dF7
bOitat+gcbkwFrTsJa6gQZzTRs0WtYoX/8It6qDBg8HlKIA3za30VKcIUZx8XdXp
okouFxSs61EofaA8Tb1+Tu2rKG7IWPsNlxRYDpvuqpP1HDRz/VGuCMqDUf73JvHW
FW2FgznqYYetdknQOE1Dw3hRoBhWqtqjtiKihb9fDWLq724cxI9kluBUe1XAnmEH
D9HwvDDlHF7Uc0aBdCc3GYzy/YiX7iI81gm5W/MGHTQXHNAtFue97omNW3xYzKE+
D0WvnNK1RYZZhlu6Q13MyzwWC4XBkgVOSwsa49ihBG59apaanmbQBX10oJ1/KRJY
oNJfZwnrXeVbDJCU9aWmRS9pvi90KvcNv3FjL2m5bzkOByY0pmODf4uBlkLAF/0e
Fv2dGnLFURzEl0tXzc11vi2DnqOnQCf/zkkph9eaxu8Q4PPFoxeeA6tpRuqiUW6Z
RiHT7f2XWyXys8WqXAadglAMoe8pdL0gGYzvBAKB4+b4yftU+vrKlheOhMt0HLSx
sb7iogIwUcLxYCbdExcKNSFB52Fz4lanwM/iyFmEJhm6h3egl5JL8k+69LDfRPFt
xFaFya6tO/UtZUHCnwqAjof+iwqn06dFD5dGUwuyRq5CaMlNZi/9lhf9AbYGaFdV
KznksAj0SrR78J8CS/CCLzIPk2wQmBycsPGSA3PWYDzwJSeva8fd+6/3XBAWD8o/
l4869vy4dGoLZmUjEM/+WlvzxhwRixbXlXxGBjwnM5mRuJpX0Eb2iecyXMOSZ24D
0yIMbPqAu42QCYu4DpmrGcSHOB48SavwL8d68VLDC9cAsNm/PFXyPPluPZy6iy1h
3zjKqJLeCM2h9ozhF4uByzQLPZ8cIVcMJklNPahRkMHKCTJzL3jIEK2Nk+iKozin
1z10QOywZtm+oQFcMe8HafkRE/n6Uf7xKQfbT2yFAv/1D3dP7cCIeYcjWtYnqM2x
5e+xn1jQorSdTgB7FyGGD5GiDvyLcQQZV2ntBnJk+Y99cnXwJxwfMHNXDTkUC6aC
uzqbY2xViTrvVocGevfo6eqemLNLMlgNO9gcaI4b9hZjWtIvcYdr1VrtpQUc58Bt
SODV/hB0Em/99B6p6vmfH3MxAgGTAzOzqpt4qPUvOVhBN6YAGetj7B2+k6no3op6
4c8vXiBHbOWtboyXwhFbVgggakHhjesBkqG8aJf8NOmR0rTbp0eV318aRxYJvq+j
V226TL0jXMUqva01NMTvbbS7QBJRweZwHzuasHyF6SzbS9vDygHEbm8Xb9zWNLiP
ASiTWcJKyxYkaqUhPrVvh7hTYccFC5e5Q2bJyN5/CYcB7r++cXeeyntcMlSHxwkW
ZPwM8j0nNmah21fUDEMsyCoe8wSAIhJIcp7ZG01m5vJshpEr/7M/5/PDmd+v4d7h
NWHO9Ak2AnapJOLPFtALSQhIsCeiUu0/JVxth2yHikgIkqRiXekpfnyVqMAP27FM
yX7An2t7OTvF41KhkYnb75PPNqbiIbSLmwWVgeDDHh9cltCav4nGzl/2BI45WNDM
TaDwwLLsCaUcdaAE1+3RhNm877CL+ngU/8Xpw/ClduQiDrjDJp0IXMBJwtqBOwoy
+ThKV+uC9pC11WEZ6uDuAbuhsPQKS6BAEWRj8m4ylZH8sARHUend0hNLxmO6D5iB
d/GRv/hlqKXHcnPugfLOsUDvOkD4/Nfpxk6ZSkoN9XhVNkjT+KFEzzlBdWaKHUR+
wHVqUOQ/eowff5V8j8Wv39QpOsj1O/Cz0FPTp6SJC+SHuaQLox7udYrYmJznrzD8
mSLQlM/vqE1Mj0Yyd5qUdBs1tkc+nB4x7K/allQhT0fh1rIvc+GQ0Fqhf1aaPEBo
xnGE1SYaebep3YVyize+I0wa0jJwNfxJL77Q8ILAg5Y44Hrwe0OeGwuikNx3bjH/
NVhRkbfg0/GDJoz7RXXcdWjyG5yBd/H3k5W1n4WiA7n4jm0ZC2e85ZCEwWypkep/
WZaCZichLI8mBt/Q+X6cXTrdpYkPK3rwNpX9haIdcDpFZkkAQAbLpCSYE0NAMoQe
tIGI15eEGHx0pcRkNABxv0kXahVxfFCyre1ArZBs/Fhydb4KPQbc9pb/vHQZaEVg
clTDaWsw+63C692kivDMLKHArnI0JsGSK28ZFQYysOhlSpCCLTmdRt0VumUyabzm
AL8YZmS9bwjWvAeBKqSMzLwTYPA+rd4u5iA4qJHUd1m5sw/DMjdeHacvocemWBhD
Iea8LPXszq7aW9pFPmRQjZjycS3D/7Y1I90DhIdH/ngFnY6OAT7LKO3ZYMu3MhYd
XCarsrji4GamWJtHIw4Qf1QBg5kUjpMqkbm8TE8dlt+PmUMLqQfaVZl+t9lzSne0
2R2LTuT7214ywiW3rzxwbdvMXUh/UrtWZjmoi4xEI33GfzbehaamAUG9T3NXdmvh
LbOLhjAg4nj0bWML3Zw/s8H0F1lIBYbIuJm8c2+PQT3Bfr123r5OSDnPvmM/PGSd
4naOtFNyi46sganURu96wWFmqFSDPrqQNVvSpHJOUwtuarQVwzDHEI3k5ZARyQo8
YrF1wZaOqK7sCHcqTfotv4rQ4mZPBtFFIGI8DKnJnytkbIrpC7/7qj4InOmrMbWV
TLwntEdPA9poyRdiEi8KkzQhAIie6A9S5+DqPiMgLeWb+3L0rciVuGqex5BF6Auf
oidNYF/ipFUI4AvjILv8BjbRe1YxwyIwsCugAufML/ig21d8VZgkEHmpJGgvVF6N
to/yQd/IqMgsTpsXDS/PGW6dQV1XBYbFlNhVkhaU0ROYCcrq9f3vQ1DIINBmPhRt
IaamWe8Tp9dXbCW5h+jZhZybu2yg7JbdCtNL6Z6XmOXzFjoQ52hbLh8CMjuHinQx
LB83RDjajNQp7wqMv2vc8U9ZzU9k0+V4WA3l8nA/sUAqSyiL7Frrppz7SlQVgOhF
8ItECW+TeVLQ23151+TXnh5caBOnHSb5yXRygPJt/KbNYd+dUG9ktdI1mTgFgD4M
T2r2mkDqvpYiGsKXuvwWtnwDOMO4HaQM84s5b1+AbG2YigllUowEivllPj0yuPup
5H9nZKCwnl8t3wg81jZFqz5UjEMXQC3ra2GMkpaXzdizRtkbcI2XERkkJqyZvsCM
z7NxKCb9hQNwWVQTHL9X+E/hskTPTHCk1Uxrkom6lTiTMeilxJemx8kbMTaQnO6U
V/4AbVACTsah/NAbPUr+HpEHldUMj4eauadiG5nm/KMJDbfHeVLo71PC+tKWZnws
MrIsXrsjAB4px2Zzl+1oAnXMRQkzFWdmnv033o38VZfxZEVWj9TzqaEUSz0pxFh8
k8mZy83KHlH5HsqGO0D7GsHkpKsfR79ukWoErlY2jZy25+beDeJiP4mHw4S4NW+X
epBBFqiiaAaPTMjCoat3+xrOeZRUpFogxWGBfGJj4Ow+IgPc75VR81IoG1dzQqWZ
QhYJUOKIf0ia+EjgjoVDKQCVNUabODaLcEkBH+TO2yHL8SGNOOTbotWaOY+N7aUK
qm2wRAmN+F9b52Sx0N0mHYSCb6oE3BPuzl5TOPteTun7OFRIyR9mv+uuMY2pRBB0
x5Inngmh5r3pqw3cWcrmEPocxB5KqDNtUYXFQbAIKO+8TQi+jy6L0ScHeRGtjp2K
hkdkdkkcXWkhNFaYFZoPDyt1NDuAR3il05RWZrH87B22URIUULxYehX+qcakmfDW
1RrdJQBpfPEM/H98UuUThnA8BJq9omVS41AW1DfRMun4C0fJo3JoAozpufZtS/8r
uDKE30z8i9huqzshrwtzxL3IhL4PlSHfYfxzmEgP2L+nw+pngt+U+A/HbExPaQ7L
y97NxqcRuxxKqUTnOb63HyQUDMCK4jXOj2T3+SHUOprTyofIBnYD1rApOwoiQ4fj
Wn3QXLsxNZmgDHEmxG34/ECaPUZksR30RNXRRT1NamRUAEVo3YwcGry8pzsf8yhN
jiZ8Q8ax2zRkC8KssSoUNdTEpSUWAX90WeAFz63y9wXXZj1WXRVxXLsCii0P7yGj
gWiUY2HhvT12Xi6zMqp4Kwr+VxdJYX4L46l0gukI76EPGkaSYs765+9ejUI4i4GF
ZZJp+ZLQ2JtP43cfHZYBCrz3+Nv/sYieK+JY2tH/gtfZ+VBqtH/cDTGqsQGd3UXY
PNPfCVl0s6WQT3tsXmbNxdaeNkm8yUTLnUKLkrTjG/iIJ+Uy/AFssBD/7VN7U97t
C1iqIGj4HqGIsJoAwhkTRZgbn5uy4pS8eK6rcs3+JVsNm7yLmfE7TqLNektk8f0g
fHkp9KDrBLTxJneNTY5LGLHTa0ikI5t9oKmMvKsQUGIyomdUGiM30EF95G899IDB
ZRmrbnRC/PHmQeMFn3IVGXac32QNfDf/OMgxzQmfpwvnhcJqBRxl+4S4mtRTX8wm
GevunP8Gr7qr2pGXSn0wFmcT6uOOThrHpY4IviH8NjxNwf+2qXLtQslpYR/75Bma
t8b9ch73zER57c1c3aJnZ5iE81QACSrk+KFY00uCDDkSF95mkwTlMYtZEHvivipa
H3d3lVb36CPOEFjdEJUUdcSN6sMEIIIewqZ4PqtyQoWXYJ7zwxndo7EZ2RnZBwu9
QwXwo2fVrEfmTLd/2kBuYNIup9FAax3tcoAfUzClUuGDyAHWRxA2YTOmef15KGFS
sWlGwD7Ts5fE89mgQppgisQaoczZUtXftiSJHPMi6om2iDHZQlRk12gYjMupeGCa
uHrT+f/UCUAmnRPmQatv8xw6kgy4p09OlAspwenDA4O1loP1yNFOORPpQAP9aMwd
sAPHcDI7l9R5gFWH42tFX1PFas/dQIR45c70CGaEKIei2+a5HUc3eGAaJLdVorIX
0dXudha2muVcCc1cM5DMZO3uWgMG8agS0KdKgbZoQKbfsV5jo1uL7M+N2srDFXly
bRAenfyF1mDgWxp0eRlXjduSl0O5aBUAABfhRGCbLZCqr1mdowORABdV9kqLV737
AC4qyxopNDY+DSVlX1QVCOikXYaLJPZFGg7a+3KlkQItibhIyYkzGNOyg1I8ETPi
XlNtT3WcWZbkYFbFKuakiaNc1xTUSWgas70w02gN0oAxM1AuK9J270DBnOea+4C+
HLU2fyq3WNEUtmOmU/Oa2W22Rk5SCm4/nVD5brpId7XAMWuFczxPts9tnDmH4t1U
F/nrmLEMlvOGHWdA72LxxsUsH5D3/0afIEdOjIh22liTx/2sp3BQ3BQjaLNzTJLU
KgwEm9F50VeBnmpSqdht9hCtP9fpZKf9iMK7RpuKz0zmd4mzkGWCSkcRyPFpl94S
eM7Oserbl0hAGmIwBo5FrGx6Rrc5NDTBpLrbG1QcS3e5yPpqeWwfh+kPVVWv1Jcx
VKQ44KYBL6PWMguITFn0Xn3ba+h+cRzT5V5QMO3lwcex7FyfeIa+UvsSMrvMukwA
ZADoq0LAq0rtWtzh5ncKuWlWXl9vy78BpKaTswkCRvUMSMBDdHBqdxY5kex7fc3f
tl7OZxbLgNLLRUzWjVJFL+gt56r2TxKXaEXJ93R7+WeSGOxmOYTohhkRYqy4cpft
SvUnDVwY7ojcJd9au+jj6UWcUiihiQVMvVW9snrYLliLOKREk8Qy5hKjglqVuhDz
Onp/CYwFrs6cX49rcQ5XyztW+o801djSKSxsqMsHCpuweimsuvWSm3/s8R2REEWH
h4amo+0gk7b6KkLwHW14MgHzK6HdKvuI+TvvXvn1Z+Fhk7DQcfSdUeU/T4i5J2EH
eYtTlazuOnr8E/jImqbdNcQxCbikXyOA1IrCgwc6ZK/Hhkb6g74EuHAyoGBk8mW4
4oGwgvSqJXScez4HP3gCr1aFLUnTx/eL34Vmgrvdie/SyPBUUwIPeuPZcTLUhNrK
BjZ2HG2sqUl+NY8nA0kCYlwwiTTfiuodU4OdR63ngTT+ZVK6lMChPGzl2TkFWtw8
b6Fh8pEWRG2aRdJ6n12p+yPv72UQZZDuSJEIAMI6dNPu6mbs3iJOSQm53kPYDkAK
A8D/OleBX0MuJ0zSun9jeDrQua517DwKE2fIENituBcaSfYNV85blBjJAz8H47Yg
T48nqOPEfTOCSJ63G5oxKeSIWkHS/xz1u/hJkWjW/qiJz/NrN0SKqodjijQCAkie
ndrYk97LEhEqbtvEjnTosq83ulJ7a0Rj46EHyW2M5v1/bsa8qAGZx2XkuDFjyYOb
yHLBTB2VnpUg+AfDZZz2zsquzUuqlFIpUgoWBkOqy+0qvKYeH9cc3DlLGEsz6/sJ
N7iYrAPbivHndRiHwPz+Vx9QdBn3FznkCZXP85I5mo7JrH4sx2HPxn5G/UqSSBb9
c5K32rgRL+qUNU7QTJSpGUXtDrI6ttDBjr988CquB0ui0Tbf28jj5Ilb90YODXMN
VDzyQVzyd3K1JepPNQj3AWc+Tigsum63ebAiv3Mg4XiJS/cvRfcP10/31CPWRCjx
+rlAIRJi45mya7v1b+9xYpDG6+UpeVhtscbzcuMchO+uL8KsNOYzdmUpq4blGIyq
u6J/27HN4/qLrsgE6Oe6M+ghXyTS9+jEYS4z9x1S13/GTa8Vqu6oJKVS1al5mb36
XICAB54ymdR7jy3xo1KCS84uF86wdo5TykJfT2mh5ChEnR6f7pnBacqSlMXFWddg
3oAHX4yC2+LhEZ44hNfGiXjG1ZVzyre09Nh0r0HM6jPnnTgv9wzoo4SG4zkSF47p
PkNd/GUyJ0q3O1pgnwXz28kvu0G1OyCp6GrhkdC9LCkXCiz7oP35TpVgD34Vl3wT
ggAHTOo05TDpzR7jIPQNEb/Zrte891LL9Ex6jqQjMf1Prft/dFKb8Y/ObQMhbfDt
TPYRPV83j7DE18syN1zla7wRZzivS5hoFUSgUbx8qVwyZu+n+Hxzn4dNDNvFPngw
75EvZAIlH+ffNJgI0PQFnXmb5RpsBRblZiKsJyKFyV1pdXKyJFZUnliWvNXc/TBc
QIh1oNv2RiCsIOmmC6SfHu4GLXdv/MPSapbmgrcsHtjRedi0/X41jIwJjuYRmIE5
zbn/5acxNlXTAUO24B0uXqOg55Z78YS+9EnbPY5Y4PdqA/kqPShEJqqZ7s6bOH+a
J+eD+DXjlsRMoSk+qckYlt8VchIUO074rjST5WOh8iQa4eyR2u0cjXWfVL7lssB6
OSL8MFgfTWcHAh6fiwA6mdx2YDglqSZVa83vbEMXQT562dc78SwaItH8g2vvDKdI
ZlrPmD1OQ+B4IpM5h+Cp+TmsBQTxTmTkfKPUKHlqf6/SxvTD3dJEcRtcAZiZ+PJP
QoQtN0rXEism7Ua4UdGFylHxKs6Aiz2SzSOdSwcdu5GaYiNqJVwQRZW2GGn9q7lb
+7QtB+eGmI4oIjqXYh9UkmYr2TvzEB+mylCCydYX7FWIyEJIwCSvj1xGdBiMI1G9
zZhLycmHHtm3veeHpu8vjR31ydJ8wQ545SDx0I23iZ/hgr66MUTH9OKQAJjrlkSW
Yso36uvHviW2NLJc7T0erqui3sd6ALJynL8gh8tQhWKVxDoz9I9NlgXqwI91ELct
UO/Dtv3p21S3ZND9OJ7X5OBBEkn/KHp++0ZheNaYrIe2Kp8S0okWC9fin4K+9UHl
eXkExSVRNc/Vjdhqz4P4l6QWl+0YcyOIqN7xb+Inl/3KYJpRnLvai/mbrTEDlpXB
/cxLsd7MQjCLzflC0NLVBYho8ahZFAuDU2ctgJsUrbyrCjbHUAdWs0Ws+48Tjaqm
/WCF88EyJ091RqxdbIiAj5usvtLyclbi0yT2aiQnblS6UyErrS/czeBGcVqDWDJ9
0lSmkLtHId+caKc2P18NGYaV4PMLoQk/9F/t0I36exBM01QfJkF/r9WCMvXhYf6s
sR1FqEzlQ8RoNqYV95wetKAdW0vU3lTJq94vhz/t6x80UsuGCM7fAh70HyCZdUfT
fjuQ+cwoYJ0IZu8GmSgYiRTxsWCuJs4kFtaOyAR72za+7vgVl3OkzzruqAMdmqcr
hEJznemnNk04dMQgh+giXpS+JrWBzHxHsVkEowB8V4NSND5ra0O3jrKUIVzQ8hq2
KQ2LfgH5i/QInuLme1MldwDQfuQ8A2pvefUnfhP1otb5scIyUSf5w3yApkUZLjur
JvNI34FAK2ttVwuHWnwLwSq6jE4bwjvKKFDf9K8D6lG0hSfGcXKQuuHOhBpaAca5
Pd1HuxXZJA1k0OGQ+JpuHO3a1KQo8D7PavmaV8Hwq3Fl+/tFNLIBwhlifcHejMyw
CTd9jpLjNqcMfThyfQIzRvdPlnnm7F0Ut9lbI3SrnHgGR3YBkE5tlFVwq7lV0dkH
13x5ozji/fYYJs5vZ+JkBBbve5AEglFYVVTP79/sXrXVEz+Ayhf9GPug0DUK7ocA
ZKb2BBbQulTmTYLDo/rJytk5T6KrOFMuccmUaYvfzZ1L5HoP8P63RGsrVPOmlQx4
wItZJvHY5RmGiz97kUvUK3kBNoLWpPUP1VpjRSGi+4lG+KquvncnHPFsURVtSX6f
opX0FydyT+yAWPMtbXLJrZsx3EX8V6u2/F26WMgsfg2DbwgRBO/+pq3NfrYuZHV3
hTSzdpo96DVGovkw/0bi3H48saYlhNpiuFJd4mqRBVme8uQunQQvph05abH68/xn
jwgsoOntEUN0v5niYwvnqH9qxTek5XBSVXJjARIXTk7dDO17uTK0kI0+h9jF1Y5y
zB+zOvCpQ3mApX+17RDzLi5sNgSVoo6BOw/nUqD1ZTDMpvqgQryrdyUkxjB8twCR
x3fZA4/l7aT209jmuE1WN4eQCySMGSBgiDj8CG1ULlYcVzDOgbgd3/8ye/KUYC1n
0niPCWABUoud4E116PeOKfIc2a7ImdZ32KuPJPM5cfAQrGmdmrQ/yc/qCrVIXgpm
0MT0Uv/l/jvBjaMppEvonE0FvH8BDO/ZDl/7BEH1Tu9wkLyTkF0v1C5jh5WbWzMN
s5jXy2VjvrVXJEm4qPldj+k6+TtyWDBZ2ZOIcTAIkuOsUVOEqV5dj0SqeO/V+KcE
Wsqafpr1U/n+TdgvwkRr8odBDiiT3dkckZRPDP9S2d73KnLg+II+EDr8s+iiWJem
JEWFbH6p/4PbKTSSMXjH4Py/0ESg0U9AgynectWgukR7kx3zB4WxxCpA9VGw1cIA
NhHX/d3x+VFg5Mj6fdlw8lo4BgRh8CoB+VFSavS9Ho/lV3wrDdWBMHyhc/Wv17ti
bvWgJ9PwmBaM+PAEDj1s0vnUOT/km+mF6qY+HzOO75BY9WwNEWdsrc/+YRysJwOK
11Ttqf//rFCKVrJi7NBkuU5OtvfcAfFcQKzLBht24SpG/FnMfrAn7/TqblCR6/w4
xLQIJ2lILHjvtkDoQQQe2eeZKHtA+GZIQfsamvW7zuBX3VXXUFKErxg5/sSE7SFm
hqVh9mx/TRfigXXeRd55riet9o0qDFynAMC4WgYkC8WBKUG2plss3B8HXC9rmJyZ
bcX9VfDSPaA4iNpYeD6tgiHpbxQDLyHMlxERLPANBvAth+vu4LNCeKSWO9nijeud
0tcNvMwWpcAWk3ZKteLKz/1/Q1YzjQvkIbiqsmrTgyJu7xWlglIlBhchXLfQrq2/
gwxsYcsW7OGYJhOLgafXpY/n/yNa5fdlcUH0s0gLSatCMwwGoQfEF/3YEXb8Lw/Z
maO0i1fKzLhsW8+n8WlQJ5YEzKP93+xcU46O8iT8HvqHdi1XWZ5IgLpTAyuOg8qq
jQLg111uMSo0GiYGeZjt/+r+GpFj/yuXbxjmgWejhqn75/zhJatWHAmsUNYUo+UW
i4OKhRSLR+RiwuSoFRKx9H5/iINcZQOYmlECBLITlcJrVPtaBePY+VGnIJgYjzk0
PWVB4i/vSaqtu40t3f4PnuHlZcR9fZtrWZnZVrKDNHyGKz6nEXA9R7GrbR4+DZRL
mox4n4kfm8ufeeawxDgtdAJoJqPCoo9pWElVHVbn+aT10hwku0AybQmkm6A7YnaR
JUar6dQeHPc5t8qvMkofUB7GgAvIOoY1BcKW6KHhjOUfYhDoI0P2pDlaWiPjT/pK
AQbUuSgsij+rqe4I/6vWG2QiuPXW+Voom5I3A1FjjIwkC0Fz6QnP2vJ+onnWjK63
xuWwVLnP9tTefPAeg7xlBXUeETaUqeUjV9/J2Zn0ZrbVNySVXgfA1JFbHyLvuxp8
b7wE1lz4yPrVPBSjgRYPhEbRh/JmWHVXvBq6fBvxNaPKonpqXd7KctGIPzG8T5g+
Td2tkUW1lfjZe0L3WE7pcRy/ISY4K8GNBgKDGiVyKrzIklsU7zHoRMsGhMB/QBQB
BOXoOl6itKgevFzIAXzP3JKQSSM2wAZAXj/aMeHDYdT1QsTh9wauhlikK5SGTPMJ
CQsBhuIugIjc3H4522DTHZjFEQACXo3Vkr6qvQ15ihPBmrRrxtXSd1roSpCbniW/
VoK3LA7B2LapYCD4wo2l+KuirlApeJ3GOvp7zMf/0CyrQtOExn8u92sS6amoypvn
66sRnEiGIDpQVSlnNyP/VYbm/3J52D+UMbsDfKdTCDDDQnL7UnMcNhHAXpHnDCzI
8x/gcEAE6tukwYlU/ZgIyNlxYeuSMMYM1zTU5314rUtzb44xECpeqZeDFDAci7Y9
68vZ56j1rKH8XRUGva8qbNg4DJfIa3CcLVbZAPv48SQX+A4NSuWjJu7KXs1s7wJP
dSYH/E2tXOxb/3YrfdaK5vKLaPyg1jhqnjksPspNERjLbaKB472b4+klguGgM6No
gkNYnssrAzyBs//6ROOthvJH3CQWg+rbUeKS7IB9OJSu9wr/Qpz6rTnf9BQutSPm
Kock52NXyXL0/8Q5fuW0FmFGoYiK8rGLpBdE/HbApo7Fzda/oRWMNw2idz+n7uNS
8Vikb3ojAHc1WIN6NSjuWSweDKugU+w/hsgO+us1AJ/GMEqjux7L61TlbP2uSC5g
eR9XiFCLa6X3elBm49WC0Qy7Oiobu78EevH9FwmK/ipuZM9NWIyUk5jo/3Jhdywr
FtGIYz2vIYlRggRxkk8teoHePTG6fvZ4h4UlRZc6QvkzSVExc/gAkfGye9jiWpXH
7dVPQyUYX6nHxlnh0+0fmvlaPx4uMESgH1/5HvariYkOF76kOhJex8ZUD/btVqaI
31UlOvyvDG6wpMSqhijMlz83gj0tEaIAVRqvad4tl/FlKDDRdOHOkTHChvRl16N5
j2syG+Xrqt9ywkoMPK+5wcWo1WHdqc908vC3N1zuhJac0Xkt8o5Mw/65GeZXVK3I
taYt4EqrWwqu88KGMnlsqo2kuZTNhj1Ny0OfjX+ufF4hIZLFXQhHBNmIAuEHpsTt
bDXNha/6hAUZIC9xGEWH2igOe4xUylhennbSG9/KOLFHsIvQaGSNXeVs7lwTi6AX
L9knmSgKWJ8iQOpqXrACpRi15KfCw0FCTQuqgi+KHou0LxPV6UU3lFbwcFfkOelK
nEbedIeRIFcH0yLh9wJ0+1IqH8LRbsRXIkuACRoWkO0ouL1sY20XY+kHjTPhY92G
JAZ2ajYbHbnuZsuB8j8HAYFu+FiBcoGt95IemWVopt+0Er1SrQOvSXUfFmUSUvC2
LbDmh3oWKr1G/Z4HOb9BjX4ntxcx56VmpTBS+YsZFQxr02ggV8jn8hn2eYM7VDQu
MYRUuPzxGwY14gDPsbHqytAH2hlvgsNiWUNXTzFgsb+FTRdciBVslDf/EZGzBRQN
8bQwu2B4lo27A5mGRGMqOQn2JPobStf48sTtOO9vgwOxfcEoaGAbFOloHGiRpyOV
FMedOetnm8u1aFw8BsHXnhoU3flmzCb4gLflmBjaEDJ2n2WyyH3lhQieTb8Nnxss
yRJtr9Wu6AJ2VXHY9TsgTJp5fECqBQahKmPjdvDzH8Qav9XOCcwJKf5GIKdHoE2i
+UfMPV3UTAl8Nt8PGuv4GTk2CldxlaFWzYr2b84LGQdUBOgws6/qQr7xgDWFfgN5
jXTWyy7HAA6JK00r9lEbiV1fJGacnRjk6pFdhBBthrI+boqhFOcwnzJPlVnrxiXa
G0VU1fDwMrF57KvL6fEK1M5JqeeKLHY5luQh2mIi4za0CY94rgdBNl8YvJJ4zVA7
UIklJ2Za8cZ3stuU/0VbRY0DS99mymD709Irq+Xa8kL4C2nIuwpOPs25Ho6X2nGO
VkzPjtGzoid2G2YtbjNiixDqa9+xHhMaimTZmCGAQREeIsIz7UsM8z5rAPhSugAZ
Ep9NjnQSvLjehJlro0Xa0Fv84lV0elMwrEjs91+ivI6SOGXHApTlU00naNqnlNBJ
L5Rkst1HcWTd3i4BR7RqJ6owoXKEtb4l59gDmTA90vJkgiVbzeum7pCkvReRdzS+
9zTqfDIVoW3Kis2lMK4c8ny8s4/bERlIznv3drUIsUqVwTpa0jWQRL9FBhz/Hh/R
gkHVg5BmhR8hv7qu6BcE9oU6ido2uhxXHKha9WwcFMBHmOyfwV+JKOZf0u76Z4zD
KDS9DI7zrf3H5VAfIjdYjuNWa00FfptC77tVOeBtMKspjjLARdMAgslebdHpCiC4
VjKQzbCWUbSBcHeAf9G2FtoOSZUMeQQiKp51YrJK8MiYAXIjnHmHQ0am1Q3SAMmI
kwcCUPpu5uoYnzw5WVGkD+rgrHmoRgc418DGEDpDADKm6UJhLSIZYnonDV9fV2Sp
qlS4Rzlvt4eHBuvTzYoj5OiK5qLpf2GEobXLOfV7gDTxJ+gNcVsHHHx7Tab4lxXj
tHp6ptNLWJsrJcLe8GDP+vfSfjhH1ojbQh3bclc51S89K0XRRSXnfn/gFjToOLkM
BFajx3no0aiBNe9HSEGkAmnu5Atqe4W2VbkThm0Qtbkuq+fiXm0Ne420F3A6S5ZY
O66y9bwKBi6Zfg3pxgLz7vKBhOEjtuuglaf7EmfwM9t9yov2e7dwZq4WAIq3QZHt
N0W3cPzh8tZQqGXPcNmMd+nRFef2FR/y7AuFORHs8O+XhsrJyZKgKRta+rhgPOgw
QKhU/H2RVrCxSUluRC5LBt80LbgatcqtqSYJLXpf71TThbazWYCht+fI0giMMGa+
bUy2agzV2ggsx3T0OyLaa6EDgjaM0HmcENuS33/9OKOJViJwdvkyCdH7I77MC8Cz
z6sfWDTeXNkltmdKD0jvXZgFAmiNSGATFDX6plvkS77gEX4Tpf2fgPIFNeSyVVm4
osVA0OPVHdlI/rdXoEfM4rEUfRfgyrxWYSjYJZ0rqaXkCeRHAo7IKQOhb3Wxl6uv
hm2Fo/+PSyLK57Uzta/l28iR9PUjiZeqmJ5LLRMABbch0Tmc8pSWGC4OANCeIEKa
Jw+xbmpKGuQ6jN/Jr1qNiWR3OweGA7t1Ya7bmcM7x5k+TBTdLf0A8d6Vvnp4nmZK
gxuNhRkcxfJENvtDs1McFNVoCYqArE8K8NwKKcKb7813myhnH9ZEu+8rKjaYKapu
6mq4R5Qutz8yEWR4E7r8knLgWGhj0im4GD3705FA0Wu6URiVA4GjxUBj5zkKJcNc
/Xhts9OklcqMqBoADksf3Hv4We+v1ujmWqgc2Z+tX8wBKuVaFNpGnoniPjbVfsZa
siFsdZi62IRApZpZbR2hYZGY9I4sqVaGGXM4vAAHDpwz9+ienrKVU9CriFKYRnqK
H1pbWJH9P/+XQUQVTfR087IyJLA1CNDAwv0egXmUG8Us6BJkffmL0lo7Fsw6rczR
of7E74+txk96SI1NIpLumnmpFh6HmsakdKr0YIaOPhnK+yh4PB3Y6cmp7VZAQlMY
rp9IRlATm9lu+F+wEuHxqCWIE0vutulDdLgMO1j2AzlX2qj4u04KFsgnpweKCI/n
GTfP5NhgRlg4xO2xev1JpUllzeBEPDKd6lqSloqGdWqD+cVAnTxQaLG4g9zg8oPH
n55lq2GM/2o6h0hxzMFYP+EWqLEfMG3mYn4ehJK5olvWUMxuExsNO5r2Wd66unm3
k/IuvxGr3ynK2KkdSIeY0JhZ92QrlYqEASXg8MOZ4ifN9IknXkWS7K2LgrUen85z
vDSUCr/7uLcMBFULDI+Czzuqc1sp1W7/oZtRHZ6Ar6uCMGG8DQuzC8XukGnz5PA5
5f9l8phE62ziyilehOk4M2ErIOGH5p8CjJPgzG0MLwJdSvY4VUA7cPMOpM7EhexN
68mU3jGTU2J/XjrOSJTHtlEgSIqAAmnM38m1EBIWsLucv5RD80MFAprOIOyZNx36
mTADogZcMeXu94gP4v+CjYcUJzPJPWbp0EM5PQTu5Fp7ZojVgYV6YVKMuuCOrAP6
PpACjR3yR5WxbdCyvGXnDrerNwye7+18S1STaGwA6Wrc54dwOE6xdfY8Qj2WO+Q6
O5fxgPHQOvgpdhMF6JZUFdkfpSY94er1Dm8Al5qCQjSRNaYyHeMNrWC82/OtGWwL
5cGTq3KJ+t7Z2T5Dg8Tj+iszE9R3vbNXi3imUSW5K8bOwdDVMGDMQN0VSMVxKvkm
pKgbN2s5rA5j7Bt7QjcXbYlVxsJP42Nuww7n3Vx5lduohLd9aA62k1xDreQv0K7c
nlc+sFQvpk9hARcolEhUibAJ9fT7K321DPqGVhs/RCTp4sbGwZQwD2jtvJOprIgO
Nzdln1QOo8D9EGEjkSQsT1tjuhuB3l2z+bGsq2px6FEpTLVKrlw/h1tSzBUNoYxV
KYK6hCp3LuWfMoySs/Qs4dhd3r19X2ipbOaIEojzqPXrc06JH97uJ0DYCiGKvugb
IPRgTaeMa0i9wGjBiPi264R6l2HTwFuKBHa9BJwqS3R2G/hYEFgR1eTEzbA8hXKS
SSNolO4hupOib2SEzztJVNK13hzul87i1t8IYl776srg1fy2dfi16Bww1um5PTdo
VSDfIhDgP5LOTEPwjwTNcEx8q+zn5gy/CKblVekrBHPjeuhfHCD2ntipyiVz9MCr
6XVaAYPTUBdTpUUHnUt9d24DcQLK4ejJIPHMkbxdsFVV1HmaNSY3hBiy93ZQb+nq
zvvc0Mm7m0qZ/kl47A17aw2ijs56V7gVUKKZPlV6/aKrexFnKOHKqtCeHfRFR3fu
nhEP+nlV7OsoDTzpAsPw6X/knF/MWi7hR9q1t8D0zq4sgom9OxFtMt4/q0mOO9dW
V96AwVaxwUoMyT0IKyWTrUYw9bFmlFCtEx1OECuYjynnI9MLhTt6iZmswEr5yjL1
RnRTKCYDWqO9Ch4ybSNdDuokPtelYAULYriX7Wf2LH7POdvPM5YsNpmqf4ZrW9pp
XD4H3/OxcRx5n+/pwh4K68p7RrUuwba99VeCV21/VMaZyviMJNWcBCphf18IHJn/
eVepKHd6f/NJWjFQzBRgoRPnTSXRV/5BTbvP/W1IdQ4sxXuNgY8ikh1tUiGMq+bx
fBKTxQNkMAK5dKXAakMbg8dFSyHWLtewP5uYhjF1y4SqWYpdNyVgf6vuSqEWxYM8
32wHRKKcubeIX1hU9n3epKnaY4LBa8ODenQPyICtbrZImv+uYsaTxNPX/da8Hi6U
PwDF37eoj72kOxLI9FajqEKIj0StKWQQDBwIGnPEr3v2Q0uCKUnBgP9seBVfBAmD
qLZwpKGueTlMFJ+qpMXuX6wlv+xHHOlUXRDHeVqrsNsYSQgDVXbnKCrRSvHSMZVi
MzoFWecZW8XqkHgpv+Uwd3VcgIY9mDYRn4qOx2yodJLMkPalNy5ixT/lgXSK2z4u
5W19pGOc0DDhpJ1sSYy+P9tuFjENiGIR+wqx5EzDEF6AzbteAF+Unwi9hgIy8iQY
zh+hKF0AnJK1qU4Uq7sTIHHPOX3WH1ITa83JVV6cFnDI3xQYhoSpEA8HIvCt+JQR
OPitrD32EDXWOmmCYe+xY8vqiVnareGAeg6kOAsZ47eAQGRJnNkgg5o+SVRbzKiI
K0oT7rvl6opRakxSF1dZPdlxOE09kPAY3+1z8PWZifPYFC2iHsjp3lCWjqavKroO
CPvEVih1f8uCKO62Zr9BNm0CgX5SLpY9xmrr7p1GGUQ9eoM2UK26QxYA9P44tF5V
w7lTN9yQ+E1badKv72de1IBhpcE0BKcG6bC91y2bnDRzAKTt2Me79f4OKg2xqAD8
/prk8oi35SvvXkg4gpJJOlkc6IeMOsqY2XIFAxwf+eLhxN4Y4W1y7MhHMyxVegCc
v7RY13JLCjnZtSXUR1M8nVnWmwlIHDcn8NQ2aF2T9gT6igTme5DBux/7bmFD7V4l
G77x7dsrWX3gyCNBzkS9dXbkP+MVuSiCKpW4Su1s8knAF1y3LBGO9FHN32/Lyjhf
q/LhfWNf7Q6we3MnYQXaXEJmomyqZLy0S3p6M/iCVvNNM6um4Ht5M/hptCiGok0D
96w/MhWb6JDC7wDcuxkDc1lic4bC0puO/wMS1bgsxM4h9dz0ZOgWYUshbQuGytnV
u0O4y05UVDrxNYPrNDA5UX20kWP1UnIFgclhOuNs99xI9EPQ2k7BnXDfaD7IKX0t
j+cNVtK3iyUKRWDjtUd4egdVxa//8pZYzmGTpTn6Jel1O1nV41ri5fX7Y7ixsvMh
CNL66QQO/AkNNc3vm4uzI2irL7M3HKVyb8/2bxlLjL7wzz3VXkKbGMmaLwqPJ0bi
Y4v7ga1McVFwDMfPrsQ06VlbfaCFoiy4Gaa2A1f0IZ2/NQMIZuiFRWh1a0BFc8hU
RYpd2xnJAXj8kYVhby9ma5KfQlpEm/0+MUMjPRWxemWBeaUtnpX0uDbQh9hoScyo
0qaiRqvslcej9N5GPZqwGEI5WybjY9ZUX/rMa+Z7uryvBi7E/vQloKPbwZOSTufE
THR4sH+iI2h4mutsCojgKTa4EZmftWBFbhpW56/JoArWnYXzVEwxQP+4gxzzfu67
siy7efkw4xT0xa2h+acD+Z/Gz/q9DDC8zBiEbJEJJ0rfltQ3ryxhBtqt8orEnE8t
iERvkBJiCly9giD2Io+YWQJ1XhIox1yvDxKLbzrzzZS+LGBt47DjiatviLpgZ/2t
rraEkiegL5A9w9fuLnEOvGSIdyO6nw/h2g5s0BkNouKZKlHt95TjiFjn0Y/eYG0x
HYHDynYdSUv6DqXyI3vyMro+mcNJ7un7hKPUHjUSrTKTEsOc0Tboa5b3MBVbIv7N
uu3JxrzNrpwIERjT7mPMGPaIgNvEoCcEpehAvedgII2iubqnnWw0AO8Ztu8zzYyY
ZuMrS5FvauLDOvIfAZhCyPwk2mbLsuBGr+RIB89xoDC0tjpeOiTjqY+xnyfUJcig
5c30U8Swh28S1vNnKlYLc1sllIrtCH1nOVuTEDy+WTBWN+IAwG6MFiEDX1TAip7p
W33DIsXuShpoohVc16yhhfVrtxNxmEojTlLsvkKHM7XQHCUPxZ17NhNw2xOr3jOQ
IJB5Av3lQ+XPevOsaQlIudyLkzaBuz5Pz8BGDttznLvkBzhT6+rVwMqhE70NfBje
C/ActTLiwJcyJvdfdQge7bpONV8MzFynJ8exWNwJEGe/zoawqj3qN/vlEnE1NeMm
Xv+jDr+qbCAiKFHLqIMf9vvIsWRBj/KybjtKcGZl+m7ZiJF/IbWsbkRyvzBbnj2A
XkbnpatuVvbaTQMjDgwjCDuoI8hOkbPbwZIA3U1jOGhPHHiMDAqPtgrZN79WGqfl
b30FBNo8zo6Tgp5+Qbkt8cz59JgYaqWcvAuWt5T8KvW8u2yhp3T1MG+3I0b4F9TI
Ka+u9rrPwe+kCbdt+2pn4OCVPfAMU+lu9VUU2iO+Y9T5ntIINT56PaGHuiU+5Rcy
Mg6YT2r4AEnEeCGWzKonLByQhiL2loAz4cDOCtjU8LoeeqdfeKmbB3ZqmUshqV6L
zsr9jCrNICVLBWtoTAvgZ1q3q9xz5wP8NEU5NXy62yKS/JGv7ux3t3pmDLVVcRJi
Xx/mEhB7jS332uiZJKTKbf5vfQwKKom4ac06DB/nGO9rKL2OG/gH+kGIm2o+X74s
+6hpn3kzjsG/ib4aofknASrQ4tqT3qDHkwzmscvBdXJRQOaYwIBUmC/Vp8Ga+74s
7k8kf4UD/rRqQu/xoJdcuncLehUMEKN9fayRcwuK/acpC7GStUct2KJxpBaTeEMA
tPA+nLDJ8JBTn9HYWYKcOwiGSJa+9aqNmbEjKAiVPvMPk8eYCb0Hy0yqyKJ2j4Lq
jtorcR54bCZMM7xQglWds5++U42heDu3/Mau6B+bleDSbJHXs6C+uMvDcus92w36
aEDeXEIWxdN8qeHb89+T6QDG7RFmy0+CWaPPmqITpbhaIsM/dzraiEky+1tdl01i
pxdWG+sw8Jv9nqHqfU2S3j/3cojETmLe7hNdDoqCvpmbnJ7a8U8+4um+SBbIwh3w
5wZ538pm17xHuV77AR7AOZH3D7fIxqvYKEzlTUX4Q4S7dokChEv9wkba0DnMAr0t
iMtKRQ1RpM5vbTu81mb+lpiJLL+y4qjKO2lsaiZJzSdziuteJEW9oHscWzAXN1dN
UFrS81gmrS8pIkS73rfIGq1IjwGK9RuOWEurfURns0+fiyhnaQ4XT+GQrZm3FS3+
RszvR7k9m8yFeI4dbXLNb/kP3YsJ1MkNNNCItGRSDvz5jgVDiKacaUJes6qKpZCg
RCn9geSWspLgRA7tlNUH5+QAPC7uDjsgAfhwkXau9fnGnvHVMVBUxQraWsMzY32h
07dR2QZHuWuxLuRkn0v7B5qHgkbppypM8pDPNLC8QanbTV1wJW3DDwx1GSWNT6Zb
SucMm/zGaQeN2kGL0n2+Nl268J/L2RqBsdp1strceWAYikx7h7erN8Lmd261EiMM
czUpl1b+13HOFnBa9kL7qhQY7IgGM86kyLFfnoG8bNpUNmp7SFUbSwBFY99R5ziV
jFpjhTC7v45OCBeZxVCKUvYTXQJCB/B+8KbyHRokCU30XhoDdyE+99LZX7jt+8Vz
eRkkZrhpaE0lC+4vgV5EL3c1aH3r2WkwYbXPhfzUsjS11rG/7nUK1VCJes8bEXxS
XxAYT+DXNn6Y43Vh9j7zIKROmC+Qz6+2qpVFmwvc94Tjow5S6/1CaNHu7PekV0Kr
7mMKsEvOmLLCtPjG4+/0+QVS7OU41x8bp8P2GNjVdNFuyqWofesSYaDX+lEQUjA2
mCJNK+l2kqMMuLdedE00c4trQoo7GjWn/RH+cvs30ZmUvGxRwv/jNTri3DuZhW48
NIyhNtaxWuHFKF4wOv2d86ovHqsa+N2ms9NdxOUq0CgzE/PHceH26tzLzuJQ5ZeV
aH+fJ9z/RrggGRP55QeGD884rPuuS+O/KSwDR9yi8NbqU+Uy7ySYHF/zb3KdIyXu
GmEaQVJJO0UDiWzq6/aDxCuC+vB1rCeRn3p2U7ZdXj5oJTXMEiWvjltDAFSebkpD
RZj5TSgsXf+DKgOHyDBpuOSDqLjt5sJESupR70s22+fUNZG16wLOva6t4fe+oPi4
xu3jRT2To8uTYVH8UZqL+rnCbQ8KoeDHmub+nfNuK8AgsG2A/Ol+YmGrKs9dy502
9uWteI6OwOV+uRpFweHIbtYRJ3cdL8M7im1g7o0506OdciBEvKyFejKy0ruM9XJ4
+pxSCAli3cZFJq+8SY9RPgPb0OI/XFCpznic0SKkg7LCVfjWTPcruZ4RK/zQlKtu
zjJCXMq7m6OjKrMyxGNSaDXmmG8XFOPi4N5ieQre2DSBgMZV37ZnqLse9CJIHdnC
k9jHZw2mUl3s8aAqZBs+BEM5CiF8/d4c6r3bwzeydiTW77AncXJrBlKW3DtxnM2j
/EvXNsdIryrEtC98bYL3h1uNbVsX09V2A17Kq1YTotxZs3iCKh0EfIRKIQW//7FU
mMjdMH05o34qNfu7wjmBBX4NvqzYyZfVzkNeeDLYmZN1wyeRlC9opITMyxD8YlnP
E5TCMRd7zobIPPXBxzaGUubNzkMEOQTGnrlXZ+MW0/I20Po8pZQhS1G4xU4vPzyK
ojECEvsDRxfiSP3sXsNh+0gdkk19mGKQD1PL2osQT28Ce8pAyohujzjpsjhYVIPU
h2mp80Ynbe3TrraDPFTvENMRa3sYrLQnItFk6Cyhdgix3DA/WEY5orAij+X0vNWJ
HMdN4rSZxiHjnUb9ZC2G8EVjymT+HHxwMa+Uf8MK4S8M+Xqda5YqOasm4azGDwn7
lnebJHQ2shZ3G0xE/7DnCYjIGjUOTGW2s9NY9KFuIxqJFKLtxjk2HQw3vl69y5M3
7aRlq/Vn/muEainjPoOSx3pxrjOGfCV0TXDoK1+WG2/4RrMHl3fwXpX7/6lgvjpd
Dcr6aSglTZs/hJuIGCmGzFneFqW27SVKs2DGRflq5tkEv+2UvZUU/QTXmYVUMhbC
bG2Y8+9GfjQ78Krvc9PqSn0GISzr0W8ernJb9WmCrX600bjd8itYwm69w5aC89YS
49XsQrGDyCqIo6o/+GWDPXn/PwOybb7UqWeJRWe0Oa/ICznNu+MOR5Leo+kn21Xu
s0eiLvL47uLZU0fq1qw7EeyXrhAIvUQ8w67j1WAgAJV0L6AFgD1g0aeoj2E8J2Ky
K/S+wdoDuwfI/hVFTSuZVnt/aNpr6TF83QFlqhEnKAe0D4K1oSVcaOXh2DvkXDG/
3hcY/cNVKy3/WIS0Y0B+3siZHVfXspxDS+0nkLOidyKHlSsdGRjj3bH6cr5E9TBa
kTvewwW5aw73M64NHtIwifmiInuFM4jebkad26r6p5jeDDMbKgA8uQAYv04+M7S5
jM8vLDxA+4jXtQuWmrvC8DwHBfjFscbDi/Fv2ZjuDhTgKY6rLrBaHaNYLDjdYvbw
bslDSlKwxmSvjZnMB5z2hZ2XEf1x0MCNAfnbn46+WOYCS0456gDyDSqQjUCVIcw9
+Hf1N+A2Nog9cePzcgA7kf+QN0HzaVOWUi2RYOiSLb7VhGqfSuOoZRgI28R6nyFu
UDHOXd0SHJHo3UiUPVNmvLq+YHmTCKtor/rqb6TSDxca1CZN2A35sbzBUo6zJvph
Io99u0Q+AAZkMJaxa4P/+37h9hmGwUrSO08NTgwvSG8zsqb9W6nOV7YLeb8y8fJ4
tasLna+qUPaMPjzgSWrUhrVzR7W6hF/mCdHsmnw4YFUzRzXj9oHE5Gw4BuJxA93+
J/38sjZWhYS9DppSZgYYsKvVeBkL9SiRWAc+suV1Vuz4cHugqlQ8JehYaoacCodP
vFjX/YWG1HadzpwqI/YAHA8A80i4MOWIQxc5Q75eYQ41+H3TwCyl/AagdKhRHVm7
6HuFlc5kyEYcJ6W327yo1HJvPqMVwBSoUi+U0GvhUGF2kiT9ICtpPTVfMCThdUu3
B3blItne7CQvJANbHXcNF+G6wMnhl4DMnZrXQnHFqMvUU3btsxcEYdCFgSYun5m/
QZ2mYe3ezr2ovQK0+hWeC/0WsIewRYZUxIqD4EVJOWuF+NXWHQW4wqsC5Sa1pWVx
CGDvqiuuuiseGAAg4vlWoXdulR34djTPN/FjIuc8+M+L0m7DMPMckusGyJGTvmQN
Nf+P3Ki6hVrELEgIXXCPNua5Wy5Rs47+BlysBNADNVyfCp8ojkmTnpk+U5W+BJHL
xiHvFDqxuHxgXl2nS6t6vkFdFzjcs3iUQjZJdUIzJVU2EnDUw0+jyPg9AoN3Hvmo
v2xyv3JIo7GZ1u4i6wENFPsreqtSkP2/mJx6f/HCRBb5vnomb7kPQKxVra71RWvf
XKbZInlK8hmDYI+t+Z2mXvdXXkFO7673F2hrXlJHgFqb4H0E0p9e3ZXV9dkhAaVQ
EBKJGQ0fXQbIir2RVP1UCCH1w8r8nbGlcrg0QEdy8WN+F/PidZBwqqfxkOkht+FW
BP3lcsgolXclVr0d0qN1MrZAus5fgVlpE2ZvFJCMDOoZsrw/h/zPYL966ZiN/NEq
aCs3RrN4GcAwsIHc16xxqgJaZzkj3TPR+xgHkG08QGkKR+Hu+80RE5cayo0HenA4
y3pf2ZG/CvMbsH6A7zaTnXJhkm3jjPdFz+OlrIsOTetX/q+iyr2tb04xA0tEzMrJ
A9OxN3vNcOtxcWodNQhEccleCObkyzxJghJVYNdO4dZ+cfLjRuggCYoGLDY+Af5K
CMkjTqc9uBIEKeoRDW2E9ue1Fk7VqUFTuviGuW1giD3U85i0RnSFaAX8Ed0VqpcW
dBdA3shnbMIqNP1bOqR0tfvMn87jT0Z0d4Ic+L98oNYjWY7GIE1G7gb7ATto6HN+
HFF1C+RoK5jHpptBzFZtBEz5PhlPlVm2bStasAwKDMc9zJkhldcplfEKmcGXjGum
FQPsB3gbU5XvxDpsYqwEo+pFuzQipdsHJg5oCusuORVTO8VF1145i91PufY+RhX6
OjbdBQunIxo4/usRsamxef76u9IBoqyw/CRmr8g79Onmgac5mLWjujGjKD38Q8/C
JDbTmiAQuszpDD8KeFp17Nrr68FLCtT3VsItZYm6tDz/Dx+wcMrzDK2wXeKb6vAV
uFMl2iDSFaFltINMfYKVCm6UnfCoTAtFZCkXMBYSFqViKX/92FWOJm0oQTUxFGZ3
+yIArWUCtNKF0MSdajamS2/rS9/fpSlmY6xPRxm3XjQP8u1VdcE6+qd9eJrRHxCC
A+RGyprNoBwjRq6jQEFdWoD5DT4aX3BAd7Zod3+NKcLec0HzHxb6l3m/Oo+h7Ezz
qSP7eHyY5afOtoyUc/DCdT0V16wCB17eZxB6JCVZuPaw/QIjjv8Kt8bkPc+Z5mrZ
sDBTEkgYS3nmxGH5Sc3SjeqNctTlZH13ZubdvYO1DfYQlb3Vct6gSdF4i8XqPDs8
HiYfeYNBoBwn5pAt9PwL+v5GtU00s33LOzppBwOHQTfBFmueYazfgjUDAtrNDTTB
2SghpNDo56czVp9rC5bR7sgCKX6wSUALvYnUeqW67ENSX6zofOiLCmEpSZkoGNnE
zAy3mDianldJ7U2F4gp3xs/8+kIGB02baEHLkvLjrByhc1lGlpafdE/iCRHkeCnW
N7BiULExLWWJ9eqDoNJOEaMqptuPYX1V009FpqPEAK0VFFACegrffqLkWJj6xiYd
1zvooFhRG6CeHD64a+XD0hXP94YmU2E4hEk0Wv/a8gYFABKXEzbUlvq0BLT/3kEN
n5T8K5QAEvBRAm/1usXGl2Q9Jcie+aZaQTzcQKE3IZ/QVeTUvDYt5pMBKWyGPmLU
79X6XGpD3nOm+N3EMV0fCKs9PhdLzGXCgKc1u3nnYKf+jAWnas/FUEgej3y4K7Gu
zNWVFb2hQFEZKjKHlIzv0VJBrhciMh2nrerlcFRcZHrG5m9IdM60iToDQEjbOr/X
LE6tlwAlTYB23XpknYv/pxf03qA0omCIWFVlqRYENKM7gy2hHPdC3TURHogfot6U
ConrDJqSVLbHApdwrCZkoe5+0L7+oJdo1hVFIXqgpVtW0DLH5YWVO0ijXsEnDl4J
MJHG/xh2LNblGqd9wT3rW4Vg6TA3AwExzOKw5SIAH2DR2l7RwrBnbBlWOxxccMps
kcYOPRTUyoxXHBch2Z0Sk5chR9b85TGHQZ0h4Z7/oEPupenWGF/+mCXTV4Q4KyvY
EuwwPi0czP4IwJhzmBvH7pgUWmWPIcWKutLEAQVOMhw/BWs2pp3Ji2L/JKM6PlPE
pUF0+6NHgRqR5N9PuoYpghlBj6oNi/384F3n9pduTV502HNj4YuSYD5AVrKokxT7
Ei7yUxT5qUBTkmw6Bdkpy3rHjnIkBoq34s9acpdgshPdcj7ihdOty3cXP1MwCGFl
q4RPmVgQEoTOJ2ctJyiAaddsi8YCUB/xJzrNCu1dGlJETzOc94OsBjTWIeWml78n
goi113n2SG/M5wtsMIVPO8CNsfeYUY16slqavhsUpkpyHo5uwyuJYm4jRDZeJFkN
51dC38PAtaKkv3IrRQ/3m+VQM+Z5EHY8SFMSo9uY2MHWDnQcKR/q9s+OEMGWQqH/
mCT4Ro5WSBRyD4TFXYG5zuYEIl83gARb7AJX70auLVs3uSumO29LgNgFc01hHXGM
cipkvNmUU+c81gGvmE4eVhj9OZbMynhZFCrzw7uGToF/RmI9wtPSOrSOoTKt2pWe
KcSP3ve60S00F9ewAW0ND6dUS0rSGmXoipOmPHg8rvfSoCYJxOQ1y+d/S3oLlfx8
Gc5XydIQulEkiSjNZ6kQdzSH4AAi9HWdNZ+igHln3pAcuHWDbwR4tUDemnmOkr1H
EDLZkmI4nGRMMtU+KoXKOhe+iEkV1Yyj5DCp1MIfDbRJBgWDAW92i47qgURSmr+d
ixz1Tjcc0b88X2zn9lEvVcSPBdlctaUOUfXLGPk4bdzeWwgSaCgtwvN97WoNz6Ec
dquBCMFycv3SWz6i0r4V7sUiuc7kwJXVYa2EloSODrv7aKhIfpd5MtWZPWXY98r4
hkoAJhE+a9NizlRRpO3y3SaWl9q/FEZ118D7VLB9WO42sgKr7TC0avDVuRzc1MQn
cL9nAqplbLeNdMy/JOvlN1dKAcj+yC3IpLQVdIIBXA+hBdU0ZnaGE4v7x02t8zdm
1SreVsCdZmW27eTMhxTwYVkjpLo8HmEOlMBW+VzD8RQ6rsnLcD96fJwnH+ZZl0AU
kNaLDWL3bNdLdfGIssGQ4xszZeaIr4ckrs3ffvw0WNjBke98N0BUdQD06nQoGK39
BZPR7DoBvk0UMWPPQBCFyF/H9twdFaIKTnA6aHujN4hvLUUUeb+3I6K+Miq8wlLM
4jfgxqv6iitWVngWe1lYwdjyVjwC9rUfHTsijavrG87CNnRkRsMlNEmoC7bwgVj5
+yLC875xD27yiHIux1stN/zKUvo8GxNL0MTb06Iua10tWUdXMpVLHwEuPQdnScqH
42KpqaojsQQyyIdSgQAgcxr+dxYcVhn2oLBsVSDvD8AUjas8t4NsZw+WssTXEGdG
gagr4KotBYIcLsMNhBviW/hlMaOmDkbx25B7JvptbfzJNJ59fevRRzjONh9fyFjh
WsBIL8eF1ebDijnHgPHO08Vqwh2Q2VxO2Rt7j8S1OGxYEq+yTO1aSeRIK6LA7aCM
oh91jsM451ifyrGxdDL+uPvRhEnSVKueKVSy95ukwQ+h1yzhR50dYczN5oRHA8W6
1IDDxvl1ikqTSX2L6Uk81JPcMhcGpaNJUkUb0AMYLpcwuZyXOGS7dKXxvufS8mru
LMlEM0pax3VExipoHiGGsL5S3MrGrte3krEZG/XN1d6toahUEBwa3jD7ETc0j++a
hp0NqAulH/xHkGIHCbT5sD6U+nQwxWN7BPguz8fFpgp0E4+DcZ+VJURQE715V9Jt
unHtmmF/4338homRGBAUy1EWv1CujjC4OlORY5e3P5sDS2kriv+ord8mPC1Ra4Jz
bvhus+OYnKs65plm8lyhk3c2mSEAJN+ZzrSnwsOakduMwLMv5LsXE9Wimt3UuVq5
+vQ0leRUwx/L4RRTuLXOU1AqQliBQk3Ban38vMOIxU49xnlvqNhrKkksB65m+Mb6
d7KUB7y5CS8VnCxS7bbeAkQNkqKEwfSR/NRb708LKwIqalcDiQOFoeK0A4/5dtpu
QyusbCzFP/BiRCmfGndORAJqiznGTu80cLueZupqIaFhg5abg3ncXX3WgV0dEaJY
kWl9z31dViw7Jq9mc9QYMwrNDHyGmcTWxeBqBnBFPRUeJbu2FgIzIj2ukjoxSdCG
w1MoZrULogN3eCrTovAJPh/6Atu8eeAtJwKHWuxAH1k+CrXEvFHPYrXQEsquMokz
YOcoHk3LgyS4bi4GoJ8gl8847kQGhAc9aHQ8cczcXd4ljGy+kKqa4mhr9RnMCkzz
/jtpz96qmk/iJF5eGdd9LmO5iTo6oWZTKHOhWSnM8dmQ0UmiQ4563CbyXv8G3kHQ
WbNIxLV/8IzaNy9f6JlSIVPa9aHo1YWZ3vvKPPONwESBYAGdnSIywPNDlfc8hq+G
+MdmSbwi6WTYZx3TWfxjI8/bxW0LPkmCzFfOWPbP1UTwhx5wIlnv2FFIwHpB5+ab
gs287V2irk/vWLflVUxchd2Wacl94iysQGPnFdyu8Iesr68KKFa18nPSJaTdCpGS
d0KigUPPVTXwUkkYjXbW8GrYVY3tWwLHo7lNuivjXveNMTXp9Jx8R7AhnR6nzrDw
c/O49ByOi7B54K/VXG2VRmCHCB/SWiJ1nowxfha0U4MwYysnudtDFNp4xf8KOAht
CD6gPq4QFsXGy6i7gn5O+zpULX0xiyBMKuV/iFd4AmI+3fKasN/eHSqutQ3ZNw4e
uddzerfy0U02hq4VQn3PuljYdu2EGzlFoeWFCa137bumeZsaCxWA6KuRZTSQJeam
KyLty/JWr/B4Y9xS+JA5n9paT7WeBF71tmo4Tr8W1foK/sF7minibYWioYgtQK/m
N/TOBiDchSrjxvUQP33zqYMAw2Wf087RxcPEm5uSxfg1Ap0MYBrj3MCqcMDKE9fB
zcppqmLmzxQDEqNuDaeTVnaRbxU4Uv+pkmN0AZCF0rWAAtdp1A9z82xgLcIJqCvU
Ir1ogQ+wgJ5xAw2+z9inODzT7rxrWStaQT722xI4bXEW03u7a80Ff6Vrp87r3sqy
HnDE1WqLR5rNo/b/CBn7AQYOk2zWrb7W2PziZpsIUnt+wq7iV6OIySOEa+4+eJUq
//x7In0SudqbYj7Ag3BEOvJHW+TgMzb4CNOYORbpBTHuhcEJ5UB9nd3LCnI89Q7x
LiYIlEDnQQ3plmrlbTNqQPkCDkNVzZYA6yYipM4oHZJT1NdT5IsDL5+YR4i63Fs2
31w9EioGU5d2J1X9f+dwMxMOgHd/rFsLalDwiK/LGlwoFEI/1XChvQxgdjJpE0al
XnHS7JyIOFdGom57sbOBblF1z96JEH1LHVyie5gI9OxwFKlDr8v2AAXzQgyk3mM4
U0TJE8O5YSEmPQYVlGL6K0fzBJXKeaRskKH5NiFkv+ttf/DpfuPzUtIieSdaDXwl
01ZgEWDdwEXk8eG22/H2z8n87E2gWa50JGGzJJV5HRuT1j7y9PoG4BtwnThSyaEM
I5KBb+NMIKyqdI2kNaXEt9Qr9bPNbBjvZe0einJarOk7H3PUkd4HJzZQMz7C4cBu
IWdPtbziHaBRYQdLbEWGpQvtK7WvuI1YWNbqlxARqfmHaSNxEDLL0ZaYEYG50Gol
FMWtzWaajWAKrzD/JrIssHb5A+muLAOBhgtuOq8jHPOFOjMyh6OGbs/rg53l4z1u
ly8DFs5LKePC6NDwHl9D+ReaPK211WuYMj27VtUrPn22faF9d4WG5NKbhRZfm9e4
lckFZ9LL34zWeOQung/Bho1AkN+t2V+tKZpwgnQfKtSoRaDXOrF2N9YCi0OCJBuC
mcOCnYfk684p9lgprbrnYGzIDObhk1jLCGFEcLiS2rthr+kUsUOYEqHoT3pQWNd6
20HuiqbjcaI1olXq8i3kw6v9x/3weyfTd4VhLTZbXSCtPdaqmwKN+r/YeP12+HYo
tNdrof6EJLJs8Ze29vhj74Ijj5IYvwVbtdS4XV2e5ZaiWrZM94+50Z3wmFbGz9Qd
z6kZ7qCF2Yqol6CXBKeV/BWEsw/jmX+GI/VhbMUAcky0WlcohxA6cgg1ev0XFwMt
gvUAcnDmUBbszLEUOJkH+YHUG822In24blH7aWK2ltu8qwFAPstvBnYjpgYZenCI
aZdoaJf1ycBDMnXE4csGONtvWkLpJS5ka0wBNqWc4lbtc/KFO/QjjEZpEvdvZTzQ
Bh8EhqCMsoVqnRbCXtmOtGtK6gzFtR3p380TOSXHiGefJsjs9UTypH1+rA6oyng3
VEBiFT7Tpe77pMVv5HZ+/c70Uq0zKZJ4WdYzjVp/lmTYtdc7VRHT06W1GuonYZ5u
yn84aaz+yba76xbdI2ojkInr8kpqadoFd/H1bzThAILCLQXrRW5BUiu2GCFZ7/Qe
xD1F8AdEXV3IkaLyVjYQ8QV+ybRHPvIuYg4Q6RY6D8khYCZZahOksX1u/1t9DzRj
lNvyicEF6XFyREVzGcm9tsi1KO5BoHR35uQmm8lRSXwFvNUgL3ocFx8wPc3pMboV
wmDppof1DcpJkNHVozHK5iHaU2TTI6DeOICP/PPMk99jWBPT/seyV6XhNtDVxXdk
+SF8aNCVLL8Gp+YnQ+XVC3MAxNJgfXbqBufgkOXj4n8pjN58enupz42Oe/s4sJqS
eEOkeGj+bvcNL2vuZgdpsWtTH1+vhIRqz1y5mam7PcWmqrTqxfQLdR9ccl0hWsFz
3oFdEdSeaXlM+k9vGl7z/1Nh/iS471IPs5+e6KpEdNrudhYuOu0gEncZtBZpa+FC
7pxXmPQK3Ra0na7jStZ1lMUwx9ycWiaojMKmdbdWK5Rh1Q4QlAZx5SFyhyYI0peA
/xvlwitoowgtBGurlLRVgz/Nbfcw9aUMIAaNHnBw8x1A112lsD4PCtLPcBDf2v8z
rZa1Z3AaqyqrncxxG2/C8oZ+inutcwrEtxjIMGAgaanzLpx2sSMK+RPURakyCwHE
3npbGxrIN+CT1vlJnonqaaBUpWtG1QFmd4ClbiakcOJx0Gg3eGlPV3Uen9ysaW90
wBB5qjWGEK1OEKirT0siKHjF/eUEvy/NPe90BgE7vjkfcmK5hhGl+wTKxcWj9D1K
/uC3Y9UbAtLOg0qcBjucWloInIAT33uyRqUxGWCPfs0EEwaSbNs30ACzqy5clUX4
weHQVvcZWqRmzc+zDtTqToHmV84yMdRF9iBmPppHjgT+DxQ/fPJeO2rk3B34zzvR
i68PyzmV8silvWvJgsggHD5oicmtXzmjBNJBXq1JRpUCiq9u7BNpE+jTtWH38irm
V5WY9/AQ9tsg5ROYEKatG8k/IByEnaYno+Jocep+C8uUbSKquGpND72PwrzxEQHT
IQE+Mgsk3a2Ksi1qEHHo2WOFdM0a14F4mwPxb1n0ulDFCZ6Tr0uUTSFM8a0qouH7
2phByTiV7ljhvV6qw2JkqbL1BkW2Oy8Hzmtbf6U7XqDIKdSSuhHhwKrAZyuWmrrb
w56sXNTTsdCKiX7PZrEKBs8aZ9PWHiGTrilEiYlcGnMz3h224zXLjmgBgib4DTof
bl19jUuZ6cJOqDr1zLRtfMMW2OFo5xsXhYmQATbAzhpRqhGBCO32wOIz2+hW8bAV
XcvYPagfYdRvI9MyuYzeZvfHufnqbj8Km4yjlKW7V6k3uV+n3o8OpGqAd8GTCayE
cA1agG5Hn5L7SbGR1wopfL/0fonHGzXhT1aOp+cfkreW5dMCws0GK1j9sWl6FXgg
zn7y6yhv7XEEUR+basPt0zhEJ72PEo5SsxQZr4F/D7+rNRkGxSogYyt8LgtKY7hJ
Na3+gdoodh2zUPOJRyIKlDzPNmiUY68LDuMbFIeYiBi5uszwYMKnhpmEdpAlVIM4
julmhwItVGf6Hb04X8OVVwiTPhEiB3SUztDb983X4UbTCjLnokLY6X4F3wZTu19p
6OOQ6tEiUt30qbHokNoRB8K4HL2u6u6wV6govfvM5rg6PurkR62/pgmhPOslehyP
jyg5ws9VL9ICDvlxFaAtvxj93/0s49VfRAKq6rE9jRs+fR0NZo8Almb/DTENpn9D
XQEf8kaain2h0vG2ZjaIXeRSEtbXMRaL1GFdsPWfmNNcJM53FV1bfKa5z2VwTjz+
F0x/EU1Po7yIeHRMsfnRc6ZL8a5Wnn8u3t7vq4w/YZUFeAhTZTY4Wpo2E3AG/avb
82aS7EALPmMEbbn+K+JrZPCBp8p56SuVAR4EXlJpLOsSvHlgA93QBPBbAQwL+3+b
cspMJFRs5/TdAk19hy5nAVIADw1QwxWIy0L6dz3X6dS6RbcsunuuCY21BE7GhR6Y
XcEeeOl5dt1DKc7tDxxPvErHNQ99WT9ppouwVoFTai3DVm7eyB25HCqc7BYX7hRX
YyEc6miLO17yhnh3IRR3BtRm297sdID3sYNFAm/0rpuZdw91vGIBhBVGKvsHY8se
+XRJqEktAHMe7oLhfugKMS+1ZlKQOqTDJhiNNv+heSZ6lBCzqKeeAqKef9jzwz/W
8K7ra8ZbkjWHe8BIB31dV/jxeoAwbNtKVMO+zY5jck9axhiY3Fxh77FsltEvrGNH
a/+J3RHjpS4PGOZ9lKLdbE3g1fiHtlcyMNFmoImWgda+QXYwhAItB1sZOh9k9Mjo
OtO4h1YeFSvtyvj0eAv4czuzsHsBTbzZ6yVkdt0rWB1KXXT0acBNitkZcbZHqlbf
FMuUU9UFSBz/N9y9RFe4uZfBXzsHyWyFSAVgXX7/9tFi9P0leggZHLpEkQ5D/d6z
QbYb26bD9bmgkvFKhK3hijIvhxL4dmWUE23KTIV4sheypO+5/aMOWrWAhYWoAtLa
C9G6A7CqRFWmtkosIKrxoaDVpD4SzcNUNU5LTC9ycyuA+bn7DKXidIEocN7b4FXn
bQf8qeuSSaXg99/vQf13CssmWM0oEfMskSf/KwUKOP+4Dfsp6rf7pXOqfCJu83A5
aYI6B+Mf42jwWKq7EGit7l2EdWgcidBy2p4t5614XJ/Xg1Gaf3QC5SKWoUcxgRkj
quTZj0nC5re8OEt3DMHrXQTIOI1E+LopLu+UrW3b0kbKNkc9U2X8MBF94WNEA9AN
+bSYRcthVgaHI9du6GYCskOfUMnSuE1QWso/4gG5vQPtNAZI8rAKAtIWrtqv8Cuw
Otk2IpgwkiIF1ctBvgilqN9vS8n5wMKErS+1bU1ZR/9kl/jcmS2ElsEQPqVvs1YE
0CUCBmnNhZjSU5UoMrGeE1B+20lhkdtKBkkalPcZdrg+C+XUfAg0x7zYfVFAQYZA
QaC0qReya9yt0LmYhvX2oPu7LYg0aGVwDjyq85ruTHZbuiVRlc5+MLFD7yYWe0Xm
4JEz4WNGwJWFjOX6BoQ+dlB/Tzz3ZPnrbIGvEz3oqnkG1zgkVvUHSTGzEg29uAGL
amEiLudXCOpI0wkZVn7djnxzv8Kt3BxxHvyqofIVHK1JI8+crLduRyjhLSlbvLsQ
QY87J40pnH7tTaiZEvBr4h+GwsDYhZ3nCxe52YHnzWrxcPGZI8j6tNuDJyjyKvIR
pfXWhIMPGXvDR2fcN79c5CyYmDbEwFrQ4oEF4QNmcqivLxhNiQh/VIerxWdpxeYg
UMQfSPUM+vHfUMIBVbwmWhWdSGKVRSBVCH2lM1GJZkRWEWJJdqYdZNpboM9C90sy
f+xtoxnb2FJq9OIaEfXLwyO2D8RQubsLXCDrQDfbeahkFePamA2AtfW7c44GbGwN
BAdUn5KBkaFX1NRvDG3cHt3kZ3DvqcqL6/x+0aPh5+m7sLck7ic0og9dhFtPBCHP
dzh7R3CUzHdP0FBz1+SvtufxtVdzZOfeiCA6CESpXNcPbR38khRsOfcqmINem/w2
Xxc0/aBW59GlBawPiN3BLjwrTzAFuPoeFYw9NHGoYbNa6EdqWo04SG37tysJm4Ab
0fI1li5gesQbhNVggufuW8E5hNed8mldW24dxNGXuSyN/0qpVq3MHXlqR1C3zBwo
LSqVZgMqQ9ggzunXgtqcIEd8Bg2apMkrqv1a7+UcGXvvYgqxo+XK3efOjeGl/qT6
/Wg6WTaOj5gdSZBBUukkhDsMMsYHtr+b+JpFFnNMAKN0ACC1boAimQKlffoinu8x
RJTJlFS22wnhdJQTIUbDpa6/QEX+l3/IBQDvWWBHZ22AhAqfOXPja657AnqpELa/
aE0JotnBWhGuTFp3+nwLxi65vTjcbhFVbyeYkic6eogkSC6YEINj/DBpeewqweIE
rPRGfXOMiShuzC5gZ9q2E8wD/y5sxldU8vjsdYRVnzBqyeg7kXmanVqih4xry5o6
RvId/O4Upgy5RboRJd+F1quyMS7Me7cbGwtrnCgNzyV9fMYbrXkuDT6GDpy1UozW
Oiz+YTgBsVwy+ilDaWLA0OXp2qRXLFaqMjgL7A/m3PoMzput0QfYPUk0oXsYDFmb
T1rqVbPBr1iWoMHmFHsAy7wEzrjjIExuxa+grbTgIIGwBq6qrfxQxOfdg7yZEYGm
2BCcA5GPT23Fnapgyfkz5+xJc60++vxxGXu1Sz7FDiKWQAzqs4tIvyCGCw01cUHc
30BQzsf528PL04d0Ryo4MieLZVLq/9Ffl9F6q/qD/R+vQ6BMXAZNzAiBDHtDwEjn
yWHyA/XxLxVSIF9LXOPDf+xz/dxjbX9MIteCqppzYWGEOAUINvQjh47ITuBU3nI9
werLA3RGeNWNEdKmxcaaqYxIj1rIHxzgAUJvZJnIraBM15VE/WAZWQeZ5yKeeZZh
CwmFKjG/foCHQ0+wGwvJDn4Fm0jEkeCHkX52MBJnf5L4j3g/Uf6F8YZ9sMnVqYFr
GG8QktCBrY4nwyhDLP67QZUeUiG1sWfzxjyF3HUukqwo5iDY8NumT8IexCc5FLMm
Z5csGLc+V0VlvJ9tCJBgUyE6DjkqcEYyp7HU6ms9/wvezkfi2ZY+Vzi/IJi7Sof4
gmobY4R4GV1nNbxWXrcxwJbPhm1s7QNc/RKJfVuchckZLz6zyZ4rNucp4MqwuUua
L0y899VYE4AsAir7df7znujlHxDR+jcJkVTHlUeUCnBihZUn8gdkRyfhmZn/E2jX
+Ef9h7zNEYfTcJa+FtNV/+R2B0CVsvOtAvo0N2wGfi+hLdqk6F4b6cVIfGE+mE1s
aFWJ0FszlcqP/O0YOR87p96SCtZ+7KNVm5ttZBrQpIVjyWJ5xCzO+jbPMQs0gMo+
SBJn4Guwxu/MnfrbT03F3BcF8tNielKxnYYzG6yCD47/2+1zjX81fzxFCKC3pEx2
WiB5WpsFNtp/LSauslUG6w8NbC3UyiyMkhnnqUQuEslA1pkxjSUWCm+DZXqmmkK5
bXrlTCAEzxEHWAwieHq9P/SSUpzYbhYwOWYWmyu6sTgiufP+F5GFAfjfvkM0/Hvn
MDdkO2//3VN2ouGMBJg0Ui7zGqMCxn/oDH60heZLYeQ+hSBgeQegysOqIi2uNnBS
nlb88xjNLIreOn0+veC/ojgUDl4IzEpKS8nf5yUfOCaYxyjYN0YFCSluRfJlFeHu
/8maOuQhjt86kAQsIYaHdEXiT5w60AvoElFyuh2Dwrq/uSXGtHLB7tjraGoMdPTO
wWgcRMhd/ukA1SCQGgQ9/AOQ7p4I3QnpOWmL0dEpDqbJKIE8YjN6kD7+InJ7zaAf
OcCb0JU0BAUOEZEEfxpGn75/O7+gpQmJ8jO6qmji1Er1aaaZG63hh2FmqHiN2Yd2
vb3STksbfCuXtdCxBVIe1rcQdEig9TyXK37KWoqJCg0OdDomwENYWmib8cPBoegv
ow7M0IsgW1J832+9ykuQOTz1xzUZdH29hHq94I7KZOsgMcdBioWjqtn34oGEjJpc
jnYXa77YQPdapfhFEswag11Pe6/38eg/Xt+QoUf9MFY+eScI/qeR81j6wZo/P3Yy
Ny0tSFTh/jVbOxSmlSgarAKTRPdxoQVorABpiwJibhFcOif8WlHr1DFDDI+rlJOr
q4q94Pl6hA/YOktmP5xe6DPKipg/Pu4DPphaVcoNKKwIrYfOYgLLV0J5Zkoqp/6f
ARmpCOXtjUY4EFoWSY5s8GxxlKUwqKuiblYSgACDsPVhXOPNc+GZarWMoumz8toO
qZ5V9du1n/V0paLoSf3JPTcfkIC/ESTxicPO8bmPSovR3z8yMFpDXYT8sdLsrfQx
uVdf7XcsyOjcyhxHx/v4f5XUq7Uoq4yhpHlvhVfCmPizp6y6djo8LY9xhdhT9seJ
Ew5aDqjwGUR+IxcAijCDQqOCIBxrVdJeAg2jq1fny8kI+2wKF8ZJsfclbAp4qfKd
ePkN6dbgb/T92lafPTIfYm2+T5nSy9MnLgq5zwgpzDBgXtpaZZfKR6r3yAxm3LfX
DR3BW8UCtro7jkGaScUD+GSYaB5FFAIFbtOF7OP1TVA1cpm5O+c+AM9uCQ9EAD5o
Wd4+5xXpcXrb0H3iqQCwZp8jvO9RkC0K4yribWrpDjvIbjmc2w7VdHzoRG7s56YC
w+xNiUa2sTkpiHoDPp9FkKKdqxInKu7yOeQWYgLWivg1Ai2ADqOeexuyHK4YUv9e
KER2/oVUcGTehYAxBoqadc58veK3zrIhYQ70b+MbVCZY3UeoyM0CkeLSQnrbn+gY
Wye1XvEHISpMR08ztZQnO58byg6qrO+C0vlC7NKf//dA0xs+ZB+k6iqGlWEnQSUf
lSaZdSWjLUjFSH1VVAlR4IA3wDhR+22UK0xwWFjApE2i+Jkf1y/n2IDhJNJINOgt
6FDYs6X5EHvhYP8Iuz4RDxx4B9b/jDP+9zFzwKKYSCMV2SpRPIjpIroYVdZFzHfn
4ZgnOGniTvKMdGDko+U/Oqe+mQQCbhLbncdsgUvlQedOzyNp4vyLxd+7gAQ6H/zP
prOohQQI3SIbuB0Nv8Wj5/HhaUbnCire3su7l9c3X4A+3bq4Ct+geLhB+2ahCJQf
Rm+waxNyQveerL+tOm/5wYshGro9RnRcCp3R4pyLiSpC2xPpCQUFG9BGXMjVkq1x
vMXh8tpAU2eH75ZyZZgsrC6oAJEVlUi4AfiENKk5T4qZegTGoNOpbgO3gCTiHIbU
gQO/9wMsCcrW5Tcfo2Gm8bj/KQ+QufnXIlMDQPuWENIFs3gtyCYRhkLaTNGV2Lik
8XxiM5tkU3RS3r7iYL8asTjUqyOTe2GLlgjXsPZXVSZd5c0D2YX1IiSXHL7iWuUZ
cw1sf7w7yi5IEmUpj8F+WBOeAV5wclGi1do7IUzJxysdkoHpx15C49+Jt73ApVQw
DBOhSFhFnbIV12UuJKKVSou+v9tsh60m4GvqgazOFQxJA1oo4c2sD2FCSIBmedNg
NNuBNt+97zPyzC/p01vqp0ldWw19o5/9uYeRAAYUScik9t8rAr2iBgFHgAf5CRPD
RDF8fu2X5cawAd0MH4RURNhoiCPdG0lQOO0jhDhSZNvTW3RiU50zr56/c/A64oZg
gCMGUD/lgyduUikXbcYFhhgS8M3ZuHavZxnQTtsjkQZFrX300gX9gW/2Uj5qtGIJ
oYni/DG28nLXIgOe6H1Qf4c3jC9/2CBJEhRXZEqcTxvudv3Hksz+l/30wD7q29D5
lrgqvqnyNckStjAwUhGfu+LArQg2zJ0mgn5jVh/Su/o032lYx3pcCO1/pWjbS5I8
mn1pNha6h94S1IAleJt3bYgQFH21/DEyD6bndcQz/UEJhI0Euyv0/3QWTfPuR9Nx
zV57xH+SpR+l7iAMpcXxLEJQfJuWrMfeSoJMXRN/FpW4/89TZwxwIm6gb7+8c8Wp
fwD7Yq0gJaq9QLOG24DJlD7TxrtophPiak1YUQwaDGUQKHpCfUa73Q5g0Z4HSFnf
tVlh6VqXhpOtJrJ077sglY/B6TO/qfCM6Xr0GKLT/pUDuercCu+KhJVumNxEqlsC
BRRnD8HGDchF/5Q28cMzrHWEyFaXvZi0Dv7VlQFCZ17hGHK2ag709KBFg6051rU9
Ua1rMoCWayWBuZ3r1y9Px500IU5tKZsOM6H94O8cIPInxu03KDYA83ymSgMMXqGD
1xB2/a0DQ/UNPU2Rk156d5kMPtWUkzD0XR66t3x97qebg8ldkGmNwZnynrtTGN5h
hww+8Q0fOVDYEv8oNvcFtEj5vU0miz0ZLsS2CmnqAFyvJ85MRY+xCkoNtcFhryaj
W3yZJPEmElQs4QKm+juWS2H35YzAc6SBMSOJ3W3+nJYBzpLe/Sp4m177TqzYD1QR
/5Qs3SGY0nM46ijPTp+TxBKCciOmUUbe7+S1zPLKTOh5PlL4DRqrI+xH0vP/gGJu
5D54rkfb8r/fFC3mQs8RkH2PDfTOfVBNvmRqbYKtRkyhQEInjS/HLJXAZqE/L0XO
LYJz2teSuE0qUmyKQF1yiXiaIkUfP7BnwDxSaJ228159TTIlvzg43ecjQalf2ovK
xBqPY88xrStX6N/kUgvIngh7FBVRWGpRhnGCRszU7GJJm0CYdaIRtp4f9GxelocF
Q++xUb1EZV+KowWBz5OA6LxBvk1pgW5VknfzHl812BU1VBmi8BRnnbHdkmbBylTa
oukcE54CMPvQHYhWSGUds3fLDjHSv3m1Wd13FMgMu6jnNgfb4DNiM4ZPpXSTBbA7
PUW5U56SB6YHHamgyDRs1Um5s4KG5JBjnZk33/5tYjsLhj3M07k4GbjRFrXzq7H1
VoP4iH5SJ/DknhIldR//ZjLE1FXl4Piktk8RmzKMIJWxLYspJ36IFA1Q8jgXpW3p
r3VJFFIs+PlyYz7KFybtnLFMVwba+95Uw3gb2B1RMzjeqUAcpKvskUSXoSP7Fh8Q
ayepBZcJmSjgCsnBwVrhmkGGK6+Qac78vyRX1zmL+svZv42RHxK2imc4wcEihVa7
iVaE6IYC4apXiUeWwBz/tsnXSoNLtHEjbacVsiwuTIHMSo6H/Kls/6v5w+huBcBI
lWVbvZArHdWmL14l+Qx3tSbeWgzpTLo5i5NvBDPAEFq3nGbjLgd2SvjZYtcjiVjz
mOu8umdmg9xGBvIEwUOGbu6yXUJOlqk8TlKd9Tq4ss9cW6mFQzmLyzOBgu3IMgGJ
5UjF3gSIGai4iA8SgnYZdBmk2Qq9aQgM5hkP7sRFDx50Mzo9OfNJkHg6IcpsFfPn
R693BM4qFolZ6w6hEkYLzqqBQuTqQM9fIJK/faE8IRDAiCIlVsAlLDOtm0fuobVS
w9PLQizXLVrwb3RMoAUdkI4n+4KmKCPAdqH1AE3iUqln5mGs+sV1UTsaGx7ORCA8
pBGQu8D1tZQxJPcGHa5XqrGVKxZy7ZWa1KMazbGgdv80WgL9Q9DVAwjx9wW8EywX
bLI9vJkzdYo5mi+S467/Emwci8+8ZE4/X0uA2toP3GYnEpqR0XWLICAfHz0CQyDR
KvuGsmcofxAz6h+AdLOctobJiPSkW3sT/iIuYelZ2rqjMI68zj8fOSjSpHmh7LV2
GQvO7meotpXj9/h5tjQ4l3/wJTj+fJAS9lo7nm+H4zB8QCE2XAwIntNwQqghH852
gUvSP5Ztix3rqy3Mwu5NbxnzAlN/qvMa/WtcTlGJtRMYvIwkM5XZJapBckDl3dcO
c7aB+L666xNBhsRUzL/flMtv1HRKLJWsV+o5DP5YZmKYxRNgLkR6SE3kl8ub9t1W
nzuuY0VDmwm6EcdyJDt7KipL2vh7wQ5U4LDqLq2sNWMq9TPaslETFPoDdjv0kwkO
a8DS3IrvtGP7uw+cEcTH59xDATMnHeuaq5eurHMmSwO5Tc+cKyc8yvYiQwkEmFyX
51A26CLrXRIuC3bLGeYwzOn9yYNdDwprnYekWEgmB92aju6CcPbnJ0GyDgwqEWT6
jGBvpSuD5kjvgk7dHA/W9opjYQcPxJurjrOycE7wbONZvkYWwKxNC6p12Eo0Xd9o
/2GHwIKECZgBqJe02WzxykvW6S/UbPTa+9mhluEgo3lmFfIwMw7ZyVGbbrk0sVlN
59I4UrUTY5IQdfdZ6GyWut4HNpBdgz9Y1x0ZI0g3avTxcb7tEXDtsGWrdtO+7e7Q
P8QVF+N4GWyBNhau8si0ArajbnKtw9QB1IkR/8Dg+HASfyU1OlD6OVFMbKn500gv
hf1FGRMaaE/oYJBtB/m8r/E0mbJwmxS2WTutSW0G2Y7HzJg3tN7e5XasWh+PGAGx
hkbIFDGnZovfAS213LlHp0rq2aOb29kOVjCZDZKqWH5GCgxmo/6PwzOIYC92WJHp
3t/7AwK5nYYZysV/Jrh9anrDJRo1e5CnVFgbITKiQm7SuJPPud/L9Lfr7cCpxmjx
GlqQqVyWFJgNqRG8f3/MktBPttUMdZU9aHDNis3uBNTDhJ9MpWOeueQHYiPO2zuo
/VuYYIvjT5hHrVWDA0NUmBGwotx4G0hfvRP375zPGz/b3Y5yeaVb3G/7NXCBvjGY
yYFcYbjVpr7OIkmZwdjzFBLx7aflUobK/zz/eBbHddd+0Myguh1c/e9aYPdl3G8e
HmXHZrxqiYg8ryZh1wP2KHpkKTTarlkg8eQIEHgP4Hqd2BRDF4vw4fnFwLzkL3FF
7X5rHy26VG1Z6sA/70SoiN6b1TouN8S5e3o2W5245uuFY0PudRiIUWJOGQ6MHbLI
VZ/UISpSdChsUgCxmLeliO+M+Q1HaT0ew8u/imHerrirIa8+rAcMnpYkJ0jxRe9Q
nyMJZfMlXmKbwS69Ep8zxTJcMzwbjzf45NMMdFcIp2bIzQPdL9MM+DSwFIxiATZn
HglMVrvGUuClocaQ8rF+iMXsSf0YR3V2ms2d7HN/FiI8nTQvprLT4CTJwNuim7qS
yWF4n1l0/xCrKiqdtu7KHnW26elsepvf6jdg7BTpPCR2yD8su8GW+41eXoyrjINj
UzPPZIb1DpSY4UUTpE7Gab8DXJ6xIGVgBN2blHxyUTimNOrM4Cp8G8Cm42X6+HNi
i3xtzCBCa+NAVPXwaxOKnvjNpvF9rIZOUqqI2GnLCeDFAD3XiTk7reuTB6qgpHL/
Xi18V/5SSMarRhX/0RSvVSRFpjOYNtf12FAfm43UgTo6x3QbNHEkZmuF/oTgz/88
ZXDStkhAxZNVYzb+xjtvE4UomM4x82Cx6Ot1XsmvODj917Mf/+9IFVaxy1I9Isvm
xftIKfSIzXsGf9qG8vL0ObvpDqeKVBfso7lm4Q/4RwyVmKLYToHG0gGOZ1Dey+X5
oy/WItVPz9cDf8qoucaojEmc9HpmDj0Yt3UIHPKN9RAo/x/hSShLIXNbE9LaOLXr
3ndW0fG8b1kjc0hyxHxWJXHeqpsQFzwEWxjldhp2qXDlWbD/XwxIGpU8bhAempoz
ltQHIL9KFZGMVZgQOLfoy0AveAMfxEKsaOWM3smM2dVEHd+HtjiKaFNqtR2w+bD8
qYRgAkFkZyrx1gC1+MkSkM0Lx/GHg1Ytp+o0fwgvQ1u28KxTQZ+MW7zNO0V0H14J
wQQOSXoqJQfesnFNL2f/tSg2O8u6Fj0mTXJTMHX74nwozEbBm6uuxlchwX2K+1bp
UxKYEFSz8qB9aGD33Cg2EiELUJ9SBkV4NNyYtJlkXFnNInl1xNhIDiN/nv53OGdz
uPVVHei5NFpHwDOKCwCxg4/5MvqZeREafo6A6f0DeyyTCRJUfPuYJzPYnrLMjgnN
UwyH0G4Xtug8XFQP176jtM9Be/0r8bVksBJ6D1kYtSOKJbXXKelIHIC1J2/qk11i
TWdkZ8S//cI+sq4Z9yNDF3yzdix8PvXC7zrrM1xcGlzYUS8/rKwT1MTVKejB0DSP
TXYZaRq/thie/Rm9E3hobzdgRlGrKOoFuSBQqUrmN3Xw+QizW9M557nLkmJ8GtR4
M5D2r7Z/385FdlE/A7fdRtER96SRxYjKO7zeq7F0gL4A2Gc9oCPnxlBw0JfBt/TE
tWSWnK1YpKOgG190GgKXkg4t8W54JNVrquAw5mAmfBeP7n4Kx6NuVxwrw5/aLPeL
uaKSjQFPgxDGG3mp8Gb47AlpC+UfQwdKmPJYossDGPQbwRWggZxHxrgLB18x6gsV
UuU3iqTSV+HC7hqWGiUBZDM5Yl082vMEWI1mGNtwdQYjSNL89HaGOTXbhn1tZ3/l
7CP02xFGnF9upwicsNPEKsjGYbYyKPGjDv0WyI99fW4D6BT87RIWw9QkDZTU5f9l
TUTUPOZugramqV1X9K9yfeg6vp9PGdDoW2iBKLZCxcbM3pZNOM/H0ANDvkokdllP
pDxxvXkBMyGc8RLs9oB0xFIQvh7iVc+5vYdGyL6rSvXls4WoUIcu7LRq3qUycWtr
y5290WypN9YiKQlNI8iuOCUqFq2jEKn0C8pmwe7g6nYxSt7RcbIITcXag0Zjnnfn
v7xSJ5TZ0ASTcxDQRYN18LPhO9Eu3lMAq+yhDC8/+JISWvoNvvRZuh8PgH9Sx2vn
pp+w9zP/81AGwbluoys40SLk3kURQlVkIyCsZEGwWQ/zgFWl5FRSoIzRv5n/FhVT
sXGuh4IGhQVBaGXMXoteQBS2La8vPeopGxgBZDQ8q9eJfTk+MQI+wfg9dxgjkblW
3eAXVHUpPSUFTUi6o3kyZbEq7+PJcOTRjSNS59h3LnseOS8MICx3PIylmmq7MMmf
i9hBUIMu8nyZWZxwstLUVc9oqkYSqF7o2kc7eLv9d2c6QPCmP7JbY/7SKX3c1hJe
qjy5b3PwPdrv5gJBECBlAlVl8cdxC2do7Bwt5MavgWNzohbgj8GMmXvQxcjnTgvW
mbvqWJKr+KZRRw5/xrIK+VWB0eGIWrbk1KINMBCCoGUSXNhF5Wusmh1SU/fb5Fpf
vVUUn1yCWI/jzmw6/107Nvx9Mo3ubrDik/PRMoumrc//OCso9fN+3YJZY9NxGBiT
g3BATLZ8T2aTHpbJ2PHuqtspFQE7PdvBvV2dH0pZF0NzXQsFzhhBSGndwaDKfxxN
ZaZoVKSBRdD1kHO1WXM4pQuBULlI9Xq9X5GyPCVtQSc/ZT8bDipurzOT7OWomtQQ
JHd9tbi4E6m/eyXTPpixwZyZwPatpM7fZohjCodPweJlcKlqgTLm0zzha2fvKc5r
FBt/pdGmf2mz4J30nRXtTt4TObtiZHSfC3XLZozxhUliayTUQLbnu9BqgTazVtG9
rzunfUmX61kePe80K1zxGlE2hQyPfvUU7dbQvgas4n8eTadTn2Q5l4XHydwy6LBS
eva801ATGEvhgdt8eHrD65GOFNBFJVjU8bUaO53CH3p4QltFuHWgDB38yY67WnPD
Iif81ZLHmXUKF/sE+2+lpRvBZYg90AvY6xQbyGLSI/LKkpw+Ig7Me9GtCxAPIX9N
nF+8Gv0F2FSv6pSkIPNEGyZ+s4VKGLjS/Dgar/HigcOf+UlwDJv8AsLfqqLiuV08
Lc9/HQtaXX3k9cZ+jKmWx/dISjOLaagB306NFm+LB6K14kILSKAZH/50mL/Zp2Qs
TgnEIVgdHxnWyglG7iCg5PhC/b8L1qzDq7wdzLnOxJr8kWZ3+huZ9PlO1pYGRgR0
UX/w1l5TT02RUwoqbRRtmXNjdW25bl5AkcEAmM4LPG7kYYLtR4t09jb4kWwp343a
qOyv7TDA8g3NQRXLG1K4hnHx+UFsbWebc0aDsPvzCkLoNz5rol9Lmrk8eAUWc6jd
2xiST18hkeRj9Ky5JHc/OhqF+NFXRtHhDaMfijqJzptgmHSEaX3iMt5QVA89DAD5
e9NNoTxXygAsbS3jyjgHQK7xpGJHXWkc31F0u0/JBmwfA8VqFAJDSBGApjLHtY+i
6DxIvMRVQPt3120VTf1sL+Zj96B1OMzJCxg6h5n8ywagHWINwkDNL4SLVryDDYCw
P3VXmv/+d4lPYqnibwhA9W/ERphJhNnj6KQ9Yu98alLfr/tbvEUUdR//1c0p6R0f
sMrHX1Mtu6VzV75Ne5haBbcWt9l4oEOBBpaS6M3mNR5q/AvlmNTOj/rgYNTjmlbG
Y0DQwwOB6HAmtRLLimro2fJxCneSEqcsxiZkTa4RnktnAbWBWa5tustn212sOQVX
WVdfvWzCiVbVnmO/5CXjUaVuTnA+hIke/fsDs/rHG8+QeFe06f6MmpdVCa9O7o2s
uZ0N/9cLV9Vsv4LGJa54V2KWxjIVCNmQ37fXFhX95cKYtbPUR6ygaUAJ5Zw60054
rDA7i7t9Tb6J6hWWVUQ1OQaMuPen8QFGN96I/pwrXDDWfQWSEagcHuKVYb2pDr0L
hZkyrSJAZMYL1KQkHS1SGnMvXw1Lch1IBUcoqDtmzKtyi960bAATXpiappIXn9wj
MuwdYIABcotcSOQWGCPtUJ4A9xnrLBah9qUvm5thfoNr6luGMx1KWLUfaBBotMpf
ozKWlpW3XBiFLQM94W8RBuX+DixUN1BzOj5L1emA6STxDODG/QfO9ZBm/ga1o3Ty
jbugXKrQWDkbUeR/AiBNi2GOS+XutEammfHM1njKSECOmZRYZndiju8sl0bW4Gda
MWN3DqMpgMAX+JfVeruzMDdC1kn4UR3+tiTEnyUl7nTwIyJ7twjzcAJdS8AiHs7n
ok7ELPJYc8pDlYXpZKeHx/u1f+0MDYiy1He88oZMQK7jX9jpXd3hYMMNLDg5SbHU
FPABt41iaYFAizGAciFai3GctK/TGcDtQEkzyHnz/jtEA4SLp121jab1xIKk9loU
aA49OZrudAu7zj2YBDLSnHTpgn2LcvUNVNDO0FwLV67Tth9Kvdnui1J6qDwngR58
oOzQhHVsiGXzsqi6wVqUtUOrzdC1bBoEJe0MgUrrc0nGVF4tfIzcbf72mpCOKMll
AyudBshuICHU/w3Jb/wNiVZDnzbnmgyc3utKKpljupsMYSDLRF7km0Z8fWHBDo4e
LyySkIiiOHrReZObE/4JSDhatd5PFXPLIhmSWGkxfDMQcc9ULamfI3lSxz0QHgvf
x+9/+JNHP3J9eSjERM0gtSxUDLjf2vbMgMSXnwgKSSWqxTdeJawDEBwGI7dwgNHP
FEMSHMNvW9qTuhZiJGdGPCgTYF3WVFu4hzNZydvMHa69pGThk2eA4c7qeunc4pLT
uS2AqN1j+VDTJtQ0ejn8NCFrcC55wPBwjy4cyovDfzMoJxVp9hJYmAtOSnb/9c2q
sh/1RefCSJixOWn7zyWGg8jtHCt48TKNw3fcTnMjhPfsxIWnxa9tq3ZR2xcBvM6X
Yqze72VdRoOfBbZdUF2mcWmvmiNsEdUSuYRWFITWe9We4oISC8WrVsEsejC84cnH
13muc5lqhURD+5WiEfrShWqQfjwzoQRVRL5n4iNhAkOp5fuGZLtsGIFBZUpTj7XL
bqtA6l8DX8zBL+twwE33ddXnx+BdtduiGJN8ray5tfaFur1KtGSLzy2m9mxUY4qR
5Dme8CGSOD3SgdVB8BiibItzHqF8Ga1AITeM8Bs7MAOZlEDE69Bgayzpq1Yivchx
C17RilA9L3/JdsWD5+mTcX7hq2oH8L3aGaHVWGq8z7VH1+0EWbr+X77LJAbtmY0x
8lLTIQE1p1fc9J+xtYRba4BKFSzoVVU2LAaCzhFbaiaKDi6Hxyb62g+WLqNYf77t
5VBE4Pni5ZadMu2Im27mdmqouGhYu7g+HqIGjUuRTr36toUdPa2pPqFWesgibCaY
US44zjwjxmG+awLreymd1YMyKE1ww7D02BTHv6Y+0kaTllwUFWOuuN3ZiUY2wPQ+
av3cJ01EKSWcBw2e0SSit6egmaPN37HIJa1qXTrSx5Y1bob6U52/K4yYDxNuRguR
PM60q+m/CiZxOXc7zQ/B4tnufhG9/KDaCblVVVejjbF6z+jJrep1+yF2ciYZS/pM
z0VkrX6Mg6OuSTQmWJxSfoEQ0f1DbwZN/V194ddG/TSADvB/AaWZImwiIxIBVu3i
2hzz+grEr/dsAJFwckDZcJf2Fats/USlXja5gxWIkN11smqPcL/m4G+o+2yVqW6d
06NY/1XKC2J5osqQTAPD1j5pbvLsVsX5PyEKB+Xf8bdqxrw7i6oL4cHLxtn4QISo
HsV6pZvgFnGviTv4X/s+eUJHTZURi/e2D+JWOTaR2DtiZoMCQtkubLsGk9MsBpj6
Lu9qDf59ZjwBgB6UGp0WuM6F7hLtlhrz2IW/z4cxXiCwd3Ymipoump3qb6maikGj
rWuDdIBIeDJt4GKK+/SaTh6OUcvVZnNlWLzNMXv3RormQtRyUUIx+namgunQCG6l
u9ksUiqUhfu3tqvtZ4xucOUxsBFjaH01ECM9xkIElrG5Ys6hjTHEty5BvAr5NELO
RrB+yC26PDeXlJQgK9Vlm0v/CfRKf6iWhVEDZUkHX7Dx8NMV2LvO5cFsToBa3uH0
qaAdKHQ6CKXHsWyUEl2ZFynqIGvAWiXiIaum6JaqWFOdsyM29WG/3hWTV6NRP5Zy
rBQ1zcwgLvr+bpA7SdReoFQbuPgw12S8HxT+YxH9SteNLtjrZMEVgZ9L8rBZwGOk
TmNuyzM/HJCEmUZ0ORiaw2bv0aUl8VOb/jnv4umLCKsar3BiVzpM8glNw0BLCPFO
WH8VRoQWioKLWTEZm9UblTEdk30bbqOqBPZrvu3VTYH4b8D23uMosk5w8IDKlfKQ
AmZsg6FLsyMyBKl9SW//+qeHsrGaBgFBdevFvEs3wWLohqEc3+JWLv2tqiE3Wb/4
PK9NAzMvdPV+OYOntr+2zPFsbu0OYNnO+BGpX0eOlpaP4Bo0/peqDYHXTwCj1E4I
rBN0alUiIXai35RzovrUvp5Tem6tTqKcroeHcEoEbN6dgYGOhheyAyD979XTLSLt
AATbRAgznLduyq0hIFvOBZTi0G7c5lahPlvsCGRkTiCzIshPsl73yftiHHmJCUOW
baRjsMLMUEvSozMDU+AjXYAh6UzhKHh0UAHIZVw6apIwq6lZdVOqw6JBAD0RPlY1
nMphUdFmKjPgEMJN5e2vzPR0zpIFIoJ3FMr9dTPhNjgM4QYWrccToJg3iQm8Hqxs
CgSmVlAL+b0mDlxPV1ZNGRXuavcOOyEn6/nVwo472Fgl2NZteLP8w9332BsAjOLo
unS8c1H5ZqogDiAU2yhGQkcJv7csvUjQt8toI18va4FwONW6twvCELXlChAHIYlu
DUZzDXMsIQkYXHB7ODL6UHoYWYOXXwnvgaOifWVR30BjzCFPcYg5UzJL4FlkWMnN
Dq8lB8Zyc2CLBeTUZC7HtdBrrlwxnvtmnvXe276XryDxYhqbz2A8CRFan9RCiu2P
1olcFuNC2iTAaOAvTG/aSNLaKWrhR3ZUW7O/ZgpZuASQBeVjQxRmXa2SX+PRiZ9L
bh0+59eg4iDxR+r+H3aAG25tIvZocxGfyGTSCzd83gp1MMOlzM99T2A99cweTMdP
5904x4hJbtuWdBjho1TV/GVi/EAnmHek4hHO065zXYn2yVMPibeWfLZrGwxNcMeA
mI15hT6sdUr8M7wb82ey0JCxVYTj54A9pZv2EScmQdsES2a8xpjRrF6za1wEvLi2
jz1jIJrDwFJwCvvdMvhXMrGMyRUfnmDO/Q9fy4CBth0kDU5duf9Ctzc1kPuworGe
+/t9NjY8Fl5Xa2gxh6o6+Lt1ivSY/lYNVcbQJnOQrEQwA5vCvs8ArFBHj9ftz2Z5
MFsGIuWTETaGZNc4TZgmOh3UTpot0cchdNeJPbfs1D2DMkgRSQ+ArNzRzqxv/z/t
QsfoD96FBxjUgmydInHa9z9aDUq74kN+DWlgYKdbcCQKF6/CHRmktRp6BEpp5Kji
z2cbZvkoXYKbNw6v3FFcr7PfLTW5seYPyUkdaHxn9A219G7QWDvu0pLNpd5ujXeG
5WvVWBgBvLTa+jkNjW/OlC3rRfzLqwVMjbiwdSdWMLMG9rOvxGWi5bQkXkyGCu86
OArJUAeVZmSDireq7WfM4yGVkmtzUEv5LdhrgcdrBVNZHg+ThWgCDh7OFlzrykQI
rUa3afIUWsEwlaXSHtunJx/GOejRgopTrWwqeedB5fUtNNeKE1rmWMPQGpzFPEv+
xtQJF2tQqnYZlQ+A4tVvnQbcnbJBwwwgpIzOo2OQX+s9zSTrePq/O7xJVHj8QmCK
WyqMTs6SPzf7Cgcng5queRDj2Q1ijiE3PlBmq3eFgH3fMgY6SOhgIXVMPFiipf7v
ohbrVSCdo+5lsxY4Ouk98deuMfiAjkD3qcVtBtcjrgduF28hP8F9vqE1l0gnzSJy
Ae85vARFPkMdFW15JLWcO61X9Nt5fmoMe72uPFXNGtDvJ6RrnV6pMlsXSbtuX+2/
l771o/UKQXjz8ZHdfuigp/uX5bbKEx52EOcTNcTE+TEPge5jKJQES8pSBWUFHHrN
AbxLamM+y/NPcNTIk7TlUhsBDa+ERXBsUbBjDlm2nAJrq8Zf+RVANBxLNIAT8p4m
JCrr2U8V/LHmo/Ioe/zEbiRN4FHGSFtVe2EaMV357aM8wr/KfAwAVJgOBQtruEYV
/jR0aX7iW9kJu5W5SAVCkKW/XdMj1ZSpntJhwoddqj7NJwBLDcUmVZ1SywBq29t2
WpYgf37BQKXrB4sEODAhQDBp6C859E3vpHhfgWYFBr9H5h2DTn8bCn991kXCnGx0
LavB6Q4JJCHIU12mJHvF6zlYYDR5pxb5Jn/PuuKFtnSA9P3PX7eWCt+xMhZlhUGC
FF7QwbJFqeJ5SdMHF1TYzc6rcnKofMC7Nbr0EP/5wZnOFIaM86nglY7bGdqKAZiV
7rvcPujFWax/23bO/TTAUDW6UOLkZKT23J0+vlOJMMF5CwK13gU9W7cc3NnQkn0Z
CBKvzXbr0yLlTlM5cP69yA4cV5CgQZWgMAdI3nLzcFT8hFdARXKylDtinXk2zHtb
S0/946dC2Hi1BzpBxcg9CFrg9DnKTrhnLspwrtiWSJsFKFVESgz5rstQDSvNSw5H
DZL2SBSnclqNKPduBfQbOnQPyn0J8Z/UWU+seKfKUH1InBjV+O52E8fZwsNTphNz
nIMGAOx7YANsUHQtkIosjsGh/Fc998A1CLHDapbW2ISsd6RTfCARoDFOobu2Lb3E
UOIGp6xuu3ld0sEGbVGCxj79dQCsRTyTyTVEQ0QTfKuUaP77pVtfNN0/dOknMu9T
KAGdCjN+mqxqSLAldK26tKp8nmk9yXodLF/wxa+V0RDUC64gBaIu5RdTkglcQVNg
nDv8JLLvh5oTTd50FipPooxpCAkMO51OTXuSKYwqjTenxnkaGyYtnel6YAQ8GWgS
ZEOjxnrTG6hAMTTpWjORK/JtmmLvnpqJDTnHazof1AErEmMCaf4V4ocCHN+XwQhj
1RFFak1C9TWDpcjmb4kZMHIKo0Q7iVmOF8KWO7ujTNCyqgp/m9ADw2RBQeGjF19Z
f2bzZoPb2zsSy0MhabcSz8jyFNLgBsNDhvBUASk84KRbUYu8WqdUgmOgdSc+faUL
MwnD/SoXofSbOIBVdBSx1i9P08LUTGZAGhAya8dgralzWW4jqmNyGr9/Zz0vLBPP
qJbV+3C24zqVMFV8YfhpQ5WYrdn5RvPbO14DT71vX4NU6fjO/jtpiOBpMiGQBFuY
YiQ+5MMtJiO6ReYFF+X1RxiavqjWzAqAVlH8qsmRxc0PfB1a9PxdOWgNKAPqHqyf
nNLk7rIKY2MPGe1UEErMNF+8gzJZcQPtsREm+E5bQlhiMw9bc4JLRym0A32vvClJ
UBCv0zV0Ka7yWH+lGBpBTrMfMqCoPvT+UKUT6MdoFIkqkczHXO6Qdj7O2pEyG7Ms
4ISpI/KGcFese0Bxslc+IKDOtALFIjw1xi3Hhj0XUlB+Y+ekLPgu4MtlRsJRbX3W
3MnL762N6ExeTS8Hx0ZG8mU+wG+66Ev7Wtg5AEKWFcdGO+lyR+iLYGw1ECSkdga7
3PvouRVO+E9MQi+NPGAHDPpFv3ZuO+1y50J6eHKMRRlV8lOG0arF7pMBvNjjWe/n
D6vtZoQYPhkkbj2/pIVPG2l3btXkVqQoNz862tMyeK7/fsJ5VjKFqeB80EiZykob
CVaimRGVk0KnZKLlaKndAURj/YjvhSthX28VxVztjx3TLXEqUMDUwDDEeKP5qxYy
kJuxOc3GFDoOfsojQlUBkLG9Upk1nKa5shSlaILygdjiijtiVPAaXWGemPQ1bKk1
yqoxVmQw0QPCRfHt5C6cGCg+JwVONYBGN800FV35K2I/flRx3xLoGQgtdsNdx2n5
rSO4SkFs5/NQDkp28AeMiQyL7ECwQBo+mPkyLlYZ6CDnj0LcQvn/1MMCw5ME++kH
8xTU19hqaRwtXpIGXhOe6h1u4VDwEe+cI4Btqgd2IRFj19GtdWjkTWvcdEC8VwLy
4MDmOsxoYjcWw3F1iZzOP7Hv4ggpWA2t/v6wDaRcsyFaGdi0pZr8XfA0uyu6U0Jc
pLl4SJXK+WiGsPHxYkMJxSKfRZ7IphCDW4Zr8a4bBzi/8yI+REvNcYQzz/QVax06
ww8PRaHm+8eKHUSLwQWJ1IkMhUwRY7clN5BomPtFM9Fp6kpVoO+D/ZgghMEowh3N
8jrVGldrusxDeKmx7EYBblLNYey/ifBn+FxA6junLEks81VWQvp0/bvO2P5Qx8Qj
u1EYuRfKTMb9b2F2jempORGcplJ+FJn4nG4gSUgwO7bvSOBTjcyB2aTICsIAoPrI
ar4qHDtELrqud1+Vs1rqA3jnnWlu2ybDZ2UmdUzHLy+2xXJlO4aArj+3RE21kO7g
Iv5+ryVrw4TTSVfgPeAq3I777+CCr6UbMksrxnGnBReXrVjesNKH029QjRVKKCPl
5rHx6UKDPNup4CY41pANYEBFe0/+/oQGncwmAUmtFCmE949qlxGluHtf9ltTnhV+
pIviDE+APyuXvwwKNP2yhLWy/cexAgIyd6wRyUKakyDT7xdK0U2X11ZJ8zv2Ybdt
9igh23h8BXqKHq5/vlefRH444ukT2kcsEqCbw7jY/hcX3gPbGyRpa7tKnlx2cMe8
MTehsvATWy/uMi++b01wdwihrIBFF6krPPi6jhyF7ijvOYLdYwDDxJQEiM4GTZh9
aM1/659u1KGENJFMc03yr5J3K8IDHsMHP/l0FNC2p8Hh9aJfdi50aLj0MXr/Yos5
qfoOGj8YGLyMwGPockaUveiqinWxGQEG8LOtkzCIA4XTceev8ioQ3TQZg9QXmb9L
44WjfxiMog04NybScOZG1LiqDfWkoGvf3WmL3n45BxBsuPatOU+/Qr/hgN7axdoR
ZogREuxralFAw5fT6HSC5Hp9n0yAat3DQL4nXjuPRSayOKFekYW91x7ej3Vpfsf7
aI9OqyebgTdn0Za8+cnVvJDZ0JQl7pKOP/x6bSkyCdAb44RQrYajtJ2RJsW6lb7u
0Cxr3v5oFzaKhnBI8JWTjyJs4jkCq1tjMp/Sm0DnNfos0do9lUn7MseVnV4c/YfU
cM9O+9XhpVc/btEUXNkUY2yZnCEKxWQegLvP4HEfc6/Oej4EdVAQnMVxWCPEa5IY
J1iW9mYnqMQqeGX+9M3cRXGF0FE44KDAZ9/Hr8w6Ew3HQdCa39/ycA2VygE2bvDb
dsgmOxGnBVkZ62VrG/wxk1MIzl/tvkAn36hmlTKcEtOhkM5qABIDiaVKExYNkbHg
6bDOq6h9PqbM7L3g4YRosb/y1AV+4nj/pnL/Ns43XKPpKfUXyawsm3LgV0yBtc1v
7P7vcz6B6e3TP6fP7ZZvr5S/vAE4TlNymc88DHgxH9NjrmhW0L5ZIhVvCfi5zlX5
RYDsLVE+U+NnwlSaWctKpMt5JLxdhW5DWvFGnmnAEHMM6xjJX1uxHpwSmlUj/uhf
n9JyJ0GPpLb1xHUfj3rYU/PczDIVzKmeggQrI/Ml8T44etHjGDIi1QvPY/1F+UIL
Fq8yTcrvpponZ8p1vA3VfTqGzWfZwO5wiPK9/QfAJWtGd4C6ei1M2iGcmvXl62dY
XC8Uv/CFmG5WVnhSqD/kkX3rZRPIena2H8qX8V2cyyE75panD5FchO9pmKeSTRGl
FR2sDh2/ZjMa35KZrlKxsEAp2QBwWij0wG9H5GnZ8dJcdQxmzBzlhqiCunoGwKxw
pBLQYVieWuIg2DqzM+vT2TYMOYSVMOmluKcnIVgG6hlI9XgWoMBqSyCgUfRDn9j9
5P18PP8ZXUbrAnxNwIt0LLTgkYEHZL288ISBb6Xk9rLZkAj2yzUVMKqbc0vxpNSX
UcdrkSw4NChQN2+5TNXVKqOp1LaUa08E2n8GRzNIePcc+tAL53oMSu+TAZxzuFUJ
q+a59lga4iKDlpCt7SKoDBEG+FNY6JqbA9BfpmqjCBhGLcr8kOthkfKN9SgOcgLF
sAZyzzUesAbU5/cb7cqyw4YK5hAzBB+tptQttM6Zb+4TSDYcw0ANDBLfCQ0FXyiU
qZ4N0ntajx3F7tpTplaTanae+dDNf9z4gYNTUOh4esJAwoBfdXDCBWy1diyvSpNW
IbX4axOE3a51OXbH+efu9hg2fvneeNhFmrk53IpAVrmGvB5w1Wci96lMA+UK2REy
rc5TXMR4AEdjW4pL2TiQnpWt1+bSHiXPMb1HsKEh0naK5hhEH2cGDf8kmqO9+rz2
J4dJWvAQ+LQFUueUN8OHEcNS7NXqLLwjgCXQqA20WH7r5I76w5kF3BRK/trtIu81
oxIe1mYaygUCJdoOofHl5Yhfwy/HrOHZ9BNgq17BF92GdZZ7z4IKsJDDXD1qcRuB
nx2QOz4qsaRjRgAY3RCYqs/vIWjL1G3y3QwlXTDMuP5TdGLo+6BsOywALfmXrJjz
huriCSPNa4mKuwwZi59pQ7/rzsP5vpTC1YcU8MUxCn6s3EnadKzqMUXDpsKxjEUi
7v8CM3lV84E2VcpwImPxanXEnZS7K0MtmPbcMjX39/VvPksw2vKvs995RaKGwGyV
kDF/asw0Dqqu3lVXQdiAKjW3PsjdCY+nPGPqH6bPf0d3CG1h5Wa35zoOrCzRc+FO
NkCogu7eIPidsFDlQfaDguSMyl2V0Yn20wqd9ESvX8H4Pgrxu4CJAXGTd089Hr/f
7UWfVFNGHiPaWCkhBWjB3s8mfcGGgnGQ5E3ofU01wojRm13B6ao6ThOhYlBQpRpZ
u16rxBNXrx+xTiDD0iNqR31mZXhpFlHDVv2zKJCanwBOuiAa/z7nm+OqIgQO1oSu
qlh4eLiF1unvfFk0Rmidxj41ad3AwTDIgF/RqYNWQgw53fdf1koKYbIE2UP8UTjl
waxhzjnBHzGcRI3yhhW9m38nmlMXs/OMz9MQw4BURa/RGBLT0sTBeBghDEFI0nFA
CQn0tNr1Bejeh89ra8lDrMxVV4yR7FtUNRr/RO7V7S7M9Pk6WSJUMvXvhsh6UCbn
hyWQy2xcH0cVMIvEgQeRM0r2D/G9bsc+ZLyrPZHCrxX91uwBeGptmvv0oVfHRmsl
TsunP7P3XqAAySXy9huQxeeXlUZIgwBmjKacNsEGpYPqac0TQx3gX6ZB6srUOyVf
IsKvf8TsqfA9kV3V0BncN8/1srTW7mfuXNhuNunHPe/6Bz9dXOO+inSXNO3tOLVJ
29c+7MeTcJ+xXVeA6lfHhZFm/BYqogNQYh9uNmtS1bA2+pwL9VNt5K9s7YoE0ITT
iSFE5lvXmThkfRZ+nAt9NUXFkNKmNSZ4x/7/aKHBO+3A0HfF57K768Q6DNHRkOOr
39j8IQ5opfaHy8NtbsN8CF52KhIS2hIU3uuLzMROwriZgDxbbnLPjKBX/TFugNQp
iEF5/z/l9vo2ImaJgh9NhOOEQLa2OHJqY+DE+zHzkmACGMTQJdanonAHflIXnyOL
SwrOTebsJ4tKi60nC0Rkt+QxkPb5fXkH/4bj1/0AcmEqIIkj6MSNgW4pVaOl4n4+
3EJHAJBEr08vO6FGhxEVjmLvu1CTNgVE8eu+PxzXrc5ooAlIHD5bBYWZ5qy/nhTq
i8xSfHBETZI1QI4FqIpvrEWY0fEv2h3teJINg1BdL0aFKnebm5d98xUQ/+WBXMtm
kL99YTbQCrvwXI0gVktjlvNS7E1S4ePJrXt1VSejAqFbt4bUv/RH+ArEMw9gpqxL
qRvLHFl+TsGLxF2MQlkRyR3is6X5i7iucmGxEN8EvPWtTPYPTky/usN3YRchSG1t
QYd3baPZArdbNuOD72wXZdjWqgZzdkI75ymUYva6nXlwsY55lLq8uv3IzK+PC4Au
tujLqemDARGz5AJPbA1LcTz4R3c6EgMcnxDTHGDnXzL3FFUvt6d2zZec7FkOqEyw
aDROu2DFdAdXmDGYf2vH6h4DuTBegCMa28JH2GONJAE+NM1TmAtSchltASbiYZbg
3aQMvlYHB0GHPJv6lq5KoJUM5domZUXp9LrorYKQmnKdvd7Q/gX7U/lgoPr/CS0t
Ru9VBC6xk8NxhWaNEb6unE8w/kcd97moWhaHlHuPo8ikdPVq7ysUw5ztaYxULXOS
Lx19KKGsdpGKILa/zsMte1nYtyGfkAOs4x4ccGygFm5f4wGX4LFwm/8e3GtYP1Yj
dzL5OU2SgpsG1/RELJSTDhfNdPY6jSiDZ6sHEdTrT1n1pIEqu3UDAW5hw54ptoow
kFW91wqKaDFyfFoWCrZbbDRYVsQYRHG3zObT8tPAxQtjgwsonw754wsJC5J1fyR0
62goYpelziBhs7kJXIYAX1IM9a5FqzBh984WJx5/+pNILOxep/Q8AH02XhGvxXAz
GXJSuo/FZbsIrsPb/58ohO8e61eznmry6DFoG1gqd5sdEdAVog6ZJgbCrM+IsrRJ
2n9zOWn5TCMtJjb0X0qbjMO13M8dFbqZSMsHw3V/nVqVXYsND+Z0INwWHoLkiz5b
v8SrbD9nDQHIWJC7NeBq3z8a0EkycdeHb5rkEpVFIoR5VbVy7Z5xh8Pm3/8QOXit
XcZA+dlzKpeV8muSn8597NswwrrsR1ZeQnuk63LubJuvjdpmfRwPOT+8qEFR7UOd
vqsJpgQYqqEsmVR2MvatCNWdopFRCNHlph3y9mi4puLVXZtikuBHm6/xs+o1Xubo
7C+QCUlVyb5fkEPpolqgbL05bi8PsZ9NmyzezQW0IJcuonWw+sW4JFxnvNBebYYL
CzB4PyPcp6p5sMPT9fyR5YtqD61fhLBBwY9k5GWfIcxc/v7rcpoVhu435jGxghMk
yxzjPZMgFjA/QqwxWgZPV9TEZfH5GGQSjfOH9w+4xDudQqKk0EievTe98I/NJ/0n
EBRjrUMhWLDRYJ4za0CIdi/mvphlh8Uvn2OMt0nk//nHo5hTOEmVjZC6BRGaXDBh
V+ScqD72Fp1nvTBhJetQOygVA+kPCjbScb47h+4zNACSrBYwR1g2VHbt1pUeIa1j
jemwBtEZ1z/pX90us6it8jAZt1lnlIbhcR6RUHQR6VWriLg41zW2nUGwbFKIsKj6
qM9YI/g/gITG866MBxzLlXxUKWWG3uujnu+/WFGiYtPxtFkN0/7ae22ezwPU2Sxe
r+gc7K3H54sNneb2GAohjHOfWdmYUzHKv5DDITsThCJpS2jcL8coTp6Nx29FZ/eF
dnXhNA8w/6mD7twfv1nL9KPXkTFa4+yruW8NFsKZHdZc6qUH0BpxmFcoe6YGhIWX
MTteid+GsfohQU6nE5+Trj3je9OAfi2RGg+rk5BYWzUq40Vvc6kfoyYVqQTZYqV3
q3U3u7A/tJ5kC0UKHG1fsOuB0PtsDXmwEMEpLK1lfrZLMyVlDByIhfhIT43taPZq
VvRbE/Yh5/XXKWs96DowoPhSm3VM14kXmwPifEYD0GgFfiiRa1Fd7cx6aWp2/G12
AbrPyQ6d0KbxFL/tAhU1e9QmbOgKy3XrMrc7/tByQznLfcwxSQC2ZU3eCcUV+EeS
OJPbxWFd1vOIYsvy874cuPUB/KFD7y1ZZSl4uBPHZKVQ09IsqFH8eEn1eYOZDFnx
eijbjsjfV+9N5SmhLSuwI/Rwf8q6sVj5uuBApBphooODYHXGtI91KLxb2kGX1CBX
X946tr5c8Wluv0Mx5mZrxH+k0xOc++iYTHVZcGDhVU6b5xOK8VLLEODyBW41Mbv3
Ex/h5FEBEJx8t6YVHm4a60jJ12emRzY2pMaDwLAJV/wVCe+Z1cH65MId4YNoTk3Y
cnL5j6WW6kzNT6woU4b3+CAAecoiuJXkHxjgRFqlbN/L/b+FMrQQd3QTHN+VgY9g
kXTGzntNqF4UVt6YFJilENIGfx/7AdvVOR0w3naDKFGLoWA0YlbGcLz6Za6ujBfT
BFrA4O6toT3UndeJpuHNP8Ind5ydzN1BJbkp+Vb2hinm2LEcLa6ZEAykSQyTLKuP
eHJlVWj1VRf2K0cLMF/c5ZGG7nAgDQ51hpoPV3tR7lNS6fYw1ylVbPbTO4Zt9Aur
PExaV255S3cXaiE23Va9knArukkZDQCmADFam57lpW+k9VND2Tzc8w9gmoD1ICi9
a5BGmFAcRTLyUhubw4Xqt5o1IHN8KEGuG+Qlsn/729Akzg/H/Zp9UZDFhWQNCDiT
UMTpH4DuMYLKs9K+2Gwi/9XGKaoB9kF4bBsb8uJGTpJOaW1UM5/IkQM8zBFHqZq5
3V8B//tNisWqEZD99CxnI5in+IzVN1i9f6aODlcJ4riyn3cFME/0Wr1bnAx96kr7
nwFrlkb0bkQkNZreplA5a9ct5laympeuJ4CyIY9YiPfV7O13K/BmuDuC9Yi/4lbt
1C+2P3fK3ULJ3c52hj8YNXO21jDLAZerA9XJILIhXsXlsBXYgQ2EeQ3FWiLsA5S6
CW/56EJT1HEUcnzKkphMBYvUgCIimna/0BVgxPSsy/phTlgSoqpI/lvOZ3iBFd2u
yNy3HytUJAdjgJoTUwv3hA9R/2lYN/eNXkNq6pvdrDkKK0KEjZoJDag+zePlWuWT
HJpf4HkTMaqYFHdn5c3CRPV/ztUnh29xo8m7EQKySR9VCq6gZwh5nDHdTD58Ro9y
d8IHMlD6/0Y84ddr0Sa7qv4Qclo5uk9gEQgSPRdKyGB9R1GavYAoXERFYEgMpbkv
l1qXCYdprMtD9JtzbUoNK4P888DOGDtCXn6m6cI9lcihFnw1ApjVZyUrX85xu8hs
wFlbAXARe2JnXkXhmac3dnUdwyID865RrXlcrqL4ZgAvyZuhWFjV33Xwvn7uE/X7
gEuDBcTsIK/GCpE8G1uXmIDmdAzujiW8TYChEgoLSzv7XMkby1smi6Jpp0wo2Z62
NHeiIDyzhOWLOXPiQfy6tWVwvi9Xtk7jIfqXuDUduii+w4c3M6KtmRQlte1tV+eB
tMKNCjfQCXrMFPFd6Hvb4fc4ZcYr5pRhsYt0AD1PHAwlyMLv6/KONuIGAtg8i2Z7
OXFVcgCzuuQmEMu/zP765SVDThDDv56pY8sRynAxdSNPVodMN6eJrwCIrWP9X5kU
MJ3453MecRgV5HyTbRuYNxoC8vl78Kvh+rEvlIWkUHQUWisE+1Gay5e3IKILopMH
+UwEuejyZnl2c2X2mCC4mvh/AKvyjn2i5Oq6SsJ01d+GPycjOKdPRVcScGbyZl76
xhMsbimAbhvgi1Nub2TyI+kzZVg9/uJn+JcvI3CWG+ao8NPogALIQK+23/hRnXoX
uUC877/NGNe87YVaIoG2XLQ4zD9B7vhSUf7zCQCd1qaatgSky4n96/9LqA8+I86n
SYJODS9sJY2evrJdzBNG6LC8OUTb/Zl+IwKz09read1v+0cWj/pD+A1YTfhXGlMI
zwULG9cE4nvCjTYwiKWor/0/x4t34NdKeOxZ0NVOIZvF+qOXlTK+NBVbnvSKm1Dv
E8KPT+ahqXgOjMRzPm5yndTzzIYarCmHdekkEk3uMXiWa05tLrmXQv9YeOB37yzy
lqChh4g+gDy7JLda56m4gp1NcLyeCMdR0UIamR4rc2mVIjqtxUvSGTAB0ArPE3oo
rFfOB2y0e3pKDoegs4TuzjbvK27bmHvUbecQXn0coB2iUSOGjpA8geKIHHOZvoQf
3k8Nz8+JIOy5H+4/6dG1dBYGuKx5pGwaOFinJ6Hj7iDQowgBK4cx44K94aNA93Aq
dtX6/uzWefzWBs9oA2zIYvP3ULnCKJNIdTO/KCrAZCxwnrevz7TIlp2o6YQmMQua
dILgXoSJQM9DjO76lq5hm7NKLoib6Hew+RmvkUvUoJfQxThnD/cDjtiLT0SmHTij
bxPStab0A15+/sY7YWf6fgKooPVyIjuncvswOTc5RUybpCTsXeKW9GBp80Rw99Sh
LuS4zndEA2E2rMcZVtPJRPVCBGjSroorE/vPRfQ7LJnZkgcvLc5mNIfkxxI8L20o
DtK/JhmIQutDCS3Nb5vKQhgq54bx9Y+14PNxSgFhmrw+ulh9DBIUIX79Pfz+N6Cr
gCNnPc33qbdc+VMQpd5Nt8txdLjhsfpe+P02BrVImeETtK+Pzy0Up5uOOZhiDdLt
DXG8jLCtdo8zC4REmaxM7rbNvqupWJm5m0os6z8obbReg2zWMp5sVeqgxZRhg+2j
WFMlh6OhFdHnyNhEMAjjF08zAzt8+RVC71JiR/cXCLNqtE6xe/hz4iJHjJcEiJWL
8Mk7cphCeSeEXzk5LrrrD+kPKMDvaXA7ML3YKD9VqkqK99h9Mlk6aH5+et8uRr9c
UUIM+VJHAAreut6Kd4+PuK5St0WCJAUpF9fLMpvkjKXm8x2h3msZfYrHkeLqOPd8
0yof7Ty7Bx6bKGu9acp0My05PBqL9nDaAuqe8V2laJ4shNVS05zuAtTBQJwDyaAR
b+U5A0RdSfV7kBx6WCVFduu3X0DYj1/Eo87mNCR+ooTUlGWyYQZB+ZmVGbMy5Mbm
7h4KLPE2fmzgaRYU6PaKjDDAHfoXEwTAtnWKIuEDYcQkgTSMOf8VnhC/o0mnZ4aG
a39TjOpXJSkT6KAv3YcZg705tipgU1OFFg0nddtCwqBJoWY7DvVRZ2XKyBWAy6Bg
udu20lOHLOKNSnthojaHnQj6DvhCqsI45flu4BGRuRNdlPVieDTgrO412yTw1roA
doxVHssnA451nXwdD6EppXJQxayZR/Gh7aDwaVwcQDMcXS0nDY3NKMGHF3zdqunl
eWykmPhyRxgCscoRQLTyF+huLVXboEygyNyL5BpoYfvx6XHgEi31D9ApPdKkp3SQ
YL9KoyzjmtYv2wuBFGAZk335nJXlX6BLfnBGRZ4/6dkvdMMIode5iZc5OmD/f94m
vC88hzoiEklX0kgUsmzAtHakHm66F4tea80nhGGVb+PkVd6D7iStDCrkd82+hadC
mzcyvUdZygzJBqA6hhWIYL7EKcPgbqLLohL+RXmV4yDDpNxD+5ibYSdEb2XRr6jW
Ko9vsF8C2K6Dg3z216pS6LWIYL/+w1ycWiZKDoW1wtVqU/pSmKBuQePWfQ3lnCrA
MeHg6SfIkN08WY6Qqb9ceeCURez/zvhH4jPOXWqWftQvZy/ZwS84s4P+2LKdsi6e
CyHGMyNImwJSs3iGzlXBCgxiRC3MjsqYjwvDCGxQeg3VRfwn6nphM3lfhov6BPL7
FxkDQmBBH6etgCmkcvn+KBds0/ivUNY0O1Oq2ISMFNOELB+e4yK99reRPw7PDUA2
EA3a8BIXu6geLYL2CeVIEFm/Rx2JCMV2YnNV6rMkWfjIqb6U+QyCKJ9swOGOXHXZ
tTBxj2qLN0+1ZoHgCEzqMoVx8Cx2kBLL59vxZCxVEcsPUelhdCE6jKC8rkhWKN2q
wsnFrrTevMAK/biJzUarinJCaBuyHlmrzQEcik2mA1z7ISBuMR3eXGFSZR65sH8T
W7g6RMolBYSLIGK4BuWDtPVFXhZtZaf8rj/4CFxKGlsrYikYz4+SENKzqUIndUF0
j/8mqZ03TKx2nWdhC6Fn2o/VEHshsZTdwKgx1NTfR3ipu/n6+MBqI4JwBQNdhoXC
8OoSMA1tzj+4WEVqBRUbHYKUfmJlq8rh+GHLEoC0w8/lJr4XjaZrbPPDpARLSpE/
NMSvCF3dUoArcfirsIVeBU5zkecPRm/04PjBUIXX0j0bHHxWiTmhQpuvnQyWR/em
t/fQm/JmtftsPzwGp1INR5L+KeGX9AHbR8CHPptRP5Lyxo0ydoQiIXplYguytSwW
VV8A5xvzgwiSGcR7ajlr2dcrwfH3wYzYt6jwpN37pGqS5p7vpW+y0V5wh0Bb3aI7
q3XbrPwRO3lDV4M3LItfY1bbnTmqfrFNpzDxo2jAkvDAEDyUAgx44CvXflagmL/x
7qcLVF02/jxvx0T/1OeK6ERaP+2sbNrbFHEAYhySxpcLEZ5Xi1PVYeYtYsFxhsyB
a2YtYEsaeBAZTtuSxHaDHPku+f+kL17BvWqx9NNtlA6EvyZbjBC4GM+3036JjEYU
alr43ygkZ7WJAY8dPh+0Ljo/FN+BAw+Uy/Brpki8gFFVbK0YApJngP4+o4VN9xmu
jkRrSiLaIr7W5Mi+KkSA36EMMAAzu4VIJ2mjmE/AwV/JbZOW8s8iPAvF54Gysb2c
bbR75zk0TPrxtTGYvQBM0/FW0kdJ31ogBllrbbAS5nDtYlwAagu7GEcx64jr9bfv
EhayhVdh2aAYI+Xjt7uX2aUw25m0IuDyEOC9ZxDPqDvcrHBxS33nzQcrCGWTyydh
wpzkrazaQzyctR4Gqb0RGC33xT0Jnknwk26DnEyIt3YmXIZ75mx0HKjz+GBSfKga
O1YJ2x+CCW7H6yPkWlIo4ukEWZYm5r8c0aOg2lOrtrEkfVrFX1LQM+/JAOszwipL
3oRlDkao8fsl+Be1ojIXDIn6f+Xo1QKeROZaoeUoAebzG7vAf9M0uIeF0z0oLlE0
bT9VUisqw5/KMaiEsFax6yiOrEA60T6oo0HhOQiq0OxEZAUinT7x/UVtz5ONOqAA
tioPevt/UzLzLgMbCM/aSNN/5KG1AnzaGUlezdrK4FdCaEmYnbWjIHY4iN/Uqgg/
TqxD447d4YC0b7feiBE4ZpMcwWQllOqxyhW4/gHTzPhOoA7VqE2utDda09pptwKD
ahy5Fp97FfJlh59OeOLgygd8ndFVYFmPJ70+VHxurAi8PFIi6YNQgSlhOYQbU4Z+
8Y6u2+wBgDDYO0FrptQnCLfzFZgmYcA/A4+P6Xy8IiJMozbS3bq1jwRrQXrGm+HN
W4Tn5AcxI0NWvZbv7aP1HtlfmW2T6s06NNlVC9Z6sD2PeFGDg+BX+ibqJG4xZpK7
BZS2M+ryoNaFG2bsiUc9XZN7qcya0+jeXLfOWPKmJRMln5gwTgLf/TcriSNMQLO3
xwdstgfc1DkgTj9yiR8MF66g7hNhjQfem91KZE7tK5Y6K0WWViCEa+2SdobfYJSD
XxxAM93X/rrachNxc+yqmx78RX/PwFx1v3XvwilP9iukfbaRfKaxZCcza/Sxh2FU
2HEJZIGQzo0qORufok4+//4zAYkHwgtwM0E6BT8VvsUOHFkXq47Ri1P0TtdpeRiq
m7To0lH0vKyOypO9HgGeZLvzNBL3lHdX2gnl1mN5ddbwPk242lLxRvtHltq5IWae
B/6RTih2aOJiM8FhOZVfB3J6c1rpjhkBirAnP0ODtc6YRTrvhLEspJNKetdZl1z0
1h1VZo2KX4+TY/pXW7atlWQavQX8wNl5UpaahqZHuOgwGrOZEyJSfus5g1wI6ue/
IkUU9/pWSZZhBo94J8pnip3tqZGmL0l4efEL+Dpu7WyWJuIn/O8ILCnZD8HMR63i
PHrZZannGV+2zyoy+oJvtVtvTjES3NHMEPmnMgab6ainxUNkxUrI+n1iwFG4YDiA
ruqP3VpyzkmrZIldb/akOHNixusZaTaMxyOn+Vm5+sYvrpQYC8Q0eolgjbi4zyKE
K8PH4JsNvc8K8aPpFugS0TOnm9CWP/a60Ty2oZGfcqBUdiyoyV5TRg5HoX9BsJma
oArzi4bIsrTs1k1pKnovZK57qlF92yIUiIKrqPJW4pZTquQS3BxDXiIg9/Fw+9Hy
GnMyvakq1/2IDaN7FNPU6BXAVoTOVT4QxHpK5X4Nky4vuNP/7hQqc70DyVmJ40uS
h14Lh+req+bsASPbF5HFnDeQ5Qy5ls3H+ZelupXjExf6TcImBs8CUf6Rz25LpkcA
54Kxz1+dT3rQc7+ZDrwG2M2eB4890QqM3aZ8SLn/uEE8Nox1X0GcsL1AaZDaahA/
9oNwZv9zd7a55NgXebo46TVS4s4gWD8slSBL8+jxYB4BNLZ3jqrC5xgWGWHJHof0
WCWeMP0DiA8PUenlCqMEkHIQuQ5Img3oHIZLe1pmX5eIZSI6R+hLpU24Vhl8NlRL
ZN0Fs4qAF8FMlzQ15E/CThJ/mIQlja4QrjOVzOr4tV2OMU2NB2bb3vsgUfdAGUQw
U2ONncuwKTtbl5py2xQ6kUvnueo5TaISCOf4rbV+gWuBqI1lSoZA9l9FKq0lFsW5
VdMOp4l7k/bDHyYGQrMZyKffkcSkRGp0NDbiGBZzybHqYYTRfkl8AxNuyYX0PsrT
MuVRvHUprs49dhuhhKEK2OFswXsgl6fn/M0wD/WVFjX9bEwhvUqFUOYBg8aneAj8
3HCOBBllUW5trmbjQ9YKML+jZzWMMX8wMTDGIKG2UTjpdNBKitg49GgxmZs9GgGb
dK/D1SMBINICEApO9b+zyfzU2sjV+s5i+j/HzlQmGPLDFwUQiaDzZfSGF98gwFzM
HE6w4s1Jq57SMCzQ2zBCzOfw2HO6pLNj/podAu3CnXvpNGKOST3X9qbxRfBRz/Lf
U243j5Y6PJ/pTvg1FxBruq3IzztVkiR5vQl6D25ZC3PCXUmsrUlJMk8o1ZC+fNMV
umBiU4MhfVO71e7ePl6Sto5xsf15AcL1jDDdJOB89PTVMcQ2Hw+6AY8s0r2/XktH
KPk3Av4D0EigFeBiBPLQmERnrGRyrAbfRXqVW334K/RNfPLECCYQJ2jisgfjKvm2
cC/rG0m9M5TSW9jO2EdemnA3C5lTGCREImXnfxiQFQno2hi4K8Kx/Rt8033A/eqa
u+SA2lhrCrtdd4LAXMY+7PLvK8fXOyxSKfU43M6JBb+jfhvgqI6O7rR1yqHDOgrE
T4QGX4YCxZpN0JDQOP2fp2kQFlrjBJDsPynzZAlRgo8L2jyiSq7iAJC0+xHSmYeM
NHjmUvlMH3w0dOJQUvUjpsb8NTKTpyfUYAZx2M1XE/RZ4pJAqtEB+nAWy1sE/7+g
p9I4lyDxS7pRWa4Ks3cc+H4UPK2+vOmK2wj9YwC2EZeRMDfiuaYZp0FeJDT+2umu
RBNcBCzhKhjcq8M7saY3/9DM64wRdsdvOTtRCAvOzamy+MCKNMmHIrplyVQZNoW9
RfczBQ9lOMJ9t9uqNu8D51aryfgG1xSb/IUChitFSZ6FXyQC2kAk8/ORQ86ghIKz
qirbiGhvwPT8sJMnqgZtm46sapscn0DGivut2Mo0zVaguSMQofsyx/TbNpflJZJQ
/cEhRkr3WRD7qVHhm8IDwSqOSVqxDEfZlLS4RLj1c1wu8761be5rbCAceuU0dNfv
hXRstBl/qB7wsCTvtK7arTYjs6asJKTJi15qPJAmbxJE7B4UXw7vf5IAuhHpTzwh
djdQ4q2w0jF+5k0IOij8Uc3E+r201zDd8WOCgyqi5t1I0/UYhSfOZlRCqK+Y02cc
8vpNxp/oXfyVEZCGZo5twKxW46KITNWJIP4/nqzfcfq/why8v5JAfRgD5k9bhg4p
93/sdwSKDPmPCHcXYTqNuBKeVpLsq2B1XBEtHs9w/7B31iMNY5JDHXOt0bG9TWxg
t3fJ5mAkEqlq9VIjpS0AqezvzgEs0y4wn2VAo7K3O1Y4mBCuduG/pORS5cfF0UEz
L47nKc9louZAzm7UUu4LoNmmnNtyFlVWvLoZey6FFX2Dis/nIKic+yBUM2JmUl7s
KzppWuJ8IGUMmEO7RrWpZ/Dit27SHtek/R5sTt9jRFIByXnOgl8JZVBj0Xj2F1dK
L8eoG89B6QqI8Vrv0jFqX0eEOOZhY1HAsPS/YKJPUdetZ+vGZ8f/aKdIHk9Wf7Cu
883bNRxNLrf0tGjgu8keP5NLsVGunCBHtG2hLQuKZe/AUyQCmC46sO3Vbr9k5xis
+ueBj1GTIJ8qw0X+JzuhOqaiM1tU/cXu4kdoZiZFq+/kJq2bYdMztn5e/BuHnUxn
x1Fm8UNZjUuNvFh4F5a+UyG0RkmZbG5fVfWkKCWfjlfbnYY+GyLJBMrRLNfmRfFx
N/P3tMk6x4oS9lyRVrfpLE3zcQ5usLcqdr20iBWuVArGuN17w/o4FRKeYkB1oavC
EKlPOPNNRvfKzinA/izZNuvRCiPZM9c7uDfgho01jd1PRYezvOiSD2yUL3QqWhNg
h+NzJ4febB1qr1C1BjDnHhG1EzpaOlHHyXWl9ihszbKrmPw03JlC99b5h2gNlbL4
4CpavtG4jnyBjnBIvfZ71UxkiuCuzXGvFhdwvtIQoT2uhM14tcJfQ0l0j+8s41tL
pY4BwBduwYhjA2xuKFrv3CIXvYAwyNjY0HU/x/QR8cneWYuXUoV+Q6in4xPBGNbY
fevZU3MebQWFQzQ8wNHOiIn3uuLUVcEXQ95XYvZouyJ+fPZnpBRyWs2kzpcVLMFG
FpBfuiMb/hqOqfm+Som6ktIf/HTQParM8Y+ZBMNzxDSv1eQT2mBJpIjEqOoBe2t0
Zim0K3Uut8dWLRPZC0PEJmGispPbmHkO5frO6XxC+vZAZ/ALjmi6nG952yAvkxq/
U5LzFYgqukRJUQCu3Fr9Pq0r2VSIBcPVrN53f9CHM7UwDg643Qskj68veSP9bIou
IfBjBXjKd9B1mpkiUeLHLqr1Sx7XdZn5ekkSAsR6k/OwCV0QseNyUvTIh+xV4Kmi
Rt5HQKi3IjDAisuqUY4Nxru8TrwVc+3+fJ4kekUAVCDthovOJlvnezfhvsO4djoq
SwfabV+uR4X6Cg/Pcwk6n3E525gSjGVOYjp/I6BLWU3jX5PM8pw2hAT+WCIr5Bfi
RCGob3gbKDDLpavV0DcAcB8uPVAL2ErMh92CrPixovvnmr+vtlN6hawsmBoCKM0q
F475b9Dyy4uVt6bMZvI8tsKe5w/qteDKx1NBTHvunWpmKcKCVYni9qM0U6y4Qirf
cwYiXLED+4QuQgMjpMLcltoNLqaLeNbP5sNSNIrQAEV2PK+OG3kbyDHSQ4RTGP/w
ur6kUwFgFpE+bTq26d6M9U02wYAWW2Nv9oJ/o2suubdlOVdg1dvw/XdO1ecq2LTr
tgQ0CKyRKoE/Gvi9QHloYbInQn9I1THuL7NwodnBLFKV5xMp9oOvz8lIJ8Rhq3kQ
YiDMYoB8Fnj+iwMJcmJpJUKUWfbBZW52vzJki0pfHdmR9EygDpXtGwvkVRdesjSq
fB7rOFif/WJwNPgKQHyNJu++yJUFfCEjqNG1HsON6bhSWsh902ymKXytEqY6dWdM
bLEJbAFcknH/kYhm4UHAu6GTq/rcCVZJ0UGQSKpIFjb1v4k5tYX4O4X2PKKq5JXU
Xr5v0BYIpxYCGDaSPALXUsgdjRDiGoyNIpUkHVKZnJ2kp00+MJQr+osH58gM+kLB
jcsZv+1qvGSIlnIip5l8kaqHgx4AKnXKIJokyfuNoBUtzqZyWrks3Yn94Ba7vu85
1kQ7PGdUrAGFvt5xxJRzB4aQcCUI7Knj7qgjL8DcfuCyuQ6dKi9oGim/wXLSE77G
qrqGzyJHb5OVFsVh3SFuZy3VtTIH8wHZ8KsGTUbdeI+JChfB4yN3I4y+G621h4RC
byLLUDw9dhqgShXAF7qonY8/y7ixo1dBwRkQqdtgSTGbcc40q77cFcBHjvk33GzX
AewZPhZ6E+3FHPuXm5Oi6mNUxPOP2B5Mw6thccKArt0/CSB6ofASRHc/4MYHZM4S
DRPXrdsi4NJQyMo9Ucn4W2UVZaDJm8PgoQhk4Vs6lYBwQo6vx0E9d70PyebLASpi
RzvxQLyGShgVpHJpnIx2O74Gb0+fn87/g3SfWjAFqxnO9aCpKBSuY6Tp+5L932u6
kPvrKpSHyhDOqwK3gygGUQ1Y0U1pQXIq/6eNjU4hWxRH1gkS5SOSXOqhClFUk7ut
07qLQCtvdDKlpZKJ1Au7rfdAR/+qt4H1HIjLJ8F+h/KHHRfpg8Wr5N+WC/8DMgBi
mVcPViLTUi8o/62NfDuNlOSO4Ef6eLAW7DZw58oLjB1zls342VxGRUPjgpwNdnM8
4GtbcuTscgsqi0rwpAWqkLPrRuukWYhcCj5dw7VclXAiHqnemlF+8Klv14Lb9pWy
4bhwcxRtfNCvCJYncvQtRJ3s9X9jPFWZoGR7cUkg22d6AdRN7vx4iFF3VEKHOl6j
MyPJJ83X+KlJhZca5VIkcKmWDgFuWYEe3TtBBxqcgo+6gGHcrUnLjIFJ0QUxrJwZ
ak+RFsAVZHN7uIxMuL50d8S22sakFLPNxJxQmdt/SEN6GsOn42sYqshQ40AGmStL
zjtYFk+ftKcO20SdH+zezw4HnLkwOzPBnYobwhXFuoJbcFRPRIbs1xQYTYSknYQx
6YVywQYsqJDrfXOruI+yReb4BmZK+L/gfuZv7F247wDMidRNDX7Ds0LY3f581POE
nJIvZNGuw0Jx+mxuqTCSXyW7gWCOAgLaSMv8VTVwWufI9arVRttEgHOF9ES3Vxs9
KdMdAGNSirb6NIotCZONv2f4zssXGftua2UrX/10pOLvuvfW7juT3H1T8bzlL+/j
XIs/LbiYedxGaV3PoUTDwCEfagQOXK8/fLBgijtddKhZi682BHWfOmffScGAne+9
Tmo4kysIe/av8fBHjtQ7y+3eH5RXtua9oqsMD95aY3W0sFfjz4EQbg3YpKk5wQNp
faPIVrx29Jra+Fp4pWEnsb/AnjoBeHML0qma4CoDuCEZfsbxfqxPmRxZk/ulQS8c
tnGef3pOb+2cG26Aw8dGsDNLVocbm5rKZyRm03EC4HlVIv3TT9dCBe5PzBEi9jzd
e4rQM/G7dtFFhWWVUco6ZlUJXXrV1Hnnl9eZkKo0TxgYPc63068dAwFB0gwVPHqG
u1ls64mIMrf261zW6LCACMFiAVO9pdv5J3glh2adsDhNunPdQCFs6azbEymv3yBP
eWhA9xEEZdEs7xi54xsQNfcYOjUAItbAF11AySw4S+OaGOZ2NbDryUwRie5WFMRm
4zDr25z4Jcf+GTYaqBhsZRq8uZVSCeuXsu1Op/pmqKBJoTDdI4QFowaMe8uU818W
39eUqnAb05SOCTcu2qBagu6OP42CwhV1CbAtbUNKPi3c/rP2CLmsF1QZzC1DalzV
JmzHpUISFoCdXy2FrlZBYj/FL6fuqQZ8umv/7xCr33Spuf4DVjb0EwJCjQ4O00Aq
FhEEJvMVMcxKrYIJuFEyGmotLb7kYFTOgLXMbCLgBJhdCEj5xQefmYv/4gmXFeAz
PqUsODaYq8a0FGqkp6uzwHmuZXvSPWIFZyBOe74jIOMk5jIRGzFxOg4e10zL/oYF
o45IswuMEKQg+OIeTVmBVHbuD/Go+tjaFuKA+dVlEWs/EMmLxK4/g5cNjMzGNMwS
NMF21Kp2oonDr8J25WzjFcYQbLB8Lqx8FzxMf+je0OvHiPGLuJQpLvWHKtz6ELze
F6bIVgVu8EgOv08X0GvQXJU8lRu9LKWFhBs/dOitlrTQ4Z5SVu3JT3PiMlmi2Ubk
T7K+Uk/xl80SdRgTiD7tV2UEYD0zxzZFEWwxYl/70CBfnTfgAzivLGoKmmmesTja
tOaBxb41tjUU220Q3y2z3zW8DQNhFYNN4ss9jCHhpxq4T2Ec8wQcmdtWJ4jhAiqE
+KqchaEgpa5hwIOIMCdiZEDuo6jTrjCUeWYIgKVcNeYJoTEJSPSV4IJBrnQ1+lCv
Kv6qfQj0bSuSPBrbhMUIZ2I0Fl2im+j9cS90fAWyVorR5v+MCBXI0I0hN+5nL3v+
NrfyPi/VfNl4PDzhX3dHX0s0Pibiey9sP/0R5wdXBB/mYikZBK/AS5kdqlSUNFkg
lDMsOPIXzWhavga9BPv0u0kNlX3bruTelB5KbnBBuZf8rquvTEWur/h1by04Ae4P
I9X06qs3YKaBDoDKw58r4VBB+7Mosvq6OGulDFlXl95pPaF2psZG6WBi7evrQjaw
lnwMKC+X6/Jx/k7ddzeWagLxZz7oePqNfC7lx9sbhDC09CT0+Z5Jg+FCw0L2FU3M
GaWLlUPl9bNxLDM2MHaeGL4glpOl/wftjDkr/bYCkUQ8pSqB9rNMTX6C+VmzPvI5
vgO82/moSPx35s0+sf4SiIUCB2/ikzZEYTs9nT/6RCmqTYkNyt4OgEVWVdeSUlln
oaO4dTuhQLXvJtI3JRzj8rC2wK4tKJI7lRSQGKlTBBdS9tLyb6lnvY3y1SMmUBZ9
i3JnmJLuVQDrjJaStfog6tXNAFE6UZQJ6nGYZCYuVdzYo0p8fk/9wxTflHLGlogd
sw665NRaeu76SK4obMXljJ9H2D0FNtsYiaQG6sB287dp3ACME2hnkDvgRQOPt0hg
N34WriCTdRc7X+YHElxUN8Cd8bGwRdfdAvHMkKtGYugGCAuwOMbPWhwviNTGxeXj
b3Fvgb6MisT4dyx48SfwS/8wumo52rl7mCe+B8lKOaKB3bhzUph9YHjlhW63/w5L
sBmfWU59US1cHL7GCheSW6ZATLeJi3sz0s9rXpHNqEikK+4rEOecBuhkjlRwdzfz
ifDIs2Q1IXom4mPdf+QbeRgbilmd0VKVF90e6fszfpqio873NqJafYa6TGTgCCI5
QQu93oN7dHtHM2hsIl+FaJ6sN/biO8wnPJnyalTp0dZ9jXgnaXuHqZq5O7opoAUO
AyRMSMqT23E3Alt4Q/e55GfrBO+7vsI6elgpTiwAxHU3Mdi5LSfdQKzfdcdhK2PG
4bNe+lHPyCz2cmnSAD5ERyOPgdpyr+7PKsC/kAgKZhX0+XNz0Ayb2hJDd90YOq1n
v23vjSz0AYbn9RunCd20hVD5a52E/ZDbwfjxpzDSG8XnIdL1ApLEHH/l+cgLZwGR
cs6M3B9CoUfMqK9PZiv8cKodZeMgsg54A9O5m37p1GHj4+NDWt3iYeGcQvQtTio+
cMYPR4lb1ngzo/nNn1bQSnl5vOi6PmcgB5iTr8xh/qrWhnHJY/CHYmiUw8LEdX6H
OpcKYa7lUodVSjBQgubVewm3htZmbCLPrDLZZoYeGdlk/Yyn7jMHCSuIXPCNM62b
3M2wIbl8Smjg+vChFaEphu85nKcrZeXpw2kVyhalZ6lSBxyFITeqtmeDs3NWGdfX
DLjFw0gIe8rew1B+9t9h7ETsVu19j3DvhiSC1IdNZJsjbYUFTRLyTgUdCSI3Czwj
A6OCnx6PsvAEUOanxxZG9v7IdirFJe7WeIsC7H1YRxs4fO8eeEPqxpHcWDZCGZPT
hmRd62UiogRBJZKeJjRkHA+ssem/SE8sWdqO6pokc98UxxLiJaxjzpDiaFrrpyBu
QNPa0wb/G5RiQ4mCTxV86j1/XV22cvnXMuW3Sqdl8EcLVJ7FbqsaUKnXb3XlbWn0
eGVMFuNOTn0UXNh1quTfKO/Ww14D6+JBLTY8NNcI7LJepH5dZ7qbapwzrgXfYjMV
ww2Gpm48rPezDnO46EtWEbXBgpQPunmXJbRaLl9WUbrAPGA8+EnLd7bJHPh0/44v
j61URU74hEDbEzO+THZR9O0DXTbOjPxqN1f+A94y14FTcpA9N2TzpYV1ETBUa/R1
8/QEsLMZ46Tb6lvEHnNpCmAXujx3GQsj2w4FLncr7/5eyMeR9ILYHXRae3YVy5uS
O/SYLmDL18usjZdAUP7Kw/Wv1cxS7s94biweV5rKz0H3Q4F9LJGKJnmIeiaNYCu1
qStaXAes+ylSz0wNG9bA5YbPCwkPPWb3U2iNjBNz+UHdmVOikeTahxsqUbz7JTqG
ycoOPIi+yibcTAw/hrgK/qfEJnFAdPUfSjCTuX+zv+tZKFPhC8ZIqRAutoKJhP4a
ikSPHMEa5S/XClzG5Kgn30oNu+QBl9ih6XNZ9TSFGMwrGdxJDRa2v7uC7zZRub0w
6AeysR5P5LEJsNdvsjRBNg3vFxcIKwYqXoExMX1wqwqvMg0ovU1bGbNZXh+5YfGO
/C8ogLDFfIufrcRFiZV5D8bfrtTYF21bBHru9GHp27pXri3Cunsu10DzatCeusqL
SIOvl6mqqn1+de+EIS/OeL2CfSlDg7JSrvNAUFwCpHceI++sS4Rz+tFY4Je/YdBl
JS3PJxo2H3GGO0a7akodd3Zd0Eend90OrV4zmauOw0Q/ONHBObZ4ja0BuK0YKed+
w7su4VzAkbH+GMkc9vjT6uABeO1wi3yDpL1nhv6aO7qFcayVSf6uRDDwv+2kAWEi
okZCRNBdWfdNEYpQL5kvw5DUk9T+BOokVXjN6+yR/e9yxaRLQrH8+0iCPPqruHXe
tjtxigvkJUXhkzxGWHFFPdFj1zBwBzgOfHMK+4ob6zFZpcqHTBzz2ofzNU1Q5470
njeva/YSbs+wtSVpftzLj9SnadzgjOpqQzGNZjnfiakfAcppfE3EYlyqIjy2tq0i
3r2qI8p35I4VPxnVT/sa+RCWn5sfH58Ve+KaNiWinzlf8FRTpBvHwKBpdkw37pq8
z4BrlQPPFRh/dahqlwkYDYHGVnIsd7nJf/o5LMi6949v2VZx53o0s/PshT6C56aQ
divGQlJ7tvr2d8ymk29d7+dIP6a+88YqSkHgrWwqdShq6kGyTMelPG7G7ADIqSl/
cC7BsJ/Dwx9iGbrBSIYUMuWJ8x8pwuq9RlhhhlIL+sMrc4ATsJVsQ/FR1x/TfGL9
qeGKWQjQUE/WjfDmXgf7hpPHlvSF3Ghf0zWKoPWTTFTbxoy6NhHgU3r4SRAMMnkX
dobi/CdoJrENU5Ymv0+3YdhfLH8AyPQtQhjP5h4ZSYVtfKuOANyWJ0kG4n62RJeo
Q9ncPFfXiexJUxnsHM9YBxNYv6TOVZgYMkZbAuArW3a/TvTU2DKmjWeJ228vXSzT
FZhj8RF8Bp+IUMCL8feir7S4pR1jK1/8EP/365X0D5Z82VAtXlTfCwxBSnXxjMuK
PHJ8UOruvlA55CbOv6VJIHB9L21jg5WYcTQZgB7Kim7RKYxS6x6YD18qG0HkZIpY
ggdORQOPDCAxbgzJuKhuuv0IRUYuS2C7vZ5z17JRAJXE72TSypwM6AeNveYwMZth
0tW/ThUXhKpTH4pemErPS2CosprPPxSNIpv10JNJA29e09CCgTnt8ypFnWUlgssM
c6g2JGK/JR+iV3nrwJQEEy4CcH4GgBHRP7/ixe17jEWY3G7Q1aBr2/dnY7ijB05G
f8JkbF7IvPaR5P5jya86b9cTTg2+Tqac6vyY0EPDoho6xWA8LaTOuBl8UqwCHIYG
En6AHLcS+BBFt98WHdBHNmye9L1yx+VdiKKA5rOz4OiXXwHpRpFPqOmfXZLz4JvU
OKLN6s1noP5LM3AR4vHq4Fk2N0pJ4ARFIsxJxfJtGODq/yyyHQ0XmOZjIvqEdgMG
yEVnbzjbHuAuz8oAY019ee1eSL+k7eYAytFmGSwPIiMbRzILqRa9twMuIAchy6DT
LI476qjf7qSdvfNyVrkoNdWEutPqWjRcgYrJUzfl1MJRrvk8LcEwMoRZw0gRnemy
mrUT+9NdL+/NnppQU76vyqUbkuMDbE4ZjjKtxOFKp4WRGz7yZYGjW7IYeRar1dpN
QxVGU28GFo77Vwhhw04JX05Q4OSHJLw+PmLFbsyuy+gSWBTUSQx4TZpFtPiGNSlQ
9v7GEEZkl1ZzmNfthRwgay2HV8D1t3yoj7O1ZlNqoTDtai87wCa87gNz81juI1bB
sutF9FqIOfBPZja+D3x19gi9yoyG37y91AEe82LQhDy0qxBaS1mm42BCkVYWeb9a
m7NUojd06DDpghX14J64y1aCDxr7Nz+pIOk6wfO7rir7u2EINv7BXZOPCg3YRybd
uQ0I29XS3j3/CsAEz4KKMiTR7xsuJjuvJ8TYFjo7JdB6Gg+gyJ+8I+CU0AmwT3vy
1iLAnuNz4rvhL7+Faag6Osyp8qonWDIsfLpUCosbnApHzWOyuMsfbCXJrUMN5dQY
cq8cAOVEMz57dfD6mud1Jccg2ul07FNKe381mFudZkGitPv/oDQMH6YVKqPj8fY6
aq6fxtJ1fmNQbtto/dmP92yZN6wKXl9cJdA1qZEpgulnlxS8qGBTSeiZrH1LSdh8
iQ+azWN3OHyoqEuAsi51Ds5RGgxYbFUV6UZq83hy/q7RQV8yVUQ6SG8jPEfc31d3
dAGh/Mw3KfEs6U486KuDcx07NcbOtL2JfO84Gi+qPnLg3cOc41QETnbbSVFuQN3Y
b76OBgKIbrcmoasiv8HIdkNjohwFD7evVhep7oL3sCQIe5K126JsE4ix35liVNyw
Rkf241PmtGdOPMfeAxI4awGUo/QkGYgWREseB4mojyopYMT2F3EBiS65NIqqzJUx
hMHPzP7HdIkxJucVgApbSYg6qHb3+kCVFSmtkEkmpWnE5PUs1ayYeDjsZMxhfA8T
4ciRzWw4Hwdzd3DvI9HPLYXO5EsyLdHD0IfGNIqAtH/wD/Xi5rmk0H9FVTTfWEB/
efpHZ6LlDU5/ZSQCGHnnDM3Sfb/KLIRZngQjAPWMGAI8rlkHjJc1DcK/62GMAsie
bYxhlYX4ltkxO4xyU4tG2oZhv/NRDioRERXFSoUfMClNzkIJ61lHmS2SQcQ/c32D
jtn/my6mDQ0G+zOSS1QGzrG+25KNZS3h9lj9QohjgtV8UOlytaEH8ioJywZ51oo6
XQ/aMelTUIPUEFM7tblzGKGREP3f/dpTcwaWerKVCBDjfygapbLQLrPWUZxO/q3E
1uVBWD4/sd7kTpMJk2PiqtRvFF9ExZd/s4PyXTEKaSbFizdfGRLmo5aRsu0cBTl8
A2Mq81Ords6RpWEl5Q/0emmIKhWjHFobrGb201iHyZPLBcEuVPc17a+KpO2fjEgp
4JUxO4XRXNxkgqaXEnC+yzpSsQrEVs/gUS/eW7xq8Y9ubZfBoNv4wrGNn3BmZcxG
J298n1PABTRjS2ZV9PQvkxjRxvc2lujfJszvbaSZhvJwvoaUFRAiIVeTQ0rs5guz
ozxtvvM77++OkblDEZlkYLaUrshIFYrMkT9ASfjJHfKldjI9obQGcoYNg3MG8mty
RJ5oa/9qm2q7okbdTLqbIe3LgtO6tRzOOzSOX5bzI7r+6CfrS91GRRgz+UH4ocZi
EU7uVFR5ATD1reOoBSmHqmOF2oQjea8vOLH/2UxpoW52vaJZN7YteGhq2VWA0f/R
/kSA6OCeAQ/8/HwLOC1M58G42JpTpQ1OnPh0Qty0gI677oaPGHMjHkC8T3t0pqIi
gOoLe4rv2dq501KUoDsHGHW3nJMU8j/c16Fva1ci2nEJGeHbWYkNN/5OwtmUo8Ks
hwUnqXCEwcnoAZ2GK0Ig6flkaf8QXXx4IqfGFJkLP0lEgk3sTy5Qonpnu+78dqvf
1J2IMCFt/SWeAGUACl5N74uB+GXbNgvoRrYdGYqSZ7dcsh8LxmiLh9UHC5TK5v70
GBZVBry+xXcliJxVEAhD7tDwfjVlSNNgOSnzDSMdd2WXT3Hz4m8uiVY8XlKpXQ0T
Ilvw/Ib1NJOMNislpZTLsVGz8bEgPUqDztY6MlOMt+zJV7QhDYau/e2x2WiDHOQ3
IW92bpBBWJbpJwPFxPa6O5FIJttyytLkyhNeTWz/Sc520rj+4ksx38NFmzh+RW8q
K6r/Cfys3XjOxr7P+14oJfU4TRI+xZjE9VF1+mV9nlZ/w+QQcl5II2qGhMifmnbY
4z7oH6Aq283uSq5bc5pbYYxGCk59beU9+6p7rRzmFh4AwxYRBamCmmh4Oj9lOUEX
tGilFtuikJfpwDvBZ43vKzZl7PmHMqXqmyYlO79+3Ond1jy0BRL2ZnH3KeaJcXxJ
DTJZf0BT6/xNF37vUY9MoomxOmKttNGtjki5XPbMaPEiTFdVPKWZAhFfnB9c71gx
C02Lm8kFTIn/f8fSNU6vNluHnkmx00jOSeiaBRxv62Tu1CkK1lWw+KWC5UkZMtfR
xlHBckjV2Y9gE1GZmtm9WemaTJcN0F7EgSW1mCAXIJjTuKQwCRcyuThe7ZB7obmO
qEG9qZDZL09+vuukHg5DU8QsMygoFAB7eC0k4riCTt/LQ9/QRctanXd7iD/CFFUu
xNGHAORT9REffss0sYodUq1YdV6WgsDAYtxTeNwq5uzQpb/2YuhXrbRef0SNrMlI
y1hdWcr7VcRR9I83SGSxgKNYkY6/pQlhZa8ViyslRImFrdzKZMyOt0yvUiT1YIN+
5R7eyuYuI/0VBkJCqbFQYlFu8I3TC4AWVScKT50TEAW/XQOuWzU+VrNXrRNpuOpb
ZYLdoax/tRkgCFu6PcQz8XIMMEec0Ev+u+xcW8TeKHSMq7IpqYe63Uyr3WKgZerh
O4g8ZmDOpsn5LdTdYBH/X0eTLzc23qZ5D8ax21Q1J4ReZSOzrQ6J5e0WIiTgGzpR
eI+Depxj+uv9X/70bT6pR8Q5dz79kCPMvNTYuEXI00pkZBSJihPpnHTvR0Yht/uj
i/hc0UL7GPpTsq+koWjMPpXRmYwPj6b5hMObQUk1RvexR4MInK40P3sXDib8vWMd
JQd2UATCnLGKaFf9CCvye2CnlRaZShPSnVk2r4WXsnp0x0OQotyJQclZmwJKltPW
7z4J0AeGm0G48gH0Pr3gIlMBOmyKQQLDLEj3weGCf16tQ/hVdfv/N+fxUCtJSe/G
OXibV2ijDxGo412Zrcw3TphiwiEpN9UIVl9mGPVDWRCaTp69FuUlX2Ej6FJ1IWW+
npZ8hKbk3vwtjZQVsuuj48QtlyoY3C8ROib5fi9KnfZakf/56BaW0GlGPIeReXf5
xnYWShuXJPks+856z6YcFkqAgH8XpPcQsousynC//4Wi5zhyvde2FZGi8C1oHXFO
ba7W64//fiAbzul/hzDqbgNyWunaDPaqXwP1Mgb2Ski6Opx+eJxv89Ar57uJ7EhJ
2DVkhSkm1Y5WefVyQMDfdvyGm6e8YieA/69OXHV2XPLUTc6z0YsyUwLfd4VLpMlC
TwLey8q8m4l2QRtIFRPnf6yOS+mrbSW7bKmDHdEdV0jz+uGtpyWtkd01SjidJ7J6
AKZNAWtN3Mx46mcDjk8gzsHg2BqYBFkHRXEILO2eFGKEECC5bDmRFmxCOoWkxF86
aqWxQ0JVBgT73F1hcIypoFzh1V6w1cWyU1OJruBBVoZg4y6nXKKMFkhO7ecDI+JG
D7payw62I/W9x7V9jsm9bjj//ISPZ28zBW3DtWuiclYVhmH7Z61ULM4Fq3vPFFLn
pHLPL+HL1rpEYLZ/qtMigDS442ytUBvCa8dszmdYr2e4kigRKyXiobgFPQtxvdG7
22M2I5y1O9SSoL1ff0vm2GIjAQEiXrj0aHFfD4N98VagxC5xxM+Iw0oKD2ndKwzL
3oPInx4cyqBKBSfWanjF79CIY44aMMBfzc11XjlXskOXXr86AP0V5FTCB6jIBPce
8UP7FZC8S6K6hipl3wvW5K3LS4qjs5RkwBSuzPnebPUu0jxb0D9Q9pu/S/5LA++0
/PzWs8VCEiUGZUXRPcbfniJ/+aBLhUa9xI3YuEGMm+Y2PD3dtoNHvB9Lt8cslydC
rW8pq3yWqbjMvPlPfpOCKYJVf6btdbFxkyFEUJlyIqMukhc+400cUUaTdke2FKyx
LP7caWPMsLs4AUPsLdT+hXz1aLrM/4FOy7/XJeLk3115JhqYdiDdKwdt7Dlz8Y6P
wNV4mA7rEOM4AyJTSY/dJvCdNbndLcRNMUw3krwhCfQ9ob0xLeVsUr9dZy1it/f/
c78YZDT6D7imZg3oHdb4aidkvv6UXTl/3c/PMwERG4bBmzCYvOXScUkGX3rbTIWC
JwduBY8IsnnTTG3yfXJqEzVWltC/kXkP+b+tdScmCopT1C7nKQcBvyp9dYL87q32
VQl624Pgqhj9iCxpaJ9qWCsTGHc9cXrPZGbU99peKcfyykBsP2u8K7J8SYiZf8PS
7RRlLYR1GeJAn95aG0ZyKj5Kk/9SsWcTM/Gw3CDcZ8W4v3/7TE/Pwzi9gyFFkDQ2
b/3lGizFV9DybOtivO85ckxFubocp91zrocmoAWsPxIR27Df9kz91mODpkKZUIaV
iGnqGHvl14zTVCfMv658tLZ+SFpPeFj9GpJUReJAdDvCOqSmB5Cc84/nFTMH2J9O
L1GwIpdcue31X9OIKBFDmj+4e2k3VWIzYh840XQ297R4LxWP2/jlm7L3633/rWm7
GNjXy+ZziWcNNPKPtYqWRyOghq8L4RNgCG19UpKtAustH5ojAVuAsN6Ors8K4k0b
KIV05hGibp9d2U00yej399iyUGuEiFbtJc2B0Xu5wt3rWBV0pCiEyZp9zzG7/WW/
/2qO+i/L6rSEWZKiW9QuiVz24/+MH0oDRMGCyYDl6CowL1Rkuuyi/03gqVszpK6w
TjxgZOpzx+95B/mdVPqs58klFThNQ3rDcej+Pabe1FaT8Dmtg1/zdLYC5ncxB0VB
dsWuppwWqyZjAzVJ3elUL283T8rFIz/R9Lru314eibOsf5XdpUnurykfaziDz+HH
ABUl5PIhOREoFE+JxPqE1uDKOE5qvicXzFuVrTPeQhAY+bWzGWtTsEmnk+BPVFZV
L5pb+ODLEdDKq3ywWqtju7Jhdb8dIwsaVpIH35md/B4GMYc8CbiSMGFk4EuaeTax
nLcbO52X1ez2zmGCWbsOgnR5CSrh5O86RXfXmmq07GtpaAdDjrY7qP7P2AG0DN2b
qwfyHklBD3ehcookao7+Wp5Un9dNisN0kz7Xl+BmXw9s363FRAS59e3Dkp2wIPOI
Dw+WRzNd6fA8VAfjQHkZwDs2xnZuet/lnQMz/x/IjCtQsgzKNG5e812J+QE0bcen
xB5GZC11qNf7dfqiksIbNqZVNne0IQ9kki0+Myj5szHbyCe6JUTARrtYutYheA+U
rwbUcz5KPXfPLmebxbcSo1HdfXtKjDHiTnGlzNaK7LuXzadQVOtgjPBp7+Y1h3u1
0f6tagEu2F0fEPVyyZCSF7gc+qyQH1es1L7klHUPIVkC+xrSiF/vDm+n1LrgQCDa
DqssZ/IfbBp8A4+yhlE6fpgZZvN9L9lGW988ZWrYIp2kAD9apa7nxo8VatZddZjP
qB6E5OnCMebqAxDmJ2dE3t5wKBdnTicYC3eGt4Ul1pogtxB96sHVYyZU+ZdbQ50q
yVmNvNY0JL6Yj0KtOlh2enTL7BAqO3/U1OXyWK4NQKcjkgFf3xtuqWl01nMwtWBZ
RFNJtnLUD8vpQ2kzd7UwvNSSRLMygcLcbiOampfuka1UM2IhEZyj00SZ0uQ7Sltz
vtHet8MyVmzdU+scZJEXjm6LXpem4mP4ES+0l/6rgBC8xaUg4SR5ssxHvRarCuxl
vud8VybbpfpmqxwHwix5zKPwC4GSgiwNfcntTZJj22GCtecFUyhdH3aPXOGAAd32
NZ8ib8LGnCspdhS9KMEFNs2nKGVrEHURPoHPCy3ATNecP1Zp3F+fmg+27dmhJH1h
V3G0AVHAQ0Nw7FMrnA9fJqo0jH00ncOhZSt/VqLrvHzjiLuByaCxPwio9T4r8V0f
Pc4HTnXYMed8hvWzsgI1N7VYMSmtVJn6cGDJGWOhwk2QvU+a9mMa1iIc3qASiS6v
z2BO2SimwGFniRviMzoj8BGqtdfL1upRqCfZ/7MYhZfsW4fu0ik9awNLaaQKY3mk
LU/2vLcT+4weVOHfz2zE9xaFsZ1cq82JDENK8PZtGIxP4XFDRIE88AqZ0hDjbjGZ
L0e4d5XvLvLBBtI82M1Ec37ua9jmvjJO94+/FC953vMRC6p6dx6MjdktmqKW7P/6
4oOQEKM2JRfrT+D7l4o1vgT4UjBOsc+zWM5ae9tHp9n6wNwiUyGUqezOjauOubev
ZMXz42ZWxmFSaV8CbucMD5Wb4waOqtA+n8vB1Q5zn4Lxja4I3KVnJlkbVf3JbMhZ
Q8d4+Y+wN8YjuJ3kEaA/RZ/MlFtyps5A6dWTFQXkiGzO9lmrPi1h/H9WeUS8a2CF
5LC8onkDP17OZgIR4r5wgnkJh1nKByDWpiud/0fyfaxQvJhwMM0cxGBNhta8nSwx
vvbdy51zLyB9FcsWOUYNA7q9TPiwnEc/plk0f1DBmBsvS62rZ5JllG8VEtEeW+ru
l0MhLW3Iz4VJwO9oboCVdWSVOsGJG1PJ3Og//9D/HQh+AdP0hky9Tc0VoHFbtY7v
ud0B+w+UqC+4Sual7EsA52hu4hdBFiGc844KeOD3v+fQBfLJzj38KwGMrQpk2JK2
v7nGW0zcGSREP5wJZmgWPpo/Wbi01YcGsSvu9qdyOnpFhcnCxZvlnR+11C1VybhM
O0DGir/uCRVrIl9/D/AR3zXUGE8ielGjhu3RTCq63t+HCkLqaxGxBEQd+r0A9/rV
E61HaZJzvB0GWACwlRAQfEfvJyInMNWR/Pju9Cao6FGOt8OJ9KYjv1FJudfmJNAG
2kNoi0rGl6XmZBD4WixkytRwOQhkwKI1uRL03LnOXKFOiXsFzxOZaavCkfHZkDzF
gLjz7PzMK7qSFvVRgPqoAH/y2OIuqCPK78sQP89okIOUkANnAe9UAgvUNFPjkryr
3B74MJcuNogmMuMhp3GCxwS80YEN4WQx8ylYv92qhaz+Pnq3bIyB5fGsj4NppVGt
FXgiIoanfObqm9xLpcVUshrVPisBVkFFmxfUTV4TfDE46nAQg1UhYeAS6ZCUA99F
jE/7JriusivMvz5LByDo64xeW5t9QC+xkCLAyGxesxR7s9S7P2JPq0pLmB17U11O
Be8+CxjUl9vkcTM/P9mu3BvVL6jerMHsCtMHfkAuScVS/MofjFxxOO9ylNdvS3vW
pMXtHxSuA1Q0nyfeAq1jfXVm66ubWy5nRv1KhlLl8+aQvnLOFjEmvyUbSN8MpBt7
FmKO2Ohtij56fyH+lcBC49/ASEUTgi8Oym30UBkEWUl+5g4x0o5PwB/UUfbgaQiJ
iMBiAY6WIBtqYIgGgDgt/7hJx+8XB7vZ8yweddQt+56r7pJoFnHEb+XBOHxWSJ7s
duUec/qx77dfJUwoCi0RiHP3c0cd8pAfc2/QoNqUaIXl7v7iyCy7iKe3QLBdicWQ
2GUt/EyRYq8TI2oHL9drTRhs793N/ptMAheirJYyB59lh3fnvEtuaSMfd3zq6FhK
DrrJk+zl/mQEEaPueYYwAX7tpV3tFmgzuJXDtenXqGxBO6NnemCxXyH8612HMPIx
Etb+aMGREgAjmvZejLvGYI4KUOfu9PL2MIAXwVTyunJmi3Uh3Tjy+qkaYirrG10N
IisHVo3qGqAVCTPLL2vGHUyVg0DN1fLz/E8dQI12zqVKxAgnnxIHHoXQfWOhNRjY
eYrkv2899MQEKeIvQ3vG+z5qKsbEXR6Qfz6yBmRQc9pf1K9llU0Y86UIbXS4zIk1
MRzWAWXRDtHPzarM2JrvHjyM/qJvOOVOnozLGGoMxmRMOuq4xO9sLzw4D5iP6Xqm
W92U4RTUDVMtuNSYGEmlcoL9jwFjFusnBBl3H5FvsXTNeeYEu4CWp8O1o9KmKCwC
WF01wZw4Hk285ZF+Bnk61oMZuCtGRb1zWRvqH6cv4VeLBxb8eV0riJPmrDG8oHRP
lZnoDSmPVrx+bZysXMGOR0AvISiZ31C6gZnt1h2OPitd6VY5HQ595KFXeLXqoO3C
l2gnp5c7bPyOD23iU25KNk/+ZKHzsxSzy6QgB7duIokDWReC4EoVAPOVREOXpD7W
AF4dLw8YsiR51Q4IPzqQ61xZn+fQ18dqdhQWKBSPNUKH6rcjQwofVLrYJeiNOY41
zckZJr2mcUmGvTckNKPdzZ1W/W5s1OKIppvmznPrA53qmHILbAVX+W+azNGwmcaL
fcbqeDhLu+i5VC7f8BVPS4ED6ACRpgmylAabokyOvj9lyApJB54OKqX7RjtDzKJ7
cSwF6izMgB8PV8uTPaP/FqCYfRuyFOeJvku/PkCopsJl/9tz6/mxfVDG7gXPkv28
vedCACSW4lZ1I1iNXbqLHjvXHrteJyXpmCqO0Om4TLXqyOWghmGI4+nfvr5Ynhex
8XvV+cifrkLuiHggiZ7pMLDhwWRcUE8+Fiyn+d6gatqdQTythU+OT47ddje8ze12
EmjmSjqfwGgsjoG5jzsakWtNFeIdO7AQhZRJWS7AQ3cOJeAWh7LJnsNmyugCJmVh
srZkjXeU0rd94GaG7I2NtRjchl96wjLTt+EFYlS+WQasHQpgcCnHNNt+rmrQRD5Z
Of1I7eIwc7P5FSq69A3xOjVYJNDci673QvjoK5O6y/iWO3YAjTFStsImXtjXPgUo
536eC+3X70L3Ga8qf81jldbMzdsnI+o8AdJcwXx311az+r5TmE/Fy5/62YWCcB7l
p1IHaC9n0TMXYyu84aETlzV3O30pOMz8rGeOT8I7S+0vfHtr46m6aSrbYOlZmivP
dc6PCU9Ao1btujng81ENA+KiHChu+20WnG9IL/Wb4OI8VQLzG/EDRKdVrmlR7MsL
jMDlBTkmfy+COCT7oBQ0JZdLlty1gXRgq791Fram9nzL6YqEqq296UU2ZZnIxzeN
b+tb0YDiUg5KEhI0xOmXfUEz9+McW17bPJSx/4l5uGBAA7Wkbh/ANEGAcEESGVtY
0re562aVdZpMUO/sEF3fkWVgwfsVnLXTsExrcRABUAkhtFk4npF2BRL1vm+l2RKV
yVfEuEzVC9/wI8BCypm4xwCguMeLBK8Bk3ahmCk7hGCWS6GZWznrdrlWEv57VF62
HyoMfXxpRnUsw6WxWkQ0kazhhSViV4u1M/p6tOsAfs4z2E+yCVGy34xcOoHUmwjC
TeUQXbT1WS8Qre88Dj9e0ZKr6H6o1HO77k9OyylTMGWmgdw6KiRVnqM7MKdjcEfL
eBKSl2J7USM8aSUo+RFvcwJt513pwyNHFM8rPtTx0d/oKjmp8HLKKi0B6HeOXmcP
0B/QXfm28DDop5uBFeF49JkzPP+pvYArspAXMDkzdYJSbPp/NpT3HJxEcSyOZ2dd
dclqx/tV+KCICnQwDizu2tY1sjxm4pjxODKFT6vCgLbJLX5BYv6conKpcMYOt9pd
sHnVJiRXeYleN3LcxGOYUxQdLc0OVLvKigLVpRUKz5A7EHYcUiBahaQuR9ooG4CQ
EGQ61gTtCH+LEqI19+7SOUtvpbpovGcmnNfapkqQwezaCui/Le2W98NVVGZc+X6g
rku2FDTxvN/nmMCQVK3mAmaTWrj1pUTqrCpWel+l8cBigZyI+45fIHgpbU3/AUbB
b+cmVgWwWKYkif56ZfFTXYBRsQN75DWirvwpO3nmjdhLPRAf1m2+oCLEUHkFEURz
fWxyjt03rEjAgHNKab0avjLQJOtlR7OZx7Q/LuaOa4YkviNGRZwSjOmOmTi0LUS5
OtHmXe9jdx35AuYb2LMi4aRaqDW7ig5ID4o4hgnhf/vxZ3OcUS7jLV0UekukvXI1
Aj3RPAGKfCqAiVUi09FJUoZQkT2oefA+u+vQnYqsjzc20L6GLjr1eIQco9Sy1HJj
NRdUk0OBZ8wWOmFvJGp/cwKbyH6EmtDMni/VyxSOeuJr1uFjUz00uHGOXQF5nV0I
I4o+VJBzprKqi4+n0ncj6VUwRJjLT1Y5sfL+oEpZjdD05dyiIZTO/A781p7NAq1I
nh4l8vd4A9PUo3k47M2SYJrl0Dw0o0bsZJCse2xHP7/xkBYAInxheQBJXo6I8leo
e1Y0tCPToVLJdKmca6fOT9UXBdOZoTJMx2tiJ1mbPvDicahizIsq5v/XNVKnasA4
bu+XeHa+sqLZYJwawlSB1L1PQRVjjPW30DdxXlYEybCC1ffWFuzdHNKsd3tfqRqn
mSX7w6Gez2Pw8PR53akyNoOIrkfMlg/tNMUFIEg+UCaxzgi+rbOcRn0v45/frj+k
33KAWglA129adDU6T/dF/YKtaqeZBfY6jccuin6HUmDzsZKvi1COmQMYn8UoE45b
z90NoQEgka5g1XPoOVuSwBEAcSU1JNOsX5cjHq7qB8uktFkQykFnsn0z6vnBBQVT
DCC5g1XK5DAkFf1rJ2Xjr+Fbu+++tEmJEEUQeZgVUg9vW8uLs295xGhGJAEl30IK
rNWyDBlIrP3PiD0rhjm99VaNFT3C0G3JpfGNradlEvWGZX0QiLe853Avs5KX7PPd
EmC8cOBFJ/0RAcgrF3uk9ltHMeAFgGEVFbeQW5Dc4SBCAhtA97iVT0saKe+jjXrI
BA+IoSximjMGWgbmSmBVwIeiH6oKqzn8JXAZAyJFIZDa8IRh5eH1FrNp6jea48tB
H51WQ1rHr6s8p9jzaVcHedzJ/HZ8Xuy6RHb6DbVe9dEIukcMwPdcMDmK99/i5CN+
Sao1pUffcQDvDMY6joqOTsOonTgasjPIl1/lG3giLvcLfYTyPh9AMUx3aY5oDs3K
cT5lLRpPjYaeHN7uSjWOj9grq0IWSWcQgFcUpr1sOwo50+sApqKJCMAvpzaxairm
ir+xoxAK3CFZmPXEOlSV1+Wi5p8B3RFSZrv7HQQrL/lAx6ZMb3Vpic7vqRuFi5HI
qzC11uEWzxMpRHL4vPNROoTTXmrW0Lv8Wnpvrzf+HTuBttYvWMnuOrofVQibr4Cx
6uhByCJyupaeFowavcdwm3VYDf8GHculcEWWoPmVVKSkJAB9lU/bdqLam/k5tqyR
6cIilpDytQRuYb93HgQxJP+kMRguHjB8tOVYYUis85QgoQQFJDpSuqNV6VG8pYCO
sTj0Y4nuuzaNrNq2oq1NDGbQKepBTOwowybqolelXNf/FHz/oMOg+f8jsYwN+s+g
7alRaG/N4LWqeV+deyfmXl1mDA+wbq+vBOTJXGCiCm99nrTcbFlyPwM9bKK4ay3y
yZ0zVZm6uTnZOtnMgB2tJwdMlJ8xboYN/ZoRMrWrSBwy0QtPXNWjz8s8LFDIQWhh
zAh2RzLWKwS+6KXpK8J44Sl8l+Gorkqp/Z8zhJsIyaE0jRt5Byc5k26p03o/YPhc
2STZrfvalfzMcuWSKriM611wlvQ78WTweM53BxXRzd3A8eUCAVrYwq2z4eUlDjoB
jquQ13CZQNHbQhIr8GU6Jv2xrcLnEo43fLVvfvikpd+77h/EuaC/2tRU8ebWMRES
Yop99J+n19HS9VaO/o7f8ufHCYWLXUCItaugA+ZrH9+4sv/7awMNmUSrOAlLexBB
n5Bv/5UCBN3+J7vqZrSN8YNkdLhS2Uw6LDinjsrGYVQ/6MXstljQv+ikiNiPqxZI
eiH3kQklj2BWnpfK8DmE82VW5lbdsMHWDdT+OLGd5CWhtX6D1zWaRGkkXnsheI7n
N07E4jp9azcYotsbpM8Nc4iWG2VNeAs8GQRCKGBrTUWz9iEC3HF6VGRoJFmsaIn5
GocZ4b0Rh9nq4COUHTPG+z5/avsU9XbLdMXsJpttSiDWgQ6KLhNkcFxGXrK1NjPR
ETmDYb14phIvGkUFLkM8GGdYK4a/djvJXZfi61qTLiEMv244g6CqD023SL2NgDNB
g1ZS/pFYfdqlo7bXiDuccAs6/WCvWdiHF+/rpGfh9CgJty/YIE9YWrQbtsKmW2eJ
T9qc43Bg1sF55vSE4NeWeSofCFOaBm2qBDq5rZfCgUHWD8ZNF8NbsTnzRtXik6G5
ICClMDUzZushg8SSLFguzfdxZIQUy1QbuBFM3rMN2+6jnMdZ7z6gyLJSEyEP8A+8
kNdyb/aPlx3c2mEBX68WERLQEclQyD7QVOf4As4mMAdcc4tKeT6ZwnTepRcjNJMy
D7aTRdeQv14b+b72vrYsSZiGx0BwOBV0j9aRzTUqTc2NPSC/iyy6/KWokC42hojQ
6IulZjnYX1k9CdBjViZVhBOaF6FAb7LB8LhJp939sqkAQ7d2E/VUc4uY3j22DZ/g
qIIPNkZeEnhrBhEAk0gH42+F1xVoxvrEMpz6ncSahlJ0fgetzUIR/2u44bSI95k8
o+XImuAkzytZM/UPSAsdSo0RbayYMXZsTmUsdaXb7rDIRRN8mZpqvKonJmArr3Gr
ybD8yb+yh5F84k2gC0R3rLP6BD7cLnRNK2JNSkfdT/RAJv6kLFJx7Lx3RF0V+t/O
KZ+IpRyi+iUPqgxXY+5KhRqw8yidVsxIKSEynzhkBiJYWo2EMz9Jo+0YKvf0WeOs
r96UPWIkb6ssSzjEdx381I2xv02TjJFgAfHUznYiBLw99SuWMX+ex6grTV31MfHN
EXRcQbQWaqDggtX9gfFPkVx6yHUYG8s9Wd1thdbsKNHpkUby9TH8pJpKCqpwXIEL
YHBeefkeybsAl8nrvJAVNlS1E4dK2ydnznlYj5RGga8V1lx6Zdl1VMR/qXvqpGgA
diQsXsofAJz4S0r7SUpXs45UbsfQhaSoLeAX1UYxcgUTuk1VW9l9JsIdQOJ9UKeb
ktF80wXij0jAGcDVojHQ8xXzLmjOciOOaDdZceV6tDEp128CRpgUgXsM/8RRc/vm
IgnGYzi6h0Zqn0bTv+hZMjnvYggYAgwmzkhGVYQMtWKPrOdFbOOAt0/4XPPAiuFA
TykDpNkdEcx866eUFjWa6FVnqFNQaJor5C25ryOY8bn+MkHfr50Bf1fEEPP4NLTI
+JmmbXoIbSH+IVoarkMkOvFBWheSkpXsGIS2MrTIrSQdwiMLWBkYcI/hFfasOGgm
QOl9VNPtVgsvPA7mU8doNWFyfPCTksIbI6nBVe6lRB34fg8JRTpilM0K1MFlOM/E
tI7lwTQSPGhJQdv4gB7YQcRLavmCGPwz5N3jjJ6cMA+meV4wvQzMK8LYhMWhbARu
bXwhp8N1ee3YY0340XCiH1ItQ7nI7qYPETeoLy5TxQ/Nfo6r3K/uubRI67WN7R0H
0Ls/yya+c+OgVKzuT+8q3HKEvYJ4xCHu/ru2Uw5ARBEpGZO1mQp51p7Ed/HFCp6g
QVfCJCm95HRUaZ9seLyuf8yesl4Xu1QEaagTVEGgd9AJZtCVQuLSok92vHRtAb+Z
z2sdItsPO1rWSKp90B9Yb5lH0ckkwsm6aLsumCowvOHRjn2atm7DkjC+rg8Ch52s
skhgcsxfRLQ1OUb/Pn4envl2eqkLszkv9tcKD0avY8Vo510dOkl8VHvHGqfQhuB3
oIy1i0ybDlzk/3clJ4/ym6giDsEsFdoSc8vil27zQ8hpmQ21jxlpRwJ98hpWwvps
0Y5VXjvhQUlQ00aWS2V3rHRwPH+4vglBtwHYu1RSdL1hXxMX83FlSoZdzXLkCjs7
ln15FtCg3oKSuIwqGWOISQDqxnMmsZjqLQjp+JysXhKOBO/UfjZ/YeW/Q/Rpr1NH
AHvlPO/rcFjDUMdZuQ8gXPr/6Yi4JJ78WRv+6W8+2mVx/hZ7C8AV/H0p5Uxv9cAJ
gfa9a7/jSne79YuCZpzGrnVDR0ReLr/xhY44+OEEcqQIR2kz+Uc6lmE6+MWFw6Qt
22Mh046Hyq1CUJuMJDQgbg5+jGqSHpeDNvoIJNJIUHDGX124qn8lytjNTpcVuklt
AnPQOzc4aw/x+9E/w+xoWcfVf4vR7H2m5OtD8YcfjgayrnUOJuprldycob+7wRrC
c1+iu3Ulk1RNnXLdOD9wO6ZxuNQ3dtZtgFBviLCLb5g9EmtykVBUvHsvweOhhP4J
3/MZuFZyoxn68Y0BHYLC7d87SLBMyDtLCRZ2SmjoEdOrCghtv6uPL72GVj+JEgd0
cq69JIyJC9dA0GRPZ+Amw/SW5GY7PtQYkFh/VVDw/rzhDIo0oo41Sb/rKHeVW4Jn
Fn6okA2/aP7H/Q7l/PIEVEYg6mFk1zcpZ+Hq4atW3gv/DqtGkFNWm98FLusdDehV
auVZkqixLD+k7Dk9zz6AhHYjzhwH2mYc4m9iF+TBNhL5HEaeKgVp5BSZQBdUVN2d
HEQ6wkSmC9q2Adn0Fp4sLEl7XuOl/6eGUUevdoj34cNbFpA8k09Ojam43mdrTa1V
ufSDPlkcrK9D08Xh+kQmtIS1btZu7MWbRnXo5CRJJi2JIUyIOWRHr+UMIwo81qw6
Alb1Tp+sK0Q3goiR+vPBeDiWDfBpVom8NZvamZBUPDV+X1iycUwIYCj1s8m+Eu0x
QmrYu7JURVafF6iWnKUtwFHkV4M2oMzh6vRG2m54qo7A/Ra2/cJDbIemuU0puI5l
NWBIHPvA4/+7KzyQEv8ZuMDRGwTiMBYJLylLcOD2HTssx9U2tGyDTblXFmfogVlr
qa+OU0I3cuUGADaNeTpZkDWVLhziUYbUFUywSCeCYU5QSjEEMqk5P3pCQsHLPReg
I4JsAe0XLByjRh5S/ZzsEO1QjGggq2eOk6H2ZVVoMHDbZunBN2N8Tiud72z1lZ03
rlop0E/IPQCK94KxYNRRuFe963PAvSWe0zrsNFvIl3XFaD0fmSMRWRdLZyEaBze6
0iF7WkdCIeEhMnknURJUFfE4XQDoK10tRNf6NlT/qriCkfRbYfTjiom4UwDlCjmZ
gt1qur9duNjdAtE7cbixuP6/nk7RfxhXGdof4nSgoBcVzr/GG8WU8flng9EYeqRT
XRSC+WqKJfiHNdnch1tU3fD90bobl0dYGAhmR67y4vZMCAqZybT2QsTxesUXG9qm
4dofxZudUyKc9nT60sVWk0u+t8bur2qTR1IJXXrbA4UjdlGU3vrbZvle29X68XMk
IoYfqCAu2uhCHyPrXj1zS3jO5jm6xtIcuCfxv1gd1Iw8t6pPQaQJX7do370sSwrp
CpKfT/uxXEFLZ5pAA2RynKCJfNr6+1gegpnNOfJCGedFomY8M3hSXatmo9RIYql6
HdExZ27cloG//gm/ZFoAQsQZk+SNNqDtAJw8ln+BuyiNvH/ezjnlE+O2NNHMASeL
PLFZNwViWi2yHeSiSKJY52zBwOml+y7r2SI03Un2+Ozj8IrN2/dZBjbLH+c2llTw
Q1IOIufoUUU1xDotnRxRqK1Wm+PNx3n35V+INRtlceApZDDvLxRDM7B8+fbXVjxu
g3u2SJ7XSB6n+qPK5g4t4mTfJB+ooi0SPosN+d3H08EKFCQh07fCbVOEDlKZZ76W
zsmG2Z7AHzET8DpddwrwwGBr6i60EX07WhYP/mnAmZOqSB2li7+iUwarUZ13emK6
JYYxmWEM9W9JvpT5R/xkKcGUHp8GTyj743S/yBQ3a5G2GMlcXonmeilfY05ISpku
LljcxvgQfhLxO5Cqab1bPFmNVUJhL/V6L27Byl6ntBAOPfCcerzhKqfEsLoF3PyP
cN2PiJEaAV0R6+N+ecsJkebJYpezkxKsDpA3FneEM5WfwWChv6Q3Nhea5i17j3Zq
TnscgivFWVHg4c8JElAjLIJewD5FakuXbpd2VxaGCJVpCNfBUYE7G5jbQ+AFoDKT
auH4CzRiwKEU7cs6BNY3vthLwPrbCK9bGzEijgCe/uXxhFUoySIO/K4s0SHTTn4q
LH65zoPjOH1ikRy2yeDxPH/Rh5W4nzdHlXSJMxVtuK9+/Cx34JXn/mgsRrqspm8A
W5IqXMgNQ8c5QKK02hmVJmu0dudZLFuUm2BoCmiHtIBEyNJFM/xeIidO7hhseG8/
qZZaRno2xUDhRs4PIGq5J+JRFmGfT9RLz2BJXPGX2A7/kGXHr2NUiWJxQxm3q0Ee
nIh7TDS1Dryr7+Eg7sDofPwpDWuV0M7ylJXimHQUeRDtaDG2Vb+o/h04op64Fe/9
calABfoWFB81E8/0j0fLpNzsONRlFUf9ZclyXebYacjErjVh1khuly10MLo/MFj6
FVfeljfMaQ0VybhNyLI1e2blwBTI3P735sAlMlzthq5rT27JTYSROA5ju/+NxkAT
CeAKGVihN9bsX4GO03HegVQ0buSGfGXgBzXTV+1mzHUTpQVLeSgxVAxbJwn1Cecv
NVnvYalNuvsE63489N+kZvCoY0hkpwjdhfloSVzjZNI+m1oEXygEdtfxlL1hsnql
BBWRRc8Xzdkegpc9SaCcyudgfTdgB+DfI0LDmTQn/zTthc2SHa7DgHfIhrnhAq2v
e9uEmg1iG8G4D6Bjw9OKW7+Ey26g8k4QkuLfwlLGX+51ZEzgm6G/TRGfmwEusMfV
JreSRx2CAgAKYQb1K0DBnqgxztWLqh9H6EkTl5OCxcZ7gu3R5+e5nK8zHT/4L2Ir
pwCHlHs433O/yQw13NNSxKDYw3AijpPWH3S1qYITx6Sw4ihBNunbtmjaWan/Br3f
zzOBLXtz5erewrtS5tzmAspEFwaIhJmgkZiCMTkE2C/bLlKvSfdS7qW3GRFoXCJR
/U60Pnf3umdj9ASMkkdSy3/owDScL+Ae+zQww8djSQ3xF7DAu6V7LTeYMjNrSIpn
sPjrLN9n1gF78OmFGTdoWBO7J90r8ymT2+OBhzUjj/+K0nOnaLpJvV3vjB9Hnhp/
caHscAzeC816j2zuryRygP04beGNXg7ngDUvaApb8GRmLdJUZLB5L3Aj27yXJ/Sa
E35pmvGBzdblrkYehT/HJdbyVv9D2np+n9TtSXBe3Ql7HoWdDs/r8UWky6+nD0wd
eMIbsFFHrdz+618mP0wBJ79C7Iw89oMh9fJWflM5hUquUrjYwlqVRpaTrjJnhRP9
x2KkgKT2ayrsgwjfm/9M+Mdt9s8sUC50o7XXaENZ7goNSetmO9C7txtW41KgBvk9
gTegQy5FaqYvd3JUGEiRt2FzYGe44FFJFUKSCiX08aXdFTFA72Oz4tSXm7Ld7u/P
tStnZPi0JeQlpWTuNPlFlgj2Eb2jiA/svwOjfb44AeRD1/qj1AL3YtZr74bv0Wq1
2ZjVHnNy/BdCig9aaA/hMgyeN6TlHO8tfGcPi3QS17ufmigBeaJTiI/tl7QR5uTg
ZYd1mgjSsUY0ORI4aZHXF0jm8J729Jz1qbQDXOcYod/GNSfTylyKtsFl1spZ97Lp
GOOMWBbd4wO0xzwy0xS53vpLW7sBytcU1OZqTAxszzE+Pb4Lj6PtdPyJsWcpLsmz
DhbWrMWyIP9LDhwsM5NBryHsIvXAcsI/G+zgCLEtBHFbkYyuUgVweo3K3Jbk2aw2
EmJFdO2VhJYofWlHLa4a/nO4cZuwcQkKuJoSGQ+eCzIyScXstEzuG7dnWJ7q3Dbl
NumlH2gmHNWd2KAAoTBaP9oVqZicR8T1FM5A7WjZs4rB6qk28VGIbA71KAZawM74
I3Jcu3t8BOk0ntWN7L39wlxGx8GS7QUe5pGCD006Vc5R7qJRcSsqrr16TdX0DSG2
8pfd3yQHTrLPYLACd2wpq1qWhLKI/XEm5qxeyvTzF3XqzwUkZTveZm5Yx68hRu3y
QJg+PugX2OMD1pIjPzlfhfsgIvk7MQZ1ENkhE+jnXAxokmfV3YzdMPTrLim+8VZH
jtGba7q8ghzL9+QgEptYBDQEtw0qYxSa+98mck09QHRyLmEScX4e7DKXH45wGQDV
ddJHCfUFgZfLi1B963q8gZd54llKGYRd3bCVSkDMPLajB2siGNAdlTe/Rlpj31E7
jwmWmoKRtjNMfVLOTeh5/6BdDsJT9oW8v/fynWAWpBzbTC3aBnOVpG1p8BezaxSz
aWJFlR3QKqAMg5VrOvbr8g/P7vSTAqdlMC36pBLC3wxvdJhiYOXFWzVQDCLZV/lK
eXu4mFKfb3AC2bqfr1vjDiugczGnNB/gCJDE4Y66rjYQVQ99gMbNNaeca63bmnXZ
MFm5SJqQRkBP4mOtbqzg/Z20QeQPGn7gsFZZZ7jfGGoHuwNOjLkp9eTAPrpjAVFQ
O0yE0G9EXhbrBBinVe+TNx9A/yNNRXSjWPlISA0z8BnzJW5Ueplr7DZbUEhF+zQ7
NZpB3nUELqXgQ4auPIKoX/zOr2Ml6hGwlQQnngHzEBHhCGGiRYXAa9AebRxEjlwq
m9dBfwkfEzncL/102YMSuPHkBiPeveQuaOLHuuG1gyAGnSrk36Hp8OWZ+be/LWdg
U6t/keuusitRRhaNdACQ/V1HoyJL2YT4Xtu8BUODGoiVRnrP9aN2D7XdTTvMMsfE
dHLiHZMjzvFQ4orh0xqW5jl2vYVBDyNgbBgd8PL6tnJUninxAGItWDjVD2zm83Sg
uypHfSZGugE8rwpOA+pj1C3CN/b+NWymECcAeYRIP4z0xxpGt1x8Tn284jwn/jZa
FdKZF9D9taX8XxHdSKMLL7dvEgcpTtf/+ILE7hnpT+6Ftx8rGWp4S8Gti2OWvduw
gYd5rPCpf12qopYJj6TmYPLcz5qZlZzudFAKa404EIqOexVK0DZUOCnfFqrn9xIs
Pp3nklnCCXbVT6KRsJUmiIVkztfnavV8m7MFy4d1q7aDzK4NSNzk4dKLiMfC82hO
tbXPWuHcFsK6XW1wqdzog/pOOkTAMgcJWKEyxOZGJe1KpedY/mbVgpKK23bkph9S
KwbyiCGo4pYoCeuAyEWiJt/T+hsDszuIdiC1VLJZpTskSr4Kjv4sSdGP14kBObdd
mw/L2Ai9qwDsRyDYIpn5P41hqKauS4XXlJ5aupjAi78aN7zgx5SsbuZPhPr7U5pE
WC50Cs2xP/GdKitvaQHVfusGEhXiN0MtYabdWYF1ACDghHKMabn/roQJyd1mlsz8
wnRyE6ZjCWTgBeu6MPleMnxdxFtenyk4TzHN1hkJFt4X/sLvJ7MLtoyH4h7wjS2Z
6T8G0v95hucWZ5S5S8T5LiAdHnsVssORAlxkyEKHsaRnd8/2XuaJcXkP4EK2tr3+
biIBVpwXhvb+b5F67Kuf6w6/TCGOvghkcEcpIC97c84GMAATEdbFFYymLJRM+iSu
L+zTyaf+jNb2i4FZSpZC0cfI/hGQgG0MCgw6nBP4Pfw+8+jaTC84h6hsTzHPDaXM
1o8Gy5KAgfhkNi2KdGwC5OeEyRCk/0qPVexV42L/zEIDRtUOAYCbs0wGvhDTLDOR
HabrFZJhOZuaO0gKstiQRZivKQa+k20z6PSppI7C1Omp9XFtjrHcR/WRWp83T1XK
4PzbMUSQ8g79WKHpLhYOmMq4SHcYTK387X9+HK8IEYQ6XVNXln3HsFchNzNgBa07
t0CKxLuwtAhn4UsmOcrQqClizFyC0h5TL262pdHcGmpYw79UEuIuD6IC20T0bHVt
hWWVjpj6CwMdiv4HY08imwzIh3WtJzderNjdZKOMDq8yuBmmrTxwSYLwwk7pgIps
dceD0/RXzdLjy89aC1sT1fIyndTsuQu5ohy4XkEh3i7nMOtkkWrpii6ElPKJChse
zxg2kK4YdM+mzrSYnHAT7Fs78iWVTxb3F1WDuF62aAhSf7wX202/U02fv4lWHL80
DIwBTPHY0Z3k+nR8UDOBcV39mtvMyVFI5oQRtgxnFfpItOI47vbHW+bn2bPH6cqA
/w/EkFUs3mFd7hQMSEnWyp79jhzBznzuxHQkvcL/eVkD2FlKhbKhSMcv7dZKSyzW
Y/XHPlkcXRT3228wdN4vfqFo5X3NEfzzU8TSrdgHoH2IcijNu9SyMML78ZnTPQXt
N1iQHuGjTJGggNVRJ0qacIhMaTiTZnQGP00H0bWeQBVbZ3iTCqSecab9Of8lKmvj
MpVlhQb2+bYpE7hzwoL1LvsO1ZmbHhbSX0uT11fCcqWLbGyspPOQj/TBngTZNFIL
KYwHOKCJlg3rogQfrHphtJuwhsLzusnVl/hmNiDTqbzRf7vR2CRJSwbwmYHYwRoO
A3uC1YE4y55lxItaufDf7lQOEuSyMaPsz3YHHhb94zga2msIVMq8HD5td8Wzg5Vn
PN9ROBoUQf2nc+FkR333hb7efe+iPk5U4S2ldYCleIBZtRzBdFmHZKM2fbrpxA6W
nF7qFKzkVVvV5g2DxTjuxjHbQt8l4Rp53if7S3ON9dgLTlOUOkLcNTOLaV4IEJSX
LgHKbb1Z5CUkobymqQvPjSsk/f2LEFV8TLOHcrMWHm8aZ7GX91ExsxPxGSpHnW/f
Xr92aYaMqHgmVDP3OQuZ1C6+e+oNYsKksciLC+YAdwzFeP535XjIuEiUFIqQQgNm
FMV9v7TLe62aFprz6BqFt5mrF3NkpCce88GVB3ZAV9JUtXm3/tK4HMFdUqsGKtNG
co+s5fV+K5PyIxQhF05AmT09naCXNeEplWH30CsRteBkh0srJh8ixSaE/LREoFn0
UQTNzU2ndf6fJwZPCDvR06QGQe1INTAV1KSsEuR35M/eNiSzQHsX1cr8tXOT7SGi
P6i59g+CLPVcC81BE4omfyZY61O8SH5oexYD8cvjApGhYuXqXJir5fRvhw+nQhhR
zcfeoxm3BfYo9+WfzkamZXxWPFCuXUExA1JcACbq57+tWIF+czy/coKJxN/+Ph55
iQR2ll9Yo5YDiWhLNXycnO11NMlbtS9441uJvrnfPxYFyQxl072LCb5UEMvanwjW
G1gF6pde8kna9phNkxy8uos2JWtKHxESqQ5u3cLW7smutmwMgbUAaWho6uQliYVd
lBaSCl+cwmJW99mBTzCFfTdJgcV2F6VGSdcBIj1avl3YQbAaoDGiekdt7sSYFVP9
PLoezut9TLtXO36TLK2z/Ag/6DNXb6//Orw1bADozHcnULxRmCt/47OLYF4HVGsJ
Nvw8P5SUZiJ5/9fv/qvAkCUcGBYDEzZV+dkucTwCZCzsbEX3wi921lVH9bdbiwOX
kvQrNg3ToTj2X5Jy0QcRLTx8yAjNIFwPFQ3aqAoBI0IVzXXpMqAIJNsTY0j5caWH
FX6+hgccG/4ztLRIVtosuXL2wh58+wEVRvXzdjOvLbf1igbm+HiooWZHTNDgcHxO
3CY9KUvvguHI2YojBdiIY/Yqy7GwPBwcyF5QmtxjzCuBhAts5HwDAcPa4951MzfV
gSGu4P9mPRKAOpChwpk9Q2KUhPc8K5zfs2SDgKzpSR0Ab2UhlzlXak2wttyeBxHr
fhIsKcxzpKhI00BiaqKea8hkUxyXBfY8iJZdtKrXUklwdjtxGqISLFHA75lRd3h1
XCdsMPoB1QA5Zx19haaGzcAWlregMV+f1u+ffSk+0vaM4qHGS+rO6Y/pw21yGnO7
ew5s1YQBYR4KNHqdTmPFiJdrZcfwwZP9MRFFIE/hVpnNuLOHOitddz/lTzh8qKHD
EKpXvSQ+UdQGOc2uV/+kbUkHox9xOAF64HK3mt7Xmyf+gqxkfMYRCivKur9+f4kx
KZOPrgcB8kLneNk7NJ/j6SpQc84/B9/GBGXg8ChKwCFwJsV933Hw8a4K3apqc8be
yZPAc6KK6ba/ObsM2hSDVpy5t7xb/M3cAgmlsQYRh85drbdFYV07oQtEqv/IXohl
5s8+JSnJoTxNhy0n3OE5YDa2iJKnehRWJdI05FnwdCyxKMkkOXWwFgMEfJXlCQ8R
z9ySHt1v+HPN+k5PfNJy+KmC3EjB7skENEInu4SaMPDBOB/Y0N6DaCih1WShmp18
an3C3o0DzKdu9/cOnzMvINi5+5HHYAdS7qWqXUTruRF4WF+MO8zj2tdj1eYi9FOS
XN8cFZbztgctRB2cvq6daq8VDlojPgDd7bQpLqcfhKKkGm/KYwx+RxqF20sPQj68
LezsyYwMpB3mE8MswQSAuUXNaER7JY7mguFscuDVQ3Kf+wq3eCcOMVc74fPXu5hA
kR3roGwIXEHrsvMy3pMxUlTFY3IRl5xqdA1nJ/S8MKuvA7jQp013pE1tNi8Cq7t1
P9M4bvj6OV0G3VPlcbEN+xVLJthP94s5cn2gpndonQopt2cMwLRwh6iYlynbqlKA
xQFHYqmy4h7eWYS2GIMET9F/XwfrT9Qks1SH9avIMPtXU2k5lr/itnVstZK60/0a
Z+Q0FVtFSjtU2BBGCO3P3w8OzzPkQ3x3Jkp3Ks5KzoxzH3TcT8gtUr69DwXME96m
BAQd086wBVw3RWaoKvJJeeBebGI3h8l+08s5rT8+UI4tfozbv7dz7OnjLybjZEe9
s9Q43LI2pR17mHjma6WUsyc76C4kfjZESPq2U9/4QjhBrjn3Udbh/RnVQovGP5ZR
vm+Juem0L4GiF7PwgQsfJMxIxEpbVUDKCDtuUBtluyrsBtPlbDkKnCwDvi3uaBM6
5WFa5aVWNMitN0oGoRa01C2x2wSJf38PeT1VHII4bKsDW5N6wCNBCztlFR52Yi/3
Y4KCZ9ISOI3N9wWKuA6vKtUgXsvv7sawpC+F0/Let/hgfquh/ybGigIaoWF+H0Fa
Q+JC9K4G5H2tymF6Qwb47A37jQ+PO7ZENFGdsjwrbijXMUwOD/gYM5oKGvYFT496
KHFmEVv0lKmZ9NpIxplAbOp4/A3Brcb8wPQQVSf/upQ6J02575tuNCLSZnurG5IT
WpHvjxufLG6SiHgTju/eUdsLounjHmH+Ba3N8PvTqHRjb16hoaTQkthbRw5lVwND
hXshpmoTzMv01NdzDrjxogjUxbHBM2Z717glV4mbBzSScdQwexQBv8eMIB98tXNL
I+io7CAby9imPR/HJDlkiZ0Hp9uA7NAziwx7Bf9eELNVrW/X4H7yHRC8sDAs3hu/
n6Olu9MQAX1t4Auv4bCnct6YvtkED/lawZWTAUxtVddFN6XCj1yFbgHx4Q83YpJI
eMbQPYx7a0avfbGUdh2C5lC9Kkh491GMD7DiupOJWU5CZAoDuo1eejEasDv2wJ8K
e1oYNDY1oTS889bGPaHQnuKeZ+08WPquC1Bzp0RpsnK2s6sIrHnghFNMeO4S9i7L
WegmddBuXy1PcRdONB2pWA7anlEVsAFxUUhPVbsxnLq83HYGsQQiwqcF+fONEWmh
4sQM+ypGaWY0yno6+qHDZBlnsNWUOuKVV6OQYyCZuHMpSCIJYA+iGYkk4PAUbOJ2
OZ1gf5X1rHGFwu2JjqX11XQS0MjuycII7sEmuWJcpZnkBWwZ/5RFcqVPpcQpZus8
UcT9mfCL+WtZcZPhgQIR+uiPnwr0U/QfpLb1gfnueishBl4KzQSuefd0LNY8gjKY
Wx+ViRBHV+CfFzJmuxiZAjOM9/bOQTsbzfy85JsdpnRjHthDv4NlmHA2dIz1osTs
RoUABKx2JayqShiF/B3VbI2xjBbfg2hb8WLtPl0ykz/ZrXfOwM/ZeNhnp+heOU/s
yGT4p1cq4NLKHEfzxjoRysHUrmVOBL2l0jJhq2nUjtPrYiPRH91orfBU8RGRMaxh
s4iCIqXzumoQaxE50iwLUuagII3TSNjxysiXOMSzjk17Hgpudn3wI9Nm6M/j6qlm
Ml+rw9pGtr5b7zVTkBTF39kS79+JXnoQHcjbv2Ma13qanlCTqQSRR2XiUMIweooP
qiECdIVPY5OXgpBHrS7E/wqFIBILrwYFHam9n4+6NnF5rToVF+LbXGY4uwu0w3CO
M3u99U45WV62ZBpX/RD3nUyaFD1ofyKloYuScPUql+OHuuMWviZpp1xl+1f/fUEp
MTCmcub0XILIY0QIeim4Z5tH7AU3EV6EioLrCQcqStZlu2yn/akyQsUOhElE20J3
fNb1U4ZolQd4ykNH5FVwvV2A/6078yaM74VAIxqYAeS99iQl07sT57GB+ypfGVnn
PrNWzlQ1KUs/8QdYBIBzWAP1/YM8RytrRqlVp2aZOwhgBLjf1tkBsnscE+9R0IY6
qE3ggDGNib/W8iCw1AxL8Of80z974RsdsQov+vWuQaibhm0DBQs1pgpvBn9gK28y
y1OWjxs691dSOGXV36hT+XyfCY9CrfZWbLwlZNotW9ysaDYrMmYy/xtXxAlmevn3
s3jJBQFeu55MpFyG3+9EThgXS5/5l2zFzbPnMoqUMfIrWKVTCuk4lUOEKlN2nIEu
kwE0sHU9sxyEdpBcO/FZ4EA3cY+80jo/BCrrFjZWbmezkGV86NeFV5ZEWOGZGLL8
ONqDhTeUxxHWLvgL0KPzT2mIWVbzuFR/bb2S49OpsIsk2amZIdbaWwamexjrrnvf
O3GjXiL0CPfq7OCPUdGwR2unDAoXG8Cb68c1ApXzKwKQJHWjd6d4BwBAf59N1+eX
5pPrRXIiKAhC/5VsqVnxaYl8FRURRk8HAeiHXiun/1Sz9Li7e08Z1Vm8A6DE7nlJ
hV0TNJFmf6p5aTuvfUcRhbbD9OSNh6or6ZgdCW4p/zuXPbmrOcXUSRYL4+W4BYN+
kDFCItO8u8QLG8s99odt9Lz3mYjrSYCVcOXZgqcKUMASKEAO4UEZgMMaR14znAhY
keIt+llNgEY+5GD0sgOtNSY7AfgFgQ0r0VZQe9nS5GXLENvNuNG9g+ORGpwTjj/O
3YOPCR4zeXB4xPqxQTqEVAgaRCJs8iLxeapVi20HW1+J4v8vO9gU26PmnOkYWwMO
3cHemB/JB2Ndk3m44Y2yhJg+wMYQeg9+vV0i+kYFhxkmBCmOepIXBUudFrT1F3ox
aKwC0SW9upwMRdcfZKnItLaVMiVH3sQgYy/AgMkNyJtH4bp34eeDpvCCysbObGd/
/gLRLZYzEZrWNmAA6pd+iHoWP06jEUNcK3BUBWWAHjA5rQMo00jAzKjw6qPgKvLZ
uQIrxbRQ21O+jrlWcKMUHyyozhRbnwGhlGy4nOtKS8p/ktL82fXuLvP+5CccRhW4
J15OSHzYoPgUpZbw2C3GdfjiZJkDMU0pSNnwDCPIw/1l2672fI6pcI8Brje7dfqp
/YKdU6Zgtf6nH8sI8EEsf2AB0Y5/nDXm8WuSNS9+v8sIrJ/Ps9sCLtGI8CV7ODnZ
RpUMbzNbBQc6+AMrzhbN61nK0UsW+HKVMqfElrd6+cUJrUtiacmkgroE1t0B3DZM
liJPv0BYeJT191IYCKQRdiqitaXNqXZn0Ap1gHhG1MHCUiRNt+vyarR0XV8n1vcT
Rdhc6pT8UzUBMprwlAdUcAAe7UMU9RR4tfdP3Ebl0n04FoI9a+6Pg6VUKK9W1MMb
mXntTR/YAFX6CNEI5RGSxLC2IqK5G2uZ617Of68WEJHmkCl2LqXsyuhNzEH0kz2r
COn2p6EeaJDvbA9xBIfV+7MVaGFZX+1WO6G5A1JkSzmLug3uzi+t42Kx9WJEz3lb
fhhq9I4Obs/BUKFJT2mvWxaGFMjUvZthP36/NocNqtTSDIJDwK3QXLfQm1ykNzzx
kyiPaCCMhXcurNYSn2+FOVgDu96oTJeXPjg/Oixpk6DwBGcggc6v1gxOiGb6H1VL
KtapgNt56fILgIUmrABTg+g02F2PFNQhB7HFpDdgetpnbqT5eUrIdu9K4Acs5zF+
a2lrF8cqJ33/4wsFvjhm1N/bQ/zq3AnOcnXvyn9fy3HFzPKLyLCA/4Uhs9Zp/wiU
R5E4w8eDtWLS9k8fTrdakzqCITAfOvXucIOXP0cjSRu1KpBbOjyLI+fOSDd8ag93
YTTmR1qpCmvcZjvFuvriwif/dh7t91FjUD3lcGKncMnGlA5OLO7vDzAt3OPj/gsQ
8mHys82OYb36kXmRn5idyVUMUs6iHyTnOCqIyUrGnKhjUN3fYSCKc3VJyBnYtzIe
+KS5BoTMbDNz7fePsCmtlM6g4DyGf1YZij/p3AXDNbLPI1S7PlxfESms6eMEXfOa
rmYO8NIjBxLrZQprEyc3s38DnGxOX7iPAHg6+XVmnuzog+doAHGpBo9zBnidcT1c
N3iqXHkllR2RXtq02Cvu8sOZsFCC4Dorl3rWBf9Ne67tzsJnlr5wI46823SgBcGh
6ewHWJTaA9vCeb1HBb3Wr0NN8crc84caJVc8sseuzkBw3kdP/jmjroKQ8v5c++50
dEMLloSAqO74kY4qUxiggtjI9B7tIFVE312mx84SRhXzlFDm3pYHoNmzqfS0O5G3
bZ2SQUrSnEX0I5rENjsW3/N6eu6mD2OWuIh3hfeZWEYHCDJO0gcTJ8JUE03BtV/s
J5PMjMvuYQLVZubUFO4nJb7euGnKZlv8f6lQswLwXE1xJ+BeXB4fL31NZXivrsb2
WUqkiIHilfGaX9IPa24XXsEyULiFIRSgj/dus8aNk3HRvVv47cfEvPUjtDsUOMOL
wDvstq3MXC/zBbiFZ06uHLOksw5NxZtTfdI2q1M50RStc4l/fOjn1mGJzNjGl5GP
MEiFDHjac3JrNMa17i8XAS2srrHfmy4L4hJqSM91scMYWdreM9Xzk+I6J/BupQmB
IdatQzaD+8LBesNT1xfActVEH74/fkz8afgHY/+U7mcxt0FbU05454KgtXFI7JL9
gpxY+J5YHCOQMNejGduI5PjPqDzbjtGp7dIG4uxx1z+48nrkuq1CKiBVgfrxoSoS
SCFnz7d+3QxHKghDJ2H4GS0ysANBaNGgVD9mbbQ5x4eIKNng0JUQU26aYbBmH0vV
B9bXgdp4ioUbiW1pB4gAp7dF4SagKP6FTuyhytBeLxaTp2lNNjC8G2EkI3m4IpAo
RbbU16VBfkjE7Leet+5WszBHuSzZFpD9VeY8gq4pHdb2O/cicAeztFleMj+/wZBf
Hv547GoyS+Qti6ShD5HMdx2+ApvZYUzmIiNHsoqF8UXzd9nDgZTxhL2OHRUd7Dx4
BXnG4bpKW1Yqu74rmFiymAgkdqBmUxeMVG4sb0DzvRHpLPkiBs3GhXuc2tdr/p5y
Ut5LYi5wSlNdR7XokIrsmwtTbRjpeez0EPKl7NtmGIC3iFEAczD5wHwZmJpZh+vS
sscUII5VI7Kq265vUGytlpAPsy36Zel68f22BSApxfgYif0Id5P4SLoVX0rPj6aE
ISNsevIRmIQQSvUTU2dY7XMA70qwnbZOsT9IDgyxug2xN5tCtMjj9Ln+zzksLjtc
Rzjjmu9MSov9dbLMasWk9dfDxbkZ+l7WDJE6JhC3XP/dTgeJLbKyP9QiopXsFqPf
5aTXYPWqbv90uQGmf/gyRhcrz2Upf8pjrk4bR6hAaV6Gm/VkrlH/KM9/MeN5cTX1
61+AbTOmVOGd+u/ubYiJVIaqvNQcaI2bjLJewnzmyUNtgYI9QK2h4svECg3fZnmM
MGlQ5AVYVqV3lITjQnd08EyjbBJRkMLf255RvHwppmlg6F+DPVtralalnyZ9t6oQ
y28d206rphBVAqVX1+F4z2ttL6/Hnxau2FYvsNH3PW/rrjK7SLGE8SAF9cDk9hE6
CeqgsrM7uaYbqWCVIpe7ljzUxA+MBrrhtqCBst1uYc/cEjAav6/MUnvtit9txdGT
YLG0qfQbgDiuvQiABWBGKidhUPTqPSyB2PDIDG7Vr6hOuARPj3f5OQEdfduqS/1n
UlARTr0yNdkAJ4lnrMkDzqHx68LpsGGziSLT4zuPl7lM4yATyKB0Tg8VX2lcyhkq
b7P8E4UIkZf1I6Pgk+8SfB1ZFAWKS+790m5fM/G7fjj0hkZ3wi6ztGLxONCehJ88
ICF97/x7jnSmxWjNqVH5jm8AC0PjJhq1QjSp+efBEDeROyvCpJw7oLJoB2hBTg/W
18mdReNT3usnQokgX77HZHys3CpwQ/177xSsJhxnvGu3wWSV83qiPBYUrKxT3EV3
yOJUwBDgX9zGHKMO89kQ2UIj4Myk1l5FdF2x8A4XgXfVT5WeTZ3L7uVY769BPm1L
vVB0LDvRK4vpvgiHRR1Z6jeQjeJVODVyu7dJsXzhnycANQLOeNry6Kiw5+4RCyVD
1Ln+XmN1xfGBT+gamJeE0bHE+01RRvcvsOlKzZ8LLHaC3OWGV2WIHX9FG1sU/S7y
/Qu8DHXadcuIdortklCAf3GwMEgSam3H2kx2QBTKwDwPNo0EXvPn88lgpupA8agh
GPMjBdCOG+M1p4rew3trEOWE6jF1D0Yj+kq8YOOEMP9G2phi/YbYWeAP6aPPVCTE
bpYXL5Uejx60o6TudxhYk3Z+i6myAU1uAvzWXrL6DQhb3K0tSx7414FJ+nLsb9d0
UIEDwr2104GVcwXXsFw6Zy8/effKP1HSqUNyzs4yDtQ2xO2IwkRW94Vya8rseJXg
ksMxteyf84pJwFZyCSMIL+lKnb0NznvKXKpiFaCkSYU+sz1PbStIR85Rs6gLZwYU
fKM372EFMD8pjN4Qh8sETBzKk91aIxPwHPfKmG9eLT7jNgLGFKSlLW7fRaR9Q4yT
9svJ0FthfNk9/4ulLlHOCfk7jmpTlEt01SE3rvNwzEQZSQ7CbjEZPF/fyC99JglC
HtbjdHJ9Z89gwHL7BCXPbBlRss7qzSzNoqirA5jyncG2upI3swzZrjeT74ifUNQ7
WjTo2RQPF0AQA6Z4ka/OfyVfK4aBxwBx+FCkUuJMFjY8gj09E7/URgAbkPmjU0TX
e8Kd1ui2ej1ngl1dC62x8e14njToo0hJoRcp88CmZX5eShs0npgFzgZaD9YeGAnh
AaQoMQnHndEnZnk9YUMa5zZfI5BS07gn/7J2YXhsD4ha/lr4+pZvirgGIuBJSJYX
jhhUPywZcGea9HnG7glnPfMcujzWO0fRNwjqrgOhITJGS8Kps/tGc6KA1jaDB56+
nE6Ym6t4aawUVmq0yVaNfelbMlwI1mgjka6nXlVuMs/XA62QUh7/cP5ryDlYpJFG
pAlkCT/9VBSVGySBzjs+sEoj16ZUb5ilQvdTfMTBOlXLDU56zYWCutL5MMyFC1s3
avNzYYquNLZmYFSsJItd+Ik+/po8IhE2ha55veubB+DEbGziG21mZTfwfFnLLv4r
/NXd5u6DX8iwB5dwHDNyVzOleWOS+NL3QUDJhreG+t2zH/cHm1aUFKxfDL5mP2g9
axlOO3I6at6rS3l7uVBVAcg2WvcioicXwUOfA493hABIgdOAYjafrbJClpFfZaZr
yvMeiV80dyl1D7KDByk0KTSJ01pIKB66rkKW2dmH59nNm2oKZ29Mnl7zot8KUXxh
K+Of6As7fOUrlQ2A0mKlvkC4k9MOUqjCyhl56FPJDT/Qd6YnhE/k/vuYl8BsGf6e
yLXF/J5HOUUtLJKVbvC0T34FrqaFTMj3dCMQ4Vo0T8/vQAsMGsAVzTQ/BxeRLI5O
oecu5PqdKKAGK8Lt7U0NK7/D5PSN90VYFfJC89sYpIiFunAlBmHatPbH30WaH+RX
qYyk0G9qzdZaRJdM2InLep0Y2wJ/0gGtWCQREMOCwWjChs8jOwd3z0ZlHdwVJ+vC
X/c6YPkIFDEmhtXi95yl5m/7s1DJinlPJ974j0X38I4MHADqW2fVR3zvI63QqfwE
93tNfQHDHl0uGuJh5+dRHf9vRcsZocFOa5NS7wPIHV+UFblBpSTGdyLVFJ1xa5K5
VS8ELUjgCoyHQ3SEUu6AK219s+kgbexRzYiYAPffMrksD3xnXQ/rZpcg/FWSFz+3
+/LQpfWmA2/5dN5879QrLua2dFQDdHBBzxq1bXZRfuEdL+XLHwgTSCd8cn9tOYrp
0gMLBH/3Po9ZijQrfelixNZMul2ZFQbm8Ja6lzUMFyPj6Uzo/0Owdzb4+mUAr/Ke
r5ox2Y9sGJlG6jUOjBo7inswroTLZy0SWQYK7rF6WM03Vy3esA2BDl18nzNKtqT+
uFwrpXQbqNldm85v0FKaXeV+I0gfhgwLJ940/4/yiOUJeLqxSM6GBhnmp4MijtE1
nU/dFEZCUf4vgDF00/1woDJmgEKeelKGQlOcFmPPsqhdHHSG4vyO8JMWqf4AT34Q
0tEUVYZBMH3OGFj/ZJNgkFSSC8C1kexcmEY/5wcmSGqLl6M0w8EurDulY7z0DltC
yuYwlf4NPjUaaex8ZnLZjFWMKiK36En0yRjvznKfkS/ArAx8ueXKOV7ygCNl+io7
f6GMz9HINfWDwBKa+8Hm28aicobFJ+aF3wJX5tBrKWP6uAG5dnGpwI552ira/Hes
WdtKvvQIuuTpPRP+NYkZCo0fEhvecNl3lIuWqfC7qATAcQScCpVQxMKiLkcg9xaS
DqG6z6ph0jDnyowe+SlslBtCfaufibR8Qgcp+pvmZyXSKlwpp9zbi4pze6YrVZ13
rZA+AFh8Wsm1zhcR1WATDCU+FWl3wdHQ217i48GGB5f3mE7k/clmUmwx3azrRLST
HtjVoF2Arua+GslqDypK+EFnIT2cFPRPajTKnavmAcdv1D1xl7FEJjwaDueX/+cZ
6uHcvVAFdjhi1uZS0SI8xtwdPuX06WZal5CRPxpXqNiIEK5KiBkrIRfsX8iAEo89
YvMiR9cnbCO3BSJnm3ALRNDKlorH24sCFuQB3w/tOCHLFp0PF8uYyPL96dAev4AL
+OdD2mzToA1AOztr8CS4mrK6g6ob0r+MQRyFeFEwV3t5L7ftzEjZ0bsaWYCU41x0
zd3VqYGLvfKzt6sjQoIQo0AFwuOns95XPUi8KxubhK7LJexpT+k25FZDv6mDaqYD
cR5DKKuXxSPODNKAC0Y8v3eIZLRscZ8sEBrfapmkBgV5EXDPkDS+RT81prQhsl6h
EiOH0OHHAGl4TIlmAngoxKXfb5OTpAlYOZsWTMzXbgHYRNzeU8qnW5aoMHTUYcDP
CSz52nWnrMoHsvuhlt/Ro0RQFtx4znOXX5m6wgtoEneBYvQmjtFezj+vqM+GVpWd
OwO1LV5mXxRv8EpTD+2u7A96eUnycpsI6KyFYmdA0y+pz3nWy6YTFnaoA9VZNArt
HKSTyGSfaJ6hKvSwB0/VKQDQm3DXNeQ3/cEgxbvVjj+dmq65QBvtrOZOXoM+v2LF
aRCZGmk56BqqFl8K0HWFWQfPX4jjSoQyjv3G11lWjzjio0PeVWM6hqy3QxVhks0M
uZXsWOYcYMtEn0oVnt+NcrIq5Dts4ps5aPRm9aKqSznLMF0MIND0ZCfUSzAPXHJ7
pgaHl06vWCQG9ps58SLfusR3Cm4WUmGdYWZaWpCQY2Gh5YYGFS45l2qzB/UFYAPt
qdyjk453Y/7P3Wkz97mpuLHS7ir8ol7O9AJfdCO5UUc++SJsLOu6oKRXFUH/BVVV
LyKBDKsBc9e4dRZo1ozkTCxsez7EHqgJncbJudbKA8dP3DAnYpAOf3NEmq/8J1p5
rNCXdyXm74j2ncuJd7Z+REM/lcYkKWGQ2iDIl1mclCNVEVwoCsrTwgHJywoNNMK4
rKw7ePptj5lMCbxTJ7R+qae77tsAfxGGfpY6ouAZt5ZT9SZvF/snDRHpVXJWRA1i
p3dYkfPYgGF9ZL/hKwtZkXtfYsseP9GKMaPRzuVdZh1E915pwBn93rfgke4tfkRF
ABxyPqfl59tE9mXjPcIsj+VRBBz6XVviCY0Pjv9ljfR8bmXAmUdHfLFbHwsLhckW
luySSybgz+LHvoYbzwhAnVyR6b9S2ZYCLG5iE+Dw7nFN7ang+mNjZsDZDk0PcT4S
2wV0dKvKIy6cUs1ufkv6IVbC19JYRvJH1Ccjnj+CxZzQhKafow4rObVonLsRha4I
d8TUSnr2aIB8xnnb1eKJ4k5EpKXdlMsHj64AyoWixfU0hK/rwcUs7MeqfgCilTD3
qUOOsPDxMOpSkv0SfzOuXee9I4a+kMrHVYzhb3+ujml9YY9E0ZoT0RHCxVbtlJYI
6YWvn3wYGrFhC0ZI91MYgf7WJ1Nj2Kf2dlc7pzivvhLPMypTb9L1WZDIfDM65rhM
VT/8khdoZnugzb0uyLcxTMTRDOodn/dqH/FxgF6oG0nbO0FPAndQJXZb20kV0Rr0
z0Hgzpdbg4mYvotcWI74zLsJ8aLZfRFcQzwUeOUAWqU9qky8uB9T4ea0oHzR6R8T
6/SKHY8ZyUSa1oUwWIZu1vo3jMsYzTGurX+vUqhjWCzWXK5agBbG2460hbqNQpor
BHut0Ib7JVFrJHQWOF1CeGqjRJ3+BybY2WPg8MrauGb3QZPl8Sj44JBzsmjnrUlr
c56pjkCZQTtgtb1bRkMLaB462F8Xgye0y6WFkUwadKatPkSo8vnHuUVOmI+OHIGD
xWD2MEalRmwqr3Tl1SSuk3l4IGyGSWk11leaUfL93uKNRpQxi8X16cRyltKLnBJH
NNUrleoIB0J47Qdzpjlkv+x6r1wB5ThGF+dc3F2vOVarjzHJOLtIUitCO+ugZHlX
Mn093rhRUSOy237iW2B6SmYr56kiqxxXPIXQJyjmF5FI9M+aCLjBY7apAGvdK9rm
rIXE6GnMUoDw3kWYef0/3tcV05qts4P5xADxVDNyZCo430YPdXho44PJoppRwfWj
ATa+N6OD1xVC4hA2NZLdwLv4n3ER6rY4muJUflTBMl0iuGvxPD9OcvP3sbw5JC0k
j3eNMTl3VzssUMNsy0otapVB3iBIe2sMn16CrNU4K6sFe9lol0OPkmJiE7hW7xVr
VVjWRRIk76uHReS9oTQE9gx/oNqpWvHKOtZtP3RJlF038crzqx+CVXm48JHSh64o
+w5Z1Soo5CerVdEK0HZBbxuNQXdeUdUvIxbv+YesQBjvPoV7TFDcI6TXwlsm2tf4
ee8RPq+wBTZ5qtaVlunE92EAw+J2TtVuVQr9gwRJNvA4957IdNLCFLGEyefmNkrX
R4iPowC5mLVyg3E5Emf/ZvUHr2OnA9Vo0rcGvbW3Xd6epdHHbxyGpNrnxsnpvdKp
RYv+qGiKzIoblvDVviJHqUubtBzGmHpcrabcrariO6WPuBZ4yfqUdF363s6hLlmb
Xc8qX+ssn6c2JKbLGpDWdRIzjsVpuR+WBcyC81qoiu6TRoNk8BGiwRNyjcDWpC64
tUQ9Exh9drDdEFlsrKW0uxYvhZZY8t3ENgI9EwbGgvwLH6pwhqKEKHtSj7k/HmB+
bo5YhF4Vm44zflYtQyqBPPlRBLuOkDATao+IkkstQFbsXjhjSWSxDURsVWTRDjx0
a54/n4+EHEQpgQ2tjUCNCTcyuCKTudMVGdEIzDzHWHSZY6DL8zvXUA0YPH5n4iXz
Xr+YobWKG0AUNOZkABHokiGW5q88ccodpe/xL3d8RNtxzxGM7GH3dpVE5zOtDlLX
yMSNjzdtRMhMJYfKBNlMqMdHrxfm9QWXfRuOxs6R9kbTcmHssB3A0Y1MnNKOjBqo
l9cPs3IDjMop7/Qoykx2lKc17qgG4zjI7Ziay4g9SghaMRsEk1of7cDX+Gl1pgJX
m275to9/CTQ1XoIjc5SQHRh+Qs5GrBBLQcfve3SET7tH4v5sWvBrtWA+0pcUFa/1
1wwQNndGG+IPhCLOatwI48a4PpCxfgSrtzODmu/UcDakH3T1cpcedjhuvxtP0sBM
9XekMjWwduEnWakUUuaDANflJKsDrERXD60/qA7aUsefWdMRC4FD1b5FOM5Kix6P
O8lqREZHMBN8rEMCDXokOYrhed/vTjHdmFBgGGtNU5EuKfzHoYhPdN61XzZSRjNy
IIGolsjSc/7sJMhPqz5AyI4nNBefXXtirE/xcxbi7jIpQKjnwH4bWMhjjbfT0cxU
k6ECX7x6R2rA4lmtWR+gdZAaNE8sLxV3/5u4JMradPNvjQmN2pWqiJ4c939TZK0d
Lot1ge8V5rGaqPseUtqfcw7NNbbEnzTx8R5ES0mhvrEQdxXvCDOTErut0A8XahRu
vIPE+xPxnYzjzGP/qL3V9eeJDV5qyd4W+rj8N4r/wpZ/jREwbvheDLbsHG7rhPUK
RGUUPm76uA7+jc686tm2wPtiah7O3Buy/qQlbw+wiOt0YvLQVoScdmyzhdGpktIB
ctXzI2KgG5HPfmcP5YLc/05Ae9OvvT9MOhrHESOrCEIm4nNeaCqo+DGchan7n2VZ
Qb/HZfXH/hkI8DwNaRKX02iR/TdZfQKUYKULVUe9Or9tITQSxHjpqNpo/2POJAcY
eNQVVLf1B0FWnwjyuHdO81watWgxbPLHqfujRKyOzAO+oFUkV3HHN2fFuYUlrn1W
VXPxF/CxQl+ZuEu6sbcgaZepDcKv9escq7gCcb4R7ZaCUk3GByKuHkNSrvp1NB/o
55wciRXOWCXrZQnd2LxBA3nlUypsGQzJK5Rl+/VWUrMWuHetI+V3mbeiKav2F4Wv
iyzTsZoJi05kx3nH8RsN5XXvLae/k81rssGU3wIJ6ZTMrBb80qulv8ZZuMik1St4
EGPhr5AQKVmj04zUQdWPkQIDszf9oaqK5TbPL9kysj5Te0klvkJyQMpYZGWg+hc1
vRn1Icl8M1/NCzIy3fpVZj4SjHCBvfyyBsn/TEqYyl5K39Ni+0U30vnSJzuCc4Dd
e5qnBjC0aqwfZv+P3XGaHvuBLDuHEcQt4eGf0WlJ8LnGT3xJ35DKW+MHwJlJ713K
uVgw+WhEp7ATAWdcXyjgHT7jfPu/acP+PZej13gJyOabxhcppBng/Zv6/WGGl0PO
IKY2wT5qEuJLHxWKoJFxK8XFX0c8Jv9lZgCpLiE6Nv7hrh3+P/75OYRBKm/A8RQA
KwDnM3pkkMJBqYj/bTs48WJtWpXAlJ3sROmJUVTSjWpf8hTtljUHj3Qgmfi5PpLL
DOMRjx4WB9lmfwReM6e6cq2gu7PSruTGiKEIceMmvsHj3Q4UCo3Xv58k5uz9v0pX
pnoQCjO1Zr3F1RY6n7HNMQiCx9QDaw2C6c7yLwpnKOLFy2G5HMkcLP7tm/IpWfgU
bLaZGF8VdC7uflu6/5jsJYWOze4YLND7MF00zF2RJVsxfkfW4k3mrhs1GP9OYpPi
JNXEwY/+qZRceW/QOFzsPQqnmYmZ5TEJR5stDtV7hD6U+uG2WKV/lWV8JNfnL5YC
RDLBP9HQQG1g8WyVc1l4yQfxbgcGyqSgOULDHp351xhusTmIiA/qHZdpXYhq9sn/
cjDcwxHsPnLF+OoQNcBhFqxZ7QFkawlKfPHGs2LYUeAVXpDdyTtc8CdxXQjc79To
kiWcdB1C5RvzDa6SOehSKuV62NB5NCby5ZjyAYLsmnppibjy+qULNlxsEaCJnzif
YnXImQ9jQ0VtMBItc+lyZzof+0GcR79z18QTO2xj3YN9Dn3tmsEaWmHx1DLLADpB
lcvp3onVdtESUcSnxJ+cxVvfN8FaT5q0AE+VgQWW4ZBmQQxXc96bHB6e1I9ixWK5
SWa9HlbV8ClMYXwqGzhh5kvCtASIn/LeHpWrVye99qStY/bnuH8aAAiVjUt0c0ai
Gx6sh8VQPcQVCQyTawqyzaJzi/nFZSGisi+3xA82ELbHx0HuP6nvPdC+mI4pJ3a8
YK11om/CoAtL8AM04RNf3CLR2QqCOMUWyZisurq+X48MilPvdXwO8sNI7eywiGll
GCeB3XH6haFS+2b8cBcPU+1hKZYvfeRR0BP0kR/ZDSDXBL1Tb/c/8VpDewBU+1Eo
raSJEjpZ/B7itFATmjV4Sr9yBUpDoAeLA1FaPXXQNzUzIdCBN4TRZUtV1J6dc8WS
wiiTTHaDiAzWZI0S7OrBxlXpHv8ID69oAgdcTrw2PRymGmLNizQERaLZWcF1xJie
OedXFNv8tTKHJcLmdy5YPC74dxrXcM1vVlj0jymrkLtAvk2G4AIZGZ4kpHFw2RQD
KAs+iyo/FjODh21KNKkNogw2LFOoAOCT+IeTKrIlpgtxnMy94MEFsrypOZF5CeVM
vjl9w/1EJiawKFnXIJ/cc/bJDqs06LsehHKUMhbldPPPILrAR0WWMx32SUaGfnEd
mJSx10WhtiaRu6dGKQdx9eModESS2SKUEzrVZUM6S8/vAw+6X5tFBT15IEci7iOW
vOXIHUESOPfVhuhQ+knkRdL7uLGP9C6bXrBB5IgBxBqqXA3dnQ7kp+j2Xw78qcRp
/Loln2wqCrpkPmyHpGSIyTBYqMW7whqjI4UJPcqFbdx8yy8hef532xK61ge6JaSP
xsXUj/77DpwJJDueMJVQ41mwgfPZqgemzPc018Wq1FDWgrPLQPzIqLo0pLEG886s
pZiCCqksAZ181GfRxLNlZKCGghgCZxFDj0QmK78W26vAoXZBVYF85GbQZ4Q7xw7X
E3N4TLb8AJe/VQcCQM3YH/BMt7NU0s+dIoefWOScBf1x9FXuI2PQrgHiVl3TZbjE
6TcBeJfGiqPQDbbArC4RcrsWnbxvi9xUTTvRAEe/Daplqe2o07DH2sU4Py2PzQAk
XAY1SbwxXST1iMphjDXU3yCAwiTm/+t4CJVJ0AFixT+YoX561X/GG80o8gEfw5Vb
m/7WtQdhfNSpIbNrAqVm0NbjWQSpX+bjmjJpNYQuml3bxCOVoaJ+pbAw+SdRLcvC
LF4q26pbKieBUR0nmTwAvq7Fiee3xs5iW+IWJ+4uLXUtmz23oottrhUL+OS0zP0H
N63taCM9rsjaOZwEhEh2gOFX3ZtBQvwnl76sgnFct2N7tI9fCRN6Ry6ZroigtKBY
jWRFElRp3Doph9XAfDcpfHLjZNujaXHa+9Km1kK39drCqkORxISsaMLGT0BdPcHq
CBj/ZGoGog6co4Y8B8LqK1uWceXNa9vSUo7F7gep2yllhD8Ji1xUxZGEo7d5egsN
vpe9ruPXjlX9SYLIuVxX5cPKHviqRjNiz2ynhlB3dMrc/TGmCtiBZFaqF2OtHlYz
jyQ+dIfTYwdAv24LPQZ8xzh2o8qxkkvCF+6W6oaG+6YUZy5HE3Jricbq4YOPE69C
STSRKE3RYXxHL7+KxwLkwKTQv+dDJZWipw4Sl8wca7C4amrlDnRkZVZjOsscIBFK
+b3tiOEu89i1xgdLEl4wZ0gFqpWF81DiWVrsPXunEUUn8gJgZEkpmv/0Z/2q3GE7
yQzG0b1EGEaLLnCUe/NhDpPVmnnPwqsNsOoYZGC7mipekdYmApIOfwABX1YdHvlx
G+FhPprOoqkKa0vQap01ehtHhp4D+iZ7B5mjGlljOQyQJ1BccQO0XK9p0BSoECDu
lC7N5D2SeFcnCOluxG9OutZM5VWouuZuZPKvg9wq/aAlUZSmNSsG4H2M4/rLbdA+
yyN21Eiz6+LxlGB2vmsFJP26QUu3awtseieSOGXMOCsqVd/RLF1a2gf7T0l4erWT
zbI7zu4sA/loI57lUEzVb8WX48cxcGt9d3kNTaSYcNQNktXyJJN1EGfF1aP/lvrT
mv4a9uHzrm1pAYwWVZAoGti60r9i/nRoyh0Zvus59LUm2jgaIELXk9YzS44RGx5H
g4JmY2HIXGPBbCqRg4SFeSl4HNYepCWYj2Toxgmayw0RXqE0C+MSUJWFErOxTpCP
tITqGVJJKDSZMPnJWZS+wOuzu+nBXPHswKy1xk2R7iSQtUUwvTxpOCTtsDR56k9k
pSySYyLLD+fb2PgVAkdY8Nv4OggpU7yc5k4fa/O4+tqxHm2W5ViAuHIoD0MbhTxj
hpV9eFbusnvzdZC4mI24CnnYqMmESHljWo9xGX0yJ26m/Cr9+fYHtQMgRB5qZczO
iycwwTXwoGUj9ln/J+43ToM6DeB9ja+8A2Y+COw7oPqggyRSTSKsthhScD+Mqcwo
6pEedquWs0/7rm4tBqsTRF1YH+cG0dPRC0KaQ+KnvUepEuxCPj4/DFy4VeWfDm8c
Ub1PVmdjImE9SMxO21vdQmAkjGTlBWED2VoMJwwpdEjILFI8oliY5KtdGKLFnt/i
xxAY/nMl+cA0oLnJ4b0hXdMxN+9qQxyQ9BX4DWojHdb2CfQ/QPQHzvb7dMnsBN41
y1QxTx0ds+Fh+1143UZ44AG9yoOlzSiQUsG8ROdPwdWIe5OxG6WuOpw0pD7NUrKK
tefjH97r06oO3gQv1/D4k909Xgu2O/3fo+/3QCzTo8ytmKGVLRlqgUmtsoBeyViU
tlaoNSgV4P1sqRg1ruambfFJdzkKcWFz9Y6s+k0WqSL+yqMPAqlxyzX4EVL+IxXp
1INy+ECOn0BBUY9cWXyq+sCuhsnSFAUXSamRbximd+b/LrsYb0gNtcpcWTQW7hsO
QNZvfm50kvosTw1yKqz6CF5/E3BQL5xI42abD9dzzBZ13yX7MZ6fdIk0cjeXZ/Jr
hOZTI/f+TfbYhqRlqnJO/2zb4uzZi5FLZavMNZbgwfKNGui9RlCJ6I1q9qWycn0x
KiYca3HCbyG1+QTOgOMPTZOBDWM3jiN081KCfifRJuEv2MZYGIH672VaOSBEoplT
w7w8X2BwKKbXlQITwDNvC61OKAu94oUITbMGkFAiXYlbJWC4/wNXA6McoBLVFDXH
/F3reNiXzedmvHwR7mnrwiyuK5aiDAHr9rCJZvOVWnrCuwIsmlMXxNuYgVrNVgxT
J/8fc7KwuZv4JcqMv+hJcYvhTI7RWD9STMovn7NjrF+cCnfHnTuttJom0hb6nSWl
t+U/7h2r3F2tf7zCDWQlclgoY/8pHIap40W/wS6t2v3q8uMhN+6PnEDzhR65pa5W
nn5j6zExZPyPO7Hlq+JoVnFsitKqU8sXSFz1IzHa3mwtKIBMFsmP7DM4R1WEjgUa
sQnBq4gHEbn37RaQ+r8DgpbqUKdtJ3o3sWNXFKPbA90D1g2jDeXy02ZpnMeWElUg
yWH4W0fqP03dV8eSZRUteSkKiadj3jePDDE8NIt+rI5BG+V18gOQLUpuyQHbWcVM
wEIic6iPNn17LNos25QO5RSfXHktbNO4HqN6PQs/jzdLkLs6t8GSk07QT+O8wSLo
Y3xXO3/a6jZJAVirOXZg4jO1FPWGm++fgS1sZwp76hQaZoy09gBhYA3hLgCzWaXw
P9gep6kG8HSyfB3+IQQhaXTB8ZVAlHc4+ub9atMRDXys8vNv5Y2tuufTiXHNquqF
5WGUbC7elZVyRQ/HWOzLEsoA1Q08idqls5eu8NABsOc4ol0uWZ4zPz3v86/f37u1
meTq0GVlxnNchNsjIeIqdbY0mS0P+mL63t3bN+sUFXWwAiTdu0YUfopoG2Gup4S/
djMmvAYMedXJk8BQdo9bqFmc8sv7CMQiaSdYHl6jeVJIZbrAKGtGFcpkS6X7WrYL
J1xePKAjdblgcq1RNTuOUcUoUClltZrOzsCcCUUq0SSDep+1DSrbg2+rCw90Reeg
QSQmZgLupmDQgXDPFzZeaZDPGF6r0aBazAhlFPd2frOd3dFuiddiJ0M916wQUnxZ
hnETvT6PqL+ADma9PsbLjdkSyOwRpxtbymC9Ecq8m4dOD5UvHENs1XZ3dpJ+qpuR
1xCgtgEMpcVeNQfUtRQAY7rEX+Dd4IBUu49NEAPCQoYS/wR3uPuajzG409H2a8Bc
RMTRWf20dMUhTMRMVqgi1mg0ajjRjSj9xBhD8LVDzpeloMSJS23xs1wUM8T/wd+K
Ddoh2hbAijUUaqOiMXhwj4xJV1I+nYb+riu7RfFsv1sIAaSdhb3mxYgX2YRMSuss
G/I9avawVqYF4+1//1F7WqtqQf3qEAigwd2QMzbdRwu2d+OpqiMjJFRsr0EzyzbM
YxIkERppzH6A4cZ6URQjnypbV6HrKWpKDoDwc4v48j4l9oyLTqf1NXD6Ysh8LYPR
F3asfVunpV7E7HEH1lzIQG9cTVFDZe1gt7XrCko6+eWrbd3sss5zx9+EnbakzXK1
ARPuGpBUWYAvETITGq1pn0TNGFS3HFFVZX9U1cBhI5dYW0UT/RLLhET7Sdnozraf
v+a0TYShsbFusWjjFO9pn8nhOUE9KF84N7CdCKLcvwYiex6gSaJCVehMYsliX2b+
AmqTgv5daTHxzMef/r+KXohL09BD5ywwdqlGNNNQ8Lu/lDH58FPuUeNAxyGQARJI
JyV1vRDzSglYT5O704YgZvrETuiFjU8UdKcStTdqTLmEEJMe4T76w0F1y/VYumPj
+wfCSxnZmxIrepKI5up/FcHOdzh8WE0zOwOHibtxFYreysziCcBUTX2QPH/+YOFY
MxEQGADbc9UoINkm+gA4LixwgDMK5IIRe7O1N8lQVQ27kqFQhDcNQ49XAhA95OF5
9i1lAUDRkesgsyVlHxKX4XJsqz7oF5e1R0UXkgqyTsKRBn8XTx/AJKEmr2YgTFsL
EboHT4aiL9VmzcQ8VGnOLiLXSNjhvaU2TBv6iXjs7TieR6Eia+Vd/uENbaKfO8ny
yKJx849BnNkIy+CRmPPWzndAvzkrlyyQi0n7N5Yrd5kuA0AQd8Kwre0C3Q/QL051
hdA6AhytXK/W5MRe8vdoG2AjMspGFx1o0ll3de5J6nkeKUM9ksb2qF8tpAyx06y6
S4u3ypOt+a8gMp+8Xm35yHx77M2ZaaKazxjRxRTOi4+30uv0BWfHmZ6N5J2xmtc+
+AEqWr52adjkFpGXdVHkmRPYj/AGVKlo9DNf/zPEbAcibTdE+Opl/F6/1ialtdjH
VxMEfL/j3gfWS66ojbOnvUUbgWlBlT4dM9vvmf50KWyClIqbJrQQvGGS3HZ5kAm+
xGFaLKyo83DCGFFlO+AebML7/fm0frhzvryPZlPaHr33P4StcajQPYLqgrzDYaa+
R//xc9AGrgc/o2nBEXTF6qn/uVLY/jRqdss24ZKnoAy3tmZ3HTqEH28vBkfz2qPj
E/8heqh0OtzFgT4SWB8ozbnVHKbDIeN+MRFtgBxS6MAVicOD2kcyH/xwoA8bASlw
+1VWtz5+FR4itKmN9uPfLXORH1nfioeJbVN7bm5E+xWhl+eUdIM1pTBlrs8qhz5y
vc50E087j8lLvYjdItCdeDVN3MYSiUQHyRNlrOH/gBaBnsMTQ/q1yqIPzpi/l3+M
+JoIREcWjUbDFgcBC37T+8TMn6/suKxGjfrvIZB01U396AlKSDWunoYMD6BlAGmA
wSsxujP83dWY+ktSPOxPaXPfhKdzXjOp+EDChdnN4i32teXdTqXM5TKZbv/wwSmX
Av4cjg6SD/zTTzOoZDlpz8kzObp0neGZyU/HIENoFJxcCBjgnewjRHDcbOhPSpWC
PbJgSRqgQ6qG4bjsBmyoXJBpY+y4BaJpiZWV3KvRntsg+zFYYk90gkOC0RLS7YRI
ye5uYppm6mSyuIPiKNZz2o+jlS/Gma55LwOG1ZTRWs+W22tSyq6OFQawqW4XBSW2
irvzP1p4mrCRE1Q8hX9XOOQ9wG8I0jQSF8sDTQvhPJsoEYpd2LqZeamLdTcz53f4
cxpkrcD0MZfD+opXeuT1erBAFGX7kSeJPAsN0rZQ8X0kBRVsoJzm2NMvDZTzjEMW
1ZO/s1BewV5iw0NxJzt2Ir575YSywRwoAyfBsuIgdjOAEb4iKGccNduFbvYss7dW
/ZAjhal8ogzoev8ySKhNK/wDFhM2fbkt1LX5BPQE6LFM06m0piYCVM7fyMUrIOyG
ewW7KOy1IlKugAn3goyN14a81J3FB6TqlhnZl3himSRGBl56I9+CsMmWr2N5/Ygc
7/qaxtF2/mo7BKGh2xON6+Wpf9PN8zWD1vFaZvkh8WRad01GiVTOZ/1gBMe95Kow
22tTWzpkniy5UpbGXPRfUGXGqYcClk1jxoCpC/2KsAdJ6wQ4dzvOpnIpoYxVzHmA
0i9hTqIQV8mLSnJ3dTUrBcfs2dyRcpXOzd+81Y7q+EQSrzTe3JTSbqf3LoqthUQo
pjVxVYDGn22PTegem69k0IAJlz46HrNl/WBw4Pg5kTgnegs2SBuZSbaENOxJ+vqk
GImxLmUu3ZpjGZ2G969IIQC/aKUZGG4ltWATJUovK9KTmbedfwN8+r1+23oxxRkm
7QtEkVadJ0JzUlPoK9fagsBtjqyBb3bKjnRcORXYDEfRf6fvypqXcbtT/yQzhmF8
7RA1vF1SPjGh69XDeVgqebwZ76IKEE6/mtK2TzqEkLe4/lXvqaU8sJBiKd4zGoH0
qmwp7Fz6FBvjPwS16xjJRpcQEJ70HO3THsAQsSLQto9ydxL7WissqWulm0hw+Q2U
gOaoorjxwm9q2lPCBK6z/Dv9Y0AbrVzjB2H+mdyWuGtrJ+vPug12sldVtB/HgLPP
DPpyu5J+cq9Gz2HixXBRTMjT2AXxvAYufNkv/WnWvmC9tMAMSo2Q3qAWCP81QJ0h
A/Ag2GZDbrfMA8sAWEFyUbJWovDVSJOSkZXb0D1I0TLAH1cAtA9SMHVWK9Q8mork
n6ZS3sV1YToIiQyoq9K9HY4ruj7SE/UORZKE0gIInEuLyhrNZPDLE9qVsHf6uTgs
wlSKKkR+krdcLP7bUchgmOF4rlGMO2E7LgiAfaKWx68wbXMvIFM/iamMrN4OxM5c
DslqicQ8voXPjZtI9hqkKTsfY8WSHh7LQm97L6fGzWqKJtj/zWreOM/vYuoZzUVS
KcwUQvdYJCR0Fm5wYcLQ8s8JDCXsjiQxEamJoS2MYA8FSUEUuKqueICItqMOr63b
z80tNr5LjJJU2JcFacELyLTuw9M2ajzJV+I6+LAR1Wu9/Mp1mTWn0hOkqDBXki4M
B1cWxd1ojwrf9kFxrgwCs2zn2/ytzwW7ul3oeCp6Lq7VYghnrVN7dX69TFK+wwFD
PjqR669eiYwQRU0/IXk6Qg0TW9QDXlEJYVm0uitBv1IX6mzzLYsK1xjiJsVTiqBe
OERZa95OSow4OIFU4R8zzLge7oiZ5INQ8VPDMb7L2UT3L/wiRwuCRtxIJXc4/oVl
UFZ2GG82gGwzs69sNsk0VSMd7xUjABzyGs+x2kZxfGgD4PbKobAbtPbKnfxEbGvI
u6HP4OIpOLg1orI8ZKRBI16/jRyYvXNtEa2WUrw1x3Ke6l+6Op0cTHK+ocoxlXys
eOeIMQ9llsaXbO/R5mlzrDIrvjGdw2497T59YVTbkhY654E/Y1uRbWtCyavCd6qz
9KYoGQ5AwgjkiHYm1LU/sKKGjJuUU2lUoRuzyhp0YE75yIxWN//4zYPMR/pYiGLt
DoYVFVgm4qKkstf200WNi5BNvwbOPdns5nw0oDMD/oEddnplpeVpo3KuaWqe7nWo
+H08NzgJAoQG9YpejNRJHZF2ynRTk821I6zGrk57RnPzkuReGEaOoPRrzDxSaAMY
Z/kVboJqHEYFWzfKrlnkJ1qMPMwLcaY8BP2N4p+HRDKcX8SnDZXZ90l9FeCVJNai
Gmn+SrqBjzJFqxq4XzV/vEeKaouH3VOR4b2d4fqE4S3xQbQ6YjQ1X1kLy78abPS+
zn5sFGrjfs/S8wS/Z7ixB4gcr6ZRj2V62zs06P8dSi3uopU0Kf5mJ+/CfNdCGunI
b2lWz1L7oo69spDfKBbUQ+c7TAXMWoRav3pHPYg5rY560HWNmtDyMkc6b4FDXJMl
ltExGu8e1V/O2UbP/lCfDYyrKjEjkOasjg4aUYGN8V0FrrbrRCYaeNEa+P58V/c4
u+XZ/kddrG7YxwVitwQsdqoUSqwbv1L285bO5TkX/2aZCskAMl8fjv+GDTckKcwb
PI5F1dkzoOpLsp9AD6OTJBiQu6t8PdoMDtUIxWu14N9j+fecQN7kN8edPCezG3QM
75sToghWEU79u5acaL18tiVAy9gUrH60n1yFqMtgtG9Rd/9czyCH9Mdz024FwJmz
0GtAw6GthxyKBT50ZBD8h/jKkYtLg8V4mkBXR4U+YFYmsf2z6uVS9P6wIC/b3LdF
8hvHByYVmdFbZY3MNaR/RWT5rrUPYc+fK4qxpQChdhTLKDnNqXceJJblIWYCKDko
njm4Z9LXyHoytO5iwdgn3Q5Q0wpZU+LCrWLExlee1kyTyihXXJrFUkj0pO92vHbd
JtF7pCQMi2Ho4lQk4ZPZSlcZy8D1K1TdT/eAHnZxEtIifpweMf1Gs6K1DWgXdpgt
9CQIb5mzHbrtxEzsg41vwJ6sF3d5Hgtf+fk4DQGNUPlN6KUAK7g3tif+91qNfzI6
tDF2QMeQIhZTJeK5vRyULf6MrWNkkJ5E3IoweoJBpKNslkBcmx6h36y2/QiucmA3
CYWcLptRsVk7ZpYbPUDlwua7N37rl2FkgxZQ8I5LSEVQbIEfLoseb8HeAnDAR8lv
myK42qTQoNE84lWkHz4pjNKFJ+D2UQsqtD4S35J9SkhuPwPIvp5yzcgOLA/n9525
+PVWPMMAHEnhIsczQL319DMLWQpWehz9gbvIh5VgPHqeXG6aEXGptxTPqV9JH6m2
9xgDChKXJOzzjl8Z674ebR+SXviYqzWdyhC4bGfOw0IC1Xr/DNXgex9zWAIPF5tG
J+OYvM/opmJMrEoGX16Sxa/l+MHovlC+MRCw8ppN+M39dmV2hWMbWfjJ8MYfqLja
OdNEuUENI+Rns6Itsko4h+ZOu/97wJfFjRo4PBBoZe4myMA9vIgDNEUiltmQsz5j
esUjPN8/x5lzSqnypdPwoF9AeYxcDNVvO9c/EhyHxel4fxJPNmOtGQzBO9ik+rlm
AX8R1/ocetJScgb5Y91caeWOcsosYPj7GKJFDF5VkHGqd688u09CKNgLub1PrLDI
WkaDBCqVj/oB7FU9UlF/eg37m+3DvRv6U00QdHxjvXW6DWcdUaFP1G0MYWLQODKH
2DJKA+oD5sbFrS2yl/LQIbpqlN8hwZ0N2ZBQosZoeTeN1tzwIU8OsRDaYCrPU+kn
QEFcIlLJZDh9uQlL5N2JvKjIp8MoWYOiCTxjyLYzmZtsM+t6Co5QG2f6irF2014H
N3CdJ64LsnCKpxIFnwxa7KhMpXveW1gZ9uSt4q24lhOIxQjpW0F+kPst5fnhMZ8O
KwviSn7rLb3wgc0vGlVrMg1wo9L2b8oX/p8zkzRulsERswtTbfBkVvdBKLpLM/Nl
jivqugLd5+dji+JylY7geq6bKOP4b1Dlu9xTAigvN8QBKz6eBNmKIzZd15gKmYH4
nJgms/n30e8hYINlOmAOX8gusUrB4z18kUKuZaZpBItvYJgOu4/0zm83+4J42bSL
Gy+w/DPsDeF9I0BF7/vJwx7SqFXrs1DVBGi6L7JEYOtWHm1Fw54sCM6xPUDsHye7
EAw8RmOT6cHxyTRI3jQkoCSgJhUO/tR8l7MYssL9iSNNCne208pu8BkuWKpQtfeM
0VWuGYdgaJyWYHFK0i0gRSzUA2G6lrNBpf1EhCs+H1sqKJ2kKBjDViopt7/QohjP
Eor0G2l/XuUxMVs11nh0imYtCtdjexI1WqtNPFxu5fTg4Lv+W9XWZ5DZjCVoCkOQ
3kvJPmmlOpRYILca5+2LOygHj71Zu+6V9CWgNY4cJ0H9yLGguViR4Ew6xgfCfjn6
Ya9nEudOCz/dubJd2kOJ95ozBfPU6yGmenuhhovE6kmYkfLpjpKh4PQlFsWz0cYr
IYylhwFx5NiedIEChWuo74RffuNWao7OA+3uAxltJQS8ApBnBS2KQOlBK3QbsDrh
kXk2zzX/FBE1aZNh028+diQhTKzWxJxrQlt/8MORYnpxr02lCbGriBq+XY236+e2
mCIhPsiW/dvzRhEhgdFSYKVwHvGPAWaLX0EOdYE4ZHSX6rG99dEKSu+muImYfBOf
/HpFhn2hsEVnubvGilcnLmZRB9q3I+RMx0dy0ICjv/T7YPyTepxFar6MtUUnLJFS
FzlOql0Nhwe3AYQrjz1DwvfcQ51mGRAGvy9qYfIesE72dysR2KIEvqhDKDDAZTcp
A/1E58Yj8b+Ye3v20rOauT4X/vpMnkKjYJ5vC1v6U1UbPpJXg6WJD6csJfQ77jUy
2g/qMocWck8Oue/i+7jpybK3R900vgBLXRcev/I+ccin/whHMTqfy3+O/d/VuLSH
bAx1I99rN10NgbCrACs+HXsz8OUyQx8IcNunRrJtYBaDMz+o3O4GIAZKOAJFpzDK
AJowJpvY6XAU7VCQ4S+f5dZ1hlLhdSGyR+LIsHs0tcDw9mVjb7fRDukKgETYRDk+
SznlJWmYkHOsrLzgdhz7sChw7xD73RvjKMON8NSU4A7glP4kdXQxyNMqqKCA480k
g6pxv8xh1zoboWNpk67QVET+r5Ess9w/MVf8YGxDCFvveuGTb+zLQayYWe99Jv0T
pCELDtiAQCnhw0n680orSS2nkAaVuARecPsGQxxjOyIQsoGNf1KyTtxxlGY/eRoa
IfyGVqHGChX9JVs52qlXWX3vcHYQvQHHi5Kl2FeulwBgcZ13QvVUONlnhtPrvhmm
MWS96jOsenwxGUlXwTu+f+OC3Q9Q60ttcnPE/9b8H74vnfSZJrpgiBGAp6iSNdVN
2kcdANY5c9sZiHRRSgGAqqnImgEMyLnXtLnQb6FE3sqOrNUuktNMMcXTBla7pZWq
ARFte2XskqERg4iDWfu35QLNMdiWlhH5HbFVYcHcHqGIrXBUZRwSVCk35A9/0bnU
e6Nq3J4AApi/57uWQlrYbCUCLTozQunuigWg2PoYNGjL+ODGesdPAXvfaF2KTGwU
yz1sxpeLKK0ccM/SSr7iwkgGDj8pnD6quqcKPRowdyaYG6h3dbNuU7Xqw2d5kfBc
1pCnhglSVynL3gTUPGgzNhQzWi1GpWFIl2HnYRhjR5/NNzs0munADefEtfElmyOp
NBqmbVEsuqn/CdaYR/9/BH7c5rttWFiyOadi9pqTjVVPM82EhjHNbUfJCtMBjAvP
r1vOeL6l0vD2byUQHbtb3dKY+xp2+4R+h2S/Q3BAQ4s+K3TO0cRuJpOtr+UPd1I+
IkKxNmn7Ep8WcQzto+y73ZMgf3pSn7BdB0sKs/9ddwSqTyRGjjpaZS1e1VP8Iu0Z
8iEFbBSH0UGJ6zvc56veM6qs53n1VFecU/SKY40agvkMdciZuyP4usGHLtIs9xoB
gYAwEbWe8hMX0OgcG5nKIGvFI8bBrYpJd/paZLUsXAvK9f4wd4ItfkdvDm3QTFMB
wz4t+uUa8/2Q9bBeaietgaYVh55UzttElj9JXuXa8nhaEMuWBDuO8ilW8l/5Ih0u
untybl9sDbF6Ey5oDH1l3DNjbjLk14XyKrMDCfDc7+oz1d1KjQnuM0ELuW6pt0za
wJ5CITDQb5CdTLhSLgIKLPZugrdxJL58lmmvQ+os1szJdTyDVWlCPQAxtRPmloLX
0AFdwdyYMTn0rQKai4CjYKP2eSYFTmYo9ZEUGDrbNSjbxaEjuMoAE9dVlfHj9Ld1
ITv+RAXaloR7URAoEOFMA0lbknYcwjd5K5T95w0KMATKM8T0PkhLub1qJJyEk1jm
24FLvngkSExclEjtmZsebRVMOe8mAS0Rq3R1jeYK5XjWTSnM2ZttiJskyDdbKiu1
UIDWvL99rH/4+4aKy/StU+8NCMCyeg9Ij4rnezdN1aM3BJuM+Qrg0/5bh/yy8mlz
fbGecmxPslhv7jPCfoyqHCO+mrI1QAT59DX1SKiBCX9uylw3Puic9bnJ2g5w8Oeu
KM2G+P5bnGQpjZByHOpymrhsy1Ixy2NC+0BgEvgkJlFDE3R/+KgoelveGI/7JNnS
BD5YIDzRif9hsi48gRuztAPf2VqEp/YrZrof+J2tGbc2zx6czTAX1JlN+5mBHl3U
LsWHqcpDSY6nMujchlIcaT/eVH/7s5Aj1Yi1YrarR+9fYd/K7wBREUXYtPU4ZXYV
zwKK3hLy6xIdEgjkubT1+hwc2sZvmYQtjmOV4tXq/0K5XTLnA05NOQun7b2TncM8
WTFEsG/r4n12jrHVYDay1hcEFimxzsLkIFFMvAYR15Xb5zZn8pL/wn6kmcf46CkA
clG7dzBw6rF8lAf6BFs/LqaNFkzXCvdzqqzJHjs7BVfItqLCwAFfxTsD986NJJkV
/jdqL/0XpsKZcppeLYTbCCC+zUqONCB0Qj3zean7DmexDAqLqh/uhsoF81/GZLjM
soPRvb0UGk86C4CNIsg0o2PHeHCJqvHSdEVOJLau7cWPnGPK3Ue8pUdvjZWt3N2k
bhy/hvQuaQvPT2LlvXUeu8P2QymmGI3Wl25n8S8En4IsSY9fH0QG0zp5lGcw+pkY
qLdLfOmUwtg7cA81w6i/qnTZid677OuLuIkKEBq0cflPt3yzzjbAnNuhJcLRDJm8
rUWqgaXU18zrrEHiE2pdMofzOZLKMyDps/RoNcsqztCiD9p43FLoh/9IUR41fruT
MFxCO3DRVnL5a1FjW3VPkueyLMqoXndNLdrdf1fWfQkWBsCASxc30xD8PeytB2nM
aiRvQIRUolOXTyduk+ed+yscFfVL5HDhkp8ER/Tmao98Z+q2JEkBo5k0231DrsZo
BiHUINHJS+X3GfM/V2IOjsjVk/8tWp1R77drhzDSZluN4rXZdc4UgkNQSSGGFpNZ
PgqBao8qkyd2Zd3WN3SlfLtSxIT5kwTrVlscJi57ZMAnwWm2f3gbIE16cPE07ROf
7G98LYIymbKYLDZTgKGu/cDgxDxXWMpO4Q2JGao2GbY7GbLYTW4EtqhNocFcSTnB
ZC/Kk8fZyJMywwUGOYFNgPy9jeFH4KdNWJ4h9yt52La6N1hLl6ZXdbqm7WjWb6sN
fG2kMRSN1nM90ff1BwbT0oOYg5UNWhae+/2HoSfZHGwmDSynO7rDF3+s1Bzr6zT8
7n/iITuaxfUOEHDMjbvtvLTpG1weiRlWuqa7B5Q815Vs/mu/usnmxm6Z9+UmJjtw
CEsQhTslSDM45PZeh6FtYGatO6hGg+OzXIHg5j2FjLElpGms1/fU2nf14Dh57KXm
e5UjZtIVKdSSROK0BkSILs8EJIdb4lPZA/urq69JBQwcXftoJRX+eKyWVYy/AdTi
0l7gkuFI+rJiJskNstrBzzuqLNcc+voFbfRHx9LqQtpGIFbZYnWuAdRHGC9G8qeZ
IFVwYiDc6rXXT0SiLEXsyBZ3e7hZjvXAmQgDv/8VYiHdgALQHAyVLL3/Gb3hPGuc
IzWB7z8bDEmyQmW4gSFrYL2K/Lp7UpOsqIVhPGTev4j3UDPaV7pC2SqLRSOX5fOH
F0vFa8zXtwHhiWYcS/KBmzVWYqce9q4o3GVY00nXY5lhz9y+IoMjUFPBQXRMaGur
upCsHHjmgF1osZtzHbY5nfvYegw24yzAOmkwAuUJCqb1OECtAPznzHjidrHjMFfi
3jxNgy4Q26Pg5cQXndGvQJ59SwXYfoGtyNK8fYwCa9hG8EioOww5PtbHa62OwYi0
06ruFXYMCy1A+D7BYsLkZ57vzA/Q79Thlw5uXCX7s70mXseenL7RGRixwqkn6Gqd
Osc8NgfUaUnPoLxx/3bOPB9xvd1eshVLZv0/a1z7uBifxemCPQ1f7RFso2ShyUjo
ncMt2lcOzM+ME9I46+xAkmfKnl/5gOFNe/fNhfFn9KYEZFsC7I8hLfzqdOAcOiSf
Eo56FnRpkb714AE09b/w+JUjZTno6MfczEDGLHRsEZcNPtmRQkItRxnMj7LcD2IQ
OjgTnu9B73xGCzJVnZAF3jbzifY4iyfVAwuuVfgC9ftb/TFsnYLkUF1A61JxN5E1
SvoXykB6ByGi1BWw8yxeJCRSi9RdAZWzt+dmOjNB7Vo0KrGIMpymNWF3oiDyr223
4rNxgtXGzxNcWLQ752PtbWHEJI8Fw4SDXDKSB2vCl+U3nc4quie457d39tgToFlf
NWdGY5h0iZb7e9faaN4e9s21+Atqdmt4X1FksTm1mpoSIpS6CtnTwSMH3bWaBAh8
ygEhS/vg9TnEib4CT3Za63QKw0XIhvyFx2vZ48ZfFFvVKH3xlkw/WxcTJCMQdBzT
1uBiKgQbHeSSsC/QXzelZG1C0KpodT/T2WJ2RSxCdjclbFFask0fD7Vsq4qzMPLM
3emgMvywUPnR+h8CFJGwQVWAb8A+BSbjeSHpNPV5izFnHrlbZV11soHhl9NDJ4LN
xnSoXyGi2/F9z3l2yyuRybbrR6HWykfcis8L90Mq5y9GcsBD14zPcMpYqhjzMdTM
ElAgWHugUmEeFn65PmS0aDayhbciJyDFUg35X/pNv1kptDa9O3VhBDj/vUxlWWXT
S0JXDIpJWBCExD1z3+UaO+1K0pq87hT/7sj2duYBlRMNE+MpJ3s+KFFPWVwO78pC
zCbhWgDUPMPzZdF+etVcMuooDPN24o3zqdc6d8L3P0tUKBHIkWO5DeIecv3suBhk
MxGplQlcvg+F1+/VgTxkb7WEMFvLx3HQEQiGRUWMtckMhQp84M6s+5CbJ9ojyLnR
3DUnyUommfxpQ+IbhOs6FUx8AJd+khIgvhDsMpfgjepq+a7cIbqItJmEuR2UOJy/
MkX8Ba9/C3t2oGIUKhrKBUGPnQzGrrQTW81B27XXuYbC2qOyGYZ8ECX9WQloPE0I
zeAgsdqanen9Y19yIUWAxPGRA6wYahPwFpGt+bPZWLrqEDfAV1+td6NSaVl+gU14
W7/VbMMOUi0nw1m+mkJmTHYzWx4Clrc/YRDUfXRtGOS8YrsiCP6600ixhfFzj4uz
/etTpb2zGSubkvQjInpoQmdYHN3eLuzbfp2AuyuSigEZiHbW18b3bHReksA1qnSA
1Hq5/MNl4M035yxYA5J0FWqlbhkI9TIaD/FrWis/6FpriueRH0Mm8a2CfXoHsCmy
l40LrIg2x8aJAgF8Q75qca8P855RHNLEmNzyC5LgCYUaErhGqEuweuW5vJVeyz9g
+feJ9OxWgkMjnRUFdS3tKsP+eUmBYyt37hUilBb4e6B+FjR0lm7G4dL1QMgB6/Aa
d4yGGMXxtCUwEkuSIXmZipCSeMTQyX6Pz5RrCXAsWmP7bkI0s2f07stpee2ZyH9i
gzNZPv60FzJIYpjzZC3Sb169nCkct6Dy9e2FGqConIrJGZV0ZLpsqzVDs0Wq+XV1
gBAvObO2uNTm7gwI5Wrf4agcSqZLOeZAJ8Vb4VxKnBPsEgsphw1deMNBsdddskbE
WYjmqZ6ZsfJEALIOIXOJvKKgJlBZxGsLxusetPnDfugEs5/Iypvi9trsNOHW6nMS
HwXHpNS4BxI1bDq6PgwnIUfI5QEEVBGSnQDgSjf/SKHCVSXw+nVuCAGRM6uanhG8
xbgRncH1XpGC2jMzbgHIjySgppzDY87PqCHXDqVlF+YVOxPlA1vMso55U1XuGn79
Qbno/Z412nZWf+qrewaPSq6as6CcBOx39RqGc0/hFQfMKPD6WzHx1B846W5ZrXaR
yD3BN5Sm/EkDdTX7GYJRHV4tUOYdToTo3822/F1kyCsfDK42IpkI22iLshpOoFsb
EmietPFnEbkKtx2m30zTX3jMpa/N2nQ1lOaHceiSsHrKC6+qF5Vx4L1N2vrQP+w4
S62U03+s8KbWTFyMAjRErWKZkhXq3rCimYz9j/+dL3yY88r9GBapW7WRj/vHYX3Z
+JE/Xyy1gXGlv2IX68bCZa2nnY4YRfycrn6hiu5Or9F4XYZIYOLTN502etsjE6mC
pjIYUi/tiX8J0+y0eexWJ5nj92in77T7ruTdWedZHBkZ+UodlW6JXZoTylt+CR9d
gGrZKEatRq2imIPsvgxMMPH13DTcMuEiiDFitJftniyXjG3M8JM5JomNqiZ3NOTV
qfkb73X+pBqExQKbfq30frsCrMbqpKgW6fP5AlZKTzMJwka9VUqCCW6e57BWiz0d
xLsztQc6HWLcylSw6pLv8o3TUGKGTZ0PUC8FyByIsRM3GNDV7Mrgs98ABi9+/tbF
g7hAhCF4NgLjzmNbRW7IXZA1YWQu1QrsTWP015KW4eODo1tCUJ3K8YxSn/IZdLvu
BBlpHoa3D2fuLQ8yDxDX6W/TDudhYuasGKKoomIlpUFknzlaCr2GgHPg7lezlQKs
X0FpPxHme8Lm9lqBA0Kwp4Yo9ePFYrPHwZcgVTEEBJ+O7pGfpFiY688ZzMkupeOz
jD1eWkvm3Xjg/3q5qg9d1aZBA2Rv+aV/WgyLOxX0LhUBfK5/bI1tAv/evHcYeMOu
s24mkKw8chNoH8OtiDA9F9hGzhoLaPWgVIAJs76Om7wVBSdLYLcZRZ3rmNDhAGpw
hRjiF8bhPTnwhmd5pjTf4ARBhelIX6jTo0Tbs4kJ97c+Xi8UZWnRASlAU6Zpq/J4
xXCi/8+DXT1mKRxszowsaej+B0lsZuNqGqs2oqRrc86h5LO1rdVtJ4CUYkBW9Gck
bC5HUGyvN1zGSwy1JvMiY9kHhQrJeqHdkG7jDyCQUAO3kPlNUY9je0rxIT/eyBv6
6cV7TJsOywmSDKi8fHcmMn0gQfuOn9nA1LEx/tZ1jUxPHKyvBXz+vqNtAfYJI7Ir
40FYmW7iKvVNJuEZ1UUmp1F+viW31quGufUkVuaQLqFz41uKA/HZtK6eJmXmuYXd
/rrZ4Ozh8GuNxDPmPbq9nlpVIxz+CuOTrjt52Z+Tu/6z/WvzHmqpOxshUPBB0iGl
QmvMHoo8C+IdNMJ+1yQmOuXas7aOZrZ00whaARaVkCIOMlbwupv56nvybd0hGGNr
WAaI1pRtkEo8QqvTf3VBh0ZY4M6lfNak0q9G2recn6zJ0CtX174eQQhLxoUzFme3
dWBRU6tfD1qmnhXtKFHxOae1sBSJgznVtBloIaOnXdg7Vpobaw+ntgxlj93Ok/8X
4GrCr1zPPdjC3zAZcPrU5iKroQN7n7QdSc3GdVGEOody6489wuNe4LmETyd8TPRa
XSxx0Za1zFTQ6LUU5bgVUwvF2g2s1ERU1HbHdw8/gxHKvUaSnctXA210erBb8Y/6
Aid9Ouphhde/C9DivRtBR0728syTeQ9MtuujEEAWaH77F9heEqyp+7gRXqPULt/M
X+CbEOUg9GaZCfAH+2NG00+Uex0g9wM0l4K8FGF99MTQmNsQKtzccDH9ngMIElBr
T9BMTrv/AVzH3lOcHt+rCfaiiDRJPf4busTJnYEvKq4zEKbbLLfdHmkMakAOequF
Qw3IybeAxbsJ/2Q+kMNWvGXTiKWrojw8Lf0kr914b8t2sxPFTU5/yGlXnmHzw9iJ
sxWemnN0uKYCJiOJukVVsHCYVr+XD22v5Mp36uG4wZbLBSBItnORNhwXDBKdPPnK
rtta7iQhCo1zVWsbmy3P+zhvSXEqJ1xJKZ8Pn4iAxhWZj6PmheWyx+XcEMYUMB16
Brp/+Xf8X23sYLJiQm8WW48ciovOxPfT2/feHxZ7ZUfkgM4wH2TYNkjoJ9oRzcfa
ZtNNdX7T35ZU89VxFr+pcuFrNrcof7wzOptb0lMc5ZwPpnDHdL0gB4tVbzlmMCke
69sJ2G3dpk3yjI/fbnAnFmKi/55ZE1F/z5s2Eaz9q8o4miU3RLVJS+ELk8ompZR4
xgAZHMTx1HKsDJH9p2ZBIVi/AWh7Mfw7Xv5Gs3/tbVdvqz2qJssON3EBMyVAEfWc
PZPeGj0QL5OJZNFmTPOvEZ8zEdjMuyCKMvF3PeBYxNUGI8Q6hpStppBebiAfWCTv
U739IKTpqpiZfcFKAVvCTJzlg14uuLWM/RG1OWbUxqdNjmOrYaGEskmSd4g7mU1j
iJsmYSQFNbfj9F2EIMXv960HUFYRLIAsVk2uyUL9rQMl9sLTXVhMBFDgXgXeUvq8
azKmGwlCsknd8UXBnRPxn38/QpvM4XVpa7HkaFKixB6dK+VLF56GcvBD/4Bb07wr
aZh8K7d1OBBeYBqCWOKqmet3CXjM5bWCMu1mt+oDHYPHIkRL9dD12Xu75NmA06Yz
InIFoNvXeZ3z6JDj8BUg0jdfmNGNCeUxZIcUb/8/yjGYBzs7ZugQzSaGTPRj2llo
HEJQizbGyJIu/V2QqJfyS3a1hceMKWx5CCwbHlOnYROYzE082O7Pbis8fUqFDqvt
51pKfUJsrbBY4r3QR/S6q0GlEWaBSUikYcV6Kevhq50FRFmN+zTIlJVhwef9VuIf
slN7Bh6CxHchR1yarb1+r9sW/V3ppQ5GpnxMrTkFNlfAid01WhqDbQMNg/Jmh7n/
m5iZh0TcDbIMFZw0XKn4/74ZUXsfFTFURRU+YUr9F6Dm/ZjwwqM6p18PB7hhc3Bv
iMPwhnYfQlzBWKNx0LCaKcpvtpyhH5AA69PPd8YWk410GeZraMBaMRpanjiU4Vli
bK/WS/uB5OKSmYY3emWgjstH08fBhwzaBD5bWR7ucGzmuq/ZsQtXH5V1AIXkIJez
csx8LBs/b3qp4wllN8CqvBgwJJZWcFsPH2GC4pmo0Rx2yAj9WBd4/7tur2KXc3/Q
DnL0FA9Moc/UIv4uAFoG7nhzx8yv8PDJy+2VcUp7r1YKH1VzpL4QmIqkCPJURefb
kfHrhXuKE5EmYRZwatTPbgNjKqrDeyG5Hrd9A+A8yB68lfs2B3NFm7ln9unx5pvX
FUGUYYpAnXNPoGNkOs0afNQGaiioTZRt3/47mamsgGpWr6fUK2U6s6PUu7M6nY7J
Kj+7irub8KAGhlNdfxBpTQsO/9GaAgIIMAXmKr1f51587H/kqOAN1a+0PETMN5ub
stBKxnpP0K9ZAk5P6yDVLCFlyazrh8EYcbUVj9l9b4xapu5kfMR6ajHMtnDyECEo
OU8ukIYTPDjxHd34uSgovDOy1TJZ2cSx6gg6k5Y7iMGBh5T1tOmHJytJ+1C7q2sV
B4YVsj9KFXfBcTZ1pjwIIt+pMPmBcqDrd+1aSBKzwZArvDIXEZcUGt1gXe0QN8fL
lCNigw0bNM2O+CVHmfwsETossn0MNxeDM7eVWlU9ORrO4SMkMnwzwmSWF2lQCzcK
sAjBiIhApLsCNGc0ixOsElt0WzqmKzzVcGavNVOrs18FGDByW4tzcUqQ64gVQTeZ
hmTN3zNpwBk2rAvmJwClVZasG6vh/jPcV4fZ0vYRiZ37l/ZIlEDXKaSdPCbkUpxx
ADf25LoZqf8UmUxXvHv+nVeMRgRZluKnOJKI8BUygPZvFDdGGHtmR5Fw3MpEzCiR
JXJg3sD3vzO27PCeARzu7StL+7tIY0C594ua8RyNQ4s8rjz7e6XA1erFe8bVbfWh
cmO10MlX+eZn1H5GFBOios9zeuRPv+LfNaWpNBUwqdmEvORbb+TrDWl+pLSYzhVt
BK5EVq07XfZg9mtZk+hM/VFo5ERtdhxWRhtU/VrlKZ6i8IXqsZFpVKBgiQSVWGuN
8lXBDfMtSTnE5v9gr+SU4OkNEkV+0IGa7kJXz1gktSAz06UUzPINWMz3xrJT5Klw
+ghVO60JLKmFUv7+9FNdBf1e8iLPjHI+fVvUCuQTISp0Rkse3amQS0b9zVj1Wlz8
00h9RfCpqY6rygcJOlrICZNLUb4Eq2wf5AUx17JCDqXrirxtQLiRTs/WYIkurKwj
0qYBHQo+47kvr9OrknOaeCVxpkzQeSBNrOYCXhGW+vRj4TOUVXocBCTqJqMIY3v6
VuEl11ssdHjf3zgnfPxZq/TM3iJWInegWZQYkuAvKMyDrBHKptM0OmTbcnxj86EO
N1ix9j+VjEtXktagmyIxi38vEU8bdjXiLIAg2VUbjFsrpmf6b6tO7DDoKRURvpna
biRn7NSUJOfKyyXaLCUn7hCvXi3fiUSg452oxMWCedCoe+C9NAjc3+/9BXsc/zIi
Rvcz8BN+TBX77+Hko/b5f5nYTFhUws+OXDgx/xEOkk1Xu1Ink6nhp6Kvs4RuSpDv
7pbEZSSoNe2ocDvNxT07bSiytRUV71cfKE3Id07cd3EIDE1pTas7Fo13K27fHp3B
53KzJDARfeRLcdLYxo2Ut/HI/uNSngEN5A6YBIZYfTrTUXE+17Rcajz1urDmdqF8
p6PFYmwgyDJDadRvkubHQ+WvwjcNN8mfCBngUoSMCWVsl+IZjtOvO0CLCnBCUNaJ
QxU9kI7lU1ng2tR9AJTSwLa51vmv5oiQUHbpo4eBp0D0b7RIdYpuoqvnlOWJTxE+
AvE1lOESmynWCmpmxiBg/pRehvYiWORLICZVqp1oQQs4HDCzkAO9QSwT/kWghUFm
UOnfExgCEe/ciRzVy7AiUht8OcxIz5+SujkknJ7ZU7/3CP4Nd+LlaWqAobCs5zRE
krd7FvefYoPVn6u9Ej1fiQp3JDqXzoNdexFj4SVoo9r9g+4lYyB2cpHUeh505UfS
EHsmrn36aACfURuSjB6UCv2j5xhA/AzKCABS7SGOsTSsow1Tio/nZaFOAaIVRizx
07YEpU08h9aysjBbF2XO8kYgnF8TKO8/xFrqYzgMLY6ifH44E7F0NePKVUyRHyV3
Ikxm2Fp79V4zGcCytMPwboC0qLJZ81KL6P6jqCHR96inuUx2y2FjqJnNTSoi3ygy
PlruzYiWHuapV3L2sNmPUFc5nOTOGNWoM7f8AGVQhZJRIPGImIeKR+vgOS2R+dWu
XhB1vHECGbLCRAlw750XpxFwp6tLGd6lDqcHrwdovfFRdKpks5bSkDwpCepMF2UR
0YC2BEGRru0UH2N5x7TuwM9s9DFPqD31RJXnk8eys3FuXenx6aWaM5xBjw5nHyNu
hisnDK6NTR3vBTpedC8hDgtL4kaV1lclavv8zSwFvMamwchMZQHQ3lAxze5wAGJf
9vvB4siox9S+RJWh/zBesIBlj/xT8I85k8PTgoDjKQPPlAK4b5IfaIxOF6MQcgBL
yj1TvQ4mOw3R5WvSaxQvYQju56J6Q7WaLkAPxVhf2fXiBbfPCJ7LH5qVVahYojjp
2hEfk6yZ1ADGxJBZrRX9HAOrQhF5TgxfVxgRPL8aWzrpQ/OSUQ6CZfAcGigsnjmg
zdOdZMaXRBxUoDQdf7yjGDS+y7wyto46XaE3H2pzVn4i0+S8ZA9MRApOWbH+fufa
HtiohYEMuq7H62FsAIxPIqzKPy6UArTirxahRDfTVca3Ho2IQ8LfVTnAXxSCBB6O
rYNu3l6MAH8G8KdzT55/h5s5quCf+49jhkokwbxHiSffqkqFYYGoglrNBa7o+Wxk
9MzujUum8yul0DRQXyilgi/EccofkkuLD4FxpLSpVC6ZxU+1GQjNP820woilwFLc
a4AdPuUjHNDdh+L7cq87RNl/yCJvLCPCE+NzVo8d/18PTdMi9X7Dbn+yT6I/PE2k
xxN7oqDzyfhGvfsZt+XJRWj+IbhUTy/AKJ7aNA+ePuvQmfR5BhW6jw4eltqrExgc
rQFbfO6Cbu2XxeztEyZrdEMQFrGOe48vAc4TsGTiw51YF6hH1iHJBuvrw/t6i032
a5alAJUxzbz8tcZg9o7o1UDq5aDm0n5X+r7i/IDeizAuz5LcGlK8+P++Kb0Uz+Kt
zwNRdxXMFsiSmlHbJ1Ne8PQV+9e/6DE4melMhcbURP/Y4W3JzJXCTEGwNk+HNCJA
Qmxcycb0rUwYpzJTk79C+tKKXJbGhj6zutCWPmFyT9Qws32qz0fwcZHrIudUTrA4
YNtyjk4Hudx/v0+qkeCHFt4hYpEwpN/eap+krWNtDY+WglmUgsqnTekayDABGAs+
5mYxOxlxTWE72VkMeIYtkEo7J1i0RrT7P+pZXoZy36BdQeDF33u3E2Q6cYSZLg6C
g7XzfcBK3bWb3gmTXIB0RXI33BHqHHPlKWMSfSkK4DlkcAn5lnndmfpcbIQSvAQb
I6EtYJEhl+3yNLypls2gN1XOQL0GWKiyydxlSSMVUS17TzLoi18RyeX6sJtGnLzJ
3ZOVXU+X+rgYm7RmgOvaLYb4kFfE2ZKuUS8Odma+2798Az2FcGPAmm07cHBNAtKS
+8O96ZKcK0XKvNvEJMALgPl5OQhfFX1Sv+Y25iA1P6cAIM57ph5ysQEMTKG2xwcd
98r84L3pT+XkzQMvNnOnuczlEJXv68g4kbve/bLbExnVPak2GllCmww4dMK9leQf
dLu5OZA9XA9Wn1EH+rH4H9u2M5702oKNJPs4e9jfoA/ssxGFftO6iSOfZVWIcg84
ofpgbZ1HzD9ywFxibCQSyOiXTycC8+AcMDmKQeTpoTJcAUV61FRsb1UVUspyi0ba
BaOB8meYozidRLhuvZYp20q75ZA3R3IfdrjJBuagk+ypMo78n5a+5kUZOLf7lD5N
xKSiXtJKZZ0oTlVrcZbASJlZc6rDQ27CpK1jIafSqwIEJxRZeB0aJnNAKRe92buk
S5LCV1yi860NzkOKe6AjqAhnjSJznOrjrW/ZOprDR9BA1eOUpz46cshS+Jf1Lh2H
D+VnyGnwD3IE+Spq0xWFyEj0gtABxL8Z9Mo4/uDGhVILDx710+MR2cmXzPDbzui5
PYXt/htfYGbemX/XwnAla8c0ev59k9uqw0XcrKX3lmtzwxn/vb92anh4uwZbgsIV
8FWknsivIZXx4ciQa0uNJIYcAxd/9CFiHDevztWi8D7FhvQ7wPrg5FQvlCp4lkMk
Ed+U6frjcbzChWnVDUIEQ5DEiLbe6vEbZWXA8tJPmwjWQKpnr31IojxZhGF5EWCv
djF+RR8y7e/QpYnFhNIg32+A91UYTLmWCrUQMZpDCm/y7Q0ZHILnnp9Spc/nSf9d
IsMiAam7t94p0ctNwZXBUScYnZwreaAruYxQ18EXobEwELEfXY6x7ydSdVBViAcJ
NF0fVlRluryhIZTJZjn5+imMFTXYUcS7Yav4C7aQJe+KKwnFedVMRu4V4KphtiTX
2feBLSodKIoqLCqJEWKCohOR0hhaKcQqrgBX4LAuLrKJestjtJKh7pGl1Ea8SOe7
VbItRBI2TGwHlzoVSmtcxyGoDgolqb93lyxTkPfMiwBc1wnyB4It7V6vi5YmjBwn
dNFqmrfcZtdfnlIZZCQiqZtaH5mHP0D4HKlJrNnCHVrdMiWIFcRUc9si/nahd3nl
4gkP+D1xAvYPNWTHz0PCsnsCHBk2MPfHazcU8KUIK2ERJtJIuiiPSPQ1Bq0DoG9z
sldNMFGU0yOeUjyy6FnX/o8GGL0S1hRD9vBRJVcGoFsPVYahkfaYRwX+8M4uxFdE
gyMZFVazPvTwpAf8JMUIvya8sFn1nrcHXSCpsivVXvfBgEcmcCkY/V0hloStTxps
ydZMt4VLI9KZy6LXF9vKjirAY11nR/C9576GNYYWI37s7aeOoAVJc1xQQGLwOfop
6CazJU7MDgaWqZnUiKlhSXwC3HQoCmXtug9RaHO96Mu02mnQJmW4tpG9ROKn6DGj
L1ByUYYwfCAFaMl2uzMOCnSc8A21/8L8s+n/d6qt3rT/ca6mrBYCGH1bklmMy83L
F5UsxgtJnPicfeeCpC1nf2D0Ogk+L8Qw/yh+3iIG7wePJU2WxA4g5/+S3DhPmM5s
JeFIs6lCr/Eu8gxB7vu7GnA4uVWPXUwm8ScRG/AlLYjxr6CLdgSVrK5uXUL3dnbs
hwA7KmL+ZAo5z0ac9ApdXLhNxeIwwGBTESJqv/T6yiDwDYEQO7ApgCOn4xmErSjn
tEcWJoLx45AiP8LWyxftEtIpQAt6trO/mxWEXrc73eBaf84N/I2nnY+/HGoZP55H
96dM2jFBjAsKItHpcKea85FcjO/4v5Dhwn6axT6cR+xxVeAO10GzP7agWO78/p6Y
B1A8vTUlDD0AjGkoy+xC1tO+dQzwVaxkelix0Qqifi3LmyWsX4uD1mBX3mdbl6C8
9D4hhLj0HnMwHRN0Bhf6GYhUt84Z9RcIg9/77jyv3aziVWuDFP3IW2o2laIOVv2B
YnOOoyHyUZZUnycpJrgsca49rXegwFMG3lFCveYt5oqIxmbSUkFb/UeUd8q80zeH
P4I7J8u6iByYeIbBe8rl6YxoE2x5uXgCxb8wj2gc3LQTs5I1lBnSz/qZKl8iNZ5G
dgBaGQ1Em4Og+GPFN79yeQvw1yC3XfZBBaldF4Hl4N7FlIi43tmJMbNoUCGmPTBL
HH30seP6CE1+UkUF3IgvlCsGCLN9tROeMYpjOKwo6RbVEWOxPT2txuZ2XN1TRPMk
Gq7fkQDRNcXyYJeTuYnalt3ipHI9ypD3vs7NFCW6KUNbTwV+/VpMl23Y8sj+knuM
X6zkhrKOb4nRnCgUwAGf7gL5EXW988QnZQDnj0428pjL9NHxKJN5SKRP68QU8HTN
xT0s1fSgG+QuvPMqC35kCkT3XMfeCzHos+g1jS87mXxbNPNpvKeZyXosUhEaoWXL
3GeqSpnmafWOricKftL+65kyglUekvsCpJ3FLatqkQpzeW8n+2Iy754K5jBXTXmL
JoNK6zTvD3hIqK4zl8N9ynXxRTUnmz3dqaRT/ljnEjUY7+H5V5/PztAH10KIk5eP
hN73DWLim4RHbr7rkQP479s9S7YcHeGEL7ahPQ4Pfk4t4lMSI1+BgvEh9mn2HSg1
UhYowyain8v7kwOt+pB5eNec6+6cJEOsBgS8prnlwkWecnwui2FCcskfs142+Z7H
j8E0LWuO596I0JOOhQeSPNTbhQMw261rUEro/g5e+SGMUvurZluVdeQUWo/RM89O
6ZoeU7JvVhwjNn6zofTtrYk55h8qLOCA1+2KHWkY1NUVQFXuCWFMa3ZxpQKpQreO
vvcbBQjJD73b1Q5LkcTuqU0eqrAiiYZWKDc8oM/3i4c8rJk1RuA5Lo4pzrBW6jSg
ETVY6MLmTzKUsnjUP+R7+GCL/dM1JF8jDSPe/ZpeKS61DqiHIMKiQSe5yBeXHquw
kjCUHatSkzrPEN8fAs2U4h7LimykpN2zyTtiLpmnsp3HFQC+EjlZZitw/jpVSVPy
KG1JMc6tZXlnhfN0w97ALw/vJ6n+Ks96IQnK227IGQIymBW7hPywx9eK36jXD3Ha
LkZU8xwhZgKxrPWlQHi2MI8UFb0dGLkvnKXezUfB4CyYuCJEnebk7SKWWzm5QujO
7t1pdZgivL/PHKKa7B57XEIdURvY919kiLqnU5pddnQZa5CN6cuNjwSy6usQ/Q+D
ZTvTNGvcE5kkmTkYE0HEVAEZhqx68xb2rBCDK8flEIllen1LFPU5bdU9S4kvwgya
pCwHchfBMb9o/leNEsQI8vdEz7mrdsG++CcoHE0YUYVB1ZzeNRbj1y9hqUNeNaGB
BKWb0bTTiD3ndBZjBYo2mZg/Wsh1KAO5cya3nufnX+mEYpQgz58fpZvrU3VjpYH9
YHyXvnsVr80/9Pwrc8ttPKvmHjPIc2UjOT8aOwTo5uXUo04C5Z98G8l2tS6lTKfR
idqux28Z2xN6KQo+iWdJBK6xl2oPGDangEy185pCicWxsz7xOeYb5H+P0By+9BfA
R2kB0BxUUQdgUPwEJoMdDWSBXC6/bJd5QaQWlXZZeV4/aWwVXXYQGYvrafGxTrat
jgV+ikuDPW7HnMtz1lh2tz31nUB3eriUt2Yyt+RwRUQBwCVuT12aI25g/81HXjNa
JGq0yECCDFQ39D7EKH2yDHBw7VXDZi8em/r2bDz8KAtf+/r7Rzu52g+AqDTGIsWu
1g1E/Y/dwO8gaa2xyMkGfT6HlKYfSOqVJoQAvVSabF5/YMdyxefELup3a1rFRFl9
pOCSBReufnjUs0vgNBMvGtLSENLMEsH9RnC1vu6AlI+ClhI2b4CEUsrlOe2QwcmH
7ny5gYFXyPX3+Fd4QzJ0mScZHXO8JPwRlWS53UnO3NO6qms2mnzpVleLI7fIts8O
1W/GWoTa0d9jZi7CXgM5U9rOGuVrsER6JJJQk2vjWws4UxhXwRmyGqGUs8EQhiSV
zKx2KE8BgXfVi0LzI+Wwo4/OJBFs8sT8pj9mkQS5+GsyWZhuMwU/ez/B8DOG+Ces
HtZEDgIX/jJnvj14AvtpNMktTeVUIWQqgvQhGOrGSwNj2shCNsC3p718XRJacUvw
ZiKDRMU29ccx5nv2J6zsRXXGXeRieWe85tcWDXCRnUdtnIL4OxWXz+q2KJvO/SwS
f0n3l598pVqQhWeNiKU53Xdpvn1Cn+pJxEPv9g6gtMb9eHmFidCHhVs7pPqsDx4t
HsQ5okzkdsIHvOk4ApBsTGMdw425mZaWVYt2msM5vtPws1g5r8DrF/lvA4+ks6UI
PZm3XPTTz4ZXm+qoBl2ztTsTk5ORzJ4agJSyb0wqzfTdGkh9TlxtGNx5zZTpZjrL
+4Jjz+7w9ZNdt5WwwtbqAfAQSP/mZ8ETJQLO2YwIDhhTFvFi0CBlzPjUa0hWOyRw
6KRyiCEkPOc/P0oODBKsWT1x+0V+ZTySHOWnDVB5L3k/RjNEht+7gRp+mXODvNdK
hkqn3Y42w/yiOM4xpm2h9x/zI7drv1Q0+WXRj0F1js/3OKdVbXRPWrxtmD7fOmmU
77GTCD6vU6mGMQNAo3J+ztBducGnCqPtGBaqlzm+a6vqeRj3MIRXrkRH0Zc9Iy+R
IW3nv/bAEnZyk/WksF76LuWcEkZFkiFOX5Nr3GD+dbJ1oXap8AoVJ/Y3YBOT7nUA
VSpxJ7VmxXhC56qaGa/oNaFtsVYAkqXrZuXlcRytJte1sH7GokDUSNQ+nQvtYgpt
zvOfOpiiZjigAfy//pqFz52kg03u7uOaXqyUrAytznQixsBwPgsT/Ml+YG6Yt82K
XbuDHJlJ3r9VnlZ7Jtk1KbwGpbI92AKFgrtxRiJO9JlCA9C9d4NK8CfNAlK03krb
NRcSRitRscSQ2Ybon9ssZlzBEIznjfBl6qjYGhGQk9Pbj/hlG/7ez+yNyKl0Lz29
7KEAf833cJ6tAU+2wLcPuxkfsCOPXmIQ8uyrnSUICqYiTb6LCou4COA5UBqMeyVX
Gft/rtuAFGjwk0no9vcjEYuuzvWc3mymw0VM4Qc8sOU1DrPFwJQ54HWX+PzVAWPz
d2/fdINjMN07Pi9/fSd9pEfBBnIwdnhJUcFLlBpFjTqBRH7HOM77iZxnBmS2GtY3
eo1pmhA2SsAKfJoYICXNJitPzxhD8hQPM6RJn6jY+BWgb08nZt3z5wzsOr+NJYrX
un1pBg+MEZo/9S242B2jMnwhIEEx5ClorcWQ/uj2iv4qy3c1Xuj5IUlkKaWvAKUu
SdomWGyHx+98zSo/JpdPr2k1S2wbWL7dHkqMmz1cUdCFnCBpgCwUgkjhnh+314KF
5gQixjDsWBvuZlRuq5dONod+T9OTE4RSZu2Jg/3s2cZyP/pTxJgZNiExaDxRB3rH
qZbS85j/bZ27sBNjSZwycP+fAi4n1d3IZXz1VOscDCu8QycRy1xWWKJD7uf3/Y+6
znu/yvruYXVfAAw4hG36RJIR+fBruKdDXhHzqmv+W2L6PRahX+UBA4OR+35tJAu4
yHHdE6YpIGjAjgciEKuL1GXGo2ruc7TL4MMRm0Nz859QjraXseFcI0NsG2meypep
9MyAR5hDXUcIvlfiYwEfzvzRDjVCowLO1IWXK5sKoHPEQlh1YZKmBt4W/DmueWkN
GLKGjLTbpy+dbVMzRe54wjFqZgXlyU95kG3tCwXYxr9asbAXeYMwTtdFuvevPZPc
PB0f9KwLFWt61XeodoZgqWerc+9/WyJkRLJd9HCtGivOPh+1C7kXLbwfmXmLJ6Yo
Ff4oPWVt5spci9EjZIM03A0bNlor8S0iIpFF1YK/ce1VsG4qn4t/GLCgCNgheUPE
1fAbE8bKHfJM+aW1mnX3YC1LiEqxsJ20fLimAtB1r/w62HUZiXA6lu2s1BhI5cYh
dJJAdIE/VJGiLEUOQ+igmB+LGS3UN020tnQKrxRsuLV8tJJVxvtaPx9UmDA2LlOA
JaksUUQrBfEqTyENDS0VPK1x/VERogKYdG9rEjrsxcus00ZKxuW7S3AOSJXKNy1i
tqI0OUCL9kMI+iYYXrn03enwmD0aXJyCVZ6AmsQSuezx2AHKdePy8csj9CfmBBNv
4k1IScyArMxh1Q/PMbw3+bvmVbzdtM5DMsCwRDgI086Ac0JZTlXRZ25gozzXDJ4+
o/q7bDklhduMKJa+i4HFefqp05EwuumImDnFzqMUE9OrF5i4qZcM87ymqdTO4qCx
eU5IG8nPV76WF+YCQcckPaWPPVQohccdiCVGP6B2vnUaUxbedzb45vMtJN5LYbIZ
nsEjjfUAyFoqefv0prA/FB4neDY+9TwwdYICSMQieaFD8L0H4otYxsvA/jGkwgCk
8hzdaTP2A03fIdlGoRRVEDD6La6p6UUQvXsTnD30NfcInaZ3WgxdyysYnWWEEGiL
NKqdef4D7GNpRPUnHBxlscNMVdyTuwhn4K+OKU4livNBdMiAnTRVRhMsBpIV7vMR
S3OljyL+vxFqg3gpMouMKTOpuvySSB+RL2z/p6/X0ZSia6WfAzaObZPyv5SWQteZ
vIGQ1cwDYLCDjfLjXAoM2XiztfgGqUwrbUkzIhUEJUwN3U668CE0IPllffTwVqcl
eqU34+SoQ8bWIFPcjIpeyXdqC/75jMcd9BI9OD9xhzub5IcjBMKYvDmOhFlivEoj
fx7p5F1tdvbyZoS5wdPGUuBJ3bkdLyeEa7npRtCDWpMX32aGUief8iq8lSuQKkN+
6NiODDdyeBuA5FobksZw78RNze/OD1/kLlLZMGCrJAQfOfOpuTEfQysXl/lxk8f9
+dmqoBsyCgBh1YeYYeeew+W3ZjNLPAB9ogxI1kI6hmg7p2dR4tFymMbymdvWLZ8L
s/3KkYU5eA9yXZFQkhNxsbNvxHlAwQy8BNXVo2w+88K0vadY2OJSKDb1Cox5cw0I
+7OYhPb5h8e0tJmiut2wZFpfZ9JPgXcft2+FjBm65/nwFbzsgdy0yY2OQhivTmRX
KpOO1Mpx87YfzOdH3to/2KzuFu10zsjcf1uEzKIOteNZKyjdstmvLSOZQXeTcOn8
vdJqP9zBCt8+Gaxgr8zJH1qG4T7wN1bEGG85r17n+RN7jaUgRNg6reaSA2xrsks8
IXgr2RCmzVAbqr3II2FooHIJlQLSC12GQfngtAUTw6eEaIgSzBi6oYiXwuyjtRtA
zcmMFMTxox/XVBEkQQY4u6UEAXpl0zcSHlswljt4EsakNbnKxw7ONJgOrbJ1NnJK
WgqA7E54x47K0Nk9UQwRxFrM/rGqDeFBqlb5SxeGil7wleB3otx4IswwEG1tx5WE
+HzFSY9PkzKFnrd+WFhboGgRt9rksTChH2xuQSU6/jfx27qF77+HjfwG/qWITMhc
brOyMGg1HrFZDG/ckS/hzmc/SRtU8LhjBY1cOG5EVk5krz9xZXd6JNSqDJgtM5VX
Ac+atvGT5yRsgGU4FpumDgTBWK62GPmvY5tXXpj6Hxr6r3IfBkj3+ot9yq7Xmnb6
co54+wQ7NSWaQd6NcCFkyjx+reW4MguNDMoyCAKYAFs2xwGpJVYvp5eNj3eN4mmF
eF/bbtXAEpWSRRQXSb5ZimoqrrWJMaTYWkjHfZ2NGZ3+l2Cb2PzQFzv+VwvG50Ii
Psu0UsPuV1alCIwk/CM64DQIrO/41TZXrvScQiCJpTtGhGN6ql7dnQ0PBxH9CMFt
6uqEXQVAzkAywJcz0CSAMyynVz2uTmWW1380Zsk5Hw1Z7zD5uvswwasc5nkdcjWd
b1EItagizDlZHUv2KP1uh9bXZVKfyQnNM5xButy7o6oWydfU1/tw65vRPiEZm5DB
aXwXV+itkf+buAxYIifjq0+wBfgYopAUkr09Dh1Fm0ifTT5nihxvB76W87XXclWN
N4xu1il4kwoJvC18+KKnLuYf5TXtDaR6blWKAhd2yh8p9D9KEh+lVAnRS+CcU0Bo
NffiyvV+/MiENB9q5tvxo0+l82tdgl8jbYxSl2l420uY37DKH+1k9vWl09oAILZP
USfusWhuC9G7mD2mUDmPROjnVH2gwKM0El8MA3MLYs1asj/kY02bBtvqu57YtnEE
68ilgR0z75f2Bg8JCIlYtEa3udEZE3Ah2gHHBR2+i09NmHfMxXDOHUBHQoG+SEG1
QHBotxW1nJ3IUPIxyh+2KbSz9wL1rXOlcKlpql1EczuvDJSSiKOgn+kf6/aKF1ww
UST8JA7yn4YrUZyxqAjqHgu6M/VNWDisyuAuDj/QdXpGxWJ6ageg9TFdD+bbZOQ3
6ELOFVEFV+yBQil6yu51nr+xdmDhPtFXJU9i3CIhMT9Yb0mBh04CBSVDmaPxI1kI
iTnxiOn24lLw2I1wrEYhgjmw7nvZi/ZptdqGQDv0DkdUYDBRFpFj9HLp+mxHoTbS
XJFqqncQo7r/oqJ5VGTjwSzDCsLHv2rySIpZpRdj0NePt3cOYGS43BCF/8oZSpHM
AX0w2Ll1MJkHITu/VbepUCFB9znrQLCy5xNkv2+8TqcwurjqxicY4rm17HQ/N+UH
gKv2dvmjpuds8I3bpv8d5cf8NWV03sgl1dh0y4cFQ7xKCpF1ffcZ6J7lkFIkXTup
l3X67YpMQaitpDU00X/LPNbdSg4KaHlHzC4QyRohKX3kY2X4M0SFDfNrQsUoSkOI
S1u40gsMNKZjbwbRhjRZmzpUoM7vhmi768gvQq0pJmJj4vAmWlsxftizLBuZfhXr
ttFaxak0ASq4jldT6hHaheo7f3ZDvdc/QAzuV4JxvI7uqX6jg33HuN9TvWxnK7Zt
9brY3qh/ReW6aefVb1tsf4DZgEdWyrY4QDQ2LFxRXf9DQQfqOaR3BD25CHthd2jy
lQuHnUNZekBvzL5p0viOEkBJJusvkWHhlcZl0g4yArJBHS1WTmcyKsH09FbdfurG
8zo55Nx8zO14KPBqFTZlK9dhutXCrKduCyjPDuQWprxZGUIkOHbQKHkFNB/PHwTN
NkV3SfoP3QwOwHtWX0qsYQ39iThGB/WcjGBVmKnKfyLrOXVpMu0Ucy2oLAcNY2S5
JMov5rXYgqwRHPo4FWFDFsuiiBBqqcrIcRQ/UdlnQtFzoe3a0npD0331DUtKmfRm
a37ff+K/2p/AoSWSC6XtG4Xv19bdeksZe5+PYIBzReYyB3reQtWCVCPqGyQMqKa+
TgOJ8Uewy2QmUpn4POv9ZkabNSjaZrackae/ctsgUOc2KmKztapkzyMdGewW3nTe
R8chyefxLRF37RO0o70EcMFyB8dZEPijGKbfMkNviFWsoC0EG8uISPgHibceUhGS
WJI5GV/P+XpxOy6H3E3ESIglJMAcFzd8onFOaPy0RmYSonkjpP9vL2Fh5YxlBGMf
PrSF7GesQw2gM3F11fe64MLY5iSLxX5jdhit1fKw+gVNq7NY1nNRkP0BDHcG2jO2
c1bLhfQuY2K8B7fT/ywwb3Ia+01LbF8XStYjDDSls/JoBRiHnvzC390mukhTsGaB
aFjJrIkZjVoVwSnhyWxvQUuG5QGNOb1zGGcjWAh6Q50w9tW6mH+qouT+Od0LADvL
k+mUFVaeeRUwBqbhzWGMTW5nMheXsdfVu0YXI5hnzEz42NDlTdgYCKvFdcDVVxy5
mZ7JIdZbV4p43kZYo9FpbUofChnerf24MeXmYDQZRVXg3cA7THFruxuDXtaIB6L/
KK61YcznHBps0nkuAiyQk11qWc7qX4DgMCkepZfodewk7nwyTdyHjeiGw/zNsUVV
YC4gZPq+rL+k2JqHr4kRpWiTCkPVwL2TfN5q1RPsOkGChv2sEL/rkvfTxTBbEwfS
Ku6PrwpDKqqcTKyb4nJmwURRo29yvYOT62Tx4+qSkzpbt21W0gRKbjP+wYvBbNlJ
2k77aVPhcpfFqna2md9nqlSg4wfZTHnjhTFEjHozwOKYy1V4veBmPCTcQq5Rla+O
MJnZlSSwisji0UOl5HaOgX5SYQkiDGkdHi90rN+7QmXB8jz4j+TLpgIG5rbvPU+P
+JXaXgq2JtDY4790AH3hRIRgc+V6wxddQJ5nJcnXWCnwb5gODzJ9GzS13UKhSrox
dASva75b9J/cMd24T3xEaCtORdjB3WxAPB6RzZSVpjQoAJi6+QyCGncoLAXgxz18
Q5rTGmNAT2ZtphfPLUEdtjRJZ2ufcoAJNWSX7kb5vs8Nrr7Z1rEo2I+49kV5N25n
9O1u4KrUF2fVIgYm74jpfRuND9XHJn8QTXh9k1P3IdhVyUqFCYkUUmH10y43bwfR
YR3405lzwxKfhiA3duz3wA9WR4nn6H6rjiDzq8j1NkH+2jOdjoxcZLbnafc+mOHI
Qv96bO2vbdiHIqeW1Sa3IvKV67Dr1cyZM/1WgNB+JpHMNUMwblcPXjvSQ8b6aWtV
islNuy4PIjKt67xdvS1OgmWOa8ItmNaT5NPLX5fYfQkgvUG4KKJoZV040i+dRalT
buIkQCvX2YAnkhAZJz8E6r7Vk6E9hZgKqNr9UsiP57PhAFEaTBjBdyZAplVEKtuy
WzABLe5a1eJhnWewNiilfhhv0KwBPUoUJ5hyOnwRDkEgoC1DPoDqkIH4bXVbz4XI
MsVyzT/Jr2DMNX5VohzEKDPUUctPhl+Ibld0LIBGHHwc04SMexjL/VLaqkPXplQt
EP1/YcdtzNA7AxIw940Od04WYJIw3jc3oix8Oi59UPQlA7OIW/dGJoYKNVwaRgZY
4Swz1zgj11WQOqqpl0bbkvYmsBKPDO/YMmo95pWPdkAE+WZpx/3jfe6JXQexyorY
jFHgM6unx1BiL7nsf32qrE39NKlaNEUHQcr+pkVFGTbyukYCI4XndSUvkFoyR1cu
16b2FsiMe0upNge81uzV2EPDJJqM6Dz7FcyUx+44dOilVjkF955MMlxJylveC/8J
5qtwixjAWnqcwagVWIn/0s0paklnTjfo0r9M7bX6HThOLpBkcZZI4ozlfR7QSupe
kMCppKRPY4sh2LWlyg2leIfuu3FUyb8RNOjoveZK+x+940koC0bjcl2AMKL8d6y5
YXOFxFJpBHZz/GlBdw80ZA5SF7iPL8XN/QL+MrQvN2NPbM7kPmiXJQlralfTtBqV
3wQBY6WPPqYcn7ZASfQoLEFCg1sOlxSdhOqtMJI4kdP6cuCNp4ks6fFFl6sBsfev
ePhTBOcKTMODVX0V20+Ej/sp/S0fyvt5NNCyGzrKCUf0VD+G+r9Qkxml06tV6Bxv
FyXHLXlQkav1xBOG/XHrw+eEwatwPZ8clBQDvaKYdIJdHdPiWNqbN7l1QyOhKLxY
+e3GYj7qbXQfi62lCCjRYsCxNJdCKOuYIBJ1lfDGvDWdYNeLnuuxvbM1Xr7USTjz
xkt4m4Yu1yfR44D1NaQ13piUC+pBRqU3m5ELG93w18L330+XrszWbNswCrTndCmD
g43CzrU8lhG9yEGfEUPLCeEjgf5Aun374bLztnoo6X9y7QOGXtq+g6wNVFYhbinJ
5AFMFNUGq933ZR1zjR57s04RxCmszfEe2cHfer8aNq62+Imm1Xr1jTbXlP64ips/
rPKt3Et+7RL5X9W3CfhRQYlCdFNb56sg+j57E+Ed9o4sX0tXzcUYGl73hJ1xSh26
OFaUWzS/Av0A6Y/bk3Upm6bMZby1FToFGLDgnlNbdKn0gT9Yhx2c3jmj2fv3rB+3
3TRQ/XRM0GNInmlLgzZeXyqQ4uuzMdoWvBWc2JQ/VxFdba6hIlrKY+Y5UsHkPQ8Q
I4mWs3rbHrCmukJmVDYOgxOgp538hN3SpSpjcLJ7YohzWUlCdpMXkuwORgWYT0kf
uwtJcLeNOopryY54CXOPMVA6YFRch+frhJRR3MEXWlHY+gy9XMy1wdW7xVrhO+jS
ElQVVGCGXQtYsdzm70JepZ6aP9OcWtIYElI9+L7m4gA3U3QmgXfE/2r1v3bhbFp1
k7f+Da7NgGs3VzYcngB3XUTTdlUDJNVnheuLr5DqJ5nRFzKREzRnJCrMzXyp6VjT
06wOHfgxpanoweG/rH4oZMDdMvMS7h87FckIRfq6ljflRn5mFuT1k5Vdlo5mCHQ6
3RayjbiK3h6AHuHZBlbsJqGL5h9TYp7KHzjyPlloFpMpKhLgDB7OruquYfrgGwvO
i9hpCl3aABvdZTkCC7xd2xSoKcrtQ2HyE5IWS/izlGQ2w0DsP5pkqjpLKICQcnqA
z+5qSrd+A/730SMoQa8VnHT+SFEay+bdNz2102i2cWpCrqt2tZTNfVSkzkY7Wyiq
SpdkSNNwD65p8VbTminrxiPdD1HrLCxI04MKWr8Dnn0rfXIz4eKpKj9+ASuhi4K/
/Mynm0/5u60o3vRX3wGQla/9obAPUiMr5JDvOP2v3A0Cus1n0HWiqLXWXO6gQLs7
ajFDNxV/CbV1M9GnZcPB3r7nrrvBmoCxTdaHJ1/CGfHTnMzTGqJl82uKjcgcsVOs
iN3yJ9vpWiATHPtPZsyTooq8OFio8AhrmPisOHho0L7U16A33LRSJzwzBkI1QuFs
IZV2MJ/E5L2T1zNlw9aiP3xu4GC0i+eGuloUS/W4j1efNP2lcFYzulckSj5s2GmS
C/OWtMZ7i4WkP7+nuNqJYdJ5PCXeNv7m3+cqz/Dciu6sWIcV8QeMh/ukRmSEZvt/
aMYFVmLDBlk+Ug6HbaMSGBybzGTUGtmeTzmHVYv0LrN1ILMFCb/3d4BrE5yY0pgj
wui0+ILgoxLONiuilh+afdek0+UPxFA1rxUyHK/U6SS5aQ312GnjKqksUC4KcVmG
zhJWQTtgzE8HfA2edwOfdtSYjBOtzojH/jhI290/KGEgjEuc5GRM2pC/fiB6ljAg
GDSLU1dOH5X2pPhf0LNxCNX6riuUXlSckD+VSWudiUOk4aaudqwYG7MjGWGYNQP5
jSHu/xFVzPVRMyq2/AY1TLUvouMLNaa/MsgaIs5+2Sir8oXxGjbjqLovT5hn5tAS
/85RTioduAr77ELmc+Eeg66oEACUa+RtY7rBjPJg9RT4VqRGgYAEMGYjRiz45FX/
Pnse+lpqE2MlzkDU4XwdO/qscc7vile2+wKiOJHru7qV8cUrInXuQRvEkn+zqiVe
q6thnHYel2zz4qu7eFoLUySGIGQvkxaG37hwzCOzUXf6xbRG5LaFhpSIXRZJyQ6H
39AWwaPfsmQbAYzFTaXoemr1loG6fOOJ0HTVa4mDNWlfWxmOOLnlcZ4F4N2ZYi0w
6tTezj/j0Lv5AxvFt882MchcOxfW4/N4RxpTIqGc5Bz54ltvUMrcd2kbO7FrnF/q
8GcNbwdt5yUSjDxA9IbA2b2ZraeHBPBIuA+nu36LUybJ2MjSfaBt1YA+nMseysjZ
XBgB991JFCEy6Usvu8yTukd9EJv7ZbOH39ma/qzHMhRZhsJO6TlyK/AmJE047xlp
Kk/zitVs6no2gHXeQXfg8SqhQHXN5x9O0NdvnHpD/KcLuyMAxdkiymZ6uKt4pjax
YiTXhSlPVhcKuLMm2CYKBJ8zDo1KqcTXSNAdk4X8nurAOEWfo+ZH0qbF6sOHVmAM
cbS4Z8vEwm6UsC5n7UjO8Qe9R2QBY2eXt6XRuj83EORNPtYb52gD2z2X2MhG7n1k
pMTBifEyCi/AxPlIgYsnE3/Kt8TV0nQmDpSSr1bEx2bkV71UThGmzQ9KPTQB2NY5
HpDxGbk3NqTbbyBitvdCiFKiyHjhKFLBEMzV6l7IFJPPdBeoXST++We3R5gHfHVE
SL1rAbF5sOvWzeEE+2rtIaGH99KIoauWqxDGNn5ESXjY5ot8w6t16YrhZpucAKtb
w75PjiRWIPdr7XH8OPsnAD7XMYWPxwdHvYLAeE9YCWIlGuL+qmYS8doCspNdGq7K
N35xE6lgqqTU0PjTFvtVru8+m02NlVHcqDvy7x6EmHLJj1yoWPFT0zT2f2/IRDGJ
Ji1bQRmvPtYS9azKcn2V6BysjLNKqx8mfKhUmBRbTtlCndYkiiksS2rMfrP0+12u
ieEGs6g9ERJ0CBkCkn8VaQ6ojKnBqAjY8++Y4V+b9IYKD4lEiL/G5k1ngcZd2JmF
rr3HEldcwu5qKhR05mFlT8GoFHDxerv7rOZ94PEaSnvVjIpa9CP4ZYpkuH6WGPrN
FDvD8Xp2CTG2snogNp2W2pFdRwxRlbQmAR70kDlPSEXuSz6stcZFRNaYSRDIPIpk
bkZCzEfwel11106kqxKXlIGX8jATuhLSjiFCfwo5ko+AMMRO8VlZjpaEwzeFLuvp
eQ2jrgi2LCSsJ2ciWJC25Cr+PYyHb9o4iv4czL0ai8iWDKtxVJpMMww8IaXRALfj
CC95ONfGAfl6rHDHO48zLDMRbKEjlNwrySyVb8ds6fR4GEraTNFoaDMrfXpl/i7S
8Jjr8KYusAD+btZq+iP7/xC38YaGwuYe8mFB//TUasFTiGXapM3KDxVu7rs4sdtp
ZW2rfuwg3YU+iPBgOIf/KoHVitLy3H0sztxwyNN9D2/RZQOk+jo/+A87ENYeH/pO
/uA+YbyRV1Lyyben/K91tIBqwIq6oMDC0zN4FckPKJHGAlNrnJSJ6+T3pM/jApg/
QQ4njtBXukBbG5hXAWuG98TqNj713n2v5TD7eoMDF0JT3uGgemY+AWageFR8jNGi
1aqMDnsyfNQKr2Ut82i88IMK/08blBpkhohoTqaUT73JyspnjVtxTzHJhHrfBySV
p/EQhPIMF3Xum7RVyzlPRDkSMrYZ/KMyOI2Yn4ETEOGXwl8y2wd+X+7vw3cAK9ah
ZDAxcd9SkNRAaDA1ldPFTWHUadVEAFzIwdo3uxchdrxPHKw5yzhW1sJSftPkqZaG
e+wFMCdPKlKQMUDKDg0UWm0dlMSp35yP07Dj1DFQ2TYZiI1jx6u3JAU36fIdGKvT
lturErMrokpvjj6l1gHSpzZuEsmLVoXFtEF39bCoicwhUK1NlIHHFyygdoGQJJl4
qNVDp0lP+jZ7H9jo0MH/ROpr0MIBKaxOviMmQRa8HSu+7UYc9FeEzZ9y34aJJ0+d
nJ3AdCvx8OigFhgHhwuycnCfMHNASgZcqn5BK5O1FB9ULFE24L+r8wqcyJ6ZwD6N
zy45RcKTxQkirz2cBIXA9Fc6o6aPsWgAc8DKHL4TqI0CruElOv/CZX2JjePThpuH
vzD0sQhgTNGUZoEqcEeLW+4XnBlHDb/+vjCC1qHf4XuK07T87idNxGf3dGl1DI6Y
utjCy8ndzvAgKChLqxLa2xjRqXZWmgjLTx7fcwt9MGyp3GJZLJ6mZ2OmDjPTJhO+
gpVJ9mMWxkzdCxToV5orzA2w6zrmRe12+70z63hcUvmJpwOU1cVcsH27rIC3GY9M
UcewTeYN3bXTR5aVDbkxPTQA7Zc87Tt9zD97yNsUHvN/rH+SdTp7dkBxY44d0OzF
h2AiGl30oyKxfED6vF5Ywd5OKu7QNtpHKbFTSpyEuTujjeUzKoJhbZbnhOpLWJm8
4oA47vsZe4aMiNn344UBO41TG+4OVUyDmjlI0IPb08zPik52gFTHpjStuopWoXNV
Sy4mxy+IV9WhMdv09xV8tInuHz4sC51UfXZ15nUC6xeXlnqNLJGe/drqkJObwGh5
ziMXg0FV9RCWDJNfR8mPHL94rx+DA4yMl03x3mMEHUyROD5+zA/xf82Qxj1NWnlt
GyCB3ySiWOxgQ+u80gFwudzxEPfky1W64I6Tp234aedkB7ujFiwnJ0O5urB1QKA9
XqOv/N5prbsEF8Sg/i1SefWfSdg+FX4OeNJj9uJYZoEdTNkgFtsL4Tj1aE/fO7qP
3jLYnl6u26jbUILchk0k8u7Iexf8Pz5ieZdY2DE+hQ3pvKdP4Yrm+LCJEHPo25Za
oe3jZSPFqxMFK0FWSHrXOj0mrOZ0QrwF/OtBI/T4j4DJcgakgvtWviN7Q8zUKscp
1rH33ZubLWPmZOPe01OOuA9/qEWSVp8iUxdOJD+8vprAFEcOlfnf9g6HqvRYzXG0
CsXnhEBDivxeXmsbYQG3g0dsJpiYEnk4V+59iBv4f0xve3cPqAKdOzLdvwvT9Ywr
NpOHLTc8mxpK71jRpjIEQIPdvRd2uTV4PqTzRbYOkM1CRpCdxl8LbfxBTwTI92BD
o3Z1jofs7XO50H4TcI6YDKHDSUXXYQhrr746oLjMYkbRciGIig0EMdTUg9Xweoq3
iBy8L+RK9R73D61JIoQIVG5SpeH+MYEkai1XtzyHpTZ9Hr9rKTFuzGmlT6ApdDan
9/TkbDOaHKX4Z4Gm4N8czSKEJQD4vrj1k3+q+/B113882VksvEx7uucCX3frPdbO
i1UwWINDfa9EjGD3N4+DqANxim0mpW52xfuWpaXNQfaupBMxLnYjcWXyKFLCe2qO
3+ABufA97uDpNA77jW8yqkUZNZyLOO9rUNjZdM0TEYbwYoWIH5bjH/qbM8wH6klI
v0mUU3qN5HaxPtCJKq1crPtj4l2ZEWjNuKjug10YeyRwK6FMUH1ANEr8oas0gb8C
SDmzRufN08yamvTmUtHsaSWaEHyrnD6E2tcgR44EnbUxY3dCHxwRImBMfNrHgaP1
kZQvSQVG5PxKe9Lelst8OWIWsL9QtjuM+Em2powAKTWDpIyLNlaZ0klcJzWOhS/j
425nKaPZ/ZrhZuQSi1HJIMLjVAg/aKoCJKaMdcU9xVUV9ojuM/jGBu7ZsIw0U4l/
gXbZy3ZldRtvHPo6/gMJAgzv4w6961pDfbVZPjiN3SJQ823p0IP+74+2jLMN9IUM
HVjZsLo3Vqe/25P/TgjYwKyk0dSyviiKb38O87sYHQRI7Gl6nBu3MJn/XT2+D1UJ
n5NkB0qvhTw0tEPU3m3MIu7bOR3W2JTR9GdxmZB2u5xG5BjXsTP1E1CQAvHwvC6R
kcDw5H9Do4pSxZ8xmNuqqDog8L2m2fW+x+UBnr8/znwzPVQYkMJpxSnTnvyPXktN
Ce9UXMcfH0nSwKIIjaQ6O7ySDJWnI7DJxXgcg2MnH97+lU52fc+DI4kWZnraxKEy
1dcVQ6o+NSzQvccJTZB1hL6Bb7sFqlZYZXOcxJc45Xh6OElTRZPHnW9w6tIDXamQ
mcN5OmVaP5X8Nn+XsVnx8vS/29mA7nz57D7IjqKts4pkpLXC1+oM7qZJE14bQ31a
Ehhp7TMXBYRbN8M4UokyDWyYFqdI+cw8V93pSlCGo0rYEHhx0hAmgsgz/SSnWNnc
B1yKDuHYaekgvd/BXRp75+eyGT4bDx8HBMLRJu1nKxX6EqLVlbFxOnqdsvn47nit
uVB1ivME/mUN1AUkd/w/xhyCymUpZhhEcrGcll4mcGNRaL2G1+XZB4pv+mT75EXb
y7nt0lFbWsFVxRWtmlSPkRKFvf7+eZ0UfsO4bk0m3ty1fSe2WRY7AoUD0vCe7XvW
kec//6fiSc3vSgQntQ4bn7B8lDq9EarHAkG3mMRQ1/PIQj6zt27HRnC2ycVQfP74
yjyE5RShgjbRPH1eWnma2lrwsCvoYCKVOnHUquelfRw+KKThDfWat0cdO59zMTdY
TOFb2cW2ztWnR6DiDHrBXxTxX3DnJ244JlQF4WBU98uBqaMYs4FSeMd+Xh+jRK6f
PtuL0gK/fwI1uuSU53+2WgSN3UtMFSuCm2/3i4S8BXo31qvjRutdAAkot8uxrIQI
QBq1P5+nQl7xg0gO1NgWk/6YaaU2dcwwc7zBE3leWjKU2GNSr39F8v+GwYfX5hPN
FqdxxowwBb9R36wZEdvFmkE0XJQo+5UzblYlPE64Qe4PJ0YruauQ4kU8RFyJsKKL
vjB5elQknFLexMXUrJHoatuWK3JmY5NaC35s5P66LRx7UAMRZFCGXcK+0O/lO/wb
wqgLEPdR1wN+KKtHPjIzzGjunN+Z8Ote+XAYaOAEH/7oOs44INWH0X1lZ16SXdw6
8AjaxwBp/eRKg/B9/+LMdnSNxqC6Vtx3ux3HTuFQsJiCH9Fa/+JDDcqnEcyzLCTv
M+Qg55DOUV81aExFb+1YBZQ0riBIkRHzDVMQSpa0SuKsUGJ/fXOmbDLa/fBS3VtA
UnAiwFCUwS7JW+mwc65V6CeOe2XFBT3EKQs6T88+SzNx8OkF5CPsfZchhHMb5w7V
yO9k/sNM2EDc7MpJVG9XmP71rkWmIa50V+uEmL1GdoliRW2JUxu8698DLMXQryhf
7SHQzKEcXJ3M9YvnWl3FyvNzxOFMVSjPZy2oMuRBCuIqM3rXPZ8EiNYm9a+N1Cr6
gYt73TwdkyB7IFzK8UQTLxtwmA23hT5JW6ilhzh/frXKVgZX52eEdg/0sA4Nc0pt
6Dapen0CazOBVgzPGBFCV8YUOomKm/QrGv6oSxnRHtdnLeS+B3uBd3QzQC0uqMqa
oqWMvQfpI3cpR6OyvAqUwua4JYWW/Em4bBhr0ZdMCmnFKEpMGxisXjpTmNfHkmDP
cppMwxugZmPekFeppm3FqA6iktn05la5uXT0CCzgSLobIwUGIWoaoa2CS62br36g
wD7z45VokmGnlZr1AjiTRl5m7N27dXWhCQ3ENo4Ae4WK4/zGrrwXtwwinyliaQ/z
mYIdDnhPcFhOllpkzvuRYqfRC+3o/+SNP+R+2K2KAkS/2Ac90GEiR27IoielCIxy
QF1pxZJvqHr0NWKZy3wqH3CfnFJ0iagbGOuPN57fAJ50O1v9oxQs6MTI/3ZXUTuf
nDRKkftVPgTSQH+zKGz5kiHS5JjMxyJpSqxhSR06Bgnc65Aj04c6d4VFOWFX5RYe
xBUxIFGr/yjziLh60eKtnKzGvooLpwdJ37vBe82jf9p+zCjSSuhAZwgTOOvZ8lmB
di/Br/QrScDV6zxw2iTnvqjt/4pSiTvHQiwfKJMatI3f807HOuCNWxgEBwMhXxEI
VK5tTJ9J8PCwxwuvyFhDC4qqCRtpgiBiMwMlBBHsK5/CO0uZ7GmJD45yq53M502m
c3R5bxPJRM+QMEmdt0C5edMuNXAqLZV8vNOEPdmhAbhXE5U9yW9QgS6CN3ems9PQ
ffSuVvcmJBWqXcDPPiWX70i8EFCl7SsbgBM/QTeBCBMJu52R87Ts9Fy21NUwvwm0
fYsiSpDsQsUDayUvhiYcC5oSXUi68/PMRuCApM6XhacgXmUcEa7gDIYEH9XDgMXy
YSkkWW+4FBkt3449C1WPke+gtfiR7cQN4iqMTMy5A6FPe1fNhOSffiE/xzAWzlTp
+TCWCBtIIm5kzJHoxli5lv9G6QKPa052oAG20ygRXOJosSuWm6Jis9X4pPN6czsL
3v1Qt8f0kU9Ke5saW+QPu6ZIGxTHB9+RqC4xv/JUIW8y1hHgEX1IKt4nfFxMtsD4
69+RBv+QDnDUgKVo0qxw6SjTeWZ2E2V6YvoafHnPOpZa7TxhqidSzZeCjfW4wtN0
ayL0jwQkPBrkw5X9k/H14p30V5vdQ0eskSeQ8zk4Qtf+d1Srj2Kx701ZAfrzvPkC
whN5ceFbmIU15gOFYHclhx9e8bpMtKKrc411/SWdNlBTxeYojbkypibQcLJcXVDA
sgNAs3mAyW9ucmnLa7i3HXBnIv6Po08qlzBYwVseoHIWc16sDDQJLdfK/u4hFjvZ
aWj/NmdV5bL1V76iVBnH3a9Jxm3OW4MO/m2nWM+Hi3cqX5t5KrD+1hicgTWBiqXJ
HXnwGsC4U4YUwZ/uiPXB7w4eet9jrtaNNZySD87I1d6l9SVRpi08g0IG6sxQA/ZU
SzhcC7GwWNmZl7uXxAdcnpDFRu/7Gv/D3lGqGlXSAnEMTdQWdRcS/W1sSJ2tr82M
nc0DkBKlHv9OcSzsiicL+ABuOaHbUdEMXvTsKSCSl72AlSS4bFMZuszE3H1odbLJ
4k+oSN9Wcw0HWJA9nD1iePumVP1Ta8GhUnv58P6blEPsaClc/xn6+GcENbfuwpUV
Lt4x47lhDXUPVtvDwEvVMx015//+M7GqbLD75ClHDooV1f8lwrRwGeqBKA4DiuYv
7JwjZv7il58PxfQPdtE29h96/k207MiOxOKIuQhco3UHbcwqws6Lj0BzN+QFY+Cj
fuMpNnuysU3FxNXQWT0H3yMUC88YD+QXkDkWwd/TqVBqO/Ko8rMdhKvOEAWO3Bqp
Tj9uN6bbeoow6nIvBxWZOZMRgftcI+STrqEL5/jZVuy13PEe1zUsLv2qtQPpkoJt
MtjC4ySweMHf5AvNfvrqBdI0wrRZb1jMPNmgcTKIXUavsuesjE07+61d1St5wdeZ
dKc438hlTrpvQ9sXf56LYXREO/4vOTG2zo/Rb/XE1qTDSlJikj1YboKsuxkmhL/m
OsgqQ9q1csNw6L+xljTU6EEwWFQGAdlXlR/UOwFlCTAbu5GaCVJJ6MPeVcHYGeXX
M8wDu1tOnRvdqZsKlSOPNT+0gwuX508YmsGd1hyKTXHqAV7dFtfvkqelkdXDgP+U
QgRqlMrj/GRaVoGMNktqgu0Uo8NqicIBf4CPrpEh+A8yGfctIWSsy/p5kSwM66xo
bx95i7DKk77tIEA/S3F1u9TIRC+TUbYG5sTxbiKTsMBxeelpqNW78BTPt/BpVy1G
VBlVLR9FODejhs3u7B+vR1WZA6nVkvDdKbjF+1L44mw1KEzmla4t+eVTJ8ZNX7tf
MOeYVExoLbjSG0l1MCqotnTbHPC4zkXXpD2D/yEmhnccPFJ3yY0giur2aQ0kWy88
EXCOACFxMEWOXaX/y64JgtyGQ8FpUCR7Bx83RtMkfPbGcWG3oU0GoQIeRtqXOg9G
fOlZbInXaT5413xObQUIpxBFZChDdzEqNrmE0xtLPUi6N2IBZoBx/tLxFDhZLVil
2SkT0Dkl4WrPyBdzXNLR6vGtDJ4ROBb7g3FTB/WxSBeH5tHe+iFkD0ZBPWlzdzk4
ACCAuPfFiioeDtrSUuY5XLKcyIURdwAFZ4I8BYsXPvyW9UcDKYMkI1sQUl5vtl1I
kTvRjlOcCm8K/9f5VT/wtAJofcnCo5oThMMC4NlzBJ9RHzHmfjTdNr/rkl/ViJwt
puxwrW0iiKy9IzfGdp0eD2laOiLNWRBgPkn+BI3pn1IbP4DGE9hAFwm4Td834s9h
b0r1NF0Gmr8uoA2whI2X/SSwMS3H6gbKxfBjeFyDNUEGQdf5Ujt+XpUYv+hjPbCR
1ohOmouYo+7A8hJIiTo0nFqVLn5ao8fs6Vfdi+TVYZTHajRZTvb2uDDtVmmJ9k/5
vsLe1CcXTS3ZvdgIO/gO8oHsKfKrMAnbZDIv5xEVQrDMgmajs60WS4Fse9QGqD7x
ZiPNNmXAIQJakWugghYJa5DNzN4wbu3DFFYU9SyR5/237qcth5+WWo/UE5tJMbzY
sAj7EfCZOXI9kpg9X2K5qNbmvAk0aG6tSsqbb6OLBrmFW/8DCf/gMKX1Ymeu+ibU
0jkyvB+Td9B652MHgZ8VltGsp2+Q+Q9ZX13QDIv2M2jHS7PJ5Qx/wwcpzSSB95jq
kk9uvm6R53FebRS3+mfCeQr+dZS7AZ91qHiIJlsTBw7rrikaKRRQcQdecDOz2bol
eVj3a6LzJLeT+RsUjesiUMCoN8E6ToWNZVESWIMbawOpSRpHwGZXxNRbeVYiPKlB
ZJnjDiWdc1mHMf8kxhMeJKMng46s4gPm08Fo7Ik5AeSrc299EXK2fPrWkCPkKUmm
EOnd262T6fL3nlLIrYPoBOYz+xs5F0lQpTYnpA/UhXTOznhA/KYBqlsuXV673CmP
D0QPgkonrlQGu846WJDOd4eL57ZX/Il/QDkglfssoDJo6Ch6l43Ssz79HOPUNDxU
U3Xx9G6+9CnrMrKKduC3H4GqpqMAyivwWsgdMfcUBwTLZ8kyEvyb/2T88NHDN2XD
SeQLKsAppHHVUp8iPRdmjr5RoUayHbKOJBTmYWXYf38TsADUnyFEnMPMstWPBTZi
kzwvHIAMTD7qALKTyvILztT+4IEJE2LOYFEoVcb4YoEnVOVIRvcUYZMbB9qVmLbI
bfUG8DSmq6acG0ho+PNZDya/FhxLmgjQGF2CD7aM3Pc/AQXFF74lmDFbeki1B0FC
xAq2r5ew8M4st3fyxxXHKt44D5F5NDbWHh6EvneZcEJYwPEHboiArFJnqKsyvzu4
sXKbW1X4daAa98hnruVyeo0IBk30EiUnUSqZAP1qsNTsbFylYS3JyNCtMQJYejwH
ifri+4yYsADpb+M6W8NEbnRk/scTp+eQPD2OINiAUrXYlQpjY3qeYi5HUQB8tbRd
0TGpH0Dzbr3N/Z5DzUF9MTSt4evclQhLTkBo+8rzxpa4wMYsozginIipsaEZ/1qK
zcgpqWrhK9S1aaYxx1UCeM1yOmfuCljqPRZp5R/oWXiY31a/zQVoWQpp9D+dZDC/
uo25WsmLLStGCPlxTyWG5SijRmaXaQ5+L6Aya21mg2mBQV1bI55Zm+uJZmD5xdiX
XkyVpBfFDz8l447fYDk+4TDtgaC2QTiX+cbz+0XlFxKtgQt7ZU7PZBHPQ6inVObt
Lgk4AEbT4JAmcV5VG374HKZyjtS0c++P0emPq6iDbMR0Rk3p/Yyng3qfJTp9xTO5
DecJXkyQzfw6yTTL1ZBO9w0T1rUkVYzxztVy7FFoPBSWmRKAs0OZ+FkR0nOwQqiR
9U7vL641OByiP8Zc+g0y+0gjrcr0oCVibod/TA6MEpJmqgMxsyTkuHIA81v3hkdN
RhwjKZY9CiLzOKRxDKZlwCWuej5VLbZpvCgtSOWfAncaQRdXaI94RNuRfJNSawH3
JCzPddFar4AvgcLwtv/JAiSiRImwrSfrL00nkam9jvTgLc3uIAe1tSuXc4UO2lE4
NgQXfnjMYrEz94N+0uwkyqFdd+oT3ndV9lh4y0rlbxD+jAPXWc5l8pu2dOKSXc0T
UyG545EiK72/FC6hTP4c/0sJ6zA+kb5wnwVq3JIsF0cKXVnD8ir5NRm0ro8kgYej
x+Iu4Br8vdZgqwu/Q5OwmFpAQrWnP8+jPAdJO1zGXTODo2G3Mv9+IjVs0CoW9k+n
MIi/eXiLSSD8xcKw/d2X4KwPL/JITdnKvtFeHF0mjnfjq0JOsFILIEwUN8v5GJDz
TZOPoEY38Fg9j18W2o82wvfV90bXuZZ5hFNwyBUWBzxWleYRI5yH8JgIC8WMICFn
XOvqQoZgbzR8E9THXQJlRgRbYPk7ebWTrFO7VFp2w2wSI1qfD0v/xDgw8gTtHgjV
GYZvEPsymeVIWtKfSAL+q4WusX/fNk/DG3/JmN4SIe1rK81FeopVyZYxSXpMDfh2
aulFrsE749oDAKajuwwrBKfhZNMCcwLSt50N1xC/5YBjLB51iF5WrQc9x1PaQ6St
+Nu/vta2NuHzMENfFwYvnC26FIlPSATmratAQ13+RQ3Rw22ymHTOgm6ymbDvAQuB
VMyq1wkqFawkj0NoB/D2Jn2CLWcB9RZMuhdQqXYT49mEwmQNWKfnqdZkHy8wdOFC
HdtYdV+jvhTsgEZVl3m5uVZXcru0PH83Eg1pN0Eo7ib73xUujlq6KLpniick5X0c
s9qOstKT8iptEDtI3wRgSUtdC0AN30uX9WhoI0UeAgWqsUNwjKF6XOHpmbUgC81b
jsrsx4PprrJpIL8U5c5I7Zvki8JWa5p+qAfkx8N48ynlXPxf9TGtHcBuJcvni1WQ
Iz1NN5mn7BVm1jrMiu0mRkYtq26Ff3ZJS0vu5nfnBrSzDEFoA2v/9sJg+ZFd8XTP
JnuyKLHXnJPGxADTEZ1mgOfGID3JQWPHeWmDtnYH3zrpzulqoW+tYAbisVAbjJhn
dCXnOQgOGkpB57nwx3ZrSa5yqGseOZ7VNEU+caqfwHbHEpGLpfXR++8nAiC3VJcb
RFfBhbVzrtQImcB+V73SyarvGRdyHYpSixjzFFAhZVr+nuLyTBRsU/oOJFTsiRP2
MWsl7xFBQybQRwRtcNkEloEX19lPP8QsYwo0VW3K5Swf3vyMTeyAHUwaSKT8PYrA
ZsvYbJ6nk8ccidt3/CZIgd3fWo0U5gZcILaWS+oNIiwzTwmUHNIFjZVa4hIXYb0N
Loi1LdV+RMfEBJ9ahfEV/A2rryEIM2jXDFgLHpC1NOEkmB6/nKONs/F4pUexOkXx
dY6j/xi1/rtpB5IbhTtMhaFqd699a0N7XExaNZ3Ii1sMN9ZtZh9TnfuJei3r1ZSN
gJ2utBIMYdpVd3M/9STNmwclh6Z63BIV7SshEBGYDI0Dn/mAStXiQ+qFvMx40rM8
dkZqx5YWKsp8D9Fwi5NbWvkyhuTg/rPno0ohK8wO4uMM/Ioe8YxYrPQHXvuIupJg
ak6HObYUfi3Cl2nTZa2QXrcVnadWfj9N6SEuzAwj8bmVmtU0RXNd8K8n551vwhSI
VsrG910pCNHiP1vD67kmm2uQ9tOmoQcHlnniFWYBQcysVHbTaqBG1Nt107LcDjPd
MdRSbsBveYuDFjQ/eNJBubTVozAemQWpiMvhsh9nF7YDPiW9QBZoCGJBUtmebcc9
UMg2nBpsVm9oxLi7BvlQZuqNWNfWdAdiEbR9ZEBuSywyt5iq2+eKG75VG+ZTMGCM
1Jd0sK2ogsc6dbLXTMrKe1yz/NM4LWXbv2RoM+hnmHMrxX4Oi4zk67b+GEDepIiP
f9XhSlFeefSVb9PxPYqbeFkLf+LYKYJwjvPGSbttrUGGlF539Rmq5EKcTxAEtsi1
BkL4k/QTVQOyhGX000rto6Bfi6RhM8pp6ocRDmyHsYIW1dFYBDoMVoLV0pWxH29v
uzEAojfbww90nzl+JuUapAN1pJvT8HCRo2Y/ddbn3p0lnqdJV4nu7nzvFxnguEmd
urRGBicxNPZZZyt2JtfTq/JL0X5fwjhDXucLy98D4MAeLFi9UIPBOX0FaloPuoON
cEIthYY7DZTFov6sERO5VCBgO0a+pPMglyjLBsaGv1fVWIsxp8FTydYngwUtjBh9
eZTejjWSEYtuAuC4D7kpfj+kGNZMOeXiAelZjXFePKPrfEK2Shr/V01A6yjcalnv
0Pju6y8ebomurtoOP3DfNLJlUYLBlNCvNefQ94ytbkX4J4LAmi9baieOhB0iJZk6
sLMambBCjYFKGLsCteXip8+/67HHxN6vbiVncSqm7SdmHRAMp/8xBN58cIOw5XZ4
L3u4ajwoloG3brax7ibHj3f/BxrMhUZpWeDGRxOUwf4ZhCE0fCFXn5IiSme7W6IY
NOuYgWiVdNZ2mNsPZITopB9lBqeDwl4Axh3GcATFCDm5ZfqVLSXiPRVw3RS6YM9u
bphMvIT9h1wFM0vEbJq8C+LD6X1UmwlIlkF340IXKbvt2fPCaR8KrksrIqrpvEiv
MbI2HPVav15Swimk4cqhvHDkYadmKrLrqndZ1H3B7UfY4D+Y8HqllpDg514keI9v
qJYgXzGs+rlzbaIJnFLV6FF9NhRPL6Lz0xfAEP+zIkEbjF0v1HqjU1CBPY5OQBY+
u7xhPW6ABzZCcSZWa47aWjqyX1O9EGBfhVNkfB75LLm2Cv/UsHCFDb8DEJ3yfF/2
tcx5etdLRejYpfyH7KsXt1ePUtOTdrnM5ddBoeYOXiq9wC1ex3A66r4DIUEhOl9L
swUA3ru8cFp0tBbrjK6reNRDk07z8zQQ00RINc1GyUoY4liMD4Etqd1VBFeKwP8N
obQBG+ZqvGW4y2ucHkQDnfEFcPi0OcitWR3ldKTXL4+H6jvNAmRqSDxMmxGgqQ30
bH61a9VOBOQmM0SWAB4pibAzzHts7E4urlLigiYSroeUe5r5jduW3Iuh4duw2W9P
S9jjjf6UHQsSbl+gd0Dg2h4hu8KhAfAaVGjM4TlYMUtyIj2RRaCA/+rJfE4+mix4
IxvGL/zTH4P387DnCcp+XMyNy2DDlsXYXJ/BnSmzHTk2kgus7mJLhW3WVimg2dG+
6teB21ygWqud/w92Jjxs6t1bfTWNztHjBNNLzdwVJgq3hHgFRJBceqeRypwuqTmp
+h/i9LOH5RmJ9D7Cmzo/rf0UsnFWsEl4iv2CmpzLdbav5RnbtkQcyD5o71ThVRLz
fdbK9AV91m7DOH+uY4XC8nWNqtfqG7iE1i0QwM5uZVNodD0Ho3PRxV1gRlEjQ8gC
bJ+ndGy5rvl4E+M/no0h4uhG5xBqdlB/9yfQqhGe+cedACMHx5IL8MN/9+efbQJV
h9UgfC7FvY3CjF/Jt2y1BCYWC2vit/EpW/PkXSLvjc8hPAaQu8fTc5UFefktNtm+
r8p1MrCeZyc+f6WrsJ3PUV5N9XQwRKyz/I/TeET/A4XdIuiTVKWlKXXMedXG6MP9
xmHAlniyS/mR2jNLLsQvHTHuqvJZJu4WjgBwalSKeFia2pk4AKaQMzDoFyNBzsOW
T4nDy8WRnWF8VjEB9yKKM1ccFSI5hHrLq1SjS9V3l8VsDWj+s2518Q62Olw34xs5
2p4v/oXwiUzcaYWbOaCWsoWiIR+F8RgvhyQL3imO/98n+CMxYFYfme3NM6jVOOok
BxLATXs90i5QogmKj9VcwAXFkoKBhlHA5tnaTphkKiNaOMyCbYH9DoPq/AB0zccj
x7UDKHbQjMtvks7sAXKXFuBKRbNTjJj8v7tE1VArJlO4yMbWCxLswxmmRqx4xi0i
kA2IfgMlJgwFCWpy9PXOfoZSa62gTPDWiqCzVHPywq7tviYL+YaJpODe2TPeoFsT
JcJxeuAhgQwxC8kUnnrzmsMm4x110i3LRClbZmyMmwuixOkcdtoyxm01B3Ld3aDK
bQAaDTcPdkTupmJGeq4Z6GMHM0xdPvzWIQSyYj1W/ZG04cbX2dzFVpu09KENkFXa
Vnuw64zVK5DK0ZaqBh3zDuhzSHaoMDk89Os3zKFYUPoVfWWdg6Qp9XeLrNaSu31J
1A9yFsAYhy3IHhaHCRd/38mwfAOiVao3xBQWb6tFziRr1G8JoefSJAm7FWKABqC/
SCSIUxmn4nKc8VwDUSVN1LV93ZvjAazsBzday58eNcKhIHNdB50VzP3tN10lBKOE
yp25MjEOe8q8X/+e4E3FTzWg+jJ82skqWsU2pBml3UqV5uOpeaZkZGmqKDzCvY2n
QzeB0FdMbKD0ToYFtn1nvFHL96F2rgdHRm/Ad6HpA3RvZTsYltnPVtFTppBj+ixy
gL4PEuVacEYcfj5o7cAUMf8EaZUt0HLwwelZeS6dtM9B01CRnS21jS2xvLl4S/te
FmWPPJ6gEvF8zGGSfByDNJOgXK2dcOnYfFJuI2k1sewQVC0KPdOvFbzo/9UIO+Mc
13rmjFVeHns5DaifdjjGhCi7jrEd3r8tksxGsL45fs1sy7xJ0ggwTY24UJWpKmnU
cFQBF8GHnFBbQDvl+L0++KyM8hMeD0IpV6zb6jMLjFdZYXmLmoypjh7pW8CZdnE2
02bZSpFyf7vC5S+l+1HUCbEuMmL952TCmCVimm2RmmusTIhDdCUCYuTHIjFoupcy
OHwrz4DWXfuO0h/mz/rmUX4xTd6rsjcWT+nCGsAf6o2v/jNKT0nFmDovJcgavFex
6cQSY+7lfL7koO+zoH+fo9HLDwXuRLR1kanJ8ug8QqTLRsvPxiIot0YD8zHSQA7j
ZtbRz5uqvkvTpzWfuWCwfwaX64cArBze8bbwYxZB5HRQ9MBoGBbaBfPeYu4BXW1r
qbeg9IRX4hWOVghelJtMePmkF9iJoK5bW3iIAPBnwzCcCuv5sgfcLGZyYSqdh6Qb
SoTLYJzkx+NDM/mzGVoZ9o0biV3IkbU3KWVJg8gb92BqhnaQvioyZxoGHqE3A9rK
9cX+rgZNKXj5di7jFcTMTjO6Byv0JNcmFDMfwYMUojL/b961WeqP9PEH/lvt7WtV
umZIuEX6lpxbEJJotXGJk6mGkfdmUFlXGASO1oXu0gj4yy5nP7eIGkCjKFK4pFKF
G3E5wYgDhKVPPb+eIlmkMjaGHcunNqPcKe8x5i/IKP+11tt6qCq2fWKo9ASQTii/
e9hDs4EeOBuZukBU431xe4s8jbUsQ9gGpxyyQERob7Rn5i+5eRhiuWvc6jzBElLe
btBscEwCRB3PikzY528jkAQOosLY190kFt/uae78t0RCqR+dxAr2z2yskLll76Pi
8PuSNJkTszUJHNnLkgB6tsHskDSBG6n1xJ5zj5egzkzeYAi229v98oqFTeQK0ugL
vASSO2TmR1dr3PIJyyRW2hM0TFJ5muduUXRYJf31iqNVo9iupZhA5hnvlIcGIyd1
y4S2iOTqLoMLzNAa071lPtRzYT0jh70mpIKMmAJjVekJC8UT9dTeFBnT00+cuReX
rfpkHeJIMqVOTy1PW71uEY9E/DZF7nm4PxmY+ykD+VO8waq9k1iWdti0vLvTT2Ce
3+zyCyRfxTMdQMtq9NJjtp9TZARLlVPWIKIDb18X6mRyu7vIrLIBMa646fPNLJFz
EBgCtkVlIClPvcK7Y4KrW2Nq2yjCoMTvgKtddck8FcGiegkS3wXIKiIZJ0TSI6NY
Lzgo5J54Bgohf4qXAFZLDl0n8ZJovyxXSRcZE3NOmzpYHft6mUyBzmBv6g/gqmvw
7ggWMlS1BNzoG3QZx+WFGyvq8BTICn4D4xMWhtan33P7KsB+aPjbciCxx+IuIVdN
BIEYXzY0q/Nww1LPOng8/3rDnNJzR8asrBpTgThLtfw3pNkFjgBP+eG6GGjB7mig
Cb2oEwTI8o+ivR9aBI9VfI65dYpgtvuCk3esR7Yn8izRPbf5N1MKreLf40sYXaxP
U0QSSiGC6jhvM/EJMCFo2dErBY+/Hn97hXokyQG/0hZZl/y0qZMSzjCgBQU9MIAx
4k33vqxL0a6DUOWiPEB/yJeg9fTyukF7PKadH5UpnJcizxj9YalJEYLEiQj4l5Zs
nm9o0cxyq/lEq7SKzgnt7CzygGT6hEaP2qftMd9zx1WYnofvfmN9fSfKBerrlYmh
zDdWcrpYSrkq1A0Ma1+KDdcifOEHEeJ0Q6rAhVdCypiiMLqUnlYy2Vwurn/iX+SM
plN5kXBKdSYARETgS8BR6Z4T4SiGe3sq79eDuzMz37lkD92Udblha8N4hL/bm0FS
KtLwfYFBIu0rAcm8I1WHKx/WwvUaubeB4tqgRs3B05xi1FJew2D7miL4TIX31zqo
aMbZlT+JF70YPXhd134l8NDPQ8ih0E6yLFORyUgQJF8WXA91HmDvuA724bnCVazE
qOoZSa4Qo221xhTSmseh4mZD/nQ7dvKD91O7nnnq6mnM72v8106bAQCVx5WCeVCm
uWX0Gx7IdYPMnWEsjj8qTR8LYb685LrDa4HexOIApD0gAtfVgASVdwq5JXKQ4+cj
mpA0328IOTQY0WfgQvEmAnzEB08Ou6mX4vyRYfhpHWtgNrMdIW2i6MogKGQaxeqY
FvFOJs9cTFK2o5zNAu4x6u+rUZdbTBWkSR7Q+uLDndzY6OQTwPYssZTIIgcNNOUk
PhSJO3jk4Mm7Y7WK2VakBPKYCxFYpxsO0QUZzAJahWC/gBl1r8nicY7dLTd+jlsb
+MM+O20B14pVp8UsSFWBvx8SUgOywkPxlJesNnTojr/Ts0FE1ia8oPsG/soYMMtH
H4Z4wo5EI7om2ZL41kpL1gMjNcS0e2ZhnbINYjoRQte3jBzGfC04a9bFMc8OwshH
/VEFdsYjOrguNbJZMM7rIuFDJ4gOReYUs+yT54jGx4CfCSCnAwyJp+sadcNv8SUg
Zs5aCT/Ik5Rcm81vwyHw0nqfE2+Kc6VWUqdptf8JkflRIQpzyDqw2W71F3zniY2Z
mM3e+84lek0b/bYqztjPbhAf3qtmtZzPdPFPb+t6Mha0HwrTD9oEjW3Lwkzm4+cz
Kvf474hXMT+T1HMY/HRiO+KLNotkNlTUoANOMjJ3N8hWQhWFO3g1njRm51iKz/pJ
h/6DBV9zqoDMgrrvENGkN5i+AEvmowMMuTL0Ld+jD04O+WDPfuW2R0KoFptNrhke
klDdIhDkQAMaJewgaLg/qSJnQ4enLp9NuHlRMapvdKjR6FzPL+YOptiN3vZpNmv9
NymHDb8BCDztveAEOKBniRwTe4XKjpqkJacbmPqlHkJ4tQiVCXE3twWIv3OiErIk
JNPpFZlURv5gqmvDqDvAMljmpX92sABceY3jDTXrc0adS+/pFbQxsiC9K4Ghu+pn
KPJyf6VXU9JNf3jgbPXcbuBTyA1gDACsLZHJPL1I/5kQNpWESPuJRliqOUcui4Aa
cJyarkOPBZB7QS57YP7uvsCjlUUogHjLQ1qULh+VHt4bSukyPP1dSqRu1G9d/Y2C
ePf64aHQOJlLL1p0NBdA6KTU2QMOQjbQvImRvYxbfwTHiVJby9NKRbDC2l7RFI7E
KxuVoUUnRj6MLRtAh46mu0QFKSU6DW/UOpaHNSI8dZhG3cwbTCXgFDnB85Iz889X
gYy9HjVeUGAxx3fJg+z8m+2Gies13bTxdWwtMWjPjEythuUz2KLDnpDOhQyODJbN
7WzHrNvncKg6usRfdJ/MklTrk0cb3/tMVqxcQIbLOfGk47q6ElLI7vywGR3jBVPH
M7ZaIhPNSdsozzjKRjgbItaJPGogXXdKYOH8Sk+zkuqVRaXbAn3c+HZHC8TDeOL6
cbbWBNn9Oykc8ys2Z1K1HCZjJindEQ6c7YGYyI+E2j2tr0oAp6c2QMjQ+pxzB/0w
KXpSQ/iokQtKGVKOfWVP8F9pPdzIuK6eBC7jGmz7LNc3BWohf5q4pnp7L9uVfzJ7
v1hY5bZrpChM853w6z44+640EvnY6a8vmjyj6w338Hyl0tmHqHIYeyp80uBGCTM6
chcR2jix35heu19QPca2zRXjNq6uAwGSMjn67fu5OUy9BAOG78eqlwQF2ADNUZGf
RUqMnfdcmQeCp3dg4vrLERBMH508RdLj6sPvaFxAFQqaYqyISOLD4/fYXXvQTAr2
kDWDBnJAkLQ/1U39B8FpzR0dTOKks2T9ndlYri5ylfqvBWtR1sbKadB9sJiv527J
bE/G1eZFNBpTRkfG8bQ+lWU36l/mptEInyermanM8lfa0Tpf9O4bYAstD5kN0n55
VmhFhMh6JSWuTXIwR9iwvpZ8Kd8BIUA3GJQnVn0ZU6ULW8BQbIc1eIgduB86mvYj
oi2DcyK1Sitig3nhv6SQ1JrxS2z9TDRhd5jiLolJDAH7h/YqhTwyMh8rR4Psjsez
ZDgDat3p/bhRxyvV3q1tTF4mn26SxZ20ISpKa3VgWrbhrCTp/iTOwGmJuf1xA7sK
Yx/eFNQebvYRthj2ZQO61zBkFqxgYN6Mxb4RFD2ceTi/wok1ECSXPvh97MW818y5
DfCxwtjNjAZeCrt+ZCxwregFECcNp2x3puslxBj+FR0Fmsu2IL7tkGtdraUaGdzm
BxxzfZ8AlLOzOV7kewFyDunbW/mSNH/krvSi8pVLKrioAWdCUHWe8iIcRZavwwKx
omTtyg3PozuEnDxId68DPTfHe9y+AWE4RGBCgllyy23qe0VD41NSlxBWDkwPgnl7
XdMC7ufr47zkcr/JgQw3boXuUr1LEogGyNzZfW3wVZUNSelXRkHEIc8f8w5mqTHw
5TeUF7dTWGIATijMb0pVY9W69CZain1eidvdjYBvHy0snO7sfkJx4WCO6YflMi66
7BUwvU3g1KG77AQ4M0nozQhkNw8/dZa+mq4Clrnh407Fsz+1Rq9XBbdGWdEmwJZC
2stkYS4FeT5/jwuoxvU3wdq1zJ+MMJrpz0RmqQpF2rBqjMCUgFGpTPuogxO7b7IN
gIbEKIF2+nlnXp9f9Cs6VkBRTA42DUAU30pBhJY6wv7LX6YjgmbYs2uWKiUNdNd/
vviRM4YJ3g4VsGvIyBEwfpyqBFgYzMlW9NFqsEs6Zwz/lhk2UoNuk/VpQY8F8WXb
J3i9rpI+KDbBlBskUcTlUGZEhwnYcG5WTD23tw1p4lF6PsEFGNjuyi82Oey3jc9J
HrJOECifjVvh5eVqj+1h6qKvD8DH07GfTNsJi3vgb3qg7dFnivZbUMwdVRuYe3km
S+pZUQKh2n7j7rwcK3l+5/+2UGwYDDTtmhZF10it5idK7CS4dJhU6EUai0UQTdSN
POzD9pLP9OxbOWRMwLdFHsJjtDwTRefqebv91pG1RxyNoRZI0P/eCpHaIMWZagq4
2auBgu0mwK5ZAmjIZGCc+OcvpbmBnD2Vy2VFguyKXyAxTPt1YEcftuITUTUaVM5l
9bblReEEEEV6lmWe+9Zf2pH5JtVPcrxwvIz5YUyCRAs5CdGb2fsZywr4kdbfkzoU
7HjRh5BapUcSzwVWpqo62UnTwoWQNiEdm84d6TvoCMQaJ4aaDcTjam0ulys2Jurr
40ov7FNZB+Zlw2iBgQMz7Lu47pmYlWbUWhxUnbDe/QjtK9eVj3I8NtlmOiCVlj9K
cjatuYzu70aqVjOr7V2+nBSBT0EYxuLG8VjfAfT1zCCcl6JJ55TLZu4rqYnsTXn+
MG2jMxrk12GqdmWRtsW3BuAW8WLI0RJ/5vQMpIKNSG4gbmV02XYZxe4OASUGhGt2
it2nOKP0Zqmyd44ns2N8vvH4uctUwTgBlwEnZGs6YtrC8aeJVTcpH+CgWIaBQNwA
QrhHGE01zZIuZuVrlIBABOvTURmf2WYnnEBk4oPZ3Z6fVmlxLOCledOaZh5v10/M
1yoLKCFJK5wTO0zFBL8VsaTQphKfM0J/b2589ojOzya7Wfm+/k+Mso3RAoufDKLU
L/rSX4e1JDtDB/TLOaF6swq6p/eToqVXmbFTz0+F9zRCcP4nkusQ6mQJ1zxmFANE
Jndun2rhlbJRaoQjaBfYy0ACcbK8r7tNua8l0fXpywoCYOZP6pmQP1VErvFHIRBE
MU/pggM2jgH6wEPJ+XAEw098pm9NRj/wB73H1oUKGmpJazdkBGu5W8X73wJPiIsS
44vAbg8GPNWoI/ETc4VrBWnZVLs0en5Do77DJ1pBsYHalEBCoWQuPYCGZtrEEFAU
mgrmErvnI7TTdI6D4vIZSUbfg0k0z01E3jljMJhSDWVt0LuMAYQ93oS5SjE1JLmU
trzlGEIeGz6ekTqyqm3rIspKzXinWt9tGXuLdvJt4DrbLh7wm7MOkr4TY1Wgrnwl
GyST/jkx4yHfBnKWRiYzaCa+JMdz8oIIOmhS8xtcEcWG2q4WgCQTzqG6tgIY2Z8h
is2PuC8CmHcP5ZjaTsVvrnO7rTChlNyM01DubzTHS8Q5+/m3DT/JkN9s4U73EJe3
5cjCDsoeqV9GsdPbcHWnXeIOrTy+SKWA0irp64VtSJ0LVDeyLAuBtYdAI+qg9Shn
YiB4cYcwzK4tjDt+VXvKmCv6PaRCzs4HjC7ybT/TnW656aO5L3sQSC8b1jzMfJl/
cmfCwZnhvJ6K80rTFdpfwFhyMaqY+LH96FDtAjoe6tEaQT5RivNrm9lRWNMWGfEq
CrcL7aJFlji8hjIxCHBfuw5cy0VKCamramaZmEIzRU3H46UTfmaFz51EJb/E4gQy
BSPy6vLOrX9s5bRoumRnUQYKO8j55b90qcVBrK63dm4we4EojS4JSwPhR8HOtIQx
2A3LR2RYqB514dnjS11e35bEsBuOgArf2wdhs8jJwFahy4Gq+ZfsN7LPGj27MN95
gTLWkp5/Ypd1ul7BZXLON7zWBecp4rMc2mvmAoLn3smXRctMJFz+NkGXGeCFMzAD
BLosrpKQ34LgusPvpRX+fwsYOalGDawPyBuiHdVozRC5w+LOPr0GN7zKq3VcGi1U
C2RDUL/I4GmG1bodFn5qdqYJz4mF2eaPlVfT7NqDvYIgY17VAFEn4FR3tGkRF66S
nKTUNjVgNPlNczWcvXLR/ranF18WAn3GKcUMUCnHQGAqb/lViKtRMoHSzIsfs2rc
9ljmvBVyEdwYPbMk+hWTVLU1rA0S1COVAq7TkZhsHRF9lcMZV6ypj1dlp4t32+eL
divHfytZ0VrjnNMRJ0PASbv80YFTXz4AKlN631efHsvcn3aqHw3Z5CdxGpdt32xj
zsDuZ2o8Z/TVV+Po9c00/hr2fOV8WnvLzrq3edqCyoqjIVdiHY0zwGSH6zcCQolp
TsZJXzOrVxLUGVB3ZT6Kgu2QPTM2pI2FpBi3mmK8yR6bIeA477SUZkbXyR8g35+Y
1t47tOacz+W1VDnvF060cy2ZUqc+OGG63mjgDqlKx2H99RvnIuxEihM+Vr/Y35wm
4nXR7DqmkbCnf0d4g1OrLex2V9NVPTbBUPSbgKy0Eq1pOjwa/q5fRwsGM4Ka+8za
0pIpWpp9/u+EkjV1VUFzGmKlq+RWEn+iFh9Z431keqU3Dtvu2oUwOx+kSXAZbq1s
4ucY38lEM+3uzyGiS4eNjY8kyycE9kVaL6dAaBlT9SOVhBFWqLYaTYoyc1UpFl1g
bew0QbyUmmWPkHlc7TsTbY1xq/TnrPzFPOBwx4yF1kVt5QL6I3nH+/PgN8Y9yTym
do74FGANTuEKIgVP2yJCIL8ysFo26SWRYK8WBknUpHnqo1EhWpOwMMBWfvsUNBpe
j1+oRNjV97WD+dlB2hf13SFown9y0xRv4QMAnZ55ZY4k7YxKs2hpU5oPOcEBwihf
1iKa6nu4L6YPZkKw6SZvTJNRpQpV3IbsxtOrPJX1Teuyji5VMlTAKLoVUqD46ULa
UYhAYHM191jBLIARbqGXw6nfXVNhXR7VBZKps+pFj5/XBsjFJ2e/rTv7CLKffD1j
3ck2VdV5mlqMdjVsTD6aNwt3XmzviXNRArxA2KbWXRh3Qux0tvDSJ/OyhFgd0etx
Y6zn0zDPvH3MGWmuLSOo1O1Jyr7jPazDEh7ohtfcrxLZj2yWkRZn1TD5GsJVEwVX
8Ouc3Qnntk+nrqKJXltNhlIZPrm1F+gQlYNZ2HV1R9gqIVXQ9x//s8n/6a3ZoSPT
Xw2VN+lS4N53xXjTT0xaAcibxccl+UeGfcfj+5gN1nw6yU66JVVyQJejtBHQwuNi
E794YtY7EV6sO8FAAILLghi+qZhiElnFPlS2mDvYucqszgiwi/Z7ERMOH7uXegq/
9LZspftYQGSsIz7mja8DWvVUQyaMSeyQxVqSLWX2S8zOzYFcUdoCUaX51sMV9g+x
Nph3dFBM7u/o8VO7HOBoWCTRH2ZhsZSz5QRcnInBeGdn90oVPOfZpiWXuxT6Srv/
/Aqc+gptKct5b4KMMYZM2dWQTov4tk0HvUqyFRaY/TM4Daq62lVv+FIMG+lwEgyO
sg9MOC27WyM5+3qK0jzQyuzyO728t8lTlhMrT1kS14ATuzstBp01G67Y4lFoGtER
BFJYiXv5gPHnQbDimaReNAAQJ2ZD7qYcHVtxu/+b3PT9Qj7GWfSBOI4CJRWZLKOc
Ia+YivIdkNtEMufL4pvbO27LoUEJgi0cVPupYfwi1nKhlvwkqNLCOj/torwjNCJ0
dujG6wZZSE64TRHxKr6HpG039n1Xfzd37eQB1kaVG7taCxhBHpGyq7NxJJ0rnSer
KDqjioSiOpimze+OZKQLZi+T5Z0QX+pl2FvT9XDVxAdDkeRn5vJjqvSF6gGpSIwm
nRPV5FTNVxpcrASv0kkmbSsQ5zczoWsPbEjrxN2sedOsbccwCY+uvREENariBHRR
nnPsyU6ZNHX68B7cXMTo4/PSspWJ61gkujD7XLsyFj0dtm6r6YE8m+lAR+i9bW0F
p7pzGPSVKcI22WjOnRQPC2YQ0BXctC+6uerkYCTMDIIWaoqsEaZfJxcRa3RW3yFx
ONB+98mUUUoxOBjVFaxA+ZSLKQL4mlGVGPyR1qcEp4wooXmShoIkc0QzmnfAFh5O
5BBVd2bzRB0NCIxmYElScUw3Wc0h0rMb+166ywgrxqmpF3ljiBbRbiSXRh4EOgky
+hC6cWPgPWjmmEq+8JHFttIj/Xz/siJI8LO+gewCjUQNRSgBw7fyXjnaorNChH6m
xUzDJmdZb7kfgIVsMnEiikuqkcb5qUuJVe7ubeniJt9b9bow1gvGwXmLykzvCiH3
J39gE37/2l3IE/Y5cjjv1cA3EuhKnFy7Ne3BeI5MwNuQTk16zbrpxit6sbIIO/7A
bpxC7XwMp6suEOQI+OE0t5yZ7c01l69JJJpJLc+voi+4cTMVYueivCGo/lUOyeZm
WPoPXniY75p3g1T1U6lHNA6fjMNJ9frPKx9iDKAiGnpFgae5c1wbyzOR51yglpXZ
7xARUe0pFE9Tw9umXi+QVCvIL+NHtj52IJIgz71mG+Sp93kLud09KmLaG60lbhRA
XugsbCy/W5Z6CpyqUqcqAO7KFo/4zd/f8erPvXDyzADWUA037/C4+/O0Xj5OPNHJ
YLQNIBy4FMBjw1VcjSVw97CQdMFF6s1MEpZreJAzdFUX399ksE3wsxJE0ePIRoUC
QhDwCNe2PRfeGyQ7qgdMWf1aYP8ELA4pparvVWwy/Js3h695TOmDMlouhKW/EUEy
o0QBnl4awgDJtZrzptWjayQlfKlO86Otp00ndLBQIQ0wspqGcRORGuSd9TzbeWzH
X7DXtHrX3X4zzknOuwHbSAvtniufO/n2s1ysSeQR/fM9DYRMP9orkRvVcf6jhwqp
ZnA+e6Nte1dJwxobGI/AifmkqwY67YsapzqM5lv3aJyaGS2QOGqTYYDykZn7UIx/
lZf2mwjwwn7F+xB12vhUZ9X6XioxCM8z1UcF9NhTqvNDuX6lNqTc25iIWfkQDpCw
V7+ywggz+3LePa7iIVGyhjgvofV3uH5B0kibIEzd5JcUYrG61dmWK8boWhTalKwC
STU1SvH8gDVq+B6AV7LiMJouH2mTefzO5raaxxWP5/Bap3qKWxQKYDWtuuRWZoHR
Sci00adn+nKCZnWuP/TJWUiFGhGYcZ9iWLx8W0U0tdLxT+T7eVPXTOBHdqcd+KcF
nyf+L+vtIS4d5434CakptbzxJODCujyEpeMQXN+FZsyJNx2nfysyPUlTlD9lsIUN
VMo4QRx1iK8oyg46SzNxFgbPMCG4X25Hu3BAnLeYYaat06rkbI7cCxRIPVzvMwoi
dsAFNDnjvcvEvJRaXCaERL/Dz3YMA4irHD/WYZT2HDpbTgZmTa3VJg6NbAi/ppOh
yKepr3WX23b829OUdEEDsUUu1OMFT1wgnLPzlmwtAXnb40E9ZQPTUyi3R/Voz6i2
hox+p5Z2Mi4qLDixfTp0+4pUOtMg/JRl4T104lxVuwFSe2WoFuXNA2TNEXhsb3R/
jZFdj6B9atXGpaLuHitc+gA9lVf3POPEQ7l4qkI9XZQFKADlnmwT7ddc76TzXvUj
Aqf327OeOBdz64y8N1NI1lNFIFl7OY4MWxM52OoNM1ygdlXAeYH1wqXGH+0ZSEdC
LvDwybFEMnvo5ZWD9APjHlUd8TdegLKmT4OpeGvJt/0CyT05cOaTK+hkDrDmCMoa
YRuDFaWzD/quG/1nnYX/IjWMGWXtu/eLWIcCk7vcnHoA7TazoOn0AjKQab4/lp38
NigQdvu+FuhzoaPFq+sCZF0uhoX6H14bFvR1yPV3YLV39I2qgPAETHpHVaLeTfQq
9wMzNAndP2iguKVKcnenQP7HBYCUMhptb1AHbHY4F8D7MkFQkXWQ3dbN4jDkn7Qm
GzryZipIAlUw5gxR3tUzz1CyS3BRRrbbxkStnx0LdGNqQj09jzEQNuvh5yxxgcST
wlakcgR6Y8/5eJWignf/4c5c+NVB46YPN+/t6trrVqMllGe6tFZ2JJQVzuK3Ix4n
hAjzjkNUPZiPhVzGH1QfH8yUqfcDFfclPu0tazstSvBuLi1EiWE55wWINcfUh6J/
fOwEJ4xxXpsJy9DndhgnjuvXw43ypx3YQlg6xt1PjWeD7NSQV54R21iV8aY35o0a
/Fh4VNqdYfG6mC2Ji0p3aZetkIy1jzqnmE2llZWa/V0ddotiqhh/wDsVV/PMu0YL
Du20KQr/YOwcLtgY70buCmBk5qtHhfPyAp+N5B3xKBVjUNYuRGL5zRmmZlKupTp4
1V/t+pmMS+H90w+Ahz7pZdwDg+iqt/7VaXYtjffnX2y0Uv28TuzXKxWmXJj/c5ix
7DoARhdX+G2CIH4cmCjIkA8ny53d4vZasMO6n2vE0QMK+b+xniDysjMWypXwXTTy
g01oODGB1WvYaE2qNGo8ISb6TRLwib7ol7ZhM0tTQqozzLCWWDJ44au7N6FUgiAz
XnfMWZE+ItRaGmNnEUyfx/oW7km+1MxpQUrCcagu3f830AfDqMGG3ERnKDMuYFCS
fpOobJdb9xHjgZRXlSzhB+7LGQql+WhxqUoFa+S4zU8K0d6Ku9N20eiVZciIUYkk
BfOZDlBkGjjtO4yMO+1pcNX4KICUb2/VfFJ1Gi7+77HDjSUbsWlFT+6Xlkm9VJi4
YVAOHrMG4LKWM18PU6EFQOEZAdp+JQL2Ewwm7BqRSaE5bpc/wjhEebj5jP95S4Oh
6Ampw/+DQo6Upr7RnZVL8KXAPvl4i1yQ+xgA4TNUYuH8DOW3lD05oyLIo8hJPNXu
mB0URvVbrD/jrGNkIGBtYSgqyshqe9g2rE8X8PtrSUo3zWlPAp+wvDVBr5GX9ytn
vxU7xzLPvktGk/D1yAJEpqSiptEHUtrPiQeBh3SEbSV6pF0mYFWnoBB257YETBem
NIr1M44wxtOPzvJ4YVjQRXTOpCfruw9WDCYT69Wikc6kb8c8SfIfznSoINIX7bNL
P5XvZg05Z1Z29hL6VC0k9Gl3UEx5mg/zL/yJcW13J0MAParzipDDYA4Hi0PUI4JH
jsxzX1ItJFYNUcUriuvZsAQRFZ9IXwjJv6aM+wplKHCl1vDvkYjku46FKyOlG6nX
ROBaoji99kf6flUyMMfk/D7dg4jNFv2JARX5XGnneG+XpwAhKAEiRhVNp+jvkxJy
aLCKznhDVKR4Apxr/ZuTSqmNbetaBc32nFZaqWHYQTpVbJLn7KGTeqpWQS92y4+S
v8a84b6E0EFejV55JI5vq0hicFa3K/f7G/kvbYu3p2cCtsL+FCME7KWWd7r4qLBy
1EPpKVWOqKYAQ+jD1R9T58CWUP4BviSs4z39AIqM2HAekbxaKw90fiqsdctWeRxb
GZghXwQI4pnLj8BEp/i5D3ttotd9xm+op+R2biFN9EzT2bNmgwTQ0E+I4/xa8Wt9
Jb4gqgpy8AAzvRUAWWfACqNxSUAJVAgnlp7BJC0q9alHju2FI8nN3Qxp04pWzo3u
trPtwdriI+AK7o+ExJvtmoHROhcvsJIdICg2Ee2PctOEhU0/NHFRRML6uib0hDuX
3Zouy7bm3V4PuJctj+8ZKO4dgAmSs9KT0dr/FJG3TkDbllOBID1D+TriICUKkktQ
SgiD1lngMRn6HvVxZcBfvPqnOdwygukSzrRh5N2+8OZn4bhmzvpzNWThJYVTXw6H
MKwQx7R1hggCIFqqtXM/EjDZiSoMk7SBeHtpMO74j6VpNjk0eFaGk+bEh5j1IvbO
TGs0Bj8HAPboQ4TQP+Lltt3iXIOaxSF3P7HjiqLngqaRUIpGPk1euGaZeGSSIJwS
fsAQyBv5lmpDbqY9XHsAzU6uyKau9fdJTuBmVSbW6siK8f392HgZ0fKqPDDVGOdT
JljVfwXUOPyAPMuKRBjyJdB7n4P/YnLZBbPZsFcTW8XYuoQlYAaDWSXgJ5wKSQhW
ElvA/Hf01oZ1x9A0FxEja2+NTCehX+SA34XvD5Rw0w6k4Flr34ewwICAG2zybIRn
KImnuvciTGPh9CgX4asIYIO1rPogL+2S0c0UKzYLcWoZ4yFmkzwI52SANQB4TeOo
5K84/rZznjuAirvvH6Nv8zHKSBlWK0ffTT5KP+32KkB8DVftB7HwD9RxogMzMhdQ
SMy89ULRJgzmiPK7Ljh/ykocNt9opc+N/PY5PqBvlkg1kPyy5CeUkchSZO62QXO5
zCHiXtX3U19bPHFRhASs8Wniw4VHFoj9nf30aAbvxoCqwr07xEGKgA6AKDLmVXEv
yLTd1nO1DK1OrIkpj7tPk5y2bQJ7E2edVLeY/3J70Icb5+P5r6Loh3OpVAf92sL9
uHw2Fbyos/m1/qHoEXguc74RuyMwbK2Fu44Ss/YPxyx+XJRZksDRrftpmLexGeNc
LyZYItZHMLvL4EyBKDU1P/nlwMfwh+i7C6uVz/BJawOG/1644IogN1oSXfPsS/X/
TOs24PTKbP4mfI7POZMEFCdzGdqiyqdeKfumH5d7XXYgZ/elJC34wY0J07Upp4rp
SkQhu49oKB/GRGOdPbspn/HBTsVkRfuO8MdwmF5FiVMpah/rNguptScWmQGUpIA1
f5xhs8pIavSfK0Z8HvqosCR12TRc0X4XGWWXgg3rJsRd1BW16hKeUvHUq98cgjA5
OSS4mruZLZmxVCI4bXhWq3Wy+atI8EnciqNWITZurrPoy+I+4Mnrt89KPxkfGm4N
qNHpLPZFxqKy/yb3vJaZUU5ElbI0uxXlIujDF49P3duvmyszF1Uo33lmlNvvZPvy
rnBhJ+amdWkvC272htyy8rW8uGVq4P2czqKMqW31X+LSGuUaViW98d0T7AchGGne
MZIPH1u7wWKqJ4pLz+8yOtrYzhRrgWiE+e9YLLi7oZoJ2vdH/+ftonvht6tu+f+E
AmRCzWFGqrbDXYUzEHl6T+TEWJtGiRREyyPuJaW66x3ISzvGx3pVtHL6Vzf5s0/9
tRBIFmSXGKjZpRGl66w11eauq66PxHIIyHkAyk3Cct/Ae19GjrYgiCqnyrBQYuxz
PFjDYRMtRpj//Bx58+/OD4NTVIo09Kts8aCr+aCH5GyrlsYGfTYgYKh25ABTQy4a
1Zx4Y+wJ9LxKGMYz22E3soMc3NMHhEBKnjVDuWun9srBQNooZj9VKbt8GcqYIx2b
142w92JzNIcCETdkWKdWxJJu0vMN5Gl2JeMNBh1C7ostdZqYVK1ecBuysj000KIs
MM13lKpjnoNgXDxEZaXufYMe/FiLQi9zeeIALNc9QL85aQMGS4qPIFWLT5H+3xl9
vInXUks7OU/Vlg9Y7D+7vJWCZnle4kU/sO5B86Pw169wMWy4Dw4Xk0AR/indoEx3
ruh3x+s91Gy3f22jCSYUttPLNN9Nk1Ls+2NfXsXOlb8fqthspBE1eT+tz/Dl20Ur
wc4WoebQiBzA/SRiEVjEbYKvvCjJ9aKS6kfDbjmcxewDFop9YSycOLmcb4aGtBZL
eWIA0DGV5EuvjpynZFEfC2BGVPsTTNaRuHlhYkCFjnHntVHh7/8vZ2k9gagMI1bJ
5IwTPLfRE2hd1mMhhC5UKbLgDivb48dYEBJopxY1yWcJjdXYNFK+MS1qOHMEfA3E
I0jSH6BafbesPdZj04Tu5kqe/7+xP38OOvluLljv0jt7+T8pTkm4m9wXCuSCJtgz
ecBrr7mLbAki9V7u0A3CkibLnqRqiy6v7o41E6OSSkHJByXssCwRtyZUsR7Do3qb
ygwDL1GUmqtdv4CDCyLrHFrY40rXBVkGXe7LZxcSEKe35xrJhL2YO+uSYK/f1DCX
RutND9c2ASxomP4cKCVfeGun83sc9UMutswGwP0E/uo2cQGp+vZAVKKxLWVHPT3F
ThOcwG1PBYuf1VfJrXtsIxzSETcZbiwK86zcOAmgPmU7GShT8BdG0OVFbePgBXpL
/SS9hF2bOqZDRihhfs/WSO2065xdHeWQdNwlGubHRl5BWZAUIhB5+bDD8OdAz8mI
OVxvwmnve7YSK3OjHm4rGUIfnPjqP7wkYxxAqyNp/sEicrvHh58ZdWAI0FlNRsXa
1OfQCFTAp0mWbyRZPKr3uTDcXSdUAEX78xNG4lk1Xh14CCZ1g8yLCZ6eLaUEogzR
nOxL88fg/aOPkk05Bn8p3RUoshB3/9abi20WUfEa8/nDGLx5fDRJ/rBBb+dSHTr8
RLC5AXFpllN1fzAAYMna3BLsfucfR/vsimdI9+EGPrAyipY8LGqPRwF/Vb4OZ2A8
6TcxFJEnzJj20II70dKCehkDg3QzRkICavFGxFWSy5d3dsuFamidqAYkypJ0lSOF
5YNqw1GdRZCx4aAGfi3A6pomk3BP2ksCpx0xy4UeUQLppWzfoqmNfoKFgeskCvOc
KcXrcse88V8o3udK9M4B/us+/zWMUt8u7jlx4t8/TvsJJwq/D1C5A+m7jexM9jbB
5E1fORvXpvZsXHIwWG/OxMih/aziFfG1Xq0q67I3YrpiZ/2OaY0i2rAobMNAnIR8
hmqUC0IGY/XYAAVvTWEiSMdLuX6SS9QcIW0Zy0GSj/iqklmqyed8oG6/MKGK+wbn
sPSRwVPghFl7b0L9Zf7rL847+kQd2nZK//PeMenphEyM7foDQDd2GqXfV9rxbf6k
+8aW/F9coL4jHzNnuOPCvQiw7hjhU95va/Zv9ggJ4sU7UX1aSek64Ar2oj8fEnwx
8xc3qeKZB01xKQbF2rSgBrUJ7mtOPfloJv+gLiHOkLWTS94FZO2k+egyIfgbUUX7
ogzi2X0Mhi6tJNfwD+Bm1Z2B04Aak7Q7WRbaxY9pjM40r37HDwldPIB2Ac7yAqf6
7zofu+/c8imYOm2kEnQCEtpd3LoRTXdxlmXwuA4NDpB4ghJDYWqbl3t//lHmX3AT
sJ2kbT1nkhL3vzNJDYJX5LC4jtBkF+ORzdFsyylksPP+UyQGnSH1JAu6SQkEaJYX
p4g+9d0ZNB5oCWF4PxQgrRZiICnQZQjzpxYzy8MQKSivnKAkw8bH5SXSVzwBxG11
FYl1bmuDw8QzsFqEPOU+kAdJ+0rAQFhp6ja48JT8qGuPhx7cjVxDapilax41EtST
SW6Kfb3+0rx3U+B31pV+TqUAqy0zXlbPgjlt5WLiFgiQdtqSmVvyiNK004PEd02M
bNvekcuU7ks59qsQMMLYEikZt3C1jYpj/arXZENAt4q94FSWY9QQV+sG/7HdqvRF
mGrjlbAbrbXkIUknN4mdGUo71rZ3GYbvzAYSjBhVVlYvC3RNMVu+v2t9UyUHF5yx
w93YFSGJoVUKWuxU3g9PKNKO6AWNg2UutSHIqfZqFkUD+kAAigly0a5dCCecAVSU
M09Wtho4Q3JjYU3vh67zJNkMhyKTVHCGiAwv6ohZnqt9E/8w5dALiYWd4enUnJRK
YWabQCF9hgjNDpDw//+y5MMyttaE9WpAXvPOYJO65dQdiwjMnAGvgRF8iAqzVRBI
47uKTMM1E0xa9S2Qm8aQpSJnUOU8uRw9czq0mFKPIqnqFqw/+eASyqd7mCtXoO/O
54l0xjAZGayPqSxXt5fP1/FYwfM4/sa9K9zZCpNVLr5ZFl/hB8Fp43MuF6SSRBcL
o1UCX2nQaJch0r2DRpf9dk3YxNHrxSS/L1cq4/Kf/VTISxXijx7BFc0GfxGKZBkA
iMGs3RvOUvXfGUy/R8s/768NralB6fpNFHGrJ76VKe4Pzu/dZwVOzOMK7+5g+nLe
4kboAkCL93qEPy3cSyV/CeEixGM7qdhREJlQuR7NfwS3k64znRSx92bIgtwRGOx9
iwzmkU+E2fARGWVSdtjr2Ug4Q4MYlVI76IOv/c1gzfHdQ31CYZu0t1y7fpAX1SM1
zi2seZwaFCyYF3aJGeEPZbm15sbVDF+lxRqkDr5akEz/Do0S5b/baalPtWUu+X3I
NWOa2Q5/LvuGNZeNxQ476CpOqiC+qfyqfSXtpgi5hIzdc+kzPVdItvmViRkwdKNE
ZcbBSBWUuaa8m2MJfdzRcXIdghymq2f99G6jfCqetQG7YVhrfY2AaMqwq2+23hR8
eyGCNA125csr6vXmtu/hWRT/c8u9dy3eM/R8u6xIaJ8+VqEuj/E8H8WrbJonEz8s
zfXkg+TST2ueUhUWpvMP8mm0t9ltXINA+dxDFhmEUh0Qy8+ljvL2S+sH2Gf7JGg9
bV7GoQyles+e6rwqDiBhzaqIwBB93HxOfTct5OrMjfDYqJKVsoK9pO3P4Nd5pEDe
emhJwPALCgxjbbqAGKe7TuMKpgQCMP+MJ7CSZswOgfqs5hJGRdeyJI8ZCGQ4g6Hp
YRg2SORug+5YCmO0kKuw3oB0kXlRCZu1/aWPlRrcXCjw+hGALtBD11L5ngpfm8G4
v4nbBWxTdSSvaMiMFlmoRbLMIy0bSg8/gK9egN3/rgeYlFCZLZUQtmaVX9YKdr28
ilARhP9fCAQTI2cyoP+FzEdCNFEBLHCf/UcoV2SV8xN/eQJzw7APQ95MSGOogpf3
kYoY7EgsQ90alpOZF9zgRQaAMOhYZ2VTT6b5FKXkeGSq6Dkqbb3o9jw3jkqwN+TW
xurb2uov+kuztUAZwrX/rEvuH/SvHteEU2Bmlae78MNiZM0GngzNB1FYHa4rUEgi
jaN7jqyvK03hWGBnijIui6/znGalAa6JX3L6BhuhPiEx3q5qX00OZH+UCSCbt2O3
31n0TzxftNdg963FLcB3xag5m3Uv+Ncbxu+RraEM0AvEHoJ+vrI7q/Kg1N5Ar5yy
Y1aRv9MFPDl5gmvP+bHzJe8nQ7uJhQp/i9k4ZfvvzT3XPUacqL4B1oaE2vqP79d9
q9F2uugIpE7Jn/9N+ATEplMcbIq6GDUxMsC8oTC7c0USeHXZ4OKGMkvxoR6b9Ki7
We3gOcEaPPq850lBRFWHZj+pq8hD8Odg/6uYAl3Y4i+5CdTcoKDyxoxKk2uS8LVP
HaW0EDvTwNXShHDRAj2WIgBNCapUVskPTQQBXYG24foOtMRvhwPrpB7KFT/xQt4i
hnelIUooHRHdzwiQb+gSJkCyBYR7jKlw5akMTWqVMiu43yJBBZw7iZE6b/oPqCD0
5c/99JfiOpdCQO7EF4RBt5wOYt/4DbLwkZRWm/bLtO2PxrJfF+IsYGYYJQhENhPi
AY5VVlU8Bu1b9/vRABCbB+9BAbIjACaPwWugpFzsole2ijch/CYCcEVgBCAS9akJ
+wkb7p30cEObK3t0H1ma52oINvbLNbXmqTfQuz0yZMbehUNtLmDqsmx9kw3vmZWV
lMe76F11IcAlJDe6uEyHC+rQKjFDK65PA+FjNPuXvzuQfrDc+bs9v7v+60mFWsbR
zPAc/vu5VuWWdRUNcVgzLjdiome80YVBbWDRvf56dHLow0QVUHEHKgEQVGRHktJJ
nWmHW3Vct2+ox6uhKW8z3RbgXEdKvwXqULRGnR8Nbz0pzpaQvowjCfRcerSHPE4N
SDOGnEekVP7NJu+wc7F7nxNQsjnAG8ykACxxwUfl5rpcetoUv7eEmfBOZUJCpI1e
+8/sbCe0NydES1vLlWx/6Fb5Qk7R+gDuDTnKtcnAyzLRqIT4xF4flHpNAjOR+QDM
sdfiXt+zhGkQOIdwEcEf9v+A8+ukdSv99Jb1koJ1HAXcgw1qWgEcTqnKy9m+dyft
0bAEDR8TqglEHof4/iAuUEfo+EVY0/EncIwSKnsnt2hlh97fDAZKYe/RJdfN4QwQ
wCtlTR7tsoMRx7fr1fkhb7/1Ojknt1hCjBlrovO9gTzbog7+XijmALA0yhrCtSuU
M+5YXMgrMkcb4DuTOITYCGbrihYdke+AdujGF5mlEH2s40oHLdFPOZXXAnbjAM4R
Q350XL3UUtfDQVyUuQC+ncH8d3JcD+0ZO0AKsgYSwKu0tzy1QdM17EUuSCjyhJS1
/YJYdChanUF5RWAtAq0zc12oNWjAQsdrTp16flF/KETgdUApz3IDJCMhYSEc00fp
clHcj6x7ApIkx3oCugaUowzZ7wYouEt3DTGrRDiKX+HIcdAJVbkerDht+hBhM1j3
tW/7d4PkBtEwqWlQFAP/Y19Ca3ZGEwYn2HvERfjDHEc2/lo090Ys9dtugCGirzmM
EGDPb4Ag0FsIXYuCNKfBW8qMAb4Xv1K3lcxBIry68Jcjh1jiPr8EfiUu1+L4zcfF
F6t8Ug7VcPrb0bMJl8aN2VpHAi8DATLzn1/FYwpnuSPs/4J8Ualm7x0D3KKL12Xj
hX5yDyrQuhmhxgY0SQzCmM2rtyDRy14CxWQXGAoI/8/Gm88GqqtdoNZrqP+BCI3X
m0QuIONZSJfwz6NRw2Fom0MCBhmQkZ72LEu/cHo2OfpzufPiTugWmQE46ByjTQ6c
jGgUjuU9S+pBW2ml35164GO1I1hK4l3qCRI5DjCSxLXG9vF9dkx09nlX+swrbmRs
OVygBv4V7vwJozF4rcdTQE1PoXczO/kalYmfeuLzn40ICtC2WJKDimSL1kcQBMfv
RNlh6J0AUbHXLlxIG3axlcX5HGveEWmo3zl7mWs2ftv8gBzD4l4Lx/7QvS1drKhe
TOgQmPlAgJET55DVzmpAKoGBVVd8zWTBMQEJ3S7ehnrZQeIPuT3DkgOnkguJp1WI
MNoOsr7sEqBlwPxQJo7+qXLIzHjy2az/uFLg0gkFluG5UnxDxjW9CMXq0QqVSXE2
yUbR1YXFBJjNiW/7fr11oqYlglAU/6dTAUL2x7nOTlAjv4LfibbUPVWeJ1znKz+X
8XNbFEYkeC/vIGo5J3GqNKKl1RyJ8ELrwE++MASLIL3xOtC5wP2ZRQbTbtd2j0tE
qTOfG9ECpvnFRiTqYjUg585XoY9X8eGXsLi6xHAELLmFTYAzm2yCtsYZHRSYUoiW
JzMoQyPWmbthl1Uy/N4H5VE8UA8SE8bKvYI9te3XHRRENeNBtplpBKtH28b6ZlzZ
GGWpGnqPOelRxQSlvHMrtd04MgdZ9pQbMC5EsHPJYQDlJmAJsc3qxrt/YnGmVxeZ
+soV3vZSN+cKvVf8sdpHiegn/704J26xAAykD1brnWbSG5eOxh5iZ7V295OAevuP
zO0TYeykdqhVC9xdav3o+JDoJ5md7kL2hCgmTbsb5wUDuEQBrgg5ILllT+aaofnn
r8D0cgnCKwR0gZi/hoCsc5DhhV8J8JM2B86peAOD3jLevnSgC7Cq9m4tHAFVWm9m
HDxRqcIrS1bBEZIthtWeDEfmsiCbkQ7oglnoqE2+rtsiC4kQDiqZzH03MqEUh8q8
R9Bujo2uIMY1AlUMaxRc96TnCYfJBkzAH35gXNnkJTg9rrSo+MZTA+USggWEUHUY
1kpV/K96EZnXw16+1SBuWWlOJarJ9gTCNiFyjRtlx4F6ZZ1kmsYrCMzTP757V+r1
8evn4CLGyZb8eNpBxnmObNkb/HaIB3O4PwK3y9vsHEQlcFu077pfAx81I44vPprz
8XwfVlqKRr2csvIkWuS9FXm56y1lvLudDWTz7FQbowv94OXSuH7VdXHErUIaJRtp
kiJqUbOfIwDPlcZVK7vWA67o+gi5vGODfSbDcljpwxNm+TiXYqUe59Oe+fqAO76f
W4/jiaWtpVAUXqG+aYpkuogl6kGuhevGN9iq3Y5ZeDgylUYvNgqAqQpcSnURZR5C
qik/xWVWNixZQuEf7kSvkWbCQoKquo8LcoacCIxpIj/TEsmSd82CPDLIAuZkEibA
pHM5kuEp4qi6jQi7eQ4ygf/sx589m0cUhgyr++rVwsw9NCDju4uh1sbrYjmsBTxm
z1M7dqeYE9LdgHSBBX1YclVcky8ATcnfI88gigWnQZR/88dMCqk20sneRDwAGDB1
4oYHCMG63f0Y8HmdJWkGg/mL9VpW4sHCOQ9bE1ernlzEe0rzVg/94wTf0hZxRniB
mqXhWUZ02/7b1F/sQRV0Tpta9NHfXjkEl7X/9K3BGM38fJp8CHxd6/H4rnxPAz+X
kn6H8xOOlPzizoVWEWGUBzSv6qgkgoqjx321LDwOeHt8JrFVpBbDDncNbMkPk9KA
+0mr7jJkDfHLyO/0QfG9rdL2Obo26SKrfV8zTkHCuYwCyeDxoERZFXFRIu6VketQ
OEOy2fWlm6YEf/vvHceq5+eoYRGaO3eU+1KoLLeeVwtYj3jbjdreQYtZFwoj8lx7
v3NxCrK1tuvjuOzxukrB9PCfjq+4s+qwdel6BfBBthJpCwMY2HpDEPcVudA5h707
gTlIrH4LzHyfZ6my6eZ0JEaRGBQJ1j7LqAe6lCF/xuCKkL3KSm3r3IX2o4W8CvEO
K1L7f24HO3sITazFeD4OCxRFEoXIBkZi0bHAiFY5Y8X0Eo0Ep/mDAL2WkcJuWrOk
B2p4ZDkQO9ikobKLvLsKmaRxPQk+71tS0PsqJN/rtv+CTdonOSvcVmMo6/89yguF
FGwkVzucJzclbJU2m0iF2RpIcBadLYj7I8sxWqHc8Httq1mLGdA56Rl7d8He8YYh
A/WBTL0qjdtF4hjZskBht6jUKfVilXFsFchF/L3MKErfoAFF/7Yfnb7qnqyaMeEt
SjPmsZXbkqvoV8LAJuJWwJFq08Lm90yLcsJ03CIGKWXptwhQqz+82CWo19HY4Nm8
h9Ucnpw9q0mWQgrbI3cb1+jWLNpaedS+1GogBsdBBWk8TJIsB531jXSbxdQZnM2j
TSfBdAz/zOgIm/7GCx13oRQMtf5zNM94+1uiZDxjgKCODfAJMB+x4P6pyBf+gPQ0
96BDFZA44IV3xP3WSqZy1jJ+IoDfS5LQuCB00r6kn6dXY1jESdhYOuV96RQEO2hA
6XFId5gKIpIrd9oYzi3M4zSnYvOI2+yY2i2dJXk0PhfJcPCdg6AYGO/172EdRjnp
9UrrNG7ToL+eeEKmnfthJBUMwZuLLFpoYenIy5eeR3FBB/9hrQ3z8Thi7in/z4ZO
XtXet7mw6PdbDLjdrKGkW+E3i2vw8qUS5WGDkmpIPJBsinvXYdrG8RipXy4ktVYv
DjRE/55HXsFSOe8FfzOgohShYkQ2RqogOsAkiVpHFVbRvpljxVQ5/1DjgS1wA9Lr
38Ycho+6jxDH/llaSoJJnwbi2mF/J8aj7FWvGVajDlK/jP04/nHG7pp3C3TznQdL
K+4atvq0RtpiAlxl/lZLx7VijkFcWJ764oFmNBuvJapIioMirQ5X3QWFYKsEHiUs
fKEb+R7NaMdJVxCPZ2RSBOIrl901klWFyNpXCLWyvRjL3H0hFTJi/+3VXch93I1y
T/IbMblildKQcJiymXffZoNn55S4x5KNPHLJqZZT3bzLuXRtMz79RW9cwj/fM/mk
OUh7ipVmRjvTNqgOrI1PL7pMG6bFl6wbgCqNKWjAjy/HdI2lSgeuOZicVV9pbncO
RDu5k1gY44QBYuWkEOx7HBKf5Xd21Ez4r3maTOARBGYGlxJnhcuI5zIt1FlSlHCs
Bpdi9r2hEWmyYy6l91KKSnrjZ8SwjjoXHNgM0l4BiteTZTnoiLWWC3VfWLEts7ep
SNY1926bRBKav9bvLRRbYUito1y+DIfYEb9vsW06905L8zK6Iq6WW6xes+/+VDSB
re/hMGNMRVJZDFHoOjZUgKbflemY0wr7BB2Ww4enWN85N/8SC+jGFM0kpuMQjVLy
3Fp/qLxC2Xl2C6zmzTesVpwbK5cpsGo+ZQ+QqRODI9rMT8TjjWWygOpXThigsKRY
TlFjgjjt+gfP4xCKd1Umi3crsTzdTkX55/6uqLqDDm6ngCUfTpdSsC5mjwmSh5qP
8rZv+umHelV/Baq3p8sQx1vSTv3whjg5zZupCAncV6yLMeWTl2EwfqZrxCZHpE2q
Yz8cyY5ZfKtswghiuVlf2Rrwb+FwJQVuVBSOtPMyYIocxawryj3JQNtFN5oFhwJr
y07klKDv7NdNcPvvBMbi8w8QMWHafx5uCUpGkvUb+9cg+EG8Uk6qDY3w+oyerlLR
R1Year8LLDU5yYlEzyLzOlbi/lQIEIYXLu5ynhL51HnhjAdgOwAdmVkkeOC2JOs0
ar5xQuUgBHVPUNJj3rb4uu91lh5v+eXpp8CcgmOBKOGShsNirz4+ANub/b6u1kbS
/gfOFp8CyoeglW6hnJUBiv5lV77n3RXj68iqobrjDgTHT2nJAoh6HrQsvvAycB8i
Rp1eOdHhExDVCAxxHd+rs1RhHSy/qcNM/G/AZPyWzONvijMMBigepo+nGXKtOUqf
n8pKHXXxhSAdD0CTjZT4p8QXJtDA2XKzwEApp5UQ7XwSziG1pNZfDpeIYzSXtc9/
UuxsDgd0SjQ5sAhu+bt1u6fhsheaERoRZgQIeXMUxvdYG3/AE7YHYN/LOssXuKqd
qKU+kHfgoWFTmcDg0w8/a91u+EEfN4NdCLzepE6afYEchmdFGttNY//lebTHn8jG
hpwhE9QkvKYWYc/ugIjKKy1P8jMNK2otuCNwkYV1t0nVCgL5dQZ3jN24CyUdc5l2
gSps0jsMxD1k6Izof5kdU5e1fsxXEIAJVGd7eb6MVdfaE3DUBK2MFL0snTJeEj3N
2hLDAUpD4hFNaQ9EEzPBwIrxSCPMGnc/sKQ9Ew6W4kTSqfGJPoqHxk15abQaSB5s
ST2fjk1VEdTQBmaAFnafk2UXjIj6j+HYksA0+6d8nC1PERuSQDDnUx5nQkKQk3Ir
VgoUROGFaAzQwAB6gvZ3E1t/aB0CbU2TonM8O+zeK15TXHqakUmpGtQHVM9htesD
7lg0r8vDcv9T3HJ+3R2yFNUMr76tgeN5XaLMbfDKxThVtxZuctGsDx+2/S+gKBJ8
IJ6/AdkfyC7Kzd6wQhARNs9k97e1gFaxK/FHW0PEGsdMIHXMxIssBenDtu6vf6y1
ckKxuIgzdILYPvdF0f0a4tSeboKJ1dxogIfk4Kl9VWpwxUrEdFWj6MwhJMtEdoQc
1C+3Uvy+QOfmtX3h6Cvw778kdxC2pLICnQ4K7M4ZVtHF/sZ1G3qlxABWrWpPk741
ECUg09W9etpdF3v6be0GppHSQ63FsjnRvq7iMZM/R0ATiYyNqQv2f/hhVUHHAZQS
jqUN+QAdMNDnWK+hP7auXhrZL5V88wCSG2Ege/ECbeTdrwccYkoe9PtEscqgXPY9
1Of4Nz+IdwPk4O4JMM3fP0aclm55yanNCXg2bhtnA4Nq945BTgVEtJqKbT5dThRZ
KvqDSrtBUu6UICDrTX4Ckf8LZRurOOVvAIyzSsVGgEbUgw2rcSSMKqKCwQ/rkqM5
vIuvNcxFeXieKFVofLIk+3OucgogOE1bsJpKJyIVNoh+4Lv54j8az9xJnheMjodf
zPBURNlm22vtX2epS9plxIWVv+wWUXeQPeiiNWWkNGvcDFfh8S0VjGJKgf2SbhWM
FOfz+fwFT5MGj0Iy+TSc7d6vAKJD2WA2Bo60EdTlL9hHt0u0/mlE4EDaMsveSCDD
bfZXwj5h0jXlmafQKGuuC0LXSsIYtmbRlshXNIz2AbSuAY+e2H9z/0cWU9QbDqAJ
UrC/LDhGtQuO3EUfXwdDfw1iPCMHymy9qbtJCml1GI4Rh5VLT6rSHN17Y5QocLAh
/c2iYDazNeuYp1OzE4ph4AjYbOlfC1JfCchn/RUKCZ6o2oa9uExP8J06Hkck3wcg
a/ECM5T973cFD7TwvQLJiAFoMvaPNMld1JwLbGZuGr6A9d2ganjR3s3hjlADGHRQ
J5fDqdQlQgs9VGheUGoBukR5/ehoBk32DvCBgeqDBFboOaDmf98MtMXRARtJ+hip
Cb4MwEpM4fi9WDaL5+2TRjfi9r0f7YILeLleflj3cJagHv1obY5g8Bm5ZX6br109
dYTf0LapdtbKVUiMQkk1K9szdQmWeVfLrICf/IB0paHDCl5TSCh0afIZWcnvUyBk
6eCh+2czO8R2BQfAFBvDkg1uDioTcUnkTuSfp6SpNU05OGq/savEzyEf/o2SuRTq
2Jrxv8BDFj9Wd7vWmQ5r2n/2iIaZTI8s7o8Rngy/IVIuuBNFj7evhuml7JmUV/Pu
140sJiLmEdlP7ZG2K9qgj1VpWtUJDEzoiYOjJq3Bnei7XFhucH8m4lQLhhJ70snZ
PjSeypYEGkebMLkeQIfIgpS5yn134IevhuNoiLzNLgaWc3Cu4ulHt5UDMCNFmllu
xohyQdu60nQv+ligbXKb1QShPKiVlU/F+go3UU1OQE7nAL3ZQuZJRraLyJAmjDHZ
omYvSKVvOMm8Ou+0+fvKMOPH1KkBb/FPu6t4qvMw9/oF2XZYRFrg2xNufhrQUeBN
sKm3kZ7OS/cy8aqBfH2lLhq2Cp/M2VBbm6kGhyRoG2ptH/t385/Mng8RomSs8rge
Go0iJkEt4eV8TBQ0pCBXqDoTysvWJTLq6VFr2U+lnPYXKGZTkkk29VVYdGRcHcwR
j2YuI4rEWnLOHWDWQAPuqQUn/fsHjl4v9cRP9YO07TmebzHc0uwJutPchEio5NqC
FwrnuDlDe++lnMafEXw60rbwNWu415O2wA1VgvLYpGggZGm0UQGSQvxif0M8zAfU
A6ZXLNBlNxnAa1RMnki+8VwCLS9Kf20DCFHqQCLxqNDg4pZws7Wi4tFmEuEBFJMr
5OyUEw0JPmN9fjgN/pJ/8odP/BkxLKXLACTKWQOYzLWHCBcQ+vhefOvzzU/GVzb7
5lQXEL6G4SN3Qiv+k7lHm1FcnjHfYtCD35VQ6m5j68KCR2Ofyz3La7srUhvbAMtk
WRpewzHbCkqQc0Z63XspwqcEwohDmoLpZyNZpG0xW3ONRxY0XxUm8Xt/WgOne/B7
QJ/2EEdRfY5IdEJmYI0vhcW+DGwLrtOD4WE6pRNGOu42wgkivRkM/SWPXlOWlqbJ
OQ/hmBL5xC8xOzYn9SygxMSgLnJCwNJgoV95QcPYQjUnGM5LiVS2FUtsF6l9SKad
V7FISEealDVP5GL634tcElF4WlU6h+nS9LGo0kzhzEYDN/3wQvNpBMEXP/4vPKzx
IEkupeNCdfWiC4+BT1jZbGGcMj1XTWRLcwMQOfFZJw9LUcUQkd5qRBsmEaP9kUmb
UkmtcUGvlIizSzLyDOEoCJUKeO16Ct3rzK2mEnVJFVZXZsYUzF+3tpRLIXxDK0rI
mY1+LrJYM8H1mONEg1jWH3H5L9dJkcg07f+b+lw1hyEYDFryYI/Horb3qbuqdGvI
WbHyd+TBwDFrDS3yqQsXo1TmNxUT/Mq7EuJo5yFcqNl3R5aX1LVeD0O62jit5fo2
LBRhpI/elJ+Ps1P0rZQRkKDYyILW6MoBIlYgglUpMhhPX/hAlQhypPS0DrQVqp8I
Gk19ODw91TF9DFILbdUPuMxvPit7Ay4/+AL4VqlzMOlOnfcw7VmwMEATBfP0ed+I
EWkZkEJkOvJOy+2SM7A0OvhDi/57ikNJ7f5gOuzEyszES7xQQr27ezqjz5q9URki
9sw87iegs5ooiRn9n5MqVTfUblua4Ab34mK0FTp8SL4GKNJnydylchFwkFxzh3qA
UzSBU1QXM9N9CilUaUBNbm0mtN3Ep8BB8g+lUAwthK2ab8zsqcfZDPiC7GKaScE3
w+sSXJZjEw06cqKfnVy6HedBSGutZaLdTpqrFBrT8s9vUpSOAbHdNfC8uZ14BZEc
Q/ZghbA1nF+w1uTne8NfLlgdNdd03qSP9scAmkPVGmyqVy2cBgHKNLXU0qfzWK/F
jTFrkYxRwqSgD2T7MeNOo02YsydAnwSuaZ9Qj2qWi+WH0tB3exOG7aYsdnFzVgiG
WkY9nPmz3GC7U3DNR8O3DLUD2Ll6PjGPHSql6wPxbPDRPfl0uO8BkzjjeBc96i0/
g6xaOxJFMP++mb2k29RAgJtRCtb7A+eGExgR5HDAJp4cBabqVTcufYlHBKXzXPsV
2t7e7X3cg+5V4FUtHaMY9fpNbn0dWws55vA1PK2JFMx531rCQnki3kaWhfAjzbBH
3YAv2xwRka7GIiegngAurjWhjZ4cMMeUsnPbqhC07qmB/K/7yXuC+QA43azzgBYo
oOGpKOxWz6VMbhZvFfw7arEnJEI6MJ3wHsxwm8xKeM8R0lkZ3b3U9gINbVFgNKRg
INs/5JmXn25ucv1ntGoLBaRV3+8fu39jZEb6PVri6SKYZ8aTHmLUFOG6JyrDRGpX
Osbs8rOuzkmDTVU2s51yeYdUVNFKjbOKlz7HfuCeRueBnlhE7WgYHhDbZXjP/c02
J2L18wezvdFf1O23vvdcjrNvtqA53ru3IQ+1tiV+IvZeStzjAClk4jZ6dg8AcP5M
frL9Ec61m17A3k7lDfmLkl9HUR1m6KkaEOSHY9NhB2J01gSyr8kQXkaxCOYwwDex
D5vnDCTXS+x0RszCCn9Tt34I+ETobojQ6ItoMWumwzh0MS/Z7fntUcEopCs9qEEP
KSjXJ51dLSNaZxwcfg0dmX5DBjOprQ1YODvIC8qD+y6ABRzk+pZYQdAuqBo9z+96
+gA6rCnpP2u8THRfinwxcUIjT4/JAz1E2wm0f2JMsHPy1lFRxBZUfgyQ6sXrMXkQ
eXKsUFR9bHvkDWaYDXv0EIvWod4nknMrsVd06wiGr8Mdpln8nfZawSHN5ElR/HcT
elAMxtsJag/A3UtPxogZYd1YLvM42Y+7B3cGDoN/GQaJk3GdsaqpMo6RurfpUcuN
QIaTlP+cbUGM4Pwa/fdJAYm00s5pEvLfzhOL4HpiOo7xSLdsrhRh8sYTCOobvFiW
8gxPg6sndGDq8cOjoJXsUIXQ2/n0mIoNJiS/TaXFHl+uONo9lh0HQum4faZBkZXB
gRJ8S/smekJGtCOocllxKeFHONnFju4IDNYU/uHUwXFoZJ4Z5wIvUdhKhtT6QLOF
X4ugxP6j9sUcj8ItHdU4NcdrVaxlQdlHKpdY7rgOknIaX6cH9gFuL4fz45/kpeW8
xMlrBU1JNkdf0549lU44F+2vLOwtZlMbwK2jfszrSdJbnow6vLd3KTRr6zzcKr8q
uEM62csWDgszWy7uDa8oHHAnVzvrJ12msSy1ND+r1zXnY/OFEs0ZtmEJOefpUzrW
40EM/oNKNU9pFIthlrMn7gbEKd1QsfkzhJiVtTlQ2j/9l7L88l5XCtdZ5ERxlTel
VjFDY3yRQ1egd5uMeFqCsl0afBMdnOIZ0RjczG7C3HL401kCYcgZVN+ffeVXYiaG
8WsW780Ih/YbRzYneuQP6Ro6Dly3Bxzc80pKQWxQnFggwbvVpHazMyEZs/crJnlH
t+Tb4biHts5/suREFYp66+BJN/uMB3uHi0EN7tcyt5psS1ajiJhSXFNHUIa5naym
ZfsFSNevMQzqIi7xGHuPLdtSMNW19taV56HWXWXiPbmLKvvmSBFNiHAjQkaAl+4Z
wIHb1M4wYGAwTDjvWa4GJ4HDh8D5j5N7A5jyaii/jVIZ5OZviT2N3MlnbHxyJknJ
eFz6suY6STNH1p2duqxLUYWXGL55/5+stwSBVQ5/AV8YKHk7ooRMrYx9XOCqQYKn
LTeEBrZim6s/SK+/J/ANK0jSGzjc7Hf7uZr8CuIozMtg+1UbI+WdhYx6bu9eR6MW
tRajIOxt/FM8/JHlAEiC/lT/w3HmGfTuFI4j7yGYy8xXDhYQOZX6sSXEU1wCM/Oo
hHrhG0n8F8wnQ9o3zBhj+AUkUvX1mMbHGDtrRJ4KfIxBya3XgLZuAbsmNDcUXZi7
n34ywjZyKxU2zn8CQxfHd6R1D1HzgovVPl4qOjOqYaV/ZiWIXBrjG25FkO79otxe
1PxIrh7I2hSTBp4uSswnQICjbkoNLqyVC15fysKAQnxIyAIX3vhTg15JByC7L9AH
cbmg9EVzEEYwwyjUn44iB9QWclg5TKg3oKQBSLq1JFs5TNXRxTP3MwpGUfHpJ3Ei
AnMcF0HTozhQybEWrcXQIXtxM0VWfdvX9PvslRPJ+URUMylOcNTufk3rS6IjdUGU
+7NO++nHXKdewDos036CBAoqEIH+tsJHXQVBbvgY/g3vrGSb22E08Ec5OqIfVuNU
+p0wmGsMRT2NNsCOS3KqPXddlnkmMXamlKunpwJI4F4KwdNzv3byywodrNjaLkGL
XOZQGPKazTtvaUEZtQ2Wnr3njApVKlrg+RHsKQkZfJX9eCJVs0usZuRe0ZLuYmh5
WYexOaaGB9ZJc2xO6A5nrxua8j1+OI5Vug176JbgmJalOuBzp+G5iNL5TGC+SNYe
goEYGnWiaAotXI7uY8hcrhVzZFsRVf35h3bOpQj3naHYcq+755fmwzCOXXFkAQ4y
ygBIb94/P/id8EGvWtEAgx3fwCjgQJGSVTQUfRL0Sa1kK6YXeaa955zh4iOHnpd0
+eTNLd/lPJ7fecyQFhrAukZMXyo+lCq2qOcCVV+qUmARyKtUY/5THjDCsqXcnN89
TMFSIMRAutMy9NeVh3m122fGa6clOeFyrkRs7Fr+/P+C7k3gwHwCsyJUVH1MpVvv
EjGH36Tb+p0wqVMN+o/Er6jdIGl0r1v1hvjGkcr3NwPcVTFCrUB1GyqmP+0qAtCx
SVKzAqhwTCA4nBjMgFaRnO4fPIHBpChcsVDA6IK5+fo98RKJ9rqvFDucOEiZAkig
hE3kIxzKCwwCtv8yeSFpXG2OoOeASWmkmx8nyUwp2AgKWIKsSkOaJ6TTFhRB6VQO
EOcYkwg7hthEt+uFH9NgH8ZV4woMbAyf8tBO5oXvYG82IFowPI8pC1faQMAMcPGe
pNWLJUUCjOFGssFWGyhFVyeCVlvLsRYRbNPGRJQT6hCi1a8Fq69iqyw9U9nOTa2t
TKavy5u0Lu1aguu0aBBHogdi2uyZ9RPf3/2Ix03QxQ+xBe0vcCBzKsV0IUzCzV9a
fDBD5pPYr8CGopUDfbOuazgRBdCXCek2baklzE4O+uzk25yIMx8kJUMfw2UOwry8
8OGix84leFIN9jtQjgqo/OCy8sY/UHrGhCS62KfeVPfbseQvHOvcWEOD2ZCbBKgh
fyV+q66Zg5km/2e39pl00WeTU0lc0GP7istTirE0VR1Q0zyYtZbz8tAIp0e21JH9
OHZzq+f695ITbdLqDjelTz8C80QbePD2NAW7S9gqeWDNh5QGwTgyG8AQ/jWOko5t
ondA6EsjvoBrb2CrzymVi2/EBj4US/0XfHAaDXv7MScemkFss9Wjr9/C0yfEJ2Dr
nC8KpCEDkj8QZ4TaE0Pho43vhWeq3DuB3YHgL8jzV3AMMO8FNilD04dZDIMZmInG
gKM2eNFDJGzF1ewtNYWtg37AYXwuPgalF5OuDnR3f5r9zyrimdjnK1jjqZL8MGZp
u+Jlt6kzutSrRTN31PpTClzdZrVdik5tRL21TtF7Scn5NSkONT0WT6XqbpfTcu+K
Ss9/sR1kV8WchrzF/6KAnnwTTfl9tpvEm7QNEp1mjdvlur9K+QIYWDr3xkY7yvb8
BRRwf61NKpMkyxLBp6ZqJRIrkg99phUTTOyXDBjRVt9cKlVZCoXEwEXzxgGTMWx/
FKawJLLoGDyxhR5yVP5M+60AfjMrx2Cxh0zKHWIpQB7VgOfohytZcuynO9YqprmQ
TfAmV1azymtCI/tB1eeCBscfUG3+Z1u0Deed3/OubTSUWYC1ULm6dWKn900guggr
Z0mjalC2UI5+dIUcF2saRBZ6N/jiJct+BbzF8bgdrTH8jp7Q9V3fatFoDp0TwZSJ
PrV3QeUhmQ6Ov5smden7Qdbnwv6BWsAWbHQTSSZESNkW1KJGMk7R0ww7zUlTOD4F
a5S0H08nr63UzrFs9zcSeZ2giRDExJJO+ZJ5aB3Mg3c176J6SeXK8AvS3uHa8H3z
SYGKleQIlRZimxGQEm9Xds1PjXqjpngyl7dty4SHpkWIAM9dJnJl0FwGaiWYByXY
dNZZoEmXnvmZRDIKhuZRn4B43cc5OEwKbglmj8N0iTTkxj9x8Fo54g0wEgo2PJO5
M5ahyijZ7EzLZB+wDzkoi5/8hVzwrRl8KJ68P/gh81Atj9wPxL1AnytdP91AZ3Tf
T4c+w58siDl1aCtlidvF7EM90MXtXi9SywJq5QZoAXc11NSG5JGI9Q1SBmB2ufZl
5tRYDess8/EUpCRylIRBbPXIw2LixhsyUqMA4RvbSKxX3zqECFjy8qxARJKx9TP4
UcOpW3x35jysLupZFKsprU0/FgBoSa0J1yglO18lHbgbjYaC0pQGGidLNY74ATMu
ysgcBC5J+46vxvX9G8nhK6VaEj5YBoUmppbZEq/bpqyhWOmtHC+qX2d2StbeJdbE
LB3mUq/+7OixeNSOOGC/Xcl6L6iEk45QGQIk3TJR2Eu33QoSM3uhm7XZ5whrRuz+
BZcEKXbR/xY0r9UsRv9mH4pU1m3t/HwuXT0xvNKA8Pohp6IDi3LqirKOimoaYnj0
Bk9peCyVvEyJRgrv1NkSSQDFylGOMaKmSz9yB1Ptv6Jy5MYI/adcc4wWJvbBJVZE
QSdgevGIo12gIEJNUZHQ2Fa0tjSpRUl4sgdLchuqhYMHbjdeIkHu1xQUnGvEkJJ2
+1AIStOsNguq0rINQ8FDOLyLKsUzuqm7oIRvz+wpQRRoRQyVLn6YRtHQKXUWZPC4
FfJdRU1JxHCn1H9INwBg/7zjCAOcQ5kS4u5GNBSdcjSnT8U/1p1itENLiWyjhqfa
OymKvbjB49rF+gnkzcEfC1Gio+EePywVYupV31J+J9n1oBD8SP8dbJxuwCfXf7Aq
lyIVT2uu77NcATOenQGK6n74F60gab268w3M3jjIGSz60ECJDhSrbBoCBBBffNSX
0kAleKRkGkUa2uwIIZ9MqbvBo4HqnFoO7flOUVDQl9JzkQUcFGAQXvRSnYxSdgCe
XMOM9EMvTAeUh0S9wzHUREeETrBhnLtdrT9qpKj+u/leutKTIS2HhAl3G1VaiLFS
ADV0mIJkwBPLrKLYt7zVjKE3bBta7hj2Uu4x8SerR4ctBKoyhQWNqoGewEnPPYIt
P/H32gnPlYj9CpPwc/DAYQGNL3MEyO8/e0nHNhNqtvzvJkkYVToYLZ7HLAKVMHJL
f8JvHZqQS1UjzA9Fny2drAA78fx7UTaDjjAXwB58xtgqZAnEvdpkIYYMrXwoXNBe
AmxsnM4cyUZVUGus1nQ/5v/6i7TXIXUwlmlSyZGx7Q1TvkP9/wcJQmE3LpsDNYvm
IIR+85JOOWP3hLNkub64gLPPnlLdv/luWu6g+g5KvZrdqIMRThr00dKJLGfOYPS0
bnxfactpmcNipxUAKd+aJUpo1oDx6EKqJiPlOgnq2+dBUbV9YBxCsTh2WE2UGOIw
H9Bz0bh1s9BpzccLFniHCr1bHBLNc7UDcUEQ2OvOtDgE51pvop6//owZ2nv+MXTu
D5qtLYGMkf/nSyHn5k1a1R9ruwGdKo/O7hUnBYYrjX3c6zTLx4xpbYBQ3d7RgZuQ
IjKoWZEZ0YKXC7iQyedsp5cmfmLHHPs18P0H4PqkECDuMBFcvzmhpmMZULn1GE9B
wB3X86p8ZeScyGw9wQVdyitKvZbSMsRTJBcsCcLI8DKDbYoWEUxQlnuNhccCtJCT
gYqgUlWH8TrlNUPhklhSvsrWTVePednggImvEsMX+e1yUIeOzlZ03H2UBEdxh0+M
moEr+L20lYbKNwR9OLUTNhls6yuXxcDDTN26+T9H50QQ5g3b9DyUuPweSBzzQP2Z
r6qe+alszM3ZjexENc1VoW02D/yPh07zaEJI2Jvq2BtXr+9i9Wk4tS7LYrn/4Msy
3IdjQY2ha37KJVYmzuQQwIyVjR/BLV9rgTV+rJ7FY3ABWCB/7yfIthFixRUtV1OH
FN7lF2pLEO979xreUBU/Ik1MncISMLBLzTMYsdJiEVmwp1OXZnJo8FMxPl6CTjCY
2LBRNPEDOx9w5qpANocVCirTnPnDy6gUDQLONomDUyaN7Oay0ZSkXW+KpOh+cZOY
UNNadpUZuP7Dq+y/14mo+o5ioM61EBqYtnTPzIv9/SL6Xu8HZ53xsUUPwZ9NUaop
ye6GCZYFBG+DSpbrMFtMZCO5r9/uNn2gley3kDSsWRvbI7Cvik93Q+hXkjhaE2Vk
PC2Pkf6DmiHPWVHasW68k5sqPqUbqBAAazqGyULZMnS/jl3V3u+/VBinoI/kRyeC
NIVpuuHJM7Us0fgAj8Ghh9VMehz3JiZDqzTFr27ZU0/irSrmQDiuwi+37Knx17Xu
bcV0rlj7toVwUCWUhdCXT0k4ukTygmU7WyryYMHj7KCqwHPGUw+2fAB9EbuIXOTZ
D7MxaUfQqYKLQcfD1FXbJ9P8F+ixp+59BcG018a7QbfWg9cgWmYCkJXZQm19lzd3
kCSNfRDa5SVnpWdekSm6Y6rq7sYttn+OsSvmy+VulNS6iBe0/9qr8qoZ4GL0YpGP
nQ1xrI+a5zB+PR1hSVZbJ0oOm/xt1FqboVsZyt4Lz/ZRS1+N2xX8m25j3eFKSqUo
UWStdcA+fqBqpz75XnN2w0yh6fROFYbIXRytOX1WTg0XUVvfEbyEnlVjEakbyLj6
kN0B8UfMZP6WKMK6HB+URmKwoGnzDTynx1te/SSyzi3UE5ke7py2fymUmw2hoQR3
6nDLDD81oqwALwRD44hUiaFwqmgW7SYvIknpULfPkV0GgCET38OvDnMmlU1j9T5L
9The2CvwCpnfcJ42j9ZGdzGWQH8n6rFAUBjSKlnZAkDM+jGS9trEHxikp7F1sQNm
bpjfnrXpK7VfDBmMTIUIxdBL0EmBqDC3sZPR7PADCT6mtoIUoo5xUvj7Mjxq05pT
9v3pO0d28cNUk2E2rUPjuZuavywjYZ2+Oeuo/eSxSs5oDDTKeExfyMggaEcWryWc
WtKdEQj+FpmNr+CHd58ADV5C8688lmNLrIdaAv43+oMmXyma2+Qn23ADvqYLVT0h
oOnjnT9U2u8dKtCRY7y2n/GZOLOInFLv2KaGtAvyPpst6tS+xDV+gBge24kLC9WK
jTLmroVPBSZoIEcE6lmwBYQGtMh4LLaCmpB+KEhNQ5Rpy4cbTTRs+cyJRkLDl3Pz
X/QgqWJh+dze4Con9GUk++JcHJ87na8TBOJeGlFnFSNaPLHopzOviHRTd7yf4B7V
V2PFMaTyvDBK4nJrSNhSceYxteYSzz2ZD6LaSDsLj107N/z/+dDoNmP8J1T72Kit
Q/H4dsn7TzU8+8SVHWT5s98AB/B6dR/xWHzicVtdt+IsdX5UOS6tzwa8hKT9+3QU
gnIc9tPpwfwBpKN+hTx/SzKj0yZljyEsE1tLHsLwRCE8meClPE6JQCcFB6Lt1X0g
niK0yK2u6SrrUJBfM/nFrPvaHT31XcwkEedFgPoRiN1RncE6vc9Hb1dGOrWvPOXJ
haqzvjJfvOJB0R3CYocSL9fX1V/R87B17QfKbgA842ykL3rZpXYMNOZoU4O4qk4L
MP9vgwu0a0wGCqmGaVPGv5ivDIocjnTl6b40GgdjBblYFTFWcAagIUb/+k9+gAJV
dkza5tLXkK2Ytd6CXX2wfDRwQZYb0JZvLkc1Saqn4ey5DjzB9lrJvt8UdFvSZI/g
TZPuE7RvEFa5p3Y2Bc+ZtugIrX/hKkkKwJJ4vKHTFv69PvN0UhFwolIrYDHZM8gf
U07U9VXQRumBY7IOMY/DlYOm1mv1JpHjWO0utyFRLq4ULrDd5i+v9cUDutpcv7w8
Uqgj2mh1RvuZa+dzhNL2XYE0UjpUW00Pv8MgKJGi3zd/gPYtqAXquxIrZN+/wV5P
6ys0PC6FqIF3ATHRkzlUKFAPTVfX3mVc1BWfesNMP2Znh1jBF03gyuvFHfqyhCsI
YVqtnxdQpILCl7D1GFcnkKOBDzBYqcKutQEwkavfZUws39KSrzxAZyuOvmkMs1Gi
9nE9+pDJ4nLGEb0zsNkXzdkWYI2KSFBCZalziPFHbfjvuzdB596rW+xOYQKgM8HS
xn4ieXmYZbbtu8ZqG6Df4K46FQL3PAHdkMHY2VRbBJ/CFjiss+w7QIBYZqj+CJn7
ofZd5a5upQgvXVXs5nAp05e7Vn0Q0GjBZY+J7wfXiC0g9OoU17RFsGY5tK2rAzLK
BIqYVqVx2IFbqnLlgttsXMIWIVrDIVw/wExP08K1fQfbvC2PlRJlCszsIgQTzIyu
/nfSV48y8WhpYfpP4ughSqgM8AgU1vL3c4IJvYyPI1HyP+uLFzolaYSUPQncVyo3
+lhqtV6OtKmVhUSXlCn/XNiks5ToZgc48x3dzRC7iH0y/K3jvcH65mBsZpoU+Je5
wO/AhEwl26D+QqVkRrwlT8aMmOj3s451NznWs9+h6k0FQEgdRqAoCQDeOKPTt3cs
kvM0HXwTvDCsTprTFYWYDLbWECxccoKxUtLonSdkpeVQbNijWm8Jp+DwwMaPjd4+
z4f9/YfTCiawlA1rIEdKiJn4444p6IshwM3QJxpHa9ODfEvP0JnSos03+pkyxR6a
Ec9POPb04eaY1HGlCk4ELiwTXFAmy6ZltCWvzW1T50/o86VDd6BvPxSNnlGwGxKQ
r+WuMuSq5k/hz0M9xQ1P+ALiRueT4vnnBuhBsZn4mXDtFLu/mzn91v4yyXtPlnw2
58zaP113qd0bec1wgS7R8xbJWRBkXdBSOSOJHuUvymosxxzFUBkKP7SrDx3mOMeT
NxQNkZg4EnrhONsvdLFpVlOoivZIvMqki7la/2rO76PNvMwVKV4F703HjSuZmcBd
ZJPCa/H56WiIfy5KuUKGb/GCJ1pF9j9Kmc/Xgcg1i8QypvSOIKddC8zdK3JmbUu7
SgnaGRIg/uLPH0iG7xkwvqlC1RK2915LIEhYXdGGGY2tdGuuWaRjKbExEy7p0gJY
wlV4MvtoNqlAwLeFN3nXUYwl5Coy1GH//myb2YLX+QDjVlvEZzHz4945AUktUiK3
MGaDi4fMBSj+NMWYCn9aahd4xb2oZz0NLEXrPTD+zJNaaTi2NJdiSjER3+K6OsLy
hTAvFB/Kp+tvrr6aDWA73dbd0gQ555zI+u1myBBnQytPbDd6jlJ1JwNydaxgD95X
DGFdTeKgjkvSi8kYBkVUUE38+OV7IQO1vxQuo1objWlpiSvj6nCOpX90PHoVcNSa
ysbK17QE6hdJV1QvgQDShKuaJKIP9c01OmBufYKfVy+4yjuG/sXvRZ7xOYtEjRX+
qZ2S36Oj8DAdWByRdTD/4sdv1eM0zM9xJGOaQ0gXaymw1hYYfFGpTPlsw2jxUApG
oeMeZaVCgyPChQxtmChHUktlkdawgDf8fFG9gCMR9ITURHltCOZY+TrJctgG0BoJ
r6ghYvyHmuWp5FfteOsN/Qa30yuL/C4aeLhMPi8yzDjUVFqHHXTCqOLedJcEeC4g
RuOK1SFiWryop/iiT//Yg9E3LUE0heRKmeKNdEghGHyqOPPTlz0Do8TR5e8qqPSg
VIN6PhmxU6SbezpuLYmr/hbYPhdXWxhachaG+KyQF3yLLjYwBnmmtFK6nlqUYLk7
NLBfUW3Gb+GvF3FJ9U58VjjBMQBt+uUr2II6fCn41vUl7Aeqo5frtQbGz0SehThu
zXFrikbG/q0Z2BfFj1HV4C/NvLUtQs1tFKJKKEmEGmsOQBF4ybJg0P3PKqaKQ8WO
BQasIYkTfD0KWqlBlOsvnp0w4NcSisqEviPBAsoJ0wSvdXJruNGMrXpkwQDChPH2
5jeCObjAszcekVMK8ZnAEWApTmspkVR3pzgFYiN6ZuvyTIgYDG7XfcAYUXb6wfzv
TdGvlsPnd+nf+jxrR+Ysl2+KK1kOAr7yDXzjkTt+TKmxQdSYF2VyJR1RnEgU8fsO
UngwthujprTyuhzWKTbGzQ2Gh29z5WxHT4Cmg0UqYn5OJI8R5nyr1/4YqV3ePyQn
DcoenpUqcJTgcxSKIgVHBUhFEL+jJqrg0y2vxwzVQ5xcMQr9WIdpubQIWIOZkjvp
Q3SSPn6UJzmeDj0cW0lBkoPL6C8KOLh3ogbrshX4muQSwlG5qQG7YP9IaSRez42u
LylSYrvcfMqVjQKIBnTLFozn4NGFRuensojFvL+E4h/RYP9diPfs0z5qDf8cY4r9
TTULywgXm1GAFOGYEpt9tvVOCv8sSfhK+MA9dE9zICecXenkJDXGzYNi8CK8by6h
kSvJ1ONfcHkLAqDQdPAvXByohRkmHPV0enHklmcaevjNGDuzdvYGv/qpZ+s7sa4b
CX+7H7LZlf8OJS5X9xXJE0K+6U9QUqyE/aKgkRIGkly3vwBPawBluXJUhAe019t3
qGsBBgNCFYuv2gJ2BTApsjADUB0tmVm8EoA42s+FP+VLc7IOZRb2csty2OTvwZ0p
vNtxo9ZSemtZPh+CfzM72DjVp4STN5AyvRY7AZ64hZ6de+uf39Z0CD11iffgzw++
YfW1vbusDMqa7BSNT29p1sDC/yGWM469EIu3GuJdoDg67LQATzK9rmVuxjAT0TOl
c2+EvDJFPV1SZAdrn+bl3QEVxnjZkUTW35GyUu8XEj2iYS3TcZc/IZ0esM7OBR10
ppl/bqUSDaZ0FRudSuBC0nKcuc1ssqwYL8XnudHX+nNdsh0rerd/WLy55veLXHjB
ZK3wn8GozlYNhFopwBV82ExwpbYcZIA2YS2L7sP8f3+7dlaTgQHD/3I2jgaNybHt
WedafYy5KN1taAjSlrLc4D7XIKw8pJj6tY9zn8lS/1czsMI8K2v95nQCxdTCXCrn
umGsCNVmEx4Oc0Tp5bmjvyOX35CB9t13Vi2N+vi6OUv/QxmDOPjpz7eBF2b9RRed
cxn4FPeJhgCC6i6Zlo8DEjsFG1OXjF+j75OumQ4+dn3gWIwqnDYh0PGwkb7TaFdz
uip8SIRLa1JPmbIOfbtl9KBIbNqPsAJzUD1IkAkT0YZaDHfBKNj6uIc0KezSC4YD
EJfpmeHmvJF1pcoP/Hz75csgthETPQcvdFDgf6mTWuKydAG9A4IHPGeyUS0FrLQC
OkJaiDd2+rfu26a+hGitG6lci7n/ZOrYeGZsqXfjTR5DtA7aRNl8NJU6B93oQMd1
UtAUe7S3P+Amzq12upMXUQqA92Q3cbMSYLnPBvwUTFlftz7j2rVECwcvqus3l7Up
X/RKX9YaTTPtu7H76XAAgRUI5Tmbc0Ag6B9mz23m4jP2PSsFBbN4xm3fKq/QeaDG
aOoRdnhXky3W/3536W8P84/AQ8GHWmu9Te/u3Q61qdu4ckB9DjRQsZCac2SwP6z1
PiNVirCM6D6Bssl8pexbE4wj+vaGmFRpWXp5f/fy0sxLC0Y8qKuPCb93Cqi1OGdB
2Yl5Ams9U3ac6Oik5R+MLbzWJ00+PWA3iSTcvdIUFNuogS0n/90qXbBFFU1CmeGV
mOcZUzjf3Nt7OCJP24a4KPzCNk7oYlkxvlgSMFfP9iz5Z1tycBaiVuf9Yzp/kjpr
b/UalMD3Wi0p+oQFeID3cKwGfdd9foIQrudKWHV2Dwyp9E5nKoEsGLWfhFVzi3+8
kjelo5xKlzelbHu4bnLkPK9vlCXU7JIT2XpD41Lppvva4o4qGQPKC4MthjiKG20G
YjBCNMt7OvJk2yksOhojiNldhYZS16bqWHInJA8dyMS5Jr9ZNsmoJERD9VFgkJpN
1c/XLZinoKfu/gErp8TIj/2ey4vHsRgBAqKXqFPnBheoDgxrnc6vuW9XxdyC3lZ7
nOBjVxk58nDAtQ5+On8wDcGRFvZ7TahfnYFw4Y5auqQ6MTYnMKDwmjIbsTRlIaqn
uWkfXNFNCtGWMqF03Xdf9G7EVrmxeJhixUBLaxk6Nh7YkUlffVcyY/9o+8looaXp
DiKIa2BZj4/Qg3bFD9EKfBNFMEyHqPY9oBrba2r5Av9sWVr5munLbSIyoS2gCwSX
YxKdKnoDjY3vb3Vw8ngYUf+PwOjV6Id8QPjR7Mg56jz63bh/FlMAgdLJnSF1jjfc
xJAll/QsXFrROOoo3qtnkwG4wGPukHs34JLDtOVXzEs3eNO9mGbxbR1+of1Ej2Nc
Y/aN7LLjykJHcqaIj5SbW7YG8Nkiazp0q57BLOt2Y3tkyC8FxpD0pJncDy3DFH7v
WjdNnp6s4PnR+cCgNLVF9swu1Fhxjq4r8I7csOrjnT8dHQilYinwtwxF0EX0nHP6
5zFclwuUY6Hwkz0PapoG8IuHnsBCgUnawipQ3fISBjV3wtDQnfCm5llfe5A2e4v+
p1WXF5PUkjEvz3u36k3nzWTWp6GWHC33xcEFz90HOwsYqJ6K9Ec+umVxJK4nSxnl
X6ddc2oJrOSFbUEeCkjjuxBUaoi3NV4dG4IGYBq8j/Bh3HgI5uLeXFwZbAzzpayH
GWXVpQ++o+wK88QefH6RBkXlDL/r0cd9ltQ+cM7y0hGfoZ4xGtO54RQcAir3LS72
8Xh6hiK9ppI7Xbry26EaMZr+kYf1r/aB+QX0XC4Ma+0BizlkaIJJQPNUI2Pighff
rWVWOlVKoCPIjBX+9dByj7cx2ev3NQZ/XhryhGqT5MQReGnicjPAWTvB0jNNn8Z/
g6lZ5H9VsrAeyruiWiodE2ntSgGkmuOXgEkshB7Ahi7LTGe58aeNa9vtKPOH17tc
w9oast0I5GU+ULMFWnm7VD59q7mTrUdvZoCjqb6hNZgYU+kB9LRsNdjVsrR/qDzE
/MZEOzQayuCAt/3uWTBNwKMhW0Hs99DCYDorsmpj9CWtQHyawf8FVdL6WirLZq3b
64N+ZcGOKoKasRD3JRp/r9WaoZYhW+N1Ojy703h0FsQhvhFx8LKPS/i8Whh91Rzk
A2F2PJt6VAHwob2yCIhC4UOJq9Y63bLjy9SS/99oV4dZAWBcWdKdqwtw0OdqM2Xo
dwpYNwJqG2b0HAgkXnOzgvPHHD3FeT3McZ+Emfkrrmt4VtGAz8gfB+vfMQTySyBx
dyt7mLU3K0GBa1XfamM8E1tJvwbAJpzMHlUsKCJpZhrrQb2OwoT3aymSCH2zbgny
Jnk+BzOxZmsizuNdfESuQbB4UZAR9K22reC8rzul6S69Mdkp5j0BUc2cy1DfDrrL
NnrzGRDzzuP1KXnWHU8UYfdvJxu21YE456hRgpPUQTrUdQwt3uEZtL3MCBtIJd/o
3qyht96A/59nJCVmu0139uhc1hlk5VLqFToyzd2lOlQBzv/PSqxw2Ua7Krd9dEbp
qJMDErUN0ZmMR2Oe1GNdlGsw32LMb253fW2e2v/FlKXB/QxQVcHbe7bXo1zqMxHy
FyuYBpBHFHtuYofXNdwrFTBRF+Kwpu9GxhExZ0JWLcmYBfuR71WfueBwJVsT612J
xF30p3LCrXox7S/vO4wrw0PXUnGljIpKt64/XMKNe5o3vNFpbcc3v5ejKmFAaOdM
tzzsIkAXRzwNAO++cpNtHdvI8kzqOuO7ilbmvOlJAM5rawwZr+CBZjM+ccmbtbod
pZXoI2nlNpSy3yA0UevSRlkmGnQvoNCWA/lmy2JneOU1wCqs7rVtYfMyMOsGSvH9
tSy27z34ZoSxivUWGr1x+KUGWYHsqPFuHfk2qRrKjQpPM5daRtDhiHXWDebQpWaO
FPk9jd2oUE9hxJjlPRFnPwuWiKmOKsiJnATUUrszLl88QXX/yeyvw11kzYZ1MmnL
4j9DVfQJoYOsLSll/UgC6QhwLKwDEBb6JfzkgfH1XcYEFYFUx90Qj2/sVadRTtvN
SLPvTAQZEJQxBLCuQCGWSoQ6DKYhGFOMMlSSnCm/rxHaW27F8dtLCEwEjXI29cL/
YqNSEJqmuJhYVvARgW6GGqE/ieOtdSnHzgO2Wz8ScYfCdOUj+xb2yHx5nPqatbI8
VF63+ShWqDJEWBeqUTlXtF/djBmsnEtrOjseJg2/jflNYV7HplGOFbdeADu+X7Cj
bQRAHA+HiJ8Km7hD/JWkxnA8HfkYBuKuamctPl8mySIXbHzDRPDvLnf6oRXmGRpc
Tb6bSBHlnXU1gjC59eHEenP5BPJ93X22cNHoh8z4DtlmugYapxVYqOpj1sPW97/Y
ehXynUKxN7uO3gVxHFA3vHhhMejWgW4fPfzZTVFBiMOcDhCA1JVot1g6ErXubNZA
hy6ze66N2cD246fLdfSuYDjmTdb4MjK0fqMUmPXHNJ9gML7q0dIAAz6xpdmWaaYx
yHSEBANIvtVWPBF5DFDNTbSyy+kuux8+Io8KyjN34xoUrtFGunuY3H/gJGCs7Lai
VO+f61ZC7H/a5KW7q9719KTgf1js47SE/yzhSa218dfOIejEy89EF8EgVTU5BhXI
PhobwvSsQpzY3Xrqvte1t09oisu9G01AJtUt3yxBbJJH6ODuwkxdyaz0Nk9tcNdu
qJsGMuMxl9T5Y9VaKCrT1rFomsC7qfCG0/fGoUuxaL9hw/4xvdBzcb9AX9O40noV
7+YkgLW5s96QSicI0fYvcTicyXgjqB9jm4vA3n+h7goPeg+B+cMNM7a4eue7yFqs
PDyr6Wue6Roo4kOBM1CHjLlQsnE249am4SvUTK/cUeFgXc/ZhMVerjd5+g3jvKHY
+whwqUbwQ3F1wZnibxrt+jeoyTkuD2VErOGnTRjQAIB+623Qf6zxtRlhtrJIj3xh
eD7n+F+GgxaGSFFhoDOAzw0E9i/X2n7a4fCuFXiRPUEanDULU3iU8pBufb5S9Hrf
Qa+1vmX48XGra5QG0YpvfCYkVqZjBzhwoEy82/HWWuMcFqmT5sys1PJR+2zLEMcc
Wqqb6/9ewO0Yx+7OCgiCfKQglLwab+mRqrvNBLjTxRHEua8YI53Bwg6Kh3quUFCC
SThVgvND6+5xepQ4Ia6S3kKILl1E35PPdr3FlVyYMTn7cxbGB3ihQqTIfS2MiehZ
PBiCZxC9qjEVeiDcaofzEBf1svhBzb2rhB8wMGbFzEE/W+Uw97v3bLQpSjyHvHgv
5x07g//u3Su5QL2i8xFSOrB7pWj7O6+zlROThumqrDe5yz4AQnw7yOYIIpdt62GT
tirAOsYLc+d2GuSdJk550Tuomhcv9GBcXYTMpWGFErwVW3hIkN0AdQoX87MUKsm+
K7N0LJXy+n19sGiS060PNLrUI1FU6TDrZa6ZR8HI/yAuexixCFNBQNzgTcwbIKLY
27+/Rzz5HeCKc1CQ2fCmdAgnMPX5n0G6a5kKbNvFPyMsOvXAnQK7lfqSs2tTDWrd
JUP6LN3g8Dpfn8BG8QCpzAShepvJNhVUJGtnICvXCmNEAjdGgOKnchA/xRHURXwS
84MKRpSYEa4PC3Fyf1z1GibdwXGUjMGAh5fZkFjjfS7bZIPnAKmFgcIAmTuCTI5M
sm7HwLsfJQvVrLnSQZV6Q8bLuZZwlFJVa08CzXKt7tMpcxQPyQR9kn2WPvzLMGpq
XTifm6J5DGCkZViTW6GU/SrZwJGFFaH5OBTiAjysH9dBuWFUENEIT2AWGs9m5P+4
ZrWoVxyksz0bPVcNTnAhDOOHnhQEBhhnG3NAOHY0IOlXJGwgvJFKp3eLLJ4RBkfA
KgYYiGOubGuJdGyTRiw2JUb37r/EEN5fJTfFa5AIJF8BRXHEzLZBoDI075E4HnIF
jraFQ8PKS/HLcgXmV6oDAj/DL0fh+yeCLzPDBvBAzem8RNsAYXariC1iLU5SCflX
4sGwN9XHou708XA/hp4XX2llE2dLB60IPgj4hvg1djSXYDJ4MXJfOL9YbuRF9oJW
AKF5Z2I7sHwdFOsMH2OH+R8w8pU6eY4odNLSZm7WMSNtlDiWS/Jo4Fo3lsVWjf5R
CMIpz4GJ7Gnet+tbtD4jkzp3agDxlz+OmDU2Uwsm2IG8+BcqStis3hvfMLh80KN0
Xqb3WR7r9/+axIdGezcXXGxMkysKJRL3pbczvAwovM91frcLUOoF50fDYkP8Wpfz
PdrIZAgES1QwYJ1MB1P/9mddpshiM2U3D81TA30+o999eWGh7ceqaKhcGe4mE4bC
FHunWKTvjDp9vkD9qZ78g+z/KSVz72TLDWYy2MfO3pUSGGQ8KumyLasyM1LUesXb
TE1T9xqgThiInhk3ukEmddBIYreKcemRKqdaiv2spkeJw8mRzPZVHd48tVDvFf0V
dWc8Ptx/VKY/jNinC3jvUf4yKNi3M2oRaHDkB7c0OG6GmdvVRJEv6dMawqxlPNix
jcqCJYpc10Tvn07daMxIPp23txrr9Vrzfur/PtteR9JXTlsrjv/IpMoukGYg5Dgr
6gx9ZDOPGfUx3DmRRuDP/9v/JpLKXbYmRdiffyVNyqP1jHvwnUWVCNFLWdC+EC6Q
6F85eOSK62pIlVPPeTvckGiOoZgOMaTi5SbkJ9kGMBg0PGbfOE7BlZxpBZDiog8Q
b2XFDVUleACl+bNMb8i9ZaJbArCdQTNgDhuInbbmJfr9OZmJuC52IrsKSyW/CKbi
Nzdj0DFEuHPIOtXYODvuJYTVsh8A98AT5whCxNAGcA3jZgJ/D8g+CUeAhNPW9M5N
TRaowuTkgb9rNe5jayVwRuCvoa32VOmcCyAbQHRSZKdId+hyUYpGVH68j+CZkXQ7
oPAbzxbm33CovlM5aGCMRWHYdXmGzy7IdtK6OskiBtPQiV4mGQWPYkBb6UjnI+fQ
G82LYe2bv9Ppd5YHVvGQRjm53h4QQbNq+FJynayI7A54DhUAoYaQ7HE0RHfyipPM
RcPV8e3q2VpW3I066V2NyplYQ8ZSmzbtg8BLl3XKJ0TVoAXL97L7P1HXcFqPkOiE
z69fP4JzqF4l1MHDJjd9IZt10DoqwIEV2PQdnquBcpBFDaWPPFiDg+Q7tI/qqCuE
Yym78oKrYfpHmaof59Jpx74z+IGZwzavjyQv+QFo/i+nSqoCQdVYtH3qRz1ISK00
daB7X5D6Ug1HN4OlUZKxdQ7ZRvvkiJlzvl70yjW8tHobRnKXuEAYmi7vxuUjf5Xw
MXKmScazGopZ/zvIXoA+7wjK+KbzgNRwB7KWlhjrskVKgwakpaCvmZCGXadj8Z5/
Pa895CHKFHL2LGE87NO9h4e8IViehG14nukBU8nONcxdZhLOZKqPCeV6dWr4I9gS
eLUa3vn38KkNzoRASSlmhb3OUsP/hBBYwzdZLHQXqAJHp0sUh//y4dWbs7rWLv/i
fh6zwTmo8HAFDFFujUDjRh53/49MP/Jfr37dmN0KECJ8A1GVcGZGiK4B1YNeRh1I
cMbSZxkgn6BYInvMIE2nVHFHJR7FkJfwHZToKLv5ocFzuiF3/sLFXKVwv9AsCoCv
/ArEo12AKElPTuJi8jQM7Du/MVSTe7zlYLUIkDqYSXmccNVz8vwj9l7LLfCdekZE
SHKUXoa0KdXN9BUr5GG4FXq0meIKYs40oVAJKfwKLZsR+wfZi7XqJNnbxoAUw4hX
zCyzRrJzMWHfyNPTHAj+Rzs0C3BkIjZwDax9geTuHw7VHr9S+LLeogBqVDbN8xGw
IjUyqFjJl9MkFYoLcNgZZSNRnE/LkSMFoNqJqmDj+kbYdxS86rZujjCj+wxh9Uov
KzBRYqC6T2SgPZTkvxc3Rf9VF1SDSWW9BdbVR2NZ/qwn9rhABkTN0STdsuCEHSFp
VNMR4KQqQE24LRyDodtBQFpoYA6EtLv2Ju7ykDt4wX9VpEPKj26uDWUQkTk/zg+E
qnsMxpIFQBRBmBD7OVaWGnp1RboCyXkoZdTTJeAGtuEB5BBpGSlgb2T+KAfbvM+n
JLE/karkRNSFK+DFq+2e7SRZ8A31gEOFylOIRgqCz3Xic8EAwDjRM1IBxr0wUCgM
oNUrp8GWT2UXEjvVA8KVbmhEvSokCTA7Hz7SVj/Q1bxCb2MAVimrvTSXWNvxNxTe
J9i7M2uugfwjGjZb60OdkHpmTfrHPgi0LGNeBcnozB8rRTKsGWnnLNKnH8uYsxEV
B92Tuyi9j7+PVu/D6tIuHsXbTpxEdnaxr9MTkAoJM6f0x6+nFqz8lxVE09lNa/6I
R35A+ybhhZ4zrccphdm9YmMw8oq7tLVSLgZN+GFGgfC0O7nOYaxpzVQnA5yc0QcB
2o9Hq3SKd/ZZfxFkEb6qdhTVojIgQWayqh3n/sN6PDWvSKgMpCCeVgBesHV7KB9c
vEmg9KocjUW/IOWLl4AxOK0ZWrDHjxbSwMlgEYw8zjAwYzFb39l9gJ9or47PVKCZ
VCvK2XjWYp32QeelR9MKIIwF38XNRE8OvEylZDX1KQiH41mnbDUeotnKXY7UQKxq
0lxeNuZkSroMv4wBQ81/iDJSazzkEfkEU952wUhyexNzcAj1WhoQ3B29+258CrwH
Dgm6prOKcXtBGiDP7e5PPICOVwKJ4ai6F3KvgTSuDu7B/DnUAfckEWFqWc4isBWX
nBFfC2zTLEiK+/2OugHpbe8DmhU1xGcYmv2oLUFsZt8fsX9XcRHmd5gyf4lJABIe
r4ncEoOtE5/IwyUXMSqFGirB+ashqIySe9Bk4S7vRlPtjUTcygeUjYAPiChh+CcF
0k0NuGwtEJISMfs8yK5tR+OBf9nWXqUqN8KlHDcSAqONoV8JAkQyqTzvxXm3mTQ/
JwYBqyiS7QHJnIclLdpG7uluOV5DSX011OjUi9ULwJYl6Lmc3fql4B4XfwLDGQ8q
LQ7eDOcqe+1GZyz1bArs08gjKVHl6YTa0SRCaZnqwKP8DC526BzTDp2DqsRvq2XO
Hgr8Rn+RHMsj91zOiUi9UBJYOX6M4nEhQfdDeAPo74RhZa9lJgqQMRRqcBBvO0q8
lL3I7tbQ7XOy3eqfuCyjIfZCzwWpH6tMWmd/mtISb41cvBngndnImymuYu7JAx0e
AMmUZMnCOl9+gxCh+TKYg76wha9pynqs0CMAMce9r+fwlnNzwQE9aCFiXZZ4fsOT
p2ndkB0QBmRgGnj2UPLsY5k9BG8G1CUr4ixxfRdt0xNhPotJ/PMwTUJBuQXYf+Vq
KglphyjkpR0ObhnG1sMplDMURrP2meyuOj2bmyuTun5Bv9TDwcpDT1ZuZr7A3P+L
kRd8E/Ljx82HNlQgxYFSBqOaLuOvb9qjXVo718Y2aty8URhA9pEWARl2TDvFS3Oq
Bf8xOIEACC/5iUFYs5UxCOiqimgXBtLRDytqKkkV0LL5owwYAA/SLdaVyWJE9rNx
yQzRnnuQ0AGUqkAtutW2BbE+/hGbjLIrMznyFTvZs0YS7JNNXl7LCR5HMeDsT4Tk
CFTknqMnP2CJiVatsWYBkwd2LPmrgNV2KXUAqLyvBu5zqGWOflhEsa36v0q00ooB
CgPhI3iO98hnej65itoqWU7JfuD/GPviXSq5TInMjWVpial2DdTDJUXeJoAHyBxu
YQI3aAoUFZG+O9J4sUGDZoktxmMwZhXe7Df2524S5P+/X7buDy2WRTib9JAi+r+4
CGneUAC6F79r054pUcqZwFBRYqL7iMXAWSX1OuNfdG40jM+H9CgaSMD0PBmLFtR4
jw4Jq/qQSaqWmFN3Smfwix5NTCWoOZ5sQXkRM6xopidoM7yKAseZIXhI1PBLIm/r
05V3jVUH+s7YZ5CuQvTgrq7PJlgqIS+JBCJfJ2gKOWArDhVgXt7sSNx1xqv9b159
tLvTg4OduD5HVzwmOSXAYCIAl/TKqBjDO/WRDQbTzHDYGSraYTHHy+40Ep+MzOjv
+5Lzk2/ODA7QNBMAIDaZ4wGJFx7Z9QiIZwQHLWU/1jIi6Zi450m1xRKJkAWrHVcE
SovpPbI9Z1fUkWiH6rlA6lfBnBqqpmUqUwidwbt++ta2LmaHATHTrMd99uSULbSR
L1AhSbQV9SfpUmNNn1RsHEtgsDnpX82pJLinTHhjxX1xyKxJPIT3/y32ClBRDwQE
57783m/M59zVMONzvSv3J9xtkCee0gLpnP5shDPxg1zNwR9VhGcaDwBtxWoeDfVZ
LsIPnth+q/aQ0cZV11bwzmuvTptpErfHJs/IyoIdXipAO/rJMQNBry/MF00Z+sus
4g7kwGxbuvfZo//KeM7oOLnVSglcqqWs/xiagDGaKOFJAz7BjE+Gofkejq8qW3p1
J3Ak0R1DoYa0K///aWylLRdIjxCLl/z2QeP7ODQwjcfGbJKLGBOXOGpvOarR0rQR
lZYqa51Emr1i6mereS8/l0annr074p2X1e4i4NpUaB8rGbaIZ5zpnAM/ald3J19j
h2MwXQErImXx1Z0v1UbtHAAniEbASgEN076U+BiD8z3H7eNdTaIU7VdogrG7n8FO
Nh52mkg2uZU0RO55SG1ycdRMTQthhtKBYWv3i69ZyGCHCAY5ZLdauKlwgz9laj+Y
AKtq1010jT8RWNkHCJjqUpVV86q3YcRdldEZXn3pH0FnQGGBEnJA3zyat99QBz7E
aw/qWzXTn0Ce+KIXL2TcYxBdVKkrh7rbTu9UN/6m/uBXnhKqkkFD19oZdks1HSwC
foRU1gYyx+RkY7AWhNTQkNGi+uJJWxy1ewinZdndLEUrD/MUv1IVK6il2w+lJRgF
OhxESfVeCrqDgMbZIUPXgtr7wshKoVM0v6iTpuB2lgSB+HldpEVDERWfvmh5hPKP
CTurrwbZWYXJuLUe1Onn829U73J765ZBFYEpc9VdNQZnTMYe8BTkUpylpBa6ZBuU
ncHypSuABI8U8LOD2mqsdQeIY6vrd1hYRrcalNwnl/o5750JKioe6wbl/lAycO9O
5TMOB5km91gbO5FUJPbDVlBeUUAKOxIaSh5DpMRaPVHPNkrfhq9gXHAqUOmeHooN
EVPpqYkTiGSYf1g9j1xIr3czDc8NJGOEFBxLalN3kEjfpI7uay+3dYPb+w7eMTD7
0F+Y5c7j5Vfpy0c4O/EECLX34/szkqRA80stUd03CuOgOmLgnyJA6b4Y53sF6G9D
+vYRw8Ze4+IH3PLP+IYodrFfKrCpYXdQwqdkzefFDiLafhToKw07t/11on3+zF5M
sKHx4RO69TNuRJPEvkXBCa257HUbkRFpXks6uJ6WaekuldfU9sj/NFHRNsXaw4zW
SZW/R/5sWqWV5a0nInpESNbMVsEnKVQz1ghzP2/afkpz1TITyVEM3fNMwhJ02Alp
g0wGPqHFMiIGSvokL7Ox4RogK0d/hNn/NioeCv65f6ipOci77j9kWG887ig6DodE
yfyB0TMNoJuHjs8DYXtrO7irocbNF2xEQuxfl5/p511NIcz/FXQYhgyNJxSxCG3i
KT9H8tl8CjOafnLR8jhxr4epZRAQAAGha3lSB+Jrp4YC4HFL8vR/Ee9mLiC3PCJt
gd2Tb0K86CaWusSG+RcZkus0MTUPJd8ryA6SGmZ8O6B6UJ5BiWFvr5VOWIhiXqP1
rVHn15Jgbm5Fgwi+WoZc/Wu2WkgKtDAgKdSM7Yo09GX/RwzXWMbTzWGAeqQByP80
89sJagVVe+2yCuyIX2SqB5ISoXn6CpszYcBWgKAhVutSCdVuBwC53SxFdvPTN+U2
utkV/pl5JlgYGFD/4H6dmBkrewpsxMG/I2UxXPlORCvYcqdCukGvEhmetmd4G7Ci
i/Mfw1bjT8IxNet1xHhIAKa8E+dtCJbrJ89HL+UCZRKD9z0LA0FagVEqbmqEwh8t
+XP+43fprP6UmdvvMl+QIJ/86pfJUaN5S7kkSJ02UmZluB67KolbpBOCTd/xHzOS
YygMnTGxFSkuUqBVGUCyF6Tyvl0BQmyGsN2bTVGtEL+7gOmpUIy7mXCjX71b2RNy
JIm+8pHnEDVR7Z1mnBJH+5bpJk/03X++cl8nGUH9XATpg8Kz3AS+PuaREv4HmUnP
d/0n7qZAAjEHDgEbV2X08f9keZLq/oPG0ZgPYtrijtmQq4qGFA+OMbBZxnAWvO4A
CN7ka4Ew6lssC0JnvYMPVRoIisj44YgPxzH1r9W0QfVVP6nIeZ6sv7oNO+d+WQgj
XCwIC1RipqFEEk9iNWaauLF3PRVLnNyFzySQ86IKsoWoWUgm9qLIuRb/8ysHhzaT
LJ4uyl8E+8MXJaR3m4t94JPWE694fAYxat7gI4kkI2VH3JJX8sEJjxwE6MKPG1YN
EfHO5FOxOdrprrY8mi/iXCfCR2G+6+B2IGyp8g+L/tGfWO++/5uBKqS9ejTF2waP
RgVmlcQX/7Hagxh04ZRaDxV1Moo9vH4VwRoosDuH531cIcqkr4XtkWCrF3UQFVlw
JJgmqu5eYwJWBqqTBfMoMDM2JJ5BXsNqAayKjcJ6i9QoCYt3Hlan/dlZYKOo270n
kgEHye6tTAgRJH60bzbDhY+gvC23x14EsldOALbqNSVgObva/7zAv/OTiNPjqGWO
h7wIX8E+UNieGvwwDl1D5kqHofjngVQwbS9wWdfmhBBObgxUGR4+4bCv0uj5J+KX
bBNfZ+vIio9ssYXnIFc+HpA44Y8ABpeqss2KtXzXCeRv2sFysrwbSSl7UbD9Wcdw
cCWbP7yqn0flCq9RBP8VcHRHtOjE6jNb837QEOcNQYsXH/naiQ/7QTZwIRily+Hi
o7KgatlMbbJ1m+n/J/JmnJPO/lB9XABKX9Lqhb8snhsubJSEIvpQ7f8qdBpaImO4
NXN8kHb2rbvIk8XPfzDEOHHcNobGK6jFd2yy4YMqQRdYMpU00XkzTuDRSFbBLm2s
EKmqVjFClaP4zxD8RCU7x1N5jMKtSFcUUMjptrg3FiMNZqk4zK7Qw+Wa1NnqaLOu
WnmY5bGTL4jNQ06uHjMELDu61XbwEZ74BnfkCrpte3PgCHxnBznjDpif+ibzZ0y+
DmqTgaxgBcmokBP1pZW36luAQOfeT0ANgd7nOe+ndGFXoXOMuDDpkinxHoAgTd/L
gC/Ek+2ywqJjJrUmSIyPstzcW9Df4prRK/3UlaJ922ySmRCPvQwKxdPzmsfvdu7G
jTIUc1egvIiOPuVLp18+QHU2A9HoYpwOP/iY7OJVGFwXFFsjp5M4uAVhqnmegm4S
r6VbUpzAhoAxNBia/aQeNGk5QaPVLtX2QOy6gnca7+Xtnn7haP+mn5KO2obsWmpk
F/tifsYc/sSbfea0GIJUvClIljdu9soM4DNQKu+9koC9rcgnw2JVrotqRZOc6MxO
TjC6yLEgY8DZyQfZMJMVLFyHAvb34BYALzccSIfsvKA0MPWsKBZgyCj+qSkv9Ica
gcbUBbthHd0ZDTtxGPw5kgPPBd2LMZHQIlrRqmzqNluJ8WWxUwV+VcxfCIi7p9xt
3zCFTJuNPwcghFTRuzmp7IYBAbyDZzRw2nxeOFfvUwVnmuweGw1dQVpXkdWiKb4B
dbyojCGS19QMWpQvB71GlO3HQw9mW0jY3sF1Lm4B8iVJNE7KtTScUBo/q+420QRg
ckRKPzHck5hzxBDLtKYrR7LHFqGcfdH+5Rnt7tFk8xM6M0omilWNMRYK1swk3CAZ
pjh7oeqBEzoo0wLQFD+uaHmBkaQ/e5Rul72HdhslQNNpVXkO8w0DFis0397rYuM9
diq1yfaN6//M1ePnYl1wrsQWHgauNLIj+joEbH/B0nAEjL736NOH3blX1qb++ZcM
ngYJmfJeIAV5vUYoghUX03Lk/5W3//S0oI0hFIRoSyRkmGP5QAEccz9pvEcS7wmh
/DbCGniPGwKTLRU2t+W9js8UIhvltgXbwxdUrHwMF1qe5w3ABlBNZ3jSJHduzkba
NNeSsmYkc+4URRoKxjvDmcA0joclqcmc58+W+akHeKwihOfM86NPoxmfBChIAQBk
i+wNvWuFbgfZ7NqsEZEpzPjxER1U4gBMZYsPl0gkHaKS/MJybAGLLmjwdmaLoETZ
59/Yqir0SyAKWxJfE5r5UaTVutgAE9OvfF1c9n98ou1EF6nI7OqRFNmJYC57YTE6
1Kws0cf4TqY7+x1ePXVdSlMPDJ2gyHo37YaGQFlBprJNWslwVjO3OjcRhv4KwfYZ
k6yu1Soio/QI0x9RwR7Z1bQyAxBJcN49zIRFWRXHT4GVHF95ZrRNh6Nwil3GvN3m
rViwZT44eNWafo6CL9VYMqXZxpEzm8pgRYkeXY/bhuyA7LfZoras92z/Gc9t59qP
iKiSlIUr+Xr/Cbo2tTUrnNk9Ns+jqLvthqWoNcItmrZogkLko4+yjo2Fzix+fB5b
KrW/GFW30Avj5l1/W2a8soJOYrS/j+3GWXs9PEeysZFrlQpUh0qM8ZTM0co9XICo
XDy59/rLLuh6cnE9iL8+pRmrc5NSZCdVLNW63LnQlMJwui6fSw2pMAAKMzdKCqTP
+iMEg3H23xMJpdBza7UW4q1JIes6pB+ZzcywC85LRLcPWmXl5J/yDazgIWKgn1/b
hu7NxJf9/YhvYz6r8pdrcua4bk40inhieecAHROnrYg29wYKq9RnxnHeCCuM+PZH
+ymjzPU8txDvqjoZwCsC54MYu3fXK/DAq1skhyo54NLGWj1XzFSbQmwA2sFQAVL8
O+8x0Fj1Ur8bcZWuABFUdUtLGk1pdZoBTdC1C4mBt3YCTdfHtHANyAILKi37byTO
vDwFvlcGr7yLfXaqvqdZR1mjiUKHS2us8n6qBE7WYxq3uQ8HD8E17yvXTfhgSp3/
u3zEgl4Vjo1dc2EHTklSHz3hNVKNQwgYBD+x6Ws33bgPduZUQsqO9X2/TWhnWjRZ
I0YpvhYcFDxecRuuG8IcE0IDjvgYi/DomDslgqKU1P0JYPAsZsmoXm00TBTxVeX8
XKBo2nsvHltm1AMjFBVc7d06+2+cmOjcThM8jpzp5KJ/QKPiNc3Ry4aPOS1mFYI2
y8b6U+LBTPUpHVkhLSlMBPHJThr59ys8M+PWp7u/yYS/nQiYijciHiFiT2msx/g7
N8ZIle4gFCUW8nSiTRDbp/DVdHVAeeVAON26y4HOnB3ossj41D8ghW4xfB2XLuL4
EW5paCELGJYG0fpfgkkOqMn3tFlKHwkoUUcxei0Fg5NTnI7vgdFf3+ff6pLnAHE0
I2rC9RNBvFePLetck9XFmrd5JyMqugzQnpA2QiYlH64WgTMP6hw48MJjD7RwrfCx
4TFY0fONk3yoyYX/TDzgnS9r2vRyFgT3fD8D19eJF2ldn1YQ6V+O9mko1Ow7nAH/
TbkiI9+q9u0b95UufdJFnSIqcABaN95LTVRKWAGGUL5gfG4P/7rmqKA6ysTbgDJE
yRfJMNIAeW0ghskKaGCXpC9IaH6mmMg2YyKxHcMmTgTLxy15ax7KHBuRY4GLJaRo
3QShaIKySYJgRBWXCNclWm7fRr8Cf/iXclcawC7hRaOJ6UqU4V7pIpEs0GGsj0Lr
bRH6N7uLo94M4NzYyPJ+rE/3bcOl/dQWIR1anlVTuHSvF4AFthrNCHTfzTK4UupK
WRaQF+VCByDBOy542xjziQdnBpLC+eCCFS5CLSHUBV4XzUyRSwIh2DFjs0NxyhtX
XXIWKNnIzsGJpPpGP8iUFv1FTUluKT4k/wW9dnZMSPS24K/QUdlntbEwQ+bGbnvc
6DVj+CY/Yy4YVTK9B5DZR/Qyfmms2OGvEJ8m/A58g9V4u8yXXI9qUpb+StvgiWc8
AUpTfiVcCrLQ/JCn0a38M8zOH+1MtKXR/z5vOQa8V8Z+w5/WxHNylUf3GomXfA4F
qEgV1ilbxd0WVyHOscweaCcPkjpNQ6X6q5qWCeNno2PEcuzuTEfVOn+fD8E/YHPl
aEOaLPRuxHVPmoco+Ku99n1R9fV5WCE3Kph+v4JjS9dZv34Dvp7ne25H3olDvS7R
06rDIulfSHUCJl0cluh8BZXyJjZctqddf1ap6euyWG3O02jAStAcxZNHKdsFNUEO
gHl2ASlDQlJ7dGdbs8rJc13ojopWKVAknPVr6erQ8S7P14NVeMMJeRnIEYtEcNHw
KsY/CrUWWIvC+7GHUZiOMAqSB/9P3jzbvbnrJbcp9t+bxbPyq9KHE0HgrffPLJnK
CxKhOEh7BeGUprSczI5EUsxerYRYxsXUooOk+Vz88djaeNj4nICvyEn6sCTEqv4O
7Ylckzcd/lZzaJjcHgntfoiwm2VS73DC43HEnusSdglpAa0apbYIEM7piMJfIcos
p727bNes/ixrtNaAoSW1kiSo1bpG+/08vIR99KsOVHXOllaItdiBcTQ+bogO+/WV
hKg8IeIPhPkefrb3qNWn7Q5eMKfCTc7X++6gpGF6Kq5pt8PzvWsU8kFc03f7IbbC
eA+H6eN/yPhHBVR5vEAD4xPgLj70eVtbmXeofXGv5eIuu/AESTtIn2Rig3UPZ0q3
Fdm3NX2ACEnTOSYDoyGsiHh1hqYNDm7evRPcXJBFUf5stbpWbH1p02V8QKWCD+Uw
/sCIWW8RJt/36qZUaV58aSKBBfO8TZFsiKMfWXhSlCy6WFJV9+Juj9RHY0b+aLfi
6rSqNJ8wX5/Wy54U6HLmjJJSalgeMqbxQUK+8y9wc+3CHpFIeebTG/uYIS7XFElY
V0HRiisBvqMHhxwBnKhhQ7l57UjvVDAn3EwKGIMcI4aMQt87/HVavYJQ0iWcxSno
ioiBZxpEfTXCSLgIojf82GIUW2J/uUH41EAWr0FqAxcPu7vB5fcTNQpnpyhrJT7X
7QZ4kD1FyJGE+6LPDAyM0sGqUfwevcNoVA25JP0kPGgnXasyxx+yct+9roz6ZG/H
OVrH17Q+GfqG3yU99ZLp5Q2uLQlvbuAzrpU2/+4WsMwYmnYZT1uuOC+OkhlFe2v8
WoZwLJqS3s2u8ojzA/9t/IqyN7GmtNA7b+xJXaImZcHq+zAd6m9KUViqEjkJhLjV
z74wnXEK/JAxsSj1SV7C4nOzK4DziT2W2z+PJZ7zLN3R92TcNR2RdjazuyDZy+kV
5SxTOOwN2o20t3LDVlGglemIws4RPqt/gfkCcAp8y/O/jzQZTtL2rkvFWAgtKEWJ
ZlBvsRfT+YNCB8p4RLkVQa23bMsN37wkRZI2fARZx0O1heDl5ds+qVvD3ulEL0XM
Vj9ou6DO5EwhDWJ0vwk88FeIoVsF/qNuX5ndrYGMBqNu+AxiARMn4PiqlezNowlr
K2zB3KwDqDM63e4dw0XJvLWBBBJrAYn0nI1VpLv31bC8zPKcSumo+DYXxSlb/Jvw
zlHurBzJAHBPJ6TIR/773aNT2JYKvH+NtaViW0MRhLAaxiBdX1b/JmaQlolyCEtA
O7gF3/WhhUSf9XOGbhl0PfSCbsTCvbDoUaP/FS/RyIDwF8b1ChVwnJ6ZNXR5Khxa
nC6aBSQJ6YPCDx0KQP7y8y1v+Quqh8e58WiXQzCFPkt/j0WueCXzO8K1SgaYMvSg
1iK9BQmru06hJzM1rp+KA73MpPKwV1zZy7elITwmCrQEemnD7JODoqwii4gVCxZ+
QTn8pP779HpxzupmTTpQxQghvb09KaoKYM51z30XHr6uGZo5tOrWKt1pvohfpNcm
7kQO1oi6Is9MAUZhMdM2RBXFn9mrG1IQ0X+qVWMrZl1KwjOX96FrXWu3ZTT9Oak8
nGalDPE47aWVJC2EEpMK7eGhjbrx8CaJKZ+v9jzhfgpyi4LWknH2XLtegKoZzvwF
PAP6sRR9brqg0aomFcixaeeb3FU+LuquSvE3gxmiyabkPcQVqhWx5CscgZjsY57O
XVz/1K+h0WkZ6Ivo3ClUX89t4JM9Of2qDvYRhv8ZaPt5cdPhhvJwY5C60gSYYuTG
JG6AK6ctBw6/bnD1MwAhJ+0nS7aTh752CNZxzlE6HFJTwbIuG9ISbmLGxnRM76L8
ueG0iyMbaJg0dzk6Gv4UzEdWvO0tCA9rRIesH1fboL5J3QM50koGg6bk4O9FYsJv
gWOZm1W8p8bAUfnxK1ISk22YF0iH+EQv4ctjptI4TBGlBo9qHzZOqCEd5ujjARvF
C3bI8jcFrOYb7jgvTQ1jq1Tg8hyvnUY8/wrKVPL3kLGB8T6rlKB+3930gz2fvnmL
uTgNHpaVvJUKWSfNONFObkFefCy/KUST4e+vN8H+Vc13M1WlYuMBycFqOt6GnKP+
2o2ChFIJNHVsAkl0eR0nBn8NTLPjFylgJR28pOQkxfHWbK7cfp2RX84vAuE8YWR5
RyWxbagmosP9rKkKFK3qveBsa+8yIVZDSlYcTjtQvG6aG3cdBYR+BHDSinq1+ved
Y/Kfo5+6vnDPjQL3C7++YpqFF2iIgDJaon2hj+BvykgszWYIr8NsykjmrGiRWa/m
yzVZY4uZiCtdGiVXg+nbTSjHyR27F0ulIXumc6RUXmUchQ/lBI1z0OldUj5E70Ct
lhN5BxEK10GiEWFSua0cXg3das1VZFYhX6HwctUZSkPG67kGWwI1+KG09XMfk0HD
oo9ia/fGNLjYxGkPdilYjroYRurhiy2Dbp6DwFZaGNlp++ntGXkdqsgFOzO+xDwQ
7vB/EgOjEIKY2Ti8ptNj2RY7xQqMBiS1V+nWRzND1KE1sUYGXjNwpJmZvXwUQf6Z
o0gEgQhNLLVJGTwveZG7UKHKjhYXPiAqD0luFHFJqzCRxSY6VrlmgqVzP9bvwMJh
TlWndcp1gQ1jcixzCKDY8Xpq68a/BFsDxLrLoSbUp+jqJ1C4GG6ldmKOPYx1E9k8
ROlB+U+UeEXgioObIjDP/yGn6Rwgriw7y5uprwhOwFKKjBX+P8+MbZHnYtVuhEtE
0rAf8AN9Bxt7DU2ftTjcAHUogJzZWRKzM7SH3vhLW/RnQr5YtfLKEs3peabe4oQZ
Vjr3ox/fXaN26OAN/Mqjq+jE/vnOSCgvpMyJSyGNkiLMmpN+tMtCC6eKVoUHkw7w
Gvk1++f3wggMNvQe9kEVCKsQUkv3Ef4jTtTDWmZeWSEWQiRbyB8QDbGy86cecK8e
q6z6dzHMWa0Il26gU2jZzFrLt4nxyr3bk119JHW/qVUAGS7y326/f90Vugqf//Fi
MUHab5HlLH4T/0C0XMGMazOPlW4P81evyJABkL7KtJx+RJP9r4JJmIA2itErJtEe
UmZ3VHtwtB1P9ao2DRLxznb7Hhnkl2eUtyfKiJiVzd4xXT5uiyZQ+xX6C4PUANVp
nHwE2SadzLPbjKYD0TVTA9DGmY3wy+1Pa86d6oxisXGLUs0IYqlM+iY9zJqmaJRN
aOR0rIhZqfA5xkRkzL9eJcg9QSWLkdBUE9CzCLO5xNhD/Eu3fow1u+H0sNJmJKGA
DUFzQ0jnYCBd9jk6XMO0AGMddpdckwgmYuWo+7I2MlhiJyaVb4wGkoSut3wl/4AD
KkKTOImOkOkm27mtUbMm0wSaWU5CdxSRNMBVA9LKfvyZJn0ZqatMhsZItdzHzebm
9oSon399cLiH0y9N1Lvh95jn2LBdQHtGdNmIGfVcKFNzAvWoJqNFLoOm1AGSzXrY
PzPRzFko7xDCZ3KByKiznPD+QoOOxM6LH96Ax0yDISfoNASFTlobxCLVwfZJO/7s
bBJF6j2zAOssw78RR0XHurBTTpA/fVUzHAvigX/q48DIPYC9gzB9fwbhW7hyk7EN
YLYNcYjjrYTsQcwdNVSFn6XysLaX7rHEFg1IVuPxKP+hOowdDjlZ2OwXwBMStG+F
Tb9+z2tQiTLYL/FUwjqBQ0NuKRoAYU/qJvnBgOYtP+AH5Ab3kLXn+tK7OtCtypCW
mu5vFX9E6DGIF6HauaYcZw2gRo5IdtR/mEwqhYFP8WNQkrfQNn0nSeZWlDaM95w6
SmLsR7BdaejcDEr2diEwuPk0OY/ytDAGoKQDjSo5CAOVCzmE2aC5BU/2h3mX4xfx
UvPSl1+QkeppJk6tKkKJI9YsQ/96JxwianCwSs0ysXHjdHH/hApQxrEOPRcR9zwH
gMaRrxIR+hnSPkd+ES/7Q6iSt7p4yZf02utlWOvVNEq8UGwbBWDtuN6sBaIclqIe
HCox6JGD3IxJohiJTraicmnDKGjGPLTzxmEKhH33YOQ7KdCqewD+46eY1hl/GXDT
XIoBSlRFfkeYY9m04cT0hBQ9tUJWwmVfA/7KbjPjfR490o6pxNQRCJAILyaNKOgW
/g/s+ShddX3o0SINQb3FNYeoTK3UIPvEk67a9o+24EXCFjUW0ejvZDN0OxvPh3rt
U4sCCstqPeAH/wkfq0oDtLX8XjZo9c/xzqIOOjWZXZwSueEBPNJfhgQ6mSzJYx85
TusalkB19A2jPbxZ9jfaQvytgOQ+caRA083i0rnasrlYC7RTKLMELhdhkVWbtZ23
ygIus0VPvDKJrX9NgMCssKaGm3mHidYLg6pdioLiTdT6vYjIzuBML3SWCMegFFc2
qevWFO0TFIrGFzF8SPp4XZ7JKeAFjvXJZTXJoTCj8feVrW32oLlifPLlTJWy0y6O
vql7wN34rOS05OCTWbxPYOJ1g2xnOv1vnkpoTO4nYcQ4bJbHJyCV8TtcC7nE7Ru6
jqGwMQXtRelmtCNEI3FQFNtxmjg+4kraiBFg05GEYdWyVux84EDc7ESsSU1L14HG
oMi3ajHR0qc1VfYFgCSmtM+HKD/OH8PvTWZsa+GDMlNzGtHyww5d9WT+jC4xxPnk
2aXLHYDh0mpYKJrXIhr7MTMzeIatR4kHh9eQAisJ54X7rsjDKs+9IlQWDSeXOAS3
wBH/4jlrbd8c66JFwi1u1MdRU1AY6RtBXHWIQuhNDEb32KVHGG3o8qbBSXHwm+8w
Nrej5z84Ht7oyD0b8/SNdI64S24Ya3VOY8kasdj3qCDzbMIm9rkhtl+cDIh9SNLB
hhi6LwVck1Kb++/2fO6esNlP+LQ7sML/fyzAxnJgBtLPWggb+I9FGC6NsY4D7gBX
UAzEAN2Ev5ss8HBrbvnii3UP5qaqr/oZWAcxPGi5lsKMuRnBiw0uQTo5PA/uGZlG
PN3hDaQi1P1NVxTlwLm/cPyNqJlyvBhRXLTEUKIXxx6xza5RpEngQLGRkxIiMSbi
JLHqxx3FWubX5cwjszaQWnUZD0EWyQT+e8iOKWV6dxsblhxeJt2aZ1H7PtglLP2f
GpUG5DvbSsewMSDgGLqtviJjj+4QTD6SCEe4MKvDpDcXAzEe5ZsjtUdvujm0eGvQ
ymbx6/Azt4Fe3i7K/K2VBCg2ov4Csc2q8oc1ge51p5jHdzlPdoBHARhcePQMFpkN
AQWhrwxHvxwm/t/L4L6PvXyOP6Ao2Dvnbp1rE7p/pZy16vFiE81xQGYlRBG3aFJd
HPi/OHI2r5MlaJigBOU6gagmnKYR1BMWw5g4sNPla4fHz3cFO2FXeeIpuZEPAg2M
W1RWeLi14uZtjWu2yo2gh0FDXTeviIMf5+3KdxChw8YAOGmP+5xUZmPC6ziEYRv2
Uvi39CZedrSywWy1WRNLAKnRM24/yW+CtPQRrIKqjcMrydkVMi6prNyjC1rZDRz6
0YUrn+vH9uqEHGryy4zJKSSD6ZAa9kFlnvlYmPKHgZB+3gGUMMJkojSz3EIc72Zc
g1bdY8AH1q2/JiwG8FlEo6twvk6I3+13kXC1KoXTp/yhVA1zRtYBhnz2YxL/enlX
y3xXNqZZtDlT5sNOglm0coBUG0wq1z4ZQn845H8POLsp93/4dFLHMs780XrjFY35
1k86NWbsynpivCRHsGZb+WwlyM6SYzqWvONQmUnmzB+g6DMSZoQ1Y2U717YvvwvO
eyzB9XbhXbATRIyWq/NAqeiFIFhewngnA8VYqGto3LbVXHZULyLjBbRaB7RZP5+C
XgD0n1nwzfFVCcH43Xc+Ct/Nwz0rjVmn4x8ZezMz5beFh57bRT495DWPSLGTmQXL
GaI9HeFxMNnDZqb8ENMBmJB28X/0rf7W72pf/NPoicseZ9YVxVbXTrTCPwglgjNF
nnC55llIdRNaEnuKcBFTrCDFgdglA/SVfeGU49cU89ic/dCHRkjNBIueTjaeik3Q
NiXWcycTn4qgoQ9j89+xMBIwJXyaPEd+oIOe5gJkvIse1w1iHJUuWd0Rh6Yk5xuW
ei9MBtcD2GhCjfiu+X+aVuPhUvKd4HZpZAkrvZsFqSw4ifvHHpbqFVVkp9F6iu5b
9lHV9/+Q8LlMdD+d6T5LkbbwCp8SjXPhOjrNVEQJzeoB93k8DYEvK6owZu0aan7t
dZN98A3HHtIhDmqWTXj6Q5wHO3FbTlZ4b2zAJOFRS1H1UQ9ykF5Wodn8LC5uE3Hx
FDfZx+H2+62k89/6YdnDtpqmEcNd4QQttlNLBWf3n1FsmrB5aJQS9feUltxnvySz
NQ6GY4KDHPihGqSp43O0J+pRmkpOo5SyqHmWyulyk9sPZyCMJbdWB9cO1EkN6X86
u6nbf/RQFn9dPUJ7ZBKjA1SK36lwjAcR8qUwsR2cSG3W8KWJRQpuqVVL+oNhkQhc
Opvo7aAd46hKBK8KjLpF4pjWaTSz9v/B8RMkKA0NffEH9AGT4w6E1Vcg6ms2CSNu
fQqxtHTGfgnUad9C8C7tiWcmSWKgIY55DpI4XTWXfFZM2T96+hQP8ww+rk6NxSW6
pesoM79AxuUoyAwQGd9n6bEEIVYAY3BIYT7h55LjaKvq6FNcQHHgM9t8ZgRNOUAT
iWIR4dTVudrx+O8OkIzOq8s0qb0H8IhJHNAMg8ZgNPtdXvqndzbRN12qNCPeBVcL
NZgmPIdGN2AhK1seiqMfKlUUj8n7VKaCPDShYELHlbz8QNknhu5WJvTHFahhvu1g
3Um/bQUS/JaLTKYuz4dxHtF4BOZopU6B3wkOB0qDGHyEhCE4XrxzCOnAGJ1OQ1ZE
z0IinPCxh6uEUsk9Jx4D8U5o7U+jMhQX03pdJq3E/nJChqqrsqb0TE3kDtidSDKV
Ea16AJc26n28U+Mf/5aRJxvL9QUdtEMUtMHfCtxMBXg0eLqD4PDXCFCuxgVPi0Kh
pKwwexBbBecYlQvyc9+jxtOL3Q9H7byOVSm9NvYd+ktT++lbjj0mcNgmwxu/1GyH
2yNFaMrjXAThYKX3n0FySIG6D8QxiHFKsM2ncfVXojgCHqDkbEjqPpx1jBs5easD
YoK3G6y3cgbrVMvd6fy+yBfNoYYwsyMpu4I9PFt4hKSkzDxqHLXBc1uKY81O97sl
wWUvlviJJA78kkawGMeI8pyqWXlUUtLM4kr1gRFkW+H27CTAQ9U+Ghk4flQcjj5V
gSS24TueeD1kz4Hk97OevlEPGIRB788pZNy8a6p2qPFUsHuJhlKLI0N10IddmDoQ
/9KCYHBk1OnQZxD+jTckxQHoKOrfBNKraLtKCUeQ1cs2otCPNJKCE1DY2bxXSSmL
8BDLMLB/QUdysIWhEB6kyGVXaJb/tMNGfELOo8G0douhu0YysCaqFGcTQnvPLtif
vjVoUXdjNa7eROWR64qQkT5rsHFbEWxiYJMcEwInrNL0H4y5eoIG5/LAc4t1bKtV
7N3GLiB56JIRHw1Ke9h/Otm/z8/AI7W70NFETaPyX1O03mrFZeT5xU75do8eB+kX
YzNOc7B4P0G4p4bPuK2GEDvDM+758N2l35tAE1ErD+LeHAOlGWuUVBGIIJbbb7Vu
uqxgyZwPjKGP/HneMuCuco71UVXDhZp+XV7VoPLwESbjyi6lFxoa51Ns9atJ5z6C
cDzUr1oKS8ouhLzvLG+uPoMRfHOi+tj4WXgECJi2MivON+KuH+XxGw+1BR1NEbrd
5OTw59+a4s1bx59jL/ICS+aRFuxPoil2w5GLAK6AG3dFUEIWi42WL8vRHegbR3qw
V46RICYiwiuMQ9vQtqNP4adFhspRA5tcCzZozXpxuzXu7KOnjsNPz0NSfcOssFWl
MWY64/Jf5IFK4CKvaofbWYUekOvrhwcgsimukklxt0kcVqgdyE+ISkLNNcoxlVRJ
rive3cAc2Sk7xYN/66tT/tyHmCUJCGZ3XIUMZ/Jm83BVlqp7CkpDUgMFDX8VtnoL
bFQBBR6FROk3yeAmSlwsE+eeMQK06RuEStO6J9Qh9YFB93q0z5LwcO+LBXVjrvaT
JRv3DQjtz37DUmlssypEJlqxf6gkyTiiCOKdwIbNQqRhdsCXElfcqee3gARI1uU2
BlKP6KPKvRt1Prb2eIRSF6tlicI6GM5efYSsdSsYvP3AMPzfO1WZJPpke14D2pz9
sdFbCtNuWQHmX8XlOREeq95v0y8sghyW+cjEFgdfaTuG0B4YdT4wB2sVO4cwxYda
yrrBfP09Dxho6SRIaVP8Y1f7jWiDjkRlpcVhk4rpQ6PIEKQ7CQDXUwpX9w4ARs0/
eS82cR7jc+2rBkGBB+HTdJ1xAbttp3HLMKXlhBaUPuIAn082/fH0QPlFkoI6unvs
LAEfqFIGLymUZin0ImS03+sEDCnHijqnNyKWk4TQ2uLE+y6XFmoPpWjJ2VBY9ijw
QdT40yVnewv0B2JWS8EsY8hB4XVr7j2yZdexCsm1tWTOdbZQQi0nO/v8xCVfm75h
UcvVK3CFoxNdO6F/QQl9eMVgO66Gl8XGqWP62lMzx9rwXvpvex2t+fDf23kxlRNi
jbLqthFdUOHfQSvb/ZkI0ZtPKOvky7mDIlYfzMXWjAACYzAe82iQ67vL8hI+WeJw
qVhK98VHSm7o1XlZzewJcT4zOU/rAUa+djQ/cYt3otSe4ugQhm6haN0PpfCyVGED
qx5+v2xlhgH3Ig/mBdSfw/CIFv9gZlrGJ4wNcO2Mw9bVNfd54/Oip4sGil0Kf/FZ
1OY0+ws8u9DxP3n8ZFhio23qRCjOXbOLzk984+sXZ2IMyLFVM426OFdX12PnyBnV
vJVgo9xWxYxDTIJelrqHtIB6wtC6agD9alY6vcwbE1/jI4gtXeyg9yDJ3STiQHOT
mCq4tRhN3w+4WdCBysnfAF8n0/q+QDkRXtsVEFEe+RCMQv9uKpW7j6bPCro4+yKm
dcee74Amf/5b8dtNJEQkxkIj6f+jTGjp9uxfvkmUXMITSjVSiLubXibUo32ZdWYW
evA1mqAnLSQF9L3UopKi+UYiXCNEF5UHz4L1YFM8sh2usd9esmiUxS7H4/k8QFU4
x3uzk3J22WLww8o08mUnYfHZHOiB43aKaEAmXBmZl1b5hJSljAWTME/Xb+j95+ri
t49to3qo+dA4/6G8JlV9KLz9muLhxmSx37+vsHe93MPRi1S1Qgu9BMrv616Zg2V7
/6JrmWDtg+guSe4+hqCdqx0WKDQJST6eiuMCwjzIg3FRNQaD54KDK/Wbj1NN3nrj
EHYJxoTGHUqrr3VeicP2o4UGPhqYQF4JGqFEzrBZJ0EFilwvpnoEeoaGHug9UlnD
ZwxsKggqUI37KrGrGr9q4osoh3WeQscZiR2YJ4rIMH7psp6rgzQEwvIgLNYD75nF
NgRxuD9JiEJYqzcFzGFVAQsWQuuoKUr34NPmKsV1i95izBiXN5jpzvatyktuS4rb
QCeJ9Swu4GSZiwp/a9IPZ5jUvlzijfj62X1q0tplo/51S+chLpuwOM1XVoR/BljP
Fn6QMl2lorITsR2o2d3Qa+cyT+64pXju2zDuHjWVYB9mytDsVl1V6xHmP6yffqXJ
eRNkisP6QJSd+1y+NqDJ5cS0q0v1INTE7gxyDo5WbI8c8hGEuktZjA3AchDi76VB
GIh8znmk7BEK7q/8ybSEVB0ElXpyiqpDgWhjof3d7F98SL9qcLK/1j3ODk8k/acI
f+fC/ZpGKY+zQLI6sBojWaQE/hWqjM6joOn5ZG3KUcTz9HxmWIGatzXIGPRhzfH9
l6N9mKrqnY/kBnnbf3+OdawuoR69njkTNn0n8r221yhIjWhcl8VIM6vnPcPVkGOG
1SrJigICOkBOGA8eVxM5LdA1DwnkZn91XVujQn1IXxiz9EVJl9OwVgtbsJapvodF
9Sf9Y523y05yCvFpvfNS3VAkOqYoJCVewbPG4CZF0puo4is3jQlKdHWfiVr2vX55
C3zEpXvG01iJqeyuWazc2AyBB3Ge6dK2WrAtr0p82VmMd6kGf01ISoTn9UYmeSyk
72rh1ytCNtYqaDFqoc3iW8kQab2+mWhlDHh5Qoghp/p17BqePAs9TIlVF2ovfEzu
c3mU3l0WHIgQbbaeIAARBEwGAFMVj5tUllWv/JbXy8dLpz2wb4rUq8892OghfXuk
ZCbE9mLNUuM+RxMsbxONx52Ni0wbjP6conIZQ4itd2sXp3Rv9RbloscjpdWCGZdH
qpbYIo+TFX1s6tUqrLMuXGnQUWYV8Xs1QD4aFpAehUr9Kgmj/4h5WPaRoKzBD5r2
s5lEvmivjonibO0TjT3hIyuVygGvNu2XibnC/aXrpIZiSwWfHLITRSlT3ozl0FXC
Q65CFBc+2JG4Pr7eCw/VuC+Oqd/GBkNWoIf6pGq7k9hGotSEHie1sjCqJv3inJcs
GyLxkgJEPWeEEP9Cve06P7tQls3ftHavMVBo3KNTe4lwQu9zekp+gEXn4FlnXyTW
aO5Zh0ObheU4uvh6chUYAgvVBrOnEeb9sWPSzJHap+kf7bnaNBaQLnH7PcwMF8n7
Gsf3Nio9blOp9USbtKXtSx8FOVqRVmkm0FX3V/hoVaybaLs3jTmhkOYlANUaW+B8
/PPXbWdY/Vp4BEmodYlYr17pu72qOizqLc/RLjxQYDPatiE2OWO3C8sTnyLr9u0D
B7wvmSSxFa4jg7tjJmg710Jrqnz7OHG6hBQ6ceUp2wSiskdAyyVtIVVOlCXHzPvc
SPaKicNn2ze8YbN2NJEOIGsdMvlJ/gZwzQrshfD6EippX6QOjlWt3Q9oZuAvX+Im
4ZcliNk+mcP83Hgd+dP8m1hBykzwfKcVYSxN8T9IJDT5sifzbkLYUlXpaUK3wbsP
BcX6dZnYXendFU5YNZyCptATJHukxMqYj+r852lBaAjxu2ZTC70h256IFomYjEhB
dglLsJ/yjVgMJTrWYBiXBhC2DeramwosMosH67fo9+bKS6Y1eZ/8pjBsv5jlgnCD
sAQcwlmh8vupNAiWC21a+KLFn2hTibDsJQVkARy1Mdz0Vq91bWOa1QXD45+M4y6/
QTYAca6/RzDboMKMDP0wlgYBrcXBOwuIEkE2dIiSpMMDar2rugWKyzz6XWIdtpn6
nlBhw5cdP8F2rb/71+51EhYhDpZbShOt4D01mwWQUXoPrtbgcIzInePRMEKbA+If
IamOSLnHDPArCrF8UgFBayI1oXYkSKXLFZ57q6/sqxuJB7V3QFZ9ONA+PUdhh5Ke
2fVYWebcejmNQcknuu+OhErHwcDDRSfxlgXyw5ArkxwQLHVRN8vi9K9fI6lCtSEa
SKs/HZkDWHDf7erDLQYqA6onELhxNNKrtz2/sUQuHbV2KyJPyXBxSbkxQdF0SClb
mN2YVuqzHVFw2TIVkQwho6yLejeBaKkk9EeT0NzkhJmtaalNN5rFsqXrAuVX52HV
OaeLAHa2cccU0la8G1az2rl4i/JlIPc5DdqpExzxyPcFzkSGWLT/im7qfLCPp5Px
paIfzypNlCaOWYNLPqYvmmXZcpJAvmcH7RjpNm0qHEM6n17mzOIQ4vFbpuXW5Ndu
6qdv+zlcNyMRX80COtl+1PIxwQe4XaVRvPGu9mNy/dOMdmjgVLiqPs3tbA3y7/Fh
YQsUavgBDdcDOB8rclCkLlFCwM6kq+TV6q6owE84DlAIRaeYVeD3HqwqQZyw342X
iCP8Brs7U6uOMSwzxjyMowzU4TDMkyB3tBdQ0MBJ2By7z6u0LY4RlC4kp33UChF1
Zy1oVgEX/38FUD6be1od4W0GagYftUDTHC1M8VNgae9skhzm2Sy4e+/AdQi3CBJ4
TBjuZiHv+daSs2JlVFc6yMmBqT84E3N4sNfRRSvtYGI13B6ovTkeU3xzwwxpa8e9
2N5D+b8jje7SUxuxq6n2sAwP1Er6GeEPfwZwtgUkR52JUJcwjcQ8e1aWQl9Qg2AY
qKvDOQyqspAcEdLyKhUpaOqic7mQBJZVBZ7XzzwpfKcsa8VfeESFBITVJnbIUI5o
fI/8C1TuzG3/YhBTpOThpmPHGTZbNhlVhUyNNGL6PHq6nU6qLlFu4ZxuAf0E63Pf
NtS4QtiERpvhdY6BrL+3ccEM7i3AoN3EAohP04UlQ9v1R/Ts2/x2ayfpkf1Rw7NF
4s/R2JNrJBvwgF4NIHXWWsjpyQP4r4O+XNZ1pckg1Liq0EgE4vgtW7TN/oc6zwD0
UuuwSqPXZcXC67UMB1vCqXE98LJ0jjvml5M1LDKF35mV/yh7Z0QLfQTO70PJ0+ix
ZfxPQsuZ5KiQdwNjNT7aQ8jjQSFK/8sHHA/Oe9R7bdHUHyvzQTBG8hBaJ+u2bG6S
fqBefNw4FlyQXWF91GoV8/qGuaXtlrrPPZr1CFqIGaYcQF9OHYAWGTtjvXXtaB+6
i2h9GD6MfNLMdajeUefCeSXhdYJuBPtl2REpJaGH4Vg0MjIDi9A/kMm6P0s+wQzd
lAsPPcMex77L3rWAgcwYukUNecGYCWiwqg8N3iWhPn2FMn7eVuOLnMsi4WL1KQIm
Is8RbhWlk5Cx7dSdPDAotnp9qrE7Bcs0BIuYg2y96BKp8eqhGr+oBM6XFEYe/JBu
5oFRGOK6ZJQzi3ZcktaU4Lh7pBEfi1X4VjMbExM5uB81i2fB3uHawe9UWJrlti/O
zCuxnZXteTXnHex238kOSoy0b43xXjC9qCIxGO2cNQN/oNrY/W8dVoCKSKmzKPgs
C7TNsvwH9KMkZwhExk7wAtszjJ6elvmt69fRnwmFlPyvyWJR8HonoedxB2sPGDCA
gzOrstOGx1hGJ1CjWWPoO1NGULZWb8SN5xyFye7obcH1YVGaj+KOVPIyMDvws23g
BwBMw5dH36b7Nbw9i16+fGecXYiTXTZgmELhhvctBvYqSZLxyikxbHa19WBvUhNY
vsWEiAIVdN+ZsyQdPoeQKqQopAHh4j1Su4Jkl4IiCHSZCV+WZkP2bamjoQC3XSMn
ZscbfGNuAwbiDlzgQqEq7bOO1kshYVdJ87cVWAYbeOl+KRpT1jn9ZB4SQPCIVGzh
/j2jK8FR3Olm8iOe0noj+s5XSdwp6C7cw0AD1RjH8OSNXEc+7OdesNEuh8oai8q3
waYrfvgufsnVE3MagJyfj+x0MHlCqu3ZLFtao6moX5Rg3KxT9LrKTGiOMngBQLU1
VXUQ6V+lr2hi0SZaBHHyNRVMxsFW/2dq2b1Phu0yvGJ7A0Fi33ooUHTLN5zMV2WI
ox1V/8I44XtKx0z2oiuqLRTzRk+qrR65FmraWnYlDt6eqkRIcQPTs73TYuruh4qU
PAx6AK4WAnXGCPN31HaUaHCSLIqVMB0ptNd1hSPpVfA8pkw8sKTBwGG0XayRSfkM
Bq5V1F3ftSgzrC52HI0vTzIghLHXnkk/SNVZ/v8wTRttTMFkth9xjU5ZDfYA+2zg
QQcDU83w0Be1rAm1l6tSWgx9S+DWWDtk2kXnjIk3tqpzJMze+ZDsUa8BL/m0SUqA
ujdZlgeN8N3QGquT1LHUD9p9NF1akpL+Aqbah9xzQu6e98cUszCVuAhJnYbxI6BU
EbVTBW36pR1iIQXS88TO3FCLkihRC5Wtgdo4Wj17e0mT1lWl9UQF3nZlh7MFAZ1a
bow93/xvmq5J7idr73DhobDAZ8qTjionr+61Oq8SZGLnmyiS06cnVPOI6CvHHQBF
u7nMq7UOpTwWlqRkKmzKvmGtx1SGxbCnsXCVLFtCZmR9OKV6v5KdIV8TwskY7UNh
kq0m/SX5s2dtY5pS1xQih6+/Q9gZC1u409E/YSvmZ5DsY+xEL1sW7S4BFGidzVdU
EkFIj3TV+ROxrYatrXN0byL6aPjXVVaKxBRrqeqZ1QiStfqj9qtVN1ju5/xwAmUr
2Qj0AouVapKww2+FDepsvUo5XI7vwaHkKp6IyKNcYLY29XNF6dHSmh2gFqXxqdVU
VYkUopOassgDYKwhP7p2t4TvwdyeDtq1DQnLL2/cDjaKFjq0MP977quAr/aYVhU7
m+3lS2+fyJj4eW5zZLUnUK3EFDM9wER/NwAcemYoPV9832Pjbz8Kzg5qgjGFofhu
IOdQFgqRlSweKqWt59f0wONzsgnERoqSU57h3BNl760idgFkR0YtQubdGnGIvcme
suk8TmdooOhUxN5oDwpXh11XLftUCkuRt9esWaRHT3KR6XcJxP+/SuKMXlnzPXIe
1nLLSPIhxHRM1pErUsAhAsoWoxNIaUccStoGY6m4jN6HnYc5jdHfu7MCpTn1lT5F
T30RyPdXet1HpmtD2EazouS705w//SfluDDNmGdNqpcn8Algw+hmoRdy99vTChh0
bjRl60Ycssj/n5ofkwcJa492qI3lEtFwJD9Au6CKbkkGy4NTlKjZBfMEMZ/C+NkD
plfkrs3IxTntYiER4xpk9dXDrnpoiel2L9tfRHhhr2+ZDI5S/K0mfQYk7F+0h6Bh
sz9WAlngDvq5xnvBoEl3QhCQhtwANRDs5hOnwZi9Bve65QPNGF0Uft+FyfbMTyF0
LGCfq85X1Q6DdGR7t0aYCHs5pRDGvRMwc0VN/dHDh2jErUTqRCH70RpNFZYLQcWq
ZwlGEfJCxjkpLiQXx1/4B8UFJZiX4IQDto5Yw9bnz0RC5JBhhqHqqUykUYhXHrkI
XF/AFxL1k50so2B4HqvvIGcJvp+tI9kpHCoSfgs0eMMbOa1bJQuOEJ0a02ekp9Uc
9obUAxHcSPTI9HlmbhHjW5qdtYaae3PN8oZ/B9Q69yI1NTzqTl6l7uqHuZlbVzGZ
Cd6iMFRAU5aYS7tWsu9b5DX/GGQVgv0+9QhzTnBFHl9PAhAO4Lhxsu37kucECht0
EKhyYL8bdOVs7PH5PI1q4B6lhb9R4Yjj80oSDAfhhU7u6zCVMfgiBbWqx2RGMCcy
Q4QkPaJMNcVkYMWLFkTDhiVflUMFgA2SDkIxFjUYTmHgW0ZOzeNooCPt0b0EVPG0
X0FVSaPO9vEvw4WL1Ox7IQ1vFL06u9QaaYfMTTgEad4IWQnjor8TYF8PEsmk1uIX
FcKl5AyJmUZLpwEazNhZVKN8TF9cpghdfDhGI6YcyE/oFd9gOLDmijTAvtsL12lf
RTDOnXZC0cVG9IFs1ai6zvqBp1PvAuartb9kpTeysCZfXMWBX3oOXV/7rOH9bao1
CpT57lgbk0GrbjnHXrCnb/pa0SU7MB7FOz7uANEVZb4Hc/ffmssTvmJjghpZoXj8
1IBJ8zasHeCpuupoXaPcM8QyisPXh4rCZf4qbZWNgQPddzNOHrI2vUR12FUchAPF
bU9i2UQ6pzAWNYbfHuqwsWDdMIrwvErQ9Y67NptpOqQAf/FZIEZRWmnYbpygLHMs
BGijl/LSFsjMNCnaftB4lU0LJNZ/pX/CA9BrwpJrFmBwMOwUh7ML9Hfm6rrvaS6v
Qrs4eJGIvI/v6R4RxqH+A4DZcA1iV48z5mqJGOcFOysTBslno24ec91qAj7RgqiO
4OwtAuQL41afmKjb2yKvH8d0pEllh6L3a/aBs7Iu52NRKhrQSGVA9DTC3PInADMW
S48lbAGZjCVaDgLWS+ugkg0UImS8OcjD+wIe3SsfG9ROSnok3W0bUMMpBgLK3Lu3
8fSbhj2XF2emo1RprvphavVc/bU7BFioOn56CKYw/aNuytSILTtbNZ5NdVCHM6Pw
Y1qHsBMmso1+OW+X+LBs+CfPU+GIVfZQCBzaAmc5x8FG2FfyBrL4MBziwi8D+9ek
KJsI24r3fh3eg2fQ1+kq7H2VqWLFm1hmxUG/P0lggJXdvXTIwgX5VV3gJ4XyzKJ7
Fblb31ALfCkYpytbJDty1nqgFF6UPR8ze/mUFKXgMmHKpdoUNOAKuyGyTD8DDvgH
F3h4A0Ur8U+n/fQLDLdMJ6AqTOPXZl/zENCT7EBh2wsqnmi9Un2smtZGWct+w9Ye
NNXe+qgdAb7NWp71FcowpJdTgpU7dUekltOj1yZoGhznG6E8GrwGcD9yfPVRMixm
RVlTt/SME+hkxybQGvf6/89R4N8oVWeihM2y+siFvD0sD1fs1rzx98EaLb39vGTQ
Ka/kS/zYLtHHXplug1od6qKRAy2aQue0RvRtbwJSksAOOTG8FBh1S5CyAffkbnu8
pHoHpjX76J2eK2eowsFh9DnHU8A+YALrcoDBlrlKB1tWySo7ODfb59fkOgp/F0mM
eKzG5Y2bZ4qg/ghg2cyvrvSdE+klJWgqKAF3Y44ycwzP2cbLTcL6by2P2Ct7oZ8u
mN80JJBbozshUusMyseNx47j1SSPj5TyvO0kkRgE/GfumSJZV0v0vbJmIgLIYlYp
T0SJJ4L93Xgr6k6DkfHN+GB30hiHa2pSFYaMJZhH/mg+Q0IhxsSflWJeYwCgoyJN
M/22fFKVlWdPVrXShcTSmHNNEOyxvGpfDE8Kwkqkpwm52/qhixaeoCapUrBfOZh1
6IMqifgC3CIPIjwWniu2gft3t0MN3xH4whkcUi7GBxEq3jLm6YsWZHXoq52lTKBs
ND2VVOCuvl6g5ZgtQpnfG1WPgWir0pUUtwRF9+p8ZzW7/DieztKeH6oTxETTjOAM
DY+X3buxZ1zsZEx67dKxhNIevYCUuezGY8uhhP+TVZBnRsM9Zqus5JNnEaq6S/0O
6lPuMHM6VFMj8AkghPJRAKRKCJM2eIr1HuNaRLZK3XepkL4RzujFt73bjJ1b9fom
/i2rSG59ar7Ii3k86/HkU1391MOQMVs7Dqw955AAwWYju2hIsWYv/zeyXnoYn6c5
BcDqJoXndRe1jMVZg8QsP17ezbecpgeGglryb1vWuTpLBt0fUdH4X6wPmH9jTkDH
dAKLeh9hyS4LKwdWu1PIc4nPcqJU01xBdhh3kJ/x2il0x5smHBGa/ACkP1wdBgcx
QRsShX1jzBjrl+P4tPEScdQex41heibp3d/6gpl/6kS1OiDQiRPye7SZLaB45NjG
CsJjBGs55pnj96/zHiyHza9zbfFI49AGsG7q/Dp4Qc+1NaqxOp8uxOhbi1g5Rmh7
IzAHh2LVk31XjH1pTCG20/CDTkzdF1WD9ayhsskW8Ed/4p3OuCWeSLABIujp4k39
PkRAyqEA6Dc72zNgg6m2CatV5FhuaQ2nGgdE+tU8Kjw9RIzNeNm5jn6dkY3YOXFB
ByB0B7/hSGwemrLPPYRNuVq86clHHufxzm9p8SpniC2rHn7uuMIUiT1FPM/jmYLU
LA+D85J67UY0+d8YDpVJeOhxqQuF2hJn/dtvT+hHOmZGHyycK0+iebsMBWPjNuux
pRZBrZ8c42YVVm1aNDa9h40jcrghXFRJQVOpkn31Q83inOYbYkxnUSoV4LVOrUc+
Qt8S5rpO2p7BuZwZJpiX6LieNe127IEE3QGH15H4kE3oTNEMpPuG7WskacDPLNPO
ulprWbNU2HwbZUCxyQ6TJ0LqDLIDzTOY2VQz6yaBW01piiTWRfOhzC+/AWxsBXUD
YDnvjzHnCQIAMb2Z6T5/jKWzM9Sf3mGN/m95BRbd+j8Drcs9MfG9mx+39HoVtTK7
h0gCWrrkeGXn16bwNHd74cfGxA9TpsIO4pfd0u0pxC8Ime/KTk3pG6mb/Ro3JbCf
0Zq/7rbVJYadJONs8C2RWLMrBVTsTNVONOmXByrbN6HD+BdDjj2jgJaIXDE7/qhx
L+4sjhvc2iRKORR4bJLwCmu9Al6N/w5ktug3WT2PnOCCLO2RKbzh9OgH/y8kGJuK
QCua1ppJIXubnxg2G0jRzXWWtDJLSq043lVeZqZBcR3Vw3tmF98Q2g3yUuSag4/u
5ZEaTa/uu7PyJccT3KeRLuHgZVKMKh3Zg+IfkxYDEWORMRN88G2QkinVgL/OI29B
hQcm9LjK+pFaisFeO6YS9L21XyUgE1zvNhHN30Ra4iB3Mr2cdNJoWDoiVZNyACen
KhRTGkvhjLgg0r+rp5lzBkoYimUXQA9tGk86/nu2D+IMjvds0EnCwfEv3jIi3pR8
Zuhr1S5XLCKSiNP7W31u4oHJyAVgAv99PpPIjeIq+VTTd+pi9jJEQuWrtUKF0+1g
JuJogevQ7P9kaMcC08mhUYHGuydXUcJk4eTbu3VBTzezvrvEh+f2yQG1QT1cC/lf
BKjFXCqcWnS/J6TJ4J2TK0erUUB49YlaPSK6aezg4ekD1Mh7CRwq6fPZT/R2L20z
kvyqbkBbuIXM7FZK7mUP6AfQALj0xUtc+SI8mLTTelJkCQg2ubdcKVcRkPZVTvPW
uRffKymUNTuyoKcaX6cfeWBWkTu6r98DWwXqZI/ICFE9cou/DvFfjNOve190hQzV
9N2MoEMjIHeS+i68KO+3CD7BBUsXxc7r6dRyhRM0fMlHvXrH6ySxdEpTPWI0Pxnp
7mnMF4tJMQ6sTRw8yLUjmh4/bxAotftG2f6nksO/U7Nae3i2cghvikeWRGap7Fyi
R8J3gvEfQnG+10q2drJTY/DF7sHUgw/RCvoDLd3Z+SWNdR+VyLfLq1pOkMr3a5IF
Lc4I0mhDoYJcOB+wNb6nuPQu0zQ/xGg9OnUsur6Et7oIAS79pRkTXLd+b/Omcx9/
J+M2hEu4dcq5BBHyFlDbfCjilt7kx4IpXxpLHObC437RZJQJLl0P8xGg6IeJpxI9
xiFz4tvz5BSG3ZGNFbDNStBfVCRtPFcEXQGKWWb9cOomn0Mu+Fja7bNKqAyGI7Fd
vQ9OPNUmGC87emCWP0FOYyf98fiH3oPL/YjEEIj8ryb0cJ44i24v6jDd87sQBZpI
GUol9/4C/9prnCqWnpWZhz8pIFN7saS+KuAFEuUZVDA8mp2Eo0LgybmJB9r98VVL
3J3e/vF2jGd/V8ucp4Iziocg2XWERf2g69MqP6xZxvtUVKozGFe2ZDy61iG9dIgE
f8N+ExFKEUWUVGSbe7L7/pCedMwe9WYcL/tPSS5Jjx++B2/z3Ofdsym2DmzmydiX
8SaN+o2cgBRlqTl5mSxNdzdSSr7s43xvSg5IWywviz/5xhqR2a1PLDrCfe9xJsuX
BEUUmqrmrltcZOmyorgABH5WbLIc66qxnZZVze99O0FV7xYNrJVcgRAbROiUKyqS
ido7qgV4CMIiMZYg2GqLomVDv/zxeb9dndzqDYYUpREMyzq0zj7zg6xVr6Q79LEO
bvQrbmIIEBQFWNLe+y3nxGrBhSYCLA5M4Hh8Qpf9LXFjV818l6auG/w1UtV1gq2l
YHUYJvm/W/E+AUi3wuG3uq8Vw3vGATg3gL7+H8qLZYJl2gXDb46/7RS8b0Bx6PI9
HSEti5+k5o73QgDxnbJIiEmCJDwPLmexo7UZk8Bz0qipt8tCEKLpTLtzVE6zpgcI
lsvLERkGhlxcEm7rSxBYP6fXYlycJ/RqqFAiXjL1Op/Ta1q5rHu1C9Vi66S8Wgjb
EbiKRO71iL+PCS0+ukGmGwHp5PI0WVA4vPaXGjP7iKaV92TzbdYO38pdm/4aM5/Y
nCe3nETUgD5sDbTsN70KhmrzUh4xkFb4o34q/yjXL/a51271zsubv0tSYYrBqx1R
uLCHsSwSL52FzNM4EzRtgTNMUGUWmBziOHw6kj7b272hCpwEYiT886ByDloYcaj4
Ct8zhVzhpQ09FidW0A5AbALS28R3CGdAC6V4UnquSpRzcoFRN4rZB5q8siEKHUOn
OBuSMdZzhuJphG8aYHnxi6RwHySOryHyRD4wOdVKFPjWj6/YDmjRfMIoCWP3gtUZ
sRsOuM0jDKjyaie3MTv8yYRV7llWjxhT0zZs7xi71qnm6yXnMiRoy5XPovQ7E88A
/5D3Ec4l0VF2YaMXeWflmIMG0iwuyuu/WBicQVOJ9vt9vq3i+yTZrMdrx15mD5gq
g+LmKyJgkVfVXqXjT1d15gsNMxfXmgfEMEicA9Nal4//9BzWbYhipQdnYp3bQqa3
lCm8kiHijBg28sbhq0+urJdX5PKL9NB1bT/U6BFu4zsRQFx/mtuqBjKkVHk7BSFn
8tEKI97IR6Mf7ys/TnZpq5xunpuG1a7yMrSal5q/LJVKOBoBr/PmKimER7JSg7lP
8V5yijZ8ApQDo845d7JfoaGX/zd52VU8MYsuSi1HyJERTGSSVWuf6TDDWqiZ0d0t
CLYlb9t5mZ4B4CxJezfpO/4sG0WyW7FiQvWSFtZmhJiQnkwSqysOcQAVz5W/N7kS
I+afd8/vWU0PCOMSlyDtLBcsOsAB+V8Y+bm5t4xH30cxvTUTo6sPStUpAnX7Xsgh
j/3gdpT+WWD9/rWcun6Yq1wowLXJIS3t+jg6pGmx/JUAUF6lQRrsyyV/Aj1klkTM
Urw+gpXh8KHNXQg1Lb+hwPPlHb3M8r3mMwuFmF2Y7KgQ6mF1EHc1o83Ic/Zg7V5u
4OCjESsyWDp3BW1jcMtVnHH0ywPqRohyXCYEufcOnjlxWS6D+Kv5ccvAIV/b/n6x
9WFAvKOBBhFYQJPVxiO/wMQown9QMcuQ5h3sHUbKS5rNBTqvBNDG10sJk+A97PE/
F03nGUOOtMlASM2c3043Pg6/+LxjbpJafe9gdVJh+XAIDH5qU9tHgS5rLrNcAL5P
NSvVAurkjLrndsrYtiMNF67JDypgO9Ymbv5x8mXHJY021ZNaufUaJ+mub7PygDV6
FJaQu6RcC03L0LjB/iPi4TQXUiPuP7eQd6apomkJQSvn7/Glg/L2foEj9N54EL4o
2A2Yga7iGZgzCwA+fRxQO2urz0SCoYAKsj+5iam2fFm7VoKvwFKBtLNCURYzPerL
HPRzsDeNe9EclGBtVEMkrkT7ESB6jXaK7tZs+dRqKnVBKWlZTaTTA86ETG6fSM7l
oE6lLYERCS/yRoMFsH2y8juTlaVzfuUA+dJBBplD5m2fzCcTwODs2tYPe3glSo2t
UB5tUV43ZdFNT8UdnKZp7t3LeqhZAc+tEi+KY5OKQ+0QdSiWWvobb+YZ1edgYU4x
nFkFsKbnbWqBLnDWC02svn/L+0fWybgUlFEZ73TqcxBDoZ4JYRspNUvqv0TBSygc
8R18C9jI6P9sNibIJFXJsImuZyXNy9SiQFvUwmyJVNHPYvjAu0ihfHVEiTyENZ8V
+av6HGaHcE8tft4+uQ1xKL1fCkaYeqoFVffhpIIG5W7rQe+rx1qwYGoc4yBMhW5C
CLHDukkqbSbIp8U1jC30Dhk+9fZOW4KqZkyasPUJNzK4UkP+Oumi7kSJWAtKlYqg
DNRuaKgA+NpSS6MUvIFfQZ5iqvdn2+RZxYwPVq1dGeWSGUIia/AKG6rmxN9qIIEn
2BzaibBrw5W0jGU31JsQSDX+UDp5lE5UhkBSoH5Rzrz4bucSa1GWiIK+Ztv5bfv+
X1Wg66EdMHG5C3c4FPFML/PLZs7lAkgwuMdaQOVufvWmncYB5coaQo6Lk0+nPmET
25NmUezA5bcqf28cr60j9dbLXIygH88tWwtQnhrys80/h52cRUWjayVyJleUBPhP
ccCyxbkjeVxmJ6ytN0PiUMyOzB19/sEj4yOXlji9HH56dDpw0Rp5HYRcougGA8/b
N6JNFF50G4hZQgyh8X5Wfy2Bqll0WcSxRd34V7uuEFOrHtCzVnRhGMUAvZbgktok
g0PG0IAN0uUoKCYCBajdlTkwJMtJmPyvgtuZHm4/r3DcncmvJs6FIcmcK27h6A/p
8UueCq5eh6+CwZyTiHWchpJsWb7Osopuv3qEInFM9OeufhP7FJc8kTo2bQjGKobz
XmPAkz19QRD4TAsRgWveZOD7LaBFC+zwQOpRpjnXuRXrP/tSs/GoMu/vgAe+z8Qb
vLPAkSOkW7pKAw02C1EugskuLdJQ0GXXTR7JcskNP0rKw6CAsPhh7AZXSxudpozg
Xb4BhKhvQ3O8lG9ML9rkUSN1HqZV/KNvs7x4gfdUazuBpWHZArDH8gZYg+B+F1Xj
Htg0fqEC4oR5DBNklJHE0FWPGazEZkd5jRy6CQP4QH6fQFEedjNMRDVUf/V2oxfl
ebmlq1N9a7EoANstmt0G7AuVO/2VJMBCkks+kq2bpZFAhHBUt0cob9XhgVfIgqKn
MLePQSBHSVKrWeZ7U0OsP9Df9dtRdmQM1yZQ7bt4axotI7e87Q6QovTzjSUbUB63
G2GNDR9GmOHpdSqfGl3zMa+sqOuF8/9+MtKA5+34OPtzjtGG2TtvyM3l4FZSfwGu
aGxhI1H9vnRSAqK/ow9apqdMXcJsmQe1uGCbkGP2BXH+4n9MhTxM7Frw0OgjMlvc
FRVeTQY2V1GFucogTaQxk/oDBj47bYkJmVXl16Q3fNM5U16u2NGHuPR3x5Co69eD
8F5HzYm1fyxzmbST5Od+YuFNpO2EASFYr8KLUhisLN8Tpqp/GYcLq9Fqf5aOK0yW
R8cf10knz+SvB7AcKf4gZF77+bm1Ybt3c6SF6mRUxYMTWNYlLrkuEE4NYCVvoEAr
Ye1n4GLDctt+HT0SJp6coEAurMfsMn5dWzQzWY0bT9SscsbeNzaXNnhbucZwNY8g
BaTjMheW/nNDj6ySQoII6RAYdu0JaY7kKHRD/gUrQiPX8LJhJDw4Nk5lyydKQPe0
15+BXlYmtGbpxkgiChUhXndUyj5xA62T9RYnN/LvFjMiVL80/vKllzhPPzQzYjDZ
Ylxx6yeMBRDY8A6nCW/kibQSnBucRwjtUmNRUxKS5XY3Lu9vcJIrSwrOw9zEOLLq
ADjbaDbNdFBDwH/f4wzOwoENA9QVk59qNnT+raOHCnVWqeP6ne713F6g2d1qAGBZ
J/hq73Y9UUkbzqIu0iGP7j33e/RLKnpf4wf4bd17Gc1ycSRRl75aEi3cPDreokGa
JO4MMesQy4eNNcq4lpw0PETi3SAjO63y0S9a7RLrvFpjYYje0cAA4lhxTDU4xqHL
ZvN1EJbZfzUO0NnD/3HRHBXPoDO/mlY6mvtEZdks2iAyIUGLGY+0cNMZ1NsqdWwx
WM33GjUp/IWL/HHuHJPp4nLySiM11ydaAxJzSYTErCgjT1wM7GeWulHppLvylNQH
L/kcRnwVR7tvHgITPvYTxPqDVx88g/aX+imOKm/ksrktIMg92K5IZYazP/K2jk+w
xD20Y+jmI0/EtabUE0X2A6Y8lV/Se0cdp0kzReyfGcO5WTGRFLXGgg5eVzwy63Dy
cubs+NXwhhkfO5jo31zRHH8BXYbHCIUmsWY5u4ouNMhPV9nObgdwsQnZVP17qwll
9BZ21xAWDDt2TF0Nz1k8PnriGPU3elBeY8rq2ZhGe0H0n8xkmFSGa/HYYDXkNX+n
6plfypAitfvbCxZNi1lwmc0uN0gFe2UZovi6MODg7bMHntLdQhrLYFSC9jHfS4jj
3aaP2z/nAAjclIs0kmeJNTrM3aM2H9UuVNzsGhixLtIHxibydoAmv2MHj5k8Oyp1
2QvioSFwRpwIUQEjAdCkepupittVg5HetayceJnPeX71A5fxnAUcVa8OY4RO/2DJ
UrZbTq94ROebZ9Lt2mo6sL4zhRML+U7/c90cHD9LLESXwoWkznKUcMqk4tsVmzy8
RDlrAIYlxnNgZW5J35oCdXdBTi4Wztpc37MBHJbRKSitLeIylHBi3O9w3+U6C5Vo
I/fXW2SvMJDzOd0VP1Gc9uESysPSHItyfXMvGW+jFU2wJ+zy4ZFkuNerZq912t05
0tbXQGNAQJsAfxkdhSzk+CbCdXFSCQaKH7B9c4j8z2j1Q8P6IquwpF59P2k5Wzak
ncgmcg9agejFLC2D8jBZckHf1oqTTtpEKHDPmm1xWVoA+CPrKjeR2BJ2E/Tp6CQC
bycbvXzCYa0h8WgHPpI3Ed27iyx8okVP1VJMIIRiulwalJuF9XDU1zquJyJZlOVi
YEXNBkmT33lsVjFYWJcmuHoj83OmA9y94e11RnAY9VE+xe42++GaVu9M23ApBdfq
HQoTK6V1xd0FZQwdYSP+A/OTrKEMp3j41/8IJchnoYz/PTVUcZpyiZfl+yFhi/ax
FECFB8m7Ox5H2nu1cXSWRMIpHL91u5rXj/6n73OlNelo6RU/2goCPTkwLf9mcboI
XC0Y878WuUCMQWgmMmE+WAr/M90LlP+zcET/D9nmOsVqvHuCIY0r7JWYKrPTI/VH
QZgdY0M0hkG7QpYs8BmH8903TlpF2JOxFxAzNY9YRfvozx/PZF0b/aRyg2hwym9d
OjvWHZVgL+uL5eiNwtIwshlzDpURCBcMlYIcMiie5KI6CSSsLdzKUxudGrGizvFi
MWqquVFOecKzNS7f4z2DsmmO83mVrXwL6H6N0so2JlOshNp1omOAks68bPhrFQwy
uBBdanc7i/nwO4duqpjNJi/wCuhtrkV0HHbXwduhCBKqVeaJSncSHPzNn6SoY+Vk
PUhEfO6Nd22mOL4Yf7xJ8g4LiwE6uMb6icME9fXdeiq2GLa9kHQFELx183trM6ZV
vpK8nbw8xYsoKdGH5G/vERTzv23jJfS0axWFOgwtxlkvdCOxHp+UY+eSASO5GvOc
xG5xwIJK+qGl4OhpBvJmNtW4nNnuFIFcqtA/fPTvUNt/atS+xf+Itg6x7Y9tnEQ/
Acq0xtW+jbUpBHLynjAFYB6n9QxOuM4zs/OWKQF+jiABaHZXe0uA4zlxPAidQAdg
gmyAGI9WEP9BJEkKUTraxvp8uLzw2bbExC1IrC/BpLW+hsAufcBstTOiZ8fAQvfx
/tZdqZm7rWd09rhmqZi4ces38k3I1mtprU5RaRyec1K8Yc8pFzg1BUdnjTn00m0L
7gIyNGxjWdEUo7lvE/qppBr4gEnqkfzccHVpoPKe5Vk2gAElPwJ1AQ2jceG/GaLw
Hh+1FKpLZVwpnMtyRS45qdlv5LL9257FnzAyXI8EZyE2ONJHm+2Hpc4l45qEbUf1
ZAEFGjG6OfyOKgzdVCRjGZMvuyhHNkeWoHBhcyPn45fVt14aTaG/cVwzBp3hcVBj
9e2wdKiMx/eFZ9esJvtW+7HQ+9SjwqvGEA5HngHPu55hh3jzbjHOPPKHJLUcRLVk
A/UIClHqkMQ9kf90jKXjSD99ga/hPGrBJgcZwOi/6155d0inGYvLQlkSnjmsugTj
QJLTa74iAm3AwC/+7n3lWtPblWQhJDrJhLQ+X5Em9aIwQAfWDW4JeATmcAWbY9pM
1Dd+EzJ+DyLJ/8ecUHFmqbsj8D8FOQDym1nj8ZPleIrySUIFYtZEY7PfjZbJzGjL
Ly1EEAdAGkemAoyuYCpOFgeQwiMwt+e/4zoJFnCBZKFTbGCIThC6zcz2hnd5+8Q+
xxpgjLdKyIA3J2dx7EHVRkDZ8taH8Ze2JUn+CMGrfUwA/QiuJa+n4KeKnS35ZMKg
EXpzX9EekO4jCm0Oez7fXSNSg/jU9am4Zxq9PngkAEGmByJpqbeGTr7Cj+BB7Eif
zzKnOs9YeRibZO96jcmOLHbofDaaNK6OBBJondzyfMliD/+7TvyXOMfJLiB1AF0T
7ep//XyBE4OQqqrwqkqzIA/H/Rv9Tjz+EfGAmAnCRVPv50PbNP0lRxD1Q6s0QJQ1
5CFZ3duK3nEitoqnJhjIWApk5NO9Zb8Dy79VlOAAioCXt6QXmYwWYOl5HDMBUzVo
aDnQUjSS5B7faxCJ+ZvFgyD/XBR0MCk0dmrnysfoj9o3OVAezVIvRDaTe8xXfoCO
/2L+UKracYhDMRKq+l2Pjx4DwY/Bydnq+uYx8t6l6lmoDxomK6Ym/iTFerHDwRTO
umwyxNZ7+mFY2/IOFpZ9XnCXxjtRWoEFw5cKQxoO4wSu++BADCZaNO34zn4tSYLW
RCC9MDLQDlCYS4YALM56bmGSfanyfeFXH6uy1LNZ9rH9eXUvUDmuapYBzY3Ff6bw
xbTqV+162bJd4pK96CbKCtCCbkBDXNwjpqvO9F10IQ4AXki14mA/KRxBlPkhcmBG
nV+8TC42zLS+/JyLD8zZGZEFO/wZSByO7t4w6Fxm2AcLYGZy9rmD3jcVTbquigei
FNQeN8O56S8Dps/rlhCDpA+1qEoFy+jaPOC1mTpAPo9ljmvBfFlRNRtUMDGsoJyO
cZeacQIZbneIIvMKZwQF2Ah+W1gbvvNyTDg4o0DPpDeuVYdPJrJRkjn8i+Smim2V
3dQgqV3tV/bow9RlmQY2hAVni9G3qjczkdZn2tmGwj628iCH5mbt3pFo21Ix6mDg
BOCB2IMseruJcQueLKnLrBTpfkEtnDQMcFb+/AqOcioFcXIKINy447usrf1oaBaS
P5rbEMrleaqXf6c6NJOtMKcPKSPNJPulABBWWb13j+azkuT2K9sO12LQzvIuSN/Q
P71PYdQUzGNrjTjYr6fU2Y5o/mEAVRHTQSlo04R6x0gMIr+540YT9jVJwDRd+AhG
XECfU5hF1EZya2q2KXXjPmred/aIGN666uEl4zSVGBQOZD0iaHqzD8QaP9+rJtxm
kjp+6G9xrHzcMqTKiTxM57DnH3PnhW7VFvTSwDt59AaZF0kK6/rHkTYpCtMwHOxf
l2oqT2vyqC1V8Iw9cQc69OC/IraJvuh/xPGeglFgvjcQ1BFlVVePNk3SfAG5B5p6
XbzYuTYDY/JwJaCOskeaFKI7EYVZsaed2GHq8LqgDacuGdXTT/4wmZy7LcXo4F7A
ev4sUJJkC03yOcVEz6QE3y3seVoo5tZ6LpwUsNs1ARgHn9JOYUMVZMtHyDOS9hBE
4d0+6ovgSrybKPFe0OOS+D2X9RiBXE7jZOUzq8HlQHDKWkQRj9rwtxBZ85qHF3Uc
9Bq6jrFdThavmfqp7JrHls+TNLBdSTLuEckZDJGcsxHj8zO8lmALsbskU9mYjOu6
OoPsmgQ0TWdSSDTzP2Ej4ZAxumrT93d85h+luhHutBpAGbxKnWUQ8qqjf7K8EP6S
VcdVRh9qw/xHpIklx8aY2cAMUvuK3u8D2YX4PDo8O/yJSOIP645bn2dLfszXAVSG
rFj3P3i5N0kNWQ8FXgHN69jk7P455JVsjXuvsFZMCAV91gPCJ1PwU74Z2VisSLEt
CgbsaSlOnMGBvSR52dJ+YjR02pnRWx/txC55M2xvLAgaDtAs6/4i06vdzMninqAx
zPZC6yYJ+q5tEKiqZeAuBuBNNpNPeYdnglqgXU0XuwxPhkknO4ImJWPPg2rRIRZj
Q5Ji4G6iVoxaz+85YutptFhNKCL6nV0G731ytx2i4uyrcCUU7I5wfM5XFEySkGss
2NaEpml7O4kKRHcE9Wl4yjriZlW5X/RSxlVCjnIDFxidLEtOp1rgx4YN8c3GEckc
e4WOep5O6CWx2gmlCi6bf1ZGEgphT9hD2cqcsQ37+xNty0tYXSKd7G4NwRogxQl5
+JgO4LDvSwV/g5HPEkdBEU1YWTe4gm8tEWjzHMDbQO1ALeaBXAJ5a6PsL/CZTjhs
79PvXJpuLi6EmQP46QAY6iZdamafqBrMovAMDlTz5lYLySodsF2gIoa/53WQ6Jdm
DdS2h0sH8tsJuCUD5j+jA7ohOXZdEf3TiTzSFsaksouAk+zdHxIJQEwFtyvZ/NSE
Us7/kpbQh0cdnAhwsps5oPwEfivDAAZJwPm3y3peukxKenw4+wTDJ5HXjd/Wbu4V
31pAYv8krKKFifX0vr43TOfSXWOv6M1cYOsugQ6GD23JVhCgob27nGrgq+jjUQgj
5nArL5oFP3/ThJa/KW15bJAxXozm8WAiHxcNWepAmqIp4pRMLOmYfrLZ6J5r0yEw
b+L3W3SodwNYfnpxPpOlDQAUtnVNRBeTQoXL6q6/OlmJoQqL70Gj4us5UPEjWG+1
FPRPvVfLclEsLWEt/ZfAQdcdh+jMgAG4+wsYbmVKdFiCD90l/9CR4S4wvEkxTSOB
aGvEpugmqOa9A2UnyEQ2DSUPtmB957mhtjFxeh3DejGec+bGwqYuRfbWLzvxyBtB
TNqINHAYuEcDiuBaSifsixDsxCu+Jsl1XorejepXcbQO1xw96PUSGexv39VkBJAp
TkOm9z/Fgup8ae/5mJ7lOxEi3RIOsj+5bazX2NYdsK0E9yvOcYEfKh1pNi++i58p
qzWtfmwjW9KxfvFbPw72+vS2/9f28OKMveELASVRiid9cOfvEHjxQcI5FQqM3ISY
cbJHPVBbVU9cCzT7qOTkUY/Xu01LHRxnEI+i9ipSGEbksLW6yBwWlCWiszpIrjHr
eythRuX/XWpL6hAlRlYqZa/zqjUvh1Wmkzp2h7f/7get2AbtCnc+xqESrw/yLfT8
nd9qCgwP6y8exflGnrsbs2IUKJs8erru0U48STQcSUZKe64xO9VA7SzpiRd2VI/U
VaxuchNwWWWVvqoNYsG11gzXqrJ/AJwP/Nl32x76YbSHhHtx54LwKinRtMHKpj62
Bud5ewGvcoZeCaPgLfFh/4v/sCLdnceudWLWnZ0/cgLCGz/xcAvr2RiJ6y7bMSK7
G8ro9kxOmqpbu0KDM42RgXqQ+d2VpHsxYAlVmimn7Ocueh+udnAfggaXXHJvFfa7
vXsMibr1i268YzW3/zwhh9qEkGxedDW/+7LP3rauEd6smub8zRZ7czSieb1IAwFp
oafRDmqeCMh312RGGsQ9XJZ3T+4nn2/ENz/tKENpMlzO0IPKTgslFuH/Q5oAevN0
enqOWgZCTae1uy239py8hRpybtDFrAzhg8UyOuyKuICd+MBzD5L7dD8fToDeTwPF
nXC9u/b5vTTfxBsAHMl/3PmmU6+vDbflcY1HN3O5z6XFtc91n/am6nlqStQtWEQG
u7xU2kN6l1EtZiQiibQ0sRpSsarGE0nSHOV9wHK2QMX9sAXGmZjS48whAkVPmKJf
i4yQXM1MNacVq+A1irkx2tbOGRm74Sn5/Grg7vC1Em1FLCz8vs1CbZMByAfA5KeT
U0/CY82NUDEZIEAHQoIpcoh2iZeMAXbInbpE9HnGVhEbEDsRWcV6YcptxlQOe/qV
UE45fPNRuX1XpDalT247yqRS+x4IX1xDsvN5jowU6A340RLnQc744wWdkVuMaLEJ
LjFJi3+JdwvlexPC1lLRnXO9hgXo1tDqYfqWLP7jQcG2iSe7sQMZTgsh3WDTehRz
g+OMTM5plrI2fSb0VYTC1gt3AsF0mv8nUKl4G11mRJq1N2vA7TqRuyF+d9bj1e4Z
1g/0Wpjz8uiZUoEHazJP7ho7mrWKFB9UE2ctZv/ephT4DP+a+1bUVsj1XGUVFTEC
l0p60TCBK+SbLQWdI4txmRbsUQJaYzHIu6sntER+VCpVFEyhi4hYuGMWyHl6OLvW
8wUlXYbuFOxu07I/H2NyhlkI/lPWJvZhohXTnMtHoFUSC1xOQNmEc1V1k2P+twXT
ah/7IJ4DN4TX+LJfRHrTKGy8pX86wEKFHeiR6bsDCdFk7czJPkdnTtlphKHb8lod
NPGdmIjW1gkwhqIy2bI0oI8nLiniPY8w76OStCOXw4U+kexqdAXDplFXL6w0Z0cu
9n1Lvfjl7u/neuguybA82CXesD7i3kONWzhmarHQdC+4ZtzpZvkY8v4dekBjHNot
tDkASUyqe53sBAr1C03h6yZTZ8A+Sq4QSWji+F5lDEc2hf5ARVTMLTNQ6F5pqMMD
lc7Zw/RQ7FaB1F6feZ5kDnFan5Hvu/dbkl3g7dkKEYPWZsyf/y2ElnSYkrAfTFyU
a+YZs5CZ9r3EWje4k4IitWUj4BaxTKf7yVuEuqF4zlS1U7AxVd6XM9d6N+zLDN0b
/pmPK1S+JC8yOFDCSYr2Ivd8z3+slDPdpqAx769Hut5NAVAqpuaLTUsp5kuskEIo
UtcxadNESE20BYg7vKZj0Lqdamrf/aQl/n/IXBTurthRLd32Yh7nXZHjXRpfvd/n
5qh55H+zl6uJE2VAyusBMKogBfdElt6svBUmm+ZYqzeCqqV5pM+RAhrt0m+Givvj
SFaxofL96bmavO0uefZvTOcL9oP3l7mqFHv0zmwWvAXFwi/H9cKadwgIjDN0HJou
utFT0ofNshQP0mULC59aWwQYi+k2B+2WP/tuzsGpepNukn9AdmpdKDT358jw/P8w
yJjPyHM/LtvcF4gbOgI2ntW4ACZmrL1ai+NO8W2Ps7yAgCsRw59U982sPRg5XRdx
ZAZ8NvV0Rsd1xikw1GCthCyAh2wA+ND2bwdtWg3m1pte4BmT9IcrnD4ckUqC5ExO
/AI3poNYZ1tjJe4bf5ekVMUbbsDHL5lIxvNCHY4eHEgL1786lAVutwh6MzBh8Riu
4gV3emOUxNrVuj/3vf/yBX8q9BjEm8zTl9+qqZ3ltx+bk1Ec63C2ER+pzrL2rtYb
pxoqwiurEX/tGhNAuwW+5vjjGSkpx/6MUbtVVEzbzGlUNAcNvyTUEs7T1CW6TIFP
UTinQjlUyg1oNkuPEiSgOa+9VSDACUqhkkXZM+5p+jSdW5EUWyOfiDk45QFqZ/EG
lLyncma4Ymcq4dkZ+lINKK0WBA3DOofBKwquMBKeVfr3VT+MGamlZaXR8uoe+CmV
dR5hjNxQKAJ/xFBnYr+PKvYojcM6ZSL6UBropXZ0jBFgt5Ymi82/Fzh21JRHuNqY
LEu3M50OiC2pzPYMAefVuY+HTegeNoVBzjCTCGO3GJG/Ss7d4eKnIv5QIHJTWRQs
tcl8J2w1RpJ8lHjBrP2Y5sm15HIRIDKmQkfyaoKJzg40d9iXMr04tVTRhPuc9Fkt
R7DjGfv4As9t0VJGEjfUjqp90fKIQYIqCbkXi+/c+kgT+3yN8OtTJhmQJK2VhkOg
WbPn/C2ai4MLrs9qvhwMvIVDT4yCWImwspZ0e8ecupHbV13XxbmLS2FLsRiDA1rS
Eon6GbjbNqCp3TKwuVbFbL1X7qUueOYkJzBxoQ+BtBpLIVL1SvI95JHGY2z2DyOF
4pRif+9pLU4JeIZdRYIOICGFfZX5aQwXTULi+RrKtm7fxNcm7YsbNXO7IRUjw5LN
Iq18ZsifZ3iAd0gqJ69tsABSgGZYS4yqSaOYEO78+KDlH+PH+hJh0CE1lmQvgkct
Iz7rXvIHP41+01JCBBJjXoCgFXyj6E3CqWI8NJU5nbhstsglu3QomAF1SNHedmJq
7IvqCsg64AsRhLWsjOv5K00ZG8m3hqE5DfeYp1gxLMowNLOIfCVBO2psDnvnihE0
rwjLjj3xrLgo70QQPu/dG+bMAMwX/OpTCnaDWeeYAFdy6hKa9aLO9qTXa+JFm7Mc
4w3vXWRghrBSn3s1yYc+5hm9rnUE3YCVgCKNF1NGlyMFyHfB2Pb0oOC4e4L3JBC+
GbCK8fdevgLlMPuZJAaxMg/RKSkBQ8f/JcQMBGqh00Cui/U9ROIH/pliTz+EGK7w
uk7erUn56GelxHAvltziszDVMPEyz6D8nwhSckp2XwVaAFlEULNpREEPmoA81y7D
KCGL+goxiZik7holrwlzGTh51wPj6IL1aq0eunsnNIOxTXA35ir6r3LHIpEKfkmy
sWS+Eh1l2krRqN7pqE2m1c3f8wntc3hAvzSR6bOlRkdl5VG/YXSVsJLI6uIhmd6p
Li5gSW6izSoedOU9rlR+9UGfFxysfiCFVOwhy1C5mekigbtTvHjyxqtPpIgADK7S
Mii3LWrXXUQ4kf5tLYvceCkphNXvM2Pwml/0c+prpG45BdOKFESFBKC/tx50kUo9
AI5O9pvEOD2HjN2HsfPguhT6z0teMusHeg9yIuZzRcdqNDUsvr8yFa2jlTVSF/Z9
f7Lq62/AG4yZDKfpC8P2ULITfB3bp1F/FvaDAtf0ia/d6T1bm5gbL09dx2my4ZJD
2vG/xpib1HCwrsbPyL7MkLx6Qf6N0VYxjIiZjyu4eoQE3OrjQ+0ZaUG/ISbiZHgb
l2ZVquQhjGJ9QDKUimpkuCw8k0aHvK8lGGQlJyVYa5u0PaB24j6KCwQAPdxdoONJ
YvLAFA6Sc9984y8weOFvTaUt2lJIpikn3uAMKmUbgK+KHnndN8AkJOiaRC51Zuqx
U9Jjrxw/UcXq06XCZNKVuffZCq+J2gBvuLKlnmsKeWgYrnQKCqPRdu9pn0xoCAlk
qpQp1VugGd8BdXCIT2OAjA65mLJromTrrlve2Q48YydhLHWgAaObhZZy4jDmT2QG
oNknSKqK0fiTRmWqxLnKOme7dYij9iGn9tfi52BqkdpjwtGWn6o/+ciXOtQkSVch
rtBizrxDhL59WWm37RqxYViBr1Iwmd2qmKleVPcZWmqNkKbCZ00NeBC4C52fK8fq
C55StZOGRz9VtD1XP2qBb+gyi4+2T8MuuRSkPSsaR94U+Ryb63fFftgdx7OMNrEe
RBtRQrbI+YA9K3Ij/wgDg0zrLinyvUCFhhS1JoAV7joxa6WOPNKCZJLc3lhE9G5r
bdMyn6+u2DkrnFNPG5tAnerXAmAHhQl73gcdEZw6WdFUO3nTeEDIcYf5XYPr/JZl
E7RNVl2YTxYzxTxmrsCSwC/DbHNGxU0zJBHticQAAsF8MSAeY0NbE4dV/vJ0u7ZZ
nzysYkWqpvkQstngptqmgvy8rG3/PEYtDSIJyxsNu99/3mhuBC9CxEDdROc6m2DW
DgNcK59N1EodwtsfeDBkZ0VHdGMgQXXB2EAA0HLXwDnqJ5Hqv9tK8I2+oTWBDBJl
M/iHDh23scYpDqOAJgfM8X0TOO8FHGT2pquGx0/19ZIjcGwq7oLU1/QCUT+wsHN5
+ToMrEmTMfmfL4JDMcLzH200KizYpdqVifGetswCOZ+HLKpKkf7j0jTD6gMJbUie
Q7CHFYbIu6zMIayvHBkX6SOfkdsEQ7O36N0vldk0EFUPSIjohBgYUf3TuMTRGLS4
zphLZxrMo9MUuXNYHIl9eGvGhywwPGgELxradkRx6kSd3yN4UVTaTVnauvRkou0O
OfDnqzUKkCQO2D7SCWvluplCyMc0GLAMXwvGIH+iTHSnXWTVLemKL1iCyEFX3P+A
ysUsC6QLZKspzF6tiNrF2eisjZ3ySiP5SwgnaB2Td1WNSdDQs5I+Xcy1ztObY/wP
y09HFFKVFj/4sv+5iA0nhAnEzdaf4f/o6Bt6KzbqkLXteEx1WPBcXbqfemDqolUx
JosuTDKq12hZ0YcoQx3l22GVw4h13KfI39FV4EBlimLy+yM3YsBERzRnM5hYJ1RY
J34+3X4j/CVQPyv3t52lik0jodu/a7gcsvvaP/3A8lycCJpELyy4YnS1BTtENzTH
2DGjKrNEdfqU+xQxPaUJsezqwGw57AN7UovW3x3tstZbPdHRdfvpjQ/YU6CO844+
xmSlCIsWtFaHwd+DW6Mw0RCcUQ1lKVlmtXyl2CjzHeAMIgRNkuPbRNUeyB0j+lds
gTS9mwfIXlVQVsAZZawRl4NU9GKobVAUQxsHaTOf4oElla+xfP4KbMw9eU28Q2Q5
A3PxyjYimdOTaJtckpFeUANxp/uCelnGathnsLHFXyGNQaWnnrGEcunNEZTJk5ih
6pl3vXhRnaZN9TcNUkc0fqRTynLNdBkleJG7KHP2FNuOQp2klA5Now8+ey2Ltv06
FoJGB+SwxcdzXiGsveJFb3tUmjp7HPs+eyx3BRxP7NuzsnKbwsXMb4xyVfUmcLuI
7Dk3x6Qup7G4P65Vc3tcAgGJNALnYILyklmPanp80xoHw87woyMkKn23PG5YGIKu
4qqL0rx+V2hqlza5zY8c/svWgFVXZXQWFef/ChfD/pOk7Kfe9u2QnP7Nk0a2aeIF
nwqCljc93DRlWF/XDyL2/x38xOu4yh1cH2TPFS+LgpPH0l0mCiGVENo4/AuDegSy
Acikurm6KBsBzX9DnX/IZMFbiQJE4Vxk3cNjDdEgHBLBjyLLsFWiwc0eB7sy8CLM
ts/Bz9sIDAKeDbHSEabz9ExC3vPpDhgibSBzi3A8+FFnN36e2I/0arvubFeGLG4Z
VQgVZ4V6oUV0sGGmmmbuWlZhcHWjah8k+75rnzrPTQe+Tw4XEeiHiqMoag3pRF/o
kzIhFLAvDhuI/8JM6xzwlprG8Lu7Sfx3vkwaMdZJGaipbHbZDs6ShaN1Adnt6kyk
hftg+Fu4BnnvlEV7fhfgrWnv7ffQ2i1ZY6BxmwMQstjuL/gZKXh/xjTj/Nhb+S4t
I0Cwr0tRnR7N2DR4ZjBjw4O5aCbTgubqoUvkKh1cMO47w6VzsDwIXknHJkQN4Tqr
xRkFRXO8UGcPyWDnHYVD3hr6+Y3CJI2JX2y24y1K+KNjQI2hblLpmYHAItKiajC4
dNVEbngQGJZr+oklnly4h81sIHGgPJbokIJj8X+TNKy5CQ0Ts36IvyIOeQRwLcjV
wnNIYSLeK5r39NHvou3SiFcp2In1ydzC12ohNmRfc7ZiP8kp/Yu188Awt1pa+GUG
rDnyQXeeC0g8ga+MHKMNytYWEuHyup9yKzMow7LxDY3PvkB10DiwHKSzinDo04Rw
RdhC2WvTQV5isODEmgslinGiLBOrYmn2Fd27ux+5w2MJNG/n6AqxwewnJd+uBSWP
NUC4EDjYxzsEsP6QE6Zu2Yb1bqzNUr/15JQytk7yC7iwlC53mnIdeDONmz9NTNfR
5Q7Rzifci8QWdXrDNT0QA75qRVJMbhxPWEGQ2MnsB4tYyPQF4JyrJtWaF9JI8Zus
C5KFeH+gflMxqpK93hzJC8Bi2NGw5xmrGtsfjmLgvOi6YqK4N126uGW1DBecqYhl
vQomjNfqqwoiratD07ncHv7sGjjzVee417b98f7oXyVg/B+oiUE9GD8/nCuc6BsF
jdX1uj+BI6aAMHEJKhPTUIlJsBK8qBX0aGTWzJN26nZu8UPVq8l6tu3QRRCH2E4d
zINIsUaWBQ7T9hWerdXBnQx61TXWyE4yvLNkxMWFYlRixZ+MmJVOO0je4CJqdW7u
KPylfpwif16Cg5zoQd3iDsLkJZRabh/rGs5494KgR2wtrx2Fa8QUzhHEQAJwFWtz
gO6DCPu4vL8cPeUtMoUaMbx90JdBIbgkkkIJ2bu5cQRY0ZLUaAfFnzy9okg8OgBg
0r6PQw6YHtFuWtYqS4SKqxZ+R0dx+PXnYCCd/N71e21nxuTKyDus25sK3rBdOMYl
CxgYfe0sGdj0xIJoDrkb+KSHLAj/NtrEE2npISEeoCU8vFELcscoUrFPPBPv0OgY
18BFNs4DxEfvx9+L9zRvjLqrVG1i1KynN/+cSVrMETZD9N7MFE9N2gKmfSlVQwjl
tGyw9AAW3a16CTqDAeGZH7tRciLdZr1vhCI7zBDoW0MBk7efV90fQfaKYh2F017n
YVnLNFkrrxdZiSODpOrL6Imk6+BmrXd6TbLg5obCRX1MbLJtL23rGdK/C5+cyKLL
FnPjxC0hRL6y3t6zMYAPruiI4qGEaLO817C0s0Fd+jULjxw/MGYBjFuglmPK+Ed0
+1RLLOSe0NTrL+nZt6lydxeZ1h4mjBRdvmVsmKd16FpKPET8l5NO4hXPbuMzsDh/
+WFCnXnjXIzcfumi89A3Caf78jipZ270gQbRWA711OzaJ3dsb7rs2v7IJwxFtmmY
v0lA73DLcWBoTdAUgM2PM31F4mFNc7VDg00xR71MyP6YK8giOGMDPhR/KnKMx8AZ
VbnemfqMXts+UgpP9ABScQDcN+/hwcYPNDEwosjXadE/d7rT5y6pVvw+eR0IhHzr
Doxj+NaF7I0EFY4HqqvWSw6vzTBhyrqmf0/taZwNHBeKCvPo9Rc7r+GUHYC8ny1O
62/+iBR/PduMp0pRnSOHWVUO2sDoH4HXm6pm7Jh/jnxWi30+qVAIqbn+v6cXtqN3
CjeIWhdnzWpz6UMmxJCbGo1UM2SUqaRYLeAzoUUysrBU3PBq9UT23YXsEnkKiksp
4NX5PmVjtQCodQcZyJUQMeoxrx5zNxziQp86BNgEgycDy8IUshoyMQXHvRNDtuaf
nb8MJRa9PfsxbKKoNORD78iWapT7eZ6i+zgiOhdch3ESj/WCob1FPUK2hSYzCVqH
QCqmwN3TvDTFNch9F35jtVWzRIEOHwip6LmQD0zPhqlBsRahmjd9bwzdkhuLLZke
E0IhN0AE7ZQKsbMixrR0Rrs14jlCQqywKECjwfZbEzfxMFzKyV8j4wbwdchtvwU9
asYuUeynZvahbuVUmFJ6WsFBZCnFPzCJ2Yuw+D8J1YCyJgUDkN4iPTXy52LogQkY
1yvTv80cHbNTpiX3HIQQ2HXVxyrVV+tULVmlbcFkJFWxy5ycwmQJgBV74bT7TYk5
z8UiNDlj+vJa1JAZtK6RILgsmzJsZGRel81sljvVojPlOqA2J6jS0o8z3Z/KiwJx
nmc6eEQWtMXoy3d4hCkWHIWMll483GQx+ukpPCVzhIHl5pJfXaGYONx9HA8mMouH
rPqT2YKUMbMulxL1wHihiMHct+aVzWbYxs4szd4HM/5XG9ZbegN4JDUhVHGH1CCe
zc6IfutwWY5Q01QfJtc1PLN/Q2o31+4or9jQsU/rVta2xdDY+k5lod4QGLpbQHWR
tu/PfTf2TNQdc4ak2oBd9IKpFTVWJj2JRAqzmlRszt5Dut4xkFOjp7KfnMeBnaVe
DO/37Pod9hRIFmGaEmCfBExbi/J1dLl/0QwucBz07Toaglq0fEot/hsiZqfX+08d
34F8VRyt4vxbWlyYHHKbFsNradzezqQGvTK/uakCTbuiGAN+xmXflb1blMon13VU
vrGTpFOf844w1XbuRaQ2W9ZahwNlEV8CZS68bx2wd9JVAU8CM9m0nxZVlKkcgT5R
wCA5Hj/jBBYBK2b+6zxOf2pomVmGLLqmDKMTQ52yymnWLpCincQ3iLB2ZJgzj5hC
agASeAt+IEM4FkLTfj1Lx97xQlp6Z3TbRTlz1YAmTsWkXvprjJbOjWD22u+ik6Sr
N85WR3lzGn+JDLSoVH6vz7RAfTr3ypSfQpMaicAw6xP6GKnD7/xNdE+ys/ZbgbU9
DvHR62EpsiyX3vhD5gMklr0sXNDL4nN/hfGQDVOMj0V8trfAdS8ozq8zTVibCMMu
6uNFRWa3G+0G/Ti8LT2/Q2a7M+i99MPIWc7VPMDb7CbTT16WMKLKmdIeRHEJoIT+
BHKXpQpzcr5CH1cYHnPZ1lzAcLIW3WETg2kBNjE4WseWPLsPDQkCKWZx69Wb2f8O
uB5C32aPRK4jOfGJwt4J5NkeLaJNfx1Q5QZqFWoCwJHsSEhW4CBFK5x0QhyjTawE
ZLXmkdU173hrTHYi+NJ5/gOlwNiv3vaOVtYLfAikRrIfvE+dSCJrZo5qi8RgtkTP
+Yh24DDeFnpMJ+/wK2cludAO5ES0Bdvra7lVVFMeb9dAGtjCH8XGUcCUgfStZmhj
Gs/zFgUqxprswnNqtZMWNhbboLUFDGz8Ila81mdO/8vJT8kLdRlAEi7zDi8THAz0
shKBtxNXBAAZrJZ3PM9byv6CtkJIv7WfpuIpHpipNrzqeg8snuhzcmTLZVzyLUnC
gUDRh5Lf37lzLx956v+DfBrcggVBy3rI+z8DsHjgCiK3lJBYalUpODF/bf9drMfY
ApcIAosnFNo/69mrBHymuRSNEzecRpnXTyPy0e+kLB6+1Yux+MR/h4m+4ar97nBb
35JTtnNeTJh+xGB9o45inqAHl5It1YJixKInPYWImt69uSBsy5oHezWGWvnuBMCz
etRAyFyyOznlsZIALqNw9eCDFUIFOanoW2S2yGu/2/wgaMxJOAAIYXGzifdEfhKP
S9nyIpMpIln+VNdNHXGf/csDOAmWy72t//eX6ImEy2I/FJ6kyG84YGeCYxxi04ZY
bzsiTj/mj/AAqryBljr2ZvQQdDwUFWXgbjztTStDMmOlJtQw7VEc/zpHVLtca+RY
b36pKVgqcr6iX8UEG0YQg8QVpmMi3YMLUDdEup3os8YHNcVtpiLdLjf4RExy1Z1y
x0BIUr2g8KOdJGqcqse41R7g56sowLAcGlyqI5CFpLgWYWj6qv1aANTOoo59uFpE
xjsjeY7lu8Sh8quSdyZzsmzUGG+IpfXm0o8wQU+NHI2mnRabO0cUxq220C15AFzO
MHnUhaz4oZQZAmvwezA0ycneu8aZI40qlyUJdw1VvxgbKzAqCRkuJTbDSOIDZxhI
V7k2jlRtKF3ERccbEKl4hfwkCbUKdMdUdy7lFn5Kz69q2l2qsgm+YNcOf8+EH2gW
x8M6kfZsXGEKqg5yiOWQFP/h8T0hVNrbpozRZZwclRcIITyUZbHH4qyuqfrMZYJA
oKmUK27oVmM9TCgxSFPH1uatCtO69qHgg9v3aoCtOZ3lLsZJjfrFWRcjGwWl7Qpq
LyPZQ6Vj/1H6u9ZEs+pEBhM9vI4+krVVW6Nu87Y1R3rSSiK8BIYCj9g7UI9JbOog
C4HiTRVX2k/p9Way5E3eNEm4nuZAmhoCBHf7Ge3vaLDAsGTTJcJO0Uz6WwRWZUbs
yd1dS/JMhgumJMIMD8e0nJM6pe1LEY16V/fbrOodoykSdn+vws2vGCLnPyyCGIV7
CmhQXTNLjBXSga2cP1470zhgY65w0/pTQfEmJEi7h7vM4VBym59rEsSBC9hPZRL+
ljykgxwha71K2PB5yy6iPc19FbRCL7Iy0gte28r6mfxsv/wSc6V/JRO2UCH0tKKv
ekaUWczwJQpNeBfi5UUuctfFZsetspMo8e69xQhPvX0v+T2QL1wTYX0IhFhGwvvm
wj0zphSyZd2hsBgfNMtWB+ALJNyIt51VFMqoG8PUoSzS2+e9/OsqgYRcT7o0/ZGz
7XhTW848wgOylOkgVgraQOWvmRbT614ROA6H+Rj5zJyeSKph7lo9nMyP7pGPMb9G
LyxKv2tbNYhvxR4ZjrhidsZW5M5rRv72NR58WMYOgtD3iIdQhvrnD93CGbNAmk6I
m1N4CEjq7QFyJwqFj28k/99tvIIdn68NGKv98ANSXtaSsdL5jqigXlP1KJ/YND8M
Paen+rPHdd2+wwwCJe7ENyLb1ZFfz4xoZNoxWQMkXyiTj8WPGVW7/xal81N0y4X4
UHiyhvvLgjDeP3X3gLkGUS8KLnkgWeSYX9Hlp8HZbgJNBbfWqd/ZazSXG5UdgW91
Xo8Z0YRGULyPpj40bOOQukxJt1TtJvHp7spguvG5WhV2NBETRJrpJDXmt/PXYr3a
Nf4CxP8/1p1mv2vUe+hPbdvjshiXLb+QzOFu0ruDIgEw3xjtcfKebrJwd2VQIRJ4
leh3GUnhbTitzYA9FLYcYbcksRd6NC2sdj8Vc4iFUwfDu0bzKiXf9cjN+bk9sdKh
1c5hK7iB9CTHeG4p3MD61pnwjbvoLfYO/OONv5hB7LSfG9DYXXxXFfDJsAlURRcQ
UWGKh3RuhDqWB79eOHSp/p075TL+xWFXsz3m41cVIyYHoRHGzUVPpMtmmB3JQ8zE
PZP3LwWI3IxrfSjHxLYYxcbGFJMIkoatPfCBOVitk6UozQgnvQ8tGSK0pzacBg8R
hZq6zygXk+6xGpVAy6AwbCm7QAOHBgcVFWYEfoaXAXS4E7d9BP3pY3ATTMLIxBgn
T1CB0qi6z1Y58NzBndy9Ne9KazTNtu4a5bfvkZwcbSYs5HdeNrGSzSLAAr+yCuwt
dTOI5HczvmtZYWIJuBATLkmnp5wNvoytOyEtEDoG6L2SfCBn1mpvsODdtAqe3JIE
6nBdVPMSMdYyzV5f8ZBS2gIJiAo9SsSIYCxPdj9UKYQ+E1vvWrwUL3H5NJCtmTqA
f3BlXFSuf3N6ozFQHICWyRxZJyGNhitUd0pITENf4KJCRix5xsyMKAI5HeKLsFPM
wR3dPQe9s3EH/peXHXOnx+IEmH8Nlp5ymjrCj8ND2y+I+IcyGyYIgtpPaR2OJV/G
+NAqgWNIw0ZCaVUG5IMD+NGP0JjRjo1JZdaFrvFfKkwlaL24PEYQbonfyeJuald8
JPHI3BdbtBH7RCPlc7Q2Ts3J8hefFkQtDlyr5UjSk0PIBobGdwgLXkuLQkFLgx0o
TFtyLKVw6fSfYgRlCjV8K8P0O+2WEALQ/lJzNkgxjmCjcSVOkglpAIjvAsOkdr57
Q7OT7/6pefiaFwGw92o9JjIgqVRWGCZ38GY0/21m9Ds0JmcXUSCHnxVEXMcDK9fe
mh849unDNuRJi9LjtXAByGE+U6I53wyBBEOUiGN/ISkvK1U1NcJ/19F0HYcsb2Qc
eHMfChWvP/f8WcmAUiTCPkitJm3J9uNqrXXb2gssbUim1tEMznIJO4OvEgA/1mjH
P/v+xIrTyevL+SAK/Cq8nqA4X2RHXjkNWWipDGJG/o6PVibm9l/4fS8jCuiy5pUb
fTwNNeSHGHkKqF63ijFcnpNX6CjYdLNc7gTm+YZDXA0dIxOk+TTc9V23CgzD/G3o
b1mwvE65ulin/BLEAmpjG7Kl8y/CKPUBlyq+2XhzNmEz/NlTbmZkSWwfHVjIM41S
q7m8XDOQwvssZMWCv41Hoc8ZXmV6mawwg29BD0vYLJ44/7jgN2VdDtLA+FJeOYXK
4JDgZTQ3yLMt1TwbUQuKoa/XWvR0oJHffjNsDilHGMQtbfHcWrQLk53bAMW10p/s
9lEAxuHiwa3T9/WzYyTJxCSh1foUv2K68wZX6zmKM7PpK4dtv7njEubSW9tHlHp3
8oWZKpD71cWW12111LU6UGkwHcuhXp4oKZU59Ntjgy7qCOK1yHwCXMSz4GXzWogY
g+BWEuYW5fxX9BczNHRKeiliaftzGqDvkXbnyroKgyJa3Ysf8dgTfVVBkl7E5Wnd
ViGNu8hiR+8KjqM7svb32f5XVNw8q02a4ekarU+muu7zYtwnQ9idcXRudCBhaPxc
rHtfrpHSUr2m5CTncgjBFgYQ6UzrrVB95spuPoyP7VvQhiLSKxQauGVLGDqmEfIy
LL7qBH5woldN9wnjRRXrJQz2F7tMAbCO2KKB56JaIcxAO2/Cmoskesn0WXUP9gy+
1fibw5/KHGcfMnAnemmDTFy+iYnUcBn/1Na1lyUulxHr1Je/8YxP2iM/cCj46Xgt
NfYyMTKEBPZsAGdMj4Z9rV3/QiFZg2PHoOO+QfUtxPX/0IL9TgUWo6kzVBkWfal8
nPLjpPtIocUUzgLGlRvSWS7AvKWmlLECEdXYLF7a//S3FZ0ylJhA/yRo/TMHz6G/
ecwLQWVMYjBLcs4e06RDplnZYxYWogiiD/lhnCuX014yM/iV/+IFqnUMQzlC1W6O
XRGBuVoKCOp8m0YRfPeStbfX/iBwZ4FwGLcC272tK/ZMmKblZ5Z2pgkf2WMNwz0c
D9B2mpw2POoPV47F+/m3L5wLK4mkuAfGzwiWIVSfDTWl6fvsoMKme5yYG3BEGZ5M
WApLyOhRJg1xciWE7Bpvr+73CqC8CME+oyprcbXFSS0qoxu/8KckPMzAsDFux0PO
Hh1/6u1aCy1uf/H+SY7H0atHLJs21PJSTagWxuOHbO2zkzHmLkHwMPEUxIGXSvBB
6YxoIjdpikaQGFsMwa+YRZjfa3f3mPdwvX7gPZTIo9rNdL6NsEdjyH4UGlfcPx++
cJQsJdZbqf9e+1bZpW3GdQIzaomTTwlWOKqYF5Xmv0jjbQzEEueu0Ei24UyWJVEU
YLLlSuWLltkDgZTO2/6GynpM1tTBJWNvg/foeWVv7KgPKPBUV5YpBrDFYMO7rLCk
vsL4QaIccPaTgKXGJT70xs4+BzGLLu509U0BbnOkAIydjpMpoB/jD+EsIySBjill
TVz0RA+tcgRoz1BEl7L7DdECcNxKUJGkoCUcPGcXZdhIbvZHdMVI+7ZE2J0IP42c
KABuv2eAf05WMeVEhKirU/FPolaLEti8og+tiOF3DPPXDu13bZWPMoYhf59KbbUU
LHqVmI33bLC4NJQ4E0CYVsCIvu96OsprRmRnC6VZt0lYzaLRPrMG/8k5b6LqpeG3
z14MKpuSD19AAiBQ9u2B+GCM4s8lTPZZta4/d/h8vFZdO3kWdB0FnVdhhF1FmPS5
8duVH+C3UwKrw8TGAelASXRxCPmVeGcvPvNCBvbwk8adqo0vP75uDrn6RMRMyG5x
bLpO2PN4ygGBF2pNO2mmRtLagIjA8G0E5YJ9bP471r3+HLuENEJbmEJrNwBRtF8Y
HdJDiVMmpE/r8SMxcCVKN0ajJOa69raV9zVX+zfXR1S5bieIRfIFa6kt0O042kI4
D7O9Ii5zsiGEOOp5BMA/nhSqQhkMgDy7XmAxSU49F6Sl9aLHziOVOlPDB2/uRFx0
3mOr77LOJFizUdneWN5Z1szw2mGeRyzHxtB80GAttre7znp2JZgPS/+rIo9xrw1e
V3J4+oTCUKGp81WN6FNmEKWA73LQNwUTNHLuL+X4gx/fFQHeFwO16QJCgj9FIIoH
AANrNtN4zBnlOvzpDnI5+9F6E+7wpUNegEXxgsg3Z9OnoHOWvo1A5JNn/OIT+a6p
5e5PAh4HBhfURMCegz78PJ65NAraNKYxWg380rNHdCITdCeLZZIhNNtdvpnuqsrH
yE38pel7ZYsW44LcZpoZ5eym9Fst6fCxxXsOD6i71RcG5163fPRs6502Dv+XcEc+
NvIhfo8xIsxh8iZEteOHuJVIoGlOAnAl4j+JN1fxUQH2JQXtqEhuyXr0F1Z8+qUG
2RBgXFSWfOH/L7kpeE3PwT/+5KjMOZjt6QDz/2U2tMR5bb/jIm+kJM3BIop6peEJ
Oy0JEflGyoN/kwxSSIAzymK/GnfAmj4GXKzduxblowXJf2aNzADgqH0X4H+SRW4t
YKXlX5fSiZ9xVCSIphEDu3bvKr6GZJmmDjKltuvRTxQJPlsIRz4MaNOT5PxQ9/oT
jBOBgV3voJvNlqK8ny5F+9JGUsDp8G/oq7UmczNZFAL8gXGDejvRuUHSYzaELe/N
A1T010ir1OP3aLMACv/vGNKGAlbUxcMWXqMJGIVkSQn72yOc8Knv9AKNGyPdYR2J
Ema1uez14U2z8z/YW6QgAtbyrAU5yemb5vMGyrI7oateFR9hRHNnPFb1+EQdqeoD
LfCbY4tnfpshCGULcW6z8kydQIODdgwYo8frrLnACG9XMc9w9AKr5JoJQejClOVU
+XQvrak7uYKlmvri3kEoT5GkB/54dlqwfnqH9+dxuNMQE1j5qGv+X25c5wkQAcxx
rKTTU2kqgqQp/n8T0I7TbFdRRQ5YQbvGW5vQAlKkWmTDvhYKWtA3hEkSMKnDi/7X
AkXIEPCq8v0ehmDOLbXbtNcK71ZF7NJ22DkNmSpOjN6YXl24xWunq4sSbH+qqJ42
uvZCAHy2Pf/zB03FGuZcPYN4JldXhy+KYFnk9R3ypsOXTke0PDUJavTfB8U4lEZl
eCn0lYswfW9IkG+4OTA0Z0Ca3kR6LWfcsvoYE7ZE2zmSAsGV8A6vUZsDJS+aqSYg
ZLYPSPhLaOU8Cz5QLPjxlXUB9b/Q1uSbSH9+fWDVgkE7wvCnwWv7+VQBkKzIG3pO
MGai1KbDYAarS9l7dyM65iM+f8kcO/yt0Gf8WmL7PbESrMfsV3OzsUeFbbFNTkNB
TMxmwnRmDfhOzT2wnJV7p6qN52UJxeuRzKA+IpFQF4NXNihAjOG9FFrlRi+X+a8M
6H2jbZAGzA6/U1dh6JN1sKx2FLcjCwxImXlf03b2y/ABI+50/nkkhS6gLddbcVCL
I2qZXigDhZdSYNO2/vpSYH2jRDwQWseMDpLs+UIoiL490YapiiiqctJlHeAZVVT1
vjb+7tOigGCep91WQA9bsaEd1xMzu10rLm4DXcL9r5Nt7s7rQYkw/fGzp3OdR+dy
vTIOgWsB6mgL6lH20JyprIpG5K3eDqc1nVEeiF2Bp6rcFA79FyN/Jxxf+E5N+rqc
2kwLaE7hChmElK5/Y/H3L4qckn+jw6jtTgABHEaEJ2tELVgSzXWv7PduPb3iPVKP
eTJU7tuPeikfHmg4rtBcLfNbFDxhzxy2o8ANCWsb8bjqUc7OucpabKw2DdoRP9gF
in0+KDAg6Kxr9ggENtO5IoQ8ByFRA2d72G8v4aQokJCGwvta0BAQK6IExYI+H6Go
Rh2Oy4m4TUQyqht51/xgwV9AHYQBnOLRa9jOPLc1KfPdESU+smsnWlPrjIB9D1nL
0DffaMNEulFqVbFtEqfCmNRVcUS9uaNu74XgVH+eBIGiUwtLDD149CyOcKw/sBlk
hpOqfwERfVdlz7zbP7FNpNv+/khv9ZysSjo8K2hnUf4st2gAcfuTi3KTjf45WdvX
B7gEKPtL8E8dSARqfFSMBukDo1NW/ajW30Tv9xzVoctz1olX1CbvyOIBvAXe5llY
EJlsWhz8baygnLl7707yCOnYhGvX6iDWE9PFfDiqVsSb4F6JLSXL97WbES6+6UXe
NiUWQjJorcQybFtUln9tKru3/PBLgCxXUPyelZZmb/1BcAFWDV9n6Kucg5IUHcGH
5No5a1lJsgYOBKI/SzoZcKE4CCEZrC0CaMdASjyCGBejDpyRZqzk7s2p55fHbQZw
khQ/wJ0TwRsH0mLTlhP0dIo33uTdUmUXoklry2ZMgmuHB/Ae80cOU2tqZ5t2LAjR
yVGQxVqipO0Pz/EBK+0yWr2ykL0L//U3kYjHuyT8+LC/LK9f514trf/ovRHlkMfa
jLGSsHNrXjouBZvbS95xRb5DdVsengeSuP9X/cJRqfRiUX9vtagpqlZJb7Qzizdk
+y/4w3zp6RMkiK/6grv814onWck0dhqSRc4EglV5Nx8CibXgS+E6Z55zFfCy5PUA
tfmQjjAbcc8L4j8b3Gw1HUzJeDg8hYQu1LFBwt4UrFczEtfTVnveqtoKXJAE+mIj
+h7B5AftfmU11J3S5Wz/P+H6Yu1BgOei9H9MXpvjFn6/qSYbpiiWFn+5AZAjEsFP
oGJW4cqGceXs6PLvAmQGu010RMqHBvkVfUWOcRcZXZpTW9mV4TotrYQkQwceWl+x
UvBadi4yUznPgv6jUnWbhEGONEsTaLiZqMXX4zD0IiZsUO2xDp4c/UiJCuN9A7sh
2CI2BZn86IPceLlQxkrNEzrgV+mygMo+nZIDWT3Dps7bbWUB22IlxvwVHgBSONe+
27vjQz4mmoIBFGVa7c9Te8GFrok6lHz6IoL4yYKD2dSccixTh4/6fo+XKl6eXDzD
YaVpM+tlj3+R2ftT9tV/sdzhZBU3Bz3tnm69un4u2srVmg+hm4amGy8STv9pc8Z2
ytVwdV76ETFxwjufckjNFfCMs3evDK1veFCMZPjNT+1acDoGL7c9asJ1XXLPL+61
GrVDXh8v1W1CMbkUYllqbffFSlLT4FZkcLHE+diMsV9w0Cl2QGnL6LQuo6QXG6+q
lNJJfQ77CycvANET/4Xk1vKwbgj1KVuF5p3KWlOvSgYRzQkcex4/qlXohsUQdqxF
5+mqWECQFKkS5tOj5gFRGT8VtELHCGGaHlssauiq0f5fb+xE0ItpchsOf980Nib2
nvYimV5vOjPGdGea6rhbmAw9UG9E2t16+MkdjD2lPG+ZA/bo4t5M+RG0SBuC8Xu+
EApny7LvDtxhPzQ7b5vRa0IAKgVL47SiaeibX1c5WKyqffM45Z8VzyjM6eb2zFK1
TbJhlu68j0zX+7Z1p7/Cz0+BEMGEsDKFJX5KYvByaxEmoVMe9mX5hTeqcwla6m5M
ZnHnc/sLTc9WnaGZ2rxxl4L9zXu0QvD33Ru1wWzDKSZ1rmjHvs57akIIRqYGAX90
V7sx3+gUss+Pn76CAbEehGIQhn2GrBvqsjdDSBAIS+PkjBKEQNatIqIxtnhFd9rL
IqM7zy8TSecnxUrG2pirbrkGu1epw6HJl2Atrspg0TeA5/+W3YSmJ6SJajL6mCbb
4JXHdr9b4YQynso5JCyqzJo8gnSFeTIlYhft/It/jmtKPOkv/qsNa1PxPW/wr20O
pGbvZSRK4+rXHB0IcWnuIPl450o15+8okrY57LxiM+ATrZEfFRYgr72Zn9KIPOlo
yMDe6KrAgq7KANfZ+2Rrz5E6w8wxzMeuPRo7ZbLBiKXHQRhetEB4spl9sSry8Jem
nm5HGuXKpcQR1AhPgCm/woSnUWnv+9V/bzDoUfJdxpUYxPGFnCbjNGaoFFkSntl5
1v9QPpgH+HrurCTTrnwzFCkEzwwTjeQZFzIWaB/foPIEtQVru0YkftfSAu5UDNc+
4yD8Dm6Jn72TUlGiClizfxR8Z0c1q+rQXVoA7w9LwpF2SkDqoI2uukI0ypmx3Oyz
ShXEpxjYJewxxRDgio9e6wiWJfV2he9ssoDkxtMx6DmAnP283G1tEx/HlcxUFxKL
RsvnH08MK4HIjNKFIKxmFtMKeBCZXLO8Lg5wyoD7Lkz4OSrZFOT84JyuPRZ+mEGp
gQ3295lqiw3lodt2srfHaOQbHqzXYS/RszPIM+5dFAFsNcYogTFH6qfbXpMusklC
/ziHXFVFG1icFBF2LFAp85LT/5D1lMB/Vp3MvJPSJ8uXcHhv4+z371h0X+isY100
Dwz1LZ84rb4/ApECucdZ3r1LIrXZbcUOk956t3t/qv9/CKAsJg7C7yg0fCpEWvtz
q2qXdIcihcf2BELKZ1LQimY6lm3ra/cjc5fwMSblfaJoDBnZilob/BeXUUiOVDZn
Eiat90GSBU/wdsBnQ9LkLiDVU9FYAP85YUXL8gL65G+V86NSsvjE7H1TyHJ100eJ
TFcVFzDegKdG8F0X19/O8BT4o1EAQkAvYmsgvburK55J6ZZN+gr+Pnk+PZzbDM7C
qMJXHODTaVnXC0HaKgwzji/9ggtthWlVrFoKD4ugogiRvjXc6gpfKgff+0Mg01II
CAkvq7rRVoh1pRK5XSkJUCXzRQaRBMf1meBUdFb6jswqVFcSG371Mx5hJpvH3KRT
x1jMZgYWVF89WGWqjHHXGQpR+dVudqQJ22tDCL2cPubp7hhdWGxNOfQclX2xSl0l
XYcG3HLPPj3vFsDnjua5hsG4hxYuCldLweD7GaNJ7ccjOhM4clONq5NpUX8mulrt
1Zkh142p8GJvqgv9xxoPj9kR9RwEyq3cGBYPOWKBAXKFsr9aLYHOyYEf5JiuRLJi
aUGtiaQGPHMpoPhqCzgfGRf+Bf/b2RrJIFl9WFLlr2f8INCv3RO5VvAB4eDirLA8
hpW/ARsoJh5Kjcg3zuuW71zn2xt9Qt67+Qu67aDWWq2Q7d10h82Be+/EUAJB0uhc
aPaPBJa0PunmALFsfdXQugxP4MO0Y+meDGUeGlGjhOCKxiYJHfMvWMctVVLaGOCM
ibtHM4pqMpGGUapG2XboBPPmidDsXjge4tshqov3hLm5uHzYle6pO1JsFVcPoaVk
Y9kB1wEjEQ1dcNVGt/LozSnXb01NR3JfpXDFxbzd55qayKZ3XVHnR5S1rC9v9PtI
pQ5bcp6sshYjEiXO9ON28bXom7Z+14vxE0QRdGJ2g2Py6F9fLOjj6d8JIF4bb+Ix
wYN+Y/RDnBzl4bpaouhizlLTqZd4SZtzHKNAp5vjaH7/+GSuJLSiW2Oep1shr19a
hsqG4HLHUW1urSKXie/gwPOsl+uGTBQ2hAlqsugIjbsO3gQYXe2UhHfkXubytDeI
v54DNwjgzv7EQyKv5nJqa2qmtf24Xx/ii8Ysrt77NplanUkQtfNCPkk1SVKcVa9n
6v9Hjv5dcll0gI2ODZ9nyeUPyzGCwEz6tJjHf07+QvOp9a8y5//OeRy5o/KQpehF
xchI+iWI8S6mxardrMKuARVdMBWQYyM27o+Pcm+Zus8S3W4CsMdF/g1MnYWaWB/v
bYoONWF2JAOKAYZJzwBeMx8dk5MRsSbhI7wIIDyInETg/oqZ32UBa0pSUVWuD/72
XuOwdOuhM592f/2Y7qFgRwCcMDCjoLxhEy2SQngEqO0PcB5YMcdPAhF+E7V6EKIu
/hXvlcptC6hUu3Xks/WD5mujX/4shi9qCSA6f1WdP8wj9AGk5HN9UGX74G7s5eSP
k201fJWJhzhpc2ITXFemr7x8fxDEqON2g4fsT3YH0IumazaUveJXcDy2t0FcW5hl
BQzh8kXIeASZmGXtBnu5PulPA4CNO868lnE9xV2TfdWlh9PtltJzahsBJ0+9xcB/
+L20IhWdmiOTpA7I31+45iaWbYLZzkS/ikDny+eqqjQQKrp6mCVFy+NikgdqCJ9n
kFMHFrFJPAHzy6FJZ54MbkxwSGn5g7Lgqz22DEcnLY+5Ea72NTE83ujjEiQ1s3nV
vLg4X1kWEPP3vne80zVZpMr6J2JtcHzqn5XbG95A2XmZZ1fGTxjCoxtrHaGtE04S
LicYmv8x00Aqg5opIhlr2s1T+p2e+aLlafsKASUVUBQpRag2zu7BYK5GR5Dbcv+p
AsGiGAKY6ULq0Q1coWXJr0TpIZKTt+LeraQ1IDD+ijXd70+/pYjQJ7U5p/RL6BpO
131ZZm5Z3516L59geeeNWTlx3dbdJIGsvBmK2gVBH6WTOtZKvOZ72FXJ4Psujhge
w8TfCV6qJo7Fqmzkg5zoDUqBchW6mt1NGakbXvRB6K0x0FF+ij+3JaCm8QnRvNia
+w9ev9NeCL63JDDOng+/gNCxUJCq8dWNduQkbKeQimLbMJgnbomeuXWQJpcJeZEF
/gTeqVT0Gd7GH5Ej/1AzT4lENlr3xHfAMdjo7yaoKJAi8funt4Z2NZpFC96SVfs/
yWEYEjQPrUc3ZObxuCAedcC8D20NWX8DE0EKPukRcDteqJ1PNaUNP68RzjCD9nLL
lO5FQd98C5WU4fdxc7PNuBVXOelqfgocrmGRKPdoEUQFhCMvEHM4zsFSwB1a5m0W
cNwaye+E8jdQiNrDX2C51gGmQ1AM8gkPxgAe4bO+dgUpIXkWn8a1tZQZ12e2dGz8
gujbEIH3/K+i/s6SBeug062aa80BuG6ZEYwZwN/KvNwyj8mLtLaft90aWSTzzmcl
hj/YaPdEAAgjxi4dATThYgyGKiUFNeVs+jhbgAB0bSMw2axqYPjnoSI1FeUfJDFj
JjzLY2nhei+MH4G14YY6Yx0hrwWHhtwdk2RPyY7bIoaY3mMtnVn+T5gPed7J1a1L
wEs9nht4AAnMt81MMfSD2yO8m8u0gp98BHdSXrL8oy5PZdx7gJOvWCg21f02tMWC
faHFmcJd2YQWrYK2WACs2M8g5iGnSjJOucc43sn/CoyagNuxdV4QYyN7Sf6DC8t1
JaWmXvh9A0IHLhunS8C0SJj+b+t02Nw5ZVlQ5SDXN017S8mP4B9coXxcX/WZ22Fc
dg3lIFTbMF9VI+dr5OqoVV5Frf6L1U10TzSCfBwZz5Uko8vyxyAyqRisUyGzDVga
0li4HDo3gjz3OOfFK6tptBki8IOBTRxumnIKty2vKUvGA7VmtPFZLf8acvwXMKlH
B3wWCyutfO2wHp/WksdQgSUcOtSVFkJxgRFyGBykQQKgq4gQP4iaedrszNXnEhAy
IqQKnVrHROcpqG+Rc4LTvWUjxByH1MkPmk8FFIa9WQG7cPv6V1jdOjEYtHVigTMF
/aDn1Tj0Yzjw9ytQI5Rf4+ansZg6f48n+KOqr6HJRGjgtmL05Gf665QmGvvww7pf
3t99zJyJe+o3SmnacVX0fFuWrS93pBKJU2AwdZTSKGkvHVl+nUIEEIXKLUMWpV+r
LDMWzv4TuvKmP9rvnoQGMszogMDAMYPBxm82YPV9fGmHB4VmnAFYvE6J6yJq03ld
R2BTXl/17SZ1ZmQnTJ9KGvKABAfa0iPV3B8Qi8G3m4d2uJs+wmMELv1Pms0c9cDS
xe9/x/m/qc13D6c8nIbNB6HehMTsGXW7KJ24Pu+mufELEI3OBrt237TpDqttgRML
0U9wsYOLCG/8IdJCR6luqFUukrpILRvRwcmJ3DDt79iV5PtKIlf0fHuLD9YPe0eC
gjKDJHxDEUbttFPnG3DOfU6Y+LmzX2K8d2Wv00eHvip/1Hsnk/wDb275ljukyEHF
7WRMuIvTymQUjDCgL7TT/PKiT0K4bT/S2SMYZ4B1OsTqO6QlG/JzNNumBdPJQXTW
VPun9T3YrUCijkv0Uf2N7dkUQejDqSV/JO+qpFhBqBcEw6/Ty8hKYoMpyD5K419V
6IKYXAJB+SLaf5Q9jBeqnWjrtdAkKu6CEglTQkbhV2wmm7TwgpWP6qWbdO45ySE3
v5ulmP5r8kvZDOC0cqnhQQ6dRET9IRy+Pq3Z3KGqRiGTfF9wmWerxpWOiMHdD0n1
Lr8XMvND36hck53Frgj1rOkCmAXJHnccrtYQwipyhCu9Oj8YWHNMc90Rd66lvwHO
nkQ0QkEb1uSB0SrqzCCdq1ESMUW/+8VKyjsj0RZwPb5bQj3ol3yYe6WsimmHz2ES
8KyWaK6yc7w2/hY5/RXrdOKu/1RqIela+gA/bNt3kctKD63Gki6lSDqohMLSjmIO
jegHCjYSR0BpIbKFuVlGXU27ER7xlAGA9vwmQgWckk9YPJAtdTY5UZznUrdCILdk
B8TM2n784UU3TCtRfVDfayF6peJxeJ7rsiRF3WapM8ipjwR6I2La2LaHvoNXeqjc
Q2QbCqbJ35PbHuoVEIvHbh6ZVraFI6Uk1wX2/6moWO9khtRtBmKCD6JK2rVjXAKT
rmvXmgLMaxATGo1hL13Z+QUnEiWvDbJpda0DXoHqgy9JkHCnwrXA3DJ9PqDQyGoh
H19VkT716nho25QJNaG//5yxq48d/sx9yCdE5WwVXz0cDq4AQucInln/YkybD16E
0kbuAUc7wHM7KlpMpeQtyVBRs++fscV8lUjXbjAMXhxzGibNLtVdk+Q7aLrm9Bt+
GfINe1JPqRJSDxjgJupqLt5pump2OL8ClpkDx6X0sQ6mOUGvd3ZlW+hvCSQEfpxs
kOWc46H3fj0sJiHVOEN7XzU4Jc6tZFsHzeLBtpBTQJ4krTkG/ZgxDNn9kRXZ4BgP
wDN//m3LNvCCEGvU4NglRsdVotCAFN3vsFtuyCW3pYsMlKpxvzbxeJZr3F7gEp5D
6i4BUTulNigsF06cMu9jCoa/sYdt+Sgyx1YdidK3ytBgazTasnM85gqvKa8aNemH
eLqhIzb+5fc7P9DW1WTjN6C88imcdcQYVPgEqzQXvDz+Y+HNah9MPxrHkPYYZMTc
00Tp73VIhEXGemxyN/CoW6//Jw8kjTLVQa3JIB4HEHPdpXYpDc1jx3s0uPBmWMAH
j/pUCCIhJ7J/opUjQ9y2QlleTmG74QfW4pFVo4rWEO1WFBMEm/YoGsAAOyknPNMV
nKgv9Aga5cJcvbU16D6H3572SLIyHKln7INF52nAfiui0WwGB+WaPOlyG+64RrTe
N3lGwxtpgNtJuLt/s1oWQCRLEj7SRuBskLN1k6eOovTgFGBf7Dq3Iy9xPQRoq1FE
f+pjdEb4NyTUsrTDOkzlVqmQogtjkwPyuGVaGGK2d5dS4E64iN8dhZf4K2bs5dyZ
i1sIyVoQE9gV5dNMccREcKdbKom8JhsYMuCJxUjZ9SFUJCexTYg+fBxI6sptvSdB
g/+wPRj3gwRDCcqUDeuFRHuNf3xMyonfon5jUNTDrD/qU2tGPDXFoWuoLyjeTW5R
2zkh+ugRoQCqKudh2c++PFxrjiHvqBzJX61mPpNfWNUNIdECklLU/kAtaIp/lX6z
eU35mlAu5Y/awpJch4AD6hRtOhfcGDzYPGhAFzpUhuAwN7TsEFK4n3poo+sezFTc
s4MHXxfMHKv8bHHZ2wGn+UoAJV618vWroClzK5GXAlv7ywDXgctGGjN/GyXPzFkz
GhIWJVYV+nThkqkW6aTVQn1/DrMtL7fp1GPdubbTq/emUfS9O+Uyi/zBDveNEXU9
XjJR5T+upx6uSMHJsastkbf4VXvJBNuXJraO/LngLrBCKa160KBB8b7aao7CPPnk
PbmRc1uOTd4rcJUJTU4wDqwGqvkg+6e+a5AHvMx+iTcjkxlHQVdEPLxQtLGY/C8r
F7GNYLjXi82pqYm38JqcUDiWpUaIfzvrd+OEg19/Kpuun/Z4FDQe5WQv9RvXbVON
jRKYtOVyHlwmYMwnmOpI4WoXN3SSuVxG3jzgQYRk2QsBQbDzF9uHwek2Vd2+Pk6K
OThiWhOWqUZNfaNauOeZ4ReCR9Zwnelb6ETOIYY+FSwW9u8TrJj4IzjXU0luWIEC
WqtKFefA9HxZLpi1lWmurHynhupvU71L7u7I4riDpeonOIwzwib9hMJu6movXMnI
3X029vT92J0i2S8HorAH44Yf+o/kQDEp4mo/nZN4H+28LE9CSDTaft7tLqK0MjtQ
hfNnB3ff02v2wcLkXNBIxYcIBoDZotPH0s9/Gm7yQjVAvuKeRJpjSbTqca+9st2Y
S+phh0a2ihb7xq4sSjdrrTSE0e6fw4INzZZIoFLT0UdOqegNS7jOsE1rg3VzKD3J
cJeHvAYkIw89hMIAMOOVnkJcxNdD11WVdheSenLxKjsAKZT2arahNY11TaA7/Xu9
dPlxIYYMKkaQXJn2Az/E2uanFq6YU6tBQ/BuS2PluAbRAnnVaXP0l6K5+zFF6OTl
+UxH0ezqSVd4Ev5A7sNxakhEwoWziVAI0TC3aZDl9DyRzpebF5PoKCq4xNuiedcv
kb4It+jwg+KOi2gAqmnAEzXrhpsHYVAoGsxbzNo9WyMOBLenBnNwe/cttTS6/sZ2
sBvCHww3VYod8ccWKqkVpRv1tAQwCOhYlK1QTFGkiuVIKr8PeX4uuuII1mNZGv0i
NAF+tjFTUFWNvbA/8XhNN5OsFL7z4yIkGJmdUfSVLVHvLbqD8Yp72YkTYXSwHXVs
K+W1oyRwz5NfYKsIyTMyPIxCUmG+P3pdnjkdi1FUkpTplHh6JHXsRc3s3S9xyP3v
ofxDvfRTeaqAd5RmQb8PQn8WFovwY8QxRgduwD0TGR62a7iKpGdnsYOkHQ81ilx8
RZXfwZqxPNUGGmQPSz7e0bMMnQS5HHl2x4VlO7r+FfKsSVBX6AsO5odoO4OE4T5z
tmQ5Cc9k+ylmJOwhVWlfOfclRMAo76yBhVA3JtBSzK8FjT2wg44zoOcynAmXyN78
86+4AVeSJ3/caJjv3v+aJkRpR85l+izROrOqC9qF03bkOJEEJyNG1Ctby6N5/4zX
DX1B3pGAwjszEQtu1UdGgJxkjxGHpMcEYR3A47tJHszBP5gcVpZJelu3sb7nGK4x
UFPNq4eFyyxSq9shGb4V16jtg6Kta3nlZtEN7kfHVzBfi4WTSxXpWY6kanEYFtmc
L/2ujIyZNFTpYRRhjMn626Tc+vjcBMgo3ruTEVfN1H6hQN0oipBnRYDrBGrMHI3Y
s7FplLWY8pt9TMQ/35dWbhFqP4trQMRZBJsTL6F+DF42h1sOGPK9zROcNGm7d6ZR
i6yfS51aSSDqmbJ2xfceeVB35VpxSkrOQETUGJ7Cx1/ltkrwpeUGh6AfKeUW/EyB
/TVdHXaP7gU+ZVnZ8rxaMVvVSlBlPBqMQWbIeW73g3FCNX5KKK6dUAEH19Wlw6oP
x4i/AEl6/ZUR/AzA6iCc9myAnCzkGHLq5v/llTSzDBYrMUyfDnTaJS+Ix4sNBstQ
RlKPLMwmxyk43y+CP4gMG5A5e09tdtAxDTpSWNT0cknHSQOZ6X7wg1iAvEa3DSNs
3w3DFtrcCxCexDhQc4I49aeTpQTexTEeBO30AfqczLcOpHsLMkly5CuibatJY7zJ
ekRLYfkICxD18rqfLaQLo64sTj/55ITQkAUkaFBWDRM9zUIIrXAPsvl+WpFS8AXJ
RXdB0VvSqQI/5ylmMvWnAz9dnZv0l8WAc+/H3q05yCvdF5/m3BE40vhI4aCgTFJf
i1dSllpNWvAXrIqmQbW5mFm+kUpu/4aDFgVUgUqhMUXdOovOsiziYds/qKhAYUTm
XomTliHSl8OG2YCkE+dQR2D2bq9VOaZV9RKNDrfgtP5C8KRrwHXkSYN++zD4c5ep
GpA973ljLYohSV8gSsUpLVGSfU6pP5bVJnlFaGITkn5JwxFHuVI/LFF0HPLm8uRi
LjOnztxr+1J++ovBDNnyLQ/sCR2XllKLytkdVovztc/TSrwOd7Cmiteyskuj5Q1n
bWvVidmIoG+ZkxSGdjojj7WqFNfsVITmz9duBXaFlyY/OyF+lnr4t97C2pgyQ/+L
z5q5wfA0OS2qSksKSgeUnOC+g4Lwn0gglWFLouvT0/IYYfJb1Bydq4Qm+Aai1igT
nBVQxJjzHaDado7YOSgLr0f9J9lFphTJEZl8tNr+ZzIIHBYYysaIjVlBQDWt0gXe
HIrw48pVlx/4g2g0rEmbAaGCe3gvh6URizJ+7LCsJv2pmlmhhJd7Qb2qEghOxyXc
S5PZUsvnWhYb/LksKEstq38fVpHQTXHFHMVg1u7cVGykEVSvJdVhl1MeE5LDU8ZP
IiJ5PxiKGBrinc6S5CzHSS7DuHfr5WacEpX2Vx+pzkI6gjY0+s0lTIXFF7vmHb9D
F6zNAqRdU6rJs27mPMn+TtVekQ930jMCZCPGQWvfr3T6rA7+qhwhYFZhIwFnxW3j
Wpl01q/vOlUaTbqnKvBIa7zATt1pehbNWGsHrCVUSNtFtIeqNt//l/nMY0Jos3wy
TDqEXTPmZ4oK8dt9mPJ4r8Xi9tyjdhBMFAgA1n3uKODccSgl/cuA0RS/7aujmg/s
YEvF5PuTj17bMbvdnl6Y1OZmpuX+qtvvFTdOUvyjuT+1E4qm5kWwDTgirTvAxJXc
0Ho9B4AKWLD+a5MdSM3p8YH9HQz//qq9ME40cXbpx2cthcSSUeNPoE43WX4hD8z8
Qn/l+zA2szPxrnzuAh89oH60gB0xkp3nq5bo/ExoO9Xqn9wB3W36/TKsKs3zC/Jm
kvSm1fAuazt5Mcolp0XD3bANDXjImUjJF5Q5a9P9NvOKts0cyHATG2vRIkSlPdZR
7xAdn7/pmDgMzsX98bwElz+vstrFYEWis/Pym9yZULqD6sya0hdjkAK9m5/CTDKY
A/Ox4yem6Vo5H2+TvnFxYyD62DkbGn3Z5K4GrpBXGLK4V0j/vxJdezbAyWWzxb5m
uJv8PMT2I/OUYdkLgCP2mcle15EMGYZMnz43haasQOsH07Y8xxpkYiNxuaRI3Vrj
ls4oVmjlxmauPhbY33jHesJG2D+jtb6mMoyDDpPfuXRVaT4ax+Ox1ANyDkBODJ1Q
zcaGK5JTHBumksN1ClhxU5LCKNXQBDFJ9nG/UdBFoDPoGinJPMXMtc9gW3O6rb6k
VIUCMXFIN6Q02ivqGcNQVeiYJsPi6MOgeDZs9DS0C9TAYWIGfD4VoXB+UWUIxLXZ
/iAqxcd0PGxzAcPFPI92wNV7xAbkPtL37re02TdsZpLSg1W0EvxuBJKEkNEri4gE
CctajoU52JzsI0jHlBx8nvc1VMCwtNeayUl6tfBszMhjFqgkabu6rYFq79OzyehD
jOB03YqrGI1pxEt22oWLFuDvpcrRmGrrV9kn5fMOaZwlYPfQqYMJnW7ydkQe8JtD
Cct1HGycN2kiZuY5lNzm/VwpUKjXB/17UBxnaQSGuKG2cPYRwCo02hFP+kqg6vMD
9PrfvVanHqqf2t5ZzFjuJI/1i3RpBYLlowhGy8gzP5ESyAo1b8OVA0leFEKUGcZO
nYpxRGS7Lnf8vjD2fPtoPD3aX2l1ajdWOhX5QHdS5blWY+2OPuFkSoEVB2wPnIyI
qMOCIDUgcOinMbaHtWchSOtIfaM2MVRxs1rbyVbS9nVW/uLXGS2dRkaK6nZyXSzr
SVPvXdaDxcopNYNZ8Z9eQxNMpMBOkEAPWftgHIS3hPuCboALMyG0DTpE6sLiX8vs
agYQEsdBeCwrrwJDlHL+dQdHxLtvQxrj6pzYd4Vcw5c4JHMEjf5XRXqqA2XKVZYC
2/prF4gWZMeQ16FsSJVw/rNj0llzRMu41R40XFYqCUTaqOGTs4HzCKr+SSpAJLSx
LbfwVZlESNIUpVdNeLNMzoWtlK7ffM9Z8JlWXLMvg5phFxbBjXsUZlyaJpo057Px
onzrAT2ytO6uu8Z0TKAohCWTJBxTU03MAi3GU6Fcn7Hf+VKGrD5BO/509Nk8LwNj
ldd5YM2qO0YEkNIvO+EpOatHKiRJcvNcgi54fsYDvGnSBuP3xGfBC3m6OhUFFVvU
LiwyPu+phLN8rChekiB95wqyPQ6zoOC2evTFflfQkBex0gd+E0qM8mqSQuZxFxw6
2VbYlWvMlgYeFD2GbANZCu/f3+tzzjKPfErhOtw3c6ms1hqnkfHAeAk1IAeeL7b1
ZLjCJxjnNjpUawOfJrpbiNUATfAHnawr7yDO0BwID1rSvvYu0LnUUBIWXm/+tfY5
nLHcHh/eBlB5xmEfBPzE0rbGIQa9RDfVZJezyL/v78HEitq+m7TsaOKxPJPxH/sQ
hqzat7PkuyWXsx8lK7Y8UgGcKtHHfqDq2EPIsUIn4GO9MQj4tppFMoE2+d3xBgr0
6EPlvUziWf/zaP5dU7DBaNNBf6LnbwK62ubf16yfA6hrwGi4SM/qFvwoJ5ZRClJt
2fqKH/ngTDNwjZtQTzcxIouLgrQEcY2N0G8UdLVCWEO7c9a7UjIUOnzZYtk3LP+0
237h227OM4UgrKLBQkC4QkDmglKv4K12cJK9RY9ameEc8I39OXcNnUmPJEJL2ds4
C00B9XFaNmE/ndL8LTq+S+4l5a6wCCzCnJ5l55nJarmzH0TTqhrhPm3/DQLIbkbT
LSC/2gURf+JgLMBAVuumEZZ7wt4H8i/z/u7hFa76FAXief47s/Fyd0ZcUX0izvTP
ohke5XBNYrI+SIzMiqtwYXXEZnDpDUg5yowHxsaLBfWp3z0y+hdilG59p7opEkiA
HeWY+vbsjr45J7oSwagUEPgfGnqBqYJbos17h/nfsyYVNYc0Qde0gu+6Hs7Mv9Pp
cvS50OhC1vbzUTP6zbEBXj7YgNKMXL6u5YRRct5cewom0vBltn64YuiDGzqBWxY1
uScEYt2SUZb41ZsmSV2nQqIoa7YxcotssfUaULcm1s6LJJT0SmxEWsH+R+hNTPkl
78eQ6f21dIp4thSu+93+8ar7FJ9n+vkNkOb/P+lHAEoLinytTox2yQ+t5Fd+0ewL
L15Ze2dglNyq6pnYY04FJ4VGK/yhWy158Yklishz3BXCBxrQ6sn34IH9ucYQhj5d
ywP2wj73RdjC2KYudYbL9TYUWJ65wLEn4jWJyCdmfe/ITr9/l/NXnZ7sm505/J4W
gxkogUP5/b0y28Lmd0FRZXosFtj27JWGhYAQrW03D2RQD7Mu2ZTL1wDq/Nz+otvu
qM4PPbhrzVjMuKq07OpedxUiMvuJ36pp1AwS11A1ldt2iuPDWvdg4L4LdmjQMwmA
7jYPEUzNrb6xFPHmGXfr7TNVBbZlmkVw1tt++cx2lTGYkE/R2nqjj/97iCV3eg1A
qmPLOuIaURPKIx4SjWaQqgy7iFAMdHkHoyaOdfwUJ622yLMy4uiYFIUu1skhjkRw
YBF5QP5m95cb3bLz5KpCse0s+WkxHNWgDwsXPNFmVwBV9uR9p/3TOcH3Rhd9d29F
uNw19moNbxCv5TPp0gweak+GuGG2bQs6yF6EQAgGYFTfLLT5vHG/lJ1RVQz4y5Aq
/0frSyl0UAZGAts2IRpGGOOIBjDouHgYhtZIVH7sQH3CqyLQA5VE+DAa3cg5ziAO
MM7YgNwhnqNjJygfGuRe5xpTS2pzcA5xQewuqsBBumhNOggaq9gatBOJGGVieUrI
R2jAEuc/F1lcDKH8hobKbngVPIZNiZSkfmlP4YkXOErhaxakNLww015/tgEYc+vm
ZLl3wGHWhUmC0rm+yPJ1spgW2jIGmUaHinN/AprRLot2jPdOt6/CktV/qadXYq24
841ao6uDA3RyDUUP+umC6WH213D1offoOIRIhKUjRDGobp6CBccKvwWUu3rky8dF
8zPmwR/PPGM1/4U3vISuU7twptXOSE04Ql/+q+RWEEKVNvwCTVWTv0YY+voFoPrz
es+p+YrUeWts304tWJjADpAJQl7o/QseAatRRsTn4gDcJPYA0jOnYLGWTfiHdmy3
d1FG3znZ/1Q/sqUT+coiFWAXo8PhrFtFw8XN+Rex2sHRxPXtnsc7GUQcmBwUCBCC
o84FQjTOo7lW7AlpJma7cbjQiwdN4gkOhB/9nhDVmv+NJ0jtmDvikrAffVPpt6NE
ji+eVjJAR65H2sdYLswdbHdE4h3oJw9HzIDeMMq7DCc+WYaq0SzPm8LdaBimmffm
qX82mlg78aUWWTzkdfAaTdqGVmhqO6nxhG8QkHlQOysHwTsq4anRRNOeHBE1xssY
WIXHJSXaHKRMuIf+Yq9e+JlKw+DBugGT6h1dOWgK9J6oapyw1BThokARLcXGih6n
101DGsczW0p7zapEvWxYZrMz6TLRyS3I7FHFJRW2G+ZVEkWHcoE55YE1Qw46/AsY
fZcvzv7Ba+XDn8rXD7X3B550rX77/aHuHN0Pyw2KqIZJa5Av21xPSSafKAFCdqmY
f/WEyKsZxHXx/GFkFSjKav3oXdAMRIPdpjiA5bhZIvD1lgytuNvWPquM58bmSnAB
MW3BPGFzbIoWVCwRvf1MloFfpC53oH1CE56iwQEFHWl1wlkhQERu77HPShj5ITf8
nQu2+aJOirv7JmVMNC9Z++h4sunxhiNlBPa2B8H7BV6C9ODtc8JfPF0JU1XDZt49
RQEWPkakYk7PnMArdihWZlXT5JApxcZ9VJpF2gkhdtSr/QbyDkhs8yDQlKL/cZfo
uXIFBG3HF7EhJIFOZErIY8WYFodDE/RSFS1jLGKlkzlaaQxSHeMYl8TW1nsI5rfs
3ow0GVXJyhHOqt12kVBv6lBTCSGnLQ8BETZu/eZ5t7jRoahin4z2nViHjtNMMCuS
d2EkRUF3YVRLjoVwsQHpRMDkXDrtsS+Ax29kK6gAxlQpiWuY3vuKDYQunVxVKV3m
z108ETiYwLbqPmSQl5FtQraMeIkKMg1P1B6NnKp6UQpdIbfPIcLDvGyHe32PhfJf
WsUJE7qrNCsN90noHg/rI6IR5EQEKk2vw9LS1lmJJYxRkgRFu54H8CkafIGB5YXK
11GbbO4W+0i4AL41qFzZA8t3pDgx6VOIXHiLxyun7S+sIBIywmW5hMB2/oxvjx1N
oxqL/AsCTOPezF+/z77/4/A/QgP1A+3V/6Ru2RJLUPJs5OCocTSzLy4Ni2iahsHv
k4pJBV7+8UsZKz532tFzhzG2PJuOgYu20IxBkA9y2TfAStU31y3bcSkV9Kq9hahO
DbcHlNtATxz3GG3gUBeOsnu6pCO9/c0xEmoqCvopn1LWNM+8jO6bRCUfEalSYGRE
6tsv4EtFxJ8agIjwq2nelgzVMF3JCGPxNYXJCjrpBFDxqhWgXd13A1XqYZXd0X/R
RK/R4pusz4JvK5VR7kc7Gw2PdGmCthdx6zYOfgPeKQ6s1DAf3ePdN2XDPiPMC2Qw
9EYIYu7axwAWaClJ2fCW54hhDsPW0rmw5saTdWC6w4emMjXIrghfR4VthEB4ibVl
25EFpzOHQwiYvPNGmqHueWMuVPUML60BETUbVaNMtbFxTDepnQXkAiehBPYojuOB
1P5hzUd4XkkiFCSyRj9dtKASiV+YnmfiOUhsasL2chVgHT4cFuf7R009cPc/DxDJ
IUGiqHmlKrtjuDKXQhdgXe15a0theS7oMSqRtmMB2iqr8dH1NVCAZxVdJAPCmMoU
CMUmm3vY8cPD3nbwJ00CbI6u1xXmUSTCGOWFixWqdX6U2BSmctlJDBWDjY9gqRI3
WYU7DSGMeiRcBB3M5YbsWJHeDl8MPPulvDBziLNDPsOrsttJtQts72FJdP3hQfA9
r5eND5j8v2p0WuYtrwZlHTaPIBJPAGHdCaZmojSH8RA+dmHYJF2OKaqr3LQOVvaT
nL80J9G218BXjLeanVPPpiiuLHPef1syz3w6CJZqAXUwM14gvFElNqAynp3a+Zuk
GOr9kB5wMJZD4dfTnohw8ZZjkOsO7jS0Z65vPE9U6ZxqEKeZyPiNWMjY1OvuDEWL
Uc4kL9SoWh0XiaC23vRFtMqw9VVSAMstEzfGUQt6nzUT+DByFEqXSAidp2LefX7K
zhnLsIBnT8kXj8QDAX+XnB14o4qLSrLevmsdCjSwVse48dHv7qIxQRAcsRNfA8b1
ClCO3RsbJgxbveFswdvqg/6ebOPMJKhkOtZVn+O2tE9DZFZYsu1HqzYhWLRBSYFc
nvWfTast4PaqxgVtLTV4zg1T0VyZc7ZDSMKA8gfw5+jOVBoYXpwHtMyYlRGH+WQx
Wm2o8KZkMfBi9dcaaRsRSi0KgRq56WmE5PMktHI3LJJ1DRxh8zVW133oGgmvHH6G
0Uw71Ip9vhlKGGcO0uniUByXKvWM7AQzpUJbe4rMTpKf2WYNeGXC/E7xwK5WUzxR
B04UnzxLmAhVr2Gua1S0lzZZPc9hqr1QZ//Clqcc+q5iSHhCc+0hgYM/a2YfV39y
l9RSetbSNAsgeydd3E+5oT05HwKigD4aX5g7cqLcopQxrQKGdyvs2uddZNezTryT
DrUXO1OvYtW9IwM5XV5koQbZ4Vd4Id1gbS+b15KoMcUt8dE7tJOaLAhKHE0CwdpN
nSpmAGQ1CfdN+cNMaqjuIVVWooM/QKc5yGHtGwUAmXkWHs7q4yrs8Y6ilC68Z88p
V2T8+nQMBlNQGlJBFh/9lNRG7D2f8wE2R9zfMKXNp4dmoUPKqK6zGVskohiMR/bN
Oz41AEGzLZRsqYqPEjvM/wlNfjPTEyIV4GxOqrxgRYY+5qMHbFgwABTW4Z02xzfe
bDRG/xi55QggJPXxOk2A+vlTakIE2pwYWHU904I91eFGlqpyuQSE8KpaASbvs4Lq
ndglNm7I5Sdm3It5xiiZxa+WPab+OcUNzX+PLtG9MsGZ/oN/VZCB0AEu+R77WKEF
EwDtQvLe8wqphiVcRLV+Ld1a1tl/r1qMW0E8JyQrlwXMYEG/17E9gsV2Ld/BFylv
iZBC5T6KwTea2G4zIhh6BrH5NCXlx3fL/GHi2ipWJ0AoVLhvw/Fj/+zQgNM6tnOS
65FH9UqNAZFVyF1PAytSvOqBWxAjtHne4u7Oc0iZMFA/qHSxj6dvmeuIxrRIlOvi
AF8vDIdKURWCo7+uQzCo2muBHBDdA1kG1WAr2HanB9FDk73nC7bgtjeIPAfN8/Zp
MhTppAnzCQIp188s66si5kLQGJbNRzawf3CQTj01jPJqchtOXPX+6eYmgg7KD0VF
qr+qbM+XGcxH1WUKbA1gmsrnv9dXuWeRzqTI+cnZbpshxkG4OaM26X4zEL6UfSLq
hBpuY+g/6Ftj5cDgHCtD5/q1Z3kwCHBo3LK54h/h2WbI4Qf/qQKGcK1jobOwZcrg
K1kYoh37NWkAI47ODT88zBp4iujZ+jV00ZG2nNi1hkXpYK1WnAu44v9w5PtoMVCZ
HcU60DREBTyO6Ya153LGfm2YBGJRso94cxeDX0OORB/O1cVwjWmp7+NYzPBktjIQ
uR/75rTguHxS7ZkYrwZ2bCduznTbTylKw97VJInWORuxz9IGBwxGyMYaY+9gswvq
Qy8Uqgm31xwOvNwdNK/vlAktSgcLxFMRjluZ8AonWV6+eaUdbAbBzvM/WdUw7K6S
jc+71Cj7yxLtpDAEZm5tO8dlJp8EJwO6TDfJIeAzrRWNm3I891yj0ttzB0iTjSIs
zIi1W1857z1QH12NkafnSmA31WGZBvdXXoXPB32EkMheEB+6/kpHzDL5yBUYM7r+
UiezXiUaUQ4+pFlUQty6Lx4Mr8ddfPh3dVSnU4acEs5YD9OcObeOEz028eCQPCOZ
IJ0a/IhDwmiS/bPjPSdDzh9FKjnJY40UtZFbLXlmxi8EXaSkMPjTK29UsaDtB4pd
oZAbR2arhtAihUU2fYakSNOboEBRhqH4IzOGsSp6moDNPMujosOqOntBqy+9EmEi
TmaCYXfhuFUfbN7wLLpdBGJeFUzYbIUjfcX7BhOAVv9FLfhkg/pIiCfjulvYJ2s9
zhSxjGtGKvIWh5/drxWXoy5hPUMg4ejJhEv6stzWa5jf1M2RBWFfFvAvUAMvs8F4
+3RLLFidvMaxVnti+yBUsxh61dVmcXMm2eephxnQrWdCTPMSsQJAxBfXu+wFZrQs
ibVIgeKsDC/WfTCWnmBhxne+rSuxCkP550AxEXDXHzj7vCkqNLxchtj1EggnlJmm
NE8hJCizTud40HfCCJcLAD+NdSYVmAgvFPNDmOY9ccJOydqOc/R17ePYPVjw4GS1
5RnSj1eXAGXBs3bUl4IaXI6FkqfRFj1q7YwafSPaznVz71h+tHUXlx7kraEj+tAk
TN9jKkDK4DQXhiUo7/rj5lUYTkZKS2K8Hgi4lNlxY6X1rhqfhfhmB+LX3eiHZ5VJ
9/bCn25uOkt5iZ3zgDWW4vuIm0DBdu9ni8zl0IhlNCUaest57+MWBSTGEek5Y9+D
Quynetvo5lZIl3WBuh72nIOte0zp9I8qvQwDINHEGSv8oWfckhQlOqsVQcWh7yxe
nK6WbE2qGiKKFNNut7iPQrcQAQkmJITm0t0bfwt6//tTKIjTywB4kCCmKBku4PtV
oBi8P9K3a7FcXUQ4sbfDPz15u7CzLc6dCMYmwOwpnaGWMcS0N+cybR98zXeOWYUe
ZDsw9K6xdZGmw1fKgJNplaz7SmLv2GIvGJaAhc48Mmfh6UtX2D1sJPiOmhsTaAWV
8L/je8nn7horVLu9nByHrzH9X5QQqH2vnC36XnBm9hSw1o3lTUyd6XqRI4iV5+/k
GyY4TmdxgwkFDjTMvtrvFrVlra7LKaXZN4vHH8l23Le2eoFhXTB7Qjloe1iMo6j5
MQf3kqDVUDv7kVK0p+QG0OpBYgtGTYyZ+9lOstFcGbSkWZ5qiLtN78FUeWJ1sKw/
sDrJVMKZjVwVj37m0X+ygu4JQ4RixzX0uI5GgFVfPS/SSWRJqIYjWW9t7Zuq4h2d
5vbbTSqbpKSyB8Ov1XIH3NfP+AD6Gv17Bs9cGtSibFx8FVubsDVXvcYoS6ECbMK/
tV9J+Ik1gge4AnOV2JjdJ8mJkzyNWHAjj2DE/8utcXS+Lytbw+aUEGF0xZbSXJEg
bhQBNApV9QsqhEXXAReAqTrCSbC/8WISgHidEwM07unozojdshsnfyADR7Jib821
eAWryMma+7hqtoXq5ZnXi35hurGPk38c3s4r0oXT39wtTNORYcAiud39xZfJu1NO
Y27U5MdmH7LsXMgyvP1Jx2htoNHuwWKSgbZZgCO5iqik8BlMSJMoqRpDJletypI7
uQHZW3EMD8XbQTCOppRE52FFN238EfDiKo/1lhfkl5I6BtoycXcUlNI+Bi/JUMxa
H6PDDuck5ElCucDSblvq2+YeB+OSB9qwDVOJ5Dijf9kY751letBwyw7WKqE1+vyY
K5leSLfBBq1j/bHKP7DWBEwdYLn4lDp16Ye37gn3qYmf4xlaQxIwj3Y5y+OikDnO
IM44mnmhtZ4P5Mrg2ZP8zHz86sh+xN4pbGvsJoGSVQUZN409Td1YeYjeozIs2f+b
5iQ8Qpaiau5zMnGBdUdGx03hQ2YN7FPhcjsISvjKdQcx2IGP3bE4Gacw3kbBJgy4
NPnNZg71BTf1XhyabB2zXHLNAOWorpkURq9anvdBefODYgRzv0aVXep37QaFGLpY
8KyVleMXjU5Fsa8RVvceWTjVpolHKA1P+TlHQZJBNFnBGPpCKOmYj8guxWPD3Jdc
tE8oVelsE93HTvnEuYIFIJRrnO5q2HuH09mzRBDlvG2o7ZwXH9MPx+GkmmjArHsu
tbfkGnmYjL7Gk9L58LBI96670ECoEqTXw0qyr0jYfDRG/PQXeBU30V05nogPbCI6
Gh3mgDZFpb9V5w83WhIsbQnwaMTnJ5TKCVXbUPPjDKjYlgoqjyRnr19qKg5BkJeT
/oUbkDrmUDG/AHfAa5vNr3wb3Q0wso3rzM2Rj3jVL8cB//4qem/LUpMr9PRME6ib
OsZSp+a5lQGnVZQg97bx4Mw4okqqw1dWV1o3snRio0SkC1cWLovxLeIrkk2tbWMo
ixa+kY+fEc7Q5DrXEZqkFBTavyBpm0p8yDjkytzIqlEn9aBBruH1CztyiCC2+6t2
hogmchcBhHv7Qz/MeWa15M78DlfKat+L4gL/gknuJ9BGpvWpPaK31TszkKBOuWz5
HtUWTqeOrQ4asDsQnKd8sQCUOmS2goJuqM8TcNeiVm1JLwVlg1k/hh17mLIixL8y
mHbTV0a7nWfT81BM/+EW3JQZwc6QDewgK9GuKAOQpYPPUyCT7vryMuqex1KP2xZF
gBrEK3TKsJOxETe4eY1VC/R8GaLtUOzGqb9/8u48DvAohIWqcDppkMEq/4KmVVib
Tdjhka2O+qwABnkYRk9edFjmaVXmN9GVRmThAQglS440HMPuplw7OLGkf2KzKaYw
XuWaJllbPe9Ev7oCntfSDduSzs3SmLSG1gwS6Ys1aT8si8Jy4UMvYFNAVidXdAGB
uXI3QhepzXxoM/1mab40zun3VCIN+G3DbG5+A3yF1YWJ3FFEBfifbmCOmF7ecch7
j8kEjLwKVdjXLHpDi42Vis0Sesw/mCFiCN5/dyHEgJ1s5jUQVQhGmyOAZRBi95cK
qSFKRCNBYmMoANpt6QQBBaZXGSNuxqddF/Za/+P8S3avweoRgwQVgLSuQ1x8VcKR
EPni7qnxsGMN/j3gEH+H3E1TdP3tS1I4atQiwF3K7Y0ZEv1xviIboOn2r0rgVqB7
XrdS7AJi7UzI/ytbeTPythr6qctsT1BGca/LGngpK4+MBp6GkSGzPw4xlhXwuYmP
mK4BYcAsR6vIqJUtmdOzYgKKTwdVc6/rAC1Gx/IhIYBi0vQWyyCGJxSyCI6R2biY
eghzenAgD6e/HZK2qpz74SjaWvUg56cYDvrsqkHWhL6KdFBpngzN0WdCtJKSacpr
K/qy3kOgCx1i2DnzhqPRrx0a2ckYfXyhgOpEylrhQ5qXPniITnqxW/rxVNhZEJi2
N1akOU3ov3pgmT5FapLn4sVmNbbrzfGeE5am+FvTaqRWL7za0VZa9Y2+IdAkiaXI
oALsa245bZkGI7vwRo1+tJCAkFXv+xH2wHAjqwWosENbomljdXLDNuovnwrlBZhL
S8lC9e2zSzgD5gK9WMOkj9XlBwS17kyRmvsTXK3t36HAWpI2GfX6yD5v8nceNWpj
Wy9zdT4V/VzSB+HUU1lF5dkP/b8NCe0WDrFK+I10+JZFUJttETXAMNpk3HW8+nKe
E9auY2JHpItSeUwhhygNOP1kHx3mlkqoNjH4Gv126EYQSXXdjeknUimyARjRDCrw
TBzB9DIDLu1wK1QJi3iDCV2DIIEWt5Tcz63rdhVYe/Y73D2g7Y7auASSlHi7BD+J
IYeznLvmuczgy4BR1IAYhFGlySEjK19s6Fu25Xfd6Mc7ehTJYe1giFDmfiCwNqA3
NCl5agKvxkcDQ4oqLxk3S1qBNcR3NAgy/OUuKHlnHZe3zJSFYhAqmoUcR3iQ/qU5
FcKUzB4kZNnhgAaS6/+LDjSqGjZZEfjcWQZfjAhk4+P6TvaFjFADMhu++eLKoDca
MUBvPYTT0wecVp+q18s8e6rynL0JmHo4RJS4mmXiTQ/z4A0KpYuUsjJQsidLhKjv
x+IZ0CJp4LJoPzCn6sd3o9aAzZiNL2kRq7eiESeaZPDjxOIgx1ehuoxAkH5+WlDu
a2mMNg4fc4Od8JvdSj0GwdqTPDNnn3bbkLsOIAIyjDAiu1HyH/sPML1W9DzrnYj0
jKq1O/E3r7DCZaW/Ofd/ny7eSQlP2NlHd5yWyMLmikfyFNKIGssSTpzG8goYccjj
OZQ837e0dodhOPAedso3M8Qp+veaB1j65BaXzEHWDzpLx5v3gl1xQqEsOTbB9VIe
hmahkOKPx4xvhLBsbTcRJyjba0CDTVzJCPahCP7WoVvZDlQFVQKz9/tjEIccNadh
uLmQzjqY+Wkcvzl8PlNn7ioXJX7WJRVyvrOWCCzwFIAyEJH7fp8LlGOMuPpkG2Ds
TbCxgM3kBecdt8tUOl8KYSwWymbTvSgdIQ201DymPFWjx5HAsW7K+1z+UER0u+BU
hLZ5yVYU0PYRIZ2nJaE4TsBlHWBoKHvydQOXK1Ph/x+4eEIo5nMoL8C8A2UfutAg
+/FVjzQvUutoE3lhe5v1E1QgC0WaFr5bQgi86vGsnEMhLzOv1gsPSullTzV2DdOK
fRHUudo1DJ4SrJHEvphd3cELPgH5RCcEpkGKxw9T06z+8tinGX0jdQeiLxD3Kyoe
Uu5cAbAQJDKJexGPI+7FtJyEEByBTMBy18yD1dIadowYNLrBrmnlKnk+pJ55vqNQ
y4+5GNESMVC0MdJfjKHeRKgOdUz6zc2AI3n05+cG6pZ0cNPFRCR+JtWYd0P1d8b8
4pIjOkg95dXEUEVSZeplzpGZQXGWYRapL6+wB/DgwrGzcHY5mqnilbbW0ORtNL83
JJm/OF0X/IPPSGB827Ibq1yiPuxYvmNYu+8SCXeEDxBV5Ux92CKMopuDIgXyxpw6
DaXxYyWHqH06TdALVialsEfi+mG2+J61N2iRo6uMdYhXpggToqkGCnmF8diSNZVQ
AWc7oa4mNjqJkdNd+O6EM03Qi4/mmw2H68Fv9VPN8xVmXaCj3QkXhhSMQTBQYZg5
764C3n7wCCZfLBVMdhOzWBiCB8cnjM8ZeC3EXe5BG6oSQfzULkcat60vI6Tk/RGa
GjHHX8OQhNY+blyIJukZjD00M8KLA3xa6Ub6IPPP9uh1kiJ0RX2pvptjb+uWtHYc
CRLotbfR7it5cV1t6NbuzESTZuMZo5ebM1EAjAV3rElGST/BteCNQbEzOI7Vz/OS
T4+f9krchpS6e3TRZzfqAAJMxGidqZ6/UCKuoXOeKt99SypW1TIBRD8GccRgoleo
rN3XT3jHXJ1BDQuC9/ej2XUbbGDDQuS4en1m4eGd0Gp0jwjFjzCsjK/xMJ2yfl9S
rAcs0/r45zqqjOuS8btFM580mTgLc+liTIbqNeFNlTT6XeSJmYY7PcG8xy7d2ZYV
bp1Z6lpvayCRQVMRV0up31CnHJCgGDHqYq+u4fbSeaqOO8aIncytyDKWkC68JNfJ
n9Sm10HN7c5ewO5H8jmfA/OMOtw8Lo8axFg4PHKnl+KwT3B5vlMKmo9ZV2D6Ellc
YaEagqp2nytXZiTqEnw2Mr5tloZlAPgIagyYjhkA5RwPoFQmC6KDIfra1tR2ksG0
Jq+JIBZE6H+pt3UeVDOU8jIQPEe0bTS6yd9OMOo85ErXabB2Dhfuwb9ScsHp8YxY
uXsouTK5dvEWBH1KmA0S+V6uS8sfOSidyaA46Csc6F0tNOxxfKyiV30VXOicrAo4
Gm0vy38YxL0M5yUl/hB2T2j9qiQFOuh4lzQB93HLFgzwihBFcgL4qJr1Yt9Q9Mdi
2FYaGE7O2uiDabuksm0DM3Rmnw9XocJnXyWJaZPHX+Gwl4bcOOS5Pxr4jKot9YUN
mrJwCUojRMyouPxjyMg2JZUagLvR+RftVbt2KASNB96N0piRX6mKa4Gr71TUpvyZ
03or6HwpEwuRdyn4oboSq9zZihchvveW5Xh/wMu3hO9fYMioJklynwuvdbQ8Q4UQ
U/kQFz77Z9FRg10Oiv8wSJ+iO0EgfpMU/uGBxnhybepyxGMmUYQtO/HcxaI8midX
8vSKtRysWcWhgc2Le7tkloyHKTYyvbDJUDpOzt+Wp2z5ot+MSsVN3drG4aXrPnKd
y/yyfus+dudib3+BD+Z2ezDFS/aIcFU6000Odi8z6D7p9pmGnACRtZlrSWp4qOq3
j4nQYCF/pvkADnR0AcRVCS63JpCV3ArK4r/b75cMEsulPsQv16deFOmBAzP6OYi0
a9L2UaXq529JX4O/VkjXGGUyhKBV8TqSCFwbHhzM/+lGDD9/qe9XyUpSMMQCOMor
z19yzBtSKcrW1MowGzJE939Usb81fwoMjx1XFa/JfNm1gRGAeG5ng7sqnbMkkxcx
mZnyfFDy/wEhqKKA0vlW2KJHF+yI9gh2BU3V/ucQTA7/eA3Qw+jW2nto0gdQvXXE
3zKZ1dbIIJi2PTOPleVmBcjvS31Psl4v3UpOJKa67TfAcZVMQ31RA6evSMQl2Qqb
F9dHxR02HEEJ4ETNeu7wb9XR8L1RG2PipSuZS5mo3X8ntzWQmDcxwQknQ60O+Ao2
j4NsQe0h0m85Ob9C51LjC5LplVibWbqNpl1Qx61dPArXHyxAayQejSNIL/LJYCDm
H088zVwWtLOLJQu7sCYI/4XjMrJ4G3Xi7N/wyTzT9oxYePBbEGN0crGmX8hqHi0R
+FdHhHpzX1cIub/FzFyvlMr3SHOZ4/9bY2NCrEte1tjsBemy2ffqUeA5Xtbtnr0H
Y1IPXK4ghcy09sQsSNxR2JurosdpZTjz1drevhnSup87YcNZSmTa0gATNOSs2NJJ
0a7raVbWGFcxvDgV3ZElUhE64Adh6mKKi9W7w3aQw9xRl5g0dKltex+nNwET9BkE
guvdzXPx0Q0wYNS+xNtXDRx/RhzFZvrd7jwKUVB8wExWTBgn1ADwZ+g/nCr13rwT
pJZNnnMj3tiZMNpErn0kOeriDGlMO9Zjp9m+FTvwbJtE9Ig36VEu9DhW1eUKOFj0
Z2Xt2II8nB1r4uBlFFB8cykkGpYwYg6HWJyC+C9COl0Npmco6HDi7g9AMv9usy+I
nS0TxXmVXZ0SyCRlQw9BLiDP8dXLWNpDg7YmBzse1TH/mwkrIEw4YX02jnJ92B6D
JFgAv05OtojII0BfQrb21ZUlNViWxuFJnC6Jzhe0n8k6KgyApEf34jOpY2UEnrSs
PtoFJTJMSQKkBq/3wtLGutdoBWXNNDIfknjRsOHPyNC4yGPXAmyEdVRIlrbq0vVG
ZZOIyskxQu0Alzui12CXcj226ZnSRmvfXeetElugqb5ffaHP9ojAfSCqiRXn7jN4
TKSvef/+C/DwHUEzCMSraik3X7tUzXemOaRgiuNWmh+oGpcgLg59wR0H++n36CE4
JIhBtZVK1bLB5BtwBn6FzceWwqhe7plYOE+cEtHNkGgmWtUf0MzbtP7kAMn+9MVg
30GXBFVjuFw39hg+/PCGzH9wBowRkfdw2B6E/5CudIxWWSADRZGo27fAlgcnH4p8
wwWSZ+dTRs41YlO8nncn4qUOGeFgUu0VIZhjQa/qa4CHzvfmdfRoBKURQOQe7fMK
g1NnS+yoQL7elHIm5bBFggBAIFzXCcJ/JbXcg36np6EVY45SVJRPwXHWN/tHKOqT
OzY5A1d0Gvgf5WNSAmBEqbW82qD73pgCesJeRhE736Y+dupJm6ojy6a7uuRj9H8Z
nSZMt6gy1zj5HxlaMbvGFq6JLXEn3pTeNq56a/UbSFtQ1yW1gPfOca99/8MbCGpI
Ntdo76tsjrR/B+YR/1NM/mUkSWpGcl4iBq8HuhMryJd8llQF35dXOK67ClgDAGgr
+egopB3RqU42H0Juu2IECN7Lfy8EijuOjDqv0rEm3cQNUMkCDCfizCttC447QOx9
T7Ba/+6C9mxHGbP38AQ8RjK+M5mSrdEAvNQrvqyXuHbtE1P5Vr0mWJbGDeRkjrc4
Hfg7gu5woGAlerpGyHUfl4q8unkDoWO2PvufZn5niLe6Kd3fYZVito4HZ8rgSMzz
Y/o7X6NZoLkDBycc9JvInpEleBtK7uV5z+N/u1af5hLb3WM7zCFjwNB3613TNBpc
oxAQ8lNzMMhX6nCGLP2EpgF7UhA8+PHarShSvDXFmLLAi3cojJt08WvUeHd1fsxW
J955fK9Zo1lz1tJsT+y8oCyydde7IgGdmpVZLsoiiHBOaMM6MLg8D+6gq5//SD1t
aifpjgjaYqKLEwYzQlPzcAIQGU8usaRvI3OEMQ5H7RkrFsvGJq2vmL6Fg0vpz2WD
rCxeYoxWiIXUvUMvWAsy6xb5K+W7SmLH5F+h1mZWTAVU9ufVQl0QNDtZLNF32UMF
7zen9c1zjXq7Ua/Yd3LIJHgcByoTiBMmcz9R4AdI9otcqQxfSrKTtbojiP6OisfJ
qz6wel9uRhuy7Wqy9hLWaIkP0ZTunsjxmhe1IcJdXvF7G7fhwWN7U2CkmgmUK2s+
7vBylnLmQWq77HCJZeZ3komzN19fnO23AhvEl4e+5GoIY/rwojztbfIHvMWnYheh
8I5IbC58JsYhTQeErFXRzANjrlMAh6txcLz/98rIGLNQPhCQ3tjWbhk2zKTqQvbB
myZlpvY3iTfb2X1ppfeobcYJXFzYDfH06iw/K39yBA8uOcDvxw0EgqmipeUOjYsg
6WbPrR5G8+8fK/ixYQmG4QcmkRBwwv6nSgSvlxm0BPwUitJu7P6Kh+ZeNuSi2fa2
Q1OiVzeAMr68BoFWXAkhOAG734Ou1+GZsrtiRcaocO2KsFm2gQEJl6A9thYq4+dj
Hw/djeOwaW5cXhf1aVYn0ozxzgv9ZxXROFOJLKnYf1tQ08DgWTv60AiPY/vKvs4z
Q/LQuQIQ89Bqnz+/NUaPP6gca+jwnTdnAElTfwnYs08RGO+2k2hhh9zTFWCgqs26
zsOVLAMqubtneq/yDTcy+FrpOsmyEP+1Izekgt7/VKfYI0hDUFME7AGFFzLmZzZj
JnpsIZXKI7wKSZs3/qdSpW5H6fw+z614KLt5ryKTHLZHS7wG1PvOrwlJpldz2iip
/ok2IcRnAhNp97On/SEmi5x1LsXgwap1/IsDLrEXD/0goM9NjtzNul76W1063sJk
GAm5Z+y0txa90YEc7zK6oemOQFR1UshuSCPD1/gA/A20e+qhX2A701o3zrUOSGjr
WKkhAQPmDjyNraOh0iB5bTmp56dtoSBaxUT53qN4LsDP6pBv6yiiazrNk/HqMx/P
Qw9awqF2QSm78hNgNKe+0VEotY3AwY3ZH1meaUH4aQj+jTs0FSAK3TDHbqDFMvw2
8W7iM+R9Ox2hHPmTsATCn18vjFEat80WGLf1847PHuGNGqS0/lLhIkimVFwP7PFe
XCLxLR6MAMQJd0/UdeYOinzhAu+ms+YVJx09rcI2qg2BeA1uqizEnIjAMuYunSkU
WhJ9J6QQQLYOWT7A3OUtvVvrDkqr00jm38H3MQXPO/23B7ZVYsdu20O3+6MTXqmO
g93EnmRzdtH/gQtFg+/AoRgs18gRsW+n2LYX85XW+8bW/ppL3BHkPe5lE6MyIOok
kxf2flBt/lVgj4SQXeeYZ/E9u8u6O96K8Vp0SHRIdSSdljSegN/Fsx6/wMk5bknx
/OIr7XzGJ5/kwu4Wuz8zQcqXayfp+wxp8QhB3RpmA9k2Qtbbr9IrO7vpr5F8/myD
Xe0fHaw6o8Dj2VqpF4Dd01E/rX3MF84Uky2Oq9e4FgE5PGQpnjb2sBELM54iF6nu
byIuVyVOCO3BsA7+VoPEh7BKFSjyZihDPwGJ2blrSb64sYu0Tno1aE+RDBdBi/FH
W01Wpf71tzU0P0ErMDcYb1hEkWcpenBbFMwtTHujjgpuw9b5BitngZCCMuLwd6Q6
xluXKDoyUeMIeWH47RNH7UojUIrIlwZz7xkHsGbp1cHL8EAra3FX7/nXMHLGWu3e
sp+uVUR0fLys59MyukrY3dVwSmGUrzcYhwwBqPgkvYIzZjyS6CGVl/8dTBKag1D2
m8x0WQCJFvUrofMldy0pyU7b/jnLf62DjbD1YnN6gS3kuohY2icyegFtCmMhvihh
oLxpVXHlDAFs1zM16ILFwUOfyXBMX9b2+rnti9ppVYmR1NvxKUWJ3ZctFO6xfg4p
8K1YcjIJuKCW68MnmWbrLr9OQQ5iDDlRLTo75jVmZkNvssiebH1X2WU++3sP9OZS
xqEEG5TeF0F00BfUVVCeFz4qUrMCI8SWFNQMJFrAhSWCxxbTn4mRikm9DGFJPpQp
UHuZCnY2x6tjkWGBovGxElcAZMXvamRQBPkhPvjC6vdLyOUAULUlOmizlSWhrnOM
DL7EKnEwbu8fXiAqPCXkphRIncTmRIdWn/iB6ay8yIKKzWHn3iUyhLhc6J8uX7FK
P474HD6sPiXBFiLpOgzY+23NDI6UtvumEkOc5tZNnWPNaHomBMc4siI5v/jKDjJn
ujYQPWft29x2UB8jRvPxhSloii00p60XX3bBQCb79Kvum5c0C+6av9TY5x3T3+2H
JRxJcwxjPaOD2pRgDWSeltsf2sS1oH0ODBfnZ0RFRWmxF0efcp58YTwdkjboeMOl
xphTSsRzuMNa7N8pdq4a4bFicUA7C8kIKdxf77eMuZTdKHQDDGFMF9j2Ig4f00BC
eriRendHz/AlujkAfnroskIPorUQBZwlLGfmJ4rRTMdy8D6KUfuZDQN9AMjvUT7Y
lF5TOkO+l7TxslXhHuo5O8nxsl6ZvQeMV2AB0OYq82gLpjZuJ3pdKqfKOivJn6FE
jDjHHCWg1Ksg3IyTQbtsufbRNS0ixdSgqVoTwDj3QYVtVqmf6ktUdY63GwCDq2eb
G58p53OGqDuvBH+7z8LtLNxtvxhr9HHa5gD4dZ6il4sEbKgLX8n+U/62IrBeFetH
V8qO6sfu7eESiducZuVMRWWVsp/9Wd5sSYlDJGCQx5rxCtGArJ8SUutC/PdSdYQE
Ma52Vg8numRfNYZHmbfFLc5OmXtTsz8J+llCRiRtFiHdVSiQfb62m9geJgP8cdmb
hV58tZoDnMJ8kH41TyWxCy433blxxgVJga1nctNgHaUtt2yqNRIUaT8+7FVMijxo
CpxLotv+0LokUOv94+hB/TrxM7Ck8+K+8WdH+HVeWBPhQlRtjz8/ARieaZeBdnT2
Sx7oQC7cQgQ6FA3SRlkY/Zc0W8FO9eBjvIZMO0GUQcdZ5JoiW/kz+dYyXqOxnH+/
nuZsg2ARslGrLfzc1Qvxd4lyurh6+38GQlSx//wAm+dtPXoqGdXVPg3erWEt9Pb5
r0lhN2LoutMMn6hJ/yl/g6Ms5Ee3m0fjU1f+JLSU6NjtdTBleGRs4hJrIQHQuMA5
7wtdPjwC4wwP5nD+QA70JPq1cFu2YXTihe/PyA308gv5oHkW/YMYee60u1Vr9t2u
LCO8hVH49kojRHdG8y9qFr82oqW/e8q5UAwMt3tf4hmdJjiZKvQUqmNxrObc1nLm
TY5ZgIgvhxPYLoGW4swzusffpVPbBX5ixRu9JOHOkmvydCDaDWxIpaCrWg0X8o4m
lSvB8GlUKdpBIVds1W1IzbAD21uB6IVEBSPVq3DkXlvc/4l1aQC51UW+npMYacSh
Yq/dcWvJ1kCsSEWIxjC0B6vZKYGxJC8CfpdHasLwpsDtjSCZd/aK3U7KeUKTV0md
UBVi8M5OmHhgm8R5iOfDUebRV6ojizt8NxFfPK+XqijVNLiBb0EXI99S8aFeKIfH
Tg+MVGInFOLfGhPm4XgAgEu/EAes8+lXAHOBQEXodOw7uzb/eWMkismvI3XhrmZ5
pS6YHTmlIAaNjsQURiWqDl0ijcv3vFxcNq6eTBm41vIOu2LyEqlL6C1qT28A1Uzq
vdwX3CpVY2j1f7ZeFgvYup+FoOLr/nmpQIHRRDNqi6yJpzTfG3MxVhPVw6UqrOJ3
LbAuI34CA8uTD5kzIHFCvcGjdVkotBwKPDhpOXcZq+ECh+wvpl8zfdOeAGsmPanC
HWakUQgCcsl1DhJ2PKLsB7msHYXRUxmeEukiKpbRa/6tLmmQRq/etss9+vT8YGB+
o60zEymGpDu6k1EyNT5t85BLltuz+60QB1P6tPvraONS6s/sYImeQGD/MvkZgTQI
m5lLkq3U4pfgyO4jhxgZGaDmU1cmp6PjWLHYJeOFBNGjfjaSY81dNjLJrg8nG4iQ
kks67/pdBfDofTkqobwpwxTkb1TEXJaX4joHxIObwuSYFyhI5+qpUEumseNj5ST+
DIc/eCIXcxx9gBGcep1AudRBQXqxA2RbGmnOH1orTcpY4DJLL5/0+RWeXdlj5gjB
Iy++ySbzVaz6MOyAE26W7dB1peTlwCsahaGW/Ccy4EyloN6fIqsf3kyv+F2Ur8Da
JexZkcdPqVDDdZ0SF5thqiPqJVz4mlrZN9MWDUFzsBplIwD2mNhV2X1CQrus4C7Z
XumNOfmMUFAy1MHnwdR5XTvRsfBsNaLZ9hV3diJ/vdux9Wj0XEprEbL8XJ2cRxMX
CQPAPYLH4Tt7oEII6rAA35KViGKNcyu+YMjIiC7SC9efB53Y/OXcL3u9mwDzPPSb
vyNkCXRrn84T9pfP5cunhawrfSQAxCHY/FmnKmhJ0gkBaD7HtHZPkJQFAD+rNrP2
XwMIZ+uDJoa22yUTZYQCYU7L8v5TU/MuuFBkr3OFnIGIrF2aWpsaW8qOgztg+Ka7
wOO8n9ih0p+iXgQ2FPXkD/n5tWmt0+eqvA1gvhrQrUhWzJd7EiifYGRVHSxo60rv
8Tb38tUmbsLskwxUIeR7S6pgdrA1BiZb9iI2KSNgfOLAJoiylPXvyAaogwWgrLcJ
1bzk6oeDKWj+gSX+hpISPOTWTr4tnJH1trHK1ZxmgaP2xfemisDjRQ8iwgUPoYPq
G551JRYEo4RXb6o/73uPNIOatY/JpxjEYC7M1ZviPx8MQzO4ZTVku4xrDhu6z3JI
E4np9SF5mr588bseFfHl4CIbeVg18p0zS42HQEZVsimQVYjV5hqWyPxfP9rAeIpv
ZC8jVmn1nin6gQgjvhGCRsFliPAetHS6YIJ7VQak0AhwFBYQ4AyK9EmO8KHjI0/b
iLHEpKZVPfceweQA01HlkKJMaudyDYgmHjpk/kOtIk2SM2T0/ez6a9lxlSTOwlJZ
bKgKY+5T7J9M4T/qGEajKb+wp5AOhNRnHnmVot1zhFX/9KDwQBIxiaOes+KxU+Yi
NJixU4OGEgBoJ4ju6m46Zye3385HVYST4rZdxqQPAHw9dEeFQpN8ROtm3Efuz1qi
/hRJNBKXKc5nb2RqVQXlpW4YqaRuGyClReDfzjf2E/so9QVIe1okBfzSCSFVm+Zf
+a3H9yOfrjTwSGR+hfF4JiTAcMzYY+ErT2+VykxmICSJGciK+XuX7TN1xAxQVBmL
oXBKiIhqvgc+cGTCrzq7dOhyzuPOu2FT+YVtgtJnB0JCUgIteEq/vth8cuZ7WrBC
nfKpqnGK/bLW8xOi2KFODdNuUjWkL1+81tFptIOExVt/bnHnriQg1WbfpbRKzR+k
Ymp66fYSLySXNLTyuAVXzUoiGw8XGKUmKKLAIJeR+JtiHzNlyZMNX57ZuotZYzfo
5hBi7QA5BiPaLrU9IROmpSySkC4kG2HS1vU0Its7qLedR/osji5Wzif65nu7IkhR
OQ8Qgm1CTwUrON3lJL4KFzCQ8b/Xo7JWhkSy2NVbn3XXRLpRFMWnb2R5mTLmETGK
25fDj6lu1IHSJSDdCoSe7uEmFVs0Jo/lKI40p5OCYZFHzmTN7icf9KssQb4i4lRz
iYxyGAMxJcN0f0RYzPwvwslrFo32mStnp8h2z+CGx5/iWcyuzBBvfivpPBBgkK5v
S8ClUG/eMGsQfjY5PhiM7BAxMmyLKwGkdHwEhw+wv2+4KYNEa/HNlrDqbl9pIOsq
klt7ZpwDfndhidoPI4DEvbgNr/L1jBOQhxQRmqCYys8n0p86NLAMd7gCxCBtGt8Y
QerR4hztx9cJFRSWpXEmxrqic7vQ+UQa5194XN0BOBJhYIG5zulii+tw/WnvwW9A
2xoNibPke1bIOBvkSXgUl0o5TKA4d+9GzBHbe8/PGVfhjl2CI6Zs5WKH5+h8OtEy
nnpAZ8bzCESiX5WMkmb+gSnAY1bS5xAYlNAR1/IkTGDcmAtg0+T+2lRu2nYa+IPY
5w0CMvpxWahodzeuSAA5KBm7Dr63z86H1f0aPiIn+DxosMbjvrPoYFy6XB15xuU7
viyfGmE5aClJUvTk4EDBPYry2brsQ6x0BwGnf9Ai8ejCJhMPGdkAtMIj4lS3bsEU
K4B6GQMvFT2dqnJmDLPnFvVpHYfdX+rV3YpKB1n1HObUJzqd3Q1sKVpaptBs7IVx
/zMll8zT37IkV4wPiMPiFDZiJjyQa+Vgv7FhUPx2CFWGy35tkebGvrV9Mh2zOGl8
49scMvHV2EQja+jCZvHPeR3HjX6obGZPa7gaMeGHfGSSmBDv2qE5iWivWHP2EJSR
JV5xoV6eSIrOERcI5Nu4zMPCo4MhQpr7QchSBNpt1mEftWeH6u83WtzSVNOiJnqi
5xpDNNgKbkZ4TqZ8zKQvBa1hLtJKJGfYfrMbbj/tCvsecYCat+VllzOHSPwzZAOy
RlJdXNMUeHiwELgFj/5zIAuX0KFFJTQq+9wIcO2mIPklScSZlPOQr5i1SBnDGFI8
sxfLKmsaUvQqjWXi8c0uFrV7dbelGNyRonBnpWzU52r4i4biVc4/njTnOnYXAf+m
Pu+QtY3uZKGN0UbtIdjapLxkEtZhZZVuGs2zA+up+AC/WRCh2U6PiO/PO2h1ZOcw
t6IiYhh8AOjkyGVmFCvkBCt7guTnQ+6dqd3B3bUMYkt/+q+w+aG6GAT8dCnoeWsw
HxJY3bgA5vPIj7uadfK2tqANnSI95txG7dFS/6/0lMzIIXfJD8BWoVHd7r68Wx3b
w5+abY5u49d0yt1F4FnsxgN9yQoNnRVAz2jLf9djA0A2oP1rgO9obq0eB6/7PC+O
jFOoYE4BLtmBEgajjBeG8ODYU/KeO1psdnDLtucRWbLr1C+Lf8qTRQp5sZEN2kO9
mEFABEytk/93kVAS5Lu1qzPmFaXrp5utZJpXXxrJQRqXwYE29bw3cT4qWS4WWKK0
1ywtPVlINfIzsahSquCzXZG69xUQ+NVvm0k2sRm34DIJZgDMK3iTC+OH+Tm3wAYS
hnFRgUUUo1O+9xZT2cWU2lh/3P11a+3VQw+4GDipOUEMM8dCac/iOdG1yIwk+U9L
GDbvbx+LaRtFU0hgzAyur4Td8+GWeLFAq25MBC8g25i1DpCCRFswms544uBhdXqW
4neynAJaL9C27F2TfBpG6y9oPBSPRbamIrKGTizTeWuFlcMi+2QtxHmQu/LwwRGx
Qwv25l76sLESmOsT5SNBTyXeA/6e4hhGH2Y7oBP/n6HQr222e3XaxpCiIZO75Oog
WZQuZM7TtRiaxlow27FH2Hk4sKOucKnk1lN4j6JK1n3iZVOPCt84XPSyO8VC0kTw
4fBA8qLX+p8fPIgN0QZI3Rkfrxpiq3/cvsN+vsmDEA2YWj7F5qavKodR/nyUFuo2
XqpQ9pMpr67awoUtX9YWMTZahWRzuoxzeeTe0pm+lB9eTCHyL+8xgqFZl64M5azE
3oFeg8oaZCzbJ9VCzT1rKCDQZzkbM/9LCzL7JrOPqW4OF9NRm+qWTFRNFNVJEFdk
+FkSAXJQxU4yZuQMN/8OmSQ/kJnIA3naiKbO+iymR2InX+ScceZImmndWC+BzLdH
16kf5bsEgbqedVsYCnjzthtEeVxDM5S4VV6rit4iuxBnaR84Xol3fuAhgDhKtByl
Hwh6pUd5+6u/8KSvjjt9u//evw/P55TDoNegTUDWIEvIZp+aswfUbCV/JLQlGk7u
1ToBrs4PgIk73onue0C/eyhIzR4N8Np5CnCAxDm9hcptoxPi2o5Mk0CEJFyNhHIy
wNx/f0btGdeXCR77yQ1suBBYJHLfq/fER7PYGgE4EWfDWjyLvPl6yq2RH3HFz1np
yG0S/nIkl08xZH/hGRQOuOvX3KB6r0pTlzMXrFs2p5qcChS2wCCtS8NVkixP+qOn
m8v/guUYLKqqgMHeXFDqWkraWiYT005eUt/oXOEZi95G1NHAz0+8+0kkudWMN/Dv
hZR15ilEgWSSHVRYsbaM7V82VC0ckSvvjbT4six09i4AyTkG3xXLEmA1vBkf7qoj
+/AiZA8nj5fvQcbt14Bhr6s15uKQtiHZIneSXSteodvZDNacTgF+88mqGwDSe4ds
1tq9qeuoD0dZxxJveptHMyfi+0ix4CwvhZY8s8exrpc2Y1S+GAMp7018vR/EwzvY
oImYAQCWcI5P62+eX6bzjZRwM4H6Ts13e+Zb4C1VasQSuTfi034OZR6PTvd8/r+z
+bK+N0PB0nx3gWFmpR+1qpcPgpS8v5XbDh+lsxhBdHQ6diO610yvrIq26mx7+VGV
aM+xPkLK9yyFEXL6DYpFx2STthxS+mQOV25AgcjP/1lvMF+Kex5Jw5Ydy2GQxqqw
he5G2ZL1Ef3Ig4U2H2y3WyU3at0zYduE93tjrSohf262I9T6YbgFbYYuJ/NH4xND
RIfqsgViWywQYMVxpwbUVSyuYYOtej/4xPJJ4LxuE7qi+ic3RBS9RX/6Y4LrQz33
PuXhEHVQ7Rf/sy+lonKGl1AJD4Lz8Lj6Is7mBAXnwp5/mziWKvBMIZdfgK6RG8WT
IYoPVcMYavduyMyjRRnoJfsli8m+q03UXAehQNhHWcs0TDbGLx9bc+g5K9IccObA
M8STIgpar3B5DEZ1pnc6wc53ECITDV7SqgBI1CLp1AyvZjCpB3VHbNZz39BFboQz
DyxvhBKU/V/Pq9hTpTcxt/4hmeCGsgpOyyW1iO81Jj/jOul42iKMBL1VBi840/Pf
cqt6KHAYVbMyQ9c27oI6uianvTdJLg6yV50kgMPG5N1AECeGCnFMovWdea11//4Y
yqs0SmzYttxuex0yIEgYF2Jj8L+PhV0cyDSSSpEs9kJ7Hje3u+WYYHK0FBV663PD
cPpThw31kN+cB6kWtcB9gblVI++XvHyuVLw75lF/oBzmC1/KqG9GurOp6C+nmUMD
lAHvvXItwg62NVQfhJ4i4KBS3JnIiJs90Bre/uaU6Oi570kvJzVPtK4jz5czfM+e
/2/degnHjpmXw2SkT235tS/Y1hjQsBAvKwBng7RI5qu0mkP5qkowAPJIttAZnjLU
9ctb3KqbTiM4FZGHALS8ryczqB2yJ6CX4/yS/FRvCt0f3sraTzKRQL9GDYTyD/aY
acwSRya6x5nxsKyOGmzLtvU0S5Ho8kbehqrCMReb+NvGxkKc3B40Wu55khLm8kMv
g5Z2UxJutGuJDEY9uY3bkznv06PwZH3JVSsChjNIbWwWhYM/k6lCQiJOTLbhygTu
KCOiYL5f2Lik+bx8zeAS2rWLeEonDmGcDGNGS8LsAuoPAue4WHsU70XabmnJacnb
gbSt0umwes/7akg0YOFRt3Y2DoJIsWJ/nt1qjvl+DpMlxy4T1lTa0tRzRsxq2LqF
S5+9TS0fBH3X9pCROicy7OlnH7HldSMy2Qc0g9OUzc89lDLGVNaJJefD4AawoRam
fIGwIbl8ZHAhwe1QhoGXxve2jugDOlaXw2HU02/kbzny0MO3ZyNbrmHxdc4kzHTh
9o+wyQq0BdB6VLwBP8zfdscSh/190hycjs9K2ZuMzPUnPlTdeqlK1kiLdhC8LdLi
73OjkDHUyt1SCJaB8eTTXS8EAbs42FgfRHx7Nfj5O3V+XfdTqCyGNfkivCUByDTf
CYsL/jC7XrP5yHAVdlxkXwX7+DzgWBkbYObEMEl9w17Uk7uLi13LrZ984QIwb0UQ
mUUNWfeZTvMvZrE7yNO0hDkVNHFndG6NfADxHXJja+Z58T9J4b+IEy56GvB/JeGb
vXVT5WQWx3HIj3KQ0CQQbCeLd4s1AMGx2ng4Hhd018TgP2GL4FdFpTyJXISiC3GT
vV+LzXUm5m7V2M9gK8dxpGg0lWyBcJuv7ErReOKD/tZE5HKJhAeyUv+SsmKBgT7h
KeAZ0BkJv1h786+0zIyUGPD99kf3sKp26bKatL8Qs13doqrEp7sPRR1sWPovBXbG
+0KTgSu86qkvYxHaGO7gX1820NWYFSAMUC0bs2wNL+fWsQruQZbRyezCRcyAuMv1
icyei0UnB3v8t4/dPj929sUCVX/iQc5f0BhBlzl3liFHeHiUCX0/eTVADKEFdTcC
hPmjLk7VUonJNqkFVhXXcwC2fy2Ga3P71x6lSM9Nq/sytP6IqPsNf53NXkuOb/to
KQCOhn09WT/x7MNTs6KpBDdEanyVrXy45pgHPmxnZ/e8EOAu1W8RQE7nZbwftXKG
pK7BTMVGkonEv+V1AvOpdHspnU72Gqu8bKgN9qYZY13NGooPU/a2NNe+gJFV5FHd
PXZZDGSge6oICPe6gtnnlSAb+89b2tMIC4Qq7GtQOUfqaTMoOdX0cD1KIp73sv5n
nG7omYhJ2tkscyJa0qPzdAap3+KOmDbFwBP1d6z0vyYQG56lJvd34vUekfnOkbZ1
L5y0msBZmuzLRR5K1q1cGouAAikvEM0PvY7Y5sl5am4RtUmvh1tpGaO/wexBHVmP
xVg6rPfbiDiok+DqB4SaBx26u4d8O+qQyx8FxwaetTxOrvCIOrACpody5drFqgwB
aaCh3Vnq/+4wAsPPX/H7SxYuU8cfp0nvUs2UJytPibXYcmXbp+rKMfV6ofC50DYm
GcTMvawUDbwDDzYhRnn9coQH9j61Z+YFMBRc+2DM5ajVx6+EwltqREd/35WH6Ray
dW81zOvZmMljmoLKsNk65Kxpeoqp5v6+SU0PTsaaFlxV0tBrfFoSLqEo0vK16fXn
jI7axxFoU4annOjnLUgy5UgtJTyMpwOLj/JdMnNYehX4USnv/5E/1Ef9yjEt4JRJ
vXA5qSh95c3ADRxUGMY8NfXHovgPcVomi10qhP22LLP6zBUzT5WTd1pd4tUL80xI
G3huCcblLqHsTVHu3sSoIv/9u97/7K52XCA9HkRhU1E77IOtUz9TcWmP4Tns6rJC
f9Jxm8A/i205lAq1oNqnoIXyH68i+l9++jLu0M79V1sSgcU+7buJSphUv+ZIY/Iu
jtR9s3p18vkRYIEFDoISHqMMQD2M9YbaNSD09jG0dSDUE7D9JXEYvQo4tqUawImC
k8S1cdX43PawGlNk667KhGLDUmdl5EBbFphGn1EztWmx4ViJTpo4Yhz6914MQBMB
9uZMsPIbSCh8hUd/hWNfNirXguufVHxXDoyX6+c8eOb2tnRrI8BMBzdJ1blkRdll
4fGE6VvPJ0JE9RMvibbwLvb48mHHirgRUhotjyYtxYdE1BUttdj7KdwMNGhh3C7z
yHEPdU6AK5KinqkvB3nAgsMHH3yjkEe1gQUt0QPB6nC1WOWAQEpHvI+dSkEV7ozd
E/7i3c4yzglsrKn70wrSw4pwDfAM7prsM6xMmDVjRkk6tph0QYEooR4TqVkGABbq
M5KRN4kdKSvwsO5RMrTuAhjQ83PwabFoGUfEXbaCUSemmN55uvx7sVEPJPMLoULj
uirFt6g6bB+LXv7dcEfDiHkpZHtyW6xyxvITKICOchx5u43VLbijDKIZpEOCiLry
xQWwTE+FOL9MCZlUbq+AV8wHG6hhHO2MXHCLBPjSbzpLZFKZqX9LkOthdDtjoIN3
rifcKIgQshvLTg6aZflQt1xTnvhf1XQrHcrrg1SRAyS3eIU4yzoLlqqq3Q8wS1nf
osRV5EJsKm1IYDgoArOkbX8Xw88v7G4cb8/i9K8GAH+bcsHBDaXlg0SurLP+3AR7
ERnfigZo3Ga19d/x8Uj6qTA5zVMzxpiqgnv39HgXbL3HNissnb0aaIkzW/oPHLqG
5eFyawiSV+zCORJtliqkDmmsia9k/PQpWVUEvzhKQnjXJuyQeCL/v19KRVaR7I0+
oBcuNKEhWw3hrU41dqXRRkvKd0XFlKZUEUwFtHHhEvIlkPozpVoZF1KjnnFupe6w
0KnagefFGvT2I8nVXQdFu48cyHbhabyfXZKa9Jluoa5cnGZlGAiSwhI4hsRoCygv
V3UVW+n340R6R9fRcomUa8rAtOHlic4hCKLp6z1J+nML3j2NtR3AKKInxwZae//I
nSqxXkQ2XIRamI66clB3eHCJ8XGFQWFCj3CZ2qCqMezsIzo+WfSK/xkoB5rwHhrk
0rwHygQeoi5kS5/S+4PONLvaIAbJ1MhBXHNvk6eeKfiTZtUmgL1nNB7Dn+NBH+13
Qz7fEx4ZAbSwR/2osVuu+GTSAQk+B2PsAEIfqJzBoLuu15JxHRbf9vrAIg57N6/H
ESX2nMBi5U06L0j+nhHT3AlOP7a3c6pN1idOYr2IZiS9DLrmxHIVn150ULrKpK04
aAEO4T7/ypJut+zC/w6DyWUtn758ZIhkylzRgtA5JCRCEWW49/WjFnW/a9YQzyD+
xXr9DV9+BITAk2C2ErVSRrbpnC5XnkPwSabi1vQGqAxBEqYWHhBtvc5bXveXE0eh
R+5MUylCqINGkSAnO1yLw923WPIw/ijlnO1GjzLmQJlSyXtp4ArXHtrxeb7L6jh8
BKF83i9ADKCkHIVW9du4FeHyyOIrVGloFbYIyFbGlCmu+4S9eV91y6Jt8t2RK3Q6
DenJ6JcIiVbsAtaeFe26K4oQIek9R3zXCfIm+HP3WNe8iNoS1WyXEuJprrttr8us
AC8ma2SR3dhULIp0kZRYaGEHjhVuMcyocN+FuXMTr38KtHBMsMBh0FTmxgbu5GEV
A4gGwWGSgzaUCWmI95zkD0fZG6Yw6OfOiFB1mGFdA0GEdmhHgZBIz0liKzHBcM7B
MeWUhIRHPp57HT1Dj1gqgKR3rMcTyzev9PZv7KNf8W7+BVpcjczPN727hers1kCl
8tPrssLJ24gV56wpxzYAmQHNKSozTze8ee3a43hrg3C+fyk+AJTRy8Mw5nLvw72l
MrEZqyafgtMmeJbIDbmoLVlE4UG4mb7WK/P2OGS6jokID4J6DhUIZ0G4GSTFXUqi
3rRDRkU4K46/96MypY1qc+ET6+Sh0foe//wrZSrwsr8f+d9M7emiiwZ3SY1Fmbga
dQN9Kt4Jbat/lmptKltYetIXzxvzf6cTsl7gctgGWOGWrMot/vAiPdpl/iFd2ixf
GzlBh9DPi01tOBkQN92uQBsuIP09CvDp+M82RFMSHtMSvJLpIRkv0SHPlTR/f8bP
KJyKUoRwFbKkpSMmGo/2+/LsgJ9myRHqu8NhCNnK9h5aHm+ljpEuzCSKXCfpWH8Z
1omIt7ERZDS7poRKIdF//rUEkAT2ybPI7p8pd8WLOsdlE9cK1U8vrNYVEUg0rVL5
xD/gqcq2CTcWQMCaYpvqM/6sUK7K6/KOH+TkFvf9civqUnCWQJNm9HrNZzCtnjaA
V2NMuwVf7YJxZMKXd5WHQQ2jg+gAEhwgQIWncbieFyuUSmdikZQwx+aANKzuxsIc
lGeu84pXx3E7jjGyt+EdHhUqCDUdduEtkw5ANjDOe1Ys5GiGV4YNoi/v0Bz4nHD0
kWdAo5oZ7ZB2qoAO4UGyzTkJC/AiXvZyAgUBQyRqtmqzqTaU96tjDrPC0gEwQC6G
U/2x9BUskq+r60LOkhEYed9FKeibJ1Jy9qK1FT5NQobwxnvbfyP35wnTOvj4m3zS
kR4r9dO2aA1lRfTJlrmTZcvnIuRJg8JWEtGkolpLIozFopw7OnrPILoEcImVaPfg
lHkE6y08/4NA2zJjbWCcSyYaZJk5jNrKxDSLRrGZD+mUeuyZfZXGx+3rlszPLtMQ
o1+ezKo0w3R7a+Z52mWrJooGmylQk/togh+rorqkOQjUqnIe2B966D+nEiA1WSLS
Jygjag63xt+mFtRB5bS0VlX3IHMt2XNI5OLXSCplCeLHRuPbdg2fy+4peKwl6OTx
VJzBsb+I0RtfPY9M0+okoYC2ie6yUX1Pd3JwQ2lj6DC7oUwUpmIGXRdNGWlok1iq
bBRAMQ/hTeVpb4gzu5byIZ6tPW7gWrgCBh5zSnNlpZFjKwqmIFABg38DHPbo99aQ
fEy6LoVHM+AjXSUPx3zbz/JlxIf9ek+Rp4d6aKA7cjEo9LtF2QXLotrvn09WlzIs
YsCtaKiWNen1SuL3C0nGdkISX7ZlpeX+5z+2ET+C++e/ucegLTi0m7X/v/WVny4Y
5Tkx3Argo3D/b8syLoPtnyfVUewtgyoKWZVfJ2e/JBYblQ2KuFGiWYCIOm9EPyFv
3JsoUGTUhY0TxAf19xcdCecksVpEsWnUx9Gk7tG4XP9/u9dWtSI8COoS9na6P3Ww
nNzxPzufOonnX9fPy8KJVXT3DELIalvOBb9LNETHElpBZAXGUqAAFYjX41yIKTnU
ybxQu8oG+X2ZzULHAhiJHobqWdYLChN5OTaBd6Cv7HuJ84mE8lYCnrS8z2sl/8yH
WU3wK7Q1fgaDP9CKbr6OLQh9MRpbGApkRXFP5lyqxrhbhZyRFEmLydWSfAtTxk4o
NlZxIcBsLBHKNQ6nOAKXwegjJK66IoXEJGF13mYpocXIkeVoV5P+77wF2jwnWKdh
dxl2otdsdjoVtXWQNyMYzw0tUa8q0LNV6dAlXVeoLXqkkob4ikPWkMDZWWp9wxVi
9wqGx5jTQtVjkP89Mao/Z+z7Uz1zNyF6sbq6zqdrB460HT8TxLWVLVyAImG9i+PD
mO43HI/XNM3eprqu9iUznEh7TTDYSNVAUDWjac9WujcVNQ1cQFORDo6EzgKJRDkQ
Qv1pn1qKNsG5pOtFC2GR5r6lmwPuYDlGycLTjMaH8AWZ7dVdFsaCQxVnaDdaudxm
yRwEe6jO8VTKVORaqaKlxmwsn7G67MYOWYN8J6zg9+gnBJqQ2nskne5Pwk8aF+jp
XHjZt8NqBMutw4ahGqPVYBjWyBxEOB3/hEhCQ3upi9o4XOZ+XAcEJk9l05xEEWg5
dSj9VfNAFVs9QpfGOORKoPXeRTKfIN7xwHfbAGg0IQIPQTBM1/Sck4BUL8qLfbQM
ujmzGyyDmrsaUi6Tunh8t+OzJgdkdCoHLhaKxZShhg9i4UxUkRMpvJj41RGxRRtH
drr7ecv17g3SPB7KW93uNJXsR1rZ2c/e1u6QiAbqJaC5+85K5Wp9/o+nS1VZPWb/
HBPJ0Y9fvPQcmVAOMwYoflFXC8am0ZV4rAbIcZ8Sps58lOg7BOkjT06i1K5L4f+2
h/89D3f7Y1TxBlEmV+XXLyfrIQU9l3oJWde+UyjBPz2VouCVoOYO4128GN40bb+P
B0db5EJFFvDQeFZ38hMgElwuMa/dUWrrzJ/Qc5YyNG7b6mJClkETMopj+1MKY+5g
yVz3XcOEIW1z3Xxwqcy+Rc2Xk5CgFJTPdTYVSDroW+GUr+XhrVdBVFIHPbwxqBG0
CjlUABbiHcTP2+KT4/M7Vr3CADiuzsYj+b92yAcKlLZsCk9sU90BEDxlUZxyRHFz
h1T0iuEhE6DafErQ6yicQNuSvqkwOk3UVWvqZra8K+v8J+mPwqpEtzKcPFljZN6W
Q5qpkowuvWJ3gDrS3YVuWyl2nlsQvc6hGD2jEKZmVTWM9nx0yZbaqhMe5TOXFzQw
r41o/MtXCqAXkF0JhoeXIYuRQYv8H0zJTVcUu5yuK2oJcipe4b/aP00/XQtkE0WO
HYRODiwo2kvfs6jucQJOGbKEj1/8EIcCLT5xonI7J3dcxa37IpfsicVySv/yD0Ei
Yrm/EQ6o6FfogorzRMpeEoRYwu0qsU6GFPTHS8vTTFZJqVCSncZ0CntHP3bxjnAs
f5C1LFQ8m/ppDNFwFN4zQa2lj844AUyq2dKrZRq6OVojQHK4xrJUBgLeiuaj27Ja
aPE8/IL6pCEFPx1QmrDKLe2ha1FXKqOALSMmQCTF6lxSexHW8Nwy6UixSru1O9/n
BZEnOiEAZdb5qGc0SgsB7nOrJ3l3jQ6WiXcnT/GMQIXAgtP4zezwaEPm52ucFhKL
yVm4RQY4S2ucS7+r/UlgzEWqiRjZesTtYXXEJhnl82LzvGVXsvtz4dDUJGO3Tfvx
LqE9juBgPpkZR7OsuFzWFP7ZfjHM415ILCwg5Dt5narFRosfOF70OVwFN1jDHYPe
3CmUz9yAv59zlzU+sJRgbyBSwzHuQjgpUYYaHmugajCYP3Wj9u2PlENuXTHSeIB6
xxpzayzSTHEAN426ooFBkWQRp7da9eu9k4kXJ18uRZrTf2tFGGmPTpCtKluAEuwU
FVcO7Rik/C5vmQbWlmEFMgTqacqz8L70puBhtSjDls9WZ7jEf8nhvhnudBQq34hF
fLaz3zprD8ny6UJA9a/C41stUy065KfzQyE+Iiq0yxNohKjKmkTFRT+IQ2o9hgYD
mg9jJVMfU/3YZYeM0FBRhE09BO6vdUZysIlUZwXT/vFC6uomWh4ZXJVvxhbMYZtv
TKRzq6nJpzthXCikQCTHZUdkLtjvH62aAbJj81MkWeOKHH+b/eQNkanuJrtwsp9q
0zaxkZpD+FNwnBh0XhJB3hAA4JTLgLg1uTbwlgwjk+vNQNCulfbHKNqRbliTYJ4I
nHqHTQGjWM7R8mM3hJG/rf1fDVd6ZJPphEqNpnNQDOqAXCAJGLPrOj6b6YK3y0n3
PvQ0vFkMDTipEHI7T4PP2P4//c0JmFJ05xMFE93XDAyjprEoUpnc2u/POEKYyFY5
81EAK6HQB/8jV45viFLNgNdf7hY3kUdkaiJbeKcuuhaca9ZhNRcMkrnJHU2qls/4
QDSeByQw+ErOy6dAtrAoIMLjzGADe5WwtHQjULRphPOaqCAu8edpp8Cak+lWPd6W
vJzzlL7pkfpksvz77q5zAIhsjVn/wpeC6TeaVOB+yBMtfEeVE2rzAy2k8lxYURIZ
N1yjaJczXIWMHM571TT9mMaql/lvSkgvDAtcPbMM4m8gc+hXJK3fs+Via9gysmQK
ClVaqaM0HRcY+Go2W1oqoSXzqprPvJcOEyOHlIIw0ouI9Wg4wVRH0JWr4avIq2vW
oy2vfhiWQExkPZcuseIW+DaoPuZu5RQJ9huy1s8tNgYohaczB4wRce587qz0B/1Q
dRaxb2Fb6ZaoIOnZHE3eJMaQFRAzR1LP6bowgbpp/8aiNo0/szs+P37owydv1hFT
OclMoalT7eP2y9AEk14yaoap2i6rBURquI13h/DgDLh92dN4PmjG+V2aTeNaaTok
x5q4kNPIWiOdyNqEgu8KFy+DRg5+x8aOhIe613xfin0dKUSzJahcBMbvYpQ3QyrG
ya6uC+0TPmrmhn3fuoPu/xyYxNpv3l0UaR6gQWqn8YJaFiyFZq+CRPNp+/RxWcW6
2bgdbtYMvgCsDdZiFsUpWvXjFZobg9N0Hk1wbE8d4HOg7N82CVNBMrSmBvniGmP1
Mp5vXj1fQzWxMkMNUlS1iTbuEhHvbL9S1tBspbygNj02uVLnt6iTeSATN/WtrLWv
A/RyPZw+CdMLSXP42iWwWfjeoNJzJC2IfgztLgB7pJyY7QK9bm5fV/M1r/g4NpWi
hEK4KAv9uqYlb5XXOl+zHlJesZ83KCeWwoQTLqTulCocxST+Gv7oEB18GELh98U1
O7OB1mGTfR3MDde7RJOMt+4VcjQo1/c2YaSbI4u3DBvNSddhDE7lPmSj0/V5uQ/W
FBqTXIWBEUcstl5o1J63T4s93lDhJRTeOtt09MF2AsxX/niO8hYGK75c1tmWFv3x
7K9J7Snd+yLmvWaYpdgWp+MfDrVAr1ljuXGZ4XLyLOeYR30BXze1XpBgJaCFVp3Y
sHjwSBWV63t5raWcClNW4BtI67ahhPdu/M1isKnv4XScUP2rTOZDxDLesbEn7C/m
hyEQFZZaUDPDvAJgHIEcYInIA7c/rgAsSY2ztcioUXn0xLBWz5C095Rxr5OrDAlq
enFXroXh6/Jv4tTJ9nRHDTkf3wveUEKY7haM8FgsA5ZSBZwJIQAGa9DC/wERRjU6
ztOVSwK4+PsWkI/jdcZiszyU2bW04BAgk4nY/op9Uuz4nej0AFnn5nurlRJoQSN2
829EhBhBDKXzHKsVuGeaLYTpJ0hadYPelcRL3q/W9jARk63sLrqw7G2Szt2JYG44
7pRV/d4/HmGWNhBSZs+EuYQ69IJCf2r1PDDWEq1zY824fYJBNDYzAszkJq3raOrw
9ewjsAZC0Aozv1ym58DIiSgjLh2/ZliqclUSouqwyMK2DCeStaFulV6MEDzW1QHc
7P6xvX7eEcBH8PfUkrkbNSB/w9XXw95yuHRMC5VQxILzcu92Kbs/B02tCKX9y2Jf
6WTxGe8ZW6HoVOt59dwChLaIiOIiW1VCpBFWdi4HOXS5hUCyM8gvb9rC4i04wAVj
2z7DfMmgOSvDH94d/XxLwaQdogBE+Nxb9wm74T4jhslDcV35m4gu0ePbSM5cw+El
j9U4X+Pd9ZSN5ZUDclbPbF+HpSVMYyYA1Mma+wZwBUeDbKe1Ec3bf50Xys4SHZKu
gkJpaVYbk5aAO8K6DmBvQV6VhqM21YnMLJdrWwojnhezCu39iDHMJ7ZOEkk+jWFN
WnsO0naQicv6pZwI72K2LqsUWhKjNAHr9VS/mpAX5D6mk3aQskh67VPF6EjeH/M6
odIoT0Ho9csmPPTeb43wl+5v1Z8rLvqm9vIsYb2jl+vyHGWe6wSWshRuFpJOD0Yi
8Obp9mryVRs+r5vZYSzF3724rgX5wx38qiXFiyACtYwLn+yJ+CL4a6LbW7liqAKa
fEvS9dI5N8ddN1Bgd++7mxj8RzYQZUq6Q6aMkLNAa1o8c9Yo67wutzY7wKBRDeBL
8fXLkH4gVfiYe2u1lG8BDL2qBPWtIGzT0oSGihbszfIexPnybLCjh6OaLWw9rfTm
NP0prMlPl/16qcAsS/GtY86x/ByZfK/cHk/FqBgD3GhKUBUMOIq21SUnmOEWR951
tCRBgYLWSjgyRC4SK5UxbdL/20iSZs0vjRIK8lyfKeFhJ3bA1dP92WT2sePRvwuR
bg4yeePzEXND/P5gc5HRcaT5MYB3ANd5Y0ePHyLnbNOrTMfU1ktQYb7Sl1jBgN/m
nRyQqqDW+07Kxax52LKH9ySWrkX7fFP0f49Txsr7CGhSaZBpu/rzbofkll7HVp04
PeZLw6tFNPGXtlvo7ab1o4D3utavgFMGq1XSNc5FmR+eeaeIzJzS+jShhrrpuUbe
YKOXlShTEBtSzetYMw6B8M1Da5DnNLAyE04a7QJRhac1hfYZW6Yu6hO+/WyOgt9H
1eY3jbgDgq9zjQw7woJ9erI5ryS7C+iIatJdG/3Usy0/TfnAkUR5kg4Xk/VH5k7U
5exjBu5KMJ7TeODrd4j8fF3pNlfQt3BmpDhwNt5POhrZ07a2ilQi2eMdIhCs3JB0
p7W16v6uvxx/X785XO3wvn8h12YP1I4zCOZ4vhaywN2ywn8op+u/CJjifhxncddN
ZFZAqcVnKxQvIMAHIMM9VX83zRAK+i3KNz2ZfuXhyK6LMgmVf8Tb/yRaz2s096Nz
7bUUu+mB7EUvRgCMW6vaJnWNnDCTaqNM0XLXQUYuj1JMNla9qU/B3jByDSEwNI6+
3FIFxsuS90fhbPKmGPOTN9Z7q3X96ykx3fsxuol3sA8T9/RoQfEdBwELSJkxaYaQ
Jusq2VPl3ChywQ7Ao/SDJ31pnPClcKXzBiUYdrp7E7UOQ1PTjxJ/J0sAQHesNnZj
OE8L2Ybqe2v8FArLCZp4QgnoxR3ulzkbGSg9W0fL1WLBBMojGDZlbWKq1mzgo764
PjSLblfHKvpPriaiHPtau8Kb3anXYlvLPlykt3AN4rVMSma3VEHrYR+yA87XpVkb
9BiD7tk+H7uaaL2JW5O3fbQp6Frk4brxIOjkKU1EbkH6PwuMct0UmkW1cGl8/MN3
krFZP/Te3a8CCoVsxL/iL8w8ls6vlfb+L4Qh9V0wpKZMCeJgyzqna2qffDISKgzF
H9uIjun5Nij2mkwGYevuD2Iuw3S3oJ0/u8ObMn2Y2ElErPXlWeY/BGhFJVgpax8K
PpcRra3I9bQccXRVL/7s5YSVs9jySG5T4kZLqgi2rwMrSJOdccpId0dyo8a/przp
xZkydGP18Vo7Rmh/GdkyTmuMz9ImnudgXmFhzQ0Hfgbs7Hdr7QG6H31JaElbtSNc
EwvYpb+pPxYqtIeEqOnvvGte7pdLCvDbWBBjBHD73ivSn1C9W0cGRFUw97nHearT
wlszZdiXDySf1P2lxuJitwPTU+lCZBTRtJRDgURDStIdj7cj5PE4y4B/hnYpvYY+
Kv35ZTNwqSZ29w9H9waa4M4GYN9ZisiLowhe3VoehYcEjjKHtKytO1OsTEnrhqBa
QPggPJfMhqn+0oQqMrQrizzeLnkfrTAQ5u4STwF9FlQq8s/ZHg3kveuhK1uDHnA7
ilP/vVBQmLWrcRRcv4w00PuvBreR9LEOYfYS3btSHswDdbqDWjfWbbgZwyNZzsgh
NiIDcgkDP8pxrb9nVZlUD8AM3WqR6TJBZIJjr/+aPXFOdXJY8KVyqfUudnnIbF1X
fY2iPZhr8sAoWWRuQJ6mAr+6lvStNzIpAZ2lrrmIUxv9NbJrWcSNg7BHiBmCHsPV
P60VqpAzAPTx2mjNNw6PiZOOXScCKPaxVG6Fb8zzf8O8JuTXdHfxi1pcuNZ2T1zl
e1freDShp/S7Zmy29jUdlnOtEFTeAkGZo6iXguPCAxOnPHUiuaI5vUo/C1SeTvFp
52tnI0upVh6Wwqlag8B6d1J4mRYXeGB74FxXf4M7LHW1Boe6TpITAJhGirZzfcQB
qUQVU1a9LIy6/M/CCBQxkU+Jx7ZQjxCX4FpkX2kWgtTUR74bHUzzYYeFqr+0y/jK
2S2NWO2+OpNm8KrJpqOLKqA9QM/hDf5pN3e3LfSRZ+mf21lVXhvry9CT1oscpIdh
WIhrnSVlUUHVMfY9n18bLFwW8gSfOj6Dv0vVpVLMZQIwVg/uGsiOC6sqvwN3mwN3
zMqagke/tYauu1WgnAlWDy3XJRaedo4XMxuGBOWPLtiyw5kYjz+9hQrA4t+WtMnF
q5urBSQZp4Eg7ItyYhn8/fm2GVy+H3aebTX80sbLSdbJtZH/4LZlx9vxGCq3LjGM
dShSff6mMr+Ad5CSZgsQA9emuocmSFESM6HXdGJO0RpXfmltjrL27bQOLon1ew6a
yxRcpgyHeNSffud//rkv/TkdybK4YUOHwoF6QKDQq2dF1p3ZB4Vjj6AcYVTIyidg
pewKNLdsxu7A15wM8YrFadhW+DcvXmRtGO8YOaj5dJ7r3jMXY29GSPSxPQ9mYc+9
/aC4uRCQsUOS0kLcDtqBMjoZmErkzrkSkUMBaV3Wvp9V5YcTqFVBxNGx1LtfMBVH
LRXWTfWX4ekFl3FzNz7I9GAi8kuwvWQsrqGGNoJgZQyzgFynZpWbWAYNaXk92upC
7eoK8YqCQ2TM3qpnQyb1+YeS9oQ+yqxDqUcw8fHWmXGBcLEQe0XmzEwq9g1dLwfH
AlIrdoSKfJw7qojMDFi3SAWwn13IfAwF9ImX4r8ZEmK+LZQ4LHgzbIe0izFDgz58
a8v9rMq+YmJ1zG8bBBVudh6i43bsX99XCih9Ka7gafHNaiGJTJqD9HTfeoEjp7Zl
S+DdfLWXDsPJrYwdwahE5gMizDpADIgTu9pl1KMC6ZasTPtrIuklBX0rnEkFTRyt
Tf0Sxb5LN0mZTfbPGohvPB5pI3CljWkLgfXo0nnCfgWau+l0KhF4v2qVY/USF+B4
6F/kRIArqyGaPlThFMLzmgJLBPvlA/eM147h5RmB3KctJ9j4EbfUJsEncgAgg00a
VuIQ7GdsSXU7pqoF1o5d8bmtVGrunuuWB6JcO2ak+EKXPOBGBWFZDdygZX24Ada/
fsOXFWTpAs2yEWixsKpz8sNbty7ED7uYahFtDmC1uv36ppfl9jARfwKLN9MmCTcE
6Lx5yzaPQh+qsYORvJ8zsOcmtZOmaia6G9ezvmEy2NNsChrqmcPqJuDRBRyg4Mx4
R5xrbrdVKKVjxNzvrGilxIJtOQJrhoMxPkgFj/gXGuvv418q9aKYXeiE1SSvA1Gs
qwQZFIVAhDioSCi4LP+KqKfr+KGEOMVu/klnddeAwTcnU/+YWZmCHivGvXn6T0dj
V54eOwLmNt7Q/pD85oRCFK7+2upH8vaDh1C6pfqJaA7DDeMTKqGk9tP/ztWuVBM0
vQLJY4NT1HIEhH+I46N/ycXqQrpzbAMjFf9IJzeXKRRIhQD6VjCEtQXzSpekQQv4
zXRtK/81XONSUdOZLGXz9dqS6wmJ7CuYSx/bG7BO8s1MjPXl7B85RcDtPYDLk1B0
qn/BlsdFQ4t+Sx5xow98XJC4dFzoHXvqSTDvaViV9Nw9/Mo+MFaDlPNO4UEAPcAu
MlWIy5oyX+olMlGPz6k9OBY8NY9Qc0X4d1iNwsEid2D+iSEJYLqQAGSsrgNXe0wA
9Wc7hhNZssiLuRASHwMnBid1ag2SCQyHk/ta3KqUr+eVuXrvdFf8OKcwJ+ZmctFN
U+FK/83QdsEmUhBftXT+yG+2ZOIy6jmpl/O9m9+F3tkH22BxXN6bJ9BgrTHrGrPs
568DioiJpVtXAr5XUhd3HySUyLOC+51jMQTbXkT/bfhdPh/vI0jpyuezHzJtAJFJ
hFH1Em+zbx7UeFxlaeurHFBdk4QIQWc0v69/jmuciTcyiYTHRgXFYqmSUE53GLG/
QiVTb4Tzu7iqzmmCI0UnhbG3u3dB3bww0OaiV82NSBHA2ldOoHRIsnPSGLLg3PRv
c+kyMYuz3xYG1mMT3PnbgnyD529MB8BnyqD2Zuf5RIV5oUfr9QkjmA31T1xQH7QY
gFOxyyuz9NwE89oz0d4Lt3MgvtuJoDheRh4LaylWFLXy7H4/klMFUiJodl7RN2GH
HjpoLVG1jOUY73MJf+0wA87ZzBhd7jfVJKgUxEsDzxShzTSi5hUAwmA5eEeBwTNd
Q5NxTXXvNFCXrrMas55XB1+0pdMQ9FSFHM61CNtOFyANhfM4sH36VFWTQL3sniLM
YHZXdiNSQ/Sa2DJuDdsbL7V3NYnwmMgqPk1Py47vMK6N5L/HfVDIJWBwlm/KQ2yE
0hVbn6HYrDQtIGYc/W/xDPXKBJEQjmnHvdBO77yc18lqQkEkxP1ZiiCdKQgTM3Za
oebHQeBQvsv9B9c5rS9Yd5ALyLI+3zO5mzc6iXZS2mXghKq+Th9GqlICGMRnFkMg
qElTmiVX7oVu8nXlHNZjQMryYRw3RSeaB3G8a3FlvB8exUkwgEUp4DvPGje6JtjH
pDZoXs6C2mphg/wTEZ29Qb6Hl2uCSeWeHMowUSWYA74t58nk7QgcxE1Td9UBoZA5
QL8+u7EmyYZ/w/drYghLRfzX/K0z/9seT5WUMcTNpaQRuxubvXPaLGZZRuy0PjDz
FGN9vyqKKWFHMcpQ1UYGsccACOOF0Y1tKTy90UeBnbZGRGy+6yMi1aF02RUsIG3w
62JKQpe6CFih/wxBilNn3u/+MSWfNBVaQUZF+KsRkeP+FkRBgOKCGoN1AVm6VgDm
/KH81JDCPe9/J1UDBvw2zd7crctUL1GQtSv9PHJ0Xfxd9u3fabdEJ6y6GPlkyuAj
8UXTmUdCAnKXMT02GF4aLwk1IClafdDp/GPMSWbYYsiYAsA/uLY22Z34TOBsR2Hf
mZxrbt+RbxWki8Y1LUQqGBFm5yLRgw1eLyCFOYCi7/hVDppZ3JbzMaGtRzQGM6HQ
YwXC7S1iy8/XA66bFUU8PlbtgXgQi37kWRZ4jFsqithtw5/ky+/gxI+euPgrQjeg
lPdFTmx9+PEcAlwE4KZMpRU2xlKdorcblhJ/7rDSvEQoy/k1yhTizs4tjPPjdPNx
UFaIyDlR16St6x3Kljc/UiycztXPlkDErdhBao/zcpzYVDoHUsgo0X+vIXyDm6MC
+LCvFGpv2IkCcq0BV7pkBiF9jhPD5Y+q39U78YmOM4HPjaMVbF7p+8w/CWve0LJP
CNtBHX4/9K7d01vGBIwIN8mSmhVahJJePcrqBLly8O+Zr0sxlfREou/+9VGmg/jE
1KOi7/RXTaY0mU7LyP1Igkgg0uvm5Bm6dv1zdwG7AtOYaz4Iu9GZpcOcevnHIh5z
QWrKAs/pGStx7Cw6KVrnfEDdRgx37U01TI7fIUvHxtgbJ2nvcwOVFBwmneRljWqf
vgpvmscdcsedLI3FdcSZl/otRKadYbR+6h9JNgTqV0mPmmpFgSlY+cCI1mmMgOkq
KX73+N13VbDdoAwyVwiOPBGPnE5XjRii/SGWWplNK/E0RfyS2x72LgX8v237y5dx
fCZE5gAZZVeaDivgVr+LFxqu0KLKWCwnf/d1maFqZT/WuxMczyJKwSiisJYkvaPF
qbW+3fp9wOhHSaRa6glsOMLh7f/6tVKy4L6WW5X23//zpCf4Lxvv4C4SLFYSvmNq
cXdkAtv8g4+H5z0I14kHIbbqyHB+nt34zpwfSyqRccnk5jrXKBziPvQemEdKf6KU
ldyyWydX8AM7rD/qn1Fi9kfTk/dePIbCoEqKgXxi9fgWpggJ6FkEjJ5L6AMTb0ly
YVBSWvV9Ickx0kzGA8LRI1F9WBQ/dqDdSEqEcamDdBGyZj/cZks5gAWVp54N2+LF
mFQEEGN6nCesxRxIYDFwahy0rQ3mdJORfvhhaGMdON1RebgrfAsPrtDl/8qdmK8l
+KYfSdKtY6YjJvaCJHzk5gyvQLg1KMY8nRCpxHxR3VVEV3+DZ1TPJ6A/uLZaFgGL
vFtQhe08jQhHTNjD40lQY0QWpq5XNZp7q9y1JscwZCclN9Ns3xaVwmvbvJ1za23/
aHR3B8JrSoT8K8B3K/3V5j5uzNYR+WQUmrLDfn3mM1a+9wEaUl5UoVCODJ9P1hW2
jG12ZlEtdxRzYIHxGk87/QdyVMvHZVYgp3dvE1H3i1ZSa5PU3qOJVB8MPz58H6Ee
ELVBqGDHHOlRmxrygnU+mViQ0pEzacoIaT/tIK3xlgoDLpmhkYmQjc0I9GMdCmEh
DvMCJ621z8FAK5DC5J+J1ZbvUuyCdenumxeuC99PyIL9DDLmNfbkCUP4/VUtS/aD
wcmrSgUCFKG6gwGzacumRbNpbtLZll9MhoA84t706Mt30/q0VvcgDOVtJTbDJM2V
hWqdt0shVP0aPQzlOFCgZHPocDx+OIt6dgO2fQIQbwWd20YQVRLDskEF8DbOeekx
VKSrhuElg0qFJiSHkTrh/VreCHnaKnRGuqUg1B/UC3lMyE9hLluGvRnVB0rXCRtT
W5M4dna9W134MIjtCrfLXEckG9TIxNHPbMuh0lJbO68bh70rETEpT2DrJy8kn65b
Uq9Y6gFUuWZluluLYPX4+qyvwpijb+90o9yjZdqn/a55c+QpxFqz43cpOuBL0kCT
b6+tKMvHz6jZAjzLmZQZlqAGEs2Y7XIB+dtib3iaG6UsqQ7+lAPlEf0OZJgRr6xP
uLfA5oMNF+JdpFzj8a9hhslZi6sQdYUUG4hn6dhXhvn8wcIkeD2st4uKG9pPTtFu
E+oEBSwoFxtt5/y51L3XKqKqCdG+6ry9u674vZaBgBTNnG/kYDafFLE30UVbNBll
7FUyNuzkVd/1qcTg25JoiHbgEZ51DAqwVP8JURwSVbNqD5VZgXiuXE3WZkRelgAr
m3QLGBV5dAewPjGCJSmjmMOlUrv80Uu6F9m+1U1MxSWApArDpm03qgA+f+TUA7UX
bwn7nr+mjX21omZ5z0zMk7wzH5GWnt8B1vVCmDHX+gBJqi919tSzmLKuWx78cGsW
aiNZ6+QJRDECHrhxTF5p1BJ9cCEBptBDJpzkViScryETXQwBBgFTDR8qr6mi3CyF
Dj4CnbSaH8oCcRfm5aY/jJWXjuBfZBtxG+doje0gsslYbJWHgETMz65cOXx+9/Wu
cctO3GtpmQrfPcoU8h8UpU91A2v0bPq8acO44Jiny2lpOdcxpK86DZUyv+8Hxw1n
q/nduxAL2hqydAchi+QmdDOGZ+SUkQ9uHmXy54NArR514Ju37jgDX1R1SPzLjlOw
t/yKi85x94VPOKxoKJgapPm4C2cpz5oDH9MdlfihPP/kyCz6yJCv6jBMaK1VWypC
KzGeoQVwXrAXwSvuJi2s8wh8rjEu/MSiWo6kyOGQm4EFfiu144kEDJB9yLK9y0Dp
97d+oUlAQ4gATYqtSNq2haG8QzKe4YVLI0JkoBwIUgbBi08cR44TqZyQ3R757VAU
9U9s4UFyx4DfXwaowj1N94h89u3TgPoXRhHs+osYoom80oS25Xa9wyG5DNDKuamY
47tfyLud1ed1ObfhRL/RIAadKRqgkQFFJ5EVVy3XTN/3pUtOaWnvXuqHcl1rLXv2
obTGQrvwyb071uN3lc/a6/pl4TUMNJ9CN4NsVV0reZDxmRkbzG3SIF/qDu0dJwmO
H7CoOdlU/aRn8Z/QUDJu1EabBjVvh7CHWsMxdlZtvk8SdoyJd71cZOpVai7nKo/L
IhwVjg2Ln16B7O1jUkTP7FSAsKwXglN08tKPotTrAZfG2fFaXTndvjA16tfPyNcM
SOKxwwV0BOlYtiCEKFWQLOWaW6NhO9kQ/8aiwLmJ/cGI1E4EmBdHtP71UVSmFxtZ
Xls+Bkws5bNXThgR8A/1kaqNOjQzuff3sIBaRw8z8i0QSvUxkphh7Gygr6vGl7Fm
t95mPzlw4TBZl6zd8v4H8rsrJFSCfqRJdpVB0H37Y+LK8ZBHGcw8Ta+d3YYZn4ni
qJQcSOZ2yBMPvxCIg4pYqCszUjlFZqFk0nLeXeijSGDQmTWGcXTparEM0TqyPwzJ
reB902CwJQtIBciMSyfvrzrftmwrifW3p7Mkscrmw35h3uKAqOVMR8XwW0m0MR81
CLZ5GrG1TpM1EwulXJw7Q86LXavOUdSFl7j8Rr6QYwcj1f6BmGl6+D4sizzAfDXp
ryiskYhM0OmWh8WGZD8FpqaBRKn/D9/RRT9UNR2smBhoHY2ipFsRqn3ln56uZTAI
w+jE482+i0LL/2vUZdMtGKuxrA5/cMcW/FgToOJWVhnI28zJbGbLoY/ZzDc/fYxY
ExrDUum+CWnCGLvj/90r/L5Rud6i1zf/KAapJk+FvvNBzvkDFEgskuxUc8NzGIsu
DMFglXyDOx8qet0ucY9AQrvcts4tDrxkEnW9hoYN96Ejoef3MSa2DBDNNt+A6y29
ww9y6RKynivI6zq2Pav+N40IkSOcu4j4gfkZhmI3hsqnY8x6sA3v1g97vUOBSze8
7vtmdFtQQrcwoMFJ/RmeZEcQ9xU/Q/4W16nX1kxypW1S14yFP3/Jm7T2KvLhqtlr
xnUL9FaHFbepE5koAYup8AMWmGXLnMR+qKlxsBMPDYnKYVGgt6qcsqa4oskbhjNR
GzyeHjiXUUNIY0r8XMbWf9HQWKhClROE+2Nbv22Ebbrnz0AMAju7VO+ErDiMxpm3
N39ngEarbQm/Q9ovAqgp0As+joGJRDhKORB8f7F2bw1RlTUEmVA8TAGKyKVH8fRU
ANz5f/PGcSKIfFX+wGcia41XN336bZuROuYfcQs4599LH85ZoZNceHXAG9jnwkc0
tXnDaug+8KeR9UA0dZdYpvpLLKU+2usedKCt11TK05Qa4hQrixQ6i0SWlROdBfIe
xWzM/I/cCSuTVvdW2Q47KcUgjtKSqnHkZvMD4RJ1ZfkJZDz8s9PmjJNVzX3UjBYN
MZWG0JxW1QkvhEutcM3n87UeJ0WipgPo0WLLpnlUXbCM3hA9FEpZtOqwL55GAJQu
yPOJALTHITBJYxhh0oLrNYzbeWmiv/h0l7wgEOlNakv/VecxUzNrhU+JhRVC6mms
1SzCt5F9y0cCe9BF5nfYGs1V3Yzty61OSu0Kgxq7tY/I9BLiN/PA3LKujoC8/jiC
BXZRl6V99U+7yABggtplvETpkhb6JsCEUPNlUgKv6SgiyIFitffjUbptmXme79Rv
j0xStKYewAXOrxZg5uffd4CUmzHjPRKv6ES7EPSCqQOUyt3MSUg0gQOUf6dvN2IP
KfPQK5MrZqBjftRzSmbMMIbt4VtDwTPykzaHA2P21mFFkTDsz3a30AEY2Kva83qX
UahGU21Mumz2xWIpqRLiQJvkVM1kBXYszlQWPE5jJY6epke2h3cWqN6/4T32IZ7j
zU9a3IvOAMtGYjx5aOwYq7eNevIwlDvazplRBKAtru2HMBmjuj4FPxI2bKvVk9UQ
hHl2UZHtwiOlBWV47a7VGc/yUMynZy7M50BDBHdD9CHr5hVQRifx3Q6mqSvYYdvx
hgZ5tYEkTETlpJ+OkRdoOM0x4jplweNmF4Py52NqS7LMjT85TuVgyNhtAOPUwA9s
10/qDZJS9+NURbwBi/07DgikLSGMag6qCDE9OQtYv69DUU3UoRw/83W+A8Sak98l
ild7b3yGbCnhVMd6qOt872NbGPMRW9lON7qlwjHJi6Jrd/WpBPUPQGplcm5WP6GP
yDVKUGSmBZIKyWz3yVF8+cHjMtjZS4la8PS6KHyJSCGJZ7H3r6V4RjF7jNK70kiu
G8UwI/VYwQWngpbHx6PQi+Dd/DV/zm33YRk1P/l7sII5rhOa0DcXtsCvi7adIW0g
n19IZrqmJVtfMU3Ba1Xr/Si76XSmyvzIPNGAuQYQ/Qo957wA1VKZI72Zs5oO7Pkg
c0vTXqlqVQ1sh62Cxh+8kVAyeBonpJlL4c5gmpPParMQuueGW5Gfw38yG8uY4OoV
DlTbW7Re4ScOOq36SJ0kTgzSZXbBzIAZwUZlZtb90UwRVnNpcHhTTj71VBJK2hCH
34nfKAly76jR8Buhx2SNRMcJBDqteDEHoqJ/5l5U+RU5GffJl0uhgGbHfedPaPcD
D15uPCCiEEmGKAOQy18eWiQcHgRAEhEJbEWi8gCI9WO2bXoHuqv/H8cvpX2WqkE3
NSdJ6ow5qu+/+VPEtf0vgc2DQdcfzIFWJYKrPo4bEm7H97EwranYyN1TINU3ieAq
caQV36hEqwPTdIQpXLhJ325/5yH5qYErXJHEavx6t0Im2IuNkSRRD/VaKt58ocQF
ck3iqKUzgRvrK4jgW0mQTVV5Pf1ivds/MTCHWVJhuhdLAPU01+0V5LgjJPJ5rvCn
iMyPWDULUKJubZDsJfRGUuCaPZDZ+pZoIjBv4pnOMoU+QAXfkAP856tBgVLhJq09
EyZ6uPYmoP9aqMUs1XBfTlq5C73xzWw/WC4tcWWSEscjrK3Scn63KBGF1K3fpIy8
DcGquBiom0KL/gVDaCeY7jQ8YdjDN3VIWZqfYBKcHpTEVyAXgtkMPw6pRwcKb3tX
xn239CdJRRHGjMUQew47In9trpYAAmH85Sy8bnsaqAS5T0NWVfXM6ZvyjA2y/u89
PRh4LHIH7XuL32q2QrMyAqqNhcEGe39ctzsdcZ+qMWwz/+Kj+JfrolxKVJgwJQX6
HnYvvZSBGYHPf2/1CT5VtRtVXh67mnbiRXExOSh0Q4dTTBUi+Uvc4bZ8S154qj1R
F4Fu0oD0vXmQC/l47XYNwmNH0Vn1uN8dVUb1ZfewMTq398jxnsVPWwIQyHj76CrG
6xbnqm8rV/ADvRM98BAFja4tlfw7yttSNGvYVOEoyU4u1VxnHkw4aQ4Muo5birpW
LhwAMh21ZDV9oL6yOdkKwFphculABfE9TrNttZHKvKIg3bMi5NkOoZ0R7i8V0td5
DNDOqFz8+RcoB1PEr9eU2CUbsKAT+g6bmAbYjpmu4OYJAUaCfgz9H/V3yGRdWCK+
yPCzOAeCzkh5OdsWkt18yoNfdgW8RBFSgUMQw1WJzokh6qDgUkR0lvU0mgp1gdwY
GaAcfaSJOAd+HMmpUwdUI/JhKJVgNDeZpkAIKGUieN/8YdXoR4fFavZjTz9JOC9+
eUi2VjPB8/VtDqXsacATM/5FR1jjO3wijUcXynn30A76k+jTCFBEyDffkjATgFts
w6zRXdPJxNLY+oXrH5pGNkOdW14SLSH+6yU1WNVbu0PuvLfU5X6IioI4q8DTNiY/
L/LGXXYhizug7qSprDLSiqpTo1ggqCOXJyqzHx2ML0BKE4Aa/osnKYHoYydQgnF2
SKjG89heYOpG+c0K0ecNmKiczD9/Hv5n/xef9+b0zzrMVYS032RsivzFxFYJCkPe
18WR5mXNpxAGmnuNPBJHRCwjN98WQ/nTCp2LOzvaKsLXhcrfehmnfkBfkB1ozlL5
61p4IFFaRtc58nJA59o8kYhmh171Oa7jZJ+bPlz6ZJDRh0ljUK3fjsYDJInw9QZA
+Ox8kKk30pwVlgGxEPsKQhW5pWJTQia6lgwOXtFv/5xam4OugF2XZrfSJxmYwaC2
cmkLKtTQg/YgMbp0RbZ4Oi/4Z5oiI3escYV6BjRT0HUJMjZY2CkaLGmspqXefBml
bSQY42clFY2SKYgrMN6dRPyHCeDNHAvfQSkbVtBUPVfyLSt/fsBrlqlpQyhUahKh
c7TRo7vcA5SQpaiwSzx0ZJxBbZwPKqqiUNlrfD3DdEpNs7JSKHbdD28IKFhINBMB
i/5Qqcz3Q4RVdhIqSJtyycWlWIwJoqSoJLGnZNY8rK1tAUxsVPhenAgvjhh6WOnC
lxVi/lxXrtmeel0tZ4KCQtB3qzHbcBkijohpug6YLJp82JbuPdQpM0R8PqlB78Xk
/jbk1v0yn7+Joh8vXfIXo7Qu1oSUYEhLu0oPudg+d0W4pAOJNVH+h+232f9GMlqG
P1mwVnE6Nd59yUx39PWuQ24FZ2xdsPcwWCknHI0qZAe8aMhWh7FDQGfjlU8jMskI
u+9hYJJR/SI1usqVSRG1mrK1gzvnMvco00M2LO7bZuItp621bDP2xkBH5lwISVve
Kcoc1Mhr9+4LErHYhK+GItVxj/v9bYrLXG7icNbUiVG4lKq8lmQgFmktEvgYlXRl
SOebE0rneavBSNSn7tvI+KKGirxe4Wj2hGuICxJyvnZXZLFAoMVujKhmnT5p7JJo
o9TD8WmZfItjf+gdpESlxEwx6Ij9NoNeRzZU1D7BOyAFaYEXvl69EC7vKp7QBKH5
COzEjIhbDFfEfWpTPJujIqi2yVxWA5eR/0SzeAj+bX1yZA26Va1old92fye1eJAy
6hgR4KJCXz21orunTlYSRRjpoGIuf6abEDuc3ivESaz3TMRUnA1AA2IlClYXsT0i
awup6rbMHIuCY9y5UT+okbIshWBvS6g5DRIxFb6ykr0JeSf0EZ5InDB77GMfBQrv
9/nViMDjcOUnGRshVP4KCAfFxtRwLJyaLVCrEMqaObqyzpXsVIX+8rwadXojGxRv
ClsS4y0P90nAtypxVEKGisd6smpS3Q6OR5CXA9/SdB1QbaN/xdkpJAf9Tr7GcWKz
e7v46AqEOml2JPN4eGHeO+erBT+iiv4466pNf7aeFM6n5KyuLnlY1uTlW4GDwXG4
OTjRVH5FJ4H76AHM/afDxL5A+mbwTMNKTgU4IcGV1ez+cbJgiWVyKtNiYu13OESO
QS+vy13ITtSx7Y37Vuo/rR61b+AblDgRFPgQoB9wakPIx+nK/UkourEKrCsEkj/6
lh7iI097kSxgZEE5XvJ2K6PNOrRvC+E1Hv+RbCW/fZMeUgknyazqPw2KjQwkAs1D
4ERZWsd+nIYfSOGV01xHyWoxyJVtcHauUrQSyCWlL39YMeirEgaYZBhjFdUCmm1T
wVxH6cxB5lTDxnoTQOVb3rj1QZYue1fU4tKJpzrH/X1ep7Ed5vB9bV4bbd6A6RWH
NaVLV4B7N2Siyypy0EK+H492uPjChzfSpqaVPCFi1UBc/rKe6+LPvFdl2dZa1etK
2/CRo54AbwOAS2AdN0iot4+gaqIT63u3M+wq8Q662mJ2CPZHyKi/P97hmX0HUTXc
lB4q1sS/iGk1SruCtFgtJAtt9jPzH/sh2kZsRxwytr5AvMZNh94DPHb5Hp3keCs0
SudE9KZ7k3L2T9eFUHLNif44xlWZAKMt2LU7sHYzXFQ46hCVNs+2R9d9MNWKX1ju
sBS1G9+jGwnWoNFAu9LNA73V68DffA9qRaSG4SxgmzSS4GxnIbUOp67nodwCOnsO
eDsA1sUEBIvTShO5ndpbhYrEEGP8z7kZZrMSrn8uRfvydHw6E8yWdhk4b61fc441
u4LY4iDJm0v87GMQFLJJTdloHRaIv/oKSQePvpFlWzk3LlG2MfVqnw4d4F5sGKXz
bRxwG7mxnxUv+CdsfI16mWofGwEXIWAlfC1XDi4rXFzizGTlt5S+txJchIi0kVur
n495a5q9Zvkx4qcB9SeGUwwJyBIMbUDrk/QsNlBi1Sl/tVcJSq1OFJlLAdZZfFkU
vkv3Ajb/UHFxX4CzbIdwoBH9LyHsSlGOsNFt7rVhpyAVDNz9ambNgsmYfzbGGrFX
r4cd5hPTDUITLX6r965cisJBWTaspNU3lTlHmfKZUJ/AKpCtXMv4KXS/bEF29R2p
7yU0HIz/steRgbIqjMuPK4EkvyynOblW6+z0jdmeS8P2k8RoI1TKp9MlWMGPBTK3
gsAYA8z8o7VR73AFtOedJZTEceII8rshoCGkhMjstFcHPZh84oZoTNpdoPsJ3Vsf
XBH6Kp8d6lwcNU4yyHEGhn4crzUvg6aherHchXiHisvP22U8/m1Ztw4bei1n9/br
OsdIY0VrRtxXWsFu1CqfhX5nJdnlf5EePr3HVy+n38RGmB7lHnwAYblyPWY6d0jO
DRSgj8VWuBOr+KfjLvNRDD57Pr2d2fpJXEX0mwXMWO2D75cO9WNsrZnhNW6eROvJ
R1Ab66GeLvirb1NVE3aAycB3kA4fvrrdsANWBNaG3hzWgkmmTl44IcYjxuqYiq/Z
8IpeCIFgdbQC3xbg0Qvo6PzjPsBLwa31/GlpsnRMAc1Gj3hHk3aBFXBdXj1I31l1
jo16AehGB1MhXOEVgRT6mWBIB2SGNuwPawkijHMSc4yUxO+nsFAp8y3/fRBjaXOE
aG0wVIxLrUUE3zSSVrxcA4uXRepP7SWHE2BPt6B70GZqrA65p08/aS0GeJjzVaOg
x3kDvLUKySPq5rBL+xhBQfPAYLBfcytwS0mV4u4ejotPP755dD7p42Z9T8Z/RiPG
jTnEk30tVIYNELRI+uoGYX7Mt3KGuT+bdU4IQ/nafhzOEQ6O+aRG6coF0nNipbSC
62dcJi2vOpVZ0Hk659C/+zVvbgSmatq1I0VJuM0NHgHW5UdQuZqg8r9vvz3O0wfN
LAgLgPTeH7Ws3UP9kR5t0gFBbYl+Pl2qGfEm4NRWQ7eBxV24JJ4iUgbhvZ2yoa4o
7Vt4raDrESxeKcRJ91KKwYJyYJqEtUgkhp7Ynq1fEs1F3VGsHnGN5Z12VxldvW6C
ONhbygdtH1K+sn3vtXmTXz0AvcNa/wtuRRrMgQeDxuo6mRvkZHulDTF9mPNsMxSt
8p0q8IdAHFF7lUJjioLPejb6C+rMM1BpxJ9xeviV0M/5vc1erkFmjERWz7zVDGEv
dawkwsx/6ec9SjoiMqTmLH2fMmjwBcBZAXXX/NpUieMTfTq47jWa1A/Z4Qof3mhK
o9BZBtCOnrYtYm8bZFcKuJidNcOrfMqxCVV30qzGFGzE2/eP+UHQLr6OzaHh+lAl
+GqoB5uG0Oi56QZi3gmjCbhy3GcCafL6h6Nou/0QVaXfN1kzu/3dUFugv8rCrdCN
kKKK9+kdNWTvaz6DDbPibmbVFm4VlJBQ0dEkSAtW1XXdRIzSEWcQq0quY3XGvnRz
m8zHhmz5BUFTVT4F8zVN1nMVth3YbTeZ1MsDLWB3QNndlv/d2wOWt7BYWIDX23OD
Bdui7jRfB/eqCV/RJ1tbJzSEx0/MK0VNiLtGL3XaOiDmVKkcnk6VNf104GQL4nxQ
3hIaeL6Utfcjbf7LI8r3qAY6p+LEbd8x3OOxO0b2v5mJQXG/mku6OZjlr2+dngqn
/pdt16JM02dB4S+wPNkVb+YfGtUnYPl3T6DC8aJd8m/M6+54LBJcYl3a4CpVuUeh
BRCT7MEYTy+fG0X7zIgZNPvSGk9ymBV9Nspr/E0xs7M5bGj/d+lSSWkNaWHnFDsA
yx0byR8RFS0mzVazBQJzyS3cgOb6riB1cby/v+t6z8T6bX1lPHsuzoLEz5K3s5Hz
9GnJPzw/39PUItkTMekrs+hZ24QBMoZv+dpRN77n50lzEhCPhw5vY7N4EJbCTgeC
606NGA+lcQbS+Cv6JcYBat98ZGdLI2e214ZJNZCT+ekit3I4GpoN0PPxIxo+a/rT
EjxfoE1mjy8po8QFvzr2YAk3kkjOOq/jRfyiXaqEzrAGG7+uRhutiuOPPkH5MqQ4
szzHmB3NKlHV1uc7XxJFZYbz9vMWg+xumS/llUMxC62s1kgFRPMxJgx2mn3DCEMp
3qxhivaAR7CBsX1Fl89M7BG2iNd2EqRQ/rfhJfCRyqSg1b34npoKajy6tPpwphV4
loZCCMlVUmUN99MOlGszzMJngpfbbteyeoCrJp/RCwTQab6H+Iv/K4mbK0PcyWJg
/cRiT4at8gwkpuXbvM6NAS+SHS7zREBzPm+IzAb2ADsy1wnSDKmgo4MGBSzp/8IV
yCGNhW5mJudGXhfi3AwRQdfvedASqQIA1ZYIQPLRU5d90VEtrujh6XmZgaO3cFDY
TRWP0byZutm5R7dVzYbHbJKlXa7ZV4khZ8MXw4g8BO29utsjIqp+o7op5ZaiUBxR
zjM5Ybm7LNTAV5A0xscCAf5ODBuIxUbO0AU8XpgFTKHxVH+aOls9j/NtLi6NEqCi
H2l/QAD1QuaA4r+pk5AuaAPpht78x3dZcZ5ceBR69jFCdVYmVaNU45ioaxVvBUL4
dCdmEesm9TkSmE2mVnZGYVHILfpGeXHdUd/P+eHtIAXlprgRQ0Byu1eOKRhC3zYt
GhEclpXM2QodS7qzTrjeza3SHVkkT+z5yzSPTUVJPmSvUmJwzVTL8/9CkORVhr8b
T/bq4Q+yOFq0i40f3Yp5Y6fGuAX76ovz0mF39sqSdqVO2XOfJakfBUhCim4/Odcq
/W8KyfWRvBh6sU8NHjI7KMteS8JrWXJVb7yNdghCcKhe+IVAQqo/GFfA0bikxJbZ
iqPTKc44WDNJfR/h3JD/FysVKOIAgnLDKb5wHHaVX6P1qqz8QAZJfkCVPGSqIqlz
Jo+dTCdA8WlkuTjji6w6uYw3cTRRvA1XcLOTxQEMMGC5MmNNGEa+W9huG18gL2AG
Mv+bYj9r5iYySyON0nxYtnjR+FADNGgqXLB+rn8pRMlnfbe5wg/owTItAq6lAdrh
4RMFt/776rJwEUW568YWwhcG4jeVK+QBjtIpmLN4spxCqvlfjhu6sx0Aeqz2iPMp
SieAhazfjoZm1Y3TINFTan+GpfgzJemOjPCWv6rG/QC5xhcHDdMpTt8rYwV0DOHE
Gbupd1FazO+TysO0ilVLcqKfgizqSDiF1W4DtUevQo+t8M9RbzhBABzCSL+ZOFkg
VZMI0rSkC2YivHvTLXUJQ3tGgN0DyVI/OnGeMVyf7HGd2wlTainQtmaPSMUQsulc
6sbcM4fVTnPFBE6+XW59TBe4OdXs2wSDbCWK+XRYgJYwwiCMz1EmTpL3SmCw1t5I
4PvE2j3iTiz3FFJP1h+APbocAq318EnyMxKQriV6dwJPHKVYCvzDX8O+/Gsm+Xzu
uiYe2sVqNfI3tfSgjafYHG1rLNxyJLH/RiWugfpH1nO10bm6tTtqYNYoNxmsGAWk
oAcSb+WdYQE8Ob7FUc4CBXhOc19yVMSutvytu9YHWebmpQFRinwYri2v37+HN9n3
vCD1OQw49v5EJVQLyiXBXSwvCCoObVECqo7ymVmP3kk2ZeP0hh/WI6jlBYV2AbOc
mXXBRSzT1V6rZHm0uSNc3h/Px4lQiG1TAn1EVI01sC8Ou/1IOt3kRWnRgL0/JRYQ
c2UQnA6Cxx0+177QE6afC8dsBcQmASLxfN/+nbZ8TomZH+YQlcbUiK8WsXPaFKtt
RP1Q1Hhp3T9kcLl7VBOylMh2ZcEdP2g+7k++IHM7CroyRXPRaLZg3REYH7bKgyQ5
c3Knu5NquGIuC1KKphET/Ph9pZWkUPdWBk4UR/VslFp5smtPR7Yar+ybxggBdHYt
IZJ66+iELS6FGO5JxMvPa3jS33TNJAgEh/b1KSFtGVW90UxW52r7kek1WKoguBWA
4LHZYZNEr4exp6DcwL6fjjYuS1ob+pXnvE/Bwl87/iUzHgyNpiwavDYiFF8Bsn3H
DdrJzxYoypkSv9j9QstvVkj7ty9GwHZyBSS3Jwe4m7hLUUdW7kOMXZIJ/lR6bCPx
IqJcbrWSxepRO4m1ugTORNTzqikXrnJKTa+NqQhoKs/VDZ1oJes+a7enXfK+aBHr
THMVHGfenuw447c4REM0ZWweWG5wHOFTQXGQIVzvNm4JGMeD0EdPOSYlNHVLWixj
iZy8T5GSST1AmsHMeBun77ZtdmFC7ap9By3lCMiR3hbQi9GIAEvwuQ5M70/yIcqj
b2mwN3kRY3vkITJc796FO63IBepszFRq1e2hQMZYn/Va+C3baZCuSutLYZ8CjWo2
96Eg4TJpEP9a6S3h6vEKT9IYEcbZ4o7bY/leHAog61ytKyg3NQVFmzGL0F4ecsHd
ZQ3QwkfOzZ2xtMqhn3m1fK2YBSzH3WcmvqXQUDWVPXMSS45tdp1e6gfooNhYDbQ8
X4aDKPXO8qGH+JyHPRBMnu6l+g2UA0VhjFdE2qvS2k267kZ8l6S+yDSEJmdFGkM6
iSFrrNIxT/AFeTXUoC2oOHbKjydhENa8zll99Yu9SFSw4felZm/bNxuLWuCXnenl
K2UdSVW2xF5IuT1XadUbcWFv0JaxwGVBF18KMrMhYsk5lOyUFT7FOwX2denpKQHU
mL41mKnARc/LwqqQDmoDIjQ10dkydyqmzc5qDhHSl2sB0C35UOba0acKIrKkCRhW
wQgn4/gQN8XEPL/m09VWaMUnGJWaOF3fxdKVUhSkI+T4KPwWz97ZR0vaO6JdNBsq
dIz7BFNoYUEPDK2TT85JAjHYaLAht5zHZwMxgVWOK8jmvzU2MAfyXm9UFHefv3Ik
MYdqUKnNzQ6v3nNtrs/NJrLL1xEXleSnZkskiL7Qx2aTwJNXcg24wE1/xM1MY2Fv
R/dfh7FelQQ3aRGexup+EPvkS0DC9yDkJKoU9oVHQb7HCcs2HskzHHik/gddhW/c
9QC3zLavD9kIMAlLNNICSI+YQYkA9h2qtdmw26V+mLvL6GodPAFYQBLBGPLQR19g
zaCNm5ZRM7xyvEl8aU8Ta86zJvSuXDfp8HPcv0Mw8TGo2PfL7JvS8UCzMToleneq
vppQkquVFl8Dl/UAQaH73Hwf5dOBRETYZSR0xxsA8HbY9Mw2vlsFp15bY0rlLYO/
/3EkMdNferBK/yBCxg6vYNI2HYKBlUX+HnRY7LD26oVFlsnOF/F9opW/pTrGwK+a
LTLbWQidq34KXrBYO3PlFQ/uRrFG7doJ4xBte7YY7JH1jjWEG4563KqmTHpWdrrx
uhtabecBqRpD2riNlCd6x9h4ZuJntk1t8fQR6EJ0JJGh6OYqkK5pc8USMvYf0NaC
eubfMRXmsa1NzrjpRa278JDLzRH7R9Fb3wjdHphXtADCoEVSD8Zsg3LeTS9Rh4dU
SluM3sqmNIDYH6GPBe/DNI96Fz2LWcwaEVW+4ElDNC4ADIe6GsEiGmr8ySvvtoGO
pmMaiF9UD1p59sv7ogZ3yacLbkLJCr6YLO8R0pJEpLAtqkPVv9zXhixByZu0Ogwn
6HkpGffX/eRFxVl0RVZ+sAMi5kolecLJe20Wp05zy9KhyGEwaW77SNUcl90LWOxK
Ec3bZCfvhFCqbGhZW4B0A6BZcyi9hqhHSpvqwwWRhjz7PUuRfFA13+BpXNCjhokN
6D7EcNGW30S7j/JTVBBaimFwYKBtzg/Sd29pidteRZ9altC6SkKmzO4Jar71NDA4
KdnmAdYbcanVrsEIhuePy3rHEBcKSMKllMSPyWnyn3t3EvlzMNhcMl3Eix5RRW22
KC7+Vn6qz+C7eAgd1LgwTfyUkHmaKrZiQjsQbia1ocpcYX0dDoRsnblQ1nSuJw8I
J+6UyUT4XK3vQ4IRMd/l4WES0Gj+sgYd+Ema45F948u5fnYpdpXnzmcWvjI5NxWY
1/uiFUWsWtiKFS5GxiE3r6M7FNcb1CyauEcFOwfQl8FCsHBJjMbooD/GChCuuVnw
LpRlYBRtSwItg9h99EXw70FgoTOuCqS1n9aAR3HQwowCh36hbEzXSkewc3endjbm
eonCsfw3BW+0sq9r5o8QPWlAcU/ycpYoYUDXXYtkAqx1mfwlVQM0djgVQOrs6p/O
Uj8b9tneWXP5T2IQnBmIzpinCAHX3QqETQ/aB6NgwQ70xDXcXzi/8HWd3l+mEmGN
ng5yT+Xhm5fLwDepv6cexbOg8vJNMB6z64Os6TYcpfuqQCfJPp4X4NoEuuoTm94a
DLPCIVyLOpd3bl7kfBZxMP8d7zyQEAn3iUS4jLgMSxDCKwmmLNqE2vXtrY7nbg0t
eFDWTxRYfbBE6hAfgACN1+WJtTeOkIn5rWbBa7eOR7oSV1Vbkj9c8qPFZBsFwoqT
nj+MCjv8WjL2WwlcNu+Di/or7OLJd3QMIvjuK01V4WCgW9zLWKqvBakSpWO+E/A+
PQiEgllnSmeODg99TrILR8peLN1nUDSpa1TPgkDssbqBPwvv7jc9OVwIcHmVxDx4
ZEB+hZvsvm4pXBNoFueAGlpew/LFy5nA2OtDd61/hTpihPvXQt0ecpBRFg65AVeE
gpJ0J1HjclEunhXdcgXdCG4E4MbIR8ubHlMBrwU3h2bYcWhOeueMu8xCiyrVUW9K
Hi/qHK3T6oSHiMXaxGE/BW5XNzEK+pyWDnPA90l0jNN7UDcaA5yiso2A4VXrCzS0
TXnoCfEl6IDM3yi0p91CM7xRFzVpvYKYn6bcf3H7HAmN4ciwTrazzZjwoPrmHU0V
02MBwxlbIfLjqakUFvEhyEkXu0egYVXmgdZEcW7hL2aNrlb4iV6/DkfziJDmbKeA
/E/q2C7rdBwWPxwsKV+DnaJthXC2HsazW+EB8ntroSn3nFbbvGpzg6+ce/8vIsLW
ec7eqkNtUUO2V6BOLP21H4v57yF6tdeuDuNrS9rbAKCp+TsWj1Q0WBD/WZd2Dq+m
OAmOuitywR260BnUVXIfoqAJOWyEvP5yb8lsY4A0UNEKwAzN42HAfPLVL6My7I4s
bEdf8B9snuwwbCZ63Rzh9JakMusxyujQJV5OsIN4NrkCdwfu3E27+PvgrAUek2x0
zR5namXmmHQOf3cRpgKp5FkQdQCZhW1lvqmWAuWxo8QsQy6DlAwIlBsNSXgDJV2j
AY/3PE7xfJaqXFxC4slNSYghpSdBlHDoxXXZLuA1K5bp0kj+rBU57AshODhOl9JI
hvgqsulzQ5dltvvaY9fjD5OWM2SAGJjMz6vVMsu5QSzwJaLm3XIoffOWRZWJebVG
Y5dn0j4LRX4OH8ngZOt41KS3y0GhlNt0uZ87YAELihYQsaf/XMSUsn0fbk5sSELV
six/D9MtPlEuECkyburpgYgKeKxxLITm0d3urBcrsmwkrCf54v+OxC146uhATLuH
EYzsae8M9SpofSQAHs96FNoBqZszOkAZWPp34/BSFS8PAQNanuJmgrzf/+kP3TyJ
cY0Gwpli1R3dutFh5O4tG86jWl8hkM4VOGujkMbepy1iP5bE0noxcKFEdiiIu430
4jNGpGYddolpbjsBHqq/cSN64XtuY5YooMRyt9ZzQurEi749y/ibPNHd852XFU6q
uDqCaxiLREq7hgpHn4csZNfVWquBEbgeBVYAf4yQ4A4CoA8Ff9f5zPj8qi4KOf5m
JC3g9jCldQVe7j2p+4O4qMo8b5DQ4xhWiKtfcQgEx1o5C+tEZ4YV5oWCWZtKHSyE
/7q3EnMN6q3tfU2qL8ZzcvfCLZ32YjC2SY5jf5hrmZyQdbZf1nrtaD6Yk+6UoDQm
eVeMhJBSuWOWk2xNhVr4aL+aXXH/16hs6X2U+jkEbSs/sXX5RFKGEP6W4X5YoENb
zSZL9LgrU86unw9Yv4aTMtZp/ADATOEtbIEOgbIyWJgxNLZ1oiCNarzUq6bagpL/
KzCyeCFNM/DlbTlNwVBEUfGwhbtvsTKtD3U1RRPDFuBZFDwM9eBtvT0xY+KFaEmM
Sc/vi0xLsqebto8ZWK9nYuNZ4d1EwQawAyVQK/gAwoFZX9mfQ/ubGUQZnZE5xRGO
LFPgZbosuc6RU+xMXWcnFkAb7gcyx0YZSonw7gtzcx7VtkNlSOPTRn6aXffL61Wg
lk5D1GHb1ar2dddGYgfRgmMyCH2eeqIGl27o1MN82XscRL7LhAL6MY4fjy8fMPY9
NLBMGsRYnBpDvZNQHc1Rytd7tBN5dg/5swKMJr5fUiIaIJXC7RMxy2njPLc6AXkb
Ocr62iC728kIN0hynq9ChZ3pSFXKY1YecLXS4UqVLIHOg+uloW1ynf04x8icZlvt
9Jsx7VdYF4lqvKA0sNWywGmSv2cUBWF+GgDN5q+r4nOOksRjvMkbVn+xk/gIuiJb
Lp5rnwYvywJ5L8kTLHWUZ+wOcMPp3uG46bWfsixV/GNQMIUd2UIpkSbO/vwV8+Cr
iArHDMkbX3U1JNVJSVIeJdh2YXO8LJWc8HIqRmxv54zRORV9V9xYzb/xKkZ/D9bS
G8K1dhoamcuhQHj6gcwbm6G4D88Xxioh16MaQnjLlL1rOqU3tvbWiB8MFr4EVLMA
eRH1h/pal1sgNo5nEdWM2Sd7uX1imdYXuEjXtynUEfN4xdm23qv4gmqqtUcpybhK
s9GA4BE3EQVRAaANXGhUzrAWGuQffmP9GRnCHFK5P5vHSVZMoq++/pDtGBD142TN
VNyb8VDPtgKOsHalhfB9eGAH4Dk3AcmSwyh5zn//g/W+PQyyDVxASNvk2MCGGMTG
a4DDGD9HRVF34MK3iUIsKo4+6C91R/OmiN/XuXZr6cHt0bX+rZojddZhGGSLSN9L
BYohh78TdFfdVxIuMrUaUM6qO8G9AuJ8Hnd5LYX6+lOyeeV/YdYJLnYhqxN3ubYi
629S4U/mryl8Z4yUcqomJu8c7bPtCeZsHQP5Y3XtcEu4OAsXONG+1EKu6CpmVNVU
l/3kazVTWaYB/M0dQxiAEzvPhw2p1K3L5zwZPDTQbRJTfTMT6hPHRF10YtAvwxCe
O5djTzRd8cp5Z9XuuJMM7RgOq+Ri56UJa26Z4JGvG6Qv8eN1hQb0CzF0ztImD/J9
cSuluEpT7CkK2Atbo1pa1MoC8vlNITthgHqcdDOq7WzYVct9KJoZkj+avdEtCHxX
ZLGsFaeMngpCynIT05NppS9NKxtoO48FQJ0ANhppTcxteouRD0DvQ+Sc5I6MqMWt
VK0C/t6aJ6wyKoxVT8SeiX/IaWWNSx6CCHLHeLfH3r08lBbDU99bHpVLTkSLciBi
VwzapQ+3T8Aw9uIEA9rP0hY+XKQW14fmgTvQ7W05R/7S5NqDCSugGULIOS+xtJIl
Osgy5Sucg7kyj/wIpgiTMFI7l3KZ9myGgxNoSocTGy/h6KyaXRzGrRLXaPSDTg5x
AEzdVdChMrRY7kLLEI8gi22nAgATkN3xOnSxfPCzVJm/MNikc6Egl780oX/xOFui
TOfMyMo1Dzr7Tz71EU1ei/T/S/0R7WhiT6Zi/sv93DbfcGtbhnb5IX2tAB6gSNAQ
rKHcmwwXSmtayDnHKTWlehdiD+nQj/Iotw1xzkS7ApRC3WobBDPmvhR2/jitwy/t
sXf4oerM42I//wsLn5kE4o0vwGfJ8GMP5W1frrWXVu9jmd7AMNSe9HCGc8gFP1/R
VBp6T8WYN9Tf6bipaihZLdoBk/6vlLkdxvIjoiqLYv4FsdoQ/G6tOi1lKWkA5oXg
/v/+IOZfGsjluRaDk4YhZ6SRhzVe8eVHDSM3A8t0NDUP/3pbDz4By8oIuKR2HDOU
DDhvTAaekMMFeQ9zCoelz08jVcKzyk2mXIj9TOkxpokFBcRSoFcEWk4/BPiMOZgX
I2txqWB3cmjJOhmeG8PoS5rZP35qEy9YaM3vvdTkyhUeWpxujW6hoSIrR/Emx7/3
GA81lM1tp4vEaFwlJiV25+Pn/nnLE+EF+r6TgCGLWGdsZ2oF9ziWV/88BK9DjVmP
FFEzn/pNw127AlCawyQn7EddtsK19DlgoUw9/IGxcgDJOwd7qqYdbPzBMiPeyNrZ
Vz8Wvm0IcZhkptfuvWkpktKJPjo39JE0FDalRCBCVBi8hMRYdoszUzIBae0SPtSt
KPTwwhCFnFJG7Kvf1rhGgihTLj+Y2clOmB10BgeGFgV9NjijSga1MWg9Q520jbzZ
I2BE9s64JcAMU9o13cTYbWx6qoAYIENHUv9LtlGnFgMTAiBO9bQywV8z2b7rX9eU
W8TO/PhtyWj+TI+TaY5cYZaHDttmr11psuZTF+nEGz2DpAL2v1YnH9v2otHdNYXP
DfwuHJ/85Dojw02Qq/XoAzwX1fiziAMBf2dNMr7cy5ZKxHl6rJbkPXnibHM6/aSL
wrLZacdwYfXPY9iaAlOdIXYiytIgCY8zNBveNlIAXmgHbl/77Yq0g0aRS4IDd/uv
M84s+bv43KmTzPJmKGVMe8cywEbvT0BVEDAdFB1O18goy+WBtheuEVjCltQL9hKk
wPJB5pIf9fe0lenn6yp23unIIrOLI77XCN99PfvGXEVL6MeX9Poy4qMQNxDZQ1E9
g91PSEx075rcYPPEKjw6mvYwwUIYybMB+QDkBeqBaFNg3m+zejro/TUw4oGKu707
KXubYIHREgdqx9czOju09TltU62Lyf1rjd9Lvc02wByChfrMUefyi0f3P78EcogX
x75cnkPrG8ZlMJXrwPEIu+6FPwUbn9H3So2AOOfOLlCNrPNP376MWGrds7gSYYZ7
+ASQ4nW+QRE5/rYLQeFfUTq3JW/kkUPuNZMpGbeREAoHlYjHZlr+Mmr1jlTwt/+g
BN9u0Mdljol2LGe6E4a3UYgb3Y47RM2WB2CxR8pCQlt3Ra3b0gV6aeENweGgBGdD
27thFWRA1GPVF+auZWZVVV+/lOxXtB9g2qQ//1E8aS6jd+3elCcPU3Gf5OS+CCz2
b1BVNATl3TM+adZd5UkeSGh3k0uH8jtsENd0zXpMmQbFmjHnXjEpHvriBArkZtIP
yD3kH4cGsi4nJYGjKqZNdpHtUfcD0pRTgQQHg2UVKdHY8sdOsqacqpfsI43lmxuf
76ifc4CuldyfMItbWDArJm6EkMNERqdFQISteZAvaDNJrw86jn9BbUMBvAdwZ/RW
CmiAXbg5XDSEN7VBHCtitlu1lkv8OFZXLpEJLIOMfjDUKQxcK8WZCpW5STGgHMMR
zYtqic1pB7PENHpY9uN4liC0kZRu4ZUTFNw4pRfyxZFk+tECdBP+MV1M7h1Qwtj2
+wLhDzmN56wU8htUmtu3Pph3QPKoEtpJwIoojaSA5+ciqH0gus83nBAMdb+gMqzz
tRm/Vt6QhqNd5c8mBDjCDpq4e6D677TFCCYHKjenYjzPK1GoL2Z82akPaEdT4MZM
pVvWOoyJcoeR7usXXBSb+YxVgBqYP1l2e6axCq1b91hZz0J64vlsXzvao9uqiz5c
B3PbvXo/7Nx6PuXukKs4SQ8In99krINX/+w3+FX2RDGacyoR7q34yHlTmuvOyo1J
qG8PZmfBHm58DLDr9AHSrDgMyFZ/rzUKc467HMzvI//2ez6IaWOYGoplXYOB9WSZ
I1JYuQle/T9ITj/XVpGSizZeS8J0Jlzy8A5q2Y61nTgNoDMKoqDUY5eLWdpQBJZm
wiSKZrjzRI8uiWeAGwL8Fg9zNpcKwkzxyWNFAL3aL7RI/cJkc/wEYT06Ij/cPxy2
1s3bywRI2DH9q05Ba3Dxmwa1F917+JE6hqALpC6hY+rm6p/abQOdogB22JzXZADK
YT007z0vbwt3KWeNbORCj+Uy8XyH2+5SnJKv3re4w8/c+H79ImZDhQaPE5YXuMPh
lJTJVNAN3BWrvSvKiiMUHpIcVdmhufvvUnvJ+1a8idq4LgjDcxgfLcyWx0mLfZP0
uS2tcVJkEFT664ZUKhkM/YXI0EfckyjNl6KAzB6KB2TjH7eqWzfP321DQK5+Z5Sk
lN5MmhM1HasudZbQYLb92Ds/tdsuoICeMH8OENDTL/ZYc4N0F5r/P7fZ+bmuh72P
Qxz+O7ArHE//hvfvmxZ0zSXJPCQz66ZlAO1FgSSlxKT6BwmEAx6AIwf5RhpNuv5n
jzEgT9ch76fmCt4ymD7AaL0H1vCZtoyTtZprUtkw1M4jf9sIMnN5dTwTZ1Hu1Ad7
m0c5T4+IMZtZ9axBrWRnUOsJTMwKd1CPteQz6fbgy6cwhF/GPpjY4ObSCOAKTwsq
VtcK+NLY+I6JC8bGL3X8ZFBggxcogb1wFaH5ZzVXjJZw28tIL4VAq8/LXRuuy7LR
hIkBG3Fqov7eYT5S99l+rMs27EeZDjw1M6syZyNJwXHq5MCCt7mOELkHFss0hFoD
vszqIR7dTNiWLkyU5RXwD84AAolLpMajYMqOW6mFA0sUND90/ZNK/SMhO9wpQums
m01gyIggHgSGYXZnhK1NIY0bO96oxGp9kEZlfOXju9cPLlywT3RgUFnBeSJudbmU
t6XfkzFUHAFPvVeCtQF51pq7K+MDl/4i2y4BwXNavKjXa6TG0RgcIPbpOAvaKQGt
yMPcgt5O6jE0VtHjnwkGPeI7gHm093ETVBzfkNs02mfLWUk8FYmtkZO+xDnW2rOI
Of2qHsQT0SIDDaDZ8n0ZNV6tYRUUOhBCIqCchTTUoRMb74Xf8ha/7SDgsH/W9yVl
3NCTO89F2uqPA9FxufgR4uLboqbgw4HHHatpxurKY4yXzmSf6pnXu+6swCh0NvtE
u0a+AxoU5C2A0Cc8DrrY6lSQJ5VX43+XCY4x9PQmq6F1JcrTnPo1s8I9jbfZ2NiW
ibyOdhrJoC+HaqKsHzzjjsT83LrtU/MVTnBUobOsSYRe4cMO4qeje+7QFxZ9iuvb
x2XMbysFBhTgBxq90UF6djtT7H1e/zm3Ke5Lnp28QurrUElLkQmwHcExZbRm+2f6
Zya5CC5MjZlKv3d5cW2ORCxEvkckU7GMW76sKinEnsjg7vNpgP8wmKNjwbJ7kqiC
XU8FZN6bsdDeHxC8gYZuUxxqjokadIUEegfK2oJfbEFGM2RK90pztOSjqNMAaKZ4
5FJrT/KmuXShWlQW/t0SsEFtLItJ6m47yiH5xvaA50xeaK2SnC/gNkUBlxnOBTTz
xuVBeRhXzdiTXDdLTZbw1PDsrlOkz83FadtwKODuQ6cew45RxyyfHn65ad9FhqTc
oWDL3HdTp4xDmzZsOuCRV8ToELUPLQ82mf8b3N3N6Z4EwAuqI6oeYNb1m2Thoo15
3wP3k55Q1YeNmYcaIlCZSILTGSbCCPz0GhP2ABqVsNgxpVRBMwLefiDwqPLscL49
ChZTq8ZxIv0rKXazDq2ibZ/yMaERzWsvZmZSAJy+NcsgohukQTKA6dEnczFkN/+O
wJnCrpoRk9ZrffexBpJ2qE3lkuRzw5Sual5KAUiIDrhx3DZ8egQIz6mTfQEakiw+
ZzUyQXwbzRhs9wXqxtM47z23yr7IEIF6kgjL/9WMIckMFqkBieiFvNF62Qhp17Ll
pCTXxdhtCEWcGIQXtNUmpnd/Pla2alf+nvX5amdx7xU/Yf1/38uHPdV6luwAAdbY
ZcpMiB9YpaE2WNL4fIn9K8OosJ9vK7F/x66qw8APZRKL/aJ6paVNbkzI+vu5cawp
tRuZTnRIdy0LG6xCScmIrwy4ZZrqj4vX15RpOnGsKzNr6bdMmVhJdc4j+F8aEj6L
7DLV5gL9gRijoJBldy3MRD7R+hi440szDzpz28mwKmD9xhmaMr7JmtAnrLParVsl
HhKfNcs/0cCljnoTbZOLwIXyWudrXpRRQlQIaoGQQup1FVXAklzVLQFlSdFnByhi
yddevfjZ0L82q/DBT/qsz1WWFbBfUfRTtuR9d1YMNi8voCRiz1DuQeu2xMKMGYbV
oZqtwldf0TGyZYLvgOKzFSTORLNJAkrSi0qpr7+oHfsBdFRTot+MaB/Qc0y8qwC1
oGxG4YdozVZnW8F8yI5hkUaXJNxEbW7YNvDHetCxTx02EPbBsJ/sljaot5Al5hmS
zMazjM6pLvdpm4e7LmzwSoHYXLPk+bCThOv88j9weGT819JkEn+mtmk++BdDIjzT
LMxitiW82Hh+HU1VvV+/9OVc6ffMeqkHAL227MKQOGjHeJoAfVHuYa7HKa3aHlup
PSCTPjw2GU6ElDhERFpNhjKUupTrKrWUm1OzLvGNypO157zSyoMxq2RObvjS7b8C
qGkbvIkkxND849O3Or514jD/3z7uu678LihwsAs4lkbLve5Xa+vVhGX0wuzJQ1Xk
5nGodWhKsOgDd5eRySRh0sezO7i8+NGrbpZlL716cX5yHe7Suh89l3ojan1RY2fL
EBM5B260ezehI8K47baj9TDMY9AndOK2TD0iQO1wvtZE3XrumvWqXL69Ivd0U9OS
f92oZnUs/FZsb0+5/kT0klJ1MFF1jFdjk2FJD/rPpEWhrlD2oxLz+utfl6cJvX8h
6723eANVzk4DeyZRkNHF3KvXzK89fredlk36V6quYoxvd5xuuI+mCC4yT1lnI7xP
5Vdd1S0C5BSTHH/2QDeH5msR+y99FfVGxYtxPAEM0dVscnrhzhWBynzQY9ac3ylt
36MYlZq5DYfqaH3SUXcKjRUQ7/gl7DE8xLCXVQ3PQT+iT156SCJ/3vbAa9ulsZct
bJEQ7ZiW6zu7RsnM4XDGEEZjmMY7GRt7GyDTPxevg9pT45tgdV8w1/j4Pi54A5Uv
Q7tQtjCYjoXHCwTQOwu/f69wPUSIXy7IS9ifZaL7LO64KvcrSGsuJC5yXqg5CJpI
SQ5WYAZk43df7rXh40agF/XEr840Zn2hwKCptJhpyLAKGz++11Gw98bjM1RJMB2G
08wVsrPWko8j4GIQZnRv5VQrguZiZMtQkX+LRirU3LH9+616PWXGqADNceH8lGHe
NU9tHiGLtP5jQ2gksjDChukCgkQvU/Vw6RG0PGIoZoH04TXnhOgzEibQw1D6Si1I
8eXyOJgXSk/DLB0WSReGH1ReNKNb7h4CDYHdb3z+iuG2J4jOzKfDqflWl5SIdQmP
8Aw0EVnRHqf9fv47CLAaoyw27J2gfCTmRb40139UxDNo4TYdcftKbldzU+N/wTS3
OzTyY6Y4gbgnryMHV2ZCP1/JG+zOL7X0OXu0VKTrxfm+OIepwQzQ3JTle3k3IyOM
resT1PFZFevnkHUzT21hza4DIIT932s+F7595/XoayBrYKvPQdVbrJ7Q1M2Qhv7p
ujl3Ytkxu3LAHbOl1FWyUNhzgsZYgYIzM1fT9jQJi1leMBKel9SWIHKiJjFrZL4S
2jOv8W0QcfMiVL62iNhTCOU1Gtc7yre1FobnSLg/KZj8gmSSE0boixogzY2WgM/I
Owolh52TV+dLZBNYGdFYtRw1uZku97/w6BtjUZk7hXvNXFBRvzHbh4Qsg+ZgL0g2
pn95Sj77raatuL5n3v5JA3qnSwHInKufkHo2McoE7mL2kfSl+PKa5YJa9kF9aKy/
EmDrZOMzdCeLnr9aaz89F5/o3XKDerBV2vrCLQIkpEj6C6cr5QpByta1HCZUyywa
PdQbHe98NCEIhFjbTpoXSOH9IFFqugjY9G3AbR4QRozN5faIe0NNrhrm+CKkiIPH
29dc3IAGpIM1vyPPD6Xxq8otYkPu9GoAa+Q2byg6PzvsQDEmdP1Bk1pZaYvAHVpf
v19LDtPiTfkyDqGA4nCbR/0BZ74QD6iPJWM/uYkYhfj6qlBRuLNgX+FEwO8VgrO0
dYprz1GDdPq82J+utHkjNw74s/jPVsKBnrcAYgib6W7zWEOcP3TROF7bMvC+iroW
dEFrYMiVoZmMOxArK+qKajoap2bmdrCdPuo44QK20D+DdljsysuhUmE42TjQzTKJ
XXL/hQp5Yl0ojPaSfjerYExaZWrPL1Cbp0zqfStlUleUe09J2Z3iKSa9XW7KKPQm
nxYD31sbufR0mS8s0GztMZRNqhqltmNN1SPpicJYuFtHnnGYo1d6I2KZ9yiIBP0i
47IaK5J300DtEUlgyaAYaxgDjGYRXoZWr8g2DklPL6mMWUg0Pk6rpYfdZXRR89C+
msZQvchWBXWPkGObRB5WbN2ID5maqFlBJ2xkvdaZbPp4heYzvanIVqyHUub1rrVn
T4sXPH8Q95kDe7idHH4phlSElghfSOZCXOPv1+qSNE5o5G4/XKStmvh8wprLcUH9
b+ZjTk502sY6KFJbyPuPRgVlPagp4djFYLK8xFnalpDExw1OI1CReo1myyOEC/xu
ZPTMbvTDn0tAmvN8XOMHPKhviSXl09Y5YWCBwgS+mHDnDmd9Uc+jz+OGlzMuDd0h
Hbl48dsIKaOIM54iniYMB6EjztScK5x06u9lL3zxh5DyABtgVToYj0a1eMijUVRb
KXVXSjztTGKJv3S/h6tSmDymKnEJ0yPLMp6JCdx+AO3Bclxp8fvtYHzufmg2FiZA
RIhnekMyENDLkltT6RuGu+2qX6niQTft1QQzCrvg14chIMMfDX3BaEiGZarNtVKt
o4X70KsP2SZ4867jR/j4RznESPFjSXEvTWKroGdj3vZMNSQMZg+6lhn4i6IFXCqX
0jl1GmrBUe1C32uhzLlnb9llTFMuMcPbOL2zQZTxmvgptXe+UlO4qru/0WlgVhb4
oxULR/Vcj9VrNfgv5XLyKUm4pYbmjGwvY2otwDyfH778WYJxf+CE/z5aZKSKG9R0
rC2kxkF01BnSgiVHd/yuMVeyoBVkkpC5EzFMUOSkhiBaDIHhL6juQcd5WKWrqw2N
jx5TG1DqPKOi07fNVl8MKrzdZGakjPvEFqeysnuCGrHFHO/VLmSQ4sVGGE5obOZi
l0pgyLzizi0xOSjATdERQrQSJGGycLzEXZDp5h+WgDypiYZSgObaF9FiPcXqQB+a
MFdW+XPiIixuX1D98DhbMRefR/3tuYxx3DPdw2+mmtuEWFK9BCs4AolRmdQfM1bR
wU8icdiHjlyYH9r2peozCvL9X1duWtBkXOLlN59uqVgJZCnKsAQ5kUwnhtIXN5Os
NF456SQ+elPR0syO4ZvLRAh+ct43ClBmNSQU3xOckB8uiLBiNFGpljxkmCBdV1rA
TqeoVv3r3JFpsJ5RaY/A1ES40OsiuYCe+sl4ZEjnoxMsKlfJZ8+bkb0dWQP3HZ+i
jnDZ7r9xVr5hdZL5aZFz+2S/247AKk2a/rK/8W7Ae88jD8LpgRllwwBAIB8PDXbr
SlP64Jy4Ww5SExUUPoxQqD2JWnJ8nsq9GqrI4yHVGUBDRJ9QPdNWAwvMbVa/ucVZ
kzWa4YCylfg1o18NGMGnglyEJa3L7e5dcqgd49VzPOBUn7b9Xva//BQjYUAe0St7
OcFAg42PTRvk7wSpZjnoltuJBmrcgzScAiknw69tXDp8Gke7TfLHXFyrQOLTtOyZ
/HJvsKgTKSP/BSx2jRckkgq7CW+Kd+wy2dTsCanSumWBFlm0LlffTIW8zYx1XQjX
ZZf7nI/kGUz5BopH4Wjg3B1x6ixAp8l0QGNvquzd0hWh4R17mVS/KAWZfmHBr3qB
4yMgxvoZfd066czOQAK1RS6234VhL9sWUEPOVvs32Bu+2A1fcmdaNszn9rRQv9SQ
9F8Kc+H7M6dF+vjcuiWuTDkD/qtdBl5wSKEQDzOWrp7rxr5vr7QIg5jpMBoMWB7a
WtrjBtMiXVOnVXVyemDlfPfjqnUQgpDx7zUh5o/0oSPI6zAM6A5EGADBgpG5x5Gh
pXbW14/VooFSO4tnzrhX3Ci62uoZA7qvPhMw/qMZKw1LtS0L23dvzWHXos0khmch
O0fehpkJ2HyfkTYR6JTVsO0nO8hSSNHay/tZpmo3sHWj4cZqM6aOA2MNy7g6l5rz
VT2aRNV2F6pa0IT0jUiPklfKuAeDjc70+iem9n4faZAVFkGmuBu7jVBwJ4gmmjVP
9zX9Sytauem4B4y1XI95gt95G9OLmO1s69UhKAt4XAFHQT0xN6ByVd8nkyYl63UH
A/fxq5XGGncFPrxdSyGnROBQPs+mGEsmU57qUhDS0rmA7Udl4NAaIVZtPQEXXHwZ
kfpY5CEcLewI1HZcui9rGbezPu7v5rYlZisl2OHL+GJghbWj6m3SDwViXg1PG5an
X30RuH0k0XAaXJwKgIf9kLopRxMkQa34Er1fPZRGvaj9hmwuVI2tclimu6PgKwro
ChvYHZvQFg/9Tf/EcnITSKgeeRo0kWY4E430jBmgYV+NwPz3y19KfaQMXFU08R6r
YYWgJ18Gz1xX9V1ntuLvrGlfTzDF3brY7TMPF4ZKI1DiFVpseb6SsoH4RzldVrjc
IRODhaLQJetF6WQkjXyp4cNKqkJsTR8E8Z2cjgkT4WFxArsivBcyLzJO3z1zZK8x
HycLm1/N9LixeAC50nTtPhsGbA+Ma9KxVMdekpEP0j3zvROVhJ/yRZrfQcmX+6bU
CLw5489Lr8HAsrieFnOWV3LzvssgQnEZcOz5xRUsYwPX15xm38/4jlzYVLwguyiG
lhnbWzy9Mkyf6eu3d0Xr/ZnTImbU2CA+Cz4Spygc/lbrAZpGBRBZypQA1fK4hehC
NHfRMSpaPCfIowkMZLR0ApG3IOLY/BXQAa5awPPwXc9zKcECs0hnb2mNKDEQ0wJM
Eg/yz86rSdO3S+Bj0FRk4qGz7QWfASmKeUaYMe8G5x+3APshUaJX80D8GaFoBuhp
yijCBwldkkabcaYqoJDw1VcvTqiMsE5uKaL+D2q60LGaQHeDqmD7bZeL56Vh2WI0
rWaiybowFsoc9if/aNmUpf9s3RfkxM6HJnHpbUyB75fnO0QnRkozBrxfbTdQgApO
pJxPpEqporVLi90TfN3WF64rBx5P22e3SHiRDpKibC/rjwyi8Yd6S7nPMNz+IiK3
8SrAtpwgxJqgbIU5kmh42xfHqg01Yr0KKAeyxPUIB515bTDViYpLiK7ClzVaV78A
knIibYJQ9Z4GxIOqNvI6bEGUKQfdPgm43L8kQVw6zIeI27sXAjcaA7aVJJk8/H98
TPHFR0MDtZXZfxuYqvqQt/8EnF5PjCVi8VPYCNJoaUXZSSMf2u8M9r5jCbek74YA
PSiv2WETLyuQgRTAthcUv4t2VwRpy2NYbSg5pIR1gdOnPtJm8ZY8q1rryEunn5E0
tXRKTfL3e0awzf4KKp79SlYJ0Vq5J9rfop3xWuqxxqIkK8OKrX91BEeIyhn++lfZ
AteLce0lLsAEsiduAUF15zUwyibraoOTzd/H9GIZ5zBfKSmjWsyUDo9LouaLLqPU
CDlFBoYFp4aSecb98abqWa0zq6eMPV50gN0/mY5QqyEQZ36l7qjnMfJXF3FxMSgb
49fYTX/R8h4HZ6Ad4ddkjtlgZAGyUdJ+bfgIpFG/pFYWzZBow8oLoXmtBUzeUnL5
DrAdbfts77/kA0fc0JCO92HfO0gVIf19+Y/V993hg/DYTiEkotBESdvVAMLTAUDq
FFDiODyUjTU4hLDNjY/XSpJ1kq2klnlipkEkOMVkCZ4Bp/hsn3udVcHjmyhJwsQt
TST+yMW2n5Z5JU9fbWPCuURVEieYnXNEQPkO/b/r8bDoK0dTjZW4X9neB00zB0yQ
qsF4EVIuDNtqaRiGUwRU3Ljc2+8HtrYGNeu+BcWMolYdgHJK+0uHsPqocia+6KFe
QXiqPV2Fzjx9y+mqJT/Zfkdm1rDvZwiVbMAU6mh61mNKC3bQP8pOoQrZW5BhW9CD
wNTwHWUGQv0nLXAS5mNoPwfvRzyp3Jn5X4OayiNWwJJLR+hvci6IXH0T72BgElfD
jRaHXhwFp8leLYrwUS9p+Cp9N+3zp02CnJrjYqph7l8miqueDjhQYwe1hXoBYOjE
n+HxI6gpuGE6A4Yku7Z1zCtG2sy1rudweyjhYmYJWpAPYQROEZw8PwDoAHs82KFr
1KF29JDDuDc0KNprppskwmk+M1YM6ZnLEzL/TcSuHJr8sj2UL4eNBBda9XWi79ov
93/iz8irSaVtrpENFxqBUAGEFozt5AvgRsBCcqau2LO+QW87pn44WP34LgnyBr3G
8wljbP1yTD+UZENSePtaxaJJSlWNmuTa+APqp0IloqTC3aXNfhXsFmc1ey/M/RVP
WjhOUFfzBms5AWe59RhMJgtxJaHIfOy8pJMZn0fsklSmE6gmVqoKbJcVS6k36KSu
2YSEz54TrwSE6TQYkK/bmI9WrruJMKYGGv+hRdoRIT7okQphAz3Zbe7jch2ZG+1J
cXdMEqJsGAoC3p569ACu74Xva6+b5l6I56+R17jYab3dLNaHYvhXf26HzgCFa/G0
Rqbu/TtuqaaQgh7aLMoojU72XiJG34bZ0fPRT1okzAbK4Aq2epDHnGJQwzQrCkFV
53e7Og2AGWTaHT40k0gL1CUYPL3leMwwnqjSsambQTq8lcWUoH/zjhFB/eUnCO18
011a/OgBzlh7Cppv4n1ESrg3ZUjjdRZ89XbiRIt43neU/aCnZbSurVX4kknimzlQ
Y2Knwk31uaIMGTP0IZHsReup4P3FWtUEVtEY6YQ7st8qKGJ+XblaveVGHEESlSXB
w3ahHjipyU4oXePth7slzBn+Fwjdm8KUiL4ePLHtvxmyYERA6QvmcwkWLvBp/GFq
+DuHlCxLMCFVpklSDBvVY8dQdxjtciUlQv3yVJO13eJx/wi1WpI5WtmSvgBahIr0
qWTZ7cqVpyeosuyQhxVj3Gk8axxJT0z8PZDk27l0KyqJVj68swPpfSJLjFw+vb/N
0h+zm4dfW9V3FMXy8ignE7Oa4qcRhWXnJyoPVpDPGzTaNv+BDWyGvBP5xVBfywNR
jC7KpJuGBuFfYhw0GsbxrI8a/isVztZVDv4VVbXQneGHLakqby6HOUUGw/FKS/7t
Qt6mUd69qsFjALENHAkP63+cZbxj/hZ+XEwjhnqUzaaTvLbZL1G8DUjtvgjrOKOm
uLX8M2ljQT8UCVssdrVoVGaXNxlWEhqlSQEo/fmAC2SIPWbemMLsFBPT0qZH+/Q/
ezBL25vQbKrKcEYviScfmmYufIeSAsCq4QuibMCWhUTRuA7MyDBPaGMqvFjYKzHO
XXvfzGFbgNq7DF9p8X1On5fIbtu+jTcExXCwZWHPfmX2cQFyiXZqaTdaNHhrha7i
D1Uw6NmnDVU16cwW6XwCy3wJJIYors6/CQXz0hOb940hz3k9uPj0Rxkj1osyBT4z
/hoDtYCHBygGBRN2KZma8S90svivrTjY89xKEHZwKA82tAeWSo96r6zpNSZPL7mV
6azpdvunICW4AhONiRu0ocm9rS5MyAQd056zFkElKUiTQCU54wMZk697Zu7r29ci
UlMcVziIjPIiTA1aGmlZ8QElKaKfhfI+lsXNz6xG/XxK084enj442MjqVyjegEA9
5Otzu1IfjmQ0acrpFQwRqr0lNLATZUtVRNhl8j1f7zWQLuIophczSyTXTdf9C1E7
wdl+CvvHwhaUuUWNUo7C2Wc/ZjymUT4i2DKwlUDJ72wucZBnt5QiGc1qrTx/fQsP
iaDq4cCv7kVcxTsPH+MgPA/fqrZFr+FP2/59hZTxzrG90E+RRJHcJNgANE14rFru
FC9P7pLwCPFwaWU9acei0ixrTMDLmk/iv441KbhYKYFSfLFXoio2ib8BP/7MhO4x
ecnBvVNfhKeR/kdQGxrB0Gy6tz6OTjwzBa918uebBk1xyLpeg4na5shb6lI5LzO1
OjorqiMdzjCTrdm0H/6NOFK/GVmPJknuZXIYn1XIX8qRrGiMDnBXvwV98B+CddJ8
T8NnceuxW6XJmhv+v2czxZ9uYaDsNs6qKOpAq9MpjOrMCaCzNsMHQgKo7pJpbPit
fchZtcXR1hFk4tHnoEXFZ51QrMle4bX8Sov1jf3LsE/tFYMbITkFwcGODH4A71x0
cXdtrEnQ/tBZ9jr4MkYTRb7DVdZcfjqUyQB4isJlaO6Gwrptds4oU42AkYYqFJcE
vGsd7Ltj40cCReHyxg6UWKpvPsjiisNUZu3P3Zj5Il8cs62+/rhmep1B8ZaNSCeu
RjS6DIXwi+Ts2AsN24+Tc2hjpn3MM9KHMM/M89QMcXGZvJ8C0gXgJbTZWRM84Zf6
7ehkAcbKyjNkhmIEHuewMx7UMYLIvAmvUXK8bd6MJuYNR4E5EmPcNNurNHQxYTBh
SlEi3UPrhMazG0or9g/EsT3LJyi+/hihBgm5fjGS15DCaz398x+MNURG2nJi+tQq
z1fb4LWO2y2nD31V/ubiVFyUC8iBle8ZmjhgwNeUZaO/Y7n9byVqXS6fAhDfen0i
9XsdevCvFSLz529VoEzJdNtEm+uoyi6xss5t2z8CV/YV4sOs+2fuFB+mxagg3f9w
Ket3gywWs1HTiRjqcJ7cKC6Xktli2K4R57J8lNo4+iwHZcXPjh3AnTa6pSuez5ar
+s7IKGl4soHQQDJWlKihoD/mDfy0bmUnYoJ5n73Fz/nB3qxngZcbV15Zp05809Nk
TkbJVfTLzrJccxflJv1ZextKyyvdTPSeZVV3QMKRpk81DPQLvrx1mGCgyuij4og/
fsepvs1/hQ7DEJX8xB9o4bp2MNXcDyGaU0unGBPhDF2WOpFJaQYo4YL8+2VELQRZ
WI/IsBIgd2k+JAaeg+8Pi27U73cdOggc+RueuuE5NzrY70NUwP9KT2f8n/5UG2oP
fGNZr6ODTcFMQKBDII9pTN41i0nkglf69YG3I2je6uI0NB3Y2CojAHllR3vNNkPr
oOc1VahicSNo9CKdsoQP/ycsTt8Xt4EJZnvWOOEUKwCbuxjEIhLWfOqZJTWlYlYb
OHBigG32pSDQgjHbEsyButKxqwcwt/6fHlXMA4Uw3VgMc4AOlV7VIT7CSqx6bjvH
8FipOilKAYyUKGzvpBx4Aa9sX3CRKZ/VEPh0wJIFtMYhAtaEco7ZRPZQgcXc1QRP
+JGQtrM7aXXr4luDvALrDfEd02a33ynw0mn1TOZQFem68IqISYeUiR+/DMoIPoTg
dazA78czE02Lxfn+CJ0cbe0ePdNKMvsVHrHN5sK/vUqBNQAgeNrE2C2NGIWU3X1K
RS1DxPml07ZoXXz77K9H3I5mkj3PN4Tv3kSramgTBt6z5iv4tqShjNVIUCi1yySu
HpTBHRffWMKJHxIB64vPZ9KeTLuBXV8ZxR/CJPXlGU8K7NlTnRqUEelM+UK6mX9Z
2DzbZWMvp6zvqEjg/03NvaoVUWlHZzf+6B/tDH1oQ2+qcetdO66N6aJmdag+XK0N
37bI15rGLb6Xn4fGOLLkhPqSMOA1BrQBT+fLo0JsrXq+EsepOjyLt7jH+91YS+0z
Fx74dMPgYCLrNJuTB+CR+7ljgwXV4jUZ2KIO5RnvfYpPy9Rk2OARO3snEMeTlcpa
UPZ2j2Q+GKefutIZtaS1Im4xT+GUbwCZ8dst1RFjEKxMrw9/s93LmdTdputVVSA6
5m4c7I/iI5J5vqO6F84b4U7ubVtswqG2dD4+veZ4ozTDD588/46K2K8Oh0sLR+Yo
AQhTGHmVbIIscAhgvtJi/g08DW7ZKUdw5vLCRtI9G2cGnm64JgQdJAJ5v+8ml6Xv
i1oBzpoAmEPXEBvHXZcGLf3HUzuuS571LmPyaC1/yRNsVdsKwenMcdG0QEgt0Z7w
pK/7Tyd2JCCRfMwrBJxsq1ppH4xW7NgIbm0nltQ/jbLlcR0BayleJDY+C/Z45Gji
5ctaA8dJqRLvc6wmhqsFxPSFAKUNbhVe8EYpsg4p+yXheKWXrD5Mc1ZCbgKzGARm
if0fBNeoQUGGp2iy4VIJV9fMlzlwq5B0lnPeeIelo13Q/n1/Q/vDsaY7oM392n51
JelfhJfr/uDU4Iqu1P+PlzzG+G8gRHmmOD9Aw4MMnO1Mc1OP+Ysrfy2dBaUJ51nl
Dt2FrvnQ0Joju6GMmXyvKMJXs3GNage8g5rGkzb/CffdD510iFU9zIX0rDqFLqQK
8Yc5BrccquQlJKmIKvBvZISFo5TapoI+O2vWKN4F1HE2hcb5V9JbPEKeeNUxQxBV
rXwWd+firT1yk5vVAmFjMpm9G0MSke5i3/bSP0oOKJlp8a33X4NsQdagn+QzR0lU
1oYK4W2rrc7c3LMlTPk7vcbdSgzFNNQoH+uQ7iTxLZIxaOm8NtrbTBSHbAdQmlZL
iojyL5cs0yrjXrW3UBbQpGg1Rsddk8l630mJ3C1M6hggu20Pbtt7M+1WZM+e5QqQ
0/teOzqU06jJMhb4O/O9ZdHlU3lqIa8pk1bRQQqvBrAbMAT0MEmdsNAEpgKsN4og
B/b+eTk0dk0TgO6LKJ8+TDZbcYV6OD0DS19UfV/9mcX0vm/z43I6NX/HVBbH7Bbw
iv53Lx6/XBOUc6VJdexfi/LuOTBWW2u8iX1ZOA0pezxnvIzsLmDRyr3vhB/R+pNU
m25NG1Vsr8UCtprPChEL/DGbzSOOZlyiths4wbTqs4LOqbf+YLJlQAWzVdiFnIgm
b1N60wx7Q0C/b1x52ctJmJQo6PvYh+ru/ug8wc9+pa/NYXXogLRvCUKJlYZszHmo
mjmqhYHss1mF9SgkkSUcJz6PULlMAM+RZgbBc6DHhaWskxFdjmSTL9EBlInF34wr
JND0uTQSXjBkLjOp0cL2TSwAMArDfLji5WbvH7gpxsRWx0x7l5x9tDh9z2A7V8sC
IiDGFwSekE13HOiQBCK7QmwwSBPKPZAXvCeJD4uxSazUPyFIDbDVwOnApWqFSf1Z
9AlhPfl+fH7nrTOKpikTnpUXIvKgIe51TuKdoUDfk+xjZpCgICcQfWfFhjxleOV/
UTNx8WQaLfkoZIh8gMT9XBcR8X5CRJXKs9fn5lAc3qrnQS9YEYwvzxvqJwa3qduL
FUnQxuD5a+KggKWC0D9hfe5WuPXuTv9gJAujTTib+qoyG1P7xYPNx0wZzIc/lnn9
NQn2RNb4vg7a0MRDoZlb8Nh9dg3OVm8zRpCe8aVeKe30q9MFF9m+nLabwubOxX1v
YZD6OsVRqBhZB+EboNbMBmVWYtk9RhbB6BLyfrDtJ8bK6koMStzZvYMf7/OGT/bm
SLy+TDD8ntlwbUEbmqzfHdRGdOFwazF6bmO1tLqfBBndc44Y0OGvGcl0f4nFCX9W
NzpL4FFowBlcVHLJ98wta8evNYye1jv9Nag4VhAywZBnwlXJQUX/SGFNMtoUfWMV
hqQBZfLPwDmzOfvLyGLGQSjT7CXuX9YEpC4gCPSAA5oPeh60Ft0v8/XUMCyw1fW7
TJIyD3tbJqDAo5VA/Erml2uUrUfJo7tAq9orpkIoped+KihWeLy2SLTe6G5tZlYm
9rQeAWPEBOHFgAlVxxMfoMEPFuqSavJNRlSTySlPIYZbF0JHt32Q4KItnA6ifkSw
uvpHAXt9kDXw6WemfQi+0ydV0J/YBKY/jIiDFuAwt69WdDXj9w6qZAFskEmeT5wC
g+k2OVzr+uqgAfUIw9YKA8Bj3iDrqxYTU6uxqR3si7UK34grKWJwcdtgVoKHbxa6
+E9VISq4yVeu5bEzPvh684bRuMaQwbhIviVC4ulp2qB/C50Bck99IJfEPuNhU1lQ
Jg7ONQUW9l8p0UvQ8Dl1gX+x62K2ULep5RlwciFiFeQgZuqSewgrefKSErJ39uBG
Jyb4Yt60m6gLNNnUpJvG7XSsbZAu5Yp9qYy9ZjQBNv/b6hDnU6Wso23yPYEx0TWu
EhO01ECPceyyHXCQEXq+jZcSUCPZAKD5y7kVaqyHnpRnBJXSwKwE7PLJKH+rg/c1
FLrKPIspNulzrtZy5dNBBPZ1ZumpAx+DdUpqSc8ef4hY9WU6hU5wTGfXf6WRmXMb
IeZg5lNp5dpbVtw8aUapn5oPkl6zjAG0kzEgzTII4E00N1y5fcI5UNz9f7SKTd3b
SSTP3oULmQ+JBqhgTV7KF/pSBlijh9pcVb66eX3OCj1BjOV8sc236tTqpvcF3bRX
c0foPDs1XYeGm1SgAvrIr9XTZS8UjTs4FMUaKJiXUUR5PTOHennUUHqOFjZDF11r
Fc+2wOLLu+fQ/OmC7r4rdP9h1aO1r+eqM+dF8j9/Z68t/geCeNx7qX35VEUbNwL+
TDZYYZpAdsnUJQIcVQFE0VqOvY+RyGpF6ojAsYgd624+V8sqzzVF+G57UF6rmBmt
Oo3rddxDsvUaxgJlvlL3QVEwAVW3Pytzc9DNvV23OIiRRJC+zILnb10L996wBID3
gDLbsxXTxLGGTLN/Wus3ox4vycNP0xYZjpSzObe2rFZyBMK8Wk28XAga24jGQ5jT
PCDiDMGZbDhZCzGhvNsDSTG9smQgYl3jn8av3ukDWE71MyGxf6FJsTtr/faNaqa/
JHxc01MNjSU1XTDr9khrXXYYTPA+eK0jq+kvGHYJwELi+H7xiFMKPxlOq9A4hlIw
hbB4O+jA9dainBTvpMpfFkgM+dtFGVlrOoVATGxzgMDXjDmfY56/H/tOTloviPT/
mxKrhQFG1heEjlhmajzf3FZLnveHfyHb9Xvdn9Fv1iRxAHsJf0UQ30L8M2P3AXMB
PKz8C4p28UCV92W/hfRsRaD/a5Bl5CxIUEO8qLiGQ2rh1bAtVCZkl4fLOvwmOt69
+oKTFf9AGps6H6buu0hbNTW7wSNuZO/uyHf27bzifbtDN1EnpN8cpsQA1bkQ46Iq
G2buHY0K+2ymdAPz2S5K+6T1RKvHGlw321qQOP/jwOUYLhPPQ8H3/QbLRlwjz0p9
I31b1xVtV/Wa5dDHOOPHV8WwfAWMorGlVamfT89I0D/2t96GQrkHzzNrlBL4+ipI
p9DQjtMrshUoCDBUaOJjeYcJp7aRp58nRRVUuuexy8FERksMYsQyvo2E93/Eu84k
I91/040yZYOstDJJKCGPJ4UTQ1QbSJZkxz8lsHhKe2Z+eeeMxSe6dBZ+yE3/THDr
xWe7RdWqhZVe39g/0v6WVocwSUdRrUyF8NWAHZGg8KgHY00SAKKe6yW+MlDn01N8
Xwm/xDwPeSsFx+zANpCZRajlHH0cWGnU6x7FhA+UAcSCNO+5J8bymnQGqHQ3XPn9
epZgtFDzd3ZVGF+CgW3QSkSP50Ify1GnxrI/X/HqJK3158GVYO5crIpKYS+S7lIr
rMz6/HRwD1rjWu4TBeKjRfbs/IsSsg0RxFyX2L61ruyVqea6lRUQyb6L3OENXdie
hxNEbYG3CX8NxCkwQ2qkiBiKtf+7+sRK4UyMtydsK6LhGwn6lzd7I85O5Z3AoqFC
MG4HkT1Ks21Sy7sPB5l/wM1m57RyEcib6siw7cIkXGRSVSylVd6B0IPlei0d7wYg
Di2f7R+55VVaDXMcT0aW0SfXDfanTpDWZiNIdbsvUjiozWSAUtSVZbxMaU2fRHl9
EvhZc8t6JLmifmviM2PveljcJJtMXKmQrdod1xqNoVhNAaNp3Nc+Igj+udkuIMe5
niwKb6hs57ivytBmoAWAurgR1s9xtZYwB/sKOL3fsDdcWv/+WqfjIkAKfNHIFOKI
tS+b0lzJd/pTjGOvGteo0BQB+FTGCSCiMICs9O2LKk8KPrZ7fG25/jIIIqrq/B7l
Fp637rL46jnvKu1tASkGHW7b6Cx0oCbag8Q3ZFcsBxM3vw1K3PpN4sP7NP/1EitX
J95UIZTR9qtSqr3VxU6ugaid3aCx8tEvlbsDAAy1gcU/9ouc+hAYZAaCr989/cDP
PVBFOjmzkyyBAQwcNnKT1sHLMptJsNTuS0qMhhXkcSXoFET3a5zVZ7VCyVMHztUX
PSWzAQJt8pmA1qqDdNnHbePuBVAg2ZFfOQMBJpEYNCUcmddm5zL68GMYkKKHSti+
LU5Vtg0qFj0rzYQ4jmIv2IBG0Ude9B5SJ0fW0oA+JT1f/+SqYxih1IiKK+NOtkf/
l1E9voeq2FXeIkSxm77lsbL1XMZpgxSs3Af9vhBLogP9ID6O0nulCj0DHGYHUnHI
XDQJKAicLUPFXmX/GetQg0A1Bs+pzS36F83u7RyFhvBIKyzLtHXDnlS17oVfYzrM
o4m1eFoZP5lINTN+4Gule2bOQDNC0w3wtvINRoe7pce2iOS/u22tpT9FzZ5FUqGA
Mrt7zGCXVe+FfPmCVTYwIvJt2zOX5wwIcMOlt5eep5Rhh7HkgrGlG1amQYuzq02H
sMy0OBveDiBcE9xzljVQcCzsLp4OdEdXa5qAF4Wi9WYD7nMPIdsd/VVUn+NCsrdC
ApZCfMXXH5tL9Ene/2BUTzSkyTSGBjY0zjlIz4uU/KcxQ3h8JMJ9w6E5rXlGUE8p
V2aBuUiD/3LHIFsaXhMbwg8CRJ429YJ+4kzEFX3r3HZDtMHWML9oeaMMlhdQX0OH
h1EMs/kCU63KFUbRBO34Hdozr5WQ5izCwMXww0n6N7eXPzP3qCA+EULlOCp6ZfKo
kj3h03lpW8xz0wdg4Ic6rlxnCBbYY5/CNpH3Glwe7ZN16e1vENmpTqT8FXKuHxOr
wsNx3tmMoQ1+qQNUUAOS9yhmjE8cLvpyy1N52watpurvxQ8mkn3tvQM8T8OIYoB0
r2hZdjkGMoNIDWInErdqiUCHF/YGoUZsgZ1HAL1iMhUADUhuJ73Tcwk9CmKaN50+
khoZp4OCbB/2AX/ktf1GZmhf4Az2Xd0pNOs+5LGgOtayFwRrqqFcL58lxBE6HMGq
WkFxahYAyLOWkFv/b1+HKnB+2MuPorCNIQMyV/72KX3rWeMLyJ9fzPkKWvmYpDmF
GSjlzBkRVJf4RNauTDToYS7GTKAdjmAw9/+Peyzu/iEQBxpUDXdVPThALd6Ls5kE
mMC+j7+tp5lp9vMiYAwRRXhBCeuEPa3yiDm5pjN3CKhRXS8krWcHAX4HFaYgojyn
GSd8QnTxp0uo0kHbewLKiPHylK0s0c8PrgTUzLBBVHAl3YIPxQMKC6yFl0C+3vwh
8MaR2yY+/++OwQixPRWn06QgYXbiT2maXoAB9uZTQl2eu3fBb3z/EbrRbRBQ4D+N
0Nj2GFLGKdbeXiCsWDgxCww0H8RaWXkEOYtK8Wg4wflq/MWmLP49p1B/8+QSeac3
6REZIXuC976OdAcStnkvec/ihsf60Nudj/qd3RAIVjynlUQqY6iSMFhFuvgsE30k
PcJuPQ4tdzWWF/1aX2Cu+w0cEYhV+wjBas9LVG5p/OFKnMQtjMzCuUZj4y8cfW+X
fW0DafH6wM0JhC59sAcgFs04y/JEvBdUZqSy+6+TXIhl2oI4FOMaTM0MQCSiBq54
zcyFKWuge5HQ3H1TKhXwwaN96f6jKdvdOXXutopSm74nKVwbMKb4lTjwghDfXvR+
RnOBhDB+ov1JDNyovf8h2IN33kxaRempaVBRcbp9YnYptOuAvJE/OxXusf8FBobD
BXJfYt0nr44LMAvQIFhG5fnnq26SyJ0ulvQOlH+H9uxBXWlKgCYHiifBpNSGsKQU
unskfwAgwUogtjRXnd/PZ6mqL7Ou8Jlk+H2ZpOmAlbpFZyZDt1d51X54AAwCrENX
KB3Tu4U40vfzHyGEpGSRHuyvWsL4c/hCojfb5j/BjV6q5wrAmBgfC/3iAeTo9s+o
gOTU0DLVs3LIXuRiHTBhvIuB6OpZqGLdUt20dNWIDwwzfUdZZFJy2w69pCKDs8cW
h+MGdvrbpJNSHkA3/8qWl7GIvp3toQphnD0YWTxfGSVTlRi08tfXQmFY6WMarsJu
DD1dc5GC734Z0g7Bt+YhjxxbW5lSuUrrGOrutLh3x8WhstxXubjNwPhqkZ9iKSLU
1oj5bQPZ9tuxoYtewMeF7u3vYJhQ1l2H5hXoXAcjU1aYWyZcfcN/gcn0WEPdafKX
hZ5GV/WE+2AbHh+3p2RFrB8Ot+VPDS8cYpQXWar75btjP7ur2xB9fQPZMWaPcG/6
AkAhar/qiN3U3KFbIO3xdjtoEpPcKY4myFTnL5t4yhORKwmRykeRcjYr+lMZXP2C
RUgVNpc69lhRIq6pk4VKO1/Wt6SCxMI6HV+52FJGVHbLFLAXeHBv8FFOzRmnw6Cn
m9R5OmKA9oUQdBz0n/zTUzn3Np/opfAgzlZcfAZGxIDN9SqqIiaNGJ5UFXqxEpPF
Nk6LUOx2kciTa++VwX1X6bb3U51C+Ks8kBaSEQpw/dQqmHWpQ1h30WbTfGilxc6/
Xf+NT0MV2hzsUegLFuLu8/g8tR/ItGKWNdMrOlQBWbZ0XvY3vPJbRrzkHLjh++Uu
DJ6hfaRkkvVKySap4mkCvl6YL7UqOVnhn7QUH7Q2wWIOgO5RLl0C2XVtvvrh35fG
ASTNVZKDnOGku73CtAXE5tM7VZaffu7zmQhYcJuRBvfR0Xbdr8ePe7Upi6AiHUyQ
+OXYZxkxhaYeyYTZb6pQOJFVs0bsF0PgNcVrsxqQXjvy5Xp6YyjVf4eGPEAEk77y
F4CPwuj9xPE8/66H+HUITIKuORpbibBoWRxPMACjKiPb9Y1IdBNnD3/8sX0AMkom
nLkeRrGknPn5R9LZwFcxZ3qDyX3mCLvTSBrq61SOebI1Rt3wA9w0EiwLI262Blq9
nilZRdEeZneWxkO8A1AL4/eHP9yx/SyIzuX6zbxZD5XhWIlY0BaWoC3huRM2IqZu
U+yTFpfk7Bi4Ovf3klbhFUVeJ9Woem1ycfw0cf81svhaswtKpE9yLTQE+3hKbTWW
DKGAvYrUeVKeMOqjvmtMt4SUy9xyTYssA/ilBSJ7nixPIYHamS8xBIgUMzZtILTN
TzmGIKdvFeRw/EhmWd3Drhn/zv9vkY82IB32KrUKna50L/z5x6oAc9xrMbYRekMI
gy9Yuk+tcp6h0LsipjaVAhX+4j20jCA78Dgoc/C293ekRp7jMhPSfHja3WOvHMFI
duCSuJTUN1SD1yVWpLDXbvk51xEGZdunJ1CbjEflY4d5iJ/u0H5O5bp3fdsZkhxI
05bwSvW05NfrS9mJr9E6Om0BGGmz9g6vRDm0ZPU0r+eDlN9YcQb8Hxn9KyZVgsSr
eYllmS4+TbFzGgPVtl14zMOc1WgAFV9wOOXv/Xpzt/aTAjqnTQSE3F28cc+zw5nu
vrpcppoJfObHhrD70ySggrc5Vr5HwfCnXXlI2U+vZtoJhJ47R83KPna9xhvSqy/7
4yghGs1kroAVHqvsmNa2iy+2iboqjJrSIfej7EZUXgA3N496Bs/xQNCrl2zboLBm
6wugA8y61VZmLK58POPXyfRyCimYV4UkXdBsQ6bdcwVnaTQtuDH0FmFWrWYfCsfH
7ViowBb0mYyDYpHQ4zzvVly4hBP7j2TOq7HWLOhWrmHnFBRAQFAZrqjwVMPkSmgu
sVdTNzEH+M7B5kYAAEp3osBp5gOMArtOyYLlJfZzPiyL3locjTqFrahwGgWF05mM
lPuO3qjrTJgWaYjttXG3Iyfc16ErVPNTQ1ns8dT01/cm8aiCCEwyBWCBPSEQh7sM
Zxmmijmzg7Nk6LjEUf5QkJ5zIYK+/12Z+eJHBdwScDPKJ01NfWoasxwzgqt/3voa
ej2aGIa3BYVgWAJY3YUBFe5DnOoOvcEjtyp+eDQjtBs1CK35+aQOSTuTa3RWkC8r
gGqGdve2P+slKX0JVZSSatZ34UOlJhAb3R+btojZu2if5UK5FC+UjdMZRc0E8Ynd
NKFcBuXPce3dvlqovXVTnzkV5GDGWbsXxWBjP40LXZA6qDNLUSeznwEsGbxaN+PT
zwuJ5WUXFmxUtmMTRluYTOEs8U/L6Zb2t3sJG6bynF48G+d5SLBe8ym6gJa2XKJD
PTcRZeq2/nk93nkp031VCZsag+BQtXKAIsVi3tBPauqhI6EOiyPfOxE+N7hSfXqg
5EMvfmLkSPRsn3z3N+mrgbAtoKIxp1Lxj2RgeZTS0R5RQOH4gLoIcB2eQaj/wFIk
Gy2uvHBx3XfNNZOroRO0j/xCaqooXkMODC6wHI6e9dvR2xHt831BchVNg4kSFQXp
MoJ6ndD1gZODEKXgkLdMf4oHTGLcbKmoe9Q3nKKh6IVSsiYvv5O13XPE3ivMy3l9
wKUVGLwd0MvvcmzYZb+JRWHweNdsdQRd2buAJOamnV8Is10uXz9UNcoU7DU8G9eM
EB5FIXlYBtUjZTUOC6FWT9Og+83NA2ahrW2K3+aLbJxOdHQ9H2ZWaYXpQ5u5lWQS
MIgXmDw41HTB5VcGjAkLtKB3dFgv7sEsL/qdYigFbPwONQorBmnRjD/CnWg0NmPI
YPGaz7XCJHMa+d9j6rEkKD08pa6XmzaTEcdq9mpDIpCm8IvEV1WOz1yt6Kdqdwzr
GssrdcXK2I54aM+dcgMjl2dqD7UK3577O4mgt9bewTyjVQML61Bd8Rzfh9EDskyi
Brl3R5At5z+zKo6maboOHh13KOJVwk08k9uaHD7bypcVjOIILfwNP+0bzoZr0zLr
ljkyRy6OyN5cFg8us6haRu+K+dEC8a6PnN40gmfLZECfZJoC+w3S5fCnYkbEolS4
bIo42+Q+4c8qEANlL2B+UV58fFnn5mleIx97eaKVXmBGl8BbiDqK9lXfI6FdjbH9
tyOiMosIRw9Y+gsvkVaKnqB6+6U/QygCsw18wMD6HFSDIW/lNc8k9qPUEMhZGpLC
Oxa/wrusYRllBoYD4vXRP2yZT6EeI+VzsSY4CpfLDTGWXHQPTtBg8YoWunE4Kuns
wr4qxAEywOjF4NN0AtBBeYTziwT1fptdQbbb3QfmP6F6CULoi7ZrzASYNaqHwBCx
mHEwu8NoYmFQ1h/tub7MpoizJc+XWy9Wl5lJRG9ukQQ37eGbfFCkIRk1nI2z8xYk
DJMz13E78VQHswQWwEjjArYf89y3GUwus6/dm1qBJRl/z4vasvvNmFaefKzX1brG
Qn4Qc0EQByf7aU/Q0NWz49WMl60iR93YTCr5Gs8CUvWb4Ay4lN7G1vqgEUh+DOH7
hyR2sgfZMqB+kkXtx/jJ8K7KCFDOEhSAbIUuw5eCJmHX2akJeZSoTUiQks7CjQeZ
QrfrAjAD/kNz3kca4oMUlIgc723v+yWFmEIWjvEayheae6bHsctooExDdpG1sUvH
hF43D531W0yjOspecf358x7bLQ+nKY9WZczt04ttUPoyamDfM5qI6/CFx5N3iNo7
VesO7TCjp2IcCqDHUSuSTugYM1b3mCBnXJZmUNJtr9TD97QdEF9LVsq99oJJ6gZi
GLiyy8EwtBdT72Pj9npiMfd+HZLI1X2U7y53QFU7Fky/DYz/mgVrVHQ3c6Eb5ZdZ
EE5OFkwd+PMjFct/IkLP7hjP8XxELnfXSak9k/KSmj34fbF3Pt/5ne+Ze0ggtEZn
Ji/y6qPE0eTEv12rzq4vCH69JpIm5EckrhyGUr1AC6YA/7xZAbF8N30z8Fdk9hyX
DjQGnePTtL3NXuEwc9IzRVHUYg5Oy4nL7rj3ozQW+Otwr2zTz+EFYNm3ZHDdgWvz
+FGcFY6YFa0esQr9OfWGHJnGL+8JUrCwLt4pVrA39sFzpryqpGVUcqQsa1oQzcmI
rU9yLPr6FkgXQxCf6DEuvItFd/Izt923KyagI3E22Bv5C9S12ACFIMpwUWSiSX8q
G4rw1I90FlEdXnLYwO0ZWAaAqLvFdxsPAepj+oZDcRviN1wOKSDM5OCZUQBnysKU
mFvOx7X8o899IEbQ11jRb4XR2tXRJlZzwhJvOb28HpRdkRd+Oxp8u73ay9jdOqp7
hHUJb3mbZ3adav8aHAFbpSQgJrwXMPGlAlOFw7bcoPXYDDgL/rop6w5DoWEQ0uQW
tbvxAE9RDtCrooDyePYeqJpmm1Qyc9vNJyXapz2etFfFvbJXB1GnBzOc+Sy7wB0V
Y8JUWBC2cHcXpPdw5/z7UZZBx6xkukGCs1kgj5YrG9Q3cQ4kygMAAxiKq6GJPAfQ
j/VqOR18lyH9k84Rqo6waK3cmghqRGYgjgpi2PxfoH0tO24u51Fi8dHlQUy0fEmL
QNb6sxXk3E6DyyBPfICNyg58SqpdeFU4Dwpz3TvyLhqjmVfBkMkGPdSmwlIwtLQh
rem2sxALNZTDCbERkbGfqujv74jR8KCQ8z1cWVpg9vLmWx6GEnUCLe6A9VROMHlg
hlHa+U/62oZ5Yt4EEdw6yRTJD3CyYR4adoIot4YxRm7xY8MtEPdmfcAQz1v73RB1
R/4KYLVlUkTiEHoNJTaVvt26+Pa0G1DCtq4Hk6mTO4FSOhFwMab0fpHQGo2y2wgl
ol7estR/NoajkdGKclzDwuos2a1Nx4PgSuubnA/VvpL+ZmXfcLw+7cHV6SQ1R/Mu
1x2lScutJGtZLNxm6IlB3le1UAmpnAwTLF2BiorInGnaP1Mj+mmUhXunjf2OlcDc
kd7KFVUGmPfidXMIDh+3hx6hnJTwkS/hl3HABAnykYK3qRQdGRkeRUmw3pR6sOFM
OiT+P4rYDFKHKJGWUZn6h+BT0nwWoFsN9SW+isI70fkCh75b4VA9DEtn0tAOhYoD
Jen4PdLQFxOvZbv1zyNa6dpTHtKH3+0yVK0hlSCHp3zgV6IgtStkR9c8zCZTvOFI
HDs6hV/mThISsoViNqYQLXWqnnUS9fSkXvZOdvvwL518TXbZhsMp17VGY8JAbsSU
MRMqyXta1/IkfiNT1hCZklniRtz9tdkDIFAMkUNRX9FJaUWyCZVSjSIUwrbSO7tN
54+YUGHBg+pq+ONlaVqgJt2F3/QCczMgDYo7X2+rulWtxsdesSHNcBaisxJjyVu5
vwoJUsqfP5xcI3BB+Rs5wnpPg+Hyd9oH6y78JrmuzoqoLJUaWycKsvkkMtmpVU1L
NQ0DSLYqWjDfLBukdq3gwUfAxtugM3xenGpHWtc2fC4unSqjyHoykEVkKBe846Vr
jknLU4Mbkzui29uHAnwm+PYZ87sBWHI/NNhD/K0jkG/qB3J+ZhSix88wkCywsEWw
P2igqAkqj77I7MhQBxft1yFspxIeICS35gSjQM2DkCSNj9INmKcD1FaB/HW/+wts
ntn9e5zOG8R/HrdA3L8FN5J9odsYrQ/Z+jmlarTWHim/1S7TjfHT/YqMU+gk9VD9
hAwZ51jpAUpbVo4CdCeEa5cYlMPBGAZIIYG0bTgCNjNUnuQ3/yyepERGwYsEW4fH
LyoOct+9SUzm+qaAAlq4IRWzirJkrdclqv0RDDzHLpo0RsZaZJwsgvTYCbagOHsN
NReGMWO2njBwmQPZbWJbbE7oIyBugv1gDUgo6QRvrbBL+NYE9OUEdoy0bMvOgn9d
fINd3+qiQLsKgwTLqb/eAxkQOV9SMnFEAe9iVtv5SCLqEld4ax3WxUBg0O2VCKLU
pZdB6bn+uxrG2wlTA3f4XoM2eB9dkncci9IPbG/45pTFYgKkZVyA02EhdgIIBVnw
iEHmLVBsSEWB+fC1dGmPPdL9C0Y9ZKSO3PyNqh1Oa1BkgjBfuyJU6P8qvi3defZU
PaEGlFoGIZP5nTc38s4msGsTOAequQNaFpQ/svYLjBmTanY0Pco5mFmzQBX8Yqhi
4eXHOwASQElEUdqlBCpcBiDLNAiSMPz6STNwhBSYfHUQVX7zc7zMK9WKDH7wUeqe
gxleL8Nyk5dWfm4v/1uUoV2ZVFgnCHDFoZy9CeH/8ZSo7y47PheW8UbDrdVOIsVM
JOB14T40oVtrQOmQ8F3dYos4fEi/2ZSpMK6AqtY00dHgQApF53xI1Tu+pPrQbcBT
DBOkZOuchzKiEDoNdJgv7bzh3rCoGYUH+45xERX0tlPF2Ae/74pefZ9Fvgu4qKrY
Hpxca3LSIgV2ClPSy/JllBAkQJBNTI9EDOmJyRk7HEi0i85X16pTnkQ1WmOFEwtm
PaHkVQUYsIXEdkMhQGUR7RYN0lhoxDKFmx/rrG4iYqBYcpXZ+6nrpMGrDeNWZIUl
oLw4HJc7S/1gXiFGW5peUcRNz4YmGKhgUIud5rLWiNRItOHxaZByFu8psuWUk5ft
LYvz4QJhmYOGcg0fzQmFeaY0w03A4gIhbyAYajZa2lu7R/aFuD+GrQx/ZaYK5yT9
Vdh7dDMHOeNw/VrJV06nL8b81J1kEfvEXQeSjcXQT+6dx1DR/m434jkZyyt8fwdc
eYXBz/CMbPpAJ+lAQMLzehQzjzVxljN7sjIrDL9ce6ZXDBLxDHymRW8jKQNHJK6g
s4O+g80c+9tlQZZPL1rn8SkrhLBPAdGgEcNMSADdAsBVeNkoPeY5zcoIPO5PAc1H
yyDofOLZAB62lyhXQiGWtFut0d4pDnUaSyF/+/VWIQ8Tl4PEcfPva944l2IKzwWW
ot0gNF/7oR7s8D99hfaUuvvgJRoPBaYc8aNp4siX7O5jaQuMn+INy5aCV8m3A/i0
cIxbXc6T8+FAapBeP/PHEYQMbBiYsei7E5kaC15GdkpfrPje/37FqN50lsYVPPts
CRoihp8nzhhUNcpD4QE/o+k0pn3kYiXd/Ck35iE2fOuhSLXVxuu+NHFVCgpKZUNt
jpRteaIteOdij5mqFtKJNzYpNPv6N5F/y03EUrWj/9J22f8eMOewgb+5zQY2Lq18
Wefy6Fxe/LYEketbID+BiUXhRayVMjRsEfKolmkNJsA198xJhUcjlPR5wJxFn9We
E9WWx6IyfwsSaHEBUtVVmLHvHSimGa81QN4h40JTAyRTjnoqAiF1BEQQ6UPSeElz
iNl/5jU98nQoXpPTk+pEJwUpsNMX9Zs6db98MQQrh020P8f+cYNyyo1rOFjOve/Z
BejPc08Ngo+7NUi5BQ5JmU7uvm/Z5VMwkeLzVajm+sPTaTgymwfcdjaO42r3fTJb
Zcxk+KN8/riUmtBWY+NCPbv3vphYohPlFOf1r+rReAcHdr4goKUVT8SDKtAVVQY+
6g8o/ktsiFhAUbYRdPLOggqYLykIrNPg1UueNPn0FjSH6Iih48THzWtId4BDCjVw
UbWDpoL+f0xeoLUISczukv7tOi2bAzTcD1pkPjf/joIh8TsVeKoOcK++/NLB/1HO
thxFJ64XCQoLGERJ+WBPtl0R7xz3XnX8/iQ7XxWCpz7cfLTeF679zUQyRRuqfFo6
9sDhb6nO/BFfSOliH1ffqnNzDzXt4lgivxPx9lTSbSAqQgyAV7ObJKVtteleQt9/
8I9Ci+x72KtxDtLIi/kyPkeXGa77A7a356sb4g8bX6kitWkto7hchE9zfZAvjFfR
IuU/V8w8pKYSx0bkOWoc+RbzpmZuRUriNb6h8Ij3q6GByXprbLCJgYDYO69Nz4fs
OWauyNZhzpFq0LRDwPjqUBF1GG4TFlmS94uuZoAPrcuMdSYIvHF9qxcdgTIRrg26
UV7JbqkCdWADCy4lxRgCx/6YcWheoq2F10dJH0onAZZXBwzt9cRjyA3IjrMOQnRk
z+9S2dNoV0J4x/EoysKC6L29oaevEKHSLnfLUjELmQGA+DR1k9DuYKFF3QDNFlVt
0EDdsRiWjwxoLez7vouOVXqTUlf2Uw5Hmy69FGlzZkW/IcLZoguTGimuz+IWQvCE
wnF90WxiE+SLMBZ16iIw+14Fw96PV0RuPPUtdey0on/wFfuz5sAf9/Zf7LFnAL18
ITh/PUmsx5Q3ElAf93V+lMq4Iv4UWYAPiVEFaQV7bEaLxu6T+ECtE4PWtBUVNg0l
cOQ5V+j4quF5P4fPh73qvPqv87gOL8sBIESXwH05t0aR4OZvuUjktWqbpSXHxKVb
LsEQnsZ32cbSuBMtc6dCZzAwDhbneIIh/viGN7T/+UFm2Hy8GYmWVv/zfh2I6oJ/
y3osrBoopkGYCMLrCaC2hCEnLFdKzNd4xdr/wVjBsnKdEahR4BnG0m2/CMAmTWkH
Q6yYSDXHkkb7mIVYClErXrvxrzuzYzEIql9mLIPNUkKwFQkm//cHdcCZ+7vXqMPl
XyFa66+WMHArN8Fc8KdceJAYF+m+3W0cre6sQF0hzpKIf/2iinyjRzWTWiIt87bi
uM+ktqBU1dkgXbyLFeu9XSoQSKxWSTwHCs9yApflLPrpmjBQVMgGiQr25qt7K8Jy
1am10le4/XkSxOILDynnr9NGaFBWKnHvkrL5mjNr3hwZr/DpDccqEW5MDhq2eKps
GF60o6FQ5fLEDvkRUeefG/c49fkGXcjgQHx2gXmnGuIG0p7Dg1FoSeefNgTKe5tB
YCSpKjhePLljOCkno+XxnqTGdeE57a5hod73Sriov5DuMZTrKSSJwCpqGCcyngOt
qoqSI6R776/0moKiE72r3nW0L/0bkut2VdwZdKEoOtBirG15P9xOTR44VjkZ6sRp
6e7u1pyi261pIAEVYRiFI/HMOEVJElC5nyKhp5rp914fm8v2JSofmJTIMwRXHG7w
cVqaKYkRKFAA6XddNFuWGkcLWkAF0JD7jpTnVbkQUs9dE8KFBFYN2heYQLAcU52R
j2EzbelUQkMUFX/azP2Ln7h7bpHd1Z6jBl8AZF/tTPV/7Fqkz0hvm/3vz1SGzo/k
Rkbf/gNI9dJH0oaPDtLS05EKFt0v8KkxYPXC4dAQEvLDG/5hgmIFbO/PzVRjYQPe
2W/IaRyGNGHN+YDX/QZcwArS7z/rA0UsKj5h3f/cn8tmTLffwxM+ylZpLUIUz3Kd
jBIZdtsLjBaHBdAU/k0Rs9AXFmM1gWskEU9RoTk/IydZs8gnyLiD2FDdeMsbaqXw
v5lokPLddAcwCFT6clfAn9+YwX+XiuOLLC14g9h/p+3uC2uEmEAXC8kniWuWjV1k
2O8QZTRXi13daf8CWriNp6QG17YLIl50THK9Oxv8U8TdqP6iAX8BRfOmM8eIRFiz
DIw8RsJ5r00lMa1Iv4oNmLDuqRdNeHKkwEWaW2KeUS5/Ai8ceoauxrPVnky02+8O
42Rh+2EBFnaxTWzYwmkx1ET/5VTgcytPgPrJlJZxNZxTdRNtwPXVOzvKb5F2vyK5
siyShZh5gbDOpSd/ghhkZG6NOyFgI4XbiJq+HdMBGpA2kDgpVIBqd+XSe047lppd
Sfmo5XQHYodJTBk//ZhtItZA7slImt+FdSmE7TLHk4pWKZ8A62mIVF8/nBoXa8YL
akNpuMXIVoEN3Sirc1Ma0M6dR+UBXq+/VuBAHEzYHvJn2vGTQrGAEIuVvhaV6CK/
TmEnb4Wjz5wX/iIkuD/mKnHmZGXK1XLVJrgsSR4KDKoi6/8nHW6PnJcZQPYdIOIr
WiTHNVQp0ILlO/5/02SIvKLr3OuudQqQ6d16WQVm8iK6kAfLkK7HotmHukjbhDWL
ipuIDfWDVzrO6+IHzvEdpuy1lrKb6WgGrv7dST6nX2CFGDhe8uV9Zr7bXkVnT9yE
HGbUnnARp10dAmd/HOz44sLOC7xsoCEW66pZPr9FXBDIA9nLnHGgJwM5Raiz5llZ
Ykga2FkDXP70O3gkDH7X5tmUSqpyt8Xtd1WmpWeu3YAtiowQbI/cJt2ohCML30ae
CJ91r0MDBDU91TehJcMho2PMeEjCQ4U07nFBVFk/RAiNav9BdguvH62TvFGkFkKU
EsmMzsGhoaCUxB2I8gCFYB+oDpN0XuWh0Exlt8eSFihMYZtGtWnvzXrmEJyQw/nl
SO1rdr6hIk6JAkHZ5KMKYQVDe/DH+xkgPPMjW13UafUCsaMHjnjgKabiRtcrtb33
KyGbbRblTITBalhPW+rgis8GVYAvMXAocCPC272wc1Ilrmbw8RnhnkU7F/43ghOy
6BEpNsxeCJn9KtCzr65Mx3Kg3dBN8S6aphXCH0nuYnddvtlHvJeUzEuy/AcU/M32
VfYA788fTeNFFlm5kKL6LcNO8e/SHQCFwHSauf3vT9/36YBL491Ym9ARIfMCYu9j
RsdNWDlTtwNIRa+cm367qf5w03agMLlQtMi9vi6LiNNSzneJ+RJ5GNLTptIogGkT
N86l1t3BUm8P7Wo06kgq5Cz8aamCEUcawaul3pJTqWe7VAx4EvpAxNKJoP25CRZq
Sj6JOmgyPugBMxsXmwhyk368kzozmcRcokA55Mqfwl/aAmJLnrsgKvfwQaR1yNvY
WyTeEtfn3lAbZhEYq3H2RTJAghq9ctDbqkRUoX51+zXYMihHainZMelYVlHq+f4w
WskWIOszlC7wPoSOXPYS6mXR6+XyMhEdO/xq0LNHX96rDcnXllzGlssnOWb1bntF
EycW7Ih2UEvU8RTJgUzsemK4yJTLnOcIHp0pcrPh0UozJ+LN1vPQ37Dwmmsd8zrk
ZIR/77+i569J3P2PP6fPL6PjyUloUT0Kq8uI4Ip/yNv5WGXtwkxg+oZgoB4Enl4O
Lb0+aGruUYNw1GSYGqF9Nipo25svgQzJVsyfQuxsFGe+d0CqsWDW66R4bt++rl9X
WGqs97mxHN/46gfdItBFdI6kfeJZfgndtQ1uiZGec6Kfu4LWXn1MoDkqz95DN8qR
nNSv+gALOmoD/4LY2y3KzVi0e3BBQVeQm168a/CIR2+y0CwOQlhiRl0OMLWy81En
cZON0N5HnGNzH583AO/PUahCo4HR4sAzOL6hIwm31xRNyrO8BtmAN/6HA8sEE10T
Dhb8ziDf814qKyFa8vqn3ZBhHVpHL9kA49R/Yq6i8UvS2f+WwMk0lmOtQgJR2uzQ
DGbV9zwvdfnITbhEPD1cGePFcMxGFMn9a9h2XInyRp9myFpaq5qbSGpVFVpy4l0f
9/h8lSMF3NZTgX66d1WT/wu2VxwvjNtMxFy9p/60yEisFlkKfE5uc2InlKN5gcbp
Bb/mBOpqp9tZvc1y3fNuxeP5mQgg6OduWC1mhr7HvZn2A8qFnWxuUqk69j+l/jzh
jMrsOxlYVY4Bx0VodvWCaUm6yznJ5nL28Aie0A4cX0SKxfXhh6xgilIpCkp3RwwH
+bSxIzmU91DjLq7DanLDurJZqvKR54SksfquI5OeDniGJlPFM/LtnXW5zrvOZlco
Z7pIrJNYsQchf19EiX8/qoLuLvCdhy2U4YcOtKTxZ0iut+N1tlYlni90oxpkFfY4
yCPm5Fgtt8lz6m0+WCvPNiIYdwq/SQw5s3lZsGCHGOX2HLWjoCTUjl0KbhpdHT7i
99rVXYvyvGU1e6Ki/aUep09h4LV74T8guz7zsxpcBap2WK3JTFshUQIGUNQO9GTu
Hsnxw1Ij3HrRme+a+SAi/q0Xkfh9kWw8huzsGy1FpGf6/kyp0GLL6VZ1uGR4ikIG
BaxKK66Ur4PaABP4Gg62JTLHiJhCm1PnXUDRkiXHGFG1igmyrX3qK+UYZLRSEHJX
lfCstQSfxzTQdY14XXOdGhIc3TCgTzXoeBlb9MgB7OQSi2kGwMYPTWGt5Foso74/
8mnH0oLPosUfzu3ZI/+F+slBdTi9TwwOUKQfGg0tUk382OtkNmnzQIytqDcQE1Z9
kCFVnRIAMskqxCZVNat6xPiS7rjT2aibNwl+W21eQPtePQ3699JV/b2Qmy7FVToa
6RTH3E9Rg2rF6bkqMakDayRfvsOifDUpSfWvTDwJIGsPCpmAVmGub7OwqxLaw8Nb
02Gc9+lLU7u4bCAC1Ip7s34an9fUv3bNS+XIjaumtyhEqRZHD4IEJSCBYHb2d5mb
SbQJgdDAtgFGur0iTFZDX4a507IWUaxrhRL+lvTfN2+f1rt62aiCQLP8BghxsRLk
CXl6GZLxJneoXTcAmUO3DSHTAxaofI5U9e+zId8pgB9Po+OsNQd5Cbf3ErSAwLkn
uRPX6FdJ/Ig6Vp4s9d320UVaEGNcjKd03mK9+Uor+u1KFdRJayxVFE+AoJMtVNKg
DN/svjFkM9LJL6Ryo47KpYPAVQnKyebl/RBn5PAmQmn8sFxrjt9KiJMOWc5rRhLJ
7TG04w0efP6XzxQSVTbl2L6lu1LtXLBh4SQ4Oyir9X64qyZrK8C8HSnasJFybjGK
dXpSMa4Nwve04TGxR1n7F2Pd5M7oeW5pjzZTVtDoTUpF3iQqVkgd8weM+GWAibLN
5SszT3RuBSLMwEVj1ye07C+TknTQrn45CKDJydgeB+veMDP02UEuYP/qFmKUGYi6
VoiJf79CTMKTOGmzhkA5ItmtYJuVo31fSSG1YYHBmroKvjyvZkzPTDt1OgRRRAbj
2ebBG6iEj5YHbFd62mgKaogds8GMty1VKMbpsmA1JxhquRth3ugCN4yedy+NtnPF
BT3D9noNI8FlG+HVF+GNU+Ec32KcHayGCdl4hJVs3cRHOIiR0LqAWcd3xlqR5CJZ
CRXVr47UpOjczjyQn3fLmX8CVXTPt3f4F3VAx3XxarZLqxVKs1/vYV6zcobi3cob
opWjIfxOlaAiwHXVr98dCQ+e7lZpOKPfH1cFlJlAAMQsofTm4B5ufqgcAVU/fUZD
RBJhgbP+XBT8GLMj3VW3WnL3Qm60JgTcBjX8O/nW+MDkXJ+WyEsudW7jsvdmCAnG
SD4T9PuoHfNQ98IsopZItd6X4dYS5Af3ZYse8z/JggISZIdqYskhkNSj7/j/7iCB
MAZYKZFsI2sR04L5y2E8Q047WoWQI+ZR51CU4htqG2018RD2uSs7T8nL4qp+TXGU
lWvKRBMjw3J/UK48eU95g5Tumw2V9rQ+RZK9IFaVVOHNRQyXaoBhKX8st+JuOuBf
1JhUlV+kRhcJLyVr6y4maK3rNSBQDiR/MT0m88nGFkHysOCnS3f+AZhs5WL7KFF1
Bd0D5ChKbcqwBgq/Lp7rcY9r7+gWK/qRghNuNvet2ZtbdFwPhNk/SUdnhTJ2YIB0
9HktMjqq7oe69vxm1fYrXDpX9YmnIWlxBWhdOQVuyldHXH2b1kf+naE45oHC7tmw
1K6FksOBtZOXr5nOY5U8oX8YvmjcajAKASwPbp79rDAbhsF3kvJowtD90ZAatdbP
byU6ERPZLvWJvqb90zhFe6RIgrREj16VXNgJcAaQ/s+ZVzHpFEOoqG2pKFdbL/vy
gcPvcG+ZTuPgHJt6hBVApUcsllT/DfCtZbcjepcjPyKMyXPcgVXbOpKROmDG20ZZ
t3GY2lNTcZt01siRiGoSncxNAAmNcJB2bRxYqMSfvILty/CTFcchwUEY2uzxP1LW
yJ/D3d9wMdud5qs1ZulpnDXGkE3ewP8JUSW/S0TPsz+AfhPuFYfcQacOeolumglr
TDYNFcZKg6BbJxXCspMQD75DRCSdUHaJ/WJ5kGdpjip6a6/jLvxu23qlzR/NSqSa
ydHX4o/YssaDt9G/uienjHDuUY0g1pM9poR+1jaMsU2xYxiu2bI83zGR8eeBP3Oi
FlBdwhl/MBxCxJeMrsKwdBz4At3Sg7kM2lyvooea1sXxE8yFu5X+ucF+PqsBqbMR
ENyPx4EamWNk4Dud4rEo44r0ifAOTkzLPP6PzLS4lvJRHLR/hkk3MYT+9hJ0DTHH
kbbo0CWzdHXyA+MN0aSIyT5dRlXKF6jmyWymOYEe3JiqU5YURWov87upwoGbOxDI
oQic9y1mer1e+iiq0jRAwmssV5z0JbfmJKqv1xeBhFBz+tb0KWz6VtBpDZJitE2i
w3/QzPNzf9bq+Q3vLRJXxNB743/0G9KIGGzW4EYhSZ4QOiRliFEn08rEe2/+sVgR
/3mwmAuQ/oql6AMgy8PLywdnCyzSaNK4wd9kZ657Faf0QUQQcZMz+7DHdNsyQPtF
wGYu+WHB9urYE1VbM+w+Bi1gP5SRCh1HY/cy2Js2U2XQzTnBxPD7l+kg/j1Q09Jj
w9lYx2J8NK9NK8Qw4VRiFnApAG3UDzHEv08j+QaPycFPWfOpL6CxnVzKDDnMfqWP
qgP8ljGG2xSsLzFzzvI3qiVPcew7F4vq84u5SU7aRlIkHJDpLCjMHVVx4YuxebhJ
LQISeHusYz3bBEzGnenfkd8yD3zZILmZBgU2KiEY3RFLmjwDd+B1FwvjJwVsBMax
J9oh9QBI3IB3POvR2bDb1clks7BIKkkNhQ9FZDIX3YAkWaUgzoJBSigfOUL+Akee
EhUadaLrNC8TaloapLk0kcYlJTP6Vhr2CJXu9o9ima1LU927DeRwV/kxqheqxWMa
B+3dY2L3SdaXMLaqExRYmQz/+8VX4dqeqNxYSuzijRgLfEe/gE016sum0+HSZp0f
8FbDqqxwCCBZvcaA76E1/B/3gI5hxxxSx6WVizyMGMxs+lJQawJCltaPke4nhu9y
xTU+r5KnEqwOfkOslYdNP5W9dT83MHEL69MzZCuh+iwGFtYkxYoWeLc/pSJpZriO
AX/uTxuudQekrWwg3Vmmagwf2WxpFED6rE2tGFvrNHkzBPEM46DxrExR8QhT8SnC
hNZ/KSUIwbJJF2QBDspg3e/KQqMUM9ZXfs/JH2QB3VydUL4RIuJQh2CHYlOeh2/6
o/pgh9ZKmJhdCGuz1qO8QmDVNajWtXT91ticW5SavPRVlU6Z1/+AJaH04goErKBB
OHwjpIMmLB7kI4osI5t7EbhVFvUyrnK4b43TSOvruoo2GPuVGo7tORa4CqiMiBoJ
dlZzRhCFrJsxHljs3cayHAMLwg6p4hYQuatOQTujtzR60vEd/P7oG+Ef2koIiiRC
DQnv2LoBPx0/1cEd3y2OQqL7SFu1qdHY6OQApZI8sG8icL2DXkKAYR0JDeKVgv85
O/PGuoI5sBiqfFyfWJV90dXGV50XrPtJdmxysesoh1zOO6LGWh/QIzCov8OPEv9d
7s4JrB3nkSOoO/8ZS6QT1aM7LY6Wn/6i0ry2BTlNLtqhaBZ7NL/qUTwP/VBOmuzA
L3S4+bGMIdvaJVsYzZqsCc6h+q4Cqo8yGrigmR0w8gL23xLWDBOPWJicLuSygr5o
6p4jpNrNuX9sZFArXA7QLLW2HBDeqyR5GV7k5IepiboMIXJBq04Uu4eG0uKtl9eS
qgUfU7L2fRAURD564dbJBe2mjpy/pYbz5llFLPKIUXyVqbN+likAcXahymFHXKuC
9MucILlyssT5yZLLXaUiDDg5RApsqZAfZafZFtCztuyY0iXxxxMyvW3U8eaSlS4e
djgFSlZsJx7832Mljq6nuMGRrR9VuD1N5TeKHhPoetqlbT8rTjZKjyGDJ+7P8jno
R8n3DltG+4AAyxYh7bvRhkTmu67V6hBjtwXrn69g20JcES/jELfkmGu6se8/mLpH
mW1NcK7+2ErNVN7yysB2bamtaEk7Q4sUyJdSdgMVpjN7ZcHLzZyQc1jSWu82Uo1C
KtqmBmjiDJS8egtuuXoUOeHtto+S6OYfX9HZ2N/WjHxpMu4xA0W+EXMIjuJJvz8G
MSXbjfrGwuPfIBi+NCK+UfyM1XRNcXpWC4cWqiZpF9mQ37CTKWbEkLOhOMwY0V49
Mz10derc9ruYIepOwYI+Qf2hwlwIyY7Z9tD3w8ojoVA6/Jr53HZQD72OYozwqea0
pMI4vnuSt+whLb8lIf4k8lG7XWkicjjez/Efc5oNh6TW0pRXSLTqYxd/Klmv+OCJ
oRCwlbhj4xrBgSO1CuOpd1sRhs3nEH6FtiixGqj+GPo/o16dLHvz049aY+zW9jL2
n1zbuOHGvwVcFX79QoHuA/bgUsBmNloAnCgSunkhs2boMTE9NFpTdC4U2cr9VHPz
LaDtsnHmcKfdIM3jKruVCIphfV+SaNivkulF3RpX4/6amvf1KGqV5R7o1v5Z+C2T
0+1HGRQbuM9GfHWpFGz6/oeBQV3DEIoL+vh0ek6feeWsOYZhIQjIOlxcUOHh1aye
0F2gMspwJYhxK52upLrbGMaKj5N8uxBBVrB/3VW0jT36RQLryDXgfxOVc6mUU9C3
x6lQ7mylnZGYq3+n7Un8IocM6meFEzxiDNg6eVBPnjXGyGvpCJuKVZ+KmGRVXlZ5
w5pc+SMZ5xDH3evvX4JvkUnXE5cQnaQhz/SF/dDWY8iLYMBXKRvZVoi7QkmeyQRj
sf9vBIKw1YuUobZ/blJ4VGpKaltAM/Fn+dc2e43ijxnxUQkyeTiZDMt2QMZ+FDzu
fTAAMxpGWjih7hK5wftlOD8zjbfbqxNQgqT5fMEZlfx+rlADENTSsHEKeILvRaaT
+ef/RG8MX7D9l2tOCUQ7leH5vj2Ok0gQpHMEpXOasfesRHZgZFOeiuqw04dRM3Ul
WpLWeoq13m7KfoKcT6gcr+ly9Cbnj4L/3+mPm+p4hXkOQ+RwvteC92kuc9aS8p6Z
YVQ3h0VGJeoeKqo5vKFr3Xv9BAdU4GBkCidRX48OS8tjHEExO3NFJIuPdwQmH0dE
taTrVxa+qG7X7/Dg+mRkiucE9CwHOPrXjFwle7vqNo3INqCEqkvF3pQZideOoxy9
1RaZIvvKOWw2vwoJ1TYsC020SAUhwhJA/pSOGlBOJ3jAKuJhmVQXv/E1GXRloQLq
lqjZ4pgX84lqo+Fz5yVyZ/SCoGc+QIMz1DqK1DyafySSXNMlplycKvsQQVuHK8VP
UjyL4EJ5jYHKdp9Mk4l2+MmdUShZPi1vtZVrJdbvY9fLAuLXc597irswC2PBHVMm
VgicC5nXUKJA3zIKC8jIfh7SAX3n6ikoW0a8HER4iTH12zLQ+uopcw66dBYaG/bD
QjoczANXam16zhkIVScK6JBxTI/JJQOmFlBbm967jy1rrRiUYPA8r46f0GA5pq1X
wrQ3Lx6hrBuZW0dcr28mmsQANlNMI4sfupb3ZvSFku1kBHIW4OmQsoetYvhM9tmt
o7GcChWacFbDPYfHG0UzPtuirnV5+7/2Dd8nIgSYaE8Io/u5Lma6LbkDmtHG4IIX
iadX0x46NJb/Mg5Pzc7O6NdGsEJIw7hpJNqnMPGQvoi1zBpQMTqEFg+TRwW8rDB/
UsQIFwEp8UGqu0X6MGqi2UgTxU0/Rz1vLAKeLG0BzUOusJvreh71iw9n7RYaHvd6
9NhRTQqPpglZRuXtPz0EA2epujHnVSTH+dtoRgm+lckOwe6x1aR6Nmhualp6SS7+
7ocKgoUblZPvrrxAurJrtuhSeUkd4cpoP2gjMYiUfvNAzIyUHns1XItO8XKFeMV4
hLY/uWjnJw/x7LAC6ceCul/U8u8kJfYbDS/QdFN5wJ3/ruNVmEJwHbP++7nwjwyF
KUcdJ1JGMB0a9iT9M1Tcc3fi/adBT7eZAuuPGKHYQPMvYU3UINkurw3tKAsI1ORR
/38pfJYZUEH7qO46nSj67gRRLC/zZp4iLR/YWEMxtioE6Ix9+k7aXS19LGa8I0Cc
inxSyOfDkzbmaLzqtrfSjY8AOWE/c3eHDHLGnLM7bGT4phkN2oZC0Mg3Lsfnb/P6
TFX2uDjMSxuXxqtfjhsO98BntOsyoNGOJjkZCZEFiMP3ISsj7eh524ZqFC71616/
/XuRNtlejyUdOFu/li2xfk0Osc9WKOAkyzIVEcrDwbDA9x1PlPeC/ZYTfXxahGMB
Q0kufaz1og7O7524ahAHNV6hth99OKsoKS7qwyNGPoTf/MNel4kc/TksHncS7M0R
AmvifJbUPDAxxCoVJlHlUk9Y8FtZetKUkimXk8zO27X2m+a064k+lmCfFq4o4ufy
xPq9K7z8TdZ5PtTzByX7pal4Z3aTKBA2l40uzGD2J9hMvlnS8Ac7eXiTRAOpWH8n
MBp1x/GAvjtSWNm/g4lxO03Z14l03Iyo0rGs7z0JAiXDdiU3ybyNGrZ8oRpdeChx
YcSgp4ytXnlDl7nEW9abmpfwRrh/wFIKITuWGgcfINJAMyrQQ9nB563Nou76XBpG
9IrofiiqdTDaOmSP45J8tq1J2jPgZgiC+c9rWg6Uoej4kMharCttTh+oe6UyKv99
JX7JTlYttU6KglwWcEpPWIcIohSiN745Rw5xr3V6clNYiUiwLQAiwG4jrdnXqqxg
nGXQmC6xIHfrQZW93xN0JFtK5GhGzib90naDdOedD4E+52QW5jNBCah0gvoXGvdv
5YjROxUpnUXAAIfqH7fOyPrZb4PX8NY2ZXzTGgoKi9IgQypCGf98pW8iPP6T9Tvs
jg+ZQWWQp/oMWMJj5L6gtQv787+Ok4U/YtYfIQTDv2s9su9uF6/DfTyMUbGEU5fP
EH2Efbpu6cBQGPFR9kgObtd76HuJowCuFPDIwvQpiWkLjuqDPG7Kzh4Ip36t45j6
vKN73H1ooH3rcMM1MwxtNOtKmqPrYs98yRoc2u8ptzA5B7l5Ia/VKd+wzurKzUP3
tLIt9JHAblcNbT8FvtAd4/BC/nwthKfAeibumBbV6yoGpWLcQWcdZ5DCsplbmQdN
GTa8zdmEUpqKNczd5SknOklHDQAeAC+ZSqq+Xe69Xn4cFm1HmrSeBhitXmDW9nDo
Oem4PYcPS3X5gDCGZS1knuccPAmcgggzw+LlL0eW3whTd2k5lU6vsLBX5ZvX163l
xtgL2pUgVjzMkg9XuFZ31tJsyb5BAx5x/PpZXBjwSPZJm5H6WgtmREo0a5jQFhIl
ZBAUpSCRR8YazWN+6esttkGMQj/5ZlDFwG0gKQgCLHwCCbH0qvoWN4I6d7RYyb5z
GrFgQxcc6NBKNOx207CzPKssDJNuMN/93uprYOP617SLJLuVdzqttmgViPuMps0B
qaeRkgFkU4fHdoLu+X6yAgyZ5B8sahGKAInlIl3v2kwzKbzBNi275EjHYyJrFYcJ
1hBgJcI2joDRimr/T+bip1+M/UA/YIZB6IR/B6lZtfzaySzS5aV7guVZGmdlMzv2
ikCjAqN9PE7eojr2lGQmRUBgHEsCj3cYu6dUPBNXQCGJxmgeGGhTKblxQYmdGznm
ZDFRiSWe1QhFI9RnIB+3EK18kVYZr2jj1efAg/c4C+LjYvQ9MFVX9ucfYyRwLF43
QuQpyZdf1hGQYjtaXUjRfBo+O/XUFY1pOytB3cnt6vWL39L3BJgdYbCjpEf5e7IS
lzQlrq9/ZsEskuTIcU2wFJu9l+GQGWvAATqzfTb6lTNWsArDKcQ8yiiOreI9zoDX
kVoKasfVh8rye3GBrwPTy0Q1crMrYtuMZTtQJGAV7wq6KrCEtivx8p/17dh/vEqc
Usv9eParhBSOgl2O/LVUkmbO4xg4LI91VVPgjFBxn4PR85RWJzd0wDHkroh2vKuc
1FdL3TEtxEXWsZJajI0M/yREcZwJ+qxhpTiw3NgBvR5kFHXbCe/rVcuFGDSTKFZH
b60pnkz0lz5x2iGwIeT7ZBOdIB18T6EP2zaMveZbN5Zo/57Z2mhc27nB7NGNt1ae
eVTyo3UghJzkbPxGzu8lGGQawKqOHf4AbJr1SD78a2+d4J1UTDl4TkNqSxNmxCnm
bbQei1G3N98xFTebgDqNCRRVIH1ttfOToXpR66f6Lx5wVCmdyjPisq7F8KdbNVnx
T5hs/WQUCpWa9SCR8zttUqSgTr3bFsKozsv4Ppjh+SzL7hIJ+9aAepPrr9VrkY81
3PsRv6lWzqVqFsiREwyYp7ZQg8FhSRiZsB0e5Rkf5rklinaxqZ6yseaAiV6EwsN0
gHnFv1DeNVvykNkBuPs8Rnn0o4gNb0jHM27ek0G5b2g+NOFRm69q/mXqVqidLjWV
N83m5zRDNlPRa2CYdLEHedCCz9pJl01DKcCmBIkfz6BV5DXQrot2faVT8AN6DAKN
FtM2EK7lxfXEQwmrHth/ujOPkCaQwd96cI4eZnrneN7S3g2j0pwwBS480PxtZj8U
pi/4LV0S0d8lJwdL/zMT3WOx98wwVpmMi5rpk6HnO0us6Dyp0yP1PqFaMqIs1X6G
8Jb/wdcqQdceiv5Wqfu+cX3MAcxc0mc2HseVdnzcOYTPlJ8ezBKe0GnWLMllY7AK
rw5XvlKL0OYYvtVhf6DMQHmtC5zZ4PDfznzvSzzyqlh8OyRRsdbebEsi8n6Irk4j
pKzwbefvU1L/anJv4jQDuntV6kjM19WRz0Q2aUbWIfm7//WmdxZ8QNnHka1fS0F1
6nkF2+80pX0XnwCF2FTtnD02SlYTBTsNzmT2s7kYB/WLELv5xDfLhmvjSuiHSvVQ
wahqzcuJlQUw+aoLArYA89XBOriRPwNSW889BvXZAszOrg2G5OmTQ3nvfDsD7y84
9w14BYjN3DGM48y4ZM/GYweSaoQrhieldqwfjw9ikCfADdWw9L2aSYBdKLAu+hN5
ZLKScscd+xro7prG//YWrmxKpGzKmLmU4Iy9qyZb1NoG4YY2PYq9+PyJVRGSzEi2
a8ba+LsM9wkXHuhY+B2/vkovEcrq1dTM3NE5S6CPkolbrv3W1TQaRfhlRcGovQXS
wd7gP19SVPt3++pqSHeZbAMMg/5xcUl15WekuVQZ68cMvQa+RVoqzzo+ezD202/1
QkXuVgfqqopoKywALslTnJ4ekUitaXnbLgHlJ/al2uTkHVBtOYSrk5enoiRFaAfB
7MJpmP+vrEEaLbuw367US5D8FpNY4OsXXrrMJtkUGc26DD1tL6yl4tOlAa9wOxxJ
+zeIT9RlZd0TkZ/oysZZgRdm+oTSiso7OxfSHSS9V/Lqx84Vc3ZtF1WVCk8D1ckA
UFih43A9Ks7vJWfQzItAFA7CbOQsSPG56aqtL5owwqax4MtnGmGOs85rPXrmGfKT
QGC2+KCN0dHv1mx1Ir8Qza3hUmnTyu9tBC5qbkEaZP/h6iexs8JrQbO/33kHT06o
pLYUN1fonTEjkVWqREAgYH/b/ktbOgJh7Wl52z1dNgp9+16dfUaeZaZx7aD6radQ
VP9jSZ+xfxs021MRujlwxx8wn0rp2QpCYkcxHtQsq5j6t6/pfht0PH48CEiIrugh
kD/IUfT2PTcuqvzRmAHICa19wOa2FM/oSywGWuQtkHQw2avns/+Bqfvqhe7JzK4E
3Y7XVvb+XAtVprcHFBxQhkELc2TXQQSS02zZNilwBVAJTqPU28sbyYnJhlKrcv+M
mSb3J5Zbi4XZubJ9seb+D/d5/Wo3bveHStsTa+m1USix1ZEOh/SjrYyKohcAoJN1
BmMzHPBQUEaRtAYITRIg+b1T/EszihANfWKhkrIWQJQAx89GUkzZ5iXMJGN+8zRv
HTECNkbsZH1YP44asKFiIhbQoHFnW2hvFZKeX5zrTpM9ApHGGFLTnz5ZUoxiHfgh
31YrwJCirIt4CKZHk+c8PDx2KQ4Q38WxDpu3f9PZTElUKDRz5skoVilj6ac1cj5I
GLb77tLFu4A9klsB0kyOjisxZamSaZYXZgLdvavKx+VxVTqvvskpuftZg+jRcbs0
1vNGt+/NCRzyJdVDRcXcJdfuliuJ8M5Waler5IM8jjiRNT7Bx8RLacx43S/pCON6
l0JaC7LK3n9noZPHC2nWvhdVWp0Nm4YJ1Mu4aq/pdQp17E/D3EOopR0fV+DcGnuk
5WeepcyjjADqbOY+/zBcfbWolc0m+TCjfzp2IarhG9enQP9RevXg275Eg6NfjQ8y
Wp3OT2vRmyOYcLeGQP5N6bOyP6iaWWwrz74cfwOY7x/JY4wX5zE22lyClgHRNjBU
YO8MzXJCrIigNvCWzk4nVqIDPz6kTx7wRCmBfRbREeRQ6ck7DaBPx6iq6HfU0pme
iSQ+hMnFvU3hSaUQN9+b8z4jc6TFq9LOM7lqRYSs+yDcgVSuEGA1MB0W40eD6zh4
xanWxseTrMIh3N3xhC1LEV1tDW6n2uIWgsshS7eUWs+RAcRjH6Bze575To5T3fuG
Rok6UctH3MC3tyURdz2n0PHS/ZfTg58CzrZ7GP414sgYhgEfAx2n/pMcWFL9HFHu
fVPPJ2z30USRrFa/OgyLxo9OhUc0wVQgyU/uX3i+HIuOu4vxrHJ0iSOcJX6BAcw0
kKhgZ5n/tsTPgS+pn502YXWYEhUDe3iLB8ljUrYTU0IHjNsm3EBM4MVvtd/4riDN
ncWSAEaUSWLcE5eE4vJqKqaupNOWyRvUt95TlbuV7yh7yL+6dK8HQ8Kyu1OqhqdE
SwDlg2L2YZSsCQuNHZEJaY+weavq45KycRLeZelgtTzv2gHXLZ2Zjb8+OmGR5+zG
g+ciFTFRNvtiujvGEO8W5fTItHXpn+rBE/uGo4RpNsXFJFrLZsCOmBCtfZW7POUA
H9hlAUX7L319UwENUvHm17SyMv0IPYg0t3b/LIcOe9JxqnvM+uBZKO/JWNfiApNX
Sgp7ZGlovHDRyYJlMaLOhWD7PgJGnw1eE9lNwXQadqfKMCVvMWpVCDng2JapXVNA
/+3AsHzDwyW6WjVwAn2WEmzyzFIrk8ZcR0Kxr7ab8iaqlNNcyJAS0yQ0l08XH/xA
wmuhrgYEaKHGbEqt9Q4AqEOCYdSLqsYxXHWDwh0J7Nvc/um0YdzNQcb/UWVeJWjm
JvY74Bm3Ao/L7GFx3d1b4wnRx8/VGYvIz3Nm8YBVnS57PrFJJR/Wj37tE4HlK3Uc
lldRQSoywICuqoOgWA4hXpS0AbzGBRfSqxdSHSDmRcv0FeQGfGahc38lJHaWhCAB
5I7l3YWZdSq5kANja82XhIyGWqbeOZ7Cesg5weLUDchaIrHV1Df3fkhwFLvLgdgO
ZiY1+jKm2iJKwJXuDPhkdERpqaD3zRrV/1RM1MfOFrM349g3+tZ1iH2+LI8qBw9y
5uP4xwWnDlDwq1C7R1QlgK1WU7rbgveA8dH+1iK5unJaXHMCvRB7fjiHIYNeQnDV
EczzXzsmXWXN0BgCLHWuAHZ2q5vKmhPhSkYlw9Yb5dJ9Km7mL3/fzeSfpdOoM+Mh
qhOHMKpQYyb8sTixpTdrOdL0NXwnWmVhF1uPiXbDJ79G8w8gSC7ZLKBtLYJhYBxA
PO3T3YmYZTngFqXaHf9V2boD7nxfBQEmoY/gVBOQCdACT3FA8rbpkmqxCoFN05yN
+79bctYvgsEnd799tsxTqmsFGgnmNM1DcPtI33tZ6ZSRf4NUj6MExYIVBmHtNyZ5
MelGiEbE+E9LIEDB5uvfJZjd8CfWZ3xOvh+AkNoI5RWOtB+Co8EYxCyDvErxqh12
QiXnD9m7ZUg2Adxrfxc7y1RWl6OyZce+m16k/vmtpksfINNM4YIRnfHsIoKAIOox
q0vBWzzDgjc5uhk+EjrpzwKfC+GsYvmF0TDjlD7SuhcGgBvSn633gTZF3sZuoLO5
4O390/1X9ZQGnt8MDIp6u4YSP1GrSjO7tP7Vb4ZGbEm2UQRTnumW06GKePbe6Gq3
8iDEVlyQR0dcYyFHtGYg6Dujkk1UvfgG77xDz9KX9fX1HnEDkHFdtBOQKfdBKa4f
BNG0OveXcjA2h/gZlObH7WS8h9UXqV0I0uFStUjf1B/weJLxxiSVWig4RgL3s/oX
HaGppfTSlCf/LuDbTz7hVKA4JWwd0+fu6w9P6N/7rwyrANz068aZPjbaFK1jy+pv
bVxuvh9/j8+qmswzaA5miWcu8wDLaBHczcUTuFU3S/JlaCzSmiXiLn9X9SDIgFF3
I55UYWFL17UzApBOwVlxJojOGmGAfvsj6UspwVd+DbfCqq59TLtwYvz5R00jpedh
lexEjLfW23Uq7X+W7MyX1c8zCZz7RvvHCELiWJjjWX8TtwRBUAq/IlYncONEfpl7
K4jp41XtcnFzeuyesSY11dop4/cys89Xt6z4K4X3VDe7HjhTwHFFujgqTUvRL3UE
XsEOwAI5/tQgfmAwsfUnkAoWAUeifbsjW9ILW8i+da6arBp5BTMQsMe7v2Y993KU
/oUqfPBcQw3Nxr2v+NsTTzFBN1qQYUIkNQ94IqEtqrNNQadmaJtwdE1EkFpMk3eO
Z2QveceHpT8jHm10PpZ1br+9mANqZOfYIbIh486eKBQsmmPDrQEAOlYlrZOZMYZ9
kmfyBlfxy3xeraXrTOzL7xZlQkry+rrEu55hGEbYIMay1TfodeXkjX0E/FZN9e4K
Y0BlEP235S69+W6MibIIc1fqggXhXIyBjBIbtSd5LfTCoX8yhEsPBGJHGGgNZB7p
yn3tMTpH5ngC1MRHmGgrcGdpAKFr14hdfq/E0auYp9GdZdQdl2dqyIz54IC9PCP0
w4ueGZGLabmd+LgO6UXnbKQQI9g3K2R5z4rSuPHWVEPjs9riQV/Soqm8Z1fElgIy
GudhTb5RwOM3zfHSPLLQ0vUmyoBDhs4DOiBQ952HtFB030m2/yYVwIXmBKFR/lEk
vwknYGRzQZ5CcZtcAxwfrhCyBYMUhv0r+Aiqt6dznt1fxroSN9LNYIpLpRHIt9x+
gmA8imHW/VAP4Qww7QId5p1DilUbFdicO8Lo3ASc08nEIN/Q+C9RE/VYGqU7Uf4U
BQBBJ5jm3MVy3QeVkSIxbhZ74qk/SUad+gO9rcDk7MQx9P+nFINekCD52s3NT5J8
D+MiBKyhNk43ZMWigT8ajbdlVYCaXmzVlDOJQ/aSvyHz2ffZFm3Dfnzsimb/z8wy
IPWzTPhrqdHP5bYldWpVZelVBePMOI2/4exftR7k6kfnfbIlks7nk0l2nDd7N47g
cv9BM+nqeUPAInNxvptzfkdlQCeMMygI+dssIFF3M+52EiUOW0VSJ1AJbgNdy2ZG
6ljobdcZE8ncFaPz3f6rSww0O0w+OPDDElPuZjO9hQkvGYBySpZl4mI6sxQ8sn/q
70hypzrP591djIv8AC2KTfyfH5Sv6bra70nNa6GxH/eY4wKGWB0LNBgk1WuGKmvZ
QipDdyKGqcUAhNcukEUim57p0yvMYOQEyBL0Exa9TsCSksbFnE2vSyPbE+baaSoE
JM8cyL3a9lIBzWHEKBgjkc2x1eKGIyIDcuW2VG3RhbFUCjBgz9thPehkVpiyV3g3
z9a6/b9iWUOwg7wVwWGqMfG437hk65o9pog0N8VXEjPEmkl2kfSza5AhTAUA7jgT
jY7QNL6bpttHunuoTQzn0RVdjd5GCWaoo56AJ4kgwyZkBUiH72b3Aw/U2Y+J3+Ns
xhUrZmCtsT3sQE/JWzxaL6ciftr/hd5+XYzerNbgRN4WIdaX/EAdwRNTtVDWQ0EM
E86QwJUgRFEdXdQ4t3sDOIe2cdJXc8hGsy4wBlDDu6iM2dSSkpQZH+g03qsI0td4
nooEOLuL+AGICq8dy9bqHULCK89CIYkdw4OIGCnnBJwpVzFUeDKKFNYyeM36u55c
M82IqMlWNhfgBO3RBNTAPA7uVeNvWHC2AnKzuEhlQmPFFtE1zodeV89J8g1JOZNz
Dl4NuXGl9tv0nEwj3ACtYkYuaE93BCDpanoFgkI2q0cnuKz1sUXNeySSO29hE4Mo
nBDSwXsVcRDyDIgE/dnFuznaCq7h5g8o2JYY0NI4lHDwe+EQhyczuCyeO/NuMwST
Z0XK2ju/X/pjVxcszIxoq7bzmaH4MA0ihYTCp1PO6yZnmwlfc9NFh88suMtBuOXP
F39XYEZs2dzfM09Agzd9ixY8IopYDIb2pNFZ+GvTZ2alkyq3fDExbyujo2fXdTdK
KYjGb5S8mXZsNCX/1uh8T3LG1g3WmuhZFmwA/yNURGE5PKJttG7i3XHi4Vxwhp1x
xnANvCipMCG7QpAr6mxCLLKeup1UIzCardFDcZXnTUymCKmUfgWZ3wNErwFra3AX
lKzsBfil13cFInBMu6DSYbTX+3TsaDOJTCOqSU6KUh2QIld+BNDcmY6Z2lPGyA4K
/LDlYSmcWNmbEJ0bFsN9QUu8g+5k5oUlmkiKNhbnqOWhLqISjTAhfMfYRvdaPvSE
2k5Wloe/RGCz5O5BVgPLEE6T/zPMlv70bYMGShBNYpjr/NcS9niqq6XcE31hxLcY
1kLgqQ48/MKMTz8ywDz5o+rmvQYNhYeNlprYyYEdzC6m9MbR7RFB5FDfpL3OxEh4
Co+YRI4gZMmo3MqCYfd8psEdI4aV6uvBAjaqoYvrIduXLjRQ5pLOTpA8iZ4wB/FI
QKhCxQlc3xnSkxUu1uOBLeHrM/XS/3nNghV8NHUK8JjTg5sdrHGlsjmn4JgFpZXP
DOB0zdGR1AlkqKdJGi8VbvnhT+b2rSLN6FZF/SnOMUXggwAItc+q+SwG7viim3GR
+80e8f0gDdwPxPL0Eb3uhuhW8gxv5kc4N7QBihQK7dcy27zUwCVQRjFvER3Rz470
6M/dELNEW2J8omMXwegOy9IAgQIglMG0B0wqtU7Bl3zW4EFysUS6eAQ7f5SzXiWd
GJI30gWR01hexgd5MaOZxWiVGjfVEQnUpytlSQ/Uddt3Udi0f/u4WUuso+nXjBha
cYvMfvzHUtQUOh1soksN2MkwizB9XxXA0Nvo4IsmbwTlJnFceIPLyW2MDVeT9/2A
xlbweFkbF6jmrg9EuzhWX8trM5aGFwnvFVNK3mvLFjCrte688ROA859x70hREPqm
QJ31+mkrXFNprs0IoNV7Xjm5am6gj/Li7hERDIZ1Q+0dBtgSb0jOHULYGEi5RRbP
9k2ii43Ug0TPsF8Z9XNpnwo+YQqvLv3JiWdJ9tEJ1XoYRr+qHd6jY8adsdkh+FW6
z/w5GS8Xvfs/4I8EkXStlaUMrcRlVuBy59DIZqu9e2dm9MpKKphA/rx5Ymfd7BMT
cRACW4ni53FBTK1eYHdInHJ1zamPhiY/HgtOUpMmoJ0dJUeg6SO3OsBsKnsRC7kv
3l0vYNrzNb1oXsh20//swtNHKfzpuz6zd7f77vjZRsY98p4JNNO+e3U/JkKEljwP
jbZv34LVf7BxKnH7X2hKR2Q+sWnmnrpzODQYntzVcPJMNasOT3kGpXy/I22EWR/g
61/K+V/LLK7lzBe1yHQsvxjJrS0fg3YWaumnfxGU21EipLZmSiERTAsJyqTTBwXh
vEt9K4z0CrwhJ8UtYGMGmMcG5AlBFhyXSifPpO45kc2zXvbpsn2qXZVi/hE6eUJ+
2JGOzk0BU4RkTyzsCnbU+82QpCm9DgaN9CFJFw6vIvEJjDlGyAQcvw3I4njCfNY5
5Q80jPGFkcHQ2KfvRGL5HOy/5HqdeNVJykzk/IPUwUIRnCK4Qztp356ftYOj9FnI
zggiHI6m9pUJkpNxg9GYZ3y4FLiuyld03bzPf4CRg2gjIHgmGsFMGlD65yp/qftn
gvr3CpCHLrDzKN0hi5QPr2y1TYKkV0YBKb1Gr1zrmMe7oQQnZBLS9heZiKGirzkA
KZmGoNwmjGCDF92QEHR/vc/yxPbcA1Tl699Dn0z4WSYzD9tQYAMt5kP+nF64tt0J
z1vFcqRpo9spXoNbyP2XS80GsTN5M2O84AzXvzwPB7NK1Jceul+A9ZihG3xPyVSw
yT7++vMGSC/ziFqVgFwFEyUNkSIM4wXBVqGzecvtnDF4xkioxCU3knk/xqORxcb/
95pIrjYRuH+iei5GilxhtYB9wNahvLP9+MTMKzzuzhBgCycl95n3w71KJ1g0B+tJ
7LESrKcjKEryQ870D+DB/k8Tk4WaJ0IbDiPFvtdXa4jTvhAODzL/SDRpqm/RyJps
/vEC2ZEXqCNupeWJDj1cV+sYIaCVmP6raV7kad3KtjkyCyjjeAtN79ZYzWuYGaYR
kUO7U6Emay/PyYQ6jxOkdoE1hCxWI1bBNGjK69fK/Bu5fdkkeAGFfgcaMSAYRx4X
B0AjyMtYYxQi5lVpvBJXUDtsdnkZbr3ySGxvwqt1Mn82HzXWp5FVyijH8DxWjj2S
gPsxboI63TQwXEEOJF6pFZkIvK6GEc9Ti8Ork5uf5/DvjKJvW0RazGWyKc3/FDAm
9GNvGAVxUrd5TcnnBDCO7+JFTXOKCFYiQI9bWCBGeoqLglS2HvL43n9CxNlrUEqa
PybCDj7ilBL2Xkacdz62PL+mm8THPIYUomMndLnMlyOT2wniJAOM5S6Ge4xtdKat
k9/KswJTdq+d2NbiFp2ylOri4rFFeQVYME8c5/ME8fwVrFEDK570nnAjBqhtzrol
V9Jq2coe3LSdUDHZJO+lrR+YAP7dBKUlBlA4reVywiaGBD20HDVdqaw4DKYvWSvC
pjQzSCcRLkRlTHiXiSDb6OKa1ltXyfbAs6eSWFM4U65/xCMFC3MAYL6arMuWsavM
HbRLvce0lI8qYj9rCxJLN2k8m6Xlsh7BBYa8dHfBnWJziWXG034U42NTCkaXbO2F
q1/sbrGX+9eJtElNrAxJeRVZGkD5KU64ykdM8Cb9bBK+oc5sOV10242g5aoVlXw5
kXcc3Kq1mqZjBOu62bd/3yrV0XJkB1hFIdAfP1fTO+Oj1MhORvhSiVuaXB4ZkR2Y
Og6C5FExiZVAyDEp5e1a56ocofGg5FB4jhKqB+QYuo45KCZwlrXzpbDpKOWPvTBl
ry4k0Odii19BQkf0voWMUbrt1XhJek5pwB/5ei3kxL4KgSNT99Y2UaqRd8TR7Nwd
b3C6kU3P0xr5JvwdHRs1kTfw7iYxXejcdGZuVcGVk01zsiviKgwVOBHv/nSkKi8C
UXIOHTDa8swZ1r8r2fcnWhT+Uppz5illyHUG10cSuLDgE/KTOrBVcVleGL53RfDY
6QN5SxypACAtUqNtPb+MIWIoNgTzROkXU8JDxajwSQFMf4l4ifLnQG/ByjiIvht3
dY4ZIDaZw/1g3eFNbILF3DbgO3aaDycaKTSEqiWb6/feTa0rnXBHAmx7aBTdlqqn
itu1pprCg7HZtsjjBq4E18/ofBK0+jFYp1AoSsLBZx5I9aiORSkuVNWQpINPeBkW
KNToGt50ZcmdtUTlaygakmALlJefflli88v8+SIMTFgWOuX6vM7KVdIhA70x8C0R
5/HnONaiHuXMMPrutrnZt5M6D8zOmC5xrAruvXpgNyHXD/qtYRQoQK6QDyvkksVD
yOFJYIbMH7i59FEiymYj4kkbgBsO6oQqf/kwf69eJVpKzxXcscDzjE0YmgU/l1dJ
0tTZKRKBUyBDz4ys+DO94ofyRyQyKnAyd6Oii/jRXjNwWcIh0ZgC1PWOxwfQQkG9
mR3zVj7N3vfallqmgemf3o+1WLPaITlXoZ8YpfKs1GfMYDxtYxrPpkPd1J4VMD0a
LCIUg7iFbEELi5eMVtYe6zXISQB4tRbjyTP75z4IOGT6C+ehmf31UbRDYSCn+se4
cNM0x+9eCMIuXdgcuNO4Tp9eY8ESdeJ6H8+C6XS4lNeNUhFaoNTm8I2ueZRkqrg1
zS6sd3MYccVQnDPzKHDUheCNPxQ9StHoM8AweTZPozUFPZD4rCVvgyTn3DgvIhMY
+x93mC9v9ITDtG3q7d/pC133vQHP/EvySNsd4F93JBxvuVw2N0pWc0aUE054Pwbi
7StGCru3zf1ra4bFBYePJVXjA4Mcu/BHeNq9hmGJpUaT+ojQLnA1p/gMf+Db2pbm
IF1rmOE9eRDPDThiL6ClbXPmlYdvVm/BbJSd6d+DJJr3luT5YSgDO73DMLKRHCKP
C0/6sLOiYvCER1Bux1P6WVX1sdjcElm6pqXXBUhFVYKbIbIjpXZv/OC3Hn6tRLft
3ZRL8ovoRr82xZ54jM4iOpkyqA4scOHHHCwjgXRcdOnSkjyR1cxaeODWhJw6cfH8
jNn1lYeOlwli8sRkWytsJOMAOrxDg8u6nL3mONoLaS3rxmH0qxttl5hIHRhG8aJx
4h1Ph8O+vV61SNZumbpeGBBQTfC8AF+NWiG0o9WlgtF3fgedF4rb2GMNNHbQnFYj
7vu0uLyNhERjI8QZG+nNAQKXLdQBIO2aUoDELgSL7ezPtCEFRJF4W49Bk4T7Krcc
2o6mndaBWCMHbOxB3ZtqDA+b8DkgVzyRb+u69hvnEBBiMQdcowkh75Bn9oXaOjb9
OtHpc4WlisCQv6qs+f2aRvBvSrz88ImzS55IrO4vUUsFFEZGd9HEFNYQkpcp78z7
c7GKpOgPYQTxLva2R6Iiade7LH4TY+CuTpte4T6Xnh1m77+HCM7S2ZGkowSOPj5F
Q1czuUSCs9WEOmYZD/ACFx1ru3WPwjAgCw3u6nEbWRWtdWlStYIi48up0cGFm01y
F0e3zviuJ/Ek3bPea+EWKbEnFri8lmVGZZQ4iSzZyo/wVdrNI059kotzAVrjonq6
D2nxm1TeG1LeUSl9ZUfEeRnLeEZO/NGsAatvjCiPlqqizkSmtDnXpmKfC8MxuTuQ
LyAJ+nArnEpe3fIUUginoRxu9IOFYaULyUij//HrPi3aHA6bL4tRBruX5MEHLnA7
Y6ILYqbQXuHdqM+51ZtQiiLQmGz3gd4D6Flvp1NfjHqQWjfn2e5rA9IcBscliQ6P
tsM0uUuydyF/xbdcKouWVlefWk7jaAf5SpmES6GfY5gMMx0byyYYkBBt1AMphXCs
oU5TZjsfoKaSqqeUpnnJpdIbCZuBbgR1KbvRKRUSHFXsoBPjSDxPFn9kdtwDfjNP
lN1u4eeQtqI/IIwVnvqdc93/s4CVYxLMaOp+fSccow3dfCzRoG9JS9a+PaFyjnwN
jtljZGtNApbqSxdj8u4tOTcVrwwp2N1Y4SHvJ2HX1DNIMYt34ImpwZ22OeMtAmXv
r+K5BHu8zYYduHJCLNtmSfHBi2H18VsibEK9JRy6I4OjXrQvSNmffYUlQKiQoR38
mmfvQGwR9oETsnE7l7EA5LSzlPXT4KPrDbZz5D+MMJT39IjEwWUZwJ51cs66cd6z
7Z8XBSC5MOE+JlR3eaRBwSazeE8qp0MSwgm7cp78J4go1aQeStaRhbJoyguZgAFj
C8ow1A8/ArRsltvuy9cL2YjHRGX1hP0vfhPyIiZZXmkWbFMDYsQlmC8VjI+nZ6eY
HM6ICoHlspinW9QXJlDcpx/YvlNQibLqaQB2iZps85vN1BPWGl45C4moi+fFuNgT
aFPISG3LDzZjZ+KwZch30kkzn9lr8uLGaGIvqizmB/cYiDNaFp+Nrxix9iXA4+TN
vDivcoyq6pDnD3X3HjSd/2OsbAWeBVqsosCfzYrX0EqKmrhrSIb6c8iN5CEGzDPl
lELUqPrY8gXQqts14yo6rHcdlptsL7VqTSfgEhEMxP7v9mRhuJnSup0BAktt58aO
mT7PbU1hkEgve0F5honC2gs8+EK4ZUjQWKfUF1Xd/+bq4fqwt811SkpDfasFmDmR
OTnFg2QCDMHzhV639fW4H4AD/K2XGd94cIcGrHB8GBzXHbNIZi5Cq+BNZypMPN8U
KNjRTgqiGRaB4fIhZbx/xk1L/xxmOa57lsFGG7mTwivWJPm3iSlx6KffaY+IOd71
UvSUT0+AlsV7BEzs8Rs/RytS6FLcEpAQ4KzJm88dIqLCirht5qlHT+LRSsg/ukdv
RlxlmiOAzkoI5G/CxYWc4b1jwYPAuwul3MBU/TyjEt2xpndzqVUNW31SoiiKSebq
jRpjVfC4j39lmFRhfsxrXWUMIJ52FusM2avfGF2wUWgqplWgi/bV2M/WRyd0MxG6
4OP6ckBy2ZiPXPSsvke6SjP76vnvrOyW1vH/zBWHuzXKAbRGWi2qrmU949By1AZV
mrudtyQUPDr/srub+NSG+G+Brc4iYcGYbjvpGccbFZi6NR+rFyn3VoGRKNVAiSsu
SJd09Dyqn0O+p5CbJHOH3VI9lUYpu+FLJT/9latcxZygqc6GTvIyN3+XgdYAhZ1b
bEeRhvfe1TNQoTYhz6O+c9nsBKR+ht1kgBmdFp8VsAmEO4cNrLdHNPn6vjVcTCPs
v0er0I3y5jUusqpw0YPE9CGY8HDQJeXvca4u0P6sgCclMV2enNh4KSJuO7XXy8XV
0cQg23hSCk7ayQcx+69rNuO12hVeSZo3nUWgnILI23LhqVyqErEFbt0BDhPosfD5
2g2Gj/ICkzD2YFiBTkUtcFc2ygsFYH5cWekE/QPl2QiNRZ5LvXMfe06p/1yJMYzR
LSZeISvXLeViP8hOxGpl8uOw2XQiq4Vp5MYMUlztwTFRceYDWtAZ7hCwTFXGYgiP
C1tUfWhf+oFC8axipHeO52+0LSSOpURfHb38O2EVMmihRlmlU6UU0VlQ/sdx4BsA
JbCcfWldUPGyHFdzuOKRX7DjSfIZExUXhfhI9kubCl2g+TuLVXQK/usnVIesvG9s
HX63g3ifO/eE6S/+S8DgvwWa10mFa8dkMgkGQgt+lLTqbeADx/jsArfUQiOm9nzB
/sAZb7sahu9OHq4Q/YdOWriRUPsWxE3oh6vYqZ2BESTxX85c/rQCxZ4G/aoDqtuI
+SIQhlxW886wFRkHl97r9olDYZuTnMaOrMCYnkrwR21+G9zqOSA237RHIesPOHNG
hXjcPAfaoX9cf/JSyDsqTi2slUSSCTsN2qyWZ3NLivrzbAMDej+cLdDj6sj1R8+B
Zk2Im2AcwAvH+paCyCGWoKH7CovIbAIz0OHLc93fDNd1OElw/Hr/WRq2brvlLF4q
CuwOrzfYbeN/SIlWNxkuxiStClkD0oVfxyWZ8CGFn6sNjf7FP4tWinKH2r8jnOT0
NqiODRd9kNooTEM3kFXsRd9jTJUhYh5++0GAsZ6I/Mv8KpOfhzk/DdhMJTVLbUDv
WeN4TyVElBfnWkKify1/BCaNavxi7lyy6yNn9Goosp4j7+mVJiPI9wzAG1G7j9KM
JHhhX4QV6NSYjwZnjWvV9mQmKiS1r/vDJ2095zxWHjXDwM9uuEaT4TgwmWgU9tjp
FGokxGjzi5u1lFg8cta4yTNKfiiLu+Z4ltlVKXRp6JvbnVpzblvTk5ra5O8Xwcv5
oMtGv3HYCqmRcFT0NR+PpU3Wfo1yeD1pILgIpszCc0U1riRgzKJJGCMc99sKamje
CoMgNaYv8rr6CoIsvy4WtJpswZRo6xCndexFnFZMTaTtExGH8MibbMW00vysu1pj
Y0F/yhyQYtPbV0ZLt6tCnmfsGzJQ/1dos7DfrNLGxjVATpcCcs95l6eSBCfb3C2d
qsLBTQdNprNB/OMOF7cHRzGX4ccGAfPngsQ0f5wJdrhVahbVCuW3iC+4VqTsQHOd
VPWvH31c2lbRLXWvswnD/tRMdDALZSGWvE5+fU5A3mZBZ3TMmpdeNKhc+viIDIey
Q18B89H5//eSY92PixKg/GNKKEvuiZ2bAL2D7x4pnZEJpNziq4iII3uKUTow13a8
UhJsp6grbMtOThu8EZSEk0b2t3c6NGbVkFckkzDxPtWUb6oeVZiahPdVOsNY1ogz
2H+0VCx81/ZaX/hDitz1pFpjf8Br/dAEOlvF2vugEKau30QYApOROzZhlWzJMJHK
SBl5zdQU3E6L84HAS3NkVyyYO6crqijrEwoD/B4Wt+OG5YmkY4ECqUFXSOhesCHB
YlFjMLMx0CMziBykRlXw8ZHrAxMF2pyJC1s98Nv4JFO+XCieB+pyMwdpIWhJhPOP
Hwi7zAHAercIbG5dbRh0b1oJQ+raQXdCeTXwz9mT6vL80GMvcPb+KJX4xnIwbgkO
oc01Ttc7pNpw2Yt+s8KVolLakl6PwkDo6xgJPlDfZtnrlx4KUVSaRrHXd2vdAqhk
sQwnBTSWc/TZ6smiSHAoBTF31xRo+VsUwyUxDDjVPCLrAM7Um0WryuDNfKo1dvW1
uxWuf9oZv+A4VPSeFouVGVJOoYHXTZxNbE1SPg1VDIgvVsWX1l3ajl6sDpf8sOpZ
KnHFIS90A9gAK8OrJ5mDADOv3VPbguHsU6yuFYdssyFCrAB4x1mPaQJONJmVpryT
S1v5S8wuiEwoWXQwaDbnVSm/oGoQaneYUaiHW99wAUQuePIGrgNk3v/Gus78RhGu
FNYlqjdRk+gVdRuzrQ9lfF7XOkaY/x48aRWHis2P9wdvTFKEu33PMSlS7vCwrxY4
q1eQ1PN2TbGCwCri2zZUxtcen+qvNUHV2qpXDh/pdTJ8DauUfHZc3xnfnusMHdnu
ajCcXqZ3C/W91Buwu0llbjCo0dE0rESUOW+qeqTJFEZ9EkAghfgNaRF1k4wvTEF/
Pg3OkCztmdrCX07o2+Nd8CcQjDWjsShmx8+WzprD3fXjYTdGyoERH690e3gF7dFV
/DNSPhkL+X3JiAHZ7uoZllyYrO83fWlg5xuFYWLMOHbAKzkIEwZ1S+FgMQT7VXLG
rsFSeG5Ct6lNO/fAiilnAHOFfLOwb1UMfHNQVSkTm4leUGdrsg5Lz5kEI8CHNWaT
MWpAQNIb8+4+XIbYCrV6HThD/o7xQAGSO4q5KdS4bCP3R8uF66oRXA7ONdRLmuSV
BtH5Y2ln6kB02JpPyWc3yDJ7F3kG5xHv854kAwESNxv+IeF0SH9oCTi4Q55xQHox
IaXLEd37FmZsJnYEA9oI2EGNXlpvuzXzOBt92mvx8oKLsgF5gLn/YNxtxe/hnvMW
FlpBYXOUnREV1l9Hi7QdQ4wfXUc7DrXHHW+fgSL/dfG5/t+UYVIjf+SZifzQGuqE
rgZRjqxAaZEixX+RynlCV2sKjyxhLBfhA7ux7LfS5ri/e/AsF2jGEjWgtIER0+BC
/+ByOZB4JKyZuDhoHfK8xu2DHwD3sMyP9rHNZD+IBpXF7i0ICWGt77NOeGfJS0GE
XFFymDKjgU6Xr8YYsnKxZkusqqG7yX9RPUhbUc/ukhC2XlINAxklyfBudVC7O5TA
VgSYvMi+mLQcxH6MEHaYVUsPMemEqaKOJROFtEYlYYktm9gz34/Vuhjox7QDMuX1
WFM3Hf/+PJd3w2fW8U+6yjxJ2dSYotTs6qNKpI4fP/Q9G0SxweoCiNSmmzR1xN8n
c1MFYxK10PRaPrAj7m2LO3z3D7bQls1tlAM7Vk/L51sudTeumVzzFrlaNkB6JFvA
H/4SdetuO/8Lu3g/WKGgDUfp9S9h79hS3p/PRItykBxlkM96NnULJSMQt5cLeski
9LPS/PztSd6WdQ0mX2FigS7kj3JZW1Md1bbmn+6oxY59eiu6lhUSmwCA2dfDcUMB
4aKgvx1TqEZXWADYpwMq/DHvMR1v+qfZZPHq3eaiM97lsSp+zS2xWJVraNGn5lR9
6rLHD9UHzj8N1Te4of08hc5s/hyzkqMwylAD8M8TteeaLiN9k8EbwCrVhJAnU/Uc
W9mDKwehTWkjFksBsKPbsgx6mgKSzf8K3dAgiG16q5nTBsY9uilyFhpl/sh5SZDf
+BqZrADYIdi4hLNa0ZoAzgXyA/1WIBhWWMhsOI0lEwx8ygAehO6M/GA0X/RPVJwg
I4f2v5ybgR2nb/zCQwGY6pVbxCeLe657dCcLlZBk0dTKHqQw/rd4choAhrcbQR5a
BRDSiF15X5Rm7XV0icl9XD++7LHsCzfMbVcF9XyowJACCCpNzJhtrIWtW7cXQui7
ZHTS9UR8qhecsPfEvqXZqhDHXQXOTsnbKz/HkOejVbRT+ZqJ1itafNtYW8gvke+J
Z611fw9Auy3lRGl+NnFQO1ts2xsAdV9z5gN8chcTvS7ZWOwxHPO3o8PabQkl3wW/
Kr2QH1i+7egmMgQBm4eDRq3/BXi4Tv2rOBCB0HgbHqWWd0i8Pe0hmVncQkDABt/4
dbts9ZdFG4KI+YCo5uxNi663kJN2wyjMo6eqXVknuUFA0jNxk50fyHMuvF6iJzSv
TB9QngoZFi01dDRw8fHfZKwe76ryHJv1TjmchsPIxuBZcrru6I1+BWNORicpO6Nl
mPx4OEXtJ4K/Fl/m0SX1KE6kNnqicg+v6BdXtxjxP0rLGJSXFG6FKTKRmkRLiDpT
jNesy1RkIv2TPsRYwOJLt58aJ07pdAnZP0zVQ6QGM8O6ZFpuvcUp8/YP03N1KRQO
3phN54oNYofM78NyfbzEOlSnQI+Z/c7QJTAfQIdMdvKyCtLrit3agq0S7V6EF9+n
hCp7aesIMzbDzabbi7mDwvqgrliuuNt7xRLnYqNJP4UELooKrNK6wtrL9aVQXphl
TJVPDn/qLMyGxufQYpYZnbTcCpmx/Ik5JS0vbRXJfHjzyzYEAmKdbmI4vKpuZYrm
N7k5kUbXcQaXLfkYZ40O3fGgqh9IkViSmJPwCKZ7v3dsAECWpOs7uaSWRjlzlk1O
FhUl5t42/LBq6l2dH0x4Wcu0du2gaZAWFY5h9RMh4xkDlrKJuR6kp+M/1cYepRfy
gzEY/9+yd56TDhNNAOWnm+8QJ5C7pV5InQqu64oWS1g2YRbwPcyu/+Ls4jwJHUR7
W0OYPYKX0QrSUzv5L9MrO2ukWMkIpwt4FWc/M2ZXlDK2zHBoaidu++JXEsM8kEmD
ATWS6AZ3cYWHIB5E3/4PMvNAYVhTaZck+hA4n+LFrzLKsF+cUCBvQGjHpjWeSox9
GYNnsSLe0zgs5L2aZ5RO/w02Ru2mXN1txj1h3G6Tc6s6QDL5b4671sK2gNIwPWNz
vqI0+Kn7Uba1wkTokAFOK/R2vcmSZ1ncWkYnzjY17/dFO/lBUSqra6/owlTmoG1u
bSuxldegQz2J3joyYExN02bIBNnLuNWfNvZRYrQ39Dflse6ZA9OC8vUoFZjlla2a
DKHNyXPbf/UVaj0weyjdaEqsFvGcLLcP3VrM9GEzFELgEPqzcMO+JNPfbs49fh6C
a/mJCvVHKxLKl1z8HfGGPAuteF9+S4LKe/xGPX2eEoiuXipmFeOQvhvhKAOei/ac
Q9xPwnYKGZMwKOeF1OCvkib03/sXD+LV5pcOCtQlpMSLlIdqfq54oJlFjV6xXsPh
qrIIFn5HsA1WoNsE86HQmoYDoSjdJSFs2H8ZP+B9tmA+Ojmo/JXnx2CuWfKFj2YK
73oYYbcVsiqmdZM4p2FFM+FN7R3llrx9Z3OYRXFGX1aXW3pcD7vis5wngFkPGZFV
GsbBL6jgMO1JD8+wRaEc8cEdWpFOhJ08Yz9Zho24V62i2qy0BY7Em/gdMq0g85ga
K48PEUar9XSsbiIBs0bJCTEzId/mNlLeLFh6ootw6VeFlqb3Ime5ndsu20zfcfUB
d3Md+8pwr+98WmvSjmGVwE4QyM7OpiAQjS4gqAMdXVHTbEb42NW5NuuHj33cHDCG
qWbuTyEGecTMGHjmzp4ycAxA7Zt/dc6k1Cz7wDcx4cTyPHQZphv9beEKcoOQdod0
YM5IlqDjUcMAyOKGtDPRIzPO9P9CZR3AvwKUB2uL0CLSK7N9hqt9hTgEn7Lld4Om
NjCL9yDMBhXQj0MkTaAyEK0H0M/xlB8nZy4wmATKvQxJDyug3aBudKPvsSK+dpne
WcGKFYKabTSfIpD0SPW7e581KbnGwPByFgv/8Vr4ddnewAbhK5wD3mMTENk/URL3
AxrLWel73C6oltiPQJKLuXu1nmzgGLL1ItWpPLLsG3erHNZLVTftBTi7oYSdGQh8
ehJXhTGP/apWHs4391Q3tvo4vcFfQxQJFPLfd1+glfI/pFc8NQGdli2bU3g3xjh+
ciNTt0JN2YtgyGZOxpG+HSxvSm4DXnts5sasAZpH1a9paLck7oOrYL3sBnKCRehT
s1u+Jq2ZeGsecVfoUNkYwStcC/2VKU44ahFZMzIZbEWLSjU/T7s9kW8GBY1kqkdJ
xeBlOD5oCCD6rqI2wGY9in5MU9sunjneW0JptbBERpcnBm72I4ya7RHAO/7bnq5e
j8gIdFzaIQIEvIp/wrVDziinPBGfAxcEzj+UnMkKQKOG10zJAzkpPF2UVTi2wya3
GLW3+a8j3ySeRnejD7V199+QmLwR3AJZLYDjyv/jskzi3TtYT2g6Cp+FSfuMe64J
9FNYwB47NnzCVm60jg8bKulNb8Pdp1VlH53N6i2LbJoDXH4Ij0hggl/OlDJcVKaa
2981X7Tj+cddmDXvyIYvFlP8GURUs6RlYZLNVGXTW98RmB+CTvgqBOJfQvbWakPo
AOhmxBXjXUtflu0JtyA23V/Y7Jh0haqQMcpUxUhkHKbMaN7hFk1iODFCizeaGduP
KQrUVcFpjtzv0DYBgFMZM1JJIn0/hLhOXPyXkDdLFYridFBO21nKKkQcugGOvx8c
+Y4cBz3dJ31XSwrHHrmN+nq8PKBgIWSFo4lPawzQcG/ixxhddBn2w5YUwAnwx4j7
5Rc1CQ4lLEmJqB4QjgaherELSZMzPKxTK/L5xPs3KF1AJSmbCOSxOEViKiMsrqHY
N7NT9Rzaud7FQh0avM9sCzZbengAnBA9c2PQEaeByxxG13r913rTVdepc1AkDKOu
UG8fP5WVCssDCfhWUj0qTeyHQrYMP8honkmv6XafEG9Q4suvOrZNQcCb3/0yGPl9
dVhL7lo5X/NCP+VTf6Of2FqLestaUF0AmwVbR9Mbu3ioqkRK+G06kswwrfBysx1j
75vcohf7rna81n3xgSTtVzytp34vtztv/UIOV32cAKXISdxD+FVmaUJqNT3/B0xv
vr6YbnD+2zo9FqFVwFSMeUnQ7QwTy88jjwG2YiUEbi+MAXDRRnHkYcyH8ay+uflR
ajtYoJSVTa3nnob8UTmeykytnbcT8KuKSa4lMwjdXWqYxX79U08TtQlhAPHEMzdz
5eURHSEN3hkeDxao8m7WKaaA4/JrL+L0eHjtCjWZlb7PL4lhdk42WyGVasQtHEbt
d9BzWp1a/NTzWHFQ6Gq0x4ZV0YicoIcs8NIBIj+n2WICew2YFqVZL+ZOQZ80cC6n
m0liyxTgSW+e2d6z473GbIEmamemipDccUMhzjixD8PFAKuDI5CjToR8sIUVGv5G
sISrkq5Tos0IxexxC/ZkFR321LwUg4V1YzzgXJBqHaZEk1h27APV4ydFsJHkMlj9
mtFI55yxMBi2KCLB+GbYPgKbSuCuJ2ntrdPca+mp5e3AHga3pi/irhLnVr+Xle29
uHUILVLgdRflsr5d8y2iUraIjqBBwCVmMY1p6VaAN+N+7JsrFTPPHYr5WoEgjj5x
tZfOoPw8iM65q9joXjrMeP0B1wSj/r85HYaGfbsMJUkcBPpmAwU6EByPI4LRgulz
X8uvcyTabZsI42nRRyG0A20e7Hc138mDzbS3H5qhiJZwmkx82VoFNj1fV65fO3f5
vdrtH06u+egL2Zflj35bHE1UK9ko8ZgFH73uBd1WBGgIIsp7CTZJbP5XTn/SXpO8
y/y2jpGOdTxcCOdUReRKNpISdhorkPOBTF01eUbxCqh5pau1ceklQAWj77SBzvs1
OpLYkjZf746f+aH3dYh3sFBBUseJL8MaPs09x7LLcJMb/4Qry3CNLEqe6odHNflt
iadM/fmi/wRb6oyFPA/TfEYUGLX7B0phI5XZhG3pnVY6C4laLrNJGKBqQmvRSw5L
hGjGcNONqaMaLYTvLMjhfPE335yJK+3HaqRfEz8dLmKgKxLdWxZp2GSTDo1KOVJ9
afs93z6Q6e0d9HkmA4Ypt2kLcpWv52bIr/e2huvnjIH03RIoQpRB3h1laJMBtAI3
Ad3GJbozPZKBNzJVechEHXJ7urSN5Jd4x2I1CQ81hc3X1kg94ApQgcf+q/o/eWcc
jveeQxo/6tW+Ak6T0An6xhd9gF65M8uNIhh3YFv4DV89b0smAcYV/R1cJez1BpAI
FMCXfr6hQycYFEB0aQVoamIkCQ2RcZWQVkAk5PYgBD0P8shEmn9lWgzU41cxHoAa
g8hx6sxWCi0K8emvGC/ajlcX7cuOFZH4qmao+XRejRqZSOcH5CnQ/kt/LXU8ePOE
OEGedHQcps1RTvYy8fjfvjV7HDlvx4naNbnwel2gA4sJr1WewcQa4xv3PFXJ6A6H
1nvQUm4IhmZE80Qy8ds3UCMqKQ3A+agWJ25jO0g0qB8KdfbSNqXrWRMZodj4uI3u
Zrv8bkt8b4ttgLfAuiIZHUQgr8ERWzgAjVeHi1fCgTC7kmIQXTAHqDweR5z52z2Y
SOP+HstWm0v7uWN7qbjFng5UmlQKtz9hjrTdr1p29Tt93N4jaV+v65CjckExWzv/
qGOjfRjaGMcyEXU549w1xRpkXD+mQRUuBkfY6FDJjpSBgIwx+ifuhCBPUq/CUKvN
zJH4o91zW7TdM2VLpt0FWM9fpwk8W8GcrX+g6ThynKkfPGKYnPMKuLzuODey0Nr4
A5qNCtEPOqxscVYnd9ViZQhHQzDUwLe9g1YeY6+oE0GOZFjIMiw03ba09sLDtnDw
3xfZk7d5G7lDtb3FRQXos6pH0KEMVxaQu3BtdI+utjqsvHT96z/6syPOL9G3fMck
0HvQDh4pc+avhRD0bVMm6gvw8d9FlGP2XhkldN7zdRBSmqo05CWwgFjxegNoDyLr
34QDJVq1j1pcqdlo3FlCAXx39TPwZctQOFDWUdrbXINA3VpJI4hpW2ietDVAJwpZ
Vru6plqLsMqrMnf0DHW6IBdTkEHSztll4eeqYsVOK6BgRnPUMPzbXefbxcJenKLN
SQpYhJINH6F2dmJck0gAUwMPPz+0vW3R5TEG1vEtRnCk+i2OK0CryS/VqE4J7jgt
6HefIZXcW2PrF9An2a15rK3kR+vCsxURxkq8WOWr7KSELb7VqLM/unMasdpoRNEP
evjJnpv+zPUlZZdq2W8EaF5mEl0PTcMaBNg0SD3R8BkW18MWNhMzlZPfn0PVeFW2
8xdp4fRQjEviU38+IOsjYc8eEg8Gm6O2dQepD8xYcFpvkM8Q1nfT9qiMrytmaP/y
1DLXN+3JxAqFahLzXSl5BCiw563gaOYPet4+RMT9Kx0JDD50sPW+DycBz9ljHcuX
hqgIt6KwUWmfFQQeQNa4jPbpqKF6Bt/EVPedak7oTXyMeaBpVqnp5Aj//94fNk/y
m6l2jgODhF2tU2LHth8ZWO3tJqvBXaWZuxO55V+a3Ybj9wsgcHuAtIx8OICquaDV
HSv9RW+DLq3tGZ/p30f9uja2Oe0x7fW0f1MPYWpagehniEGCuqDICviazn5i8ef6
C4ijk7FHKMWc5GAyGxIsRPVtaN3yTMxMKtHIgMSB2PrlDOR7PMbawnEy99t8N5eJ
4U9SxlsWIIrsHq0Ksh3GpruD1vn/BuaRBX+O3GAtf7DCuTrQLn59c3fHcFbnS/u7
zoYU7hqF/3+YhmebsXpu/OYUIjaET4R1S3TfBxRR1XDGaWryRjGsxe+rSgLFPnM4
1oPGzjW4IK7diuTfQwo8IMyx4AvrTIwMj9n8fqOMpF5SP2ph14zD7bS8eIDClsj3
LvRRyCc6IOEzCNy9J10ZvPwqt6ceK4vtKZia2oA3wPiaYOGh/wtAkXTUEAJUdE/U
Lls9k8V1+7e4+vsozVknLCXrMyFFSvvbvuU5myWDR6tfIrcwB64uyg1L3VY0vY6Y
mYd3xm2kuXWBuZSGm39/MQ/gssB0HWegjKkGTyML0Sc6tkxPrY9/u7QeLI+BhDiC
AVH13RUBUDU3fbXA0oTSnMSDkpRrNeZ9+lWNaLFnDbsP/s9azDQdTByvKNiGggso
dikcYH+2ZU8FJsn7R+bhxkdFEcNLKWN9c+B82qXgikPKApwzHKlj8xbtlfh+qnPL
UsOVu+gZR8e9Z9wG/9GPPUtJ+TWWGH154TK9DQncYwS/GpSOh59+Q7tPlaw413/A
A/KpnK54bsJBt0d0o3kROoFk9fTzGLoD5TcJTsrc8NNd7oUL3WmmOIC3jaELnNcH
ABbHpiWe2HMqmlwQF5EsWp/3clYFiPjZY9+d2mYX8bFAndzuH0fmfaNH6ZXEGdDV
77yGv5bX49dBqlrbu/IcAoaNSJk6W6duq34zj6TkMhQ1t23cO9cm3QR0Xs/7hDZY
d94RfUvXX8xAZz7/SjXcFsMTsZ5Q79Euw/WeV5D5dbVdBr+n6C4MtuU6cI0BymYC
bvERNREY2mbku5cKcfcqe0Sg21QxlkNHYlS/iID6u7pgvw3yjXmtB4ly/6P/14RZ
ZoOkI2rNM0M/798C8eJLCeeDiS6fPsCM1Vqj/fDiV9+NyeJg5KQduZokrJphDgxw
Os6UkjYY6+9wDnVXXTABvWG+Wq5utMh4dcbBsDIP8xL9a0qQDnjoSUhg7WEilVKE
940P3gUzurkgFLNsf4NAGACnYjpWEAWRfgREvjDH+EwHqQfXjrFJptM0/sB7xT1+
FNC5ac/jq/aF6EFhD7sU5V1GxUnkG9Nd/Fa8znYAdDm9w1lhu+IfiDE2LR47Uxa8
kXZBRV6VmXCAMFCJPCQL8AgP4KX4vsTf5vV29ID3C4uBpUus3rfDpK5WU3oNcyKA
0z6Q148Z/ncQ3wlcCO9oHrgHL5cnkxmZ0NvI1iqMxRkFQ9gMAL402aBPT96wVBEE
S2o9LpRrKFPjymZxi4UDivuvVC1RBYCp/b3kR9MKeom4/eeM+Qj7GO36RoIA7/G0
SSSY4gxmLRi8Aj4yxCvr74aXJ/81+WyWTpyKbZKQtvm6vWYurG6W/eYvhIQDHPiB
7yqhuWzGio9VL/YLF7+i4P1GzM7bQervEc9zvT7mxi5Ogs1+1/9lLslB6GYcpu3q
Jaty4z0jybS2uXeE3ueXkz0CKE66lGxPl/HiWklwj0gYGjXXvJw2C8n7wFofHqjl
dhPz2o+L8o34CnjL2Kq1etwzKi6G8TYVOMX6o7Nm0szRZVDCm9PzX5mQvDWlBl/q
w5J1wBXbizm00Zw2pLVCQb2WbxO0A5w4RLpMNVIZaZ0cw8z+Mkxx2y2ci+/r9d7i
Csx/jk2XwOSGDv94weAD6T/leBjsX+BrfrL3CWTgogEGt7u1d8DsEj/nhge2WJn4
q/8gEZS9AEWU0Vv2zMq8uMWdQ7Y8ONdm0ikJAQT246K6nh03R6yXohPggnQ6Sr/6
lk3H+Om7Lh5ZvIxkDcC8NApIjadi8VDJYpGbsvUTUmmyiyIFbrbro/cWJWMUXTsa
WmisARIELBwaLgPDu4UX54PdzYrV73jPs1tbYCCpp73SqS3uwgF7E3SrLwkMznQK
nin4Sq9Seyyjdb+myFFZcDPpazoC1x4mLUFL+KdJS5j0c1xdhDIZ7IWkLTy2sKkh
/TWt7RdWq0S2LeRr4NajFcJqc2kAAZxouK/pC0LFWaJBH5kY2TGL/nReFgd1DAj2
Um2cyKcRWcIa7TmrUbuMbge0ocMzAHZ/7SjJmlVwfuafkcs8wfTjUmjvjBZYOXNJ
keKW2H1HWmj0aNFxrf6n+cBOHGMjxMqXMuv4lE9CTYHpMhWZMMkmj2r4ARcZmzQt
DwXRHIug0BCR/14y3NKUYuk4VAMbstouISoz92sKzhxtrEjbIdDf6P2Shch5ErvN
nuZbIEUAOoO53m9Hk7ndexQLZfUsSDSfez2CcctBjBijiPvWSv0GIUurepC2a4dl
FcRUGFaHiBFcSVN9Hwm+Ytva47wnOWgtIn+Vqc/NTFMSOJNDtyz57rE04Al8lpiV
R2JtqfRurUhlyMBNXnH210GsdZC9fOXUGTLNpcseh+ISHNXl+GJ+2psyC1io6Kq1
7gkN0AvFTnAaIHPqUwxrEgj5kmz0ftGE41g2ZxcO9d3+M7Q2W6c2T9nmhTI4BoKJ
ssMvPkCoycZm20TrIO6S2JAXIwW6coorbJWW2vZaeE8WmQsOSnVfHLHmBdiP+mj0
7KQrrxxMnSH6PojMmwceoE49ZIiGEIgQd59FHa3/wmXHjfZCBsJCi9dr+v5temq/
SQABxv7gGP8ukfVb7J/b7ikjWqeRd9KuVCDQgmiJ6X9zOI5htUxS+xL7fLt48As0
nJnJCzWqtpmQ58SU6YRwvnlyXWEySoA/iuTz4X3bUe+cOsWDI74PXGV6eRLRby3n
zDkvBIapVcxn+xSwQpQq5Od4S9T+rmhJBZArJ9d/MN9+pAls2hPjQNF/y1LT4egH
+SIdyN7ifeuOWkDav+JZ1Rvpx1h7Lwrlm2p5SFtuUyjc+5WazVws9DR77jtf47Cs
zc1oI5S1qOvcbMIKNIRiDxV/xxN93zifGAJ9zYjzACee6j1ZNIcU/WbrJFfTBq8B
bt1STQu/Jti4i13YgRGDIdr2aCuUhCTmVHeTl7ZTQMcdwB0LfcEirL5zmknVzMm/
sPLeTqY12xScKKwLmJI8UTK69xoKj18d/gfG/KNIeZwZB61cKZH3Ssj0OiwikMo6
w3DYstu/D++NfXRDcHI5ejCt+JNxiRe11dNeVFddX3eM8svlXX4Dgc9XHuAZQ0jB
jgBycurtUmK/L/iG504cYuBPruev2NF7PxZWorC63aRaRIHStx8ir5LnbyrCS/j6
CUfPvdgjaDIJjr0Eqlnyn/1vk+IzMOaJutFIS+LGX87t68dlRH/9PZoVg7pwUR8j
eK0vkVTa4YecbmJl+H1EOMN6nksHQUTEz1bxLx+KuV2RZXzGOQsjRzcGSa2W45ZA
g2IJ4u68D6M4Z4JdLGXA4lSU/shMXZnRaAynMZoY74+Bibc1p7TzqupTCyGVXtBs
uOnIiPg33DJXEVUG1HYEFY8Aleri4/aUuNWJWWgIQIWyQnABFEdf9AIPqaAMdfsP
ARN0z5A2N5oHvMjN+JNhoPM86i3C0Ka4VJaN1nvf2tiNByHJzUa2z2hfDKUDD4Eb
+SnW6iN8L0VcUFqY8vQm042PqbOQ3ES6yrjh8FtwfojHKgWwHwAG5S0aspwdzDJl
4+xhjMbjTUgXsfLcaMmLv5HuetM1/y6xB+if8Q9ntnQv+OjUuGpivjhvpdjBP36a
9Y3RwkOKOxOuxFjl191lJ9TbPzulU+fO+wJRBefHD1E8zFViKMuIG8su6YopDUNr
lRWxxxhlQU6T5f2I4JxUP/LVsVNjfpiLqQRk+v2Yt0R/hsUMNgxEeb2eaafljNKA
gchJXRjRAp0xqUbta4qRsbn5pLZbpRA/NPIEgtL6XfJk+jPUIwtJWwVQwE8L2CE5
wcBGWnPX9GiWR52rVIkk2C/rKooa58hidBysoYiojLqzB//NyP97CEyMZkjAHsy7
eEQ9m9Ug1FtSCL1KBSfzMwL0mdRbSxdb60BBUm+ttxgQWYKa1FiW2RNl+RKA01/a
pYpn3Yk7/NEu1B1H3CsYyz7qeiyP62FmXS1lBfaKLXJuJmxl9sVJUM/0CkwB3BOX
bX0M1wbr+kbxQP49XbFYCVbUF+dXgEvvjldsE53gpvEEUKbg94mgrIzS/q2dOA/F
7EaiSZ/mp0qe9asV3gMqXshzA6AQjf1I/z8hbYWnp6mQ4erV6ccnmulgtbEA6BD5
mD+pfHDJA5agZK0++QkrHSctAGpspxstUIsVZ4y+vzs2LI5bj6UjciDnbK8eKoZC
KdCCWAu1jaCOVV25DGVTXq3180Vkf+dMeV+CBRljudgTjWPeDh5H3LZPUw1LyJcA
oXm/Rf2fSYVn8Y93kFzM89dXmPy95hrGUJsK8PyIGdYpTLy18hw7iUmnzujuEdHJ
IqIUummiIB2UXo6VmVUa0CgpAUCpKZP/Cjhg5u9AbUXHpUmZDrxcKeC36qAuG2xl
nGypsYR/UV6D8V/91QVnPB41KczmdL97bI1p1yNJ8QuBkh+jk/7uB43ekiHNRtyw
35e1ex8jH+2Rhwd+DmX+OW1WSpz7Xnf/20uwpFqunisBI17Gr4k0K4NIyRX4Skxi
F+ALvNWYmrsz0MKyxTqG8836ebno6rq96UcpgBVrje0DyDGlJ5jNO+Zv2nBFVSXc
BJEuAL2vjPnv3iQc1ZeKzy0MzDLaEf54AzP4Iw6uFdj4JTsxRnfFeI4IP6K6at02
qnrznZnCml2iteaxlYVycwyExZNKMkI0m5viPurOx+CWEExOssoOWl9xz8xpYAlg
dyD2FQp3KXtIanu3ZlsrcAChyxGfkEydhW6geW/XM/tpkOo/Ic5mN2vkRxRBIQb1
Q9HOcpqopbml5HjX98CLTWdhh4BQFjaVDWUj5nT3v2Mi+i2Q1ewpIGy7m11/JwXC
ZsCCjrKdc8PshcZjkFnZfIud9E+zCg080v+iCxY72vMfCCU5Mz7QVecaTT3sKfOI
Jx2xPD28ngmmytbm36wqyE3qTzxnCbtJ4bQj4UjtxnPmufOV1uzKjPa++yfYZYR8
SCEwMVNB54t5pSWcmIs9Sjq8K2SOK1/VoUSVJ/vaUFE43MDLpb7/NgMX8KJc1M8Z
JbdR23pkPlplQtnOtDHjUa1AzUcAHbedw/5phtjb8iPS5zR+wIQNFExwE0cGdZnH
9bBr2oUC70zXPAeUoeoPo/SgLfsGhrTvCvCMO7AGgl9sz3UN1qA1nN66JRJWvbWe
A0rvNvJLz8nDZM1c1dnTYykxAogSVxGv+9B+/tOog5aNeQ4tBrW7+L1dswsQEgsd
ZD7ORgCDBg+Eij2nBNpI9gZUP3u390sYcBPF3bneLtdv5rVUeleSFQfeDB983L6H
L93ifTXSzWC19Alqhd73AKJMpErBtM1VTn7Iu72EXChixwjEmQ+bPF9PlckSRjtg
ZGN0QDPiC6SHEaoFkxFQ/9gaVeF6fBFloq1A0mcn6ZJCNUDbdBFnLwEjpunqcVsw
IE2oywxhrU5EhTwCh447QuQN3D6TtdIuUEkIS674utWtnopKt9eU9PJLSzTR1fcP
lhH5cSSuBQJNykcrK+kTnnBRscdeTyggY1YhGU2sqH/tmHAKtSQR7HCkWsZzF+Yu
6ff03KYnzOprxztyZIz7RK/1Utl+CTi2aAPcvRuFBD42DX5OUPCucaNilwl2VXJ/
ZSYdoc8UECg/9kR3hEG7xIdNsZ06tmIh2OwLpu+ai2HhyZNwlu7yBUja6Pn7iKsd
KI5miKdBqvv0lINysXM81YfbbEKRMYe8CuzWPB26QwTIWAGPcv80OTykbKChCpeq
XEg65VaU3QQYV5Y3NuGwixAiSWsjMIMTl+kJ2PrgCN5vTpF0DyW3JrYemnjVQUb+
cK3LgkC72wgSSWaoGpU15q/EZLVRMw7f+L0L0aCPfFMsVZHFLE5KlQgphxr22n/L
PkSb2QV7jrf5Fhl6399XrNzgfgPCOWrsLRa4Zw1vNamUZi/9K49LmSNEiy8jHrF0
xqOugNWYODvrEp3TVhwf6QqUIKOPKhB/Ex4PLm4FstfaqS+r5eJ261OHn4BAjEJ3
cOui5hjsIAT8gwGZ/UCPbh/Zt3m42fMaN8RFcqKGnGtnQR4dL/2HrHia3WPk/nVp
7Tt4dKcgUw7eD4aM0Od8BoM6NrGqmO6z+1OgbYPsiNdN7aWBr1DPLK9KHhBc7iec
EoygNJ8x4o8BdsQrhSIQhZLV/xGzaCQfSGM2ez+D3j/mMBREesvd0IewsDBHqhcW
XDT64QVetJpX00Xu9BD+tmj9q5aCs3H9b4c9al/Y9DV3GXdTqCjSoHLREddnCkDS
wZr8HK4c0sXuVNlov44B4tzGq8JN4xhtQvCIOKTLzPVhJLoSLD9WmZ6X7N//y/Fh
RfTswZztzh7K8f1vzEZxpLCVneRqBiLKeGZ9J/bNuCQY8jsgdXDSOAk1bA7iuLcG
tHY+IkydYRpYzXcPyalAZyjyo0AGOfpX9qLIs9VVoioAkAKvt8eaYE74TVb2U+Af
VN+JL29p9Ra8RZ879RMcuKQsbWq/ssmb8SZKJPsW+N24qysf9Dy0XVNs+1zh5F6m
7Eg2DGlUv1o98iuUGY4rwEvdo6CFWc3XjYDBgNtF0BKHsENtv2osckMSRmBJtxzu
VVrp52akpbVX/JhDBQZDlUKOVMWFqz02IeF18tWaobmm/ZzRcZRaRFg4LQWWsWri
yKu5U+Dzz1LAAJz5DYR7SGA3HUI2wInVWKolTnbqskc3prGehogSW6d203FlnU+1
7AgM/wIfwAC8LA+ui4z6UXB/G0IGGbx4YEf1/9zmmVm+duGMWhQR6KgwCeyRyzGY
ofB22d+eOpWS3OgLrzd/qWOoLh7flXSlgQRCPoUolJspZjD13RtVFKaWEgmNbi4b
p3h3b8j9rSIhgVy/57NVFRAYVrsYOMRMamr8fFRwCOk0EP/1zQuiRbfS99+a84Qz
EpkjvMNXsb/vX1N49d9uYjtwIsZNYuW5p46WbHk1I89BprMHxCwBbQiiPG8oFtEE
8asAbVXkiuKS1KPC0dQcnqQTKhMyOIAkn60GxRfDqrb62scImZ9V51N89s4fBXmr
iLSScsqg0ZZ6yTqfRr75bFsy8U8cDxbfhurN95Z3B7MHFSx/l1n315LBisnZ1rvQ
zuCGwUnaPyRzW8sMsxxI8jrULaNq8Mdy6sBK0ajXGt6uOOvrFcYUfWq/FB8E36v1
oq/E/VGCb+y7A4qk00yeSw1e0awvB5nnwUgaE2aQcsSEqY32h8SmxADrT5Q/d7AZ
eR4y/pi0yiI4mihD5D6EIsL9plhAAp5XzEoSUhZTPyQfZc2jLme1euw5A0lLoIef
GLwrsCfAHFNAYOpWXj+a7eAXEGU4PEJwuzh76la+uumybO7XlKJ+14OEpSQOMoOP
Knb6Q7REUjmfrGMqcvYw0uuCQItBIJHQ35MTEkC9dkMA/De4RNzCBhbB3xqaSxJi
Q4yQGibGWJjwyLILA5OeaFsH36gngv755OrrAvhYO/VtM5/h2fInCock4rCPIIsn
HUemGE3Rq1fzTQkz5IB60A4ZWpoTD4tHiuc6e6fcej8BghIiqYusyoMoHkLov01Y
BR2ukh//3LgMdUBmGoWbZbmOjreE/Zyz4kcJ5CfwXHErMo0eVR9UuHjZXs/3cZuE
CP0uqnMpM1F8Y/m1dEWu5hD6jerEsQAh2txt2NpVrL2+oa2jJripFn5ecXBTT2SQ
rIykS0V/yy85I3fPDEqnEww0yP01xCsodNZJPdWjzDv487U+IiSwXIbkhvWgc1e1
Rd+/qphv4mRiC2pG94T+hlpCAfh+sKrKwc037I4F4h3ySNlAV2FmSSxWsvNJIgrZ
wx9ljXRksxhgn4+/WHP+92dIfgpRVI+OMfZIEe+xg2uMuMCnJZQ1Cm8gzRgbVcg4
GxjJKmVgf6Df/bpqEDMQQI60BEt8Rar6B6zCuOaEd42nB60d8vuOgj3Zx0wnjPvT
O1LuTUFWjwM+Q7PjzzEO8WQpgcZeU/nnlGdEsmo8vV88RH0N9Pu4avmGUQ/JvCG2
9Nd8PRAlBSaI2vW/u6GZAfAuX5RXHz+J+o8ehaCMBQB7NlqZ6cwYmuGw0xlzJWwC
n3IbsBD+SCJfjb6FHft40zINpP/IhwGneFsInwpJ2ndbxp37HRSfFEdnFFh3X/fE
PwWJbN0eb2xCc/JRtsl3tDuvQX7xqWyL6Wb0so3/nYWzhbtBKG9dLb/J8q9EqtkY
6Gd6JGV9PygN8X02XAx9tnMHPRco7N21UY1p5RclFgyZll0CUxz+Ci6dOuZPobUL
yE0GAndi6hhwACUmH6wdlGukHIutDUDplAbtfj73ORvdqdXSidiwWWz7Fh7xDDBC
2yZUn7EDB2oRBdJf7nJOPvx3C1HioRLFNkqJrA643Kb0GHfoY9QbEIqnKNZq3CsJ
qv3rEKmSKspvVanLo8oaHJjumeuKajPHhek6VC0sE0BciDaKjYHyys3ujhOusE1n
wzaV8gBDqx7qFFcqDjxmvISnVPcbgpgZBuCqxHhQpKf/OMSQuxZumpxMaKNyoYn4
s+SOUV25mzvzJP9OA9mA1YYKu/egfQuL7+iPBoAFCgBCZTl8K4h66lCIUdqd+Q2E
lqMb4nZEAsHYGq2TxgHNzMlUr9cR94O3V7uOYUoAF9NOAaPZWTRaJy0m6c/R2mPU
TayrwPCbqqc/2vy596VPTH6NbBVMthTOV0K5Jq3YgV9nyC8KFqaL517MGHiB6NZJ
brNNy72m7RsWVUsn/i8UQG1LatWgAZrhZLwVO7CQzPJA1G6e7X/PyEhvW938332q
E8ieyZJf8ki0FzJhINghu58ylcX9ZP+eG3YzpHfZ1J5Yf9EwanDscQcAlX5+YhvE
+NGtAKXCwpFL8BoAriBWxw6of6/StrQfx/6qY2wi8Z2CRG7XKaDDJqnDAkI4b7Kp
iP7C15RiZmO0efxeIVkkdtjylry+doau1c7h/M8UJI9l0pAJEwdkAproTRblwQe6
xDWDQawcAgq5dmHGPqszYsHrlkISkCOdldCe/QRmsV0TnFMpUYVmErMlocCUHj8F
ScpZS5d0mYEuCSokiFMhcVAJ/Iap8ye97Xs/fncELREGfiw4efaar4EyrkBAZ0pr
mmGlJETa2r1PbGUgdFH2BwWmjxH8lH/ZL1AhdoNrKEg/k9V9mWLkYNU5RsGIo63E
s0maBA37xMoa5Z3Q3mqUcQi71dZj6okOlvjQkwZKGLJ9eHZRf6Y3pVHotDAfXLyI
co4TWBQbXm/ow21Tqj33nuK5FVL9HSJgkddil7nusF+vEuOHphxX8I8uLD43coUD
Z8jnmGOMQ2IdCTfvI6KAc4jbJ+HdrV8FQfSzuoxO45RHCPsd2ViW1O5XpLIcWFMY
qKch7uwQzMb+IplMqdA8PPURiTtSJG/rTSupxLVAFRqhsMcr5pTv5WCA8AGXLFDC
ZiAXyVaKva+y06N1H4TwpDnQQI03CaU0vaFGr2OljQiqu6YDGVx4jGq8yULozDfn
gvdkwE8jxQCZ47UyaV4SIETrCEOh+VbmPAkdiObYTzFRSQCWDV+tdVljTCe5xDur
5l68tsioUNHyMqcfeMi6yi4eVJsiH2Xa79AouMEkkipu1YxJsbh2Daw43En1/PFh
78r3VP8qED4wtLyXgYVi40jumz8oZBDXZNfof43GYbcx+AYyvOCdQsTdalX+fp4b
oYan+ooviKXM89qf+wdHlo3AGckx2m4+v1T7ImGchgSn5T7K2sPDJwOyYypznMgN
OOZvYuVvN2L7LfEaLp0uFspIQViPRO2PDVodrqdYIwkCf+bs72hNnbZ53gBNbW/4
S04MsVV8Ln8cVLeNlADOt+efAUUHVhrNBf5/VzzwstgfXwGVti9nLk+3+icbH5uO
IROyy0Cl3vFe1ViptMD51S0fm43pwlz69sSxgn+75uYOLGs+iggUSqpxtk5lKPuf
H4G8+8tgMuL1+uYNAPoFRl54M0GNMJqCpC2zURpUOZAXOJGxZozaDrkaSeW/yGYX
PlXGGMzuYoSNRzy23uzxQAcr7SxEefDWHOonhU2fswkC2Kk5Y3SXe+yFv0MkkjEY
3RNROR2zb5DtshLlxFwbXlB8PD2H6L2TVHfbjH4WLtKK8cbR+zsB0DxZcfdFQCvn
qZkWqIV5/Stcwa4WJBV/m4wY7eDIZjxesAwkXrnD4rGrYPRoVptki/6RtfCOJQRL
E+cwo+Hth8Jx2esjovUZZySRHNBdd9AbKUsdxMlTQ6ucLTXCs9K6NdOq+eLgd/iD
duzxlxv72mbXt4icksbNxPbvwxXYLFLTvO7OYiOli2Z30rtlOCOisFQ1zQgXREKV
TiICjd5WgsWJx9t4EUAb6xXRmLmnvmX+bR2NVtO2kglrqjThq9ekFCGDKIFbFLx/
jwN35eSOtPXpTflrnqUjdwoVKy2ac21GxOqHRCwnvK691YlfDmL1hnM3iSlzywzW
eI9NyFkWSCGQedQD6RkWmD9zBp3kmTVn87ikyxSPhhQdZTPb/GL2sSiApnnOw3yO
TMFrpT91kndkVHIz5mNTQ/YL1r6O89X+m/uajcxqWXctvpRFj/iZBeacb9Wtx5rB
sbm6wwKsOHpyT/XVoVz3ivQ+PeAmjrY+9MtzVdwL/4XHv2G95JNEmCmyF5uSrvBi
VRhDM3/T2H8TPi8SjWY/0T4/gPApSXssX/X6PS8eKF2wVlk15ztfVTwkTOeULt3E
BIwTTsJnc+n9qUry2Zp8nNTCFbVgajWElHhhMPuUrR4aTH+fEL20DEsWx2w219Qw
vXsF+IiPWrzNwAgZMG8t3e2DRob+dmwMSJbPnzwmFYU6ZPx30Bgdbm4Yn1CVdji8
w3ZY5Mf6txYbLv4RbwsleKaOsDryNQ4tyl5cxw6R9i+C6kPl2G+D+i81HM4JQQ2N
cZG7aorJiP05AtM5ZGTAquY5dM+uAuwntNJReiCMQvEb3M+iZ45MJP6g0EQgG4lr
OdIGX99WXuYFewWnOgtwMicnp4YiTT4nitG/2wVeXYxWwgKaev4m6KpPORqVAhDF
ttB05UaFKrLhVqMDiOfd7ldC7BJ9uRA5lOduGuIMmtcEz+FEpehp4eetyGRbxmSc
WM/1mQz02kHNBNwcdkcrZVsSmyLPVmBnWRr1q77voJ+12FxTaA8CfulJSlhYDLeN
KNopa5TgId9t/pjMKKDdkz8krgIQwTMOncamAL6HGsz+IUTfaXTsi4lvWd5KkAOF
/f2CUzAj/nXtfAj2cB793P/Gyr+J8RfOEcfDCMwECpQjkzYnIp0Mmhoo73NiOPF/
csU+pMRIXg8OLw9VnT24pp4uGeh2aaq2OrCOVzTSD0zkVCzu0HL/zXtoNuni20Oa
dcJXiMEaV+TpOW96BBbBFE3Fwfpep11zrcb3/Pt5E+mN/PrHcDcFRdZnAJNQW1Js
yRlIJonJuY1lhdG4egBwNmAyeqpqU+dCYVWTZ/nU76qLM/vVi8XsAtZQY5VUsBkm
JWfCvTOMq14f3o/lLcRK0ho7MI0GwACam1E/VxVmwTC4kmawUiRPWHmN4C3LvdVK
dz8NNXsyn++6khBwwwCcdKgSY+Q7NsZEzanlh4SPPKu6BdyigH51s0tXxWyxHCX5
eYK5DA3Jvb7TrRo1pPonmLF21Khu7RAfziHkoSBT7S31UMwuACa7dbv5OqChDWpx
zO9nddHR2+kaG5sNrr6qnUyFED0XMR3GLPB0mPksZMhlMLgtGCJORzkg+F3ZLx96
hMTW/+QA6NFvuewgRn6qidhV/pJm8RUjjHHQENghCAlhfgUiyz6u/tvJvDPZexBX
6QtiYHjYb2kIBbSaSdEWWnliE6s4WYpkP34souVZua2pVVJfbaZ/+zegYBvgfwUO
NnSmuMUDI9wysBj5XqX65+fUAmAVQrAIxk/kBEhncA0LNAz0ngZUH0QoPCd4s7ay
G4HbLPcr+Mo0Rer0trbT2620D91tXFCfzEiOZYV0SyBQulBNCbgJFryNWpmGLhx8
IZqn2oX8voMz4aZV8pT4exQVfC4g4tOKfnXxa30gHJm/x0APbY/uLS93rWom4B8k
3oOvCq2YAUHmdQPnsFFo6Yen1EU0e8ix7+ky1He7PRQHk914DlfXYpPH57Pa3tMu
lrLJbQi0upr8Iz98CrGOMLOKRugx730GNkb0pObEP6QZRzRabrHEQW0118V8TTDf
P/X6CoIwfcWlbt8iIL+Cnb4/NzWiZf7BZA/8A4L7itymKXXFlqYaRTcGvsqcXc0k
P2tfxENotKY/wqKiTI/cQ41G67KP8ZzCbMehnsqvRrFbxLKvYw9jQtQ8JfkEtB50
9epqoLN8b7gc6ZdxB+NSQkBq8PYEi5LNz52E5Dx9BttkeVvMuMFYVhnkbMloVVXT
m5ZKXM/g3i4XA3E2Ri/poFSlqJMYEmZ8LkSFslR6oad8ezKdXLgilqO8vyxzY1sZ
Oop/CFzqAzqD7ujJGxIXw6pztJPTo5xKAs3W/tFVshPc3hTObxNB6vAzrI4vBk3/
WTOIUJ2Pd0uxMCjw0zm8gTKTRD3wLyI5rc8GLDscdTt+r9lIDRSbyhmEPf/kAZYI
eTMJ/ZZfub3D1Xswmrv/TbwmWx+vw9wdh3Q0FT+3tJA/pQwYeMIt31vMOlL9KUqV
NCIB+We9PaRYnfsOKK9SdCtkZaNuKwOZBR/C47JEm7VJnsGV2fZrtjlfVHvlxADo
toSyTvcgEbR63JuzFC3dVtg+aCmPBPPee3BMqnVGaES00mHUPJTqTftEQObCMhU6
oMsWYL7KBQlgPwpvaIOjcKLGNYR/EgT4kzTINUjUFn+9U5+xvQCGthA+AFFwwONI
H3SKaSJmklzY5xnaY12NMulW5k5NJqi9xX3SxaGTJMSh2E7FJWZzlZ3iKqCoY8fn
JMBn7R6WWB5hWQky87s3ydvPOuHLLS7B4JGxxDKOb7ddQKcSXo5DqL+1K/qOUhFx
Jd23kpwlbtqE1lSaeMTgSpzDA5u7QYJRHmp/KNDpPuSVBCctGY+P4+eZNJriRygW
zJyCmEh/ts2qjxQ0dESkuRav0CfwX36IAzl13xIKpClCRpAi5GKSxXM3bWau+5l5
c90ETmMC3tmSBcIFO6beUbBpVR0nyICu2PDsdufByny782nmzrDqsSSn96JHKKya
Krb5uJZqiXmSQw3eZrJyO+df/7KlNkoUE6Gwqn8orKScYfkSGi6ef/I83J0fDwZ1
6gNNBD9yoX3OhY3hDxMfbOXltDqLq+5K86whNOuYZeu4mM5Z3U+OW1AuM+H9JUy/
pq1KbRmRY08Vf8YUiNafQgWSB5HPC0C+pag8r7xC0an1/ThXZG7ut6oBLJVS1RxB
wW7EbaV8xXQSU6icKVgiGwr/9De+butSIqCNvG2qZVPfpsV3KKZyYuibAuwDc18x
4j20VL3/e40qguFwWLwdKsXCHAtqD+sUHFDTMyQGf2RL6jwiwUVjCyODK5pB8AGF
6yzp98jy9psvr9ZjHCDDG8/ccj63RjYmM6buRaf8Scr20iiCXuZ3LA1rOaGsUSnG
R34iDRAOabaxaTgN2PRWAtOBGxDFhmoBOfeHrfAVqLmIWfrhJKapnsfO2Gzyh44F
u2AGt+vKuUL2qjYTM+GDhCIp0u3/7eLs85SKRBSR8XgOmKf78gCY5S2nGXBPX2VF
uppJT9bxjyct60kjj2u13o2+B8aJJ0FOuv7lDV7o8hS0ewvmZYHhgkv1ZdB1oK2x
1I8lboBEfmMBN8FDziHi+BJJcwmwfuVMw+V3QFnfTK4TPqN4JRHke4RsBs0XE3u8
MbPujDe26I4hAm93LUb773Az1kZZc7A+EH4NvYjYyhw4wNYl9Th7BdQ0sRvEvCK0
O4U/BRzwTgAnO4AugTzGniJai98/Hpw2MNNnPMriLb+IWqVvYoUQTER8oO8p8ZSZ
vSiOdgayOUdOKJNjZETS9RO549IJ1PdkB44zlP7vlj2uGHOzN5eOdI291ynOWb/M
LNvHzgShXZX7MjRs68ANmqq40NX/Y6UQj1azZqQ5wZ8i86qzZq/KO9xwcIqRA64G
TA0HA9o5Etmx4yNwS/iAQVCXYINYMzyotWllmKWeNVgk9yrGumVzvlt9akoSfER7
NrCpLRtK9F1d/8jBiP21xsKvPumSzi7VjHUw2cJ2iydkdPECjvxwB9vvrJG4r203
nY9o9bLaUt/cZF/y3AK+upLLWrjxqKpzcoAOAJiIkict7tWsYbyJVGHAE9Nz8T/G
MENwq+DZOFjvx8T+2/jlSF/4bcs8F5aeAjwh4zmJ166mT1ZJz68aGjah8x/1Bpf0
ID+A5Hzh8Lv+rJsk/hMXvgPymSx6sQR5RYwNS3sWet/9QU4yeATWe/fIfEFcb3Am
DgvACu9gv7jm4k3yAawtWwN0eL1PVHPvqrfc4QHAKddQh+OLgDOMRwFOSIkSZBrg
CYrz38my3jXCPYtsigqB9r1IiTQAAizTvsoTkFF/AC9SasZ7hoDKGfGLHL2n4WgI
t1n0qxRVWh8zWuaLHgH392c4RTstb+BweHABbrMQVYDfHQPkGw425aIWeS9NC3r/
ba9w6daKZ9O4oTi6UtENj51s/NjoHcHDrEZCWlpusvFshQcSFMkQfQPY2oI9HgdO
0b09S6Gt/79veykBd33cZhdiM8A2jvP7TeAxcV9y6fljdQXHSHPPGu7XNHCg6AaJ
F7lvFK79gIIdbo7qcnkk7lbGE/9scEBNDPPKprsW+LcdG9Dk0kLumn5AoC+nN6j7
WgSZOR3kPYStw3r5Bw4AtEwjeACnqizWYlfcUsnErCS0sEZP87GymCKQeapbZvAA
T5JoQhIowNVCUW89JdkSo264XUbGksT84pefloqHqv1+j3XsgzRohwwb+qWB2crn
LZ+QPIcVCS4mhO3ZMa5wACdTf8mV+N6/v1j/qQgGF5ZdqfuZ6/u4j8KqGqYUda8V
AuWwV/qfHRb4mrR+oN9Ei0t2JFnWsNJN2jaaa1Unp4r9lZUO+3bh4nAsWuQe9v0K
aY2d+sLzGE5v49LJf4di4xfSI4vicpWXECHAcjMhUO+pGqDE3pvX0/zV2bQVK2vC
XqKC8kYsoIJbpCh7bi5F8CciZj9X/68eGrUTE9S35Do/bfO+XfvgNfEGqNNqopCM
01u7y5PD18rbh+rrOaF5uyOGo451SVHURABVAOp2PsJbdYiN1RT5r/VmRcQhDKe2
2p8SKh92MUWiZMTLj5sG9IuhmTQYYXmuXH1agJ+Es6FNFVD66HEu5kCckBviiQne
B+H/dGqLVILTNgtUMCJ3NcLj8F/W7nmnR7F1rXeQ8y+hDyCmDiGJAd+JJqiINW0A
cv0yaPVGWkF1YDdneJa4bX0PZDpvta7kF3WaHzuBc6HFoWF1K8l4hNZVYpS+JROI
diai5AthsSHvU5PQQhDbZhaLSurGxtlMmwVx04gf8Vm7EL1Ks9x8VcvaSMDITzNO
Q3sS1MP1QwTvW9LJUn25JbYFzhSg8kQTw/JzEqst3zEcxUxDBdxlcdht7/110hqS
/tptvFhSXvqCiglzZ3mq49HontrQSUNRveJtwZtK14Ri5fb1jfPT6d4DeHyzdLa/
H6l1PtYXCGMUSG/d6C9kTJwMbqRb5fPH/fR8kcosBIUDZc1C1/j22k1wEoN52sJ6
s6gsKpcieRzPFJ2Y2PEUJ+5iWx8ZpBNZWG4RxzuQ3RBw7mhDF4E010Dzee1jGyW2
zhze44Hw5dubLjiFUNaDi6EGZIbhEXbCxUwh0urgeMQVtHijjoQb9k7TE6C9IX82
X42BSorXR9o9MZ0t2VB5TcmsQjzl6zaaX8CyRuq9CkEhfWWLNenq/BUu7SKJhJtx
H2BSwoJpjRTSekhYIavGiLM7AmXhsvLnGwFwoFzBM/MQ4IZdapjR28UoGdgaSoaG
c3xo3NkE9EWTp0dqjo/LqL+niKCUKtszOBq8S+/8qEHbF8pcQzGPfWEgitpBjRZr
fJpcr9St/3OTjE20P1wpJoQQBh8Fz3E5URKUodlBbkPYOZuJbsgN6wuy/xVsBKjH
jFy4KMeo1lZhAAszAsd93V+qdIpjzriSQw5hWwNks0GO1t74N2u4MXM6vrXeP8bd
vZ3LNqxqckUtcrIORndRI8z3hzihgr+2Y0lFUxppz8zno/iLQwM0oFHUesgTgmw2
fLxfHEq7HPY5a9MOcYtQ9bb+aJAmZorerBw2UtyNdSaGP/r4usJZtDP5/41PmytG
a/ST7hZRGr3S8+FKjCXpjP200KsLt6zjcO9LzfbFeNlylFDO6bIZBfNJdOx2iwKQ
eYVBb4eA3s7gJT2UgTJKbB/0A9anvWdgM3ZE31cX4JUZtOU6G5RmB1h55PmcmQPd
Tc8ogeAY230M4lWS5rgvXFjaqDm2XbvAdpOkgPuitsDY+mKJc2tTArSI8Jm0pX+C
phbvSWLfSrjdCA7Nor9qJll4joGTi5DS1lEbV0k1mS2xJCY7mJ5H3woVKDXYySbG
rCVEoVjgjb1T91RsMxrLHvioO6DoFM9WU5GIrF37VD1qGv/P1+9ZLdF7fP+32ica
XvhAQgX8En43rFmsPRF0SgQaIATKtAFM+9WVg6lAtIzmGyGgJ18EpodCLN9itJE/
wsXnVtLm5M5dnEUBHPFY7AsF/7jJsgc5K/8oKzHxf9ltwADr3KnqUE6+/hly6ufB
0CKFDamU5OL5tYSMV6adSrk/KxPNoLRcxqJjwA0iN1mARAscwZ1f/g3SWNmm+8dJ
xGNxWP6NCfwmLApuVR33PQh0Vd96LldhqWfzwRoIPMHGP8z59HfJfyLtdoLqvsn9
48XNO3iv7s3FjP6kcGQjHKNkE7Iv9zBH2GtezGipMZdtTAhCdSiiVS6JYSW9swFg
pQoFHYUEq85SETA6RZr9aYPMzHadfG3g8BHtIW1vPIga1o7b/TlXreRt3EZkkkuH
iCLvWPjh5pWnlbVn/0Xb84dfk9nteQUEhTPk1nzvxhdk4BPg7IWW0mekCBowS19J
B9mGKHf1nvhYPLL9jIb88L2DWRXFwSiVuQNAe1uB4zvsYucQ6Ahk9CzSL2YMVoPQ
0nRENoGlaufpx1tLk3exrH6f0muh6uHX6fhev1SJXoux0N8iilP00AtmeJiekb2J
X8Hdg9V/hp8AN3ifEVnO9rTbU4n0YXY3QyFOf1H1yjspFdYFigGge2u3Hb6R63G5
XayMkTWNFWB69yJWaMxiXCtpJqBvh+LcAww9I0k/I7cbPEnMasVhIcnbJ8hqYQsx
+VdrKI8vqtEskg83JaFdGNT6hf0KPsWU8HSFttxGW8SCul5eCuvUM1m5R4011PBe
2LwbIKILxrqdJOgzKhrSGutSiZG4UcGwuSp+aRUeO2n6cY4wT4qk0uFZqamMPF8B
AL+bvHQIdD9yt3ns8+r1Qd969yFBc3iYFGD1MznO0y8soCZlsJXbMn77IESRA+Ln
gok+0v5xxVtglNFt4+8Zo2Vz3fxhbP/JSIHMNpmGwHcUSlbiI3YFwgzF20UFleBh
Zm843jeTDQfHrRxRTT+qs4tXuaPtyGC/ceUB1IV77z3XJQeCMK2VdcQI4XFa+XPl
VdagJxYE7eykUKYiMS3LOH62ZKOCPdjljBVsLpwPimdT8zAoLs5kNLSjxXhohQFo
rn86w1lO9Y1zfKcg3lA2ireWxdhBnky/tfRsvQv4Y41d8UZDoBrhOHMVzN88ssf9
6kuv0BEkBbuhyxz8ARiJ4e43MefJUk2oqzZVGPrIaJn33byClDAa+xjrUvUO2tJN
ZNfpWCruP3R+NE/RRwM8ZK9VwWZnCtqGyL4y9oLjCWTQpn+/8rm5JFH9Bi0VzssA
cf0jR+T79AIkHVqVLTtseh6i2dwW6eJokhgKfIF94tdMvDzcdE3apg9CUUvw8afi
3DCCtBofqTdGd3q9N8QwSM7zsLjGnzVed904XMpx/KNzOoWj6K9yZloG62LhMFC3
XenR6i3IGpKaBhgWRT4DAJ632xbYPIruV6t9NRtZ8FdvSEy/AQ+3HgjOcCv8d/+N
OSltXvTojcmAJleu5tAKwjRgOTVsd84UPLUX8IGXD7pFlkPmZKTpIBOzA9pmhIuI
3YcAvZiwkVsPDgolKPCCvymHv2mko7Q0psZeOu1Ec4tEtuggIMG/GKXEOTvce9Cc
m0O4sVyX3kNJhkv0aUkwI2wKk3iyRfHEy/03sDzxeKcN7xmI9wMhDwTsxu6+tHbt
tziGpEloTd+2vJkZdak1gJAgB3sqHto5vfIH0FAjNvcQDVitsyMmHN5trnjnKlTy
q5suAalGLK8X4iX8Bhwbgl59WuMOtiao8ONOQ3qtEYcTJmtIfUH3aosDll0ayAHk
1KhCu8JGbMCbl6xcHpmZuMIQsmMjviR6z0qDdKSoiuZCvCWIZkNwdZcMvUPSw64y
ati7aum+mZuopPF5A513Dr1qGsULkiHm4yfHzrNhtxi1Qgq+/oiOFaSq3nOO881J
uEEZ3oFs5KmLmu9GUrLm2o7+HHG8YVwdYgjN7+VVkB1vrL/TM9pWeLDDdJwFSwPY
JiA+RE+q6fbLhL52asFD0Dz2X3h1vux7iw8Oe1ObwEF1Gm7WjaItvzDqC36caffe
3062FvQYsgFo/5Z1LUyZQKwFBW/jGs3nu+3f+RIBmuNCpUF7ZfZ8M5BqPmuROaeM
zZzDVoUfBltwbXYZUEwyq+y1b2WgVqEX7Vn9yE+55ES5steN13LkhxavVXuOsMoC
8wHu1looW6OvQIDcbrCcPza8leleW4h4yTKirWKB1yn1jybr1mWQ8amuCpNCZGe+
pkNbQsrYkev4cV04tW0Iyvml6CSJMGDtKAt47U0OiWpe4ZuQdMkiDcZ+nO23174I
DSFrVYeiKQ39x6SCZ0CTQLJ1zkCprbfABo4FgFCE0Y4RZVthbJPnsnl9RA+BfnV2
zAILuguf3oS81gWaDxSjJp+G69lK8k8Kq2ViCc9rbkpjvAzNoXmIc6xHZ58jtF6r
DYHxMvw+G0shURXd3sE/g6fyu7gW84bllgigK8egtOfwQpy9e+QX5cdSLZTwcHYN
5wLTUxsQN+FgUZjTZqtfBZKY5CVkLYKE7LwP+7ybnWuxiNUZkSae8dWMHyjKElJ/
Mel/zD6hnpwFPabbBr1uflcUqWD3MwGvLVz591a1mizbyt+WPoX1QsKHPEXRQRtV
9Zv1g/nwVXW1aXVXUr5fDiosooZsVWlB0Zv7qpxSdj+GzHMJ5SCU0FClyt/Ah04o
hxsMDlCqc8mQWQByEhhKl6Bp1lPTJQQ706o36EvTqguoLgmwgVbzxJnAEbuv1dI+
y9dxiYKdkUv4U3G6AMcabzMcgGthSO3JTSIf9sSMjx6Fmqll4Ko/IbSZ2ffdPBD/
wZAXfsz31iWoV5vj7hT+A9xHU/6heIa3CBCdPpYQ5srKT9mBvbCI69yzyZmAyhSB
EQJwZ+K67UiK2Gt/2SMsNyZ0sVdAo4k2RI+imJ7k1/A7a8qH60XimUr3MNOiSWNc
NJLQweUxuKTTI6tuoWogr3LgZrgjnkTCCE1w/dOYKZgpaifZxdGGb2DOjVuiD1Uh
DkUWl5xLiHB8OOg7lJFCh8zL8muxQWocDpK9kgwOEo6PcDkLO4T2E2frlEAGxTZL
UIOx7naTJdOmPb9bjG0OqGLiZoHZNGL+Em9X67M546/mdlHr1niFyaF1oFrsiq8V
1KkyyRlIPlNEBWPp3ydHw00cG/qfP+jRO1TsiKVj6TvSUkoleZqIUvgakgKpb+sA
GJFIBBDrkW8D+zuZaQRxzAf1G433bgdxzEuZOi6KRUhseH8d2rZY0mAXD1tlyb/2
DmYZdwIHKA99uvqHu6buclLtdx04wsFdrgfHqe/DJKwpCx/MZrdveOdzTbLncTyL
IAlkMmEGqFrPcI34OMFF22DUEyHv8Vctae8+pzANNh+l57rcnCWS9PjIVpzztb7t
5hsPK6GrgcWtV56pWaElDFECFchQxQ7mwSrEPkiakCUgOsitfrrKQ40T/9LX73x/
yN6aLWKZ7EY5CjmQUsEZmJ8uHRzAg08sPO9wpOXabOpLu6yMABx49RjiQnLSB71V
Z+2l4KMGJvIBEmT+5RuTPYYYuR8t3rblOQe9vmLFFZ3L40R+M/aDzg44jbyM1kJR
AF8tVe3HAMfa7BZqlfDM4k9fmjr0BiuG1JSgGEjOtXhtV1nYti3/Z4l4jMbSvOOS
Srf3Gir42bRAMv1HTGcnGFh+v2S1vOhhaB4oNRhy9ggGDl/jTeJ6+yCftjtExMu1
RqdKy2qM9DXIs4ljlr5kV4sfRVyzANuz29RL70VGlmt+1/6fS7oaBlWeuPsrvZBi
dLyoEldnRBs9og28DuH97IuicY5C9qGb5T3LlIJreLlfQC73BFt6ezczCxQfvO5P
Wie6rfi0pmthjdgaj8hN6AIJiyZtPTsfsslVn1VIPPAKlReMzLmg+7dpAjvpeR2L
n8nEFzugcQQxn59SUifYS4u9sgvNslpTTW2/J5UzhrhF8em96rQrymOnzCJV/Uj6
/pVkD5xE2rExnB38Va+UD0QDAGC8zl8sYSRANdELYowrj+/Xyx5HtWJ05MdBRwoA
Btq6e6OAvJaEtqlQQvgpw3D6jc7h/btZnwbTdQn9ZCrLbsVm4Zb5IZm2kLqgvq/j
Bw27aiQOvyQ5K7C18SrrpSTamY2TCznSOPm81zhLSbviq1JCBVRprBK1mEdV/N86
LE6s+EX73dkBVm8KQbHbA8+weVwkaMHc4dbI4eEPiItRqn9jKPZM+Ei3rlfp2GEo
gxVu2FYEu9iB3u3CamQnX6lkzrT6plxC9gk2mUd3rYvuCD+jfnwdsh6hrEYr5CwS
9ArynnGouD1N2iCkDBGUG7KdwvA2K/f7NYfiEVgRJTZz9+au3bYIeGNevWCSCgu+
hFbT/ySxuirkB9tiQcizl50GCsil5J62BNjlYgeWMSQiywecu4lf98KBMXsoHpzs
2OJNsDesuHS9D7dNA5jrxk4utKCg8EP/Bv6tTPv6J5HY+2+tWeXVg2dZKt3Zc6Xf
/ysqVj0dTmxDAPiuVIkI16XQgKgV/FoSvnUSN7KsgxmnmsR2C6E+slnnABeWI5iP
1LUqrQITzxBwQtM01SKuoP7WdXX63stGWphN+GPLmpzDd0gG88IuAHmZ0iD0VhTM
kQCcaF3NvuR2hSI52xz9if/tKu/9/YJ3j4V8KWJ9JSMcYunfH5rX0Cx6sZWs1pe8
yHCQ+dQCFwes1gaqPMHwQBVQ3cA3fuZga3QW+7mCOEgvYSv7ssHeAZYtc6GSUqGW
NouAZaokPssAObo4dredL0xYQvTzWD+Y6r3mpcBnKl8pjM5BkFqk7Jmn5zAAMB4t
6bisT8I/OoP3vq870/Lg2nQ3nD3Dr5q1cF84kI9Oh7MmXJUkE3XzoIvyj/ojuZhc
Uapc9+hNCIDxrDtiODcZBKGi+5SE4GThxABjtewcznNPnooDuEtiE/5BHB0Qv+a3
N2Bo/jdXxtkD2tFZeGePkEyCB+43qoW3yQc06Kc6zrExuhct4fsUjf8XG8cXlJsN
8Fzphc7YGGQ2ggjkSAB3oRCIukI/h3+BoYKWLBaNXRl5vVMhjUVoWJLwgpXgQ7Xr
fDctGPRnr6fPYwCajXdGzD147pY5B4e1CeSM0L1DFuTj5Qb97GHw9dEeLZNE9+TL
02EoZRAMv7W5VLdpuhFeEP2t8wA92C4Cv8uueTG3V/XrixE82TyimdBIOmXNmTC9
p2gL1Ga301LOseRGYm+UVkJeXkK4SueHW8CdGJZvT3x7u14pxSoz8cJOzX0wch4m
yOqeZ7YpVScVEp3dUIIFrZucbz3UBxtP2MzAVdcb2XNLrp1JGDFLnLFSJQNgUjXZ
uARfyXVsk3/5D3jw1mEYTK8dRNhqj627N7K9zR3JYxzn12Ka/39WU5FqX0iWryDX
FzCEXC9vrFJLeIfRKwXYpv8OUJ9XqiWW+PDNcwDKPLtKfwizYgSuhBpwMDJngb6D
HsIgNrR7oTgfsbXC7CWJtTJ2a475CaXslTgrjXMuswxg2wwYXD4NGgjDrstCSfBf
75vaA7llUmbk5qZjet2fMmQeAWmNOwSt8nWkYPWiHr4NtgG7wkA+igE0fX35n0vc
ctcJMhhJTuS7CSqsPdE1HP7+q/Ue8ZkuwkQ3ud6kyb1ir8QZuypau04jeE2ewfzg
+sN0PX4prwBN9dxP8MpEhczcoejMcnjWgkmqejcJ/5EU9Ow3tYfisHkkkCalvF/Z
D5HGSrBAa7nAt1QQTY7wH2SCCKszGCGZ6/jgJRxBX3wB1cOgQ6vbhKio8z5T1hMD
j3S772pFKeUE/PFuPFiWv2BkJPrf+mlnPUezK+DEcITj3n25SaY2nYPLGES4fXLg
iit0L/XNIcNKcGfr3KPT83uaV0AG+RbocL2v7qnJBWXjankOPm6QgKDkxs1w/L2y
VMC+y/Th8l8wYrRYmGuPQo7YXrDdUbHLnE+tErGCpoFTXviBAsZ7+MYGzV4C/+ti
l3CkYsMxsrXONhMc2cDxiriiXTRbL6Q05BNHDV03wqs7jAAmEJ4im2ASMWVbBz4F
Oq61xBhhYbDLxhb9uwxWX9CdQpt1nsCj1aVoXmfpyB+66I5MHn6SOTUEos8edoIR
xOoBkeEYg0BqUCSya6/Xcy1D82dypPbgrUl6NnY1NJ4faHzs+EfIuJttqabAxJs5
m/C9FvaXVKQZ6WDixcuCAxwPVikrDcT1Aqga4XfqJ55b9zbfzCq64ExXQqedSQe+
mfnQz5aC0hGxXqCa6EnV6JUQcO+Il0sCaRwj4PxIRQRZR8Q0CCR2ASnHQ49ey9R0
MIoIiCDwbhwLX6dK8o2XC96u5CDt65nb+wiKC35uYCCg4W02YQipcxYGmolnOiQw
YL6Lxso9oYV9UGCf3FiYMA1Irahr7Oe6fkMWuJni958zgXfECFpJHuHaLC3pbf09
4fXnPZV6kPJin99inpDzA9O4fsOEFvpSE2UQZRpUPRv9YEcoLZzQVtfjsBL88DY5
Q6dOVBqvbys5oUvd72yGGXhpBO229aM1sXHdFprsjyMqakpHHhUmRg/90sH6hPq1
4nHlV5CPX3mZYG+n5CGIlWXjJ8b38PVNIqNjpFMyKOxbbf/+Wog770HLNtqq6/Z8
3N7k6tvvlboB5GspyaMzjJG00UtY0fVKyshshaK+9+3Px7508JDjsdhDBmSmQt9V
lmbrkwpjUTopj3nOKo5XzWRVlwphfzaqypKc61zYh6iK3mbFa5kUrx6aNscn38iJ
CNhq9TPWxs8QnzlKWttJHV5X8PaYxwOnToyjFeb0Ao/O/D12QendH/AMd1BRz/Bf
vzcnIT2Bw90njUnRWZ+bVtre6323CRItJcgADCLBK0da4Rrot4Pju2NzkkCUSjrF
WotR03KvUsRNgjgUaqfs4Oj9yW+3+idKQp+vaO66UaTbjDEZmzmufHSw4KbXLNxS
4pXmU4STKDVcFF6VlFRXi1HBTeMEWX8bjaROv123Ri2LFO3bU3j2/dz7Mbs5Oukd
d6Z4qFZAt1m7yWEpczXsXmREANSdyUw/txCvlSVBlpUzSTHvk8e6Imk5PntQJ2pL
ZqvyqteLe5IcSXNoi9eaCaMv+5qZb/UFOcX4igDq8Wr5zkFsPyJeQjOSSHkvDJYL
T1i+G1K/AlPSXPabsle9AsWBvImqvACCb58M/m219vQ9TftycTil3umy5Um1x/7e
2RIcqnICoIVQwNuFRPkkY92ZDSKdYHQQwPoV8ABCNqdd2A0rFmkojMuNO8Zv4KqB
qkgO2++f7Kzj4uTwcU3Ki86ph1PzmsRiiujVXfkbr4+EsDZMxqASfntsqpQ9LjUY
X8aeHaR7v1tC24StQ3WiwSOz9+cqIVWGh9PwNLaI3GY6gVnWQJvOdF1sfX5E5IAg
E+BdUTStwoQMG6y6SbVGvHpVPMa/I+/vyvFf9o8dTM5pVYYhsJJqWKDfBloyD7U0
wWH8S00/spfG8IYd6Q5heHFymuGt4duXTRVIfBNaASPYsmbxUXv/7MHi38shEKf3
MEZ+U9w6D3HCX6U/aIoXWPifGyvWXlXU+abZwHlAru1vZa7ZS3qpHWAIzX3XNLfS
kvxiFHgX/Jm2AP6e0O6LKiOQ+9XegtUToSzLGphY3QUgn+FrVWRijo6Fg4O9B7be
pJMndqCSowvSQSn4zjR43uDyIFh2enxrPO9AB/WMurgxvPCVOU15kJEcSr8zJ6QG
pvV7osOMFgwc6l3yqLfpMrSHAM3P5YtilX1BbLHnP4LsCcnQPQlKIszq3XxEc3fx
P1R1fxPfKuDksQQCwg6iNa7v5OoHiW41GB04W+i/MRm41VWWcKArajoZd7X2otfY
9gY+tGq7yo444EvWfDpZSY0NzXtgGukrhNH0ACeLcrNzg64UHrCLUy9v2nofwj9G
W7w1cHJQ9Vi1XxxdHZ/c8ynHATUYxpHiPErsTphh4G4QHvgj6/zdTzBcuUbdmQ9d
F2aPXzLo2TG0T1grL7u5Epnd3GH5fYv1CNOTWqz7Dx1l8bKDd5/PXjp5Zl8KEJFV
wboa+A1pXxEVMZIGHU3toUalDWmUkvyz8Q2X/P8EAOV+cQiBysP22mQ9wblwYYTs
US0efcDClUEA7ivjMdFDbA2H5bE6+wmR8/1hnCprFJ0UVtLTYqvQqwxaSOPywK9w
zqvcNyFjsWiZg/6aYnnfmyNJTz7cMGTeecAONay7IpVGWUJ4iHCWl3qhFHu3XE2W
MQ9Wf458SPI3SpBpm7iRpiNbmJhAAVs44fFmpsOWIRtXIWcZc6R4bUij0tn8wEYh
4fxTsL7y+iDjuUJjW7i8xWLidIEkeKTx7nmbWQiAiPiK8IOigij3XXNzNTWYa43+
8Mjflw6iYLjgtHqRAkXQBtjkLqhrmfrV6Iv83jhGNBoXHZE6AJDCwSZGszCQ+mxG
LtU5QtMosPlFkHdU6rXDupEOAIYYLBUuRHiczUNMxlC8sifpNZCGtLt+eeizIdKj
ZBsQQPg12TdMIEKU4CFEGFIlg+HGS9Eo2xkhpOtvheSoAJ1NbGRuUOrPvdX+9Q0Y
5J4p39OXoqTT45AeoRC9J4lefx4eek/Z8kFeWCAkrIADg1eH67qMPDjmQkj0j3qa
6gWr6PM3WaD5DLZFN728M4g7JLmPoq11baIXWnsDStXoQB4QmJWRMJBXpVBDcLQ3
+o5MfETBlxjfHLtzfo/jyCr1xmNUIYzWb9SKADcqau/POMVjR5lKkWsh8Jrq5z9e
2ynF9kUihfAx4RJ/NTuQJmFPiuCmCRjogfVjkISn6F478QEEei2+UvmPsVLrk4wa
/nQP1JVt17K0ha8L728kxbLSmSFYLJURhKuY/da3y+ft+4VO/oBwkC79dAZAt0XH
1cd8Un3myE1XXM0SaqQHHp6g2olYcjXKoJKQsoTsTo1Jo8AiVPbTxadmLcHutmiG
NG9H2GlhNMc5xeKc6epfLROBwb4XoFpNl+yq9rIJgSEvjcAQe1Z1oocB+zOq8p+E
iAi4+4j2Bx0PhwJgeKLlbaw8/tgJK3zOpOqDN9Zx2pbNhmUw94GJ9WpgnnHJK1ae
Wj9UTJCylU22+abfo1zSd+tWNF6wzHyRhfBRW2lic/tS9vzup2g+383TVtX/C9ut
UkKLfWFzornn8EbskuWRMM3pCoxGp39ryQlsSzLwwdseNpd7e5ctGuNYh1odzgAP
PyKV4rw6ogB0iwCy9mWRU3yuJKLB0jfPNdnGX2LAp/sW5jT2ryXCNkHTvcJ3Tme6
u3l8GDPZZ9/UJgV6+vJDTPhly9gmRP+rqb8GUSeoR2SGarEVZ/RLXGDp7Ct9WpHs
CW0Wu53RmcsO43jkGdz787mIUCcILNJ2vqVVmigVH0TTSwglbkeSPV0lnL/Ql8Nl
Oivo9cap/sQAOAHKiRdHmKg/wNZp0c3p+2Eri4IJbRWidtwMnqpsBgxjcz8k4wlp
uf0Xc0KXMluY/wDbvwJiRY53ihrBayhIZODA6DsUeJp0KX6PMx40uL/dBYsf9Jo9
Bez87NEp0e2noWRuhacLbW9tg0+5PUhiMXLgpRUZofJ/srK3TW6YSSxVXm4rxcqK
4lwj1qyCVd203G1N+B0YHS8luUeCPQ6yaL3OTxx10lmDNwy3Da3f4FgzoZjpdnco
d7S9TPo1jj6TOwrzovCtlwFeTbcGW2BT1Mrb/V2XbLGbXkI4WsezMNIXxuT7RZpW
SAdGCI3BrPOr1V8kpHdrf0fVS2dScmETFn611sYZkbrp+PAGXq6dantn/EHaNaGM
wp+L2gj7GY6Vx6xGtw9MpWZ9PXkWw0bjiII4AIFdlow11eSzABAsA1nXU/NHmN9k
rQHtyCZanKNydvzSCw5OBp8KUiBw44fSFemON4g7GUOS0IQcXQaPx/A/PGmTTkKA
uFQvxiV+ZxocMGk/DCL6OVLqbwq+FCOCd0HCoGRdpyBGO/NuMxRWUqx43zVTe0Xb
fkiGczC0Oj3qNGlUK1sAtQC+uboxd+wwQLmUI3j33TQPW+4ZurtMO12R1wIQgJvH
VsVUpl2des27JU0oxWEpvHDDraw8AybeoZmqL2FZLt/m3OS3t5UKtL2VLyJwYxuL
uml4Feszh2sZtpybv3EqgvauDqw/Zyi0UoTzqsDyUyLcyULZrU1goWhSz8+uvatC
47B2fcHymuDd0nBkJJ3GzDAn3UrzzjK+P8CnFWgdnuKxqIro3LV9m1VTmTiPOZR+
pYOCG3YsKPiankKXM2Jn2maSUnhW1vEgU6nEHzcfma3GgG1pQJlDc/IGwMj3xU7C
wxQc1Z7DadzkhLPEoTO3FO5XGG9EFHk9+VtBl7RUkpLo1XqJMoAQwW1CYhRBq9eN
O5xbdP2HVSCkZvwz3GleQn45L7aNdllxcOQrc26TpIan5L5avmKqIGGcwSTfG1SV
Ks3zINgCwGOBFADEMnbvthVybqX9ZrmkNbcpOzDIjihHlgNYDQyBUCM5Zze9r3VI
JR+/e0FC4ZOvGLIdhhGiQULZbqmN6DxdOtVaCrx6ABgwHqI3Njvwb1d/d6H3CK6M
YXMfoOvg46wQ8IRyvTQTAGVyAYMX8mpJ/5CxgENyLvqeq5eU0O3hW4bW1LyimWEW
CYuke84oGApisYclIuX7PjcDkNUnbOkpzl/MELq2rPoJEkkkDNbqya6/vy7lL9QM
qVwEFABRrcIiC9Zq+hf24NgIFhfJM4Wh0JMVvSfu0iq3X/Ivm8nkY+GMmoHd2gmI
T3YWjfQMPT/arB+jDW+y8IUl0H/biFp6t1brLqAS7+yD0hDSSXrp1HK+cSnhPNym
Zj7Ql8Tr4jeQPiMtjTKTKDOMX7ZOY8xrqHFFRvmTUP6hYQcKBmjcy0pZ/LXILbQS
aGpEXFdulvEjS48tRVpBzf640UGTc/mTjKQpmXvgsHb5JYj7D8E5bI01T2lLAtQO
eA3N/NbMsWoa8lNjqblIRr03QR3ug2TyT9lTUJVqa1n/WF+3MY6V19v+Ehy+WSYk
lB+xwIBX7ZpjyLUirU+4S0cN8mvtAhq2f2CInxlGzsy9t1kUYHe+taJD2e0Dfj+o
tKkwoacP+2HVTVsRr+HbwQr5liAyWtXKpDMznqNZcSAHP4+43bivsZW2yPTEVJa+
8/5LGBXpqPl/AaOcZ6FYVYU/lm/JSu48iAv775k73CzXSjQ5pTttBIf9HE6Tpa2q
s+F7SQS9U5YFPut3TH7MATAJcZYutXEXM0pggseOlScTYnaOChkddewbD/oxmvE9
32FEmrLN9VjmcHc/4IiisaZWF6FVNOXVICfSpcjYSGs+QKNa0xZCYo8zr4MsyU6S
7oMZuPrjS6ieYWG+rYlsnwhWsWpPBXWL5/RhbW1eKxSeEHn5QbA+qSqlSffaiS6u
NMa/QHFv+L884iNycFpWn27MXFzzT0mm+pu+NbEK7TDoJhAf2Ot2x0sa04eVPjZ+
npv+yIiKDJMCndpYQIkgcZhWHWVvzV64ibAXHogvzaTtiTe4Zh/dzmcu6dewYx3Z
NsS7zqNso+c+eiPl1jEMOf3XS+RpnOHfaJpnarSY8Hnb9g8sTjxw1feheZMLFadE
VJ/25oPk3JIFlRItPomEbM4un5/8hS2ESiIlvATwKk6fXnOAUnw+06Da/KMA3Y8u
WzOD0baaEe7TE07n+qHXrM9PzBKEni6NShxse7E35X9gVZ5rmrJC7Nak7HS3qtl0
JqNVvoSX5mRaFu0/CAq6K76b+znY/0Td6N1493s1bUM9vg0etBc5AngEioiALAoZ
ii4eETdW9TozzH06BpCTGb9aDS5+9AyA4JsEyyYR3jv/y3YvI1KpSk7viI7ipk9q
E8Cs9aEpbsowg2TVLbE6lcaouPdhELdTja3aNCeh1OGPPry2+KqXnu0nzI0UPh9T
arD5brvVZX7K2CiSyYCBxgjzKMafBml0XrLSpqfjChVsBKtuSB0R/6FdamPje2ud
kMT9QClDFh1rKAITwhbTgVpq8Jwzmq+ZVkWu1cHe8SBx0DlUJVF8aw/ln7FtX5ZY
Ij6+xFlIfEdU3wv2/4Y2/+l1tD+gIJQCnwF2iizPyKnBdFX+A4+VBCEsNBM9RF9D
V1Fv/mrfwmmn7hlNJgBcCp1uCaineIvDcKwn+FcxQPt/8oPdbMiVDMczKPWNpYj9
bhIMS9ys6H5el5fRb3YzhPVtXvfo+gvKf7eTlHTOmsJIVyFRUmBouOTIj+44xu2p
ve8cu7W8+Qa4yOn7rURf2XOmW/rWVnkoYFLbKF2hhsbz8WQN18CqcW8IuZOMoAop
p0+sQEhylA4im/woH+zMSA6aXrSAmjDEzHRF1kNJz0AwDEXxPeT5DiACkXjiRWwU
w4AXj13Ap0Mos/L6CuNNWmbuCIUMBze0lwaHWwCaD4D47YxKdnzuZ99crm2fzDUQ
F7hdJePIAbuq7TEMMnqUDg/cNi2vD3s8KXIiu8lOq77HMt+XYoBH2jnpXt9hXel+
lv5eES0B5KAkTrLmtgagKo6BRsTPRwHowY2xnjjoCZ1Gm/22fBuw4/woiluC0WWS
NgNE6svWg5h0QSjhzkrzaMolnh/R0na32oc+VjVZ/Dg1wxXDrE3zMiJo2n18K69M
ssowTEp6/mI9lw02k2IhstDJ+n4P8ukzok8EQu0eA94r5xnQbyTYrYi02swiuV3R
zxEQ7ur5T+nhqgMoLPm5PZ9CgLV+cOsD07owYLJanqNcpn2L6NANHJbm2zuDon8y
Lleu3zMprxzZ8RwR0B3+fuR6sWAqWeyXYRUNszjCU+WD5KRDOgalR7d3Fz0QDQ/D
jbXRsQrlkybqH1gPz9MttpH7bdr71ARdF2PYz/XDuiuVBC+Ek2q9vIy0ZsJowRH4
9k7FFobDXNIz+xHk5f3QYxo5Hw2hw6FWon02+XomyFUKFwXhdX7GBd9aYKC6PjPY
I3XKtTFwOLo1OkZb6mI1CRPMTRz6UO7F6WcZSj3L3kiOpfdeMKXeYyd23qlrUk+z
7l6FAwwK3IMJ2Bsz2KPMmB2/Ieg5c+tam6cewrEcVQAshQRWNAWWV3FJrIo3vv4x
z4CoChYtyAuYArP8eSoCZt2jJD8QeUlWyPqVPnVszKsA9NIKE2yj7ZnXkzAopQrN
UqjkuNVu5O3l71WqseOX4XNtScOhZojvtPC1JZPvSWZN0cYZUXDzK1QFQdG6oskk
9Uv+2+UAfD+AFpL9pn0cn77/E/3kkx2f778B/YA81WN2b469Tud2hw1KjiXAF/Hr
9mg6vrSh9hzdBQI/LNcFPT/elR1CZCTIV+RnOMoU5TswSf7H59eSzKVPqtwEAGEk
/9hHPLq8lHTyV2H5aUTnFY6Duycrkc0tTgbxm7uQlZbWi9Sj7cbc2ONw/y1gc3tg
oo64PuVuC45DTbempJumFh2VodGhkC59OrXmSrwe79o9+HnndIqCiRUBHBA71Bn2
hKsLdw8rNWcguG1TdS9fSlNSbZtENa+FzGoC4cKzob+a89/0LQNGNNlaltm/k/O6
zHZ0bkxL3yX3+oqrCGxZy6z6lT79vv+PcyYlGijLE9gypZp4XYy36ahBJ1qdHBdl
iW8n37UmgQ3PkvR6n5We8mNu1O4+89CSywamA5mEDk9goQ+hf5YGIaLoctZKxNYG
nmpWnnFgtTW9niYXXqoPFtLF0bJ9nv7JG3awIGrcSPyuT3Y1qrJ/jZvEsbBDmpIu
KlwV6Y6g2Dso9jgwet7VoF5tWIkR3ninI2vZQvaQzNrSv+xeRGILFnENbhRBfWPT
v1abmC3VsEi8MVKb/h/wKDAgTBZN6nV1Pga5VYSLcqtnx57AVOYeb19M77WSgRE/
AutAmUV0YPudQoCXCsK87NWEJtiSW7rAiREDa8atuBVWPb6zeCa2Tg9Zn6Wev1Ii
eZeov/vOxqW4ou4qLkauWaqSPwmIDq950vtIc0CAUCUC0aLYMwEAQyeTAI0DSRwA
POjCetEtW2fDUCzQDzkqSy9ZoH3olxLpAHD6LS33zPQVpkPHJVnkDT7QLtE2jFXb
MXeoSuqcREJTUq5dy96dPblz8D5JaJJyESxw10oPV1uNIeVJNW03I0pWYkvmi4J+
irzTdk8HFTNwQDvpbxJ7GBI7F/K0AxlmkOJmlqydQJlpiettsCxWZvx1BPHO1LEZ
IJfsLoJ0MSbCegFL/cSffkcjlN0VeE6s8y1quVuOOZDXyt+rdTAP/VYQIFcIwlxY
ibL5MqOxaVHl3OPaCKPhFznSYWtlZ/EExjdrXTTZap8BnsLviCiPGFKKzym+y8+P
pVhI7tMmtFHRje/XqVcICTNr5ojv5vz6G4uWd0Z2hx8h1VPYwnInCo+XcgkfwWCC
cbIi702RJME4XsxFoav1480pzF2sctLDjvHast4p7T+Tolf+3PT9sodHP0Uhfp+b
HWtGKiNWTQM0d0PUErbbRTqwOGSc6wDcPoYh7LntND82e9srHm/jvyIRvF+9XERA
rbUw6LinXHAZ3h6SRjxwtU57QAPx/KcnD0+zkkT7DdYxU1p+YEu0lisQJzKKjrhB
IIQ5GmZGJRxcH8WrrQQtid9V786mVJkODPNGGQKbM9YqvWGmABHU0XWX5k2bJst2
SIZdEM8v6livoFfk6xhFFydUEvNG7rEJJeYy9WeqId8YueHO5+VMZVRUHGTJ0isY
jm3Hl7ggNb3eMDN50DSPLfS5iYGEHsfVZnbGut8JrXI8AGixDVFmX0vd1bL2uNTy
1WZQuYfT65ywWbYtEiDRXgYCHejHXn0ba+IHhXfuOP6qCzbMNuIxdInVbYNKoP1V
zkMsEr3IWyXKX8uI3FaTR+xD0uNK+DGhnTaAcTkcUy2SDftM3hHDYjersDbZlXPQ
0Fh80ikHOxHlpHBLKYK0BRJJmK3P2xmcraMZlpQPjLXEC2XwZX7qmCqRe+UXthA3
nAf/QsT2YYKCRBb/UnG3NNLhcH+ev4xnnCZHO6/wAvnlx6nXeMFpUdI8K2qpq3+9
hcoenlOOyTu0pkfEn7VnF3ZJfVmFlgGtYrQDYT2yMHlFse6xzCpdhh2tb49zg/rW
rIXm/R8CRLq0DSigKc78D+VN2gD8oOQlajyxYt0c9+zj9r1QSQ9iza84FXnqK5bv
Yswc0A3u9qPZQvtJVJ4pP/hCL/LMIZZnndpYvkuxHykPkDpwIVtZ4o7k9JHjztct
yrLc3p7LnXvUYkDubnxYgop0m8lbdGaKXPM+mWTF7Qvk7FveWqQ/cUu5raj8r+V9
5lcYipL8xJYuR469uKs+samgGM1w5QoAQKw8LN2BfqilQQBitLdcVyihuCSDkDe+
4TBntfTtZu1yJWVnX+sRSOh+XUHaP69+OPy71XynpIkAcXuQC0td7wCIPnMmjHVK
r8l94WjN+xXSe/wTVGVOG/y8S9mYWFvGnfpDrvElEQ95oIwAviWPDu1JNIeWuKbJ
xqJkoaLA+qtTWWp5ibHb2n0nnVCO+JubeDSvkvzs3t+ZyH05y5ZM5zpQJfiWgmg9
nJM5d3d/xB1ncrqU7SGLrdB5E1YM/D370+jgIVaNGldeY6EEwW6jToU03aO+Q7bk
VdvtYkMR0LFxg1YshwxbnlfCDfJkhalYf2fmFo6AUqwbE2/s+EITycg7z+5cw6zO
3xlMKyfAw64++j5GZFpWUm+dy6mXCm6bZbsQ14GgkLbYRaSqAB1XxoH9OB1JrQYX
sKW0MAO6ynwWltYSb7rTJqAXcgLxF6igw19VjQp3WOaLAAfahzrbcx5Uf9ToMsLl
r+H8Z9kXy9LbIVYDgLylj0sGPvJIfuqW0hFloWFrOq+bQQCrSB5IZgnkAJ7H8CNk
ncL0r9xedB8FdfUVY1pAFfDys20EDuqpa7/hEoD0F3X3sF0qZ2SG3uuhs6nnMmsv
QIFn8m7GtylUdTkIQmf8eqBPacfsLCyqzkG1HYMX4QafKQmUk5f6M/DZkBvI70hy
t7GmYbMVK1RU6OhpEE7zwFrmhH3goUB5uAKHtaRxCl9XCoJL59Do1On352BJM6Of
JfHGdcB7M44ihiujPQI/X0t0QCPdOntZJjQZNs3pB1lAKcHeuiQwxhMITZcaucdS
yjWyhhLFS0BXpxTyA6UVegtPfIA8i+YvP7IL8FSOhbNDI0NjbnwmR7Cv2vii9IyR
y8Hy5M7fsA/0qfPwA73/Vm9uMfo7owkqveqdtqfyu0WS32wZJwKhIuB7WSwILtJY
wkECafDYNWLhgzHHtoKudootUgppGXIK2hFfzSIo4k9AA4Ejnc8E3WZKOlhwpAWq
LI/jKuJLnbjwnUr+md3NKgMM7NHpX3kogrpGDbVIn2eGIJdFCcfu0rd0iOxc0tmV
SM4F4hRi7VmwDQXeWg3N73Ae4XSpqYu/fr3Raws92w76eSwCIBthEd5flK6SZGPh
5jrha92LFQbMGSf9ig+oBpHjbfgqriSQDSZgRg1iPRbVPTPIJVYOvT6hc3KcDBvj
1zeYWFfkqvQDQWiSfB+RtFohsJqpDO6wmQfa7MARlRKytJqSvDY63OYy+KljsQw5
yf1x4HPtO7DD2FTXE4GyLjFykrxT+n0kjhwfMLWQtstwTNxWbIeSz3EDMLGltsHa
zX0Qd1EFdm1t9VfJI+DkG5a2sVpIwtTQZUV0vPvJ5Njjp7TVElRqI1NWUIrOR7ZG
jnUrqG4YTSDJ0e+pkaZ7t8QIHYGK4F5RsGhxBrOfLZUk4iosYgrOjfj9HLalMR4G
bKgubJjPn7j/HMEFKgdBkrHC6s1BVxQTrZx4onaO+zE6fSn79HujzVKs6vv1izAP
OZJk4OX1eoWVUeQ8EAEsvLEuOXsNGMATOFnqjZYTpgpmdy6j1g4WO0GeBU2WSSrn
LDTwWRAnCfagjAdebnOFJdsxq07GXJyrh63RpxAV8QMZ0Ffz+Pdnpk1S2AvM+MQv
zz0IlEAcxhNdWtE1AObyF6WE5C+ESBU310Qt+ZrRMze/VFEFxYWwmBrfbk3GF4do
Z1BnL/tOfEYN4wT0W9Fg3Y5r5jWvFZe0w12oHnKbQmw5MrzXCAajc7dV+/o27tfG
s2IqtroBaGiFLUjrZYB9tTbTdmu7bPxdB2MPMvHPMO0RcJjEMPEqJ56gJ2L+tKiS
w2uws8gGlf2861heexZ2xo9UXjdnRuQ2IURH8CYX2a0bRwLGaaHT51nYlNh8MFco
mgTQc1ER7whL8MIAQJDu76yLZyj2kkOvDHw+0vDwJnU+KgO9Ojw8NFCzZGfsOx9H
CvRMp0Vrfn6MN7bjBuZrOwbyR9938an8r0VLxnnoN1DQfAmWhnw5FoRMJMmoWAWQ
5eCsfErBnu6uM/C4Ut3libwV6tmzOulg0fdGkg1MtgX/npgrZcMC0U3wvTWQuLJq
YZlo3KbrtfS9tZKGVRU4FKiKm/2doWk5EdO0F78uzIuFXt/ljMaVjjZZJgf7VKSP
4uUHgZ5EZ2i/Uf+t1Gi3e/Gk0X2nqU7OUKrZYok6dkc0T7PUlsBKhhp/FLrOXxTn
ixmpgMVWI4K5GaK1vNkjhzQrmjl3dWPOQh/P+TZzdcK9VUblkyQVZSaANcHz6Pz1
sDGBb2Oe1w8Larp9ebh+B+S0CvItYlIY29XxmpZSAvTouDTffrW8d/CHqgQVrgaZ
BLo2hUBFqtmaEjZQfvXh2QUb6RevAZBrcA8gsuF4cXGKqQ98wY1z0avw8UwHGUmS
iL/jAo51Wd+bIOW7gZML4W+f/cdmLl2i37J9Fhs86CAvz2QZrW6WR3KQ849gTyoO
NE7dSH+HV4MyODUOymNzdJqTiqlZCgDIibaOW9MeKOF8pVMg7+dKOSTQ2oQs5v3n
KyNM6uHPsG4vcgZDbiV/MW1HYJKsjrO5MhA0sMayQn5U107S9N60foXD1rqNTWUv
m++S//rMNP/2uRseyzub3PMMe0sJ09ZMLCCWy8vyFmcwiQ26KHPccg19UanfrKM/
s7eZ5IUX3XsFF4fV849++2vym7xYLkU+ZSRC345mMtTAV60uUmpgy/hYlP16vkWg
Vst4Do1n3rtOb8Tv1coShA9igimSIR3rGa/libG/eQZKjRaWGof6T0zR8yZnnSWi
sRgxcNqcuRBM9QpCWC6MRrzfymxb2Fkw8kV//LNPLPughuUMja1fhgqtanoOgS4Q
n4JnqBk9o1P18hLWI9LKr0wQXCoNNSqEIYvILnxCDsjPkYx0bO3S59crgE21WJcl
0NK491heHsrM1/YCPe0zU1BONoAGZAYD2sWmgXvgpZ4TGDNbjBRorwPKhgl6xgE/
sDJ6YFPHbHd0kRF39N5o28Gc2+jHbrrP48uS0kYzzb7ZO1D0nssQy/XuGjWDnVQw
hSOl5mNpTjqHHJlyPppzscySjemAN4QKbLXfMNh1ZFceXWR96pMeBkRzrj/gBB+1
HW4LWKSVr+h6Nki+S76PoiMnDuWL9tQ4/T0vCpITysDT2iQcQydzq3ySyn7N4b14
EjRlBblua3D52NDRCHCBkxSStNnt28svE2M86vES8nkl9eeAGRY4qpeQDCSQshn7
SxYM3hrI/pnAWpWEY9i2vLytBgtZKlL9YgCx8NBcQHaF+ZDoey7+WmZ9VLDxXfSN
xCdPLlJT+eIQbKMTRpWQF0QMY8inVOD56OG27mq586BSd2OUsMmY1FZANqU+/953
qxmwN/2PgY/sG2BXtQzKTPpk5djvqNp1g9qr7Lo/Nabu2Rxc/41lulfzv9Sca23j
oxpSVrerWxGYzm/cFvkkVJH9S/2ekobR306u8bISh1ASVdTx0VBJL4yPvsDR2aMn
pndu1o4Wnly4beOqpflNVMi0fYERkt/l919Ypi24ITuO1RWwxcTtxOOGfkAg/LnS
W8Jcy31vRfvn4YAhyjoOlkxQmNcWH6HvUGxz+wG90ExHEKxJf+xMl2HplbAL/MIk
USLVOGVCoBP+oyua1yGeZLV2RhpRaqP+na0RKtrJ+FtHIp6kNm6oPLw16pPZwusZ
N1uVOFllgPllK2C3sCs/zKadgdb39T5HrPptHStZcbCy4BqAzxEICE4ZdTZK9kQ7
Jmq5eF9Yi1REOMd8sEHOTb9jyhV97nGmSr0QNnlw0P7qvy6bdbGpZEtvBkvFWERU
rMKxay9etTTf0gzHu3+nOIXSuOq5TjFfQfjZZBWy1N9tyB69vkj5eyIu+i2MJhS/
p9XdYNM8IZtAo7aSdCWvpiuJIxi9gur/GDI7qjSK/ANkrycS7PHwPwp9Yy1PJyRk
2Ebm2CNK41tkxsNv6SZSJ/ccsGLbmLGr7PP+1N8eXsw+oScWKwZN5UDegWNJz8vw
4ygSfRMqoQCIXBZOLCmQwv3KCX+4PdC3DZdJO91vyMcMHMiUOYCHC5qR5I5pyLpa
UK6M8BT2oeM8iQ66QPd+1iWi4CuYncV0THxDwIE8zxB85xeGW6ADb1dfAI/ZKZMP
gYld2dS5/JHVeO7jRXSgaVQdrkDph72a6hI6aKoCHPXPoyEjT8C5DhAJM9Jh1bL6
u5H3skZRnD68xx8KrMeEf1akor+FGhqrAjftS0XyH1yOV97KPxvTQMBYEUk5erl0
sMK7j7qui5Gsw+EyEBmCQzhWZ57kqBwQcWeHM52GShhf8VvAelAEYkm75+/rwNlx
VR99DVjjuDWscuMwJ9gBldQQVt/qq/oiQ1Hy2SYx7bTWlUGVBCUZq94ZCdfBb4tx
FsecDLGbE8fNIHE+cyVq0U5UBh+ceare9TP4Nqu8LKNgI7iZMA9qtaN/ytRZlGTv
0Kka8A3KOxENqb6FTItD+jUSIS6tWE4I7x6DzaIG6Rqq30spU2AxQLOWT3lAlyG2
WJg6SDIC7I612wN2Ir67UwnetDQNeTpjfaE3nxoLvSymcWXF/lAdA9SVUdpXhLwn
P/IoBilsslRH2jH/POWEBrBNrtuc7zxWadkE+3C5M7ybaHmOp1VNk0LbkncjazGZ
xZaUjXxfMj3jsyAfD32QFJ+aMP6gn/39RjasP52bwfPVM5yeNrGhQZ5K2jGV6ihE
s9X+WbLmiCobg+JEK/Y4LHJJABZjRVkixXeTvssk9rzNrwh4DLY2xB/07XEhrawT
d8DDJlX9Ve8HRcrRSnYmKKBnECQLyLiHGybAlcBwY3HKNzvHONguZkTcTKKSHqlb
sCS3spRMPgnyZvNRaU/yPgu4PO/ZswVD4I5bO2fgy69EhGmH8Efj2FwY2zfxhnqN
pzI/WzvRb5YM7AT3QWL2pWl33pAcZGHuKQXTQ+juoIvG/EIJgneFwGJJFZqOB+UR
y2kb+R9zv8Z6GHeScDVWCK494dv0b4uILnsSTfWms05/o7GvTPBMEl4Nt3YcYUGM
JtgzfNGTFTRH/A1RbRPS/Eitmo6UvgVO5hDfcNCA61NIv5PmBZnEbwCCzUNYHfGJ
he417RdclpOBpUcD01Ls+JhfE+zmijU/Zdb0/P7/KF6Ylp9KE+jsL0QxEA07WKKz
VKljhJoTx//OuijqNkEkjd4SsugP3tb1hqbtjpIg7rvdo5BwUkHnpqLnisTRp8i5
yo889Xbwc2fSW0EHfPd7OcafBNJgXtgnXx+5Oo16CezLgqk8lk5RGNGCCr2aQtj9
4b8rpqOASVVVaoqoBbvXZZxzcmvzWmetBAawvBGvl3PLUDxd5ruo5bgLpfdez8nH
ZG9TfnQxjjoQmr3u3pxDSX2AIpC0ZdSf1bcyMxG4ZEQHXholroY4iKOZPkhVffw3
H5NY6sirdfwFv4uJKjohbitQvNvXXJ7TiH9XSzXeqMCAFCbgARTCvw+iuMJ0wE1Z
9KajntjexrrIdF9VRRCVkT0CkMTPsCnKxE7HH5iSW7My6b7IbmpSMxlsT4UJVDR9
nj1SqdKMqmwDHqMeT7faTXbIDIDVeKo/81bU3olLU6VC5oMje9xeLyTYhetmbK3i
849JTwdzpffmnmLghO64YrrWg9jIpG2Ktbrt7vlbnCywfb6xczA/1YXxeLcqoCT+
fm1PdUjQM2NjwW3xZSsmFJfKH7DUigS+MwbI2pAmztfNtDu6BW1O9YvoJwXcQa1c
V0Yr5ws31vGPTlE6JyShVmXk9X7L+aorzDqz7VUVACC5eQRUtG+AN0m3WKmMkiul
uTqR/tkiMv2kXoTYNqfzdT00t9kCYjJTaQCWdWd8HdQuEG8llEy1julchAFqnygh
W2E7U9U1K7s32BsaH3uVDRCjo6yn8VL38lbE6CCoXjE2WMw8lZhOTaEZypwdxIax
WvROPTuUFUuv3i/ZLZhw5c3nb+Dg6IKPyc14r/hg8xEBdAzU7plsW3KIDPyD3u4a
ghH9UhDJ9HVUDqrBURGAPrBIXZFj0bkM1EY9ZaC3alt8CZTOcLpqsA4nQM2vwhE8
tAsIfskLXiE5WyoP6+jA0k5TlyzsxlVtzmjysXgJq+6b/yn8VVJEyqPrwCwPaX4X
yFA2j11bg8GM24tnYnNtJhw/nmQ+E5l2F462Gxnc7wwwdcLmQq4IRsdsNJC7CDEg
1yWiXWtRXGIX9XgE/bCZtEntY6SqxL+mTLvm4VSuj6RyXt9LGXofKYfuyHZVWR4R
VAVsgwA4HR3OgF4alzXvm0szW+3IuCGRsgdMZD5fyf+5Dwvhl9aAj1rTwHCzhqYp
sZkt0jDfwR681Z6Tn0CQ8Dwd4m/PccFW6YL22sAndeoTzEWQTMZ8V/xenGCFRypW
59Ax8wyNS3E42vZq7Tc14Nz4bI3WENvfvn3yAKE0spwvtAfggvqgJKbWWLZcKvpl
DUfI4K5oVyZdM+GJzM+NLAPHrzAgMZr+kiZcDm2jVp32tX+WQhHEXtV6QjaxVp0L
iIVA7Na9XHo+5hwxV7EZ+YDjHkW7uoWATxKo0M+vZ2upZYJjNKC1jr21svcLa2Rn
fzLZFAmvV0E/RmfHHT/fWzOF4gB10I68WVH+S4aJIDlP4XvxI60x+786mJjf5N4S
VkijZx5+ne9G5PZ7/469BI9Z74cKdBvqnT9hPizHZ7DnUVVE1FkHEdwAFjWiuTM7
/+NTaWWOpB+5uTX8tIpmgUt1cC8CuI/LuPp6QEXdXich5IPYA3npYK+44gvLvtii
klZkHucvQSl13XoIOAHPS5knYpleP+8EDUGFAkSgZWc51sxCJZjpu33WNO0Esxn6
K7lYo0KC1pM0RBC07QR9GPJNZBmPLFReuHJ1C7WSAU7PIvez5g0kpm8/g7QAEAeO
qXWVROGrnBsEW4Y/WXAXOqLdJtRz/C8SFJy+3gE8Jp8pdK5Fxr8Bp69nFdbBmMkN
Zv4xYBN3LTfJiVUvq3qpvZ5W19His9dze9e6QXr5nkovpStsYBD19W0T16txZ13Z
uw0SkrLlSTVt4jkAilw006qzX0qBsAaF6pX47DNrEtOsWA/NKv66XuWma2rMMKPb
m0d1ogFYaUlUjYIq1le1fmZ4uKFNBFYLZ2uWY3394kVcOH32jG6n72rWizh3lOZ6
GKhEC52bQm3FJdK+9l0ZQ29P7g5APCnG2A5m9G7lw7Zcewt194aScxhNfNbnfz7A
jfvFPx3RKmMd0hRewdrA/1I3qZBYq6/eGENzuIc9kcfNXP1/C/xj8q5alQGvJbBi
IqOLAQ7eJSGhqytYPGx7i70Wuha4HzMEY8yE+3KpXS0REAQggajZs0C3a0fFy6Hm
mKHXCCqV/oZdw46lTV5L8M/OEbz9YtXwC7y2jDz/+X2pp+Hx6HRuPs/+LJxG1jUM
NDhIMVwVeuWB932uy3v8jrTidHxDkPAJYyahMW5dqE/WrMT+zU8woShdKVLMv9eh
+vxpqtktl6tdF5QZR9gwlGUS/HPr/CJK/nJIE48Vsrb5w7BQYq1GWPb+GZMFyQ02
qcUOX6PbbbarV65uynWBKbBL8FxRZDa1N8J3MUV62/Bu+FgD9ml0PDtDNN8vhH2E
ZbbDfWfISoh1mneQIrIxuCWy1qbJY9cwVh/KwGxy7s6qm3GBNvdMqqc0pSbwDIA6
6aMx1MXwGgQs9KTtOCGOF3CEmeq/fhu7D9RY2VRTYRKX2d+lWNlb/NzAFJJJZiGC
dY7VpamTM7lbckRGcRFv3fpUPi7UlBLeuqBwKj9zlajZSb4xMEg8B0TjQ7PgUMR0
eBrq2+XccBEopSwzYnqQ9N2QYp89+8x9jXaZg151aSxT08JYGX4T6+1gvnKOy4v1
cY+YORrnVvKGGJXY29FMfVHNx5yflY3aoOgHkofY5N2oaAPSssYQqvVB1JnJaN2m
rMePDfl/M6PIBLv28qTz0grYhmQ96hX6WfN0xWlSxBpcwuiJX6/UwNiKIhDCGVqo
0PGeVaw0piHc/FxKlDvEM9JDGzLBQ/0lFa3mSgMF7MhWyEkPweHKf7vEabS/dpfe
CfsXEUrv4pPuJ9g0gu/yWCoR7QbQZT9RAfk8522I+8FbGolPAedJsDTr+veTnsEy
NWlGBSrbBuRjhvRtkHwptD20zfPaet1+UVTb4aczl3GDEnrXWQsZl5RElM0RW9Q+
TIXafJFDGVN/9dGPATRRG57fmURMmrSrEr4+6b7R1QlyJ81HrUcYfuLjTneDWfD0
oZepQ/EsIpwedyQ1HxvDB2E7HTSWs+sSWvD2V8XaskP/9/4/1InCv7a7RhGpknoO
YfSS+UZleZHVDzvYoBBvuY/Kf4ngnawq780lssMnw6Bmrq4tMxN3z1zVK9ZrQ43A
pCbptbTD9m1ysUQC3eXu7CuXNF2AYIwQEsdd216Vsbnb94LsbvQoX8u91Mfl4/S9
dFao0DWxhP7qXpTaXhTSFvpnHwhQIuI08bVFVtTxG62/FFUrugeyLgTMv+SPq0dk
GOoqYTzVsnD/I0jBgi7zysXQE+jrT+OSXQH6Iy8qX1YTMKlbdjoY3eqm61MDKEle
aO/Y51NefC1MhzGZz4iw1uw1bgXXDoGHvZN69wOYTyeqWMQetFV+qcw2GeC9hE9y
+40WAkZ4zvlQZzxKjeqN44ROiR2kNw/oiqUurJhLkUfNc0U8z5Hr8lmTSFcCDBCu
QiIZeMoVB/DFODLQC8saZ3g1W9UPB5t8s2UbkIsl3WUnXbp91aFXlmGRlpbV14v4
U3AZ4YIcXd/NPesuxWgfFTCy66yB+mmQn9Uu4ept9p7i83KS9/pLM3ARcZdcuDwP
sTXzXElCvHRVOQjMoQMc8R5cjrhj3m8xclEvpx5NKc9zD1UUCyNL4ie6VfgRHdil
oBJuwJF9IKsuqh5gz4aM6RNTnyjFAoGOe4q7VmItsYE9dn8WzKF0ddVxou4fXGBV
8bTuMOsXVzJnFvrNfhZVyXt22Zob5/om93swnKILM5InsenkitchDP4rNLl2wmeC
vCUfpXufiMR2EXK9qa3BIE/SAOfCpX9/aV+XI1myNA4GWUeHRIGJV/kQ2TayoN8b
GWLipgDZ83NU+ASJCUNeWyakYXsOigL6DraKDfE/MTtU0pCnLQlLFB4zXZARslko
zHZDIDvhV00H96574hmBpXn/TkmWdb4+MvWkP308sYu+aMNj7g0Mpu8Yzgozjjzm
3LOd+AGl1KiSyh6OaYeF7Thr+0XD/F4bSeiEYk7/qivAhdgOz1x9mX1HQIdqP4s7
vEHTMAzMyLnJokyNbUMujMBTE7etPjasJZOqLbT6fRarjj6caqzl2vg3zNjev3NF
87wxRVODMyOPLAYnVbD+t3K5rBJDtc7NKshNrkoj6hJBIBAuUtTseCXgajJJnv7W
i0vwSlz3CqL9b5YmhKpDDusGvX79WjCeUvJoI3rvjuyDyrbjWwFLo7ORNwPq35N9
5/iSGjNtvWLePeRlsjabrQPf6EmJ8veAIsdQ5VrOBlf4ycfujzKzq5uWUmtTvQUO
uqt2mq/1MJRkKY6JOjm2kRy939CLt5d149lmMCBkRf/2qIHOpEFIZ+Uuv+Vvk6VE
H+G/HWc/Xsbt/wirxaGsgm5LENEVWYJoPTgMOjDGGHgAxkTaySQRv93+UQtL2qOS
mZiFBgGyi3y/Cn1iZNBmNNmpU2YL+lKqrmn4O2217+nhNDQeTcWYMRj/6XbQUsbD
ckNkLz/fcW1p43VTkoffPrmYzoIDpCQRwsoPtcWv/iQPqse4FsVM2Un8mRN7XJA5
Z0JaPx2LY2rYVe1PV9hC2rFPVAX/9v0MfCS+8dZXyzSa8UIs3Bi+Z8xtR00Oz3Pj
0NmwouJvvPOMhH33r7uc1xJJ3fOApi90nKpn1XwEF14Wm+4Urw4RxDW+MlUr9U6z
+nBXrIbToRVUNokixD8X6rVIVlbeL5bibCmamMFK1skTKcEuOeR81kw11pQvMmmi
Xv8nrBuVgC3+ZmLyohkpiuPLnMjoy47TwpnooKYwRQncvZLPBSSkYlTHvSmX/9U5
p6XAhftfJVRR7LKac/LSrA56IVS99Q7tvufTK9oj3JPjQdqBNK9i2NpoiT/dzy8a
VSAzacYraJyrcdr5TKYjJMnfYiUVWypEFEj0ZnCflSYZdBxdIN0m7E+Dnd4ApIhv
2mfXxIsORHm8qIw+zlVEnUeuCf19ewbXGt3eza9blksO0oAR3iZhNSSa9KcPpN9S
9JNC22XMxbAXWCi4xSTPMYzw0mikGh9Kx7ktMbc2EPEY27uFEkX2bFRvM77TpNxN
C6eFTXbQ9O1fhPvxWGKTx9N2KpcW/xFDzj+leCc9LUtHF9pN70oWghXCyuvL613p
Skasvh0WNNrwL9TK+vJ2WjRwA8hWimeI3dgLoZjLrxJFQnkjpkfj+47BmnVI76LR
s/RJ7ycLo2fXplaZgT+kx/H6XYx5tXiXSrzwtPIvtyBoFmCytfsu5BXimmalv0Lo
LR87OZy4S2B8zcY4076jQvBB/mNGbX1gmwqdzn9S2hZPAYydq5CIyZDBRt+pZHY8
qkkqD+1tqiHN3/DhiE7yzYnebDHJ9vrouOoqMBpXYEaiFvMC1TsY0m20oqiwGmzD
uhLOuDAlTvHoXp5SdpS0uaPDno0ctNi2s+tqIO41E3hqbtT1upHaKtWTSnHhfa7a
YTKL9MsXNMftByqhPHiS/fkVYdYeMPAQXUrEp0bd2MWKB+kPYbq/Lw25B/XkwqEI
b6AsEWxHDILpcvzHssJNayLwaW0zRwBzr+qE7ylChIpS/DaKrl2ZDejUfG/ydN50
VYvN8kckM6aZ4w+6HoYFbopwAQgnCHJMYxYQZuts8pLjd/DYNfqmQ0sqEQwFmy1q
aAUiwyUFxI47T8o32/Nh7/nDy4yab/om1sS0irvqBnQ0ldRoyQiwXMGJQZ9iKJfx
wTmAgrEHnWoXm/NPBHAU9KOXtSrggJ1D6X7jOswrHK5pZAmrCLj7MX5r6ymtNdis
Q+020TbNv3v+F7pOF2+lGq6zwzKGLYZ88bWmLRzcP0NhRDwGCMHTIEadKSQf6ZnI
fXS4Gwj18cevzO02kJQJgzOIeBh7H91UvMjxYBK93fHXSTE8sPoudGipDLqFQWiH
C+tMH1bQAzAGUDm2/kHaqTP7rq1hXU3f3C9X/Vnptd/2iuHchSzV04EkaqS9Kk+7
3nVPeSiSB+lDIyJLLKJe6r8+9sMnUyqRcmanmpgGBx6d/ZG0Yq8l9PWqQa/woFXT
1snRssrN2wWRhiQtBQHaCDJ9bhwwfMsB+NolGE1A/JNhyWkfgPaN/MbbaTErhJYq
mMxiNz7l2cTA+UwXtfzEALPyHh43uqXi39yISZlfpMW4Glch1c0vfukMg/YLDH9U
4cM0wyjMC+I7OJFo3XVJ/XzEWkUTep4srHOv0uz6d5TMF77XrU6RRwNp/rG3Cg7d
3FJ/PLsd9y1RzUgFdqOpb7Rs/xV3AQH1ydyo3cXw+QLgLOrQwzl6rriHk7IGng50
dJs6BryIE3gnwZ61XvRMBqrqzU9G0+O9m0IQokIL0FRyZRdZh1jmPjG5mHf9Tm0V
+UfF9cQ21DS4Caw60YWcwP0e1usOwOznre8c4zYN7REd6L3zfG6t7I3i8WxyPWnr
MOvhLqXEKS9NSKq51CIL7RG0glSm+p4zozSG7MX5bzJ1ITWze2VNB+Li395r9Nqa
EY9p5TVJMJ3/m8eGDpwQqqLwxa0rNqrLFuySDqI6CQbkZ0JVncK62a4D6YcUbi8K
iQwU1qG+Afz54W7uoGeMguSLUtohEahDzSAO0tRA5NLCoY/10ZzrAVeRSnGKpMEZ
6yD4MUe1aDSOGzYV+Ey8qZmM64aS0O/8ViXDSz+oNP+TINxYJq7Vq0HUuRWjceJ9
Gi5rImQagP9Z5r91HJLMXzDvPkSG6uDSxryZnu36T+MBbQYzva5X1H+gzmW5YozB
ZZtY+8Mv1NHcJe4mhZM4W37nlSnOV9Pbxt1UDGyG7mRa/LXp8+Sv56qPCEhcBiw2
0YH9HN3e+0HwI0qShe1moG2jKxVRAaM4bvtEpGePOjK2w4h0Cm4hx2JexuHEzK2I
9tiFQgoFPFHPODEH3B/SWoZ6e3W2LihVcS4YfLeJ318aFwDUNsnyxbD+VSbFHD9b
qx/0Zt7LgdV35Uwfvr3p2YL3VkzbmGOakLAOpP3ooIAN6kyhBdFdAvLEcN2GQuH5
inewg1gI36vUUYMN1lJgcNh6CZQSQeJ+LF8N+nboCm28ovtXN4+PcIwMQCn6JKcR
LiteK2YfTxBf1Ml8WmIzauy4LuA+pW7+qm9/xJD2+iQQLaaSGrky9bM1wyPH8kJF
VMIjn/QaeNMBtvzw4HJkpl6MoMsuO5sqgGpqMKykRPqsM4jorpV8lcXfQ3DbHsub
RD2mTxdq1xJce9Fjzd9OqUz+Ui/6+1Z2/wj+NOAEmiFEHLHJauV+qfKVslFv48qh
1vjxxxDO/a3ujL5oEmtjpdh5b6Y2txMjf2ZHZXC9YLtAm/hPUsNlEBkNpI/x8s0T
HUblqGWQgOPyyyTVKhDRA1apzFTa6xWL8FpmldpmRu72qgsch+T3do2fYQNokb97
Mbb+/ES94ltdsKRgI80enYxxlNPvcj8XGcU9AlDnmfgZO+yQZWOpoXVmKzA9NO+B
q3l9WaVTlHuDUSfRlJLBhRkQvZBKz61LgfmIhZvVzwz8w0JN6qGvBo9FXEOHGm0Q
vbYd1jTWJNlp3mxofoCah/wn5bbKtDiF37L2K2/Nk5sgmaBTSd5tD66OVKKhcW3G
xJchc5IJyrD3q+HlxRhHVTpLs6HuMg9Zfjkjndu1VqaFIPV/dtH8Y+pt+KszedZI
S6bqMdbtfC8delHy1FH0TCwa4hIF6dIbMox7zaCrn4DsL0B1Ka24OZYFc+X6zX6J
kivAFa8uQd08epihWCNdS/QE0Q8bodLQOSIe7LsEJRLQ9mjwKthDLCLmA1UEgpK6
HZptK0KMdRgfCyC+fyaUcN2jeF4YY/VXk3UjKjQjyJOxitMz6CFOs/Ma05MNbhg3
P8uXoDemZ5esurxwOK/ZBu4gWXkHG8/Vv5HnXoCML1iRBtt2SVa0tKXSRJ2Kkb6d
+2yKp0iMvh9QDBzKpqk5uupTo0J3ZDa97KetCal9tpuRqzcIuNXrZef31k0qgM+d
m7XomfRhyM6ajSZ6GuPMtv9omOFIxs+gSPbb/qmjp2E8dqnW+yTi9T58zTEzvEmX
z9zQzGYbGInFPZtwjpHvkT1tUh/nfMM+9ZBxBxV0stRDNU9MQiqUgS7HtcRjCiJO
NCsoqo70Qt71l0dX+LsEEYIIxsVTPmlCYFTeB+ugamCR5LXzqSmyBleuucd34Des
V//07dxoM/ipie2ozJPm5QYngU5E8DrVlfLzoi2nnjCmKlv6OJVwU/FkKkWSNItZ
ry8iONe8kVFuQtgjznP8AZPv1sig6UvUDsrPjLyXocw1/HkK80ybK3GA5C2u6zYl
XiRV0rn7Lk5mNTe/NSwzUk+j1GJAEyD7FK+b4Vs4FJEG6BbrYuIOoQ99tssrIOd1
liE65C8siWIZ5DScGVtnJIhmel+Bu3dK/o92aEbMh/LWFYntAx6VzLfHjxYCj6zZ
FFq9m0lIyJBETb7g8nu4jBkwe6+ihkXAFiZ1JTcrvkJC9RDP0njSbdONQq8wlNlX
uXuosTPBAmZeclF2RieE6bLJ/QBViAbZaCB93cXn45kP0a7sP7WHlL9G3cYkuzuP
gL8RHjrKEff4IfuWvqgofCSNxdGwLfKKSGhaDliM/jbNH69GoulzkjULCAcMlAXW
nE9+ECvPK/gRV/X3YPNJmnHaEuvGQuXTHr9ZxRKogxKKGqWFTq9C75G16i2tunQl
Yy9j8sBuqvuP6OfbyzfgljjvdMLcqV40y7MPrn9/CH5GleBh8hKloDc+bn7CHUlZ
XChC2bHXOxqBVzZtOTzFwnXwngZXyCssdk35Jq1klwZx2ooZX+TfihXG7GZ8N30F
koK7moiQ7+CONu9SMinBPDAF2w2ZcFr+ju1Dzgv1rJhXYUA+pRcZjln0KlOp4sHf
hacfKAk2Ci9U0mth7qWEYp0nzRy6XtR/NkIZ8PmYcU/J+NUZ5MGDVws/KzSos/QH
ZPzqpBuU6fZqXRrkslP13CaL+KzE0Zw15zxBNoGOyCDURIZLaWQ7Wd13Kp0k+RSu
t54OH82IZmx1arvLrBn8/51z6F/ysN4clqLh2oWtQ9+i5/hzj3BPpjrcO4ebdUnH
Xn9vVj1sqYL7NAJo1OnSFCubmW5gSKwnW+HjvyyoHNfY7zxmLaWCuYVZnjIoIzQ9
J8kU2I7wiE2vwhcD8cea+fUk3+Dx7NW3jGXeSsc4d5hzzm+B6x+T7iJnJ+33qUfd
nY6aMmWiQp8px7TghrFLns2Donm/Agu2rm9ARX7GLB7zDezElV26S3ImfspnEI2a
Ksbf8qPe6xVxElSHuGsT99efKxXpx/dFCEAxUAy5tS2en0H0GlLb796r0ZtvVTJY
L1rQeN8On/LwdYI+b4GMsqCr7y3Fi3lNMR/mdLNub6nUswXlNXJT8ZL26GjOY15H
OKErMF+Wv9tq9r1BJhhGmmErZ+GL9o8ysm7UDtOOyZFxDGPREGjMoytFUp5sDddB
ruiTSjOk1886ioH0fPb+0ZAurelOeZYyW6EJXXtvZDkHHOg1+jQ0svokWBQ3XvsT
+yw5+DwnvZBqDuvr3gjMED0BN76zjOi8gt+Ke/xzd7nxxAK2rbTjD0LlXAA+8uYg
kmn1uog/96DwGwg9YCX4yt4+nuTXX33v6vDHyl1XHDnKW9kcKMBQV0fJX7EH3e8t
yJVRZCiV5hHNmE10XCcaNV1Oo3KgpsVFVv5ocD9wVpWJkQMvexrSC4PvngPHTxco
Gtmg3ZozPNvlvNmvunQgHo4cwDOpUxqVD3piICXF4vgUCSzgoI1LyS526KRoCseX
l58b0lu1KuOkWSnKoSnqHFTEqodf8KP7+Ne0/vvvG5cet/KGJ+J0Ts+9C8tJPfL5
QNJF7jPlNcBNmw/zaOpzmVdsaP8F6Xp4yZdtA9xgI7pEoVWTdPLC53LSra5gCrnu
TvL2FudVuM8PNsrDpWBkeBTDGFKo4BbRslWDFLAmJO+MYqJVoYSSAvjURvbXUF+p
yAQwzzhRLQh3XECyfpzl+doGxHgSZmupK5XzQ5XhezaYqE2UB757y31PW/L0OVQJ
YFY3K8byKmAi/iDHjCvyZ+PiwHpvHwWVCf9/RtV+i1NjejrJJ95laBOKnwzHMQwY
XRMQ56KtmU2a0qvc9imjdM5EwiwkT0xe8B+nxP6TbFKoXnMvQ11l6YfF+28DvjXX
yzDIHjs4gI2iu50dWDg/zkOKYzUxMSiGe/ZSM8BRncVdJbL8EDW+DiSkzi3WgB4y
54laEL4HujsgSoOiW2fXVFh1AZryWyegUQ//qPMMMyAFesUqii/vgR+KXUDenbgV
5itl1p3IiVn7rgyYpNsgqrCuBu9A+U+O6wWzpRHRrWL6kmuZ4yhbrplp16jAZZId
QXG2Rl/zxiC5ODcmPfppRRlYc6NiAZnjOgKTu7kD94w/TanbWWPAmDrBNAtuImgv
Sp/qdp1+g7W8Yj0tdozXdlDNJdQ3ZG609B+wr1pcyx+dpX/tpYiFG3dIbJgNGRA5
nV8ged4p5zlXhzsZ71vl9cbip6mbOEcBYed84lgjiloHZd6zBAoED2A3NTMen0Oa
HPiNiGKLfLdb/GIC1bKb6pB5D3iXzus7Edw5E3xIdbaRdVraG9Ka2CkzkRx4KUsu
a/G/VHjjIwyYQnlzf7Nq8jRnY4eGgz51XbPgNFJyzvHeO6U18G8NI2V0ZgilzzEk
RsVwgDDzRsW1KkRvV+ALr7ZhwizzJLiDtJANL5VO2B+SswvGiEBoXJ0E/nL8zEnJ
e4VluO8U+XgQoV6b4ci1AcrPnlLTm7DYxNz9i2ZOiDxILksMMx60LK1eUUk5nAJs
6skbd3VUGeifygaNI81u3kh30VZDw042DGItERXG7jTZxqRMaQ/Z4QL0CBlTptaV
EIm9z2LK4TW1FUYV7Ps33Azl298pqJ9DybAFc/uXhguJpb5tGicxolAEiVnCG4Cr
fbOt0DNLrOu53hac1n0Z083shbE514R5uTIE+q85h760sYq0Yjh2PIYwxYSbNmpA
kqNwBCsPHk/mC3pZCOkt3XTFmAHuB8X9AQ3vn57zLFk/h1NQlp5IX5diZ0IBY63V
+Qhzm9IobebKNcRGD66mdVi+hN3/zjqZiY0MCTY0gIHW7rFSdvub490AXNEUzUKM
ce/bZ/u7mdmVsqRxqhS2Yri42cmivDPsqeWcbQ8AIJotQzEk4MGTFK9PwDy3Np9Q
Wz4KSpMe91gnbfH3F52nOYF5gEAtW6kSU3Ssw8zn+br/L86SiAJ2kaGpMogCNwiF
s/Hc+JX6faYi6qdqQhHFCEdPcxHINfC/lRlarypM7yuWJ8uwJTds2XV7ThRyC00Z
LXnEGhnEeiW+LM3znGiMN8QZLUtqdXIg9qW6MHsQGuSJ5SSsXbvKpgVZXXvhdZIt
HLc/BEAATsbE/wfpJr2mZPGzs0niAlcpEtRqoMZya4Im1vrqxoLJOv9ulnj6YW3m
a3P27V1yGyh7ta6Qs3O1jCeLqQgeqyra9RzCVZH4q8U7jbK4cCoqkyXK9wdJEKtC
iBVnx1QlFjmI8eFuX2/RdXd0Mq/cOlNYqOpTwCkpp3PEYR6KBW9gPGaL+0/h2Gg6
6VhD/iWfhHSh5I/BFrNpjKLPqwu//aRNKJ7O0bN+yTl5jSK8vRm/5sFq72zLDPP0
glwbncemLYYpBJyUc7pYqhb5J5xHoaj7CqwCXKKe9F7Azou8aRiB5H1CnRVH9NtH
5Ag7/juaDYkaBpVWHwuKPgx0iI1rMd63g2wO4pa5jqXLtz497z5Yper1bjxtrWAb
Jayrv8ss9+hT9GBjAr/mWKNFJxrBsykQEsToRKOaNtJ1ohVQ+k3017uofrDDDCuu
M5bp/glXyob8y3q+zGi4LQaupGDTljAAU/sHJ5Zw8ac8aXxPHYG37ySUs+c4eww5
BZbL37EDl0uIilkHo8KQuRUGGe0EUAXnH72DGVbX52GlzcQSPQcmrSUdFLB0bCBU
hp/yp1Fza4Inhxl4ktm7LWgnL7hdn3flq+tUC6dKYOWZCoHMvC1zz/xXYZINVazD
qRUML8lXGSihXtUEEmaP4EzzTNlt3ixCEVkwzdKLHvgkP05nkZ1YQBg7DcgnYuyq
NhQvZ3rZFu6Fzox2gsG2DjjAArkWSXL+4rgGE03Sa1hYDo/s7Kk0t/9vAP3B3YKQ
7s7w1jNGIwLxkhUNjhCT8hjJ9QeBQlGAqYrFXlVgijbNe2P2C5G/2QrLLLNhjUXc
sOGVsBk0EPRlp6Z1zRS377bAhWI2BzattR66aXxoSYR1aMQKgry81PgwH6J/gc2O
Ri5O/4MKy6MgB7IGB5gS6YAFlZNlxPEexSTl0oD8bvvoplQlUnEC75gfvjCpyzsn
EahMuePdODETYMsDa5G8K9pOCMFiDVjlG3L4b/C5PDoj0NF4cBWjbAdbcJyqIHz9
wipAnC7cVVXPVGE0Alf1vXDxrb3lrOrbPF/PwGv17WuIT5QcbqgCCtDzu1qA3kKX
O01f7v96OwxFUozN7Mf1Jy3U4CiIlD8RW0oIBTQyHx9gAveLoa6bfxDXoqVK4KPO
ePMACdAxVX8NT4f52OFW9JvPY1L/CclUh16YHxc4h7T39Wt5yutkH+ABgi2Dy8nU
wcWIbatxKEnLya+6ENL3AtiurGirE4pmU4h7Z/ygVqbJ96eUVNPkIPU/OwFZvm9J
jtnU6u7Vk6zDFPbEStpdkQcFW8XQmtT9bekSIH5hL6ayuPfRuw7ZTuDV/As99Wul
c2nLvBC/g4pd/WGSbMvEv8p5t9zHaQbrLq2U0MHFhrSLTY460VdQqWiVZykkkSdo
TN7RExrylWQ4NdmqqHsxBivk0DcyIJxSUaYRgSJvgdt0kWMxS9rKV95ZKp743ITP
PXl9XQ56hZIBz7vhKPCvAWDBKcLG7BzzpYCes7cKUAKR3ySkGimQ65SXkgN6Hzxr
gkchg7cCgG8apUD7arKMYY49qKC98I0OGHKUMZQXaR69zv2Xe5g8XcY9DoGfWjmI
BCyMspH7JqVf43cQ9H2RR4r2bQtwqTUOqEq1L4ohM6eV9U4szMQrpEzg+WMkuAmi
fAmZj0Nlxta8rd+I6FiqXXFC3qstduaS/+ebwS38h7tolyOB12mPanXZr0KNvIDL
XHtiO2CHiM9evJa8Hol+1HfUF0ekxK+25g6X9w0C/pVDaiqsI1yLkcdVIoGqzqSd
0PbD6p8EYTFoV3RLUvKhZtz+60ilI+7Aa9a/S514kzIwnmjz+mgGB+Bk/Prp/tPz
fGU8nRuHNLpsNfUtXly0RCVnOPe1pY1hZdCxw6oJqYIduDhRx/hSgVmEuw7/itkJ
bcBrSjw2255KV3qVJO7D/Ek8xVpxvLonpW/W/xaaEQvSVjVeLpjE6wKk9BwTsg3R
ZaKp0NncNynvmsuvg2TpVk0r3svVkeErxcEPIl35MoHsmL1VPEpyXIUdkbQjYGE2
Y6QIS0pVIe58+EnU7fUfn/x+F2CkLxvzxCBalx/hOa+MJopaP2sm5LpIejWGXdBV
nzycm7p/z1A6Rju75wd/Dc/QY5zIAysVPxf9S3hhYCFRltpKWgb68Pj/XruVcYz9
lZv8+skU8DVo687R6G/mMwFamCqktNQD3Od+j3CBR1MQ0egAu688p7T0KZ9YOd46
h8+AtjdlytQnUTFqO4k7r7dLf/mjBVoG+yFt16KxdCaKONC8W0sOejiJ1+UqsX2h
k4k4x20UcHddt4Ovc/xEO0/Y8aWH6Su5h4JsfK+dz0cGMzyhg6Vs2k383hTIk/iv
2iFvZTENmXlxiTnsU3uedPvUlrMb/GRJ9XC8MrSr0RbbeVr0a5oGIMhy06XhUKL7
er6j2XRnqi8X03tROpHk7GPi0cpJahYXS6290py7k7enOuQXDXOZWFM2ijp0Wa0O
XKcay1zISv8S5VDiwG84dgXN0T2jnl0fEbTKGiq5s7SiVN4ErMUR/ZfFyqmIDr0F
5VT8RIFqLqJ3UoWGCxaL6BprXoLdjzadeafyfrAd/0HGUkrrV/dPvIueY3SggGAt
PbqtFNukJKBO+Z4zg3QU3gH3Tk3P3MGoCgqrW0YJScmRHdJgCVozKSCza9OsYRdM
J5sISDS2O2DnGRK4xUcv9cs24Xm9wFGUyLYSNNGifPOLMUN6Fs1HVYrn6ZUzfJs/
fThKZKfZ7bpAhy6Ce511RlKHBwjUJuzAkFH003roDdj0wQfzJ/f9nHunEKaRSkrQ
RqwMGFT5kxppp/VMjujGGFwJHRA2HJcxdFpYkS5t1D2uV70MBCd/CjXvHjg5AjLk
abRFdxC1v0fF2ZubJqc+rIc9+qnqAggfBkftBsx5utQlG3GZVkHBUcxw+qF4XH3C
LncmjDtHde9Bq05edElgWdaL6a94mMlxlfPvGDd3E/tSc0M/4J3TA6c8oieufvWD
gTmCFp8DqLpGBJ62wX8UWQ96o9l5lGkQj6mbuOfcBZ8wqKqMEA/bgWIWMsopxopE
zN457YxKaJB87aIV6XsM4dDq6D/qfTuIIVzNvlSBKb3QOLkzbPM6V79ot9P24/te
581jdRdAZHwGeXEteboGbaPGEZIk5oLGTESIH2jDqfW1k/zUdOy6EwZVIvPGUwaY
t4bZX0I/nedS9L2mwwYTtRJhhASVMTYFYLMVdX8UisTnzAQ7+SSDbjUqeBDPnm6K
kSsX2ATztWzyGAQWwFzcV9IhmPkOMY5SOlpbUHjb2DYtrh+alQJx44p1iam3ft7w
CZSdmnCgZ1q6K34zRoPUHYWsO0FjVgz6ZrZJwZZ+Hp2BbTWvz8ZQNNXfOjt4WsAb
EEPYJ+W/Pkudvr+P6fpE9rBiKXYqUqslE5oCozUtV7k9Stg6dv2Y8K6dknQB0bb/
u6PCCzwVwz/8O/U0eL5C6RArwHn+W8U9+8JArWTw7BM96kb8XlGAXfqDcBY+8+YK
xBcyR7QGrlzfXg54/ix/CFDxKsT6bwWGgydjNFE0AKhvHvE3ck4fcp+paKB5nnU3
V7V96DROpyP9lTXNw5sQlPaQo7XCEs245QX2crn4dHrr6D3VW55qmnHjMjExJZ3T
Zd4bS3/4VzeulwpOHZfCPUQUzfY6DE1JW/qj89FTOS2DxSx1X//gBDuUx0ngCdyk
G2u0MHiNy/aF8Qm1qclbYPS4zfRUgZL+0liL+vqpYOTXhSeIJe80jW+5Z5Lq6zpB
IwnCs9p+4FFd+0M2Tuwnv43gR0TwYWHh0YGfTWk8pQI3YUD/f55IN+706D3kcqsJ
+/UyLTVKXdk5nQLCN6W0bzuwbZJ0JeowGKpSYQqnHlR1yU6DNX4jtCx5Rj2mu2d5
/I/fdBvw7TQ+xvm6HCP55P19Z5mmaNrvB2zWgKlT7/7HG0rzOvsTR93tsyck4+SD
p7ACGYVQjYR09O4mL3772HcAO8PtjfWKhcKNTTFLstN1aejXkY3IT31dl7pO1BKn
G3QxglIhPuLwU5Vj1GAl/d75nyRjYqkWrQArDom8f7Kk/QrdfyJ5y+Why+Bb2gC1
BU0WrXEFk4G4+k2Bw0WlFU+n1U4L5Zaj4Joo8h7XDIDOCZxFpjXbATuYJjMndvBE
zpp/JVE+WNfJfx9wicfTNlBixTz44nrQYLYT0h8J2kcY43evILtXoxc9kxFuaw7J
KhBlXW68Ai1MsfT2tZY5m1nR9uY7+VBWQgQYf502vxnTuHavIph/cLN7WlWcp1Dx
fuvgjXJWqL3NBL0eHnighRbqwfsTmQlrSsrIhE0l38CNbuxmcOEz0kN5qxkH8w2w
G33/PFfhCaskGb36LJZwT3gDQmXcdoIioxN0rXrEn45KIefeFatugeVZ0nlRBPcs
lPJGd6x+xJn38jXUwdETn9xeHi2SIxY7M/fZZCEz2S4fWE5eLIL4WFOo4qPSB6by
5xP3W7zi5dbSYVflCMHV/Gw23j2DV3hpCfKOIs53aA0UN0ujwRBporCueT2msXsE
xxkGIC0CyuzDrwiqHFE/jv1zD+6ow76+iIzWN5s+Oc/CGbPYa9Y916rNq0ceFAMH
kBvsx4XQMWiBFE9P7NpBncv0ltzjkZyUDzb530+MWWVOECQAA6GybOc/8H0xUZUx
uoEX0+vv1cW8Vb8e/3i2mKc6wY1FTrwVy1BriMKzWa1BjzWJJPHPgX1eWq+WrqC0
+HY6czheN+Cx6G0mqj6MzcJKm+rL4+hiu9ZUe4FfXKeaVmJVJ87rzMKpYmSMCQvm
w6t9TtHx80c4svvWQP5loV++Xcita0/rguAfejzSHNaaUGEx4Ro3BLtuGFRsbo3v
YzccJQ4B4GGb2vlElgd95ZvOUX/vuOlhULlNPO/xergKPzkg/v2GwNxuyTb1lxSq
KNajU3Pfr55ON3crE0OMAYUcmlgRZcPXLa1XbrDw/IG/slFuQ3OhenoyYiI9EZVK
8Ht3WOprGwNBEBrt906zai9SOrz9h2XYp5i8TLBGL8Q4fsvYQtq4CZt7z5hLdTdH
/8TO7LUpqq9PguBwfYQh5x+LloJ6IapAatDhIjUoRqK/ktpDwgOoEkP7iXj6R86N
QtH9fcjSIypQigaco8GHEKq9KpRhoLv+UYNmIvfmwj2TD1+J/5n6ESqWsQnI2m0+
Z5Xt6v9dazNoGlKu0sFEma5/KWI8pz6Ih/cbgMY08W6fLlsHqZJd+2mNGC/7M7CV
JzZPjoR2AOYpXeHd9GBHTfiklgaZ58fMVrWcEVrAwGVoEASL2CCW55IvZH5vgYMd
1hlcl9Cvw59ocMNMF56fnL7f+dfhr3L8uY9WCS9r7KecRWtgZrHAWpW1E5OGtGac
3Wx2QiwOKRx9YN9q/uN4p3BejJ22k0AkzUveGvPbb4AwvIq5R6oNqOWftcOegVf1
+Fc/kVzz+Jszlo0c8C7qeVN46CW0e0HYV2AgU/2bk+hULr9XNBgfGxN1PJ8oC7C6
Ep/4TRSMxhnXroiZilLwJRpgbrleGhs2M5B01nmqvkcrl/L7tgupp6PAv+00tuTk
NiOaFC+PM6hq9CIghZMutxo04tVuE7zegmrYM29GRlOIYHcHeRli6AJWB8LhqEZK
bdogaoWY9wlfYerWF7O9EfTQaDKg4dAnnKJuy1/DwiDgerY6dTd4lt/BtK4tmuP7
NR291CXwOezQW6g9PPE4alphJxSZIqUVo2TnVmKkwi0XYzsXob1Pto/ClAxbB3/x
/1dY6V7g/fukomnQsu6Sh2Wy3a7EiCSeyYBoWTIglmWgrR1+1jOpUgrk6C3mVLvt
d1hp9lWwLcTnjBjBCFb/K10n2mrUK9RFm5swvvw+YNKuiIq7FbpN+vc8FYKGVxBt
UpTuyTpLphTkqeK8kJoIk0EywI2hfQRKOA9mLhdH/dnizWkzhkQ8UU3l9ubA04hG
3kQRxTMhWXrh0lANNKBMtW77bxwdj9kh40SHpi85S37TyA8lMM0CeCYdEOALPj8/
wtZpnC9EIGPyfwRqkxg1Wf+hEuaYfW5eAEmPzhYRJmGRFAHkuPQyLCJbhUB3j37n
bumAZykEm0T/QGUVAe8yE8JkfYDs3Tr31PBhH6kAiS9mtM4l+pMBitA1zoLh4X9b
TcpHTXQGR8sfQv1ITx1qdmGjtEWYgxviy6k+Ie1mGeXkqooZABAoOJ7LoU5CndI3
72+3hKH88uIp4UVP13aSVp53uh2qglOtZx3YGs9GTormknLpnxSPkmKL4A0x6gXp
0/EAfAMhHnYQ8pnk+lNuSFNv0z4gzvLWoeAagrSPmBkIYVILOyUBCSQXjZpEqYNO
cXEYPN7zbnuUmvt5+5y9umx+lgQpTo9Y9D4FojIfVpkKsNHXMDmdt2qk6c/a2NCq
YPIZNHT+7Gnq0n5v9eL9+EsBfZAMAEG0CREKIbLMJIpNvNQnqlgcnQaQCrWx3sLm
g1a+libCkdITh7QylAGgihCMH6JqtXhN4Y/ij8SAeswnt6Nh21u0OpkHkDEp5jQZ
2yhqH2YpunS0yi6XMiRJDbeURiKjB1e1RiQWtMRMg+Jtb6P/wIfnLfKal5K//7Jc
XrlodRHKAogXGQAOdlCuDITpZBGgAm8c5wv7S/bpOCrKEwCGybJYjYzauR/v2vJ+
XzKhwVJcWlHEdII3ABwcQZEInl8dCoa/VkYVs7G7RNqlm/6Yag4Qg91K+8PoHEek
iFVV9OBzo5Rw8XhsvBw5F8eVhZTQqLN9BZhrZ6jcSa4VQhuhtlRtkbhguTM2ljqM
Sr6vI8S1axaBoF9uCRaHwWVv7Nb+K66jlM+smrdPQhv8rrgHZKwWQs9E3At5gsqE
IJ6pT84bc8DOWUZeMGAbxv92lD5Q0doRRhN71W4PHJ/2yYLlxD7gqrUmaFhQuLN8
5kun4IxsjSvE89q9iWvY4muv02CRjEG3v54Ob8wQaibNKS6yFwtG9Bkb2wx0aV6n
m0uvXPoh9PpOuRh6R9imJLdcC7ypgRcpzqDfErguAH3B7BwMfnOiRdhHy2YwPIro
ocS9xSiMheFalkCwsLTFfix8v5Da7d8vdz4WK6WawaWWXB7YYOinIPOF811oVlgl
nt70lfRCTSh8dRel4obqOaKJ4Ly9VZnFd2dzCRMu7Ryo6q8u+vGgFejz0ucyaoWV
YQO86pnvwktk4h4EuDTQ2gpsgdCUXN3L6KTI1vFtkPYJZlBe+Jgt2yVNzOWOCBGJ
fNaEXbdJPg+dgbaaFAxqyTAENBb1SUJ4hdyUSJQT8G0Fe9YT32nJEbJz2Q4yK6Qu
LmkTlhg49y74NhoqhPLaSMb4fDFB676kmd/kiJX4PDz0gpfIdPEOgKQCslK+8f14
wntimghJVTjNO2nRAhmbe4UBNkbu1zKtaVKfbqlCaFl7jZDEYzH/egVH9lErNlNs
cL++JZ8ID3FkOCna9tPt59EWnfLMl0lOBD1T7MXIxiRGo4vnG66HTEvTEnDDYdnS
v37Jk35YV549jSFWK2Z46iMuKB3w8V6H9YDKeYTygnNaGUOke1dqnhmn0x2iZCOt
TPZQaR5noRs4eubnFFpLqpEJ6okvqtJZfwUStO7PeIrsKn0BAkxEniplS1mlGkv5
8i3OPxBdM3hQuIV5B5fXQQAZ9lAa+IRUB01YJMPNfQN8nOIQ44VI6nOnuH3jk+Xf
5uncXEh+jNwn/pRTs4hx+xan70GsswANQ4MvL7dwpwP5bg3HimOTtsFT+HNmEA2p
Tj+nHAPdNCGjSprpGh7QTTiM6mhK5/vdACfsgI7hvjlua1uFzBrYWVJU/YFaBjqn
Do6vLdopCAiv9sgfEWOc0M68uWjCwfzrHJBvMsuxCE06iMvZ/cE4LFT95WotZ36W
65XSRXEhdKm2CzTKDi5uHzyE1z+9Ib3VwbuOBLvPgbB2NX7Uzush0nYIcHxVIs29
7cjFFDx5dAQfRVSWnD40wmuKeDr7ZZVfxroa547Sc1Hz632yaw/xbBVtaG374dRp
Suoom3kwH8QDBk9+OV46TlxsHRflsJqAc5mkRHluryplLLBKGl0UmflTsADGB/FO
TZ2SxhJLmXcv4AwCTwB5+U7+cnwkyAVBoRED2s+UmKUmbkNZwrejB/8lYo9R3ag1
731FcPn/m9AjVoToPJRgPGtHKTsTkv7+p+Rqf4Bt411lYkwhZr4j2DweH87p+xye
bOcW+gBQVVfv/Ck/ACXJ4OwUoaI/qNT9eDinAE8jR/TSsrspx3lDJPTTmGFY40pR
H/wGjWRrFG3JZSwNGmQcR8n1X1MpRAW1CQG4E5W3Xgw45LbWiJdCItEP1iVznsQ4
7W5o5bTlg/ctpSTcDTbXtL0uBy3sQiVYphNmq7sXHHRBY/nevz+cbdRK6hNbg0WL
PR/EwupsSCqCPXd/S9XfWVZDv7IcZ9FhYGdwN6IpbS6Z54PhrXzDSWGSQyPoQxqr
8Tu0wUjT6L61WLgfPZIZNOQ8LXspCzZYVZpILRnvgqxB1+dRCxKE2UyPuoX6wHem
ao2Zh+PAxcR2SgdJ64rJxeVEhNId4Cq2a4fke7Awj+yzcXuQ4sD+9ev88DkiRqM7
7LgmJcmOsZUCjSEzCd1kzytTgFb6rPiwsHSYR5nAPprELb2q0pe88CHi74F9qrey
TIASJHE2gQuJup88UWiwy8ef5ncJyUhg5EcknmQRK1e4ZeK61gGMy0A/K4BMGi/n
AmYYYzJkUX3orfDIFmuOa+UIaTCsHX+HXC8rGmvSLWs2EsEUDZYz6/8vX7hqeThG
Omy3E74WLHYnu50e+WtlyIyiYmqEEr8VLLP6ZzVegy1AyMHOxw4Pu00MDPAFB5wy
yPJiuklAyqMHX1xswYrUzLUgNPShZ7+S+A0ge2z9SuH7kikdW7EM20BwgmOPhY06
4RSwMnD55QbSL5END8T/86zaA7HqwmfALRms9JZEYV+U4GfDbF0l/9qdupDaT0Vn
Kd9xBJ5OE4EIyzmmtte0Wx6P2kTA509uhOk2ltY9hBhhKzWE/Dooi9bN4iPAtTMo
hEG8Z5wqbKedrxotaW0PPfD7jH108e2dlItx5r0MfeDMGLs9+Sttyq+ijTdbvYSQ
PqVnNgbZ1B9caoI6J2LYhyc3HqURZtaFqdB5ZsGRufzCtY0kPfHAmW0VPuhPQmqh
7aIrJCciFbQdGTVptjQPUkCiRNH/8xnFWrSrueTdnj7gCpCSgcebpWkXcJVkSCSh
e0UtC8uYd4ic0aTbZaE44PrRL0hQKhtuDstY82SnUnFq09lXZT6a4fDi+wmI6tV1
RZF/qKfUsPm2OTPS1t8Avr5rou65y0EKZi7+RzXiFYibMM43wC5k+0cOfAx7guCG
ce5+za6Eb2Be/ltphkbmCa2Pxo9aczx3o0+U6tOoeKTgQUejrGUnNPgDHJMw0HL2
SIk7xO17/Z2kg2aKCF6Eyd1DYYZELukupTlGtEzh0jFw/ykX+vwROGxiAEpGVlSa
h8ETT+0F2odfnMFEfY9FFFjsyk/vFK1A5aIFbLNBUqHV2erWggdNogu1XS0gqBKX
eU3iF/SImns4Jur4onu3TBYzZVfysRFGyMJH1AqG+NfE+xopnVpKdQHyCg9VCuZS
2HUeMpsBOOhbOgO62XhHsBPYB7cu5TSkmxM/lgAbg1jgy6M/1Gkn7ByhhMqrQiHP
WdyPten0VlZrfITbV5d0L7St00sbpPgTjPFQt7ZvCrghp6uZbgzScq02Ygq43WqQ
MV4sTZQgkGfLQYR9b5PW0IP/rmC5c1fSnpnykyBYnXKmLU7NhsGhKiOT2ITA5P2f
el9Te5p+B2BzDCc0CDlJyCbNxORCBomv/GCMRNgD8WgAhFHa4kTJMZKWcOkRP/Ro
bbjJGGWK0lH+3yHedeYPb6IcXna3BmI6v1iCm7tnKxrGIj1OnNDZ2NmudbpL1wFW
M0A1iuMudjlZDMw+/bVhmw/Te7Jl0uRZRyQlhDcW8H1oiVWgYNkAjyYK9DH2CMYe
FpBzcjM800YyCQ3wbVpOaMOXhmnXtwJ4YlcfG+fXkxw7aVxzWJYahHmIOR/ZX4r+
61GeCQ8xB/CsZXJ3gvSq7q3KQiHzeJhT7/Nm6ZUYTSicoQRt+8Od1/WUXG6M5LiY
KqJMt79Ld31ScXJ3qsexJP2QuVE+3JmPi7yEA57ez8c38bEkqnzoVEO2rkqvWAyL
JtGABl2b4D5sDvKoUI4Hq7MYyjsSfzT4UGQDO/QoHkRSedG9WwLOZUTBIbF979Qc
wvVups0lQQ4kKOMhbVGtZS5l4uFNf0IaPdUILUHiEheZQgPNxajxNn+JzlEgmg3y
Sez4on4xpyKb85gyfLbMNp5/tNfETV2n9KCIrUS6vw/NC73BuGK+pMAqeO8t4Ne1
GcgtZvJR3nRDzLuAQGPHsbj8RI4gckvhLpA3kCrLNT2TDiJx/CTKcNaSQJacPxQo
bSYvWD3y7+VgeovJ4dD+2X9nTGGRFYMDQyFVxLfzD0X1VnwfZAQ4CGkRvJizOS/q
s1is29j+nSf6VAAm+ylQ3qJC6qaCLtD4H3pYUsjIReqqjk8R0J6TNuHHbv5iCPvE
x0of6WSTvvWPOEDZK7GOwQcI91J+F6gynnsRm5bglMQZITwyLO+bnau/ZJa/aWdw
fIcg8cLIRlDlJFgLhCIc7tG6X5O+IHWvNiTgCo5ur6KQCWMmvwfqznXg/H0P5Wu5
6TOjVdcMXIuK5XRM/eIOoxMopbQ9jxVQJjW3srTZE3lbD/LGouzjoyZUrrtxW0ef
GaP55K0IAr2lgFfYbty34hHYJewgxGcGNdClarB0E1Sj4tzYzIC/jENscHpHuF9v
BiZupnNHDTwcG45vfR/ZGqYXpVktKAegOQbGsImKwLEiKd5dWJ0n+7upW9mq8zWh
06v9wemYNrmeqt9boLIVQnBz+D2l5aopIHMTkAYCm63/FdTmZd4SVqWHdMsZf0Gd
BxL3krLGxmaBRc4x+DNWQ8gQjdU2tiGaCN+0QYz3nqHfhsHeoJyM31QQg+mJRxS8
XYK94xKJV12WEb6q6CBYXl6bvC5qgcip8FZCVCUOLYejGLRFm70nVrvq6ZJaKVS+
+PBUkHfHiq3Hl2x+N48VqHvcoKCsZ19qHbtggnD2aGJo/skPTyLOTr3GDlNvBi5s
2fBdZhZQwcSmwuYpUJFImyei9F8cq8HPclD49B9U2FauqJ/aXDwUhnM3Qbc1sBfz
6GGx1P1csOQmeLKAnSjOBjKx8dt9O0V4NOfeO2idtISRvvlc9g+cMm6wIRQ0hcBv
4SLjV/RNFYbmWRMmSyqKDxZuzC+am3Tu2Pi7aaxvAMvvY0cxqwPJSFnxEbKDvdRP
V+rHAKlRZRZ3dSZKx+cPWg8tbsxVkiLVYsfqL3/R0zFGr2CsH3PPes+iuoxlOjHF
d7Vj5OIDzr1Jm8prI1ilVRFCU6pjJOLUZtEyNkw8/Uh2ONXF7AaviaIbYYyJQfor
WCx7nZ4LspJoY1oz96x+umiT7+08988nxPAN1o5Pz7pDgdKDkqRb4Jiv/rYdm/mp
hZd+S+xxReASAkZzIibxUVa0ydYNgiUOHQLKFI1u5+LohFwZHq8QvIcmPkDAvtXj
8fxf2f1dGZ+jN4U0rcPHGXS0PvPJOJY8eeWW5XkPBAa2MR6OeF0lDxI8NBLlgHXH
V9EWp4mXXNvyGbC0PGlie2uoPb2Xt0duEpFecUE/5bO1pAddqAUihLFnr6w70Tlu
DjTKPTh5uXacwOC8Pq7UtcA/zFtICozCp4HD9EPQJGX39Z5cVBGFRK7HFFc57neP
7K46gxXuFRwN+SNA/Q3s/nvEVKmpoZT35MVxMpRFwnIc4ut0HuxsXmE6rohXpeqy
SfInWsTLajP+Vjo7pJ3Rv6F6nMEjHBrK5dhM7xr5wwv7k5UjZYyplwJY6tI+AXQa
KVMyjGriKcjyNIK8E2eQ18II8lezrLsHMs+o08NDcObqVDKBOmU9/btuKau3HlFc
fQJ9zodoCXbWy0arB3ZgTBMdrYLzVkFYK3lbvfQUsi99V4TbiFXFFgu8MEBLfmai
TfY2bY2wji12BVLSIQ5CgkCDtyJiTCgWEMjT5gej47e+yHZ7faMtE+2XrTk/WPhT
HPidB+k1A0ey4VzVZJO7ZoagMU6VyAqAYTsJ9sDQOWc5vJ//dULzFSrg49YvdT8Z
2JbvXLpoBSLpBrS+SA9zzqBALO4/n1Sn2ublQ2XkQOEoT7KcVZZV6Wkmo94RkzVP
WpUphuiGF6pszyE2Sbx9C52KXdQ5c+PIElk3G5ymbSR6buEkWiwvA0n0rLLy3w3O
Vcn7Be4SnaITOXOLwjtjH4VRC5iUqo91atTnBCp/ivm1HVSQiFym7WrZjtSp/kPw
TA4OnVe2pSSoFdyXplk0oXhGNOjyGhZeZuiElPoq9TfMevnXay/Vwy7FRMAVOVrm
evVwV5F2kHtBiV2M4SSf+WLp4qAzNJpXSqPGWbsxJso+Be32PhE2nM1jPOWm0AJh
cX6+P/MWH55AzGU353c8tZCYvS5vuFCePR5eoFyTqXFwI455bq8bUMuBjsLmw+fn
iipXgjiPT+4XdWh4Ad235/E4nHsNrbWc8SikBMt3ytapLvULofvaP4FLHG6SpNe2
HgTn4ahhRaUkGziq28lBSJM214gD2JUJb5VrD0To4z6ppDxKT/p2oLt2wlmgz0pb
7JjxUT880K3sHMdXovznGL2aNZAyoRsp05Cwiu1EgTlkbDHur5UqMmftpyWqGx+e
nYNNgsdCJQJwzG8iIlZyOODGs14n8ZIkMb7phkhgwKRaq0WfKbvSlAEm5zhiII4L
QmWWM0oR6O6JhTDzpkpSu7Yq5DySWYgzaepfLuitjgYRUkFN1rv4uV5IjYKYgfz6
o+WTOBp2Jva3fhakfKFpU8Yvn6OFDglWVSjCIBkUKgG+Glj0y/ggRiozBK3uQPRq
MLoM+zfEZK845t67I9D5jZK9dD/iIsnsbsLX0pNshknu9wOR7SqoL02VqEpQfMXQ
lSsNtiqu+IMvvPb8zAGbxdXVp3UZfTNKVar/SYtONwTG73/GVwoG1qWEvQ9qr3bM
jDzfnyDVvf7kf4qu1JsaCO064YSw8W4H6gOuIZgBzhjZMrIPOIKCQht4tMWC8FuA
7yydX/ltwN30g80tqe7R6ZK1ELTWv5uCxw8Nk8uny5OlKVOHbyavvhYzuEMnbe9x
Z5jkjYKTcXrW0GP527RzamHW3rqcquizZPK5SFXPM5NEadH1Fnm5/5E1ti+5nxyl
yvmYweVPvhlTR57zs/rZ7gJk9VOx4nAToCBKK6MBQVzIqc+QkmNEYunfm+HlqvOW
MGpD4zed2pqqoXgBbGx48oK3hDDNob3CyVdQLaX42oBJG4hU4TmauRDVr05ejd9U
DDJqqazhWOxiFTLxen69Ii3XdPJXdHjPSHbEvztHqp3SnevMKoa+zsZLUIAcasci
VvzuZjtYQuSvX44jnbabEdUe94sIil/jFqmTUYHFDhbo4mtEDQnniDdrhNkmncGx
AlMEUuB3GROatQD0Mu3YF+LED3BXvH19toesbP38bjURMxr2wT5T47HW1ZFnA0Hx
n2k1WkDxP8HJj1D/f24PKwTvwkObHIQkkPdiQRboFDx4Ed9bYXcNF9it1Mv1Mmf8
8oeWd/DOCgRQ52RmBBE8G4hBwVLmyAKayWCbPeqqik9rCmuESakxo0I+RguRxZMM
AR23uJnyc6vtGlO3eEe6/IUZUvXStDZh5wfmmR44Ohg0DmTHO8jalcfE/HZ7WmXm
54O+oJ3rdQUTWC1g4RRGE8JBHU6YqIUMRB/nlVrox9OiYvi13PPzFueH+t7b4SWt
Kymw5qYZ1lgaxXZaxRamu6nH6zjdi+fc6glGKHV3yDGRmMgJSPujJvW7n+68noK1
pvVGLTbyMw6aM5ZxicyqgAHMu7OXSPLMCX67k4EWopaNmmDWZMeeievgtIt1gCyy
bf7dIItr+MDW3JK0DUxTRgdOuT6ULIdLfABZRrWJSawYxUXOdeqz4rLHC2zfToIB
TDG8by1VG/lLfe7PtJKt8XKoE55QyC1L9diKcUM+oK3lAjamaraY8/5hvJER3Wqu
wi4tt4P+PqmLX2/S1pd0TeC9aOMKcMt3gkn9o/yfzciYVq5lgaOvFXKgvFl1V0SX
J8RqDL6gmYDkUWp9pVPM7Ku8J8zH452b4uPC5PqkcdYfNQk1BC3CurwGvwLT51I2
N4XGSzX6aVpL55uY7qH6LriDWFEb8H2bXZGQ4t6CNo86ciAJc9LFqFG76lxCc5kD
bhcS8WW5F4SNs/DMCy7/ikjSoO9wGVr9IMB0KyD3JAnSm6lkHkGjsKEI5RZjSzeU
fjV1LzaAixbTxcwp2S9tCh0rdThvSPuynfsP54wNeRoW+/th5oR27hQzLrTmbxnQ
V6bR65mRuWlZlvk7uRoQzIorU+8O6R7YboVhTylsPlwvlK8Ds/+jgb4TEO+BQnAJ
TSuU/Ry9B7jfwMxhIQPuiZJ67ZjU+6YVjqnSkFNcx0u1yHLO8dGi7WVi0rB9/+i+
wuYz2N25zn7WcSRa5+g5GbKLaAgigUIz3M9X9F8VbclJSmP3WsjWRdxdSLWyxBV/
LADdSd0Kq7aIACZFc14br7GyfLDSAT/K0iPf/TRhSySACoENKvmD0MEojIqB27W6
1UeQkc8A877FiExydgOwCt13/n0XcO55bC5qsFsoXvn4YWfAHaVJMVcJeew1rIps
EW+h1BZCHERpNgWsC4mTnoLHwnQauUJTU8Ln90vIBeFUDoqbeORGDGEvOzJr9396
otNl0z4GTndpCMWb6Fbif+hHseG4HOc4uOnPMh1/vXAT2V0Y5DxG6gX7ke95WPjH
ADMwj88ff/lQGYB4R1uXJ14IbFnusL8cBTesV3xLSARvCVwrafUQq1QcZvdEOgZ9
M4TPZl5ESUm9Y9GhkVcvV+xztb0D+Tk0eqPFod6iGA7xCjBejM5pbQBKfsvm8M5Z
q9cE5QWfk02SyL7PDBHqBuEYsNTETU/Vcs6UfgU3RbtNHHOWk1rRVcmyoKUfHb3/
HqBMJrbocM8Ueu0s3RIKfacl8BpmbENhAuOQbNUJ18P2PffgbOq/t/4sABhD4SgL
/pUQaJ8tAnLXZJ9rwQW/DYwG8zLEGZq5AAOqFi9D5HzwzrAQzHYiGv3cX0uM0hG0
9097VD4QZHntq+8c4DTeCTnSTEqEKGmRjLLuPfp5C6JnJxJXCjOgUdkD+XOy+K29
4qB19qSJcZIHp4DiP91fTEOC/UTI5iuiMx4Y3gDSNbJaS8Z0wm+hFpaxNNwiwGgi
T0YWDl6xlRK/LNiQal13exWKhoY9zL9ON93o72fPBjKekJzk7pGBZLmPWWni8pr9
M+1HEQi6ErLeZhTdHN+MSr7snnCV4b8ExE1Re3+3TTPmrYAcsxtYrm9S2uS4p4Hc
NxvJFTmMzcG0wMF8tId2egI4QKPICg8m3PQtkLJr6k1G8h25/E6acgwAnddsV0l0
V09V3KCh0cf6wPD5s+sh/vDD4iY8RZUg/Lf7bhtSXPPwOGYNa6TNtr8dtIfF98+o
ik+48sjVshTnLY8S0FKSJY79pZc3BCupOUTAWhApI5K4kBMnswz77I7+G3Jl5Y/G
OI+MfVjaG1HZofd6vgYYKas/nCzdviraMWUzDCfTZwIwYNowQ17vm9WviZW3Q5Gt
kEmQeBZYFUERMGjUTK0L5GW30nTPzPrYq76Ke8Zav483rVVJi9C07+J7GT++E/y+
b279YQhznHOwRGdm/4vfxZOOmDpR9Ejn8qi+zSZxP2RJPwu54tLH+KymWWfTLZeS
AqrMk4FXI3RZCiEYabxLoq+DLbGyElKL7q8qd9kpvtivVSVwW/434iCzl+IcVsjA
vHznliH9wvVaAK/yj8VVaSaDK+ralifhU9eN9vnM8gz4kVf8/Zzeyy42WrvCdM/l
Xq0oNcHu/bLWkadYxYJ0FBFl2H/cjCgnQT+e8Pm6sSSz9tDrref6H8tU9+AYO+J+
Lcm/5oTj0ug0PG1+/TO55v/XabT/N+qvzeBV8fwGMlsuomklEErHM2Xx2Luj1ItG
C/WGKug6S4LVXCNKO6X2/JCXM0n0xEJ7FaBsoo5u4z/Q8RyV3aPyY7B3hZWsCL0n
15bkeSzQnV181PRc4wj3JVvlz0uWKgGO10QujOgP6YZ1y15f7KLt/7ttiB9bVyII
4pyW4QHfALpfP5IXlekd4BdpAeTkhYWb4gbqlXEhj1gYeKpe94ktccsoDfQm4Erp
h/RHxQ4QPbSGmxFwJry1U7ZWi3fhhO9sk0L8y4h2ocKJyec7BE8IAtnDSwJq/02Y
5Gi2n7mPETltPoBJDcHuZTnNrXrDoqHmXeZBk7h8djYtcJFamN6LA7PDCM6mPVzn
6UfbHr331rBlP79N2LkakyTzVTEqtAsM9gsZ1DTXdhgk4KitjFs6EKWEdRUgwAIK
BHXjKbB/8mPPcTSSH6o8g87/e94hUb1tBJPzVonBshI3y+7x3QwVvyc0FM5vzNj0
NSMoIGDDZtuyUn6SeVHgDjQgnedATyArxHf3dNsxSL4RNKjz4OEwa6LxzKquGQok
Mcgzn41gOX9qzSxz5dKK5s1cizFreiOgMQKre80Gp8ILRnav/Mz5K0iMLONpTGXT
yuRWB5+gzVjmjzzCji5JC2aytXItP0JCRblkKKANwtsX7lPGIV4Nwhg0o5ygbex3
ZGZIyKIzf9DsyigTinTAB+koOZiUEM8F16S98NLmos3Jpl+BzlA4o61bh0QBcbdo
Ssnf2m2/+vWa3ypTLREKaUG3bIM5VJY6fbK9E6z+faSKATEQVfLS5D0XGu9n8POL
n8FDlKeNZicby8Idw+/uvkyjJUa+QxLGtNKdI7df9mGnlwfF/MV+ucWMUO+6RNox
BcFxdVpGVyhuglIEBo5mZg/HA9zO7VAZFfCglyEw8mOnep8R++gvYqqqPBvuMGhi
7M7KF6DMYsnMXv/kuInVBOdbgnqxVHW7RJve3mNPKBI+e4wN25XPt/p5jEZUcFNJ
bwHoRUKqm/g7ZfpLioOMZJHhw3Cn6lD/Nt3zpCgc/vhmKWMm9qjexgfd7eElQCKH
P+Ks7mL685K8VbundH6q1bLrhKlHcSceOcfpojQFeZTdMiySxYofuJjtmjyJjtzm
LK/590kglYHt0xH70JU82U+Ko2VwnaA41g57eg1NNcMxl3U5CNfREkb0lBOU9Tn6
h5AON8xaDVlkYQa+hRXMEZV+dEoaYM7B4k189EYUMuKWsSj6EtSf2hV6puYhWm72
Xp15ztoPgvJAbu3SgCeYschjx/Z26svSibHKL99Vvkzeyysh8OeeiXEgXNmKDYXU
IrRpK6UYD7kooWkkOrcaR0340c8BKE4gDVpHUDPvn1CisL6ZoRy9eGhzNjuLTyBR
200BF6YvRKvstorX5/tuhGeehiWBG0TD9nuMZd/As6Of7H1xRXGvMcVwbpX/+hq9
sO+tBUu8Y31H/RkOUnwAIdPClm1hZV8vPw2vyBpD9+DOudDY9gvswPFbjoUKEGDs
JMhsYaUAzmnTLZKRhbH95pGFRhx4i5XqQ+eZPjUvdBilXg76SKNq+YAxYIe7Tr9Z
R2ddBF24e8xBdUOY+7TJuOLpEWKpe5byT65vHKIjN5B84phFyaiUSwS55LkCP9v5
k09vqqd6WQOlvnNg6AWyypZTGCj8W7BE9y1k6CICPN8LzS9EhBw6/sWIoXOQCjSx
7szskYALB3eWmwOL301Z+fQjgCo4biFFhZqZfPLM1usDv4V2bCGp3/lFMYhjvvIV
bwYEY0uPxGkYFH3LAc1IBcoW3oTvmTMWVjutPi7JVnysivbcSPYZEL2kGwkDbviT
I8JVoO0Yma+tY/ZQim0Jf7XNgyDvgIhWNpTH0xXQtPkAyIWBrnrJMCCiiqXAcV1H
5GxL+b82hNIFeyYqPa0WnA/Uulgg8ql+l6USY9xjTdc96NGVBXSWKUFBktIcg9Gp
Ty83y8dWwW8iKDI+tYXWeEEuzzmay5DrOeX8giiv04EXmUDVg4ekqT8X/6j0l9RM
q1v2iDrWdGbVbM8EqoxCraDG7DGoeeC5uvqP5Rlc1wHUCphOeTkcEjylRb3Krnd3
cFGO0yvCc+IINtccP6UCq4Elc9ILxEL9HzuPSp2pr/wEIQ8qCQSjeM7W7Fu6Diiv
I45zNI1Thpa7KNI4Pftl2eqT5fSI79VcmzcqCZIFeN8OvSLDlYq9hoUZ6R6sCnHm
emgGc4fr80JR821ihUE97peo+MQPbQpa5RfE79/A95gOy1Ws72qkwkT6yaEhfNLs
AHupBFjBS2HFvck8fqiNFlMQzBpNS2H5ItBNW2+70PQPdktYpHw/GrNDFHz5TxuS
FDL1wNNyhcUmuUVn8a+a+LIFAuyH2GXqiDrifzaggheqPTxolUEN7tUQXqNjV3qt
SOS2kbn9S9jBY9xL4/As1vrm/p5tm/arid+zUzMBA0Z9IW3DApTGHA43GV5MEyhS
o9hkrD2kYKuB1MTklfb1is+AJ6WOUBRXm2YIvtUJsBdKzFfGvf93Bjs8usQZ/nQq
40IWH5pYmx5EFPY4EGT82aYONtBMJ7lefWwgyvTEIxcgI1cjSBLSxu/wvYK+Tm0R
m9H/FbCyeOAdzMo6IDaczRlkR9SF+s5SymhcEcgJff9PmmB56x4S5NZ5lNN4Rg/w
okhDtfUxCWIdvFTa4kZZt72gzwSpcV1C0PeeqHB/YpdhBlgDin6Dn24KmOlwWhxM
9X0ykpgjPIo0d+/Rl1rO/whnAt6kRakbw1YvLWw0OS2HiKEWFCDOtn+25p30W85g
LHHSqCIFQhCmTr/623x8O2tJ+2faNQsc+N3Zo2qtUAZZOKHlAkfn104uzI4w93Xg
NNDRAVlJ1sT9CrXUIkeZ1zArvDq1UQpw9a2SP1IkFP+3yBMbdxcybCvr0CyvHey9
bJ2GpXr91Be9A0sW9nqadlOONW9GvcJ2sNjjBTgCvHgvznV3oZwBIuJ05GxgEDic
qtfZaLCDup/53gEv7qswtsJM0114up8LJJMPTOyeqyqFkCYqEKeHYtZ3vX0H1HDj
IJ1//KGBzt7oumNk0GBmSuaAao/f/+I0RNMdCggO2UG6ZQRr/DD02C1ST6S5bVJe
cxjkb2nqwRmbaDQQRLBfMaoBQLLvvWnpJ51UMJ8QrJuVzOHnpt6CmEZQYDGa5+3l
NSxPyW9n+FuzuL6BYEoZ7ig0Uwby3MlhVNkKiJ/2eTbAe4/d3WzdfWSy4vVURyCM
bm5SqgPDEnwXEjfh15daC/sEJ4s4p3mKqQsKNGHlmJDr906qYOqMJDNxy2sJ32Ka
Hzb2e4i5bxvqW9mq8qcPrgmcTrCZNh0dLWONncVIqZfI8Dy47ieABRatcYR3I+e5
LJW36FGrSoLBWuNDdCsDZdCl49fDVPJCOS1bZQohYcufxrvQ0qWcmrBARecD1lSr
Y+7xFSYfb/iqKTkAUdtd1uPpMbJau1+fR0PRoo+cJiMzCTq2Mu/RBn4HK03KuYAs
34mCqryENPzW6n58XUbn8bFOLlc8IyF7hOVA1zQIdpyXqJXVTfhr2NnPgQRJ9qol
fP9wvri3n4u10b/oov5oBFGVeitX7i8q4H1ewIXjMsu+FbxX7MZoID9rgFQzobIO
0WXE15eUJYYXAZAv435VYu4YMwqhxli0xYPANKG/WXLzrvfaEUMzPa6ntGuJWxeH
/kG6uSx7bDDPNa3zPK6teuZPYMQInKfQ9Y8xdOij9GD2G46elYGw3Gk14VOYKsqd
nWS1UgRJRFRewjwoGevBBxN5ud5cspl21lVs8SsvNZgxzgSVh3dpX2BIp1OMytVf
YiEZmBpL7l7cJuRf6WBtqw8j1tuhMvwF6BGlykVLX7z6U4rpsH2r7FpIvTkJh6yu
ts38FSvqa3JyyqNtO/9Hvt0fdP+jj6GviXAYrdRJo1Q9iQW7fyx9FiDge9tph/5X
shRyxrlSq9Mwzn4cUlrjdhgvXVl2FuSV+87PhLiO8UXSKOLZp93mYRPUk3Zwtj/6
hufaMbBRd8LmH5LEXyetsuQbF6rKf00EBQwB8yWhBw+p9EAthsn+MU/t6J6TgeII
wqzBMbm0qoLZWbDI6hY6NLPRK8GTK6P3mqCR+Hi76GQvOEBd0J3jxCY717rpI4Vz
miQ69WHE7m9ZAVDwQpygZ3v9UnK8sOEW6bO30lIhPDg8wFt/2YPgHa9Uh5FDLFCj
Q5ukxRpfHENunckaYIaF5d0TnSTjxU/JvIbXRWXvshz0CMVRmB4NH4jL0l1vn70M
LXvuPNEw8yWdo4zGFAiMhDxt1WD/ppa/w1hYhKzuwgayP3dswNRpIrHnbJ1eVvrv
anVB6YJluWufYNizBMl8e+BHOZzf8kvfBlQRtJiTcatEwTmxNdz9KVl38EutUeI6
y/R5oAP/2glMMiWGIrN1LP+/C4bmpgqyz6RR1VZpgMSN0AGF2kaq1JsEoLKVOWLd
s97KR4TChc4pK0Dm2MC3o1C67wF4+phdoxM+Ns/bqO0x4gf9MygdsF3h2SO2Ms7f
9CeD3o5kADcezjcldkQbQwUPooxEXUS117nfruEgbNiNibQ5b91XIf5LsB9/OJQe
Geg4q0EO9g2rktG8etclA/tP08uSBiShsJasf2cOwWW1sGpraKukuSdKn0F1N/c7
msu0HnjQjUWQQt7WUrbXrz2SMthk6j6skIKN1Dqfya475dN/A4seMV1GagX8e0oI
v5/h/ZpYfnKBFIyQv9FOzKTVWHKMPCXljN1cmdNpsGjDNciQ0qQPOySqqGWhq0um
B4BICqor48DQ5fFLuCjvaVmscB0d40DdepOiIWByeaFe+fVPFhUnmqro9zOgL5Vi
6HSOVGrBbqy5kV5Rgia3lMgSV7Uu5Z7qXvduse9oS/0tD9/cx8rFEkS548jieTMK
/3cTs9PilETbpOet7611//rycLUXU1kEo2fqAeXzrEMU3ZFbG/Wawmzud6EVtAXK
VmO+ivZUsFhzmUJTIiYjydLP732URCn3cYbKi2836lCsH266FWhsfdjpsqCiTmVf
9LwwT4JVsUxzpH7WR0QD+mdh1+QQmskdba+Cr2O8xzGcVth3rrDQYqxy7PxxD45w
s45Vm9ajhPGXNRd+XwEhWcHrRdO8WyT8GswlrXRRBKmKTaDojp1Rus9r0z38jyA9
vtfqd0W9vjSt5pDa0NWG7CQuE2EF5GfE7fI/ls9Ph8BPxcpW+Bo32qMYy9cz7q8d
+BladnA4V5pLbfpRvetW/eT5qM9pX/kBQxgOERtzGSETrJNvQZEo2+z9Xg0ulAtr
cDDgWnAbiX9g55CkANjU9qiZOoaqfvLnAcScqvV27XXJ+uB9kpkn94HeTUSNG4yA
AIhGsDQZ6pxfJdGBV9cfs5rsadkXb6MRWKqXYLJ5U9avJdRyoW7dnDjYjKVzZKZh
f0dEFuPG6kgyTukdjTMxNcoYj00E0qT3jNgA6TKUMwMe36LXdR35xYRqCLM/GH/y
hFiU779tOSOEzl8Tcbr8N7fXqg+D2jqroKZSFjLwXra6LQUQyoFPe9wMWBrVsa+e
/liFhVxWPFVI1+dFnZn+Gtqe8hT9iaExTFWK64xD5o+quiMkAZtGlbsa8hQ+Gym0
QvKcDluJuYrjWI+1xzFtJ6rrnVzL4oteh+3rKbUSN/BR4a2PkIog5+gyZ3JkijIv
KtaAxeb7U67IYqn4Dhqc45yHthCx788H2xWfKirVS7Q01JnEgqVjCfM1zMRbOhVF
H0+BVovgzSM7qnxY4ZSbr1jitdXeIqIQPQntPmfLWyG+KSy04G3BHAScdqrW/1vF
tza6vrO1H3gqYyv7C5W0Irm3J4H3Qfp4yLVIllu+wTK7JnhopGZvPSQcYByB08g1
fVo3WpKP0MG45lVPTc0UP52AGy8fCQmWUeRmo4SzSRmve5JB4QIpwxGOF9PEmv3b
PTzAjQaMzsVptA5JfMzvsDRG2yKflAH+ymw3myP8hbVZ+QOXy3WXotvIzWoUlT/e
pefTvmeM6uNFtrS5KLHLIxcLxyaEoxNMafLjjcnWuDZ6LQfhtWlDEbGr79pVyA9G
cnnRqdJiqE/3D+qxRLA5JOgELMHGOBBTHP8keGpiQNlOV7+FRZMlMs2XXsDnzBoC
fQynJfa/Kgy/k17o0wTgViLjM+h9Px1KWccHucJXf+RhyUOY1m48ULRmOMFvNwTD
lQ5N1jtuydTot+6C5Chh+L9O8sfwg2k6ax1G3qtOS3DrOoUx7WBi2bnMcGhC6AiQ
IRFrC5AKX2E1w/DxCf3PEXZSBLhSLGVsxB0jcPNe+Ip2f8VEx92eWKrWHEVvuvTe
Pvenf1yV+dmAyymuZpSjse7LlbwEWBcmwNCeLCZeTpORhV4vOVSlGUkvGQ5vY2Mj
4+t+A++7cTO7GIiJPJthVTIUfavyyKvq09+U3yHqLYuSsgloxBaoQs9EMux1qI+y
x/gE9sysyWwVLa9Y+EncgTPZkkiypUFllOE1sA4vSXFFbqgL4k0Cse6wtnz3w37X
99rIDQMFUv8R+J0mvEs+iDqE0OgMLfpYr8+MhW6BweInj6c3WL6pP7rqyFiV4azM
eh7NX3GF/YLATQUTuqwBlqfKRNJErQMsqxGqxgA2YVBkntYfk0jRx2lz/YKiFKC8
kCQgvfgp5UmuCS44odS4oOKW80YrT+I1BqosUEnbdZed+VfmXZOQKVfvkMA0T0ph
Afyry60qNBWWztYoz4fTkc8nBal38K12bOhyDrfYP09qV4TKjO+IuVLNoiHuXJef
kvzTh9rfHNo33+0zO/scnPGp3IDKXsJqKSdxNg5tT/Ui1DdNLg6r7iSzPxLdPTUp
xvf5NiteotnkoHpRmPhYAlB+svV/SZETbajaQ3UjFW9a0kL3uABIh+XydOnAZF1b
MzbVBj4XdzYd64dTUt02o65viUY61UAIvKUa1q0nOu+Lt9Hx0zoWaPEwiIGaAir9
5buqL6jGRKulSeqmVKmVZA3xl7BipZxb7ODE9NopJEBYSK2sGF2mtmllTE324tcU
QST6TtfgGj38w/ndY6TTx9wc5v3AKGQd/08Iw7M2TrMeGasDTXy+s2+p4PCyJM1a
REPcqasEjbdo5q7XnRH3juDmUtm2xDCOWW0ZIVZh90wEeFVs46OitNSMtCbZKj5/
qOgXpKdKc1HmA4ap+Lg11T9z5p7qSObylnJAWWY0KnhSrlC2t022R/jHSrhysebN
lQNGpUdB5zO4dadyETnid4V3KadCtxl3h78/Y7xla8cZgWMjSe6MguGHOEIFwTad
rDnEgYYg5MSkR9W26XPrGbVsiwZggDAtjD3mGZKPA11PzBtcQFAUcGaKtRKUhLmX
hxftSb/lgrBRJ9faNqqRYnaaWr6eyd2D1CoItOQQv8tlb5Q7TC6zl43/Due322PR
4m42HzqqiuTzSQz0ppPxLZ+j8eJrDHL4JcVpeeM3+CvABxVoMfFO0yTSVXuUzfNI
PkiMlzKyGxJmvNIYKd496q+xyXu3N6IXzmk8MIcpbFAxP5KFIeEZ4CFc9O9RdFhq
E7AaoO98LOxKS6Cef9iEfnFl4HwaPKGqclueIaUpos8bCtcghrfXC/MvSQIbT/qq
6dZ+wN2gy07RLgYxhq45YkLoYeQhBxEYKJb2hfx7BJk6NRzv63iASs5QBPGxzwPU
naBa60Vma92QDpUvP12M07Kk5XbuAWW71s/mTiK9BAPIXbgRLlt7Gs5UT+MfsSBb
qdJX2eIr3RNhyA5Gs6aBQ/82BQC6SO7KgmRsi20LVJrJkgT/HPeVY3ZJSwC44hLi
lk1oszIDHHo0VlyqY6LrKm4L5k5rfPfD87Kz+HgJrP+s+362+aFY1H8aXU8b6/Ch
B9uQjnDcDQ4rCBmoSrJ+oQYqsdbi4l4EpOuxM/csCeaja9DjS6KFRvzqizvJdsJW
1wb4HbRgWOpAyFqkeyqJS0guRpZh7p/4B4fJqgs/c9iFNX7zOQY1einrmzsnGKwk
Ja47iXgtw0eotmHlMot5La9DigR1Wpb3fyV+OvmjiIk6zWUtefz9M9fa9JE0fTA4
in9L1apdaBv5qkBh5UTn8SYK5aOBduIPPlMq0ncMxvPftPz+yM9drSo9cQ6qhSYp
cgb7kkfngRvdHvVBd4PWmgNjGKBMglwLPHe4lGn9rzp8GJ4p+CNDiu7qb7nETElH
K0ja+Mi3036G39rzJOa4Yt1VNlZjrLsvOGsoa5f9bZbFI6RkL5otz+9Uswj0bMDy
OtzkIuesWMD9T2nc/N+hwifMGkJfWIcuyqvxz3rITGMW17Uwgn81WZOYkJZPmgKV
w08NrYsq8NhBp+rkptP5bR58DhpbE8mG3GheoWBwYX57MzG6OFGZ28byX003TTHV
y93JqiGMKYUo4XGGvSb9KLxY9mfJR9EHZlFiMfMlOdnKDPtqZ/ujcJKaj5UpzuJf
QFQMb2IzZm3UlPRd3qVzuaM6azUlMwLWLuehQSKE7b5e0FCl/b2JM7ii7PdiSRLZ
YJcwb3yeqdjKQyL1iDTytgpRFv0KZglaWcGHT5wqx59bH5HpN37gw/Ts7XCw0pxy
t3jBtOG8jVJjwca9y/NEYP3e6di9Uq7pwchpQsgzgPQneImqMQdPfVTTfR69bC0v
EdLqeY63UntucA40Cgnl2KRtvmYdNvkKUclGUghdFCffnChMZeBDqllS7g6vzROF
SHtkffigFMw1y0YeFFa7CZ4pKz5AtBnOhRiNev9U7HLhcw3EcT/Jc1BTa4A9jxKU
gowGx7VV/crb0epIk3xL+f6r1H80xkD+x3kh3QVxtOzkrf/mV0zVdBpP5KHet31K
1P3JezcQyzkuxuK72SqXykb06PWsuQijy5YPYhK4W1Bdd9W0lL+f7ifDoDeNd7bb
On4Ay+L6cSDEI1h696U5SM/AEadODsUEXgjl/tThxSgcdRnYgaQX/bO2+g5qMIwF
1+TJqnNjj4kNTB5/YyHgAPPEz20Y+HKwSPa9O3iyHkLtm5Vq9waItieAthGwGXWI
LXKCE/fXHSrqVJswW05fgW35TQcg1TmZgT/INgkVhIoPFfSluhBez520c2FhRwPh
26sLtn7nB7C5FCA8m4ID1PF6iLmzvEbv7oxwupgbkOHTRwoKRkllsfiBnzblgZdk
Mt7vSmQgyfKlh1qKCgAcydaUuXJsDFnGdzCYoxSVd6ZRIXDMjU827LnG+a4H3UvA
7QD7aK5/Ny9KtNaueFhpWAY7BGnlQtWTKrN4z4uFEuBEf2CMp00jvXB8stFIJGNb
BMwfpFdgn/iA3IBJN24CZJDZdtn+xN7iI9tsvl5epp3aqAxJ2PDVkMHNaXrIsKZS
lLbAnquUvz/R3hNW3kyp8FYJY2gljO2bAIs2W7y1ghPa4KA9P6C9iT6aXxwDHpco
kXY5I4GhTAO60jblqbR+kUsPfn7kCZCClx1p185pAiDArwwk3e+hmQwaScHIvxX7
fTS+1a7Ldj9/I7MgPDsDYLGT9ln2jr6AikmBej7I9i9s/nc+LKkGp01qTznGfg6v
9GVdrhUKX5J7067ghnRwOkWb7ik/Sqq3DLmkgLSGNOJ/DCq+F+ls7uyEobVOIKM0
GciwCIXknWx0tp7jFP96ILnABVbBXQu90Sv/lnJDEAJ6BULiTlhjl9ueXyPOcFuP
oNF97QAbrfsd3O2WoEbRroI8BqsnV+PgUzgU+1/6PdW8iFy88KX5dRc1bCNnOGZd
wsBkW3fVOmY9cagJ21FeRL/xAJfpYgmzE0L2XiYD3N6t69b6yQPfc9HwW7Vlx68x
+3pObrCgkMNr/L4K5ln85G9medkgtdFBD/h/snUKo1MALItzFOrVwwysmRPP0UOi
+DZb6zG/SzUdF/jRWz6EQCT7XyBdmdRcLH8GJG2kKpQqIHRuxTMRyMccPTJ+rY5q
TNoq4uXW7gvT7yTcuTpBRVIrHTTn4OvcxSrNxRcAAJLxxU4EGtMCsGpZtzVnVJKD
Wy8lfaxQIbohHbh7IfGcpcF2qGmszPlw68F4GWdl9pHU9iDYd2knbdVdmqcDcORD
ao+MGP7Gf3FeS2L2euw7sHotI+P+WbmS86L0WbTM5qXvLOjlR1wXFHNbkfyEdTAV
IrnbaJ2z/0NZ1zzQPKxBoXcYde77FYHuObx0Sl9+5NR3eKr8U2uD8tv0M57qj0Wj
sxJ0FGwNxnFY/zSxISc+dM07/jezG3SL1vPnTXtC4O2TG8i34pvWsBvIydhzWsV3
mIauaKwWvQGJId/i1e+9N+EFoT+TUTRVo943qmHsm6E2H9fKDibQGfOkPl3FGqXE
7jugfQXXGarHqvMV1wM71iswRs1gT5KhVx//mr0yJM+6b+xa30xKqxRgL3e1P6ev
N/6FrDwit5blBD6P7DMUalIL22PTH3GW7Zk/ruIK0HsA2MEyvfGoXAfkKXf9+qjU
3G9MPTpYFl4S3Sz6jwSELCaqIAcHENomfqXAbqyY6sAkuEh9Mc2lBpGnVY5UyzZv
VfRQbpBv5zAytL1rmAz6w3iOxRZJt/Z5XRsFpjwumj9F8iZsh8FA4Faf7bPXOl45
XDF/6844bIBh1eCf5K5ANKnwlFxD8fW+3vBArJPCoJyisGzsnNHymu+nOn9prBB6
meKFChIQWyiB6o8jdfESx53i1YbNaHmC66aoyREBylFYX1ZbqvJoMajXgFWQ4nO4
aywTMmGRJtA4kdKI3rhQf/M6LWf0hbeCRZCDF/DZkjRlwVh9cI4jIbNEiP1C18Py
4/yiZDXCJEonMQNAevkKS9dJaCjIoNq4XG0qpPVAFHTKu1TS+HV0DEVLraG2VqNt
eTlCxYFgdH4huk2WmLn8lqUyeZvzcwwfXwW623GJlDUk35bTW8ITgw7aYNZ8E9f+
rKkbDKMg39Rn2WPNMiDn6Is/k2qXSgnfv78eb/kWHclsdDNGkFjwS3LtYdYPd8zj
T4ni18S5gCWqfc/qGXKfOMjRCizyk7pDhed5yK6zl8cSQridWy1WcENN06ds5o4b
ArmEG6dZawyTkZ4F2o8hTw1GaHpMIRGdEtuTN7PfO0kJTnwzfs8nqGf5isP8TaLf
+iELSKRC8d7xD63isukWruwB+You88+iPI7D271OadpHMaHqmoBkRhvC3zjyTwD+
Q42+va7XCn9HFh7B74Pk47Ye1DL5VgVXFwmJ18rcMQGXkOOb4uX1R2fR77U+fOpj
wYkbdNDQeyzI35URxPaEGKg5bLLIxdiazXq1U8P60FgtpoUET0i2BEN4IcwmHOAm
MNIT7NLUArBGnlBsoIFBVOBI9FlbJp2vPyqloAc+fihmXWAStepEYyzptikeBg6C
+9ItHVnULK3v4iX/xbOQn8gTIh9tO0sIC6hL+mW06F59NGAhSmYOp99FjNI6ykfN
/neJAyqdlBo/MSKQqLodLMO2teJq6RURg2zYVFeihqvcYjTPiVTaznSuWBJklYZF
dK7Y8yewMLz4mtKMbubZyHb1A4vsO01yAfGghkFuLWgOisWHhwBZ2dpafZaYNgGE
hDLRfk9XpBwHuYPK5Fv1UK4Y8Yg2wD1L9I2SitDu5uPKcF5LKkxuIQIFr+yhWYhR
5aFHs/lVeRLy7adeCfZhpVhc+OjA/XQW67xH5dzcQMIS0KBJbmM2M1hYGGqArIQf
qrVVcF2rfyGMbWr6A04bHsQmXeetUAeN7eLTk3nBKrscEpPNscMptP6Guh4L0QwZ
kYRyUDtvW7nAnrq/GvqUU4in8Q0TFgKmMCK3dR9e9cUU6JVDPAZRB3gBx3g5Vzzi
wefH1uFxWn8Y45iunue4TUVef2oi3eZ0QRZQAmx79LzbS/cpTbF8i+Y5PW2jprGo
XJ7d6uA39VoDRvBIhmfT+w+aeR5O3iKNPtR5K6VtzSk6UFi08gaEOd8FdEKgZiD4
t0ah7hkMlCKDgmtR/Js4TdXT0lmTm63FvIFvkGccB77ZNWVNMAMt4eCfTMth/EIT
Q2ZmKciH/OgPqIPUFknZeMDFyq2WuolV2UCMpp2mTM7Lhbvkxn8JpqFk1bHZ2HeQ
zp8xu1BO6S5zh8ywXU21rd1xWzSph3Zr7r80AksAnCbFzioDDX+sQAEEFDqKrtAd
Jbi3F3cYyDwoiNElntEU7cNAl2agWYK3EJ58t6vcFSg/qm2ficpqCnlRygimRQK/
ki65pRpBTNjziUy3WJLJW72n5eXJFFZAU4k9JsrBXpowkVf6JdA6oLuYYrpV8QZU
Ptbp+Dp25MV+sd7I5VvsdVGw4ulTT0n4CFtH9SLEAih35L3mmQMtoR4+QzC291bY
l+n68Q9D5HTI13zWrB09abmiem3KVl7l2t4uLH0JdwGcWTd5NbnB7ATuQvrDMDCF
GgKwLwCMIJE12IQVpKT4d3B+XKvrm9/0SpY6x25drhsj8IeI413lWHu1OK6ZmdaZ
TIbIE6O/50bnQhpqMt0MHo6WOBKjokJUXWAHBlJHUVJS+j7TDRtiAkxyA0kCNvlR
MDT5Q6+OzY8AKYfnfAxmTJCVWG1lwpYH64vRj4BHbEmgxdIyfBcfK2lZmFcg10/r
1Ew0uE6ywfsHjlT8uWGXzvi1WjjLaFuwZbX43WcvPkPX3wguDORKPOX+Rd1OpxnA
40tEpBCUmiziBwYwlMavSoNo+DwYbkKp/ps5dT+2cCrsrTy0/4dhkrxy9DIwkTwK
n8FgtegOjP6ZeI7cdgJb6uuTF5+VRrq0DYGVRO2QYUsLH79cF9zcP2y1JHr7gpmr
pHOtmB0I/p1Bw0AbdBuZJevUh/r4StfpoIRbRrjAJ5EQuIJ+PQcbLZNPlPVs0ECx
96jle5YFE3Zqov0my1h0ECKUWHrmVCPnpGMuLuwKomZa0c8927QimpWRAwh9gSII
EEnFVZ5gjBrbKK2bUEDZ6pmna5RZO1/1X6fi9mrgHGdojxEiyG1Ee4QqESOFGKr1
dri+aphdMzLb9kolGy4RDjESXM1SdwmE5CjW0/f5O5ZHB4obbU/KEIV4WDUtRHXY
h507NtoGA5P+8Eh2PY8ypoOIbKRvbXOnsIxdW8dmELk4oLA6RQBHoerw13rhdoji
7PeNcDky2g7ZnQlDMlUi/0osEriALnmiW3F37GetjkZ2G4hew9asPuMSilqLpLCi
EjbhpRgThEd6Y7iJob9bRulB951w3wfKvui1dJCSpU69iFEBfnnIwMLuEcgOPk6z
nmt/+wi71YkpkUhMsTferRx5gDzTM+1jl7oAHvguZmgaYFHogyKZZdv+wp6tJyeY
DXcH1VYS1u+hBrCqx04JZLCIoNF/atQW4JwZGSfN3kDycNGw5MPmJASed546NlXp
Qg/uuI51eJj5Fq0cCtlY5KqrmvMpGi14gm6VWuqi1jhRali3iJIY8vpoSoejNSrg
ThC+OLuPESwcPM5JeTomjt5BhBvES5nzNabEOhgmtzCGDtgE44RQoaA+DuWznSW3
d6f0gy8H6EBRlKYg0QaZYm+Ml8HZK547P6ZfCdOf0wTJf7wy38XmiqpSBYt6O+jy
BlZwA4kUKVc7uRsycPlVJaR24TyrGTeW8s+FFrkKR5CcGO5s7Rw7VCXMjYFyypmM
87HV/kmWpIGMhPLT9MNeyW0jgonYk5Ufl78Ngeh2h3ZyCqXYRWBjKUAckoAk8/6f
p4qEs1/sZYeUtRHzO+WeCRjXOBaLEN3rU9p+PWsaI8oqWfYElXqab5CnUGfB6iy/
NrPBHL/oeVg/LVYvENI55h5AiZe/9fGAf3V2BhEbMCIT8cE2HefOs7L+7iVhtTHd
REpu29Mr1aIPxzHn3onBRERStGc/XlzkN4KemwM+9gfXx3lgA7iTcBeBgJh1pWk6
dk4q1nQsrfAQge2u5ikzkSTjcJMrPcAv/FvTr60NvfgsYtN6kJUWsxKjtXtXgyvT
pKKJYoPOZAiOYYMpjkzuFOI69seMAsivWiRZGBjiUtf5JJ0Q4f5N8Xv6eSYlupY9
w3SAsR2K4w/Q0Xcu2D0HDi1+143IQgDsBob2rbk6H33TJRvUltyWiywEG2ia51wA
BHt6vpeS4hKRNbp3BPwOEGAEJJUk0CyIbu26ZUVt3oUNMLgGX9LXD7iuedgenV2H
mZLnIJYV+/OB9JWlIz1dLiqaeIMBVvKGoTE1sX5oH63vZbXz4REHDo6EHyoQ8nz+
F3Ux7KP77d2ZC8xbSGHyzZH7zT17ybyG9QzCp70pPdRYlVHwEnJ32P84Foz4r3IC
g3Hw7BAhioPTl0EITP5ucAjb5wwpLFVRcyMBo9qBpAuKvIdZGMQ3ARvJ/EVfCAv0
T1hxQfv59c5LEcMl845KDt1ZkI4ey+N+bj+QzKx/iw0lbnHyC/QfkSNEdjETCgBt
lmvhTHHypUDF6QNFiSLeXJ8OEtQvMGdC5t5HrfMjyol02aLplwMWJ8W0TgmEN5KM
8RIcM3hliruLV5VoLyIimDc2+K6vdOx7aWkxJnnk1jHFC8bVrAdq1M1MNEJkdayE
xK3/PPbUhE9h0hRjHLa9Kcz2y0tlmr0eEVXWQ1I5k3n5R8Y+qA7CXtSgxdioKnvn
X4q00RqlYk5x8+qU6jDwz+Gjibx7RU1wDP81RZRdHwOCHiw4U0SOesRKqY+mZVLz
xTjKgtXExcam8K9y2++I48hNqAUdZMSeJz5f6LDvlHxMmB+N67818LNyh6slL244
rKOI+FcMJ62fNx2jXs5iJdk5v5nrb+3pBs+11QRXbLuayQ2fvr1l/wCs+sp75IEI
EchM33b7x+oM4DPReR3b8X7Unx/Q/b7M3qyCOhg32MBNLVPYmWC6OvZw6oUgXjDu
+1Q6c3MUd3QAtzSDV+tymxnzoje+/UBmWK4f5gy9pcn1yJ50nbyMYqMvuqqqJ+hJ
NfOTe7l4gvl5sfR4/oQPjeOdf30EkxCQjf7Z248Z92plCWxYFKHsBnXjPGKRVzR1
oAJb1qYu4cRg1QBXXwHweMB+z7zhijyqqYoQjIt8zfaUtJYrbSrM+eBMeC1r98k8
MbvOucKQ4J0SVUURdcxJP40pZeDn/zIkROKaeMit3/bfoh8fQfzJAIMORRtxogoM
EECA9nSGBFHxvvPMILf8OvkvhFMh3ER2t+utCVHSF1afi563rIpv6KO6A5yX39NW
ttBuWJydZAZVnpNs7JgoNUu6GEqmNq1yXBj8bibke5Phz1FdNYtc0HZkN9Zed/Rn
J4OwDFe5nmO4FZ2sCh06zJ+PyyxIB6nkVGDcmrmSuy9sADgUxTPV2lbGbQ4R7eN0
e0DAM9Ii9pjBN95U096ZCFNGEkzrVV17OCFUAAcrl42y+5c38eMAmXDgY6RX+BKf
8IWY2OBvX/DNIM9kLIy0/kaz5VVj17jtLldYKhXxkSKUc9ap+dZ5ButdeuP2zYaC
sNxX5r0Edz0AR/iRTBRlew1F1k0kbpuCZ5IaWBsyxAFsgUKhHZaPqibsqvusQg+n
4vXsTbvFfOEjwvHq+45yjU3hn3EMQf492x56wpvBdxWwk3qarNy8EU5o+DqkEwR7
8M1RE7gxpOkEw1nPwDWV08WVfm7MRogAteZ7FbNh+nQaeQudgeP/dqi2U/iZLlL/
QywbYPS3UwQ7fUP2I4wYFpCoSuFFGDHcXKKOMO/wLzVWaDAJ5x4TeJ1tHBcWn3n+
tUc2ZXA89FnN1WrQRZXlYWu/QkLFVkfQlJLB2LLa09KayiLKeButI87xZWBJC+AQ
mb23pcsfUEZgU8TSBq1E5/a/yGzlToAQo2VDVdtPi7bq0dnmcM0oO9vfkM0OojBb
KfcI3eeirig6PTs3PxQAtkyia2eRRaSI0YM5Kio5un9DxACUjbDLSUx7qG3YN2iY
qm5S/h5if6zyrLgLQGUpotSDu47BJZrhfhEw1Nd0LnKfSrMHBR85rLZRhePwAQkr
wAkS4dYmFXEkqVy1fM4a/fLQM3NGyVlv9RlZneeFyBCMnvqmljjj56WIp2/fWfPm
NvRAlmYx5reFa9FygVthckXZ5/47j12eNeKVIfY82/2mRPi4ljlCE2h+qSam/h7D
uehkTqfA2NBpktxhNEi6noCBc8/50cCSzskIHHpGrosTz1sPp0hOeiHs9YUkztWj
VUhCyhVuuuWTHspgq/6/CbEW3XJB3mu0eXQhGX7/qjV9NEIcIRLe8J5iZF3lmjfv
AFa9kJqpHBREOn0bVORHZSu36DbrAD/Cf9v0MNXyjhbRitvThZIbPuSmytGUl/oy
DyxyZ2RMVtizT4iqcqIq1iq7gKQ8DV0MOXDQuPSPgnHcSRep99fAMqCzuCAJDzvx
b+wYVmO9w5ksbkeFv1qhyD2z/dWSQW8sXZG8qnPvKgUjDGrsTZwgHn+hY9oUakjG
OWx+SEySiExVSIP1MN5YsFYyU5fGnE8a1gEURhJl+0OwB9U+DewYIuSC7EtpRAkQ
BNCbT01lpBzTY24rB/KfVJRxORGyua6v9F2+5WeL0t8+MCTS0jtSKAjWOyYLaPlU
n6XChZk85px6o6YymvMBHXxXD8SqxulFZzR6O0O3o5OlKP6ErbRaNRFrjU+Si7On
e15kk0MAqSh1r0fITY+MgU/d7GFOXwmjGGiK2ZJnXnNfXT3h7qfiM+h0Jl42yk4q
8ACxEWiA/I7XX0Jo6ZSN8OGHGl4Z7PyNHFB9DiDtzE3VMT+N9QMNBHKPTtU+DAXT
d9ybfMzGB6ORcVEPRKw3BE0X/FT/z7yCn8FfO7HZnUk27ThHn3c/PN1sa7TKw68o
BIgpPeiiQcwFdex+IENCKBZQHRwRyL6AWFww1rPy3Ok+I30Rx9s6oQiQj8vvWHKp
Wjj0Zf0pt7atnjLTGLnhsLBAJY6oobfyECbzInu3TaQV7oq08F8eiKXnpHpokKR1
ERAmJbJn3ILrz2u04W1yWoFVFjchXuwaAWCPJc0PkrARdlP6L3nQLDIxWR2X4JCU
rC5thJV0T1LwkSIoZiCmzMCkd/IW0ZU8rhAtp4GFVRCg76l9voGD7XcTaJiM4+KL
0ZoJzVM9kaMqT3hocEK3s7CpEXapTl/4MxKSmnxAqSfJda0J9jm417fx5ElLIOuG
gZ9ZRXcmxTU1qex9aAMcnCZ1V7VWMN47gm4RH/jM72NZU8px2LBFjOHn6Xc9g9rC
/Y7sQe1FjJKJmn11oPfYSEfA85HrpfuC9CHKNSbODaqFcXmNEnYnyffksJ3y/6oC
iAYJwUbz98oTEVgNDv6wZw7JvTDX7y8ICimgVulWUZHFKwK2rUUBFGCPHJEhUhPm
i5v4WHwI8P68GWgn6kPCgVqjY2rqSnMoEl+cB/S6c8XIDQm69PTtqag2UpLZgaFl
tW+p5l5oPRfPldPaD4mj7z6TO93USn0iEZ+t7klUG1ltYHFAzyA2FXcxGcT/pFPk
3j4pI6PpAC+z1rGpJ3A7+jNJoOjy7MM+8NaqBxGvbkZZAjhw+R/RdcJ8jrc81c0C
gyliOdHiuM7vR3ceAssQGTZJ6kzsXZv/BF7BG6AtMXMVxgHMkC7idycSQe3w8OyE
pinAvPo4SOftTSdhik5SGKwvY26eSAtyMpjF9+wwaSbZrYXHLZL6BrUkU4DIpXhR
sp5B8CkJWpSUqgP2D3XEAP47GcIpZaIRXCr9tRalMQmnqFlyTLhGvHfBjZkNGved
ixGWzbRQDra/on+4guJ19PeJnzkLmHexogtYtEtZM0HocMPJMAHv+bKeDcdipijV
8pYih/8syXKO6IZIuH2SMczBPgglkQvZd/guizTeZyy4WuqbETssaLnMtiy7hMaD
xaz7MmPkYdRsXdNAub/lZj/FGK6VyGptRWbNyHGJbYb0aUdOA8LtpWTGmZdoHBbq
rzWjIJn1yTL0rEsFBkN6+fgLZzHyTVKt7rQL/dzY5EUw+/EsKXlGZGp+rGUhSnjW
H+6blB9zjh10p0D5LSDid1APemijmz2dB2tXGTvvSGl0YOsA/Ec2unavYcKEykld
lKzLauPCpYXv+rBcBrcF264YVIOX56iKJde7kMVr1gu0XGGpa3pA+vrC/YVhR71T
WthMVKq+m8J0mpnwilP/Fzoeitd/ZnlFnCmVhUztAxm6S4t9H9Dr0kRldQxZFq59
fmVv5wsa4UnePuqO7c/diynmYIKXFjUdKNNpCEKL6a5janIAV/DTshVGunMEzZfo
ObszvHKhADtha1ucSAxwnKBWbw+q6EQbNrgxlTsg5J1d83Y4++TYAWaZASOK5A3U
5dntMOfX8kN7H6snGU8oULPY9zqmnZdUHzUFxDqj1DV2zWFCK9hVu7rVb5b23OsH
TPi2nRcpRhsxXUtt3pGaWSIE7hp9ot2mUXjl7C0BTGgbd3A99R7awiJnNmiv8hKX
CdyA/NF62jrBsr6+tAq4tVpJK2HhGzdikcYO82LLKfw7G/rLGyVTVdyVNcxjAcRK
TD2h5x2RJ+KMMya4DZF0c3b7crOT4uCdq1yzDU0IuDkbSINEvrcXNcLJ3km3DT3T
1kCEnU06uJRO0pZOWbsCWy6WBmZw0CTQlUW1hiWYhrpTLzIBWGwad+BQxxDuZioV
Jg4C9ofoibPINHKURDIsk7ilcubH+HKiYyOzZYe+k11iL1aunsRm8XiSjf4qTuBY
2ZavvAZXxrFeQG5FP/Zz1DzcW9LvE+0Acf2xoiZdTPE9Ruu29XP+k+Deur1vS2zX
UCEp4fv7n0hRqBN24PzZuyCRXghkCXcryTUxVPsRZhYmFnoPnXEDEDUegU/hEAKi
1gZgpBir32kQyN6K1xpxFtyYFWrA5b1s0aTzsd8++Djz178WEkSwoSfCgDhUmt62
nByf3VQN+Mf/YE+y5su/oqUF/fK05sOSIJQIFxr66Kx8jLI8NKmv8FSiE9Mr+J5x
c0Kb6tgtRAyY9phQ6MUSRk0EKIaY+h+Hz++Es8zJPUkohpJ0Bahct2F/vdYf2ks1
Jpy+u+0NmiOrWHfliWKQz14IKb6wcaYP2elSgn0SH2OG2shux8HSuB3tdGtGcBD0
X00XY4z13EsWtXx+Oiw60nlOgR6ndDnKd9ZaCHvGrPhFiI1t6TOiDwcfUQclR1/4
XU63mhNF6/t25KEJY/+NtQ0Azi23U3zuEDKgnsLn0EwovmKdWJlCEeL17HUIUrpm
ZvsjKm4nrkksFBoFtjWBP5WZGykHUgTFLh0NAmJ6TjLghyim/5JdHpxoHrIeHFvF
NVIEQE52gZAg6Lbq7tpz8JwWTttX4OP9zY9REhRqFTsFImQ6oIzDbIdNzoSW24gh
5dYk2fQz0FDohjBjHXMiPpxoiyZtbDnkbLhA3DkYHkbBbjxytrSSDrJN5tqgyExE
xywYvEXo7NOlP0zoSQJFifvSbJQiztw6M4SDERPcIiVu8Ik7ulPQ2LIljXGaS6Jb
BuT1BTYBil7kTORGgUsgj1weQtvfyV2Aisnz0jt8L+dhb+5NDcqjZgwdn7KNbHNs
Qupzb9MUC7SHc70S84oikXySdUdffTuo6pi60QVcNGkqYUwebfAMQisrNmVHZnPv
DbQGDp8ZbBhOhHd4btkJlFQPC+bII847rpXkWOSY8msJeQRclsfwZPd9o9V0gohz
wg5Qfr28/I6PnwoTMWNpVUKn6PiBInCs42mFbnuDOAaSgRd0HhjK+JlwdC1hDb9h
YoZK3LBHGvTDXvbOp3gCFDuKHiETBAb8RnjQga7d4p1Bw6f3T+4kUP/wxtOMRJT0
Leu3OJvAw/EQhc11FlXKMslix9bLbjaeor9OK1Iavlmg4CU8FacagESGRxuSvPSI
kn/eKeSXLrOirheZuvD6ogxcfDya5gWh+k/xcdTKajfpe2hgwRGM7XRhu/RfM+8S
za7GwWj4V/sT4Ie4qMCs+1ZhKYpacZe+OA8StsxcPOp8yzwhfyUU4ZmQnpaxPd1s
4mFnAXY+1WpeWVYPCUzYm8f1dw3TSKgFbpHfvwryc3mN4x0fm9SC+Nsk2OLSvvlU
hUtYheDxQjzSFfsBNYpAtlnVTVFe4mhod6HR1UZWYWsDKiYVGILpdILx/2GGqxNW
GuF+2itQGXmV2Ta4DGmG3tIpoSJuxbdKQuHTPxmiY491zJFNqYf7EvbJzrEQN/Bp
TN+YoN8q+YJSHlzdkAwoRXl7EAUpY/nNU2HUg7uS9Hck2fVcOg5tUcyZf9tKn+to
Gl9DvBaqthiWBT/hQIYo2vpQxFC7fh6+oVcSsHkmdHMv9zFHVc7P3jAg4zLfWigh
3OhBZ3mkfl/mS9GQ0VkHVmI0hIxTAQW+4DNzRhqyvfdT0JBt5MDBsdJAd1Jwmkxe
M4PNPfzRYtq+6jQAeniqE9ob5bu5WppV5x7ClgnwvOB8X8VXTgtAt309bpYjqurd
poP10TR7yupw+fjzuEoQU/P9SkAQgkDTgsO9oGfN8UpL1ONRcIkxsNwtvlw/tWYF
H7/B5AFtEpHvNhUZl3oz/H4CC2rlGqTiDznG530OXWy60RKNXIFOKRwViknyuSd+
9deFpmDOQrqEcXuEwCh/LOY1LELjVfvoVYOUoQt2y5oGBgm8wzdfmE6LiOLM0OBd
wZOtE48Wr096xHt2RHStZ7oXeWa10YH+qF2yj8qDms7TNqF9D1KG4PmM/vOoZ8gm
ts3h6JBf+gcx3X1S09bRXK0YZMwOkxghn6tU1NtxYTX17+wN9/aAnklZsI95ECvd
h426PtOrKr0bpT0IRmcwPKGfLY8RY4l2LYTW818oGniXEfYwkiUR4iPMMG3C0PL4
TunuxHrTMQa/FJiZJg3MoPJvpIt5anE7OO8kLtaDbMx3OlMAkYsROzWnWPIFiFiq
KOKXsEEAM2kT08QQRXCYvtxqmBh6soZgWLlmt2mknzwZWAlIymm0dNlP/mpu+2qn
BmOIP80I/sqNGQU2b89Ze+EGNNH4Ei31+WX8yHz2o9JPjM1gmAkSS/9GMU33QiOj
AXNwUN8n08lWQeZLaZG0kbZ958JBRVmxerrTO625Brrx96JSZWgZW9+LQIWwVrh+
qji+6/70Y0aynemG7xS0wKq/ZKBPkI+wPNSrmMkpQYqriPUA3j48MhmW3K7eKfPl
7cura9LYCOXUe+5FLyOl/FtKq7v8QIkt2BWycLi+qGXhs/273Ooa8XZIIITtP3T9
4eTClFYsQh+d5HbGFPeVJKAuGG/WwqMcszyq2qJbPpc3ti809xLUP/VVryf3vRG/
rsMl7fLAOWfT3xobNNMmiUbppVhyOxvUoWN0M8208SQMAkgBXNKydvpS0SyFrwNm
666KMIpEDvaIWTanXJiw1JRX786rxCJmbgsmDH/SSafpsz+nTn3AWhfGtnmgf0Xp
mXAHDgM50ewURcLGKQTAW0OneTC6uoABIcs2xCJJaQRNqm+fRpCCNRCwYDK3/ekf
4z6NvWuuGqEt9tsbiCW6RrrlOBkrWKqn3t86aqrei5XtFpsgtxKvTRnofRcpFDD5
7RF7BVkae+qX3AjLbTXs8WsnpwS5mbu5JjLLonIwGrnB9qxS66CmMju3/Fm23ybr
wEtMZgOfmikoMwimYkCeUTP/oKMt0yTBtaSrumRZqWASLQr7W0qxKNbFrfji5i1X
QtSG5pQ485VuzPdk7/hTz6PKGXWLskNYsc8/I7AX2DZ69d45slWP56zxpKBHsA4N
tZ+4AZg5FZXd+S50NovdfbZM21qaDxmQgpm6Y34ANCkGrN/QPW4LqiKJqRZAQxby
kZtcqKDd/5lSbPe9R1pqDjCyQ1B3tuVYpFpiB8sk178/Wkd2o53rbq0B6H/ZIhOy
MiNSTnM7O9UHUpY1bz27E+9iRY+geHSgR0m0ZLSRy7L/EPL7f1YRUcjPCfSisUku
DG5YPaS71M25ZCYMc1OFyQ73m/fc5COIHKJacdLxt2PuUimFDUQM63Ek0SZbJaoA
+xbf9YsyqKEQCVi7vOejPHm1fKRVCFfqDc0+eU3EeQis73dpKDwVlYgpHjrWS3f1
23NhY68OL10HNuz9yHj/GkXZ1nuiEq4l7DINn4JLeiQ/TjrzwSxiLBrmExGel9OD
fooJq6PlwtwztZ+/ZH3n+hCcaNhTBOwhzW/CJiVCfyV1WDw/PF6uVlfR1KcMNTBU
Yyfh0O4XZNcHiC0pWZHMmhxKRZGpryBhAmgV13gMYHfKD4FgwbOsg/x0H232YEP+
x9eUNtg39b1B9NN7j+saUDu1Z3isddE+Pmi/WV9A0VgzlTX2d2DKCwgcp8e2kkLq
fwlV7SPqVSvrDSUrg+0Q8YELnar6JxAFsZHrMd/zeKtO7DjMqfFTqj3JDcfSJUFD
ArW6QyiFLIDgAr0SxxMZjdGFMlXO4ufF20004EFBLbPn5LDlT+ZABbB6ka7xfcon
6J0OAkrXcIVQvdQno2gWasCeymFWOPHOvtYRgKs3tMnc1dTeLtTpUKDrama6Ow4G
i0/L31b8JV9CWFV9lA214MaEAHEsP0/VZOD75NIUEjYcNEHNIq5D52xri2FFE0yV
yMxkStg1Tul89dMVNnx+dRmhQY75w/wWv7dTiHfwc5KmG3S8wMiXc/ev/YJqdikh
awNP0AH+L+BcBV+vZJHEHDtzmtY3r3M4+C7hyI1p+3kX1/toRYAz4HXG9re3IiS5
yOome0efvffVtNBlNNGi8OMv058rSYPnyLTRD9c9ygQNy6FdQfkbofrb//nyi8ji
q99dr4pufSgL3hlSwd/1/DgDLwHv3k7Ba/wyyHmL2+MCwJfc45Y3GMq48NGH+L0I
2dVrJkyqP0RPrHr6sUE3Zn2EJz6dNGQUFyVkJSyO617032gSffZQn3o45Byj2kwZ
Q9fpMOf+uUVHmhsWxanxFE6INxbekxVhpqgK3ad5lIT2fHbr7TxdobNnU4M0kIfJ
KCadwfIgz2pgXsoYYTQIkrTDJ0TVWe4xWWMdSQdOaOHwVzAnvWzsda7TliGA0rrg
JloGIsE0V1AKJ3fRnyxk0ljCAoYhpNTBDE9Y3KTz5oX2upnniXe+hCgqxix0sPvp
TG9o5kkan9LZkXrRjway0sV1UEum3z1PSDvNb51Wwrwx13UB2KFIAGe6u5CWOogS
4r2WWAXKMxsqFwJvh7FYyuf/qZBSYuHTHlRkcTmy2mTtO9D7QCjYG0wa4AiiEx6+
TF+2KSgorgwWzlIM7BwOv3pAOfnedg7LBxWmcEX6HwsERbcloJJOrBnGQ63wN5iZ
woA/SVxvqawKNi0NYqXYVrWylU6/0PIBNWhpKx5VyAg6IGTeneXowdY192t0+wTA
Rq7lXP/Y73TNmNx7TJkzyXcDcNdK/uBGFxf/Ak7+dH07/pkgl/w4XfgrVsMJ2d7K
1G0iQNTM7ZtT3PUp/mWUEmQX6jyEeHKpmXh/Vih/YuDT3kw6KKQuiXHq6CKPc1sn
MmGFJvpBQsiN/Hv3dGX7KSV6aWghH+AqFGpbtU90z44ZoUhYwvtaG8GcvbQkcnf+
/8hzxGwxrf28K4w2Ezt1LE8sV2wm8gKV31Fb9Jpc8HrdJ8pvlyAnIWu5FP3XAWbk
HDlkMkXUdiZAn1Cei3Ty00xkH0P97u5AGvPy/UhxhO8Hh3GV8Hj5+7CE4PR9isoN
zmlx5fskHUj5zCMN7spOtEi3ehjRo+tRLMUs1ZpyMLD8tHkdDejeTr59tAdTLiJp
Bd5JZDv0hGYuREIMHDxAtEsd7kVLzR80mhgl2IgpY5FLgK5YVyrikfU0XLT8KWjI
fxVEO4bctElabgtO6k4zd5rxLupUiud6rVm1bEOLhEY9/1pJO0rJPaCFbCqEgJDJ
1HeIfNhrHGiExfGyiqB54n2SclCzVNJZWrO6VR50XrNOXeHewaQlBdzMitA/6OAf
3wWdn479AQ+vom08HreKSMNeFvSyZfcUnQUVQ3jvlhJZMfJMP+k2aT2rLgVaZDt1
OAAcXkrB54+ngdKxDxedbGjBajS5QFNRLjkldLABfCofTJFf7ucyJZphOvoNz2bK
86NC/rAJ4A+9IYN5piAGlb7v4FeMb/BwY3gKjyMNMy8m0+lkzjisq7N7VpV5KBU1
mvPLGYI3oCmS0BtIwoo1TGA4+BK/jhnhzgF+kEdpqHdw/VgBKSq4EZONtgBsqIqx
lHF9lAEA0FBgWeI/ai1eu9ewEwy2FgAj/HobzWKkP8xHkrfVoR67Z9dRzV398lgj
X8HDmszoYfv+9aYw9VkSP8KCG6eqOLyw4ULlkNJuLf33Och8Kx6YtF8MGd6yxyAO
j8k4lV4PaDjlbD8394uJNY6eGBwwGjZ5NKju81WVtOgECEXg8sHLy3r9WVTdwBKY
Pa2kvn9uMjiex2+FkGk0a5blReDl+ufXpCs949Q1jE9HS58xa6/7ZpC2jvaEF2R2
FgQo/ilZLvN9/LIAK/eG2VFFLWkTR+Wvnikh9RmvnCwcrQBNqKDjDkxsMw7DD9Vn
KJE65BNB55M2fhvGWwT5VCqwHASfK664VnIeo9XnsJ5tAd36gNyE0PvTAsV+72sV
9zNGgIq26u8EHg1BeThCXztuA/yKGdtiysZTqjxN4okS/Ts9QEIVNZTTyoycFc2J
Lpin0awYPF0PBCE16t2G/Nj4fay+RkLIqIzgcav765vg+X4ntQtL9/uw8U7jq7l4
nsM5HoTfvR2OuhCwYU1O34vOnQS5a2jHjjGzeyng9zn3YjjAdV00NMTGoT9VlVxr
7wJHulNQNGF85IEpK3KLQJRCOaq6yRkng9Riq40hg4QztInBXJF9ohkkK7CJM8nL
2PEbcRwRR7j/LNNI/AwJ26SUu5OY8iQ4dZOfiF1lRtNqnqFEHA8NvBbh6qSE4v0W
6itId7HcuHhtUkN8JcRhkRz4UNQJ1qgpouW9Q7asVmYtQp3S6dMApKXQ0ry6l70y
sqnKkM7mnEkjAkEcS8d+Jw1sHXPA3goGdwif0NW8pKyJhaUziNcEgNXBcpj/Tb+I
oga01NebbKKPdpxFL2sUNN64tMzJ1EqxPTaZFrhN+RFFrfVEovhznebNa8WY6iyA
/wHn85st+GEq/MMY8UDYp55sCoU8Q445pfS2enRS+75tIYZwIUJR+0sS/Vn4p0Vz
0+Ni4QA06vtbN+REu66DG0p/5PN1rH0Lu7nfA0UMwoU3WwOAlKXZYskwh5qnqxb+
JT/7kPH0MD5W4JHTXSqBMUs6UsQZkXhAgceFxrbspckl8HPv0KBT1noyBDfqtg/p
zan8sDqBZbsHZbykVjYDeu0EMFYya3xLgB+Tmldq3jw+DdUgShGhSHzI8QqSavyQ
1N5RIrzYTawr1y2DD5tTxHIE30J5RICzb30WgnhtZB7HdSlBGLfKkI/nq6B9H1Ow
LfQUFpVdhRUn6OqZ91edgL8G9B+s0r+vfCyEAc+6x7lO/JFeM4mxlNwfvbnk4vfS
kINsmNx1Uto6/XNKVT1i76DjMYiUSbLhF041Rfkxn3jvscbiQdSAJd2ZRH30bARY
r4QnJXmc7IWPMvm+vF6+jgiiaFqg+mvQcu+OQ3hBmiY17TOfPQWwSkAY8GbjzqPT
2VXY42FH4KcfKy0lqKPwlHqe21qlFyM56TWxYtPmZBdCoKY4BOi8cuw9Y23J2nDc
RXYq7gTj6ZkmKo+xv/T75zMvmaIZLVUZCQTlw54BGJs2dl7JS4eLJ0jJ9mxwamfZ
c7cdKFwSIhBQqMgtK0rJBkPYxImFzrcm3I5HKZIL/MftbkOgiw8ZrFiwhK7+MGLn
asP5QxAZv7c60DTashoEMg4+giPdrtCB7VILQl1b4b4P7J22+yA4Kh2Dp2YrgXIM
n85j1uW4Q5DcIIeVZ9XE/ZGEln5v2wv8ORcBIw2FCuXUvliOCGGriuRPQzFhb/VW
oJ4DNaEk5BdbiKINR69w/TEXDaeBKSPOMo7uoZAqMAL7xb5NEqjbO4bAsEcJXALc
yXuGdxUTZv/oRDzQcTYVqAhc0RYplVGZDeWKqTHcQZV5ytmw2Ipr+eRsn6y5lk7c
HTbumuUI3m8DAkfKT39/AmOWnTJAuU1mV/Q6oMqZw++chyA+ieop+BumtUdu6ADu
DjBi1Jc540dEc1ohNNdL5vKRNPr12khvTeIiRxeJVDjJjMSDFaG8Auz9nOyTLwLu
0hVOBsqUm9b6hsSfG7prQ1FGt80cCQd2NRqnzIhx8kmIPB+jZgSbKDdFy6/fHjXd
hI79nq6bwai7AlOcjnWGpISrxzdBlYqp90TjRsjVz+ahRtvJVGvtA7QY7w+FJ/Qx
mAvByjnF2KSr0u5poaK7Z6OnYosqQx/ztwbXegIoG+1wuPWO9/QRKMOylqHddm9p
EWklvObD6cj7C1M0FQMTMSFBRYRfL/kbd60aNkbuNx5uVnBme4nhqjUa9Sck4gly
kQruz0cvXUagEgXkKZV6VOB/94VS4krNRvJmBo0hwRhlpc0AbzTzvEUn9C6n3nTJ
yCGNB8mOJAlk/CntLif7Hl4NRyLetPCuW962Ld19z2d8Fgv7uzOzJgNXDcMztPHY
us2QDhXVTgxoKIWqroq7z+rZ/zwBRaJADEDJ5ftzSly88u7bxZvK0J04PiTDnLFy
UcurEJcCqMI3OsnN8D5wPWThHX950BTtpRF5rkYAuA6EUyanT+bc6N9zTEKPWWxK
0oemjtxEFGhxZ7TNLuaGf5Wx33R/sZjI7SwG8G+XeIKvB5J4bccvHkQQFbpvEXpf
adL0zL8+xu0yLbxKkIacjejcjWKAIMK20EfYgP4mbB+gyzz4cba/f/pCyBxcd55P
hAW5awRuwG1v/Xc7uuz6Qc/djsUYSGzdQLOU6eCbOIoY7tYoczDV2MfSqgXXfojW
juS/C0RqTjeUak28hXIsoT5gE6XdOE05/3QU4IDY2b742jH9CasNHJacncGxS47y
oApFpI8IWA+gvTdO/8Dggc6Ei1b0Y/sGnISlnNQceE6znsBLHFjO2WB5GdO9PoeI
l0zR6rIq8v5UyT3omUxPlgeH5O9Y8ktibjLxkXht9OBIquLydyi/lWQ8fy6i9fJv
msd8D/nuizimEErtbd+os6y8cBC4BmHa5T4jSCes+4jTJtquBiElC7uXNrvhTQUU
HAXFrDi6+2D2bG2HbeETuwqOCivYT6S0JjDF8S2x7ne0TAhkabkNklh+PcSw1Tp2
OFzzF1WUvr/ObgwljiRsn2rOmh/jUBYbxWdEdcbUk5Ov7p42QP0An79QpEjx9PFh
jZW/+00XdlWH4Thf/ihB78jJNIu4fAjbH93f+z7beca20afxCGSwsvT1uziyeQzz
l5XP9WhezVHJP6Rkz4rUcYujMSIbX03bcnhYc+fhb3/8UJF0di88ajhGBWuU8dON
Pf81Oo83c3uS8JYmqi3tuMQ5j9szOxzvALOIkkh+ogQjVMMALdvcHL4pN1Nhyss+
0TQeowaqfglpM7BFm0h0dwKolSag5lfoo/yu70bVHgteyLputW8uZ86HG/qDk0mT
ncczu3jCS3sQ1Tnc22IkiSMPYQ3e9HXcZrUnwPnyHayvdjcho3X8Z30m/DgoYG2f
/zuCyeBqu0Zuq6BbH7WLSun7HiPzvUFV+D2DLKPOG5mpwCeJwusGqLv+j2PtTpnq
Mu8ypu9lZgm06ztpGRGk5Iv2Lo6RerTFIcMRVjuLXyu1w54JhmR/cQ03KCh4KCwS
uKsFr386F7bMpJvWoFvfuJKPM1zdHYshVzhOjPeXZ95HonbVPCwUnzPctX+YXJ9A
2NAoyewVNgNpddzyjMlCLNjlAwFMVJRS+yPGERjvEzUP9OwBbXGm1sbyj8qx9gK+
hG+CVDloXfRw+ixfvFoxREvO+76zvdoaZdfTu8IAjEJQNXUr/d+5b7aNHEQEo4z7
onP+Gxf2sUZK+HfYLM96l+GDjlc+1Lspv1CKS/m0GsEHwWCnHFxRzGle/A2X6ul8
03bZiycH5i9alIkF84x1EgLopdbx+VSikEns1SZxiV+ceS1uinIp/yBnIAB49XXS
MZPDSxc0cKv3UqGeALJweHV0sassXMkSDFllSddFK2JjuxF422lfx+2T/uev+K8h
M+c1SppAz0Xgi1v66MdAmhPeEdZCpYqz3en4xDUT8bE+c5SPHpxKeyTvw1K/yATm
w9WpXC9i3Io5EjgOiZCwAkmz6TyJym5ceN4Uaw5XopduJ+PH8HJ3in2WwkkMze7s
PcZqpU0mqOlLTD6Cdd73vKhq/j3ge3QdcXOtxo6xO8KWIDNYHhgpLW4sujRpOeWj
6zq6pck42slxLeAV76qtGE7i7RteIfqVbfjPyUD1eipE7h0BQWSp9oLDIeAt8s4N
KjLepUlw6ZbQ8LYM3q1Vwvi232vPWQWFjjtstDxQyJvpTwOczRNMPBu49kEYJs9i
9ZQEHPSSf7hczQBCGF+kQqr4clNkvrUsSFu0rn1C7oHeBXxg2j7usmLDXyM7wPGe
nBnWpPwMuqCy/AW5dHlhIOcdVN4XyJabFmMs7QSWS4qsBLnOxdVUvDWZYU0r+P6H
ripyT2SAYp6Dwe4iiBtbNlta2iCVF08fGdxJZ4zD/sX5XPVXelfnK/pPfydVoWB/
vsYGst1kJXOc3L5+GrKAbabPae6kg8l+yODf557jYSnKel76txRcBc3GCcqjmh14
9uOf2kurBsbvLWUA6gO6KCuTffHmPNviRV99MiVMZy8ngjf5IuykVxr1zhEUTh7m
+apWeCg6qOAWqtExUrpxgJOKTvVWFg554ZakpH7UR/gGDMg0aDBYwA6duarMTOdC
ku2DiMBIt61tc6iZr16O69UiTB0YKK7wS3GPsxkg6WsrUp3nx+T6aFMgNSolTQWX
urU8lmBAsyU7TQ/R4lI87li1lHALYD5hNjKb7Bt+A35nQqxZauV1G7MTro64a2+b
2rnwLsp28aUYg2MeJNc09ztr58RoYLcbozUxhLgQfjV/MppCTmKa6QRf17/RsxXI
0U4PPpqx3+Y/+9UcEvrSxKJlz2fPqagsDRye6y19Oxvz0Arr7JU86MB05JjhLtye
opPHvCCBzp7Z07l/QB3N/xOihBy5P81BNMk7G6LJWzTD1vg7CMYMoiuKrsisvom1
Qp2325ui97O56qkC1P118zpqlj8W5hhkulmb212PsBINGjRQWDYFODPWEJZ5j13I
WChMeNzCr7HGO2PNf+M2y24q3aYD/sLIg99dilZG8OOyYdQ9V6vuinFE9IcU1bN4
8JLXdLyRALkHsJaPkCCANQIpIjkE60exqD2+MVv3VxgisHuzwphhL0qcCpvUnHZ6
bO7fa7oYRr6RI75uHJDrPSdRYhAhjmPTpqLaFa0PUBpat0bdh1CUJkO515o6sUah
QcfrY/33bJfS3ML2fDUzUpdUDH6e86CghqM0Nj8LbcMlOQ/tEU3ZQQ5oHjSCjGgh
d+TZKGgWieNflWqEOmqbB9I22ji6aEuNZN8bsrV/HSecBuSq9+kmXMPoKSOp54ih
YZdRmlTmKgH0L01y6TggD6ih4Ok2jiV+k6KQ/217yr2z4fI7LyR1nVOHs6Kz4x1Y
42bF1zudjD/3Ac0mV6jvytfcGLe55b/Elt9+tWqMatXkngg4ykzfXt4UmsKu8/tc
mwurihyphpSrNbRihIokw6X1vszSN7+dFnGw/7bNK7KEmIAsk9GsmPSEiSS56hhk
XKCHQT8J9oFsW64Ip+a9HOWdZ4I4KPedEqlownnACJwCf0WyJgUNYO+xQaDm6dtA
JCXsPURlSiyGFwEm+wzq0eQ6GE51eiRn35qbvrbuIDlf+FsHbtO/wovTrQs7BiWf
EdP45kMucta/z+U9ogmZRiQNtA6rExgdscm/dkqFtt/m+t8KgKKMteQ7792TUBHX
QbXASaj3S6nlIgthGBkMoFKz7ngFZsZHrHB64ofqKICqm9XrmPgwMjUzUWPUa2+H
2FFayPO2/peT9FzGoHKrym3gx+m47emfSv3KhUyIX6rYZAIwg5dmrqNg01fEiTzA
eJMyW9/fijQGrRdeWQr/IA+NaTu/mN9r0l1KdO64EgsmQarh/VcauQR+/vf0JjuB
/OPPcSCM5U6wxU4G+bDr2FboVHEHFJU4v3zg/rx/0pMB+bh5xHa73HNYPgdfpoc3
D7prvQ2fkFHkbbYXwuVne6qo0l8IlKTAqLUgWsF3e/KWgM6opIpvA/eJIaWz4H8r
+mphme88JgciyAIPn2Z4fInKQtd7ejkO3ia0jxC/UEeHNw2Q8YI8dQH5uP1LsStL
IYO8FjGT1ju4p9Wds5O6X0fAo3/6lA3xr9KS+/Vtbq9AV302Gd/wWVxIYc7yeTCA
mv4RtwwIF1dqpvzejoyx1sO06n1DAFlmXJbxO82CwoBtYlSBw51hE3cnTjBfcwfs
V1Fl7dZtSlfRuqwH9WidDl4WuqYuYyp5UBkGdNq9COLcUqTeqV82aZ4NhY/ObowR
gnxWQkUe8c6Flg0lcH09VUApnNo3whEfnc1l3THCvM8NxOl3R0Ot005Xjmv1MxsV
/q+7r2VSOPVOhbpOSsMWrsH2BMW/s25QJSpF2PThVidCqL5eCjYqvEN8AwXXnOLR
Dgp0jzvQPQb+tUH7ymSHCdbHYHSgq+39uCFlgHXKiAO3Q0ageDdGCvwCZWbErdYG
hoQEnemMgNkp/BGDxtP3+iyvTC1ey10u9WkXcaIe8RGxuw2ZOXmH9YQJBlRgxQVQ
q5B5jLZ0N54Nmy7l/gW0PdVaL1O1MR5joOVqMXaPU6UzenyGfjvgxyM0VDQ39nwq
eCKpX4/41kCiLDOCY6NFncgrsSzuQOT5S2ONIZfHngwtN7uzarKltsYrj7MPKZgN
iy05FGhTbQQwx3lf3KIwW3nurEl4zqVi5Ui2jF/LMAcR04R/LQWCdCrXWLNFNySl
DjfEfjC69nW8Bi4Xg3zuYG/UGo22C4bh6JZ6ORJxEbCqhl0V0O5I/YtGud2PPP3x
NvAJGXZcBdhS+MAbfMlXI5kML5gWz13xePLuYZdRLbeZsFKSWMCHdEdO5vKE1W3B
HsfT9zvnMvReqD4pOGDrGE/W68p0OeUJWk3tBARj38YLbR7MJum1u2tUZbLTlL3r
FrRh4O3zO8xblCV97NwM8Z0331MwXFo7hqotDapYlgoY8dbm16/EtPQTPhcYMG39
nUpHDbw8hTGLVADZ4hz5+AIcjFrwuUgDhXGG9kl8kPkqoVsgJADbfG0bFGokiO3r
qjL0HU9J+HkZ+8p+F+ThZjLByfkeEWeKkS3O4SzvuK5Hoa/vgcbk0UKLVdETBEuz
jYI7HP0J7af45/ALN3KYLYMNZ60GgRYmjCepJDbUOIWuLMsFAT/xRhYsiN8l5RAk
/O4ay5kF0FN9LPefwL3J2bWlT13YyfrwpTtj+F8rypf4V0PPyhlPno174Jd69DOb
QBQPLpHmX01UTOt/gZX3+rT2v9AVYlNnCW6HuGo2g2Vk7ZUgBFZSDOrBRhoYAMof
oFSIVgEhc/W7zPGidtLzibi/y+4MVBe0nc2p8RqmX6sW+j0UA6SbKqLirzkisRje
2qfXO8+6SUMAyU7GyPgbk3IVFldKdHulFV3hI3zsjPMY0C+VvwKLYAaPJw1tSv3y
AzgJkdu+lBUsYQ6jzRZp1U7jit2s87Scx3rgoLY+8sVeWU9hPV5vINMN/ZuaSOno
9UPuhko80polphwkLxR/W4ljHcJM4zokbAeRugMVy4uouCIGGxbU8VuRYdSBtpXz
MpT40AExtZr01idFkQqwggPDBxuKuoS0yyQcOcyqY9VYXxOMlOia8+cz+OMplj8c
iiAIf19U0zsq+3Sjy8OAb6z0t74CUVrhm0GjQXxmOQYb5TRzuJVrWs4HvF4hWVbJ
Pgxx4pvofMKcpBDKpdNsyg5kttDsr7e0uUThXZTdu+qOCnVDirtr4Xc8JUzIgSjm
lyqxHxQ6JfZbXm2v/9rQzltmY9fFx3dzHZkLznimQqkGBSkmTn3xkRQxaoMMgenz
M7QiYimURj6jU5Kk/9He3tNNIOFKol/wYQGp6S9SeRfOVlFdcLDs8yw5ZpFAgiUt
n8BRjQWAuZBsPpbBTeD13CTUfWpgcNaODBfAU5zmVMKq6N2KVnHHgpeGc6IGGJKo
tAOY3ywQroOegMhTVCJuEL19aQgRg+xygYKtj3vrOdkim2Lsi6vf+YS8ucn6ykFH
6AEBj1/UzUiaPToclrYbwK9HmdOdv00t+jZ0h7pvIZcgtQ89cXjdCJNbeVZc7Cgd
KgA+EMwVWdZmrPUv7i2dh03y9kwN3Wj7bAr8Bd/P1YF6HhJasP2UWfmIRAkbQfIt
pUX441CdVuNKtn56bFitdmsvdDIKnlUr2l0uneWXPHq6vOysd2njeyx0x/M9kDep
xc747KYKfCVSdYGj/MpVNrqXka0X4SLb7jonNtqQMUaAo/xkl4Wu4JEU+WCukmWO
31Eb1gycZ33IPQt52hEQGlohLM96h6wb/j4+VAVuLrsCbdVBdpmo3vCZUJ8KbqhK
gXgUtG8phd/AJQ39rPf1T/o/Mo12llroNKsFmZUxvCNLia6m1viivJy/8oLw0+Jo
CexDW46UruFwAVXfBlQt1S2sQNZMSAKFRRtUBRu0MhoLO8sjptz5ZNv5CW2woPFJ
ALq3LUiaGvb52KUKCTuVm81YNJHj7Hm7A6tG6TRPHlSWmoEm1Uvx4axLm7GierAE
VB4NHFxUiIjjbbwd5FalML4b5+BZwLTyw7HEqo8NFws1TrvjIjbq0HF0XWQ9D+X2
0v4ryg+3isu9twrgtLhLhTl90P+btUCyrhnUXnbT/R1wDKOWcewRlVrv5lzTlOnj
1n28sZpkRuvc/+Z2BETF3Drkl/nKKOBqzOTMjXlB4bcbzNkzEpj/f/1a87yZKY4R
sEMVpLbkwqzLTOge+2VnsncJrfNHrv7JoRDEryd9plDNYgac/TOlLBq/0mpyKqOd
mU1R4ZASD9AzHAGRJ0BrTzXIhujAyHTSS8e2rKiLUqLBQmUSxu+G0wvqmhTB0cqi
FaQnrulxa+rjaAqMBLWa775VL2G2nPgBRJE4EArDJ1E8JOyCKONov1ivYnIM7AkC
NjDIMQN8Nr0kYHBza2bFdxVQPvDp09FOZ2EkxshXVawj84IFj8WQ7SQOPzd6LuXN
69IlXvbnfXCIiQcVwxVLvA7b0x4W1QkJ/ktve84IY9wks0fS/hgu3d7iHlZGfCbq
lGOxoMQYa96thcOzjtJdzlE8WczYy72NE55Z/aNp2hpu/Q8+Ea4xfQlPHs7A6g8y
u2hfcPAtSGGS7VU3vq27fMZzTRFKLotaC1PhDfUv/OMLOL7I/tbiakk1Icru+aHX
p4wgL4zkr9UdsK2pnBfT5CvVkcVH2lH+FXcryEt2KCf93g5zKrUQ5wnLCQND34Fy
nUYgb2CiEkSGfLb2Z9T4AW8tpp6uPdoxhNmRfkEKPpDk6o5ADEDOdHKWwzJbOpEL
oWfsk0m39pVxVL+p65Pos3x09dlGQeplUDF1hqBEl5cmGlrIHxN72xOwEdG+5Vi/
4Ki6Kkdh/ePqGbDuAB94vUokd8Z40v91cWaYElmfAJChh46RpZP/6smZT6kZzaxT
lv4WGJopPvVCGDRy5+wFkGZueyhO7kUdGtCd22tZn4UXP+eM66d96t0iLWoIuFDZ
lOfOIoSMmaEq+zGi2muvHLp+HYvQgeZ7sR+bgzhK6I5YvsOTgIRiq5XDKiAt2Mk6
ltBWZAKDaYlVv00KBq6p7LQIHH12rDgYGzj2z1X7qChRegNmTygeo/d6Is0Ev05z
JeZwzW6biopDYzW8PJMIBU99yXwUMwghxBzLW+7yokcfFJMtflHAAvUTlFCOzlyj
4dxBQDz/sUwe1os6D8R61m2dqhMjZfwFyu2N/gMrqrx/g2ny2F0ht/XAxlcUTnkq
lNGyb8Dy6GDtxwMYQNw5zOb/TgRVGq8IW2aWHZ3ErcfjhCoohYzw/iiufHdflGt7
iAnBstaV8ucnxTkCHUXEc5yKpd/IJkIsZ4ajfiNDaTJBrRePbb9NqKw7cv4ND2TA
ERd0sbhlY6uXzHUA2MB4AlIicjTWwrU1zW46pfRg6vyOuXLpcq42ZTokqvLfsOq7
1a9cUn1JK9PI714kl2EfojueU7VvNnGXLX5mCPjMs1AnG86JXuGQNvJgR9Pug9ZT
OwjGSZ6Jjw4Ppg8UgrlKvkfW8U6tM/mj1odGkl7ofSuwUQ51+xJZgQLt5QiUJMjp
X9mVM1DWhbOw5GqcSU7Pg7L0w6LwsUTwiWEMOMU7WYudCbm/xptRgkARp8hPNiUZ
To+wgMl2TfYYl6D2fqjeuFG18KLkd6Sdg2//ld0cwvYYqaOZIHRHU3Pe1+q4zaAf
J/6obgSZB06A1KghgfejIVQcIo6bZCtc6jkOpfTwmEmiBEpkUFPoxo/a3nNWrIja
jxW4Hev4AYtEe1SJ5svQ4gyBWiYBx/8xlUfad1oXZDeRWEpyWNe4rIqyKnutS82s
ffUTKuKMmnGTgNpSWWCoc9sCKutUcrLrM7PB0OYQeGTu2Jw8peS4+KBUcxFHEeJF
Arsf3EncxVx0GvEU+0FNQcJexmPTS/YoSDs4HPfi9ZLbQht7JKqd5Y5Zif5OQFhj
pn+29/8NJbhm83mOVNQllgRYLC6jzPnGhzlxSy4Tm6ECsoGF/6heA8mQlyKeOJSf
91i3C1QPN0Sn3K11+d3taxMRJICnVnnpbb+J0652eIoXABVPRZPJ4p+dGOJFryVp
9uB4hvD//gaWqzI1IdtrkXKWa7gBbLTIrz7pMLdIc7xLHeXpBky+3TZTPGmAAtQ0
pBsJaqvmOgrOui1ZyYNESCMt8MPP+fh3vMvbCAAO+TQJTDUWlwHN0JvPnb7KY/Nt
AbWZT4+pMuk4pjcPrCkgC6pVJydGzOj3BoHlP2cQMfBsYSKNzVt9zyt1OP7k+rz/
QclI2cOYeQYjJ9dScu8LETB9JPtUZdE1a0gJx3zSbblR90X+wZqQQmIUV/dzh0pU
FxWOk+OpULVawzGj30Ylpq99hs2p10R3vK91ZF8ctYqhUb2wpfN+Xl3Cqlo7tmWr
wnHbqaMCC9+/84fJ3bcrl0AUHVSqcAoylbjL6rijBtATMUAc6ZyU0WY4BEoyocKd
e+yeuMSEH03jL/XM9StS723b5R4QdifDCv2K4kNZizM5TkzcbXBs/c5GKlYbdZuA
dB7L1k+5vTUMwIvp06V8N+UI/Rufs+hJWf+7jRQ2ySru09uEkpYWUrR6egxdzHIR
CIuecn8T+/baCADYLyW6iR9i+0d9Uyw3AsaaAs1QMQCilZMXE6yk3c4PgReCgpvn
PPE/e16ob5lopXM30XUaiIAR4r4W4eAmgzw3/aluiFX9e7mRauWfreMKWuiuYkZM
aljsbZmf7WsjEmMw8J/FJk3DjLeMmBy3MvEfBdBwSPLxNw0lkh+Z4CYeB9gPfwpC
JwEF+mx9JigI3rMlHOJaRs0Ar5e3yoEriMJ4yksEPe9Jeqjc6ifNmpzmoJ/t1Sp2
UlxWmPGcei47TkvGdimx+aVYRzoHf7yefIENiJDlHMpG64avjXGGkvoV2Xj5JiUa
zZUIfMajcJDHw18OWTnT2gJAyOg+lAxndx8pYQAQhlOakfOuRMIh3OddJpaZCRuF
4YiIxN0apcZHjqmtYUP7mGbik530I1Di11MOYX5KYEEYeh5DxYilaGnTjz8J8ePp
a3oNR9f39MIOfNGq3IPbW8GAY6F8ifXU4bdV8g8zpmLdgbCUoP0eIroDYn+P1Du8
sYxCo/s4hzQ5HtIlI+7iJ/JkbnLOsKPCy2tRuptXe5vH35hqJaimYCELOK8jXoHq
iQAOTuXTYWNlkv8UdfjoCfgK1077ysZ+LXErGATBurywAybjbHBKv8XezB9nwbwL
jC85QX0BbEKhMqLWfuieb2VJbNjO8MM3lMMsirRo90Tw5w5l9t6rVCtji0o02Z2/
T4sZMx++1pUnk08+kDze9wYN74aVm/QI3d7p/CVQYqR3Vu2AfN3wmDTz/Rj2NhAR
GomJKQ8O2q2FPpFKsZF51GwHETbYTreNw3rgTpZY3u3wcHNAzBgR5LQzi8YlhYDm
EHgI4gBa/CTbtmoZ5ms32lNCNfYcpef82i8H7CeAt3iWU6av3z99796jYVn0qrH7
e+a+ko52Qx/r/YPAfUuyyZJ67Blhtez6SnejSReM3IuNlQjXuDnTE89mvUNiiGol
Mj91gy+06DXJfIDKyfbgdcWZZW1uKCkt0Edf/xeq+QsUUdwGbNeiHr8dOV2tXpfN
tAFxTR9nYRiR40jQvuDZjVKRhzO8jNJNWZ3QW6o55HVw9ZaC87ZZ5Hid3EwstBwT
/bJCFC+KhdQ1f7RO2tDG6OBzzaF9v86GOlk+M6N6M7sNP94YHQRYAPX+WW8NMKk9
KINnj3fi8fQR69+vRYfWVMWMdD9s3I9C+OFPoUWZ5THzopaOKt/yynJEjAeixhBk
P08l5PcwzTBgaegJPlc9v+uV1LQ418crWOjcoc4CXzZ7r1fxdm9O73X0av35cJLE
gK+/us0DihuO6VqhA0w7HnrPJysruNDxh2vLyVJJUOHURqjkHP1XwR68TIrlrzA7
4kVFd+MLeS2tqJhnPJtEeG6tjv9Cnm2np+8W56xYUl4JT4TIAvr9tfoY+7Fdok2r
YXM++n1Y00+WThtLZIcQV4hrin9svXO4atr13vq2pS4j+IkBUSa6od8JD54P8tQG
PcZOOMgwI5g5Tk+52JuDRuJBInKI49zYbB6x5J7wb62+RUfLZC9eTl0MiC7Vfoq1
IIyJIXfntHl3jJcH+/CCBvtQPBFUXSGSJUcoMdrDEvg+l6aYzhvtdVL7G7jKRZU1
HTybdmwfYAKO+3sRzjmDoQUMDc48P30LJ8fmso7E6V8KWaH1otHRmLtH/dpqtaFl
Gnx0rGBoAATe8HXgSk8Yvcgw5Qk2sP1Ym8uAwohSjfXfettGD5kFkZ8EbYtnNwAO
CLcZYzljOf5IEFyjlcfWSXEsmMTxReIqiVX/fLPt0ILlQJTSoZjSyJE044wzudqa
NrIJ2pD26TVR3yseSmkJWQ0uFm7DN1ySDe/KpSkcyu5dIxdfRJPcm95quQSA1/km
V8k7ckQoykGJLC2U3Gou3LfOAfx6hB/mvsfT0LcizMR5QKi+fV8yrf+nzuB6IzXT
jlBnG7B90hcQbKNcHY1euKaZQcB602B/Tog3N1HBRjatHRdOC/O1uXNxdabEx+xH
UcWNJ+1vqmmuME93Rv2GDPrzclGarqSC6rz46OrtEy1nB8D7aCZ1CTyCjNut4pix
T0Kveh/T8HjGWIVccPahtm+tXUTofu67etyYehcplz5F+W2ZS5S/Vrg9NuTZzC9Q
I1p8DNTDi5NuPGRtq5c+NKfykO5HRfESBQ0sDK8gxhn/pIH9piL13NWbvBessE1k
EZAV0GL0880VKoWkYkKqpT4fOjO/BoniK/6XPhTKCtvUUCLJNgt2LlyE7ZZdPijr
kMSrlqt71HK2DCn3BNicAavbPun5N9ogd/QjwQZY57E/z8jfLpMNAz7OyFJVvrs7
KZ0XG1ibzOw9RmLuiSfToZg7Xu9k5IZCb5Xt+qQ+A0L842anQi1sAcToZX3/HKfO
ueZS3F9T1yV9PJeqYbgS3/s6NbsjBUmS1s8/jF5mqkM8sl40fTfcdqZcMt3Hw0o/
iLuwO0yxgjF7rzhxUjCdC05pT/25cTpGLMv/PaBDvSJnZA+hCupZdyg1/RKzYaIN
bEiBF19Ppj6iur+P/nZS/5P03w4Pio2utUg0ev3I5FwxzGg1s93IDQKyAISz93Ah
IDqrEEuD7rx5kME6p/QeKGukuH4D9UYjgjibOGc8lFA4v2Hc7sDaPX+o2Wug12jk
+VxffnzSqdsoqrjJ//NaiYONHl5odv7C0bE7LYJHYpJvvx1ADHRJ+kFCdohYURL/
BwEAvy3S5yAqTwioAq9o/pER/jxEgQi6bvSnvmG9/po+KRpqHEo6Ssk+WKWF5yB2
tWUW49xRHieTnJaB+3skHwYiq5LQ97Rt935x93REeeMF8HfZZXsFDWrsO4lPSo4F
ZiRUdCJCE1KohxUTuQ8TklBxlw4Rf7/L7TEcN2/Fzhi+r0Ws+dyeVoP5mW9QJx6h
ohzcxtsHrAN8GF/LU5ju+GG5MxMY10wJwiZL9eUuopU83aA59WlBB3Bng+xUsYMC
vqiFbI7mQW0ePngicKXIH+zO4QM5mXiDbTMjNoFprStpKRLWqk2pFAsr89kMyIYu
corbt8g9dgxvl+ywaGo43wI+JTajpub0IbLrEOieXb58ziqWJELPkCVU3+QDk31/
sdqNfF6NArFoPQJkD2mmTXa5b5LbNCZaqRYKJmnThmgPDKR7+0yADjmF/6LVSahv
l9JQdV3h61n3JK1nof2qv33JGeAO5nUO3goA9iTuF2ZH9BvJski+7d4R3tazsfHA
/EBg8eCl5X9rSwWGCWPQEhtW9cDkPwjvFNwFgv10Ko09UV2TkHPGjU7Qd0si6Fpe
pc7ScWKEr66Dkjx5dYnz+S+Yvu9DvaQW3574aXmynyJ22SgSLifjxRWfQF+yk/lU
BvA0LZJYmGXslR10yO8/7OASPU5PBURC7O937PAdldP81BF7CFQdendA0M/ylNee
GyizjapJVzPBeRe8unOOkBALt5QkKV/EnpIQ/kbyWcMP8r4mqzF1wdRyyIaHNwoL
uf+MjMp2xc+iXiOaKEGCIuZYokKrfeVtgMXrucz62hzN+jNQXUEXWYt4yhmRnd7y
Mp4JGw2xBYII5Nu8Fg0spsyWlgUWeTxunBpiEwGgJ7wRUmLXt6ISMRHUZqXLMcxG
O9CmJ1UPeCymhMTEXJShQ3pdLrJ/u+biNETn6XKm/szQ3wqWpOrGnZIKvXhZt5Yt
pMhYSyhetfVPUrD4eIeJcb3LiiEhwOh/YXcAf1T6mRKc2gk2GkTaJx1Qwn0x0PcT
0Rsl7V4LZ1tIahps3pxqwWmTytOFcuPcSfmJesNku2UbTfHDEwS6lZgtvVeO6DA6
KLbLodzPQaMcdodRvvRYhc8vNCqhnegtYO2FZyVBiOXyS1S2cxxMZybrhjvohpv7
zAASV7o3NgPAVhC2BOrV6H5FArFzzYEkLheQu5lokOJBzJ2gFZsPd6VOG75kiXE3
FMNJBGeTsTRZuT42KLHMW3V5bA6HXan458mVfgs0n7B8tYan0bRhZL4lK1Zl1EH+
hfFq4R4W6oSdGBPJ+Ae8FWOWQ7W7uGvNYizObpMATgQw1PFqxZXI7VnwTNp5feLN
1iBS/6F09vFo6liINedUFYI3wuk9jC/CCrH4og5LCOdxcDrFp1LN1O/tQd8pQDlG
MHTmT4txHFzIb2U5luNHIV1tp0vYRss62QmcYYfg96lTFDCboGiaOPt65hXjqMdF
6SP0RIR8VEw2o/8lyf03EVIUTYMSAny/e52XK3P2FdA+Zp+k6vEM5YzfmqIVgQZB
5/7HMxSwgMzaQK5DEyYhCvXbFI6a2/YzQTLlU/cEZePvkQgLd2l+om/nk+yhgqdK
82D1wqQjCKHBlN2CG1+5x6FHqBAUtaND6VoQwoneCSglh/9uSpzMMm/XP+PEZGhz
x3VLqIKNsNI5qP+PSAKcIORzqz9NnNVIEUwU1lEJujmKQ9V8mAIQT7YlTszIEyOY
OHMy0TtlwSUEqZnGKKiPiHRKWG2LXESkcgTAkErLjzDvcXLd3OWiJTETARkagIpT
QWpaw/+l6F7EoZ1NRTJDpC74C5xkvGfLJ3oDb+MZQtVPQ0zhcoB5bjgz67k+dMII
3BbijxA8NL8aOQEQ8ZAayLvNwWmICfXvagZydNFBGBy+5NRIgJiF/uMuIpDwFEX9
IvefgRT40nsiKCp6kTMNmvMH88SD8cpcRemzuSIsz3kyMm8gse+LRGzC9AzniAlK
wAL78ir7U/Wo4iDTwww9vg6a6M1KsQF184idFH8aGCD2PWyrQcMjmvwmvSfdIX67
DokdjCO4NSX+pjEu0XVwWoe9tPzsjB01TmcSbBeuiTQ8MUhA0KjdrW+jUYfkCyDZ
gzzKpyDdiK6jcWN5tYkn4l8GxgCkktZ5EOdNiVm5ybRCWXQubFNhTcKtlOe+lwz2
YOGWnTxljs2dYZHERRUkAsakSc95zEH6FUwJiKpL2uqnNqsyHuPYquUTbnxENpl5
j7bSVzKHUFGRaGOiPJEXNCzHGCGvra3lzkI1dFMwaYhMyx1+FI71VsQnm5CdHykv
43fDaquI56IPhdQ1sg+x97i7WqpA4/s3Qky4DsCclymquqMKeepPW2H1a69AO0mb
OoeqI3QruNZR5dSy26eLGnSVPau5WctcY6aOEsPOSby3mK2C0mUSfGmmtqhb+Y2M
igLpgbMc27DxO5acWqZHQfC0MZvp4OAA3J/dweKRUXw1VXffnHMQ3mN3yHutLydE
tmR6bPMYRFsvqLmu8x+hpsO4xbEefXXE/mUXkCvGpcjZ7lCFKGACNkwMd6HEbY+V
4NXaspEU3cpDD2RYX2OHE5cpfbNYCW69P7kS8UawcLjT90PqLZ5Qf6RVfx05NpON
Js37N/OLWWDm3OV5/0OjGRs3qSF4p0eyF0iZ2/vaIyJzhodJRcdofPeWfeMi7IpL
6gdJZuIOIAFspzJgty7G7lCq3Vvi/tn2zP9fyJ784YhqNagPEn4wh1bCJLZgcoBE
afU2HLDAFb8xNcj5b6kRs+qDyWDor/H7REZP/059e11tE9Sei/gdmhnYlaFMQvS4
w+OJdt/TmwhjrnfMjI0LaS2w5TsTsntV6m/TXeHJ091xpBR1oOKEW4RRVPFU/UI9
bUbZ84TDPnQC+Frbfd5PhQ9xVpkDqmTwPA1DwuEGS8Vg20QbAOP+oTxGf+VzvkEu
Alaw7EF5bFPK1ZRSZa/3M7gX55yZjLyrTNBrvcstCvnbOzUokIffjvnLKuBfKCrw
pWv730HXjeovv9/ro3ozSiy38fnGMZ8HGcOdzdG77OWPGfVX+nIRe71uPo/F1Eco
PQirheKDmyuCX6KheiSdUtpC20SpgXJa1KbApb0T0kNQy2I0/QXdlulmk4+aaPll
rPxj7I5xUZrzPK+yC7jvC5p+Nx2etSAT7pNH1qYfuLiTp00TfGzyIIlKjv5MvOjs
UR6718QA3RBymmgEjHgF9klwP56kUff9bz3dWpiR4iW24vPufL07fjmbopQYp7/a
iM5zOy6XWaqjW2mM/8QX9hvdeKN7Kokb4AG2UR3WyU0cBHMhPjpK+zW+cAtZWjZs
Rbgl6cTmJnuDgNz5kz6GRYlLnI5tUC0rnma+gkqY5cPZOd5BxgZb0OBIGSRTsxqR
iSKLRRql+FYPyvJ0Mr9egGlxizYS50lHHkz6HfFBVPMMGfTK56haeRjI6/cpRZUG
v0X5ad/jcM4jdPnNIPm16U3/1cf9ANXhuLGIhOf1AnKSFQXjzG1cqxxd5Y611168
9qnE5FgGbT/CuBVPYu+m0svnP4hm2d3rd2UtjlCpqGGh0sd2XxDCBoUCrTBFUY8o
GWhPvkyEAu+RCedwsg008wuZepbsRtd7z+CKCFXMPPoKox3EfWZd3tkz2ieSQF5D
WJUDuAp7umMLuTM9TBligrYtL67FXKVBCWahk6taJcLx6ekXotAmdjI0OQuzG5rn
l0vFWHsHo5ALJofwKx0pVeqlKdLrUFE1SE3R71ReJcojRppyEDKz8dTj9ZkFRY7p
ZOhJQIjqO32KpmAKWYHQCkGJQmbmDJV96zZXYpdT7fTX9xHftpS3DdmhTexOfbEB
wqELy7ygv/hV4yc0dsAMm7DyJMwFHwMLeE2HhrV036sI5DNZdYOxBze/uplkV2X0
ILs1i1Ok2ivel7DROPvieLgC8r60IQi5yBfjEsuHGicMh4JXiaBnYXhqB9FUrTUa
3ATDTXWeIGzFrwC87duxOPhBcQo3/W2z1pTL8JYZHpv+4CQt7VMdDqLFo8ynO2vR
xEg6yR1zQaJzuUHzUFfO7IXHriP0rUfb6CWNIE+13CQ2RGZcM6znoXTjww/a4nnU
pEUN3GdueSlguRMNJjAvKg/5yDJyqHvJzsMggyHAYiHMUKWpWJi6lDBYvIjTmHcp
O/PKg3FjDBHT2iVJXifNpMph+tT1srXFVhQ0nO9rymbwhLIAWSshXmK9+s9kpS2w
TpZtZnIHAboO3h3irRLBp2C57Vm7+gK/vwTUebRMKOIAIn72lQ/QTV5YiYFcYNBM
FcntmTNKGkqKOdv14k9736IsmH5iJyncn+ov6mrRFJxgOO6dhfW1MVRBgL4IECnm
r4hCtpWX+fmnQmklRnW9AHSirz1LU+Y6adiGoZtET5W0sE0uCX6yWi9TSgmKEFcf
f6DOErMFd5N3YmGRJ//dQbBlBCoSmPnubWL5Y3KNbFDa0XQu9n8VLoUM8Xbh4vdb
KnH/a4G+k5AFxiTQRUd/a5b9dYFLjO5xk6pbSK7m+tEPDkHmFiCVbXqdQFqkWVgT
7jpJVPc2lN5d0FaRu2/O4uKd2AGymdtA9/Ub5z4X5KxSpHll1lihwupEvPcgS1wf
a/K22zR3YVknfbysxaZN2aSu8BHwjVbO3GgD2gp9832jxO99nT3k5m9WtbrPRgC1
owzFbLnpbJ7f2+ZmNVu/t/1jOR4gsgkzRVizPOQ1L0h0TaunkL9KR67Kbyzmo3Cg
9LFQypGwduJkuC5fX/iBpXx6CEkyTwE3wi11zJ/iE+tMhrXjUZGgwwjJvWhZSm1A
g1lfEYfGMSAbZFsmdymRc0nfWzSYtUNRXe6xI+4W9xOUIOw4KdCpTuEb+4/dqwYs
vn6BPown9ojpYvLPAy7IVIneVTD6hvZ0jfNhavfk5xnXNKy7VHKBqPWCZn+Hdgon
e3VYEok5bChdaVg7JnPyIwAIKFiMDADY7SNZaGOmMntWOEAIb/Bgv8gi7yLMgntP
lbBbE7Edt4yijJuKrPNkFTzpmwNkw09GCg/EgfVfFHVDk8NWpRfQtfTm7RKhndPV
tvBKQRsA3TAW5x1ty0Ie1teo5h+mID++2ynYUaueICOjmiTJWL7HxOtwx90hsmwE
1AL5DYMAQUOM/UR4yu2T0zvExbRMh4uka5tCmfLM46qE9yZJ97skfk7jfm/FAaug
Dyiu/oqMCE+Ik4O1DAo2sqEJFoVCyr1DFJOEmwA0eHEmdEJivcYcMJ7u5Z7Jqeyb
723mCpdnLuOSvwFZ3fKuI5Vjs9UAT675CEw4zE1ITjVksJlxUaFUha/IaUagjxU7
EJSr8tFLF3oXHOPl4MPNkg7AeiHI+E1RosweSZYB+udICODKv0hgOdmNPRDmZ1ao
cJmy5DzAnrbl658WSBmInipJWWQmQqNziFapYgoe14rSRQ6zgd2as85eaqPe3maQ
2Yeg5Ul0gyFKqZMvij6YdV9a9sEusKeXEnLSGaPORoy9x3pMxTTq1zvxEF2cmpPu
5V3md+3WsymWCOEJZTXfN7cCfhl4MKufN6JXoW8j3X7uH5FaD0nJLna3h6R86W2d
Ib2ea7TJc+LgZmD0oZ+HGjyOw/TjFpl1LZqWoukTIVF5dVBK1N1EM2AZu8IAZ0Zm
qyDildPeuyhwrSvMAb30NwXoT44ac73ihCMCmYvbGipk1gnJRc/A5ba5o/FU7VAZ
9HEhFVa40otMQ7eF1vMmpFFNRYwHnc1jkoiUVrBVj7Yu7Cz2S9kItn0cgTEMf5S8
o+tCIwPFNzySwc/9u/oIwpV6199saznhVllRxsJ7SNO72sxMH4IhgAr5dkN9/0XQ
QlldpGjTrJQj+Rf3RfQarkoPrCA+VHYcGK0/tLPGSMKCqL48kohVCPTpRxELt5sH
/Bybf/5hw2oNcygV6TfyMN/fstdo5ldM3rPeI0SxBqbFf7A7mAtIuTJ6FvxU+dlq
zinAL7kbvZ7B2Cjud201jBOiLPuCHa7Trs/kvErPGQh15pLWTyl4TVnPgkgBHhYr
8XiHKcBWBfYL+dPLaEujbeBup815lVIUOyzht6Z8oNEpQtjZPkA+WjBUsTUBQkUA
dEJg6Ty57Si7e+aHkRp86MQmFDO6cJmJiNmVK9BAsED2z4fDGoh2Oeo7fOJDQ1QH
T99iCQthYWytSShL8HEzCMctDexDyNXSHVn5a96YJTY9wc3YG70Mph551vMDWWE2
pCfa1h+HTE5TZjqURotmRtrH0eyK1qIynvcdZmQw6JdiDqkBi5Jfc94g0vtTUZYV
q+sbN3ZeCMKiQHamjA7pekuQWEaf15J3PbxaOrwfZfWs9rf1GQZyB/Q52ktHTB1V
p5VgUrFEP+wMGWSLtBsI1t2+L9Engj1993KVDRl28HWDYzeTDEkgjipPxO/yJnPN
pmnnO1GECUVl2A9aZ2mb4VTsgvMRfVEnDfV5on+dEqSGTbIwLfwmi8Bp4oiDkG2h
+QYmVDHhSEACJ+vxFb1aZlSO6jUs/MmswUeemZKKl0R95jQEiftOyfoZeozYHCKB
xxtw6D0FpOcEe6Mys+lozavvbEOfroEGSQ+wngMvoz2IYvm0DscITrL+yxeQ+etY
XKJRyz8sX3fdYb6Jt5XzTaJqOcSqO8Fho/Y82IceSk0To1dDUKJ5zS21Rnj6viq2
Zd2wnAIvLD6DsJ7m6NL4IZwnkQOv4zTZ2CHfqszXQxNFmlJP2eFiTCbFGu0Vr83o
X5V/wTV1wWQ0KhghzrrOCkNd6hwN63meBzxMDmuEKzKA566rMdx/iVER59e+wcSv
j4VXKSKMADM8DUFO8STecKpszF7QgYLIX3W2PhcoR+ivoUdTglA/9R1EVmQlHQt6
CH9v7rRa4+7VDYXKKSBDXIgj5DpkZfoO+b3Vkp4IIV+rP4oqTuCd0KpKWZpiNQng
QvBl4QGS8eDJ2VIfhSUONVBDd0LK0m5g7YAzySE/ap7L20sh7IOrhEjmXIWhgn9z
/OLpxpL7aSF0YDstFtu6NjVs69tuLn87GffGHbH0DPZu8SYPDYmI8gHW9u5gFLyf
evOGsfOMmEYprasZcOJKzbRPGgpJktoDva39iRcioqSaz3SONnicCiOZuMa8k+HK
pkb+3RW7XCh747FS19suiDseyhATVrlNih30IHZiRkk2POPEhcxa/K9Lp3156i6B
i8GdnK9oqiE+320oGqBtKVuXY5ysOFgLzM/QdfdkXdOu+JZ9zCiXSwnIVvdiKhIF
DYaPANJVN9W7tR30BGgJtUYpwDBLXEV30uw6DEWHq+CXXSiFDk4Zh61DPD6vnPdt
affJY0mjFnvcFfKKcHltNKELNizw+l75IUyNWjPGmCoCKv9tAulvAmtLZ3HNG7VH
fz7rt+c4cJsHS2PciK1x8mIN7GkwJntjyf/MNdQ9tgtLk52Ior7TWWpn41yZK66Z
J0gvfIGcsfiiTN0dyScgzSIKEGdvBOOUeAPuvKoIZSaV3I9x+BeY059TdUIRsMvz
Ga/5Tom52IJD1tZQ593/vOhLCfhjhp4x9p1JjC2+M6OlQS7e4J6s43wWZ99gSy0M
OfFZW+vnDLeHWW5hVTnSfWlSdRI58dANiiAWBnQakfyn7BHVCiNofwhQnH9YHA56
ex/tsdJLnwRKXzT1Vvf3X9KcBxknF+TCVGnGOEajWoFFQBMZlA9E4U5U7RcApV0P
zlrZLj0S+KDGRHNisFVDwbItRcYT32ixe+Pc9o+/tibmdduIyTPEO/2H5BEVGCiS
9HX0ANCK0L+87GKxmqBDRORz37oTZBHlSnyPOEnER7KJnh2Eun1nP/zC+WrmgF/l
cdSCpMD3NB1F67ikZOPFKexlQMs+f4eAKrID92BrviVefV7CGBNNSt6uCc2CtgCy
l/5GA+Fq/6wR/Bbc9M1WEtevKX5nz/0xsw20Hod1xr1/pvAyUjxhmzuk2ZdGd7ct
gswLupL2DtnvFMc7Uc13fCxA8VUvJEKTyb+Zy4cY/CKPpkfDxD5/mPibV1uayuxD
M1aYHPALqNcNIQgBzFfrIzbN9bDZlrsd8/ZzYdBfifAaoJYPQgBX6hBVFFr4W1lk
Ly3VjiqioH/8q/SbZlKqu+fd1WpKPA6f6BH2gJVFe/9u3+2pfB9IKwQ6SEctUkkK
YTSeg3Tw+HZWEYjo3KbS/LRysSTLoP36WviWCII066KFlzM+U8QwG2bQiTlyxlIi
cLZP/yJ7dn5VEwuISe8mx3wCEM80OuMrFErL7zb2C/aq67B6/v92ez0rlrVkzuuT
2edq77hr2mQy9ch/oZu8OORix3nZgheWpe15UQQDdevT4g72BVve/+H5jNPEoZgb
jx7UcLrIU3XsTaFyCENyXrMYkmzp2TFXgYch3m+8D2lTYzmRr+sSd8KulGoRwdUF
9fs763p9Qawt8AKBI+A7ogzw15OGfq0QbiDQO2ohqAloO8KE9Xjax16ACc2n5sCC
QCMDSwaZCvI9CPc0AO+WWRzxa274ZNU7fTRuIYGQKeutnYYxZ6at26lBf1qcYw6r
usCiSXVk1J9fxfH0mCeNgZvS6fj5Vb5AzdHoVx5aZ8/k5nZW3sVl30fim4QeZe8P
oscyfz494stPLT5h397E2uPFHVpGJlrSy1agiYq345aWI1oTKDJXvlkGdSu7cg0u
AvfPyquiGL+PkFYVNDuQRQY9ssLLFcftIcDEoWENz5PZ4Z1Xy+asv4TsMlbTiQaO
ocuWFSy2ECEvzKN8NO11QGOQiLp7Efqy/t9LlywPlW3x9pPEziTJK6eJcBrIIxm2
i6GwuBRhkn0evt141GU2taf6yYUYsuLE5PUwUHn33UkqsfEKD6rhLGlcT6EkQRtJ
yK7iYD3p0XfdWU26kWZtkfriseJjR7I2QyuM6Oqxu6z5JmB3r79rxjHdJDrwqirv
O4keAjr7itK4J4yhlD1YStcP12kGRc1HslLTgQyhkvutoDwTgZI+0wBCGwEM22KM
ptA6ycCXaFD3xpw3oc4wkxKLY5Vj1zF7UBB6Wqu2SQHprp0UmnOAZlWXDopvX6TC
mdZ+Mm/02EyqR9GJRG4fUwtcYa5zDqq7ynVuGrG2Z4ATutjXidtlDNr/CK31Ed7l
QCbNIDrjK9xhIXRW7UKx0bn9M0EcQEM37rkAo3Hu9H1pouiGJWmIxYimuTZbXylx
2WOgN1ltvP6Q8TS6kPOVVlNJyghNmJwE7y+3pODlqkXssRtJ/VvHPX436STOhEbK
VJk5MLiixX/uW0vVTJG0nvyJX0uu2jiHHWPcbJdL4tfCxCK1omOEeYHNC/8acLmd
az3jm8qzLCxlaFw/eH4fQ5DDMr+4lTCJAR+o2IOYMq+z/TZM1UhRc73U/T9tkBjM
9ohWuMHlvRVkQ1iFGHf6t9KQE72o1Hp40kawqOhUL+L5oaI8P8Chts1fBuCWOxV7
V/T7Vrhb/GJIA6EW8esb2OqxDFbwwnwqYod+6B8mnkFzU7Qcv5Bp7W8ax7gNZypF
mpV1/WGExcTdZiM3yq/5iYjijr1mSajH4AGoDp5VZ3i8lyc6lJ1QDGL7bCwSDHk1
/pnKc5r2Y2n7B6TsnxzGmihURDWcrPS46Ic2BtRAzNiLVz+TEa8Y5s9QqCVw3YDe
X8BUnsOs+vkuYTpR0PWr+IuWDca1pgJAZMAEJtzJyvZbnR0vg3f6cQ+2MwmjvhDL
mxGaEGEbFqS2+68yBPDP/lQ6pyEiW491zFyxP9PwMzsEpCUouO12VrfAgosRQa53
H3kHNtwUbBtHx7ZzDGqew5f2kus7vIBmQ6N8Xu3li9Aab7OGmaVRZ6nvd8WJ1694
CZ7LHFBrnksatECFrj7MCgqbreUYFG8rJT17vCikFPtmNbSt/x34pON1VtChPN+s
khKYnfXOQ78+ndSFxZEJ3Zs4En5vhtGLTp6kSsioORAsvEYWAQf5JqKhI38qZwx4
dE7NOtuSDp6DglCOTTKDZwMyhdr8KTpWgd2DirxT1ZumXC+07YV5xCeGI/qKDrb+
G3LzNxOEHr+cCVaYlkQWkl5+U4rapWA1wKAceqkL8LTyXXkz3VOzhgE3eSh/exg7
dh4CBATDBF0aWdiTxBy3Vs3d8p8DXeyBh5CHQgAg/vlHpgeQHUI43wGInjRDHh7w
V+EK5qoKsCTzAqTVo+h753bz/JpjoHmyT6d7Kp36vqasnMr34vglvvCkaXrAH+ln
wJdfpLw3A40PPXfmtZskjRAeOX7ZVBoNBP5bSsTTJR91Q8hACd5Dbt7OdmXr0XPs
HtCu5zzS9NXij/Grq74K1WjRV0kXrQQ0H3enT9yZYr6BqCsUbpZpFQqZ1lTpaW54
6aBsNgbrsPWXkha9l/nib+5vlOBlz9G62Wve8e6uHIMW0gIkDwUCnLK2gYC+m4L6
wDnkct7OTCwb+p6Jdyf2KkhnnB1r2+Cmi+oVbwxbqWBxd72zxFXcJvZni/Np2+Zp
8R4hMdemdSKT/ajSo+a2j+bd2B9rm4OAHkU3dmvfZPsWdMUKzPOfWg0PABXJmNyc
xM95IBJTMVOmMGfRIYq/U4tM7/RhN0uK9yqSQZwegenbG2pXArxw3D1FLoIi6/cY
6R2o+xQkXpXqDmb40HK33wbaIyxN2EbKSk3m7NrlmAuQRE8t5CZE7gdkYKjeAr/c
B9K5JkjEKYOaOyz3msHmzd2XD9ZZoxN1Kkg3O2c+CsGeWh7PBmt+ujQyijsJ5Ud+
Gc5EDVcnE8HEAFjxDPDN2PeiStZzOS2KNS410m6tKxgIaMskegP5RpSTQKrd/BwE
Zw3zV1igBHR+f6pFIjGM4Ls3ng6yJiqaK1rwtj09jzBRt0IMpYBlXyINczp7ZupV
znFIEXb6ghF+EJEDdCzH9g7OX9IOd0vF7bezFyIMcfk6SPplEFMToy9qcNUgcPTu
GLUwxKdbazSv41CoJJT4Lzuo/vrO1xsxihFhAemnG+fGgv6YsZ3rApfACIxQAAT8
rphqhhGRU2yixxwnyNVas8J1O3rFmTL/AsWLRYSToBmKIKniWwbMCTod1z6mXlBm
+KwqqWkxhOt+7t1h8gYMljhL8bx9mfkV05cDok8LWSzTztFxjNGmgktKqdOv/jpq
lU0MroYS91sHnFrtR9ttTusMIwQQTAHoKJUHl9vKnEgFDWxDoCR7PC8gXSlW0ygH
FLvWSLTV23p+89AsXnPzLLvO/sHA8ZBhQsPraDj2Mk3PS02iTgK8rnVkfTsmTEXV
MY3DwxbsTcPPhqA/w4uGXpAlUyR0Owe9qpgpL1dTd3SPPXvQlJ8kR1dJ0TEb0WU9
xXMtCc+jrWqRBC6j0tdbLNY41pjscbNQwCwJQi/zeiavUC8jZLano1BG2QI7pMzW
XH/TejQDlbSOV8JWQVhvBvvfchUWwNZayIjXhJr7eV+j7FvG1TLh34o1KG6TMDn+
XDLYDjitxjCOkJvT/vKvuMwSB5ziKm8hMS9IP2se8z4hMa5h5MaYZ07mwZKXdjR6
IQt1b5u97nIOexksk9cN5ZJ+V8M3lFOIbtheK+i9cPYSQYgl8yJmvH1FyQAjHq02
fTI7D1A8UqqlXHU9Jmr/Fu+Bs/aUYYS6p1aMLyqXIc1KdNlnKWeaZGzLIeoAukRT
qCjTqVjqXi2d6L7GUp8OHiOBXLYbreLMURejMAlRlCtiYUuJ/sLrkp9CuFsDvlDW
1E/t1nKLZLU3qyKAM2tl2SEsN3MJX0OUQSEoNWXyP6eiSDoHsgP1BXhf6/2qlxaR
vFskn+wO2LL3aTeSaUKpsiLzRW1LaZ8lGZub6XL1L8LaU3rzC59oJaajIXZw93Uw
LMyaCsnE4ZpTBosYPchlcx7nfGRZjQV9xX6fFyW2CfmAOES8cH+0DMPgDMXiyNOJ
jxCfXHVe0LDH4/VDj1R6QB0XWTTxDOr9wctfh0OFtjyGipKsAzW548tZBUuyIW+y
IIbOCJCTnWUt4y/f0Xc7RUBgaepDVjjwYQqOG5fiNgA/neUuaS2GkVD53lp8+jYV
KzF/rGME6DK81XW3Z/DbyNVW5oRxVA1KVsyH+FgWN0d0visawB+KqrRdMlCpfuyo
A7EvR9mN3vMc2QKii0ZW/oQReteAKEE1CcThAeVDIMUzFLr5eEMfvEBxME67SVjj
b68hj0IWZFSNu6dg9A37+WGXKkdtMXw6W0DIlSSo9D4bD03A8zfX7TLRiUbPP2/X
dsyz5gy3B6XY8mVWGTftyd3ZWXCPfsPOZThtSgesigmUV0u3m5iYMLKzQ7qMDOHo
7SomptakVHl+gMjeV8EZjaXHQ9S1OwoFXWYmr1GCLhk/auqfqU4JciUgIlxOP+Z+
wCSX2vPq5m3zQ3tbyvJU0IGmm70KPDixrXXrgniPSVNEiZqhM1ZqNJYLo9e69/3g
3oTkjrCyDCPDCgG1nVM6Yz+gELH7KaDg/aReYGhIoClX0OeGW10ACQ8TVKS/zfAC
BLbiDODNcPiTlBmg11ORR9FNQ+AVuJh0HJGrkrgxVGZ/8d7T9ldQN2ojog3+oxaV
/VZatUVj2qgHTktdOw1q4oe4qoN4TCBT50LIu2Tmlrvq6MFfeT/OnmXDEAdYPaYu
+6HmEmN3BYzkGMWbzR40naKBSRevp9Sxawqup3d/edGfs1dNjZy8cmp9RSvtVS5O
VG05G54lAM/wP9y9JlUUb1RDCv1tEgae1x/ztH1+w2fhztgecGPcjvlj5FgRwUvG
tcfUA81jx9057cnEQ1ZanX4sdZQgkTxlSrCsVPzcsNpfkoDeCyrjXNNclCvM19i1
Ji7WydAD+29GdPoHOJcV3yG1fowp9BrI+c8ocf1IczzwyrFbNBv18Fs4j8aRt2fN
+SPZdVqv1Qc2se6FuqLo+XAz4nxW1Vp2D2Czp2R2gRwRl7ZEgFRI0Y8B6fTxdYdp
GOwPtjYG/T64IY8VZor5RI34sr5WTypQ1RyLteDeipricfiSgeIWhWRleHsRDK+e
MMVC9s6//cqFLr7SkZwV3v/VUwZZzqMTpNDtHpzsORKwK29u6teMl/QXIfhmdde4
sEQeu1yPBsMUaItnLf8G9PCTL8nON0VA31llKbeeDvL4jA388A1BKh9Grrw7tcgG
uNodicKxfYHpN3j5SjO/NCcxU4S73TvSSX2X95cS9etNp1qrWLVFHWFrn7/btMbk
kCKnjYFr0wp6vfZfnfw9YT8SML2hLt8VbSPdcKLIFp+AYnbcwex1BOQ01r4WSLOm
TRtXtEklQAGiA0sO8OYhcq+Uck0z+beXIvwcc+jzKWCG/iLJmxLu2XVIMssUyXRv
EVUM9qKYXwU02tJ1IjT4Zj/mCe13LOarUMd7Mgene/f3gu9xGDjGHJzJwEcVM+d9
8bzgzZ0lLZt8+KGl9ZssWgv3FawY85i48GXZvPKysYpdassi+QC9JtNayZBiZIyi
T/ddXlNoLcPUv6iZTalidfbq04rQ5bcGxRHfy1347tX0OKrA4QmpWPm+fY4v3LJy
OO5FxOMM/S6zDOUJlvgfT/UsROVMG4bvCivwSSV50Un9xAAiHk+IvdCPFpWvwY8q
a+JZKHocBoYdzgbJdeH7KTt459h4Q9/eov/OwXOip2yhBM7CQQhk6oXAcdWHUZdW
IQzw9OmnnLqIe2D4MFQth92pZ+WGR7w6NpBgfX9gB5uCzZ7Rp/C/mfjXuoOsdEbC
2wTHWVwX3mEFlbOVnhQ9erl43Qa2n0vdwl0subyDXBd6m7rHDZWHwJoVBbzNGLhA
eezDHHd5+3Opz0+6elwyT2kgIkDPJqqyMteIAlHczmuF5Du0BHRvo8HbDrUh3b4Z
XrZpEro2HBWEtIpDhZU1tX7o2GtFo8HKEnPvWeTbBFnAO1hU4ja4+PCim93lJrV4
0jA8CoWRBcoEZBEW5T7ZDrGDH0//MiSN6nr89JbZ6uPguEtg14y1K/S73dkmonhY
CAMvJ4QoaKIRL6SQPSyK26DIi2tdZMUuDRUmqs6jAdMJEGECaguMb/lyvlGpcjGp
naTKsHKSV54G7TZJBYgL1uUn2c16atGdciNLQwmJ9koVfGNoijVKV8yILbhqYPG4
WiQkpFNJyTIEV9DwgxBqgseUsofrs9U5nuMXjyLaT8IHKQnV+hK3SdqGwJg47aLH
lsS8gz2aKGP29yNaJ0isknTgFzB9y7ZbFztnZzcoY5CBcVVDxAEcOpaKlQsmT/68
kzbMXLetdhC0AIrAyOqTjalXCOsxwCpqJSGNjtEOBuFadahIEfT8qwUJ/ZolTB1Z
p64HpSzKQnaVznCWdYqoExwTgx4jgE0klSURpmaNUjcvuxvAlor3FGWpMEth4Dva
YwwcjCGohTEG8KN+wQYrjfZdl5VsfHZZeDEhNwW9YhAEED50yl3Xwej/27c2DYVx
QTcCcZ79K51tNqgmQl0Qh15XU4jinCI4xacLp91JmJMOZ2tFlG2T0DrsCzXStllY
z1QYDVlmx/1/OKORiJlSJDcInzdCuZEZ3P8YVgQlEFx0yl9nTWgzoFLzEq8a8bpm
tXZRKJY4YiovMNtf28xCy8Cb5p/Ibe3BBhhUos8fZmZfECDLlSM9tnakvFEcwDsf
tTJvAByLxyItn7eEC0NBREDWzo+5Zbg72IBIYv6iafDl2DBVFB2ywqy35RpVbISo
+lVjPk1C7HvCxCX6ax/ZceNRM2MG7gEoItVpCrPC65XWP6IAZou19Y1uPMa7wSCY
L3Dh9wIty7jFKOsMXkZJ+GmggizevhM2Z1ddlgJ+Xy0ClFzq2Go5uv0LNUu7HXo3
i3YCCF3ltR0zNTgrEbnccJTLGqU1kNJfWeWzFTilENqgUbBgL5JhL+kh7arNuMQj
kTaJdI2yIAcJwLxcNhaz8rCf9PdUZWNcmRFbnxuevbY44xqiHV5+2STf/AyH3q3Q
Il4d77xK5LVz7NVUTzoEgu9iHC2tjALkzBeVVHk79iNU4mGVgsaafGcIBEfCixoL
ssXjhs0ox1Fbm3kbn0CZVmef38kf4M+ffh/smOM5Hbun3CpALp5PtypAJvF/NIQv
DvIYxdII4leXx0WJbdpwv4H1RBh2dd1SCGYKvzFARlF/q/YU/nhr+u+Q601tp0Km
7b1vooEeLii6ep4+h7azUFRSBtKkf9SLVDZcc772y3VBbt4msbBZ7O1R3u78V3W+
mwKF4Gqq7jeGKymAsRwVQV0IZ3fI1+5NVue3GWO+B+qsaJCF1h7z4PjgF9eab3WN
hoxSxwNBhLXWnHUoiiBX+zhtx8Zpv9jf43VI76zqgHEwYgJMSmbQmfOqXwyuOPLY
tHTNeZtZk14k/IQAs0D7Bz9gOmFPJyVIW0WGmiHfk8Mj4qs4LQSeDskD3raVjtNw
6lfoRU3Un4x4khYe5kbNp6YIn39IcL3nFv8H9hjhtlvBe38N1bN501cWtulAlUmL
byWIN5wlZv9po3RB0cZDVJwuwDhnXiGvHd89tDNqJnmw8SOlWLiy9ZD/z2QcKHGL
rDGpalU/g/rgy2ZdtBXb6NxRmzQ8AE+UMl4eh7lncgq+0eeqEXZgroId/KP1f73N
u8zsmtgYR1+rSvH7rdqDP+svgCSrF0vVzVsWPcT7j50XPvHc9S46lM4QOF4S/71J
ZxeVvvOZkMUwGcUyAtHeM7IAiKw6TSwunbaqH6Ea5kXiBlQV8u/epZfSbz1o5eT/
qAjEWZKK4KtQQ61MbQBOOHOIErt5azkInUoVOzS63JbzO3rf3ZbHDkaAEYyrH26i
8szt9qC/+467DhXbvPLX7MVWQo4bTJYO7hDk0f4ZlHvZxUtBXPcp6dn/NWJoRPPi
lQ8ihYzrFCM3/xKDUqr+pAOiz2K1ePIYfiajyS4NEZdWjoV5X2uvCzF1CtNidQSC
28kwZjGQ8HFXf2CbG8bY4Tn4t65i8RX+CHd/JHFhtRmLfTrNJuh1hCsJJYm8qhx5
VxLlggu6xmCbhvA/rfEHYYwMv2L5ZOkrszafUqP1EFb0h9hC15qKOUg4q38K47qK
C64a1KbRMd8WkKMBcgC2WtgHLIRrkPxEgtQbAB28QXBxCCXVnvu22utnfT2m3k5v
PeBOnT1K7Uy8sbd3z3hhvzBxA/kGaHHfBp/fnNEd1JqybDtkoUAkgDgEb5ycu+6W
6sByUdPjqfoRPsa25aemqo5XH1lDmJgZ3cwCpmwoAFPWyii6DV4p2Z3cGZdvNLjM
GwOpjmrJkHUOB1bOO/UkQpFEyHNB8+8K43h1wtT3RjWZrE+3XGFZczMKWpwmWEwk
UyrWhNL20F91ocqbygv7LQUkreRZxagj5pzisJtK6vshvSaIcDly2ycoMFKKU2fz
P951FpSWAnNNsIYvR5f6cm+xdQK3Nx44przH8D/axSHJkITbxRePffC0MMqNdfPS
gauuOq9MPJjlBMRI88XNiC2ApHpcWSMFgtF8+t2GfBjbFgJJWeaEQXx+Znub5OMQ
ZYgv9UQ2juabzjoSCAOii6rl8t6O5k//hs3p2QOwEI+RWBJ7Aa9XYkX6ctb2Iwu5
N9NBxCowZyK7TI1xtvZ5fgqVnDeVG2LHwJPbV1x5Sj+wAQzbhek1Mpx+yzi6j4FZ
ToIMAlQ4xNQ5VPeqmHLx/BpERJ6al29/pWy9aqQSJnRSoGUz0BVl+He/SOHT0uHg
AZFqVDED1tRKHjAcZgDKTV0UFOgb2jwaBySgbgai/hQslkFhflLM6WerIx5SDRSz
68BOlv6iUj3Ev53E7xz3ABUCQ7HSVUo+CHTAxBmMk23XTIJi5kdNBIwOi0CBS5vd
w03qBpIheEYgvYCpCf1D6jgaFfKOSv/MqHg7uZ+fCFEpXRRNUKamYCA8tyiQ41u/
d6ltceyZ+imjjYdLEJLsUZmvCpSP+QQW776gkMiRoiVVjVZFhmQm4krBxc1+C15R
gjQWP6/cQFAXt6p1s5ackpmFMOs2AeWPqSlznbX02X02P6MYvrOB40mNlAioautS
sc+oAmEQ9dVdBvBGpckR58XTEx/h5vU5o8+xw2VYBWNXsD4Z2lG/16w/I1jJEIF5
6RrqTEDFnOQTGgJaljzGXxq3lK4U87iIxrvfRPTntqJ1P3cWY5x5KMZz1LCERk11
FOIlZB+16XoHqoBt+Tyrx33GFH19yB52pWfppfQ80cOZNzx/wIeRR/XnPJj+LzJg
ZsqD0T+wIwEN/K7Us2DQgaCuyKkD4/c88aa+cmtqcHmJ5J1MgzspoAyHarOY+t2v
/+1kUzoJzYre1AgoMg22RxRKMkUqEb/SloW1WgK5PQa2KYzFkHVVY8dzE0KUiEYm
E2BflGOYxKz445VG3yEbBZwqBJirQ+Rd6zP458fjbiCJw7SOz7y40uGNNavjyUsw
NvcqE4TL4+4QF/xrijwKOoWa5dhZv5I6sS4/SJsNWckRde7JWQeag5+0wVrdmny7
e1oICZ8dh/40jTFtusHEGXqJGjASJ7+DWcqZ13TaNQMZX4n0fzj1zIH3fBbrV8sj
4sW382YjP6grD9ZMhRUYOMb6djehxpZzZxFfCwHaUFE8/kNdkI5to5r/3hj9Cc7U
Ob1eofKBhAfsAaJIr9SI1XucjrRcgg9z5VPxLMDriXZSpd9aJzX0y0X9/Xgnf4GF
fJ3zKmimIkJz6+QrLGqr7VAz9jZsQX9vp7EEP7K1iUtSmE1gm09Lnb4QXWR2sKK3
m6Hv1Gk/gMpf6NuIO0ZY57Fk3DB++1y9SOUep6tXT/iNtfEWcJFlVNJpvixmPn7j
/DTzQ8yibmPmyScnZ4OTAfmEgqON93wTB2ZgBJ/riK5ML4d/T8bxMj+BpAdzUFxA
ZVKvipgHLUBx6CnLGlEieRyMzNL7YNJfeigjKTSxs/u0AXqZ+W/EYXJuY0ojXf31
n3w6SHJPqwUjEi7MjqOILW06Ojthb8/LCYg+dOUkzfHOHG1Id+MOUwKkD5A4Ovq0
EQYDfh7ZGh3dqeeeN272s3utV/Ks2JPTkN0LBbQjcWCycxgfJaWquNyb14DFa1xC
4Dd+h97qkBj/U7TJs1WvB1Ieis0gnyKAykeEtWa5VsMUZ/ca8oltx3MkZhimSsrB
DppQZkkhVj/tr+kiwHKg6xqddewiYuuiud/Mn2VZzj6HdEvxnkMlF6DNLjOTcLyp
AxR74izf08YklIM7Xgy49FsmTCAqv7wJK0zpugdTbSIr+EebZ8jHSqCoEWWAM26L
ie/IdZ8mJteRcQnvjOsnyPDitoyviBFx6vKQJw3y7eyq6gBYRD7rnLnVy092dL8f
cIyZPK9OCC+rR4LBXq6/ZUyqHJWXQEjJsfelLBaXNKMxtmWD6+sdSZzN3gFvglDk
Lo+s8NWz2olgivIQDviQO8XHlHWUzBUtvrnouaeEUkGpIQ4+8R9AMPeK3jJXO5Cw
DwusmbTKO8+edIZkEdQ3HKUPcIJzsdidapjpgQuQbQeAjXr0g+LCahyNjFlCJrZS
GrPM86R9aMcYxvRRJwzzB6wcsszQqzDJByG2CyHSqyY4+ZMe7PHlTHT0l5opdPbh
dc1kWCU2X0vooKxe/JZ/fA3MYdiwO9zUkApb0gElWlWNXs2xKN9LKDVlu89y/9he
JuUp0t8lJLvS9RgkLO+2Jl5ucFtJbsdk+1zVCHAZbZMo0vRpIFz5w08uSZLqttIs
ua0GAUwiH4q0Vt58UKAiEBFF2IxvSwIHJaTbzQt3xiOaMP+QX3KIjG+65/Q7f6ZK
QQziHf4urRKevXZw/LPT0kcFL1By906F+MkLZt6rU6lo55Uas7oe6yK3CUkZHiPi
HDNjau91OJHbw/T5qlShKsfQkSUQU02I5Aey8iXtX4Dnp8JATsl2TAfruTvq1LXV
yRkRAab0vTuuvvI3BSG2gdNz5sZhnLpWRGWsAzKOwLzSL0mTs67+iDgNnTj5pw07
3wBW04pDSZlq17SQCjLSenfGq5uzkxK/laVxJLQZ8BQGWr8J0Eu8XZTLtZ47RCAK
6D5kghG79KaSz2wmwTJWZ+qDzDehVxcyUeYmAE7cvcwdt8B+TRTTtQbjOYzhLliI
nFb48mC8VSQpypw2XvMYytJ+catY8Xf0zdPQS3Fq/VFjYOvQFexuNEH4HlLJv0RW
dpaqzaYZxr0PLbWgJRDTjqorB3B9lvhoHWfyQIMOTO2Yt/dyaXqv0vGCqksp9vfC
67ec9gPdAqe3g0QOfxmJhBznedlIgdVl8FEVc8DYF1bqAaGQTYv8q8uHnoVz6e+T
Um1clCIoE8BWYzYvxW15qxp50dG8u/zyt6+52iIUaGlS1vfO+xR5zsMlYeG2A962
D1LrPpwxMn+2HTvxQx2WQoQxflzIO3ZCAROz8IZNKajM2sz31klIpDQn85odFv/4
P3488F1Y1gckEnjKBF6Ne5XqBl8sHSipTg7JwGT3FnwFPwZoKrTcMYYvXt9R48bF
YG8lHSDBtcF4ML93NF5Ne3wuiHIC9klWF4usc6gvF1LfZJYRyLPjPkNjrwLNQTih
7K77l+dZM5eJuE1hDDfnZJ8e+DJNaUOPRRDVecy2kajyl5J5Uorj0OQyHFH1XoUR
Uz0jJUCsRcv4xhOpiboIZGNuAss6Y6CMB57iG0HGdfb4aS6oZ9jYRUrRRW/YCQ37
IpdrhPFDHvQMO11rb5c9h4kZEnstembGKMWciLooCHNDlxAar2FN6tdhUj9UUywz
ELXaggWzRZJN+BAAbe4mxTxQ0FzvzuzUJfg26VMTHHbaUZ1E00i8VS8PBiedVskv
n5Q1j+ZLFwBCPlPj0iADc3bIPWCNmWA1RZc4Nz6cgXcraeZehCaD9zeK54rduQiH
VQRe/jZahbukIIFn97yzZe+nNOAdWb5u/OmM/juXR2E2aYRCETrTeZKKRHLouHpW
w6+ZBNAoHxANL8sPdvU5vFLcj5rK+8fK1ukuwx23UKz5vd3gz6zJXvRNHSPpmXiv
SWFvajCJpHcf/eVD2uMC2R0SJBTKFiZ1MBoPNRL+XIX4aMnWQR1o5wJtbcPgt/Z4
xnNd8asuAicCnyHwqXtq/GTygFm5HAW0CAGTOWtv3Np4SZ8Omil6pVV9KMd9KNE7
u6MAo2slXBuyESPOjlfpIWHmfQtC2akFVPEbfcrhZufax+oBUbA87ID4s3eczTIS
eSk2V/7hBkYWX1IWeFJjg6b4gKqoDRaMGe14HtMbFbJZfbOUL9dqaxLOvpJyak+C
LqMXzghukGMVhFt5wzmE7ZRRx5utuPO3WLJ+6FVZKy9bNxAAY6Uu7uyLhbsoPsQt
mBo7cvD8wEIDBPXDwKUK3ebn7BrkveyEeU1xOJWLsWSRJB92IsSeezbtORRgLZ9c
WE5vZ5IpsZPQrGmm/Mn79OBrzYoHDiOAtoBnlA5L8d/tsVYrdG5qkf7MY/+sYP0k
BP1VQ86Jem/QMPhSOyEME212+kTbmJ7in2OdcfRoNfs0pP63IGWrk+xRF4H2HnYR
gWhyQVNQqEclATAKTUq+YSkO8MndHY1dYzaIyGw1/+5X2pPpVpRqmWMGDhgVjJm0
8bXQKZbO2Yp5NEqgK4NV2Du3iAPER6qCkOWZyuvxLKr+Mf7CMIG/Cw8V69dFp7Ws
ePYMDTsduxh21H8bpbIH43JYVhFT23DL0GbWB2P5/7bGOBfLHtEIuY7mKiCGjhQJ
7x0V0O58SWBbl7RKtd+LId9BjPfhjFiTZ32TpsFNbdDDZ4Awrweq/771lHsSjvv9
B/HHyMZTAU++nW7dbanqSpBVhvlqAUOlCwT7FKyJqATANKki+WNNrPgNVERBsC3P
gVUFZEV4I/fvKENJkqZmu3Uny/ImpC0YDaJ41Y9NwQmO3Mb9Hhum9y5NDR8SPB2d
WQcJzNRlYeqgZwH7NB6vXkMwxM7OxKz9QH6QOU9CpPBUIRZGy5X/7vMVtNcI40O/
ejKUoffDYHCTsya0amVFwFgRz8lLFtg+LD9n5FjF27T7ZH/DxiAqDSV1hEqWn4Z2
aaCOxHj7MhZJkR/dx+9dC/ZXT2+thbF/U7qZ96ZGtc0fNQ8Vuy6P4Nrs4CnYZ66U
/8/BcyUfqLjIF++F34KoSuNWxj3QD6Q4rQpp48kXbM+nM5lUlGCmPxXs+OFTWGsC
ZhgzgK/+aJm9QRmTbOK8lAy4sYgp8PuSTSqgjWTnEGrsgqcLLQEi/9C6YDc4MPvJ
KGvI+MnD3RPe+bLK2RW2g8PTfyoWwQWCkYucor5tGxKr503oavlUff4nnKQX0hIJ
LT851jwO/EqBhc8BhoP30C5bvVvFzBbFTkvgyoawR+/cljNEIPYhJAKq1FlvUXct
jsEEuwHpyV2rdaVUfF4ZeTzI3U6Iwvbdjb6HaA5vG5AVwCuylpTqeuMugFpOU1sC
ZCn2kW2PtKsXWxiE9Ek77gkbwY/Y8fql+xEP/W53BaM5ZCRxEhlbpearUB90aqcx
4/gVHKfG1Tf2wXtLrckH+sxcyz2pcIxnMicj0unS/SCh6NU9Tk3jOl3NCpjlm7xU
WLEEKvU26NqrayFHI2rs+aSKVNzKGuCVlTccVMkKT+4Si0f2b7tY80ID1eq2fB+e
6v6ig+BKyPLtPW4LgiGhB4GFtMHPnNxsYGnCmgg4W4hzkbzFFyknQskq433nGhkR
qJTM/uEuA0zDxiUPrXDPTLKNBoO5r5og+A0Kg7zGkDfnZMfCTnW/pMl2LVSmYmwK
Hph0vow+k+UN9h/AiQaT+1JCmiaJbTAiTpKmQ4yYY1ZUGGtEpxSgmhCoEpZPlOAh
NFKrnRBBbeVZV2nJ/xKPH95ClqsEE2VJlm2GjaeqP5GFyI0FCsRDsvImvVUX9hoy
jBwlUo+vyrRPCpQyVGVMWzZaTYrcfiaKXumPLKtTOtp32HR9NM658XU80SMta0pk
R5chdABD5Nqid1yLLOcla84yTSpugy8WTkg2DwdzaFhpaSEigXGFtfGE/ViUrugt
RzAjIDeVIoKBhx5xO7/wG+iih1XmhjHSshy68z8lTTQseKkh9K4RnW1nPQZo2YXi
6ke2TeR1zsMkBLbi0QJoyZ02/cdqLxs/odLvGxOuKvz7HCr3fm65PojgBxDb+Q6b
eE1u99VCLB0Isrpmox+rJagU7fNWNNwNfcFp9sysQgpj00L9yVWfjfe9SIduZvCh
NXEemwCzf122HzRIBFmStEfxt2KTP1jU8E/XOV8jZ2nRoM81ObrcRrAszghSubg7
7lQBBPzpmEW7N2zy8iFv6i1eVwOYKrq7pQNG1yY6xlNYFm5Ntjs1Ge9GCFYRRK4z
E3pJ3wtTYmfMdelK0Bwm8JrImORODeak+AdohKs9proOupiyUMcUeyAB5dr9827V
xfA6SVjU/7ZObHrq5OSNQ1+jEup3suVDbyuZZL/GfU1Lb+LWehlux9VZelumDJR9
PGQIOeJdDpY8Tzf13DESo1zHLLnnxDbWbw7w95o4bLG25XmIdAGGgUbslu0TUh5g
TJFjKljFz+lJtocAWZgmIPNjgOZ1Y8K00m5SezpdZ+S7D06Rg8o8MprdZnK24rcF
YwCFMHU57fLODV+ct8SO3Gh3J6+Hof+jCzrr00UoCy03ZlmdSPs5WkdB466A2wLv
dDuHt7QxZd8aq+lU+sD8bUm+Om7WUwzXIl5gY2XIrwzaOq6RXa2cb96eCbzxfj+I
34Le8lqQl7ctdD51exEDsyQKGHJoXcVcgvvjlCPhX3BYO3zVWQpInjdQxtFNO1b4
XPMLuPHqajS0gonxKWRrVjxi/WbhKtQoor7ES/qhEn7PSNwyTTWZBIQW72GxdyLm
Zx59gd62TWJDteW085RpReT/9br+4XZHxJtKQyJhM4MSbAID7xGUP/DBt5Cu9xu4
HqNAPN/rpzWOukkIbEgABOBMTudE97gFiOsz2ePKAqq/P8p5JEvIpJP3oR5dmVmq
IulnqiKd8uSW1YAGMTOOOt5fb4fVyOhnMwwaFILeAC7KPFT9rT/jb2W0NY0m3mfC
YPmEAHB85gcI0RKJwNchiHVpZrxzy4panHgNtoytxzNyjVWTzqYATkC91QjCliGK
QIL8/BvZTK4Hz36o3EXVTdEE4R3Xc9F88gj981xNHvilouizseHNBy80cDy1xmv8
9fP4dYOf+KCviSBT3g4BRZfgaGlW4+yYj9AIE6Bu+CxPlS2Xd/CQP1IhmPd/7tr3
31apuV1n7G02bbbQTjLJWi2YbjFBOnUpX74A3NQqUUbBTp4Ze5ALAuQLYNO5dYAr
g2GGVecg7WB5CHtLInlwPaZFQ9Lf0NXaUXYIS5w2Eu8UdcssPvpJopmaf/Hk/BMq
wR95wTbsxC3wEXBKPGsikrPFDy03nWNI8R2JkhY9L1O7fAuar4VGCk7ZtujYssM4
K8dVpi91j09Gv6IitfZEtuDhwFj8Pw/9M8/r+tndar/+JQembQlWMxir59GrLbsU
CK8ApwD1avZB5MjCBjWrgQqLMDY343aq7O7S929llJy/Q073uKrP1i/a7+U10tFs
hqlALI+ubbdus62JU1bq7PT5cFvgszZLKJ8MsvA6FIj4Anx4SViHEBoApUdG6JgY
ZC2uZb3fHPhAnJTLOb4KOaccAXWsaMAUtL+6hu/c9cIQgDR2BLEtNrOrhmBj4l7v
PpOFhoLKrXJvzH07CDmat/Mj2bl5HfHG3GHgMnA4CSppvtAkwl8vQrCecDt85bGa
OgpgNwSg1yNHCam5uEoYn/45zB3c6uZneIxafZIG3FsKwgj6H4Qg7i3NatQe1CEm
SSNJ8QrLqOxJvm3CFZU5dGlQxJHVSEsNJ7IVedIDhDIWWsMzzKwoxDfDWkk6jWUR
1Hxes8v2tIN3bd8PnQJta+sUXw0hlJ2cxwWd7hh0bflQMF0mNZSbqJewmilAa9mi
sDUVj3Gq9gOqiOTl1WHVpD645zzZCeIjGHQbnCiEkmWhvs/Ao9Lpaz0toVu8PUIc
M3UxHC8IQdtggwcYVo4SrgTkDOF4tbn4gqNObF2f5GW/F4mM2clYuBJ4ax7qpbdt
QbCwHvF8pMbhLJX3ttjDKjnkTXc4Lv1OcbjyyyE/cZ84yAwKzEwB9yd8MRCfJ1wn
8y9xVcf3XqsrR4T2aDx2fr6g6QWAAab0H+BLEMtkA2+dOz+vVtg2UT6cxu4452ea
rHVmjzIZXAVnXXtYK6W89GcsoVwAlepsHWINvSIYv5EHAZTD9eq0HWbky+fn3Pcd
NHIhTSKPsKvqYD9LSLrtYuOBJVZI5TP7sa8YrS6SSkAsDSLsU/ME+MWh3Wvx6fWW
C5f/oixIToFWwvctGt8xH1N9LXpld2+q+5T5Xn8uho9kSB/0cHynfeIsuiM36J9J
JIz1FNMWO+dspj1ijE4Iwx8TUaVxusIeVXgUG0hHyWV/pOBFmElfAlJdNngjW+Ro
L5R+aq3ETCKYB5zpuWWvD2yYdQjJBvogfQCgQpQQ62WrH5aIa2Ao7RSCyfJ09oaH
w5meTg3AUe5pUhQh8v6aPU/lTgyV2Gj7ueUXPLovvSWU26n2re/sk99onOjacaz3
hIpCWZdu2kc6Us2jc0JYcaUZFZX4s5vlL7TiWlekKBfb4HZevwykEoTQnZWjlZ5L
6fgGn8Sf4cLhK54c8hgbKNgdLLNcsiQ/mJ2L24ckluSrEC0mO5CnrJYAlcyFGhhz
b+GHBvyNFAR2wQrvWLruDhy/n29x54xPF7XP3FTGQjupRtvBH34KFyM3aMRqpDZz
Tj5JWmlUdEeD1DEAWj4dasb+AqoMq1nyROd7Y+96v/3vgLBD0EichfGepGNn2G3q
XXxvKZnxL+kURJO7QqpbDwYOBrZqNqxHSHpBVlBqtA6rcFFMa3QFG33/z/4YX/F2
QzcKj47d4Z0sIfhTgjNeYMGstVaGUrN/LsLERwNmx1UbWXxe/HGlZOzNEwwwT1uM
BY7k7KitEn+HEDcvWHDSMWYtUqXujg7WxLtqz7rLDO3LHn4wTeL4EuBJRt4ApwM4
BBfapmdEwg/a6Kr7rH/UAaQV2IhRF6pKB1SahkGFYi4oRgXcwCwMR8QzKVvPQR7R
/Fe7FR9ie2MinJUOAnUvnfapycFdM1lskE28i/cXv3FWltySKNw8JBkKwv8AYU86
Xfig5YGDMSYwC1XZ4/OFKNKiGgRFsMQpMv8vkG/lIU6a+zztho85qOQ7YhY1I6UC
NK4rMG/qnnWLuSYPwGpr/qnDR7aGoqWH+eGm7zLcRIZQjsu3fbrLnfCb+/AP80gg
i7DyrR6/PU4Hs/mFOgVCOtohoqL8VEQev3sfroI182sMokRK0OfqwA0t9JDixfwV
ZhI97lphDcv5LdVynbYA1/AwGGeaasGCUndUOy3ZE/vcX0FOYbZm4QLNcNBGysti
4TkSSCXO61u2tHGuTsidUY6GY6dNtHxZ3uYdZgnmt7cEACqEbDVZ25aKBOy5Gk0p
S21wUi9wqTnvsp8gROFUWL7m7Vnjfrlq+Zatg68T3HL+Dfa0AwbTSZ1KfWO5hzuF
f3rsJvWkUKTxj/Nj4I8oTLdeiLreysBEZgw/v+aWCcfjMKIBU7jiefbzB/5L9aN3
nNqaXAtlG5qyCKLgzaZJrWPTAY1j2XB3YDSryknePUXWxqDYnDvPE2f+Vb/uHI2x
pAyZJ2dYkjVtWv/+Y+p6FFN2rTzlKx02Oi01pgUWQwqJbNuFVUFoiO5wLD9kjbk/
2veKfKRlXUdJZpftTYvS07KVZQjVB9agGLtT+YyCMu7sWZbAR7pEVTzhZNXPF3Sm
90rpa2BqKwEv6ekQuBknd/Tmv8T3UdlYYx7u9HYFdfcbWQ7Iasj7qTgI5mUSfPM+
+PlaBHB5NzNOADMY7spqPvAK2ypHH9bM0bqbzAk+aMM1OlhXulqlOaejzd/ab9dw
IaDilIde+iFbYLtbvhbcV5ODFD/wFV6WOEjsoCM2yl+XZqx9Kef2QuAZ/vo0CoMt
HuKZ1+TrPmlFXCiYGfClq72v4K5gBS6dwbtayg0KEm6Ijz0jTrWlz33cBNqzXo+e
kfT/F4XLJ5Ym8hlXDZSq3VPVAGo8tJaw7OS16LPkIOevgIkGrOiWmc3aZhF7YEZp
J7XeWG3mlxynZ+uSZnlO95jKZjwOxMRCNVQ2T2LnvCrA41R26T04zNK0I/nbj/id
5XywOK47P4Hnx3xaFtI22tqZe3JpGrkKiw1MMXpZPpS4eHWBzFBl+cCZwOosyG34
ZTgVK/bwCf86b3WVmvOOgWBz1Bev8yaeCHvAk+PMhEQruJQ5/Gfm80On93egIDHw
BhDbMNtaO8czGZrzpb1WbzUtNArElxfTQk6hMgx80lNXnXstetRK+dOmI2ccK0to
D7VwdMOSUAFo6Fp6ptlGXHtJygNoPI3Jml4kGh78DxNEkB91HnmF3WzzW0GO0drD
4a+tz0lBVUZHBtzhckH9Qzukoi6wwI83zTXFVrzKyzb/uw1ECs/+at439kX9uwwx
h+oEb32KRDOdtJDLZeB6HeJFZXnL88QcstZ80pZhrBxSOkh+q6PcBYGIxBrtH9Pn
FgN0Qxxje8K9gyZdMDIrBOl2bd4L8uxNYV7BUWtaAFWdR20ERcT9KhtLGr5NJelb
KqUZQ5AN9m0LK4LzUNlmmLEm8vpcgza2zCcoQXd3WdBTyhwAgWdqbBbbK5wt1lon
1FcUvyVW90PEs2UMEnLa55H1wUcLLGQzmtdOco5iX4aBfy0z4YvKYScSg/CHsHZT
C3rknlFkauPPasHus/X7PQWAAiaN491NeiPdHKvDQCPSiKsLzzC2VutCf6bz/Hcb
3w7JNwAEdUuaXRgQqPmD4//O62V62S5krkdYXj6tXOlQdMp83mJf8OF6/AlFJ0Tl
rUKflT4/3CvShArCRt26T+pbxq8IVOOekaPoIkNCGXWTcSkk65X5dK/8tDHCUYHJ
TBe8qpRmGBBurV+kccsgEwDr2otSyY/ujsyPuFfgcD4+n4Xa6rOfWPz8t4fmIUHP
v1ynKUL/knNl2Gwh3vNJk4xtJphpkkZbpr+7DLIqOZDo15oNeA4Ol0b/7ppe+SR2
tMR1wQAHcvAjb9ExKSS/ybvm4Nf9zYgAzXv60pojAIUPo/Nyl0srJSGmI5f//GrH
tfu9xdiOyoORBijNxHB2cVI3lIhAffFmjIrbPTmQXegUTU8fC1LRx1yBo/Bvnrac
9QnLjbSRibKsZPOa29gYcPsKH5F2ywt7vRlF1ldCDKD9S9OBBBw0Su3KUndXWA+q
dwOo+QexJjZkT006bsDN1ctQPHHSbgcbpvdJ9kj/st2N7gr66ziao4BpNygT01hA
Wz4tX1JhU8V0LidWHSo74gT3b38Z4Oqsctatf8V8orh06CYSoXCoQDLVIgqWS2NA
2E3Pd+2DjFRShTgAZUJINUQOd14saA+UYjRP31MONpId/WJN3Re26bpwUv5qx8Si
LtXnBkEreDfl8PzUVCR/fDWXRR0ZVYsVMU4CMF+zZFNlJIXIC26ETAiY7uyGDwgJ
14YQcLDJ/ol1zy9YOI6bLvLrcFg9rH65uGD+ac7alAqIRV3xkbxMxCFAK5peNFpN
AtsfGuN+IQmPvfF3tJRqaZh5CdZ2Lqx1HYt2sB8UnoQ6N6X4lcOxN91+KNyo6ge/
3/N9lfPYbUPZvnFxaSih0bem65Shlv2n4gQA74ur7WYkUCRl/7zGfZX7N3wdebSG
4s8b6rvHdDQHH0K42+GxEJx4nqAoW/v/CCBQGtaMtxeSSrVcYI0IcPWbRep7tUtN
n2xKhpNO4Xodr9c/JPmavDuj3N6hefBbQfeEax9H4xDA9HJAPSFqyNi1e9YgN5Zx
9sj6uFaBeAwbdxY0oY0DKzYz81HWCVzlzUd2733aIzItNLjHwricpsgIbLaruXoH
zJarOu6y1Qf8kzRKB4TgahSdhyACxt6j28HXrgXHOWR43IGE7BfpjNLHYXLS4sLG
NbNHINMRB2cFH8A7XMeuyDMZPc8pEKKVj6UABEMWIRvpizzEk1dxBrM5p2IQBtrW
9ZGkNu6xISIPdGChji0uEaht7xcC6GpIrw4xld2WEdscVOiMZ10wOOJrc+7iaHhC
sVorHG4bbP1wtbDPJXKefgh5XEvXjb87reTPOULH6/u4h1Rn3ysvJUEsZ7J+A2pj
B127FfkKmgsAasgmHjP4kRsWwH9MYbxPHLz+8fjmRLs5iXzu8ZqD5ntHDY2SSzC9
iZz+Soatv2ZFo+nFs/L/zPLUlg4bGoLg/pHktG9qbuSu52uNkeNa5DPP9QClbJLe
jnThS4QRt64iHMijM4v7htA9QWf5GVMmbkkBnkGSwFzKbkHkYhMMXA8uRiPn/21K
QayICRT45b62aUMFx+O1G4DkGdyZHTjJ1u1pHNGF93pNE+jVrGrNXPWs6BlCTv0P
ujwDsdryDW7cCppRwORPfjhLrpz66XQKxrOKTQ+7WsaqE7IL7BvyK1/v9Xisz3kr
NIUmYhW+ebQcQHiY1QDadltrqI4QRqX1YL4Cllg3qg4OMnkhKJ16xhiWChPgTQc/
10IfdRfeet/rAJlQJDlYo4mnfMnt48UfyjM4eu0pZ0qb9pRyfIjQPgawOpnwuob9
Uk2qcN7lsNSUgO2jCZQwZ4S5jaFVeObpYGjftiJ4qb9W8INrJezOFsGuxHVnCklz
X0UcrtYzQd5cQm8NmrKE6OPSFWTRBmNYjDTYMpZLPQXu0fzbGdLtvOcC9HRlvmXS
QYfzNeuf7+vc2sPka8NdrouN+t5pLKuSV2mvf/URv1mbgKgIR9w28jr/rUx2wITS
40pAHVBcVLk7mVBp/I3PAA0o6h7UBgUkhYWOsdx77/VsQeVVDPkTI7iqjrxUk1xP
YIkEDy1k9I/RiGoflL/vd0wNUCnouuYiZ0h+gYr+1OxwME9m2PGQKMp8htPqHya5
c1ayo3Mam5Hk/mXali5u5obf8ShEBQ2e3gd18r2dipo4HNHIIkSfYNcI6i4k2C1G
Ie3ZdbibUjR6bdoWn+K79MHbF6NLy+4hjjXMbPUliAgj2g6NhrcCM0ZB9fvxczh4
N9qSB6mlEmWgIUNBBMCii8Cp+LRPtu88uk3HUSaieJ7ORMxmbIMh3Tz8jHIKr5LG
FB5EUyLGUoulcGlXA8lowF236iDqUpb1VssDYG4aIpuXFRAGMJ90sFrLJ0GyH4gB
GnOO6/qMaRGKR/mhl0maHhLbQTP+0Y2udKlBs60XAt6jBO0A+f9ZXEYIO8lOSGwY
ruSCT4SZvpTN7l/bXi3/I71Bw0p615tADNlq194RQ6WWEuQkNnDhSJA9Hs4/eUSp
4ll5brAuGJGjMSDHhYYBx1Kl3qhjMFnMbPi6ZVZKxPgS/75P9DpmWHK5VBnC2IGd
jgwzDKoI68PHP8UiLW0pIqjpOPp8NL++7NHibJTSN/Rxgv8tztvdK71+usC9MoVu
UTYzyL8UvQAnbbmjRCF42Ux7PEyqAiGYtD27/iI3yJwkZI5ZeUVcltGj12Wyy7vQ
sBcj1TS1D9e27hXCx4KcP2i8AYFj5S3aRkTRIOrvmodio/tqWnSFAvOuyNS7KOls
PdXpPdlZtIK2m0n6t+PJehJs52QD9lIKy1HgcXE7HIMAjGOFa0R6jznoK7cnv4ub
IpGLsOV6Kup1ochmApZgwCgKt89oxAQwUo5TGwJNx4J3OJ/oGmxz+xxCITiQBxSC
CApSnggbISDpKLCFTZO+xHEMWZ5kfLsyRFpWBLxbBsQROcdO0bS03btRpsz6/R2j
FCEN+cbSKWwh9ULXfhRplu5mGCknad8ZNviuuPPjoyCg3UzRTAF5xtrdhpB8C4td
gDjaL6CIi9iEufh1KCiWwIV0Po7hFec41JFog4BZh6M96f9NZX3E5+soaVMYDjqC
FZRI5TdVGKnKffw0852QdR3xfK/LxoRfBAIBT+9c4HX2g/UxePQIUPXpBO4/Ieoo
/jvSHCNE8R7/1HFAxGaMqQH7iu3b0BsJsOVFLzIgl01uXqJJcVI7x4MNP6Xt5KRb
IDwd8hR0zwx4TpYIkk6bJQFjiMzfIM2mq0Y2pOL4f57dYPg48IKnF/on9LqrA7e4
yFRLMVL/4xOQGAaBj+Mxuo0wHrbYjaJkxPdvxO906T2WkuThrZXCMurkeyitz3sT
dRf0/nE1ben5z62PYW6/VL9i4jcGW3yJkPsrkwWCD8+dAtGQ/P4vFZfVakmktgma
JR/Z0VrzBWowyAL1cKAvvlm1cUudKmkW30uv0V9MEI8tIYfT8LiXmJIdLzAT85j6
WJ0icxXJAXczpWqXR3fSALVomjud49DrA2omOv8j2I2+X5rj/n8yhwXruKPoam4Z
O1oojHVSd8UMQyrtRlz4RbtU0QcofFelpa9VZG5HjK44ic39VzR/jg0TzFyN/9md
yzzfa4Kn94Rx2wsHAbAHB7Ft5hLlCeWBGs+AIkshdr774kBe0aD7ddRtvUjbZ6xp
DYCs66DhM9i5Mue+aahLwpcSXatFr8gVWmDQJwJnO2Gv0ztr1+kqW0La9cvWsn+M
bqcABvtBzONO0RVUR4hhm3br7/jhdse8eLzp1ifiDX6kqf2gh4mEGlspl5bvgFoR
QeNpELLbz6crIY3rSZ4RsxbUI3JFWRUdgGqGL9L39R2+yqRhht4f6H6Vyxirelxl
U4SHNJgmoNg1XQYgAX3ymsEQ4I4ogBGZzwbGxGwC7Sq+ucaIWkxs98lucF1ewqm6
kpyvPpDAEaV4rqGe27kPw6W9KcziXUrzEkfNXYiKy5utE0+I+RyJOjCiNRtuZ3XV
6zXpRSNmeHA3f0bWDkTWEerwjJ1Wc8gfkwSnAFLUjIqTUDkgOU2QRPPirx/g9y4S
MayX5JKu3Bhbn5yj7Px0Zlb9GaWnEzHTM051Zv6OJBHywH2jbcxjfE72qGFQT4FS
tgtUN4YzeqB0fS9XBulEYp/A/j59hDCeBkAWdHvyJNHoNydnYudsR0ovrB+fUqwc
ctkfvqd0g6uG/1InPaeSz3wrPNkhdAdObQeIGWSsfdhVJt6yAGjD1XCEHFKgkYGJ
Y/Qt5GEwDbgWQLu6awhKVD/PcdotZjB+goOw0xL8wfq/F8BGMq+eEKxaAyLOEb0k
Jg5SQDqb46u9TGoHviSTESpDxOsBL7Vuj4MhEI8rG31/DcG0E0vOIBWaM5wzxZ1G
OvkbRDVeSy3KMs5o+HKvhTiVaxNsvLP+7yFD8HVtJIc3w3c1E/+8OKublnW5iFPy
Dt2J4HH5mrddHJP3ijYq2xRH9H6J+i+wbPDz9Bj74TaMk1YLQSBy/shkr/nUJXn3
I4/HarZHtBjBgvh0/+JBXBSyg4C+BUafkUzV2QRabNAq7ziTAK+Y3P5t6QIK5lYG
IKyWFdmXxgd5EimnqVGAhOy249SnJkG21mkiNHs0rBjPn0/45515gUlNE5FILlhm
ASCWP/I1obezqhaJsUIziOEsK14pPYt+s2i6XyhuIfM1C00PsvSlm6Y0+Be47o5k
WbIlTmSqHWI+trmT8w1ybhtL6FDdsNm8srGfqCrbpB4Rlxu4+HMvdoCMam1UGOHJ
F9+J/M5gFV21Nv4M8PgjHfgvAi2MStnvKvXfb4Tl0rbXf/WIEG36cHucMmzRJkv/
rQf259+9Z5e9pSvXVyAfparn9NTlqAYbzRRg4Fsq0q/guqkbgHOkCKlvNwwg3esp
F72OH67GgNBlLIerJ33OsBwnkyHDklqJE5iYJvZgYsKDmvYaz4/eDT5gSQPuwIrv
QrYWsSYpNLqB1us9Mmwhz8K/d0PI0E/R70EaVMt0C4W8WQDJklDfFmoGWssET122
evr/bHuCDYm5xu3M3w3k8h7J2oK0RiwVbd7xtTGT4Tnz+LFHtOKPmRDz27YoQFVi
v8BhDthBF3ZFSxzrJDIHuSiYv6rFeGMCEnMqJIvRZg3AkQYo62dExDo0G6OFz/9I
kOcY3HuYqyDrtXrYESS2rl4Kb5sJ7GKSJwFNgetNpPHddlR1lSSKmiuORh6Maj8e
nCQsjl2d7FpQEqWUbQLRp6M0+efss9UB1adxY5QpEJQSA2jB1hgTXlknh42G+kaK
jsp924muhjKbM+r5n1Dqq+dsfT7qi++AH/QLfck0Zp/+fGfU7Tq0AAp+NGeBIeG/
YbHjV9L7rY7aE4zMcBO3QfiWpuz9ns1XqUI60FJYYw0wxWfTF1SaZSh457ganHQn
ODT2HOCcbIrOQB0DfFyMsaQ0FJf0l0hq73BR1DKSqP1XbHeQjHkGW6HUCadmcGpP
TdrmECJVsdz9z97xyv+86cxWu8WXZafAw0mpYU7RBdBdeihkgYsMXd3F4Tbo2Tf2
EuO1XPvbKF4xq+fNg2lNgXoihLE8GpdLi8voD+tTggFK0gEdt83trOO9xVDKVvLl
94/BFKvFMd++aMoHIsmr4zPRqbHOghcA1+EPVZyZP4F6Tfq8n/PYKbQqAWNJ8SVi
li7gXynayvbkfp+cViOldXj4BcbL6rxm7C444Y8RMfZS1A4j7haN2gZO4Yuk8rqQ
HPLv1L9b0tzf4zfuuKI506GfB/1VHDWpwtDkGx8mQi3VTnODyJGC741ye5YdLeNn
QZ1copvYjifoWYmmCIwpGbK89ArVhneWb3Lvq+etc0hwKgOO/qsloKJmVYPQmuko
ePVVC76W1XLQLmRqCb7RZtN+twdts5PGCEH+/0KHJThwSI1qCoMZIcnq3ga9QlWu
PheqT7pNEbMainl5heS4kD6dXmZ4LHN+2gMQGBpeLn//8zcuJBqohQjIcm6utczX
4z8p22tnyEC6bfFBeOXu3r1aSeFM/So+QbAtgrgmd0klaHI/RE7gP5wSFi9VqyH/
fDHQIVPfbQoijtAtwjvZwm51gXY9coVIDpOVRAfLQMxcM3Ld6lBNWb20XqzquCyP
2xVTwNbk5QA54bOWTiQaWEHVgcHHnVPCQ+1KQspvMIRifPd+dpN9rSSIn1lmy8Eg
eEdZNlXAeBJgPeLQ/N6RFbeyvDyAXmOnaGx1G17p/uDAHsMUGCER5HFfrLN7bfrT
ERsAnn4yum8L3hMyUQ42OArkGkOiCR/CKIE7ebtyudbk/17BDTw+qYvmauJNbWX1
8KpOBR4JeUscnPr6Y33Tz4FKPL5cNiSwoAAxa/fYgTzaEIS6CPWcFvJANEMcXPUw
jNthBcsSFKsqXp9XT/MgwEp8n4SfEnb37KPNfdt1y41gyfLb6f7mb/cCepWQ8DUw
/Qsy78vpK83v7tZBkSBwdc8DLeby3CPqMQHrLdGMJgMqwE26QSgEuVNhbbDHTsku
+A7WNeVrqXJRIkY8k9j6/Rhi+Q1iASpQpdnDJwIs/PSzHIBiPzWLbbUVdFatY9gZ
Kemu4v2NSNEC4atbJmQ8zilWPo69RTSky5Rzg8xcHk1J09u7CynAS0TqiTmM9MsI
OoP0/W2qsbUifgGgTB4CDFbGTBAvyk3cTVJntLO2BCv/UKxAclhHlBV8cf7FqxTc
Oo2NLZVWuSYRrdKrqInenjW5KaNBkcMkKizvW4r3PyMrNjuo5g1+/lKw3uAO74zV
UusPwC8h5dqQBralvwOGyM3Nj9HRGN7fh4dTc362dIWieUtFM3UcvXnIca71L0HI
wXycrgt/5foBVLw+l1k73CAhua/mcTh2gVWrndAoi1hPMXii3c3BQmowif4+16hV
UiIa8mNBgppEEPnrsADuvWNrPfkXAxkG+zosgNpGZXBvR0F334wuXvRaFQnZ1xue
rCMGFYSpsKm1Adk4y8itMlWZs1fA4PdNDSxBPH3HxKWBlePfzC2nU+mt/qQxqnIP
P20vKyuWr8VrdvzR/NB10lTgdX+j1wEty0IcGyD9g8YSAMnynvZc+WRGy6AdgAhS
mBP4L+5SkCbyJ3hc/zeiNXNtiyLWXKORHAJO9HxqxGXlzOd8dbj8/0Csmc3ZF6BQ
d+ueCQvkemgJ4gNHxBn3jZBkgguvClzKeLebzzH85IGn00RNNI1TL/Hhj6MUwA3Q
IXtpOtRagP5Jrg6g0PYxEmnPqcbRCqzjmAlF/JWkNKyRgkixBK3nIFT0mkLueF31
qx9Avo8p02TP9ydLeGNGU9qyDEfDkTtpYuVTT7PZk8PnzWtLtiXn8IBpbmzg+Fio
7TJBrqz1apgmQiDp2k4oVd1AWTe268X7Z8PZq8nAE9FTHSApdHrysR2sk+oVBGWd
PZo7N/L6eFz74Iwz6h1Vrfqo8m35GseTH9wwdP0g3Yg6rzLsLLyHYol5XcUyJkfF
hT/kxB8A+Tpl9Xpl2KHD79zRkpWsrz8IXyAke0b7LM+G6SvboqgzkZXlex8bvpR3
7ZBupvpH/UEAg2QFJ2df72Z2ToxcdzxMbRmmlGoSk83Z6s6sPDJFCX0G4UNsWTZB
AG0J7amSab2SmMe67lbSqWkPq7hN+uyIc6RObb35pEIEMUI0pENIGtXYDzcocEhE
tF0T/VXYdwIkLf0kAQxU85DjhCahxhQc0V0ifZpCdxUVr0JJiQZ0NuLGM69iJZRD
ta5xd8L2hzxdBV82EjK6Z212cisJbfEe2GowDwylvkT0hJ2PXOGrOxIL1bsi5VU2
bvic0vSi3ETYJ+XtZTS0uD1X6qWGCws37el1yF3lRJxdRBfqnZMDxPpxAdGTZ/Zj
VXeS1F7KA/A3wrNrf+UtiHWhWDMzF8x8x+RUZdbLOcmwLKavuwc7aaLbL/y4EDB/
+ZfVMX5hm/w/RoB3tErFTnnBEgYweN0HFeBxPR7Wvio92fk8zTI8BGVLku8WIfwX
EWnhksh1zmB7B67bx3490F9oLA9/dHOYeFwA3sefUyjHLCjRgTZDTIIbSpC8M36n
RhPa9JZn1Dz45h7jmGRNcpzCBl+RhUJpfogwlrlG098k9niUiGBTtdyv+rNHoHZj
0TssefxbQcCB9UYcVxw1fwOegUA+XuHTRGqLQECwSiAODpC9HS0vKh3X5XGMiM8g
yblcvKAtHRVEZQNt+pSFttt7OFdPkHVXwmu598ZSK3g6AkU6zPOC5IoYRqec7jof
U8UQkm+mXUom3u5TVECO4uRyRxvgv05wGO8vz6z1FSo7geYlaNNKJqu08I/d9NNA
T2cLZZcKGHzWKBCdbzUg64b7aCXyROefGoPt1NYusfIZuk38GrraPqtJu9sF3LaD
LOAfF8SDqPlkluhT8w9ugvrzDDN3U+ExcmVIEztq2E9OGIcdaQaB4h4HU7KKXhhB
/RsaQLupW8VIKDQpdyEiv2Yjg9Z3aRZHcO9dIcKg4R0uq9DYIiWk4/uAu+QgT+k/
oqh5HZtst295lMv6b38/Kw7AeifmZ1bIcBdVxQYyvQv1V/Y0cSLJre7WMnJvdc4H
db8wmDalNRsLvTnQll6nFUBjSdXpgY3DtuzrKzRs1DUvV/eCzCLCscOEtkoNagqa
5pPtm3dG/0UeZZseho2TaOEtDAFi6aWiRwueJNoHsmfM+djoapkvhas+rKnP+h1y
jlKvA2Iep91f458L0sN3ddEgUDyDHy0+uVj82tHzoRrD78/sevTxnszfg4NJmM3X
/JcIJoTP/cJHcHCbyOhjx6heQHU8yc56GKLaWuOSQ1AZVtLSAjUVmwXI0PsrgPrS
xZxkCzkdlnCufiQ6UpecxGuErAYYbvKCtFIAiGXDsLt2RLk06pPgH4Jylm43b/fL
5EntLPxEsZbZ59kQwJ/y6oyQN88+7q5t1QNTxI5Q5KZQMw1l9fzXBHSz4zPCDfFB
Mb5o2VcLe5X5EZGao3N66FN7Dh6zlNGl3tUJZ1iMRom9At/hu7w0jPzhsFW5DDC4
p7jtuY0OMUUtF6U3+ReQ6as2w583sgDgXzDpoNm69BtMK/CkOVE3QAUeVfjHt6mV
lLJSFaFfR47H2lZ/yfGw0Bx/mZd2IKVx3otEnA1yFiUZopJmX1zqDtWuTmsmkWdk
D58zka7DCQ5NGiRoQyP4U90v8GOfDzo6xxA/8YTSi8j6OSAMeJbAXktwyknadveb
m1VMTDt6bZQxVRrHiTi3vbLbaVycsbhGJv3ieQvEYp9u77rp4wVxb3w8b8gqKOpB
OyJ5tXZ7I7eEXq6myO9Rnv+e80ipTAq0SVriGk3KpRtb+qdFjReMU6Y9oTejQYqQ
ydO7oPvvFf2u0nGPBWNNJziUMavqglxU827ebHTXPV8YHwftRYkYkzTD/eCF04k0
HQir/cPOLbkT9Bphl5DKJIhQBPuUmjo1G4M1rqIMN2e+Ein5pSBhpi2bc87/vPPs
C86xnUTOyMo8wXJmLI4RCU+qvF0td6tM97c7yS4z3/P5eouEsFjrXJEMM2qnQ9jw
F9Sh3l+brTazLB1bYN2aNn2JtLsUrq0j5eK05mpIvZZEKlpfftamHqyX+FuhpAKM
xozEJckt9eluKgukicS24ymOYkVyBrVmGQWbRNQWrHyhJmDAqB3+tyRVll5S/z6Y
Eyz+bGN8sVNN9FprFl2qQgudo7Se+/bX80PnulReX3VytFM7oIrsjK5L/DSLoTrD
1qLjMj/ngxBA4vNmeIhmQeVzKF4AOqnAqYPo04TFFKIxVCsGUYt19os+4P6yq7/v
/bm/89HYUnfuKqP97fCU7RCoT3/J3bsmbo1oI5hC26dggV1ksqgOzmzipq3iy3zy
OSpT3lOKFSPjskeyujXihu/5jwgpx84HoLxD2cMpHVP1zodmJSnyug+FVgEl6HOU
xr37QufJWkmqUBzxWPJjkS2OVTO/bNr6JjmoJ3tp0BS+emYxzCkhaNFfxsgHXToY
1dlFKW8fS+g5JAHxfdt1UDH7oBjyGBKVrvuAbTMwvzjgYW7AP9+2h1PoAeOw/Eyd
UEZqaDuzhQTEL9WZXQ8acrLYcFxTpQgnsOzabi9yEgzdI1f1nEOPLtRgLiY9/ZPw
HvpcXUbAUfHTY5uZucfdeFcd1alEa5U5fP80nflAPgfUc18k7DMKdQGebTmgx0Qx
E1EDqbPYUHf4NQHCi//o9l3FnlNO92oHOPpWIbzYAD3hryq4S92lboeChjsVYU4H
6wWLgxnGKFucAUAUx9CsYZQmI1qwKcRNoL2Hd0qZDnjrS76140Zgj1bLrYRABuwR
1jP7dgbRXGE2f3s7kOa+DOSEJq5GCW5y2waDacCE5h7MWTukGO0aA4zlsVKe5xgm
ej+xbJT8I8FsDzqaol+6oSVfE8JoPy53pTDvSvIpG8XdgyHAoUHDM5TmOtz8vv3G
L98QSnhBxVM8ueVhG9i49QgA9ffvUcx9L9cfjr/gJcelTtqMu0MsoYPkULJWVNzG
OHjNsufSkdvIJwR6/YPPPv6wnj8ocquIG3SVTc2KLmVhgih745wgmvlvE6sytwjV
xAhGt77EOmQPosWL2Z0mcFnooefjKIsBzI0khaAQbYtDJCIB0w9haI2x/EWBqOPV
HN862T77v0aXP3DFWpDSIaz0eRwr+c/q1exTMipDrbX5o7ejc5N6GPfbZmYnfluo
WIxWiFFHURvcjLXzScsF8fWdlqhPr6Bl48K/2v9mSK7t7Zl2ZDM4uo7piI3NSnND
1B3kUmY10Q6d6+952MbDzT0pY6ItWYtYWXuyrxp53faxJ+61aRuWsn+Oxlmo1u6s
iIPJ7ktSxbGK7wF5lh6v2NzBh6AKxTHhD70OgMtG99uCvrszKP09xu4BQTcjLS2I
ptxam0Z9/xABfbSeV9nUTn4FvaMAK9cpxh5kZJnNF5N7yt4WbhiQe32H0mxkJv9H
rzAkrMD6S//ksobPe962VwNiETsbpS5f7ruHJMg1yZtBvI1JveiAjqXXAqyE0ULD
IiefweY+iqequUjv2g0aUAjzeVfCAjJyaNhGxAxSoSPgicu+Oe3uxGufRNZFt+HV
qMibDUTQ4p7VUl5kI2u/Bmk1cXWA7VqWoXmYtUdK+iOpdu6gvCRmZWmKrsw8Hlyt
rCC96I8574exCr8BY111b5H1y4ZlTZ9oAAdoRCTX7I72KS16RmUTuPjoJQ++Jxs+
zxpr3kyJ2BQBXfhAzaYg5SAS5/dji4DCU2uzmodgDf1mhusXdHaF6yCTSceZLlDj
WAh7N1C50W3lzgIpA2nD17M2XNhIN1TINXFVsRni+l3ksRmub1LDCA57fM2Gn/vs
MzDAgAh6Hxd4fvsTOT64YNiWEakCH0ZSugmmt6PfBI++64EfDBL18jZvWRl9Yud4
MNyqEHnDMsItAuqLPtJTTQiRFChrCvnHDDJ9q3d7g7DZCtLvhoexIYPFSYwFRf8Y
EareFHRY0VSEvorgHahfZZrlE7ex2SBXFMQLxpD6mp6YJUDs3NdXoWjgK223DTp7
Czy8Z7kaK6QKJUoAxYdvtyy5B9lWMLUa9SNWYO6FnJII8dIJmCGfyYMgZGaWb+3g
cP4ZGa02HFCpx8H9buLOItfPwD1TBmlQLlOqriT+01+JCn7lGL81GKV7O0mB2jht
O/DWQVQ5DXD/st1V+K7m60X18lqAHZvpwE0Z27GCvHMTxeUO7fXaOpS31Yi0IPzI
Vh5LWYtLVSdHvolGRO2aIFkCFbTuFT7JZjn52jiIY/AlEdY8wwzzRf0JgHnc13nM
dCoSFANxPyBSV3vHFmar/GDYG93idvaZ/gSSDfnNlahMyl/DJaumUfHmWfS973c4
JmtNOJqDE5mDEnquZBOhZ/K+IWUwRbhVUnul3YssDXYbpj3RyalJdTGI+l9nfJlS
/671e8e2jFOE+/a6cGut8PDfM7zlqhXG7DHlghXbH3WP8JL4HrJNwU3zztC4bP9K
2tO53umxVH5h5g8LBwPl3yaZbPI9H931lJXLUmuhrrVG8hN7MMjsl6ZsnfzZIrcD
1wS6AqACkdQg07Vc2DkJpx4tuD71yJJLVIfBrumtRzMHPD0u1vnNKWSkq7ilSS6X
evAPgBknC4W4TUaQM3mFPjHF0PTPZcm9A7eDhakxLQ2z3dU2tITwhXcpSrXk5IJE
1NNEd3+9xkls3yAzzLsLB0jDQf9jJvQHOtgN7HTd+lp8AMzBuXDlr5YC30OAxr3p
h7zokBkIkeqRclIHjRwT2tVL+2zHgxdJaL77I0DvxMCeTb4hT5Y5IdD/XJlFTsmu
o0EfRZVW9JSpxzvrQZusxQsTBZOo9XhjYtiAOqETHYWVPw9qTGEHtU+c2foaAE4h
mkcyJMS78wuyvwfPMbLuDsSs0c7QpOnM8bJ7C0pSCFRO9+LQ/gwscJs5tHASxyoi
lPiEY+DwhrFc37w9Z6Y8zbjomP4T2/GXaRZDQFdZNADuk5jFzphtCnRb2PKTrjAP
eUzt6wKCQRidoVGsQ801Ndve35Bm9o0a8JoLFeEGgS1+TivY8H6JzCwiOS8moDKh
4iAG9Usu1DQWSY6eMA4JPaNs5dNrjetVVxH6EaPLKlpJD3J/6m1iVGtCD04SEEU/
ScfRlv34sOHdyNtovoQA7rLsWj/nwcWf/3EflzAA5XFjXsqwhFVtbA4sh05LNr41
Dg2rzUwcwgXEJB0Gc97+kLAO4Gv9LkXIFY7/EatEz85CebIv9lYjcslJk1fNbSgX
LRF8kE92oB9da5L7b9lqP2WXxcy4GT5PXFMa9CQurDN2WErmTjzD/4204yBgrvhA
cFK2o+6pdc6a6eiHXrWrMN6eoEid3Z5dxd2xo5ReZNDrq094iinCvY0uhXiFqKq7
7WGwZWu+naVF7VZYqI+n5/2fFwlCDlesa9GStHtL31QztfzDi7NxdTzbcOIUwE3i
pf2z+15TYl3RAswY3Y7J8rqxOmBcSiqHcegHbWciOEIoYIpxb/1sWDQk02XAeF++
DftJf2KPguZxBX5CNAToCh17Wp/+PJJsSUDnT6h2FH2QLjxfGmRRE5wsam741f7z
SAN63zwp85A7QoRlWTyDPDo7a0shFDTgSGPxmIJn1cMbEC4XXID5f8guFFl3alZp
Vr9ec4N/ovxPjJNeXna+sdrVoXOeJZ72Wxr3G9znTIQiUi9CaanqQKotTPNaiuVp
mVwKjcHhOr+qi9GoUeQmhB1H0GTSwTytItsjwMeANSwmV6gyAygwFmcrp6FWQqHp
2ioRST0BxavynaHbG42DSO+x0p+ViZ6aZkuvTFROZNdqBVfUX+O7EGPJYTmI8+bK
azxAJIDR58sfY5uGx0o/oiHjYItc9gF1BdiwYICtg7TYTdIVXY7aBMWUY6qMDZPD
JFV/QDyQalqGJiyjOr9L7LWebiebZ+2q3/ij/Tin9+WQNKJj2qlsTSpkqhcyyZvX
rLxA5RW0hJTP8B5bxb9vPjtFpsgJum16LmECfg9Pdo8rBIOWKv4M4qd68EfCRJ4N
Dk9QiCrYKuWArtg3u6Gr5Sgutj5UUPN2af6ofG+4rOTFBmnIx4086ZqImWM3rMMx
bQ53JE20j35+iAskKq8H+OBxZK4lknyngFrKvykPuMeyaLM93j0oGdElUJG1TojE
vdyt2mAhG5iGuIibcNVimSeGpTOQp8k8yF+wNqDsOkrPVOMdLjcuXvpAmO9x2DSP
jOz5BMVZBnGknDMMPuNLSjoYXQMHahooVAhncZ+pLyQa6gf1vO7Lw7pgOBduhl0+
Dy95zOaH8RkQMPbzdNQUoiOaDwfJnAjsstwtyMB9cNXeQYMGG61PiFDQs1z5EQ7T
aPCsQ3Uu8CyFybTTJyf+s8v2D3zJa30wCG4Pz6zSnf55CTxicxjNrQhBnnC6/U1m
yZygHROcYNda6fCkTC6dW4LgbeGOX0FwU+Yr4BkK8WFaNnt+8emjhDTEjyPkdNYx
BqS9MEamD5dis6xGhOyBmfkrqKBPdXkOw8Ixt2REYmar8mr/Hp8SMLu5QvIucv5Q
2Js0YpCM0htfrzO+BLrZWf8fqNLMueiZSF/c42RsvMg+7FX2RZazWFgj/XR5zbra
IVF+MJKfaKTHdXgH4W17V9xw1cImGekqYL1Q9kJVRCKrRtXA8fcS0gWTMVqZmEKc
ACVSJ/bAb0EGz92LV8XlJcqrwf5qbnBUSGvzL6tLKpiUnfx+l4dIhmvXhTR3Pgwo
la5hQhyGj6mR/Mmkfzo7unqvBsAYcb0A/2h83RPBJd4WIeza4oRTe7VY6DjbEBrm
FFcoNFzLNhLvGoMwj8fkE5atmgJsCdzkez0R3cq2Y/wTjjOySke8AamE3UuSjuL1
K4N0mkcwyuuMr0sDf6iP3frCsj+3dLxZSwJDFTIu6VUgq/4Yoyi07TUSsU9cPdfw
0GcYBkt5J7naaDZvkBQUeXPDGbX81fDUcdBbC8z/DdTozQ0C0/GHP2od66Er9Fu9
PcbpwHgkMSf2pF2zutvaxWcunDfRkdB/fCLmLsfLNHKsXv3n+WKFfPBnoE3c8Iby
vbMoZ9g2uaJ2mSoXE5hZBx4sP4e8ZzT+c0hyqWL7wjZZQSaqk5kLTEb4B6KQ6gXW
YuFZy6ljeH7snR8caKiHzjg+OlXgbLkSrgxOiJVtg6wVNZQm5RMvnIZjfGRT0I4v
dauTnJRdCd73IfJMJSg0EdZdkYJMR0Q2Tfkzz6IRYIhz5z7r1xohn0/MzTS6DTmS
swWRHZfyM5Eoi2+lUbvyxSNuBUEYeOZaQoqy0Vvrny0PBxgGYfWknvBMvfybE5zA
y52l79UJuRZk4cfxU8ZKAaeArojnt1gLho4mI5hf6SO+v/R6Lfb5Y619dJjletAk
Klw48yVXg4RFZdDB07fie5WJ0u+Qhyoy+HRz2gkn+O5zsmOjTdUNavoAZ7QjB+bD
2/dGQDZp/HZDhqaa2mgGs/5PnUmZDenJi75htYidz6m//+Pejxwcd366Dm/BhVpB
fF6RFQnhrmU9OV+yVV4rLoEBPUyegCf5dt7zqj9kTz3Nq2xkijeG2F0xMhGmTqmY
cxniTDSGa+QKiN31t21Uh6J382nq5UadYzDD2LsA/yWDOIpecoA5y9FURp0fPUHv
OKm7nSjEo+sA0LCU44W1Z4wd/zR0Q0sd2O0rHTYMql8G+W5V9ORV4k1u3MnCFBS2
Pvvb/mwEzvyiftKmBxvFDkJyDqb/AKJUqL7wmpiYnngce44szHttvOWIWpTTiMVD
AjcKdg7bwPrkOVx1n7bmtra9Dos7VGKto9AvJT98K9wtcoF2KqVC0weU4Qf3E0nj
mk45FNxQvCEWjwt/MBvdq8eN5Tgmb/kP6HZJBM2boLyz9IXc11kel2yQ9LaJJBtu
Gn4E2/HfnFVAbWl0chB9/x4s1tL8o/tME3yioIxpT5JodLhzrewaZUiZIyMW9cP6
TkRBF9PN2NNBDJeLHMV92BsMuZ3JsikaCufWtD8TT4amoqb+48R2lPE7qYe0Q0DG
esmtdPs7V/mMe713RaroqHRE8N0EK/gRMv6LRKPv+wKn1YVucmy0vhu0JoFPCoNS
ILzIvqWmzQUchPjb924GYNR7sqJfC65HYL9f79UiH5EqGeNCpj9azIljoJH8LWZz
E4i8iURXSL9OCEOBkFyTjKg89mLsutnWwVC8lhRqb5ncpOFiOiFdVSby/FjASti0
mRDJdIwX7BCeJ/O/9vTpuohF7KLC3D+QO2bdiLwoPQit8fHZchJMTurar0wwz77A
I6y4vX47AfAiAEXLIRoPY9l85+svhI76F0cSCNCLhQmBLSjlRVyQ8YxNg6cpmuRJ
k0a0jdaI6up1XhAH/SUu4YMPoUUaptq4eHhMn6o7eqjL7aLKhMGbIMiThusswkdQ
BDgKnROSNcNY/m3DejEm4Ep6MXxiKzHBqVJvaIlpNCfP4op4ZKhS/au3OwExz5i+
j6u1OBAA9ILS05N2JFI6A0OwoJJvFHr488fPy8bQd81qe7iiuzVWUWXE30iDh0Jg
G4ICARe0lnGrhp57ox25DcAPDfZMjyXqqJcVKkexUEFvGGpPGSWUdOBrgPnTBGm6
fK0NDmkFEnIdk3mc5MiUc4lpYC1mLG3fB103aQrHuYfA9EyCpR1j3zFc/zdykHrt
+q66yNIxxIEvoKudu+yq3f7gfjpAV+kNGn+gmrnWwav1TqYu0JOEErGewmK575y6
N/Mm5w1kMvNDzF3cZyKh8ohiypMo2BjYBKbbrrIhHF7haSy44gaYziPwU1vWyzI7
tcm67aVauugN+WkiubgMu9p9VQOXQXvjyTpbrmd47mawA0QbLDNQpzP+TJ/Ps4LO
4hZxOsTt+Ob0WzMKkrGKNtkc0jAKJZ8hN110lLgn63OX2fm9SNumUJysro+aCMdX
O9AlcrWWtFS8dBRc3NCGhTSFHPntlsTCp6e4EuTJC7DPYYY9Ksgzs7at5k2RGYwc
6O+7/2B4Ns9BFggPkvMoU5Nl6oElshsOaDz7aPJ1VgupTJiRfoGssCc03v8s36P0
P3f+YnxcuVTixn73Jyo5+lDyefFtNyz51mpAyBC0bQ0/Vc/9BbnbOf3R0mpa9CaE
Z7yERoZ/KXN4nVEljUay5ns7gLBWgDfMRrsORHQBMOJKvcCArMJBXxMV3uMUxXAy
XAeG0TfWaIF0fIcK1ghycOhqbH5zUC9tGTiPafFFfnZe9sKw4p7IKBdxWLCzwrTs
gXkzV9Pw4uon9xAPvg79sBbTao+YFCth+ObnpK+7XovgMKs+RpHGKoI93fBlzuaJ
0cMD1MnDiX2BhY2dRBsRMa7MrAMJEg+iSpzqdTAPA8HNux7AIz7xXahW6JwNeEzo
HpMYXofi1KkK8p26P8vpWpZddjSSv8wY6uLOIrRGcdHxxZc+Ni90ZZX6t4jMwKv6
U2fEBUwe4fCrBp5bg3PD/T1ItT3UG+DFtnuuhRdT6NaOCagWP667pv+Uh2PGhxYA
mN72s94zcJu4r97LspCZNgpFg1PVs7L5udwbRvYUkOUsTRSTOzh65pp7Z2Ofdq02
rIElQjKOsZ2t7EYrv+PEX5/+pscoAKKAs5Nc+qeJW/AGZ+7K+ZWPu21XY9DEd6Zj
5CBdh6O9tZ3I2VYN1uA7okTsOwAvZeiZIurosNh3/3CkJuurf+XRNDjS+laJmQN4
xAYL0wM4B3Rr3ceWxqE0hnzLf/nJVNtJ7hcWKU5OGs/eiibxptM+XUSGZaAOXcxr
fb4BilixD09sAt5QwnIFs0lEtAWULpI05k4A69tI4CuJRNNG4CwZNwZhPxBdp5XS
h393VQRR2UPBo4Cvyzt+AEO0c1p1JcrTatH1TNIKYX9XU87PdKAHTmvt8PazP0iM
aA8kHmhxe6PjYkJSHwYMpK77xwO6e6OeBa9MbVO+VaAcl+qu2Mk2fSguFfY5gQ4F
bWRxVViwh1daCog7EDpz97V2HoU3ycF9/Xs5hQGFTghW/bsKivoltx0Ex7usFMni
vqKNoe+VzfjlNeIxX05pFd3qqZsthUnPWXo34bmYTRRwlQavpUeddql5BmNveIgi
Jyx9RCNGMx9n+uMwtyZK6Z1jGoql6Lb1hoGrK0mBqnuXrD8ZwUxsrmrJzbQ6Ft/E
GflJ7vZuRhLDvGs4Ve5gmyAXvOJNMO0Xn3PemGkSl7Q240fKvoNPPrGsfDKYTZIe
5PZBKXEtfz4ONsj+hZxNSrY17A9S+SwjL8g7U9q1wH3BxJNkywkgQ3AzGp4onYpi
tVXBCSmMh+wt0jJWFxL9lrsggBD4sP2rKro151Iw+4lRR21NM9n8X2SDjmPuC3cS
PuTuaPu2DmMcLLx75rRQiHNuQuZAxADyCnc6j8fUb0xl/SaArwnuUIf+Wl9i/B0q
mjuAb7PsuVsCGC+nDShLJIsV70IW8YD5fJRLaGk4+/QN9WhTUAQgcigNQodF1Pmx
BInPolgzWnIYBeCyoyS818PgLXD33uLdKJ04xTwOEwqI2x5vGD8ANYE6EQIvCnJ3
Tl1SFQmJVjtzINUA7MiS0cOoBVEK6KRDBHsUABF7uVGoejg4BvHFzOkkeBldZkW8
P8E/mW3ErPSTGi5W14ZPWMsCjtQlt1XOYN+MaFAvd092KbhZWnu2QVUfJyso5zPX
ttWNxu3rsPb+pwbDH5NOA63XGAL2skHqtpwbGyC68COWnf/NMDWc8y51jNj7oUgL
A3cg2w1S2OZaBpOmIsBFeFs+dLlcSjK9cM6Voq6bi38viLofXKjBin2cJI7bkGMf
3u1J67DC0bNUBqC/bIea4bOQcNFOwgrykvH+hRPd/9C6Z5e/z/2+XkVrDtrcICot
tALDzZv68KeBhyhwolyjHUX27mrPWnX4a/gkp0RRjRLabl0DffFhsheOfAJCdD4z
W2PAriy2HbGi/GBSyJ02U/g4R6WbU4bVxM2ahlSWWDIJapMEjBcEJnb48RRfQdou
Sy4G3d0xEFkaxNkV4uq+HWrWrEGdsPkmVpdmz12fN/orA9JIePVCzQzNS0uTj5dc
NJO4rKVM3tXKTB+fgCJV3yjbn2Ove8RQTCGEO2UY3JeEfmAU7m75I2K5W5UX1gMZ
75o/Vt/rCz+GPkb8FSgCwsZWQnzbVFYsoHVYn131aarp7nDrZ/ySk6VR7C9zRQ/f
9WOjW4fJb0U4h2HsRC2nxocJeuqR0T0k1u1/2it3BoMSnA+4x1eETzxozkFlLaFS
MPclpbp4avIgvOGeUTHqkdyB1OqGJCnmzvTjopuLcF0BiOvGiILUI7sjSy9ZwO5c
WCOZGN/sXkiAm8kfmaG4/eMQAKRBeAe1ahRTwaEDEmaVBDq//8MW4chynA+HCXnM
rSejQf87yNy+tasVEJA8RcM7tudh6Lm0sPuQgtBmpvkwffOtmZ9ZCSQljusmCqnj
zkIXmQYeJEG6QcSqfX030KVKIQw0hMMTb1vNT3hFZSeEBDlPaf3y1IZ6Dhs8WXei
75qbHOJnKImDoT0EUviaIZYw72q7rR8ekPQ4z+MtZH2+sTD0sYmJycErUTNlXTd2
6qagxYdd90H6p61PsU+1am2JsOuX8VsBwhoYoHlmKcWr/+SaoJJda/QSF8rFop6q
P6axhPwJbpQkZ20BUDB+qmCGcUr1TnaRSULc7NzCD1Uc+Z8zmfFXtEefLuZ6b/lB
HSfgCRXENuxcQ616RaXVjO76enORVb/1bDr85qmduMuGXBT/ns7n0mGME28hRJmx
zNhRoobdlOSKGcUdpy8ZYzc83+Wx4iOtQCEYuvR943cKbbWVf+CQCvpl+gMe+NzH
J2XscNRkn6n/s2wDC4BuY9CXWECzKxYQkliVn/bFt0SwuU0gYfWwElYMRaFj0cbx
Oea8cm6mSXYC9XVWVnQ/le6kFgp7+b1nCYi67Nrw5qEwWgQ6BheXUofKDW9svRD6
TEPgmwMJqEaHNU8aYKEsx0He+UNdwaIFSKSPjWQ1HWWy7DbBXV3jbLOsC5KgyGDz
JIZBpJjW5lcnYnyQZH+AcxRXsLSKMHhj5ykc+bfXEoLUz7G5tVxjtGCokaYK8+3R
W5eqvIBft5WyKBCoFiV6DCsMqpIulYiqqJyH0/8I11kJ6+qqUbu+PdzOTO3a3SLD
yI7TB5I97rytSWfImURw2fHk4qcI203bOaQi52ZAsCNrbpJ+qzPx0YQPip65wIIS
6WyA5162uRhWwCNHCOxkSGlztaBL1n40Yd9G2To9zjKxXSnXUi8qmPxeBHxUSxpv
4tLOfgzyY1/gCU0erXD1JUp2PsJMm58RHES4Tbk5RydTVXRbF1hm5HAkOGGTCffx
shs+fnGWsksq5Na44ixILsDAd8fpqkGXSh/cV1DbMmfQJgIHH3cvhP1LDS8OV+zl
TF3irIQVCwr88wFf2o8Hkopv+FMhHy2iUZCiulT7njIoj+7fcfVEvuFkf8gh0/z3
NOXeGioQkxI/mNCipw0b3M6wgLVSDz1IMYwZfPe2S8E+lCcI3YiR2Weox1vALWhx
bElxlzaDqpSjX0ruNiEidIYy4LRX4pS/CvrpIMQ8I64MuybnkPiOzK7JFEK/Ypx+
0dO5iY68WdMrf63a5JvSYyj/c4TbQVGawVgNPsI3Vs73i622B3Oe3oXeHKaGRajn
yFA9jMmtFr+oNMjS3IlPKZWstbjOqUGHI1Aed2/O6bbK9PgbavzaIKXLkDEW2DpS
6uo2L9lqFS3hmKjwXMNPOvc9uIf+ztEze+jsIchs6AxVO1DeGXVzzr/+PF71ooSJ
QzzjcnV/Hv9KdmTjZEos/74nSVrPPo7ltvYmOeqNwwqJgFI/syensDtS6UmtTiIG
yO5D+8v8pvfojbD5qYJ3Dny1mOZbx61ryF8IXJcUqyVR/05/otMkMsuNH6aS0WKA
CjFXTeXczkAY4fa3i7WYZw/9/Ts5AuNQ1WPBp465VvxuTziwKlV95g/1uIkg9SeC
a/H+Nc139CeT/dbMESpypBS3sjsfvmRjVxZsm4KHs36qMB3Cjx27Ts4OpIwfvsNu
5Hu/GV/kWDT3OkNzjiLfR0LYQXnyALvj+y/Y81ZYH95E9wqODKfrOZL872h4oSJj
JSLGg37luN0Q3LNjDrE0kDcl7zn9ZwLoEK1eOntJ6KichhAJGdsntFzk2wzzeRgB
Wi2gRUrmzZomzNpSIEzJDdxn/q5tfWufdJX4bayYBydxDgMsSSo31lJjlxXeh0PV
SJtB6zs3Z+nfhyLHcAeSsUBWnGs6YfmXJamDSwyGdb2D+Wfyom8CxoXHvPp+zx7H
udvpCxwkjTWGRNdG0Ym2lZUbdENmQtzbxZOH/y7uq40NGWLItCffBY/JBcz3bgdF
0zUneNkDnhKUBbMD4tZ1kbVra8kxwtJipa0xHDH9VJ880U1D4HIdtG6PuVabSOic
5fUlkfE7NyBhfeBPr3QVHbQI2prohc5hGV0xvtI1/mOuP6/QRnkkjRAqVrTdEZ7j
5Xk+WYCeJwPNSowVQZbSDQuC/mZ4yBj2p58gtl4oNFzxNleJOeTO85/HZ28UP1wr
1BpfuE1owhauQI1I4yYNvXYKAGG/uagm5MXS24fR5akfawJhPCpjg56o27iV1j3s
HSr8uTeKqccAtppOJa5cxv0VjkjupJ4wdR84xjbEMxYNqrMh/O6n3UbzP4qjKCRh
d1nK+V98JqoICSsZOvcLlydBIvhTUVy/9wpwl/dB+UfjnEJdFsI3ekhHBQ5Ijgw8
6Ktqy2VQDfQG8SfGQH4WgwlKKYzaPHdx0u4fxyItUqjfYmt0+lyHmhWAgj8LW+xD
ae3npiIcq1isL13zjwvu1z6opJWn/2dUWfUuZrFTHi0YnZMCncof6yetNuB5WbNb
1/xCqhBBp6KTX/bHyaxOP1NoxnBe7Pz4kVtgp9oF/B4EPKC3dBwrY7ziKQvFOHmB
otbdY6QSOUQdORaY2R0Oxui8wKgklV3TbXWHize5EWM6P3/It9Ol7AEr5/KS/P3i
oj+xGX7ws4CBwpXP9OP/aWxCiM17YZqUISX+cF4lUc7zZZ0sADf//l4L3S2899jv
pP8VKJeiKaj/1GHZjZmQKpRn/2xf5SHQheEHul+cOiPihVa/55Ww4CtoYYqLxk+G
qewPO6tcVX0PEahDfZY2iuweUSkPBBO1z1lhcg8wsaIVyhmVvpxejhJgQBOJpRlS
nZRIxbzr5aPATk0lzIdJczCbOWJOXdOhrUj/hpy4ZvU5FK+NHXh9H1vqpL4EgRF/
4sFz8XmkEAvQ9XEFzUvf2heG9MrFIrUb2eM1KEsQQG/D0W7yqMWaNwKtgJseNlKR
cRzaWlgGNDfTw+QnX7shfONT93h7AQRpbimdfKAzChHaKAOe0INqXtPoOcBuaPTs
Bp6XoNPYM+GQDaG7+qyuYODxMMrxm4D2SKMtfx9fP/yx8u/Ney8eLcIEEXoh+0U+
xjBQxhJm6qKNE8m0ZVDuwghdtjVjqRiBU8DCyzMQ4FYfC6yZllhhIWKxAv5Qi57T
iJ2ueMQHYTX2mvBP5b93GM3qdKrrkvgclkqud5vtsk/m8te0Ijl5j1AszsELM6eO
TTqziod0dWJEpQENXoCE9UzE79kC7ID8yOQs85zPNdKS+KBhTIxoREBQoQ0YKy6B
JC72b1hhkfTX4OWZ5gz84oehz0ae0ZJmFpRRJ+o2nNQva3gJL5/H4OaALBXEyP+3
MYeGaTzvcaGjZvGAE2q/9P6vD4OKJSPGPfXpErLRiMf8F5PrGPt75ODEtm+Ehl80
SPhhIbvrIHYXxZiByN095Gchx4p+YxXt0KlhPjKKmRTWzW+VWNAwIeb4vPZ0nvXp
0O9P6AYA7/aXr1b6rGyYvtOLmMAbRAsaNPC/Ws/iwSMwwWw8B5GI6d6uisb0E+oQ
628EUpqzlAXUX5AOXEa4L7FxdZHa+8VbFPRGbJ0+1sw8ZTwF0wEBqhj+h3V9+sMX
K+mkEJOODG/zzw1RHDnKhJXGpX4ir81KgGNEi/3vIwZW06KQwHv25VC7W0bG6eqz
pe7eFiFRI621KOBOIXyoPDHI25/u+pczyi1Ji7zDldwl2dHmg4axw+a9eSzjEt8b
kQyc5VA2gI6+rzV9JZMTx4Ut3HRO9ueVKin/7tL3sWEvZpMsZwGZh+YZZo5d2Bin
X1uzJ/AySWYjjsvrpQ+voy3lkklJnVnmdVPaRIKejuphIOi1Ke1p7JR779XCsC8K
sE5xQgc5hF6GJIXJoWduKXRpFB9q7UUGlDyQWhTVQKFGHzFpcYxW2/yUdTALx0kq
vB74PeyO10JUhKpdT7w6TdoOxURuP4RWRpPXfh2EXrHJ0TzhqOmC4mZGwLi/TTZr
RqxH0ic5gZq+VAMbQS/rfdTSYETSfWGhY3koC9BicMijeZwsOuJ5SKoy+4vbhMug
fNrvrXhnsGAYj8HShqrxgaOB3srYYDJ5kbJ1bqy+tLHJtWUiLiiStNzCFRpkdAR9
7iGyf6NsF+XVmU3ixUx9aMg1jBmqZWPLlrWb6QxUdWQ9TYT2l7Vc0KNs9zhlnjwD
/aSj36FwtUkNHlzoYJRphZbTza+OkkwliHiupqNr1oKvIZ5jCxzWr+K7K+X/aCUU
U5n+XABeuodxhepKm5SK4Vr8oHUf0FSfGre63KToqz+Kzljfcxqbu9ih2JMCbMCV
1S+Yo9EqfhX1DPrW1hjCRA68KHsqFAASt0r6k+/nts7aJRSlTGtMEryrfrCcIANG
ErBHGd33PpeKDEesrTCg8fmVH0KcYhHxv2bAanDhsts1DsVse1+VeATn91xyyhWu
+exPVWq28IapI3AlP6Rf+M701BbLedDgJXqU95IKf/IFZsZfMxOwD7mzfQHTxaub
GbK7Wby3EmdHhXbuorMTNUUrnQ74geFYb4ngRv/f14VY5PM/LHc8ZwH1t6egNKA4
p8JJYFgy5Dxlj6KsdnV61Y7k6ZKJAlCwAIxPnL3J4RcOUC6n9NS7JNIVcV3OcjbP
Nm5AHME6teV4A0RxKhliCJ4TbqIRQ/BsTPyjm5OAQp4QlOxrcomI5Cvs48OsB1S5
cox2aNhyTPyk6d7FO2tYl0qw2KAtHAExA6vzvxKcgkxGE1geT42Laxs74HrqBwP3
ZtaGOnm8xdmMrGFIf8PCqKAOIz6IE41ecXVlbGJVaV6Vgoj/J44SKeKzP9Z+X0B6
ZGrDIck7DH9oObShkKQo5b8DeyMSOwI/MgeIoQahBJeRGy+gXZOBt9u/XTdbBD9s
1c/hVJUlsa3oBm7SIvXEK9BrV/8+CkX6+qLxJYbkJQpLOtb+kBJ0PAmTgh6k8Lf8
vhwqZM0MK1lMN+ixiPNsRS8lN/5IR8Q5ltLi7nMEOCWHLj7QxriB1b9LZqU/NXit
jrRKarHiNRqO7i/E+iOkXgMNSeAYRRDXjZXOxV3EWvQLd3LjeJewQ7lVC5QpGVIH
uZWtHAiP+8l3sn0sRxWVxFl7wr8WYW4MtmCyqFOtA6v71aLRGckX5OXVmkmXK8BB
q50zc9MeO8dyaLW3Knlc8MpLltucDSGvnmKSxQqN/VCWa1s8DonAddJdppE9FgsM
B/GMuPwdmP8dCZWstXdmF6sKjVdPQwav4edeMry3J9AnWs6Rb+jfQveIfsUJZqJc
OmcI6xbdLwYiR17ar0hjw1Jl7tsMlj4DsaKfShOBQsv3/xV9puEuWdLmTZZ7gT+j
F3ZPbPnCyRQ+iSg9cxzhNGxtj3mbAhXFXlKiq5jiyKdb75T8YNljg114OT/BID6X
aXG0J/l3M7S8xME+3UeKyV54DzqKumJqOf0EADoojrT6qr8cpXufOLXA55fBAIkJ
gk+u0bRqZWiYho8xcsBQSjPiiF5Qj+Widd6tV1vwVTkF8obCjcnc41kKq2TfO0p8
kHcnn5GAauaGJ25cFvWxkXFqQzpmrX6JF6Dho2otCxV5H1COGS0sUU3/eMywlq6n
vehqKLgLyebJLwE5N+PA+A827ytT7vkH5YvhAt7F2NTANKvAl3lUttE3Vh6BB5Tj
lLHj8nenZJPQvNcHENtvXpXgbKN3+pvwz5RaZtsuCv6k2j2ozfkhxE2DKP2YTJWn
ejFPe12hN57m1pQgiZ2u6NEPrZK8w/AJAL+nQNVlRhTaOvoqxr3AgZqqqefy0iot
F7AEPLinuAO7vG1CtH8Uq0io0n89yvsecf+86WzABnnEgC7lqxV+CEDcF3XVi2W9
pYjsUYLfatDeMuLp+YdTieTsrIlfro7vQpmJjo4Ibl/wxuztWgsp1bxsT5Xveo4q
WeK4gqNGMxuusXxH03YBM4S4uoMvYwfbURWdJxWD8VEV5cLJqdOtTCcilIs1qaZV
Vrax1A2sggIOVDh8hbJl5wq8bFmKR7FuxSWFROnCgyNlNNiGDDWkUglOD3Itz1kB
qY9lwKmUDhghXwqrbQQ/1e8/bzkSuUP77ifGUqZMXsGy2V4jEYCpTfzY11EEWl+i
bU6lLZO07o4kxTsR+rURcbIl5vxeAovyFxOyanG9fFUjAUwxlbpLpazssG98nrQc
Y1PUilgkvuIIJd66XIXcxXmagw/srkrh439Y81513yOsiHvanYT3HHhz6y6Q/fTX
oOFHoZZarYDmaapD2jGgT+egKBPg7QD5ud+g9zZNCjWjo1CWFxHr3uiSOlfsamMt
OpI4aojIUZiOPBeiiB9JD6AKlBzIljEKUDw7RgcmdqDq13zECcCFtZNgyB3KPaYa
AgHUNrp0xhdD0h6p+3LHkSSSdXUhxBWlo8iLEAwEi1RAmxJAFV1tsxwhvjmZKl5T
oM1hgInXfaltUYTWphey48PMyezRoAFFvdsyprvhYaAydH5K2MkfcA7YenoKruEh
Iz0LjvJzzCWL7Q1eYh7wLnzc94OtCXOBFG4KD0/qj+2iuTAOq5YD+0S1kgc+2Mjh
MWFcDSbJ8OPBBYwP2ZxwjCl0Nj3hvQ8LTP/maOMTcB+uYoxPPW+s/mTWzlo+aNx9
5+AgjsKTdZFqtf2r+AA7SWCbzSoP4OZ+fsi2Ygfm8xzD3WZT+/HX1+aXWrAdWI3S
UMzDr8jCWVkzP68lxVtZ/R125BRQ19ykeDLaT6vSf7NywHYiWMHhHmC7W3ZJCLDS
cFI1tSkPkUyiz7rAdJXI4C4rxB4vilK4FgBZO0hwgxf3oITrDu0Pp8xv57L/QEcU
L9IzmyE8M+Xs7yswQ04IdUuLqGZX16vuz7P9fYBQgnUdJ0TW0TfJ7QuzuxLynyPd
3nEc2Xq2qmtJ39E5uT0YdLq0EhToPPguxnBV5FzHcMaoHkka370ab1yKYNKSlOYi
h7LAElWLzVE6iS86rxosyfeURk+//Ut/2rR1Wdpyl7fB673FrxavwIrrtFmCwqn0
Qtlp1FkZgDQrB2iuAcwCg6jd2xKQi6RJLbQC0q8VoLpFnZkcJ3RxswtZV3rr451Y
kK9qAzUnqSxx7DCo4FeryHErBYs0rJyfCC7drnLV7mVDzPr/9Q/H0TFZwVv1huv7
JHSoZb3l2AD1duEoLwHlv5Bw3aQieOpU3spKF+6hfV7Q7IFz78HzRfhViYiwVUvI
keL5eX1K1+3JI5soBGCOv659Sh3yyeh6U/yQQc4RRtbiqqL0UODuGmb58ZzzBWv1
C2gnf7oj8V4yUlftB3m1OYdMF+hKMxrp7DVeL+Ypkda4cI7zYWvxqZG3aVPW7ffk
L5NNlBKjK2YWujf3TiRQaDCvkTzs62rrDuE0TWazEV+htdqaUozPWaNkvkxVbN3p
FDbReUB1v5IyJSv0H2kZaxjqmD3Q46uANsuSha1kQe4j8e7X5vESvj8Jf+p9yl6E
e/ceU5mcpETaYJ5fqqi8ggsTo9CuV219E1VXLAFSXq9SeUmxE5o2xW8nUUNC8SXy
nYrgMdojj+TJ4K5wZuS5OMDhZSN/79KmqYOqUqVc5KRMVfdhYij02f28Uqd2eVb9
oHDViN4r+i3cpNS8WeamqeQQ0GKvEVRf19bzsiqt7LEFztx/dVjKDlket4NxoDm6
pLCOlaoXHiwNlB2Ngt4Z5bYsINwl1FfkwNe/1PwYoJDtYOLdptswDxCoWrlsjs8K
Kl1T27klUgWcspgWcxpZQDuChKkIrsIRUCE88hgEjGe2V6VsEfw3SZ3kZIy4j7UV
UchDRWiAs5F6hYVaQfCilVY6DjsT9Ng1qsMfNxc/aa0Ac3kHrYpGzb7WNdta7puW
IYURpy51QQETuc4Udwz/3xPVwcdMYZYoYObh9vc08q/DjDRgBW0yA5LbY1rwMWns
XFY+F3wl5jGHwLUFsejA6VSJ8L7t2sWpQyvv9kjXsyMD/0i67vroSEZfqa6pd5K2
KFhAd6u3163ErdXOmD7CoBklpGikpwRXwRc5F2SWVeprh2ntA2RLGYWcdjm4hm/q
iv6x054eEcRIpGla45TvNN/pvLUctHxQHwPQiWeskIbUbzvrdB6zp6B7Dj0YCjzA
lIC6x2j3t+4lSMttLC1ePGT4/cXMpWOAt+vvXHlT7gxp+KAH59/5Qoga8wo77nJi
KzPSeKNOd56GnOc593z8pUddEU1IiXpgwJWo9bAI12kV6nZ2Tz/KIzC5rgvXsO6J
BQsp9T5vEYq5LkIbFEzJJGl3jYbDkgRYqZ7ZXdJHFM4+IVeKFse5JL/1DM/puskM
muK79W0B3f7eG9w/WlJyG9RHczzZiQJa4o2gvp6tB1UR+fAUxCvoafd/UJysyaZL
o5ALQwxaVuM4Fw2kn8Y0Q6CJGj51/n5Zrme2FsIVmT+Iw5oBYLMndQYVF0WaAW5V
BNxnGQqFhihqNz5W0WUplxhPA9i52Itg63VIH7MpUVp8CISokBsLEDrDJPhKgVR+
CH9H/ia1DgAZX18SSc9luMIrauh4euqsACyxJs/s1gFw83LLHfFfvA2chuKeVqNf
hVvOVXOeOJ8+ccfne8UYhhhxwiSlPNKhhj4+Z9WnvYSX3KeSwpInxcYqMfmRJ8tN
keDcplOhnVGarAa0nRkrGRaIb8yc5AUQ/REK+fBJ4u03w3Q3i1wr9nw2ro7He6OQ
kRVC6MNDv4WlN5+Ri7gi/34mj07OMoeLhGj6oSC1J2x02Dxe1dItmsKfNQsIZoHK
eSPk2JJCGBsYp4V+LIqCHUMzW5yMzAIL399t4lqSNsDNaimbCwnms25kKoz63T3p
MHwTnqvxIhj03nhL13jntIo+Pxzl8DCBgy1pCsfu3faj0YhBwyJh+ZuLkYq8BOb/
M29HJksjnUD6oJLE3RDts7a/sFsX59mQuy2z5LyD3v+V9AEVEv0rmGv4om8vFnKo
t7nPiKgmer997Ze8MzUpc5XPVqiDw63x4/RPqZMZY992xl9ppuT1HdKXRAE4sYk8
VEUwEnuuiRgIdmkIoK+VgAlPX51Die0XbxTUtPkRuda8FOCiCG/ttuz74YNuf2/8
YrGJ3NkGX6gx01rQxhfg601ti8odvjAs82C6aRfDusACGgfozZRMniy4exrCZMl1
zjmJMIzOmugDEx4s+e3Ghb0Lpw0aCHaOSG6N8GyBL2Mh/i81oqXVNmlqG2Uop6oW
YELw8xkcxSbsMGj/t6sAFw4wDG18CTlUppYh2a53F+LAq7edylme2Ikx3B+Vb6TF
3DhSuuAXem2nl8c9QRWoNHtARsTg/WtLxzgAqufBESs5tsPxtXYhSkFSpVmC/+UQ
wrfusp4yJyrr3rY3sPcYPFJU0/TYS+Ch6DF+YNpERrnFO5iKwTmhz85mQWuFzY6x
72Ov29vS2mpoidFiQCLjEO6Vc1g/mayVJy7HuzVkjSrWMP+zro1WgX7i1+1JEAI8
d0a/DZxpP3d9armyv6xZnfZLXcQcyCzndT19rAx6jtG3+HW/LdKdVB7QDh/7tQoq
s40Wnx8BM2Bvk8b1L1DlY8VQlz3UQTeFRPUF57sonlZOPauCqwcM5w0i1IQp6jzb
YSNGgGnRG4JzqjVRxR9vbwixJ8YyAzJbvTEVj08pXMGiJ6u1nXVVD81tZH+fDc6u
wpQyzYHLf9myPS04xtG7gfQblw/9jQej6Thl/qQ1u1sfcoUfGcMqKa6/w4ujwkyR
m25otXCEjlVvq99UWNA0kIGwFll4M89wgveWOnusTzkGkEBWiQ62JE4lq4zYyoA0
xEO9/8dpgI6ibIHDOWMGUdt2Y8BVESp9B2p6wSz1v97931jF013GQdtkCCTS4mP9
cloklB+j8SVnSH9w7hLrhjlsZLjhZbt1Y/rtY67rLni/M91FYZsua0XxaiI5dJkf
UsV02x2RNnko1qR3mYXtVxWLp4qXKsSXo4K/XdtArMkNfvtF7Nes+HJmAKaz57X4
FcOcKNZ0uf7+4IcIGUkf462K8k8NARuppR2rhWLX3FqJoXfEn6GKBE0JruR7v1uf
hraWC4VBYsOU9DwHisyDHejbEy1wGm0AYk+wmCk5BpC9/DS2PwUGjvwhG4G3Ha2L
rtO2uXjSR/PeamSXMDm19cRceNoqXUwNgsG2HqoCU3e6PNxC8TwZfEMYpRraL3V2
QulLz/QM3zwUOdu+obqj6f6LZR/jU+1jHSpgUctNOOkpML4jfj3+WRkNTrJuQGUr
ZklBGZM6c0lGn9Tn4DRJUU9hsNxW8Brjc3ZWN7aaEUmO0V58MaSmdWx/eI1Imk/R
8u3gdb9ZCKl2NFEpuq/ifbXdMDkutXsHN2uikHEKplJ/qy0o9FTu02dWT3t9X4RH
Pz4iCozeRvmHJCzqBKOHrwe5V9/J91t6NFqfpSxA4kIF5kB6f2AylWTsPin7v1in
MYiz62WBxU7rCEk68i77jSK7CbrdoyD0467VYCDKwXTHau7gk8kVNJiHp1N6UHa0
3o/oHMU5EGWMSAGXouRfOeEcnv+Vu/t8NOytU6m/zx0brx9Mf/bpRdGkpFjh6iJn
QiLKEwkLUuDCoZU+1xqlDqgHzZ2FU1dTTVQmcxQgrOA+l++9/c4O/8my/zteZ0yK
k2BGVZZLWMiuKojgr19WifaXAk7od3IfkuPTHSuCmLWLGIQSFWHuV0K2OHShoYYO
F3NchSYvJBKocd45S6KYuQVHkbpuFoudtKliA5/st/8d+QkmRktF10FE59B2VPd/
ar0izvdwEsHvpDSjyuAJ4t0d9+6TnBd6Q2fLE89ZGcy2L9+bAqi7hw8pzXvUXibm
mETy29afO3v/n6wO6EWDH+oHBv9EDy782C3R0P06Pl3qei1ayZ3O9PGOUo3tTSTX
A8QC6n41d8tLiOj9Spe+/NSKMcqxzSxwCT0BS25U70Z1BUdbZMqDivv7MasX4eAD
On5ztlQvEJnCwDDkD4EHtHk51sO62D+HHtxILgKVf3JTtbSTA+alJvP4qYljUCZl
3Utmwfi3NGu8jVoIxQW1fkVgJcS4YOEjWOPh41hjPkDNGUgeyLH0CG6CybIXIOHI
XLVO6fOt55mWSd/+fd1eQpI4JEcR8CVJTaO0iTWqZZbwgpU4lupk+1Um3jo+NAfd
oVvHDH30wj0/e6qmpPjq9wq1oNnaNbfXfY5qslEH7131YG5ghjtCnsKrUvOKx8Yx
6kZsTE/R1MZISFs1Jy1hD0Q7Q+nNQVPrQwA5v2DE/GzLAvn1bx0/Lr8ucCIy9zhp
rLgmUNhCkBp4WN5fg3O3N8IW94Zy0ATmUIOxIV626o3v570BO+3HDHofEQL321Xq
waqPbh/DcmQekQOcC1xzYVxWMM9p/mYYMJvihciB1hCAi4minyRcs8NqO4K3Nyln
AWGD5+E4oxg8w/Q8pscavdOGZYUaXQXymDgFh9VK9BG2qVtBB7GmpueEgouAEza/
xF4o01A8IKEnwopkBIqSS6yecpwJdx4In0Io+56irwHlSWDvUqrtWaErxVxVIXqb
RMG4JM1oKr9rBLwmBr0gGfdrhih7+byIkUBhVkQXJuMrzbFvseMrJExS5JZ8xUQE
zWJWJA76kZS4o4nQC1cpxUeSnT0XKkO6a94o0iQ8mjuCXbQEJeZuBaVMD9U89rh8
nydu0bzFqMcQj5k1hlNKrYcGz7o/+P2krphf9iFFLGIrAnJyh8ZK2/g6N5NmSu9c
PMpXkOrSKieV6SgyETZqinOjbuqWv9hdTAoK6AQ5kRLW5K3hjdeEylk6QglXWkoN
vlDP3BpXtNkaZi/7mnc5vBXxVO47crfgwIT3kBqn4fildzwMfDdOeGvq8jwIpWcf
0hqrJ/mH2dX/RI1f7QEOf7xzsKvt3yo5lD94OTxXd2guWvxGzRItf+y5oS2EgHNg
rbsOI9Iby1Ben08PdSLnRzOZQ3Co1iSgfASdxZbaZ9574kxuYJ1AmB1g/WSahLum
bbgeFJMI3vehiZHTbSc6Mm7DYdCijKytjRt2FiyrQS13Lqyx9oePlRaF4b4YXATo
9O9JR3BX1833zkWledRQz2mhhA+y0P5yD9DtSbQIAIcNkJhO274KxzVYSzj40TGq
KKNgJ307Fmk16AKpvAcwzNox38bC5iNnUaL1tJ8U6iXdttvjc3TWCWrZq0odf2gX
lTRSqTmzuaTLjMcISGuF8ygsevR3rfHoqEbXkPjPwtny9SIotT5tsB0B4YfBgz3T
5F8u1tplG6dcjqKQyqjPywIlx7R3/q8SOSUshgyM/1Cnr9noX1yU2Ap03S7ZtdYx
AxOHjl90ghYM7LDqHkVjNUvpoxuoLdlHrrUzUhp/+7OFOLOjOX/WrZvHQIjGns7V
DE1SAB2/sdXmdiECAqWeVrvsclIEfXR9D8U45MlHPWyREXsNNz+ihNKcY5EApIYY
9i4MlZi9isBFThPvbxasx14ssD+MudOOUIiGb4VvscwlB7ccMmT7cuAkLAF7drfZ
SpwhzW1rxDSCCOZoAMTovq1TCeKfm5uc+TkMLx8kdF6UloyRU8WYaL5WklWizVgB
tjyLQYhWgpE1mlwVMGwbUaAtrsa2GHwQHoz0YkPk3tBm9aZb+cEr9ejWmrZag27L
xjVNV7Zs4SmnoyxZUH1j1zqfLRV4/Q0X/pRmWTLyeq9xjfzO1zUdRiWKfCMLA5wc
1iKnvw2H1HSQ08yJ/nCA1Yn2NDl/JMGu8fnXo1hLFhgDxsVMWpEgcQ4vgoNQRV8m
hUMqfcXelScQBPl8SUZWpzsl4iPvbRfJ26QFOeL/iO8D2GeIelpJW+iUI5TLk7eO
QHVjvpQ60AxGcYsKmmnJ8iQOCgbNu6MjzOptHbR6W9PI9Jm/f7QtVDnFm1AuJNcM
G+NxIB4kTo4NKhgYLc1MHiMP7q+xuclpvpIs6eHteJC9VhCXiW3Sjy23Z3jIWOtt
WX5sG4xaqajEM1F7oEWAIMm8qIyDuiKlq+jvvXMuP3gfZ89uCMkeDTfzi494c65q
kCa8xhb6R2X8k0zK1WwbUU96G55oeg1koEpbBWVRL2Xh+H8ge6QVhtFbuYGa3TF/
wPqq8YZPomAgTtIWj77YiBy130aGgXTq4BVs0DhivO8PFVgGKVwE8/C3dsdZLnvj
eK+0rP46vRcxw52hMr5tYLl+Rji9JvOWrlxhw34uM65tGvMbt7a2xMveIOj243Vn
daEKy4qA7RdFE+8gUYjmj1nyS1GOZ4dViIuwPFAIo0kLImm084XtmtXNmdUv5VOG
bkke1oruBy3zv7cunuDf0c9ZoWqO5E0j3hpBBEPoHRhaPY81QsY0RSgWOT+P1e/B
1KHr/POUnGMob/HIza/ilzfuDs7NY7WGpi20W4hsX/sDtOkDu9qkDC/gcESOwwBE
lpQLqOKhskC1vDyzlGcv+8Uou9acmR+ZRetE+DqYGQbuo0etNhrC1ykK1weagQ9a
iiMVLLOZOPfj0IcJiATZ3Gy7vbRHtWXc6nFn12AHes9FiTp04SOWg6l5pY8/EwXC
akQUius7dArn4lw5vymz6jHQgLIcEMXRUmy11773lYxGuj5Z+jF6iBbAailr1oRP
c2inJqNxwCehUBrN7MSkFhj6dYSoziIInUm7nEfg7zA26CIMNC1mJXXqB0eko2VP
V75h8eM/ORbPGKhhS1ydd1K+FqGxJEC/k7i/iUcAbbp5ByqkGq/1lrHxUNZOWPxe
pPbb3uoBOCRA8PLGZUX9LpReq04vtcC+2YLOyEBSQZnXq6vj3GNgVq254Q2p+GTa
Cfh++YMGu+cCVf6hea4Vzq7LiGB5TxJUqhgoeWlsErOBnOln+/pQkB2rzeADCkws
QPC+MoiXHh2Up8ZWxT/S8dn4waw7FaQwGFuW4c69zST/iUbCN6VY4VM+oxHE29UG
7sA1CMci4eIzSYNkNXs28G2GEfyHUDyATRcP5S9LW9/UQh0wlDgi63fc1yfR6teg
X09lfZvraXQp01ShPYd/MybMCPg6Orig5N78lCNt+mPtpwuWSHTqU6OhYRqdmSBq
7lF/DSyhCqlU2zVxC79r6k00PigT31/V/ko//Dim9N8sYyTJljAjCbipRSr0K115
6POdGVsWRCQaUhPjGwo7dwdr5fJJ3ylflugOh7crAZDttJjXX+5RfYZotJ+w1QXU
94Y/9dF8NC5a3bmBokdzmZ7EFpwlbthNbJsEujINsYj0xQcQdxsoQMZS2xNiF3e8
5iZvPG6EValX1E07iWss/2ZzTh2MuzltoGsenz/6bQbksKBdulB0/IjW8P9UF8WH
RUU0r19jKHz3lwNMNHAfEXaSLSkL6QTyf748QOAQ2GZHsY6f6GKCd4qiWG2osLAM
xaRp8PZt1eyTCImz2UYzv3fk70SsddMT3OBk0EKMwdbLnsi046l2oJY02M2hg8z4
NaN3eEmqy7c3ecYFzyL8e5tIHn07vhH6PyFuuCHErgVk1yJnncL80R7Wy3LW703q
YHRnYnqpwgPT3Nte5luUuIF9OWUtlhi89O5oAQoXQfCoRnIYMQco4HA2BDC6J8Se
f3ybW9zKPw30C63rgy/aCSVe7npauLDaUhCFkBJ8c+mYGskQB6bjKXtJnK73pXgb
gqXIvWK2gX8HHQUw3L5+01LbU/VP1ZiDkXFywep/kANQyyrcePAhwxkAQ9txiL+7
7DPf0e0BiUCGGC56RFA2cI2MjzQ/ADCRJLfITVvm4vFHROleQJef2nujB9RdjDiZ
50Kkbkc7kZD9egZuaOFZAI2X0FK1mAenhgICMI3f8ltmM1jv9zmwqnWG3PMV5pD+
1YlJ26l5Diz76JyjCxNwqaboVSQ0Y20uQtQw2tdsivNwj/N2/BpegNLDWxS/EAmQ
Pg9/CIKV21SJMjor3hDgxAIsLwNU84hvhxPHKdU9nPy6wYDHs3GeUCPVaC+X42oR
KXnAUJkJ632MOqlguSMvzdNVRZVO530FajAfKtxFYROnex3TlkSNPCPXv/k6Axiy
Yo5gLHTOtvEgrx9oiM0rfExoti+Zl6rnPxV35gi/qnwLz7GVAAqKU0CJndIce7fE
0ZB+Urt/IbivXRXvDuN9o8NOBmGabKDcZhUgP79NV/qkDXBV1aief9snauN1z+1g
+WoAXOalfLduIe+3ymmcu36ShabB+m5IyA4HSwmh3uWGTbpMkgmt6FPWGx2elUbJ
+ubvZd/GBJ3Vql+IoNQETJhpi0DcINht23vVUykpwS/2kDVSyTUmQ2dlJKEJT/Ne
o6htaseS4vDPE6h1DCNDFGyNAKztffzCaW0RZz5fmgy+xBH5T711sjnyS+JbfUZF
CBZEU9XkNUbPNACAOojn0JrCgd91QTQdzL/CybamuuOyKepJfAFK5VmPNRlbjJbp
4rBOVS9ffH+6OeGpMSNHf/VUBwX4yiXy09Do5vf19dkavd8kqpOlM3xJ8vxleYVC
IIa7qx2j7CMk55XwzshCN7BaRqN9hhEN7drheS9W/RqqU2guOsq9B4eUKRcEdIY1
URd26ozpw2iWmImYR5r4PHjiNhuearXPx394IzjKLaBvpl0IPL+460T0rha6s1BX
n41BxSbqkSgFuFBvmgoM5xfZPYo6TId1bssC4Zukfm2gJSDSO5PP8IjOn0BC/j88
hqWM5Flh1ACIRCkhPLtWyunVwKdN//zX/LC/WrDdhjsaAtQJfMykHitHn1/W+a1i
ROeOEb7J/AQU+n9dfbq7VaI7W2xlnYyRqAkvy6PPXvtJB0vIYWUFGL8bv2u/Knpu
70HtEIbAi2sn9IT5s6RxGLg/D+kXQa5kibaP23wUiMcpz4Tpa4WRUDXC1t6pF9x+
QFDOyeo10EuwKZC6leG7sELL/zjNTf1S87t3QKrTKh0P1aVzWM1Pw1+rJHTKaetw
m54dRdfTePB7Tt8GsOp0ieR2FkOKQlmCtARUqnL9FSzH9456Qvig27MwWtMQ93sV
JE+/v7kVkxt8LxJxLMvdfA9XUEwGeTG3bvpJlhYC9GtYil2LGyqA/BPN9cRccNsT
gi1n0l2dODcCVnLszdSPy3lWd0o9+OmG6uiCoh5K8F5K3ca8NTPS6atU/LI3T+oE
mXfCkwvK7xWa5sOEuqL7LfHTJPOfc+UmxAZH1S9+YeBC6Z4aa35bItgdO1Yzux5Q
QGtV07dQSUM6BhyUYhdip7Z2zo23dpORZI3nkNCgw6cVyeAKMZ293CINH2/CKBZv
iPTecSSH2PQKbhLoyasZ9zL0Bkd3pYKIcr0lu7VmBakOkB0NHhbU5wWOkBcNjHbd
yNKuYAgEFYKzg/PWHdHRB65/1IQVMUSkorgSxik834TTSuV57Dx9ZdQ0UlAFAOGz
2m2Pp7TRGdwBIDaq4Rl8cCYFjMHCGeoHHI7+DqWgw8VHYq31M0OjeTCiRM1cpfwy
6uP/vbDYdTFoy9CU23+COnNdy9BkLEMjZiVSOCnx1NoOxU+ph+6W8yH6rHEK1I28
XGBNWYJFIhw4dGqleouKB/Pkrj8FJ+5JpnpavCy5B8nKAR8hLLSUPZ9XPEmm0tuJ
hXwDcc09hU+tSzGEMmkHJNgC8Ucxc4iF6E8I+h5I2JXOjzN1w7yfb2Zlm5SU8YUg
69V/fCcRqY0aLTNW3uS19zJxRscB/8dFg8QLCHXyJOzDDB8nDlNTDv+3kMoNRbDO
XC4+mODc5DHYsZb15vEm7Lfwzz6D1/uk+273b+lC0cg/LzdG0G5lnb/AZImIv+0a
+gsczLEB2+AGB0xcApZvON3E7ba7eGYnwqH6zO7ooM4G6VFjf69Xz6m4Sx2RSzvT
yNUkqhugpuV62Dp8tBOzdMgK/BLWxW0VsgB5XMLBgf38tsz/LBtd06WzZ0kN69Fz
97NotEIRZoGYch9ZQxfge0EEppb6IPoK412S2rA2Zv6G7NBoyovHK+5GFMsR+JEW
ss3RwGPv4uzQU4cKZJ58UI1GsGHUVk3LUdZxJ4V2oWokgGS8Ya9WsEsYTRuEKwft
EAGvG1kjLkE431BObOrFogGcce9p4qY1FZLLM4vLc8wFn6XYCdQrGC9tnOkXfM5u
R6FDlU1pGXhbpM8GUojnlxVuXqf0wrnODilFqR3lBsMCrtwXy2zI6CTI8BeBVR3u
cSkrmVTXd1el/Hx28J7Ji28fXYqQ+1Ni552IprO09VuebEqNjEIQsbMTAIXXcWTJ
iY7NSpUrQtBxCLpT24dNz2UyUwfUViL14l++MLev67MJoY4PTiPk/yu5uWpQ50kC
eyDXZ6cbFumq092rxU+h/U+ZsKiH281FHhfQDa8BfmnRPp/YOdI23q5te7N7Vh9o
g23CSdm07E08VPAuRp8Fam26NzmFfAh7q4LVL1j+QYaS7FxhYMZiAeJ5jXHAk0jF
wumdlfPGPSLMkh1RkP/DemQI0l0SR6hTDRxqdX+8V7IaEHlo4SJ/FZFZ28iyhD8c
wmwCEZnL6JV6S4xw/VF+pzHKziOXvYKyDbO0kFP3sX2VYZJePLjEReYIZYMPbTct
LMM6zdyZQmKD3Hk669FrfD+5ERBftlKcesRcfmCNPmPOj+JqrKGyqX++RxFvIBp+
6NJiFgY8x7Hr2AGSCiT+M18b3ZV0XYwEUkcdhGv8ITsAPZy2JIrpXF3b8C+Gh9+G
+CtwRNB01VjR1hoLc/GskUMOp5YqLFz9xhcY/L/u1Zpzy3YKTLEWxU8rHeT7jN6t
dg93wksKrSK57etBAx4FnagE/jXNjg8nJzzTHH2wRthDlEwn/FejRxfbWloGVj91
ZF22rq4HO41JgDWF81H4cT3gisbGlmJlREEPKEybTEVuk/Hcn5bfJG9pnRonqVry
rTZHypTTYmD6VTK1KhcXenxb8nPs9E5J+NxDPxJLJsHqq4Jzv7TQ6l8ekr27GqBX
e+tHNzHtPzfdLW3rVuGGnHYiRAZ+iNgsmIREnqLF43E3r5YqQ98wI9sg18+ifToL
UF6WsGXBl/h/C1UiRTB1VG96uUd0WlBaIy4kRnF1//rQX8Cx7YCoxrYIxD0W2qGe
8yyVV3I4nrXoKNcPuHp3B/wBircZEbWBU8hcUDaSzqdZuUuKy6xraUAEVYFJodJ2
UzKP/VSneWs11teS+VH8LHZYvZHM8icELm6ye5C9WSDcLatR0yDs1GDq/lEO/z8M
wWBU0HDk+OXP7a55bzBndCQP7ObvUUN7Afcw6mZPZIowKuD/pBIPaCyaxQyhdctl
9AymDCtsRRdigunC5k8oNB+ZJ7jmy27QpUoQuTtTz0H8xWImSMEVqSUlOl4LjzZO
+kT6YBnbYMZWoQi5AZfpzpXt3jDVx8EkroW3FyqesHDDBmymhKFcHtw34n+ia+aU
VxIxpEyIUCJlmA06D3BzMOw2kv8PDxc4hr13l1rPEfJ18RHo3mphZtLpSjcNiWVq
bMQz6K/Bx50DnOp2fRD2CzBogK+QlY94O8bmsgpqyiqRwnLuplVJJGLHjvCZPcxL
SVc4mYYV9rbgHCDYRCbMYctad5TVImD6yVFj8Ws1bI3BT1odWlbmElUlC/7gFbGN
22ah+0VKCi1x9XA0exZm/f0lMyniIbNpzVfa0HX22t+aNMoiIVxk5DSHm7viMXvl
WaKbMw/3qjLbMm/sT+mFqe5kgm6JYdMaNcGyNm9Cw1TyqI/7seP6/l+lIQ7uIg3i
HdYgc+C3tFS+Iclkh19BrfryX9drwH7CNORPOAQsONXg8sZvUSZtZwqpmFOgNdkZ
Ci0OrBRDS+4VujYyccrqBTy549GhAml6K+5ENyHFW3EH43+8IieFFIejMlpXEexS
nuwiaWWUJ2/rELwkZBzg/3jXHjjcUG3euueeSd0Ob4G4s+CLMMiFQIA38ocbQbVR
tm+fdnmS1e6vpooew9/RfzJx5lurEwfh1uNoREDR3EjfDTotRzOwJyjxRDybA4bC
kMm1v6BnrFVO4BpniN5+rSDAtuKlKIJ6/vm3MGggCkVyKgy+IkpPxaMiC62mTU8E
rMUTQ3ti2zfKaK6s245L2dt2li+a3ZB1CRbCxga8XP6AF+tMHRqQwcoN7a1lOE8w
Pn6xSHnKbJ454abhtAYe2mQ3DvToTgFBZ6zO5DzlK6PY5lQznWsh0Wb8DPnXXZl3
23FcpItLqlQf0yTpRk4B0Cn1ey6G3lKu9QeV6R4rXxcubeEP56tzCf6yMU0UX/Sq
planRPURq5YbDKv0wqb/hiZToCm35v2Nw2QTRthTzgu4fgoOflZIBYMv4mwpGvr9
5OU1pjP1lq75KhpvPkkPWY8utZ6zL47eGxpsE3PBTQM4i2DUB36nJRwlmnhWQ2c0
IQ8oCIT7Vu1E8z5Y2vG7MyPcpW8HrAYZnHBHhcEAbP8d2TqllJraZHNANtGYDIud
V/8Yp4XaI0CsonlK4bOJeLlxz6l8lvyfmGGvfdf0ph9x/7vQbUezm6l5egwJzIsR
qakQVJzPsgT9X2zTzvRrRXRvFLQiXkpICZVaMTv090Bp3ahwD6o0yHh2LqqsmvZK
M0weSZIF4WTofsQneDrge1XdA5UAtchHcDGf8Ve7v88EorxeZpemFOXtGZ4MQrUM
hF0NJWP0Gq6eEnOsAuwp/KoLQ3nMybCFm7n+VPN+tdOtBbPXNYxurHpkfiFlEIpy
nAiqLlJ6PVdo0KKRjQLNLffh4xRPzOj3HZFER1gUDZdM5RaZhh7D3nrUHfIEPPz/
oZnh0BAE0mgVj84tikvum0NN5DjL82MyQLwckChvfkLCARBjN1VEdVxfQ0xKfKIp
dxGiOAesLF1qScRZQqNvfsaGqRd1gbbvFzFTWImooE65/SyhAoXwB4rDlgjVC+8+
eU9ebxOB6yje3+SgLJqvqA19UEBjRK8q85omNlESzOrcV7rdSjK/oiVdN9FaS5Kl
HPRAGlBlG2i0bDZPfAJHw997tv6hEa1iSW1j27HJQbTa2wG7xgpe7NwmVKzGFIoM
/0+PK8JTunYjEet26aHP+ly6ZCXndlqXwGx9cCbrY77oQcds3bIDyTU/zDcpLYrS
ObH0rkISrowUF5PSGWOfJ+/c/0gwZXuEfTelCrG3L6CiDQqT5+ujMIJsDrnOkytR
9+Ei1UpCran0UfH/jqs7PjJLadDqYbSehG1Su57kjXGTYmd2AueIQzcccfRruYa6
AIiQD49DzW0YC+eszgvaLkYcroJ7ic2E6r6PRrc+mqH4X28Jw+ZZ+P+AEl7IsNMh
fcI2z+4Jtlz+6K2/YjrcbTpiRdr9ActmvOrlnpUFqTESXUBifPYfSwWw9AX8jSbQ
zoEgdCVnZX+sYmqJ6pIqlAWnONLLwno4Swlnllw2EUJZMD0CyvF1IFgQkbqg2Lv+
sZOWxzRN8IDAmafRUQa8jZ26rUlzHKnsiQgoAMPjJPButwoYT0ClKq9Sv/lzTLpj
XF6UZKovJKyqIAXlhpYi0oMZ8pQPhkYaZ8lga82d3+pJWADCrA1TxlMaunwSqPEo
jb4xkA5LSsmfDZ+grdVuUy5lTAV7CPdOCi9czsjGvKv4VdoqYk+L9v2uqQ9T9ui2
YxM1FgmoP1PnurLTvdDxJD6iMmVpfWsN3Np1o8U+qJawqELJqYmgsqXkm6R4K1lj
cBkrMfp7FH4j2Ch7rJQDLE0Dp7R/zalAGqPW5GtdFiBSmx1Z8w3fc5vbT//dgwMI
fFNWoUIxnZPzQn0xi5xgleh/SnTHr9jdqKOBoM6pKCNDw007uAnKIdHOZiEvuCYg
B3rLEYq37PJenC3NpOlKMQx5FZ+RI+Y7BELZixvV65oyShjjW3jtfnh7oSXhMk9L
RpmtNFWAGZAdiq1Vip8cTmsXx8Imo5ez0ftjIk2+3ASIR1EgxQzCV90c6wuMP/MX
x3jArOVpde4U8Y/cNJw3LqrUZUBO2ezZsPrUynjw9bzcjexPq3ii0nNpQXE49dJx
VO3shnmG5XyzdDMHOAxyXNPZG1X2ptDrZxI8PXBL4YTkbCvdivD6Vra6UI0DhhQR
EYlTxI/vcbe+MLiK5fI6QgBwcyZ0bMUWWhcrm5z+Nm3sKEma22kgjRQYQ0ueTu3D
EawE3iTljSdmycjZjxId1gdexVBO5LFSpGpxpz++KOJWLsUHqYUSUXiJO4eVWIvR
30wVnJtUTUkJVuz7wWt5w8Q8qJ7IqI7XwELJSQeetz5KyprIZ+rRv1OA8fV3ONhq
xR40y34ZOe7Yf4jsSRVBXZzlW88jSpBL5NFZieS7fYzFMi1FXpe4CzgFJWb0t/f4
sgSK0Oka2SgcMjZtTpzi+ZTjptjIa4ny5SlMFlCrdtNmaoxUYMAHnwWgfo2UROdx
cO9o5nEnZyqVfv8ozNs11ANjWHg9WFM4OvqBaoD7/6RkcJinLl1Q0YxO7NNHh14I
5NMR8ORb7Wcu78PDZDJwBglvnrwuAyQMf68mhV7We5xjU9HI0PdPM1qP4aF5FuZb
CpZK7B1hZD3VwvQomPTUC5WdAE2c0ezIqWEHpTtvWkx5RBdu0x5s+Ux7dX+5Kw5T
Vtmj+98dzKIv/VXS6HKHAxxiDSCPbaeoY05AXKbpU3HF+uJjWF5VEMq6GsqYIaYu
y/PIXOyiWGeal5i94Xi8l5B/lqGGIjOynja2CZ1dxj7xRgqUqft9IJqveZIK7sH6
YwO5oGTGkA7S7ubWds5W7PMSkx/U/wGeU26s8AvbC3XQyx9QkOrbZUvchD1FHobY
tZnZ5LYfNeVm+4pUO80kTaAXhwNnNiInMALcF3VEbiJqJIdKB+EH828KRucSVife
7p+5RXOUUAE2ivJBtwvrgBOnLhIN/it4VX8b5USlwf1BnpiYyVAMMH0ZyCE6hBAw
wnJCogUk8uJ0wrHwZpUHHghuda5AZqe39nrhZMAzHZFkmpVYzl969UnWajiCwZwz
XSrup+eA76T3E0GswOXnnFr0dyCWaFWnfgcA4TPZPZwnuJcaudEP3NUZVCgehsoH
yTEm1CIE/o9Nh3bKa2subPy1ZTQNX0UcwtXy2YFEootvtvxBc/DuTAT4SpYVrrBG
J93xTYzLYorUTq1sAV5VuCNAED8cSFtPYqs/AvqOdp9y+klJzfIW+GhrN7BqVJ1v
T6jcQlNNWA5sm2PQnEX3IDUYXrivvptEibscaeCCWexug425BU7qncX1o/NknmYd
/nQo8HjAFYbElpUaTHMGSBY4EC2U59XzjM6QofzfNGA0a+RJfqqHpDxpBtpaFf2T
TvS7RVwvbsbQaPKQuQe8nD9TzocyFtntLTttWqz/FoDI1cxI3Bu7sjuTSv4zawRl
H6tOZ3iAhE+FsblNVZfyb9S814siYh7rvZLgc0DnjyoK180RUtUKGvQ0sIIyM+n9
eb9yWtXIEWv96dmuVa/HGHVcCv266lW5wcZUfeyHxoS7bwi2l0+6ouFPaVfhn4Zw
gIprmT/7CXEma36jb7tDcjXHYNQEm+/Rv988/TalEEvcltd6+gg3svd627f3hTjD
yw0Whqxzgr5zcqvdEPYLdAatoeEfcXIt3RLR/XSXHN+sX+1TXMWHJxjsPx7F4tA6
F2WGdQuLCp9mEkP9SMeK0lhNy7bFYzzwoOYQwTzDfjXEDhJutGwvMW4dZ+kdLD9m
yd9U4vdRQQKE/sjVrPVyfXuPy/wuVXALFgvJ69U1CRSO1Y0n8+JUoH1iFVW5IOEo
XPsFldKt8gXUJlcDMY9dwbP/dTgBhMA8h3nG8AbbrTaDppmKuBlmEbm2l4jzxIdj
DGvc41Eyn1RuQMmaqPgsoFarmmLuh3K2yysZqv9jRYmuPE2qKjVZXSAlFv9f1sn9
fqLHx2jYkCbCp0mWvr9BZxGPgeQ18BtaNAi9yYY71Q2r6CX7pmSz1UEYOnE4/Ap7
hRxnYoSvySNwQX8hyWIF5w94zLJZjxTGPvyAyMuGpLAYo4fnZwdw5HNYccsu3YZE
KM/oOgsh9VDLIgr+DMUL08jxmWQErxpVV7ldkTEPyViJb9JTznxC/HnxQ10xW6ey
3jZ8HKyjqeoEgJ39miw2kzYbOfA5cXSnfGDRf3g9HMdlWaJ9AZWKsbeumzH7DP+Z
AQykhOHvpe2v7Ux0VY5Ed/H9+Wlhxq8frSivKC6+MOzvMYW6zrax9+9HZSbx/aYt
dDP1cUsQ1PD81S9CKahTB2+BwqADtoWTVDcbIpykr7jyOReb0HihRtm5Nsp6FO68
xMSVi7IsvW3uvufvnP/knvp5Wc9ezLTPZvwNO8UC80C/CNsQMSHyP73kaOX+pXcD
B4NdMSuVbY8HC0nXRUrRM2qcsq1jHslpAEirHuaBqxankjRy5IJG2YuVhB+oPXG1
n+0L+h1VbpIo9gqC1Ofil1yNtQtMPRRWyHty1iizjsUvOdCI5B+W7ckeloNwksbV
UJRfP5zd4LvJYg4WOQSvnMWwZlTDqN3N7scgDGPYf8WCAHDV1OTghX3jCE24ZQdt
NNo+oBE/W4c6pXfFhBQAy9WiXYMeYk456iEb2zkmRrE3Z7csyReK9f5Utnig/eUp
EzKA8b4zZJl6tVIHuNvgDRDoQwyg9MgDxpAL52CHKlgPsdWUKo65nA0pmNacV6jD
QIIidBprT2kSm9QsB4N9d1LC2/HbfdwB2G4xldYCKC8m4NO/D4/OSk2o8jrEp2LJ
ARA0VfDyb4x0Hyoj1X80YXZC0LDiMjCwDB1sTxYp8T+Bj4SCcpZB/C7zYYbk1A4O
myd2M+oiSUl/B4MwfiyswJzOyAR+i7u1MuOKWQTxctbZbvaKV5iQMcxIWrcPsMkD
bdkl64rlWlD1uhqDtuJ7fXX4wd2CeYdf4MApM5CSUbtwYCyT6OcPAcxtl40nOVHD
xNF/lNTJ0orKDP+Zsv13utYdl2srrFOjg+a+o5mGVEHtFC9Ucfa8t0DBoIOSKBvy
NPdro0HwnY5z40hMa/Fm8svwpvGCfCpn7ye33lhIob/g3zs337Ywu1/NrC7HTq8s
tF6HNKP4J4G8KLr8znfxTbeg07G1lrM42jCkDASwMPrHH0uDwmW59UhjwuPVq3TU
h8ZQi1wa383Bo6oaFEsewruq8EwNPF+JCYmIZzcK65lO+3pF9lcaR77PY/+8obe3
LEgB/vv8Rq3khuCdH/VV/fjEssc9ikIDCMkBGA6+yx9U5Rpt7kUYoUR6YbADoyeP
lbJMnzvIkzU/fCk9nk3AycX9M534An+nsNYwJ6qS/rnO6fhkZN1Jo6pJoONa/hpy
1yNyHQDd/drrSxiEINig+gNUrV9hdhOkO0CO3Wloi2SEwlnQ4GJ9XA8gk+yNo5tx
XPTnxLdreRiF65MYuD4oNWaS4nnKPpuwe3ivn3PgUnwJTl7LeZATmEZ/iE2pmaZY
ucoVQ647tgTyYRFK1IysyuPTm/CRxQZKJwFLjYWqbowfTDafkFibuIesGgOaalww
/J3hzBAZfpN7xG7X2OGvcU8+edo/mUjNg9sDg4MGA6k94u0LFW6V5InzbBIOZLm5
bmdoUigHVfH2C0pz4jeAikaq5bvd7Z+vVMNiR3U4cHh76nPlqWtQW/lc9TFmA5c0
EyGCR13ATOynB96hvrBNaXpy/T9ReSsPs43QhBte28eDupo+gOXz/HN3FGayC3zF
ht7uShweXs1r2oemiSYn2M8SvehtLoNhEvlJpZySYVweG7SKJQiR7wU/XO14Eikq
25+SadjhETIpQvHk8tMgJPoDSSTCRTs886QLjXyEDQZQ6AH7w3hO+WBn5ll1WVN/
PuoxWjarcT/tS2qNj+iHFjs57UZGjz/2Pet9ddpXGUoDZkiSiISwlpnPesWUxHYD
82ncP1+zIotgx07FZXW2av3/Jd5ymR7MfIMn9h6jkqr6DKwT6+mOb4p0FZqrChyr
PeljPSFkA0CbzQg1qh2l1DPm8LDHQsyUTRx7WOMKA6vjBeoN7MQN10+sgE3krdDj
t1jf7VSHWqteNbsZs57DxSrYsTLYlwxWAVMptwcbKEJUwBKKtlCMpojVC7IlZUqC
/hQSsdC6cXpWKM632Gjj7XLioCj5Y7MJ9Tr/H2Dg2rAxnJMwME7FuXSt7fWMENl6
4yP605X0g+e3iiRhVVR3ERtPzGFB9E4AFSusy96RnYdrRfAaqdUE7LGy1wedLwfq
SyszHQBhxjfDMmpLWYetduoSH2zhrs/xDTzLJbzWaww9EVaT7eeUXlzgvktrtUh5
SzO5bTnETVrZH80Elzz1bkw2QxYdyr9YP+Cf8pgjwz+2VRyIUR/8E1wYoAnNqtNM
adEOZmQsqcJXi2T39VnSk4J+WK0ChRdcJs6GeAr9v3257X3QRwf9jk6E4DiIJ4jm
GSAi1rzW7Xsu4jljUx5sfzSAOuPiEDKRjrmUImz8W29D+mvD59nYvjtYEMD64AI5
RGH1L1NXYzLXU7s5h2kA4Gn2fJIXUXJpvy4l9xoDYPt8dhnOBulmhpSdKpmE2JsM
SebNZHQhqSpv0FsMOsQb8oo1/NMySo/70j6qAv8m01fi/Q0pFb2wnT1jT8sNb107
vE26fCfc1z8lH0+FRPtJOe40NIThvDSXR3JyZ46XTT1yDMgMM+4LFzhdayPL+pKv
RTf0/3bA7fE4oUmNjb1PsHURnDOPOsdbmtzfuNF5Ns52GmTSc2ppALyNszbXUdKW
g8O0ngAfyEhhaADPfR/O1zAd/qKsWBrdja01LFsnAOOB2tsNdaqkEFnxpl+y6EB2
PpqO81m1eYBs8bTPYV1IGmPTskqTm7NzPo+eam0hwGeWYn3ZANPfpAGxe9TQJQmB
bXK9Kw20oEyH5/unjTkPYUVbSyX78VQ+bNIiOgkp4jEgo/SvnW7S9ekdSaGVbx3U
TDJGwJhVUcK9DFocy/GCkF1YwgmuRERQQ37L+cplznB5FYpCY8OBsmJ/v6qyHed+
3OEP/p7WxFIeRuVbxwXPiOliKZBcz0RU5ueiTlApqeGUedf34WN0ySYOb1TfxIwz
P5lbMg1x+oq87DTpClzsZN5ALTktOPgJxdg8VrUvzXpFSBaS8uI6139TqnAV3Siq
g0hIh0dbCSJWUR5KHeQGwqrdr+ed2gIWEBJDYon+uiAOXR92YwqkzyKujttPcT1X
lmNW5DDet4Oplcx9d7rfFQ+E2yEsKsZ6BWVolTZPUVEPjEmLpaRhHhfGVW6rKnSD
vah60BHqXt7yrwUCGn+infLY0JeJThCSPwxaOVS/qVRdLERB6N6/uN+jw8IaPnRJ
P3moXloalTLODWtwFX4Yhw+c07c8eCIYJOxn4daV6UHAPgAiITpOaWY3PUo4uUMk
ZGP89vG3uu/d5oQeStqoJH61QS0E4BRWhmZzPnXrzKi5iwAH71rr4dx7YGq6Ltio
O/6dlgk9C0+kvWx1Wico+6KdS/kW1zBy/KcLdd2r0tUCFGG4GCq9wWOMuwzDua4D
fL0tC/eBwlJz1nEs4TQkG4lUZtmr2gT11zmBj0QOL/at09Lw0ki79phrxuCJWbAf
MBgmDPwGbn3m2V0Ha8zp+7fcJfNZetYk+AfPCHvqG2C5Md9ziAwNYvqa5TtRi1cI
Lq/f89V0uTOiQaFtm6cnspWFsJx2slGdXPUdZ6S6CVfxT1NRa2JOvNbpEURmaG3S
BMs8RJlC9jnwBYomXqtcnoIQRTircRNoPl1nphcycI7gOx6RCe9zZiwgoyxpRoB8
ceWBwVrmht9vPZF948p8OFw0K5pX9URXuEkq9TFfpwEjMJL91+O6Ig2Mj+b49LtT
q2oVwsdXfB6KcH6FgdSm0XHIdZblDBN/fYz/DuPriQo5jXmirKjdV9aqfqYyY8IQ
uFEE+GL6r6Gh5dzNDItXofss5+ryNNy9JvtZpyQDQTsf5XRaalzGU/SDFfBGEhXN
Kzpl1XcxMwV7inWkfBYB1+W5K60O63YyK1hNrC2ouDqxSZRj5UD/XvfDny7+3Zpm
NszVmSe+/eEaI/K/EKhFBSMLCdGkYhbjLmLH405h0U3HdrrxUhvzdpdZ7Pl2Aq/5
3V/r9U7e02uwOvqPWn9hUnVcxuVH+ZK4t5j5AO1DavFbKsdGkVaxLYHTzEdVWfEA
yc9ZlOW/m0AonakDmFdzXg/MXnxeAkePvezmnRw8wX23KVEnSk1aelLofSS0OE14
gAOJClMlyvksbf2zgShyRS1jWOR2/F4A+Hasaish9R+7DBzFvrZvI3msB3W6C+oG
Chn6f1khFQfD4E+GHn96JPYM09RLAfpp+3XbDGGuio+VEQOVqAjMyLWpseFw6dIQ
N2QDnnNDy067mr0nrlS7Ziaz5KF87iQcntxXUciEZCHfG56NfrexPpwsYjJQHIYm
lX/WHpCTIX+YdWvRCMASzc7M0PQzDNPlNzzmDqzHiByF2ltiIFhLXEuFbXpZWwkt
F+GzkD8icypDcAlc4/LIFC1hd0jTxx4Kz1HXEBxZoBUCLeC3dtAb0rTfNO56ZVkW
iet7L3ebEO6ydQlVqTMkixSlUl+wJsbVvvCtC67ZZ1JcMmUw7etO/V2T1OaZ1ARH
CiYA2a36GXMXJbumGXEjHiM63Q8c+IPX9+D2mIcv3r0gmX1hhd9Nmfp82USVvA7z
RbmWXmRD5BiWYsLP2mbrysg/7gdpyfHzIu2jKImiwfNnJHYm+cm7Jp8NH8qzryCj
9F1xIKg8GA25iMXhDRI2CSfQql5zH0ABNEv0fW7DNDY6NUbE9u2clXVddF9LnMS6
ACP9IYzAqtX9br92ioDoYuwSYKJ3Kii8oeV4rvPqosV4dbsZppXoZxfmdkUr3MKx
COhXmFq+p7ft3NTAK2HnK47cMBD+3Pob/XNfjQm2eIRtY8TXAqfvKTqh1lmxguJ1
4D6NHMGM4XMI59WdJgXm7hIfBsJpRjiihwGe2X3pHH8K8vtqNTYdvifN+DR/7VKp
Ts7M8w918p0EGGOb7BOUWdRvNekDr1xQGU1u4vqUyvytVdA//2brpASmusQCvNNJ
3P3VQpvbYMRIBbMnO52VGWxesnegp1aY6RE0SnxcmAJm1zicyk3pfL+jJ8Win3AH
9cfr5rdOYDWBFLYdA/P0Q8MMsVDe2TjXp7WQJti5CaZ+no+aColRy81hkr8EPPEj
zsonsMbW9LkolPFn8t0naAxIq/yRIcGzsOI/i42PGPk+nkN+L8RYjXK9jbVr2eoC
dAcvu2m1efFcBW8m3gtS97+kh/OmW2Vm4WP28ofrBsXN3CfNAN0jjcKtAOgjbk0S
pria9CoPjHhp/YhjOaC0ToOHBNQF6Sz48/ppcLRO9g31Fk/OZ1GaSAeUffJ7hiw5
OEK0Bwvc+1qdWdfoQWeYYLArZL2JMT+6hFUMt6Psopz4gXgW6zA84ANcQ8K6uVGj
5YPeGIDnwlxSBvMxdgwIqxWYYTCtD8ThfT0SGGgYS/ox4tHi8AFip0CulmAZAfqm
Gh65GIRgRLm5Bk6G86uEEiJIKi8W5sYcGraNSdOPC6/3KoEG0EzZjU2JTTtY6LQh
9leM8+hUbbNHmXnkNNdaKwmWKZe/l5F7voOXs27YbU+xG6y2CWKVny+fg6nD9YF9
BrRqZp45vGV0YkllF+iPQin4b//VF4UYScwc7LV+Q7TQbXFKBvSery6GlbEAdpxO
YNXP6jtdTn7r9kHu8R5dYHwmxln5O6aquAT/g1QCCdCXkLoUc4EDVb2m8XKd2t1R
qO41xbDSWR6ExxsZ4g/ZBDSF7TP5ly+sQN1XBB4kTQ4jPTE2i1LdkG5ONoP2/uKq
rjj9sxQKYGYPPdHFklHaTD6WxmSzitJLLbnJl64YaRlZnP7LN3ja54kgcktSXStj
W9fuI6Yf7GV1gUXkA/n/kx59mVEqbFUSZrHivkXljv04EyEFbNFebwODxQrzK6DA
hRJU/iiibrEjj1BC6e0EeW0nVEvpg9ea1ur5F3ZwLDPHDtS+rDk3roybckdYQVfe
zsxVa1RGDlPPtepAOlvC1n2Am7U5MmYbYLD4AYDQWetTthT8Yi4xQiBUuHCSvxP8
jQF6D3t3Ys1t0YYCj0LZVwFunczh60p8Q+cgatcE2nOkMJqPODWGMxTuN9fVCWqQ
jIgHLfrlescOnoYrEFg1wMhAy+AD8BfDQ3gEqpCZXyMjVjexytP1d9v0CqB8wHW8
KzJmsyjfAQn/0j1V/SrGLhWdxRZX8LE2xy6BwqGTUK+OjDui1OrDRHEeNP+rzxbg
3wjsYD3eTSXyYooyd4e8i+3MvamQz/0Af5Tm95X5v3uez+ULxf7AWFldADpItDEr
pn6yeHqyBtDVJUHVI1h47NHHu7bfzCD5hcYW/Emu7OZoIQyfkv4aWOs4xcY6swqe
x+MeBjE6Q88qY/To/F0GdW8YnoSFf5PuqJrmIgKL0YROKmzW3dJSb7h0LQPexEzX
hnDwDucPbTe9YvQhMn5NG0tI6u4RQcE2TFE2fuMCKTu1maGFXjKP4laWbjQUcNaF
kSR90hatYMSsMTjDc8/8edzTDiMNVH8BbjSo/uGQGqGQ2Yrl0nwrQdvLOo7FFXjO
+HHD29MfTJhAPpyHdiOwaFXJ4was5Oyli8cBf2pW97lCz6b0Y/0hv5JXa0rIUJ48
grn3MSRKgv8SG5AwYMPykHrZOgZ/1GYXpCX8M/ny9KDPo4KdRyofyb23LWJEmLhd
xeYzSYS394dkqFNBCVQbuY3TPeWh42l0nkupQDYqI2+My9WgP2LJqjF+Hjt/wF1g
oNsoNt4PN+q4VgpNMe8lVGjr3f1oKDR6NaFeUeeP/ddESHG2Dgh88naDcbsDtMfQ
omL1r4Wfp3ZbC+yzJNBrZjtzE4BXcNrCnMAWSGCcpPYcz+nEBPE46cdvUw81GEVL
THLrRwDsAM4bxNckgsxijNxejOzVJeW4dMy7239bPbuHZ9sU2Xm+b4HsI2kn/ncf
pBN81UUG0t+SSQmpCkhWaHJ9s9jQ/kAcLBh+etbDmgcvhjV6hRhFpjAuAAmZh+b6
tP5Kz1/W4mdYarpcI+RHs8cm3hrSexs3Rniwn14Cj6HN8vEaZyXc9UltCn7y9VLV
sqHGnBmQ/+WdbKCyzsIN6jP6u6j7707z9RdLurRb9wUVMBdAsZr9ZSzSEqYoLaQd
lnAY0Z4voH7BpmLqW2+ticsNZPcxmMyo9wpSh6fiAS5GrdxsGxs6J4Bm3wZIowIh
qbDv2zsxsLtBkN7lIyMpH9n3azBDp3G5jQvcVGgfP6/GygDVUavbLPzUdcAWBViO
SNtz80ku08VpWocY4SLvXGNr9MfmI8fdZNQtqYIl7nhqN0NFN3XxOSHZBYCeepNI
2iOtgUPTR1e5tWsAwlx+S9u9R9WmUgqek4xZvnRzS6aRRyng49oqhEE11Ncc50zl
4ihgDj/01ft+JflcPVPuiEmk6WaIvjaAg0C9dNggQ7COu7FmC6Rqiv8FG+NgVqJz
3lElvuBaNp+kWrw4Md/v3fLfVMrFiQDHqTQ7aYKPNPWszDuHR2LPMG/Q0apmBu7Q
c/yrcyeQArI6km3Y0twy2+Yqy0fxYrNdcDuag0/u5b4jbE6DpgAJay2euIGog+VA
JVxP5OJUr0YTurtZk7JRWNaR03PEtinQLd1tmurZ/f5ZJVvKHERMW3Vh8rH/9LUi
P8Hu15AELeGsnGT2zl2rCs/Ca6066ybZKHfVcly7pagNCmXaLk9LW2Cpzf/9yzUu
GQ6h1G+qUS6RNnSV1s2FaewMANF+ys5+XduASSdHQRV0dYGpv+D7c8xQV162ArND
0JlEsptqzBsOpMc6nRJRRyZ3soWue+mJmTEVoHnjOzmFPk9YACc2v4XRQjL7Ywwx
3OJnjbSXf0w4PhlsA6Z5/byAKinuiint1ckcrfulb8+tvX+jzp7BzafDZrq1qKyX
3siHOjpVBf0YgcVkAOxG8alfEcHBsQs0fti+/R9aNwzDUeEnBNPM/La2yYJmDDi9
IgbLjjVIGi/ZvIhcRNVFV4J2tJ6szwQLXkxZREYpP3qY5T8KiKIRg7fI0OVIWr0y
xUhDZ/mturX3G5fdPJqS8J6VAOt9uaBaLVR7JoU0J3ZnjatxnSbFfVmQHO51Voz+
Pj2foS9/gkSfpcMOENpWH4o8oD/7zZHuYwdjQL5qeVzDrs/vRiZlGHMg2XFLlYSW
AqKxA1kePHWoPcQl0MGFANJVtpna5u/6bbmcIJYm+3GrYPClNpLxqwjW+SwrAuwR
7AQQPblN+SHY79gMmWJ0HFn8gOVQ7TmFjtSTRp69ah7YquLEmR57sFFGEfqNo3VA
bAetqHDJBEBU6+cfV0wr4sSOtWVjYA1WastUfpL6YJRRKIAPD5vDegeDthrXcf+x
ctwiJ5Hl9GUZVV6PDyTiWEuX+mUYm+oIcPesL0/nvkLqOcyTgsr0VvbNwyP1taQ1
iVBAsRYAkZOoxprdmwY4emgjGUD1V5OXyGFionwCz5wQeXubozzfap2MEQgpxcNw
bYGNDcbXWLVLt1etxARhv8823FUvJDPeUtDEYLpzGBy++sJKBQXXBNqRznqHoGEr
aMh47kdu/0oEisM6qq9KmcioJlZQgMeTgLfoFYPG/+qeK4YnIaWPc867cW+grNPg
5V8G4+wy5m5LX+q1etOw1GATYW98V4iYj79Oacesbv7j4VMboFVfkuE8NM4VW0Ym
gMpVd3kteUsge4cb4CAx9VLj84GyX5doy5zimKZUobRxiAOyAaXg66siKQTl+Smv
M6vN+mwXoD9/rUB0a+cbBXvm8mA+6D+8iEibTvJe4kq23qOYuucGZm/90r5+vYgL
b8ra328C08UzV3XhmLQsVCkIDqEwdu9NekU8Gt66q3qbJbiZo4xTD3CchDv+QWl/
FJ3x6GsTtYRgLqHnCVWpekK7LG3uYnT1s2DJvm2ZozQNPkFf0iDJUZzbg18WYy2d
Rjpug1RepLObC4GKIu29jLqxhxw5nYNTBtHeTdsDEUb0pTgxdOMoFYgxlbbKdzqE
khQLyIGfMLjUr0hklCSPVdItx4l6oGnB4OASyAhEJsTvAJyaDO1UHNO5s2M5PMuV
4lSGAfGxHsJ0Rf/cUr8Gvm7zb5F/YoWmmau6mMfStxL6JwBcYW1FGrPO5PtBujVa
JwpRJLJtRjau+UVbpuAgLTLKwOzvdK1rjCqHbHSXNi1ZG7Sy6nygAZDzC1axDTOz
/+Bo4fHXLvbRL46sxojKO/zshY41DDE9cqYuD2pQjqNuWarbCkUxx4IRykdCdsRF
CWJ1jgmG+crv4SJsfRHFWtmUN6QbIPm7YBVF+7+GG/Rs9MNGrTygI68/l+w1YMnp
ZJCMs+RAMXQrE2yZRO/8u3osvY7NREpxKATp4bnIhV8Ag+6kN2ohoqk76ZaX+qmm
6U/Nh6SPjRgb6GZ3do+BxdGETGynWAWmoNPuC7yFf3Z7aVtPAXgCLK5kUWJStYUB
XuBkHtarN2czlnJrQckoR+2iuMMLvR3nkgi0CqrH3YPGStVLmMkNkLBrfJdSiZhS
6fXVyYS3e0J+/RW3quP5yWwVUYKhDCq99Up2eR3S+4OTePm2GoVmg0za3vLEGGZL
i8I05TYTB3NVgYwjlW9/AiZOprZjbPfdzs7x1Smiy50vKvpt8SgsqYAMzhSIZKIu
fQp/JbYdHTjXCUm6DEzQP9PU9pNwNeN2KeBjzYnQNR6kDu/WY1C/4X4z+qW71TAg
jC0Bx8w3nwYcA4hwZHqM1nm2uwb8ODkkCCKtfR8TssyeE1U1y5XZDIQweO9NY1o5
+Q98VXn0RgPQEhdDoltmzDMx46mLa1hpYFY2YQgLyohq0f573vnA91cM73DnvfMS
QX/5FtNNY3m/ZDsm6uHj40GSbfE93aoX021LuungV0zOIJR1Msrr35M/pJ82yRXG
kLC5P7M1xrUuQM/vm9ux7PuyPGvmaagBzTBTfhsgumOUZJyK8IbZrYvtZg2ehKJA
+HTCKbYn9sM/6WcTA1n9qHlzxz4skBWNm2ID66bsACxfVbzcYdN7yhsoClMT2Xl+
Bdo6g+VYi2ifTgjcNSg28lRdpU3XR+tURYmCo8Bmk0VJSUoeFp3QrjXUxrpnHHoz
Gt8H+xdWdwpqdPq5QzHOrYb7CNK4pAzM8pFj+aY6eJ9jKr8Crgds+jbcaE255tFz
L146z/sJ8aRMazsa8BWCE0tDpB7hLkbkWqk5lGPXIObMDerggxxF835kKfovWgfB
LymslNzhZSTbdqew6Si8bypWsYUikLrTldTMOWszc0/0tr5ydyxACBiYvQdc6071
NQWG+EVeSkZFOBFwqU28amtIXDTGtQYBn+lqrYP/P7BSuGTk4scOzTUtUEoPNRG+
P9R06ksjZWHl7OoXmaGGZ3Q55I11f5bVcQUOS4Gq5RCMEWW9cZMmsZUrFzofHeSg
C9pXi8kQ3G/7Q5gMnIo9XD+CYWaEJNlzPw9NlYrqU23d7RSbWLqYF4udEYjjgZ77
mDh35cNswIZ2srgVhbUwf3ikSSTbjztwVL/99MZGEEImHHa6sS+T7GctyaUuqIVa
CDoSUmxSac00o3gzNpNajVuVMJcaUw4DA927jH3Rm/KAQmEGdLSH8977cPXFEonW
kPGbKYJa9aDvQdJwj9jAVN6C2HsQ0o5Ydr3aNufqrbNVQ+C848f+khTJpf/K976v
0mVF2b3K4lfjJozqPHQlAME0zXmHP4EnW+nF71VNUt1Fo1UmxMbYzd/xo3Lv1aUz
X13MAkySuIKz8pUpdZiaszTVU0WoCk6mKwP0sivGxrN/t0PFjdugkf/bZqizaWU1
OTy7VH0guvJ7jtl8v1Z29JgUu6ASfgwujdWmXgabjhqWMLjtxBGxaEKB+IQ5tk/4
BGTi6rHa5Aek0pdZVqHjJVp2aarq2xDEGGxrF4wff1MAvSDHB25O3Gw90yXKEFKP
ZDUbBBWy2FUC/Sgpw6tBTrt88L/FLmq5nRBAgzcZNWa+keRT0wd84hlcnrS3Yjm+
PVRqzjqRXbH1vJbQ00la3pWGDyRy65hcZ6FIaajrtU8KC4q9WD8Xh3M4OOu8kdKG
EmIMNjke6frlUdelCxos7Ip/CMXzeiwAVICYyGSkHZ3G6soGhG/lDW+J2cvUHrje
X5PSd/K3YLe0cZlOMHTo4yd+0m6y36mLGIdugoFaPVZRJclOy3QZKZZw80RBFhpx
ajzSAW/nO8mFrTdbYO0LZqZmytcoIYUTytvkIyPVBPtSg9IQIRWOdDbt4NfKYTQq
IyEyVNxiLuvgHx7pzUND2UU0dZoGKhWFVylexee/28HEiy+quDSb7pe4eQb/de7x
rI+ZyrVUU7ApHyy0Jb/gqwTb4Cy3ziuIpj8Zmfer1vkAeEfglZxRRV1i5H90RLvt
/bO1yLtK9pWoZ70dZz3RcuVwStT3j2ZjMNUx0cqVTfYiHtYpOZyW4bSf9k+oneJL
PHfFRlxObtZItzHKe9lGw7NjlVt9JUEE9Nol0J2Y+hAOmn5daPP8bbD4qhShXceT
jaWOwv+T+KnHTBX4oOtfKcrqIekgagUCLn6jIvogogUumrQas8SCZZc96JQAc9Ck
PbgdxJUCm34CHY+OP25ub54JGnWhUcNhvlexfQCvIclLlSdpprDaEzFN3c+0n4h0
/7fqVObV20QLanhNSXnHfWRpY7zKUrklLQyYG4+mfAWT1s8OO5PWP7ldjr3j6CNe
oZkUUcQPf/UaGi1kJvXQJgYaNuxCbAvGusU4C8BlzSRRGR/wGYPwgeeLrGqVqsEI
RHePJWQUIa2suDwe8ma6OhxaE3HCIdtpAHMFmYkQxMS8ZKLLLgcNIS0O1kCUmcu5
B0mtNtHDh4x0TJUQJbPTbUi6ifYrmeJlf5zE7dv3he1uz+FpdFXqGT+54FG3L8zV
FPGu5Nn0Dgn3RZD73flciSWhyIBO1Wv8TUAxlnQP2zDRTObn4jM5lEyigRoT9yFw
rSqvzh9JuKyE7WRJVLyjQab8Q1qUw4wUjj8FEBlpaKotYyx+kVtY3yTjSVhZgDhH
r6co5cEcypSB69zxkusiAvObgsj0zK1AnQhrAkzmFKkfiGePeaDuKYN+Tewq5zxK
IK1xh+mqglbAtjJ8EEcJmJwKB8BFpk4b4QPaoQTcRKVwQEV/AjBcH6AudQHxozAi
hyklcFUDVrwjhiCAknWfuwwGwcvMKDf7kMKdWpjba/msN4uKQ6/aNW7OQVY0pjFi
TyY8Z2Nko1hl9Cap7XuiDsRnSvgqLRx/BeuZ9/EVIeRh/7jbv3sqNzYYQAlZMFp0
HxZsRSDf6gGXsBTlzYPGGJW0bFJtclkHrpL4g6SAAK0Ds7azmewHC33USE3g7umi
+dY8aj1Zi2fOnHo4BKlUluqyOx0jiSuKprf8SAQND82ou1oRxBUcej/hpNapal3M
bh6pc0d9IADYrggzyE2f5PqxH47J0+MwelY83K5BZmuz/B7h7/RYQJpOwqxTXokU
3sQcrV47qTuyYs0jDENZO1fT/o7bTFjgZxjPZi9y9N8tBZ8XxttQIEiy3zSmWO58
HuTEC47ELunl+2DINsF3xmIvQsHr8l2tawVS2f42rYk2QoRYyoaaBp+JKXqgcUES
iDcsY8Z3jNLFBniEAB4VBypx3gcSxtF11tX8HXM9PNOMTEV8jX+V6gxAVPSm5vV9
NBaodhzJXXSErDp3W1G9LhiaC+rLvYF90f8o2SAcSbWlhwjFZd+3pCbj8WywQIOK
rCBAS3T9MHKukWFXVV0fmqhJXc2i3MDRia5LSfDxaJHlE0PQT6ct/unMnCAesu7U
p1g5a7iRddkY+CqCUJcqPtOmIbJAZ0h1LSbYZ5hRkUx2j8j0NhPKSo9eZt+NnzJd
hjKKPPBSzB4ShyR3Uj5zyos+DXodmN9iTk6Sbirc28EZtcfVzriAzpwdoB0iUvak
zRKFfwpYoGAfUuM1qcP8+HOTxF3rcbfeYImRHL0ITKKXN6KdyH+GwuDsyl7GWT+5
yRHHnu2N7gWDjBmnrjT25pUxFi5gsNhj6UBoFgREixNm+UFPLkCNEE7WpUvDHFAF
V+15P8PPATp43qttSZdG0Uq4fA30eMAw3dRBL8srI8409Cat3YAbHUidT038zZmQ
NZf1LzFPsRhWNrlxdMvZN2qfp4i0GOpG+fjTMli9TogFf+04aCQn2q9OWutiIw/G
tZSk43FBWw6WiZ1gb3IZR/6/rleK0LkBPnMxQc+pdNtppzv7PvGsK4+b2DHhveyR
JfzLJMu+Lm7ACrKUTvUReYQwCtGY0pmnyBe+Nzu9hr0SgcUi6bsuj2LE4irLl1Il
BeeX8YMNMPC9RnPFGVSfXmKibBGxdbmp0/77SKPRfbQnGajRXmyuTYOTM/1bSlMm
xb69qg/kYuh5M38z0wtPVJeUsEb8Uri4hRSnmtIvIR1FF4IEWgFg6angkEDG+zjk
s8WubgcVdkPjldx9S/AyxLQyF10R8FQNIGnrrf42HMyzFD9+BQvrdaDWr7dV+V1+
rFryCQ248iBq/ki6tVLebMOSllm3RDq2od9OixorByMj2WkexlKzvm7HXrI77/3c
7lEZaiMF67ZUtmJGZdTAv1r2hslguPH6nbFxtZa6qQzN40G/cPSVtrvjHKUifx51
+XpzG4F9lMd/qVljhhdpYLqUOvLinS+vqRhVGIzLfE1tuIUFAE2Gxj7GBIv9OHKw
U1Hn/V+NQhBuXWRPfpZs+NAyju8gPUDx899Kl2Qni8fjT8tB91H0MamG9FnQ+wSu
/mfxOOOB0lQ9XxAk7Nbjau50PVOsBOtwdc2IkXrOV+FpDi/R8uhcCJPTvrXFnRnY
MiZcqEwz9JmSnkHXib9wwEDdhD+xKAIBLIz/Uy6LPImLWmt0lG+OXuET1gvmCWxZ
iBxCdoWWJbN1o8PhwSs/scKNfalnk1QBnT5QVDDQBVWq/oVX+fZ82RgFvMVvG9W+
WQz3J0W1fzPwXtxCBSapx9ltxbPlVTrIVK2lb6vqImt9rYlbyUTy6v9Yfz52axfI
HltVQ+WP9VUicXRCaIsAcS/eEs3b9sAaTP8W+h3doEZkdGL8JI0rwORKZ1y7Xf7p
yCJjUKC9x9cF0TkZvEDS4TjVmOiwwkLvxBf0AFrczXA2TncCa3DrDdGqZVGv5ecB
IKQUeATionzkRY4tBwhZTEkPUGUv/pGumvmsuUWmMU8y2KmIUnJ7pPsqQw4PwQ8x
sVh9KJRqYvA+BvkHFbHhC7ScMZW+O1goJ5OfG2/i4X4fqrJkbRA9Py+IPMYTEW11
5MNxMLuMIZSkmj9oichYVlObrRhX8LDNa0KUDPALB0BMCUwtHqx/4k7IWFVi7WWX
HpLEcnE+UnUz1heQwtkG2lIasd7TaJ1qvx1mLFd+HtDCUWcTYVbUwRs51Z8+dzmO
Xi7Hi5+g1u3oHq54QrFiYuXrdyB2rtu7IUp0AE6Xjm9O8ZQJNm6aW822pSHl7E4P
aZH0f4NJq/pBTjubWRr/uxPj187QgBzPBhGSWgWVdFLTBPkT5ZfGxmO0fPfPoW2h
sSRiXkXYUC4ykCUI67UEVUD2utKcDM+LqmxMZsqp2ZLxeqb7PXc3ogOns0YVqyAb
HBME7iC+UF4h7rGQFb6uIfR3jjA3B/ITEGATtUMrBPM1qll0eW5MWM/e5sxeF7Na
4c9yIBhTK6TylH8n8eYYwWTIfZ/wDfBY/lazIc7UwDfen2IVavZklOtV1u6sK1sP
QW3jQlHcAK3xLTp/sF9ivzStvHMxw8lVRtNcEhAm5A65a2RQHMAMbZvAJ9C+k7fy
n+tdebFTzNi+Er/JHaNI1UkK7fXk0cxIzk3mIrSs1Nl95+nKC8ePA3W2/+Q9dPEU
4a3+B9ISat0PrCYfXg60FV2CWQx6K26E+Az1SwK76P7twG8DL9KcbHtk1yMCcOpr
kQuNjRLYmyqR1QZk7g6HJ2er1hz6pF5ANVayQIOcAqDQr0Ss4DEKvVrqBoC7OBnT
8D43aJHSljmMQeTdlXDq2w/hTNc9zKn5MXhHUe9TfuU+Xvzvb/frLOQn+YstxwHl
9NxYISN5jpPTI7pGWVBDrjnu5bBVu87h2KT5oCV32I3YP3Bg976OWfFt120iCREK
iBF73cYJ2JA/nTD9SH0pvlLdehufHYBf/HhIzSEPUeMXTguX76Kz6SIMfYF/fKVx
XahxWO+mF53Cw05tSoOth3MN6ZSuebaXpMptfKHXz4KY4fT24lvbQ45PKRDqegZv
EygXBP47hDEXbKQpwssIR/kva4HTwyRfQlvJE++rJVUzWY2iDGKljGJ6ZBgITQSf
l2dR9jiAVT7GA0oid+6Zhu+IVqn9eWY+o8BPtepS2Y7Jytw3cWQcmY07euWdr63a
aWuth6exkXMapPsNHDdnkD1zx4BA4A+pxjhBiZNWTHNF0CTwXROaTzS5eZbXGVlS
Zwe0oJRU4T9/ZML9utCgcN+e73iadbUNvPFwoKJVkgyOdc4aK6bm5D6T4Bpc2KPk
LqnvSMymK8eH0jDTgRMzHzISbB0Py3Gh6ARBBPxzQR4wL9Fun/OYQ/Q+XHUgBgCM
xZn0WnHcs+9HrIzV4JHVHGHqYpfPM44DEoIVMEAAeOSikVh2XuNWFbaGGypELC2y
lMxBCQXiShani2tXRE2fg5eBBztWPG4TMmXAfgYUzpP+x04nvR7rn/V7owEcqiq1
+97nxq4b5N2b9+fOEiRGIjIi/EFwvreGcOe4SQlGTwE5LGUour4+hMNnqx9fXBcc
gT6t+5IPeE8Zypm+GwPg2b52Naq4626ESzvpgXaFg3W83A4qg4yqkh5T+anj7shs
9le0dPFbHIcko2Uzkuoz/KBSGTV4Ra1USWgeSff2rFgCv56/RcqRNM7gTZz9iTNJ
9YbHksEVTHt5aAW5cP2fO4phee3RIJmw2AZo7jP3ILbbMt6AvBI58rKNLs/RMRh9
HZ92we/qD6VjWUtCPwb5CDibsm/Uik+e6tuj1d6H1UafJ7r9fcNCKls+kZ7PENvW
ZKCX6J07cmV4L1Mi+5HuQGjf2NQ9d5G/mCAiKeuvZVhNSvxxsK51pWWEG2CkifEq
OXtIRIf8Am2gGYnVfwM4HX1tR7gnfLH4qZIEFesvjhseLzveIBFtkSPbWuzMeHpd
hVt8gYXNVIN0BuNNeyYkxJuo1giRaj96bSc9ZPhQJfTJ0LoqN2G/jxiEpiT+KBEQ
atjkR+4+HbM6Pgn7rZnsJvLCFBcA4wz9dc+QvHfrd7xno1ux9maE9TNr6OwZszuC
RTMnwuFlsi64VNruEArGS1ZiBiKhetVwcHN7+Uo0r3TG+mD+sgCY5yZjiPo+meOR
56U/QEH7EKW8IwXIBxky3qkIddJjIyqg4T/IPxc7aGkYSPtPjovtcBRifSTfbw1m
w63pn0pREh6GM3J7fr3sOE6FYsqWYNaJFBotAseiZUEDW3YKwO9gIc4Np/9F6czU
gwhDYVhJIgRQ7IpJCuL8r5Ib/efJyQ24L2H/XNks3HIsbO9PEvsEarGGISSJ1IGc
B2G5J1a/IK5/c9JPw4wsHURkQOwkRn/4HIMDdUCEyxDKFXXU3BC2R6E536sr57dM
LUa6KtF0yjDw/uBcPh/4QncPOevJs5Nl/b9VKZ0I1jlt+3TDszzC7mAQg5bX/Xj6
xuOWM7nTAmNikuvy0EajcCGVK/5PilPgh2Den1IsxyP7T5XwMlX/BebHPq5ohBKg
BSaftiimkq4H31cGto5mq7vGerubFK+RiSuI6R3oITEFQDU9E6e3oLT6eY4uam4o
sWa1QyUZQ2tqRSv4vD/QV8hYoPPeD7Um0iNxVyrc0WwW7VuM/CUViREiszRqZE5m
GokxR0xjit+tNgLrxMIUG1TNPG+w6wdUH1Dgz6tOpzaJeoCghNMTXJfEL5RUDMzw
uH8Fub8CciCrLZDEU7X+kzG/QVGa7mU/+swkfJCEKw6ugEWv+KBK2QBf1CYO0GgU
TFy5QdHP5lBl/3Ojh7BIj5Be/nUsnewoogNTPiAPiAgANIMAfAxMUwqn4ms1n3Fa
elUgp+0w27GezUk37eIaYOlp7UJ+f4iuvcRoH1YbBwZHLMhfnSTSn47rJvf0Q02g
Z4yPMTbOdaPRgiX5uTucNki7qQF2TLvrhvrQVUSc6bPjujKrfb89TGWj8+Pr3Asn
Cdan9GlamWQiMRyanVA/kFqIIbURKimIj76L5bEkBNH1fB/bAltNlmY1i0Pzu6UK
c51aWs1fW+awvNd2CL2fncDkboN00EtRLYwDvLmcnnuf4dElYmBNw3hp7yHSLlbh
g+lm2EOPxSBfNM9DsGuZAzaNqa4Suc0/HrNWRXpLoEaEaKUjyDVNy4ZPSJYf0Plo
lqHeVReQaUO1+1fZTci9gycQzsJgtqy4Dlx+evmRt5gzC1OHnTXyvH8TlkkD6WcD
gecoiONcFtxWsnT66fldOx8kwNJXKQ/iVBYaVoO6dmqoEUKf+akIumOzih90mOv2
woLCT80Oh1nNcVVYjJiYPTqvPiHibBGUETDBo6Ko3A1lnaa5YjfDJLzVOQTvl3VO
OsEyZmBX7qFq8YQm5FxlxhdrTd5tOy6a3aD9xoO8t6zQgu6ZIRx8kNetG01n3kms
C9wOIo8lqP3OIW4uV9ikltE/XGKNvhDdV1Xq2jNJd8xhvw/Uit/lSb3UO6DouRv4
fjHCZla8CRyHlLLhmMPwDJr/gxXqFeGA/p2+kVbzKgiEUj9Zp28OmJDKxV5aVA/o
U8nAJ7d7+o07BRB2Y8dGfSvSNZnPDf8aOvU+VVrshm7tMCXYleRy4o1jZm6I52Gn
CCH3FrZHlOrsEWq0CQdfEf8ME9d/XSFwrtXBzuSmW8VTGw8LgRNFc1rqjCrqxxtZ
7UTfJozY4hTjVi7UbaAy1ybi+brkzKFT4yKISmsE08EutuhnwGu68Xi/HKiXXSqu
hZX1A8+Nn9iyOf8xP3eb7Eo0prjBnlIjN56+vlx4kfv1mHPEioiJYiw0m3WVVA1H
PkAWbGEvOvu0pLdnfXqPczuzdjf5g9sPzv14UPJWwn7eVouYHm5UfvF0O2caDDRY
3RukcwURsaE0RjxQBsZcAjdZ2mCjhgIeqYwa2s3lpgUrGHm79hLg97XRljE30oRx
vylYEgRKPwEFDAO2sA8PN1lOipwTtSrnSvFDC2dc3IAMN2jLYBP5OKrhB8GJoAHl
/D+Qb+Ba3uj0PL/Cqja2CMXKzoFAYgyGUZLnaDnX/T2lM3LEtHy2DXiXUpa72lIW
hML7M6zlh80ymlPv7yi+6jMYH0xKU/35QC5P3tNJnt4eY8lzmJJMqOXmoOvJrpSZ
F7cb4QaJ0Lb/6LAVfPHvMOkh5NNRtzNdVmR2LplxhcSoxwW1H90LKxWCWooKGvwx
M6iLVDtT8zSC+vWso7+FUL1tdPeaCKJ40WARS9q1wP1X50PWhe5cMy6lDWGDl8H7
+jxQdACNdfJkGGFLr+GKyALY7G2a0D3l/S2nttcU4hpNyPizS4B5V/kB7S3ZjXno
Wr5ippF7vivsVgZ5Zu9daod5KS3qG9YJVLlL5nRvt/BjPwL5Hy1x4eN1FsZF293m
8BfswkrUNFr6jOJuXawOQR/08HR+IFKU6+m4t7JoFmKF6GMcsu02AbiMonxIngQT
7A9KjOyJLJMhGHDwCvTOljywrraQy2FiHJg0a5XV9Qj2tzQDR1U52Y/vBMwWougz
mIsfHoxBptrf/1mSk4arkmFT6Qo9YAVbRUJDvBUkA2BIaCRyngG7IjnsxvpFrxG1
5r4QrqJnm3fCxZo8nIuXjIz3Z91YG6Eg1MXZkjYlukra1v+dvmIjWKE/Sy3GtNgc
KdmuiKKP/PiiEWlvJAcuVNMhTWPd/WbWbe6q1zUcjTpXGqUElQhetKzNUsN+ggUs
+3Nv+e6HNblFDs7CW5/J0lh0rVTyUDqythaLL4C6Zbemw3jU38f1UwvxvjbNM6J+
THoh6JwAvEUA/qOUA4fyY6ox7i6+sy/GQG3mlBjAl21O/aOvQiibrublzGn1vi8I
/qy3xLlmJ+l4fqynbuFd48CX9KT1CHTN4Q9xPj4MRFmOhz1UuDb4N6e82XVk3zWL
UmNezMqtKZhV5aanhwP5k1AcHIl3WVsDVHeXLBsXTmp3PaRWwwDEFCf3QbTLOLov
Vp8R6+myDsyC1HVNElX3j9GtG4DOzU/Gaom+MYtGzAad8ozqGX5wGdShV5RT/GlH
Ex5gz2ih4uAWgnCBcw8bWh2ntUQhG7IG4HPkz8K43FhCwdsF3BJMJ8UsBynqb88f
ib5QG5dPnvcrw4EOhy+qtd0DHPnQckfHUKWiRa2w7NFXFZ7XcObsoA/XF6rUALeL
gqpzxPim0e5d1kw7O8kBpXKyDWpBgcdJTdl8ixJBxjQ3yGWwfHxDKFbFLUtUUlQa
nR47f34EQkkeguQcos2TFtEbjmAOZ2xi3S+EGbAcj6tUxPwIiDsag1dORh5ghbkF
lnv3wvUm7J9QUBmpKzk091hsLDTTDnIIBJktI4Jg7VDT4T+6fEBg/61l6kLdqT4o
xSwx+Ph/BsAtQklmFu9XARo8kCFgGwo+gQmysbe72UqtY7LVoAj9fdu2nsk3aWID
lqpfTgwdCKq3iaPEhAwqVzOrB0jnX9sXEuLYE6n3N7CJVh5oaSDRt4FVUoWbUprg
T0zLc+KczIN3Byc5M6s4q0IEhpIyYv0ITTfxaCs+kvF5CtYiv38XYQyYXtE+5J91
7Bt4zE0JVv4oVrBJTu0w6ktogfdtIuLN0BBa9zJfRB0IG52SCFwGmw8KMc7WGHSY
wI7DolLJrEuhLmGBIlQXqopQ2ghVYvP4x3M4kTaa4Nh/meAUgMJCwfhEb7QVWnR1
K8K2CIEATRtP6QHMLOEzc/0uqY61uLcs3uGmfbDa+Sv7DG+n2NO5G998+DlZ58Ii
Qy0kJBt/Rxi2gA5++5uJqPT0/4/Jg63G5qjJDptxTeD4PHd2/lPp9o82/Wt1c9ps
V2pjnm8gp0QsUmbnBhHCjyctnceu0LKSSpVBivNev8EbrBxYWMWt0jgGvnCrTmQc
qGqug/5sdtIlLS2yqHhjAfZ4LbvlUevaId3ky94Crof+SmmACBUC+U8+vNX7/Gpp
sjpu/KUspdTaK0YE1vKTh5Yym3vgfdrY2w+8YHWU9BuSDyXqytOJlBL3lTSzu/ae
mseTJf5iL+Qe6C/5loWTlRclHmbt00RTNR7gtU+wVL7aLzsGFq/ZoMFntu5Cb7Ec
KR/BQ/BquqmfJdDoL1i8gowtr4zyUaALqSICUtD4N2yeRkq5MTuMNaKY+kPiMlVT
wQ6C+vl4wiWutJQy8e2grKDKXhIgLj1zovZQHZvhjx0pMqMHn2tFl/XSrFuWGVHZ
ogP/JKJzB0CLoYdcychD09x+dAnZwjNYMtlLkFxJHoeGp88fw+yPYOq337XwbzRX
BDuDhd9wSLdWEWQQ7QZZxuR2bepblyeoQpc3XhRf9ubqjoIcFI0Nt1n1UQLKfVIN
8qrYD4Zw8u9AFP/9aNRBrxiezpwm2bo16bO9Zjw4cpw8PX1klzSfaWwztAhP8Lj5
8SgnEY0gIgDC8PPz0ldgo0ZeADaWxr5qYxBjbXHaPbhARSrQAg18AXUJZIgeBAe3
65eVeVsvw/E+x2nPwans0IXefRbX9dGlce2kpW8/Z+3Iov2T6afp6DvfG2RyJtlI
wPpxgb1s1obV8wZf5S9Z1uMzISsndZq3CjP0cFLciS4ICEC/lPiTeGetnIIEaat/
G4yUiZnq3HJW69eCfnyKKOHig+kDU5VKZWvh7sx5dZcIE8AZLkCITCZr1lnBzBYQ
djxS4oPvY/Ma00x97/MnSggIib0pbQ6ailVnZiltzD01Rhg2VM8SZYTR6iHac1yv
fXKC+HsM8sCAqqOLPMASQ9VW+FjyWjW39SSxGZ9/z63qjexxqRdCwMuKmS4qrvQW
4y2YZ2aydXI/Y9PQfdxsMp8SO6tRZgn42wcOVAs4lYUZF953MkiojBTqvD0lRmzp
7KR7xQrzrQEjg+V9OTMxNfjfzZpvMds0U4MabmlfGU6pGo9bH7qBL/jtCurakbAV
huJIu8InpR5KH3Pr35D8CLHFL0PrXX8Tuzn+UdOaD+OYaqrXTjHkNw+NJdzg+NyL
hMC617nfPPpFP99JzAd3nEKN7saz6r0Pj61FnSbsfU6hRlef88nZ7qcXjyW6NlhD
UtJEaS7YKSONnu5OYbaLMTCAx7TjFm8W0ORJpOtJXGOl/9I6qMdsvQA98jHHUVrQ
oufarfkXL7KJ9Ln3UCKCJb1h2M6u55GiSqcQ6myhGSOUXExPUFOF1qgt9W7NGSFt
8lhV9ginRPqNj0Yeh3LiWjKnMXHE0fGLxl5XjWNvBPOS5qnubL6UDjMLF09vcRDt
syk/GnH9xMo6v6k83rgnqEIm8WdQQJs17yy68uGKEeV+ACyn713zGQR5eJi56NFe
PAeH96Q6tocETZ5DM5oFM0wFZsy8D3esl2ijpxyRs1Fv1lsiBC82M4zCF5cM42Iu
ukPIM43Y/gAUqA5f/ZAqHl37LF8uYNcWQQI2T+N4UfU0V/qSEUTGuYQFc6cXKgBb
QvxXg802pW2K9Zv7MIu+T4sM8NJwiFedKPTpWMlM5N+aGyzBlY8/Z7olWyJQyQ5r
JxFcETeR3xk0CEfm/Sb+MDjVtowGXikwcdCTRG4fyCVDthRM6crsrZa/NCknQ1LH
pullB1bWC6pcdBUdnjYFvR8AOl/hWMyFKczIjHRvmBRUEAHIpXuNAmtAZNkTOUH1
z5MzfXUvOr2GmwZR+ZCQ9F5dneFqG+TOG/PCxBbXMAc4QJCPQ6I/bLd+6hwfjCuf
4DO1dfQF/0m1VWBg48SNnyJwBn57XBuiN2xQ4rkaVcJfIuNjIudMe8fAwan24ZGH
CIR0Hrz9qRgmc89X9vbAMBOmZwSQi6bH9m3gA5jSgFcWQVdDZb/1GRSQuL50iKPV
1iG3gvdSxG01bXKOA9ERpfQT3phCZIJCI9sjOycs7SN+HKcnuUxHvJWLEXRzULnO
5seDXdrGUAv5pLKypKiWB3VMEW02PurDdjDjtyaas76fQImGcbN7yALWLqLQVZSF
alZ13l/ArltjLbtzcpzgbqklKNw4dbPJPKQVVIqyjEk1iU52ed7AXnQA/Dm4pn/7
2ifPFlQFzpUZuK0JTzOWb2hIyH0eSy96jpaVcHfPsnSVwOXeFjb/dXxXnYJYm4RY
cnU3uTTwutz2JyA/KV5LvPSnai7syrOcOe2RSJ0DCIGWeiLuT1z5TI3bA1CvfIJV
UgkYCCL+vyNRdN0CUh5O/XY3k89ikYey6tWrm3enUYiSMcFCCNrvbuh37ewXVTtj
pgD1fF5u1O6qsfiVB6PIW0WOR7ziISqvNGyvkrVHBhk0riHyldbHrJSW/Fsroe5u
j2btijId225Eir+s4tDqLLIsZTF3xh4HBMy/zk3vOqLiBgiZY5SHXwKUaG3qg186
r9yBc8QYnB9xv++FPG/kFxnlqZOBs1s45ADcbojEFsPTNYFwLj7q/5S+QrIBYUM5
TI31QZcJ+/53mYiJeEjOXTrzYCVSCbkF1mFrAD1F1kIP/qgOCo5A+cQQ1IIwtfR+
XQGYkccrnu982dzhF/gcFEI3Y82r+5wfE+IyJzOfC22yavxHS15jqQAWL1jRz6Ar
SyPZ4jfLM6F4TDTzhs71QbRZOSpS0Iy6ZYS04jDO0JSfo8LGJtvJXe+uYF61NKDL
+EYDkPT+KA1g5tA7hUXp9xmyeMHIwDhoy5yNKJyTPk3T8J3JX0jWFXUROWQLPHfR
1LbvvalUymF7zuIG8LTZLJ+f6MYkT7tH1BDM9h5loa6PBImm1zrKGC9s6bwEhgtr
wW5TzfkyHkPzWS2V7IKyB3ozGg4fBeTz23iSZa9XC3iAskXqAWSEf/3bBAEEQRHo
MtDMZTSXYN36KpQKLjAopleezl5LIKCFjBbNmhYwC1K4G8n+oYJn0GAtsN/+P17W
AD2BP4wAKMnGX3SiHDViwoqpHNrTFjDQO1wn2Q2LuS2wiYQbzdcgKDERkMPV/uaM
HfzXtVYQInTkhyB/DNyKm44zvuNG9tixK9kGabJqtpjZ5R421aENRtzpE9PReaU7
o1jTbe3cgie4ttNnlLif032cAKycyBTp9yESDq0UImpiAGWpHp1Vq5jA7ZIAX6/9
1H9uZEMlXyvC39RDr9hG7NhulGMF4hIQA3ZodkilB31wyM7t4H1aTXOI7JZbHHuM
hSbsRqMvyKquxXwgT7PbWyRUnr8eT5yHylkGK7WfJGH4bprlext2I8Yn5FGu+hSd
WCOIONC3DCX+4zQSPH9LG2X/epRtGwvqzQ9NpU/T3RqASKSoNO+bPtBTM2AmSjuz
2gQsd2v/99+J78lvHR2CdynaRxRLDQQ+iolY2FvNr8sSuvItYKu3GUcS4GGoePAg
8gxF8GYM7F16Uv5tuYmjURyhp6v/4RcPDSnHmZ8jtHQ3XkeetAsLtrdHzDVkjhbq
2ukKseUrGAGErKruQCBKpIV0sk/i900M+ko6VLVcvxf+oDNuXq8gkubvbfKcpmUj
yzbvi0yBU5vl+6VZhLkMS2aB2bL6+Qd4gmlUaz5b11x7D8qD3WKBqmU6Ywkv3Glr
CPIGhaVbO488N/xd3J8Lm3HXol6Fq449mmnbn7/NV6HJPtbNbBJLbRd9dSMkB7kK
fWZlezJo11sTanVa6topSUaXwnp+dIIOal2oExdekMNWSAs9b01el4fcXOcq18Li
Qm6mjjrbo5Z88n2IdU0fM8xhxX5vrwQeEH6G52fe1KbRaGQKNjn1PfIiE7SMYcKN
2RdboPauEgf4S6+P5+N3F5QmXVJ/L/rXrpTwZZjrNs0i9ByoJ2zavaaTUj2R2f/0
7dhz0yxYlnbmcbypYXZ61AvxlfYkaSuRAn1rOIvAR50bzJxoQ5CSd4ve9VCLw282
aYHMnuMMRtgsYu/e+8b4sQKIEPmZ6ddrn2JCm/HMpbXydYwFcUoetyMQ7zmJIMi+
fZwBVPu7/G6gfs8nvauXopxiAwtaoFvbouOnkfeJiLFbOX21kO7vBBKMZfICDX9d
f6wold0QhVRKNtzxIjVya9vGjGGIBBJSEHDx1iiqtNJ09EiDkOofn9humAYAwTha
1VmpROToGJyqD+GVCnBPc4G1lHAvg6SPV5izb2vl+hSGXGrSgh5qJg5ej7CGQKeG
AlgAYg9sOu6HckZ8qykNlP6d6Ba7TFHhXa9q7kDwhys6uUvDqz+Uqgq4Zndlh/JQ
sGA87dmAwzGCi/xs9Hyowb8CTF6X4qI5UBK1oLaESvjSNmvxKNRabkaKzkBl8RpF
lM0xxq9+sTrh9v4Yf9TnftN4Ldb3rYjjsuSGP8HuAJMi9nrhDGD30gTnIyninO4/
/PbCIs2SqyePRwRSK5MhYk5R9J2yMWF3nfujQvwvozq9b8AIsqO24WYYBTFJh/Sr
E4A6nTuombDZXniY49iF5HmC+M1TUNbJ0UEo0OshHtgP6S+hImXicJ0QOB/20CB6
leIDPy8RFZa9x1ajYYaJr+eU4M8DtlTRoozYn3lVo+EwZ85VkBIo2dLWxQr+fMVF
wKPgdLMai6F6Dy7wyXVUqtooq+z7P0xJYTNTY2hQyvRTP503nxQo+tAxAxqKgsvW
kqV+y3tkQk3+BWl8te9othSoz9SlVxP4GS2mIBI2lHcMKYvys9PJp4x/YP3ooUFr
1WE2c20IvnPEivDgr79iafuFuV4B6HyCGTNPUupCnsYQfagAP+G6LNlZCWX2XZ+W
faoTsPVWyDiS4AlSPiCTq0pBqYIarrs1aSa7U3QTysuIseoDET89qICVm9YtjvJl
0JVYOn9E/OERjgC3PIPOHCTkLkZqb0OYI3noOPU2ZQzCxb3UuF61f6w1Vbd523NZ
XWzpH+4rl6s5BRZNmJrliDgr7yui1C48jbREiNJ7iCL5VHusGHHuZmzkMrKNZndY
BPw4eF0kbjCJKd8Co7Sx2Tkf/DlJ8iCJHO6Jjv5K+5qh0ExGe41ZisBMawSVapsk
k8vAYMWbCf59POlsau/3WtYfhoOnmCFRz5VXG6axi60l0kDj7ERZzjS6joAJMkq4
L9SrayMVFT1kKi0FHdXUJTGSomP9buwbm8AM0cGVzNWlbCWyOQWWY0FQLK+dBw4M
jSwYNABY+9huUq7DQNYP1zxdk65r6/hKJXMw9JcpuGh8m8B7gAuMaT2Y0BhvVK8B
JtydAJSNoJ+S8GtgseJgaXzf8+nxcEHZqv+LMAgNbFj9uT3q+afHvtXJG0FNulUE
QtYJbgY2jWsuIIPPHtgku0LuHb4oaUN6Ufg1/VkVfydXitoQQWviXxS+ORRP5t6o
5zZ0p3XKak3fZtG3zNT+j0g+v64P9k3K/XsSy+zB5Y1FfP+DIVjGScXw/OFa8wML
39XFf7nqph+BDQNQldpuyZIAg1lI2M7YjGvtxIxTutTtsXPV42MCMm98j4GC6k4d
wfc63XajVuCratqcDawCe7ELPxTowden8VNNpfL/2GJyeymY1K7yYKwXpIohvppr
7T9TEuRYhU/8QcBAx0tSyqMhPURE/kZvRitCuUJS1DSEoyWKQvGtuVV7akfRBpDZ
trdcw6vTkDfg47VCDMkWI13JX92Zuv3n+1LTP+bsNo323LLJnF4OVhlfGZ4YZ4fz
pB2CBFoLdn8zVUJxUzJmuojyCJR93Y3gjuUj4oCm02XNKuwOf1sXHXHZjfe6EB9b
9cY79JeE8U9cAhKfWejbGggQ8WZvT45q8u8AJfOL1AZD2NW7mB/NHrd2+Iyu7y6N
DtXJYZR8JlFFMHiE6jd6Zap2GmHQFxMI9f0OnoLFuCjU6fV6PrX9HFM5FwvIHEQC
ihGea4aRZFoBDxAbgmWuXXzozJHT/KGh8tU8eE47wMWvAIvr6toXltdwigcxbvrw
URLs99x/d1xXaRjUc6/jqlEDYy2kNGYFqpha3MPIZjk+nmLhbjgJRx15k/zYmevo
3GZHQB7ZxTYhLxKwD1LINf2sAW2qTKmwHkkqVoEMckXppeCqSTU9uYTvzUEjsEQQ
FIjRnzMIxOXhGTHEdhgjRP850t4i/W85BHjPlYd5tQXgNOwOaRWfkNTUiI6tTemx
MQGbn6clfzd+QQWqd+XH/9/ZK/6vD4va2kM4blguWjoAzZ0e+nOZfpm3UIV52b1T
zizZI2mQWsWP+ecU+4eoJMQOl+Pzoxx8TM/TLSeyQY6GCieSNU5rPimxNTfmwMze
l+XMP2m0gEpLgT9d7q1Il0jkv9nZ+phLA9dtxhrXFZEQ50vzpVoFzRd/2VJZRsUS
n2ie96TUYPpiORCJeAov2qqcg5wqSM4xKYN+8U4kIANGMFVWZV8C9WxfaEIC/avS
ZP1F4LxEn64kjkKR2O+5hz1Pzlm4yd/OC3/hoYDFLYif1/0gcdt2K75PtdDUQfop
Sqis2fPVFSveIqjE8vgo5UlkDoWYl74J1xo3N8K9sn5+7VYz/j6MzjZmpUApd4fV
b9nU7O4mKLm0uOnpf41zccCDCWL50H1UwPrnKd/gnZ/rcGkoDFjevOzcLTYuccMX
SXqxbaPD06ezi9MuE/G8iv7/6Q8u1YyvdXoIDI0oGm2eYXkWFW0fDmvLOUlSpzsl
iBvO3+Xrv+Rj3aIHLWuY0S6EerCi4cYEoAO/1O/D/XOM5t/wuf4TrXi8JrZb+ipw
8KpQsx2zaSIrQSUk2lHzzO9eQsvBt/BfgZTAQSRCH3KGaCSnY3wUrdS26zOtlrOs
80O/Jy/fKbjh4EXtT71XnHMJpLal6WX+Te0InSOlghvDKXCPPI3HpwTBApm+PnRW
1YeJ8pKunKQ64DB1VC0TelsrOEHE/WkRUfDsyUmoHiJvMZDl7sXi5K34iGWZoi8S
o6dSsJkUz2GaJv5rTP7M+30/dfiQJuSo1lTR2WPgCDY52WTigz7dJng1xXElKEhU
a7foJCvmxRPR5hCmkhY6NzTpFwZLjLoxGKZEiO1GFdXgUg9VCD58VsD3UzZQx0md
B1dQDagnG2ccHuv900tzQclavQCnKhyoqzcbcUoqLvMyDrgHcOjKzTQA+D/xhsgU
MOcepzPpCVU4jVElMIyPP/siJ5oosaxtMDBhx2nModuMQKNUt4Ma3Wy8hghs8sCC
Et2URiCoZI0xVxiT8Zp9TB1SchyOYYd49cmBOpWynM0Ua5XogB1NaI3ch4iVOZIQ
Gb+x4MYYAAQLrwmJPvptYPTApsoOcp6VskOLhQXBH6XB6vktwv3T5BFaHQ40xyY8
4+gMgtODq94olTlYhVgu9cyOHLrHlU3aN3j15qDukJUlK3CVBcsr3zX3JOyYYo0s
X7DmfM1UVXH11r9/qd0mgKc73EtljzrJa7pdpRW9lLN5PKfhIhWiika+Nbi5ud0z
xDUgG+Sb0Hbf/SEO/HhnRrK7+zEQwtPzevHuGpi/OvqYaYR+phwpuJoaRWW43axR
uB+FU5kHjdDCEFcFpZVbsUkxsNGWcGcFDTjLhbfEgYllmPQ65LDXVsvpEFurRT9O
nHq3E7Wj+aJkWqQHQ2ZhnMbSUGX5Xo5q7274oEmhWW2eN+e7hT+lfrttNdCwZiS6
qB7gsHviFYWqED87OcDoHVEi69bwdjYVNR68ZEq8qOXUXXROLhzdnWO08HudYstg
f8drT1Qoel62ijnf7W2AZNBhMYZSdus20u1zHNvTHDCmR/j1B6+PqgPPbGRphcri
Jt1mehuO7dTADKvJ0jm6sZkbbZVM8rGn7cm/CiFhj3EKuJddEWeD2veiOdNpUv11
gBvjtQV5abLANOgU9khXeEbIDIcofLJWREQbJe2EjwMgjfTSIbHXxZwfRrPwikbA
GNqDIm0ACI9KePogENDj+kC72cw3zWjYRk2oNG+3r8MJjy/Zq50qa6UprKGoKXR0
pMgA8GpIbqIEn8R+3MFLjFqLLKHnmI3gVYSiTNB/S4RD7VCbrvj/h+AoWZPFjFx6
5rigZpfRf5PLOI09yhcgCh7iBTTWlye+Ty6Huk2vKIlToL949TkRB2exEUo59RAb
QQeZCnR22XjQ2v9bbdbiDg9OTTXemTWX35qDOBHTIxdg5e8fmcZXXT+hpM1NaOzj
gC1Aivk9ad3dsQqMzd6TxnX1kBoqAF+Ey4xv2Ya68whWAHaZK+171uoqX2A64vKF
3SqjHfzJRiuSCBewb3ilo/O9IW0n66L+jd88gOnSBck0kgqc7OA3/9cH4+Dwcsxy
M/iaFUHoFuOfI7WPJK2NLHvwWJDew3fcID6aZKrTlAjBDCT4iz2G33C2vU2BcPcj
758EysrRtZkfOUao/FSwVdTekPfvN7C5o1lWxiqcur1naywtMbyV6nWNbiz6kkzQ
ifb8B2DPncjsTtOUlmVBvVCD81sRhO7KafjoRzitirYGZOHS1H8fSrgvFMlxVqre
Tq3WVf3SWSHlA1GqsXUBYwoxMIgKWJCjeZi1H0NJt+cmVHwOjGtBcJ88S69+Ws8b
+9xtOAjPzjLGscCKOwZvTbSbhbDxNSzy0AJmYCCfAqoZ9yknkhBX9LNZMtILBzR9
GjZF5m5CBMjOG7MbZfhEJi/5lb38R7o0IkCoSkxQTOLltLvVtM7cGubb2bBcOmXu
CyN8hqxCQjGHPq1GTzSqMj/E6Wf6Z4G6ZBtejzsc9GBd1s1MJ5UfcERXVRJSNPpS
8s1C3lqKlJRraa0vFT+a16A3cUaixaWGVnwx5d8cmwUEy9FLnWEIVocNRU3LN614
7fDYEgWimwislYoPc9TJVD5pUbHGMj51bp8T2Q93BUJ0KmskmuW/cIz04yZdd7SG
QRO38vK+XXmBkYmaxT2ktjNcd6TrUxfGYBkQkpUuHQsFlxUaEJTSRLZ0NSpB0I/5
N+t+HUJYhhRiihVmbr2hXPjIgG7cXMX9CqHSla9xyIlr5dC40IcGwiEvrJMWPU9o
XJpn0FZQCcG1fGmLuIgqvHWBWjYem5Pm4AMGK92QTh2R0niqi+fHNFrV82r2CC5B
rzJ7W6IitAjOepkVw8ojCjwNiJEXFIBckjnnNWjwJ/uQCppH6cewL4Omg6z0wXcF
gLRc4ap9AQkGIuo/Z/rPElCKUiNVUD1UD1SauIPMyFN+yJkrRfg8ozzaejH7LUT3
1MOLAgsn4GWOpgKPhnSAdBTFNS9hY6ato0+A+rak3S7zI6v76y4dIyvD5fMx0aQ0
ez0Y2fwaewbWUs3N5jX+WpeVG/TaJnZmxmFLeib2wVgKjGS0j5swv7a95pYW2ADT
ZLUwo50DhuLti/WQZ+bx8ByTaesPhn1SFb1KoraQyuqhlscnyng1VQOeCANxy3mi
U8EaAKoCj+oqdcLyumAVap63Kaj727UJ0s0iSvo/Hmfofb73gMHj6bjXkzXkq7Yn
azpx5yr5c+M79ZN8lFZGmI7uNNp/Dx7CVXh0WzV8Kp9SAJrQ5QKykIngJGJq1h8/
3buJweePwPhyrXliVIj7uWDXUgHPFH5K/5oxqEBFT7eGY4e33cAuDwi3VfS0HKx5
NhIKYkazSmk2G95pqF0fjBUiuRw21tRoUzIkBUDonw+9ld0xcRE9lgyDfVFhxnXZ
nTpPmNkCw9MyfqAPYJqn/ijGDOQ7Xy4QrdfF1F3pzc08h+Jp4r4cP4hC38Ilv2ci
hTLvM1UyH2DTc5Dc0iK0vkrvAJo8T8RWNYqbub4IjEL0zXSwDlNmqIsV5gqjYSqQ
GfvqC0Su+XY3H4Ooa2za5DB+P+bt+ULWq1/FsTEbKJ+LrMsKtS9q/zx/9O937y/4
u4w3Z/f/BLTP2zW4NBQQqVFgnVr+MQ8TZUe+Hc1slSMMAJ2yN3f/4LAXEn40MMp2
syztOLvV04tyTfqv6v2q3Aw0T9hCFUD90coR7Gt64Rwybp+OdeHdC8UpZ0f0TDUs
8zaWplibF6R7RmIl+062uNyO/RdmGetE3lHvM8uUa4gm539jJAcKRtPBzAWknAPK
q/I7ufQbZu+6otf9eSut8MiHzZHM7OZQG3OqZlelTlOhx1iNxJO0vhHekNqcaJlN
QZ4geRii3WobQ+9w8pMZTi0zGRaOwlqaqFJ6/S40551y6Bv5dkAmSEesRhLX+WVI
g4HZE2iLkHFeU38Myh0iQNUZrIkhnDC4Nw/YjtMynKMux/ZKFXYe+OdGX22XUdP3
F009YPRlpTgwzHrMSc3P3TRZVNLAIs/DipbkVWLqlbMrQ5o5CI2JNVhVr4N9QEfI
lzG13vGZraD0uoM01CSsRQE7vn2SbJSePAOibghnaYXQQWJkeeuFsMDusldtE4kd
iZ/+8WfAs/8iupoPkgsCTACIwvEav+AJLOTAvKq/DqkeaUH+sDDpf1QHX/xxs6Ux
ne73eoXNEtRmsd3tdRgfU5vX5kNL09tDWjGpKB040SkMqh2P50IQn6ObsoLitP3V
hUd5Xty1JlIeKc+wtR62EpXmioSv0d5q05CoO4Tgcwcqekf7yaf1zzkbd9CrNqk0
mE2upx506IVIwF2PdfFlznyrxdy+rbMmPocw/fXTfS2oQeV6aljfuz5kXhBPqCqg
cTDQ5xgj0o5WY52/AtO/rdyr3rDVqVdOBFbH4G+T0Jy7ddl1Yrax1kgoFYgbBVFC
XlP1ocmLoOV/3itoBZAGR5rIs18DbjjhnEdu6pvXo0ieqUuRlBSGoyOJhwjM/TNG
SMbu8hnvAxx7FwZXYaXUzwe5NUsY5KPkWSbYCYM1DeY1egBXBLNOYW33jOXEX7gY
g5rRw+tfofmqNwkYfl6AmEmaNCk5UZTM/c6CW0caqsbc5lBDSussGjQbgvJ+dSxu
pbEq4LfxzDMi1AIy8NWZTGgX9pQVX60OrPODW2zBMsc3EHk53MbUrinroXXK/jG5
YwEaUxE3ac9t/7cS1ChoMJvy3TWJzCgejhsNWw6a5hLhKNgHYomK3hrcw79sPCcp
UA6QfRyBEMzr6JnL3PkcnKPVnFevPdiDVyN0VvCK+zRNOx3dC+XOSFDr5UL+Ux83
Avb8e/CbbpcNrW2GufRsIa2Uw2GgHNAMztcQzma9aAYtw/kUeci7J0C1GP/xdOj5
usop+uuEhn7MW33KyrgzOFVnfSBLFtOeNsnvji11YSx/BdnpNBq//+/gOBwwRvts
DWJ0n4i298hhAf/XJnqNIR2dChhqaXxqqezww1iZ6sBfgSqYvs/aE7B7WwpsSQkU
5AA8oLxod2E+75pHtxuNiJhnJgryMYnKlHReV5VomIj+J/jabtXAPzP3FYrdeEwQ
9A5BE1YvulYOIyh+P/WiA+bK2RmonwmQ7q0eFTENsOuedcH4y8pkG8IySBcdw3Sr
SwA8nvigcyRP6LKJ1syIQpIRhlr4WfPJo+avV1uYcutLqZXcBODdSP+pr8ixTHmy
bCkAQPWmLb+LoeuV3SW5hTnLPKlDF4PZFDaqndQ0xtruAhwszGzeioMueU6JVXqy
KquNfaprC0WxcCOuTk9arIL1vpsTorFBlNC0D8ZznGgCCo8+pE4MsT1VcUh3dj6G
tY0WCh2IShA+BoJpQFnnjNedku91dvXtzqyWfGgAdZM8FCI5619dArJoUBRv95q/
Y1sMahX/Jbo+epGPW22Txd+h1qEqDk6J+LFUaNY3LmcAMPbGplzkDiwzJFm6GzJq
a00ZeVX7qiII+UojIiQ4j6zGaXqYlDj4ZINHKRXNT7K/aaaMpcQ5GN75oDBmR+R7
qK22vt1T9MURRgpL5kM7jgZUHNGqLIt0b6ctlrZzXltoDCarc1bJo3QbfQcYnkQS
HyqBJAH8u6DFNIMv7N8hbqdjVT4Xyf3ZlqFqEd1t8BgdMhO5SmiY7giWJi78IaaQ
kpRXSDzAnLgEc7VyF9mvvSN+4ZO7fRnyUVN4OgwRE/JBMrziuKAMzDj7SIWvOvku
rGyetOblELQK278CaHv3pTZGBWHLjIN4xIAbGQ9l7S1y59ZMTMDoJqaGshTbUMuE
aj0/H4lH3nilzzZTf9aSBXWqIWad9K8z+RlSiKMrlQwennk6m582ZAYgN0Jl0qCS
wjXUEIjmYj6+IdEclKqsXYtM9APl1N0ri6nC66ZRtgWGRlfwGYyOS1O2N2fByM2p
PYeo4RX1uBwF0DJ1uNigjc7aVokIO0PwC2lgNLEoBJ0iI6LF8l4gZOUJZvd3erJr
o7f1UYeSc5CdGFn2Zyjp37I2RphlvhIVOm8b1U526yt5HvAM0kokVbQ609vNRXk7
Q8bK44OtYkw8VVWpEB6HRM3nBk3bClq2yOFmOMjlxZu3Ykv/ONjDBYwbSAorYXtI
qHXC9cV+NNXyY/t/UoiIEaCOtdtTJzbItjtZSiKuYOc8gEuukPfFANMSA5l2BKsr
/Wpl7Z7O79qUEz2RcLei4s/H+WiWSUYMQc0FmrQg4aGOApS/6Iy0Ng/SbEwuv5oV
bX5ZxcU9D/N0qqdLn/geKW2iY9X1mQjj8tbowBWOMYNLPR/EY2f/m5zSYKN/pV6v
mD+azJfsit0mgrsWTt5yZ6ITR8Rduw6W1Mwa8gEPgfz7tW1YZeURXP2kU5MB4z5X
CKSLvvQ7nDB7fRj/4+fnWwLB9fE08L7nRI2Ml7FoUj3xw8RG1XXk1r+6wM6ZnIpd
7yOwJNFCdtrihhoAvNp9AUVzS1t+B5tA1SuQsAxeZSiDoWRACQcVOHxTetSGkcci
i9UN+toimP3MaDPi4xecEUZg1g+VI+v7dB52TohlemNC+XdgwHX/V4nNbhzcFFJJ
aH8Oyo/3+GL1U7PCgcurKtBmf9BNiD4gOAEhIbzIGG1EttcZuiKYIn/3TeHc0+ZD
1ZqCSDB7JAMM/o1TsM87y93ZJ92/lzlN/pisJ+RSLXLtR6N3FSy0gSx69+WysUpG
oYwl3ICWEx1rtIleXBUFuZ/l9jfJVvHnp97/0b6oDDRSxkRbmNNKgWYzXvEwdlTk
HQrZLsLNgiIVEnYZqoL6f1BKn0ZES6mTEtXELvTifMZxZNZ9Oj/H6Pu38o1DnhDu
Xs7IYIIBPy5xmu857VTdbgWHb8fnCPH423wkmOZYfvYS5rxzaYY3IoVgm0CN21xL
qH4XZlWUDY9DwGHzM5eg4mxCmEKoBWRO+FiW2IzlKhekKjbHoc3w3JlYtdVtyLUT
qmLIl1WES2Vh7bfdsB+S88g9QIjP29OOQk26U8psR3K6eb2XEB73Bh3sr/tDuyCA
DQeHN0I6HqPQmR0jGgmWJugVZ1ZE/xvufXSJPKBLH+pl2GI/w952CNNonH3QiNGR
6snHZ2FHIW4xtNzzdqOF99U/Q8Fn6RhyrqfWlSIUMczBMhQhV8ZImmlzq3Lf72Qy
KkyLHZRfNjoTxhhgUV/RTb23nz2u0OBGZLiNFpYRPRnBiar3dGCtNcaFbuTT9cdF
AG+jEp74FIZeObag2N47lTRZg90TIOsLHPj5YSd4euEAoIcR2IOxWJGYlbgHgKFm
LMPHuWynHtJ0FAu5jsA5avizKz6jPvxtINlRZalW9pf1JeY++GnqA8JD2NeaivQ7
cT8dpB/HCKBV1YwU+kkv1VVCK7ORWfrsV6/jZ/KVl2fWXawAi5ENrWdOO15LEfY/
4wMtYfXy3lLlXmmYXP1B/UsnN6vhsOSkA9oV8qw7aAQhQwapsCgExSki0TO2pSJ6
qMZ2l9qGLBHFB46OwNA9ex4WvEf/0iQtO7SpkgHHUixCd6wUXR9evMKO9n5bujTv
wWgTvTC91T1+fb8IItQrko1gZ7xkd/5jdRaPPn9Ju8Lt/M/uuf1qOXgFXPyECGxF
HRvCdg5iEB+7n5PKuK9Q3/lUAE3ys6iCgzXrGSxMfL2eMOknATkHmz237YkyQCLF
Z9rPJp0h6ltiIbmrmdO9uulGnMvq/iioLoqAOEsXeJankHNSY7wnGQ1s63zuBUq+
/PpTaCZaDHKn1aZoVZvKxT8RQpFnLBjsPT240+hc9pE+JmPIYiXV06bfA3dGCjwL
1m1j9YCaUNkXeSjm6mDPU/vtUs90vRC2QBJGcQGd1rXKhrYO2qi0NHCm8YPOBaVl
N5A9bxZOiDG063DxtUiJUd+YceXBRerUcTc1aRTxgwbD64scAQZemh3/DT4E7ZtU
nNvgptFPoeqTwwZCsDkFtTiaci/xQ2NzvAadbePY4pmGO52XuK01xw8hSi7NLN/L
3wULewWoIdpt3+zO8GE7lHKLs/bv7ssgr4dJiWWp6YMYKJkoWWCbTBcc9SZKp5cC
/52iDaq9+lNZ9lFNsHG5x8JPzqvYXim9JTBBeI5t+v3UjYXG/wzTdWJrJqw2pcfE
ZacOfYriIKVXxDyN8F/Acr49araH4lYoBbzPOh21cAcWz9J+MrXFytAtZdcEtRSm
FX4XuzslbZZ1pxJfrCjfZvSnrVL5cap6ntb5u8HAhC+TR+sP2ugQS3dk2mAWq61+
EzSKbb0UbUhdZA1aXVxKInzvhzXJYOkkXcCL3F16EvZKLNsm0CwHBjU9wfukgGt8
XwaZombsq6nIcV8rBAEym9xdwqkd0joxGC7v8kruZ1fyGVtfNx5AeXOFS77cde0g
bIy7GEIa3Avvht5yu+2YntrurWf/krq2J1gKsjZtRCQIXRRG/jaXbblq+1ebyWj+
OHSGb+3gBb/ZSzZOrh/cbOgYXObysjzq3CcvBhQyPoDDoqUfTVy4Z1NGq0FUdzgH
mgv/tfHPwYA52wLN2OGrWyqbt96lEXpZNTN4deugLp2eih5B6Uc6jA81jdD3zNRB
4Oy0H1U/TiBOL2n26dCchyJ4O7rJKI5h7Lg52Q2FObzWzyM8TLxqtgH8ctFmSG7F
acsxnqp9MWZt/HLQdwX8nIq6LWR6JDm0xtHdvrEoKO0ZL+r59IvqO6V/pTPp6xca
Gey+/3CNimir3sAUzhbgNVXg+QRWEPItWfM55lfy8mr9m/kiogR9SLwC1qprNngx
uLQC/00myQ+E/uIV2KzEs+a6WGgtQhSpU7jJXJZ/hGDFHxnk5bxOn8ZyJRlF51RC
kzI6NHFyyp2321uWD2cvE0P5CDk/GbsfBQdxBHJNftJu3MN/T4aCPaLKbr/8U+uc
Muv16Ot9GM1o7zy9QCpK0CaDtn5VtBkQrbTHdR5GM4wC4+BNeh1NjYDXleYWD4W1
YSiQWBhHYzNWWQnk4Rw5hdNpEbU70HIrA8ySvhwrZJTGyP2lCq4JDJGKsY6r/7zo
gqicBeZlGz31f4jaCmlrqw25kdS8SvYLMAFUeGMTOw9ZDR4fbKS4hFWHHm0w4c1k
rHv3a9m8+pZYf/p2htqtr+rezFEHilb760fzxtnvGxsYX7pEGlx2LGdYczYE5868
bwxFbljfnG/KXZmPriKIPLIw4bhASRo/BH+7mcZ1HFEPyZ8pFq0dQxosjWq4rkKN
QTPfs6OgNCzXFTCjUNilNliYrKtIe435JDZk39hkLQa+EHAUPNR/I0dQsGwJxDET
63T4h/4geHIL7NPEvzMajLVCa8f6EgVtwp/Cp6zJCwmeIHs8tTSvYDr+tW5OObe7
NtCTvW+4Dt7QZgUN+Qi1m9Nkv+rkrGmvSwKXhzCZLS85CoKtE3TDMRi95PxFrYTN
z4nTc0rx18h2p1CoL3Ke3cdMGK5BUK4C3lhP5cpKrdip9D812Xzj6cAH7vwa6qro
RnoVF7UKtZCa2IBdbn0moAf40Rq84pYqqk9Z9rMBaxAnlfD4gZ9DakWfkcryVIjf
r9NU37XmVR4LX+X2MHlzH93cWIHOsb6KGHa5x4pJbpwAVuW2/vPJH6Y0rggkrcLt
YpSyVAt0ZSK2NPXQ05MCi/GGP4iWI5+sbeYIbf8jtsiHE6VKp9O2Ru5qvK5OKloi
Qf1yvU6iCJ3wPWNhKm9Z7l1PpXGfHUAOcZ3+ooiKb9pHbSc8yuM6TGzwOhOMt13h
zer9mBUnmOfGOrCa19lQSGwfT+jsRccwEj8p38Zm2nAAXJZOBD4MnAGrNbnJaOhQ
6wVOkySt0/DX2sj+V3jb7BbOoYnoxOWZmZMftkw5tgHiAE2dSUM6pTNYBrZzUabq
bOlITojmxnWr+j1jBCFxsHwE3GrmThXdvu8YUmBc/cfTbvpbQF1oQdsLTG6cfIk6
Q8GOvUm2Qs8AUwcuMkzv84xs4QOb4FZ9vCjlTgLMfmyhZDSZ+VKHXYIgh3Ll+wfn
6KdKcVPXYd0pnx1XjRpUoOv9trQD6pRi5w+avhDThu/BVDVZRcI6lkv6x2fTqvf0
jrOic9H5oIE3VBUuTlzrJdLlMw7Z0bz6jGF43aWC/Kiy4tado6Q61O3wOVlvYBVM
2JrbuhPdYZ/noxOXZBA1o1tfox5L6Ukt96ep4aNqakPQldL52XMeyaGzrtvUpAeW
gD/HCSvgs9QGjRgv7HhhywzgtsJO9eimywTNvi3Q1W8IXqynkG7VjEfCloPdQlSk
NOx6bEP7686sNjQbS3v8rYgbADu5z8Gc747UtcRs0J2J1WuAaMYq3x7Kyg0qRIne
+upMKH2x1ISKD76sCU35z2vrExRzDbi07b69mHjQ2jXMJGLuxoYyy7RMEmswX1+u
KBCBQDgS0Uwnudb/Iakz3oqYdUkLw88X8aTvkX1LJX28BtB0sFLUs387IhbIjo/J
yNQHiLqlP68ptYqvIFahn6uCCwbBu3N2bDUEFgD+K9HkaMKsZD0h3fO0oQbtjhvW
E0DLSH0EI0Snc/oA+atKvARc1+mLqLM46L0d5PXX2AlgCg8okVpwqHkPTe/eHfDa
awoRfTCPvA5cmMtAOkbGHPjm+i1Ru/SAhHkRrIkUK/HdRVkp2ecLS7qXDwSfefjw
6VdrYl4hAW6EjveG6VO8ZHeCRKRlbDZYu1XioQQx+MGvdIK1BuuE5rF+Rhjw+cp7
9xAx8jJOuhlxUpoJkt7ttcFeHjUr0xgsSKjJQn2qDYoBPWH0Nu4hItvzR3ArS/i6
vgNllgj1Gp493nCuCPX/W5dPWl46ubqndOPPzo14om0PZEDmFmeVsmlRHEFssvYa
w2I8oii9mn905D/S2yqAPuHnA6HdGIx+TyWJGdCK22JkOVpHXEwN2bMpd+g9qAl6
WporYafZR344qBMi5qfbt0L8ysCT+yfS/sWbR62O185ZshJSyHjku4e20QCv6KVJ
2Ef4PZr3YwjmGa5jm+XdraD05erGtU6IjpPRN9SvEzzoPxdmCj5q3InQfWIjClfL
SeyNX4AEqqtPTvKjITQ79nF48YVk4xEPxgF+OCSoD8Yx+Cp+UWUbrgmiITeBlRME
OgaphXi/MJaGlSpo0R5hc6hvk3ihMrpKf4Ms7zF0qg8X7S+67NN5iOZSlCbCO+ao
zG3Hc1bmKLeJl9/pENdKqY/xoAX699rp5y7vqY2otNFg3stqQlb4ba18xZEvjX8x
e+1rka5VPzAu8Lj+OWwG2EdHae6SYwj+klLVU7j6NZZ46giKgrWlqUntK2nKfLSu
hdrPsp43OlCCTSYGJcsrSaQp5/ftyT/4ZryuhLGRfSsycBJPWVZnK3t2hVUn+xqv
wgLfTnE6k/bGxJjDVGmTOH+b6ZEAFl+FGFtD7zkZ//VBa+VJ6JETWDFRlrEzeIwS
8thdbKIR1QrK1RifjFiPPFb7MGFy/9OicT7hjOhflARocaPWH88sfr30AhtudYR+
EHTa8/39L+SJGyykbRDY8rgDB+pPN4G0nL74xU0ngI4xiGjLg1LzWet6kgaGDe9q
Fy7J4HLet7VWep3q9ige1h4LBSKfcS8fJZPeSl5J7DCEbJa1MFBDOb5CvfIxqwTC
xXzjSCygYNCADEIfzlt9FY8y4WrDsXjBRfUPN7r8aYh9eew7aT35oBpske4wm9vZ
qvWJghskA+EGT1Hdc643ylJ7a2eFi/o3L1R/5PuMqbPnD+hw5ts0a+Wpt4SXTzS1
eUPvd7VYi8WpRW0dmPRmCUs/bAJ1qivuLLphXAgi85CdNB8r9mogj87copwfEIKH
+t2As7N9CDzNMi1xx9xDNUuI7sriTz0QD2NQzpxsGtShbHNvA3WYSVIgo5l9pvq1
biwExRKFJJQ54NPXmZ+0QGfwWt/1Icc8ZuvNM+6QIjJLeSS/gRwXUn4QSF5ZIEdS
cN/paiHl87MLcJIzW7c80muzAsfpHzfDJycA7qHmAkstdNrPooaBD10eWFZueGRm
d10lHL1IFJFx9fLFUMrClW//Ays2zDRBECCvheX5G40DcLCyjfZuyMqXO/CzqiA/
Ntnq471cLwAmZd0RUEVBdoIIoDglDYGzvCsRHESQuQk61ZUWFHs2fkaQgVXsF59A
y5PZ7Z5pPVa3JdKDdX0p25VYiTVFEelZA84uSRE33rek7duj1s2ZmffRQtUvXQwR
4EbFPeXR1ZjccahSNGeSAFFfGqTqU+OsHJ9LgT926xyGdGzMSQJU3Bl8fWfNZ/e8
Rt9ShsqG8+Yw1Dh0SrbJWr5GnkaJSi/MEJwFlVVRADNWQ3QuB0/tjbY6Q36S3dW4
JwbsBr+umlQYimwU3Clsc/0URbon3VBC5OnUT80N80I+p+1LaRfC9UZxly1kBaXY
UgatNnbkHM0HciwbeMYdyaDQ27lFabIPX56OlrydrYeWn7iRWav4VvYTrKfi8kKe
pTAXx7icrX7Xgzlgm/ON72aJuxSX322fJBwFEt9v8yoBy5As57+ZQOkw1ZrKDoXg
RWfi8wFMyw/9BhfNbwA/RLZcWswhx4Dy+qubIdoEm01YEtLXsNFw8piE9j6gfGF8
0E0xNelWlKDXO9giJbDdshvZAe34NrfTdziabp5zhDjz+XWHUPluCjblG1aDOor1
k54EbqxwmpzkNRzao9fiVb7JwpCyzmIwP1pqBBX1cI780V6DOlbsrsDHE3VSijxI
dVCMX5+/6/lil3Tdxw5zG0njyBp4lIjEu3YaRrjrY2uhBuKeFhos0OTfYP9d+F2N
bHirty3cGM9atg9y3/0/QNaMa5WUW679cgCW9BR4GNrBsQlRsWVr1HNz0179dn3u
9qtWIJKrD3BFMpJQDwqVMhCJ5FWijqcjxx0cJRMfKoK2spik2MV7eqVrwJE9h85n
n9df7+yaC3glhP4Jc2cjM2pYn/bSAxytXj98+WLPNT6PLNtV+NIiaAYfb3Es+BM1
A4/7X9P9MN2hR8tqxvu5PBN6ElPIJvzIn9V19WhBui85MyeHvDcqVEli6zMIb+N+
mJqoxwPCKqhOLIsopPs3nI3FNP8K+vgMxnM0N6n/UA6MHo2YXCE/hVZ0BcC0Goa+
d1zC9QZylY2azUOIktJe0y44TU6QigwFKdqk2yYbxk1MCBl2jZar18lsZJfPksAo
wRYcBMK6Ui6T5obDVf+FCvW7JQdOtOl6mSnIL8/17B2yab02DGW6+wISu/VJv98q
ehuo6AS9Jb39k9g3ZDwX0Y2Ri8gVpLBa8Q9XU6xUutuS/rBxhNGvb5ubIeRFTNc5
43qNr8czPP7trptADg1xe0vqWOaRFqaXBCI1aiivCQfgV4zVSoZetnn/Hv8CyScT
JryDWhgzln/oeM0Jw3nCwhFfem/VK1BskOKfpCNah9SMGl4jhPwYNR9Fxi/b03g3
BOfMSAnztYRIPt6qz/KJUYTCLGQaSmhJN1nqcHVUcVsj2/jdW/XSn1thxXRIM20c
aR33AVECr3GpYPiR8T5xc3uZfgozfbBOqEBHyEvpiTuZWRh+EjY5E0/JpcDEd4JU
Cek4TTxiDYN0ZOL9vpiCrPL0F+uIiAHxs5OVhFy31oQmMEUqQBH0xscmWr7WSUJj
aekCyefGoEIE/iXdrZhbRWCNifaDwoYCK7IJ2IcaK3+f9SmxnMKwJjwKZUnhmNXK
F2kbZqUX8gicIMTOhxsepearUnqdeyFkX+CSgTtxwUGgY4oipYoDZK/WFfrkkwE7
rqs0KwEF9VbaWbcMK/6Q4P6VSzlna8yqS9LIUN981N7HM8HhUST1HqzCZem/hQ66
J+LEkQGabULp85uP/4dIeZFMvqPe3THJJG5CwkoPuYj6e5J+CCMAy65ZblaXsYGX
OKm0gIit9bygxHOtCATDdu+ixmOhTiaKTowOmiQftdmz0GS5ZI1R2j40/dki60Ff
h5P1hAcUZNBUciuxjDezn0uaVGQXc3g2wiTykJmnVxqc8FOnME99zUzLzu6M54Oo
ELix0BfUFNVywYG9F8r8KrZmNbkaDHe2o7/yAcxpuQ/X+PEaPexYraWFpqdOL2MN
o+EFPweA5Q6dJiiX5YTlZPYHxVfHQC8pBSYt4eu9VIdboC+dkdKG0vytleNayMge
wdKiteeC3ZR2w5FSnQflN0ChHGJBQ2pItLk3hCnRSXpir9qlvghrqOtHxc41Dn/K
Pb0q0GOxA+vMPtnKxmZ83vop1UXcpT5E+26Ydmamu4gMLM00+287r8bedRXTzLyd
kuVgxnwyd4FzvO8uZ/ttS2CAtbkIAsHkq27yFnGWbtJeAH3Go0ctJRBqvipRxT/O
YbWShOgy4iGe0ki+Fkz70PLo778BOnB0PFML4PrnYisGBpaRxgkUI7fPDmizWvRC
MPwraQVpdvTLa8oECKqkwYX1FczqyipAiVR1J4VLKXSqCf98NTu5VivKHR2QMFLQ
kIXUowv/uzZbi8DGzBFxhVOnGWgo8hVy5PVd+wxBtAeb2F/DI8mPUIdqYqTjt+0Q
1JWfVXw+DcN8fkDMgWRohsl0gdW5X1fIXp3uBMHij9L4w+VZ4PShMtTSt078rVVr
NeEePu37jRXpKaQ3Nh3+Nw8GhlZcb/Vf2JoOYJ8JPM3MtgKQ+Ezxtlp9pMlEZ39R
smLdhDa0rJuBs+XnzhJr5zbXSQaKKshd2aLrVQTwD4oViGogdsTBA3Lk/z+vaMmS
e8PxXWOmCLSggVG/w083uaqRCJL8qg+KDkVQtWxsuIbLt++9Tcyc9uYdCDDDObRS
ZuYHC5GshRR+F9/jr5/ieMliGekqNvROCZNuqyoeTqPAJ9QLCjrZBmSaL/gAw8/v
KkmqFuO87C9sjwLCb8W/rtOevV8s4DsbSAs5agY0Qsf107tJ0tgnMeIHxMg5ctb7
u/4cisonHflC40Agm7HvugH9Ve4L4dTrOUI6/8IoXDQXOX/+CqkscOE29AaM54I0
54AvrH6UNnrwuMiRu5ResAfUMDbfyzPnhPS7Jh1FpfKrJ50VIdRd3HpE3A77uHHb
am8KgUqFD6ZG8uXrPlrllvISyhzro8u1PY50zU++kT1khNpnxUiPqMl6l+WPFeoV
w2a1+j6zo+vl+3dMP86nW4STh7a978hZQktR8vBadYUvYXnOgDWEI2ZjsWjc8ezZ
AHDoxE9RAt4eFi8RZIvOsrlINVK/FY742SvwgmJyiGkrK8i+l9mg9ncYsjUrY893
+hfk638pH34pVN7l9AX1j6hEm4KrF715rjeAAXZxqpI3piXPzwCRBC5iLsY9v4u1
13as/jqfIIVQyNJibt79Va1CykrgnqF58KIaHyyRHzANZ3XD99v4RX+rwQnBNvhR
1RhW1uJXILv5Yoh2pcaBEuOwnDMSpicqmT5Ia/SS7/jjKYQGfGqFNMsFij1RD8k5
Av3m4slcB28B8AwyM8AL1y67w/dyQZD4lPCMchDXugJquxJ9Kwg+dy/YUxUCzdD7
/0huXaySb+2RLRnpmw/5WLI5A5v2kadFR4e3qK2OVHLgCzbHTxBFjizckhfMS42C
GbPg2B3s3OYg14JAnEqX1htSNq/fV5sPgX+V2FHr3kha5bCrwOC76UUYRffP6MQ5
y80gAyP1gDcHuQADv41ChHiVVcBWzzwU7nGI/ZpLPaHgdDe18fmG7gHbthxqVIDL
u1LEeFpTRvPUZCyyo8x7U+Jv2Hshvhsf0Jt6L37umq5UPpsY7rn1bSQQusAimPGg
ZKC5k5iut5WC8OYQPO3w6LuKj+lN6pmfvsuQ8eri0wWRLMafn3xP+2BRUXAXtzyh
aO6iaDhExqIbT84owCED7WSza89ncUCot0ygN8jaK6uJyTBysrU5Xb0yTyBla0lQ
kPsyOQxfJyP0fi4oUvT2proAz0a7yGbE96NvEFHXRf/ee2wrdG1O5QgsAkAO0NsI
Eaz+0PZ9ZvjfUvgBBulsJs/TV3g186VCMjD5E2qmA6mfvuoEzpGQO8PCiDdzuPbQ
0S8rlc1qjH5vFSy+2Zt+ceUK6+jPpXmAfsB2DfYFjJLiLFPM4W9qUwhTX9NkJ0Jm
WX2gVkHXc6w1lviKQgm8jRt9Rr9kzoMxmqfWxFqAOX/U8LIsaYv2y8U9w3uDIfkq
85v+ADJRT/8mMJZgTjhr6R9MRsfChdWeey23DWSporg8DqkqXSaypoaD8c30aTX5
M3yDa8U3OD8s7CjNZYbmBCxwrEJDhoIpttexiWzt04Bo2Uh36WoJa4YhieT+FVev
kfgXBRYYfSSLHVFsgnA8zAshJQjNNUBZpcSwjp8+twv1x203M4MMHOQAdTySNK2b
7e+59fhRhyd35EWGcuszAN19XFBiUytJXwK0x96brQqTNLi+qBmpt6XaVs/vXNvh
ygj6SmmVY8hU9ZGlj/rty+81vI4jwkEW6/trakhETp85ryaghFTz78o9HQ7Lgew+
VKQVNstQaK0EsyBWfzSOzVBRMjFgCRNgNxv0z7PiKTnzqi8/v4ndCq/NiQpcoKhN
eN44ttBfwMVvvuF4yF8DAv5JBOr1nsjXSsUhmkV0C1Jcg+abmKbCLD9qBAOeCrmx
8AN/Nia3f7oXc1fBRPhkOzejGe5Ju9gR51F6xDILU878bZasxRA6gfgeN7RoUWVl
6i889ViR5hvMO0SDG6ynxMPrr6pA7dD8cGZ+ZcRQMctHUA1JmNLwr3PiViWXytpi
g0PlNOjwfbFFgALrbCfXIvhdk7Sa3/vY/2bi1Oq6joJdsGzbRVivYpuUOurRhCQu
HsuTFOxLkntWfPv0dw9C8fpncQCbgy9Pma7TlhSCvVH5jxyBbquqCV/yIJAgTaS5
Q4NkEfmilfwKfWywC88wppkZTLNoEWX5716hny6I+OGNY27aj9SUJSeU1j4PaxQ7
nC74deBl1CnEgNPNNBsImwz6xvOJhKO1NBCuN1B2xb9CxLgY7RrRNBcmb4rzkTnE
9XgkxpaVQHxdnJ/tpEN7TnXQei9dfqUmBz6CP0t/nB3FFuxn2IDDfqeHxjjCSj2g
AAae0S98sup/jtbi3VuyE4S7wgjpGXFECQwbQbZndpCjWImwaFoZp73fV2EoQUhQ
gu2ESGW3uXchPxhx00J3wJDLx6WzFp5NeKiU+dXjnSTatDC0vBdOlkdAD9XTVa9J
1yz/6NqWUjSRtUMVpBS0G4wzqkyIwUsoP30+/9el3vRG8IOacC3+Bglz/80OV65U
iNB5p3USPwzsoVrVGILn9FttLrkcFb8eveprTNUGS7Yfs+BeTbGkn99RWmYwc07r
WP43A/LRhmHFLezHTeHX3K+gMhXTS0o52lcY7uAe5qGyxH4qXzQ64GSM52HWJu6l
CmsIX0l96mDbtWCxP4YLoqjY997mNfpvozLctzbNHVMpjU+2mhcjEhAaEFfeZ+Ws
i8Gqqn7SzLxepKUWPSONb0lA8O6GQEJ5JziCJkmKAJtL+0fz2N2Es0LT+1Y96JFY
wplkcTifTl/NFkkbGcaDZlV49O6M9N8IbMjr0M358+vcUiHWSLdSq6TOXx6+ypf4
lH9gH9ituh+VW4pQQUsjIBO9w11WpYtIcqrFcANJGL8FF+VA5uVYvI3RYgOBFWLF
M1q9YN80zKmKW9V1WpuMMPdohMrKCWHZbJUECDdCf04FsdIAXsC8D9eMid/DoF4a
pWXy1KmLfzeGIbFwF02hSY97qILP4cG4nS2negel9e3cYkfifVvvTdR7NzBKXOI3
AATtKzQNOTP+BBtFmZEcK9ftG+p8nJ2PWBtx0iVGh/wetF2NHb5RPa/ujNOqRivB
8bwFolHCbONTZ44PLV8psCxtdZPUPAe/fJfOwgdRp79xxH6fi82yxPj7txTdhZRk
ex3Ac7Ra+QFFVfswGU9sWELPNceXV3lYEn41jlgQSQT9fjmn6brCsYyDfpWFpIDG
5ayuNbLur4euNuHY9Tg/ypyWxuImGHA1CGpX9vPWtEHOwloIZP+3HrYg5PEjGvMA
pgOLqv9IjPr92WVPoseKFFbu6Uu0/Fh6kQVVhPfHi2yAGiExZmNPOjg3oiziYN7k
+UXkojEz1lFEpJg7hKBpxJ5gzda9yhkeT4/vcf/E5TFKUMSlcqh6Wu3+O9/uMLbQ
GdR3Gb4SRsMAEewS2jrO0q5tdm0RAuRt3Xn6dtstaRAara0uHUFFnOJ1rVhLrJxr
Gl/lvbtKoy2OtrM3yCbBarytF9/gI88kDD2dUODatMRqYp9iiIONbKqG6nIayKCZ
FA87rIzXBiFXzw18BSWMtJ9C5Ysin8KUT8t7mvCz3bGmF2Bb3fVEg//V3Mci+Ujt
zfzpoay3wU16dwK46s6loIPcbT/mIuq4tGIghgvQHBJdzdOCqBfomCaiOLntv7JX
LrG+CZCxVUkOTVr0oejt9f0OKc84fzhmR57/2wtWeUiCnl/TvHDyVD99y6afQV++
qSHo1btMQ37enx14VfnMEzK8nptiC6MznJsOq98oVXAXA0Pfoc/Q3OSFcerd8pdg
VJJmM3xMaT4AxGPeU268WccA6tIagySoMlOaOd11AeV27CK9F5hdxsW4Mlsawbpv
Kz8qMrDKO5sJsKek57LIek5n6M0uPClV4MxplhITG1BmBC7FhcSenSMQhUxr5Kor
2jREQO3FCEKwqMBd8nizWTQcIul3M/xqFYXYwo7iGcGkHHxyODLzPbQBNf7wLlS5
TZymbl4cXRYnI7Xj8NkWeRRT/SZOyPbwt6MO9l62BHsRS1YZfiJ0ILzz0INzbgyJ
PK6B1Xz1oR7c2aT/Eoo9WgPRAF8Zws8JvrBzr13rE1iAWjeM239gQatzw5wFgOgh
a/Ta8nmRdsMD7j4vvXiXEz3OfE8IcH4yijpBOF3eLCQV2aH3QUuCq5Cl28JkweRj
IuUV6SflFo2M+k81GfbYWM4x60Ok973ikjSSkSsDFRlwL/z2agPbM3F5BXfvox0M
zpCPuTb4ECu8b3fZvcBQ8W/vIXGGyYw9Q7JuKL60/B1F37Oz0T+5oJzyHxJjV5jj
T+QP2RspXCXh69kkMYuF1X/Yxr27JriDIQtevWLMGIBm1DPmvdhz/raEQf052ln5
BTF9saJGQOTunnmebtN7RGbkgNl5NV37ThWQjEZ+RUHadAj4wBjrMEMxgLZysjs7
svjf6sqatyBpcvw7qSxOsKGoKSirixcP/dgeZlW4ZqarjPDrwHKcDE4afjp54Zx+
EsZVJbqXXSLCai7gpUdUIT5VJQ/gLlyqvwIg1iyAJ+asDOSDtiN6YSSJ1AI+KRlw
+iNoLy+Ma7tC2nSLzWaNJJx96PxJzRkeCd/1m2W+8WMqiZe74QukCImOGW/PAum2
mUK1rzC6wnn67c7PI3HdqKRuFKVgpRABvKNBpw2Ua+AsP5po7LHu6BJecT4mOG/Y
yF9K/axhfckBBzD9N6s4MiMXRR+Y6TAsiZfthYXzajwClzRJuZtTHTBfIn4H9GMr
R9sUChjmUj/Q7QPs+IHE8w/ltcVX7sHOZBZuD1nvgtE8LgWkLtBIF+MQB5Htxyj6
qRTH8cF/q1doonTFB8SOf2S3hIZbFdhF96kKfB2h2VWOv0fUHdmwrZ7P4qcfMQiH
XQr0KSS0m+BQohpMGNKFy3h6E9hBerhC5HjIVzwhVVnykLKSXYfEmtKEIi4/t/NM
kpWyD75e400l0EjZPAiJAzQfhzNe/cVHiyBQTi8pgkBpzcJf9oXdm7AE+cv4J8he
HNAs3j5v+Eu14ObTall7MV4i1nCVxwnBZ6ckQzNtvm6gz4NRQkjCMZHVusdzhTvk
ZBRjAXg2E5hZGFEh0J4nR/htk+CWJeh8JEOncETl51Y5LvhDyquj3eIMVSLY9K74
Ks3bRlKfLjo0M+bcQWT7eBABoYCKgtlXPVqojle+sb/8YBu4OANV1wsPkTUK4JdK
yPrUDCAOzsq7m6BhJUCN7LT3MGHhEEKuye9TRE909vl88d+y+3L/VaGPBLeaph08
wILTkza52XdAn2e/T8O6UIKHo05lPAXGe5L9VYmkmwtm2yYpNDb04Fu/+Jj1mahB
BQ8BBanXdRV+6jSJbrxjq2rebjbQw3fs9nT+SA18KS0diPZq+yozGmEG+striiV5
Fh8cY3fwOR4IR6zCGsSKdjS3d8Rie1kfslspabnKHHUV6KAOaGiATWMCbtYhBeJO
CQscBIPtLNKa3A6GVjg9XugnrNPsvZgELpc7xKdsRg8CcmTxBySxNe6u8jEjsmoN
AEpny34JPfQJOgeD+HRG4qq8Ex/aT9DzQdUEqnb6gdJ1XS8hau6AcqpC7wh/G0ST
B0UlPrxdtrsPP+0RiWJn7gQWys23FznzO4Yf33Z5nu05UTshHtV2Aab5RUvKBxv0
4s4tM2wOm1M8Qv6gHOK/32SRI66d3ntxBXdzSCqtlkIhBUgF5rVKIsSotAvRxzZ7
mp1P9Y5krlBM2fIqqg1REl1ZzZtw7pEW6OvY4aV6DiuZH95j6r4odRzZf7ImnhMZ
a6p8nP64flITT3UAiojXECMoqSJbdeYSnREQtD3aSu9SdSx+lwNoXtuQyJtf1eu6
89/beor08XX4g6KWYSFKS0TOquh1RtmFg6XM5F/IgH13ZbMxJQZenEdvdeHq461i
qD9jWqQ+Et+DGaYz7yAdMmSSixVxgXgbkyfnsSHeWspfygxqw7FAS4HwvShQMC/X
k20vSMElDq1HFpelM9cLjGaqFR6cl70ZJv1aa6AvzKK05LLiThLUZblg+HxE4bT9
siAYLWRsmTuweu7f599uxL71E+ryrc+2D91qUE9oRq9EzIDXE2Q+oBpAe7U/zz/E
t5sjG5puNbJ6iBE3pMHJn41aI7oCHIg1uyKdHT3K3e+CCKsG6U4Cp9vbK5dr66H5
LWpa4nfVFj2KH85exlz9aWbp7USJv8NNC/vYzzA+80zmcVBguUuhv5lnaFUmZ+q9
BT5pCN6tQHVeZN3KJTvQpmLys4dVyd3wskwtlqxLSOwiIzx1rJz7KTNxf4XO3OBD
ZWUy9LNUv0pvFPnHqdZu4sWFxo3v5CWIYzYowGor3wJE4O49CSxpvpM0TlQbLaFL
RXNs3b7z5CZk2klTOXJd6eE1NXE29hb6tScNIStRMnvnHzIQA/u7YGGD+Bl0cTGr
NCC63AFDxIiHEqtixhqHPfZ6jaXWEIy8ed0IdirH1Vq1DLoIbRSwO1f7+gp488fq
fX+TT7NvA5NbR+pL3z6lxl+NR+hcCy70bHyF0N8/wKFZsSMfRA7M512oNvtMQXmv
F/aIi2oi5Hz8bUod4JkOZsZTo0Tc999FhLSiO5kO3AQC8kybctX0joogqKyvxphD
uMks5y2lu07UC1vwleHHFZa92xrqNUFxn1oxZ2Sqr3whGD1pIW4sHIMdUQbcNDMy
/3eNL23/3JaPQXVcaDR8L2C1YFez4Fh8qLUqTvdLM1oP4wwyacDNk/iKtGVCP1gY
9D9I5/18i24CBYB3YAWAVlZUHm7hWMIqo45JJZGT2N68wYZuACA2UuXem23R9ouL
tWRJ/J7c19DTfFveFOYcBc7Qbs85xdfnVMH9DOPBuT6hbc887Fhc1sVUYV43FLpg
mR5H7sr/M1JLzlLyRo6u4ltq4mz8Wfu6buECVAFCjq51Gw553Oo3bafgQCf2wHtO
Kx23g0G2iDIXdkPIsoMh1fAAY03gff1Heae9V1PnE8H2HhSMwOhup+Uv8KQtUwk3
3fwhrT+4CRsuSLhpp0MYxV5YaS7rEh/9y+S0v3xIJcbJG5LrNQvIbmw9+9IDsbkX
edM6Jg+f5U2evqjSk0X+HSv3Pbw8s8XLgVlCY4ZEGUiitT4WAnaVWCxbn9qdNXhM
sEG2oLQB0eoyw4HsvutcDAVDBWh2WKxzOP+PsghEtLTU10CbUip8Lq78vlG2qwN5
FeFZpn1JmtOdWDCNsydA3HdOhv2Z/BQJuVZ2HBrnkkVJfkCO+Jt0XVMpnGUtrbvU
JN8Zh7bLBXcSbMeqQMBo34+2TZMqHNW3m7dsiVEjmLHtD1amghQgiNkBbxCXpk2U
I5ofnrDK7ZDqH4cWxv7K+6wfhvEKPBnwFV7ea55LXvZ03iUKpEoH6xkgVSCxQaX5
OllYDYXiW59sol1dMZmE4WwJtsH5C/JTJq9dcnWYNMH1kDISMKcaPntvyrPdHHGW
4hiTpmKdBsYESgOunQmTLlwFAOiZjvytQ8HFeQdAYUca6/DOL6eq44n/57azseG2
u+GS0l66aSWp0E3dJM5/+e5PRnPItyuaN+hCmaaUtW7rsftCcJjWoxgsQfGZ5DGe
2DjuaKLDd8VVjcCnxIrXLXjoJ3wEr4hbvF0svMk7yKSYCnd9rBUMTJRXStw9m8W5
+nAHImpNDnnCw98kH2piNTPSk8XRm6vyINC83yKvMQeaPK+/LEhaf2ofZWERu1ib
vo3qmlI/o4HmUU7blxk5ga64UYRrlGbAdwLmTeXckjbeLiITN6CQFFGu7uOV8lGt
23Pg3p5O+iW2xVS8f/jhddhiI/uAjghPwA0Nhs462/wGpE28J9LSNnE/DmC0jg4V
jRk5ZhMM9wG7YhqQumWmbCylV7Fj1HHLXB+6yekM1KRRhewyl+d8P3TgIK/Pk7gl
z8aE7N4tDmvGcvu/dcVq8NomHodSRiWg5b09TJ5EVoO2qL1Ypgf1f9t0X6fp0dAq
Ev8nAMWmxklEe97OkC6KHo4C1ja8pfExMrM3b3XrmnxUafnNUn2g3R8b40J4CXyQ
sGQxQnJ212M+kFRPIbepQZBP79ab0boWJDWponchZJ9oR1MuhoOWKB3uxGIojf6G
OJvydOzGy7Pp5Q/brWtwIO0wAC6dvY9pGj028HbVF/3DuC3vLF4pJvNNYXBrnnPk
QcG1o1BJQMx3r71X4sXAZ6Rb8HK6jDq7gfpkGeP5YPG//xPVrxX+6IoC28NCmNnH
F1t+tnbiBFrjWVGf78XYRjubdRjePkyoUn+b90dNZRy0JjQBQrYpqM//FJ3SbBLL
KN3utLjNxo8ZiXqwhRaQkbQl83mWjxY6rbhJpxuiYImJlEZ82x+bJGKcOLXcFZw/
/jdHxAjVyELcQ3maENsg1sRNQwCYSt5qe8RCifSFXHe6mIEJjXGImEhABbtQofkL
nzbc0ggO5uNS/Pa/fM1am0xx0PVb1l/TkFeW1BHf3JHyHMGw/SccInQv3Vj3mNaJ
a9MYNd5jNKF6vSTwZU/g04AVpnqoopMfg6TYDAx4NWLP8AYe4EaQW06ZR4o0OB3H
lYX8Tcrl7qNHMMRsZ9rlN0j8QOYMfeKqEaq6pSkn7BXMrLx8baqGeOC4h6m+kIcr
59xoL6zfyV2I+Hqo6Tb1USfRIsv9dhXFHqOWdtI2PLh8OIOZPepVoBW/00S3hm7d
L5K6S44ydqy6t6wE6EfI4XzTRAmnmcGbRJR0r2peBulx7hkdPWXGZl/pgoiwnNb1
YPnZH7KOCP55H7w9e7hF7LqOTeDnXe2uuRdSYzl9X5n6X+UAuaZRBBIoUplEOncX
pumrZ/aQ0F8ExZwjNaMlcq2QGJ8JEbaupMTXecPtkN5EzYWgBX9+4UdqXwpNdwkR
7k21sQKWqhR05auPzKYkg2vs0Jmsu1SsdZ/isD3SXcjY7FhNqqW9AUZ8z4225GWS
vmHwMea/DkVW6vcCO1BESJ8g7+Q2+czHRB39zpt3Q5q2K7FC0VRX3i1uL9zrSPbX
EBqBA2W5dPAr214eESGowEKJt2WSpCJ0Ox0DbPOhjQDQ5vmM+P37Xd9o6iEvA9Gj
7yHEoJl4bZY9H78KEKeInKDhVgN2GJlPTopAUaoW6NGL/s2AF4Gx1rPnmczq8p35
W45q995t1ho6LNpspmsbCK9icAsPWMjmNiucShrvIDKAcI+/eBV4cVZ5MUy96kKD
vNNZ+HhU9i1DzltneyZDjbc70UA8arKbIspp9RJQ2jE+kLaGfHccKHxiN+S9JHIG
88cjTMJit9Xs2WymiEIsoB+H4YIKN+0Vii2eS3BStWlR/cT9EXrGe5i6BhFL4LCY
QXG5gv4lUxe6d6OUOm90Bezix37txgZSxuW0RPnsngShcJGFz+hN+GSWdnLBQ2+D
3KZf+Y00b3tmZDtvtUndXUUw/DABuMiNY16t/7vl2dJ7cxIyJN2XGKqvZLxHLbCv
bdeqlaT+LeQepQLw+iEFHGAebaI8cPY12kBpRCVcNKnAx4W52VfmxPKOyKzyaf3u
hmrCeK6sOm+JpIRPQM4VY1P5DztziT+BqorLx0FXXfJcQqwv61t1Y1iZl3VpbXF5
QXY6dTyMXvRbeZhk+w4940IuVt7Fq+puxu8hrdDYGcTvf06XuYWkTwecOlT112JH
yuc3pOd1DxteZf/WucCjXGduel5XfB5NLv8gXYam6ghriAjE+ExTd8sJL205FPlT
G2zClAflw92jkU3NRxZy8wCeBax2RdhoauDt7PS4nGohjxlhqLh77Yv1JBG655DA
xo4+1AyXq8vGcVNAYzq52t1VHE4p/pux0YSTWNmH3FY+nx5dO0iuP9iXTv9CQaEw
lLdSBRvOJNKLTQsHv4E9jLcsQn4n2IHxPp5evCJifUZExz2zyz4pZZgWLf8ZTz1s
NRovpILQO8RmEkUZ3ru7SroxsAyW+/DSm6u+f5VhTWTHMXRcZ18SKLzVlILl8YnK
9rkS3c9X5RQNzzXngmzk9MeeDty9nFxvwMFSkRB4QMx/DZkEPjK7atjAZXthLS+t
4AGML8SCU1ww1Wp3gfmsY6GdAIZA1ASTh6Ky53wkk5w0PNfu70K630glKfTKyu2w
jAVM1fA2tzEZHaisIntiqQYdq1e6qtdFINahz8X7y+nxLg0E3Aglk7nJJ3I+JLZO
vcySfUggltMGjD6BB4sKX4xKX2DikEf4KkX14XXwKT7FKTVYbTDbP4gN4A1rNx1I
jwmr9xI/NBTScPi/nrbSUXQgj1TAr9a7+PdHl7ScAKk6Sufutbpx94qkmfShdCQ9
20IUpxfq+3RfiVtHFgaPfNUWCpy4xcdEO1KOgmW+ZXhhmiRCCPXAr8dm1DMgxbT8
IxkjhX2var4cmMR9RXAZFzIK/2T2lmluT4JrFk/1p7lABMhwNPXd4cARA/kffvsn
ojfxdCpxboKL0XGBIqp9UhXnKarfNX7EacxwuJbD4uhXzW2bnL6c4k1az2psm3xI
EQBmXMJIfvmFRCF6g4B7U9BM9rKhakG4pAm+fCvAIuvsO7B8gN6ZUCIE4VGYdH8J
0SSDGMFi/fuDbc7vVz4XsHsmE+R5RtMc1yTb+XG8G9kqAkMOOgBORBrs35k2RhIS
h2KzoD1xLxNRpXJbkeFMZFS4gWja3fPEJ5UrJjS2RH0ziPqM6M2G4rNOiNDOlP4D
CvXUhSYYd9sgEIMzNeyUOXGTtOrRygScr3LZMA6eXFSUfx3PpNyXYHMmKBgS4sau
2MCjDk5bifPwjaWmdpNQNWYQfnkjW/ZzrpihprZTCHxmyc2klCz4tZpJdes9Dh5g
wlUod2GLGqpq4v290TTBRhLlj7hZFJMfpLJTYaO2WA0gz2JoOWDJySY1K7VkZX+A
dDwjDDSzZm9pMc25TwKiadelCsxW5ByUT31hlxBSXvyvwZawtBnizxazoSj6J5Ri
x7oAA3wOD02/886mLmDKzCtdpOt2A3IsAjubFgPB4EoHAzn4CyJeapdR/uwLYt3N
4a7rCvJ5e+AFwxfWcM/dIQZJc/xXixHXNLrKD/omzQqyfFUVOA9VUF1EhIRYr1OD
FLvpmU4T2PCGwubTZ9OKFWKpatfAmQ2CKaCCSq6HwtrYahhV+7e26bvomE1rFEIt
QNAgGSGjlbM9li6rQmzovwT4xvls5C2eSJjgtRtC36xEG08LvJHDXHaHEVLN5y9f
Q/lFtUjrjdwUBGqoPUwpB/nIqYBNP6j4yVrC2Burhb3ddTQz2TTvAYn3ZjEFrb8N
Gij+2oD1YEqp0GeYA+QmQNZQKpVb1L1xQWQjuSsfyNOicGh5JfUI4FLTZ4Wj3dwa
sdudlXDR5/yM6VA2xOyVDQjYsky7S8MU8FyhHXAnZY5bCKG5Pv8sXiTiHM53FVdl
I2TMl20kj8PXd/6Bvsr76zryWeeyDqLWg6bgBrYDqLJF+5LpOd9hQ+4ByNH6Yrud
IRm4M2xXvJBe/SYOnmUlM3JqeRFfayOBK2PEroCHIbG+myZK9uf4pPZtcPRttLyY
AYQWfqIBwjJbf6PoAvdybbsWbAjRgpmwBnL2NYvXpJ2VHS+lH+IXYEur57lUnA/A
B9xMPG7Wmy0VScT8fUqtsGLo3IyknZUZNgRpNOLLdCgX42Q0BQHptfz6eCkMAx5I
kKMjKAqL/97sN0V8BwRELKq3lGCZbYM4ch8dsNDKwnOZXaLU7X9XczuKZHlZCmja
nGIgKABrod/XhBRmQp8aI1X3WUAqnf6YymODfCc5XkCo3Dnv6zKvc3rvm8GZ18VW
pDhgLeXbZUmDuoUz4Di8syNILIHhMs+oXVtiPwB50bygZIHDyYAz1wlc84wuylF/
fNxGgcJSwkfrEN9d0i5GsgqSZg33hDDh48KHf8tRQlM7vTc1/YdWrJ6mCKdBbX4f
3ePg1Bz/S8frsofSm/irMzHpuGxZinOvYwr9m6tsL14PvCsLrJQPpwgxuAzvYBus
oq0BQkc6nyROwEfaYqmwj46jCSKhXc38jIAP89NR/OkfAMh/kAgMINnfjZFneHYg
UjJTQwX16l2zyrWZ4OXZcv7kxXacSqK2OxQSUQndZoUXkc3kK8RgGIZCNZoZ27yg
b9nscosPPRgP9sgvdFp1/+vS1ybj9N2cYpao5BpZehyHE+YbckO/HF6FqRGkPzHY
NdHKuJxbR4272HrI+xCjcUovyQJtXEisLQRG3u1kTcBmsJDlfBNlbUVU0sKZXAmr
6v8imq7C+1ZWTMKQIUCkFWKHAKW4UzZOEzA0OoyIq3qkYQeX8OdkVSADsotydbmY
X+LovzAU9H0gFlcNTCakd7ZmT8U9v1TR22xqejOV8fgfygZzcM0SdIm4JRhhuDt9
YkTP8zlBkwenNfOmrFADGWgpZ+IA5O1FnEzE5nGTQpwKOo64mvGvv3bJKZpzBTFo
dk1PLd8zxV/edK456kDY+5Omszw+Z3NiD04hBcrySIpyjMHuS4wJChAUpLYmyg36
VMdYw89sYYPIUmO0K9w5w8cAx2fgePsn7tB78e1zDy0jV1egtAIW14kYvRgZX8sN
qKpwRc54K9YWQApYeYBC+8gc6Ow6ywf22kGrXCkicXaajs4GxN97IACbgKA8kMGF
yBCp5qNek0TtP947QGw/a/SV4VtpmvYLCxD2f75BDa9Ht7LOQhMDu8i6LOwq4uKZ
SfeOAOrZgyg8JmjguDrBa3OC3KEtRJNWeCCyjz0pO2VMdOKZvnB76Tmopf9W6p29
eyqe6tMopdezDjkjDPbQQs+8lI6S9Aq21h0Q52WuZPT44MphKerLPepO949qDYgk
gR6JAZhPWcuswia5+PSfxoRSEyre5nsmM1CsRDIfNjPGzHjB8KhHMJ1VIquoWNSN
XtqAsYEjB8VUILKriEn5SZv6+HLXHaLTdlxd68/j4B8dC348838FepkH4U89Izu/
Dz8o6MGT4Us4XJ42Egr955cD7uMo4ifs26tomiaUMD4X/7bBfX/aDAdYU6mWGiQ3
KnCXR7GxIDj8TfxVTiQwaNx1mEQ68h3Z6mxPvcg95v7jLdJg3swXCnmpVXdtJ56w
mVKM/ybFiqSYoordwl/sXCDYWTav3YPrLlWVAqa7uh5YOd0oNckKuU3Pwpm4hROD
1mqzxFkWVb9VISos7yVmyMG7c3yO2qAXrweeefZbqBqepazbt/D86QfwtN5yvA7u
NmEo8lsOS4c7x8gy1r0/vQdbya/v7QqeUcMG71c7tRq5QZjRUAAXFmjq67XJDKFT
aqeLfPUMgIeK5sZs9knAKqtafdiN7rEsg5kxfXTGblZIiNIT3UvZUQlD/QxvSKfk
804Ff8GEjNP1SHOExrXxFGLu/2WnnYUZUg4BZA2KM55PXL+cuwQBvV5F9YHvB6oE
lT+MtIBSN9QjhSY/88yaEugVRWq5DHIoxwZs/fut4wa2jrl1B/AO3pt0tNIQKRUe
B0n1VzWspp+aQ3zNbWsedEgZEbeZSYLnxxJUCXzxy/WbCZcoYAQMjznVH2XwXFC8
vqGgrsU24mzBJnAnozL3yswLTcu3fBGG9uMLYT8yVta1m400oei4l8n75eV5C6eZ
akbENNOCxOG9MPTKKiajmQp0oUxTHYsXgros/BcboFNunJWnqQxWjRkffAr+mZ7j
W+1+Q6Is1pWJs9rflK1aDWz81LQJyFuMZGFqMDN4G5z6+2xib7oDy8RhBimvXe33
sb5TnaOh1RFSV6UiiDpPLW+fLGgk0HJaxDdcch4rrsEci1LXPKyZshsVHiuyKw64
AaNpbsOCNrrrbdqdj9Vdq0YVmJqZlj3CG+JGgPjB+SUaqmANg8TOfHGRXNiMu3w2
bB9s6rB+4l+Xc+4JhubpBaaSGX5ul4tXLpP2bYgBIHD2WL4NusKt8IZ+CBvoFr1q
9TO+7GVqFx7t5ZSpO3FxlIXRYKZaQnqLCzMHKHrViuMjLDzyaMse+8uQfRg5GGMG
Mvmh7DrvsN/kvs1tpij07oeoXQyH5cBPA3bLJoFh2zzbV1fRF2cxluSh9tGMsRR9
Ru8jO4Zqf1O3IUOf16AuWV/lHGbPWZjmjugb84IpOWhVoS5Jfw9mhBOQ54iA7j8z
XP3ZLnC9G/NwdlemYYq9kDru9Ibr44U1//5Xw0l7lSGFcgxNXUvqIsY8AViCFUHW
cS1JIC9E3eC3X7RLOo8wTmPRi9SFfehtcGCAlveRceSPGx6L0lgpqN2xmrLIcEB7
ID4gxANGzDGnHlCGT6v5LkITFreetz7uUBp/H7hZdc91TAh21E5HQVnnUAq1YeLS
sPhgjZ9oj8mfxhWLk/JGUWw4atMAL+LCEo5I41rT39KAsYi6SSDZ8wqsZOUeG96p
frAMBxBYnh+pdmya2Qx8mU0AlFqq81SXJNrly0A0NvUl9hcPqbzVPJ4hFKl41mIN
fj4kbm8vkQdy240LHcVEdmT+94Lrgd6ndjIRikuWuhKRMLe6Ea8CNCyza0gi+Rgw
OeNEBJVAzX6zWz5RD9qrDKTDkEFfVPI01uU16L47pb0ntN5rcR0drcjDBran0rW2
yaWScJlunp4VLZ1kluXpjQRUBe6L3ZgN1ZJCP6ubYjfdmCc/wdjCIBJ+kFnwDZqk
d0Y6BUuDOuhi/U1jYzur/eMdLNW31MOH2MjEUa/bAJXa+KTM9Fqhv7o2mkpp3SId
iaajifM0k3h3fZzNECbuhbajGmUnJhxXny36u7PL89ulfGBwDbykJqUyIQIm/ng7
M9SPmGX5g0m6dAHe/9QwTBZC4HpkthWD7Bz98zHD5RdDmeEtJY/qOxfsruNgX/TP
2/5V5vRPPXuHXbbmTbFjSX0M8ye3jfEupJDb9eNHvfCmGd0jVLI92TrkeArBLg20
5sAj+raI+Ztr1K0zN1PlWGYZrE6L+NT9HoK2xZF9O3o9P76gIubt2kjLKcgnT0yB
rn6bHEEkKMwSJ1zJ/hc+gRMiW2P8cUIHVq7aE8+/U6mFy3egp353YIxkiAOPLwJo
eeb6J3PKAuoL12mX91p4yPaefeL0omV3LDMuoFn4StF7vHQ0aKPLszRAXum5PWFK
cFP+dW0BlNnHzPuXucOlXKs2jt1RT0tKrgCB6gd5JFjVVLNyga5YhiacanYhqvte
4hIyOtUq7jxG3DQmfSYYypDaEsVkEi+/K/Rdq9MlN37wtvS3jKR8831r5tE7ygyV
Un6ThLvBtMENw2stY3QRX/yLpnWlMXaSwF68v06+BKxaD/QrJaxnMnIgdiou0hu8
6cgLZ14sEUjmlAIPlDUR6ouP0efJ8hFFM/4uIU4+0oa1rHIfn257gMRproBAzd43
IZyCZzmxNIvyH8EPX9z15IcApOkv6LXMgwABF9Q3Kme8g6x9s4eGZZi/q6GeLqsj
zO3aIfpop1LPB1k+E79I/UdctQ43DMLH/S9axJRVlPLEYjp1kyw3UFX2L+wMASNJ
wzzvjNDyseiiQuqNzPwdodRb2dWIsiT2FuFrw9Fq8vU+Q01c970K9L/PFLqP1MoV
Y8a412jixbOHtSd0uFTfpUfuWLvFLqNL3WNgLRn7xOXJvC59PyYx7wP3hizFm44k
8+DILcxATZoVsSg5OaYHPOgw0oaZuR3csRMVQQkAYV98raWM/ZP1QuwNIR/c4NZz
63hJSy3lFkfSxr0VEWnxi6H1acgwYnkEgHE+YK7p8CAFmQmgc8IxpmxtYd74rJkE
aWWg/NXmlu/b4MJI03aI7Me8IjepT0YoEWnrtqEtoGC3j3xBaiJx6Cmc14CTps98
+Wf2mKPXdzU5u/JkipnCyXhXETjDb/9Fe/lapDUtV8+UCbmzxK2Xuj5ql0kJ45m3
qhbDFyzV+CJWjxdOcxkapxHAl+ICFTMfbQjKKYsPwlAlohdXqnBPcb6DiySbb5HJ
8kUWcxiig3PkHVyKxeAnM875N69hamKERIgOXrp5jajcHRUtAFtBRlJfwN2EVnIX
zSJWr8XK+tqUwASLSKyVKJItu5KVRKTZrRpOjuyBs0ucUiBGcdMV5OMNZybml8ea
ezU2g2kWReBAYliQmVTcc5NpjMmw/FQqLSudtVdCpeLRzlmD9MHEnYiik1+idQmt
sjvu1gWAg1skTYKeV5cco6g4caajY9mgvEVtOLmPKZXEy5qh00Ucgomy0uRpA+P6
5zHYslbNXGWbwpkyqcrfRhOsgn1noJlMCNDlNbN73kO9mM2Hbv8gp1iZhqVeVc2Z
b1e1mgEtliOU1WapMUjzysIxl2iCH+Hmx7/ULKVfLSbxe3OdYCbCz9TsxQH4qLI8
0UxyTe/+K9UCRkDuqwJMXZPhG2yCJgsyGubz/NOEDYiK8FyOAUMWrqo2SWFGZ83s
0m0KbhMXNaAMywxGgNT1oBb7WmiJf8iZzZ8nuxBgPCKWkTFDJusLs2RDQzB6vgnK
m9cvahApwbzuU8Zk6iFhnpvQi56LmxUsiIdK0v7upyh9OsT0pmgrSHVZ0Lp5+tok
fR74V3bG7zAoRGWSbrQSXcBXYLGleswvzngqFP5hxzbJbeh9T8WmQjKSgqJzo0WV
U+fN74KB980wc9PIBIM5pOYKgRelnKZ5JN8YsW/AKdaeWFoa5d2bDt6DWeltSz1x
b8iTN3Av92i3yH2YKAQBkjZdT7tQBVEu3bF5DPFRHYlKBzM9QRAQhqRYCLMWqjPx
ToPb+YmJ2coBmKTd84C7RupRh043vSlpPMTTZJw66VuLt9edFozsf+GZME4h3odc
AufRqdIyIry+9sBWgh6ZW9rcLFn17VipRxWPqQYXa7FLIM3nowadDLtvJ50CUwCt
rNVKL5uUwsm5j5tFZR1kdcHhmrZq3qBtRM9zJwLYouKZpO/qNLnk8B7R4jFjmp/C
MkHGNWan3zFyn4VqELm+J+5ycwG17FH4eFfW+MKYYH3kQdzYVCH+q7nzw83OHdsb
Md88Z45uZLfxN3V/FyvXab2skpRRv7IxtijvlqXPPLHD4jtw+vKYAw8ALAGvChKF
bOwFNhMAiNX0O7iS8urUScOteG+vs5AX2/WpMRppPbtGuZoNMfRSUH0BNcJS7ChC
LkyXXmYF6FdTX7r/0S0FUZoKbM/bsrkmvDUhqIcqa0F17CkFWMqgGPcqYldIXMba
JhdU29ZnhV/GcW/kyAnTav75C9fFbeNY2vRHaMNg+SMqi5hXHMInJ4SjqLVh+2gr
Tg/4OqhC0v07UFtAeEg77GMKffKKel1k46GjReyuVS/h9WjI5Gcop4W316X7K9CH
qbGqf2zsV5bVms7Ce+683Y1eIDlk4o/qBNfMS4IwgZ3HJ/Dmu99u/jZELiTukCwz
VEUxvm6U46QbuUj2T+UxbW8tRrJOYqrOqMbFEzMAHi4IJG6FhjksGLsZWXhI549A
HdFB7C6BAa5q/ViwQwV5vaL09dEXgN70sw3iGKTpH8ZxT9OGtHuOLKdbt2WsG5ol
l7GzqLkkpUmv5QbzB6DHUfUK2woMjUVUUuey8DJvycsradD4q2Bm0YGkwgIFgZ1h
8ckVPt7uw8FQenwXH+/gZHmUYRFnIMuGe+HUY2qMwzKg0PEh+zRoqxU95eNCmeaD
54kLW3T8HA47qKET1zcNX0bHAnSVnBFeP9bXNZQPpNKYfX8iG02YtsM6sToB8EsG
gjhaP8eJ5qX79JTrbaCgGCLtqd5fdnOHK88tj8Z1PCNSRAdqwKpnpn/fS41S5hYn
F7Qp3fLOYFrk2DjcJBwPzUd+DG2MfTTIsl/RBVjvZaVzos79mqnRtZn3kAtNufpq
k1vKDBETf9h50Cy9oycUWx617LA9R6Z1FD0OUWD72jU+Q5xWso2H/uLP/Iy9BlrI
VFTctIZWcsibGbjk8ojFgoBmpeAJMHYfOqkzZxlpbkUWG2ENqrhquig4PboC9Dvx
bPb94gwAYMXm4Qe4N7u2L0ozU7ZqNoWDUTzrBGU7kSE0IXmtykbAgiuuB0FN6uHA
b4XVIW5sfguL6DI2lbU4MbWKeit4HIo8nnbW7HOoJolqpzKJHh2dEnLoaawh9Noz
NFWO9pjxBs9yOOjZQQ4ykAORbTVM2wnWqQYXCe39gIyGruqwRBaq5NFXlX47vX2k
dGXM+bAgp/tU3WmIVgf6u0uAc+kdgLij7HtAyeoKRPlYP6+9PVA6+VmODO43IAvo
dvimOWtXY/jftbCRfmVaLBOiqXZDau5KSSIeecfyeL9a/ppyUySp0mxOHxZ7BV/r
rDp+S1LX+d5YYUae1ZbXgh2JduMLCxpKzX59dtSLTvI86Yt08DD/MyFtf6iHyVL4
SkRtBuNEyzsF2V2148IaJ+ZK3bUWqu8DTOmPYVs7EaS9xaA779/ckBbrnUKA/2Sd
azhTiJ/KGdJNtmC9FYFLLz3WiXKpiCfv0QRZPXhYfbSVU5mfMQG/L/UwNfIPkhQV
hprLwIv+rn6/97q9tI+9Yf8rKi2uvoe9qCXgsVnEaW4G4Z0tN07VAw/iLvRpIKDc
i7ZpRxPkS7Aq6hFLyn7SEKR0Uh+lOXP9LmsTm+2HDogQaReF4hbCGTRf4pZ1ZlG4
FrYAGb7GfiXoTQ2KCuIRjc6aAE8dRSEtRf7+wIJnFfzCq0dxCpyqZ57bjYykC7vD
0YBXpuJ3eRS/qse+X24kqFaBQ8ILhUZQfCVAGHXJEW1BQNHGgQSpo65nc9u8joCJ
jk7SzcIvrC8ZQC5eVheA9e+cSTmhCnvIswePGcOx27ccuG7xpfVUvMShEgZWpj31
N0SC9YnpAR3AprkycSfr2QdSIb4ArjkiU75ezwPzFfrZ9Y9amsG/+3q6Feiu+rju
6tywgkVUch4IrDK+G2V/zky6dEjYHA/Q3CN1mHGVydUeW7Tbl93aC/rzHfqzxlRP
miklXocfUlR/J/Km0Q6KI83mdPgkdYc7ZHQoS6vkrGXK1cwNzUqXFCD/B2/bjcVg
vmA8MVI4ShAPyYYCiVa6wJf1LqYVx6FHzrgjuF6n/srK2JWP0XSU0rWDR/jss6Yo
new6AIB5ctYJt6yUm1IkJX6iSRpGTqP7FrYjHGiBLEAb6deSdMscmddxRaY77VLX
8SKcGir6GN5LmLUMYLKMc5jHl3doEmlPzoWTnI/6Zjjm8ECB1wvs4mqEnM5MogO1
TS4vLHn+IYXG0m1HsTjta1JfROz9bZqa/tPlJp4EtOVb+QAz0exozC/1wWiedY68
RwQ8XW9alW5QxeIt/zQyokbm21rHJZsNQYpmym0F8DXYKN0lelCQTJkOPQ85CfG/
cx13qyY7Jwwx+QuP2rBj+cv6WUarg1wjWKLX97tPjEaI05Im24Hhj2CKAYlurJCf
MOiw/Ge3LOea+dWBdhyihD3sfIe4AzPCi1QAq+IO+YEsj+ATrEH/qnZTmvdGw7en
R2etgBsKoHDT3zf8ITMFtDn17sULf5WmOjdFafDWMyGSHplRmAqvOBKsXNg9io4O
oIf/VhNfSm4Q1ADyr76DQ9SkXdEdefR+N40X+yKUpmVCQMTun8zzFBdYUDaUS0H4
v2a0ma8Tz+cGPJAW1p2QA7FbH9SopRJrkWBqpO0VTSGMPvAddcW1+e5g40JP2n3v
yen8z/i3eSCwlO0ZuBkyd+TOSKNQMRSgYBuLHWAqqA+XqThji/NI1Quh9ILMWZA6
LE9gzrmS6Li0rKjmqEBBw4Yy6g69Wuea9zi9Xb/O7dbjeHwUcyyOcZlkRA+c70al
V4JTPUQ+LzzOMHYO/DZVEFhkGg2lfIM+/jqbLb4N6RNkTDVK+ZybSAeXICe3n/hE
kEv6pwE7yv68/1Sjv5QG0sM0cU5lhxEzUVjlDxpT39dHUksrSkx4Y64xQ5VUhYUN
c0Vsm7yzRe/uNjCkNJSOULRz/iLdjDk1m+OTKWDXbq6TBbJ63IRzUwZJSAKvp2m9
If1ubjG8cQxy5zT6KV7+0LYRHjJby31rVlcQSAWcf3HLZ6xJyXVLooJGUExLpV8Q
DU7sLZthy29dcQjk0Kqpy9agnvyFmZmTn3tSqXed/XYrgxXPeLaKFBPf8zUE7voZ
7CEjCkw/E4bWI6D9DtvODJpDgC3wcox6sVAttCsvD4F1vcjCrwXsn8neh1XKuJlt
+g5983RUGOs2bx4Rdt3ye5CcL12ig8tvrQ+1TIzBF6htzlilQGuxbTMsiJadjNWX
O5R8nV07DJgeYP6v6GkjMn5u31yFan6vhh4IUuxFOUyw4es0+ehULH7s8inoy9aO
D2tHYhgW1+yozpsKlUuTgpf2QzyrPIwu8eJLqInmuYBm8WhHunGgwwmikjR+tUxE
KgUJQI6IkiSTqwsBre9+qg29sFo4/ORpyQGAFdUo0JoHeQD9HCFIVzY2nn2obSjf
V6dZYJsDvmPhy0r5PaBiiirh0G4JYlhd39SyvctkPjr4oJXf51S/WxcomS9saMdT
z9mjtZbZoJo507XC2wuXIZrddgm+crnDi5x7vr+PFP7Wjc4Dci1F9xo4atz00QGJ
aJto/t66UTQDIM2wGQe2kPh5ylfxdGDL3D20l6+rBIMLwAMi7VCfikIxi4nAO3m1
Dn5lY9ckbqJ1ouXXximxFXKOLFrLo9u5poX7YuvkZhRRhl+CQju+44kqoFgVtmzF
oYM8az6j7RgxBIHXsKd9XfWlv0flEeZN4bx2FpuDCGcp/tTL892a4NPYaRj80bxC
vLJ3+V12rft4nGMn5FQ3NCUm2oSoPdJlpVdEKN5PAv3rOIiyXeimMSf9zE/9n/2c
R1TTruALeG2sFhKTfd0BUh4hQRpJLQQEm62RJX02sn2Qk0C3ywGNo+kjyD682oTM
bwup7BN2XbqwpFosg6eieTXq4DSfas2L5AEi7s0Le5+n5SECUdhbamIWFJCsGszh
I4kiJAWeaVENg4mEiMVZcMdEvEpxtxdEG65oE3vFEX04BA7O9syu0YpfUNYpomJj
X3/tiRAZJgxSf5LHodBoKjTAcxY5LEm9QKXcb7cMqOIsjHBMpHqumnGhGFQrXBEP
WWynS37Op2erXRZJdo0UIrIz0ws58gi2Oo0j87MmUtFL7bcHf+JSPoNZ7kGuUZes
i1DgdiOeieFMpgTqU7dzrLtlbZ0pGKbxdHdaFL7VRvsRPFZ16EF0ny3MHEfNpIdW
+11NG7TxvsupKi6riY0R8LppZaPTOi8TkI3GZ7s7QeEhp/Juj6yLxw5uGEXbeb8n
kvsmccPZKGrKdvh336p8Zi6UN9JX3EJEYnxkfUaG5GqLTejWN1p13daf326lUFGM
vTH3vRCdtxuVRX9+ga+twNOuAoQs+sI7Cf04v69/6loylVObe8yMMmvdy2PXn8ly
4DoYjB1kr76nsQPPO/YoY79AuN1Nh5gefIsc0XYcHVo1HGNX6RlQpLddiROW1hLv
DQpTMjp6/8ZtW5dCb5/6ycGG4DnsnbDuKgZSu55SUV+P/LCPglI9vlf9ypshfo8S
eysKrfjtc2zwhqszZV8gAjH++sxbK6jGSjdNgSI2uIYatqZusTuicMo4XC9ZFAZ+
/rootJHrJ09zLDZ4XAG6QrJApgG8ynfA5GWoVSif1npvX4+/qWwaFgP9HE9YoEJo
Y7vVfZc4Kb1DBqqYsG/n8FVv/bUknBSPD1QFW0C80yRseFcfbm0eY5XqGXbLD0tt
dOvt6SttFAq6RxfWp31Dzz1GeV+WnQV7iPiFaz4B1BYQpjkflC0M8scuvdpuB5f7
VBawvATR/qbr6lm7UKYuu8OwQG9MaSoKYgB6np6OohzTUUwGnZcdBjLMSgkR87EN
Ge3yd0c1fcdLQ8qjYZ7xUIypqKo0OKJ6j9hIdS6rYf9C2384cBOkJtMtoL6cuBAQ
pfKmbPpbQYjL0fDqJ2m4ZyOdtyel7TsdIwaYTHw+h7CPxAfzUwnhtaAHdh1UwHiw
hGdh2Y+kOsUTot62wHXrgiup9phzvyh+O52/KeLoP5++1IVdjb7i9gHcsLH80+X2
iKAX9uLAYriApr4DQhSDNSgir/OjEsy81k31ViaIqSwVWFyqw/Mdkep8VkaDtPjN
1Mf5/5qQke3Z+ZX8Piqu7FkjLVy/Vv3mxBddCvyUEjC1t4KBBSd9JT+Oh5Ft8dBk
KwySI1PtQIvU+s/KfSjLVhCVjiDLwZzYar3nh2MBYDD3YyGEKbATHG3NElNys0F0
1QB2E2hXNqYQwkV0ANT3Kc4vabVeCBfzeOGjEtmrLupfNp1yF3Qy///8gTwrcfXy
HzNAqaq+hMpbPPM1br79xuEL0/NQ98OqLBzbCHeKSx0wd5WwQtRK0YDO1lOmAg65
ZrI4I3hjPh33xuCA6RMvctNxrJZVwpl/0oq1hkt3ie6T3PdN9Q+CvyFBR7YHHTla
XLxrCpGC/icYr7w6+js8QOlXRFAD0NN//EhlL8GmMJowJZiiBqyKqknSHcRuEFvV
YxTG88WUUcnbA2BkEmjSwcIsyFhj0BNPJgN0oFZu2pORCe0D5NvXgHVLB6se9U0a
LcHISYuiX+xhDRSZSfESxQBDjBLfmk+MIOPKeZ6X2WlDMbHDJVvtJmMgvfk2IMoW
wjwOUp1DeQCh4XKYfMnn+2p5PjjrJrQ7wNJQ9pMm0+SA47H96o1cyhichMk31VgE
sAacAyReVMzejW0p4oo1ty3leWiw4ipnPA1PmfVWI58WGHep11j+lEkokOcRIxuk
dqYWLouJ/9JcXhmZs78JUmFN5YSxIFoCyVb++euMyNVyUTzD9p/PSQpyu29MtFmP
VLpuOM065XKFYeEQ8aMBQpzKBZYd6eTMHU+za2DIarSTHYueQg1tMqCuy/bWvDj4
MTAyjWppfsxwF/WDysSJK0qkc9OvTplcloEbT4gWYGOjXHxqQGi3WxpDwCOmuRTq
rRKo4u81y7nRgwJDv/oNRvA8UvqfXpJMAnboHtm8U90GUSw9gvU7lZRxdbavX+NG
oHD10ngChsTzr+kekNY6LVH/bph/ujIwm5nbKMuwOxICZ00Zgf9b36YMQcMfkXOH
ZFf0PXAeqkifgOZi9xaRlF1zXeSH3quOrhXbBvhFkBPUS16qqpGwlvlx3jDH18xN
KHH/EUjH/dvqdzvX/AYmoGQsyA12bPRwGzc6MNT2DjbG7z8TMU0xoK+gj28lZ0su
VFu3KGFnpXwpRsK+C85JMw+IqmmOh0evUkHRkLuOKcvJua+ZammNyFuYKVDMSEq0
kuxZOLtXis5L9S/OZnF2OGqBKfF+xr5532AZ3k26xFL9QnkE8KJ3e3CUg1Hc5+tu
j+oCez7w6L0khHaFJfAdeA2GiV3mCqW/zK9AchmipcdWdaD14/dGSGcOa8/qi4hT
uDWVrnKvkOOiQFZApvmRd8QIn9Sd+KlIUx0xOtM+gjXoV/xHdt/pIGK63r81/Bzt
1Gu7cEsuZ0PM5X2azROwc8srdnTqZIHrTmSWlukx8CbuH1kcm8svtdyjTp+AV3pm
88qS0uzpcgb4dDX+rqVb/1Wh2osaIaSJ6EQWn3bx8b3IBlFn9zB7REWEDm6CAZkG
BRAlKAA3M3zdOyxZK6+Ri1xPHhd2OXylnQegLhakFvsFMBQEvAi4VHqsKZP3R/T2
PKG+TopA13WIyXXGJ5hPOEfu9+JX/3TbK/Qq58L8zgJdCt6KdqY88/1BtxC+r/ny
lo79heNRgpc4diJ3U2TkE9I0laD930ZGFPx65sZdIfk3udxjjXDKwJTWYr/lNcks
GhpfyNvKd95pt5sU4btLCitvf0ljwSfkQnz+Wm5M/qcTtzDnl92Ubc99+KF3RcPs
rT2pDj6LIqy0AZil50DLYU0LDw11DBri1yhRMtc+KBq/0DLRlEaqxrF6fl8fdEP9
a7g5a1JdQTRJVlFEOE+D0KY/2iFjqjM7C8x6dEWJk201KAOrMqcCjyaC3A3QkMqO
ya5yw7fpamzuYOoti8/5aF4+YvZdu/skyn+1d5BNK/rPCU2xnUCQdZ+d+pRhfQo8
IDIDF/wMlRyKeYnClWM+ONs1ulwuOYbuhNbiZhy9n43KEOH2lAEiblMaKqPNG7Cu
vPjB4AOE50Y3Ben5g0SXm9jlFQ87Z8QgYJLdtXczKMf8U6nsALu6hGc1GI8QbShO
5sQbitW1sgv16MXqRFhEE1j2aIFxCulEMg4GHWHNE/gLPs4uCGg/Whz4mQtuwHUp
ZT7PbQG7O07nip7sNDVAc63b8xL/durBJcVGw4Elezmy1Ni9tZpbnQ76e7U745+E
Dnb8KmkdPXL8WzH8bX2k9jOuPnMLGBrvZYrwCRExC+DAeQtAB8NJotp5mAMFJJ4y
Sh8CNBqTYrOXHdiBEBtqQOE1qZvH+OpZBCs+W13xmFrft9t9pRd6PoWSpwC+ACCF
XyuEZ7cWh58ldeQLRpi1ahyGzww0i8U9h0x5fHlFYLrxRtXUuZmVDsiZhMpTNUQE
AqLOzbW7DdUuJA49tT0ERPhMj0TZJjHrY1TPz8Lvbb9vlR2/XSPFkTHFysg3M1/x
NB3pLK5FJeyg0U0aWTf49EM1kCozoy5fT5AhdzJ3e9HZyEOPBrTtQWeGee/f+45e
/SxiYcsk7Bn8pl39U0Gmm8SWRQzWyqNmR3vwZZfGH2hwiGSpd+BgnUWX+P2vfv/m
bwIkzPRdOgwQ1p1+RrSC1VVjPifEWpcrOTrbWbqQZcVQ1LR8z7XxCylSWgD2zrRU
RaqYBt/0S2C2ai1J/BMNRlS1mH2Wio2Td04QI1AVz0MzLs467QX1VVe3wmUSH/U6
aB485feUgIzZ/r3bejI3MHeVgxD1e/C1N1HyFXpvSkoC8Y/NZxQgJGe7AHAAX1um
v1cf4zabJlmDF4rEdAMNe+DzvTBk9MeeykcK87ROs8+pgH/B/F/tiDFHMbXDD14G
uXKynOKDvN8oNoIx/++GuT1l8zMwCCi977sjK42hUBa+DiX/bbZhfBg+EBzpYZ8h
iUbk8+b+MB1oKyIL8YzHIPPtRKaWn/xj8N7n4ZgDYZXRP+/F7pIYBQ6KVmMjCyZg
9QYZm7Ub11yioHuIAW4DcOPwZy2RARhejuj789qMZHuupkKMvlICZdZuGwXccVU2
0d3xKvyBjgZ7trYfB2epMrsGYBNtrrW3C6Gi6K3i9fsX1qymgR0bVXa8mubSam0t
iJ5I8ieOcgVqTsPg61e6jXAWvQeEJduEu5I+QB4E8kq0mlokUduwqwIMDbBCutDL
0V/NOWjdWbIp0kOt5YymZccvpSxmddsto1XkrivTMuwoLFp8Fds7cRiicizWg76O
y1q82JrSeg0JdtZ8ZROP4nCmZaziBw97OcLCHG46OVaUyp/vKiXK7B45Hs8wxgtE
NMGZZe3Xa+mfDZZ5w3NPFOMo43IqWrx7l9BlOKwEHjUX1mLQStBg9xpGyc9J7dtI
cbeZhK3w9j2TLPyYASShucsAZQ3xiNtaiyBcXjeuR1xYvHXfrNMGghVpL57I0HU7
vsOSQvDWiVHaS144cq14gxQfSvPI3oq67rgQlUWxflB0sfJSIbbRZSp6W8/f6sPC
tzxwNMO24e5cfxMbEnIeyuDRKTklXltWGrRqPtSjTfzKeGcU2UqB6G973bse+lnp
XJH42a7FlYhTOL9MnbxIHg9xhNcUDn4R+SrGYHOF0hQ4XSpfVP1xG06hGdr9x+ef
oBJPnfCgwMOPIgt/xMLTCig0Isy0O97cQdWJz1Awgc91KPwcNggOYboyKG0OM2fN
mk12Edu3N7tIOjRIQkh6ovZosd7bUhlHC2IulsmXfj5yRUHmDB2xmhPqrviYNkSe
rCLYs4BUtwAlTXuvbxcp3ML1dKBod2GM1sP8Tw0Dwfj+QaMAANg9T7XnL1OjsRIc
Ags3P0W7EMc+ghPF/qZ5uoCYkPlqdjDVBJEoKlT2La/IgGhVqloHciaGW5BEIjOS
5k54FlnbkJj8Rp8kpEXss5jWP90yoTlh/C3NVerRa0cGfYhkykyXh/oRlMzu3gWL
wN2k95Rp3gDd3HK7GgP1htpeFiOd+mOjOTsNDG+uzJWI8zqEXLwUMCpiGLu5M9B+
bvlqmqGrUXBElNaXjIfBDWU7StpYcJFnzAV+Ha+4FN2BgNaiUOVhywrQJ9SdkR1T
Mq1FBUxc0a53nh4Gn3wmxOWhPVJGf1sPqDAklWT+spnQ0tpb8rUp7qZqmS7gzTO6
MkbYk+8a3fMtaObPv7GWwH1hj48ZrWZDtNYjcj5Kv9kT6bwSvFsVSDjwwAhbPjan
oC0sMvMobtuwLM1F/AjEGL5b3AAEQ14uaTnGTnsZYaK74yR0ZgGpzUUppupx9xMM
ET316VpQ8fkPFbBkVOdAouB9KwM2J/nA/2Rew8D+XU4rdtbP2Fohnuf3vYAm7bhQ
PzmMcvQ2Duh06EUVjYaGG1pg9lkpKdgOcT6smja/Lwvc5bl8p+9JBpFl1nr37FOn
qqNgJ9UwGuJXoXofscnOg0vXFJFEYosRcNay6K/bYHHbZpLZ8VVFRToalcVs039S
aH7bwbJNWIrioigLa4LxnPKo8V12dWLMhOPnEKuihuEvhGzy/VxtRCYVx1z0EN20
ZBbjX+i+RQCP1qs2qVlo0hrTuC1swaCWu9mmxuCUjINjgG5QrsJOJqov9MfqCpc/
NlRG5JaQHi5Q2RsGjztg08JwqrYcaFl20VrVKrWGoGzUX0TcniSjlZ/uU/kxIMo9
VMcajpfEg8ZadzYAAgR2Rrr8XE9c9cQ1/7EFt57FAaRTFfDg5fE/UsEjj6L0b6Aw
P7s/JzgZcdyGeTbMC+m63RV6xT0fKyprD+oZifYLhPika3l0gaiTGLo9/SiKbYAd
pqud6j1bvILeT3LNp9DUOKpUsLGpjmWPpZNF18fubrEdOpwntOt3/32k99RckX8u
1nQ1qg4eKrOfN4Xaanf+vRfrPnNY0JfrqYazKKKIGAjDwwoQ+x6CaRTzjZ3Jbvhw
7QI1DrDW5MMDSzoV7ESG9fSIPgBF57H1GQIUxGwbrlAnV7ZWhnlCqn+49KYjfjrj
QZ+EW/NDJXcEZcAvExC7zAhBJ5NOXGhuAc2L2cICRrAbaPgYlUOLwdxwIbyYIw36
vIpK00FdyghaY9x+lFV0c3VlpFsQ83cYFETKaRkNTc09JnDIFWPOrifVMjZ/GpHz
3tSmfTCj1pEX5vnTqoCWeaHoiith6+2J+d14MsMTurugu90KN/5lS+NYXuX+CHGL
YubnmEp2GiOmGJaVha67y/KSeOqIOaxG9l9dsxXCUIw+YAl4xg1Z+PMfHqSmKAXD
u8D5JXC4dEZ8a6KgM5u1ALnU/a1uz8V2kIVXf3lW98DeWnrHvzW4+EZahi7aFPW7
3ikMitkk+Xkp1SCW4fVL2pPBKxdX9f+wM4SvSXi7L2KWFXDosghfcEBSYtS9ucqN
HcTpUjY5iloX/6nrwTpFS494El/s7xb6Fjlv0INaGys2U353J1Vxx7mSSOk2jJif
+AHv3f9qJMqzESYkP8aV8qN8w7rrcuHraZrxDE3ebxzTnOg2ZgSsnN3R9BRaZxTK
77T8lPsObcmNzJzFXuYAJU1EJuCKA4xwspN7g7IivENUN7QTA/NbpxBR7oz7cD+F
pFBUtLT+E/rIxMpQcOuZbpLM+6yVFdj08Q6SNySiClBqsUOWfK/DS9b/Ohb6s3By
r2gqWfE8g45WwdRlNyc5vdacE8/4hJQDs/CxElv7rrPjwg2r+RY4Q/dSv1e0zjq+
XzWijjG8FwZxGESWKVpAS8wwGFdONII+8np/CSiREPBGZXc6qRWtfdu+j/DHF17x
s1JHmkIWHpiQ4WgquBgfPJivjUuvPFLF881neT/FyJQG+7Nt1PWF0rbPrDwL4f6f
b2ymQhQrXKeahT6MTy7bjlTboG/icAHW5HV/VhLmQKhj/GOx44qJCBCk+JY6lPZ9
ze7AIpHvFOwDUtkZoul7I3dPYxfoGpHtIg+tqArsDdwDFDZFNLZIvnrexAraEYnA
qXOS/UUU+SXmvnuGcqePi6E7k+SPGO/MurpjF+uUFQak67SUgplpnFyjbbTWXUxM
8V9mp/7FATsfFr+lEDqeAXDoeQUanCRU+98XMw3EGceI88HFRNnRtNICnbaQSKk9
6qibTKoo2YN9pKaBSFdClH9CZ+2dpXkCE3Wan7Whdm9rRNV/Hf4ibyy60hMNz2f0
YlHAIWaCP1/p41JpCixBwuAtqwKaryHFgDidM4HrtctzNLVq0OQXngZF9eOCdaLD
WreLsnW9ZM10lOh5Sy1xMu2AQUpw3oflHkTiMXK1BrxJ4fIDofVj9aYQKNh5txSM
7qNBqqZYIewhwdoRSySfB3UO0EH4RWMmaJC0iNu5/e8nF3N+PhWxIKhOrP0Lh7cv
41afqrIFOfKLsPK2D4VZ5AOorHcN6KZV/XRB8eFjsbzYLEgFgz2czPfATywao2eG
i1+iM8q9bJqIU7Y6fGSkJJc3RTop/GQeJzG7jJhDdDXqDMNkSth7++D9SyVfLAqu
qhwhQhVsEZ7NAwstlEjSj3XJ2gWn+ShsrCZ3KW/A0lZlVwhrN/lwUiU0+Vbot4HU
OjhKFLsn2cM+fokjdaQ9wqWKFDaHnOr957owE3qslyhR1i8VEb1aWfO1xjoY7o0B
ab76Gqt5w7ZdpobNws2pynwvtdVOEY4QKGLDIfzFybX06lHox9yiitnL4r9sbNGD
YMYWywB/JJAhePhqnBQI1tOy7V75r5ZV5Gssy/26VDw4Lyj1V6uc6aDTNaliHU7H
zFdbrR/awiP/EEwWKa44cAMk/glbGWD8jbfsvbDRaEwrSNOjTUlxxszES/7G7ji8
StxYJFO9h6/q9BMSkfGZ7EWkCZa9k4ZjKjBI1sL4d0zD056coxHqV59xHgs5sOAK
enASNcn10KqbuJ3lGrv7gO9H1kxw7znSK0V+3qy8GBx3mogmKmQQeaajA5JKMxze
MZ6wBQcyaBi35QQku+gcRT2EUeAPrcZ8bIUL0UZIpJudDvgQ30TWZ80QeBraulZu
HE6UPAkOQUgrvzACPej9jpS363PpyEDmwVJ6wq0W7KyadSQ3IU8dmXusGAsSnC+e
7OlA/etC38+S3C8vVS8FYVPlMKgYBugYt21kUmPGbEAqRH/+zs7mhrpDwSf0mCBr
yeR6+E9zFN+LPLN3wuLYglTAR+/q9o1vmkpOUqPxMA6YpLkoLXErzcPtijU6NtzS
ECGIris0v5niF+Zz3MAj5XCCXSm+jSR3gIqAaqqHnyEWvbBOlm0R1SN9IzluBrqO
34d3UC0B7wuDEloz+nD2FhXsHJQ9mVaJ/4yuOlMRIgZ7ZecwprScmjjHYCn4lqCw
NU0KSqll9Q+suFw1i6M3DZPO/cJD8jW+LPM6sVmz7N5qSg0ds2pZSSXBX+xujWEG
jFXXc9NUlgMjUG6Ouq53xEH9n9qFcMBhj9zYf8MqAkwp9OA6ZJM5jWsIrY+M+Jzp
khf0LKSGRNRdaXUa2O3eVBzdL7eO/rEgtikavMySgS27aqHZ3aHW3h70DbDmzoOj
mKe86YJLlyozuYrroisoefenB3cX0fDVBby74LK/88i1cWeq1UYX5D7y288SwxAV
biwJ7Qitwzd/muD+U+OGdzvopVZxke3twip1f9DXtY0Xu6t6LgKNI2FqFCkzgnoD
7iBKoI1XxyyCbMzDZMg1dvr/tTbY12FqsU3o3C0xtIcJQtD+XZLBfCsPyJuiE8cF
FWCB6IptVNmNY5t9fbUBcy0LbNHcuIXGjyenuQ/5RUjrbGAu9j8OW/SRYRLW49yi
XADKaNO9airBeOiVvoCV1yORjRdPCPrrydKSZphRlRMm/2bWAa76CSlg70YY9El9
KA1Tnxjh8Zdwgs4WuR+BJ/XCdnGQ5nuuDMjfegxQKtPS7KWAAB4IgWT8esl8wHbp
Ji3iTo8xFEjNQbA8z6E4uaUKrP4SPcbWroiNM1O1hX5k9VF2xkAUtRPV3n4V/Gpi
ww9jrlsIpOGdbr4GpHoOuostTSwq9fLXnIjfnktMLDN8mn6pw6IS3qFkyjSkEw+e
cnKEkc8WjIhxU95OJrlzO6lZ9l+kFBVPUNKadu9I6BC6Epkqab5q1DAnVxEFQKqK
eAzNZ64zM9ZaXBwQvkjokSkUYQXeLH6Gc2Xr8mxDNlH4qodtEi1ANztUx2wZQFwi
+xmcmxFwGovYb9MA/GP/gVqtkXLZihgTPDq9pZqV88UREjh08w5Sj0aMhaw3lx8g
rs95tVIrSXjv50q09RAeS3un7WyktiIdbwz9Uij5bglcHH2auUdBBGjNYJOl2VWW
N/c/Tkv8dvG0c9dpa7eVvTAm1KI9M9pEfrgFA7sNKK7Gwvlrg9DJ+B/SyLgCsYkl
s2q9u4++bQcomArjUhTVaXuy9Sz6SXvdMG6swvfT6gFQP//4ESd3SCK79wll4iFY
S6xWv88RLxCW2671Rr6hqJOPZZSTlsutZcSThW8OUdOuQ2XAhTW0wVPNAF4A9KOJ
q4Hy0ERJiOJmWNfeD+B+X1Gvh1fnvX/GzvQTmLdADxyRAO12E9ad9URYI71MSy/F
Ely8ciE3dXfAgO+O/GoWZMDZsGusWaKENZlSWA1/R/ntTT7H21pCzKw5sWqSjh8w
XMdsJPeb5IpDKdDXed1Tzn0Ypwh+EoX9SUuLqNdz6hzgHnBm+XqL8SOoLOOQl+oh
wgK9i7baG+D+zmQPO+7F2TQkyJGgENaxBBd3q3nZHJT0OuL3kFf4gi4p5pNxQOef
FHIl3frdB5Xy3+C8l861rM4FgVUdR30R+jfrKvkNz047GgBbWN3qQJKSe1ikmY2k
ck7pU2jngYS8dM4j3ozJXSJvP9uYAxUYk/JyK47QuHb+r0cFmlXissqtfX8IO/0Z
YlSeeK4HPQXBsBUe6wsYz9z366gGsVegX8JjqjflEVBoLUuaXALQVl1L3NhNtEw9
x5zWt4G1zoEr2ImIv+AawWQfzejLfnameSEvfg8irYpFV2qRoTZGQT5hIkyPBOi+
ZzqYbPgbniGPYXUUEkenTzS47jfNEBpqOEfCK942YEYw56UGNCoGml1MB3TBgv/V
BUHaFO6zol9myGS1fwYz94FBm861uZWz8B5AqIVa3MAHOiCVfh8dLb1mg9DkBBoZ
TPk2CKcnpa+rGXxL6v5W0LhN+X/nZhyswoOHdfC2LGrzY1rMlelkQrLUrG2Ug7iN
4OnJ0pYwI/5SlWkJ9e9yYeDPT8PQ7hvi/8AUiMK/UPEPZdYXGmLtbsEHhLvIYT/3
eruue538xHJo6BGZWp4Y1ffvfevuCDxYsBECBnORfx44CYP81r/bnz6pPbBGhxPZ
JIIPWgp66ypCRKioej/G3661wj7Z2aLwl3APfR5uY9aETrHRg39X7DyPj2tVXSWd
zhSFv3zt4ab1prmC3/2Ew2uCY+9ggZZkvCyDgqM9+49gjWc5F1RuvXezgHAzvvjn
OJLbohM2VQOxsd5TJlmYNPwMTFcqlj+sn1mTfWn4Ex3YjJiAPWEAKXzH+pBF3MkK
0jv2FUbtWS73U+BamR8vvim3u/6rR3g5iUd7pgLvs1c/n+/t76ad4z9UhD17TEs7
zZk341fhxbMbvLOnPsaoU6yE+R4B6aH80Sowyx4Iy+VFb8P0kWMdQO8fTU142vmk
xg0m8Sj53w26+TxOZCHbf1Njt9Hd5p1LtbOTflMwSiVn5Q1OwKxz8Yy/qKXlXh1q
8IpojL2k8QndFgPfNQEwVbJL7wDa8fau+TQs1he1ZLnme8LQLLALGsTglMrSJCR3
mNYW+Fer0oYQwYIiX9mRRbiuh0Y70f22/eanpBR/8HjwRSdA6VD4p1kv4gUN8JFE
opClcNHFj8kCwBb1wvyrUOG8Du9infezx3fSHNF9uUkwk2kWN1/nJpH2wcvJXAUN
yAsvU4JmgjMf0EQT/5/clK3iiLUzjs0d63QasnMxKx1zMOrSQnddmemvgMlDcyUm
VMF3109sIA5H/Lu9Fc76qj5lEo0Vac7s/JhswLosIcm4AfRjunPtibsFjEsS4W3p
kzr1kX/ka3GFM5Xh+2lpd2TAdY2K7MDQaWrivkpy2QWH30L/NdEJJgLilOpc94dM
3TMyVBcvvSYqjz1RJqH6VnXXva6ZktfNy1dO58ct67MVEDJrtXIIoelHk6fGGeGn
w7ShEmX2W5aS1XXSEuCJL6Do5Gn0Nu1CePtVvckOJMotn5EcxTZCISMue7f2dRDs
ZGCF2vpxuW/+HQ67ZQPbZjyKh2T2kZXnUuF97baejmCladMGJOLnZGMJEIcw7Vmm
ymV0OxDQPQTAZhcTL6bVEpbrptb6MFvgrY8WcYq27tUee0VDGCyzVRpUA3n8Yssy
GLwJC1qVLtlmbji5ja7L1jIYJ7NQmSaq3RKMecwMhami4Vfpz4mDdPunG+n57YuB
dpYXg3r5CeN+9YhSuu+I6UazO80Mne0dKMGQu6KS3MFYEqY3j40O7pNu8WdYLwtP
deEs7LZ17RDii2gH1aqIt7XqsVf/c8PMGkREHnDwmLhHLsyTt60vLJjUuIL0NAgy
auSnV6KHRoFEWHqzEAb2/EOuc8ltvlSN6eyeoZktQVLxjwK9dvE1rJZT4LTv2ji4
BjpGL0hkmtJiaj09F9KgW5ARyItznoMwXzcFYdGfbmU1a216WTd3DXID5zvngNkV
dLruiJCDNvx9NY72UPBQrGEZRbg8ZOjMxhLyYN8LDGGLN1VGVVOFcjzLW5zG1Bo1
tZEVGedoONE/fJ2rZBNXTcNu+oAWiWLCY3RVKUAN8VPf8WfjglHhAjJX4IuwE37z
ivP5tPbX9AmXu8l+HH1YqY/lDwjY3QqKDpZt6OzJV9ri3YuVR8adwA1Pi1gJPaGf
GI5XDfO8K0RYTMcaB/a636M6cw3OFU2LeslyP3xEcreDZUhCJbQFuIlMI8luP/2W
awtibB0voZVC2dkVMGlAtCVbJi/mCtVv5X8fxF6aUWXqZNtfhXVjav0L59E9WX/p
cC6qB4uePkzIAHRcYjpOjk6+TV+2qdf3lLd1dz4vi0WtNBykKE70+eQfsDz0943U
IPJ8sV5ExBEVftQ2xyNLz1UBQq2fGLN6No/K+AEAGVnYMbweRjW8vX5sOHIzhJZg
8SpnHuVJGh6sWImpGqZI14PneU6gzN1sEGNaEtF3Gusfxg+ATCMxgBo2aoTbqCEn
dVE4xJ7pQSq5wdgcGzTb/iUZ8PZISrtvxyQtUj5EfZeH+HwQcm0W0qjt8FKUqMc2
1leymENokOqaaIdGjny5p/y7rXTd2+roEa6hZR+jCNaWU17iR046CxETNH4vd6eL
ON9Bz9hgF41zPmBHrCdTxK5xHEy9HyL91Ar9KC0tS/BYMLY0BEA84zAEZCfrZ9Bu
0icIt9Z56nH1I1jj6cSgRZkSn0De9r2Ki+EE7L9oRY6poH3KfyccAjRibiuO6lrG
2cyl+HttbGhZrOhGKXlY0viHmQWRX4pISExRdNPYr6FaLw3AnXPS+LAyLKP1fGjW
5JKyHbX71rHm83lu2I9A+YZOlKLPCJBvSyx40taam4Y4fhnZf7P4RB0Cr1qW1Uno
PpqbsepnawSEgDi7aPzf3WoFAZTwr2tKf9ScCplpyLzsruf7Yvj6IbZu2Ak9ej/I
IjxBGmlsGJQ8aZyvGQXE7Q51e6byePRv/hHkX1ZGqNwtlUkWChvf+AjASXXy26hG
QbpHSe47E2bVZfjb91gUJgjIySyiF/F05YDs10lFuZfwtZTJs2wOmccjdHcbxNvt
1Hp4dQpZpHu+MEfIdJKSFRavO4HOn0IKT9ppLHghQVGGahHLhepkm2UREN+GChlI
97Ya0VHnmWF+t9j3s3oU1uh+KGi5j0tN+n9rTVcXz/PmlYMsJnxGcLg9s199Mc2Q
Brhz1xaQDANxbBKlrCeLMmhF4J0ENUFzNs24JI9HH8NxZtQJ99BMRuzd+EFcdjuw
DEBark3dAOdHjNNzvggr5Ciw9pJSzfUJSNPygvLjH86DPZx7x9ZCa7KaQx9Qv5ZV
wefHBq3XZfwV34NxjR17C/EDRYCrlyUtBWwh144Vs9wCox0Iw2XqRJSboFrykH6x
ZQCutiff2iCAltg7PaHQw7+tn2UGnsLYt4Vj1WOvnG3hy7kEgAWKJjT0IBowiYNU
CXjqXKJxTOKWkSp5Ty//goLG6oMmMGfC7w9DZYpqniD3ESRl8mL1BP6e3oY1QpHz
AFTrmF8RDJ59GMAfnMrXpYJ7diu/JNT4pG01+8ihoExs2JolQBAICWKoxec2UO2O
jRkGuUnmDRwDrwh4t94Vv5EY/RvJDVGG1hzsT/TIh0f9dBuQyCcNCd1fWSopmyn6
XxLq6HI7gBffxRuGzgivBfYkLAcI87Iszd5LbsmFAJBRt5KPUVf0Bc/5Io6r7qib
iXglXyLsagiMA3DfO1GUEOBrNoyZ/O/j4C9kw6FtmxXcqhBGPNu6YpHRwNGDJfJU
kCD9QK4lSs/G+H1JXaktByKccKBXe3onwUPaDdH2I64mGoSWkgozNOiHBJuTVQjq
QZmVz2Y7/05sFoMuRe6F84tv90CXi0wzHX4mLRD++BA+EkRu2eYyz8/GoaQklOCn
LR3ASwnTzUz6NeU1KA0i7KM2BrCGHD6hF3UZutKoZDaq5vd0TQCjjxa7M6BMEC3C
Lo8HxLVsh8a/EnyZlI5G/+4LKxiflX/450ArEGu7omVVnEjc+KSLEnv60x3Hbmwn
q7xWd8L42IJGM787eixw8AciqYWHas0n2dt/fU7yJ0zXBfApMYbS8h2+bbYzYwdx
821saPqwPUEYOmyhwe2pxATbbGJ5hsqCBCrkoOFFFMO8xB75MduGASRotuBfOgsZ
bgp2Y85XTMPRz9CxqKtyJXYhUzUnMakOaDI4czKnR8SZBSsJ5GRVB9XaQ6tS3l2n
ff6DvVkBl26jOIcGBbCRZvsEDLFFoE5arinMN92CBaavTWTKkpP2dyDVxRezH5X3
J6iF/AqZcwHqlGLYz8QYScO67ZWE7sW4PnSVb848p5PIG8SlH9nhByAxsuOWk0ON
RziVHrVfZZTJ7vdOQstokSg4mT0KUdLU+G566NzLY9faoGrRPWC4FvROaI1H2L8L
5anRrJyUlq22SrPAv7epDNE8BhCmMdsCPy/+nAwbHtW8YmQNqU0I+/CG+dju9wSw
Csb2a8rZbGmC+7jfhBU8TbAfCkHOcCb/sCwrnmBb6SoMFyVDK7URFShtQLe2vJ6U
s0oSzrUO6caIv3lgqTlbB0BxVPFpP/rAP5v4noX3OZ0sx3uVTq2Y5qMOpG3CajYw
WqmRp39cmmSd5RbpCfcu5ZWcuDyAEyecy+wyeu+h0VLzSS7LEZUaMoThIoW7ttd9
nIkYXnamweI8xwjiDmCctTuBdqTGYOtLwkC5cd2DPde2SxEQR33kM9Q6hmnGhZvz
UcwZ+tnQFSdTnSqkbFsOR8f0M8bMIFDDsJRCggRZVyqtfIGak2fKqk3mjJavI8py
UMAfaN36cpDNrPlfbiB/zSuw0YZUfjbdv7S2Nxmd5U2k2ay38LN0jH0KA1RP4AxP
qyVek1D+ui1JRvXzzdqKCyYQVdD9DPfJ0ek96m4NSMHE7rEJgjbH6HZ9JGlob7Vv
5ZbkAtPBPS9tCmS2shRH6Nyt+cXTj64lJQTWP1B/KZ1QYPrFGXmbfNhdjh/w6TG4
xDwZ9RmDyBOypH/oaL6Pvr6the2+HBuSfS5cgaGmrsg2up5NZOihAFJt10SS+SHH
vtfTwhXt1s9ZMavlhzd9Wn4v0gDjYCtarPCbYystP6Ii96QDRt1RiCFc9RyMnlTZ
CXejtTeUa0wcBCYeae5x9/UZTElWr3BumCb58wP5RqYjfeMgPOzOX5Bwlyfho4xB
RV9ZNIsgq74SBSmcWlsU1BHyZHOWBT23Hmk5Hgtd5EyNQpAI2UJFO4iQpBC6qmp1
BOrHlLIfgd0UIdjbQ4tpH6qz6tFlFy2CzRkjUlG4qs1Om7zL0GzuE09Yku1YyPBw
GDjk2S7rjqiFiAmnJXpTNtwboTsAXIbuZKTVIgFQ7p3gwur5mv+Xwb0qEsG8ESIB
3A6CWGjcKKna562M0hIjbLy40UsT2TQTmaAOrkhGfAMOUwV3PrfpjaFajnvy200Y
yqzDODCaveDHGRnNWq2ErkMiOFqag0NNqF1of5iIGKsadTrBf5Ro3GU8iE06NqbM
TzDPrGwOT3Jc0JLOyFIXGxfAAUKys/vPo+pXWj8INcZzOV5aolBs7qsInbeb+Y/+
K/ick2Gn7Zv64tdSzOciTv3ST1l5kTiksYxn6e9gQcwnRxqo8VvUV4h5R1twac6o
/dPTsrYiuIFTTeIwT/a4mpSY1dzI8F3Xp2wYV4HhtJ+KJAlSpvvCfKJ1bmu43S6M
gdCLdyN1PLZatLSXuYvIu6Lw+b/trR2pXwFu5VARar8k+xzqeBVB8d4+y/QV48ff
IuC7YcePK+RPU4xf2730ST6h7o5RZERI1uRRlsqzmU3fbg7GnMnrrLi6YvELL9Ez
fvIzYbATmVejuJ+YGzKQM57fFICqodcsbw5D4Vq85mlQzsPlYtM3Ui6HZ2rDbS/T
Py456sEaydKCdjc6LhqxaQ4R6qrZ2hONCv3dwHS//JtxJp90mqpeMsfUWPfvvNrt
0VFo8OvdVzVomCqvGyjKM3BxGp65HFBCVif3j9BaschyA2tHYs0S0iiBkT1i2Qbg
Qq/4on8ZwhGk61WH2hT1GyPMjL6shyKF6+lZfjeN0ROTB1cwgybrvV8uPil7hh6p
jStz/FS+/tRQMZC8FUXPuo41lZhCx5yptN+yTXD+bSEh7frym16MwY3Dvk2th1Vw
78Emxyk4QJPOXvYHLL3Nff8B3oY3ctEs1DNvW2L5qae/KUnY1OieZmeaqnm9zWym
42Zrz9086siHzPqz1tZegscRPH+n+cCcKdFG/gnlYlozTwpBMndmEAJApgut+9IO
WkgUBycGRUDURcEq40dr595clKumRo//AqmqFlc0yaSulTC7WMgXOsYSbckf2v2z
YeJQ17xwdc2fKVKfb28+vounqegF2+E2NIrL5VWNv0InCn4Lp3PUxr39zgOoRUGC
T0os3DPLYByzDnpvhm1O7evx82eX+oNsxldUf/8TWhzMwBETu2E2Lk2LOg+jSkNL
lNrV5UZbaVwNGonUCCLtVggTIIdB7bmlXpaI6xWjjh2bK7ihpPx+OmzhHTxI4DKq
nCFGjxrGiaWDae1A54wwHAAEq08JVGRMu8seBHsf3HRncBIADtVAmhQJR42Safhw
ToQ23obMdor5HZqfF1NdXP9oPjxWVmbr/6bl1sv+VcDA+vHXeTPHOg8VMJyP+qbI
GblCvG3Eypkml7VL00hF6zrzsiGV+KkPixkcn5fzoRjHkI2eHoiLZBZydtnkjdIL
wqae3kh5lUnr7ej4vyUO4zRhPi65WJLZSOQM52cojQ2DkK7XewovhclHAnpyK1n+
3rv0IUJDBFDGVuM1SptNWL7iT0MV2kbvNTI6je5GkJk9avarwFwdJnPkMFZK89i6
31U2yKGC7fUM//gbLK8La65kGeM2g7M/0IHWWpOBDTX63ugPgLs4JvTg9++86sfY
dUSHfs4p1dr3pCOwoqEgVnPvdue5awE9h9MsyBKJ9CWQ3Kj0T00eaVw0bmS1gyOg
aAyq0wmMa+evc1VVUcSiaHU/xfdTbOECp6lof0pXH6sa2FLqnddPVyMnHRZIcYtN
iHk+9dWbTf0d8jmcf/JUjk1/sOo5yFwbcJpzmO6nvPkUKSBrSDsPzCySr+pVclti
ZyOpLzSigI8PFzg5GFmbJfnnpQiG3Eg+fUAXfC7mU1sWDx8sOEEEeAH/GvFK3Uv1
ZAlPl4mU/3hXbB8sMKxovdzJg2XU4NvJ5l28OOzlNT8M7B0TzwaK4/KnNXn47o6y
9Q40A8wE0nuitwYcxckS6W1QINqUJ8hq1qmquSqbN9xNH6rzzcCCJZTkD7GmO5ua
qM9lggbrELMo38BMJ6Mx3AXyz2Jr2chdjh6F8k4/GJZUz8t9uBp7pswnVgFKtf5k
asrK3SW+hwBrqMCATuvHdq3vdnTs8FAPaLMaxfkOpQyeEBjbkKk9QxvT4mKUA/Yk
MMYvSW/CUkFkZ/5jgP9fxNeT/lY68ORnApnfck8DKh0+98bomfwoRYnNUpj645OU
dS8iWdIEzPra+oqsNs/D2UGMcUtQhHgovZCp7Ceys1RVtO8ciLmd8g4BVBzWH2m4
lHzIdoyH4PKn6ZoMDRjlLK4lg+Wee6m0DP0pQ8wdy01Hq6cBEtlTKqH9nQk/2vzy
bZKgvj79wrBVK0sqiTpb8Hu6Z7xOPWgui0EspMbrByO/hpLSunTGlh9nPf53bKW1
0xl76HEkunwEFWHw8nHC9gjiIClQhYdajbRYiuzPZCJozI3HQZ/zxdXXItGNylML
hPqhInZRBdDABHWqZc2fOzulgnaX3CN8JpK3fHfxd2ijvin6VpZs44MDxWNig0M/
pVPstsv4g5s8R4HYOcVtt24DDeLT0uI5lSEiRId15IITFW+P9JQV3ZtOvjmDI45G
aQPU0CGj7h1fxk9LJWXn0YgQMftzNnpBAzY4L59nqzC1iG8BSDDB7OpD3P9WHlFp
QwVme2A6p3DySQPI45kd2Dd0e/rXrzUlnkOjFEkZd5iKxmFvKzRR4M/vD9laoupy
L/Odja/y9QS0YWrnM6PXda+iKCMPJPJfM1L7Yy/Duc3nnv0dwP1Yzasedet7LvZJ
S6JkqeKxBRXseJUCEId3Wca1yEXMQVAttGou/bx8w161Orr+gnthyh4va4+TS+xW
gY+CafzppOMU15/ergBi3Ph7kcklHwMr4GbpEqfYcXlfEjqhoWnqXRRfoCPwlFM1
rxkASTAvaGlbv142SWN0bO/Q6QkJ7Ke+wN/blF00pm1v5GQrFWNXMfH2PmVrV5jO
TW6QvSOPfWj0mJ/DII70anux9Vb6yYDYuAvtrSSpnsjo5FUfVZfsn0Xx4BN+rSME
V86XMchemypJ9tP7Q/65GiVIylktRslW4+dqYqCVcE+3yUgwDsvidmfJVwiK9YJz
Gf4LlPmVOi3GHb9zZ2aIXOu6rQINplI0pFWVk3QThRSnrDENhi3kJPAYl8S4wMXP
WRYFY//ecnEgi8H+Izfz9qRvU7stFHpYy+Sd9tEfwicoU4d0p6zGYZUtGGvxAaAE
lkBsRNTgf88RYkzdMPJcIrZNg6Tinq/O+Ki/lIIb8MR6Fp1F4EMn/z/w77XHJPel
JVUH4pGityzubZVkazB3TuMrAUj9YAKYuf4EL0BnOeFsOfn75o15yQY2Bl2qGgYI
Neke6zLZ+PB9UkYfdj1OiRrXQeJC29CH/mdWMXlhWStiqTG6DBUcNjT5ag9+v6GA
49pViGKHGPhY3NsJqf4GomRS9OXshba5xo6cPLxMGD1PT3zIvvrG99in4lM9hIgq
MT7nZ/gruiA0IqU5WnFVx2rD83jrmPPzxZF2tr1fP2kYTzGigAA0tnONq5qW/NJT
z6hsNdpn9JdgcgNxLBKXUn5niVvV3hrK878W9W7SFXzTx3lMnibF/SpEaAa2LfgS
d17wZW5e4WgYhosbDPzmL3hdNQLFtZbuA1hFLVCin7zoXYR9zIRnU6uq3bUzbpa2
YBywj0cezlo433frPUmiRY9sdPkFA3tWv8UzSUauqFXaFTokCMwk9DYGf+vDE8cr
OwBnn1aG7Xr3BChL58me+1kSqu+0fzLTzqUFFYmxZBEv3yP7uFD/2Tx9INm/p8Q3
aQr4NyEsBnoE3v3z98/hPVTreAVRwNmTxMo90h/6L3mfwjR7+F58mDmI8FLZr/Uf
LfmGQ39FmB8xVvZPxrAc5OQZIqpkoRpL0mf0gGcmBSsEbbnD/4S+dX1mqcGyWgvf
VGhtQ5Ss9lyas7uv2P/Q4Q6entxAwAhkak9rUlPfKG8x4rDvvw6TtMl42ofVVxi8
KLnmdD4f81EDbIlYu3V2s7Cm/CUKCWY2oijTjPEAVZxsQBPdgadzgEbykwoxNfGQ
9Z38PmyrE7VhHlnYpLJh4g1Tsx3cBdnw9NgdIlhS2xwB/KQ6l2mJZ8SGqPnoZ1th
x2zrmhXRNFn1qZg9lc1J4bxL/P2h4DpNu7YmgOMss/RFZe2E7Vmu7OMYPU4x2APe
CSCXeGlpdG5mxt87O2itOajTk4gGfZmHew1ssh2bAfvhQdMNHj1v1jOlrCFNb6FH
05Y9Q3hTrfkeCchPEDA0jg7PX2AUMk3Z6JL2RCdCzT0q1GwQSbL8buG7DThlD0ob
xHzw5bL1jAfLfj6BMnaWdVa/rdP3XlZSckSgY+SZaVB0/Fs0vPoclFb7BAjdZk+m
G7GP9werRAkvUmYrc3vgP0deX27X7fwZzz6tOnguZAn5bA9fTpEiX0OYNUmxmCgC
85PeT3jmNZxlejwbdPv7oS93o4wn7EvQ7SqVnhQKz6VZIjr+ClgxajzKtz2xhUE+
lH4DOPPUqwFdesGI7f/cv6xKV+NqVJuj7CQVddcJlvM5feRtMHpfDc7Lu2NQ6fsp
09LukguJ3SM1LVWZcRO0EzItUljYWOm+fMkiA23Ho+UlOLLeki+JEQnBUhRm+m3G
V9TnRFJDfx6Cz6HmY0Y3Hc5S0pjvcH7idOCu9xAqH8IFLYgDOS2NXAkynMG0bw3Y
VcczMYiMePQXwg0YN4Hbr5k7hbx7AFifOSTgOBpRht07SowreYEDQ5jGfJsRbWTY
VIlJL3SrA1wJuC9twQyISwR3sQWE6+AwER6FhNEf80ZRb72tRZ31y0PJOCwIQotH
g0zsj47v5GRmunYS5r9b1p0bA5YQOZ00tExZwVO4AGx7nwXoPCrJCxu7D5A4/a1v
8nTFha5bjXssaXRw++fn3bScKbQ+uxYM/pq22EcbZ9Q1txS3d4w+FomuY6YRurm8
Ipsv146vQoEPZeUkx5QeiKz0v6yrjC/hfasSTtChgSq17ZWZdygJ/8mg7bHKc7C6
v8HyXr1kLlDF1RsMBDyfJmd9XTt1uD9J8H6UgQMJoi9pbTbK3q8Y8pmqorTSB6x9
xHl2VZe9V631G4TIa9YT/+Ejm0cPuhHJPiBzLFWb6R+5dn/XOb/1R4oONc/qjiWU
82kcuBZq1qlmh+iuV/ix0441j3LGf0m4yc5/L+Re9mw0ScGHXNoovxg/vXrnqXrk
Kwhnsq+HdAsXea88d8vhHBT2ADgReD+5iNlN+k5HMHSw04hU4f/JhBwmhsUYLFgG
klauIJE5T8LGbY6a3lCkylJwT5VOiLR1Yegip3LA9/9JO7SazX9F/ay/NdsknE3u
/GqXLXDWg+30m/mfKWXA/92h0ix5AhiUQsYcnuzQ4uxGRrqClqjNm3nOJabHxv1t
rFXRtZhDejJamuQiBfw+F/hpWGV7GocBcPabRl8vcFQGjd5nmbnDp6Ds4WGjvf5o
pcFUJkdNz2f4yH+bOwyzkR2Jr491d1lMhwKWPBa53r9TC4H+aSjW1U1jB6AaC7b8
QJuQGnUIhN6gmwmdJbe9vMkshkqQ+NSKoHfjfJiBMJXntxPmyNDhwxx0X/QzXC4R
DmE8c5/pVCYL9iMHWQ/j8//G4a0ZeYx/uvGKgR//aeKYhx0PlV6hYH2twm8ewl4D
UWdUzew2LHvZalevCcZ2Pofe5k5DFCvB6F94wXymnVY5JpsWUiPJQpMlx82CruDS
zeNnCuOe0pbm8pS340BQMt0LM9SjiKXraebDVQ51VgJlO48el1RD7tNxhI4Buk6H
xrbdOzIsp7eye0unMCoBhO0EhUTEVALgCnbdqIrjG8q1QM/q/FkLC8EuUnx2f8n4
T1I4S9b1AtVnWJX42AOZIIv5xiAuMTi3AYI7kN7PPfTrzWyqMwytE+c+os/1BNQM
1nXza6tDrg7j/s/CWoK8/g8yC1FG3U0NjCH1YL/UylIIOtusYr6onl1EGOP8npSn
Q1Nmpj/NvYvhQwX+0pDUD6EDDbbjVBJR4oMHisGwZLYPWJFGiMewkO9p2tPXqgzV
fHOK9LU3NchJ18gioYeT7eIyak5nCYzXS4WEkyrzwiJQ5aPRTQEDdW3gyOOI2vMA
hP7fGZ4b5Ev1J95tiGfOcl3Xl5BoOewjr0r6sSOP7mnSc0ORZyIMe2K+aZOwq06e
as3smwoq0BLgXz2AHTj+9onfKuXUpQtooTBxR4/KuZorxolWFfu0I4NP671CsLwp
uo8MzmuNPfV+NVATVpYOJr9+hD4MCebd7iDW7wApZB13lbDsjUFUOTblXEehxabH
nJ9ZhD2civARuTUo272ozMC+P0YOimUhzK0YH32AWQUaKJmWRpVN5BUBw24tKjNC
7G6SG1RZXcT4q7zsDoRg/WBaVvZof1UZm4EH8VQ8aCY4GoKFgo3+DaaWA8gIvtcc
7mAdZhIouwGsx3+w7pcXR3ZVinVLyxSt3gO2A3Sl0ECVox1zvU9WzbNP92oJb+qe
FIm5O7XUyh4KC3nk9OiphvMD3c3p5/KzvpuBoDU3jl11Ad2L48SLfANYemFTj90A
MKPzYXTyOHo6EDQSJPWCrqaYkcxDqu3RsP9HcAenDW2CnUTFv0UaeTBcHdGH94zD
Xldyiyg5tW5gKimK4P6h5Sz3InH8qYassTJKLejM4hs9DMxXsURTY5QnLpIOs18F
sTkWo5My5ukz6p4DgrjUQohEdZkBZoRDH/zFgTtyPlkYcI15nVOElKVT+0vrfZ/c
wxLRA2b0V6SEiuFYGu3gDkO8VHKtMalBjr+z6NE2W0YxnYxmHzt504J3wrTkR+NV
LxzAB85uKgSsVoHfAKoOEkAOCZvFbDLP7OnQOObzqAOIxL8IKchB87LIBVQOGb95
ovuuLclFrol7nLIyIO2+BN2Xw1uEbTAdH/7gShLZ0gKWcroWOTuTChF2+DqIT8eQ
+HqYmrFCWLX3yKrKwEbS4TUI3BH6j6nn06VmpSIakGXEC+Ql3sK40uRUcYbNYgvo
G1i0zy5yC1ozjh2fJqWRXycqQSYKzrqFWMmdYd5Pz9+bGeRygRu3FV8cpggqw0RE
slbMBgxc6zqfWaLPP6bZ0zXSWhQnuB1z2jrsf55KyaG67QiznEdw5lFOVlikP/v5
IzkGhLr9KWmaRMkEDMCYvNHwlNRkO+pVBGVQDnsgiYgcDDsPy9A5Bpxri26KEQEm
5ZBHX6MGjnOwqVgHH3fusHVU7XVBGaVIV0/SAMBIEgOQct7iSV7o0eaBtxENBw27
s4vom0XrWLOHOvBEXR6A+lFZrU1nvsM9wQC4yQGC3H2mm1ENr1Jf+o0dEE+rpoRc
CQF/krEX0iPZusbomS9ODJh76w7MNbkBqGoXT121XoUAxr3FJG+jjd6H1812HQK0
dWsUJ9ULnJUIJJ+s4kGBTsGLCTzqyx6dYjWGopPRYzx51w/WC745lVPQy3BNMVxI
yawnyVO43epLDLKKRxPWxHziXYy8Jz2VYJxePt5ULIsO3/HY09hdUHqPNJGNirda
tNll06v1wdyAx9cZ/xaHrvXcFxJkR1++pJZUHuO4lCUjMNu13f/CdIZtlRT0wc7X
u/dtYkatHXFi9jYuo4vVDUj1AJSMi6HXY0ekGh+RxGfDqKs8mXumucAktcn9ZyTv
4pHanyEtsUQvS/6yWsZ+WXCOyPMiNyqSyFrOxHg0zdkoUM1EYXU0Oor92N0TR3Nt
3+yu78r0DPyrIAd/6r03F+H3DHc728dKTIHDPSLWRg8DkLnwYxAsta5b+LDluSkO
z5llghAUyhdUjJJpE9+o58+fJZcOoFtcnWUz7HnHwoWTIFVZD+PYt8Vo3ybjEaE8
65dlYQNOTL9aaQKALw7dHn6KxZ7vPZjv+mWL2w/1AMdZJTY8oPZ3HIDWR7uEvMeJ
1B0nKwsH3FE6I90bjTNcUbIIMdfyUcTLyiOH9IuA5iNOp+XBNwr8zpoeLHCX2iY0
4pvVXitK/MysVKUx3dQZgqMz319oVfE6RMLmJDMTnXJreCyOL7BUiwBYleF61sSi
6AQ9+EeFMsqChMnBZ7++bQgeBs5Rvt8OBmAkQ1piUde0Mr4PSbG19whetO1dKzA6
vHT4/svSamafVuo0jBy+nO3JXXRMzto6pzY5dl46ADXZE7g06WlraXHHZ5Xq5ZxB
Zv5uiWvFfdXV+mXZSPHu00UZGl1MiGphm4RdYvss9YMdyGHrnThVmdjTOUZpJfbO
4Nh2ym3QaQPf3PMB/vZHm2nOs+8GsVXR5vGNhG9KE5SrbrS3Ot3Z65SzCIDwlpJb
1YxqU97hKhvY7Jc1TLKSnfG/+YK5pSBqpvY0GzKw+LknvHiykb5XzCe/0rFa7aF1
HWLWK/u9yI9MSbuRXzVRiQweErYg5PdLNP9KrWZFYlABrjYY8IZffYJsSti96dHJ
2I+Xt35OabrDtmH42ZQ9s76h0A0QqPNY8aNyD90JKM1bYgc7L5N+kP7I8Txocrp/
EtPWAUBedIP8xFA1kC75r0um0jpbqK5j7/+SOa86kFX0Z0XEZ86vQ3Ah52QvPkd+
ljfDBd9c+m+q9PLoyZgc8jn4l1NvOER2vocsooVZiSWcbH9A0AkrSA5vFMalnAHl
EfW58PO/RzAv5BJLf1BRKEJGEYXc1LD02Swp7lUFQ59YEYN4E8wsSPgS/TbNhVJA
U7utGFvsgRVXz8BIcHtKEoO9JD8I5t29D0PlffykoCWP+JSNrrX1uFkYGYCx0ajJ
+384Agykcx3+Ms6C/EIi+zBjBAHUXeKs6mfoyyGGffo6Dw511yQicdA/OqMX9ox1
HiKmWlzRcscWHb/037/XgKv/PdEkvHFz6/M1qEduZmsKdH75RXM1NaxHHnrEMSDI
WM8IL0sAG6/DO1DoASUeA9SvhwLWLNbVuPOeEofRsGB9ZgGl9X2l35V4ODqD0ceY
ouPvdVtUoM1sNbkkRu1C/gSv2UH7lqFyznpBmy3P3Zx6vGMfXQHp0rP6doagJhFM
mHuHvqx8YNAXeJt/GqaOr4gb5UZRdP6xyIB+kIHyvl78xQaaxfSx8lAemMPIkjwE
8KxRYEeJQAiWgAy1GCNG0RbcQJXuHYOZCWG0QE5P4buHTcW5IHDqjb7wbCbaJ8AB
5jZZryFCHLqIwyE0rxvWHfS4luo3cr3B67jMIk2pqHZ3X+jLtYJX2AX9StzU0XeX
CNH7CAEjqedi4KO3XGxNwvheNRB/bPiFnz1msDOt+ZsbgwVFTFD2u2mM7qRY1A8+
xM+yCVVJivxgmK+c1gnFMm3k+8EfEpKdaJSSSX1i419G170arI6WHpAznmQTyMOa
HHOXjxiEfam16O0Az18Y99JuGWxwYdwOkZTWBq7XLYI3XgYJUn3z88EDgqfrYLI0
plN4AOzAA7inRgQDKcu2fEIAKE9dkYh+vuFE+TXqmb7vJSkGnVNG+VaZGUrkprgT
UFkMgv4Gpjnl/+PQa538LdgBk+V42VYl6owhr3lfMOpBU1E4bqRDVyDDQ5yBcDYZ
a2cOdY9WB5oMtIbmvmSmFH06eRrteSgp6hPaMDSyJq25N7TKHxVKfpoqfoJz8+xf
xAYngqJwKF2plAbOwHwYrA4OOWbkm2rSIg3W0NHRtwpRX5RAZye6WxMKMmdhDm5S
lXoC4SoA0iyzh/9wWemFBtbqhEa9xmnCQcj6hjkrBVX/Voj60sE/7J4+IgSnXKaW
YVLW5guwcmoiucEtAp/KqBANRT7pIj8Sov36lTLTPQUf3QTaMecOiOUoQm2Hck90
xE1qHQpUGHlMQ0g86fMBrkXUqXBKXFOI+mNPCtVjfXSljzs+wcuXeGzc/lWlkVMZ
eaY9kG3oNAx5UNg5djGKAh5NhoFd2TL8vWnK4qxvxqQRwtOsc2DIS0jAVLr+H3Lk
0mV6Azge+KNjnm/yZk/W1iqSd4oVr5pEWMf9ia0JwaZtOizxOBSMkpwmngrh0wb1
/xObDovzfl3NATM047RRYhYV6aA6WVyhcPKDqwtp4ITUXfNpQx5mL0mEwwY+vy+X
Wx72WCOESBC9wJ7cVd+Ufc6NvPIbSqk2Z5BmWq1Ei2MwPoq8RNQzx2KXXqtZXL3c
Q/uiikOKC6sjkHqDPz+xisTGH3/271BBxKnSHzkAcAKBfyvxG/zoIvdb0BHGgkm3
uf7HNV8HdGgNZXm4Jttw649THEjM0WyBtmoA92PlipqhU/VT8khbfoj9qIz+Yyhq
OozJFsLkUWWiNlEC938g4DEkGmXfgYnsFCcH63nLrESVujbht3rOredyJaD5pnyw
3niNiM/+8Z4+/akO/eTpfLDVZD8GumqYcw6u01MdcbMNxgKETpkiNo8DrmSvVPaf
c/kUfoqpOF2POyyDR8udRjcY/b5/Y1EUkbO25TbSHIF6A2oZf6d3oBYQN8Uy3Fos
sa3uV0PpahoIgBVunzhxWguckKvDamdifB56gG5yoHVXisIHhFqVy9O5PQ+viwbO
ABahSuTTnQ6fKVjgtGB3crus/iDVWTk4bPuPJILrrUmOavqErvOgSx1fQSqrDMkh
S19PvTwi9Nl0i92fjCSixU+opM2UqIw4G2UKLo2vGFz9Dd+5O6M1FBxz+nzq9n+E
6AWrE/YGmvFzgLiBuCtCIGC+Ds1qUJGmPnAa6GhceLMzNh5lO5XC/R5DdFWrGqW5
TT32l03/Hap44cgggVqaHG7t+B6IovvEayA62cKnh+jV7RngzjUy57S/QYiHCyxQ
BOP9b4jRNtesIBe66N9t6Shes2T0yeb9nMJH8bkJcaK5nT7M7Jba6uTNaEx7P5lC
yycnBBeC8Lzm4RAZWz764ec7x+B4FNxR8B0JVbzS7jF8GjVLMlakMXNMETii3QVS
wUqNJCuf0oitZXR7i6VBlmHaPTY7I8M64jwTTUpp5cLvHE4mTQiz0L18IZpAV/yu
RVgKyKcozWt3JLZ2GAECJT5j2aTb/G82QG70E3ezUgQD4mfAGz2nw3SGW9FxUYXE
txNjaIUdolL18HAOCU/7gJM7mgRdI5D8C8dj9Kb7ep/yOZhbj6dJ6T94+AtiQL4D
goBpW22Zz9kEWcuyR/nkiNFM+7YrNkJ+QvOCfHp5EvxCFZHSXZXRQsbVtPKbFhMi
7hSYXDEYVnTJyWlModQZRLMagIT0pJ5PKQFEKUFEHQzfj+ZmQfVPf/7BeBNqaqdz
OK1rbLv1pApw+Am3Jk8iR9CKc6adfaD0yKJRJe3ZE1CZMFIeqSNc4t8XSkMV6jhh
euKOEd2i9wAe59qfYKt/j/NBqdQ+fYRI7hkyMUYgSwWOiWmGR2BgxNfglFtRjKJz
GMOdjSX1mU2LX5toADH1zT1E+GD/5vMlVchwssy0A9uHa9oo/Cq/b90Sz8uZ//Oq
JCC9dUkWxpN0Mc35RxAMAtSU+dJiZa8GmMJRccDdtOOqkeom9jKOhFrrL5axFOmn
G0q7QwKtTwB20JWFy9eZU2PQALIdcb+bRGXNPI6z/2ou1yIrqqHmIbbS/ME9OY79
3tBJpxxPF+4zjp/An27NOf4M7SDmUSJ2RM7tF8hgRKIh4l+EShQCd/2EzZbtSyb0
IUadqGDE9xfy3RlcUB5Uki7dv1J+QV1mjY6hIXLrqovw52PwMKaTklWU0HyZ3+ac
SyxxQQLWLxhmmjmVftynDwildPIBlgs41n8i7YtM4OvJnLzvn9zrSZOl6STdCHQJ
SBEy6Ic6fZpRT++CFHh2qX9KZDVXe80QaN8f92CylELXOoo2UyO3CqhJeiiPbN2Z
M9CDsHMRa6/jQCAlfV3dXSpvO84c8HM0EYI3DgWaVHmV7URLll7M5VA8zG1d2i/3
QXdGhLmzmqqrVIEBrRvyjVXfEVx2ISyucVLpg4Qq0+ZV5b5LPEJJZLFWZy9f9iFu
WUVp6QlTVEpjVQqkWY7grQx8dkJRVtdiZymKuxWkfqLYBcFipIGVWmuyyYUKarTZ
5aEH3B+V99Jv8KIppGvXyu+ll87LfxQd5iKZ7C+d4ZK2yJks4M0Q+TWLn3tPXlAO
yGO7hlzzn0Y/BUtbH65046ceunupy5kQ4AqRc0yXvQRLHvdcJcp96P1pbbW1T/qN
bLUFJpdj0ZzR0FuwVT1/bIMPknL/o9yU+vhLM8bhzUHceUfN0jxcOQgUP4aV4tNG
1JYrI2fV1fwJgvXwEM7qlb9JfhiK2uGJIRUu53i4k9GWnwNJ3sanp8Af82zJQfNA
asvRKOi9moBLzkvO1zB4f2Ypb+N+VsZkbZ/FEWUgh4UKqodt6RaK86VX6ZjdcZCY
T+WsNz5i1p15clhc3PG8rnkJhWD9fRaO5nHfwAhWj3z2NSxXVdHZ/+YS2BsTkFon
dldVDQJiCfCNbuCzfRGbtpY9vLwY/vqIoY/895DHSJayCfHTOLvWAW8L0N79UzPV
XSBDz9emo7CMO08+3LoPx9gzfoiornvoKb3uqQ/2ViQ6kLE1qF3kibBn8sgKzLmj
sGicEti5CpVTBji+a10uOIiJ5Xc2XHFna60rDKDu9kDk+elgj35G/VcZ+ksjqCY6
BYtC5dl5GR/2OYBNJwdBhIipEweHlyB/6WZTW1IWd301NhgbXwzqE3/iKKBKTF3B
WeF3/1hdN3sD0MkNQtp6dkfB2uV5+0R7HafJCEHZQsbLkbGM0wB5hC7cX95ogqco
RaR70iWWrR6/HhlN53pjtoK/ddp7o99v+4DH3QxUBJ1PxH19mMnNKwY7hRbZvMet
COTw86oyq78hrx1QFWiEcOoH3BcZ97ioJb99LwRXgGzzH/zgFUScCckLjqwIvOQi
/HN1e9YyMk1/cMZNz9BTS25zpw20TAAkcr8uK4TGyVLQMtw8OKv4XsU9MIa8zlxD
MWuzbv/vfw0tRXbLaMOUvDlDk2W2NReg7CQ93eAEo7pYRlu1cLuK8xFkV+z9DOlo
dMWNGopvNu48SSohwJKk4QJ+XsJ4D7Li76iuNDdh60ka1Kb3VP98IenN9FTmRpQ7
Yq0RhFtRDUmmUSUchPE3spmbYuAE4vV1WoMmvXGfhz5Zt9DBIJasUFZbmWhE8a2L
wxw0NIs5QJr7J0Bb95tOT79sOEpOsNtMWjiSm6RbuUn446Bo1IOKT17aO2+cNDHu
y+pTEYHSeLSBzng/wRzkTf1WmWElzN1TuXVGdUqevq5+JsuY7qyaJn8G6cGPiYnZ
bjMFO6yGqhAc3XI63g1Y8/yLoPW3x4hd4wIs0Vt96EZSPpWBmBtrwzkp351Rl/jR
xwhffksD7Af4+Fx35bQI6b/tnvW9c5KsrZLT0W4Iq0ze5n/V9NNNxngWFaU5I12d
8p8OrVRl7WzMJIzIM9c53+3ZQIBK/6fAIMa+J+wykug8HKQIsJkjrZVJOqPRQHxT
JFM63ZXXeMEyOvVDyyqpYf0rJrALvTLh4r6Gq5efiej6NPaBDT/ejVVHH471/oBX
npmm27iTytE0UNKg0vVFlIMDcYfoDBQKkp6RCj8La12RtC0JYZyb/zZgwNON6ElE
ArbGhDccntTFrDI/bOhOq01sBg7p3jTZf3zF+gUoYKGxpnI9N0xIxoI3Sok0GrDO
jbMl2F1QPhQu1apCWKO9CVzXNMxXxl+O11+YsUZgMpTcRcRAUGIwlqMYKHBofSkb
HM347kuAeN6T0/y5uImbc/p9LV3X8BYuHiBVm1aDil+6syW8Khb2p1iWKLvvxeon
Up1pr8l8UT8c1YkwQWkijXg80o/A9OcBwAYqKlZprpdS7Ap8ddY3WGiqjY+xxxDL
BJpw81060huCCKDAOPf6aVT8Zb75kmDvCEK7mzQ5dBppjPhX/K84lVLqxVGJ3jxT
6Tts9kUJJnXp5KddjYM4OHfqxyATEJ5uwoQ8IQSmp+ZLfpso/e9PnmN/2cLd35VX
zZlsK2t7WqA+F9QQKQvnfjR8wQLiOPd8D6BQg9XZLctV+juBnNVcoXTk57OQuDFP
ill16KevejVbagFvCave5MBS4mZjiCWD2XwvDfu5oNXcVMVIZGnIXF9m8ZIIrZ8h
S1FOLRpzy68/OsAtzQgVkkB8Zf0+NGCJ07B1PE+n6n7czpY70pzmT2L9f1hj1qgc
VJHYQNNgGYrmd3qRPvGyjELChdU6XzWfF+YlecqiwP5BPhjJvymdxNXaS8ZFAegS
SyR6AVQTQhazmTsjx8xjvQxYwGfQ0dPP3KRvDd1EcCJWSsYNhNpTLaAqZJ5iySVh
XHDaHYdpaK9jtRqz3Wbse2wEz55T1BtwiGbG0UbuD2E9nVo0GvkQp+K70/FvQFnk
eP7QYLpVCgRGbT5p7vtfMIodwbVJ7M3D0G39j6f3wNbpE1/Fzp2RjNdyfBP4+lPl
oh/zdJm9Th6AoFvY68wrqicl+OnragDSpEv/sVALJZz4rNGOX6faCXxru8hohBrE
NGzlp+LjzNu525oyJm/3D6DeD/+cNbSA2dVHrAA41/FjOL4tEcWoggaoP93KdcF7
O/L1H5I6VbCpje5NElo1UFzdSDdUcwAndzDqZRgY0uKgKLlWnU4vjslGCWWCIJ11
toG9pBWIUgSfa5nSdJivxRZVxUCvWG2jIJRSTby0rjvQNLdqecQb+q2hVm21K6JZ
6AgB1zXadHi5/m/UfrS1I59n1Wbfkqss5e+7pSkgHVjJDutPXJ1D9jVEevm1ZCAf
NEUmtCcw32yEsqWT6UZFdneqBg7ngVTmi17pTs9U/aWKLlTBoSk3kKyAVl1ftDo1
bZ4MCHSsRUiOdshgVd6EQNtPqAqhOIjWmTuLAIhE6drkV0rYBm7Bx49p8hOHQdql
9/f96w0yWTV5t4fZmoZTsHgZ3jR64ofidwIJPnFgmWJyQHNuRrp6q4bpOtpk6tgf
57aY57DEsWuSeXjjEGCWfXoLqGayX3YSjQqa4Afl8UjxCD95gHI6Iy4RGDVkpHI6
5syYkx8VeQZGeR7IYh+ZIqBWwMALbiIVlyeYbOn/CnMTMYMM85dbK7bKpnWKdiCE
t7/5vbzRBxIs+JBlKT9boYydewAC2J1/XVKajhKce2h1YRQcnxsKUmDOPGA4JCaA
WwIWOqJcIXLR3+N3m3Ig+55nGuNFLUTiAIR1nxtaM5Ro4AoFx+6njJruf1rKNgQH
wXYhwsc/3q3cyoXbM7hWSjmjMNcSmjM0qDOTf0TLKjvl+6Yu+LsSslfUMcpHC17a
9vzMqjq7AVTFveX2b6C9ZeirRWkquYn7YCUTyq6yTTAQOnudtmp+MizC8Ng/XHpS
HhPQp9py3A/T1M4KzkyPJkfC/+2T5c9sm7Q8bqLtz5omF++SbY8eyP3AkbSBOhHM
NI4aBKWp4Or45592Bez/FqDeSK/2YghWWgIiyvOTtKkzVGzCkvOvwn5gTKVZdYRB
Z6852d24SRGIQGi6Lg38u4pm8JF5e49b/3T8Bdti1SWiOA9rxikSNb5khoCt3EkB
B1z0dnKuHz6WEg3TURR3aiFNxrupRPjK2eDz0nmnq9CC/wBAyFfQ1xM2EAOK4hsp
1rI7MUPwHOQESruh4IqngyQnHtvs39g6usBO9d1JyUljFQLd02KNFHXBNrB0vRi/
rrE2OrHpvPIIZlO3Y3UahPG6t11BdADqFSZVHUz7I/OkTF/0gd551DeZPe2zr+3h
r/VTwNnpmk1vhJkN+85qX1GOIXjRajuAkaUAk29q2Vlt0IPVNbg6HEwsK9egb1Oq
DaB818ibb62k52CESGAa/qkLIZxtrGKrSF9Wq+KVYB9eLOK9h+b1QZ5zCF0qXqPk
L2I6Gbc0RgDfYQFPS6CCrn3wWhltC4oMaxEtdilChP0WGaaQRSt5BMI/xGn7uVF6
QhBbXM+qXaNg6xXEMlaGgOQ0O+qqn2RIq3+uo1lTlB+lVlZmuV0UcEZz2U98bfRx
B8cb7CieTX/+nNYR+nYe/YoiLg0OaE+nAz3QKfNLhccvxZbBW1ubIt40OG03UnYf
JaWvFzFTOOZBy+TodWFuHwKh0hVAi5V1ePovX9GytmcZHtHhLFrUUakcvYHgWuSo
PQ/vTvmJrQ5ry8wRcIknvVmb0p/8BjDVs/s1WfgERewtB/tXSEt06S6TWZ7PBpk8
aNum/VOa4XVkfO7YAKblI4wpDO2fEG5rktqy56j+Z8i0nuuU+oHzkOOmW2s1hQqo
7pC0aO8MKsQ28aoeW5a/VLdO2Vx/G7CGrurUzDeaeZ9D571ITgSXmYaRSckCh8Dh
/+KcBsZR/Y70pFA23Vn9ErJFb19e9y56l9u1UvCjhdGAwvXF+KN7upTiQ3wxPfwV
bq2csae+mQ6SJYhzi51tQC7HbF5T2KYldOs1Qd1xK7TjKH4lOfMqwbKCktV/okJo
2hMKrjM4U2v/YOyKRYqu3ThpdttV3uLXm0XeWhbgNYbe8JycvGOw6g3yath3oU2i
fAad4Ri9J5+qIleVSAY+2pyk4OC+89RPEKsQpI3lFAqpuPxN7V6+LCzOula1lDbm
BbfmByuiU1W7vM7iAx8EMqb0HUtM/FR3OOUdXDZifj763DYKAtMXPovA+eRT/QGQ
p3L9HxxcqSle0CYNwSOgdj5GHPA7xo/HnZjmam6w7Nb7XoVuQn085/d/mlB03o72
7xZS+ULwx1YBPgKwSbUFph1VinMB2V5jte7v+5xfUQVtUQICQM29WeCT1PdKsqVe
EED0CCkOHRaokOAzK8+85KLvQ3hc8sgrdgMET39AkzDVfum3cgaT41fvMRecmirx
QZfgWiYhp2N51ni2Uyo6/BTQt9H32MTBpTjH2YawZ3C2+VO5NpPPEAysTJQ2V+pO
UyyfV0nxSXECVcO7QrCezVGiJFEVGAdlr56BO60ne4N4MT2+zKljl1uEe2DyuebG
V0ARxJ7RzITutKO1YStiEyAyowKPJ37h+ALtjS+Lu73YpVuMnubflDl2qzuxrv7P
nb1c/l0PAa3DsH/e95OrUpJp2ADKXzQlaC9K+MuWVyBCleFqYWY7AYT6wQewZgFS
rRL+CyC4fqYI8BYQZR4P97lcz1+JP18J9e9CxM894cWxeAw0/qH5qIP0m1y8dSyw
IMrPbw8824w8eb6Mp+k3lka6f6cR2iX0kw8P3bIOowIcTS/tOSnvnAVe0xComsDo
VTttQ685pUnt5K8DBRY/t+RuKSpvDbTvvi2BQkIjNcq44ylF75Pz+qemQs18XX+w
vcw2rzDKVRi7gWXLiDVFscvkkaUeo4KmiQaN1NwLsYnD8zysjOEuw7F5SYFrNCT4
OuBVymHdVRS8ASTVgfzHXECQqDAusa4b7gBEHDV8ABBj7nKWd+0MozNf9w3XOEuK
V4HiMUBIXJ9vRax7YZuSIViolTeJzSIyRu13xVJ7gpDT+Bb82Nhm/GsoQA7J2rDv
RLGzVUhj/KTORByOFdPGpcM/XJI0G0EJd3iVrRmwNvK6EbewjRknhhPO22q/7bO5
DlgOc7qqqNutyIsdkR7bC/YDs3V1RwAKJbg2qCeiad4IY1G8vxzF1ijDlUJ5EDnu
RlLatiC9KiK6IbMIH3hM3Pz4Xs9hhSQnZ/E7TzPzgXb5nr0s9sNNrYvo36CKQhLa
N9u43R85CMduAXOwtZ3JaMvfuc6/HmlRkCgHGpDd97G1yIYREgcQ0Xy64rgGvHYe
6byRKH3p8MRsRraoTrl+WQTrfyZ9n2dni6y4X6SiQwfeMhfF44APWuCVpIYSEMj/
IV1njaID4duGUXB2kZO5khTYR8A2Ojh1Fe07epJqnS6z8b2nPzm3mjfvJD+l3ztM
dPjo0IOp7+PA9M+zUbqOkC8BCmQJq/SkBR04epOZpcCA2QCYfWNVFTAs/etgyIc8
uKKeh/8uFVOu5QOY/jb2XociAgCpbo9x8G6BGcdsd+3chymmHuYywXN5xNKsXlbG
pEwjEaStRcJx9Jq5ubEWVHkHsuKIcdKhXYMCZ5Dvr/fm+ubVVjVMiq4orLeJBdUg
guftCD6ZiyK6DHjkc37PsS7qbvIwXsu3Pdk84dbYo498W+QD5bPvemBsMaAQBhfB
Cx49oJY+xS1AZIj+ZOpP2BIiWrHuIQsiilH69So7krGLbFNiU9szgm/3xwkCrHcZ
EwSMRghxfa1F0amGJAOKp/LfDf+iJqaeu255rum1TkbqDZrr5ukkcUszJuiNWvV3
OmSA7oItnSs/zip0Ba5+OTNRoGfiNtfPRiP+7FrUJSR4i2RyuDpc1STqWBAYqswM
ux7hm5Jgkr2AI8Te9ui/cVXdu+0KI1Jk4qjycFKIe21DHiGxnYfWDfnUKOJr4FG2
LRY27G9r6p1y5VWi7M0ZaBg5Yq7IuTbJqRhgGSSD/G3yKCJYYVMWvysjj8RGoHIH
fjIel4fRB17VPuQ2EJx5A6AhPnkwebviIYG/DL0nbly5dGK4sz1930aTNCLdumjy
laWwLuoJCMZRa+lauJro7PcuM364xZDRnwe3yQhWB1qLG7fexNjIft6Cwnrmrc1+
3o/cXoltbW+XgF/2SHFMDDAwGMX0F2nIirMdk8qO5Of6IAY6O7tCfwdK5APvn/D9
SkrXo1SJQeg1rKBUj4w5hp6AR/u+lshBX4mOXHpYNN13S2uKmS0Q/tKuv3Ri0vAw
cw1M0lbKA11aLGKPgzrwHnWOCdXuim7aVjGKYmFm7hsRNKLrE0VpF+SFdF0E2MIO
XxY3TixjS1VTH741o1U1+MBBSq60rx6QiJLNFnnJVCA22cNOAJrA6Cj0g0kbP/qz
AaTrV+9pOGnxMBzrcWSsMnn0ASObz2oyPoPmj7tlAmf7CfsZef3T7qlwgMrIY2x/
SXNd5EJ+xIHNeHREUUcefl6x0vhOyAYRc6CR6PY1jl9WtWtwSRO1u4+c7Ir2xvmG
ewmWe4R95LD0NgBe/ZdQ9tPcadU3jEoiO1nq0lPHdupf46gw8sLkvD1O0lZUq7nK
S4Xn3v9AU1hY8yonqPtWq+JpKMdBv9J0RWN4nhzG+l0auC1oz1sOznU43e0OxeX/
X0/zEV6JknOfACEN6epUVFCzBNJpWjin0JvEhL40p/yIniA58noXGjgRqpVyVor8
v+9r2gOyZQak/doxKH2M6tiFvXhP3xNyqTzCojYqJTVTIPrtL04xnO4rtXkMeEA+
35UDQr5xIEMpw4gh8TKLYwXi4vmnxhrHKjPAsW/FL6zIoKnFa0vqRVMCYzox4ICs
TYmGmiGrYEoc6HkuiCYm+umRjjV/9c5YiQZZoXWJZMzxe2h2IqnNtePXqcogMcVL
svJHcpbHghJ4nEM/RXXyAXZXa3T5qVvE2K4UPwgG5JVv/yghVLPCPyHExaM6DiNt
ee2qMovNY5J3IFwqw7hRMiPyVN1R9eRwP2Nk60s05hay1Vyfzb0Rrym2C+7jt4jN
hdbwr7H3vBjtgL46hyQ+DMDnoitAcxkA3mJkhtDGCsgAqtb48b8cImtzAbtvnG+l
0Ykm1WwmmdowC8FwvaVmFj6HHWK+mCBaTbBtNzfe0buIUZN43HCk/bxmBHvGpFdD
FXO0JRfdKrO1nR2sFoExm30oNwwZX5uDnf11CNLd37Ga1RBmNjw0q81zxz/uQkv6
wYVLBQ+QHygzsgJfwysju4PSLnZBHTq58QXJhL13EA30vPrJQywMquFqmmkJblmF
FM0wntT6asui7gUgETH8a/Zv2CHw2ZsQhlx/s3eaQwJkWnLUgijWdSz+/5/xh5tK
9ctrV0yQ7rup3FDZft4pEY9jhJHJXi1d73xRRUmMlI2dFObeyWzc1gaG93zUZ908
1C1ltEYIAX+Na9rcNW8+ZwhaBugxPdxmCcmhKFERYY47NzgvzVkzLZL0oWP8sELN
mkSpSKiYjSSTk2G6qYbNdQvzUZOA2SjpOBJuUk7491eZDenwxzF0gxcAmDfDN8K+
Vo1H53GUpD0Ou2Xdm7L8kASeyspuYCKOBnxnDzlclQ4QAl8SB3lZtkNM1zphhEJP
o+9QGpMezVcFj74CKeuHCn/fBiL0bU0NuUaMribI21z1XfxNOPWrBThwtZq5REgx
DRIDK7hq/qxAbpJzy6qTrMp1BS7u60GVmXXmelKUAS2LpJnAa9+7KNbJPrw3rVTV
4bSoUKRECiLFxV1LlG7lhqjbG6WwTrlrT3YYuQxlH6pmbsZZm/WKWL/iYPo9BM/m
qA0ox5fi2LTnMA5KytcH2CLn6bAQpqHDv6iwzstUime4vrmvj4MnWLs/0b0i8ynx
3xHvu2m62iV7R9D7pZbFRed2jolkdy8/YuYJKcsBZlzbeMpvIvh+SPnpeBoM8A2v
LH7ttVvTkRbVZ0PT7rrWDgUx327/XSPabN/JtUtmVfSN8gP8jwZ/I3xbHGGTFOHv
d1ai7Y7rfb4bn6uvjSZNqAEjMdhQmOXrEOM7SO2XZx1IZw6HSXYAygHByjJ2dzyr
wwISfK6QHotztfcO6IswbrjmiL00OOb2n/x7kTx6T9WuoN6DKynHo4gF0RzbwYsY
7YglLt4Wxct1nW3yD19wS33gd/370/Jw8rXjDlIutbEFVxKCW9qUlZHFyf9sSxxR
GUJl+x5gp7hsKRrnbJ1v7deOtD90Ko7nqIQQ6+pMGzngpf+mLZ2ol6+ouahU8/76
Kd/VK+p1J1e0ZieOaMp9qYGujODNHnCteCFKWnnK4Stf9trqcjURLiz5JbqAypgP
RCmIvt26GSFY/IlQYArhqw2z/mTFWW0x5lJATmRYuy+ZtxRuJBuWyclhELv4Ih6B
CrB29asV/eDqKv8jM/kRAtbLv+kj6xDNEN004MPhV91Dl9INmVoj3ctqIc4Ty9XG
3s2F9VtRy/JeRjPRZy6Ahtj9rTc0lIttQMszkZYFcqf5nEsDf5nOMcgflDEXQj+I
1t+ebmWIfHLBtF1N8NCD0hzPNO4yFRZcM5IlRLb6d1ydGLQ8/xpisNL8Mz4nEkoE
7xitD8mSKEVRoB9Y4YNQiKLNV5PLXkcp/edoUN+IKDjyj6+6gAKfMrWzt+W9E5kE
qxcvnAD4RtrOZIym6DWWkhElSXTuAwEOCB9eauNJmXn7GkfKt3rj2XvBnRS0r1uH
FUNbJcpRjmAsLDW3sDJ+Ro2rPkxrvPsXpakVkcRgmT9KkdFJTgy/wSx56EtP1LSY
uUqN8efCK6EGD2tLPmOrblnazV9cxq1Elmo3Ud+C/Boyc2qyfHHkaJFhcNfHZs3q
6xaRlFbW+cmgbqKMbLXg2nZkYRXq7ukTK7FpTGDRycv96kcNqZ/0Q5NJKvW3kVwt
aQLarwRGCUVqfYuodEzzPEHxp8rmygHw3EqqSMYHi+rGatoAdncd4TOJBKKHAzU0
jSrpPARXo0K5prGMoVdkG1GRoI+doCeCw3QSmDjZlmN4y20zb7PZ0mb4tNjkH4kx
ZSInRVkqSt4Zet8LQ/13KTxkwMAIqDeD5oXgETLB7uRVH87Cs03ZjvOVSWLVvpVk
4HOCpeGlG4dcVLEPXOEWk1zF9e+O/scMyTYwNlnRrMDo6FQh0Y7r/E0UY2x0buJt
8V21GoOhPx6jt7zV6whk0TCtpEE8a1aGA4S/5Bvj/3FaBZKdBf2+qU73pFgxlWzC
VT7yCGLPtojqw6lBH9xdnnGW3PspcS+3KfNiXYDDaElOEKbL049Fl0p4awNPoA14
498oQ7HdrCpbHiwVPWCo+t8c5QmWWlnVt+L5Lax1F3fysXGvzraG0Qgk150StmcJ
be7XjlfsUSqxeUH7duFwAcNcApFVW6ay+RDw9jSk7ZTSHiCY6aF51dp9kO4S3r48
lgwNJFzxjAiwDExkoOsld+JYyL5LVMyiIn+WZdOjEoXf4ubcGt2NamMavjzFbtXK
fZkDIWQzqfX2UBHuhG3CrHhdvjkeKvMVZSC5IHc6HvL6D7gLnBKRdOj2Jp0tf+Is
S/zj9OYFOiEfwI1G86B6jIOCXjB86nWizQs6yBijKOWnuidD9QywI4GUkjLb5SBy
6x2EMYNHfRQobpQfg3klHeYLUTKNZkz+QMcNQDFiz3YZ9yUDNcuxvEafGznywxgH
aFQpZDKo5YpDK5zM3mqRVAyK7UnV6Hzgsdgi75OCGCfuU5b3SWA2LoYrnZ4h4p6M
0gl5EXR+D6Gplj2WgRtVTh89LdLYSZ+2Vznt4XLzSe2IHt0q3iVYwXS56zchHnAD
Nckcdj77g70RWhf+nn9CJthgne5GDFbqGmr+z0akBTAkh/LEa6ktSmAobYXR7cq/
XhIXN9YMqlGWkb3s++B7wg54AlsSfbkq9YmrhOAS81jYBrVZyAdEQTnuBOqc23wN
upqGNQNqKjU5AlhBZ4Q/iuCVX0FbUTWfl2W7yundRNffvFOnpGmX/MTwh6ORjtCv
B6J8k7e3sGjiCX/9KaDPcfDooctxgHFejZOJx06avKAD1MYqWXwJbCdhfszjfc0J
O+QcMSk6jA430H+4wf0iatPv+XLZDIMAwPL0uHURDs2lhBHpJ5yW06VzWj3OH0Rw
zP5CLNpPx5uZ+35wunw+QpbN+FgNG7TqvP5Lbf/nk+J/7ozYL/r6hxn0m3ItkeQO
LGRA1ja0Hnp5tlWIPeO/h/VAGeTeOxBQArq+1b3K78C/3yE3dqsjIVcn4yS4FOwo
DIAmwurQLGS7gIjqG4IwUjUyHH+udrPTkNG6CF7941TkrGHE7HJwnCGwOGXPYwXm
ptI6y//z4SBUqM9m2fs0nOtXoNqeRdOWhWFr4kCqmCQp+OwfV6SInibDSuBri6WH
w+rrdmmb2Wtnf8chKAt+N1zxtNqFAxlg+cv/lYuvl+qFwQRdApEDhPY0tZ40Mi0A
C4x2Z4EGi5XEk4vODn9L63yAr+gwMUE40yDd/s5nU27dXN9TqwlDV5tzah1oJOs0
E2I9XK1J2qpRQdzkf0m3ETYDK4ichY5+npVohmo/FmPM+lyoQqPYxHSdwkzCAB5w
IUO2sd/tlNujlkEG7dOd2Gi0AD49q837KQqa4R7tVnT4CNIgfdOzM+67ukK1Exv9
QnRxCibJZ1oZ/A0/WYSUs3Xp0os2ok/v5jPO/iUQx1rqMYX3VfzCoq5wdrkn18nG
rXA4Bfkf5mF3P0G4xurRFXRxbVH/vcwquivqNZkGcRKCHrD8ATAX9hTT54vvtG52
TiazwODcK6KZ0e0yzJ7IiCF8eWJSrG1Qw4zL55nKPZ04NujKM+L9wzukwRZE2DJq
sq5VgygMzcCvz+LSEJPYV3gWBwVulqW66OIVMAxYyQSrtwOPzeYNTG/LCLGZFJkn
SZfYVPN/j/Z6wR5UVRxFigJUnupMRnBOaENBvIUjQdgj8AnlAjG+o12yx/dqUrm8
UrY/wpfXE9elzxQhaAFHGBuZVTLoKhUsKETX8O7VJ1oKeWX5LDlRQg+Qcpkm1BHa
n5Ac/BFXaJM5AhV5KeTesSJtZgrjEKvFTWqBNW1QFF7cONzfk5IkkxQyOv/mEeim
J+GT5YLVl5SMXIJssmajbBlm5XbuU0+bWQegHQrYRx682sL2wxGBsHjizJUJmscd
NJjnqqHor0YIkyBEWUYjwLAXclTO0QHQzqY66roZZlD8RP6azA0Rf1lKDRERA50i
rLIWG/DD4GjQYWuMHzW0A7MDkd4xNWk6fRem4iqBFnjZfG/GNRXzocqHbjhPoWGb
hc2Jas6c1Vc0OBTQL6X3R+IRnfdiNR1oNemtR0oULxEb6cr8XEGTDpgJ2iXh8RmY
p3QuWq2YVuySENki5fIYllQdmu6N7N3H69D4l0i2uTCxzQNn2uAT+75CVr7W3y8V
nzgHPpMw4R5CFkQdQBc3XEKDH2UaLYvrIuJwA2B5TS1NeqOGwBg/t+VDEjqDHGA2
4ijxEqhO7Y5+yULN/FC2IHOnokaEyK69pvFfwrjqA0TeV4hgDhS1Vrapw3/PaB58
VRDfH2XyutmJ23TZyu0H6a+hI/QxZEK0cJGe2pZFE+HBYGAu54QLE8bdxPNjxydc
YTExsr/pvFcIoeXQGCwEx8woyu7Ykfmx84SSdrSTmDJdGzuQiJ6ZF/bBh8tuF/fJ
XX/H0Gsp4lFjrbRwUTdpfyIgQFWK111hDD7x28TU6wDlrF1SWFTW0ANBKp4AJkjx
YegA03vOiLOPVAY64gl6hA0EKRRMZgDkmzNNomRvaavuQUTEnlF/2GHdiVxi6QU9
osXMtlhN2MrzZ5c1NpGHkbDatdniirrm5/p5Ujrq4tI37HEJtmElNNIOXgj3bPPe
DYN6DWUKzJlEwpXR8u5qNwRtH/6qVyPufPybSBCREowKy7dA77ggB9nD9DBpvHUt
ituLTuaEOV0mEjxQTqiqnIkfv6xALYrweFDGXVhRdiAo4S2u50JRZhNVAyc9PrGU
8ZBZBBWhc0XVopei4BujhX+6YHd/gTjOuc7WYkEL6ZGkp9Q285qTIp54PWa6CtTF
T487vmzssyWedZ2vA5nUDPzvOuTietBL6shn7yL0/lmQOQVGKViyPqns5oscCKnc
n0f1u21t5Op8I4dL4ZCVeDnw256zOKcNBkg8hueGHg404zcE3CGfJlmWRZIE5PqJ
EeHvkrzurIWmcijZ9/ywbvcWDNoDWfFA1qLTyrQodrdRN+UK2jx/5MBst+Cxi8TZ
jEY+gL7TNSDAi+7hLvdz3uj+RUX2m1dUII6GBa8md1yUa7Ddu7a1s4PcE/CRu4ea
pZlqMT3775OIwvfDVMDBqYMlHeJMg0h8ojd1h2AwZfXtYnDYFXhCm4KowwrAqDWz
9wNlwN0N1sD9HW4KzrFp9kvcWrBs7w+r2ljLBlvV6/SILh+Q96WjgUMqlNNXaBO3
4VDrF5LXjRIN1XzILZoY60YVymPUpifPcnkUtNzrH4vNSFhmRhvllKbgmWm5CUuN
gxCjGIsqNQPFJoUnd6bjlyhOg2Gbs2s1PL1SwOn4reJMz/0kDkD9PNTBYGYRYXxt
MbVrVfq5uLiC0FXFmvCK6wMnhHgmZgDmMsdbSHkEtIaX3m4kBwIcufnOiflH8dZy
0puIzqcCKs98KZNwkxpP18hOEYYU91yyiHMLqz93Ik/j7bSzrTSu5JU3t6v/OYH8
IcjuGzgucbD4d8kqmM1SU5t0DLU3OfJS6sMH85kNW464+qUDRKInpPkNN9B+uPje
MoOHa242yCYx/WyYA54p790yLWE0DBXPP503Tbvaq956PKau3mIUeRK+Xv2X8tGr
negm6Vjp1LnjNZXAJP7FX2upYcxdXjGoJAaphBi5Jx5E/VkqtuMNo42UxLlJmSaF
5fxh8gyaoV1D3os4XaxBkWmtTmRo2MPGXiHR8q1ie2lm63YeUpncT7wOvuQR45BN
hkgUiZIF3RA7WlBLX0sSJsvFzU5h5Y9qimjqmswsTJeKwcZRWUOVnpoIpQlL/BLi
OxHZSyORD/v2tEXRsZ5grFQq+b0HRHkLboeAsSTVe8XA3uTJErylrMLgZfvZQewb
CpRz0ycfc1SP4kqHRM4sZPsG1LvyK51bgwlRd27J/397g4pnQ/TbUev3HR2MS4c8
glh9rOK/9versDBaAkI+huDlFmo7INhLlUL8Xp/e9qT7idAfeHwtqQOHPDLj3ubS
N5SLvNdr25EkRWWhhD2gqxRH6fwXmviQuMcu0JGrJ9v7NPy0pckie0ySkELrNlVp
tYVUvQVfqv/LUv3s26xVYA7xcVldiC7tRZ7eTDwRZgzjqZ7nRTxx93Qcc4UpxXXi
P+SFMUeFS2L4iyuHNOjQ1oAwslDMPfGT/XR23cSRTSc0qKZ5d3AIEXE/3ilBH8Z0
pZrBbSid91xALPXdGYs+cDEGy+W3jnJxEk7J/bFhQ1jb9jTSCFVN4yCIqFrhkl0s
7LeNL3klV1/+HYGY3L5dbrzmBkj6EPPRowMhR1h2uK1FpbV/g2kBPO+P0HGaedEI
agy14WjnVWh/Q9gvcIO/p8lWR7L/UV9+16xdiPUNbI0V44K/ccLxoGQHyA06kb0w
JKOs+TDYD9NLjh7S5+vflrk++pgeRUOe1eaJ1K5F+ZtUNknZflPFut2ECMUP5QbE
mpGuGFCd81MgDIfjVqfYCLD23JUKa89wqQGof/u7LAmCwu0h7ztpvP6FaSPiZRb1
ydn0OI6/iPjYNvsj/P1Ii7U4ZYTtdl3RteY+8AectGkNQF+WniRSO2xq4b7ioIO0
tC0f/UuHAbOHQWFMU/DFMnKdZjy4U1rcXN5WJUwTC0tBW6usfL9GKeYISelmDieo
YCK1kitiut6BzkmY1GJ2bler/7ASm6x2+DajFHMDRyrR6NXswfrwheTSdCg7js73
/ugdtHORFiWwgYVEIUL95e54ygjcgHnqHNYcvtGiv0ehNgSRrFZg49xOEBv3wMgu
LyWJQEXNBE3DBn7dXNVC5r2rB/pfVRzhxrkuqP8dAAjBd+w1I8mjhApb13zHyGYU
h39gCbg2qF8V07om6sDYZsIlSGZos6NzcKEl6tgYWuBWDddtQfgudx4T8+u5HhA6
tZ6bAcJDK2I01G0H9GDa6dXWaRFVfmCqttLgWaGuZmkcAXNnUsfKnEFcmMhsD6KU
ly/zUzL+fqB97/WPar7AGfcOVsNsuOqirzkTXMu5uRLU/hglVgzeGft9IA8VdqE+
w79oSRHdFn1dbjeI5xd39qk6IYwR5rL/FInTDbeso7fgeKJHhSC/M9McNYKLUeoY
T4I2Tmz18wDbZ3dwZFNcFlqVuXZd8UG65CKuysi3uXSAex/4dy6jjE+tmgXHX3GA
fAR/J18rrz+txwJczENmti4RWL2Agpp60VYmbxljH3QL14B65f53z45BLUYP9Ngp
U5PVRaz4ba/V7xR6LMhBFvVTi2g6Zoj1eQ7gZbfXNSNicUHWpIMVRSAtlgxxLt4N
aHIyBkJCiPJNIU0KMwzRzqmxy9ZDLppSfaBqg6oQiayUxoA4Azck3BviIQ7BcBIi
bUCrt5zbeFBL10oCdFATZRJkl8lwToNBRGGAa7kUHnaAH26bFqAuXvqCPXXtgT2Z
zMD6rww52qnOR+nv134TuHuYART5Pn2ticMfT7dV2UGAdcYl08WUnz4itM6ykQuw
7vOYh/UH8UT8nDQJViXaWrq/yJoW15Ke7JF7coXeeNIpnJ7KlcowFshVFouTGiZt
ZKRC6nTOIri00NrKV2Ad2IcwWrAq/sv+CRfBcfHvzAysVa6Tqm76Iicz0Oz+wRAA
8crYl1xdXguY0YU2KYBCtsDNLt8PUm9VZNHyaSsafTNIs1n5fauvHtiCm/cciY9e
eLGiYqlrHEC1tsLOcTrppLwVBdUgHaNLH9XWG8sf/CWaEoOt/39rWZnkycSz6A1f
VDIlfks7s9FVrwPHsj9I4ffanTQx930pak/S6fz0scRhWbI86+iLm8jFRDnVuoed
Vh1cC7kh2heLCmEpkhKg6ODCUmFFMgdtSkC//xithDYjfsqzr9u1ejMo3DsVwF7s
ugVPz7FrMREyDg9rw/mjYRBD3nREVS40wIvwLQb29FbmDdokzJYEwcY69/8uqeVp
uroECJ16n4Gn5bSpOsljTEx70PJ9eOKeoKRJe0Jq/pHRvYff92pl5yRRex0bwEJx
S70kYyI8MWSu1f/24xbWBEIcYh6fdChIMXOGDvEdKjsq5KbLkMpllnCJ61BUpNX0
hc2aaiE7HwaRV6ANPgtxwDM7Na1dcntgTmePI1iCmWJfIy0UfjMw9syi6e+yrvCr
OiKmoragf1wz8JSzWjsG3iO5PjiiZjnL5jrRVnOAaqldQ/WpVK+alQ3mlxUwK93u
fJNBZCoHe8IpFaqUjPHKoB9XCQa4ucVZhA78D7cvtAhjuCwsUtMmT7IcZhWAJqED
4tIeVp9NxUYNXGfGBOzPDvODBrRdK8oqIJoucWDBPHGrf0k+IKZKYkq5eiNgZuQF
ASfPMHMYmZndR5jsUumPbU07Yy9vKu/ZPr2/hagaRJ4Wmmnj+26IdAnyQZ3ROJcH
EDmQGqesrYVlU/SZAxMYhqiGsxPZzJpVhdLicGVjuBxdht5XIopMJuXpLhtCw7vp
z3G/S/hKF+It61x06rAK6J5aVA0+J40dKE0OFNZ8ZpxgDVfV3HpMGlw0kVaHq7rO
BCxuKAB2425z9qjQYiz4bHyzXq1XYXOXw+OLDQuDlY/f8P3evKJQyOgLmQu5QJx9
VpuJb93kEeCVww+F0Fv7bFuPmEB3xcs6oRncHCSpflK0dZCIZNAIulEK5AudYVTD
WYGSW2E1sle0v6a7YjHVV3SLoqbLmLIhuEtjT2zaCmvMM0iWYWC5SPp9/Snh+2en
KMDzZ6HjJQ/BAb9wPviH+d6hShlzoRpklUuu9uU5xxeTPd97A9wTywB0axmlWCbv
Y3nbZgsxGxuZlYb+f2QVh71eQC1oaDhIKIzOgZQiH2DLvV4avsZwGPrs2nRL9J74
oq3m0pALSKI+mmmvW2YL7wrBA8rjp0doPqHME6zSoOD7RWDi5msxaP08xciFV6YK
bqe2//+frxSNutHf80y7DyC6mkH/7A/UYjeMcHbzxlI5BtcBLQD7zJyALQcnNEJy
y5dpMIXsRjaJZoichtq1OqsMGCFXXsg4bdUWdEkzdbZMe7nRb1XjPmFOpLVZJ0E2
Vu3LvXIxtbg+GIplemypGDOU7t24t6ujuwr+2NV6cRBRNhoOkh4/FJ0EmTUgHMd/
nBOWc0F2vDozSWSuO82+ZvG/XuHb2tbWFgs8FzgAYt2MkQVkjoZJH0FdX1yZpU1S
Y7jkGU1fYpMu+jzjPsBmkso8Gq4vQ9iYGX6y8tWNo3Lg3VpDl85Syqkutxprt55N
tX1oZeV4bklB9zqnzGoe+acsYafik3IWUB8o7U6lvpkOYmQO6qvDFkr5JKjdW8B4
LA57z0mJiPNshxQhpR0n/ITE38Jk5pVCoIEeDutZksIFQmH6Hj/rhLcnwCLlcoHK
wRPJO1LshbB/rFTfkj+Pe/KZlq2lrKcbTzojg4gmg7a1oY90Q0ziljQhJcH/B8lM
k7onnXYyK9cPuy3hbnkw5plkQVjQ8DV6WFG7m7xe4+IRbMDhBIwZe33bhcK3of2h
kzypS1kF65lML5IaDhzJUnmgP7WkmISzkaeQNPlkQBGnm4YXnAv7SY6/ZS351WI2
b/bytjCYOiFuiwEljkUlpKCR0XeUxwhJNYw21MLMpn4R3qNeOZGBy8aLVnFscWF8
eQLRaQkynAnQZSVOB8Pk0BiV/+dApKJUhxGf4UA6z/Dztvl/DF8hoTkbwoKLjqiP
THvCQVCE//OlRrrA5P5ILWYB8bpJ9gR11K/u/lnUkMVq5hzQROvIqMt9EpBMc0Rc
J1BDwUZ70rYGBuYBVtv6VpCWekxcOJrQv1cScrmiVteyN2MyIaOhKG/gMnF/OJru
wGdYKDeDsueTfq/f83nRMOl7qTt0AuDc1Abtc4YTVzpApO6+zcEvbAL+jueirr0O
/ESe6SkO2yJdd4/VcqpIUSHSc3vefh1XZrLOL0w5PWQ84uuTKBC7v+ggD1InHbgj
HRiZGHx7lB3GHZu6KQwaTPuat5z5ThVrdLsZMyNtVPCkpP3nHoE0xbKYuwEU/acI
fA1BZ6/lOL2Ka6JwfNNxHSL9nCBQ+48OJoXAiImaXgCfzk3htVHHil130+ovn7et
mXGxoEFjIV3nUNveuQSvW5EqAzPVQ0VhP2Eqldi4ecMOV+7F9gAk6fbeHwciovgF
4EBQdMmEOwBDRnhG3xCgdt1oADrv85/3gJR3zKaAq2AslTAStmDwDHt/holwwYEK
StblJxv3Ch6qPzC/7gNarGQmWEP96FqCjgWQ9RB1EMnnTwBAwTQ/ZQ58w9LWS9kB
GtbiAuHochcplKP8Fqh4O8HNe7/e8YV6wYmuIgb2cDUuFo68qpH/EuF5QtkviBtA
jgbCAnzj5xmO7lzXrD/Wpy1CQCs5FOypMzg4t6Cmh5wvUzznHE+95uAyVoEHdQWh
LcDKGE5xmKxKO4RoCO6xY4sdaT6aWWzYLyRzYOo7ZHoYouz4e/aT76JKs41zdF6k
EEZY3c/xyONNqdXZzArYUpYCtPKN3UokFr6r5kSc16OkFrdnZmOjQ+A1fLUZQjER
OGm6CccDDga2Atta/Gq91ewbOzBV9XcCbBmaOUc4d5bEM0evic6Tx47JmdvOZTsZ
IxqyeLyJIXZ+U6yBV3l+YTyOLqYyC/obk+qFgeSyDaOjTxhvJaMDjk5Xeb8pRjU7
lsxgNnaHIOLbytaLFoasfp9IdQOM7WG5Pkod3O205q4nNlGrnQi9HZLDmUUTRRO2
1S+R6/AHVMklM1vv4zGSa9DP81sEJJJ3ulKQVJtZxuZJGgRFA/91hBXQDW2s9VZj
9HtC7JMJ1J/FGyqCyv6BD10Jf0K2PXmGhJOXpMFxF8ZsscGcji22OiMjyJ/nQpVS
9NkYylMjhzzRMqvOJo+UVE5EDGUMePcrBifechnQSO2WXrd9UnKzc0UBkl3fZT6V
OXHvv3O9RVkQQLtWmnBRBdYHRSS8xvc/7ky9r6FdYqPd4ruS2YMsKqU1fxyA52y3
9NJSyc80XgDy626Y7aDbEUgCMSfP2u2lsxYLbVgaDHodZi3eJiJy7OtmPGA8iojg
IXW+0yJx/rn1RLXclqdHQvndS/O1ujhAit6N7BMMdM20bGhB5CmYcOw8eaa6YojY
BsQ/NAmlyUbxiCL9q2xeTFDu/bCUnEuZ0rvbETt1S2oktXdtVcuJ8aLGk/2lzJE4
WxAXJAyWOgmQHgvNqpvVLbbyl4RuDouAccJfs+bE1be9Q0923oNgWsMs+5CL9xPC
6hu3n8Nn1k0ckGN6MHHq9PmfVHWDorQB23QVrgBb9xC1LCb6ACq4J2itaKH1zsh3
NK/TuYKwtcWrHIk44+CMa2or2a6qHvAmacm/OdFQxtMRI/tkL5f+qX24UnpJtb09
2Y6hJumkDLEmK6KOGD/tTwTVZUFfSmtGfCJN6HoImQ1f0BSg0Jvp5OkClXmtL6HD
t5yxtQpy7vPMLdM977Srd6iqASY8prUJ1HPliXnM3QOvLVCLfyiadoDGBJd55P5j
B9h8yfeGKfb1SzvIhKE5ZPoNghZEqIfBmje6ACOzMcD1pHP9RlfqCOdtu/x39Xpg
MYqCTztjS23YqQBVTajzQkj0EZFdVJfjcD/eZfKPN0zKiK0h1hpBAE4oAxCDV0Wh
4M/TKg76y2KMOULp8iwz3zDgUe4KFdaiGwY5qmYjB6SCZDfEe8NUd5o+PGpXEbVq
EuM+IZBDicfHq5ogZqDgVkUgfHu99pXJyVM7Vdwri1vgn3fyvaPi7kUOKM7Pnprx
ljYzUm/+GaF95fVLH3o2GL8+ITh5nGOgU69r1jTIyS7Jx8R17jpRRvKU8YQqD78p
CoAalAa85tZ57X+4ddYba/zEv7CWOFHtBlu66TLJR9EiTx7XU7xUIc+z4qco5iI/
hwvTMQdIZnh5z4WRngOX8muxR5jC7Iq0pWMeahdS8yxp9NzvZWN+inzH3ADsw4jt
2h3O4zb4Dj5AstTx7GKuZgauR5AtvEGsZgrrhItgJj5RTtbiNuQDgkOnLy+Vuoo+
jwmXaeasLnNg14Kgl3TBUlQhGBwEaAMrAFZcyFXyiLswJDCllWTJLmr2mdsESH6q
WedH+NoahMZagLCXgxzSoJkqFiEqRLwS1sXuLxGrIrvi6NOzCf8QxszC/CYA9ynZ
d48YiZWgoNLCg92iQCMubc95Bq+BQr6vaBOtdaKY8rQqc0+77w+DSTf4KdrnTdyJ
I7mHXc3ADnz8F9ALZdM/jvUgRAwFl4dV9Pvl3wTdkzq6idq3YreTG+hn60fAHl0O
80YkL/QwVWzwTfminotPZ63XpZMBYNtON/Eu9Re2HQmxqyVWqnjO2ZRF2gmc98DO
IlcfqCjIyRvSfs6uiotN578F96FOZlc5MRZJ+oFPhklMEKTiemNFvtlBBfKZA+Iu
gX1Nabcus5RuNExDhVNEl0amL8BL4Kcku4rMRpntrubfFAvXdmerp37NLQ3hi/W3
sQZauO1gjfM96+vO1ZlcNa3KGSYEb6aPrbS2sKeUO7rR79Vtw9e4Sv7+hunp62Bg
0Oxa74gHKC3sAt/PH7e2XMVT8dRDXcLi1Evu5FD71ADBwHomaI66CA5rv3ZWzntl
r4NsE4qDL4VmooVQ6cAK88hr1N5+sBKHz1bM/saxv6LsvJaZ34lmTabcs0Faa88t
ZMPcRl2ahTR+TZ9zeWbTTQPaUVSHX97XHTV91aHEt3ZPp1MFw9Ibt6fT9nO/eEzn
sG0z4FlVH0lbol8t5fztzHqwyeC8JUROnnjD6B9aU3tFmhssy/YhrZB7HjtWxN4V
o7ZT0jPIm2rqozgFL/Mz8gIYussBpEZ5XPmFjs5cUEkZRGrzbDA4gvu4NJh8duoW
Wr5oGkgSfMvR+Et8E7WCHVp+d4muOfT+TK7mfRpUoSGnKw/JlNua/x+3G7NVDw8T
YUjG14AkFv6SCX3lLICNRm07s9+fIqUOQ7GpU4F/vVcUHuLsXsomfBE7lU5Ln36e
cVxo/igGRySvnNlytzhWntwvB/f16tMWIaQLmRgLsVxFgZDmUYJhwhVGVSzc2yH0
lX5z54vApNtrpRLvh/Ue2c1reSwdIVIPOSirvXJ5/YCoDTt6H10YVZB+oGoY+jmG
3cmfTjPJdLmFKsTteH0uQgJLfuCnmOZqLmECDlOTR/NDTbVnzOeu1WxDav/0DoBX
2I3QMX++n7JGQIpUzkO2TjGWaGxCMF6GVyb+EyqB2sabhRZkZjdfcSRWe78EeZVG
A5Wk5TrZTe/BZaDqsriVrSs5DnYIhC0CcEGRnIldq5iXurKAwF6cv5+Z1rcXCpN6
wFE5S5oGyu4YVuE/ADHH1vLsz6NjqLxygCzZYtitagP79NWLa/1Dk8yuKJ/bnVcD
no37T/wLWCtuIyK1Gaj7HCruDks4mpZevdW8v0JeMMCJqHSXj9Mo0rbthmrkxQ7w
t7qzEWMMuTDSsF57SuN5DPTs6gGWbh5HG+MMEucbfTPqShwpZejbWinXhQn7XESS
hH1SLZ9TkQ5b1Lvtcd2JGB9kQCBBswBHTP0RAQDFHYqP+TtaJMJeUFYEPnx00nsC
6lCwsYQQceSiNhJJEUpn1QI9FOvfBTp+UfaFo6BNfr4lTt3x05Rv3ayekvy4a82K
DUyeEr+rxEGYb4kwO1iTtkQa2tazI330qgM06BWH/iqsRIgRA8CmoCRge1X4/tv6
bWZFz87v3G9LE7OTqcKMEkvxXkYWzRm2DWP5BsKHbFbuED14FvTPEPigYDAVGk+o
KdD5MV5u8X49IH2XVBvs/kCGZAbxxEBES/psBoJV1/D8FE+bHqxz7EK2O+EGUOkw
AsNWTBih85gf/m8iV2mTJcqxuIHr5ly7R66kq4k3WjfQJS/xmtJeSlHH1HenAqMv
97hnC4Z8JgtGH8ccxvg7WxMcAxGFZHeQezqV+l4CIQpLZbHGZtOwr/xkawR/Bwu4
1BYWIVc9wxA71Y5XyWKBLrgUnaj79DwH2f9o69B+Om/J+duiKCQz1Ltu1qOy8deT
XxnkpIN0A8YACXvZMKQs6JtM8edXoFWQTCUHRBYd7YJZYsTnxOGfMnVU8WFEpSoJ
/39FdbTjTEJ49EUOSGA7afP/bBD0wmW2+pNeVIT1H9s6Ss9MqSr+6TtzLU8JbbwH
6jPMN5LIJxSI6+z+HLKeYOu4YRjI9v6e3wgqrxfoi+Vd8s6AtDzSxtZCDJboyfzd
9vMgo0mudD+W3KSBxIz4OezkQ74g5oImUymKO+6b7NUZGIYgV20esBuZK7GNcxG7
+nEsQwpxsRqmcY1HEk26/mzgoU/XSGx0lVLtp9tg6SpnYjKkZ9GfU8Ni1EmBBmNL
l5CP8s6Df+lEIN14JijJVtdmURIG03UrSpDM4VeIYR2IG05mfaF9L7Wx5Mhzdc59
JYThu3oZBIXdqfxu/tspIac5Ab5YOardxBoWPqWG7vce+dW3zp8SdXSAZPL8jcd/
9HZUNnIvclEeHK0ldATrpFmMxMPKKHTPsea5Kum2UKiBphLzRmqhzmkmKxv2IsKy
V0FWFG8sceohV72rG8gpqF7LT7ajtUu7qYdhYZztwjgrDIgDnKk52gczV/Y9h12U
TpIW7+13ndHHrWd20y6aKIWpcQgbmNW+Kw0le2q1TLD8WJiXscW3u5ojjTD6m7kf
+7zu52dJyWWUFDMLal2Kr1BMpfOfK2bftztM42lrLHEYnUQ+P8DCmAUnN1KPMQgv
cgSR9XZw6Aaed6CG+UTNclcynIvTzcM4p1r79zuKGBSCpCj+DP/ms8C/cH0eLm1r
embfrCysstRv14LKVZQt2T3+ruEK0LYRA03/DPrHKevaL8aPLK8mRlT3hg38YSFh
m7db5EoTv0evJs6ak1tVGoKiQRaOs4qCEp4eCAHEpMn0/46Ule+Ycn+5LIyy0jQX
wPJ9/EYzWtKNVt0NTmtnbIneYNRayM96iMmcl/GFfBoZh4uXsgqvaDuuFwL1CBds
4oYwZn3rLGyTBX+ljncnGSRya5Cv2Kee+R7rPzs4Hr/4LoCqCkRf8aj/J9KBv3qj
vXZ0RodABeL1YeGy0r+rhZr3l+SOLYytZ7fViBYoY9pjz+M9Ycqt6BvZjlHhhMM3
EidubhnWV+j7XGRGRa8LSMJcRK9xUs2TqUj/Wcr6XT8d7bSgr1Iw0aZ6zqoEWSek
CCS/B5LJ9FwfXtoXkpNi3SNsxk2D2yBANZrUqwubpF56XxvxaQ5eBb+jJZB0HQQG
YHlh70tvk6z9kMPhhuUMNypHaNxMqAD0D+di/9M4jtBcCeP4TA9/qRoZYDdybakj
4baQKiLJvUsJEoAzVnFWIZ8bdOP7uQ5UjvRD+UmsEMsKuNYs0OKqb3W87WcqlG4U
ijkW4qwDNafM4YNqDz72VwcA9V6vutqXPjioN5gzfQeI9vPjChAigT3enQoujXWV
zcGAC9OSd8C9rP860CYxI2JnZ2bxHCDY4gStytZ36rPh1FB++cjs5PFrLQ1TAdOZ
gzsmUuE8M9PCXAu2Akf2yfBWL68v24MQAH8HBjctLsKKnALj0fkg0WLCoWfl/Llk
nRG9JzBw0+HY3YSPQi1Q1w2AxiQ7eH8zVW1h8tbBcx8a4DeQ0qeRaNhdI8MNU4Sv
N0ewwPHQuQYLw4pRMVcbfqgKyyXEYR9AToR0qysEqpXHdzBLCa83ijlr0G8JJNiJ
zzl3uXIOrDztnLgtHbjXCsqb/1husMgAc+fMlSDlnDVGBsgh6Tk5dToodgUFJ9tq
AHNIGsrKKM1zKJ0uial2opp3mBDPUQVsnW9VLwwLAZd4PUCmRIr3mFUbMKoq2NHE
Ycvr/IVSHKw83LQsJz0CE7TuV5sjrum8Xj6bcwnDP1GoIT7pI8tKdMXe48AQ5dAi
oWRItKfU3u6LR+4Iwm/BpNGfzBD1sysVF+QVjzRalXFIHgcuPM27GoVThR0BjERB
+wKbvOt9pn/ayvK+/P5miNfDKdWH/5/ap1zGssqcrX5td/P6GnOZ8/XjZd0fwCxP
E6Bv//2ezWK3TbXpctGtoqXN/5goSo9XxfT9QaHfnwtzzCGqNFUxPOjVvmq8ndr+
gvz+MllDdVWpPU60d+rXy0231nZWS7gu13d1jDa8H8VoAcM6FIKRUzwVUMo3snkz
EDmsIh29By4owfUVcKVEndkoMNf2Be6/gpW/LleCBwMI24QlrkLQU9qxL/V86ZkZ
J0JIChkl1vzpsDX5gGwJ39WH8JsXJeMZtZWHpbcN22urPsuqGmJp3zh0XrOZTusz
n9iT0cMVLZVlz5uX+BvsTnRJZn1q/Ex46r51qq7DFZDJOTS7vxtiDIoasRqc5cpi
HrrOVaDaZ5Nc15mz9x7aEmJmuhSjZJBUojVnB+irxP3oy4IzvwMQu335D0Do5OLK
mKPwfP/8RnE4Z7X3bmvfwt7TJnZ1mEeazeTBnJSrEva/A/DIqdCJpfhdWF4s5ojl
dr+t/hV0YKgGMkJWxUwiKPAMh2KtJTfKpOhkuMhpjw96DUPERFXZlMlymFtHZTmT
yG0miOnr01s+RYDI1ALBd3zjkxSoN8FM0V25mfsDxMl8LM9adKYt6yNSsWN9tafK
Pvg5TSAPCthQnZDet9ooXTDO4hBHwnCiaeEuwKHbpl9RrbHTsl0S92Ab7jSQZxhh
dddfgzEte/ZMuBLl0rkE1nIQNfFivRxRRqD8e9Br/yiTNsYqXLMvn6i8ymunruMT
DiT6/yI+zEWLuwAxQ6vCjC+6FOW8ZNHUjuiWiTKflJ5FbVJGAg0wFmSAoSisIxhJ
e8iTT0xfE2v6wXcTBlBLv/iUld2mGhqcEdcMCCGlBtn7D/BS9/OHtp3t4KDZLB4w
IV8iokprrHVheg9eMjR4i0KHEbu3MrzZP7wMSv493fK9dFYGDhhXx0LDEcWyX7LK
CS0wJQqChAliZ6CR91PLBmsPu7APg5au3y8qj03WR6mMLQxvUHe1P2MUfwaD3qe9
n+zQ59llpEJn7WIImgaFLksyUAGG6wGYM+AXoFCgzALqPGAA/uqxz9FACTL+5yKx
C7akQoudXYAEia2Hu9YPrPvhe7Yfd94NaOowaJ5CqztUX10nEupNCgKb+NxI2ijp
y0W9l+wzZnyr/ZVutE3VzlkYpaO4Q2thuWy9PHk20UZhdQZkuXaHOKZkDBpyRo0z
Kpeom2clAdnIdWcODE1eZZClyFuFGi5UKzcAvvsid6zyFAEucERY6ZL889NgNXe5
ZzICuSc8aazbWDs5UiJmJ1aNz+R4xY3CUzMzZFPTUkJ7p7juviOjIvDLo3C3y/XB
l3uoyISfKPwsSNXA0AIEz0DzVO6QtYBl2WXv1BKVI6GDE6G2nw9aCEnN7RntTKL/
L8E4PT84YqhNuAW61gCT3KfTSPZIAHsUlwzwgN7gpiOjM9wXCwv8WWj9c/ImAP0i
P3n3un1qKVa/ch62EjYN+SnezBWFxcOxvfZCYXmlfLWdYjXMdEjDmLm3ic7X389G
0N/WeEM4HhaT3aZOZAuTTaqeXIk6LoqjqOsdIxuqIkWIdo2K6sFUcrcb3rdFstKK
aMZvZNQcILVN4UbKnebHbj87iORd8Q8GjVAZM+FbRjTORZh4U/ihiEGHDO4fKbXd
yUisiCCduWFPWgu8nTK2B/bO9F2g4hX7II7LcCvlMPMcuKoiYgZGMwIxfuDMtncw
u8g2NFMrwfXnyDKd5q8kjFR4VhiZdI3rnKax0+MIr8xRG/3WmOe/hA0oQ4+SWTjV
nXRhw+3yLlqvQscmfCEpt5mMx75iCPmGZrWcPmWOxa9mkb4ewbeUxPedyAYiFdTy
If71XTv7mIpICljbQp2orMQghGr6o3v0h2iCWQ4n7g56TdKv0SImgY4WP99mB1aY
qWtgTZcITspv1dKoEsNk9S4HsaALppA/D7BarPUOYNnV4rXD7HohmyNvFWRrNG4Z
40y12v99CL7O6EKSYGEj674fSHyqwOEA7SJpqRcRAa/nuVj01M+3U/ibMvbszaDe
hfGlw0wN8HVwE609P71chteJvKWp56SdjClP3k8D+THoG289d8A2Hq4TSUbKQeCW
qOsFEeDanlqNrOSHXUJGgHmisccbeMd32sxXQNBpcS4KtuupEJahGo04SpH/aw18
Gnsj+5b0pGrrtdv6e7HP9C7Q5WXUGm4/hgY0YHh0Y3qxkokqm2ycrrsiqY79TRhs
4J/+HG2v+nuYHFIK9OsZYN2UpfPxALmlaOuFdUOEc9sXv04hYazxrjbwaBpUfJu6
A4a18NLz4IEsZ+BvAnWA4GOVskia735fqYMlUPVkjN+8eSLJAdd0HfIXzjO0ZCgq
Ca01JMtjJxaa6RHjgMLzkodXrB4viRgejH8JrDTmGE2+mSTufFTfHd+1Fq1PtvB3
ZVXsYbF1Jjbsz6+kqlHh2giOxfezAS1XLvm4QLYpYXzF68aJ4PLD6Gpd9I/SHR+r
sjsnpCSFsFHVj2/VV2i3SiZ9eRpUXCdSAG27u7YBCxB8x9SdMwR9uKxyy4pdOn6c
7kybOYJIyNCJIDyft/58pJz3I+0cI/DrpE9EZxUR0LKpTya8BwjxFw4kx9WP+NHh
wNTIiLUfn+OO9tquShmzA9+EIDAj22v1kkI+RsDuvEgY2WvzmX/o8vk+aSaXCYQw
pc3WNsT3HY4Q+smgt+OlzpjAgQe455aApB2v423XUiOKmtDotNtEUhXiBUQADxiG
S0j5cPVcpk87OX+Ja9uT3fxsrINDrOEfduG7lmCW8vt1vpdpE+Yd0ga8MTwpD4i7
GGqTVvcX/9/l8OrfwGSmRSxV8Dm38ZPwclp7c6kjSQMf2Jw0K8nMYqROM7JcxSad
TtvSsDxqz9E2rZe0+V4OhsXoL+ZUuCVn90DY3BtrGxfCbrmU8yNE7qph2aTmrs7W
S9puiZk9TezswO0gdGvhDNvYWoi/d8hdKu3pC5uzo4VzN5dc5mYYYJ/6tWesKxWO
Xrl8gpjdnvg//s6eLzpjCY6Q2fF1OMELMHnmnxFYdgu0nR1chO7dDOr0xxeTancg
JKYZEsZPi3J4w7R1mE80DPOcLsneKWfvdrisnzSD0vKUpu35z2gJXYqPtFCSRTJa
5fFE3wvZX6Ycn0Xrff1xXPIiM5rtDbqpXhcHyasRu6ksTojKw+6MDGnhVPlHigyG
dNJuFKVSiI/2EF2VHUvAN9dOu9+atbsEZ+9MAh58i2qqXohHyGPWwiTZ1e4gt3tF
L+YRaiBl7l172bHu56sKkiW7g/N0v+1n1FW29BHR20QNBjACJwiqHqvGW303xx0y
hTQy5GH/pqfRoqikAElm5uiqnJuv5IScoHo4DrzEI9KA5AuvQir0YukicLnKKNHb
SNVwBMB5O+vEA0XDhJ9NdzDBU3SHjhl8InxJAp8tEyI4SbN6yEisaQgfRLnezr5j
xtBoqprGOx/5kP0SUQutsCca9VjdBFNgT+xbNCkWNCBxqudAwYZnXgAk8Pa8JMW9
PxTUsquXAP40/t818OFxshBGbuN+LYqU5ao4lN15Q0W2Sy/gEx4MtzqR55wb6vsU
YMxyaUddZJ5/cMVrlr9zpXQ6MfawSS2TcrfOx/ZFvf7+OkOJMSFGzH/w8gCNO9mJ
1/PcQ4KYt5qAWC1psPxoDk8R7T01yGDnY34h5WQKkzVL+a5t6Enog6TVZYcWxoYG
ttpdl6+KT5jLUsjJPhezPnFl04MboIwH57U7sDoLgNyfPNEUHpdV2E9wV1aasjd9
tnBfn22XeFmQZsZn74vDE0YTuseWnZ7IzUDG4+G2Bm7VHO9FdqhfbALlDzMMl+RD
UxqWfFajLDVJdjpxtxvc5Lxjd8aPrDPskVb4Zkh2v+HD85XWqoFnwLXHewJApUQo
8A4JrRb1B3zQwm6CiTMRDQU4x+W0/oc3TBndS4itcEe1X8UVCygJ5Y0EJ1x5b+6p
+2C4A+TO5xIZkv7mCbwQli1qhr++w3yD8KFLz3I7aMs92JoidQLyP0nXvhSkyj8c
mFXO0ib5UfXtikdyv52u/HIyK+lwzJ1HoCZZWXEl4KoJikFwhlZWrpn4hLPXG60/
Wk+Cj21po+ryeDv/128hIU2aqSRWetyrG10SiuhDc2rOLiYDHFTcdNVBjj+2NuLC
hT5lUyhpfJrV80Gd0sOgoVpLY7CyzzjjtUS0UDwnIrv5+xdtcwrJfMAOCMNAW6OC
n5gAijI6kyRwD9MoXl2msddGzyOP60ynjDabIHynKQ3htY4BSMpMqWiNZ6nFfmz9
Gzz53PFMDZQGv469PeDzMKLZ7iOKhxL9zfP/ARsbhrb+cJfv7cQanQRzTUi9K+Es
cCHIKy8hqYQpaKveRNseFwPZ8OKW98ONPBKBwxkq3ck3Ef6OF66kWn5yIa97Mds+
1z1MiZOB87fsl6KwNMJnN8m1hHFN8MX1ZX4dKUJxSJ+0wxMuhH8Ng5EimHdck29i
C0ib1SMj9dqQ1J1kSNQKF5+HNNL99+PhKEsqNON5uPy3ezkbCkaw8udKTRnRDSgL
vs/IGI49TndUAVya5kha/NWHdNRrTxpNii5gUjgv6CaPB+uyMTqZmVapnjPcQpLD
3V0aIvS/hOltOoHuaPolyHxmDECell0uYK12B5WlOB7NWlmZPyUmsSgOQ+/pEpWL
CWxcIjkM3BCVpIVSrKY9SsUt+TR5QVueYFbmQ/euqAt8B0jg9km/kCKJNLf3/FmY
NZAdo2vhA60K/jSphcJzwPgXqoMRw3rhu4zoojqM1qfGbF9rrWKDfmBvZO2G+0lr
Am2L65qKDT00GvGtwP2kbrVlbbRctkYGlihyBaCZ327i2n63n/1tVYsEUCuRZnem
N3EEW63Rjoh64F35qAvbfb9WY3qcKe0btUc7uze6vsgQKoJQ+lv6tB1HPgaqMK+u
Ut7HHpObTQR9Uvm+KCPrfqmyjvGb36xN4F4uijyl3ComKV7WE67b3z1lvJ+woLTc
gZcqY9Wi9pZo67NyY0WHvKUXFa1wsxKNQTLBJfWvpzP2Ug+ZsLSZG/h4O+gvX2Z/
TFsqRj7z6HlbZnz1lGzS2UTBv1i6KC6NLct9JkojdUpOXH6UDHMh8tzNLEnU0DZs
51mF9GPPRVOpcMCAZprmq4kv9uZu1eA83ooCYUtpT1Z2aUFoIDC/Wskm6EJdx611
YEpy/U7gz6XgiXk4qadJsdZ/9QYuHlsMFxymw7uTG8YHkRBtLS99HFQ84QdLsM16
htdEB8b9z0zVXUe1eGbUjlhk2LJ3ynMSab0LGsKc8T+7CSrjtaTzT5Cm6+2AKmGX
/D3ipqeLNz1wSfB9iLuhwX1clCTxoYIj6ikdvJdlLvXfFdeE6/TzKbAYCFJIdIpI
YPlu7GPisQiudTrqv17ETOg01bAsgCa9CQoE2ybgZm7fxIEIyYwtbAfp4I3rQgk+
PeNRdzGgfwdDL2oIp5aQO/cHXbP+0h2H3E/xyFhl8bduynISw+ZcpX+eAwj5k/mX
koYvrfl9uW6LMLjQcrU+P7aXlLiEeOBK0i0kFVS77Mf9lOLgLGBnGOX4z5NtKmtP
rsSYiYXvpCzPlk16qwuvOIhCLc4qov53vWRufbixcFC4ne69ArtE/Yva1u1vOyWA
G3dNGs2utg7hUyKNk2NRn9EXWYktp8m2rTg/B6CnWgkg6D9WXXHNjggTseqaa3YN
bh1kZOEi3IbgcASLQSqvWgAl/juO+/3NNNI39Jch583s8WFDXClipMWUp+NMJEts
cTmkpdGdFA5shq1I8LfzZ5zNw4jolzM1PDXpOqDGLcxd/j4ORBt6tdbavWtk3hEY
4uqSbW7tlYc6Sm1UEFkOL9TQ12kgvkodv22D7GHWy5TYolhmMM6B03GohikZbBew
Hem2ZSVE7XXfNpV4bondg3Y4c+3uz1or6lWjRu6aoHAgJEpWWXWIJFq5UJWCfb+s
GCRuDNLAgp5M4Wv+7cZRhclEU8ctQCnWZAFKnP3S/5eV+HS/whqi0IeukoOLZT3T
qy9jNrqV/sDozF4xazlpybxiMgUH3352VElNGugVBJpqTkX0yHfz8EdACcrLiCRF
JiPeMjQ0M23vGuHNnRXHA2phppdFutI6DPsC731j+FDO8ATXp+5bVB8vgWaL6mEg
/OqRVK4BfHPt82k6lRGyNrqcL6fyBuAZpLJscBT5YA61XSJf3XM9dpiixVuOWUB/
s3Mkv5rj3n9lV/zSpHqhdbJS3E0oxtb9NL/hsBlEi/PkF3VFrgSB5qelOkxQAP5V
1/ehN+AGzBGT8qwRVR7U2xAPPiWkmP79LBgxH/ed3W9SV94PRa4T3U+0/sEWlmtC
JILVIp2U8omrtET8O7LIA5HUrXphhCTf2traWn2kfEMReXPuN4ySZBemFAKOF4yc
PQqt8hY7bfuFkz+QKYeC8CX4ETX8CGAwAqxIbl+yd1ZSCnjLQ/dhU4siYAEWLxVZ
I46wNXJ2BpqvjBnDFbNqDSxlRaRtMfGURffp/5BflZrudRcI2cfwEIC+ia0zKx3w
rsO/wFpbBj1YqRcCYF8xw4rt4H/1wJVVDuIrN8G1uhp9bvM9a9F+7a1I+cEfL0YR
E5H0YqtxKrKblC1QCu9kT9MfCUHx9kUBm9PGlqUG6wwtjmxkOetp7kl08G1y5Xae
1Nu5XfBqyTDVJix0yNkMREWkahX3X4gxb0KhrqISxGEFDB8LHL9JUeVYfd/Yz5X+
eofJs/XXTUKzjuzu5jt0UXMdXrQrKmMLI2ibfnZN+Us7xZD0acNlJxR3K8u0fA+B
XHwTvCNZ/wROBzk69Ltn+jFo8g5UCMNBXPYyf9aXvgGDuNsdGvvPcUg6PdrYZIVE
NEc9C/UVSa+wNSbVmsAwDw47XzdhYSYOyUI7e7jro2Zp+YTPrD8uqD+xv8/IkFck
7+OSt88JFdNaMIc2AEL3tnxxyCEBA3WyBKScgbf2kzl/7meuXbjd7JGld4QUW08Y
InH+WWUFlhz257gd0Xh/U7317kpC6nfE5LdE9FQldt9AuY+nvpnwBgmB+mrZhqeV
+njNjUgpA63E3vnf6NWCHpiN3L4E+Q6yrWO9MqCpTlWjwN0iohcbaEhl9WsqTxz/
fOd2KHqwqJAy4vXlluMGcpDwPU0vzsJpJDe9rqicqxXStcpFzlYTgBlFkuvBtIFA
l9217fH0SobdDEID7JkvePDkoE4IlhxtRTY2/+zX7Rlucm7B3iXan1+8ou+5bnP0
rcTM9HZb5HvksSxhB0K+9kKoqT6QPQ+4kIT473+IKMyEi6fAPMEMR3g094pvnZWu
GkopgQFwXlPbRTFaJzXVf3juM6mqCzPa7YdEuj7rt0XN5iH5YewTzKCxAZzja/se
sBH9e2xqL8SiekdOkeHpKSiIlfA/epqPrD+Lecxs2eF7xu9TcNEYykTBIFrXhXyt
iivpbg6vIOckgOxyleAOpxBda16POZxzjhp0q9o1ToKkWbcwgsT0GBTyosp6tTWF
rqT9ao76Yw/87vvV7voJkI01IVQKbF+ev5B5NeYdGStICqkPlgHNej0Ge3a1MEAd
jIApMy2ZespCKocpJ5X7uw5LlHcv6q6J0dEX2Zn4rzhsKlUK4gNW52SACbSVKMFg
3rZuTPngUyWKC9qXz+lLsX3kL+2C23CWCkHjW8IJRDJRyHZ1Oe3rz/+f+5xsYLGY
f4HMWwdsmUHWGwIX9wQxJ4APPmxCQoH50A71Hr01m9qKSivuX2HzbxQtFiXrRNQ1
vfGr7aN/w3kTbC1UcbWCHr63GGD37DgvHOoCQ98E+sV6mt/7rVaa1Fc9bbbisSSc
Qdd4e3RKCHaEKijR96nPq2Qc3OV5J7aE7Z9EB6beZ5NdqXpn+MHI4dwfmFaG64Nz
VyWccNWYH+NP1H7w4PU3N5Nx5sSJTNdiyWvho/Iw5451D1fBYLEeXRC35H5fGy5+
0Hb7Nub9Lz1dt2veOnm3X97Bdb7VeaI7PMeLxcS1TFodeTKOgpLth8ePsNG26b/Z
gNOpbpr60/dihadCWMejTXF/BXPghzcCJF9AVGz/U8/f+xTxapYyxuHUzpXZ6lBy
5Pd/5cLWFX4DYWjkPWMMGnT95Ny/fq/bOTLbkg55QzGyrLVPTwOvpxoWZ06D1EEp
q8gPKY2mGC5I89m/fCXeEb/uQGv4ccADrE2ACqj9ZE08Zfcucd+XOxvCfL9mZmrM
sAAzbsKzcq8Vjrr6/oxMvWE7263YQWLKHnOUNsoaPBpeyO6YwwxRLiOIPV4rUMzA
vvFKY3MoNEOE8XRrAdkqf3pZ6mqteemgq6ynH8pcY8C75irnKTp1Aw5KLvLix/MD
SMxTPqZGGw3So8zNYA1uhO9zW3ffmqHO03v9p5s6W8B7tYugZzQAXNjjRTUxRdPi
6nQvAd94R9yzX/dxfA+wFbf3vCJ18Gk/j6v0g3kuPy6Ui8FdrNlTXU4x7mBJE82K
hiIakG8MsxVvF77yaWaQMTd9OGMiBklqESP/9sKs5+VEPJl2NL5iW9we4qtNCi4q
gO4QGJhLkNkfFMMuhYRU92D9u8It8FIc8no2K+oiddAMX1/k6GR7haiUWtEthTpN
/jw8eqjSZPE1F87N3/mCx9dYTkI1EqI9hdDyfNlzFItvupZzWC2TO8d5CO4KWslG
DOSyJ6Ikav6uopuBBwhShjmV1YfMbSiGv+6+bGXCYHwWWgOPAeVF+N5axMcHx7EK
ENEtHd+Q3DSM01xeKLuVWZ+1g9lPAzNewQgPAQN37K27H4mTpuW/qxIVmPBKRO6i
D8zYA87qtBVKE6GG2czplem6jgRDIJjfdb6vr4GdyUHqgYvFgWFjqrNEYIKTGWBH
9X5+gDeGnSmLNLTVRnbMdVvBxVt3oPjUY/AFNZqlPB9PhoaJyb1gL9oTXdPQex5I
BmAbBYe4mXpYl3vwiLnuX3BdbiqfTq+9mG8UpMZdTQZb0IjSnzx1NtYgb8Ouyu3i
MhLGBsh404hQO4NIqycZz9q/V9/Y3b2+0l9jrEjqCdLqYWviVUxnXPL2zs/yEqwQ
qqZRwbjDyglJZKBGgFH8fCoedkClo0nCOCzs7IC/94sguIptiT1gtxanIT5RwOnj
NVW0s5oW0vwQEinzOnYCYnSD42sW0te2qqsWLSuuTt9BGNl3XJGNwQ32hnGMGMTa
x7Vf4fUPqvTU4ir4nZp0LHNyaB7P6ofczaoisXgpCBqnpaC2nCU0FyzdENFKbjwu
bqayRMhAgTyk4ulGZQ4YkzB7gOFV8DftTw3XBRYtcZ2BLSiYrV63RjIXx2Js9GOu
FDLP9yv0ZPyDaaFd8By1PvPoSv4uSJj6vfcJGx6vA+InTTDoVrCRMuGcY4aqSRZl
7xlwPevnFyImhq8cE7JRwfuWmfJrbTJRALcUc0+Zuv47l9+JaO9f2BZT0mOMOgDg
ctla+sukazzDntfFZ0AwaHNmHLZkQzX9zHrfJHSfFtAFYdEo5/jD08nA+G8gK/VE
rs5SZj1wnqepX+SzPjPp6lWoI2ATCOkGxPFpsz6Y9CRwj8LmggI2iE/3P3Ya/CRC
HqTNSHNkNI4utNA0JHrFkNUGtEYf1MU65AlO/mnKuAlqJR66p3WamVP+jNnSdDRi
ANbU7E/xH8RLdTV8Y9Amut75X0HpvvafMagmjdBJTfPi0zcB7elx7+3yDCmTU3z9
uGiKl9rw1uDu8ZFJvCZEMkZ0+3YXOe5CcPFe+Jcu1rDBs8aq/qip3J68Ubc+QDdy
YKJhWU4eS2HWkwKYaKsVuqswuvtxb59I/1ko1SyjSFzk4HJTTSkbvU3IPoApgsqu
3/H11emPQSq8yfgbYdrgMRHbKGOBAz375wG4Ei4FsGvxQCRUfmEPyX6MpTKLTvts
LmWPVRxlDCLnpOkJmnfelfjStbhnCO2zdMAKmsbyytyfzR2OrbrZbgDuaakEx1Mp
Irx6LVWwAESdwACZ6nHtNCdKtZ41Hk6gmcL7Q1CWqt8ONFWMv1cp8ZzZJih87RV0
ZTEDBbLKv+bnA/5nwOt6NEeX7+cUMS3BQpRKavxmRZzXmGj7b8iB1h/T7s6A+CE7
fBLuWnBvQOn+mguGUlL5ZFXjZIAwIUKBTPeXIhEFD9MUFqLV+5zt2zFD7gC3Yy3u
reF7Twaa6FKtbHjFAY0UVNDV1VrRZJs/6+UBzhj9Ys+FElsQt3Yhv3WdgAmtmb8L
Tcv/YDW6G/CKqhsvU8aYKYs4VJiSW7dM1FAQpCrK0lByMfVATQZU5qPwzognL5HX
rK79tkzNn0p93lhi5pt/jfWOtx4uhn0nw0yuhW0ivlU0f1D8HywRTpQK5jINwGEr
CbVpzcA70WDBBAM6SKlK7bkbQD28HW/8aMrLPDCnQ46EBiZ08tMXft11Yp3DB2yV
rJv7rdiZZN8nxB+R2n0xlEFDCzI0SF/UX51a8sIw4oyoAYTJSqGbr3hkx1EZqFCn
E5+/QeuslevNFiVdq/YFuL5G/FU9MeygSouyp+sTA0rAtf8LlIidYbsegc5iZYtY
8A470dQjuBZCMutlyaZZWAYG8wvCWm2vsGzU9Ay5nPo50+aEbT9ZlGKFoB9i6G0H
JwiLk2cHWAhHRAOuvQ+Sn2RNaUE1EGVOZIyLJMKfhcbbHjRybTZacFnlw8YMMM8X
qRgZlugrVRDgU4WoyS5qxLfQmmbf/K9pcCgKhhr+DIOwcvIarmjD1DSvNRN34Kie
DQ0h3bcKmRVnOqIA+oAV898qPRLwGk8FAShf1DIPLYdxxDp5FtMNcSy/q7FQdosp
JCRF0VEJMaZRS/BlkSWAnMlkV+aPQk8kC7ekawOuu4Lip2dAUaEpnMFJBNSyOcVK
V3aDtxen3uVefhKvTvcMWOoYBOmD2In+qTkQUqUYozuMaDy3UfFybcsIct5lc46y
MM/Dho0ajuvAZb98bsHIMLpRnFiO1TtevvQh9QOfZgyHIxLFzzmWNjfS+rLSyJR3
CgpaLzBg5o803qadUSyTfNQVQR+fPr3j92gnM8D2tdnxnozjfsBeq1l5i0Ctosb/
35VkdRcQZVlXBa1W2sytsCqKaj+H6eF8nhdJKpsoqpUD3Rv337OL1zjTB5c9lNRy
VMHIUV8WzjZASST6YOJoFxG72YfwVuJPJMtObHmDseK7PeRgIbL2c3XTAG1vJSdD
LTDuAFnjkrkd8I7ISPbnBgbIPH/HqBRJZqZvt/NevquvrlVZsUoCshnkLnPzr6K9
TynCuFmGYJNsAshmHgZVMAAXchZIfeMceHBAxlgJM5LNIK5iuibCzmt/fqT1OUTH
/9Wf4rF/Uiio3OpwMLXL+9pjNrw18LNjbVeLPSp8hpeD6KlqbYRAuS77xFoMJ6LI
9/AUFKDMtVgzFaiSUpkXw2KBaswjsVXIFhgl49HeNuYjXLwP8hUmN8OUTx+7y4lc
8rL75Xc9Eem8yeVG9Q5lWDnZqfs/j6tOEYqE+5pEGQhqiufMGqYAP1cMhqTiVxai
xmsIx8O97T6rrtGAEgw5lNAbX9bDhsQWXVWbF31iNRYuOXuwOAIPhegm/VU3b/G5
gWUaH/tcprSFHihpeuV5MDb9T0drUpq/1u3UDwM10Ye2KILnyiNEhgtwrIHnIGew
k8gm00DXCqQTAFs78ymU+sKj9fEJfIJ79Ii1F2zFpVBN7zYVARgal82McYpiEls6
F/E979glutBOar6PREAaRIku2UcxtfORuf99XfU3yuuNgGjeeY3Wew27DTB413qT
NYtOuZgHhPqDMXoz5IehwydofcW0DIqeDbuwv1zT4SZKN9OXcPDSnWZmzijLh/sb
6UuILBnqaY+rD9KVbm8wl6Ug4lI4Il9aS3qVNqmT02eMlrap88PY5Ti/5goHbaiw
Y1ihgbagPT/nR5oU4auMiTjsBqCYVapP/4/hqI8LwUQRVqanfp1TT1v1r5lVHzm3
9JzmkMIbpfp8xnLyEsqnEj9oVGjWCuN5dq98AZAA87AL5/KzFObkiXtvUHk6Ql7h
LnINnqLHIWpwvo7U3pxMdZajHEv73QPwmHQHwTaESsFsDOWHufX0+TeeBxuq80/5
iekBVxADaIH30IqokoGJiASQybvy4bbvY4RX8CotKMg8Y6OXuJgeqMxlpzagKa2W
zYnNPWUcwWgsToLYT9OmwACwf8lsSdJ7WUK1EVsOnmvrYUABryzIH1yjW4O9xwmw
8NVvV0cxhOvXXY7TDB6Ko7/SkrHt+m5LjGIJS1gTBQgmVZ85Ntm+SqTL2W2+j24z
fjkrWQkxWXYDiaqcBae75oSWykk3xcUr2ISgDeTHIg4uWAHCQBV5cuUFHDFXCKX2
fPepI63KeeblpZi+nhmX5QcOxodKKwWMmQzPrcxtwVXxS2DQ38hBAOWfOdvfgCmN
8p0a+chnRbytmfLGhlPSiZ3b9QBINI81IolDq1lONTDHSmCa49sKojIzCtP3d1av
lULjPdyi+17Z/43nGDArewlTzObBIpLu7j7LG79y6vnmBDaKzRXyWzZX6jof6LrP
pQO4c7UR69S2Ky50ar5d91ce2Pod6awaxHPSa1uLsgka56halYLpSwEG5s9FGZYk
W2QFI2dD4ztIAlhbsN9NQ1L8+z19j/+clDN4sMEdzAL1JtMDmVT8O6WmMObO5wzH
hiLUvujIYa9rF57TgubuBzkA4jjnHYAdoSg6jWpAPqAvUSgFXllHWEHpo7APQudf
XzdfFySmVQbFSbQFeMytZpJRjte/hZKIY0eiedJWZbWBoPKrJiyCMWOwGCzfT0Ny
Uw8Bd1nS5kKD/FF3/2iDY/oYT0Z1FpiYy0jb9op3YehOUZbKIOToMqD8A3A1tJat
y1NTz7kCLUxDQy5WkLtChEkNF2qZg3K405KNftjSWKKw6u3wsLR/4dhfSjd2frDA
dCG0Mk4k2F66NsweK98FyrXCwrFTlHBsrnUFkMptdX4B7vVEYCNtkfWZD+VQAJ++
o9fOH0YrR5RcAs0DzEmnJNOEaK7IZdn6dt1g61YCOwP5VvSvqImMBMk5WIOqfxgh
Lc9lrzKC3eK3KYcRWTMbIrpaOUV8ApieY9VscXsBaL9rj68Ywwc5uN5qizDs8dZW
r8kvGaRXoMQCHT9GPR/qistemvxLyEi41f4fR9AwqAjodt+5dg6RGvV/RF5jCZDb
ludPXsiFBKqgkPPQKVodosVsvAK9wlY1crVuuHxiPpte8ka22Qi8CKFf5lYXZN9+
BXpz3+e7RARZmK1tqbEkPtbFUUW4R7uW0ScYjnAcd2jll6kRyHBjzBrSWRiPwbS0
9RudJTDGHsqHE3wK4+VSuPMUMK+KbPk0yJbk9A9M/7jZ1eph+t3/xpNoOjFDh7C6
bnBUPfgVH0JGDUfwdVcZsyAceqpNru9Y72PHjJx+Tebr5V++SK8a1KTUSS00kAhd
2FbgMmHLCpLIndnR+/rRAjouZex0H2jBiU2Kwc+7no0rvt4sAV8lYewrTNBV92Ry
PzyUEd99sxMX09vurZ8tLW3xaYetW7d4mCRYw83zV/KexRwAOMqAC8rk+gHo1Kfi
Nd5vmZMgul/2aAy3e/hPi3ol+qPsba0lyCJdgqkjoXbe/cHtrk2U08WH5FU18U46
dccslJSHwML0aATmRdgoUtDw7UNa0AykOfl3EQGycaiRdU+SrmEBwPyUmcrNURzd
OEKVx8dDXscmbcl4BAEkTzTmK8LbIr+9Pbx4xTmrH7pXOupTQwuP+C817YT9tofa
MmALyEtD1GEVzV1of4LBIZUQ3qZvft+kP1tl835zjkY93F7xaJyJ6scMfep47Exv
V3WeGwI+2fBG+oeeX7d3LMJWLdjua2r+hXXCNF4/pMFHYBZpTTWSedrRBvpTLisv
n28qsKKMhy7MRPxBOq/4mdCwJoqf6ozezgqXm7yJSif2P9h38Q+l7o+hoBBkfuTM
C2X2PjERWgAI3iGjTn3DD1wn5MjWfCc5MEtXdCMB5dSUfUm4cbL3IYJ7Q7pRTbOk
anEMyvJ8amooqmE3bz/i3303+wdMLnf7YLdbG0HDJ0rJmJYmQsPuKe5BcPvFeq3G
bz4VkBCKRgepCi+1BrzQGia0h+8/RVetmyGefJCgZdn2je30jxQJJ7+sbV1b/xz7
UGlNGwvOdpfv/zwWO38+M4bBCEgqQV/OZCDSRCdbB/TWbKzwxWXO3b6KCj8cgV+E
QIPmWNxop0/VwVDAMjYT0+A8XfoNG/XEKzJN+YabEAF03HHDazm+NVNKg4300i1s
Y2Hs4KDDiui6mnJgFgPyrG2JYx9bBwWarOYo8SXEKHq9k5chwuH90uOk/IIWx4G1
cBz7STaZYEpU0jJsde3EU3MFd2CQq0SP2HPHsZ+Kl1c6L0ediY5kc2OQ3pEwWmgi
YzemacPNqf1j1tshFVVpqxW3+DcrYGufE7qyiQ+uSc0awMKi3sDv3eISy2hglRge
u9QUZPcGkno+0a2WVsKwJa/WAMA8NQ2MebiMoZ7q+RRukVL0KzUWbtDYCkrqvgtC
WbzD1Cjv7Mg217CQ76v1NEjex7e/YX6whR1UrOJ71V97FEpA30MuoYtOF6LHxUCW
MJaf8mDsh7Xgmjo1Dyz7YGKzX4vJucu5gyrjVLFTNC9W9Hoq9qHfS0d4nIVwNA9U
jHGoOSGPXURUMf662CxtSeg1dKiJTko3IqMBSqIUqRDe1LoAgRs6eqKJ7ganSG/B
RfQRt3YyiOFnvmga1wq59L/2WNcI7ySwPKGZQfUMTi5A2kNEpwhpXBpWUHwsctK5
Vhxj65Nmo+P6h0Yp6VQrX68+zZkLn0p6fLbBxYrh7ub0XLwLqHnW/C4nJ3UfWhwV
UKgkHpYfQ0vrJZSARC2H+elCA7zqrZ8Que79CU5mzH9Ak/n5hlYnNxG0y1GpTI27
+2SPTmT5IK7QjB+yfhVwocVD+38dUQL5CtCTClhBJmFUbuIb2qLGdEjZBdKnDFfJ
/NAii3WPvfVqr4WWLoa1GVO8JoS/+KZmHWwFCtdo91BCpwjlYyN9jbT7fRC53Q9k
M3OuJTHxtnMXFioN0lAMvnn6nKpvZFabXMZPoq4F5HWLwuwYFoQWTSotuTUAodXt
VAQ/2LAukZl5qEwgov+FKDlV7Z2c+L3Bdq/lbV5S2hmdyC1uza5B5tOlR72Ew80A
1wL1YBCXgDRaLJv8a9y6/a0G2T9X1EtmMCpDDNeYWDhIjAkBcNJwYAGXp0Ohw5lj
j+LtIzMIPAvYAb+2fxc76/s/2OfZwn2WYBAX0SC+tG+YvJ9TEJCnHxDGGFfZfnB2
KS1qi2RNWIXXxPlxdJqHKACkd/Mi/0v7I4fVXWcYFk/C/HW8aVH3Fi52R7RIM064
fQE7laIjYNVtPEH9Rcqmqueim0kzsNna6C305X2wFwD3Vvy2NLeUhoGUdItOA8zp
9n6u3gjGPRKbu2/MU+6pISZ/VopRWcKsm4gEmD8wqaF/XZxxd6roViCiyFmb2mbw
YY/W4ytksTyCnsCS/UY1W6Ax3HAbpei+TAy8Bh9lAs7aQgXzoCrUUYWWEjK8e5Hb
BUqI7aER4GJOePVUQQHvnwL/8BAPGeTLFxTQ3yUr1XniI/3P13041kYC7ERUHUmt
WsAFq5vQWpAbjAuoV4LS5X0CEkPrloY/mRlyFpgBSi6jznqdcN5ueWHMI0zHETSs
AMHcud2xM10kQpkht9MJuMNIIP0jE1vsnpV+2s1pblCV3qbT4Lfk7wPbge7wr/Pp
fJa/13nHidj0TK73MgEpfDxKqGOOMZDUwyvjQIkA5ybNQrTumnHGRh42KoMRefwb
t8jVlnqfpHY6JCdAK+AyVpL8xXHi2oFxMh+/CjKGsJL1vkc3DVegcIrcoX5e27Q5
0ljDl8HHMONsq637EmigHF2VVhpANXSeFgRvAKadMxPnqI57HPDB7sxwCKef5w9b
AvYU4PhTcSKN2g7nvGiRv6TD8lTruIaJOb5kkgJpWV6DmmXNo8p72SZl7qyMRUkp
jPHJulEa2/IMboZlvkAMm5VAOcmWmjitr+EeIoZJa7p4DjN9VDrPOm0/Z+NHhZh2
AL3Lt2lvroOF2ddpIW9hVKC9ui5Etyi2Rg805jHk713XfxJtHnfYP9QhIGcn2k4H
9PydsxC/yf0ywENad1BC0tu+0+lVU71+wU6DGBF3PhnfpEe+iWguYE2hmmvS9yUa
hhvOlTZq7p1z/dCNRxl/YuOBALAM1I/GFGJVyaBaX3GbaWfIy9lUOYGGt1vhAOWu
5okL4owSdPjJjzHYl7CjjBXeDFprtmfawjk+biTX/Vz9QcM4U4JPzBGhw0or+L3/
fU2it3FsPa7jzC0OoEhLM7cL6wY/LF4UrHIDVP69naebUsZruMbi/snCwqhygiEX
fLmQq/H3I8lLbykzNRlIBv5hMd0oF23hEH2jqu4lm27Lr76eYMeQRaXYZTDgFFz+
E2D47h6dpYK6LeDI5ExEyIrergUQXNlF37+AmrYSQlAomhQgWhki6GBvM88yuryy
zxxIi0jj9WopAV7oVogUI5lcG7SJHLfkgxJ13e0F4qEJEkHK3A+79/WJ4WFFieXf
SMskG8gzSCpL9TcCVaFR/f1vcqtDgVM24xUNJTpgBf5WZpDPWO+rRdhsX/r5u4zd
YC9Qrt07v3FvcV79kWGLEmBdeWt2ZjyctpvNABvMQaRIHss4hcR+mW/Z6NaVKqlg
iecebvjk54hny0X8ZrujAyhTA2Mb6APyqA18npbXUX7HlRoCzrQhNUhQstVA87EQ
PWo9FiqiT64bfSNGV9Yfy7pw/EfdnvrRUnMeVNMes19Qrt/5FH+mRaJ1R2fiFi3T
XUEk73htnJrq0DE0Gh+z4dpFQys062rfd6p39cz0T2w+yVBV0ObPfuuINSKxiaHl
6uarZKgEkUPyArOtPG0iv1mvderoiVxtOPtrnyUUev1hx8dIuQzvX3rx5e/Ih2s1
2O+w4lYC3UL8xJyxW8NAFlkTpcEksoY03+jObwHP012NRl7GS+luEdywik+ax8ZF
uybFz60fnzfGJs18euo3qji/HonsEyCHtoq6v+IaLAN+OQhF1476ix1A8x41mUO+
v5J+XzRwdL+VR5aZWJYQ4NBo6faClOg/OkGQdiPh6YrXz2jcqHzjsyf2XrBKiYB9
sbfATRcOJ+uYcN1BmnkFkqJ4fATw65a94916mCC0C+Up1TSwk139xFV2swKcdyzy
jmRqEwRDgviE963Zdw6D71h25X4PrjEXo1kyEUrhv/XD346phcPSCstTKEXxDlz+
ahHOQx1yR3KgSBoAZJ6MT7Bf1Z0EkQxKBT/FzBpzcf9t5H9zuUaeNGJNHroUj/96
50AgY1RUg5Hl1FtEvCczdxAHLzYP9/IwfeIA86f25eUc257g8akv9M4+EhlOxmKw
5h6fVHLsGXL1KE4rpwSWsN0clCN1GeLUEEGz8lE0hOp6wVa/hH2uHNzxCjn/gPcv
UBJ9gcbX3P0urIjI0kM32dWeKf7RQMgommtVrEvQQf1cTt9BgHcUWnA2J7EU5oUY
OwU1a3PxvQPm8WX4EjR1SEHUY+3p1oxu2tXuHMvY/NDu+Vsuq4O5IQtTCGg6KH4M
J2s4HKfErrXQqexw7i8tadOnD5zhS+L8hsl2Sr84l5JoBFmiWEB5D7ZynbJKHT/F
Ofhrn2hokhWC9fRVejv1aQgtgrHoVIs2ecDOGf/lRVdP6FUGtr7l3Fmtp0NNJYc0
RLWISuMez9Rf5R3KmEOUGGOeGgZCc/AFbHX5ZmMQQw4OjTHEV24pK+qrzIhCpwo/
Aiu4j5FmwtMPEfRtLZKw+PF7H1x0LWLVwpJ0PP8O/F6HXMY9A02cM5USoWCcfe+r
vDjRFpDcZnvIypxbLOcZrpWccIcYNN57Ukzoy/RBFOHws9gKGM01V5jRrZta5eWD
r7a3zhjrzqdXOecOr6dmpvAT0ulQJfdymSBlrbmU7twn/fsKKJ85sda7ctOdX0Yo
s+dNVi6Hl+Bb3mQUk8yew+cfYI5BFM2GgP/4EwAK5YlAy7wbWszlCol7R5wivYiD
vbsgjvV4YXG7LX99Xp4WAckvrBks15BbQnQExJhSxMPR6q3mxBeFgJL+r81N1bd+
eohfewIlabKChlEr0a3XVqT3YCItUMmjCH+mjg7OIwrITcn8KZdfTURHea/yDEpj
VIF3icu3ckqVWeVuyrFRqXLCLta/QtoPwDtFU5TZCUuzq+kFk403mimIurVfPJC9
0W15GTti3JRNdSVEeClniLOaekyNl+hlEFwXPSuOE+rQD3fw71f41Jp2mizpn2ne
e/uZp9HwPY2nWB5C6r227Sz0zjCweyzsmn9F4F5FXmAE9n4BfeEUKJltqD9Mn56o
Me0W5j3ws7ZKzJ8UExRXsZ535qh180KAp2xfh+zuFOqQ9MbtPxVYl2Sh3Psc16k7
Imsmzah7eBt+wI9/X7YNSrNgYD467+sFL8rQEzu5apdvZe1F6OoLT1vT5AF1Y7sy
juE9hTBndQZLPAhmYi4Q08W9GJn3Sl7iI0hUij+Zh9ijTWtNp0mf1Iv5drmQoqPT
fj47F0DtjkNOoPX8TURY8syUFCRkXDEpOarz7TNe7aKtFpUB9Sm5L5fZkxkJ88+b
lK011xtx8IC2zaqJZL3hujKkPnz+pGQBKoSfYolwktE6mhltNzZUM6TLG6HU61w+
3yGCVni2HbN+jmK3VE4a7LqPtfLGcFpSmSK21Gqxb+a6axAWKH8ZcOqn4XYkPxvs
tagFMngGwrbySRdPYPqgS3e4jEflRhjXp+3uasLmo/ztY3S+bFjPoQDoBqVXUm3Z
Hc/cz9x7WOamcDQGU2lFE76zc8Vd3YVaT/Ut9Sr5C5uDzTzG7+mxXC3A1mXmYSZg
4xNFVKKu/4m03Rxr0j50aOAcyhPI2v5FfQ42k2ve1PlZ70BNzQk68Pgg2Rv00pYU
9ZeQ69fbU/5kgJi7pnRuKtYKS1ZK/5cIDcFbwkE40MQaGZEimi4Ed7vmbTqQv2uH
sLfbDrzvE+P3TDcpMsWy0Zu8XoZ3tIw88gZPKsH1P81uf8mgO4X8c30E1d9V5ezK
QBPi3F2ZSSOIFDYFYsiQ2In+bndmaN2BISalBrDfGunLO39zjMOq6xFGEBnnfqVH
UG7/9gByaaVeZ4AUIrtp0EkIdhq1mGVU0W3Cl7OGGOHS8UixWmxutnE1Z3afkAvm
tlOU/kn8hYd2YJEfpAq4/KxRE7TWFmZKHTtzMHaLTOs80yXeZhv+I1UedEpnWjbq
B3ZmxcbHTLo1YCirHziR0OPK8Nrq9Xd/lHrd0NhH4uh0pOKGBAczZtLC7rJO22rd
Styi7posSRbMjdm/YSL5c0FD4U8zgqzKo/wjRhUKEuLkhGSruiF9Dd3DUxcs+ubT
A6TczuSW+j+J75d1rESxdbDDLxaUmhunMGU3eGwl/WMi6k4LJbIBfVS0cFwEPxKi
zj8nxulUqdo2omvox0nW3amard3aH0xeId8Orj+wPY3wV5Q/mZaR4A/1IX9G5BpJ
IJkzwBSYZhuozQo13/DPueweeNid/DL+ubKRASro8X8lt+Wi7mhMBbN8cwXcoBWL
5DnsUkthx3Mjjg2cFjYlR986yLJNmaMBpfebGIQpo+V0zF3kLRXj3L6Ngoq5cadO
johzUAbEvFeyXpfbuKEOeX+uhVYmKgoNg2wU1/8eufKgH4gDVUlD/kAIRRl2SMk/
zXSMccMKy9BTxLH3Ichdu/hvaxHRrt/J/9q3FA4ES3bzLHRAMysavrEyZ9T59xLo
GywekcC9s6hYb7tJt3HKoAfWPPUhBb8is7DFVuttVFPxz/25F+ftN+fao6GXk5D2
aqqWxGJobmnb+N7W57iUoctBHYPZqzwn4/lGZdHXWvmu1KTvhiC+dWKN5XjmtSHB
rJoRJJzUgkyU+spMom6eLWfFwhtqX3Q8r9vF8wN06KgA1pN+ShkO/aWWmFY195or
oev4zhjvObuEzd/UlCcKZZNvCmYSt/MRvzWOA8aNL6f/3hAYZULOk7BDfXGD3ZDZ
Gqt1ZPN93ABJLqtUNUynzZEh4LyC2OwZk0eyuZcC9wIrE3ry/ljTppisGxKwxF3Y
yBX4oeXWjAEoDFhIlw6yp8pZhL0bpT60V1x+oMsUzwYk/U/3MG6uYJVytgIWFbby
S7gBTliQajZmH0wvJN+V9phfbZgKbcuZ9BThMN17yoWgSzyurwZVCAVSct3vSjTa
lh3EIcLErAo4f5cRRBJ+gUloQY2ciIZGDATFjCruWr1XHEA9i79vh99vjcJ0g9Na
j+5355ezSkyY36NvDpPuvXfeJQQDPVQFyXSSll513E4KxQ1YTAhQIFzioZpZDIdb
Pp2Q7JQAtio3v2dPO0+3YnjakbDEBdt3pbNBvRCd4C8IsNCY+m7K8u07xG3RW8HV
41al3M8/o7zyTyjC56Be39Q2uefMYmxHw6PwWru0ioipTb6KmBlWDd+OfgwpLJHb
dgwm7xFAa9PGFnAfPw/bCElwMIzZt9jtzNwQcuE7otKpa9mTq90wT68vnH4usg82
bDdCYoMsVqrnCxlahAhNeMAdte8fYTZVJ8KY7hSE7wxrHhmhrValShEwYlkCmCKl
KRS5dDLO6VhWw8TjbFTewMhxxP9EqrS1J39N8yrtxkFIWHt5jG61UyY2qNBPtzDq
3HX/9VK0/7w2nn3IQOHr/j8Onephhsni/n8M0mmvWoF+B3Q2AEUrCZQp6WUOSU0X
kV7aCUCJd7RSTJ869apGTLIBzIfzzroaZw7sPw4k7Lq+LRGT1A1SEmlDc4UQAnPr
/JtJqMa1VHu4i1mNrQADwj87Nxs8BWX8/ahjgJiQ+vrV66vL0Wlrd831EFwqb3cN
xXZJROenLa4avGNpM31OuWg11qNUr3fma0582N5+COTD1cnPbhpm97xh5pXmJoI+
Zmd/zeKoBWCI3PCMZHgINc3bil2rxKY3K5O6iqg3q8TxdIJLKBKvZMohz3Aq98Uj
IX/jGUAMML8rT8cn3gpYBA0nYqvcUKkuSjoEwH9eV7sPKklCGdl0/5yZ9T/P3xiU
PWP8P3RXxXuwGRWjNSL+0NFsZ1RDn3Hg99JlP0o8F95RZp8DC8b94cOIrjXgh0En
LyylxB1APpwa/VemMlKt10+REOo/MqGVtdepOrMSWX/RzFDPh6CeS4bukkGJvt38
om43kKSHVH8CwV8x/RSkRgAZPWAI0lJxVbZlu0hQaNFs/7FDClpON/3nnkl2pHT3
hPNd5okapEH3WQdAwW8AAFlxbGoY9nnHn2F9NfABWMVwB4ZZ/qJVMIo79J+HMH96
RLXpPoHSKPGOK+Jzm2eT9/WJ77wJ+2H1njtLj9vV3zN0Pp4RLB82LIJFaE9NAhRl
quT1eLVauBMLIIjEmPr/odeDBAkauISzLZVYsG/I+hdx5s8W+9/IaRIZoXB+Ip/E
5IBAScuLe3HzAyGUKqZ2EBcrgbE8RTZ1HmAgYaMqq/QVU/RlFC0vZumYHCtY3I5M
CHD8NWqHTV3y6zkOnt7a2nf7LO66UFBozUodqbwKGF5ab1oGnZo7UB2DtrHHbbAG
IXNR5O4D68twXaZZITnd4Mg9WaVf8Rtrqn5/BWen55tSnbneqWSzXgwVehGKZi7s
2WS9rtH/zY84hJRKpkvVBIdeaWQ3rSoyL+yQByncelapOOu4iNFNNF2X1+/o+Id1
mM+YXafLkNPzwUeFPhq3aQjx8pmB/Ifw9TQqLBYCY+3Oox2esV6QtRhRHIa5sfPk
j48yTzL9XW0+qPr0Ysad+ovLi2pTv0qg8IkhIcgs+ekw5BC6vFXI7W79ckoz7np6
HLztXbTBjlxUuY57xkM3MoixZFO03Uh5SzADI37VPXg3A2vxFffVLUt3myAbgXJx
AU225wbN8MWITgo2XiJIqgtU47Zs6sbIy5MwWCDmiMXU+Gi5T+hNJvVG/dbxE/nt
t7IHfUwUJk3ovGeVfXJKY1jyjI66LniyJYZfrM+YVwAgin3xRcqPgUrfnd6sNOtM
ZSwX6vCaHfvCzejcjb2QzuIe9RbtVBK/EGnWNcEWnbVm/Ey7ueasrk9QwTso7HRq
tPuqA0fsw0LNS81xaZSg6JXEzgoe5ynw3Pkc5M2PXhs8BR0TCMy93+r27Kufbrgz
KKsybMtIVKj5i/pE/j83ot/SXdpkWkgfvhNGxdnoW/LOqzjcwFJvrYKGEgfLBB6j
xWexx1txoTN2oi0xp6ZOBsIzKzRzojw8E2mGEhM/a9y/DwG87OjROKpMmw203hGm
pYw7hKJTqnBDScm84qMGqyfEIHwzsa0iy7hHfD1SKKIvTaiRXpfUBxslgTFRhAoM
5QG/dDBHNoEpRkHfpZAC+BpRdaTJqtLRPmSHDsK2z8EJ8p6Z912n/jjiH+i89CRY
rMeJ4pnkkiZrZE8ftBgiNNA0fJrNj8BaEu3YgFla8VKO1fxwk2ce5H3urcZOzA9J
V0G7+xFFpKqUo9nttNqqBmH6RgVRoF5jChYZJ6OjX5EKZa4DJ3c/+Q4PXNJQ4wrc
X0bJMVLSXTRmllncIU/nKJKs1TGEx9z9Q4qx9L5m93qBbnqryepjaZ6h1QaRBmjn
GwwujMskaY4QKMAajNEaJe6PV8j9VyP4qglSz1YtMh0SeZJ1m4LEWJEN4lcPuy84
nmHEeQCP5I+fBaOJ9So8RxD+tMRTYU44mCMDbDqaUVAQ2SSv+EueVhRBqqwHpJsg
5bgnGUdEK1hx8vl3E2GQm0OibGFqHj9JgtQBAH7bhAQ+CrtW6ac+rix2bjACiboR
sbS/njou5ksteQiArF35O5AjR2hVTxTD/Lazew4+weHBeh2t6YbGYlZugq7yWEYP
6IIGrEYdPYkbKXcrWWlHmKNTfUf/4KA5i5g52bssTN1UCGvUeoKzMHv4TXN4/oFw
+Ghh9khOnGm9wlNmhemQMgooh1Dn+aov8W5vHpqWJorD7yzhtXZsR1n86C0ZEcMi
jo1PVAyK+X3Wbwk1NHoptZMBlBCXHB6j+IjBEZMOHJ3oIjMJxt3pTHbOtMtLxtUL
GFniTGyGrimD2xfBALdDTb8zHARZYKqFGW1e5azBKf+WZGyLxf0mIKaewMKO6Axl
fN2Mcoqkw/8vaEBv5b371PwMdhc7entU6Ny71q0Jr6EI2lmaEFiwvEwRp8XssgYW
Yqwswwir7eqlGumNgW1exTXHg72DicsB6uxJSDvnghV3mGj3gU1vqWaNMx5du4uw
O8CzqwnoyHQFfeH0fxf1OxDL60LzLmUW2sADx2Q4Y1dCXzsKkoFHPoLxNk5HhBDp
czyA38BUXlakqMJdvgPK9QOjDBhG60rgkK5wBxI4t7LdxxECLl0jXyCnFqYyxx6L
rkr38dCki1GYqgU5XlRd2fahS8wrUGKWasQTe0rmmqQuAsZuEnsGA0WxnmqqebFw
VPdjV3khoqiiiDcpL6eVzV+tXLYsSF+E2guTwwPtakSF5ihvuBhvztOfaok+Zzut
sn/6a8bAJFtLbM1LsXV5RjzmA+1SFX5dX0goA4PtcR7zYdrU14R2oYpttgYVrBuz
KdkMUZmPkZ2iHSvIGP4NtSFaEN0sw0ZY+blkf3cD90wDIXwCeu9pntJZVdw7Gxec
WpqaBBh+YhCakbBSq4u1f5e12H3EgtVZWXMvklGGgWb3OGxX+yBZs9EVyGv454uA
pqweNCTE1h2IA0h5jeHOf+pq4JFW1//NysytYoz0Gczps6hOuuDlLl/wFwlFYDgB
bZXcqlYSAixsjCNDE2kSOXH7eZel83Y4tbEj/BlsmRxtipWcDXkC9Bb6iTalA+gg
WVrm5m6AlLpnR7zb0/fRanfTXeUL3C/eYvnUntJoc3MdzPqhabbICnoGl7hJDVJ6
P6AgjC7tfclR9/frS5MYe5vNVm1pVf1qXH+krAuSwpk/zdCWN/trSyaWsiI4mCJr
56kP/iNcp/4O4hAStgRPJUcsWfprBlnHSv54X6kr4G5Kus+Colh8ymmpkEPK+gmG
s08E304ZHYyikDdY0fA2lKkZan9EgxXW6UVXTj1QiMgGyMa9ZXANeX7Gg0d05dK5
Cw0pfUG7X69GKZfmKB8j+qj40lGwYK0Ikb8aXTD4gz5KTfi4mVQ6kyh09v/I91qj
gP8kVxI8wj62kR3D/GE4mEIxhryS2ibOk+EY5Y++VhAP8GfrT8gybmZpvdLyGBGG
mKALxli/eqUAUZqN7dwp/xZfZW4VbH3/ktqmtCY4e9erfMG0Gt/ITXHkyZtfjUKI
IceDRXrUrG9M9Kpw0DT6jB/NCUR39ME6uXeYl64C5+YHHq2WBXPLTnZCfbdFCVNj
NsMR9MET8sJiUeTUlYI2UpADEtkKLvGhZo4q9EndyZ3DcH0Q228QPfazeUUFbenl
3z2fPC/1bC+vk7sv+J69PGxRdwpd3zHq6eRqXgWOWjd25FqE5k/KHI2EXYq3s9JT
Iv8p5/GitBDcYwwQHfGdXJ63VBKhn5FDHdfqzUOMvWwBTK3zvt5NUCSxebKYh27K
bCGJrYRuGqz92f7ncs42wQxfQTPgnEECJr6PZz1SGx/bn0DUDSAxX7X47l7Dk21W
bgAY0rkpVec9yDK2kwZMfcL+DcGBDb7CGaBBZWhCuHF+w1HWtXBW+640zlkSTxps
mCbakFE7Ve/NlA04jVRUHf5r5wX/XgKuJLu9VIyyqonDqzcQZGT/J6pCaKtMqign
HWyFvlNBTEJ9pOLYnznoJMlEivpU5iFIs16rvtBxQDUZ2T7OnPYL6f1brLqdeFzo
fkaaUuB6Wh4MmGoIRiDbQwjSCRDeCyA0DFNUFpixRh6RBRCzg7v77dEb/i1QZ9MS
ykLq9W7Q5Vxb7/vtmFkG8FQxCGDPc6qz4ovB0BAUkvsJ1+Ap7IFDUrFcUZT1Jtit
9C+U3uxE8EC6wAtJsfDwM7K0Waxla+PFofsKvfJFwKZUiNAIHNXNdfWyxQKPHCDK
sNHEYkv66vj8pr7VHu26u1MHcrshdbPWDEVTY73wWwaWFL2BU44jpMCC7ZWckeRH
R1DUlB25S23U1763AcLgqgkhl/VRm0BlDUfN6h48S2zKNfnn1I8YkY3Q8fxjZSXv
YUhq5JvNOWRVFXNI9N+gXeqnRNXYdu6nEOuxVP77RAqeIsUTICH5oRkP+oQ443Ll
hgvt2Uw9fmclQzXc4srbST1DB/IUyfYVBLBGHDI/a6mlCN5dr1zfzElODjWhZZxJ
Jl0KaUDjc+QK/LVLInUq2QjZXEMs+/0hMLYo1UVavfmPlt6WQGOCj99C+VmfZqus
wOMUcYe3QNsXRoAJXALOxiPYmRrqIEf7bzwnVIvFkc4xhYtd/V3t4tu1CLkKFUTH
qV2kgXN2HtKz3MZGS2ux8dfbJ9G3yHYvbWczQkVGcsNZ8t9RdqLdkUqxTgE5+nmm
SohTef8l3hbBYK7GeqxdmX/n4wEG6NLCwH9l86Ka0X9ggBxf6Sl2O+El9qsj473Z
CPDhFFdYxhl+ro069kdwKoD7UUj4a4eHE32P3joJ/UzfupH9WX8exGjwtNmbl9Eo
LNio23oR/TyOcL2kTofEMwtzAsvWfGL4qMCO8VgGFoycwPvQQiO/tyhzglQhy/hO
wUC5RY+3Q0k5rVzljU0zwQE4AViiST4Mo6cUuLhKIHsDYaJsijimVk/7qhSSC3xB
eb5zP/Gw9ZPPq8FMT7i6UGOJVztBN1n/F4ScjZVvjeIF8vdq+b955jsiyTVuau3o
boJF5Dsow/cXw9QCTpdLeZrTEyzfjxhYSxtvnI0qw6Wbrt6u2RgwBCLtL6gzOXxp
Xz78JkbRRFxCGk2M+Y4iy6oOMCIPdie+wVWEsVvTu2hL9r+knqeGJDFbbT2aT4ae
+v0z+HlGqXts2VYzNa/h8NrR/yw8g2Ih8WnXtYmGluFUoyATByw2qOHzYLrd6/2S
M8talA6Qv0h+UuyI9FSGZXXFLGwicEHU6LN0seEHdLPG610Xbl1xh5HR9G5uHoLo
EvQubdg8mOsRt2tbrFNw1wQG+8cX7/yCrRMy4W7cJ+VTuU11edouWVDYF3Tt90qc
W0pPoDRuVC9hplt5ZjHsUBIJCxrv54Q3I7CqEEI4KT/jMjOzqqKzy1sNYt0lgU7P
4E75JdOtvPzSPj5JXCw7vqHKrh9rrRs9gz1M97bwRE70C7YNMjnTIMyUnBlB31U9
v77GpksWJXyFNUNiQUrJbtIvyWDLkpO+J+msfu1z5dxq1bkLqG+FZrui1ehKEfJZ
2FfVVF2x/RQusGeacySSPRugkCI2SqUx9f9pUMrR0TdqmW6ErW/hrts+Jszjm2kk
PbBMY0JZq/QbNU6mnTZIG4tjqdJ/t6G3lxLjfMIoIxNuVlTo5h+2dgGrrBTn547C
lP7ubZpNfFD+u/w+X1ikmvN/l+sbKDixZ+0MAtpSTa7XAlMYyn7ocpOZP+lYey+V
AKpb8hd31IgObZeqUu8KXEhScztDw3qyVbtDC9ODVKjghiLKPrAuiEfIH3utX8sD
sHkUfo7wpefn2oAevGZJme8YKVJBS3JfPgmUU/zoyxblbp+z2jER6VzSeTQRB/ev
OdZUDlZmP6bgl2Gl2wwm/YpgYdZB+6XNyD/pMtuL1TFlWLaMnP+jvgTTIoYA32cZ
3kcJ51YvTEqd5GrtKZV87IkwQbWFbIe+DRvgEY22toj1yjc3q/LLjuv3XJWc7PYr
r5Jm2+ScB43BOiQnOOmt0S6JZUr5BO1fId65TsZxOtQZ2gwTg2n9Nk9r3pVThGiy
wKtXB/Qe5Drk/Yycb8kV8GDiy8o7B+qF4O4Gt3GPa1jQ5iJ1RuHf4BlZQCJjyaRA
mJlzJNb5EBJhrDi3AgFo0pkQCFwRwr2r08+Jwv0YvS2fK6bXiOjJVd8RHJYqHTsH
iNDo+6Y0C8o4xHVyUGyIh1XJKNOvdDw7sxF2sIDQG5V+5mEPRNDm738eJr6P+jPg
NQw2kdmDcC07KvuDbqS1PXVT4n856WyV2+d3IaxC60cDF9ks5cVmIHWdDBlU+5UT
d0iPaZgjsyLvFPEloxztnxTQJBclgExFcnlQj2KTLiwdokqf4A5LrUN/dNt+YlZO
PfKjQb4WXNiCtr1WDIzXmRhTuN2x91PBBTyIXkYHvRBRFkNDEWBM4CKrqCEZzXlf
kbhIpHan4HzcpaPwoSztQWmhy8cUlduq+sRQgdT0ig+063Fm5zTxI42X6LJ45bfU
Ir2iPsOdQFszBI0sy4cZvLbbOTwvm3upBxq7A3Q/k3/QA88DH6Z9yLcgje5JVtSw
kigv9mOXHNq7a8nbfXcXjBcgXqxHWmhKaopbRBU436ueTF2zY3I96y0vjHbeIVi8
+04+tYX2N9B0n4Vddf32DWq56SEf8+xUsxX+ZTHXMNbOji1GXqUS1YkKPdX0ezkt
KeC28IEiQPEvvK1E1m+InkWCcDpmub25PpiSKAp8QEktSEtG7uVVvzpbEY9hRX4d
BFNILghvki+yngWuLOtwXAgejJXQQA1MHGJf7PrWNPNtSVcRPd9sQcX8DBA0cMb1
lKXYpW87Eyn5W9ofIH5X/bgHSdYAil8TPwL9/BGBAAmdPtM3Z2nwWYb2pe8aBMjo
tC63tJljwu/NUUApM1YVGM+nvNwU4/5DVM4L8MEz++dsC5e0K5/C6ENKtzkR6T+v
vbiCgtrNSjvTHQhAquVtU1EcR44pi+w0aKsmmMFGxJE19qry6/bH7gZGVwk3DvjT
ZFwSdmL/CWBta1szu4/jvLnJBUsy952XYuxq0/XqgH7TMh4+5XMaZbn0v+LvHQBb
XMboFlk7z5p392cmD1hsr/MzpFU1/2ZHbeY3NKwWBgVUpf9nP64YIg6Hqg/wU8Oz
3Md3pH1l1vv+YbcnMHn84HLggKk+nZFRn5LCO0MLcNqXt58OMUhTe3GXfCEE94dI
NP5220D7z/tnCT2G1hcE7JuEazk0JCf/8en4D+9ELdmlKkLz+alEfLlCwUObLZNl
eAhJA/8PdtFNnDGcw0DHrXvh9AUSnyqdjHBMvKxodId/7Mcnn8FEIsofj6k7/iU7
wkEOR3bRlpPCLK9+IRnV9rd2zB6aQmhlh5QldEpIyzaXsbBX58j6xsQV2NJNop2+
r10LURTQttdT7u6DkneXHVkXVsiryRhas4hQUHjb2RQvuUexpfnGzCFzpF906trA
6OntLXsSLn7BLsUW19LGTPTfiknO4322+FLk8kLYO8tV2QqhBYer4wXS4XEd1oPO
hfweBoA6eK/FXjBkn+REC3NdV3tUJuzDqOxfkSh58xUX7cjrmi60mCNVdTWwQVwg
02zfKPTsCiUUaApcibklyLRYQV0TckrncvNuLMSmNwbAcFndoWz4MTQBbZSqRUwd
l0qHKvDqKt7ihpbb9zXYFLFz9YiSTI7JENV0xuOQyq5xv363MXaoDT99EVVeZ/lb
bcC4ClF81Q1R1P155HI43KvWIVTenEg15t/7TghuX2XpcEL8TNNBWbJm/i6zJfo2
jX1uXq582W7ccWvZUjMsEIlc3rEkEFhbuZT7OfpuG7fvx4if3wcxfnwewkQCxNm6
IU9Bs6lo02DDFP6+rPCkL0/gdNqFbie9xCa41o+SqqLzipwa4WLISei+Pls0R83q
uGCO2/uQ9w5SUOSB7GEACWG8VOuh2l8H0IbHIzbEroNMb7leBnseHrZld7g7/CQG
bW8pg2hbAUcFHsb2IclSJRPM5l99D2arj+U9tqAZ6+ECTfYrquWy6FvRlQ7EiGvF
PWTDtbQA9DfjpnXJEt70KzQmvtwRvKgjf05A81aMeoK/s6X20RV81d1nuVx5vhMT
Hjyt9HZ5/4z7PlJJlt3CB/HcklQQeQjK7k8twaW1mRD0VtS9b2t8TnZBaLS5k+YD
eMCM7syhurNQgncYbQaS+psqUrPcnlUklD3pW4oUcnau3Vvu0a/4xGgj2Dnu7Jxc
+QJgNUkEhYGTz5GvfkuDCOWuiHfQiJi45Er1EtNiMYQoIU/AoNSx6EwHurj+al3E
tHQhQEQubDoIo7rr8usu3oTKVxRV/F5n5GqKMTy4wj+S8w4svU4GQw9BqFsb5RdH
Yqapeu8Osw+p0M47d45gfYVpeY7aooX1WtdptiEO4yMMjRg2fjdGiiPOcJL9CwK3
LUCk5zOQ4b8BjZmtOS2qFqej707lH3glE1bwAdvHTFYC3keFNgxUwiVY79SD43i1
PUprQDyN2bXDjyEC1fQZXiE+Wu7TlUNpWCYC1jkk/CanO14FZg4WCSbcKAjYVWwq
1uQbF83DhNzrfN5fMXj6z635RVcMEnLVqtucdVnL13gX/xEHgWmLSfY4s3HkaN+L
LYzacL1KADXM3v6LHJypiPfhQMvnSBGlVd22AeHYu0t26CLOoZ4vM9iYm0uqtGpX
1R5MEVLb4OqwY3/QZgvFeZBgF0Ibdr9gKpLAwKGRYi5PWxPX3Pbd5VTl/fUI6puV
8fibC1dgxXki9R4Yark/kxlUq+OZ30jm7B37XNLV8IPHn9eHpw7J7sy8G5kTvQ/W
+YIS5t9giNCGwip0M5M7dNoqE5kmCPC7uq6o4m7S45P1tj3fPBdZAsH0PRv4gvkc
Rkm/7ZYOl1VUD1RfGFQetu3cRXSYHUkFg61VK00bHuZDfIl1L6fGu5wqdLUR6uuy
7MCrBnbi83rXfbU2ZfNTAzzh+VOE9uEx9t/m1C9jfm881AHuTAPcybJnICG1BYpI
RKlzE9mm9of4JoD3TQ1ebvZXi5n5htk2x1ceXuXA1kR5zsatAs7gHDLRCcjKJ3Jz
HMkvfyDg9ENvcTrSpcSHPRKRRvur4e/+msRYqbvgiH+5xQVPo818R+qLEMQJQkgS
1mAPsEkTupApINWxiLbvpj6wTbmb8LCNfqra3yvDyAAxxYmTb60KRL4WbGDu/bkI
jznf05I4YUe73inOxExeTcLQzfCk1WXUQK72fpts7g+fl/tpesed0RYh3/nYj2UQ
oL5lfJl0rfeHVD0Hqbhvj5i0otvMfYIBSn3FpAqGIvHk7TL6y+oSn9sQqH/1vj64
UEe2GGIO2/w0LduzqEYq0mlo0IJ1XpxTfX+ySnP+fQ4sc7M/LaGGqKoPK++Q5tN+
5kFclwu3uTncKwQAJM7AK6phIwlxz2ZC7qkAzFrYJ1LJkLTSesxoCO1IZC5IOC7a
zHiWA/z4fRLe/+HUL3XpP5jDd0nesI+DTH/LUIOl+p/s8HdWPf/Dh9zbFqBxLN6T
pQZMTBeRNpeFxj5E551+a7Xw5pNK0bOO7MDF68pFV2zKF9KpUcAzh9S04ZUG/uvv
0tRYuLh2jI783aftXTrVmqKNo2ltS4cB6g9owrOm+QdXKMnLgYrrIoYXjrhCxuYJ
rVm8/+PFp9OjDthlMHX312A0XPWRzQxhdjVvQSDViNS4/XkS/xQWjxXI6fJMXPi3
dXZci6TIAoHXAiK4AU6LiXHo78Wf5+22cuX8MpBADf+mhh/FHJwsj+eaqQHiRgbH
KGjeLoSmw4w1hab09zHezPLONLvK2NNzA5JEiBlMJLdioXdBKOmstB1QnASAhsdp
nlqT2mWChWUxdxLURXyi0DRcjmmi6d7Ah70HkOdNpugn70Yano0/yAmo4HshvTwU
Jla9e5yp+MXNVG1ahgbW722QFvDg5E1DTWoF7w3ZPcX900Jh+Y1nLLmIKaQHOA6i
UhE8s7dyggiuKDwewkhiLZRUsKhtRyhqHMilZVzf0WgvzLmlYtOVQrBazJQII1qb
R/9FD7MWfK1BtSbIO36Dlib0AskeX5kVGNC+mlcTASYKed9u6zpVw86ERZ27Nw+S
g/FRe/BG+MXaQgRpFC8qyaeUQKDiBm+eppNjYMtjuz9Oh+VeYC/Rw46FIN3VC9PS
keoleGNNBxl/k7jqAtYn8DnbdSp8bgr8qdmtWcoKYLdOLPNZXwGmvwHzptQhTbeR
Fu//Hbjk6DUxv5+Q7dwNf9RaPudaTDyEPJ53T+yo9noi3ZwPK8Gkg1V9eq0las04
APK6ggienOV1vbOgNyWMXs7nrbGMrvPtb+5SNBaKUekQ9drDzkHjwIcvusGN9bVC
uRSY6QAliAWeU6oSkQy6yj6swzzUy4vrFBwiV/hTpC7KsoD5THhczcPiNC/jpSNv
dTlb5oEnkRzrdz5Tu+vbjiRk/eYyov5s/R+vBD0itY2edT6lqDVypP5Du2ViClY0
LWNOc9d8JgAU7I7G6mlnvDYMWBUeRnPD6Y2W4qV4okJNWs1Jh98idO/ix8MqliWX
h2dLPVLZ9aUMxklfSx7v3w9yjro4YeznJjp2z6HeZLzmo7WnjA8FzCyzpI5grJXV
2kVOYzsxGTAvoB9pENeT+SujKRgNN2lgpoMKwg6jhVZThc22+Zwc28JMy2Y1f2Ek
LJZZVziSZzU0h40JDpr2ruX8dg3ZXj5HOKLFNrpZEmOYXNwOAHJwIG4wwi4nYriG
gp70oyOSsPgeY0rhZrm8bTMyYL7Z0ecvJE+Hf8ZIUAD4TzneGr6FiUrvJEjVreGz
0SQgO2cDncCy5lu8smTBEPxXn2C+aGVhOa/6GmXEte7LC7qvWxBY0Y6Y59bCYdkw
heeaPkk4g7ofAzjDrpT3Sn7UzcFygoGxkZ0lcHTfMm8CN7wt005d4hTJhyGSG55X
P5tqMf49KKVf8q/rhpfO24IE0O6oASkYI2KD/QC/J1kYtBabR99BH5Q7jDkL/g2I
ywyS8EkF+DxzXbDjWl3WXUvXtoFcnBJZ2M26bKTyPh8OP03RWjO8q0P5Y41HwIZL
9ZRiY5NwwQkvjzV+q5v7n8GJMujLnDQ3xbOiGA9Qn2wgO0Nufzjj6sKkq8p4ziLG
whaLyzkbw6JzW7uPtG5IR/0QicR1onq8UGJAaFerEFHHZT9Bf6ejGbE6oos0E9Pj
SWhh8H0hxLIHtiia+nGbBFWMGj8Q6fxhKfemdUKYoRL36or1X2qe01IvyJJrm6kF
b0IW5bnpmyII/bjrrFATozszGmJphcV+hA/5OIbVe/oStGJy3ljTgjoFCsW722jy
uXTMaMUFoJ5pX9NiBlpZzindWPGOyeCnggIeRc5fBF57WRBklKJZQwUSREvS4MKD
r4k4Xdp2T3fBSfGS3+F+xfoTH8MvgIblqiV3PYVJktreUiS0YwHMzSpPDV2oZoYx
q0KJ3hLslG0VRjvQkbMz3aZfiT0GCGzm+BSm/lZZbjqu2rf1hN2rwMPv5mkSxwwx
AttQErxg7HrViel/6hzw7apkrJQx++LixKqkerH5YHPNGZHi3mtI3drxXXCoNd0k
+FnO8bqGL6/5tzyJRDzkrObsltKAhbiOMMd7NeI7/4W/8Iod+/dX17yXHmx5rzuu
9oM9ShuT1H5swurXX5FmnkI3KEROLDtPOLwRC5mNs7AX3+7si18NZf89JbPePDxj
u5kY9ieoK23HgVE+0iRJYj8viWFFDMT9l0+sXBTaHwBW/CBbRKkcau20Y8eyClpx
LKhRq58k53hlyxbxiWuZwLk1Cyms5Jicv+BRRTW3/G7Eg//e86tD8bd9FuPF2oOK
TLyaAI4KTAt0PwYv9MByRa4GpBSWk0wN/OyRjV0H/61HTY/JltMLnlo+zHwIZ5rT
NaOdzPy/rTEE7otp0Gkhvdp2KgcvWwU6tqsWWsKuAQEsa4ckfR8lrp10KvEpjBY/
WGkP8ShWtdD92ICBrjzT4M32X5zACsMzFl97GTwwisHkwoyWXmJe2Q27wrks9MdZ
vNOoAcd72Q9PLQJBrbf54OhzvpTgqdCYO5FwTUsA5aAY16l2RPyRfFMxp4c7uqEv
SRH/83Xp3f6rdW3O6WKqtlLMhEeNz1Uno1ekBAZQexhMvQngjN0IVjX0xL6Xa90g
ee0pDYJQFDnaT0ePn++R6Yy2wA6yWmJO43xWtNa3x+QH8hMxYfYdbQfnOLia8Amf
55EhY4ysapcjOkVFzYPrquLbNi3/XoVkKDlfplfloujEooOZeeOsvEpqpKcwlFGU
ODNT8FLxhAM/WU8cy1a4VwJj69IT+BxdR6iFSykeDSl+Eg/MYmbNGJUeH15pkDZS
ijKszbV54PvflmS9n9BbD9qan03241VwakufffqFalas7uDMrQ0i1pM8LARzfoz/
2wLpK/bpurCZVRuTxTRwRkIWWYfAhQ78fq+Qrl2KN0rhe7iqDXR9eI4mcJ6LgmIt
Pvb6BVP8nN3ThqL0ZcO/R3adb19EbyB8xdK2UZ2KGsLUCD7jzBeqecSQJk87ihn9
gP6F37B59EXLD+pXMV1sKRhM8aSnQhDWwj7FmtvfjFQJOBNIoPyVIFDaunDS37pJ
ZwD1mLtU8vWGtI4yFh5ouZWYYJSsH85tiBXHdVUfcp9/LxwLTfJJXduSpJC/mMuA
XmOWDm4mQbmDhUX28l34IO5Q5F/Q6V5wCnjcVQq9eyD7sZ1rVyAr+gUlEN7ctf1K
3xCB+CAP/wiZg4ybdu4t3Nu29ASMjkcBWWDScbXhKjVDJxxAwMiTJKBFdvPSzYAj
5DzMpcYSyPZlcJFBZRnib7M9vIX0+336Y9cNCCxtBxDp5RAP4mswgJmAiJYNqR3A
sKMAhuk73Cd0gAg3l93CrqcIY1ZrtAyx9LmM9yINjt8fX5H/NTKdb+qAB7bhvqJm
xkgf0stEv4a+m7IO98sLMLR+6FWe7GJsyYot3GJsl+h2ZBelxApxG57KEkUPMf3f
F/AVc4c618LFesffFLZfIV2Jd2lnx4LCj1g4+8xTiBlYRcbQwGfoUB5x5CyHY6/h
MSJst+HCEzrKI54BjgAM2KLhA00lKQcWnjNlE6rveK99FtdDCZIi4q2rAmVoJVz0
r8wjtvfSSLrOrAVp2QejIw9YmjBKjl4MYD9M53vNtyQha3WJE49+tBmODCdXNJLG
HOysOTwS+J6+lDot+n2Xx3qVYJFkmdlVSah6aYQMqpuWH0/Evq15Ugq+4q0ra+K7
aoi/1lTQfvlvN9TZDCD3yzx2RI150y7hU13ybDgrQ9ssiACGDkqVivh00v4W5Vti
2Ddx8bdg8tKQNwwgJPe0gP8nYayNUBVk1NTzn5hByt6lvK6U3OGeDHDgJ9AXortF
DR7r0Yb9+a7LhLxqtDn+NVVKbxTNCBs0lleDlGvRL/HBtQOO3W+MgjAl6pApncJt
qyE1npXqjX/xkM8Pi/nO6jjN4fN9lPbE6ry49zQSGnlm4aP3iOR35ozB+m5Gwxab
gdPVOqg6CEhP+7vL8h7fdNIaQ9uStf4e9eGPdhcRQWYerOYEzhLIwZIdfztsT1K3
N+vGWBRNRWQewez4x35gXCKQSwHaRZxZ36VDvrgOlamNk9fyp7YpUhUA3Tg+Q34A
G+OCd4U2gVW2vjknxjFlrm5FnjRxM35fCJtPr90dgzbUmnbmzhz2+fUPjah0h0nu
Y0IoqpAE62dwNYtD0lQWUq+KEZS2I6wCeN8xv+FpawK/E5jAwGZbjHKn00iTriKW
jNs85j2o/6JBCZ3kSC7xQV6SyqTBkfpnhr8Drwc3XZq7fIxPfFCpwVZ/q01uXItz
pCjQJBbQQz5eFYDRPM5uXzmiE+9Gqiu2qT+MqmtxjgF97Epf0dRri9e6z/CF/J5V
G3Xi7ip+ZlwJpbKUMXNXroSFaRX4H8QxnkS5plhuLXzk8mijld+fj5fZMAXDgfnA
G2XcNpb/TG8P+m7UMI71nvo7oq6yaNybn4T8PeQqnSshm8rYLPoo4616ZqGD5Dpe
dx7tpRLlZrkndqTXFPnatoox3YPBlaHSbU6zqZ+YLyNi7ZEDs2WXjBQn1Fz+/3+D
mwGGZljA3w+63cCG1htMdEqDYveBgU80pjeeCc7pbWBePxM+ZuRXuZEY+fFmeWuo
Xxwvbs1wFOMheGgphy0RHWfVUx5uaEPLFwfjNdiv0vtFvVbvOi5dhsgNCqK4b2uo
2ROJ4CKQ/Scm0TZl3wyBlJAmt7vtOTDn8sUEdFPgimKdRf1fE+EFvZ9filT1RfnR
ut4ms4G8iGOUiB/UeKsighjmfiBMkftAqN/2Ruf8aFz3bSWD22nuwELmNmddzl4v
mEODSs2KAD9aYWGej+Cbp3q1heW9FiEg9T9MBU93JMcpzx0SMjLzgselYG86hV4b
cP3Bc3B8qgg//PdHXbB5Ieaznz5yH22rRVQTwRWb40hTScG3XKyMbWSBNnT8lyCf
mtAtlREIw+y6e2w9KDRc455aH8Rzn29RU9QPY1JSHjWv+Wspa+/nEE4FuC3qNc7B
+7B24vVFa9TFLFIcjeUsXi0ACQsoyH5Yw3/tXE8LVOeN2Ey6wy5AA3Uwv5cn/ldm
MGSY+u57wXcpk8dF88To777/n3QynFO8Pr43iYZer0gmdrp3npyB12AhroI7MgGl
MxKI3DphkVpmYy4p+LRurN0dRl5/uk/RkYUAcJwfhprbX6qCGDk8MQDaRot1LfY0
OC28dIhak36beK7/fA1Vr4Rwy97wcXcLMwkKq1OiQwhTuCOQRaiMzx22GSl80xgd
S6SQVRGPKknYZ1hfUwwKSWjjcUEHRHE7UMV9rwubp015tpZCRGGzVQZHhgbSMW+k
vFZ7h96+zyHxzS7xMA7AcZTj/sWEqOE8GeGA3WOCRrNW00sIgio5LLRQbe01hCoM
VjYiH89SkLEajZEaqeu855YAlvEDoVDXp9qt5UJoo6FwUB51zGYTBLvmnKeXDRYG
3buJ9pmoj1EMg5qEU92p71JycN752ZFQq4IXSDgc28GAMvo4TqJ0a1M8vu82RWu2
Ikgr5gF5gulMyQ6GHGggKxMmMlphobLgA8fWJ5bCaQ2kSLKGbqCj91UZN5u28BQd
68Ne+d3yQrXE4mx3I8YoA7x0SYy/kNd7IY7jAalkSrqXLU0XnnXUd2J6lTJ+5px3
f+dkgOJldpAvFs8+OMyYHkumtXRL5o+dclQHwkIRLganiuhbYTKdExq5+d7KVyh2
oUQbiye8dAsMOZRLDS3jx/xVqcMvj1sa7dVjY4IMJdjnTIB+58e8OdBeO+Z+Plmr
mtb+U5aOvgCsQn0lbVSdY/iujb9xdLHBfIK7Lu+B+Ug07d8KKn/87JJLCLb9M3En
dxDp1qfO9D7x49lGE4E3msD3j8uJt+3s4+a11HhNGRe+TxX2iqO+c2i5z6K7BBFX
EBY5YoqJShE0B2iSWJEs7X0JFjqokkSPnF0kFI+NNlfqN5Y1asD3Fe/CxL5ALBPN
HgSM2xUfMwUMuiB5C3rllyEmrROr7jkZ6D3qSaClfRWbSZtJMnRNQYZ0fuagEpnr
syq+u9EgTSryQ4MXv1fILrgOf1/9W4HtypdSkgxYX4c2JUp7SyE4jisKbe1eMUWb
gBHaue27uTXnUXUpx8tMaQ7DUleTrBMk4pQd17vz7J1TAEU+VtqNTQtEJV5wN/Ot
tjPsZKX6wfe6E/VNAMAADkZS6Mp7MU6PuClyTl0pdxURUFsaqdCiXBFKcMf49nOh
crttN6uN8OzTyKrgVMogh78luqCBV8mD4pSdvdHkW8s1fiHEN5Rwk8tP59Mvb/fp
vFSOMwiozNZjMlV667zutx6YYEiXAt1iJEP/JVG0DjJ3VD2r7luiw8U0DCDhHCUr
UmRVHJDDV9w63xyceYiHTAP+VabdwUy3FLesdZ+seZPLgi8m6m1wRk7OQE7faT3p
D2B6/bRnSE3XzG1hJnZRg5wqA8HNIE/ZsGTFIe5w5G+dsWQMkOyJ+FzsL9vF4IM/
p6T1QSopZAuIjVyeUXUp4EfqjtVK11R0o5ejPQOhWnPbNCNDwDZ63LF2Eq0WOYm9
Zk82yOoDpgrStNkNMjIVx64bBhKNWB7hlwfs1jRdZDg//Ne5Z5YwUNYLB2sGDIeY
jyQU8ZK6hvPG0nw8WB9gN1rxTjmujYpToNdfu7CE+pjT8lrQBlkYcGnOuDeAS972
IZKkiw0mMIVqALiirtqXMGLVWZZs/r26QmWsqgF30Ux3EAbR8zf/MERxNeRt6xVH
q44m5hhXhDf/tHhxnlpj+qdFfL45qD1ZjPUvasHvHCSxpeueSi3ZCu0zZxnVVg04
4VRqPeWAdsJwTihR5mC2dX80PysWQkVlsbVKIB550Ny/QVPkEqJfhSyCGzb5knPM
BxoC8qvQR7ZGEzCSR+4jGXlZ9EqvNIcBgGVqFpZAEBjAszO6GCi+MnV8/XDTgAyA
MjZdyWsFfgLHEFveucMwoDTNJ+5aZssO5L4FU6xc8UQp046U3IcL+NBMU/1yWXlg
mVK/9w5aZZfSNXT2udMG7qEC5WaxlTuN+6yIl1xQcYTeh2eGy8O4opEeva6HJM7x
tHiW4Zjuo78u6MqoZ15VodrLLH/FPAvX20wL2aN9/Np+gaicWpLs+X+QfumC4e6W
ZEqNJvYvW4iM4ov9YDoHZKsj+MBFZrT4eejXjXwz7vGeC5MQr2Ki3oViByvDMpAg
X++zwL6T71vu7yKMOY5a2rVhEY7g0jDoPd39Yg6ZPugNJ/t/hWpKC5b9KhWdOrGV
g5tgEaiO/4OZ03AXW63Oh8xZtnRHJDPgKhkKzEClcMRwKARINhlPtJIRhLNOSUH6
uo6v2d2iZr/ZOkkPt971QyDiHZ1rifBEan5lVbAPXScpVXImp7upUg1L2qgTei+L
Zl1reKx5ZcDoBcI5beMV7cVoKNgu2PZ+65eQRFmrvFq5LV8W6aVCMBXk8XXBJ8VR
U7FXJRGfPma+dmtStlPDP98aQs6bptKJ8RL8J4nQRQiRsaeAD4+ep+08OXd5MI7n
yY2I5kZCQQpog/SfnqWBbszhGLQkerHjwQMDLVfwNpfNMtPyRtzr2/i45rjUPnaz
zqcs6VloQnntb+/Wdbf5xN1XXCmH4kIJLja5ERZOFwkQzAwcXUlsIPBwYXsQqCnT
PYx7xqLp2N63yDGU/K6u1qTOgEgezVFj5VxSrjHYBLlYN0SjaJFtciOl3nOw/58S
4+SUnDE54Avm3awTsYLtowmzcS/m8atzPT6N0jddQlgpvjOX8z8g+OZNePF3X5/P
Z03RJMdfetub5KYhhD/W5wBAWocNa+xpTHI3JQlwYhH8hUI2UOodrZ8Fa6dO0/4h
GpLbS8PYb9OHQJVE0HGY9GQ8vD9wUs5lMT4XTBTTOD73Th88BqeSqsP86RuKuuHG
7d0h0W/i0zfWvRr2pt6blFdjXljb8DokuTDwdKFiGNzu/0Y+UrJJN7YDGJkDAzzI
uE7yyTp/LbJQhFEyGQJmQUiWMMqDON8LpvIHVk3Yx4cSFLe7gYAThed55uRGFOnW
PYEFoQ9vfC42LuBlFvMhdlvQGfLSUJ0tq+YyTtp6SPD2dExlhct5XHKAtv+VZ3OG
xgv9PrfRD62T3eyUKvVwREZwCXNzoNWWDwyaoUAsDffo6QyfFf+wg7vLXMl++6wo
Hf+7sNJbmBHsuPoPELYnUr9o1f3gAbrL8hbM+WYmnC5XwGJBp73v0C7c6N6Wizy7
BmCi5JMsQniEToDhxGKpjZ/349B+8bUxMv7aOtU7yz6U71HWXIASCLbXd2ZTdtix
uloc+dsq6BlYkwLnUhhYYRWWdsltR/DQLMRtzFHseBb3yFbLoxgzH+qRI19O+qJJ
A4NZJMNf48Wvks8Edmq5nUGuDe0oBu+6ANStTwluDoQw07i3JHLiCw1naAxW4FUF
nKp8ZpyerE/baavqCitrI7KD7q2eZOyZOOsCq50ZAwO8wa/+oZ3P4fGRmKKcIXXi
KdT0XLfIyoRNAM4RbguFmIQmJpPT22VlW7Bilknodb3tk5eG4pt/AJqTPqeTSaRB
JQtrxsoerCT4dXtK1Y0ZokvT+74fx1nea63QSgMpvM5+UMo+9d+VDVANhpyP9xIF
CP/L74wl73emTsCTio6UnceYNkNmnMt55cy38Jz/qU1woRxVPDsfWUdh4xfxKZAy
ew4IckAn6mjCKu21NKNhDmWdgG2QcBhjuY0mxuRAli8q2c8dvdiaj6V4u5jNIYhM
0RjjRb5C2YncjjKi/DweC1zMEVUDwSExKMruSzp98vzbqMd5D2/zstdjCIti7pMl
qLmN+QDIQ7Jzw/81O8WpMvmTpgTwJqfUorcqC4pWWLxbNLqStxlAOvwn7ozT0/b6
Hcqys4Eb2LZR5jUVDyESYYTEXkw2KXebRet+BUs52yWSJoQc7wrclqK1JtJEpKgF
Y2FIJisp8BaZYjX1YlFSQu1Li3LhM4XbvBtN6vzXGoQOl/xmgI+eAc2BxbsocxHU
8KISvcddo2Km3dsPBfBq6QsY1tncVopYz5AoVkHooBdTgTRUDJiKSH8ypWkviueC
bAYFilamslquuVNrhGue9kYnlo0LTfyWRJNhI4PObnVuiHQywGAk/G1jkHFSyBJY
b/nJvovM9JeDX+wdrjehlAqseMcfKjCG/Cq0Vk2lR7AvqUoWP8zLCGoQFSRmnaQW
qdcuUV2GjhOs9ZgDVdo6eVbhJkEbm83okF14KJmJp58+H3M71740nvnVpZJ3Cmtx
TKZ8vED8TMrEa6wtnppH970MjESkyiOGjOIx0kMxztfwj5E10jOUe6G2/6Rd2LPU
j0FiGnRm0B6dvOpzK7thGzxuLxoQNMpcUZ1elZwvQutCIsxMtrK4R2gsPfU3PsZI
srlwVGpSvE19IQF0CkcD05DPDUqVGNYnOwsXbce5Zj92mp24piyFD3DN3c6PAuwA
VSqz/UYyxwZsWFAElf2rI5Z1w7e+34y5t3nkeSHQUPRhZmRKUE7CqXci9gstE7WW
QW4msR1WbYf6uRTnrUubrxljFIuQA37nKw5Pi67XyJotqHXebzFqWvtnFNEFqcg7
OxjNSdKOuhkbMReGz3slEbFtxBpmNTt1daONnO+E46a0y/Nn/pyrQHj80jbLhJFv
K2DONIT00ThVMwMuszrN9TCjer+7qLs86yCFfgZwk69O1MAoV64UMIiPApovTl+l
+wJJaKmn8Fd4GTho4elKgbFoWBY2yyZJgvM6YIoFUCzl00gMVLISmEZ4NicrJ+aa
7lyu7+4XZMQ1PU1G8uNRjn8gEyh1sdBkOGrNK+ZinjTJyuW/KY1VR1+ncmYGuuba
BPiQYVVeIGo/K5ZeY9v14R4Bk2Uwb/19/9iI+IL+Gs7j7ictTAT5NBz4Hm7stfz2
MCGh9ZYARdX63ThnhOm9km8UCXoJTwxpI1zXIw9SDypImYcPV6C5Tj5LFx45bHqR
jWDgzHTrQsDMUkGxM3jZhQ1b/x4XMc6jq7WAq8Tzd1DGQkMu1eVQe8Q3tvFmTNNQ
6i9DnFVhepQPWKJRFZAp9XTMz9Kg7hc8Mm1lddhoEelmSVADA6bpLQVK9wnAAWIW
u8HrfcEPtmejguzq68EGrMEhmwyiQCJQDwdGZPgTrNBcx+ifhyZmlrWCvTeALHLY
Fj3Bb7/4z9HN89jfEis89oG+EbAbR2edwJAIRHJJATfhv+euifP6aJqoToXFbUgQ
U3WV3PYX16W09CAQiQse7GROQ+blO3oUlOanl1hxHm/Iu1gDvBkOVrVxqZkbBxw2
BZkTiP8w+Z9u6n0PpD67wlqxQgLRGSOSX8Kf+Xly5TqrZ2Bz2iR/GYOwlZLns2c/
38iH22zwktR5F8NsNmI5G2fdOe8Lqok+bi1LdSPqU9YO6lRPpebHZZK+r4sRZS8l
+wFGfSPyM7Ald6hEvar5NkEgR9w1RDnHv6ZrvHbBZHhkwAl9GtTMK1ND39aZh77d
nppzgVTllg87ML4WySIxhKSfgsHK9IMVkpQBqRggzQN6SpD/VsFZ8bbTKlnhp9xa
SVndrsp2llovfLvx0bp7Ij3nynbfEiR7yqnNblyERQrbRdvX17rtJBd6XczQXOYY
pddQOJLgJ6AaEuzZj5J3UTDugsMqdxXHfSXu9MUOpsbrU9Y/1NI+ACtHrAWukdVt
uvGme1D5Ohj3rvTV0OrrcKV8bObcIB2MjRnr2w4ztM6d0mWzneeRYu/Ey3gESay5
4oKlYCcHuiVcYIjFucw4wlVjSY69c833TmKACVDr2QKG+1r3uLR5+P5ujTFJi7Su
YfHA95ATeiDrwM+h0hnDut4eKC3q4DZbvmZqthbCQEekxTC+odAcH5TsY5rvPyh7
0YQpfCTbls/fGZRlyVBcDTq/EVAP2QzK3d0FQMnj1u82pGQddJv3957rZasFlJqI
F/kX9n1va8XCcm7wnBfE+CCo3x30gWPdZkeSjb7aYrHoE1Rqf/ASdybck71Ksg87
ZYmr17QaQQefnPKItRa4J+gWR8nwtEVz72x49go4oONeKSa6PyZagXqyUo0Um0Mp
kTy/I1qJPh+2bXNEy0nYtAxlMHsWkCTASzDKKhn2rjvbloyJDEWPC0Pgz3M8OyBP
ck3yjwKFRr4zrQL9hXulGyxwH//IDo8I02K3qZbvGqzc0xmDtyiHmbuhGVk4KAbC
eLODHJdBvPm6Zvl4wPE8Bcxm9PMA42SbEVylJXUtWANe0woWDSroHv47/dMbvk5k
PsY1P47LlGeBVnkNmkTZwmVUfNMdg8npo4VS146ndaCSy7PQ2JiYNLiB8KnBulVA
tllyznq3D7ss38ITPmpyPkUMew2WhJgZcuM8G0LNxXcRVS90/1i5AdtQ5DNdRk0P
6LBQr9ZXU7LdWC1IUFug2Xv8ZtUUgSKauk6d5O7Gl+VYiTzv+9i6iu6WFwbZiZBD
VTN/1LQD/04PK4Elb5mfqYql+GZJo/h+76T3dp9wvd/mJkl2s7xTmDPfiDTz8hxH
RhHu0p69keEK8MlrMwH5FGk8g2tVIZU6BWXrWPhbOldLCRyXUx8ECN8Ij1VD8OeC
MbdmAvnnCYdx6A0jlSwuBxnn8w1yvHAA1dw1wPt3UlQorvvbe55GlmT1hQBevIv5
FqyY04y2nynLZJF1njt1fLeDS9Ol5/TpQApmykyT0cOx3bc24ZsRzI6f9M1F0Tao
KSfCBe7ddu1KnywPG6/JoUeCTnpThg4290QkNusOf8Kojaq1frgcnVZyxuch7n6g
0Jj2WW2BRlDyhzag0aOL2sXVkUptmcaRUVZFPB/0/P0rnp9cBxkXKM6TOZC8d5Sg
sxQQb72EaKlOCZd3b1uKLQPZpS5XzWmiL1VuOHrY9/3Jw2FDkIVsRT4xlg+kOmvU
l2/hgGhiU/2GJG85z91pNLY9/3HDmOUxSgFvOjzjY5gqfyxzWIYo19Jzm8c9G5Fj
RHMxH1qglblfOpQ0+fa16ivtlKuP+vIg27Zz/WHOGPqWYVpTCncRYy/MRKOTA8uM
4l7euy0gsFBjvE7zUkpDUbatyYr9YvIW/ZblF5g1PuvFrfZSSwEDfi9HzZw7mq/F
WYJ7XD2Oo4gkNQmFVWkT+D9lm/NO+/0v1KbTXLayMaa8jj+lhj6VFDkwXDE5sqgf
tqMIWIqPUUaLBgKuQ7bfcDNaje2MhBkSHKxJEmkP+G57UU9B/jsV1PIyVGe6r/us
q1b24QL1Td5TeeQrHJTiJ8DDcVz/Ce+M0uDnnM+mvpQ9c1uxLmG35TvDf0HhE1Ii
I2L0cOPjhcMuO1Sl/3b/uQnYu+KQDpppmRjls9V+GiYm2d2c+ywdj9AQYfEExgIU
XYvS7mtJEqszlXWGg9cywF7wGDQZIZ9xzA7+o0qyCvHJtE814xgZuN5EfyAoqoMi
VkjZ9QW156V/Edh3lmLUUNJOLfx6d8qndTfPeJwE9/L7/h97bF4i48Xuwd4xJ5om
yHaF/LszOuQTYU+z+BxuOl63+4D7Cb0JaU+KOrpyqcrHwGflDccEtTeuo4ztAmRf
XHCI28IRGTn5mr4iEikW4HuK1CvK8aNA1yEaHCc/DIkte91CPQJAo8keO1eQPPkk
c0wMIwsdBpf0JpeiK25dajOG3coc8XI36bV64GcsgsG9u+l2Om38gfYooQO9bV+N
J6ZwPUED8ETSRmo6mBZr+lmXiVPEt0ahsY4c2EwX3dQGmVsad6B5vHp7XFtuy4KP
VP17K2oBX2KPC9rKgHO3ZuroYR4buDjc0W/k+6oZVDhFcu9v7uDSfo+v69cudYpn
5ealCUT/hksE06S4q+Hhbhi8gyFC+eyeq6VzCwvGjmz3nq/pNt47o7WNbyvtf+dX
b7KS57PlXyHZ1XkiKyN6wUFgAS+C28cnlHqk1KAE2sPaTLv+TrV2NRL75BSdl2D+
cB/zflhEkjVA/NibbOPC6gPpiQkZNuVJGU81Y5U3NRExrZBBNJJRgS+rk+kJjW4z
v7DUd+qtSqABGmxn2yhLNb0+WWOQDbdX4FotT/hOI3DJJXxo2BJEk6bomQuEarl0
FiEoiz05+oYYxm1gRoDlP/XVsSEHtPizo9Skw3spFwF9JX1/bwxymxdzXqwXX/kn
Xz+SSVxNJPU7SXy1uomVk/b+C3uiA6bVzt8q1TIW9wDl3YKcYJTK3lFgGj4xjQF6
g/LIT7w0J5Ox/IjfiO17xPFt7durRUMchC/DHSqAzYO6grDL2yx5lM05vigdulAM
ZFNKeoIWD9JX0nOA8iP61HrDmfflUiJ2GI06QfdaOnAx5inPOQxme5MoOxRuOc/i
Hdgq1dA4fL/Kmbwb955S9vKi5dUBOQaCX2MRcuSa8+4eeLxHleTOxqPC81/gRttu
PpFkDicfI6wI2Zd7gjX1uCLOc6O6wuXX1v/+jnG4Ub4Q/TtVwVaHe5BCjoAv8jYD
q21viEHAhcsM/h8rv1YyZSZNX3iuDKRYzvWVH8vakFlsooBT+u9E6fltSQxWw9gR
Z/Y8n7ih22hRYCjSYpzLZdJ1VFVhFCp59xbxeK8BaTPR6nx75EJG+W30gnrbErH8
fKgNfP1PVfy2jLIgL1h7Yp4tsWtKRWNtqxUFFtAWaVRGtY0c+iGBCbwiZYeLjHLE
7Sxa9uPJsMcImaxxviUTx5efSE3SNKf/135RRY6qTQR5wIek8pmbIIfO6eA5Ltwb
lJpoYw/8FCP6FX0JeEHZodjZ26C4FaHL3/Y9bYYpCXQCsUaTg2+nPCfMOHmSZvRv
F2X+ICgCdvLu3w2BGbiGLroJYwLbGyqv9RqrdR3uaE0gOdgO80x68JAPdJWLAlDD
tLu7Rxy/lyjhXexoVh2tERbKpJgpvyA7Gbq9G8Fdp2LsdckA92QyoVhHggnjZqTz
WTXRAeUyBZhltJEp0NSDH6391mmIdPlkmfJTLyaRAzuayZgoQTM0U2k0QkurR6bm
5o7BkVf8YxuDUXV/tDCz/GWXYTfOjG0y0rnLWN8+ACrvCzE9XlcyBbgstnhc4TBx
msnKd57OMSVJqDb/cjoWyRaD4AEEA9LW3nhcmAE+BbKwbVE7n+/ujy2ek/ukjfyi
LWrw829HeqPbg5vtVMr7Tzq0B3/Lm/0MhIzIBgwdwch7rfRZL/QLWutMmLOPQvV/
dz42aXbGkHG9Trv1kh7gSmcM/belZ7ABw2hoDUYDtFptd5SJbgLSRmQAJQmmkcKs
/3SNy+cX4yWBAZD5SSdoQbK78Fu7vPDuE4RalFgUP6lUx6d/V0ugLk7KBwclF85h
qKDVYAu/niXWYx+BstG7DHmgJbsGPt00uamrIoaG60mdnndQrBmTnj0un64ZoiY7
4TDGwngL/cE6E+xWXHxFAihDyrC27Iwmm8nwrGtA48VY0On5SIf4tVcU3OtHDqLG
C3x9KSZEG7e7HcJg7aIBKM6zKYlhwz8IkHkneVbYv+RHyyU46Er51jyoLncWBXU9
dEImgTibYPxLPYKcDOfa8V++eLzUiIkEl7xo8G19yN7dApGMl6Lptw00MEwylVyV
CT2eBsRgVtWuluKHEp0cioOR3FkL67MHf8cjPG+hPwY27cwu0b2YeSAB4YWddHBD
cT4HohV4wG9oI0VUX9o+0hF0/SaMllqFK7eNrgsSSMzv03B8Jt20XuH46DW/Gvbu
LETonk9sl9WUZhg+clpnFiXtaLO0FTDjZavsd493/OEZvMFseEXhC7jtpqA4yesc
wAsKmvCC3FyMhatdb9ALIi/v9V4xq7DSTRoX7tZcWpT/VA9vxSE6wjm0VpKYBf5U
rADJp5BkrNgQBHeCqDjbDnx/NJwlSTshC6FjvH+XiMhOewV1FnsQtK9v6MD3LQWZ
hdqeqVYO5wGOn+ZswiFmc2GZlByz5aLALj2fsrJLT0SPvGn8/DWHottaLZhfaO+u
zXAUZidjiYPkRh2GEWnuo+vcQTXoGgs+yB8K0HThprII3PxXi1xecU+n34J6UG5Y
89D5g9pQjogVXoZz5DuHeoJ6B1D5Spgb3Vt6yrp4NJFC1US628XLgVSQs9Ym1PtU
WhirwGxwx1UIMqWOdMb74VTqGZ7MR6aLReSlqwVZLCu5ktCBtt0PVgrY1Si4ftaC
UZeHuaM8wrMgSEPlLsXxbh2XZxxbgsaubfdccTF9n6+i9iMCBR+lQTa0fALAxLwv
7VeUt0CB/BNmqNHHOxNdExbyIx+9IQ8w60CImp+I3AI1+Nk2McN5I+fYHOKFu/Ty
la2TVl2EWg55kUk/cnBD71HjWZ1YCgQxldRTXjF8rA7G4oImj4elwj9LeE/2AIo6
uGS1NnTDSYi9nk1J5ciYL4aGTqeP+zMF9Yc2CF63zwjiuXqYIkpvTWHdshcGx5RZ
/mQs6Rgj8MNsavAqvNzDshzMkMBR7jrXd0EdI+EHqsvgG12obXcEPWd+++YKcvcV
mgAl++inoRQF6SufVBvcVdIgLhiGKX+OdDW8BnPJDMUZtRZyzjp5CmZNOiXmeVZ7
3CnrT2ljZD8OvPCNpFFd9KQat5xv2zaGkWHlM13neSW8U4aNBK8ZnvnwdX/VAIhR
SfHmsPW7mHdlHQwlVTtv8ufQE/7hllnwTYOhMZKMV+USFx7WM8AS4R22DJkHKQtC
OyOO6lq33t6dftLkV75v86DhQEkRdZatfobeMTVAbuS1ub3KHtKdP/y+hGGVHVB3
t/B19ooErNt+a1zdGccLbHqbDA44WcxApJbGYaP2TbLg90VPlSNhgsvf11UQSw2E
9UGOxQXEO6M6ohKcmm38hJlqYmY90ImDYfoh5o/857GsuMNSK1cNjq9IkuPkcfgJ
Sh1ETbceieTnhtZgSNZszxJ+zOuwOxow1SRqaJJy/LbCDpHzzR8vTQEVHzxLaC7c
BhL4Dyptm0920/RrPohaqp6CP3cMrFkAV9hZxUBcvCiaUMFNqEidTPKF9Eq34OwR
MNwVZ27AHHlkJpRhfB3UU91B5D5Ts3+TQ8Q47dbQ6wINIKhij08IFrmfZL2WCg7A
OreWYlnVh+Dnt68Oo9WNlFJV5D0meRTBxLRDFmz8Kmj7VKbQc6h4ugGod3q0YmVZ
s1X4+G1eCo8LeRScj2x8g8qKk0XdaD0eyChEATBqElPZlkkogYnL+dhVGWA8gYqa
kZHXc3f6dt+aXOrMUTbtylMbXiIuz6TLUPRJfhGjxvQHgJUvepkSQAwWe6tM5xx/
ZIKCWASctj+PoJG9vJU/oM7D5IrE1GKd8By0/eawlEWsnQP1KqeVoDTkKTcFIUey
8PVWzSH996aKGkaRLs764R7Z4vFB/xYWYYd2xWmz3OdPOqTjjU0/PbKPa5WWEWZP
fKzXR5nfyZYI7mgcAcBV2Qv1t/2Sc6tCUEOA80xAx2NNupKW4wN6WcMYsNC+MZ/w
JIA+mpKjidyvULcnSPlOjL+fq0hhhaQ0N5LqKYhTjqgBEjWdmpr8sYOequdUz4vb
zxt6ZoShjprhtuQmA9jkaDAXkuhPBAG+tXYT+h1/1m7bzQtLt3CzHDromsOA0plp
4FNPIjythyiX54qLv0hS3YBR50LkVBbKLTP4/FnV8E9eOM5iwe9hb6xlOfgkpJoP
RkKulWC6qSpc3qRacmFGikTUiIFOwplqZLtiDR2NAJYHJv8F2FJbSbLVOjr/4WQR
9ALG5GfAXiaFWgGwMbdlN+D/zpDwn4549o9cvID3ChSxqSbWAuEBvWK30htt4G31
iC6c9ytAOnkk/1rivR+hfadnPNPE5ZePSujih8mESbf2bJwgUj5cpjKNuP0JARBd
uAEVP/nXqKRZTyHlH9uw61g2DLOABHb4bo6vPGZY5PNZINsOBF9Wg+up2ISvzF3q
qv0U2qXf0Aq+YnOrdKw00Qqi4vAd+ZqvD2kSHkVNHoVhAzQGgDgQDczaKbfRGj/g
KV5IBBZcmmIa6CUKRu9ng7LbVm1v/KcVm7/JG/UaKvODCbiJ0eR5VztzaMlq+mqJ
+wosEyAlFkY8ukNWmhkjw46CwdrW1hrK6Edr330BG8Jkws46rMbI7F+73gszdjgV
A15ITG6oYVeXPGojx8waXnedrNjawsKgLVpOXi3zeMdOXXmsHaiuBRfIqLRNOKV0
o6TN/0XovS/tMz9xAnn5VXncuui121B7NT+GWxctqG6Rh6Ld2UMw8LsgHxot7ktf
JBMxXW5eyCc7K02MYYDF8zNXABMBxpt+FXuVm864N45w8uv9RSLTWEoR2Celjtm/
BOnnjn0K7DpBRKYyNO+CyUT82tenJvIYSheChCPOgMOQhHi0ajpnPUQqlOQL9u/9
vJt0eDAbQojUik/YzVcsIV1yKDclaOLxwnG7ckOxH0uTvWhgQ9moaiM6KCUieHb+
63E+RMLM3EU15gnEpDqbKangWkZM/X8H7u7mApSmgrG96cGKsQGdUS//nWBa738c
xHqIavA2hrb0Ey/0dQzxrNfKPJfjjIOZHzF8wFal2FjyDV4e8WLnkAkmi2HmrnVl
cpqy/ytvVc3bc34wKAlOJjgkAU3lcWCURROd4Artuelf7RcrC2+aXbCTV/H4vqwH
TPVNxruD/UnGT1v23++HTDhx+Ycf9LMtcMTddsr8IUhdJrmsntM7XP9JQ/pzPMyS
WxYz2PblvPqq7iw3y3snd7ufiCGFHzdtKmLHhO/QeuFZnJ8q5vfTT574+lzy9dLl
eYjaR6bDy35JDKTO8FeHgZFv5OsAcKZdJ3Li0ecfZTWrlnByYisg1+YRAVgLRA1y
NkR0moP1+KsM0VrvbmNPxiDSHOZs5hPlAp8ANWr5NQBATLuVKqKofmaJD/gtTrhv
kRQ1IIp6tiPgynPc8i0e+mjzjxxAFgj9gR+BnJuc7rEW5yDwkH01d9Nhs3WXc7OB
KnytXKM3PXnz8iq+NmW3k3fJ6IhF/I3vb4pVDQ53jSdYyy1hnnS2QiaAD30UlBCG
XnnJB3Ldy4kiI5yl5wiXEp05R0GTN6r2a+GobijMhccyQoc7C0RUyJy6E8xFpTxw
FD2FaEQ9of7QV9lBkdr+XDYdIpXSFi88+wy6/irx1G7kkrmtjo2Qyn1oKfU3GrFY
rDaKCzAoKTq770q9IWRl5HOioKnbUrhb1l6FL7M0sVR3djpX7Z9+jv+YUY1HbIti
PR+Ya1kThZhcAdvmK6zD6B0c6T5cPbo+pO8BiPxrRYxm8Gb/BJRR7/wURIKLq/PU
v/cOHuA1TUVTuXZdTchBUhqUnTVTFRVJf02DvHWKMD1D3bG+Zkaz0Ni7r6hcVpMW
Hg5exdW4drwRu5o9E1z2A5z3p2fykGrTFzSlc3U2v+G7xMnfhcoCR0Y9nUSx9fb6
w5s5LoVM5+fpYwQKnG+7htKDQvPaHshtiBt9lKtvXuLKg2vhRR+MKsbJE8HxdeIQ
LFDJVb3BTszyNRoB5mdfEGAh9FmotuwEq/f2AZs2UxAW8h6f3BbMbQgSaQ7ojRLW
Ynez9EFn333Fqr+SdZNWYzLJICL+hld8Ol7oWPFRRq/eERPQ0qbJsT5XhsBy9qXs
miyoH6tLwCx28bVhwX6ZkhLJn8j2/+adGWMyQHiaMHHNudGzVo8LHtHYrJMq5UKt
+N8glRMY2/mC368qBG5Mv4lHj2HMArXlEh0WfL83C5WGMnpAb543kwd77Ngr8fg/
YDzcSjma8ULVS2xorXmk6Jxdc3Agcs+Od585wf/b9+TCZTRnCyq1/SPDIge3F/Hf
ncHRNV4KVIAJIpWJOTbahxoe7zgxhP0z34kYUhZ2sYpxxV04V8jErR9gCP7zeUL4
VFNBPMxYHGnMrhLgf4aILl6fVrUpW7c+2IDNbiveDUkZbszKLQ+vus8cEjII6V3S
vf6OY+4J3BvyV0Y2LUwHDgNrwIdoH3Eycg/IlzdkrKQONn7UdHiaK0qxZdfTD6oH
b37BXaYGE/R/rl/kAVcWu0DpjGoizwOBTVO9SUeLr1FrJ71HGg9zF1w+IJmKBru4
e8+NDH9oqiGHp3E72h4DlFZlwhZabV8B1p0ktIPXOzD/95QW0b12TNvJtilXu/Tx
sWqhmcmwwi3MO4XJDrYML4yJdG5XstyChYzUs7u+d6T4X6oOZijRleFxBiMJlua3
Ap8qRbHa2D/2g+ghHzT/g5piprSxm2l+d6NqqtRtuqxL7CUGAMgOKra8B0zvMkwO
mnqcpUEv7VVx/H0TMD4iQPEuRwB61QNxqC8tlSxtBGW1Vv4HO8HEYYg2Dhbc1kQx
2dLxb2DohWSz09ooPBonQ2I5jfzucfkcL28H4ynifRR+JE7B8PxC/ilnEDVec30y
fyI9+4EW9/KBks0cj2fRf+wvGqKN8yDh9rdGtCvJ+b1/W9OCO9qBxld0jR3Kgtpp
RLNpUD5ArSNSfFXkxR11Zu4EB7RTFokBrLQxQiw9xcocd/TE4ud+K0apikmdDn5A
v67NNM0EwUHKNE7iflbxnUE7Wwrdz14FOaKmKufNg9Mb1uRP+W12zKLG4mUzVtjL
zDmZa7kkLLk1iklJzdEr2w9WiZprk7rr6cRODMc/CdvHL331oFdPhT0CHoTlIOxd
uYSsVsPqPYsjL4InWePyzXFFcre1HvvvSami9MU0QQZ0qReagUdSAvYDjq1O5d4Y
W+sZ6fmBb7psNS7G+KQ5xLSGhxd/01yEaCcHhUOpLGGrZFQW1xpcZD/ROmyG58pm
nGfu4RX5ICdAJpXKGmVodmWAjDaMrSm2IDNPh++h/HeFBC8rOoM3S2+uHUM2RnKf
FAkSZnIHF2RaHQ1si38Fnigf2Fdc53oG4m+VkoQ7uUVOJo1ZYzz+Ickl3jbARcFB
GNk55cPPK5hkp3ffO1ZqDHz1NvX2GgH1zipZDntueUQ4sPHIawY6QEoGZeG/M7CA
5xqWfd4K1mjG7BnXSeylxVVOD23RZXbWs8/tdcBOHUHRO8tIWKl0piSzsp020Z3m
PLlguQFuRGjyEWbvKxaU+GO8Q0ithRDObGBp0h+hZRjwHl0svo4fTpiKdRbozhST
96aNtvNykQREBl1PN0Q9+CXHoSVFII97WEp5tJ9+a2RLDVK1C8bcqOvnYXNepbEP
VXNNDE598EQdqqw1Qv0pTiU+9VSnGIxx3JXtEVVGFkWn4B75+zREoz1JnLmzSwKI
E+sVtWE561x9aZLllZQEvTj/nF/ls5pGEQTjdd1gOEO0pQnLt3BvzVvKuoiJQT9/
FPUQU89C9hP1Kq33doWh3/UU3YOKlsgDAzsk/vjOnZR31WBG4BoxeVPGu2J+hjRi
yvit4GHxL6a9pkimDxFRGPBLRPLCYb+WSqKXYAn8/POIhT0KzaGkD3Xcc+2pI8sp
iYw2gwcUJzM5gXyzqZUD69FX3iVlM3iFfaMf5VmmcZcxtltgN0uZaHqqaoMNAhH4
1eX5j8rUA+KUuQi2ZtEiHVHD9f4v0nRKYoHftm0++FLeyUZumH5t2foJJ3z8B0gF
PGoXjQ5RJbwdC0xLJzm2XZ1totBIx1LAb2YqbSyQo65GljtSvMLrm/3ZI3G4su6Y
zDtLcfklkYGnnwdvF85ZP0nUFtQAdiZ/f2GTbTX7Ya+KqXQYlegOrTSY2HwOn0fe
dT+EZUhkfxdz+QfAzTfZygDugUZ1P3Al/iIfWa98Ud2ezK5BefLkj5N36fLsS4lO
a7KS+PXfDflCgjcMrWmBfN1v/XaL4J5DGIZJU5KdjvEHz+2JAnRrrYaqkN7d5MYa
YG4f2C7miVNIcdw1nfi2vvvqUhDrzhtHMG13EJ2HGRaQzxUnyh5tGP5q5ieM3lKQ
xuqodR4HjfbYenuCg3yKnDHFwVmfsfgGSnCPcvZJopBigYrP8lJOikE9/d0NAQ6O
wTcy/EcNfJwh629mzFNDG/FN8qzBdC/2dOOocGUXExJzo6zRC/e6v9WPmsM1ORT6
wK8KIMa07x+05Km2IWvf1hnO4fVcp9AJLx0hqu4kg7mMXNLhx2lllEJn0aATkqso
ZvZxO1XLObOR0RMD0d1xEw2/8Gfmw45MO+AgJgEiG09NcfZ5zfeiSp5z1gkjYyMz
xx2h6O3RowcZOYYhBWkiVUUozkmUmCkESzNCX4TuxaroSpTsptp2WNpRSOAkMBmC
myzeHTHsn85szC8HUmfLGFQWVNuOB9uPH6QP5D8FpwSEFP5zjnJ+g5wpv1vshMSr
2ZdOi2DgHp5TnVpatCgRVLyz9n8NaytfhXE51yRM7AwDLGZfSYGkrH/V0bMt5JZx
e7l9FzRkI567REjj4jAykzYqbpmNnPg5Kic5XCJ2B8Srie32apH48iKj+fXwz5lJ
NTINMqxrq/qLX8c1en0cjHfIMc3n/rdUU+Yhr8jHoloyAkQC91EiNB/fswuB/NMe
NshfrnOsl9mYTU7cV/K69vtcFRsx67Po4KqyawiYNK+c0gBnOuGdzDNYsrSQbOzk
ya2OYDbWBuX3BBftrRcricgofFuDhmZwgD9Tl2S29ymr/CLiqMDq/k4BQ6aYl6+k
TT8rtbZ2S3L0ddj6CJQ/ZTsIpm4gqQfeJdRUnMpEuVV8wm2cbBY3kOKqpN7094nX
E2kidgNjOjY4AfY7unfNADWkZjcveFRUXz2FoRL9rJ00Yb1iw1j0nSrDeZriX+oh
FyO3ijXp3xOou/FOZe5bTwllQdnGe7jxKuV44WtTcxQKwnVQ+xHdI4c3hN7dHQZ6
v4Jf+97gUkIQ8aa+GUNn5MmYJ8zvTSdd4zUhhdFoD7T9jgCkHxmZvdjlYa/W058h
v40a9FVddPub2ApnKXO2PPdiZkPA37pQ/8i1bA96yNYVFtMvRyDBzd01JgnoGqQ0
lgs6PPE7wPhBfir5fdvzxPXBpmOgpopcl9zggbA09JMZ1vA1gmp9fCHGaSOzYKi4
ckZs6o3NxwlU6fZbPOLn4Im4oIiWfjbbDVtyqsgYjID5fXr0VHDuNNg74N/EdfrN
6pScQWhhEtZIYGFVRTQz+i4TcQkHrVhhFy2tI3VoNfTx8TJYW9thx9EUT8eiuPWA
NiyfKgjljeFczlXxMRHcmqr3EnzO67Hxa8LwIYAFUi5mWO5aTp93PJvLSAUY5FUV
IAt8iAh/8pN2xpLXAfVlKNY5uaF1Vx9Cdtd4a7DFWpg7LRbqdCvkF0n/aFk3+F7O
wDTVSS31KDMT5UWCLQHcoLroXs0V07CbSCnfZqPlFPA8pnqy+B4qxevFpvxD0gsN
6RSFEVBF8Bi+aazav9ELCNF2CYpzkLXjOHXDLjgkXYZODWxEBkDdteSgDOQs48Hx
ix+DvTZro55YMI4yIGn1CaWthOXUCx4mmFOnhZm1ldQ0YM4lbh/GOxdVunwKdhiT
9AASUNrEwQn5dkzu1Sl+lLPbC1A6i3C5zl7QImmzk38D6ce22wEugk8HPsODVErW
JITmvqn0ZPrb6E3J/T5yEfS8FF4ntcrl/vUqQc5Zoa5S5lALorAVkSZs6tqKJjcu
eTJy6bhn5vc96Pt0LIzjh+utFGGFWegETors3MdsCM5wEDVFrf+5gaXZAfNk7jPI
JW5P91VbT9LeW4389d2sbspX6HuOA8YrS5+mw6NVd8kQwX9Z5BK5UaimdIYf0B7j
YDgHHvM7tyUTuKvTlAytHVyzOtIStQRvw14Wvs9LYBKvvlUaLY9VboDhFnYHMG7k
IU+dY6LoHHGoKRGWNLHi273nTWwyEkyvq/6ax3n8g9iG8Y3lZ13EM+y5D+URu90o
LOh6NZ5jbrXAt/kIawjoUhDxGRQsPmzGk2MLkP1R/thL+2PGene2SKA/XkFri+7M
PV2mJCJHJnRDuiHmYo9APE/KsAUqnKqnhR7j2gise7hjOyYU2VcWIZMBHpZ/l2l1
MVrbIQSToS81P1/2wGrW1NnDOR/jRSjhcwrwfOfuc5wNDNrf4358e0VG54xdFPBS
bgwpL9uU/CE1nIiDx7ErGSNk7aK7hdrIAR0PKHBmLHC5t0hybSUj80d26JbRsDgX
QJm2GIA9V/F88d1doDMbSztaWtvWSquNngNryjyA02KoIZPJfpAgQuN10gsRvi/4
+yDPs7U8yBh/0RSXLNkvh0Le3pt8PDfs9G+lczAw0Pt1UvugsrCJ5IFMfwTRe1aF
GwV1BJzxobVNQlpIGBUYi2cZIbDWoXQZJiOK3uqU2smqyuQCQkqPwn1r5VZqfOnM
kCWkzRZS/KOoE28nXbF5ktuyWjzHW6UdxDe1JfI1vku1vcEEd2qajiTQppvxA6A0
uHeuMhRDKHJ38LSW3kxwlx9YmWjHYVv89EOQplUINJNo89H9gOYiAjQKBJXfH34p
H8pzmX17TOiUH5RtDh3HGYKegWPN/NZ+oqn2uaoGR5HJUmSMAGyLzPFmyBhf5h39
goHZhDh0N2lu6+q0HmSfXieGIq8QYF6B/MZQK3tSBSzxK0mziJsyhZFRZlInp7fy
nQUWUxZNT65BJ5HMfnqAaWFmNc3A0DvGqkq4K2DaDwLanPp92OIM5ssFks6qoOnI
ckwQioZMwwh3SQV3pjb+77I0WETS1ZxCmwJ2RZz3DOu6poEMWpYy9tjHp71IxSIl
HbVYu4eaFPfZEkBA+ehSvsXbkC5SCy8PmKU4wEoz6G/wGhfnMZ5G5zhIF+3D4fhW
w+GGARhF5cMUOys0Po5nprZWm7MgpNOnl2jH0HDTnT+rknetfwPQgW+NbBZDKhDw
+ztd0IqgUl1L5LcJWEWW/0YUL+SdjdS1m76VsNQOdbmBxWga7XnFFw+GsecicwNs
Jwfvyqw6OFVLqNCXOhKpuWfX7aV/Fx1aHuxzvIzoGD6YPFJkfRbDZLlfZEdKHKus
q1uZ5BaTUKHwwrTwOurzfobVeU0h3uA4TBt71SDLj2Q36jRrc0n8KL5eqItDS0oy
uwqpiQBF+kj2uLw+z7Q5zyzSeZyz+bPoj+IuXBanEzRF0VFbFOVGntGfgazZIyVl
xqJR9s6CSw85VgOtCBkcY3Mk5K6g2vBJjlPv54IoGGuaaPeBNvYYOXu5VhyAmxAy
MlAegv6oep/t7TIiYWUU9gOFYjkh4wkRyddvV96kLyeXLL7YqVVLbe8EwyrK1j6H
LJpauTu54BldiY4ZO3fqa/Wz7mNzBBlYUPpMdidcmPLVScARjyCBXmkDRW0BZ5WE
gsU3S9rlDwJV7b8YbDOOsrOPEBEXlar6wk0SpgPsdDFl+hDaXDqVTVo1cOhQbIt3
9PSdVOYwB3Osz0AwCIo8/vxR1lsyplS5B/oACGj36VpW+q+qQEbwc5cowNmNzDNA
e3Wrmcl4RMGb8MeIugArqFcB7vA7xKzD78YJhxSdbbPZvO6pzot7/V4LO6cav/jl
nSJy7Ed6w+KGDUEF8eU2+omPjFkP4RtJg2WBhhhPAs7NvsK3GCd0y1TzM4RjvZJz
uQheezJd/pc1l+f6Lj07p2mjul4VFsOe5tut65VZZmS2R2440OkmGBU3iDt1B1dp
UqxX1MJ7W5Ip4cOFYKG9WmxITlOhYVvCFrHIcDuKFao1CxWuLdQKIdCO86iaMSlI
fGZ9iTS6F7jSj/f8mVvJXDEl9L5QRjsx+ust739wwsGucXbbnu3uXV3vi3EmHW0X
UUFR92f6+aZWXl1W4xnfW7UctBnQE1jSHm8Y8Gfh1WBpxbeD/ExqnKaxbUyBtilz
Se/pidQ3DKwbcEUWrvrmMOGYDp37tBTwVlxsiDBxY+Irk3kYXwGNNIkIio9i0sJh
XRmITIk6lH6frPc6OIhzOBqUKp+TYQBn1YFxmYqq47Xh+X0JscueD9x88ydZj9me
iTb8JtE6aUraKb7YvF4bENzh1f+XFFjd/KJSvwEJEXzb66rl2pj7kK9joFeQ1aQN
x+UuwPUrPaSxcTrFVc8emygIkN65TvdCJHxnNeG8GuqwX0kYxFuvHeZXoQ+mrFEZ
UGIjW2k94fgA1UX1Xmnf3YP8zA6rtW99o3HKOpw1ok886tDKF/6Kf4p4nEudBChZ
enl2E30k4sSFhtrj6svGarB2aFcDqWOzBg23duW6KGAR2XlYBp1IPvmP/od3MqLv
AMCbdMFomSCz1jxEQa5XIsUxeb9I9PfsIhJ/18OA1s+4SWp+JAjAsH2yqMDL5MhM
iZCm1wsQ3SQNG8ecJ1eAFADEEongfgtR4wROXFyPeNZWqPwVvMiOQ611psGFqiVc
vaNnSsYQ39YLUIF9RabysvJ5LNbShHLs6hwOZGkxI4/ggNmgNuYCRfzaweoQQxXc
ZpxW87JpQhUh696NNi1CSG7PY5hbOMZgr1xvsGB2MkGJWZac6c0MrN+voKNBNNum
EeNAkSiuTCAK4SjQ2u+F8e5muXMSpzRL3eQ9m2kNcgGSuMPAL7XRuuq61u9kEs30
PRpfFJDbvN8GVqHqNEelD9YJdgBuEEBHI5zoUI5l74TDdLONqC5U8fAuFWd9M8OF
f8EIcMCE3vsw8MqJBiu3e455MlErz1uUk9u+Tec2/P9SpfM9ZNsZko9f9U5WCB2a
6Mjx4j+yISaJdccMeiKDo2x21hA5Zzacvt5Grg2yYMBWWwT4lLcw/NM02HkLe9fs
fPwNOu28EYxWWGlOMg44EGLoAEVYYXEfEaaR5q8kWjC2rICbUrm0fd5E8kcgwicE
5/a+Hvzxw2eee143/6QQJManwRl5I3wBpgE0+DiTbWdzo/Vy4MrEP/vhDaiIeOtO
YJcMYMmhoKXIoDYQ2g2F9Q4THfQuZChsyfcssQfWmhh5K8Y1snZlFv6sHUVNgWTE
kuogBDt4doQ2SD0blMF1CQHyJNBZkMThC09cYu4RDpp94C6ZK6eNEfidbyjvnB6q
0IJTkHElJa4uFsyuAZ8WOyXuk4NoVRgxXqidEGzlA3QM4wOfBCwfhOVwjTgMnjKC
09JSk4DfUSiFEBqupVo7NS4o19LPIUKS0h+1mBFJ8wP4ujTCLLAoDMRERVB38Rua
jPlNkCQRlSF49gJnSDDkCJCe7ladtDEnyTPuyicqYVCORYvsdkOenltIRCfMAuls
MxdRo/20vWJp0g5y/3KmvdbbDTkHT07HkEjqk6qgR8bPoEVfPUIYyBcJJMxmK7t/
7MZvqCD2K5qzE7jIkQkPFRo0juf62NRHsfmt+TTomUARb0uPnc9jFLKil7q2U9P/
81TOBnvFyDL+Bo/ICbBV0vi2o9K3VOORa5kmCPCW9YJwBmP5DkC2y4M2TBVUkf/3
vl2nOxiC2/ZXQCUBCP6lBtpLOXQgsBX78vTFdZmlu2mBnlp4IZk60B1IUbGKUegz
MEc5IT12VKSq79yxaQNJ7Y37rzhchJlOJO+5C5ypI89eNTCdUBnBHUConM49GCZl
XM8dMj/wtG3rjixlwQmhE7T91H1S0mU0tH1oYl/SBdGE/K1wDS1N/XdmCd3lm6f/
B1SoHQ9YMdSO+Yo94lNAaymxMIQVctpCAa2bRh7r+VHb3oyGrubBWnkc6HGpEzSd
LhRASy0Res0N7IrBoYP58TnsZMg8kJs5wNTfot/hMbXglSThiLexHJCwsnDBLiin
uahVfo2Clbm1iObICdLx0LzBCvXlZi5wcO3+UQnt1TXyN+UBdi+nYQX4qibruZ+f
ZyQuqZcmvsjfoTKp/ekPiNFFOS2saoiDOVjOdKpQySTZo1KdV+SN3Mb70oSUnz26
JHtn282VNQ3KtwsFqvrDZvgDuNhPRsS5hxt2c1Phm4aTZg1eQWn156LiTzNKXGPO
os4dYnRiKnJ+TpkFKdLomReCRGIw8ktBqo8JK9X0MkWYX66kTuidSkLPd2QxttiY
MBeLJ6Zglb4A5nDSqxEQAZpAAMqUa5FCZB2Bg39IhaMrYg1J/7GnzHqO42R1ypn1
H8nMZXZA3PUJ+LO65m+wsbz1NA88ZVIBI88RsbROKlI761vtOnIaMxYYgveqsQip
WWUqjHKQHedO6MQaWillhiRtd7AAGF4b7dJIP9xxx4WIgk6+QDFwuNHiN2GVPEv7
mg2FBCdAKw7Ej3rY00AZ9TRvILx0B/rj6DajcTiEeCEtO5dau4Mqvihv/WwIgSQV
r66ZqCtRw+GW/8f5UVv3boJxQZYaYMw3Z+f1dZvsaNhmKlGET5rRvwltiy/lrqtc
7F1AI5EsVGx7RGad1cf4yE6HOYo+kGKMujhhohQ9JgxqBsvehfQB7SWdHmct2w8J
3/RBm+7Lx2ViKDO+SlYzNRvHtTzun7RYHeLDb8J2I7ExkH6Yym9jMC7klkkJ9xgl
QRLXrpIOeZI1o74FkpCdCB3/RC3ox4HGpk8fw6VQfPO9Pu1Vuc4ewyWdwbaA9v+q
4d8yF7ES/ya3WV7fJ9AbLiC/9jArY94QfbhaCiYNWwxqRFiPnni8vNm9jIcjslPf
RU1vMF0tebNEzqJ1YibVNla+q/qZZ2lTcOr2nBbIW2eqveURjn5AvUjfNurPLJOq
7U5kDzTyd1ttdTO2MHr21SBQcBcdXsJRuDPHEObPjBVWJXpHsd0bALKYwNbq5Gpl
VDiLeENQbf31hCCYrbovpeFwzVZtiAyK7CSo8wXS4+DTWPemrAGbCGl/HZ7zY5DR
j+p7AAgNhYWr4A1FEgVHo+aRVCz59oXEw5Ug7xsC96q5uokjSWBc5wI3tw4KSBLx
e9OYi5tLDkkg+gSbF14isc4E0RMHgrvmi/KNZwVkT83zVu6tJT5KTvh7CF38Z7t8
U5Pp0hWZrv7MywKjSJNksTY1wwQ2fskIYOvfKUbzUgVti9LGhcRKyWmnL0vrOEsr
XdhmbfnhghX0wyiPcBgKCkJbPFM4SYRrTku68EGxe8ulUPKPeZICyhU9EbLY2Cfd
TwYhBzVmlCZFAaVaKyE2LBHDJ3Ypg9u3V3zT+czu5APF57phAdKOJGqd7loYXrw6
64PaMB0aX/ZaObiYWgxdpNfYQJnhA3I8ScYUDYkL4DYKd9sLbkZ+nKWAogD8hHNt
2GZGTCVGoSrbNOxF8n8tlNT5rmpKMOixRmTZ9nbVGKdhtm4taGZJKp2/bhpAWZuB
F9vKYM80burqDF89L04uHQZafa39TVEzPNZQjtfqU7/zCLfv+4uPq5AsCHtUANmO
0w4uT/nhVQIyBlXvM/fNbTAesMtRsnd5Lw4vdsi0nQM9yWKO3GaAg+F8RA49vBNd
HGge7wFS2rJ6//S32na46QgIJtIc2AvoSAB1K2Eo1gLZqDm29ZOvMRelVkOShp3q
QcY3J/tLacY/Uj90pVyqR40RZ7R/CNtl7vrzUuRtbXKTB+aE+QkF47Xor4kgP8JI
vZ7bvjF2oE3SyOxTjLO+7Aa7kJsxad44QbJFRc4DZ/7aKozMJq1ZTgzRmqVPFW4W
l8O08U+lh5EeAS6+IW/FelQ6Hy4D+fqkDGPKA3GGJP8SxvISDgD2TaM65hrpVUhc
aDsWEH2ZU77A1TAMHpGohYVxxBtEVzipalVdVYdzbFVJUo6n5XMmGqcdDQArl70A
2VzKmxFkjLfookmVock1SPyCzK+39g9SA+ZuFjWiFniF0mRKmbA5KJCLzP4Oo4sM
LSdfgn/PblzTNNjIoPsH/WuiGkX0sv/67kLaku7WrzC54yee14q+EiY3YW7V97zx
M2Aahg+dqEkIZqhDRnpD3c+uN1ZZnBoPKforurlLsFMK6jjutvc7jkswN0NHo3jN
s4OIZv447PrlqLJOCviMfPnd//Slxn/GvZkHrCP4DCgICujakGVPGGMgrGOAPX3F
03QOJUPg2DssZjEnOKaqXXbPi/waMgijUfOHJGMOSk+JxhdVPs65QIzl5TZWoHgx
HE3ETo51neSWR8JqqmihMN39OwEi1fz++RHcR6YiDnZicdt8uahAzTAe0DJu5W4H
pCGlwiO/U0fW817IWe2rqR8SgKqrQJNLCkTrXkSzdL9Q9I6tXUMkkkKRuZNoLxU+
YpBTPwRywoIzLEQWqwSTYxGHMPig/HFyKKnANZ93JyE9yqK7FcDH/DTgffvkC2nx
WaXvwpFgDHJhWUiQTqAJ8oiH2jZBgwADNF5PGiX+v6uvtGFxobHuPc1QU+2FCAGc
W4hiCa/r3/TckvfMxb1PAO4a6YTgE8np6VtrXRChiLwP5uTgweo1qnWtxYPM/c5D
MXVWRhoCbQO7HzCs3l3trMpjpmlHkQBuP5eYOSVDONPZwKJRubvQaX6xVQ3xBcXg
k+EvT99eTBQ4+Mci/uTz2gVLf/AAkyu9Hxw4DKIPzO6mfaRb0DU4LrXOjRi5e37U
t8ufUEW7Vs3bROm+ke3inpWyykBOCsNyy/S6Pu/y8IZ5YrEMgNVfFVS4jd+AjGiS
13ONr2MwkEpeFC4MdEWWodOfyrWuWIuU0dijuwcZYI48atGqtq+YpZxsVWmS39NO
9MJsHNPry7KMJWjULd0FKJnK5j9cO9QIyJQkisy0SPyeM1f9G1fVaZIakq0gIToi
lQslWcn47wYn36H/SheGTR6qzY3TYzrtPuGpynchdMrXGhS4Aijmn8U/AS1o8C/u
xbGX/BI1FKKLAeQZqW6rRw4Kv1MZ0dGsEQiyHP8I1/jdfU+ATJNjI4DcijQ4/oWB
2x8ism046wJNaXwwkxBLVzOM30Uz3HYYljDN3Mt+/tjtyWTmb09Y2a24Ebvpbt5b
09p+rH8ETvZh5fu71Mla7w/5gf1B3GOO7kc5/TzKDzOaIeP70/YhhGLIh4z2C7cP
sDCzBnfaTV6fGqUMF2OWVMEDUxsdiv+pkOUmq73UzxOk6/PKjvwE/AKySHDZbqhP
lcZJs7zN2672wVJEz7yGdLOcPMOo+YQgOMeJ1egWl2oVjGU6Nc1wReqUOBuPstMF
A02saBtcQREmWc87MErLbOj67z+bCeZTnzIlkynBpdOZNyrYnLbGD1hyrLQFUQas
oOK4WBn534LqgJQB2DEJ2VJRrL5+EUiEgeWomqowDh7vRIvnx57OXGz9SQ+sfXxW
HnS9yEJYGomP7AV3G1GdHtuD2WYWvNpMv58Phe2qVvyJfILKKONlUklz8Kb0KwNh
jvKEFMiYywKOU9RtOY2K/kB3BLNourBekXkdCqBnHauYLOpPVjiqFn81ui3Z/pfg
ThM6GOhYevmhOt/WAGvY3YVhVhIyu5Aw2YaG1m7/tzYEifjWZ8j7jH0kHSfDyoxR
wBC0r7nKZFGibR+HzX3uJ3LFC9DA8G4FJ21YcCW8QwJ+BQoqNIAjyiTw26ucc9vW
s30oQt49wYJDU4juWFB4whpwRHsqlymeNWouInyeF3LusZr+Xrv2o0DsC+hI2DcW
DVVontDPtZlmBxuN1ea52h1CvkYgMP8JT+kZjrumZmAUjvD0cNgrfl4sXHse9AL3
znjcPSFu0yokTB048JK5yixLzcKSb3iOpyOOLdKvAIBzAhF4/yfLMNJidBokNGCP
s318CkYj1S74euuIT+RoarRWqP/O9TdfVHuSkluGUENFdLxmPraUErNAOEo3pwxd
ybbrAYBf6qPyVaUQ3SnKqT0McN4rgC3mayI1TeuNuv7dArm5M/YqJ1KRWblTTG7p
1+NCggjHLBI65gUbeD1HhLxdP/5CRGE1TuNDnO+u0XJ9b0ViS3yoKeZGYXDBOVFH
XcH03VmguZmcsie7erSwVypCu4aTRPplRfQTsxv9IKGTbHi6kcV5zhWRaEbeKQ2J
dKhDlIioMjtyTyQQ72q1CI8MdJ5h4HlrRbOOOVJ05/ljZA6qJdmDv0QOJxbIKn7w
QPDWIv2/IfBcTgA1rPL2SoEiveFFGxYX7JvelnurmsmujBnoFzKiztBryyYM2Lnh
e4dwRf5E2WXhzkd/O7Ige3w8hurBvdSVod3QQkiVZ+fuEY5+PWX3IFpUjLKHd9JF
z/JRpn7oweWl+n+i5szfsC+1/5VF/EOfkWUgVNkQ8zUSnVY8x99tp0c+0QleSegZ
6xP+DRxgHxe8CrisFxfbK6PwwHrUcRvXcl0ghpimgYw9LU4tFUG1tBrzD9bWrOzT
PcSZOeKvROz4ImsNeYjViYIw0Iugm3BKkaJ0ngu/Bt+T+dS3LafJSNMGmi7F/irr
r7o59yzshvLZ/K05x7ddTfwspgNKtaLCXHUfSm399Xvph1KHM1vQwtVR2DZ/f4b1
+r7ee3OzfPI2QqdmpA3PVK8PDRwrItk5ExZ1lMjRHC1hT1mSW7zwYwUmOH+MZWvX
cJJegxTNn/g6VpAaJR+W8rtjIfLc9eHybItejLGU0qpnSfpuofVIrbdc0amrh7pq
n/HFkMWGzG459BYi8vj4fB1uDe2XM8sD+ExHSaJKvdcdlkealO9AuLu3lbsvMqdb
/riiAs8+VMidStL1AQunzXvhwhqrA3Mg6PN5JCAVEQDH2ciQ0Bop1wL+HOXEvpV/
kMFupwkFzMTVKES/ivsfVFc6XeyLTybebeNRNLyUohj2LV3jIPjFYtd5g0isx4O8
IjK89NzdN8zx8njQK//ZIDDpbotR6fQaOrEpI0dMVm5TIYB+Pt4pEi/D4d53x2RH
dyhk9mu5h6j5zXSDDaGTdY+W4kO4v/AKv0rB5Wgu4TOIn33PSfhqGHI5pv1k5++7
QaSI+NWRO6+cdDXIxAUhYmGkKInar9y43piLRAEYwtB1eiyO7C21iUIQqwBfJZVj
uKysm0KSrnQEbmrBgunhxZk+E0NKf1nZlBZ1lwgutnftRTGD4fzUV1XZ7l2CVk8J
VVPWQ48FKzJHi4PqV11jY4AJV1iEAYzUnGQOMYmJ1TsIJVYx8jmVObW3O97cZ1V2
PnhgQ/D4mbySG+fsCLoQcAzcl8QZzsgPoTiyZqg7BihEDLBdkdEbl4trlk71MOTy
CJMciqi9OgmY5RKaWXaSeg/szdC2VkcHzpC0HU7jMIofFX8GppXoeX1weo7V80cb
zVVn8OMaaUcjOJJMT7Q2H90lL1nJhiPTXUfKo6JnQFhoU5hELVwU+chfGDeUdPNY
QpEA1t1RUrxwKsSkKoATHhngLrJMp42chz2PT95X5E3w6AOaoSulfvAPd2+qMhZd
J0TqEROus6x+EMYviKcJ3AdPbx3L74LhOKpvLCTqSP/+1SdKh/G0FTqVHnKw4tRu
B40mSxDMwJzScq9WU/8YLL7yFFm80aUKNK8/cO49ZQBGX3jTBHq/asA0PfmoNgSg
5vY7G1ppJRwri7dOw3h7D12zfUjNK/cB2RAHq0QehIBOm2CAMj2G3K65nsoRmdjD
KvHSLkQA0z2awKbIXM4i7FGSHyeqZhL6mKTsd7j1j1rn7qXPSgRyhGX9UC/4dupw
xVmw5knXmcjaYKuFrxfiPcPnGFH5oh9YqqCkbW7EYlsF8ird+JiAuWMMBgF+EUXR
ZYehCdP+JrTKwJBawY0SDj0CDW/x4QBBSOq/TlPt7R4wTqRIq3pkpJKvAZc8bDac
lfTqPMUSBh8ZIZKrl0gkJnFqJQ5Di/azbAph5c9wCNazUf9ezbphuY22UohHHNPv
VNUAuyFEYfpfTb4JotzvfatX6Rp70VzAb/qk5MkwVdRGstpouRxSukoMuNGlhWo0
rvaIPTBHzLFPOaS/7VxNuUKO45aYOpJ26wzcULFo2aW+ukO6hzCKh7qTq4n+UbEZ
mWTftHEferyJj+mKT4peG/gAtMWVSAc939CBqbUu88bQtMhpZ7S+IRn/Nal7/Tge
lzKBOZrbpYT/f+lFcVwEwURLuezB7zs9qyYUKrYk6QOatD4Y4W0dFSVooCcCbvem
FOmC+Wnv6cAiODUKm6gn4Bi6iWUkkcQHiXbd6UMC5x7xUsBJHuHfDO88gMlqn+fZ
xvGqgvpKuODmGgwi9gV1SdbaqgpuXtaTwkC+tlUENSnPuCjQdcIstm4Up9EBQhXX
l0F8BOxw//ERQrkokE5UPSRGppn9Od0VTNUV1CRZYPz6OKlDjGa+darupIBX/1vu
4T+EEZ/VVk4JqYFjSYHZBsIhvhz1I2YS/+BD+4UNHO355+Yz4W9chzxctG5kCAS2
TFw/Qry+4Yjk6+Il4T642T4d9NsT1XcJrnxh/GTwdpKZZzloJu93ztJ1R4sTAbb9
wOsQCJT3NNQFkBuA8L6DGFL9BvDhqPMNcqKSSkXCP9Q8UT26DmtODpiY6jjaHeAB
qa70DIQR/tgSJMNuhxRie0+KeFhrvC8UQSoeipSGcGQhmXNTDMx7vbEeYDLwYb16
qQf/yDM9XqgN2m2LvOE1VOtOYRymKmXJPcDeVjryepoVGMzf9yOVDTBs2ZUbwrem
R3tI42GZ/gFrDXoSZLXLSceyjlwqCDoUw1Zbe+bUovIy52O6pIdaYP0F15Guzv/v
t+Ni2zJThb7y68KUkUV+ywofXrsbvlw89kUs148K0wCXSyUCneV9Pn9k+LZ1vXzk
3QjbN16H5YrelsNnHVTNIK+zSBkjHQVmege2TmPXd3LrHPJcVHd0X5XeJcc5WeWQ
ynAIb/A4P5fSRQNjvt0IEAnkPwDN52N5S9Vqkn7tyEnHavzcZ1n8WXBrXnN88lF4
qlCc6VFDOT8h9aBxGbm9WGyTKej/NjcUOMkqH1F/L4m6zUtvyOQGYZASKPo7tlCd
PZAsRCg77C1eGoEjAd2socbpwwCLH60wPNAZq/K9Z+cml9WfXIz5mAnDoaBX4gTA
ue70rXfwY8FGVDE/HNSQBWPAkgyNX2M432EnIj3UyWot3pmpdjz9NU8VIE1hkesa
NXD3pc9lpAoWyZODWC2lyT6v7Id7pVjbp2YloqHkztaXR5YhwnuUM3WJwgj+Jpyq
hL1CXUD5fZNsnH+Bz7h/d7DEAuuQFa1n3K7XR5Br1sq5FGR6onaHVbAq7XwEOOU0
vbViWy2dvGFAzJ91enMjBLo0bk1mLA95GKGnioSqECNgZLdr34qmOoLXEbL5r9Pl
PwjD8Tpocwrl5pnlX5E1ZerMEFUvPRsSizYuujjZOXJoxOJfyTotSbqwaytc2Jio
DQtYGNRhMmIcdhls1LVhoAKIE5Fr942qhIMmzvoKcTO0s87eAIZvVtCwdLKMrCAj
/Xd4bm1fIz0OI6uCmc0QkZvgCHgd7wfT8Wu8lGhJjdTrS/rF1Oe1jjGN3tPP8TVf
beASxr2EC1YhQLFV2Lq/SoifS31I2L89uteYgKci3KC5SmU8seLPfgWiU9YEvi5e
69Pa7UN9+tpOIVt56+KQPPU2TaEH/NBwi2cMOkVNp1/iu1mWRfZmbKgQzOIngYzW
DI8Nto3fG8512KccPnJYG9iNR+UPnGt/dvlIjsZzXu0GLOAXZyKlZlv6PI4VanXL
RMVGjRc5y31w3KAnQ8Cd0ch0ilpY15IFoXseMb31KsEJ+pMr4BfRQKmIgY09O8TE
sUMZySGzCwZsOqZL+YhF9uIH4bVGzZb3L3q3zXItcETl0ijI6Cl3FkLL5SdTWdi8
rHukFwutJVzRMjBX7+iyMTkvav5L2aiYyhycwrEXZrvYCGRlVjgndotqrGStIFOP
YYw1qfgKRjXimHYYqXV5AsQ42SJsc6xGE6lwY4KLuB9sY9fF1FmtLvtGFIRKEJFK
LKNnAyrKMG46+Buf0gFsZ8AAuJcySqy/sczPTMeVEQjSeGWHMSUi9NoV+MM1q50t
TxgfJE6n3cdKJheZkUW3IIpkyOPnVo+3pch4IwuHxBXypRtA1bcP//GZhOpwGir7
yKhD2F+7u7usn9EyO4Bo/acI3eeAEmwAZNeYvRhtRjnW4IRysyAs5NG6XTOopaDJ
SUoVutNLvU5QA8c84Pc4sSrLjv7Fc84dmxEIeVS7X7AWw3fUn2D9sCJTY+FC1h2f
4veZ1bCh4b+blCgwtkUqphjLfu24kRFMpi9JJIEV833vVHTjnhO+P3YGU88I8ZcG
zOmtcWyc1+Yr1SuyHw6Ui3F6vxKZKl+7tgueASnPXGqXRBAwlT4gKWwwdI13P+of
DZOt0B2sluNnsMZzBuqrjxBsumKhBqHPZKhdo3vH1R+jqQN4AqOpkTbSKqdPES0k
U8GHkqU8tqc9MUA3uUhmGdP2LsDc33sQtvQJnXB15mKtLf5Bx3VR5TjN0A0I2yR9
3bm6dBI0VTwdTKuGWTMV6trzSBq1L0f3uvGLisxX2FfRlaiF8OP2EWCg+mes9+sn
knKtr5KoulptVNigmruhBhnONCmwMufzsv6ueLf+ecJ1RyDc0CT4jwF0lxNJ/+1p
xfZO2O51sMvHtWaNvEMR2Z8ZQ0ygz1aGe0roSayQO8s+NEU+0yVpgShV+zoi1euH
rKPDxTH0Dkjud1NFL47R2IT9vV/qFzc07xbvHHoLyv9ZcIkRz3R66CkZNEfEq7eF
a0RAAfdPygOFlPl4u16kg/pdBGJEudbIV/gZ/Rk1Xi4d+DDg4rnFA8pnm+EZn29S
mXsZN0AS3pDXFVaVLtFojAFEFQo9Vne8o53CCgQY+X/6Tmwx4lA3rSqkPtk8pK66
ZlQ3Y+Kn2rVq1HyuTXTdIR5Tvbk0e7NKo8fGNtV92YamJXk5ojMW5WeXku6+3WEf
9MgBDoKuighoAl7AbGhMPdhPn1TQhukSKl6MeoiCWRwneIw6s+5OAUH1midjkmYE
8UJXF8/av5yzzGilm8WQWirVPWPFQqBLnINRzJsWvUobGosiUzafbDHPGCiWBqDZ
bTMCH5pwhHP/r0N+i/REBvFsvVdlCAIedgv9YaOVi4Ulu86WTGUVXd4Kvs2xrCGA
2FfjLKOulFCIRLuktuxwaeclGE8vhGfvvOQT/pw6eT/r9E7rtmEwitYi0g8YA3pR
/p7hOCo3nzJJbrHBPy0RCqXZYAblnIxQtO4AT2tmudWmxxYx6TsIwyq7oH2nhuPK
DieXUG89itZIdxH/4Wz8s9RgQhFnqrTcRYTEmgczsIiTHR1LRFWaF/wv1C0PSCkn
ttW0vlzVaETwlvbkPWhug0m8d/6iELFCmeswvi6gRLeHe4ksVa/6nAAXBhekaxgT
QdwIUw+HPhwJscsLF2uiwQOgEGQ9s7MBE9HflbGd6FGT46Jm7cyIf4fLl+0U6RMr
L6wCiJWjoc61oSMoRD7V+9SPq2Oi3HDC6MKQTXwppEAF1SX2f6nrlcPL6Go0yBFX
VH+9hz0vAeh54HcCvVQFAHxXz+OqupS65wevKvHcNBvWZ8b1rQv+zgKQDjbDJK+W
kONwGyclG+TpZscMQ3K6CotVkWy6FEngRBWcGCd6lNb1JKtIQ502Wf2bSkxGSJPX
LFCbWOFbu+/ja66Ag3mtQJHKconorHtTxoOIhcCkpWmYvOZ+bR3rN+9TABVz9Hjz
P01xQ2HlwlJHw/GcW3n1pnDq6ezQHw0E2Q+7GAYFkdwOYmtNIrYpYAhnAKdIt0Dd
CJ2v/ZiSK9cV8F4oerEuYnHVSUUfmKG7EITi6rbRNNXOTowR/0sJTAE5zZWzyPuH
Hm19wx1mQTuPbXa6dlirJA2HfbRvDz1ezXG7Gvz5+8tiX6bYnP99Z2yQBUm9pVYr
cTxlTg4Lw65YstuJpxRcoflc02rWE77+e9e6eLdNf1kA7cQjyoLzn8KAUzqU2ifp
mU4bqcWdp75wgc14CL/bZ7RRhxbYGcTOvk/pGmA24shWxsR/OeWeYhDxuf3iEzxk
h+NRHWHWotHCnRekAoW6rsK9TN5cL3uDLeEZxzDbSdems1c2sAAv2RMXlxcHHmdP
cbqE3X/TM5QXG+NaTtOyW3nm+lJcldimDRN0aMn3Sq8PAa8CZ9BDArPc1JJOH/UG
CboVn5q6gVOsq+86vpa1C6aucTpDrpc8H0TRtTmG/avfJ8XR0kPvVrDG5G91w5nM
T81fo1yDvFC25LXDaHUjCdFMNrPgaoYpfXVIOwPyuxbtktKD2Zd3ociiclQWW2iN
1p9bP3OwiHhFKMUpmBJdbTWs4CgeDIgrnjcOhcH/vOfT/iJ2fVs+HWQLw4WOSI9j
JsD8+prVh8hikgfwb9UJZ0DeGkYfq8QtJH4KjuHLXS/s5CR/D5eJZ6+DqvDMWCNS
rJDysOdLjgsilZn2QhHRmJNjuEcdZ3p3Ybt4eH1tBzpj96Wko5nPyziFQ2afzQ+X
rgVMOgp/5e7x2UFMX5J7Di3himGHZiXVqvE5qxTPlWRsNWG4TOOHYQgdj0lIhUp8
bWancwTq3XCP+fyrCNsOb2X975X8Ci1LeqRr2K4K3GTfqiC5eon03JDC27Jtvmdh
lvmEHS2IbRIOtfkXisQiJ0IkkEo/I7ZyxCCR340JhUBfgaFdULEDgVA0d7PtS4Yt
dxh7vTF3s3pK0HBn8oL4U9iVVldjpMYuofdfTlvN51GiHB832VkKkzhThJ4KG4U5
2q03/XKawEaps3uPVf9C/vnB+1H2gbR6xWKKHF+c09d+VhtN0B75LtohzO8Uz12/
0mrQ9BK0q3fIXhuGrMFSZSLcdOjg78jFuQpNuVbKPob4cRgig4UWSzC7cWQlLG1w
9Mz+GxlCXuKskty71mDVT9u5fpTBWk2y3QrRmk8cXzn1PpjW0akDgRitubQ5T9OO
x/nSztbY+8ERtpoMrP3mH4j18OTiC1iTtn4j/tGsZddG9Q3X1QDgYN/BftvQkgkk
YTcSyhlQaPHmhfGdjY7kPMdaTZkfh9RmMx1Z0l929ljgT5O+JlbI9HMu82s/LQ63
RJgYSzg8VgiVIOPhC/rW9Lle1YdFvz/wb14OSS3r6AyLGFXfdbukjrIRHcZIi759
Vz1wC9Mhzmxhjfozsw6/aX3EAz9a7S+Qu1+8zbmRldU8na2e0YQBBkldxlImX9wc
tSSs8eScWqZn0ra/KI0VNKg7HaEAaitcIw9gxDgWMayYAjWgI+7Gr/czrm3eu6IW
OtyLqEJS9ppEfH2TEfs4RecCxYwJMDUuErQwZHuVOllqnisYZA+5bodzCqUqOWNf
2F69rqORteDEnn1Zg34aos5D2+RgURaxCgkJU7nPbSEQOTUa6+svh2YddvoXHJjw
/otqG/DOL1qWWHHGZaYuO0wnP3ZFpqYuh8B353Doj9+KtlktG6ddzxt/9ynv/GSl
wEJheeXU0IV1H+xk8sRoy+8LBAnZcD7o38uJMwEZ7OtktXfx9z5TzdYZv0uzw1n0
pBuFpYFulRSItkiwfK5/YwCy5qwlUx1gMNviICEmGJjF8uQJ7NQdZC+u8Jeeap8Y
s3vRyDAVdEqS/CdLXKwdrT/ciTD2os30Sw+mno9F0O1GIfJQsQuBq9bimRGvv295
EBeNEZ1PMQ9D0PHLDhuGS9O8eKLQMt0Rg55IaaBNGPNx31Ct28A6CpGLsAW/Xkdg
TWNWURI7442Mmp+ZPh4cB92Mu/YykT5Voq1IYZl35Z9FPQHHDHF7ax3WHyfw+X76
mKi3oaHQpV8soYLxZciYKopDTP4FyMv9TXSqm/cc7OIgC9I9YfgVJxDQk2OMJIFB
YbqN1ZO+uhEuAMz76o6raJggaasLn/QakykAnTeE9Q7eALN7MIB6b9p7pv/qCp5H
E1QYLDVH6qWHLZvn2JMVtWfLSbdMrn5/0USqPcnrQg9ct03hh/I3H2EPwWalZ5Yv
xd2miiXudu8CxcKyJZz7HZuwkRIiwDHqh8I6NueiOf7VoK859FYxWFlsE7t54t4X
JDbs96rbZMG+N1/X0rOCXkuHKQDxqfmp67Gi9z/na+C6OppQv9t2Ewjm5sQAvg/k
oZBwSuVJC38kpgKLsQ/7DoWJVEvEACxoC+XrG0TzxuzY2+AXiZTZLz2w7M+0WSRs
6goBKom3uZ8tjTukzc9xQCFEt91yif9LQFbHiCHgVuJ1mrQai51gpj86CrWviScd
J4KPIV93BD0bep1p/Yyzm42aCX1ae4tI28LT11S5M2oPcmMJzxGhXUYUyGBt+1Gd
L/GnXiNDK0ODW0FlNTkoEdevU5e4asgBHh9+UWXlt+/2U+AdVFvLso168fvxgP9P
HPF2gMwxXQkNSWt4Y5DxfNcHx+zBV4kRhLTIAhhObnWgo59euAW5wXg5KoLFsryz
5uCmdz980zsz8nLziF2iBpWn+OPuKULbmbEoiZBx0yDzgW4vM6GZV3FQfxnaS1KF
JfiThTbY9TQTZp8QApTQdH8doGVaW9pzptiTI4mgraJgR4LgWlXACTlSDAUfeDS2
l5wlk3CXwhaDUnaDi6PfoarS596NCXmTHiAYggSKJq2dIc9RXlmxD1bwQOkFDaoj
jZfwxf1QAk3ue9AJG3GGdGXCW8EdKaLekIczz654yTrhHktwOFVVt1dQx1Ji19u/
JZtINwJ8ZpfLfHqYmKbgVFK18gCSd8OUgW2qE4FueWH1o6tS7pghdzKXQx/1r+1e
/Xhup2nqJlHjWnpWZW442tKORs4DZ4gGExD7MEw5fYMizBimODVW+7gJtGHj2pZ2
Vr+Uky5AG0y1riBjbV6p++4N6XLmgis3m6+0sn380KCbVPX6gxsxBJsAXxWoHcKt
1ReL+VlKq65Z9uLWP8NcNq/jVcFuABZoLFnHp5UgEBJokV/3Lu4Xek8bzhJVEB5L
DPVncJNq8q+OBX0oWFHmMkvPBfcB452/Chzyf+i2RQ6UcInupZKR9rMEIwGw1Z1P
Q3lrjBnQc+smunKINjZN0j7sv7uyFTLxz11V/eanLG2aKIFnQo36QVbjcXYodRad
0KXAngINzYFpQqyhxqVtlqr6iqr+Jq9s7DtEQLsEhm/kZk/zLN0E3VZVkMkIIMdB
plVD2M8RSpGlqfmIdUirWPJjhPRzKNY8d02hgyrJRHwAA4SB0izUNpVFfmkMbZM5
MTj9JURR/DLEmT/rSuRNGEn5WYhOpMqeyaSfXzilBYyoDA0+8QdZXsH4VuTqz7vr
lYoie60Y7zy88EUfOe1XJKte9AC467YCxkueYfmgXtcVy6iNiB7FHqlJL9P6V2u0
tzxYH3z7O4Yt3xoQJxO4dXK7AhdcwDd6t7D7+oKeeIqOJHO/UJe1KQsXmJ8LS6Ob
PQEmt0za1vEzUlKeBNr1S1y+8s1gvHBl57qN+ZrMUfN5m9IyYfaPWEf6HOZy1QMb
qT8Yu+3YbHx8POZf6IJlx1DpfsVj64cNIJkefTk+mj3Ec/n5ShfxMPYT5l03+qCv
PxvM2vLR+VS8tLdGJwTk+tH9UA1jmtaHwCIz7CaHIM/tVUepM/+3XKxsnF/56Dse
ISjowtL8546hUdv7b3j0fhusS3OgjoC0ArNcCei+ju51Wkixj60/1YLn7br2a9nA
arwe71ATCR/B4+3MdDh65bcdRO8ttjAbPserjKJ0qH2kSabICol7/TGtp91U5AM3
XhO3aiDfx4vqKi5IQU0wcqWWlm49Bwsbu285nH6hWWOTsYEDEfYDsiE7EnNv6q5U
xh5Mnxi1+hiERQQ814C6Bsp4n7fPj5qNGwy3NfFmXQ645oko31p7GQ5rJqLQtLsc
iexDC1LBR5bwJXcsrRBoaVzLHiAVbHiFvgDIW0+eOBZ22ztfoVIK1ZmaxCRsT2cJ
zr+Z48A8kdGq9YjG89m9gY7uHleZOc4sbSbjR2D5Ed5sbJ9OOEeyszxlySiU15Ey
xMe94JFyaeK6DlJY0eaj9eeYl9x2UKb7X6+hPd2UVKupCdB9LQtoOnNanFFjNqtN
aiBgyVQ/5VSeZqvtBjvURANvdJjaOvVtgDVxTofICpyzmwjEw+HVcliZyCtLZI94
xpxS/nJYZxSZeMdcy4HObRsyxQEFiuoX9tCUXXZJR+kFarCvBkvVKYJnZcBg5Vos
rHYJnDmwWh7kdrxvsw/sDcIqbaJQRRtDbs+WSXfDjvunsdrOIQ3X/hHyiv8qAdyD
BqFKWa1Yop64sd+Li9wH+V20p2lXaQZgtNL49PAeAWEvl0aH6ABpy5zVzJX1uC7c
wNRW8ZJAiDfVkpL1L4aY/0QBtRT9oG7HQ8BBwTqyfdaFFAJkg9hpJZ7t9udi6Kik
pzVm6EgKGWqSbSg2wrVnahiFPBOdBfNC1Cju/+8VZvBv2dB2gd4HH/zClXpbshEA
1C1Ux45Mlc2ta+2u7vXajCxV3/R2/+lo0kCh6GXu998xz6T2Jb4KexKhYy9yixTx
DMY/u+YyAxysUUAFdXiz99YK/RI939klufjtRbRStinK7u5qAFtLk1hleJraXqSV
TTWKQIHUO2ecEXkcdYfsU19PD8ykKsiT5SjyWL8dXhocGDNx3FyjXVrpOucwpeCh
xJTbpwcNBjaLrfvFsmuCYOHpknV8MHFl+rvJNF7VUc3jzNXToYMmDIvFg3stBqCE
4EyunpNgvMzRP6Psu5+xZAe9RV2Wt7YV9EmEYuyEjlNkK5cQrUvZDo1cL3SCiTjD
ivdst4myzxxwWRQI2R9waY+GGo5aWt2yu32401pyYf3ZZHh9OCy3qoTIMVdEsm5v
ur7Z0v4ZlIpaQNv7wQwUBaFMurPObxLG3EZ2SGrkOXG4WN2R9mKiTzH3wsRJtJsd
2TzAOdzouJcy0bHaXDen3ikVSXW/sQmrAdhtAaLZJ0UFk7P2J1sTVfB5OWsN2uuH
fjzHE5bg0NFPpyXsM93nl3xHHJWCLFEA9PJUtj2RNFAy9yeYk3sGKgR/rBFk0P4G
uTwZGW/2CbJ4AzCnlWM9ewc3fN+R8JDLluJS3QkGsDTEHE9BczGd1yGa7QIviuDr
00LvqdxW1yRjpxOfKsFrxOwepGNYuWNsaUjtpBuu0P03EJ4MEFEhiCV7UT+krbdg
Ke6ql2PR6bwzBQ3lO0nYpbmfYK54pflBxDTUc+sJPQjLkdrLRwwtLON3juKbkvTr
EpmLTMWS+alO9crKWCykmv9opmRNM3L54S+aIIO4bsZeZcVw1LeQ/HRuiB9YxKRV
YSga5HkZMPYVvxV3SLA5onKBZK3fFeCytQGpP4x7nA8ktGnWCFAteYgyi7BbA0SH
FRUE6AuoG3HCf+ADARX688lJqH8HO0vdONXQXxuHhv85va3zNxiQff9hmWyKAM3+
3sYApxoSDX/DPGC7mGa0odwVkKb903V7RQT0YZc/DhdWZJxB5ZIlOuHENZzWW5M8
0uVhFBGjcvNu4ZG9oEvR7bYW/SYC5UDs+M+xl0spqPUm59vE9vHL4250RIl7f1xC
RNTkg9a4CAK8IS65Nor5r9ntlNF7t+AIZlDcttXStHxZSCDD57W+Cso5oAaVxJcH
FKuaInSOoLBmYZ+EqoG2HyNQdlTASkQLCmbXlyB0UM6khfvWnk4LIEgXwUcX7qJs
sgbjCXaR8E1BQAAzU9VjWpb3teDZ8wttYLmIMw6IRTCvdASkhM6wKJd3yFpR3REL
Bcdfb7BR/K7M3uXaw53kz3wARcT1a+n/jQDS+utLtRlLLj4daHTWzdEM3z828Di7
f8jjRwtgkLM1ius5TVpCLweXaeQ8LLheUrIE3ew8ccQYqoVRqC5ZOerjURy5FxfK
anUkiQaL6WHzu+Y/c4BZa4NrCgnnT6+HLNvx/nBxw3Krn68dNlStTYti7qNR2BJf
QsVPbQW4Ht1HNoKlpT6hSEinVNxy8cwJMA1ZgnmWDtpcaAqB+M93jpB8DfAxc5bm
vzPl22FH5/ZPqMJHRdeRRXov1IeJT44KKvcLNKNdMsnzU/1HFGH0ciN5zgcQKoWv
CryLbBdRglwsdnA95/ONHDXgWgyui35ho+AoIuJMU/sqPhG/nilYtS1yCre5y1Bu
DJaANoRi6NgvLsprw2i2ZH+hfW/Q3i0imCSHMcp47CSUL8kFG1WVHSuDdhymglZD
mb6O5MSkPXv9bM8z9OagQi86QP67gYvyGJ6cZ5iocHfWpYn+y3zWCCAo1DWthfOj
0d98TFVQByBubCyXPWSGv2MeXXZJpIFUjLvILK8fHMvtwuKH3TON2dKeU3GoI2VW
/9HOql7h9w4yhvIC0ilImK2hhBX08nk/snESi+tjjWvFn7b4djPET9yLmTmSMe2r
/e52thpb03xPDBOfNKmnt3P8ux4iu8gqbsc+Jn8xzvVukEKXGddqAgqVBlKfSTsM
4vCcPmZ3NwdiS63dhMvXh4uAX58nczjmxsS8EZE49b7fkOUvSYsZCq5FT88Elb8m
vabv3peD+4A7WFmZuqHy0391gnyBHy1RBuRFtYzf0IlGYbV3HCUuMPRV2Y3IO7Tl
WGHa0VgPJtLIpaVks0VM0vQ9s8vcrVC+mSoq80Dkr5uW0RdeSoQ6hPzgmIMd0r4g
zhSFD3pJp1i5mIt6G+Z4kRNWKIj3HFc4usKG3zuH+DGrHqi/nzTn+kzZQrmmgyVv
x3Yr0NYMEoilDQlVmb5U2uR/Fkhl4aApL951Crj1LFV946xwIi5Z0uAKgUQP19oX
LIcqP3NkBrl3h9huuNmvTI36FOibmP7MSHRi+wL5GXBIISQukMBH2WE3b7dzcQ64
pdkU29LEOkU7ARWxTDvOvxsX/uq6GYhQs8h7mHqWXywTDafjJdwwB7JXDrVLiCsC
AuwJ1K5Vpum5VB1ZBsucm16GEQaFU0jyb/P2HHutMvDtptIACWqr1V1f1em+o0TK
FSyvYmkFYQGaQvCINVlktw6ltOlOs+xc1BQT7d8ftaIji/mDkoIu/6lISR5/Fio4
zmTeSjyw0UYYKiXWQfcXXhjzvY06dE2wb2go6ntu9bcJhEOQBHFdOdTzUvUz+5KU
0OQtP7RX8yJ/TPfQlFw35/zicSmEIHrcc0R2OGS5LrLrJAyeV2H1udoQByuIFUff
fRsDjImXNFg6fFvA/BY5VgNuSLJRS+SQfC2+jmcCjhSP2aJu+g5t0EZqDeBe4LDZ
wbaEVpW/cLt3Z/sB77Q94fjKwHobnzgLkj3weeEdzonRzi05UcVN4ZZrpDdOoKcT
e03om8P09gxAGngHNlxX1/lBBq0iLXYc569W85Y8XZ/2zY1fmjDNuzP4ZtOQc/88
iPpxVesknKw5ycQMS/bXudyxfIyMQekIuwbrxiCfIUDuFOVVdtnHYJj0dhcV4Hw5
LtZQ72wtPAZvPMkyq+x7yzJDH4weH5Mr3CVk/eooPaiuy09YnA1apDWCbjGoUNqf
I/4Goor04ptUeZIYSLIxZcF5blZCgTRpJUGrug95+vAp/ZqF+mtthVrvdMTyaNEB
zHUBmWnvd6NPO/nI7SzNSf85jdoLuQiC+PsSCW0TA0MUkxsAjk2PEEVHwtRS7JuD
OkVqUDL6bAKTdXGVHLAoFk6RVj00kVxzbYl5emtT7lzeWw/S6o+eqU72776I+rrs
OTNECko9KoSOzm23JXHwZgS0+fJIn5zQh6Y8Oz0fB6ZgY4MkEBPM4An/AO+4a5+g
cYhRquK6Anuc4eQ8kOAi3gnuA04W1krRX9DjELEgroJTM8pH9Us3prZ5kCqwstM0
Rux6Jz4zKyY2BtAACfgIuJYcuqy23ut34Ya/8E16rEFiZwcK+FLoJ/3wYn0ck+Sd
YZv12K14uew3nv6QZpiHcM75xPFni0A0xyRdn7TjtBmTEVj6tBe4/LYYNu1tzcnp
yglbqO1ViUwxlRgjMkQLCmcwdCpYGDYvC4E7sH0F+RQgriU7I4m1RuDj223nIDgi
naf9ZhRyTub/le8GvL6De18v7p5yHv5ZtNoIJ/DT/JFR/1IBRYlTdaijbzqzHm5P
N1y3nL5+uRyVKxV4DpfALuDkigYE6WtUudL2kjs9ph0lPjXOkXxZt+fbEPwTWmae
3areQ7m7WUj8Vzki8IdZFoPLphBz7+jUWzs9V9gnwKTMizmijN2HvbiEs7914vzy
XRWYAI6qfBxUn+pHBWNYBrOZLyWBBCSurWXWmlWv33eqjYj9ebh1v2t1AttQ6K/y
jZCOkLtaX5gIyQOf5p/roc4f6N9UViQLuiMne28Bb0Pc1QgJNkCil0Y+BjJDPQzV
0RiecM465pGt7lvgbmbUBPFY0HY5nu/z1GvsKTyV2N2lLnYcXxON4Xz2d+/X1e51
F8tkQ91A/1inhPKlvWvAuMdrJ3obyElWJ0rpNuDB2aHhOrZi9MydE2BAEoRTj2Nn
pEASDNhsdIe4L2WpwYLIfukTEWikC6CI1NvTvnopJnZck8Qt76j5F06RDvi0yBPd
w/Qoq1Z0ONANW7U01NskZXtfDpEeYTldUzYznfR53bO8vTZ6etEMzVQd6/hht3/n
2z446f0pICpr/PmQjU5mwbfZO96CQTv6IpmnLA32aSZbBdzbT4cvoMS7PI9a1Tgy
eeFq5BXqS6EKPElIkwKX8+t0AhATSa90AifI4CxDem4GtCFbBwgPdfp/iTco9hdX
0q7FBsicjg68YVb3nX9jYstXsvLI15/4ii4kbblb7lIZ0EXqG2lFNAbJ+D5+qjdA
rZKwMYJxA4tfI2lQFB/nbCRcbzSwXGcQZ+7YhymETTYNTEbeUszc4jV3TcEa2Kju
aFdIQH+oXwrdBzYaCHe4mklOgy4jYmiqp7RJKVH/GYyzRqV8al65dGyB7UwYqVNn
0f7F6PfvBTnAhjthE0s412TEx0KNP0LeOao3mK3B8Ol4yC7PCAYskIgjoGfPIeHA
MR0AOJQdIIcaomOhapFoABIUoZhwzPV5AfkACfsaqevmRBDiKW0VlxSwFZDUkhQh
+nQTOVfX3sPNk6OK578LqsSdaZ6Of4PYDyQPlWzVa1gSoNL2MfwHw2Ar0eyNzl9O
mUODfg7dQBWhrH0gbk+dXuZxMNyMioDS39Wxq96mh6/2oakNXptOlYy0VE1Muj4R
qHCjgDyKGldYmhlRY8NhXScmfJrM/jenSbcL+r+FVkUbJUlGbQW7bqcfOoR3CCdn
fda3hOpOvFrHlUq6VoD/dEesvSMrcxp3rDv6uEwpo7e76fQ8QR4o0NMT4EVHyjji
jGB8dsSMzI8nWjoF5WGDTd+rE1ncLeitKbfk0K9Fkwpy7/SITHC4LM8l11+KAwAT
dlX/e/1R3Y+olhHrg1PAIPLRhdtqmlblR+Q4g9eESFr4S6BRut0lT4Xh4NyjdnKc
bkq/HZ9l2RJl9DiEblB+jhYQYyTwYLMuBDPdnT11oXSxxmK8VQ4XjMUIaRt0mIEv
JWttJFN5sTIBfVrCohvEHIs3J0w6wp6MtnDvS8LtEq2iRERSpUkJoIy9qIZoIhy4
RSJHgGXjn+vYawRKnR/FD7KJ9xHAjVOQWA0lxQH+IKFQ6jHJF689t1yaVYo7AJy8
2NlRBjDY63Xd29cUTn61zDj2sWCRAAKc0sxppydO5AfO8CkQFQ9zlgLEyqmNz4Gl
KoBMmlKkNHgxNUgp59uh+rtyr8f1RoKQhyntlb1o14czX4UYW0eJ5P12VN0AuWeF
c6m9WLtWtQ6TaQ3fkKxbXL3uwjg4ASNA2+0oVvgbMlcz5EZNWB6cqRo8anfXDxGP
8rlwrA/ENJI318ZX1voAMpqd3cTcv3RYCFISgFcgY/rykXZJ1MchYC12cSInRN4I
AxSQD/Fh5maRx77T7UO9CURCOhOUJwAVCCjvU0/FlE4as5Xmi2cM618EyJhqBYfF
aycVZt69yMbK8BHgVEZqdTiwsm2r74ugIW/Fkh2FD4tXTGsTqjEiG4AQ9bwoYrv9
nlxDt1jCMFED18A5vO56HzqJ39NezpRGVV75cv+uQ0KrCNibEldYbQrWq8yGJjaX
8CThJ10VKp+Njsx2S57T/G/Ywb3MGWKPl7vuy40WExIyuVi2IR+KM1CG9sNU/Tm3
u3gjnnMswj6cmOGpgm9dTpL7H5NdxBdki73im3H3MVpUfxUorM0oiMGCjPmF+soW
Fx1je033gdgmQCLvhEVGUMe61FldL5zaAB62AAPw/n9Plb+uO6IoneRPC2PGTXYw
zvg6uTKa59FM3jslAm54Gj7LyGL9yeBxxa1uBNA7TspGI/c6I45SsWCQmSISaXj7
ojFk7UawEE84lxnJsXGwIMseUjNtRvKt3jRzm54vC0Xyni9EVoSKnrNZCGQZGiVX
N1aL6ZCrV1kY/dMV2K0ObrciIU1AAvftHZ9qQzxwLQlUYwyFXSqQJEOLKPhuAXwh
1zFDwUm05+w0nnm4DHXahzKvU40ZPvmrPP5fH9j3JzVW1vPnUAFNRrFE9sniVcyz
3xpq2KvRH6uHBE+z5E57Nw25tfiMjYoxMmXF87hmLEE2ajmwoItnmqmY3PvaJRW5
AyLMzSQOcQmhlfWGZVQTr2eq5JDJAHUfw2ELW6tVMNEMvvqnxF2r1M3J3MPlr/Qd
oIT62l3QH1vpTbmjX976/zWL1SvI2am8YPDkwI/uIjV526z3lSZP4NmUWoj88mIn
ehq/YaBsWlUsbc6M+ry4VYkeRxmhmzA8upSQiG+F22zp5A15q/DUEM4yt3bzhD0D
tE51PsKAzKS5nI0v55FavFpvOy4zDvaxtsy5vbPz4TzjV1IHmFIdXGdHWFneGFy8
Z3RT527lGe+hSBO6veJ4/D3MfYjCZhRzXp4YpDwTIIy0IAfcCXNu+Y6cJ5bipZEo
D1qdJVIQbqjPVvTC1KmBocUXsIDQB1icMEF7MWvsAQWSeWw5fCYIY0DivHR6zjuv
dor+mXPK8t06/Ooz3pHQK4s5Wl/RO0jHsLVx0M9NpDycGn0RtZZx4Kd1O3AXBMG6
aYieCFcFywZNbVrcA2NJzjnxoFk1TEuFr4ZXKtfUUXLpwppjsAzMcT+C6mtPYWmj
iwWs0n/NYSWJxgFqIW1DqYoH9D6EuYc8+NpJNbxYlKmhPjhQdKBY99cGVfxUYyTX
I/Xe/VAQSTjdMwy7QSNwkg2yDqMn664PjcFwomyzsx2CP+D+u7jM8x06K1zmo5bX
ZVzZ5ixzog4tiYRPByrLph8mt9hcyRWm7xUzAqw8KW+0+NTh80Pt/NuxlTfosUqk
JnTHmJPxwowZZs9fSOXxE6HTVqUfzthYbkgpTsn8FdZLL6GGrhzh61hcKvhZ5PsK
q3l7cXT5QlrhJPBmDclLwTzZWsRHXpbJ7W51RYus5GFE23950K2SX0F4sBSYgSw9
zpMqh73fkpmOK4/DlU+qMN+JklravbX8C+rWRKWBU5l+o0o47Uj6STX7gOZArq3E
Z7VpusKpmVT8MMOV1tUFouDSskv88JZRZbRPxdlAOs8E0WIlS+lAYoAv8ij+A+vl
kkdmiC0GgOEnjv3Ff7xz4WjuK6zJZo4WmOU2qh8bFodkbOXIHkNIBifruGCPORYY
thp9gTsjjhdqI6G53tY6UphCjyszQ7sQhkWeEVS90+/iJkDRlwkaFrDJ8EVj45Zu
m8i6o0ZgutID02btGvNed9NX0olCFTI8+jxn8kg7+VTdm6Gtkyn9toE2l2ZGVlDJ
2PymCJnn/ePNxZWfH6mzfRUtGAB3TqmGVu9VDMOmXIRKRd+YrLUnZ1lTQUVVqOQA
pZRV5dWyLXkpXqYLndd89n8DN8gIfJLQXrEzGQ08YCH2ogEOM/tRz798wBmYMDwp
+41oLQH0Qvw/X1MZXotXUuQRWnqlPddvvXxcSeL1LrJYyWzAr3y3LWMKveO3Lmmr
pAW+BK53RhusYVI4S1wCqo+dnvEr0aXh8QKBMFaYc3+Kbqx5P96eYi7Xz1cheKE1
aKIsbdMrugnxY19TxacX62kpkyvvm9him65R7OpR2nwAE4Sny0LS9qGPXTqJw2m5
76co8hClHDS0/6nnpodANzW+3jNxO3AdZsTTCxjf9j3/7MUPivKrnAO6N8BR6qTf
MVhvv+UE7vJXrRD9MkGI7Tv/Aq/mCxDuHnVCi+AoUBiRQ8O3OjOA7OYk2xgzJTXm
yj8yXbw7O8j+lE0sDMZ+ZHOdKf+HcCPJRa7eiIikitScnGuE1z2dxq540xWQB9VH
AQwAnZX57XQ8kybj2gTz7GBBnQjsJKyfWyEfB+tOJVmBXftg4srEAy0iZuetHt6R
83frGrh5YsOpGu2MBs84WdFDRWfb/QSQjD59RskmMohAOejW229uZCeGbJIfSGKr
fLjMcwN3Xq05TK/8SGcLMXeVTzDCe/WNOs7ieRCtIXFBG2+vi1hs+9AXPqaEF0JB
Z4JaQo1SYkCBtcFuvF5EyxVT7WDOhErjYWEmeamjbONxkVCYXYxFYIo9iMY8ceGc
vFGvH7/efyC3Wuwn3WsVXkHURwmof6jyklIn0bD8QUa2u98NTgKIlYLPMQHoQ9sq
Mt6HUIWv8MUPa4WwKF7JL67GrmcXNiudQKY7JQJv5b4w4Uw/taFvaDHrUBIMhyjZ
0BZroxRi0VOF53NUdURHZiV2Ha25Rn3hO/RAw89cVSj8FigZEabvyZa4f6MZqcxv
meZmbK5fpl5ZGINSDbHogl4OL1fcq422y+EXVS1xT2k7Wry9m1e10QnAYXiKI61H
T1/Eta/lT4Jb/y8aADW1VYsiyzu/0+3+CAx9yxmtJyIqhXDkptevYbj5WbVhCQJS
697lDwG2EJdCmaBTOw8Jx7dt1a3sS7lZInHwMTgmb9JWr084hHxMEwi5HUf5EhG6
yhz5TWfPZ8t6fh9wkEKZcZVZto5oAd1msMTWoc8cVn2SrD1i2huA4g8RloUri/ue
SIGFw0hb4XDMZVHoAf1br4pyigoAgLCayPU65wrADmjr3fXEF3eH5o4PghwpUgUe
65F91Ytlicdtd9SiKKHu4bJ/E6WzXKplvwY7AKSUReCHq6GEJTZ48r7Z9dq3IXeX
y+q5A42tAD+KL/xGTfQ1pPuwrobxPBI1DKKei1D8vWf8/PUhq+Je8j99mPzpKK95
5GhJKipUUMvS/Z/gnqnFh7a8A4tN6AFOmbj5xb4+lkae6QF/dtyOhMHzfaWE9U+C
TwGbJoGS45Ex3aDz6bWCtBWGUvmOJz+ZIgBTGmVjfVYKSfJ/0jCEnUhd+gDsilxJ
Z6Risf/H/2siTATq7BSzLpxXtsR6P1vC3TuJmSuhZWwY8h4QG7cZc+2+4AYXsr2F
uMoM39ngaxpq3a3hfRjhTuV1hODxLbNWoco6ktaDkvOT80iGchFwG9vdAOLBlYR1
1EZcQWRE18zUEUQWMtH8MNU+0NfA9X+8FPf5JP7bGQKJQP7krG8mKN4D+Gc95YU/
wFFsUDTtOROc1xY1OSEdYp1VxlM6I5xX1+4H8bPa1EdfX2Kmp2fDmd+3+MimFaAk
9JwEFW1A4nfS56SrmivKv2V1C9gakvnzVohUIWwW1Q+/eDF2bP6rNTY/hQ7jnnfo
JhQcZvM0jLY4bNcMzWW0AYclhOGQFx7VeonwsuEOsEVDo+DoZOjjIG5kJ/l0Rosq
gsjacp3ljFz7P0pdJGLHpdt/00QPpANfzSAuY876nvl6p8TTlmEKbwBqWVN6YZLg
178423YqZqb3YPaLByVbaW28wyB16dj256ggRHu6xDo0wdojQ5HBn3upV2aZ5i1f
IqXodRqG5ibZD8oSMAyJq79BDdcNs4D4Oqj1yNdEoC+VhtYZZ392Sgp2g3ShDfN7
phzBPmywKfu3/UBGylJtgx8sJ9B7ELkuFXmiUoA8DGaV42SvYcdW77/N+lvNXp8z
RlfJBhgLhtWy0Mnq/kZ+otLKOWBUz3AIVXou/8QkdLPh3QRNoE5r4VksxXZAaVBS
obkVPfO6T+CuOvU7Tw0aTmfXwkxIRr5LGvBgFL9dwtl4wsuRy7BcRg2onFvWYYIO
EGhB1TNE5HEUl67+SrnR1CpPMFYY8Jo2fDmCHB60pfoC4oUebvYKvPAM5T17iC/Z
CGDu5nH56IlJL5BcfpsEF8en5wJGw7EDPyTo6fMJ5Gt7DUS06LtmxCYfeWwJDCPE
2YxZSCfw+jr7m/0tbKlr1P2kbYhqFZhcbHKmm9UEGlLiwLNR9PD/GnO0fWmkxoPH
pLLvZgSLiD4IdomRbRODSrB0xbYo5jT6gluXCuKtG4ReOQb/jHXQB8Wu7vJSfMc6
KUXjNY8iAp3TkiWebezQS05tbo+0ux6+/ohqAkBHFL7vgHLFV7ayXhQ3vdFxm6bP
0k0nNIskBggQkuLltA99L41gwr9QrB2B2/YzaV4BHEOaafBBQtEknwIHmRoXQc37
xQmHbBGkYSNPweGCDV/R3S/z5uIzyMee7m1WbsNwtoN7bBLjSiXB1gSWqHsjvHRi
8fZ4a+y/1/uIECLkHn8pO4m1XleVXB2YpsjeHBuzWEGV2ysDaWU+ZgPhns99if6H
Gty+wkWmNiXd9YpPPwgWitqzisQG71nVYXW37gRnRNaMZNJHfc7ncffvphDqvtzn
5TKvHlEoXyOBbLGB/+6UvvOiSsiKDGngjBQtUfXitXedSaIhkwCn/rQn34yJ5ebG
jswbWlHfvHEsqBDLPMx60Kh8TXxvUmtNb3K3GGBsYQEAJQe2p2mSRxCiHoyVI350
TX3sRCcR556xWYkZ44AmyGJ+IaEykWaBI+pyNBfJQwmazKlFMkM09s6VOw+j3t+N
nBDmogo/evaAX+fo1yunvgjO1ja36hf3AVar3ONlFYaBAkWhlSWBasrlsnM3VjcC
qPcbz8ms7XO3VPxspeSvfW4BV9V+98Lr8kTxfrnxQotRTVxDqTYtA8cIigkKbEMj
YzybPs8oqYPNhxFth7rjqekuU3aDRCHzV0jDu9Kb7WLV1Bwptj8pdFXCo9OwHr9t
YVnjJIRhuvxbrlNAmaY0O6QlsbMxFl6qFaVcR/YjxCo5JDjv21sgWIdargySRube
wUXGr8mGvc6A8eYJusbZt5XImbHCSbbWPRxhO9WQBm/oKiiJswD4wWl4lvnfYuzj
zjlYBTGmafPQSN2iui0D25GbQ0E3wl0ZsjZb+Hb7s/iXOB/n0QB7GSLUyQ+o+GX0
pDvmxYFSIw0J738xv9FvJUksNxW28pi5w6xnSF6TlehBl37p8RT+mbXq5hznhn9l
qHwmYv8IjU93XXIQwejBq3vUHJQu6uWZKcIxt/juaGjZm1UseUHflVEUIQmvgosE
+DiDevFZWJYRFl/wCpe5tCcnCWJwCXQl6bHta5kri59U0vy/frbKuIM7GO5nF5Sn
Ls1xG+8MhZrwMP6sIW5RjyhKUmuyNS80p9psaXDX/f+tJAk5FRXPIilWMRFJj3o8
mcN6f5xrBgkqAt+hzKns9W4EnKrr/YEj2bsFUtp42lXt0JMNzxPNBE6kWYzxqmma
7DfZS1riNzcCiyqrKW5AeWlgIJlelxf6XPlqrqURtuSdBKvoHQFpFqq3awJ+E6Sc
2vaaCXYap6csfdE2kDXkS8Vb9+MKG8EinIGv39oydnFRb0MNgldUETURR0S/kWuN
uLUtotb2T96X9P2PoPA0iFJc0zFF3GRDcmL2UFPlf7U8EIlvPstVw65brCiKzozp
8Uog0Y+LNeSats3VDc64llOaUll7QlYV/7wpvjs3ChJhzX4qui7H25L0ZCYFRHtT
5S4Ln+Qvv68L2EwCZ+Xt3OgGQuX9jqzsuSVGsxoXGudUk2kULD3D/UOKUCYtTSmG
Wzf1rDC7yJdQnBrPH1kdYPqocuBclFYlSTGhSGNqt/uuNg5FvOXoL8+enOF6IE+5
WoCeSAsu3UAPfdXwBYjKROtYDP4WdnXckI4FVrGeW/n487CaRrxZ5l291ItikVf/
Llt2kCeenxnOmhIhEVvaqTQsmbMNUil42wMtI8KGB8WjUh/RHiy9qY2vKSjavBHj
1hlk6ODm+9/UD636EyH5bZLsYrym1yZDXo5ukwtzPgYrs+Gkn955Y4TJwxnpiU49
DZWwI6Da5T6eFTlVBO2HeOD4VpQZcevWeO+NQhzd7KxBSVy9FZkqbndiCfWWWQto
DysB+YR6Zdhuc/hGBf+cu730ww4mBS/rXBJvjvBkqeSdKtbTLRNmzqXSKtGqcs7M
0HprCY4RgyQ4X606zVua0DwEnXG68WtRFvw3kW+66SWtkNC3s4sA/AhnpRyiwwEm
rt423EDN1hWRz0nzgaDYYrvemtTNvH/CCqQsyD+SAj2ZY2yYON6CGJ1Ok9yWoPku
T9OS+cPk/zlcvTFh4lUZKYknVeXQus16ZyHSwCQW760m+yigz30cAm8u/u0laL7F
hK58uZjWiaEeVJUT5GMW6lhefhX8cC8zoUaXyVc6Kyr029L8yAhLl/32jVDK3Anj
udqjH5mz5jqtnU/UBfobSfNFy07IEAfHAQu4uMPVRzf60iiY7YS6IXRz3uInAhPb
Imji8gOhn8o+MWC/hT3SSQXBClE8MKtSe5GbFY+T6UUvltYcXmb6/qP5hiiQajju
Obocnr7n7ep3sOoAPb0lyarw0mJo0VgqoIdtuVM9SZuT9a3few4LWUUYmBy4+ai7
CwvZ1VDVHTyhpwA9lNUkyqTAJZSvMKx4XHTF3lE2Bj+Xd1zpPkJNdLndsj4yfGOH
rhvSe4EBgYhqRi1LaoFQne7hMb/HqGnu0ytm6mK04rGVUfCKUTb1HXMrvjdr0sET
XY+Htif2HfrgBARdcEeGbUp/YngaJ/57cqOV0CFziBAwogizLXGxXWdM6BfzRxUF
LGRWFIvCrqp73v2IJ0+M/opmB0sBwVp2NWZKbR2GlM6paD3LtsRxn+iHAOGGcQzT
u3odR53JUIWYobV+y0wYueCEQrgX71sTs+VuaYnm1Zdz1XTaoDAAhuBtei7FdEr7
U10hXJhwK8z19UlRUQrZ6Sg0Rq1x/9TxzLOAX0hY0lc94LBcNl16CT2uuKtbH/9N
hZveCAXzrHnGi02LhmAJoHDXRecGSIuQhZGX5WE/nikgdViajEI/6hnhaVCF8r7t
GC/oHpk9MMYCiAteY8+DYv15Bky2vzuJhfsNg6f5RlTex4lIzOoNcGeB7PfsRcli
Z6lWWIcIIygraf/VturJR9zUEp25CQxaGqU92T/XPg2no5fdlyGqvR/OWXqROpvE
GVUw2MQ8SwlwPrEXrfW9bkmSBjQ9vWm4LtArtfmBKfbseoUH/2trzWzAlaqlB1Di
/z+OSVFlrCTIde1D/oEd0BY9b2L5e/KqCal/8UFATP/30A7fPSWDIumjEXiz3KZX
ExYbzqLZ6f/kK9xHICpSrQpYCymMpBEvWXcit5q5Qv7MySlfn2c5NhyGpFhrstyN
Q0zSucLnKsR2lrv8aC0ERQYd0B45tV3D5KQjRVUQ8wkKPA25nLUeFZIMOlEYZRUD
HydE2sVqq8XrTYo0dZdnO7MaMywJBZZMImy6HIVCB9cbYmdSh+2QfiVAhk3cuNfb
zm5MbQ+pBkCXzfSmoO8b+ly1DThD5xSi5aKSE8Q45foOiWGft5OEdMl2tRwVSTuG
XEGdSE/OFpD8BpDRK9HgUS9NNAMmmnns86EHcGrgJLXKGE30lUrXsyfdSDFauuiR
qRSWkv3anAV1KQjx110ilkvSCsp+mGL4n1Wy75uAljdt055m3E4g8Sft730zwIp+
PegZS4U4uUAbuI3zAAqC3CljFE/DER3N55gDu/atiNoFImhnu7+lSXy/fFQOwHRc
VZXc+Z1FlIClya5qiDDMikZI6U8p0MkHfUZenkNjEENoQU4QPRnf5tEhZoc/l5WW
qHLwQVDEbkmkRtkS6IKiYGo1yzoOR0vRKFQCB2uJYzsOqEo2wlMQ/wdJk+LeDx9g
09g8QqVrE0nXtcGvCLAXCCq8gu6pqaK1WqQCDMCRtlJpbtgYlEWJ9GNe1Hq8QL1Z
ydB7ufSPIZCRQ6Q+7IGlUYkn0wnDd2BVDr/0LUfXj9vrIQZCbZdgtf1eXP6jksgD
MbrUFzMAeRQt0vxXusqwg9pk+1/fKsJOET3T5mD7MbVN4qfUmZKdMxyzifkMXDBG
jk7jOwPJXssN775JbwlGeK+ubF+HQ/L6n9TgdI6cT8jv2gONs1eeXB7qhgwj3BCI
K+S3xkCZZoC3PH7b8qAfmcdy7TQ9FlQhzrS1KjrK6xIy6FOpHLgan3sMGYngtBo/
ZWA2rsW2mxf5J70ABUwoaJcp6VKxCRpTnnW/5GJ86YbSbgEAE5aLodBAiEewz50y
925xlZ2v1gfesvXBau46Hotuw05qTFuArvj6cticgG0woB+KGu9LV6rjk5StfVWr
t6yWQcsMW0XbtrUJfEI1JYQtgBLTdqw2jkUkDuPtcrV1IkG7d4gTy8W2vsitJ4/L
tVWqd10glCQekBZwpXSKCrV9Xm7EhFrqA58RmoJXbB06aFqFi8kZyKvZgIL1JyvJ
YjKf87SRJpyMRQOzlrb+lZDddm2nKcrN1tL64L2brzS1chlcfIU3EHPA2nTA1IxK
VtSytF86lCa4W+Lw0yXU6UIkTCFdLNFo8Q2OMkr+72E05ABFsRMMKath55MetWPn
cuFvVLPSnqcKNia3gmTtm6KY53LX5Ez9X2pWV4MeTuiEJjTWvSRWeG95hUDpKI5i
GugAZ35JROWT5sZCRDWVZ2yw6/gpZiy2tbFXkvZQgQWQh+sFjpsaDLF3IPcnJjsv
L8WxW8GaiS8Adaj+Sqh8qWJg6boKIe27pcFfDoh22z9YlILIN/mxYY+s3aNnwsYG
l7tGPz5WE0+vE7oMXvy/9HqivfTBKHs551zbL1JDvOIC3kKol+1XyZWAGPldQMGJ
LMce4C+NPIO7DCW0s2uRZCwZ8krLuQS3EGed0+FJE7qCxAbEOCRSEMMx+lZIAvwt
lM+cXFuxFnerMsuUxPFB0pStxgYN1aPTlcWexFjqOC+yUDgoktanKmYIjEAHPINJ
Jr/0eeXZvE44T4cxgYe/5QnQHMB2S3o3aNDuEkoilIS9nQlJR0tA7TY7pQOd2OcQ
rtOlYeFKAB7JIV37DHUX4YGVpuKLrlpXz7+e78Qz5wHBuf+L7bqbGTWM05WZVXJm
WEHKA8t3wAPjX5zaClUyyjEbNqmUfzbNXr64bN8UNjrleVKpElGx7Gk+CJAj7E8P
zh86aIsEMWoQHVZG2YEpZ3KLk8VanckLGwh0RBVequm2DcqN5Y1n1jp2fKKISd9M
W0hcU4yO07c+JPC/llpL2DqHp6aXX8YjQdxAorXwY0FLpU1gfzG871NhHC4CVo/x
nBfSGQsLY1uBvPnbGHszFOvzA6q8pWkyRjcHK9T9EK+TAzK3/6vYbqI59UUPTXUx
uEzPj1LnZixL99hnWNecEU1kIXnjsIbx5Q3qz+/NceE3T+BqlsvcmKWFSkC0Ksee
8CeaK+v8NFRBzH0qveqz2WfClGOaDfamw2R2gEnpFXVjZmu1VUxUVlNT1n7aCqVo
LUWjtml1DANaDdc/CP7VJmp0t2FH/ZqYhXRQ7KlCPLswUUhjr6tCxsf6iMiS5zN2
ys0YekJjDU24S/ClRqFIp+L86VSU7W9uU8lB+ov84mrX+WMzXY2ufFl+vQ+fzxqs
GrROLIyN2TQw1malaVSQAtBaCiMiAlyyE6tHaaXviXDlf0x9E+447B6z+z38EPnc
BCuxeD1ChFvjiznN/Xnwv61Qi3z1wyJ3oEIj5/jJL1bhFTuADWGNTk2KmvBEugcQ
fXk6sJNFlF+dQ3Mkda58KPTwghm+1TrHOLrho4T11oUM1rpdKc8cNeoY0OMQ9SLd
URC+DSQngS7KKlbrxKeDK234eCF5vlvS4vrQsT7ozuTnPdULdpP7Yb21ppkAmKCq
rG23VmoBvr6KeGhnBIgCvacVQZXn4osBv12sPN88ccbeyMa71iIQMDSVFe4cOYul
Q79JqoCyWcdWzqnkW2lK/11IHgONpnLL64rGesW36DVu/3b1+BB2MXXAxMOofxsZ
hmkyOqEtAiNNWyCwfA1+uzwGGfH56TDzopQ66hbq7eqxzRmUpoIceHxjkLm/uYVU
IboJEY8FNMLVChVeypZSdOwt7CS8awsQNXO9eWKoMyoV527sPCxiUg0W6uWCmufJ
6rVTgClN+lBoNP+q8r72gy8HmcOI/qSvhvm5boFmwIfToWHDwLtgBftkBvlmh8E/
ikCSAW89Z+L5O/qzrgimtFiqnhJMGPRd9NpZvuoYd8748Ay9IEreB6WyYqgn0QAL
d0kBh2+mNJXt5jTlRFUmfhM02WdCuKA1VoOVfJC0EkJlhEWs4Rh3AKWoEF/bnsG3
2eI0VTFF95saay9/+CS3fHaNIdtpakDz4usJYP31zZCWaBGVAIwC1goN3cR/QT9p
K7uG5GAEYZzGJ1/9BaghcQ2wsnmVh8N3AVLxeCAmuNX+EbeKYhzgCrjpgZYS4bEJ
zk98Fech9KjA6fThNFJepTt0F9YM6mfNOGLhx0WBsExTGGkfiaKF2HhYaMzliILH
8Lf+geNC0XEsXyOkqpKSTYM9nlJjPOQvGe4vNv6J8bUskxCLK+K8CWMMa5/CrMUZ
5oecnb6JkMERXpWT794LGpkVKW3WLIzS/StwQwInZ+BG/m+M4sv48D+dsmyu4LYV
+5pDtYYleGwnEFsWRGpIDtPtoO6DsgTfloIBv/ToSJ7GCRWr2jbJPkNnNZb6wKhF
lwY1XSuxO35jQhk5eG1m1F82NS8YFiCBW8GW4BW/tcD8GNDibMsNrLNyRqWZD2Ji
qEFkIGybonIs/Oug3UmU8Urc48JZqMnK9321cN3D6upSIpvp43Z9mgSfAiqI+vE9
aWmb25P+dZSMZyavsJNsIbUEt9YMq3FgZQz2E15Avv5wRYioPMAnSsFbv3AgqtQQ
6/H92BDjnV3lxfmEEvxZSVQ3oq2ZjrfF7IOpd81++oz4yPoAansNTDrdV9+lQY5K
63PoS1aHV9VKBhxLd9V0BIfo/qkhJ48LiAft5OUshSkrn8TXkZnvX70Zt3TuHZ6W
JWKc0IuEwsyVhznwOw4RLfJoiNvL95ST9MwVZjCE/8spmX22RVrLuoBZjellDsjo
T5HTyxsHpkjU0q3VNrJndQ/B2d6yok7LIQQtbXeRGg5ZlDeKAdYKB5PBLT818jPu
IqO4054Ov7lqSTD6cO2KfcOdQuWYn/i4e0stGWX+Ivr/y7yP+Si47ub0ZelLcTAI
Ir/BsRw8++lc+g7p5KOIgVt95zcOHzK2Js2Q/cDwtcWJNhvtWAPuxjGT5oWKXDsn
YTpXVDdThEW+EtBr9Ky0Z39NW3CFv2gHnH7YDCrZieD60xOC8S9zlGcEDFuisanh
IgZcrV1ibCiLkVCSm4yQXkewBCLJNpjia7EPHkWSjLlvnrfDSIGLq7wYj9Tqvh8j
zJoFk1GbZZZ4k0wBXBipcYdlNVxaFGEhoZnhQS9VdGRdlA19218948odjmQ/yGmM
xXrFoE7dS+6D8CrQM1QtJTMJP965IYmbO6qMqMmx0UcHKdToqU1+hOMV0XBGSBor
WavBF9847si4BSrDBK/lJaKvWyckNRngVntHp3dXRMTyUN5wLQv0Idsj+lXlsmBw
cPvPcz1mzWIZlji6A6yFUhKnZ/c1ihKJCtXULvnRvwVS8HoErrGbTdlI/2DeRuVV
bgyMSrF/HZhxJT0yPBZD+vcAB096t4nZXA8JvKZ47C+wnqg5mgTVxwts7gqcZpn4
SLO381ZmLC5dUcdM03475Wo5V/4CmYfrLmpHF7i4HYyHMFGDDfC8lbLGNmaouEpi
Cc259gIr2osYplzzMvndJFrYQ25ENfr9YGVEAUHl9WNyFC96U6UOM/padSehrthj
2Ox/ODjSCJoyLtMI8RjWf5821KlpMf/4YDbpiCZE7VKmq7RBU0Hdc1C6qnQrBXqJ
m7C5g89Z3fq7Dg3kEs6k1J2n2u3P3GDo7uiIuQ8X1TKMeM0xju17yl9oiWvu+v5O
qrz4kLRIiSXe4RuCLXKAoycR3DUYnPEUKYOcGvzdUatMf1nMR/AVKdPANHyhYH5l
LWKU0uHLr7s8hfh4IVK4fVcodhpDwWzp7uuIqqMqe6F6usn9+kmCZflkgUY0gep6
pMyYkzUmSqxFVzaqUwnP0ei90KCBzvl+HG/ZO/M4vMxMFPnOzzN4kQBlEOiBJgOx
LD2fYnTFrUwATkdnJJiylhgWes75E9r5Mk+C9ZTLqBEQyV9Y4zj+hCPYl6V6CSSl
zwuWdegv/nNt+qWkS8xZ4YSM0XzN16LL8fLUd2a3pZrx2Gpa6E3JEk8fASRo55a+
aiQF4VHm6ow5imNaTLPx16xIKQKCno3Sw5FTyCuL1Q79BrgVMZeuym6Nttyr9vl9
D/EUxu9ZuhA9UEHoH1lsn6a0LvlEVARjs5StUc5K4hNtQ1uPeUQIyfuiQI7bP1rm
gu4HMxBj7PMiJTAmeI9Xz7qyMZ7M6FQYYpKF5UNPWnPdVGtO/ZmrnkUV+yt92+bZ
RX6DlN/ugkSjADn5tQFRyFAJHfMgmWpa5M2KF8ByjeF531KxPv2clDVicDGBqlG0
6s05Bu/xq8JVUXF0hs54gbxuodF6VAjpRCBPH8t10Z/b71QwYlxh8+hRee1wnm7W
oa3ap8k3oAXXmtqz4l9yg52g5OvmvoE9ldI4uQHk5APan8V8jvc3ikjywQmYr7GD
y6S0CtU9YQQnd9owtSUPAQzbYG0vnFrGnByEd86O1KSahjdcLUYf7K089F9QlR6H
ZC8omAfGQVKTvnIWtAcUF8NZgvY3DmePpr+Ui0IgyAu8oRqISp1DApihDFc44hB4
sIcXGd4NoxFsJyrGevTiPSS2hZchAcqJBorB2zJMgas2wVNkbbmS1zFUNEoO8X0v
m+mfZT7HICnON9+A4i1PKggUHEFhvs0Pw1KTd7DNUeZ1j2z+kJrApTjc9n7JfbU+
tkg4J7JUDcoPUlLyZ8vuz0zhMZNbMmrjTi6Mp5syso3rrSCf0iN9ksRCneuqgXQq
RU8AbbC5JA5whdkaZ+pm/sH11HQFq2t/B9Rca7b358d02PhoguRmbTXlIiEd0c5Z
l1eT4OTWV85TsDJfaNCBnREWrXBZ7odPnQ602Xpw1E+pQFtwG3vxPl3k0C/deps7
gUrYr0OKKhB5BRyr6PTWCpY197WD08PIXMNsNEV7zWYTDNAzi72QwQrruDOOUO4G
RNpQ1ntrRlA71Z0xXCNP8uABRuy6VWC4xWr9ypN/YJGQ4hzYsV0K6EDpbzAO2PYR
7F0CAj2a/1BzieThPxK821N4YDbCMKnXl5PFQKOujFdY54JZDqlYKg3fjy2rl3s+
FHJbTDCigbFEJgaUUZppRu62eY/vlqIW2QgC8/nCMzep7kX0LNfzH3c8LPPI/gM9
1T5LrgT/kuKdcKZe3pOBUhSgiQKqhlP55Ze1tL7uizdc0g0JPBsJA6QUTbE0jT8b
pi93JageuH9jFc7t1RWaxZYdc2bFvW6xQ52bond80Q8bpbCjCtvPF+UF0fbIzs+3
nbUKNoq3TIAoLURMhF7rG3VigTYDvq9Sz4kyIJbE5gFeLNyCx8wcqmtVYaSTAjWa
+pz0ZpqDYI/mVdtxaoxhkrs9dmGE1tMyD5QaSwaeFF2EJlA9Kh8zI6t4qXMB1Wrx
TZXvuhDgNRp4YPA9FEkFnftmT6IAShCPHi5KsYyRvjFXO1R8FWlCBlDLlGR1jWsi
yXfoQwz2plSlKh3lrOs0qMb71rNc+lPk26psp0SILys1rcgkojZkhWnJ/j96Q3qH
4eqhjPp7lBZMnnLAtg5KmhTynLLdyTwxjNloNojGuymoAVmQW/kt6HWHm8MqpI9a
DIQu51swZpSX4rcdN1Ud7/9uFpc3WjQH2GaFYAsgUY78bSro/5xRhiERYBiNRJA6
VnQkyvQ25UmFjlQF+09JA54rbUE3LXzA2Q+lI7jrBcYdhXrx5b7idJzML4er8m5k
b85uLSucLlwBKaczZgEH344GzGV5cWLjFpAOagHNSPEPI6fZc5HmOvB/ZOsXFSuN
iOQ0Wu2Ndb4ea5ZMB+GRUI2xeZYSGa7RHux7jr6A0/eDbJ4SRgPRM8SWeYtk1uyv
oD2OK65h7AOGwgsfkdlWFOJrLLsPHndNdEagrYhYYOQ/iAP9jLl6UdzPXJPrXlZW
XderuUiwHBZkOs2a83CEcjcx7wcIyZnJAiANECYmre2hU0NS2wBkOoZiY5Tpu30J
fUEO0+1+9fUEyMi0voicalBguJh0OnrhyQ6Bk6XNpD+jPlfkHdBsWTl3kfxQTPqa
JGM6d0oWUT+cyAzxl3vnMSniNYoM9wvl1Qqo3BPxKPsGC8d/pheS6wWOH7bL1IS4
Tgl67igioOnS3SaG8zBeNTYTbm7vLvgIKdc3gptZgdnev+yTkWJ4G7hqAGEnnlJ7
542R5l8FYPd963M9dokt8V/9jPejRVgR/Kgw4VqiWCmjE9Wn0jT1QG61kUAPgBgG
TRJVZSquJMAJ4be1rShvoZiJ+SB6koUXOVbCcswVBzzOZaIMT3Bg+ptjREyL1tLt
hUzsWuLWOvvvKbk8ZCB+cPTduq3QCpydyN7kzP0F0+v2LxnuNCSRM4uZSIbCKJ23
UNu4oSbhRL4wIvl3dussArpbUVSIBvNQ25ewkXh/i4Ik5zi2pi+1ShLsgH20monT
SLxSzR40++c6zTBhzE0bNke9sH4ZAKlsYwyDg1cAOKiKlU8KwZLfcLhMjAeY/cH7
9URm0RiFaMcMJHfnwsu3bRYvIFCDW98zky1SKOeW30Mcy4rOVYGg6v4bKzpKLE9D
uUg0d4VPMbFcP8jhHBYOqDQMBs3cD1N0xeo5gTt2PzNlkqK9RQKAFJl/2fhyYVZB
zgQwCTN8NxfVDyD2yESDfZCWgyDkkZ6IKs0g68IVkR5dWNusM5fZJtvJN5k1o5by
WYtkzMzJh6C4b3Z/42WzMy/OY3SCXs/+K/Ne+DUwT7aMd0jWW3JRBV7SI1BRL3ot
dlPIVp9xe/D0vKsyYt4Q/X6SqJ4DFexvePGyZ5YVzWmwlbl3Iuf6uM/SuC9HiUfI
PZXdMN6b8OMJBIDlBiiyrS0s9z4Vd0DQ1knZc1fILkyVR6wWtvdCLc2Ksiuz+uaO
K7v6Q36XzZ5c0usdeGFYcJ+9D3vjry/NFSGIvpXVSwr5TGn1YKnR8Em/dh/OEkYr
NMOeRNomA0wMkaswsZlAdoejrSxv505LDVRdxab5zwGN50j0FnWX5Wf/k3nDIS0x
g/zFm+PQyiDYo340BuHxae8avP0hBwu3qOpgdcw9pacNwSH0VFO5NRl8JLfTqz63
3VodMc35mSGOrOWZ5ZdXyUr3y/sL60Ywtbp/VtsC4fgpaMAhyF9nLN7P26MRhNsb
CkEIIXjP1SLydVOw8vBbxblxqmnQrnAi+2a871nHpMAIz+1Ltw2xjExKS0PhqnLP
tm/R5AdgqKz25BbuoptSXoTWU5tzgL41TnascIOlMJqoZteCu0bjRkGZmIREj85U
vvFc0mgQzschrAH+FxvPhNHqPrvEoowtFsoOQZ0mfrlQzT4AoXp2Di53U+tKLQIX
OPvVfH7KVuQyODk7O+6lCBqJb6XrB4h2jhxww5wE2ZsT9DSK9W1GKNTp5Xl/weC5
haPXDY9iaCsxaMbzV6NyuG7jlfT91JZNX+oR3A9LH4UFiDHtG/InRvvl2O6odEAK
tD9Ohamc1QvQNKDDir+mBcvZ0wlMzKojeCbsK4xls+e0qRrpVSLowJioqaEAYomu
dr75IOmkVM9bxFWwDFXieFTFPuJDV+DP0trd9ygqPwbF/Dev6zx+SqMimfnlI5IQ
Xmz2nJYs8QNkYKAigvJ/z34pjI4fjzHq1pytJeZnk2u30wkTttvOlX8o8dOo8Rn+
K8Z3QvkTxkMSeRsDhgWSdi7xuzLQX8DFRqPRYg53fjhNZ1VbMpryxCYkzm0vYUQ1
f1VjvL8EMI2Qu+IgKHqsGV8ZH2t6oUyn6vNJo015+4ZDEFvTEK4gCcq3SxCg3Fyw
djedIyk1hPrTcw8I1PSMX2vde11wnNsgVjAvoNpPtdNSXVonA7CbaLjWQ5vBdy92
/5EmGPiMZwPHcDyg8NAqqv6lF8ZsID23+GUv/f95QNTDytwUIpy49PAyGWCrZjte
JSSo4ErM0d8NItaItOfj/mOm0lZpyJ+5PfwLhVQKBM9bnLreCyTPRxBUwazxiADy
BX15RK2Q+ApNSeGJtmKRd6zj05/8vo57rnEYU2ycUiCYdS4bl23YAmfHJn9aNzv6
+ny2PwK+vKZq+nNT/tCBLRyqrq9vkkoF+RQMRfif7yiqzIHwSXJeN1qmukG0oGjX
B2wDDC7xWA0XNzsCIFd3mgauiyyCY1JEB9LuJ+qRg7Cz1RRp07DX0ceOuNnQpLSZ
vokA1MiCEa6GT6Z+BaKE+L4RbpOnKcmk/gdtxbecntOOSM56/5KdOY6LknvWEzcb
mLG4NTNyEtMckX9nPb6eoGJwecLZPs/4ZCQO319OE0MjPNDKSCYL71G2ocXgFvhJ
m3ZvsGKjXqw2Cwg05NlVUH+aXBSgEAmcojQd9BYj++Y3G3RufNpvZByJnapMu0fH
H3tlCOqDPKHsJjyBkedYKz2Mu6Y52XlTMAmmgPHJIp1bsI7/c2FxkAcoxfsGFIgo
DDQzzsygi2oza/icoySZ6JfRV7yudkZBXNP1efiQBPiSe2Lqv8phAjgywcWuE7+6
X4NFFhGPSRv7iBDY6ycFqa+Bylk7O/P76Z8Iam4VjMKhQrMJtiOF1+i6u5S3trty
eohn0KZb0uDjDVODkcHgl9PBFVUJ4pB88RwFMQWe/fcuuXs3/SoXxZhHYkTDGkDd
j78s6zbtQnvEnJ6Gz9VZmVV+u/rQrsVbFWzjIbh+wz72YoS8svEKYFGLZ+oo3h6O
YRRjAuVKG8Slz6Aw/9GZq+BUIIhMsGAfAS+nCHRzYaWxCGbJ/McYpVu6USS3PBle
6TeHAmanJ5lkUN51ZsLKVSVeL90/F3PRtrv9h3snJcJxwWDlt32J4e6dwl1ObrR2
NXLYTnbaEkVqLoKKoTV5VFHiLHB8qB8hPC/BpPaWclt8N/JHu7oqnB+XPt+/MsYg
TUYGxWRwVXjeok2CxIsmusSJrLMwIDvrXsx0Xe7q3K6zLguDEmmYXjz1YalLEaBV
7m6PiyBAKyNdwodV0dQk6P92kfKNQwq5f9m1gn6oxDmq0Q/uw25t+ITAnlLyr2KS
nKRD3tKy13xtHEXzNOWVdyE4ulcEHKTAxPPwwcN8Il9IETAVAbq7GYw/A4T5nwmn
bcOxu8+1Uf8NUe5B1GJI/I2kUGsHZXui/+5qj3Hwmh/aZ6bnL1kYR7uPm6CIlZjm
2BsZzdbP5dsizmNO4jed0SLrlZYFJNWBwCi3M+6avr4hxqt+zlO8jDScHZDISfA1
tXXMus2AfIQ/E9PnGsAKd/iJS/m1IInNUCwrDUc7xcGT84Z+dEi0S+qemmAjRjxg
e7StKXJ7u+ctz9mV87yCz7L+FDgJbZhE29tvAVt+XmsUcc5xkbvpSa3lJMstU8Y2
ySQ+IA6KYHv53ssN+XGrz20dmwuIfNBrDPlO9DMMt4d7tpjAvdgLTUPpnSsoEhK4
F6StZbgHVWq8IzeWWS9Mbd7ELrZinLyMN4yElYRREU0kyQ26ohPLB4cOKpS+9w2l
it7BiL+W2z+qooV80Jt0r3JN7B9VZVpbKRq5ulxeNjUffjrImIPqCbBwFC7veIoV
tmRa35k0U4uTZZyH+RzLE7NzXqSFjJFsZyjOClqKEthtsTJbofNoE9z7LPY/Rjt8
qomXf/mmFn/mJlZOPhwURtwPE/PP5gr55Efrqnvdeoxjnvo6qU5A0osQJ8I31PC8
dO1WU2L2fuxZ603nP7Wb85k/em74H3nwQ2aWDo7dSLqGQfsQTtP4rzZdaMljfSgS
8kHx2uoWCeTpAH2FP7eyDyiY6li2GfJ0zAF7sGKIz9Rf7qe+q8/69Uujp/c6DvIv
dZwf6nmxZxMzlpLwD1Dzz+PSwDcPJW956TF06uOG872EvF7dEJhC/3SSE0ziadeU
Ius2n+JjF88YpUeNq2Q88MIvrwhDG4ckFx41jByXIyMjGuBZn3q1UgjG/JE5wIFR
Ud+q2tScrMdYAyVDWGI9mnSf6ACPK1P17ep4Ds1urLCIKgRgWW/o5g9fnaeW/b93
isEPBjsKeRN1/WykK+IgC5o4sEbP2MpyRX1CZtqNvQX7fO7U2gUzD2Q5kIC/c0Na
zKenNUeEsPmMDyBK8mzTfHvWPu54ZF9zy8Jya0LPPWl2S/B4AIgFc4Dt149+sycU
VB0LPIYNUOY4UFjenLCRRvOw7hupGJ+hlcSplSnMSfELcrpr0HlKLlAjVRJFGQdk
DPWW6ciio7xxTNCMOTjxamKI068ZcTcAACbSha6VCCvfYCcygsoM/HX5QBOT9gc5
U3O+wAt44X0dfN1PPZvyrVW7BcBuwOaGOpfwCZVCQq0fsw7ri2BMGBb4KQAWaRlX
kOjD1DBNbWbFgBv3H8NomoPgZy7vfAetAyjXzUSQpImwrZDZiFWBV79BcuvMSOV9
K+NbuLhyZt6o+CXPw2r9DXLfTwPnjm8xhIwZu8I5W8usj0BPSj5NSz64RBfJ79b5
7cJWE8Iz0FvmvP1gNKP0zGfDJdPkWHvA/gTa5zMTvt1WlHA7dt27Eaef3QOwDfrE
t1KKHneICtx30YH++HuvgADg0atolDcZgyq8mmkdNGWmuww1OWOCNKskipGyG+lR
pQhsVIg9a9XHpFP26DBuvxYer6iXqG7i1MLPufEKS3DqiVHkIexePrO0U7yv8GE1
164GHa9llr4PIiTnQ6veQdAEdYW2kXKJ2NuhtfGJsrJQEsqKEIWG0D6jJz8eISZy
Up6i6KahZ2Q9LXorrJCdLvgVBuEokRujAhL6sAT0iPPsXRsSCWx+5cTf1PbTOuNy
CKrM2Dvza//Jp78WCpGuvQMGEWrEqgPW2nhxkxkOTzw2mWp8/5qXFjJggmzVP2Cw
7qZLBan94QmKdnpJrJGZKXnCKqghX6q/6Hgd7SEVhUFAf+TblTgCsVzZAmB2Y5Xh
j7QUw54JaXtwWaC1acg0CIivdsTRLwvzu9+Vw9xj5Q4626Tl42zaZeicw8trbK2i
x1x7WuJUXhEv0XtiCrGvMgGEuATihTUV9zOEWrOIXOVURotaHY9Dy845G5DTtePd
Jb6GobiYH4W1HjIa6g+2js0pIXruxjAS9QMLRdBNIqVPxAYPIMVQpSq7h2LZZ35+
rd99Y/urgx1toRwxPanF/vyM1rp5QVFwn755OFjL4ORX6Nqg1x+QBL2xgRdhvdT0
TcebABg4Ku9JON080q1dhzymiI4PsZ3wxz87l41KJhWs4hfS42dUOCpuYFtnU5AP
5A0IuyHTDvx56D3BZEsAEU5jIaWZys9z459eTeZ+gQfC5078SEm3IepMhOPASVxl
bLGTO+BbO7xdUywNw21JxwJiuFJOaOID+AxWzYyvpUnFIeolet+Z8QeFlUAJgxz0
XecJ5WxfQDAOdMgdYZddSmv/GF9sOtwvAqZdN/+QNIJxTxPcOwwW3a4OnZ2aJuRQ
KeD6wyFvqFGpQxffj4s1SSf0SjEVwCZ9GfdsIRHftULhQYSvZZ6IK/RzlFXNYA3u
mLXaOFEHDVxcyMUkmCrxgmX+tGcKBb4poKMzZdPH6vzOA7pqLF2SZDQRe7xVXxeV
oGSEi0gxbKMP+2xlFi4L1NKEgk4xxtjgsXq8R1gMP91Pz0lq5Kmjt5ffbu39YIgY
0EFiCOmdgK7z+shUU1Vms01iFACgEd22txv2h9Ov/Bbaaa76h8gC7nDPvSt0f26S
3hTBA0pHO/Ii65lWEul9AZxSjesYtdHdCorD9PFbQnOLAHxPky/zQ2UoNrmn89Rx
TZHdEEaaBR5f8jFbXrWDdv60xmt2SBdV43HRREiDOKHOW+pp119dxxG0Yp3VIc5M
u4EEL+tl4pMqmzBdWUUP28OZGiMxWjiA6SYVzS3FhvexNSyV4oE3Iw1rLe3d/YRO
v7ZpKfSKGGqL/8h/unaCOgONAVNfKBuYhNulphZmjj99644Mgc6JngXNcvDXcMfD
P60gIl3Jh1rQ/5vmhf2js7ExJ6x2nxYs5dK1MzUs8/f9INnDwnS+nxaoHft1hA7b
bzR+V7cqr9AYyQkA7ArpOY6OoQLQUvA6TsogcFxWNZHHbMF9NCfOoCtaiL8EVlzw
zQdBonVB+wkIF4LXOrXH7FwcA9hEXPQ1GEuJ97ps59ZD8MSZ/8iRd7+yxbaTFLrI
teX5uTPG0sE8kG1jHe+Pwop1c0OvnpOhIo1L5SdZqkaYi5v90i39SIXNUofNg87X
/rrUyKuYiisUf+OFwqREPBxSCmUSADBEjfgRJwjSurkjLNB/Wo/1A/kBnZeuTAQj
BWtJF7lFj1aTplX1bpgypNiY1vnBV2jARvTuEmQ6+V2tkfOkMIYw/0urBT+1ouYB
2y78aHniKAmpuP9eikjDNvKjNNjYmL/UUUL4+97a9sad/JZ3wGYO94cMA18V1CVI
wfCsBt1wYDEKz4lXmvl3rPgFODv5u6A7/Xu7ap41XGc8UOcJaKZogJP18/ksiDAZ
t5XH2OMrYBz4TJkZoz02r3kyjUCHiLjLJBnIJEqJRaLXMeOBrdM5CxzK9zsYhEp4
GnHbL2NqzNdKo73QqFHhqKM6Cd4/3DGD+BljO77O9pkBHj66FAbFSaHjHHAOZcvw
DLds4AMBy3Zx+wdY38xCDC9tpwfcGNJnaxp//prTTsaHNe85NfgtVdHhyaypVjWa
wvx3E7ear0Mc6+b/+lmH1a5CSvcmK5z8lsBLQDWFNQduPArfZLgibj+GB/89xL3B
vOcCaopJwZhbIJ5H8i/9uxME/FiyYMJ7SvdXM3wum2iBohxVQz9l1TZXYyydt5cF
fqjERWBnmM0PfQzGVAUntfqq9xcKKp8cVKcOF5mY0tghKi5pdQFhRRMdnCunmhU3
6AEHQLq665WxDcko0llDR7GqswYnciFCjf2AI0EJP4JXr/aXdBH4GfgHJN3iMW1/
4iOMWs++FzMNZOk771nFlOvD2Ug1uhQ8rvM1KwHCfOQJcN7D6WrYh0ho89n1Z26q
ju+cXl2dLJrQlg/+a/T4fchg3hl7XNDs3AEaGUcvGKq2jJnqBIkWe5c/YdaD1x0g
cdZKV69Ndxmr0ldh71lbZqsqugQTPaFGVelWSLj1Lo+4mARRw5t6W3RLMeC3OWcz
8IdPQo++6pHsIt6D0SertbKKwHrZk/y6joQ5Pf55l2ZyAg5onBriq36FIYApgprl
2RXTa/V/A8U6/w4RhYn0t6MFuBzu+emDhoF9WgLfS36Xxmls0cVisjY9YAD9apsI
BFXgEFcH2CTxL18Z8S5oBX/U87BOLpZ4AbZp5a8NpU67IYDwK8fUoElCnCkp1ibS
ehyhGQ/pVPQhdFurFVAvZHGp+LiMQJH9Y/IA270AvJHp5ObHiSZCsg3k7HZ/cIA/
YGxLIE3rKARyNqLFJcJq8NSp34EWFPTEyrrczN0q1354QEBRpbRixDLIMpe+EeE/
he89Scy0R72apbU2/O2BcmnG6FtFwpgpKB3C1Uj3HOWcocNunRmF9pgInDqAwB3c
PxxAxLkgxKvusyshzowJg7FoyrrNvjE5FZuomAvcPupjQqVXPLlMVkOKgA6NJBcf
CEdDp1qkVLs/UYPweH/svJ4KFBKGgOsDCQFp6oHuYWgJw1S1Y+GGyGoTfRK5IzXz
nEXX4CmfFji+fRdLmejUoC18sms7aPB8NTKn8SBM08Izwr/kb6GZwywQMPE2cgyK
+0MLo5kti1CqJ5MsyR2jUE7ZjLWKe35woeMpybsw1ANOkN0ZkqiaHHdP3qhfozVr
mQexnluev6l3CB5mRMLUApJ6GA0i3BZ364Xlt+L/GwCFxkPcHmooYdwt9q6YKpgF
Y0OPOvd9NESbqiGUH7ZNWlR5t+DbLqMVO0h/fOtaKiwexGhmfI24mkeqpdJvBgq1
MZmGuJipEg6cc8xorF5l0CGlCreVqAa1Br7B49YJDmwRV2X1sFI+kl35+nkfhpzm
itE+TiTzenKAmlbC4AMO8FsCjS0JQYakhUyq2i0CLsJTPntsLGjytkCTLCYz4TI1
Xvu2xCrsa3x6VqNJr1nuJbCYAbamtNdndg1oZt6yrLmulSUYzKSUCl6hLDsh0HVk
AD0SQxVVBcmazU6mAWJpkv9zFev07/D/efl/I4Ia/oCx9m33gL2bf4ePgI1sWDum
/aBqvqwSRx95LbE6lAia7XgtqK6X3jivGzPfY/9gQ5zBS6+Ww9VftaN+gxOrwjGn
cfcLq6W2rJyaFDIfin9g6md7bJ0pRl89cdWePjoedlC8uuY6bPUg98Zg5hhe/ejK
MjY2Bu67WWWS1yp2oZw9lTN+JkN0wxzHqIyRUpOwOlkKZ+6MvZ4h46hQze1KnKSs
YxS07/ANm9scdqUywcRIToXtlgQGtY5tC1xgnCyo3Lofl1UEelBucw7OR7ign237
d1NBBcYvJzWEGhjkrx72u3BXdCGROqCGYpeARihApgvGCBPHb0BHgrP58533bI3v
IjkX/udSXQdGaWwCY6GMDE/eq/kLQvfR6OtrQldvFKPXsIqsy/Uo4RRKmEXe4S3B
+CnbZExolhswH+FXnojpmV3yzrt8qS/9YGNF9gS8ouBLRBOd9YINzTcShTQ5WorB
QS6dXY6FTpChlhOfqcyhET6suv/bYv3qeXm6Eud2v8jDmwqjmKwc/aDa2Vq/PeV6
3ox/s4oQf4l723Cq4u82iIC6Wghyq8fmX7aiQvOXXJ/JqXT95LgNzv/pTuljCXXg
c5vk4xelRfqVeq/Ru/SwPjWivRhvvMb5QcIrx4OozPyOj2F8gxXOjTLCxcgc4WwK
6034BeYg4JhfuzAGID7Ffyl9U6myvMtCDRfzxFtuwJilfwKuhe5mTjRXoMnAItYF
Tgwkp7AjhAY0DO5dEzgvu2DqcgBsmvpKWMBX1ipAJNoB2b/Wj+jb2agto4SR1QHu
fqhO4CeviRP3bRbleNaTJdy7nv+vQK2oEfAvK67jLfF7HRMwZkaH7RqkOMZ3xvP8
1L+8Q0EiwfjWiQIEomMiexBARH/IGD46j3jOzSabEH8JUJLeGSUxGAMX1ZelemXK
ykegraI6jF3Y2alNtKQO9rErluNT4P1YZAJOHpdBpfBhSiVExjuAsVRfwzUH9357
CKt2CbkZEdIsZci1IUeRmbYOZqpuergS48X0MUsbLZMsNyfTq0T6bcDSp+8P0o33
WmmlI+9pZtyL4NjWHDT8199rR3OXZEsilzXdRYbq15GZiu1VdGFQJzdNd7bq0+f8
njhCstCdqBSdQEYExOQQOS244CR42G5T6HgSCzo5BgeBMf0OjmHXtf7/obJRrh4T
qYQ+taR4rvLq7UM9mmeCw4oBrXIHzOmGkXbrGMWkPazDYEoheQiJdzsyrU+TN3G5
NlO4s5rn+9OwCgLLh8IE0zB1pySWVhqYTFkWlb/1X6h0kfy4nxfNEjs2Y7FyMMmr
E++EkWbcAeXlrxGFmRW6oiY5xIV8zngm2vZ17d3HAjoGh6B2BFNQwafmovR41Z3a
yGGLPQQikMtjt4433zHxVBguLPtAAhI8GVh3szbVDaR5GgXBOEACX3/p9Iv+qW2F
4KQwfpyBlnBWh496OQNNITujmkChUKzmGMCrhDGxw7I/XUmT/OF4h/Jyn4k5AU9g
Iz6f4J/B0yCtqaU9hBgk0hkUfrHd8khuNAshISUU5fdPFVhHl0XcW3+iZrtpuliC
tGzQXZorOgOG31itBjY8JqggMcLwTGBKpeqbsRdp9DlltcBxOWRZfF5TFFszq+zn
ZSQ//h3Dvb/RpP+haejidsKcwUTcst/PsHwPnXS0zV7LNFM4f2tqIta5ZOiKdzDm
+IaBlGrjIVGrSWNCCESjSwEe7q73uNDsaOBtAnqn47CDtqkA8dDoCvcayK5nHdyD
lmaXExbSUjSoKaQKAj9zWdGKkJCFxBtkEd4umYle2x8Ok9Z7U74HIplgK6mSst+Y
acrZnfD/2f1NbneuDqTcPepwceWA2lEy3t4oIhe7DXLsjUbjhy+IzPp1M/3GyRS6
Sl9crdN80pbsjD2/OOM4AsY5njy7Y5srAt4WIerKZkw95lOieV67j4c5JkURJPdH
6SkPhAsLJcB2OQlPHdOICJZa8UXemlnxyncjgUC0+AYzYGQ2O0nxFV3kvRICuEof
CJnLVa+ByXefo1JWXbtlAYHVHoHSrJjgKm6cC11GtIxLC+6O+QJU2XOBFe6f3sRv
Y8Tmq4zFuMvCRRnH/29oisJTrdZOIwoyl7YB4mnJTcNjSX/zvA7xjzkVZuqjfu1L
NerXhkcwWkWxaZTMYaAossFX0yXJVDQ3/87XzntltP7YYEODs3G4R0TDmI2dzTEf
qcPChu7g177FaF/lGor9U26r9KYVEuPfJ93vOQJTTl3D6iVtCzjthjb1SVAVc2oc
knOFzyimvetGy6X4rQRHPgib+kXOLxgkqQByH7vLkx4o+nMIDw5Us1nDLoGUmLWN
/HykEMgcSiN3XEMfg2/fzhtvdAjw8F6BzVlJVaIUVz57Yos9v/RqHXvvtq8jw3oI
rX8itYq9PNbGjLvKkhdedq1fRkV0U475jgXvUmI02GcQlaGBkXwDAPpGtS5fxM9b
QgK+rX8SjXy36p0AxaFrIbdNlJgaXMWrUGOwSSydj/sTHMR0DhpgIe6HclC9lkUz
hKJ84IDg3HTc/UykLriBKB4B9PmmOD+5dpabSYWJkUeeWBcQlciqz+BoQSvihjBT
2dIjlllHwlpdbodGwEpJL9Ks6+bydjxOPXH2LOutb7MG3hJjJbQoR9QSKI39Rz2x
jbBq2MEfnKi4YlUypsHvuZO3KcrMjQNoXvEJLiy/e8LiC7WZI9dtzMIjfz9KKlE9
L8+HfeRDYLQmp/Gp554mgESUoteGoB0VteZvlWZR5IF1Facb/BMKDuPiI54GLw3a
Vgzn38+mN39KcRhTw0TMxDNGqssoNXlLvcH5s3DptURo7thvmqHwGU2TwS77IEeR
zvpqQ21dONz3igKR0H38P5wGAeAUKoSOxvi5md0DgYWVl4OSMclvpIA0+M+PlnaL
SCUusL+XZNTWtDi/bYcQ2xXGo9dqwEP+fYRsKP0uOzNgnOC2gbQuP21hs6DWa0J9
MDOG+7sXex/uMRukkCHhJmIGhCv0DDVhj26heaGv3J7cdiq7/qW+GvejytVOvdmD
DxkTq/wDTDWU8rdga92Xq/OV1RwVGx7lGbFVVf2McFZQ+denaB+EuEOaNtVv53yL
KajJQtdffb5eN1/haPeDLuBphjOXwyQV85QgomSlGLhFsi1m4xSlvfdafeyYhTaC
vHAI5ziWoJIw1pcSAfHCzhKlLYeH+2TsvYGD+rwhlA1YOD4mFCCk37IBTyb5QDFH
ALl7qWLvZYmbNP+iT2MiF7ZSFXYz4lpAufGUir4ikT3s4Nv1U8h6KypBwgpUzA76
XgOGnC0s6KpJrXuKZcGK8XIWoGMzoxW4bOC+KuwN9nPrBUjtkipSuFKK/fdZmyGx
jDtVUVC5A0Cp2n8YmWMDutizTjgcQZRPXhgd5s4iNR83MSrmajdfpGz3UgRRCiLB
xWCJYo01teAKMCh2sjJHh8U6QAqwzbYqJkykHMeIez5ZTxKArLFNOh25l9By0uId
YpJJb7nnBi3FZt3OaqqSyLLbJvsJI4//ZxIqAYJEbbJPXxlMI1nN/BmPPIwdrjr2
e2t58xTVak4z52iV8aJlp4nkWohivtXuA1dLZcHXkSVskNUov52AV+bRKTnpgA83
z/TKd5v2zbbVhGsLJ+v1zH6C3bLYS07sHc9Qz85SR/GS0nuC6sKwQp/WBJYC6FKo
yMWGqPsvWNpXV3o0g8Gnmiu9nOhUlbxS7kaktFhuTQEBGKSQOkLvpFvuzwHDzgUZ
n7PZ6koTdcrHF3Jv6c/xWjg2avPmdJhWUdt8SMtNY72+zBEXGPcmooTM5lDmdt2x
BFMZvWmhjVtjQNC3/UeeMxM4Nugy+gbqsIPYxtXK+GgvE9/MjAT3seTtSoWhjSzd
YtgrfFzNNrNspOguZuPmrnIRplL8Q47aDnzUwN9dD+ph/jxzvOK9oWjccTI+8uTl
MccMV03gAK4hu3cbK2MSFoJMKTOkufq9ZCQAzK92kL+HlBjZofO50Tv6PBDa9Adj
ydpUbcfp50sfn53o0OYa26I9KqpzOQatXf7GFIz22znyaNr28bWX3NJ/gZ94S3LP
uoUzKmyDg63jnJakGKkHamVEemYQa1C7dW1Ol7ygD5yfRiv63myzRd3JKHB7DCvO
vFHV7B7YfoAdSWUJ68yK4n5/n98Of+pOlvofNY2kKTMz5yeuFrEwMdIsVfd0OZq0
nO5+uoJfek77WG01U0QVbe3M7uya5uyul4Xmn/5rNNXP1eVXG/LufqvsejGFT3Ys
QdSuf2R/VtAaqJUNDCI2XmdtBoHA/D6zXh2HN41IvnauYW+xwnfnjvJ8w3KC+33+
TelattxKc8wr19tROuLlGLWR4pG+O/k87rNztcFlF4axEeMEH/Tr6FE6wntRq8XI
hyj+EozHr/pNiG8QnBhLqrmhzALeTwV6YrraAYV0NEdPjxIPrtjt6+vTlJeyp2vx
g1OzFQ6kSXDAdmgr3WbMwYba/VA3dwwRCxJ4FOBkVeeblxiqY/Pz7m3YttLhCUyR
5cYfXtKp1HYgr446BNF7BY99u32pR5iZhldVERTwqhAZsYqOAbvvHZjefcYmV/Vp
LqStSZeramCs0KpKsqamBLrdBz+QFW5ulmngxClhyeAjcrxnHaTlVUQFOsh+fMEV
iiUfADCd9mHeFzntg5SDaw0N1JPscuPa5kqwctizgyy8xVHDIiRk1Qko3ZH5mCLk
qeuVSJ11R6RqlNaZpXhzwP4tpOXdCcpSZ/Nf9i4Mpn5wV2bxS9TLyAarbkGbAaCP
V9gObdPUGZGgXWfn01icdi6aPpbMUjbm8qmAOETcGhUEZuW3EzHDWMWTtZNbYhMu
eSHQPpXSKwThCf6R81vAuuAYZI6eyFjr22MlPu9NcsNTRq2leX+RUU5SFa61ZI4x
gXvv5YJEaj6ioYYVRo9MpNKWLcbaD6CK+Ro4zNlgUHzv02qmEV/zretctSikI4BI
7tSm3pxmFwPliAkX3Ng7vmV1KcSeuGMQg3ueg0Vvyo/VzVzV9+GXAkdQuxEB3hdD
DPTOd5YBXntD4rvrkfBtBnRYxBSmp+1SZSyUbxIHsKiNEZ5OHx7bRFnkXaa3se1T
u7Jf2hAAGOV+MujsvZ+I4CQ0OV5Pa0Qc/NP64H7ZFQ5potebqHGmA9OCtZVmhis5
CZTK1DCFl/UznKTXTyhGzqU7TNpoeBhn6LOxplWKyLX2CUrSB8jsfsolfM6yFC+R
nKzIwUIPRFTtf/KwXuwJGfYANPSerpqfT6AHIWWU9j77mEOScUXsgVNEFujAk930
cyh9PWYGcXVt1I5Rb/Zv8Rut1vTLSu9yjalsYey7+qfVJDruCEAHAMHu4NzOCXIY
Diy6tLKD4JvhR0QsMG5mlSMjam8UxVnuSj41oYOuAmpLFBq1XZP+XS7R22zT1uws
y7Zc5IHoNAMw/SsSoXivlWoL66/6wPvfqOI9+Y5sc8hysp4SLKLxD+yIDodIbzqG
bnSAaob86OZNKaJrlXSOc9YlD9/KaDhXfNoKcABPuYkAzP5dKrkVnqWomcLIs6Fq
/3ItoAFh+n0Pr8Y0Sn6sg/j+TwZFJeoftcQTQ85va+V1pHpn4+ptqQ+sPo5Lv91l
g0AurPmHPrpBwaQkFd/bFcYlPVK4qz+yDmyHrlk0EDhm4OdoG3wpqFQwlizEWswM
WGor6iL0ZWYXqJ37QsfvUNV9RE8OYsnOoJbsnXk7sFpcwSDIsyMiHhzBxlg3+CpN
pfFScafN7xWyespVnjOxpY+DP4xKKR7g33UH22h7i7+4l2CjsxGDBwEy7rmOKlF2
sWaZBfR9KBVM3AvAAbOdHRSusxb2i02g9SLUosrIGjK9CTLF7/d/43fqKjdiPaWd
MZ8OnN133w45pVj3o7tqtqCffV4x/aumkXSXvKH31HfB27xcNfNMAxLlMjBgGKZu
FyLyelX2ptBwixvPsmrSBX0Osv5oqkyE89ahEDFk9X4zm1gnvuvQD9l1IbTVe642
3doFMRns/xRFDU23zOlNBIdTt+olcPzj4g/5OxxobVxdnzaYxQEQjVDb58ON0O3M
72lPfUVVEag8i1I+Hnac2XbxAnrxzSAlYgbqMbhdlfasJgLlFYDuqTEmPokmwlFl
zFzZqy3yWYBU553p1DOPd/jFv5R/AdjBLXElnntfoxuNCMVZb2AvzPKDhNUGq7gb
aJl7Hj83zsufC5r6qVFEuyajd5EMlhOAHNXB2U+YMcrg+v5op+vIronOpUBdPDDz
wf66GH09H6qf1j4y6H/apyhhHjEhnsr96mpN5hM93JjONVw0ZVrHVl4LrqUjVwrq
Rr4yk8x1FK2qTH71xYOf8Khd0Q8jajhRjS6RTO3MAdEMmWdiRIAFz33S96wYnL3I
q3DAGLseaBgw5AAbW/zjVyGyAtpPV27+Q1fOR+FzRuUU9Adtuc2YYR85Q42gCmgd
rDzV2+0M+EgMzFGckUkD0HJCQOK5gvJmdAKfFv9GyT2bW1fbotDY+87I1KvLMU/D
a0NUDbgZXH2TOF1A2dKI5MaBV7M7hACGA/O2WZWQlBj0en+L7R9ykieYUB+Vnt1R
ABDaMnmz9oaaM2yGNbSBbj92h8GdGQPjE4okg7+W+BA0j3SDDDjVT5Xiis03z9N4
T0HX+3lctMOnNcNrKjVy3mPg4OJ+vRS6KlKzl6GO6Pzo+F+DE/u+FY1/mvaXCNyo
6NCTGEMAc+32Cl1iuOPj6NLrLIFd2wUjj6TPpdXRbU3qNAnT8s2TOjmtD29ekwDB
sinpc5KNTnD551fQvgOYaxZznTJRTXtQ4mrq3me/2d364DL8rbbaTDJqJDDbF32F
EqfiZb09Pr08NW8yA9nwElekeV+7zXgdi/lxaQXg+t8UCw30/quBRoTPM5cS07ju
dOaCF0qDd4yTu+arlvX6QvOAeBczO14iQ+Llddk7CjDSLz4119G10uWYcDDbpAXh
k1ZR9325rnnmPS2ANfFz1oy3Be7kTfR9yMbVz3O7h6vUya8QHPCXeezgKAAtJF8K
RzAgQr2W+jOH6nHv0ujukRi45IoFj4okn4d9hjHs89SjHNlU8sqgP2A58SkwpzSP
mdIOh9D8GW7vXdYlwoxRX5pkUG8RFqG461lthLU3IKFSVu+/kJAkcMPY2R0BNWFV
CVDcZE7gQe14j8nmV8QX4GuzFZ+bdiWoj7pCPMy8Mom72WDm5Zu4p0u6Ou4DEKLV
ZZZNG+5HTbzhEI8NhmM9EUbNrGwCxZdzaf+1YFxB8lZNomCA0RaM4ljAkS/61s02
fNgw10C1DArLhFb07kmATCiwOlZ2g5aoH+8u7tgSEzgINGO0cIOWCG6JPAqNxGAK
+mpCbD6GnMcX2m8BF8AQTVpH+94RXUDhI5XN/wTVvBFOqaPl84l85XKMevGI7JMn
WaIXi2YGEVJWmALZpsIzgqYrk11e5IsFra5bVKB78wEjlzZwgrRo6feL/Y9IiAAZ
Jm+s518ImlzrVxgWYLR1WXo/IzvdJGmv/+JELlqTdGk2bim2M0UE7kALrXGbuasT
EJ60m04BwQ0UGPLn33fO2lFzcmBzNLKkUM+s7n0bjZXZfq1TrkZmpCbIly8z6Xha
lLLrzRBO2c82R9is2Wbe2zgp+BiihcWJAkYG0mfMx5Na7ozj2SN96mL9sPU6QHGj
2B0v62KCRwoxN4POyGBI8h5vMmPPY/77ij7uARcoIlsAo4yGtg/9MnTQOA9LCWP0
E0TedHlqECGxP1Ht1nAj9OVNJNHZHnl9Cq3WvMDZFl9s6SseaZjZDR3iXO1ZmBwv
h0pnyX5vdZtyu5Q7ray4mn8qbY4v7ICQYcuSehwHpMYrmGg3sdrb+W3yxFM88Hgy
I8ECVzWCOkfqDfUvjwIHNwVFSIHT200WG5Fcooq+1jHDNgZZVjdn5CMXdLu6tIA4
5SiYAErjHJljcf9LLmHwWMSmcweQmjQT5bsOyvENIAuHuLlmTus8a1L0t/Vu2KAL
p93YDjYEN/v8xbqyW8WBXQKdjUoCnvSj9M/ITFQsnVXvSU4NBa3G9ODWtv3zLKmj
NtKbUWGIkObYGBvGcJPPxa712GUJEXfuntwRb+gYOzOFUidtSDwAayYizlq/Rcs5
+zkSssn4yHm2lXXKjbpjBPnPZu0H+EkYsh9vm5+4tKzB8u5t31Hw0gz9h3FGgl/M
W60DNIcAQhlosPu9APx+tLBgR7hgGxwSJmzmavH/dOtKVbwnvbe5VrYLG7V+zxOA
DoceIvqkAi6im5Qyw3qPmFOmLRBX4T4yoSm3kJN2IACnrTcd3LokhyQgXuPO+cdS
DglbSmbM98FFs4oAJWxRmSnhf6RjW8eSuZQvrvVPI4GX2Tcj7vWtr1kXtUcWcpQB
SPiR4LKurrBG3BgLZFK/n4b/z1vEqjUXgtSYWnfx8niPi/eq+3Jec1o1rcoZ3kku
ktGamsbQi4PJF2bu/bXXnMbWC/Mo3V8jH9WAkJUvbt+OUrw8ZC9RlM+Z+QKHl66G
b/jxgJo6ix3J9TszhQsy4jWeODiPmNw3EjwUzleFevoLOYEVgAl4qe7fo1hoX18N
+r/L5px2spgST7++VqYQOfsXdudTFuuctbqyQV5nta0rF2V3vIwPOpfT5xqOOEOR
sVdzUTqM3fYxqWjFu3ljA+ozINmhbTxY/48N0wRlNVJUBiGPkkzJpP3YMyjKE7ii
FcqqsmSHPUGFpPcjNZOKe+qkaaHVllK0lItSO8Ry2t4KMj870aSl73E20NIJ/rZs
VuWHP3mHxJTlQjwz6jYtfSJCN9qwY4V5Ebz1knPO8IuYEuEZmhm7djh5DEcSvvqF
E8nh2z3aKmYnya9pjEX3FyGixylQ5nmBUfEgDb7RFPuioXELORyi8IPOo2C3HIzh
PUUzz+vbPZxphzxsfpRSzwJtnhtGnPLRzF6cDQmZSfbn68rivQeiJC8NxM/TQ0zj
L9iTKt9+VdOXwtLDQ+6MUWbnj6I97apZ6SdHY60lonrzsGerm3V62STXM3nwCVKs
+686AVVaEQzllE0J2+HVrP8ySEfl/B6Vg0y7ZF/Ffacu9+zO90BYrJnkPrSzd1bf
BNi7SrfM00xAVP31+RrYK60s407bMeKiKtFaCB/cwRPfbSL52GK2PnbvxHPVJM8C
Jf7S9/WdVtNBfz1BemWzgJOde6AvekVaUHJBErH2T2s9ixjVP7hUeAmUh8pAQkQl
gMysKQtIvlMn/oOLD1/CFamLehERHNbnTh99pqhkaiV7qioqeNQRXtyBwvVgSZDZ
5dy56jzvpuqbjmsAoU7djbGDO6fWTSl7YxJyJhc+taY11AgYlKPYNzIgDcNKoXN7
4pmHFOAbzjvYibbd76z/nBqrdhl0J0sN/Uu1YLLQQshFHV6ifZ8l6Ucyd/AYPvxn
7/bYTPhR0lHq0+heTXh/zZYgb6hhavRFR/WXq4LZXmBHv2MgsRX9Or58JF1Ynatt
7jKSTEjwio+e5w1ojcxgh4h8poK1XNnttxn58l7OBPuzlSwN4H2wGpYGZvHk2P8y
Mm5nsV2Z1nt57SP14FaJJ8wIt/hUpTTAhK2JDXkAHrGrUCzgtX1neEv1nMQC0yjx
ruF7hDGB2oo4cKLq3L83hj5aW7Il6DmaAdmdPJJi0qEB9vnQW8uc+oT3VquGqGZh
0KjZymWccvqxfrnC+2b5XTkhqmpkY/e/gmstjtX7quoBZiUvDtaobb3q3oHCGSNj
TKHKb8c5efE4OQI1dpmt3VVI7WHHQNYr/WivO4OyZAZopg22in5Hi6ecAqitvfXi
BTp/PdttAevLmIC97PnOZpiQA0YI/jyMfX/WeYszbVWruNDpRjOg1k+oXM3UC6/A
YuKuKAIOezBmgOWDQKjdIWwSAayLqmVy8ZSKWQGiO0AavZJH9sK4Rf0neJY/tS6y
OmuZXe64V1hX3ee9IKF42Q6oUR9K7SjNepzylahAYimh8uziq0tLUqBBAGNIXHFw
TIk1GJ/pbaoyNbEz2Q7lM/t/sFork1cHuOxrYKBIcf9uxYnToFuArn41rtiZMSOQ
yyXoj4ywZlOH645tfu2NJZVNg+MzwKQ9Pn/4nUU0MvCWAJdiknTjXUOoitBlA6yX
RuIpW3wq5Db6Gqo7m6cON8ZwF+jw6buYf8kOMMT1N8E2kDeN5hG13T2k1fgGAZkQ
8aOhT2MUDsGxexzO8+gEKKaOwgJflzmxvCFtCzez52VbLItAHinqQtNbHU0k4H1L
ePyVAnxTok4vGwxuSgU/3VX7hXw+/AUAhJB0j0+RF0Idfir9Z1vIQxw0ykubw7vO
HQGkTaBWTbPZ1PnReWzEHYvQXu0j5AHykDdyCM5fejyS4gpu2Xz2KoPJ7M7EABBV
jDzXEHwvbbeIjARRCc2rQJaUgHoFm1OnTcJWfANhbgcOnS28HOwbf6uAipHRJ9cr
yUFTrBB5PITd/cLLF7qQogsU35cVDr9MIZiWNZB+XKwsGRG/HlRPbMuN8pxkGZNx
1NpGPpFx+2gB7kcTRrVETwzUhZivXpL5A9TfHwjC1ltjuPBrjWKV/ZVdnhdDa/fc
SHU6TC5BBGb+SKA4GMC9fJDvTeJR4lb8Bh/IWoXwmmscD+PHbqbo7m6viCo2YzYz
j+L8s8IFIIERnQ+jAwh8XEFk529nENIVc9my3uRAnXvsZdZNOhFQeWpuOwojN5+7
K6b15qpTeiw7khUrj6v2a1Fg6JqzKCjI+3mi8Q7Jq2Hfmp3FJh6XFTGMfnVoQhOv
+UiPPrEWA6BwEuA0MsePMxKcjWTftwbHCBoQ0zB5ua2BRzuKA+uVJxe/lvDvzi1m
5Gen9k4FEdM8eFrA3RyeDYg8t31yDP25+RSGnnaH2zcDPt5JFM4C2H+TGL32vlzu
qeo6RPbgv2sr6y4N3oSurLUFcc+pAW6IPNvhfNr+ZNDHZI35aPs4aq2Ssw1vBz8X
QGnlM6QxB6dnzhkHA4IJ31PMASlLgX/biAZ81qSaW4u7WQwZ4xII4sLHQIx8hWxY
GWMrdALe3iaLMp1DJCNVrlz6m/t04Zxk06uvcYThzK4UGPS2SA6YCJu1OzxX6Z32
g2IOURtmP1i7G5FWUI03wjdrJyOWFVBdDD9El0lHOsjhpAM4bk5zTN0r2ee6CLAy
LsZ10OgLycE4+/muA4h8bKVV2vBtU9EBnwVLuUkg2Y+S+0W18y9g6kNaLauVL0kH
NSTIW7ZkLobkuQr0ZwB+597Ez0zRvth7UAdCexUoYyZGjjGPCufW4ksKMMFlECTm
5MIrfIOAwTK+rEVuCcnxyCu+ltGrZ9496L4xJEcl3+yuPERPuwb+NvIBc438+Jo4
NxNvt8/snMVshhVPQYCtbL6kjHWiiKnRZvfU0l04BqD1vmUY3PZklTqvzOIoRoxb
cd7VfjYTNEJqOt5h62gRVB4I9nLe2lAjccOuJ7rj/b8p3cDU3g0w3ZjUmwkPYizE
03FyJp1X9Fp3xK1CfVeRtw6X0pYFGRQ0dU16XOvJ1klV2BjFfFB4ivocOuO8qqZ1
LjcTgI9VzUwuLE8mFMzQ3K5L8so2s9cLNUjwiAuzvHPe24jEZSm5J7reWHry140y
LMWIh1+q1kXhWkRR/MNcwp3JwJG+k0R95kBCcsSji3D/Nxx/s88xYJ5mAUxKuOmz
q949souziXF6JyX5YTmNfsXhJRSlWGlV2ktS98WwPxtIf2P7GuLkuvZvv7mE3qkx
cQOBGu/Nu4Q/+ZSK8pt6YeK2uZKWgD+Eh0pIzmq8pwNjXcNz6chnzMu9Go7j1y1B
MWiFs/DM2P3e3we70BfmmhtPs+zDXchnSw8zq8sR2GmeQ/1hlfQF/OyxIQED+1qF
tCaMeXzGByOsCH6/daLl6Z1JH+JWEu5YPQ9qTxVbEAvmoobyBxEawkf/DsBTkagq
/NeUcgTMjPJWSjuQ+0lDF4XjajAqtC9yX6k2CaKDdSN7jUhdRhHoGpH71AIy7E9O
2xQhvtj/dGjQuaNTAX3hOgAg8NVZmjKGtZt+1/zHT9WVJH1ck8SCv+983uXYKo0d
k4tlhlmdAcKxc8+RoooFpNLx+81GJpw+mSFGePSGc3UxLRfvuqgI3HTEygkWgXZc
jINbT4u33OmF2YH7rfl493NPKl41EbZ4eIvJcxc1v+cjOuV1ECcOWzZUQJOt6tH/
OP8a8Lie2orOYo7tG2pr1NHCNbvsT/LsgWia8LQCxuBXvsANTCbaJKihIcU0aYiz
IJxzE6RAeOfDtZvZD4nUdkyq7qX53FWG9N63rZ63+w09lH0JOlRi1AkAhB5hqFiY
rQw8Cwx7pT/qOqNMJt/w9/I9jgxNVeI7Ebsri7BQUR919uDoReWTqgI34mtb4fof
EN5Z+F8f3E0lyQalddDGQuYoTvVCfn5Glz7W6kSvAo0RijKVT0tGSKrXN2mWJmkq
/hRoeFOwbMkdMw8bdjHwmGUeYeNlUPhSFcKry5relzLHoqZWsRXs0sCPQBXNqbZI
dBEykUs5Z5360mmf+mqted3D/jxNZoWY3OTzH6eqS4UAV1jbrGUwFkR2LKeVEMgm
/VnZXNyeE3V9QHJ5RlmKye61+yp6qHpcWUoVQyQxXdJsgRiNjSbZ+lmbqG5nXj3K
kI8zYxTO/zPPwZ+34LVl0nrndLAn3VG0IOASiiHzVxyHR+8Wj2OBWYaEAyY2YZpf
5s8JCYAvMk77lYbpmg+h9MvzWeKUIkX7Z0A1W+MMlzidlCem5mSSgVawr1SBurTr
Ygje3rKK3+mCsEA1KaCrvg8BCbuMV1iGWBlHctxuhToyjQDQfnGIrwR0tDTPPMSh
5SfZ+L36wWNe3yp3xTJM6hWMWl6sGRgqVZA5KaGy2H8ogRz3QUJ29HshVFSyWjfe
p5vbxS0fW4b8LEh8IkhsDWuoOF2xIwri8rPILoU+tnXnD4FARzG9AhJ7otSI4coQ
YsJzpFiOrVzArcJF/bB9/s8DT4dLMEcNeLzdD6hKAmARg267JS+vYOw6J8Z3SGQ9
lLAwZ+9EQdgFD9iuzE+szavHfFDVAymlYfI/Zyq5n8EODxVUBw2qMGvEkoe66j1j
tODISrvwHwjhpq093Q8nV+qtRL2Hmo16jiTRMWubzQBSaf4jqAtow6x5AQM1Zy38
SWowC35/Ci1aSfWXQd1GzfHSqbAI3Ox3wEcAH4liyuShvZiCDGN8P7aAZSETrR7d
7ih0hH7D9+hoSEJmg/om+e+o42IW0G1uavQDxQZiB2uCLPnMfNX9crF1VzkGYTnO
zADR0aawyNpYCSNEHKNIMfxIEtttO4ZTnO4Q/GgRxHtYxXqJC19hy0AWnOfbfzzF
/mDz/JSd6c39Zy9MxVHPT2KG3V1S5FqTykcyEo1qlN9S1qmXbGu8QUuJN2EBU0TH
3TvmjQ7cxAuX9wzIabH3j2z3h2hDW24vP+27e4LNMtuzdCsZFiFiTiFZDWCyuy43
UM4q8KZ85pNkmLNPsnYpmxzbNFNkJ4XqiviasbBMImWiSKpiLaWxH1af3tPOoW5i
FjjqWBXKRU+1IzT93CA9NEGVDAgHAFqzRO9AHySSnhIjIfOT4nSd2EpoRDbVZLDf
sP7exKimuOrSGhRKnbc042qCkGy6hyOJgnS0xLcK23l6Mnn6rcGYn81JiCk0V8ZR
kHcA5d1ZnW6Gs81cpSKOeuM4ZEcOU5dUFAy+jklBIsgF+fq3h8ohbefuz7+iJa4m
NgKd9QOyJoiUy+FTRIavF8Yq6QMfrDZS+qVnDYTQuomec6xjRnIw1lU+pALcQMdF
ezUbUYrslecOi0mI0XAwX3b8kKs4r5JAhfzXTrwQcpIbnozLgKjk9aqIF5kBHYef
oFlLSOMFkPeACS3THvBQz8ifbvSRx6rJNgAs785pfkckRt/3BwUEkSaeO/73YvW1
egRkO17eULV78Qqz9XHI8elIETi4Hl0INaHbmEiTUaj1szrYExltvTV2lEb1J+If
9N10a0Tj85C5ev9/jrXPOWjrNINFBCAwnOfPL5bbnlQqD83Gvbj7a3Sdmr68X5Hs
8zdJTWaGC+WfbvEoOWkWfLkpx89mI0jFtc5WSWuiyF/Nwb2vSiJJdXDLetP348oU
XrTcSj1Et9F6DP/InhI4CRCXrum7po19Dx9wi8mPZlXqFCftciFjUJXPfU1/QEyT
qqRg70nGnzyy5sPYycZ5pg3ZnTwNGdELDNuM7ZGau8ItGQBdRrldTheomQJNmOle
ZTwamBq52/2AOXq/sfgLYwWOySVSr7URYgXKEVWOKPVW26shrt12HxXlxkHOEIy+
a8takha5mxDJqkKLNQcuD3H44MFh2s8+6Qe7u4KG9TDu9LCjOH5O3IqU+3v/6Yn3
envvrvO1VxPcrUzJqwRjAKwppPbxX+XUq1+9D/SLqrWfqDmKPUqcBDB5GT5IdFRN
APepMqXcaL/jQUJ3KaC9pvfu2xAysJ9nqw543eNBv9UNyZwlGzByMatWOunXgYRI
rivuBotj2h6jGr68aWuw65liueSiZD1udY3mynBIqWh+7gjIlwk6vQBZelVopaO5
WoWOo0Lrufba0zpFlg0soSgcJncZFhplKyQzsgH9VMiUnQbUj1TYJLpUtDymxMG3
hC6oi0hS97LZblIETY6a6EBB7/u19IyTjf51VHIVU+PrJoQTvaFztVT3Cioder4Z
wOTl/IR9YcTOW+U4xpROggKwuyC2/2ZaSqHkr3bWNBsGPw0nBDksbLSry3YUXUzR
/HSeGYRsSa3GALGcALmHbfB6DhxaONmStzIX/4KnpKY5WD7QMOfyZfPa78flIGvp
UVZOmHVU4vyCSb7Ya/sYmeG6VMm9vyrR89hB8d7ooqNQ2mdIH0gyHc7ES6O6t+cx
vPz9soLHYWtPDzZemd3D/RUPhxvUdkE8ZU/LLCwqRZE9veQSfGpCdZGHhCpgooDu
1qmre8AThyPPN5u3B/eFaUfG2jgEwwBkGpGClwQfraG7/HXFxRi8nnYdxS5LnGxn
k2Ks2Z5Js1IHIyrhuy62VngkE8KaUTrPJj7lrsCaEjFByc8vHnb2a6guyxUTwH1K
S28e0af+Vd8bQSt2PDVUpTZME5OtW6ej0bOMVruoV5OXwoRqiGpP/p/N8FHMKbZT
Ji1BaeJAoDNCIr0G9nUV+NKDvTS+nfTlPHII+cwDpztJS2j9ngdIo03VfMwDOsIb
ucAXw3lmmD3wwKRajzNPNhFMVC71rAb7xm6nSgdJsOrqTVFNlgcPID39EzAAjGI7
YZmKObwSr5BjLwMdytur6c71axMGyuOCkzugHP/+IC/no1zcXR8L56SgsxwYdDX9
lLYwWCXOMvCX6CVfFHC3LeOvmzIQGK3LxyiDxFfTmarVGXcFFuLMDUqMTEis0HvG
CMuxw32n9WccrlU5bJP77a7ZHdyIodkOME8R6vLrj+qU8DZjLij4Sg0R80PdK19q
Doy/BLZMQfoPGF8HFN7IngI/QQsrFW1wORQwwdZLw70NnSoV6e1WXIgd5TXvyc1H
XGBu1WKQxxPNOzCUimZRim9n9NkC3A6UCBoIGs+PRTt8rRJbktCae8gMzyuCVfEt
/WVGoj3z1VedRAqRb25ohYPycjTPeRYhKKfNKWXkcMo1XAGrfmgH4fun0iLJWBW0
g+95C6PhQjn2ZmWyK+Fs1S8auc84+KTPV4vzWiMrvIdVNygEu0+ex2F/nnDrdYBO
BBzw8O/MlgPL/6NARf3kaLZsjrVSqQ0FaiUz5B/jv/9sj81u8bk5Z1bMejConaXh
h9bHnkgQRzcTouf8VFJHRx1dOZYHextl5/Ez7iAbst9z1FBnpmzRNudlD4KjZMHR
aRhRX9cEsVXvAoC6hjpcGGh3MUm6voa9kIav81joec6IMT2ruAinWpkewiWbCdym
KLhvi8vczVGLoOtsCmYRJtZZV161koZZ6wDZQPmndF8Fn3PERNuxGRSBABiUsHn0
7c+qisqzYKS4zAjbr8wf21Yrsm2xF+OdMhm+k8Y7oRPVpJRVimy71YARiY3pFsO9
deRzHGTyD2E+VDA7ahzUpmdF9W0vt7Bn6VWSpyFUbnnBjuqNBGGT6DS14gOsNtxF
t3eLh0QZwsbwRBkz3alPJwtp8jaZObFo+1jsbOpumGl6CIYIExBib1zCEryxPDTt
v82HiqasWHaxXB3ApTTpWywiVaj1X+ppAfJ0TYmlYq6pahPDUcdBbTSCz/7gZ3NR
0P549aW1SXl5ok6rXJ4VqJpHvIliW2yaZCnuebC2S4Efau5N4xKGYsUS8RR2HwTQ
nCMrsHmlURXfWFuECJH4bP+sMo+mSe+2Ub+NvzPCVHyJi+Pdx29ZABiHZ7LDB2sx
9vC9ju1mSoB0L50abB9b+lKO8X42NARo6CP90XxjAOnXdDb/heFFc4eDWGLNmQ2h
tS4AX3FF5ToQ34J4WCRCzeYksf2govBQwYVbcpCD5IJqDk0rtjAR1mNhGbOMyNKA
eRA0tR5idby2gAG1KqkCtivudpn1BSoo3KZgd8860hdlMajtxtqYynTdNDwwZtvW
/n36CUzCXAJ1WFs4GNJcNqIvwmhti2x5O6Uiartp4TUkB8brJP5+rJmuCz14DYpQ
n6k0zBRA2k+NcMT+uORJRITTMqSFcqFXit9/2hlAuECb74+uWfGgXuLUwkAraThZ
lmyvnOIDtD0Ec0iTkAuS7oP0Yd9kXoj09fFrZQTmKCb6v3jzHURR2soQ+APxHthd
9rBKeSMSd70rSXY1a0a4cpKAW+Y4cGdLI5FFkObcbjczPHGn5MXIuC/3oNL1Xv9b
LzCd1iQtdABxoz20Wqox9zkMUjr40RkWIrYLfC60WrvNX4G/5Gwmtmm8gdg7TeDH
Ks9X5fBAQfel95+usMbNasREv+pFu8awAahEtd2FSEWqxSL3ZBa4Il4eJiT1iYoE
cm1O+kZ35urYAM4v0j4gAHM2rBqNICCXPtCFbTNdv/ffhj6HdfZXZHD0GY+dhsVw
2oSAYFAFWIZ1ZjHUVItB6lIuf1giSz+5oJDrTnVq7u6j8Ftd5J/JgU7Wms9OTQhr
nMytvdlpV09lqMM4kt9HFXEAKmJhX4UCLvTkxyi3k8hTFAgpU97jOnG0Ah67HIaI
H3yF+55n49Z3p4T5oQDKnlKj8WRVwElJzvvZroXL7/TocRJG1XWOj5ox2t8bHS4k
Zu4lIoYKIqlUcH5GhkgLCN2WhpSqGwvAOVt+BnMQIKrN49ggZKasddywKjzabbvs
EFmysG+/q49zGLa1R/zWnX9SIQ+ox0MbRrMhSaHZvgY1dWQnqrclUjw51ek+pTql
pZJbZ2TyZRzHG91s8seLe7io9tVzoGEBsXBlBgV+PTTzc8Qap1c1IRABNsCH4mq7
u1ZmduZRWlEs0QnOXYuoxbULc87w5U44x19aBT0Zp3wJUEVxeUImNWB78O7hxZOk
kKwhGXnAcaytJ29c136xGHMSGqfXMjpvM77O3I46YpLM52kfrv9rtLD16UDkgmDi
SAJKN8+R7BxzmAxQpqsnH02nR9FNAXxupxwVvmcNTnk9ZslDN724N+w9sRmnL3/z
luILPif3XEzx3IW14V6R9pFSa51M5rlJ0+uuL7b46WWq/OlUeWJ92fQ2v/LW+d02
5FttGg67pIzE8POwBN2Wfiz1YomLwLS3eO2+ljoqYHhE5UjarcyxYA26k4GzTY1w
o1UAXDjXWTejQFu1GJO8w4emZjJOz7E2S1QAVuuF/344crn6KOKVW3vXV1iMBlQX
ixBIzYHa6cLR9gYALlwe5EFUkm98CELVDf3a/TLSY+rQkTBTw7hhqXfoFor6QNtK
Il7DWdBUp6va2pLZOCix7F1UhrZFKmZmDi+lDGqwcIqK48kZmWAoIZD+Lba6x6pE
5MtjZyfUuro5uN4QylVtn56inFLNQR6H+Ljm/nF/tCC0c4cOAq6fOM813w0Y87+j
bKQzrZwI7wF8QPYJ7/qh3WSh14o27ZbjmMKY0aNrboJBkhJlswKpJARoaFx9QJCK
NgzAlt1p7bX2NU2CFHAsJ6YxdlG7ylaK/FK0iEfFMdi2bUAf6yfVdob7RcfrRXiF
0FOYuGW5uUEK8kuxA+daT5Mkg9++zyGeuEk7JjC10Wr2W+69u9S45ag1UmC7iJ5K
h07nH7HwxxA2UNhxV3wDT+ly2NPvTcD6wpiNeojiA+o4RuSDuNqXXZq5eiy6y5IR
Aku+Sft5z90Z/0Pp+fqEakFJF0gsz15Km7k6ZZLeiwiGAkKnP/4Xp8OJlkfbX+7e
n/jZRX1wK3foXV205/+mCKiGI4ubSksoOWnXDk6axXhE+Hvuo0Vu7EYtNgg/oRfY
yq8MSBdoBSZD+UQbeVNdK85Xna1GHxRWuOzQzmwUabAGa596LBIVivpcHiObWvGt
cJA153sCzV/WgQ1Df2HpJ0xOBILqRhh/T1sgc2f5yj0sPgKVG+PxxfHoL6RqmYwU
TwZgo1m4fHIPH3jOTDD1120S0ylckNU0VYb3YWC8nl0lyXlt2quXYIudIGiopr7e
QLXe6HYLDH3nSB7ej7Ajjlit5f82dnsk1HxTYVLc7PFdgDMl+k2/vVoB2q9yEPAt
ZKZZ2hUNUMLEyjid1QldNF3KO2FmaY+AcyBB2Qit0dX/NFz2T8KcEoECbGn9x1t2
RP0pU03k5yeVqKBzF1+d2CuLrnyzDM8KiVPF3W+XNcneqXlMe9RrNq8sPrTO4gx2
l5Ku46guWFpLALb+yvb9r+jW6QAnvZoWL06b6eHKnpRHVxRgCXXO2bHaP97iFT+v
6KFwWIBlGc2Ae45qHJnYqvq3OXfjZZTVsoXrzBQMgZxaJxUVaAuZTj8AE70ivEbK
wiXRKYQo6y/J7idexcBpyNMxksTUJ0ctIOqol/SHim/WuN6mDOOt5sWn/eG0s3/R
pQAGi6Mrtk8Jc8bjv2CYpIHRFdVBNmwUY9VjblSQBq29ieYUW74WFLh+RWgnwu8n
c7rwXQl/JevpUjewdp1qiHLB/wmyhQkU14hHEetrSNGEpfxtsGOnX4hFGbB50Wcf
qmgbl0ucE9AsqtqScU9h45BpJ9GwbfgzPOjFZ0659jGV8pd2fWCSSKwSK0nBC57k
1Vlbo3i9/pyGEpG4XhvdN6nrkIVCdW2LK1VLoxUfFvpAuaU9VoJ1Zs3DKqtCjprd
M7oYJNe57M5I2qb273Ga/F0jS5PRUylMKJYnyUQxLFsvwQn1n59ZBXOYh3FKBej5
0Elks35kDGUZbFra7AQO+hPOvcJDz4PYYb5PDP3fmbJPytVg3SHjjbO0JzyZ0rXh
CHpUrIxoac8OA77me9Fm9NBoy03or57L8sCn0AKTFVUMdtGPZSqbLafdBhAcX5AU
GToDoT0Y/Sk122m+49yU4/IPgVJhKswunJBfA5oysy294AHocaMnyb7GVqbB8xlW
2qiOx++W4LgkDvlOLK0mSpYH3PplvX8puXphd2lozsegVK55caOgJ+2oYcN31+Vx
tnVrxzK81UskqIahZ0cFc7Y1jL7tExezfSDpx40HggeR+Sp+watLZpB/M5wbkzfV
S878A8494g/eFXp8JjbXsczoy0whTsRpFcK57zdC70An6d2KCo9Q8OHklqPmjM9z
8EgzIdGugMlQN3WovKSuSX8IlxOYUTsLXp9Tk0CTu0BSmH+2JHcPdvS+kYBr+uJZ
T5o7/Ug3oon9UbpQnBtX3GRn28LFEWt52E3dS+TlVqQlXrGbdCAFIXDtx8ObAWZW
CrMUj0scBIcVLEudSqEe6YrWprUA1XNRKo6FrSCzQv4ds2SDRIotcNNmDVwze7sO
U/io4aio6zoHtE7kTdLgjEnVLUsNBsqkLTg7WcPbR4eI3ql0fVyh9qNPSZUItali
HoWmgwXiHb/zIbLtdxswxGpNSBdY004/l+nt+w6giyEi5bLx+Nr5GEUtUlSZONpx
5N6uWe8p20jDgW+kWedqyN09f3YPAAIkAnQkw/BCNw/kVUW1RRcOwfnmVtBEhd2S
cItvoCNtJv8wmyaHUBvIBo1F/ftmoDipSEdH6p0LfF/y1pASLXUN9lAaP/5pRNdY
e+EK61sFXf0COBF90Qf1YpQXMcnNp3CbHeFR23oHp52HB9r/Yv2jv7lzY18VPe6f
GIHXXYfJAcqXTCt2ft3cGAGOyXe3dcFNb1I/DMRrvLvssmpZMHNJTqDbalBDRR88
RwXYgPsDvLhco1J+W5PDNR52Cn0UAGOqnao2KkDse8yVXOQ8bnf2hVhwI5FhQkMT
bd7HxzGitaVxQBNSCZKO+dXrqiuc/T0r2E4Wr72UlnoL4pRc2YsnY9mfkYNmoXcc
8vaCNzPDCQNuGbT7V2gfLCRvo17kwDcs1x2bSaqEZHpjmpPM66VKWIcDNR7Vb1K1
Bg+QWLJia5PZNadm1uXyEoU9/j6M+1d+NbHUUFtXP9ug2ktP+Yiy3H0WU3dWDcYJ
HtJzaRoKn2lhVnFV2xLaLPvrHAH8cSfKsumMxt0q3zVH+cJ00CpASTL3c3dPaChg
Iq5qlFFlOeOdbK+QJ0PoB6PmallGV5yiAXSJPZL4DyHBiej/dN0rk4BYh8g0475R
oQ+dVeo5s6peD1MSphcD3XxPT+NcJXWyvoKpzDZiF2Lf6b1ApMqhlBVsjf+vWiug
+sSs1Csk1PSEhLkWdqejZnFk+ytj1K6+fYqweujrqAdIdhZIaEL0FbNPIFoRpTNA
WlIJfX7tY11wIcjZhRr2LcdbflfPQbS686Y+pfoH6qD0+RYGIVFdDcZiuPPo4Gux
QwhGgG3xEoViBxziHZA6uG17DS5hzSzPslcFIho0gfGqlxa4Fyfq7REem5V3v8VQ
/QVNJJHtHIBGw9nclkNNuMZJEW6bYEuqSDJM8i5SCMwT8DOHj3uTTE4V3lGxQTbK
Hv6HWHs6YZRMKmgglUW5MrrS9p7Xodph2O5QqzH+xXLIQAp8gVHObLL+DP8rvv4I
U4YFlZYeC/CO0F6y3yOBaDtS9xCi+Qsm0M9XeqIXW98lVUDYerepzm1nqjIz8XEK
VtfRrvskWcSJv1kZZBc3G3id1P0m6FBUkvgWvBXzK5j8SQCDvy0DqPvUmwx4+UJH
6EcDGwfzgId27H9KW1L9+x71iWT48rhGsLkP3kzh21K1tqohGZEPfXfPDEdrVbDk
f3KCCH3bxv0bsZCq3rEDEu48UTBfmxI7AGSh3e2HCnvGpOmogT2qp/7QNdQW93tS
lRx7uYkrIGqeWPM1JtnNYPkfutRbW5VW5hKnmaBFWKffYuYZu2nK7K4/sOvP5O+B
kD2FiCpPHWzJ1Fw5oDFhM3wq3qCJAW/gG2FU/oltpwmIV9yiwAKMaKruNuKT6F/C
8lKW1iRHsIuMK2FaAYfXV2TxD7M5bY1N95P4w2QT2C88l6JVm1Ci/XhKfq76dfdg
kziIjqMFCqw4arj2bUPnuE3oO4DwEm5KTAxcXxalLWFQEjSciTRRUEMA2v3mTRAZ
Y7z0E9o3CONZd0vpOVE8LNg4O5mu0lmrN9p+WU3bcdbE6DBHvmMw+N5aUDf2khrd
o3SDVdd7IXCAV6RXFyI1hFbOQ9DXJhRJDEqEF9Bdg4wPNjgKGgd4S2iaYKyd17Yk
sUsFNawh3sjPHJPDrItoDai5w0z2CYkqtbisdLD5OJdgylVLB9S2zW1ayXidqlB3
fqNIOkCa4taIM5e4YtO2mxuJM7NxLoNWwqCq5xp1Y30Vzy7UrJ6p+41gVEcoL8H3
uhQsWRVmNxFiAnjNT6PvAQ8DhdZ2XIYoh3I7jsHpag2KIJNXzDT+/YcPke+dWenl
a1eugcldKskW2rg5ThSAcJnQYLNKGWigjezkZxgB9drB/17w8VXxBhiJDp+i5dWs
CfwafLY93WhBLSHrLcMnscwgez74KNDjKae9bUKVI1fkWyt/PTrjGbCEdK+/dUBA
j4oLcFD6+uLrE5ZbhTIUS2djeh9wbUwxEd0B2H71tJnVhmxIzMT1dPOxoEkttnQW
8tY6DXPOIoRjmOYfNpybPLLDDwlDDZzkDDFLidUNddPx/0aWXbWPRcPr1M7F6XT6
9L/27DFSCA2u3rRnr7raGSiFRVjn8fLouR8q49LB1M2bbp7ldMG2bP1uQfGnvBft
ijKMZMatvzjhGXGsZFZe+OEyEMc7VA9QreckfX4kyfZkskpb4Zb3JuFNamlcSvo6
mtzX8Pg31OEvStRhZ/jsPDl1zt19aW8qhaTna+SXiJwoiFDPHYQiFpxfuZb3ZRK/
TjIhLqw7Sw86aQBIwhhc6wtXqHNW1OHAymxGEqF5/+2Ar+Y/RCKNn1Ph694JXcDd
smrDz4fn9Mvdhcs1APvKiUkZCB6aUW+cx46KZf03xf02WnLtfhokiwhkhDxQpRnr
TM/Ocjaw8+NtTbq23s1+gHroTbZl0y0sXnNVkMnkKZ337img7rOtfCmgBf9wLgJ7
lDDgEc8WjGriSTkjY3eYHaW0NtH1Gwe8MevrqIz8E2rAR2bMlZoydzpM9nc7HgDE
Ry9F2XbcTU93PNGE/1RpLOAIEVc8pXgkiMNxJQ1tMQxvDBLLVDmnMPPj/14sL+XL
PRQfvXSo7DIq5LvHfAYuWJtKAWu/XXC3PH4hgpHKMrfuHGzDrIgF/z10jqK+3MCw
diDo65wcknSwAl9qEIKasDUZ8WN/OzmDbuoNAYDq1Ni8w+WwFWFsqiC2tbRgnQkV
SOOa1Lzncoc9+eT1YjvtUDfdRPloC6YWhPOAkLKvAGKJlKXcT1NF5Ay8K6o3Npqr
KedRWIZIJPsOFChbVBeKbHn5WUn+B8pJZldB4/e34anj8/2/JpYGA028JLby/ILM
Zi4CnafGJmeBnJFxqA+RVu1jHecJ3JHMXWwIabPIHJnFTwitX1jrZbvBKYbe31P8
IdJe95VOYu4Trn0Mm6P8hylaHvLWlG7mnQTlTa6VmlF6y2Vvus9DVXcLkAZ+BpMj
9hEv/xOS6RMQ9BrIIhnP73/giPssEu0RbSy3eM1Dnb+g6IC9VOnPG2bDqQUTsqcv
Zo57HPghO/kGNdimT3x52KeksalovL/PvDHuxm4sQVxjD0pSwV6Xc2+JG8qzdSy6
o6j0YPAmo+ct7k52JRkxhSaZ+5MhOfaRq/CF0Kz7zfC3vKGbkuBugIz5IQtqfymI
o/RfzegaFOkL2MIckPT855mw+M7yLyDmnU26vYMLs/ogwHGx4/xP0rmw5F/1HJiN
KEFApg8CL3EKIDTzJaEDTO4afQBzDGkgXFZJK0L7VJeOI0mM/oyii24akV33T/Ur
5iCkEQvYKTGs99BVo1BeX/3BrwnTk+FYy1U9m2doY42n6UsgeZz9yekPUFoqLwe5
skyrlcJ7UrhdClZdUgPRDQbjoJK7u4mK3haeJFtHUisv3fd4DYGYOweVu+XZ1MzL
Mow4dtQSRT9jRy7jfjAR1h7mokYOHxfyNC9wmueA65wjSkFIWawGC1XlwKFzIfIC
myVLpCvvE7d4R+7bCWRKicb8gOsQPCeGZcjTVMmvfyS6EZQZD35kYT09O2HOkQgk
RwcY3aiz8E2G+JgfxhmoKnPLInCjfZu25I85jDgCjnSGVr1TIS8mserhpeX+KCdt
gGzD0cfWFf1Ir/VHTgiJZQyA67ltIXkRrrFuiz7vaGKGyP+cM4QNFGzP5o5ZZP2R
TbIfjjB22rsYKuQl52Luplak0Jb8i7yMi0uHe6kh1o2PpGuBXVrg8DB6t9aHnJae
pABlcktSDegFaA3XzD2STrZiv7QNqNJ/x27GFbapCZgArkjlvzDs0RGNvpCVNq8i
EEEt4h1UUanNKeLAkk5XS3mgFf0FRDu/loMFktJcC+cFE1H+mcYToGC2l9s9K6CX
RiSFlpHu7NQemcQ1rgxCXx5Qo4D+cJX3j7ru68oDMsPLbvcOzLH9XDDOFDPHAED1
vKlqT3WtFx4Oz7hn14gKIypEnVJtSlPrZ1KLCC8EqMMPyrsJEHumAajvZoUIaSE1
xMMdR6oWI6N6DJ+xdNxa6Ho9QDusLOhb/1qrx8katqJTn7Bl61k87Y5jOcjndUj/
Gy4tWdduFseVDOTpCO9dtFuC5kurdET+j9/mR8XZhQeLcxsU6WS9Os1nZm7TIIp0
/YEMFVOfNuNRtSdkQJRgUUGplpCXyRtGojkOushH3HRb9N5g+0I9mA+MxmWMlp8Z
RRgErVHOJtMuN65IQQ/Lq29LDxNEmUb2Dz4QMidjaP1ieHpNVjhfRWNnZRJ9A50g
RIsTsh10zFlhs3vtDQQ5ot54RMuZvrRCo/Tejp6ee0aN3exszb6HE36ClV6E9coe
zBt79mYh9819/fxNe//f32IkyV0xqTXgMx4ZZ0FlazwAvXMk8OQUT8l9t3cx+ZYl
CpfEolWZiZrVfe3ME3Gnkseeb23BuGj+kF+KRJnz5FVHqmvf9s9CBodkeRKzjzQd
q8vH2wZILP6QFedE065R2yDDS9c7T9gaTj/RRSq1lMhu4gEiPYHgorL0h2xxYNd7
mW9RLtamzXi0dF+d+iLwNaVnOMeCAr7ai4wU7oz1JoMyKqeqZdB7W71SPWvq44Z9
h+oIXLNqu3NHDSo5/3yKelFzQWu+13z8OK2O7V1+muPLxV2ckJGBldw7bbZpwRky
SjR86NU0CVn9EXWSDw2lOxfGh9GM5w44X1vf4hHh98N6ioBUewDUwA+NrwW1xSTl
rxYY02XwueruWJUG+hkDoOKZPKb19pc6PT5yQnt1QS3xli1KoNiLEtxUXuTo8RIe
KfsZjmh9Rsc28ZsvhkkeIBkoMDHPcoikUNyaTvFVZNZpx1CJ0zcxcmGiDdz3DuvU
0mMCcKgFSsv8riD1NvN4vtiD9ljdmbW42ClC9v8Bf/S9WLuv7IAkGG27hZa9L1VA
l94kvho1GdWjj0Wjxk7yW0k7uCZSo0V+GLoUn/PNAqIbKcCuLwMl05uyukyzFSiY
JWDcWHH10eSebnkaLGbNIjO0i61Jp02IAXvUz553KNxwIW776vZLd0LubnnOniBU
pG8BT2K2apxgwmzOdhvJfZp8iSF6Cy+vWpkf6Wexyn32Xt6+vdm7p10nq5aQJV/O
JSlnu5wK2fbNL6YnosTT7Jrz4C/i2zh0nHko98Y6z7Pa0yZ1YqwYWKwK6IZjn6yi
+JfuwVlNfgeXXx+5oYzoP0PheRWTHLr4DpUb9bijjnxMo+qh5hyyFT9VnymuU9je
j92tMemHghwNM+pOab/DxrRcQvJY8wc146taz+9sfUyZ8q11dMrh/W0PU7Jh5brr
n1bfNdL+zVac1NtvaJKhC5QNQmYWu9sx62Frttnpcdic8a6GuTWaLzAdVhqrWEcR
m4tbYYT8sOfsnVOe82RQjX5A0amlZ9tWwN4aopZYYG3zlr6zdBUQ4abuF+QQAhxT
SvArZ/aznRPR1jBM08F2IfAqHGUFIKvviSjpSgFN1asPcw126BFPtxPaO3qDbsOv
VRnDmvUKOQ6O0ftJOdDNI8HDIfXYq8WuSBTyTcftKBH69eSCUhmEXMzOMu+IMTox
STSS4lLm6BoS5D3MVuv7h5jfNIV6vodw/upF3YCy5AWLcgoPmRt8p9mZKuMRmoZA
+WAUOgF9LXAX5+TSNpSqM/kAq1W9Y94OLFT/jqB07fNucxZjGU7Vx5VCXPXRij/Q
5dHpGGG/rPP2AA0wuN7KIOTuy8nOdB24nPclKVUxfOGfoSTtLrRFsMUIurKTDiGI
/vGEDe4+U/uijDTvNF+oEoQmA1j02Kn44SXyaqkQ+tT2qBgH6qyn3IdDdhFJBqcq
0+scLuKQnpldk15RZ+j+AyC4XswSQzA8uY5+tH34M3IqtE4SooNvKc0R3j7vGcQ3
HiFWk+E7lTCRZBtmpVwrBN70xsKQX6YSX281L007tCgA45RDxzD1dwolXc8KU0Yo
WV81mipP7RhTPUp5DZfoc/xPrzTdTzL4bxUipBYTjzDliT4sPytxlOGCDzGybFaZ
+a2ilHnT7wxtWlBiD0HPvk0DZmhjUzks7jMIXiIkWF8WhkzH4SSnRfhr5Sjd/Sr4
89bsqVPR/f6fOEYyWu2MAuqe1G4VDHnoCG6qdUlVhy1brYc9tnQpkHNpl0b2IR44
Pgp6BI8SsObnTp8A+w6oU9ubBhqWgKJg0ulkbXJWJjyA+Sh1W7ScUQH1mCNdKHC+
ZTFhQRp2KzvdNkd6PwvwKERoZh0SqvA3rO7Fxj3bK4fifVAnkG/T/H5AKH9/aL3V
x2ZxbmKW9S5tUs1/H9L1nT9YRyR2yY6Gm4uUHXF3tD9gRHqdfHUFH2shHRd3QhUF
X93K+dANjRTr+f60avlR5uICK3Bbp4eahp6o6YfDrbiR8g/EqUQQFK+/YPFvR9hR
ibPcHTw7QnQpIEmhmJ0qLGY1uCreeszoN2+GK1b4HB3lj4KkX2G0UuI0F+4jLPhL
SqKLdrDG/hrwjdaCcU+Po1aeN9W5f/CEzPyy4FurmBzzfABTMhMhT7aptmTM9+od
i7NCHFSF64jxQ6lGBueVo1LLhb4um7JwsaccbrDo7ysGinSdjNaxxejrV7f/kyuo
rYlWCEvmqstarmi58nSf82AUeQnP5a3lHS8CUt8wwxZ7PqTfmLjVJPjZ6cgC6a+p
RROtGlX037pt16iHVhdfooprVjkSBE9vg/XyFkRPLwUHDzR4F+QrQXUu5kLo302V
ABbyVKa0pPfZRGn8AnAx/8msI3rgN+din9RkQGtKY5vt/mxzoQb2ie1EESexUU0l
N9MairqDF/I6tLAOUHVpEioA4O9qAwzMbD/VXrYlz9Y2Bk7gmOToWDetoxqkBUXZ
pkUudXG2m9JbhwfBJJo9GCFhL97Bx6M1sS6dO88ujmBTdlqnT17fNboWXQWiK7ki
mveWAWW/1gUtJwY3FeKfOYV4CTAd3i/dG06uWi7qjdwvxW9vETb7/NWQSDLUQpmU
twGygHurfQYUceDZJ4FfRrCCnd54+Gsp0qrSRqET6MS1P7F0a2BCymwZnfkusQB9
dCsYR8iWe0JkFj87kcy/Ok9zu7XTeUjd/pZFKNBEqeuW6SZdd+/FDG+wN2e9yACC
xtzZHB/pwkDjehKaUTz5AXbY5nMWHADhRODuQfItMPXntL7h8dmkUWBihfvWkV0T
+zWRFQhoN2kI3FAcCs3OdtUTHxUR6wW/RH0OIOgxjJfKX0ywtAjpBI3s5EBoTfRc
422cMey9Y5p5gn9BKSIMjy9HzVWmS5CPyGCmFHKPgSDZgybgPjktx2WCb3D8kMgG
dprHOs+J4DMKdwaeSiw+TetE0sIyuCb33c/UAxiO0gdmqPf0Ul21b71MekkhYfwo
tOVFPpGPgIAHBsrCEufe7je9nLN+teKN72Jfh93Nlw3gsvVbQG/6rqRzWvuPUtAO
pqBgyWyhg/hk2y7JIJe17YYSQfPIK2Ilt+F+RQ9N0zcSWyG+7442vFvCAsh0/tXg
yRn6RraV9zZU73edv3uV/I0F/JNgkoc3iP6MpiM4g/5vaO4+TaBIrTdJcpM86l/7
puWTLjjOD352Ge05sjAPHYR0MiCjf3Lqzs5RY817KC8JizmTWrFgVwFwvGe2M6lU
jCr8Z80dt302welxYxzwDcf0xCyhwj6yJtiEwhjMn8KaVIj25Yd9PXf66/Vfe1ak
iRkX8d+cx9SNuKnDQBuIY7XrR7W6p7Po0lQ52/GHR6GB54RgnxddDV/68XEIasj7
8aUc6RI/ktCve4cggEgvplAtdF1OYKuqpXPdmZvgJiQ3dVr7hHCSMayBg/Fd/ExS
YZsYuufGK9HapKefOJYm34K3DjeYFKglW9qr925K8DMHTACqCfUmCTi6g8N3oEm8
sG9hTa2pPupK1kQqHTTG0Y17RvGNFp6mHBOkiUJomuL3dbuyyexEfBWzgHK+22hM
63YQ6rl6xoa12dqr331gSWmi1ZS0gZb2Acoj7s8QonqLcbc7JXALiqFMMMOl93w5
alyx4XB+Kml0qRbMEHf1OpRS/VOxsMNqOmtn3a6HN41KfIMoYHj+8/xk3Fq0geBX
c4jWLOBvucOB1eoOKGukcXoJ08AiPQh0+K+SlquCI1/djPLazGRsuiuTK6yETYwg
9fiwlItVQF+Jh0vSyRQanun9WQCTPoea/AQXeURB3re/uTDDJ8YYRlPph1dzeuak
6TC/5+QB2uiIWBmQWml4+rC2YrPtoGbtteLAv+p9hO4zb2e9F6pEBhKWKadreZwV
rZuyBAW0sCm1CzCafSidcGFcJvapv4KRexHHjtNCMiy/txGsGki+EHyFTCJipBto
aj0hD62mMxnCnlQ6igk9YsNdLS9nQMUoc4EFUh8SZXPDlazE1H1zBliE0IxCLUku
qHbrFtq2WBVLlR7wfuRp9plClQMKZiXlWwVyEdlIOEVMbsrDtUJw86wgZnQ8IBuV
U0CPDc9TTC2p9TtbcyyBB8RBGvgOw0ehZASDCYfC4EFzUy6HT3laU3jjRyqvwqBR
kdg1Xm0BfoonccnxBy7QDSiGFR0KAqYotZ5arG4BWTxmThaxwKybBzFjQubZbw0X
bgngEBFIlRH0hjW+8k7YOjEhR1CzOp5vkpXeT8tXd3I8etVgwJJokhnUcR4TB/YW
//LDSh7IEIDYYWa/e/GnJhghwfspr0bu+aez3NPQwe1PqlRBuLgCS6BkaaWK2suH
/kgTw5QDPiwF9dGC9waRGgO9sYH0R1JH1GWT/3fA1SdKxaFQndzqRyFTo45ASpYQ
6HC3DStDUmdO1t/GD4PRH9BDlaBW8Za+TMHh1CeQRjS1WR5GXDtZnAnRfV0P/js4
+WgsLmNc+796iBBdBYs8aw5oM7975vqNsuKYjDu4Fk/WATl0Sr53sDGEfOiCkfm0
bG+28DI3q6pD/7pbO3vzNfahjDB/dAZEvE9wRWm3KFuluVlPesnBordblRn8tsme
XsZWzgBb9ZDfrAOpW84eJWrmJe9okU4OVlOos+vlSE7DL+wafWynNXBpzlMuMJEL
7ldQiC4lBLyu/p1otugKanLTvcLCRYUaDrdC7lJ01LIH//aaj02+1i9gn3Iby9zQ
d2CpR1bwWUE3hf4PV/eTxqVN+NbgnZfiCqvWPAzK6GmF6+Cmo5cJvr7Qnis8DUOI
R8fmKak2H/98gwbLMqt/yuXG99z3Cvm+MB+fG7giFp4rvmor74KCe9Pld0PJO8jX
JbGWlFPFzAMnMFnY/ZOBei3EBkuJYtHb1Y9Q7rbAflfNmZkz4USF8f08a3eZ8N8h
0diI94HvXjTvkhcPgAR/k8ToiG+otYHQu3i8fNlV5l1bejNFc1eynEVlkaum8GW2
T0cL4fxpaLlEwJdSXOYanIwrKWZR6dmg3/y+2g2LR2Vz0YXIqfNorE3kgPHUQAQW
k+aruZH1KeirSTWWBZ0pgfdoj8JcQEiHXrPtRPhCzPXDSopiMHjwYsyxa9bZnThk
Cc6+3RyfFb3eobp90j6LhNPHEWQelaAMNWEsDSn4wYl3Uxopd+7dNXAT7l3NihYL
MrM1NQxXt5PK8e0bx3dLtgcA//aDcI/XwdPiWh9+SN/e3vml3wAOY1l33ed4tgy3
dtmErgXTVJU8SDvt5VBCNX1kGPRjABBzg35ij+mZAGxLkdgOH56wJyjNFiKhZB8z
VHnNzJorzpim9FDWlLDhsIu/AAlaezNQl4ozPIzK2uL8+IodlzHpbU0uVBqJ2WWy
aFR10mWrbagxtl9Di4oQYh6CKwu0Y73n5dA2hEUnLr8WMzq00Uo35KwuhMJ8N/fB
OaCWd29FY8vMVphUxMjo9uBaDLVKyQXwKUwCO4pP1usNSCQyZwPavO6l/zQvoqed
5QYiJH2XPrHVLIA/YBDwVZt6Q11aCwUr5+2haO59ou6d0REE4rBg3hih76yqrbGt
O9Bdh+nhW0I+FM+5rbLj+5Q31M/ePa4Iiq4qeQCsr9sdmYVqhWDGvfPW4kV0xjF5
5fJ3pVIX8pDBCGwT58HByPxXIuttKBuuXGJMt5duOdtt9fiUZXVnEpfkHNpp1WHy
u6omP2joDMkmd2j3CPoJc3oSRVylcUBEBW0dV/yAtr2ie5aBV33KX/B9CYpeQ96b
Y+G2quzVXMcirEddf1kx/Gmsa7DV9Wsufo7nKLZofAnA6gcU9GxffLCn1kvKu0BQ
xoaQ3c/aeUbHP9CD/OhKk8KWPiTQ+6NbDjukoXxkGmSBv/kLAwCHOmXr/5fuswPn
2sWkBX9psn8Hgabi47WUbyKwm0Y68G1+tOekQwdKDIJoGonxt1qWuUzHp9MksJFf
rlU6HsDHlVB7zE4CZ9471dKVXEWpProFUGtAuECoImRo8q9JDSaHPDURlgaZrm8r
T8itJCMApf7FE+1G3nv9jtmUYhdEghL3HWvuevuTpzOvVLO3Nfk1EzlIbIroMVq6
Lf0IGiVasZphWto1xPIoZDooaKfx0bdF114+yFJ4XOfJAOOELgBSZusKOj03plVN
bfhT0lC1Xqlw2X0ZIFjSX4auwLbI5krTIzqu7IPm+R9lEK1rYETRtJZVZzxXXuI3
c8aJy5AzSfSfMSdSz2GnZhPUGtfgdjR9Ku7WwvipEmeZYrxXDVON0X75OYpcXUqh
zkkAYABrgnTl0qpTzYXMukfdpYU/FLzkhJHOyNqBRzrSfYbMx7aZzS5p34sO8EG5
iErgXuKNsEJRq7unAsqUjNvEbl1B2Tw8mujSwRdwC+NI9Te1+QW3278M87v1w9nw
JH48TJXBKINRcG3peAkIwhuCrp2Jy9QEn16ErNJoR5qBtXnNOth+IYSg1fUveoCS
OTpmCVE3t+KWce73UVMz7GhyR/IB/aaYBcxayMK34XKrlpKEid6urf+wGr+KXlha
ezLHWjHNvFDVsUlnmd3+48GT4A7TTBVp7MvOtZUPc+6NBlmyOt2U8d2GSnF4knUB
5HTnSmP132lIoD7+XyQ11AtIMiovKqnjJOHBwBujEXpvZ6Ci2oQ7HE8QZH5/5oDD
13oRio17r4zeHDLp+0uOufLmLhVVNR6M612QnV5K+SiTZ1bJUrA858kCNyIG1kaW
/M0CPWEwkKH/oQXmIOPdMKUtRefPGNgbExIjNwZMKm+Wh6LsZsbIHEii1pUozVcd
NXO1UrqRvLhgMwG8PjR2Sbmt9O/NKhXL8KJuBn2yH8yxSQ3fyqOENTPkqjgV6JB5
3J2RgsZ6rZiL0eOSl8lqbN2Zl1vuoJ6UHFzro9IPoFUbBBVs8GQH/L6CAH/eHbus
lmnG5Q9n9id1bnpw7C41UcpzdHPfNQ+3orVWnLKKJViFPzwwC7jPy+NXZ1eobslW
wXJnNIF2PAxEaO2QhyzAWKCDY8s7hEj/J6Pyob658Z9Idv5Fbmska7y6uUnVr5FM
KUUm0cXMYhwK4bgdIXDG2fIxQLoyyKBSZOin6k21NP8qtGMpN0X/xw9xu9mHMwsY
iUXIRZXHYSnVYezHUTDeffWqjpF/1AqkijIA80P2cfCXyyUEocbLRwuGkVrS0MC0
9t5NsK+eUZDmgQgkjOJlL7m+Z6eKRny3o4l1d4rA/F9f4TqDRI2nMHn46KX+gfVH
3+7Pt8u67IJHkOjC2wY1xq2ve0BX6aFpnEvy2lYm+FEWDmGBp1NzW30qxm/yNw2P
3Yzr9a2ch7XjD2JxTpizsT+uVEZ1HsfsIkpeQyKiwMvUb6Xj+aouclKxQTIBNKVu
f8x3evsPOLv6EVD5pCnPrHClwQ1mqtRxUwW9FFgKfecLDzt79d3o7ZzSMcf9FtAn
T0ry0jACoeCV43Sw0m8BcckkECWewqdKOTHVKVRXYyV0TrFQsUCmC+OBpSSFtgHw
pM7J5NSjCoI+R9eEoAOsrsy4tEZnhM/W4Nf6DeXqj82D9fK8Fr6ldEv6gd16bLRr
bNH7+syXrcyQKhHMgInCwOh23PC98/cMqX2tT1W9g1WdJktaDVNS9YMFIbnNiK/S
zrXLC/1bF/2RiuCo0tlmgt8qJvKdKfDmT1/OdJP9URxNB/+yudN7gpUJTrrJVQZ/
EhD5ywJRAeZOYDncYNoJgmnoEbplez2S9lOBoGl65Xet4m4lWHIPuZHbdESmpuw8
iVVda2a6LgNg2dE6toPh/wfij3F9OEfN2cCkn5/GbGShTt+Op5r4msAS1/6dWADb
BpsgUxr2RlEiVfvngT+/2a9HfzXEEAl7RntQUR9oVMfG2Diq6+XiXew0ZfpeKe9H
BdkCeUlijtiLehOpifUqkA0oI2bFMB97FNhI9aJMur/omSX+PsLEk38zUv6v1Dp5
mOmOk1sNLhq8KvtkNmF6QyQBJG2TqIvxh1Q1i/Rn+SBcUbQLslzsAXUqKKT/rq7k
z6PFdQisE3aB5weoXh4mP3XZYcre9XRQmSw/4jwR1+/QMZiQ8jMSyIXbMKumABub
zgxarjMC3tQx1DppoB+Z27xPkFpuIRJA8gUtjDXO6KMcwLXfbzfJPNpL1066Qdui
qSksTLOiqwIon/kKFuLjJEXlG49jsKqw0Blwsl1ybgbI1cvCaYXn6fDGIC9r/U3N
W6fUPv2aIgkS6xfBeMjQmzNFPqbElUNYXzfXnuFlOO2RsguVAUXDc0GtbymiM+Pm
NQGfN/9jWRSTKwa7foUW+sDiK09b9XKAlZ8WMIcY1kDLFOcEjoZg35nCOh9uMpMi
066mq56Tb9gn1gqM4KqF8jUK7fQ1dP1r+YKXBP4JiO1r3Z1gBlVMWR8WRL+m0mt+
9SbBZafvS+jJQMYHsA7+KKEKILptmtthf0ocffs9ugJ1whkCwciOTvl5MZMd0sj0
7NpH//Vfomd31c9OAFuSseOjkOQmOPpUz1ftkYqrTl/KpH68WFDhtxF+4xb1sd9O
pYP2JD0QohsACOpe6KcqfXApuL00jMjDRWElR6a2RdPk/R7VGDrujFIHDtdU1Hkz
y+D24MRuKuMdToeaPmBAXaxF+MOhR+mMcmmyEq1cfHQbYIYDZi4AhvoyMQr5udQO
z5PuDicgOK6v3yx0IHDiRd4SYaCq1BnVGF/uxTlpFFcNkVefUNEcWoc2YDiwytYU
4iuFBlCatTrvKymOgzQI3BX6gGE0zjyffdEyV5qLECQcDZp/S59UnIimOcekBffy
S7/i59+t4m7Czave63BkRdipyuGDAISc8kBKqwHdeB9fRg7sVi9ICKyuFYxrbAla
u+VMB4Ij0J9sH/YeM0ddH6jKJAsEfbPuyQRWfz2tgQOySbt7eEvJuiwJ1i2FXiF/
fvctCj/47Rg0aQwOK4XW4t7UVWmHFZZUuICPyeB2Ivdd4f731P1lodfEPISMkftI
jjAIipHbFNNbF1KqzDzmjHQJqxfHHF8zEEj5cK+dHXGnPMXY40alUETt5Pc/RZFe
D3j/BFJr+XDlZAqt3X1QL7zPwR6J+OrGc1yeOBkFhqmcK6JuvKfP8Z4COSz0igFJ
c0RYwzTwbn4rZmw8qIOJPcFP2+Av6DcCV9Jx6ADJ8UWFBAs/w2eQz02iBr7xPstM
sKGDjHCjR2Fos4eOGwhAS6P6yEBknsEr5utc0qBifJ1U2W7PQ0PTFYsfjPbqJla6
FZcDIz85cfWhGYkbi5q59MpUxa1fSAWjOGLhq0Jyb7HHu8M054LCQU7H1wvpX/5b
Ayw904TdExEq5SHRWl66u2sQ7sWjHQiooM+SUifOtbCNg7GSQSMgA6y8/IadFo5n
TNhkzp2V3PUXH0zKI43LN38hQKPjGLWnkVIxYJJQexV8K/cYnc4pmW0VqsXxFa+c
XKCU9SkSNep3Ah7SfOgf7YpDkGRYGCIg4sFdK28EvgonfVeEwICfAGzQbnF3d3SG
5wRElZU9ROrTv9oJqWLEcHgGjD8e7eJNAy4773S6f5YnGou904aqvoQXM4fCRZXo
i/zsSYQDqaaPO67kQT+23cNLfEuNCREluVmXOjw0wLPtUQodEv/JhU/jNTYWsQYR
ILTb6E+gr4WEOyYI0vXo3RBMRheCrGd/CXMMnOF6u4dpwAs+4H34XfT83LLqLOJV
HYmaxk81LrxoXLHUaBckEz3mOnTwLylzQpDsD3Y9H+apArueMaoitW0w7WywDhOI
32NxuM4s0lSQifwvXI8UCKySHxLZYDm2pl6pTySSoKGDfSRlv13rM67+siTXYxzZ
VNp84MCB4Dlioydgp47dct4al+7ANMSegY8QrtH6Krcw0rJaQ5U8chK3QIoE6Chk
3owl6s6C6qLhvzLFj8bbnDnavdrgrWvT9eCDVNN2WpDzyHqAN43WNTSKHhq28eMt
tOIeDxcaFwqAMammD5SL98ktzOtfrbwYcGyMxgREh7HtEEBztcaxtrIseo+/D6aC
Q/kJvsA25yRnk9jnKkASHRzrx8uV/lr/9fMjbg5KtkDZOeoz8a+Z0ohGtzusHgc4
Mpp4mEBXcSrVhaZ+pJfUalibpoQIqK6gpyTX0BX/7ytHn1P92Nncrc6W/5Bfhl4p
tYCutomr+9qzwK+VcTBCFqmP/F4ca4rlCQ6W8ZAEtWe8rIgLzaQViYb7MSLEOQqh
WjKnrqQMHnLULyBe07JdZY/cFWyp7YTj4EaRE1tyL3OoMJ2Lmd+axMYO+Z2SREWr
79NxUNfVrvvxPkvG14lPWjTKjHBGul/08k+ObJST0GxRZNVcNVLg08jfAseg5JyB
X2MYSAYzd4m7MAoyzeTh+ZXPTLbOHpYXNTQT0QsOOFnKammHap+2uqJEzTt0VwKF
75f4Vo1GB59vTrGfHZf28OW0rBDF4RLfIoQ+65V/swCrXCRiVGM8hK/uFlYMbjsz
NXQAHYB6oUssGEQVV8VxVbs5cV4JXqaNjpj2GgpNgClNkyl1TAXzPCK/aLsqORXr
Iw52qtJy7Du2BRM9e7vpviINMeIOgrvTdeCHRtFh8OZfb/Z780pkOZnGwpCtXgMe
QwtX2lBDzHvW0e93SFq4W+q17tLjvfnSQmd83jN0ac3Ma2tAtFxvzGFZPAUoMJ/q
b1yz5wLcTfhS4wyP+qW4WvASwgcwnZo+MLQc9W5C3Julo/UMRDAJH+qpkMUy2p1s
5OTrirIi/wP6Rt+CXni9p6T9m791TFxvDE3n+1xlIgc0ooCEf1QHLIAggwV6C6/I
RqPO6QuQyI2vDoSK2d7j4efnH3RHHXj/sxyNsn2ayW3+Q/Zw2bQ+3EtycZHLvmnA
ZiuauXIm0NjxxAFm77d94IfL7Zeu2/CJo+9pZdXzBu8XKZa5s7e/w+evF/ncsIxT
YOfHAsiKGaN3dzMZ1LB043/ig3d1FwKjh3sM6QIcRUacjimx3FkXqFBi/odBt1is
9wADI6ijHLTkC5GKw8Itc1PBUk6UrD9f1q6mXKw/Z+wWHe37veauJsee3Tt4Oumx
RWErbdWHLPwgziw05zO0pCR+5j4nuRggDKC2BDkS3H1yrR6eylWkHpt5HwvLd+RW
L1JjCNWDQXJEchCNLCC8BHopQORh9g7lnq9WUJRPY/ZzotTNvkcK/FoGSLvAIW+j
dusxLvs0k2Jof0tuvD9iHSb/7TZve3aEl7G+MMEXWIeks2jHhUXuQGx4M5mjx6f8
GbOchD+kT+LHANulzX2wgYwy8N199kXMu2Q4dWJ9XUeJdwwHefOrf6PhyxxW4g0L
NIr5/c8fAl9wGnfxRe35KJi3WVZZANOg476AHmP64fuZOhyG67DHlzVAn1gjGdpe
c9sUTSjao5zpjcPY27o7CeQuBfhP+2eMYUO2TdSwDdITncGI7DCURLFZuhCUn3c3
Fh9PQjfFOOBEpMTj2aj1j1X7t02xxSDqFuRWhYZ0Ku43PyXqWRuYKqdyiOHYiXmj
wW3OkFKlYjDcS6qF3baAqvIWsYEBawOX//tO0ia90+1PKVBr4y6dJHn4F6AaOGhB
TXBtfR+Pyo4qgognpXoKB1754UB5zC+qKKATPxwChyV25nZ66tu5/bxHzys+23e/
0T3QaF9Ue0VtVzjE9RiElbl60HuAE2Uo2OvXGWRlfGDelgGXNBUQxqm2i7N1bKeO
6uckOcvJhgPVkMzFnZ2/hVaITr5btYQa4hDaBX05Gr2IB0pWBCXjLeaZPkLi9avT
1olS9FsWhkNjXozs3oE3GJLn7EuxnzvjVFhc9bSfvuT5NFW2v2ClB73iMiclcW4m
wqo+Z1Ci90ln2E/3IJffE0C5t5So3nqoTivuzoWh2AUiPdBWcknZVZszM7WtwYDj
H6eJKG1ZgA905KQHHu+qb01xGnjGEpICqLrR+7DnEZXfoQVTox++2xuoickb5olL
fERqgMC1Vv9C8wy6aBFUU8QrB1EuHloN4N1utQtKe9+J78macyVFrw4GQpPS7VUp
65+b+MWM89S8xsiUyBsjHzqgKY776RKekvL+kGJ8uAMrniT5HlpLIugsKhaaM4cl
+AX7DI2fl8S4FnudVY3lhQXjU2n1e3THGGeg/xoR1qRHzpfvaIe6GQTo2wNeJltb
fXD5rH5A6nBWNaGjCxxMpNqwIWH1/0HHuUwLje/rl37R59g65VXMUhkUfgrt67ip
WyCCZAwLPRAg6jIJGS3TroU4CncNzoNTt798M+7rzVjscqz3QTglGyELrRWDXreo
sG0uw0oGExMr58rN6RRcUl8ELYwbosXHQbk7Ldkf4LRVH4l3v1W0wYsSwacV7XST
bFsAy+f4HJaRa+Qxqia5EVv+rEkMIv33dd42kjDeBjrr79bojRxAer8H9RIFtV55
7zuz7h+Os70MSJuJGBKCJhOMP1DsKazqOox+QNeRTTJH9yP5242gSnCvTU3U7lE4
UTccVO3lgHc8tgNPHN3wke6+2R4EHK5Fq09iAvRPc22G+zOfUf9M7Poy0sAXQwYd
laMIS3E9z1+5ubShiL8IvfaHEa/TddXr3ALn3wdnnpfjyhRon3zlbsuKVXqcVwtj
hfC8MJO56IKdDfwnm3rrMqwMosKUqmiCfUUDJkdQQYPqn6/YSy7+je/8UX3NKBw3
HE9TD1O9ujiTEf0HjdjV3Etv8n0pOaDJsmevqQu3j0HEoMvc1cc7+9FSgDlbTqT+
jPVHYgpEReAECILLP6IjUrMY44K4+cp6iY4U3t8Ao1i8BboTdpz4U/8W19mnLv4B
3Z/RRnFGghdmClgsKto7SxjKD/roFj8O3bB7PrjFNlaH5kCK59ehj43yp3xuy7K8
AJop0kB7ebEL49aH9DXAWD0DdyFamygMiZs/HUWuLyp3zmo4gDCmCwlNQ/lZM0K/
gGcjYfNlN5oZ7V07utjpFhYo1nUKPTOsmrt9oWY//o+MsfJ6AcMazJHuP4RMGcMr
cY+/+3XzdB6bCU8afzlkKOWDVKiVumS1ENkBOYwSbzWzUfeYaAeFR6H25PM/8NAz
90KU73HjiKUhAXEZbwQQtLV/ApO935HXGxzoztqeiL6qnmaVofcddXaObdgeIdDR
o2w8ktk/Wq9re1133DB41vm7GfAQIz2uJLDIdv6HqvYeezqMvj1HJk3DN9bHWXQu
AEyxmdTvgzmtXCvvDWPlC31sgweXiYKWZZz/gmL8bwK1D0QVzCICJQCN9KhNAnJC
NwFF+GQ/IewZsSqIzriwR+KN9xDHifqfbTfqf1qyM1SQS2LBgKFykDZRJYNDRjho
LFRIMAUtc2zD/uWMAOWhhUhp/Wti3aipEilF2nHPQNThVNofJrkF2vqU5yRKkQkX
zervrQL1Prby8ZoDYZ5ymuUXjENG6ZnXPF2q5w1jPgRySALkyEax/BNdJwno2t3/
4GTq6i+5TDQFg8CvJuySLOI7Yps8A+ByyqUX/HoySrsVeHaoWbbwVRTDJycb2zp5
9KyH0apvxfxutACMIcfBRzHYZ3mFSn42yor/ZZuyZe4t7fhrJg9LhPPHMPclBJWS
PQDeXDvIhsLzSND36dycrVUxsU1KAWg1Jyk4uDzu7poT+5zO3DheB+hqrgwgHXv/
VfEw7RV3/UZiJtoG47qwqIWaPJcx0sMshD0jhYF5oD/pDNZppenmeAulinT8VC7g
eVlB1S5sfcEGaYRNzIeajxbWRCb5dhBKkPcZtsaI3UEVdxv194c48+nttmZsa4dK
Ho1F+pxsBo5GLg+cIUmgz8njCx3oO0XvYwgYf5IqW6L4YZ8U8/bcxnGiZKUYWrxc
m4CV0fVQU2XbhpqOscw8k8bTRNO8SyHVqBI+TQyMPyetHLSuLi/kWCRgIwVxrAHa
iBSLwhqihsr76hGV6ZQwxsJNe+6BoWdGVUQHCGJJlKinFGNxHg1DQ1vy4VyT4vpQ
EhPpLRMSFd2J2ltjVtNu8kWgfWkX0JpmLvl2t2KEy9qDURoH5TnEeu9DWLvEgDbO
ROshZnww8KgYFCLsxCLjbYnS43ORLJcZJpQ1qCo1F5TTJR45399z1p/JsOGYDviW
AfoqImi+bzLvaiCZPLl/LrDlhFwUiqisXQM8HrWJlKdVyTbtrCpujTi/SGPO2mW3
uOAyYbRZa7Mq1P1GHoaH21p992sfzl8uTYlzRiVX+dctGU++LKWXxSVTyB5SKskG
kMw16XZ8AtXaDl2pQs+AKdv3BUmmbGyLTqRyuARGUTPxJ5EbBYLz7qy0VhRco6Yr
5sVsBykohn2jeCDN4qWzUCwokquJg1MUPH1H7/jHynfSCeboQe7keHgtUUIxg5rK
WrUyI+/pT7uTT0nDYBnBAHjN9xKle+Zz523fEE6DO+oAN0ea/ueCIe/k1fT5NFC6
eKzxIj+hJSm2j5sBGjoCCx7U8o/Fh+5tBNwWX16r4ty1vu2ucvozbz1QC/DLTBWm
Jh/1F+KodC1deUrFqcxn7BmyGt7Cmt7KWMwM/ctyAfIi/mvENHPw0LDTd5IB6+GZ
3zrH8HkQh94zWNP73PEgjwMkOqwEbc5RtZZSCxZLsgZ6JBt0fxwd12NK1YbEp/vA
e6iZnxLOXCOZVQbzRh94DJCa1bZj4LktlsCGEcNuOxZ7BIBSOgu2zjmpX/0LQMQl
qiveuO7O43GhJn5xhMaojd7e3fr2v+n1JpJK+3HqUyPGrEQ+eSSfwGCqAI7lcMHh
2jmr6i0D24XmL1mYKYGTPJtl8K7sC9SKUYXMvs1KFFWhmqJb8DX3+8OfSzkswQnb
y33nr7Li9Tv4X1B/vr7I6N+e0u4dckyo8/TfF78iyAw87MkLxhMENQgT8uQes5Uk
uIf3WVxhjvdku/STjH0S3C5Y8FdiRmRs2W339p8YYWz0SPJnoyQ1oiPhP7MLzxHH
ZUXY4s2puWgSG1XeB/fFC1KYHYPvY9sPNRjxuqCvalt3ONWKEtFKNgXsxvgtzBSP
CQ6Ekk84G5ceZBR4gihHqmboxvOTI6lxC3jSxcupMdN0K1cWIKhkCUiBE0FPHobj
LRWv0vb3GOmSDqFLrN1Gu6Me8aoozb8Xmmo5L8UuCGdipPj7dtNwYn6Wu+12kegV
hrrn4Xfi6h/ETgqRdAEWcJu3HzOQ2Bmy83dPUpZLWnu9M7zEzTv94toyfgQNlWGG
7fJ9AX0paW0upQ5bcKvHLYc3KtHp5EolEg6tMwCcyyNj4jWcVAQLh2WxLGPOm4rw
EVSutnMWGL0f6W7UkoCuM2akIcHp9d+EMKp6THYegF3h5c0eeck6DCc0S94dO9jj
z4OCPa26k+JPS3fTZC32Z3o5ThdvcWy1KcwehZZx9HB4SsPntsTAaB/pYvGUAxbt
0HyLd3Uf+CbISf3saT/BbWbHwMdNqdR2WnFrPWFH6OvbcaYr4AviFtMugogQoNOE
h2ny8GRG1sc/1QQEghODARxGx1Y+Ihl491Z87UpLoocClpeyx4m6PbwLFnoeaxT0
++NfKIkVhMZEJu7YJSHuulJbpTAWoZKN9V6UeOaBXqiJw7rWUpeEV/s5P2AynNa+
GbDn0U70p+L+rADDFM75sVQgpo02jwne7H7b3TfUlGNKd1mghqUqfgJEyNhx8SRB
DyIMYSyNo9zcgzrj3WmCe3RcXnPbLgI/ygemQlnEas+ArsqWm483I46mgJk34ztW
4R+T94cPFKnfLUmQKSKpurrc/W6uoBZZFcXPhymN2VB5VQ7M2hZ2yRwoa0irbDFX
qDFifvk9m45WoT3a2im5+qpkapaXim1YKmWoP/4XBAa+uQ29CMhBUwXQRLBuXkz/
lz+EThnw0wUU8nNooODQp23TiwkuKDS7d+JZu1uzJgNEW+2PHyOpP2G0ger4eknq
VYfVwrjjjwFVBqW03DUpspUQkAE3c6Yyx/j1AIvKf33MtVInvU0XH9KpNiZ3DDTP
s1dasStjVNVTd2xMeg1mfljKUvlCw3UtpeBtglV1PfCrczoyyFfQiL83xbpGCI6r
aOcKyNc7l9/wAooIaR+2JzGIXLc/QWqFetZGHIOiQ/b9AnjufaxrBsQFP/d1JKM7
cTKi9YVAuT4I1fd8Q/L4d8k4faEgdqnOzXxiRni+PTdpuYGvZuuQjkbgGL+Zbfqn
6ksH+JjktGxbFo6j2RyJPJ0lkps1DK431KUaZzT365lRPv975ZiXDlaRD0dRmr31
Qr/4SY664ql0pNyimOK5g1dTLKPJVz3/5C1jEn2+inx1dhb/oEL49n16eY9I38kw
6EzIGt/lII7eThP2qW+1Ze1G8foOfPHs8oEIZMdgIrw2A0jvu2nfToJ7J7Gyuhax
0sFGau+IkPeR+Kc0djgh1NhvnQd1mJxK/y50ln2JgYKa+Ncwg7MgHQqjypwb4ePd
vRvbT/fWETqW+OUzouspqrvRPvNCVG4FmoH6oseleaACDvm3PetZGSHRCcyDKmLf
jZGjJa2NfVrTh7ay9seHGGLvYu4W2L5pfk75iddQyorkAIMgrCvocHZQG4XvXw8X
1jZOHbac+YWH9TlPNFI9j5W4qbLwMeWKJzKhd8Btim/Sqb+HjKXmZzVD4EZjnKyb
fSQ35qUlwRcaRGE4DbX5pg2TPG9/1aD7v+hYT3ViyKVojdZyNJs80/4IDWCAAu1L
Rx1CBAAj8q0z3jqs0E2PPU50F1qjj6yo1KZQeXjV0m0WpXm6/GUvCUojZZ3zLkS2
pKatUeJTiPz6pJWi9aR9di6XxHniYWyL3r+ysHl6+vxvPJ0WO4FwuURACHMzF6vB
zfrBZHhFOWdrpCthBY5qCCWzwlee6ByWhUui3UuzXDhoQrCM5UHdsrU7eWBYMJSt
SWguj/FiMlYvQJkbd7kjPhIE5G2wVhI/Jiek/F/MArgbIhZ/5ywwIZ5zr58PCjmx
3fUBfdxSvl3AChh11eYmjfKRCrrw32c0fij6c1WLzlhpbmGW6uSA2pOA6uMwGuQq
71ILBWov07QpWNIZRuTRrudlL7PJH+trHKlCsgYd/a3he79jfgz92bqzvPWQcB9q
DqL13LGBLixIuOXsAQDtMvxGWH9nWiPzrnVQJO17S0n4AGTiJwq1Sx3LgIdebi+n
EbtHgxb3zQyY/vySPh93KDPW9HWIO3IvlW/r1NnZ9JjQTKM8DxiTt/K1AecWNNh5
Ic/FsNd03H0uVO7PiOfx7br0wE0zxvquAAU0FC+6LNbAFHEs6Dj2WBhG7SVALan9
nmxOWHyWAeC+COXlCctZROb9GCTxrEqtNN0O87R4N3mivEk7zr91fYUwhweMvJje
tG3ZD2l9L+Fe4rEjYtsoBgOz4umxKGuRDXzHH7veNhA5Y3TDsmJbHHun7L8HW+73
xT9JwNymACBojW3CnfrC3RzXV/LG+peGBnkpLWqNCD3PFt6caWxeiurMvBAc4vRz
HtZ8+IZI1kwMMOBZFWoSgFE1sargqSRGnspedHglvC8+RFh5zQDkvGI05Cj9Tnkd
YZsDGT2HHHicovGtLjAVc+Srm1HHb9m1kEenEN+8MVVxmWQnajvBhvQWTV2e60rx
izOV4bmnzhTzaTR2u8Yl+DO7SgOiWRkbLlp2ph0lbMO1ODdl2bQmwlyBMauvSpzS
jU/b5dfXV9RIfoTq6GMee7FlZvd+4sgup3WbnPYaTnAaiyl5wBMUp6d8E3X5vogT
PaiYkxrZwChd8n3WXBulLvBdVrF9XYTm8/HfKwJ3W19mzAsTRyGV1JRoz1BMflIb
ysR+aOVNEwjy2ovcX9HdIZUJADi2o2dp1Bg1GJ0LzGR4PLla0cVXklMtkO853I0W
Dp5o14/9VB5ta56Bv3u+Dlfiz+KtJTXvdmRYOxTk2gLk25y9ph2xVPrf/Wyvgw1Y
tuBFiJRt9WiqGaMUJD87dU3VhMq3JWBXzKMk9Z3aQfY7kgswZf5G9IdbAEcRvMWp
5CGwK//nKgaP97lk5roIhrR8pdQqZCpFvV0UZ6kA0iM8SRxYeQQy2yOHAf+orKI/
w5rHIQGnUm0Is8Uwu0GDJiMkWyhnknmGQ03R0d33405B1vIpfc91M6zNKjbvB6AH
Xc0tZ0DzzqBYLSSwF7G006UxtISU9OyVS0/LO1yzR35SgdRW1U3X9eSUCs+pKxAO
PCvUapWq7BxSqEn93vEpmPhh8Ll+p7UeGTqjjM0ym9uZVIcgC+qRb4ZFXEuQJApd
QBqx7zeNvOB+eckTl4NaAqdhn2oCJWSKQVwI+E1yFnoj2vuikyV2WHAY0pj06A84
KvMZv8ULy/BmbY0CrcbsvoHBpdmdDlVRXWMQZ88HZih1q22tPiwvrpe8ZFb9GQHn
C3SwNv5mILixqFjzuVC92CRnUn2BWoK9i5xv4WJE+6S5xEVPOqnIkgpMiYzq8hCU
RnmEy3svhxqUwKHPVLj6gR2mwDk2Ww0V+wdJT/NXVjqXO1gbF/fYEGecMmp1a3bF
lWAimYwAg2D2JeN/oVWTHNMnY9eAby443BwL04T6c3/byL619gOUEh8Y+uc/gx8T
A+d2oDeCmkcZBPd/HVjz3vTg1PL/of7i6li3uydamAQELZlbFiheA37huVBjCmA1
FPvhM+O/2Z8PMxQ+y1RNkGPC5I6o7hHf4LolzbR11XsQbeRiaORl86qaHaUgqhTt
KYNwotMWHpuBDCG25UbO2BC3caOpX5E/hN1yvVoB+0J4iKtCT+P7WZbTo9n4m4Z/
HmEt/RKlMlKevO0ZROnZbLvtbt1MR4YWTcySRqPO5+XAmq+QdM+++Rrqcy7/lAYe
iU/4aeIPbqfkwD++Ux1pych1wpdmXEhRCarkgfbrlRWr1PmDkfPIaVsMUxgnrQab
neYzU3ztZ9Ez/D4hE09bcmZFQxQgplJIsnErcL1Jzom5fqXcI4Yn6Ew+bqEy1ava
zXxZK7SNhK98uUzfxAZJAhnNZzzN5K13BYY74ByiaJlrLR/vtNfQaHlxUuDqvxmp
dm+KFJgkuLvR3knK5MQbc/D/+MZDlN6ZVAUnS8Iy2aUvOh9mtOySI1OBgAfQo0VM
2cZcAu3gwcPO273Hy2fdnCSLfxW3qLkWLnxzinCxf/36srZTx8givSHp/5TqKs0D
FnX0zA5Vwfqc5ufjBFc6z0D4/LcjIwnFYyz5PS/P0OkEGhbHi/A9dmjPVzQ8l7ME
yFrHuf4lDBuFKRlBtI7KU2lk7w2AQvzG6oDPYgEY0+/wdJUrG3qz1JcYCWLivQ1K
rPbxRnA0Mh6TUsU1Ct8AGcYzU8JJ7xfCe9pvUyU9t39LVyBedGPcN1SzTCelNcYc
ceVwym7S126AX6KSsggOmaAtgmIoVNtI5szVslHR+Gys07o8FrRkN4sDSd4GVhCe
RKYMxMljwNEaadqmbp0m2f0NITzfJtrNwMyW1DnFZ7Cdgpm/1P781j0e1Gpt5J4a
oR5RU3UJCMB2M4e6E+9ag20CgJtly7OuoO8GmqGaS19nMSz5YU4GYGBDv70recva
4rYJe04/TtPfNGuodg9RaVV66wUZqrZhuN8LvXtRrIJDcui7PdyyuEKoC3vj2sal
SnAc+VcPw3l7zDqgp7sKWX1gLvjAA9wCJ46NAckCyoW6N45SmnwIZ3x2ql7iCAof
dRQ2t3iZCDPYlm7PvqCufSZRJ0+3AItBrNDeYDqX63pte6GgyJIMcBiAohTxlf8H
/cW1eEVWJ/htaspxNn5ObHsdVL/Pdwu98Uwk10hMAMRMAiGxn2dQfgMDk5o+o8xq
WR2mdQnKtwRmpzw7mYEgqrYVL3u/k2KjAmO6X5+iDj1klPHZZHRPfpVc1NvFwx21
E8ZjYA1EKYBeKeEZbQVCXfb+EvhJni5CQdBzVVhLAebh6wOsMUfL4u9aoeDrZDkI
4OL4bOLDNEPZ0wPHkOvKSUufudHFRsB9xgdy/WL6Q90MEm/DwdI2YQGGPaUVqjgm
w7UWfuKxCmPLSC2KKw4W0e4pxTVz0kZi9y8LdtupxTNQ/3BTHUoXfwOqmIfO5STA
wryrBSujru+XrLiYQaRzA2XDyZlPKm75mwo6U8vCeHuIcT5uIv+bA0QE+XPPOFT7
qiqyH0R6Wgxz+XvhQlcmPbuKlhAuJpTfpanKVeKh+nPIxE41j7lrPGi0wQMubPXr
ac55G/5kIsbMo5CJt6tWX/aAvwXM4Ae5El8wKf4NiC+JjurjHHiZklchUHet31sF
wmkn4i7ML4Nr0TqgAX4aCtm4DDJukAmHO5bLZV32qHM9KnWEoSURA2GkMafLPkJj
ajyEJJdFSqTVHP7ndYfkPnPAcn6mx/5xHs6UboiYUQwNzXhLDeJbVmsotaHYgOVr
CZ08PF1ztVs2UoFNlUsSeEKsMagcIGGKmAmZDW5iP+JNul1Sz+fo5Bs1qQ3a1Cju
0r9M1D01HprnHFNuYqdm8L2htGZbWXBktC1mZcUPDKd5RAR40vMHjPbUu3IL3n+O
TotsNHfSsMDgZamzcvgRNiI+Hj/5P5vCRP3iuPLRHl0K8mgUUXNn/mlxuPFyL5SH
CCVCBXMYu+yJNuc4xBApGW9x33VPXRxTe5nA0CvzqY38BYlzaKcsOAUVYeKcklyG
YS1DPdGTqUoiCIAecBtYexW/4BVvxayn/JZZECV3FPts4EkkSLCrTZo1qxdJgDAX
VVWcp5wbWLkxTdfRlANB/atoWXAeNcmDUFVVTGCmCLzlzPcJknQXRXe1yflNB1Rk
DlmVCy2JfmO3u4EkyX4dyrOhvvLR2TW1C/zsSfkxrehdwY9PBaieg5AvtvnCG5t2
xV4GAOLuDcuA4oPQ5M/OmMGpeSGLev5nGnKYPfHv8gbU4PRylLbaIT+n5QVmXERu
Kth9rk+/UuQ6bF66OqsP3QYsxrHqq4iphoZQ2/b5MOEae4YllbGRxBh7iD7oOxPc
DqCsKzfSUrJhH1z/f69tOMSj2wCMxewXJ1oP/G0qI3oi2hH00D6AvqT4N2di/ozj
yI8QELqCbvq4mWQXBoXr1pyPwEWOmLs9x/4E8CxOyDn1bs7zatlv6xlfW1535Q8O
0qLScj+W/lDLJOgy6SWUo5P723YO0c0FmmNUbGlaWfs4ClaJvJOaVYwOzDiI8w4O
OvlHkdxHOqjlcZmjVq5kTSpCHynXwtEs9od0RqUbsEppGNlD438mMATLXbO8Ed9A
gjwurJdA7lBIajuMzV3LzXjJcJEOMetZGCpB21JDiQbs4crFKnuAzSoI12t4d6wa
dtvAO7Oj9PzWT3p4fpxPhHNNnNEzHw176rIKjQXGxeXOCl1Vmcb7H594To+6gK6M
pOp5RVWrLH2enz0pf6SO6+1motVZq/V5r91JLm3TvIsvFv1iMvlqoy5bNiTnkTbL
e6zkg7A1oywiQZecWKfwE9vwe+gPrnYKNlqYDk9CKPVXqQQoOaUa5lZ7JqwozuvC
bYUSRBQgUXCrzss1PPggX96K2bDwCLjMKW0DAdtEo28IuyIsDKOEpIXV8Vr6i7I/
GjK1hdx46hfmIFQpU3Sni1g1YyQVnIF1u26Ke4BNh0fmm6tV3BgHRifT15AZQBzb
uXaWayj+g5TezS0qG+Z6kBKI2VHk56gRmjP9isYj1FHX6NyVCOkYTFBdHvY8R1Ei
zH4HE+EwUU6nRhQVFabBBluVLuAL5QRFD0MDFyUKISXlO7irlkBSlepUXP5ujSrx
tDuc94Lc/y1mySZ0fJ3XIw5fyScvN/011hCZI5LQy6ap7JoiBnpT4444osARn4TL
+3exx4SsVaffZ++nhrqAYJrdz8i4OULv26W8R+JoTqNHZVcdM8JKBe6nHYkFEifX
2bIW9KPZvT7EKeQAzJCWZ4QPhO12VYaY9v6natexe0gOjap5SJL5m9fBuifi+qwA
y0pptgzfl3rsSBUta+FG1NeQIXKSXmN34D2Fr+YBeNMLhWQnU/3U4jGhWee/kNXl
0pVGbeuDAl1Mr9r4NqkXmy0WTZ1cw9LNzTqbmPD441L/yNzNH9r3vyhKDQE8Va+P
htuXCGMrDZbLgW3/IOtzFVA+M6W7w+j+69tpp85d85OWG7505pIvj2+7Ylvm9XqW
lo/lurXSN9ZfJr34XJ7XWjfv1/wsnbjycYMD86EiJ8jcqiSK2y9MMi9tjpsMOgZs
3YD5qVWoLU17BReCGjQj71cQdn2Xyp07u+bZfkcAWX6E9WOdwtmh8vQ+mCc7W4Z7
CRZCmlX47eSFbvyNq6W0V2Jvz+UWw/jydEq5mn4fX9L6ErxgZZ4YisDTSJHiKgxU
mCgpsAqGubT5xHtEmOEHGf7abK5SuhK+sUrSjcEGpyBcSB2D37mGDo+F7Xe8Mf48
SyX595z5W7c2jqikbKmdEiEH2i0M1wb6s3sDamJ/OhlTow+F80tLHCbNfZQ9Xdx6
zhYusrMKImdmEMmSzdbW0D61bJK99fABK3Szf56DgODfaxxX2JY8u1y3oJ8gRgvT
rDFuI8VzGtaUarMcvtal1MFS2/nUOmZgBmjUhKHudUf4TfVp6SIAUUykcq8zLM1A
MMG8HEiQQgdj8zwM9bEN+0FwxmSU8FAFy1kMl86ASsUNS2Xa5m8C8FAs61c7eMMd
YCyxOxzwDtYlOlOLoI7aYD358Yihi7UFYoDXFYU1yWH+a7Vt8TKMkzh1Hl5ZJrk7
TcXjgvJ8wqA+VR6zP7B7JSCgG6qm9k3TmgSUXfP24RT2sUik1LpvQwM4tNjPBMUd
0d07ffUnAAOBKOg51kz4VPvCPzwCmXcUwFCDCm9p+P+DSLuOqcut4RDcwByEWiMf
ZXQ7gN64tniGJBrEMgxLBC+e5Wm4SmiI1nOGfSsk1rvbVkW4XggnhtkVhN51Vq2F
Op5yq5liZC8hMfyoF5YwQvJeSwN6TUQMlCnLPkkEzfE96nyD3lOHeWZioL8C7A5u
58AF8frycHexQqS62XA0tmlGWP4C0N0SGJqp4BwkCflcEzsZUIiPwVqP29amak8l
3gUURpCCY+TmXrtEvTG3Fw9SBEAr8CRjV8D/zpruLC9C/jZCeArQ9xB3WuRHh8s7
qzBIGZvQ6xumLtmk6ukw0sODkFfxlxSDNH6TAxdOagX6jfne4vg259Jwvc9qJngS
dDDsA3/F71Rba7VES4OgKKuIdp92JY7gRv2j1YZr9trmi8E8jWhU6cpotvZ8MlYN
9diuo9efmozrNMpNcaRmY+v9nk8nfVdhD/kTHKV9M2lH9IBEpHFpb8wmnWMx8MCk
EjrEHEhe4pG+QCRMVbk+IhrhP7i0Nm430uGgUsHWihdKV6FATPZd+Q2iit4CovxQ
LPPMNIQ0kKK1JBqaftS27A6Zjwanr0GCyRWopqrPTxR/y1Dq/Omi6ba7BFc9RdwK
kmjUptcT3OmjRcAxMI36tD6FlaZCPewdihn4kzZyCqVorQ9iUUQFmCqBr83qNQYP
e7QwhQ8r48g0M9SP97ffgtTaoaK7f7WSWY9VTSIeXGw532sQQKDnDaZeTqHbn2EY
R2biIYgCn63a6SzonaGTkXR63c2HcASRa0F1PnFN0ud3zg880Eu7Tg1hengN9BB6
lZDyeiHfzT93waz/OgjbzwUlL/Uzfb3s+Fkh0Mnxo/CTrBk3tU+Rk8Ny6ZlK2XyA
H+gzqUegaXKQ+dEVJfxvSx7ZwuKkHjb8l9hN3H1sG8aJyREXPJYQiLmVrlikrzyq
L25/+E6Dnt+2MIgJ5nrz7G5JA/1wXbv0PPF1vpVGijz5cazkKBxlYTOS7QsFhY9T
D9Tjc/aNlhyg4dbkFIRV98cYmFAE+nA4KG9NZVhW3EtuL6KoLkE/dvccqhjcAr82
lcvAZ2ydRGmZ8gjddamvsPS/HVylqUO94//4DFRgyqp46vXYSICDCsDxejyR/Vds
Mrd/zYVPbt1tv24VQWEaufPT14SU8kSitCA0TQG811QHcI2xT6Or/RhMZNRr3Kt/
OxPuKelqOFqNwYGOS4IsUlCzF66FftphvoLNEFimmcgEp9poHvHNN9ckEYx+cOR3
rbERXKqp7SPQ40OX4brHMR7V5rHu2NicLciZZZ9UNfp1Hct/TDOFbgeoS8BitEL+
9eEUKkisqXOXBEoPP7+xyTp1XveJHsMVZmnOnqhND/Tr1x1JZLjP2wZ7lOQiCGLW
FD4mBDhJ1d34/03pylktoyv0aCgWHvfNdhSkcLOWPUTHkUf9g6nsL4aRB/EfL6WR
P4CLbFDW9F6CNBLk3eoC1u5DgSgMl+3xRH7WyjsS2uRP0gcrO1qojAzKrsEeLAl8
GJJ6KbMHgPFey8y7XZVYiySDBFxZEqXpJG7xBQK/xgUKs0v8+Uj9+O7UHFRNepv1
Xv/VQ2yF6qQlBgYJRdf73rwwYbfGsInxz/QKIsDBMqNpDS6mTixc0NhmTCDJj/VY
JtnhoNYGT3pwqT8s1JZu85H2Q8SsorMODRZOeZ36Li4OpMJGg8kFuPGgukrZbezh
z4KBIJ0h6rJCpgRwvLmV6Qu7gAmKvTcYaUtWEH+EtFoguJ8WKgKq5gN6dt4mxnci
ZGwyp6U9r9l6+FX7mU8SM1fWclI+Inx7X19OnEjX8Azkh8gFY7AptcToFDfhJ3Ao
laVHfgtrNLSA4udmf8Qv6YHuyNNp+DClJJ6j3NCD0TtbgD2DtiMJ8icGJNzuGZbU
+1fTCMeJkkK/t2rDZREL7f55FPNz1dBDHeTzcf3Y+N8l8HUv8yYHpnWPYEkKySZT
sW4EpCZLOZ4bwM9Vm8AR4GBv6QX/jpp+J6ugusW2veGEaNTsPKEqVjjGLlQ9Ug/H
ENZQA9gNSX1s3o4aX4VghejXMhKpywP/Z2qGEAzOwTv/y3FWkxviKg370+TzufGW
+OOSMH/oKMFPfqWVmoi6VkiS66VMrpuRp5tmossX2/3LF9KTrJYEDciHbyWso4dp
ojlGw7KInh7xk1iBMqeK+CQ96AZveXzNk892ZEJ1W1FL8tYOy44M8mTzqPo0WEUD
1qA1gOPpf7Lbtas4L75QBNfbi71zljeRSWkdGeG37s+U3bhrJT4JyZ0Y6GRR62/f
WCyBqhJBn2f5Vm7IZQK/qdK/wpGGpV38R/oI/YYhM77WBrG/32YtNP6C1+uVnZ3d
drrbOZjG6+ZDTnOEfqV/QHJjumbdh6fjloVeB8pnWZB+/AOtLn5Sgs6Dfh8u/Bbv
YCJpj05AewnmnQpq3zHZgLYHJBvm/NjDDp0YfuupYG/q6lXW9+f9/qyhlXAQ0VEa
DWnNPKxL9PR8KGYyVRQqUtkwNztZRa2uTCWx217542aUQJ5No5dj+eFgUqpBwKtI
2qJdyPiBZv2b+wzPnBaV4b7lmjIYPBkJTJ0sMWE6r+eE1gvEimt94ryihCR+gsAm
O3wRcOdaFVHGeFnokdvaBtdPSGFYzsoEqtMNFIrxqhlNNT3A27Ssuqkb+/rMBfmT
+1GoIFT92S4/wE8Vzoplf93L0i7LaS/GRoFwX8bFvoW9xUWRhpT6A42jROfl7GCE
wcK/tbCZR9xocdzEbp2OgPlzxyG1gVHZoIEQZjEDhE6fzVj1USUJ6A4fUes2IW0I
gJebLxtPOyU3SAnT0DIWZJVw7cDx6bHM88jnGQdPQJrEhmAuXSrWac3mwryNA/ns
5E2px9LmyjJomN3v7o8Bw5NcNK5wPUyBC1lFAPwUz/KKnSFOb28vw/DHTmKf8UkT
Jr1vmUFhZXWTh0CjYU1psbpVGK4qkAW0tESPhHc86/oFdDwVRUuyIJdfGqFjNUwM
4wwAFQ/8MZDYGKnLelf2SnY4lnSQGk2TDoFFMY5vaqtjXa7hBzI0KvkfA8DZZqkg
+W9kW5iBAy3ORIArWnjiCLSo2ShcQziJIdpH8HfFi6NSwp74q/1yQJAFm2XRfQnf
+L/A76/XVWMeTd+6rVtyq9hBZ5KFSVuHn3Ejtfb3RE+AyzV73bFigptIyTc9/rTo
4ag23LWln9YZ4715O+rkljNBxo4A3FffPk2kJqWQFkoBGwb+cDGnrLOVOidXg/dM
Wk1jDghRBnmYlLLl69byJv9Pv9+Tal2Am4naVJJ1xC+QmG8VCqyiumnMNS1G0txx
UpxSoV8oXKWkl+nZuGBROq3zV0jokFDZkZvs6vKOS3xgcxTYXKZgj5xRPcFtvctY
8WKq9sxb2QLjgLQy0eU1VeglFctKhxIbDwVz9f+YHwwwv78l474r/tBpmxrDEiYe
Y85Vqk85su4f11Ai5rpd0N67sE2QdFKAyDIFTDCp9t5RjvUYZHoiLGZNL43zvfaO
qrU0mjnyZ89+S/g6QAN6zu+ibMmdte6Bo6m561py5zXfbWgvcFB5AJxKAgloGavc
Wd502ULHy0fv+4m3NWFJLoaAHctvf70uQ2bf7LxxtaMMq5NHb4h2wXtTuVr8qiuS
rZbUJt+IedIwdkovWxq0fM14v5HRMND5Z8pYkssffEeN4hwQl7Ap814frEbCRTgA
rCAYDTIMM2RoJYQqVXMwRPCGjFkHVg1Al3bYLr8ajk1YlPTeyvZCj/mqT+5hsIY+
qpu7KmlecjZ/eBQCuvxxrK+3G7Vbquq/WW0AKyEfyV1731Vy94hFai41Uu6/JwSv
J/EHvVZf6a3tjKUjUzZjEJ1WfXfQ0KogYabGUcYhynUM7RIRDk66ncjBt+zV36bC
bVLMMeiD5Ik9DRtz6gWoluFlZ5/uYte/V8I2yFmvUYmvXUhjwmg2pg2V4RkqThUG
e3kFwbdc1NbGT1zoTYMdCOKtXc0BXDnHtvOw40o9d0zEH4fxzPwlTSvKpCWRtx4Y
7vYG3pNaqWPmyNdd9FGYYW4Md0/f2XnYpUxKh7BuQSpCZrMyZl7t6tyNqhPRQUdK
kXhJVclzNLFSjDXRVFQFqWQDHzJesuT9g3G8wYnbQ8BTPe/E9RBY09BcSN4/2Dp6
kOyuSQ7XKj6keDSGFTWzIbdQPtmOAtdFoln6ecA2Iroy3uRCNBpQ9k3Em6Az/U+s
QwpezzpqzM5yXOVbRdXSpLaGtjsDvtTjY1tp0C83HdynXS9BEWso+ij+OehdThfj
zLUZ9s5vAT25r/kA8o62kCKHXqXdr1r4TZBm59oG/AUllspbC+JxsO/c7HuxQFqI
+1rHhWdO6vqbwZQsN8MDEYkDFhhXZoDKfRwoosoNvTcjp7TONxK+yeYiifB0LYgR
DR6Wc08RFJzt3m0rufQKEmEtyw3iGXEZJvMEpoAJN/XxAj2Q/ZTaQSjCC026KTa1
IgsiPh5kyaWKx2p6EY0lZjCtJDK/zs4+7gMdstd9qHSntuwDdZgYrpIMJm6kRWLA
SJVWjI8qNLitPsWxujzyb8Lrck1vBDxcfjzxrv1Aswpi30kzcwmISl9M4XrjTWhg
wvbiYU9ig1qtgNo8VWyL2HWPj3nGldaRqPLJJSAM4XRvwamKvDz9bspyuqH5RF/B
RSrskhvDczSXFN6lnEfPMK+ecupr+LibDvLFcpKOqA1NrqggdrS4dUrc2PbYssoc
L0nxQ2G+ZWmtvk2PBehXQPTgkGXw+nvaUoOCeawe0AqbNIqJScwx3wHtfY9JKb75
eL5pxrpmUKUzyM17Q5qQvk+sf3PyizuCaJwkFktcRdLdcaz4pI/Meh6XycE8uBBs
RMwzkaliMzT14bwtgkH9IYDro5YLn73NQuDTdGQ6po93IgEdwPeCNjloV/8ST6cj
QVKeF1Gvb3bACXn4wNRDbN7zPAGcERNnkqDOIMVW+iJPVyVuqx83TRumNDzpD/xa
MBBsreg43uUqcDBXGB5HTknczaSLZPEqyFUyOSFnj+l+cyqqRUrROrdv4qXAMr5x
zinXTb/lL3xbSFjV/9mwbev4QzWla6dViDNtzqMYR7Cnbxgj/6llLKfNvVZ1qGpR
Rf8aaaimFstg3wmoszJbkm5//flzQedl1Usu2a2k28sy6fO0T8xewK0jwBKM+7oR
zGZIKCozXRVqh660Br27KdVkdcgFO4y9lTnepkdVzvAn/r4vUs6c36y8cGrPwOtp
XCaJazhccjCw42YFV+vas3D4WAoQe22+r34jFJNB2xeoAftNGxYXOFypKuTegqL2
ruXSn6qqZ2vFU/JFYIifBiJNHfU1ebZc6YTJluqZ9H09oMOn+PyFDj54v2bDj01v
8J9p62SIipwN3dUlfKU66qyI3cKqoVODyB0NvPP03lFfoall++/KRwLq3RZPrkP8
4MRyT9FETUU2A65gRC03tgbBclGi27HN/UWwAsrjQINRCg4MoGiZ3tmPzqenFKrG
uhP7u6QHsnuOT9s3ctOs3RByEmXYpdyBd3r7ZLUTTQLhs8b4/NfmIOr3tCNL1U19
mABMLKiGJCP9MUaiQj3KvQq8mHijjEDl/zFmkMFDntLtzz3jzTvFEtTCkmhtcTMP
7uBFL4F9k8zbHBZTW6KWAU1aFexVRVyYGS5Uh2F5p7uBX4sXJqVPNxCTCocKdjCp
slowFp9Czw9DhQzDFOHLgdR3fdCGIUKWheYt1dPy637FjjgDuR0DC5ty0tjvGOPh
GngWmbPWqc/1Ed/KPuamVdJCTPkgcIa5GPSFH6EBcNPaC9xrJgAJg1rLneaa8QWo
l1F5zB5QQTJqrutQQKblo8OxwHm7CQ4tECVR/6/KpBb2/Y0ZOobS4qNQ0fcDpwqr
Syuz6CFcolH5HcLo9xT48Uurt4E8lpsIOzLdJAltd928RIc51lVwgJETZvVkGbIE
/2g3fmuuZ4zTEvd7+6JB5d0pW4ByY5Hvov6HgzwsATx1BgXp3bJZBEa6WMTiC7Lj
jp9jhZkJWFjKUtMNsc6Hc556chqtLUYGADl27DTXQwmRVGBA3lAD+LQolf8azKjl
Sy2+XZd3wrHIW/kbeVcHWKFfKHsmyPk0BF2xWzO3ezCV4dgjgAftGgRF7neyT2px
u10LXrc+XDeYpgwi17yR6CTZKtRGLvvL/iIVIjdEhB1OqxyWICmJsfgVdbWTtLCf
a87iTQtNOfS7dgxTbLkDmKBT/Eu35bUQQsm7I2cxjoDcJr25rm8L/GakrunXDf3t
eZ5UUjhQYvWCNbuLnJa/IUPsrhRVdHJ9HsvpAPwJ3xPx8IzbExiK8nwbnerijQS1
bXd/QaBfWmIRZCGhO0n6gNbYBES4d2YIvUKJNPwwcPgmxI9ruekEWs3SzywbN8bq
8p0x6SOJAFMMlO+URBlpM57UW4KBu+JNfLlAd55waKUqStpg2zMlvNGjZtdjgkxJ
Qo+klZenlFfVBfk0TJHw6WTlv391Fo6dzdUGtN9y2Xa4EhKVu8N4GGT/0zCmLIAr
JpmmEiWLKCjBS9RF7Do3HWlFJhJPU23HHilsUv3PeLedjQCW0tHH1MSur1eFFiDE
VoMly1N9AoPdZwFhJGCpBolByrckXrABFhJVJxAmGSXbMR0jzaLa0nIc0jiSkUBt
pVrpe3nAFAn9lbq8sCdpBy/c6Vdo/z+fR4ww0p44ZBbUq/iuq7VOfK9akT1J2KVX
tLryW8pHk4+UPmI49Enp3RR/5YOlxrzl5KB/4zBAlowCYSbXhck8/mkoWSrziLPO
iqsAiQJvVVQjzDNQOdYtDCn/qCWnlnp6Hb/M6rVQlRsMjhAizBPthOemGgggLDi2
47LMKwAb+mRhJdwE4hQ+4cOFS384V/yBI+ZCoLFDv5SZxFRcpgtKXh7mc8lXAtf0
RNdpg/8H1SykeyoHILKlWiTiNbXOUgjTLbyWqqyASXY8tVor8ogIlX6SFGdxud6H
HV+Sg0vKAvZVxGXnDjW6nuZr2ag095b/rI5PY72xWORTHip7jw/P7EWZeNefpvKN
ZKtinQHrpW8dFWw/erVifQQGXxnSKim/PCTanCRblOUd7UvzueXh6MgwGoWZ9q+B
TJIJaQVl0/m8hmmtAwhpKnGdy+1jXNF9IDP6flrsg1rhLrmw+1ck/ZBFV2YDllvn
imd6gWrq6oer+xAyL63JferF+0rg7OXmNI6qMYpw/PNRpbxeJKv5sg7Bit6ObOV6
C3nuuNMV3v53XJFKMFWdiSLMzip6hCtIHlyFfMey6Ke2wkWn9Wpuv+5KevqFdBKW
ODyc4D3UqjxoMGRQqjANNS3lAZKhM34tmUW6VQnM2vZsXDamVxUUjBwEE7Bk2byP
3PGnDtvMNvgk4qv0U8V1bnGGCBP/92XxJ84D1Hudpxhoha6DEullfvDbVE3LU5A5
AbNcyDVPdzvC9NHCDndTwFERd/CrJp+GdemTs3WpJjUQOs705/UUX/Jhx+khbEwt
uuwScSLaazLdNa+qbCjDraCa8xG2y0WnntsbZ4zD58S2N0F5mQpKBiqUskwjTc10
ZJqscRLfrrT+YTpge9DX9qgOZjPSG+os2cVsfEk9tHYcvrJcFaRvNMZnyTj+Ds+2
CPVrVTrMxJuvoH6cFIqiVXkEEwTS+FBcUUthbAcUkgV8Fnb1J0sXIdby7Nr7F0Ot
swBMXpgNE+JNTaO1HMQ4HxDsDTIYvHk40rZ5PhNi+c1g7KWd/mprWxf+UCTKmuTG
hXG4bRuX5MxjZzTaDDEYZQaVSOoAnbC7iJ+agYFZiq+F2z5Nmdrek8eOHjrOCjWO
H1wntfld9ugR0HTlEjzgMd3WdGAlpndgdhTm7es4/5xyPSdSr6RC7cWZe9d/GSls
OcON3zjoJy/9FArdFDg+k0RDZQouNXVvFWo/xnwg9WrDiXU5Y2G0RDIDRDCvzxU+
LVVx7IQ49bbehokPtGcDBzdhsPjBiB45fay+sH9jdJOXePXYRJ2T0G9udGqXZdyi
+nQ3LQ3Lgb76coJ70C+mytvwSG0JSg6wq7Qe+21wfJGNHTlXBcCRzPeqkRVdfPPa
HwhNJ7qnVC9yTaj4c/NeEBJusYiGlRtn8Xawq8Z80hOdQ7BDZdmvb3U4MYtvieiU
vn6QwACDjkKQD3d2/xIWNfo+717DVW35zcTrdr2f7aAxuP1j2XIA7ILy+hVJn0Fz
qjI1w5DfE5JPz+Ts9vvOZHiA1bJ3oIYkyu1umUmUUb+XUH4VcU3p94ULMu/F/+9G
7rme41Dw6cAQz9UnspaqQ1q+wtSGNvBumWWgc47wi3MtbyosuthVQQY1XjIJqBDA
8po1l2YU743fsn7yXYgB38fbUlV+WKgDS8mHMrJfHJ5K5C8GMpfilwWD1OC6exAV
R465XkWmF0PJgp9ld5Xk4K0W5Lako0G2jgV2JLzWV812dioCRztm3uZEC0utKSN4
E7yownmfJtWfft+cvqPIYxrhl+rhWTY9eEq02CZxCRczSKL+5gNnWA+K3h8M4Q8o
STfHoBFHm5knRvQzrhbL5npEDd730z8NCns/HfMkwj8AZm5nVp1g0G2uqcY2qP/g
4ILNU92WqzmiQBGX2pE8ZWDMeaM4/NFUpqI3Swtg8UX0DEDJc/2UGrzC8JJ0NRVZ
i4x4EZeCs0u70U83jEnosb/9afSBoQ2jX1gKfrDDcrFGNC27UicISQWOXeURyx4n
J2nIloSc3h8V2wKM5sLYhqhrUGnFahmdjEdUu7hr7h3iDyQs3mOsuedcwc8mN/iy
d4/FnlkbegeZHgUy+thXVWNcNUibONJCWodGsyyimhbzj+HEGURY+sI+xkF9asZq
+D/n9C7q6gFQawZVkINxvNW+6k3ZZmWTmCsqkCFBH7wi0kbOpbbLVnPj2OI6TPIj
OLC611GJjQ9CaZY+8xAZl0kQjmfxI6IXQDbyOsXtvtYITA0+oNaR67RaU6pg8Gbb
wqr+uJMnqexcITFPvqJo8jPiHT74YV6dRRX5aOSQQ99buF1Qpjflf39/vhKwoXHM
ViLG9E69/beNI33PHyCXKD1e6G7bwwmvCB/pn/8sgI1HVQyMFvnmEojjruUBkBMj
kdZSWrv2g77vKm1Yk0npoMkU04x/0I7pdEZabVLHR+NIJJh1E/CAnBVSoMNjsstl
EuXXQGb8L3DNgOvr5pwW+CZcjl61ER9jrPp2gtQtP8D8DmTzk5T+2qUbzEx92bPi
DDL43U+66LN7rvawLpfLx6TQURXrevxIXPqbg3l+SaxTNsSYMQI77/ni5D41cSwC
CL7IueL802uht/MMccZIhdiNrW3uE7v9YguZY1hl6qdUMsqmfcO8/aLmJCqj9kYc
p1MG+a7dS9CmChzHb873uBxn/2KXedakA2SHqWCpi9N8o4ZCdtH1d5UUkmT9f6fp
d3xfhYGHohxpNYfy3qAwX+PcskjHTz1Yv0uO1IrRBZnPZuRGQN/34JXdS4avQSPc
0McYmuF5KM4gfItyT5oo0RyR7Pd5k7tFCaUY9Xl2wQaCJ/3uZI7IrI8V/fYX8i68
pSatLrwBTjoIsE4fwVgSdDPxA1Gp7iJ384YH22N1dFYHAro1VfXlD+gVtcpaH9GK
/V7MvCKOw7MAx4h9FGUhhzQFFbNjsJV3Lglli35QCgG6t2KwQLASZS8aHBzFMu5/
uKkZo+YD5ib4Hbskcrs2pd9jEUNDaZCZrkWQX8r7C6QaCwEXoJk8ZnozgKm+RIL5
WOg+bIzTsHiB9BebYXA6m9HXzZGX82SMHAoqBBOHFoTeLB5S3AMrcKvGjQzL6pVX
ppdpu8ohE+TeiUHxF/KGgKh+92CsHflil72AS+vyRsWTQgi5m8y1/F/brmqNHFMT
1fYpq2Il1Wpji6idL/K/xx4kXLdOo+UTq3ljwcKwHXmcqwfo51BivlT4qehEuODm
WC7XZIQDba7pEDHVnkuiUy6JmnApct3CGtuCU/SiEkOxdjjR8OA+ixAoU7hpEiPn
RO7FhTIxcPDKrjkMy2bMyH6LNEX0AvQqSrJj5fHs/PrAeoP6RFvUudHf0c9JsUrH
64qIdeb2NEyVsUTaT6jPkY4aVgOmIoJQFpuZBaaDnWQZ71NU+H6vmj2gnC6YQdBf
tGwiW//DNBEGnFdu/5i2ANpoA16W7DelMYL2aQuEEIbMfNpltx0oSpkaXFV/1N5e
+hosf3hIOJMDhAAeO1eNNg60K8vDfeBBjNNiMlqlWjXBQLhn+PyOZGkLtczXksHA
Mgo0EFFA4YvqXEWta1+sdw1bMdkG7JXcJWvM7EEXcAMv2dNtKW+Y3NNwcde//9MZ
ERi+LT4SWM0KD4aJx9F6ZpOpWCkbBocREVWCrHtChSlGKExql1nJ+295+uvt+pa6
V0VgALCYI8Ij1RV9IxWNnpxu/29mLOQs8ZdjpANSbua/TzE8/9ZbSa5LAStteSYr
YACY33B4JIFhoWusKgXcRtBX3S9FKOm+nTiCHao4CzLQYZgVVVFXIisnogkNUG9v
1yYGZZ3Vmk72rUURFl0/jbQRmRPO8GCCKzRPHhc5MPJmbDeABKyjLSt5dpOsd7R3
hRWbZcwEUFoDbL3AT1YmzeSU6MXRA20QbKC2Yy3zG0BkNYPjUTpUMBnafvbRx9Aj
C5bndjdaIkK2z302f/VPYzlr9z/p3zhgqBn+qUrG1lMGCHWsZeQxtSoSq2EC58//
6tjEVFynH9u3HmKH22agQSVUwZbq56QTwtnX/MCHDNK12nMLffX9WmR1TIRTwran
xJ1kiFeT7b6hQ/YSNFXBCl0aTMptN3nCDu6IDr2PE7gPO09A4dUx3XJhqadzCjc9
mzprwAzWYd6gGcfRwkZ0ANhsT4KUgQc+oogzJ5FEka31Oh3Rvw5tfe3ieMNwUP8G
PbXImdI0NMVLwXGPFGod1iPJFwuv8acZ4BqjSUNWgLHnG5TxFxN6Px10z7UdIyRU
RGKzb+5tfijqx8WnMJYrowo03MUSj+Ykebgk2gXMG0cAtuO6kdthxWSjlv9YROqd
w6lo4V9FZGRkBPHPaJzZnpI2CB4YJd0KQnq+sPT690o2eLhs7+FU6s19f61nh485
i60rFqenAGYqe+WftmImq0seMZP8nZrMq1QGCCCx88uuLsg4A8C/Tm09Vtmapp71
sKUYLxobX9tqlgUQDVO3/pa9r7UrMNDFBjoUeCxjGqKiEN/hgPEyYf5yi0pwyXh/
PqjjaaCOIJweWtV0KPVceYxvS7qhkfnuEY20ySAvdfVnbv4lwnq+v/dlwq/kdW9I
Zq2BbqxOyQu3Zihx7oDYu9hEkRBVdxOZ3o2IQoAfn/MvJV5GifilTkwBCZz1midM
qk9kHqe/27vhLoG446uBpS2T/dNWt4CpthDcatx6oqgqEbu9H8ckpEo4+Fgv56uH
8Fi0ADcplC8+f/Z3Rzvv7QegjrzgVO73awIdWOvs63HBu1W4lVQ43OT56Oa4QsKY
Zw8HeSWImVg0sCZE1RR4MqMkHswtSCJ96/oHqHhIXJwD5cgrOqIFUoJWwfXNohw2
dBFJ/PUVpfkqi1ib+7cONfrfuTXZ6B8Kg8DdFS112NfnrqC6ZVdkC+9nuWnC2PdY
+4i/XivlwVIZtMBTl4vHADY4tobpskEaF0gqaALEYPwXL6YaYG247UanDV6/Eb1Z
LRQwvl68QUJKgnyxmLEKgn7InmdsUQMFLb70kHUzTEYehcVRSYcBU4vjmLw1tZju
H9UDVbMq22XPs02Szug75s3yv68UebJpUzTWTcBhKAsfLXcV+0i6+Ba2jdEEnwNX
u+RfRg2iepencXELIvl3PtGlR0nu5qh3ErilL4qrxhvgexxqCkGvE16j6B2c5rc6
M4oAym+/AZN3UoQAPvl3r6iNlMmp+7YjWT/ANlVByoRVVNC4J91hohRRK096DJhm
D/UpoiqxrBKGYLMh7b7t5Ud4fU8NKSH8Okvbhaw4DBUQW0JWWFclt74PM920kopH
m4VDPciRIuBHl6LOHPP2X+k891VC/3T2GuQPAdHFY553b1G6kQsPreI9K4JCYZlZ
lIsZHzWLPCMT9wUPWYj+eOQLiEV/lfZSipnJR0R6wfJDw/nsbN1x1pB+ECNt4exQ
2UAL2NIsaDgGYup/LTqyy6tlySyKaoqE9Q+ArfYG92EfFpX3e1ewA4xkphbMOC2K
R8fEfebFC7ycuujUy8pujn2qdq3AkpH9/fKd/q7VWCa3tiX42Gw9jIeu99nzSYzS
70saafCgX6Sk/NEAv2+sU94ExubRKk7vHhOxCmgOC1xvypAcjGhpLJ/mgdDKphDp
x58yivTxsemfETAwTTXVEIhSAxVncUZuoQoFhTeja4aQSlpFTxyzvg4D8qvSMIcs
1+vUQc69NvWCxfDlcdIPsMycJ8DfR7ZY+h7bzbPgftKuVdDcAgNN05BY01OtWmUL
mqFFEvAakyU8wpMwt91TsG+wwk2yTzxMUPe7DpbokxR6ygXuIng+Thmciq4D5S9Q
risRZSpxfNgxu2aPh0m9LtDq7pC1KRuLFgLSXvdVW8yBipGfK67NA5Yl0a9QNA/F
kCQHHb1nZEB1CQj/lPMyCE6vFhTLCPEDXZr6kVcYdXOji8F8UPWovXhs2LZqomGW
boKWMbn1x57qIOXbSmU08Py86SsZ/spy8/7Qo8JNfiAAYwYAh7NjhlYZt18/Hwab
+Xo9M4wOebsa98wxXJNNG9cOpdCJBsA7WBhizSjqf/ATthpjZpGVwgBIXDGVFuq0
RQzEpxq6KGaJu6NBs2fCvU7CaqfaGnt46oRWnzyORjgIDVcS+JguR23OcmxZL2Pw
RwL5q5UbXbGh/pwG/IgR4uowFMOjzTNZqkf0yJTyST0qRRR9rr5mkLn6nwkwlkqg
hqEjcrL3466L0i1EwAGdMsenJhzVx0VFA9Xq455qGr3TkPwvMG1p1ThCBHzoCgU1
WiO+7SVgQlSM4YCLF6ptqAX4MYABC6EnS+LiGmCHgnsaFQSAOa/yfiDVwedUBSI+
Q2P2M2TazZkLzAFtVE1OP1xY0uJd6+K/BLkc9EFk9o3ktjFHNbe8z13kbqtJ9ue2
5dF63QFB9y0fhoim1B0ns1GEM+k7+1skbDaHRaCWgk34qGS0duAzYZmJaUz+i0r6
/aJYi1TX1Gp9nWXWeejKxj4fFCpUbPrE7jsZ1beCF9JWCFyhJtK/SE/E+mrqleCd
HXqaUja2ISJif/hMJOeKxMshJ3eIFcDqStzImj+OmoipAGxFGsU7HVkNqB7jWp0g
TKEL4KkHXgwtrZg3lmPItGH8wLIUWtXimJs4Lgs8NDSyBWuOOEAYgOjvYebFUnOG
QvkYPna5QTf3EAlKtSCDvd9QomZA5I7uDNZmy9CnYHfisFVUuPupIFeutKpEh+Xi
ZmPn1F7S80PNVTVoQuZi0/EGGbAzv9kUnzdUrhm5Ljs69lXbNyJQtO3V2y7DbDCT
8Ml92h/vfoVwUhyyEyyrHDFbHOtYSRGBQlViWjAlcfrTF3MQwufn1mjFy3nychkg
zAkp6tvxksJCw7tQgyx+lCtgyWRjzq5O4SGoizT9s2m49Vtax6hRfjUWPWzsUxuv
dEdZ5lpx3pgjZ9nLyclnKKxCyYKohn/0soGvwHRzLSUeiylA+TSpPLtcP46xksvh
sIbqbU06vFFyDc0tVkmK3TqvuVLyWaNZRKbaXBzD7U1s/mDd9k8oYoUW1qL2CqkE
uTNduikQbPC76tPYEfI9B0T4LKxQJXrKBAUKPxRqiyPivwGOWWD+R7ko9AyqJf8l
ebuTwUlZeQHQdEfHpG/Z60I6N7UroDhYJJN3DYyUDwMcmLLOUi7bHxiJsAi2wqIk
n71LkaAgGsTGV0cmNQkBAzORJ6jXLo0b9ZsuSbjo2y9w3ETFrVRc51vYfvvNW26q
sIGm4I0c47Ku23zJB/NGTxh9YgDFYH1wcoO95c3PRU+L+creFeQXc0DQeCWisxlF
EDsuJ29nMaTgND2I825aDmIgD2yOi8lo7TiG+0rZx7+bKq/MEheb4GAO6mk3mkdj
HM0dEe9G3/5r/iEBBB0tasaN1t95hfWBtXpeDjBfUArxBZwZ4cTClORsxoDWDvIn
S8Jih5IJE3cEjvlucz5JXW5DCjrJj5WFZbaDHcNQe1geqB3By7Gs2tU/NLY6TcD4
QqVyT2Yy84vPdjAoypEDNnQnc3qZrhATRXQ7Ds94DEdoj7SUTp3IEIVdO6WPfG4o
XkBuS6hCu5unRm2ATYTwpo/tZ4SIDom22gVa/JItwlQoIeGjWYI61+jPjBX2ehix
q+6/2NK2YHJh8q8FTu0zS/c1deajS9tBpS2ThzwRH4jehtXZ0icWsJVcB0FxvxUS
2MVUETFWE70EC1hwuYqYNGEMvhd/6mb0VZTRsfNC471+CpuDz21LoPbZ0PX4pcpz
dHLIxzG8tOPn0PeS/HbohZHL0UEqyCEH1gb3e+QWP7KDsfW+Z5R33UgFYsFck4gz
A8UcCpjoKNv7zpO0CK/dRpxg+1QikO0YLRWUe9BLbl7l2+nUDq6Qc65tHMcvxvab
LLOFEn/la5KMuoXI6E894kUNv3hYzwJFfupXXY8G9L7XhTZUBnLt7KPLDdU3EyYs
mcUl59Czz9fpOMCBGds7zNI8AZPzQdVrqdGHoZJvhE7B/nm5tkNNbVIyhSytheqE
RwVyntfRsrbArNGNVH9zNnyFVpZuCw0pjqbSRgCRMvspjWoyAZFFOeMnzZ931gAH
DaDe+sIrLGEjM9fNDAlwUdX3mm5FMcK+BQKtGltPxAK/m4cRniMy6FOS7A6tGpCB
KNYHvnWPyYDgY1KfACGtJYheUdVOB41Rs0ArJTMn2H1d1yDf6mggPQEu+UK0GeGV
IKvqpY71Bv5UkEudZxntUjSFaNMp99Xbaiz+P7nUrcdMo5dOIz2o9x2Dc3ujxo06
JgY1g54t/6GSy23e9z+ALkaoDHv74QgWhYBKikdxqfABcw8+tN9VhvOOwfdJALtw
yeud4lAzo6HqORtIAL01zEpzsYLGl1iDnITdon/q+KVdy1wL+JUffwonV8IpsBqP
ViVTc8UsAZ+DnCRCdZ2FZSz0Bh4uC3m1FYWEitTIzAZqZkgdDHYWUqPd8Ft5jzic
Jba9NWsXGJIfRTDBX8ZH2OIztZX3DwQAJYG772bC5Jl7sHyk9T2b340iBTOIpW0U
77Fv4eohDdWa0S7LWUJ5IHlhfjWsUB98cXe9+nHJ5rqKbDMNXwjABaAjU1u6v/LY
sHPlKU3/FR+8eT/3qdrg3g1Thu2VkNYgkfIkIGrO1ILeoVS+wKmQCaGzKO6Imjuu
tcsOWckqvB/CFEI0dh285BufqT1crXGI1om/eaadsPLiWUxUIJag3i3rHlLxIjxv
m8Oob+5Q8hYRu5oQ1CH3qGcgR39GRJtzLmy5IlcLLVBcgaI7rwO8MjACBn3aXXhD
QqtpQvygpx4TXAzQhuXtxhYFc42uUiAQp12Ep2ZTe1dN+PDP7jF9Xf3k2cFLfYD/
l0gsdSLtKJ9tbMCtn52H9g3X2N9IaUcUIagqBE7GM62NF3pDpJWvx7iUVru7K11k
bRpljxgTV8Et8bRJLJWlFb4cCxwOctniB6XQBpkPMOV+fKpz09UbwffcLfqJh9HL
H33qQqcHgh7xEbbBGi4NGQJnC4fuCaDI0k3fCvh9RL17zq35hCT65pyS59g/c3VT
uYI+GGAXqQq+U5rVqlTlEWoFEQiJK5bMW3r8jAanzDiHe86t1H3DgSV9WFuI8Mt4
or3lfPrKLLTuPfHMY9M6mfuiO2OIoe7qwac3dIrVnotLnK/f5rHoS9+FznIlWVpp
XUHCx40WOYsKscpWkhtneyJXWfojOVa+9HCnjCVCETzwepvIv9QL2XM1GnONlClF
gbLT1dwf8ddhCyAu8p89M9M9ZiKVTi0X6YZaCMSrYBq8kaJjAhWJR/TkFgxfn96l
uMTDH2Y2shJmCXKaLrEb1uJ1jcEDkRl1Rgvt1kMNC/KK4rYwfB4FTOy0Ovwh/vE8
IFkIrTCRx+NRPFuFuLW2UEftXWfNas3n55RAhnMNAMUWBfIxdtBJ+9mtR2xTAlbh
xhQze4JXqUSZo3OSrmdb/MJWwbraIFlI2d5vUSmXVMW7CBPB82MXF14uv8/fVEhx
PZdXus+TURMX2cd0Is3hjN7gZ/Nx67yNmHhozIzwMO6FLcUu8EYrliAfxPCnP9qI
0iNB4QQK7PGrfeUu3SoYjLrFwMD2l4zBxW2irpmmxTsi/0mnCF9lhfa4aQf/VPKp
K9mAihUTVbKtUo8g0CyAGqiSuWyh3kmYC4w3YXgDtTf524Gb3wrG1jZKmLEYzMb+
APHFvCENS2qJuUJClnWX19J311sm6N/aTFGrebbNFxYeGKttjOtzTDFbGQlznvtU
3ULRTTYIUq+pjjsSoYrhps1qRaSpw/8tq6nVeunTr+xb8pQmgfBwlhutL8H29y3w
KNs3OAkAsbStPsqbJJ0RCH/svH1lDO36tajVIpN0ccvmsP+P8VnvzUpCpCI7fjNW
hqe0AUmHOOCEh7EYh9Yo4M8NGomA3ue85uGxv4BDpKsV7wuFcO5mbjSJNdfzp9/B
Ws4W/cLWDTzM9+Im5YUEQaXPkj6/a1MSYOgu+Gf16QYRBgJIsa7Rw7LcDT1m6hnz
ECJQ/jKEmD2gdovTFWbvw4AMcaF/7dfs8cKP5Sh31eSMQpmcvNuwT2qr/VMIW/5n
t0sqH/AkzLzvvb4PUmXQN72HI2Juc7zT81lWhweueqK2zMD7VWyrSfzM73FnWNAX
+A++IPa5+crJypZNRCM4vwP/SswACia7SiPoNBmcarqJzioWOk51Kf5l+cXANVil
auyLQddl9LLj8XDfs+6ErRP3E3pXi3xoJkxAcg4Oy2/FGCILlHg/aNiUogRY+gMQ
D0Yk0CzbjRz+mWJTRuqISAK+mnYdK9S1F8XZgsJEM0Q7xE7rQMc7il15MNI0kJb1
IwA8WRb7aRQY0G1RBhxE9aBnnTnCu5dZ/L9EOQrOmCiUe7jvBimMT6PhgOE6oyeK
wcaMG6q+BkkWFZQgyA4Xf8mRjW12KWNxmFIbYPlfik19w1czG750ItY4XTBtLJZS
Wr0x0rk/T/O8a0TmQyfjgIzeszMe4r5oftsN5O/CJGu4aKBAAmhhG0ruNT6UaWyo
ZAv0IunrQSvV39hkDF8Oq4LgzJC0Cpe37C9MG0lR+ze95GNwaWN9ibdAkFrotvYn
l/kdgchn2rNkccab3ptwmXng0/qQBe+ae+h5GFH3b4xn+3tih5cXCSzxyuIF6eLl
4iB9Xf0WYIoA7s/VmbVGkg4bgbVRzqvze+kFfyyW4IrZ/XAHpcQ/PJJ4cEalTI0N
1nJFO73B3auKQUrluDxe6bAfG8ung92Vwrbo0ixFJffCEdhi/SVAxoLrMMqPJDuV
/sh1yw2lZySvt7LEduNKaLgaSgj+O6skRjd21okbtOUbVn2sO7yOnkFIrlfAXD24
wOOt8sojfbd8N3e6P3IBOqT8e0zh9MVVNvfSLWegQMsSEeL/qdb+rayUuBedOd8b
/+pKLBmhQiJy/6VyE9tWZjZuFXQ0syqr9b61qmh7ApIhEJ7Uyh5Fo2X1UibpVwmr
x2wq4Qy1v45WyYxyBcP6qdfoAYbwaIoJQ0wMOoFcNrzvI24CYSkgMtA2glgsFbUT
K2rsom8ufbTHiem7vV3xGma/Mm6x0ldYJaaK3fm3FhLuo9IOUDaC1r5w0d9etIWX
2iUcTyQ4Ut+sGiwh4So4sr4QlXzE0llRBq7uximuxEtBR4pHHjlrbdPyawqU1BzU
bpUP3LQmd0aNKbJQ7xE05GAzyZf1P7j/sScUGjHVj8uTpVxGhks02j9E1129ccnP
NS6gbB9RmhGneAauq/TyMSi2OBkSZFa46z0yg36Ef+SM9it0HbA60W9KqQDr7KWW
7kdwkdNif/6jk5vjvzVjKfYX4sqYqs8lR7b5IosRgOGgUvd7TMko7HDdjJ/kV4+X
6SKjgium5BNy7QHcADubQRBm1jOP+1JbJtKP/13rxXTeVVoHLnO5Z0FfM02LHXOw
Mk8uPcGAC6SrQ/22lmqzjT9653LbWu6eKwhUKbAgA/eRcL84hd//h05pn9teoFU1
TpI63YetXjC6IoUHFf276it2b0qMPQCGzvDsQbgKDUD1D0yceNR3SrutYRm0ai6v
6+fJU2i+/9EuEvaim18Gn6Uo3pWrCwXN2Xeg7q1BNt5UBGJbU2smFbNeIYf8P773
TGG7HlVIKWEokII5n+p4tYrrBsfj8tUuw0oHmM7K+vWve9FnLDRIQl8BhVhe4Siu
YDHJDIgA5fp45sjc3guSsu02Jfr8UBVu4p/2iggT0kvh+nIVulb41+srrjjN04C9
hu8Sp4wEy4JLa1XeMujLU13KtciA1DyfhbkiYzATVdqIHD39dXNXaXQ6byREr9Sz
7fftYlYRhPTJLR8TWLqZvV+KqvjgeQqgDQuorTTrXO3LXqvjHYu8kPV1b+41cHRU
t9bWRALHJQgqLzMOsaUAnu/Y+zHn9kcLMoMeWALee89pgA+9Drczm+rGYHtigWGG
CGhSVenAhk+/Gr0/PfG+okG7cdJXx4NoLvA86LsKLAchS93xlgeFzklFr6l+z/0N
ZRYGRO2n3Og+mDm7OZr7BY8LfuYUxt9hEj26RJ6fPp0lFnX2EmO69Yy3idfuxlAY
HC+Rm0ilT3+w7WRQgjpb10j9IwNdv7gBtPwAF9Nn4EWjVQpeVjRjrATxDmsaZLCF
2OLARYIM77xb+OcPW3nZV366NWIEcxG46kLzfYg60OZKKz6Dp3FNYNUqa4CIZR5n
7O/BXCjNRopQU/PKEA5U3LNDBgzWC3m3eKY7hUFFsZJg3729rrQCh2Gmz1sqw6au
06KsLjn8jCwP6oHYtWrOYGdR6gTahFAn/DYocDTBLAp6gkQnlEAFwUzRd3LYXhiR
7Bm8gvTeqw5xScpYb25X6nkdWeTPd+wiJ03k4YSjBABcjJCQrrWRu6m/nQNYaikf
b/Pvty1ULBNibD7QBp6LAh6Z7Oam9lzEi/zbzQNqnwIoRejtKtodhoDPsNEzWc2n
AqZJqNSt03YcoPsxIMRIvdp8i5yfMDQQjrhcNKSc/MBwDfGytPCI9asWu18dT0cV
dpCnwcgQyMCcVEB6mvDot4Y3e1vv1hbsBnk0p2pHRUh8dq9kvcezNyQkW7IlD81C
pEUxy43NEbD5jjgVdu7J07Z0mV3k/2lx5xTgC8JjwDQJNYGj9+UDE/FU92bHDNRU
iFA8nSt0lO9u5paH+m7+74OsB+C45HGu39GE09lZYfTRST3NUIFQYCfRcMMON1OZ
vRZHwY4nmsvnovMwWohgOOfOMOV9Xgvw2L99aQy1zsiR4yJF4cRLqFtI0T/DuUNX
JoWTpRdgTMbTVZIQbeSyQrucu2h702pvoy/udhVq1FiIsxyU6LWy4O+Wh9HhjUDY
GUOohMWYeIYbC7nxGhoeRnFH8D2uoehG8RxD7QthKdSGPxyNkkxlBu0UeA4S4lY5
HwEjBG/YOHe/cDkq/QrcDmsXdpq2fHyrq1eXPVdXVVQg7oRirJGpsmcSnbl5x51G
wu1FCOjCJeRPFPI3BsDJR6EKIka12E0qAfB5YS9HKtRsi/7RYR4o7gCI6erGhOtn
H3bwM0NrJwZbPq3HNOhxQ7HW3BXUEVrgvQdMMtm+Nmdli5vYNKtglsSfqrxwi4AB
pwntnY/3BiG9+XFIiwETKwb6wS2EfzuEBpMjB5/dIN3edB66vNAgjzw/YacdR3K0
VpKrh+G5XI/7hldEnemDgQSngflGvFrLCRC7SunWTXHKV5ZlqNt2cz5QM4ko0qEx
gdtGlwqTXbVqisE39hLhYEHWsflvuqpxB2orkV+Hzlri2Mat6EDTzCu0txdH9veb
FHI7DU5ko36T0CdDN3YIlWruLjOo49TzviYVPm7mogT9tGgfepIiQ7+XcbLwCtji
9/+yBgSC/tzzKnJb5KufcCbdEvikOddpuEJfuwN3SKnHPgI0oG5W6nlkQ07LFN03
xEGpW+ZiM0zpr+Vbb2V9lNzIBJS9f4VpbU2LbEMDkT3xma1vnV5kvMOFcj6S1xAO
1yvxGI7mxPrRVTzhsSuo+Fl7548Fdomq9XS8w/LeBJD1YqxeMR527V2pce4Ca98v
qkO+ecvp3YssJN414sRVIi1G+AbIPk3TDaefeXIzL8UnbCVqER5lUMSuYgQfxE1M
U3qeQ6P91y4zol2lb2zOAgoSSwp5WaB612xPgg8K4doyghFLKhZYnnw64HHrmv4r
4LWn4+tL0jgPPtchnVotOpZRw3n/ufKy1BQ/VJc9gdVmzDhTLehSQJ9Gnq0QUkFl
BywkhcV/FFPEAVyfgB7Q/YW2EDXimIYtWGg/kqkWWBQICfI8IFUUBKLSUD1Hdl9m
BRUNAMi3wK35wMdktdTRela4cPsk51L1rgxUBXLTZ4CTkXI87+Y/G8peNM3RlWLR
Mne130elwBA48z7ZiPCpTu5ymuaERqE2958bjSBC+gd6pR1Z+Ack2lVLJ2m0fEQB
FSif5VsMSIQJSY0VK0ZkxXYSV+MeeAHvXsde5O2qygs/AeBJH0VFRl+4eS3Kb/7T
T6Nd5Rc8coH78QZDZfxr2qDYwQ1z5DYh9asuLsWYyaeBQHo6u1lAQH4mgmZl7yZZ
1vmKSn6sveQOacmrZmNPssXffzJWz2pX++xsySrWNwdsdz8D05F2wrn72lDCTNf6
GWIqLWFTVr4mtMox4WQfTmGNadjlJkDJRmf/xZGoawYC0sLQzzglDtL0cPM1rbnQ
oDK+1IWocRAeUt0zklguTlpsSRLBzRXcwnqtuxZvzEjqOGJNP3K4DXx1v3L351pd
MJojpSUD0dIJg2Yjk1L7LYLQMfT6KyFuWpeXO1lthykejjzxWukNMo66E8JwsVgS
wl69vhz5lMFOCvaaCjjaSu6Stw7Qzbm6e9em+F8hcSXkpbJpgTpDB8TD+UwcZol8
LXIsqkQJcS7pETc6aaYQrwbRierCT40EmII2yAtes/ilJ4Bm1xT2yq30Ixxw8J6m
hB0kNPASPmIO+omqk7bzGq5AYWqsf+IdMLl+WeEadArDTHN+ACpMJnIDczRPPOhx
RKHN3j5PJI3r2DufE2CIDddGfSkxvgdPUs1fD69+VoSXRkgLAe58H/KFFMvoBbjr
IqbJwVb1N5RSiBV0MNC86iRcdogpl0J/0NcpKqJVAO1G46whxg7Ni7FzrQLwwTSO
+qZBP3+tjvSOBUtNym8kA7TcE60n3DqHp67AvtE+Uhd9Cl7t8rahfvUSGELMXfrV
ffXkkFgusCJMwfaTxNG74stv/MJrm6p2Ax5YzOCmTdLyHHRxsooqcvfAHtl4qOxv
xtna1be2HhwC83FhODsdSNdvhHAZ/1VzspyQ9HfGObg3Pno8QpRJhWdg8lNlp8wJ
7RngKq7LL1q2Apd0yzuI3pKmJIli67iw5g8jHDCcbhz4SQdfadP+lOwrYYbDtaeI
hHbHzPgME1o4MAmqvwO3qepuMWFil/yk62Vb7JdrHIvVL+IXGrQwrrZi2ZJTtdBx
E8b3DuV3Ys1ZpxQkZEEKx+dOujY1i9rWj38zPVaFRB0jR8z9ccPvWdVQNxWTt9JG
y2EkV/uvocpjiUE7abOcuQ1dKkl95QfORnGPiQiawMPtnX+Gin/uczLx/CkiirlH
plt70tcAT6rGBjXMlqfmJGfyWJNtYJ8DsdO1tfXmcf/2NeY0gOmNzgEgQMLB345R
nvfZeG4mZDwF/Y9GILsVyp2+T9P1tW9il/JuhF+rSgVYkZJfELF8IeguApko6CY0
iu0eD0Fz4cMhmD0ZVy+RR4bbqy73b9RBH+4cCvAKfzuiufocTvMcBFWvz7cfD3cn
coP42XdU0PczpwUFJxzlGZNFv4iSmygUXp0nHGfBXljXSHBHq900da0oUSJrxcsS
M5yTtNJf5YmdqeVNi0o2aUuo6X57pJk0x1x2CkCtt4pMCiwvTDppb5xzJFoXwa65
2FcHSFH78/PeFIILRkMQkaE2wci6BdMg2cZaWEGMCcNlXzg6yb6PxNmQqPaSxRjx
K4aMezrlNNJUAklm7Bm9pTPyLJLro14TyskpzfVW8bTEnmLHyZ9gxZMGf0sCZc3E
gQ3RmP7W/naAsoc0IQfD5F67bSXBOpHnWe2bXSX1Ru11BMW4BTjftz7ObqX4fEUD
GwgGT2ril3hQDh5Ei4jYcV/TAyFAu3o99jYgppOCKf1+W1bP07G6fDGcVutOdNxz
pAoWPsxiPbnzYa9z0SffxTXY4VS5x5m52EfYNkpeAksOR4WA319fcEqxk2n/uBSZ
XY4KvimGm//ccHhoqFV9PrVUwwNxuAU8kSVfsLPwWZM69Gy91dunrkiDp4qmAhkQ
j3zJaQw2D1kj4WS18P41RYI3W2m3Waf7VI2I64vOBUWu669hmZHrEuV09lpxSDoR
su6TLbTURWhcLmgzZ6c9Z4d4qRs2lUv76MCSZ6N7GQtCe+M2/A+5+ckTsq610j4V
9Of2jW+NRkzp06NJNAnJu1CwHIugO6r/cfeyHefqpErDAFp6O8Dk3761njc+fRi7
dT/MLM857zDsX18goVJ0VeNMyVRiDDj9dCVP6/tQ5bFGfcnulsKaM+BXsWQdQFHq
T780f2ZkZrfPeAKTtqdruH8B9WAVUNeM9Hglu88io2LNqHO0BtdsHPWC7NFrUsBf
q2bhYJB50Z+rsroBDGkLgLaUzKIPPK7czbeyIbOQtQd3oJ/Gq3AR2UQVrqf5YsjI
iCXy1Jfz+qdCvttl+lClcfmGZhjn/4yvKifQtLywRQUl38Cimm5dBiyW4ma88272
05GC7zYZ+xfLvJ/4grSid0pIA2CEUaHVrGJGkfNG3iHjakjBIVRNYoGlspjQarw9
DJ3MIPYWr4WEuL9+lLDiSIQ2ljtMkoOKiggWPuSSSxgMDRYvcMMgDAlLJgBB64eT
0gS4dcsnnJGn7gf1PyLCFoLN+M5NkRjWo257SlUvFbtvw1fY0u50Z4lbxrTOLMOc
z673r2IKg+d/KZagauNwPD3E5VIEJuOqTQzgdtd+PhNcDXY206ouoLZ6gGU5czGm
q8/AHmJBz1F5ALgPOSgYADr/4AaKh6WhJV0vfLNUQeAJczzj8/TAHSTdyfIAuXBs
eCeMIsJMRkFj+d0kvxdbAP0+hrFM0IcJy1hmshlgRHE3UfHbL2AbWQIDYXFwjGOK
T62HBlhHV3ti/BG2Ui109DFeUhGpHsSLVN/P2NNefX2u0zqTOt5TN2fDcxR2Nm+T
7HBQjiJxx4Pv+ml5AyHoco3SSS+/O+kK02qnviVt+7YgjZd3prZTwE2fxZELHumJ
NmI4SvzulhO0d5RuSH8D96K39A+UaFztZ9eXnan5KYqbJiyexbQ8XrD9J45MPR2+
g/8s4fH7niI2rLDMv0MVaeq6L0NCeU2YA9XWydFhPX0yOxwS4G/1k10wXfuQBeJU
Syt2UW61KY8mYXLT6PUfQboH9/KFC4x/SMdzSyQ7ePqhz1CV2e5z2dt/v25uEq8W
VFJVl4kRT8tZVsZHRYIN2soE6HD3SezWtj4gjZ9+MIEz6F+f8QL2Kwd2MnJebMit
8Yq5CB1ngo/AnuW+VDyykPJ5ZFLztbO9ql70LS5E8XBJ85jWnCF68xtiKpWTcVTt
14mTWiEbJOdZcYYwFaknQAEW+ZZYcdGqzl+KKCjYxAKY5Bl+GF8hAt7nUciXLygw
NJm0yzEe2H/A/aczhIVB4B3ZXrqHzaq4ajsklHAIrjAUCluXmAI3aA2uA3teLwlK
7uHIY5/o4LXFC+DXRoiFq7QZU+XmUMf5CfEiT/APTTzzLuv711kNNvdy07cFApxm
EFKddA4K6H9swbU1+RuT7nts7LRcdDIzzj8wFSbmm7RPYDL6Gm9GkFmPMT9Hs7ec
lMPxddPboBID06KzQdhsn9W/Nqg78v9Kq9YkUjX9FvSurBA/m6SCWrA+VwDiRbxq
wyHCBxKDDB8B+pdzTXLx9SOsu2zzqw4Cwyyh7qBmPnCmyHvUWSv9HZgqYbDiVTRC
vZxphcGIUa8p7jd1QSDc+gmNlI8IEVNUdKM4rNN18sGZ2bOHMmHcS/FStv3RtvYy
jEOrhK7wUYeC4o4QfPMpG4wWfu0UC4A/nd6gvZdGbA+gnWbeGKS274fyUUKT9d1j
oNHi70IwyAPEQ6eQINergEGpj8sOoK2PiwGFyydo/mnb9nxESmtHHfhOf39yRr2s
dKIijxd/Eq7v9H62oxM1i+IaTa08zr5EonrM77b8HlY0TGQLLIe0wbV3z77zsdkv
F4x9cUAt3kS626uPv0uLtDrNdxhVsXF0R7Y83fpt3H+smahJ7+YyWYRu5b6nKPYV
yN/bj0/opR04C+pXdfIfMZWNPnuqj383TjIAdIWSBQHuthEtaN2KbvBKsZU23Pit
sVpkC+3PZ2HXawaUivnvSop2nDoFtqDPcXLTDj9y2RFDAf3qf2nNVf1etMb02Bwu
0yjPO9lOpEUdsw5v8AtuoSNi9LOWriPiI8rXAkAx8BL5EHl7nij0io+GI4jK7DB1
LkUSQw6rG1C40pSrobAeUf0EI9Sr6MRtfgsu6qWNoM3U8X4g2mk6uKiPjEOKa/iT
j5aJriTkNl4W32wwUYsfbeuKZdhEG6tyxVbUlHYrn5tSeLlVostjT1r9LvkFbMWK
0uz9rmo+rcGzTd+A06oDYUj/xagKQ48PgWf/xGEmzEuloVKcjmHG/F//HXQYFvfB
itIrmd+AgsOFI5n5BAsZTO+J+D+Enecrp0UhixSm/Y9KnbbYWdbnqa3HvXK3F4us
vbRbshAlPJY3F1+3NyCvc5yObwndS3O1+WcKZeraGXYIQq8eWKoGz8zhhvrmCAp2
fk5rihBV7euRLiE59CRk4pcp7maMGdh/xd5oP/n70ysUcfDga4QntP/ystkmydsA
WViidl+LfLUeJ2bjrQ1dmhXEEoAJlU+yVSBWT8Z3a8MlkaNgqRAjfqzALhpznOen
x6Kh/aV1BkLikXBbXBQWPbniapfGHAOrv0Kim2cfRwi4sQ7AZ6EcDKeiFf0SAzA9
tF8qXwAohEqHyEtIFMih/83bDAb1IE09qrvrAjeaYbQsFfhdZhikXdzTPLKLWQxe
hkphk7/NwONx8Qjd/G5BiJKcvHhZ2qd1BEOLmXIff3RgEfdsokGmguIaLH5VG83Q
OZMBY7WdWVqc6rXEEcntbAz4eMvNRQcTzwv1Hhl8aGOMRqtPhzED0bvgPluAzeCE
b8k4xp6VeKZmK6TfbzKpJLccOmjKTenqoAWAFe1zDokVM9oBYtuufkopevepN+8a
V7UHPzB71Gl/shfBq1HcDy4LGgPG0IorgDIKDojmuRC541x/vK8BsS+xAFJtXmyQ
RE97nn8bnRp6ILq4a7t1euUL25HxNMdCGXyRPNNhg/MRcxkijbOYmyooXRgx1lfA
8in+SKF+z0TY7BA9A84MQJ8BDC4Gzth7w4RS+lldq9cyzV6rIBnQZ8C4Aea487Gn
WvBeSfEYu6yEX+vzYV7TaHFvv3V9alxhJXOvtFPMos5LnQR78D5xFzBZXtG5bEGx
4Yqd4t6UUIx/vYUKtJSNr9w5HzKu3Y9+EY0rqRNWQHOQ9wPyC4JW6jSU4fnN6xM2
p+jvoSAPsXZ5FYbdE4Q4Akq+Dp1ZhLc9a6xffpMhT71BCuK8vK+1B///NsPdjsLK
q7KY10uUafuSZdojNMnh3/ufvnJhzYVC8Ad+ysO+itvikRj0odcL2N797EJkLJxH
5vqii/PwJx6OzZLRI9aHDzrxfITGhC81CzC5hA7aAxZkSPJ1HlNDM5HRjkJyExSj
8U0A73KZSBlVaDI82FfpoKw50k+V9Er6an4tbw2l+bJrPQuJHvOQdUdkHlpm28r+
y1Vng2B5oeqPhnLoq9fHFPq8bFv9i1DQOCK5W4Bwl2aX4Nt7QC9EJ4SjEnf1Jk/i
9HDo7/isOpk9ve3GH4sB/WaBMSIZ3hyXvgHh+7ucR7KssgBxtrQMDC/4PXTKhuFQ
sb6W+5PpJcXQdTnKGqZoLay848A4ifBJ8pNfVjMExY/YFq3Gwxr8w/2kmCfA1Wsm
0U/wnIgROf++ScgHKEoikHm6zVXmRh7rSEHfKixPTrIn8zgHZmRuWNaFvlnaZ9n7
VCvhAXEUGEFBClVvTeZCYGYHARP6owtN2PPtzxjrvqd2/bHS0B11O6PYXddA0uxj
h0BBLlL9VI5sAiBiVr8F0h05u2g/DDYxduO16fox4k2KakpZkTKjl7mEr1GxoXCc
aWZmZfIU83G5BCRaeowRX0QGyQZoJhlDjlWM/FkbfpsovYJjcGcylos3vBWhMI/8
ahJosLC6VOwv4Zxwv7oG8HW2hmc6OjLgOeKys2BawrhVfoil2Oqpd1a/rShIsbFB
YXImoM643CG9uHSo1yZGEvp+Vx5odGaYHUDiZMOqxfFQdlRTpFrOz/cOBkUTHahw
Qz2pD2AMeQIWLYHD1+aboJRlAXxGas4yG+C4gI9/jxL4pTefcrd+bpKilOMJM3nE
S04nFohVNrOqIKtUeDLoddUgqLYMJ73sFrRixAhohv3ck89QLJhn2F4tYAd7kHrl
sEBCjfI/SD/EOGwFX5jQnd3nmQl/2CYl6871dmFxkJ6gbppgicMLkcd4AqXBIMVz
niv1RfTGRqZdakd7jU3n4RJU4TDs4HWsjMeSQ6AZyWDuquG7pDTIAgUIxJd2NEf/
NdzSnhk5meZN1HqyzvdQW9bz53Lef5vWZuQXEo24R+QDPYyxPDCF3O/V0S2FYXG4
XGHy9eiR+zFWRosMtRahlEYZo8lrcnQfAVuvWs67e+FkFM+ralZuYEwAQb6+qdRc
r6uwHMgNer9mbOPqfwK4iNZRm+ovrojDE292U6MbLSw2PE+cs0OVuwAN6qsdd1yR
4b5fkEokF3JEdiD97dJBu2+rNBhFzSSAzOsTsHcnPcXEkdHCJ2C3zT+TwvM1yueh
9qznGS8eLNKVbkK6j78EuoiyVhje544CSXLNR9Yl++XYgOFRpyPn0evObxZ2AYy1
rrcuYnpoqTzJKTswtOfwwMgKSlR90xC5jJ2Tztla73Z1esUQWFeNQqwoKNVEjn3z
Gclb4yeDFeWzl377YP9iEBR0fAxX23xC75yfj0EfJOk/VmFzMiTUzGsBqW/gsB31
vQdQjDR+iUMZVs562/GWOJeG2D+SbU5cJ7kE90WGfnZIVFUzFP+W/fJReqgNQ6E8
x3z2ozBoQziFUAjIbSGJ4drNJNYKh58mDsBmqSptRdkZpQ00h1xq0RnzFLE/Ff2+
p+JZYMdWpdexcHDVZ0X3uBVs0z+kat6NDleWS+hvOohBZqgX2S1D3kFilF2nqa2F
5KUUmo9ewBQ6P9UXNbxCIwVtv09aOvUnGJ35/EKdhkni7LswpZoOFmU6fVGJ4ZCa
D34gf1lIYm1IbDRHAxzCdv3YQN1yxT2Sa3y7lOK4+t9v3mPLyRGcGYnnQSl//8Eq
6NbTfHlA32TwuWTK1VP/tGH6T3yOidf1jNAFd74oAwO8LlBUlxTHSO+8Gw2paf/S
L9Ph1m6I9w3olqhxv5nxBkAq1zWbyqDYFjC/bzM4CxvGMBoBo7yaXIr9wG7zMMKZ
7QxdWhHKE1oCCJdvxSjUZbDTGCktk9ruse6i1dZ0u+wMvri/2TX7FpkpprtPVnFN
vZLocqc1uzxjYlIq8yK9xkrLbLbkSZoXCKrQ4t5VrBr35XO2T6iRR3H7H6+kwlrf
uBaEWUpTVBBProkFDV6UoaP0vWNuspuUoi0DYbxaMAWtJiwgD5XaxfUu1cz7uLz+
Fo7MbeweyF+GUs4g3GkndcVPQHVSt/doLyqJU7SmzBRAndLZYiCV7oAh2V8ZANwl
I0Gph6gFvdy1kHCqnAH7ceJr/cw1swIfyEx06HM/eNphAvIFmYZt6ymPQkZweYxB
EeMkbQx5O1XbQr6TIpA2pX8QMkHdEzKTczU92haU3mozPB2+DNENIvnIdxWuRTik
iUBbAlr3Wxzum343qG0w5pYLM+0zF5MAVBGEPbmPavnJ+JnUVF/eE/geUiG5SAUG
3AoZuFVAWQIhiNSD5TF2AVihL3ykUyTrEips8h4FQfGxuCTrFJ3o+f34PuAYPtNp
jShnLYjpQg4u/DPr8B/dZOFH5UQzTuTUHeSh/HRRJRrC9VzsOBCycH1p68c2bw1/
nypXfz7A/FcW6ST9SKpVb3W3D6nfooyND47WWd5PED/MS+GgoZXO0LB9GP0lcXrU
yKy667Hk+ehXJiLjWCKIqkd00DRugNStHTZsiyfdnHUuEOzISzbU1piFqkaGYZEt
muX7GH6puIwdQ8SW/xIjZeCLZG4hCbnSMV1TXLnfq5Zsc2jd3S4cObYFNWatx/we
niEuqyJiW5mOBEbNFSpY1I5yTdLQZhR+Pb2MLKpc+Y6R5gJXM8jrUO/2nDqSgmUn
HEh+4QS7jVo/9ZG9oeJ5XcZbRRvKNzGWgXTFXPUBYQ/Ll7gsOswwajN9yr8lemZE
ctFKSAHAP5RqqZrpKQR3tGPGsxcReJmrux8r5PLQA9QJpniX9gKhMwhcMqnYu9ow
MatFb0OYR4jQMg3t3brD1/QJoNweLvxzhCg2W5vj+bmOCStf5Br4NLPD/jnsKqTj
gXh7LefQfP/rboBvLFFjvbUFXj73oLVJIcXZwshVhTfByTPMcNIdRG9UaEBKJ1sJ
l7kp/tDORJmWHPZs7kTcp9c4eziQ3uQvU8p6VxiRtpgcsYLAjee/TBb9blhK+VdK
UwJTj/ck+jQHlRXy5ZK0RhCWMftnsTN0bHRbKUhJxtV5IA9DtsL8oSABj0IUDsCS
OwzerxoR4NTQA2LPNm06ZP1G4MxrkbsS6/uG0J+9bu77bP/knobjRYxdvBZq1/mb
9Z2GEeR4qtmYlqDGksM1dhMzJOB0WMpSlgmm6La4onn5Ct1Uiu5VCUhQZb3BPyrA
2P7ejh7UhD3cY+ojOmPxbpKATZZkIHO/9j1FLHNb8RyWgkkO15VnhVyQGrTQx8xJ
AQ8T8bMv4mSROCH+ZDerYte3pgF0J9Xg9nFDc+QQyUJV9Kynn8vJ5WYv9bIHs0qP
qUUoHNDll7JbGd0418r4JBF6rhrvw+jAClwXFfu+WSUzIN3XrNfhdeZzzwGeqEDA
OYl8jqSti3JsCs6UjVugK3wGvdn0v/jcYadSZ5zp7ug7wUD71HG2ISbEcB547opJ
LsnV8B9CHvQp6UE0zfiLY5pWlYqx82Mh/m4afFl/Mh+rrRtEba/Xc9aOcQ+MsNWe
R0gcE7BXFi2hynwacxUM5VaClLgIS6gjy6ODYQTEg4CbYmB2QGmoHYhY+/I7aHo5
KLYRGbMIOSAJIjDKa0cfLnBibsSndYXwz1bJpVKqUpQqYVBq3zO5uOKr65MEbcPr
Xokh09kWW4xUu4VE1qOSsbg3/FetSlDFb0fGLC2qZMr3eRcpAKzMZEhAG0DMsn13
0A4zXoJKWH6Sv2gpiYXcV+X34seeutbrXptON3hxqTdd6xT6GINsBRuJdXNf3Z67
Aftx4dIFMQpFXOgOSkjqjLMOFUSt7L9jgs7BtP+z6VHCwTdhAWHV3NWFOUf5s4o+
R9b+5qhjPffWbN9gfXFZ9OMCK6LY7tVGBwBWL3riIMWlGx91JxV7NoEXZJXMB7Od
yVojC7+JVlH1k8282+ABMjyIO2nhqY6uk2gt3IpCqyNA2wKiBYpx1POUToj12bYS
emI3PNyI2pohLeCoODXn4zF8Dpf2RkOJRZ8NijsDdzvJu/EEDCqFcjNUc/KaO/DS
Hmim22HYzN6bMOQ216tLobYwphICigk/yrxGHACnC7i+YUZ8fXAFhclJfwJV48Gc
iddyJR9x/wfxF4hDzusmLf9wowTrZLGPG1EkE8WLpd+OBReCa3aWEULedMKsOaRX
byNMZQqT17dP5aOtug+HW2qLXY/kdVuHYAUvdNf1c3SrUY91cctLOul4USke3BAV
jH5spvyvvdjxBpJhvSwY0MdkMWh4ioAhGxdUN8Sr6gPO9+F5kZeLf76X2KOHkGNS
O4bG5CPzucsTm5+4QrhrPa3GoJsOVivuU8Ws7F1FbgdPL1+ewFVYORm/9VmYUwVI
eIL94TSq3A023iJ2Prn/5vNWLz3M1TlTBvTODS7Yt4uZ+tc4b0GQgFPQpYL7lsWL
30B5LqkPZn17JJrbK9SaI4+1FWY/JpeHbTuoD/YBX1DasBOp+d51CfUMAdlaghME
u29rvoVxFtErYbVHciJyeqiEvtofA6WK7T7H3bcOeBkPp8GmuwipEFXRQWrRUBjL
pUXBIqQFQepIAs1Bvx3LEgu+3LZKN0PFncZorA5CMN07QTTIKtLeMLksiEdEMLND
Qa0rVkTMWE2GZ1Hmu8sPzqFGIVjPRx4OI+GkT+EJR8292uF8hvdfdpVUJm+8I/jp
aGi4zsp0lAzf8oD/sa1TvafUqSdTYgTWH//o+qT4JEPSlG7wCneGQD2ak4BUuXE9
XUJ9zBDpUNq6isew2DpkliK6O3eZOxA1Fwm9P3sNimQXZn4TrHLtbXrKyZUosafW
5sD7qvSk+zVs1jApghQZuPocfZkjg08Kb1kE0AqaGR+64R7AnzmhKq7pkQzkyLLr
RsBDZvo88pXHSYrcjdSaum0Ncp8r0Ewohoh+Lvg245RCxPdybVR6Lo/1aP5alImX
+ndlIcuEo6uhd0QiKxMn2ZIjK8TBFcMl3hZNZ/B6dDPsQhsDiw3p/4LIUTdVVBK/
3l89BlUIYhQaxIhCd3dgItLlGUg5cSS93bT8xjGCsT0IUOUhq78Ce0YMNMWKmvoy
02KvLE+K4JcYQUDQYF1k+pfHVUaPBbscyFb2rzbYiKjPI98OdaULUf8zf29omLuU
dZyflXTRjwQce1z4y7PjQ2wk0EacYyEDxZ00fXU90M6BAWxStgMWZAJaqG3r0Ler
x3MLjxELE9ousBNiCfBSnsu8qiIEN4mW8J1I9XfK6OLzWZ/5bn/oR3YT8wleHgxQ
8bPg54uaWuyOJxHH8/kTSKDKGGuSbQy6Id5c0Y04oFuwPnqXcwWe5o+0NNbM+YmK
ePyiX8vTEOY0eA5DM5oKnZ8E5fgoHAnHMa1R2OF+ai39B3nawoIDFipyfgoR0USp
2ENp3pIYX6kd7CY7oMxia67QdwfaOhByrikiraEfFqAKpNFRkjTEHkU21qwPCFfY
8LyOYOLw6WExRbx7YeyKmOgaAoma+Urf1RZX+GxgPZVjpoWwZ7yhlSQFbR6KqCcP
uIqJsnxF3SR05wq8LOBDYY1QOpRyJeoE8Ei/WsqvLvk7YKoL6MfnPbXM34LSBK6Z
isLwJdEVOBVEj5r+LuArwXUVWtVGN85O6BMyFvbPuP2YqUnRFyg3g9ZnrrELqaN/
lZ2PK3h7EQYybEhMfk9qDsm4UsoXiFjVstO8R2JkscpsKx4kRk5EFqzSNv1m5xgA
IvgMEgo6ty8caMSv2KbB4n1LJVu55VF5QoW/Os1w6Ft58IRutzv9LtInvvs3NbFU
AHPN0LYn5y8L7IFF0sN95CgCHY2V1uE+OlXZCUaY/NJiytTug4VY7bmWjBHYgCPt
eqUd2W8NsKMcU8ZmV+hS38yH1TrNUD1s0VrQFsSUmI+ca+YIuOAkLnJ4tyd+pXJI
ruyDguSLfs9xKHQtV2HHd/xqEjpkCAzzQ1xsFDJS9OV2lb3SaOHFUIreTtbZ/swy
J9M154ZH/MF+P7eUIF4ppXg0UvtQz3h3sxIk+sfd97QQ6xvxd0zEUIC8odmvCCZu
b/MbzWTjbQoUnVkqtJaop8mo2Mv/AzTFuWzYzj/YCKly64z5YkzUVq4qJ6vLYpGZ
q0MGw/Yf8vk4hZ0RcXdqtdS/wjYecHOIAKJYkqOFy2umSWJUUYmYiGlRBgvJQszs
9T2G0CRD8UBLSP0hPMXsKpjB9W13SgLQfn39JMnVZqayXsKfoEWkTKQdyACPj7wC
foTCvrk7TUCGauX57DtBUTfGFxdIchzghNobeMHZMUsjTqTl04AAWLyzBI/PJkgw
K/kw1tYnSgj2fqR12BlFoWCP/B2OrFGJNeMxxwTCiMJPjjQnesG0DcTVMoem51Vm
SsOgI2x0/29wQA2QUru0a+/JkKjoNW1FtFT6JGpGVeFIUlYSO3UfS1cbhhiftB5t
4KCSgFtHMi7U0eEzgUwqC56xf7KHaIGM8qXUYlTfHdCkapOxVH/nMnApNxp3wB1l
+0p8F5k/b+oms32FmWVIuqM6E3PGek3jBQoKkbODr0bOqq627Xkkwz2fFZajFffT
6q6rGVy6i+AP3OZiJ6P5nikMzxw9Beq+8+SFpGj5golLdeKhuO/RPe6615/T0zlN
iYvskIu1e28g+/Uou0oAbR3IWvFBMhYS3RB2FCy2PTxmNaLt8AacIlCwte5e/PVk
vvjnazr16WQMzZVUTjFtUh6J3EVBUohot4FM5TpdVMVvN3T7nkh8QUJh8VkLmCHV
YCQn9cq8rjtzJnZN5ACX2OpKr9Vh6bf5bQsekDlG27+nPx2XcIK93g0DhKaV89LP
MeN3WfANyyL/rLvd9jp5efpkf1nNXD7Nchwie4hhvDuIJ3hQX9PGinH+Ll30M+6W
R7e7ZbECYG99WkSN9q2XmVBYgdk/YH+ZVKJem1b0oE3NkTQY/PGnmtzaMO1IoZkv
M1PKbOqRBdsrfvhXJYCCRAta0Z2D06wJO2YJlkzSrLI2tRiXAOymnSBUIoyx+x8c
SddC5XT3YbiWeX0X6uENmwOV8exU9xsm2c7tUN5/8UbOO6PngOuASncPcrMYSFO1
pZ6dVS+MGTG9yphgdZwwCp1MdsKVALf+d3Z+YqNqP6oYXv5rrACwF5GLxw2Z/05M
QvWpcQ4+nbVyMRhbFexO7GIC1Ac60+d2MTv15S7JBMnhJw/Fd5DMKSFI+1bW/QT7
osA9tnX5ZN6AH9IUIhxamQIjmAvuxEDn9p8h7QtsBy++fwpAOzecpWPRWCDwiRr8
ihFC4a8neR5QK0dugmXXJDAqTdoAJZZLFHNb85yX2n/4S5ZALndMmVPGIu/j/prb
/mH/9FLYU9fMbJzk/PKy+nHqblG7G2w48QGNRaKO5pdHx+6yHpot43OPmJdnUOh8
xPnoB8CiqdNaPRqDsIXXeXPxb37qM/zhv4JaQrGteMbivQRSYapRDTn8lnQe/pJ/
dhuU4wwh9EdmdDGxNAEk0fnYrLMATUXDt+h1YibX54/1L1bI0FI49QMT++TunKNw
KL57jgM4DD7lo2oRgicAxiffvEYYJNUcezgOXqQl3kptFZ3ShPjh6W7o1wNawRvX
9CuSFgozSLd7Z07x4EIH2dSj5nuvL0J2keIklMJ+YmM6oHRm5sNfaYVi9ta5tiqS
1C4J6/+35bIP6meSiw3Rg/2NuQAZY7ITD0kwbtV5o8fZ2e+XrNQ1z9cWkjrBMTsA
c3cXdBi0O5QDnxuvDNpKWEUAtynVj66Fgo5Gih7p/CEPopiWamNf+EiDD9y7hcfh
3pZa0Aaxm/xpyGAg1tZWdJOOH4MZtAFT2FzCOeuNpUJeZwVQyKTbLHkaU1/IT1di
i6a8wmmhTYhj4OP1sQihr36bpXFb+MKyHT42g6CZZQXpkaVERSxwTNX0l0BCxnrB
Uk5El4Gs33SxyUlMpKHSGW61gj25WUrLqAtWLWR+U+9ndEUx0kpkusLo8JkE9POq
KTS4SR/KrP7iqoo3rEszRZ72AgHuTV/N6n1fGIs73cMWI/GDG9eRuiVjBzMxkGfc
8AKwYUApkEJwmPIhOf8d8JV+QYszTMUalmXO+B0AbIpj8tRXGF77qG6ooCQAo6DW
WBsMA6p+fpYL+48p7CJ4l/idpFb9VBnf0Foe6dcD6Cv45weNcRAWM9Mb0XsaiaAA
fn7b6WvDA2NkZp7jDxTuDEhfjnT885y1KmBLQKzo+D88UIV8hKbL4mPHFv/w8vOe
fj/rUbqWnGR/H/AbKrB0oTXfyiwEkxZZaXzHMIrYST7Fdf9L3rHxS8O4hCOJ+4LM
kyQkrYNkvRHN31LvTbb6LSZXwvRTuwH/pQjiKZT0/4N0y4+kEydV/9MSRwqMPLjB
+PM5qK8HFCo2CRVf/3v2uRcbUYg475WrxmobV6jmDDkN+wpKeBSPzwkJOD5ow9ZD
ZJ33CttKMZkE+tE8exwNbiDgsO3oieX+Up3QU6A81a00jHqzTGNmttg2gCsCM/DZ
LxOF9kYS8NJCT/Vr0j4k+MDjV2+M/p6let30FURtZcigJnyT5LoJvOUai7/ZFCRl
jyUGOh8LD2zCPn8fYOKAAYlAuNb9r1hcC5VL5vac+M/2zKRYYGnJ48G4S20kS7Cy
STz2ehZdWjuOywSWF3GEdFmZCvR04kSOSpz6uT0l/h6BcvWvXAfYP0Xy4sUwqQhp
mSgrVPA6tv0ASNZmSfXQ8XC8nDOrXrPldYilyfeehOuP6hN0AAXkUDOKy3o28zCl
sHey730wbuQ1ZauKFY0z6vIms3EjSN8o0c103U3zvAH0vfCNfjV7MRjM5brFLuyi
Sxi8hacBykC34TwtuX0EAOvzMG1O+hlLMxQIFDkL+V13iJdl76+kCyJuEPqD/sH+
0euD4+HrEdW7SRF34eW/0Y3VLZNiMx7zS5DGt2kyH7gII6k98/CoGSFE2GAIsAdd
ekklwytpVrkO02EnLsZOr6iEAJ5LQLC94ogOuCGZu8RVfvag0MHm48MUqY0iTkZG
0+EOJl7Ynwfj2n4OFWnaOd3+OCD8KbpE3aTLOMPDk/GerKCcYl0yJ7U84PjAGFNJ
RJQjFExzdC6yRYpkP7t5quA+KnBZoyLpGSCexmMpcZ3Ne0VJq9SKS5ff7sETF6Q0
tb/aLjwZhS3KjNUk3MVIU96ESKsyLTJrDsEU7k+Hhd7mdgFQIfozUkL1ZQ71Atpd
wIJ23dNw7TMZpw4iBjLv6ZtGl/NHezF3xsQOdHQYkur5GiHXDmzwpc+q+mt1KA4o
geZ2UuxqfuU51BAqI5P2J2AJvNFs/UxdKXmZlevRnFBgBcf5U5STSLi0ep0L+1fv
NLP0Q2fb9nC+70cHQviqUifMpa/tUq/cXCa2d7iG2bjvSykLRq2p8ofuofSf8IA6
WuZ0jVQcOY5TjeEzM7gLxeXLsbFAPkTSnarp+g7Go+royF3wd/igleB+qkEtPFE5
x5S1ksiHKpOSzpEDVyjRzzjWBNWFMBFCR29vY3QujeCRtyRQEpA7r9WB26olNn3g
1zaxZ7kueOIV0sHTg8D28Y0TWGE7/SOjnqaQPQzViXnXvWBhrhZPt6ExGrHbjsgu
gRGzgL12toO/4NbDMK+CpsuAcKnNJEGJJHliwe8ishIG+DAucwQaj6QmInS9i8uv
TadhnCKn2OkVyNrf0DB4h8JJIDbBV2dLcameRGSa0rPuk4Nd4qOGZi0njkqfZndf
1Hx9fObdcW3qymLuv2wYLNyIkuHHGVnro1pk/M8CBpCT8uKhexM6AqDSWVSsbEHt
CRBvuFDoeiqXSB6ax/iyxHfRoiVgJMrpLiBXF5CtXUzGmSti6FoSNL5fSD5jB786
UkQnJ8RXckbYqDktmdha3rpJvcnDoQmNDadTth+V2IkJGfgiVDtvU/OqbPkb7Kb/
rNtTIZe8Mj8wC1/t0HqBaa8mxzjwUMCNxANNE+Sek2BdjCc4U4AAq+JD/lnwMfaS
Mczeu2k8fAXQ2odhnYH/FOFy0cCrSlnMEiMhR+8CfRK7KWbEDy7xElryGxVvw5JA
vwumZ3qHGVd0VR0omWQz5H/FcNmdYGIhnDrNfoblNgUNfA5g2ohTaL6LmRW3EurF
9YfTk2ohTKN8ac75FQ1/sDHcR7kneg/InqDN/1sbOCSi7oYtDaUOGRf4T2emjft6
kGyEfPe/H3IqqhR8Z8WV2vaALVBM60RZSK/0ndoAktmk6pc2RiTPIA+s7mXMG1B0
mLL8DUF0yLnGWhHh9JmbxJEWU0cquFeXUNxbJeYWaWowjko/tk8kHKWFhY4DqH3D
rDQLYbPru0xae3o01wKN251KO5ddgYE7awiyirBkmB06aoHE/BOwdBC5SU4MXiA8
XTTbpYpGF82Zgy9Wq7xC9W/yesL8yE83MmJQxifPCDYnZnHFpzwBcmDNovi4OKTT
6dD2nt6Gm6dZ+WoLdNuvoMWrEh3yuAztn+EYew3NlpEHG8EZS2/tYK/JsYlEmOhq
D0P7ZQwmnWU8oHvPb3DRrrFTaCqfB4EJy5TFvrs4X82iPMNydp2st9jo3C+QJe05
bvnVWNyv1zmMzqj/QidYaOeQfyf6kOOP7go8l6kgTdtc75jPwkTIKdLyC4+sQEgg
6tb5ab9C0GaWklRRqNW6Be5zxljpubcje2+IEr7YBkhICR8YVQx2k4zytDhxx1rf
b+1F5TQP5u9Q6JD8UJvMM9WETb4BlryUNSDMals5TpJNYtPZofvPBqso8YHQF6rG
2cacqR35p0zTCj9rsZjMOFjP7/7TSVIOZu6/zW7R2qjJsCrKcDfsJBJJYB5iiJ0e
/HrHt+4eJ0xPJysCV1tcxtnQwiEWebnbpoz+kt97yumgnqMcfPS/Gji2wAMRO25G
HCX2DQFUBv0uAsNfyTFC62uPb5hLTRWo4XGJ/5q09U+nseeglpA7/uYKg3IwSrqT
pN7zmgJVh6F+rVMMROIqzBAEdj1DZDmr5tse5DZEk9YOlO/xknW9ivbd8BfwaQbS
cB739VEV+Ch/JW253Oizq1p21TP0ZmY+iQDAi8ZCY0s+phyKGV/fYLQTdJR50UDZ
vM0B3jyc6N78shAT+gFDOgxhd3q2FvEJY95uhPNeKIApsruk2aHzHwhwJwumxDip
eBjsNsdDniYA7jyWkpweQvuJRzevO4Bw6wutBG42Y5XtbjMTKtOV0ZMvf4EYn4vs
hKTDkZHlJTO7B0Dh070BOPAZuI1XJnobCOnmagm4fVdnGHXJAdmPnwe0mV8AMXJn
+oiRRtBBBreq5MQdqvBEUEpxJxZJd8Rbmz2HMYDXhMpmvKeKfEBl04N6JDZlwTAO
vbROdtYxfX58wJGOLmNqLDJDgmV7OtuiwgYmIFORMklwQuIie/rwTV9Pkqrn4ZlU
cDtndGY7I6uQD8MYqPN5riRKwZcDbPEfd3ZVxsdQ2B/fUmP+24WQu6UiRVdpxmVb
IDsNpqeHhE5WAs8MAOoO2jSeBp+BPYYZN+YqKW0PtAbn1xqLT9vlPsEUlLdj4bru
OcM1JbHRs6DhkxcChK7CSrBwXyfqup5lTG4//bK/kDi+Sb8OfLhLExMa3/CqZE77
lCqsgiMR89qjc0sProw7ToFbsSTiMahuhjxMscwEgiq9nZugahnmpd3UHG1Hx4Iy
CpgOKfNSnLImw2fSoZ6EXL/DSycpqhhTEoUKdY3ASmLUiXV0bH+m8P+LoKZ2ng/b
aPpCI31mfdrHkk6g2o/L9TBwNLJZGU/M2lJTMAxJhf0eNX/oN3AT3l7NBg7DKXEz
BSjj5vqm2qJw+exqyxyo7wTbqDvHtFhJYYueHPzNtpk+7/7TzI2GZHAn/nvRUdB6
2Omd6aj+SzpV00+AwtiC7KD1TH+yCxoEGu6utPxv9ybM0uE3VUI4vJ02VVsPG3o1
sSrvtiQKDkICdtyfpSW4KVrjkprCeSiqtSw4pfM2vXkfJJFo1t6XXwRJMuEdK1OH
n+E+F5sGdCIrGHsA0AkFt2YytbnOxpJJD7aT4/bgHb00AdieCvLzhR/h01LjP6vt
LEot3UmV2b8zMoE6FEyruqvBZc2ylg1gW8iQOiIAQ4yf+ev+P0E1/xlj7bliIQmo
YEaS3fSoVMogj7IVtoMp+D5KGiUmvhajpfWBVJEevrj3sso+1aI0iRf+PJMnD2rM
17eCbO5jqvSxeA3zi9a/zQSo/xAxEVfNu742rH0tNtrPyjlX8YOBn62+VHfR6Qdp
XrgnsEkh8T3v+aLbvoPLzGTHvqMN1rPEZZA9/arbktrezJYC5NxlVrCWh2m9ANZ+
CB7Fu4gNAqbiaXWPx2TDob1S15Gbg/iEBRMHKjPDFfyPy6sFG4w7wGCwYDroy59Y
6XWsMnZ7OtU0xMIOM7bFbJISzZzGZ5bkXn1mlJ66YX1in7Q3VPMK5W7Q9Ew4w5/y
d2GTOoFVJRrGDaWAuKtVECLX53YrqcKx1jFoWc18cNPikUF2gngUpNUNuaRt772Q
3/M7q2sDaiq5NMXcurlQ+Amwek/e5p4tJ9RY4kKKx5a+5BfpWOsscWz++xgRCru7
gBSkTl/XCrNK8xKjD7lAhVDS0TD8p/zBqhEgsi3WUuE/kMAlfcawG6jjBDh2lIXt
GHz/rkKdo5XDDA1vsBYZXysKO2Fp9P7tOFK1du716r/X3xvNdoSdypAZQ8CnW5p9
GdV75fgL1wyixcWYivIwpx1ruEz1Gnv39dgM3qddqndaD0uvIZ8geKjypZCo+cy7
gyv2VXw9X8NNwjlmHKJ7Iw2HsJcCcGY1GBSMEZCxiU6LZYYHcqqKPMQwWYLNt0Bp
uwcQahlQOgxpNbn+Csk8yLu1JF3XKeo0q4JA2rxQjUQN0/dQynantLbLww6l6cgX
yz1zwyX7qj27HTlB+BSf30JfvGzRBqj8LwUEFSOCDle2L4w+xsu8blvUJSaZx/Gr
puFdsY2Qbq2CVPxX4dPvk4bREj3A6WcS4lliN0tJvLUxWb6vRIXKzbh+i5//eg0T
0P5RoniWjjX3h69QbZ6csLf2Z6jfk6RPlmt+cQWhV0H1gWLNl4tZIpwxzENfcxtH
g7bGLJLagVwqJkC/27YPeBQ0H22ANDrc+FPuB1YFUSo+7eEl9KOJ8sJhYyaSCcqF
yW6SAPFfXyCPzUA9jPnZMXzjwPbIUN0JwQMj6/3lZT2XkNiMEqwn00zOZ12sDMhn
NyOL40sh5G6TQM1eSGhTIjjPt24Mr/lK+miWF6KVUD3BMf6LU47uYm1sCTATEIBf
BvlBRbLJWXAoptKNvWRo5QcNKzn0UKZm9w0tkiVUq1UOIcKMfciaNbBbgKoOUKMc
hsuNvMRreVqtcayaIBTZ1T6UggpqJpInVW9qdow4zcjhnuzvoB+0zIUxaaCapTPf
wjydYigrqQlFkiHLsFGBxYB1mNGE2KShrYUGJ2VSMpmWcSv8Sntq5ozrCBk8kIhl
LkttRYZORHGHtTa7fTGgM7ezlX8EDDxM/aJoZ3pTObvC3Yy+gFgcK2291S1I+OXX
pWoAbXXl0Neb4xVESdOyklMY0wGFibSW6RuLmPDXPRSrx6taHtNnZBHse257zVdZ
7ShXnF3o5UhbCZSom++yZE1zDM1pPAA+OrY9LHpxsLjqjhgeUhwwB+3BSJgbnSVw
aGx+1uXgr62K5l1LUEO/3tagBT3RWL4AxxGVikPEnxCYCYDuhZfRJhIFo02byssH
r5kRtRmakjF2atEM8aGVxWjH2sO9/f51fRK2kvl/KJON2bpRMzqDiyvqGbVUD111
0M9EtuP1mjwe9jG5G8GY/PnJFl4tS921y5zoR7FdOfAvrQSQ7QlQY+6Vn5wula77
WIfLdsJlxhyep4q6PEM12/g7YcZBRgH4YnRca8CdhC7ddzbGyapy4fgDCuWF50qq
AUotMWA6sReCS4FIyaw2dCDuTka3qzbkwsb4VBbxMS6OeqjEiaLq+Nhk1Irgf6x1
OhPTo443OK7BLxxOJSrZKl0RufnJ5q0IPVpV6gzsH1A61c+MMZXMDc+AP2c2O1eS
tzMSnu4bexebsJNYuyWHd2Xop75P/s7ir+RGS68N3VrtxcLmg6Ff9YfQH1RhvvSt
YaR6D6G0q+kTs2/beJgFhIRDwwYKeUJ+UmyPePA0m9zrO6vCiCYQ/7Lpm4JHrOoB
wjFVv+dU5EwnkkKSIKreWU5KfpTMlgXh+G6qVdJ39Pa9ALhqb1/DhswCePVL/t9x
R3+KgJkuaAQVOvY/qutg5lKQk9tdJO+3/6AAVHDlWrUgfM1vWBw2yBmfBfvs6xhn
pKQxUza/pFTSk3mBKLCsqyG+UBc82lTh/ygSejoDh1yaI+fggol758uemtBkrXTC
054/WvOAPiAYEvSH9gyP0dsbCvAGvcgkeTwxthS/foN849xBvEdG1uCbfNR2oDmI
nU/je5+pdzGOJeskk2UsT0cTn1KAvpeSdmxsscd5xkdfrTzh+rClphW12N15BE7W
zXOnAEoyQD8rCoFPkrrBR9Ed99IIJStcwydLO2QpbPdfk5UetlhCaDEkh0+TedUR
4+i+I7E7ZrDFIQMU8h0kQHk//ghCDtUYHyRN6uANXUHlOQ4rb8ao7aAwfOCOY5xO
fzNmUZR2gGHaTmQzjS4ergX9Sw/rQX1wgrteB8DivA5UMBe2oqdk2bGgSxl1U60x
hJdgeyzx3m17hiAxqcm4147W+VkAnavdK8KRrJPtC1u3TwY1HIomes0jRXdaLRlW
g+doL5Q9b57QeDAzfTZlDGgvruU6TP8NoTBM4PqG5zgyNx938ER7KxiFMzFxxF05
wtfZqlywcus2fYswl3i5pp5IiXkO/vdIwlE8RCW17z02QwDLOTdyfqp2+3Iemrky
MXiaU/xURC2mHW3u3cAi9klEQIxzVbPeChgGNsfjFmwt3CBK2CglVD1vx6Wgyj3H
wcWV+yehcwCC6YJBe9TWHIlCcbsfXvq4elX2gD0Jo+0IquLWNR6f+fYfEm5pqeIS
Ryl70/5UJNzn58AW6vsw3bwPjraEYwxsdIuBrnn2+0w3f5+h7EIcLyugYZPL51DG
m0z8JJCITT4/vqvdwLMxPrfVn1RRQ3C7rUMDAj/AwuDw0kcdr2V+4C1W7tpMkxuR
mjDfNnnHpDY3wpCFud3sQ3SgUu6Q64V1ZqPvy0NPH/30fKYRAXpQxmW7ImcVvzFS
uoPKJRdsbjmMsNFTweSw8eeWhTCVaZA0LKCPYOhVaTF0nG75LWYDHUaVjPriJK+J
st8RReB+wFX75fpd+G3iGD9MqAfUhl1+rZx0k0o/96Po6Efk1PHrZeBjyn7OUOI7
1DeCBXuHXnDUmoiLo8h193U3bf+HyaEV5jyUZ5saFmAMvpSljqhjaqdtDMlBMn+5
GjiLkMwFyzYHbtk7+oUNXsOg/DsRq/86GWZS9m+FBaxO0H12xlER5ksxfs7/aXoU
HolRGeiQEZkc4nvmI8yE/vCbCU/OLs9Bh8yqklYEaMihbjbfwLZzKiGZj6w8oXYl
pu7KGHyAixVg/+PAW9qiNfKNlGPpU4a8CWgdJNJixS2+DCF7ZnH/9cseVI+Pvfgi
0i56Z6Ys3ZU2YE52S/fBR0YCsEaeU0DVuBoHu2KqshrIRGzkHXlUf9FWnIXrKOFb
HDnJsn5lrX+JyZyp/7Pq3q2EAQBT+zTrIL9c+9FSe+JVruW5lp3FTqRSM7cXe/8C
J8ORZf9nq6cQMek0tH19s8tGZAPxaMzLqpmD8ji1bBJOHqFQTkfT0EMmV6btEsol
JvbEdLc9EX6/MOQuxyG2rHIVMAntJMbLjnbbyAgJb3Q4r2FloI7UHIOauz7gJi8r
BFzMnXTVuiCvFlOWPTOnJjsPBzvpGTbc9zzE7ylunhA7tjXngbZfuZ/bKbl5Tn/l
ZBOH3tiAzUn9y4MZ+IfCMjrZsW6yDhyS0n1UP2N837kOc4iCJSJSGPHkbP+OEw/v
dqRA8goVnaWfNwsEWl/OnWM6DoKPV3L9uLIV4LujExlpowos09Dt0dv5phwLkV2I
B+AA1G3b7J7wgCCysE+GX8TLjF8jssZeTCql3VmC1x5jwCqX8No9CAyFoX2HEXgw
qfHty6hrd6klEfHtNYL44Y0QiS/M75GbAWTQjdgQTdgoUBaRbebkxUVYirsJGwXz
9uLpVa0zWPn9xRKpXzfhMXspXy4Mbb77zuWpCC4wEaD+//aA6pf91QX/1avQBiwJ
LVG7fc1XEdu3QjHFAa+tpC5UrQmUVrDKuHgJVWYWMryV7bC5k9R+H9wp+eieAAYJ
kND7GCjK3ut3nJzhSR1DEbd4rQOHHAnDuS/p06JqVpAhVs7UIH2MTtWIIxiB0QaW
VbmGE3fssbUwNIuxhmH1Xixi5SxC0lkKTZapQ1ZqAoAv+j+NAs5Iy/4SW6ZkryIU
Z8ZaLKCT0Ce721hOgIjvcRCSmgMDRNaO6Jws21le7AZSuI3UHgGyprfvER1v8nHn
7bNWxBhETe5eAWCRJ5RVgDBeUN2NLyP4JZM0XKSawxRT8cUzYULasQ+YXR6ZQFhc
e/L55iUM7mwIPQ5xJACq/Gw6jLUvC1Aez+aKMiz4y+5qZJ98L6FRwm1p/Aw+spVE
YPqfzWiybJIFC3mm1bZszbQ48MTpVdDdLUImTePYoxPaP61E2KV3wcsEomXVOtEm
aezPrUKQG6AvZfDpw5Ot30M7lA8KlQaMdrhRLLVRj7Lv+36mnoWHJ+CbHVBTaSxP
rTNZpIAGiM8vjReapnPAwdPqZFx5/uXWGzoM82kFhRBldx29l9RJie1TYR1XxU1x
cashKreL3n2rC/q9ej2maUPkYXsm1sFNL68KHT9lfKrTrHPZa+yYMUe945Dam5bi
H7OY5IhYlYO4N5Bmha6N0VjNflTN3KjVEV5+oO4teBLqSAgSOgsQDsvIsWlH0QgG
JGYsE1DTIexjrTfcVQ67xxgrf0DwZK9+gbjUHE3Td6cNDE0UxH8k3hbm8FNTxOzM
KXaL74Sd3GekKDFy79GtBglG0whMw6B7UvvbLgAvzazaaZIeYupWHIHqv5NRZM4o
03rUxNASe74+KfGRHXafCj1sl+xUNDiyfprxfSCv2eUZtj6MPAOXX72D7t3o57TW
M5Zc7j0KPh/VdrxhGvDW1r1MJwO8SVVLseKhorgR1KAjNlT6ULZpsp/a28QR0Xo+
EVYG2R292Oull64h37SIwhe0AziL7HIjjHN8KqvDZOkq48xelV9tXte5ilMY6x4a
6jw3ejGxpjx7EdFAEPRDnl9xo5TPsFIwiI46KNFwOFAWiGVA4MsLHfLsu3BVixP3
LuZGog6oQY/FpphhueRuoQV+neVRsf7l0kyVCp2ejZMecM40WMA9xEmYfPn6sybW
ewXfaBWXg2x6/u9pSkzmQrtYfwrmkOOS18VoCB6SyWtHTiJ6AOe2U+2pBijMDXZt
4UnXoYD6lgVPbdNkInL7xIX9oDGTrV3G9jf2wJguQY3IFzspFmbMU0AjV6ry49h8
p7Fk2OZ9MgzR6MdnENLRukpto/orcQceirK2rM7lxoREGFqEWGh9iND6TM4Ne8bW
s+p58b3zj01w0yqLPTOOlRYQSDfFKnDWXX7Tzr1LAkyp4pWkUShA7m9fYrUXW+5q
mr6MbfQyUXJAJAJ4KyG4YagI7tgdG/uGr3tl0ShBr0kZ93mcfATEpLocEPMke47l
eNSC9MMq8HKOiuhO3ailmwpO5kCS2eD84seFKTplYuI9/aSuGIksFUlRwOhazHRm
IRROtOBM4ldtpoOmzp48zHTaVxeACZOcnzP96vl+198dNMo/E6+OpNWZbloT8tno
s/VtYh5+cGIYXE5IQ0jicFqoij140J5KK5CKCawVGZ5JQYQbuyza5ZgO64aDP42u
G18tOxATADZgU/Eif5CSIFHWrjQ6nhr7s+AHlltL/MYlln5aN8BEEv/t4xrEeNQu
jl/tcU6OmxC9/6vexcU2yBY7d19y183GCVUL3WCD4UpbpPPcv5WsjmdA7GAa/wLa
BhOy3PhLt3Mki9TfT9KbhoI6A6YfDWDReY8NiNLYlkYAjSDtTdF5JAeGgB2ox5J6
OOBuYAm3Yyejb5XD44X2//nIuTfebWTuOv6cHi9VSU9aeiLRa+AwifiJxhdF4UmZ
+viUN0a8hh/lPhsPGmFpJrl1/1zrfzFJz7oaczG1AVuwW5uDPuS9jg2s2YS67VOB
8hRbctD05u8r4J/ERA6HRvQoYICljtPkIIKbYw3/V+7w0IDbKFNoZ7Jkb9GhlZnk
QgRnAKiT/s1Xe1zQHil99TKrggQ+l/RJfxdF6tSa+5aQ4ir4thFA/WGAnnalMOAO
cMN1n1bZ5PYdm2oA5BWmJttCFO5SYN8KZRsu3eC2rNVnEKJC6fO5Ha7G1mTkM24t
LI+ljznPZKwU9Bdgih7fnd//VQsNRBFVDlnm1yYNdHl9cCRCpI0omIemL0pBCkV5
+S5LMaKbS+U+K67VNT75fDHMMvDUujH1hoTwSAPCpyz98BdP/dSncCCZZ91q8niV
6epKWdHKoXfddj8nV8REtHHyxTP6U/8B5cr+gjNRdzVCaP5oqrPh2GeU5aNTCS4h
R83DMYIpGOv0pAnto6PkdsCYF/672hJyPjzqA3yVXBUssSs3a0qrWN+bIsV5Pmom
t8SqoOPRux0fYKDzT//ReeXHcNafQm0zT41PJ0A69UHB70T07a8ChFD0dDWhMh5R
5XDP3dYK+Bprgkke+GPE7PNEjtxmM/vk+LTEAvLV709+XtFiNhAcullqC5BCMsdV
IFpQ4pipakUdzXMU9q0Q6ooWO9jGZQ7qUdjXe+h91CAMzsp1McWHpaoVleD4xCb0
5zE4aH2dQTZ6qWo/ZiC1PrEeWbM98QrhwxjvNJqG2Gge48iGS5U+vbkStYULywc0
o9V0pQCo+xHyZH2xKixosoaZjK5Y6Mng0JHWi3SYgvhBe4JhtP8NHQmVMdzOI8Xv
vk4aPz/+zFwXR+98dYeOi0B4EiFxlhDw3QvAQ6PNgfFB7OVlP6IEKxB45WBynCSA
TzxP7RVGaB3GARPKxSQb+qTlrNCaNC/nnXLnK1PP9WDGHtH4a8TOKm6BHpRyIKos
r5ZBVOjs1AFs0+ORm9oUNH+RvEMeMFxrgw6ZrnpG8uYfhtBHzR1nVTe9rHAFjmS1
IYbqul98r18RVoxMVT8ft50H+QWJsTsFOzA67QgUpg2aIilf+hXTWi3xB2DADAdc
I8R5fB1DX9c5L/K0Aj86yW20mP0Gm5fAm5si3Adz9DGMRoRgShG1mAX7kTGEnFPj
GkbLDfW0fj/o3MyikP990+Jxpd3hQ0RtN9qcoMXRxcjdi4R03qqkCSB6/ERe7kD3
g8ugJFEJoo4F7HCs+liRFHCjMj7vUMhf/O8ZCyAZJz7QHfnCxOlXmxn/I8ptbnRT
63NfhDtcVVij7cfazXfy7t6vcU6FzEjK1bd107ygrfGE4CXezbNVlmMaltZavYvL
KiojYxPPnC26UgbDr134ChNhECyCWwX6gNtCumMRmy65FLLDZlTuJrRzdYzgSiCg
QkfZCbeo1nawLjdyi9/dbaJQfRj9l7PkVT45seCmR/utIdebJZ1/UV4aVU2WayLi
nkS2ZZfGXeHOyHCBiwSInVtOeQ4eXxM1AgQFT1ZNv1VJ4gqfhobMTpURTV4vO84I
H8JGuWKHpkTnR+mSweOaoeMk4gM5jlPgKWLiqxOMNOJDjhL2dRV4pJ+Tep6ZcVOs
b9PSz187SDzZjPGZPyNNS2fmhaymRkQ8TkOQDaJkUDSJqrwws76C0BpeW0YgA4S/
Pn9KGu+JdK6GQ+qf8X64Gm+irJpk1Iz4jr3FOP0mFKu6JsrZ7N+wk4mz5ns2WRIJ
1QRoIzVAIheSImlRGmK10Qw8odWM9o4dUanSJfPcu84Bqkiz3X6vESfKuRDFZAgU
JGH8X6hzpnzLJVlTLfQ3WHFlwCwZ7/+EJPqyMASxjMSyv6xuedDPsq+qWzsYiHPO
3WH6tX5VVEIDyVSt5gxUsckVy69Qega3FA36fDGKfhC/RqjxjbjvUS56E9/yizZP
z1jQODyigm06bDxQenHoOUO/MVBhWZTd8n6SUw8S1thCuUGxxLHyVg4E0G7JnoaA
Ew2XxYeZH26sj9ctq2tGuBr6dNStOBj2IWxph7sYYXW0D+QjTbfe8DMFWXDRGRa8
EqxBvADnniFDuH98uF0A67m3A1jucrVn6ygXIcGoJRhrJcsdEgLpxi5CUb1Vt3Ng
scuqDVYeh3IV6rUIGm3k8kBXYLaeMUaDXbrQhOmp2YJ5jpJoHXVGOvQtUxtCSydX
ZWODMW2Jkzj4f+Q2epwrwmJT3Y9YyLI3pdmlcLjIMQwX2ziJkfQ0WL8Qj78KP34U
8TZ6yk5jiXL1T6AhIiHJJE/PPfU4Jkn/QQVrYdemWZws8yNt3F4VnNBSGmVZC0UQ
rSun3vEHK5Rykr4EyiXCjofY+WPahqXwKBEWVjv6jKNvu3x8OMVs9VGg+2+K2JFG
YJoMql9qYFWWImDsZTXnG70dd/JtuDwoI9kFtMLTqlAvcg2Sm50dzmj0dWgoqpHg
CJez+b03OGZPQY7FoVR+iN4C0AtlNSarHhpI2VifyEP/NW3/UHEZwzzDXaal3LTm
c+rrGBV0nEmSUIn62B6HbZtclJpyo7zgN+a2gTIiD1dLcCGO6FWVJmPPkEVk/9EV
Y6poWhROxJXDx9zz1c3LAXEJZyslARkDpp746dr0Vw24VFniQdey6c1CpfVsWU4v
92aWkFeejglBoM2nOITS/TOKpKNSls6yYqjOc9JQg5RSGNNGRL+eH7co6WH/x503
BlCDbF2gU5TKCW2xO2zlRI6BU10oyJyoEQG2osmdDOpi+lVRkaAtbka0NGiT5Dsv
TjOrXmuRXIp5DvYKqF3OTj6yBU86C4EHonTtSMnGgaGOzFDE4zkbcF4UVTp6kwnX
Gv+innBWEge8xYIk/0BR6oP/aM2OvX7pC53MU3Li8lF7W8CvesNep56sJLHQxt7U
dvTfzEXceW47oqzW9xncUczSApG5cXHWdl2/Rnk7/rVpWHI/KfhKlnCsRZSrrj7v
wlWjDo4OaONJE1eYSy03n9r+0uDd85pswAeeb+eABhOg36SKzPTEX8kgxIGBqHh+
9tHqk9rkQX+RitXDZ7TIXf6m/HoU1YnSXPPBB/HCDkViaTPKWqQA8PQ7p2D2IByR
tiQqANlTo6DujenwNqlVN/l2bJgW9sJBXGbeMhKn8+spcXzsEgfTwBntDa1oYFuJ
FJrxNJddFcqVKEwNUd5SMfSUgvU9XMQy3SjCFBwqDxhDYbb2Vb4zW0HuheUtgeub
1dzxBFfgGIkdJaqV21164hfbMohrYpRGLKxW/JTXsnedsEG+dBJv/P+/3JabwfUy
HtQqsFI6xXw/32zIl5/VEE0n/Ih/8SBgGsToiDnjwRb2DMRbaCYNE7ZGvoN2jpQI
Gxz2XdPeNW9IlPhX++ez3mvRIwOkssgIJ0AlOE7gJx3VouOEpxklP0IVORxuMop4
CZz7FWEuRdqNL5IMxtxw/DAg8f/zpTXS7jbGWuq31n6e0TtUzDpuFVdy92NPTwuk
y6tPjBL11WMQuJBEeW90Nqr4SCNvI9pEjGPwrjvqbwhYcji6yIsrHDrQDzmiCBag
y9UfijvpWE/zSShdFyLbPwV8HOhqOY+PlJDrQPitViOWcD6bsPBsmhwFz4VZwRG8
BdfdMxJlHnzi65QWw4wlkUU65/9nUpZeEZ8HA+pzq1ZfGuZegV7i/T3d9CRASBxi
G5GNhFZm4tAqTjVj11Sxnc1Xhkh/FA/SFMmxoV9RL5v9qULt7h1vV3W9PMu+MRPN
NgLNbzC1Bfe2BZb68ObPwMowsIK0dyUf0Xcb6n3852HB0XtkktrP+1BCuv81YnHe
iDcrL8YS6kvGYH3A4THGTv3r265FJ2aE8PUq8X2tvlHgVRyoaEXCkcfcko4VeOwA
o1CmLxzmrsPLhBT9zGZsQU3E4JR8t4C7Mk4xpGCuHZEWS156Smbmq76c5ZPO7nqD
ncUuNVmouWoI2xOcL/T2utYME43i3LuX9G38qE7MuP8WQ2BTKS/rrNR8+exmyi9U
41CT8rcMsJMSNMEman4r+AT/hfI/BH6l6kQKIyuvT16ftcR66d4MS4CVqDwEBTFR
85Yff6sz5VzsBx1FTWAXCRJC3mo5Amp83xVjdX6NOQs5TZeeNrQlWPzVqlDAJDrq
2PpP0BnfdNLa3N6gjrdWIYR0Y2BRxBy9npXzdOMt/VoKUIqiBFzij+/6jx5dgyve
Jqi8MAWd8MR6TUjCampUoWXy7C0oi0mqsmz9k/dAjumcf8f0U9qrnfFj+aU2+H/I
XD6Xjqik7Z6MjfkidJKpLA8sq4qu/6uo0NGBpikAWFAZiTXx4cUueEDmU72XEeyU
3Taw8bjHrYX0IJjQ9cc2vpKku0f3qK+C/DdvOLfDeFcOjr+khMSHXlQld7VUsbfe
kWgpy1I1mqXkWJUXY0quk002uW/1wD0lFRpKwgbKOfm/4+/Uc1BBoaZpaaK2B4hL
p51x8S+e4W5OPLGg5/w4tD3bsbvEEYq8BmHIroJKgrOacoxxLzbhTrqu3cT/Ntk/
V6Ry0S87PdGZM3jzcvWjpJMCfubEIrUli6vnMXQReKmX4vUUhzTNwRZjXcpu/fgF
/P8BxjLPm2UuYyCTumA4gQ0koWhbBjVM9KjQtONaDSLPK/MQaQ81exjI+Tdi/5rf
fGZDoNCNAZwwvhO55wixyLCJyCw5flwASyol8GDkzezYjigE80tE+7F3+q3nXJB2
6yQkiGz0FmMW6ksuclzlLqt4LIrhv2QWZQZ5DwaOFMx2zxAS/yQ7M0cteN+kg5UH
PVwoUU7kov8IJLrDuUoyhLdWley9Sfek4F3ZwdzIFdh48oK0x2d2TkExQsJQP320
HeqqAg/enDrYaD5z5Jyei06QEGQ67ZjKWwU6BFpuPPN0yEaYpVPtzyNUQ8WlSgox
qUpXGUSBZOSFn/WZZPcBeYBw2S2DkruJWL1rk7SIcc4j5R4Gw4J5AN0bCMYMWjsn
QVY4VGXrEnwkbzAIARFfTPUHDEGwGmqjGoat8y7tVQMy3WjvwhOT0cYxKOB8MfBY
wuKNVyTbj25NXwf+gYi+uyo5HSkn0cncSD3wS8hIsYdyYl9+bDq8To15L7FXBeLU
30QpDD43B849P6+GxBgZz6i6UHlWhUWfHcqhjYbyGcOT4MWIW6OtmlCWEXPe6otU
dkQVz58VG0Wf6/RPAM4H1h7oLfFIueBd3oHRiemkuPkKO0v7oNsIqYtDQG4H3xS/
ctcWYJJ7Y3QNUD4vJqp9eQlCJWwWp6xgV2BA5+afd16XmXhLwCUZ/F5bUfCnKaS0
STkXK57Hudd+CvaG7Q30GoHZko+eHS+GkMsaV3hOXfPmkWbyHSCnP5l/YFK9eHRP
RepvNfErJIQh7rakjnGz1V2Dq5B3gUXxorY3eN1Mx1xonl4pqifEsnXgg9o5T9pB
DnHlWAqfvM4S/b/sDDg/bC8VBme/Xpf0FLbU77Ufyr8WPzev08tnhI+rmCCSk6lr
Z210jN/63hlmJlmVmMXcynUsyDIxT/VHFnTqOXGno9ycydoJWKxEjSUgC2IfcpL/
5wrbylqkpI1LLrZtnDkySAXx602xNqH4QL9u1l7HqtbGU1Og/Q4qlB3e8AtUgM7q
WQGq/kEUT8Ufxj6lT8KMrqGMaVYMf5Tt5iw55MZ44cjUQrZMfUNWGABK+rBOwYXz
/TJnfVSDsNosfw4J6AcYyTGWT8p1qrE4eyplouAHJq0dtDSVUkIjzn2BF9z4ch7Z
pDJFQ0tItb4bv7Q+3uRrJonErUL3DqHyMtLPMGrp8I0/GhCdo8Vz2GQkFyuHBwOa
8dt2CzoKB3SqYYwmfRm8ee6xAaJvZnoVnSPkPoiVe1bM8FclQ0qSTgQLoVBx4U0w
v+pNyTKSjvEK4wHB9HQxjrsqu49ur4uMFTEaNz4Zb6iXxvRf9WIpaFKL6k6XITI2
nfsKd5dIST1zrrhZdK4lhpRK9luR474qxIGNkeFbnTdsVn4mF7/TYpGj43q4aejs
oJphMTU3bMDZJhvSh0jBmBwFNTEIYTp9Xp/yyBibQogfrpJ3XpZsFgYHkMISurY9
jzzYSQZE5oqEiCtBoIvMP2u5ARiciCdqH8Pz9gRhx/i292vJ5DLT3L9i1YxxokRl
2QnR3aKuuahAm+2cWe8QrPGrU0YTQcSRAvrjdsc99/WO8rNFxJu8pA8bCyP6FuOD
J9DPP1Q2XcWAVAGFNtAPKWEwhhDtr3VIce0HP7UdLj4dRlKvhZQ7LnIz801Hbv/k
f6pM38SzMgVYWYk3dmVvwWkG3aBFdnJzq1I414tFi5xWSKjBGr+wF1iG/yE5oVfX
lOOdqOv3TTOVosap6LmvmJAnFfmBfxwZ2Dj4SOhvDfkevpls6clcl2K/TDMaATAq
BgrOu1vTzoYgBj9brzU6bOkn+NhWJ03tWm3p+jZ9wR08vy12mUq154gL3ah1Fj/f
Dg0S/hzx7XXtXgCY2ukgh9BplWLUbL7ulUArxP37BwofXZVj+8de3RxPFHI004Qz
mIeRBBbkUSS8IxelDca8N/dITtazwi6AISqKHcBRVIFRA28xGEu9xtjwhm++7eAq
xBtDHpQ3CO4L0KzDtJQ4i5az7lfO6HmFyRXPMd/gxswJtLD3nnWo5n4nv4mKFRqC
flVOGA3SC7fFco84m4Kl3fIbzGPFvsOigBRR+Pff+l8uz82hu1T6XxT71VzcJtd1
wht8tiynbCKzABytZFdL2P5u8Dq4TT9lyCs1TUMV0AIUOJ0Vg7TpT1UA+szzeYdx
qskP4A7aQVmiaglOE3iScwmL64VinMXMuC1Q4Qx0IM9NckfQztoSiif3AdvPi9B4
qtgAp+/NFuXB3H61HlIuNWWmXAzW+O0bdPcsZ3zfp3WZCGP4H7St7GGzvZm1nyun
oUgWKb3GcbW803lm/2GFbyHMT+0d6EpzGIGEPMd98IISENd/b7gzL1aaCkCTsnzW
8eGSoweNd7OqZ39gOIqF1ZZKmqJu3G+eplpK5/61xqDxDMy0OQ0Yx1hxPa9hu4p1
F3tt6r1/vR0dtQzq45MT0OBYI/0i1HPFrOGHCVu8dKo0egBR64tU7+ZnQZ/DsMw7
uuIclDG2+Pwur2HDeePHw75OcxAw3ZsMQk82BaLqRzRiJSC6V7w5piQNmMbuvfaX
gvDrbkh+WzhhX7Un79ivqmKeMuzOvmeuwXYzcS7tm5YGuiaNd/RIFCb2Eg3Qun0g
caMLYnI6PXcXNYXnK7vkWjyN0pLUuAxIsDORW92rbXXW3ddwaC2qk390Rrl7SSyo
iEW88HkQflcGtOh2AIAERV3Jqr8NBqCSW7HqPrpCbIGKLYsFtEhvaTYEN++8S9yl
/8A1Ha+V+Zv33rWV2C2OiDiLFmS8qbBh2mV7crgVuUCrlPu9D/9e+aROe6lRno7O
46Vf/VKr4IS81rlUOtO+M/awuCWqC9fn26HRpupFHWSJVfHwRv9KOdAEYEw6745z
idmFdboumPJg2UMg8nPuB2O2j2CZxGQJh+HWQkHQFh7cWl61a02q9B39kdGdoIcS
r04lkXNsAYaACnYfnSgouhrHqC7qW3vlEZkQYzZmjU9MSMLX0F3ppal/oZi4NjNf
qTsLfOMxBs2TcVHPLUjET2SNQViWn2+xYN9qC3FfGmha+C7kOKvcLqEn3YHXQlcP
WiXOscQ085QBNsX6YWZ9gdVQI1G6GtgTUdMKQ+iuuYgGqgBXgYpuNpLsOn2mxSMi
+qEfCqd+CJNOyMcfjP/LVp5d8YIJI4Qwn0x8E82HDEttHEIrVXlD6L5pfQYHAWD9
iLWMsMe17RjXs/02StCAteNzW27NGXthBuVjmQ6OG7RaOgcyUwKWCiPfSk4tGd4L
7BlmLclhlOopKgG6RAsV8dAN2f7byxnoLpHq4iOgiHfEsrpQ2BJZWeEgCbpbPbgI
zJ814Pz+tsoSdVRjsyRmaJ2yJhNM9FbOHovgjgFUP6zzLuBIjPOgojQgYJO63a9B
KI38TFNG29FU+4279UexwzK76ur7etm27YICwPct5gx/7yBZP3S0dIasp7r07KWw
Sjrg8HJuSQeRLOFSfuhsjZHrYQuS4UrCYpZi8v7JTf4XpC+ZHKElmmKC6SBV2/pO
J40IHtAW6KFYvFMUP0FyBpSb3l3xZoaxwirZ8zsH4UGRFbWaGarraCaCf4a4kyj5
0Xj6RH9Xr6gSvyiz5N31uKoOoUs4ZPKmkX7wzd+HTK2imVAiGwpM68dvCSb9i0DK
s19XzPoSRAridGbQj0riogsWT/uWH8dP2gz2MFIZDTS1aO+DHcWA41lrRPyJy3fw
ofjW79eSwmjAKlngCO2FBz7YUN63jyeWLH+hjlr9d3MWLcR7oivWxmypNyv59APo
AXn8sP60JtfyrB7DlSyCMVQlSjzJYnU1vYTblxDWM747RcDLBBrpZ+YcOSkMbY0y
CMr8c37153LD5mOy+Sc1QJx22R7cGFeEVpogJ1d6ZqF0Ht7xb3Tjm+Gs5HM03WS2
28g6idC/T8VDn+jh9vhbgar/LAqKMJtOUR83GX//youQKo9EeSH+f9yPoT/wokAe
IWAK2cycH3XQcR5ByfKpvtGiGM1L3gmCOeDEUw6DZBV3NkTs5GCKRuEHolR9JDU1
z5WNCfWqem4StIg1X0yCI1SFPFoA846Y6VtnwjsypY3qDVYi74X27WKH1VL/5Y97
jkpHqgtIWpoqKBL+6jH2u9TIk4c0TjJFT8PU6dR68d0JMlkf/K5vc5Ux4WnM1DtI
K5xgcaWhXN24Vpm2MlROfbM5WBPNXToksfmAqye8UYZgcXEgRzcgkjoJiALz/Qpa
LXLXZLVadET9fUCymPRv6Eilt+I43QrcIGX6+ZWd0w7TX1N5oB+fIFGXIvlKpxp2
FFXudAhT3wk5sBt4A3e0UyNQQjfRALZ3MHRTR7hpNg886B3+g7KU4LelEqNOkwBm
i+rodKv/9w76+yM/dd0cF9lkbdA9wLRKlRphUTdS75pP3dV4UH6WrUt01ezhfAWc
Tanwp0drHozySeonsbONK+vqbe/H+2Fzzqwkb+NJPfAj/KcyeHQP83tGjrlfYLwz
myKnoebqxQn3o8g32Yv0RA54L3vJMXPi/yy59IMY8ohwuakXu4IvqckEriOYFJCS
8vKbqVAg1prMZET+I4nLP2OA6bdRJoTv8qcGxX5s3i/rLIEhQOvbaIXgYA+57X20
/GuXmtR36yt6iwxa7xIU/LJRiaMIQNAjVGLo034z59vvGNuSSlGoWh7ZL1hWByVA
07VqRBQ1nNf40ivmzb5LUuKXs0m9Tn2adbVmuHJj04QyVJ4z+/3EKmIv5IvOmNnv
S4zzg6hdIDfqnHe8eBm82ElUUGJg5CzJKrSMioNopQ2uUgUL3iifBvGGLl0qQKGI
VteCiqEerFEbcdFDemJhGsSLHo2xI+Rj01gK6hjvoo3nmb4TEAlaJWiGuU7quqDK
ax0u4mrA0qJWNFuBegFDvlbzLckC25PcRD4vMUDuA0XlO0jM18PacX3iFN6aQT22
Eyfv5kl77TOmGdm77YeGxrGsdLclQEItZfTNjeCdZ2uO9N9qDDEeu09peheLXstI
AT1WkMu9amKUVcUpvu/gD2e6IKVWC+1nMla8e50/SfwKwa/22vlTRi7pHqod9xv9
qprIAcvcRjAeskhnDaYOkzbr4jO7dxKT/iqR4ILhD/G5enph9l6ThwxvdVvQXQQY
YnLomteFIYDwyFZtsyzZV9Nn4DKqu92j4/IPudltypAhSrh5iO4TQjiEmGUn4mXI
gUEZe7us7BQqTZjXamUGJ2mG+dAsUN/EEtOSiq4fgpY36EBOUOs1xSgRfel5goWC
Pzftd/O0+JngbdemEVvfvTBASClbMzT/1rtstCTwzBCODoLELpIm7ZROGY0cWXJq
W8dBIyPNP9H5bs+/rcnx7F0MHEPZdL2mMA4HrvODL1zdI0TgXSaCZtiyPb1CexEq
dAI4QBnzY4QhB7ZT24xguitjnAn11tdJACutQqu6BFFVFMmqrSwKM5z4GZ2yAD2U
rA2T5x8cBbF0WdvCLZXpinWwk48IPDxtGRl/uxJf+/5QpmWG9qfRRADQj8rPNa46
NUhFlX6PWtBgnqBop7fbw9fHMuAtLbNHckgdLPdyK2RUtFh59hyIPJU68xNk0WEr
6cDOtAVM89H/+dBOsylJHgcdWctoq27JJt188Hacc1W/sDsbZseTetfy6sHYeX4l
zNAtyzOxIButaFSEP2MMwzPolkXVjyaPA6/8W/VL32pVvnCYFlq6hSwJqUc8XobT
AVqjUB7QrI+5wK0uTOQ5huLztrHsTg1FTm0kdqQ/rT6r6cw7tOA4fKa8DleOAwFv
E1aMIhYfFRTCYcvEqTbhrtodnoyjUhTvsl7rbJjtyFoxPVFAbKH224SgkhYjzzxI
wgvvFLdjfJHi8SCc5EyEXh7syoYWUWf3BqBfZrfrhbjI05eBkwM/6eRYEHKFOHF2
K76LZySEJUGlqjONxznCX1cjvGipwHVEGStoE/8Gs5RpmUquiaUSbOirHxubmp5Z
hfeLmsV5pORBRS+Ilk9+wsrcjCv+7G11wvKqsXWdvk4tX/giXWd57Ob1v9YP7zYV
8RkjW238s5ogJ5d0fYUFUhgw1Z8dFmkUQYzV9/W3e5urJc6DBz2lvppf91Tb/wLf
RoeKn2HoEc5mMnittCnqIP6oz4mQ0aJ9LMwzZFUHP5bCjpXc+4c0W1T6x/Ua5osm
7vnmD4OpgOuvuBmROokLQoxQPtRunuunVWpr8Vwz+MIp5SfdzUcsMqu6dROquIwA
HyYF6Tbgpoq9GXpXVlvBZ8iCcyBypyfkxRKfpl2SZOhxkwrcAHS569AuGpLgF8ed
hZTWgMNqJJ91I9umQjLrmJQn2/Li8U86bSNGkx0LHbF6IbcvpVUKTmyLGxYTLJ/H
TRaNhmrN6U6yHsZTDrW0w20mJYnbTTddthEW28iD//5h19UMONg2QyQs39J5153p
yT54+50Wird5duCz1CpfoU4tSYviRrBrZKr4Uo4yJdP8xxPBz48yR6VkPfCh3DVd
xxu8FKnSdgXSk9pL2ejdtHpyzuURpi2oyjcenOXYjWh9cFRlXua93SVjTrPcsMzY
0R5m59Dp6j+Ao8QSMV4hCNLH4O7gpI/UYnVYNcdM+NhJ+gTZlcK2/tSfjA2+onuK
dR/vU/Uz7J+n0u6rMMOCIrh+X+xVTFUYP+1zys9YGWlknTCoflV3xjQ0u0LkXzeU
YL3ME/lXIgB91hjgwDbZGEIvmHr7nx978HjpRKvFOicuw7RKFAtxGiYYvB85HJZh
Pronk/fC6SJdsZ92WziUdA6ZrqA/GBDKhGL+h5b3H5vl6seM7PHVZ5RUBE6dl5By
+ns2dwQRn5Qn1uS+VW+zkn2X/qgqdsAensI65MM9LHoExi/4jVnHrEQALMcrw6ej
DGQjx7xQ3MY0ekBaS1ORsngoG84vcoYffIyzZWvHFCLDSFtHPwuz1niU8xpTBl1t
/UbGHM1uOmQBtSughpj0breaw8vH1BrmH3HzqSdnr8EUm5eoJVDH8137rC/MjTww
Db5gaZKR9tzQYaO3YuG/3L+BSqA5uinTdq+YrNI8jLlh//srqsiuAkSCLsqzj0Rf
fLjgAgBfQGIhzwB6zV8J6Y7/iDvNGKft1JuHnMG9jvrcRQpfboAGR4idIWptlqjn
1y+Z/If9MHuWxyn+b7i0wYWwpuaUEEvqRSHqNhF6vRSDGjbo2in9jPOUjDjlBPCj
2MZK6aPgGgmK/S56KbRac7PI9bCX4zhYvbL6c/1bpUEbvRqfnmldcwZy/tlaG82m
W9IBI1bqVO3FRULjEv3r3baFCa+gaphG2j5cMJFo+0kQuWP2L05D7FlAEDzRlriL
8IKe3WU68YzE3s6wA+0fIyO2hQYmet/aN4Fh0/RMskMUQy0TGkUu+XAuyrohue1t
f0bsB84qj5zIwbV1ov80GTlKCAq18YREgPAAZrnbUVe+nwZMcmDEMemYYzfUeGdB
+S3eAzDmYkljVL1xXswZm3xBixip6jK6oFbNxMv/JgzvJ61SX3jOu/loIlLamL7T
4QTarvtbNf/Y//0UCDiqBJ+DfIG9MznSZJGrBt0yCTtwR0QzELlBN5pT6YP4kXNd
yp+Mr6aap0AQuLH69IfjcpCgM0jkoyw+moxhsrdYdX1H/9iQ2D4YeXHakF48pcSr
q4/qmPThquIICA/NgktJLsFFNf4GYC7VMp5kNQY5yh19S6ciPRsVTypGFbGnYRYa
lr9Z81Nf0jPITibyHJFtajmRotsrEvbfPtjWxgglOlZcMJDS38kPoGHO/1Ps70AH
OLjGlBojhWXraidFbo/ma77uNW1L4z+P5GiCHmYKeKpZtQyynnTCFmazPdbua2Qc
sxt2QSCkzYMZkDliFTt3lD7Gu6+LRqDPotNaVRpj7TmidYRjcHbL/n3DkGJD5GRe
CPd3iacZCfqRcRui5iJy3pwKV3SluOymu0FFHulx79iZ1GGrUUlBS7K8zOvsly4D
I7H0c/WfmtVgeAcm7YqzCseuvLYv9RcFFjM2ixxr3FaCMZTexccxWZtfnhoKGLDE
JvFlR8JglbXRT1tihMJMSxxRm+ZpTmmPA5eXfevpuYePhDr3FpcZyowRFPNFTZve
HhMkM8eORAP0sFjqRw9Lrhq7RlCCT2CTpZe6KCvgJGC7bBQNBFf8Y3j3YIGGzuNq
ZsTU6isXAwEcI9MoK8Lxy+4VMFqZpH+xg75IkBOcVp9d9eonSyk4K0ipqb73MK9o
hEvCYS+/w3kNkhOr8xKpkB/sIbuJ8hU/OWOmfr8uLxdVWhJdxR88UuRRDg6gUc2z
7ImbtsDvFGWz1Y680pCSmBxcRAoxU/zfJhVJyTcXW2Nq3dljKqVvqN4fsNClFkc4
SriFnV/Lf2FwMjRzEbV8UcZtE4Dau/iTB3MoJX2cd3hsRAIB12EHCrC3YPdWUMto
MOesGywJsJGwTFJRZd4c3IwIQYSbWacotmZ0pHJcf/u3IBBo6/NvG4wlDENDHFGo
kVXJpLDcwzXrhctGHRlaap/xVty7eAn6kNhot/aJRNCjpJlt0rdNP+mo6CoS0lI7
6O86HQ5FW03QBc4wgZBHY8s9g8GeNnFE/nVDR5iZs1dr0iSgOb6fDNpmuZSMDcCv
rNb1+13Q4RbveI96UgujEv7yoR3sLGnBcke+x5GiM/EGBADfOeMVvbWgw/vr/hxn
xal/MlNvUhzlSTCeaULZdBLLPsze8Bga8SyAXri7i0/VwMl0qJyvdTz1O/lCBgZ3
j6mMXIkrYBry2AnlaG5qie/DnfabXfMmd9uzSL5jsZ7QIgSkVYA1tJrs/TBFok2i
mjCTRBCsOmWwv6LSUNu5P4HbglIghuTzMEr4z18OKcWf94ySK58Ek3L5QXCnWrtY
lBijJwXi32FLEiBpQnbDlFsfguykwi80eAYG+KS0GWg/l+dywwJp5Kl9kBImEZNV
CLtcL+wMiRoxbVXQI6ZVmF7RwX337awFipXz/t7BovJ1dlMPzcohez8ivScf+y8+
G2M9zGbyuho1U8AfgSYi3OLYE9ks3XjJ3g8PTBWZBZD0XS2/iTy6nwiJYuPvTS5o
AKkKOLX63sLSFwJgAwboTgnjbnc63h+QlQ6tGBNcsWvW+xXkzcT4mJ1hSMGbQTkx
+SAePqeWWHbBvUouJdHAbFhXqVRLF6NVIa6Dgazi/5VsUT5BBzzREkqsFPD0iskj
bG+fV+bf+Qm/iSixuD/lfk3tgoqtjwD/u5dC8RI0ZFCecWe7k6Wq3+c8mBMO+q5P
BFHbEC+q0u16hQSqgTX5FDgokXyFcpI9REh/40RBRQcBDmEz3NEABi3OiNKR/UGI
g1Q1SfqfDYjs4KV1dZt8Go+l4fWLfyHC2d0TysuB1wyBBHd4XyewV0CEnAitZfmy
F2JJY2YPbehIupeCQ/e0HD/CKyZ4tpFVyzmRyfOyHMxmFH+L/EXV6V/0Mrqu4lSw
iYgyNjcGyxCIy6YK0bD3ACZ4MIhFOYyX/To3AGW88ecEsI4k+VOqDp6dUAah1ZkJ
vhoX4urf63Vflmgzf4Kmukd+oicwGD1inchAjwhVBq3++oDIXX/3RooakXtrv+qM
v/0181mac5vBy2lYiymcuiI37VsE9JgEnOsAPMshgImucIjCRkMA0DV/kq2ymNE2
6JDPdf7FCnv6vKvap47TKCsrvbNbwmeMpJnDUpHrvtftDHplwtG4BlnXL3RwGXDz
3WS41gfbOv671gKzwYqx2ZIXVrbUuq+JEDc8S1TSJWlmtzhxAmg1KNAEfn4opvDz
6GECiOFb8iiLJZVg+23RVE2Y2PKx1Lbsdn0SeEM6rDWt4R33jnIOKWa8Hd9CQKFS
Dia6QKQnp8oqGN2qOLG1gbtdYgcuXKvIATxH4CB37JRHmzaf/i4vfj7rgvDchhQo
St2BLGlUnhzygZ7t3caHo9C6t7FciVWy+ejkMVsPN1RVQ1SeBPrtwvkXDp6W2Rw/
g1vteaheq8UI7+JGWJ7plnEchfUB6UUdnNVx8kHPMhXxGQAuZTOdrFdLgdQOGmCh
Dj5cY2gai11YCGGdIdwixyvOakWEMGAAH7Hn5tjY+ibsQzs/J+f32FOe19VSlGm8
2e0cCC76U3ZDqEr7xVvkoeN1WuK57DCGh5g3BIi1z5gFLMAYeb4YXCY1OQWj/nC8
XdHpk3Vg74DcdfNLNLXGW4oDeXGW/aOz5x3HmUxUagQDPLaInXIIV769XlXuwdeq
BAoFCDtnPTRptG28BZejgqyl3KlS5yySrKB/nPxAqiJqe0HZB70/DaQyEW9T8O5t
nZNqE+xy2HlOG5tNUyZ8YjArYSmIvfEtk6bOXBpm0u3RLdzstfrTf2/B5V//8vzJ
jmxN5c1N3ctiMUvsKBjYJ3xfoAmBCUy9GbVR6/9sc8XueQKfbx5/pieZmToVLM9X
1pzGERz3HrImuMTMeh94R/bs7hNf78VPPt0j9I+xPQuzZtMdRg15lz4o0AwliBum
xerR4JgJtwLim34mYHmRzuyhBZDZTgfHRESzhpHYqDo0Rz59ywFf3DgEFnaIXqOz
i+Dq5ZP6aaWL+ExX+5v8/wGMBM6HSrHMqi26AVTS0glWvU6k1IXlmTuytPmD6eN4
IqSx9+PHebBidHkyNEszy2eky9/muaGBVmDwOEKoKx38gtOOVM2iFAs/UcWbiPED
eA6E3p8uTcyvRyuVP6VOj51NbpXnrAeLswlel33IbKAzEafBks9vAxIJ1dXpwbFD
mmQFqZTjBgpISy80OxHXQseDePEPwP08liGlA9VjEd2iQlAKQQ3WIBds2l/FV/kh
JsZpXbqPKRqRo4B6vOHMVJV4of1yNEf5CWkHL7+ACln2hov3TPG4NojvFJfJbDBV
W71kTKzp/sTSSREh2tzYtV3NaXVClZVZ/A1v5TRtIqN7skw0kVtjdGsvrfOUDGog
mF6cjjzQrBkLSp7cmIKtb4QDWf4ycgTu4jQzJsBSrgScNr9M5fo3VEmbuqbMMVnv
LWlgPzICl0mpvowf5/fa9/e+HQcVJTV4380DgFtSRHqzxqXwSYklTs+jf1O9ePTo
/RzjYCN5Ca6HaEeUay6B0oq3M/RCV64svmMCOBhyHki8V6rYojNLufj/3awdHXVF
IXWysprs/1d4cecSQJwJAInW6H6L0aMxTfwJ/+0olgHJJi/exuhLTAiZtpgyHUG+
AD1s8bbuHUNAkrGSQBgxHsYdWHlRC5RlFm2DDku04Rcqo2keCYrE9DDw3T0hN77K
Xo+yrY0063tYNy2CF+i6RP/Vl8bgNK1ZUlHo+RDM7/n1uUF82mFh9DgfHhAP+81t
qmA7VUf24DVQk2c2xoxFF8shrTfE8bEeo3BfPipaVagpqDHOyey8QxMD+UPURp/o
h31zHRMjjdxG8SVWdwR+iC520nnn0YcmGkJM4PIENO7aNM1sdEc3OpgHfOux4k8/
URnqdNtx2G2ULyoz8jQgg81Mp36YHn10p/R5OChIw4gCMfanfj7S+n7YmCvw0yTz
CBPg2KXca6EUazw7YCfMowNSQffx/Do6qQ66EFCVernotk/RMh+5Bef4mkJ3RfYM
oHfCICrBSH5o5HOZkkFssReMlH49RT9U2RryDi7CfwMQAoBplORcfFc3NB7DXxr9
odSyIaRAz/gFsN8yz7QhT0FJ5qw1IB27PuNyVRE2i+Mm6Pn8lIuPpLTopbbegzW0
ZhLu39vJ/R29lY9B6xQOpRvc4znCJ2LtExJDUbdbgeUu2nvc5chuiKgx+1CRQXk+
i9G3FiUWhwXmWO0XDoM657y5/850yqRSj1srtfrRAfZV3/5eumHwna+g4JTbE2aN
naRFjs4hvZg9Xio7Eb+2sLRcC6Kk1p2j9DKJ4WG2FDu4Td79CYVMJu+K1G/xChEU
hExcwOdaZSaRftVEfgtf6kOC5lgikFNB6h64Lf9StTtE+ugEMjhYC+GU+HUDBwZ2
upkuNC5xBBu7PIcllHDagYLuikA0kbwtCpxWsJ/guBicMGBBnZltGJ7zJ1ff2ulw
YTFiY1EUODA8KPqb9ejv91UySydHh5dusXEWGHpQHJPX++JLvDLB9zMkYl1Rg8yr
LEspg1qc7cHFs/3HQ+zTC1hMpNbVNAlWYwekJiIX9bcyyGffI5xs7nvSK/CqWvoV
5eeoX2ynvrF9zSN6XvSI37Y0GiCGTTfeaTiKBv4hh70WHGWonMbLiEmjhZRbhgHa
qodYcvFW0ChsFbsxLEwHuZXOva7bgMmoNr3NdtTiM83J8ZyED9IeMH7i+ce3cNTB
IS1c7hMn3qeuHg+5KTBo38t8G4V5sOioI1M0BD3FDXn11hzLKVCqJm/j42RaIncb
QF5lpfhfgxdt5ONVNJ761ZJcVvcQ29ua/XLwyKuDIfDpTTuqCxg0siTFF4cqjQO6
vznii9YRaa0Curs5sn7DPMDkH+eIJaE9D+FnZvLuUvgbQG+7wC6UCnHoGhJzncbH
l6OEDHvoNKgU6BOZ73keqkH00vl0vseVGbiB97Emb4vo9wlShy5uvH2KIah/ZKRf
gAx73UXPgv5xuMhSyvFOAqsRQ6W4QELEOF5zEb2R8Pd66HGN1UhJL++zqU8+fHa0
U6QPnkUUlLfYefttOPe+9qgw18lNofyGL2j0defNDSyLlnAFRPgPsfk76uCqa/Rn
ObXWfPxEUPJ8oYeTE+P5yT6bV19ewboOE8USR9noV6BVI7jcIlIZBeQOQ/cDDA0Y
kJrZxuAq7DLHzE0p+b79yb6NXVk2Q6rLcJziNy59s3C40bz4XQZzp9E9fF81rhki
em4dWSRtzmz3epACr1sNTFDewzXi4MNnYeLNyptw4K5S5j7MCipOFaoTPsUiThqW
RLQ76DGSH12W3pLBiQrTHEVIPPcb7CfE1xR9gHRiJrVSJgTF+iCMvz4BEtrPveEO
YO45vikR6zx6NzdFSDG6cHHP5W8xiDlWTfH92Xa0swJFbVja3PcOowM7nxa8wyow
EcdQFGaNgSDbseXL1deGrF8uMMfIYIG+LvYu4vttHE5ZwqCBmRT3Xx+S9SfSOg81
lrlU0hVucc4wyYsTZ3dU/1SAiBk2hWpPDqX5zGpDyVoxhm2TlhJ7oYLfgBZJVje6
3VtVhtZSnHvmSGeQGwfjWpYD75rZgWxd5piGpzeRVGRqppxsIl2SvOa0bnEK693s
BucKeQvTM4Jer83Q9Fyg1rmhyvxHbV7APX2Li/Q67omj3uIcSTFfKepCQ1HwKqko
bv7e++tUAKku1g7ZkIlfVRCHcT+h9VduDO5CVSVQmhzYFXz/cB8xzSq2VC5lh4pO
JBEVL56FutcmkmzHGDfqRdTsqBDoeGn8t7JkS5szxppurpipgThaRtUX86fuAFlS
AqNUXrM4f0boSNn6WVKQqBXpH4XQYm2keXdNXQ/TGA5uHyT53pJVJLfNKl7jIwBg
e4kVIZFN8liZnT5wu9Hvsk5ZirblS14cfWLy9myzi2q4yjwwyuUCy+oNqGQ/td3e
vqMxMlBkEcR8QxSCRb1PELCoufRREbqIlKemuxgSgd7fAkvo7IKhj7SXMebv0CVp
Rhgdee4yVTc02qUXkBG6xJKg+hPQ8wG4Kdf3beBgqddAxIuZ+YThTuqE9v8CcFVU
sL54AZKWRbwZ5oJXjFzfFzvkviRMWM5AOiX6+xp1faYQPiEQviSrSvTodCrTdIZM
cyuq7qKg5ELPW+gW2V9o7SRKWGEwAD1Jf5onVJrONottEyPs/o4y4LogPc0MFmbF
M/pVVLwhEGY80M2fcpMHyK1C+EhZb2/v5skne8+K1CayyMHIFPqgn+kmyxF3ARb2
v+BZ4ofGjFZ9HTWdWzEr1/gqPTg4RTN06RFR3ZBDYno8fv6ggexNo491VKDEShPd
oNapG7HMd5B15t+cTg/JIFBoirLKmMMZ05XEjRiR0CnxCpJr+Kn1sWK75Z+GfxPa
WHoL5iOQQR0X0QCcGGsj1d/fhM/XhwjD7zLdLpDi/A51EwA7/M6T2kLDHv5YoZiK
IggWdE17kB3xwJMOxY4pd4IQTgF4SFCoPTdIIQFfTdWjyxY7B6ORl7pO05CJzuuQ
g7w3Q3XoFFQGe3R7Jf13lWTeRQotHsOPHX1pVT7WgkL7/RnmBRwX6J942x6TVezH
CSe8FaKkg4rqBypu/caJseB3jGUQ2c6I8pFQGJMBOkM7cKykrfdEnKv3A/rUCwoa
a0Foaxq4ncL8TF1Aa05f+qU05jd/wYT2GXcDoJ9VXn/XA86kx86vJ+ct7lyCcfOx
TuFngFvK/aSo8vmRecZq9VZJWs0EzUJeeF2Sd+g/eV8zv1R02c+8thBZWfLe82cm
cwXweNkcWF6zTNL2r7/RICSXr7VkkAr74Me3UPtB6eJgTNbwdFqOMWCpVgzdeGFv
1HJRqj+w1FPCGg0SJ5lS/BhovA92KSVSoTpuKnBRBDC24FtJ5/6AEvo13z6bLxTO
SpWJVwxmMbHZNZHgsZ/xmsQozzyg2C8K2wt2HrHyhobmIxR73A4zLvyJWbt50GFJ
aum1/uF5hXFMHrsIG0fL5RYPeVkDsQ8oWsLpzNleU5UL732afLXqlDRPJUPGtDww
NunBCrm3mu7a8YN6dXjAY5ugn2p1lWyJG7PcXwGcB9l0xCBFkEPDOWiukpJgiqQ3
ceW9fu9fnk34wMKJu+54gsQd4kLvm9T+XPrOxG5ER8tRpcCWaqJGaaXtQHzbgphh
ECOTx3jxc47uCOOnHQABFUmoH4tclvZZCBH9B70ykoBIleUaFWZ10N/EXs7H8P5W
orVQ0FnSVERKk76I97RoQZGGNwMVqU62KfbLHJwsjgF4TOPOaZ4k88iqv82P90DL
uhGIIr94QHVq+JM9OG2wKDcyWD59f3ufqcOlLR69MmSrjRbxXZXdNj3ZFZriHgqj
aWUIPDVcTAYY2PB7XIQr7V+uzx+gfA9n4AVOv1UyYHjd45oJhTTssYbhPIuEJ2R0
2B5shDKYuvoPR72uvjvhoY3lQ+ES0lsBdvkZHmzdGqBW21mO2IfJ2z4RLDVE+6W1
AKxLul8HKUxpKHjujR9URiVJRF0ZC8B44zKv8VsCb4NO1j1/+XCSBOvMyyVb6VQV
0WcrC2TAHY3nIftoyTfkQn9fnkTMcT8hhGTe890RjvZ8aLzspXB4ki/iAUNYPl2F
EuH8h/06/Lk+8nQmz6OA5ZYGfHZ7K+8WzwWg35ml0guOSZWvBgmq+SLw8yCJl0Zc
YQFFXE+aTIn4ZNmXWVWJ4lagT/JNQ/UStSKiPmzaQgS/S/NIvbRmwFsuxDmEXXbB
NObvYkpfCT5FLps1KzOZnX9nGt0g9RI5g5kt/R3XX3gonOCkOPr3LNmz45UKTWmp
xZLfhtGsPZkzIg6X5P/AL5VQhBsBeuG2xYkt3pXsIEYQg/o3pW5enSDP3Q2ytAA0
DJf4Fb+RZ/qU0EwbAQBXVn75U8m4a3VDhg5J3DqogoFhbpGDy3TRFAWrpcCbsZxr
WblO+wzPz61E26/UDKPg4Zkj2Glpaci/K6F2Xz6cFKx+1fWjDlHZQQg51dW8VBFa
aeblfPdBa9DLKQKTcEwaZrjLioYIWV4eFF0eDlgtLdZG4HpcHUFmXv2WrrM8fISX
ZiUk2ywxfJqA9XejbOAEjEB2PKFKoky6yg5GAnCkRXGCASLXjM2s1hQKLBE7tXPa
uMx36+8gsZKAYiJBQ04fJDTFPk30IfIKFahacrJAFEUk58Qb8oeUykIVQ6wyZCmd
OzZX2exwZvASDKFr4goGHnLsCBkswe0F4rn7PdVwOtZjmPJQLYkIr4cClBreDz37
I/A4JD25KZtARfaSQ2R9ljqCDN9HhKhm0LLdNMOTKA5P7eweWL/K1AnEMJpfCwDK
kqEraDumxsa9Zoc1BE4Zc/9Mp0ZToCHyRVX/vnYkcg/TUuz6gdMx5qWalP7SdDVU
NriBu0HBQIn0dEc94B6hZSe6dhlfbO8qkiOZE1SIkxlQehIhRHrYCD+JlP/7BNXu
owHIe92UCJuhhI+bOHYK4gLMVAbHT8pqIdbNVMrPro/EV7UZtT7HydS31/tWiNQa
9h+s77IdgQ5TnyUyX0LAJ4GkSlK5Bd5oHQDjZRG5ve2RUh97gyM1XZu9si/apT8z
jGX+ZsGngQ92dkzuKogvDBi16BX4DLc4+9YhGenD+AoGSBFH+cegPHKDNWyLFl4H
xen9zPD7JcHlhtIBKl10dCcU9miaMHorTUCdFcSACzS38/rKrTInx2l6S5uEPvM6
SXJOovcJqoNrphdWSB8TS69eDL1mUVjA5uWLB3boNcxvF4SaUl4M7Pu0X4DSdGYR
4CYN5lxqAjH5L9onhTy3p6niIPvUZ/9htTyKNbsLnarq6kuWQdHVwDl7L1LNjprT
m3JsSzEWD4zs+5lxS1jXV6Claz8HCTycuquMrn08mnwsKxhE3+6K+eYE1hFJXoCO
lzxzIOLn6TaI+Jqkkx8lPiyot1rwsVeEI22jCzn2wigF2i+se8869Qh61C6ybWf3
VJkou3FMtzNVZ/i5a7DEdNIssf8WQbgmk1AUvB2rrNoBT7J7Vs1AT8QPg+pA8fDm
jUTv3LHbu34hC7PYPLbbbhbiPfcQ1LwClPnYWfMv3dYbz1KlJVTPcpHFJDa53yxf
58y/YL8Xcc5obq2EZHj57S/pD+680/fkaPydArA9JqP7OlQ9pD9CbcQBcfxWHFlL
3oj/zSyYKLO0YSy1hKxK5VyuvfuLXEK4bH9o/C8ZPRKGRDBqtURk89y9yaJ9kpn6
ozUYaxehEIjss5DiO6F2AnadZgd6Bw80zCE5hgGuk4NlY3SbQPZdRM+Lza+Scyxs
aD61jbAlsM4n4PMVWuFDket8YYrF1/+jCYJ0Sha1cGUccAmpfxm9QwF1dAIiZsXZ
TwcWPx75S5HQWNWW3EkT0sgjM7CS1f/4Fy0+Sxj/Tk4N834T0UEN9JamkzCemb9Q
jp7SZ+GXB1kdZLEa6dAsMVPjxzkYityMBbVs9EvzMfMfu+hiDh8E+UKRBGiy6OD0
d6cpZIFvcayVMpIT8z1yfSwAh2ZY/0qvtvVNqt6nEbzXFt0FhZb8U8GtTw/7cRn1
xsM6257dsVbQ4EeNwZocw4NMkk8JvO3dGbUlxGcg++O3BmlddNO6dx9AUIvLJOUT
2Tcr8qMm+mse1/KzsEZzWFcBNgJbj/Fi0NZmK+gXQUmlCHKct5v3bn/j+SOt10bU
4XoSeagMiqPG2cR0xGv891lghakcxUaweDksjsEyIJ7xndzZZ2eZKAVg+NDxydAk
iFb3rOdrwJmUxjZqRgLXAZmM+7tUBHqcoWUebiEGy8B8yVFKpU12VrUDdHBz86Io
1duQUDwxxWxWxlL9YOLRgLpkzFJGdlm+U/G58BL0kEG6r2nEU/3Vk3gUFJwGUuNd
ukLm11L5Q7UgH7hXlphvwZkzI/O5zEYp8KyO7a6iWgG+3uXBJW/eNce39EYJNMZX
YhhxwS2a60PKfxWfuYbh3hkoGMUu1j0Y5XpjWrAQpaUZc1Tl3VtrCdpt6vaZKMIn
E8hsseloS7oqEx73kBbzvu6pd3lkXqMz3Yw1723CcPCP1Gj74Hth+j9bb+7yDTFI
Sx2+fsSSZVLSSY307rzXh5rgu3IC4jx7Ubn3OqitBxSFIaN2ny4EBjA7BqWlAFV2
FgvDfF2aQG7UiI5zbS5omr+Pw0G3tAAqES2p2/i2SmYl/Dw9QAXhIDcBMWtMmcmL
vBztaXypLiEO6rQpHLLGcV6PK0ZqeHFKcv98ExuVuhKitqBVMQ7xwwSWvYJBbTPS
JgiTXMY89JM/OEB+eP9mtAoBQvj+Ffr4XtwnywC0XsMURQKtON9IYohUmt+yyFlM
U5BkyV9zZmZOujxfrYQvxbHFuRtqTltCRVBXiH3MKReyIZRzuSyB8H9wDneWyIHK
px5xCN+6jTo8Tu8FyAcktkffwZQjVeKykUf7YNVUaTp3+O+jVrX0ggNNqoCy1AVD
04ymmlT/ggA+v0ZQME3GWLgpbYgqGZe4RUo66RZiGdKRXIhLlxPG1VWR2pYSm6ve
82Ns6Aar+Ps7EMXKFptn0mvzWEYHV8dmXMzO215UtejtGc5DeIGcdBqAqUQMowxt
I5lBnusbhLB5b2M8xz5/b+AglYaA4wCDmNk0T2vq1MBIb8LmAiLuHQrqu5dBmOWA
/OqEWDeDpZTrLLWLMuZLIsp8SpYb0G+MarFO2VRM5FSkmElgzDl8by5nvOdID5yp
sqvQ0OR88fFX430dR9WuB++WBZgPxfh1h8x1jscoSf4r2dwAhg+rkHJlmm/BjImt
TkXrMSIp2VaFNARo1PA/zu/F2Kc0NwMf43wgBeuSZnfoTjAFE7hNVnbp/n5NrJns
4dLTvCetJcpVDIiI1uusftu/GoJzN1P6nJEakYauckDd4dydu/BTDD/l3BtjQh/W
TyQ2QEQNtEVqwuivJIJTP+HS4HmTdAbDYmYVCY+t/97O9lSZ55sgdJmJOc2X+tYF
TXg1I62+Gox4hTQOGP7sHsNzb1YKWuEX0TYwOW32yTvLMIbc1Ai69EY0PzEs3deo
oMjFHc1QGdeAmezkUdWWMX3x7/w1/mTBBO/Atd16g6zcapiocLs6mu00tJyU5Quw
dURCtXuDI6/hlLmkPGeibMHU/7CTCZ+rFGw0xbnF9sLeqs1MA4w5xZZ7XAIjQJ6W
4iWDpmObwopJySlDaz/XshKYCQYdiqVTXmkmCrb8VQZ01qKs4W1LSsCphYfzyj4i
i+anD2Ag262d7HG71MxNNGmUTo8dzLGL043btoPwEVk4U+Z6r2T+8sOsbmrNJxal
sv6OEc0OTaIXjA2uWEupy380AhA4y9/oOC+svEAZXYVTZpKFIUaKv/5RZZ2XlCyg
no7jwYYb1djHAZQ+LOfr0xCmkKjHPqLswCf/9vtFycrZt9YtdZ9r8yusW748aYS3
YC51ZYi3FWd5yUee1/ZUQ/7t3UpTnSNW08glK0E0dfC8zS3Emh9huS0EKPEvX0tS
qeSKiMOC7lkUaUWb+boVD+VyhOhp23de8xHsm0dwxHc+ngxBccr2KvkICTUq9wy2
W7zXKZF/mtGNSIns76sBDC9JR/VhI3dK4p521XoVR3ER9feQIyciu4mQWeaO1wUY
STWLKXaHKiZBYgFDYkxKyilhLbZjDE3Nt5thjpiLFfOqGReg1XiJfUHGt0/jFWn4
fJP5js8k7MmrN7EUWOiCkc2n5cGyXfoFgKhLgNQzu2D15HX3vW6l8+1b0ze5ovxK
1JDHxLxmoFZ3jNo9Q2D6V4iwM+aPp+UWV1PZjTzjoJmQaAviThusaGJj0hKZ6a6w
7sosW7XDd0e4FgbhrQkl/wS9RGh54zAr4ggpZ8Q/tz2TNB4MQn3nQPPuBIHtxQaO
Ri8ESC4CN775DFsxWOJry9DHm0FDY8NAy5ro2XH+wVJEcjjkxKUm6qiOMc0BRkHX
sJ0dUkadJNJ4hgBm+PNP5/z2rdJhssuiJVnAUNboRWu1cgCs/XrR0lh0l1BA3Z50
52brBDdp6hMMw1rw4FnaSTw2I2+V2znt/oZN75NoGXMazNXzHJD+kDQIkoDiVBvK
wkKXz8hPGJ/nK7mnUjw2QCkbAR9KGpBcIug46LYRiSfvw+BfgHoWtAswdNsfty3C
O6JSSWPhz0KokTS4+Z8eAJptaHmTOnnVfS6Z/IiLfUzQddt6us2ouq6WV7eVy7wr
lCMPND5GSWNum56JD1h2K50K3nhkiNT5bpta7pITczmtXcF570vHJby1RAbqynnt
1/amMy/GfV5h/uDStJfybAETtRu6e6aHt8xgJAxq8Kki6hxP/WqlftrcOU3181EY
o0pFwTEHmzD6CWjjNJWk+8OG+4JnwlmfwweTGJ5ipa3Nvuc9/SRFApMOk4PqJL5x
jLp580Qzs3C2WbES/7s2z2lwXzh1TQxYiwpMlgMtq2gZ+fxvEbryfm8mCEGtO1Ve
38w/27s79vV5gi3yJ2sIoqwcJ3nMOD6NQj+0mHouMhwS6fhK82UCFiaQ8o50PJ0q
XWx0CQ3BrOx/fm7AmTxe0KhGvWoWMfNRKYywyfLTwdHOu3GoiydoDVfjQKmbgtMC
8a2Ke7KMAUZGdXyGVMcStkejL+xy7H42I252oGAQJabBgGLhrqGVOkD4CkDDi+lQ
oBQCgp9L/gUx8qxNzT5jNfj8ZQLW4BILdmqUn8DspVS+KMysjK1lMCOLCQeVkuZV
odJotFL55HlKVXWxkTeV5Ix4TyrF3ktoRETS5Nwc665DtZeJFfiMmftudiTWAwNk
eJduKzGAFg80kmB1XQRCJG+lmDJlGKOV4C6u1DTkE+V2IIUcuy+Xazrh4wJDtSYU
bEFdMoJLMj3Br/fCMMMBiiaEyX/ZgiFwNhfsuoub909GyeGeN9GohKLbgqeMEbSK
WqJJ1IJ5J16Rlweh93e0tS2W8n0NR43m0ISBz6dOgLNH7TovTnOeVP0ST1uzErUK
n5pTdVnHIsvVwdYp2FSZABl+onbU1L9SS2yM5FsjNNWDOMNv06U2gH3W25TPyAY9
rhmGU48L3Fd1sszcCOa86rPQqlNqOyK4OXQC+WxogfCAkWS0e7yQFExu8qKAbbds
z5CCOPS+QYMX4jBB9De3SgP2KG/JvNkK4ByCAYV8NK7+QFnOD3jn1mKxG+7aStcY
vOMJjSN3l6ETJycfFdyPanY4esZ+ne0FlQYtcBK+G4snZg4mgp8AgHEY9tp4TwCe
nWSrj0OpQa20MnFFw3r6PHqyBJzISda6t3XMHXPuw33pITJGpD1zKZctuCpjWmu4
QgmW8ymgrPEsCblr1fUXzMIr9qdh/2Sm/FLJuQT1/d3gfIpWpO2Tk/0gdUrh6iLM
wzKD1oov0iG7OPtrEMCG/FL7u/Ynw5D2tWSJkBmjPln0QBh8X5v5Lo+jFDLVT9QP
jEbkMJnY0LK3rqrZ0mb/Hr7g3sq2cNK93Y4y7WTtU5pR9/6h1Rx0vsJOtvV6hq33
gl7Df0ubvnGK3VCBYGbx0HFVgHcY9Tf6bJ/+soI8jasppZ7sE08K2GecZq7Ss4TV
DFFI6w9NAv49IrVrFpx+b7z0AsDqZ14xAchIryPqiULFlgttKxvs7knV0ZHSOGUk
reDjwroe9TOGjiJ77ZpIHdYu2LyI3jonxqQC53zEMGhkmgkg9WvzcwT2zhDBxr2S
pcOR4+DquqC+y4P8WB+YWRfF5N0iRAl/XagiYibrhmiavkEoUysXPsifxrFjAY5y
aGNJ3B/QhtMGse+KUEOazC1hahFaz04Lm1SEFLU91kD6IDDlIEqQaLKfNUXI/k7n
/RDoUqEUWXmHl74TYc3gzJLijqm28CEdbmiIVHwS3RyighxzZtOIzAy1ujkpf/3a
YyQjQc3VT/I+meK4cRripIRT32lOlT2V7abI7GasUAFCQo3yGDvzuHLPPgOaaiOE
M7q/C95rtA8AKJ9h7U1TnUHcAb+GhG0L82Ic1sgjUS85d8cMr29dYLDzXWP01W3k
xxLEgsJ+1+a7OU5osemSW0Am57IN6/ToIqdv40CV3+ogPOE6L768gPYEH7jUkaHk
MpnktluCT2CGE0mWX0BGKaclHuCVLgEf7v/aIYOVs+sqpH1a6KMZP7Oc6Daiwnqa
50Tc3Yd6++qq2FruT4gxZF4McUUobp7vMp0usxl9J4bMvhtM5mGn03t6o7urYqW9
HuG2MEjSpv8Tale13NyBC3lahZ3suQjsYs8hf9UONhUmaKIbL1xJrGB1Zga4SxW4
7+xWZFDXu+fJS3JAz/Essk08Jf1C8DcxdlpgVdqgG6Vgnt66qHJauAzatyKXdG1j
z6InklL8lstkzLtALXcMgPQjV3+ROT1HMBMb1MqV4I/40nPH6Na4uxdVLHohv62U
rrxa5vJqYYS2k7dhRpiGn/bZmkyzMS640xs8kgpI3Rrl3wVZUAMZNHE+F+Y0/Q8z
/6kiS9dlDF8RE+rlyB1j//NQNIHN0nMxf1WA/+8J0YVBZWitL8LiDRCg5LLw621p
UPCV5HTDwkrpgYA92NE0UtQ6PVrkvNEAs2fsyjzcRQbxv3i8neTtaud1EOZ5v/2d
XOTwd7ZrTa0DAt52v36Ws+TOp1ToSYmVxkagJoY9/ecUb7MtQLUDV2FnOwROrh2P
pYr/onV4Cj6aJ7wPXAgXlmN1XfGXATtBFh8nTpG/2e+Kp5hpfaHsttc4xnerV7c1
/TnVyCi+PRq0Eq3aGYgBR53cv4bR59nYhR/GNG0fvHxq8QPD5TMHZ3c0pj9zp6nT
1Klo9/yawHNWhMyrgzRh19ulIibfj2fe1kMIBjEjd4pG8lnZlimvTXTxXgbzzR4e
EVhwP5WNgt+ZMIZJ8raSF9NTcihweOmpHID+baTjaCs6DCnqkwCS7IAR4KFMK396
D1ADg5aP9AeNjB2HYb+Nl+NPQG9ZxqhbtnrvMKVAGU3lPai+aI+6bmtrgfqgdGqt
SKMDIz32rTautr5nhMfdpjcf9K+k76ZpTl08g722HhQ2On8W51HKE5KEh7R1TNCY
yps1tkN97TXO5bvezBW51kEvYAhnqMsD3YiE6LpuNr8ocRTju3G9JTCQOkJymGRU
b5BdxbhI7QO8KF+JVGol8SyhcfVxZ/VLVETa+mbuo0FGWPQ7uHWEfOi05pvWoeHW
jdw6Zw/ot2Naf9pqFPlQmZCf/uQ7HHk+2IVyguaBv1dRcwRDzQgaHowhK/AsOwOj
phqnPxZIqwtmRJxsT6OJ35sOr8ChIUrZ35iIp7DvImM7dlHOOXTfRWOFZkWZMImL
PMPWiAZKasX1pOjOlrBtTqB8iLOIEz2cMdJ8MaugNq51k8lkaWgdV6EfEZco+lPJ
epj2y2jrhuKyynSzGnN3SGbMr4eYd5Q08Yzf90UggkAsaH/657O1pxpBNlAe3yDF
nl2g9uoaMaKx+6JifD67s501gj1p5OHMQh0o6A/WoxhBcL7Gt2pUPWxSvMu/gVv5
O3uKt9mvl0LgaCytTl3PC829PqqHJHbzWJgd2d31WXcmc/i4JES4KThsMkL1mDB/
Ugzn2fP3qhAuyP/Umfa3+uneRoMUAxBsxu3QMwXcJyAZHrgK6hV0paVx2g3vwdWS
l/O3foiFZ0tKx2eWsfPcE1DiRY+ImahEuE4xrhkwUV8F0YAi/booWF3vXz/0p27Y
FANjlBG7g/KO99depQkHvfPj6qkc5ownFoviyVYVXCZoSbLeK061caRXdxgVlNdP
TuJhnEWsqEz1y5nv/kTQyCrvYvPfxipLgPzWJ88Q/L39qO0sUN5QiCTboe84TAaU
UIIOTdkL9Jw5LftBttBb0z46uBFZqJTsF73gWj0NVPGspJHcKhhUqRqvteSMYjnw
n9QX04xaryIf9iOC+xgBJW/83cNntWxe8nShfE+yqc2ISE6OOgBc12EO5mVXn8FC
C4LVsvqvnAIMMpleC+MW+qQMg25bVlLmj9hz1FG33myqQbLz3UU6HlJZvX2wFZIJ
ScduYx9LbLkManEmMslpXUc/2FbILh/rrYqSz5Y7ccIsGtJcKonGXbasRXCrRmQ2
Uj6VnipH3r63W+8B1Pr1eh49226W+X5kr0cm+ahfYK5SSzKzllygOuAfhZXnMO7E
QwrfgLdEMHS0PL4tDgfu90+/ab9RC2KtfLQdtYOfJsgOJIHVY8MwhWXvBGRTWpNd
Dbf6+3meSFI1+7hI0J4M9DgyI8WQPPAhWTyWINe5luKDSJChTA7EoJtLV892osGs
3yHZFilDKEtILnoOc1rkpPNUa04ssKsPe25UueE2+fmOnUR0/UWONzF+fIQ7N7s/
gaePO4ROwAHSr9KtOaKAzvw/+L6hG8SU/bmqMAqGEtwUPJDt45KU7Kd+kriTagNc
FHX+bYoFTZgzayEPE5IsTYi/ySlO48FIjV4DenJ3q6SLNnFmKRAKQQxkABofE8Q2
YC0R0omUlZ2/s2fDtuS5Ch0hUHhVG25kNRlhRQlbjpyKshF7AFqRW/YuXwbI6BWj
ot2JEUUIQZLjwcDFO03RAHACb/rfGSybLLpQAFakuV3VHrKolKRG1vYy8ksZy2+u
cRYd6seQth86tGdJxs8kN+tcHDvBgh41rxpdNSxwwjYAwo4qm0YZsJTVGW0RTJos
P/GxFWpk7dzgvSz/oZ012+KWg3+RhQ6zNNWUhV97hBN0hFRvlEI4Uni3dTSrHrxB
tJuU5bO1axbs/rqyzAqUcAVd4PmynH6qlUVOqSK8MHLCQPBtSP1zOifWOXDkQ9WI
gbW2zTq352QtTURPaalkJ91+HEIeDEXnbayrV86Zs6bPyDZDOmwKYXmwkC0YUpTG
APbSvMwGjRWvVoOchV12fV5RaWihKbPG3ib5YOHnnmf+TxXJZR1V8THHPTXR2+1U
im//nq2+WC4e6uK+6XVn90ND1Dp/QxrPppqdkgPBI5JB9sCPRfAHPF5OrGpcQZ35
U4o3MYDZv/Qi/M/F8mF+hOLI1MJJy+sdieD2u6MpkxdN6051aT0Ouz9J+0b7RSdf
mvIqKJwyo94cu93CgbXsZT9ChwI52Sz/dC8N6KHaCBShisCYuXeZef8POsiukvga
Ffp5RjEtomgvIgR3lhMpR6ovCim4Sb/Y//l6KEWa6sScpcd0VzKBV9Wz2lecuuJ8
szUTRZu5IvyFYY5IGZVT9s8kw0SvChDll1YDBBV4fbNiGN+AGZxptQlqmg8Q/s9R
aMcnA9Asg2kvyX8cy/65NQEbkUIHutxQtx7KQJNaEX+D5ct8iGCw6nic8zTwFa5I
Yrq9iNlCTYeaJ8e4AwY1+FOQXS6zzpHwFA95iDavLijG/Jw2HDxYQcacVi4MOpFQ
9H9NLPdYrxfIqrcIgwCpf/vfiI9FrrLOKwQFIs0pDs3IeAmXYPR7BY/DA+vf0eQP
oA4JQNP3MkPKPmTfn2BFtITAqwgJLwCVpB+ARAywyquaxZT7O5YdCBo6iwAiS0y+
Lk66udgMPxlIW/vz2ajnmTqeIZw7TG0uuwz/8N4shiLhCfDHMmbRkoiKxkbp6TGh
Z1kuErGeE9HSOJIjPdoFr/paMK1JCykh8mPls07PA76MaYAkAK/3uAKEYraupeCI
dc5ciH20J157+TQoX8u1gXJXgRsMWhA55T3VTsuGUiUYv9D5PKtIo/JIS5Vj1Qrf
2RmoL0KxSKKvdEPHpqyMMo5/xiqimXfQRdngB5tHdvzARovmCujvdt4fhDOZSukx
fLOxIf6m5mm27QDb0G/h22QzOGWcvidjazEbdpQYwrlDv8NNtJsy8vOXZrDBly3X
g3P/aNktZv99fZ1wEKYFPklqUOVZgResyasasuUg3Ru7jJm54jQAYCoR1LMkvVUd
54RlPMfYmg3rJVZw3/L1UeL/aWUOtkzl9et0l9KAS72RVzDifVg2pAnvYXVGR5A7
sqLHk8E8HMITgzIUfZgMYybsiadaSc079+N8iwE2+KJamzSHLJVWaVkm2qVmAMrt
qcO1zyFBC5h9Cghwwc97llLN5K9S+BGka7BgYlF8C30WVMgCw41L12PYhy9AMvCN
gAoFdo2WYDMyO+m1XeH7585H4bhNCG6tbVZn3dGM1mxbw2erhnYQO4LBTgFCuyOf
CZ4bh/Aqgnu3ffqr1FHGdo0E4pWaKUGYioMrMuRDNAH6rWHmpxUMo8Rt5xEHFE7Z
9+x0S8F2jLpZJ/o8AkAspRsIHQ/6fcH7dz6k4AqLYS/V/0ocpUtwNtqv1Y+v+Mbo
nd32fxmF3qpXsP8XPuCru9SejEVP2DHBzXqzCt3nlJCU3ZoMz/1e4xH+5DJQ9at4
bXoxFKPzMxuentyjMhnj2bUTdWTPHI98P7HffVn/MNgnyPUQ5xkHfwAfu3WhCjKk
DHLidYmPdYtI2xRQeeLsPAhaTFVIMJdaMGxf8qRGLiE/ium4Ztg4ytOoeTrpOR32
Vv144PORbPHlT/KssUVEPsyhMj+MHaWRlcZ2d9u4l+sypW5PPBZ5bBB7KipFIsaP
oYxdgxasypC6P4S1kWVu+heP3NeIYmNEli5OIMr/ldpFPXucktMXuuOBBlKiJybv
caYZk/8fYXWqAQ47zfAamH3knoYK/fQ18QuxqHYusJqlf4+26/QV0kMt/phxQaQW
V+AyiCstsDbWGHJkwjYjUFQU0zltEiRgb5nNcobViKl0bOw5L+EsliRUfOKGCY6x
2GrU6ix9DJZ9P1NxDjppMdiHAkHkeNU+F+pk3iJE5WaM5+xordb1dP2uiGhxT0wi
AtltC3zYIkAjCFMb79hj7Y3iOo1/lLOXRF+gXAjIPt4U4muCu3Fm2ttQfczRGlRe
qBY1MJmB8FWbV7vOBOdJMwPuNDReWfXdaxCq9h7zTLrraEWW5pExv3fiwifUEXD2
qXGD/e76JxWRCNRqAFPpDQKe0RuAj7TSrvdh74PGQPX29MpfoF92bvUe5V/ptdQZ
Ml5nbXhWu/TDEJ3AQrRU/L0LK4xApxyrmJce1bjq5D5nSb2TgrLzkHhjXolmnCTW
N3pEfjjj04RHH6FblL5k+KDloxe5HVhR9u51Z1nFfvEn9pvHwrfWcxqlTHZAJvaI
3WQxBL09W4HICT8qulr6ZnvvpuC1XchOwogvSi9pRCecuLgMgzyUnrCm/9yq9kzw
AWQY5UMRusK0WnGZU+6s3izn8ye47/pUSsPvSLRxJZMGxbhWMKatmUV3ZzDehTL5
M2kdeFYW6esOkEFifKKtnbWHIwD2Sabmu4RiFqP8WUoHh47CkXCTknezwCC12sET
jzxcfi5kJkdCYPRYqhKkRt8usOwwuGpHw42EE9F4/aBrX6tye9mfPt2tQsYfC/Ze
CtdC/N7X8dlJu//j6hVnB1EVlmxq+1s77W7OQ7h7nG9HqBBFSYF6ExkjoYQMejpy
rD6zl589qS8prWoUmZzXWizdqcLF8FMKbfQOq2DMnasrPX7S2PZFZFBc4sD/NuxX
umOYMR9Sj+VGIU5zjfy0IlJUQZu2wGzL+lQsV2xeUnkWgvqoTTxcZuS1gkOcLtQA
vN+uD5AGyau0IPIC01kXrTuMovVCIgXTcvQ/SbWzT6jhl6HePXje2feR3rUaan8C
1g4FBIGYVzEHwQobTpFr2i9plLnS7id3jZHAmrFA7BhflhbcVR7Q/pg+XFLSuG/W
HRsWI5fwCjTUQiBrrm8/Se+lrFB5tntRQJyPNL8QSajPUNP80M3OXp1cSVSv6+E/
uSekpGdhf3ZR9naQGBK05DX9enNubJ9bUeVX7wFLR1qhPofUXJC1YcaJQGw8srw8
rQrZ5SX3EHnTD5MZYvVHZlUA8gtWuNLj5krxgU03vAUg8/pfeKH7LDDkQqP+sPVl
ZUZkWtOx9cOI/kIFNtxwzwme+DJNt0RbEkowRNwPgXzIQ77PWT3Y/SG03coEx9jx
buRPPqgPLqMJQu5jTzNgeX1u1OEuh7MxBEgmwTRWSvqjTFzQ2S28cEH6tscCnbT2
wOYYqzVd5SXYNICPa6+RTyGcc54wP1TfcgC0AsV6j+0WoaRrLRK9zY3bRP1XMeSz
OfD60o38jdmcvzddzsBnLGL5ezeduDJu7UNRzynRWU5TWnyzjre3S34WI5IHMYV+
CHkibyViClUoaXmdFgO38eI3a6MCoZaBE9NPTNNb6DN+MyY4y8VHzDHA1/pg7ojq
v6Or9k978tYqAgbS8fR9mO0/hu6wtK6+c/6x4lBoUc5RDYbMoWokeb4Lzu3jCSSj
MDTNq9Yk0ypitlQ4Jh96G9zR+vKNPRJ2u/2QVWwClGo8KRqAsyHbUAPzxn7xsNjc
cqzs92PqVlAK/P8KpwLilVPE+es7VK0tsoMt62U314kRAc0zSTN2lG4QAvifK33u
e3lHqUwYo/QCSKuSVZA2IIeRZ5xUAzJyYAboujv1ApRzmY0WohlIDFAZObHOnUC/
4nU+B9RFddRbEyG37Fpc3Qwb4G8kAyEPpZtGUBy5qmX82D9jnUlhXGA6pLSJDA/0
QSjFqA7bRadiRG8LsgpkBOFtMDOLA4TyEsoGhbI7pqHkH7cXke6lv3xNwnx36zoj
NFvb1VNBdoulK7D04YIRlO1cb/ooeGTzRfDK+wWZ9xxVU5j6w02imdZI02ZHQ5DA
fEp1Zrch7JlbkVpN3W0zpI0z7Hv88Zr6NBqtr2aKKrZD7difZpTei+sg15GpumJk
1KPDAF/Nupeq0v4UvI5i3ngyK56ly4+/IIILUUxo//PEDUGTpYJ5Uikki2FJRU4O
nJFwnruU+jc8vZ1sUbl2BXqBA0mJLBKBwN9EBQYobCU9nDei6FSO12SShc+AMfqj
9BW+DgmB04ncY6s/jS31YSwmzApNGwHVX1azlYrLxxie8RtyIMdC7qoFkOmLnwmQ
ZWB9LOrHrY6FLcFSpYAw35ecX06DHgf4ikfWuNUJKgWShUeclPrPC6xKxeNOQKtw
qBbfAVleDcKnSi9s7S+9sLviFPlpgDxcjKPRBDIqBHTjBpym3Rn9N8Gwdu3LQWoO
bBcE0geiomA6c5oK7qZU64mKEBe0OrEOqO+dkzxaaMI3co7Zi2gAR/jyWappyZ6h
/9r1dcVWIIxMTlYUyr6NBmouZUXaECfnvzzwkVnW4jJ9lqxicN6iiG9VevGWMeCY
ybnQpNhqfHCOB56l3iMuCWuP91upkm+qh1F5p4zRxRodJ7Q7DGIWwTzDMolYvBjm
I8Kj4jCvffM/OQxQI6gmQHA/goQAfOmYNk7fftFR6Xe2eA+IfbVqlvkkPIZz2zc8
YIB00WXUeMwZjoDiiytFwM0/354s8fUOGhBtS/0CvVXqd8E12dZHH0XjUID7pH/2
ayY869cVtIlZzqzj9eHzl6rzSDGRM5yeS4fwA8f/FBjhKh7MdRRpv+oslXvdTOLd
XsV+xx74YUmEHoeelVPriSjGG6htnSYQRy4UD7nmgfjhTJyP6QyACOO6f9pW2vDs
nzNpdfh80SbYGfWQ9NcZvwqCpsW9KkGJdvaJLqLJlPCo/pm0zdbmUyYPchsMDfOn
pCk2TRXYtKBGZ13czjaqTPa5+pgY8ohJ/nAXq5XrkONJeHol8+LSfzZ+jQ452kr7
Kk2AwSzGeHzXhJAIr8ZQOD7aqHLJe1AnQaFW9/QgnRXGzmp6X841zgVJ0rbbyQz8
YgGmOdpvRZf2oUYqRemrMMXekRXnuj0PBjhLQVmjkML1LLRRNQjomPOEICmvYbEc
KLfzS0mqjkd0tvtj2Ec83BGYcD64c0MPei4gZ5GVFVURIbzVtr46MLzZ6QJ8JLeU
0O/jpj+oCHAzMqRjLH56o5L9Mq/JIDTB0jIbZ6UjZ6zi19iLcnBfC/hsF7lLdvU7
gAKtubsmlUA+gL853wLGb98Kk1WRUTizFQce2tJJ36HGZ8fz9+RgKmw9/Ym4NDak
YiJ79QpWavmvxI54U3NeElGgC6yuyEk643QQ4CNkOnVbxALD85lGsdBkcKlp5MAD
yd6baUUPH8zk5+3YUp2JqExkB1XoF16KfyrSA9fkmvR/0Sbu8fjdJC8fI7gRYENn
r6Tm5bgFvJ7MuriP7NmL6zWvslKWYFfw3C0jiQv5gIGnNxQg6ZGzN/O/jbL1B8/r
Hx7SwrFeyhjOuBzRuG5+YOtmlWA+JK39/V9WjDnGUGnxae/WXnk7tPU9ifskGjqp
9/cfWmldA+ofSYA4az9Ldn0M5/VRgsTAAG8764HtPm6BJX4eEU4cIh7yUzvb4huu
luHyXg4WUId7qb2MEk/SHf7fipp+XHP/eRhv6bG3Zm/shyLe7AH4bdrKfGol7W/0
MP0yOFvvcl6cq6vaq2yMJsuKXYMNP4Dm6jApglP1phvcEqfWPoQhA2Wj2kIrY1Ex
UIL/lDgfsrt/INLqfJsYSqBT+ET6arbi0jkzWm3wE5XY9J+dJbP57enCvgjh/lvC
pyCtpUwjqKxh6xmY3rnN/H9jdevCZFXN7lU0pFtqIfI7BcXmOTWCYFhqA0m00QJi
p4+n4FoYZ/pVPGMS5yOslJBkjp2bvwDgsOWytiPAboshcOPbBNRD/mSGfXAbohRk
YYttTBHBqALcvTB4b9kNiieSfqzGZZQgNujUeyera5Pfl3KnQDmPljC5C6jx4tgV
9DMsPExUGBSmngMgogO8EkCrUwluDZhLXspIeldhnm0Qf2J5bQxhqsGSpRLQiq86
awbCk7CESQGz+bumqnFHTD+lo1qS5IaeTw2wJpD7H3500UG3yanVIpIhfKfsZI3j
4rEdwbav8CZoW3Y0v1/58vTRuasJaJZyAhsrmABB3wS3Sy+2WdkYOhS9+dck9Gp7
kPbBgd9i6/CEyCbCv9N0bDQ722q+YjrIh13rAXAL59Yc1UrZqJxruOBMoYCiRzTo
KI7VGvksl4EGDXGSkxqNMOaxiCKiAspPncP9FnqQ/mXHFHn20DsBmotF9mWw67gH
iWk+TGCqI/VrYVtAKiXCl7Wni55G6c8yrgv8wvZrxkou9QpoGzCzv+XZki8rTNcK
LgiXSzr7Dgh+baBQkIgbmxNzwN0F6Ta99q+yCcE2ziKX+kgPVxbVjJQDincQnf3I
0e2BRoAdttm/O8PQzj/g5jC6Spj4CbuuMEh6Blw6lrOU5vnY2sMRRtqaL7SRo4Do
NIVJ83mad21el2wXlQKGseJxOyq2YUkXac28y1PivPyilXbr33qTXmwTG1l61hhS
wyBR1gukVDwXN9jCZ6SiN2sMEzTjm/G5vrul0F88O4sERBe3FoCz+e4SeLz95Eu1
VVfoRscdC4xmK7ii5o6FaY1K5YJcssHPQ8CZb8Q+pQZNvm9//QQzgvL5Hc8uqqju
DtuFd98ntidKn9a51E4T9Tq4Qp3GGuJckXZOuJ9el2ndAXiLIZclllPtbX067+4L
Hjsoa7SMfZE8Lorj7hmnVylWv7G1syoziKajkLbZnnhB3mvY4ehFTla0IRf6uuAn
KcaEj/m+qJM9KgsHqy+rSFIBsvYScEffjzQSkZn2pIuQR1MNqgDKbd6FFhI6yCZV
sTbNrjuW4LlAz2NRrzaXsJmtb4nqPQEgqVKiSVUWuWEci0O7g8W2Kfeqnw65ctsV
zYS8oc2Hl5VHDQVQ8GDgAG+2VnFlvAziC33JF3rwjlC+OlNnJBdP6B7J0MChYDiV
8Yqdze0Ms3jeI6JwX7J+VqVdRu3QIURlUOAHYKEu74FSQcQrbyTR66ZsZnztIjFs
CQ6IWj2RLTVst7fELmoExNvKGAnt4s3D8drV60zzHef7mjNli6zLdmNd273gkiIp
m5Defk/OMc2bTWZqz3bJekr7Jv0xw8dhMeAmpHJKcqzni9G1u6j+QWedi+XQMfso
Oo0ykrCQRlwZ5b2v2KoqyVhmmF9TBs3x8gjct3hjXtsRLmf4en8BalIQmwGxtz+/
U920UW/bs+YiEndxM6nBuWf0B1ufPMCp38Qgg/1vmXDff5hshs9ADng8YqeM3P6f
t5K28IfpGajdheNrYKPV7oaJtYWH5spf/QhwkzTabC69P2jSGvH0qqsw3GWy1c46
eDCAMUcxguCu2r2zZEtl44W5bO15kY3sNKytsiO5uPaXwcbN9D3fPQ1F0hd83gDh
x2il9CMpnAfqEIpDFOc/bevC/O/0X3RC0T8tBSM0nweOq5p1XVgrMci5/0Y7/iam
VJN+qeTECU5D2Tg6q9M5h0BOipP0rAdhTzXBAQwvOk/JUXiQwwQIgOvWJ6FE698O
FtJ2VAEwE0q4F3WR/WcnqPvfwl7KjA+AiMIRcR2u/wGhbCVQh+zJexwq2IWwe9qE
XaiCpLWP3OR3yZdtb+2BUJmdQoJRgA+l4vTWT9xyYj7BFfY6sA+KF1sxxC60uzWN
sjMTI67Ty8NmZBY726su1WBjdVaLjm8hSpDs9euOSFFEUZX3idck3v56OrZ9ICRA
y4dKKrqJkDlVqABu/yzuUiL58eO4Z9Lmk7Tk+n59iopHAMFgcy3xBBq530jhZHaV
6voc+DYqwqL1Xt9Ms9xFF/9GaKX448OJpcLISp9WgdcX6u1Bh/h3UesUR9wQCO1I
KwB+JwRS8H81nO/OHeiABc//KWMLOMbnLyELVGMMxdkndp+XUU70DdKr1rDiCU2Z
8Qdenn5ZaaD+JXemQAaSwNJmTVsprpXnKUsCYpxX5RWD065E9AVfrUWlsv1USSvx
D/n0DTRGrjYX3hDKO7U1/KcR4hjIVKc4eakwsa8zH+rweLOKKFh/DT9uWnMyBuim
l+xA+CE0YFJD1ZRaPdtZsuoiGNy5p5hpXTUs3VVM/5lE6FboQ0NqzDbyjanlxBCw
xuwRcRGvnfrbIbQU1S9LbJJIAioV8lrjVniddzKBNojuC8zuJlNGQ/ZkAm12utQG
23Dtohy/Ik3uUjR1077xI2n6hMrKiyGTj4b7yrPiQESBQjuBaAGNFHOjHjvZiuW0
OjLiVdc8Mvwm8vP1VpolFujrfssQIVVXapGfoxxRfgW9JABYbYmRC1IeleI+O95x
7qvWwtEa+5Ny+MALINCczoGrrNPG4o6VCYw8Xk0SZJU0aKBY0LquSEe4SD63K338
G8dCf8zE0m8n5bFsiXa6BnZIFm7qS24U/dGAW8g7iSBoJvJXNDRZup+IqyxJ3Xcw
+ssBgD2Y7az+3Fgh+cnhm/0QS53KXp+9VrdUkuxm8CZFFui7nRBRy8pHItx4Mcam
L/e35PbJBiD6IKRKamjuSJcujzklArjY0XRx9AxaEAPIx6UjHj4cZ7K4rTgD3XT/
wh7Nh7HP8XiyxX6Or6Eh6KtThnFBc+nq8XQhhECHXQ0/x4VL63e8VVgTirO5mBv4
fGeKaJyOzaZHekQy2boId7olPREw6tKd6kBSTn0DG6JpgGMZVLqS64rNZyJeeIto
79pknkAAG+4UnEpgVfdC2ioC4YP5MOOcYZbwi+HcBDN0gnJeUdefTHkVelApHYjp
tx7tlpTHU2FxzqjL7PUtkl24xpIlm7F9/JTIRE8sI4R6Hmoam3vHgJVAxcSUhk6B
z2UBZebxdgqtU9k+ot+B1cE/wUXXxR/XJNFSHbqE921uUvZNTJ1/TZcI/jyX1vYY
WTIz74cKrtldRvi4/oGrzY+l7DwX5S3h7pSQXpsuYA6YhERfjWhkzVAmGaD0lV6V
fKLhnu5y+HXjWUN1cLKkIUPyOvR1Pb0tJ2CCIk0ZYlBbllApAc19ceYlDg+KA0PI
hNWW94N6gpMbOrS2mLIWbF0Dp50w60EG9PVVH41K2caEOC5461p4iVxQzXLwniFo
O2/JiZnmbBQ8a8BC8VBH5y8zDunz86Jg6Q2dJrWJV/CnUB0Kw+JYzZjAeRL2PE9l
L4OGqvyqL5viJZNI4X8rP1KYdCN9iLQuNQpOAPsHoHt8E8mhUxYMiepw00opCf+a
bQ77PGF4NmDwS9BmrJQ0W7KIQWO4DIY7PYGfDO62D1DCCqvzVTMeB9a6K1yVkSKp
lcJkFb+ZE7ZCGzGG7qfn79OlCAq97+YSgfB5+kOSyN+5En9BS04zO93WygLyJxJN
ZVvtIAUkoHjpvgW69zu+Pu53wFOLFDK0uV/mJXWS5EAxobUFllD8L3IqEMoXgedM
2G6BwjKx2rz/7IK4DqEwH+9dtt0ziAQLcz9IuzBXOJ3dbnsv5c5QSvVnWf593T/q
+cJvM0D4gc4zqCJMtqkhdCqfXnkjItUr+5CB4LOQk3FvrjpRcn/4j+bRKtLEpPXo
JdcJHP71zxAbJY6gNhqpq7Pr4jYUkKb7C+fqYdkTvZF5MaqhRq980I3nGoP2SAiy
KCh5VNPYtDfxS1oGZ/dn8mikNLmDG3A9tpxZKAs23yzr1S0VzDEiLQ3Lfm4vuK5j
1peOQYveUqatz5Jrl88Y1pdGH7PIv5zzln32bjfIeQbCs9H1XlgxL0FU12sEKu9J
W+NrFzMvQf84lLZDtp4zrE1Iil90OX/C77ND/CZn7AlTIUVG8a8VJTFC8sZHmx2g
Nkhen7c5ILvNuu8Zgu8KoDBtKRsVCPaOWgzV7+VAK4GwOcxWXhyT9ROP4i65J7Ka
cphmWt0gNkY57fsHrYx/pNG/8ERlGPyZ5y4+x07Zv6UibTJPluXgXABf+TE2TCY5
YeLOWfKF5CQUXvCtPdaemhwYdxkMvi6TPejPYjcjGzV8El5o2IWcotyD46FHMj5e
BuhWOGFaHVeEVUxj7AQwEK64JSc8c5bVNx9hXGppWqk5d7OzftLOCIZvyttDhTr0
QwicR4F/clpgvzAk/jTLYtePV/x8DFDDXhJpaMTwSSa4aM1ESx3TwO5TRBM7h0So
wZmdgZEH+LxfHH/Ok0LdwhLgX6hwLwcWSfPgazTVLEttxzTHXFLrS0X/KKWODA0D
VU8TPYpdvVAe1gA5Zm9h8C1fgtGKMsCI3uyfqj/YS+PVxTRQucsDi08kwF53Q8mT
/FZWqB69lLgUJL138cATH+1d9g+B4+ynJERXnr2taUuGq9ywv7C9NSSgLM0l6Ewj
zsS7plWIGq0y4eP1Uee1iLVPKN421Ij6OK9xahKp2z1s6WYHnznoB04Es70x2O/z
zZ3npIMqaTpKLiBaqZ7KlY4e9RYIRyVwBzKcMbkAw4PxEwgdY3sFnJb0J16T50mv
4VGgr5TqLv8pK8jDMRLz7HSlbcKefxQSJnwFLL2b+GUrV5+NJrGA4dHGiR5XaUkd
1OM3OxEKdA9YYPbQV8Pa8RAhzpaOS2Upy19z2gzC5dAYv7uFTQuVsC77tIQMpkLm
MR03UavhTnvZedp/V2zY8wjuaEY13qxqUOFRsYZDKhMaLDDG6tkyocX/vrpPo/sZ
E55Po0S/fp++cf8Bec2e6LMZF3dhIU+PRmsAjHNNqCZb1fCQut8WstRRkdre2W/T
APc8H40BXDLOkVUP4MQxA2JzvcKp5GOEihKya+O6UW0LiDSoOqMuUfSYuda1+RO0
HXfVOWKCYlSJa1IBVv0iqoi3PU9xckP9vrSVw45EYXPZ7FOapM1i7MeaaqLvtj6D
8y88mWkQv4VC4ua4Zy0rXMsdSLIGHm/3J+0zPTXWqAsGlyF54vIldaJryvBnHkNT
pPY8mvnq1jTRCPhfeB9pG3ifrWOwMLtzLJY1ACVjK47Njp5s2PQoI2yzhAAkfi+n
HlPCMA/BjhIncFdlDUNJvTpNIX/tCMU1YgTuHqoeA2jmzOoW5N1J2AQwoNhFRw7l
MXNOsPkxivfwKp78xfZbcq+o961LpENSfs9I3FJjmYjoPm9UsmjiriuhGCB/W1Tr
RKeUDXg6gP1kbJvNHhTiXnkVw70mbHdfXbWVbpiB/1IcgH9cpvEp2D+21N39SbCh
ZAGJhyD9sYda0E1t68uU6trT3x6iKoZ0VWIzOt1mwO+lwY9Ye38uMb9mWx4oHqZU
xx3q4K2r6rhIAdWl9id5RWBQoMJSD+1nTU0c82AQw7qvWlnYVMVphbV3SPnqQwAt
6S1xa/WeVkc42E1Trf3kZyTjTu8ogmnEOVxMpsCV6DfvWaO4i2KVldjTWlb5Vfp3
uYdYAuhszCu+taFVx2trkG0+r+Ri7LZnLjj2oABRpKfNNoPQeaWn4Oc+MWutt971
J1gRdgWsSz2r/Ht2lu9xaWni5DwksjsiAzFSFee+ziA522Puht7QFZR1MmPpYR8K
o+42VhRUxaxhp7h4PaGlscYPV1w6FCHYTTK7fBEImXfishBYcVF+0p6fb/pwz0FN
UI3OKorMM31AMOEsOAe4Bj8GfuIhRfiY2seR30+D8l3r7GnurP+lL87xtuNGrjOJ
BODY0EA6nBYDP9KYjJ0RNwgvcZTtglSMgF6X4IxPB+rI7OV7lhZtjzjSKrvESMZo
CkmmBAojtjVHX/wykvzjK5/6iQMH4N8yE2bZKbqdJSWQB1W9l60RpytHvyLZoElf
0WwCl0nRr2NTMgM+eOb3h22rAwnDZY7Trx+CNyaBGlbq/QRf9utJ7c9BysfWZJoe
v7JD+03/D89ER+aXV+MEo7xdd4j8Fvb8hUYKXkn1nRjOETgFX1trCBvh93M9NwCb
kXaYFoTHmqflFmnX/UyRqtBD0Zjr4Hs3PybPb8BJ5xX7/crVWgRexuz7m5F5a3uG
wW1W1Z/RKcez8SKClwfAiIJ6uIfpP0IrhfA+sGDusRMXUi68kZ2HR97NmptYAHjJ
13y3SArAxJUrG4at8720HuSoZUoLNkiaFlLU0/cu+JHqBUeanBHeUe6U5CPIPsEv
R1a3Ic1MzldOGpn/9uioYPGWuaZ+PQ3Ceq6Zxr6wYVwf06SkeCUuRSSiS9EngoKR
BUCqMpCRJymbdZQIfxt86RmuyLBMGBGc6NHlLdfBVT+4Canhru3MHntIzpZNYEG3
+iY3vQfP3wuLdNiSoI0fBWiA5A9+NpH8fAbNmXSt2ef9OqfwKOyK56eYkKYZmTsj
b3I+hasQUKWB/wfC247HajxcmoMd4rGqTGYU7labAFjmIFJSZ6sCRiyN2eqlb7NL
3t8IQUlx6mkBG9WP7fvma45R2rrLVkWelYpMnzUbawumeU0XbMZkBKgaF4lRx83q
Ze4Uo6s3gLb8XIDc2UWMGtTtF22DYzI2fn2NI+DDmXj/pbAkD2WCtm6V0Qv+TCxa
ncqThxMH05HXysokAGmzf20Ns6wzNtOngoK5cqez1FLr0y0FGb2wsHorsw27V+Dv
2tGo9ixFcJRzXVho7KRMm4RIQLZOXSdo+UljNmP46lU690O0eoL7enKsjCvGk+er
HYnwOcbzYcu/2TpT/oczhtgsH9TF5/TUGFV78cRhdKq+LLNyg9yJ8HCEIRojkgO9
x/8ajd0vandKbhjWq/tZ/G+moiEgNw5dm7IMuIuaZipgxUtkTZfJ0wDwD6ezVbwj
Mdo9ztfiPj3jvo5giigblD9rljxi/EFKPnfGVysG7dWGFKe2SO6OOC21hy9FOMra
XeW1q0aSlINOhCaP8CK+qbnstaCXNMIHjVqJ2kxRzuZkdN3gbjHeHtEJfkZHg44F
jkB/f6lTfrBMbM1qVnxyr/YVprd4C2h/L8Wma5cjMGWbw/YG2egelYifd6x+QOVg
ZW/p3Rpdu6Ok24phJQKZUPJ/wJLpUIv/Fp4QMWOKBXapEknKKcrZWx8gxyGQq6qp
JsCAI5Gg7gOG1UrgHoZ20ymWsRZEhAOv3W+TwLZDtUS+8mVhlZ/80C1B/yybRXyW
MKzWuIjDVDdYof4idFX9Y/goQ2w1vvkNToYYdaKIsr6efNSRHvKI9qHgtIzhuRDu
NCwH6MX8LokZuzgPY0HN4UYVEkc1OscTIC1aiVYdNV/2LW3JOHAcvnTzu32WsLIK
aLcgj5eFq6HOUhz8fq6BpKE/u3DcuoUsVi43WaJjrknHSShPtUwypEewlhvnhfiH
+axAtfKuaVFAPTyULKnPQo0Kas5Ax3Ux5noPmhDfeltIKW8OTZrqEjb3YDrn2w2j
Aj0mL9Sp6cPf3s7dkvc/poNZ+TxNDhna4odEDFVjINmNX5K9ijHi+CV0qDp7NYWY
LPGSmGJWYf3l6hY0Q3eI60l2gX23fPB/ia8YEd5mxd/6hTnlJXXX76SR3+P00OC5
MtxDbqd7V72CkuZr6/wKTPUYKFxjsK8FkjH8hz29PsJyovL1cBIjtq573sVy9X/a
9N8Rx4pY+KHUM9QnjLE6IMt0jtwCTKI/QJxUbMrQ24V0KUjz9yvVfdTnKKn+lCXU
oEvsAEW2fSksOf4Fy7ThV0rnoQkBrok1B5sssVRSkfBKZMJlSiRyIVzYMhj45BPr
gSO477g0oTHtKLbOqvKTdP2ZRRy8EH0Uy5VyRROpmpGUKwIOR5D1LhxTKvbKjw5Q
vyiLx4322UeCaaZ0J/1NX1ax7gtOwmfJ0fiQxcFSueuweCXD0EQy84t6eoBkbAME
1LvcRTrSL54dtv+NLDWskXpR95V7gbhoKucuXFxgBvpMzoAup2K46bPhqyqoUOym
IdClO9zH8/rqIlzSNFXV3wzIpkXWaiCkDznAsNdbalhDSk0gI41TKY5PNkCfmj/W
+5OPNlS1ebQ7WdBdAFZ4gGtkbVXUP5W0Vx4o0UXWzL1KnfQM1NZGier1+0kKH33A
KVHqd3o4+aDJj00QE+/vROe3BDBpFvIUoLbadD4KXfh/uT/JIPl9VLcK3K3/qQwL
nge/sO7L6YMomhmAdI+BrDczV8/uDYoJqRTWXku1EqJsvY1ADiLRa0eJ66NqOoV6
lbCRe1eY+CAvHUnu+yvquT8eV9XsQux1+Mz7IoHAg0mDr564VF8bKUD/EZ+c62Ko
R/nrGUW2JJMKm60LxGTf7W2aodPsEySSlFt41wqrNd7+0lCPmmVx6MedMJCeWVim
KLrosK9tsMneOYUfLoqgIGsrA/zjdDsAn/XO7+NFjRSTQoYI42y9v6M2W3vR8KHm
JzF3JIFA4bjTAL0ezDwr7uCzMUYJnHyDTLEw0lejEZ5bXYHNYeGjqXxO9o6pnHiO
kEa4wE//jGl9wtdjw7xtfmjCF45Ku+N/9p53EEQfIohQjL1ynp1xxHzYcEEYv8oD
YMQijDM1slxhgwkGRf2li9ivxmt95FSoPQhFExKCWfkAoX1wt7FEcAdKM2cgf4rM
ZyC+WAjtHowKlDRSBELvDXR7c8KEDEk5D6zddc5DHGoM+dn84kcQ/+sgY7Rcl0z0
YhHAMY1J+PtU+qvn2PbSOFLM8yvIHFSL5gUnhU7xl6U+cW35hVT/8nF8xqxztHDs
8FNV87hZ00xLAgjeNNk4fD5muVeIvg2qzQyi6DVfZpIvEuTkhd7SOO08W2UE/f+Y
qGWGi9yeBqc0bzun/hGzPa8LPSSviZgdIL0Wtm3BPz/+STO/h4cUfWSS6O3RfSIa
nAi3WeZTUA07MfkGxP2ovq7HOI6iIzvMD6vmpImGVWFB+Sh4j86zxcE1g3WmHU+Z
nHoB9ldo1jogKsyM40AOpI5xb/wWA3+17MwDzFsth32DTEwkS+mceUNUu+UVNAYc
a3KY+bSa6/SWu24gKzQtnL4TV9v3Ysek4dVMQoo6D4pQvsQLFUfIzaidNAkOvkdT
/Wi7QBOvQtCgjfJTII4XhiCLQrqYKG11VGMBEscAd5Ej6P6SsTNrxZnTTdPblmvA
7vfSmeOlkv1mZh3s/bL0EZFhn737grrjMQjGoovb5YVac9TsTNqcCfcsA+rusWY0
2b6SLDnQ8JjqdogReZ5E8cYCScELeRXcxsnXxr5sS+M5fkJhoWxCDk60+O3KsAbs
dZAkdlZl2QWxq0+8KHID/kH1Ch1hGmUggyGod9TJU820UnA967MDrSYThKT0mU8m
H6VRbKL90OsLPAkcrsDX4w1oDG3/HXXTEXjKU00uUfDqEMFHPECOYuQfjfrMCpp1
Er8ecjcgrWhhgQfm+cusv1cwCtXTt56dSBFAhTaIBmGNmmhDTBU8RTABlOn4T76X
yzSn6sS7fpPgZRnGSjFludhUKrV3hqNQxDvqG14SllaJZBt+0Wfv2MVj4eNrwONy
JF/vT1w0pFsMqg24S9E2/zwoqRhWgj38tOCi2P790GO7t4vV2hVVyYaLCuLSlNBo
emTQhFnnUH33dIR7bHgeXwxycXfqXzCqNVy1kN1AISNwHzwi0CtIisIYF+WZxqxV
mRw7SpXBgKbgcmFAM0IpRwXxAr1gbrGEgrWrSy0fjNctkY4LMEYwztEDkq+qU4NG
wPg4T0x9caQkqAOFd4lkCuchGFxP6QYGS4mSktrDnXSsm9CfGGrI4/mPvvAnKEVz
d0FdZE58qJVgh+w0l74KlN0BIZdhK+z7wOpMvjmhZMXOzqCW/DY4DOmCDwJMbTYx
NX6WfYcCKtSjIQtL3uGP2p8dvTaEQ+A3N2SLu7zg8bw938BBa6Wmbv6ecwNsUOLJ
kI1fBZHbflTWsl6xVtIVY/jsCJ0qZWTaE7dcdYL0eKDhVt6qTXPvZ3nFXqUgM4dO
l0BjHwW4ftFBmks9cNlXH36k7bB72n3LdbcP1psXh9zUhdNVJip9Kv+ARWTq/2Lb
Yg3Rk+E/djpvT6l4G5pDTBSNntR+PWoKDsl6oYqhbPJ6lIVqfsJpqGID9cwQfnIS
aXqRQ8sEY56ZjRTAvtYOd34JEDsAZywJnrraCCjlX7CkYdHP1656+KFAH8efj6kK
2p1cTTFnOpiNrqC8SAsjOSgYpJZYVQJwDViktLy7GueZl4IzcwgrSnRtoyOSSJHY
HMgaVABAyg0PwYowIaPo5VQQuCm90jXP9fw3W3Y7eIMPF/5ILoiQgsFWbu7pk1BN
YC+zrY9Btr2pBpxWo1MYGP9TzWPrmg9hNhmxneyPGRDtwQxBOSErfTTK2zQcmfm/
qacaQuwOZUnu1Pz8nzUmoD5CcNLanllen9UEr7tFC8qSzoOAkTddRWJgOfgWZvR5
6mlYSzN/VSV9c//9+eGNhCpKXzDCYzrU+pF21Jha1XGDCYD8lNsUWW/0Tc5QC513
RUFecYLRVxSLPRVS+atxV39kzCK1gPwvBCTgR8HDsTrq+zwF7UOnZ4txwWNs5F7d
INYV0akDKB22aKG/grn7r4BUDOv+O1QtFy23eBq9dm0BhhFMm1DKeGueLNjfaBtm
6OMKCrP5F4UN3wXZ2zowABUdCISc3ao+4NMPXPfLuJE8fS5gjNqlZH7bsMbxsUCd
8+dxB9yVQgq0OkLWN2DS4IikMR+qPPoPeyQjn6BL24a6S2i5SbzjWOoJWxwuOc08
XhvpT98fTXXL/GcqG7jQqYyGoLSTKu/aD4W34iKnhve2OEoJgrysHMRGDZe9j5pt
guHCwvGr9uJlPmchHM1Fste/k71q0NvNIp3DF1exeKPaPQO6CcLgXXhXgPrZbwGL
+Gu4U+b2IQCZBIzGWeBDwcqvn37/V7pWjZl4AkjEbyVOWB6cTEqy2M1V+vo8BVgV
iPNzf5IXMWwx9HfXfWynhe1FWSsQYAJWS56vRO3zu6YTfVEUOs3N3CjOE97JlrKT
xt/XdSmpZvGFTFHlAM1sKhMdOxAeUncGokqJFtm7y/AJRZMZ8QlEg0/HpseA6gdS
UN97G/xgMYPkFVxwN8wy1zMBpXAKf4ALIW5EL2NpCvKflXHlYbbzO3VjWYx1+5L1
ENQqwqxBu8ywdjHD7vj0bhxnUBlSH0z6k4KhhFU7C4eRnbfKGDUulOWppI24hFW2
S8aVKaP3hK7q6QzqFvxuElQuIHLwUKo/AV42rGdGVQ5ZJy1EcsBEok+uSXgrfX4x
59w/V29rAYkedpV8XaZxWpVIAUnuESZ4DFag6Y1eMqZjSaNjy60ME39NNf2JlhYW
UhoJd3SgdyJ2e/8MXrH/KYtibQBGohdRu/oPbnu82oKJe8Ie7SvNK+yj63iybvfs
vHV0Kz3ff8lgm0eo3uAMjkYie7yTA6Eoi0Vc/jfgTZu4JmskDUwIRDrXGYvrX8kB
3RRjNB7m7FCFCqbUObfUWqcj4kKBuglIxeH0Uw6PgCbyIS/QVdhy1MqAbr+KrGVz
bsVsYXNWNKkr1caaHKEsN0zvwU7rGKKVSi0/OhEqmAT9FEM0JWWjd2S1dhpsnOmH
LswlqQi5Uv3+rhEGSWR/LLa1NQpeewtP6CF8CG3C8mBKDCDE3siJLWHC0GO7nGNC
+/y427bLRSFrGpU8LXvcyuCw4+lnj1JX+bMrueofm7HOQDALGQh4X03yU04PnnqW
i4sSW5bxVQrO2ZfnTf5rc3G8bgyIYKxBd8r+0MAEBcz1oNrkkkRTrbd8tg9A1/D+
Wyyo6i1l4JJ6tgpbzCAHktvFVHy11Ipz4r3zT9uDrZoxCv33RCGhhNfIBvQNvPnE
/ldVHapn46VWEm1iZB1zoFWc86Vw++5Z6Bk3XFh1gX3GNN3dW/8pUuiqivjE7ZU3
0gQUaSsXqWPL9GxnusQP3tKcuHJ5lEOdXsNKLyuRmWVtE3mWsgzsU6dv2vUuAhQT
yi7Iybn/pO81+0YU829f7AFi2IXaiiQvPPIfg6oks9pFtuvnkkrB2ctFjwfnPGhd
HhcnfTpgze3CKAN6Gqp6qHMqV90ysinM2o9KoNwkjRwWbCkjGrk/oprCQH8dEg06
ge/vvAO2Rc3bIpV6fohCuLWaxvmubxSC5Rl+qsy1thkIZ9b9RWILS3eSfBGrzKQS
Ys79k2RhGWK5ln4r12ZHqbhh6Rjy85XpNRkwuOKhwpTCKVl4rk0lGqYyVvvcIUKC
N1S6cNK6uM0aG9w0kVw8IA9gncpn47eeUMHevsmNZRxnqZAH3kNYngCukKmlW10j
RwQMnMdUGywgO5oYDrtTVbnTPZ9tm3ly84alAX/qUPG460Zv63HKKhR42Se/w7vQ
W1eOcrxKqjY70aqD3BkQ3fGDe/xLLRZ0IEGDJrbCTUFW90wp3wzjXxS+0EWGUWBM
xtmkFFpi3HQgckHqxa07IIEbxGSi9tbKUysVwZoYN+enJJDpb8YutjZ1WY5CP7ZB
Y8nhMkIMxCDfZCWag8k5ZfKUPpcgS9YDEFYf20CG8fdf8h3te1kn4kdHfOyidxZj
h6omDfhf+BhsHHxTI0ZyJcutmYrGGL27nuZlHOJSnpXHr5JSK4w7FTyKR4xS1nPv
3LCnHj24YOgM/OTuaWmQEsmUSlazNNbVM2rfyhU8QCQ77v+qqBTvDJK8qPsgagWV
4p3gNsd+rnlF34fX7ABtIL2lpSc8QWUb10fu0Zif+1YGUKHitGLHAViCUbcn9dUe
+r03Djvy2joL0veF83s+H+Q1yv07gFI0bfUXtOoclynbFHCBrb7dCY8+s6rn7ull
hW2LRlVETzE/SoMkle3KZIqhO7Wv+vcaXDMnYlLkySSoPQvYFRKR9vNMRsjTqmdb
tByGmj7S/g30/36lrPGFtJouvX2bdWbYjX2LXGKgsp2oRTiH63RqGkzdXSCDqfvn
Dx00GOzy/8hZCchfFIPAvvUR3DzukPKo2J4Wfcvd8+Cn1Ud18AR2D8CjkgciNvn7
4xXgm3YQ2hW8QyTcIoXWq1HJJ/2yVAHQ7R4XiYATE0SSQx0u3mOgF/A5oqCTwAxx
VKT00QpykQNZUYo9Y1aF6JoIKjfq1vrsR725Cx9/v6SWlzWjcFz7D14cMErL6U+u
wf8lpxa3NikYAECKc9Xsfat1Qk3246qinoTrswjfEIZi6AsIxuKdzAz6/yf4uw++
i+vn3N5IXAb1kHhSGq4RZ+xotlbEQATB6nnlEDmMKYC4nsB46viG1b1M+YpubKbg
bsnevya5wMbvBtHpdo2mjCeenM4wFxZ3H/mkpGqVYZS9sTwDZyEtawPBKVozOvE7
lOmbwpcir43wbZAKokekEkQzI8luUZKJM8ziKn5Ss3A4lGh4uXh4RTk7ipfDZv5o
DAgJO2NZ9V1/Vf783Mnt5AbEfycGsiOF/TGtDiFspNF3xKd4XzGcZ96MOj8582HA
/K1LpOGtcNnIb1cnTJOQGvgFkwgxZlAi8Hy/TI91mhY2GQ3Pqj/NtGKNtmHk2NjR
ST8Oo0wEj2NBedtovW2yz55RxcH0kCgMWYllm8cAMLelWI8njwWsjPOkf0pDtFrt
5lsioHHM2BapdWOH0TRnPYkIb5Tf7pCDzwfqlhD+VWhPagBas1BOD9/tLva+wwCC
i4ngBZJUFIqyeAVuTlQnCTBVuy0HJh/Vx1l9CQ4sc9XNiPW13UWX3roQGr3IE6PO
ZT/HJ1ZaOnYY64olK9/ZETKTzR0IA7004yRehTLju1EAaDvU+3aWfWUm62+J6a+g
FAdF5HgVSNl+jyPOpJXQHXK5g3lRXXAbs2sVQhjqwLPoROI1FOKV3pSNFNxvYgej
iGLawVHT3n6VH/W7h0wSdH63252sfE5nsAfUczfRnmuceKHh+QjlXWk1s5/id9/n
NF3MpEqq3mgafcMZYVZttYr1uZ+W77ebDq+smIOLlbP4ugc7x4zFvXFKiF7PCMyf
8/szzpryn39ewbmZPvR6cqtxwST9xusvQEUlrRRED41HWny5yDk/1Bb98F18dH3Z
CaBPy2ZJnL5nExoP00F3XJFRicHRIe8BxYnqWEwv1huvYVCTafbGUM63+doxSnSk
UIKYzxeG847ifR9cGyCR+Yzolehjw2KWQyeiZVm+uTfT49Iuw13dZNhBQafaK5mQ
c3xyhtvOWfwImyB0j6If6SgrWuq+LNy5yp5sC7Vh7nQIqUhlZpslbGF0GRkHje8T
uyNatiBRsjgED27GArDMONyrxm0kHCg1v5LWthI5DtMMGhZobbmS+w9FZv48xffa
F9ilhyGcyctpE7LwPzq0CKrCT8baOSlnOKpFRxn5/VvlIJDsF+1wQKalIS+qCxVP
9NQz5VSZy7P09jkRc304HS22NjQUnejDBgVZrNl4jp/r2ToCwvuT6Cozg0l1B/1u
zztfWNb1GiDM4L9t6S4FSwmihg6GfEEwFDyfTdlLegtqs44p6nSLzGN/zSW83vRD
NfFrw87/TbPYWGP/mos4GNWwIckR6gQ8l5P39dYZZyngi0S0WZhXMRg4hGZe/oHm
joqbkqZmQfaKL5GWsQyuCUwMbCtnRDUOkaBip6c0MSA/CX/wQei1ZMq7Kf2tFGCk
7u7U1ZnAeEQTNBEW3P+T5x2qOS6xObLeaIQ7csN9QTe2dO5ZuoTxLjpB5fyYqUT3
lQYmqSIj8V+P447wsuSjThaZ015opLkPDHlmP7jANoqHHsDePAw7IBfw3Np93ldK
jdRIdKpeAl5/8Wxemllup9F0TndNsLu6ivI1DR5odZDReY7HqQ6zjHrT+PBbmYZw
8fuvRYi31Ja6z/sB5yPIHTnUI63fsVT7e7SnQcxDa4+b3gsK5zC/QbK13GhXDgVl
9rnx8H+nUGfzyuuqB2PG29ZrjNHbGg6r3hlEek8mgikvj8UonV3WBn+f7P8beg09
3tqzJV9jVdyDleSwQT7llZbI1KJGcRY7C+t+yybk93ZPJHZ4DoW0yFzunL/DY6B+
A95cExso4lYLFNLWyK8rO2oYW5mIZBoVDF0yjDLCZTn4pDqN1Eb/4l7XnP1rhVjI
GZmsC/HRI/9iIivQgiuuRNSEApHwdU5q5BbWI5LxlE9hdGMuqd0LtpvAa/F/jgAs
Ym7iiTNwIc/GTRiqGj4iL/0i3g8AZ56ZDhKIcpOKhQAwxYsa1CZBEHQVMe5gcE5n
ZdyUai/WYpXTtP3h2R+HiFdgIA3rUTRKzoJ9tL+5WwZvCVFdeTdg0FDYgJktRuwz
ACEz2Vsk0KaU7e4e8JfzExCfD5IkBvygaIdF9GlFGnO8TRD5vMB6Vsk6hH4MAe58
+jg5LjLz61H9U6B7TzxYP8m83lei+ligcDnAq2qxRGhhbq+Yw7vCFgtCtFcKg9u5
jwFIAJE3vmmeh2sWcDzSppOjiRsC0NNUIafQBp5RbWMBgEiKDVQDYS7bbnsUpQiN
hGEBkI7p4PWJc6q3jy0OYsyh1lHBbUyZyHGpFjf02h3Fl5BlkVL4i/TfLA745C/p
DVYa8tKY45aUg6WGeteSpl1QvHBkCYp+hGILwi7WLTxebfAn9uXqE3EB10WR24fe
7yd6pMVK8OIqboHKJ04jfBDF1vujtfRZ7l9UXq02nCApg8hh10iPrRyH8MxFCykd
MHdsG5YfF68wcF/hTlsWjT9cg5USzGfZUu2ghsRb7VRCy7U2zO1TfhP8xKYrt+xn
70WwFz03+1evTDm935RdTUCcskRXKijhT2cnO6aI7Rht3QGPq/AQzHkjj7vD4s97
xdqwwHb8Zea0Ul4sYbv0B31Fb96u/qZCUF8tKR5YD0nJZhR+zdUdu4hDhLdmWFbv
4ofZB46Db9roINb2LYn+4y80NYaXXZzpUniKf8vps/Lxj8zJrajik71U8v4vcj/8
2cCVUtdvYFbwnBUdSyJFkZ/f4QgLYb6+Gg2CT/zM2vAjcOJE/vv4ECyEyDftL/Zy
880aa0Rvk9AlwkDfgrN7oL1qfWCO3L0DMoUS70h31DodjySKBod2h0Z5lcSuXEdV
Yy9JYJOKbG3wFMm2TjUMNH/T6mmabVCK1pgLxMNQppdKqOPxg/6julJUziGt2R3H
E2cVFD7OmKS/abomZuAHM1yTzJhTYRfnrQwemPv4yewnLat7IunwijLyoj1SGT4R
t4AvJ1OZNcBD/zEoZOgI50GhsvL7X2jBcji1JSwLQM1SXTI03LmVmrRfnZPX5Mtq
GsG323mnjb1Jf9YZclu2rpGayYDUf0Wb+gP70ufsJJDTchjjYjoN3i0ud/tDZAot
kx8AmhPx8WknJUiW7CsgVp1+TacjYfHeMASXNyjjhOGl2H7/alSnUEitk2I5wkwN
kGlkb7Zw+A0LT/J60cqo/dvH+jH06W9cRytISjVL2uClv8LLUHii8YplkfbrqK1T
jwdW7fFPc2QjkZzoYY7IhkaYT2HJX7rRKhe5MRki4FVt0UmK90PHxahHQW87fuPT
fCj8urjBug5lB+PhqyQdcRrBhsJU4RYgwJZsuo88q7Wutc2g4nk0LP7VXKHQDe/j
CVA/Fc0ko2fMQqZVq3E9wfOlVMa1vEgLn3NR0V9eRIJeX9MolseKGGU6CNdzayyv
/bJ8XE5On9t60agYUDIo/ITvLZ3fYyAcU0klMQh/4OUkEYH7P9MmwD9GFsY5TEv2
but+0D1cta6SVZTQRdfgYZcBKFt9LEGlUndgBiUGI2KlKe4h2qc5GilLIG7PD+ga
1hKSjhH0NJ2ptPfdfGlOJfmLVwBoig7NmsFyb7tKygAGQWkC3CveLqwr0OgOcNLR
HheH2vA32n6IUbLtDMXnMkdxQ4TlQa/y6HAUGblk0uSl2qIDk0rgXSk3lFgbWIk+
e7x38qXKkVNhoPr2FXYP1aurhGnTp6AZxpcS0mLLOmWCp06OaE6la7kXo/Y8tMb3
Kmwk8o85xoYOZsW/KOkV9vM20K/tlj3oYYyiz2UDg4azuY6ETG7iPb6Ayoi6LBFy
U8Sqlj/ABqnaYqKf0Wt6BAwBhHhF9fPGkso7wu4F6BonwJQKsFeoZlDsLgYlIU3J
oMat5la3knyz5Q092AmuSnAuXheNUWdY9cS/K4Sj3Q28VTU5vO0xsCVYmXiN+Q1g
g4kBuheuP4ZZOg39M2lBFZygmTStGW5dAMNXWrACy7Q+BNCoLx6EPEvcywzQwxUh
Atjejii11/akOainQ8XzymVgr5k0r+QrVnebmuehe7LkvVnv0adGACMidItTmDqi
4MoTzTucg/fzFvU22FB7FLsB7yTOcAlD7h9mF1Cgg6fG5X4X2JPqqsFTMHbxfcde
ee6nAEaB0O4dACLLVGFkKbg4FuoBHziUDDo7OiduWqaxv4wFIP5AVrI2tlNvkApQ
/YGQ3QXDOoLQxMv0VDktJpNL1KNpO6xuPY5QADkaMX8e6innOSEEl5ix0l3MhdHJ
urDvCrqe/RT/QFMZ01O3pZkRQOfZfj21/EGZqrPtOkkmrn7pqd22POHLe4naxRBx
v2+w76hEUWloPyywXSqR4OGYeOc67hitdGDKQs50NOcawVLtI/eMoOOZ7dpK6izO
RYV5Vxs6ItSGAW9kC6VvUf+MmG7vCRORyLoXV3S+2hQ0Zips/56P1CQFtXj/zzwY
Is6VZQn8PXW8kRsPkjjSQPk3f/W1JMqlHX7tUK1sebDWeX+nKBEzRHYioGSmvhCw
k4fzvvOplz9VE9bgE62uuTMrcQVwWNAG2GrAIYbrnSCSk97q55Wl638gF76q6UxF
nolHn48/u480SXIiEKkH7avifSYhvKyo4Og0AeAY4Njvx68M1oRLqxzrq7XYLlw5
yfpJFFgsxYWo3+vN8oAvLA6aXaMgzcL7vJplnH0sQNbrt9UA5AnTZFR0bG/Vnen7
5rn09lu0yllKopDfXw2mGYg8tuBgSlQYRcaMuv7HBnzswZ5ij0QgeLgX/ynmSXx4
jXT9qNjIYShrs9W+TIdfAvyDfz9kHMm1G9U+/zaec6d+Y82C68zI5/EzE6BL3SF2
6yVjhr3btmOwWkHj7xESeJh964gM42LnKYeP2kie43VS1cdqzL820p7c7d13nX2J
KqS5DfCcqkZ4iQc89rVnTj8gyiqddG0qqmmgqN3Z0llA/1ZqQODfBWmgdADJdDfr
8Mi6n7oe4rBMHlWws7I7I0BNFygCOUSc1Jvnr8Z8SdH1uEFDSSs8QBNjThw51R/6
MgtOhtTGpK7F7kKETxPvMcx3I0ytfZPASZBws+KVgIOXBMv3dgUlTX3ngKoHyXnu
fBMtNPK6nNLM5I+vHHYBu/6ac541wa1IYU/J2jikT5aVNx5R5UZb2G5i+WYV7P5h
fgxqjw4D1U2vNucdLR2PmQB2m2yPOCDni3sLvt30TSNz2e8YftJdo1otDsk/IR+m
6xIOkPGrR39XzKBPZgfVt4RpYD99xj3l9shs0nBy0qqZMPcwIJ+Tb+fE6f/ftVKq
KzxQq8zpmd1bwDKQaf1pR+yh7wP8X+MAwTgW1NLMdFeYrWigGsNTVhgYUxkgMp7g
3C2+vN23pwfd2BU1mj/7T2c0geKGagCZ652+CKrVGmcCNfl6YX8n9uzDzscFUA7n
oAviOVTSTwrHtX6THNSY0DYWTV7CTnNLPAI3puViP5ASnU9MLtIfSAVz6W6EMPJK
P/e3BG+U4UetN1bej2vHUz32crTEzEGSq3fIe69grCDYz5qGHApNdwaF10bpUdqA
GMEqX+IzQ8OFsqeHKKqdGDRry2NHkqtOUmaFhQtPmtqhSlUxwAJ0NNKozVcr7Ci2
anQFjWCNL6T0zBngYRLQoLqtOKuz6XMQKI22McYMZSiMrWSz3kQd4x8DoMEEV+jm
u5YVkZSI7FNrD5VprskmUYhu7IEoJh2B658uDkh6llCjGDwW4dnElKZa4XMvT8XF
RyK+0DJK2QU4Qxy/seNf+TG6KhjnuwUzeF/PM5a8d4WqwiNpOvJ1/zrlrS2BaQi6
x2W2Ua3lcKbcEyA+cTXwpzu8oyms/xsP2RMHiN1mN/NLcrErOZodvRQ8dSAi+cQv
AzEmpB/KBQfNx0WUqfinPzjlEnyQ4WVXgygLVT7czlh4XSz820cp/YOSfd7DBcgZ
d1p6aPJNGODIAdQpsyKDCjZBZvwpW3VpKqQBF2ZNLi/uiXOESUtb7ENfTmcle1C3
SjClscScykjUKB9S257qFfPeIO8JdnaZSMEZLdO5qBFbF4MgoabUbpeYUs4O56y8
42X5wFClVfyrcViqaY/Fa1C9FLRzpnF/h4y3Zl1nVQsQfSmzz6p1AvHM6dD7Cfw8
BS517k6o6BaFXvNdCUwhJJNHnL+l0ZeLfLTTvMbuniVxLpbQaRuGP8DAIP7e8OLL
AfC48+h9dAmBuHLvRot54KWcLU6uxyfX9PVdJiVEvLTrU3pXx4J36Ism4rc7jaEs
Y2wfNPLauu2gU1NmSDZf6F/Kinss9bCvuaR2Ip83WYcSlG+AP9Scvl/Z35FPGSYY
7fdzghPBh2aaCEFcXDnn3Jw0IT8YA2Z+WHimRDtjBPcRhL3P8DIZA85x7U3R8N2K
w+ezUThH/opMDbYacc9ozGpbBeml3mEY6r1VSzUIJIiq82iTsL5IvCrvvzJZzUjO
//hgXN/weQMqHgOMjNE74YxhR8XHqSgwIjbdXQi011RvKGxenOLNO2LHjGq8K6GT
CkMQh7ov5nP4mVlVBKZiQSo//mZc6PXGMEHsoH7k+5f/YrRH38MgnM96AzUNlkhu
UGn0Y+5CaFyQpjx8X3V7g0rDU4INASGV/gP0jsl8mfIPUalfUWgN3szxZd4xaaab
g/7qoD4SH6cM9xMXkNPmPrKqLgS5POTBuZhw65XMMQbnnoOIBcGal+tjZrCTJ05G
devsNSkpjXPeOeo+vsIr+XApWxthgftAa16xREUfkhepU/UY1CWegNYYbCEU+wqc
lRyxR9Ft49DV7iuUEGPMCXk+4Gbbcg9wZN+5iTTDx7b+ngYMadP78AX9WpnyKLNr
9ZXWuB29fD/R4SntoL7riPlUr1TkCNlih4vvQGQWWRVRYgaFVsYMKUVCT4xcbK51
Memyk9TKJsg60sIbV1MvaJax9lOTyn/WOMFahmslarpwfzTfjeBQa00ZFMW/bthT
/3rUDPGDgHbgShG+anrUDpRdANDPY1wuxcmxsmg5Q6z/Fu75Zb0uLhiS1roU2BxB
u1s9sm+OAwYYIWW8lzTHkqJdB1R/z0YzByUjIBkPxGtNJga7A1Lkyz71R6a3hqSL
T9aE4dwoG5XycY3n0MWR/kwj8kSwnKVQmKbzgU9+Bv388ke4QvafmloV1R1UYFEe
UZ/vQdDAejyHNaFMRGpCnuer2JK6aX9K8wFGAYbrFnrIuZvWSLmvyv/gTxuKMJq+
m41tMiNSC4ij/J9QyxYzzZcUZDjJZKZz6TYBKVALbrNYXtfXX6kfOm9VF84uvnaK
vkTfa1rTvuZqU+6e+B3dU0vW2J9AgVkiVre9PWXGw+hvHBdKaSSM6fE6l2axpUwh
Ql+OCPRgeFqpVuH9yqCUgDaXPAMxxdWPXIdkty6Q2UJGUP8tjpfdJ2a5i5ubf54N
bu7u0QU76LTkX2ld9/ht7OGjMcLxUgwS+55ywvCLNCZycIWQS8Fiokiz3jLhyWIK
CAjT/fOuPtrf7EqIoEABlOAIWDqtM/eLkEU+e5byh8wT8WPjI4lej1HrjGIlAMEy
hZry64U73+YqsI/gbI/NEqS+JK4v0nACku4x27BLLTdpf+1ZsbZnJKfD+xbXS5lx
87NmhreiDO7wTf1zzNhoUFSNCKc/O+cq4luhpYQR1vq2uOLtZgshWsogGlrnfq0V
K//GMpxDMzduXDIm8zfpxcXYDJuuDVHZEBfQuRhnyoeIxzEk6S6fdQEhTrRmEhRV
59jcddIjvaRDtSADQtxtDqEIjMBByIz48uZQkbyxdfoDY8RQPVciIN5JD8KXFuDo
edg8+rVB+97xeMWMl3sD7GQF5uDJdcWmTfp7qrQF4C5HBssgDBqjs11eI6proOND
OgX0JdnMz2mRCOw7v7V1P3hKhI7yR31fX7c2nJYP7Lh0RQFuC28rARDgYBBuBe1C
bJgTRq2qf5OIMbTjL80XCuP7HVre6RVEluTGWR/LX8pCihJR7ixemA8JnVZh9dJo
FpUib5xZ0YCyM/DWHUa3lze5RJNME7KSvZ41R3lCoKRl++mB7BnUZum0cYfR3Clb
zG/tRDp1cSUtft9Z36UVanJTrCk7wqGgQdnVbh4CFHD5VfzGOGh/s7hEdjWtWnyl
sdaY8g9/vVNPHgTbuuSWkQOOpXNGTRViSvI1G2bGLwP9jUVpsz2NZoKxVN5Br3Dn
MLvegSfKgoVnqfzk5sM8EADpJjb8m1++klt7mpkUDea0izfl2Eq3Grz7HEbfwUtI
JstnapVNbN3xC/Yi6e+SPrvnuuxmrLB4vk1aykc4pdpo6n/hYY+WQuejIcj9CBeH
9glT+EVJ/h28PCP3bEEsr0zXq1/r+fyrPNUOJ22ULDTBgwG2R2/Jq5t05sscgg0H
JuR7rlhq0pC7di025S8iFx4k0s0dDcephRunxPVt/0H/Qe1cZHcG4zcGZJogCtGJ
W0kxP/XWKSfQr1INrTKcXat48pwS/9e7JR+tcDA/UAnsJJDj4a6hOrt7yahFOa+J
lcrU+v0qgFeuxle0i1Pxpcursk9eEF6UXFSLv4fibgpPnTuxlIaxZTXs+N8b9n3x
3rOE4QIYwJQxCvcc0Ngk3msAlku/cmTI1WIzRExElVkhGTESaUVWxFtXhfld3YUQ
5tjpz0pN8TQv//9G/2dQL9ArIGnOuStf+w8n6aINXhR0FBebJozeZHXbEQwRsp/Q
kncMRjCG5DW1B80xHF2xlgh7/kImYnqOJee3y1DMTEojy8PlBNdD4iPLex0fFZP4
o+vL9GoKyFfPeVGJv3wwm/cwGNAsvt3rRvgv48RfFttRsqF37baww+qSmOuCVjl1
nqEwpZALacOFkWcEcqVtnTs9n51XVVMCBjptzEonaf0NYB1Nxg1okpxiySArTH0l
NQdpFbxvcWSRA1q8iINHYvmTkGl9163OUeOxVzLhRbw8IdCOysw/zpBR5YmKb739
gCW+Usx+SGGQEcuPDU1rErxAi7uxaxAsm3OFimHpeiO7/yDe7Vi41uteTnRKjMn/
q8XkOVJzoKULbXbhPhGdfkxXB4hRwqT88P5ILbIBgcm9oc0zkwAahCib3OuXzbTF
lcGqPgbKeRoV2Rgr77M1v3rHuLr5zNmEVUx6sK0WJDd99rMKJm3gEQawoKa/aU3V
3dxBwne+AvWD6osM41MYcuOvqGkseU+FTTV8abnboJEWvZIKDRrY7Blj8eibP8kv
tgawyPIIvsNV5jJ+Z6OwIe1Lnas2hW7USgk+LlZpf7ePTsdUv+5AB3cZcdC3QOL5
eWciLknakbLwNiES0MvF8g36PCpBj+ji3c7KYRgL3BXBqiVYpCUNpqIM46cSVp5f
RRkXNsV0haWMJtBdBjA/zLe5KaIA8U0XvclJh73KfT8WH2RvRs7HAWu1PR7Dl8hI
to/KmXa0KLUxU2P3kEUid2fN/0hpNtb1Em+EV6hNY/RXw2oyHTGsCFcb3Eko5Z84
v0l0qIib/BvDlsFcK/UlZd+E9lA8RMTFJeXLzgGOIh9rETRjAarBr2L8Bjgg1sRy
ErhMORzk81UQG76QSDXsU71ZfSwvN+oxp8/OPkf5ChdElt/g0Ck+NfzKXHtutMsV
TjMHi+RrQzAnVQjMtBBZw9j2Fqj6+CrJsL+vQJD29yEAFmHZA/yhDfYt0dCzXKI2
iahgq168LxqM4oooLNoeeNjw8IgLzzxk/4EQ6bQILAePx13cWxMka047M+gEjh5P
4180ldv6hiI1SCXaOWFE9OpUDznEDmRNq9q/0ngo2fZYJd/3CFeBzEzuXYkCBBFq
/qb8Sgq8S1AChLD4a/E1aKMFWsy4fHmx6FGaxbnUZ518csmNx7kUCeKm++S4THD5
v0AC9KWC5muSd3EFOUxtoxsEcuC+oLoXp1byNA06rFXvNTUGCjPrCjU3vzsOtVXN
lBfxLQICZGCMfrelQAIxS4E+Zvzc02ekm1Qa6MZE+sEGEwZKrVS7qEk2m5hbkJaP
VesKOw6ddeORTDNsobe8KBJmQlwq9uQlsGHxe03482jY2m15+6Vm1xKFByejNrv4
mRhDuM8Nscy3WZ8FBW8W/+6U5iDMcZZYsAEsQsqtVd2xuIOLWfHPx0okT4WbV9AK
CzPADw1GPJzx4T2xOGtDRtjr9eLlN7aLzEZQHMjR15JiHr3gnkrawdAcSMVGGOHp
X7XP0SpgE0GB+H2NYG5NMW7tZuHfAySteoa0ORjA6slqainaXSMw3xzBsxCrRIJB
nTWKC97juKdlkUKREI6bwW/n7GY6ldH5wu76zO+OjsznbyD+jhQxS35kSAzOU3ac
885esV/U3ne6tiJs4wdToIXb+XjnPX53p+ISu1Zwjef9vEbkwXYn9FjmVllF2HVr
aSDo98MA216NJ403qYYtl5nSGyacCC/aK2Gf6lepyMoCeIS9giVQV69c9eObgcn+
gYsBqkuSm72G8xUIMRw+0Yhj1HuaiTxyAIqPZH/TLTHbl8NHXNEhQhSK+XvHez3N
m+F1M0waG28EvCmauKOut012b/tpq5B4RiXqr9kk6JNu1a/On2KZTGPGJlu7Gyz7
KvJT3wkTYa7h63X+FrSsnUdzttkeJp/hjEdLhHg/Rv8eGsNyd2hdJ0BLmfBmdga7
EPAgreBVvfRFjSXwXGikgt98Uz7McZhO/qXbZ4BoEGRSgVo7wZ/BE6ZoQA8bsz3B
8AmtU4k/YvhFwne2vAaer4M2k0drbXRri2UfCMMfBgrS+TzZQIcfRJInHHrHrioQ
k4uV5el+yRw0bj1Hxh+HhLmI0uZYl9A0fQ4VAOD5JFM44cYPruvCaZfWQi5NEM9/
efayNb5t/7wvRyIcuvDmisJ8wF3qPZe32EtLpCs2RvaI0Ado+bdwMQSq5+y+LS2K
D70juz/7O0aCGk0ybwlxrQKVIvT8p0aDBDhOpeddMaXHGQvsm30l2i+NVMm4sGNH
sYBfONGblZ/R9cJ3kuN2Un4fJ+Dyl34I9K0gwBaYEZCzA83SQiONTqX1mFGKJBTv
VPoSgiRocj2dk9XImk+dJsTb00yH+C9qLh+2Kkq3yY9Q0i9WjhgZME/CNUoutAcW
VFJrmRYQ4yQfQywuAKfL0Kn9rX8WkSPZLDbI44n0YMtYHBh4DqiM5TbgDnoFqE01
rTUZY6ph9+oYdhjbRxUVJrIJ10ahDwX4nnOMRUR2tabrddZVTIaeNmwbzVUJas9C
XlLvGIY+PIcMpMVqgQhIrUMLMm77D8HbL+nyzXyagDK0L3Ez7HNggmchzRBrMhDZ
YFYwu4ed3dVJO5QTCFJB8fwM09JKaHpYaS+qAaJmWoaOssppJI5hkzyAFlkTr9EV
bTI+qq70mGHwsVBKdyeiiZzU9+nznRtUPPlNVlfOEZEbTR6Q0bjIIOXXfgN1R0h9
GRsx1uUx5XptPn8nffUtMGKew2V4xRRZhPhxZQog+hZjxfF/PwArCyu9GSGH/SjH
ZWNUpwY3yUy2Ov1+c18H7O1u9e4ziYzXoe/GGL0bVfduqfXS/9tBWlh/b9MsUkBn
n0KwC3ok+Wc7LS6PRiJW+ulCPCALXqsQt4xFYyMPHkgOWIpxJxjkAlvlzPpDq1Yv
lmtDwHL66rfhhOuhMjK1GeF0VsAzv9CInODqgD1CVImll2tIfpczOl3AGQwPUKQB
tfU0vwA0lpDF4dT5PrNKXA7Y0ZmQhVZOnfQfvDIwa7tkV6IAzJ5fyEkOYXvPoggE
Aji/wkE1Y4PhZr9tHsuC3jQUlM2Yctwv54rPfsREI5oRVjwtEq0t4pqqrCxoKnv5
v2Rs717JJ3omYp1AWZte5P/DUaq/4daLFWMvC1HlS1E3ecG7vRZY7cFKdHsATbWp
mZoCcrPKoltql+nv51HV4VBQzM57LABHcawxkEMPzHPH/2QOSP/0T4ywiAbfJzmk
CIWDbqiH4lbd244KvQOd7IbbaPAtrvQjkSgyW2G0THhYPfvZdDJbk1phEVXFnW2a
PX84D0gkoAbmFidyJNSHcvZRp+3i/Sg9VwMndJ+GGRJkk0v+YG6iv+80e8gqEvsv
ywdiR6mB4Cv2EvKEaM0g7m4MZ/I8AAjwb9DqKUlIexFAnWUuvOyBpZGTKuMZiQFl
C7LqFurphfRJhuOcY5U4CXGkUmODiADt1LsDxcjeUH92bVRgZEyo6yDotxBKT9+n
NF0l7ZsEuXDU8b0zV65jjnULixr/RbD59lOd58SrLL8uFYvMuqZAYcWJQofXMjin
hQZ8sDThSEQBjhhSrBjO6ECy1GCnneMLhYnKoPTPW7MohJfcNiWjOca/qjeR9Wqg
ZDG89j0VaDCweil2gauGyNuG8JhdAxR/DtxUybCNs/ZNksffBf9KWHY6m8z1CiCQ
QkGUJwcCzSVG784S/y1mhCAyXDlBU/V1tEiz7TuQ4szPlVKtxifLwk3F7YB24yaG
Xieoo/EIF/iJEJ7AUtU4MFkNEmsy91D6JyfoCcYEwNsEh5z0tJqG10BbEwFc8Vmx
MtueD4isiqeRX/igzPf2OD6+ktrQDkFWfBBR8z2x/AM4p8V6jRkoyA7uQIYmGsF2
P8A4ili5ylUW3UDDKNErEoRafmtTLO5ec+6kvLbYsQ8YziW9/fRyWtMPd8wawGap
8rod/zSUh6+obbB45QCRFkr64q91SMCrvMYFL2euuOMiKWC7MSzC8FAnPHktobaq
ivOM6cEG9lrqPBlbPaXDvS2wVr62Kf8AedmHQWf9iW2/k/onLpjRwPdZOVC2XLxP
1/sHnTBxKQGtnutFZGOfnjPUZyaT4WE6MfDXv7V4vZpkGCZvv0udMvRpOYNTmHG1
POBmLfRKWSGQ9dWOFlA71qvoAqQw053XvHWAtFD9CQQsaaPWyDidt9jSACxn3PPi
PPCAo6BYU5TvNKpkKe7Y4hT14ql6JeoBGusItFCWNlkoF+gfvnKTQtO/pnIAhMuC
zCKe3WfXH2a8s5E+YvLf/EKp3xJHRxqfDRaZN3pb2q8hg9AUr1RKPZxehzzXz2dG
LDVEAzkGfqV5Lt8DShBodmk+6qFnAMK1pgbHaDkfsOqhk6iSb1vuw7ho8ua3mCPU
y1QHJrVt+66Guplm5HrU+gq5FlwZmoImu7TjO3wRLoLU+lfKygIq0Kk0ZW2y2wto
8Y/FqVEEuzRIZEA2Ene1+tbP+uvIWlvlKpIfYe4WUk71cx6nTcViy+yuH+FKYR6y
T3cyifUsIPUwnRzKQxLKuQ/bn4QnBUrDCT9RJFmCJLiJ/vz6iyn/8TzSnmorgbON
q289ZDDiKTt920vrIStNYb0KjQ9dRvuEu1wBE4M/AzVH+yxXQHnHQ3r7K8iE/y9I
yQkiX0RAHCBPT/U4yK6it59KHFm9tVDaaqajilZFL9aS1E2EsRL0jnnGjZrx5lzd
hWXX63D3enV00VgvGj6Sn3xiJZ+rIYATGrmjqKBunOpqpe0m3dPSV6jcDa5iTCHm
8pdtLXt9W/9fd1PKZA9HV1nvHNuhtAeoDVN7uCESL40PPenjEVPd2cYsWIOgnDct
pEhLEqB3+jkc/GpRXiYU+PTR0vLqeONyNr1KmxOlFoLU2BdnYdFf/z5BKwRT2qWb
tw0j9oFI0xOJ3keQA/0ZhvGrtAV19eVc34yZKzKg0Ki2MRQ1pzNel2JfzfLG/KsB
FwCoKg3J+rTrcdhvciqW4MjHFJFM6h5PCyB9RE0GTGl8rLHQK4W+yNGDBdtEQORd
uFq+8v/GcA9DiPF0GyO/1p3qlBAa9yuk+2DtoKepjjIsZh6Qk8VCs6d+4OdMFMRI
FJy6Njj/y3/Wmi6gdgb4MFaNNvAV59HwhSTsgQYXylBUbTkv7dDGvdpoyYWDaG+D
Dg/g5myd3w4pt5SKoXlxA+zDlyRU/Uu6Y9AJ4+yskD2Hf99WvviHrxQhUP3l+phT
thTZ7QaJ8bs3q57vjSoWd1j3xNhKDuWXEyI0BSOpBqt4JY7Ww0wUniI1QJETTyxJ
5ErNkaCTs7/xsZugIpg2E54uQ69wbHSC7hpHWsWHLs9OnZoLhtGQP89fGJXYQK4O
LGV6DMJggQR4sYx8plCNh2OOBvkEz6SvLC4jKat0lAg3mY3Xt53tWVfLtrb58kfc
BbWAr1WiR9k8onrJ6fyGcRm9KHA2YXBUubFdVM3SoiylVak8i8kmEVeb5rECiode
P40FgCABE9O7qQM/nE3v155CmssI7DL0aQYe9NmepIOAO07Je3GGxnXvp1fgyNtD
KiJTJ+JCzCUnn8UZ/o5FKAceEQ1RD8S0Lp82Oa8x3pIKdzHlzato98Ly7uDJ6ei4
75TitaqSQo03IYEyBvKOGXAoaDrO2UIhOS3iMgFVSwDBxwa8oIbSlLnu/kbYFwvy
eW8TePrlre606NKgQ8S7Xc5ZvgxFHmJ1MiYX5Qdj2QOQbK1Ych/YGfuSgp07fp8t
GVNAD8Vaim4Btp1WbaSpviC1UGG6+R6+/gE79H4EbGpVEM7597U3L7ZILs4Pc24G
KJRC1n9jeTS3AxIr7KqjHLs31JrzbHBraE7V6xmrAkUVyjCxA2fef65YhmUt5SxK
mQKdOY48Jj1bqFq5Uwc0WWMsmqf8M8q6wD0cvEz3NQQebam8IFbwI5e05yb6CTtx
M/M6sRfx2tnimUfrxB7qxT/yg/zU/pEcPxoDOn3Z/qCz37ouen9NdlcHQNuyImQp
eFmOkslkdBXxXCbGKmjj8pXBO26FptKP9lBOxnoKaCoB6Kkk1LZlgR5Tz6+43v8P
8ddVKh5+h6VGsSnLl1r+iCQvZ5a5Glx/vSTDsS9I1Ff9syJU/LIdavGhZF/8ITto
kbo5F1i96xv8S96uYez73tOeJ/mB2v9a0oHc9KTsFMkp449hZlWXG2ckhqpqbRFE
SVYWypxK/AQYzWP52UV7aEuU3dmhr4sTPaQ9xN6lHTJEynCXvo+TzE66vlT+0s2l
i06wIFrt/bHRxAnf06JzDtOiJ2k34Oq1NIrh+f5lUZsYbmcqGrLAGKs6Ygtbkub/
oSCp4oyKA/D56JFvppE88A9luY/Ubc+EKRatB4TepG7sb0YNTRbh4CO6UhGFFUDZ
6nEA2QaKgS0+0rjOcwyODwAtgIwSqM7iWaLdPct0/b4jNGq80BdDju2Smi9Q8zhW
9f3HIciQjMQKSI31EF+kYeaVWXCGSkw66aBsy1Ip1HsPUhYLsc4F2T2V3V/xUNR8
tZEzTW3TyrxkXeGzkLKOVM+JfHkSEfgPYa2N6DiMOHpHwmX4YBWN8L8pS+YHFZBW
srC0vl2pJzACvQRuDlKLl7rLSCAIQUL7R7U0+a3hKaMX9D0UBxufZ71z1pD6eUZc
z0v5SJ8vcWpcZr89g51jL3P7ydDTVFh4lUAo0TerqnMmoP0IIFH7HNUmJv6RAoO+
ko9XmY8ov1dRAv3YLSx7CYHkVQxQYsXvssQcOvcm5fnNqVZ2JIu/+buDNej2D7ir
YWCeUEeOSpH4BEcr+BgVW/306XQlVWWqoeadAwZFN4qR16h3d6yxdIQLWvK0e/qq
fwrc8UcQaOFfcs7tTvcWdt9UzUZS1+du1LrTy3FBlOTulrmfgFEDXzrBHEvgxR/F
B+DyTO+l3S4jE5MpQsJaLNq3kZVAdn4fAEsKFPsTX6+IxPq/N4HmLq3h35J7Tsmg
sxCYr5pfez4RYvqEUh/JCj69hfdA1aa5eMD2D4s7DiQL/D1gRXa+mjQcgAGMk6W1
ld1bczLzNiSoxlyYoG+MLpDHyi8VPN97Bs9Ktk0dmtNtwOo16E414EicyiRtpjPm
rU8Z5d6Nzsne5ZFi+zThwQlLv0PLUd/hovqa80/qMSH6lpNQUhZxT6KzFRkRmp9I
j3jQ+hE/cOIka92yAIXdT8OCScP40zZFNr4s59c4kUpe+PV0b09jvmBU0GL+9iDA
lwhZMt1F2uPh8nMdlfAZWvSrS5d390mZ2SxXdRM5EXlTpoKGZpFNT1xtWmGMW/s5
+kHqzVyWmGXlXhai+MADWIqmc31kASCPRnH/TzJevj0zgIw2Pz1xmAYBcsCrQfdi
crNqB1pcrPIZ59jl2IpMyY47iD1atEBAAW/YlEhSl9MgtVsqiZgn9EFRbWo9FhQn
CSO6pRyiD2o15QK5HfAD7qP+LFWXiPmNmbs4oc8/X9zNWv4KowIgyyC+AiYnUpyh
QoAP+UfXyE+7Mp97wGP40r/kQ1kzTj3oskerOuF+J9jzsu5vvmqnNLiwgC9X3r0A
r43gxnUrqmH6VJIMmzoWFnxGfE7eFKhxTItM8sbNrcTPQM9J28LZvhwZTGIDkXrK
O692MAbP00vvVyBxWJbcHXwm/T0bY4JxD3TkaO9HkJzWXwzKjB7+CaQ2TQrGFi8N
YnmXWiLUm6LrFCARhq04P59I95zTha+rItm2AuxY85L6XMeXe8E2s/M/Chykr1fT
8nnxiV2GAQuKTB+M6BfZCBKDb724wrsvXGvyasqPW8cmUTiMWTnhYOpKU1cqzam6
n+J4WjhhM/ykIUODbhTFeJg1sXzdo/Y0IcrIF3MWtSEZ+i2txSmMunpsGEGEUDyM
cB2O0ITmIlPMXjZXgGW1VyEZhCd6a7LK+2WrDTOKfDlRmcj0NMOQzM44V5nhoKkR
SVHZPXuFZgLtgdJH9NIUUsm0mLTp5V1TCf/Y5i6sefVI6+146conKFx6qfAWNvVc
nZjz3LYhBJyS0tXurqfFZEyoodnPhZK797c8ZGh5KGIuRKHGVZAi/O1Brpo/PsOm
dj7J9X7zLeko7VQred5WsjvABbV7nvNuSaAqm0o8ic731X3rpbpxGwjcF9Uvo/LR
gJgdGp7r84kcGY8qi7scrw2/9k8McGhLw0oSV1Oa1mywiNFLlKATz1L1WkuHG5Dw
04F4Iv9c6riHkwdy6HeehueWS8jJkhdP/dSpQmcABJW8kN5xt3PlXpgpHYkTg18l
/C+QblY04ZuAbTbt6MNrbn97pL6/tdX7n54HhsBW8D2p7ZeGtHPQ5gzJrexrxds+
PviDwhWF5pWoiHce53RVmPlzjYsKDd8t1cWq67PHTrWpkR3CxyhsB/BNEQ4x5jDk
YbEgjUtgRZ25G7DjuAlP2y6SZncODWgryHNG2gV1yUp9QrO85B7MeL6OD9cWjZfB
gVCIrB80OefRu4vYix9tzR1ZqwIiQLfc9Q+1xXFfBR7K9zYmUVwuFlub2F1k9qXz
NfOsJ67GaX02HYmxI2fIZuz42vUL8pcPchUNTlTRu/zDESMo2b9SCmIDggEh4Yx3
E+qo7WyHe0E/WkVyIKfoex6uhtFEhoa2I5qphDa6ENNAiCBm49zb8sTLEaJDfZ3i
YJOlqlVsnHzo2zY7mxclo169RoP+JE20NtF8HlTI+SypWFtRB2uGO1L54YJ0KT6q
qgSVM4el0QR3jJdreS79ujUTHqOX4IQ29kubh0ixeruA1kjqp3a5+6k4/BcjUYXM
CM3Twb7MISWkdfGEsBC26o5LAYnillOXcd6tEVIJmYH4XGJB4ED2Cw7yaAmjWV0k
pvi6YWakGSmN1ule+jQztbJQ07mNjNZgfwKvUkzyrC7KxVkenpsWt/3WYgrqBDNU
PBCnuAX5sqMfopkdzhYZ1zlu5BaPD3K0xedaiBbkGdH4+xE8v4kfAQfEdG4Vd123
fW10v7+7RKeO8+54aizB1R0Uakk/1K9hZTYf6Hfubqjx7SoubbwiLu3IqoQa3S7B
jlDRR1TLgwKfJP4Kp0YYbvipIBhP5jAYPFt76D1MHKUrhnlK+MoxSeLNOj3760Ma
I6tpzNb7s2tPIR4qGlM0TOj8b4cOK4h4CJNXueqU8bWicH3zmLbdAcFHgYMk/hie
4U+xUtsBJYlTRIFF8qlVqOdzakh+RAoL22Oo4xgJejpkQL3wSloF/iT635m68yPS
y0lN1hEV+ujSS5Kw0ZxqHRHRfj9YyLypqU+EYIdspnFMtN7dlq8H+JTDSgJ4i+gO
bWUVDIoG5suAcygrxISbxkHYd7C+C1lWBLeFa0dZrW+VQ9NDZ65x5EcnjOU7uUKD
OENaemyNcvCrbQiV7n5ojXMOPH6GiRK060wcQEx2MAuCTZDAY9JrrIZVldLjemHh
ooIreQchiY1Z0uEKJX6fy86GPQrpEEjPShcYb2qc8Ydwfqvj0i/LYD2aCSIEgClr
a5fRMiPXYuXIMINj7aDAY78bghgzYmV1CQ6mSKjdPzNVKsiGAfkl6V3FkEXcS+J8
T5aWoYyTXcrhsiZRRaicZdJC6xNPzCOena8h1C8SuXli50/P/KdSU66EeLLPUYsK
muZwsluJIkRlymzzo0oLXoOfP6IRK4YAS05NxhZjtUeYbjAwqvcXaw/ZXDtPmUwn
bAkb/PIXEMk7sLAz4EG4sPJDQyWTFuCRFjmeHZXjsGiqYc517jxc2y6ARJVK8iog
ZryNjs14Fdv1J389nKZtxao4urL9Go2i2aI/OKbuS4aBfZcwk5FWrawdKU9VRXpq
3gG6IO0EKJ6Lda/CBjT5Uwt+rGa9TnawEmN17FutwVC5hBWo2YgBC2I8FfzVeTVI
RW4OHn6H3oDopU5dNzKb5j3HlFwW113L5kehj3pV/LUmFhfV4uAafjXWFnHN2Wnm
51YQ5hloTsSvXcwpYfuso9C4QkgtiBdeNYfn1ZcDoU3SoYmhpa91cUoXEAeJBOGk
0g7buyguI+GqdZRD0q9kaKDLF1IoU/MgjKI0OevoyeCUKOMyMsQCTk6l+p1fCrto
oxjH/baLQE8jZ054osP3nytCpfE8OYBKFb/+zvTOUW3KOr/D44JoZcSs8J65Tyc6
3GUaj3JYqmOf9XE6V3eW7go1ii2NCBP+PJPnD7NCbF/RXSgH2RdV6Sf4NFAwulnJ
VSOHJFKnf80UZjLm5bzuf3kzmX9j7wQEHdtaGy79YPdtESNVrXBqmtSMknncWtJH
eHWfnHCCjDcliQKY03vBEt2jC7zIHvv6sPQQqZmpm0GSGnnkYb9FlZQJ/PZL/nIt
Yh9W3VOdBJUrBfMkn9gwAY+zec0xtf2dwRH7C1iEuKp5LH0xXb0Z02iG9IPNIhT1
+wJfPg1FU2leJf+pcALYmlk1xg7PZ8oIQIZ48wfHcmovA6ZhlCyHfW67kdy1bqeF
BlQn1U2L80J9dbFA+S7vnQflHqwA7oTJmxvcILMKqFr6cFl7Vf7I1Td9uTJ4mWc1
aAAsJ9WCxEgAXDGvWBiFum9qNI7QZzqUjpSmO4NT+7hgC1AS63K1k6/czPDJRn2S
j88d5qrFlaiibHiFC9Ji1bjU2U90tTPtrGPEBvPggd0oopxzdnqUb9eezE9oanEr
3ibM8krcxDGBpRZJ7mTWFCfiX5z/dgZSBVCh7TqiLW1pcn2khy4kfF5/QilKWT7M
snSvL/CQjPoWROGXbhyfZqCT2QFsd3TKv1ZnTkkm9L5HODfWqd9mU3bMX1ECY7TH
XFTPSNz5GNy1eBjs3BerxzHUY6QI39kK9xgkj0j+vYFjY2VdLs9PNqtRlD/YxacB
5O0TQHS0+U08/esOtSWU+r/qmJklB5OxDAQX/lTtuyjARYK4mj1e7Xr4nwtDyvIe
Qs7vkmyAhftXoq599246SJhBKhT/jeE1yA/WHwI1+/KNIWRXD3n3UOyC5uv6z61G
c9qw9JdHWr9wELv+mY+wpiwFA8RBFEyXWQtA68k+mGqDyxCifHKnukKmIc9/jA1x
PwP99RfNyjlgtPa0vtshVRrGzb8n3MD/hGyXhrnEEVLH+FzU8BTXrrBUhbmgRwb6
VyvNYqrNL+mpwWoy02Dxn7ysNcR5bWNXQRG791gcIlhPvTMfyR9WK4dVk4F+/szU
bm4CAK8g/7+sARM+w2Ss7q0amXFb82dnGPAYDWeFEcLr0at5c/pNA4VT0GWkqsax
8i6Rut4qH/Xe+nyV2GeB6Ka2jc60zB0ogh9iqTbYrIqUKRYv99HsNnGtWMJqkaat
E7OUyk3gWUPagPSF7lb2lV6Qlo0RTNxQnzHiB3z1GzIdYbteKWvqNqm4yU/NQYUv
iY/U2NJRY1bILqLgq5w+EmWZem2j1quBVhJDTTCp42FFV2WHcn5oQ4dIG/t9luKa
+NIsadVq76v5YwdR681NKyKv/sNGPf+PlskJPQkCO8BO6BdQhKjutqBG5J4KVJYv
IOrK3p/R8u+T+TOh2u0LegAKzs9k6EBmKy0gNvExs+Fybwx34dCWwYfrHmh5NF4w
4ZmRgkYbOSzlnhrZP4ofXh1LrcGzbn0OI0X6LLRZq1+rCu+i2v94dpe2y8EOAjrX
So+X0CvBmEVj6wy8GPyjbQXERSuNIXQI47SWkcNsTgCqaP2WHPS0UMj2TVH9fNKw
RZduptk8vfmo0egQOcsLjCxX9vTBDVjnaEmaGEJQeu4sk2ojt1FYDNiqwblPAMx3
r5hXUd+vIDNDN4xa36AcjkTjrgRLHKx2kccxRmZ9ipVbmOwE/HsPtda83+uU9MAG
93zpuLtGbij0gaQ0PE3DeJed1daFLN9RhZE4cLQIL5lhCtGO7nSRETmswW+QT8bh
rIQus9uf3H4R+xum5H147bAtrJtBpd7SlqZGNbs8rCemz3ikVjZT2zj5jKTeLnwJ
ROQvoLuVVAoYd/MNcGUAq27QeI7ONpKmmLsSJ+D3hUHno/m+iv+k9wJX4BXYAkBZ
NVGamn6kw2AdBQy+nH3/siY5dhwFiF9ClQ+dTObGG7ScC+4yIgmOu4pt5o8k2B4j
YZa7qr0WUFJbBisQgwCRKyTDrXW7izVOKrCmRHVQ8isN5TJBM6emYIKVyWnX62i/
fapZsWVqeKaqRTXkGyxiVc4FbTEn+3bq7imA+U9ApMhyXZmwRVsF1B7wODwQS7CW
3DzHHdn+qZbrC0WinKB+U99s10la7Aomy2VU5XLu0ANklx5+8xzQW+JuuNUatOSg
ISsKGRcX+ufgVif+Cu5BlCp6FlgTlkNKWHU12LPwr9n3N3ARk0PagH7XVZSZr6To
ZPYBNFN3x2rMEsWuSR+AbXv43fE/yIr9W5K3eyKZs2X50O68EBvrNI1iD1tKoeE3
t2G9iQqko9rzDfdVPHy6Lw4kXG1mfGBIVCqfMtkCEcu/JiUY5jhPYwI/ja3HIvek
cXo3UPBYPxaAuyWWjxpZlYsq56So2e+3APkX8i0l6xqODMNhmYefU3UUwyX9xsWH
/y35UpDzV3MDwYGCpKWTB8G55EUnRCVugha0+n+3tConfUumg1/K1hWAZGq9rwEu
TFL7gv/6wHn0osoCjs69dMDmVan5t8mqmTr5RR74bNgDFVLSoJnKWWKHuhT2TACG
ZfmD41UIOzbsnM9lFNqKpWQ8N6HfTtDzbE33FSoBtbrHc5RDjCC5F0iv0YyoM/qK
VD8WixkBLaPuvUn7i7iIuFd6RWP5726hij+O6dZ//AG6+FesbQV+J4KrXWfdTsio
2620XHl/qVJGYKCaSY2e4NqzipiWLVQ4ycMxbeeocZ5EYOs0tj+/NFG2VoV6VR3E
HRiV7EwqsUWIR1TbA7sUV++RHuRpApFQkA8q+O2PLjBNM8MJva2229BEkzwo89+N
BeqEvlUvJP4HKZ1zTarsxMxbXFMjV86i/iXIRGRzFwMGmgW7D95nEbFr4Q92EkT+
7mtHEwbx9Zz+n3tMonx0nArp66u+NIiYBiVkVWg4xM1yPRskYlsLlLfts4Bf3fsJ
SZT2vo1rPIVEc6icuQicuQydMMdp3T10dvyorxpVDk/qHro9bxnplHeFt8yodZ/8
3/rzlQF//t/fU767RuVJerjYIaktO05VreOwI3E2R1kIYhHZPVbueHnSvlVvuZb0
FWrgO1lMaysiczHsM2EYstQKrA3jdGE/Er6+Q/XXPqEwqGVycH/b5V7U1uLztA4f
xdwJF4I//iHfGUEybPxudC1LkSEnX6oM1h4yX0fdCUBgwvIKaw+jaZC4+ndoW8k+
ZJuCRfPXBpLrB+cyvhtOil9tfwg/0/fCBLEAxwyaLW3jydG2JVU0fYRzEUkF6ZVq
fxTDqrQooTcTcGXVFAigJQJMD0NIeYw+hfVcQ9d1XgUGGoewDR/EyUE3R4I6BSMm
3VdX0BWUbFVBjwB62oBRVj1Wpkiegaq1h7hFTueE1fGaobt+4i7KjLstLAqRDNHp
1tmPVeSnIWxaNDkoXYnda6b8M3nXWv9227wuly1GgjpC21FLh3gCJtf2GQ5ZosFH
W4flvUdkoS9RuReIcFqag3GWuIqgvJhDrQltAsJ2XHKWnNf6viUwEbY7bM0heWik
IGC6a6//UvNcU/RV4hnbdVSCJjs3iYwnARJTVNJYRNjU05fJ4pU0/skttko1bDr/
TK1cSbiq0Ksd19FACufZZvaYsAOFp8GKShtYeqCb2pO9h3j5At4dHt8WXFS87Ud8
VfTe27SwYeXSG4vp/gu1iyaaXcjAmIC0jw/n1qNyKB7QXdVwZfp54rMM9B1cl194
uabOkxtyQXJoLy5SGQg3gIsyzFMaGMS66ssbEhTbJDhqy/lcZMVfDltIm4XMtGWM
Nln6IlT+gvoIwrvasC9V39vhTrtckJfNJZMnBvzAx+KnlglcYpWeUhI5VjWu0q+y
bsgB5hSPmDzmJDmrmMCSyLB86GZ0wb6SimWAF/8kehKg5774H6rikcFdOMwJ7T+M
XO7WkvlB3H5aaBUJt/nshmurXmObjCI/oC09DNN6JdxQPkqIWKwVKqjwCwp4IMYd
5F9YXInk+1DsI/uUvHY2zVAQ7QBjPUkG5YazCR9zpoHqWC/WocKyLG8gQTK1lo0W
OrB9nwvEFU5uipp7t+Jqh78TKs3uI+EIO68je4vhdAvAq0SvX+sAPILmxUa0UBBp
6U+Idm9fnHHFb2ESneTyG+UJEKMV0XKeasycr3n0f6satPYJ2X7WE2gTzPrPU/Aj
JWFmVHTsFjElkZLRwcdRSAzmK3A5QAa5B0aA8nlV8GTNheML3ve7DOjd+syQY1MP
BJeB6bDXb+SPi56XhMAhG9APG4hgjnVscZZdak0SGmc/AjhlQbsAoVqn6YFzKTE/
EtVgqhB//o/5yWq+iu4N8f9EMh5E5eDyAr7UWlFT3pzR8Sdbmk7MoQ7p2AtyyHSP
dfGPadMW+YD/9odvrc6Ir4x2CeZ5vlAF7/Zz1/N9tjGZz1UX3KxTHLmSdlWRbwwD
KN1vCecBuFBrtrsZGAU1K1XZmZ59W6WCDWcA9tdxYy3DMnvKFDvWItrDXbkC0SCO
6Z5GRlWv/ZEgtcb7ORpSo5TqyF/A1GvIxBqQ+zZfzdaL98/LwySWWukmWg1jJXPf
LbEm582O/jY1g7p/batFpv6wGPmk3z139UXYDLBbp/3OmTw/QBTVtuDxpLNPl4Yj
2XwaZCqegzw08Z9Uk7Sg0+2tAwH2CM4Gm406CPK+C5zkGc8xIQwI4SdNlCtDqXIo
qdBWt0AzkOroQFypGYhyQIgFMQSoy5ZR5fS3nuMMLwVxcSqy0iJoeKCEGCyYhcca
ur+lgOu6EZ9kK4CC8bNjm7OlpWiW/O9Ee363W55rbs9sodur6wQ1/k7jAROMXC4A
i7JpRGWi9tCm69DOcovzAgAw6BLx6mI2oDjDgvytrLGT2xkXmbd4t/q7zIMBdGVw
/9c0JfZ1o+mriPF5bmSaYLTeSpjOOpwPafu9iJfwj7AHZct87JN3u4vHPRq2LT1E
Ecp9IocuBx/kZFlEjOjdnSUacUPhRK+VfEja3BljfHt+5CD9jdNwDE5qMXBrtWq2
wBsVyjJBDMHtA0VMyhu4ADq7lFPdwFazH3zV30mqLK2n9vGOOveMknxxt4IcgtU2
LXdEC032vIN2RfU5CMzFcuoUvi3REf2AOs/geH4bHPmYPWBlK+kHjmtzgonQtqjy
9xLNcGabpdiCErgEncsAo8T1aFWKj6tDtAvGhZNhewc1YhheOb3ky68LX902pIsS
UleBXVIY3TcwfpMJeJsRDDZxnOOAK9PwpvLqTpjAKmrpbkgGgf7IYfQTmioKFjkB
gZ85OutnXAsOD0RSaTmYdbVkYX3v+PD9tOSCnxhuDSVW453V4kwgZme4jb6EQQ3D
7A9JCoMsHm76sJCmFB6CT4kkThkv6Wx82e606XNfClEYr+ZpXzepC9zGA+il/rRw
0cIqVOOZRquyBfIGB6d1G5a5pIhY9bbuhajrC2WnD9ZUdVLFzAiPRymZNhlRP+LZ
YBuUTwgt8vgrxJqt8lSlB8k9yrOX4jYD9Cq0muyBxA9goNskVXYqY3NeTxc+Iy7y
c2AJKDrqfucznBTVxvXzN33WS/obijXJY7Aqm+gUGqWgOpo3Rx0++rJef4pX1wE3
kW/y4iXwspsESo0sRtgmLe3i8mmofNm01faZ6lDGIoQVpROdkog1EuUEOtkRYglH
ShZvALjbIhNhQ3CYLcesBBfwfeqhQUJaS0n70OxSeD9NFpcMUD2Eh+iI2osNbgfW
4s9HH1uWUqI2icNNaNq17f5ha/M3iTN8yKxyO4wrp0WPdHDCGnrO4x4Bg6bJFHD2
Mb6WzQu6X1mm900yBI8y/7LYAl+jdJrJLkpkchny1SNf0EhlI9GOaeOiffzDssvW
d2UhyzW9oF/Q1ke7ZhfnXcffaGvoiZT1aYMRrHuRshqRZ9btUbe1uwS2IpKuA9cw
oVPLSqLqACK/+EXpCa9jz7re+82iw8dFnje9hkJk/BnUSZ97/3/40fLaNaUHLBhX
f6nYWnDSE3dIwyBlWb1UHTFCw70NAQ0eI2wfr/f3J/LuctAn+NVnwFQwqxL3vYoy
GyxGBLvKcvXG25yKJ358R9w1nbTo/gijpItdjfqBMHZ71m+5hdkz2r3/u693Y4R5
s9m/ReuMF9PSf+K3rgVCbqs7v0C18hJZmqPT6PmKAfdMIB2e3Jh9QGL9TctYnhMc
gBV1dqn4V1NIXEOdHXySEpGI8iPuNXMjquEsub0N24qj2FMC9IXr2krGjQizgTYP
a9trIAQ+RdY9gVv5TQI5dHn8HoxC5HAPWQYda4EbzErJRMVpdI6ks3+mtFzfei7V
tOTmelobVKbLnF3B5JQmSN0A/GW+O8KurLehym63Q056N/mfqqv6hsr0hfgTYnEb
5Yfypg2YHi5y74OuZgw87N14dD5rZ9tv6ojIjsj3M2yNeIAe1SFwUNpz3GKly/8g
VnBzzeA6Q0qpB5wpLgyTNiSelHISsIbH9ztEF44cBrrnOOVLsDjMiR9O49y4bvJz
PfSPRU46z8gwzlgNb5M0hfehdBAmwvbzy7VTPYEaK1+sT6aEG3pQDwoRMYTGEsSI
RERk4QBYnfZRjELo4W5dKmAwaxH8vrhzUDRx+sEeHqG0zvX2OoF3e7Ui0DpKz7lW
24JjNCnSMvEQta9Zeu2zj1y6FMjwrK641nOPpokLzyRpH04nzkdKwU9GxEstGeQr
uKeJgJVLXybQm5jvpLx0Ou3WgaEyO+M5yQRAbqxqznr7UckWOaq9UqkYTl4FBOTQ
0Jc78CNuVkgmJRgRhUDIHoKijjEXbQyB94UchHwqx/yGI5b+KDwFjSEm1WKcDCsT
zv7J0LCKAYnptYLcyyASctuMP5HM59k4WxoOh9VQAgxYw1xfru/fgiP7+zsT6QFy
6WvhnjuVPiuoYpgrhRyy5g/W8Yv1S+AObSSphzpheieIF+1JahVvcTYMo7T61jJz
Q4zp0lxm4TLGFBLP9mFXFFIiwhavZ3FznaRswVaGVL/6o7Q64oHwDV88L1OyVrOT
XpZVaq+iIGGRphmDVkkGG9AMIef9Tc1HbAMg93ny+jJVf0JE1uCzKDgO9twZUusZ
+9pVm9V4XgtbXowzWMjPQfOkS5joGQok0uznHZUSLdkt9bycKWchQaslQmeCSHWc
JXOzbJPZDpbZo52IijM4BSItQ31wqQjiLx6TMEzVno1j0rAabDa9/MQtGyXozGRQ
h41rbtmoNv96tT12a+Y4s70wKF5O/5pL0ckJhtNkG9ZSfENzbEoJQ16QPBwiVbtg
wbKHhYG4VMKwAUjw0wXGIXTZ8FkOy+IiYGN4Mz2a2OHIcYl1q/rVZ3Wl63mh9I0S
4BpFZfwjnhdOoIJP0Cl4JD9aUEN2Dq500kYMnQbAVYF/ZpdoD/UrAUq+HTA8puyR
9pAj+/dTIxdZo/gf5HesWsTiby7KZy7Vt5N7nku7h2HaUdrEWzCJJXrgir3jDOJt
4Ad/DANRI7CzQE1kGj5j2nYNrKFa6LwOapgBgJkT+HUvBkzX5WsszI1BcIjkETNl
bSXPgngsV3ggsPDcD3Okra9WXM+kl0sAPecMyQYwaqWnturI3DPP+ZqsHRzNTPSx
qZHqODFJfbHSWnL2ccujMWxX2zQpa/tbgvM7KC1JofFMeHeQFyaLlvq0HfSHzrpF
3zimrMHKg0Ow7i2VlzgeDi5y4eSbLamlXy/QFPK50KOgDYdO3wBi9d8zkxk3VYTq
orMUitoqujGEKsH5erjIvYBIeBdC3yWryvoLw4NA8yoCp7dvJNm0bow43pxH2SFU
EzFqG4nU4aXtvZDsOefs+q0TT8wnwgoXoTzkcMJpWwUNOrZBxTzwTbvd1+mjMVgq
MrZdMbJqbndr3J5xMvvekJk3difI6gqrmAxb2Rl4cQS9giYPmUS5aAq5azfFx9Q3
YRpHo5C2h9pX9ChlEPhdG7cauZtJtjqWMeYFwwW7oEEy30o7IDqCrqXf0Hnsi4mh
RJPYdz1cRvGm78QYXKV1aVJzEzFwhg7+GXlmCcpDGuN0B2uW7ujaj3kPHmW2zsDm
OPb0GhG/6nhwX+AeZKWHubva+wTY28x42maJHTa+knyk90AHOVI26JRFctcAEICu
L18fJBe5kAMbOMJ80ntPKWWcYfzLVgJ2uJaGpKRbj5dVlR1yaJozgtL46TcPMXlq
wmnmr3t9vrM3CubVA8tft+PpYzhfVyiAABkaBz4vlqIxNvV89/iCQI/mhreElGv6
7ykHGVtkOgEqhpmXARRca8w2hV7+wXzidI/1oHUH5+jv8FrErZzGkC6LrahNf8ri
xHvxS6XcrJEV4of27HKykjM+sOA7HM+UyeJBwz2dpvyuw4H5ZwOdmhp3dyBFgfhd
tSdFOxo3BgGnd/Vt7uO1ZFuptO+G9T2S7JV1pBk9QfHiZ9UWvU6l9160D8562VlJ
ug4a+Wrf/i3vD3swXmBNkR9Jq4z7UtZPFq5lzb2KoOhMvF8tUrCvpt0Mh6EwrvTf
oIilVwfRSK/30xMVUjBzTdRAE9GrRirMZ47a6+vuHVs3bE+X4hNYej6tl3ZlaRlc
YNiRULQhp0ZlIPlvZ/ZDliuaZNOea28ZNWbCPxBc+uKIUbI9+FLS31/Vq7TugNRK
gYPFC7POQTjwBJxpszDC/RXLZV5jxaL6BYyl+YQxg1XIkCb0+++x1hirlrbvzU8G
yx0xoBY5xyJ2zp8m0SoVU8AXPqWBp8u0Iy9T2jAZqTsq1RSE/f1TLKdtEwcyM8bz
FQSvbg2wFW3SOOK5NOGay/eiGDsptSZ6v/DgSBnTs8WA1W9WaK0b5h/UY/5jVw4V
sZrfyCg1oZb/QhNa99O0DxetiE78ReFOKYFrqC2A0jjwvUfs4IQFkzaVxgjO4JmY
rMhEAuZILcPvQXxPf7hq9Hue46ioeT3TIUjMVCuzRU1Y5+PqfGek4scuI0GP2r3e
PTREYBlDGRa2NENlG/45lkCTkwVmk6VZKMxgDAWS/ZA5TVjXZUOS2EBTS6Z8YYEK
Xl69kfl+xhN654XCFULkl1QOxJ2+heJhERtXL9CnpMYbXJ5x41n4sllGPWbceqH6
QRpAHLR1t5AHPCsGxcgNbuMemcSw5psTa2+ZgWXXoVCmLs7bTuZ9irYIecLY3rlR
NSxWB7M3XXFBJPxvk+bFim+ZcPL/eD4Vi7kt+u9XXdWUwlMGiRzeO9ggWVdmzqO9
210QXfo/wKjG0ia4h7V9dmpUT7Qu+HS1+ZgzMw/aQ5ZuYd/AL8lWzUn/ahR2I90H
KM+xpFd1+pa1XnliYZssWej6gEV09pwxdsei/AaFtSwDvJ3fl1xlt4w0k4JMGJBy
+sRmaojxlpot6NClRv9pI8ddPC/5MYjTd/GI4X1/qupYytVjTIECEEDfBAAa3eV+
9Z5bDJREccJLQ+p5Bp4BkHN1k4Jm6x12Tr1bE9dKRqo5HbWqnealv6gk1dMNYUNX
TaFssyEwZmbERFsqfPLSZ6bUAThvL47fL8Qo1WHVCj7usi2NyUAsDyyB1shZSYeG
QWIC8dwPEZg9i3LqAgVpUA7JRii6acXhUotlEWY/aE1Q+h23wKoWEO0Yna6aqdl4
tJGf48FFkkReUtGd//vgQTJ/0yfJVIinTKLEgWIqcrJt9nUYqYogYqQDQZF7uibd
sfpKmhYOfBnbv64eUcP6U2n9unKjISZ8pov7Sy7egCVBecaO6L8d/Q4PLF4q5D7/
aY7Cq0PkqPt9Yu3GoiXL5MYzdr/8U2D80GeKYzJoGlbzFXnP4EppYgF+gFnRqx+v
yR5a0O87ppEsxBsiHLQhW9W5fHBsESqjKxIMcYlVsJ28JUk5hscxpPVyr1S5tMaG
OEFw9pGFtvYYszOrE1NLLnvYXby/57x85CKXMdPm+IJIwZ4yFhDc5gI9+p1UJs6Q
T7eTEbi2Y5jX/1wlTHtWGlWgIEJZ8wKHQkVOVr9Y2rla4CychhLyItTVbQRDCICR
cOBejEIEkvxILbQ7qfRh7KuH3OS9lIO+yYUKhobJy5tztAJmQOT/2cpvjqaPDA8S
YnEHyMaBCcRwMtBA+qiNKdyqkiefWAMnt7+KXONdRfIrxS421HP4xnBfVVFgPXK2
+clDLzh3fZJY1FsPctuQHCPcBAaKqtZQgknOE+Ccz3s2AQMED+ltltLiGO0B2+dC
LHvi6VeKqAt2o8vmvQUPfxf5Tf+32iKTxzj2Mc6rFkfFwhrWuCpNhth7RFZ11sBB
lA6IEUYtDqxvMiFEHdP/h5cmnLhZRRT0O74bKG8L5sZutuKXKCGM4+R+z588xQLj
wjPfctbRqaEXeeB47I4MqwRpCkLlLjorJb8Vao5glAN/tgEe6prBeio/y/1uVRJz
JmeR4c2urlUQt8rQjBL4YdVj4Zt7m8cDnXIMC58JPvfnzqDsnLi3ROM0of+SOQld
J+cUk9pTEkovLrE5tdlzL5OX8dZm3AllO4LU4kA6nEL5uhH40FkJHTCe3ZzrBl+o
k7yXSL53Qxu1bLFwPKqXzJG4z67chxzNZoxMc/pX1bZCWWUoqNkFgml7cxduoDJw
p0i7o3y5BXZyquw0I4f5NhJmz5O0pjfcuGpOprLgApur1cTXaf+xAzegt4XHRQLL
j0NA6GD6Ry1zRTrmxXlt244I3nBKSnzsIEAVFK6C9EuSVJkizLY9/yTa/4X+T2cL
uCmx+w3a40nexMIXMZ/ZHaMtZVYMmJyx0dd43ktRZ1Tvud67/pK5LFAhjEL1oXfE
XxBtwzaf5Gsa8wSjY/6KPFm74pnY6BknSrZLgCefMXTGMOFHEBa2QnWEpa+Fg+x8
+Xi+Qc+c5AmHoubCeWqix9VEKPsaCPc8yPgEIQmkaj62cpL+Mfl7BKdqU8ygO8FW
S/lr/i0emGCO4mmcqgRVlUjYvYytA1qNsP/woPfOn4lYgtjysSWkagDQLb4rHihI
gd1R7lz2GJu7yDwtYT39VJf1APWPr43w8nwq1gG4eEJNrsxziKcBL4F86KBTIbbb
meWJ0b5H66ichZlNNReG16AOYL6Amb7m/WAHmLtutnnSP9AlRmcxHHAdKrlKZZhY
Ud8BfeKHt99+WxCotq0wCk70s/4kv5NyeP2nYoiktmmKpzZ7EX4ldsgRRDzGbR3I
BOsg06mcwhl4q68KyVt/T7tjsKZTe7ii/uihwyFTWvm+nlJHiZmi7etOi829HR4p
kZzDnq4/TTpdD9vpaakjdAAGn/7vFHbs/v2XOgp4utIkcwhisUEUbBpbeoozPJ0i
Ke4MdBDn7dH9LxNI4gYpOrFdqLnuwdrwkKZHdjA5ml6a6CJI0mlSE0hdIZMF1D7t
inks9Zqejb/qim+tz5XilAZLlJjYYTOaYj/rPZHfj2fGzRWQhsFqdsyKloZoYoNY
XEsNvC2a+Aw7U1pSJ/f9v90X0oosRuq36WNdv0pydpJGp6kaaCcktG6gsVa1u8Tb
QjGZa3c3abN101hZwRscIZxQbSDxYTPWlY5sY2UxyVriMkLce4/HWPN1F6NFLpJx
IIxVkA110qiPtD2fN9R6E05dE8MJTW1SSsiBuuhckk5weVtBEKjEtxLEVqTF4v3P
vC3luIWMxLDz7IVTpwWCsVGnWnGfp8OxjXJ2K4rhPaMXSHfLpCTXFWlgX1JfEVgh
8MXZpObIACuCeX3obg1fzWK8katNnK/pDVR05Lb8g0gEAqKmFellCNJy6hR7fvYJ
fPbD3FbOsoyBNDAqgIzsJ78aw+lX0wql6tJMJRPzv/IKHq2i1zgNAk236yTapwrG
jQrY7lS2xLDAgeEZXiwLmv43xZURRnZTQOPRrz3sYFwGKeCfygUl6bx4W21sARfj
23NmNiRUIgCbUq+oKnAw1WILGSyM4FGvjyrYuViptydJ5KQ/v7sSn48u4rYua40e
t5izPRkMtbYliRHY/5vOtBOyIpwzm+K8JDhHM6Kv+6zky1VRT6ckvf8Qz6MWdy7Q
gH919tAMKMQMg45TN8x/4wFpJqfGNJlc9JY31SZL4LEaOeqPgPKN3VdkDe36AtmV
TUlLZieT3ooqUh8lKCiLH41sEwvLQlCws6ZKTZvbk3l9TkJqjiJPs/6Q0uVIp49L
GPiE3jHquuWrVYEGrQQu4PI2izWyXwW3NzKkS+kmK6fP1BuBJ3J1sht86J5FUWzQ
QVi5rpaDa9bOEh2U68Ca8YI/vBqshT+0DYWDeRrxRJ0/e2IsALzhZ3HH/NWxfkIR
qGcj1spuxkFFja0WZhlFD7HYfbbaPExSHWMhbkS4A4EE12p3JhcLMswbAbazGDSq
UrQVd5TRfGFSxkUR3H94SZUY2bAQR8W21EEKUtana65TxoHSn3GLFoAmmanfSDEC
4B2f3i5ofUN0pEFTNbmt6n2xnhYF7+bHCCG6FRpnlXrf4bWUATMe70QvcOSziNQ7
KzKOf54szdw4KBS41Um4pVMVRzHhp/GPih5oExy7WpSdSHS/iWcsBlPu1IrLBQ+h
cXnwPNeAw4uYVvy0U3TRuPHinckP3BPBBLA/nvfUwe2VTZ3beImPeJUFRmFjcZao
KbWpft7MkOwhz77mpPft2c+Y53BPMlNsybfbAwQ/Og9M1rwn40Hi0BLYcIaCIYW5
4aDW966G/FlOE54l+o3JyF1mFc7g1RM1xITN42SKXI21j44gpD0/dv05K3tcvpGo
vRqK3o9MuB3r3hWVGJx0PTQJql1NszzscTHWv22Yaht832bh22Cqjc3LMakZRXth
EqgokGqiO+JzhO+Fg7rehrx+XMn+tU7E0SL+47cUYzDzuTtuH9NjeaQ7F7YLaivJ
zy5iY7CViOpRFJ+8cj01nHEJEi9GdCGDxfehFIIoEV+C9cfJ+6SaCrFxA4Yz4WTg
AVVGsklHxNWcunk2igp3wZU7+8TnE8LHORrSVAa8isLkPCYgcNOHYzglxyxGLbzK
KjCpBVFZ1faufzwV6AdvfhNvwdLXaDZdtCOKmCrb9IcLfRkM2Ryp0NeHvuWh8+yy
ULu/AqyCBvJby8BvCkY25XZ3BHqjoWKUkDclX6aIitD26W74HBNaEUiPNcy8gRjL
ba/zNH0I3tR51z7ZWq84l9n1yL09Y8/shXqmRwV7D2g7u/vouHPel1KOzhXamqB5
ELx572KciO1TG6/6DDu7TbayLLuQC+87IpW8jvTTlNoX4waB4wAyiXDqPQL+zAP9
HVmpfl7uPUtJ9iYyy6jXocOY3j0/8WYe3BrEdYdvgC5W0TBQe4ytv1K8tFz+bKYR
ZsgeSVcvmHzp8Ey6z//fkEHdYFjeCPtZxDgOfxNbcq5bSbnR0k7gv6z82p/sBU1D
lB8im5NHap9lcZ4CjtKK5ZxGClbG3qctEdFZccVomLrkvqy6VCJxSzQS2YltDfG9
Jx1TCSEZDV7Kns1FGTIQLBarvS563xxv+zYN4ONc9WkqWWVRvox9C+DqVqLaFFX9
Q3tuTyeMJVqbrVWuzpF4s8DlZE2YEOOO4mziDJbwQMOSvNGN3hm4uU+hhGHIaVSh
GLR0vYpX6M5mWVnGhQA/AbTehyXbF6rbUaEuhoEfykgye9VKK6wTmlw+8ho7Gycu
LadQsPMSHV0x4jnaz3pnynyKp3KciHcPdgTH5tGU4RwNoi8KAJRbcSoFhgvBCWEx
+r+HimmUhI6051hktU4NoCybyHaUTrBYA9QJpsIY+ad1cb+fHTgHBsJ7SpTkW1BC
T/o8wUZEWoQi36nEZniHgb0rQTpfebVRdL3Blwj+f+ixuuLWQcxF/Fa6vc/i63NY
9btTVw9XEWUbNNbvh+BrzW75pMP+lO4McGSBcjnM1eXIkvwo1Q8tU53iZ5q3Idoo
0ZgozCM8hkg2Xn6lta2HmsUF5/k5yElXQH9nse5+/brbBQnRczmcvNLQEoVS3hCo
SRTYUaXzFqI8as+aOXvxXHzzHomYu8Q8eMKcSd/Qo8aoTK0sM8PRlDIAVN2gtf5n
rMXQOZUlv75VG+T7VLJCcCr2F54E1UWLa1dJt0476LHlZVYQ4mlxKATWPrNf75nV
iPkKTzlqCPhe7edbcednpMPmzYfHkRwoYLsaCglRWnU64eSkosnfz+Y+q0rdOxQz
60To40zYSOngOq8LEKlStkGBtrhUuLeoHzP/isfRui9lb1Rv+kHegO54dscO5EvN
Rvna8qokxFdV4PI5HSqxOX6EAtvvfHH7nX3FqMp+H5AH6w4tSkCYP27aMIwTF0cl
2/6EkBxMlsEK2XcwDLtu2bLAr4oY9lQcl0qLtWgDl6uFG8rXnu6Ue2ulVOwCGu5y
kUR519PITQV78k8iP/NAqBIOisCyqD8OCVn4hGXWhHxgDgB5KUuw2E6RAvzJCj6g
Ksgldqt3QuROYrWTrD82gMF9ejA43mYy7OLDBQAAH23ElS2wFOSzHGVjEVCL5x5Z
4cVArr8OXmGmUclJek18MH7wc3lyh5XY/YvCFsiVepdm+5ePciRGur7xd5pTOcov
jx3XPN/X9h9s4fZkIBTHHhCtzDTt7js1gw35zb1zhDR/HC+jJPJLJWawqF0QSOmk
+TZN0YWQFQGF+e6xyFVz+++X1m4sIq+hgBkGePzYAA/kqH59JT18KKVQcSv5t4b6
Uq34xC2qo/YJtDDV/04jFestkieiCj5ib6iPdvggWB0M6eyZBWP+24FeU+hgnYtP
oNkwFQB1wzj36dpNGqXKYMr47XhFDkYTusGz3RS1WaiZ+0Uh4+boAUoRVig9PRgV
BUVAyRSEOSligYzhl+ZV0efkZXqRUOhNDr35DsnN37TnX2UADbaSvI1m/ZycgAXg
BMrSl2vyYjQinr/escTbpoRrfYNyYYw7t0GjWGkQxJMCOn1EeWCPKFS4NNN/z8Ye
mA/QuDNM90naHVOs76O8D6Bkn85if4faXQ+bWWf/hWIl/is4/qZQFMEc2zoNyswv
Z6olJ4K/XXPa2SOOjWs9ginJpYwbu1NCpoItGD8E52LCKkcarbhG08PUoGLnz/t+
AWSS/cw996B9j2rbxUKeooAeJBYz9orHCZNCeFuOQ/U5y4+WMALRblqqtDmGpASt
htUQdnlp7EEVTHxjQEcj8RuJK2HDZlEVqRj/XDuHUAzgWfc3PhjEqjbW2nMO5SvX
pcrxa+7mdEKwiL/mDAkFYSvNxIknbXDjxBIGS4VMNrayUi8mCwePvpECKfOcPltq
9dWDSxwpBPpiyTtOKusMWQ2x/BWstIIxLC3Qil6zdHSp5nikH32aSZhhdKDur70K
PCDM3BdmL5nkH7hS7i8Jzi4KyMMe34Ymzh0L9K7ko4T0pRHurymgQh0P6AQdkTSs
vrvt2w4bsFDDlNSBhjorDF9gcNpAQtf6NDUHwHJo7/XtEcoXHnxS3qezV+V+lNR4
4IdLifVKpYp4HGhDzjyq7wWeXn1in3rHrjJhni3tQgL9ToXv48wjjx8+Hc5OS6Zm
BzSZKPg/RIT3WckkDQ7tb2zp/SHIyGD/nrrtx3dGhB0/JfaxY7lyUqNw0uIaMFKJ
uNYM2UTLWMh8DMGC8TogasY/Oi2G8CSylqL/+TtAcVTLo8Ux+fKa1Wv2kmcltQlY
DjLh/+6vHukqk8aRZhbdhUWyBECAnxuQ5xrxjEPXxcnZZx2OlAEBoRBoa0+tYFkU
E5iHCLHR85LHmSsqgnRd+B5jiOhDN4gBNNBH3awrkYAUlXzM5JcoqVLxulCtmar6
harDR/fQRxFnNWM72CmywKbogl/7Ah1o+an77RNRW6GkEXNCqzXPwdx926ZHMnJm
snrTgWiZillT9Ktm1uWutIRkufqzwFe1yD0lx39zUUTE9+5HX9XYn0MqP7P0LksF
puOH4nk0OcvonbKbZQH8WF5nX5hsrnhQi9d+5DZAxMpFo62GuKxY8kh6SrwMMV2h
zfJGyPyliC1QZ90iUodiagL9x5tJTYH2gSre3ENtJSTbFfKw2hgzafOoW/Z519EH
8ODbO76N2EXS6L11Pd6s5Z4xykttVNB1SPt5ILSui/fhZLZv2H8+QFCM1zDz/d2d
3HDNaL05kfQL/r1FwA/gJF3tQi7u6rYCrhSuwaXKx1kHNBIqDt/ebzuGZtUax1Tw
nHwg903yTJjaT+Mq3AcxZevFMOxdprCvfgktKLOOg4Xv2VV47DY1dytbOzeQBdga
+NA+Z+02vgukkRQBBh536rw94g1a7sxGoBo1qo7M1sxo//Y6Q7A5HHn3NSTljozL
fhuWrGAFRqGXrL9FsMlD4udDwAFrelsDl4czY8Sn74KpOjtMWiWWWOTM2ImvNyWB
0VMGtS1mjpRVJ0B1OJ3AkoM6lvZGISnq3Od6hNmKfZY1lUuYVwRHhlADCbFlLYkx
a/IpWOxaKLsHru+J5VQuhSa+FLiJjqPjczQK9/bLeQCd8JngJabWEZr4amppS6Vp
iIELgZoh/D1/FB6CbaNjAX16tbGJBvusWuOPgEI8fw/eu2ggC5VAVgCICu5nEGPM
KdYRwvFAgNmfv5xtjBDarEuisSmcWQ/RzF7gN6lZ73t9vQ5Nt/2+sxEXSZmT7k8M
qRvYowcMYibwmtBAQJvooTbt15s9n6P7S7Xv82Lr8XGe2bLl6W1XUGHYSGYOZPqT
Lqw8BuTOJ677lB/QQF/0YNWowCdBHQWjFHe72UepiDDRb6VV5G3xAio3mEaWSoRO
Pz81vA5k+erLlORXXs84/6SujLNyLcLHylfruLWo6OX9x9TAG1DWi37UYM2z/KC6
argvJJUM97ngRbAOxfGEgv2VeGUCeDpxHKGesmC1dKQ0eKAGKfQLbKkeBp1py9/U
GObshPkWDmlu2nj+8ZqBwl8YC1lUpbcYVjrcDT2zzX+dZE980Qgx06cZgUvEETzT
4cOEq5vWRRBkKqttrnDoJKcTxq+x/cpKzOVnXTchx08dX0YDHMUefmWhgWg4nEyk
Bjtsyr7lyhjmF2t1wJ1vVS4LRaFSt+rBfpA/uVN5YIMtqyzkWhQeU0L1w/9xNXVh
g9HALAUvEir61MO9ZD/3wSzOZSSlj7Y8tScvqTmDSvYyfiWxbp+3UmnXIQe+9r3n
4SrhgjNFrqFhmh+awCx3qiwjmGmmyUhUch7jSGz3iMERX8ZdVjr1BsAbsb/sDoHw
BeodcOAxycKAhC/uU9jhiNCnHyTmzK5LrutUYweUlhZ+ztMDTgLxY92ue3F1Flaj
sZUvxESZJ9k06tl/xKYbzqDx51Ys0ey6siaoSG2l35Zow3lkZ25PlKJNzg0tYI4H
m48U/67CJ6kZNevKXQ+JD2z2edlGXXNj6sfkrkjT1AQ3lSGCFFbGhH844uWtbVSX
aW9lmfVvb+GAENX1q8P4so5+7YB+WS0BAhtwRLwBFUIsmMupoU+vcOAssig26Rhy
if6q6s03145JcCgzjGDb6unn1YXTNGJEAnpX44Px6UqESgg0v+v80+GhAhQl525k
mdU76oafnC4rBUhT3BQAo4bPGf8YaBwFer+f7OGzlZW2lOsRwSOFZe2mvpq2Q2Xe
S5coQAKLHMzWOOnwyuYS1RY0n350dDoUtNkYxgk+IZEWCrpuqRjHxIvgWrM2Vk8a
B40UYRKCmXCAzNVAeKEs8jC2ajhjZc9B8urh3926thNcpdtL52mxKXeO02+HZxcI
RMgbgJCsNWV2s5pqZL3FT0hQYylCFa3H7bWv2V5G0ptxCJRwy3d4XptbywuVJ2eW
6BCNu8x4AQO3fTNxI5o4CY6I13uTRc+6Jf3aZZHFTGDCrV8sKptINq5eSCg18uoV
xKXyixI/mIrRo7v/rLpVEZggL2iJpm02LgXSsfK02OunuuKc4vDVbQnE3eJrl6d3
fzR7EoGAsPQgbIjvits7rzBb+K0c1xtO3mKRyPQ146IyO41KURXZsmUvnL9x527Y
6F/LvZU8QYyn1FqgMOFgtzDWAK4sLPYiSmuSiLh2jCq06yu8KeuBP12+7jVNe6bg
fTil722hynkpKQLhrWt2/eNuyb60I1CEVMhS2cO0WlL7DdUxxp2FVtRbnAhmR2HQ
gst+KNGwifW39JW2qvinuO0Ka3In1af0BeCpH2/U0i5BzCWtA2m8PEECOM8GV2Ml
sFcjEr4MXtk9pt/bEIP+z8lpOgG0yfGvit6DyvrJmGSi7PDNI551Osl1H8S7bHzU
/WB/oegQjXAf/c0+aGOsbbm/nO+JKl5NwnYhegKmI93NjceEqZcNw9OXzTsZBRgC
W4BNESgLRsX2SAUnbRpNfCRCWW/5HS2zhfMK2oRadSjeepcSM3UjJBn/4GZZnvld
SLnxL0Z/TA8vvleZVg4Ty/HJlurRq1DNw64u0/DSLW6SnBk7z3NhvGBku9/Fp70l
46HweRNH8DHRt+O2w8aD2hZPVeq4pQClpawuLSVxVckdt9/d8PuU8GneATDYdDww
+xygR0yRPQIa7c9wMkR6cgDD4hPOIeP54cTTHi+IqSEMi1m3JMX2L2JUUZ685QsL
VnsHR60MHY2sk2DP2VoXtAXYOED4OUAsf3ID2MSDlnYpx4F+e6svh5k8dNwbIrYE
V3oZcPVClJzcxLXSGswlMSCgDtOE0CLAlOkWEKXiYWYd5y/2aylXAlh1+yNtTQFs
kVbFcRyKqupdB9XJgs8mau+pYK497RZjuJNIwS1Bb8BZ9RNlBKGFzfoWZ9yNLKJk
IyC2D8A0KCW0V6ApQHh+CepFau2K89/AhOzWmbs8dNV5pBBOuU8fIk64bhdYiaIp
a4TAZH/AYJ50fzmqH0c7+8GSJx21p5Ai7CgxFTq3YCdOO+vgnnL6lQa4/mdNFzrm
aEyV3mK79X0EVaEzd5HtTcE42iR06h/YZu9BZB9atsq0Siq/ih7wnQK2KrbDauDl
bbRNgvq/CaTW6do12LXTl7QEyyPPMQyeuAqg+wTrsAbAeFmIpOvVe+94MJxjHuoJ
/xUKpDtZB+hSKfUqnirLJY3t1e0zsuD0iVKVS5yfqt4xVeSG4lZ38IdXp+G2vQx4
6WfS2PHVF/qSJiUprfZHpyaQ6LaWvSEdpupIH0ROrE8MC9aBuXqCpKysfa1XMJMs
ipa7fWbLoIyc/p04fz6F62azIpB+Wl4wFLsGYtS0hWlZ1VG3CBcd+kMotJA4ZKMv
7kspInZcdSGdH2hGsyZmNo6xXYq8klto67/+f/EhPUng083YyqPmu2kUSioQy/yT
TvKK2AcBQaS4p+/NS1EJvv4K0KpllWhaWxemwcuICzpPRZQdrEdmDEXtAvwU2V7x
ERLjzdYvdViPbyMPiYQvtL3+RHhNH3jAiGBvIvA4owzb7YQtAC0oiYesi/NPyuT5
528CcD56ldLxBC8cgds7qG7f0PSg/FGEK2WArfayFp4dMUj8FrSxazYEKKcQjN5J
TUHViQf3DzfrImNjoq2IjBT22Rw82nfK66IWOZ11zmwDW+IHJG8rEy1ZZpPwyXUj
n1ZToUujzLymXK3Pdb37kx/p3p+Df3xw4+PC+4CzTJnItfxFuATEWwLmPknHTdEs
WW6OWKXn3Kg1vTIucK1b2+FqBlCX6SkNZ5yp/dqytk/mNYaOEU9F9MacSFFgGO7M
xp9umC0sBQhnQ2O9s8txZ7/1/1N4dr8KpHugzQUAOE77nBlYlK0irTAqRCU7qCWV
RRS+iswjJ5Tf/cnbDkfWFIGYewn/7gytcRaUlDQLU2MBHRBusS9Qxuea5ruYR1jA
sMye+pUOkKzODic6dLp8cUyUJ3qd/9WSOnkgJ1atLACPSXeQDdEleGhm8xeVz3fe
7OaLFCyeDtMbWLiRtGQ01sXuBxSTGa5jqkjvsfHawNe7kSmdEfvH5e56y4WEAz5z
4g2oiJd1Wsf7aTEBAXJ+28dh9gJbbfzJimtaDzEASeGD/Aa7PBs3NJrKnli61d0W
sE4f0/jCLG2aQ+AUacOZKDSqTTesqvWAvsYOuIMKiti+KmsDHEWpUAULNTJzlkfM
u6yPrge0a0OcG9H8wT7cUARz/d76BvyAU2sfBivDE2l/KFjoB5ZKDrk4Q3sYtqZ3
ebMwA5lnbhLONc3kXmf4URelANUxAAykUJj7z5Km6q1UNcDUBzji0GTaxNSEWppT
vP2pnJSLp+LPx2DJcuTmH/RWlMkf9FkaAL45I6JRobaQRp3Ob493nSVw4z/38j5E
tOaFG7LMjEOGUn+CkTl5axMY4lIiU1sUDygPh57G3O7/jktnBs2sKe8TmBBzxJaZ
cTjJtW4cDR6SpP1+tQGA4z6q/j++VS2SRHioka5YM+8/CTF8j4juV40UnbdBzopA
FbFrffrOWJou/V7hAxGHgZSciP1XoLLDEyaT9k93v0qIdjKXAaePY85a4Qh74Kog
lPKiUwXNPNoysdDCUsaG/Am6IPINefaydHx+EgtqLp74LqM2i8rfFzHQppnpWK1j
O/SGB1HFeAYk438i3SQbbQYskNYPY7D4okiVORQiu0+U4ksZ8yuX9Tmyjrw7RCgQ
ZVObwg07rd+o3Fa82ElsLKjkyvWU1uHV7nrRnQh/zEybRGlKHoc9F/QxjEMo4qom
AXxc1rm4Vf+VGcbPKJHap1wBj+P08fHm4UURJpm/fghQMfZlbBkdUrqQpTltbPan
q6E4GOV70UZP9leRzQ22rimWQKRKg7MLbGh88lFz1/NbUqciHvc0JtYpYrahUq/N
2VV5TmY5qF8lXMwA+UZLn8yWzq7yi21K7v2/HO5v0f6W8WuT0TZilGNchlxa3Zs6
M8Ni2QK3EkX88I6jyIwnRY8ZEV0Pl6I8I+E7LqG9uJI9wDj6AWjmG1aqLetTFMaV
Q3WrzKaIgZ2TxE6jnu4D+rmh9lTrGqGj6RHUFUU0xgdzb587/P75lU4wxVFkLMHJ
CsXgy6QH+el4JC9sXYQPUhesue9E6wALNqYRjbiX64awE7U/Ojh0oeoHsTPqXq6X
Zkp9OQO8LuxVe7d3xh63xGloLMeDlNxCrZqighMJYRVdBLNlNurEg3Jwsb++ASM9
lYFXitORzOATT/2oWdxrn+gqiYNFlAZfkLEEnHsl3Ra+X6kmQwaSXSKfOYIksOow
fMZKISiRyicjVOr9CoVQtgU5GGf9iSfTZBksdRrCtJ5jetMCy+qJzASmYGFPU12N
cgIF7KjVKoHav8dbvVpRLlmM2gOGaPgwEseZCpzTMfuJBHQrrYn3RwMb9g3gyokI
qp3uL8GbDxa2cOa+++myShL12aTo0YVql5s/cfgauTg1rKk3ApBXThOzVkgzS5YN
Tn8Kba8SAMCDouhig3vDB7VY0elvTnhiqhcOAbo8qQsIiSt3uhwdg7CUh/9d+U88
aN6MdZxyJiQjjU+VsOLUeelzZUJSa6VMI5+DOgQ7pYvsWXOvyM+Gr0pTT79SAVOm
ltD6orpPal8zg6I2GJQ59D6ETyKM9/cJYoMpEeFTI84BSKcecHOkt0bkQFcVfju2
okcZ4NS1MJocjN2nekbesjQsOzlY99qneIZ3gJ+Zd1jZTLv30RV2CCyfzR00KPpf
7QXOgq0IybrFNVsRfumAFnIHM9Hl4Pu8tEjirm8Vxjhor5Txs4dPM4OPEdiLu2LE
zLOfgZTNbaHB44Qk1a/bpmVlqCOZQtrNLTCMlgErWbPi6/Kzyn1WQ89YA0xalVJ9
fBlA8D9I2FfDglTKudZTCxiDPJveJMTgqjiY/Nyv4BjPE5VGdIu2ak5es17gVtcJ
u8gBtYeQLzeRkgvZYKSZleWb0mae4xdFJzFmH846Yvk6XMBgPMZfXj34DOe8i3n0
O4YIDn52QUkD+GXrf+VcjAxgkwv4DHZYJQLL1yiMkmQIThrSrnwad42svv0A7vVL
StVQU0+4rP4zAUJAmbLwNzECoe7rZKbkt8p7khdR2/mAMyv9tHaVswpwtSwbr9lI
eqzzUhgbUJtVS3oj7gjH90JxajX8SKQJQQQjvfTbBN5oN0vvuuddlXwR8qfwmPv6
TJWT3//lis5jTpnWIIIzYDEIAbhNPoPrWF6KxGSjZwGK83knPj+b2WvUfmZfZJtp
3NS9AWSkxLMiC/2TxaeHntpV6yD1yX+Oqcbe4oWdJ2goapD61Uy6Y3QYMjj/a/Dc
xMB/Jks5pVjJ5iNB4ljQwVqB0z1NeYrIP1gqseZYZ6liKP9vkusqsAeqaYlnORLN
X0if1Wo5Z71RSi8X2er4WCl61jkZP0AueuGWvklyeat1SeGoP2jKBDpoIbKYcT6u
TorDekN3quLpHuCrhriXbUC+K2+5rwr0Ezt9rxeQEql2mAmmgI03qvsgRojHmOuX
lxUAjTPvibLhWRI2qxX3ZPmknA+wJb6kGZ7pl6ojaGDKV32Sv6qEGutZK9YSJLaA
C0seRJ7B+mzEXERr9RCxTGQILX7WoZ/f5o0gN36T6E0g7Y82tWOigJq8Iw76G90a
PX3yiZNRSQ396xNOqTQSfE/5QMSA/TJI3h3BBNJDprjXali3NDO5ynLdvsyYAVKu
sSEOjGEDTMQ4SIjikvwHrl9jE89/4DSC27Mu7tmeEx5j8UtkFZgKrtE3f6RRKID9
HrDuxxC0Htl440iqjLPtvb6KQfTfbZGB+3rKsKFWLgRIgoTkfxvE7PHYezF2HsZA
7y7hxJnlCr3XE4nvYe9J7D9LVYcJOm2o7bgoUvmayVQh8MzYF95rbXqdIq/8OEqd
27cy4rm+bEZwZYW+ngdZ62Lx7/lDw+qvlwQJ/qmqoPU/TAgS4OzgPVg2feKzf3nG
hvtjd7OL5x5HYc6lH9nbaQsif8V3CLB0irf9yGThK1FYuvrpsxo/6kydsqWq6BkO
5JGBv+5vWl0DSVkGIUpOdcd4R55B6bK4SPP7oe9mzBna0B0UM4X/GoaplHbuUBRm
rRTZKeQudb/YejBuWOmcpFntUA5C/RE4HEN9bFwPl7zaOn9J0xRRHXh8Xc/8N8MJ
u/2ivSc8It4xamZZ2vTrdlgp8Jqy8wj0hhoztV9V5Ps1w/GJ/6LASkymOR1vOu7F
RVfs2PlFOfCkGH8dICDYYbVySx3SzQ0kd7gLjlL42xOpNkVFLUYC1JIJIY+hHAqF
XIXHN+wEyAerwEvBi3f2G+9Fpf0JFKcuBV4fL1i4H/KiOcuHCVAgavIPMTMK/pCr
QZtTgOZs/qCMDpzU9JAKNTWqFGnJIDsxt2ULFu6iCiATneEkLYYOsKjaZmWrQVRg
IgqnC2PWAMu6yGPOJ3058VDNiGfD9hiPhASB0eUUXiELqTCfOLhJAu1AkVS9eGT7
dS71vbzXCElmaore9453K+4pe/ZFMfW8ASk5us+9pUwbDoVi344F5/13S41dansS
Vm6ZVnx4WKFzBYiGgNLWo+DHtz6lNZBdJPsT0QvS/MBh81q3OAEkQvL5HTI5g31z
lxKMIpI+MaSQFHRk01V67lmhpVBJSHaD2cSSA5I5/OUWx/DPDKk91tyBF46ihGC1
S0opxUu+ntIAr+EIQ0Foloa0hLyhzgwlFV9DSYo0zcL64/LLc1iaxDcHvFGbtTZa
5x7pQq8ysFc8j5L7QB3D0fe8up8xmo+p7NirvqQVINzRBPAiIe/hXM4GX/uz/hLM
QaIE0f4JunY7zWH/ux4iiZk+L4F0ssUw2KpiK1R/6AVapPjEHhtlImHQbd5q7f4l
spT7JbshDrvtxCmGR/pPuOVJrh78Ws7YMg10bu85pM4iHQnFoLSAi4AX4go4XAjT
yb8sjDrjkbtL0HJOh9TNBlBTuZa8YAaN9siqLuzNt2GIDS+phoQNESl1ijvPvgjW
h6HFqVOKk8U+WiFAj2LoOxvme8NpIRhF9+Yzhtps7+jFRFEvXsdPt6VQfxdwjx8Y
/ccETT8PmK2Lrw/B/R4FbnYZFSxsOxMCsxNHdlp7QPefCABpljSaHXwdVcGTj7Qi
IXcwHKYShjNG06rEhcMQbhpCDw0OlPzZcxChCCn1v777dQXZAGx/MlSCOA+/0Rcw
kd+R+j8rYfg/ylG1CLtsiJ4bZBTqEp8yv1EqSf5/V0hij71arzZw9hEe6mdpOspi
7x5syFMpH/OxEoNGNKpZ0acChhlRDmnGPhGvj9YadpOTYHUVisbrmoPZkAoCJ94P
hJ/5lsNwQ5DYPV6xGs33U51GXQVOjvO8g5GmCwXONYFQSSn6ydjy3SAY3c1MpLcS
2A/8ySmEOwWrtvMocNHscH8FVUXQ4aFAB90eFY2K+xCyd+baNuDxvhF1DUyA1EPQ
z2iPVjNgTM6hQe0ROrIfj0H8p9+XTVr/77t9tTCS/nZlkn4pfxlBU1RdDp9GEL+D
47/83Abz3ZHkQrAjEIk96LGFmUSuFrzpp9seCFSyYQxPyABbwDwMOIrDhwMqNmP1
o+zZx6DB5XPvfrEkmNn4QVmDYadrny9WLsylpggvwjta2fJUH7paxRrGsWzNrJY5
7Br38glJ7l5hZD9zB5bunHPOAsQltvlmWWnZCYNlI47VmcLJUpVjddsI2TAWk1Uo
ccaMDBsGeQ7+zHVPXF8eQ9SWGFNvYcRL9oEC+biapTXJqY+4ygCO97w2+0teBI5X
7VhOEhKgX+ehTQUZ8UZe38drz5KMdzgOXQDo7euCy9wJgxNrj3O2USbqte+3Zm90
FJTiqMAKjxYaWppu1sD+zOFuBhXp98GHMhoo9SKlecSE9GSXT75dGBZrxsowoY5T
VexE1yyvl9S82W4sPWEvVnx5jFZ5tFpGsD6DCbbkFej0VIKegtf0VcQacDK0t1C4
byRbvqwLjBCZ72AvLOaFvcB1j2Vj8h0GWD97CHXQyoETuFVwBrZwzZepp03U2aez
8VysW8wS7AUx6pWxH8CJiIceNbBHje+24xD8nluaeJwkyAJD/EBsda6XizDeGSMC
xr8DGyzbxQ7/Exp71gsmwUauI/jjMnWiNpXlOd1Ja52dValgeTwxmPoOEF828PoF
FkqiljBtaCXPgZ4Zzhkf0Y99O/kEP7YHntb9Ow2q4JYu2R2a0ZLS+EsAhgLs/40i
y4Ahf1iSW2+azzhpKrKaWlHGarhAeSAG5xrwXvrb2ezbTfgw8riaUNKIJX7rcPX6
WPRAFWeQcLx/lU/6HksDoLqkLS0GdnPI4CVkXYyI0G1F6JaL0PL4xGiRSI7tQde5
QR73KQBMXhAt0n40JRnQxGm7hvztX+mZcMgW3tYaeaphuO0EiFazgXdmjAhJTC6X
PzPsfFE3uY3r+Vmlj2YpaK+VSwQAW9XR3JsjS/KrmWNCh3bhzW7txlaLzi4c+snq
JH8dmUj9vrTi9L2g3ColWzkas4TJ7DY2iCfLC/IO+pXq7n5yrUmZIBhTVndVIipB
aZ/eKiBX8mDqkC30DPZjMu7cPh+DYzCmmD7yQ5CF5Lb60SzCisOgDO30GfNctPdy
TNPXO2Dw1Qk8//dTSyZ3gRegD3mzwpNyu/7chBT5AJ8GJzhig3GNWIYAwVrFkYfC
AEUz0cn8WB3j1RjlLxwQblcnfIlLR+JyhQyDeiTmMGwBhH5KA9jvTHAbkKn/Jx0B
0cTd4qiowb+oCmDvwxtL+z6qJXADKGDbo0cUL1eovlXgfEkkydW1omgZtvI5d1uO
GqTvJbIGda1l89fRnYetBDuAIhu4Ta7IVsAt4JC6WCmnTbnAdo06qjs1jfYbQ53l
HNR39fWMQWjc3+l9mjdJdeVnvGtKhKOYF7NwcjzKLrkXsHMBfsLKq5pxlc7yjj1p
emY6Q2R6s+ETSbxlD80hZuhnu7/tmQqQWFdWBmJAQX8ArYLIBorfUGrBj1aAa/wU
QIMA0xLBzCmFN7DAOKyfPHISyL0T+xDERctZKdkZUAQMP00v1nAxuEqU6cbMj+3V
JepmNwT6P4RsjfYsTXdzOtJ15+RZRpXPwq1Ymot6W/H6naMJrY+jzXHVUh55s8M8
G2K/cTLqp9E1G8mbT/LUErCcNZUUui/MpjXSX+LblRr21d6KcQ9BUozvOwS+uZqc
Jygb0/oyEArs9KiAq64bisQ0gyq+YE7pafpEfdwOSlR30gVmodbMUt2w52PViByx
Y488QXxhbjYdMmM4oOSLw5fzO9CJfmfc8r1G726FsAeh7yUBgMtFpBraGwcKOSwD
8f6rrAOaCv4/8DmQG2PHmNcCG8ODwnMcFrw3sp675xtYceQINIQhfuEfdabSTkgw
U8h4U+1EzgLvNXFyX1Jl34m0djutK2XG69/98qkKm6vVOpNMt2+fJ1fP2bp0vR30
Zcr1pZ66qi4frsjJ/0IQzzkQONzWy9RLImJ1SEovXX05GlFqfNCOal3KgvFQeAjX
e9vg2rftebP+Upcs+HwYxa3/o89FoJ3yYXz+6sZa6EmkncbaftRm5eXIbsmxY0f8
kJrgukyYvOppo/oVhOf95CHD81OQtiCmD8SSzKzJqRAapAvU/tZh4fvGN/TB2uov
bT75uFkKmmtebRJBxLmMZNL4oZREOiheQreUK6JP5b/jd9NE6BgOUh3aVjtQr/J+
4eECBoFySclDFTJChwf5SyULHUM3ACwHa7+BNm5Sw1F3QLTYbRntLayy0Sddyc8h
tlwJiXHlUxrmzgec1gdhihSUHdV2b4xB05d/wPJzSzkzvknSTveBCqlbwdpdso+D
vAyUmxmB95fYnYnhQSGz63sVMZzxp5+eZetbBCVfoyc4uWU5Qm5KbECExqofGx5J
BdtB5iuoSoQopwOOKCv+ZveJdienGLpNbn7eBR7fHYg1/2kZGEbI4FAxTX4G9tBJ
PuH50q2s9Kh3af+xR14OQa+GG/uND6s67O6pMrbYxpUI3xuGb9LS9YBEPOI/OJ/U
uB+dz6MtfJyrnOnyBCLHZ+s03hY4Hzp+nreI1KuaSef5sgx0KiKdEfoGOzjVjuVx
1ywKd7DuOBnhskGiAF9NS+KwRiEOKZHZMNpfFurAz4HqD67k63OoVadl+15bzu7x
lMxMzpMqxTBg6EEvx0sHsomABKkYqKsudVw9o32uZVm8lADy7hiUkIr3XHSzirXp
o11ULVZYSr2D67VUPUrwV1txk5/15LXS5zYLqknS/l3ZG46Db0D7UGiYjbJ/n37t
CBJ+KBDDFuejBz5uflYO3oVfRCyiIt8J2j4wBBKGx8Naarc780hIMk1ZKsDiQupi
29OxD8BldD0qLuWJ1amXnJUwlQlGL6b/Sak7IqZSTxy7tezMN7rjvPeOMECLqVhC
TZHiVXjKzORnDwtnb/blbHguw5o0+31wOoqBlV+d2QzZ7u8kty6s5s5yiB/AEMAD
SZlvcM992gX267oi2F9KVMy2e3m8QK0wRhcqW/+aegOL0mbS16sUSPZI/4KMoezZ
D4oKuGWdCzBkAbN+eaLfNuhZ5qlQUaVyHzlATtWc/st9gFprD6nEkfBfh+zICfln
1wPaUBHAWlib78FVCUsD2mPzlwiFuo9CPQUC+I4f93JyIOfjzwdqnZ33HweKLm3d
PhQjyJkGcP7Hkxvi2J/tx4i3DlPT1K4t9v1WzVzQLB3UBa75Yk1lGUe33diExKdz
XLE02h9iUwCFa4XxdRjfR1PNTZfxCGNd7fJyRJUUV8IgKXODgUQLLKdfvuPKlfQL
jKrSCmJTjSBbXgR/0tMQdKCScGW8x5S/TyAjZ8sZzYv+Hez9Y0C7+Asv5HNKd5za
zCNvWj20yayyHT1ZQU791H93pwDZ5Cq/A1P8ZTaAU0uUGlVa2Vf2448ahtpr8A1V
2F8ivgZROKnntyWkfIwff6Hr7ZVAlBFvofxqteo4dbxx86/lzBRCrFHMe2FYWcId
rW/f0aymeb3W1FdqVnLIsAcmBHtkpC5LOiQZjBkuHNjN+5uUnfcoJI/2LuR0mZPU
9sHOxPDoX5zjhh8oJigjQEuHQ9NQ05fXrRmw0PHA+yoZ00GBueTq2OmHXhgqFnTq
H56FuZ2YhfA3TRn96S1fB+HMKRkA0lHZLw6gkfGy1m9aQmnYFXHHAe2s0z91pC/G
hjwvGo3IZCS+/EtUtUxhEDDWQ7itqM9rdoudEGv7ve9orEfHpVKkecMHEm+Ah382
EZh86dUL7fSJuNUcYJDDi0Hif6R/lbLjvO8K/6QpCl2c3vTHcBGteXqu9q9qSfZe
KUIKA/9gSs+B4xswYLv7nKud+0CByTx4tHVvwdRQTXiuXXEAuaqF7EogSuVKAVU0
ilcPKDe2wXoOaIkaIDu0kO1agh8F2L6h0ba7a98ahN6buGG5l0Pe88j5AD0ZKMLP
0ngr9lzDUJ9vwGAeLBlQT6rmQJ9EEbS7nNXjz92J/AmeS20Nld9QYhPhkLPXctiW
RRbtPoHqxYYq01VwJc+0q34YIgKBTuwRrl3iDaft3XP27xV6JXkIf6+k1cq2ePaa
LUmPgEKHdGLjw13qexSB1I6nxzxJqlzHohHY5MP+fHGheStCbYfX+UjhELWzkr2b
Kq1D7lOCo9iGXPYagxiY8V+IcGEwJyg2/wXqykaIaQViVzBPw4+bAS65KhctPijR
tslY0tjCT4qX998kyToYYdZrnWflyVlBOJ2mckGJ4qXH3KW+Ppp1uYyK70DJIx7o
RQTH3gbMGzEUrA49YxPbKbvh+EelO84hwKySpsFdLKraBYOFt+gaeaWiy4cPTtGK
DCCzoY8Fd9JEbYml9cvGecSkoLCyzJXiFeCjy2YgraFAXzdZJh9nzlE0cQqO4Jv9
XJ1oBcK2Fr40aPLDnr7RaddXfwKXqgEqOhD0SMBNyzJGUc2s2EMhvo2aWg67bnkL
FJoOFUv3O2GUfFbGc/vFptenqA9ghNOE7F4tZ+9M4l5anvFnQ4fIymftxmdFiLGx
tpERj3f47lt07ZV2inyf+TyUB5VzbmTViurI38zbs5QZ8uyZq1/V7sdMluPq5UHX
luQ3ORcyyPXrCOJqomdfw9XSPfppsenduwvaawH49jGDK35xYkQt+FvnVpiIPmaW
C3bb7bvRm3mnZMKdulNyfVdqOCy77/1rhM0QQx0yopwiOSwWjtDAiaC/WGpXNLxE
PHHerJr6E8BvlCiiDNWeFMXi/a7R7sD3eSIcx5o0hzt5svvPu0Zq/7e+6635377M
DRfrvpSY3rEWVV0gm+TRbkY7yvC4osuYA9SDmftp8WM4E8VNrcak2HS+BYIC9UIk
TV3YWuCuQSqdRnDx/gtOL72FeLXtPiplUPE9lSD6LBFsFhIrYZFH7vBXotWYVgJK
l1bbGq6LGvmiJUstW3X8+VoI32410qOJB1ZOziv6fdgt0OiOSL5Xa/gMJ8VKppVu
iLxlj8zIg5yK1litI+ef6IrIj2QhE1GSG0EjlhtBeJ0zZoZ5stRxYEZ65EPZbKp5
JYW/18YpQ+fndXbnYNytQzD7X54Yd4BJRzHcI16D3YtbjJxrxAKaNp7lnQRkm5QK
75gkp/6VrVpm6mvgujdcJabiKgqDmcEy9IUX+xBXkUc4GvOfC6B4Anx2Rj6qDJyP
jtwsOKq4WcI7btFirfDWFw+huKSO8k3v2r3mqsP5cQWzAKoTqBJ1LKf0lDvAetKU
j/0fy5C2ZFQke7BCseYz3ig9Xr1/1vrTmKbH4ktyYd2pBYf1nWunPNZQL14flAcB
PfzGmBv2NjqTxXjppoevEYc7Em5ivzNdCaj/lQQeETBnljcWNRagYcNzeE+y4bZi
ALzFuI9qv3K4sFsr7JJyfqb6LUdTuqIYlIHWvJmVFvq1NBc84zqL747qK1lVk96j
HYQu0VSogivNKVEjv+7W/wnhBlB0O9gBunwhabm+gTZus3C5DJ6NZxuhSid0dp7W
DDxgQb9SEBHnx6cr8kRXPrSn/aKHQ5R6mVrGOiJnJ8CTdAaRJ7veCQxPH1y4319g
lNbK1Nq73ndgq/Lf/zH2vm/362YP++9xKadwRQszm+n+KMiTNdd9pI4jbHXdsMpk
FRlu4LfztPLfFhzq9d4aCz8tGF7nBvZ6UdCszCOS4TviHNWd6ZmsmJcd5gKzb8h2
QQRxKYZLOudZWpl2lRVRYyj3Yvs3V0kLHA1/W7eHNGDD0MRyf4628DJUjzY6zVh9
d80ei/1MxzLCqs+SYlG2Ej17fpd5LluWOvYPO/iFCRuIwfT/pPA54ax7sO2Dvql6
DQkjQjAn5ptNLbyquNJ9Emd7fH6wEhMgbdaPY8wyPsWvtTPovSjCeRMOAEO8+GTx
GL4loNjIoSKarcoucBO4cIlTWnU+g/Fp+7643KTyCVguYaVyo9fZAmxy8c3cg1Uf
Mx3FddNSU3KywfukpWs6j309BA2G6XMoOnZ53gh/d2jJtfNqznzk/WazNG1COUFl
1xeg2BRvykJPyzlvDTozVc4pUH6DbLmoafpVK0cyZ/1O96YlxzWGHf7yKbS96OqN
46l45Yim0RLvUgxUwE2ZK/Kl5n4nudQ4tewbsXcvmjDFgg6XJIeWgV2domMO+OQq
ThNJEG4CfqDBPdJEid0P6MEl+HG8YAZ2r9fH0AwDXo54pCJBPwGH/IPbVD25TUAs
D1YvCFVAG32VfMGRkqXJxRSKtjrIRVD2KDOb5Q77ftys6j/+/thzbqYHpXB225Qe
ywGj1T1ygbO8njDgayVZRUN6a7ehAd6D0wlQFNdm9o/afoUWZ/035D9nKbYEUofz
bi9dR23FZmWJjr0vdBzE6zQJMc/yXGOhCLoc/+Bbxgw2o/RRR4s86r5KHv7tJvH5
T6Nebh2EOIT/bzb2S8WcpRYTk02Yi7RmJkCMfSiHaW0g3Wh+Ju178e75HcZiDhTW
MGB57YSojNNDJzz+/3spuz72jOUGBhus/mZsDA45k7CqiWjGhcIoJQ3Lxbnzv8RG
nqsBcxEn24QQBC6wQTXIgYLkDpk4jYRnkcBoGpW9+Ik0SU2o6L29Pcf/nl2nWLvY
r+zWeQbAO8tRUCs+gxybpFiD/jv6sDMUoDOBoqzutNq1Mgm8aXHpBDCDEC0WNROV
M02sfZEhXD+V+9qWTObCcdh7fnY/wb60wIfNUozCWUenoEjkqZsBPg4CjVDP8dDl
4hUuiwW2iPg9QEGJVFMTu/zkAQ5oJ+1YHnw0WZ2VC2VeNj+G3uYYpd/nOcRct9K5
JZQ4uBdiQwEwktNWCJpAG8H077iYAq1xox9K6mSOOvWiVFyp90u9Ud6SAqHL+ZMX
UQMtqDO0K8OMSAReoC8LY9StIKhmkDCkYoQkHf1dwkLeOa4B7ygXutnzoZKmfiCL
MZ7/k62WTnMP4I2F6+T3kl0h//p/RvYFfoJymuoGMTKP6FxxhSLY7wmjpV8aq8tb
hDK1G0YfDGeilaXlllg30WO+cndSC3WsjyAOCWmAg+tZph6C3cXbVWh9xkQdLrNw
D8DRddeHsxoN7gdjjIWFrtO3sYr/8aCoNxqSyzUwbq8CyWJLfKf34i0pfcZj40yN
D251XQBWEjYlv5XQoeIEpDWcFWyn4WmDhtg9FWTc4+g3KGqweGDxIiu3Fe2qRvmR
nNsGhNeW8oThcynZhabpAehzi9s2/vO8F0tM6OZ50575B3Z7cu8U7RHKOXkhsk7w
otlqP0/FkKRoVRBPPKhQFNTDwLyVtjFL6aL25cOMjKlPIRVU9s9OLu23Jz5uuLz8
HvyR0XC5uhPfQv+OeykE2xsfROgY4OZtnfcnyeq2rCNQXrdxBT1xqzwo3Q1K2117
sNSL0lOz39WCAi7+Lx3h037uuSMChbHgSFs23o2oT/Nw3t0nE+ocWPG5T1+oFAWA
vq934YcLmc+/sptmx6FPVM+xYzFFxyfwfybYpJXckYGHdVtBLaH5DAAfk6K6EOqj
0n2ZRJOrrc43BRHkxFwP9EOXgglZbTdt/UiE/iHtUQyiwBJlOMOGVKcAeRWDjUZG
I7YxXY9duRv+tOnG5cRA9aeG01LYKBndTUBcDMNGXu0FFoUdQHseENEjHABxVX/p
mP8vgmsbyBgvCDCX4dLrFvKoWCCz11RlN6RgbBhtc3VRY1BqOdMvdbEL/5LtmXeT
OTTUncZwlGMsKJ9AD+DG0qaWQo6dL40pbVJy+qpzEe3S8eL4tHr9GmC2BO4Vl7vB
z+OHa1eMgpmnDmXcs940JP1/4xMmdup3VXnh0fOyyyMdCRWBPIicjIXq+i9L0sHN
O50LMfpbJDYYAEz9CoMATsmvc80hOyQtN+HUOvh3o29q4mji+Dysh81H2E8jJUYn
iqY50Sl/dizrLewryqwWKt/mDp/zUT58jgkpK2DvBEYrYiydYhLE3mGiQfV6x0xo
3aWrYzLblJmjPpgGEQr3aDV7zSWPEeFp1TXChuOMq4Q0jaPNn2QzkD/PdV4x6OF5
ERmiEVdv7kjr4YlBcWmLVTNqGELYigV+8Gq8TK+Sf4T45e4ZAf6GyGcgt3xLzjdq
tnBqv4mgNe7vYqIG9uaKYllAWpcSHOFY+4iMt3MJGCdo+9yt/QaCEcZg6cvcm06+
y/OBmydjxj8ncpc2hqCN4XjuT2a0a4kIfnYwaGb4zuCCe3nTdcV/zMtGiT99AYwR
/kwLdoi/wHAgD+ALl91g532LrSXC/tF5lHxn/B4vqnsxhDNsrdpjXJiu+WYq88j0
YlkFkznAk1WjzpdPpZV46xRvT07wpKKg/gYRCctj+iyKmXGjxKhkLELX0biNvRa/
gq2bsRW6CPpEL9tJR87jZ97MTOQ4Ek3WIJSIbdEe4ECdi/t03kmsDWozAEjNJvCe
/N9wq90b56rpL+0DBrweu2QDA2LELE6TRwyinRmJeXJHAyjocSeBCLiv49t+Lioq
GffgayZnoGA4j9/G7IR3iEuJ8cTUCOs6Ap77w9yxFnij9EF37v8A/nRK0IDAUUE3
n767H0z/XIHkE9W/tSnIGZt4+aukjRtyC71V1J6x7PyNB5B/DYLjhhqA9mVR2wBb
7/3PrJYYvClE6XX6VBza/U6s3U7UfMk0b5ublX3xjCKQpuTQGSqTAzjNscH2VN7h
poeiOeCpQb0R9/Fnp4esRG2fIqFIKNyITzf0hGTntfpjLaE4N+oIhcCIZgW9nodU
27xcSj6yoZrjKCNeW/dyAY+CpK9Xeht49NFH/sW+FSM2WCnnSTGVtFsLsKmXu1kF
hQnwTVhpStbaYvtr4RTBptADpd+CuDv97MxwXeezXVkr/J9UapPmgDNLzx2gl83Y
WVaHcj9M+kRfRAojCTT0WadYJGPQRd/iDUY74nPxVTz1bEDuIltJXP+EOSVV5Ruu
aXNUMN8+0emE2IlpuobJcx00k2bMogTvW5vBA7SJSQX8Wi/PcUi4QJRxKmU1HO3a
pxczID6EZeUhQXEE9q+9+9hA9Loqz0Fh3etCxBCYZw7fnqWie2M/LBBL2u8hZPEw
zGXkyf1RSqf+i/mW9WLWv+8rKiC7jqyTyD+CM70UM1maLDa9BpQpdJo8XoBMos4i
JBGp7icbTQTU0IMDEoGHzM06/wVmlIH83AThuSzFVGcnXwmiQuQHXy6QkmVjCAMZ
xzBaWbDccsvVFxOpW1tGodwH2Gjptqi2HV0eWHY4FPU05YUFX5o1e+rSg737AdKt
r6p0OfRWi8f5xl9xdFXbQHE7R9KrcYRVLX+2l+2ikBz2V/5GeLVrZfGjNhMtm5sq
uqM3Se6AjtTwL+V8IKOM+IdKAsVGE3k1C11DLAPjrFodeveIj7vJoxQaJ207SDiq
NRk6GxYMGlE9lbFglNOD9SjR6CDlcgv4Qt4brQP4LZvuypXd0/3MNU3u73K4Uu+V
7hdzsOvRf0+c4Kpf9mqRbHMmxlvQ/ftNUypX2eg9TINYM7v2oRdpilIwoqL68Wkz
0nxpFvJpbUWFay2wv5vQOi1ygtyA4ZBUFPGrHMSHKYXI3/s7gE8YAmw0CJYKj8LP
PRaev41+oPymgCYMdOtcTzb/m+ttO5K/C18oL7H6ac2w/R3uIeK61XklihXeW1U4
vYM6sXcslJBoB1ULniHi3JmrCCPnW2sAb+dV35OeOYke75NmLZTOSMkdCOJDd6cT
dSRfhUHE0ZO67k7CkyjkHyoOhaA02AK5gRq1gMqZKALgd0HA1dApxItMuP3MFIUd
9qrNuuWa7uBRa7eRz9IhsSo9Ohw0KIER27oppV9Lm0YQrZVa/j0B+EN6SvHVG2fU
w3CdPtEpQXnJX58UxjyUZ38tj0H34pVJcYi5IpyxNxsgIHk+/EKgT2rqgAbd+BOA
m0BA4QAyPgGw/qJbRBIGLrZz8U1zNNKB1OfiWEBw1v9zZ6tAyl8wNCOQyI4WOREu
Ek7WTqQBVyLQRlfzIkUICw+MnkQBdC+nKREUEgrTvhWtfDn4bAAns6MEc7sB+M88
xhqccN53eCx8FO5rOax70Y2zhuReEX99fg58qHLe+vKYnfNMSNlg1onrzRbq0YDm
hC/Z7JzSe+yOf/Gbcgl6saZZo+vAo7qrzjQQ0xg5gV9bYmSJtL6tN+b8WSgegex/
kwr+zxh5zHHdzi8tnM2gwCRG9zXouEcTNDEZ2ma+bSg9Z8lfRooaGMAm/ok+iSo2
6pe626w5+SiukHzNmdrDM0ZP6J+CbeAuORf4NQWxUA3RK+zHEUam/KkNQ30gBB6X
u4p3sOUUKMPpKCYAwcWu3NdbkyIRXO8zUgdiYMVhChAxaaMlD9KKtH9zmLvrFV7A
QR8kwLP9x8Y99cxpVSN7ZXADEgRJVE24nXC8hIDEg3jtDPDKP5iMvXNFYYQmwRQv
BXErhSgo4MoieZho6eXi4BRMhcwI1oWf01Yhi5BEIRZOuF9A56XNcu3sayVex8sl
YA4nHf1jb4A41o5ClRLPQPToAZSPpqPb2utTG7lCeo6PzlmL6StMuJ3yMQAy3bJb
MkcswHdaavTQhu2LSrXeI99hCuvw9vvuvZVS1kUYyvKqpFOTFvTJMSLIyPFlKO0z
pgNPDvhFLFX/eoyDFQOC5rY5dPVfaNJI7p+8Zdpe3vlmQF7FgN+pCQymNhQ2Qzcf
rAHZW5Yeh6wUdrmSklIOEr7t5pVmbmNrR6wuFvqGgeoese+AbFJm2hj3rEIXKNEG
UdgwxWwQP9bQ62B7u5cgFd4KIlBQssNzfaj87qTlgBdPOHEV0Tne2naIxYdzbP4+
Ge+9UAvu7TobVmerjBSVpxdhyPzUQ2L5tttTGnBgybw13KKIOZL5s0slAWutGIBD
F5lxfC9BWIyZQCBDbNGZvPY3sP8DRU6Hy4Aj+X5CxsxlSvZfMDUiE4pu7tgSg6xb
hm3iho3mZJt5cI+NK2lzG5tD/SXV8ji5UbENQYRSJy5DmJ8A8NIhqm8S8TyKtlb5
UiRAGEffXj0B3sOKhd403n7pv4YKZIKMCm9SDtkZiU6p8YgZdMFGJD97zQuBW3Ve
gk2wydbzHpyG3zqgzyjt+lC3BY47/a6KeCk4W9vN/HHXd8UlkSrs+Dj2PWwqW/5J
97oDetOd9G+lcy4EmfM+ifYad6zy1mO2MN1x3WgmcJ8AxnFvBNMOM+ZymfXSxLxY
BAbD/5MHIkFGDI90TMJQrQexV+6/1Yx4MNjRZEJDmllGqDxA4d5w11ZspmC+s5wA
5qQ+ibrl+Zn+q3QedAUpJu5LiN8tTaq7bOzgV0qNQ33FkI+Jc91XAY5XUe3APyfh
FyT3x85R0LLUGgRGChE72hFAFpPzsISN1Tgsng1kh8RrHqnOOCSwVLt3EEop6zyA
QtWXEeALae3p/3uKpVGp66uEP4ejOOKAbKdafFoy6lnDggFyhUMoI+L/Cxcx2ZH+
tTiHYnLlMPG+QN2S1ATlZtHQ+FQr/I10/YPD9yW6CPLyFn8vs0OiKkJKt8Aa/Rgb
V1htamM/s2qNAdaXytY7DY+BNpQgMWTGFOFqUpv0zqwZcu4Ql3NdH09vMKcXF1GY
mxQnbg0E9qhwbITA0EBUT+prrj+KpurgNoiIry7T57DIqsia66aRdBMbmYpw7rKX
nMsbeckG9/a5jWvUycf4QUrN+n1ThjxzkVOv1zNWyP8sAb8RU64/La15KL8np2ZF
FawNbeXyAZKnDWEm+TWTUXEPBElrlD+HrAR53YDA7XiboUWlrU4XW8Ukg3vZ/o3M
tHv6JcIxKY0ewvVpt+PYnYBzJAa2pArXa65wGMzEwQO13f1O5jCRhzfadj5Ng9mk
175Bv6N8/2CjlcQgbAT4MdnT+qBN3TUqTh9R6QXSqyTQ5BHWff2f+o9iLu0EbJiL
daLh58HDDx9x9Y+iOKybcN0NTF7c/qdAflHtLuk9r/GqnhUarK3CWNhVlN26SHDo
tXoA+aO1h8WxFNY6HKjO8Ug6zlAOCHgrwYym4IrwE+2wPGSm1ap3924rdyd/8ER5
Oi3d9f/Ce9StKrVn3Lc0yQKiAskr9N0TQrRrHyj9enfYxHGqK0sYRwg8Ygx7v3lr
wNsRFTGCMXdPapVqfA9IZWq+xDMC9b2JAnRkFi1LPMlOH+Tqojs8hNgmCQURf1v3
yVDGWILIu/RG0la/kgo6hULHmA5zzgnsqJvw6nKEpWdvvWWqejW6Upbe6BA4LHIY
kzfBQtZhsRxXNgoXk7+FrwULxV21eSc4wNdSbFbk2YhiVrN7BVmUUhGBaRta4VJj
l6gFKEvSKTpdtcfIwN6mDUp9WDJzESObVWxxQn23x1Jb72YonuMpRXpjpekzjKjY
nFivCLAbMPxDkOxxSUHV7NaCrMh+kLR1Y1DFdbW90SwY4LkmWy50p0Scf/psRcmW
ywYOfNNx5Zg8RQHtmq8wS2PMyVi42I2LIn5gsTTxaBWJbo0+pptXVkST0Kd5fH2g
g+avNtwBalYVBcTVPx8cRrNRZep2tOcvLD/DWR7MpX+LsA+asm7xlX98WpuR2K7I
y5qLXjkCfgqd/hhVERZh07r1pAL/QR3faKine3gcbwCIOeqPeb3HyHerBXvegGSK
Mpz8uGbw7H3BSxYU23nXSadl+OD5ScMdzqb7o9uEuSe/KQPvlW2R3ZvTyGmcBF1E
PB/oocVc5SiLD3S8475w4DpBy7cL9nplvIhpHngzlaQvRovckKFPQGHltTACGGA1
lDcsfFg+W/ioV0F8VgzCHmmGEMVZGAUtY6+TuSpy5X5fYx7/HFC8eNUTjgLX55np
i1b7AoCqQqYX1RSAJcR9Ub/6b3dhyRKC0ubNcXZ9X7v+YupvlAgq2Bl2fI5NqaGi
N4Rxpk/ODM/edWtlxZBDBmlxCVKSxZJly1QB+qDSJHw2aCX4iAUtc6VzGFmOabzS
+aQGzh+TSyqs5vt5hAfOTCCMcKP2DZwphMI+4FiCPcyfU8N9S4cPBQMZmWf3pXQA
NjqjBzZ2SolE1V27eB3OA0Ea9d/hIAGpnR2kIZ4XF64yoM2fRI1OEj86VIyv5Qd0
PXpX9nSDTRDTJzZ3M0tBl/DqgPDrU8603HZ53rmUOB1o15iGVDvPHP9G5gjrKyrY
OmrHVZcw/bbtf4dM72dsAmwOoxedEymQDJ2Zh0hdBSFXDsIhZQHwLdlCvdBULVj9
Qmeu+DeLlRsHyLFgUA73nBheiWzHe8g/bwyvD7LRI7edOtZ9T9z7r9+n15HJ6A+D
g5M97AQ+xoMin02e1Kovkmq7JNBd/uXTdKl4oIVMl/2L1pMPp3XzQVJ4AsD64byO
wrVpEqw4Rv5QAVaq4tgVal23t15v28fgry0gqhOPaQPLWF9guc80chKkUa7ynhZb
ucEflFNjo3GJSaZP6dNwCmLnJs/csrTuO4x/F9PL0/+DoISF1ZGXxdxO4pLoKLbj
cgiNgvTu44t2jdgeUM8rpmIPglTesAIZF8rrrbcWeA0084QMeyzFxbCDhe0UVG0t
elDkZFdYAfL368bet7usKfNIxACSE2RGU4Obdt+jteAVeP4GuMon5HZjy7Jfbh+8
dOLfz/jO1Wg0Bx9D5BuNi/mdt6/TdDz8BQbW5f34ME0Z7aMLaQWhl5LlYrd5bC8Q
7XlpA1rydqAJuh/UVZOKNU+AmG+O/hRnF7RegbvNy/Jt177qz8uyn7ZHcE/Ksa21
rDmvSTJvHm2mt3OrGcijOp17ukSlRKf6reMFnNyy69+SYyS7A4uJhCkOqu+2LMxC
PcjijvG3jaKXtTl+eI8LCpWglBGktKL+CFAzaGM3u52wccAhHUOJ3mHOm8+U98S2
HNenSCvPzFwrbBHgMdlPSx97YMrys+78pRkWP7ktmR4RsZtqhV1086op/4k0WuXq
Ps8J4/mG7wOHK42BZyOyl4V6VpS092pGeU3si4nXEijgY7kxD0HpN3QkamLQyKWV
VqB2kKdSYp+ef/anX6rJFryT46U23orpS9nmP98gQFYoNm6C4+W+E83b0Ivye0wv
8UbcmnVozMcq1X8rD5dwQeDNk//W79MHGRn/UpgltjYdhY9n6vcWCGqX9F/8SMaF
Qc7l65Mr6bbUmSjbywwYOL5YeFI0ajLmR6VPeaWWmf+TVdwZ1yZvbWUuSKnvz765
07YuHi2W1F1CWXrNHP4g9KyLhJUtcJggkJ2bX68t8fEs7v1fc9jC04A1W1KT/EhO
Ieb35DlDcfZ5hQf3xcM0TKLJlISb2rxOE3zONn0QoeFP8itxa/czO21APcBA/n+6
txYa2NIzLir63dL9Y7vhyQ/P3RmsLwXy2lU+RnDGtnLD1zKPhykjB2unaBrPAebH
XNYrfttvWsA0t2auHGF3ij2bYHvBYC2Kr+Cmd36l+6MwLROJ28TYBNV72vGL0e5/
uihsarwcex8vpBed7U/p7n8G5qIhxdmqSdaKRxaEGAo1y0KDRrSQp18uhb6Se63S
jleXEEk18aR2HWKa94uuo0mh+VLk9xPaeI+BlxStDHSMaRogq/TOaqNVIEhbC6bw
JJ4yN3uR6Agg2cYTaNAIaDbxwlisdZUsXm/bV2JYv4+F+OLjflLGX0cyaeoLM9Zu
XWjQKCeYA8+EBBJeHtrP2azPxLIJhF8UysX4nWc7DXmZ87iOfmV3izK3K16gDqMZ
0/Oq2D4YyVgzSOnLeFNCZBLim1RA1f3cWIPe+teKGdUdYyC61HL69I51QODrT5Fl
1rkOMxVHkd8f7bCNjPV/WYztvvVADM8YQ2lZ/8kPAqr2rb5kLT9/KORpg/wKdmGL
lhzsfA3k6QIiXFMBheET4tHeyUW/v5BCCOX4s739PRXk/9iT3kPTAZu2C+O87TLR
arA72QJeW77UIIDqeBq19Jr75LiLgehV4vt69FLa0e0LEgbFqR28qmQB8ItduVwX
Dvdrf1FXz9EjWCkeFx2EGnkccwpnRQAbNMWAEb2fkowKllVFD3r10wv2ccIAoAhV
rPqS4uorcu3QMPOVGbTUJqUbO+tZA40PVMzdOjZL6IOFjxh7Wm/PKNDlLCUmoej4
/BJ2/+rPInJQf/y8fTYYgoU1OpDRSQc7KtBFOu3/dSNJRtrSS/PatzxMMCged3OK
qt6jD9BsQx/p06fFvtLg0ZyDzQmGMVKanB8Fqh0UnlrKHDoIT6XmoEyvnn0w2cHF
Z9fKVMpOacCbQgzkDiu4sJtCxvNnWPoV000mqi0vKWVyFMrZEHAo8+ON/ClFrJL2
ywFu6u0zPalzdqJ65LlsFF++4Lgy4+n9tDHeF36A4/ttVtiBW0iWzWgO9ZkFHe8P
9f35vI6w9pZu3pCBnALE8edGvsEmss6jRqq+4r7wf5DWxq8B5v7B4tnCx7ekyslq
V4LzZEDbanLNn2YrNyhmDRKx8co+Vy02fcVVbYVcVwt4jR8uUJabdeLHhW7jVVl/
ERqNrcrmXaniKGWDEYY4hOBqEZr7m/wuWKoNusEV6MyZFYxS1EbvUqV8wS59+UH3
OxRt4qVbBSPZQ84Ymv+J4Ql4UL/bjXrz5AHIEp9CULY1CGnbnkxSf99yA5MlY94F
xT6eSief2A4eUh8lTPD9ZDBwymhrsH1Qt/mUn4NQ/ica8cxqL7Mok0RZ0hYw5bng
8XMxeef41TPxPmSia/lSjMb+Mufs2IAs9dpB8wmYAn6L/+CfpOEkKkTmagRT8WM9
03w8DihFQbpgAizXUfoR2H4TpHByr9xb9Zox+CreAjSlHYTVJnK5nJrpjOsQjF/A
Hznm7WQTok1aOVw8tMbfSkRS4OFjupKqnm3QD0cW90FvTBhUh5MdG2SbuIdGDgH1
P4GnRunbeFL4RyLp7QvGZyW8ZxLb/0e5JGgjW1HBOVUhvefOta+yWBVKuTenaxQc
tEKGr8Jp736Rxe5dPX6PU44DT6wg/hzotW/pSVHkNgYdOn7cQalfBGOyRRDvjpRz
90Yl/6gitXDgkwFfEoFDysT1P9/fvnlhhbmoukODTC2vjDVD/fnA2ZoOWxmPu1Zz
+OPUgz57FquUDLbJ5lKTN9IpyozAUl/2HQYyfF4aG+R7xj6olgHYCoA2bCFnDMys
wlYHNq6zpI8V4/rKyP9yirpyHzwrx8lIu+pfo81NvmC4bxluxOFLApBDhpHa1Gqv
lIICKBwYeGEMKqJxXFNgYRYSN704yB0NyngrDoXeGC/D4VP17wuhuWNsclU4q1fx
wUfa2FGvr0xdI+6UgtGBXSPOau+05h9VeQ2Mc7l31BwcZoqZguJ9h8NL0A60L5y9
3tr9720tKiAGzd2Xo4HsgV4Oys2JlFO55RV/tPRhkH7cqCr9POXtpakWGwkcn3RZ
mPirAY3RcqwRIZz+jYhnQj6tFAzx+duSbAqAvhwZvbIuROOnu7BtoW6R4D/oq9IW
1rrYL+N57tCE5sGAZ8EGnFQV6yLYQ6Qk99vijhrQ1WIomtfu1Pg2gMPH7DwEAtCE
KPnBtoXZoPfU3Clm12cPN5uNwm7jUX2qFMRtndlDiXbY8dZrUlsLM9gE+6unsG7d
mAtw2A58jyyKvxQ72sOBF9JVYQ3n9lTpaka6/sNHQ0fO77n/PeWaJ5QxVXAbujc1
LKWY+plXk5d2NJ9NZnvwhgUYkKNxDQH/OYCFNN/ch7mnIXVh63v5wn5rp01CGamZ
P4meQwMwhiYAyiO1KFKZ751K75AubyfB0s0LXKFgadK6W1wzlzmM/R/EaZdrpl3X
Hs8xMTVNqG+LEkXrfKDah8Qzu3Em3lUwHboz5W1g15qFh+2dIBo5wG1LxawsOlWM
XMN4A78gLuQ4Bq5htDNQav/6ND38os2p5qbjezaVfznkZniwKUReXiqqUG42xA8V
8m3oIZ7dEGkT+5dr3O3RgRd7x+/i0YPjTCRLCPfw2OXUemF1DapPavkcIjT0H4p7
eLU5cZ/esBFR8MR+Aztbn++OvQFcBcFhhq7+0apWvEbPeaT+lFDQkvI/KOzUa+Is
U+HH+cUom+bf4GAo0roVN0zDmOUSdtR+4SxmPzmIJM4wsNtQcc9KpgXO6yZdkzVF
OKYMphoNHCPn9SKEotrC19J0CyoF1O3amQbdPJVx3ExcKmsx9SXII2y8zSnFXS1m
UP22bFyK31+dksStBnF+x0tCNV3nPc+I/qr01aCPyvQMS/ICBrFCCCkb5i9+8VhM
0e7EJaA+J693Fj+tI+juUf9VG58Ks9vJ10pojUkINjtLT19Q7+XS2znEN0Dk3Qsg
DWfI5dD2w11vTlEvtdDnh+nXfyMULjET26GSPZFXCPNgLAr5/r96JH5PFCnFtNxy
jtNVnH0k3gsRE4RA0lslFj9r8x+cT3vpcasRy5+nPcRWhZK7uB0c4oEMP0I+ZMeC
cQQVQ/rSP62evbDLNCjCt651su3yYJpNeZ65Zz2cHm6rxLbfuB/qTS4bmUek2kTY
gDCWBnMY/+uWAAoEl+sa3s8ptwSh74gdJZFDK5waGqgf1bWFtGUKUzJGK8HE3ke0
NoM/IjUV6iJAlZ9vaGQIUYn0R1oN9izHBXeqnLumVhNcYVvzqSxDW9skzrKZSyK7
8B1HsF3R6Qanel8dNrIKZHsZUrUycPATZrQFN3PO+P0PFXhJDAbtc2e8WL95NIBs
lT4pq2mPPuLvL45UIAlg4vyEd/eCaKW2H09ouRaCM5fXtw6N4QkIGLN19293LORa
arb27QluYsO/rzwcEyh5WZcFSJ6M6P1wiAglRVMEVl2XFvZ9W5KJ2zVrlpas+6FW
M3LCzxkllc3WXgaYvTq6DWvsnu+Fxcb8Xm+TxZ7NqUgdmrUR5uHknt0yfWOBNfCd
QDKuZXVysiPqcIMjJUV9l/dAbHb/Y1od9lGtVimiV+OofiB2pZ64BKSp+aXMrmnE
Xwwoc8URWqdsEkXfTvU8qNY/QrqtigtEehzmzfB4ph18cuqbiKb+4MrlHkRhq9jU
etG1LsMHFBD/gGoAC/eWsMC9N1qJ4YaKlE4kdo0nIg9H4P9dyz7luCyF6WjBH2Bf
JZOHx4r0wFqsoW8E4v74VkkuIx3WWncwcrNRMfpW3qBfO6JfUNz//yCyS97FWrB5
3N1nkzaV7cFMLhtOaHyWS66FjUlS/AUng1lBcqhC+eiKei98fwr4Whu74g3NIgWY
34cFx2iyHfYxo0PAGdGqp8HUKZxmovH35tg+oA49nJR69q//PNQR+KaeyFwkAdbo
atGv9A932o63YIS2wWvnoN0gttjyB6YmpiAoqbF1iofNRafyfcvLml66Nhexxzrf
ndFmK84VoTFm1ohStibEmg58dpwdykw4fYHQ2IzAT7piJyse4Uo1ZloQ0OBv+OUP
39LhfDfE3etS/aUc0XkwPlAg3IGwcrtYf98VjRl0SOyltbQ+B6n9p/y9BKLfgO2R
fyFtoUsM8Z3m183FbVLJFoXH5D3pVWI1PZ2hap44IO7xN5ja33TNV0gpRRAvX41d
Rf37orA+okHatC7wWwLYIGvqYDlA5XDKtqPljmcvvikjts5rF/+89Sau6VI+rmXc
ZhPHeriamkI/vZP6EnkdMq2JAQYTHBjxZjFGWFw1wdjge/JPS4jKP0kf7DaRW43A
HQH3lPvhLVt5kve3yPS+4kS8PLHr0xLIdAdVhNtgCZbyW0Mo5KHfb3S0wiLX9A78
2vTHJRMa/hKtJs1wygeugi0UvaP1UlNjacsOvcejp6kGngjZir7ia41MQ0LFimlC
GtQGAwuJGLadKkBTzEW2zyUlSRQYI2QeJi44lrYCzQrMABlGREiV7hng1RyKXSnf
yP1NcCL98S3eYSwqpfYT4A+wVk016ZK36dhClFctT4R+mNh37BwFmma0PH01Kp0D
+jBNkVI4Q7PkFlgqbITgqFIeZOR0Ip8RC6LCUf1deco6R5ihVbSQSDIEljBox7Ic
orU9/seUmo2Rj5rgJipDYlOOoyxP5ZseT1mDAVJdLN+ElUyPMk8ZhWuAGPXiD51n
g16+T2tTPz9Vh2vS2dwpaLY2bT+xag3IJWtyHRKBMFQsVex0gEdgiNnEv6y0Qfqu
jqbITmGly3mv3b2jRoMtU/JiL+O3JR1PFC+ziewarBd+8fedtwvydspOZKRztLhT
9CQUrdEeT40jhq1gwBZOvORYub+6KS3//SwtP3gG+URxxEAMgW781gwg2DG4z/CO
YJuJjTETipgYcPmt7BMKc3DaYdC4n4AT6tNp1Q2dQnfSireZTU9zgFisVb7r5R8v
+YrNgpS9n0z5A5Qgfy2QiP/JvUhPOPDgOvE4kLPtVsZXwsHiP+q+lyhIhcyWOsuR
IilYltzvaJId6dczXBx6oBfBaHIa4vIvEB70YI3vTEvS+6A6H2OXhsZnz8KkrGcS
EYDfQGBgWY9mz64PsU7MbDy9cK7ckyG2f9HI0+v3Gqi/NTnDATsc7ujHRPNrRMNU
LkPXPIgWp5N6TOGqDnKk0E2jnDFC6CI8YLMeZBuvVtP4Ixnbn2ecfllfWUYhMImh
IBmR17zg+AiM6Z+5BcKMtlRhMECcYPUgUvtfc0rlGZ0FopUbge15Wc+JBXBlVrD8
Egao0GNwMCnymE+ZmoMOJ20v6qI+6LrCPxXUNpDSnsfFhDxBCpL2JtGIIgyM8zYY
Ld4l12vIt5lcqWMTbEaZ6+8sBtIlIIQUx4kYeVtwvDm7LxyHDn68TIn3v95MsD4c
T5QNvlFh6CBVPf46w0tD2PDtADtj0RPl5BpIzkqx5FX3sDKcKTsYTrSGH+h+nrWI
EWaIIW/H9jnsc0xX8WPPF4GMLgb391ELCwWb0f0HqP0tXFkCKZ4F0lQKrkwoLGp3
+rtVoBjUE5mk1b7t9kdH3mbaRHi2pLoHU0p7odJ14nWUiJPdzgKnK9fb/freZP9c
JxOAppU7OuDI7yNkW9LPVvoNb67dGVz3nU649HJZ4S8ArwAS4SEC0nQ92a27OI+u
sea4rBd9WmmRnmIxaK+CnTmHzQ27KHbvO+JtXweNvvZmwxy2xSymCF5uYi9JH1FY
hzE+2Nmd+90tbtKHTTojiLAsI/f8EUjeImVvkfKz41RW4t2+Nmq1n2vV0EdbcGbh
16HQ44CZOimGRGmrIQ5wvFjz/8Efmqe2lw0enYyCowSdecm/dDUsKwnllIhDBzjQ
fVwWgcpP/l9XPn2mh74pVHvi3sx7AQFPls8rCf8DVlpanuBb4JpZzQltVhunL/GN
RK7Qupn0xUELK+C6hhd7/AyKS2xJ2sYrSWV/O6IhTjKKJb4w1bHi7Oq+n/7oz+4Q
jQOGR0q/bnWh/5gvkPNhoiZ1feIUPLlqSXu4FzPu086FIJ44safJw7GMuSZdd40U
lKTLzvfig1VfQU6hfZ91iNGjfnxRH3VdpAyrBl26QdaE+RK7T44fxe2Qhrr1FtlN
Ux4Wx1EDSw7165ATLGWrRLWTguDxE0U+i/TXPMYcIW43ccFKR6DoVmDxEH77BrD0
dsEns8FI9F4/AJr3S1nddaKCaxodTIt+gCHANeN7F003YUOxXtKwa9jyD63zVBqp
9GOZbtQ+frghvyuOTnwSOe1KkLBvgDJ2dM1TobmxSQWjAJtY61ndZfsYDlVE0ULh
4y7cEgMGqcx7J16nDhP63LFp3XCiQYY49S1aTVqGG7Zf8mirF5ck+kL+SYQT46re
WC/4R7p6rNlG/d5VGvRXgNRMYlqHrQ0lvW39WmRPB8xL5/cCuXo7grQ1FNO10cv9
K8bQHfYDmddltYpwLYjnaMCHEbfzOvX4tRxXFuC2Duy6grb16Ipx7NLfay7qNMdQ
i2jZ2ea8O1PTjYTWI8H90em4bgti1+pTZtUOz6pzzHXIWW4uQ2dddeO9OmEwslB3
YLZuuqbArOZSdaqVqxqfj47+K9018OZlAPwYsang04yVOdsJGLe7Y7lRPmJorzrF
PV9t3INo4K+AjbrAN5OyWYsbgwncd3v0OKFSnV/YGNZcjVXrmd9UcmgQnPZsEy+h
9bnB5dBywcHlY8Yx3Z7ukfC/zA5/LWb9RULmDctz6p32oY0fDHndCfHKSc2jVFF4
R8wueHcZdH5GNGT5mcwJuY5FvYaRAJMxpxekjmeeHLDW3sk1x8vmVGoK/xEBMXij
ksjJHBQW1IDJyMEl6iYYd0dP1QOqb67A/LsGfzZNuBaPglHLuILvZqTy8f2G/B6V
XvApER3utqh84HigD7rGRMoQPBheLdiyW9/JRbFEc6GjLsN3QG5LPBJgKXEl0sPa
K80j9z8abtPFAnWUS+RalE4GLAuqaOOUVKwF6smIrLM5Tw1sHj/olI0impIncoXM
9Pf2dwpU+C2Kqq4iw2D/3oWNHw8s6hF8ORi/v8JjEl9MrZFPZWCAbOKFzsfrG2p9
HkHt3roIO+wi40+vNq6eyiON1T90Lam7rdGUytxRia2tzUInxfjZ7hOcP7d+bM/3
SKYgetwoSi23YaItiBrAcUMfCgrlkB9Vh64bc5/rpIphXNPAK2+IR6e3N4G/XJBr
/pTYQfbuADdBuXOCXox2sFgo22OMHlccszzy/5K+t33HmUYx5wdjuDdevNSx1gjN
e03lQMqx+roCAr2hQTDn1TUAHFOhiu64lYbb13bwBdpqVqUd8f3/L1XXLeyjRvp7
C/j9VBO2aPS7ePuiwdhqANxJrmZBcvjjPw5WMDhMManWrqaXtkk7ySmnIMPZiuJ+
2DYVxsl/l8ibGMP0QfJ9buxy5/spsqgXYJ8S5JdhYC69zjpxVl2eV3Ez1dwAigcd
ccKyW5v8rPl3qaqjNGujWP8xwep2+a85f5rzr4I2VwcZzOoE84qGdrpg+cTsqDtM
+lA0K2zC0xQJ13tYUrL1akQCH/vva/GhXdfwXZfXtc+MBzC3fP0ZVdcRuoofLapt
PV9JZmNTI1/yNTxDoTo6EHA+5p/nQ+0lXdHQ5Fx93gffqiOUxoYRJ1cZks0sy8kL
G+Y87YBoqlnH7FdspuC63ju8mcWFz6LXocA80ygIKiOeTFc71+rsLCDi5TiI/DR0
gF1qnfZ8iQIPGi2/O4/iyt8stI0pOqqgNTeQx/Z8B8gEQU+QVMz1Fid+/S8hYCD2
sZD69Wt9iblEu4VZACyLkbN0BuN6E45cnXQxEYsmxUbZMDPro3o1hX1mxEvvCLCZ
Z9mEJhqE7p3NwCHQ+bH9Nhs6YhkFhY6aq83ehi8N+SaOP2xs5nLPk5N7GB2xVnse
CmKUNpIYVjH0/Np2roUCbb0kgUsYWFJIOpTTOCUZTbyJf+BE+0NrG0aH7pYFW5uT
gKJzLJZY3PHNe08m+z8Kfd9jdDW5GJt/j3pRtrlWXXwD4yCKT3W4Qrcf8QVEh4HV
re0ppUFQuoK0vimE2IATBZaqGK6wjvWZQgLf+4uNPiOhIaGN10JlfKSl5XMeD2ED
Nzsb727Zhy8uBZ0JXObXKzU3NS9VqYW5DKUoYfhMOS2uN37kAvsSTE19uUqseWzu
8IGmiHO+0P+BtqxyicoD1/PxuncdWVuT3FInPBJ7Ec+lu7iDR66FwMucb/AcrwJm
NAzQd/Lgr50oNtbwzt/FQkr6o3r/52YU2xY+bjbI21yepiUVgZE6aV9SwfcJoacC
WdBAfadnLn8nVe/dlUH8b4noA4Dxr7V5uWPO/i8IGkr78CIAU1Qub9Mt50m8Zv4i
3U9hiuseJ+LOzDOj9xFXny5leUYL2G/NkCzuXChBuj4vM2K7kggvEj8dkiaYNBX3
GgEqJ2/WnVdMqn4I3uqdisHCJME+ENB1jzgiCt+zd0pyOfb8rFoK6Ij8qrUEceR9
f/Uc1cPRce/gcOjfl1elcf1ARRqEU6dBO5o6mCYhacUmpai10NXKbQM32DfoPxkS
ICi4KAW+Kz1vrmVh92E9PI+dtpjQG+ckkYmNc3KcO2/hNw9Q/3d8X2R0uajYA42a
TgEg2QizPezoyIk3si9my9olg6CAjhZTkqNYKdfLOc4ij3yOTd7S/IyYl6uEOx95
wmqDsj8Tmchet4/FlxeUepM7uMmOs8LQ6gdTPkWXKj567NZCnvy4/0kYARPXtaOf
qIN623nzRa8rA6ktf+wstk4jQucmQAdcsrNtQaorPRoQRzojOuxnPultOiU3AKDA
6OQ/5uG0I4f0aH5ZmjHSvOcYhGeydgD+5Xhczda+VGxz1BwAyo0lyy+6J9KLXpOO
TXr5OwKbrZdLgew36VEQ7g5gWYD4ki7+qOjm2IoGzqzL22NotDobKBR+0eIoLVK3
8WWB+Z/QUkMH+LYGrI+qrYjq739jjmAAFdHY67dEZTRZHHKhHbG7Kchg4G9cTb1P
azlWwYvVH7YRtqhEVdb0LaY4u/ELALflePS1Axn7BiZUa6eyZjD3tIxSkkdpC42z
E2IIDHD9F8e02K24oMQJzScxLm1xvKDInkFJGPI7L1V1Fwl843hmrLAs88r0npxl
jXTF4clBqqLdoLYE0XH6Z/0A18DeOHGuWghehqtUg5oFGT0PjCaDm4+9tnJ2DtzG
TIjWHsylDth/T2LrdgKn4VTEEpj8WaCv1pZyE8zytiSo9LGVtJKTuhMfVufsk56s
q/UkuEYfq5cj6uLHzptE1UeoXClr4MCsGLVJuBz90tXikhLGDR4cL61gAQjisAa4
ZFmbObneeloTmY5UQciJlEp6T1+1zdVjh++IlxL2up8fgET8tg3O1ujpMnX972ry
iOMpw55HgI/C/fDv0I/ldM6Y0WBelKPWGcZ/vUwSWo/sM3qRwljrv/dRCF4Bh4xZ
7ES9I/PZ085dSOJd0lnKfs1gDwW0ult9X9tgDiOnOGbE5XnzF7O4T7t9UWKIo7Vx
AtZjMZxadPjCxCXsalMFvDWQuqi2u2/IWDbnNLZqbEolNSXmIWh4dlmlRdu2lVyy
4p7pvCRvWp8af35pKLeoL+7ugmj7afdGG+Ow2rybgSuM2q4J8SPlluiKCST0k5nw
x0sYhqgdqd4tPMsEe9yh87Km/twCxXO9/ud/k2tV8YRWBDGkFta+zgReOIp+547L
no+WPe/k6JFz06m2rSA+uNLlVor9YXt/blyaKyWL7h7f4bo6smKexMEbtXtVhL9O
XMfdffY+p72uFd/GOiW4n77gPViz6T86Ls8vTj+bREBcrxLwZ0yfb01kGSOdTzAr
mfpTsovHpe6yvFftzFRosLVEMD8M2Sk35R2M9ZUFWZY9tuJordLPgehEs1F0jNcf
ae4TD1619ti9VLvu5Z9n74Jk6mp0u+BammFtLLn/D0zG4FJr2S0YgV8t2uVcWGG5
IHq2VDUkG6ovBKGIMBBY1i6KCg/pGamj05eddW3Qy1F7XqxAFhbpqJaDCHj9xliD
l5aywNDR5nC22D92R/OOgC/fZM5aFpchnDkyBPst1ESeQZi2wPY6YdQHdoEkiJfP
zxVNGDzBjtJDMWtpZL6gbF/UODejSAjRKuUgmmLAuGSVPwj08Bhy8Bz+KVRqHB9w
YG49QJAFCTjaHinfBOVQFM/jsCiCQuM/PHDMlez4qf0OAEougxJIjysC8DPbF9yd
jbVuDcgFcrUlnYnSQkLNuxbnlAEE/0zL+mINxEJpj8PzA7dJUdooOkMUUGD3gKFN
Q0t4HQ7k9ql5Y96gkNwX8wrWi01xyuJAZBp+2pDF055DmL7LI/qivTpsHszxhLL+
VZVT/iYNi11Km1qgSF3hpqSaQ44Brbt5JFftza0cKMk1kn7MOF0UCGvQkfjwFOP5
mVqD66DKbS+QXfWDfL0qBEhDLGUg7CkY23/VufE/NYQx4pDQ05whbhIVmCkHG03T
SFC8M9hxh+CwwF8kVNV2zcmPaw5cqIrH219IufCO7v5L4teOhbJ+bv9TC72yuGKD
PyMqj/hL3GExzMbQJOc43ffN/EKivi+8efzNnRckXfnviniidwsws+XN4OytEnR0
YumsHhuP7hFZmzEpYNZ16rSS9DoKTE/AD6D00cc8G7c6l4ELNjkduWLlKFTH1Rze
R+Xl7b2KMbnI3c6nPn1TjDZBn3MW4qKMN3kWBDdcZv+9oH6pef1ekW8kgtgiUNYm
WHyWhKNjppmkErRAj/eApjVOhnRTHBsbNnZIkflU+nCRcm7ze2Y0YEn0d3WWN4Xj
k7ZntOthw4Dc2KNt4/VVUu7N0IG9bU4sw4fWT25KkNUcivdYe7Utv9YWjTqS8Fa1
/JU5QsuQz6zrcIgNPdPQ+qYSA/UqTSrIrSDbAVQ940cDay/7EVjO6QID++Be18q7
1dDB9LHxw8z4UEob4pgXe03L9XLh1FQinSbxEVi2Y38sEViYb4knIMBE2TesJDYn
rOOApkz5+dza9EtTZa1Uh0OqCwELfXre4oq5Yjflm0U4o4zKqcmfL/yMSHhJVn+R
4JlfdO4fdYlbGIgDwsvTVD51sIVattbptNFGhG0B1lT5q1Tre6R7xqF8BiKMRqhz
tUfOxZGlkSRSHpzMVXN/WLjTCOG/0EiBkGf5Xm7lHBi77KhM4yl83SUffG5VaN7m
x0L2ya/aXA0k9PI0hxL5a7LHoyBaioZOShU9g5oqkSMF5Ou6mUnB8aGDd9AxUz2Z
e3aZU2F3uM2xOWM7pDzYttnGvNCMJP3u9VU57l+PXPTwWq6VezhsWPkJC0KlxdCG
fujr3JTu5XuIpPZolzB8MTHPJqaUlzzA/xzHunpt8sQyyWOFKFrKy+j6KZ/YQ8lQ
euX6+/cVwkc3AIyEQuS3klc6qJndLoSp30609a1gLtuINU/91wFN/jQmLz0vF+8g
9ro9R1WAaw+t40lFo5w3DLhmLMbmCHmHQCNJk5cOkY8Z82ZftoO+jv0DZiuQSztt
0KlUnnD2LiBQ1AUW5PaDV8AQ1pzRQo1dfMDQu/E8oszJX8Ij/0P1hF77t81nhXie
YMsv4VY7W1JsRyTRMEBrjJ7rEfblKJbpyZY4UE1nRJEEC5hJFin7VIwlz/WP3hAF
LBNoxPLB2i+Fn+OHWW1bEu9Wkwb7wysFGLqTSX/I6zp63ujZmFJL8EGmI5/jwDj6
t7l5cEpFTMAeXIcx9mrZHBAadRaVZCnjF092Ai/WWJ0yrdbK2XNtoLakgZQYmHfT
NqZPzawpgAG7FxMaz5yL5U88RC+aes0uvfbL2esxGOB0skmDbuWdbeoLeI58ExZu
Vx9GmwaJJ55oSIOoIZ6i32zF4djmGOmfr2WZj5s9j7RRkwr5QG0zS9ubhVK+Yjji
waJA44cCexsZhbe6s38cy4DHLBEsVOaWmRkhnSEuACp99/jhMynwOOuPzinYaGo1
ItvZEYYHrQJZzF9xZT3/x4Rb7ZBOlktbHbL9xcTQdqS0ptygvvrOL0XzQKfYB3iC
mhezP+RZEz9/BgIL0M+FZGWbuS7J4aXb9alR3y26uE75XxekNTvqgAG6HENvRWqt
AMYEc0MsYETw3PPxal9FE8exoJj4BvEpNz5/V2xgMSaH0gtmwcA7bGo4Cc08ivhG
EF2PIktZ8phi/3IZbLw8NS+QquusqzJ0onODgpBee4ez5++wKJQZ3LSFVNzL/DMB
Cp4wES4I/VLXLwFszaQRl+wg4i9qTRcvieSqsLuFjxSanlDPgAx98MKI8c/vlfTQ
phxbSlztIVXrToUW3L6ZFoZ19UwJWEKWhG33JpVjxr8oNWDJk2TuZLQFteP56vNY
2XDv4t5TS1FAHw5gLg09oXsdLiPg0VhbcVknrbAvokaUgoSdB2bSoUJPOoJ7yDBA
0utR28z1hmX1PPqxwO2cOXLFP019w8ht+I9pfXlBks9eVA4D/oi1LRUmfi5+D75D
4jsna9mtQ6yLB0qgNv0syLSLgT0OVQMvFeMENhH7AeW7sFblN/hoCOJ5uo1zRXu8
InFEa4uJm07r0urI8GwJKp2QCXFRbM5rxMdWtLaLiPaGpOfhCh4RQBAyJnoEtgsp
I8bYIts1HDFdxEoeIyc9ZecC6ZU46vBMc96Hkz32XIzEa3dZEb0EqAMGSc3MN0Cw
8s+wAnxyxEGPoANsurXcxy3oRJn/YdsZZGaHpV0Wwt8v25ytQtDhsUlAWDYfYlkF
HOem28ykNo/tpnFPZoJ2f3O7sj7JtorBmqPlJw06NOI7p2qTMQI9iVz68AYPrDF+
2u2NOFBRjjPFLXxRLdl3wr2qww1ppaUZZ+dQmgc5Vf88rtf4iS6kD/uPs8NeD51G
TLQb3i8ao6//6Lra0/XWvei7n8P/b15epsABULi8R10Weag/j283dw6o+k4rUMFt
8pKpu5mrGwsKrNriG4+lPDZOZgw52MBRsWJqLiH1kgqtx3Whis89Q9KgpFu6Gjvh
NtO69PeevYBOc11m/j2eISwQfBm6eCMjuAgWM+jHaW4R+3wrAAdSq1fXUBhEvxwB
ex1Fuy76ABzuoQ+Go+xX3CJeNqhBbIQKlxgZW9s0MUHCv6c4FwG52iWrfGkp92bJ
hyUT630HtfXaD//MSPCGlAVMv2DwYYTfa5zeQm+MJHrzTLmyzoHE0yaFBsXB4Rje
7ECqo3ZOYx7FxBLBr6eMzre+nCZEdoaPy2IUcn0PgLYeDkFROf+2Y76a1wcz1Ptt
0iXfQqJi789iZQPwBXdI6k2ZHDWALgKLZCdspN8bmUrgotwe4oO3hLItXJaVFMr8
iGVsDG6C9jnjGQyHH0gMHrhV64sc6WHka1PGFnHuxkH11BL+XOh5kOx2IoxXolMd
O9BfG+9sMu5aUi07+3I1sKTB9/0nbIWiEfBriSVA7WcmQp1ED5aHLa27eo6fjvTT
v7msiZryiOiaAQIIRelHBHn31GRAlLnhOV5IRE7zQez1snxXihZPunrNyKkQMQ8I
VD4iM5LcI1Ysw+n3Y6GybM5l1wE3oRDxD6AJSnDDLsGvdiBSu9yMSLkNj+GUsE48
XJiTARJeXR0tZ4/3B3ZLR0nFd0mK2VMw72yKlmCDYdlN6WqJrni2dZubz/sp/Ynv
Ggdp2TE5r0ap0plo0L4vBzDOh+jHNqqV+H3S1IDsKTsu8lo42PH9RS38/DjvEvA2
VXh5il5nTevml0agAkKJA1SiRRfL5ir7s2HC9oDbr379CDv6V71EaWGeXfXBSzm0
zKXynGIVVZLvAcobe418/1RTu7wN1p9bOKCJ6EZUuYbZ19emo+FkZTsUBQ/+lHWZ
shS/FxntPDji80QF3fjhl2MVImGhJMCOLmydvYM59SPKpISlLqOw9ZxB9AztNeuq
yGL4PCnC5SxFu/u1R4Aw/rG4JLdi9ECYAKP6fB1zU1ajV9aswsNVEYKcD6qPmj2j
NZVBfYDK1/FmKAhOw3AKTYkaJsb2aQfHxkRh/CMB9oan43SYO+DrkjKj0wmZzL1U
fzADJCn7kaiKJVs9XQjf2cNaervKN+1476LfQVnjjj47kZH7ujmtqkuJZz+3ILEl
4d9I6PHoj4KyiwEw+sBlHXv+1ESWT2GK7I9J6mevBIJk1Vk5HMv0tqGLPbEKaUAT
X868gwlt5Ba8Wz5t6/9zLsr2JQ7f95E1qa6F/zpqa68PhMKgGVp6lwVdRAq8H8b4
ZxByI7cKQeWFG+nAQP46TQ58Lk2KT3vVXHkjHBHuDkY80JWjeoMNcY+yJHgnEcoT
GPNLNYzrzxP9QMys6THC01z24IM7Qjsvylc5Wj5dA3TTThRI6F8IfQdVLM8wb17s
SurWsyBycGMEYftwopQ7cSwMMWyQLok2uAGH0/63U4NrQa8xEv/4yc23pfCQR/xF
pN3L2qpQ8ezwoyO1mEBgnVjFUr4JG16faOogi8/fRGqb7r+8TgupjnK9bENMCmph
GYXk+ML6u7QvO0H/fHCKRjnZFKvaTC8p6d+rzkxmACWmkYMYMH7gsCl4ywDWHUJD
qohhb+ixLe22Ojr8vcW9GLnZ5mcdJdPE67OO6eIEdlLzt/DUTgaPhhZMVihAVEZO
6zsqXUuCnziLo60u+QcT5ikUu8MvqwKyPp/O7ID8bgz8UR2kMyyxMFW/LFvlRlqM
UMuI78XwHwMX+kbm1r5g2q0XKdkOau99zGNdGnnoqD/EVfzedQmS44FGnHMcczvH
93Q23/vNLAjOYVvYxrGEB58utIirGIY+jC0eN/4C25hftkfYzwc2pxj02tu05xcN
Wc7931Rcu+Ivz5ovPjTb2BEb5rqZWdlVKOpGm5qjQuXn05DsdQoEwA3156PwNBMs
TG6aLptUqbMX2CqPO15rlB8lN/XDYIlouSrYh/gwZljCazYS1a9G3bTOUheAV6g8
2AcuNuWQamgVhe02wgjZYDzrWqv26y/Pf9DckcNF1MwRKFEwu0nuyof7HEE1BlQA
48TCsj9JpkDdaA9ajh1mVZUK/CT3WGIWLhfuMuaeQIW7KPrl7iFsYMRZfrFXGgG8
6GswSa7cS8r+f3bAueulWQ8tnbGzHRP6z789f1L9hHs2OGg3+HaQkXqUQ9XihWBH
ZmBlizaJu8KcP3IFkKUMFcwtwu8iNsjTry+5a1SPeBaikOXSPrCF8bpImqh/5/dK
vQJafJ74QbevJkVu4iK8d2GSqGX/6DxS/qlqBMtBZQ6i4EBDwuk6fgyp/KBdPZ58
JTFh2Jrh/dYqi9YOq0y5TtyXmUBkcTWf7bxNAjM1pSYPPTF0zhRCtxYtOn9M1SA2
bc7v/Q8c1mtXnMXY8PE4/n18hGRqpsBQPfFbzqK+QyO+PJpz9e8c2KMS7nyHkt28
rf3MfVBFoHVg+Fpppfq40LgomdPA4SLDc9DgVm7nC3LYkxZ6ySQBIIMTKq8FVoCH
Co1eHGNGfoAZWdCi/QHvvZpq0em+CoBfSbgleqE3qvXUWFTEmSqyDkoUudoiRb5U
k2kxOCZ68AtUo/dZ1A13FPXygdvG+wZG8OwuIpwHA36WYPafQJZ5Pci7IeUEI1Hm
Zjdy+ZUlliW1O+7Pdg6n328Ht56MKPh2RzZgJqFubKoZ0MTEnUmUbd7c5uStklBb
kZkQgeTYNsIT3l5/gw7FAMEoFBUIGMg5a/9enwb2nc2Q6l+v+bMiifVj9GqmW9et
t3xLkIiKv0PvO3H0NeOg3qQ81rffy3nUNQNX3UxTADq07wXcmjw75X2Fu6Nd8zxA
x7IeK8FFxN79tcduHLE543mNW7wjLb2ZR/NSW0Nh7gz+417xF31WM/7Tj/7GZhOJ
cj+eMUzGBkvPdvYle8GzaojF3+xvRkPIR18PBVRy9e0AvQZ9eF8fx8lAdYxuHO6x
Pfsm2wSdqy6RxyEPd/6fYQnF9488EOvUPKv1u4pEOtilvuLlyD94UEkqLgkI6W/+
gaR88fvfzSLwhOp7g+KlHRd0WdJbnxakw2BMNZqiyqn87pdHWVITuzfozz1bc2MF
rG9zFCdpQUTqwlJT9OJ6kJeG9vUNx9pv/MoeUw6706v8KaZjZ393Elt9kiVMUOtz
TVU+ejLY5nGH4IOpjNrXJDsVrEAO31BgHsQjjNmAP5gWDzLD8N+hNLgSjWS3fqqD
JHhIXBetKVuMOGG77/7o5AmEAn5oFI6/Tox6Ww/HiUSxxROHFZOUZLIW03jN34xE
DOFU6XgW+B/FjxN97pih6fzl7q7rRtKEnlEqkVsHm+Y07QUYoAABUsqlLkbvoj6B
i11N5j9O9MUBj9+Fw6H0mv7IaybfVVWwfeOcxkdmPudKNyynUifTRQbmULjQKWLP
TaZu9W96q7kaWWRyCyroMgrGtJrmzZSJLzbe+9iQlAAUX3LXv78F1rqSJgI4q/V6
luEv+fF2K1lRiecIawaBQf3F8s53S5UkBfmHePCJ2zYjGAxbRo4Do0w66qew6TGm
lOUv/SJncZbAA+tVYxnksHSRpcUmESt7yE9sqQLSRgvZm5Wi05rf5tEoaBA2npe7
QewSztR1mMwYPDaXW8oXaaniPp9WoFs/0ERyTak5d4qmv30iXCyumkdGMaQ5eHOQ
Tfpkd80+7nMZlpDbDq1G/jax9qmWJ4pCb57g2vErVtTPvJBTL+gtGHoaA1KZnED4
fxwB7S/WZ2Iql6ZJf8zI9Wfvqxz3wPa3pqgh4mhzit88WXl/qJbZe9AgP40v0T48
Ov51peAw99hKiSLAY6GRIX+GE/JRuuCussGbUNR/eoYt//eO7KXcAhRChODdDRI1
xRoUbaA9AWVn+wZm1Z84kcZRi7w46BkNXtm2aFuMsINGdijFCb9n5R7a5gc9MLWv
ESnucypPWODbUzexBI5ZJOZgq9pkCWYnyC9BAJYvhBOEy3P+EiyopMZCrzYAz3nl
lC0oYPOCg+717M4zALA4GDs8NQADTlU8GGQwsQ5WKbRj69K4stZBBQ9A+XlI/OBt
dS5vZr5NB3/oFdnncQQZf0W1QVGmWdqPet3nj1xBeJff92kRYbKUpWpcVKGiYLI+
ERkKMnSzpAjeQJhTL+EMW15O+ufZmn7VjEMgwVhb7Ex3NN/5LlJXL1WMYYj0XFMZ
dXjrCQcLelF59NwZ0XqNXlDAweo/gVFuY5xAqpJ+p4SIXuOdBDXutcxXzEQnxD0j
dmt3CnCFU4rjlre/qzlRY7LsOu/0G06wvXg7RzXTsIApAppWmVu2Z3nzkRHKfZ5I
miPM7MiddSMZgJUT98hviUgGIdtR1mfWJ9AG6N9ZgCdvSKQTVs/Hs320NxBopjDL
80R3RTAUwavPH0cU+JG1M6Vl8dJUfhxp5i7BL8yddO7W4J0ss0DeQMEiPeSQGUtZ
ZlxlZWlU0+8Vw0RwU4YAH5MIyKchxs06FH0dnUKD/k61HqnJiw1BQN1jzOSvMEqT
Ji51UM3XFrhQkv2Xt20okiSP0PFDteILBFGFVi/d7XFfo9oVoKTUowrzJCsFhBTz
gpmSLqe9hFo3D9STQ9rtuquX/FelRq0ymEtai/Sx9EadVN4C1Sv/z7VBNej5ObbO
UrqmgSUGvn2EFyBKQ14Oxluqoa7N8hspACfIHfRvis4CwM1JAcrnrM5REAoHGP89
7BYNojB8dMAAIJTMpvqH3OTc0FjRYOooF34tYDVc5nPDHf/omEswm8rESLNch+Fa
61fehU0ZjNh5jnxpRP7pfXkGYbddcj8vIiDrsKiBgVJQqOC78iaNC+l5HQ22q/Of
RMeluIVUT419GNS3yym2Ddy9mQdDjlb/VAPZqgr6GawRxP8JuIaoLHH+lFicIet9
uifXofCzZBmSk2gUULNcPqURyzCwA0BxbTZ8xuvBVd7VNXh2QxhDvskjSKRgWc/d
k6kIOKuA1iOE8Q1GqeFexQocM93m1IbXJyORbW0R5ly6vQqDjPuyJE6FFFLaOPZZ
tVD8BU+RoifM2sxvTWyIPOoHFTvFn9YRrhMeB0lqTjePwQ/lDFQ+G2IXGOa6jxVy
xdDSU50PnPVFzUks5oFQoQuE/wUK9ty2KJtDXT0wRaBj50/quBLqtAW2YjvkpNDg
eZ8D1KXy0VHUFp040HZKomvf+ZDOLx2NQPgh3Jve7MrVRRu8HjahlzyOf/yXkg7e
CerK5emTZch/lyZQvRsz5fFs2qhnqTprkPMBxeWss0Q+rvfeH3Js5KABt4NgCrm3
9Gvi5NoaYPPrfGyIUrcfjPosljYlBLxwajqj1oWAhVa7C8mkBBF3wOffU5NPOdmT
b/rivv8FRHED99rG+2HYm2mOy1By8TwPxr93M1DsSfJCmz0oFpcb5WKz8JZJeyg1
LkJ5PPdD3hN5zkW2aY/9D4rOjiHm+NchP5hw6ZxHVGUjcDXIQSa8Kc6fuCggjD4x
YMdlylEAlNETbjiFOq+VUdTwWgpYt4nk4zFHNNxyw0c/srCC3OmDUy5SgcOhyBe+
8YtzOXArV1e4CZAS7fxAuwtj3iq3usCrT9HbQBku2xNXQi5+61HaUnGYcJ3P+hw9
6ZI8QhNbAcJIA8S5SiGwvjFTgo65+uYaoRM2bNyqjqIcYOOoGF/sLqW0pdhCW4jo
DFpUAL/j3wsR9JrbFot2HF5jU7arO4piKYOFAafXyoHubj/weypPZKaS/mW9Svr/
uxDEYElDrujQxj3wNYjTJYt3tbg8x+fPavnM5Gc8h1s1xSnfUYjl/GToGubhqjxS
6bCNoujIl0foVHIBuVReiZuXBLYE8fMXPRlu06Cb0PXkneu0jVSCX3MKL7vcIulD
LbrC3dqhI3e+IKO77tq3U5S+pMM95DP4dIpXVFixidldIJwqeOiRTo61B1j4JUGM
WF1zn+m+rbMfOxuEQ2BOE69j8eHjw1iiOOS5G0ZEFQjZNZ5fzG/bp+NeTXmSNnbc
8zydjt5PB6L/jyWr7ZK4oKoYOVoB13fzYY1La/VhfX+BnIAIEE0sDT/eZ4HLXZ+I
ZbLiXWhTMEg4Y16OQisXOZulSabugCD3D2Pbib5RVLoBHtdvJfKA1MgjsoE67cLI
RDObBDj9IeQOysUvxL7q5feR0wo3WRE2Z30eIvzzu7Ni6vSalrGEv1n166pJd0ZQ
HDRjsqji7Aza82CdmYXxBgVymS1u0dWRaZ9k2OTsMv7yH2kWlXLZZWoXTJHQFv4p
MZ8QeZG99XI48WBwxLPEky6XJqKhEdIuuRkHNwX7X3SU0KlRqhw45QD8r8Z6cT8F
Q5zvsFpSlUeBp/pNlTMzxJIpXPwMvoDFgcmyar2A17d1Uv8chIhkd+Mjg8ZRfSJY
QsypUntMksWB8r8GOs3vOuDCH0+VN2yIYlxLPM5CD+N5oeTpTEdRP/74euVDwUP+
v9cpP0BOeaAZiH1AmCPbHcMonuHRUpx3EBJNu+j7w3UTHojCCplF7LjFZL3N6B0W
EzuGnUqWZFoIqipKxjEwWJ1wiGn/zOce9W765wIMhElx8HlZNCeOOKkIigKmsZL6
WvuK5qOE/2VwrtisSZ3Zcm9ds4l3aN8+pc7hIe1tOuKKglfavfMYZoS6sf8TUIRR
K1zCyA/65KFuMUDZEcBK02F77HzVwboriiVRL7hiqW6psbF3HUn1D+OstfkxgxSO
riwAJ5vELdW5CY3Wi12v3CXoPi5qnoqjQT6jIxjMs9Qcxyc4eN5YuOmKHJPXl38h
6CY3SLfmhpmhujjXjOgeYm2Vo4YwntKq0OHbEVblYuLPgUadI/OiHLV31nUiFRxC
VUUoXC4cLXVuk4soN35id7I/MQjuXQCXGvvAysaAUhRRvMZvm6ejZkjvbgdRY4sU
q1ifmBuuFeLp8cLhe8QLSQCGwGPhG9f6qYXy73i2Uh3yZvq7OZcCqMCKwPLMgYhL
wknuJyu9bA3eNcwaxFBY9GZTnL0nZdB/MH7foSf6dGksgfeV2qm7lNAWuODEtsGK
ekrNcHa3z8B6IqrdfKWpbb2UaihfQXqBTASgRoX2izYP0eFT2kZO+UL2+thlGoJL
bGws+KzPSN0zCnd8NFvvzSyqjKx3xXBzjg79tbSQ12QHp3XHawp35QYVUhpFvWjW
Z4AwICcKldF5uGVw7tRjjv3jerAHQa3WqyvqHHDpXidiYZ7YGot7RdNlHfwP3m0H
zHXvLZ5KTuHUvkzx6DuK/aN36pB0XfLiS/fda03iHBqPTx/awXalv7bPbNlU+YgB
VQ5XO90A42p3wjRklOkor6IjsxO5g0Iti1+CIS8c8H6Ub4j7u+R6bGwLQI0xMcM4
CZZlVXvAUhyq3Uydn71c3J2pNlRIgKctuWBoXZDPpXoyW1DCThZMgszg5hig3ejm
x2teB3ntAHcKfY7a5PuN7jwNzamHpuOktcTkDeCCFLIhZuwS8qM40+xJLfGXRi+y
zHwVLrK8t8OLkrNuMi68fgcDvJnJl+SDpYIdjf/ydcRqGifI2IgyvlQNp+0MZeCJ
xzI9iePm/jp6H3WV1bZvuGxmjR+OUmt5OsmQa72fFfDg7ujcBMYN3513l+MCVVtu
ZoBFKECkl/KA4glQx4i3bct1jr2W8rv35tdc92bRMUbor/RqA3D79V+Y8m7BD2/t
k7DeqHC/Mj0ZzrKHir9eilw0koHgO2CIjAiLKXf2JVGYDY7huf9jldoHZjpucEDk
9TTm7FLNmBeM4BpPLJHUAvqdYBRzVNp2Nn4EMFxfyoTQEx12dJoDETkzi20laz1n
a+sQXECyHb4ZBegW3u8hwyZiB96vy2UcqFs64bRh6jv8u2MoEZ/1ZXudnxBhYAi5
S10jJ+UcF1czJzbK67Ck8SaPjlfs7SMq+XHqPOYzG/JuQrD1deE8AjA2p27ZKNwd
Miue3iepnZA1/JUdRZQOFOT/d6iOKSdkBD5LnERl/lLSsOXLq+6XMtciBw1LSpua
RIN2A9S4Sp+xVcPlGPxSInt24xTMiv95UMXP1oAJFu16qU7lWucd7u1YXpP4PwVM
fGxHCrrJPUgGwANEGbReS1+wjYIChgUMhpM2RLGuUXCCh3n65z+T5+sPU8fpon/w
x8pyxosWjjFfo+PCTuJjHmcS2ajGedWXwfaf3Q/iX1OjPbTCFZj9f7b81Ak1XDMn
QrGiTACyurC01Yoq3CPeOOWHxQUzeEyBsV0DJlo8Lnwj00Ed0c5swjz4h14aZuMP
pziy1/GNXjhgDjTTkmE+ldfdu9khewr9cE4SnlLedrGH2mm08LgMlLUQozwF2L+M
AFvEL4U9QE7OQMhRMbD0B4AD6VJDKpK7O0pzrLVVMNAb03GnIVbLBTmDrFkpSYoC
pZckJivlkM1/o+KTZy0+KPAVGL93ktxGSSVjqglkpToAKXTwXGWmkEnjK9oL0gPV
qrUddwnjdCygwB2gU91Lj2aFD2VyHRRvbJN7/vApBcmg00llcI57OB/NhBkWtLwN
GCg+G37ZlHmpoNCuTQEHwVeDOlw7lNlv+BFT4iMF1Bkh7gFSGECiPropKOzhWDsL
PS4DBw71BCaVOJOsSES9x8SMKAK3cF5L/ovmuxkxAAvsovprtj4K9WXCInQR0hZD
W0osSUGEdLu+566VtmX/rXl+x8m5wl9HvuJIjsz/XXfLIXwMhqiP99Cz9TZhN4dR
nEGrclo2Z6crCcmS+btOnquWW+ucLoUzZxoNVfOTA3yWLYf49vBmi/5T+WmJ6v0P
RM+NKOqeGgMz+bz2ZuI+/xLTpiXhlYp1Io6Okl/SgJtJ4Aul2MKDGnSHT1BWq+7y
okU21m4BaybwEFWTsMpHupLVp8stNrOz6uRzawAVWYNH3FFft4mVHWWBvlmj6yZb
2Ren3mhsLPlqIPB8smRi9RPftlwweJcz0Maz1NK0DvgfwvCSDmADsY6R2/BTIyXE
CKl6qW7NBzJVTmR3Por+XVisDeRuXpqoZDOo0k7Z7urQb5QdfjWk1eQPe0apQImT
erNCdZlxxjO1pYdetSsWI4Q0vrrZQwDzb/rvAGe1cz7RaUWfYtTRLh06puJTEhll
utxwvtNgUi7VAhSkPgslTWkaDCRkRUoW/9z7zZ329krR9goEzwcr5QH98V1LqO4w
y9swQUC7zx7liDN4MMmyXMPerv7XPdKsNpv8YL0T9YvKneqtpj0hIyHX/6msB/OS
7nLNu0P0MhC7NzKiljuciKvCrp8XAAg2opIZIZLeKaeYqr50fC1MYIrDt0LAhrWl
OeRQJA2ME9LEdGeXghMCdcu6u59sgagTmE+rZq2WMXZcnkJRwDoMaVyjzl6lqVxJ
S6o0nqLS8ZcWGksjD3NBXAoMv2aqENF5iurNo7QXp10GSfmZ7F07yw5uT6fn+6ZH
uMChXzE8OVPr0B9dE2/hA43o0eXrEDVKJiUVTqmfJTurvdZwSbQP2qNjnUCvuOPg
YzFJhwB7OhZzMQ3iWtpoKU8lHQbNcamtIf53LW+/zL96P390XmM79VNgUeFAN/DK
yZDAA90DDdMYhiMN90FofDVA+/xwCijVfdeNQqSrZlI8Ilo3/6lQqjT9fgT96Red
s/QJvrIB7rBZBBcdeTxC+wRxTj4KJ65VECH1TyxGSxQyr/pg7kiCwp+aqwccTj7h
IGsitvrjZg+fsg7RsqQISPAqRLb2d65qcgmBSeSSQ7ZM8nKMOyzTyfiB95f8EGUV
mTi2wO6KlGUY15cZ9a7Xxa9cVdg2XkTlimPhHUy+bX7Ij+Awp9hGSNjTQ4/fWiGy
4imBuhNMvdYFBnrnNEIkNZ29Kr8mzoi8fe1NdS48Qxl0VE2h43l8JFbYolwb+bUL
H36KyLJe6xbapHQQ2zzZKBKVM65aWesAQgwZ4xS/Qyy5AZtCfUk4c6t1Miokkl2V
8L8FPpm+U44Z+zZGbo8mrUSmSDM342omuqkW4LtXIGHytjptQsu7RDGJ8uTv1Urc
AVLfkro5MTVSzAY/HoMfg/XLm8c2xlFzsx1iyYh6EqSsj4DXNdO/F7zwJCA2e5cq
Mj7OECDh+N6EVmuUYHSGmaMEgZebFPd24qF8L3nSIxAJXIo72mZZ8WzVXmfJk3aL
Uih6HxMOJuk1HhV48IgqzEiLiI7DAOBnV4jZG+cirGzKw5rYUn+c+cjuFc2VUbpX
/AV5njaT9Hs71kCQfq+uhaJQ9OE8/Btgh+vM/bY7bRqOvADsYLlaYezzlwtiY8Af
9vbQAWfKCUzNdkwlSH763Pr+4ROmL3OZvfp6URMiuB7QTGXObjUa7LUv0ZLzW7LT
YvcETGUbgfd1IHh9e+Zy3T9wNlFaarHlbQ6Fjy6b3Pzoc8RDf4kmGtrXVj3aEokx
ryRquxTEO+X0CGh9TJIkueit9o92lwaO3iKRzFOdnTlLcgiyHVoDoicWQ6HjOORm
DszBp/Z0cNp1qOgpaSZLOx556Nwr4vnyUVaipA1RxF33pGuEbaeUjlUNA3jBZ/8O
tvqX8YJ8M2wU/HlXxc8ecLA46oHk1aFoH8X7qvG94shecm51bokQY5TZfDDAtR+u
BFsPn7/9f97nktQPz513sg214CyIsw2fiLMH7JLsE03NqvitQI3EyPz6+CoxgDeI
flvgvvZKWPndjnbO1rkk/Q+AQypcGG1BHy6bPIyJhqgWHFaGrF0PmeaxZ5TjmJyO
lf3U33Hpi6D2WSDZZXhwaxMHkst6E7BwZVe+0po4tGYzI8oWQ2X5YcUk/UzDjE0I
7KvPUncGwoHppL0h5m3BdH9AC+j5ULga16ygBbzX9lGyOYrRqA8ccpSf1H+KXMA7
BGX7WjSHPUth7IbgqJ2reSd6tlgMoAaz9VazS4TkFE7p5Ih+zgZRJn5Z7qWx8ddW
OogB0ntPycp4ZQHkjxEl5WjDlCEz6PzvVcz1Y1j1eS1gB2r7L3Z7auz/4khwMgg0
kFOz2IzZHV6FbQzvi5grgrp73Zn7pOXPtcrlEhu3nTVJG2TfCNSMW3Av6lp7EYdQ
kZrpmSwMO99etfz4HFmWe+Qpc81pihgB3qCJ6frENGoQMGIKnGLjtXr65KtYWv6U
rST8HVZzEIIjNkW+i9VXsomBpCaS2m0WH1exLUef5DKOFL0gsPPhWCiYaNFswVwE
iyq4Ts88gDasIDHpL/Fs/knTmpRdR0T4LsaRZ73ZO3/kQ+405zHmfguX8B007HUz
cBp7ZdC3ptnDT6f3HFucxed6pJcuwsybaHe6edoHhw1IQw5wFigL60UvuoEoMW9K
4KKi/Nn62CKSYh6r5wSIP+LthsCRSOiUXMKlnAz5K78P5LeBfLLJMPakZZ1QvMro
610bYDHL5GDY9BqBF+rJv49R8QxhvLF7VXifAZm5/Wu1FkgewYeWlO9qIZ9HONqy
qaFDCayk0nXDUQYX8VCzO+m7tl+Q02D3aIUoc/InTxuUGy5zM9TBz4rUjXoINf/q
8F2wgYR0pmtNN8Z/7s4KBwBl7VMH3PGoQUHarAh/nc80ClJ08ADN38u+1WOk/M/J
BRC+TvbHOuVaIVLfPM1yB++OyW1BaWJYhCeyqq6F0Tjs0+dyPF6cikmjvjermxTj
feUC3OEdGas/7xZ7YIvQMfgr+C9ZEALhC/36EUxHPzTUATdDHExmKDUnFwh2F+iB
JGprDuHyaJo/Zh19pEGS8ZSEhecwkjMStBo5fF1PVGdg41deoL+buIMQlxNLEp7k
eSkdt7UbowdAXJNx/f7gq63dmOtNNmzN1e4hfn6JH9Pz377vZ8jVVNXbeoWzvkaf
Acsmp2rkQO/aa5M71eJd5kemv0my8NCpPHYEh2cmKZFhQZPbVa3lZmerr7HB2D+7
4dyBvV6j08jPbU5UISHtkRsdy9JBdNp8+hJPSbp6naESMpwqVGUBrc51su12gsR4
0fBsoVEB0dChYUefkjoNIKrIXNMKQua63kW3u37Uqm3K0ztsj67Oa/DlXtEPLelc
kYTkaBhFNV9YGPlAkL3++bZESjfAthst8KjvnJ3c2Ibn5Qv7kBM4bqIPaynep32W
M5NICa6DYajLyz5qw+jqZThMjNXE8mryPKs6VQb0LluJTzctBoSPbANU3qph8dbj
ZCYJfCrNFwue99toS1ENXsPZdJ7WyAoonjaOirDnwgNlt1ONSL8LTIKvsN7S0jYN
FDRmqUpdZ68+Xk4JwTuf1PiW6Xd7SbAxqQ+ZcWu9xqa/lQhCYHn5yGD2fc8IMUVB
ZKBZihyGdIgfJqGllekB282xm+4voHHJ3jisJ29+Eg8XDrDTC+wE2d9UzWP27wPo
1cBqHUXGBfBL90vL9av63pxx3f94n5mKhqvMYqQt0MtDkLe2NkFzvijm6x5qxy+Q
irvU7Nii6StZy1tjpdlTISva6c9vQP0T8agDx7gYKfH6qrPe5ssrndFl0ca5peUB
UrXZ8zxi0GVbo36Wm3EgyPOjXSymCJSAy88hZcDsDg+qxAMoUz9paxFFZK3PD34J
ylKuZ4VhsstufY2kkD8vfjdrYx30R0ZoXqRHJDUVL8Gcr4PJKlBIKrhvITuqwjcj
GxbLjYY9cYxYB+/uWGhuZRbYHTthElGswLLT6yU+4I8n+JSNM+G6pQ2Anmbc5AF7
/fbwXixwbvr/7ntu3ZF2nlJPcdk/a2gjFBjMF08fC3+hMEE/XbtMURRheSkdnpeD
D2r2V6L+B6IiS+rM9mNfwGYyxV1KHI0rjwq6s7ieh84FTlCCIs+OYGyT789LTUcc
1hCq0XmBC57nkU8FcyI67AdryzDckh+ROXO77W1snvA+sWhy/Fm7M0ZSYDvkxRoV
4VfYdn21oQ0J9IKzLA5hrp53KxjDhsK43g4SgkRVx7/UeM1sw9Z3pd0u9YBuFtBH
pwtDB+Ur2dP3m82j1hVeu/4IbKxmj72QAzbMTHJGJcxNo054EtQ3HBdIVjRYVGth
pmk97CFqo40WdHYKghIm2BjiGZD7qP8onWb02P2lMhKc6XJsENMQq6H/s6++YQ6r
GwKM95xavUEChkS6nr1LB7aGBNPNeqoPil47wG+QAULQ2rzPAsHfCweu4QdMTlDp
P0vyEAQPgsajaDpPxAw0fDj4pjqEt+YPe8WAhq/oED4za22wQvT++Z+6PtpvFWOS
87RbUhMxWo68a5I2xifT1a2ahQ+cnj3x18xHU/P+1dMustu7K24viXxAt0lKhEs0
YcQog+MF2gPD46ku80kwxXfVzckA69qqRUKGV/y/6YTOkSp5y5Csqg+1LdSvkVLv
pWqjQr+E3VehnDhvO+BlzmQXWkmstUGUXT8lf78a3em60c2UrzT0fFyDoWw3Ic+J
nIckPEC4EjGY5l9/zbxs7XahcYd369JlFlvJzptpdmEbeR3d3opoQD3ECB2fCuoS
fi6IOGbKCCpF91uORCNo6Sg7b34pGMnMINOwTqvAxXjbeeBRsJ+Q+lHtyE7k0o8K
mJbKNa7IxUV9ehcuLKVBCHro76yP6K1XbprZ+fHsYreMfFvRWsOVI8RIrgBA1jqJ
FfZeIkK0+dh6aetV0A9Sli9MjrcEk7wpfFEqb0HdD1qvphSThT06EATLV/BtthB+
qAlJnP/bvXci6kEyXbJ6/Zdb4jOVUrjcJx2n4BGViZJe+BJCaiXYRppokMrGZOuY
b24jy6i/0dxdztfzMV7tfxWZXpHvr2suwFA4mD6OsggMjCESPWEpBPRlD/Y5XX+J
uNGuOr0qFkbq+f+JFePx2IFKRqB2u4ZFlJwCFikzl8uIzW0iQGFSxD/5ZQX4OZ3L
dEFRQb998jaN4yjquvEA7+lvPPFXrvKkw8wLaBWpm4CMjWNgSHgIfjSIvyWA+Id/
w3lhN+w/4kDNh9tbhr0Z1eGjBBvDEUwLx8y73K57KQemrk2VdZZ1sAkp8u9JgBg/
N4NZlf70kIfaCCh8jQdqGbJjPZBpiD3ZcYLB+N8ZiEqhWfxmZW/y4Z2JEl2TBSjQ
9wZ+mCeyTOQqXIbiKIOqRgmebdpwsuinxEZZhFS1zZmDfAUhgZyoYmS67eTH5/sb
ejOv9xVMS62M1KMwsS2xhge3kU3bpIx9Yrzorg4+U1izgZIHEX/RIY0hJ1OgKGro
ek/tLHMSSQ9mDtUQTBvE5M5dHZs6Scb9+Imo+CWBtSGka3VRwr9vArojZ6U9dSaD
HiOyk57dlJfN/A5Ul4bPJRzX5Ah/cZVG4mbQO0Sso3DUs9IOKKezo5gZC/w+EsbJ
ni4Nqf45eawnysCL37YuLUtCxkOj4v2SKn5W33lQAUuX/6tkvfRq4hKzG50Ks8cj
IKlAf8JCbp2KOq/PBx/pABZZg+w6SVUg/RXrkMZBLuL5vzFrAd/7TmNswrt2rQEi
LOkFe4q4FAaqN8Q/r1YgueqUN0DPYi8YYjcSqLvXzOOf5KzdjMD5ZmubfIVn8pVu
r2ddfJPY9xKsqCxk8vzJGfOyD6aMEx2l4WXD8cYlnuj8KsIV6ulyc0LOoJXj9CFo
5SAhuagCmixcZOdbTdcXAC4llYplDh9+pQrcLYqAsWXA1k52hrr4LYTxfw/Q2sdp
ccPbc0NdYyN2TaXpCSWmiCpLUpR05NZ6dlg6qTpPpd3mDFpRLK7i6tRvGrikUqNz
SgzJzhfv7ln+aOSPSxrXqGWoRqnXjARchru4DglGW5CdQDb8KhT+bLfMUqBKnxlM
8D9Wq63gqScG2mR+DPGXR3LxEGcDnyQCsEl+pEpnqPOAXUpcBwGUw+Ka5Pul/2LE
D98lUvz9g/nmP6jlDDEFlZqwH/9rhciiatRhlZHnK0A7J2dCXC/ueGfAAh+d0TOz
WQEejxu1cxQi4poTJRUbny+Q1HZCLY2OwYZNZnNSgkxcX8r9xC5G9J2uuFHKupHl
HMnVsmoD12/rpkbbuC1nyY+nIa8vuSnlJsg23PHBQKwoOh7OgO5aH6gXyqFK3+fC
ClemnSLsvh/tEh1WFUHU8oaRetSwg3DtsVLGyXt21H9J7ZcIrDD34h3l+WXfzW+u
3NsscvGs/LCY6z1L61aWUNT/RYA70ExL/r044axmViKZ8J6cxJCoOZpht1E7cLH9
AfwBq2pIddwBReWyrtN5pYkGHdbLglx+BjWHwMWhIzywNLtGfVmelIyIJV0VNbQi
dr7CXYLLAP2yM/3ohCdVRJTeqwP1eb2ocIKS+xlVFrQRVU46wk1OI555slsq2L7D
Z8CgGJGsfSHvztw+5+q8xyzJ+jurX+mc2Tw7CD/YN6IJGePm2iw0Z/DWDwX0MzGu
FWX/s6UjlbV62BhWKIc8tfqsrOT/cngFx54Sez7gJl8pwxT+iSFlCq4+lvoULfow
NOipBb6eAUgvLqce+u4fn1rjg3+K7ZxF9XRt4wwgA+SiFLptbzMXGzLluYd/F/h8
a1dNi/dmYGocMA4u593/Z1W6c8UhPrGLn2wDMqcOBCqYwBSM9G0OQNZxh9HkU3y8
PO80mpVWf4cHv1S99YmgIJ9XsqYksNc6BV/HzWapUpxv3siETF9BY9cHN8gBK2SJ
G3ZvNdidZt3MHRVskVOYZgeuirF/ZJ9Y+J0vT4BCDMkx2gdkZ1R0mkL4snpujIf7
vTtuQL7ynNt12H+9RmI5AklwV4i00+Zboy7ii+d0js7aL6Q8FcpFAYCQG0pQH+Jc
zXkiSa/4kiJaUa2WNru9blPAjyrxAyNdG+uBojW/EV36v0JWVogFfWBwfiT3Cevm
iZkEUFgsLE/dNw7V/IxK6Gfal8xVhHU1wA2TZ2PC+dn02++wRoww7WYeIF+Th89t
PuOuk2eUzEW1w5M56vt/ogpOGEzr5LQsq1Ug9Wd+kI5Ph/OG/aoBTm8ZtaQDJRrM
0UXVX0ZhtpzHtY8KwKqSLLXRou/w39Y3ZfiVzctj4P9+6hOVdJeVZdtHgTMMuni+
s43Z77+XEeDrjuB5j3IIBilKLuUcCUyoBjCWzDCLxyTu9OSZi8COP+MWhVnuqfGj
fQPAFJYXLCzFI5jhZfLO4LH4Chf8SO8lUFuKB997z/3G0vJHhkzsKth3cIcwPmSv
jATo2sW98FTLGpf0V1vcGQ+LPStxIS8ZZh+nek5j3zrHyhsBEKsDykfUR3ol48PJ
hib8Nr9+VdnAh+omEe0YxbhreMo8iCe71i03zqcPTDcNVYI+DfFf4kgrCtYVfb93
aOZA7wKyy+IdZIWgx2H0Lu3lun9g3TKwm+zBtvTpuXv8mmsn8JCr/k6nm9jdUm7N
jgldVGi7gtIjsvANud7+rr8ZpGfYF8w4N/LLG2k8hiSkyvjeOtWMiJTUGujMhoq8
4Tc9pZ1oJyhD5bD5bqNfEICtTBroxDSPOzeqkFfW70JF+egXoMr2ECefBGOz/CBg
bmhmTf7vp+uaxRWWlvhUKrYdYw00TL7c3PlbsRbEm1JzM0SgF27z7JI0feb8jizL
/EwX2vzCib5yrb9pwvWdjCyox/lnw1Qo6ZVSMchbjuQjmSRGidcLein5OymVqXWQ
Mosnq5+SJcF3YprcNz+Dx9X0IYXILbF7aaEZgcKf2OU/rf0e8sFLyNr+/CcrkNVc
UfFWa5W1u2gC7sWEiXblIS47HIFHYc9mfCXtseV44de5tgSePA1JJb0CRYF42Ngq
bbQzRfk9xwcHQh+JZSeQMdnDEJsN7Bqp6fkOf0/xqdVRUWh3uCyOg3IqbraHizdr
JJxo/z3iABT7XoXHJe/k+0I9W8iOc+vdhP8sZJWVIvK3LmHkgFwA6jX/ZF4oSKK8
j5PTBfqSeJbFDqlq0LoYX+fiuTOa0DJmtvBSJ1c5XIjI2NcV9PjNiAWsdWUWiSy/
sDOUinLtjhMYfx9NhvDcwxu9FlezDOwa2p8hQiOUcH4VmyuFt8syzby2AQ+OqjGd
SxNj48ekwK+ZxMqPG6npMfrL/8RZopuaDmRCJLnGIjgNaangWnh/BFQNYXHcxSIU
HQ+BoIow11wJxaitm6Im931tcKGp6zg1noo5vOASaK0jlf26x/raM4p4Y5qNhzx+
lDlvMLZ5uXzfYnw05AGU3XeEUVf7dHVGTi3Yy4bK9xBpw9izxFHUzMvUvUzxeP4H
X3lbKUbHbs10K+2GTJB6B0skCItxpXWBhMp1he2EVTYPf5+LysNDpzPdnAZYOYQv
xjYHfJc+jJsoTTgaP5F3M9lrJ4DEVAHCzB+iuu7UNxDZl7nID4/a+hP8h7gEV6fl
djsAY91icd73jytz9vogDdo9R/I8TrnheFKRSIVrsiL/c6G/9LkQSpJkwrOFOWtP
IHBH7EbidGetlJqgGlNSvGRBEU9FrAaYJLQXRqBR1igTwzM2vfyEjQ57q53eUQFE
4Tjq7aMo+dab5mXM8lQTPAbsj3f8wae9xQI5AuXyLD/qIhh2cnlK+ac9sX0CEiW7
AAvpMcehwKl0FjHoadZwbikpK8Mw++Nddux1LG9rZiLQpt5ZdCY5rTkMyLaAmpfw
mo//hjciHZyRR3UswolQpwAcYwVEYPzhtOQ1yrCMSGxb+Yhha5csquhxme5qq0Go
epmkZlCRHMBjH5rpB1hm2LV8ibtczQirjFrd1XekhyvG8A5PWIxdIQrBAaDpcgWJ
FuafYTd+M9P5mSA5rs8XFxvZpfW4HM+bOzZqdYTKtA1mHi6GYginHI+TL3txgSCt
WJGlQyOLq3CKAtA2r1mEYmyvWi3DnqLiUzJ5Sy37wJL0NUUZhXDwHpi2brv+0TmQ
hoeabsW8swzphmNCBfmNPzlL+Mafz1JR5NKAY8vc21BAsH+OmEj1CEq+cCfxJUD4
Bt1//RyiEzw45VbUutkPMSysY0vdLq0xIfNpQzfGBbCcivi/YIY7xyo6DnwXO6DC
suTalU3W3hsjRnAZv6PY5uKigC23Hwk7LISRO9g6jUw5XaWmquo2aFmzAcW/Sos2
Yr3hhDsXbJIjxfmsX3OkFbd1421Yd85XcafKF2zzmF8j6vvyX/QJQRsEB02pwDbz
tsgAa4/07BS/ASO3Igjknug9esHqofFRTXix5bY5MN8GrKihnWcz7Ej6jy2iHj6+
0LU7+pJbSKJimVVqxv+IKkQ3FuhTJ6N45yJFUZa0Mj0sUZiI+0EeVAK8bkYLrLcC
uq8xDYqNFp+RvQuGQS6j0UaU1iwpMWy/KEOtTCl9y1R0qo8f9CQ6QgF6i7IqJRjN
dLU6dEfl//4aEofu2WRLSXa065uFaPoEJ2l3FlOb3JbBL9vP57RyHQtbkwwfFg1I
KVK+MVWAqCMAASPBKnwxpmfVmh8de4MUuT0obBP3JB8YknTaXSqiXETdla+TKOSz
W/fBA/byYQQihkuZ6GYqhfff3YaULKFEzTqnYPDvfIQDw7iDGOsYpggRavWMcw0B
e2HWk3pfyzq0CxZO1zzzuyxWolLce+zUcyqJWbTu8INobNyTZ+mzxtDvAFJESG8x
E3mvWbS1e6TiPjY0gwPxL/FSSETjpA5PgAAeBt7DDuoGrz6lI8j7rlaR8Op0u8Hf
aIDyhK8raGUq22wEGrGrCoiLURd6Cd3a5i5FnMBFZPQtfWi8E8D9Uf0ARnN01tOA
e8P8GJ+j3m5K38iyeEnbF6h/EORgQ+DHe/iOsIgyq9ZoRjw4AKV29f1+g6M5tU+T
nQJsCfOJN3XTv6bTxVTSw/fImjyT66BIlJ3Z+DdlFmtP2DU2zoJxCAfhulCOCTYp
Z75aD23KpzqHjK6oKWGDM9DQy7wxYlECo2jhiHA1VHkSmvqVabKkJqGRLJ/mFwlr
OyyyuX8DlLR2y2Iwm0ygGMn6Ybx47q9IAlnWZ7lg8mKpij4VE3OJo3WrCmcWdY0a
+8AdehNl+ayUVEMw0RqA8ZElGVrfcDweV/Z7BB4R3yM9fce2Pmmb+ujm+eHJAO57
l6rg3Qb6obdpcfIIxRL6AZgN/tsgOqHw6hj8M5N5RocDcQeLrrOQjWtzeMICA/MK
eecmNJg1ePirCNnz3Ieb5MuOsE//xXPg4Ln/SL5I6xYx3i8cHMiwDzReSE7cMH3h
02rHAnPI1UfJfxnzxKQasKpZwAMD07SU0F5eGMr9UJKxkgLmkXMoYe9RMIoyEIyJ
24j2f24VjFeVfQvnMJ5mkFJSxt3u6qU+zHH+nHOlf0fy0J6Fv7k8TO67rj5oJaMz
3Zs5cISrgGSsteRc4iNH/MsThGIDwGoCNhoY4KgqCafkHKJVUY0UBkVOWa2clijj
ly3EigToW/HQ7wQOpnkMLA1gayE+lyCpJJPjrCtlzbc2ulBBxuXOB9VG3XUG5Edc
B/CvlO8BoXuClK7mCD7Rotv06wpkfPbkTJ8h+RN799Q/bJ+pgfvV3xHz5+k4oAgi
8Ya/5S2MM0IQ/KrcgJwpcNLlklvMW8gYrHJLvMZtGhpQesgY+6zxuxPe5j3BO2iO
yCgcPVUDjMqaan7KxFEgljMxRvPT6XVpjRDV6QOT6XpBPHiOgF5+gyzc8pghVzg7
da01FWMJ44+P5KNQ4mNx/vwq2VHXAOKvnA1lZUf+lFAf3nbCZeAUxr8Bin8hFNeO
jFBLHj5orr2hHrvcuGU5kMOt1iFeP5obinhuHJFrHnYzozvbkub/uSQ8moLHZEXT
kNAGrDm3nMg1twfkyUPbIXH1k2S0++CBr89FSkQ2HHjOfITrtJCgkQNDTAN3C+6W
1dI8icHzc2nJ0YN36EB+eGNeTjqc89IaC2UOq0n+zZn0SHpaU5T+E/4Augx7PVaN
noMIPX0kqmNF6e6HOoMJtaSFoZxTCsFpg7pseVxDF+XeF3ewx1gareCOSJtCMo9C
enYuikrprW1o6EBL+Jh3ubV3DtZpfibIAcsVUxiGY4TDqdly/9lfe8dFLaiHGMLr
T8ke5LQzwNklDilHOwDDIlpi+rVBgFLi8ZBXzVgX5fuYkqABIGPVeDtxP8euX0kL
0LUk8g1w6b7UudAeB+BMV/E2XjHeblPYYTFrY0JAij7e3a7kLXNXyHWK2sDjOQE+
0scVTT0v6oPsnbUbny/Cskt8HvCM9gvVKpaAmp35UOIHDGszeIbTUWacJpGxT/2+
K2iiR4IC36fw5mhG0dbX/FQlL+RYmb9KAN11vldfONdVDkcV9h2kGQMKNxtSnEz6
jxQFO0y/B9J8KKqiI6VNwvR+iAgTcU/5NbaQxcUmqJteMlnObLyQfp3UyPBMDJRb
ErerRJxr5clpGr0pI3EpYH7+dDT78RccL3n/gz6RK4r4KN9QuhIDlkHG8Xf0NfJN
Y4+UjWvbMTCmhrC7a67uFG/F3waw7i5KNbBx47xoa4XOBqbTz9tS5x4+VrKNmrZC
Xctipi3PCZDNcx47VidrqzKqLGSpkJyCNolvp5cEpOzVI5Efd0KqW5K6LwJ9sVW7
sYXBTk5BRdDL0/F7dofzHQGfboW32LAvZDAWyo4CStiHig2eHYcmHLpC5NlKDuCg
5ZsWomqb0hR+Ny6VBEQhPUd9iJPH+F9t8v1sv13HK1HG5ZJafYfoeoe2i3Qt+xhH
p+nnqm40KcTd74NKdrIkDSSmlYuugG/eC0UFKmyuQznMt0Hfusa48/P/Oss5cYcK
8MrlBGlAnH/fjMS9mG9K/AVgd7VwuxiDh/PrHxAyaVDyIs2WXNhPsIIxjb1cTkJa
U2/DjFmbHbjzmtNAaxbxQaoN/Gv05/I4OSoDs/kpvM367Xudzg4mQU2wzY4y/D6A
ZBlfSoJCTSDGYsJcncSuscfCS6ay9P85+GSCXq3zeanEXH//jeTr3fmGlQBaoRqN
MoF3Lywz28H4g3QaajKfN9vxCFuQOklXj54qx1Ho64erIhLltYq2pa0FxLye1IzX
A+5VYEgm9xBPhJ9YGp87UgO/kZUXZ7iJ/rMnbwUAf8NYt78JJeIQKTw6ajpkDDQn
lj7iDt8jgZ6qezEyeqgzrbzQ7rYSOzLQxgiHcPWhFb4Y00YxjPDYhuNErhog/lGK
ks0NwK5OEIf2HfG1W33xwIVETRFNOccYXsN4X8RxsZH7WGFg7axPis82TpWl4DOT
+WBUlJ0cg3coApWdt1u6X6hdE0Z6T131gMSTh4tggi8msgq1XBf8PEd+s7sCTaqw
q6qvCMuIrPIc1yKBDH5zB78IbFDMwjCp03HWkdIWD84m1DEBa6AZMoDpLV+Hh/nW
0AfsV51EkUe7kFgRhPJtheiM7NxZaJgiYn8pFk73Xs7HaSM+dkov+OWLYEJrc0Wj
CLn5BwPaWZUJrmIDvBfYrVWfY5BfLw4VDP3K2mSzXm7joqDUpwFJRr3QhVGz/N9g
u8Bc8qr6Xi6c63+wiIBFbB/TJUlwXtL2UFDDzem2V9EE0/ISdgUaEvaOf/kC6CMi
psld0kQxl75+KfuYU7mp64DI2xVTKrREmnfzetO5Jh483C3F0ApQe3zPEEgtZJZB
w2w0U2mgtPruFjrW+/+BU7eQI1DoTplLKYKPL7GlmZAH3aS8aTZ0NdbC0rtZwML4
Fhg84R8kQqDuw8gBhW2dIJRWct15gHPE7wJxyJRfV1rP/dUO0DrV+6JsplHBMbqI
8hqp/AuSiCfb+XKc1GrU/p3sQ4/YldtuuHiOL8A7xxSDw1vjkAy3WM0NXQpmR4qu
mQFJ6Yc0InPSRSC0XtJZ1bRInQUgodY+J5+eYcza/4Ovi5lvIRuuhCTfJyinXs1r
VnPqMLDigpWoYUQUH7bRjb2HchnOzpzl6vodb6Ah0+bO4ltF2tk4KYCB+0Oog2PO
b9qfk3LbSrNuXVTGV3+YhfPbNqipgkyfBqKnwah2nJeB4vhIoN/J2tb6SE5dqy7e
xSLqWikN1L/qk5lnfBQV0X+foj37s5xRG98TIthqQ1C8jLf3RrIJo0SC+K51Le0G
rMuJ4I9mBagfYDoUkyjkQeYKpVKUbk/8NeKZutNrvuXh1MsIAEICozu4GsRh++Sg
ha/xU9fjZilpckV9yiyXA0URjeN42DMeRy4almdshTc6ahm9EPymmKRgd7uUmbsW
mGRC789MTDxt6PqYhU5GOJKnR10AOJhfHHY1B/xvBMHrw7KGDJkBjgg8dsubgX/a
+or5z2VWELMTohL3uKPQHkb25y3Lpf42iXgUPOtdywWyoudzQxoqsklMlj0HLJaH
ag3mRLp59b6tj9PBNTLi1XAVyr9bcJfIy7euQQNBG7YwMRZjEtYZ1vLDOmcBYLb8
G+UY5sbXhp3vWFWDG+nBZrbkd9TLmN44/+iPuIHUDljxs8skmuX9RL4/CJr9ohVx
QwGLfjwtHwWvqSHYSEvJ7QdU+FWe2Wj4CIkwGXn0Ecg3Xkoyus/piuftBaXZpD0J
lflBzgJtvWbLCHrvuW4ms3KJ+nytkR6EFAa54c/H0kk/WK0mmiqtqrCB6qOYN/5j
IYo55JXIjM7/YqhwkCg3xEXNv0KVm+F4ZvVv+vz1m92rqANUVRS6cMAIhr9shK5+
E4WHQmZjSIh02Bt4iYaV7TBj9/P/vcAK0yYAVmmkbFb5Fo9AN4JLkZXJvDuwbcDx
EMmzSYYyXlAMVy4Yap6UsmL+CqnA5wFgNMcCFR6wEiCfej4km5AO3Fa22QvGEWaF
OI9u2ongLeP3+QYVRLEax7ea5EzFkmXf71w+eT7aMwgUwW1uxm+XW9ZsxLZ6sUMJ
GngZd0RKPYQhcCxQm6874KmQbJgug6M1+FlvtPG1RHmvt8htqyIP6xwe6cr4RtkK
5sBmti9U4D185oPyPi8nOPqFMkamVBRUGkyKp6NgbDmMPYt+8avbnvxLlPwHSnWO
eIYEeLS5puZj4Xwfmu1Z+b4nopSWTa7pQyWArjJAklZzywW9cgiUeXQ8ROyqttS7
RDD+lIZZuTWi19kUt1U39Rdexg5kZACclSLOddkZRIKpEouWEnb2NXi5iTp6Dy2I
TYrKoWeMeDTaY/FT0o981MyosS5obbDg9laiBfcByloN85DJENS/3zxcYpWJPzxq
diOwTuwlP3Op3EPHDIpDc5ngQxtoC6EufKzqVGzVObD158RPG3LRUwwG4HsmmAuw
U6/solGZfyCbSCgvtJtPP5WRBxTAb4IiGc+YSe6uIEDxoFPfgagOU2rmLq+BGKG6
nsQtzsMpdiqxtBXX9SzzIF1alWNc+AOzZTZTemJTdd+e6szkSRtyGsBI6YnvC1h4
1VlfTTaKqmgBbx7ZIo6G3rh43X//U2PEeyluNc/Kz9hjCoy+dUil0BXYZ36WLPap
f4gxp4e5pJRBW5ayx1qkT8+ZHB5tvP04xRGfKS465j9/0iJJVxVCKH8/0XGbtlms
Jg7f/PMSq+0dcCNWnioT2vKK0awnF6YTNUDb1Fxmmo51qtHNVf62VEXdJWDm2Ind
62SyJMnPRcVBWSQrcFu/c+GVDI2o/DSokstFwBNxYd3Wz/8UjEQ74vTt1W63ke8V
X7YdAtrDPkB5TQGtg3yh1I9NxV4sa3jLJZMbFSUf2VOvIhyAY7nqd0MbAIk76+fx
RvxUFXy0XWihxuBx8dfONxR3brPMNMoXjtFQNi2t2eNeIRJrSsoTl+Htj+f2xPBq
b9YAGg7af64qYa3beEKulhlHs1c2cYGD2mIaXUHfZ7e5walpVbTfbcai5rY6HXVW
sjkSZH5lXayE5pciVn6aQhzr5xMutSpCAwnitUvX+/dYhWy198R3qTLiIeCMkp7+
CE5/iPf30c6ckgF6StxB0y6T+nAdPIef2bJEEpIH6OBkVw3iUxTvVOjlk60EyuZC
yyN38VEgyu6g4l9xFqT5pzJJa787DglSztWhRnS41zYHJ0kNeBmKDAlcSKaVSPKT
g+aTtaBhzBh1PIMNIsXGwMESwf9XDzw3IRrxTV0kKHLvsiXQWzbvyNneEQC9Gs2z
tQpnBjBB7PKg0X1VVOV3SE5fHHUCDx64pZGIPxeWsHdlDRjcGZ22dYWRzAbsWSBC
M4YdEZoycJMh7VGTgr9Eu+4xNwSeOJfIrJvEmM2/qF8rU5hsOig9F/GWpFUMjfZs
lLWLwden2EdeJH/Uu4+lEA/XceSNMcfvRypc6KyxzK4pxjP9NAG7r/87HlETzAZe
gF1/W9F5zT+emUFQANElBoCVbcl07vp06auEcBwTZQoZ70sebkg2EboIGIU3cUnf
ygrdUzjVeT5rIY2HnkC2wtuDxW493VyOGF2OrBJDlG3Kv53YIszt6py7uJVqVZuS
IdDrMbo1rxYjMbVOSArSxplPXPk4NNnVu/L6n+2p1Rv2cGN7bgRdQJmKPeVuvYP+
f7peQXb1tpnMWKW/IYgTsGvkKUR0K28U1MaGEiC6j/fB+7km+MwuWeaRvdrEwP+O
UA5Ttdp6Egg93S99eSP5Jw06WbM25p2JgPFy61Q/jJ42csb42+4OIo9sl7eMQikv
Ku5M+NrYLbcvAp0ZB2FwaT6g5DgL0X5otcZIdmrguz2NS3yRIT0zZ+XAxaUQrY0h
kHj932USpbtCcA1efXZaWHc1csCaXlROxTd8sXvcsWJXctGK+nhUBJGacg9ev4zl
UuSr4mY52YtMuXLvUfU22kNMV50h94fz6lCXiIAcHlTapjs8HSW47e59/3HzYzxA
EIGbdmAuKDykrqxZUy0SB2DBZ87TNTghtsdtsrS/4Yy8jrdOlVaKVIwq7H5+QpPU
tWv8Rnlkq+WH4UCwtKqWSsfUNMggt+Lf/+sutBgc5hGzE1w7480blMe9UR9g5DLV
jg85Uj2KHqsHxMf9Svif9UJw89YGygSeJPNFglSopGg0G2S0CNmTp3ukY3tgeQee
1Ni+yADG6JBrsI91CGWGq8wrwvqO569e9wb5Ib2Tr2DjqgeMMxmoP3VfiywGTQQh
ZYbFM5gmuvsZEhlf1/IylK02Q0UA7T05ypN+2R0m91ACGfeALcjuXX9DEU+iwVuZ
igfioXytEX4AjW6IAhwEMdA6un79JVhb/fCKb/RF99of8omJFXXVsKD7Zviz3nCT
8iJEkV0ibfhKq1XVYeSqMKYulpkaSrMzAV6qGDUgEo6YFr/m4JVACZwu1GUcAHIF
0IB7I5gNB47w/s6cUZpE+qVXM3e5o89+1vTpPVv3R3aXCcjLQKvj4TNPLk8RzmWF
hJ/xKmMA8L3jev7Ne98+0g8YLadXUf/CCDCD1+fgCx7pKUFDl6r3v/Iuag437vDX
bE0j/d2YFtJE+bfzbuNUR5zPn1qjEbxb7vY9h6DAhasRjvThUJKP2g5r4Un/IZ9U
WmAbD0o8pWh9GOEXATskq0Z4prQwD55MRJpQH3Bf+9wt12lR9AF2pBTtg/QXwUX3
a1bD11rZIvzzh/N8S4qinfuoqi7soPLbz6BIVMXm7CsQgxj0N8HlvktjbYlP4wba
IbjrPU2D6FyN6+TMF6m0g4B51TCwCbGfS2Zzbv2TsJYP08G3pUlK74TPHQYUYwOp
oU1g8keDzENk8sz++fzkJNksa3aOsGY3PElfjekQhBHq9/+Cna+5l9PiP7SxrTkJ
/v7Au7SpeUnF0sguTxZFrOdBh+E3d87QEwI5KXek7OcdaLcfvrBuuBEMMTdAT2e2
PROAcLr2eVjTsnVr8DoFptSiHSla3lhr0DlOYLupreDspuSw6L2Z475i/RD5h96Q
9w5aOFS4miDgLwiW80OhtRYWRc+fuauJUFFPmuY/30hOY+CtIBt7GOtpud6Lwat0
Hrpudz/9ERsIW7vqgpwmnk/EJacmP3Re31Xsyc9X7EFM3IvPJiNPzjQIpz7gCoBe
/klWfV7zjLWpQNILvtjDqlmGuQFPxWGuIRYPn8AG6pralV7K6oiUrlx67W4e7gEk
qTJIWSR8phcxEttcVnKDGz/8BAoXcceAVBzOShYEvJZmL9/d2K7WizS41sMVpvUB
AXarl15HFBD09+aBmUoRAM16qbv6rrqfQUiGMFM9+aT2iOrHBhZ8a/lfrmt/LH50
lTDOtGy2QkpOOtcEEu/P0Pc2mJkuzUo2qHAsdGzMv6ozfwjrqZc0uaym64LdgroY
k3gJmv15Qs4FsSTvEBxk0sep4xQpTIKx0gJBpw+ByaXCY3jdAGroIYgUvyk36U6C
EDMdIRLJ+8659Lc3EQI4FwjMzVLM+7zd+TqXPNBfrRgYmA1i399ggnh3Gp2ZAgGu
pPt8bjTjdqHHCoW8r58RWVWDV3AbYA7PrzUl7L0owJTPdH+dqC2ypDUcY25PT1LA
1wloz2dplytuAIQyeCPe/AiWuUcG8lSrmDIVNZDOop6tZrTz2xeO6viBq4jjiRZr
bNLmG61l62p5PbMlUx2UiIJ13I4pWouCO4Bjo587CjKcwckWCOSeht+aYh5awW+R
atoqyPuHR93tALdg2jkWZ3TgKeVDgYMmzIW3ebbBUXB1JoYH2iCvR5pef4E2QPy+
tkon51Jg85zjHMUUolvE6+SHGUwsTOn4niXIKUJetWUkhPcLvDpAsG4b6oJviuK5
3y5i0DEvaeDKpbHuCm5rE+iLpSK3L2GCbEh0ypl2v9F3FK91qtFZQLiRcA9QOnPL
1gTyFjQ/5vj4Hg8zDT5rXiD1K7a1u0P2Buwd0oO2xZHDyvfE9jxcPzB2S3CREkuf
m2BepoRrcJHTLuT9zX76uJhPn83jU/DBiHmj3jGhrtk8s4+ITsmkyUpfmTEHbNtG
T+2IqnmLOxG4wz/Y/40QTNz/KLmCmnxgB9HI53S5JFw6OEkX4UVCC9WG5NQXIMmO
IGe0ug+im8FkjYQpOsroolnTSi/8GPCfnpmx9JzynaTB/HcWYPCYW/AXIj76HFZq
geoIeeSNJRYBZfW2QeYl2dWzaBWgpsOrXteu5JRBzFw9SFTC7THbGHTlmRAHX5f+
KDzqQq93/k/Go0xTyE7WOjlfFvUOkt4ZemGTvE8rwOULiQ8GST0Ff6o34xcrZkX/
jy5V5FvxendgHCunf7bDi21cMDNtktSOoSB26b4k+dOHH3vGtO6f09np2L4w6J/r
FsCEEXlaQZWSD8jhM+41RC61qSkGZvjPxy7OZwIZq66ZQb/VMYsvIA6L6CyG5H/f
nM6VrsHbM68JCjP62XIVoebePUQsZ/YmIgFhGYIM/RxWoOe8qtXHHIlrp3VNaiwh
eGV7o+sCC4SgNLUknJ0TPlTTTXA4t37htP+AsjLoEM214YbVvl1fZtLnJ/j7sSR+
qRv7ilnZEJ8NmVI+UR+UdZ5qoDmqEePffrKZ9rHTXa8UTDKjGo++X8gvYaJxSZvQ
CvZUwScMsxXjL4bGDIzgQ0qvFkVmnKVj2bhbEOxutRl+Jdq4yDSD3S0sCYPAMuHx
5xnyfvmf7sd/JBzP663FuyEMMCkmIqrGVZPZNTENhRGrkgHD5DLs1o71rnBX5noI
WQN1ZYAF0Pa7PNug8VeHIEGAqqPPzyj/dIyxBrCEEI/byc04+dpVs/aSFzMMskUR
15XL3eEQiGHl/4hTzz+9XOhQRQXiaGOqZuZbP8KASX6hLW8wQzQhfQ0P096IXJVg
jo2wZjbsFYCufyXHuoZDJDi38Mrd8MvbT9EtLVRidtJ6aQumiyHrIBbOnNv/dmDZ
F8uCcXj7EuVxTrBMyeUqd5Yk4rL/2Lg+Yp2ntPj4NXsmNYOQgIkm7nlQbdbr8skU
9JlOeHf+5BKXewwCjAZq8Tvn8UBVWD8BxA1kMbxluznMaOqrsTtXOvjSfgXWaIah
TD4E6LZvdVhJRTa72cWUZQxJ3E3CjS6LtimlsEE2iP9Vbcz8kbosqeAbzivIanlh
mYDBcQxU2sNt5gxDFspDAr8wnafqC45/v87RTTcK/P45BbZq9PkHmLvP+CozhMtp
M6NLttOhN+DixwW3wSa3SK8D8Daj5Tiv7mzCZksNckoJdy8EuElE+OZYgU04qjpC
oQy2i1aZ0G/41PzgSTsjuypwM3ejYNpYEB4S0+J5NOeb2KW+eUbNU7jMYWZx15jx
Qbw8rQdkggWhSZ4bivkqvuhP53douwMnLL7hGBLqTHS+qcMRyQYbFnR6zLNHhvso
6R0dx73utc1bkZQ2TouufmjpuSn1ziO0vg9JCQ3UhvRE5eCTOICcWqIiKUmvDPk4
HUaC2SuL+stYgslN2/YeJDR21ncg+nuyHGqUsrNe0uNFOLahAErxBxLXBYuW7qUc
sddhiuNnllqammOMrNVd88CcAYClpC+Avo80+H6D8Y4rRP6UNXCtsspVz6GAAFk7
M9TL+8aOUukNrZ0BHAaEVZONJGuGZ27LfMqPiR7g+62uA1NqUZ124WHmPO4ud2Bx
xMO2IM39OJNpfnS1RKf6wsBXmkxBZq4R3KjOsu4ffZdxB/7tJWx0+Wi9MSBTKNYX
RgkDv73Laqq3y/rz0Rj5FZpUkNXjW469t0mQwiQ4L8S0hl91xeCRYl3jL+URqxAB
UyYcXwPOoeT7EvrX+T2W6wV1K073ApjiaveObuBWjOY8ujnyGk4H71fLUZaNYqTL
JCox1Wr8vhG83l8OSD6N9qLAh5zLGYTLxBgdZHlDQEO9JpvWzNPblwWDN3ePxxT1
lsK5E0T2FevVKTjgQE00JSSCSstdkoh4U2AtmvnLUCJlhrR7W9gK2mA0SqlnZNX7
/u7xEwBAWE6YBtWnKByIYH4m98l2Q2cshpV8WXNeinM/kSt4jgvymolX7t7ubHcz
xl7cLX1/s7Q545H4piJyV4ECaIwE+eykcfiPrOcqz59dXM7UQQciJE+QNZIeItYH
Akk3Hl+lhSWQJJ8Hz9KiT0tPSxuswfM7WDH1CTNvhlM29UvCnPWO/6+kwaKjCDb+
LUXg2Q1Jmg+ch+XBiNII33+7kyH57kaIQV8JDGKPQtDPSKM0smggYwPy7rPFfkUw
uATuLVkuuDwl6NzIGz5otEt4bT9XCfykbZadbx6+gga0cq/KDW+sgQAXy1XReO3i
HTwlBHTPFkNZtFfFuRXM2VF2VIJorPmBdgv4BnrU2b+ge4VU3FpSipwyf0etbLq1
vcaRSWrU2HOHxOv5XhuoqS/jBLRHk/THnzrgpCVpr85bH4Xmsv6z6ECly3bQ5FzM
gYp+cg+f1KmQjqwzfPtOFsDQBdmJKAFprMI2cEkqzZlDmhtm4sY/cwMUv1naXHCO
i76J6FSh8iyj/qOBFDXaaAMnPPvAXuXconYoNh1o0Wt2jRGZByXQ8HKhLIpuc3sF
NUZGkotFN0UnfKfWLZYODfCvhS6LV6p6+gZWI4mWq/63HY7hXFyOgrFs8N93DdA/
92zIBsZdvT37XISnlFo523yO8nFGxYsLzhUz0pViQZvCwWN8Gfb3zb3HPxxUSVNt
ysQ9HEVKz+xOTKpBeHjmUgCV4OOXbuzX1GG41UXZ7owXdcCyCRVprXkrgd4MN5OP
0QdMehXHHa55GOUbYE1/POPP/BY7C15CszlYmd+/+SbDb0Fd6lzN3j1/YR9jsJhC
lssLyXHsn+Gmm6d1cl+BOwSmZ+quP6TnmumJ2O41nufqJ8YEYuQTW13w/1cMhOdO
nIw/OwaN7HR8RXZGSYZ5WBlAil/guLgF5bvzjIcTu/1Xz6v0MYJJh/hm8iSCllUq
zrbLPGDWALSrZDCj7zdryb3m+z/+KlFLv/T+YYJF6/hw5NZwyieNnINZ2p64Xm/F
6hlC3V7YLUKM+uiSLgS02A9OllXPv0FypFpl8phcUYOMCEO0uAc8PlMvjDw0aKCT
yuFnIkRmCNW0BxZTV6Um/8tWEEBSssBeA83WewVhpqE04IusXZ0/MsK2IwVW6xz2
9XRmC7Kb64cORZb4tvvJuF228p8VCWbnu+k+3iaz9XGltIfhDhse/d0Z+QX6u0H9
AkqkafE2L7gZZMMBU/9iGP4OcCMQKaNQWYqvBdx7ryFr85J2uA9bsVCmmh5hJxCU
+VGU2AOwU6fhX5MztnszszmGPZnK0tiTWtGI4EbtySAZ9iAlO4VxfOzTMeLj0TJv
eVb6W5oGsujGptLad8yAmRKNIh56wgwujg5TqLIJKoEsSjcY4i/TKPfyXHQPFu+l
0cHZkVv3Lr4r+ZI1QeM9NjQ0SlaVHzxghsMajcAnJqsUwJzznJbpjB1WEDANVdyc
Fz0A7AS+J2HyUdZloLJ4q/41LZZl6OJNCVImFPmIrfDRCmUZQ/vHpIY/ajTLnZi5
mxFY73oliMVog8idiCHhDDIKSiRBHr3sNGYW7SLRG7riBIfoZAudvEVwI4Kaai/q
t7ngz+rLjiG4/+mbIlnmfWiV1moQFyq933TC1N/y2Vzq2PQnjJr/3/HIXJyWchRv
PEOXwx9qdyNSK1yc5iGzaX1oXo2xHwYYGUegUX95kG9Kvu34izHmqECpfdeTtNBP
kCR3Ul7T/eK3Y7aeKu1PmxvaxVJAL9+M7IjuURZ+81kK1RyKNPmwzgKNfPlt/gNp
TthMzei2L4dPli1PtSf3813r2Rt8gsD3TCPr3l6QqSxaznrYgksxQYk34qJQqoLK
OKHlohY18lb2KUtRHxU8TFpvz08cBkY4CANOf0n83Oz3rAnZ2HADnLZKYxF99xMr
eENnjpcLAcMc6FjTZyqO3x+CmoKNFLq502bKjxjTQsqbFel0TY9ZqCcMm48FPq1H
DJmR7KGuh6QfVGJKSi3UQDMQ3h7fjqZXFTbl0G1CivqZA1Ym5+px9cTpcg6hBlnl
kZyl/pQxDIvp9qrVI73RlC7UPeTJQXsgBPKQBYrNp1aznl4hShpDvxlkR3W333e9
7FEYqxJPzR0xxXXeK+zbKmWTHxVnlbtOKotv1eID7Q6s+DvVsvz0fD7kDMwsXtZO
IhCoGEiqmGj3aVvwE5bPKpcYiGHgCDnxtp8ThMnK8ZTalHZqslt74Psvv2jtFLrB
DxKMOOAPUCIHRtkJmuoATeg7SPErqk2NhE00oz+UtWr12JGUkA7fxVnlW9pEIQdG
u+3ta0yVEpleMMnahJup6mZ8quW/rLGb1l6bOusNsjWK3MBD8WAcqXCD6x9Y31kL
XtRGrSbWEu/jzq94eK6RROfqTBAlFtVYl6bnvCm7pRIwnhV6N81ZjQTM8X/Gcx2B
Ao/nUizcyMB0pzXAlrEcy0weoZ7ifO0GWd4KOFBNhFI2Q/7QtX1Qa00N9hVfbV9j
aDN2uIbg6xQxTuk8UR9m3W9ROM6+lK7LT82gJfgvjeOun2Goxmj/G+Ekao0xzlVO
RUUrtYKeL+Tim97+ZE/FGUkBUDg/1YJlfU7LYeiKHUt35Bd7NpjhjWnLMUa7lijX
tGVL4ohbaTYzDlkmVnq/Xz747Ktg5yDMizkKjQTU9ifAuUPAD/NIHsP1OxNd3q/f
2/Wd5DoRaELTiA9U7XzuxKBq07iDU0VNNzAO2C80KuPwP2I0Mn8E37/CkE1ovMcX
gFTTeZ+EtcDajOvvUDLf9uXYARj3z82VVCss8/bjSqUAwNBLLHqfJmIJuf8aqmmD
/mqorezhZ1B2jiX2CdFCDCAQ+b8K6o2p6plK5CPPhwjPkwaICP2th6YrIMrUENTA
vW3KFBMRGVPPAzm3xw1p7NztprFevXG7PSvwbZg/PzBwUhhHYqy9/xgjDu6hvn5U
xKAIOiS900V8qRgRp1hfOFBmCdWg85rfhFnUJ2VJbq4xaof8EaArhK2fAINTS0e/
fUDTtjtvneA0B4mB152vYFazoPFMbrbychlnb0GfMwGHtwJMZ3GoC5dP1muk9P3B
7lZI2+Qm0MbhrjasJvhdXV8B17J2eO8OQIPWN/15k0QjbXOJmCDBzzGD6k0M+7Uj
Q7e3EPtCZgTV0xa65ERL0sBPfL78fAYYaoAaYMh1vpPyJ1iBecAzSDn2I4M+MiT9
bKeIH/tnUpF24Wg+2gPSBD04kOrF7jHSyUHL8SCGuHaBksOBZfjLYtJR9KELPFJN
K6ZR862xrQIRxBWv3ltncRH21fxAN8DWpQiFXSn08UJW/tr9r6y6gmY8Qyyk+2Mk
QLq3RfWRMbh66uBZYOD0tvR4Vs28OamY9OhHvLlUNm2dKpGY2XOdw53QmrMN0G/P
A6nP9PEFPyGiGlLDMjFnGHm7i3UCLAWtVumEh1ImiJqQLC24yvliElo8Qr2W7vwH
zr+/B7hI1gWJf+y04Kimj9ZrdzIAH1TtkozjcvsS9O5iv9ShWwfJDLeKbWZMEp/J
2QElTbk8JmVplZ5A7z/7yWJNF2YtQtha6452aTUYW6fnO/KYwHZ0kkoJMxqt06B6
vrMDvueIK0vsflWARC98W08gDHDfzFpnryUdlysxpEjn90UMTzQEzP7HR+qjXgwP
7JJtguv/pvup0/auSrSJKGMSdYmqdJYFeBNwq2Tf4aF02Yj5qhO01zoYU9OMZb39
70dh9xVu4OLxyCxlJapW9Q2dQ1HjeK4Cmmy/NBJZdeBDXH3u1ay874X+pA+6aexA
GP1nYyjaRg5PS/RRoWkrh+IpYRAnNM6ZZ8Ft0/XN+WD9fc406P2ipjqsYSGKFRSX
V6J3KQ7QMB9vZnxnLU7KDmQm6R4El8wgS1u4CTQ/uIu9TK9W434fxGPRe4WtecC3
4106I+b0Get3crqjhT+fYhdKUROOOiLQpfDY1PErWMdvNdG5f1sdLOQydi44mDkF
8hgpaoRobQYl60wcuO8z8cESZInmb14Zxnxq2aqy35fyaZxO4BrOgKWqBjLpSYzo
GNXv/L0vKxUocgi3ZZw5+IRdFMdlV3zjTi9MX+X2z3Q0r3sG41XE8jufFEQ6ZR7d
LgE6IU9xVHVW1iQQ4vLU/9IZ7mCaE0uRi8V7dEU/WI1X1e5E/nc3yYuJhcLBCYpD
RsDNd8aH7r2VH4lngQVNTP7YbHcjlTfvCcak2hXTsaCLbFSJ0ZsF5x67L/FZapQJ
p2KSgjBdTsDOdP0DLCIAAgh6cWtC723s55MV44ZZzoy2+xUOdMOBvGtbprQnqBPV
85VV/os6QJ4xIRY+Xxu0fZ5TWXMRAJRUqz4RO4w+hpQzKNopWBlN3AnuYe+AwxqW
DOm7LPrYEDl5eVFLTfiqg9B7W/gMsI5uWn94Wnin6gt+FSo2YP78UgygQEx+qHY7
HxGmQTcjPtCVUphAUrp0docEzd/Y+u0I1+5wvH0iAsu6ijHhVPy30ZgCM1tkmBdb
iYF8AuTYnpffmbj6dBahQiWEDvwaLD1fix90MAPDd9OEzU7NnoCEmKV5jGBChUe+
QXVO7NAfh/QNH6C+L+ZTnG2vlCKWbBF7tW2CQJiqr/4EESd/WA6MDjq3i5T/ulMg
36j84cEWfd81RaziTrmAbnLMjTciSD96hD8YdHdWkS89125AKUG0cTBU1E5fQWmn
Gt2oaiKmxSVzJFnbErCqAjzmBrfowlEKiznE76k0JKmgUI6bO3U88il3n25wrlh3
dkrzClyzGprkI0zlPiBMINNoBhithdLyPGAA4ixLl/jcCcQDrgJgIKVZTwbDjXWy
aUQDenN3pFPDVBBeYVhRieN+HE2ofkPo3Qn/TU/KPMnHs8N5Lm627HLLUgV9OSFm
Kw2iaihagHiOfZPrOdbVTqhM0w4b+8U239amTYKolOk38iJ9sjjb7S+FG8eBpzuP
w+Z3oEodTTBTGL1Wi10bJnMiv/pxnwSmMuxCoLR88rVZE0aQ3WNzUCl4Z+RWb5g6
76vqhVEo7OBmmVfYyiOqwQXg166Y+WfqiP/vEiSSfKCJpfYQnUzt16Zk48YoYCb/
KXLQ9e7uwgcRRfU3nsFebrBotMVjjBt3ZWXAsZtumxgsZ13rzL7bycsAaFT1b6vN
+fqEISUepd1irB88vLwX2W0NFKqMUiobwy1H4p0I3JpRv516+GiVNnnjCGe+lcwS
+Aa0+vgcdUPU87pqfD3yzYzVJv48mMy6OKGFMIkOlInjykG4gONCihvwngcO3/kc
ggOBsKWi7dBo4+nwQ7PzTHaYKeWmIu8VLNnTxJoM1Vh3NUsnq9pRW3N1rKQpgvv/
ukxtam9dZ7Z0RBP2MzwhOrH9l1zbxUQYstvg0h5NrdXjzFvOoUnHLpdD8xtOkf6D
hz4wi1p6nQlxbx5T5rGJHsqo5rvZ47LTIsyp7ujpg4ZtQ8pXc/4VdafvDZ0FFyvQ
iiXGX3AtZfc8wJZfKWSxpbXQGXySvaXcf98T8ASPV2wKP2nC0iinnC7O5eHbKfH0
Ztun+bOkhrFLMPTDtqph+Vpg5PSQzlzLtbSMAkn/yvhDKPR0wVwFM1dtDMeOLUjT
zxtUroc8ahdx1RS224SJ39IYlHd+huX6F97AJexl831Iategl+EcYHzEugCLcHR/
rIuOAblrJ0sadpiNTQ/z555y93EGFHlTZoiTEo2MkiVT9ZGRhXfJsoxOCIxTQTiU
N8p5JXnlKP0nEoXzcowL5DaDTnyLxI71ILzGnsLaoqcjRaMucvXBjvK8PK9E1kLE
As/risaehTnwtOibLp+eJGuOuwKwHtRK/MZ4+N1kd81nsPtp0aOXuVyUnfGkpMVy
n4nC48xJgUufQU/C2UNrS1stduN1LyTAgTar3xYVRXzb7YMZOBAGG1AnVYIWNmmu
AUuHK6QXbWFKxxgj5TSN7ZMi/kciwM5BTa6HRU+6d/CPlJxSBw8SFh1LIxtc7R2/
nMxZMb0mcjwyFG+dgpu54kdVi/VgLx5QHe7eY9WreRLAu4SEQyHGtOUyswAe5lu2
xltHoW6k+IwVI1SqcIikuuptdnussBxfIAPW+cp3x/ADsuQdY6C1gtfvWMc3+p+a
2ez3BjTLtm2uo/5L71bSlKeRnNBHgLSXlIhQQFSBKCIHvJ+ewHMJwODyBQjXRgtJ
sP9EGvM+7R6wP/NmgN7sh+/HwyvLvFUEdRKQcHD7VPvpeL+jL19dXjixIeJbuwDT
1I9Iw5KgZo5kgJ0w8MI0F5f6vCW32AGRerXTrNSWSbVb5vwNcYcobtWMZm9YIBZu
YpGlEnBMIiuPwzzH9U2mcs/O9J9bhoKv5jLqye7jPQQ5wSD7V99bxhQbIBZMtaxJ
3bE7nnbT6lgVl1pxqHuBrFvp4srPgKNdaxQTbmQl1VFcdtVghMQpxG135oOadBUA
nuteaWWMo36YD+RKZENeif5hyZ1m0Ps8Q3IElauY7d1D9sUEIvLaiebnnBFYcM1v
Qcb/3f7LA+VQCRrRm9iQmj6XoQKeBPJhdJBiZphQTKZFyBP3wJwyr4ymBHUWZUfc
zPmnxKHuG0upsIfx4IlhfyKDV44SJ7ktrNKzp5irIEImVx9PXUfXQvWEv/5UmX83
+k07ufUU7oriE1lp64cxljTqfANJ3c0L54mQx4VOM/r1U910aDjvHXrwR4QF2Yiw
v6Z/RvXlXcmT/cu9eADdlOBftbKWROnYnHKXZqqka2WyK2saqV1q1dkVWYJiOQHR
hV/+YR7f7PuRt2otI7qo1+wayIALBwVHuIbVllpVP4NqB+Y+oO2xOfyyKH4yehq9
kcYgqZck1USwiONTpqp7CBU+nfytcY6n6KQ8WMYnJwsSwwU/f2nvimHmWlL3JyFN
ax6afQzuCwqUKOw7oc4QP32Ky+pXgpuP06BvM7+aCb4HFVQDWwd4w2zZ3fOvX2uc
kCSrVmQAcJPTvJ2C3fjtMjgda7DgWAMkt1/5WCtHkVb/vuSzTWTLoETLgR1NUJGh
FnQuQWTiYhkVp6Ga68Fl7xPqKrbEN2XrAl5q59B9u5sk+31Itdu8NZxlHfWHsNn7
mZktO5fmZW8i8mKlP/Oes8kEo9Rutys977uLTODDUM7lqOmUJhzVhvCI5K31Dzc7
mbu7WWMsrkSGgBl7+/piLExcZSFLsyTzDpyxiDOL9q+mM8aik0FIt1dwK8stAHlJ
suxKddN3lJSzQzSpGaEqFbDcoDdJM+etvhtcjNjg58ANX5OmCsa1pl14sdDDUrzt
3rji0fdS88v8VSrhJPGwbBdE2uobsKz+J+B1MO0hS1z7iWMwaHXNHUExDMTH1UJH
k1W+bnY6CF7qxBUekQNpgN574OE/eumP2FLRagvTH6RPW2P/HeesSiSUrOghwG+p
yV3IMrNKaqP0lqrnDFu75Ozxyvm3l9/9X8ioR0eeKbcjo4yTkjnj3xUJI91bEgC2
3M4pp5q06rUcptyRjb1961+vtj9gimTVPGhWULPbN3TcLTP2M4Hilu+9jkeybDk4
Ib7Bf/qBH9JPmhWRR50rqPiPcCe8b3LfKy+mv2XpZFDlGoAQG2t0xotZWnd5CKpw
cX7u8LcZOxB+1OLWBSKf8n5S5Y5kJtTd2RsiY4b0MqNodMTAtii1mT0KpurvHZ+j
pxTij93NjPk4qCSvCuqRG0quCt/Gdx/Qj5SR8N9Pj4jm6k5msJ98Ji+W8nq+6EZO
dxz1S7fbvrg/s1CSg3qbSXr5bwCRaS1exj/JY3k8l1Loo5Dj6kFxWLDSdzO6qphR
AJ5LMalkCs4Qj1313V+UeNxukU8cttzsqiMlEZGRhXHGzT5Pmybqh3FTz2w9+EL6
sxJivgUU3XL2QSLmDMWcoyiL+JcCVZAOnEZ+cWBo3O1l32XCtjje6TxhqWOp7IJK
bO+1OJdTqkdbP9FsJdPIxmJBYH/xT07/vIsAU3DzK/9OCCsQ4J+FhW96un5RZocS
Z9L3cEqVZQeVQb4Qjv7YNdGaE1vm9MVzMnG5d4Gb0A1h+6hiXnsAhNm1Xb3bVM/v
64zMinvQZod0fJLhqpqd+IQQ+wtxzlRZgT9/usiYi2nJSjvklTEECl4985OUNNZX
gY2yaV1ilE6XkYoo3CavGve4OKnEyz1Y5ghF4pd9s9PvpjBtK2FGlIWFoZJ3n/rK
1XHhn7kHykqYdhNqcJj9vcpcrWWtP4CQoB+GNGI+gUzZtbZ6Lv4QF6hiJpHa79hP
Pbe2RSbC5A/TSByJgfdCRtvwwtpikqfdnud33NIi49HC2voA5580mvG9OYXd1Ife
DdGwTnJWPiR/x6V0nXwlBeL/+U5ZBjiDAB3mmPIJfuM3Uoh4z6KEBmwIMAHbXszA
fE60B/ZAhSzrvMgZeMsuxYwbmS+ML6WeG69X+7YAwegFojqbFNU1f6/nhwuXKOH7
03m443bA5xwtX/mZ0JRhBoMw8gqyfoamfcOOk1CVe05dFPFQLzYuma+Bg7KPORI1
DVN+juCFRgC5JsBxjeU8o+1nMOV7f8FnVHLqy7cLUSiRzprhPUKOjri7auJjiq6B
c6leHQi4ZeAzeLG/L6Oc2somYFj89UsQeFUF4QuyXNufj2OYxGwthG7/+XMR3bkD
ME5q+kiqEZZJXTg+/WTFTzYS0RLoijmB7uTNuJNFb18xtqDg/VniuW8w1pb27lCz
G12pUBrzaJ3/2T7IFl6LjE2Oy+4k6hGnrR+ETmBRGMDGJgsO4sqwGMMNHFBj6neW
EpDLKAuIpEfpHDCObtPukaOShzstB8Y9r+HgikeHu6I0APO+sK7rx9u7Qrbwn/ZB
XBo3Pb3/6Uam/u8rXCNzJcDTOSlCrzJThGk3sy8ZP3KrSDBcr9krDFRbydtehMjw
uZPXn39PIYiolr/Gl5JTRwaE+MVRSsSXn0gzuBwcKG75gS+FgHCttJsi6j8tQRvO
X0rLtM9H0M5GHIY7/G5+HOkmdop6URhLxGjYO1rVMNkSs5z7FKoy10H918G3O5kT
2GibuEANMInSY2Pm521ruOC2SsDrtfcAEc5l3xqg9Q2ZncmpS3XbYO7o505Z3rZW
8dhi89Bu3D3ZySXOrpFvcJMq+FWzykPWbHkrdNHg0nyEQ6084TYnp+Lobw99unxD
3WZE7oJG/PcJ1Rj4tK2mzy0/7ZznKD18fdZgiAcCTHE73+kvTE6zmdZTRaQ73RPE
12gTWRyerGOhlY2bDqV1d5p+NWW7k0m3yIDaU26rjEE4JjZi+VNYsIK32w/78ahw
Vt/QE0scleDPaH2jnO8eGB7IBrhuCvLfwbJg4Vx0LaFWWfcaRCPIPK4AsrWphzON
DLlZPjWsZbpXgJQYjt1WX+scEUlVGU2oCqF5hlOxvNn/wBotzYxXYKxoq3sQb3UB
VxOKEOKV3l3DcaV1ITbD5xLLbzgMuKtL8HzJtSfsA+pnOzBJPcy+3DAIp3VoEAoX
ucK9i5KGZbq3GrVqGGgswyy4eGrmaNk+VD0nKF/INEgrrZEU7Epo8plPfWMGkAT6
dTVc2tbY23IAIOHE6u7psNVXzI+8pLVNZzli6tOC8QcriWGqibTFF8hkPQAboCv0
FqGiTrnNsdlKJr9ZO+6rWv4u82NgRvDKXGpDzW9ZgFmiWktxq/3pEttplsBXJeok
9EVUJj7f3QXJfVgV+jkibbw7/vhF7Gj9ekNd81EcSQky6cS/bcNJgqzpLF3xdntx
lQJLnIczrXI5pfA5+0aHqj76V9omTPwG8WXJmlsz1c2xCONTYqCVbrGEdSJiPIlo
OJvDYZNOGkT3aI7kEdOm3IdTF8uN0dK0dgF/LWpbkT0GV05HJnuQCB12MC0kv6CC
xQgz3y+YIS9yBLbI0dw44YoBcB1mPh7vDiypwSOICPpOZ3YBA2glXWITxxntMnVC
bVCY1dOA2t9KZnEknPDAfWt50IwS4IFkWHwWZZcXw+RJFPBK9j8oiaYyM2raKcLh
cvgcFivxbgG00IClssi8bJ4dZHdnpkNHUrpx2EknTaGzmes2hmWfg6wjTwD6/vrR
W0sheUZkNekvw8nDeFVkNHr5XHBDqPuFOmDNnid/tQLI50SN0PjmIrvK5//K1g8C
VOFN11Ab179w1HtgIbDl2iItTBycchxPUZayuJ50b7F3gM6XveEQFz0gkoOKLMrZ
qPHHNsUg5I2+wrTNPeH8HatRh1/xDH/nR0fCSwqmnHNqCxuuK6UJQZZZCZWTdEUs
ct29HCpZ+zXQMy916wIwy4fesvwba6Z5CISDSdVUmh8IPrHmGoqqE2x/blIulw0Y
Ij43jT7E96+6OEh/QQ8Md4aJkhy9IAJB3hU+6YS5FigHT/XCgOldgikSum1pwlvJ
Yt6BupK+5H/V+GU3Id35rn3az2zs3h6yXqA5xFGkmBPdv1e4PwEexvOZOxT4loSJ
jnjASCK5ADfHc1GJxRhgFT3mh6SQHhTGCbW7FCh0aAC23AezqxKm/vyqQfxzEtCT
SZnMKfsweMwSEMmaYPaYmKAn/mO9Un9OV+hTdTNOEK01sdiq51ZF4Gafxvtm8+/8
RandikpWSz6evIcyqHhzVDwnm2XceRvRusTKKyo9NMnyMYq8jideFo3H6/VzJQaQ
9+ITIsaK52I4R+rXVrSvA1TInlbvD2gi6seCaq84oddcaq634NEgkGS0DnActA61
fQNnJ8tKz/IB3KuD63zYovxJSbWQSpl9oYJNPo2JzadXfpC+d0RG2t7eoU8ngqIO
cCSgIsIqb27Q/da/TEh4PoKnvzjd1LKngRjCvziJ82f5wtlOcI7DTB729WRRFznk
gndHE/m2kFvRsYUGNCW+GTKWILxFbfRuDwWKVujLIdroQxMtxMiPqaKnpZ7ONczr
PphqroLvXyELzHUx6HN9mFHHbBWXsgcbuGaf311gdvVj25N1UWLizSciV+pRCA8V
mQyzGsobcLlLMcF3zMoj0/eXGaYfT/bps/bNH02jv1i25NF49GlkQYOO4q3shMi5
D4J61c/MdMlGq7rJpF22ucBOubVYNUu9c3az7cins/OARzVwAzpXG6CsdaupMmlw
GLFmncgGhxHXiZaunlcFZU5w3zsfdnZLUePRwAOHEGd+1sNew3d1E2m6OyxVM4Fl
8ydlHGjX+volSbCt+tsjMFqWTBdQeAZYDynAxMH97LMSzZUkYpubxvosgXIhpsPp
4dDFQGVZ04zgHtBRXXDsHe0nR6fnqcAkR2kr+29T1yQjPPx2khKHo24mYiKimVOt
EjZqMIWf272YyNbch5K76pjQls6ROCpW/M7hDwJkMfxJK9mxBRFfS6KFL8H0vCCV
PqPVSPkg3BU/i+5kbEFkzkGRVqskmrKmuei5r2tI0Y+ggaOJpqYMpEaPw7Ap9gwb
0VGGfDKuJLgVqfJnqs+7taC/OrVdgWMde5jPqHVeH80BlM7z7oyJajjg8f+KU6FO
6Jkq/dHjWvgMrkenllvpWQxJzncW8NZCjzsem0QjRteuDJ3cQplyeceV0flvJZ4x
RJBQ1U0dz9uxfIrKuOXhlrZBsghIzZfGgs1+K8Zy4Cr/kKb9P4KFMVFJWxsJ8S9m
cakLFDylXvEiVbX/V0A+by/ytyZTOXiSO3r+4Ns546LLnModAkJvHNOfSzhHAZwX
4xUKlAoHXPKt8q+xl4c68yUkXmEsFcfGdN+BuiqKfgdLtXs4Zphd4et+/tLznSnZ
33yaU9y4Yy5PojGWoAG6zR2XtdRLXwMH4Tr3Q0QCE6z24/1vxOyS6TjwDBl6eFd0
aLTW2C13TZFDydS0Y1+fjLbig7349FIxAuq1CZYUX+0BINWS0DP2UBKsU2WtpMlo
iarDbq36bxMjEQPhYDQBIFfKveXfDyfZ6EcqsAjjAgiv+7KqDITbfhyTUTANSk+e
nYhXS5zyEXjVfEemndBs8R9YI6V/2taf8Xj+rQYRVT+1eQCB/13b+ssj7LJdibuh
V+ep/DJKSjoAK/2kRhrqN36wTC4LYfn8F2oqZdS0jCQfSThmvd3ayjyQ1suBOGN8
OOhAkJD+xssz5AQ6ivkV5fv66vND62q9lRxhIW0K8yd4uk3146moR4mI8c9ckP+P
hHdm1VDKmFjud366f12lLfHuytfI1UCJxdLnjLeUWvcAiukFMJWoujC0wc38EC/d
o012sJ0lCpg51uBT3TNG/RsYeP7eQR2Z6CbEPy5eLS2GWN8UV5m1VFaW+tYmTAre
dDmRMrFj8yRFeWaqdPEBvO+RwROXmmxU7Q8yJ9GQ8FhvbzoCFdwmnGyWYD1z5pnQ
uVhFLOXOfiplIwhAf1yOZedAW5ChJ5AVnt8sKksRk16cS/XErIhE+K7v0sTVi3rC
qqiOhpZ0p0sqHJREnAkfUuG+U3gofZZep7GMFQFR/hq+CqbJUk5BuwfGbmJaSyVL
s2tDqQur4YymzF0NTTpO+0/NGUX1j48ETtjdYLTvRn4OUQLf8SIK9QBp/KdXBAue
WCKiLd3oO5S1F6AQEkPlRiI0rBMsNP9j/ZvqKiVifwKGar4KUPSdc0JE17mLOEIB
Zj64q4ity64uy9xWoMdIufSSPRUl25haN4gZCDnx24inG+grLuazl65AlMcO79bl
xz783cVTO7A502rgJ1y8LcxtZeEjTN5uP383Xr8TXSKOkLF6dO4/U6PaHba0E1At
bDm2U/b59+Y9aImKpqsjK0oPQ5PyeJzkUn/pVScVsAHTqxER4yRhZ0BfMcvXqIsJ
s9tpLgN/NitTZMpzo9r+tv6kExb5NB0+YiI/m1gvc3BsNdYfb2Q9c94wTsg40DSv
9ygfrK2yRbIdW5b1PbuhhmytH0udQpty51yJw1tkHvL5+rjzn62kXcZik+odeErb
zTEsw0n7EZOfDrSUtiyjPpEzRwZYeCvEHFI3F1lpNAq3xVjI0QAXQfxy5IGRCLaW
ZOONvXtYVXQTC2yKoICZ61aJIx2A0sVlkxTS9kW8Q9fAy43l8XetBgBSge+2m8aQ
BTo21q+AVkiui2fcw3dQ/l18VeHgimwmtD/jn8qIxBA++QDdiFWduj+cI3Slw2rZ
NUkFRO52b1CDfGWcitBgnPhGXcj1wEUF09TEeevUXNW8IdLBSHAGzB0SpvObAJ2o
z5WDvXKmeqJphjXAPCgmyga/4AwCXiQuD08Z/A6hCSH/G3BDklOvJBzhfuweuCO1
karSoOShDU0uaw79scoNyeiynzTiOeyFwgj7ezhd3OLLYX55h7gdq0HGLyF3x/i5
RhTfKe5MrD4ZHpp/qwBeZ4Lw9vWs9n2/ZZ9l7en2BpVKeE5lxFelQ1Shb0T1fxm5
r6161JRKaE+OXR1TIUKvhttW5AqbOlJWSEGaSj8Xv5zqn6QV77DPDsjYEmUrCL+G
CVTn8k0c9fwGQcU9/e2lHg9k44WV8OELHWxytjaJEvw1hGMpdLNnMCKOnZGQXh3M
653ZDVMdfrR5TqVLDPJOe3IO/1/zcOvNITHK57wXu82uBRApW3MOsSXPNC5IqA9c
UkxaW9O0rcOjwzcyTErFFRHUnem77kiPUv52vmiKP6dgfpLAer7/aM6eyLnQDQIn
6NWq9qc1vjvrg+bsyaYtbTvJUrdH+DroydEuRemtS3uJH5cZctaTWvG2/7CsExaF
MJbEO8/Yedn6xP0ih02P2mIz00XhV+anActXz0suX4erqlh0LycnuV29GrLeRPLr
t83BLA10cIeYt4e2BHu/UERXrV7hFzh4MXAWQFsISZrODcHzPkaGBi290Bd517Cv
614rO4jkrZ1UNX1muEGqkze8eRX9Kaf56lNseOCEb7mjyUHraLenq/6dRyIVibem
IkLCRiNFfd/nAElg5ovm9DaL4H/aftBhEQZitGNWC7coJSQrB0iHHEakxpOlijnH
QZF+4fxgMBtFGRouk/vjULuMw0NFZLJBUKBoUDutD5lT0eHUPOMuME+jVOsjw6t7
hyaMG8Fq46s1sOfhRPgN1YDYTF0dbdy51TnnOsDdvk2IMhk3rFZB4Hkd1eYPAHta
3YnlggodQejX1Jm1yokkfHxW62AFh+5O6RXcap45I+oqto7FzzGEFH1X0DWf2pOA
v/rCu0qmQn1TA2teS5aovG+GvLfwWKtdF11z28R1so31lJZEar5B1mPe72fRkKIA
IrpKN+m4Hhc6C1cymtnx3UQUdS5rWlC9KJc6/t3RyUK1+gh+xVqXjPaVIuhkztM2
odGXvFhb/fXyw3xkXdenvMTgKXkUIGUojySGDnmBzhd6D9yaMTYJf4S3Z0RluRNw
uVRO7mqKcDlpD0W14aSGwN3fGjk8Lw2C1b00r3wfghY6P+lRIsSVQEOkhD/TpdZ2
xOY8cMkhxJqiixJt02IGvTvCwLdaxQHnp+S5NPT9qFdZRAhoN0K1lBB8saYmTCw1
jcV/nc9haknZCo8DASOxvVdg2u13L/WVsqWAb77BjM3JUJZKP9wS3bSbR2OGEKIO
4MWykEYyAaGICb5m6tY39NquAWO3z1cG1L8d9IClnKbqPFquuIupA0GHMNq/4rho
enheqPT+FPQmP9BqdT5mVoTbriuI+AtkBTsg4CWCEy9wLv4GZPy0ZXvpQnz6RYZQ
D2PWTajAS901IlMhSek7LlGDFVONiW95qsU9EyDikOwtULHVEpGU8j/X0DZI+kj4
EvLx11UP5dQ8VoHzlJocq5cYvslHuZS/n77I3bWZbM9em5pdH5YRfuPF94837sSv
CilMO09zvrvgbeQn2SFCih68RFWk+uiEJ0RGAoBiy5MhRxuWeULUfPciDuL+d9Xh
vtnIQSBiRoLZp4u4Rud0HPzGCPrbtsD7BOOtaf9ibum+UyjEXmabLj4GdngnyRcT
KX+SO0BkR3zqkODg7k7UBM1HS/MuktEq+7cZxrjzmeCNVEl9pouL2clpA/b0KzA1
128Lei3xPt5OZ6PTmMTR7MCgwyscgTI7Rf4TNrv1u/Sp1FPpwGZsSY9YUgwzeCKz
1Bughogs38OLnod5HwNTVzLTS8XrgAeu6OcSXYD3JC5QNgS/n49LV8dWDH8LY7tl
CJnEDgeqTtjuVigdozJlspx7jYCUqryZXFn923C2XcJCmeLgaBPey6nYzP6B/m3o
FtFEwisWBrhLjqLEoeduGDwK/PhbPEu/8fWLFdn4GffG8OpkOROxyj2iPKqarNK3
8ojzpGNgHUNgFa9N+DgIdpGSn3B0bwltvaiw4q+DFzZwV8lH0ij37eGWMS2WD7ra
bkiP6CkeihbMNRGArcrPCjiHwptEpc33xu3NC/5YJmjY87BHMo4Pwnh0ykiDGxT0
8wo/0aVgDVQCuEIAv0f3UO4VydMULfxc4kqHU5UoC7s7BRsY8XpfcLN/CppesvIg
cCR5acU0lJ8Z7vhTSZQrar/kQBUg7KWphmM0MAoYR7irTJZhNvXeRX9TN30csLro
n+K7qLnm+2LWgSgpCMwGSwZCuEKGiMqBQfOYRRv6Pp8++/bBhwgL/vrFcCtAWJY9
txpdzE45g63sdMrsISqnsr8Eh7ajVJWKTOA0AEM761P55Yv3tlhnDUJ3FWpPpk/Y
WfrZAGIpLv3vRR6SIHmVk/RH8r0HnRsZHevZUsX62zR1q/lyExAVUuT+nfJqrQeV
3Oie3nAvobv/A4Kc6X1kIASajMpuH/OmgWe76xbBQTmLHUoERnTzbaozBuo1u/5p
XM6jnuym5naqwjQKL5j+aCR8if3I/F7VdFAcAlo7pOZoxB89cKEeIJSt82KkAwNo
JRY43VzIt7Rx/+2hYCX8euOzZuJJBIfFvaWd00h4SMO+YaQ4fLexgPcK+b3HZ4KN
6KRJZbciwTW+RX+OF2r5fvVNEAGyux5+V2c8PllGa3oRaFNQpZhV293frR4lTS1v
B8tegdt+3R7umnBv+kEs9NPisxnJQJmO24tCgoQY/lzjG5vPxQ8wA+D2PK2w4tMo
zOpcmuXf+mZKlXa3uBLAn4cADwOSfkPYUuWvDFAhYimcysyzqJ0IA5PQmSFGul0Z
2pDAtHKdCOdFBWxHUeNaxs0rSGg4X6AZnZ5EUJKEkohqDfhl/xpc2Txqo568IjsA
g1/A6JD91snZENgEcOBMUmm+xxAg2yuwStx6tvj/j+aVp/4K1chhYTe4jlY8DbgW
h78ri4nBWTCnpmuaThHRVPY/ZOR2IvUTsBhJ9mbBhk7JHFGlcW+QFQwSDdNbj5ko
Wv7WMaJPAu+RHNgyyqiKnR+rTghKmTKpR8fMGGm0I9dbocGQot2v2sGfKltco3gj
sQsZmkMKypj0bW7WUADO3H50r6gQrQ3PDGCdBIlPbFPYVxd20/yA8v7Ycgj2Z30X
nJ6a6mkAMn+CvnIuQc1R/EXbyqWfCrW5wx+wVeeeo7ea2B2LCp9DBv5n3sUfQUgS
ADze+5ltaz2/nAX+xZ7Cy+gpz/VI2yvAeSTnDrjR9cRlg0YuBV6QOtT0pfEdycDQ
geK4bIuzzmmZ6ihQ/H3xeEqI+fQnlcoNjMgc+3t8MRCBlwu9PZ2PojwwMrsqtn12
fkJ4cS5Tgo2kg650QUOGez+b3lcfQkOwjWSaMNWC7bEqkT4xG+zrIzbas09/K302
CtVnFslXA2283herffVblVw17NOuVHhOYCW2uPsqNElRow81qgOzL9ONlDBIt2aU
wR0E2vTn1o2OBeatEw8DE2E+3jwyWtfeDncL4+dQdkbubdt4WTpFY66P6JNOEN5f
sB0y/hz0nG5Fw+8LhWMlfLeHKwXN4DCf2cw8PcWMmJ05G0+GGwNWT8keD5xbEISu
jqV/1tkpug5lnbggKWCYh6FeEpcKjW2n9FduoSF+WpQEfJl1EEsJnSyF3OjhbVDe
sLZJFya6SPSvwyw4Bn3FXvKkaHbynwcbchmCdBipbtvXOJ51WAi44tjGMBoQdpKq
pxoXbVxEE0eqQ6YPMAV5hglsBX6dBVqIb5lvs0xlqWO0k7d6/+RaH2wLnc6hyAuz
7w7Uh8xuTlsAIG94GgyxXETLYhPpKEycLzzol0XV0iQbFyK1stZRweS747zIa0WJ
dRy6xx3dGuAj8rWu9MElxXbfJDUmygNypFe3hN3nKrOR/U3gmy3XYSn5TluJRlD+
MwwZ6Z2xLNEjLOFA+pRXxNAPGSttomFSa8s99CQ1duE/DC/hcl6NGBJ5wh7i5fhH
wpUKeUFKysTGfsxGXPMsWzip+kREXXNrZko6XqnXmIvMFzymBoIj/k+nzYW4KXLg
tgC0TZjRIOZu47lrQwv1UlwZw9aJwvafEEAWWZtaROcF2M0e0VIUXuA5SduaqhIa
1YA0wAjJ9W4oYveDGaoRLzSUVuwnI26pTT4T7pSuROR+4ObzwPIMTZkpFabmQRjp
l4gRlE3gkUeaJucUp1yN4nMDZAZ7bh/QirZ476mY3OPlIbZNSCu5akpsrm6KL2ic
soDDKJFWt4oOLy3sGV/04AMgHtXCN8StnyhyFXTDZLx9evMck1G1Wf8ziLJV91nl
NdVorM0EHqf/pmBC6v+K/YO6InWvMd2dTsDZ8aeOcfsGX8eAdnqo0aNFhtnPqSOe
IKZF+yozui5vJCUjG8pP3/wWUCNGmlEH2GWuetQ/uIt8/ptgaXjOGU4yP2CQsNaz
TN5nw3nn7LVJtE6aMtfuFothgAOH+7xosGcK2b6GYxbHgZ1DctEoJkVvnwqb7U7H
pifLEHBvCoT6WnEpPwYMPj1UqvZfunFwZPPYhZm0yyVnKVohPBIwtWfdte3iODfN
xYfRkF3xo+NIUGjtchhi4JpI+UVezcFgLAI+B35RhJvJdcpUKenQlJ7chqI+Np6T
UgN6k5NmnoVsz0Qfewe8p1bfwnsEE/KTxj0lHdSSDjX9JFNAmkLkaq6LdQn0rNWN
mqEJW5zpJSvnt9w0mAaMtSdVp0FYBDGwXXp9A3LvH9Z1VQbvc+iAlkWDCkziptVN
WR5rMib49RpVrEZ6hRifxF1tAAsEaZfZ9u0lWaQgtZJxIQ8hpgsJwlEc6P1844Ej
xGwCn8/aUqBrw3cfSsPoG/LgC71aACszy3aKrvi1sABAMXvBRay3TxxrFnMIj7ny
Wj7cAEZQcqpCy8hZU8kY+UpjGZqVwovptVcXQKlaQB6vDF/OmWi7MGnhQqyOA+EB
Is7RDLUK/aa4yE2FNdqOrad5+s4IRghWV7yQiCmtzhmIvuGvAGn5RyLrve8W0NHs
KFpGx257CXJhwob68Rr8uIk1yQIveJke1n/FFwhtB2eawaWyZk1WXGYe+91ekdag
vTbhn+jSi6jOvBKI30K/frykpiBWn9Q3pudvzKC5jD6gJD92fSB2/mdh3YM83aGC
0gU8XgAORDtOBtKWTY0tRiZU5dcnMQH64qwmrzW24GxLadWBYgGXVWu7011i9toE
jeotBkqAQjFO18WG2Z3s/wz9T3ttgspC88eMGdLIQm6eCR5pLrBwxa/GZyCEtsDo
IfwdtPo0g89j3lj0llIsbUShjuHDGYVIMiPjHfS270zJrNUjw3XxLrximFPMupOO
pU8igAxAgQe8tSR0jfQ5iR7XvhscfBSLF5J15JuF8dlXE/G0xt0iwFWLCz7hgtnO
29hZqAgMrzAe5aZaehEDwZpI8miSmGtM6pY1YQSrK8B/NALvbW37bEZ/6CT+uTCX
BAwCuwYnN5lZjFD04b8703+To615AYEsrc2mJGWJH2tgE2uOSTE0KcZvDM30LTtb
VS/tSiZfsoKhtAj4RzQMQj8D1OnpF0+U68BsVrGj5nRBpF7psLkW+OFT1RnhIFkK
c/g6GciaxaqM/An1thXxlhc/fAyLywNdp8Q9YVN+HMwcfUNZ4lqvW/dQj2cXtKMS
zHO9DZX6qKKkKTecHJNcc092ZK+ZchW7MzZHwPqO1Gr+la70BAnwRat2Y27KihwX
FL04a6wEr/tiEV42bpDOefLN3YPSv3WA1DTznQ2prhy9FV2wevwwE0lNVlnGVuRX
3JzBhsjXb5kp1BlHj716SEo7m8e3upavSD1N/u/xfXva3kYZMKLrnwz+SPh8T8tH
NT+S1Bzu77G/ZikRLDusCkPUC/drxIUihxs5kzhl/oQPUqX/YC9p19ePjwahscXe
QWRZBmo65C6xc5N8EBEiJu3ibnK5UO3azMJvVzyl2ulwUo8Xq8z+HpJv/iHgkQNk
KKrvCBBnnBi/INUtQMEznUacWayjcWS1PJzZz43+X6K7MIxlWG/rHmXVkvOet+Rh
ntgyW7u4wZmiL1OKpg1M5Pcenrr9PQrNSaPRBAT+2W0Yn4J24Ie2YN+7H2Eps93a
LTC90LoCTHeeo5uYzeyRq7JDHvX98nKkzkIZGJrYDDvvO38vaU38WBTMy2bXdDhV
Xx5hOsen7RxJCDpwLqf4+p6K5HfJrtwbJC5sf1iJRXIldeojAtzoKVQoYrbtC6vr
M/E7VVDfSCaMnnw4TnxwBqz4yubDT3lMkKU03vIHFCcr2FxXBUL6kUx5Jh2lk87f
8rf+46i8peTQoFJkDKwXaQhjHXWdBJGl4NEyosrqSdpzGJGHnOuwbk+xgEcsnrul
os+FEG0zlhqMZ9rONJlGesI+nXccxJfzlLPg3Ew2UAdmyZuEcsGZ5uc16u9uN24d
7wPfNUl/M6Ur7Um7HUSmC56mzUERE4sAscDrEaqyYRuInRLueTB9NMmVzg9ae4iV
gSWZsswQcp8XD9xCDMCaqHbaWoAuNpQKWqUTboN3vzHAog054oi0nhI9tnSgt03o
dbQLQLz96qaCqIYrsdsa3CoXeOUuJE6Cr3IDWUf64VqGaN707UY5dQVLLDVVV6wp
mlEIeuFRlllr4KNg7jxzEQDZJ+Vi4XI/rL6Vv7a8N7g+tyERnOzEI/DTwO8L1V1t
cH940eh7PgBRqhqRKFME9CmVmBesiFgfq8UEDRsiXg9oyxLs0e5UoAlbRR7zAmId
z6n4Hnf2FHOsygOb0wh+3KmiBaSR6g2jPKTxRi0g15jMVi4aHEnSOZDvZM3LZxG/
J0ziP52/HYjzZbkgcShKs7H9WctPdzLYxcQFkWZAepU0ZWyvgoMQf+8ucObeyMuB
lu+XnkWYMbVLmFacJRJpuL5M0fT9dVC3aCenY55yjdT/WIsYTUgc+dzQx4IWTi0K
HWal1ajpsWlE/BSkBe42X5NqKBiPlgkoYNv8jtyqw/B6HWKICQFMryVzOLoixp2w
4Qqw5zc7yx5AsMVpCYS4hqZ+6dYqSovfnuPUkrXgiXz1Rk5oBJAEuvC/V5UMbQ+W
p8uU1LCQLu6w9DDsUuNMdgCvyTonpgcI92xaVJn3EkHOo9XdPw8I8rE9RFMZf8St
gKfgiBRtpu4LqBNw5xaksyvtzB9fYRRqRhbE97lod+ZQVGa5o/mfYqapq8g4GzcZ
UD4BPqGoSfhenyXE+vufIdK/xDRAJZKnp2laqw3xeJOmOs2+pPDNfkerocHifLqk
jE2fPrZlyzwqQ+7V04dcqysRbehrzhGGvq1Qv5S4lNL7UwdwYhaQZ2d/GlYHeOdl
PWgHxzej63jhNCh5478N176To+hVnG+HVJLhs9/k5fV0OP0HPcD1MCjNTlntpd4H
nukKNuj5NqLuL9mtm+MT6DNIHCJUjwJbuRGM2GAgxviKs8usHWqnvushBHnjlB3l
bZ02gA/5CruHcyPjcnYXMr7gsHfqh0qAVhFlIzY95GgpW8wWP5Rjjfpr1GLUVjvw
T9jvWs0sFISbmrEBKM+8QxLMGbHZLPSW4yhldBv5pEHDBUlutrkYupsBCOiyGm+5
YHivwQYsBCM9D+VYWyiWjHoPeymzdlH2BqqiC4BXmoGtqwYdDeCrUYp6ixnT178x
Dv4ecrPG39eATEzSM2OPHpEnJbhC/JtoZ3en4s/JcOPfCisccV+aldeN0pwWJWGv
hJiXSd26ofqw42Cfy7qUYz+9WdgLyCJZcP5T1yuVKFQmBK36XpI9rLdahH8itx4j
yA2rCCGQeJTdjqPsH0dyClrINRzXEpH82TdgAFnhuA8WKMbn2lk/Rvy5g+Qv4MxU
ae2cobguLHrt2R0OPWdK0UeJsVrw/heStJKfztTnq6NhVzzM8zwgaaDmHhkCe/6e
lsvsBdFOFO6q2ln4P/aRQ2XXJtoQn9eNwwRH3HPH84hpn4yrygU+adCHttc8v4p2
U6oNhNEbJSRh8mir+4rEsllZar1SKft+ZY8CXk71kDXl7aNdiBzL2Gpd5zU2A9qR
S7R8cDjjnSHacFsYPJxYWJZ2ysheesZis5xsN4hGYeXmPLCFhuG0WGhydKS0gV2u
lYavcs2WKRno9QFrYdev1oc7RDIUKCStFL70YOuOPNtqavKAqKpUyLzpIemZ29sv
RLaEe02T8SBqJEEi/zAxOl/EvZkCtGKdv4QKQh4uu/jSj97omGkvEMbDhfv3K7At
ml6bmpCyM0K0+7PWt3Px/NNc4gzvlpU41YIiJ4meM+vjOoz5k601O2/gNF/1mgXY
nmjayLZiDKQXNQcBd6wXvYDjRygU4Jezicg81+MQ1iIFX1t/LC6KKH/Eb61fdT7T
hGs2a8xrroQCfCwiQ6Ixz7WCniwsFDdA7+HV7KwSkz8kDR8NNjMUAXmcp0FTaJJe
L3t60KIgWONtEIeH3e1cGe3hch5S4Ggn/lHXwtSDKOdqjtHhGT4yUlTymUvBOQet
DhXqlNNiZsuO5zpuqmZvAIwpwvtG+Zx48VDNiHGamZAnauScLGFieSLVhX1nK/Cy
vszogscizGwJiTkM7VIK5QVUvMWGmJUZWBaku0IKVnlvVjk/it5vJtl8M3O6wOoF
4VJqlApXZLSo+NdrTxzSxpy6IBOJP2YkTKv3LMHSNf1H4XYlrlHZcojEM2hXJhyt
Xpca7M+dHkfv7LxV4i9Nhdn1vfhw0dqJIak5r85WdSfaZIBhQmnUMEOm8Js+8X7C
05XJezExlXVh8Zh7EyzFCqnZ9Ui1pZyu7bcYaf3y/UeJQz39qY3m5sXN5X6BG2r7
c2HqOtHW0TAGYGeCjh6aV+8zo1NEyKUcwZpT2lIGOLtkV+wPtnMKCgWv/RT67jcK
G/x2H/xNOy6kZqBiSaU3FwNVSOy8NQoLuC5dGOpRiperYl/XzdUmYIKM4+Eq4HAB
k2dJEKMdN28y0EQ1JLQ+QebuiLy69++G/aj0eeXVXS4XfN2PoU5/1SjiPf5/LpDx
F5lzs90PIrsXW0rwNbBACql2wsvUC/b6u7A3v3BBlE0fxdDE86Y221QcZ8UbFy+Y
nlEGKG6VVrMRoRnVgllSCRJS7MpoucG5LO0yHlz/7SOvy1uAUdLeYvirZxzWHd3V
bBFY1QhLHZEO/6i9yClPLu1FPDP3pbwiESkxjXm+yARY+A1TmFg2Hv9hA/UYElkn
nrmbjw8B/PnJMrJOwNEN3hjO6YKDTPYNICwSW2w4wC0axi+js+6aU7bf5UlFLMBo
loYEJrL1WH+YeZ/k6I8DONbk7hc/V6ONdBoB1H3lZv7Rfs9onF78yhRZ6PESOyFJ
2mWf38YJD7pJoW4pqgAu8nltc/FIrZ8OsorbTEY6+mZTrL/4kkOmNQt4jieotQ5I
TP6YlGqzIe9O6j30QxZdIO5exA4iJQ5yHWyZYqj82qhiBoBzqN4H5S79CPQAkINz
DcKs13QcJZsjMeN47tEmAQIHSoiofArtBF0sunedYQFUd1ofhGpDYBZG8Y1I0wCR
JWeI52W0Su3UgcE5tinwtn4UJ3Qzz3HefDAOdueBueMj9IarN2xEEDIcmY4eMtF+
YnbENKUEz8gVsWtAJkaX1AfSGwBouexeV2Zq0RjbcieTp6ZuDYgLOrws6fr9UICL
TwOhNyZWqmgAaH7XDzCgYiUhofvCumdETFLgACyYjuiAo1g2zZwGoy01T5d/5FBv
frOWqb0Xr0LCOU96gl/Am/xmZkIyEhHJ3fiT9vxAc7RYhYAznD3jxGRp/jRLoq2l
2d5+dGAdv8db/gb+oDDVBtg/HG5Vo/D3k20Uz+J5c/E6ql+a0p2Ot11PTya9JW7/
eNxHD67haTfXBjjDik+vSmhuXGz1f47m8I45m8DVxkcZCqHAQfSKAKDORkhcIuLO
oKb6Aje2dxNIEtiF8uiL18iwqKbzAb0+qpy4N1D/WyHLPHsQEZVwloJ0KFr24cKF
kiPleJxFqyNWDxx5jnth2Jc1rp8tb13zySUADNs1VXbAa78nQxN2gBayNJVeVXk2
5R43Gng/P5Xapb9D5BEXZZ98MkXPzOoNJejlLskSyI2ljHrxfpeFaBYeQy24k+zu
QSWqlUwiXWK0eY0221GOOw35gUdwappR79RdSHRvLUC6YPNBMJeT2t0AIwoOqiz3
2Oh5qXTbNEad8HE9wpG9c7wq9ZcxHJ87bJeZlRgX+udSlMQ5NvzZlJgEV9mST97Q
/6CmvnbH2JpVIhleCOez21QEFs96+vtPgwOAgEXAm6AYleVMe8Bi8vrCS/yxfJXx
rJqk9pO6IXKzuGVggeezJHlC+RoELZWpSVZjzYPx/+R5zuPklpYF093G6Tw/czAG
QHf7ziXDWpdCBmJ0/rCJX5l//l6ejkKPpDHz5gcjMt5/6lt637CQgmr4CqKU+/en
JFnMDxi+DwvauYXc3tBGfj85bgVnEof/7TTYR3csC7YzCNiaSZ0shOHERdtxgwAx
dk26raDo4W8a5Io5DMuuHrJ2jGGzR/9lPQZBaR8M2XkBRSn2zHYj/bmF6wllQlkg
rH5LlC7DhEZ/MJtA7+wjx4h8BTqMjCytgvynjzKJ702KhmyQbjUwtnzbcB8fuebi
85nvGFPVs8wB+S9F/lAf/VnOVjrMOF6pzk1xIWZtVhLrR5FBGO/6piJiqQPjjTc9
jlAZ98FLkpso5lfNj1OcqaeIWRdX5e7Eavm7vcoA7zXtgQY7sX+K/XzrvEPMp+r6
5d4jY5/Xl0zIWFj9H8P+k/xvoAPEUWwi2s7lUnSqEyFnyjMhE7tnQf7I4ktpZWDC
nT5utsmP7dD7tig6nyhjPXQHKgNOLdX8QyVKSmB/WCRXTKNqDAROLRtrt3DznOBf
XTfXRYYZ07n59US4DqlNs3KgMy324S1jY9hY6RztrAb/9INoclvIaFLw4MjAwFAh
qDjBJ2r7eVNZ0Xim/dajgHKLHsu67wXRjlDBsvyeOc9Huj6YxloJ/+C9HdlYc4qB
NNjvS66PCuFEy/bGkwXJY40e8kzSKNgMNsKMwtnNXViMs2AKFc+GVMKmYfutatEN
v+o9KUZPK6ZRXyf8b6azg9pP3wbgfQPPIlWAxm9G1G5YWNMxDE1959LsEnYXsrjQ
JnbY12cE2lbCHt/Jh7PRkXZJaRy9jlEyelEZDUSrkIKN8/1RgDn2L2s3tPLKqBKm
1RL6DkDVc9mTzvDdiSX7cZ6nmr62PSh+MXomVOjP/sqpwFPEcmp97W1t0XMasr29
63vA+GbwKk1UwYAfP0HojDUpPSM6iQJKGmnbLBSRmQKwHtEXc2D2qzLz1XEab+WR
bDOxhy3M11AFM9obUma2Fi07nCpg3L6AylwwZ2uHhm9+9Qf4MifYrgClToL/556R
Mgr/2qFA6dXh5xV4RxLAm7qBw7pX9+8QMBH4+JUNr/6Ou7yTqehhRvc+ZzRMLpIS
wVLgtSl7jUJvhSFUDC31xVKyJXIy4BToai36BuLpQ/WflIRYcc85L6JR5L5eyS8q
Cw6ndyQAmIYoTQV3wOrFfjPf0ipkHq116+NVvxShzybl/lKPfVJx8CulPbuF0L64
NewXSTfVNh4RZ/6vdWkOjFYYZpr41+mQ6AoSe4aJxcAQk8voIlnPdExTpK4A+Jbk
P+0jORRHzSu5HKPAxh4yBt3ZmkCPe69cvbyKfdxounOQ7/9VadrkWb6N7cPx3GLe
fmEFQMIpfqzNWZTy58rl0Y07FgV6H7yVC5fPfsytLDC8Fj/5DoOJ5t6EZAIDcijp
hxB0f2FYrTL8yC0fKf5n7Qcg6KYSleUFRDFOVS8PpK6wVzXU/jBPKsO+4JqzXYNa
WYHP7k08BSJMMpVsWS8Y1WCLxW8WonruiooTY//ajc1GyxH/jfseI8rXjZaUtqmL
6RmAeOzqk7/7DSVYjgdwWc0IF6hhNij1DY8a88PhQlUajkZeQeYmpDndXSGneXdY
8AldFK2UxFLun9tiw5QyIqF8kCv8SAsDRtMXItYOO1B8p5LaLXoP/S2pGowCsUY4
rllNy5aXXsdhvrKsHyXXHYc71mfgOXvcY+gU5CRU5d37BL3uT2NRLRUdjBAKhBbt
gRnaTtpq1mDG8X6wo67+NxfFlmRH0cGQ+Tf2b3YCMpVx9yvesmIgl4penfDvbVEc
YNZtGBgn3DNu2IpajKiGjKjeVshuCHG3vqegmv5a2tc+rebnapuwjTeiyC/c07ro
SDc36Wihqez/Uy9WwseMzNYfgcrLu++9/a2Lq2aVMEu1WjEvgCz/T6SKgMAgO1Vm
ngwI9b9ScbzbZX80DtjHSwXgvZ/guzqs6tslf2u4aENacmv48LU6BPDsEA/Q6DG5
VmK6SGWgt+d2YdKhe6z3PaTZCiThfmV9ja0NW2LnJ8C/iFtNxBCpREB47o4vBk+c
ID4eoggy8uIhJ6d84U7smSCMzEW2Xl7jpxd6mETuebt/Y8vqKQG6GwSDmEuezXiP
k8MRrefldoxycvxS+p5SmAI3b8rnTKNw84xxgjxtEQ7gEdVCQ93rmEFlRZQG8ffr
Jadfp19qZ1bl+dF7+1rO9U36Iu84IIeHEccXPZrPmYQu/cB8WXCIBpjabs8B5mn1
X8OW27Safyjx2ujo52cofHrhtv7S61hX6iZm3F9dR67UgWLs7k4IgTulUxXWbLkT
dL9zRKQBdS40f4FcFdFuTZxW76leF3Pq9ltroYVG2GNl+M2xL3KErzREQfuhme0w
dCfBl6Hedba2d81PAQUq/PzEbh7BbbqKbVTBdZtpDPbs6G9jkEHlPnmYZcpZ5loG
i/oxq3ZOeG12p+J13IWHk5sDw3gU7/Ci/o2Gdx+dGBjyTJmiRcUL/cho4phZIzkr
t9Nk2w4NZQw+b5JzAfrGXf3iOjHZnebv2SpslxiV6+Dr5eE5O9u9Pyur30BMRvvy
fxFd110dtXLWSHVzRC8kVMdCmYoPp5lbScckJFKFMyfPC+FGrzSkzbgBqtzcVBee
FKB+FPC3/5yEYrU5xLoe+klqCgq05oHjqpy2JIUvXce1LE7+06Ne0R9G4BU484DP
EteBiwgS0Rk6K8C0rr/xlaTLVyWWcfGC5ywASS/wLLwyuN+vvsk2zJwQnSwjB+ws
3V/vc96lXiIySb1apE19UTAQxXL26grQIbK0GIX4sH6HVlAlTp345KiDhD6sUN2q
4ERBVwBQz4fKKZhgmE1Ra7ePlUTv2y1w2LezkrX65dWunsUI0BgA6256+ISDo5nJ
dWjRwBM4S6J+YiUAaWky6VpupXYXVvTXsCvM8W4hqvSsVM/TLl8zBdLSsZafZcBp
ivvmfU3Mqmo31WZ+r/UL3aA5lxIuT0JF+D1BhU/BoKaJjKziEtTa4HsX2ZCdy5pE
aDOUI0ZHCI5E3K2hAlsbqmTcBog9Uc3wBX0dkRYqRqRreefeZ+2yK19d0wpGKVHt
0P8+2ZngogblSnxNJKtp0meozO4T5uHYEvtyys0Udrp1mfsM24QKI0YzV9tVZdgG
iHO70pVIe3dmiEzG4UnOFuSz2paFoM9zcLmjk6YFJFKT7OH0CQfLga/Mssl6fAP2
CSqQBs6bKEiHlhzfk5ZcjvM/LZaFbiRDc6fU0t+ml5P+w9qqcq5j1Q5yXSyL80j9
y2WyodjzhAlTtbkhNxUSa92befy0ksAHdV7/wU/P9kuNAb9kZiNKjvx6qJeP8B3h
5RTjaoIzT6j9tP7IA9QvPf71Jflww7VYzVh4CbkrnjnKfBfDJ9QHzStBnAt3Oa5u
gji+b9xDW3THrQ9MYgOEbqMvPbSTeRO62fKBdw9+IS4CEia35wBDSVzNE6Ubej4+
Jucq/9I8KZlq0pzcXdPxofVetskRgjRyaLlfd7S37GioVNwXLtP6xCUV2bk07zw8
iboNQ5bBrkSWJ9ytdenpJ7rzUhzBL5I+oCUa3Xc/WRgCRVZfScqFQ8Gf5ZKmXL6B
wGwE7iUe049s4wWvg3BmQSKfofLlSwLi9G5seWZSEhv4KkykSlaa62zGO5P5/LXS
ANluatv3MZYU5ZpcBdxKqJHtzhkk9eBBz3mo6p+05mi9gXAzGqpg4yKm8JNlcS90
3ICPHwWCJ6FCtjB0rpinYDoZ3ZIuh+7ibhnd827TYQ8DPDKcwjkhh0VKstwATWyM
7GuslQlCubnENW3SPlxfkxrbQ415ON6zch+/y5mggIDp1cPziMIUTyn3kepTDoxz
IT5oeRuIzlszbT2C1QMtOyPSE+R/k1SyGi+RmBxjF3RpBw4Cs13FeC49R59ePuka
v2Te31lmBkE9CYulueHb4AQWocJF3KYatpVnjTKxjmLObwDYKmexL/G8iqTaQbgT
ltPd/tRSoh4Z3ofG/G75IfTomssd2ySEAP+SDuGaIsMPljZHxKX1nr1Wx8k9BSnB
k8JFlUOqRT2g4hfkT005sBWTyJW/2XLfwg6ToxTqFW1iFXIXGPn/tJ9vqMMGBy04
HCfj7bVmsnwaDDUrmQQcYNTP32fB7tZuX6osHs5YJc6/HZjLgjYHjcWKUbdlVNIh
O2QoVxCP7iNV6GtLkoyQEfc9yT90XQglYpirHNq9Z4gIHjWrpfq/g9q622RTiaHC
huaL0G3AuoxVU/POV7e1eH2UKZBELUBcsODnO7ACLpLYdCuI8rYW26pHeoOAEif0
PtBeZDqzyMrXISZN+To465hrHRs6S2xss0CeD2ymWzksb4D7cTjH6Hl4fp+PNWms
3OWgvJpc3iLjbqXlroG791NmXMjU8x3EZcYL7fMSOUN76QtHbkZDg+4WTx6lhPRM
6ErCNjvE9nLucqp3AfSwmzHwnsJ+irabHRUta+NFhaHl1wwVj4eLJEbPgR5YunVU
WpCJnZrpphVrmj2JpCoeTow1Hh/xW2GPiog4YJItc2K/O7Dc3yCixEMWPw9ncC+i
DTSpoWroyVUJl1B9D52BlOKj7cc+hQQgzMV8voyKlMMdqfLp6V9GYfAgLoFTuHK3
ZYFhl8LIjcvV7kRIOwEoqBLmUkZhLzDN+ykss7llIwiXceKykym7o1stHsVGoQT5
2ysZWkBYdZLC834gAzE9zFrQD6ai7FCRaKz9KLt9P7GAxxeDvOdWDMdYTALK5/iB
bpcVdFr+9+rJoVqrJ92coaSwVr9zbqmqajV6zz7J0QJGn0RyYo+1mG0+HAJAHtHU
O/h773qLMG4/ZIwcSfBq/Dn3QltQjY924bu3elEJUDPj2grYHIKPQIKadCLKpVhw
KRBEky846pqckvHIZOL5HzRQor4iyu8YFg2kEMrUUkguP9hXScsdEY+x6Tp/RnvS
C+i5xrvJY41oQtoWCvMsctPlgpb3cqVCd4DuHCOLw8J/56qCGkVYOAlnBakmH/JG
5luuJ3W78zHEMRqlyu90qcijYGq2AgJkslRb/WbH7TPxdnqpqODEtUz9llWaXi1h
tEkbUogUarKTLzN208KVfJeXC3fwBk0S10ApKg4I1evpQpyIMX62BASg4xwElfRo
cJrseqBqHukzqYS+G0C85Bci5SvKzwdSXWNtNd/8mTErj2pkPiaNy15v1vWUpP+1
5DDE/qiVAlPuiOcovnl59DvcUoAV41h/6uAYKf5V8LEUFPbUvuXFpxBX/1I4EZ2U
9rpNVUiRE8on+SY5l7avYXXkkOl15t4eup1/tCrRLQuiHFWr8AH6/8RhXazMXH+j
XiC59J+13artyu5lx5UOAe7Bcdq5B4cDGdUyHnkzvOcfR70RHuTDdt79CoPYmps6
LxZzzZ34DNtLfNI+ZigFZcH+JpqTyVQINolI0vgJfujz56FVM1NA4N/y58Dhn2RT
U1SBmFNHeSlXlGwhicGEDIvbNZBnvbLmi2gk5i6/A70r1xtzmFPXc/QqNi5mEef1
+O2aALkhAmVuDydiRo4ptr6bRBpErrH7iTgoS3i9HCwueEWFKoLfMDrsV2NHaDrZ
m+U8joNLToKL5ttFMCZWg1s6eDQiWWOFBIz7RIn7niLWrjDBuuZx9eAuiQxcYjmt
QtC9CpzsTTWY4LDDHyNSjgctj09PY8JUV2KNKbDJD1c0EV2u8Jme+/FqAw6+naJ/
NOkHOwiFOe5I7bfc3trKZKRj85ev+PVdNXb42UQZ5LPhFpgOwUPA9HsKj243k5YQ
7SZfSYBFeUr3MgbVCttaYQ0K/6bTCOWVz8tZJTn6641VIpskjZsbDA0nYJDKHVOC
a/qD2x6x47M9NkqCaYaIcSSNgAiPOxx7Z07FnwnEd+HjhJbFJRAPbtHs+dUZHvVi
w2IgBfWcH6rftObaDxWl3ZBqARmaD6fUH6ihPV/EMkv9K80llBXNU6bUhZwryw9s
S5Z89ScyB6FEFJ8h1reTl11ZJKaF8XB4TmlYIF1rGXCXEfQD4iKe1sWazgBUYmGy
o847OQ0YXI1mPffYcumWn+77/94yxgugH2iexz2b/5UeNeXUcyneIcB31mErfCE+
kcQ0kS0I9qc4a95hctRfhlQKeJEjXkmLcuZqFsb5JuPC/ZBGFTmoqA7mE+bGERVD
AB8F5RTdWLKF50HSNgx88mDb10Wh4ke8UaBNsR4awwtfnTOy2wAx+5bStAyyCTRP
NYzK+/qt1TqiNfIbnBDF1+ZBbEGIJlPuf2Mjk1p8QFEtsHaE3MrE5vo8u9InAs40
1JNioUU+NCMFWwmu3FFUjMD8N4s2yyCVblrZOvKY0fqeRG2e7gA5FGShBFn8rzDW
OSnVLCZxiFWTeeoKBsADWgitnxP3Zew6wL9CPKULfKhRahLblw/qb49o2mXzwKr+
VTjOyui2lgTIsgIzj5kca4jaJN9+y188WiN7MO5KBite1r48gon9tpRDuWxjmd5w
tMcGwbs0tDAMKs4IV9shGetTJgRJ6mjAsckh+HDB/IY+RN5y3tmYLZf763BtWjbW
1u5VJJZ7OKhhXgjhctKbW4Xkw7OnyQPAD1GfQ/HEMdnWMVyBT0D5fuKGrFA3naQv
ExZTJQXQcg8KSFqxLc3GMoMGgYEsFZKiwMZ98og/ThZPCPh5uVeQSxWjtVEp32TZ
enrzhjQSw7tyannTV31wYv5lyCMCuih17gs9Ht4wLNtpurqqv0zYxya96uaNyMnX
FTJLBWc8ATQc1/RHj5NGEm2j+l/qN3x7ESwLoXaIwm8jSB0q2t84HeKN+6GBG4Jj
6TkxdmNzPyTxZn4RnsL2DlFMw/ckulTbtmf32ZYeKRGjle6fQAaShjuXthCGPbWy
VQtmrAKDPdz3jhgy04CroU7md5TD9VhD2m/x/uZ6XVWyLx6dsFWFMgRcazhFytTU
FgvLk9rJHgASmXHQKdl0U+1X2RtLbkn7SrOhVy8PCkTk1h1SKRQ1p6pNcabAvP4n
9WvbN9j2Y2iVIz+epNjE/zqvYJ/bz3GiMb30eFxWWa1hwLy5jZvDbac6cR+/rGKE
57FaLm5M5FoahYFLPZ+OSTKpYXglFVGcsBEevFjwkhBbdmBIhseWIB0xsb6VBhGK
WWQGXmqWtCyyQD/JnhYDy6nnnKJyb7eYviP6wXFc4U/4djIhAr0taZfH6ZJTxymX
U2968tNIfd942GxacEwkVKi2B+iYnQn9DQn+SkKzsHuf3UOR7KtMeBT83OT7Kvu5
bb1v14+XrXZTiu23kfcEGY8tpLOe4VsMWejw0+CF79jrftOjwFvmTfPEZUk8YMEk
7YPTfqtBf2jMtDYIj+gZPXu+3kAgJX+a/VFjRJQI71xM5Z+moKEFX0vmWieHhDi4
06ASO2IpgaXXKpF/TykmmZiyDr/lA+iVTTkN00EIBYTH3YdVMOoq9Qr12+PSsWXc
vO3Y/HT26a1/x5yfY16O8Z9LWE2bEmFwuWaUEksdiIzW89/5i4MvsUAs05XE2VSm
qrbXF14LmoAIHYwjno4BpHl7G8jEJ2iDrIdlYQj+AhlmOL6ENip8fl8DWv+TSysf
ONSrYNTT+q3GuGOOswHivaGD2k3BUGY/pdA7utLqaYb9L2ONSA4v0YkFVPv6yeDf
JwdfPf5rYRloRn48Cn4tJe9Hjrkb85/8uXWU6Jjme1Md6TD4CICip0Dm4TVhnoE1
Pbj2D3jNykJwsIC+sd+nGE3Z2eaivQfv0bz3DhVoYlz3D5llrGQ7uTSjf87mdI8v
mfc6byZrrkgvmY/h42VKA7ZxlWWNVjIlAjR87TdJdROkAAzGDUFRb4SWlQOy8kV8
lppXGJQSHhvvi5Xz3yxwdbPFt5LXVJV+uXKPHJTOJNmQM02yKZDLwx7grks0CF+b
/06YbsevptZ5VpIDqDWw/6QeVuZ5v5T6mV2uv79J0pd+PQSMFPAjV+yL+H/04tcc
vyhnlSpMoNt8iFnFrZWU4Z/2B4+MxbH2eBi4tgs9JE4gYCQqqwGG/1rGj+8QIus6
RmbTTkt+sq8Y2wGR8lbBIg/Lev755qwJJahqnwGPDqPg2SIVK+3zYSYB5WXh1pTT
wNmMrsIb4bBfi1uqN0BRmt9eCcGww5ZyLaAx3L1yWMwmOF8d45U0gJqVk71UDI7j
raY+sGLvDDNQ21ADWXLVTd3S1VUkOdbRxTDPEuBRQuPK/l4sgcPC0EMmJ9qymq1C
YsKC1YbXxHRdDDV1V0CPIAzH7MKXJR22VhddWMsBsxE5BQ6kZxyVZT940v1TJSpn
QX0g96XKAFRfMPu16mxNsO7SEg9ekFTtT2LxX5+MxVcle++6uYOXrZlxLRx0QE6y
uf8uWue7hUOLHzm0NKyGjREZF4e6lAWx4u9HhhOHVsXYmVEhJPoxyNe7wtc3f3le
CCXfYavFlj3A4tbDPbJgRCJyLA6K5ubZjn5k+6gS7O70Qtnph4zbiMQUeioRPnxf
c6Jo+9h/yw8VmhmV0LW72MeWTokRlS58OoxgT/lEHyw3zJwyTlpH/daarQW7cd50
x7zLx/6lKGTn8pAvGdgU3IQcCpN2igdHR/5OCGcTlFHV6/kyb+b0ZxUwIqQ3Qx6u
IFzXVWevlKs4/AN4A7+i8gB5iRC2A8OBI9A1KmzVwcFX0HanNjpepf5Lal8mqekk
8sn7pIkFJ4kpDScfcdGF3Co5eMV2XtsWmrqkS7VmHdanE2K0SjzQ747m2T42q6kQ
RQGxJaX8T4zo3SBU8aRboKQzmx8K1hl1MRQwlmoWh42Mg/WiJH+KKSekDMgSrU7I
Kog0Jnw+j7N+TKz+BQWRStoEZuqM7isxeYGWJO2trGJz/HUQqH2sQO1f6/v9u0q9
Kn+0U9q6ldDzQ2QXConus42nPRiXFaGBE6jNcUHJgfUhfCw6Oy31A8Z6+AIXPMSE
IWiMkrvDetWwGcayJCgf5uHz/cduuQzkyT53RaFrkgnn8NqRbga35As0PzOrDhgl
Va16r0jHzHy97fudDP4/G2nT7hxRHZxfMfSMhGbsXMYsZsQ86s3HOIDQ6AXz4q49
zhLl+9uqFemGxmOZqrfmKO4B9s4JV/ix0GorxgQm3PHheArhBJPeBo58G8mrsSge
yP5c63UDhXEq/MQldPwr2gjrRnHw4P3LkcaFBHdXd0krWlxML6BTSEAF98Oww7ax
D5HEnAOvwEf4InyKmyGdQC6ah/w8TApr7nkkEBKDGNmN4jbtH1iqExlhiig4lSSJ
QimWDTQBZftCSZ37e7yl4f59gaf6zXWNGEVayjcHJ8iqMNY9LFsRSJkJyUWl1rX8
jnCo0nnORYzA7xHIFW1+nx6U9EWRW7l27hkuAP7lU3agqMZGQf2VD7hLtkOYZJvR
QT+nZA8GXj/5M7uSiy6Kc98wys0JnVbpba1X3ESqptpqEaXdTkLz8ioerZSllEQM
ait0dn8uSJaA8r5W0zfdEkWCgnhVUVZTcxaSYZ+O3uRnWfd4tq0gWBLQu1UoFujZ
Umw4njuvWwveyCCg02Wf6jSXmBKJEBLrAjxZKo+Lunaeod3V+jaCY8M9zxOY76zA
/pVR221KhoWYjrJ5gpPPybEtZGf0zKsOOMvTmbN1Qh84kC1UBrlbK2k/gRWugeT+
HYmMZuUUfpCS9pbzEPU0eN+YTIEVP+gmYqqx2EK3IuXhXAFaMY6al43Q9t2qWH6k
TLTVPQG5c3EszwtKJe467jaMYIcta/sy7NZqn4LcQzSd7b6estoEv+9O31+2fSiP
x+AJMPTTyeILWUOix4s6EZ+VQkdHl77G7jQXtd5SebrnHYe5NrkU/dmAl9J6EMqr
vyXvOLuSDP++FqcdtYpdZm0Vdm5NotH2klBjPbZaItdTybJZz3CXMWglA9BZze5Y
fjwplt2C1W20ReAd8rQHD41qtjNOKOjgKy8ZF0BzmwVFvjBakRjpEDXfa9N+K8LM
Z8AKzF7xzGlbe7eRptnVIo+sT1DKybGAMjgMae/0fS/zdbC+g8OUosvWUM/q82xa
TUlPksWMsqMy9lCYadUecM+GYQKnsQlJLcScZL3L/7DWyTmcpG7kiqfQaLowMF3C
TK8o5tWmr52f2KaMiU9yTNqjgYp8G/bjVsTOhW/rdseZ+eE/J3hehIExbhenXeO3
DNo7Wd4lPxC7SYYKvK+WyYWUhUSjkIO7ilRSa7Wp6pRkXkd2bWzbJ8PP2fA9CawN
Or1iiMY/AJbd5XT6GaZWQ035fymYG96LwB+Dn0fWEnctDqI8Ge4YhxFrgp0gXTQX
Uq8NOIqAVT/Ejo5vnIYMNTacPmIUu4odHKjY09v44vnXmJnvj5ouuOE2l+3pEe2w
kepL5/qEJfTbnjATeVmNNqiNBrYLULc+JWXpp1WtqEWqRxrJzwlUXvI/+poiIHL9
rpQxf/nDFqMFcLe+L8MYxwY+zH6o2a+9d5LLgC1K1fJQ6MlH1unhoKxj8rAarIW1
YEYAv0DIHFVGr4eNrPXjksE6k4cPlvuxT9y9w3iQeWLBmlOHvIhBKlrMsvgDC4lE
uzgebe0yCQYfdkXiroUk8EPnYESqmxuscY6K+5DVtBVAYs+jI6IZ82zPXvntjYT8
+rXbYDRm4SE7GQofkFq3coXT0SQBu9hyUPW+WX0pTNMgxFcE9nMpVXmWKeUL4YTP
zWGWSO+gTAzxA88/aSVJqriLlIrj0HHSirPXweqzZETH9MOqZBE0usNw9IbGmmWU
jNU7082kcOl9sMvuzPuFMK9lt+mIzF2cB6Hhh02PQgm9X2V6IZ0BGG9XMOahn1EN
83uSBppRRRfZUUo/lcL/4ZZLHUUh1jPCLfw/DN51MpMeDj0NYvMqevz7AmhXaBF2
ww9aN+Civn/gsdZL0kPjhSqz299X+zl0P9mLPXBxNnmrk5uYjB5tfKRwXw2gz1WT
mBTysRjm6MOj0+txuaCdhKx7/XJ2Uq0l8qviTMCS/7kL5p/5aUj9wW7oRoKyuVB8
rHtbmCbmLg1lc5249RI7ca4t/Xv3qiMLysM5OmcItBl1FkYeu1h9ajdrkthYn8eT
vCJMWZWUqJiJ7A226cS6r91Gt85+K6npQR1KUJTin3N3Yo6bF1Qt4LaDowLADMyO
VYCbvNtTq+91e2KR+sS2WNJ2D2qavUydiOw4j8n+R1MRCm2BlrcA+YwrQrzr/kbj
e7hUcgyU+zNOk07uyNclmP9VEz/nJjWrdhtzs888B8O13Y/wu6ftchxvv/fAKua6
yzhfr0XdJy5ujMRDMMlZHoG9l+wWF+uz9fzDdhYsUfxsxFq0hVPlR2UX9y5QUyj8
4zlxzTuPJiSSX/S8Cp9S/zMH1QUec3XuAeVc4WhXFsSPBQKqgb92ohYw8ex2Ol+V
/45R4hJAQDu0eiIHhZoq5Zn99ImXERMH16lV7oQ8AnaHZYGPwhyLIQ4oTpEFzI78
HXWsWidH/QE6AHlKWnGcLwDAFk5dFhH2bcujeqnEgB8uf2rS2j1KepH6eQzPeGXz
71RQ9k9FA8PtzT/nE2jWqUbBI/CLEnxnVIVnuTjyrGo4Tr/Zsvghc3YSWUTUKlTf
/lm4W1MrqrNjuY++UPpSn4qtT4pJNEf/jZE9eyLd/VVi5ZKaxu89yP+TCo43p0Yw
rloBBWW+Lc9h5w0Xl9RRplASu3CrraWT+TkzvdXpX+GC5CxWRtWN82H/w7KKJT5S
logYmXn/uCiUmNWfR6dYwcSCP8ThlcUuPjqWIo4IpS3uAT7hRlVzgBpVRrBSSpqS
t8OoeFIAylcpuEZS9+SBbKMtwsJZyZCDQwIyYTr9mIexcfaFfo+0q9kO+KfOKnm0
nAV0fzF+9JN5ERDIynQNFEbQPi9MiGY0HXCAGj/WvuEykMgReGpqmm7UtaSYl5V3
IPeS+v8KgE2xXacXDf2pHD6huiwxKOQzyImSNpgv+c7mU4VjtL+4KrU/lMRb95Im
ycyprK9RkFOY/Wd5RqZMvdpfPEHq5AyE+KOWsWbXZEZkbRXsOALqszMCnx48ivKv
p77P4rRDxBCiWp2DU3fNoA9HJIl7R7xGMOMJjC4EWbu572fzdAtjASRhmMgFEhXN
hrz02Ze2Pgu2rQ38WzyGWzbwkunD5vu1GkrmNmwSdC4QeoZVQFcefSlBwndrN1W2
1Tuf/YD0XHMqjwbvYVjjT6u4XK9uHfQfwj/sVxZrSyVIPL+C9NyZcTUDfYEcPwSX
ZaEzEYFlW0Spi7LcS9zsntu6/sa6hSSJtsoLViWklOHI09qjNyL8ICDBBFAqaUih
K2/Z0NkfyidNbxylHl7aYYEINTujs56W506Ux8gNBwGiZ1jt6NvS94H45hYIu7JU
0rbUvbFUzC+eKI83gPzvHo6dlMrshC39oGKd/BFFFVCIk6Muh2CdUFzlMGp25jL8
pW8ubyyzk0LImoGrnTVmcRIM+hRuSJamulIhaMbt1FCNQJtCs/W7tZovUUtDHYKq
vsjUlVJAGi/1WT31EeI9k1aTp4kImtmc14FhpBOIRV+IXtBTJwnx6ngaTqeR7fIN
TLFsxtSBzbl2CqR2vo866elcE1MvgEEBqCCSODq+oC9lOR4/EGV6XzF/uRzaERM+
iXW7O/WCoRewWm4pygplid50YyuLnPlhUVJfcz65u3OdBwHbTmlKIf2aoaZg4f7j
hN+zxydq9CbGLI0Z9PlglUXgK/aKhSCQRLFvbInP/yokndw9Rb/dZ5Z02hGqv6/q
mNfkDsRCRS7gLews0N63F6N4M8Ss33pZ+SvFkJZICA7fWU5kyrTC+get2508JYHM
KIz+xxqiLKsn+nX+TEdoj8cM1L+l24+GmqdRNyZ3MnzCMyt9QqFs+122rrj3xG4e
vgGhWn2yxXoavtWcMIwLifgPybwJ5WOJS4G9f3AzwPjqTn/iGiq3S5g54ANmC6MJ
ENSpqV+IJUDVNXKWakMbjIf6Qo8DEelyS0vpQ92Ox/IoMapDW5Cn/YsIMaOm5XZW
DJBDzT6QRG2Q7f7CZd6gXe6a+1pnRWhKq6HJisaiJZjnF3VT1EpwR4yNkzKOj1i/
Raj8yiVRW+PbpqGHlsn0XtehfOLymynfODsz+oI6fC33PBUjNEh7F1BTU2BOfKsZ
U3RDKHvGWsnjEUDP+XRv4dX53XcAr4ffHC8iDkmxf4CjGrEEHZWy5WIaddN5Emop
8/WAnOcKlgc9JGSlrx1XIBV/uC1ovfTa6j4kYpSrQ5d5X4rd0Ae9HGEyvHSo7uld
VLemhXghIv7t7kmDRoLoYnLz6AhVv722iZecFlN3p5kl5HZ8VYZFuglEbNvrxO6S
NTg4RaGaqch6QFRS0smFyJmiQfAJJdkMzWmUoA0s1CvxbbCkuKJMW+ftdX0rQUcP
Gz+bWvUy8UW+iRxOrIb35+Omm9/HSkiL5voyVqsRc+Ww5+U49WN2HOlR2wOoPZwB
qEOz+3x3VAZqSorW01eB9tfWwwBg2L50lmXlYLoyqLeqxYHVpnpBBIdPK7RF+7cW
oRm4X2re0b01DAa0AZ2BW2Fwx08yU550oL/ILYDa4RNAuOgxsFGkkQ7+dCmv0Ni8
Eh6OeMnIWSekVUtSjkX6pmzc/gqeP1m25wM8VgrGLvCs0Igj/1Lw49GtcaHakfJA
ws0iqH5nGDsFtNncr9Z2DjyuO31sSVvTqdaysZxBteGqdPt7Cw3pEngeUHZed6OL
y3jF4KWoOp+0aVvcJU11rTGKZ/XyM8v8TDCVVaKI16wrp/7a83xkAHjtHJ/TZcvD
Z2XQl9YaP2zXVVqarL+NAEQ003pjD4EuNj/oEAcVGW6YJVKtEfygcZOM29D9tTo5
jns/0SXIxrtVABM10suD0BQLZ4pItBbt3kMQNgSBO6DEk/tT0SHbAVmeRwPzBl8Y
xSnBzTobelhHRFPNLVwRienkLVH5GQvmAwWtgl6nEB72SrMd8ogku+VHoY6cSvSw
2gt3Xpoz9ZWK3ZNR4spA0xoMIlhJCS0OcVaqJTho0Av4v1J+Zece315jyT4Bn1Af
Q6ZSZKictVmaWAe4awOBinghmwfZYGulxY5hBeFv5J7JEOKnjKMGsdFt/3iBibNq
dzss70Ht/MDc+X1m4hLPMQt3EiZbmTQ5PZpOLKNcWmWGiNtGqXdFnChtcAgunvPl
wJe9xBDxrrFT//I/O6g6TuVb8w3kHu4zq7LEhz+hearqq4FVtYvV/tj9D8gFVWuX
dfEHZuch5fdjacy5fFvOHmVhRp3UXCbu7F00rSiDSpHGv6RYMrd+OeaZ680s4uxn
npzoIFlFDRaDk/GjAtT1iUcFYXzOK9XXvh/KzbAsbVgWLNGV0Ywwmp8l6T4ef6Ye
6umTAmggw3R6SIJWu9q+x1rz8KiEhtzcoTk3/8MWieTdY7rK4A8kViUqXQk3tte8
0CvV6ydoExXjHl7EWX8vnx8l8D3ZAfMtbebviHXKfcXXPIuIbLninHy/GKcTVtLL
9p/Bf0TJnCe6ctRFsW/62mhMvYXb71h0POCsF03yWak2b4oWn5ApTiZBGvpWRcsd
7h2+8YnKdK1mqfJMhR0q/VCD3cUvqirLX5loKkQEdzsg4TNjw1JLqmxgxlsthQHp
1+Ap49FezEtpXnKz1v6gTfY37XDXBZfRj/b5ayo+ZTfn0lM+ezcvSaDwptXZwbVD
v7pX6GAy/iyYgZlP3SF4ctIn+39wy8k+/7Wlx+5noOaHdW5uD4JdQULsMCiE5j8F
Xc21HO4wYQcc5qxwLn8zZ/2qj8n5v/QVnnYOmqzRjo/f6DXzTS3ZDZLD/ZGO5oas
5Uxf9vSs6UzV9H4SIKWaurfhTILb2T2lpufE7eo2OWztuTuEqZ2+XkTQ064aIyuA
g541owIJKQR4AjX+DpGfSf4RdsFPRbG8ih0gVPfOjkFcFFxfBYbvFPPLuWzbniKH
snrZlbhURo6zu3/Y8urS5lTRSt1dfQq1gRrpArTbyL3tlPyXs1OMcfG6V/rJmENV
bgfmrr3/Y2vT+ZY8I8vEwz24HX67/+exJxgsG2kkIboRRQt84ncxgx7zhIL28AL0
5jwKNjyUBnEQHpnRjpwo06ppZQZnUR3vqU8DlbPsZVEbnyUvD8MIplPlWkU6v/Ly
PeXNoV8RtHp2PpChbNt+rUvghbrx2B6g3uzYpzUpBGlK5Eam/om0i3vo5BUOu6KD
pIBEUej+KfhzZGbzG+mMfQuaBWQx2BhnvOdcx4uB2TmAb5tv9Rczn+j/ald6JoII
ngnlPckvtuR02M6Cgrrowzt883kBfqkvZCchfYiQWrQeNRwShOuQ6wD/Wt5nHxzO
j6oUz+2dkdb5YVXGGN0d2azXRVxIvm2ocnP3oNwhS3bE9Ck7IExcFO1Ma2HCYSjH
oEG1IBWC8jukz2W7l+tKmCdF+/EBye4BC7Idc+5kmhfGQFDy7EIjJ2290d9O+MKk
aTtOXtN/UpstwCmSpKUGc2On2zmkPd+nu15+cmAHrVypl01oF2fYNpl5uc/rtIAd
gq6DKP305Ou+Mlf5pdIWn3RvDOknXT+GpjLtU9FoJP7Eo5sf3edXcEozff8KqmqM
5L8cms/WnSsDZ7UfSuhxkhY7uj5irgxZD2xiimjoX1VDjiplWgtfYRW7hRlbukrc
TSqHv/D5/lsdoZ+QHuOqEplkyeVJbeACfp99NfVSHRzP6Uish83se/ESm3WuUoG8
6DdkpaPdT+2wAy1k/rL/lsikO+qE9VB+GKohnCRMl3oCKnNA79BvvU0e7bVEQPZu
/Hromv67vUI83+Sa1nCwbi6mP0QaOxxW3jN3KUCbXc5XMoF2xqK2DeoautaOUCLP
6EF1YdM9vHN/oOgetl7OONy47twJTosE6cTScQbhncowRQsZAVZcJa2a1gMiuwQl
QQytpOSfQyYiLbDG3oH5kv7IUM9dyyiDhtuaw5BqgUd3pf46snZishMRxXFG03kO
yZJQIExCGkpRG1lCr8e5VvDbeOD+akVwjBfGR/pp1UJGiBSM/4ak0hAaqxxStM52
oLRKaeQ3nTr5+IKAf1Q9mGVmc6bq2ceNdyBW6wN2lad2uWHAeUZXi5l35tL6jpw5
N6g0zH/ikBEOVx8o2b6hMrTGO+OQOC5bt+bwSWn6Ow3yQctPApGwpwz8WFwFQPIY
mPXUyenAOec1JCUglVFPBSbcSsKPwEal/FWsA4HlS2CXxBRmcfXkR1ja+qNHR1F+
S/lV4QO8+GZ4mzrkwyYXCrDkLqTPmA956HpLGcpKk9JRCDoFnXZhxSzu0cgE6PON
59X3unp+sDJ47UX9/5YAXbg4ej6DwTA+DTmbQu2q6mDx6ydIFT0CbqLKmitIQOTd
Xz8iaddodp8BBWyLLef2lpf5kGWSgjCujwnd/FgMQyJd9Op/oq6qwVtzjD8jNv91
evVQw8KQ9k3oIKLKsFS7zV16FcY2bUxdTMUyYCjjcJUDlOG+VeNUMyDb4KC8iUCZ
tY7wbXtTcFs5g01tuvvMGmUv1hKa23P0kZK6uCDgfKVx2thhK5jMyINfphfMLGsY
Zst+8fqMqpeFh3LccdBG2c0lz1ZeaaLTQeH0a3woGdb+UuYd5jFgevueBJE00bWS
cLONIb1tWjcUl7LvTAx9kMtDBDyjXCoWpAz8xuPlLLEzTTVP1FM8NJomoht7Snh7
Ev9aMOplJds9hHqISXF9NooMCh5ab58t2RCR+qmc/8YgHAGrWFcbZZsNN4uU5NLo
a63aySwXO/BgPDHQbKt3K959OInILMNBJ0mF2AogKDS0UC1/uXQupiqDnOTUGwYt
Vuke5mQcOA30v4E5w4TJ2zd9oWXTf7MlB0g+4IlEoyzTbOIlybyi04BNNRyykzqq
RhmTiHJybvptnotWzZe8gtLOEOEgXnPpAcCv5DbYGdJrBIcyW9PGSRejDyWA33Nv
KbypiZbWeV18EdFL5hz/3wQgRed/hb8OTzYqoZl4PAG6P0ySsqqNpdx/hN7mY9xq
6nIreLSgmFjdCp1slK060/WXkRKQ14OEafMR8ux0MoYXC4Q92q50Pdp8KOqnwROL
Tz4+i2XyWaG7d0+w8xHbBw88Vu6AeQYxiITkOfPatKok3JnJ0x2XD3jI5Gvx2ujO
zC6HCaT8Lj4irycNbXkLpECooy7bF20WWnMDgDwrV79OaqCM14A4m35cLl8s3v6E
NcjRLhYNK4WEX7KsvsS9Szk9RUdvISilVAxHWbNXTHBSz+rr5bLp+VzmsdPOtO/b
TGHtVA7RMOYOMDA+pI4zL3T8/BIAgmX2an+5YFzN1535iDG5u6VL3qB18Ueeml7r
EV18sUuLvBrI3Zj6PZRnPj7W0jKAUQYYWprZ470CSQNt8cMS2cDIWlwruhdL7VjT
aWJEAW0SvF5e2+/MAAY6a52HZzZVO5jNZ3id9nDx+/RHYVkrQ88rI0abXXo4PO5f
aZxe8FJt0WdtrQL8lmGEqALt9byxMH3dYbNAU/eERm9XHuLSo9gug0cqYlKyTGFU
i7SgYe9Lldce7SjYIMAxSu+BL83Hlqh93QT4TyQR8V5BSJA8YHoWHVtnmEo+GLFr
FjKY9rbIx1safMMuftArDFIrk8dc+72kVpiKiGKTOg+pkHNoKEZulq/mGKRwDacE
Rgcz7ZPI9L8FR1lhENjWkyM9M65RAlNDNOf7moBKOfgxqsHPYxsgiIVr1Ffd+fNu
isoSlJ+aBh4X6PbW/2MD7/QmUUoewkDV2ri34pfFzHeQ3nQmRcuyGvmQo/eos/YN
wKQhwObfPqK6hfnfzQI40Bg2pVO8KwlS0TyjSvW5UyRhs5cOi33lnrOhaHv+z3Sn
KvlpbNr2JuUMLW890hMVeyueRYacTDccynpf6Rriu/5veQw4H3nBNu3qkO6ej3LO
NRte3LYv/u+zIdf0PAqS24973nSERoWVUevqBT8DNwyQQbsGES1WkQx7rliqoEs3
Ne64Qy6NwJOF9tVmwlddMV14vxK7au+FwlQlTUkiJf4TNzGjnMdz+Xstg5QSPb80
333t9Nd30XeCaZVWe+9woJ+bDOy+g/MNYmie/oyjuYagpnKf15f3vs8Kl2mkL7gE
WYh287GGMLIG6aBMXCFOE+ktEkRd0rpWI5xh2IL08Di+N98MW90YUcGyTqRV5Y2R
Ro2s07+F+opxcVdFbK23S2PAWXoOEAYCeqbP22M6AN8XD5c8O/cwKDnKhZ6Lwy4L
77U3RwWdOFTQMpfiJ6ES/afGtEiGIKxKyluPK5tkKnzjbaNbOf1wpLPs3pzCOR8s
7pf5EbDgf1VZGwENVyQl3mu3F7tcndqwSOHS9HgFEDIV7Ymxm1vdJI50sjKVrY7w
GMyvX36IMI63kQRNLdnoNTnVtSP9chCR1wK/vCp0V36hZxe6LuOOynF2fHHAZcT2
CxhqH6WRQkymqFNfAozuagsoSzeLJnwxs5w5QwkscHOsZqB5K8a4xyhnZ+yY2Iu1
01LnkvpfzcYyq0Sfvk+cCyoWzg1Ox6NSbGGNlJIONVkyzJlJUKbd3DHKJiZ+k1DE
cTMiIpcfvQ5VixsOXYf2b4m+1J7KVjW0adAGO7WgiQPayCwFfIOk7gpPq82p7p2w
tyja33wLfs1ycB8nfV0qlYb3nJ8WWx5djUNlxV/TJeTxVkd0PmR44JnR0EswRz38
KYtLWxwBnpjJkcchSNIQSC23whN6mhinj0ECJr+QkLhte6R2pNlG5Q/F6tHtmuoA
6CmJ7fBvFoE5fkv86myoOhKr3zsDqRpj41SldIZg+uZiBrGygWS92cnyphHjAEbm
B6j9/1FJQ7XwPgU8vpPjWTDyFICGebhdQGCR4ul0ynYgsZa+QGgqh8Q4il2oloOC
AaxIMYAjCCGoUQr+Z/sGbdODyYLlAS48UXVACLMYihsYiaaZrBo/FQE0hn/Zvch6
LZHGXiyqAtW819IKj0eUvybh5nwku3pQ0o4odo6+cxL99ZChgiGRJ6+gvAMupdmE
5pIGSL/AGTn/4jyzcsPmgCxrCIFxHto2JOcgRVCer+ox1rfmfXdIf78uV5Ku8Oe+
56rT6uHT6JYuiWLMlXxzSbyU+6hF8A+L9fROyElV47tYzb3sW6meO54BU5r8SEHk
xul5p8GmB5xoakztl1qptdgxQ1gsyYpm2hf6/vemTodH/5fZMhaQKsapJKb32jf0
j5vECmY758r1Ym7rZ4dD4QR3nvKHfNf8hT2mDMQlQAFx6SAXgN4+bLFMwNysTo/V
f8W/bMa8atuX09oggipfo6emhRi4cnq1qgnbpjkVCzPAtyPZD0JzyO46qig6Z0cY
PGXiWuGr5CqU9v77NGaNLXZzELiGHAPtbr3wgk+hoBL+uxCywK3+nw193fsKvt4+
mf3xt+D7M9Zja1W83xd1fJ5VAXi/RdniwHmirHTxSrkKgadSy5Wnoot0jjJMBuO9
AMio9PSvsZsOeqKc9EMgiKKF3ITmXtWss8wXKWzKXZ+hrD62lo7mRVpSjl087bIx
3ZUn8XbJMa++0ZEIO+6zOGg32b0Jh3+ncMw60g1ws7bHqX1KGakKh9taOwXvILre
HZ10mRBE3Wg0+6Cv7QHFyeTImtSaDwcL8cSt15t6qmvkDdLdKa95w5q7mHHmVVYr
TG61sPFfjIzwt3mtdRVS6P4n7yAy5+aU+oW12gHReZaUaDqcW5NjLX6hzSfRQi58
uWPPq+eO3IHf5gUi4cRf8wbeUb8KxG521AoR0qEIrgPYrfusDc1g3rnhmiwRyFmc
5uzHf9gfhyL046Wi7UlRTK3+BT3YW4jOhVjo67Q9o37O5+ea29eQ1fJfCDLg9SyQ
bwVr6uGF8Ot/ItbPElFUlVzkYs2qX3y0rRMDvSfsEKgLFWKeAnNn7jEmDD1tw/kR
+YmBanmxsTrRb56wvAJFhGQ4OPgoTwo8GBU/fXn9JPe60jfLy4eSerHMjqkRb1q3
K+IVrQF+mTfrkUe46L8Ap8+bi2hoAcPCsjW33iOPgEViWpvm26j+y0O4J2JTc6cC
6Lc9NqhR1VEZqoUS4svDxWdY4+BeESd1MGpR/0O9NAz0GT4ITHwidjq/KmEpUUEH
p9cPHzux2fMyHUG6sFZbTXB/svdt0B1cpsWOVe+GU+mzSrFtrFYz2S2Hjk10/Kb8
lWVqJkTETd6qgp3nEwVKMcWpkN+WHdA0ZS8yn4bbRWehfwGSNYcu0lKfn6ywO+0z
WO5Y01ltMT0YpCLoZ2/s69dlYViXAO0IEYk7PERkXr7STxmXkIQEqAbFiKhwuED7
ehXuzqUJK9Q+FrNhmhJP/F2BCr53/E00oWxdekdqsK3CZKMb29Z3aNcT4EvGoXSG
HVgG0/A/aSrYN9cfX9986KMv2WHVEAsiir44WMHkhElbDaYj6KZLxaatWygbe1Xr
mQMN0ywR9HK4/Sjk1dsg1EBz/OdvBT5cSnPTchOoCKk11tWqaZwvE2iwShu2Csj5
q0I9apyBGXnZt1+hml2YCbmyOhuN9rqCrnb0SJBalNv2OgD421AS0Gd0aJto3NQ4
Qa/n77RLhLGRLYQogPTUnPfL6/FZ2dTOinVN/pURlaKXjJ9qlGMLn23sx+SJxWNf
Ydn7vPqUQXHQl/Xj/mJGOyC0UPAU0Ic7mMi2d4xJ+Ssvr4jDWj2OezmA2sL+Ke/q
uy2ZPYNvwcOo66FQuMBinFF46DDMg9wmPxlYbxRmqGWK7NAqP5E0bWjDvSOWuqBM
alDQ6PVG+MA/h6jJt/glAzNuEGLhBx9D4FMMgR8KALf2mwSjedUYXJ+PB6Hk6OWo
jjp4dau/qDFNN7oeqe10DfpoHY1nKx/T2jO1jYnIhG2Gemr6s0BxHgdlh86jEoi9
4+T0BuwCS/hvmn4KOR/GTfY8L8az7WA3OKX1XNRK8R3BIiyz3K5sA4PTUdro7xnb
ALGW5b8NN/gnlnYsEnunIW9kKgN0BYnjgW+EYiF7Y+0WpGuFDq5EB7sn0Z7cxsQB
zKKkhK68EDO2bRMs1qWmLSwkGtSdz+cdpfCLCQhf7dw5x4IeG75+i1m8wP7joZbi
5tYq2ypC8kUl+glz74Rpv+klXiIytqMeIj/72kNMghu60I9BW/jSmcgF1Jde+Gzn
e9yDhG4TLZ/Fjdx12/0/ZPia1dw/t5IgzxGLsH2CLAowwBysSGzJFE+TxYdRhKU7
7yhx3zX3ZJZFC2mu071+OTSL4SGTv+zSrH4fBrTmf//O9GFul2bcOsdfawfTJCDk
PMbUGhfafvRX51qzpPxspwZya1kO9Lot8FIeMKjYdqAR7NAP0VpUGtR3c2sMY/b8
JbFuIrGPnNQx1s75yGedxr/8oEwBzQmGoDrBvZ+7hQPktch1VzI9as3XyiCRINmZ
yx0YdiHf7aR+DvvWIZogDNPLcUSMKTNMfUQhiOHIfCkehB4fdv9J8pfTmojUiQ9P
lL5rbJahWznN8OYEbeWcfWXzsXm+jYw0H7ut0i92NUizmip7pc4EeYkZLbdSQiGO
736bhydNm3FlGUB6VN8G3QpEjmbFaZT6A9MLk+wqvgOfNgidWWAEDX0ODuNaalW+
sCYlcADS3xn95D8bp0ej5O7MMENnfWrXI1PSQ3bc175oXFUhqJCpfHLw34yO8jjG
snUkJNk3tPi+jZGv3zIHNAthQbNNi+ytb6v1k2LYzgKD8gnJ1oFhL9Hqn4uT4MKL
8vOLvGZHGi3dGibG+ykCPxKfMyZmNrDqCjWFByoVOx1MZmP6AvQ6rvBXs6FNwyME
pSD8ZTRd1qoCw78jvtgHF8EpF5cSlz/D1exUAdh3VlgV3C67ua03Esg+yUGpb8jG
6xf1ZV3Uljp5st5I97np68/N7FXdp4ttJJ2Q0PmQHcRH7E8Yjz2ns7AzmDZg+g+M
k8gmBFtfAEj7/KBYpUsj1bNv6xc+Qt5qpHQduNrNAYubHiyfGV298u7nJOkkNYJ7
A2Zf0JTo1dpurX6BT+Bv0/s/0ydjPm4Zvki/pR1rr1POALKdFP3z3UxxeIslddZb
UTJG4nRsiAViPtRzplamb+IZcQPZM3BQ2/n5T27XYlcZayHDbjkIY7LXg6GpJsdu
pounonA8VgB33+862YyYWbTG3GMLO77o90+6h3hMOFjrY7eOxpOON7iMG1jdAKNO
MhAOVvU87tnKlBWnT6AumepmWhGNpUjNVTH6iiS/gE6ceI6mtFNOvmv8Rfv17YpM
SiI6odLJYo7s4LCoJav4zRnCEpHqg8giTZqz3rwXzzV400t5QDkS7xdc5TAD0G6B
Fr+4dLNBU5/srxzCRkKz6PQA3NQNqgXr8xKV4UjaAFOOxmJwi1IxpN4U1Iz03HJs
EDg5syWsu4nbV9UToJRrlWPBxY4yEJpfq3AghCyJCmPfL46Ft4T6enrC9z9oW32c
pJ1pIqyofdd6j4bJu19O/asei/9GIk71gSZTo+PQjKk2hiQaCe7hzZHJj7OREQm3
GX/Fr2Y9xirTN0XmnTPfuK6xLQm00PuMUqPNUMcKk7yUIxs6sJdnt+w1AKTxnMLE
cOTyMggSMH9Tr3Natee24t4XRh3ElVIUTmNw/L/XmmGQ+1nvdThqi1zowWF2KWK0
biEW5R033StYDx6ZrhS7Gx3yfPDDzE3YqIPaNv2w31xixzBgZqN5Odiv7AC/jUmt
MbABab4RZgOtiVDDPB/mRtzIPJjIFFPoIiXbX0s0qHLqKLfYAXHeM96ztNdqHBTD
oIfuywKO2XrhuKHe7EpPSg2x5uSLOvZvJC3+AFARhbKDzxpIpXgN0YpsZRC4HiRc
NpXWOr6i/kVRCICgsmO7p/kvjWssKQQuqLG/UCmb9LOycnVbhtBIzgE2Yo6TkfGz
fW8plBUC4QtJEPAkeak2t2C0mEuVlzxbH7VvfXbTsWTO/4hP2Zuw0luq1b4Quy4d
jf3EX701mDZKckZO4zw1/KfCWTYHYjjVHpeZklDhpAdrSxjTRju5bLRJMlyiHruN
v7lko5n9i3hFY3iQ4M3dDfNfNUAhV7AudEnI5VGTRTzTCwodrbzjn4/Yspn5rQ4l
1pDqa90cGM/wltX25+G0qcKugVqmBPHkPtMFQtrALrDkhg3idaOWdBwEM1MOVD1y
ecZZWy5GLhJ8HmPi8oS/hSlOt5pjkr5+WR/DEBOeGpcRYfLKvnGKC7YukrUuKiWV
LDOgKSlrUWOk92qkHHicJuTG75nR0XYaOCJP1WOJJAlQ9y3Ppx+RFpOnVRAVWnp5
6KJHORjcAzVVmm5Pvaeuv5iGJvz5rNBSzQPg7WR0TXuFLusLJvlW/kVAefE5nP41
iMqWGmRx9fV3uHTgR+GAwROrPlNdOHLYNRc0bfOma9J+X/gT+pFMkWwk6IJs4MA3
PqrwUNvgYlPsceD8fUDQNNLUzg0KxBcDI5SzVK/wwb4CyLc4e45vRruqalQ7mT+Y
E93AJdnPRXE16A60cRaPEbj/zRwdxDUBRve/KQYJvf6/hgiHAnjP0KOHtaHn3G6A
nOPSbbZv0tuVwAQaGQ0IIB5yYF0feB8MF2w1J+WrHaRacKg6kWReIMrRV+9KcAe5
BdM/HJjMZT3IC0z8kvINIc6nyPv5OL1el5O96gwveRmpPwSHtmqu2tTmlAxVxIij
IN2kLOJ0dDhptw8wHV6JaIazuhTYIQyTlakkuup51XWxOz7xaEWeyXePHNAQHdw7
NDHxW161PfbbNRjf74gg2V9F8o+cAEVQxrB3k6sPD3ZhAE+wuoWdV/Kq9XmKFk46
03iHLpJIcBgssRxZ7CXlpVCcrGvs3CMArVrlxqer+Rgwg7yAW/Sg73IHO2xPHjhz
BQegTxYrKEnQVSaz3fNC6ECU0hZRhZ4ylvPsjCZab9qYX5eP9WQdF+fDKZ/1ivuC
TJSIEsHYSsTB7+wYSBO2x3HYSbQEvTcIJv3f13/SLH2ywP7MJe5BZpZoWtpjHw3t
RI2ySOugRmVpjhcKBeEMeCAbleGTOB7Z65WwDb4UImVkIyWFYigacSNhbAegcwlN
Hi1toRTOGhz6Hz+hru8dJz9NvqwiFxMoTPJKn8kE7z3VvbH0k0TMijy8qY3rTtfH
6d31pS6VhGm/zOmorjTyIkHMz21/2KCH0FfFGmYKBFACx8NBoSVTcNSN8AVFcNuR
dqhLZDYiKpaSB4lDRRDj1GyICCJVmRUDYXAAGb/GkJq7XTl8sMxSOZhFbyV348hP
ksTzZoSHoJkyvqX4Y/ZmjUjJouUbpIPt18DUlCJxfW8CYm2W1OWprPn4nWWiE6R/
4n+6DNhn/R9XAMlHgNMJqY6r20cWjEJzZ/OnjV7S3MShHeiau70bjjGF7oQ+7mPZ
BN8wZDGQxQxcbvnBJCF22RVuCNTXwsUG4XO0wlpVaPCot6vbnzqyA+44PkHqNxCW
VTG9Ll/Dh/hb+BnFbYXbPhMVrUxT3Zbr0vmAIgiCSUzmMp6qnNt/+Hyrfcgcx8bm
+oYa2xMcZ9EI22QM+06YzhpyfxF8kFmgHdlWXuBrG3+WQQFQmIpahFve13Q9W2sq
dWAYgT9OxLDgv0+HG9ASCTzlFw7xV/TZGs8d7u2817FJVSCRAdiiVJw8nmSabv2j
H+Fd8nAOW1M4aGuKtSxQAxxoASjJodMhn0mJ2kgyrPNFTRCIx9G8hld4Rm85lOU2
yhoJ2y+XxHxXNSbuT4mCQPGfZk3kWseoQboZifcf/YnYO9FKLwTRzLGiV3yXHV3L
y55CJ4dOloJlKq7w6kvSpiQdR4ZxIBzctK+GSEGU6/zeT0o8xztEAuaNe02mVTlk
BQk6sF6TJSN62Oo3SeLo4r00HSLu8R2wuxpJj+Kb63Vt8/ANWd93ZxfGS56vaFme
IKUSY+g95CEPl/qrtAtDb+TPckUWFGMCoeTmvqAMbHWPFpzY1150Mbb5aRJ1TABD
ZxdDnp11LnjWuU7mDIuS6lsweIWpJoVPHEZviA/pgW+o0t13EMhLYFn6XMmwPpnP
bcfBS2OPAUNY0LF2VaBl4vlsJSiLm/kY9Xlcptea+tjHMT/PjkhVCXUQLsM136DU
rCyvde2xOgei751U+e6+RpOd7K0tuK6gWzQygkeE/JaH8IWWNlnSsXL0/TuFo3ve
tLwLtCo9EbpS8Igp1vnoW/MTOwdBaM5MiVi2fmQNVGHtRjU5BXQkUfijwdHHggtB
90YumGOfErnHe1dRW7i+k4UDl5c7F2QZ20eA394zOKwIBhwXfuKxI1SBc41/wvku
hyk3HTlckHm2mjJka9HpSkelESQV3XkPMhAd4GqR9RY4hondJqyt5ORCQ2/Q30G1
PaEk8eaeImz+QSt5NDfBWcTYI0cbcnNG8wUBdoW+U35aP6o8OF7ncy3tGDNZNq9+
tb7M/IdxUypwXUB6/+zL2ThotVEcY2ieSNuaEH72BrIV9p+4PQpGWzKAs5ulQg2X
kxfZTryvHTrzbMNkRyQYyg1ULwDt1YpUB5ELthkIS2WGM8Z6/5cXYL+aotLroALn
N8ZuHb6lnDrUldnA6RGyJ38muVe/OdzGWNKnowpe0girKpZHKcPGNfHq0DpSjedA
CFjWDQBFU3YUeDXk4nIeMTqiG8qAUDYOYgBHH4ZM5Iwbp84VwxboYQY14Fhn2fgs
yup+w9psOSNyDew2KU4f2du+rOq/C3CQ4Gym+gYZiMeB95P6sV3fYs6Owgjak+Gk
zsCFRxr0sDOFXf23NebH8mu2S9JPrB/Ha4ws2qSdUwEWsB1khM1EsnFp7F4ery3N
BOMooAtvSlUkDhrOOaTfzvV6nP1N6E04SX/h1Um5zh9q7ontaF4t9uy1ufYMgA6E
YemK3YFcfbTutDRE/68xgTaEycs0tvbBlhSoNYO7Eh5JRCzAiWJMgnEh5FEoP0KE
JXi8QJCSuGK2j9nTx5KwkiX97TRbBV1+lohgZ96wh9isfCJZbdWArZjnVVYpwraH
Ak3jsyV1NFYk0/k6eG6dQ6OIAJgQ+cMg/p+z29/SyzAIDli6DBIjxlAsvvaCkmIb
cY9wn+tZopo1RbTn60quQdn3TEb2ZWTB2rUI4UkmyW3HQoAtl4VuevhDpPSTzWqs
OodICzPMomrzWtnvT53w/Zjs1Yqr/tvz1b2nxH5UonM55cHAA0k39z4l902B6nqe
mNE7eVNcig1bOSxB1B7x7WVGnkfiimFZUd5n0gGUHqRKb7tDBxq/73yERrasFuxZ
BrB4Xt1/LEEihoIM8gmvugT3qYv98BV2u/rAdgbZ3VCzvHtr2BsCaW8Lg4hBkACm
Qxl4Vk2yf68aFJb0TAym7Vplg79Trh98OJjH5ajlDtI8bzKtE8Tkxv6wZWatEPbZ
Fz20CX7JB10W4wbiU/Gur4U09MWcP4nTxxAYNrDYTYRF5E7JBkzxtJ0c26h2EQBo
8XxqD3fZn9xh6LBF/gy6UUH5uOND00o0oJzcRvbJqu0PDzQTTKpdogkUoisImN1D
iuUl05umS85UNEY2gXRXa5Cf2jjh4qMl6tLYPLyULWrbpjQRmfrdAeBujvWDM2Rq
7Pq4wKIR0as/Ei3BKQoBrbyd+7CMt7L27HwMQPW2bOQck5SMo2z572f2U2Bkj8vz
0jPoeVhglcp0hYb+7JQb5D3BZZPK22Elj23LqRXyzoI4wdvbVrRikRE/nu/WfiNt
9jUyaqdRVZ+JZW6lgUoRuJNyzn0chs7vGYOtEQQuvr0kGXy30PmI5hNUsYMeuqAJ
FWsLeTCK3MvWJfQRxcRrmSo5sbXahYQaoaLSrXLaUp+EDfzCVQ4bgImvShEnI/3q
gsWTyqIF0zFJExmzveUrxHCtDuOJYdrShqj1Bvu9r1tuSuufGoxFLsvcluZ9Rz1H
mSFIXt8/oZlrCkEXpi5JIuzLS5A1IMgInjXF43sMsDq1iUr2MZSQZC2NRDtYd/bk
uP0JfuuW13Rh635NTF7uvht7MuAeGJaOTXnYWGzA6rYrC/T0L7rsTqz3z+WRnOn1
g9X15IPIlmADw6SzoVjtwmBhdFB85reJZB8OJfrT3Wh0GxjZdY7xKCHWNeIm/xkf
wVKCHnuGZmGyvbw1V6vyCAzCCJJIEZZ3xrmPMtQW1cvwLqloyR3EwnzuYmcd/BVc
7zTm/v8dijCJUj+sF0W97k7rrgaGpXy//k7Ce7x4Y3ab+jy2yIRDVsT8hs2E7vrI
y5TFvvWmMmmLLA7wtzX27rkGw316Q7gQ9anjNuXkbaUUqNamdpUZ6HdG9vs2zrSC
OQTQQtl5Ae6Txb0BTQQneiGINRcdxaWIy03rNCuokGDenBt3dixbfQJixc80c9AC
B29MwwEXMVPbORX5jB9jIhIearxTLxWcegZzyD0K6z00lSeI8c81UlwsHnK66PuG
Tm5/i+SK2EUv4UqC04ov0rtJf58V6IgJvc/UWnMpvidoAT5geM0mj541RFoeR/ZA
w9XFHfdv8mHjRvJAuOiSJJdU+fDUDDYNx9U3j1zrxRIh938IVVJp1vaW86YQfRlV
HMB0L8kytT3buBgcOTkaMw87LSAETIF5FqHM5gZrUG7QlfPR0jTV9mcMqbpvHZDu
D3QpMRLiPcML6INs8mQ/4MW2YC2ky4KLZdJfgwfm1N9uFUYzntmns5BW56nDhK32
C79Kqbu0AsU27PE6XoZ8WFUJvj6SS+vUMwl4exbL5gozH3vxtx2Hy8LMfT72Ub34
wjqGJNJ8W1cuW9d2hnZHsRHJ03AwnWqGYtgcdbYD4m69NruJpHlR4gXOnty4uuqc
hUINfzd/6LXRflpQoKkvzj1Lr4m8eUVxcLlHOoFlOxSvzPfymLh0D+/JMSZah2d5
X7AFkUAN2RJIiE2OZoEsb6A2XXMZa1+PYA0uivZwzvOCG9B+Q7xdALcZg/N+CUDh
GC/pURAXGmkQCbJGE4uo2RIechVXuopXPmNe1ZDk393mrC5FygqWkzWAV8TnOpUN
w+rZruhlJ20cFBaNfTz2tczLmUfbfQeIN8L/LSH+TBZEVmzL5Az9ik6zWfxYq6HJ
TiBATy1iP8utZnsQGYmYz0CifCZtXwXfGuqmoUK/HW0Wf3Gs+cJyG9xmgnZL8pzL
63QMs8ugornvI+j0QqgDc4+N8BmZtLMx3wNXe+H2QenF0KeLb5Qng7FeVrDLfcqE
cbtGevCNQrq/MwIcFW6MtIhS5Yhd7bZ+lSPhi4oNZ2LbAQEWlmX+MB+ZFsS35JZW
kha3vgn9OYvCtKTG9UQ9VzSs5YvKOVJC5OQz1YTCBU0yfLPbymSvr5WE8Kyjwa+D
6xcbZW6RhoSOawY611bWChw4EayfwevWTguCjVhguA8uA25+nMXOo/yGo7O4hSbG
sOBrF8diYP1p1MxpurDUjs/PibNaCz7TquFGtnbMfhEpW3RFMMIJr1Zs5RS+kzXZ
6O+Yhjxmzo+GkTHRBvCXudaWijUGcsti6vVp3twQXVNSwpjphSBXxk9uBFjot7DX
NoxahL6R5YLqo/T1GwULGR3iqC2pGU9JO9xndop45ZlTlF2Ik3xTkYPFx8Ce2Whd
kw62LVVRBIW1pixoa3BCQbhULIyMyxu4nvkoMTAVRA71TIjjLxl4ZJbpBnVBGUDB
djeuGGZg78O/LbyC3mXcN+ISSEhrMSvb88kmVtN1NHyk0F53WUq77lvQ+PFAA25K
OdeQ0kiYBv+Bco2gOp4SpYwMRGE4Krd17bfGbK/IHjj4DDNNdj2G2eYyxgVtGJm5
c1SPAx9JIrPBV8Zwa3Vz90GJe4ms5Lwc1GxKUZENB7jPwhbSRpzXTtsBoTOlbVM3
3nNgDmPBU8Qbpbx8B6N1w3ztnR/mf34J9kyHNlY4i9LgUsRpe2ghDE6JO0Ot+LIR
mKWBrCuKCxUD5WyrDeNjw4+qkIthXfgq1bGp6kZ70ozMgcUEKJ3IZBS3q3868RnP
BUlNwa3K4n6MR4lvHV/OUgkTZhZJBKZ1cExXNJ6IijsuHWTN8ul6QhK79Txug3to
ZcZAKGDeNb8x/oiPHYo1uTnfigI9f+ZkWHCfnzepItBtpmkXwpZuFWt4iwh6siXY
Sup8PQzk4N0DM+bgcs7UzpLvaUJIIiNOZgD8aQasyRx/NYgSPCxRGYB/Kux7/tfo
aDcLbyUw503SV+5nYxRxm5dSrPN2oFi31fJAPHoh8DtkZrWbPEZ1qMW+D32SZpSF
Szq5WN2A9zRKO4E0IAP6gcFWntLd83DVJraKrHdKJVi9KlFAJVYldJtUgNujwPEw
zA9E4GfDqLprj/BeE5huR0VhyBR/v4Xb5YMTQx6yjM+Wb0zPXi5gfJDISCwyWxDT
2UtEKkuAqx4GifHvvA2YyTLQwoT2gmKTdlPbX1tQASnF7W7EiJ5r+BjraZ6Gc3Aq
/+dnTLpZ57PZXAhP9yw1EukJVeVK66idslz4npNljAu/pJxFC2y5g6qNOhI/Bgzb
Bk++NDfv/qh2wZ6CwFEVhW3c82y5PGopjyhyp54gyUenJu35+oUWX8EbNKpWM28R
+fUBsi8RlUvIe15knpaFl1ByxEJvJAasS7SbzBgZ5edjBcR5vnjv8WDCChCxyF+D
quymlKsVjn5x1ePmkVghNEkEpbFWv9xI+1B5olSnjrDYYqzrCJwNgC12JHQ4hxwR
yXGLtkGx/u8tlzSdhZezvW4Xtnyf5XIbPuZWAtwFGHNmp7sm1W/xmT96buDF2WKM
7R8mXhqg/pvoUMsvgJR+P/jMXrhE+aK5C9exZYf0wJadLC3+hUqeMmdv8j/e1X/w
B41AOf6/JX2VnryIkzkCCmWn2jeWX2+099fHUqjFUTYqiQjPlXoI1EAEn033lFNa
T9LJ6JXLGo5jgIjZD5zXDLhUoryxniR95DC4vKjt+zaHCBY7reJ9MULQf7ol+8Yz
i52zVE/KByIHQp129f3Z0LUYbXmLNRcVg42tbGoh9yq26De2Qyq8SDEqcGYTFlIP
5cOY1TW6Qy9aGwet2mSkixLbIDOjqkGKvCHCgbttBeHkVMHQ+IaCsA40AQYy56nK
xshjDUjIDK6UtsqfF5pjVbE7XLS1To14muCyuNr1qLG0g0KpPyI+hhkzaE71eGkw
Qu5IXpkHBjNQDKpXAOU5woMu3BA50xSIiMP5j03iFP5/ebv8PwISNlGxsPSVm2cC
5AHm3P5hbVDMXbAaAacyT5cQ4C/2tOMprP9HLigc9fzuwThWphvsGBVdbwCw7Ymn
3DbomTaKTqXJTEXef8dTE8TXHBWrb7aR8qBPHooK3RvaqZO7h5UfvdejSUMW7TsP
wGE99N2Ghrfq0D4V4fS0UHVqz/utzehgUX/Zu8kbWzW2ppmPQ23FVPi8Nly6eamO
HISKZ7kq4bI9an3DDhQg+Aca2Vc0oTuPYCrP+9BZji+VJImxTeeusdqaAMWAt2CX
6Ye6OI+bhkf2972YnFFIHR1eBERwxtBOYWKVGXKWdnLNT8BK5ZLBOnN2JfR9in5W
3XZmG/Bnm7/08sASRatCZKjzsTLhk+M1475cLrEtleBuf7E0asOYtLYaFpFr960Z
YdLsi7+DSwAIZ1HPP80xSLHPduZGVNbDP10OT9z/UP0wkCeWOHT4wlkkZR4UuPJv
AkuPCsLxC+hvR3oYUmcy+ez0OA1rRP2YC0L2rtCBkFLRJwK8xJpB6K+nhwWPBwjz
iEQQZd+rQORdh3xOJQbtrjJRyi6/MsZJZhCfDL+ClQewo5DjRzlbRoO5jSZgXExe
7l019EmhueL08oIAgw9QOYfeMsQy+7qXkAVUA/sfteqBDV2ZotRDjt1OsaWwyZeK
GvbfRU3PGQk0Wn+gmCstofUw9hDDQVDC+jn7+HBJzQhynCUw+OtEm3WIdLQ/0ybg
cPl7QMS/oDKICXZSxrTNq0t9dxUKeIwaJez+GzZenovHfIcCAozLS2Uen5jyahqK
qsMUsn9pnkcA2qouTbxCjYqL7H4mUEBwYsrUaeLRAfkmLIexx6RMDqlLdOsWRifG
ahdRX4b0ct6rVR1OOB/Y0n7BMQB1YJinS1EEBkpN9O6gSU39WOguDnGX0tU78i4Y
DDaJPWEAPyvqj+RMu62kEElVYG+AaYrk1/lFzVuGNIvp85hfaLlJZw5IbGKkzdM4
pNDvwcFTptOTpF9bCteISR7Bmniax4n9vtnOebulfiDrTMogV+tGc0UI/a4JGSh8
Bq43eYH5x5GM44IcRf+huJx2XpVVMAAxrd3GM5dsHuuBSQov0EpTsSTW8Cq8O1td
RtCBLsExJBDFNrg///S6If1wNahY9ktX8zBbmRldadBqMTKkD1IRlzO+T9wXtxBP
SZ1rczNBHXWE5eniH18NMWVdPaFWUGM0UF7xw5gsW48CHqPYwcRzl6vOd2L7Fo2V
cM6jw1b6oCbFI6nMiWd2zUzmUKHgHCGZwwF/+O2Is+JVsxZ8eVnVrgf4v4wW5Di2
AATiBLVQ7UB80Vqt+u+eaaVetAE9SvjZ0AGCth/MsKzXdOCM9T76pmQlqWbvfR+x
z8N0y2MtZ8uhg9hzpp79APGykgSH+J4ddnZJS462GiwnQSo+etuo7MaTsOhgZNFw
6QmFk8TDmWoWnfp7nRbkMsGYZuOgra55uuKxH8xDYTXgNSx/lKNiOqZw6TfbdnuC
SkFr2TKt30U8U/e6SFjZrZpZFpsDIBefwcZGfaTrQo+j1gd/68eCmdU6Kd5CVRmR
ljJHrMuhotrivVNEwqMqrV0o6zU0HeofQF89l1rxJY51dQyPwMHiehYOQMkKjlqv
KEJ/XtYi2DYJj5tm18YefiTkNpJDQ389B8HeXUcLMdNmWxH6o6Xzl8cukyekW+Eg
eaqaUAMKAK9EsFemEE9GFy8BAhV8CEzNy5wIFK3FXfOM3nAg8ZDwX6138kKVKOIJ
Iztn3NkSfd1BmK5Cf8oV0nJg4HPmvG+TXstoAWsXt6GPIjj7+vZiMftxn+m8RV9d
DYCC+jio40o7fyKko+3yj8BSx/alK+bwZu3rLDUQfHbZ6eQFxuOj1csEMeZ8uBPy
uQjQYAkAeij1RkodgiC5heNIEKyOssFPNt+pJE3dSSE1Bhq0DagYwqhNqyWg7Oj3
lnTIdx/dHRLh8CexJ6D/ZapMnOF07vqvfeTKidWnLSzDTxf4U0El5h4w2NGDGpCo
TvuRAxCyTNDaQYAiRDoHF8shCcK/sgQ3lk/U0JU7wKW21R54+uojvmVe8Tbb+gn/
IvEANB0z3nnDjHhvRo08IPI3NS764d90tsxroaIYhWkIXyJoLBVADSM7rf3FZ4QX
sjAwT40F3mBlQC1ZlioQ2UI+H+hhL3FXQEPfQkHmqTaORstUfmiBFQrQFnsxy2FW
yF51/lkP1HqYjlpTUywLYeaN3XNJ0wl4jcYALvNId5l2jEeeb2e5kujKOHhWn3ab
EVVILVP7RVZMd1bAzMrtm5SxQChI6qZfZL6qAAy3OOZwcQLg5jKr26cRh8vCDYXE
ZPGfWTEX6RmfzqllyZxf68egRdRrHkPvnKbpl8TBGnkTQNCsICHPFYJCjdH9iIBp
g8CLFUMyuVG/Qs27TM4YBonYUupQzRVxCDpEf5pP3hhSPrQmHWjFzctYg5HFBl6O
sQc/V909i+6ZLOlsIf+0T2fD+X3sIV4Rd1v1BNQUXBG+Mvqn0jZJFtlZkQtzXjvn
hNvPv+BgKQXQmjjbcQtAJO8hojW00270a6/NGxOXBOxVh69GpKZsmCEhqKI5Grq8
vWKjiwbMe8q7Bo37ok3dQRTSEOOaXfOVFRfDc9FDCfuOHQget4Vuj6UxuK56vmSY
5OxoJunoDWtAdIX8sLTS37LhTH06XluHksIuG6AR5i0329sMUM3GrFcpTJ/EuKaW
3UQY+gPMU3u0CKHCPea4eNGuhY6wKSvjTOQy5HgrZJF9nT1fAeblNb8UnZtQPfWz
shfwlJ2oezpTOqb6XuwgPDKq/n+0L3KXmHxsXjgH4KOGV2ksAjNvZzZsKz6f6Rbo
MzAQla+q6zKeWmA/k0AuEuSVp0ccW99VmuGwSpZen7muhcXvZwq9LVfYhEP0LIr0
EAIQpsxK7eA1CQHNW/Xl1OjyB0ROxuE7BpuJTTHkWMqIk0Uho2emARkhhH6nmCgY
+SBp2w+Nmkbnwctb0OTnR8D177kkGcMV14JL65HM8QAeV1U7YpdcsGOGGXDcUsO8
zeHTJsCm1Crt++kkfssSyzPsUGDe8sZGexBJtFvNRLV1RhH+jURyD681de+UOiaX
4w1mqo60zbZjjhTY/rdKi2IShWeUHK6EC41krFVIleO1fQKfmk+cuUkk6SoEUv7l
0KceDnCUYMIaJOTWl7ZQPMaeHMRGrNEfB6aQWXVc8pd2SyATeC+s0uT7zW82QDNX
NvF5oVZROa76L/of2EZilhotUAw9vr7LWNae6gxd3Ki6j03tYsZZzlSTY6Wc3k9Q
mWa4qUSrAyL4zpfmTsPiCHfIynx4ACqGpGZ88mZIj1oHM8oafUOC5KNT0wxPL6et
Nxs2c0Yh5XyC0nqCtM3uESeIkTZSl/kOSj6PJqKYQ1Hwo5lfuV/6cHEg/449RXNO
ulMvhylJ2Bre8KJOCUKMAKdf6U1dhpE2njk6RxhSHXHvPGbhdvrg2VrQyJlBdwOu
0cQfr/6ak2+MUbKJ3Se/z3E/iRWcTiXWfzan89RkXz3zuYde7s9ZRxw7eBlvECe9
VdEYJwHcj3CgGZY3MreLowawnabtR9rLDf6Yjs0B4WUHIpvsxXFzk/X1R/uXKetL
VFoxXpnkhf3vF7hbSmAlHvuzaZCRVCMbWCtpYSQziOXxsHDrrm5DGQuZWdPQwAPh
mgHhuobBGSl0hGpVKITNL6sfmzb9zKJHyydJbVmk7pgjFy7Os8de3CWZvAb9ACwb
q/oPvKuAghH6c/OOie9p/6Mby0H/IWzaUGX3QRUbaGXYyLyCtQ4gH5NkZzwmkdSp
6abg0TFCs4mXMkLkzdcuzYOeftMZpDgSWGQOBRpsY2Iz53hdtcJLKM6l4m8I7o12
NlO0E/PyNenVc+9iSyr1q2atbeIqYtRHKfS1gggABbs2wPVvZBObUQGe6MTOYh3x
lMGUcXYFhgbXJkVhNHh4xWEXB6Xl/Eny3N8m7Y/VwsEyD8mDbdLuvoIAFjY0GgDT
EHL/R5AYdF7k+YcIXfbiWdwAXcUSXvpqgwjOcMgMaMHtOK/s3vcA/qBAB6LJ5BYS
SybnYiPMCnHHDdCm7KloLnow0bA2qjOXvRRjDpnlf+mh4TCy02CpYu06HBUhsuzO
fpQZ25wOHg7yKwAPdT3RHnSKs7rjYn3gS5jBob08EpZS7x7U/LHjV1qt0XnEHDIJ
DAnYqrj3XSx/wK7Qvl4ZwdVEbGcUAbiiOLJ8b2GCpNjYAO3enNCgPybjOFfeglEI
ym1cqksKcEHQHwp/5pmYSnWHry8HeYFwk8CT6pZNMoxgeIwTOJ/MJhZCWgUH/dt6
d/x+LG/S1RP/WmIv9vLo99Oj0wPn2CMa7v04kPc1nWwBjGg5gt5Yjr4DvbR2n7cW
G+TgG2Y4mRuXgGPHdGCNyeCDIW3YDoBfc+FNM2My0I04E+Nv3gSgJw9BDn3P/iY3
0PnvQZbYNyWZQdwuHKKTaoC4ZySd7NglX6Trpy057H5OYGDSXnpNnVioQaynyqQv
EyvbQ1SRSTM1eKoU2GLS9Z6iVtwJjBNHDxltkD703goqMrCXxcXmX3V1VzeukECP
OVYxL1tVt218twPzdX0+51cXNVKpFf9dbypMD0rc5Mia5TL3kklXtqWGKkrO+8DS
yBS3DbLnsXTvwkOmpjXI7dkEzApRzoxoZ2hhHW7fPKyT6N0sgoR0zmwjIPAcyc+3
VTyLedoTszveTJs1MCEzZS91fLYCC7SeLWlzm30cbYymve8fE3lp/TIFE9zv5pcT
yvyNmeINbV1o/KlT+H8OxJWVkwnkfEbBPjHXQHRAonbHOYQz5drHacJsidaJc119
U6L8k/40uI99XuhhRiSCEgnxjrv5gA4odIXj0GKMtR3FEHjlXqYyXzVf4ssvaubm
7ngnr7V0JQC+PYE1I79X+bV7s//COBti95HXYmq1HWKz+R/fbluWukgsDEPq3Pi/
yLK6G7U1EY8IvFaGtyCG3GXc2gmERByh2ZYdkv0NEJucS5jE0KqZjuPoJoGwIAQg
ooorkem8eGXIXIO28HhV99oSN6R//WYSIvDk7Afnw0rAefiLYuZpiWpC6m1AVeIJ
dLQLInkBLBUxhJFA7bUPKqiY5KdH9ge/d9HRPu2n6+iTLSmpRH3IAl0RaTraAgPJ
lpOufwDBm7dzofekpHKmi8z+fNZQhi7k9w1SlKt7kLiSm2rrM9hkUE2Ln83wS6qH
h9BJluB9l0/YBkPsu95ZbgRx1VMb/dLKqZb35PbLnWYngibtU7cFfrjX3uzZLQE3
JaB6/UmdQOhQyejMZT+omW6XMDOUW0mAvlHX2bJFGgRx1s1BMKSGkI9fuZ2zDHt6
mzZ3EreNL6+1RqD+4H97oCthgoWLAD1BpT8lkMyrVeWzQ/mY+AkKGMRwtId6zQYx
sZbHwJs2HLEv3bfRF1FVxCClUFqX0Mp/pgx9OlI1UaAA5qEBF6AsWfyctrD+lnuD
Q2D61HxMK2v72knjNCVDxUetXsnorURlBRqG9YAQA2vnDW0wL2cG4f5/T42+7roj
nbmbIdHF+ED4P1KegDK6oJHBrr7CncFMInlDNNX+wxwpCM9vOu9rECrnvug48I5K
dNItJDkU3toWBNsW8pcns9w1IyD8Tufr1jTdaAvLQEws9A1AhlXc4YAxdqCsRRGi
K9pIcacaeeEi37U6saLZCygUQzgKEIzenArVgLSMfvO5v4soV8B8WWyxJgKE+1fh
FLmTsNm8l8k0zvRC0VGH3sKVr1m0Qlg+S2reYH+uwf1YA2N73Ztg6y7SvzQiffaq
jQPk6xy1PemhRUuQt8KphgLA0x3OsxkWYAHbWZvKrzweAVv2Bufjy8Xk4Bk78Utg
+LFaFThok5SZUfz6IQK9p+yI3Z//WH0biZIJvbV9SGAHWt4jKYfRIbS5c5zI7sMB
LXu1Oce/pi1SzuFgFkCqwuAL20TxeAEt6hoGZvKIZTuciwW2vLEpdoijkFGcxIHS
9FAaM27z4/EMSpZTRPhNaxSanNj80UiaH0eX5NGaUyC1w0h/jd65NYxgPnZ/nSsC
Iwd4Tivz2aShdf0fLq4mQWWgVj2mCUhPfTw7wC7v4+Zs+3jFmKYsjY8lkOcL1Z6I
F9KMM1PRw2XPt6/nmr1SJDk6BPjCO4U4ayrNLK9JTxa8BBJ1ltYPb4qy+5ZKYo8f
1OEvRMqyCIDPjXA1/kPiJIq8eGlYuDE9KLLdWPE9DznEg/woDYN+fAUiP8wpasqv
CEIpzm3UFdtrSa6jdxYKQMAzT9TGMLrBbJSVb2kgVpgoJPs0kz2nxorPypsSFVRH
glXWv6uxlNWyokr3gGgz9X47KOIZY76mGUWpBa7d4uP7qIM7KAIY9bBx8Gm4DyGw
1f61rFaGXIJZYReuG8Dtk/NxuSJKu6xTvlXd/vnFKJ9GBz6eoc73pb9aMEK4HPPt
NIHNiOl0kC9ywd99rodSam0uzRfSmwF7ir23YQthogefUkZ8TUgES4vwuo3FHQ8m
UuEkbtif2o9YIbeekLcTMwgoE0Fm6Y2bQZQEsL1N9FMSla08JqJJDpCOA0D6fwiS
pWLZG+mRmlka76E55zF/oyhkM4aym+B5wNoaKdyy2Bx1mP2cjSYTqmKEHITenI+/
8teXk9pE8SIf0Qc5Gg45DdT0yUOMpukMD3tFzpgx/pU5WbuNSQlTNcXaAA4fq3dW
BjVbZwlf/VkWae/9TpkSm2hWmIsFlxqQTs4efHWgY93XPEIhDikXOEB0SpZMt4Zn
tvx1W8P3MuFKu2E2lRHXcvemP8BiasdVN4ZMZ+QFHneQ3XPoSYcsIjiu+Ukwm30Z
OulnL5TT4Q8P8fOIUZqGgCoU0UA44uclGYsNufDlK8xIkskBNyNctsw9gRU0UEUb
YJOmQvE6+rfpBoCXx87FfS7NM5Q8krIWvgiB6JBhrR8Wol6K/qF8dnpWBdqndQmN
bzB18Fwt1vU2WneQD32poYxaMCrRzE1vfLIZjsjXhdmcpRJ4QunzgoLj6kSKl0Ho
BNikEovEkXPfZ2UR6wF7FnYsoJSMNgqffqZnUDDmeUSJmNZaKw4rtgfxECVjkRL5
en15fhof1Oc/WCkfp8+SpLApwilAwhUXaH4qIIaasD9Ph6dXyaJH+i3M+x50tGeS
rwDAgtjy0JGVRw88S1P6IvbYt/cdiM0fEfZkLwijUdz3p1hl7CAoRzyX1uU4+1GJ
2T7GZ/cQVlBH9H98SZDF1mxuHTu751ld7tPR7mNAnaJZpQqYZsfRgNUZ1iZDs5c5
Te3gjypGxRbqLXYostuXeqc94wJgFjOtBchZI1OIiSbDtTNzO/lXJUkhKGS2LaYF
cijWpwiUynrbQvcl8CjtSg41EGg0d7SJUboYjyqYfDLoJ3rQrXPfzcL3v38jYb8T
z627RInN2UpDjHEHCKuJfhtITt5eDxy/zNjhVM1CQTupYZCHooVFmlFs88HAkmB8
fEYCwp77qp5iub88x6N8mVblFDE+u7SIzOjvVMoOw7IheNd4/Ta5cT9fcQK+Kahk
Qg5INC7kKWjXqPxSCh4ZgD4rRlc00iOfN7FKptDKE2PZ0j3N6YVFBjkhfnBoM5za
OISA510MPuZHkLfpf2SuNtSIJ9JkPb6zk26ndsYcLBZAZY5NQm+L9cAaYjiwp0IQ
g7N9KZ8r99L55YE9kLmLws842U4+p7+LICHn74aWDpHMSzS0Z1tyZ4YkMWKQxtNl
tzWXR3ynPQvtGv3M5kdO/Fs4FblCTp1Ny7MHTJ34RRveiCSY5lfF+z3zIEchxIEe
1u8PZVRyYVtlg2QKj0HBkyCzj36jcvQ2jnOvyFwpzPuhwU6FLP7RQO0Gq1RAE/iU
w4zftCAT84ivQJ4RE3BPQihj59v+rvQZMCRDFXuWl6Ygk+KAelOWaIxuDzdfqGBb
umDVbfnHr1bbeZKknsw4pN9ZG5ekQrAGb5mMD8j54BqPbIj/RCxlH4fngOaR50WY
ur+V0W7exXdgR7D6IPzN1i9DwRfObIKDrpmwFXrMCtstT6KwaKx3fqofyTxMtN25
R4kwbse2OFFXnFF5vBX8dbSQeCtWW/USTVxs1SPqAe/LtVKye9fwIYBEThgKCvd1
3TmsBkNMGQ1QHRlbblKVzBm3RWuIK6S2m1lRppTKTrJD+ubVHApKo7n9g5tn09CK
BHEmkibj4pBvtEoamEAqCPX+kIZce1ZCtSHtMG6aswTpOOZY1UjsxuFXkDTrvRC0
hcokK/3QZbyGTIPCbFTYg/gZP3hODLKhZwnZhoPQKJf/u6LO69rdW29qsThmE/CE
D/uAcHfX1OFQ8pstOkYVShbLDvWl4nNU6Qqv2TNeBzVieBvxeJL8uaEDC3+zJPOb
06qPv0O1XNCs0PsKanXwJ9m3oj2Nlc8m4f+13TEDuMxaVCT0IhdjgosFYY19cqrO
0CSQrM1tbPZLDKJghIwgDjlXcJ++EjICg3ePArF/zfJ6r2QU+ADHkGYPbj+FvE90
eu65gpF+tI+nLhX5mUjjkrcqa9+1dY7L7nWOY+Xh2lFszUs16yK6WCUqTT2XZKrm
H33BRJDLRcmUg7S5t7YsFy0JIftomOOnZ3D9EHQpBU7m1QqjWVQLu07gGY6lwCYQ
KWgzpWD5OxwJkd0shCUH1YU3wVv/l1TU7QTZE+5rfrIg9s6LUDEHgvE0ZyF3MOuo
jMy+5D8YWOxTl/HMsSSH6nAkiBFUJpJBFEB8rUUb/FHFfOxm1SAfA/zq86Vo6ocF
v5gfe9iePEzTMU2v/KZLx8UpWzCi64Z2E9gbus5+80+tBXEgkFP7wouut8Hf5oRj
Lvg38GQSPpyR+XiLtRibu+meAEX+jBICyhHbPE0+BdoV0PXK1GzaaN0hH2go6z1q
otq8aJAhyG2F5szEMV1lQsAEmpnm8E7fwYNnSkLJ74yETMWWZgi2xu8ztafpKVyN
axoC2hoa4+cjvep/djepKh40KQHG5GcVkP89fzO0P9Y+RDDtee1vCptZwazxhoX6
l9OmMbNNWrB0NdLfRHlBq5RNQIAwiWbiYOp4j1ONFBH6U3X6abBQ42xV+PCuZsa4
+N2GuxqyVcLBnYEjBRCRkFYhfCPcQdIEMUUp2Ne2nWO0UHcirW5ArSzjIu5Hd1QH
eIPPV1FllvAFiMwqDA7eXuL22A/kXQb+0h5e5B23Fl/JqS8lKH298fmYeyBXo1zo
ONV7olIsZIvwN4i0Temf47gLF5SoNG5rf3iQ8jCjUE1mM6HsOVXv9pGeImthh3G2
UE8U/tQC+9OPr5R4416/a2UvNfHrWL+Zz7ImCBaZxZX5GaGQFmKTCqHkaPdB9EMl
gMAIORCI2xInWRM2NTE0Zqzyn2TlfeNUi1PNAhksSL2y53tTy+2C/wITyh8qLfGW
8HWoJgojLuqdpV+roo3Igei4ly8AY4DvlR7eujeFtK0AqTCqK2bG8f++ykaEuI+8
24VwnENXyiUvc/Ei9n7Dlch6l/+/hFBLa6IEnNxH9Zhv+YZYb7VuKGvQ7jS5eSGL
6XJta8mQoN0CqeD0sh12yd3Eck1GdJ9BA5Nk8NXRrjLgxcdHONA9T/rmbOYb32Py
WA/nXfYgdC6lhg1vrdB6D0vz/itne8uqwF471DM298LTEY4WkiVmTI1azWiyg4HC
VPxxtJj80t8lpa5cW8ID/7/aulCghPm39kyFarERrSO6fKShHviA1ubniA7NFlcT
ie8TM9SzQv5sJ6/J0YXt/v7i6Ln/C4mCPfFKxfPtF1t1yW5LSrjqgRuu+LCZDtdk
/oBPjKST/Sql+40hlB3jmcz5BNwln0WzS1eHsY9E7fxzeNnwCyGFzTMb1mfQZleb
qE+4QsTHeQJGo6eSFC2E4DRqHLeYTf6RVp6zCEc2rXk4vtap3TUqdFLGQSaslDX+
D3zsvDPL2haaThHqb+p4BSIDgbVCIwctEcQPDvGYdhHyfeVIr8p+gvxSptKNxO6p
VmXNzNQfYE6+9o7VS0bpyffVP7EDwdrQnrXf8ST+8PDkR9+Qq0bIrXA4+zClZNa7
XQpSaKg0tY1hv4o/j6fOTUfwhZOKxlT6bAXphG/9hxi+r5nhzkhrf6vZ4OAFB50U
JIXfIcy3DTQpcVfz/leD5B982Nl1oub8hBGr5tdnAJe2C5Yv9OIbOih+/GcjpIHC
bcOT5jibTHUQZGq8hCttvfx0m5XksT04PzMGodLKP3C+dCbcUdhOUhMRHpVIo92N
ypmOQ/t+ByzIS8djgl3er789zUwHS7p4i8K+1cFK+xtMMrLlt8NA7RLbpkCbBBf0
oKVAtb2POQKhmPohehr8VDlVfglCvPqFz0ykISUkSMNH3sfZhVBLd5kPJxBP2Tv9
b+eGBr/NfHDovcNr1opjJRtlkC6vC/XsEz2ZpzKwwIHCqHDjMZSI+9PY6GZjQ8Qp
Faqz46//f7hrBlDYNzU9Y739aoWCAKm+xpXnlglNg0mraaqDF73qm/64OvZxkJB7
VKIEW2kBqyNEqEgmN8NXYnxvB1IkFvG/eguGF/Ei6pY2u7aMZdClr6nZDofNClKE
8xc1IJgqKQh2OkUea+VVCUga5BqnT6Ct/Igzw4VtvMf2sPknYZXPfZcYC1FjxlJA
n/a1/sp9QPzyQoh6Da5zLNHGpz0AIFAoGIhGFSmxtN7N9dycYMykS85XmF3nZnm3
xZ7V7Pfp7N9ZjnK6wQXxPu6zjZAgA3kgJLHAygkwfYXILI2lI5fo2L2ku7qyZ5YO
bKrHMVgIswR88j2xxggtQsBFyR9XfgN9XhcbTybdPx6m8hfXIDtg7ACoiVi7hig1
o9kgEz2qDxJq9bax7sb4TUrJuj+qgxjIN5AXazuOWgManWlKdAC64SgoTb1jzPs3
gPVvkMR9G4HeKSF1tde/E92UYoDmCSmhYt/eITqs185HVf0aQ3flGUGef7sBqi3Z
XdrHEjfS13ivitfnQsHLR+XNtPNnugpCEI08HomSRBjp6R+vNWRoQFAAqCb5eG9k
f/elZSik1s7afluVghopnhmGqFZMQSFKAxa4bY9QGVH5CgkVM1yNFWABJKh7wbmH
TVbMD0Vefv4iwy9f3g/kU63xp45fAz8zGYi/xeZ7hVITH48IsqrD39vfizcl3+3h
2KBbVYCv0TMeZc6RNTVfgiI5m1Pga/up4F1VvUyuqgtQN25n3hmFapnWHk6jx1dV
TDJYqEyqNXeL5dfJzvEdflXlVfirCA5OxF4eev7fZCS6YWlV0lsfg5RZ1NwAUysk
eVQEH/Wts2efsaTOnQKKE/5x6oiPA7spNEFSTOSetrVTqKC5IWjp7clgaGwcw7uk
BkZ+hg/OgkA70HDy4r0UUuyoPyr8ZttoShuSXcP1bYbCPphMSA3wNZJdyPKHz3RS
fGiQM1An/JNrPhigj31dSCgPTbx2VaTrGL33bjvY5thLPpcemM/grX0R8ZK2TStu
KYQTQd5gB6GcbcO5AtABzzQ97HhDzvetvN24P0cyvjlmvyvUDLrMo0NNKrFnKifP
PNbByxJk0HNtnK0NzWrRp5ReVBB8zBVZuizfMKYLZHcQOyKd6fHLrespQgH0H8aK
9ARKpM2w6fJZKSYVlRoOagyeYSpHimOjqABwlASyX9WF+u9yg9Fwq43rE4Hey3FO
GWtFGBwlJAxIx1YRpXxDyA0R5M3v06gi0xQye77VXJNEi5K3S1YaMwKaoFqa/mNC
8/A9kQ5qnKRAGUNI9Hu9UnIiRRipnrmk48quo/ececG6rSmxhmhwsATONAo5GoEj
Zbrhkb8lXIPDL0nBYi99u/yBWRT3snbQx07KRI/Wq0iGe1LDO5Dyb2LT2NQESvl9
IuWX1OKpweIY4rj0vap4VKhqraQMJoF3NhXWVklqpZ77W6bgbooIitaPn8hPvlQd
eBtsTNbfdFz7uC7WosJEr9X9znbyRMxRkz/nL2BZLjq5N+klsilDw/fJngxEn1VW
upNvEbitUY02s+YcM3jCmHckg/cIkuIJ9I+pXK+Z7jZXU/7DskPUYB15liG/zOzp
dvF8vTHoS7n0+gktcPUOwwI997ALi069/XPM63TYKKFMmgrTNeFaDnERiVckVXrc
8thrwtKk4gU5qAo1VtlNQve05XPM5xwpju4hn5WH1kDutKEhIMcgIXvHQ2/1zesP
Vl5xz1c3JFrrZ60VIwZ7bkTlEJzQHpxMyU621sXMQDGq08R9d7P6sGlF1V1/x5ot
Ic4kZnzWBWw9N5yJ2xW21XLN3a7LCCr6vRTdWIGqyajt44H4dPgPvL0Aik4zdkmo
c8TmcscJOmG/DLPiYePP70t/77kwfphDr/lHt+dTcuWB/zEtQ851pdNzHdly+fgC
8cSxVvBfmbcNcsmWFL+/ZSvMCxIOVXYp5z55tfK8RhNTTsTGxElO/2xmkOXciPx4
cJhhff8tIDI+v8URJGB6tmgZ4UQ/hyfa0XJJRpXpjEjeEVSvMBpJfmzbXQarxLqn
sjnKm5mKlhHVss3jQu2X2ebyv56R7FAS/Zbw30Zd3+pwHpBSXBlOjcTgCNjxwlcb
vnrJAtP8SyeAgjJy5ioRoSvNjhFMa63d9KGDs5Aup5dWL7CnTqpaB4aq0hZmgt0n
ggK/ZUmCMg/2H3H02jTQlk2e6+2ptPdc7Uqn4HcxJgOsuq071nz/g7eIEPp5kgTM
SB6Rf2ZtD/hFtfiyQrTOHM2BCRFFyg8YW6gGtTRGvosS/46iXdcckZH4Dd03dLda
Fw6qEHFKsSDTvXUGx2LSI6+nfbdeHPh21jwE2j3SZ0WfgbrvZU4SfIKLKMmn+/RB
7W3CrSk0hVQaLElgScPVuc2m9GKDKcAxQS3NCmuSd/WmPAE16ndWOZ1l4fwSzAY7
ZrGTazv5zt8EBX5xAry5wyUPmvkPvqLl7FKCQ58UrfXfvXNlJUtA9yFm0ECGjAjZ
3mh7WViAycH3glOoqTpLVj9ZQDLZIlr9X92Uhp+arv7m7NV9SaIybMhq4FtjZlNp
MWZTKT7QEjjbaR1HyPHIxhR9Xiudl+DixaAPHRMIZd1Otc2+0UezuiU0RSGEr18+
kwcNBxbyXVx9Rx44VxRuPi2wUTj/zXSk9sJ9JXX2QzjdiUwv97ZjsgAReooeVALp
9oqLJx5JjOrsbaImTDSj6NIightLefr83uFh3Nie8He4qBRGDaa+R4sZLu5Q1c1d
atZEhSgpnlRNPJQ98NfKzddeD5h59PGneczuwDeXqb9SWFI313drWabceg58LQkN
fUa0VwP4tLX6M9R/IfZLJTdh7om0+Am/mi5ZlfBbPi/nReX+zhpJKd1qF5i4Ff0L
65oe18OLLzvPz82XX/sCFJcQpb1Bv6zWAOAPglbzkzDpp7SnG3kxG65d+malDWq+
pptI2yeQ5GlweV/WHI878QqYcATzFzoqQG3EpMmy/dshuMScrjKROcvylbiF77LL
sx6YTrL0NVCCXbw3qGoF2EZHAKCnjDwgNK8i/D0AtmsBcEdJdyaC0onYZPdcWrzw
flOFMqEV0KSKkLpX79s3CQeFaNiUBDeqyYRDUII4hO4RVS3eazKHaSOHCvVQ1RcX
r3ycPBTObXOswFdp+iWN3EDsajFqJ9vqGnqhfLJwxcx8gk4VzzxKJfaLd1kBcu8T
EEIfhgnWuKfbfkXOy8Ccc8+OnGRtsGg/p/w0/R5hIfNw4I1b6wgwY8V/XglMFqUZ
DtObDiHsizqAsmdOEHxV3qtZzymNF+rBegLXMrmwbYS3w7BrDnbx29akkeyNFdKj
H/zw1Shuv4AXjjpo/GvVzpnMiYkfR7XpO/XXENCMMkaVZmijsVQbRGqdUz41XRM0
xBuBXwBx/inFGIvE0eLIQtfBIRbXwO7wrlIY4doWoEY2K31C9EBibX5pn9o/84Fz
nDs7KpgGesJZndbbUALJ2l6r0o+PuvSN6UnLja/RQtzNLLCEQSQXftU/Vs1mSA7j
t438VlEjX1hDWNbbYJhX9EaP+FdLvCx+etbsf5OA3XgJy9mUpMLNGJiepKRyDX6a
f2Q1nCrPdaxulldOpm+uxlh2gwaFgo6F2CATtvyLgtReqZ3zIdrcdEUZcx1flVca
CoGbytldQlUf5OerT2b9GZbqfcSSiyJ70nPzn3XbuiEzA5p0jGauOh15r+m4sKw0
pIn3u1kLIlhghdHSlHJjSXXdI3JHdXWUoyGtVD99F1TMpf2c072vtL787UTe86f7
btQG0DcGSXAVdPar/fbWQLuHJKM0+Cr48orseq/DjNg2v9kd7ks1CljAErXzn391
qNC0mJZ/qf6bjzr0n370AEj8fK0ZLgmgVTdOmMcCQLXf7wjYlMmMO2f1r1kTeHGA
wanfJjkB8n6S2WkQ+qrshIlJWiQBwxbjC/RuAK6CJu/EPqT7n+h+2e++SPqMTbWT
laUgDC8eeoil1NEK2GytffEgVtQ+zAzZQaGeifNQStx21e7fOe6LnLW+7pQwbUUu
jxc/kh3SU1FD34a0pEzb0FJkcavZiRbSPLnwoQAUGrbNpl9nK4RFhd1mci3k4+M3
yQ0HYrUuGb2NVOEeWh8lcJXo/c3ncLlOmLjS1QcN4lNWeZT4lXt+qvT2Agy7RK4F
ktrleyqswmY1+A4I4PUU0cqa5nXWogYYFXrzlMbgHgX8ll0tuA/yzrdRqk2r1pre
W4uVoKc7fti6IkDj5eRHVQigqR1CuLizq5RCe9NkNTTxolmrgJr0gehkaYVR6hCT
L9BEMzkoJRmunwGJgATapX+QgEHQGa3D46yqVr8B2KYt4bJUap1gxyz8q731HTwZ
7xCipYDf+nP2zG3BRdOKlNjDWX2U52iUgAR5Zs/1K3atC0bowPXjMgf2euORf4cE
VMlnsIHjCqdE4Ap+zUPbLPAKyHmICpJjEGjFd3SaWRKH+lem9IyaIJEHuqhjYj5h
av8YTJ8lHzb5Tl537TJEcxJ++bEZTujo446kRBVj8zMtfG2rtjXB9OOMqvKWZpEo
SotVcujU/AEDGiELfGcUSrFpRGy4nhn/6hoeca47mrV2yAljL+haqyYtAfEKJxMW
yMQIjhfGNDFiS20YgHGfxma9rblHJcU20aMSG1Qi91ZQp4huuBGaCBGDyUkn70+F
zDFrF72j/dTGFAA+8cCb5g/jOviDvdKvxzBnwZHIR1gSEzNgaTz8o4XBfV0Xnrbx
k/8pTXf7au3TU3uS7g520A7Aj3Jqwn1T4LlixG3+GS4Kl6a55z6/LMOxrlFoWslx
SNugGDj0h8JxFwZsULxKYjSJQl1flySeyR2KFUZT8J//xBaH40/fwQBmuEUSLNcb
Ekudsswc0e2f3QJYliXjHQSy9dWg9E6GBi1F+VL+66/rU1df9iiDFa+m1gDNZHvJ
wlbUCvQH7jIE0IUSMqld7JpWk179RJQnKtXdT9spKXlQtTW1V9QmZXdBofiiRAOY
KaEk4m6J8580g/YNUgvqlAY7E9447XwrAYQDySkFP+KOjhsm5ZOTJ/P/RNYbQke6
pJ/xLm9VIA7AaA0/XnK3tXv5v+rx9Go/pOFrHJjWq2KIHF1PH3udGFjEExVcMO2h
d3hOX3LLwtyexnZvcP3S3KfSRjPkV68Mgz9SgXYGnI9ZXtMkBFWE1rFUQUV+JGEL
RMoDSRVQIJpUrYdG6PsIUzlfoBwR7WIJaxghUGsT/cwQuuYa42sewPhRzKz4e/gM
nG5n44XyO2QT8VYtevYzCIWHELYOaV/4kraYZqcJ1tc8ZZ4Y18k4ys8SMuPNbTFv
cUnUE1eM0bMoT3JWo5gCOjtD9zpmSeE2cIaT0PA7qBL0XPqnvBEleTm3hvGsY4nq
PUMKL+EjV9BA2Ej8xsT5WQfs6exyMItWuXuWYyCqtEWo7dmkHnhE0YgDhlfRmwlu
gJwMiCLvBTY9lZF/WoX7dxRgsPERL+xHTQqxYphO4i8dLgpYiQmzvGAnBLcPOFrx
R+J59HaT7DpzxYcQp8Pt07VoSMXTYYTKLdV/vKZI6RjmiYoJb2bCm9gRMZmCkRaI
jrLkhfBH+ASPv22KGqNSjBlRZXIhYtmFGdSr3wwx+hYHExt37G+pv1ItqVsERB9s
SYf8Mjlv/ypuRUvulZ/GoKfTb7P3Dd3eAbnwxMdhMgYfef0FbcR6vtrENbj8TO+s
hSEFdbTLlHSqZNhLS4bnpJ9UjzFSxj/pf/EhYGUAAXaOgwovA7uk0rH0j0I66y7S
86g60tO5a2vtc76hYtREeiaxS2QuAqUyFHQGDLIMPHPI7v4LsETe+eVNkJc0hism
QTVW3dLjG40E9QSdfVVHAMSWsdeXukAP6/CZd6tchOGoEyyndzsYPQUfaJtG+tUl
qEuFy+VYi3kyzQ0j1s5IP+brT1d5alXMAXZfXW52Km70TVeo7zqqKKHH0EgB85yH
cnVLCtm+jRSJocrBEwDAwdMFAr87MazDo8+xui62tPpcgzkW1FloEthaQEt8WoWW
ep5+zA/Y/mrVPu6ErYePbnzTlQCdnMTkGdOKJ/REIwYrGWxr7uJJU9CWXoAtS/0P
zIZ96jITDWMbEc6xiHrh4w32SZFdtqE5DjSi1hXh7Qb7NvA+HTIrRZ50qKTNJ04+
6voJIXENjbXi07RwWoGbqyYTu6m2xD4J4UWEIcSg00UYZfCtVhduZinGy/BqbbSA
3yzgzba7rYgTcHMvWFjsVpzCQwPFNqsMgY8qxSw/8BmR+egtiUtWKd+sHTdBDGSX
SPR3zUr/QL7A8gBCJw8ANWwwiF7KzBL8Cpk5YxD1U/o9/y3hfxuRrTD9p/iNYizE
3ApVqPGeZ2W8q9kdnZCwoEpOgg28esj0FnxIIyEFmTH4fh2+vEDQcGxxwFD5JUtz
Nfqi9b5FfZz3MzJeCjJrozy6S/KMK/pTqDTnszHGWT23uVxfeHWBFA8wxDq8B8Sp
FoOH0FytRPel+oAJprwz0oJeFo6VnVvdAuzREk4q7vY4MZSXLqXAwjhOqHAU/1SL
OITu1zBH1t353SCB6CWqEFT7dYVq0Pxm6P2MBXESsmie1eFkAtEhyR+gU0BGzFBK
7tKrW5uTM0gytsATCcB0tzrlvqk/4SEKqG0dlye1nOhakq8QGBS+cG8t6tmQiph4
iz6Hee3njKMAT8/GFlYyE7J6BHvPaqjw/VWufTfqpaw4zae0OGcH1AlQbeiIwb/V
aPA4K4hF3GkXQApz7IF29hSOc/UoZ8Yrbomm7Cb2FiHYkw6hYalMFAVlJYopjMsK
P2G8Vcw1pmI49ZAfyPnPGeNt7GrhBAZ77sZegCaNC0fqWOrCZuQLJ6lcuMfhmhDT
PHyzGozhJN7LKQd/dbR7NGv7SdZf9snYqMcMohGWTRHpTUHIL1IpOCUyilRaGtVJ
o66SOEi0azP3sAwiSZM0tI3qX3fdg5Ni0wxN3BrmAP/AaDxi6LIFOLLzlxhSx37T
H4CIO+YAW4o+Skcny07KsG/aYb0WPL3I06kdzeyYGK9D1v8yrb7NQk6jyPN/KvgA
DyL9cmWcK07eoGRjTs4amCLxUsNLBGn4TreWHIGabmbU2sWgePc42SIpL2htYeQR
mvoG/UeOGfC9Qett3IqnLL5xSYZWP7Gr3wQRnVVaSFLKmX3zvGOKv+FSI218nG64
zXlX00QSkiV/tvmym9WQmwJo34LaRmvPJNdD6/xz090W94aLmVNzBx7ya3NV/fck
otmtlrluI7XmK6J/AavGA/bLJ1Bm4Wcn/pNMzX62tnbVqP1j6y5XvMIanFf4SXFc
SoM5tyuYp15tQHdtFbScrJNqghb8SzgUSGo8Ptjlt3OxhfG0Dn/JLr7tEaOau9CF
3KRkONRrSIQmZNfbdMxCFIEWCVR5nncZNO1eqgtyhNwpOLPknwjE0dMdIBFbhRHv
nMtZy62cuw6mNOkvM0x9uAx3JvLVUgJp10rsAaqlZodPEqHuLDN1rAgD5Sz8x+YB
nXOI72kH3rKsUsWSU5S42SdAGCTHSTiEO5F9ewnJ/4SiBnbbaPx8bs/rTvFY5zWN
WFSo7DfDpYEWTbgV8oBEogpxaceMNRolwLtuZL7xkQDHMphMp2x//RQEuFm2v+x7
hotCcEavaFC/ofWP1Iv8QrdFmVfxRUd5zt3E2gYtb63LijRcb1as0AoUxFq44UI5
hsTp3OP2zp4JVHH0V4nHrS4HQ6TdzAjB/EglFpgZSpRkrULhtifGxiAWYOayXQHs
xWUEViqQTWKq2kYH7z0C6BXMzOb2xZ0awfEAJlN1v+kH6eTNY3QXwHhAVpLK0p96
z5B9O8k+skzJlJkQeTj5zL0EyVgROewMp1GfNyIx8JEySD4+hEJ+MF/KvJarj8pj
mfEtKwKqZ10XXO5VOI6xo7ZEn2DrwwQW1TDQS2e0gjS2d9k3W3k5T2xdhQfgFBne
fiN9aicwCGBdhkd9s2t2Yv4xhC+C0z+DZAk4FCxoWDfmXgwEMd/oQ6yhQLss412B
fQl+IOK6zRojvmw1PwJF4OqroF744jVkLJtfYWV5KeNlxu32dbN97ghpKhP94kk5
7DMK+2bu/xk8X5D0KCcKzIgfnZtyfFOoSlWiftJsE7zlwluqU8ltJUeJz5W7kf/7
CSBvFu7qwdrKkM6z4waluzSaNrRUMH8XintwKO2f/3IxqahDkewB666k+TTtRu7V
5z+z13t/ddjTUDG593iQDrlhYBkO5DPgnk2YoFjJ3WgyIELaPHt8K/qZI1E4ly12
J3fMJoPqdgAScPeYF+QJtJTj5UIeVg7fqgLGlvU3NX9uOeuw12IgH8KJfCUrwHyR
4/ts12ygpgMB4hkJv2oYZEGxjmqkzSiwvmq6j36WP2fhBKmlxvJUX6BOsddAGMA+
gCJqr05Wl8+ymRTy30xNQ2FHN2Fdi7OIwGkot+jbd7aaGocbf2pHUXrZTMIo2oHt
RKmeCURsnoIg/WbOcyKx400Ur9+5lWl4Wzi42dClqtDE3v2MfA/Wp1kr2GYcupAo
oTEUe6LAHmnjQUNKgET1VqESLP5gsKnlH9Kqy4gJsiyKzm8GIyoAyyKKMQSfwNlk
21cHyECOVMrCLiKzYBA3NBt3CKFPxDhyh9Pca/PAOuw1g/1/FvWW6W41t/OCQcQG
Kzm1FTg8Ayp5nFHeFtZvU82DB0MQgS1djG3SpIolUMIKTW4DYcbUGWf6+g6ZySsF
0MaPjpdarM9Rr6+V+wnPIP99MttgVtsSr5l+MLhCrcmfGjGhZC0v+3Zwam2D95nx
dHhgCVnVPQE0VjAZSE5JMkcMNzaq2kE701C4KN1E77MZcxYakkiVTGP4Dv1mKtLs
Tp8FpbH9oJfDhRARh98KnJx3IVR4a/B+00jB1u3k/UwfwkKylwjQhVQiQLp4/Udh
pxhAlML+0pbFGnJ2ZAsPCLMKGgFqs2kg7p9Wi8HlP+I0S/hRddpGhSZWn4osDYsF
Uv5NUPOEeB1k1n2DlATgmwBAqt8yTXUvkS9GNAnVsfK17vzQ06cygRdNY/4QKJwO
6NnkyEGL4g2lVeXYDyLbU88UkygLKA5KUMrHST0vyIWFcODBz9oVOoCnwRx85yeF
UWcEWK+hlMujzBf/ysMNqtCxq67H4jVf9UeaUFTo+t9Cnlv7EpWjzwgSa3tjLpsA
NnO/Ie8c0HWXN+7bJ/Np+dFgikpU2vGjaV0oHIpgCG3UpdGKxtCHN58/Iw/vE9Mk
bdJC5H5IVJ6a2JKVGnhhqHJ0VyFjg3VaZINcdo9t465wAKI4cgvXK8Pjs1L0pzFT
mofzBewD3bbbiIpSYhcDcJqVbyUSfZFIDEVoDxgf+HzmYMUPHL7SUZTP4zTmjD5f
Rq2vcomG20d9aEijK2xzVTr12mMBoNPW/ne/haViVIcjiogoAG5il8TlrXbRE/Lb
W5CtZdzK41IxvXkwHlfboV8Glc26xaOhSMzvS2hmBKkO38115ZCP3tZqnyBHl26C
tpXmGCLcgQaGe7b4tm7TElKUPqEx9f3Txktpbc9RWH4sl92/vN9+7W45bMmG/uMS
Ewc6VririXsA+2E2ULfZAmfpxCpKt8CXlsD8u6XONJhkE9piQtD8XFxczsBdC0H3
WPu6NK7vOus9JtpiFUt9yYMXISFWV+UwYkzRAKi1398oteVqTaXodOSTPVEfDbLJ
hZMnTjSFfegQWAcS6KOLWDGavmVJZtYGK0a8Haze+hINn8JP2GD9O78P+4wnNHiA
jmzstnbnzmhqariMNNuvspZhPXDHtQCsUNHr1m8DrldEX8skkFVEot0q/fGgnUEx
2osjh87mGbBrtdLn10Jgd/8HwKM8gVz62Lno+HQL9QqsK8StRHBcNQWLMHxYGwen
72UZQg6w7kfBhjkbP2C4BhqjGidOJH1ho/V/TON886jyY0tovqRUv3bIAKML/uCk
eEdoAn5adwArny4YotPSEDMfwMqqaE4H2d4t5kZAN4qArVuQv+1gP26SDJ/3WKyb
2zTwjKhY5zo7CeAd6s+2IPLiWJUaeoOcTKLjWEtxuorAtv3E0nlWIMV5lBcciaSV
zg2G0dbd2kPGPZmQP3fYL0wjf/XCt0jCdO5FoBfQAJOWnkH3qZDJ+7fVNgwekI9J
WSE1jMu6fBXpm4UyoSui2wX4BJhkZAoknTUC7dTDtIEobGpRnRZc8XfiuAQsyKuu
iAJwbej4XI53TUQgTcRKHCLRvMb5jgHaICN9FOuBSe3vcNluY0YmDXIVwfJTD+JO
bqpl1pC+hs1qrqB2xnA446o6lI5ezWQjNKiINJ5u461rqoQm32OptkK/fFrevLCx
CCIVSXRIh2EJey2iQdvIcvk7NqpHR2PkxGVzhUVHqwV1vTAE/7dggarr/ha2UozA
MKG2t1orCfrPIQd/k3TFCSlwjrUG+9PJqbfEy+pmA0FFBsJbCq9I61IMU80NVR/I
aPM37DC4zRmSsQCVhMaZH/m1e1icnoAH0xLKwzv7K/3nBCo+rnJKm/8x1a+SOFvc
hjyJrDY0NowriMS7EXUf8uwfCLQbvNIMOlNSwMBwj6sTRZvRu09vBRr69m6pAsv4
TnQs/774Bopvhhoi9QSwSaYrWL3pKqO/F37YjBMmSJrnJxYZUz/hiahI0AXkZ8OP
9a7mer1KZFmZ/fndETV9tUdzBimZgSv3ow2cIMFAPfcypdhbfp5lod/pcixStuKA
fpoPNCYNLT4saWU9Y0mhtYvXonKprUKVyRAB2rWtxUt5M/xDR3Yv9YRGkVTCtyb5
tEUXvXDiCwKVoK56Sv/JXFNow53cRbVYyC0tOBGOsgkS44UHv5zzGzdQG/IO0APy
y7eUgsbPfGwUvYgcH0HE8C2hjT82CQtuKAjXGhIhIsuStJ1jwp61vxV0KXsOCJtu
iFOpr2NxWVTLSTnW7fvXPAr9jDin/lnVnCsC2nWfskpZmdwB5nD1lnS4W9SCJ/Pu
sjMvtdnZcYMgkJhO3iEEBvnlECAdl2v6VEg+x3IZYHjJFzmhqsG4wNX5SaeYvcFR
jqAeATjNXAOyk3wOE/YcdwhWcxgjriZdByHAGF/e80h/aq9VJKFFlLKtOX8xtCta
ZQnmKg3sHIEBZt1zh8CCbf5y5XK2auzZk3Ne0gsQVwYTqzDDiQwU0nAcwQiLQxmZ
X/qlyQQKvhR2oaQX9q4R6hbBVCPmNCfQYPWXkxKfnY5xdl6VnQ/0FlrcDkGT8p/U
lFvIJnsF/b/xmV4RtacTXXy48yw64iR9QeJ8Jg9h7bR6mpnwkyI/14UclKsTpSd1
7KYXocVN1IiC3nl2W7gX76NnFpzx+fUtFSb2HUmreFL+Dy6nPCtaE+aFRQgd1ME/
MneKLL2a5Wbgn4f6DZdNM0aw6FjgtP1UGSGCOx20a8hPm1zgSvHe7N+BalrLvLR8
RCmDBkBHYfTGMSPqt7axXsB1Fuezp4f9IWDPcf5QT/+/7RjvHJc28CqBA/RCmIM6
I4HPy1Q51Pjtu81HP7PgDPtrDdsqR4VMdz6O7oaOu+Ct/HDlbiUyOIBcD2JeF+tt
WRF/bsl4rul8fvfvZ6O8BTuYXVlURVh/QQ0tbwiYSC1nOREoUdCH8k858g2fG0lB
cCxaWJVGKWUHapY7vuyQ64R/YxJuPPr8ysY1AhLk/5naRZR5Ge0VnQv5/81rx3PR
k2buc3Nru7/t+tiumtFbCpX2ZQLgJUHjmd67ohT3ThSW7XW5clGA5mclGUp4L5U6
HoRW8S+ger5ULna2eCkjSElxAdER+ZqQRfSLNFCfVY9WLwThVMBta1WZ4unJ1H6s
OFvSHcOxGerxySGL9GDs/7YZmXTsEBC5PD3kXrrD5XZb5QYRP+hpVZX05q/tm9kC
f3+d2M7hUEEBGJybafD191ma25iJ+VGrtnGDabAyeCPYFYRa1B4ZSkyY2VXLJ76Y
16JNhEtfAdnz101ZCy2AcgPZoDgOQoMCmMGXD/TlXWFD4nl3xS/39OV/8PMRqi24
TGP+KL0KP5SifbsWeI8184QXfgXfni9G/sV83OtbBAF2H8VFGc02lW0Y8PAAAnnH
5ouOpXpD+1ftOZEVY+tR1zTYsMoEH6alzrLJ++8p6bW5kwv7skCHN/z8Maz5M+0U
tJeEbxsYhhMsGrSO53/jBaoDOyEMTM3c2dUNqXNrOIzxpuDKIRIuDiSyCT2LsRdD
ef9ktLRTEdKqmg4w59Zev+a8S0gWarMHyZK99ik8R9gIgROp163T6C9pRWuT3xYj
OSYMhAOsbDIrnMrYDSWsBaFBURD5ZSOdq/UgNaUWFsvJxWpaIuD3XDuYC9SnqVf+
Udgx8LHOaLYZcspjv384ZUUW69qVpD4BwUNURcN7dFBUJIJeoBQJD7Gtfuj30WjN
4pkCHjJ2GhhhCbflnSf8BlXs3p9zM7ObE47GmwsIbCtNLU7Y2rueVtjmOCkTBGBw
dB1sQ0t+zkNUdQXAlPQ8cyDLt0LcZO0epkUjcurfPmGHbz46jKHqE1WTbtHATqSN
3YA9I3KO99/aXSufBI1PA2mBEAGbiDSx3pejGyR9nyjLTy7lRPH+SZRdNDE87HdF
lyC0zEDZaEPlswhm8MUOw3DLLsZCT4xVq9RDCPJlzKVHEfjyAoI7XAKzC1hFF67f
1hZl4d7k20mufyOqHTfnqkJQKp7yn/ws66GgjnwAHdjZgL4TEc4DVgx/dfzA22nJ
PrYOculJYG9fW2XQGauwUSicU+gHGc68KUGS6klK7gujzqGdslp79V36jSoRC8QD
YmcRV8CHDCEwD6ShSxf/q2RqlVRcT7KYznNmWEOtJcQEfSvCjEND63WL7K/Ei5sT
BfRmBWLMrv21OaZPfzOPHV34BRzQCoHdzMO6BJUr0ByCZE8tIs6EbB2oIeBrTZVe
b9jJDpZ1bSklQv4y97xPH8uzEPHUd81IQAS0gXIUmzNQR9l9W79HFeAKLIkGdH7U
Zoxu0ve78MCh+jZmF7NXnixGvcc6+YTl5LteMC45LozZi7rDOxVIsR+5kH+6SQao
5bpH5VpWpAYJisLMn6ZqupjhbXuQJ9gVAMgVqk1qj5E7lotJNmlYPqS0gXfy7OwM
2iIB78Ogc6IudJ7fNSWIjJUjhSnV4+SlD4BqmbsMAsnarOQ8rQ6WDdqPreEGD/TX
8bUuP/rEv6Efrh0qFSJO879W+QBmtgTNKbUWdOzmki36kA1gxQ/ZlMLCYOawDPTo
FVEUZj0wYmKpA9NP0T5+KUkSsWnl/s5gC/3N3AlTJbitPBVZlMAWQyYF0ssaQfvO
LAxkGsDI+aUaoFPy36mEnYv3S0rItTPKwCAZIssUhWOHL2eFxcmQ4JgWPKAWcFsK
S7iI9XY9Y3AOxwQui/m0/R/U4/31PVsRks3BQodi8pPEYvwI3McM/Bjsw9aGaPAz
RekLbAfpmaJq+xMppokZn+GyfN3Iowhdmyu9yCiFFOINO9J0f4WmZ42tk90ygXBh
epgWkY+LC2bejL3MMu4nOWUuYM/Dst5wCX1M/pk73IZ+ySNqxYSD3inDCAgljpyz
Erucv3yPw7LxPwm8jJ3w3c+Y+VOLVaD9Eqpx3+1iXGeGIDZMZjmMqgECxiHrn6Y4
Txcu+OF8HIKnwz9eS3t1XntlrsapELILrIjzU/wxJDoTd4UWYKAlz9GNz+CyTh1k
nYMwQNm22TVnpG2WuJ0GI8CoplHp/pZnw5GNMgsaD4Plyl77My/ufb9c4fYqxI9U
OWUIJp1kGpoNOaXxbkc0xnTLKnYIDb//BEQyjPynsttbYceWamKu+ksrW/HU8omj
qoOffxAUtG9nIS9AtzUtLTyXQNhWnMRQY6oQhdOl5u6YsI+eY22h4gfizPxQ6SyK
nUwg9PBO9PuKxKGfR06TBIzbI1TazJpelpsjRsxJ5JnRyAOzJnDGF0sM9RFi5DHW
K9i3foDwz5XUSvSuJM2MeTwD66oTt7w/Z6NucLVgZisXOHOHZmfSnSxdBjdU3Nx4
GD49BgE+vUd6XhUmbYCBABUFkOnijjIcyYtppWujyESzYG4vHPKZVBIhKNDDUJjK
v/wD+P/NPafEffckXTn/J3qhuV3rmvXM0tFXmNJ0LWH+tR/Xd8fYfdFUS+ezZELc
/Gxs0lize0wsKmZF0nvB5Umnttms3wrhg5KX+rXh8/bqWIKoPmiWF8ou26FP+AU/
S4N0n58nww6NILVY3A9OeesLzdrzt3DRydF+O3JhQApSw6TerKvA9Gp0zmBkp3dg
NIXX7cvPzbOarzduCYzsjbCznigDDFpMMYSLUznkLKW/kc3Gm0chznU/Fi0g66ZN
z0dP+v4eM6NoY8+SH9guiF1E0+hPXcOln5F6OgIr/X9W/lgOeeusiPnSp3uZjtMb
bcoTsaoVk9HPYxGqk2O7c9e2DifPe4h/z1MWQDJ7IFFYBq66cXHL00OmfLVKjc5V
FEOswpHdFyOT+XiD6aOxjtEQDP5H/Uwb81tWdTLC2a3X5heCP8aru4COgdvuxKr0
FJ8775AjiEJYo0KkgFBZU1WeGbjVWtEjXYhcr0IJoFfyXTwXw4KhOxb/Sh2drJn/
xouv0daz44bbEQUhRYwkAZiTkIYLEhj6GPc0XPswiOdAoLNlpKjmbhVKoKStJtDd
2X54oEcFTaLHNpDcZucW6wGPjCvsudDzQf9n4TH/gbLR55mV7R7lbE8br2Ph5iwg
Uv6NQN48ddfzmUn2dEhJ4KgLv5S9xs3NVdG+M5H6kxigHiPXKN/nZOWsCE6zIq2j
SDwbz/J6pzbqGRnqPe2g+z/OVuONEIfiMeobfJs0Ks8mbQUc29D7xNs8fh44x3gT
wo8gePMgG92t4Mpeubi5i0wN8z/hacl7zY7mU0ltiYgPfD16IbFBtu5RFjPwoBul
F5GOOpR21MjXRI1RK32Mgf4V/E6OouT9einYaqb7QeyNlhiPyTab4O1KklsaPe6e
4Y89D3esQmk4NLDIzX8vw5bys/WaXdBSZYk46VObYyaLecnzjRHWLFLCs6w12G1I
4d5jfXfNRtuBjVK1ndUhlWhwmR5Ofx+vaDTtDvt9F+ufxxWtmGPxl00RatUYEwYV
Sce7le8jCmD3BY3CqSbdQlG8uYjy+maJn9LrR+VQrh48gBNk6hLzJ5TXlq3MHcCI
jAAQwWtnALsnvsv+DFeyveoVd3pdpqkBIgGt1Tf/e0kyGm2ZnkuuP/kQ6Y+Sef7D
77aBiYv0CGIFtG6xmFs2Y/3r0c9/V/R/Ohh9KIeStS+Ri7V5nZJYgnDAMqfgLTce
C+zUBVvNm9DvJ8MVYi3nl29MWjBEeHTGzxNmYpzpDq+TqPFU0uc3PTFmUmnVEBOL
fZM/LAzFvWlTqNKoqkmMwDJLlFPIWHKTFqM9akEVe0sdGvh0sic8+3lz9NF5T9D+
MwdVK2I0rBARDvlXZMPtcvfyG8LQFIhLf+j0i+9SO05sWKDaWavzKgO7zUjfu4YH
eB/pFf/ap4+Kerj6Xyh+OcMnpyULnv+q/h9ripq1HC8CASp/O+h2fuMiCbBtYGK7
c2pKX5fgk5jpcAeqwbcuuWkLq9JDXhLZxzmQaeGL+79BeRIvcD2cBxnnUsRYeJqs
RQxhRERr19Wzc30Z3vb2tgDdBMWm8OU8uqImrLGOBvexSxXAAeQdeuz6msa7KhHi
g/1+6CLHYJs5WqNFcjRWXfJEH3FxaU4HZj5/ywfxkIm+mme9PYhHGWchEPnt4GE6
zW/59nU0ZIl/uxLJRyN1mOlphBERG7hnOl64ERfgSLvvxDaHfMQZWvuruvLWdNsZ
ndoByzIZucSbHFxO9aAvPz+O0u33zpOuTvFjZc76dI8Aham/Sr0WXGLafykEaWUA
T9WaRS8bGak2FU4nHRtyV4DQEZD6a0v7vS6udy8zTespkrH+pKIY24sDJlvJzitr
Wml3Y++xoYRYTYUXn6UB0JYyCKvdNmD1+WJc1Tf8gVUinP/IOXMBUT5/SIq9wP1O
Ib5Anwbvajo1K4nKxTJVTUEsGTN4s79sfHOzgbihgQimj1a+rRpY6h9EFjZZ/MFO
37k3t7vYELAmZ4FSwEIItxbTI6H53XBQfCzzeMgz/SGcJG+oRVYJ8KS5KvQOz5N1
tfLTKfFzVlinaip18KVpbK8qa/iJEZ5W+s2s1kapZBnBQTIMl9BnZnNnRgakNaEN
L/eJzgFjE6BBbPcwAGCcreK5Hk/q/Vrk4rqVXfbB/UGxUxtPqS0HRB0vP8vpL7Qk
9Zilyue5WS39d9JolNHqKraXNcDJLvfJAQb7H2J6IdGC+7wDq6c08KPbH9QIStgV
PiYyTwapextJNBtj9C81TAeOJVhSn9no2s1aMMibARgizqNM7twjEDcOFpxZVNGn
LVgL+p3lT/huBVUjpUiv6XY8cGl+b61CeMQ+Y1CiVW1RXMJefdavX87jVH8B+cRW
2R8goiaD5Ercb7YnX6z5hmL0vJS5BUoiGs4sSRZZXSK0B0rVQKZIsSa8Pc14hWs6
rCXe2rbEhlb5KwM5WPq5bwBw48vzI/dOnLs3RMS1CCcdGhnk6iR+M6ZnSaWGN1k5
dT05jJhmYT75PJhMpr69Tc8FrHSXWzQlLiU4eStRrK+SUWCrcb4Jf2pNbcD54MXg
TNz4rJLoz5eW9AkyQOcY6JkzShj9Q6MhwHZtFYutVqCfYzD9+JYeaeor32QGF0jb
dtdkW2779DD6DlI9+JcXVmFeMlTnm9z9A51gZO0YZAZ4uSu7WCpJg6Gu1oO3SI47
NFUV8xuTq67UH+dKt560C/lCwCh1AolGPWBEwEaPfQR4AaQadQ+zhQbRNjMdb7pL
VGprJQgH8/dP/06PN97fqySYw4gmdm0w292r68hdSKC4Q1lycIVP1cQ8JelixGqZ
IUlWIJ5owYvsbDs0MXUJxlME48ohFBrbIyje/Cm4mlqr5YXAdC6U8Y5Xdc3bNi5D
8QWgYJ3RmVB8Oevah4yu6g9S0CgE/p0Y5FXfxkogCBGWTPSiMfLq/IKQ/xrORFMW
wg9xY8mOi5BBMUIHX/fNGGsvwUDhWblx3FV80NXOSyOXke3WCW1lUX3moX9fj/XR
KCnKizmloZ/tPryZnzdjQOnpqSpD5MPsY9gzQp0cm/4lBriE0awcpMpR3t+2jHGl
BYQ/f62PfUYQfakNl9/gyqe8SBaLrk0fhnSWPUZVfgMjjUnbJyDGRxVCisDxekMO
I+IkdQunbY4ogZurG2a0SsjtdAREwI6mBt4uhLF+lSf+F9/G9eGMp1uuPeNiKNyg
aFS68TCLytp471GbYr0vE3XIDFqs4P3aITwXO4BnB6PDfy2umsAl79N2X9DWQr+o
WuVdb7SS70GQH83DtW2mEYjJ+X81jkS8r/SoqAzpI2HeqMT/5jRdzs8tdwltTOdx
i4K+vdAa1LVmb9iuevs6qgECVJ3G+go0+3xt4H3JcPipYCf6OeSKsPi6Sg4jqgsH
Z7BLI2uAWr/FDmZoYbpeo80uKCWQBFiNtL3LwE4WnoWGfKKd1zrIw6tiOn3bPi6e
UW64uYkOqZSUAbd9XYQkHPqvE/Jq4qtxo/WEbPA5q54bUDUGHf95IIJyuTubFFhT
BVoY28IzXRdAu/vNonHp5mUfPVpfw8PsGoBnqX00KKEPVj3ig4VCAurMsLlD/nuJ
92FuoHHmDs+2Hv7vzXPVZ2MkFqRuM6sWMklRmX997GNfVAq5pOm5pnnHFBZxnUMm
StH3ouy8UXEJE7Rdl2norWG3qPoYK4pSvxqINJzaCIc8c/PP2pGiYnDZB0qkDJUa
M3zKsHgfWHk9Ne1BJ6aDBoCNGxH1CSz5jUNtSGZXuvim/hEIIZIGHKD+tAHQNuAQ
wrnxdwMe5rui5oOA1YGRak/dYBbta1atxOSR/LUArecHnXYn/aYhvaVgzrqg5Ez9
bvfUdnh2U5x/Ous0pi07Cb4sRrX2Fwk8iPBdFjSvhXzgGJlu/0clA5i5Qu21EoQh
Lj5yqZjeyuCZP3x6U6mvybAj6OPsj4RP5Qq1/1EPizWgEO0jUxMa5ODbGRKnn1MY
xbP5HSpr2oEukuO1NOEaLoxvOM0wrZ4kHx4gULZaABLMl/PfBxWq3SFE92f8SLBO
NfOoo8Hvj7iDjbDwvhzs6j7d1oToLqnMMd2Iwj9xokibkBEc4GM1xS9QDr/jAhNb
Lh9RoqY6pL4Wveyz2WpUomJYGDBoX382biQ48U8tiu0D2WkraZgOSnzAS04OvYyo
c5QBRVoffAb16EPvfUjhSEvsmeLOJTgo0kBCmOeiHx3n3RWgd2U5p1CGpCkuOcfD
szjiTfdTSKyqnp67tyixXYgLAs5A0wHuu+4W6qvVB09XchsQNY62Q11K3RDy5zsz
bP03bMXF111HsQUZb551g3Tp4V3iMnAXozPB4KpQBfnG6pGWLKi4az7e3G9lNKsI
7q6x+qXpta9eBT74n8CFu4/sYu53LNfaSAo4nsVh+Pw+D2KXkM4KXL/9p0QOFM6v
OcHjYwQpDA+N5yMpzYWUvDDr4OoEwzubpcqWF2syAFAJljTIMB8d8NcN2CJf7vzk
FX/yKnpQOGs9meQTsGXCYy2u4wcmGv3UkMzBFSoITlA5a8ZyxNULof/OS2U0ODLl
AllMJahQS2e4yO3HnvS0eQVFfm2hGbHiJ4bh7NSW61JQZP0/51YYpZY1IZxvFfMz
pNmmyBegrqQiiEkVsPYp8ozpVls3Gu7SJdXXFBK3E0piBVg0G8Fozr107smvLM33
kBqq8khFyR7ocyamBCNdRhq9CxqBQEb1PrKvY3jsc7JoYzeXhZu0g0UZRidvuZca
zoeyjVIoG1XEXjFdRVLNMTxQrdjP+p7qG0cVnUdfeU6S93moL6kT0l6xIR4w8SNJ
KHf5KonFk3WRCoTvZnbnGHZ64smbNRP/7cxSNNLWvtTQhjdj0kuI3W8G3SjoXa9s
CJcnUtVUZqFmTESeUwp7ZyEXfoPLbd7ScKW22Sru+/OdrEKkgKJAmyEct3c8yZSy
7wvXPgbBmidTDZKooAMaLfVQDl9B3aKK+aC6pYcJ3RnJHLeJOMASUovXjhyMyPWe
haFSW/5uFYZSkHbw06aapJlRG01a/tNjNPExcWUrYmpfliHW1b7pbfEt2f8L3INg
rCPiMWBtRGeutjSmil8/B8xT7zJBtYm+WAnzyMIXWViqUSP1e5cXRUXfJmzhDAyD
WwDmQfm5QWhu/nam+OphzfrZ9Pioijg/5mB9eye15Hzzfu4ODy3sObRNTxa9nP3E
S691dqEaKK30luEvFFtVrJdU9bfUkQUvwcqJEtmf47YBAg8WSW1JPiFj8r2v9onc
xZYrBreTdXStNtHDSzlwl8UqXhLuTiHjDh7VDyy54xP2hcVSD9N8NyYU89OSrfjm
RqS7sefZXsVm/iZCi0JySC5goZYbJ5+57Lbo0zyPembff7XmaPsLl47ZVg0EVcmC
ww1B0fWw/O+S6OJl1m51BWlWnHOx1+6b5Gl6wVvp6+2cr8VPME8/Jipd1rwNE66j
RrFGCRtiOpWa3jLz4NhjoYHf1+g7fi06GgqzC5crxwO/YF6GNjXuoiQEYsc9OO4N
vT/UMseNMrhUMqmw+vmxH7iasUhhZvYThKWOSS69qvLm3x/DA8rllDRK1Y/nquMr
+b2rgbiomhwHFdtgANBTFuyHspXZnaENu32whrlTRyrukyKNQEYwGTNl2oHMtO3a
WRazXwFDkmm66W0+gLMtf4sIOqIjDOU+ne+21F5sPmGwpawlmeA3Fk+TmbzE3See
uTaHm1rEYmqaNOytvfLzynxOxbQthjYxr1sAhw1VPwY+YkgZjv2AT9HoNMt78U6d
ro7RSqXz1S10LqqmSG223gDhGUAj56QqEVMWDQkaSKtWXK2nhj51MtIWFmragGRC
CQwP0LzOrx5cMsTf/I4879ASneLvem6Y38rE2g7OCA80H0ki4UMdvth+8XSE7N7r
uxFDKWr/Ug+2EezwAd/gR/nrFjt3dIxlpPWXULxLUdvNQEBRV27dOpbfR//C+JkV
Rg8/u4UnLQSqVOmD9fSWAX0h+284EI1LKN5FK0WaqjCHr+2WK8eHOrtZy+pV6ITv
x4PPOL93FQbDi+mZr6m/DVABWapjexlXK7+2VJSuf3/lboGvbQC7WxcPyI2rbqez
WgEvXk0YWrBO0CojnfyCYhYRdw15DCGEHBmVNYDl0h2DEBjbZvO7Tav6Zbkxeffo
qXy/eoT4IREAdwAGLlqlgYdKErSnuu6EtGa2wbRWwi/J5boHf9FDkI8/OiDnd4O+
qGMA1OG+Dsm3k4XMJjXqcgLKBAOcWmcG4GojFxY/KxHbBJgboJjCeuPlAsD/GfkR
ZgsqcMhkBiuMO+Q0Z5zabs/tF7vAKYJ1EeAnNZF3I1q/Iu9pCQFzmal71rQPfZS6
b4iwFIaJoHwWWZ3QbOgMsXCY1aNy5NnbUU1EKEXqxXx1DeUKWvhinxjHewF9f0GO
Io4B3aD+Ar5SIjsBrNYgCIa3ea+N/v0gnVaiZlYGRM7a6JUof4/NKXgwV7IGiDZS
eC3KreBkM/886cRZvsHdlZwKdVDJ/LPMHPVFtKT/hxaIRT6ioACZcspBpMUsnMAU
JEFHf02jfaoSL7SDBXWmYYeEspspykzTMn/MpAkbx6RlVWpPJiu7lqupUtkm7m6/
f/eUgEEswjxEPWJ/TxT6uh30aG+GTELdaRvWiEJRgwRDaisjzQFAwt0hWFzNX22o
YkVM6EfESqo5m6O3gbdx3wpPojQZU+D3+Hlo63yB2wzaiujnvUYa+20c8x5sx3To
HXAAT/lTmrkZuRKOdjttbV8O0JdISE6jaXj4mFUB13KKyKsjBXrNiFQsmbmsyqix
r9EgN3eFXulwCornpogp7b75ijOXKbk8ooB7bVlyuWOwY/YKBq68aN8iHKpisopU
+Fmrt+T3JN0D30eMlnhBFuTjR2TgbAAS+mXQpTfAA8uyhGFzl2FQg8HWspsGVaZl
UhJLT1+ksoGAxxFhgHpbM0h1bJqKwhXPxFVFDGdgAHTcAffruHOtZo2GDFofeigo
y+kvhOjkJrL9a9eCezW+lRCFNDogCQqg/DggaDEVn5qSRjGe+J4xV91Dy5dvDhO2
te2xNIz4bbsd0313ouOLuKQF6S6bk1sVr1KMNaL3fYbet57vdSmhdcOVXYE17o2K
79QyQkj5wB6DmTTQ1kUaRhpWxUu+p7xErswWb47uz5FAxEOxba4fwom4JD7ErhDV
2m1PbjJlFHAIM+DGHc9xacTy/digg8rQFWLQsLXsCm1F1P9uZdv1EqI5RwooqK12
CalKNTpENKiYKF/HEouu3PMuvWlhV+0cZ7NDeioR6mMdGL1FboUBwY+c4u+x7g6X
sfw7Hjip4naEDaHHGR7GUBShS06pB1Ikq+DkUTjK3yhcHpqqxZNyuHE1DE+auie9
3JaswzT5ePpoPn8qmuyGnCaET1fIDItAtxKb5ElWyrtV9mw1xvLAEAPUfW1zhw/p
YPdmJ3mzAYa8XCADoXHPQsOlWTSs/z4SsFTva7hmdeuisLnEeC6EskIlmCng0Doq
KnCWk8tARdxSDfBcTEpqbAoPCMKHSuSnhtMZHjHQJ3X3aGYOQd2tdiv5m9wylfQD
nbwODLPZ8/Eh+J1puRmStB5qgN8ohpo+TJsvTItyd0LyNUlA+zr29AKJnbKRraTZ
jYOn4zcYrYSkj524dh4hFoqsk3SGzZafowiCzE74IRMr6JjYD6FXCmPYC/G/qhAB
4514yuoGEM7oenwYNe/aiLS+jh1jahIMOtvf3heBbRXBSwCr6h/BtWnfki5hZtsB
ylOL0CfivxPvLcPCUBeskUJhhon8wcQHV9nnb3qPkt1Irlg40E/iZ4sFikAutj5J
c+qy8qmWcG6kYh2dsCZHkG45ssFMcRv/0hgI71bBPvTcE9aLk274Na4rZb/SCR/C
D/2otmJO5F7YnPP2LJikyYRiY+B1JylpeW6wJb/1JALIH7YlXqya50uUFdUo4il1
VWHR/IDCPVqKGSSBWNFPWmD0dI/fLc1b/JG3/bTbp/tHSznnRPoM4SSosg55A5i/
P61t3dJcY1RD8310XQjvRBKlN0YQ0j2jo1yHIHl0mBqAsOVMEYx8Kl0s+cJgyACg
ciZHK8aY73t4EkFZea8185+td3J4Rx07lyo39KeuTKr6mQf0+1bTdU9uONR+3jbV
PX8ee/yDJbjUAt4sXWQNUf/52MXmO2amF7TWBfmaSp4LWKcWYHuGTo5jujccLKmt
YotkRNvEcfP7BP5L4qThOjF/R7pVR7fgt7R08+JceYPaaoxj1eh/pEvbsGcU03Bg
tcYQrl7LgKJmdq2Wdv16RuNFLvFPI7Dij38Hz6Ohb/NGKhmTFUzr9Q6w+tbAs9Ad
ANpAm76y+vttuTAUB6CIL5lxdCnRowMrTzcaS75yaf5HW93zXohghJW36JMqi+0y
2MbgwvqCUetPrPyf0fXCCJdo15nwjbK1jc7IKTC5RLqDJLKNXZstJcznDVVaaKqH
q2P6w1QnglJcTKzUk7d9rUyEAU34isFv3pD8mcZHoHHj6NpfLmJCBwMo/izCGpuX
ufoJnEwLrHeEW2tosze7EfKG1G6vGBM/qZXD8v91L3bV4JiQE9k4b/CiV0uAlCe9
KZttjZgdBz2r6HRilQBtnjrYlgb6xHP6YDzhT67WY74y4j4DQ16KwK4e7tyjzkcK
F7gvQMERsBIT5dy/mnXuyC3Whpo7NgXhjSAv8Ela7cs6Pd4sX8Tk2Y7BsWl4d1tb
119+OcRbNAhC2CU7zHPnrVmA4tTpRvWjXc2USHZIuy7lWAl4W7qbWwVXT37/m5JH
EzKJuemU/S/K37R2l1pVejh8eHXpnXa4O6piiOzExPHo7xa1/ZM1XlJj3olnLWhu
YCJ66yuiI0vfED7JBFwpr+69XmjBVXggy1n7vD4EeIoImT95ZH6E4KardK+pD3UZ
+/hu1kiL+keTDMw6DCqGcKoa+tYX8//7CFHjN6+Ek6OWPalpDGqHTTj86N69fMUe
XvBnfKzY1OW+KbPB7oEzZp/YSme2d9JKUUwx/iFexlVrPR+zQHlozxUIQKGA+XTP
F7/wal6Y3WoVWVzd++DCfr6eS+WkE7LLQpEH7LLckb2avFIHFz/D6b1HEd1un6LM
8zeF2CQZUYAyzWLx44S4TkDdy87Q8uCHLMMHjom4Rpa5mm/Okv/NfmDV2GmVg3PS
tXTKH0HFE0IhD2JuFI6Cow8pxZPT0za/zEOCipffXC9WOv8UYVQNPwQE6064OEMT
qHunhlH74xflfDHXdtX+lQgV0aKZes1TmryAw+11KRTrAtJw9PiQM/uxhMYwq313
XX7tK48uzvO3YRr282RId+l4cSgcq4ZaDjws2rGA5Q8ltn2+egZPEDrok73GHel/
cKo+lV9jR/94WGSovbcQf8p9xHdOrY01+arxvE8R1Bz2d9nEYRb1dlqub55a6mGK
OvcVaSsCzK5D0jt9N3bBXb+wRWE4iyWa7Fsj1fZKMJAuk6iTalLCjwEWezg26an0
AMxo/o3NRzUyidWEiWPNjj36WHeG7nPbdkvIUARf44bbYJPbjTcG+6BXJm24UjZp
GuXDtx+qVy5lDrJZtWvp6MPI4e+A9rdI9uytPybDSArKyXFynxoQgOKPqwjPAoNT
gi+ALFjz31CZPKhmS8LnpPQvD8xeNkcqT416Q7ePSVcpjKwvjhRxWNSf2cEpPkpf
+uPAeRaTCX18PxZX84XWjpqtI6KbskV5oqJ3YylgjbypPnQnBg8hVzXqK2Fbb9B9
Yb1oiWd1l2+7Q1/Ix+vRFZu1aRoyGX+2WC7cgOF063fO/s7t+irIbKTdjv0mXaBu
XMe1rfnk6+IXaFYRO6Kji8QV8SyC8rhAypAmX5H1IScl+DzKfzBUocTBPehhUYl0
QkUe4YoyyIUZzXDvm8XgV6tjx4ZpKs/cCOxObYEAY8YU0TVrsH3ri1fhrvfGlMyd
8KOkp1cPE0jHPCaHTjWzhNKoD8eY1As8OmpcfdCOm9xb+XkhlK9aetsezfGpaHMh
seTUfq7LHtH84aQ5zCIUuSBS0XdC/4i7eQTqiHTpaC/zAAyL/mVy8YbIAOEylexQ
OmkqIdczMXG8CXH82ZMVwam8JeOL1LLqrYy3LvLdHZYpiSZye+2apqZtudl1o37d
pSG6aW0X3Aud+tsR0FmFTVQs/TFffyfXNFxA04wEcw2LCGWMQeDVVv9MlV8Rx02f
f8gkSETr7aNl0Ibxl4KhTUS2FINn71XzdDpemb3FRUlRnvi2t1i4iyMIDC92c8lX
p0soWICTRNQuclIPE0ItZOc5clNVoRQboUcSqv+e4s2elv0w4ZxHiF4qTh0tGJA6
lYQrGe7k9ljM6MPVjhTe1CxSLryp26kuoAJH5ES/Sw09Rtt7g9zNiQOuePFGfGeu
rjTy0W+XgzSOQI9qhndP2usgTtzLHZZhwSq+7FCdPKvC8k6tMK1BQcHFZGNlHQnk
XYy+aunsvlX0FK8dEoOOt6oG4MuHwjCE6Mc9bj9fjCIeZD3LJj/tAB3LeE5lRLUB
fFXnHz5130pCAoD6nAPoX8vYu4dGLUYtbcPnMwb5lyAcq7vFClUfHt7RfsxB/x9Y
ttCnzCklW/GIkYSWo0dnyYfvAoI0UxAAvH3w7hPDhiXA+gMvVck5nldaYyanvlR7
dBjBdzgS2s3r87sxHVw02+4kllBkdZ1QbhQzLsFpNTF0A7D57xrTvoSXgdKOeb4R
+jK/DFIPK+pOnqox+i2SzNtIjrQPrFf5XdEdINLQ6gHzxkPvG0MJAi9CcN9UBtx9
HpC1Hntc56oC9viHgBTHri+pc7R+q3B+c7ociej43llETiaKKRC3wjwiSw9dD04N
bHiK9O8VXaB84Q4T0GdBNzlpa6YM3t7eX8VHlGGcWrCcD2pfLQM+BIyyLOP1itXi
Ybh27Cn+exeH8Sn0VMWQDzuknCfen88QOUdq5HmrlhpvpAxKsqN0t2LpBOvpP9Mn
5K0SG5glsTOSxMQ7cQx3+Kka9CJJf4RSHPxi3tsP25209yA/kucPZKOS3jzhVqkJ
tMnlql9P5I1Pnq+QUfjSN2b9WMQdwovnSo5hEJgR5q44sA20OxzhbxdnAcg00rio
lZQxHxjKBIbuY/XWLyI4i55D7tRoJw3gHenHQ5fe/Wa6USQGT/NX7gquJ3nem545
12ZNqfewdSy1jC/hNdaZwOChAYRK03w7YIoN3GPj7UnHVRSMQ8ln0Wu6BnXmxbAE
IVowmIyfJ7SWDq46Izdt8pvq8YrHlRlTI11LimhRRocwX4Ow4rzmxKwAHAI7Qnav
3aWFp15yaMPMvDInPHpXG7MXVh/UFPkYDWME5TMYaFJcJH8n8lsGzRoUP6V+CbL7
Fj7o2TWjEujzav5wNyukrkz7irHDH++tyb1hlFLj+uPfpU3SYK98OjSFRosFJddr
JzIEacD7DFJ1vHO2XoyvmZTjfXusWc+0FePYxK6IX9hX+cqn2sYKRQdEII6VjpG+
C9aFgByCKe4lRUmTqGJNAv/5aN6yA1dqn0pv8NYMwcq1MQP0cEPmRrIb289CNy1S
yn7nSNJtSXSgiY/G2Eq6BjIVRNUdYHZcFQNOoi0xUoPcgL+A0bXkxb9q+TKQSzVL
1qJkvU86h+7W+ewUYAXvwETFrguVXfylHDlZhmP4nWI6lBid4jm7JYE1LnAXHwXj
LHOtnyBZDxW+glgQZ9Ixqo5vt8uoSC1EIp7hn1ONbWRh8AoaA6UGyCeCJCM3aIZN
oNI4JMgpGsuc1i09izZw5/r9qF/9RuwMtggk66pJzDB05n9jVLNee9y8QWBlUfJ3
sODPp6XYaHuDCUn41CNdW9hyhT3Mm9N1/nt0VpcZNaFj8IbaYSVtAgz8RtBM8lJ6
C82fzlnWs7vJ4YGlKlmmH1FbrWY5+6XMbNvtpL7N14pAC2gCkMdgBXFnG8JmP85g
xvSoS9WXIsRK+DQJa09ZpmFov/JzOsDqxkivffgg4g2UKOe8bwyOm04BoeOT0Ub6
+kaMAsckxyvAl4sDM/rhnh1VYywXHWWeXR7eZ36O7ol8nHBPLVX8Oj3FnrO7mw8u
uFwiZ0B5T7YpCwOQVDZjPd9GBM+F1NnZAu7rZCNMeKRgKTWiy91tPoxsrJE4pjv2
DjwlsqCgcFxFRo/ssVcZRZOF2D0pOXWNk2XWVcasZN0PpCaG3+GetrMn3/rmGO5L
QUj6sDP3uzr+toSIGnxI6N0WhLqJfwHQ8nDHbL55EzevD4XI0PS+1UpseaB04pPd
OQ+QpWoeu4MmzQBkySymtg7PjQcch1o/upWrixZZVrKw6f52l4XhXDQPlpr2OONQ
9/C+qS1bEcR9JeUQM83JjtZHvuyEerkqrrjYUAoewJrjh2chRVBRCSdyCjlQ7Ii/
2X07+apO/2o0BoX0/3jGXWyj8sEU5B8+s2fjeFdVPv+6ZynAK0r02yBeCYrIS2bv
NTljlXT09NBAEG4NpAtjHHSRxOClId53yopk1ilaPSlJHi4DLIH2RT4BdGHpLgJb
rWjB7S9uYmMvHtfXkGLC5c5/7bk8tNxND27m1tFdgI7OmmBYuAyEDfHUS/x6AXn7
pD1F2HtUGG0Y3Miwkvf7kPQqUzJ/LpY9YY0lFeFuSioRuc0LoUjwPCVOnQeK0Z0t
amxUI+/5snZzpD/gLxl+MMiZAX4sZIp+0ZpgApzkh2kYHJWzuybx1zOcTeZQ41TK
DD6a5/nf7DPEVy2/riCfIfO+A8h4tUSB5sQaVxejeQWXip3JViSdh1YupqVcj++N
s4v5Y/P+bWCr/iUrkGNQ/ImaghP5uuu4e+cvJReA3JLSV2C1JMRFbzUVGswhcEuv
ckQREV5IuaJtnWrEVP19Q0qf8DifZDOKBQ5Vzyt+CXW0giskVqw4XI6AqHSUrNDE
Sn/oWX08+OdwGQniILGox6xl9uIy/4qRaMY7hKJB789WJu8f52WitGNYEfAVbyR4
fnvnDXpZ35jjxKgYct+ZvSAwn8HOYbCuzBEXK6EzWE+gcGiDPOWD1QVTPtZ7U8If
ERY7yu4OBR5+Jo4Rg4Gke2JQTFx+0mWWWpw59SUtOsT9csbwSAfQ3LkNtNRS6KEy
BdW9jzJ63vpr9S8nxBIQrhcTgAqxKmgxGtLJuqpIdLZmZhm3ep092Bk1QDzJIfaN
erKaDWGhn9luY2xqHAeHxI2bbDSuI8nNqS5FVV7D+MxcCizOf4S9WSJaX76C0bLG
721j4z/5RJA/0dcgVIga5tz+KVUmcVFi+85IRIREwyFyU4NEaIDzJ3V3hVAj8LIY
NwQB9kQzZsayIdPenz+e9YvgHzmWahD+KdLNK+eInGWVUYKH/UwXgrbc/WffkFAN
Qq4qHdVQCexWK8ZObx41LFZhRCNL7ONBu3pyx8do98NG6tAU8t7XcB3o9kBKpdBL
IXN7khPvX8qzQX1hdjah8oYGEed0kN0J7f/sIJQHOhZKKGMWhIwpxMUTvc2DyWaN
Qk700UzPZoZj9xyxSNekN/zk+I252PwstXRiLt/N5ok8NggTR0SEGLLHtXcOx6vI
fqZh/5UdguSOSdwhD8x35GpN/mhvEsxlvAoD/Xhed2GEeCmMXfTBmqA7OUNyY5sm
QWPImz+5lTBcZ2r43pIYDeWu9iXfINrA+INuwrnQu4pulOag1HU9hVoX4Q8NS+A/
1HM7E3Gq0QEzFnlg8R/gZ/xh6N0KLOX8v5GMux/Vis7s/QXVOEvdu85mb4SWvG9S
HU79ADJzXJWDD/VCVdt1D/C2mgnaebGRCVYTbfcFg2x5QUfmxugrfIt0w+UGqTkQ
/yur4t847p42PijhnTkkaKDU3Ni2f7wbqMjQ9lJV8Njme77YcCODQPI1idqndzyy
r4TnAcGpdsGo4aj1XKUOG5zZxRUIRPusUrV/JV7gE7ytx6xXNEME/RjgprcKMBgS
cm/YG/+CTzWV8bImdu2sjveja/96xPOOLfeLhRzsGYB9dCJ2Ga9VOZvs4rpl6dkx
phpQDcRyFGIrJJUPC9LSmGt9s3dLCFvnV/k1ICD/GvkwNk2y9sAylwRg6e/dGOO0
eyhLTvTWybct4CKPv1eUct8fZ4FUdRi6CPNE4dMU3R0iujzlVNTPdwLI83Y1TttU
UYmKEbyD0W67M354N2qGBOjG7UpicJPIPtZdNddK+nBB9LwQapzXh9TmDSCyrz9I
zGhP+gStfo8VnMaaclUJmTCO71olLcEmFPuVuHubzYYZjJz7eWXUYMG0Z7wiQdXF
W5y7HABrEZdzL9Rxl5Ze6gKYhYqNbgbq7S2DmM6NKY5mO0A+4CLTMUKWpaCo3W0H
VzbYic83bpf5r5wbTmLhSMyBebLtGvts/zuNqZ5wQYnTH0DH5LNYbZTNtQxffA7X
tfRU4NzzNCoSxuCFEk79TQQxzbIgJpjh6Yr3IWvIv40A3lGf1iJKsoXk9wMTqy8b
XwLny/VO1jUmeLw5wvwZXqwLSypFFYomIH2p7hdsmaOB0+4zgnsaW7H/k+LbN8DT
b4wnt/6SeGlVfbh5sib/kU6jZUQxWDi0DswFUVE9ZZoBHU5Bc9/Z5VofqhX3R2kd
1Qpud9erxzAU/1hBAjGg87BtZmhSieY+u0w+YQUZPXR8vD+ducVwoWu2DqHP3Dk5
3X/rUtU5Vecy8HWxlXZFmd3Iv5A+AeYq0PmLsbuvtiaWkEaIBLSkbqIMKfdslhDe
SKpfhA8+Mxqner3yMpfoe8P6aH9Xk8bGOhlkzZje1KagnA/AUnrt2ueSk3DIucWe
6l+eeQenupz+RuOgJlgGSDR1f8DKWVPJlXxvc6X6u/BcrlghT7fI18OwwSG5Pgiz
zneNHP3Myvtj5fFfkC5NphAD/osCm9d12YkFd17TynKapNseDdeOAOUJjPMZmSIR
JHnW0QaRPInyFXNOm0Zb08UfWnG9cdoSxmXrGFVxvTeTiLv8GKANJeu3mUCzx7oM
N62m0vjuvxbU3jlv+TZq0YQfGTTni8F8Bf+wr2ta1d6u5gtrkRCgWtBZ6o9DyKfN
WOhLeXXX+E1jTp4SgFlof0UY9uRfRennNgnE1Enhh1r/bioDW8ANu0cyVMj1MDJj
SvW+TJja8CRACHeFQbSamBZiM9/K2ZuT04fMQt6OsTZUnmLyUs9pnfKfkEO0MKQ6
9SqwJLOhPr5+fOB+EbN7aZRmqlly4whPbST6TC9xipCVd2Fi/DRyYU3+wRG5lXqQ
X1K/G1+LaheuOXtk3Q7EwFh4zsRRKR0gYfNy3FK0ttrC5LGkLcF7fi7LepX4BSYd
cy/Ae+hgHX/UC5qqkZXodf9Ahjxpt1NZYzR9zIg8iQCDGkGq9rjjXenaJ2ptLk3x
p2iR8xK+FStn2CRjUJKu8I2wrhY4isPlbK78sciuRvUaWDEs3XADhoekQj7L/+d0
G7mzd2nI+fFo8LrH91rHgVfQmeIMDhBpRD234ElH+7fwHmrnpPJzZLiJ527tBoHd
XosiWF6Cdb4ofTfSy6/gsoVzJz/zu0gDcfro//u71twNke48t4Oi7tZvLt/DY5RR
ITebicxeApXg8dZoALk/0DAX+Y7NRdnniYUUdt3XcwxNgvYxn0k/NCM/p+42pquo
129cR3xlsn4jnto3jRxGFf0bRrPmtYd4Z9lJVfJc1o+JPmUecL+YRJ95nHXICpFz
4lZZThb5gnKjYcLVt4MY7Ln68/yf6M1tiiR/q9x4Kp1dv14NPf+mdZ3Dm5C9uM8s
rpuPl5lbkIMPRpHadb5q4Mm+W58tjTOS2PFEoJNQtG4vpaslvW/3+voZYTgOe1lz
LuFyEMyiRoA0fw2B0SNGF+fG6wfDwkL5mGLYGeC09p7OOGuywnmHTMmYeN9t+lu+
TWOfVriAfjnqEpNmk1Fp0+WUrgGuCRuEVmxQiYVgXW73Eb6Kx9fU5Mw+oto8cyV5
BbEyrAs/KADuqEygPmwpaQxtrn5Z4HNYUUrHeUGrKMO7AtnDYT1Ir0dEIUxUMh7D
I1RCGKhi02U/Zm1juVQU6RVhz1uTCEM0regDAE+Ux/Rz4VNSBLx1qytrSXeghdFb
AW1mwrTXl8d8Py+OprpXBduvvXo8dyJ17Yeq+ayw2/jJvKgrc9YmuPT+2WjSwDjY
OmcWBuTNzeO98FkOM0V6yxAyXBYipqh/G8gkX1/mbUBln+1A1MlCM9Go571JWgY8
4ld0vqeYW5NZ+APgp7vI2Az+MAxFNCL2PwaGO0saW60YfjMht7D0yCiYvvb39QOv
Iyol8qHdr2AoJpMy4cHCxShb6C61QA3M1lQu8Nh5EZAx1gndR8rGboVrsIM/c7ZR
c+XnGJ1ZNInaAFy3/FMvhArrv7g2Mt+9Vr4jsJrdXzc9/+0GjjnXPEeefR6fL3BB
s4ce27nirh7s6Aov3gHuwWXHzcUqjqIGDSiFVOYtCeGF3qfcv9lt1VNz/bTa+NFN
w09HS/YVH0zsND+Nyc2U2Y2Hv3lmxxxk6nzkEdRqkLR7JUcDCn1yFZvAAy2HLcZB
HMuwg/KA3bhe8rnDdn8Da+vdRwDRRAsimmC7thgl0iZnocnVrhYZRzvgpyxECQmU
GVtWeuz8z8cAfTlNHi85Zm14R+MhEFVfTy3diPiQvwpEEIN3qW0rNyUEnl4B80Em
N4ZI7HW7Jv7cVL6NtDzJtRgTvMZy+N7xPQJy1NuSoUxOu5KmCJZV15E6hoIfunaI
8g1O18tZZbf/gqgyJCSp1Yo3saPyY+zgtTy90gD7MfeRWCC2Bz0UCI+0/KuHFaqa
aai9kOYgWJjJBqmGdLwzIsj13oqrc+hqYiqXtB/euuxflGtU2sammCPyrrZAJua0
ATEne9U37wNd27XQKR+LL05GdeROHVq477r0XQR2GWAcG1GHDMNxjx+bAoY27vHR
Qbw18UJjzgDcf7JfdH1SrktUnZpnvHQrDnDsi2s/xhyZELwUWOLx2XwRUCGskSst
6nRloF1irjY5sdoZvxnjrTjw37OtreyawsvyvWSLp1gC0mCKctuA+DLm9XN5o6gK
ALnLDxEffxkzzAETIxn4wSNvvkruGWs68ceHW4kI/WVwhSgYyvKH2jpSztBZE7vt
vs7XtQ3mBpzUHxavkIlE6CtMZxN06zIsggGqKZSkXK7uJ2McyvV6HIDY+zaC2Z7t
wqH+sn5y87ekNSxEjvi44gMBnIXty36SZ/yW+fMfpqsuOLlbHR5lqrtia8Svb+Kd
caxRkjIfhMqe9sJVltgPa2rDSMo3wPjKDqXaT5SE0/vRct/BU3dz9XsT5MUovpz3
9SrFRJl5YpcuQvEeLCDBMTHLb+rdo1tYFU31lo0dyq7rw8MVwjZyyFoWVimFX819
ql/NiFXaAt9e9kC4oGr2Qs2P0gmGVjUbJ7rKl0iEbA+16Ny5f1TChTTUz319ncJ3
Y82aOtWhK1R69qeMQDnNOzApGoJazmXFuH43K2C68O4Bakc47oaeqhS3fwGwjRSe
r8TdP2ytewyNWQHLpnNTig4gTOZjr9jEPLP3CbBQsdYQfQUQuOBTpJDuBCllcJH9
ooSKeQEqW1WbRvjnY0M5zZuohqHeXtRRv3cWB7WGVI3VTlxgrDD+7024Jz00bQZu
sLARSDR13Zka5cKn4CdWmuenheTRpb9KAPirvwt7Igbf+FI6Rg2jJka6hv6Ko144
nw9tL0y7iOcgTdZ87r+8PjmwEixZEleKeGP963b3jtgkzD77f3LTzmUlGTSQMlJ0
9EhkDPDQ6l0qWDK2wfsJUpNUOjy/qVMzl5GbdZGMcxFfH7iM9K6mzASX0FRcUsGu
4s0uz4O/xNIyiDK2nLyIEf/9NajNf+QVitG8wuoIsxbHfMFN2S0mRY/u87OfQaaD
kvEHB8Y67e8rOzpgpptxsL9jk1YRbUFFhoHZIzN2XBehqifP27osFEKQiSJf/873
4s3F78jAP3Cp7h6TuYrmhi6lxsiFij/RHUjOj/YDBzW2kiMUFienww1hPQe3Xewc
5Pa2RAElsrhouWd8P0/3XSrOvML1YqDZwAib8CjFvsHB+tBdlpMtlaXPqBmbH6y5
JEg0zM3dktoVadYnxOimjSPBIw2tQjwGRNIHMyfj+gn7nAzelLMdLwaGZSdFmTWD
9JvRYD/wBGzJOdqtWgrSGsGabfn5oQzP4y7faqP7NkVlsLCm9TRc7Qejk0JKoX3o
fp1Z890s6UuCQSWUu+9cjK8N8fsyCTVYi9PX8kCkYUGLZGje80PnBFQVTwjjeutL
zaH79AhBi/FQsQ0c7Vny9uKSIgnYhsABgHqTb7BBMoOU+FUWj3k2q51Vks7lhSM4
byb5g+o2XULwSJ6ryNkkvOkmdLX7whMja/R3QG8JpsozbXXFBs47zzyi+JspS+Zw
CemaGAzHIZYETzVHAhNk85V0ImPG8D+9wz880kZvEn+v/1tWKpGEb8F9uhNtfGOX
zPiYUqWkYKpMCajyh1gvmhtJNtleGTikPXM0131qIHAtwhSr13CggM2Ku5ETbVFS
pu8diRJheAQIFKWsIypsG42K2T89ReQqcKX5DudkgoBHfasoGLoP0g5L+A9TzS/s
bZE7S6mA+Q8Rcx1xvzxRavj9SjUuNtKOhpp5mdBONQRNfLtiSJor+QWIxzYh7IeP
4zfK8I1Q9MVtwzqBhmT3aSR4yV1xLrGzjyXNpiqaUHd3WmL+22GoqaRMeBtRrNcl
rYS6ZU4C0Y8hTkqZpW3JuF3Iv2tpN2H+q1bgKjte4stG3ezqsqE0FHDNAKUTCsPT
SdioynHCT6yNdYazCrr6M4dKXjOt2WPQteqvkiZ5ScVAv49snZbSLQ2r2S//6gV8
IxPQNJCF6Ij+M4tutpO0BUUY3FdlKDv6WfinYjucgpY+nPEgIJsaM0X8ESoV6qrO
9W/pZ0XvvlZ0PW0dyGp8uene3s8xcS96fvHe4k6Z3i90Xa+KUY0bciE0VHUX454P
78bvK6Mz1kSIZGKAOjPmMsJ6s6Rn9+GG76mo3RHSlBH1Vx17PL1mfr4xQD/na1+f
2UTBNym6eqcTh2Nl61ojXOB3C5Y5BUYJXwUr9wsShms/7ek/M1m8+F27Qm7/mmJd
fsRYqa4+reGxwKA5v5I+kelFzkaK6J36RHvNz3w5SQSpbo7EQs+AmV2rreZu7Hsu
3uw0nJxLCWLAdsWlUOV2UAM0+ZezTsg3bb40PlPJoKbGNcL5VuXM78jSras/B6I7
hlMT5lqAvbcwJfkl0Y/Tr891C2DOk0IfoLM9p57H7o7yI20LAvaqNa161mnNQS1f
le6irC2nhtmpWQUzASmXKMBAhiJzhAga2T4+SgAFMQL5bTPXcDFfDtNPqKpdN326
pGtw6pr70wSpnfqcQ/MbN+DUPzRnVT5MW+f3UsXGcjUxkCM2Cl4UAldxAnqmQKZr
6pJN6UtqNhG5HAz9tudk3lfBrv1/wedrkIAsqP36Yi29nb6AqIyy4sxaPv0iQDTZ
fVLNzMJmEk4bzj4Lq+mivrXnIwupKdiSdZrMlTSctcETqZnHyLbG/p63ovBf4i0W
EtrOr5bz/MPneOAbUmlM0ZRkYYb2EWIAZrGpxT4Y75Yaxt26m7jiKMosU+2wudQU
bd/2IUDQQYR+SabpDmWvFZFQpe9BTt/ianQb9DMRz4gEwE7xVPDQ0IfPKq0BaxcW
5wPzSj5v211aHUnfghlJakUEHIXCmCnCKCXK1X6lpZ0ks8hrU8Okbn8xNbN4BTup
VuBWh0BW87zM4K0IG92HsZvq+gmtBxwQG+4SM4rTg4iK1WzqP+iPwWq/5HQG3BNu
vPLMG/XjONMFhcGu9VfOfravVAsMeBe8sK43n8O/Gu1PXhNtBkSFm7N5pruofNn+
vgSB3aiOyfTap1X9Jpaj8oJ5XiupQsAg/+PDTBhT4tlNW+6RM5+TGre0CW4sSRsN
32nGyJvkLylouZlgOngvjaPc8SHhAHCzX6Oo1xPAD9Pyqn6u1J1e32R95pqri8H/
Eg0SnML5VgNrLB3Sh74nTWBJXB7CfzHAB6KGRExJMcl7BHLgXNpv91TM9sjfUiMx
Nn6cU8kcU58R135/hdhdiNecXtui6JuhVnC7Ldmddl9zuaNWMgUAL5neAIH63C6l
Nvv+WJ0Z42RpiKMl4xqIzQTrRrkFpoSlCsBmtyUQSnf1znGdTJcTqUl02+hKHxzD
fcCA39Cz67zPVZ/k+txwJeteNsjxl6j/YIxq2e6MAE3LMttN6Gpl03Gy4o//IgpQ
5O5yA6lIa7eMNleJ6XQomiLjRDOgTqCaIPzMO7kNPKlL04Kdf68sex7G9h6zY1Gk
VuLz4pYUepEXFUOuGIp9xujcRxTI/2qRdVspT4EJ8YOozmRuLC414HMt/6vkBDkY
TWBoX2H+6s92/wdJJB8dBgoFKZzon0LWVkuIQDUUDJvZbD2k+oZISKYHrZQRLKTr
AUZyF95V7Zzbgxthwmg8jikxYLUbaYkhtfZqbTdF+KEYnp4qL5SUTmPxSkbHWrxZ
+2Hwg8BawwDKkh7OSzsT1IWMMSTwLV7mFtQVQE6nGEkEcEAmYCE/1eFbXvAGpWOl
iKRPD71vCm3LEUfI6FnWqGUOIjqH9z3VTqzFX2fTpAYwHu2tOJP0jw4BydJi3b1p
WAetl9NJGCn4/CH+eN8KI6V0rTMR5xcGOwXiyUmYtiJhF3e8ULW8a87r8CZydFna
NyysZyWG84rZqc8EHtyGw4VF8ZZAKb+8VLRfgD1XXlx1PpXepLpKhQAKbSq7Z1G+
wDqntrtIm/kATUlAZD69b3nphvZHDKgEp4qDXSzdKu6hJzDoE0g0SPCJWMniTuNR
pYnNuK5GBO7ezCFjH2xKKwlgy4RYBAYW1lb9Mtvi2fi3RRiC8gS/pvlUyE68eBoL
94HhLkuvVLQGc/cqKkk2afEcjE+3WE0W1e9M/qpZ3DEHwzbprPyfJ1T/JIWJT779
cL/+CoMmAKayHyXYLmkzwuCuuo8wF7ia9RoTs462EHpz5+XRKq0eBwmsVfhiwJzH
XXEOvjNgXE4uoVIw+BPaZoYtS9ed67MpGoi0u0ZLbfCVAhJ+S1aAC/+H/q0ANTYK
VKOXvRImBwsNqqQyUQsHpzslxN62yqz2gBtwgdxtrsg7n7zChJjDm/VJtQKw0UuB
9eNnzi//YpNhzVRFA58HGDS3TmAmk1ODBVxpnXhW1sLyp5tCslz3xkNunbeCuJDb
hQl8QQ93GGkAL2SI+KB9RuLHw0PNx0iuhh1TQ4OgdgNkOAeyULkm0SHx8mBsV/Qb
zo+8jGwrA1KASeDQnseyxxT7Xg8a9nm0/CLLffhjlTkX0iw5/BGmV5bqvNTS/g1S
78OGXpQ7UVnsx5WqacMdECrvPY1mBHZgLkWu11plA7DmwMvpsDPJwP9/qlGelqbF
uMAHRUJzzfii+6EGmS6nBtGEYXmoylwB+FGkFA8FnkDo4nxdfmrQjKmcLbPH1eD4
wHUPtSkFqkAjLcJ35PuwihFC5D8ghjTcrc+Piuf9K42b1FQx1q5g53idcMwR54Dc
blh8N/+KkhboA0tRvsk5D9zivLaS07CDP1KehKFV1wVHX1rzcxbAhoHrm3HTMBoe
xE3QvgILEquTMZfToat2yKNWAm7514Kgznw2Axz3Wuc8vbxILnY16o31yBII/omD
P9dz6ENllShW9hW/qmSSOA3+WV/Z+iJVgKVYaMYyIY/0vr20pMYeFIiUKDnQ51Zd
0DeO3lOY28jFd9N96c7juVNmVCo8H3wt8+D/7GpYG5tIepfOqW+4BgMFtKPSeyuz
xa+p1S8wyLoEHYB5fj+wwtBXX2elXvbSCTZAGdicS8fiXBPL7ohDNy1suO2UinBp
7pWsC5JlmNZNA1rB24i+GGeqFOjtMuNLaYITW+8Liqm19gV2bID4iJ4XgOUYjWJk
PAWnlCumNeLuuAi4RUZltsPN3lyzqEFitFGKZKAL5jiurKHc2iFvDk0g5scRRnsa
jBtUHKiaHt5OMVPPc7Uq3moFWsxdzOXu83tW8xHTqYwZdeSVHk3/J+UOMyXIn1RP
yTBDJrzGlDLJRGnNh9VPtuepxc2AEUuFVg3coq7ZxCnXocQRf2vbFI7mCu/3JvRy
n4tAidiFfv0w1xOsCEeLNPLgjGZdfdXm8GTuiHtAv/JxoN/j4q01MDQstHeArgpN
XpYAqnllSKErYByXbWHRigNopgayVB7KzGAzlheYRPuyY2utXJLDw1EcmFTDcdHP
/ywlGMl5CNx/ooknsQPW5gBMGyHom4Nn6BVOMn7yxMkflrDHbLxrsWxOEkzltgkl
cbaBlddcdx5KVZs/udimGqicpLWPqf7Ahw08OmHfnNSD+VEU7XkKuyLc8t9/Fwa2
Nno1Uy3Tit0Ojj9MogfxoM0ziIbjVigeqjBzvC9DprJ75V0S+OM+r5ClShtbEN7i
P4ukM40DS3v9hnXiaf+8xXL5VWBldM+xf7VemdEc2tVMWkLmU/8mmsWdrakopt0m
EsGqFGk7VEvYacLGTEIbLSG98hLMpCsUaiQ8xbfckYNMlUetWKanh2bQtswRvov+
/ayc5xo26Nqugmm3QwCohyf4J0jWZgI0DAOogAO+/EXUHWjIFeFsbLnviHqWx4JB
iDAMLg4df78BWGNYldUSJN94eoAhp7WG+NooCbw/LqAPqVuP11wxdEP0ANuDHQFP
JjWkSrcpWCzUbxLJj9FRa/3NB0ovVJDuz0klrKYmQT+29Li1vLU1o3qZ3vSzv1Mq
1TZnH7vMj8Tp9KfhJYtr0sdJgic0WZ6PA2pUM/wbV4xEc9iuQ34339Tla9MuamL0
AENCfrfTRrLd2PP2cn8lM96quVF4OsNmZOl0wxuCwhd74Xraa1WO4YLqiix1hS+i
Zj62tIoMCMPZbHD5xmMsFPzq5DxBpwzUPWPcAhLqAelt5jq1EWfKH2yhpB2p0R2H
O8psUM7PasXfMckT+QTyJxo44dnL1ytR7dm+9Xa206r/5sIy1g510DcA929B3IBc
I+RWqnK/MZyVMQ8SzY93kaNjen6kbEBE1jQL3AMshhCtmF3vk7QBFRur4x3FE3Om
TKxMidXinfbJ15H7ACygyfpOg72ytqmUkxagGIKOlI4q43AYADnqJCEXlP9C0QfN
M4xb3L7AzA+cC355BiJR+RnrDD68eLn1jjXZ4dg9nO4Gwsa+Ys72Y2wOMS0mybC2
X4QxQqpw9qTprEeLCQwRvB54mY7dI6tlegyMeVpvVbM6pOk2SFnlVccEkMbSsr48
qN4SHlAuqD1or1yTAqQDznfDAJ/Si3spJe2QYE2n/ToPU0iR4q05qsZ7dGWyzKhs
EzJQHNZOhjZecuT6mpYnUfAoQYJfS3ra3ZfVTzml3dATfXlR0c/Z2tDbVS270VIB
4OhMKVS+316G3f/XsBDBnu6d7c1rdzNT7MVe5ddNJhCug8ZpRkGAP0YaDGt+hZ/a
fh+ggVldxWShLfKUELex6fwcOaVgs5f19LiM7n3xZzlLjUWz0crPC/P3FsobH0IC
jmkbfhOQLPJoXs3DA25z3om2gR+tnOJYGspdPybdy5/eaBYDR16ezh1cZL7wxwWe
xO4h3wvCm5/N5oCp66epVKdSo3PhGcKbg7VZXLwZruLB/P9DlvXHk3try0Yop9PS
p49vvh/+Fwk/wi5wXvB3Jp8wEaIKbCz+bY4AoosSclxgWFM6o0L8XV4IjjGjkxSD
eSi0d7wgidO7kkW3UgoZAKFEA8cwtRDFQwbOp8houW8NyMCiHg0q45l40A/ETSpf
8g9s9DvVaobJduyz/vIk24DspUyi8TOfbtbpGvCTK34hh1bBj6IcCvmL8/jqjZDF
98IeDrSrL2avyqXaDFOQrJIVCkZWxflrkg77gvQuNVJYXRg7ZsLJ6OYKr2mfenzy
BZURBujQA66dZ3XixD1FEMRcjGS25EmkkPyvYN37XXej5gvrCGKAmr3o0QuxK3iS
vXgmK9HsNpZAdhQItMQakMfTQyrIJrpiuQ+nUNl6tnu+EA+Jx3fx2pUijoIHv/Wc
lq5NJ3I/sExXtreQUVT/tnP3Rm3GNLc55As5IxGLyMicELkl1ERpdqjjoxsU515x
kvwdLwrX5RqeotHTKTFTKoyTCM6TV1DM2AIwCu996tRYs1KJhU2+WjdkDh40W67S
I/dgYMTpjGuOdNx1QEsijSDohS7BSFI8fCgGutRFemYFJ98D98kcY3koGzGx/xCn
welyeMtEjp51AKrcxpi0mXkNV+gsZDktZUjG6dtMvrFyhmpU66qKVwuGU79r4lpZ
UPSp9XxBNFH68DU4jW87KJDcRNdzD0CIAcWU+3O3C9eHE2Np8sInLw0v+uxK1/zQ
FRytC+XfBK30hRh/l1gZ0P/3xx1oTNcQCxtb2n3KwDzNwn1+KpTmk4KvLO/65k7T
FBpwxYCt90fZgO9HszUoB5K3WAytfv/aeCs+xDYNMR4YjcTIDhv2pY2PvrMO2cRu
fCpNhmWGqAPiAsrBWtdMcdYgImaQIeviX46Yz7dZkiwpoQNppVKLGUXcggYJrA7J
h5uetSRoODHHVkLIFXtiHkV9hNs1nwyDfyeHI4WCV/DuYLTvVL7aJFpzsU3/EIJ7
qXjiPjWZs04DENnLFImOAS01o5kOQ7X57ow4PYbbDJPEknAhk25h0WgDPK2olUvC
U3oSDzbCXFWLBzun3TEO8uBzb3XUbvVoS++9jXoBJxvm3Hn0eVvw4QZ4HD6uRpEP
PRQQKVJmEemfiNRTg+uIbqg/uVse4tgrnrV4tu2J6A+tD1dS0DIuODeYk2fFzcgS
EnhxJ0SIh/f9Mz/la4d8XShDb9WgYOATsOH1wpBtemVkHTqsJT0HD+2J1sVrY7vP
Pc9GU/Tnim1l2QrdRwrJaiIxb2ywwpUM60aWqf5TtZBI62lrpfhsUjCQ+Jutl0FY
LQpOx0e2Z4jvcmbHN9DVXLWBMp6SdrgI/XyqJ0oLezrzgGvfdB4NWhhn0Peg+rnQ
X7qK4jnHYb16CUIwFvDM4OfojzNJx9vQBiHpsxDXaS25udY/Zid7GDVBKQ6ySRsR
bIlzLlpks3+QtsWpaiswDeZcH/ZfZ9xuOj/phonHrgVQYfnIuV5dOApJPM9GRo64
0n2I8QSSVMXfqj4GWmhonucKAFfaBEL1jFDiiap5e0PEwH86jNFu0PQ3yOcYsJuP
+9HRGNVfBxtlU5fOBAdoEKg5IC9msLCCGwR9pOKvnkRq8vrdRqn9ZyDheH6kgZIb
/4R+7fPk0qa61c/dADnIgVDwFXWEavXk7jSxiaGzae8HonXVfwx1gHpSQPM26R5P
5X7ivc5EZC8nBcNUz1acJrim/wuIgslIlD7enfYoWZGrkRKWw27eyc39nvHvI7Se
KPbPVZSXM/nRjECGdIpyjLlGZNO5FXV3Jxcc8i/QdJEmrVsBzFCgs51ccUHB6y+D
kIA/YARzHSJuepnqX50pIMmGYf6SbeWBVzRmU7d5n+AOykQ2fUtLPgPKBoYlBZJ9
3wHfgL7tET70W/69nls+NCo8fgQo4ni9VLwUSl/bXnMUqePRyom9nBYhn9P7ajET
4zZYSzkAu9FtNLeMB4gx+6M9wsgQBpXfmBSoBTVJ/qkmJ9BUfvKs7HcBiMAML9oi
ZFlz/R8qQ09r9RyTf5jDDxPu/lUYFl9IsYhl0GnJDS4FjeOKNbFiTcFcbNaMT+ng
7mR9DJHJ5qHHM7tLzeqgdOJFqFm8+t48n/rgYT8ArswElad87wvaiAsaa6qieHR6
OBZ4rTMcyHmo2bkX89DPESkOol8+hJw3zCvquqLpnw5IW4HoYTTqaeDMAbuXSm6j
eOGgKdTbuEQS/a2Rn6YgqixhVsgrzKmBTmn4z9bV7VNqH3T/ZRxOPB12VDMMO0be
T49xRH1xDmRiiLpWfoQIfRzKhy2YgVMsI6Md+vSS4RSOkVBsut/Pty9opb0ouwIm
E+IEFHFdyF367puxyqxml0uXEcKhywkNuDl4MhQZGQn0xInJcRkmOCw3jX7cbwFJ
C1VV7flePHHaCHvSFHhIMEbL7qIXXY+NfWKMxALeYvP7yPvO36dGM3rEl1YHpj4R
EVyQQ7/2Dc9aAzWTUI/yCafAuxR+9UjvaZ3xo30frML5AUi21S+PKXfMSXyYSHut
hlhR1EYjsSvk1N+G3LWs6SR0H8/MjD9MgmuRXOWyosyP8JGsKIJODHZqLMHQiyEp
GDuc3QTJEJwUmKw1GrIRaUvLvvYeeUdYknwPvcD/TwL2/5054aGWenmGNF9JKy0B
VNt5xvWJa3ij9o+o8XIu3Ba17O6To7Omk3TByrTELzF+R0NmowA829nTMWwURRFA
qL796SlaL2UXHzXiUHokQCwVZaO8Gu5RO+fYnEvYaHKeh0Oe1xA4Af8JZvt1f/um
HHyO63Gc3B9nqCQNCeJMX8oKwK3ShpzcIe7gQvnLnrDSzBynre8o02AjPam33prt
cMtD9ptk22bgtAchRnWDZ1XHb7AWFJEbh1AaDXz/Sj4F+LAFd283gG+1wyfP6i5r
oLnjmU8TaPbjonxqtI6xFY5ekW3A+liKagh+fAQcKSx9ohKhhszQqlNgaEnDskCx
UmBgiFIK9feVpFG832eTmxjhHpd3Ttb5453cNfqKp7SNzyvdqV3rCbHssGL5zOl9
hKTZUn5GURVuGksJ7ULJIGQlpoYCSxn5eDFZNIqg99V178+iNIyYjI86hYuoo/6G
j48WvMF2Cyzi1zB3qA9e8DuVIcbHQ36KZQ/UrRZsuC7j3CDzmUBPPcR3ME1D3MWg
+GgnB/DHAcpuxWBqHdKAaQuFNRhb0j0daBs3O9LlTickdFqO9+wd/7kLmIm7Z1PW
7EHMf2+xwe7NGvNq3qwRHY6FOI7eUD0r1omNgH/80r/W3QIEMr8nHR0QAvmkzy0f
EO+qeH2+566g2Z/sFRXWpreRZyp2Kbwpqwv+1D2IrAhX0C57L1V77QMSalJRXjCg
4CBdBg+sadulxOOSPh0eUARozi1FkOe5f8otSUxOTMj/ETxsHIWOugFSUpoZSmEo
fjO4CVJn4AtBTmHDrnoaW14PiEs9F2YgoLYpciurYu6DJSCfGpUKlxqlRtZTL55x
qzA2B4CSsTkG0Ax6DfR7y4ZFIGjIkznJ6dxJEzy/iVDZ4/gKP4nLLnakv62VNtp+
gzcUBjJ0MbA3afJgR/pNg3h8G5kxLG3NIZFkcnTiD3ODlAL5JJ7uxrXaYUhhnGVV
HQ1d5xX5isecMsps1FPkoJo36XlLqIo23UDgXNP3S+S5cpJglR2mqTQT4Q2LjCoI
C1gFZHSsm8yLcIr+E1m8D1T/nhruSBF+OQm6XzacSfTCg23QtnVJQQH/utyach1u
2357EzrzmizJBamE6QcZtilQSs2D/sw3fGjYINB9PIfO6nQnU7PFuLnTW1w4SaD7
OsOHJ1miElMilFLT851kgsda9xvDETaW8cSA6djCTFSAQZ4mmU5SkR5UxxWUwffr
6y0kJf4Ya0O2/i4JBkPbytwUSU3J9zC/fgWAqFWJZzR25hNpdhmOGGHxiMeUTFs/
/INPJ0FHktM6uDin+esFiRvJmuzJN+VFipVDKBafEtzISbbXfKwdvKmcTfxeDS5v
bAesWjaBguS/brw+8KaEGlJVByUB6UACgpko3WeFoEAzR5cZH8WDS6jiFunLWvDV
oGeOsN5GZgAh760V6Bs73LiOh3BAY5Q5jIf9T8zB31wjeZIf1oph9fFJk1auOLMm
Om2GfvVMZQj5JnRJolU4bIRNXbMMZfJ9AxeDsBvwzl7hdblteuSHIsOS6UTXXE7j
qCKv+sE6jzNq0eC+Nodn4F4Ovy+wR+3xKUKjkCBDQx3QhiNrALQfJG2+YCahTU7L
X89J3U0wYLtLdrK2PyAs1EHr/WIYLIaEh/zTde2T0lKNNcMBjcMTYe+Ko7zYHL9E
QBdxuvxf3vLJKb7thZuJKIUvhla0L66b+Aj84gcO+E8pn9uBVQQ0szt7AIHuoong
Xgx5P5EeAYPZexawQ6IjYj/N5h+AYPITzglrCIxMBOQQ2sk7/JuHIHjB0Ul7XU/C
L2YrYGtieP5cXZi/U7mKhIyn3FHNrvtlS1Q297MzWGEWaz2Tdm0ngBaN7y+mxcm0
gVDKUn3oKNvuUWzo1bznBbhYlWfQsZYS9j5u6JQevjw1TIJbsnz5yCjHiAIp4qwB
sSV7dSL5Zco5jyD0e4Ap+bpEULHzulhB/oCv1qQVamfK6cVL9gWL6wLZKL8BdCDc
W9ommoaW7Tk7oBXPIqGlK9tdhUec9pyZvsCY1MlVatKDsSlEM40gl6OGEP6hCkcL
0BWI0aIiRKZgKApJXtAAYgWOaHfBsr3gqVQDIREwf+bhOq88+QIuXufKP1iAj/Cq
ZhAZ+AIXrctuLj3kjhG7pQ93VXZAuoBj9h9MRa1KjKdH+9k/kVpFQ2LYWol8lheF
IsKxWjqdhTXBAErXtsgCr+f02xJRqJqOo4cedqQUyZw7cpNOks5Dd7xtl8i8Ocrx
xzitUOXcPvJtRKaOattFkPN+7QAWfzMH5azdTwx5R5MSjvwjUb2kGQADopBK71JP
IniOEU2kphjAh4zlev0BF7bGOR7QU1rj6ID9a7kqITHBPy0/skobAZTdEfeCoLqX
xAkgoe/XmVAiufMcsHipMK4nKIq8YvCT1B2V/n83hDLxyhuHOWajZrOH9ED4nxMP
TxFORCBH07DpMTWegr2Nl0oeiBsjo5/ZTmH1sdlfw1beU25weU9fjSh23WxSD87H
jtkmR1dahuLQEzB4u08/4qfpeirjti2nI0TCj87W0d5LqYyfuZuAMuSOMmDRmlSY
raJpRICDK32NHtnABjh1YipZdxWD4HpS7FtfrZyM9AUgmuM5Y2sDrJzK/OiqjHrc
o5uB7+ebo/f3OCsJTiZ61t2eATlz75ds22Km6ytj69Mbc9xmq3fZ6TJJlGdTRl2A
u3uN+mcfUtTYdk9ORGuohEPCihiOxDwcKs/VdLEXxsrjFY8Ezpkqju2pbqmWm8qk
1mMSlH2oLr4og2cG9EyPbs/XMDqwzt2OMEzDFAObhCe/E22UqUFSowaeNoGyOjUj
m9TYPFI16kjwrwnueZi4Y44fU1LDlDlE0oPRI6CzCdZkwgUg92XwsLmZGmRVdriG
V4gkcgF2F9qqznreBlUOznnohcbWEB0EF5crQvpwGiL6VSDLpJlGkcEncyGM8OFP
MUviDBqIsgrpjMopRuGjrUvr65fQgQcbooKDt/9SDgw3A9kw4ETwf20R1un9NY3r
KA89eB/ECcNUGbGRD0WfaFvO2m07TvT9iXe1jgvT+YKHLn0VFyTvMpwJEE99hKyS
ptH7mmic1xYu7IH/HJDYVRlrvYhbcR2LDTpwMFjVIgTCivSMe6Q7vclPnQdsG/dc
nrDJBewgK4KyrZUx/8yxl5LDbOOVEYMvafpC9uWK1GCrm1/bTWWs3EoT0Fpeh30I
vvnuxI3TD0KO4CmdHqi4lyo2UO8hFdwgZHyHlupdvAE7Zv6RQDievwfofFmXbDOv
2Qj4KuWdPppantjHwrn7zuxqTYIUP//Xoz/2tqkrsVyxMuR2LMVNQxHa7WU9Gzx+
56o8geyOvNjURbqMf8Grgc7bHEIBcZ0KPp5DI62PtYfVHpOFkUMXv5I24JhN5PAq
p/O1xy03p86CWcGarHtO8a6stsumHz87BmjPS/SNT55R7b0xWq15B3qhrw83MLn+
9dqzAbra4mwMeQI/COJKcvUpj85Lujv6RUEHyM/2u1xFPSyjTk6zrVVAV1P1Q9Zw
532c8RE5f9pPzum3q/R3zsUMwx38DDVbaVjWr3qiL76R/M3B45PPINbc/5BSxHSW
8r/ChPDaif74P2OPyPp7Ruo1hTQLeBPsOZGW8g5xEjKEYGyvP/HIRctc8jEvcB9I
4Hx5ZnUIhKQB84cb9aSTJ4xY2ns0LCRoZNQlZLlZC07zNlHDa8pgxQ3veNmFvqa/
MIRFXDYffrK7aPv47qDQLTGulck0dUbgfGn2+/jFyNh7ZKI8AKqd35rikLE8fJol
HMga9zXDUCJ300qzKXj/tA4Xx4mdkJ+qcGanKGrWIiImOHGUZswIKLFoa2kycqC2
/VIsKJqVDV/S8jpa7GMlLuqPBG1dQ9Q4dvZPNTJwci7EBVXY5R0lCRJwzywjwsuo
KqyIxdlQUzYxRkcizXtI6sIIL67a3Z/EYz+RDtV3MOQan43f9KSLXLmhyulBpUhc
42s7EciqBzCbE0ulhXRK/qdR2G8uFcTr/FIJQx1GjcjKRz2aKDelqXXu2V1UjZQZ
1QcPGzqBzIgDzeO1/XC1+S2QvCCZLIBqGxJUgyjDEvYYgnUTUXX6tXpDAfcsChyJ
bmF6sCGs1ZzSSv7/d8zVjhZltkqEjolIwnXAqr13NOZaHmTYFIMudRh1amKy8Q3V
AyCyHMY2M4QfXg0bQ6F6DYiLEmZ5oPoBg0oAC73dp6TXouWCG3BNjDfCY+cfY1Vd
9tbA9L4OdoIT62bSAcCAMVHCosVEbgHMMhvZKXUXilWA9HmKH9UaCj+cgixLWmON
6ylEhlE1RQQhtevYyNghRuoG5uPXajGcg7Z8NjxstpeRh54IyYQLdPAMuq7gia8g
w0Am1fJlq67TQMdR+0SgFjBh/YcKucmgP/f5Syn5eJLcnVJoNFGMZrDIC8obp6rC
2yS1SSJicj1hRCSs8xm9u2TWmL29oetlwrL5tQOaXrPk/sMLY/9YpWWow7q+dUcq
l4Zhxnp/RZoFVpj3lJrogZXNXS4ASyhxsiK/0lxN7AXhm1jpxuIWydhkVhvkQflc
g6f3N/slxbl9pDcuaFfOMMcsDK2C+YvGQhPDZXT4r+s/qpu7ky0UPFq/p0fhQAlL
QgIvl2kz1gs3u26i8rvfIFGGtDU9Q86rxVvqM/Ze8DrdgD4mP56rzDGO8lCx1xpa
WasT+HqtjffsIgoMpi/QFfAgMgC76wG34XaXQFM5ux4BFLwcbZJ/pd8+M6OD8I6V
qruyK4FWCOCEhr0823SahvvdBE0u2gVG6D5d478X1NBwujVsbneAWL8ERtu9gajB
7f4DwJP3a2hvbCPSJxoDzYKtZBE3h4XKTlaG0d+Nrcob316NLpdYkpitJqFMzpkw
hB/5aUsSTPFi1Fra6duqvaT9D5Cfu1G4bl4K0lEBI0ClOUF9Dq8NT0EiJN3c9wyX
t0ZsOYhoNsnrY7TNMhjHn/WaMJIVvVHNTeIDTh+VY6b/Ap0hXave5GwIT//L7Gi/
jZHJAKJgeMtLQL7WZIaGojpKwIBIFjUVsz7SzLjc2ublToIBBKudPetrPxpSFEUI
F9tPkIXQjMhrlMMSZKd9RUvilJjt7EYuKh6WwAJWXcAtogizLQibdglzTJ5I3D3b
ZXRa017/evz4XorXlGaM0aLjRYy9eFr8AFEttefFlB/V+sdtvjbf+Zb3vklwZQyT
mhH5pqvTV/NHht47Zy9cjpp5IMY5ywzY4DwKdebs96hsElCkGV6u4I4SLyBGas0q
odCzIiKgLy+1qW9C2SeiCHjrYEgGOFoZmFHU1QXwLmqG8pm/5ZO45GM6siY1f932
IwsADFqpI0/Rchn4VmYg7BEf6Qzev5cLC+Lu5CtPo/02v22V/chCq6LC9Hsyx2Y4
Lffnaaem7Buft1ySiXhwDWch7Hl8PUY+p3lM0dA27H/C2us5PeQoG4ZLkqLzrOx/
q/kLUoJZCye6b1Lr+feB7KqRqWUuLO4izq5CvL42NWu7/SVtPl5Qm7Ku3prs8wrv
kCKGEyhB2jSJOuv2TxssHPPxN/DR+HwgaI50yK+HNr2lltrvNgSjgzOfem00R/dt
RUrx13P3mRQCJz20aZBEKJDRnAqx7iqEuAKzvvoNag/16YAUnSVj+V3vPFo3H/0F
keh4TfzJ+NI8WS5eHthhDMk49T8aFcKLVQVIF8WgPEIQeCvGLc+tXodcV1g53pIU
2c0+Uw1hNIp951DUdMDEylRhZRxFGhSnNzHmuTJcl7fHyVc7xwe69sX0Eph8nsY/
q3W1NNR2hl6t8hdmyvuAMRO7lgCqMxUiF39+bWqTHJKxabu5rZBXmSimkPPKIj+5
q4mpRkcsIHFz1jjt327DFFsaOqvWaXGMgdfLFcw8vxh1wBZUqtF3IHOPbW4+SuS+
PpMD3hIxlxxyam8reYHHKvtOL6/RwTXyN6nRDjup/KL018xlB3sUPa1KHf7LdmhF
voA3yGw/VCDO7h3DqgZB5SflqobRzeuSWxmSd0SqoQigcOm0VsATn+ohwn7NZNcU
8nrEO9qQwwdBkJzGRCe0lGtzcSn3cmpbYLk44Yp8qsIOdHS25raeYBDhTssY6MZo
LjKvTjm1hDkXxfX6wHg9p9kUsCjgRAIgLv38x7DKkrR6EGTCeyUGNetGisgglOc2
MJ8Mmmug7P0CAgE/XuayA5vQSA1Y8/r7WmGl/wHDet2/eI8quto7hMP+Ii9jFQkU
eGTW+WEI5q1kTk48XiVAYobiyAUeKY7IcRdqI1yYAMa95yeTcSwKtSV6mPRFgfXq
RcnpPBi92SVNYllRdjRcTYAs6QSCwewW/5tZdsr50/eeI++Pngt7wBVELJ8Aaafc
LoTOM2vmrVOolQop1j56q9HMDOXrj0H35X3SZdfJKXXDcyhKBzNP2lX8w6HPpkfZ
/tiGEHBEhDovw3SU2YXGxK4Omaags2jcicbOJHBPEiPJmYdheZlpgu9pHUPfoRn+
zxSfBHfC4xo+K6ZdEDs0SBq5pqCCnM9ZA4Zrht//y+sJ72LdzJc81Zeq8VlpfPcS
TJRuy4wyonTADxBCda2OVnIYzfSw0Mto0j2y29UY6LxrmWeduGLvIMY1OJeCdPqU
GnqLZto/aHbBumwwF1o2Atl7zk5HsOApCtgsLGSBgvvFT7mm+gdloSvMgQ+nAupj
tD3iE0KVTpH93EfEy7DAMq0gFtzaIdFHObSZDqwQb1MYG03wxg7EJ0xcaruMb2My
1D1jZ0ea2L/7yYkjGfvu1W3CKukE+CeT+CWaHJJdSagweoU2muD5CppVPxHrXvFu
Npem1uLzqIN0C/mB6GHlAnaRx1GzdTsHWR7MQ1BnF/ScxSY+cgxNvz/v+M4i3cXT
LLzKZfZWR5JFD2KxNDK4g/zUBzKkyF1FagkQG1Qp6XFjrPYhKsSrCNF4DyWmj9zO
TORyuWDO2jEQAJCtOLlA/3+xv2yDm8F/wtpPxC+MoJKbqrIxg0L7hs/ybMjhWTCM
WvuTKQ9hSz9LeP1UEy+vdzUbh6OD3wPBPDKq16LtrnsR21cxN9V/Ev4NCUOy0DN3
+/p8ON+gmzaY8vdyt9aB3MSe5xTeeDNsMUn+LhDtPFsZykK/Q4/6+LjDR0Ssd4qF
3pAoEW/lJD0QWYGZIH+R+beBXfmq8o/LY+8nYdULvCmqmzwqJX61VmXlbRiDE3hc
HU90IGdxgZY9rDxcqwtxWsMPbFOidL5ct3dQ6UdCn67iWjU2L1zd4jGr5ZVtXJWi
DlAhpXuEjwwmfqF6rExsF/mLl6L5BqhrpAH8X+EhgVIsuQmLlCUkEJ6D965eeogN
gLSFX/mnjBBi7HfgjUjkcgCTXF0S7EZ0v/lfT5YoC4QMhxv6oL8L5xdnlsErHfQr
2dzI1Ahnq3YcWD02BGuk+k1oZFNClGYo4O1nrhdHHybMqV9Q+tAI7WozN14B+4i4
p+uogPDn83CTM77OR9QstnpcZjXeg2ibiHJ0ZXDOCAWwwL3CC6w1i9Kjc0d48FgS
zkOmChz/Gn3b27u0Iog3Ecl223XveCEWz3wAOmY3sQxtZ7wJ45Bz9XUBw6MjJgbz
+y2mN8r84b28jMvlDbpFuMOTReN2Y29q5yZcLoFmDhcy2JUzKz8BoF7NRzQjtUuM
E/mY1rhH0PS9rOWSOFDoY7DUM6WROdZMFgUhkKzEwhwmlgD7FFWckPjomUL7vYfd
1W66hdOGllqERc8e40UsxplQ4OMpDEK5wt0JRg65tnpBtN/tcR6syo8r9tYuB248
dzSMuVIkE3gYft+XVrWZK9CnoWLJYtuDIBWEr5OdzMhxCXt3cgQK4UoOpJsM8VPD
CEY29K1M0ZyiCPh8NW0FViseXWqmL9DdUmGQthSM6JYdt5CNrG8ej/QqeoIVfeG7
JZO0+tVoKc+PYIoHQWdT5TBaYf1N/uVs6APYOD4qZaAJ4QIowfiSjCMHh1IFVUvn
aYBTpJ1uSsZH81DEosZ8V1KQhk1XWjqnsB11s3UFrtxGfMyAkP0NOqRmxTPlLssk
YtVnHMU0d/PZwvjj38bzbzy3Qi+b/KFy9qr+JFchxCWUtamg0h2B+ssfnvw3Qyk2
RxruhygGOiB9Qr2DIAquXrOspARbpqfg1pSQQ4ByG4MQF8gG1Drol6kHSRoWPCgr
AEs4hqfXNQ164K2TdGntkA0lctWE2SdcC0EEZuFFCCTSEZEiuWRPgs/Ij1UHs3Sp
QGR32tw+6q6XiUeEsglKpFI23tQFVaKp7/bD8LfT0kl4yAqXaTZbeOH7kowbp151
+5S/gkxRTbPWhmhJnFEDlHv6HXZjto8c9ls59pxVdFOxt2P/RqbM/2yjD2qeNDh/
ssGoQSX26u7vvXldPpkYwkVwwdofmkJZAergKjvAC850WKiumw2TecVE2tLqHQcV
VOoW/GMJWlyOfInOSNKJiK3BMqNZa9/BSm56VuOiyP75mHwnaL4LsaiJGXLga11a
jMw1FGtE5Q09ubkAfBqXeCtJ4L21IHWRabVlnn5O3l5oXkDF24Doqdrin3vWU5ti
2M8CA74q5swm0iZc3lYiaB8aTcg42lqP7P7BrwDiacDwUnkIFxQfJpBvBP8IB5th
+IvhGeHsIA4JIdSV1s9GsIFIB2bcjeiTEEf1+4t4sfTw7y81GDfvnXRLM+3kp2iW
iIGsGvTDA7q1SgMTFE+s2CirUpz2cZIfxR90EgROg/+As3UnO+Zj0cuT+rh1MlRN
a14/EYjSM+Rsf14ySPtS3On98rdZnf/QHn5eKcXbsp6Mlmqoc1t5dy9qrwFmv/lE
Jk6vcXgeStHXs7yQSf94UecqFD6ZVo/xc8Ex5V9y7SAG05i6FrGDKe9dtBv+zYOE
5UG3YUeW98IAcD5ZUDk7xCkPyEM4Wfn6XARC9gr82QRltR3M7R1n5h7nSVSLXS0h
7rGC7EBMZS7KD8wKc3WDvB0GAXQ860iqPAXuKQ8w7+uJqmFr2rGS9ig8y+lEYQhw
srsNyaSsHKOF/hvXqirrcKp6Pp6qZ+swTjm4+vV8HBUWyyuHo74KKEqLAov7iUh1
9zOShRIkDkAgrJZAWH4kbq4DpjqEKO9cpKltBJ5rJHIPaboruRb0YPnQsdETv+eU
LG59iLUzC9U9CHm64AJ7QMKGy2Ter32fZ9aWH1pZOUlwcK9KrbFBFVYfa5LvgJ/T
FfipjPVtzdlLHI3lXkY9/3ojDMlQeNqBTATDZZ431tAElaGuEGk68teao/t3wOGZ
knyVlFo/x1sVIKTbjoXeuVdEywmfhnExpFnh+SH+0s2aTqk6BvVV/h1S9Yn9fcJV
7TcKQTH9s/gB4+DWxZTUcV/swFUq5Ujceqo7RqpfkV4sd/aqU2ePAbLX8ADEofaI
e6ZvCPJRiUqu+L/a1MzV5EONo26PgeoYiKfDDJhX56cXr6Jt6/QJTT4qVg3n4PI9
4unggGPsHxsmK+Nxelr6XQG+19GkRusYoXB0KQD+c94WhAd7ZWbBzSInEvDcywJm
fmsT6njnh/MPcJ8YilmhOpGsWwuuQflrLBjmNKm6an7/k1HeJl2ca0g+6/INpEUk
N5iEWBJk3eubl+qJQQpG/mna/iwzfWZbHZHqz3v7CnBfiOs4IofBimHwLia5t0V1
heH9IB4BqUl1uLgLDwKFkwu/+4t9GSX1Zkh2fp4zb/ShCUdcqbExGWfHOeFbc922
7xolyOO6uIKUnQCLuawbhbi0HnNq464oluuqRpTBaq3WhjI7znUd2AljcXk50iNN
TJHzSJvKoSRjTuLUvVhXqbHSZgqWu1oRhvW8PalT95oE8Lggw2l+nU6n0H2Or5uI
i2t4zRayESPWtG+FUU7gYY+J5TXBU+/LSX9dxyLeaaP1aH2LA2zyMH17ZYbImPQu
NbFgtBlqp++T1XHkN0UlZUtOkZHszOEz+oYYCCpoNwzdrcAYWU8u9Otukt8g1ccd
AIZhCFhiDtIch4mBRUWI5jfoZLusykuHsLz4WQnlg0ITxdx9JSukkVJqN5MZy2bD
mJg7yDfyVtayCfBT3ZQerzQ2BRvOBzT5YM0BkQosauAY0KVlPREOxT2UAl7QbAji
1aOM0B6sD9dv0WGoNSSEgvtMhiJSFZItE4YN/dxgMRYjDJ/64Ah8MVM99s7g2sFj
XRbEVD3yw08yJMTI/YPEEThEgvHhJmYtWCIzyWYartVSF3hVfI05yFHLMYYU1J9n
4dnbDmtVW4bklbsuDluKAJhg541JidPUCloWeFxRbXf9OOYwKSAnS2CfOLNIyoqO
h8vuGHMIWvx1++1vsuUJA14t/oCqqHG3Sg1dRSdeptEM3018Z84AyBRzPRf3Fd6h
HXy5HVOekm3zWEUfgQ802t7qsYIGn83yWlTK3YuUaH38ieb9FSBhNvIB60WRh7RD
aalOEQPIxB9N6L1JfcsXuaB4fjciuUVHXVsnIPQpwepQWWfV0JmZ9xrl0lCCdDHP
ejJlm8vF07LkyMXoKV6gB2gxPksGB6Kd0t/Ziv9mLlXSto8FqcmI+XNSusXHbTGq
jyBfmZc6jflJQacb1SBYHvH1Kw24BIRYwDJZcQpcQfCiYV04ABPEt9W/tLgUsGID
4Wj7S3+jbt/zybxKnUPJpnaUxHsuRK9HlWaZnqTM+vEt9Aj8BvyievX+FF+VYT2P
IvN0bMnC52Y/Te9MeFpW8CHSlup1Rn3ixpKtStp5Z/TdUYapMP9N3Ek5flyGoEIj
lDfnI8cMqx17+z8Rs1cUEkWsYL1NYfAdSSqk/827vYVszVQydL+T7uN1qWYWP2dz
k0wMAXvxcnrO2YvZWUkuHbosjOy7D/LuGBKbZLyRL1mFsje9/5kcG5G4zpQl+JAg
MSjjwzTKK3QCwLISVf4AVyBqSFbLrpH3YXmBA3UKo7b2IbY7eviFy4ZS20XEUeCr
896fgfWm23mh0lRO481sspNVFe7g7lv8s6bDGYWB7GzRNyvIs9Y7AScqW7wO8iPF
8Ml2uPisk/IikQ0D3S0hL7GTIvoRtBI/JjO80Q69emjUbvhSnU12gDE+p/P4VS9+
LnFFAm5CUf+4uKt1rG2lZst2XX2eN/Gds9UQOjmMMmokxp642VV/6/PS1Qi51fUX
50TIonBRttepgLuxnoFAZbazvTjHplV7UA693nYk3+TIJ6jK1DbedUXqgUfhdrAp
Q0Yn1ue/4Ojq73zsUyTiAnnmsvxE5AZ/SEP+1L9spefD6/2NCExaQZdPkm9d7dcU
/iZ8pIiQ/VaaLAtv6ETA1B43wbB+W7BiEZPb8fuBo5zApXTNBWI94OaLfjeMwqMP
RnzUKqnHBlLayWZ1FHtDdNpFi7pbWGEBINRm4IK1q5jj6qV2JXCCiSEXkc/jCq2E
U+GGYtldkQ0W9wVSV8iZsh1WfoTgjQeMAMdFPi5UVXDPAIslJJABOtSThPqt0qFe
b/UKuAU2J7OUMWJT8pdimKQbNcyjKi++sC/V/30dMQqMlGpDulzUulFdeytQ8hwk
lbGrBj6DLubBlMYrKhA0a/7cpIZhJAYb//+uH6OvkCnib6AnPk+q0h2+5TAm3lct
TQ7839S3iuMLm+LF2GUAkb1t4IqGLd+rBfCCL/MxK3mv1cvHfWIiPdg8eu9XmsW2
5fCJlK5XStdtEyKg71HXQRCfSbICoa2/a3YS4pj4U1geC6Inys9QM3TTdkMLjFI0
BE81rqK0MuOXPHdE0+BgsZ8F2+qecxVo//rnvUIIp8QJltC6HQf0J7QWH86e17x5
P5fm5lJ+s/iAkc7Wxf7Jv0lwgGcFSF20Aj0u0hyQ1Y+9UlmNHMdFSINar3irbSF9
v8IwJP/2PsN1OToPC80XLIk3q678bZunC+KZ28rfkYnQ+7X0euo9tBEMYUUnbAg3
O8vLPRIYZOiYkZ0e4mgvDFbX0YCml8zgWGlEjE5wSz7nZ39gpM+K/rgOqEwktIu6
Vo7BVVkUEqEMwgt8b8jBJED0/lowEAbHcGiL5GEpMgfNqd5nldmKmNtgqnHd5Azy
i47jKLYm68cgp1uRpQGcCXv7MIe+m5VsUyOzW+mQpYYyd+zU9xeIRDusQ+Jm14US
lL2kPfG2zg9Alingo812Wo16Mq5V149I8jXa+f+cxWe0fa+htUWQa8ZRcIKlShNX
KnysXSY5mkit7sxm0wNTi1kIVFeukfy25/hQi3FgxWULEpJBMa01pdUpyiEM/IpV
rn7LvrlpFEgvGCTorDRKldXN1wl8JL5ubVdAc5V7KfcNTVNeKUOlyIvdF23JKU9V
Sdwar0T6OzTT11bOqA+6WS9w2/LoGXu8ih6RXvMy1pKRAJbDa4nAitOCs2SUuGzb
jCiOjk59rsrZAqd7gyj6IWx13TzC2zymeZmTGJ3MwdfCKcsp44iiDMHcOcyIf6aj
nsmnyHHXtf6hiUQ0nZXaA44Yr5Sj1v6OuynPHnZJKxkTDGBOQvQ+RMdaRi4gfoW4
D3cH6QqckIwi50FFt3qkJZAiqwge8NxXfOrYbRKSg6lkMj67idqeHN5QD2UIAFb6
a5B6+Gwcigg44m6qEFSR9h8wi+ih10Z5PP6BGrSZb3qXiwm7x1WPctfGnJqAUz2i
IH+rVw3gz/AhXbFZg0oG33xOpNRmXuSWjGUc/kkINV2QE87+Wg02R2Rfyxp6xXit
AZvKBkei7EYSCIPKs8K/X24yoPnrFFBkURXDI9F0A56OAOSSOLvCtjS8XIiO1sye
O7naUHnlL/nkqqYCzdD3qawvKFkkhAUnDti/qqTYkVh7dy34NyPF+rDsd7YcAa5G
NOP/CWYl12qRYWhCVXd23K6neZZhFpl3vr37+XMasp1CJAsMiysUtUD/7xRa1LTH
gO+ZF+rbXrdZt45UcIv88boaOBHS3emyTwsAORnYy9zl30ZzCpDwVL+PlzPCcltm
povW1MX6qtebR38kUHyzBeBDHPPtWFv17+W0bpIRmrChG+3sMV/v63dUEOOTFzbe
11HHZiYak1eOj6IZ5QT+Xuc4bVqEaskA6p68ttVSulCBMYH+ODj3RUi+CjdhBnHf
J0z4K14rR4aDy2rYGg3OprM5NN1eW5y8sA2zP061fn16xv5atPPiPe2fMxqZlPH0
b7W8Noil+G6JNEETs3FpNLHEO7TwrbWhEuC/4SmUlYizUJFt6CBuoxIS9hUzj6Kw
K1dY7zrhHHBq7FAIQ9C73tYhRx21Nc+SX6+sRPg8F8ChANB/dhHGmwfyp+NvTQ2S
4vcxMx6054JN2PWYLI5WnRu1r6vU4YwUevNT1L/GEceLlx9dmGJPME6x2kUun2U1
pwuWZWHx3nJhHgem1ZdM8o14SCawi7TveVwvWpgESgbTv1Da4NKcTjKbXYkX1Hl0
bZZ4H2UDNUYfLeqczfhTEa0UC/GHSqMTr6dKufg+vj5Wu0opwNzgY9HtDBgdR/9S
dZhlMDsC7XAhhoL01XbvlMuoSMGEK07FaLItal1gKjjCylAMN9cNq2v03tf3e7Gw
t9aWQTsKTdDF8jnwkBUYYn6h16c5rl+2rTqA/trWNs0rrNhP4Gnki3HmRNavSA3s
H6AKao2HeSh7ZZPkjejEzDk406BPP4rIWR8IlZB54uB4qz6qY9Ievs0rZP8qAz1S
R3cYUbqwo7IvzLTHP/ZKkkqeiTAXTQDXf6nPAjkMmiolBzipb4is7PIU8Q2UXMHC
FScecTVOz7/xPk8k1o+ObrEO9xu1+68NFBiMOgO/ZeV0r9G4deL6ElCQjB27pPOT
S/D8s9rzfiUxcKP/GCnyOrY0QvPf50uFbDqDVEUxJ90vsGsR1IziggdU6EgA/hrO
GGrsJLuP06em3/B6ciTiuIB2xMFIQAHz3hD6IaPEpn1KfB6Jddcj6fwqo10eTiPH
87xN49hx3Frp4rv1tYkc8QQxYh3I6eG+xFPCOnHHhTnhS7yqTzLnVhjIgfMHOQCv
03jHJ8P9OmIHqGwzJ/asopwCn6GoDAuZ7PMV319gU3ZgUp8cdtab7C4mj1yP00E0
ZVSarDjLGZSP0qlq3SZpOE74dFlxy1t9BLbvtJGtYyzNtiFzyr7C/q6ie5fQIg2t
pYariOPEpQ4e6AtstFT6gjP0gW+DTYStZsZdktNI1iRYVr8wBYRsAoxIojMdMubQ
fPOFsTkLr9Nn+UWHaV+i/SXRgT0eaUG/15n79nsHkjF6+DvhDQNEJTMHj0TNIJqy
OxeYk7dxtGBKw03pBZb/ZkEYP4noPlAG0ihbmzS+zxbBil2Wg20Tr/os/pMa8GMb
th99VV9VIjJCLkD8EeIKxSyw905XUntzfoUG34IM8JNlUOUNqqaHl/qovgeCPM6L
GnrLDjG8Nf+Cirq/vr6AeigmZSAZ5NgEtLtDVkd85FiEN1NSH9wKRvgzRPbWaRXV
UFMomLQ+7ggYjW5rUXj79kOV0Nt84azvOrEf1WZtirY+vpQ3AF22AmEU65bqMZsu
XNBlJk2fXvw3k6tRmXrHVsSkPvFMPUuTEYbsV8SwOcsgvv2DaDpqjg7ZyR+jwgAf
5Arz0e2YCOMmpCmvMMdWVxyYM8/ceV2kOUYoa8KMkO8OxuIiIibmJGnj+MdXuiOQ
OsxN7oKjBZIrijfDNNouHpWMcmKQR8kEM5jyfF4GAlj+3k1fBTeiKrtdYJwsJqYq
kBniA1dEhG4Q5E6JyE652hhxs1JO1J46vtGmd5e6qhCZgYRTAzw7EQ8IEv67VFQK
Ayr9SBZ9U6f1ghcR+fD4mOrfaZt8EIcJPwXd/THUO/QuWK/uowJjVcTRcTXHbpnL
aH6KRZmciaxZowAkLMC+WMenWcyG630/Gc1YYAQr6GJpcgc/nKJNljQIU9HZPMGe
S50I1T6T1nhQEAeIS/84Z8RrvocXcAqYOF2/xyDe+Si65L2STzDGaDTYoqE/JrG/
R/hdLfoEik4/wY+jaP+eZOaNk1epkCZNd+J5WpQYzq4sDoSswWo/Vgv7ws1nuaO5
L2Svu3LU0yiSpYWKwx2U4jYjDZDM9cY4AkZPNe89T34rIwVcgcRKzBZ64NfLBHNA
zxq7puQN+kJR0n5wXp90gbAMhK1qwy7Uwke5YPnZ8tpWtFdmTbPN8UiOmXkZY354
Nsjbba1wYbPFe+F2EAgsEQbsWkkbS2jpgfY+d+OZSfNzO5V9MLWL/h/e3eTkJA2Y
OeHt/k5BLuEt7dBhNVr7jMyu6hpSHI5R5Wpl2RBi69fUEpHWSxMU9DlHQEofWqsP
dWKN/+QMzZkyYWL9NpS0vqNiWl4CTOBQoHDTiNeAD3EneImBKai8XOQvaRbRyEEc
O4ZOKi4czSEY2jTmYSbTNNsvWaXss4G9oS186+EAEihU5Z2ZKhb+7x9wHSGNHF+U
fmFmNIYYg1Q1ILVBUoa6TJsg9ziVfJErpFI4c9wT1rXb1SmETmbjfGm/400otfWB
EzTIMRLKCPyHb2QCCX3YTwmCYxC1ZkWyCv4O7n6eS4AdWz06eLkuKe1e680EcKrO
ZhlFE3s3b3fynFerc3cqpDiYcsdRaYsoAiOZayRNssolgdfkj0HbzeHEugM8n9Pf
vXJySbhmMMzSa5WnHgVZubzVihdT4W8HnxQabPEonmJkW5Rcj11IdyN8HKM4xX/5
+kIh6GnCptfe1p8jmzczn2v7QmpI1bZbPyECL3WLGOoaT2/SR/FjpJvEVMgnW7TY
Lth09Kzl7P6lA5cdBfW/awm6PIpIdm43Mbhlc+hheKdDpfzilqfJD97Lr1I/rlED
rqxteV55o8KokPws8MWjJ5JqNn1KyNe2lapS6UBCxKAi8As8sWvmvOjlC5wPcYQB
EPL5UXahe1NbzeiAnl11IxzNKMqcJe9/jTdl8NFCbLpcaxwf0ezX0pUU3pvks5iA
oKuhPFFq1uiLcoEkz2Zw23LnY2aQy0jB469oUdIRLuJ4Ym2nM8zrPl3DQ+YroXCc
Nz9HBP5bYJDeG+eoWUwkRadCwQDwe1m2toMc1hBurP66KfctSJeEbCFhoaxMM0Er
dPZCT/Z4hliHjN1tK4JJWOHi6LT2+XoVEMkk5PhaGPmFK1zZ0nawXUo5+RW9grlT
flJrIeENpWEf+gonM1jxEbNq3EAQnKhFPlhrH7luZZge9LcKDNVPoDVWrIjKS/Fc
D/YsIFIz7sZlIY8/DP8JBhhNmufVZ/ie3Zk0FxXEYfwB/KmgWQ8GcoTu89AzG1m4
1wHYCxvVsxgfERlp87+2F0YL2lyelkp0iGnTiG02sTuzXAgTu7JG9KmhhaHdRAc0
Y91YkKH/SzUqbEOZL/tu+a2KrKSrst0aruOoWg0Uo0s22e/chUp9aRY24MKLuxrR
JvPUfUmss30s1TrY/I4GCtDQqg6Ea+yWnCjMLlNZgCEIax85JxfxVon7MOlavN9X
qcrH8YW7Z1qxQM9e8pFmm3+1iZ2Jkmnioose5q8wB3BNVeTLR9BA5mA5WmcyO5WW
DetZzcbZjnqsN3f0CHwx3OYrj+Ii7KPXO1vifAuRlqGAxgNuCJJRAJo5BJvgZrcE
O+hkPPklyhYDQ+4oncbWjEtOf7MM3QXJ2P3qiIkZrYZ1v/4k4At1XNtas+iGdezO
q38nWL6mPoxukM/W1Eef0Dhqrb2loBaG21xrrNlCmDL7/g97nqWuMyFttIgn9IEL
9oHc5+U0K5qiQS8JiJfAHX8+CaW0QdkElQIM/IEeMjkK+r4bXgZ4B46jaCuWF5Ao
c2hAZaIlzg4XTo9p8qk6cKAi55I/kT88Kb4XQWFETie0w3ckyroMGHs66kIIoHjn
XaqWbG77gtFeWLLfn4rkoqe5ZHtAyEYwUFyoBSRI7rAyaf5CajZNzr+FR48vXWs3
HqBblsjwfJRACrey7mF9Q9Ah5HZXVRZq4x9Mk8OgAL1uFB4PXGpyvoGD6jTRPt4d
D3iPbnsfv0bVAbZNtPgs7X4ivG1e2Q5p2bAleE0wr6Mog9i40d4YZKlWXbAc+uUd
uIOzKc36PjQiwUPeP2D+QYz3h3mJuk35H62Q8Hv+vBCqsVGqwGSkJuxC3HuSWx9W
H+mcv84EcDiISw5t1UgwNd3vwO3SVt0dVOfBimLeC7/eKiNsRe9Yawv5FyybgL1X
MnKDWbhuhHtx9ex8HIpAR1QQkCrqCJFCJi3lWgpUx22Shkrpdx4PHqoaaNcvs2Qq
XqnxNk/qgnJ7rw4Xnr7k+qgCtr6lNVyj1162BLCKKFhrUP3Dn1Ist8oBq2/Pfxe9
6X0Xzk+emuDL2HA3CguLIR+UMpf5lya/ECA/bQ2vsmJY+/rswQqBhPYSUdAtvF2g
vdvlVSnTNmfAImETkOyuMLLa0OHkALYMUz9EUceXMVhQHEmq/I8zrQcndhuvAz1v
TtpXvuBqu/e+GungJCfaDadAcOZz3OBZ2Jf6to4vymoOJGX/dbPiz3nZ4XvuFTxZ
E2oHBQPUs/gTStxa0QZVorQMDk38FNwxsGX9P05LCSzK1wsBD2UHep1K8tttgpPV
acUDeIaCvTBGuHBN+jVP/2EUmtEYNP7x3FvrvPQ5dW4+1tvNWpHUZKxOwEbBN9bT
1UAqzwp9BEvvKtgdwjgBzIU+oYDY14J5a4shNWfX8oR17lHHLwlrJYyVNLny93nh
gQOTi3putK5CEga6z9h0AM48wPqXSNCCc0SbO9UKnr1M8JhNPiivLzicL3kCc7qc
JE9I1JWpAL1Zf1HNxnR//oDJIW9cWZzTqWv9JR4LVEOlNnA5Iv6EwG7ODqKJNjLk
CBAhVGCsR21TVWsNjVBGq+/iS+iZ8k9tX9uVjul13AHNa5kFDwyuYObPXxOGEm2+
F9xTZmDxZocYa8+gqvG8NqX0bmFa/GsDpf3eBX60NARNo/gns+bmSkOWOpfC+j1L
MNZda3Bi4f+5toh+EC1dZGWMEdhH7J6mWco5Y2YbgOrGbcIvBj1d+3WpUPv89Xhq
pHgCdbseR2VG79zZp5bfwPp/mWL7P6C6UtfI2qUk52LH6gK2xsBg4FFlIGVQo1Xm
o7FVPn/4SpUIrwBwT1k/oMWovnFkMMKUPnfJ/aZbXAmuZkt1Vdqo2ywLZq+FBZnG
k/xkoMa+2R2IIYwSODaEhgdhLhz7tYrZWbDqQpNgjmUvYV0zZpO+glJpL5LHnqqz
vxAJEt9tJSvVdWGzGLOjC1U4cOpoM7CIMDOyDvlDRK+oT+yOgyHzZ6SI1YmUSxLe
Cvauoy5ifMkao0a4/U1WXc/xaUTavGZMNDfe7uhu4cxA6RBHJ71z57vIr+Zh0W6f
ybG4N4JlvnoO4VGukvgp7HG43Z5vsM1LqM6iBPJGx/EjLqKVCNyTR+etGWa79Wib
VxqxwvGN4ZXtfRbbcFy/tn8D+fnxDotE9SA38pX/8tP3qRKr8YkMNbW5GKtGoZnb
htftpocIwi0T+pantXJPV0VKiCFQnXnQ6ZL0pFhqOuTSWRgy6S4NtpKY1vNwYIc0
THsvMYHT8WBziL4BDl/0+6yK8UZi4ezGSekhWwbVAOqwm6LNr/W/eMVfS0l0ahyq
rNkWs/FS//9XqN6nz8jDF1vmhnKa758rOIlKtzDLnie+B2vNQ80+wRcK+bXdLzob
mv52odtwrTS1s1TfAUBYkt+67KF6CO4xys6Kp50dTLYvaEU/f2A+S7cWyhHggACy
kjF4aq7CBEfNslSq+97RsqPV8rU0MtqBIWRAVBlCtd18D2KnyWeVJ0q01aH634S9
uypk4nTwjqm1mRPcb5/oMdDcyw6HwZ1LPrydicpmUJ9dBfnB83m3RMxN500jMtGU
KuktPFTefe1vSe4NPyMT7X5XrlbeuYcboleKCnS4MP42/BEDvc+y47hO5FrWCSXT
wiaJVmvBiHaw1jzf0z8NCm3MN1P2A6VyCaZ8twBTr8daG0ZgW6FnE7Rm1MVdMbi0
M+VenKZiKaYaCZkURx+cYBSvrdx8Tkqm7zsP9bgEJMSlXfzHlwxrh8adlgftO4tn
46WmIUGpb7gJVNzaXekkBZlSLEuPKLwiUBS5DK9scC9nE35c7KsKtOWDM8hjMMM+
x7ZQtRGSO4bxE41P/eJEXB3ZN4UC9O0Dw2hsQkdY64QWb8h5c+54jwRCkPWuR5w1
uNKG1Vr6Vvt6/iqLCcEHiVMXqjixQmCBTTI2FjXYV5MhbCX94u/ZYpyDn2I5fMJc
T4nn9gcwFDP/xhSTiXbUCyJUkbFknReO/RXVly4HsDjQUviHohO/G0jf05OLEWul
zjSnRxdjGdXO76nwF6Iu0VciC+FG5pYXkEjOvlVjEXl3/abuyvHRy3GBsfR89tCe
ikV1B6LDHtr7wVTiLsB2fo8pzvSDVa08K6/O3j91iCt+4O11Y8uLXUqPU++myabV
bXnWaj8y2I0tHu0GbHCoCVmnXzZVHs/ZKgXoQvE763lSwbJlN41W4zP7Lwbj6oLs
55hiNxnoz7hSqUMTj9ZsVZjO6uzRgo7JXSr88DkuyrBW6qGpgs/eCA2CcqI9GZUF
4Nah2E7aEpw3icR7zxAycx7lXs0fLVgXy9CulODmxuJ0ZVgIDrAd8b17C+esLlhE
9nuPvU9zAvg5CNtJtHa09Z0KAWkjZI1cW/rMKzKWGa80kXpJSkGjtlGFDTZyADZM
IxdHMxz8Lp42dnri8D8IO/N34rUvRaZ82GLBH0eZHy+Vzp5R91tB0GhUwodQKnQT
53J4YcEG5nn2LmZa03zt+u/3zHG+mIHZQo0/2eujJHt4pp6oIZAbPBfUtWEfpXOU
4vjqh0FnrrME75YbBmGMYd92bjZ2fcSr98QN5JC5rU8y/bFW3qAVB/5t8jxNHyz0
ehez1y4IkQCCeLmuUWpQQFuLuZzdSa9xoEG7USzws+ou9ctaxVkFCOrFn+fgMfVB
OQdRcrRFa1+w2dBJtAclvGOOy8SyBoocg6JV0CVb+5vXDCsX1Cignv8NXnzrTFDt
DNgy6nL2Y6grihshIDIzOX/w2+b44E4ybHMHY4nHA6vepcb47fShbWywFwAv35me
K5VBXS3VvMdw7v/0wmb6VpzwMJZASUSlgG0IJDctvHeFFu307N8hbN0O9TtpgqVI
dswG0rAcm5CY/ggG507f33J5C82s+MmUdKWrvB0N6hJGyLIQv8KpVoDPVfOgpnO9
+I2VR5bfmfTrb5WxGxrORhxcFvgneXEzsJSvNXPzcHXA52WT1zNsBDRgYp9VvPmb
FHeK3KRvXHX5tjeba6yqJmXRolPsPGULmUlhaKTRdUjGtmw6HTRIH8bQpztzsAAR
/lESdqFtoMIC0xFCVl0RQHuaRJlGtI7+YzAACNCvz8bQc74AMZeCne4ycx5JYRoS
VgdUt+Jge1VG+10lB3z8J1s4XIyC7ILXHL/ofZd3XRVZpK9xjxQN9Re6gTGHPuWs
/ojgpSThkUDQE/b+x/vSptZ2ugLO6cTW5Fd0SpKfFG2dNvvSIaGIiMiyG400q+oG
Lh92D2sWMTzDXWnJTJGBP/OZfmKLEtR4ERVxMnL+YUOWfdbOak0aBza2UnfTtDQI
4/mA78zKHgY6AboeBqyY0CkW0io1+RPto6KYUX3Q2CRn3kuAYpYJSJiPi3TqoSXZ
SSUK7QBFAgEaTgtrpSM+nJUHOwfPdUu3yxOHrYAomp9xRNtP6bEObdR1wM5vFY0Z
hsP48tltpH0g98oCfO0s8k7bk61z8KMHVvDcC+vE/+6St5HIC0dTuROmMG5QPzJX
zVN2PUTMzDmR/PhqZA2VsohafPeYJ2wnpMkLmVxVd+ZsfSw6ZoGSLWhUxlHbzxPQ
wNgPov79M8IJa7FVQH2yxNnlXLC6gqhm3pdUHVb7bp3B6Io1sq0/KwhtQBD3PMBx
TcaM7NfcmZpkgRfXjM8mOQz75mdGMrG1kgaw5X+t4itm0/6395NnMe0S0BmuHCeF
QKNPwQptvXFAoHh4dvDy6Sjxxy3tzsHUy9Hx/JL4ZkVAkEpXijRtBuP3bgcRLPyV
n89soLiuPSr+P+xhPkVnmH5p/YGUjvJAcUyRro0OKo3PR6Pcz09sQFMij3b6WJP8
PGaeKco9l7KBtLU2U8AS1OzKZbFd4fSZ75oMLhsMVP1WmuXUCNfwIrD9qVJhcHtL
QiuySllR1Vc59/kEY0f7xrJvWElV4i/i6XPS4lGgAf8euHg8BYEIPJ0aMCIUK2CZ
mpTS6bAy8r9nkA9RK4uRhvDG23FBnUZQDI9as/aPZpxST8XWF9kCgeNAAPuvu18A
O5aepiNDZUsXTW9M+wFzG6dOndkg8a3r3uwE1coP/1zcYnVAdya/02nRT6LZ3A1c
+CF/kkVZ86auELvvaGfcwFPYLa7vahqQ6ELTKq03W4zY/OJR3MKhouJ2oXusro1O
7E4nIdKxPw8F91dpTSq4pHazuNqLSM2P7X7CO3R78tG+bL4eyzcoHkmRuNtbTIiE
vYYufazfXhMSwriq1n0DN3BK29Aa4luUOC0ciqZjAV0Mkh46TctCAB8NfFpBzi2O
O3EiErtKkfFa01D++5b3H++ptMjON0bFXKcGGRnlz++h+mS7w39PAPm54tNaF9AW
h9lB0gx9DxJQO4g7Q1+2CVRtk+SPuX0F3vFOCNHuKzcfaNDKFwCEbSiWIbhzYGZP
pF0MXr8J+IHEGz8vJv94339we0criw+HSZ63jfmmgoKEtmyM21LD9DkLtYEvj6b4
OhcnzsV3Nd5BVaa5CqwpIckKdPKSnc3qrsgZaEGa+6e2B3GpgpsNEo5gUWrt8rKY
3WHEmC8GcHp2E8wl3QfiaFqUy5Pzjvpf2PtlElaezJSt8f7yLL1seSl/p9lBxFGQ
IJlYkj+P+giDjzc9n/1bxktOqZzTmjk+KtYmZLYu4LvDtZgOegAESWUFVBtcqzE/
GLgDsCdzac7I2NYAXdKzN/eg4zEq1g9oCoqLSYv7dSFvB8SbcFu0F83VY0kr28Z9
tPY2XSfSsjKD33EtqGbl+3HeZyJGwlZhODEY3hQPWj/39jfa/yYUgckkJwXlGfgn
inblRxk/YAlS21qs5tspye+b/MKuaG0p2QdF+5Al6i52JapAMiJM0pXd2wt4Nreu
8LtjmunIniZLXcWFWeuKFwraAjcOjLt/YfODjrreE/nerFjF29fa4x2qejD1AR0L
ORVg7SDjmEMMg4mUwKxx1GHNJNuAKBczIQpY9FlRFjH+Qhgv9QsPNOYpuiRr4mtd
UHbNqOqEoVsr05t/7p7h+MyZXceLYXAwWNFVNEVUD7fZfidYph57kGO9Yk6I9aDv
Bjey8C70oj02shxcMzSe0Uo8m5g8q0EKehFlbpu6u/0i2H64EeWs/IwkdpLrQVzS
kvakg9ahwxAW3KN52WruNiDCcos7WlyrfQuoVpEZpnimxhyR8U0ctwvuJfPM37mZ
wBc6cQiyMp80Mu00ddacDkiCJX5/elo91ehwDIVVuJaKY+ax+k5SmotV4OwQhQbO
cCsiPrm/pMjVw5S9CH7XqCl9Updlk1UjLg57YVWdcsFTJvg9XzQ3MC2CCMq5V3d9
1S1IEjEf46fI3cco1MYpUtvbUUF3MT0Lyw4/USei8u7PgYwE7KhyORdAk9XJ4dnp
vA69duDp0svAmSnHAU1EZ2ivHijmm2UZlR1MMvc1BS971MPwebXwuOxasdP/yChx
lAPrFQPQItLpo6eFveWpeEAiyWeaEPYaFLc4EdMLeuOPZ1W2Go9UESwsOcHQ8LmQ
H0jhnUh4OZhPG80VL82P4wJyyyzUBq41SgooB1QX82Jk3KOaidb8bsLNLiHbRm/t
5PcpnK64jIAB4SCW22cxamM/dk2ERFQv5HUbhZCfR1QPyD8q+K9kQRZb+oH1MRv0
iR140H6sUfU6JRQz4iopIzn7eN467ZGZiMaMlBpmewS0OI+3GkWSNQm8nCsnFyu2
8IbrkB+2uiQ61SsEaRF2eIFX6EnAdIrzIKEg4KZXHJvK4Fow+RQsdcusgBcngX/p
w2517u/x46LrK6sBiF9A4/YAtXuz0pX7FEKliqSuVO30UjMqLuArajAWb7poZFBW
/RNWbNRFGxt4i0wr8/peJPl/PnlpL9jwV7urTVekxNAVMlhz3EhvigEa6NC6LGaQ
CNVUpzcWF53CgVTcOOLwJcXynWhrsWE6HbSQSHAcN9AUNv9QDXMNVNf1Dax0OPgR
Lbt/RU8nzpnT111wVER773GO95sg0NHzlCLib+ux8urbIWR7lkBu4nBGPHVmyILd
cvvv0Eo1T+/nEHYddaW8fA7Q073XT8UDrJn0uDv4mLyqBfLYdwHZsB/nHzFzXvfh
5Quab63ZJ/NZrgRtQKcttm8CmMNgrSS16N9hfj9c0AyR1K/yaa8afkoZw9Ahxo7s
qC/s9HMzn0jKGcVV4IBLcDl3r4mMmx8SQzutRPwpqyi/z1KcMk8dPNXDVmCkseYp
gOQbwLEGFO6IG9+4xuFsUdiziauaBTzijIvGYrEjnpsMZzuN+l30xg2PvOP8zxI0
h0AbciN0m2pUGVhrmr7nJDDv42FVCtIoiExJGOZsQRYQZ17i70x4RrFnMbl4/n9G
k1CCxkdA6ujtXe0YmX63BgBMshOsuf7xZPFoZn393ykGI3kShXM5hX5UaAl9/59D
MXhS/DtHQIeNTGIeDFm16UBnHiEhdsF/2mIGn4hR6q9wFH/YdRUaPAW/aQ1MfQCt
TMoodL0a/gaI2bX7JS93/uV5PeCZDo54icnVUMcyayi8C9LktlP4O3a+JPPE6VM9
TfmyuLrQhLYenXU1UdIfLq7CkZ028rlQ9rafu33hCWwHWDbUMfT7CjuPtfbL4FJQ
IscD6ZW/Inx5vWoJQnBPF0xXoKfcosvT7Hp7y4r9HqmorNMGAMuMFhbhEiy20npv
W3SBX/ivUaFAGa3EdCTCkOJOXy2bzwoq45NIXZsJESreqoSudFKbBOSb6ZYYcNic
5czUjhsrwSUy3mz+/UdOLvfS4/q6PQjin4abiaWcqesIKmEqBZAYJzqMxQdCuUu8
mb3rMSDDo7zrAp5b/L7zwqXaoxszhGz+Z9OQKEpmUMjt4YUgkf3HNb1wUx9NiXuD
AoYn6NAGjY7YFJnKKUH6lrn1XRL19PmGa2eCXA/FVzZxRaxvY5Ya9CHIZfWREhZP
jFmJc0rxJlTk58FST3XYXA/x27iQVEviIajxaMs86AgY9QYmaIrrD8AqRVSgPQIk
Jd+c4tbBP2K1E6DtlqvHDyO5DvxhJYi1Slchy6HvdRkz8/ieWiZ29wK6thrkEIhG
RBpLIQKbTchiID6Xdqve1vsxpjuMQfr/F8EsG5SkSpWft8n+6zwOQxNRan+FsUBQ
JPAZpl3kDkCzN3H5qwVj/Jlu/Zp6UtDKLwGBA/gZA9+yJzDtGM/SWy/lewCJH7eR
lAVIjFWz9ep1cbb/BqPeUAy39INO5fswVuewD4A4dg3iEp7RKGSRiFdGiXT0olMl
S3fFoRMVU2dVg+hoczlprf7G/tbhDbSJIlHpit4EX5Y45CKO6eDL70OK34SfczT9
Jh/+Kc4LT/FIwxUlkrccBC5ZYGI24HL8TwkWjUeyV1SL7eFZIb2EWlBj3+fZE0G7
R125bmGqgnlVI/FS7Jzs9OCzrcuD6M2vry6ocExeFMPDX9yg5iEbr4p5mSkoK+NX
CdpU49Z1CDmwSMLhbQV2GW7yt6iO/CjWAKe6OCLFO/Jx6ZrfrfrNC7mtAzolElH5
tIQkOp2eySpRL9RAX/7zR5ugjmt8nrx3TA+NAWKhN2qz/Tx5k+e/F9H4u8yuAW7M
wL53YdXynkZ5f+HTA5fOgj35QIFNgxEvQl5MSvhopGXO9PYuYo0se/LP9i5m/jF1
U9OQawmuOj5DQLmyQ0DnBVs4qS/SADIbP60hUWjXCoL1D4xeTTWZLn5nH00HNfZi
X5D57ZLaVT1X3Z61YRtnHKTCBnfSVg+BLvSQQIFeeask/oqXR1nXDK7iUg7c0X7w
+YSDflVSD/INBp9KD16HZhqfn3fMG/RIGzKfFIYsgMRO+sQSGZ9QCDgqjcGu9iNS
W6sf1pB0DTtAZOecl6TD3ei8R225nkg5KgOHd0eSG7l6dzuzpPjvDYuAV5xx66ET
PFMG09/laRJ5iqBHP7ZcW5S1sGyELoYF9bKtW08VhOe+LFQpZFXwcyyR5rpAMMQn
2NGYzGMhVSj7zUYsYLFgFag0Ame9Y8oPIhWDaQsvCeGtqEaZBnPVp0NIkH0+Y33A
HnRF5Bs7jXrvSwq+j3iBNUzMI5kXkSosiKB8F9QEJgOBGjvmP2OBEBM0xpUP+5ye
5U4qEelT2GtFfI2T8u3S7R7EA3b9aj8Jut8Ko/4v8YreoqS0jsCOntfVM0OcK1hB
r9hcqt149pNhkHw0uOOtQnFLvKUSrAZ1vxxirZPkM5h8/VUvPgmC+mkSBIpqu1N1
SnqMxjjJ28CzdvBkXBZ+0xOfBLg2OUGl0QBDhxWfnmJeAU2Tup7YuTzIjBpMxa0F
/PheB4NLz8+wajQVMSx3Il0o7rTSVOsAXvla5mJerK/Ae7uZwSY2wxeZG9gXOOn9
iuGvLrhvQvZGPL+DTYht0OFPhkPEjElMmryusYfTP7/+th+kXjnrCZ3BUmgOG9rM
pT8sFTS+WcKvKfv6nVzm6XZPdGC4lkgwtyxRfD0H1d8s8iagCBygwzAer5DTpChx
0Zp9tT5az8o6GvoUB7t1OZk1dU0gcLSPR1wVQhsDUDCfMLZJW0DvUFvqQy9oT+/h
K4EO1w2WAA4YV91q08i4r2fdxvEu2Q54J2wfG2njlJEjZcopnxycWXqHMSjuh4Wh
tH6LBeIulaqHWNwkeog1cyTdIf70QVGGXjdVwnW/xiQwjhV32YFusP4ADsYSPddA
Tv92S8178ik5/rCULAzBUZTtRlMuLk7A/NAT9VEzXru4+kHwwyaUAct17AKVRQd4
2PMtHFQn4KymvDZcUhXeb8S7X5i75L/La48VOK/ihirrb2tMKjcAKPAPP6ASY+DB
qsQ7b9Hfa0JsFoV5eSpPJ11mBhOoeXubIKhu2KKPakSIHeAWgrekfm48nehC0/hc
E8d8arVEx9rrQ5cze2yHrNYNRAE/hMpmcPkKwOCRlWDTsR26W90wdttV+AbtlXYZ
+nOdG6ybCOpZS5PVoknn8WCJkfeez5YEBdk9+eWW31t3nxGX47/s3Ty2pIiuEpp1
21V9zbqraogGl30bUhGEKvRCFmfE7xmY9BY5I4NL5E0JZ/oaU2bAnSxpwVC24epD
CQA+E7C56m9LiOls2B20IpBGih7a9iL5um6S/IIoa5geGil15EapYZ4zmpv5iDsD
uA+yoKv/LaHsZRjP7v++hcBTkHiUfhpjpd6yEcKUf2r1IMjDgiOxEnBpnpQXJIxm
jb3ZEu6kP0qaGkChLjtevEqOAp7oxNA9eJwJw1Gf/DOW1MzWJ3o6mBc7j+b3rnmP
AnIlQaRD946pMqnOBsGULfLFDhclDO+3fSoDVL61oz5KSj0WKDNnRAuyfDquOUut
BCyqkIM3jMowG4kfhw4kss/MOb2z/peRBz9fTOsS8VFSTTpmYagOUpRdOaFAe0G/
XH0uhv1/+JgpR7ZCBrjgnb+oq/apWxtxN4Cj3HsBHg9tdb23/sO0uJoZYrvdtwKj
M91x6/NPnE1JnrhZgyoLgOjCFm5K3zo4Us4jUSainXrfOtDwnrce/AE1sJX5hvWi
6HDEpSb+9cNwk75Cb5Wpgc9i1y/9GEATsNjqUFn8JH9OqFpaPqdO2zCT2I8SYvNY
uW5keIZPbTHmeKNHaeto78i2YjUmFyk3U3zWikGomtmxdv49PSKPtusb6+lXi8nL
hzIZ1563k1IvcS5Ymyy+ZWBwlk/yKLNWbKoIrwi8nELR5kR1Hn53HNdHoTq5AiVR
YfH9wEd/Pp0nG/PnEQWVR3FfhFl8zklrbV4Ro0GQfFN7T26UEP531iZ7Yj+VJayk
X9fzTqD/STl1aiLf9F5Id2+TLD6fXGhTtuB4JoTNrtJ01YszW/6HLTbQ9z2tslKo
vs5cv4ZZ9vOTUslHws6DcyJ+HycMg4YYXGPKuuShqovfsmH11gpuqocjjGmQDCOq
+wjHpzyc/PtkCrX6Ntf+942/QLQWWf+faXOsO1e7cfOR15/Zd6xmhzY3YU7WwKr0
oXJKpohqSEptrMRyzsEVnccm6ojmFGy2BPg7e05wIY32Tf/K/wSVVZwDbf5GGRrg
sC29JVBLcN1Zwqmh5VhX56VZrprQRK/S4odzIFb3X6CKub+OWtVccAZUUpslgn/2
Q+U2vleV5N8lxVQ55CWYL03jvEPioMo8U68FH2Ym9olf1e5r45c2AOcy3E5xA1jA
p4QCdsYVU629mB5MIYGlzXy6h8agTKPwIZmt9qduPIhcjovI+nw3cSXnoRKg7wJ5
8JXXm1NrYj1vwFxYogjd6bka1PCB70jVV7NriEXXG7nt8nclguAASO/kryrj4IYW
E3x5bA5P7h4z7pUkLXSJSp0wsdpvC3cosnTRfo+XYtVfdovR2C7/vw5EoE0mML3N
LbkmQoE9vyVXx0EPYg6+mRISfMkMHjMhi8VF/ofwOv3tzx61kfkx4ovSrrovVSvC
5mC4bMY9B3ALzQYa6L5tduzdSm9xltpqvZG+bPhRiFyo73I5FQyTkSlo+0JNz1WH
8LcRpxLqeR7/nDcNjQspHYh04H8LK4KYEFERfY3pjqvsoFtr/10sbFCg+5iDU8BQ
MtK81vNSlFGxbFul6tsUv5+ULhwInHncDBj6+KfhKL/ogXY4pgNWF4TfIh7sKW/I
vnR4dyTLthbQhMw48KLKxSynh1XcmknOtBv20s1wzNkWacbfr8kqTr6z06viu1QT
cDDwmAMjYl3FzlbIutFGgUS5waWkXPScUFHsmzqn0p3KvesdrG8Z8j+qPG+IIRrA
QR2GWFNvPGaNgV9LHIdMDKoa8Rm23sI0QJDKQA98mdApTR1BElW8TkeVw1lWL0XA
AMj12Oad1frJfHrSs3BafqPUi+kbJJG6RJje2EqNxsI9/hJrXH9zd0pUhNWq8vyd
HyODm3V46BA/PVrOYAVx6pgchbhnQLBbnyp4vYS5W0R2RQtxdWTH5JaCAUDfIxQK
16IpL432DPHiDUw3daeGxkS6IOO1Xuax99NoLMwnHlf0uzba+opJfZp5j9cb+KXi
f2VzM27MKipqJdGrJnDAsGW+D2yoL/LDAyCupki1Th0dj+K9uUZS9ijSSeBbNR+9
Z1898CEcBnjiXcBRp4tUfr5cdDH4kY5mpievt4U5lv31qA5slVHwMat5j6pncyc+
c9XhRTECNFi0CvQTaa3x4WXnGQ1oV9N0j4L5IX9yCg3RvsroVDhSTY3kax9CnsO5
jrXRIqPBeQymDYc0j590qofgLyZtMldohMMxiZh1103jYUqME/tCAvNpKlUIPuhy
XEXXV99FgUAA6PhDKlGrGg6VS4aCZzbdDwlcWPEJgJJ5Qg94GguuqSxfl3wwEHbi
YOMGqD8snfE5HCeXAEKe/qG7icCm0OAzWReT0+mgvOcJYVy5yKDK3QN09X5rACHA
lLaGpZo5m4s2XJc333VMTMUxwcMh+CAmkJzk76DV4FodbFJApw9tVCWPNlvlGd09
POH1FexGocSoj8rAPdNY+upFnxkhp2RJ0pbvk7HttHejf9Uz4eyf/KjnACUqy5nA
sILPqK109EoHPkutXjacbAag8b/kv6Klc1vfWEnet1A5j91p06D45RG4k/pHZiZe
mEiUBleaTHv7Il8pY2q22R7V0bDWhLTQjIuX75TqH/J/ehBqAMVyHLye+jFuZ3P5
fLizZwzpPSJBtkpK2bhHQMWiAXyWaMVQrF0THZK880+vw6xTg7Gvg93OR9jWcf/8
b+yNy/cc6pb+0jdX+weGG8HGduRTa+qIBLYQ0oFVs8O3H7NpRfUzZqSmiHI9oGB7
MCJ/0yZ3yy+YEXzD6RoSLTmhUDoNKzuqFINVIoXvfD49m7no0/bMBpiGSspujUWg
9cJUQdmgQpFc3N8sg+AnsPiRbgmiTQ1jV2auLdHjjRNKrWXqwZ3zmbetFpBRNF21
PFHqUa9WHs9XHJP0gJL58vuPkwFVpv1PKZUEYWJIiDa/L2+ylMEr3Ciac1/+EIAm
O2p6r5TsxRN6i3f79PVb9fle23jzP9tB8rbIy/CMm+zUQgA/HRdOE8wbPSjWZlx8
WX56AM52D0/mnV4Vbp/ebMxAsRuTNIN9B3rEPSFwvDmXd8oZ8PFaDqHf7L3Z2Skt
TLDysgOnUhh3G2XzZGhwGVfxnDgT5l1g2TYlCxf+WrbgIbbf8LviZsn34F9eBq1a
z7iWzQXUnb8sJyZ8xrcgsEOqK+pZotv+1KWqA7UH3+unVLTYMSzROvpp2khgBXF/
/rw1jAwPmp8kVYuO2j5woYm1ixrLiV6nxGnJ+kKNHS4/9vCAUFzoL6oTkMGOqEdi
xIwb/SIyYH2VvYG27kNWP/2UiR0u+RCIy60Z/mkjFI2gnToppmBkRdWM5SV12J3r
3lJ29kh3SwYYUaGRQ3NQR+TrSNwpbhiynTzaaAA6V9wubzMVHs2a9KLSWOURnHoK
7/Ybt9aVC4+Nmx1e4DmlemBSGMst+i1ELAGYuMw4iFF+7RMZlxABlB7Vxr7420B1
Jv6xyW/C17pOEuJpsQGyMDbjaYq25GtRCr2g9Ab38MpagvjZQ8O54mP/evjMjCbD
ADEnFBzI7Hb0pUTuEHUYc5sFudyABa1lQJTFwLwTGNn2GKW+TkwEh7icxt6O1Nve
/lOLG+vuXDtsFYYgrL37Fu/OI5wxL8hg6KoB8rbVLQpi6Vot2jUtW7Ow4ZN3jMeB
noYrYuLVdhY63G+QN3mmZapoO6ZRdIwhg9Hv2/miiRtLwDYZZcXuheVhGEskPNiG
hb8SKaWL28H2VyO8NRtUv2nc9Cgg5vkK2Hxes631Nml4OKxQpsegnTiMYNavLZBO
HeKMhUPeLUpnLcwmYX4gOD2ZP5qCsDnZwYuM1GCYJFif6R9Mfcu5W6L7bUdnV3yO
+CYX+aNmUmsORORA1pqoEdYNqY8J3DEYljeGBd9Pylyh2OWzzRgcQ5YuyElmOJ4Q
bH7kl9OVzsscTj4tfaPuYRyJRAX06ZIkv+z5Z/crU2Li8xoviUr6PE0vFcAiOE+4
6UCg/Eki01TSNRUw8uhz/+s/I4U0KA6TTeO/+zgmERen0y5MggD3qTpdRugf4NHs
yS31kZlIw99gWuI5k0eZRQkxyphiemW4UQpwPbApcB2MDO6eZaAuQ3jStheDAAA1
lhfLStYE0bietFhqvY8gN1As/LCwi4F7J5/whoPUPFdrtYc/qmGDMDACMmgYpz1g
fDxolxq5KugYZs+DVZkxi8HJ0TzDT9ax4ahorNrZLtl8MNL1nbZQ976Oc9zR0weJ
PDpk4314gF+5GaAz/IQ0lzxcAoTnmuP0BgASBKvfjqIMRFuXX5lK37cMmtRQMxN3
6DE/0HISALzJ6cUyn5r2gwVnCh3jbnVY6wS3LdBRCbmCQQK4f/4N+8hcVO2x5ao6
K7iET/T0cIR51EzVQBjMrHzuBdA3yNXX0nnKAn3d9MAuvTzsnukIgxAw+XqB5f+B
EhyrZ2TDvYfO2iLvKTgzl0WgQz3sBt5I8FJkMM5PNJ+sg/6YdS7uffi0PM1RLiyw
L10a68EOGSeCfNl9cUQXM9n8q4H0Lt2KLkY27iwz3Xek6LoGmZbjU2tXGFln3sVo
i6CBN++nOAhh27e1vvxu/+oB/JhuwxHgM8X1lLCivtKWKYGrOiXPAmi3Ne3WaDIw
/+EMQ6EZuGs3vPJAqKouLbEqlg55FnfxjKtiW/gX2CWp+U7fKTAzij7siXZMvxqG
Qeb4XpNxvykIRcBps142JDwNeDz2tMBFSanQeEsH5j3P1nocZELJFGf01dz37Z/l
X0MV1NRoNVUNH3QWlFzcn4ZlYMQN9NQwYpKx1Pa43UeriAZHiHnpBaMBiN7czUxG
+Tr10H3fsz435xPBgbDa7dyS9WvJoR5/+fNEo22zudqMp6yd0UrJJWNY5X4P5Qeu
JLkifGSz6avz6i3cNJ24+hbJLpq0lBn3yaBJQOgl9hsuFV3n3kg6GSF4Fu4QYyeE
itYHbAi7Sm2UWXCgkCywW1hoBLTzmTVajuCxD2NDsHDEYIFCrZRNccd3EvTk4Amv
YHpAQVls5FAYIUGViicOuYaYjr3hwfPkevp9+9HJpHHgxQWlTQFZMCGbUUJAOTfC
VnuKNpeVgT5y1tHbqHmmoi+HViO0dfXohaQbTF8GC00Q2OfPgAvBHiWbhrbrXdd7
Cc4besYz6LQJscqJardqlGXghiCJMI8AFXQCA11tCg2njXZ3k3RIMQMJ92465deo
SlZ3WqbGB5qWBippTicuHFD6yhRrhks4sJBOJLZbsxWX1TIJTYDpdT/RDHepYghF
veM2Is2e23yNx1bxOyZsbA0t0IQSfy6TihmTwumN6eJuBA9auQa3CQiAiOOuWAKS
+9xBxQFIOJi9OAJ393icuJq2njSrPeiYL7i7oXAcv7JNugxCuC2AQAII6HmNc6zL
vrZX9vC00Xr+5tACoWwTWhrasjnY8qEGR951CaG8P5J/5zbvhIp/2sCOtUXyL3kz
FlFjwFm6ry8k68fGOc1SOQmyClFSgSx24eI503n/DW02nhpnQD8oU/xja19Acw2V
yhYGUl1G5pTQoWn2ZrJOM473dOPf3pPSencWmydqik7MOptbGwHkY9isOnninQy9
8OVqR6InE2dFLYNtMMZqlRlSK+w0tOG5WJDxMu6cCDr5BcspYch87owdWG2kGDHl
8ePvl+Q4GZ2tq+ePx1gf3jdNWGoqWnxpg6kGLX4uyW+1tXcix/AuOQsX6PwREbj1
mkuxH3G8MHCVe+4cBh32cWyVv1aaIEyRVLzSy+RmsbX8uyfj6mt3yCJo90qvor2O
Xi7tm/Tlj2zBn9Zwqv98hWrdsFU1/s+gzzWzfzTdB8P8zn/EDXonnF9QEd4vRsyI
9MzpGtUhGbtqVTOLJO3bcX753fxh2BXnsgcL69B1E491YoJZ9JIo9PqWL8yBi+6L
XADDvaGUWViXhTE9vZmFREGR73KJ+wh/VjRnMvlttdollYBivC9dMY4kufxS/yyZ
13wE2f1GBI85LWtRCLhE7UaaXwG5G0rO+kn5WLX3xrInb/DNokAQAXavJF14haVd
lpagcs0mB44pBK8A8pW6irPp4aL0InCoI2gxCF6K0C/LxJnU/F5s3nFqRYqxgpJD
dKgkHXyZN5OaEA5Ua3Rq2VV7Q0NjX7uFsxB2lsIjYwrJDhbk1xJ4e+VGl+vgRaNA
TvL/Vp6Kt7NPclJ4gTSkYQxODk+SLdojrLU/MK4DrFCZTXTOADuuUYla1PNWdKad
NsTnKupyohhpFf5i0SdXKCZRp3d3ICCjHiGfH58TbnZ8ZJuSM2bTpqfKXE7xQsIq
KIsbXQl3cUnyDJVvSf4xZ6oM+mFuhATLn0hxSLsvSJX7Sd0P9BEoeQ54wH2mH2d9
AdKNVMX85o2JXXFbF0+/Zb3k0z4/WFUa8BM5jikzu5FqxUFV9bunqlXF+inAin7Z
aesDjlBDwWVb7fDS9/tQz30U2gemB63xloBBaZ4WRpsAQE0ULkjyyrJ/v+3dGGtM
2SgIcFNpinvhP5YizHdP74b+RB44NkOQGoiGo++NZHEPJQreI2l2mvoNAZG5eyJ8
53U2AX1ibnCjPvzDMGG1EtfRXc6x4WggPtn93H5JmfTIAruFeHKMzpaZKn1DJ2DS
PlO5nwej6X08Lgy5eteXjmbqd2YWk1iyqjWtbwvCoMEfbxl3md716P2gjH5jbOA4
Sk02e/xSUoVbo5nKpQ+w1DPIoga5V+3bdZn9G9BBPt+nzoRJzVu219X6irR3jnC0
2dtWdIyl4dmleWL6M2cVP8EM7OMZ9UNTt0qFRpb75wVTwpq9afjOU6n1uje1Rej2
hEcmsEmW6+aO+LNI2/FWzm5gqD7OQcJV8wLb5x+sbR/44zwgSYOKwsVuAmK8NXhM
x5IBfNwX1bSjaUtAycXyThWDFGMtgeB2JHbkwsWOWTb1OdzCRAxRBMuAdKj0cEym
1NwQTxecDVrdT2DVGKLL0N/cqQjEK88H1CILr8Z+Q8GeT0Ar3sB5SSdhvkH//VmL
WuYorfo1bfdf0WsHmofwk+KaZO6tVCPpqMZBsxS7qj3GwunrbB3/iaUdBu68fa0q
211XCIgnlbFTnqS44oiG+1RYSae/oFlwJN+WIiUcG8F7kf2r0CDMgH+kZ18tMSJR
hDPBFyoz8XqewcQFsnEcgg0+FUKMzeHl+i7s0iWsbXh8xNNDBkWiFmaEYpdtaPSz
3R8eDP29ny30UVJeD1lzhlU/tU4tvxCgk06HeMqCrdoxwRm98n2dnuX9WlHmjGxu
ROy0K+IBAvi2B9pH4c0GPEAR3GdAD/MVeu3OBtPN8U4pQCauR5aAR+pRf+1cLzsp
6hBuwTAt9GX3OumNGEezsgqRDMQ6shISoWzzrk/IKA3ZyvAM1WLpqY5bhBMuFZqZ
wGpcwbs3//jK1hzvQKRuZgfWd2oLJM6kI4geOEhOBLYOcqXX6RK3PSMDQSHLWTb/
K1y/UIQ6b4nDHYQyDzUjS+hmerbqln6KMhHqwEph1YwP/PznRa9rf7pbnhR/3Ufc
WNfuQGDbaZwivsu/hnFLMj1+GwyPzsiVUvr6Z2g8y0r9t5XxOVOySCaRY9f67xdD
ssjJNHK9Aw8oZuFIhxAXCEoGlSKuq+ayP/j8EdfATusEohQSFyjoleT4puNcEq6t
LmI3z+G0Y6hY5BTlF6V0A0m2UFlc7ROxaTmQ1kp23mIqdn88WIKCZhTWZ47Ki3Jx
8AVt58Mjwc/gWHZk0GuxQ+Omi1FgYSxxFmhpWXpHM+nV5nkTv4plH9K4lyaplUR3
RwQYppj8oGXC1V3p4K8ccMVwGgQEO7R9ihhB5MzBviuiGnBQRi0Khqmvzjg4gpW1
qame3hCknBNUNYT0b7plFCMlVj3/qENrlBFdBIn7L6SZMxKvl0q8n58fG7w19dRa
YEptzOu0L66Qx/B2wR4AOZWJHyxjytk+Qb3YAjR1I61InkIP7Wn22r9AWoqEMBoA
aJVB8EkOGk+DgLad4G0hq/pLPSrTC3cEjZNFG0bn7k3hxLfoiZjFhHozKcF4Sejn
wR3OjgWrZLmriuf64lHY2YKpLPYcfyF/cE9VojEo0IIWGbckGZhkr8oeRRT0c59N
BRCL8YO0IiNfjKyFBl8EhcePfphtuIysx9YJINjR7UGznME9Ry8DnW1wjjhyYrN/
mIDPF89D2Lhjz0aMu6NdU9ogEzvfZ4w/UZxvPhTJZ18CHGcASlJq8E4SD18TTABU
8+3N+hT23SBLZng6e6mmP3r94zHrqRnMSGKtRDGVXjcHlTKhnr6tp31J+0S1uT19
NV0s+/8H7pR233h6Th2tNNTZmkqI/OdVMYDQ6kU9apgBq1H0lN0S128f5300nWBy
xM50Qvl+eOwnAtgNuQlD468WlUVcEIfQkwC42IEJcum/xVV9CL0SPDg1hVbqKclP
IjtWmvhiVT6tOzZb2ogsyYTGqfYxc1qY7gHorA765Vn6my62tS3+2zliF8gDSEVE
IzrS8Qc52w3c3NCKISmbgmaBZ+DP1rUU0E/+6txkbtDZkozq/SwVjBNEEBFlhP5K
n90NuWF5mJCdLKYuTDSI1M4Lmjhca22cqc6wMxwWH3To/84jydkjMQcxt5vy1t0X
fdf81d+22DtFHXg9X8JPSYq95QASNkyV15iDxXEWJ5+ov40VfcF2LjmukJo6tKPr
O4CLbrQMjodKCEv7PaKT4N3M2+VZUXIp99eZUzexoi+uaGLv2tuhlD0KHg/Cn04x
4bb0yN2Hjy7lGvfrHEU/SaXmA7a1IF56CNPBckLg9QCc3RZj9RpxGPDMABri+xDe
6K4rsbnfwcIlctaWCZTwSyKRtSVu/RjYmVgWW/odk9RdlgVtIv31+Ak6ndCIn0s6
mjKTqd0z3bb15N+Kst4No7453VshdTXYnimi7vcltLqZUFmr56ttre++9HMlKYjI
sIR71CT1xDVLDhDOPK0IifXcHLVyTdTY9qMv34GIpDBqylEPSmLCu0mUVoJ89m7w
mngRRwyhtCKF1KV/AjIJ5+M+pf/Fgmals3HqVZDMGt6rQqy0z6CQf0nceCUR2O+W
IFswjOXmBZIC6BBPbiXVgnvJHEvSgoRR/v08JM3fJ7d98miJGW9JQCfdT2BDDy9I
z3zPRMY9IyLfQ49/zijwKW41OUAC9BdiVC30vFIgNTjkFoT6bB6cro+ZUvme9ihV
+PumcmTx+pP+1FuHvUFWAiNJJb2XVOiAn195Wmk6BRBz8ZLR0Ysl9uB8cTSGmOMO
lJpQWvKDIPy9KD/1T84PVJ05Gk8K76posyH4Yxq6wHBLG4Wkk8Q9fCPPThedSvOI
V/a0rAfGWzlYx3xJMHf2i9ZVvqXWkMGxSdExIYyLG/12dR2G38EX+mcaj2+OJ2cp
WIxfLi2IZqGIcm+heS7LHR/AOHE8dY8Gu8mVvBYt9qO7+v7u94jJ3B5//CpzAo1e
YlqDk3EMQUjEgiuGbC5z/4LAx3oLCl7iX7XxK2GpniYtMUWRrAoi5NnSYcnPu6JG
B9NVxSabDIzP7WYSsPK42hjfwA6U+9lDWH/pAXCWc95wbm50A6PhPL7MvC3PGLDA
Fhamuq+aTTB4OiswMRvE9/XIHm3Evi/Qm9AoVffCwcQ5m5CDAuugzqUQVxSrV2yK
vhKmnMgJPSCkarBawAOPAYermc7GUTtDktmuwOwNGkap4lkJMdwdSs81a9bX7q5v
Z58xGw2R2w1XRGSTtIojX0MGgPIbDklFCVNKV/XKHSgz5b4Mc4HaX4gcYmDjErlm
8EgjcqImMIzIT3uAmyJjs9YqNeFGrVBdRAIRkf9MceZx/Tm6msXzVIqARQp2648P
ucQhtXMpR0/PNV7hqTp1hJeRZGL8mbj1NuBus8O4uDdbbzQlxZ7XYjRkrPwGWmpt
XsfHZbEO5SfRzm2Ha3/Dm9lmzrdeVdIJeDtpnGVnZ01EmYagjCd60yeIZ93nKG3h
ANRDsuLGeeq1KYPG5Wc2jQOalFzspy2oX/8Z2kdZj/J+aftzE0zTZa78evQlAsDf
Sl+oYsf5kw2AeQyio3c1EQ8wlyJSsrDnj/e4vrffsy9LE06rsbrfBTdJsg8fMo5Y
AuDxW1BV4DwKnFO0tc+fZiserWkrSCflGDHHugIhmUPMN0b5zeWOQyOjJUXnIptX
SodtxnJN8id5Yb9NlApgGAXHzkLkjKc5xz59fc1lx4QmXS3Ri2AWWq9nK3hiCgjM
T9RRZNOv8OGsbSOv9wLl4m6MftpPLSYU13iVqDkl3xPfe37dJytCqmUJA8OjnuXs
LDDCbSZ45HyERJ4mZJ8t5iyvYSJOAulkn82okREqm7thDCQKmEZUSkJc1O8k4xiP
w2xjaplOc9h+kzZRrHriJS/DQAhbbe0FKVmSbEOxcwaqmH8n3lZNtjIVlNz9yj+4
A+paOUq44PeStznwWXnt1EchtFx8VE25E0txvx9gXXKWQfmEwqlMqnIHZl9mC4fJ
jDRErfhsOmi6hclqMVYDTn6x0BflIRGUO/BtG4Ri/HG6bj7D1yX8YnRZfIsmD1xw
yOl1KdaR41ifEFTXVEya+cP94Yqed/c5HXQE/qAyjGK5352dP+wQtiPHo8oKqkr9
sA+2Am5PgdP4aadyNwj1g1xgMDgBBcb4VB1wDcefiodl6DDTLi3aLPgdBH928mWs
Sge+xQ8+ooGBEbIxt9g5sq2syUCG+iKsFjKpfMj1nTdYLVEkw0NAF2znH5nDnruK
1V/IqEEAxdAa8KMCTb7bn9hHuwVcts1Ly7iMSe2JbOaoKJle7WPD+lBZHXxBAKkR
3KoPAD6xAzbybMyUwjOx52wWBwDYB9htju57bXysOs6ddRPevvLlp7ovJh9g4Hu6
aORV3e/hhP3qSwedcFgOZ2gEAjlzxNPzwKf4YShGofUcreSVwcRg20mL90PT1pFE
nYeXca9goXb5bXRzvZ6ChmGa1vofNo70rasLAm3DtGfRCd10a6fCpt+eA6CXsiss
QoI/JU4+idHez2SRhm7sZ5ZcBbaZYHy2I6/d0xxF6IAcqYyeD9YjTTC5+ZYSYWG0
xJdSyVXIDtbeu4ij8QLs/Q0tglqKgsnW51Me7Ovm7Tvxy3w5fqQHgk0nAa54+qCC
1o/ddJlIVcOb9oB2RqyBAHpupIBU0JYq24FlJKn+2zjsEdkxjc2FO04u+7A8tL/v
1H21PGZTM3ttHndVX3FtYFWSNE+CkC5sBJGyBQ9nVnwnXXMFhioxInN/Ev/nfIOh
WcG17Myy/8VwxyCgOVh/lULMQDg0YHw0+H3OR++4GfthKmjytue/dUvl6aoPCjae
6GHkNVRpTzsDHVelMDePtZoK/78ZNc5MZLaP87Pp75UDzel4ZMe1r0GSJpwqkOau
Tt7jGCFE8E4GKQad1UPOKUHW+iTK8eDCkfim3oAV+yJ+XZ8qmrtvq8VAlIYiW0qd
bsSOa4byF74CxqhptkD7k5C22QgyutI95JFLWc9USetd+K/2q60ZlnDTPfsuvmAs
9Og16RpbjNJN/kQ4gpSc8Uu7K8MzUyBpuZvJDTFEctIgxPAcv1yp2EbZiZHO9myi
rMWt2EooTUFptAlIj1EBv8NwcjBG7FdEzqjApUcmO+rGdCpyfjGf6qWSB9H38j3h
EQorUOSP24y00Ob7tjX5k/7DQMDREwVMXAi1B0D1Xu1nt34MqCGphiEVZQ26S02c
cdE8dtmykfUzSPo8j5AVt72MTT/MQDHvUeGu1c4SkDJiBbKtmIfJyYGBGR+CRJ5E
XMDKnoxQsk3JvGFxm1zzAqLEusctf3z6z24r+2RWvMpU5NFPlLHj19smROYYa5Q+
iq6P7/9MeB9Hwi3pEJ/g8vqPfP1vn/jdBEb3D/2FjCQlFATtX1q2j579k/Om/FRw
wbHwwdMUzI5IB8c7H1bJ3edMLQBu+S7aTcGz5IS8ewYfh3KQ/BQT/QTlNJ2vW0z5
/iHwPLovtA/QRSWPxSjTmNbXDIfsmag0WVbwSFgQQDjMuSU03XyfFRpHx+rDCpae
riLe1Pydn+RamJd8ulZrCu1B0nizhBqL3QZapG/ctkDkiAR8FBAxDCz1MLJjmxiJ
o6mZoJYW7RV6cV3vFxDB1ohbUxTNeElSDo4xIOuvsZS5MBcCOXXO1K83sxPcvr0w
OH9NWh853xTzjD4+JKdI37ihANFPRwNfOXiDgiKuQfwQYxUm1BZ8nUpZUqx+6N5Q
WeWmCaeNXyDT/aZFM/514EgSTkgrcYrx2N+7M8alrfoiDXtAcaAbgezPQ7Mz0wLs
xRoay78QleXrWwBVvDDteVbI/Lc6S/PNrrHEFAftFeo9lChimBTHxheLvK2Yfp7t
GYsyak9x2/8O1ALfKRxPgX0WNE4q1R+JcQJR7aXJewnxqhq8XxgvYDZcRzd9fOhq
sHC78p7fpzrSpEd86s6ngdzOm5R+vBWMVFApSTKnXYAP6JKkPN8fttXApQgvnzjy
wkIhCHp/JwRxPDHkAU8jvUiFJ5VF/Jy4CIhIqW3oXndbEyz0BaZWhuKxmX0LQb96
XumbLGmrJmNULuf66vMCrZP2IPsh9cHPp/knnpU7IJNuP+qBMxU3Hnuw50OuZKnN
PWuIolNg9bv4vL+1STrELBRlEJDdKXtxa7sptWWMZfRcN8BKdBGGpbPwKztsP3FN
CanTTxkpEDYNY9DkFSylAPUupva8P5PcpgCd5F1yOdXwXvMWyZhYBATLbl2dus2L
opQa7fnKKQ5Qpn4KQUSmrgE8jwRgf6aM/sOGDiGg9m0g0aqsNjx91jH8bx1IHgcL
vm/i3lTDmwsD4aTcJD/pn+p6JNX16JfMLSCcJJ6R4xH+sr1WJks+ouKPEu+1iBCA
Jd+L5XF/sXl7WMXSi1B8Do8wwFb3JnOWE0Xkg1yfQCzxYgnz6LMCvUhjm/3j29pX
RU2vAOF0fo6nabKLfN4N3IedKe4jAeORIJFKSDxLcED0sakzY84xldug8c3BKC8U
DPIFH7u+HMYvNZaxc4re0BqkcqoVKVAWO+tOL6CfdZPF18BkYQUNkkDo9b/mRFIW
Cn8aeiP1orqCREVZ3OnHM2gi2XiEJJh1akKMJ/ZhZ/0yqBlcqbxc53VInK2I+gh4
Hlw+Pxnzcan46ibvjQ5MKlLa0UzxiDdyGaKaic1QYr+XXQRO4HorrtOnWxslot8+
DIukcr2uBHKSNcFoCOuSAQjhNcua4Vv0vbsKXefJqyLL+lfR8JkYNQJ5vOt0FBUi
VKAPX/2xh20DKiVg+4tMzzlrk5Ro2cKn7ygRLgtda3bwXbDmFA9BbPwixU/VdjCL
99BNbAHYDU6abl0cTxmIRgHd6v2HD2mNWjwbDPy/S+36j+hW7Uj11QyqlgXTl2AZ
hLTAgOsNTopXlvw08rvqftdJW+T4TZltlU11xKeSKHaXjQf3RhdmtvHDMvb9rhYy
fqkK1aBVa2dSl6EhoB66AoILZ78Ns8e76sIDgnwNFNiAGW9y5BNxBftDN3o4aWsU
MEn3nS0d1VPzrSF/n3pBXYpFd4t/IYOTrotkB+sohLcdr3tP3JTorrOwr1T7UuL/
kae5EscPjrorR8pbLxxbM/jt25+yMln3meazyjGYYE2cQubf8fcEimgPS7hAikmK
gPyJgSCLhAFLgbI09FnZ53bszJVaRt8CAtV+ehlLZjXfBFVKkGPY/YrwzW1RfIx6
QLQXQZVwrY8EiYWhVvSEFBOz33GfMqSObgoNWcM1lUqXaZgTzcdjHqFw/4zLRaW9
245K/2phZttw9CJbcFmntoWpZJImNrffQZi3nxv9OXeGt4RFgmu/h9TRFcTgvS5G
gFp7guR8pMlnMlNWuob567pX4sszHgx1BP1jpTDNKk3FKJCtwE8B4hh/GiydYJh9
sNM7qdnfumGQDGQciK1TlWHSXmf1IsLoetjJmuSzda64UyVExvc4O6pu/7hGoSrv
laU0w3bivTUyrOCmDun0/Uj5KgdIEV2itMuH8tZrb+y4miB5x/FHKRUDVawjxVIJ
hmyGdYVUf7hHR+HZxC+pnFJ3LyHEShITVpmAX9Re9S3k37v3Ud2NSa7W5Zfbbm8V
LhJ/AFAQRIJEmhYaGdgDmij3C8UgVoCXdz3p58S5WNMa3QhD7osJ2/0g7vozN+y4
vJ1G1Nf2BIUjRN2xrWiAwtyJHdImoOR2vjJ1OjzTQ/7m27M4XzMhJXUV031ctKL6
CZZCMaOg6GbrBy5dHQQTVuWTGPJavBJgAbWSy4ssWHPlTruenPah7I3s7+v7H8DO
3JjI21CkyPD+I6P+2TnZrVPfhzeMp6gzW7qqWT2hTZR3U4QH+7l/+Lh8Iqe/AzsS
BsOtAU6/fmIiIhINCouyQGQ2sYjbKAp1Jy8SV4UVDjwvy9GJRFYjDZndxp42pnlz
tLScgfd3tKDnRknKRd0rSV25b4aqTsw6KC147AoFyOD7qzC+zUrAqfI5Dg2HeU6M
G2h2UHEMk/q4vajNdH4vIkAiPb9HLyt7alS8lomSTSGDaC00m+rsavKujfkIPPp/
6tza/lMZJWcZgp1Auf5mroSzdqr27gvUxCr/Y9Oe3L7dXMXSBgTZTLycuvi6nEhA
lH9DAbL2SMV9aMwfIS/eUacY5tnRF9e88ImDXNPiYYqKsv41PDE9YnrE09HJIY63
6wIy934T5KWKgsOInZJHJcD5+0DMaKT6C/1mtgropboz4tneLJ/hy+miieYm7n5O
dIAckVE6ZvTRBsudwiqQPrXH9lUPYnDCxnnkqPNRP4LaCBfVWnL+hkjwHF9fYbpr
3cMF0QPr3G2IQQk/V6/t1UTEV+8JqKrfPD6ARkh9BUalsOFgabIrN04/OsmZvYnE
Ps7LrcimYTmLBx9hHuogaOBwaZux4XG0ZLTtM1USCRxI3RSdGXCryU8aYOfFWNFa
n1bEafSfkuz9DvPuUcGHToBjnddIPzE3kTJhtiUdNS4cUFoAU1AHrp99URQYePH8
rcctol33DCrC0AheTUxT6lZmptMfqwJi0gUWaNj5OAcr2EneXwHOf83WfL/u0tNd
D71tjAnc5TfFedgTr0kN9sY8ixzLj7mcdlvVDO0QhrptWevyg5g+IotrwSzHaTKB
rrdUoOsBp1WIXpGce0FAlmKF2Vbv4YzGtUqMyyFm+5jlccJcEcv6tiWYVh4sTY99
xYcjqfoXPhIhveM2IPN6HM3qnCSS7Md9MfjZqS7IE602uqTxWWDsckXnbUaxL7E4
t75Ls0Go2FCHw4Iy12KiO9pup2mySc3IMI+HtsJu5RtZeEyXT5XINxEMdi5fYGlu
tDREkt0Dw2gvYYbZDnNYtGggd/NDmJ8BEsi+lmlubfYxO1BB0EFSvyVSmT1Oeoeo
Mm8bZYjm0wEb0sKso/TG05oTjMlXY1QqO2X3LUlyaFelYKsKF96TRWwCpX0qn7tA
sVUSkTq8RQt1ToHitL8+/8yfNmWcvX/tJwfeIaIPhInVljYm9Mwesr35qaQBMtTT
W1pgby5IRcIt+T1HwSmnDGyD4wv6h3TYH8SUv3d8ddvuL8y8ycg9rg10ziHPYPfQ
uHITZEPAp5ww9+p7AACxCKpP/5meb1WSwjrjOVZe9HmoZJayWWtIu6LydqIYPyPD
W7En6/7b9n87pcauCmrkx8ENhdvKwWeUAMzAovDnyDUDpfGWGPJXa8orRi6NKinL
fmzJCRDD8r4xcqVXtUThxTb///+BUIF7xFDjODwi0aBXXYdNHXno6DrsLibOO9kK
Y1IcWLEuJAxvXXiNU+lEtocxoc0hbIPqnanK2A7lbmWh7cDJe2pdkIVd3lsXYuoi
7CJdI/ltUkAPql/O7QRyzirKCfPuYWXxTkaJGX6W202nDLYPXFeNDBiPd/U9gXNY
JSPHiQznGnau2Vmdauw76fCKlxi6JE58fEDmruPi7PFUQtrNyKwabQdDlqZtoWQu
Glb11dp0yPuEgqb6ofxgeZwEdNNYLy/WI/WvLguO0tVW1/sbZanoSCuSpYiDUHcQ
IWzhfEaFMgHpe0Hn1MiQJtAoP7199HPm64h+uLm/k8vS5NcsWNfzOz7DtdYQ7SFh
DvYMQD/ufaZ8xoP4g4DscokmZyH+dm0a+iVTrxWxK89bD27MbDCzAXG6c0RitWjb
lo2Cde3jUiVcEh/Cz91CHGz2yig90/96FkQWMErVDQl/mgWni6jroiv3RAdhxQEt
9pZOiZWJ0LYIEm4wNcrhSWznkmXo1h+kab8olT2Ydh3uPO+sY54ScuYFSmeVFt7D
g/fBLOqkFiA5JmdUx822yUZDk2ow5KnclR0fkrDcPZFFFdbJXwBy1qChHjTeCTWZ
DTXlOzdFWoNz7HlIzp1tOBFqAA2OwH0jRStWy7vye2F1X7AqOPhh5YcNG8xa5c2p
uiOEUhbZbeL7BA7GS47AL1inlexnwNJ/4nuHPXye4XeA7vqN5hTqzBfG3HZyixCR
ZtegLOLCDYhDevOcyeVyUUREvm8XlidaG1yVGtssfsN1S3fQzBGzCUzHbcXdHtXE
vTNfhkxPLi4KABtYXeod6V77UE2I7Gga4yvSsCHU1Y5S03+DWCe3/N7vwrYdXmo+
yDIfJIz2Hu5IIpzaeAbwPLMSgqNUIpF2q387JOZE38UQ5HZmdJ/u8g/TDhUNNbPz
hESgi1tzlAB0tnBYtbYiJL9N3NOK7YTGZskHlYFz0EeIKwuHEe220u5KFBiIUYIo
cpmDvROeCTjvMbSog7T6SdmxBLq8VVoXNxoLWgFtl82mpOJizvfnuh2ipNM5QiGT
KgBK3wyOeMvRS45qhGX6gICO4Dp5bTBFO1Uq7QlbGPG/9vW329cN2t0fO13iVbZG
/N3175Unh6VQ4erMLfyrHgij+3fkSUvtYHmnTn2jsyZKbXqb+IfvaKaqEn6MqhsH
mgEtYSTOcgGNB84kQY+mKyDAtO+n6O4rr0RZVBGTNux0kc8fatpm1sbBXsQK3RI2
WTjktYrEV3B9UDWxfhMwM6DdrWGNJ9yzoMDzpp3YdmLfJNz0FpOL2KC4o8YnoRFO
ubYSYF86d2qliBSpoPbw88qJN7QtbH2iS9NG5n02T7anb62oKLkovzBwJMox6Wte
CkiU1EibHRyEl8BsaI/OZEzdxLKceAzlSHnSJj3CxOW9XLY7FY7n3BSpVTldh3bh
bnI+dmcVcGPoeyQxNz5QG0MWpUUtLR73+6QQXgSzFDNyo9S5FD3AfjG0g7KUFQ46
cPzJSYut6fBlig+1Ev4e1FJX6uX8PLYD0/+3g0OYozIG8K1oISf+qoVq2ydih4FR
1JOHW4SsCtpF4z0+Q+LSZTKJl8lkdO3HDEfG+XkdhhHqkOItvDOiXKqM6z+TAHhE
/zTazGcBQ86sAdFz/z4blnICUTU28ZcXxOwfHdrEqswOkkUv5SGZ6l0/oOxtmpPL
VC230JAhSPy3w2d66SBFSx8TvE5p4JELpVFNLLVLnTigF8H6w5TWBgw5Qrrq5Nt1
wYRonFCOakSGuIYduysOrwdy6vG3amwamEvw5jn921SeMXb5SxZABqOrYyRiWWuH
qWmQNUeHAQxN35jKsVGz+syWxh5N8l1bIedih4ebwj5IJ4N1IvxP3l1tY8sXoSXO
HAjOY2UWoQj36BiC/dGoFBNL9KinJ4l07D1uAIgR2d0prWkGUqd72p+UC9D+A0B5
JhurYWZjgIZJ+BJsWkYnG+85vhgOnFlN9BZSrjGRbTXF0TVDa5+lXWp2f5U3Vd/d
I7kS+90MatIC9mjK1inIbNzSIGws2HNDomUfUd9D+bEL/6b4r79RooYhsH9c35aT
JprZkluosHMEX83DxOn/E2R+SCq8n59zqc65sI4MlcsEPscMNE8AKrNX3RGRMUQa
9NmQbIqxcQkSWS1pNj2e/ojQaWkbetGlQjKrt4nUBvtn321bfspBNCESKGGx+5R2
60ie1wYd0AXxZNmKkDSLq2GUR6pHT9MV0Xmzch35i111X4xwGHJWFl9E+d4u7cOK
Z7NcDr7zd+OYGJEDpMYS51mmxzm8lyzfx8uKTdwpkMnZlOet7pfed7LDjBBSrAzE
xFYrVC+iMrBiVm2lfo9cigiG735f3UmRUq4kEto3Pv3+cKYoSequp+A9xRLe96w4
LpVg+w7tqba7ddlCCAEoIykdqXrzOk7SCNpN5rRoFtGeVCjf8vE2n9Z0E4jqwYf7
52Vt22YyhpdHXfcdpFdJcxvqNN5BdGqTWD1sPkLCy4+9Z1Wl0vJr4EWZ8LQewCu8
jGErpdY8gOghEeXKLqZIjk/RRU4DG8hYUy5sMi3Kk59KMM8aWDZM3Eaiex9tnjW9
UkK0MCFpb2D3OCebTOWJMSkR21P1taWY2/fC2HrE6pDBralls+MdxUYmTzdtv93v
MzzTjKy7JVLnrcVSPKyO+iEU8rYgmTthUKJZemxodmiBIwcroAX1r1sxHwYCpDSS
NpxgjfXMIThHtlDwudtLPWI6W/y2T9LSqqVhS1KcQ9/fMfAj7reCu/7CRxfc1Hf4
pjmOPHmPau9xwxPMw56lxzQ5/auJh+WNvYLUzgmY7uZ0EZ27nB/OT8aMMkE+qCNB
baXTWpzo8RRTtaLPLFz9Y1H1Ih8rOgkGRgY23de5DfYXhLCp4p6JdKCoKWCU2hTK
LrK6rujUF9V0ehgVU/4SjpxlNIt6Sl66nkdADrboy431zDSoPjq2e4OR4+kvBCdG
2dK6kRN6epR81K9l+VRJkkUpp0cWSPuqfnLDobjsRx744ZDb22F5vXHoXcnGGUt4
hSGmGXG0/79gIXEQaw8hOlGJ7XIG7AfHVP9vpb3OHHggi+0UYa6gfFqpKOpJqbNU
5lUVYIiziDAc7PAw6UTt8LdM4gTsBs2Rn06VinGigDY59rkDCnBrLozaMSbMCPzs
+5ewW735zQE8PTcE2piF4udkW7IW0joyRBFsemrLdelhrEZILTO7JKtgWnoi0/Xb
3KD0Gy46EWDjfjQ+fucqDxSNs+a89AUUi4dIAdSBe6RXOyeL8A7FfQVbRdPVbYbV
V4G0ZSOUoSQQHIJT85kj7cqK0XdLrSY9/KrIFrbIl4xdu1f8Ppr/x2KumUfQC172
2EjI7pzhryQtpwMql7+IgO2UAMbrJo/mzEmsS9JoSODBBYRrYguP+f0qrSIuKyn3
4s9mV51t985qFLGoWJ1TLFw/KOiRjzdB6+x5o0mJqzarmt2Ot5RFMiNlkZspUfkN
hhJ2Impn78L8hWJphKD9oQyGhPhDNTjA1O5NbXunvdtBxASKmY/iSmYGhNv5T8lQ
SRvKKJAYKx1Vx7++W7BQ1eNTUthrllHyTo+z6YO4FeCt2R8mNMpMhJ4KqVSQxlOh
mPzHIcIvTRXoIHvvelal5widvkZlUWarvIbetClYc8l2cG7BTxEZfdButqei5KZL
HqLts8ZrAeoTf3l4FnHk+Q0QALreoVeZdaONXXC1GKR3TIqbkgSP4V0IeRAfyJ6I
iYzN67nNTlrPVQqX3k7+LpTBwBK0Ypzj6g3g9cAl3FNaMb4PsVWapjZL7UvyO1F7
YgUSBn5f45D56J9OofJNivO+xdC9cPe8P00huhCCIIZyNndwoPe28IEBqhVaxZJa
NdFVCvDdVmVZE1S70uJGJoLJ+9fecyez4gyHQfs+HKWltwf2at32TCZjVKtE6Ii/
BCVFhUtjshBcbtsb8YbFIfnnfignTUvtf+XVIqFkEdBzGI4Yjv2UMVoseQMgbzwN
eOFX+4CRcvr/fpnRWtwZMz8pGXN2G6kWo1S5Ef+zIiD2rLFhrNJkUu+YkvmkeHb9
N2dtHCh2hxzRB9agVd2zL8U8V3GiSk3J+DwkpPuvQQWo9dRzYioXU4Skf2E5M/fh
W1lcSHvWNykBJH4F5KBkV0+KDoKMSmEMqWR66TKtlHQTdp7Btg/kt6pLjrQ9EGst
yClt1UpPYh3eFLHxU7nJ4JJLMRAC8cSBi2aIje7hhzCnlLwRh1w2aDcZ0GZCWqp1
FiALTmvPOcGuk4NjrUklwnAwA7GxRmrzySMVUI7O1uw6Hjc7jN32Ipyg73JKVgfF
dAIgFFgAZJPqEzJKLuNrCbiKDxzshmuz15s6bK/mkXem9dLiYOx20paFdUCuQlfd
NKeIpsSMOf5UPU88+vCRZJtsnqcNFZqt3LEPM8LR4lS+U4I89Jf1LBAoiRwF5Ivu
m5OdatxtExoBC9Kv4GAuTv3c8OummELJzxOdHR/3pKv+2Ywzt9Y6rW0QtqqrR4db
RvWanq4rYa6etOAgreBAEMjHnehd3WYl/MlrCLg4ng2sXxclOOBlpi/sITQXVX+d
sgV/ilUkXuJT220t37GZUbRvEi08zS+cmiUIwu/jFgJ5Emj0uqNN/W7ho0A+op9b
Rs5uaZBbd3EwZGA04RhnDh7hXPd8uQ8GkExoljeuMPW7Y8H7OqWYH4PYGWps8G4L
lK80LO+wQdR2rbpdsd2gmhIeis/2LKMFmzgkDe7hMimS7o5GUiF1z2y0ALlzngw0
BMpCJfsFcztrA37RVOFQdtDjoQ7oFaLmyrAen8bSf74c5d4DbznMmZ2avP/c0f/5
AQ+m4GqOhMX1GxFKshqUB7Th/LxcEahY0T3kd2czQn5CPYuMme4t1E3I/YIsTu28
V2eA/cSCA9DtKiDPpXDeUT6gODMJVnOTKrb0QdiNxGIAd0zDAALWxUW1fg/5s5y8
yF952TnZQXwMCHC414vpcfks9Kr8NPHP9X/r84jHwRLjRE7MStlmXgZgELFoUGLn
F5FZV6SJm7UYdD84ADR+yqzYm2pmY9IZMTnFnVq4hU3K3sA/iJKHgoebTtpXbsK1
XRtPgE66wE9XpjjRc3lxIzJb24zQ95Py3hwR8yTjVwkX+TL/Kf18V3qF/OHr8wVu
QV9abI2si3tA1zaMbiSXvNLB/GnOPsRuNfVff+vJ7p85MEB326JpyWMrEF2CltPg
VIOdprqzPbPkoqreSJ99Bli6nhT77GKuT0Q8Hu4FfAfjUxJ266zVTe5cUcDzQ4Se
LlqyKDuNoncG9nFOOUELHeZAB8I+HRC1dQGo6xnpaOZCDqY8Mt6pUXVURBEmazdV
AMKlxs/sysEddHq3lAhzUThivkfEAEwKiZ9nFdu6NeNZJboK0pyYJOYIh36jNHG6
45z8mWxQJyuR1Ccynh6ah8mBmMIdLKoO1EADTFmSdiVOJTYYznCiQLklS7qSBz/x
PAYJRV6qE5My99/M0GrqCcqIFwYpnD01xcqKPZD64eQBdUd57Kue+LuEoay4S5Zy
PqLOnLhmEQvG1G0vYRmoupXE6xgAmD6re8awkTEC5gwJQQ+KAmm8j2bCAz0Gc3hm
idmmhz1CXGJWv542Lz2/LgKblKTQcn0J/OZE2BRAbCfR/up7OsrRC8XWflVLhRuJ
pAGZDf04uS7GWcmbLRVeBtg2/XqHPUVewIKwWcLdAf5O6GpiQM85O1RtsYU5fLhJ
WJOQ38aVI3/+O3nSxVIoTPem7TwWNiqPdi70DBVBAwpLh19OrkamRXA5Fr2RmbS1
Wi4I76kvWdaliY0mSSYO4BQm9GO5/bdEYm3rpLfewDETdnOPorjpv/DuiVXIfKWj
tVudxrisR4I5SG0KEWlCxTfYIOP0+v4uGK98ieZWQ5ipUJQidN90/dk59me2yn0N
8RWfcMyz7Y4p6cCUwEKnePWDZU1emtjTzeRNauxC1HeH2Ot01cFMUqLwl1910y/Y
U5JrDg2lQ7QjbiwGw9kOhkt80cjJXQ+WpWr2JRyBUB79YICc2ODJQsBtAdJ7z6CZ
5w+JbSN1MbS5e5vm/de5YpcHmevqCIX9nTN5rd+MWIMupQmT7DUqNqZ47i/n+y0X
VUROo9doOop9U+9APNc7X86qEfwHxGwV4YngsxpBJT3C+TorU0uM6oWRLZaSNDt9
h3x0J6FLUmIKZ80f0XzBz/1cM/EKSQvtrzS3gELniotYMl7LtmfNF4a478A05jSI
y100UI8xt4JcB87vkrlAyG1yewy5q+ehI/hi+3NwEoyNL/ean2s5qGhgECRRg+gP
oOAqROwFg4eGDvkB6THR5cj4bgtTQOganavHZdgnoy32Tdl0t/tzB6O6Per2SOcU
rFXTkhcTgNiEpqttR1aaPxU5oQQqbtUQ6eN76KnkJ26ByM1RcuM3vEcqDZJwTgB8
OkcF2YJReR4Of1Ml4fYTc0tQLiPdsnd6Aa3HCGD0YyLKkuTbuBzdUMUZQXdsnntX
yQxk5qvGFXY1JwlagD1YOhF4OWmzo6YbsqJaBwrOtpoRUYtYDvJRL7ZKxucTFhMq
Grj16gX5R3R2oRLh334jTd5GN5gsQul5MB1PAS6zNBmg9ipJqwhTSM6Pkd/a+bBJ
bgDEEs9exkZIpdQfZt8x/D/bkwJVW0a9gpZtCGV4fRTtB49pK8SB3/bglkxgMD+F
DwZ9AwgVikQR/YYPRK63YzJnXb7Y4sTCFO5mAJSmfxBY0Ei+eP2zkiJMWu0wyalt
rIAW9WA3P9HnpTnS8w6UOE9xSEqrtHe4MNHcjLWoF1k5cszqomN0bj8w5OEEGPKG
3dyyQ64nYv4HEXBXoOSyAlYZ6mCjQ30XW8tUU6rKYSTTtc+zeXUHFD5LdYeozdZU
9nHYL1QK16q5tbX6NflBF0NiWiPYcQe5hLjLSVeITh7gyT71WxnGSDqAH+30ne59
9INFG0hnVzLCu4KYifZLYUJ4jb2g6jkYMrAS3G+M70YGq6UvR4B4Ifnnncdbk9FT
rNz7nn8BsmuDKM/6i+Llo6+SGYtPdVMW/Nb36n1fcyAguu5uNeio43mmSNRpQYtq
Wji7WrKsAbsw3xyGvuCsOsud6s++s+YjeB4DN6kPjb5RR74l3xD8aDrDhHbmS426
zXS7Zms0eS4rLXLgcE2Unc3aqGGeC+6kMYnOHV8nKgLJ/eRqoVJXxSXc5dD9sbv9
iiaZ8AzCk7kFN3IgIRmtff7q/K0rvk3R1iN2iITC0eky0j/3Nrn58dnWfEP7r0z2
T5wx2mK3EHYQ4l2dbc3bev7N9zVNcKbR3+xPV1A8lU9NQPu3wuoYhA0pV8/QAal3
XG75YvXE9EKOObvKjGEWS9FywGl3x4rhsbTDD+y14uOUYizDRQrdl1LccpjZZrV+
ewgnWIw4xhct+Tbx8G31ZAMYjTMJ5HRmHoXr0f3+l4YwCXLi2c7z9BPEXec78Shb
6N7qg0+MeB9SPrCh3SNKXrpKTv1NXGXRkWNoCeoUAM5QhkbKfRbXW46+c6suVWxU
QqzOLX6f10LUsHo4Cb933addCz/UKla1GPCDxpgiTPyo+Lhgau7fO8FXVjVQuL1k
Atig9U4OmsE1JP5utTHdRY2zqYLdEECZC1y1ghIw+nijKa+yz157oxa7ehbuj/cm
shklA2T2OoUyPXIdB7pbTCnepGf6rFcMHwCwmr9XjTvVl75migswtWM5LvF9sA1B
k7/nzu76SKArUY3E05NxQY4ioGTbdfcaYonI7UMbz0mxNMO1yeyclQj5YS4AjeWs
CyD8A3MRLzaxdKRBlyxSJBGA0QBjGySeL9oqVmC2uDkEmjUTkGL+QvzZaXdc68Bf
ea7ibjq/SUFxw9OfQkM2vIDKGPwK7wp2VTME3HUwMF2NVyqOzy68hWUYAiUsSBgn
Asd59bqMIdARc13/X9r5XHJNbSdCxg57l5a+R3OBdB1nVTYoA4aj37tUMUGCJFBq
9/DIG1WDz9fNEy/CGcs3h+6uxkKDvdmRXMoCiS9N7VR8fwQOqSdmyy9GGDltbV62
NCifMzu7Lo2cHc8hCXv/+MR3p2veSRfDiSRaQRmv/XhpCz/DqXh8DXI9/x+n5jzD
2gPXEPT75XvR0J2EM3Mdb55ihItqura78FMAFvP7PRJX0fuPfZGaX7AeD9HwXCkz
SXBPpHwJP3RZsDHroztvDMdulqTN+Z8z/mwXLblF2SrGefTG3LnMC5PCnsBBIWNW
zIZKcNi5aliqNGh26sipes05Ex9/CGQkUOXBngfJ/mqZ3oejiRa/V9i3kxfLNoqT
1Ci6Gtx6apovOjw/s6o4XBsXeMZ8HSmHyTXVnkkX6Yb99F9dm7+DAvmalCU8DlU1
kGu4E8fF2Ff5wNSWEgPsO9SS7ayIV5AKxHQH8R8cxbE/lPOONj+/5z0U2NqH2OJ5
zSiI+4jHz4Ug8DZ5qzvPvrLC09QV+EmCwfaZhcenQps8M1EE9el1Lf5v6Y+/JW/L
z8tVNi6OCZCakqjfW7hJ2wBwx4OLCjQbS6Ku480PI1VAblm0A0kh/SKJf/mEmk1j
t8JNPN8H4jAcWZ2Gq6VjuajJuE1iLRNERKpYYRH/Baoj4Fb7jBcE3v0Z++4MS1LH
p8lvDZnDwR3+hvUmiE9SVGRU9G64ujCjYJWL8BlKnD5yNyWmQYw7OJTTZU3cDKsJ
1CEb++5ICguLSSq/mzHrANs3vEzM9xdmdy4EeF74yNCX1n2q3h996k6c3PhCvALi
oZUeWnzgIPpxWczWrBnUmfcOOdmjYbU+/cyxRs83wobcUr0EVO/NdoEDJVzz37TI
4e6s5+8CKwI9dNVbq8MU/qIMzxJmcZSpVQCT9IaVJb7mhsipOtNbhbBdPrOfqk2Q
tUtLbVdvOjlCn2Uztux2OtuEGMqBOT1tlniJg1U2XtjP5iRBeUJWu8r9+bnwUXLh
zXiRWmkrKF2quZwhVH5/nln2v7mIbtgGokXnNyPZ96ITIZzbcfwIDBToPl8Hhll3
LDqAPBwzFvix4/RVnvFAfgmyNeS8+qkJDNQYzBHnSiBK0HUiXXhgviq0L5kqCOA3
gc3OaMF2NzOTyHGmtzviGlUcrlOuHW9VRvuu0cWMHhn80tXDwjLxg6gvwo4K1rKq
0nyPsrixpjGS9Nc19RHqPto6JwQjLGUP3ymL5dbGY0eOWdQ7n8MQrkg6nr4QW9/x
Y+KTwJj0U6gqCbCOj1r4VwEM5ly2/5Q3S1ZqX7WS51tZFbOk1yLiyvPM4xphHKuL
xwWz3FtsGExaCqDEGpRtfQnRi3IUEyLpSCBRswqPMdwDaJdY0nK5HbMx3B/GthBp
P5wvYtxFcb7K1EBZ3ReqPAn1OpDQtWWcBW3H51i2UT48BuqR571zgDfeWVLC7UcY
tAsWel9tXrT4JcWtGAIRttsJwyQPnkrkgPM4SwHtFdc9CWeaKHdp9Z8yZ37Kedsv
tx4H1M7/sXEyVNsgjGwN3FcvfLFR0P2C4hZ+NbKINvWkvhRInGYPPKyajbgrAr2Y
cjPTVnxHndJDUZYsEl4tDS7ns2vueN0wnFSC3M0OF/cV8OWt4fqDmOsJ0H6Q9Eqr
sdZlIZFS+XS3kHeOtfjpce/yKYo2Yu2tvU9jfhPv1UPRiBdHujGBlWiTlX1YcbRv
p4LLvehr98NwnpcaFIL1eNEjxBT/FTqKZN4l4ZJr84ecRVfZ4lldMAfppbZ9WpWj
mGSfn8jfH7hcOc2e3ILP2WXOrMeaejQb/9uK9H0EsfVKBYYKHMnDPMhCZSMOVeNF
j5JYuzeCHEP/SldoIsPTIbrWZdUL7NJh5xwrpACGBBr9IWxzx6orO4kYmKJKomYv
wFIoKj0x8opc6vCjSBvO78VNtLkz0NDOygqKLe2y6A9ZOdPW5o9jI2rDEQ3hFZRh
oqBOa7SYVsWs7nyJylQBEFuk6kVjGb5+sSK1aTYCLlQ4nwiyEja9ujiG1dW9RaUc
1Uf4xROJnRSvdRffP4dzS+jmpi4ggbxrb7zmXwbNDs5LahSZS1hcXLzEcj01oTZq
PMlOYIc89r8KA+ORBFIfEaqcqjFTMDqS+EGCbIZfPasVlpu3NqdD7NDXzQh1FLS5
XAKR+kDfzKPHuNFF3Skp4MUSfgZhyutK3K01bXsaqMCPcJ1ZL23QKyhL3wFZNwNU
qwuKhHzsUPdtTYAJHuKuDHXyvrMuzNSMLOwhQ3T1zNXKMg1Z+2VeK1bcN69OH8Ne
HuNttLw9JeH7bAtJjsJRfH2Bp8e3cDwukYwmgoM12RHaoVaUwgLjW4mX7fP3LYiC
6e61MZizEVqwEHLjXneE30z5dsIeBWB5qWqAbJMoK5rx3Q8Li55uwDCoy83ixwd9
W01HYGxZH/SHMZoGYz90tW5pJy7/sjA0eW6YEO/xhvpGlD3RR+R9Tx0HTOnjMEBP
IFUPZgJPfozJsiG0cGhb9kbfpf8f19C0SYn2bUDY1MIxwJZEvKcG79g9zfCwwla2
RTT3P4OZldl2ylvziCRIKV/PtSZAtbSQjNo4CKDGjawvD6shFyDzt74SuKYqeTLc
vofbGhgohVIsJ66L4BrlPWH8t6MCjFQ/g18MDr1vu1yZFC7lEp7b9VIEKOWkOpQk
QZs9HiYOXXYTSy6gjcWiwfLGVKHu4DgWgZjLHQXEK9b3Fj3EclkhcSaRWa3pFNim
uMw4LHVFGgsr7jezL6g26lEUeb62u0iQlXCWqVI4aPlvTV9a46c0/eCj2Ks0GPeK
GDHxA2b6AKNFmgViFj3Fu1Zl0kZVWg7sTSP7PEoPaQ6koxX06jvqmbySpyhVl+0k
4H6Xt4sWAXiYY1MthnpQGz+4ae0zu7BhOPYNd/2wu+nXGZmsdaBcjdY2o7k8Veez
TsMChDiQovk/q7t57ZZL1rFSGPZDw6iN4tfROQfzH6Bzo54kbkkv4YpJpRyqKTfJ
xpXvrGdZyOs49I2sV3dMw8dg2etBls1/lXhGHccvY7wPcY8H0+TQYbxuIz5ELekp
bGQ9r4RvFtg5RQ1gJbn93nONd8+DkqtPhwNfTg2dvfMnNWSZsWo8iPe3Al8D741E
fIXfMxZ4Pm+0qoxwCa3kfpsTvYei5cvTTCvqPLHzPyyK6D4Mh17WTR3sGgtrqKi2
BX0q9DkKzLVgNnlD0Yz52fH0S/ZgGE44cqHuvDEKdUOsxMbCYyRb9ImfIaZgrA19
zi5JC5UR0Wq70lPj+7qbIvgCvDRuqVXfNa/MX9UW8L4Y/nHc2Z+sHKn1UBmnym7L
zPFHUGRzTUKRqeBBQWxdGT4ZfMv9CG1GViv/UZJFiYWr/qJG9jMsRw8WjjWtB55M
DyntV+W73NvZX8BF4MU9wGBpAg5Vgrzx6zCUJY4Q0g7J96RNeYB9aAbkQ7X9CZsW
EFuPAdEuRmBbWQLZlsBc+YI5G+2033A0sqsNiFbodst4L5W4fjCA05hkD49DGqIL
PgCjRPcwkKM3KGXXvcW/1EceVInyFVa2dN5MovXHpO2ZIrtoZTLSjEd0sJ4tXTk7
vpa6KWjBU4uW3B7KcBD+isZz2epPKeOQRKIL8Q3i8hZQQPRfYQxZPdS/btzmnuvl
H/XQ3pc6CvxcqT1TYUz519yEJ/k8+6ad0kTIcPSAM3DZg2d4Vro0njaF8g6zZ9WA
cst10RC8BgU7XDWTOFYjI4GcRgzA3GRALW2m0+BJk6b2NFvOrbn+UpVgdgM0vqSI
fFAd3L0DrwiUKiZJ1gCEZgFLty4b7XoztaMEBMyYy58JYQ9sdG2ANNMBkxbyXNqu
/Ko3yyXAtipDqw8NpaEYEY5pt65v3TdgpHAqLgp25VKNp9A15qekCNu7I9A+PbtO
5o8bZa0YSKBUKs3O2/owu+Au1y/9dfFCWkibSHDsuJX2UaJWq4vtLbr6ozvGeMs1
jDg2aavnzFVXfUrP1ck8ID0Qxz9WgpgNqqqQgDosIQ0FKmbarG4TFfEcxXm5eJEM
FgLGXnWKIRX2gC/8h6VWKsRLZD/oyt/TzyNie7IDM2+s4hwCLa/pFFmrHJQGAIJH
XjOVAsKy3QN095101qV5pOM5eCj1pdFjTZoxiLiEYfHrwXi3snw2QFuJpc4ynZhj
UKQLMQhS3BDWySYMtA3LzxQGzMDjjIvrlh9HHl+9Tcz+30QHgY5wnwZ3kw7dt4xv
CK4x4wkeAFm/mT1bslUEnV9Zifumv6Xz7EctnQrZrbfoUtnxxy0emTarAPXYQrGS
HOIq32CzhHKsKfsozd5Sux4t0L2hiRDgpxuvWcNC+OkCL0D2FFWV63iGm+qCU2c0
h/mV3nrPgIHX4l3+q/v3UEvLNF1PWyY3wn6uun/sN8ScoJgbkmey8KX11/cOYGfu
ph5ZclZSsXrIj9wBm5mq9c0y5elk9+ACU5R8dEXFnNU7RnWbsi11dt9H+gvDKiUG
lY9aV+Rr1Df+/yxa3kqXTjtM1NUudmCZPk0WVkqx4rFPzdSSarLxEDyM8YKVW+iC
hD7G2Q6P/oUWOIGbLGvYkz0elNss94/1Qt/mjqp0REQkfp4eXF/CNA6kgVoNeLDd
jgcheXqqrZpgc9YFxesmubeg/oKM0ln9Xj66nA9pwnpg0RwvrjzYqDgjM7FMyVen
M2oLSWwc6sTfpHownlOyQvBJErjO8NIdWypuC/2Azz/3stQL7bE8xsfJQnQsU9eP
Kqxy9vd7QIGwC5GoukbvFoUludEzDRi0Iq44A7r3qAqpJb9eU+T42yDQ2gCKefR0
2i1VLI8jtu2khjfX6jpxcQULq4jqI32Pf0KUCjdpJZi3W1sJptrCzayH7Ze/338X
MYIlv/8xGrAxSfwSGFcIaksSl3IicnDZ2wRwjc63CnGhdA92x5WHjAdaRobV1pRP
28zw/TS3UmD/SckEOweNLtGOVBfwG6uTTpqWV4eoEvsTQlftJydQ4ZiQAFsAbd5m
6rAnlgPRhhIOsdkzAzIxR4rqW3VsBChsGZTvSyXUyAE9TZ52yo1SVsvxkAe1iln3
Zv06CvFYjM0wzLQrCS3R29Jn1KM+p2FVuFE17w0QBLYD/4kzg9igGohwH5YjUUFp
0Bq8QUguKlsKbHt3BDyf2T4/UPocORbfqLRUa1BIZhakyeyJHieDrISWOvHkwmGL
0goothvR6N0UO9Kxjk47Twn6WpWwAk9Rdg0h1uXN8Q3f4XwsIKi2Lju0v5sVWeK2
RUk/day74rnxtNOXmjfppyTpn4hNfk7eBzhYFJjAXQ/oNrK6eWxENrhVgFKHEzWR
A1oyh/CBYGXXVBYf35L68i8HxZHUh+LSzNyzvjuDiMuUfGrnTZnkruOFWTVJD3IX
oEvm3v1YsUw004Aqr46Ils08vzAp57bQZr8wXF8JFWJpd26rgmWC/KQJITObS1Zh
ekil81jrXM0d41wNi5YdhrJSNjrMzMwxuKsfQJcfejXlbuYVsJtNUeP7a9ESByfc
3ncF8QjjPb8QvqS+qqgWV25j9wHnCbbNE0J8XPm9mEr73L1aJDFXinox6K6AfqAX
GzTSJouv0hUl/Ll0w7QZMPrcoha5HwiuPOt//bXy7f79iN+3TxndX5ndnjXA3uTN
3z/doymTFa9TauBztVnMpxL5zkCtKgLIW3BKp0N95bQ2fXcGthtdT2t9K5QqoHTw
QnbvKIxRrhaZF4r8qiu71q5Rav3rRwXLPz5LIWzuHFsWJrl9Pgre3P2Cy6MAFerV
e5VY31n00Ow6QJmjiv1AMSkml3z88WsIVT2hpEFjnRnLGzXQ2/kz3splcDWoNEBI
otP51V0NXT3GN4tkXoBQRbs5vZALpCyDP56KO1/etWWzfhLVPKUTK1/Yn8k65yz8
ftl6fai9EyswM35i81GfAI4UoVwbMkJnJdxnaVHuI+HjAUx/HJYSuG+WvoV4PouS
SOMLwIAweCc90CuxQH2GBvYRVdjNiL18sa/M9VTSFpWkkO+JKbJArSNho/yteiFQ
D6U4duz0tgEE+OKbbx0MqOvwUZAyh0EDiECTqb8v9D3qvJf7VtK/dPxPFxUVcUlh
N3Ca88y5kM7OtVnMb4tIT9FMLLShx+eIUKVLexXqKOQUhIgY/DtDZQmNBQaDET7F
oS8nPXi3zeLXOdFMHpPgEb7btRocrQNBHFJoPSjesthDMbOMo5mhpBekTzHx0p2u
4jo4zhOp+x3wbRe+TwK/BxtLDPSC0p0Ql+fBD6bxsauSQsV51GLPA2CxcG+/MCJB
CAydBLctERFAlhgQGqzZIGusJgUoiAK6S3NSlxo7cUI+UBNohaLyLlbwUu1VtCuL
CsEDn8dClwYmFsqYK3AJOoBKUkDUQAhAq/FWtBugIXCbzEGB+FTLdaMitsU07G/C
4+t8MJ+DpTmsd9DvkJsyByNSXgwUSk0QrTlFj3LM4ZfCrXR/YSEFzVtFjJXYSLcq
rMrEKsWZmttCnzxmR2htpofvb1YfLDJEo4vQOZd6ftWcWcz6ZQ73fkwk84n4glQ/
QErzUnfh7SGE7+DVuoA1fE636/4btIYTUTtp9RXSqWxeE4rDW9ar4D/Y3O6WWd2k
rsk7ErphSWzLCDyBUkWqyQWBkJf3o8678bO+yvD0O6fTty0+2CxO9pVgw/weeMRr
KN0/sufG24sSxy5ACCEIREM1lZMcACfymo06iISm+2aNnLzE1SMj9e/worCWBubJ
sRCHBvhGcLejpE48bPW+zNed951kLX4zgZjyYuOwqC1HYNsuVilrpu9jyU/q3KYG
BEE5ySBKH7TMKMA4bEPQcRaMPMa8S07txIbJsekNCLw8+G+qTaLzEKDyNKp+gSvh
oeQXog7tYXlSJbyvObZrkEEKW4Af1Okk32UMdVAe6tU4zE0cpIXJN/ZI7Y+PVyyn
IEys1acDOefD2dTjbJHOtd3ml+kj7iXI78MyeyRgItmPTwCOrUc4MINB/E3cptg/
9w9CEeguZwCw46r2lo4m1rqSI4bm9HA0x2LQYR7yLxm4NffYeg+sQhd3ejFD48xz
wk6PApu/0xjW4F8465hkW4pdSHyUL7ULqv9bqG40gpINLxoMkMvzZa3uHhOihTVx
giBkS6En1lYIXINRQE/Aw6ql2oJXghpXeBgMoU09Bn1y9ZaWKoglFz9vQUIuRi0P
efBD7HZiu0YiNsPIbtntpJi2mQK4U7HvEDIL1VP1iq6dcX+Ucb9+MtFCzVYxRCV9
pjJxiMZ/IyNlD1tbzRH5uFTgGVPOZ+s1KkrqNy9QASiNdKt8GXYLFSr+j+jNMfCf
DKXy5CBpLE/sNrUnzJEhOIOHDAAovjSadt4CDSd889U237mxuSoQ54+sNrTyjbPq
wkOA2eJ1CITRoGjEqyIiVO7c+bm5jWfIYm4Lc13FJ9dwVUF8qkU6syMKS6YtrFAM
TjCLCOunSwjS/9qUkHv32x5Yc/oObTqjliL7qLWZ964rP9tidzd/O8nKjlurDhkM
Lxt7TMN6LYRAj1EnqzvgjSud2U+rcCTkO+ZDQSVO4A3gPQCTB76L+IczDxwz+Ha7
lx4seF7SVNq4Zlh+LBGi1YMfXdhxpHq1IHjK24jXzylLQ5R1ZvBqmc9Z0IAHE0l6
GTARZRqWMcbIRpSvuQQvENhaXbpqTK3icgWdfr2ZtAHlzs8z3QpjwDoi/CYLUI61
Uvg/gNzgSU631UuCA3AgTfKv5XiDZB6eQRnvf1tesbkeMwsgNduRxKTH3WGS4rDF
Ct+F7xBSf0HclugDxzJRGPy5RuaW5wjj4LWWnX6NFVab70V4xY9BHhmE8msbVC2j
a/3LzjGx4Fe0nz3sOGPmtDRjYF309WxSzG27RJ/2dykIdLIEwglxO6RvaB65mkjP
xL45Vx9Cj16kxIyeQVW/izhmW4xR1LL09Pmg4O6hCZb1uqVs9U5vfaN2oTr/7bWs
U4Zwrh2ZemdXIhOdl8O0cBlC/WrXCN3vao+BQ7Xe0g7+GxIOCop/6lq9QznUVDir
ArammWJJxnXtX7K1Eu6oquTayOfGjM/AxO8Y68JQDNMRcgqB6/A4iLagI3rOIeV7
2459An2NWUcsP711Sa8Q5owheNEXa6ob14DAwMhUzMRS+qaWu5AMhI8CT1HoQFQj
V+Lr6DglrkOTtwnvWmlc5wjeY7G073CnsmbqM4M9mIrwRiVkUzD7HPTiFmu1lYGg
j8Z0SOdsw7MroVnJDjDHG3gT2lqeYUSmuD8Hw3wUR1v7uT403O1mpMqDD1Iin0TX
vzx2JAMAHM1+sFpPlos3olRIYvv1H+Sjd7Xb4ixUKa+OGJHftLKsXUexwNKNejh2
MDBhLBrf3zbNW0JPM6WGd2FM8SPRvUx33MVYR9xfqjsTLnY66bSHfB3QYNE7JV7P
I2Ym4Lme7G/kvXQT0YgjCl5RaTmjMTtY8uC5XL9MXkwFnGK7cs/Q0O061Ixafp5f
h5hPGZLbyEv95kt+D/lR1SBpqXb5wQujtj+mfWVTZEiFWSWnTJIfit5AqTKTcp0E
/LC/tR9Lm6j1oLDo2d+VnMQpb8C7BcjUKNiuz3BCHZqTjZhzaTk2cjLMpBU+O2rb
4ghbm5UZ0yt516hCMQXaL3MFbbcXH7hh5dCY0E9SsInmsYnLjl4pI5729TCp+c1P
FMvF/Zpt4NSlnJeDfqTLURck0XImhYDF0a/1A6aALew7qnms5MTmQ5KGxfX+jrNH
cz2y2MFS0H8KanQ4P7oqG5CSQD2+UJjvqgGlYzWqT5p7yYqeS2/U7j47ln9VsTX6
C1Udb+Hub7oa4yU34LnmkzoYUKgn5FOn+LK6Mgq9kncyXZhjbbA7RqXodSKyF5yu
iL96gOnMYvi+yH6I4bDatjsoQGF7+VKOMWDJim8mRkivbwV7kW09CO+S2tTRljU4
fcSuL8DIUMKTFQeKOEeMTVkEwZngch1AGslnMKVGamdUpGtaDREMCyA/X+y1uQEc
7TNh3Pq04AFttqRpeKRqrM5qo/fzhORB6dshDTkv181n8UB5Vkw08ReAHz+Vtbdb
SKMrXXJkVBo06VkBVgIduW5yYchJLpBtCCoJEP6kBm8dROlwydh8DjpBS7vmy6Gd
1kTEvDsuTrgpydWxm34Z2MHHUKVvGQG7EjvpKLZ0NFrA6l2Ijs0Zx5gGBiQj/O6Q
SI3AwGAEln+RVhx06Us8YXAMLrYPsZ2sVnDQNGtYyxSQv0ZKp05lGeysmW+ZMfyO
OqiFCbG+Yynx5adntMFCJqgCDLoaBVe2UoJuHRCDnjRV2ede4Gm5hgAg9SBG3I8a
qZyOZyS75aA7i+ef5z0AQBgOSi1YoCB9CYHUMtCItberO0tm51v6uOB1POiKCxe0
F1WGJnSDHYBNpRFwtb0jmW8ipB/zBnrZcipSugWydLkxIRvNGf9LS9BwtW7uEMq+
OGWL8ILuSCGJ+fPtN5tLYb2uQsZSJYeAMmAbn/vZEejOS7zsfZDsN23pLCZEqjpS
hLq6GgMOnpscHyby9nN2GcojfUwv4OockEvohgKc87lbJdaKjUfObqoQY3B4T8ld
Njen2B3eaIbvNb/0fL0Q+sB22bCK/+EdDK7xwJSfRxWU8WbT+afp2emuQpS9HlPn
IeZG/+42oRyOsq4LIGG9Yjpdc8hKvsfYGT9B87CaaY5rXyY5xwHQ5EttJuOPwrlh
0gIq9FT30vA5YpUm4x7wTSA1JAOPAajNTMOFLwWAB0SMoZdDgJwPsVZasFRd+bY1
vhHayNbvk4/FRoPnS7r+QNdFQmiAfXnfmo9rgZUN6au5uPkSbRLGbpQwWuQNcDvJ
HyhvnfP9EZDM9LYo4s05CDz5NTbYSnVrxZzqrWE9Svl1qkUApy3Bb2Ydb4Px8tvs
/Ieh/Lj4YKR1Zd6k0SxILmgvCmdovoGw9fIzaRLxKF014YYfyc+3aG1c7xxN9ofs
uyFQ5kZoTgsxxqUVplkqSESOvwGcSLuNglDfhHjzLIX5dwL7p2qWuozkgoNZJJFD
lg6bblwYTCgasWpcbuP3D3KWbB3XF/SBwPj9lFdusi01/ceykvVGyStg+hSXHks8
acG5LLdaePG9VF6QFmYB4tWVKzeH5FXPZyTgnd5/PG6hARC7sx/WgI9o/Ic1fZk3
n/8/BB0tHKu1aiBc/+Rc6gcpaeYoxEp8YFoz2PjDn5F8fMgktw8zuDETOV8UNm7g
9hSgRe+ZS9oai2ygspj4bwXHeqW0aFdA5gQz+xIeSstey80l6HAoS3/pATqbsMX+
udiytAA62N8NhwKk4ldjSnkyUmoXsC8BwRQ2VKWVV1/uf1/jr+BMe+Pec0L5GUIq
4PZmiVQyPCDjxex4CJ0IFtJYjhDdOWPSJnmkxEhB9KHoMuUMTHfI+NHpqYu1UEUo
u9+cjCyO7kd8PItCg3r4VShI7+CE/Pp+dzKsvv34iVz7/MbEqS0CneK7tJ3IXAUS
a2fox8evXB86DLOOo8Ma4sIBlluQr+5X1mbG50R09ZLTTt7nLYsMy4U7ZSoIJvM7
kIdsuHWxh455QY0GRYfNm2JeNOqP0ttS2q8pkH7aEjOc6uMMuwPYuxzTGJDnQsIq
kw3ORBwN81L6GqbXQk2NtYnnhpbSkIAHCdLZS4zS6UgqRDGcZQP8tivukOkV6361
Ih22UgtvFoZW+2Y+vtT1CrfjXXsc4o/S94bPdfhBwx2O/2VnsDi6g2sXCurJrrbB
7wUWjQWr3AEJJwCX61FzWx22s/wwoiapFpMWXiZpZV9E7s5+nA5tSeFALfghZM3d
xtXcy4fLGGdABhHc5sSqW0BvE6Ddan9fR0JWtGTNav4eG9XkKW136HSZYBLoOti1
IGYl6ONudNTTuZCKPQ81Yso2039Fi6zPmNF7KxMQxKAKawYCWzIFjG6/mPlPRJZO
p8k0RDohvV5Iab8PIXOVLp0k5UdFim829zq/kA4B36DJAMkQJBL4sc38YPgxDnPh
UNK/0t34mnoO5gd+izP1Wnc3wlaXysM+C0aghs/hQgQGzPnTNo9UMPd/ab/qKeDB
XEUOwNbNiGIlmeqBzLxbWtuX+CtuKn+cVZ0vVSVgnuKcfwAa++kxEcJNf54BOhXt
UA98ezsBKJzoC+4j3OkB5DHH1pz4P+zdzUXfz57FU5h3z95A+HK+lvMK17PI5BFo
j3e7oNGnF/MP8fN5P2AgQFEyxorOWWUnak5eiXD3XMwL/WChiZV0FXGAaqjnXpUj
rsq3tRuym7RTSzd0FDoCdZ8xOpN2QINQr9jnPq0j3+vtJ/xssYA1bzQCh79v4V+N
U4flRuWxpqUF0MzouIFS8ly2+6M5DTUCS7QG+MlJU3aiIz5iEvDET4KVlqK5ec4j
fq/mfgslHQdfH/B3u/Jon2mTliqsMIsGECacR6e3VBbkKHVATe1CaTNs/O9mL8Wf
vDQFQKGJ9pa1h5fu2+Cm9bEfrpBq3z5MrD/O9uBLDa6LoFdELRJbyWuw+j+6fAPA
TkBXjYwNcpYNk+xBgktYLB0o/JScUrC+SKfTaekWrmfWhAjUXoOJr3M7KYoRiEZe
57mxpXuscbbog5TQsFJNBSOXKIvzxVfCfSBOk8xXK4X6TZzH3i/9a4dANezrBzp6
G+b1tj2Y8WbUT6mtijssb019JB8QmiHX3nsEq4Yijh4s+0wFwRmlxW6yaNN7WHj9
+N8ZzX43W8hQ3xCkvNhy+8+Bln2OGsXxPKC26RYQ+7bVh01oEdyko05yE3EAu/Os
NruZDYKrpoMoHCdfrkXsr4Xehf/30HWqNIoE6BsfQRxkDgzgIanNno4Mz+GWQ9ZQ
u7zLbmYMo4Q/xqr518OhGrJoqSWsekZJIH3ygAdoKRp14b7EFDopjuACyAbFfH08
5p7M/iM2dYVp27XR9lXSisgQe/MwoOqsm4mJCIVY5Eqh170jVL7x4M40Bx6vqmAf
zhZh7H6QqHyhcdmY/GyWiDlDY9HslKhs30gnEzhzSkAjHDLMuk4m66I94cOSUU8f
vv3SxlgyIRhQdIjLxmxhKjW7bAkIWTn2+bLrMgUcQwFTtG/1K/CRuUW3MXyzkdN/
dI5NvqWnwIV+7E9iqcBqNmcec6sjlWPYeQhMcR+GBHd6vFCtTIwb6SEntdk9t4fV
VW8aT4VIxZ8dNa//ti45DduOffcnSCd07gGS1Zqhc0DWBKP1Dtpen2w7dm7hkmTP
xOx/kKmLPku7t8I02WjMKYwdwp+dP1qBLu9DgtXveZm2byOfP0rKAN0avHon92tB
JK6nkTXUT45Y+OZcK4+sfznBDL+7AoZRlSHxZnteYtqWn/RhzhDUNddBuWCqmkVD
VSCMdzeZDE1jpO+jA2XYFKWNKE7xW/W8XF1bxqaA/VGHO16vqpu5eRjEHxDpWvAI
+X8CdxbiCYQpXISJbjb6MbMnjNLhpJC44FHSe5igonQ9u+vUoLZDWVGE5vjGUPnv
VTmkqn7BQDSBXMSlQjD5fCk2X4+vzOvGDcDH76wQMa1N7Y+BhoOHhS1uXY9WZ6nK
IhurAV5XrzRlofiTaECsj1R25eAtqGMppK93c6h8QrCQnr+K667Mkruy01YPv4v5
jPtW69LzDTIdjG6N7OzR7Fe9/AlYjM6nl9y20iIQi6FfeQfRQpLVW5PsatvbDeoS
SSevAkGdntCded2MuFOId2AoFrGxYN/Wp+Y6R5f98DaXiO6uxbz73MXpO3oqml9V
1H1eXCFpg4Qkn7aUH+8UImsffPAVbTgwQRzUZ/DmD08Vf+XCYcRIfY4IDZep8yaA
q3x0MnF6Njt6uuLbVChSApDVzyINJnUCtyDoaa6XARDjmGOZuO+8bjM4LJdf7gM5
gC9bjU4Hh7ciF+j2bY46L0R0Fcw8b1wCyLr1UGvEIzaiIX8WVcZCWeIzvtWXUcjN
KOd3ASWFzKwgnA2f+pSkyDDaNiMcQJyKvUgmzF9Vu4X38KUv1qyvwd39iDs/BaBF
bR0NILLCYNMPZbxUoukndUOnDv+ztcBzLNYdW06gnJPoES5lU26gCRm2gVddQU/u
pccVq5mj2XP+QfPQ6DviT/RSkA3Aeb2KNE442pEk5ENBznlQOZItAQXp6YnEJDsK
Rhmk4hFz16odlrT0Q3T0Mj6u8w+dbzGvlvc0IJ8t+RQX7kNTp2lWZBMTZJziMriQ
RovNvYaxUNwtvtvXK9uhgwsUsnH+BOW6DDHM318nI5mX1NMX9F6SS51B4NI+sg7k
xAtM3MrXfZsyiIs+RnT1LmcxjWo9fFFMyGHrPAg4ROwjpQZuDOaQ354fQci4XTlX
x85uqhzdR2iNNOGTNz6LM3scHGXGPcQktHHEnxe5uZOrOSW+wiyLr1WRJVzmLFjw
BK+9puJHN3uAb5nPUzpFDyh8Ua3sOIInzZbKUp/96KwtWRPPfLFVqKfQjNAnOseD
+49mBqSlpuM/rsJF/WZ/OxIgUkkSB7/RrSPsHibf5uGObaGoKsQn05dCN11Xp2T9
BtVrFIhdnyuXLf0KW9ZdRwzcuCAq9RdUcGAmcsGAgcVHVcJ142udBVtEH2X4/xO6
gShpdLd0Q6JWKWm0udo/AkNCIi478EyivDClUor4BiLiG2hATVCRIN6V0+xaJSgG
4FPoxrz8Fff3yBVrbkSc8JjWYbCwrmKizWQzAunPtKnYB2jQsrObskIsB47Vgy1H
8JwSR+oJ6ulQonRY2mla7MTd49eH1Gvb7Gcmvw6eXVFKh5drr12Se3LzOqt4C+pB
mNjP7ZnLpqPPAv5qEvUlWHe0cIwJSQ7VVxEkIaV+K4tSf9WdwYoReT1kx9Sh9Rsu
4BC4BfJdn4QON3JUFcVK11UQtT6w7UU02oNFx9yIf6cY8qaeeAnvWIZ3a+QvqQSS
HIWZNN5B/6216kd5KpxG1SBEjT0mqY1MnXvC7pbf67shmhtwcBK4yqT0kq3hU0Bb
PMkxyq37J7gIqHmixz/Su4XBViLExKMQhnVFZBrzboXNF6J/MV0lt/qV/IBFJogB
X3p/enY3e2l/P8FtSItsnwWp6VYNs7FvsasI3+eXB7Oj56LjRBlpZ01aMYctc2aR
4CMU1OfcSNLmB4I3htavEarkxvWMMy7kJOjacesOHCZkHx5lvvEcFTyOj0PvlwfI
Jfnq1hdShdQoEK68qQOipQWLVVF7Oz8r6vWLZ14icUeUs4+/fHvXPs1zTkZJyHbl
XaGgNqxNPvPKa+jHUFPcUEiFsT3WtI1xA2jJY68oGhHGVeH0sOTQhzkjIo8IivS2
Uflx/HXUoD9IS4xKpvPmKAH0MLSzPgsh22zIzJ9ui1QfmA/Y7nIeKxe75BxsIrgu
0SD7/61x0G85/jrI8vnclBRWMOf1M22h9rD6bQo717u8ebeJ7987hxP9dgZq4IGS
wfxeS3is0NTNvDosSJyAMUzo4mmyXXeAV/iAVEAvFUFqip8V/THtFsGQngErgpVx
kBJr7gZTwrBS0K2VFAqXRxiAZq3QwBYSu/+TaRqmYZ3DJWAUbIf1xc8jsrTSrgmi
m0vxwvuEuYJTlMeuYe3YWGgqU9DwLagKjiedN44MiUv6RUD2/w64bKNRjBCF53P4
93EGtt71ybCKJtoGA1X2+ggecbXwPowTVEt1I6FNuMDgJ2bG4mxObgIJfVfsjkxV
B1RBGytWct4k6vtwi5O7kK2Q92HhZFdYTRsslwjGBF4HLm1NnxN0+nHsVNMuesmC
FArvNWMbBeIFWKKADDJOoEE6QMRewirVzcbTl+k2R7WrIGFGTy0Iya6NDHVaLioN
DhsMedd3xLsuSdGFKonBDmu5e7Fi4DxGFeXG+gZsIDp/cES8UhfzcnTClVcohy+T
MevG8CSCDLoVgS11i/c4lClODWQp+kWv1SQmppYlLA4wH0YsglJJqzkWw3l2tNdp
BPgyjFOyB7/k1Ca5hmY1Tw50G1AIM9DZr3/cWKYO145uFHS+VDO68s5A9a+61ikx
BNjLGZuFHNaMdAXzQ41mEC/MIJE/HWzcpBg5Zu8GKgrBL4keh+faySIkVnpfM3HL
ZnfW2FPHwOBBsKqLDh7OCbpjvA5S+HgV9Sp/DKa0NTBsWmPmKXR5NLSitTxx9PHI
t/i+wNgeenjq4lTs1M3esD7KDbH5ut2a3Bp20uYLoEGfhkCMOuFENqOxE7NRty+b
Ank5YZP6vHI0wzm6Abh+2bKcBcpqX+6FEK0rDmszldY0Ngwh1eECrNXrvNC8IrWa
i17nGxABQQcDKBwZLMoROeWeSY5U8z+FmD8NnenOCcik27BzEtrAq50setdsdX6e
YFXDDNXZypgzCBJnEc6NBwNWCv2/2o1BNMCn90ARFP32KImZKp5OShrMNjyNLvgC
x4VK/2MrNBZ5kb1+oPSnneIwHBOD00zY5sfttzRvHYq/C2ELJPAZ1Gt42SKc66MI
q6b5YfuB9R7SLDP+3WeUZDhJAepXiU12wRTnC9Jq/hBpHn74ZE3BXl4aC9DMhK+f
dogQxHfNdhjobn5yjPm04qZtAhlxyGsIeaE7ks5YFMibWQ647r42iYQPw22PtjOE
LFlYtirBvG4K426GHHXoJ9ktbPzkquz90QBLdwvBZ8+hC8H+bf8uebxE4dXnwTBd
WzR5lNB41qE8Haa5n/8rR6dd3ZVrHrzTIqDGURpCbjrGIuchbAzGkrfFh0UDqpT0
cVN4QlMCS0jToEdiJ3vUKd5Zqo/5cVVs9wFnXH4NVHo/r8jTokeGu+ExmWc1SGkq
qAik8wgvL0FHlrKv2K5hJ1uxIjYkU1OcSyZvp3s5HqXQV2MilZipyVqdYIiWRlTU
dYvN8kcfGzDv4H0NkPT4DNzjF1RUmf2dVeru2GpjKc275zcUgYXb+pxsipFFE19t
iOLofUMujAx0Q/E8OxREp5kZEqx8Ny1In4lVWHzswkWEAPe91p5UgOa9GhBwFYWA
7e5m8jjBt/o0aGzFLvSV6mdqMzFX8Gh4dx/2H6OI153o1Dl8GADlvwyx/5oEiyYW
blpkQeGxXeOaBm7dHYkfIOVJCSqX7zBv66JXdb6KQ0md9xyWmKJSAT6mE9BoB4gw
VWdclAO1Yz4a4SepmWu1LUOH4S+t81RVVDxV/Xj2BrvXwlKRgCcKUxtTcQ2r5h0R
Gu9RzFbZjd+Tq1oX8eFcf6++Nsgm+gQ2IHqt8Rbi1ZmVC2Qi0p0vxLNPmgFpLMvR
8DKUJh0bq4hYQ5wYo1mkOc1oZW0xn/l7n5E+XL7kBJMPbO49RqUgCbHebUO+eJQi
SHsgmKaafZxFmNXp3wo6THUIRW3kJkWG4ectpNnTHSjSROaPtRqdSYfQJNfqlGV4
ArNTsHuinlL8lwF1QcGzmRpUURmH3uCjyFhiI0LWQkLXoV8SOYnyVk9tswOk67G8
Q8pkhOJhcxVEGvX8g02aPd9p5XQ7C2YDqBphla6zF3veSJraEi+C/BmpTgp2ejY0
7oWKB8zuILXsGBvEqYDd73H2Yko/odUFnBkKZwjBx30aT7MKMJ9ajN9LK79Dg8tl
pscYuXSScPeK7VNA2NoxhHjf6v1tHE2EscaUBThjzsFrnVQY82azHtdNueeD2VRP
LOMqUizLs7ouD5Z0jhhQ3A4kwNJp2BqU6z3bD8eA7Av/DjnvuCGaxQhJsuMrkr4A
w/fdb7chJ60fmr/i9U5B+KOseEZt+RAYQeTlttIxasD0T1CNtmH0xiXEBUxM36ST
OdPNYkNMrVqW0Lr+RP/I148Cs8Z0dQ7fs7jxMkYimpsa19fU6dA39ONLuGuqjeiI
N98xDaqb8q8UOAvT7S5/7nDr/7iMNbxUhVsKAszOA8OI9dp5QLw3mvTduca++9+Y
xaifzEhxhTl3JpV8gGOIJm6Tit72Z+UActW3x4QKU/9lfIjs+BziKIFYz/2c7bxS
wBV/VDv5yeY5tot/IJrFfeopKojwZJ7w3BKcWWXMGdX3PmtAiewUYkvUTxKD1iMb
qXyob8y2b9h4ycv7yhaE+Ay93KZXOV+gwjfGf/DwqM1JFpw4DnrGrB/ttmpvalct
7/jdghCY9capyJYlHQRsn3hCvdiIK1TMPyUTfWWa6V1B+n74pZOL/2Ud53SDSTFx
o9+EvfaYzVXIn5HtVjrFUOCLOkY3Z0mXXDPvwY3Lt9W+fBHydx9DSCMNld6aAmPj
B0IMQ8j+KeAV/W3ZMPCS9faJOVDdOXDzIDbXeUB100P2CdJgzIlfE+D2ypl752f8
nNS76vqImD4j5HQBM8EfKp+wDXbi/wXJ/nBrsoPiI3OoUysFpquxcEfOCtT+UIpZ
O8vz7/SX5hpx4Y+kiOiFZtB81nxyBpNg4dbCnNWJsYsGlaVXHy4eg8QhXomUt78P
sj1kp6KcYSWJp9IMmGfYxCos6z37jyI3dH/zc9h7qMnMyVje+FUVl6KnCeULIPGH
H/YUt72KNVMIY3GfGrpxPBPwpsR/6/ycc3Ku2oFkOQ0SznEbqPMXxKSjpxW7bgRj
ziSJqvecAJunUT1k6XqA/BGlhPwRlKkNh3esu0ooJLbvt1zjneR/nBALmHB/TZK1
Cc2UwwTKIGi6NqLlw9mG75ItO35mA361E3WoOZ3aFUG/Vtz/If0hdGF1Pv5F8Vbg
60ctUwhoZdVDtfAC3Rioeya14XKjuN7ok1K32o+2iSKxGuRYJ0arMCzbRokCA6XO
BEoRIii/qF3glD82GlYLEIArMzeX80sm56Ptcqy6d4+Y1g2Bn1oeCbeQFtNqQJyV
fcqkxjKUQ3BGH62poXVIBZYtRnra8pG1spZDJVr7v0ukLJTfugdCX69C2ktccG8e
HVrd9k5QVhViqTnMMtEPhHljpsyMNOPaLs9oJ5Q5yNn1SR8kv9GcMlE1J/2qolki
XPuFLNXs3aBHsu5+CLSUVTVV0AiCS96kiGZg6c1SBNFJJJwLSeaaA1xsyq9U8m4v
WUM5hnneF3kLdENbcV76ZMcOnsed6n6AzRM6DdHKhZtXDPod3n49uFovoKmOMJwq
J03biLy9INuGlOWchRH7/8hBPsxJ2dmOh+YQBPhf65ytLEolwEvyl+6S06X9InP7
z1Bc1siTDF8Rpv+CLUqOmr13IU/pN6jbuc+Xwe1T69qLKkYH35q6td93y1zaj7LB
2HfS//NNHP69rq+6cRebK91X8MjaK1RzY4QNGwFKGaiuvvny7U79kesDnoTGgFEd
kZEo7zt6ylhtv/bZH5vORyyyT/bvz5NhRmcELwtxC1D1FGfoMRJg/QefW0iou28P
rEpMAL3ikjJahqnIsC8GJNF7cy55cSrCCqct0nPb+dD2fe30Uz0NB2OWLil6HQx3
h5l2zh6yuDluJkjesu+T0Wd0vH3syenoEtdNpZiCHL9kzlgkMcekPQaGqhBaLPvP
D69sHUD3CBsEVMn+HCEwjddGx62/7oZecFfVqWGGGhOJQwAa0XbYqpQJ2QCBZBUH
M61I9em+1sIytDPt0CV9tipOSw0KhnWqrBA/Lw4f+y/nwFNiVW5Cfi0oqegPLPhR
1P4sHPwFPHjUrR0jfSj3gz2hTsQnW51btWD7V5J9EnpHq7nvs5Rz2Xg2Nga3PrWL
e13V4fyZmBD8kI0HqoYiXKvf4gcOvhI0ZwsVnXCwOM6iqy9G7eF6tZRmsEpA29F+
TteVfIviySn5KiGaI7BC68o9y3dgKOcQlyULgAHJ1c3y/DFZLhZ0pcVHn+PoJ3LL
vv694OShT3GMRFJbJIBQamZ/nIsu0htk92gpB0JAP6daHiPnWaR6ngyXxIqexJtK
lT1GXPIhRbqtKVqmcO0o0Ydq+RHTZ9kLpgQYxfFwXLz71IdD63ulHGL/Englsqgv
n22zQOwXM0nhJeDgH2OhS8ECfxOKopU/630TQHFd3WN1+oATSXttn517tnIsKF/M
wiGrlkZN2GUZW8a5o4v/uvYcBgdG10QB/5dU9sdhnxUcs2V69sa/pWR0rkyR0zp2
90xf9tn/h3H6dX0ANMOVF6oOrdckdHw+8+DgA4pBd4S1SExNlOkSn9FoyDmK3FyL
Ubt7RjgvDzNF1YMNnvY3f8/q6VozH6CMzWbThzbOQoAcImJwJFwFb8ssNzMA8A3A
d2HHkM9Gy0OKxfzD7XBC+oORz1yUfX5j1BNhJhtWi2oAbfQrQMFfZwDOcE+JLckU
TXrJiIlU4nK4v/429+Kygl4aBIiGv2vAfESytm66vPF1ROMjIzgKL7YP+SmaQcJ3
aai3qj6S3P7JONKNE3NsB18ZLBLGH9z0+XF428mkQdpXkMLTNurMKp/dDPVjaIuD
3ocUedSqOcGqjiXNpAEpq3sGqNvC/s+mdh8ZuJgqe0zh4yaTfbzrmlkU+nQZltMv
M5Zz2F9SA5DNcxlOeSC0GlU7Ti/RTDX1glFPWE5KJPm7FH4Ihu4/tttF5lPkDbAj
kTwhJfd+d+QNDbc4LX0NaBzNRN8hZrSp5vQaynMrkBA7FEdwkAFuw2oSNCvBD69y
Y38cbxKy3/RNfk1dTkU/tp86MLKUxIzPcOa4wzCWgZuUPoPJF6eFO5kVnCR+r9WD
5Q3KfvsOh+4BJ1ed+fNBVwe1bbs7ilWKIdEPVxESONo+IirS1EfjNb6NaM6Tpt5t
DuRJS9s0bvFPAQ9aJxo5iZUk3Rb+pGr+sFiSqoxx4UaC+dwuUZ4u6FnSkL+qZgI0
D38DwDJKXbaUsVZO4hadgVf1hpAeopo6kSQMB7SZENJbbvf60hGj1gjHeFXrYyUJ
c50LSuahitvvbIwJsJyOVZGhI1E9ukYOkcCnxauoheRdTBN0yGKAqM0DxQtbu5LC
0ZfyoMiqMJPfunr7SF8IwH7ewMdf5uTcQS0sYqgbXofSEojyYN5Kk7UYSuSGmLHE
0wv52Sw1gCHyx3wJeg3qlU818lsYs5DFkdonsQsiNIM25t0hvIMgQ1w8BFfo0n61
seQ70hs1MM+w3cfx+02ShSrJupjw4aUH1scG2p17NBcG+k5YBiW3jhqG1Vpm71PG
USLjQxQAvNAPo/dhiqS4eexrmlthmsnh1jr1BSrJVfLY2XwnzuO/nl/IhOOLt9EN
ltfjUXhmje2+84gX5jsDLb550FPgwNZ+GKbeF6ASGAiprr1RUIdFsjQlMRGYJWkG
eeUCw6/03ht6f2hiFmcfpfKhegAEi2LmBA8TmvkFICQ9bstoWB/mV0mIC9ObR1oj
WUky4+n/M3U5lW37UlIfHVSs3WAS2iju7HR9vLQ2C7DwE5Dl8w+qCi8X9cKLWc6O
JNgYkU+YlA1p6g6h6zI5EIeFgSCl0j9uNmevy6sefa3Z5+wUpLlzN2/dI7vMgP/m
UsB+5P8i8xkN4G6L3an1gfPYk0EA22qI9tbJpkyneX+SvegA285CjwrxQfFdULzo
nrV3ou+F0zA1ZFlDkQLYUBDgC1SCIcCwSJYZlgK2o+gJIu2AJ6cUGioeVo9XyOWf
FJ74BLr81DHlHDPr4BVJ+3u8BfAswNFvKBbIIwy7EuDlj6fkK+10tbTQSmXWC/u8
LGNo2ze8997jh6sRK7cCvHMVjQZAowVKU4EYDKjWcyvIXP/P1raJ40SA5qQTp2pR
n4GQDl5BiltISXt8tuK9x3MyIRwrvTFj6T2KNgA7Q/I4jXEr5NM5Kh+dhXFuvzib
H9s0btdyO/NLlsy8k+OSu3VJrsJOCv63IqpquuxfQyLfrbk89s8/J4g3J/C5ZNjz
5qFYikzJJkXAZzJedcc1lk6ZP4vL+fjxs/V6K/ZeA+0AXQRTCotARQvB61CbGt7M
FyRUfcUyGy3r8RMyxA/eut+1O+2XE5veN7xna1CafMz1qyq8kkOcyZbX31wQBLm/
Wf5rYxZpO+0VejJJ9madFJvwssqmp3v8H5VsO7LeKl/TfQ2mJxuFviANjFzxG9JC
LmTBLiVNopi/hVY7jhl8tI7ufVFyCNUjJBqy0vOUlxUJSc2pGp/aCBkTjNTuUpT6
14NAN7E84emxW1MApIQfU9gG9vQS5l36oIJp2Fkd9eiG/kPCMfmQDyzc+baCHIN/
C/FfYCqanlZTeA/hIL5vueutXJGddpUA+7+xONtWNjqHS8LN/2GjRKRUpE/qQDzi
tDBUdjonuYAW3DBSNEAl9//42qWiYRukXzM0x4jfv8r0ap7xcrR77tHaav2HW7G7
nGKHKU+n+OQkeAG2oB49Qqx/pdMcEvEZzktrd4QkohmzgPeJYe7NZKB2FooL5vEG
FDFalAoyr4awH3lmdbPG0a0Z2KjsWE+Jz7C6QWFBkTlFcP0vbKbdfGmePHh3ZYu2
DeFbIKuEMzLf/e5vfaRN1Mke7njNTGz0qq06bsi0qSZnh/TVw/8rKbUEftw7jEXX
C3y/ct6KTMOuqNGVav04FlSh4XnQdhmhBvm0ycvDBdkzSafhuqliLOpJnQ3Pct69
p1ucJW4F1qqtCOGWWot3Mhl9YI/5gxUGppEaLjFOck1Q0bQkefPvJCr/bjjk6GXd
x0KF98ckgncNkX2mseR2nAwjvXrtQfKin3OQuOs1s2r5D52FBjubtTk2STQqasij
tPctI0iAg5gjmCkc/5FW8xiXCzQj6xAAi08yrH+UOce4/EZIb8IKIIBVz/8rC/ht
L1FTM2j2T537VmmsLjS6rp1sfqFBT8i5mwDNlrjBOTrxoeUzKuqDHh7YqwoSxvg2
xEy+6GJ9/2he7iO9HHFOV50BLzgEv8SQb6JPa1AhBTXwvHNENNjhg1GDXq9gnH91
WCCDl8K/kY6dzSvs/jRgdSW6LoOkCxeWspLME6FpIAZr8ILgEs6Xsghb52U/uJIM
VW18zpb9Rbl2R1xjlR3rtTxaEqlsKBjAAckVbefJ176cBATfNuhlO+6z5FdoZLUb
4n7Oq5Zx7QuoPtd7+v3VMO3aCGsCmK+oryKmN8+ud8x9+qD7WD5ylo/96uLMV8o2
eqEQ1VGxOYNT4Ie4PtuiYem+sv/98DKPGkHINn0krpFKoTS/Z5DkSIh/bKvt80Vy
IXbFRks+hm2l5SMB0/hNMRvkQfqT3P1KX8xmWUDhOakG4YTLwhZZQaTR+FKPaPm7
lU3cniGyYPKNnsjIN0KGMuGz8xwACpfuEc1xe3JJddJbG2SLeFfHM2A/TVB1UZTi
ouWmR0y4zB/NoggiiWscd4v7EKtkc0egWafzG9vXgGMB453yGRiZ4rIzOgrHvZ3u
DLN9f/1TC12IHSWSh+dCbgKNk3iS95qC81aSFXxgxW3B5IbbDtTrvrq62qqhYMGR
0KjXuPRTSJnnEASIkAKhROVWzFz0pRpX58STPTiwo5RUgoAoxg1l+vIB+ArLmfsK
Laff8tfDXadPzePZPvVaremU1i7NsBHZ8AwXx1V3IV1lwL2AjmsHthlU9AfWa3Tg
j/TnlVPM+emmyKaxFrdYujv91JPj/H9Vc4t8tCGhLdiEyw1iYaKZRuyzc110A5HR
4uoN283IjQn6LBt0/OTPtsEUGDkK9dnpOHz4Oav5DtY7ISrHBI5Cwv2Oa4l29R3E
2bp3lwWnEXn3RrhR1eO5Dvs5J/4fRZG8uRdvdfPPNZ4c20aJVy4ybxDCoQjHXW8b
WqnmYmkJRVja1yqhkhJqgFrGe7kdeH2Sc1Rn0TywtxUNGnA4mhiCokNU5OQ1clPN
KB/jgI+7cR3I7oIS4Ea5y65QeTvYGdKSsAAX57aB7JZQXs99v+BBuOyXKcN+lc8g
BxAb2v5Lm9FdX1Ff3vlGE3rDOvxvoZM1AlLvZWfXnsgg0C1LMgSarQcigckLzObF
44tE9Py63wekJUGM5ehlLstrz2tI52l7dU0ADPT6MWnEP0qdbPz3F3TykH0+SI9E
Hry8OvrHNMkZe33jb4ntUO0V9J2t+0JWoT8IVRw1xlKkVzww5HcI4cMG7c9WQZAv
gpHMETupfgoEEn9ZJsmbBCdJXRs0vAyRPyxT5NsukQYayANKk+yU/OqFV1/aEpLP
Z70Qrz2NyLwTDpQfbJap8vnksBTzIjYkpxp+GX1QzWWKgsqpRFjevL5Ijixr8Q/d
fRzo2pwXupra1mKoHtwtdFtuDaqIwSXkAtW6jeis+XULvTTqF90A6LztsZ2wsySH
t1CIGTrzYaVy6VhPoytKpGVK9nd8m1W/2hJ2VKvRcXmknyzDTv/7MoCL6x4AsMEd
dRvfBDRKxKtp9LRHeS5RM5YbjKxyoX9fcw52kl/seIxlsZokELpD90WxL2T5c3xP
gyXFCUbfWoBH/RXk9wQBJL3OIbozRyN8wKNedGZUu986l4sbaSzDajgsj0NYSS+y
E2uAedbrtZuw8Z95GWIzUyaZvwYdxyXgs0+Qbn10tfdSU1+gLtTbu/zHlEqrEGBf
86F8osFQ5C1074LsfEUktRfg+jeb6+1PT4SFTr5aRmLWHJoBMMORnddIyIkgUtnb
polUSYJfylh81qc4fxFj3x0U3k3qQsd5GLUVkg8AdHrRqqmHLLtFPuR5lZPX7tBg
Vu/5DKoI+Qs5OELdu2SaPQXsJF6gwWziQ1omS7u8Tgkt5aX0NtNefIL2MgaHwQ6J
Hi+Eo8YJbJtrDiOp+/rpUeFaCyV/bzAAOvCRGIt/w5YhjIMAj9LdHcxpVZDjeuho
3B6TGl7c22PJtRonYP+FBsBweNMYKMNJgHJeBZUzSKKPd+kLUGidAt2Uk0MbdhDo
huy0jyaXdQNlEbEsZq9p/LH3WZrC4TFRL8Ir3miMh5j5e+BD+kWFmz/S2WH3Gbl4
hZWtLMFKAl6ZTzVVkAAAOUBTu/C4BV2UZVx/nGkDCDLEjch+f+E7nwQKbuRuwYM+
AH3Nxt/8TCpxmSQxD6RJvHT5AEuu4jqnVpJuK9oV/vTLa5APvoEWGq3fqu6IXUiS
E+7wnZtfS+oL8wyBHmE/a/aLSJwCoML2I21Z+iWqRf6ztsP4kgC9RRRIkBnB6Hsu
QwhCo6Jl1xhjqj2Smmd6ThlTyIXKDCD8hi1Lt8IMD216rSTTgJiRdaBaiHLaDf1q
TsFve1I5/9At5j5+TD8zo5mU3JX38nokIgPz6I3EOFhtWPf1mqoWhnk+BvmD7pNr
ya6ckX4xE39n1Rs6hxxX6uFDCSOOFCtaPeuUsP6PTna28zjKI6a4b89jpN+DrOfQ
rPiGgOR2teMVVsoY8bSFwgNxflC7qu0A+cf97xyshUKHbkotdA/SXpzG1+THXWuX
71iYamzwqAuOHkQeXR3jrnkaRuWAoQKaFigldJgA7huPefibbDyzlITqlLVWWqLy
MKMl2UetkVE6ETR0DmALq3yTN8QAvzZU/kSKbzLaBbhvP7zx0KnA0D4Gk00lYfy3
iCg262J6yOw4sZDPWZpiRvuZ7+bGlZ3dQf6gC1xIT93p8EnE9cKCtGIml/IIia9+
nmdDEoCAcvW2LbZ9+LhZa7vJqFa8knN107k2zr38FuwgTTsjuKESlqxahe//Mxae
aeVgOla8tFWifnuTx+0/QhjGrn4rxcO9NQj1lxbOkhHdZtYwS2W4E5rur7mIIQVB
Jn+blDVU2tRGCpbPVUS5LC7y7hcXest29F4PacTffrMM6CazWfHvbBsh1/fNWcD5
pY4FO7nlPEuv0P9iJ4pJjDAbwaledy3Rlr07XACuh+ZMaGkCnZ6dyRDlCkwytu/h
1WC0LnyE1vr3QGd2jmBHP5kq1eiTIGAq5m8uRBiadGd/xZkWIcq7TzKWZgvQxSOv
F6hGcQT8XDgyu6ElJ7xSse4Pj7LvSn35p0e6reHfcayh1iEAwAyLodqL5bqvgiaw
t+GT3caqoSADdwKD+c4YCnfckmqECi/8g3m0hbq7VWHH058ugtNdMOU033aRGgXC
E8Wqbx6+2QsR/7o35QZPyiNgnqDERsd64UJdb/N3Ay87YIvGbUmBJT4i8X6duSTQ
FVhQLg1ItccInzfAuNWOwL3HoXaLO/yLhrZVgP3jqgfIGLUvbbofWbjFIMqjiqeW
ZonlcoizqR4eNg8yWig9lWJAFWoRk9uwDmkDJyuMLxS2wirbniJGBwt2Awkn6h0S
8oPFB+QXsLBMJI6oQRv3whtsxzheugnYB1oqMKqtSwfwV1jTFmrZAlYkii3EZ6C9
vT6hYVjLe1l+ttFqgFs/H+GS4GbNxZYb+0oGoHCFCL9f867UlBW73xVxLvihuchl
KeUQRXiDFihaTOmBYx1R8cPots7fKD0faWOFOkouu9m9iFKDYe7TW9BqV7e9IXmP
b03ZSZLjzpCh6pHcz4Zn47vwZ86GiinmTHyhHZXYQuRZKnDBScSRISiFNA3CrcJh
GAns0UgNAmlb+iIKSfssMOiyb/vXyus5VHEo1SagSvWy59KmYxOwymc+W9j1GUUD
oZEHutcbi5UHMIk9Wlv2HMDFW0LQb6iCW/8uR+bWfGbLoFD3nYa7jYwcPbCIv1C+
1DnH8B17LlMVlObwpSQyZHAwuAn2HOUgbl+URpUnVXo3Lu5uHRzY/mekEQWJecn4
hlvp3rwo00Yjnp4zSAGDXopWq+/IoHeqDxSSSq2O2jp2T3bfditefjbc5HZJG5+J
G0iqlxlSECv64vNQjCfI47TS0eaOvlJoCFOnozHPpBjFMEm5yw1PkSr3GaXQiEB2
GgxLHaICXZz/sl+YtLjeVYt0desKVQlHvKwgzp+Iczgie22hYZXimMCiek6TUW76
3PTnBJGAllLDttn6oX+oCqbdOtylczCU+Zje/Hwy0Yu2M59NbMi2F79oBl49flnL
oITenPUJ266kPXORO5KZPa8O9xGx/facYVziRCXTU1Yc0S3jzcP2+frOaDAIokeb
h70gnEp+C1eGo3dj/MKq1D5+2vgRikr/zsUk/kBti2HHdfJer2SBU1GZsleyb+bR
/EREW6+1clqkYuxPyC6+wGPOlcmwYNTrWXowhRXTxRTVsW65K1iQc3FNyWPpvmRO
L2Q07APJGDb+XNCZBBXjHmKFNwa6nptWltFCC9A/F1uJU5oPf2Bd+/ket+/IjpOo
fDrstRLaweL9i/c3txu020tCCZBzpJfusqNRWOzjhPzGKe7RR8CZRIXL4oxDrjTD
lOwbwZgZVoNJWC1a88YKrCwKDzir7x6VWPtgVOIvYVWjtH5NoHNX377a1XgLwGgD
NhuQrsgXgo7CP8Cir4cXATTPRLJuAEVuulvS9zQPloYkuan52/fALRnn9O+OouNv
6z5OnnDFkTgOW9dnfWocHYA3gJmLan65fz4U/XQVY+Yxo/+VY8l26/qKwSi0Oj+h
/Mug8BbecbHA7DbgrhE5nr1fsMsI0sRlmD5RTPIdmKyueG7+4GOFwUUDiJVWhIfB
xTPM6zoHDzmSdXnTeEwCaDNzfLangtQOfvyrDcLzW6DOsHNUrGGeNxFrRLqi4raR
pNxF6iZUSPUjtMRINj9POdcWJft90W/vHGO2folxgqRD67EIjYB/j263TZdRMkoM
YvuaCHhEYUBO53iZ2tqAZA3Ri8WMlF/wFcr2tBhYHAAWdqORW86uX1KZdmlTUmDR
CSyhgrzBAggFjam3WjdKbqm9cZrBUopLcPVGjJ1PA2q++t1bZIwq4nqDKKNhisH5
JtFW1BY7Z4hRQjuO4hUjRdbs67D/CXBkqc/f0Vz6pribRbgY7dlDIaQ1kKH1FrSC
0Im5QkgB7Sg1cNoeywkWHw7BAjQmhmvbxGyaGWkYFpwMPqbsiAMhK0RV6+MiCunO
iXgp4jGjiZvQ74OyWuYwJdSXwPdV/PO1TDFdmPq7Yh2E036LVbwTSH6HYhevxQRI
DwC+fbCN66y18uzV4pVrduFdc8iomu8nYPIGlU+p1QYQT3S9Un+y6UkqQKsS72x7
kOCwlRdQ5H9uG+r2QuYyNFCRwa3uUi81a/2WqbFR3n4MJq146UdoPSGMPEXpfUyi
QToLQ7Btp8WNn+X5B+Nx0oqasenqPafwEJX1DT3b3QY94GIja3F+1SNtQoIjXsVY
Bj3Gh7JFGn4akePzSbjtZ0fhqwVQU0ElCYZ0qbWeTn7KGiHoGu+zCRR+KbYuiruY
y63/W2fkLGrPRz+VMhOF/nPj/nqRfTcpsGRN0+dQWzu830bBeu1fYJMc8Mz0JQ+k
Zge4cwa7VcdviDfjo9+CP++qgk12QuIqal+HvZNmrVAmbEX0tY5OKyQ6WuIvz8p8
WLXHT4TG0H1mk3CGEIlE4fw09iq/poonh95H+ppMQhYToflQnU1ATsXMwxftLluU
zarPxLuvaqlq1Ms9/mRw6LfJNyYKvW77oD5ZPpsvSgpQ2UHzQ5KvtYHltxOW0ixv
YZRYcjmRm1t0xVbFzxclluLx/DHe2x+qLhY9oRHBEl0nPIf7smIg97AaIbaXgSZj
qBxIyokLkZI6pvcWK03kkZOt0AFYQjQ35wBVY4iy/LONMEltIru3mlI1SF5XQptC
D0mLYv8sIyZI5T+lSC+Q/5g/C/+01yhpPwx3udnLgb5gVZlDAIwU+N9/g74oN9LU
JDQp29UPmn/JGpPbFVDUqoWSVyG7m72lSBTHDfUWubwbqzXwP18hYaIe0NK9bLH7
rpM7kwx6nRUxZPvlcnrUq480D20RLTnDKTy+CMEY7g7vrRom9HvDJrD5tzCw0CLW
LHvQoYtSNHbJG/7I2pIxAISs256GvYCN1eDMpxLjh9FvZH+KMCevT2eQlI/vU0F1
vV/jb2Gu6YB/+zT/LaQSBOeTuITbZtSumisAquTjHRCeTfCVkLsgTpVHpjXtAfEw
uT7a/TsEuUCIk0OXJvJ4oCEP1ooXiAHB3lwvsNGpLyW6Xad7BDFgVCOvJKa38V8t
puEvpj3B5HWscfvDqOdfpKzAnxdUsDOWKWOKu2P3m2n0nsYTKM4iSP2KTUAqo568
PeDK4NqdfiENwYRDuCjEQMA/R/ON/eCOJTUidiVG+0GQ/8T7h3gKG1rpHjJRwx+Y
SmbK64EhiFTFe5iCV1qAHO1qYSSNwOwsqmLHMRAWlnCCKTp77mwwY0vIyt/8u365
UYoQhxd29DbLbq2gjQmkeX4n/PFUh10S71WYd1k+yv21b1q33Pp7nJleD1vX1EGG
oLlfVteeraCU1bFo2CqMiIQJgxKtmLXkOkP5y4lSdQivUCyPA2qDblWZRcFMbuq4
LLD4pYSFOZ6qENJUBwunt9l2/ZsjA89+jcX1pjFkpvoz9cQCwBnPrI5y3EE3bEc8
/1CTu34yMPDO/om69ymNFE5+Ivd3+PCGu8qLmxdLmKfsKdP/2sWzdCBTGbiq91fg
OIYZ6O9Gkpas9J0USEUvgeqLbYCDia/EnU0W/6r0iOxb2eW/lCg4KhbkaRjpPpcq
hmxlVFyntfcAvFS6M5ikVVPmotrck15/Q16ufdxeKj1gMPajAWQIpCReuasyPiXE
Uecb+ezMYUTgVpsclFc/KHD6XKKUfGtR9xLuME0kDxNaZJlvwZynWbqY32MzRuhu
pAMwsVLGOX4zdoIuaNNxwXay2+KvDSpEAiKzGJoykytOrNycIccNObue7yu7DCJ0
C08HtqQh+HNJR3iI2aGZkowckv520Njs+Kl/Cor/kax8hETyq3nE+MzUBN8lD9bu
I1okz+0O+AHTzF1TjD6ZJ42CCQkHMWE4CYdDYIuXN5wwVKlIFNwT2wuME/42nfpF
wKc9P06sZvGlSE0+J8rshp9JoIgAw8A7z1z/i8za1hfG9706ozCIHZKovhblnQ74
KYzrZ5Zkf2bs8kaWs/Glkb8Nm5PyGbeZei/EClS+VrWxvD18UM3G5k/P3loRYFNU
9U1mwOwQUw0vpV+/jTvHE81M0JJxWxgPOBQ6k9MUCDpyzw/JOmG+iBKQ17luMi5n
vJEM2yZaCIWI+jOePxP4CwDN6hNFvTGctVtkNXwdcGSMtuh/H0ex9IU0f3nagXDC
tNhGb8fufiYrmSWB5MN4RJzygstpfRsU9gqcYtvHqUBCPj3g14cA1ILfwZ19bFEl
VGOL4v9UXb5Qd/b79aEHEOaktdjnkzoPx6f3kgMjWT3xVD4B6uuiy8IVe7fQozZ2
q2QC/RKfWIRHsNokJfKVGLpKejgUwc0XUUZ48bzEKH3a+uIIzaPfSVxqt6qP2viD
GpjLAqhTqb+X5ytE96QTkJjah7OP0/ABITnwz+UI9oE54Vts/q4lOGyhdVz6H5zJ
I41E2FpSOxCMuaVFAQOYlr3YxgZWE4JqgLKwtRTxmFwE7Ir5F0U1yt6TKnE/AJPF
DymtCRpzLLA2RtK6Fvt8dvdTwZ5LuRPal3LZCY9J4tOfxgRR16AlwF6NNCGVG+J9
ebbREv8nM5eSMVfct2fxSj25b9QTM2cDwxZbwmsgAEOQoBxszvzvNNN1mC6BJeHe
k7b/8arZLzj+CDSyBdZUURvfnrVLDSa/3vBxPKbjcez50pG5mnS+PShIGAjR2NgJ
AjQSjiuVvM/ol0iOv0MK+fgtLc/NArGCV1jbNLi3Fw6hKtpgIxmuvNQlnL3lRmV8
LGzyW9huIcy229bkWAa2koI7vvJ4rEViYKcyNXIu1zFuc+RwyY2lnKvwDuunljXE
nskOmr6ybR2jv4gxAIiHcrRUdZrPW1bzLj1F8/Q/E3oM3tLmRJ5PpFTCHtSA1cze
eMyZCFd7NI7+ZOhJ38mUX5pjqb4IbPrJbzHK97Fp137gSO6Wiz10dBXn1q1A3WHG
ahKcsfUS1Ht65ec9tFmt9uar7tkM7ahfvKPzAz3AOwFFIcVBH6HoyvoPV4796tXS
skKSP+cGJpBdnUfvLluiH6NLKgQS+Uw0GWG/l41a2RUIml/4p2nE7Fh+yqkSXgv3
1mBHR9c+v23NikLjFbqdpjX4U53qzKIvY5eb8/uXw7hWLJ2dkexPhs/4L0kxkoWd
EfgfT1r4DaNzIvdOFNK3Gd60IaGbz5pvBEuiwbULNONoVYM7nl5Ca6DZEC9qoSfq
EMsRRrulg0eiKN/ejKbYRCdupf7hCXw5HZ/XUve4u9cC0NvbK8gdOe2QVt+Z76e8
Cs/4mOGEC+GVxbd6yulf2ErhKJGY+DvA8pUm9JnEKo+sL70O6ChmSkbT7/fU19iV
RINzJn5/LRDwYdPM7iZRXncGp7DqAF2dJFtimOB2iKOv5cBJYBOG4QDFolf3FeUZ
0QMB9ltQqFrUB6KEdG6XLD4c7zwyhpwX1/OqGcTSf7H7GhC8lWKJDM5IyCOaMAsn
PoY7xP5BrOCedSsm9b1ycA1irhB64AzGNn11AdTvvdhIphkxqPMVF/LtJu2AXaMt
JH/8Fp00QdElDWDuB0xaCyXFw5DS3Pw0o5ZjUFy0GzqCch7/bbvIU/UIbNnScLuO
gm1fTPvWufern8cMvcEQyNsRTQQeTWEbfHkWlj9PyUmmLgtwVUr8JDp6Avj7JMMD
f4V5QOwwYAVPOCKWnDG4eULS8+T+BcKiGGjsAvbm9P3ZlWQggjDi2sV7GU0mrhSl
f0lsNUYHoM8ZeoZtJDUigYqJERGaBp0Hl91sCeYcxv/xFYHfEvg20B1yrJbJ70Dv
Ce5gNQ4q6VjsRYtRwD+oxjbGo4MQncItpyPAZUV+9jaKZQej/jQIRG6oLsji0pLJ
CaTnLY+2BqpFflZm2oj6Lwn4S7DnwPa/WzJ+A53nseOufyDzX2iM8X2SWLoFg8oS
NmF6XVmYy9OIYPPuW81eW8iNU+PWHdcJqd/jZP4WPpY9i5tAq/sd5AQ0QIvToQpw
ys9C7MJF1JJyqGky4CqwvThHv8pIrMXqI5nDMDA3KlGcECK6jvbjOKiuhy30lmFQ
feyEYHdigKjj6Xz1MzXynngHJkeo0L3URknN6i93+/QXCEVTyw08G6nm5PrPNu6V
B1tuQcW3dIuKD14X+8n7Di9Ww67nmvy5p3rMB4ajLwmtc8vb+GCsjOjPlW9S+p22
NMejaQjmPqOhdQAkQIni+VBRH5Yzpt4Y2C+YmdPjVK2NABn8+790zHsU2Bayoylf
s3ca2ZPclyse5CNEa9KGq902oCBsCp7ELoaXf+pLppEmbTeqdYNmOkWkf/0TeCw2
4cx9qpxZIrWRk5s6uDHdIX7VKNIOJdfD/QsXe46znQVyRpWa2rMsUHp9tTzJXqLh
8OxpszvPN4gWoXCNcY+FLDuh1y9lQWZTDK+unN2zgP9fZF3qXeyTzcRG9UfXYmUB
TUHyJ0HlgynEv7JSSJunA6SCncbEXZ+mCJFyPkpW2hD4AW1HZdylWC3PBonvEWZc
WJQiP6nOP4avhXuxsTSqT1gCwGUJwwLfdkROQh/8wmuH9mQGPG/L5BAGt2Fk97sT
1NlgxosfouHhLQ2XNy9tfbIAGYu7B5XGAlyKJSz8b4IZop64P3b/hVJOl7SJVGvH
NXISiRDJ9I/7IhsYVqmm8ujdQyn1z8uAdrkOjl5cIz9S4ly7nj6WPEDJDq80QJNu
zRiyJqc2Ryi7SCKjP1L/4LZLOyx2/eYC+R/OU4iKu+tGhIznLjWt7NgJzZRhpmgL
KUu8CuRtObjsz3jm9Jq+Y5ykBchJ56zdI0quiM93bcTV0h9441Mnt8cjhIX9QzyW
TeI0pcGV45PZ4XnXI0aHXH4f6fxgCMRdfxeKdYi9uzMkhWMCMChenVNuv+PbEBde
yPUDMI3x/v+oqN++wDgL/bIlkNQaLXDw2xxN7D4WjHbKCpewnyS48RlsdQQR4FDv
PQbXsUUyRx4kB6o96hgmdrBF6QCvRd310wYoN0C3Tiltohj3P9Ii/733o9JFDwUR
7G8o8at/cZa40xwXWQiRMWCdIG/uUQnJDI4X9uUJw1e1KSQ9JhSZp5XdW841OBKQ
zpb+krgULkVVFNeM1WFeKPuPKqeoBbn7TwSgYErBVOWaKEu7Y+IWUzYVU3uKG53Q
dZR3AzconrbLIFqyPsfzMtugXk/DujzoQc1kFybedMNpJ7OgBqWC+x1B/Ke4cQXG
pf+Ci9wKI9T6tK7pYa9s2WJYFhJfiiu4a54wpgO3b+qksV4tL9O+tfDf11psmxN9
0gdVZ31k7/GkS1pHIs60uSeQ4909RD+Da60ttH0Yei+qvXFII9vMGq1o7puH5ppC
oJaTc4KTlvyqvIoQTb4h7QnBCV2YrQT4inETK5CYYkl5bMY9jWH48fFZZBJublfR
zw+YBh2L6ZQg9JALl/LEwtNdbm/0Y4a+6zPtrunxYOPsxibsz/2J7gSRugPXZl6K
weEJ5jUzc7jo/CrfvjOwlyDsjs19xGpeUqsCXZjio5pIO4i8tMGEMtCG45b2MBDY
+LE34paT6jdoCcb+IB7pQhTWlEMQBEVd0oCOaZybCeqFELleXLdV61r8zADglMwi
A4uVZ0qnpyfJwfMkoYxfkg62VTsQLXubrjf7/rCjhVIMef0JjobroqMlvlK1Oj17
MoLR8Wv144O5x8OM8m8hbBHIGSKc8aIN6Zt0d2XhY81sWrsYc5pPc0UnPGi/56dx
ZoPMBuSp1clcAlIAlcF3nXn+RYZ9LddBBXSBjnxN+WfeW0+y21HCN6qD+GHAZhUk
gO2YhwL/XxzKXn/JmnIB5Ve1Bdp7XP9dAX0LnpcR281JHRxObQzQaCM/oNaO+eZp
LYRcvZSUpYiE1kK+PkKrB99LSGKSDlRqQ1Nk+358yG7hkckngAaphPkM6EI69cCz
4NRRVhBx+9BWE6lE6tT/xglnCR1fdptzgpaTxTQ9aSc3URdgTuuFoQvwFbJg8zNE
MuSGJzImYE+Zx3dSpSa537mpmUSe604ZwJwOUAWGAPFZIPUUYdWT3DTMIoGJ5kFs
8+QpePevQ+PCSnuGOi+zr5BkkNqMLE5bFwFYL3isiEdkHQViyzeAiy7ppXmRwn/b
DdYf+dIbQUwmIDyyiW1BmW7P/kYyP0YAkFrqLF/zHYtOf7LAbq0mnwtJMITrGEZW
yOrmE4t4NRVQsGBftsfeD9KlrQPPM06CE5f/MVU9qTpN41QuBKol0vejgzHmKMvx
g/wAzJB1Xz1zD8dz9lngt8v7JIoWU6k8jZV6j4r3JkExVl1kwmBRkpTrAMDx7Vya
6CQOVBtaSz/2I6gDhvzoR5brotr64u344W9C9drr17GiOlBiBhyZUkb+baZlVR9Z
hJ9lIBKl/vqWcOp1H7w7RWN8k3KlQSbhGzsg6BXQH09m164phqJ0GMZafdq1qDgS
JyJ0q8QEB/JHUOPKE1KiLM4S0s9F2UkTLSNKWSWi771IpYst8vjzxguEoZb0nGBm
Nam71eGt20z3Z2nf3gWkSGBcj/i027SCAqpnLaCyt3IXj5EWxJ1CkChvC+C7pmZO
RPh3C/Il+025RW76PYUdmfn3Xp7UUzslEOlcKw78hY/fHmqWcfZH06NHeQCj8kUL
I7bbLaz1u+LRBJmGNBl8Acb+zv8Rte4kc+OGQlTvVJ4XvHd0T7bOtf4cokeC4xrY
pH3C9sg/9arr3M87jFtJGjaZwRe/lj/H8iLNsNeP28ALgVEyEtkEtod4k6JFkadX
Xypv9Z61QczUI1YKp4qQr1izLgj1w251T+s8sZ9gM9qQM7zx+JFjLisSCWkG86X4
NvEXUHmOfPI8QgUYd+GcObve2QA+3j6jekTzZM8b6EZHFyMrCTlYlQiSKOiVGM6L
+3SNZ5P6BbVjbCU0M/EoPdCgq0FA1+VW5Lch9UtlX/8Ol8DcRv7fsd0IPK2JFMVA
vZSpt1A8T5PnWNjtUnwplfqysmFeVL279JI0HAA8ruT/K4v42Gvv3p8kgCn7w4bZ
hCohjp11/8/uHkIHAg0s5l6n8VPThOt7MM5zhTyT2bQNpx9AfrYd76QsE/OXRCf4
917KmGBxU5+mW3HOOr1/dU818ITrM7KFZMI9cFbRZIbxECQH0eDoSEU80whWc9g0
Ac8YnrSGOJvzt+oWf9cwI9qX9Bbw7dnIhr2h5+Q/mK6ib2ACre/zvnhVXskj/rDM
4wszikTG8iZM7wtAiBjvsVPOnOwXGMWV/cZO87U3BcvxPoI1i1nYYp18dk2nR7Sl
P8kvJkpCbf1UXj1jkkiut6ZME3dNia+KKS4uCI6iki8vc3tFuQSgYQhhokL7/fTH
UTFa1F3sMru+JtNbbNnayiKrTdZXYbMp+kB4wrNJNk4DuyVoWx5xQqUILxwJcMoG
AHtkuDRs7iV45q3WxogvNZhI3/jzFOj3aftFOYpSUNXsXNoNpOa93pocIKoyZWPT
MN1LMfRJJYNWZWL8qj1LKO0kcC5E8J9iKqsO70Gt35MvS7LmIQMzeWU2ZXueDsRA
Rb+JE5oBvPQqnXbrtWwb5IU3Ijwk6PaRYWEKbF0ykGFQ+NQdQGcYvoc+D5RplqsL
kLd8U/CbHSj8HOnRyJSlpZMe4Q8bWN8TocmhA8BeGU0Y6qzRr1/eBSO9aFfX14ST
vGJnoVevRLbiAeog8vUarZMtGj9oMepp7UwDuNYpVyUfbIX7fRWS1+H/izcIbKLk
0jOglI6z76SIGe7ev+iGHuM9IyzGPfhMtpsZBzcWB6HumOTUtavjTcdxHA2/ILxR
qdpCsQWXisuhO+26DgqBYJ674n5px3MIPmZJOjslm+03/5xszWv8I0ZEi1hL/B9e
iia4er9P85KK52wKPvAQWau66Dkg7bYCopZFyFIMgrUDiMSuA6JxegNuWLfVyg8Y
TtVvUSID2sEuKKPuSs15aPdyvGcn/05n4f7qxeTDyn1edpJWnkucvehIiCeb4vAI
RC3jb+xh2UOKrAdgmZXkO4OnbmIQ3NNR4xeg8sXn0Trc7KjLj0c3tENmsxRm4hwE
Lwg4pDImgrTT8g23snQbXBlkPVSsJJDWnedHWbB2RgiF+jbv0y+G3ssF7OrjPEqV
HyZPy9VZjY47dNjkSrrrquaxtFv2ApD97naPDVCROiQWQlc7uHuY0/5xH86IA/WD
WToIUd9TGza0wcv1R+yMpGwI2o6vDesfF97AR7YiCc86E7KKKwUI675LpjRvtB6+
K5tE34xmPHKDyFjW2AEgx6Qy9BWiTrrHUXB18minm/D5P2GefITJiffqVJ7cu3M9
S/DaeDxuBTdAokhR8Psqzf0PoFyw2BwIEmvaeHmzkVJPFYV1DEXnVUjQWWD4Rspd
Qx8Q4S5VIBpBRCging1MGllHThez7T6kGLiChTBP4UPQ2zg9OoRF53H9o8kETAGp
qFvXvdLtNhrQDyTRlS5K2vXHf6Hmgc9x5gVRK3w6GR4br/zR76OYT/JlaDobll5b
YpdmcygnPH2JDmyq2LFXEh6aK1YR31AfnLNFco68YYHgiaj5CHoW6Ns0uSHiUyJ0
glbt7vI810p97GcwoiO64dauSkan0yyYZDxJB34O+osq0/Nh0M3lg1VTcCxon8Es
zkyvG2rmX1BZ3g7O6NWSvp07a943R7ijqKxNoeZXPnKOg+45hnt6Z0eGp/ERpV6w
t+ra7LbDlxr6dvwAvSrxUGk8/hzOmomLWzrQp2DzeGMk7h/omZhP3ajx5OQ8BlAW
OVRYQGmYqIYDE0H3Ji2CU0r+r0/FT9xpnfUSgANGNHMAxLUdWBNA7yLIuLC1V1xJ
JeY/4IGDc7jOG8S3tYe8Vcp9+xZbW2UbS9eCy7vVAJoqerDiY0y3FXMnemDMiIm+
xRXOGcgifXZ9gnXlnlqK7CH0/to66pRLI62ArrOc2Kpur2M0+zOAvLM4Ocd0c4Mp
/x1PScpVXKcc1DqLrGfyWsjsCNx8k6yKv62Jo1gYvzhL6bfITSdPz0vgIzOVe1jE
+FMt/OsYVoEM7/gu/q4farfyJ9Ux1xbN1+Mt5VlQ56AEPJa9VOhHB1V25+zGzFnq
AY5PvtUDQgZIqbsYUwT3siI5B9ELtKrTSSKe9IUzAx4SkkQzexX0U2oY1LILWqNz
UVQp/kGyejFQG2fLO8UVBLNk7I51m5lxIcA23RnsCdWmAoNqJskv4E3nggL0hV6R
/Ldtkg8YR67xqngOq8i9ohtDSaKcH5y68saH6K3Y16wZu3VZxPrv5qZjMbPMApLt
/B6A1X2l5Btqs0GmHIz0IgW1y1dAPPVuM/KAiVMq/E++BDhnViSYBcy1pSS3XqEw
IxUpmvwaBXHkiBz88aJnAd6ImOaDv+0sdPeGsC2lhBEhGFgkNZ3r7YbQVVOvh5do
QsRabRMPIjhMjD80HE3vTtR2Yp3G+kLqVzx+PDj+zQWqXTpE/PqfJi4K6+hPdF7W
eVI7odj3Tu4+We/7JDVeQg2/9Jr4e2xGN8mHYR48MzYZgfvFcWgFhHuI//mRcO31
e6SxNsyjB58CFqknNC04s9Sax+2X6YYciSg4F8BMBGXHt/eY/RudH9GYZdJArtAs
sl/8QfIMQT8Evv9oEzhkHtWgcUdazGFQZVCkMG29ZXJwiTjJYzkJs4zqacp7olCM
R4jZj1ax+QxrITl/G2jUrfmnXD2onf7eAjZemM4IIycxVRVNXpcezq9xi1o7eR5i
pmhguLfIkTpmihn9rnshTRWKY9H0g4qI8OD6U++drRC+QQuMoRKZCTh8hz8eZ8/W
xtlTSr+DAYBNcpwo0dwYG+TZN39w+ZBeE+ZUtXioz0yZFbiK721RawDA+CFJMNtp
6TeEfLsv+ZpML9xYvzPmHoEIQhYgiAkAZaSWBdUyDYBccJsewQS5S//tR5F7gfkU
M7Wqo5WRwLSmtsQIdOvLwbh9oOq80ws5pzLkatzWWhjxys6C25QxId6BAuw8slBB
pEdRTXq6AwjpSQ9J/uqU8rZQ/q1FmIjHh4asEcTB3nsZGcv2jlyoaJF8LnPdsSbu
pwcsL+LUT+7A8B2e9rn31m79QOsDK8c9TC2etVLFZ6Fguh47V4yyWPvvoe3Wopxk
4S+76sVUTbwg3aZBtJTDK3uoWRRLOLRLXU5zDZNyCQbWxFKF205BinV2qxskhBnL
V+xu0jQj+HNzRSikPD7Rah87zjd2WOq+UWLC3ZkkfZMCzn5oFqIqfJuI6fwOmic4
p5q4POLjVCgwwY03x5jjBMIKm2gHS+VjQU/hggqKzD7MNcJj+dUYRRMwqIrfC5Ln
IhqggBs6XMpVdTIMG9XpFED2zf7d+VKBVuAXelzXOERCJfV+D3gfDm5yJ4JSdduI
jbF35lNz4helVJW8ElYrgefPC3itdCnWx+gfjumrMmZ4EBTW4MUzN4wkhfbRPyhy
8E/PBB6nFUXpdFWWOuUiijtPY8/wvU1Zh3AnzwCW97U5WEgz0dAQaXuHWzGiqXaD
WUGLRmZw7EvNro66uwbXqBhlBaj4QKWu25jCj+unbzT3y6uLHxnL6OrdxzXWTFAA
BulL5V81W4lI5mjJEPZRq4EK3vhxKP+ez2BccpOV4uGCFPkT3K5alc7IKXJKIl12
ai4RHhCymMZhy/T3s5uWWWLiWy9/tGS1rPNh5ItbECy/KatZVRmL0RUvaBgw12m+
Ir9hvMH1dmICdXdO8dJ6vkA6vzV2rRmiiEnwnYMsxuweaQZhMgSNYZp6EbR129AH
mbOOPSwjmPUwTrFJF+CKQpToYzQBrVCYKfP3/gHCW1cUWTuFD8fEgt+BAX1XL2UH
6DPrYZdlPOrzztMQfkhJWywHchMvmnPyNyiy9V2nRW5ml4CP3jIE1uAj9iwkF3Nj
sc3Yz1TaPjmqopQ1sfYpAjszFPrdbArDaS+dgUNsyt+a7LWvNimUfTM4nj9RHZIo
AY//wr6A1vHgrQzgOHVCpocUXjR3Vdoubcaeks5cEqOzODY4XId9fV1pmZNst1Ku
Y9shLXUNKEMuacY0PIwAhO+jZhZeiGDCksecwvqEFRVs11cM+DV2IX3J+zQ8V01b
jY82T3wSsavHiGpPcYmH94fW/abfX2/SnrR6gdbUIvegCrLgkAzSt9hujBla5CEM
/GJuCYoABg3gf7oehK6hzgH+Q9qHuignU0C/Om9mmystfZhUxEsjX0HV4p/MkZlr
gjnyNwWHFWkH1NRe4vsLGVHjkzuY13xMouJgeHuqbBNoC1gplqVsJDRoK+mby73A
mxPpCpiFFPX6vPh1yNtFUJISZ9OVp+bsdV3YxGDSjvbfAwG7lwxeims53stjA08j
tkL6MVQCGI0ATKGdIymcueoJWtDMiI9CnJyxtOLXTRCvR+BrMrH7e6SVkx64lS48
UyJh8fu1Vaazb/e0Is8qO1u7GQ0VjIwTjsnZiiwmHMH/wia+IllUl5Jf88FKwsQj
p78tu/0BWlaDSONSKG3YjNCGX9dqv2NGU8OWe/fN2i0EK5MZwBqm2vNW5Q0sdAqg
WCbfUfpw3hhy31YoC4gWDhZPT8T1hYlEpabAmxhFg8bbL/e6uYi2x4D5yjJu8IL9
WcGP/mDnO0LHeXkQGFsP+e49jFCogxyFYmsA/TcYaUzYkIwr4L+4wCvFAqD09EgT
Nr8XJYnDWwdEq0C/NIiYP+Bojzmvfvo8hDpnOnR0jb1Bwx/adbbB3HEZeWkYGZWU
r5FEjfXXnkB0Fc97tpg4FrVJO978OW+9lEnpYGO+Jalt6w7fPDpjKjIwSOc7N/tB
/DJwseIZLS6d6aXRoMTuZ101NlTS+FUxsXwlGW+07Sl6rPTCHZZsJgQPGb/YZLK5
+g4R7F2BnJiXGyWfuMXesqUq2HHTO+KmlROn9GFw5Uy9/n5BrcyHy2Gymh1BczPG
3l3zTqk3qr6K59x1EPDoQD0I4nsE5AJg0uiEUKv3QJaMSo1CJ9c+GP2t/7N5iZ7G
kXY1+wCcKq71qjQhiF+q0+he/ToySgDu9KL4CAy4zk7/Niw4+IGxf0yWkSpwC2cA
0OJfJlCpcKBV0Z9RK/PSSj+2fZhdUcK8bSisRc10f4GeL4slq+poE/im+PhRwFlG
T7GsA26lVRlqoDK2XJDZQrYXobETdudNxYtKDseIVs+GQAogL32E+INlt6jO4LNx
7fNh7N2Az9N/cXQ3Xt947+VGPxPq0FOS3gciMDlY11qAeay0chSQoucwA4DXEdRP
jkA2kZc7kT5xReRoSbqUXeGoLrpsmNaPUs7upmw0treUr0JEerVVLNwQQBIjlNe2
Osi2rGzPqKL9JAv+igaJIzmNHVx8jYcbhvn2Pf+gvtGmz5p9KlOVlbCmjmhVS7c+
rS6JiJNB74VR7syUS8fEfN+B3dPWKmJV3BztyKi9GfI05AveFDMKicbK+uClDALV
aWNPpRf5fg6GGciLXtMMX+yuXb/prjlxnqT2AsGY390T6IUJkMjQU7bIAw8n5l45
bxirGfUXeVT8asPfwHeuR//1YHt9BuD4bKSdg4qL4RDxq7++wWC9pS4yqxribKX7
x+9NpArhhCWyOdo+y9FUbrYaKv/X1Ef3zS8SnVAKQ2NDu1PqOyuA/RRG7TdGgSrH
cgRcJGHRUVHRV3LcXWl+pSB3BGKctSqrfS2eCF/JTdSeqc7Voscu669Bzbs9/Pjl
im/pmPlk2nDbY7Csc7rZE5BeWDpjVORw6e3AWQ+TlpEWE59vul8xyc/79ARbeTcF
2Htyouz1Ee0R922svCwwRgWoU5V+h39ZtDkBhIepzOFB0tOvEe+sm0VzDCuBq/8m
7WL+AlPv42WG6le969X5lJjbPT7MOd4qnv0NINL0uYNie6Enq67KxH/TEudqMGsP
smniqIZiAuGtK8obF6cqjMzXxWYWpa8ucAB6LrHsHv9HpDb5KR9qQTpB6ZROdlh+
mWEqwP6ehnKQs19B2f8RWFN2zeObiuWD29q3jlz97g+8njDf9iE+68AyZ7zgPB1C
iSrl+/t89bQyIO3TruyAnYanLyHqiEZmpC8Svh/CXC9EmINcrfi6u2SgWjDTULDe
bPCnETh4f3iGWTLDtYuxW4TKWQe+iuEPDJTcBlUhxrEd52lzLW0Go6iq+8XVxPVU
H+z964BGKPb8NKbFSsn7LEs70nXpaaNxy1CubZnj2o+FkG/tUM9lWP4hrnshUKpc
r1/SadEElXfHtlPb2Xtat2AhEiVLbWkcuT26+Ag+D/ezzQhU/UExQKWvDZ2DQWEB
H0Oz0eH2UE0e2dQ2Spve+VWKc21wDH4QWcS3jwvjQHj4D6InoQtfbX6OTSNnOEOY
PfMpGiTaOIg9ms1+btSeo+TWLo7XOyz6ECz1iCUGX4BfUYXxT5ebr6e9jl1YEyYV
2LPYBmtv5VW3gEvkXF/umlS7owTDS2PIlWcRkUtxYXX5HN/RyPpLg5/Oe5gPbi2f
rXUt92ok31mqGIQS5X1MqAhVhC4IBaHPHk8R6iKgvNbbLoMYo/ugVNBV3D2LEibT
SVzAATX5OgcZ/6cxhMbCntJZLZ3bp+iEgf8n2gPhHevpIzkETR6qGqsc8vIf/I5C
kAZSL5qrmo7Iz5y2EiWuxeptcoNpbFjrWvwQhLHr/32cXX4OHJATNjhgknawP4+I
eET0QxngKKZkU+41Bw9NTSWLj+XJDBuTw7xv60Unf0mPlzTjxQetWGDi/E1JhZX1
3yY+taUTuvnlDXtT/Ne65eEXfWyzjPAPBVJoYAbZUiHrwNHGg8n+lPpZdkTYnhG1
4nVgBZ8ulxBYhIsBSWF6zstJNhOc7DQoXDSbMfmuNDD/QkOw3q/zyEsDjtpINFz3
mCa/sJ4HNe+ugEvr9kN4l4cMtfxnuNzCEZre0lDIznkDwym8MatfXMeb8jiE8sEL
WcGT6sQGlOZhsqokuKjtSOPeKFPK98njlB0HivY0/WQVDvl4Ip83GOtciVmL4Pv1
AT8UjnhPccQkLsmUEQe+aFbWI/gVrUgqbihbqioCbW6icK7/7E0FhlQuSUKYrRRa
tUR6zUvE6m6lx9XQM6kljmaVvoQsIaIbgUOvIhSQOF8nra6IUhjHcVb8Bg3nSvaN
e1AscAxHQoIw5KJkDca52FyRowYger8JFEFLOxESxRmUu7HzoUw5PMjoLXNjOsOB
/RfWYG8CLurgVlY4f5JBXlu0bbbMY/86geMokbbmY4cv4RTRuK1dTBtcUGNmYZTT
gusEzh+cO+iTtgN3+kOzBKCku6oyrKPofMq7uETvppGzP7MgQziC8QX7SqUQPisu
VWIIVLvVWGsSJ7B3Cx5Ffn3K1/aLT0Z+cM144xofXGFHhepeLppcJ1tfsX6FWlGk
IqyAb3I28N/SZui69BobMITrv8r7Z8/SD5lcEfadF8DmAiBAnLuqgrV93L3eU2lA
4z7NbP/QBAvcSjDab77P88io/C2zOuDgmIzPZUWk/qzr5JfWpIFhoXRoGfnQTIY3
mmpfGyffUlVI+rU7uCP57nZfgULfQAaWl+kM9qURhCvOkOtqIm9usHkelcEJbG9U
hizTuV87e9xAoIXcfeS6cPlkrCHJo8V3braeAUzTpQbjmSMWhiPWrDWR0o6TKyTX
Bf/Zhykx/ACk5K36F2OPi2ntb/ZSa3GOBjSrz8tTQ0Jjr55TnYfzbnK5bb4qezps
Nvo4QJDM2GTWIajVUYK7bycrKI6AHXJcmEPiyBkwUNUbMrkOBIgAg2ZAFCJ3yZrT
f3DBQKuz4/42EtoyZTkw05/UtkIT7hgYnYQMbjXFLfpgxHdd1smwx9jP679zDgnJ
IHw2HnGSVQrPcG2GJnenFQ0+DcNy/4dMao3m/tb9lEXy+tZOtfU73R1unmCMlnzO
ZceJ3xY5o3kZWfWPXBjYePK4f2hMxxFyJwm+6EJWMdKLJIAHv8f7iNddjB2YFuxV
XufctYo7B5bcxo1d8QyMayKLizqeDj+Puoma99dDuR7wKUB/U68XUE4+JCXRiMRG
xXGI6TykSGQGZF3MNadadtuosnmhSl0a/PY6+2JxHsV97g//I7cufaRToZcEWOmy
7GNw5aOPde4t6PbWnsfGiHRVvU6EQTXH8lZvjCyIgaCWEBSR74UysssY7Ov0QDJl
fSoJ0mnomB3+bE0ukgcRWapvP8dJ4k93nfPzPkY3tf0VjiTaC8MazOcQ06e2wRoa
nPXJyBhkRkbASImPsQ303FIOsm4CVKE6hmaO76YEhvCJscXfuIc4GYFn9iLlh4PZ
1W5Y6GGuKpOvWiYR3dr9usjmsi/htN+kTfReH/n5wHmHxPdECLCqsnMcrhoflOXE
9N/vo/Yr4NdDiMdvL96c/PH6sh/6kmqfMEnn6P1yw0qTqnlskjSmRyNXFpeduHiD
UJATWCCYj6vlKnuLqubB8IBGcWzmiwpuR4RGpqf3NADiErtwio7679XLakFKzoiZ
vcxNPsI6Ctt51OSGxz3i54PbIHk222HaSyXK6ObRmFIh5IN0Q+lVJhacqmBHJ9hS
wzo4JvsefQUTI1qoS2Ihj4j0j5jmdq4vQMjEi7NQ69uZntQPF6H2v84aFU68Ts1c
v0JGQQ8HfExuUtq3bBNIGZGNspJOoxgNk2A7RLk4rYTQPfFWBVMr+m82M8+85Q0+
YPP1G0aKyGd4GX7/WQuiQY02qavZO631GEJGUnAu0bw9GVJSfnSXrDlkkfRYxMa1
dORyXGqPmC0N73AT1rqrTLdqFAxiNL6oFVrl0Zm3CGSsJ9XmXP0drhoXES8lxnXb
1UAMglvaFWBSIsEeSWoT4blX2sumStwUhJPVCRsKbBWhSbtOXV3VBrcyKL0MEigM
3C/+R7Ojv/Jw0P/8QFl+tufKEbKyG1sF4nVjWstJ3uhhCQ/HuFA8RIjoQVD0ac1a
+YI8sAACT4WlB4VrrLFLklidPz22f9smvFnNu8ZWR67g55Pd2bvMPdwG7ZRJBk5D
L9QjqSi1sQ06zle2F4w7kXgtvpjR+BIgr6g85aWQOdioH4QbDMOmtNBF2Ak1Q/WG
J6CPmeJwTUMHxmEBinZlZuJllGv7Fjb1iWyfeleMSfzWvaK1iOp6+3bbkJJkQ+hT
XUUEwCxONDQTCjgjhm+nuZZIsoKiheKbl9UOUibajJyCq4lEsd7WwJS5k1T4w0HE
ECfGV3i3DaMjjKPXH/1NzTcNVwvRGmozJjyVvurpFZ+cpbePwEkYk4C9T4kQASGj
dz9kQ5wxeaz7jseiWK2MIl7hEKQaeSgv7NWE7vpm90C9TJIVyQ4KcnBFRQ3PBeDu
lqHRhrD/Jm0ti029ZvYzEpaG8B467WHALRs1sDUO768gTiAsNQT7wETOAuBz/qXR
TqHCK5AB8Gcyb/G/35MquQxPpPc3K9Ycwvqh2sMCQAYMmnEWu8v5bdBGCxSF0MXc
IlHtD/2m7At9cgCAHrxXf4q1KHkXWQzNcfjDJwxIorxqUfRQUc0pD8SESMAJY2ZY
fIRUuvy5VRksuwJqZUgPVDBtUA2OzJS91TB+IUL1vwu4pN5lzvtM4Mi5k0QVIk2M
/Np82gQEeZq+RegXu0B4yeq/pok5cW7t7OAWQOeqjZC2hiq8JNZLgOa9/5PvbzVd
XH4S7xQNrhgcDABTUaHdo8N9R3TCXB1CGJ+fnchKB6thVxvcuqjwXiPP3JgV51/K
i3+1RPFMZyxggC9qmmH32Gh/vrqLePSFytPjBKgHbAsf6LzEEM8fIvXu0Kzeh9Zk
F4FqutvHvjeEYVZsYHhN9j+RHAI112JWqGP8J7IHJL0+V/Q97q3GLr3M0vg1kT93
FDW41ez19Khj2+jv4p+1OMXwjNOi1eTDjm2c2OXXB9PCfVoZJcp75GNL5JIzU5Au
lIBJyO+u5Lyz5J+y/kH7/w7UFutb9dDhxcvkHr7+FqaZqldIAGsWVg9j+x4snatB
fRYwfiIaf4Ib4Zsk5TOGpFE2gS9p2FBhO0Aru40a4ptx4jXs6q5HPQy+Nkk7AGKN
Z+e2ILRhwI/heahZ8eRNZgg9tuEtjdxa+vy2z5/y3EorPD3wpIi6FlJFT/kqGD5P
/RkYt1H+lHDkFHxYL/LEgHjHaWOd2MfxYU9VXndcIZv8i9grPEHDiCh/FfN3XerR
Hxo7CQGXP513M911Y0Ctsx3XZ+Un5/tn4vqrt/ER6vQD5iGMZQFPRcLJCTaZNFdC
lkDass1PoaFzZRshFaO39sBqxG6yUQvjYDmwILgHOWZIazadh+wS+lxMrsa0OwJA
lkD5orVdvvTdif2KilXgJz25bYoGwyDNpcjkg8DESC4ANvdBDsZEwJk5WCqg+eE4
ApdKV0ApOrJTHw4b82GEdSRXqklVA30qm947b5rurxDvr8x70HbxuU9q0ZHdJKTf
hQStg04+xvjsH5G3GAXEOkt9SzCp6qOsTeJvlTeFCzYZ7XzgyDa1VXYeMdbP1Xuo
vRl8/MxdrYovQ8jpjnUurK6MlHARO/+z3ZPaFd8RyF0/hd6emZzBop50RNKqdEUK
QnlPY4QVVt38aY1nj63D7X8yEojQqYwR4dfG1KFVelIqGdYpu5Qd3dhuQKFllnOL
OicbWyHcIJGF0HLLxBAfz0X4Pu8UhYcBfHi6m6AdMp6GrS694ZHEgXMA5ECYMz04
/HFfz7MsJnR/FGebLTaH73m9rFhR2FxptiqbRg7IQZYS8Nb+yXwVv3659eke1B6K
g4rhIXYw2B/vGG0k32usB8ahCuIUN9cv+PMHWStFUi6VayQ6wPzhEUmTA+6UB4eh
UV+dveKWagR0ueDdZmtYBVlOt1hgE8mXOHhJ7qwHq/t6tD7EUo/Jt2nPkhkHhyD1
jXjfjiJ+zT7udOoaSnqsK2Jz+xre6KBo8Rx4Yn++vH4nT2FQMHk3mUorH84fty5c
t5bLPGL0WxCwafdEojLxf8kc76//J2LQw2P+LBTX+9+Zs7Si/nVkwSaa4HaL5E90
vaBSR1rI61IUnUeg1hS6rUtHbCKQQu1iRcGpNEHhzBC+WYYrtJez3qlEmlknjU4w
8KAueovECyuUpgTD1kfvjw2VvuhbSQQy/rd2Hen4fYuf0zMr4myKG0+ro3HPHba/
axSSLUGyLd8Qy1WReFyfXcM3AMhNh40Y/P8sXzUXw4jLZWsudtPObxHzRkb2136+
QKHGz/SF2GgUNvcDcoYsdhidiDPcLPg3ALeiAnsMw8rRValuYK54xjCc19eL3be3
BRPHQoRqJ5cAyov+6RjnMeAOZAvi0F0oXOfg7tJFUBGoONvyIlvbaVYfWmY41nxN
YzK53MuXyuxVU1YBnua2yXf6IFBYwaNOm5+MgvQC+wO4xTqymCSrt7dcVR655jAb
n3/0+aKKxIhlwKQPF6nRXBK8tuHK97Am+GkAzyxfFklTDBgCbYz51bAO+N8o2X75
wOkpinAgN8ZN/KTLD5b9x7tKx0H0kAbvSiNGwA/UkiajbKkTEh+8+I3tRtN6hC2h
L/tBYcIzBxM0de5G+90biwtC7DppaVUunQS+qdn8JhvUqgO6vHWMatHrMTj6fblg
edY5rc4gb/xLAgCw4rcy400EnZZGtPflqM0SKZQpZDPz9lNIJkUQsFUFw7pBkkrJ
2hqGHYv+9ntromaKyD42YIaucA1NKyg7Myz5tAaHNXd6TuMjEBATbrDryNdL1bF+
p36NrWKKRQdPyyZqKvpHGp3qk0b0BR5XGFuxRqJuTZExKSDx4RNCzm3wUGUUfI85
Ahky1IsbvPx9b82WKfpoQczPG7Lkk4zgdgVXTSwf0HH3MQRS4PLtinRuCl1i8R+0
F9JjFBuQId86omAk1HfgZZvLclfsVNW4WBRJ6KfqBG0Fgt1B0ryLgHB6Bz4PLT/6
fC4VutK2VuN3OVZpEmRRpQs/oN/0B696agJ9GzfS/9kpDiAtC9h161OgKrVedrcB
hDFVCS3Q42J6m3MA8v8jbBO7vG9ToXH6F69rtWdB0gxdRQSIuj6/1P8t/MUGavu8
eoBB/cndtBd6skQIoBUkZy/iXQ7tN/dRmzhJKSzcZGvuGNUeOdBE5mudY4BjZq02
+nawjCCvJ6M+7ire8no3OX21GApBH2QRmEYvdEi3VFx7cGnuMP6tgX6I7/+2a8o7
uPg9KrHPnApoc2NSXDXtGiP05T4ZcWcNa8q65Q+/Uk+EjeXoVRGMOp7O6CYslrVh
msWmDGGxGtuLTP0TfJosnBzVO0mzu9ObM1awFZ7hw5vM5UsQ0FcVU/sQTJs6RdfA
EMO66Yvb6rqh3EHdJplzHdk0XA8c5uDAh/m7WelJ3Ssq/KIqSyJ91aTFr6zQaeLR
vMwL59taQxaTpTe6IBUV3flNqh6yBix+B5SZgp94cJcZI7VdELYPYlzod0Sgi4ym
/mpbSKQFlbXfxMWFeJkeb6iAycTihSailJjal9Mf0vK8hgKDUOlnClhd0U2HcmTX
EBJJtXj82VSDaDXMKxV/X2CaJTH4jlGCaVKaX2HU1vAzRAAQSjX/sezQB9kFs0lY
B8ktQ9OVrvSiOBR663CmeVwLubiXIOpeabmgeOXQoeHIzrnZvZ/XhYo6veSO2ZrH
3a1fx2TohYoQGgTkGJBnmN3atj28GC6DtBNgZbLZbTCpMEXhGI6s9OyeiqKLYGN4
uBzsdKLkJMc7d0HhGO08MjqzKqsOIRjRFRO06FhFH4kacKbhmlHqNaWX1MrKKwA9
gy6GVRE4QthDv0AVq9l6rYPiQsrV6h74IvSQ2kcc7EigorjMmeayhK4M8p7DW/c5
R26f23dIQgV2/B4EzrmKXjsdQ26iWfs3fUqsHi5+xj8GO/A75lg09sqosRIm+cJr
L6R5M9LXv7W9SnmTn7aD7FwmvHXG/OZ19n6kzkpuLVnZ8O1U5LY8HznE9M/FBP7q
cMQ/V14HVveu8xg3EVJ4MEGDr9BZsg3zAeszPu2nCSokOQdbIFkCq4/ZfxdxXHpH
7FjW+ofJyIXJJKA3fvHgjbvXhS3qWY3qk3UF07zPMNnH21D1gD7CuGQj1zB6T7Lj
Ra2l3M7szNvsD/F0Ed8BXcmb/k5jeg6qWsVN4BEKDW5FEbzjk64/wRTqVwtBMdgI
1qc0qJrCUtZpfQ7AkB+KaAwnePuR1ZwPgpbz7j+XqfmCybUdFtUHUo0SF+1tee4/
kC8d+3sighspSoYRDi+sgFET4ULmW0DPvO5b0TRsukdx79hL+PjVeZZC7GuCL7vb
izSWm77Ecj+U9Jnyr9rQhK+6TLb5CnEGdr1eQOaqsQGg6y4dutRa4nuxoTfQwXWd
BPZJZUp+1qQ3MGQ3Dgcgl7N1tGTiCs4UtUJH8fobRtIQ3azax7lNh6DVghYPXR6u
PtmVNAfj6o00wQRJ8IWCnZenXvQfEOxKE7edFMPXP+pVCT/vANE33Kzge/PY4xfc
TGCzbvkvcdF4dsNKT9S8bJOrHsZHf0iaI/lhKBQvCfim4kM3GcYRTfRRgl8xVJSA
EYjq26YxbzHMorjZwwNRh0ZnzjRUG3KUJkiuzd95jDF+YN12uca0fdPQHG/NTifa
uPcRMTJhLLEcmdUWV4w7Ej8k6u/EPMDyDJzFrlTHhC18QQ+ns9BaDXK64bQe82Lz
xvPFEEAMIvIJA1tT0x4vKd6GKk/oh8QzXFWF/IQwZMeaXcGm2WeoMcrEY3w7BpYm
EexgcVsODKI8OdOzQPlalIylxJyb1i90BzWaVcA9sIgEL7IXQpQGPSRFJ/3aQJ9t
BjYMOkw4zUKmIJhMrRZ3nOsAwN9mUzPTizf7qLZQWPlej2Wn4gbbDH+exH/UObc1
V8YQFxYzhf8x+aoawCbJes9r3Ys+4ng/menMsqC7aIz2bEPVvp6xE4SnPL7v6kDU
rpZQmu2g8zlW0aGysjxSHgydjIrVwBwqQMlbQXbB44ys8iY6jhsKoTR/GpZLrSkf
wntFqtBpYCaVTuBK7PI/SMDFX2ydEMPImBhNYDDvCV2yj3dI4g1vn3yQPPWVuzY8
IKGReEjsn6bplAdw6w6Ri0CMMHF11VEuMNegczGmxV9d/DyBGtyWhJPW0omDvQ6Z
mlPiXKw/YNhz2gz1tzpJLnkGFpTaUlMDhtsDncsN0KJOAYB4hOY12J/9q9QUgu+h
v8Am+mtBPYIpKzO4zWNPW3KAc58/M/+9DZa+rYG68VuPs79tsF7ResBnRpGKkOFQ
9ki0JAfZShGLc6rsQO1nEZFNP75HMNTmfMunaUv7CiG2XjDkuNp/ZbGF4oUZwbd+
IU7g01r7aYtcO9SrswkUScBveqm51rOrgP6Mk8VliMniHEWn07rDFcqUV1aFtCLW
AL/G15knJNNgsvmWX/RexLF1nKupxEe877SBjQQMQ5kS8UAMYDbrMUd0ctCmqH9L
jDU+ZYgZ7xTAR4OlO1e8qQRDAs5CgXfzp3PlIq649fBDBBV3OndVoPUkjoOWoqlS
QweuckmB/sP0eZCMBxbOCN6+xr+hekJRt73N6dNI3yAQjXmMjcEu6OYBY29AeYlg
Y9FMwIsqGYLLNf89EZqpqiZZXvgUaXenvsviyPZ+l+PBduH8Rz190GEVKyv5AEkP
qySksAmOLwIT/5bkXuGMjaaP2zXNTSgJfizQ3AkQk5118+6Cftx/TqNWfMEVW3Z/
edsrrmzuuwpY+7AbNjMg3pEL2jLxvJ6Vb7ySD3k0T8z/rqGahUC/+9aNzAXgSWa6
SHifzjcHPewO5oDfWas7t27wPUUj9ZepYoQTcAjB+/RpFVIbePGDY0vTHzck5k3P
jEsfAcL4DEulloUViXTZEYioU/4uE5CetXXybVHjHU61iY90JRWWxqHnNmKy/8FJ
d9tYksvJ/Um2WgZ90evp/qZW06deI0gjG/ikzaCquOc3WanyrI5Q8mXxPOq8p4jH
idNuQ5hRgj9ye5L2nMSaKS3ZBXUkwmEor3uGOfVw57yQjwco4j5NnnIsncko2tja
9HpO+YgVthWladrck0cdBjhnAr2VLTfQHqTwMLW54PZ2rMHsywisQaVBjQqUR0VV
fZZzSthFiofH0tnoj08WfxXhA5Pc5B1pht/o4puIdZHPiqRmPMGqWt9CemMbHAZd
eByOmFI3FFJ+TnFG6gj1iTiTQtGZEHVqlAqISvyjbYTdC149Bqujb/hnkoO6XG32
tKDOI7pzPGIQavUjHuEiHIV42V/ps0OZy5A8Z3+zK8CxPsB5cJxercfmFV2IyLuy
T0r/qzKgjbztFs6dPHT66/U24kNvue7m2dAJpxTO60eCa1OYS+vd+pKzV/xgbK62
x1S+hE2EhvbIstYEPGyNFJQ+IBISw9jQnzwZlqEFi7YUZZCNP442CYFjisAlj0mf
MamPt8RlGfFqrQREFonBMyeFsVTV2953wEqcemTOgZ3Vnh6i5JibVYtArYWoYQIb
qauVwKRjhkO6cMHpg6wJ1m9kXFa/D30JZXppRv/c3oBdbvUQ2el1qDQwljpjqd6B
kXCztDH7DcyzFPr6qz9dB89U/WB3xYqAOV0AxwyGufodjirQrrbexALf9LcnZHnB
rAky37klAMHREzGZQ4vacA4x0Rfz2Yuvq075nBP78ACMYZ5NnwZ2RuoXrhk4WWHh
o4bMQsRv5N7k/05wZbpOIjY8tte/LFiHlAENiejxbx252eZq2AnFCze+VNHQezo7
A1+CYidgJOXIRsfWtWw9NGrqNu7rkP0i5vf5uud03t8uzOeBBr3MtY+Y6uWLh0rI
v0cG/rBCq3Rtywp/v/53kngq6SaNvQXe7xXQBRnb8ISneasbrOzVnUvG+tsl7dLm
7jj7kA0+t4ed7a4IiaJpqXsOBH4QJAhvGhrmp2ZkQnre2hwEsqnMSb14SgYyVMwE
3yucQf07Dzkv+eQSrt4s7x0x1DpBRuo7U2ViMYwAqt5dsXi2EUwl8UWp4s8wKqFE
wNbMMmCNNTvIkbg7iYaPzVw9NmskvkvcSpex9yXv886NT1UGii+TNXRABDLt/C8n
SX+tXUlOB4BGoZtldb5dJyCt9GDZVxCw52TkPnZ+1c4aaxHzsXLfB730Rcisa/qp
LfF/uD+Hvk9ab7dqL2XrBxGwXcePEFWKea1PVJaNlBZ0SMf/QMGUrDmqJebNcX+X
zzgWd50J1LXqsU+oBebGmyK7NLdcF0Ar1uzO8LBmRElmd7bVaKP0dNOh7QehnqXn
mMow2ERbzTeIoDv9zDUyGOsy4Si9WUIqhwqre/yquOcWs+xmBUlQUBT8XI9kGUlM
u7hKld+rLaVix6HNvTuHc19R13ZkZhhG0Lsfo/y/r8EJG3gzF4FvpYKlPNLE+oZF
/KZuyWuF6HpxTPZeX5cIL2uqU9fYg4aqr6I5Gaf3+8XK+KfFg7MWKLlRtm9ym1tg
L96G65rzgoUxRFIIryylwk1sHjmhx2XkXnpQ7BjRQOPjhl3DowEjXDMqz/tTDzE8
QYv26JKt74fr5y5Xq6P/obJfyuqYjzoGqmF0P2JxhoPUSZytFCahNco9svKuq3C8
0PGpmEixt9rVdsBEpKQ36pBC/ile95ayZReAPxYPIEf3uINbahU3p831iYfngT1j
BhZP4oFhlTNdz56p4oJNfIcl7AyQdD1REqTxSegxJksXNtB8S+NtM1sB+g28mTWn
kEKjLWO8luNFk3nYWF3XiNQ8becgE69noXwmbSLB5Il1HlNtcyYmGOkwZlIC5oNM
WCqWHI+bwLJCz8CuRdftx5PdhttkkkTbMHH9c+tU4gAh1MqO6WHy/ix7Y66FdKuR
i/JkMJ03CcgpKoT3QO4yWBNSKBBeGPWGH3t+OvDYBdo5VeRf0J7HlaGta6mBvUaw
L4Lkn6Q2Oj9vJb0wKQhz5E9dti5ku4kzj1k/rq1mXA3C4P2px0SPhUUQUfTNGi5+
SuwqdZ4Pt1w1SSODr2FadWfz9OlSroVCzOFJ6QEX7z/ojrXpqWfcAhnnWAi4A2H+
T5J2/P5O0a7dahzOs6BHP7PkhYJpbhwCuoUeAm8lyoac5M9yXOHj9oPkFkEvWFE3
++R5cVYq1skODgkoVi1Qs+6Cj6Zm9ssnOrpuIkjQos6YjyRiSj9QI8/m3lmwgrtV
B/8SFiAEBzCsccy3hEg2qGjpmeDb8dtb8KYeXbxCbEI/WboiId1R9M2Yi5E7hqQz
6kpu4QBvaNVI+dwkcuhIiCU3ojQMIUWoqyL/tJCkomkQ2itQCC4TCBBaEiyvNqKa
Ktx9lWEJptLGhU/rGj/JCO52zPn5luxNgVLQbMChmkZ2vDZGDis8lj+TCML1Umgx
jVqjqe+ckBps2LdJgax1LaHSPWZuFi2B8uBh7Hqd5K/wo/6g5nR7jfRUZZrwanBh
oasF0vhE3rqQgNP+7pUxangVrT2zt0DWKh2CkITZRh/esUAJdE7UWGeJA23u3Gtw
hrvvFpeDbZ/1J8/TCJS1SUuSGFURWchtwxFAxlVOH6fJ7lbqOfGNb/oKvgzvst/l
xlx0HHLR/sItFb2mxm0HCbH5m1Zx1Wi5t9Xo7kE7yPGGqCsjJgdiRaDrjwRj0qyG
uzU4QlGGRbE4uhMchyTlXxBt4bBE6H6sVUBmgU0K7XlFx8T0ieszpd3hvirkdqE/
XUm5dvddSnRkgfEVQgTH/ofGs4j3/bGTLw6u9Htq2xSoLNpcA3Hp2MzsMmzMH8rO
jS7TI/sNdVD1VvcRxsv77edRu6MbHVQsqyK8bwygNrZia6fWv6v1Co0HPPOQrJiq
wIwDPut7NSjYYYTvV/WaX8ifXKcBlZPkveOodr6bNweaLmZYNwYU9s+pihKNKpZa
C2fi11v0snJPCjYEFPKkXcMZ/snZuJpsN/ua5uPjz6MxKu5QUsXNZrd1cGic+Z3i
qJmjfkWPi2Q/uJBGED+En1CE8RjBJfcTsKZuYXRADtVRYNRoWrLF+gfHQtk6RcMH
XyKw5Sd3hIJJq5RH5/SSNfyl/uoxQy4EMzhHq9n9D5tbeDyD64FpbXatTa2iM9FP
PAkwEA3nnRG7J6zM/mcJSXjgCEuCLYPrQ7EaxyUEjFONzuZ9Cb31HXDEA3lcBuOr
vG+gytNlWXn/w3L16L9x1GW0wexRbiFWiGglBjVic15/0IOBKa6HN0rHr0YuISLe
OQuKpFhVr59oZLuYQgM8CG7HtcT0DZsACBo6W6aRfMTWLXmZd7em7fZ8woU+XgB+
sDExap+yy1wMthYLgmcKPzYp6o858ucY85MDQ6cRFKk95iMDTTxKgkyXCCORpZBx
CTkeJeQAlttumbTQtAjrYBuYBYAjDbAf5DVj39ab45ZGhvPBodO0rXP2hSmpJgH4
BTWUMToVl3n24hFbjoRW19AvxfITIPctEVxp692qrOcwhTlzpDtqtXq4S5hNQv39
AId2UBkeDkDPNkN2ZsRfdcFS3UMPca5uHnPD5E93ElV0+kyagX4Ogjbhx9hB5eGj
hN0RX1CSl8e3QgARMhwIyJzcHGi3rTDsdEFaEfxC+QO5LXxe3yTGXZ0e7ovipsyC
Ie2qH2mPSmN97sY/ZwkQCQ4AJ7rMVTVuhfXuWYtMKnoY4VcmuIoIJOYaYmSfXqGh
on63jryVq3sCneLjc0nbox01Fzm7/6QFdzDM1U0E8rXlgvUDf379fAV/cyrpE3+w
WH0YbDu8BhwWCmXstmDv2ht2Gu7Znzy/u9GMx8ONAK6yUf1sgplTQNNXqOFQuj82
WeybCDBK5IMuh4Gahd91tTnhMjxpugRIk4rfd6RIB2Fcp1TUxYt67QSP4OhnFzTl
mJ0R7moHU9vOj77+TkA5IrpDwqtz7XzSgfne0RR8go2vLdnTVBTCUitoT7XeQUmy
kKOSeLefnTrz6/j1U2isw1Ggnf+AAL5ZPH9a777nwW0aS2ybT0s5YhOTsRnLJ+J6
0+vfGYgdTxY0Pvi2m62qaISVodVY7QnJfUz6ov59kzNuwuHadq+gCz5H4Ufv/qZD
VN1m2+FP3NYywiLFDKsFBDbN5qCZFsDGgWq8MQZuGWK4PLLANnNwE/uFXY6p717E
9LQus6pLSopSusp1V/du/W+1430L0WtTSifRqwjdb3MOxQA6KQiFiUar1cj7qNOS
DpvDnivuRxSsPXbI1EADdxZy+Y+/PvYMAnXO1lT1GZeP69gFRC7fKP9KyltkOlu/
5KQUYBAZcfp3RbVztboFTfsUYyeFcY7O1pc48R422RZ7VGHd+4UfgaUQqSonmkLK
4q7DmXOiTdgqJbGVdkTRgY/iX86q9OQuLrRK9RboB5KXoO3QSeUpkSgj2flKm5XT
0kAKOERaL0Gbm9eUvMuaBdpNjv+xBAI5LkbF7S93lzBhy/HhQf/JSbeUDAhziGMH
9NkNZlfINk8d4J1Ge593zT/Tg36IBwCxwEcVMmsWOmvo9KReUQ2/9hJpfuimdx0Q
k0t2JBBgzz8fpGJLKDAQ4xanCvnDTFBe4eaAlA6lro0FZHDQcSMg9qf26Je5LFho
Tfz3D47I03YtYVb8hnyRFs//Dlwxc5mwKLG4+NdsrvwMRSfhgvM+BUEui08WXEGX
iiXTdqZ/7crLxb1gCEsNp/WVpLJtADw+zQjRtqfvbtgaBEVA++cfCCBx+A+itanz
seBGcaq3fTuH+rP7GUAsUfjyVcEUTMyWkdteop7rpt+RbKLspPhvGOpB5k4+MzpN
UwEHj0Dc9y/F9hup+CfoV9UyhvTYpzCvKXM3xDK9YdtNNRMnJNFrqQrgM7Is7uGQ
qRqpV0kL/ouIGczTJwqABwFNx6GPn/vM9wRalbZazP1x3nDM/vRlo/QmnHBk0nJ/
oyZAIuNpZlrFnkk2ebsI4vjCOKwOrqWKiF4CU+Iv3W0Fbx2iHmebpnrIvi15mnYw
IjyUlsmwwAxnEP01aV2MSdYOMxyfaPP/ggSdWYGWlNOQe6SgCKL+vJZaN2T2R19v
lMfZja9wvRsaakXpSBWWOmUd8GvuQacnHsqwZMMDZmusSc2LiqCMdJmOMHoNhbl1
yX7vasCGGWrC2txfORSJqNZmRctF3g9994FsY5H4qwzVZLET68O0KzdyHE36LYOO
O91VacrM9/QpBR2aqrXrtxYljSOjwirj6sdMrYfu6hAAzeuf+FdmnzYvN7BiyfMg
+OB7tAaBdBSPYs7xmz5dmuxJ6T2RIsyO95xaz/z+5Uf7LEdHDS35SrcQ9uE1gBNE
0fRPFFyGpxUO3bRN3o0oPUb+R0ZUrfSUD8ZmTIihBsEk0JWOB2lEQcdCvSfsyYTJ
ctcIWtBgx6iLNM3TtdjCENjTuxXv20FgT/3y/1Aa7Lukq+Cxj3eJAYTEjrqBdqqG
5cjG4qqMN3Q/h0NL2M1ldGpX1UoX25DNdkgZ0NOJgPuf0tdwO5z9ASeLhaJQ1MK8
eEfeoU7BWaidLg0qW50aHXyRPXfKK6/zSZ6ByyINSyvgffw21EAiwcK47MtyeJfS
UKJcfUAuWpbUWLPWLBTht7KqGiMq9IfKaferNwTKs3J6PIWo0k1wQy1s74z8hANK
jER65nrNoQTpUdgLhqtfe2ctgbBjLKc0K+XgU9Zhycs1aFBaVyIn3OVk2/ZI8i5/
hSaphBOppjXWm8oOl5v9wutQq/fkEHQJO9xA435RyoMsQg4/4gjM2TVSzsxyXPMc
X+vOWkWQAMhXXg4BzIdFCs4cKjo2U0t5f5uN+Lf6Ua6LGS5yJqOo7pi+vxD1ueHT
CHihkT96j4ODjnW58S3cFeldUnQo55R6NeHLaCsFd40VN2MTTeji9TnsJGqir5t8
WzbvVKLUZt6CSWbpncxnFdOhqR73/xGPrV1iu6HfBoQ5IP+E/c2vzV01my1/75iQ
n0JViebVGHU7JoPyKWoSelOPrLvXGmmdwMA/e5T2Sv+BDvoBG7AWBe+eundxEoRG
wtX14g1Q2ZMMJ+UhESImQAWFTzBNy6aJ2ImsFR30lau1h1r/wkdu9N87sbg00wzR
Y8BCj7przghnfXwoEn2L2KXTfR+iI+sY0dQ4vX1QLYCPFyXHCIrmMXHw7yzODvip
sSKoj3PLMtEW1f2HW7d59UBDZ8jleJ1el+s5oPTJBWdWstrS5aJsYpkRkI84Pfw6
YvC1zo07YjkL/YXGwsYNv6KodFRKmvqAMtPHHOU/IAVhE3YtZJlN94IaEw7PNLWN
KEs0nCUWWX3L2GcTfOOOabYojOSai2bjNqlXBZcHilK45odXLTyfKhxmYA/PFX7b
4kJJQqjdHWHKtIEKwC7NyLaGfFXoYLEbX6vtkh3r7mW9CeinKSgF8lUdAlmiVPgv
oDrIaPl/MwNRrNINVRwpVc1cMtVgZ1QJPvDuqaoMymEKI78WOoYe+avctvAAtW9V
B+s3OPf8AnXbT6fTx2fgjkvtGbKW/HjJ3BQIl7ox//5FggVvTAIQb9zOw9bFsu2C
GkUE0AJtEUkM9dKwTJeoE1HfBhY3Ht60qpSGcU5lNZRqUtNjixeupjXM6EQ4XWHZ
Oagbt4MPEbF8BnXkccT4ygwtagMyWapO349JnF2biOFgMF1Sm1HFTxT5le7fkRRp
oRJiJpKn1fYnl4IBqWRfwmB3wTWOAarXAPKvn1U9UKfvNVbVL9kenSieCOBmgRel
nOpNPv2bwSmC2/Ywb2UDusk59wNaEbShFVdyEfO3CvwslWt4izkhUZ+JINdLAWez
bMKsOzRP74gsISfcl4OL9ksvnMrTzB73koDRoFdwaSs7dEqqsYxMoF2Hw/REhKrB
2NSoLntGxyKiue7m9qWhT5s+UW8PHp/YgdSWaeaifwvoLNLXZQnYJjjdMszYSzoG
NUUHU6R3f+0ZIBFeO27UPOmqq+JDEtaP9kqYwAu7kVpCu/sMQAIQQ3hnRt8OLxhl
U7WDbUZ/LTjEqJjG96HfEeWMyDQhsozryEFNfPGObDt3VnkM4tNlN4wOUv9DYHS3
o0ibG7qwm0ZsluPm2yJ5Cks3n/YA1eguKY4ekcQLw8W0hzEjnE1x3lsS2PD3cWAZ
S5KI1ECVSrNOAop/HA6yanFSKcq/pNYCD5eBo8FB8X8YGqzqF8hulWz2DktfE7d5
p2pRaIJTd/cvcrW9vh4dsKT/7Ydj6nzhcA1gEysKxQMb4MAKR2PDeDrciBfd2yoc
2nWAYLrADAXoPbeIMc3hwakN6IossvrpuRk2p08C6j4ozjon8/PcSJVYrVwOVLFy
QCgoJZA27PalSt+L6gC+FYcN6N0H/OtwDpdd9S2KRkQo028/GMFRQMCSvw8YhIS2
JXQ6IiWT6pwFiml/NnPixo6wSiskODshbl1VNY7xSiv1T8kGPDD4cB5lHi9HgAmI
vBUdVaJ4CqqiH97O65RufwuXttIJ12ek9mSDMv8E4ezVLDZTVMDqoDWfXDRZKEbP
wFHrblaMZ1ocDqDE6waY7/tpkBV4/bajb6GLjIEkFBktKSB05SRA9naqX4NAg8M0
XUpUmDK6Fypt58Z61mgMmFz6M4a+l+0qfjYkW3NQSLLG8bl18s0/EPoXgn17/KvY
Xzcjydeqf3NT5JH2s/BmptLQqEagXl183mTWcXNGZhJ9E4Wm11E+xorbSQZbGq2N
qT+2HGO1vvk7FqpiQGuC/wvj+QVq/2UMtrRgKRLBVLQSlI+gZWG2fSEfdYSxtbZo
39eiA25xGjRRQpdd773TiUqZoIu8RWEa4ytDHN17me/HiFopEerZNHsZ3ohpFnPx
gXLDjpICtMHH9Ab8xBb2W7jyuIy8EN6J3RepAGVxXL7MUal5qz1mmOGO2N4ij1wL
bWZh38SJ3fPk0iOvjIStPHMqQrR9NUWs9ZguoSZfwjyQqQMjapMyiiD/sLfqM/hM
YVET9vIwuRa+FGRwxGdnSW+GzGNWw8VCFi8oTKak+OtypeZ8U1WNdzZmSrGS6i7i
KET9bL6kWn8FYFk07xk3F105OJfoA4NMyg2HFO0BlgffYRDiK0DMziaa6lrBKpEE
JTqg7O7hHwYMdjQVFsGu5QXPsPovYVjwpXUNMEbqb6hwbZgoVp9I9+RsRYAyQu0O
7E9b/poW62+1NlPGDcejKFqwUrwbp/xb6IELWxm5vMKpTDq179YPxkyvgYIsOu8J
h6q66V3vgJdE5+yfi5ygH65uoDxRvXUf10to2wE+fKqpTPYMkPydXqYOA3CiMKeN
/3o10mJgB5r3DAcAgAAvnfUK3U2lVdPrEgALBiz9ckh5Ts0rGaE69WEoSZA9nTJy
+c1vU4tLlpVsNALj+38YNmv+IoaHHuOKZNw4fGIWKTuv1BZgj4U3TqS2fJOMo1Ij
f83lqDihPdEhCAyWo52WFFMzI2OaM/TByYRXIpXoUE2zAB+wp6GXHkcMdE+d+PE3
kt7YIkXPeRphYRE10JkM7dq2xZ7KXR8hp1MaEIiNROOvCoiPoN03kxDSOxIeRqHg
Ap3240UEQyVS57LgUd4WjF3QAqdWannZ9CAZct7tn/EYM0A+dRKCQISvl8AJH/53
OzBOZr739N4v2r5RypjkIgJ4q8/BRS9Lp6B+C0Odqemhc/TETZQz1b944ninExA/
QATq6bkBY4uAqrgqK//2yLDnMGF18SvcxovUNSrdmOIai6qoo9mSEfwPtbmLMR/2
r1e0LPWZjOn4raU4+G9C7qNdZG6QeO28atCW+EI6lMfUIDcew+so0eibXfKsXzSi
ZG5wWceDBYY/cd96fUOY/TMGbJxflhIi/N/1+DBicoDoVMmF6pTj4385hJXbVYhu
q2e7VSgCLCtAcYzCnvnn+6Ee3nJEIUqvAkIxDwd1bRIYOgy9Ny1Nr9/iUxcDaGYW
kEL7Fx4bHlCyyUQjfQJIH456bOqxX8AAt9qY+otrZjzk6s08BDmGFVQsm6ZgONcC
LvMDli6czuCR3i/7Eu08gqY0T2AjQtbCWSj+OzQ89DYPMc9qGBFp5lSNQV65qQOc
tmm7lS14ZlZIZt32QS7vXsqt6nqAsldGt2lEYtfF45rZTYnepfh7BDzgitUMTvww
ZDBtIXl0BhfBn2QmKS31gv7EhfOI/wmWTsPaBfSjsJ9/jrbD/Msz5m0+bWTinQrV
p9S91a+XeJCEUkAdsJttjwllZnWcV6iB09/oXySJZIPOVZezWp/cQ5Hkp+ISh7gJ
n6YI3rYi6WDdXq7dgp8LVpwR2wiUgTGFdUDnEm3qUD0XapjJV2w4BiYYbuuhVtrf
D8l0K0C35YTbRB/sMlQg6f2iz0YXLROVugiGt/SeDM840mek/hZfzbLXFxca7nAb
8hXfRHtGLZc4EhIH3QKuR10SBONk1DwSacjyVjFLw1g6LpVhJ/Ohe5ucaA8gbF6+
6opn1XV1iPDCHnzboWzH4rNvXbr9keD7ilHd/HzDIYO0py8XqhkbK5XWNbfvl1WZ
DTBt5N6MHpAri4IXbcgh+1dZgBsb0x24oq/SOAIUjTym23Fg2/ko6xrp6hUmFEzM
539LP3CA7Wl//C5ITNrhmavk9iCwsDj4OYRtjVqKS3QD5rr7rqLFfs03Buk3j4nm
ssgIG4mQkzk3TuPBNfln5HBn+nOeRPqIzGxxiLb6fdtzYCLFfyIfu2Qo/YIp/9WR
092UIdnUB0hSbXwI19fFy1dUV2nS+l8w1oQzHYxx0l+3Fx8u+HequN2I2M1nmjZP
jMXs5xYlGQQF5VymA3aQjLE+/72yAbZrLccvV9u77cen3Hl6o4U42AVJ8KM+z/8G
R4YTNTS5d6uU+BpN3uCFc4b9F72vou5OrH0zQCenmD/BECv5HLpxLaH0ayIQ4jMI
ppi7mdyUpm7PGn9PqTMJQIx5AR+l+5odfWFr1MCQJ94BPngJPjBwUFEgtJJozxty
15tDi4kAr3RlhMFfOOiUI0e2c6nu6cItdIElM2CXZuk9QlPb0AuFYAKeysX6TjQi
4S7vNDyIxiVFa2p9uJ31qShtF+1xutFYuFaEgFHhk1HfxF8gZ0cthFhpKCUvku7K
M5PU/ukuWZFWvOnQjRTdsb4I7Jm5ZHZJV16ECvyQZn6ugoQRKA6hsCfaRRVQrJ26
omPIzAPqR6Z49Wz8AG6O1tLMsTRMR7//6ANkRwrcDOtA2jBElMOm2Kae1IZEyNEy
VxIPaqnIaLpbxGKAON4kJ2I4a5icQr5ef6xmN2jmxMGvukmc2UcJVMs9M6yyhVFL
cERsXPicgo1aYW+gt4e6ZspIylTLnuqAxI+6SrU5c98ScRxSDOHEOq5Ew3F3ova5
CzqUUFqK0xJScHwcy4ntcNzGwyzCJbTPHxeZzbB6f5AVySdR2+t5Cd5a9kBBrvyE
I1DNsAUvM8ajNGIXJjLKrWSiy9mbq67ekylLTMbCglQ06UFCkn1zkZr3VHS41oMP
qyEf8cX1lY7rOxfbAGB2qquNAA4dnE+NYc7Wnk2yXcMM16t84ZB0J7ys142UQoLS
bfmqXGMqFYizNWrzXNckBkkYn2QOCdiIwbAhjkz70e3GEePOBPTuVr7z3TIxPtKO
/LgHYXjGkSp2gzWbJq+/ePUWgUzR68CHlhD0Lb3i4dBUTsVRa4YCaxZOEaPM3sD1
f+J8JF76gc3G55/bg1m/eL6r6wD1no8VJXsWjD+zW3/kO3KBNTXcD3jEB6j6z1wl
XEM7veg7nWAdLt4PGckn/OoEVrjtsigoC4IfH1IVz8BW2S7KHj+8XfKtbRnrNgUo
GIYiyPrv5UGM6x9k1YDLFQ9GxnviCmHvM0bWJ8Mk8q+KUBMFqzyexdEjCplc6c7q
JP8CywulGBXNSfmTQNS8XXGacGTubaTUYKCcezp1Y7cpuw84Z9BoWFdZI6JyDn05
MR09BtHVt8dGyjCs0XcvihBg4b5DltfItPyNFmvD2gfDtG+f/FFKCy+vvaEnAd+N
cIMaj9LW8F3X9W8IlCfx5KET87aAL6ccRuzYsqOg90D8nof36T/8Fpa05OVJdHSf
/arlLJEIwmTlD/CpOKuE5kex0DwxLZ9XmO8pPShEwdOSvuCd8R6FgLIgDEqli/rt
8A3AMOUpVXg0Prvyyc47iDi8OylPUVepFlkdjCXScm+PsdQEyV9q9YERa2/w4IMk
sVeVVKw5gst06WmHkXaQq+wG7sneioiE6SmBeGNeeqQ0QH2QkEFkFxBjtMKMOLoh
96k++me+m/LabSuJT4bkx/Jz/NN2yNaUXD0EMfMeC9Qt3dCsSMmB5BLg+VY6cL6e
XYFY2nCLeULgm5cZS/aA8pX6swftkkHkgkMzhAVJP2iPE9F6rcKG19S/cShnNStY
1YZKpMPXKRad6V0DMJ9MJZewKJ9SUYnlEm2mPGTRWotp5jN2lqsOxl5gUELoXUqn
YIBng2hC/UkNND1ahrwc6GlU3T7llCVTA4ynLOn7KgyiIZM13A+zT622CHta/VAP
hda1atw8ZPfIzAgaTxf4yuoMRDj1T11iXi7RgsIoWiEekgVsJwoc66nnrnTmYPKv
nDKHKhIwNqqxtJyNO2mAg+xbEHdsX+TTMFb3eWZ/001d/s10kiMkTWQydHlKF2MU
Fsu4QImx54O80sIyNBKbCMUR0/IV2VD9NNfEmY2/YIJ53K8sbmmkU76b/HLjmUXT
9Z6RPWWla2rM8A/a6L6XBR9ks+WLVQbPePrl0Z+2zK89P3/CilIloCv+dK7KoNge
ZHuVnoi1kJADpXPAffjAmQM8pKZ8QS+WzsyxBvrvHwM2GOW2IcC+RqR2rfRfl2xg
ORPWQCYza8h1uxAkNsQMK7M5wVD6Pq34S7GIUxBM6xT4Xq9y7Ukzi146Ta46dTlo
oNrjyoSrE1xUuFj/rZaJ90IEWY/yqovgw3TLcL4EjgaEOPpU6kjEs6ibNphZP9xk
MV/vsbgfUvFyJsFCPUV0I1YZFOFVzb4mdQBhOkU7QuEVcVEWWo3zq9MXX1bpsNtL
f3YUyZoXrxIwtHpHrwNafrL6jbUqYwGgFW2fufB4PTNxl+txIIwtZ4pi/lvVwQ1l
Zp4F0Jq0EzxRq/8AIp1mQ6spI4ueS52pNlV0bZqAKQUM5CGuW+tXXHSOUu5FwEu7
IriGx9bHrLVw8S7n3ghOs2hlo7HghktHgDadFqsy480Q/Xcc156DA1lwNk3RkJvI
bu5Dvy3uuStNWWkFxRLyqjqfkNA2h66xj71m2ehEkqHIxFPcRGbyUFenRT/LmJwn
GtEnc3X1HK+vLJve056ixkSTyCGLCHNqj5w+KjpQmwGQJ4xyanuFll0mxL+pVdAN
Y7Mj/Wlc0FK/VbNvpekh3PNrRAJJUyX+PG0T38xsfVzU0ZGgVefF9eK54YdhYrsj
qtxTCbna0/+1PHlwGt1tWDAY/yekGniLroGto8wVa5L53U0wdLBvdXWLxKnyeRTR
72ZwO70Y6fVYrGOYI4CZSx3wfAVdKZ6Um32ilikTPIk5zSkyPljBizVvBF4S0DRI
w1pncqdDNbYnAQMS/FWOapZ38fjepzUoi7sV2J2B6cXm+CraatVHZYdH9jKxLsZp
D5RLUvGU+lsfpI1ZYHAffAndu5uWUn3IouHKeZk+QPk9U9xTAYdAJAePQtZjxH13
q6PLMIyv74DK4WJ69SOD13RADdvqQsk1lQ5bE3dTqy7C1XiIN+T95B/+FfKrpNOn
dH/n8zNJ6blQPmjljj0WSv6jx2ifuSP/FRqJUZ4W51iW2IiEAQiZkGkSZDlxvl6m
SKqNF6SaUy7TdylUvGvc3FWgjEjp8FPtFVrtTBLOqeEjNQRYYoXWK+LbRZ4fvqwx
xnPRM3Q5xyxH1vPnH3HAbkFXjQh1zkmJGrHfcbuECikHhObRPyxwDbbRpPAdr1EA
GemsZuAZfz0BEHY8NRKagyuNNWZZFvrrFJcUojJzsvPoaG9knZoUIca6+fnECaKV
PNnqVVcMziFEg5j3uMd5OjrhuMgolMlEiezKIL2IQwT4nOD92HKMjPAYoLl7wdiG
521x8wJv3Nadx0+S6Tnh7D8AkN3sjzJMkzS1T2du2U8MZx0n2ScMdqtOgXaGogEJ
QUJ2th77YnCotpZPrwKJBML/g6uK/2wLY5VtUTnavjSZk3aDHJuiyhr7jXL19qlL
zEXiPGOGnejEiBP7V9kT2j2YE6x6q7PimXiN/yj6DcNXyllVEt2iS8uaY9bwelq7
w0fC4UBtKmupu8gL5ISUiZnNke4cFDO2FrIxmvaxETdhQVp/ZWL718wTN85KlodI
teCS3EJqjihCUgd7EOCRZEnxXFlNhtw9/PVow+bu8SbkbyRBgE22oiftKtESCr2p
C6k/8lbTkb78ZlFgwtrl7h1OdGNFmAEvwSP291Ci8s44adoLH8e/tYJgmmjrDV9t
kdORnoVD6ZLGy7gRyVHk67DZY9CcchW8ol+tZo2LB8OXTyByLkjFLITGfAtafpV+
9elS1eYvxhR21zcuLr3K9OhyfRk+g+84Yx0A0r3RCrebCqMGX6VRaAmAQy+oN1tR
qT8lwl0pWD7ML/9yt+hsShkTUZewowgvK4QE1Y1RVlThD+WlxgtdyIRQrCyVtDiW
0c0nN/PYKc3J1oxXVh63uNDNjQLXSHjuPJ2kHDyTqQpi1H+P7PDDBBXO8WXZlojf
5sJQHo+cX06z46+DfsXgz1HgWdsHZ35EWUePj7NqhZ6snjsrjQTnlzCWUdulWg+X
t0Ewcq7oazkroWlbl0mO1/ZstR48SWB5QVa84jm5stG8p+Bx3EUGcgAHuhLLXF0m
G4Nr6/uoRS9O5jbjWiqYeJlWC2wX5+ZWdSVpBCvTIaLrqy4i2oeC9i0olWHqB5KP
JreSANcC6p7xGbB9pPbLdzv3m/jjI2bdTqchVRgy55SNQLCdPdM9/RVu9VRMt0Bv
Vb+GRMWkUt8D3KoDtfBuf9unbGwiMRnsBgSmm5x4ZiGO2mdZ7yQ58I7w1A8Q4zvk
CEl+A8Zr/irA9FRk6dMUV8YUw4ZDL9nGPWpdyttf697+AtCg1U4Uz2nGpDfl2Put
moSYtyUd4wT3mrXzpd2zbRXp1SuvcwYCCku8oxYYqmv4W4Mdk8PUlQmP8nLri/aO
M5ThJqNPvjC85LbNE6kgOxgPSYHEs5YYUgrQ5MnGtAJld0AY8AL7vn0Tu9wQ5UCF
BJV6+CAIOM4/2A2UZ+BmZCWeWVAMiReWLn4dqMnDD5vfAF2xo4EOCMg7imREEr3/
oVNhktnXFnMh3tvwlLjDxTYdfoZMUNaAS4hkI1KJ15DbSnAfXlJo95EqZFShNYTn
rIwTFiTc+CjacGrt1SNXimjp6PzqLsYt26SidGM1mLY9fqnVm78dUStMjzmyhAIx
NpGYgaJRhRfl2CgKwWovMJvuFsMMnEqn2vJC8zlTElmaAKLmCSSBJ6h7CGOJ4y3h
v6+iwFUXh2HMA1hHVSg6uCiFLj84Rcf+WzGTgwsBxabOJ7Jt6v25Ebv3L7dbRE8t
m6TcGnenW8ZZLesmwMsNVnQhYCQHZsDjSpcrdJuaNrTjqiAT3EqWxQpIaxvTbEcp
bz0mSmRPSbhRhNza1Zw2GIO0xGYOAnlZ/u0QcMsApk0avB/Lh4cx4dVOIDwyggql
6uKI5CG4r750/cF4u/3VI7He+9QrITjmRHOaZaoTJB79yOVuWC7kyVVN+WvH5QsK
1FRvvDn+eXEu+4tLXw4oi6dK7SLqmH+QI00Z7VYXn3ZPNqnRe1jxSZI+84dtsoGe
D1szylHRrOGNM425erIeS/FOUBKhVlECfcEVIYSBYlyTIux8bQuOcpaGy9c5+24b
JY10+BTAPdS8XFlVTxwCrTKSy1OVIKwyZA6FBf0bTHQ8NvevWUANDn5cr478BU7U
quXTZbLYx0B6ivoG+eZeuKqqP7PCLV3C5p2Dl0Hyz+EyJZqfE90zuvVZ/VtQozkA
lqVTGj31jxURKvp46CZCIlhnd9kDB4ueHw8Y/ryDdehZm1KLbTsInXMpLGhq/Qso
GDXnX7fP2xveh0XFrOM3QbWifZKUq13BhkPrbO8bxqWv+IN1hwK9QUuFoBhdHpMa
2pGa00imypWlUsPmBSTzOTHWPbH+ELwZfhaA4ns9GpJGt253+YEjYKkofCReGxEQ
yLiqg7MPBvfaAHFxBM4fVSzrzp7nR37lwOJ2LGW1AEBBUZPzbFKCK7bdhUq6zSMF
Qqg1LOBm0jKL/eH9AXqBuVdaY3Ru5XfyYNTsmc7yQY558dW8VYSvN9UeDhacottw
Bv2FCWkL9e8BxQ/MBH2msg/r+9a6TmK42tNCXsCfnkaq6A1hsoTn8SDvmPNAaJsh
3FqlVDUjXeDGdVJc/B9n612m/lUJ5Uim7YLHS4I3cEXSrJ6bF6gbSjuEIOK0Qp8b
Z0wIH8jSgqFVrAq9/oihjn0M7kLT3Rh8RjfN0bVO1q/DwKFufvtwpBokr//vSyYH
AdMcvoHWSvIc9yeEnAlP+1E24RtHdqTtzTpIsDRAK26CYIzwuSKfkNHItAoCgpBI
xLmw/fOA2CgCkbJFK2fVWAtQpwPrBMqgo8kAx1OiXRj2vtz/koxVm4nt9R0EoBw3
0io527orpGZTFtOhRRfNaQdnF3OBeFlB1atC4IAaiW59DM8bCFwvmo1uKZn46YJ/
v++bEDM/L7pGa5hVeBYUknZN/p2NU8CfQ8rJ1ikwAQYq4T5CNRh7Fc8u47IItUjq
GBSSHHRlN7YMsupona9DQZTn2mP8ZJ0GWHvhzMtTQZr9opn7Q108Ed9hHujDjJaV
z95R8YWMreFqpLeyaHF1aYOmiM4W22+dK11ZyXIENS3OdpogNeqn7xBRrbQAYguI
bzWVwGDQh2Uv0aCASjGPvATjsNkIlGquAty4E4QNFWFBtHKflLYRQlvA4cyXc+xD
KXalJ7FHzqyFVfQMBQ2h3rNh7K2Yr1KRyuOY5AqjsI/3ndMlK6hQkkDmMYtg4faW
5i/OvBSNxEXzQZ+9GxTUDsw5/yqpgp7XuxBkxnos2jgq8Oo3KUj1UYrvSe5xHQzT
aMMT0bYcQNAPQDiRJTcvlboMJb3LH5BzZ7mKmduX4sAoIo3xY3FsvaH4iAj5KhR9
tGr/mwOt0ulH8YNSus9PMpdPqAZ3B/OrxGHGl//o4ANfwBqNGT4DhWI/4MnIVxvM
l9AbZRQ+0SnDMjjusXmyhYRQ4xNL7U5F3qtWaivvidKpkkrB9gE/kLuCTwZFl9R1
mP2+03cALr7CUIB+UvHUAJe1Do3UInnDplq0/tK424h9njRugkGLrKkmNwpPvMcc
K6nGukEc3WZ6BGV2RHeFfOuTVGimFYnmqRfSd9Jrpt7hGaclajkWb6ybMUb7iLR1
MC/YyoDQMPLthuFuERxx4TGj+WhV/RzcPxtzpFcyfaoT2Mo0B/DTxbQGGY8pJ+Ge
oWwmxiuopPpTY8VPS/sAajEDPctPEMV3/ikL9Wg0Gx0ZA/l5DQ5YpFYAP3iZtCo1
4Aj/QE7o5QoZxE0xtrM7scr0TuzLnhYZh26Bez6D6vK1GZ8CZaoqAG7P+80IwGhE
Qty4PGzVLnGGsOOWCmGSUOMDUxH7jGPYQwaVtzAZLuFsGYLDmPfQBqlcVFN8T8Kx
8wcSd/bOvfkE+2VRpV1RCV1OLc0HkubGMyaXxMoirrzJYHtk/WU4hLNasWzqRvMs
iWm1tTmHzL/0z/X2qtJpoDOiAbK11LdbS0sAJ0JGL4fcbC3fP0I1kLyNWcGOOLBp
W1Wk+6raIA3WtSjEaJ632c36fiek25mpYi7xe2vGAOc+5aDRTTtaYFhc+YF/vj93
jgGXQ9aPcbEUdaxTqFLlWZXTJOV7LuMHRVMgXrxZd7NhwYEriaW8UPasneriy7ts
QvSsn6ONC0OoOkXX8hyT24D9y5G4tuzIm1n+9vJg6AfGlCIL+DfnfLY8tqil6zuA
v4UVHbJ2wL9mks2QctMdRcIelHHXprsDXhWU0YKXDpz1iZioVwJogw5FUXvru5zS
bCeSLGRt8H6srbLAtKOzT3CEKUhAa7CGNjvJ74pKHxrHcUve9HycwZmVwOfXxnQq
3hc+UK8H07nbIHtpyBvzj2LGJjhcXeXcZ2L7QcSmvdTTbAlMfnr5BHblWKe97Mcj
9GmQ5EJL/S14zrYD3nnL7XaRbcUy3D4zirgz8JtF67DAn9BF36iyGDMcT0xqEAID
cQk2rIckyiXWMLYe891nwU4xR20IDvVzhoo3MyBSmyWQ3T4tiR1i56nxwlfbiRda
LbTgx8Dg0qqBu0SdZlnWd4xrlukoZrmroc/7YMvVLX1XoUOmNVwOvVk/iM9eaKVn
hukmTKqHUjUoLlphSxi7ngfDC0/9C9xf5CfpdGvT+RRSQl9VGNQcfCuEvyziBtNk
2e+kGh34o0rigP53UcHHh255hfmNcq/YNyzhUscwBvbFX2eaFMLZmvCYpHzCP6kX
FAnByYNcopV1HP4sPb93800NzuJwHs0SI8XYgKX9GcPkinjLcU0S7oQGdjOpG8yg
MQcSRXFWFGSQHb7pRBNYY/tyfpjQphgLTEAHlWVg5oIZCPJKxt9aSjyyn2meNQYY
V1sYR7kD4MpwRhVtl8TqzWwOCQ6qiUdJ5iTn6ksowW7NJBY7YJOdCcXmJnEwgttp
xTMC+xwtaR+tJnxHVV0X/kuXC0cv1930d84Yh3hVJNjJblviPTDyYnDQjBkWAsmD
al2vgWAX11Q76PcYBiKhJAsrtMGUw4LFTvG4J5sXaQIX4J9GxDM9pCMqgbZdB0Wj
G5oDiBjSOMrbOTBmKKMDmqfRVY6Ocv38uARcsi0mxA34Vu1aW+sfXrX7P8+jPVQj
ko7Ma0ZYagvkAnpWU025K2FSkfT0+NjkIgpD25VG1U+npS2Os6SPbkd9lEZVuAlY
sYThSMtdAk8JWlNQD1KXg85tzgHohRocwb8itThPGQi3nyHSXdPuBumbq9YhIdZM
zbp0aTKnQxEIH7uCwDy2mTDrhUWPLZblSowuvL9ggxrCfdLhZiqQTS8fdeSfbuHk
BLTzrsNSROnfQG7xNMDIBkdi2/FDFYneBV04d4Ltg3dde3ZijHoSieWaYgYL6uEw
7AOmMRE88HM4SMPqJPWpo1Go1BD+JMNJn3YQLtVtgSdS1LzeLLKogvuY93wNYosa
HqN84fmYIaR6mdcnBWrnr6F6Xw3uOyHK1RDgWl7wTnXC331Dm9bsmbSGfSe5PM/B
rryvcCgieNSk/d9tX5s7o/dMI68GJtE9PaPfls+8c2szb9M0f9/91uLLmFcnDqKb
sZZJBLeb0N4GIDD00VLtDpgFNHlAkdudpCKsnNKKxb5be6PaTqBUMqolF2ieoMOE
LjOv0V/Uh0D572dGwT86ilyzp6OvAX4wrb7XElr6TweY/wNo6YT1RF3sB0CApUsn
OU+uy7VAQgODyF+Tqfzw1VbBXTfO7dTcsMlnMNTi+DXH3lTdPP6gZGKBJ+DS/kfH
sXuGEvbOzW3nRHlkp17W9UKJCVkKsqUb5GHPKccV6M9HlmCTtuDVzOaYlOelnocp
msRtqlC9TnhRGs5hC16O+YcIqiWncNfMdiQxjPIJaRsDEQf6kY8EoxWWVVWyCtiW
QZARQNGXisabjEGrevKJo2A6/DrWGMMUKE1FCfUUnVCeepbrwaNh8t5Cc3UJYnV+
rPEQMy3bnYjiJBCwRFDsNiuV06c+IkkYtryvNxyK536nbgH9pzQGhaD5P6LB3udI
Or50m+f9aLLkBNmRTVHkmMoLfakB9fxIPgi2sWCXJiPLZ+64c5Ye3ovJG1ojmPvj
RkKx1K7pFkY0GsW0FF3Fm8YlGiqKyp8JfKjmT6KdTlgmfTYDCP4ATc1tljtxWric
WlQ+/Jg3El3M4Ckd7rG1ZTY9cYOKa3KxxbAiTOA3E1DupctAIzvmmeQaTiKUB57v
uA7AXkBE81WpYw9H6BK48FwAYNV6cEHx0yKVF3sJgbdZwEnjrI3VXARgBpBOifHA
xnvAxePHyCBg4YOOPGhmGiREc+QqWBzSVnOJ5mDhsGaJeHpj5LG+vrB65xzgGgxb
bbDx77B4TBvdefn6pOy3YMp9SgyeH7TEEoStBhH7+K03EYzPpNIQuWhYEFPYX6M/
63BHuxib/IPo1zA5m/y4tG5J0wIJ+aEratzvxLnlYo6Sz266WR5AwdyDuLtcJzrB
5R2gJqLOGphM+gd9G2xI2I2tFeu+pP7+ice1c8EMnA0whjTh9c6uAI91uCFe5PMM
92USMWrSi6gMa/9VOzSH6sOWRZwsApBooupJ84Oce2EVASbPhMxmL2RhTpzjfcqh
xWsSygwSitg8nqkKiJqlmw5g9cISivDhS2zy85GvDJhtEguo2ICu8DdW6EPCSZBw
Cw/WsyBIHUS5nhXzDet4SvFTttep5O57ZCR0XohR1zgtfT3hswBRYK4t/tbVr0Qh
7Q51Ei3nIOWiX90RgSDNaNUaBDeEk7fUSpd4we1FiUmE43tXL6sYOVCT9gQjvWHv
J3YKpKNjjsQkQA1+aQFiXy4+CBoAcXxVNlG+HrrFNKUmCZ4XmutNPq55PCGcMERu
mlgHPg2bdCm4ncz7Nf4Bs3vtZ5H+hSBNDpfAssmC3t0eMmZnLe680xmdlgx4MRmB
B5Otn4c4pbKV87CkJKuEKTm1RxOfeIm9OAEyCp5vtFtQIua4F3thKGOvKpRlIGsr
+x1zwzMFCUJfJb3SZ7UHiWBQCk9d9orh2mIij+Utszc1aFvUWLggT+CDB6MaZA44
3dXDVVAjFkYtL2lpDCgVWCoTtBDGtQFmd5ye5EgBqQfZUFBumvClliepTL6moqlR
7WYrTosByN2aP6Jn+cx9oEPEq41lCE26FT9cnfENJUflUc2AjVCgATVG1lGBuqVK
hnKiKNCUx0f+lwnkXwAGS1gli0KyvnEeMquIKjMiObek8hDavEuVnIi5IHtpCScY
8NlvqsImP7mB8QR8BwavvJJjmlsC9EpKGYc1m7X9WFhHD/vRv9Syzmv6ToT4bOre
jPzy8BztsF/tLjf81mmyTUKmhkHXv2IqWrd6DtAElS5Nj2JciG3QD3f6VT5HLs00
0n3+nW16Gwg+JkrvLJhoRraGL6ieJejzeNMFR+OtVlIJeygoDcdLVsRu/FyE2O9X
gvbsBFR8KeUxtFqD1JmxW/KqXnc10LAp3fcIQmnvDaHedPzc9NDiNVIhPcMmyA7M
lmsnyakRxcdpWIgwG4zgAUOAgJI3SJ/RHquylvLR7n/QN3CIeLxLDYrWlC6OH4gW
ry0w88ieeNSAUp2bLOY0POSYcY93HBYn4msNnwytIQbJVbnxzKI1yGTuN/GXlXjI
VCrcdLa93JlRBLfL9/vpo9v0Sg7vSfGVqDNa9NSStUQLhAIHY6py0ctrOxIVV7Iv
bw96I3SWWE9yEYNr92k2R45wpPZngq7HFHw91Gmf7bAWzR+xSJDdoJpKJrghII2Z
9yDxEsS5HX0x7LpuRwEd7LbprYgmp5WkuWS34a3mdVRrlmD2eRi+NNV/E6gYSxsw
mc/ocEA+al9MNxxZpLuUyAMXT9Vv24JaudpSk7N2uxivMtQb42TOjvXItfSUUjVO
jw0eDDQ4DVTsaUJ+c0eX4S/2mV46+1hC52eanWAFWDlESxKtLbusy73iiqlg2WqX
xQ0/zGlXlilSnpXQ2f11RA4mbWYlY8Q9zOpl3oSJgP1o1tPFp99F/dMryeozGQjF
2mITOdC59wSn44V+KAal+7NPevekdQjjTPgMP0KJeJNhqHw1A3Z5MMS0JKz/mIM6
YAUCfGCwTZ8nbN9YxH9x5HHZyUYwGwF2YqU+9xlssxbKYZ+WYwXI7//v66dbeOYO
RaRptIWP39lBNJ/ARV2ijq9enlD6Sc0ivVjpvF8hZUxXA+4Io51kdJ4Afjbp7aw3
mbqBYqhz1e/MQgn1Lskx64K4ZS0APDWMpZTOx740+zaDokHK/cg1Pc67NcVrRNQb
Za1vvx8r3JpLo2XZQZARunS6euZgJ4kPD//Ysl8h3UeLMY3xXYRJUA9oSMRI0bft
XqZa62JiipgBa5dy8FKUshfvmroT3+ttKOjTlCX3VcPqVXD07kk/csEie1iN2uuv
FqA2umGCF/nnimq2C1jN7ITVdrbAYPIxkrAPkrstB/9XtTFJkfy+XfqwlZh7exAq
Trsc/hhN0JznuWOu/q74v/H6fPyTuyyZFIGRu1J+Wit9xSRVSE5dJgAJtNWMbdQ2
WU1yd/6WSqi4BJsYuPt3yKVP1kF1jM/V7fOnUZgWjfwboaSqvz9KuQz/cRo+aJXz
Gw5hcROBJ2V99vjc9sYah8ffRz7cSQpTUiVngmRxBIB3WaEjMxHsBYAo5z5TMlsV
jY2ZD1daBRld3yatAqIRIzNgpme0g3wS+tT5pE8lZxiE6tH1f650J7fYTvY7BPJn
GmU9/XznCXQnsnZdJ1gqG/fnfBWuwnGVR5V7BdCJPlGn/u4S/avvycwAq01hPpXs
jkCjLocFMsKS9HLxpsOBOrRKh0rcfupObQxtvf1XitSCe58DTfLCXUODDFr85Hm4
PKS9EJ52HtkEnByFMKsdrFRti2WHEvUoLotGdyqhZSNIfJYfw5HO73eAD39VAW+R
gWN4ZCYGL6E+f/U7vMngfwba6eAw4tKcBSsu6HKS7QFZbSfqHBBWlomcIVbkm2de
FNtv9CGENLXZFea+xmRtOIvnb647iLSV8megsWKykBi1myVFa3nSJQcWC9Bw2zx7
MnN01wOPFwWELQi61GfuYnQLazz0+8niPSO5mAyG8eafXEMnGfQSdiAjfUrR4m56
hN9Mk4BU1ZMrlnYJvohvYgGyAs0cAu80gNUIWu0CXqomcuqKyX6WODzCcHObyIZA
KvnA1YdvbIrcsC30jxcZzdCNuxVz+SqDgqcJlYrw3ghPKK/73npi19z/rT+WypSd
9bOT/b+O4XzBIbiRGLAx/GkxwsC43sUzMFLcobD+FPPazDskdlEYMIGuP9xm3r9S
pgeg7Hi0BuimhOA7AodpkWksFz8T8ItHs/bZzUt7Uxx6ivuysG/DHwCHKJ5eDwDT
mlspodZbfgSj1LPM9PONlptNIQgXykLw0Qgv1H1tvur6G5r24c9OxZUBZS0naxBg
3MUU7XxavvqK/64bmy6cNothdHQ+f9pmq3Mj20OCKumHcuV9NeZp53Cc5IcxgUre
R3QvMVGpvctirU1lGxa7WPdO6FmwcHieftJ68rd7fOtrBzS2G9/enhfkbfwhvh/i
jJwEYTuw+BvAfE5yWwlIbZ0G6bs4TQCPCazp+P7wxEdtnP4TftKnfSgtU6Izqpfq
pJY58bHgGNVTBr9CXtSDQQ9LEjZJKyw/HEVIImItmK65xOvvZWlS80MFCwbya62O
HG5Lrax5gBAqwoBG6CjiBKzp8lfuKgwLt8JiggL/Ws9BoHnSNvZWtSLZHJbO00hE
XBObAo9dmmuK1hnsh10v+4G6sLbBFCn/ptJfELB6LNFSodT6PjOqAIb0/hygmSz1
LigH2FjzkFrrADg9u1JGKqgJYt+e98lhITDB7W25+GgCGQRGtLTQKEqogWtj7MxY
Fg5qmWld3jRK9qV1xH51bKVYeOg7X7KbHazloXgTaaFIGsrdae1fSF16l4Bj4OZk
V9AYz4wwM2h82ecK4rJTkPL3Y26ziKn6/h7bCtrcOXTabw1n2QvZkP5Iy0zbysab
s6QuNjmYxTVZiskHPv+hcz8h3FWMsn0Wg3lHbQhJwXAKTS9Y0kdurj4r/mhYJ3lz
f+tMNq6eKIxtwduEEL82GymSWY6YRuoXzEP4pW7AU9ZBM0XT5poERDlyWSpKf0YY
Q1BHISdumPtH4su99ikm9sYLXX8Hi9stCTzZ/9NkEkQR/tjbh9ae3hytc28iBb11
NsF6CSaQENfOzPKBRHaqiZoAEt+aEqooYD34zWRJoWBfn4XTKYuVzYEHBEZOfH2s
DVpCgOAAHQgnfTZoRYh8hZBdHIITB2GA5xQhTexqbwDQ1NOi1neiJTfH22LYCuMX
a9aQkHAunqttG9LIjGlvFlvD1aesRZWOhmjNdqi8Lgd1nGfl5uOXGX7SuAGWfRnT
jHtFCqObyJiC2UgHIRgZpQ4YJl1fWTrlxj8iU/wUqyRYhRkBoUvqg/R38BjHMQT9
dcKq5SBEcOPaO+6s8iU9RQTiyyuPdtce0tP3s7a3ocSA6tNA+VBHCsQDLPeS/5ve
Xf6Gs/Fl7wDY5qx2f7F1utmhEb4BGOj+BT5VIOmH4Ztfzw17LsSlR8Exm4bzzJ7i
QTIX9XwtZ6OP3x0RZUvRfyR9VSIXXLaSsAyg098qPLdW/a1XrItLHf6IetR6BebK
m2r/+++baDF9sivOEasrMXRcXT8MezpflqB0yd/xAHK4upXvxxlV68SnH+9eY8IJ
QvzzouUbUqpq3hTnTmxACeDbg13zro2ks5RAd31yND7st2ELoYDVCLfhISx8f9xP
vqwiO7LSqdMIVs3KVrFPOzkEqfFnAMpyVbqF4PXp20RwYfkaaObfuy1L53TIzpFR
baqa43KbO1aEJakfnqXsyAZ2gTXPYucH/ZHbTYtAdoQznZz0+yh2453WdsCT6Vqv
IpnbhqSV5WrmPJGgxL0ISpZ1xczjwA2YqR/79Qv1aWrHILdu5pv0bt1eGqIcT0JQ
K7Eo4u/HWNSiISrNaEPJsey9iXT7UmqJq6bD7qdC31v3rynszgI7iSRzoBY2YoFs
ppW/0MqqXaTQE0kDqwmekl05TJt/CZsQ41VrpO7z3FT3sisD2mbxrhRf2dSXKOn3
QhHmlzrd7Ok29EMGs5ITXu3+1E+OAoKcDMJiqD3Wn1UQhYhbOx/s1xdB1Y68rb73
9a6AyxZoZk8W5HKYNE4GG52hPz01aUA1U4mYc9VDEFcOnWzTa+nYyHPITGGPyj6s
GWpO2/a43qYptMC27e+KjZpmGPgtIfb3hQ4wXnDBfdnkB/avJ88KHWPYVdoEZHId
WpqxnQz4dOTV0CwkImPPIYkxucj/j5/zU7JxPWP+FZyRU3tacoGaDt7WLcS6n2FI
Xm/rGGp7lVvjO31vWax987yL6+mwWM78JxG6TqTFZDWtL/iIxGNxTVrQrU2vW6mT
m2OTHIPmsxFIXVyglXrmW9XmXcI/+HSJM/8U53USODS76A0Dcg25yDtrOGnHR2vS
k4VPiy7QEvQmfFuu6fQZ6PqZbCYIPGIMAhDge1VbJOuPDrfhqqsd0KtVAiMISgct
yOOb6dZPApIpARdUrFe0oGH8PkltUpvg54jqSLhZp47IMsSgGbG045eC8ld47z8z
duEsl3IKU0HkQwGJf/JZmSZMmvZfTIBNChovUV3JSTtDdJuZGhbQ+g98hWmqA/bS
X9Y7/AT0SvhvJJH5dZxQ/6JvNythMkb/7HL/dbR9Gkga7hjZiStYcURbNFjoetHg
Xk4+lrQPqRo1lQlJ7QLlwlRpyFBlC2KvXXexlfkzr+6++UD1rbi1Q+ZNkWgTRxLg
WKv3yeFCTrrqiiPfSS8tGQrlh3EwA/sfML79ZDsqrRXMW3V/p0vtjLhI7ctNpmIc
34Iqk0kIRU6jPsUxrW4T2Fgz/CxyIEvo6Y2EVwuITb+H3tOmfvzgWXmw0lTx7cmt
tis7nshZ4ELfv6PMrL5ww0XmEKVodPiIYra0WDE4TItZDV3bdsHXLn8Rqn/tCII3
EA/hPjbX8oo8+52uC81fhq+JIOgCN91M3APiojYr0mZWP27TWBn02r+GnFQow3/m
WAoINJaSFpaFN3PZ1JUf1TUTdO4LpJ1gLQlkeTGt2oQCHTuu6OwyyjkdbrUSeUbz
el2ckM8dNTQX3pLi/vWHTAsvYvqfAiup0iyOuhKOFkANfWikwiiNucFfnZ9APUxS
Wiy+63EFpHO7tStz2h8tAuI9zOL/jDysjlIQW+e4sLf90B6i9RhojAZStIilsl2T
W3A7FMEfOKuXb0abtHEqvqh6OVaTRhVWVvfJjp/0xVbYJBXqkpQP1JTDvpnd0H13
sueIwsSfyLyMISkykO7Fzk3h68vF5YQwTC+vO1L9oFbS62UGAU/0BKHorQ9gAid6
dH/gCBEXr+J9Gj7HSi+9ZBy/zIWQuUqYsPFq63txFPJBZERN0FGEWd7eIq1vwZkS
d5vC18Z6u4cVhGEveBy+THMxqV+kuAeSfIzBRh+uLQoRMOxfRN5NHhmLKg20TjJA
xqfWMCYz4UXxjD2rQ69FfqQWHMvc+YV3oB/7Jnog4jmtiHl8ZWHq1eI5rugIN/M2
Dy6gKh+yeYIbirMX8i7XPuphKRQLSZSu/odbyBicvjx7oZ2t0hJEgebgXvsX48hm
tvaop/XLwtgkkH+oBUCBfyi80WenatwxlqetqmWAeFA8dVXyDQCHnAGtyO18a6dX
77bbYlCNO7k0AKcA1EZdYiOqcM8afK1drToUmMQ5UjdTCJfDHUUGWSmXYwjYWsrv
vz+4SR8bdes3jRM1TPEhkd3hIDrcgi3rU/nEq+OrTXb/uuw9XKnAEncffW7YcJj0
lcqGszIlxn7JFSidnok05yXrVl7DqcydAH5HeaWd2kkDpZh0SKqF/41QGUq3fbA9
4B04XTjb6QzWE9f7ehAm0f72k1zoDJCa8aJauuHF2FnaHu7ACEIa3a2N+JafEiNg
3JpLZ4wCm+bbgePXUkewjrCBEgn7lOrhwtflGst5OJip8gkMGkCD3mmjgyzx7V5k
xCjcxcJprBL6HMUISuk9HvKMOUpy8L5jugFBxSqKBXfbYcIgTXF8dYHU8JLb/qj/
TBnEATWjPDnZ5pMoWSFZt4Bbcoef8uBIE7f68K+JrpE31NtzRhupIpcsqUyQyoW0
lWEgIJhamYfs4YDeAq1jcdRAIe9eXbBYxyK0LwcWwMGFZZq4W2tpIQNQq3hhmGNe
9559d0OqlYOg7Iig/vmG+a1KpwA0T8YWpxMiU00qNfPUeZWXHsGekju1JAZNjhot
yZUhQOOh4AG4L+VO6DCwOzQOUmvZYZP9Kphy5AcB/+g51SIcgCf9v5wGcRwlCyw2
g7VXi0R1EBzy0Z+Y6BRoFwZgAFrpvMe6gBv1XtSO6Nled95JiolIRvDsrWATzsUC
Er6Ts6A4wbRFOZx4tmMSsnE4AR4bOzJhgiedxG+iMcncrKofmM750cFBwmHv2fz1
77yH8hxZKeM6LRjIAGtBsisNhBp1wrkahTiOC3D73L31I1g3MdEpIPmX18zhc98/
AXD6N5sKF0aOvMWh9O8+ksWxaeKReLFYFIEnIbakbv7qpmpDBIpvJak4N4iYSkZx
ep9ENABvJmzO0TsUGYM0z93C6TT6n527WbFxT7z1lyGkVmBjDLoIhLgh4tRL0rRR
JEQNxmcuuCcXpgXZee3CknuG2d3dpnAzNP1Qw5KBU423h66jyBz5tybDGxR7I4NX
MnvAjk0imE4UWBMmoIzqNP0ve5bW570Yl+KSkQ2ih4RuX09FPGcBpuro3+qUDzaZ
4qEHT66aVvKDzP9dD2roOUbL1HgMUGp+Q8plWOcdZuNhHyVHmqia0Y10aAvI3tUy
Sx1YIilVzieH2MvpI5y7qZ30aiSWWMCIJaE96Kjad0rFAOcrE6bqzlPOReQ7ppHY
nosxmje5VAgF/MP2fWfJbd9k5TgecAKd1cv9h48Ig3XI10c0iT0xlLuTewbjM1xA
xDRHqb380f91xs7pcCS1jPaNdXECP/djTwfE5+eHoe8XMwr2DoOm9VkiuZoWONO4
W2uTZODUyxWDfQgPwBw8G2mNk7/9+dJ1LVT5REHmzii8dUIa7p/+mCuY5qR7D+NL
KS6EybqAcgsuoibe0eXcsHQD8KNoZNYvtJJg21C2RMUcSupW0hiFN0D9sEDTxa11
4l+J8pNPKnnQEZkyjfhhqK6X8ipDJ4inagAIVWVTMvQ4fjWBlNc2JhVVfCA39j3y
FLe6j24DMzq/il8y4bKnGhnj+bh9nyqcJn1/6tRSatQMss/rkeKkaL0XaxUqp7xI
IzzRuY5a5lu2plq/10mgtgI5FtXgmCmYaHQXnSN2dh3WQOrZ23iKUdBHjZJUm1sQ
/57f/xh4g95I7gVjavSsW+tcJfluBsW3m0H4+SiB5FXYZQ6GplyEizkQOScHDA55
U21BqOaX51dx52KRgds1satR0RSUcwCsmD/gNgs5P9iUCYnXVvBuwVns7fdC8gE9
cNg2TeEjBR1/mPsTOeRix2ISlb7Yw+4aM72NzCQQoTRKV4QCuBojF4ZDQYlbd+BY
jqb91Zo0kambrZDLLkDm8qWv99huECsIFMERFLJhtxO7YDj98Xqs1QXcHnlBvZ97
ZmAuKRJ191Gf77aCWjQozEzfnmduHdQzyNOGlBYQoDGrr/w0/YFE+n9/aJbow4QI
WGrSPS5rWuHQypDszDUkY3F8vD+Yx/irzJtchx2Hg2ah/yykbdYECFT8fWk0ZXC6
gy+pdHWCutNX15v1oe0n6aDkszSogc2slcaajHk7UZY4t1KV3lvYFXYRXUfQ8VaF
J411BSzKUMi8ugHHALLXlamSIyqYRwULmDeLHBDmhbMzjviogOFGdV+8NlZ31W/S
jKKuA/7W3Mqk28AqYMFQn1lNwLx/socU580DRYCGtocCWN/cYYnTT5GW4qzbuT6g
lC1SI3epEGJ5sLI2ciOFGgRdDGF1bHto+4bLFrFtH6eUL53n/FWaeLAu2dOmoBBW
mOuoHTO0SqbUmmKTXkkiyyfX0U3w3nAO2bdrsNThqMFS7oh5csvFd8Eg9h1BHDYW
pSi4KV7/e26l8Rm88d/bvjyuTFDdC+upPce3e/OvCLYQ0qoyLAku6gBEyGR5oiEx
XbwKckCTjrgX0N7+DOA5Enjlg44W1NfEoPIr+rx0qZAUvR1o7Xxx7SIcAQK/M8Lw
iunoXlaEXUfTlSwhByxDIjJE9bKV7rwwJlHRBs7cqUKDzrPmbabrMuMKtnuOn1v5
Nna7T/9MmDMI/O1PXPnzHMCqK+810kQIz5h6rDh6byZdLPNTrFZolHRNQdLKmvtG
j4S4Ri/scIA0Dx+1HSUT/hcRstEMfdVMuWPbCfDe/PO6FhM83+dmescVHnfC45Mi
8sVxUJJuS/8KU9bbBdnjVBp9KA45hPmMMkAJ1ItnxI+qbhirvLr+U0BnqIS9BOd+
M8+nRQk3CiBupsk1UPIUTLYdthfGGGUSOnx15D6esMLYJ/j9yIVDUkH6QjbvuAVj
fJAyjETRn323v8Lh/6YHphgUBPLx04py3ObAX3xDKE76+yxIQHREPZUeIan183FU
YPoXa9OLpI1LLynS1cmP6ooQ3Xnm0VzqgFNEQsRunJGzY4VA4sfiVY7o+oEn8y8s
My09ofWwvF2qHyT9RV7hI9ZKUVTA6Z5o0Slxdeyhy3bW7ch37GtzxCzA1O+dn2Lg
Y1Q0le4W7HjDbSbIFKVe22oPLshoePY8xqJK9JDmjIo+0nTh3Km3vIgBSPJWV9pt
OVKHi2cnOqJ1gop17HTZGV6uEsxfvKBhvfpEfUL/owobdulp8Eq5VSheI3YhC4NS
tSCBGXR/v7WN8UVxX1oOORue2lQZ4c1TL1ZhYn/UUYMqNLL7MP+dWCiElafdleg/
clMZj7KcoxgZm/HnJFOn0ArUMYMkE31JbUq5x3cOtMOGisoRoRIo/uVlbz4bCSp4
U77DrfVT1txnAXD1NyoGILANyXX5ItDd3H9zy/xy6EeO1Fs1yxZF913xX5ix2Yq9
WO9TppUcDGUuic0qSQj9F03XYqTIjkcSWt2NOWy9LFPZJZBuLIlHtn4TtKDGWHjQ
ZdhDJTrOXdX9XL0m5odqtMKJ+Z2O6/EFGa/GcVvg9FqJDIcETaeSwUKg8MASDdZS
KzfuPDICjhbJrn1usNY6UFzX7JmxeSiIJihEpF+vDMOY5h5KwbHG1po3YEIKo7Am
U8yhAttMlpaA44sQXpa2vAhTq75+I/s0DZa2eN69wcI93UOKGWPzMUgAGNLbTZGe
DHN1Cl+BFAIqvkGtL20XSZ4b4XDzsWNP8B6EU0gv/SFCtfOj3+vlFCKIzgSYUiXx
Af5cnmLFWPaBmNYyqwc0k5fci02AQJiWNkOhT07s586uX5CN1Rx5P8FEqrrv4OZI
yAykt2/sYWzPsPHG+peWvVlTKH9SNdagL/OwLpovwfxiGO2uMvP80jzQswimqsaI
osiJrOFOa9lKrY0HRbJDqiui0B9vcRq1WzezfVGB5zOHDcuPVg+SnUl/ngfKdC6r
YKDRsr60KkxybF4WYCRiJQC0Tz3DYJYTyJkm+Smx9fruen/q9zdofrCopknBANM/
RQV7FgHe/oVqgdajW+ih0rwhYwWvl40q+mk3fydjiRq2yK+McAKogm2nBJtyDaHX
RPl76pM9D/eRSuJtcOnpcurMF6Xx+CrQ+LwERezf2o/qOmS19mjJZah6C5wSDDmM
JyG3Gny9BgoPWvJYSxe2TBarjoKdQG9fAvCpFXewEQZYr6uSdA/mSXTLi57i/BVP
lhXqUtJM0GUKQ5fXcKD5rjJ/Yx4GqxjifIMP4B/F07rsVfH83tYBrOq19xNvxiAx
B8p/K6XHjweM18OcG3K0If7XhCy5lVt0GrVwgVm4dthWoLXEZJXx6d4OLavPx5x0
gtHMoV8aEsUmEN9Qnw/jtBiJvIReHDHJ9/pxPcuITKJUJJnO+7+ecHCYhBA1ikyK
TuPOkjWVVThU7SDihOdLc7aAmt89xVyoax0SsuGxM/BXr74UWUejUycwpPAMCa9v
h6zpjGrlRVXIf6rqYAqB368cqK2pVwq6Pl9M8Chyh34/iYddL6UZ/KXmJA3PJVsO
pYO7CJnRl+IvsXTAC3uInnzft6d5FhxTJTotjPafYlON+tvz/t8LKMmJHrtkomhV
cZJFsSP2ukLBLiQb3eO7aPzWkDn0TY8Zo+xUVxXMFjcbRL6IOXbVZKwSmCta2Sud
UivNAWJo8e3Wbzadu/KM9u+y39AGtqxyfkmCo1fg8eiHWtrQnmr3ALpmcdcAFI+4
/B+kyhYNKRRyhxs/I9sXNLuSDxBlR/9OG5Yj6+Dq1r8x/6hxk0fJryxuDbdkAwdI
gyxz9aCWL4gIyCL+9zUSWY6xt+CX2PaGDoyeAXcqucPUy6n6UdYX7M4uoQoTW5Kg
SeVrAFaKnxrSdp9008VsGlUbJmLHuYPytE61pQjwfDzStmw2mZ36FZxyzDREE+gE
qUQ87pPTwmVomNT7B/S+uj/r/itK4eqJ2aAYCKtR2PumM41tNOc0OeWZvo722Jp+
5IqsiFhXcEW+JLheehfkt5eQeNQF4jIcisEGHANb2eSvP95ypDlmlwSVzSNndXwu
NtwNqBkH7q4Y+BMnafPQ8nOEOygdbVzZRYxe3kYX9pBwXDpeRkmkhbvg5PpintKu
2VrGVRmlTmpecqHiOhhnRAVOlrbit55J4+zpHCqiiV6AAKrYce2v2OS+T7a8nKyQ
LC8vu9T4/Mf0ePrRXhCOo91ll7F0MIERUWpEwt9ArDxVKp+iJSd3bZ7lw1V4kOZJ
6Q0VJXnbdiHv5iDZUCzzf1F0eGnwcHzaW6CPn1qyA2EIMRadFDxZ1TOq60kofG1R
5jXGHncw6ULthzyTX4NTINEz3XWMufIa8Ijkj6+g6mupkMgQbjDQFrFnUkurqS5V
G9fhY/9WUF5UFbnUHWX65sMbMFnqZQoo69MaMUpeRnRaU/G19JbMqXnleFP/B8BB
2uJQ8fOByI7TnDtBPpNS3FT0+19STgfW64kx1zrlPDHPOMgbb7EptY9XFC3QNC2R
W4iuv4dNArjAghdVWhED3Y6nRXu4FNW3nWHYvjYRI2/7Rdbq3OAXiM/oZst+VVv+
yf+f72k6Qqasepx/jB99eZFnDGfFH+gBgw+8jqtTTMoFTpN3O2tfKW2vt9dBRW8p
sSAcPe5v3cIgOUxTPeuKbLOnt5zVC16QDM6/usptUrsxGSSiXf6J+YKrcS1c602o
DAC+RZQK0VXwAysIaH5k0k13HelFLggDAb+mjZzlhBpnmfU7TpAveby+IBekOmlD
mGFF85hNC32g1Tw8qbgVypzaDqbmaXjX1nNJFwqEd1phFD8IoompMJ1V0n5XY5Fw
y6LiwwROCRADnMQpJf7s3D5bLkgSwfmTDP5bOOEqxGajAbc2IRN08Y2NRr6H19a7
GaYghllXmPPaoXteYoSX9xMT+2/pvF42Jr2LHkI7hNKQPw4PrAKbMvi9LbppTDK6
y5PSFI1NGBi7qcAWCwmRLLc1MkHmjAFtwGD5lX7WIzScTT3qTGQkeUs/SPnSIt5b
rvqHOObQzvANdH6mtL8SoV7YMFrVaMJF84tzMhXui0dXjX/KsyH+BZe1L2wNwnZK
kn1RSDt62b1BOFwxLDZUjbjcg2iZqTz/lt3xo4kSuVHNP5gQEI3FpWFt3gCaldDQ
WPxAhlH/CZKG/4CmV53Ehjlf0Q53ENCOoZyqSQ0QENW0NTpRISbM/fxgBvu9zw+i
F18S+6Wg2wran2oMVJEYtbHikvDzmZs+Q2kOf4seCLw7aYe4ODe1Z2XfKM5F8Fs9
2CEHovz4EdnyPGONy91xQmMtOvyI/98D4CAT2bwEEg7oCfAeYoEm8sq0egaeZo2y
N/sZJBBDTtdKDzDDoCKkLbl86M0VUxwv0biYVmPOzMIe5euIFB4y6ycmk9UkCL8p
luj7zP2OcndZPe0vL08jDOqEAjcRcpDzWZZb+2fin8elywAVPqFxznLMg+KTYgh0
vRyefzK+DKr5P81zwtgs4aOMv9BiN769NOJoUU2++CFPwuBuD0BZYs9S+gaD0gB8
OCAEJo+3LpqbF5JtMpJdNRYAZoo29cK76HcGfVk8Uwv+KyVp7BPsm9GqQ14NUDJ/
Z/rNxPYJxuS3VrQBPJcmJ1pmW2tINv2aaudC93QfUGw1Px1r8k4u8UEZns6oltgz
Ql2g3mIvjevBwG2N7IiUNGMo/BbvuWKH7HN5DPEmeS40BbbsSFcZ9c4lv8BcsbQH
Unw+6iWeya0FqCyhtZeM78Ua5ZXsFuZjXCAJo5k7Ws1chiKXudDtG/agkZ6Swpzk
mdpuZ/q5bYYfU8RhEXeENslGpCHFRsgQ2sTS00+oXb2d9gQskN6NHO8qeqgV+Yra
Ygu2Gaz+SHliC0Bwh3lIfCd61mQWr6mDQyfrMr0pr0ZrhDvtPtO9DjZpXwi9wAez
deEnj8216Mxaxhky/fesAfUYjst3ISfUg2P2x78ggpADPSmiYagIyxiNvTzWRNSF
LnLRtD+Z566oIcXJahVEwA1VRCqIWpLQsKwNtp15GyHq4mnfIH8qy+oYicnVIbIY
a0olpEu7RJmuBNPBJ0gUeU5r7T9iOb+e4YyagjecuhZOr2PCRU7R/7aeINeZc+BK
ofIl77uboBYNnXymxcyulKf2pH0MjE1s9ztgPXDGaAc12BbSJI72AUfvtg5Imw3A
elOFOZrR9H+4H8kdE54Cs4pKgD2leFxpCMc8LW+lvm+dYsNqhl/MMVFd/pKWNMIm
uxWWNnI0XzdVpdIK6UGXzjpLLfO49RmSVM7X6bcoArgPbyzjzuXhq9ft7aF0BGoS
aza4xIT6cARz2nqX2RRqn2+R9egPQsxALrNhF1P/xR6WKwPFQU7ZTeJwq6LFcS2u
gMyhUhrvjEEjFQ0zHxYAK6X6PwiuWj6e5a8ZvA0GXt371pMShQIjRGJeYE5mDyND
F3qJqXwWkKJydJrop2XSP7hN1I87Zss7oDG9NpWT2jEELbtPgwhi4QIA2HlF3qQQ
7fNgi22fuvxSwY8XwmroYSCQhibWoz25POmlO6XW5VkQw7l1S7kxa7yQ7xDtr/cy
XYzI+0m4jySt3ApN8vbSMYsCpzMjAdS8EgEaMzOXqVLJI0MQd2G+d1IWOPp6lOm7
h7325sJYhz7K85xPzVvZJJ3tfY7NHqs8Ehh4f3P1Y9Xi9nF2ArngHs/EkqwcARCC
g3a4X4vfZArTN4tsfmTxciGjZ/vnFhzxab8DlOLhKMGlIOp7XRt28nDpwziI9GIS
glZ5Ex0OI+DCf4GnuwVuvZ2vZL3jLXCsVn1bEwCeKc/nrnVChvxXWn3h1C8C+VdK
mKAThLkpnGmB7vMg1KsppQEhUUdnoUVDgkd5ZxNZB2/nh9GGOGMpXKkR1PhyBvhD
jR55hr310yj8HtB0MQgt1IdXochPxeobveAfG/8Z2pZWTQQLwka+pkLh8MNrMTP4
Uc+yjVi2UWT+3YVujrJQ6L6UEBw7lyHEIXPD9iMvOe8Cx11NfUsLMwk6xI303j5t
0dQC/88ddIvelvtmjaef+igqqHUogiPmjjqr1qAPqfyPWHgQvjdRQYgCnO01oXVh
GT24wBSQdfRlY5SJrfSm5fbiviGTWlH6B/fAHS0COcWbxk3bMxBpSG/hK2LoTOYE
1roGWf5I4U7x/FyuogY2c4AfYFy4myqc2+wTbtnDq0DIXArW7zLDN9qtiJy+dl6w
VJjDBGvCgFhw2bEIkDFySFTv/SvKSJtdhzrtJy4vJkiV0YZtd8egiCtJeoNi+6gD
xryGSnjUrwunRGfad2GeNvSsOsatMkeHVb6HVem1qBSTij4+ED2BXSEkG2aCJtLk
jJ1A6MzTFPWGgCyccXDeFnkVpa3nZEECYxNsjzWEm3F393WK0WoASkxlkiPjyXP4
Re82qPqmgWkVBPFZNl+myPYlkrsc3PX0I7EMnI7K0Szbj20R/NujcCVU+ooczfeq
h2/Q4IMlruCmiO9Kd2YHdyEhomSSqB+1R4l27HKgEq0mXuZKORZ9bvZ1HC7ezj+J
BDo4wVhjGcvHYfeo1CXEM1k1niRvBgMR9jE/V0JBeZZ1tv9h9E5FKpwfhJQstxfl
VXCBs6QlIIHnqQgZKVAaM8zJWK3kyHKLtERnUmAOjF6A45d1AlbzvoG4JJoGdy6U
rTsJdmT9Kez7fIPvy7LqQh7L2iqaP3whtLKuJ18cMx8k3VlmMZ5Pw+OsezATnY7d
Qa6en9+vhtsQ61MNUThFmiACljmqZ6ysARw4LTknXo5JTrBu1mADAT492ALbEOwv
i7GytFJ784eZFRlTbHcXBcQIf8JGhhN6Vr2nelJMbK2wyMjk/I0I1LCIoBjBxf1i
v5kdBqtcQkybXA0DR/xwS7QhRUzVL0a6nBroANJVjMjA4Q9/BM/zn7141HP9cya3
nzxycThH67i5s5xPbMCYZ6EootROwFMdat8RttPTpkOc94PyNAxT8thJlkF6Xm+i
rOFFxtHb7Z1/FzpzcvCER8EjDBNCkiUvDg8NTB+zvS7Xxm8QZwRsb6yDUj1UIgp+
SwiXITaMO2SZoteelJnWiajnNUvpoRY50o/AHit9j4sgMvPwCQDTl/jpXyCf7Jip
VhlcU1jo6aaCr5i5UArhvUuOc5+Y8xvkS9H0Wm+jaYKvtK9sTtqpgMwJjKY6yemi
4qHYK8rqeUPptuIa0XZN4C2UM/3Ww/vEow8jLFm04axpOei0PeJ7M7WGiix2w+7T
hhJtm+Z2zeBKgBvc27Nj5kAVEnnFm+C+l11KxWg0CO/Av8a2NiTD7qbDPGtWuu4P
8iXaPy87BNz4GA/1ZBi0kDQRwOYCAfULqWZeosHJQfrGOqhb/wi47AzZPwDpy4dT
EVHnDWS7kfz44ANDdiOtFGinSzOs/hQuteh1KqnKK0CtXRMKlrGT7M7ceHwM99kQ
JB2sa5yGjMm24lzvVU8utEu2+DZXY8DX1CBMbAdMI2LSbzenWHdThhJTHVjXI2Sg
Vj8ejjsx/mEG0zjp+Wxl5r4aBZAgMm7dSycFjU51RSSc89hDCEIAwizlbUGfsAi7
yp5ykPwQ98PPyLk/0sFMc1P2CpZ+itE36JtjHpcXvDvYxSWoOwTBmHfa+R6L3fPa
LvTZ6H+i/Rvde+hnMPhgLKKxnG6v9lArFS/+wbPx4vRGD9jjpzWCNIqyhUWMOuhB
xUbzAY/OMUfLo25+/osIfz1701eTbBhz236V4uhBAfQ2km0gO78m91QQOd9AlfqG
GMiEEPpBH8iomW3fHdTdK9Jn6rwuWqm9j31wNNtVR3hGhGVGVXqzzKPUv9mmIaWp
JtPzGbvjbTr831RyWfXZUMW8sSEnh/Gu/c6Ic60NEY01CaJVQybRiNhUpwImWnCQ
9n5ADiEYEwRSSKTZ2SGtsChiz+fPOJOUuOSlVYVaqKoNHpgMERw+AOmcBYfvwREe
cEWl76AEaYpcjff6WVn1ASpa0T0muDaNLfkyjMPsuF4MDu1qj+/tKOPuB7NuniBp
iwBwIjP6EIXJsBi2TcXprIctlQnEfoNnY/QLj2UQT3L5gKi7dujbkhmgPTI+/OBs
JVuMZ70mRrVzJH0V9JG7ufDBMs27SHYwS/P8/dIcNxSNUoWKhFsvKhJbtcNASIKw
63B2tZQ5l0Rhp4+y97HqCMzlChb6BZhPjnAGxVff0/FfDF6b3QI3WqIRmdd3rB3y
aILcWVWqdg4A2wxnxkF5DZp1WNjos6OQaYwUgjhFGBRcL/SB928mtanxWN42fDYt
EKMZr9u7eUJUmhma6zJC55oPaOUuJcL9mQMwVq9D7wd54zEiayj7Rhr4sevkubnd
TLlax5IgAwZtTuavuiBf+ATXnc/2qgZ1+5umAujlcGdwQCps/sY+OxsGklna+wUP
ul4Ry19jQkFPidMq5A7Fz2gIsXs4AqCHNKTg61Wex9G88nPoawN9JsZLCAuNBSpu
iDSFe/CF9OTfHnnbAoLKb/+fTks67ZHQF7rCKSJTtT49cNLS1AF8n4gAK9NUHv2m
bKzmthl/Qt8fduY5zPsMgm9gxHTD2YvzZBhha1iRg66kuNeRIcEIIdlVsu846hCg
LcAdsZ+x6hnWA+oN8WenmT/Yd2HvCFIiYN/TV83zUYZZplCkB9+2dwmf0KLgLtxL
OGNosws4iQ5pyduRHpamy/nTc9mB4XYXDQj1jZV8c7Hr2u5qAYZXnC7EbnO1LqEv
4BnxmE/w/ubTs5j8PC+xERF7O4trCxv1KKwR5vtCkVykREsu10ogNPkekvhBR8WH
o7e+YBvpxHE+dzcyAgiRk6CvtajGYan2BJdwglbwQnTCB5wVEqQct570Mlq0Zfy2
oKPFPl2n/Aq92awR200IFhRvF/YDdK9wXJGKrpsPoSfCT0ZmWl1mPISqNA8OYkiK
ixMzpR/uxPRZCunE9oRG3qjJE8H6BCmbw/LcP0LSlFfHKyS2fCZuwesBdNjaHnQt
4lKpRfPoT5YrrkjdAFq+Am4UaRkdIKYnqUibLAuwnUAdrf4tzai7CMoU3r1BQXkC
bS/V3MwhvYeVEUcz+3zkhqJxpnRmniPGC+ygf74vu8DgKcuyLi9Q4Tx9cRNIrOJ7
kd6KVtY7pagnuZv1k8g+nn90Jm0WyNjGrRtc0FcFHPIhDFKfHjJvUl3joy3kFhnj
5a9rvR7YR7yHEUrVYO0BrtvAt0lA7VLQ6bEg2WMv0SeV0/Hf+bSG8ZnUe9aCA0c/
RXzcbGnIa5yhxZx/tyQsfUvFHgSvMrWegCNGofhJ8La7FPPmY9sA7083K7dlklBU
VIdnsfzWt6hQ+EkaGUM5ulzhS14bsi+LJEcCKUscrxkgdcI871o2GFYtO5j6ZkSL
sG2/dKGzYLzsVA61YY4Pv8nw9PoxIhMYMV3isUhqKLEQ+qUOMYTKDyBYiz6j0xjO
CKQTjeNDXdQfxdeBtPcOY9kS4mK1r3tdyJNxmL95Lgl8BnxoRTFenDm8P26JoOec
rVIg/xzShaWMHMa5ISCGC/4ZBdA2xPqA8G/p3sHophHf1b54siNr2/tiuk5bQ7pE
O61S1V4B38T1+UgEvie+E3tCS5NsqVbganAeXEKV5TadmycswyV6uzCJg3kAKvds
3MaLdKh98anYCq9zKwjcTcl8+SS89pMeDRjUf1Ws733pqah1LF4PQJnHeLpSTnGN
08ZJVv0OuMExgIDj6dHpzoY9l6xha5x0K8PluAji33/tKDaHoVRU5zmp4+WtxJT9
GW2Y/0hq01vQvGhAJIqPiO9n+jhDyozOfUuCi3BxEmmwSLCsUJRy6afc90C8FiEp
vycA2CWgBEzbuzFiQu6GLdJ87HJj5JLn3qf1jambdxG9gGLy1dOJeWwtARIZIDwc
+YiN907n4QKNQLJlAuJ/KfMlP2xtJBLcwRVLNxfJ9BkMgZy+T51vnsolQkIO/Y1M
O9PNAZHuZsH1roeVexWBbD6IpZgqMwa0qZUIA/MV8dw/qIC8jYshx2mzi92Ex25q
FGj0nyIJgGJN1Jn5Eib8ZNDFR5hGbe4bc/aIefS2gGKV4YEn8q67xQYr5tKvZ5zA
+RLFFfDB+UPgFb7SQWPSRYTNPVkziKHtBMiKDGsf1jaz+fnfQygkF1KQzJXDt2bN
wJuGpeZnUsoOosU7iOcHg2TCwB5PyCpOgXSux85K5Zh4MyRxh0W1U3pf3R5CbQyC
au/XPhVtv458hshs7Vbjb79pBaVEbPY3MJauNsiyEOpghbO+MSTSk1Tle8pYhCYa
dt9A3G2D2lPc2k8ZDLfFeVPtr5C88uHxDKnDhHTLUALupWrmS0+utLfu7H0ndJvR
5bGANUdy+kw3KA87pO816rj21Noy6PgbzdtznsEVGMZ7kIdUqZF6eY0JeLJNpl/8
dblG9u+MvV+QGLgFIKchq8O6sR5Kv0Cj6NMbI0WZOGKCJCKWLoSz4mt0PpJMvk5l
tYZRg6gcQk2uTbXyz52PbvuWPJtiOlIYw9yNnXUsIlKIDIfgfPsxoZUV/oFgUyvI
9CCw4UsGAILWKgZd8v9fFN4U5EUoefM7ex9SvqANoj72sAIIjCtbcQfI5o741l8E
uegTExVIIhCBZIXdm4O2toS9o0SKYlidedoNrRNNrFZG0ScYZOpCm6+JEbYbL7Co
wuYFWLjzhi7RO99qBmOPFwMH6WcUX8arsbW+K4r0AcZAsPEn6g3vvGvrapCFvkZc
RzJZtM9LLVZX5H1pjKI+Flq7YjzWjoKwLGh5t5GF879u5nUJWw2SrqQciVIup6Hv
N4DXuH3IuSQAynFbA/5rt7eWGpMjdkbEUHNoXdckKQIvYEHKC5PrDppdpRKOhUxD
YmfDr+FzdWjCLW9bEf5m5vdhK1sbE3KnOEU7/N3NFzn8R/91oKpE7RnPJwmEnsjG
VWkX/kYMsoZ3PP1znjow4bngxzTM/PT62IlyWL9GhE62ZdFqObAvwei0Mw2y3tAj
4mmEmJmObon08FYS3uXExduRmBK+CKNbo1iRtBZmsBrFu8cw+IMyZBBBMb+UI+Ro
kAabGNOfJuRvpd52N8RuTf8ADmkSQewmWSk+nFjwtLs88FwbaoZMIazjKbeJajGO
kZ1J3nr6HZS8qkK0QTNzl+yVapTpDfmlhxkojC+D1L0r/xAnlMXmseX8tmjLHL5Z
QDh85ITskdFFJ24DmASIMzxkIWBkGV3xDxwxZlDHxSEJyKljzAi077JCEsfdD33M
d3Pv2+e2hih/otLJM/uj3MzEHfTG4+t6YiziVPQBnapTqK3jzwX17/yNrgMgVzQ9
her4Un+sabm6CuOdcZOQrKSXAsdrawM/Tjk+DIaREUUzWndE7BbVHQdInznUe6mV
wmvBxWst+x2lMkPuXKFNSRH3kBr0W9tSvrFYNxu2zG//frcGf7gfZnDYUuOzFIGA
jqVJqk1OpN4M8HjApNSyRZ5Wo9U8Vla+QCb7nZvdWpZaKaVflbprghrucjjrLdB3
e5mU+NtOybHYKVwrFqrPEJKOTxUrfrVzRUqshbPCMqaz7rvDs9EYGEBp9LjzdWxN
7OcaxxQi6XspowEEHMnKzHU3kwie7NmT2aQUa0FotYsVH64FBqSIqF8jH+kWUGSY
SfzoIQ4dTATx7ASQXDDsZO3JddasdJRM8iCK/24U/eAtZCjZIbW9O58BegPxIYfN
hyrjNF/iU7qLtVgMPfwkDpdeLiH5sKrOVbYLJ+EjtxqZ+4WMoOVhyE6U50CJl+G4
csQPTDaXau6WQuMG3TZF8utI4mOuIWqLDjS99o3I6kUrkqFRO80T4C/uvmn3J/Yr
AkrIFbp9TE3SNEnR1K0yznQgxfQ7HQky+nSM51GCYQ7MJs8bFkkQNqEXTWoXhD5h
f+VyvfS/FIoffrGfvamHw4F8YpPOQt7QKQyIpVm/1+sr+TxBbaAYoXWtfXF66bOA
bCDQ6K3kr8fksHph9iaMre4y+NrDxxldX8RbB+74fScolEPP3+9Xjrf+rZanxNe+
18THZ7O5hFsg3kCY/xEP3++AHuH7TGpY3Dk7yx8JBKqXodeww+u/8KsfWlNzpqG9
Om4hpxESNKPcJeqwe7ZM4gzdIMqQf2UgH9aN66LLQtv+sFyiQ9trkJc3/kKFvUQI
2hdYv+t57v6GPPIkhCmX1n7hj20jGgjRaFhn+96GAnZYBcB1bWtQvO7qNv7yVKAx
UWPFcOx8l7/qiBUz1S8e0GFg/oWW3/RhKU9+GyNjFm021AJaoHlRCSooIcHoEyDa
1w2q298hsQEyiJx4tshqOqin4IHtB9dh6XqwE6zxG4C7BUq6PxT/ze2cPUs0CE/h
f9hAHnt1X7pHsYXNPyuOL5kTLSTfzdmmpfvqLZFSsE1oTBA5TaYbtsLWimBWPljN
NgZaAm+bl6KFEmCEYHt8qmCoB2nH43quNb/JIqcZF0vVMlj5AqOFv/L8nJlnQDhp
QlD8A8j5/B9UCBrcPidl0oZhIWeKiEGFdMx6qw87GcH/uCJdJCZB7+T/wozWd7Wl
Zejnn2Q64CRttiMFPCenpR4zrO6+TPfur4CI8R809EVTF7n0WoX8Io76U/iQCuvr
4z2Dcsk2xEX5ZAM9lBd0ykB5ccilY4whx5dJjLY2moPNyUr4V0aCnb9UGLQPRpVy
eiBPlAYVU7i9jiKY1Y/FuVMD06NoKompxRjYQvRFUSQcSWL03SGQGTxbIP2GLCnq
I4EZ2NfII7q1kCSa0NEnU7DMq4y0JSkvWnZ9nvslSBOIlE/jQD8lMZPhtiXAfpSQ
DrWss4rdHrz/gvj6LDJEL6Q/nZxhW7wAIJbGeZZi35rbdnMrftZKvc2PibnJLPVV
tbeUhBIirvzmoxcazmdIoaUbLeTXcd1iHkRX2e8YRnll4NaMYBYvSnO8h8+r0U4c
MuTQDPknBR9mYtz5e3EccZlRQdhXYDcA9OapZEUPLlLq3KfyssDoqQiFHOFrpWLn
p7duM/DK2t2Ze3JrYEcYvo9CjHt4vZirRoinchfYAOqR1OzzmP7190lcoAzk5HAi
MUQIrycxuTF61C4WWc8Sq2IDJOnZRKbJ4V6/B4SIw5srYU3TsEuvr4dpVC0tSS6W
na8xIzUvG8XCuiS96OdKQF/5ko1SUpXs17dJYmk6d06XJ/mD4wtq0TdRNAlqunTP
CjAJgdnQn5iv32jhoF70kMPpP3F5d5rLjHVWDKqllmkW955Ga1tNqxVcbvqurrLR
tAjyICLPvo2x2p3EDX8hRlPqo7Uf4ApvZwkbA9kl5XfStrH8+V8E2P5EWQ6/u3Ih
9WXtBQwHWhEpiYblmSHFw4oQpWykEqAD9O8or+fHMGlZPnZz7gwuki06CTpHTlMj
CaA1MQ6DgE5gIOi1ZUztUUDF0BvpTqBwYtgEkeqrihOk2R1z39IRTfe4XM5Qamx0
Qdpzryuyd6HCvJ51b9Ig6Zt5mBFJMCBBnZeGuKVSV2Pn/uzyTYxtkB+fMgKvROOZ
gpVsraMEMUsAXCGvElAPtxJqNN9QMPcSk6c3jpP/1M29KGozeG9t7Kp7W2PGtZI3
MIViCTwxvYYVRosv7k7UaePngsiEW9aK7/823gu2/5zi+urk18vQmdSlk0bZfLaS
JBMnMoYU4k+sF91Odc80FHJekKO/OHwivG4ekoS8yumT9DgPYRBQsKKlOgh+OE71
tX59LmrepFdiqCJjLbOCgO5Mgl/CH+q4iMPum9wyr2XdfIx5/56QXPklYtqdDfCR
NK+4dfyNi0ivo17eIOFZOyE5CwvTMcjP5J0LTejUuIelII9PCoIrI3O13OvZdz4T
pw0LuqnrpfYBThSEZLHClQ5xHiQxdv6iZoO23/ZL+di6l+2dC7ojmEZUo7j0R7v4
apUy2TokKADomE5bby9YBuQgBbu2BVp+CWuPjS5RbdJpdXxs2dgi7l7iDnPZvUXT
LfrFcvmvt2KQtHiWtCjZw6tQ8QjbRxXXaTBIhtpkL5JJ2lpjGcTQ7cnBwJ/zP1lY
4iUIPpN62pJZmOnd2FGPoQbBgS8BANvlTXYjU5tch9py4NFN1V83Yt8ioFnxgTCD
EA+qXinK/jJRav4dgJGEB/c/oW8lhIDDQ9wktAFW7AF2RuJ/nfq7YQEjVH2ZhbcO
Bi1I/nBLnVOBGd63MChB1muZJTmf7ZB7DSje8rO4ZzRVpmxB4ZXoY0MjTqF5CJzy
m/Goo6e1+UOF9f8WuRVQ9diEwI+H/EoaIOmIy5OfiSNHDTb6cveG5LCcHCngjV9F
qTN7Fo8nbEm3fZLEpnesfU+avCp9dpG+VMJTkqb0RlEAodBzlTl7h4WxIRltFABJ
DK2LyV49jvALNmpkMOuWziG5GY3nmOq+CgfmATLI2Uv3RJh5B9+Dyb2O49hpo0Mi
Sn86DSdjs1IlRUtk4MtJg+dBqKkdh1+7+lFDywyNdLXAuTxQqlvGgNW5ClSJyPdX
a1DMbmy/xUKZuOVJEqXTNvg6ilmq9gTqRNZSGVS1tHU//fdI8RktVTHyMfvIUzVm
j4HXViClxIcbVqmUCiHRunCzdbYjtSQ2h3Mj6nvULMU4UzJ0ouNbLIQpMyfSXrB9
6ytjiWFyz4A/qBjwJOwHiG4SzxbvkBTqijCF2JIXRuufP4/HO3UH02sjbJV0ap9c
bymFuNiucQUFO2gNRNOs+aKeL4mcTxasfuuh+PNUF3dF3A31qqd9Lq7u8r2+9bnf
QBHzhxGmS0v7m0FTGKpdywXJJsnjjkYiO+lDz/B9VrilzI8aO4DrzfIkwka9te+i
ClgdPvgIE5GvRlDDJGTVIKiEFBa37Iw5mo6xPFX3cYY9JRdXWT0wC9XnaTC7blJr
LQQ7MiayVFe/w9+ssyWAyS89TjsU1uFhA97bUuJPi1AKJW0mM1DRcEuNbKRmkAws
76SogxnZopiKncPfflzTI+V2sZtm09Us2XJg8y3AmeXA+rT8e1JjKf2OoV/auL4m
aZA4yPN+q1A7/vO4/VOkn/rqS+0RIUXuvX8f+DBmuWAe/jTt2nS59xpNoNBTb847
kS7ANz0MhMRRneSlJnc85/hFgwQa36r8yR+EWzHHzDD+sdeGgpJAoxMczdBBW122
pIxdp2XdBs5ok85DooSVgkJ/G6YyDve2abSTp73dzvZNloWFkaMA31trnC17KCQR
7RAFVW3z5x5/lStweuMv0Nf492mQ0wPpdUghGjIpWNIzlHVaSwBzu7B2NCT6EN0L
sgELvW3gcoIRHMyEcgh8PhlrB82AvKpwflHaMqfsI2a1PMyKxn+ngo4oHhicRnTz
e0isHk+CK17W5Xz/isWhwmV5OL+mw4W/C5N7kOAMDb0LxiS9+UrnNfoLvgFAXCBQ
OZamcTGm09Y6Sh2UL1I1kmkUy8JbmKiR93Q1cDprgPkzWRDj2470FcM3qY7w046o
YjYe2/mm/w95ELBqh1w3Kk9+DtWww3InIH3b6h6/Wn/Y+s9Z354jzB/rCTbcM6cn
i7zcpFYHY3GDG1Q+X8DSp/IKe87ywkRGBiF5JuGKqbounI8rrUne/Z6LIsamEl2r
I86HAoGB8soaa1eQxpHQO9Ei3SJc4bPCDN/DwAR7r27wwRdOw7qCewk8UttHqzY+
EVkxSgTwxGvCAXJ8ECH8EMy8GQk9ax0o9F5w3yjLlcZULM9LUSyIY9i1/kmPBW/v
O6Cwr/aslq4ERyYG8rHGUVtLXfv2nvtJVRVDcwdqZj/VZYgIUfZiNnyFIDu2rP61
IWhC15ohCMDC5rM8Oc5lEleZrMdAkQmyNHshnaiUSqQZq4nB27dR/Nm8eG9lEPJS
2E9ayCOvyWSCrPSRg2s02Tcw+4v0fidbePdbiyJdIloFZEIkqcioQSaK2SGa000f
Z131F11RltvDvmnLf5O05kSMz0de/AQxEWatyZStTWeUHTS2N41uurQyZNPzAM+9
0JuHYsKUoNDnoCm+cuCwGBTROJQDX7iqFCsi7K1hPEeOiBPilQH5yaPgDquWOOPS
jnHqAng+Iu0SH7plV7oI8O9bGK0U30sD/qcxbkk0a9higeBsc1wdCgidckV2RSgK
MxIBAI2Ff/2UjadT9ljmF7nq9+qI0UNj3YDTkaAUQ8B1lDf+82Ot5UAqC62xnMPg
wAoyo9MVEsOrpmxdgsUrq/AceXfjb5TANo6KLn5s2LCjjsBfSaJpj4shS1Hf5i3q
Uz6l+NLADP7opJ2IVlRto7hFBO737C/nslDB5ntlFWwnWTDyUmgjKv/mscrLhI/h
pxN96npKenv+JWSwPTq3X0MHWD1DOO4XSc50dB6jhwJCp5jrYT6bQoXs2MvfHZwV
7MK+FcuoPvhmXQ3NYxzsTfTIMn7L0LmlzA36QXFmePv2ZotXh0nNTTWat/bmn0Z1
o87/IqbNRdQxcdCHvkqbMFKjPRVkZiir4ZehlyLHkXbnwRSueCJ1WHjeCYJG5qAR
6rrP4cLtYbyErHy6D3yUHxwZukhQIJwuBP4/K4Esox7jYhiTCXlhfUJCV9pLjcg2
D9P35N0cCgxWKvUBkHTlI9WxNNw52ais/FTsB8Ow+bKq21XVrw1WQ9dvSOkN8aig
SxRxQSX8wbT+Phtomw8auxWOLwTgc6WunMP/j54wJwLeUNF5nApixN2hqQDwQhV4
WGsLVbH2j6pc+LC0VHPILMqEokk4TuL+9TuAyVbDqxS4p3wDe6ilxujMFUAtbdE4
7uBJ4+9OkQHL7+ciIQYiIP1BzNoSRZecf4EY22fpChBxrset/2MinoiJW5Rj9pQF
qLKJa1pbXJMXLLPduxuLxyYxCtEDjWD9mPWx0cBa9ED//qqW9I9NBi3rWmdrBkE3
QXlci/UQ4uPytQiMORCdeFrocVWjBGilo2NW8CmggXiXHA/Dt7n+MNTK/w7XHZPU
oUMsQETj5vN2elEx8ti6wELurx2BtDBYL3IHfBI0jEtvR8SRgS5XMl/7upTIU/9Y
3CPR5gzRfwSehxHiFmAoRxoBl8QYL6NjL1eTyx2VG2TXb4riTkwf/EPRVCvUkAj1
9zBL5PoQnWZoQMMr4C2EIClgHeBIx4i3VVLVr64yy/z772YaWOFnjrdl4KxKAkR8
gVvdPTINz3v1oXJSLXqTKA1b1F4pUnpExFfjRjIy6CTTkkcox+Dbqg5amG6iTs12
Woe/QW4hDkC4RpulXZgDSqZtXgc3JQZQBLVtv96HxaPufJdalLYNJfFNfnkoYspE
uKy5rFM+0cpqVvMARxUi0+qUftxqR+SpJY0Pq9MGMmZxiImT/gCqSTK4XOfy1kff
KCsAyIrj6Au2YqyRC/Tcvg2PwijpDXL+3PVuJKaRFTTLlYbLo+9cW1EbjX0HIB9u
7xop6mB1GFxjt//8mX+jV4EcwjmDSlCqg3pE1i3909k0KwarRh+Gck/OsFTF9pNU
bjBC0l91bZWrUAW9qKy/kJAZqjVMXUkFeWQR4NLGSz9x3cveV3qvQUslBc6S5MEE
2SNMYf/o+zxarSio7FzgLSwqlll682oXh80SCHTsBlD5zlTvVGwpmuQ9DH5d5wJx
qehbDL4HQhH+ji7ZpogC+EVTnfXQHCXkSe9I2oYLSCXEdlOJalGSsnyRiVHbln12
sf5w3MvjhV5CsW6BnFU36/O1p2wzjbGAD8EKYzYH9fohmOFXPhZHkzzKoC7bm39b
hh1k5zf2eRSaU6gZ1snSIqgHPLlZ68F3DkiiHmydpsghYYrbSDU5PU5XGxN3as6Q
phZVnWvLxShXeCrj/cyGq7AF2qQF2EaNOBj3YCGpnVuIl//r/OVG5WbZpw8NkXhL
R546CVl8AO2bstdMeptC+m2xuVinGrsQB1Acof1+a9+4i3BxqSrXs7wEeBQU0b1y
TYp+eHVokma0tD7da0/Xg08VJMJuasp0fWLXsYUQGKj51mSqv2xvN4fggPR4q1Fs
+zn7JtGlwyZEiodfbBiQeDDx+bCjVo2sknHdEDvQBvYQLOary7Sdb7VSp717nShn
i5VydMc1y4YpXL+ZD0Vr9k+6UOZCXFTfcSNWSOLSu6nwrDHFh53nOm4Lnhx1KuRG
WUcul75zo45KQIeJ65ZJJnhPQQO2ZKX2QYcQl0VLUFwpsmGoS44mAh90NbVKv4vj
ZQcJQ9ssrJr9hHuwslquPprUsaFnOu2C/oQdiQrm1zkBszXdMsfPIFw+EV+SKk9v
HfLtsmb/zH0nUNH7SmTucqtOfXI0uc5UT4oKVOi7LG5PmOfVAL0TL0FnTddPbCzc
3wqqtYTz/5Q31h7iuRTM39qTB7qet4j3975KDtT7rZzWJ3IIQq5AiuMEOUU7cxCZ
pC/pfK4g+krr5cVKtvDzyc/4y/IPoe67lWr7U5H8VYaQYFqp3cSMBYUgcUCymxrr
48cgSHhZ0PxgQHLy3aVPwL3zaAb8OtNNcBUj9o5rptdAgIg5h5/0DzYzZ9Ndqud7
lxfcUKnul9sQ01nCrNp0B6THflScoC1JvPapHBWVj48l5IFu+vUl2WjGRTR/9Ozg
dFWPmzHP67LUnVb2v6hxM/d0ei7hBoTFwdOAZdg5HG1pmmIZ311I90ck7vVT66V9
ASPCLPINGhQ4OHIqVmSnBxPiWk8SmImip3GfZRD5rg25DKTXl6EvBn6arx28EkDc
b9TWjiYLH90jmNmmUMvPCiw8MQgpVvwEaYlyXJILbfq8mMuEn7pXxBqvDGhqgFdG
vnVx4Pvhp57veeVtSyo0qyU8zeCubRwYoIjFpNRWRTqgl7tfwn80cAVhpDR72ZOQ
OZQ16OxCsrq+pJPMpctuhYV7szbl+ejvy4YdoqFTXQZrb5VykoxMwFqSr42zAVOQ
yJKPkpPbagKZlEr9BZKjYfrwo3mAJYpa/wEkkVF3kXYogTr0k3IRyjnuuFxR/6ns
8AbbzN23UI/Rm9pskMk1U0kN/ncxbjTc+R8+fi8GTGqys0mcGgTd782vUFOzzvtT
LlvviZz1ykRY41zQYrbOF2mweUXFgAuNTxxSz70nX5vNIT2U7LUCTmq95iOBNr1C
51g3/dbe0lm1jy1xF6pIAiDHo856VTrwFW/fbvldDZF2Mf3dqBuEdbE232T3ejfb
JUcyVNkjN0jR2uUkQrLXdKaXHcQKGGB5uUqv21HmV2xew9O3TkX7GHeM2LRjw6XW
kzsbVbuMtgBK3N4nHwV2SjCO5tAKI9byGduW6WKAq0PXM06aOSyyPa5JeJ83wyS0
VoBIU8NYwvvDjjU6CrBTH4+Ajj5YsKq5FGKTXC7NWds/y0Q3Fsv3eu6W4PckRqM8
ZNJ0g9Hg/tMUE3uqXNpD578oqYXxAnINZ7YUsZoZbC5UbcvLfHfCaiWYs8kJiWGA
10AfoO0bg5z4JHIPkKBgpH1WEkQSBdKrUU/u4gMS9UlMhUr2zCrNj+lqhjFOUSYE
+JhehIf0xLyDVSngn9OyhfuOQwdpW8kkZ3b/D7fmQEPn5Qv5CUgfnrBax83VNayC
4OyeQYpOF4Zwwt7kuYPvTW1YHvH6VibGYQi6rHobt6h+SHpb5yHDLEVIJUP8xYxp
N8DbCFuR5IdUwJ5YmHgEntFVINs9xVxzQUZIUbSvhM7EPVvDgSJvlHHS+c5o/HIW
xX1sFFCYw4zIho2pRfDrGK2ryA/ZdXpyQFlAvSmwo0hfrKMUFiQKU+3d0YUF6c4A
GrbuM74RW3vTKWvjEbM1VTrufa3bRxV2DQCYbaVgKZ2hFnwEGVZOtk+dBMBQX768
s89jR7LPfqcLTUSOA5GDoMP78fEOV2Yp8tIexmnFVwSzy+48g9zlcu5bIk+FMwD4
GfkW9I1k5F5cDmnEjKrGcaw9bok6fSkQUkzytPUTJEPvOi9APDeSqDyCU6ENXs8J
2tQeZk5vuVpiPk/09AlCnt3POwPAdtqXjxTJqmAMK8l5fPjUyBXnvkXssbXp4D6u
obv9eggOy36lxNlrUsCs1Mf6MX+WfbHOGKeYKKSW1yJyMLTH8fNU32dEd4/aHvm8
JF72Hvx8FxElbzIobQ82/paOe7Oc3IHN0ygyrx/WToMtO/DBam+L/07g3vTjDDjq
fveJpca4Ju0o9G/Jw/81x/Q+GVlRAfYx0h9Qux5y/h23F5NMudKN+aK9J/lD6wpn
kojfcc63xEY6GB+bs3bA4T/qj1ruTOmHG9B6GWWgcH30gS5Dz5oPnUkpP932w9W1
AXAb4upRKbE5LTo4UZvDTTj4ePJrpdzTDHVgfFUiPJYIJWlnYAR4BhMWL6mUb1dF
9l772DHlAHtHIevhOZ+ito98Mmfocl9vK7bdoySPXkiVZsAEd+/sgU1HdKceNGlj
Mso8/dTsrgHDzxXyuzKCoXymYrDjFv2ECoM3e5FECF1LyGqhhho4/ITA2qrFJaM0
qnq7ogzMu3X9YZrwvv3V55nq6gvnntmjw5qTuz20lKXrg2Vc0wnWnfa4O8YNEjvA
KEb2rky0nRarmEaPnnZKA2dqRAvrhJUm2yHpJQSkhQH6qhvCuSaUi4zM3PCAqd8c
8/kDXrF3+tqOzSq4w5PAzja1SijBh0OOqKksxyj5RU7JwJG9QDeVkh4jV741u2L+
HKXLZYK2ljEBOhtKt/nq7eA9ufxPtH/1Xury8jl75OwydhVoLtav8FHz1Za56ilR
kYoy0+LyxWkd83LZ0OWmN6weoL/xxKbGYoo+Wm0Cfq1nhpK4nSp7uToJXTswYub8
H2eU8cJtt4GreeDABQpuMAVGLhMEL6rBNdCCTQii9IERGh57Qh+KTz+BRnHDYood
NYbsu/vu7knaIovlkUQEukSIPCQpJjZmPBPJeYdR0K1VDqWxM5UzGjv6ouBJTRYj
BxAXUf7pyxPg/gfNGkRMevqhL2ggOj0I8JM827CX0emltvxkNMxTvYUzd77R7x18
qLqlwcsI0eJIXspcyaEDOoTNgqMBr0h2Y795eg6ggMWBnZAEjBGG62dwCAOEugHu
xO9mdvJbfLjI4Ck+g3bZJzru09wS/ndfcb9fAanPINnESO2yzw4RqRGdYOrt6Lyg
wZDLC3DIfNi1uGNFq2C7vCEWz5Hry8khIN+IeZsnu1H+vbvfvRwk12SCp6eOB1Rr
54j7AQZDYSGZprpJLRJANl51AR+WcD551DPSTqZDJFWXquTNOcd1L5/6V8UD0CZi
px9+penujaCmzSZxK83MBPyEFQUqxFFD3ThUykT/TP3EUppZW9NMEBp089zGCEsF
DhCX+ejAZddQjGMHu+rvsHhyruY7TfjORo/cWk9+tU5UJxZublBOjuOVtmVl8vW8
+pjdGueKxLQlYR45JYCyQNfqb14mz4QnUzUMceS77sReySqtCIT6TYQs23oWDTjS
By7iKRaVjeBDHYDhu+5pAscrDUlkLPKVX9S5CCWfbN5hWn6b0+BGjmTIocYvb4Yu
jBXboj3wa47LHCP1/oS08i8JLZfeVn+Gmg7dbgSyxvAhrgu5DzTQLDtgR8WhzReC
9llHvKC8EXZ4BJ2QSimSAK6z64v4GEnck5/VuaITTEMJBIBIq5NvColA3j4i44hq
IrSxNa7izlsmxbvhDvdOGEC0eL2MFDon/oS9yft0rs2ws5rbOWale+u/dF0zrcFy
AbXywJCO/qSLKbftbTlUMtIJAnjRLyQtFK98PWdEyqy9bBZkiBmskT1erKd8EeIH
1FU5vnCWB07Q0x70P703hu/W2/14eQonw2xZDlLpGKDLPInE+zK/NUAgmNRvkH9k
hAjfpkoKaDFqqSlvSdewXnjPNKKzelJObFfC3v79mDk6qq9cbZDvOWi5QlkWWDg3
MwyxANdH5Bp1QMPvmtWqqzX5S7eNLJXxxt0AG6c/43ZY7mTHrV66sA9pBjYj3acI
5vdolp/4eGfluUkBHE5g90rPzCSKmEGzbzm0sECULe0No2cz4wfyFDGyITepiJuJ
pxJ0s0tklLLf1WEHDD0tsl4VJxzh00tQM/o6iefZEtr9rw2TzD1GxEHwrLX81AQa
Kq7Ic8n1siC/JMJ3HFr3TkPpAyeDfsW4WmqoUZM3sJkWfOEx2CaVwi2MKY/djTrR
BGpTeX0HrCxysGFko+94c1ZvR97Qlk5GKqElFiISuD3q9NMSkkYCaeALqy5cMFpM
GrAMTKfT6CoL1ob7hUDkPFLMrNEOvKJuBAJ112sMa+lwHZw97AOiazAaLokSlWjO
QX1LnDyUydWK5JASyAxTA4acIUuS5wcYuYnmvZPEV3iJ0NZYHuATKp1yOVfouPqQ
5z82Gd7uXvxzfr/CUsgMhwBl3NQ2bNwlLCpKwt1IQQW6rhM6Qi601/AEOcAi0voe
+AB1HajyQDUoHsp3Z64uDmSA/wTzqXsfpprSbmVHJjdbboKl9rXp8HDLqfRiyNxF
E+EAgmf2FFTljY7nu2hvEXKyemngRqZXrF5YILmEhKCGomiMkeJO3ft7k55pilw6
dOKzS3XOd7pJBnAhcUPOaN+1QkQ6VJucvR5RZpN4T0nUrXI7MEtlWwkkkHqLbgwB
HdcP3GOX1sZMdw0pF/TUMy/U5TyFWQor6Mk3KNlFtsFy2bm1vovKrJEkkSFyvVcY
azU2VY0z4+6dU8lQQBIltSBjvsv/ISPrSzvkQ6EHvMprnOS9R1ukqqzIV4FH71Ge
qmcn4SMwO0iYUFOwYH0O+bf6iqGCRy7OFeIzaOttTbUmQEsXZAizjRttOvW0BOlD
9XBTst6Mkrvyf6ftEE5V3u4HRWkQGXHfrhmpCJOLS4SF61XFuHThoJHjUuuwsmHe
A8FGGHjumCHICeUJWTwN2y8bUlZ3jZDPLuTkdk7pIlAJYawkHwD47WYVeJdrKLFF
auWX4d/zMbnDI6kC8JmhQI0v6ZIUh8otAO9Qwdwjf27sUB9mDmTDQF9IlKKSKz9Z
/ecwoCrXc7QsYCrF66I7sfq1sCR91AYfTCuEgAT3bxsv0bVhTYGKv0o928iJV+J+
SYvtVzcod4VDqHETSfIzDIzkSJF38mCR/x9s/MdG5DEZNdoiGml5JU69agyhVpVu
Xj/iruStnauBGS52lIVddScnJMyz0PRYc++jT0qlxOalUyXXGM5jpcZFQJeCzMBk
KSoMaUfmdcT1x2ByrFUcko0HHbyGb/+wrDozSooDdxpwafvX6aQOZe3wngrv1a9C
aIgvvZ4npIGvftLdoIMbx5d7I5sSqN4EEeu5BpG1jqW4z7G3gMLXGjial5iTUku3
NcbtrKM7GUlx6QmcjzCm0uet3ukKZ1Mj5kY7QwI5EFCG/219eV1l2i0DdJsoTLwp
vfyGIWWB/y85dSTQ/J+CkuZSudST+Q/J7WshAsO43zm1kErOrf7GST0LXc37uEtD
/Ps3Z7Omukl4qnuMW8NtVSxxNWGQlxordSjOzYaTn0PV7+O5eB7WHiejT0O6N3B+
c2qWsS3XCRo/c6q5WmasFrti/R2zovf4/8dyb+XiaONHlF7CruW2TwGjVt5j/gbk
g8WNV14QRwQjCZi+xHXCtvOlyKhwOeY833tE2yWk/PeTb8Bc2ruvil1ODK2A+yd3
qAVRqfVBwD6Wc6xzWtvp7b3fDD5CFNxmodXi9zmTaPArBHWci1gARm5iMgWSX1af
c1Crjk/ACpC5msWP8+bVwEyu5YYwtqrTY4VA0zFTYT/DspZLh/r63FNT1o4swv0i
luxXehiFz8bEBkAxuLErmbHa/CfBX07JIaaFNnaLyhh22YLqKm6gHhSQt8l2OYe2
YT4JzQ29VgegB2mJbHwuGUvpfqRGf24Ted9cN0vHFnfx/sX9ZJhDSKnaWIvbHbLY
EdXTidSOdk2rXASeqo/XpxKp/9vGo59OXSczTwWD+5FN7yik86P1H7IaoYoegS4r
wvSIECWW+4RC9d0bpa9Y9QgFLl5q1vJA+ZzzIX0mNqwWkxti29kulUdoJ6yQ80cq
lBJpsvNTNrUPA14kdsi5ESpJfCPq0VZrLhp/S477SpVXdK/HLRFxn0aMCgyPjCbj
sGmG+3Hydu9XQ6gwpgTeOZqb9LrqBAC4HACGVXydZjy2IxQ36wpFDxKitTm8o97d
SPSdmOKIGANHZW05YLVIb8c3JEXdLei8ou3ZFsaOIRuMitnT/hGet049A5GDCLl8
4CUfW7Rf2Jrn8kbX8nMhImxlVPfNm5jZK+MfTvqiKEQZPNvnpuvOgQ5m65QXHaY9
lRuRgTyTjT2TiUDN+IjHj74ic6WL1azRumVyLjK+Kk9vvyjDJzptM++a/5YcxmIW
3NUS+CulJaQfBms/aKEbeha1/gBfViqNdPr0dzmo/X+0EhjkAnRwpQNqouBA5QnR
acRKsoS1o7CTUSlmcBn+zBuQAj7ABqruHnBJjHNC9JKnC+ixioz42wlILfPv7e4H
dEI14ssbR/hW+qIGjvqQAOHmNL8X1XMfR46aLkcRuzWX3tFJ/EFQKe4Y7tU7K6Lr
wKStiiV/+GMPgtW3Eozb3C3IQODI+kATdEGC6DBAOO4u7mUFxsNzqkLn2HDpVpHY
pd4GOpvKJaa0a7Olf4m7MVZ3bCZsKlMIJj6M93bhesQcgZWvPuajVT3Pszv4Mneb
8pjOtaY+TjKY0SVb0F3BW2jhG4CkB2+4dI2ltBRlfwL3kl5KkQaVcCX8vTqTuS8q
++DFV84vaVH0xjDgyykjSbdP1/QEKt3ig/p0PwRelkyxZvTUSXCqx6j8rbB0iPaO
w4u5byYR7LMLZNvhuiSh93SUvwATqTIxGm1ncdQDxzPawMI0k2hIkDgqOhw5GvWS
lgBDQaGLuOfq4VbNM8uiw3IfMTHGaEBca5ps06TY+F++EjfbV8lifNeGHhx+Gtk+
fgo3WP2gQ5fThzCHQka1Ym5w8HnThZR3NOYkW8FgJ3vUk88BW0/4Kjz35hptZgZl
RjEdNRbfcj1Gsw1eDuZB7oft64x04WlmOOmVMdOFZl7aVCGd7slWhZqjk3IIULGZ
zr3yXxyfjgUU+hDr82AP4N4QtMjEynAPUfmlSYas2fkpk3Y0XvSHKehl7Ekt3w9s
zFJZN/Plg2leX/GFo713aUqd6qTgPQLdSz+MGsGfPDbdlfStdDP6s0kXquXqsza6
ZQySmtqQO7PQh0PAzjLBP4bQ6G9bGTJelR6weEyefEX3LM6c8vsR399MhlCTWups
sAjQEP4BPvuTKOd/SIqkH3BtiRlt68HZ11sZQt3gobSlyd703nKGbl8HCD//ov0P
q49A/6lS9IkPj+u9CdyzczR0J9nE8qgvN+cdq9adeZr1yxI8Ku2aMayM/QAlC2pN
2smr9dDvgStjt/whL/7YXEKuYFFHlG1uSkeTrvenvAVWfB1xgwgi7t5Lb3o+t3Ay
GVDmda+iwVYLD7ad6oPUsDOUv/B2ck6fOPM4Ok4ZE6wzK6u0+zd3XSLIzq8Cxrr3
zrH5S7aRXq1lFXNoq0KhVanLfMGVwLMVUtMOccgc7nE0Qk6ez+IAtR2KpHYePXQH
rkFFnBqGyMRDbVqCmA7VCbcITiV0imoUnWPw+v3Bk9s5oSaxTeeEvNT0OlYhV5zc
w4V2m+IibsJL0vI3h5H5zsbqsj5YqT/XogGvIlDQR1I7fy65U7jMQKvt4sUVt7nn
QimH/sTC+uHAVs/I3nycrA5uCSZJRyU9qczn5FBHLHQFBDxCWNFGs9JplE6C9as/
fJI1Uk45yHlmTH/Fg6TS4Iav1eTmCYqPrO7VTJOdv9cM5H90HQXQ3DBE9TtevtGy
D4ej+fzuDmY7eV0OwEw1o/zv1P6NmgkdTYVPvwCp9FpeL/8VBe9QJd5UwRuZMyzi
AzVdof9IVNQBqT6mRiRkgTUzx5ACMepowck8r1xCmwC/+yHO/cX+hcwD7DoQkzuw
12A1oe2ICh+eL1De6SHVSp0DIhaCAkf1Pwg7k9TUrYmsY83S4o59VEoHrjhEsP2l
ZJboT2NUePJpxJuBVQj3FVnEINhc3al4YtsypBy9Qj3uErtazJIh3YoP5oQuIUZO
rjd6Bohv+PCwezM0dK3OhWgDPWYg3e4/VuSjyaf2bUn9ZtUArM+c13lyqoie+J3g
kswJy8Q7dhATfVP2G9x0O5G1rnXBx2uaT5j93clOjKFztPlRqBiHdlEBBJ5M7eEm
ACIm+K2LKdyipyGKXwkrBARPjHesp9Pq+6/OnjU9xc1OZxxwxWqKLAQtvbGCeI2X
nIsUgP1pxLBL9rivtgVBMN7VBCCXNZBxQ/D4kI7nh76e6T1vmSQ8TxE6qRZluRWy
pDGEZwuIFWfetgDNkvEeJV8KjQsvc0779ogtIFCNfVn2ZOy7pXwVD9GtSm/gEntB
ALOmmyl9ZUqQCAWxSn+VNg5ASWQoX2jIqjWEAn/TSq8sJZzJeRR6ztamt74GRYiA
Za7rs4vOJgKuatmoBWnsII90Clgu8u0x5VCO4f6jN2dG+I/1q0xUeba2MKEIsDCX
si6MTVX20aKMFhG4hxD56ZHnkuEcd0gC0N5zSVH++xgD9V+CZeaDIkdaecG0VB9M
/fOG6uUs45s0V20s3xNjsSFMolJ9IOC2ubKd16ngPu5Cu+kBUJJRavgR++RrZFf6
//YNvDBfrd8aljcOof6vdksjFSBkGtR5SszBCbedkPPeLcc+W1RIvCJs8BhE66e2
g+JPj06YuNd1L243oqgvtHCtZrIAzhbtk43YBs8/300i9csN5an5rfudNDVI+gFm
626Mv5BOHGtSvKFCNECGmn8bWSgGBCJeZZP2JeFj5XeT0B6LAncpQMVhegtFSaUA
pQpRbQ9I6YYWImgwp/bkC7grZ/7o6tPALacuVdK+UhaCUaWKgPpARYOtMyYY4fE6
Xw+CtvQN2c/nwY7vsAA5nwhYdgmU4ZGOOe6bMxraeJdg++xnVEZZrr3mmMq0K4yl
FGsgcTIko5/0JcEWMrbcx6/HBa5VnxUMpECnVbBGW7rOtKSkhD2vAxOR9NK5X7Q6
w1dOHr9KeY9VGSp8PuzdcHonQ0Q2kjfJZBKA7gl7Qd9Hi075Why3m0xmKxG7kDkI
kiFsW7Eda1ZVc6KjD8mPJMfGzV38cMXFA7c+iBghX9ssqp26VgK/K8Z5dMZDQG5g
sY2X4QoPYVWW+zQ4mDelX8IZolkdYlObp4wFHhAE/qtsTGNL4CiLa+Efp9gJXhdq
qBvh+JPJ5ujpqpFjWmWLD7aWRI24edVSO6ea5y2xbP3phwHZjNlFRAlzY/kkE9ie
CJ3doyScse7spKOpeSEbJUDqMp3rD8poEzQYs9MZ0ovN9I4xuIARSQN1qIDq02vT
r5YHtOMzLpN18q7UTs1/SIunPztmYNZQu4matGQcHpbxXodvkXwxmRdejSucLJgI
sqGqAIp0UkQLIXNBSW4NH/kqrFUzFcBYiscYJgf9lOtJol5GwB7l0K+5ogf8EoX0
AkQMqXYT5LFvVkj2tvtDCHKKyhjFUb5hAg0+kcWZylDCPQ4hEHwosH7gIKnye/Nb
uJ8wuglRLpo4dnXkpjzhLcbtI3wdI2jfIFBNGG/7r+Y8I5CyEEZwkeB/hcphgwc8
KNWJEv2CSJA2jiVyW4C/vwIOX68oT98x4tJokzDhiSmI9E41BiZYYSwWW1sPyDNI
AXbxHxD9b2Dagn/V8gtnFfAidthPWMVamGaB0H5tIEVbeGOXZsPccWC7my7HT/ZD
nJOl+PYgI70QUEfC7CEsaAroFw+jKTsjfQuCb/zCF6SL/H3tNxaH/asHlMpgmfky
RBtTTAZELJtw4MRj9AuNBVjTktBXqFAF0FlIMrreYd7O7QbtunhUGHrU6GfDPEz0
gbI2eaBneijxAHcY9lCovcy7Gbk1ZeAvmypElhJFqjU0yJJIdOYqhswEN+dM8wsz
pC5wMs2rMbSo0v52h54jVY8Lcz8dN5EE/2npoRBEGiFhy+HvSfHJL9TTFT0GFsw8
4l9kHN5kGDwFjmCsofWh4qOHjrcwHc96ImqydtTCD+sWkgcZJdfaJKXmYt1Q6nZ3
OXdaGuAWdRqeHrUrJ3OuVGdn8G4/nzZbRPFKb9MMzfHV4ediDlnc40rj6xjyx1Wr
VtC5BMfkgXzalivYo0Q3487nuenyqJZtIVPm/TckJHo7/q9ve1XejYA7vq98rEN6
xXIws0GRntZRXPIdpHL75IqSIF2Z1oAoxc2OOyNR2NA4eRArlmolM9E8G3G3fo7h
jlF6ibucWsjD+XKjF7Yy6lT1bnaTTFQMcI+NXwle8A85TwOm1zYkxvosyNxCaX86
xZMA9YizbDbd/KNW29+VsEoJ6/Kkk0PKpNtDXxdIV9SeWy1AthPwa5OAh7V3FE8B
MaZWb4TMMb7BYK+zaF49Wir9q2gs2XxEvxfBt2oBBDaaKLIrUHQ04WjbZ4etWDlW
rklob+BntlKPeilEnH1jzHo3dse69SPfQOecXDYoNjBBwCL56Oq6iYHWvshc9Tbl
A3mGg/jLzRlCC/6xTMiVt4Qpd1556rEyVUEKz4STcCIkDJLInrssNMc7PR41cRn8
rBfUB1rdStD735KJ7JFXDyHOaLmEz95khYnwEj5tZTaJFKT1w9VObG2V8CmcfOWD
6xeOIGSAQwuQVzAvu102fodhBVtMfj8GdWNQNPV4HcvmXmva6U26RAqBw7uKhjdU
FmmSsDWU0wBC7Jensk5cm2Gqz+pb/FRBSVAkAnBpwom3GBlMX32k3ScP/rMs2gT6
z+ibVuZseNlesJitFwOVr0juaXgldDIkLUl3T/rRs4UXdv7kFiiWfJ41lctvL46a
6sOmajJcL5x16FV7GCbrigDcXU9aj2oioaozbFyMO/Vfq4CnbTUlC/S8HgSmfa5i
WU6ojf+KJs3k71M/f3pBVc/FnLZI2psvrQGMmuUZ++3fZUVreqtov3sZKw0vFdgH
BiDVWp6QD5CfP1kzMGQ3Dc80qJHC2UZ1KC7mRwhUBpBP50MZXO22FpyCm4pSQckU
PP2lGqk5ZYbxvl20VX/5so3Mi2dOAcvYzPhRyRMGr4mA9XpR+TWekBjrX9l0w08Q
cIDE7zqSnrJoZC4NdXfmxBXxt46VE0yoKPLp9fSeqmcLUvZG6wEA4O94QjdLw6E/
YZCKtrSpDfn8OzhWGD6E756cojS6HQF0upDXFJs4zXne+TSya/03q3TKz8VRk9YZ
3z6pR6RseRsdqU4Mt3EqRcc3Vp/zZmvN45qSSaxZxbwPI4eZlxktlqw7Cz4AgDjt
c4H2npZL0X5Ed36igW/8FgUVUhSssI4HHyKg+RerOf6xMj+l4uxbRIv1Tw0vBWrw
4r/kIs7dvYGbl+ulrVo5R5JWS5ENi7rwFuuXCLaIPWG6jNIggUo9XGiaET/L78r8
bwfA5Yt9Ptw578OOSnsNddLL718WXz4hUS3yTYpktXCSZ5VH9g3T4y+XkG8BOoy/
EiUlYTLfqV74BnjV0pVgmePiIsR9t0P/AkfOp3hzIrvmJZovjyqHTqgxh3orAqR7
BlveV0/EKeCyDCHi1LrgI8rtorzR+P+jRL5uwV096iCqEqXkBVC2oaKweG+YZJHl
QHp5Zsib+IYSSprIRhL3svBZ0p43fe+A4pepGfj68rHuLstCbxb9SjEai0F632Fc
wwnB98KKYIAk8yPXtEL5c1ET6pbSJ35P0WXU2Ub0+sfllPepjoW8LgIeIlj2ilKb
ACG/QyFEi349ccMNsQ+ZgLzo8xIWyXl8c2yWXg7HMn25m8xrwtorpfJR4E82osLX
CVCjQyKvGWw2DSRf89vkz/OzWZDEU3kyPuEjlkumhKdW9SQIKKnzfFeAsmeVcUdU
9LH6cpT0ZcJEoSL2BM6UBV3oOL+qCVfmjuMdRg4aHElxpaUz7kpVuJbLC/lUCp0C
w+yOEViS84ged0G605mQIlr73XEU/wJ6j3IDVJR2stkfilIkkhrCr/1rEIUMFO+b
egns9dGjmeth0FBvXMgX2ah6mmkcjHr2c7EtEql9el8ScxANUB/3RP9v5LU446Ox
NHaS59BE2uCUAzfbM7eF1lu0hrn+Pe2RRyHVgWYj81N7lKrnNQcWUGlV/Yh8frCw
twsnC+azu+gZs29fvNWnWH7lW8BuItkoQ1cPIIMH0mdMY8FZM+IxOTjdszaMMO8K
T7hMmtka+/2+ljXZ+w6HGM5xtISyDw5FYDLI58Z4D0jci1gaqY7jkXR9/DuNaaT3
+PMgU8IO4Zmp7O4/kbvfZlCyRo/CUOEzmIY6QGy+pWFgYCTpkk4UzdFL4wEX6OEy
xwMOXvlXYEVSo715I5dllA9uBUkVvBGNrUG/ont0FLHBDY8n9jPlZ55xOzmYInmK
yEM1aoEdd3/WxN7WMmT4pKK5UXde8vIxRVV5ZaxHSgsbfssVhae6Rnp+j3NYZvJQ
Nrt0CFmPRzU47japGlZAAFblUk417THYogek9s5OR2jXeutGm7B1tsLJceMPmakV
trW43KbTcIszlRX9hmPtnNQAPJPQVpu9aGkyu2QnCxd1dzCD4V+KSZX7WDLMDzZi
p6zy7zlXM8be0udpAMeLV7jrOWMHIU0wJ1SXk6NOMYeAwh8z5rRR0qZ6bPUS6UOt
UyG+bSK8H00eTxeSDUPIdYQUqapSOoHDaV6wwLdEu+yomgFZU/nHXDp8aaQME+De
gZGNpFKJvEzNCN9RqQ5y5vW5hCBPWFSMcLrmp7QkGpzRZ6lGJp58ETW1MCSq4vWw
mT0x6O3SOI+VoYKKCLdlSnTEuRF4oqLcLS+OG99RCLcKlvp+kF6ENXL6p4xQHIld
dKvNp62eCIry+w3PmgayK/rYH/L7ixktE8tY0rrmyAzCtQDm3UekqxULMNthv/8g
v64F8HHtUJRErrtJ9d5CYqjpk+W0dvaK5ggtQzoWjbAevEYpAGiNceWG9IgDcqHR
KtOcZH6XXC/MDnOT9QaZc3dVKWtly09boaKBWJy2iImJr0Mit2A2H+hWoy+exUQJ
JsMgScxMCD8X6kqSqi5t/Sxj6cJEHDouMBEBkVapW6DvfkX2ric0FC0mzF4hvHQm
q41jbSibpOBM5JntavFN/neGp/vQ+ln0e4BWOdZ8CquX+5oKBOGkF5SmIe/5JB/Y
Ja8ukDJcgbtbjw2uWtWlnKZzK6t/Y7y6Z1eHEBxLSbUL4ih9xGdd+aoFCO+NZ5Kl
0PgqEHXuJTenZ0URx2gQkoGehkjkrjKQnY8Q8KyPXVZDjwXZC8Qr4Zdt7jp4BpI5
4/R2m6Vny3qmeqhJeb2fIRUyNSYrSLqknkJCbQJBM9P5XNOpDvfceq+9oPui2TyB
LzTjkkoktp48aU7BykWdHwtFPy28/EbwbiThrZYOB6TWjAvPZov4UqNUo0w7yUeN
M2d0z9XuMOfLNofLutEDwhCk3MY11ZOJ58DOWFL3516OLLok9yE5yzPYy3tHXA1Y
w412eAf4IV4vkJyeJUtZqwvQkhYzCOCv10ogbO8MsvhG8Ck3ktYy7R2rCxKJEruD
k2Jr+28d5KzmO9zleMY8jVyQYRYj5ehfbfJc7CcVe4jb8ZfuBydc/lJBSr1llTIp
4JRTZEMzQ5zJXp9URheVABz59QECzdL3qazg8nnnBIGmKBygtwYlgqXjVBw6rN9J
qzoYVcBdHnTdlwC5QR9ExMvgMMC5JbXWWyCD6kVn/GKi9T1oEsIVY8+XcB+E43i8
eb3SJYCPpj1dxQgzVJpDgjXgEzYRw+BIO25iFgZZBZi2Z/r0nMhCXY9raJwq5E0M
houGXS+Aa+FI9C0Vla23VI87da0TF14jwGfjH5aM9VhJrp0Qm1AaOUzBVwc8lJRW
XO4BKfZuxAxOnt7PVDYgUeLnubfMnJEyHwEnRmC6JvylRezn4vEO086oes7tkhWV
bJglyd+m1Nx/xovA3Rf7UOfs2ZhHakrH4L7AoQHiqsZKF3W3QJE4MJXTWK1gxKNS
8CPoZyEQHnFS1x4j1HFERf01F4ABbqmCcZ3qjpI9gA4KFISAs3bzwczDv9qou43y
0Ukbo2Xed+T842SMirjMGv1yoOh1vk62HfEphTdstHg1de1XR1jVveJUvLSwmNsf
P4AZe/QerEaNYzaVwMYj3T7SEhfz7qqQxGOw9nopOOYwn5s3SqqS/wQsHh+LccrV
xh4/QaoMS4wrF/u07fFA3gqzFtHlFuWEUPYZZGS4qLUrR2TKnNpmX5GJM1KAU7e9
DzRlwuSzenU/MXi23y1dSMt/jhhkhxLAkyS4OX0kDPYM5DiegGl59Tp8OXsIwDbE
yewSO8bYd5z60QWkxPSY1oQv+LTePdUyloewsNezgm4nCepINqsvv18NgMFgjhAX
rfaMZJIhzRhj4SsMplsTf52oHYFPHU3RFLA8KmRy8n1jsptg3rHr2cSMj39afh2i
90v/+PxyCbQAZXB4Zy8D5tm3m1qsZ4gCPcFK8CPpq9F3zzLvExPTF+7kej274hSF
Zr7Q2V5V5/iJodCzjGgtArPbtiRlWim0WGWGhB0A5QcXHAOpvAKYvnXmb5WKG4oH
vPqeillb+w2ux4OVmK7XBK+bY0R6seE8Km58ZxQCWPPJxviY4RBQdYxtABX7V/3x
tlQElxQrEfU9cx/K9OzPrrokKhJQODrGe131P38Zje5RcLEiKT9HXoGRe+rR/Lee
okfiOIH71rIvgNuzw56UUYwVRzlyto9CWlydXGLNZC2dcKmwGV54iebcWvJiapC3
RvHUA4fIyO8L7TaW2QC9awC0IXhjzj0ThbcgQf9x8om4VyOUtA6pfjXvV5TpEfcy
mCHBtcluITAhq3BeJhCNK8zYubRM1rsImm5/m2W3L6H8ot/xDuxM9jdyhwv/fsi3
mz0FDH4ZxEa/ElSJldLqCNWJGiTEHeWUgoloO0ScqLJtuXv+rWBLwXuI0d0wixOl
QQqEsBoe/QZt40B9rX/sJaWHaqerWYjXV52QI9Ng+eZyPrz2mtBGJNB6VMDpVt3B
qW99f113sgVSM+wOGF8kq17suLl29SHZ5TKVxtamEjuwG4ykxMavFg+SPFgFadnF
d885KoUtU3d1tNp8rePeg3ekXt5ZrQxhLx2VuVh3RlldP71x2aOiAswOKruTEfFp
XKxkuHuwwPV9oyUm8aWLWy/oasXDkAmz+Rxb47+9MjPg9yuck6pwG0rtADV1ZV0C
7yaqTu0BQ4yP0aJ4qxd40PGR1iiTkZFvJN/VzK3uT+3zVhSHBteMaKVHHUJNJPU/
m/QQKZmYBJvDXzMSb03h1+2xMGnLyjbEgdeqaZfs9MAyAwhP6bvYqXe3U5iRrH7A
VYv+cU6qcd9pQtsZF3CcLU3bRt+UjBrIv7kk0DoKesIF5cOjdkoFn5Pi/OOkZMN9
GDXR+z7i4rRssZzJL4ljWN+4+jDxPikg03OI/D+ZxB/NFX4NaHrut1Zb5BM+uOh3
aJ/iOnPkfuSI0qA+XYvDExIljYMnMjfmGYUKOeuGdAdq7rHlv4+7/AlpQnH5Jfo9
zjt9hyxMRhgXbSXIO4MkUg+dNIq7F8HI8oQp/ul72uu0a5xHYCBgQZ8A8iZm7AMs
2uQdz5z+MYVc5hJzkWu3VbuUPCxv+gnOKBwwNMZACjL3iBY95v+VrO9+qolZhfHq
bYNXnxCiIDbMhx7h4gZIyueSb46QNjsQN6mQbnSijSx2ZxhLgRc4kbPS0Iv2Udlf
KvKaHGeU9XIYcsscOEQ2uB9HXrxpMcnAttikSJd2MiuIWSIvYDBlkC4DTql9oBq2
55oBCGiVm6hKnqPoWe21hIXbqlTfYFThoWiphOnzlSw0NC8D6mX+j6xoVuiipKbb
iG9/XEfQXQEXuNaaUuhCXJ/gk/ezXRlcRxNs/RNPhFuyrdyOSNSbYdE1pSGFRZW0
CtlkNTMCxTZUlGjVoKqrZlyFRbepUGUOxtO7alDvleqhRcShU2Ds0RntWHYLLs9u
sK+Gq66IMwrnVhlT2glEy6tWeGxMum2BgNR5FmmibtSVRR03HnAKBRCb+vcDdW5f
4FRNbEXEiCGnJbf8BkE2yCwmUoeeOQ9z+W5OfamZ0uM18eLZXNX0qYqbqpkrxmo/
NGSDPoN5u/qekQ5j8zjxhs7vA7mu+BOAn2k6O8ycADCgu0fW/vXr0anEC43+cuwH
BvK1xyLtE6yqAU2eMpv6nRrGiY0BT9vVdtF5X//ATPVt7x/NjwpWl85LXCCVKjUa
iWFnoWRIEdJyVuCKtMcJjCwgP0d79n0Ggkjb2PcEsR0Ar/DXi3rDldrK5Wxj8VIM
gkRPRrcbYsxdFSJW6g9JnNkDo+5PwxCoYgcmhyKGqFgWlZ0bl1fihpsOP2b/8PtQ
rcn2UrEz1LRaOgMhGxLp8Mi+L0EuttJiB1oOiihgVEaxbzzn2SFwpkMHBz9czQC7
ltlny5gyEtsaOwdxIP9TROe5j5EAc1oAEsxKOAwltmlKkLVFj9C/UlVo+ESTN28Z
a0wjGVawS2agCcO/Fo8opBVRwVsr5YDkQFKqEAYIwRW1Yf4JVNBqPaZsAqWNNKD0
Sby43ok77kN7wpZgzItem3sCVyXnnmigCiO+nxzumvYaZ8Qr4ztGmGjM0L68WXiv
lO8Csls2qx1GJCDsLhXscBpSojnVQxJcch+9lkyXf58xBkAlebAfd3/WUTpP6wwn
lHAixcu4bqAAkcvpN+L5wUEFiZmTqUfKnLOO6a+NhCc/YkuDYM3YzqLw6pyZ2z+p
sO1mcMV8av4GmxOdKtDqFraRiN6WJrURvABYigrhOziOY80TKsBU9LQHj4Rt+KFB
ZpQlHbA+eBx1F31htXqUfVtwOFj55iTefwrrZipad4xGfXs8J61eKw7F1QKQqIL1
WhcyJAxJ6uBnwIW6Vv7N6X35RH/T3eSCJuDYImatXhoYkv7T77PXhXWxvYsbpQDi
DI7Mmj+g4crfs7QbLjAfL99FNXrw6xxWTgyMCCLP5lpoCIoyrmCta6M8pB6rKdaQ
jXoOL7MMlygpeBlS8Zdnmah41B25Y/1s19Ha4z/CsZ8EHp0CYsdmb06v3dqtmKHA
DlzmXOeTDDCHciyDSoVddT9dmTQP807O2pgfE9TObEr2S5M0+Lar5Itu7AITgNDt
8SQEmfS4HdHondUYq4dgW/p7GHn7otaBcmaFYTd+j9XmbLU1mDtwB0OulnxyJLwC
rBQ/oK5xmEuB/qHsjtlvsqmDXlSBt9Qht7vSv8ZeiEQTN4OOzcQ+9AdnoB3bd6Jp
qMKCX7uQ3da9rlvTeIkG7G8jD8sYzX9holsF7ALFjW7pHYq3wolY0bDFMB7T4r1F
0j8pXaWXe+8K9uZw3wQa991d+diuzyCGO4vwxX6kpZH7bHIsY2G8dEvbnLdoT1vU
Y4XPoyYkpIU6Y99C8Fk/Kkm7IDoyp7x2HmaPZgnU8DIuKw3xvijFJxDSvcXxOPlP
ZJ+uhuEuwAiBHZlXy7AFkT2OJxV1KGVi4Mmd2X/WkiRy9cp4JRguLHdEBqud4t6Q
nm4uui5ddCYrLJj9p6GdxnIPBcXDo0I/U5TDWgixstUjlhtdPRSm4uom3lzGzGfB
xLkvf6jae2I6mW4880GADD1Z2Npbchnvq60Eu8tusaTXHATcsDC46zz/i7ViEvLq
03RxMQyHls+XbNqIDScAi5muFEJSqbs6POnuEaIR6CKrOch4+D+4oOhDLAmtQr4p
sf2MTHuMKnxUY7Ds1odjiBLL6QEwCluky/AhVWmRsBhNVMP3vVRKeCsG5BzQXheI
NbHwg4Vj1ofaDPXPpZMuwDBh72FBpFiKLayH4eGQ3J1o2t19Mfm5nebo7sDl4P7s
TZ620su/EiI8YXJ22Il5no49zkzqEbqIEEKGpKA7NO8JXzEWn00jA9CbOxkXq5Om
3ON4DEIucQpoqgpNOrcKFV+HoI7SsKcItls3Up+FNymDzPPYOiMgK/n7pXcVJU9R
TXv8bzUqIP3kBFGVTMpQ4X0WMnQVApvJRQabGng8SgvRdueIbWDNu/LR90ZMr8ih
f5kbfVkyYmOjAIqx7gRTAX4RmCcdlQOYC8Mfcq6EZSHKmliqy1Bn0YRMkRHDi7KP
VmJxMOI7G7H9tS85rh8HPIL0COfdBRLZAJj6b7Gria5oIGnze3BBt/936Py22XnW
IgXjjyYyonDfL/FETMc69Uxt5KKPukM+HD/n8a6tBR+fo5BUYnoXcq+KwmN2LDSd
GRdtODM6EEovjgbwhtC7fDrpRqD1n6gZe7IKmJc1fVlulmDTd8Imk6OF11+4XrNA
XyMNIiDwPrPReURiK4TVVkyx3Gz8BdJBXlIl2tEtiwqHDtP8mFw1MqN6fprUGJvK
Sg+hb6lIDkhM6MdWZ/GPdZXHmfEridD5AOdnDzCjHntrFtcnZNj4SS6Xl0Yze0/m
96ouI814KCXB4T/US6X7n4staEm5WYf9BHBhxzjrfNUbQ50EEimOpyuHQfW6xczu
VxF5cxk3bPtHY4hVGvint8V8+IYmtCoHEewX8CaAvd1f4phDk0TDkhpB1De1mUGm
eKtCjNcyK/6TSuMWwJbXfaZ3Eubldg7BM1RzXwEk6xo6StZ1sN7SeMS94aozanBN
GQ6K+9+i96iwo80ZDBKKUdDPtE/qmao6j4GnbgzP4q3TRo0FpDlar5gYI6mzL0uR
mpJikKc/9yCq0c1JCL+izGBbwvJgXaOdo1wSDxAyn3Do+iOSYoA5mkVxV/eA3glK
Cbccs1FAgIWUkMXwC5wDeUlTeLuYVLXP9THOO/3b48QLJa+rAhe3AhP2CLhYmdf6
TEyMP0NnN3faY4W/+3t7mXDhG+jF/iJxCnWVGpEvJ/rUrOulOVsaqkp8JDY1zV3x
Gf6wQ4tYJ9FBkej/48yGkjKcNKReiYkdVVNULWyo4gk5oLCaFisixL4Y7j+A3UVC
uB57aiil+quGhr41+UuelcpwI8ahCowE9WjDvsTipk18wtnhv8wmoCHPxbFj6dZ0
tR9G5r1y6ZzMY5TSMTI4kG+T5FTsVnr3zX3ZkSA1HV1sC6q7pz30xDfutXsvmTCV
DYSkwjITaC2xvzjli/ld4g0kRaoduQxWrvtVKKbEXJpTEAEMBCKT0MZhQASYhgQZ
i0lm2rWku+c6xqumw4Kr3oimqCmO8Aqemsw9tizzbO2qzn34VVMFwekpJRXtNzAs
V4RGVXxe/r4T+oQE7jJ7nPJYrWWMCW2LEl3JJsu4BVzWB4f8/4UfHTnzsFYwYQcn
nmjZDyF2F63CT1+UeZrdFB8L94RHjdgXjgMlpwrZ0j18WCJnyD/kPjRNn/yx6ORX
ZiuiZzlQ2SJAWoNP8zz77v+yJvj5iXK5b8oq36zPhheA2CV7aEBTSJ3hY5vQjtiU
OzHTyK/zk3mlBC64rzVu9ySPZgyoHv+Bi4f49YKTC+oHQPT7uSwSb0Y90nej6GE2
o93tI9wY7RUkg1opI+EHSbrisk0qxj5ph0IOKX1HbMDdBkRvVDYc+vMndr3b7FgI
v9Jsyg/o9JwsDZHTfcDDgCogD75qfQvsuPIZYyKpsmZDI1uDXeAPCPRat8xdBk2P
U0P3vPDJFhc7GQzgsX8RHnSXhBtoDBRZOnyUXa2FcjeX46df9PXIPRFLVajDWcRX
K5dPZg+t0+7Gluu6kpHUnsFrPpTBJ4JL/dfW/aCN2/bwFPg/2cPEt2S4RUed8yQv
tGux7cxSilTpkV3F3up+PuwibVExZG/jrlOJukSVp4KVrp/zSKjwKAUvx1H9lUM4
N2QIOsx8asPxd9TdoY57NJ6JeCwB9ncE4D31bGlwL7WY8If2VcLi1KFjpJGnMgge
3PVpFMem7R+5txF/bwnbJQrK8HyQNojwIPeidHh7UBHf2N6729ngSL9UH0cbqJah
TGQOqrkxE4fvviQA7oFVDWX2lG3ixQbm9r2BW+m7khhQAlADOHrSOxDL05LYHDVE
UihE1uHgfNqGSQm3mO08kRU3JAml0wNztSc+0Zta9wAGSDyvpXh5kMuZ48wpoH4i
yBhNwPAztH9ZdOyM1GFiHYzmUZlHN1c0qOtG31yDLicgRQiAfPn8ObjvM1IW6XGn
t8v1Pm1AQ9FTDAlV0jjyJbuAXXhxGSATCx3adYRT7gSoCEZCmD66hCgwf4oEP7hu
cmChZCEiyyxahuukFQrsoFMhHiXtJejm6ufEVLou6YH4OJF9MIYPJayYn8dBcCIz
JRVF6us50ICqvK/b/QTd35bKRIKFq07PhZyekB0fiZVy6BpPrHTtlHWFiZRSPtlo
2vFhBZCNvMxtZLoSUBeLYRJtVQOf9qrjAb8QayOyVBUOrRbSbgt8I06mcZvYkcEB
ZAnT93HWnH+tVEQOKnfJxTkBCgJvnriyZ3qmHkuUGLE2e2jnBmicyRc3JEy7pqZZ
/pKJvrveqlKsOsru0BD+fy84N+W23Xrp3wNJlk3WZQNL7mkKFMczSgz/K79Qw+p0
vW79Ppez4dXLklgMfd9b3Jgl1nj7ozGaBvEBjk89I724X1mXrCLbslijEOEniAYh
2YUE7coUkXdzQsJslCVJva/lX1uiFEA2QsnkFItcxS2J7r7uFFox7vXeIrwBoT26
h3E8QtAqTgMBXHGChMRIOkKaJfbVX3M3s9KDR6enx7UzNoA0P8B65X2Jy7eKvNz4
dxjk4faoGXeeSjFy0YkFfOe/bzrlYyvU72taj0p/+/KHIEFi/CG3HH7ZU5x3ulON
oaxfxzZqDM3DB5aW9dzt/AX7sitzH2hhLdv4Xd79CN3QV2fyX+pBnULK7kirIipQ
Nxvl2A9E7E7iib2orYrouzL1jl1PzB0owFNJcu8Qj1dU1haRvJntgwboJ7YgZpC1
0E2rK4bD4F9zNAFK+h/hJnjg/DDiLyX6at5ZvG7xZcUxvN4n6XFTqqwVq87DqNgM
0JR+Ck2ZW6alB1YXBHSPo6ZajZjRLsSf+Qm9Te8N/S49Qvz/xS4RXFp7ozrQeRq8
QligH7uuTyXu+LsqKYc1Gc18Dr1ll0aGRQ3GCLiAamvxz3RasfT/ZMBeUPHUhmFW
7CTZK+bco//IpoxRr99HdpvgkUwyFSEcCQriSwBGR3O+1QPh3XjGCyLJ7Q6db+AW
gVLjjudghTa96PjgybwyyfBa+WJaPsTx0wrQ1OXkhvmR6Z13p81d94nbC79XHBGf
IPd64Lka/rr49dqQz+RgndU6QU/L8ejfipbY8rO0ETz3jrpbxElxlMo6BMXtuefD
Km32cmoDEnGUUX/0E+D6vp3SkMZy3LbvuDfO8cEQeRDdyCuLPJ9ds0HH2p+y/WAy
lAQmbU2btj4fx7emyVgT0FTMWxuz3WW1sszddF8qK20P6ToXp3A/0fbq4fhwZWaN
mkJdLCm2V8eHKLwswpcBAl9/hrMFYuwAB7AVSltLbZMfn4Fd+FdSyImdFg4f1CLg
8DfjZOFPKtaqkbROzO0Q2IxriE5W8/rRYsbORT06iych+5bmCeGExJ4+mvSCfB37
OU2ir2WeW54roKWTiXHjj147zyV9+H8Va9A5LUPXah78ZaLZqtci6rIMaFSx+TQc
1r3jVngyAqBr84X8LVrHzKsCQHMHtRpoLLdCztbnG97eXIp3dXfX7ZwXd8nPwb6A
ZThDxm0ecD288iR0Fic/EHx8reMBsMmXt5Wn6n8X78MS/btGZMmSiJTOlbfYFvA0
EYLIbLDGRgKDVQcQBB5wYoKZqMO3EwnRzs25y2+xGUSpNtgi5LYYdv1MYkgDxCya
F8Zb2qUNA8EWexzIF+oLB1PFlpVCMGlBdKWbBzQkEvxDflpgZTObo/usUqhzzqR+
K9dKjii3rdbeeRMJm15Srf13cRU+GXqdRLsvFe2tNgSQ0Fv3ymWviXwgJZTpdOf2
CXcRLyfWW5kcgMzReDmBqH6nv9A/m6bqiFgrcc/kwA/rg19QKsQE1kVZJ3RWGLXM
xVLVrMTyBz0tbq931Yqjb/6ohnQBtrHc/3++9HhMbJ5pIKkKjob0MNQuFfU7YeYs
VU7oEpsayagmPW0nchWPrhQfjPFTyrx085Yp5nUp8OeQy9KuhdzVP3OtK/6hMbo4
c4jIKlBKYcNASIPtdIm9WjHGyqAvlGV+K7WQCQA6zKjdi4/eObMpZjxk6t5t1IYd
wPVGoErJJVn6FiERR4JQ3AjnrEJXdr/FdPfF6n1DZRxh19mnCpCaRJwVlhymUfB+
Tcg+7dJxE6M7VT2k8A7Z4a6++pr1JHM9zbxXt8CYAmBDJhkeW1COxi/Or6hjgmA0
NyKfJ2jsnhspYf3RbsSqLM2RD3MUWnSnqZQfnNm9Lelb9h+5DmuzwL7xyLnI5gry
8gvdiuAGBkNygj/OMa7mKGeO9/dPFNvVrRMssBMGPxa9ZZF9aTuyHmYWAMtnan5B
89nRlLviCLQ0sdjbnzjexqeZABWrsXqjC7a9O6oAfDcVodXiKf3jdA/Dqe7yoXaS
CI4cxrDch3eoZMDO1URhFSWg2zyK4qxbG4vGi2/b6R4otMtRmNiEHMHwQJEUTpNk
VUPqqwthejrZWpeaj1yp8NkWheqPJoyGF8YhXiXdu6+0qed0PFuNGuISTi5Z3jV5
Fz9SWy5LQ+FqWNDQpEUmnj7j784TKa2ZX3usKi3DX9lCq1gWPN2jqkTUC7bbuZ7g
Mv7FDB5Xt/OL87Il13O6FtUd4rREh29yN2gf5kllmJ+azuHyHmTU3YRKaolNEh/C
7z8D99TkqCalF9PjGtOfAVh73VjG6LdfwWUaUZ3F63zAVYR7JXEDR5L41zXMjMzW
vGQZoBW+2PFB/jvjMwgOmeEBYBu1PLEcqnSN6hBer4zbo3BeU+AI7fcr7UygTrlm
EfuHDmhUJj3/Coe9UUnBwD3otEpMrARYvHV/lxyuVI3P8qRXMDM485MPcFX695db
RKZGJk15UcMyavftL7sQXCTvsdHJMYiN42Ywe7YqWCh6bXEqBFD9O/bNXjBo97Xq
lr9ToA+5nmhuLMZ7kNR8XWVMlSknAuLR6zQ+QRCVBNtMqR8aQCJAE3oN8gn1PC6J
+/qp+sCFsZGjkpIMfAdCoiNTquztAm6gbZWA3jRfEnddxc6Pct5hk6JK267oiC1p
UKTBwXjPvCvi0cJYN9fUL4ac/dvTGPofxZrMtuqQ6M+U86shwjL+wATVW6Cnf0Hj
rxS7zZyRClfGHWo58Vsm/qD54wGzYjqB/8RChTvXqbRz7j7oXW0dwJGl+d6xAs9j
cnxuReUsqfVRmH43QammlxurFBWHCHmg0it24EQN6q1vQ/2mtu1kp3kK2nbKh/RB
YEFLkmyXFVqrw4xcEHmG401ZtV9t/VBnC3qdBSWRX4XP1atEhp/CN/51/L7DN4bn
PcJkzLyGzk9VrMlJL7rIxxp+bXgk/rsBlbl4SJAocFhYCu/Wn90j9EdK8lfOitJi
I5sZIh/sQm2e/TanOP0vexb6RrMe2iNiirt01YCX0cbX4+ycyJydpNw6JV2+78qW
7Ojnl+JQkk2psiyig4/zrQNMlQLJVEQO8VguXZxsVa3aida2gUhZRZnSfxlrXCNM
zhGq6+J0quA5k59YFcqEA/A9lfv/+s1/QF4xGAbaTLzdJBFaXqfs9YYFL/nc5XJn
+Ep97weCdw4KcieFKqRxos6og55pZlBda16Fjko2L2gpkG86bc2ZYkLIq6zJxABT
pyvEE1xqT7fpVjqF6B2RnfpEEk0SYdqPn8rDIKA4anbD6xF6f+NNQTqMvFHdBrSc
ZcJL1CPk4DDNSJjW0kwzaMTzw2MSWvkLBp1kxjBL3l7VUdzdoa5bTNNIBxhxxtTU
JsFc3EZ87eRbtX///5T9+uXmGtG4KbDxwnp85AbTL3xLJDbAlQMJo+BxrFqkgtYy
nlLxy7YnflFQjaubcsz+sl0vYtp7e+m361nwwK2MZo41kMEcSBTMQ77FtkDwsj+C
IdfhU6KPP2IPg9QJTOLpZ7Fr4efMun5xcTpyiCSJLd7l3gk1hH9C/lTFkJwE/XC2
Sq9CYsfTfOgXddP2as76FiGcHUmRaqm0Q2dtEc2SUpOmZDjNoc16ORva5C2Qk9uy
WtzuJ7UkxuH/dqzF4jHa/mX2GhLFTUrMXNh3eLMtDPd6/SO6LjI+ZayQvreT4b6V
CgzJsNYsEuLTxE9fvaWJaLDAVFnFvJrbTSlR5FMD5cYfjMz/PeYht4r4zejP7cfm
keWr49FvSr2AVfNUGAdrACxcmNMrRYHiVwieQfvzzkzTmoIY52oE7jUOvrw3Bb3Z
wWEosSZu5wBcyGOmfLUO902MqCQiH4pYsr52YQX2Hghu8dTtdYYogsIT8/d3qWPO
ucWyQq9nMEkAsAiZXXp0yFdePmRwOu/Yo/Zop0pP4uhkmUbhb/pQqui6CD0cCLFR
rWIPBhDQXV4AirGT3JDS3b21pj0lEfKx/WpB+azxzudyKmb2hYd2Wengsbcqkf7b
4tMiaKvHcowAOvxRO9jew8qLzQhvpp3AlCeJKLsoXiLvGo3WuvVMTmpjpFdPkcXw
CZ8ebpnf8ZNXOwAF3+m47eEZm+C+z/5cA3u/yijIhMfO3JQG534mldhSmVcSJjMX
3JJQJGeUwRxfkTlQ75cCF0vD3bTJ62pYtiEgy6AcFnjBBbFpxhx/bTH/UNla6gid
x23dNalXDIeRHvGqbvOaHrJl83+Ctb6VaeD3uipOYOvdz6d6L0s4q0yur6EqWZbH
4HrHvgA9UGgBXOwU12+A2B0FeyGIJywJMqdfo3igxabrSptakagAqSgXqqBGApzN
0bap9I08863gABazHfohu1peqxPW8+5dLCg5hsVjXmhpD+BxahHXgOwGUiOB98yb
Z6rNsjxf43MPpYkQeUrK2DpRV3YidP4ZukWeeu7AAM/PCCfrz8Y4LDeyy6VOoVTL
9568DDiaA4BiOM4kHymqLpczAP8N/5MVc6Vi/xpRQB72XMc/2qr3GOuVtb8P4K1S
uPcGuWoX/8ZXjD3KW3C6zX21Zu/CG6ujJgNrF5BYS3kJznu8kFouX1d1OEK2PeNk
Ivnkmh3s+uTdPfgzgUZMilt6VkO7xlYNLYF47y2yCcj+lxOxwkYaPclX1x0lDmMp
cxrLAGwYbn0JS3cS518x11WWbtilU7tL0O772Mn6boufqpKAweNn0+0i2lEK0GRz
28HNFV6r1hukL5spc7d1pTXyxR3L3PaThUYOqpDgNoqdd3Y3EmZl3+LLqeIC7S3C
RBMbo4VQKI+2l3mY4Oj6ZyXk5WoQ6E9aPeo8NP3UxLAuJe7ELSfsLH97duX9wz7F
ZJhDLl3wwsqRrCkZS1+BtU3+dnKyDSZ5CfELk+HSzW7YnVtib8AF27GP0rMbu7KG
LA/7Jm9mcgTm+PpMCc0HUpCyVXz5RdUGp46CbiXhsd+D9BAwtGJZaF6DgEIBnViA
h8XiZa+gld7aIvrcxzHYeAzWszkyWWd7gv48wC6P0/7BF84Or0hz+tfbSW85vf68
8c/XV0RYbfNrnvKo26legL3PIxDWYjUxol6Ji4GM6xL5QDXhIT498XXw8whilruD
JyabFhhh+6XVRgNIaEpQzxMqS53UcAugcEaGTIs8x31s3sFWP8r2PmXJ+/QgDNr7
1gooh4+fAIng9QeQPsy86JrSnr83tfWIwYH5tAIhTPV9u9sQJejUkHWiAqz/mEpK
yfJp62dYyuqLMR+BZNKGg4Q6yQTAiNJ+eK45JqxEvjWytfaS6THH0bJLgHMR2ooM
4/nyaU1SF1FjzdJPJNgmFRZLAPjxULSwWVzBM1xuNszstFC4iEYoeVQxVQT6asEI
emm01sZeXFPB9WaSu1G7t3XGnUOvDVFctbz+EbuZP7xeXcENxE71QVTk4B9FtYIj
vfoZxVg48tdhbGL91lYNG2+0gT33k4aUX9gEBKpSnmR9FD3io+rCK/BQQfTKkwvx
D2XiuCWywzXJpgnem+Uw8D0+eaDcZWlNMGe6L4sm91B1SL+ktlOEBjz3yB5ejmSn
oAixI6Tf5EfvcE0z4h0m7o64TBnjDsongVBiJhqm5aVann+CIxJfQvhb8dU+rqAF
ai0F4MvqWDAhuqKby5cw0tU7Zg6smpQf5YGqrVNXmAGjScABabUPO/OAFzP9DHcr
XpDk5dhknUxKDXUPAiWkDElzLG7JinyiofVidqBoYJAkK0iuHLs8jAT5aGgk7WBH
nMRKWl13eeDQ1/t9d/MW7j5g0XPOS/nz9oPEwqtIs9pzsqjMKThGe+yaUkHc9IKJ
R4bcMKo8ndFl/+66z3H5NFz1iI9SoF2DHt/9GS0oDnybnLtOnq68JLdBkEeCwP4U
7+OLkdVn0BEBcqpIRv+Pa2MptUTk23XThUGFe0vv7CLWmJWH8bpAW/Uv2p66XmLA
bvTYsT8garKZd28/BzA3w7OLJ5DPKWdj96+oBUBPxwFQAMvXz58oR8Ascs/Ggeht
MpPeXbm4mgHMOzHmLqyQhWWYP7y8npPmGrx/Qog0j+HD363kQ3PDm+zo9QBUGehv
PHUXEDF4QasUifKYmNQZXX2xH66Fq9D0ChdHpuP1+c72aFhV3TWnHA4EN98h2s6Y
WxHqMOfXwE2Mj0lUsxk0QA0nT0mMf2x18y5WtDGmnB5h7G9kgiDOnR4TWGjII4KJ
BIMdc5N0D6wvEPpLEc7s2CTxvnS50ccsctCXpGoo/g5HOVLIieE7blVGcRAPhddg
PcG3zLLWyaicJJE8i3CO2Tup6krS8OeIGTaYrKNyaPNIz2FT4uHhWL6POh4lB4YD
HhS/pt4aZRWcqU4GonjqbwhgPAZJzO9RsaQy9ZBBD91+fiAwlcLzOWlVPejmJHBu
NTu1kBbdhKPhFvYmZ/F22MjANBPHEtLmlSfWl8yUsUErtaE4CVlValbQ4hzMet26
99NpaL1K6T8u58b9G+VdljtXiGTB+kut0IX9wDll6LA11jyVf8QxdzV1THDxcR+v
C0LG87zuDvG6ibre4vwZM3d1rFCgnABTNLxpd7GMh7kc1sxVN69atY7hbBrjDr5u
wWT5sz0XBj/IiZFAFlJhnkRlxUvGlX6wKVGkF5Y7Ewm+SV4TSw3M0X83qQwgea65
p7zKmyyJ6WoBhg8L6i5fVg4rJAzfHjk53VKYEW4hAJWjj0pRqWDszalGZZxx42Xw
PtW8AZ5Q8tokKBECOsBTF08fsUwuvFAAIwn/mYMQlNY3/yBgb17rE8COTO6cmw6A
8s4xdyz3XQwC/0+Y02t4z7Na08SjcN6e04Y6Q58du9/mE2RNoZJG0GXYxkZ+2A+T
m4nk6NKb5HSStIdYuFXoQgn0RLlnxwIv3KYHCZpgExQfeSbnO0Jg4k+yTLDGufey
kMMNakK3DMfLoFpJh6WQFpZo2cPdq5HgcPBFGVr1nUPXmoA3Y0SDphvuRqRI1LZb
AWvxuNLm1HyYZDqm1hsS40m6uXInKp7l0Q41+RIAHIOQ5ld6RI2WHa4nvLUypCpk
OAF/OtPWa3VRXq8hxpwwnL802hkcbUtM38c7z3IOU/za72Rmhbf1SFzNi8d1S3H9
iePCCmVnO8Gl9Z7Lox1rMzjjh2lwwUT5gmbZMUfxDdX/lO0vVgqvhILD+EWqMdy3
WpbM69NLbaVrspj2d+DFtzCwVpXWIm5LuLl7JJkALja8zejl1tuvGm8ZapXDC566
o7k+p74pTdkNNAljbX2WjMz7sNsY7Wbo2+CWKaAj32qbo7cMquodRGS3ryvXA2VX
drKYYNWf5niE+0qoX5Uy84kVLTIfF23p7TU+t1kXBZvxOSRgH71VRz7vsjKAj67Q
Q4ar5KWPgdm97F4E92lgnIHRhjifLYXtfz6iEGSArNSUR+T3im+xhJ33/+RyMkmI
0ipCKEsFm48vZGu8qeFzzhzK5wa2y/R4iVpTzC/mS3YHnaRh4bffzS7Bz7Xnj9YS
OAXjr5Vv6ijxTDQvZj6kMLUv2qGOF6tCzcW/pS1ADwReElGvbGPuA2NSno2qBZzc
OclCZtQ/NPTVRNqB0FvxJKjCKPQm5jhXGD7k8npEEDA578aw7WVTfk8xTmcQsI09
gjSCPpl5iCiUmv78GUD6HpsRir4CYme6eHelRtmTEa6ctPgaWVYpbbMWJjdsUikc
TT/nWY2yHYfClf+kRHB2MIPHE2hAzzHGiNbWSrZ4EcNrdNF5TTi0XTQ5f9us/UEB
Z3FD+hwq3e32rhyfkfY4/XiMmVXctMZMxJ1MMmqCeMaNzEh8BmXUZvpbsvI7UnNQ
l8t2P2OmGQfhdv9PzxMQ0mfME9l4JUjdJSJc9xnoz9V6o69GTPx/HnCGM7XLYOV3
EBIeCpNCoyMGLM6XKNDhYpWmx34xtOYBIPuHiCPL/LxbvNNr3UAJIyZHXR7j1vR6
KlI0PlxfrCncNilb4y/gHo5S1OySluxuD7PPkOFW0c0w07Mzh+CEoVdx/FXzV2X8
jcT/nx3PidfRUZ+ZCZMfgIsOjkrSBAhZr4sIkAP7nyB5OrslOkDkcYsnAMltFVQS
h0diq2v7KO142hhSC9+dWG+bKYg/XXNo0j6aP/Y6siNhcwEH9QyWafrSOzyyV58g
GH2EYGvoJI2OgovEAwxjGai2bKQ58NrOptD7+Ipim69obkNaPrrTE/k+F1JuBSKS
TAOPYi6WS6BJ0sbCGHC2XwWPgj4Rmd5wWClztzxWRI7Wz1fqGxMjdToX0YCxwPJG
CBE35FRAPunPHk7AHVFjE7Vq8MJPHMH5tRvpe/KmwpPFFS8A5dYnpI0lclK0Z9td
2fXsRuRW1guGlKkKQ7PhPaeU/OuQQudlUgZGl40sOTiRj063PoePzUsxYRBhon0G
FxKQfX6T1oexbONjJ7YiRWk6LjQBj4UDFuyUSbD6QPI592IRdcvdVMsjYAM3T8/a
x1HAHpXQhB7qK+IeKMJ0mBsADWR0xadAFIJQBk7s09vkkRx7e8KO804wJEXMEap8
7cMFRB2atH5oHPDO7Ib6gh744AG8e7udG4mN1Tk64Y4ZkHyzRu65uGDUKiERisnO
PRSKMahEMnHWzNqWklaqXIs9cW/TZRELKxUm40sHGLjz89b96WBoWH1kXFBZjoTZ
a6CLZfrgYO5WtN3fTuzJK2c7xM8BYy9I7s02c+MRJkiMp09v2aPIvS1JUCNIp+ti
CE5++duW70992l4pq6mY5rODB4pLkzS+s4us8DT9pZj9H2DpsK/ltXjtkPe6HK13
vzP9OH+yU41O1/AGp6Gxvx7zfGFyzko481Syd+sPZdAbdTpzXOEqODAjaBEfA0tQ
0K7cKpULq3OZMBTeu2C55tnhYjWrAye09T2IBIkyvi4ubgKUtFK8cJYoVJSUJRu6
XFuscsY8XGEEYFQaqZ/vLgunvGUVeidO0lY8easCkW4I77EGSt+AM0bVyXndxieC
cUxVSxrrXZLcaJx8XS5GjgfxpyiMr2qRDt4tfasutpEUUNIZBc2bI8khkxHF0dd+
tahfXlRuL60l31iTLKRBtNN4OfYrOBh2uEotXStz3UVlYkHM0yvZGiPpDoNoleic
RbPaMWYBurBN/fGzyBb7xK6Nitt8uOL32KECoRnKJwoCaYAB97QwOCBAukOJH+4d
aXHDmrAn7Kisb3deTWCqvsNM6h2qNp63jDv/1kz/+EC0v0UbbRAnhsUkrM6hhSCT
3yYSO1JJeegPhMEYoPY5ctbmXLo40BEsQNveIEAleh4yf1CfDkEHySmQo3zPpJH1
cfa6rFC7HcOjKottd/iZMRAkEszt5omRZpUfHrmToxr/BzYJ1rxvtzCmo4cpWDeg
0LLfURzsrVnfEpzsKpxv2IUm2ISQT5VhBz7GMN962k1cpqp1l0wcQ4tulvRajEaC
SVytlB5JJq2m88lUmuHdEmz2GuZM60V2ro7FkYKqImvjmF/ZccQ0kcQZEok8bw36
0lif9sMwIwWmoZMzWU8dPN1/LYZEH8lXtzo4mq/9lAyDeUVf36H+Qz2oF9rnWVY0
spaHyi+jYicICL+ld5zLWgVW6j5CB0O2WDxUc/5jJfL9CXyQhZz2L41bxjRhQ/W1
6tsGsmSzc01Cb99ZAXrLRIl4YD/LZ8oW/cjQzA9785xHQy4OtG/+GoJqKkFvvbvh
nUZ5Rhzwpbpu9mVmxQ4cHAhnqoyZiAgTTm6CjxWLdHs7dbA6szxTtlzjR9mCSvOi
Yzikw4iI0XXVzwvkBrpSSL6kiAwPs9CIkC5JlgRRDcApmKk/t5DV43sKIxmPZyab
OLafXK1gKPuXBcE+269jfuBz5W8SyMOUNK+2v/ultSdmLJzPYPxQun5gyDt1oNmq
4gRgAuiCJ5KVqYwPfsX2owvjHjxKTLLgS4+WoZhmUCGP3TWUHC8sZp9xvr0H/btG
MxUkBU0GsUGagei0oTG4EGOpMAIHgar5cmHmD1j2mNnan5oasQl8eN4wsLi4aaOT
DoFDRK9bTmfGl0GYFidH78dsRMBJpDS49fuPlD64bCzeuds54/bqB1vWoPztumc2
i9q0CCt+eV/ouJQV0OgLPpPml054Q8+92OF/Prnl8obcHmNK9dcoKiC4D4IY3TpW
FcvLnJD2jGna3VdBoWCOi18TLXzLkGKmakTPNz9ughPTuivkWlPqYG90GOwOfRTa
syNuUWmr0k2u/tANL8gnrXKdYPUlLQ5ltUOC+vbqec7/2VxM1CrYYWhg36fTV/ZE
e91PeDR2q0ig8Mz/4Zz7KlzDWnGXxCSix5erzBsfBJvENCZo+OmCinl3qRlNnsf8
dx30iHgnJcyKwJa8yOAzisbRvFY2bGYnAAMvXziBJem3Ief7SFlrNliJo4hyPnuC
QRzYw/Dvcy+c7n0D/0m3kMiSpkQOfFPB2YiaVwuLZmhLTSXp4ERWiRA4VVRz8Uw7
Dri2WkMFd6Jp4nNDnvTm7fO0rhpUyFOD0crYxIqFhyRdcoX0MAYb3+JoQohPI5Ko
Eoqujk3s6wCSN3JtNLLIrl9BYKuacI2vaRqml77BCUa5EjzLoUMuoXA1MQC5JXNR
Ov6p0Uh4MqIMEBbVXu/yIyqd22GWXfGmWNhEK/Qh5WK4ANuZa3eIi2fwO3I49vnA
S379h/d/uEhamMMyCfqUvNXxp6zYGIQw4AOuCHN0om2h8D6Ojk2ZkLWky0zpTc0T
+vxTkISU4GjY2NjJvFNtZEKwKkt8ZY7DQ0BTRcLDWLUWjz8yyiRqnzJ8/A9XzIqH
3kdhnpwlZKi7S/LrbLK4vmiVLg80qVgoTz1nEeROznHcDNKMLhMf00SQffLDRxsa
6JYpZkQ3cm4/M4Y/LxujK57qPy8Vur3VJx8B/0+ydVGwoDTEhNxf3HcyF6k8yJBX
r4yFZMN6s2iLEW/AwKr3RQIF3qheMUpIOH2fn1AJGT6M0aVfecuArSKRVAtfB2+p
IoQaI4PS7Qg0Gxm3+IURDMz99ttRT1pSXy8crvUYRLTCQmwa5auNLAfYcXIUyNuj
jUcRmXwdjvDzru0Fcq63Xt0o2edaDEq+xEe6opAPynZSHWoTN4zWIWd47cT6YFrl
CODjBuiJppOciyoZw4WJ2caE6K1Z+t2cXRyzT8mTlqTOBUOcfSdwK2QKTcTnFKAU
zDGVrH8h+2e6RO9TpYuphFMqVxftMZhkv79xkc+fYiOvwCnbz1wToRUw0DscOmMa
/fMyDYjI1G0XKwQ3+wSISTeJCqWd4p8xtY1b6HBU1DBUi48hTcPvQUd3LiJFb/BH
cbfT4ZSevdiidMagbRMRhoBi7/SpNPQTpjeioQI/EXMdTkfxnE0JkDEdDr/sE7fU
v48eC+ofdgqBJQylPl6Ud56OGh/XaInCFqX5hklIV8R4Xp5r/7BfVJbev7BjTzb8
4ZKCQlwRR1fEMVKILnSgPHHwr0Pr6V2SLADR+xncYoJUFMo9ibFtd26VeW28JRZz
u2bWKEuaj4UExZb23IU2x2nRstvaCFRhNAyDlncF51y+cfko2MVH3VNyIrks7wAI
DwoCihYigTM1cmTvMtZZLGP6j+SYPM7M8IsVTSpp3MfgJR6ZsiW8otl/GQKn/mOP
uwwyLq1qFAMRud0thDcjVIgFpRWjIEJxDlQJYMUVm/0byM3Usdu6fjqSFGYymMYg
ycO1bFBJCSZEAzvPTspjuRf0Mc81X5YB+JLeKqZif+PzvmCv93rnzE5j5/BLaeTi
PNF4zhYMWfN3gaK65xUluB4YosSGFfK2LjOYYplTzg4iVxA335dC+rGiu9Ket0cW
ok2+PGl0X9DiFvYydtknP73Z7PhtvFI6Rko+txC2EoUe2cBF/7QBW3JDiBM1/fWW
eKPpslsMJRWS3T2l2Bodk2eADkIT8vKiekTAL07FbO+LE+2yOuttJzVuWuTpuicw
72Jatf+eKESwQ81ZJRo2yGObWeV2mtkoOp+i9J7oFhfSInUwTvZt9HS+weskDA+S
+KyUP32lAqbm3T8qfKQQofKC53Y7JGGzUnmXDl1sie7oovk4Mhpd2KkWZQLZbYO2
Brm9SeoSJVi2FLAkPHj89NrH6IMInkw4nzsJcNw6sQvTWxfemE7ph5T+fEhJNDSj
n+QiLdUjjcK+stK5SuNZTJsW+Yz7Ye6uicFjI4Ulr0b3D1K1KzonGPUIddbxtRWh
6V+5ElQNu2KSofb/qsZdHH3IkOVCHgJRsMT+3jRsogL3b+NqqLJxgZ+MECegMbb1
DhJliFISTB0cNeykXOSDGdFsC0hGN93LVuaXDSbttoxAXUDCp/h7bsKPv10W6+6a
j65MrMWEH0Qn7yT4CgQ+oFS+gUn7hbPdo1HpKB0pqVoYS/VjV+VZaAewUHJtGcZH
G6SMWM+nyqiSkk4Lxkn2VHnlxUFudIdNoV6v4yLhGFjS6YYDkF7EvL8tNGJ7hhx3
g5YbCGFae8KYIrWuJyrntRGLFHVOMtoCIRys9455p6elDYIIi3UxsWBaArC5Imt3
JJyqS2+CSZVEQsXIZb+ba2P87NetEadxVcPA3cqbH5czXHzapH2HfLzSgxtkd8KC
9oZdH22NzBLNg9AzFXLZoPzOafHlP7K466m4s1oZqEdKcILCG5NfUM6KazwKHmHH
eWT0V92v5zIatwwlIl8Cti25qbFnDVqYjGNMbla5CkYNgFpKGhCT1/29+HLmAN1j
PBS/mkH4vBDAlMFkJZuTt/F2yNb7tMkwCSFbNyfMq7WYf7HWqrRLfZgAkyEiUir0
N3bZx6LjrqO1GmqQ3Pmw0TXbB8AZTb4xAq31fUKAWQubXqzEaUACa3yRnDTa7q9K
+IYY3CDafAZKcgU5J+YiQVffOuP1G3JtnB5UsmlxhOA20vWsQ2yVPXK6NJsF4Hvw
KBZiLyYkM5OvPa6T+LyeqeBU1c2Q1d0/qrPCAPtHIUn8yc6RSFM7BCm33cAatRnj
hYuUKkACcO9SIVT3s08nD1s7FnbfwborvrW0unxzEQZQWNekSGAjM0vn9hQTepqN
zvipWSlU6XlQibL/kXkdymy1pYOAKS4k7qga8l2DSf9U2e2ZEtTAWiePPJxfhl8v
CfqUOOW0VFgJotRWGagRNVNTaGC5BHvrFIsWonRHp21jXM4ZKrBWszln8tVksL4q
9RsaMUlZasBYvIibtFBm38ejM/h5GNyzgbZdUS+bflu5bsfF2v8swfeE1JpPrXq9
lrJUzRyRATlbIFYw18O3sySY30jQCXqogeMBVIcaal9W6Njef3V0euJBCayNntut
DQtX9vrfcfPVmxtnDVQYCuSYmAn4h++lPDOyMsQQh5XbA23oqnSQKWkMdAk23u1q
EzTm13gO95Eq1XqyVVfxLgLapjuah1+FuhEuBU30xI+AJTpdW0d5nVmIZZv1c/Ne
JFcICX0PT8waxSKjyBGkFqqv7L8tugaxeT92jaGXrJ+Kmf7jH9h9NV+O7NbwNoaR
Br0w8HfjU5XUFpfovAOgwjJgyVpvld2e0Lbdb+6HtQG5ehxHhHhP10JimH9Q22wF
olKYyrrd7YgeFP/f0eQcA7A5kGgRVII8lwoJqJUEZ554tENlvP4wUJu1bkA0iiL8
4grWBn40Ajob7g5QZJyxYud2qZCTsspfPp1nggMpDgzGHtRb2s6BXGfwOUMBGfnN
NHc1J93qBsBt7hv4m0cfX6VwUet+ihzdo7+eO5nACGPFfhyTKTD6bYPuaAb9uq+o
pE1SmDVatO5JPlmnymredcUGuaMUUaCRdoQFFp2iCthW5bnoCWvU3jUmz/moN2jC
SEZk4a1uGJot74X5h7Uv83vDY3gy65AResToLZBzyPdm8PTSm6C/U5TBW4XUgvyD
pGYt97Kzi3J4LSXDRyC/mRJTcf7+uPJaouuBvldjSjqba6qgVcreyi0v09zt19Vt
+knd+rT1vv78fTjl+NglYYtchBD4FdTWKZ2KGSRpui1gY80G2+AYgHNRaCQmf8wI
6cYj6f6gq1ti3kmuh7TM86cERWaBnM2VmSllyjUVWnMPaQ4F6L4eTJVPQJtuJ+Fx
hDclXWJ3HZtsXzMxqICeja0LuOopqQsF6edgsMcysVTqqx65p6ldwMMHyAexJ/W6
F4m1axWIFvBQxtowOsXn/64/44fQQJgt+x3D9g6i0MM5SGBSXuyFab3lAybk/xVT
hPwlyk3T9G5blyqU1a9EAlHOhd5AgQhPPvn7nKanOILhyw3wRsbFX0UV+tdk2YW8
xrjWN1qMHogAbfJgmmaNecrR+rqDk3HxumV1RuNi+IhwIFXl6A7MWcr/E6vY7gaZ
O+ECKKK6mY25BhIwk992EN3znz6qdUIGxziRugiTympXJDUjQaqhgK9/x/ZVOBpi
WTIQ2CUugBSeh5neS7HIErwCx62eU8QKejJOsSMs1gNEFpbvsxC23wsGsQOhS/xT
MQB6Z67KVubV0DVuDK/8fYx5RVVk+quyHbThaqqQV1zcdVkiNQD7bbn8923q07lm
1qp9avdPfxzNgZMDwZqXJ4T/3VkrXOi504X+g7bqV4nQsOeEyv3BisZOtisaKGhA
ybjrPj64jLe96OHB5Pt3l7jntoyZMzeji6j2xJirQzoopoT3cFaCo+YkfzvOLZOk
SS3CNQuzGa9ngRbpCMtT78V7d85lJZQwisI6jJLd0dp/eWw/4/aZXBZDqu0CVzuA
5cItrzNavH0snu1XL3aGaFM+hUpzvzdltDtRDS4YTsLL/fydv7UobcJfvfUNjEN7
OrH2Yd2KprwzYyhBL73IRIBjJHS/9J7Qz2H0lIVydZ9oHwsHef3gZ/D/DNUwry2U
aGH1OIq2Fe2uTVF2/okNdGdKOfMQXwygfgkH9gJDCAOfxfJqICsh1lrgSFNcHin1
R0jnsRjr3AC0GRgp6q8fbVdTqwwRXOXIaPuS/ykR74FfAcBqyAFC/JPIs+KaEMLZ
stK8AJCshYD3ulplcvy/qoLtOgTmTpX5AxfNDI/nXNoUs/vqULnTt5QpM4v9TNQ6
VySTNe03Y2N/qOKK1zuXHsAA+qX8c2OI8vN8eacz/0u9fh5AzDe0N4JnDBURD6Vo
sJpaDSnckmTO7Hw7ZwW2jkneWb0OUHLH2efBFX7bOfseu5fqg5btat4m39Ij1Twr
YtOnG7qqEf1zZDmIX2oBqrx0rg1OUxlCXwsJvM6mCexEV+Xif03cx9j9f5hmGnay
wmYL45ap22GxLn6+5UNRUWRxkfSSCioLIL8l+49/uINve1Y5RBvQ/PveVw3ZUvsZ
MUrKA6fSpIYmBbV/atsSI+nSpgHYq7kJE041DiK6Q9hKFz7Gr74DJ8xmvX+aacCd
HGyBMkwtblcufdEWp6LcWSPuwa+Jdasx+N8cFZ6Gbiyd1X8aJ396gAf8pWowI4I2
/7cMvQ1obdYDkPc0mE9SnNbIKDAtPe58baM+0PdnXbc2PR5nYnWJ/wYa8hw7hHbX
oimjOOZKKenrxJa4Al1px0Qc1xtksbH660s6hpoF467nyIaLYhnOfnihga7cY6yC
s1pmRZzr1wjvkNjrz/S6cSlHXCOu6sIC8iaceF1DnrJOtNFiAtY/n1iRH5Bjli09
ogUsNIfPGPvphbKZa3c4wVVhmLOeTnOKEZVeKa+cpAcOA+bsgyARJiTye4x4J5l4
L510hav54wPQSHPf3QD5fF8thuDfCP0hYdCiTloUT6LPkbg8H/VdSeepVAxD347C
7q4gNgbY8r8M/C0WpX5nEU8ji2uLeOopJsraILSKZXg0QTpz/w6DhcgznRSoq8gi
8LbneznvZuRki5xvQHMx30EjgY0jZ/e0STtJYeCFyGSa+8+aKRwtjTOJ9SnJ7JVs
myUXAKZBCXD0l7Ahwzrr1XHlSiRyRCYq7+Tu7RDuOWiDa72dcvsizgKewN8cRsnx
gaJuesffHtLPSTpeOjGtl2EgckSs/f8skaKjEY5E93zECg+V62nVoESR98Ujfc5T
U27eYUvr/nHqMteSMnCOZHvs3wah8fyXQd29rADwo6w7vAcQMdYFgsXyQmmlJgqJ
Zby2cMTq4oWszAPouFT2p+oFZF9XlRZGWvEe8jzQZkDP1RE2nb0Qkj0S8LdcH88E
HzAbO28og8zD746ARVlHXx3bXxzO5NqlTy9PkIAB1r4Qpu/C+4zaskDhCcSdrC2w
2UGjdFwEepAH7yNQcloM2gZ5ctWB7vek6H+InikfHQwMs2UmdofAxYZE7p/rY+RW
qQYOd2679Nqq4WYQHX7J9qjKgnb3gyjWs6M8WT21qsWP4fWDQZYhNE7r/durE/o7
XmhB2zA7+5EUnY4UgUeyCOKu1SZAwa1oHzH4sNNQnqOhfaPlCQxvpi1I4KUV6s9e
5GxBCXWzqMzT3wGe5OlepCD6WsQnOVI5PBi3byqzoBZGTd/ys1/I8vjMUSbPvgLS
qlrZz6rvPqus3GyFQc9NGH9w8pBnv2ZXItVQyy8A+yAO5HAl+06bBP1Uq/hTydK2
kAqMxe0EdCeswikZMkBqFufgGISnGXNBoeb4Umd9wmKbIOXhM/03JmqCCnsBg72Y
iTvGL4I3y6t+d7yNdIs+FmI1sP7rqlFdoCtruv+yfyfNcIQ8fx6FdUsuSHwuO5do
+l7J+hdhY7S7L04WbhCAGKNZ5OGJnfGlI7Cv9imLGTSWipC5MFsderCx5KrgW3DU
2R0iDOX8JOI/wztsSkr+Ds63UVBs8D/l5A6mqx1iL5c4MatIO13DjilKh0522N2i
uAf1FnRtKx8b31KCYxldFumigFUVe9tqI5sClYlvDEdrR7E6zot7JfEX8D4Q8rmz
Eeu1FO7vS6oWICA1tiZd3bbGAsuPtglGDc4lJKCUO71ub/rnjGJMCvPuDBjzCxsb
y39JW7SrNVpRFURrM5pfF5QQi8pZQaMRKkadVi2ridUdNDgZ3VoW55NPydPi1+o6
G0H5+pkyzsQ+4dZantKLDiGO9V7tnkK/O9PIHV6uzDZRF/0Cy15plHRO5Z9aWv43
wPssIAgSKnzjP1rEUqn/+ZEsvu2/hbVbacFaaJ4V7bpFw6JCRtsdrEuL6dUuKONJ
oGf9/1/YwIBOsMwWJBZpQ5Ro8vo6T6Kt3wuculkNIlTYEC6E1yyZDa6gYVw87Ilj
M/1q4mC6lkluBU9aWMXpkon8yFKezQ34MW5VnMWbAvhXHGkyMXmrmysEAGVwnNtW
Hoz9SV5xjsmeyrZak7tD9/Gx1zkd4JCRFNG8bxD54Oy7utr6QuszCtty24ZAjVQM
CqEaAXtZ2kKYB5hBRJzRO3yaWLIhS4DkPmOCglUaDkoGK9zCYcbf6qP2bn/orVTG
H7XZ7drWSFCCeyeJnBNMacGQcEiR4/CYtN1ypXnkElop8vjvMz0svWNLZTS82no0
Qc4b8VeWAp0uVS4105fGTaC5x92SsT0A0V3BtYEi2e2C0bAtxruIu043GXvDE1LM
m8Ud7hEvH5Q00iSf2HmduMr9O0yeBQd104NHUmrtpKwjP0J4y2uYHpY0Kogf3NOf
UWNshaGGtEUPVON5Y/cpW1t7zUtinEnuuPPHqbW+KlQCOzNOnJt32nXMmTHLYx32
iSBfq31U/jdHKqMkMdDJ8YDnen6La+YKBEzBwaTsJJATFNY76l5CTijoHBj4CVDV
8IFKMslDND7YE2OZBsI5pj70xfglOPlwcNuTd71onlYPTO+Dy9w0Qac9azhHYE+h
VrAKxY6mYTWcroM4frpr8uPpsP0jJTpov8ThrR18IaeMDy/EAJBAMF6v6Ywp5m9m
DfHePJB7jp3hdRk1PtNsbAd0qcIaUO3MUuQkQVf5VTKMoUY+uFOAeGcEf8JnenYX
tSS+XEeNgfAQ7SOD57nR9HMwa0ARv7iYoHi96+4qCx6PmkalJbthtXe220Hf36wy
Wxb2/kL6f02yCmIFSVX6D00c1UZ1IhxZAfIw0dUNVRX8adDLrMANZ0skeOJosHCj
hpUXz4uP6F0yKa+vj83Jxsx8P+b2ZojdMXcYKhUXDgKHb8tS2Hng3wQFRFe/KPdE
KMJAtL6GoMfc6voRI6FrZNic7mQUtY3xu7yKfPQ+rpFNsKntgtMN/zXbaZkJC16M
EDa1IdyE+pN+2F/BjGiwLqr5qO6yxU0W+JS7vrKgdoCvJBp+Jxia1vu8GnarbJUo
6uIAeVnW8XcArgF/RP1naKJqyWG59AtkHTYK7fUst1yET/yPkdY43hFR5dr4Mjgn
g8CZLr/ZMtsxcjdqaMH3JhRYXXE4ljA3BdZGpjrX9MK31UD8bzZHFYH0c78fCPeU
4QCk91DOqPtFtWCiDZxOc8RgKXotbGHNV/jG1AKmIp2e/IqlK52fE8ayamVYo0xY
dEIzxouWOCzuTcogrhJDHMhmsPt0WpVJI6RIy/ySinU4YvKMED3gnFFvPnNg3At4
5P13T/K5eaWP9KPq4bKIGdkL5Ug5uRXK1Y4vze6qsd9RvOnJO+WyY1eVOefYKjDR
nD1uaFP9oe1zA1lq87hWS9ZtEMY3+563h83BEWTPlIV4IImTuV8wdpOE7ImpTdt8
Bp0d8mrgw2y/sXoXcX63qzJqEJYZSOSiSs4cte7s2AFpp3gw28NLb+/hyxcqQO+E
55VPM8a80Qr5JDARvmJG8FrdVJZK4YEIgQW4wct1NoLzkI3mYe6nBps81WMjJhaW
WW+zm0tELN9/CSzZAlokdEFri1kvUUfJoCmmNA8u7jSGSeE7cbCxV/GDuC3qfLRo
AzDnWskPd7ii+XQ1sbYZErVW4hnA/PqBbykm1Wxw770WrdtfAUSl6251/jltoZOD
Hy4vc4sL44uN3FfInDvi9WImXXjUQRr53+tfKtESEHGIcpG29cyFE/qugbrp+HVc
OB7pbV6e4rk1/HAURNe0wP/99kmGUtglQIru59EilPUBb7+/tGcTNV0KPL3YmU88
8buBLXoG/fBbGwSGU1ntVUMu0GUUFzPrNQGz1lx5cphT1Sofg/Tu9zKx12U8BW5F
FMSgYEJs1wd3RhnDUXKuOxXpF80H99+8TiyKxywSPlJxjfsR50/bWXwo4EyvUn97
yQdX7kP1f24j9TPOSSkcYXGD/Zmt0npYHoh97II8rMpmmeHy0YMLXc7ZzH9Jb8Za
kV2OliX3Ol5MCIlNzD4LNbF8CtJgVvUrVx7IGs3/1nKLdLp0UJQ8QAtlj3c6IEY/
KLfAZHa5rZL1dJxCYV16mi/Kmtc55PRc2jbwQHR9VO2hvnb+/CojipaVBLsf11Z6
4d1C2ZvM2Ss3L26agnXCRbF0EEAjqKsYMC8PD813pSKBxyrTKuS1v8NpN8K5+vo0
luztG291A/G1/sLlhcSk97dxHRaIUB1dtD5rJVsJkn+i9pUlkc+AHWpdHLzWZ/ae
aw1TMMbCYrQd5YRTAmrM83api1OLiwmM3/oJAUttm8mm0H/P9+h7yxEkc6K3BRv0
JALseDF6iSFCe4cH/d4N6nSHr3ahU9b7TZ4h1oz+7giMaU98IE4g1JMtdw5YTCfE
0+0iUICr4Oe7yj2E9CEajzvlgJkYgiJdt34wS3gLqWXj5FGoifsWDSfUs43VMfO/
HFomkgRVg5er0DlHmRJjI+pwsroCRDqNnRxjSalbq0gZMyvng9WtBf5KGYVJGDHq
jhUE4ZtcbO0V3kPRI5PG+JUd9flE8JiyBs7m01hJg33vrFba1H///RBfXuN+w6VN
L2z4zt0N4vdLWyKgmpx3Kft008G7MsopYFQu18tp3LTl8hHjEpdWk6FcK9GVog0p
+E08HuMlXDphVDgkrj0nzhWIw1pfJ1686eo771yYhxCeAiaGUabj9uN3Xgv0M4M3
xJvnzi/DZTuMYycVC5sn+KrxSS9NLgYPqWW1l1UUAhSCtWvyvMkoWpj5R7ww/i0V
S/vrBMXRZ6EyCUdKNMla5Xp6Jm1uLa+h4a6M+v1pdhCF+QFlipLBsinBc2j/Z9/i
oyKnu6KxmIaWDzrtQbqPjzvk0zQpCBkk0QkwaWp/CRell2yAMa0aB0bd+IRvk2SO
KvslX+bGEOyZksZRwxaSLt2I37c7HVWnN2JtqQd5O4mMl8pfGyCvnxUq/4M+lQ69
CI2dyWs5y6hnEEDfgDWwQsvRUWNaz3Bnv/C2GyTe2XnD4v2hXf5vwPU+gqhkddyd
N8vxIiWhRsHD421sv6TtjLeRhbBwJVo5fLVqmJnlZV9bbfOm9PrsSuJ7aKTc8XxF
rfL2PKNjRsnP9LUxTje4X1JbHGfiHPel3sI+dijm92/y2ZLl/vJW9BqugvzZgjzp
JkxerDqJ8qd/LIwPQeL+35bjRY0Qh5qdZsuQzjIqG3b0H/nGM3iG3dPg9S0aLzA5
X6YwmBoa+hZCgnx39r1tySEFL4pLKfcD8sazdgFTCUOfSfovZhvpjICG5NYiCH8R
tJgW7zFtp6c3ZoBzi9xngNRdVQo6SjRKWelyCwR4sTtmTXSgXZeThVXmXXqDCBLA
L8nCrbvSdceln6qnzxv0bFWpl+wbc5mb0dvxaktXNHXb7fAfT/3WYo1KXOVE3p2M
Pn6wQf5ECEd40gNetht0A0zLH8zQxuJE3cBjx2g0gQr5QTjoycrnGl3vOA4w4qxM
M7PdREdKi7FglwCFFKajBTGQWUaOkonZM3OTIdD5P77Zt8WAbVcRL3lu1SVZjMPE
sJMBzIeElC0TYUgiwNEnFXTLLeKuBzqdk6r5jF0p+u9HNHF/5wIEk3y/qWH55iUy
WzxLFpd3tv0vFe/tEBU5Fsnq338bM1aKOVmSwTkGM6yc3lJ1YBmgA8kN5RRj9V4n
GzSJYufyx8O9LGyC3sPjfb1o+PNO/+HYjNn0cp0ijHxxVASSUxRdcQTwvCzQZALr
ZA3J3u1R0FmgAMSJo1FKiYjCiEwkLboyORN+5uSuNAYcap93XfCvm8J09ej4HbRA
eXJWWvMv8NUGTLs32BkIc5fVqXLDq3jD4K7cx69sHqh2A0hUYqGiKlX3iyBwFmJt
0vsURHHcFX6IT93L+g/emr6gS254pkPBEE4PSiFzmWWODqCF/ql/5iFQkvbHW8fK
ebYLKkUizJ4ECXhT591Km9ZmNdpL7Ot4ceDjolAcIsC4AcJ6CU5xAiKA83NbyjWB
zlRPC8CmQkQsqaoCRq1jyHsumab/DsQwUwy2TgfHOAS3RxtEn+OJ/O/OTMeUOduG
Qaf/mBSxMOA7lfOEo3Yzgnq+Nn3xW2pa/3yRs/G3d8yApZX8xaEZkrWwumaBrMvW
wz3Ci+Knqp/EcHURvGZSTCOD9xIrpWHZq7VNF21qaJ9n3DirkRJT+cziFPA8WZ9n
m+5yfW4AcHpwHgMBRTIzFziRGhiGiR8CssCgKmODBZ57ea10G8BH/ua2cxgGwGBp
kdKmFdpTCI96qF6SOI8ofFOOBIOpCQxihlslXrh9YGnQupuu/z1dI+SSjSLivXes
h2XQxNGFg5JyhaY43wk7SoqIcNu3YtcdWwuSoeAIReuR/w2GAGWzFUWK7eZi+VYg
CH8wPlrQmbsocH6QHXJeXsgOnLClMxKN5GrPAInoHf3MKvPT5AhvJpjMdPraEnSL
qV/Ltlj1uJ6vKtcCN8OawQTs1uVAZ6HI2HkMWyUlxENfn5gjMT0DhZSHO6aFlf+e
O7f6y4KODqKS3XuRIqLaixWsmWj+j8rYORNm+XWME0K+9rCvDfNLZ3G9UIvq9tkr
8l9k0U0TuKXJsURHvxXeXJuinDQws0DOxgb6HW+lDakZ0YuS8kLl3xaCLZu5Xdo+
K1Tyzu9aYlSvuChoHfMC1elsDZRWtMQnEp0ETslrN+HLx1ORPUehTOHYI6QqRCck
p5cNhOKpi7DPEHkCV2+5u9apa9t3qI7mylbEzJf2ommHB9DG0EVDCGQhC6T4y+9D
TMTO6CzJAtPDqfMad+BvHMUWzd4uE2dYgaS8k54PH8H4S608PoukiUOQJYQa96Ah
HwJ2Y/sb4ri1PRm4yuvggkyx1+JyIQ9T54Ya5BQyyZAIaLrqVHv9JWZdUW/afDtT
lL86RNhRvqOqTKUKPSzUcsYVBWWo20HcUOnsN2DtRyjLB7RFP9VQ6IfqvyxPInNg
tcG4Q9tyMWfI9YecqCtBlz5N0ii5DGK17R3raV5+fyepB0Qx4iJ60sJhkxv9p79G
8LoSLNzpiFOrkJ8dA7Uugant5VtODJ4VXUZ6eKep75wcMo01Agm8rTIbTx0y6c/4
RHnZOY03apuFD/Zcu5LlLjCW2Hx04jOCcBnKOpf509YyyV7iJ+WjS38RaEwiaPAE
B4WJ6gsjW6Ahnipgt92n5K9UIeFLy6fUbO/7cHKtr7MbQv7n/rOQJvyfdTjs4rTO
SoFFajnflONki1VItN59Z/eSsel74zdgem0YD/SqFK4xu9BUf3zSnoaN79M7Y06R
ZxaK6p/ooXp3JQQ6dm08bDILWzlYI8P3J3iZyRwZC6HAwszyjFW4rnYMwdcC8+6Z
FseGnBYemxb1eNazcn3QAieBJBpeqCb/PaNGOlWpevohtIXDqZ++5ow214N0dlJ/
WWHsJCcC4A19S02PT9X6KCShkNAWppsQz262O79NwNqvKDnJXX9Q0azQC7MQwmv1
g9dQqIrpk1Svmo4kafrpcg0SMP4CM0QGEYZNKWcytOtIE2fu6q1sIQrKivNaT7ar
yX59R8k8M3wC1i423dOofYwAeFbG246CsfJnzKKZbhVCG71xk8iqtBKZkp74I0D5
8aQSumCMx6dtpufTqupOR6phQuPc2Hq6XACkm8B4IZSpKDyQo6kVJ6ul4388EdDH
Q87pIOsPgCLgTX7YFbXNksYaDoXHjc+7gDq/keZgJzkEqEHNog0Qflwsdn6njS0D
jUqFRNix9JgCMDTlOZnTKfwOoImNZxIFnPlWBul//dx9Mbp3vSnOCzImPTiBBpZC
aG6FJRHKje8Bzn5KZEKGr/XyumXVxXbmWFGH/WImztX1tTU3bw5ODrNvSyyJc3n5
tMgVxzOXjv12GqsF8ZeB6jN1J8J/r5t50MVNv3hDHg7cl6ir+J0clFKXztj7Kxuk
wBhgJa8khR4nPhFKxXrUphEKO6pQknTGjFyeTkQGOCaIdE/Vby+L1ZsF5YFi2uv/
HcBacDIleoh3uyJqZ/Q7elX3YXxno1hbniw7+Ph8aOWSRAMXzIyY1Rp/UadBfAfO
JvUNYkxNJTKykBzrDdkijskhJtUWOPi9CwbmOW6s8+PoGsZVdyNKG4JrP9/P1fCT
LO55AUFoJ5NHsxBakN7x1Ne09mu+rh7i3gMn0wH5V5dsDOIW0xvGVS9XJHYat4hd
QOz1NNqeJ6A5WKVCKsbr5ex91y0NzBL4ZbdFbfFLHcldufwORdMam3TfOyOApTAg
KtQUxPpbIyzoyrq4PT6RE3wvT3Y7HEhf+S4Vuv407snenCuqfJ/v76l/4YeHxssC
b9xtJ66laG5xBj+HqMvNWhPoV0uqiDXypRqt9chQ+qaMMjgLROkP56fkiz+z1AgD
UBegLIoXaNnxmnc+AlTh+qMQ4zHqNtJ2taQuHNbJVoZ02gxBWXSAu6hbdx9kmT6Z
LlLu47IenKgQZGqUYr7s+abqdFJ1SIXxc1SFQFjGjh1tuAFfB626MragEUSq/7K1
59GsJRdIYPlmHH+Cto3HvbDy3kQQGjbSu3bUwMFeX/IJpA4krvIBBvI6mU9mBcSW
75x7znINM0Ot2WQQ9Pzd/XvqVaD9RDKdpaGNS3xevJgcLMCrxMxPbe1S5EHTW9HK
Y9O90NfGXq4NX7Ts7+BMbKfBsnPESSwYiGQTDJLXXv+PphbQy9zC/cbZVmpVeGjy
qMrD549p5yUoUilKlRYdlcI9OeNDg2IeA7ejIaZzr6ua60sCUEqqXTgCHtGv3j3o
PeM/9Bf7wcvvf/xSQXBKFNqWnQbAIUA94PwOP2IHgnGFE3woorPocmKEVGqiZ6bW
RImYZXYcS+hjK8HrYFXcd9GonSiTNF3iZ06+mQEUKRBF3qJbDC5iz4njA4XN2Ik9
zjbRVtlNJMJJXwxF3t3xCE6So0ImzTPsjZtY6fYF85mRGT3HXicQqz6yN81olZ6V
lDNUoho+2un7hfrszr+ktkRtcSe7CnqtzfG2e1i63S15GJwWAx+/jEhSsURWQxgq
vAscmgJT4c94apQkAawaJQ5TuSpPRHN9ud9hxRCGKmNh7IrM+HimTaaKGrE519TO
helNK1bKv+aeaxS401DNUK2/u4269z9QiL/UQWiQPoZ11HVU/ecmwLHKqgKNe5aS
6OZ370KnMUtQbBW6gWCcW2ZLNxM5BsEblLxTRA5B0RW9iIgSBYpyT9NpAxZXoogK
FXLxPAaVoXns5AUBMfBLgPJxRzbOVwX9pc63vyD9iHkxTgRS1UNrGMEevTPb8FoF
KHwNgULd0rTCf8+grIrEeLX9969OusKUiGIDW72rkPQ75M6SoO8rxQ+fWgfWM82w
mwqXsM4vpLjUWZ7LNB4U5yhJFSQBQYiyg4xmwdogGLcytFalOEOg1Ki0Vkdi1PDf
Mx+2eK43q1zC035loYR1Rf0onX3SFUw7XljC+2BmtuyqQcicI7X8bJUfQiu8uHl8
rCrjmLul71vw1S8YSTntI8+PyGakH8Qpiju9ODkVQCpg/Hx1nJZlff3pC5QAa1jH
wEES3ikEtiC6zPg7lwRPF8vz6AISwYddjWfZR6kUe/OkRQzOqK7QUdoslD9n08Eu
PBx+0JmtQ1TfV92WxYoF0YerZFJdsj3DkSFsQGxFsJ00CdbyiK2wbeRktP5L22Rz
NDOg+IjzOatqoId+0wfVzLpooQu+JGkLgIzcfHHbUps+3peVHCZYiLipJ1uUw+0n
Y32qFufv5IVsFMPacVlQvpTGGdmVq5w9EDBLaxSWGnzd8uk4tIU/OSMsqQUqMv+T
aFJhNWSqpu3+OXfN7PbO1yU9V+ekGo9Z2ELr1IIPUlvlZWFtYTQJ3AVT6oK/R2lI
hpyW6JbEP2BCnpxMb9HmAn6YARc/8IuV9dcFs4HFIVOTVN+ec+dUhDS1lxtIMn5d
4+4btakcziUx1qKHk/3UVpjfyto2zybQ5t7ZQFpOga2AHj0HUvJ9E0/hIxrsc44r
MBMUnyhosC5cVbrgTTldXL4iaXxvcyseopyljUH0i7kz/vG14qmmzL+HhmDno1FL
l7sub748QVZ6qXlpYRXVhecUzqubW1e16mliYEjKwYv4kNVLP3MpWb6myeSOOkxg
KIJAueV8I38b8/xBT9ef8lTy8pn2/DTwVAUrLggN2eoGez0DIi8BkBhnGP7W4oOv
sX+o1b0/2BH3J/OqyvRDz/HQ3tIgxr7nKfMRfSmYJuDLsE+AwV4lVT8S2FdmbqSf
NSSgpx+4EG0lj1PxlGwEOhLTgwZsxPdIDVStUIGHNVTnzAELC9feaNFsYe4n53TC
jOKXwPPJN21EahrVHXyGz+kN/wMX2zPsMNXxx6ypmxkj3OAdjBm1tIzqv/quoObj
UpF63zpwmH3Q2k82b35Ta+o92UoSBqDFP+heV2PU3CwGf3Bnm7oKmaLW+2lc8Xi1
G/eXCacVDpRax5mMfE2obzrYnyELl2tQMZxvujGQRFZSqtXeYA+0PQRQcmw2Zo/m
2nOZ5vHUZaxeHtOERyvXRex4A9l2NNPfLGgVuo3zS0gIcixLbBNcjMNX7+OqVlgM
1hXu9OGg4kKDffwSiF6wjncRYdztrgpPe3Q0F8Qtkbz03+j7yQFX6CRPeF2FMbMo
rzLkPzG5xXs5jkRaH1oc4+BdXq+cwqRLR42gDKIYcPKKGxw0niyMqrh7K2UuGpv8
rHiRKgtNthhwrX+wdqPR+YclMFoC3994r/vDETAvaJfSrVPMGpKxJpqaIYnR972p
t+75xFCPmUCYIV6q9Aw8OtuHxBieW912AB1J0VLKcg+hJsHbYgUI/y5KkuJ3UTvB
ToCP1orDWWVNecH2+QJrBdojz9L7EOW8MuMxuhCgFu8IgIw3qubOLNzYAItfUcTa
OLbYrm98JGvUZytkF75JdhhHZqPGko4F22tLHpVXaOamCc1WinTHA1GoDmQG0bHT
NWgjm+qPvvZB/05BIDyAn3zFe4PBoCOIAP3obrjk/kbxGj0ueZzHbpMHkgHblIUk
waKKY1sToB8pdg0yGZu9bBZ3WPRT45z35R+smpqCW1p7xahe0MpPhQBVWgfapq7B
n4jxb7GSp1ElrDE4YBW8a5ChEhPXA5Bq5fuTqlwrIMW/HelYhACV5EFX1l4SdypN
ilwFaoPcYkFklQtdMQ8tfbrRZAz6zMV2T1FTte/BxB7TbtPq+i/YGgEeZUt7ylW0
SQPMcpCMNd5pnyOO/7Cz2arGsy+r0G/MFH990wDEP0ZsB0/1DA3S+2DO5jONENpO
NOH0GL9PSyed//V4p+pTWOcSu/b/26vrUD0jWWVmrZNUjX6tzWois8h17ZwoHPje
rLKCd9jQnLbaO5m97QnnRFTzoxNGTHJbGQLJO6txiy1YnfKNqgF4H0wafmNmFJLS
SusMfO56dVfTevwYlkeSiZYrGdTyBZUWyz27Wh0ryGCWq15eORl8kgFp0ouXWoOU
sZZO4rdeJMvPhv67id4VHbMtqXK8AmFKFGtuUEiUfWWJgH3WjoeDQM/ZLvw89oJx
WgR274UVulhdFUpbxGGosSaclWmPtm+xFUVUc1pJn8/VzCCLa+1+gZvziyMsiGGA
APb8KtC4yDSmfTqeKWY0qaeorLX6X/BT7mrtJFNYoWRxIuT0RU731mif0ZdQTAW/
wyUDVyMogS6niKtJ0mKv3NKoOc8zsziRGn3abl2ninruto+WKiVoLreMUbzrUDuC
/rDz+e4qA7tXcjC5djff9/nnyAy89JbfND5LgB9RNeDPBuuH50fRS0hT9UQltnXh
hWV2EtjlpNbuAFkGWI0OC1Dx+ogTuy/VJ4cIYiKqaY61fZSeqHAyCErV4ktcx20V
Q9AwaaG+5Lm/w7NC634rOLl1CGtDA70I6iGR8rXduCFtgDq0gYdCX1Djj+fioqWN
L8GxHIsSRjkZ9b+PK86maBbMjXp9OjxSFa7W2o5S0XIPveDG7lRo96A0L5BC+ico
29ci67B2tOpSfLuw49M/azWCpHlX3o7Ko3ru6GNaXqqQlLnvKBji6VHSirMXzgwW
1HHMVZRDKGZFR5DI9qlG6IvOsuj0/MBSGuiMAxK5KHMJtGmfySeuOJTzItfBDV7t
1pGGatVVhPGK7zBKx4A08wiruSLbfREiEv10nzVHOAcrwj76jlPaBkjGFFLiVVDF
4BS+UYTrtfo9vL7pApVNeT3EGRrNH3Wk+B+ZmKyhKLiGqt5ok9DqlY4vg5Aq9rdl
ZWONiJ9NJnV7pdz4q0RERtw6y2kweLvdtWS1bz+Q8zUB2z6+zhPxPuA4+vMUuJzD
XGiU9Jd2d6Q9J2bdGezCJhhEP3ANeQPxMP/jzsXpeA4vkjMYIspu4Z9zDpDNLTmS
hnzIrd2VokTUCh+eopHgJ+evGeP1svDWmPtSoKV+rxHBxaYfE5j+gvQrn0evp+0e
GH7ErsEGOmrf5UX2Q6+EymVMmspydz5BfqtW7AoPWI2a9MrZHk67bor8LFNfdztl
/tXVbMPLVFGrE9I9sIeCnYPxizhxcEul0hsfouG7XyVzX7Tn2SspiRx/Nd0mK1yd
FEa2CV5YpvqGKhuYA2mRvR92c69OXN75/AuPtE2EoEduP3JxlbnQGlYE+Yt1W6Ld
yWnnBc81R7P+3JFIxXTiur7znzfOqTze/QMPW8TiwogUTb0gT5+yj4FKOfN851bm
h4EVHbcpHvFW/KM6k4er3rc4uBs1yU2LzguobcX3iMfplZ06GFBQRlrZ6YVj8Ylo
KVGTjA8wnGTim/RKHzLSTjXvkcgz/5I68AzoVcH3cwUcmd/c9z+/rHuek41Okt7J
RVEEwMt521nKR3MeFQZysMRNOjNYTe76m1gaMjA+EPEsY0C9eexEI8Km92Zfxlk7
ZfAVuAu6gee9fz/toAkUNXjx38RMoQLJjuZ3vY4H4DfsZRA0sO+nTybzjmPG3P44
i1L+CD9No1+A/ImiNdJ/RxU8vgXJcMN2+Ea3rQw/LdU/RmmoEiieyUJzKm3a35+d
51J+aipP5j58Qj+KQ9mLIIaX0hEaa29khrnnGVip2df9qXyY4lev7T4rOg7xmwqJ
UdlbZYbtDHbNYlZd6VbTFNl5ZmFFW5uDIcSmxHQNDgXI8rFP6RorwdAdw9dKE1yp
BV8jMY21SVEyrptkuhtFJPM7hs1Dm4VWbN72GGDi6i78I1tFu9jQqOoF0ENPAACw
vD0zOjz0aSJPWGbOEHwW3j6IGy8RyMswFfbs2+H/2x/h8Mz1QmbClvPfN4xgHVev
9PQgXn0VTi6Y5FRRbdQrh+PH5Ni2ODEErCfiD8hwAWagu329Wj4lFw8bdyJLSguh
v/jugkXBJCWniPgk0GX02q4CRdAxMNO0ke4NTDjlnbH35AkGKtmtEO8m+xyQZv5+
wJ/oboRPGUcKA2VCuQQEEQraDw4p3zX0m53FdOtY3LDG3LkJACimzipyp/0GcZR2
/fXAxMHTMxswGwdlbPcE89nfi4820ioq6vFCxqlnGsNh5Wi+gu0qjDPBZc2Euvi1
pZVb3AnccDcnk72FsKOSIdqQgepc5M+Osm6BDf9FrlHUCcBWRTmQYUkqZYbziKDZ
+2cEzUcEGf6BwHNMT4mzUr+LC8gs4IsJlvJSFyec5g6LTKdxna96Cr1gQn/Z0BF/
Akcyi1sqLYf4aDO6Gt5RpA/xpVNTdD//r06k3l5tBkDUZn7VPa22+I1UzSHNKwQ1
K5HE94oDVEwYBzLS9WDEEZeZx6OYA0+f80g8imd6po4EvW8DpnWI9lufZFv0AoZ4
Lvaml9549Eg7jVQ3S4FX1Mv6FRMrFBDhMeX37vu9uDsMpZ9RJSgZOZQE/9ZLw3Os
n3CfHXdZKEUCvbGUE9TgKHRARL4u6E7rfC3jjesWtsnecuBqYONo+qdHEEAR3q6N
AYRklcn6ztYoiaE7x9Q6pSRpUFxJSreu7YM//kCJx3Gq08WfbublNkQDyvdZR/Kh
6wiHo5Zc0ZcRlhnbuYTDNSpOUBa7mBKkr/dEhuypgOUhXNpF0kSAaGIMaGMQNXxI
FrwfaV1R/QAdXa2TEf+tBV2yTw90TlvOWKP9GEZdfEvsfQ3Vn2uux91ZP5ylWt6B
8MBHyIDMCsRQEP6wF9Ry3VPPNMIYIsghIQJSbqw+Y8DWVNSulak+AIHIWIxVoLxX
myEoLq6TnxpqIYK64d7hThg5mRxxIOvfy6+fcggFAA2sfZoP914iLMc4DvKpcP8j
I/LpHcSomBbtgqhyTfWoSU2bEMJ3xLG6DTmQblCqyTpHEAF1DhEJk6HK0EE7BfE+
HW/vutzSQQJ9Ee35nZQ0IAOxYknyv3yW+Ai63Zhk2i6v8Sq+oOZEL/2V+LoKxM7N
sR6cXGvLUmJbjhvVzmTyw7i5fd/FigySyFUD8KzxUiPAIZL3hESC0l26T05B/JrR
nRK5rj2CX+FjInSMcHmKoDnLO9TW7To+PtU5SneUhXZR4fcy4XkSaN7ZhX/nuadM
FtY+ZB7FQ8oZ3so8kFyqHHk8TVu5w7tYi684Q6WMXoEXB3EwISW6tnmGrtQv55Ya
3f40Sta+E92qbexVNkMJ5FGqk/64xfCBtcTZpWkT0rgQ7fSVb34NyCwbA1Mj6F1L
K3fYHtZ0a9Oy9nHy3+dShUU6Bi0D/ve+suXnJYj0dGIFCvvYcGQpgznW1iqad7o0
+TOEQmQA3lk9dzMBtQRaVqKTC3ZRcQvGISkaNwiiYWKwbqi8rWPQA22N5yFQlRwG
fLvpe4TrGYPj3a0XRTDtKkVOXs0Z4Pe3E1ckNLx3XsoyvYM+2EgzRKFDyWC1twUn
ZkARpSzdel9o+lHeBs8idoGOkDlfNUkoHpRnZaIj61pyG5O2DPRFAgs2+4JPg7wo
Qwva6vOsoScak9oHLCZntPm8xtwpT1QcgJvFqjyklxV+zoKxk9zxmh/yGw9FK2NL
CHNWl7rFCZKMG3K9hQoabq7psW0FlTmbwoYU4bHmo54ApvK7NPlWYSxCMM3ndBj5
Y1xXwzUmkH1iOKytXILb5k6QEhFTGraJEJpNO2K3kYuZ4LmQ//txL+L7/L4y0nFi
GsWOupe0DK2qxS9wi6pXbrrWgDCi60hSxuWJyn21hWs7EaM9zwwbwjVvVPB2VJNP
YyUjQJr/dQ178334AL6x05Q//hnfT1vxmCaMFABdQHaLOsiWJR2XD9flxZBKjeAM
FekQrVrt2EZKJe0bXwTdXH36/gUE4EyZs2PHdeHAPhVOp3lqe1tEZ2hYiaVD6SSz
uVoIU/o2Rf9UeDbFsGEV58BrMzEbJb3Ly5i+EN9TGkEwHSXErpazxsKygU/KCepj
ZWAhV8oN1UN/OyMNyKGD+4tR96dCUq7sXGc61NqUmCYu/rX72OgcyLhOgIVoJtxJ
9gbGJnTDu+rkL4iJoMrHpYaSIWrgic4euQB6SM4ALXjzJglPEVAtueRnNJz7IIs0
W7s8GTv+eKa93POB2ZoRpPdQLgYk+RWpUzY6ZznGuQ0aF/ypbJzUPy5WVRGwghnY
Cd2dARDdsIqrw9I1T+a49FGaYTa8dJSsW6IWL32AxzTdkoLz3qNGXyEAwCa3abqh
JocsGp0k9ORy3I+boQcGgv2Bzt4GJJGlXTjfp56GSEh8H5NIlj+A0FJMrMzRbt2/
NzQAB5uEMEYnprAYbHLwRDGEo33FdgzvMHavmZczyGcvRuqkO/H/J6rdqUk88yrw
hT2SXjDt86ovG2jdgW80oTgWAkQQVLNaSSASUlEA9nNp3+zZrX/5BvHfN9gp/J0c
oDrdIJPDNSee8sQ8H3c0WbxHHqYlPsLU7pV/9mLTIv/LIEJpcSUFqRhXfiQ/kiXJ
F1awvctWvKR6Wj0cPigHvr4pXbPav2HUcn2n87c5NZNDk7kUjoflosSUnAnKXmNK
/x1LVzUZKis49ZMfL+Gj+oYaQTf/trkp+A6cBMpD9qm05SQZ9/k9mbrhlu0p0qP0
AQwuPONQnrymgN0S64gVyyuFlPEuOk/D6VUv7bFOa4pr57+Nimru6FirLPK19rO1
8srFRzC86RzqEAS+YqA2q0FymL4dQnwLEVO4AzW30wgMUrQzUoR9QXgHOMyo2/X6
OBybfP4OqaSdgqgSFS68huVJxtU4CilEroeXcWFOE+c5dKXse4LDw8DGk5s/ceJh
gzqkGoq9j/tBmI+NLb+OIasPWs33z64KQMO+Qy9rGIr31KxsjYJnk0WB7bnfxem8
oHLtGrbFxgMnJGxOhsb9op9GzWh5tGe+iuFb4F+eC8Rx9aAeBMGIIJjkC5AUQMx9
xeDHfA3aIiPAvE4HN7Ot4G9ecn/+EoiQcEeF0IuD5A7tObQk4m23FRzzslreut6R
HbSbHvCD2g3fD3e+UQ0oegdUTUAjbYpMqt5168cRhhvSH/iV+nXrYnApqp0QhEXH
z4nlEKzh7grRUKf/qJ4nwYnuOQ9K9jlf7jfvF3AMtsopfznt7vZp1/IufNOhV3tW
owwvtiidnbpX2beRyS3uiZAXutdWeAR2ViQhudaJ7t9Lbjq1wl9WUBvZN6L2HEdQ
DCcsRfVJ2XaY6LsPgI2skEdcWElKYP0fQ2wwr1G/3QzvY8KtCr6Jw4mCZG4EG7YZ
x3L7rZx65XFZEoddYF8CIX2npPEYi26jvshOTIjbgOkNO4kLjRaOjAeoVqOB7IXY
ZX1weu1UuxOOG/DDyw7Lm/Wq52Vl2D67vWIjQDC4iqmM50a1bXWg9XAJDYjE8GdR
rM/U/o2MsHHI4da0nfudl2D0EaMSNva3F8+hIum+dQARAdbtYt0upStppI8i6qZo
IvNRAYLmZ3WMxVSpBOQoobkjMcvAAuol+BQMpyZ0XQXesmT1RsTNu518lleL6osa
yVoeAKsR2oRP6zil59iFF8ppn2CIigYBd2A12oZaueYR/qOMTqSnd8rHsGxVT3Q3
WO33S6sKnn1OPBxtozR7WrKsZM3De8BFwsYUYRbVfd4sRdzuc8nIqstgsFglvMii
VOmTBhglIbQ7f/5B/IxenKd4rbS38lY70yFzvsr4JGFjU4/30h2x+OwuU1Os2Vx4
Ol2n85OSNVXv/bkK7eaSUZaTgnOINiQ/Y6B/N8mdK9ZR6xkLnW5a+6gUTqK9Gcgu
r7XQJk1OteQ7OiU5clEe3A4uqtReoGvJAW7s8E0Ba4ZaoZoEHxdVdCou3vYUVIvb
S66/SSDw0Ztg8TzZio5L0wZpDjg9RxD8GGwYBYQuxN5Jzql5MJPNHQG99r5Ek3f4
lFYLYMVMxI1l/vFPHGzrfXQ+Jy47ynVEkjLjqCpo7KNrOqenHy8RgNnwGc96Vo8N
tvZ4pDpv30kfu6QemFLGHPpxieUfQelht7+qWJj1tQcfQUhF7e+jEhTkeB1BNqRU
LZRqFmGHLZAG9aaI9uwDzrtr0+Jr7KwDJlK1sroBIM5lWkhKGo+lUuWyJ4Jw9zJk
UQuYztef6lvI7mJQgneidVamocnxI/ZEjcSOPvHJ7QFXX7+wwxTFaPSgchsw3DE+
dZkzvfuGT6872MvqhH9b0DqAcoIPs8oNoZnoziOtsugJOsd+qVleIOOt6kLQGor1
TVpQ2RcEwv/5pRC7kyEux7dxHMUkulbeeZpzsZ3+PJRyL8x6tYpL5vi3e4ZM8YlH
4aOrZcIMcPYoaPgg89aKVmFkaY/9RnLDCruocmmvTNjUQrK9abVQbiw1NgtlLFqY
4aRePBjLCQthtrgtecV/W2/yNSt7jVNSfVYxyEGTS9XVhCR5/cT2UqB/l6AXssyQ
6fea38/jK6q9IWs4Kx4ZHRuD2HBO924lgF06ZxfI7QQBiBySUmkHvjM+hXCuT+z8
erSWNkyTO7n3fRIZDb0B5L8v5DXmxgx+AxK+4eXNAHHLgQ4shEeU16waL2RMYBIh
G1UadKjq6dnF6ZL8iCyumSIS6PXTbN9d61Et9TGIMco0oiqTihy5RRVJ0zL1zQMt
kJYTKmVA70rdXR2VzxOsfeKv0grtmg0jsYvyr8rhdds3O8Pe2qW9EzmoQiV0Mctp
pAYcBTJDaquTkNIcqzKsyb/0/CU/H02sNvhmo5PLxrE6CzL2z+ifxN4sUSXUoKbh
EOdCZCeFGHMWF9mgfaJ4ITrpZ82MYJBTje2RoHi5u5VB03VSojFal2o82DspM77R
+WRSitPK6ba/MrEzgoo82G70kEDwItZB/kW618eOgcCWbMTa/t5aNVoNKk0Dn/GL
GMUCsubbr/0EV3qHV/wUo3lHMkvvWtCEvYeT+YQ6M1H0VKTsk94mPmx2KwNejgBk
3f1wrDhEwTtGz7wQQwh7WVk+nsl+b/fkY90nIsh1GQTZL+NmKAxB2AQ2do0Xk1Lw
mmYyUgvDT0S7v4A24NHzx0nEGX300OGoF4bbavDpQPECU52JHD8LL4w/RtwRR2j3
Z6h0S21o8VlQ0CAA7OBkkMgm2cwJMCUnMbj00LLqMbM7fz7/RASD6ye2OG2sRi7n
wV3hPJqeM+Z/hVqy+S0M9wWKpNqVm/I8s+ze4hBmyUTDlxkcSaEiKkgIB+PtiLgw
mgDsI6COiAFs4z5xnuKTmUZT6X582T9IBz2T7JJjYZolOYwSeT8Qm2P3h6U5qGD6
l6n9e0nqrvffs2mmFlGclxDmuBiPwWkD1ozZX1uPxLQ1mD3GQlHjApu6NxrP5sIp
yrbKl3NjIeskke/gmw+q1WKg/29xMS57TPjoJZUUoc+iDovFj6dLFfn+fFQRr8Ik
dJ+YWH8RTeLciTS6yUyjQ17f++qdCcEadSARIrf2Uw4tMzNBLIoD7z9na34iP0EM
aW5LTjVupbETUQlfgtCWPPbdmZeKt+5FE5AHk0pyFqfQPXgEdOulNsH0ZeLkYZOJ
ZDZpEIpWUBQfQZC+vktzZdwg7NLJPOeRRqAHJT0pkGaTtosZ1nGVdhsg1+Bxo7Oe
tZJAo5H0P+Mz0TCJw/3/jaR7c0PtFu2pJ+04QIkqcMsoYRb/sOA0WrJ9Ykf7pKQp
qans6n4I8dwRjl1VtS/uUfu2g23J/OEeiyW7TcL6k6XgYwk/fhEVVEkFelq5sqc/
JSoEs0nWUKr76+0UK3hO7CCXRcFOia9PcyKdYNJtKLlcrkhkpY7/s7lHOKJXBlLS
7tNFJQa2Ay9IFjUCXX0Zsv7SAA75125G+cjQm+bQCZ1ym8J7eJZxaJSiWz3QM4HN
BRslmFxHQ+mtHZ8zNZAfxQh5rZs///PI8XsKA3TJPMTsxa+wP6nxsG7GC269F+4z
YhbgultBJXjtRSoEy6YZJSuMVk6f8yBr2pUdfWn66TAH7IYbJtQbrpfi2Oc0tQVP
4q20uvQ8nlA5OEKBEHRhvPx5m8mds6oJh/3Md/IhoWsdbFLTTUC/ApzIvjDxA4za
8pG1HCwRozP2wxxJsfGd/K91ue3Uazc2Vz9btIW5zeFVMQqRCM7g3poxNZc5dwfZ
cIPtjB/owtH0FSruUrMEVQ4oSgBKWbuvw4fpgWqz+gFUx3hs61yd5ljfW33nuG54
AVjCWLwDjoifvk4Guy+soZEWbGLFcJNKXOoXzoCurcXnpdlUuUaRmJ7sEB1kLinM
lfX8UtebvxmSCsslBB0siV1oMWeYpzG/PvMW2lubLe6b30PRQqHXBTIpW/WF1Ym7
bVn5kOyZNP4V1qtyEirHsnZUOXxjs/5PSiTdKe4PVKNeYvCsg84VyJDq2QM9v6Bv
i+niskl6VZNk/DbTHod19GHHJAxuGDJWlht+Tb9ayhoPy0MwySWO5m8/ejVTWp/i
sveJG5h4/VLhmdiQHiwPJCceV/9s+n8OkvOGByCbC1DCL8C3OOqP+QYDVESBTxHB
EW1CYtiAUC5VvqRGyzOEpsbLfN9LgEgu/tmE4SrzGC8I+WkNRM5MdrX2ywNGBf87
dcLALETrm4wemTOlfgajnhpH8avuKlHBYdwffepmNhhSGCoITzg/WETiXFQtMHPa
T7KhdDTpc72YdBBrLqIoliWxkv9BHHRXrY038AQr7nUEOiVGRIs6ZHYI+QUcKGR1
+klIdMFJhpYVowWUS8K6g340+nGP/cRXTJO04MLo6w2NjdAs5LIw5kHTQKNFjV+H
7PK4KI7nOOYlwAKW/Wv327Od9inM4R9b8u5vRpWQ46ZPSXtH4H8giPnKHtm3uuzG
0VQq1CqIC8S+cZvE6svgYgRJF7BJ9AFt+eA9NNHc9FGHwt/7RuXwMXG60ElRaGXX
x3MrLBERnXvIJxe0gyC6lH66gq+JrX3e0PGlcO7xObmaGLRwz1jsQ/eWnDh8wwdt
sQ4T3zDdJMaqisjI9BgdUL4jLqwMZbuFN3P7vGr9AB9dehKTNJQ/OhVTuQd0lLgA
I91L/ShWNA4FxAuL+yLdvZP2uSpU8M3gpmuP0OYMGSKbPPuTqm+M3ZPZET9902YR
8YW9XXcBAiB7X4KEiYjkrRe7o7pN8t6j1R3uC/BoqBP9mhhy3SSw6X4rHXUTzrs5
EaraUTR46nCmhI0Xp3r6FAgGKaPlCehcH19jEXuNZq/11pxyKAX6ebaWGgNCvNse
LPDmzrA55QlSdclEU7TUbtg+5jK+SJMxS7TIzjGedCpM9+c3Yo0bccNfGeE0DGN+
3Q9Ey/xrRFjnpSra09Bwo+lEDjGgqyk97L/l18Mf1IJYuahraoHbHdkSPQ7cL2yy
RPelpR3bPb2vwgjLQmLBA/dJeO7cUxnmpOfHfn4vfigETrrZKqzzhd6KpZcPfmLO
bGk4bhccFEVrRqDJHH+Kl4wllGYTAKvwzaVPCFLve6YJSpPJwWAlX5kJys+NqXSA
CEaNeuGryoVakLYL2YBLCsAtQcueQJHxMopm1hsxmO9FbIxuSGvB1hfgIO9nBgBM
0U6QtK1Sgdpev1+M8l8VOPIUCV1NyrXCyIp9qv23sjB0si+U2nFUGZfK2xcXxPsB
dB7eQoJdzJVsHRWXidkaea4xLE/yGNr4r/ICbmyV2XQqdz0Pgefd82E2DSjzEnjm
HLoSn6NT1DSS8RmfMFUxNsHK54EHij/SOlgl03CxQA8skdxmFUTmOEuzNcak59R9
9lN4vX5b71W12Ek+7od1OJobjtApzCOrgFQlp8VA/mj429Wh23F5j5GBd++m8J4A
RbJiULQ8KpkPTZq8ouyTZxoJVbP0uRYhdvKt2KyMbyNzFtmxju1IZkJ4rDigUdS1
9wtsM15QQDlNbz43AVS/43t5YqwrEwy20UOIQcKwZyXoTmuT/4P+Rb/nNnhO1Eep
qHEtwyvjDWJMJLn/KIM0a03XrRyyezgpyU/gbKqUkO6O+p/8LyUud0U7srRi1kTL
dJ21iiB0EqJC21IVzSwMvb+coEJQu2MmY5JSN5tlcvyMkTvbJbF4DRwXCaWW9Plu
gNqQs0HQYfJ6nMcWXXhzeL6epNYZ+J/aq78IoTexiISGLBcudcsQq0B6VmwZZZVZ
q/nXDSnQIZOKpR2ANhwcRWBjhC9boEwksJjjxHK59cUucccQbV55Pu6II6K2nLz2
556cWFSeUvr8Nib6j+FhXyJpMTpFl9lkmdF6gFyGvmXLcCYAMsHBmWO924YS8Pz2
5Mf4gO5tx4GfCsNdTSGKl+kcf2FL/7HCMNxoKC51eBhZq5HG+3qUH6FgJk1rktfr
FFU3ug78Efti7I7rO4CZzRVsvXSLTCZpqCzrTgDZQMcO64/3KmpDWTbjDmrtlQCt
W3LPqvIa/Yx5kZXTqiSvTp6TjoeOnmvdNGHnaFj4uQuR3edlXRLbLu0hmEg1+w9L
I2tYDuCMXIEoL3ZRPCYbSzvz0Pf11bASh6Tckhq1QFzpipODAisJ27S7/EayspVh
2rvwgm1Uo08G8BrWzCA3ZxFyXgliDD/5mZaXfidSYirA/dMD4/u9rVHxsIIEPk5/
8HWxDdujdxWkRnuxwBzK4r9T3gCslkBC3JcCvVAjgkHentwg9CbDc7FwX9OysqMm
/HGd595JJ4/htJgjChymqRzhkRXhc9bkxRseBYtyRJpLL4uyxSwJVqG3PIXI0A9r
XON5dU+D+M4FLdd+9n1WGljRMZvX3BsTIRL335EWR7HyNQJ69eEEDm15P4woxJz7
Y2uf9Vuf8kAfuEbFxAZlFYYWBpXmb48W2cBaxIOkKBD1lbL69q6MgC973y14TjBp
x8gjKA8fqyRU3JXE9qJFf4esS9StoMEJ5hZaKDZdrTkHNJ8l/KDY05g1Xnhk7Dcx
AnaKLa0P+FlLQoeeozTdXt4eamgotdZCMSNcSfs8AQrZzYDO5iph2LcRWDrW4GMY
Uc59RkToQUGfA4lJbK27uqNgnI+VM/MijU0410Tx5rnN4gaGvs2NDSBRJ4kKjgDB
GWofimVJ8KTdp8TvZMpLq6vmsXozXp5WHevTr5F0KaJXgAy3SPFhevjCiN20OFQR
ujC1ornYqjLIXLGIT8Ycf+FLvrBCkSD3Pmdg9ZeMayYjcAZvui6PFQH3HFuGW96d
YFNd8a6YgYIdrJDMqonrCDQO2cOWYGvu3ozl9WhxpWU4zD4EpYRPd0XAaWwhfUOs
+r+N0sujHL2OYAG/C9Svas1+RVTkScC+vGsDjC7IUc81c2bQWy2W1B9tyzZryLcj
EAho3gZ3umpRgCJlXKCSi38aNNhED42tRmxS/UHSUsePijUbJU+Lq8hD6e4S+g50
qP+9RH36HueTfBMWkWW8SjqA77giD36G+J9atsVs+weakWpsKUD7dkoE2yHqYj/G
kWAXcW+g7g8HbQWHbkErkxqd56ke/dBpCvdOkvwVIoY4oTliX/HXG7KCI2YnRsGj
9BqCbZfJfph12wYajI+GaTXNbPrq/CCb+LTdmIdJSfoUXU+ojJNOE4ThP52mOGxz
XX7vfD21pWyXb6pD5p7VhZBlyO332tkHi/IdRJ+OOyW0D8YpnR1CWXQXzvLJeltT
a6GMu7PohM3ZTVtzzNEia97quY7syrRGikcRsPZSras/W5CUsen0skde56jxQ8eE
f9dUGeeogcFYiSDeMUCURwm4m2S3cRGVaYB2CQmZUr0wL9IGk3PCy1/Y0k1ukEnE
0DNPjk3d6OzNgaaxKmQwplLHQdZ9K0KbG12RJflAEok2DLPsbrKRESIeGQl90jKn
VgYDmRlFg4SL5eAomGO4RoqDeEyhEqTJDpT8xFS3iC9ApNnllqCH7sth4rsFojxm
vFV2NbXBGlDqLT7Vgm1Z40y0xwnoLw8G9wDmXGp+CcwV+PvWbTvEyBPDrc9sqye5
r6TABrXh1BO0qnlmARGMMX7N+ZpDRiC6xp7mFrtMkUUMacB2Qj7psPA/ipdfNOzZ
AImueZARu6sy+3gvxACvoQp4HigaEAsTuYZP5dL0M5S29eMKrq5rCfwbq+Ug10jK
3pCP8PZ+bq5MvxXQ5rLQLdchgrr6BZF5rR9xo6D7bMyyM81R+s7Vf+xzR5wqKKWk
uDq8PeVLUevpyo8KXiCqaxKr0tgfaBKiJGjQzGwok8cY/e/FQVY0c1CLit1gzjm4
hSoMG37LNwgEBmJJzcR6aHDJzYxK6VR6nzcgzp0mUslLQpGTrF8F2sGbhlfgYq3n
Snb8iSQ2w0wvwUGiDoBSBVhc6olY7kTGSzesAR/28palvNW4htJAGteZSOZXwgvS
olgVrLKPc7m30Oa/wKDOhLuKykU9FNXCaz4bXnEonrCtSTyz7njxmDUv4Q2UZRnN
G8/Z9hwThbKX2g+fsxnR2MGLY6ufmnkvsnydab9Rka1IXvaBcHWmt13mQM3JV3cx
Dulki7fSVsg4afv3hS97YetPBF48ftscR3RH+09G/EjqBAWVC/S8EFxPsN+PC946
EmxG5j1kJ+BdVoEm0kJhn4sD7np9eWlFOKm9FDmJ09mP2o+/xsBEldKiJUt/npiF
mdynU8dgdBNSbrPB90JqhKRSh+4mxUtq80EbhZPRIiaxC2VimQaKyGVxz0QBy3cH
IjyoaznYOpyQ2M/HWHY5H4F6zzYa8PVeJ5uA0+ZocYOUHy0CUaV9RjfzzS6ubmUJ
4fjFKw/pzCJb22NFWlgrsaedmaji06ujQpmiNx5jenH4hS7SrLKII77pRCMZoDow
YkokouSH1C87s7OouHKg3++zp4g055NtbfQoR+mcQ7SV8D4c69jBJpKxBS28COF3
cWZF4xMQLZiUgjccbT7g6SI2xxkQwhCN3S8Xp+HRCv0wrQJi4gKqIKKFE07tUBkp
S95TCfW2NlVApLzzERuLro0JZJCRhPA1zAtDRqB0i39qZbXb+PzMaFxFk+7pyzic
NPFrbIpl20EHZubIM42tAIDGl3NdU9hGVUw8/EfaqNJsdYw19jcJLH2+PODQp68h
aDqMsma3nNuBmQlmIHjE2mu05w9BvOgKfPKktyCuSeR8N61Tkm6nDkJYAiXSOnsj
HjV/WZ9tIJtUMErb3aIbhInrEtLbG6RRJaTYU+eu3OaJzn0tWpB/ILLaHlgE4CXi
J83XKoLMctm7QMAzXDzqj2mmHGIoOsPNK/0WMUWWcXue9FH1QXu2yriloRNhtpx3
lH7zS/K1LOeArtaphpamv/u5kVH2sJ/91vcmxaTAthk3cyIo5iwWu5kwaCmT1jgJ
ZxliFHXOIhiZzRRTVnPaqrobiAoWZF1VA5m95nU+pwt25ZYXkOaXAkqzwhwGwhnl
IRrJSTz1c8Ye21IC7wcPzRkLh17qG2lo96i5OfM9nMegwWmgu//+liYTKwCmjJLK
GSOF62wKxcNdXaqPsLTdg88IGqBTrtgGS3YvywqGAXpVXTqb4g4HKSBAHzvh+Alt
8qpuxIOy3z2rVXQO3p5abQe9eHrYF1NA5R7+qndkmQSFAFwRlTEAr7JKBaMSvgBH
W8LAJ9Ve0LQXUcS0ZcZR9zxHUUU6yBNMkV/ZVkpam9t73Uvr0KG9Zaaz+TnawAhx
mS7JLphsictqGxokoIavoV8XP+fERILg95lpA5/OIIKaGN/PYfKqThtDj6yKfGVN
z9Al5zNPaBiuJYNpQrMyoFBlJp2+3WNuBMONaakypWjWe8r4ldrezMcRJu/WH13I
1x+cVffrJNLv2CoIQcDTjtv2neoyybmOUa1XzUV60123P1P3rMoUAmp0q97wXpjp
7O/ywFo0e8YwEItdmDHtnyVkEHmdCh8Vm+Gke7R9eTkyIQBdo+EO7i5Sd+Wwjezy
Gf3BK07sPAAuWFYoHDvBfNuGrHZ0W6rHHMoZU5pgF4QneyDP41wlAJNoH+/rXs/n
wfMPBqbstMxXLNs0lwoLHNxMIifWCpLH7ArbhcXFZRN7h+JJLCMUwXGcRn5TqZ+a
gn0uGDGID3Vd6JzmsfEfgmjO/O/H+e9ozh33TDs3Hj7M4zB30sC0k1v0wCAarMir
XQjJoNVu3sx47Sn7VO86Gors8uOKhYxehqnmjAeZUK3CTv5wWXCN1XCUcSlUoQiI
zSULFviy1onIXCIwhtizg/4ecZYIZbwA6u+kw7E5cO8IHDHftIaC/sby/ald84VK
LyCnCcCDokfL0HyGSJ6cuZRNlXlHn2PIabppnDGEwQpIacn74mby9BxSFmVY5Wb/
l7obZ3m2HQABQJFUCTBPktrny5gM1lk5wR4EC78Rynb6yH5Ll2PJ3pZV0xXnOdXZ
K580Svb/x8PHAURNzcmk9X9q6GGHGrTXIGajSMjUi85gheKksut39PGqyBH32/qy
4nFS4dKeUb1N4GbhgSzPXJqGzTs2AMO0k/duRLmpacUkhbQvNL3l7d0EKWHqq7D1
BYWlTw9BNsqNdhpJ1EhV2xxqN+cMhPeBuLSM5vGLsAr88qHmtMFdtzX0shSFN6D0
ejr6DABebMHo2M1w5073Vbmk/bXlH0TPATbTCi/Zz6hIIG3Nqdh3RmSYWqG2jUBS
5KeQeOf+1JUSKZAn93xMPHkIRk2BbxuxdfDRMP3LM9L9zcZuP5vB/8IZf/3/gehp
bZ9yhqG98mDrpMl067oPEkHWWM88C90c/mjR/1shKogiEhjmxzs/Yb2E1FomjXpH
rZUTSaGhssM+QGbnpytySL5UAs5r8Hrb0kGUBTPf+k8Kdk9xvVFDWe6j3cyiF4ym
WWhA6wIQz/WSal86evPXEdrJBCvomNi9KZFMwTkdK0Dl73o608bJC/nL/pGkYK2G
Q9KG5oTLK4ZNdixVbmH0eZnKn+g8vipgXeh0nytaPn6jkWn8XxX7MwoUrMnMYUEv
QShchRSA2Zig8RJZyX0F1nHbOenlvNlW+jFfjFKcVJlimMibIKmr2MqQN9iBQxZB
+/lDYZHKvETGkH+qCFflpcw0a1mmgWnusdztxCza4CFWBA05XRRr4GS26gCgakwP
VvyI3q1RAlJkWSGzkT8bkwbCGWJ60Mqn0ndXih5VrMh6kqSCvM6bhPGSLKUQHoG4
Ceafvow2/LNoPR6sOuoiBNtzAfkdNKzhkRS9SKewBzWxUXsUbn2Wmj6aRQT9+bOo
pn4V5d2suNxRtMV3G6/WzCmt8636/dFhJaJi2dBiQryyZK1cOQ9eMwxOuli1Hk9M
ttOt6HgkSuvIvqSfOBUQ8hbnPCKUaCm/9mZRkSrF7kx0pMGhHYM3PXhgAGvG+Ihc
zKXX+gcOCtRqHRZNkS1V00TiN4pnsDXNh65Jtjh+YxPLEz8QSvURt0N0/4HeyhWg
J3DwNJgD1cXXItkvdkrsnpDUbSMCF+o2gGzg9B7eLGrILUlDN01e2wDd0CdkM7In
/bGMrSQaw+KOY9Xr1sf2ScCpXMVme7aB88Loyak2CwJpPYG3tD+gZnozZaFjZx+1
WMkK9V/axIRICavbYMcuQ5QcpDe144DfNsgVDYWRw4KSL5QqeJ6Wu8eqQY6O2Sjy
LdGYSXJegmrcaTvJWHAk/FX/z4sr+5JdL8RmIg4VnuTEXcOcmf26Yjw7yXS9YX4d
pTwKtnuRi4rprwq3AXHHKLkdtNP33q+jG1w7P27vgQO7hw0jrWE5ZlxMVojOwfa8
ww8reV3fnIwcg6Tr/QIvVCjgXEZ9Z07gUHX52iF4DRtgEAoAQnJBz9MHOT/+Foui
U5Cc0P8V6LIkRk/iqrhM83wYQNzKLXmTlCanEUhMl4sjBkU3wVWjGlVwg8N8+rIP
asnM20tcQiVoIgaxstMxOaFoya+IQTvpKfqwRx8QSbIM/wwb6oBUPo4eaGQeSsI8
EBJPPp1ut0PT+k2xj5ZMjQPIxNVU81cLsKD6i5PRSZ8dEekZT+4GuFE8cq94Cy1n
0H1NiN2r3fnmowPQ7cwBfVoPqKJHttsS8R4bp8XR6InTR5o/BZ0nSMASSFFF3+QR
2+5IzDRx2GzsCletxDDz3bfobTn6Gu7A15a9xdGrCeDjAJ0ypmlbKQn69Sird/v+
AUjJEJPc+z7WsWFdryFw5GXq9x7t7nayHuj40cqanWT0ehJjShuhIaY6Ai+aH3vT
PGYcym0xTCJAs/lrlsvIYjMbVwQSz5SWvkPv7EC8OWKh+DBdVqACKUz6xnvdyRdp
aWk/cHPL8AGshslj00duZEDLk/1u6kGc4sSIH12X55mRv8HYsrnJdNFbbKj5eS9d
sBf7sZSDCJCNcCpho0x+EScPsUzJm6RDJ/e1tgFayJbzqyIU6JCH3unUgJdYuoNZ
FR+hT/V4f1S9hdQ6+zIJk0KKwBdnwpTHP0BrdiQBUp66oAiJeki1gJFwJ7dCWrmS
SKnpQnxdZY9ds91/UNTY1OfchmaXJJTzX3ZIv7lx9lInXib1bou7BtKyxYYKwjIO
M7MEJyCuAHoSCAIX76aO38hZ1rjFzEwtnbjwM63krIGUwA05LWk7Qvp4QeBkzVSW
gz+1IPks1QEabNjU/kS8P9cZQsNnKfBCjzTTpMp4JoXYGGL1/Y1NWwqTN8lO/GC1
bHoLBFvbaVtxFGa1Qg+mZvnUm36Wudcr6WY7XsVM/JqaL8fkKARpEOl0okFHK0Yk
HqAqf7XcBY6zj35/j+7NDG5mo1b11hkmfCImlutGWsqDtTC6yQz51i+XO4HEWCg+
7AgmmiKWZIRXf4NWvnSKecn3V2uXcsOl0aLatubX3GisiUi78P9cyKrqmmorNPZy
ckqAuMpa1qG8o/vUP4seaCEkoo3/0/07nbGyeXk7KJYOCw0vLZaJfwsXMYinWayQ
E2P4gjYLgiUshgGOFePtZkm4YMXUFWMywQ2wWi5XsNFfaJbbqVLHvf5YVYYqPRvO
6KneYmH9s8hNJnxR6Eyc/NdqLqSf3zOJyI/1/MA5TpFQOGedDNh2oWkDq0jkRlZE
np1jjWc7pMGUTArdxA7wJf4YaYppgfN0OGM6zHWUVIJ8eegwFl0teTVSLAsIe4f8
0b/b+DmYWibMbLZNKGCMhODJvA7VsPNhWNZqsmAMmax19OcYpb9ZzIyMpvjs22um
YDB/nbusFbjeEgYvTPUhUbv7zstuhLTbiJOGh/gQA1brN2NkcEWsMjHDmGTffRg3
nIiV4X+CLKyr6GEzNCneaVuHT+Mepf9oxR71WdyfSDuZiwARdpVdFHBtOFc0GLcd
lqo6kwHgTIf0CvpCzuc05GObfzHSBH08la9d7Ke6RkH2DUeyzcAzvsa9wUeUZDo6
S+BM5rRUNUsneWErFzVsuIxht8J8IYqt472Cs6WTzFFmEnrxKQCfY7dmSMB+/o3m
KG+W9hTjakwMlmIuRuV6+Ym9+lU3yUC4o8o/yN8ODvb5EQWrObxRtKFNGM3TJRcw
AchkibwqRDO04aFd7f0laIiXNxAuyZqjAJqw9El9ISRLf5GJWYkIRaCMJChLrsnN
9i8gAiBMlAFDUhuvkxanixkDuEvvYUHLLyi9cGoTLwE8JmrvGDQk0DUVzPACLpz0
rFyiUbxkXqhiiVWQjzZkU2mT5owxTgg1hDB3xZEy+EHKCS37p0m+8LZooVWEvZ/V
C4kr70KuUeA8EpQK+ErIcNm5tVl47XzzbwB2eAzS0KzDw8LVaXe099B01rB/hqo8
9dTgcKyiMkWw8fY+iTbbZbSo6vn201qOZkO6ebuhc9O7kWf6vXkjoVtoIKs3bAH2
qhWLWyd2uz0PFmj7nlIWcSY1ooKR4SbRuDCBhJTm2VRzST1OdkTVTLA1pPOgdMT3
H0qBR1PgzwPi2iIIxi4YFJ2QTh3sxFGlvb67hGgMVv5wRvJp+iIsucNFvBZCGd/8
6ZK3wZZZiab541OFdMMl0vOG4cSecCDL0RntDDeLWoi83S6VDVKCjia0cN4RIlSH
bgCaDQtgjifKcjvrv5wZriXGiYR/CGyuz2B25LoUzTH7amWdy5o/IcBOfWyTa/wn
dKl8VhYm4mXe+dsWA85MLwcVA93AZ5M7XWzSwjQPA6i4l2hN6w83tVGnnqQfp0R+
oZLElcHX9IcCdYJnMSAvIe9J/Rae5h2EewdNaepun5tNOPE3JdSyOxeGu7N8AZ4C
RSY28Dm4d/n8abW7Ng4VbIwnDK0NOBCOfNDijC7rE+K2KncP4mS/25Yk9wlZp32U
7UCyj86kIzef57Gx7dA2F5EEGs4QpNrXkobE4rSD99Cm9+Hk0d4VYw04LS4f4Y+t
aNZ61hUfTQ0vGFyUx8+B4W1dh/otyuf/vNlCYnZZ8//b8K5A54cqYp2Q/B3K0sNQ
yyUe6yVibi9XzPD4eIgWzJQ0CQ3oMf+AQFWOM/p3wOx8x8Dp+g76dzyLdZR2lsog
KPyisIySnl/rs2seG9n9FcvwzdMbbywtHIRAHIR3/WaaD6/zUMMZ/WqqdjMv7ivh
zxiiyMTKjZ2YY8RvHbeemcNsZJ98N53UXDpwFjqV43KZinkpLEldR8lX05+ScXqK
dOoph2Y8sF2HgDkSSKa8/D4kliBhQ9FBMYXomTZQk3jBglmt8aNlKURNdV3jGdj9
tDRZTEU4wovtUMwunZIu7/GX5ejjb2trxUdd829i4D3frn4JaMuNecAIT3JScz6n
1I6c5rKIPpoO3pMCScfcb69RVaMzoKZHiFLeIrB/ub4dus2TAwigwsXzkgoixCm+
7MzjMXnmIwHGgEFDQg4Q1jHYNsrKXU6MGmO6NjJR2G/B7ATJIn8TeLq+HGgDObAM
qWSLHwjomAMDAikBauIApXkMruhSf6JXxTS3CoQUa3qR/HKsbEPjvq7PKkGiJbjP
8gGP+tKqFkfNLPSj70/lHgk5blXGFcS7l450bNznEjvCVoEfHsUiU5qEFUaVBPNs
m8EjF18zHNVMFs9E006nYXTZsS3n4OR/RxecSNQofaTDLlGVwuux9No1DUUCU69s
WSGurVcq28J4F/k5NZfxq9ZBZqTiO3DSVS3Vyow95IzoK4WSVOCxoRoQVsTVhgV2
CsCP7H8DYVJDgPXT8AabCbF29LVXKNwmK+YTzI4eUZWg1nVo9A2W7IybdlfTbD66
aA5gcHHXVz6623FGcFay2yitGRvgEarT84QuxGVcWfDKwOohnJCcRs9gTbjII5jo
h/yPedARc0FgP3XiLLppsopHFrW6BtiZjl998FQ7Yw8U1JJqhA+0UH2vsjNUMIWl
HCdLRS3TZ+Oo/hrp7DfCZI6nL8pI9OcSQjNotfAzYCnS1lyo1tjVyzepKDGS3J58
7FGzO7skJWZjwgX/n5EoDiUY9Svq0ch4kSjG0Fit0oFggK1MzhyFjVLbklhim03Q
wTeWtsuNeOCf5voN2kyq0hWtTY8eV2jMJUQfjNhjDcbXhE9lj9ytfFV3CQwtzD2K
PQO6bR05DJ9kfHeGaK/PDcDbGyW5knrIdA9USxRcGBP6tOsXCLvvK3E7YquW8keW
viOaHLyOFkAlU8vQ90OuUPDI8PvuRecVZIbENr5/64z/Dw4A2GCLD9jv/iR7aGca
PW502CxvpBtEUhCtt4Kkeuid/IUCF5+1jJ11drOgt1vix39gwNWujxz07udCvhca
2nPjsUajsG6X3rbjrB8P/awh7tdFUFf07JTG5Fn2eJtDBgReAETZxzqt7h33l64s
hpFdfQdFgOtC28+N5Kz4L/6/xUJKN142dlTMXD8JnLeBE/0kiCnLTRFKu7qFvBji
g9n9T+THBc9Iyd6Uz9JLIwcqGAXlQe1uWqrHWWftkOoeL6+/vqwBAiga849lNziW
5dt9BIU/fkEW8rAxTnLomj2jR3dxCeXe3WfO3Xqum+7H/UUXlGx8YejzMlReMR7O
dYn585+nbPESd7/2JuCMQ1rufYJlvs7osVxzQmIjcM+ZloioRvni5i647ssfy9k8
VD6nCFbSoHUayizx1X/zWU3IKV9WM5qG2w90EJVsxIBRmMzNBjxw3iE3v7kzQ/OZ
FpGY96G9IriXFisllkaevlP5EdbLCFXCXcOZ4RO1YR02rpfDTMSIqJIlQDMv56fL
/SZQFE97qocGr5yB3No8glU8mEsNjShkt2SORctEyxtGb3KAATp76FokShPA9d3T
khKBCPV49Yg3eUE73k1PbmLDNKDHMl+fOrki8IgePJVBCJ7HaI7ILkBTHGv8S+UU
nkzpTUVOdtVfYAXdESMYkDDgJyrKBjX5P0K5P9O+uLgls1gyxjgGN5GQrjypBP7A
V8De9TMRA8+jv/aiXnRZHcG1FJsLcn8XRh/jYhbcnNQ5m+jnovnAw6hUprDCn/Oe
fj+/V3mBGyrBXi16MXxAbHaaR6G8f5QYEVNz0sXyFgzpT8V2hOJCjD4VY5MhJCVy
I8b0ksZ24p6rSrLvpSBwPSCaxXCQdhlnel37KG6J5X1Lpb3emd7NT/6BfzFNtbbi
Q5/U8SuJqN7ML3szF+E+LBlMpehPJvChQXWA+OOj3S3+ZCO1KJ5O+6v2TzvKqQPb
Gd5GfdBIDF2hze3cRZ9JjMj8+YkqMTSxJdNvSciFxT6VzhW42+DJsRKRTNPIxqHi
GFqtNeoJAA/kmABMFoRrZ71qEKsaHnQ4zF57N/QNsTAYesrgR3nawXvxXa1Wigq1
+pJ9KA2zNvm99o4KftXphP4qHQ2n9FxfRipeEaPieTy2gKH8m/HftOfsVX7shJrM
VyyfLbtiHX2ORNdqPwUZIrFUfwCn/doC/DSdZA1UDQs6hdyvm+gWGZDkTN+uVGC5
Caj7mcc6P7yv+uEWDevuMCoc7Dw0WZbfbOVbvGHczL4HlPr/LBdG5cvjQyZXaRl3
QGmkkTitK0+aByZnH8VlqpRefvr+d2JVfv1X1ahMgRfNp+QRpsF1BHAP29MwUC+v
TrVLXyW88pPsf5uj3vXpFJfDdMLly1mPZsudU2J+MFPy46MJqRBreflBwYqxPwHU
HhdYGc180bzFGR2DPDPfvdxJVE/ucBFvyK4N3fQzBrBbotsHn559P0OSKGD2MtS6
2EB7Y9bht7xjllU2tMAkLQXp5Dqew01IK4jHhHmggzeYs4gcQpgoXx3+EDF+jHBy
+A4Zrs6un4IDWihBOxQyCjHrkFog654+QmxSSqeue9sEk4spUb3ZfjucofurWNeK
9KyFX6RMTWQ8QZOR+SMfGVCJkorVkDxM8TRT0rbydEDorJXAMQC1CIrToFdASIkB
sxagqPl8jvpplVCDy2QGwN/ldv8uY4Yn2In6euQ+X3vksuQ31ZiZ46DTfj4drIhS
tjHJGeG8CrQ+Kuz2P1OJjXhVaOv6MeT3b5rdxZvcm9lAnAJi4auik2hVAdNS5n/6
bG6bKeS5YvBcGl1cBT3qge2U7H5IfkW75OSjP6L1FNFNH8hwwNZnCntHMuRKdIWk
PwL9vf4STfkIPde/CdtKxZ7GdhxgU9OkdHCjeTQl7nIIf++BVY/4xk+b2XE6M+EP
UHwLziBJTxRcsMOkmEzqHNLJfpqSJLzG4vhTfXECTp6iBfiDUx8F/I8RJuihatUG
6gw6nxVRkWi286CWYSeStPpYA+SywNx59cGdYFG+um1KE5hL+qqN1e7zdtX+hID/
ejSRtP8dZiIENZXg9Qpe6j4KbwP6XQiheGCpxiS1f5v5vqyLacmFV64K3uXsMsT+
tD4by7aNYhxyu61bcEJXC3yVPxKl8apow4gcSG9oZi71sSMNl9OMepGZhj460k4R
cbLyHSjnC/B9NB8SRrezi6i+Od7bBxlhaursX9MLaME+fVvuiKQk7rLK5qeiMnUG
WjLY/SsvcuxJNFYrHoP/VQ2uRP2RYO0aDROEh6QuzJvDMbcTnGmB5ve8MgWNYk8g
ZEYePBdSBV65mPi4FGaBdgEbLABiuWlZEMPGaKuX/2Oz5xipz/dXqmGDs+T/3JrQ
yUpNT1RxxX2PvwW1buNUsOjt/RlNy+ORfvvBctiT26QH/PDIAdmzIec6/Y9lzv5S
5g76Or4kEP/N424qojlIcZFIFPB0j8ug7RJdYsEvr75SAw+F1MjftXKzvY7C1ZnN
LJSs1M/pcOOczzDLV3GqiFzBP+3SrByhC6wFR0utj0ujqO0MNhOcmC4WlGKh8clf
qO9r4FxrfaktCBFfqAXCL6i8NJSLBRLjtuYip7t3rpXfEV3PbqikoFBeoutG0sbB
wrqdAzsk5snje0ypJuaUg1cG/WG43OrQXj8rr9YQPqGbmmezH3tRd0NsKdWKmP18
6CMToZby4FKyelBrRVj1+ybITD7EBhqz4LDhjgQmuB5HtWJKyoC/0lPLa2BMyLSN
GN4CX2XUhN5ehaU/RBo53z1btRHXbXgVqfhUeVrk5ge/Wq82n/TSwYUuXC52IfW6
mx8Qn1ILsvIXLlBKuhW3QBZWpINaXHZymidzuir4TluAc5DXqHgmESFGm+gkv1m6
J5X/ot6SO5oGlrjGpqg8hY+iPaSvnHIqVFgmLrYuRZAdzmD8GeuEJZzTls2AXdMk
Co9uRwd8SXve6sN+EkMZtD6cM+hutyTTdXUIyQRuBFb7CuHjxz4wBuFKM2f0JjrY
2PVm0/iyYu6elUaVfmcbtlUfkxn9G8Yv+OCBj306kkknXdv4Mk5FnwYc8rfIe0zO
ilvU392rF1Jlm8mwP/bmFIswc1UgvNJfcTmaJpmI2v6EGPRWcPx9/XU3NisMstQI
QgBwFJ2L/1MvBA+on0rQcglxNG4JIgnbR6GyHbuRgjdmXZ7MQPT0bYvi6dxi+6cL
waBv1ASCnHNdMkn4MBeHtZFVTvbT8IdRS8hKci4a8U/YFS45rIstEMdU4+Zie041
UY7O06WjM7aIqDSh7GJW9lNJ67p3EA+xJ0FS8fhkc8Om7t1lssAvARwL1QBphgDh
JUaq4BP3BeCeXsb01FBwCeJzUWmchEA21PZDqwNyYkgbzr9RlEx/LFwhSNJ1odYj
DPQW0V85Oi2DFvy4CpZ2UbLK3UCV/vaBmJ6dxw9P6Uy/hRTS5nVmov3sRrMDxpS0
kVALEzkCCunCt31+JAESiaoESf86guCiBtt7NSHwYc6DPXo2Gji40/Gu4i3oAZN0
Jwwn+8wShY+1kr5iORV9dbpRZQfX32YN9ZEeTTAxwoNF9MHv8hZbpZBzuSwh5qfM
I6CyZoutJJm2Mm2MrjJfbAD4cvSygFKhT6heKCM8eQVsDqQPEXI+UZltU+F0Gy5u
kqx+DprspyOp0NZzhS/TdbG1M+lTrQUXPjRPCVc2K2CWXtzff7yJYXgjAjY3RTTm
GdkMUMuHkcCiVXFMtz9qiHKRGOiNLup9LRWkj0mJgBJuOUrGI2PlyLeRStVWxprc
8/yS80nV7+QuyiapQR/5Y+yTaiRLHjpxlaLBFQrg91Qcu4BySbL5/5RuTSLzu8pN
wjKmURkBpYK1/LEXJNFRCeB9SwxZMytlQdItqUFwIyn8RlzSxml1yNpE7BLHQNKq
KHpRHpsblAIn6oefuk1+njfdoV8El7Q+0QnvybAufZatju5PLyEMruJ2g32r6awS
gTca3tzFUgqJBE8UgesDxc968FMDnb/GRe7zzW9vxf3uCgcSMAohNFhM/mXSSNLi
vHO1bD9mNgHFHHC2aYMyZpmj9ti2SIiFazCeFjJCZO6QTQp9Y/wywKGASliUCKkL
shNngmxG3DE2tc8F2kRuTJ0bfC+CngPHtACYtvAgtnWLee3k/S1/QGu/Sa69J7Oe
X4r9Fr6d6fwCMyezPDFhKDOl0xKAio+ij0xomXr/v8iEOF8HPs+DZOojQMvV2y0O
1N2p6dF5hO3nENjQ6K48irkOKi74j98lC2Y7nX0PxXD3YDBurjE8PJejThdWddq9
NJZRen/A6htdzQLg8/jtGSOfKeqH8FtjQned9tPD/TeH+TjXqqIXQZo/86mZ/ePK
+jS590nLq+s9wb28ATb+CJRTZ3FBYOtFRZrB6RhryDxR8c9kdUdaliNNTxJneGf1
3z3odxSn20zOAxRXcGr8Zneox5WT2Zy7QwsvP3+Eb7cKAWFPwpp+JsCzAifLfuiZ
2mYd0/75IA3ZH5OxNkq8xpr7Y+wpE/Y46CyjTtUUuiL5+yGfbMrLdGwz1bwky28K
7Y+hcpt1DQTMDuENCIFxbBSF/XGdaWRW6DyEhr7CLi/R25m6LOmQRGsGU7JwaDno
P7WTWorCZqZTfQOeiLkbjNvWOhW+xoPvn+vgQRFcEc3H2cEvu/3Ek9mjdRXeBWNL
gYWoT7Oh0K97dqK/xHmRLyfhGp+rZr9YMV7azgNTGAAU66znGYZWKoQkDpR6UMcb
iCLvESPtjKMskpeqw8o/b2q0nYv+RNVJfkDMTfZt6Le9Lv6TvYBRG9enH1eXiHRK
MTsYZj92NvMNxp3KhJ8AXkDNRRuK+/JnbxwEGK5+UTUXoEREeRU+OsANNnUNEYAi
ucfh/1wNid1iB3HQwVtKoGkBJCet/UTbxGHZh8o3+sbU0XWMdQb/PGi7NLDuCSk0
FKotEGhSGTK0XZMdcufAIJtGhexwK+vGQovEOOu91KhN9w6OZw4ms4WnINaYd5ta
XUZb0pGEsJu8j9GWCmmAgKLSzPgP+NG3H/lRFE/ECrN0M9bqllHJs2hxd4IP/hve
Lu6kK/+bAJY6qK/pJn5Amay1PBjRovBOn1zr33/2dhzm4InR2vaayXFcuPzqHd/F
AmPJ1vhnZeyRaBEuDpuFFCsahgGlJsZySgMfdWy3g0qZpkTH5cbougNMbXproDqN
LW6vLkosLbmjwlaR+GjewEpPATCXVKN3ytSELf70CeuhiQJYT0Lx6CrKV2EMcOlz
5QZ65a+lFQ1Lhr2yfo8dw6oT3nHTs39w2ChBLfHkeWWw2BxSBgvoRqj9GaIWi+2Y
G7Dw92z4lymmUGF8lwZDk3IGIQcEIcuROw7surH8RSzHqnhYeWS/Odcd5dKgn1f3
bixo3hrQulHSJEuWWk++tPbXAaKFOl8oCGJpvoWPMkuXxQFzmu/oOsBMakwfTGun
BSOrAoGgJGkLQo4bN9V1XzLvWNhU3sgNr7OgynGmBpDjMf6gjNv6r9GgboMzvKGd
bIkdYaW+kVccu5Nqb89LkPVlXPs5sY7vPAIPLfMF9T1JmrjdnljfSR88uRFvTe6q
sA4VhRcive5IQn4LPk2x2kuJ8/Q2tGh48ipmXkYFqVaPhejFHTkFqhIVugoHZKv0
R4vPqR0ndp7Ig7xx//CPr8GpZL8RokNCRALmZQodM0uFqBp7KQNLxP31DyZ34+GD
dxk91UAQ2aJIp15QrlL2cG3MW0PcKucmoJkcg6v32b5kH4VC18GaO0J6tJm5cOQf
Ozy6aGBu9HAuB7gO9qJBNuJ3Os0O0E5IPftM20UEaAPL0dWtNbkMDF9Bi6VQ8Nei
/VManATiX4K4VgjM3cHVda0dx4mmjQB6zFHQQCsqOa72IaZT3COVIdJgA6+P1RMA
PC7fhPANta5yfOhKQ+29B9al+s2QBLTOylxVM8v0SFpfZ/Mc2CpMGiRJ8DKYqivl
0OL+vGP3SfnYFkK9ITZ+T3oiWEfwOxy08Fto7kZY7HrwBR43zO8DKR2WLFN539RT
PqJiXXSojkqmX1+ZT6hE/20VMx8Dx4r1iKTtMAu79nPpYCqR83cwqz646ORVnrar
MLlEtGIBaHJS+XqKD3tGlTmV96G3OmhRvjuCJNrq5gXpSdyCj3VtIlQiK8vy+yNZ
FFA97q6VKP195ncndviBhAF4E3Z3aluS3GgLhxorP7cb+eNzqpfxo3gqz27nAl32
wvcercBJaFQIfYwnfhRoi0kg2isrq8zCVF75AK/gs6ptyC4RHB2k25ohajrDYwjs
rgH9okjNh7VefJ1djkbz57IJ83hMaK5ctVIKnl82bhT1x2fQphwe+gZg8vUFcRUi
69td4wHw+wlTG1w73aFWyq6aj6sYn7Ny4GW9tEsWRBJxwpSFexkUESiVWJ/rmqoC
GDp7RMGv03vCdVDs2zKrjZkjaTSS4IUbS/g0BfppUXVky/haEDbB1HBXtkceOjeT
+P3CdJ4ZHrrALwkKGYprDF74Nqq0iKEsXhDqBhS1+3KxyNSy3JIC4Oftryo0TFKQ
nhbE0geOeCTPjtOQ+PrfNy5he2GnNavBD+Fl/lJKmgsG4Zm3g+nOs1N62K9lE1E2
IkW9nLRAce6ZTj8tPFCcAq1L4b6spbDBq/jso1XD2O9OsGpik+GLU6jy2fe51yyW
Zdw8PRy2XFkCTaLcffVbbpyv3FHM5VS70d0RmImnQ9ZS9DetImXtyx+daEbXdqBo
uiexcoUsvGAAxzdpU3x/DsGeLkfnLBTIxn9dFgmLyqnW0RhrOpCoxjXKqvW6wIVZ
pUel7FW3lrNe45npzEzRyFw9JWW2nQ1MyKT/hmG6y8LadHXjWIBeqQW4Q8u1X+Np
XLDJGfLfVq3I2T8MlI6U2RmXEPonccU5TeP4IP8vA6ISzjx5q8d4d6chBdhLAomQ
7gvqRCCUaXEfsY+RQPRnwm8xeLPCoDhA3b0ShX+UM9BHcvwp4AGvMFEFtUK5dQmJ
AfXpzYx+TZF7li8tnldiT0vEouuex3iSkUJJHiFHdyCVAUELZDDKzaguCd71hvKC
LsR0LAn0yksAnqoCAIeEiIoSDhrOQN58zqgrUnA70uSgweyJ2ZY4Clhu40KZ5NPc
JbpzOeCHJ3DACnC+NA9+5LmGnWA97GXMpotolh8LNRfOm735fqU0yqhE25QYqLWU
2noHlmL9eS1FwGc+DyYRS/frZjX5OMMyFbNQD/unsnsSjnfCgCrGBVM2/+IuBKBw
8/zO0MuuWcnXSY2U+br8oYuy30MPeO4UYIEQmB0YznVN/iU1HJAAG5ItIguP+qgG
TS4IIL+n3qWCX34500dBh59XKdQW+28Eho66/UmV4Qry8HqTQVBCFFlUEZI0dsvn
eOkq2ILklYTFy/vOX+yExNgw6mqJQeveHAcXs0j/YPsr22y93yFEfBpCq1lFljAs
6bGLFTiw1bSFs4sx00pJ1Ur+b9+asJnoV6R9HhQsCQdfPO1i+JYZU2zcrUBh4fBN
rPZQNNXqH80zsju/tV/HuZ3gatguvRWTB8V0/AVcAfBnTgH/PA550pyFqsxvZcfl
G5NPwGMYEPWmytMqjb0X4OxbA5jIq5QasXu/03CVoFgd+mpmOxmNjYT6LuS7Buz6
+htKUod7PdEJhFIF5aS5h/ctzRs196/PUt5a4w1pWexAsll/QQwGpIw6GJCQ+jPW
1K+2skNkiuWawp1bvoNA/kH4bken5Pla0HXjoP1mdMk6M8x2BV6AKuYo+5ezbXIK
/XfFiy0BkqYyzP8TtKeWfIb6XDNxTnnhlGM1GSO4tc+BOUV3V8iLTaLN+bhu9NwT
Jj46hqDJgAlmzaJKq/N6eEKd18j/SK4AkPxOXlfMtT7oPEDXtViV68M1MgsmcZTq
Xi4ZL3iIXLy7fvZHaLGZVAhpPE0R3UJq8znEMI2Df8YQmRcNbbZ5iWQgwwwLmvJS
OdiVDpMo09ToU40XuIG26ytItIvHuv7Wzs2wUuNXyfd5o6lByA/NUM8TQKj57Tzo
51O2xcHGYx8EyAg9tvTHKGWUt4JovAfiv/aWRGQBo7P7ylzkj0g61kllJEPhArXH
cXvB3s6VNBlX49gpkqFNxz+LDDvsZmnbyge0QL5FKwcvWo007NatTiFVTHXvzvHV
ti3Qy8HeFVIyvrbrNkpox1UFqF25Buu6YB8Y2bVqfNygYTpFBBZRrY+N8FG3huru
VXp6C9mkDg5bYLqIVsuabmzHEpPwmge0gYrVNK/gJ5eKzIofo/LOcmysRKyS295O
WTPDpAENqDuhkitoWnd7mZPhJOfriewZtH4rB6xK9psaN/odFjT0OQrWMrdVsfd8
bU41zTeX3dh1Pk6brJRfS7V5xcJDkE5b9dIL7Liii4pk15z/CNSEHmIXq2lS/Cuh
bz3wrwDn9P42tywttSaLlt33ihtEFSr33ZZKn+QN37HTKekQyUQ7CuulDGl373eb
lF8rBiZxDT3iC8vbEhEo8eWl6LOR6Tur3qCNozF/Kzf3oYAFLwXiarn2n896i+ue
IYqg03Jtq5YVvF4hPyY9Hya4apY/g5RQMNmu7a4tfphG/zlYK/4w5rI8SWvYhETF
DEDVJa1r7ZH0zzB+EUzbuz6pycCAaMXNMHfg0PuPGlaAi1Q4WcotSjeZhMjQsnol
43qDfg5JM2XL+MT9N4QepZD8hVgBgoxE2/gLQcS/P7sZ29Y/h9DknlKtxCkbNt05
Umqq44T4qlQ9w//5HVzJjOgYw9gg4RWt7+Ys1ge3ypKDSu4QsnKVvEjYnEj6AnZt
N5pIPRoP0SKXSpP2Aw74DoOWXYCwNY/R/LQo4qGHlXE5SxhfQcfAcBO66KJdGZVK
WmXRc+Q2jt2FVSbnTIvmLgexZd/hRtF05P59icWo/lGkjblc9CzEme2KWvNqtXcb
FxQ5vQZjzCwtT7CweQFsvij47MW+gatsUilIfj7iDbsKWKGg7QOKIHEu0+v+4Kgz
QP3oq/H9O4t/hggDYkFKKbp68GZ6mNMRYnyuTFJaY4CkU4ojgmhpQB9RCba3k1oP
j8HeyG36mAOtxNui4rY/FPJh2SqWpRv3vn84F9uI3hI/PJops03hjGoweOwL0rvi
0mSpTInZeP6zTzuaq+Xg0vMZ6bboZ43Gi+clCnRXUr42BLpWrUjuSFZTgoOKKVgR
snkqRnE78wN+KFONJVOsH6o9B63nmwKdXEy1gL3RCJViIKxFME0ZT9SoRuHIVn4v
jMUsMSfUNdL+tFdp/7UEnmXfybCEcZAu8O3kp0bVBwB7/NwYnr8yqG9LcxDmiJFH
w6uaX3/YVE9koLCfoPoRzHPy6RSn3YyDj2tPr2MEJz2ueHhVB6CWe6AmAIcUqFXJ
GYnBr5hzJbEcjpKHEFs9wzFie86NyhgaOJeoqANbuqwH52HZ/QkoSXjzvKn7bTPw
TU/sAD54DJ6e7+h9CkgpLXtHeF4KRgmS74aZMcDolqQ14+IrKw3HyQpZPQw09gZ2
Q4CNpqrmyxw860BQNJrKq4iMcP+3oVONKYtoJ8efvdm5fvu13LUaCOP9H8Ehnm92
8T8YW0Grih4CDBr7pO8Dc4X4cxl/kywILnzwuRh1qezY7yHxAXTvrcoPe1iKjdPG
/jeOn/MYRENU1xhZxyh3R//bT2qpDGuPVkrQdh+8ITubsksMFT74XF6FXtOjP/CL
a6TY61DO5eAvYxioKkXgXoEVGTw84Z4mVqaRKwMO9A7P4pmzzlHhQQrk77yOwPQZ
jCggJupblLycuGBOs83QB8Z4+OEd4KuJtBXaXa7bGuA7rl48d6uoVikD782mOfKL
+bL1+Zct5vHDR+Y/mppJTcJ+6po9f20oYurJ63AhmDDWjlgYWiT5cTWYhIs1gEvu
ygId5w8cRilQPO3geMjl0s0wJMnxGE6LKQpnKUGUdqlXz/Bk1EcGIwJVW81y1B9E
vd4aEUumDHZZzHG8gugO33ZbHrqUOWiPqGvh3fAW9BNJjjyDEPMRePJS6KCBgztN
wNUn9MFU2gloui/aXU3VfZ8FnqZhM+iI6Gl3Q3BHUdmS3j/E6456yTaH76sYoAzP
38+PQB6cI8suv7VKnSCFkhPolFlqs4ifRNqI3npG8Y6Z4cpQUgKpK/L+avJk/AkJ
8/dG0O5f2u8ioeR2rdrOLgGzT+sdW861auDw3NWP0k9wVTBteRuBPdKFuiZhGrmY
OfdfZzhxMnvGdVLWCmatXnQk+9AzxEcG0hs8LaYor69HIrLZrciL9a6nku+HIP9G
EzBdm8l4RiiYqMfme/rj/Siy0PdXx+EXBADVw8A05fc0EEUv4cVhMUlS69WMAJBc
udtA65dFYDMr0bprOu3RMPd4vQbSmZ7J8KDuQRuco9QL590wFf/FpsQ8YmuXgPzO
Sz8FIvqO71YVyns5jXjQj+q3N3J12lGDcuqbjSKvjam1a8OlRguLwdt28XFNH4Li
cwKHijI/sp1Nk4MiVWP+2qmbtrKtBQGeWhXciUbnxCEB6DXqSe603NLhMnDfbpDV
zsCY8a7bKLk9Wf/bbnzO2GXYCEsEzqu2ZC7R6L17LvR7eEAjnA70IesfdYhXVMz8
VK0beKkIzxjGnZjguZ+3yQNqzGGWc3YuRMSs7ppZGbqS/B+y78trC0yr7BotKeSn
XDUvcNy/dgjWaMP3PCw6drnnHmbVDgsZ2y+xilnxcpz84UBslI+IOc4/HAdoIE0T
2NDAKTbfkEAhl+xdvcQ7vceOG+riTYIfW9MbmaTAbcp6UGVG1UsfY6uWqIfo0LgY
tw7AdHFcZazqex3LUR9TmOM8fflFAhFQSVK81E8Ty3UdjVGDH9Cr++vrWJ4V3Hf6
1dfP7DzEjHlkMH9JMQbjrBUBWRUEy5EkNfxQLmzE6ugaknBxnMtCNj7x6bcCgXkH
eoK6q/lJWSzInvLR/Df+4vx808U8GVgJjAABWZ+A6ClhSHWYsoRVW6xkWBMiMqCy
O/qa9NItFddjBf6YfYPe06USUEc9W2j0kBbPIbEzTsQwAOKfZQ75fl1hm3JbCFJJ
3dx5pjEInzP8pg0L4V+bJE10uQ6im1HIAMnrzUNMoIcpil3BCH/OZLvoptZbYI8k
rA9ZoCe2uM3C0aQvWNVeHx66FKLK8ALg3lmTWErhbFQKcOldaxCVgGoKySYvOnfL
f1v2F9Yc/JcWrgekvvE4GikZSc21rrQMNatuyT3pv6ibr7gP3IWIoqw1AjLqPGsS
QpXG+EBGfVy8JYLe9mRQX33uN0A6c8vjiYTCV9PWXFO31HDkInSmSFzfsIRR/QS+
POzxdueandm8ZkMJFVk/vAec/f7a08L0ySMbyZkRxvDpHxwhzAPGFgjw/AkWFwpc
ywPoT68jfNQsQDaaJ35esNT9vFBnENBwHp176xe2NTmSKiipXBNv4Mg7kxi7FE9v
Yok8LrhRRkmW9PNGrJ1CFTqdQtXmDmxsIze6XaruixJrwN7Xmb9hBuiu8MmhyIS/
mm7H2ez52vuntkAsoBo3oMKde+vTUVkDmnYW4/57Ma3+XFZu9R+dqpVN4FYsyTJb
GIJu7pnefsnpMjn/eyytS+2Kq3/jyDwFqC+8CKmRdSAYU10qUVGGrAf1baV/oei9
phyu2y0dPdWuageG2u2t2PPrba4R6KUQ3jbHyIUWoNPBiIdi2IeKX3XE9rk91uPQ
3soSEwJlxa4az63lY/IC+f0Ruo0ldCZN94FdLLrDtjRPrLDkfRK0uedZhBl7iLWS
N9t+U4XJzBJO3fLc5Wzbc/ZYMgZc6cQb7j+oB1tJZLTWc+o6FQLsJoy24hOOvt2Y
vLzz1Rzgh5XRVjBX8QkLt9BXEK/6eAzi3pdzvFeyshH5nr0/IxnJZLFn6vXc2NsG
fpsj+YBZlOrNoabe98t2crEZPud4y7vWv/uCUwUW4fbIXXwFYqX1Bhr4t5CJwRmi
Gom/Ck679PxMl/g2hkyX+BIQdnAVDkDe8dj5ED/V46sHXCLtjjF4SyCvon7p0FMB
fMNcj9ng860pBib9ZlssBHQ1q/+FF45QDK8zIeKMsybQMFS6sJZUbyQXrtwNB/p0
i3riiYiqKxSaVfjYGr9HD1WP4B5v0G+bR/x9Iynk4C0sArv37xjmf+Z744CFY5ZT
GKAGuu2C8bXhx/GJyx8ryPN05SfNSfjwV0/J/9EkX7NM8EtyM7o2eWOwN1eh5Gpm
q0VsK305OPKEFbxxCLJoSGhuKzygVXbPoT6eZ5KA/rBqV2rLNBfL9q43IWbvMlXQ
93AqYB2lduiJGBNandZhScZ1NOJnbTVPDHSVNwDZp/Ka0K6hZqF4X+H80/+BjYN1
e1lIHQQ44W8E/BW339xIhSD7DeHYY8cUCb9BclFhn+m6ce8PGF/4bDqf2DFPAir6
8DvInG1i4gw6Zfg1HZxsj+lDDFteVpkMraI7izcEkQy784gkc5yJBkOaPjncyjrG
oJPtbKP5LflY+CXXDI91a5Hxfg8EPOUE4Jnkdt7vIgzlLjTOMVxWQL471/SVSmrq
rKkt1hbHisG8kh6rtXPl92PWWVupfZnSv+i1KNzrHTt/W3a6CLa002uwsHo98hEC
zS9o11Wyiu59ayMUSZDHgSeSeeixCUe9ZVQtfGMELxM9zlD8M54HqyAcIRIL86kv
WQ2pnrNdfz+hQKUHY4tnpqxc4mDCUJQHxVQGN22WpZCOr0ke2c3sSc8zbo4avUEj
xFTaDAWrqlHUr2dzA2dTAZ6fY2KE3WW7UNcFOTy16x+aKCQ5VGg5KXKZXDE4VEjY
H+EecYeLMIDcyz167Igs8saLj7OJbR2guarzT60igWvkTMqN4pKeHAeK/SM95GMW
NNOWL0408tHyZLs5pHm+6T/CP+w9R9W/89IkOCFGWYyCXrij4ZGVMKjQnx9w7xLe
DHmf3GQzanAe1aCHD2/ZHxCnOoP6wB5xXO+t8MVKU7DYqdID8/Z/LXpwWylqmnK0
B8kmEaJ19jC1QjFxJjG2TwCJm+/MyOHGJ//7Lma3uDIkNECQCvyo/OFtblu4r0hL
OZ7bYrQoZZ++3/X9hdcKf2I/jpJ3kWRJnvHKDgGBGWQAg1TKK2iw697ZEcdjStL6
pADSyA7z2dkQ2BxW2iQG3YhrjW1vKZSkzEGeFO1QzF9nFy0m3TyhaMWOUHo9Jxgf
yfVHCW72oj4wATgbz1RQ4eO0fzS83dlri9VO3ghHGBJWF6FcfegshwsoQxWOZKX9
sL3PfhO4L8Nnz8RG65z7vDSrsxm7QcIYjmMtmohmnZLwAnniTmUpUvlRIR1tLqOf
ZSyDpQvu2HJwgkqlQPWsyk6fColyFluaS2jknYd63+RNjrnpa+RXVq3DNKtm3pQ6
6uZpOVRxxFcqkz1tSO06RMrN/HTP9I8i8bLylF75y/ZVpLIAsdu61KWTAMtI/dv7
aeO9mY4NpAV3W0D1mptqNIdfZUFmiEF3LeZOVojoxtcJv8lScR6trcBIUD2+mnzT
kK95isFG1xFUsK//v7RI54ftdoiW7K+O91U1TO7mXPwo9QbYy4sBxUDXAuXHLFH7
B5atyux6sTquta2yCSX14LihUGFum+nTVZkB5K7XhBDjvYcDfD8vXX/1L46z/aGQ
vDi7IR/v146c2a5i9cmpFyyJWYanDAm6RfsKHrUBjcmCujwqUBkKfIIPSqMCoBTh
YZQKCrgLx3dahG5Vp4sz6bvHOrgfRzrHCCxMRFU61EY8fWzkyYTHKzzX0bU5DHD0
l8JMZoj0HG4uW7w4JsesrINa0cT5BUpN6vQTI+N8ulbKNEvYXGVuggBlXsvAYiwn
ylRT4rD6eJtMP9uNz/6Mbk52MrOf0YwhfB+v6PAUZ+a2sMKq8fuFqwR9vz0mbBpy
f12WHw6JOuO6Koo37JIRBwjH/6UKm12uM73dRrTZwpXD1Ub9OBftPsSg8YJuOYi3
q2I5gCR2cKXfSFoHFvQ0EMbta6OF+Q6zxb7pQ+xsmksGB3WC0iOlKaum2s8FSvkS
NK5IH+w5jcgySqrQCsUQb4a8JYpOBIdPfpG5uWLJg8ahhnuX7U38yIK6cpjeGmtD
pOMIDOs40SKFcmpfZwCpWbFPz5/BwtjOqSrxVHYsmQ6WHWXz12bWjWR1dnmMGBZi
0o7+i2dYkli6HaylgtffrbXisVUkMDcbjSJK6dHCtnwqKYPG79GK6YqtQNDTfWc9
KTlct0LgucBHwtv40vEWfcbr6vWCHvJGvxn6em56e24KLCitNMdJZ6NbJvLjMNiq
K0IvDRGoT5GEPAvaMC9on5syuANpjXJb6OQVIAn1xi++fIhaMozauXIzYeasFl+2
OxImC3rnt+oXDvp6CVjppsu4Xp/uvVk2ncNy+WOiSzVtAaao+Y6duVrifWVWsHIU
UqPsHisrwwzMLu+CCk2Rgfe9eVEGNZtOzhFkiN363dKvrd07SKTuNps4Gd/9B/3P
U9v6OkGUCGkkDSSA7ZTAjkY99Ol7bMs1U2zmbfK9m5YaMbLfDECg0xlXZ6lHMT1c
F0WVTsHv+uPWWJQWM2Q8ukZ5gNuIl9Vh92TT5WqjxakhryVJrd6DGe0aqyruKC76
e/0b+mSxhWDQV1eHbmR7stxUryAm7rzdvA7XyToDn9E0lU6DZLxlLUWfAJxIk0N+
CF+yhaOlwce4rVRc93ALBOkgin2FMJ+l0uR1qDeZW9PjzFz6+kfK9TMAMzt7+FZ+
igiTSWzGEXrGYMBhKHzCRtGLbOHDs2IPw16OI9N3jMe6ZtsrGzK17GsF/yvOkvXx
EhgIBhhwD6UufmUx6o9W0C0uhLkBn1KtAGQJ1qtE+KPvaRL/by4qOfRScFGuCQcO
buhXec9nNWfcEqi+bnbX/cKOxirFdbUKqenlgQx38Usqk1L3Btd74J9VIOrr8fWp
xkea47eaajftRyQpVT8Pgxk6Pj1Mcs7uJxqV1BGy+iY2kATmcT7BzzY7e7aILgyf
gIXMiGNPg6Pi2SQUeyXgtZU9XsOE0mXFTsewNdyXOhxmCSGt7Nh6pSIdD6l+jLi7
ZNWODcXv2coABJQsz8uEZSMkC38hhsQqSAZQElEplLS2HdiP5IojrC7gvAr8p0st
PDRqgY4lf2Xw7pvstqjaPkMZBVHZg4XUULWRUFomOETTMmAKqZYfzh59Fjv0vIcz
Ywb5h7T1Dw2Nbl/ViZDzYemNOPSmBjDlMgesWI678WjvcnDN9WzEO7IxFTmTIjss
5nMOInBrJZssgBbn/IO8VA/yvKNXKIBo1+HqT/2jX6IsLdWf5KPm7vaFcbcGS8br
Cw86z2tTHUtyOrM0JjIQbjoFRfIQmXcOQGWf8d4hWY2KxFMGgmYzEnATl63QAE+1
14K+WNmH6e7fUS4r1y/zztPbBwGLiey+mbC1o8ckt41wTPFeNdy2rE1cbH7Y25p+
UsGB5yLtc6SE3XCOYm+32h6rPcxttJ+OQWJ3yP2QFXI9AesADsDAihK94To1OFFA
x27ux3Mq8qDCQqGNwbrAf21+ukkSOEqd88i6dEwiWO4Z0XzFLp7ruXAy2IGh0zFG
/mlTxwWztWeq4Wifq+ZFk/C2/r6obeCTYf/BZYTlmvhyyRh04ozIFrE04LrYcR1I
ba/KdOK6bwP3sTxj6KGboWCEVKhxgkDQY4AQVawAD9Q3Tn6LUPz7770tIbhQdOy/
skXjxFq1gxioFlICN32tiQxtYP2bXSHRJ4jPYjiS/1pnQ49oYugDjLCWYDh5YauX
NYU/t7vCSg89mqErCG8Nmvepivl5bKYjH6RoLpvYdUrnJu154n0r338P+b+Elj9D
mAGx6ZO7P+Pzjpg0yRrSpomasyO7PljN9qBsWo5eD2WRF/3Jp/0EgNVYAa1uLzsk
1Vlm9LM7WpNss99U1DX+ztHblLNG5BN9RKEV0DK7mts0OV9IuT3olLM4OvCOyfZY
Olm9hNH74TyALWJpYPijsVMeQu6bGRti3elf+4vOZPbNZtqczxYCle/bSVoe6ml0
WzY8gqSuzucR9UvElyqnk8i896JHEf8rab/tgHDyBeNpoWPahZgrB5Uip5Ndwn0K
lJ2Ugldj73Mpa5Ub3S4G6Ts8OainKXHf0EPrggCW7bIBp6fBQO6VHV+TVJzjikK1
HTtaxdEZ4Hfdx8OTtFBcx5n6tta8tJmpfgrc3Kx/Lc+PXpCqNdFNIKVqm2+V4hPD
2vyPQ+yxCoMnWkdnHYTVgfmVqNn41m+VapQGIXf3E3lpBEqrLqEcel8GVeY0nGe7
uQa5dyeYp2eFDgyX12Cly5QTML02aIKNfiemr37L9ZCIluMTeak8aI/eq4jowiqP
SWxu0Y3LkCr6WHwO+d2qE8b5+zKrVC/BEwODy3cTLzgP3RH5GZOMGdIQwMsDj2VM
64WjiGWJMDskal7q6OTwgeD2YGTRSf/YvwVmEf/TOXIBq+Pb2zLEYKF2NjOUYiCr
Tru91O0fGnMjW3uTq18NWuoBg05u9FZkV8nBdyCyEahUyvhDwGYtDL/edFpcXgX2
cK2vwu7Uhw1OmNbexf+nB97ARo9+WiDEsQz6OJjZlE8ev7Guj0lARTlazUKi/xCW
SDksKD02nDxNzN24N7uqJS+k6Nn9z2FAVSLfWw+eZDh1//01Neuu15VMWu2IM4+c
pCaSlikqXL0pzMetMp206wGBUVrtmA4/A0KowvCz/OsBhxAgGHZbqCVDq1GwWDVD
RpiTQu+WbH7R6GhhzMlFpVgvPyXFvNMbr9mae6rSJbPp6QHwmWXVmb2PKC0dB6dT
sEoQaz4dmIBmE+Dig6Bed0ygduQNcyxjqNFKLS85UjEsqQZ8IFvo9wD0IYImBsAN
vQtjjHjUTznIRsUzZ5Bt9iB+8kVOtsUatF4pygfafrHiyBW5bHg+EpHK5rnDjOrf
7oXKTmOYYKQc3tRUQiyH4rPjVj+lYGnhd/i1qwrv/7h9FQ/pd9d24CJgqXLP3MyK
RxUMVyhmQKAKNm6VUZiGBLbT+V72qa7+Gg3rpTL+mETmW9kJQP5fHOjLjvmtfdEM
QyXZdEdoieWiNao2xvgzhAQjsSXH9mko/0gMXPn9Jx0of8um4GhWGH5EhrzrSqZJ
xPNeJoMlFqmythFz6iF1ldOc4vKZL0i3QBHqYms4X5FfkqBifcHxo4Ccq3BsItAx
GIwa/2qtRtbQkA/bo0u09IKM4dUz8a7j74XScVEv7yW7ItAgkrXa9Bd5AiQy8WxT
uCjfOJTlYUAJJtd0WKVl9HvrsRG1oi4/tTHmgXjJe7xsj4d3+wKvDV18sp/AywqR
7ArXKUBJWh+o3oQWCOA+QnbEoc4fztoqdacHY2tBKs047TBf8Kejfs5bDmmOJ55C
bFkFLtR+OTFX3o2u+Gndzq5Ic0yAb3rWm3q6uBOZTkwA2KSk7tYSutSsLMddfiqN
LPyFE+GB7tpZEEqeXhlr3LpsOIauQLOBD9RamDA5m9LJCndww7eVAB443Zdk43OY
suz80ocVl+W5zxwLH7yW6WBg6ijsfyjguG2r7SeIqOKYFCef5YSQzyjgMckWmKhW
UpxlRWtCLTvlnJytANotRb4z1XtSrEaFuM7q0tQee7xNFiOObjlOhImQi88SwXVa
SOwsT84p1GTxZlT/ylnWJ4196gimd4NXbLsk+3b+3dqsJ1B1oGg/PvyJu3zTZnuz
obybfPggP0XfQsik21YIFMHTqo1+OuvE3b+FhGcthvMMdvzo7aJSpY1dpQv9EUV2
S3Gg07AiyOS09l3A+xPi/qzuEbTuDLgywj6dJNCbjeIBtfxBZbVYQa1CLzrwqZRu
vDSeEwsxtFBNtXpcz/PgPgxt8KYjmQF2dnVhkfV0Ncup2FbF2OupIcQ0TuixRvdM
Zzn9Vt6rxfECVP+T6snkPrnSWOvjxYQGFEp8tqWiJzZtP5qCmprKkwreT8EYBwkJ
BJ6Mlzvf+Zvxu+GkQkG7egg+DT6uwUVX6go4ZqKCJ037jFvS9J6Gy5a2aBUQwQsB
XfFR8/aOOS/usAIkNERQPW+fl4nXipDhpwULAUziaRsHMbw4pcyWtqgdGZZf3P0N
CIBrkEbT5xPtupgh6/2TGvGSvYKfNQRrlyXKYbfl0WTTnRUq3sDo4ewAcJLJbmXe
G0Uknk1FlAfhz41yUfUEzrcc2rn6TygHYUqV1A3fDO13y4LmD+qpdzHOe6D5TEiW
7QpARWn2C+m4XbiptYzght1GmeyqhY+u4qKQKgs/6uij7d7ekZ1HTZRCeWjvAPqW
2ke8gXAd1eVVfxOiNm0X9qMFgeFBuWN9BedemLGHdTUXZVzXj1OhBmlz94ABdFCD
vGyZYKNaObgElBjIJBNi/C3BHyUp7myF31KaeCMakVIVqqFTw8ZoRs1CJTqx+z7K
+98c+GhxiCRn8QXWfeD8PMoFf5d0rXZgZUci4PPx9q4R4gQodfSbJNGm/fYAqhdB
da87p1wPDKX1SrOgbvZh+5dNaDLZDFiIVDjjrlkiqlSvBKyvN83k8E9A7Y9YbIRF
KwcPeC911j7QcJrIvu4m46uOekb00Nm6iayCWqup7llBjAq0p9jDpIrlX9tHwjCW
2s0XjN0chtDnE/RkQRs9QWl12Fm9nLyJA+8+EzZGVE2ZEU6kZebHSIASl605yRHd
NvrtAJrxe673Fsildq2f22zvnvowIVpRHKDcVW8iSiC6NonYTfrCPsGyKFpmXECm
wPftgsv+ds+AbWMvVl5pBz3xiSIOUmuoGWrnTRKKQmlVo7HoLETZ6LOeX9jxPv7/
eFbtZTVh/TEnaHtGpJH+La1QTLPpKFR0ZGM8owBA0bfY3lgjmI+TYnqJBZJRnaT4
DyNwjjq+EeXr+fnlPvjLCyOlOCfuSxxRSvmyP9ynnth3PWwUclbTOHc0wGufY62D
N2A+VRdAkl4ImpVC9OnRF3JsDCLDQlQ1qDItSAJdcuwbziSllJB01k/MpGnQm0tP
FMkA2jghg55IfMuVDcEKEC+4TPGrajEK6R9cmQnEep3vnz4d0j2kO6BJ/ygGfN0w
F/Y8TKgXVjhx/YXO0V78xKnLEJRgqOKMjmoswydyoY805+W0hTS8fKx1NoFNeDBz
TG4xQ7TYEJfN7zhWjnfRrRhC2S2aR0pvncXggHl2WonYE5ueKMT1kuB1OAq2RF6j
19SSo9e1E4wLI9bdXuIOgDVAdUXwfLuwXQu7vulB/LzGE6kyxmAzOcExDnl3eQVN
r5Cpy/gaUMUSZq/gCXttr77kIUUdRL412D3UmQpUAYGh30DMImGkHZCMrufv+q5D
TxKHyu1JvqtpcYfwQxPTGKm+Cm6Lhun81yoFgs7GXw+2+6MWKGi/B9IFHwy9rBg3
lEW7kgX6SsqHAEK9MfBVlAq1xR+3DFi4gwMpCtNshOd/X5wP0Vqs4+4v4BuncXMS
gAiAXdiOw8Gh9iUk+c+xfmMMZHY3S/hRh6T16CsdBZ9lJrgR3Ix0U8DgwlKU1lPt
xGeKSf1Ozvetupb81XOPbWE8LUqV33A8AyYCPXIpM4hTjYUBaGXZ6Ngh6PpCvWfu
mHVcVXs1pqrrjn7sHp+6TOyM3Qf54ODqKIOyHLL1PEGd8zThXkSir/ihQuaCPeoc
jxtGNV4U8TGPyOfp//45zWh8TqjqzvxR5bdHN5xTliCq8VgSHFunnzmZkRuEoovP
266WIyH5TGs8f98om/pDHBdcNceUCv198cU1fPbsRc9ua9RPnOX8RYq+GKLoP+Ic
N76ViYQUygD9l5gKHaIjLRILfcLi9HvDf+EIiwBPiix5nmBAoNXRmR0gGIYCBt9l
aIozF35SQ8tmQsIv0dGwwFbqETf+nmfFyhHQdt/iwpU1BtERptJAWKz/TdQRJfJc
QJmI921I2hzZXxH+2H8o9wThvhef4WoahvR51r0yzmErGoNEugEYuVe62SaakeV3
qxFXA66JE7sMH4VtR1PaVAnuWqJVH1QshAex1lrAp4TSpHtZ18rddaLbJQ8El4tj
ayGhBspMQSsNR3oafKABzRX23ICNVrrBQa7w4s3uNeF8cdHeS3EZfn38xTcdGquG
rUNTgxnr8Ixa97DUeu8Vpo13t6wk2V7Rl/TCBC1431H7ynGdwEfoCazUtekZqinp
BSd9WZ9D7O7uaSc0obg6cxAX07RuNTXd/klvSC+2un6oFVNIwYmZ1FWFRVqtPvhe
r7K4TCIPupy8xLFvb57g73mxaMrxHJI3TwX5OGZ8r2Cun4RLjZ9DP1Auf/WhNtD9
8sKMhCjeo6c6S9dAkqW9B0P5grR2f+8/P7faFu115kCHYmOLVTMY9yWWkWsLMGrA
YKHT8qbhJ3c/lPu3brfpw1Oavga0sTp0c0SgIhu4cfhO0AK2Ylh1kD9R7Sj+8ClB
WpinUxDbs29PlhGxfpKGU8mdBIhkqYZI48AfJF6/G805gdGPYMz+Y9DxIvWKYuua
EpkBi6dziDpCQTnwGUQCSVkKOYxgb4NFyqq4ptgIRsCgeNYn4cpY5VmGk1J0OCGV
on30cjWnlukfUubrdBnWDlCgkUuS2MRT64t3wENTw8D8Dt6Vwc8ae8cnvJu/19HJ
n5wejOqqx42KWAt90CtiUyKyB1urhzKmr92Woakp+vja36hzw3wNv6+Gs74p3YMw
i+MzbaaMyyZ4MudHK/+l0+fyIRM4r+8axTWTdIfEgZ1ctEjr4GHWQOSr18l3Syxw
Ol06r0/mBc6ME5F7j1iIpsqYSVQ9MNy+Y3tEKOLapVv+5RVUY41UutsDhgJsDMfJ
1wUcSC1X/G2v7wb1jnne6Vg+IcANDfGk09mkadAJsqz0zjeTgurwl8OeWEstme4X
XTDUaSs2c55L7ixC76mzcgYKHOw52fBN5tmElfKZdpCz937cBZmKwtNJhTWkCb4J
VGZzjXS727JXqJLVL2juW+e1ywJAJeq/NXZsVTswnFYB7DCv5gRx0pWRC33pGXL+
Ju2bzb+3jeaTmzONODwJi27StzxJdv4yaTF84D7AiOLqxFm1aTTsgNJyHreogq/9
z3Te9IN/8wReGwlj3YAF6EBLhi3G8+LMrgOdiGLVfc8jLXtu2J2atwZxOtcHOjqV
5WNDj1HQk3lVkP/1CXVzHpV0uZTzp0WB5enUee1ARuTGHcdWwbNiWrrlZjAG2xw3
npPD2xW05rZS0ZBoxZa7ZjrK0+kxCSKHiA7XgQJ0qhQe4Zvc3SzYaASUZzl/GrRf
VlH37Xct37zm01C4L0xoI/ErwOSowtizwuXHZW44pQ4HJ8mpv88QTuqQKbTVODqu
9sUkobbOXyDQ6NIrpFZ5khIcahodhv6k/vln4lI5ngYPbFOXUanuqtg2ARGXM4Wk
7wHuImx5o/HhP0Rq/FWd4VS3hdTaq1ky+awIBERIin8F24mAuRUk1mjS28+6P0CM
41xzMRxPx/JkmCt2rn+sz8oiOR+m8TfiIe+bU5AxqvJfhx+dAP5abX6u2zzm/lx4
1O/8kEcIj3N9ch2D2jyRN44Bu1R0MNxNE7geTJHwFdsq4DGiTjMIwkBdpIB/Otar
/lNXNqI4wcARlMHZpb1g6w1n6tzIxABOEIJIlYZ8Wfazo8jjv8IhpBC9jqXdS2jh
6/G/w8ldvVU2MCtJcxn2UbpToSEgLR10HeIWMA8p4HpXrOzxuX2cVMj/G365r8rw
VG1EplwMY/jrDOJ+h8gSnnLlmKvWNajwolWtDu88Wth00XzOsytT/PhBdq7Nghe1
dWWqtqPc27+rPdRUE+e4Qr5+TPNT2klhRir60G15wTPpwSwMhe+Q3e1J0JTTEkes
4TJSc4uLKt/9iqv0PAYC2w5ta5QnIjg2TT63gkWWH4HMyR6Maw/uYbnlUxsOe+pq
l1u8pemEX1S5cje5dBRxV9V/gem/KQCAZpbHPB21uSmAPaPZqXeMCUDUekEdNMrS
q2KPu5hgGP/JQJznBsPR7goVoYbVCRbXsHgzKuyu90QweZdPdlrBjDgOz8cqZ0LA
iQ2gMeXoSJZi51XrWw5Tfx8WyyDCKDlrqHvHmVGDbOXrRoH5snCMQKjJ4pITMtpP
sMWpKLnqPol0S8XdqzJpxbn2sdc3HqkizwuR+4Iv5X8oj3CuRsySq14D/NxKwv7I
QBep+u+6T/qbkvTBZG5i8alKuAv+DM3HVps0SYF28NvO48PH51qxDfuOv/Zd//bH
F5qQHwqtjiaH1Llfc2my0+xfP8bPUKYUJ/LUIj8fstP1EzcskUYZJPWs/GIRm7ck
6kPTAuKR5MC0NUNLfkfEKpVrXUo6Y98NwNCu6Gnf4eCpNuzLyyah2KQGVvqD4F6R
K3m0eL2FaDdlL7AHQsZ7rRefFgyHfGYfiM/sSdMcWvrOZH8wkiHVkE44r9bFC0tZ
YoDtDjrvR18fQOeEg0yCeo0sHDPNMl682bgrH5wMFW4l0t30Ox9nEg0EGppRajzq
jUETddS4KV/CNgx6IksQWASxFA8wS5UzJq0kGUE4s/M4t4yuedKOSkD2Ht/ZEtsZ
6S4r8uW2z+BMS3yLIx+H8LODix+sDiOYj58SWRv9XxIREOg/NHxk0DYOD1BD0m7P
Z7lU48+mouTdCC14ZRKT90yLXO8csblSvDv16IWbTPnGT09idxFHAfRr9LpXtLgX
xL1ZFKhmoBo1cdhByCCbbfpOw3FcryLWkVwEIGbTOqQENcNiCyjO8ZMZqtr69FYZ
TNffXRAeZzlhwk4QvUT28kmN/ir7X9HEC7cIuoGUBRH4t/99EMOrjADKNkWwe6nR
Ds+UsX8bvY8s2IYtF+NNU58NiHy99NG+lyfOZw57PEtZ6hqyjGU+/nBnGBNjgU5n
7Xbq/3EU+LgcF6kJ31ltzALjFT6UVpxkFZ39lAbiQpX0SAHGPhUp5ecmV/KVB9Hp
W1rY2cWIflYWERZj3hRT/xEtModbZ9V8H4D5aajVf/W+hyaguwfGawaa0L8hv2Su
tup9t0xU1B3QLTKW+AfX1OFCBcRW1qs1fpA7iWSeQDvRcxSL7zl4lzrJdCBYxRxh
fmecQR+pOx6LMJmMSNydul9025wHyLQt47CsW8oMqI2hBplHE2GPOdyo2RFr5fum
lpI3D1PxXIJ9SvBb01lTwq4KsdiM+Vz+PuchcczDbENy91kK1YHUGOxkYIcQUMOv
ePS6L/W3boeAjWgLLAI5TGan6BzivzlPenuXeY+J2njz8+r46Dl5QYt4r5Wct+vd
z5+k49pNaAnS709xZN5tg9ZabfqLjIbxGs59Z0FFdbzRjkee5TQxvp0FdmqjHGwD
wlUwHnNWXCwFe7ciR9PJXDkZfY5vki4sdyYVR1k/BO6Anvhx+PWlT6vJeduP3nwF
Mndde5+A2HDMHXKmF0oE76NmAvzLNIinBEm+V/TDGlKUPwi1LgpWxbnY/UtcRrKC
e6kcPRA6BVxBsgruMJHN20ej/gxHLNHdE612NXMBp/t9XC3wiIcUztMSrLPWCZQ1
rQbMu5niQ8b23dtTTHsylmwdOjXq+izrgK0KOsXkalREUH57OKkbRKQeb939Khx0
k+fzB+/fixGP2i+eEhHlzXcZyJDAsC1IPx4UTVv9HmVzBBaTXKbGo71ZR7dcneOy
CP2BdJKW0wYTTvN/ylZAM262CKf4XB+V7+gsAa9/HHwooSSkk6KdaJccz7edDUl7
mBz4W1vjkG+69loTYmP0Yzjank+Jchfzn4Cxv1VZ4W8WjlRngE71ZchnZ4RsarAa
u9PeCv9aSTy0M1qMQzdfOnS3lMfHCDKglwvdIliX6V2msrGfHFzXJYKjl9RIfujC
06CtwhG8oCWF/1vXIvGyXlY2Dakd+M5aUQBqXkE8BalghDH3hrrcZbYNXjrenXem
dhoc0IEc+1OCH7DAhwvWM08rvgJpPBdGw3ndOiLupIlMwWZMFyp1p83zv/pqkWe9
OH9pf7LzHRQJDjCb6gW8cCcXtIMAb5XPFcacvsmdEpIca07cslmkXTA3QiG1frWG
4EA6IV6PeL15TeVuoaEEqjwf1HMguVgl/wE1xIEBcwbyUn/0weM++F6IahEhQZAf
Ks9fnNAMX8JiGU25R74DWHPNc2ARxaIXMOJXu2bhhxuWcgDg4IXH5KUyvisgQdA5
KRoaZeLg2vDvEIcJpIW7sJG+g9bcfvlNd2VUlt5AlGH9NT3edld56EH0B16VCDr9
TYDgZ5/GvDTHCTOzxDlA9N01d9q7RpiN4ChVYmxWk1Hr3pFdxO4y+/8ohGs9VdwQ
XFDMdAqOz+xiQddwcE1lEBMHwZuHDv0XqX6lU3B3XehL7nxJqOm2h34mUwFZnZm3
78K7WtujzTBMz3uzTS4n7VzWoV3/F/C0y8O3bBosot2rE4wjz/+kuxsFeAVTJ8jk
JlebnDkqUPYkQTqP5guf4yjZURxgggstrpEqJAP09pYFLp0wnjZIqPBUXBhf75M6
cDNrB8OSUeDtovlpNbZ6aZGaj0ZZ08WGIt9T2RQXW35OZI+CGoe0LWcyGeHcb8SX
OOiVbLCETNZLmjB7qS6x5P5WWIDjBot3V5AwUDNxks5qpkbko6/T2j/S2RTUpjeT
4Ykr/NCouWwRBLFiVdGk39OZLL7W2Q1s0q2+MaCRudh8yQfwKlij5XzU/BenvRVH
NmW23OXKmXPJX/52+angVWz1byDKurc0QsEQN7cgrYM1IPS+L8NFUoR/mmTKI09i
CErckZ3nt3oN0ooHx1qKBgNrhGTXvxih7/nNHy3uEmT5VrK7jhI1L4Uz3oBK4RaC
GbkDmOmRJjfubBmY6cfc4t3RITGB8APyWQvL714ZDIC7sJj0XR+SoIKk4J6+p4Tj
F1KgDtOd3Z8dChad1jvDaINJ3aAgkC0AjwIocdVj2kiYE2F6Ob7snESTmW7MAroR
vphvh4mOTaLXthxrtxRw1zfCSj3G7Ve74tDBirAX+JRrh/Bh3WdZX8cCYf+k1BH0
CS/CJofG5VTNJCAo5JTkk3tXFSnsQGvXLWvAJtKgI5QKZMgF38M5imqJzi7/dudS
lEGJl6MlKoGZ+BP/er021B9IqTOByCcohVVgGAQv2J27z753nOMgiIoZWeF0aCG7
9AivmkjCO1cxj+ERFbqy8d3MKEiw6XUzaTv2dyeon29au4tJjSzH6nsevSuyocxX
xop6GDEASN16KQiRaUD7457yPQ9EC5vjehjsMLZbaVfQeIgk45FE7CsB6v2pIuTC
KRu/7sm7VQkwrLt6DXMD3iIUulV1lGS6K67JZjRKcIas3WiB6QAwXHY3gdoI5cz/
UjKs43Cjz9/hnyY/XK+axFwuueN/+jCQzf1ph9zNEGtjrzWRbh0OqjrSpy70hdT3
INpthLenEoynmf71ugGJiERMcMS2MuC7d/empYDSBjxHEymBAWWHSBu1JwOMQku5
D7fXLHTcjWqknKIATxcOcY50u2U+IhGsma5kJuxaz6JDay9IugsYLJ6jJ7Wy1snY
bF67QrD1+esQrL18yzafGL4mwJ41zO5KCoqwrDZOlCHQ3opuUu8op16/7b5XCXBR
wcj/Zg/clnqDy3V7ZPXJsIvMBZysF++2P09h+VgfnTeke3+1qDUx/UaUbSesD4HR
uWKR7GROqdSJQ0gN2Lu6TSwCZN9+3OIo3F4IeWYjXBv40jfM+p5rS2YYFqRGr0Ta
C1Wc9jo17nKpuqOU+hjv92IFHSxEOKyzLOcLxVSiq3nh/R1yhbgQCD5BLVW2hZ+y
9HWWYarULFgnd9Nt1CZd8PeQqbql0B7u5Ym64KEFnz9SIQeYMtHplVBr3/LAcgev
5pVAkydDETRn7U/AxacHa7et5cUqDPy4M4k3AT/bC5Hs4m5W60TsOkCMA8v4Hmtb
v5xuU8VQLesOXUv3BLP3qivmnGJm9bQIjUwabwsSD/geoQjz4HbHjEQ9TTDsKrFd
EoDHBRd8chPZjdBAzX+jNJxFrHY/2TsSzSmkj06e7IPm10ueWTobBDUbq9Qk8+lY
WqUn/iEglnQGNcNS/DvS8AOQXq+1f4xVk8dW2qS5GkEpBXCkKtsazGIRXVsPxwsW
IEquvTKZrjQuK2s0zUC+A3bO4+g+Cy4qxKHPSm6uCRlIFOAKi5azDymLkvLz6/9Q
UheXUKJWBfDmt64Ozj3+87u6bO2ax7cwizvsAxCJdKkHxGmjadtwiA1IGBZ04QMo
GW+AdQpPf6r7u++rTUpKXtQDeOENnN8N1nEyRdOZcWRNf9FJJQIhGj69SlEJxzax
AsrTLzrz7PrdhUp9Zc7kJiWwID1T8zlSNjMiG7TubBw7asLIF/kuvZepeCIxfUff
QRcy5tyCaryWvbaaVT++2+ElAYqxVXOhMnnA7hcaxqDUQo96fe0WyAvyMQb+A0+t
J5W4HLn7Im2QU6tBpcWr5iPLn8IZ6QZrPFwFVOYKVChVGWeCBleejKV80RPEmnwO
Hg0rSkwVZg9ewcZrcAL/CjhanJKOAhBi8EPyvAGbNzg3UEizakbRVpCmi4nmy8Vc
Q0v3YEL1J5oKG4sS/joIGDPIPhtGLzey1t3DZxW+1y/exPOQJIftmf0DzMgK351B
rmwleCvDdc8iCpVICpljgeqZxhExzRuI1Qg5Af+Xy3HJFzHoSyPxwfTiCWMp+jNG
V5Bom6QoXviJ5mtTVFtog71QT173vcSrBQEfyWvk+jYvGCsGyO2uqiraZ5DvQK9T
oBOz4YVu6NZdUTpRmutw5UBcNT39VmsQv69kYFq0iJTBq4fZkzaZYxI42GoWnP0E
/CRxfnYG7pWMrlgodW7bx68ghtp2qI4xI9LEGBKWd9P21y4tEM8hscbQTUsppmx/
NGE17csE8s/3Zouo8tlod9ql8DfOikrQm0/GMTSEPJWOBv3uzZU2J0HhNF7Tih2q
mcZlvcIt04TJqYuQhqd4J2jGVuMr1xzhsCQ4BlKVvnEVQoZLlOsiQzxnBZ3bsmKx
2u4j8mlkMANUv//twU3aEo19pNDgwuhUBsOWt+aenD+5kn3CAvKPN7092/6Ep3yr
xZdGNBAybWTRI60Yf4xHZs5HoBHtrDBJ5CBvFpswUlRuuOeP2jNvor7EtJKkqMCr
dhIxacsG+MJ4xY+ssijUKlX6FtfdQsmhNV8EHrnEJfHfLh+Rp9MUJt7Nf9jV5W/1
oh5SeDXmU0mLXP60mXjuZon0hcJGYWCZPdMisgxhB/hMOkoJmEOVdyu0R9cjyHDn
Mpj1VWeRp4K+Lct1YJFTlZEySWigJbgMu3D5VgxYbycY3xanyIikha4GraoPtxCn
7IGJK3FpRZHfjHvSxRvi0eNHpnh/Qe4QXD7abhMimlg0DQueFX/AvD9oDGPSMBH+
zjgzO2QOKP9qQmd8YJA1DEe+vqD5O5jihKyhFQwUbZPsMtzbY4x0qaiw3WDcrbpe
dHB6U/Bq+SG4RgrEjQjpp2cNX0Cbe2ajiAIKOiQdkUftL1RRV4Fm8Z287G63AMwK
zdFZ+IzWoFo1uCtGo5Pb4QRH9xgGlZlSBATDIVK4BwVEMfRpouwlPdmKuznSTTtz
b8j4tl+fi/jqzvxr+W3Bbf/AVvnD4pNA/UgAAkk7aBnzfBhPrbJ++lcXRE6r3aW9
Wgru1lJcxEUmSShzjfSfCfyGQmrlJ3RMHANsAkdofZHnXTlZ+O6Oox+78P2p3dIl
44jyRzaZ13YA9WB2fgr0a+YP+szViO/6X4nLNcsZpYpx8xgKPJByRVXRLQ71BOPM
exEV4KMU2Y9ZOWEtHcY2SXur5yoWF7ob8+22NzcQeMUzsOqEaPwsjg0knHgXVLC4
C9LM4xwU68Dx9yk8vdSUzAXqf2gfc0b752iA5LfqTw4lNK5BAdHkkx++tMFF961i
SX/4HeLbsPMkA6IuBbliFuXNmCKXaltXEK8581fDP37v6YWVpBMOeTUZb/IciXL7
CzYdTVXy2/HYBmos0VWufgqafv3ddI4okj088Aq2gx3Clsd2EEKwUZguW4nXOh4L
n1oaGdVLn2V6yEi+u5IRxW8zxWCoztDetkTg758O0wNUanajA+3nOPn1rDi2QpbA
9ROu/pGQGT86ykRrAq8TP5VwCv4SQklouhdpBSotYLH1kyTRgKn7P0etehhA5heL
QiBwKDJog0/pSEaq1GVnUW8DnxpCLWEuQCQIjIU2DlxUn0J6cvKW6tsLu4zqn5rx
2dvYzzB12WeWp4hBjtUD5tcABLLkloiQPfkQa+R2lC6ID7sHPyscDufHYVePAf2l
KnZrsciaundoCWfH7MIs3CtG6lUbhLee7UpH6ma+eJXIxE8eVo6lC/w3IthOyK7f
f29tre1e5dNqKIYIJIlIK6jc9NzhUs6DJf+EybnWqOmmPB4y1M52BcZKm2oeYiJJ
ZgzMBurWGoHXXmgSRfcD8x7QnIfBuRhoJFTDik+SZc9IiW6A8XBeB1igSn9sLAVK
ufN8YlL2eocFN/LLGn64GNnOvyI0o6omZ4m+FDRy6/1BqPozJt+Moxx6yAk6GCwh
N5H7tyQi9InMG7O7YffvUPRMTlkkyN1/exao9XLqWIHyimCF5fBKje8cvuPOGScF
JX1vBWLiS3BIVrq3OTt2sU7DCqSzwKbLlUm07ZQpDgTabrZsLDMEqb6vUhQcySIj
nzSrjbFei4bWpTQBOiG0M5kgnOv8BZTgmp7DocZM/9/Vrf/+H/+v+Hj6XKXBuIur
dExSygSx5FX4maML0j+yowhID5RKnL7KPeKYhaLHxslWGP3cC9Yk5rBPFf66hPSt
KsVmdIX4axPTrWELjyJnUaz+er7PH+OVi2YLjDw+DVc0zhNJkUjxmYNZrW3zzMGg
eXvx6EmNYd/BVvKbaIytrX48TNf3BqfTR+H18GfOcZVZcE22g5PRejZldL9AbWzj
E0AteHGqtgzkLSQl+nQCrATA1scgxsHKGYQyHg4H3EOv8TkMZUEMkLUuEP/eKWUC
5FPQhSqc4x2eu9ZuMvvzq6zbJuv7bQ0ovnhxaiUuPYx84mE2nYGvceFip2ct5IjF
C3Js7fgsXNxzbgnbvqpLbFMQYs5FOHEG+eWvUzjc2xSw7FqKY0ymn+lTt6cymrTP
8HnzHDcZWFyIKa7FOnBTSC412KROlwLOerOI5wL+PTSu+/VLx/xNwpI7tWllbOLj
okIrceFBqIevnAeLUq1P3i7qk1sISt9O+1nssUI6h2UdH8+zAU86POOQ/7FvcRoo
vFZaDswqYjslC1yYaAAptX83z+YDirwv92Q2g+noePm8c4Xr8HKCH3j7TNaxHZMv
I73p8xoW4ffoQ2ISAZFOXOpuZxa1Asc37CswIc0I3k/fqBGytuHwAWzoZj+Iqb6u
uVm38SZDktR+zTnrjh/WscHStpzOb3hAznfy6iNsTIW02UwV3WcBHvBzykcQSo9C
lKit8JsJ/3US96xgWHQyspFVXKogLULM3PrEVeHSwcUZYvkcJ4xF4Wule6npD19f
n4mccUNpkyr6CGxXDQvMfx9WwUXYhrAAiaxhxaEIEpHCNHcyFpDs3chaQcgKGWiX
rlZHwcHavapzjGF7qI/nNtLSJd3+IHgBMTZynNiPtbYcxWFz+bJtzEF96MZZ21nh
cF5bALe9fqyYPv1lsKQTrIBg6RBvV1WODC1odQUaYZz1GGGrRgZKZPZ9kTzwcQQC
UHDVnQ4gGgxPX7W7bGFHD1AcRnb5PHE8hfmCSxTL4/tXSkEBNdrdFflc054LTzPB
Bb6D5D5GJHbcyw/RE047zIi8pqxU2mX3eKQ8AxQQXk5NhY8H4d32XPDAPpg+usfW
oGZ/0kEE+/d1Hfmu1WbkLStST5ZVno81p062VRUwp8zlFNZEYYtB47iOaBykqgPf
0FpQQSpP3kZktTg20J7CKFcS4XjATwK3V0QQsFkRnTc5lkMi39sWgMlkNUszFeQq
JIiEX/otudY7/505HXX+zg1GktebzYmQ55ZCv/NFE2Xe+i3rQ+YnS969fNrPM1ON
p96JgiQgG7WnITQC1V5/XdfVHnAxCkpr6Netn86So+iqZA5TuanJXeJdCjaY3ZjB
uoVdXf6eySTw3A4soYSWFAQ7UwS7kPa8DqK3/FY4m9aNOMBCwP0qjyezReQ+aMUs
cIVm1380d46evp8NVviG4qsZVOzubWzTFYOzFcOZS5oswOqWR7/e3/VdIJwd7dOd
Q2kP557BdR0v3MEA2iBYCkGT3B+zoyix1XSOAf1116qRkbF2gDcSGFuagRjBPIzo
tIWIMpKUiMTwXA5dQhrzzToagS2u/ye/n/qfcjCCvSTlMRqeQlLLJFXzFNz8bH0c
jhnP6r7tiZ3nBMZjtdR3IQ5wbRB+1ldp49LZ0klCExWj65GewwT9CNYaRx4aoKvt
305X2OT4kktrBy1xg8ksVSMoeespDU12mKOr9Qv7SYYvZRuXsDaJourxvUygzN97
M2SHU+VjMGok7TzjEAxoXDAhH0WyQuV4B5ZvnsCqlL9lpItGi+IFQ/BZGrprvGR7
p5+SlYbOOAycPAjgKQ9sOemBSurDU5N/67Ocs9hTFpYH5x0QL4t/pBr46fv+//hs
QTHWo4z7E+DzvG+6BDtqixW+AEytG3upQy/lLK7Qe5hHuNqp1gPbUt+0i9HqPlzS
lxMExbSFh1ODJNGdGbIJ3JmB00Zh7Plq+e2EtcbyTNCCUCNmRG5j82gkZsUaExLS
kvTZVTBL8ruLTfWCJqfRRdePZde0vqR3ml6sWOk1IKa8ywhr+JXuG5I3Fd7zg5L8
5OQNarmwo5aoIEMbX9XR2lSZf7bGCkBY/45/wJ1Ok3yhwDIm8/4+i8XfV6ddH5DF
mXiggzkAHGqMoCr39E9c8R4AR69e0duqYfcH/m2FyXKBejoC/uvo1M1hTV+uifE4
4+8Lj1ky4nsEmtbss67bZwCcodsFRVAfEB8Up0u4ydnUOHjjCFjpiIiDfkqjbL5L
iTjQh0M0AYj0yudFb1cCdweKT0H4Zgevn6ipUbYVD7RTWlSmCRz+3X4NFYQKlzwU
Wh6xEOk7Mx8igi+/YQzv2Z+G47QBrvfpBamRdv5Fs8XOms21/ckngrkoVvMUTjfW
m7mTdTjyODQmo2d/OQ9BkX8H0em52CTdRjU0r4tCMJRhYfgkVcDvwm/yPehr0nyH
L47nqHnSc2FwliLKrcbjYeNKrx1Ohk3FHifg499OkKgth1fWG1NF0l/Bh5D2+J5N
EaGNpH9M5+gqFf19UfnyEw9kcP/jEMZ8jQSBbX6qTXaNx9/1MuzM0JEDIn8RHrgI
d9bAcOCc7Iio6mu4SQX5YvYhur2PiZXRhtZqw2jhIc/JFdzPuVRTwO3wRnTTh1C7
JftopwRDAPGqR13LdYIhu+9hfOwJ4NtneeN8FCe5qPRk58QdnmRfK+c3ar4NnsXD
cka1EbYg7D0Psv/dssx2bXiNURTcV40VOvuCviXcQvtoSikRjba2rXFD4hkpcXaU
f8ntV83uPiXCEaNzpcqX+q9cBs4jZclJl7JUsQTQSzGnBnPTOXOzbnhXSMV1Ali+
OXl3j9Tm5ABPwvq0r0gZczWoumFyehhs6hVa5B9mDUqhY1SmvgO2Vpsef36HRgIO
/L5TUGSWZsIc2c6fKaqTnfiHNJB4yJKnNEMu7DHTMmGZ5ZDTOjLH9D4vEyuHzkCl
u7q4yxe6H5r6SPJI9LvWbfQ0VTuQQyp5zymUZFEcPTQxg6731xTorzS81ZHDJvQ8
6NLKyxaI+IfWg/tSYXD8eAFuegZMAHGwVNnGLKq0hYu1vSDASqk8xOVQuOs4AtNe
mT0CopsVxUx1jhHciTTSGnS9xp3fPQ0Tswx8Cp4DE6IF9q2ffoAndU6Ah3r+NR5E
RQtSyA6aWcqHdSmWwkVbttJ9vlCAQabQL6MY/eicqBG3ZA9sWWZP4w9U5e16Vzpj
agZBWxLfSWb0jjAfaRR61l39wwKNyZq7GdTDRTYgXWT4bsOvOB35lLg2QMjrmlA4
oFQkOFAC+1N2i+BuRCLdknl3cJWSMnoD20M3Dk6mIhrdTN0V3BCcUAOSOezU7BjD
iNlmejY6MUuPS59S9AySPG3jnwgVFVfaa2mn45/cRRJZT9+KBbbB6RIHRurtMXK3
nq0KdtgRL90VK3QlGN/SVqeE9chGqKBNtvQeJB6nNmIOIHNdYkBBVYX8AhY0ZyB/
2Gu88gKl2ejk6/7BqQwESPlivXAAcctieh8cv/QPeqXUyEHHlUs5mBu1Z4B/LOwi
30K3Kx97Vl029QSZfHMxrr5gN7c8JlsDQWZZ2CE9yNTjSil1NwIOwfciWUX82Y7u
fO+8fXib4/rUjncgi2Ljuzsu5ZygqS7K5Nq7l/7gjuei3w2qDTFDQTBCi/k4Q1mf
Za0RkNgT4pqiKG0V+TKCoWquQWjRqIQOnzJCKIhAQEKnbd5jFOpsL86kAUOQYAtB
PipvAAo8wDEKhLlxCuwKoZNDZUqBbWiVqqmPaqVmPeVyco/SduM3w1djzc52Zy4E
LdQVamqXQtRQEH1ZCH/K2TB+Rr+j8jucTqjNL5gCG7Ce/UNDZe9SUAczOE6xbYw5
VHYtYN8LnL8gWdbCC4EEZnN7sGXYHOvdUeP+LT1YcCwwtGsQwvANBGqvvfVFLYW6
yC52X1JbJoCg9JU7q47JC4HP0Q/UdG7x1smX/mLbIJoh+7+XbakYGpOak7ISIxHf
t9VRoyjQ1EIb1CWyXylVtbNeOgF/esR330H4bXfPSeVGpw3fPbmfgWj7RfjWtqFG
nMKJGth8zHpOff/+0xjShUXyH5roA3Qof+HZdrLU/wFpqbS/jSDHA1CWDLLbqn+T
aG3CKKQNMEqnX0PVZnhq/vbG7cVIHa6nXjHTmiDFKmDdmhnefz01qDyi583YPJOQ
XwdWcn1+i2M4pEGVIcUZmyMKavyxEnhDYNQtzkw8msnK2SVywJgdS/g37Azh/beo
EX0Q8nLNTiPz37z36XBDsy7VtMceuMK1u+Lt1/8RO9DOTFstRxlxhB3PzTJBuc7O
7MYhDc6QK+SbD35qlADwFeX3vj/aSRDU4ToSPPP2rgYm3m89sW1E6wXLWNdE1WRh
anjEq8wpKpJTkfeh4ms4QPulRoFUu/7N85II7YuQd+LS8E6YJk+siwseKgCeFIEH
vI2DqZPFYBVygK0C3tz/qErqRa0Sphbrxu5bJ/Gh5RbMEcCJ2ZhwkW0ya92cfWqG
DiTqj56OIdMfLfeaw14Nmd7IBrDosdSMPxfwRLxrx2m6tSetkPZxQVpUhyU6uLQx
B9TSNIslyBfXVDb3wO0QF3W4zrFt/BZD+oXoE4fVDQAHwL+83Hdejqs27PTLSw5v
LCyFs52ItWdOIkdc7RGIwb57tmipyYME8bwm+OMS6WoHCD0sgtBZW3Rsj7PXlBiU
eOu0gdhfM/dKIEjmp/BehpZoBDdPE8U11jidhnVI07UR1aCx5OW4z7mVRVq7VyWD
0BIEzndmY8jvQretdP1zbwTpI4D/Ocf3gr6vjjpV/DyNl5MFs+O6JoRPis8AYuIV
v+/O/Gh7efERePqYWDriRhEvM70ARQDvr5fNfn6l7VAc4G1s1b9HCfgD5dXIKH+z
ecFhFXYWHS7AKkYejOrH+zNiPgfHJy9MWnfdcoF9YYDJyZBkvgkx0HRsPEW8x44Q
59vq+elPuwkw2hP4gGfqeEZg5EgOz2x8xRKeU1VWfb926Gg1xOdoyuHL7JH7TqZX
F+IM/Od09KxxMH4zU+rhPYG9P5g3PbycRvTzf4NCmcPdJm1a96DA8nfJ0GBgBmSl
yOOxK7xO3KR20bZ+j+Gdcqnp/aglJAFd2C6hZmys0c5xYvsQvP4wm1pBPARmlLtm
RrADCT3AyrPjnXueYZdU6PM0YVJgJYp3D6TqdLYL/MuYc83+m9v59S6a08dcgo0h
fgDRkycyqOuOBd/6plPOD3AIxyhyIvaNY1wD9vrzYHobdItOT/H5vaF+tfy05TPV
Ww2vjqZJWcxi7PQstG2puwJxXciNfDZZWmPyUfvSxBJFvVSAPU+DO3sdI52tkVbV
sha93dnYFunD4bEIBVZRYaYHzFnaHMUfg3rUCRpILasYXbCRPB6FxbAQs8y+mWoV
X+fGKAPso3JBavATpszt1DnHbbWOwnCEk4awMW5DxRTOv/XzvYF1WdlTGnMP5b9R
Kv08+r6oeOFDeJBqBw0649LLQGs3enXzLt5a4VDA/pAb1jMbg1TjpUdER2/X0rCi
P/5X3oI+RvHJk4s8xqDvRXg5s5G9pX9Ygs11G01xtfV2vD4gp77T5d+zSjFnvPLy
BJRfWroDCaaQnyMzciOChu41mZNAwUc6HNiFGGwfY9cvtb1KLqL2Eud6sebcjO0n
Iy3rRxz5sC1fLYuJ1Ov7C1JS0o2k2s647aFyz6tMxzIKd6qdekbGSqgj+O5iaqyG
itcVKVvbsaBefb8NOCGU691aQLUL6jRFTCE1BAnzAfIBNxl5bNUSkBwummmQz9ma
P/rJRjyHzcqVxOKhYcxdNDB+ocdYoG9L6l3Mklba1f4h1NRBvyh8QNH4uWFNf8xR
NFie9rWNwFlP2z7y79YmVty9WLtsbIe+vKMxRJVAQyQ801cGKsQ70KPVqzPyatsH
JfABwgT9jAvPqPv3Mz8CigdGjtReaaT4ARbH3SUIpe28VYWscR0RQsFv5XZBDra+
NybQGbE6ADrhF6zwfkj0d9y2GhbNlWxXsR09nK/9HhsoNvaxEJ22g8lUirCZX9V1
LHQLJTdlCJCUDCwGS/smCk4V6FeM48xCtUeURzN/RUFipXm7F6fHZJlKt0CqNbCM
ZhSZGACGWiZtUJZWdsrQcPOH84HIwU3JX8fh7/y8nYGl4VvsgtqMQkKQYO3bnPI1
/HbDKHKRsMufJ0a132NmFOK8qPA/MTefO6fEjKE9VQytlETpm+cR/TlF/EVTjuVe
nNJw8+ELKRALBKumWXD08PAMr/FdC3DYvMTJajIxrvmQHp6tGrgmaYdTkMP/XaoC
tHekAw7+SkKI7XjAf+72UAh4jr/fMTcy0CDVBw0ovAxsJQQAmtI70Jw1WsVtrn+1
YoaZCiBZOe/YTRo0BSk0YjywQg+eMxXe1m/N0Zw2xVEjlQGo2/U9Ig+34Q3XMqPR
euzk8B4IgKTGdp5VFLV76xAXBwveZcZCkKAx4beUsKWFD+/pdxxq/HnX44wtGiFk
YpJ9cw1ObdeP/ximZwyAdlmP2vz9Yq6c/9dlEt76EWfUloUKZSIzmVUqeeEkKzyd
wnprjQCFLMd41CPmH5tYw8RowfL0WEaIKFCLcR0r0EkV6UY97AkAzwVcxjNic2MD
gbgX5vQuN9fjPaQkqhIicpSf2dkg9OcAiTA4i8H0CBSqGxSfuCPN2zJ6ayrpvZCT
OfouBv0Y4D/JhNYXDvwNmP0z1KvJNXbF45/kpNVpOmv+eQINx3frf8UkxKY02XkX
HhaUkxiZ2h8P+P+u74Hx8O1en0yE1VcTQPUQ1ztWCYXgj0BG5CCRwNdR+XxjjzV/
SXs4i/G1IE/Jsjv+wQHSBsXhjEw/LRbLlWFH6bqBgQ3L3ancHLvqdBIf4Y5lL7BO
ap6Pm0xM+ZygLxMIKXDI1aUL3kC9BFEdWH6b203TqU4Z4iee5lmYeq0E/zn+KP6q
tsft/EDf5JLsPtQeH0JXppIW5rEtk0NqruHv9mp7YgGzsmsc3hfgbgUW3NhfDEvL
RFN9zHbVddYsgNgop4GaeJN+gnuMCL1Fevaa6UxRkefdZ5+AsVWCbi5xhZbpPyFR
Z4yUrOF2ssTR2C7766s+AmdtHIGO0n+cInXDt6J6WFfqWQZGEXboSqqsgME4aPn8
2EfyL82Eb1e4rjdzwJR0OP7k939vvDtvB19ihyN5kdZY3hhj9OHGxJELPh5IHiuy
yZScx13l9CrXjkijhAScMsnoq+nPYMGeTFNRZsxY6AHcErAO0McsrTY3wtXoUPpd
xmqQ5cUqOwK2K8T+sO5m0MkP4QKsm/PqSVRs+Rf97sI52quCyw1p2t1isMcYXgd1
o8dxBFqaJViGJMiiwk+1Hsn5SEQ/8PyUgw4v2jIfTup8lZdCoPq75haGgxoD2tIl
gskWrYzbDLzTUyg2IUF0nDyBmm7CJn4pMiTxkzZhk0urSKycUZZpJwaia9ko0z3T
hborYPiPi5OQEKVxqCbH2C//V6k9VExF39Y0Gd4V2xRQlD1d9DbupqJWmd3wiyrL
Zkm/5FWnLAqNwTHfOi6En8qIvELMPzK25vFjtgb8pKiU3aZcVHwRs3O2pf5GZpYa
o7JTv0aBU4x62MT1Fqlwq2IgIVNyFRNc0pGvW+hyUh59yNk+YEvThDMq8wgG+7PD
INEUK8kqxx6EKeu5pOUTX1OmYbpXTjQnHwZxbf42p8Jyu9B6lTsd5Y9HNrZgfmTw
dlSEtp47Z8HF/VDBP7mrXkmv7d8sfL6wF1do4J39sNSfwv+JBdg80TdCOi18/q0V
zllPnFE/Y1cTquER1ynzqdf36E2d1DdkphI/pUkBOgThZIjUaBJSj6q6mb2rCf4S
n9e061RD8h6rMKGxDnDBFQC3p6s0ctrK+gQ0zRYoc71Bi4Kj/ibjYHXS8e6kQC/j
4bZxh6IQun8zBtQRX0+OqgemXBEL06TViNU+VujRST67nAZpxSmuGaR4SLl/H0sq
nKng0rtcqA0VUjqkMsPof/BO2RLVvAGUVfiXdfMIgDhmwSkDsVhTi3QXw2229E7I
ultw5g6XHHWeu4larVy/iYKoH6Uzc2cMFDtOZUI97l62Csj5JOyWPCdZa82fZp4p
gkHxfUxJP5CtP3yeinq1ufl1QHbRyUkUeD2oDsGGCdDvYMg0o9V3obEE7Dvc7Gx7
EFxZDWbtzSd9U+PjQ0pRDjG+7fgUk2srQN6La7KA4BTABMwD5reNomuX0R0JIbs8
VmhqEo2S+STc0ACbFj9DXU87Z0ftgJyC1EhzT/t5W95HpVyq+htzw8n65NcttIQA
W2aDSVvD83tIhjUUaOfur/yZV5aPsCuVMvlHOAbKOOh23pLSnXYCl7G786vq/RIx
+bwgmnH8RnWIeoR6v+td3V/9GCh7A7LsDlD5Pv7mW8IgxeP+s/S1UCqDvCxTV7ml
yp74UK81Iu0l9sZ2uU4GnF7XGisQA1XaA9l+iMlkoL0MDHBnkBLNPLLOGElCKdUZ
EdX24uyTU3d0SYqJ/+G+XxoE9insmbC071AQCTWYHtVrfJZeSQQSpm5ndbHCtWhq
Pe+cgZPfSJNz0ZOI6QCTbLcd5T3dANXMLMqD55kNLfkjyuRrLufScb7esmvJ9x7L
k+RvbFIq40lPsz3cSeCEbbZojBWP1OKzpiJ07Yiq0bCx38DQRT8UvkiFF/X0yVO0
ZUjEV7TMjUcM3P42SZJj8rgsac08IZUaNHfmJ5B+Zt5ZT2ymxvhPLwdRDepGei2h
WWU3DFRf90tSzTvRgkjG2TXRIwxQNNiNvIt10vd6/2DnF2eMXjiXnwOHd6ker8kT
XYr9VK6G6kbrWCqs/H30qD+ZqvDEEmpP5uZTa2xQ3gVVKqEIaX3O4YJ2b/6CSQ2e
eQfmN9TESUCLvK8PhSU83T+jgaOtB8PShHRiWZj1FSkL/TSbBRThDAlICmP5qk70
X07J4eZL04j7pMKPk7n1x7IxAL4WbK2b7xxYKn7e4JXqbkiNNgr9G43MkwfEpRFP
trvdishMaRkZxgHAV77d6g7V2cuTlcN9srgSajtefpaUJx+qJJE09+liQNVd95j4
82Bgxgs/FdIl6uGjZtAH6EWcz0UrNejwiDOsmZ/lBrEpxcAEUEUK82aU1re2sxqK
hnUKkE8sHWme51lSsfXXU5mO5M4r0KuIdOGBf4ZUK1vntJk0syJ0DuVF1cKtPudT
mZqVkRWafOYkDZSVY24x5rQg0nVd+8S6ixWAHDWwAHFgpmWwBHUTirSvFleVpm40
iN3tPN0J9M6vEPnHqrexWXDYKczyo3yi7562qSCXhjRwFP1RAyrj7fSnX7tKwyee
5B4dnNptfElrt+yqFEh4iAimOl0M+vXImXargz4Cl521zofWcwuDdkoSYFr43hRk
UukHVlhHTw66IzvBuxzAGqOAkuS5BUwYoJHKEGHFTG+/EMwmw+2pJEVXI1hnkAtL
3iDMnfd5FTTCjJ7eN3UG8mDfREhReEsIalPUFTCYt4Xm6iOSP2ajX5GZv8Cl5jeu
18NR32R0RDKQgRUMlxWyb5YrtBxq+sXO1zBhn+IBpmNxxEO+vgNK33ocsaepu4+V
UsFJ+x+oca1RMzgswuyuQIzLKqcbHitA4YEhvjdWY+PWTXYdntxicxPLdoGWnjk7
chwZeeJE9ZJ0POFJIrumrN5Cr3y6sHnHG2op33sc3V8gz11JScCynj8ePNdUaefN
T6l4+eRWrVSk+8nmbW9Ogi7HvhyK/84ulhvMHRyHjY8FeTzc/JQQ1Ud6TxkZHEwI
bPKKmePI+dqLcYg+HOZArc2XfQqGa6lTw6NKdskB/gJOLTqvFDpfTTCIY6Rh6ZeY
Y0LPdlUPUGdl/5EA0LvJdxcL7b8HmFUC9VZQZfxHXqTtud2CaPFzDMxR3IeCiU8F
nuFFwfIbWpcafTYDNMEvXpGWVQFyr6zTDf0qrVWIJFMUgQBGqgd3uT9QHprSSLBX
/y96cdeeNEnm4mHLKJYJwCfztEXtPxGb+zAcD1YeX5NkdkHkw8HTGJHh6Ica2SAS
m8///1HhRD8rw/ztIoogZ4v2kSxDjTgAzYeO3rsyBQvBCXBWjV5BdjpsYJlABLwE
Kz3fwxPd6KalJUQVI4zJSOy4lp4XBUGaVp1eI6xZZBaY6w4MMsoPRKp/y85iaj3e
bxNnAB8lZ4mbkQoe4ii7AaHjsoKFVQBSFHCVd63kZvFbbbx5nCeaNcG+ROOyEs7Z
MhkghAqBuOUVrCsAzkiAgw/+pg7meolErYoS9x/IKovK/cSzcpL8h5C0mHDEUly1
DFUQsi+VhIOQ0PGxz6YPlb39rev+/Mk0s5RzetNZELWnJ6BZ5OR7bPD7eOHKjWT7
77a0zvkaF9eZR67cHo7Xnpj7VWoOWjxxRu0mS6kQKeT+AFNZ2ai+jORXxVIhVCkt
JnyOpZxAPi1inN3Wj6M5yGioTNIiQQlMy+Kr9F6a2EjPXUNrmglyv0NSVciCgjp1
1/wFkXBAbh3Fq2nMJST1xweJV35vd03qgbVWb8jU4DJ1xioF8MMFtOBL40VjOVOJ
than3msSsQHd+KQMakjVsydsZjBO0hbBqdulryETh/LWQMgB3Ti/mPW6Gjfp/4N/
5ZVwuAmO3OguLSpppX+Phc9HIzwME98KBZWfpS6CtkFLJ8vR6Vq8KSvqOuZnDdt+
97g3KIX/adLxVUoAG0ocgcRGUNM7jXRRRL7WfyaEn9YrQPYNczScmrETW6gvmEh8
gVsXlfYq/VTvgy7roVOhJIJ0GFUGgGORvd76iARxe81dITuzkhqB2n+bLeWGGUcu
1nvlw2MP9N2ALJK+CWrbNlcTZwckPK3ux1TEbYlWD9NEMxowU/pcTyE2kUp8ldPy
SCjeiRY310Zh8gG6TTydKeUV/1NBV7SzD9XFwl+VTWHZsJ9eWOOCxyLixJBpk0RU
e/6kIl5yBQRRdFh97szVPW/ylzKS99nzz/QrPkkrHgs/GCt/+0Xn17JKRd2k9KEw
b4eCyR3+iM+VM7FBKmRLhUKEytq0fvqoHvMU4msHrRLm3mstX289XnqjKdSIjPQY
XpYshYyV5pUf6aT0zqEmmuf/p7Yv6zirtzXq+Yu6PXM0fELFe/NIk5pggRZGfS3V
Qd2zdMc9kYXhGv5c8kplxb7z6F5VLCFRXUDq6x0SxdVcXiESaIH0dJwgZLmOT4oO
M/8g9uDhoIAca5wJtLi/J3/A8nB6+wC371yvO2AqIqi+4cQWMCA2qPzDrsGWBMcK
8HKB/+L6W+38Zy6S5bzZgwgLjt2fC1UTHuOHvDhTEHVAkYYNZnOC6gaByJ6f6NJX
Mn1eIZziBJCcTvl867NqQBJlzQOCRO8s0tjsFCG5/boRPbCqqMCIT9x78IhbMvcg
nPazJbakBLoZlOPrW0g5hOOTpiHsz8k3H/Sdm5BzJjefDWK37yKKPd67q0IpfCPr
0VmPZf4dx+KwyC18ORVCAbwd7exBtYFKxNpRUJ6l0Gc7wm6JBFj0Lu0h9HbPlsF+
y5w9UbuzNxRR0SD2Z5DjezPa5/hG0yxHro/nyMCluSL/E2CQP5+Tac8K8JqX5YBQ
BIvnnXP73qtSdVfD5cyhpO8/yJ/vR7H0PgvUlzi8mEmo0RBqFmb+uwhjuKVpW6+h
25mirFZf95sYrkWhOfSux2ZCHOTzJ74qnJoiV40XQPH/vvEAb6YixOgxuCIrDlyX
BYuMAIywzzlL8nt0T4zxx9vCqvAjHkJgt9Cslr1+Q6XNKyKBkrG9gTu+V1hWTqf9
2z09y3g5aO5l7FuhylCI/eiEtytkfaPGu/C+4hsMxS9OL1zXPwwIIlzdXJmECMZ+
Av5eKLh/g+vgngZ5+VTFJ2/iD9yn6IlHZj4lByFoceMvOsLYorZIiSiuMmV5a5pK
7DUf2EUOlib5az2RcDtAoO+7Kr1tEDdWEFYvLgNRuah0OECXrGBtuYCk1/+VVLs9
NbkJdYlMV+4BdY3/J5Z2LpNjsCYx0zPVLg8B4/+s4+w3rpFRPVjvqGFOmpyNGIgQ
xqF0Gjxoygyq4JckTungOgoUjKPEUrl8/1FpcN2dCCndRNDOb6N22LBafE68mGm2
wZe/9x/lyWxBHyq3ewp3cPC7tP5wE29TPsyVrdJbD3lDMuV5ed4RlqX0ywPGy9sL
a7vS9ATc2DbZF69EyQAI7L714Nh3Zr5GUa4IYyspIDFQrY7/bOq7yBOpoSGe6hWA
K0sbtOIC6eszphxiBt6IYmDq6z1VcaZ0ebNQefuVBk9etbH96I/J1hcY7u0Vo6w3
DftNPeGdctYza5qgTaElfzgmkf6+XCfzbD9ACheYRvbAW+c14cTaxfUBwjojCfO/
KXBwTPlBRROSauLkF/MbOd+sNNfeLyKAMkSJsdM6aDp+Qjm04nmCZiUVVRAXSPs7
+bjHvCSxix42/UwE4g/2++4geQB/vygt1LvY2Dz5J9QNBIpbE6MR5HfW7ihh0zoe
u1ErnBwANWpfVbZCCG8dDNQUWaPOWkNrTT2HuvWDePaewG0Yn7fDWgdzhCItSFmr
x50z18l56nvpD/D9uarVaVBObxn/Ca/vDMeLSpGdTr6XfrjolcFuCRJNl6is2XVo
Jdoe1U+CJqdtAtzcyJBV4yIuFy9NwkR96BgMMI8THEQGrMAldmL4RjkI94P+1zmT
s646bWQqjdhlvmM88K04fweH3jAHtqH+ANZA7PxYv4XEu2R+XvZVkXL5wrfCcXql
KaHJcUs/h1dKcfn784vlXn2EsDLRGVIJUigJ7EEi+n8FxzwCGnUuszhEDutKZhY9
GZ/HV9lruyEc/IdHXIZzzoWr1h0JINLwoWKAZP11cuvObkKXIF0n8ou6fmUTTADE
KD4Ipnh8AIPCoiM6tAaw2ImExJjCD3CYnn9/5by+zYYQ1qC50p+qVtfrw2OIwgFH
jNh5ho7MD6yFzT9/4CgNFIzf+UYtrW/Blg7dBbGK5Jmm74eoqpjf0ZkKOQglwGV5
RbC8dXI6PvAIR7FK92id5jluWyTxixTqr4eZ5MwUgF1pDxutxIyyJC+0HLzyMtXg
6F1t0vYUwswnIZBTYGHVdPH1A+9f+lMCOT64KaX14+KyKE66vXovmHNYfW4yildZ
Ux0XbAdAMs2qWneBhjgzjl33stShL8ss0btIK9ptuT6AIIx64N4wAbPwaftKJIIx
acnj1Eo73ynpE0nHy1cDKeWcMjxq1f9ckOxqFCng/o4as809TmQvecbD+3eSc8EP
E6NsZaRKtr8Tq09tVopquOmkoQXCpy+DeU4b1O+Oj9gmNePtRAr61m1B8k6t6qFt
Mf+CZqTHS57L8+HwqqpppQUpnHYjlB3MwJLzKYCBlu4KRxaLI2fH/FuLouwdKIcc
jaK8dpKFpkICx+smrF3Ho5H+W+hh6N4YkNBhfFhkCitTPb1qBn7OGBH6R+KHTcAZ
eOtLpSo5yJrDPfFrZIcd92qJ7JZ8em0GIZbPa9boS4S4stD3Pe0Ek2f+WFktid/s
xc0iaJRgkfJZFvN7HOv2f1f9PLExeTmql5yxRicTneuSxkwDmjoyXmWUptSjfCqQ
QQVQ68G3zymohv6+vtolNYYx6NzpGCABb1cdr6GoAPMurabJaelfXBKcaBW1zAmD
nqe6D/b+9jleZfiZkug+ZeMCMRNEZ8qm6NOIfPFwEZUhcJc0EgVELSGt8prI8agk
2goETui9h5NwDW1pIxen0vgXdnexXlwRoPL1pqqztSsjma+4WqRrHFPHTmMqjOio
0R4A/yxRw23xzzE6HYNKjFaHbYe9pCAgXik2xRyDL3hcCY144BMSkPMbPGPbXcql
ic9cyU/ptMnkTyra1YQ6cOHeDscLETUlPRuIfjS32rF8E5hP9Mj46VzFiOo+Cr2P
00zDhbjS26Gv5KSf6W6o1plTjkda/e1dEKUVown7XX2OEEEn/4lV/4gdjyjlZdwr
YrwHJYe8vbC7vgR12Y/TPA5oxuxqoS+OLGBxyAEOd3gO34z/jxfrqGrHWZ8ZtSXT
VYp6Xf96d/ZdCN2IBzRTsEDPFSraCsoAWMK9jGBqPTctQdSn8eCgN1KF5Am7VCYW
Y3L6SrZ9rTGSQ7yGianUfeuqUYYoUQRV31BglPKMmr4bvO2c17/ZyN7SgYLw9sXG
LVP3oxY+KYeTpLsQi6Q9xBRzt7MmsgWyX5SofBiFuV/HjxZQ/3n3W8f4WD1y6pIu
B0xQbtdw9dDOTPeMBNY8mN4CAFWkUNymFG4Tka57NWm8uvM7SrH7u2IOPwla0Zia
CHsKJhVoAhFzBjb3S7QyAQeGXTPpPC//adfD+t3tGXV21J4k4igirSoZfT61mB4J
0UisX+SsTLSx6UFr6sT1vJSWEQ5ueXeoUpjEgUoxTNEcWcJmvdfBJZk29YrT7qe1
yLiHAt979/hnULDOSsB6O6MkTem+QZAKPs0mlFsGY3qiuUlaV5wdL2htT0iOrDNU
A5QJWKHzHQ7N57SGaz4rMDtzDxlxWVsFZbbRhP/APbnSefUJZXhKxw/SIvvGFnB7
dmtQQtqgCUy3AyGjDyqJTssjVBimCbyO+3yiTiRXBr2B4Uf3jjFXvDEpPP8N8bFI
Qy5NEtzeAamOo0yq/aYcZS/fAG9+qfU38ba39WbEHY+arMtf1/fE8zaZlh48Fbuf
Gp7zeeWom107iFHuzDAlpLaEOsiAB4kxFXEB4wvNDHazB4OAtTwDtW9rTwtNVNPg
w1laxp5Xc8PIrxudPRJDU03SPcSjr4LwORPKB0xlrIreagJhy3y3+C+FYSxkwFOu
ScrY7XegIizhadsPiuJTXvPg0Zq8sAHcrGG1RDwpTpfcKB2z/8QF7RmXZAjJyGiC
zgh84CIFdoCHoaFX6EuKdZE3pfxJ2okZl/hRc+pBE0mpuvHOM+/Sm7ENHCd/ljB0
G0ck//26XCIOjqF4cstF7vRtUkEGEY8lwiUgexlml+VfBZKC7tAU/75CtqEBnLOk
Y6PE4Y0XPeWJCR8a2X6pp6gVUuY1CmuRt6L8hozHJ2OaumxqfwaPqSUSAu5a+Sem
hUvcDKESFRyv3PyfibgOCJ8/gwj9TA/yUdonswFBGkfAwvo/580zlBZ5kDtOz9WU
C0OkoNrQNCHZ4SHy0QIAdH6BH0FzBR0df0IU1J9WOquZhy38fWMeZKngSAVkxhWh
CgBLaM/8MoDQbtgEsbHulugWvm6DmBApDf4dCPhT6JBD2GwZgL5CBdNPjriY+Phv
rNJdW9TMtDq/zNcBN+lTvr5jMNS24Li6IoniPJHHdDILyZZ3paqaYu1yALHsxkcN
o3bWVh8+L9K8uulhf1aWisL7zVvmcn7tBKrno4ubrxDzJo7SNQiU1/kxOPuMB7gS
nzu298MZT3vqZ4zETQCT4HRtWDvrS8wsfOrmkDOGvb9O7wVzz8/EIXxZU/fgLseI
4QS0qAf0kZean9zSfbcvBKCnR8ElF57BONC1UNO40cFIm3vVSnv3GLRetkRZQ8cz
AJlQHuhvzdfZZf1bA7s28pLNdEvMiLkRI1jg0dcM9R2vx4LQQYm7hwMkkmRUtf/+
nvdvkCSZf7rL6bWePsc74NB9w0ARlm66V6+8rzlewcY1p2rycMiKW6m8uFqSA5VR
clvMFs9VL++07OqPQzt3Fs86y0gRSDZvSaazdGWaYi1uf5RfnjEjLHaGryA0arP8
Aqd7zoj3Dc61FhLtOMO6G+0+/XJLSCm6zHYKjbEG9nRpuREEVYAWQY9ALFw9xgap
OUTh/JJU782xEVSxTrK5oG+v4Fg+3FNfyW884DqoqAjYkoUd50jaR732/r8ozcba
+twFAUPLUll5X9tkTaHHoQvs7jAs6ZW9gqssAhYB6GnwkSTxr3/WFpcBQvEa/GFy
m6qOOPIoDjk0pK9RvEEgo6rtNRlMSA/SOPLrquraODKhwZv+ifAr1eMtW0SMVaMz
HskVI4VzLYr7f70/J2q7N+mTuow/4Dp3m2NFqyKcQtK2GHxfLHD2czTF7COpkmQB
Bgr810xJLtVsuhwl21ewVSuNVc6JXK97+A0cA038zE2wWwCJTJ8gC2ESFY6xEJ7q
dIdRe2NdMJXx1IT+IZf3djq5IgYoX6Bc62Ux0eIakq0SURQB3urcfgkLK0ftrYFM
GskxoFttJqirN+fPwko349p3/AkIAxiW+GrDNfBiu2i3BRCKQHfOLwR5QVErxFYx
YlAD7GInBsM5yLdYOZNrxY1wYWmcXA/ZHPtlC4Kh6Vhe6kWHTsVjYImFPDCcXCoJ
Rru4qleqGz0IMosOy+BMXhbWK1pF3wvoAqNnco5CTRo95I7wwrTUtUP2e4SIGc5M
C4cMZG32MmmVQTYuZGOi6MEeXW1eFeyNcIlB4nww5sTk4yGjnBJWMYD0yvbzkwkt
N5PABZWKkRkGPKKfZOoMIKUpRZAukgPudoxBGScvZX0q0wylQ1si8QElqxDbl5y6
l5A4ABscSbn/CDdL+8PZLgbhGZGu8HHy+NcVTjfP51nq544YqUgOieIu9YBPcjag
DcpBbBHvZIvHBXg80jhPfD2GH8b/X8lhZ0VojwJm1uExOnr2g+F7Zx21Jy9ClhEw
8HfiHRwkxDUqltf2pzDHeS9rzNix4GhvivLV6/tZQfXYPkr0X75nPPRCD0YUzyFg
0s6g+gul11R2anHLRWrG9aK8Zr8BSGE2N3uAnGSizW1saCExQJIt9zlxCQ7MBKsT
2L6rkHiO9FE07/vbsFdc6I7tZSuauRoeNEFAoblm5kyT1ekg1aePOfhjLCTuXdDH
nbN4WmP2w5/yo4bz7YFZiqAUIiIahhqTGbl7NRLGkTSUK07XzKml69VrC3XGt2Xn
UPCUI8Bw9GJ6rb0itPBC3CpAIt+mxQ4IT5wE4HTpBwL86yG9fFLl6CpvbYwN84cr
VxidcG1QafwoJDDds4lChzGBymE/pkOdVX2GGlV35JpdcM7TPKu0YH03qM5CAGoa
SHvQipbin2bgCt7ofelPHm8QzS/FX6VGaTEJifT63/ewVYAjEv8DBTszteDFqWaN
e0ofkLYHkLMc4UPYcGd9Q91WvUFmiBVaU0Ag3OaSTC8GtXJ6o1OacypkMezVUYKh
HmuuWBTccDxdmxAXuhDu9QZK+M9b3yuB/mcrQR2WVoLVSJZ5YBVwj3qaoB2fBNk9
24q3/8UolFeUnTiwSTXFFDaHYyiOCbbGqNa6Vs4vQX4jPtbsug/cw81nvIpOlKeG
3ZT9am6zix7gCPF1ijFJNHJ7jKipHW6S3cnh/oTLi9ni7jbXPetHC83agKVazbJb
VplskGwh3a+u0OF8KzqqP95BX/qxTrqISxHFao/y0VYAMVpfTtGw3JMtnnerkfX6
mSxBEaW2aPke2caNYb9g/JEfi0vp3v4G8/UvHnAktYcrob77VHp+forDV1UP9E5I
5rcVVe4SW7ab3ADQsz4ti44gZTQdZoN0JjP6+zSKij00ZAX1UDhSiLqg9ODTTxX5
OABqjj01qXzq4fRNKyaynDgmc5TFv0Eldcr3NaHV5UDjX6wVWLQmyzRzT+CG+F1B
+7EefMeFD5867Ig/sfkPpFYoqWILWUFVSWf5cdAAcnKfhGUCcHNwi7Ry0H6ltfUG
9NcPJ2LH+o+8PystvP5iNGC4vJQe9SFOoP2VNfBKZQYX1t2ki1iU2MA/NfVyjgGd
P9J9jitP2vgckGHfdTwF5Ozr+fbn4yZy6Y6DpcrbfikNHGG0610yV9otND8TwVvL
1KC2dP/wAaVVT4CdteEnSa2SdpDk/F29TD8KJBv8ZP3BbRIyxBy17sMdvF1D94Z/
2ChSTkNOf04l92a6roXY4TgE1Qwx8wYeiI4l6NkN9eDM2Tjb2fACCuvjs5mhIPZF
+YCKgefbMnHuON4yQ9ioeFpvpSK+Nn/97fvoWQQPefKdu7q4uXJsOXtM4IaQnEPU
qY9hCV1F9YZ45TW6YYiQhEEoWyMJHVlTmRzcUugLf1P4lGbRRrXc5vLAsvlprq3X
PUUkJ1THmX/AeUS4NQCPF0qRGsdKBtuZ6ec1ZO8Z5D3slx8tYM36Cdd+FiAPeYWh
x0DHHwN80NXdUb/EoDGsDey1amF9jSwtfW47ozlsR+vdl0FWsUS4Y+aGpUEa8776
iuHUTdX/3O2PuGQkKCgfDQL1QBI5VGhS0LGUKjvMkPFo3AQoKCKCQtDxp0puXRC0
9sjQfvxwIVLpcFthTgxxYNXvAdeEXAShcspJjM+1QJzxMS5DUDUQ7hN0tEMK8isY
IK5HIo3mDXGjflIZMOfY7r4k0xFGsSHpgZON+7Ie1LSwsTXCmFYnk4yrHNR9fqt8
4nqDIPkL8ddnknYpgdR15cLfZ0JYzXX3nGZ63pAjNhPakSAn1FhB0NDDsKjJXH9l
e5WAeSW4kBbdkFEGMDRIIxJfDu5YxUjI1ANWFPTSpu8FxWWZqIYeckceL9dKIxyo
+wuOiGSpY0dKIFfJ2tW0iV9CUutdSoyMYd43nVX/B90HyKpQIun3Zc5x58bJLp4d
F/8azL8nKSg/552czKAKVCBntBsZaQQdBdFI+FvlU3m1EgEfFq7wfQF1fQ5aN99n
BmEhE53HnXEKj1eox3/Epe6uXXqE184Pa+2/1zbP2JpyrngvZPo2f1Qn04436KfZ
2CsCp3pSsc69VtpDHeztZBNdhE97dJVod80D+LOVMmfAL+HnQXzgaRu0iihN5OVi
mBOl3H275Qv1U1Dd7EiQbcEIDoimEnWmef3Dg0Z/VHvFa63h8OAN7ftd6VThbCZ5
df7mGgM9VPg/dwVVYcekiMSdiQxXaSDCgKE1Y98W6sz5VqYVSn0shideg4KpNKHH
34XMySbHtFDauMyvUTp6adWoJ3pkZcVqO8p+LGwQIMHIwDe8IdpmaE5OCW5T44kt
7/yegiyNDtz+CTgQ4TAfeTWD4NvMZa+LZw2X+DVg6MJjeYgDYtFvyKV1UgI3dHwZ
5K6zzV62RYjmxJZYVQn7kPfO+mqatV8gaHKeBY+LiS32oA9z6LZr7Zgm2PgYV6Kl
O1Cd1IfY5rY7gbDsmG+2GiZUjBL5FD51p2/NWYlkrkhJiaQ7xHve8RmkQCFecg5o
i/eFIJtppmYjTETkV8REegzLQ0C+E8xErtC62dm7FGKmi4ijuAb4EffaDHlU9mej
vBdm9YKtIlOFFQlFmDoB7bGy/xB1XX3b7R5+SdFtmfxTHMsro7Mso+dwChE6udwH
GnZ18pH5jWXW49GrVoOJxzp7kyj2r92znoQceLEiNKgg6QE7OxqHvpnO+JsNko7k
ZrfuUuZ1/wS0cKH+xPct3cwlYhwisS34dee5ZcMuWhrCN7Uyd6JeXlVXQgbx1Qjz
ZbVaBYsc8VlRDrnF5RIZN3EdNwdpDIu+jmfc3F2KR/jTJxLasCiaiyNyMDsdDTuo
6qjeCPJzHOQCpVgpxIlwyoxion1MPOJnnsuodBb/sMq1lZVb8X9FhX9sk+MePU8g
yuSAvYUcrniI1a0rNW16fGCykNNZB302unzKKm2dqQaVQ/xpAAVpJIfwKUc0rfne
Se8KKwCyLgb9GwPpXfjRF0q3feuV5aXXe/xpe8eqUGMALBeXrfW5LCWjwlt5EvjK
f8zWgwvikG2tx8ZrOnR3je9D/gihCGjTHR6/Y3g4atuJ7fZryOfkx+PnZwLvga4I
PoGGQo5CUEyl64tuyAgUR9r3CJHbUjUInT8Iqd954ge2ijd+lNFzv7ApH8NPAAui
Dm7YBmd39vwXJpts/WMB7ljvYd26qtG9ZC1JaZkbfYS35d/+w+fncJzHHos9vbok
9Xjc/bFQ3hL3W+DeZ1Sn0oKC+YRx19yB75Vhxk3qMED6/RJwBtQd67/InwXcvFeC
H/L40ns59XB2hE83tIzTmW2TWWjA+g5Yu7fn1VFXpzKMXcsyahp6JE4ACqx+Ot/1
Ka/KvmvuW1tqpWGS3zCKw7B9HUuYbb74H4od1PcRj3hhQ1TmuzD6i8uZr7UsRh5P
AM8u4jCxZnddbIlR2CQy2UDCCg2zbd4jttdxt3KqJfjufvoLYi7YA+9ZUS49EGtX
ggDjPfsWxwE6Bq1oP9opZ2FMRk9FX4g+R5/6d0QdDOvNfqH4o8IL/VDC45PXsxjL
/ktz9cHaEWVzcOq5rq+k84ZkVH34EI5m9F/qhmX4JPWyjm6VvhejZuThZpzK4kHs
KAUVxlX3lSYhHv1/Aglajf7jjDmtwe4AH9FKUrXWNP9ZCItXVCQ0yc1M9jR/UrdS
fgr/5m2otxIUcfEslfgHt+3SraIqmuD/B1Y79ZXNhoNFp371XQQxSWfr8F+QJrea
x9ZGLfJWzV378IKLobynPnzeKyPkzvqy4S2gQYqhseOOi7faSmuf7pa0xkyxUQnT
JaXNx9x3MeQIx0gSvvuZEtaL2TWWtA5jNYvyl1MFBTpOVPyCzon+LshQNlGs6dTA
zOgLWCY3ZF+6TQnqeUiEW2nAQJeiU0TtSOBDRqS5i/uyjVdtoRFlC+Q8wRjuzTBe
o8BGqyg7rpbQ79JJP7KJENtPBOQYEvEUkAKOizXyXZxQizVOID7P4BPMx3U094Oq
apu1CfloVZNKnfcrjf2PCOKMn1Y23roL7wzdfKhEzru0noKZKVeaLpF0eUftxQ1m
okqMN7mAnwJijFidYsvAJBgBiuTcW7LKR6CT1dqMVBGoqzURSZ3r3n5EANNQJbNd
6NvMoF/QGcJX2UhZUegZ/jp/veghgUmtTG4ysVeLtB8PTm2AYQlfgxq9vC2Cm4iM
6k8pbdmNsQboqdByz2ub7EZKW1TCMPtwzl9c+ddFAiyqGXwVW6AyjO/crhPswfwz
9fdnOlAMhfRXdhnLimlQ7RKsKSI8zcwCKstualgGKzKW1nYQ9fbdG6+6xWry6IGk
wTOHPa9Itg//2/9cuZT6wyz534MNozubCvnrt2vQbjk1dIlZ55WfgrxmfsqSKsuG
qbJmzZlaCrZFW27IKaMEacWEeL3UlmtuBqJ0n68foTr8ubsHi5b1n73vjUmSG42k
7QJpFjuBqwPoYT/ZmHzjegwHCuaTuQYYJhaxdnsQrZ7S6OXLmolXnbl5W5+FG9eE
CXKE4Onu9qbur72eMOEv/vsbzsI0fgdweBgf4B1u+Tbi9RlzXdnDLgkbCxTX/vEp
ynY3U/urnQuQxapFdztihu+hmtfsPEWhKPPkG1j3Y5Tx42EPLJztwG0ubl4xznuz
Df1KCKDWhwsa9yWE4fPdAo4DeXfOygZfXHZWj5gaEWlXCswceDfoHSQunM/mDXdv
Gu5E8RH6a1rj7OG74CjZxUaI1PXU7RerW1SIkh3WE4cpkbmDCvnmdTNgudrzHzuo
HAVCKvUtn6Xrhr4QoiYv183gUMLrOx39WuEzvokkzXZBssZTjmGMUQ1T2+6UfK7R
urXgoh+NF7x0ch8HwssmpwwYHBTPGk1tC6hJx4w838K8/TKre8YQpjrHf6o3P3T8
ubPXb1jvvQTw+WhVHXNGEDFIU/TvqFmJPnd/WuYSTj9lT/4+uRvMrtIx+hY6epc5
e74VqEClSWt6STyO7koS5WsYSs0avt1/vzaSDeDNx5WY2XfDZErM5ypR7zlKzoEG
adav19QijkS05rxt/dgA6KxkXI3BTdNu3PkdWJMjKBz6X4ZLCibIwtG8eL8+KMfY
sSCOhpo50IChEDwQtawIK0iB0dn2NQAY8RIuUw/w4IuIV4Zt92bbdUrOnb27IWVh
K5WC4mr8EAc5TdBT2wuC4kbTHomMHLMgHP9vbrdDBVF6rb+6Q4TheK9t5Ml2rE6w
xXexNOf5/CGVC99XH4egeAFYvRvn8w/j0jB2+JqG67rmMfeFDDHksBSbPGKWu07L
FCWsQIpDpXm7CF9EcuxIc1VXhcY+ruBzsenZJl1garwF5j+MXTagrgkI+xYgq0gv
o2LA//IbLZuAyMCvFPsTJOuzBkK0/cvrJOVm3YksoPjaqiQRtvgh0u+X8JCVveGW
OrClPTiZUp27F6vnuWd7oF7OXXXez5DE70z7T6XH5a9L3cfDv14HwEWTke2wqPmB
FD63osCGIl5y/oHYnjQESXTXMUNCS1VVl2bkfxOz0DzjzEPxuPHZsP4LIVvkKcLT
vrz2Hqts/ea1gUG6WuRnSpk2wRAPbMoGzvQBjSfm2NGwPDBO0KPtZjpAXTDYLrkp
PQadHDRufd6Fb7gEbuzymyU1qIgtfqAC9theHVtqpiQ7l6wEgZFAzry/Pby+r0Ax
Ji0n/pHtcWTi2X2A3r2GfKPZwpwdpF12BbGxqGwdxG8hjnXvCDdNI8LN2RdPtEDK
k+fGxKVQgIFqUf0u9DfrqDhpqZV1l0vnhJ6A5bDnHCIVXyC7sM4BZ4oBHyMvAHGV
tkC75iOoPJH9hN6xAxZ95gbaOdgli78Ceee48EG6mhdozSx4h2KiJTcRJkangO+J
V6bVgQSTFQbgLiaGjUgsHIHt5B63jnWKPPUUAU4uX5bTtIdR03nsa8ujvVvqgG3R
rNyWlul/sXMgjZoFNSHneOl/GIf0OYmwqqd7MJ8WhXgZoyDCSonUebBayRcbpv7R
nenYDIgzxeBhf+rZbOhuvEgHMzj4uCtK/abqC7qhm96nT0CnQXNTwZAhny+EChcR
nSYhjkXrfJthKItaNcoZ7UAmY+U2YwY37eAwksCoFpEvSJrjW9UKGNKxmzqCalbY
0FAVYihHuhuGauJavDJ138Mnn+8qRs6QBdduU+nCCXYzaeUXCF2gEQs6ZmIFWo3R
jZXLLDtMagtXAvpue6uqAlmNpen/XPaU9lZtwap5B0vsY4NTz55mVS944hXcPDtR
kRmwWd3d1EQhQWyzRP7o/F+VsOesKXMQiPVoA0QPOspdq3uGmUhfAzMo7v1X+xyk
BLJv6bYZ6dhNpMDcxYWERyDztM5yJeoxqi21MWLfgjGZg4jE2oYaNwzbzzTvrNyC
HJiw8EL4zYebvoVXGJogHC57dGr8n1jFLZ1ySVm1eAbTcIPwT1fuyOMZoiSGwuYr
/Ymz4UKGQRTYLzdRp/ozMkV5QSPGOve6ScvbiH2z8T3ECng1RcCEDePeNzD7egeK
QznVKSBE67v/bLSmzQrai57RKHUmmp0da7j58jTg4TwJxoLYuGQdLzCNRqE7NBHl
AxNCrj0Os2c3LOHml/6UwGJO1lxHW5jGcBbosZcWgx9e14t/jmuaLOJCWypd4onF
vYrwbUcvqjuEX2wRQvYI4R5POHvSpfir03QPybQ+3+Z1NF62AV76OeNhc6/Ax6AF
7L1ZdRjjpQ8EJbFiqT39HFT4c3p72KOMpK6tYO3j2xa2pqcy5ggD7TilPTq/9+x+
OBYW0MIvQpUQd96K5zQi/87u6X5chmqHckzERiXZRo9R3cKWT8AOM2uSaVVsvio6
vV8yordECfdrvtwd1eZ9IowRVu3sd05zRjatIp95WOIWaa9s9dzt9GI0TsEC+klh
c3OWuNmqlsnVqCIUnmUe4jwRBLbAXbdpt3kzYYAT+a2QJNY9+BDeH3drZcT8vBtS
yULaucOGnPzFW9cLwAvzn0IsNw9iZMv5JtWfU4PosZo2Izrh25OmiHG6G3vs4y54
s4x2B81UgGvfT46cFXeYTdxDfgvTkfXaUAjw9XrPT316VebBbgLjj7NW6n9fTpqi
bGZfNUhvHMgthbHOfkzYEyDbTkmcDz/41D9WcTYg6Ja4GNi3SezWcVGTjlivY9nx
dgV0ztsfAJ+z7U3YHwbnLfxk09Md+4FtvvHyeNEIsZotfbq0JmRb0q/SUOZ9ol3M
j1c6S30bohwtBLUCYFAPIulIgAzxDMvFvnxyze8jMwKINwjGWE1YGExezrCGJUJd
XjixhuVRUlwina6FTi8JJ+0T1MRAlPmkYK38p8568nOlDJt28cEzd1OQBM7MFzCx
v10nkdanuF8aQsxZTQL6KxRvBtc8osvgG7cdp4Ix5aDExtiHTVZ28VAlV1kc0bYB
H2BbyGKyqwVxLkhgsxcyj1Su+l+x14Hrwrjx7Y2n0klocqSne3Vtzr/D9mi4jzbA
Sl5jL8FxrxTe5cHwaXXg150FBDVMmekdgmJJ4jIKu4QO1H0d/pbzqG6bQN+OXJxU
++emWR1NITVOcZrc0rWlVfVgY1+A3l2RXqbOP4Oe4hFtZV2/QHgd9ZH16YW6saSe
psXiTkky1Vvn3RHP7TebPu+nvPT6ZBET/56y81JaFACPH8uMg7rgng95DO0Amftt
H4OvdJWCKGu87jyY7eGhP2dbP58/ZpukVYJ0SZxfKcVw9RxboeNJsCBRMqe8z+D5
CEqcH8Vv9De2lQAUMOjM1bwkX4lZgpxWzEJuJjZfkuVgH95YMseU34QfUQfLHvJC
6kY4ESQ1fNBTUeeWGQ3oOQLTnQmdnV3KaUhBZ6FQIi2tp94SY6/LgI+jsaeruvTe
p5LjuJk6I0wUCmgOnDaz1XodLoKrYrKRmCBBMJMEfAIQkJKrtN7wk8VeJ3f8nRvs
4cI295leaRNHgqufamGBpLRdJdKq2G5OFSrASjoPQgkuWNAk/NvVzmNpNWn7gF2O
D13KvPv7oyNZ/r3bgokUg8Db2vfyDv42ZloJkszw4IA5jOtOrfZvAueEHPU3Pg2K
xfDYAVVmdaPoYh+5lf2/OMMWLwc7BLxUi4iiZ2sGLoPuUC7koiPsZ1vOT6lUAYsl
RZNXwspIoVYpxu3l6jPa4CW/s2/3vgmRflg4AquhkIXAw7oL8sEwLay+fFzZYlyc
QRJZHg+gHiz2KdfoaT4MvL6f63AOm9BkQH42YS1O9HrIxPFCnAwNTjwpmAnm70Hu
d+qKQ+k2bze/A7ghjfJbiEO45ljzIqufp00Vi93+9uEMB3gEcd//urkjcVLZDBIA
cwAju54MVTo3tPe584tho983udP7A8F7+ph3dPG84TyJohS0GE0TJ4l9+5083rbu
LqcgksObn88fGKYctgsg/KUOIMnrkHmEnQ7MYm1RZMDomb989D9rMUE8FnGrMfld
XWk2qyYV3yYSAFGWxOQ6FrRK6u6dD4sn5o/X3tNwS+GVDdPl5IviQYbURiKoK2t4
C/ZfJ8XgmjLttIvECb6KpU7UbUlDyq8N19oyW7CgvKekQuLdYQcyKk+bJVjbQC7U
1Ts4ppDRnqfbHA8wxzBtRNDGRgtYgAPleusr7Bgn73bDwN+Zyu838bZPBBYtbHYr
K+QT/c26fVBe3ILGXdvrZhJU0G1AZoSQ5QYYGMRDWLWjX/QvLtnji4pBdVdLWE1W
IQlC4nrXCOswue3WAVCeybmahDSYR06FUE7uzyhFhFMLoOUYuuD8wD5B6oVYH3tK
5X+JeugIpBrpnE9iX/ZrfQ4N/iIP1dihPrAsLNkDado6OFJCHWOgJ6Rn2l5Ar4At
uJ6aKa/LQDlkTLxiUz/IDB7/hFgOKEeme4vwsTBkeiFPc0jeMJyxgElP3Uya3ZOt
hA4BQo2KUQcq6GOuzbjdha8BZkuvi/ebdssFPBv1pzf3do14FVwuXi40EFYAZukc
Pz5lwcM13qGcZv8ZHdrsIFLB9rCy/tycfQ97mnKEPF/IPVQTsdtav4yCOP460V5H
Urhzk9KCPAa8nUdrjml1ViU1B+1+sSAYnha3NSLaKx2XEAjRkW7L7PP0DXejG1EJ
c+ZuXFSpd/k2jqPjFrs0x3vHx34XaSkwUCXlQ8X+xIFOeasY5Sp5NqZOmY9R4RVI
caDJjSQ09GNqR0cG0HMbFebACrNT2T8m4YtBWDVZw1+TnGRtIRHsQt5PofRRC3+I
bp7oONBDxfEPF/DbCZd9uFpK0ypKysUwCtEWuWEgQWiJURUl8g8mOCqIfn+OELV7
CNcYp9hIYqefhB6dq5uVbzwRheKEKvkq8knqxujxRfqu3DFvwq9mVCsInwACDDj3
UZV00UibT5VlTi/Ew6nyNSxAN3ZUGnxDETo2v8EfivOrsEeujnvVgckio6uCicUu
n3BhjVn+zth4y5HNDVZgVcBagufVlwuoa754SlmHkxMScOopEgOkosnxGswi4mp8
0sTP7EG/VckkdT98AdGP7wlY+mW3pGTJSow52NeGIzTWA4NdIA069c/R0PgYsqZF
V6v5xVAtPPjjcqF/lYFL/FpnSvS52sFlJBoJki5kgK8dW/aUNp6Z7Uj/xZrIJVfW
Rr4VB4B0KAGEt9IWmZbfEr30iLcCYIICgDwPO2EppK75i0PURz2bQE4Aj4VIvq0P
TSqcRgizEkMPfl7LUbK1m5bn4/agGkfIfMdImqP58lBt70rUXTAWj4qVKvrrYvjz
scUoNIVj9/UxakGjSGY5gjmrVDYheTH0vjiXp8FFwnmwtIeJJLmagnE3WbZrAjXP
Vm6uM0mHjYMamxS5mNyRMbz3uiSq6oHwcBaGcPb11A2TG+bZC1Zrw5diD8evg84o
rplfm1t/UIRpmWK3EIOs5gM/iYv46fPGIkPFjK4mOZlBLc+z3a+DT5o3bWuFhc/x
TCRCuWFI/opZrNAY20iV+pf369WYrS2HOF/m37Ho6NhOSQXc+VX4FwAhBftkPVpC
84cscqTA+deJejk+LUS1xujLKUzhiMhCD8pLqouXERsPV77TgD9dA2+y9uaysl3a
Pqnx69UsHKHKSYTSR90boeUkqc13iPcpNkt7dWlyPIxw5J9AO399yznmGfNz+ub2
IewfIBXM/wGH/Zw677AdUTa2bfW7osgpqijq3oBTxHjF2O69DgOXC2DsUNyTRmaO
z69d9Xvp8Q4osDsh1LjVfvUXIRcrFDRp2qPLEUCTMjGR/+gKH638cD9i6cYtj9zW
RFRYPwZQMfT+iGiuRc5fgE3UDq6oBmnXSj0FeFrmERo1OCN7EyboKclmH0V1CNBZ
JPdFm6HYGLw0KXSj7EHcUi8QxPi2Kka7xbS278NXlSkOHc37Ode4ehTCyuq6fbSi
FCaIM0Ja6glO5AUEgB6ZdMMkA109uvK2LqBH1/gpWDCzieCZvU1hVhoeBjOwuRgN
gCbIdvzjKoJxeGWO0L6OnTkcHsQoF3Qpr0tJSUbqs4FxhTx7zGtE3vDQcXcmVgmi
AdTI74gXPr19yUUcdrfld8z/tft+HSxVhEudfPio08unkRk8mJqDrHxcyLDOZ3iu
QWaX0MKgnl8oR9eld7UZ6q92Ul7zU/jHittiEP01dGzUPKnm5yteLzjBDQegL9W1
ND4D580Fy/uWP1CA9x+/zSS/8GX7EstNX5mY9vsdc1oAHDzmgt9CmxpH/Y9kxuxS
LsBwJxNvohvtp3VImTMBU4MuzWYyw/yGNmkvS3ol6B4IfigFzQtoynmuTW3oPB8m
YkOCTetrHmfkkWMHlDyMlfE0u6ITfvfk7pt5yKd/OCP22pWwb3NPG8jPUvlbnL1p
BwwuYMv7GC3a8cf2RK9J2Ch+7v3Jb3rqc8vWQoDVfVD/q6sdBak9I8wF08jlDY/q
5MuIy3ysqkg2GRq4tL8zyVkxNmd4yspcQpRXYmGADoEn97GqNK/lZO5pB+v6UZdN
79nSg1hXG3IItLzhTbhE7qQlIVxLDEhIQRMLyO5q+OaYvEmc592BRpuBkfjcHz8+
PGuppYsZze+pvmAg/xR55Uta7PKn2Rm5MKBxVKX0L8KuFpFcAIWIpIrQZnuBUhP/
X/B8nc7hZOcPj/pdL8uvBcIYfQxPoClhmdGFXErrbTJMTbSyy44TD0yuzJUkWfR3
dxaKKaDvysXcok7OChL2CCi0BlfRJviB1NtLHlyyyEX4kDPrYRksGKrooDg2Ecfl
MXI040cHRcfn7iY+tw2/Vb98C2/C8jvOqzirV/mmsSMht7cSC9tr6LxAXzOgQZCI
RfYjJMmFN2RhDSSpaYQoImY9nz6iiltTqPg2/xONsBScnrAePe5zB4cWpsA1L0ZK
07VQavioJomda+P0Df29JUX8TDtFg9AsAYQVncvXwGwPaOFlR/1seW9vK9jM0Luk
eocDZXE1WlZkxDk6R9h8UpOlvLvq/YEloDixiuvYf0ltkyVthXfB1KuLL47tu1CV
KJJcpad3Edo697pbnNQKozNcN8o8RgyTgMs9Mk/rQlb1hlN2y+o/5ZG5QH/BG5u5
/m5dV+1SoAkXn+1GldldHpGfJshw2KokvI3WSbi8KvPuQ50xWNLCRuDvi/eJRqD6
ZAtX8VZYsewwgLoN8x7W0enkn4ahH9lU6Od54t+qv41bZANKk10QPfXkpWG1JJz4
xPcbCpzOEIdEYm1X4/45x//V4hQGclsr7INZ+EacTMaLwSEgS/uka0TxL67uJfi6
zx3PsQRjXChnI7DsnEdZwPskIdTa8vaglNAtXzyP2BC0Umw+25qtfK1hEFEgvXbW
qRZNi80pQo3ueH+cV2eL6Pqa1G35izJe7zqIilBFcRTsyvz1EpopbQNtquy33ZQj
F7hrVg+ubxmESnRUWNMtDanMslEEuaLvoVcLVF5OfQdY6PZWTFc8ywY8IIhPDuii
sM5V1AiQqAU5gIetDy2vcSqqkrR+2u4O4gHr8OWZ5Ct7SjjhQkssvcHDnyL/X4j5
sXXOKR6XnArQQaN2QX2dTt8uaPljeGVr6eBBTRc4CqahyMNppKEqpyGUG5FRXQYS
SXmUUIStK1HZbPTebJPgf1V58n13GhbMvAiozKxjZZNg0QXdkf6VNoC0QVPahYzt
z1OjcF1duF1IWXxLPPQS0j1SuTrzzKWjEQhBMaxU5SmuCSz4BCpLakKNeTAMkSHp
cyoeig39wn2nQbYs+zBkCl79m/O/E8BO2BSU3tqzoUIwMxcb5N8igBVR5u9+zolF
yqyIlMAqnmrj3PMmrFslgymW+XasFOF4KUeLQcfsdSFxUbF5T/rL9aj/0vhnmK0A
sto0w6WuUbo5x+0UZTNZFb1BmxJtIYUcIXFnEPjslUHD2egkVy3kNqJ4mwNlW+p8
pBgZZTj6URSWjXPNSJkMnk90prT+n/N5dBw+tyPCjImRyZENfsfy9/ze6wfPYxfa
c/cFRtktAIYDHaqi3jkW7xPeUu3pvYcgxFjY07GO0axof6W9t9tvQoKqBaDaCsPQ
HpAQCd0X1+Kso/Rnx4Wv5EoNiT/g4ynSgPPHzCfxtqNvwNOZ92DTU/VgOi2/GF3N
pqdP3h5OE2qenLeVlmQYij8lwZ+Jn4Ws847aYNeIrVU8F4SwrcxRs9santWZ4ZPQ
4dxElJqyYJN5Z36sSQu6hO7gWA10fz2v1d+BXMKXSb6TiW1uLMIc7v3gmtNhhJib
G86SiWqFgCbtPHHKKXLbfUJ0EIwtGPpzgkBDUEeDCN0eBhKalcXAU2lSsCuGuG4L
elmGQd2HduHe1qECYpFstJVUIF1HN14iX/G+M51x767ciACF22wwy/pskUGaeIen
E3xWYxdPvTNWK83o0xMeSUZpVjDuC3PU3GK/ldZUmQBrhnoWjWSJe7CWNCVqdTXa
Lxr2TCBSl+kARd4AyuR0TFeKGWFXCKU4Jwv8Vi8FGgbP90lVPZgUudSnV0VJO9RA
KkVbBD0v75se3i/OSmkyMn20rsRmEwDFs13g1EmOjtYafj8UNyqc99ROW51yuUdz
T4mv3ZnoKK8lQYRd6vBH6gFEgGNxxehBUT822bP22xtOrSscyLEo4kz+5LN1lOAO
Ta99LMyQlTyyPFGcZYUnHUtHTBT+MIEONldkV3AAHtTNEXRt8Owc1HlR+xV8RYYb
eXAWT3mmOy7l95KnVaTqNe/CnEPH/ESqIrnsU5CVPJWLKWm0sbSaZfE8N7SiK1eB
C2P+zMo5K9oAz+yEzmhKbTBX5lZELAL8owfW3IdwvjHTZ8AUM/6/HNVGTi4nZ/sq
tyqyCaXZ/U/j0hvTLC07dVkrEHFWvZWnZdR8rOJGGBv/7nAJn+Ww2KryLKiTV14l
UeQKeL3kbM1LCHFs5Qd/YAqV2QWZOzyOqPnkHIfOWtxu/0vF8iKOLSlUGxDBfsiF
H06jiJP0EAWVIAUyDV+ZT4cFCX5+FBv71SaZSaWxD9a+Z+ab2N9it3vasKe22O57
Ads9gElLQv0YMf23SW0aiSBarq/SGF0Ylp9uY9horMEs0T6GgbFgv0yqgoJM5yBU
0ZU7HYjQ7npcCbAbIIVzK13aCYYS7wURGz6cG49buRhiemHpNiuVA0PEAhk1qqRG
c9IlkcpyI/rSKvV9gMPV10jbCHcjUcgaKPYZ1L5gTvbtGDwf/aEYCjCatcfYn7E4
blvqaScUbNQjwFfzxSLMJaX+dTXdaIas7RaVSIwVaX2XYDjtTotdFcKa+cVyxbQW
mW0dBpMbBluDAsXt6YP04VwMPhijkD528m1GnYv5eRTMq27C8H9P3W7e1ebAWNfC
ZJUILL5Pyd/7jZHBB2sAvtrMdINFInXoFhXhnRV+tNC3P8IOMrbD9BwNXDk8dy+3
0lCICzOYPxT0p9d0DBv8jXvu9WeDcuGRnOX2IXiCD67d2eAPsGfk/FheysozfPt+
Mj3v5ZD1fVqfP4DUHW0quwig71zYVXIAQ5aIr/T1qCCMxOtJpsl/a9lJp76h/zkc
ru7TIng3hU1GilijjI99NxBtJAeJgzwX3Lxz8fOZWRHX5WRsdHwVwHc7X5QQULaT
B9lK6W41JOoPKlbSJnNwa9d+YNzFFgye4UXBCBLO4dNrwqgW8qIrVj67aHfwhKSJ
NTZOyEJSLhFECmyMGBq2TZbTDtQt0YwMRAPeYkmqNv7iCdjkH/T40Re4Uvs14mxD
51Ypj7Er+fOp6OAg3c/hVDbqEsDbzElwNddcp+e38Sc51/qaRxu8p+euw9LZXN+L
l8uZjVOBhn2yT8f2gObol3ApRua3+fNYtL2FRABno4lPem+3qtQvAy5EzhU8lnN1
Qj7b3xuaX+VFKTt3FVLvIAvojSpOPdLhnJrnSld55CDmnnYhnEh4PqeodUCpZ9/l
DQZe+eTtUsRVCJ86uqgUr7ffHWOG7KJ79n0zxi5bWYMDvHzCpM7BdAsvxQi+FO9e
kkp1ONsaBVMx1fDnQqa6aNQatZhfOObzV2ELJ6YHz1PjWaptAD1VbF5WgI2Iwj1F
TKUeazWCPMkpO0zGC0kvJXzaX+K15N2AXuFq53G+c+aT2xnB51tu7LC4g+53EJYe
adJ7lcZ1MrpQAuVZW+o+7lI/iNax0DkowE7tTgbQroah3DaDNh9WkllUI/6ctHx0
R+DkmmpNqnxsX+18h1WLehdFaoPjaguO68a2vTbJOWUlz49N0GdAYyfMdPlfl2gU
UhuBJ2O63R84FJZ42O/yaMuuFyHa/CMVM4pXipcq9XmyurUQjXTPvBOZQEv0CWbW
lCjEij141nPD92WY/u8LmlheSp5mrQlc7HI0O6lgyjaxpTw6gfNXNuC/QH4bWmiP
u3MZunxCoUtxQ/4lcRKwo6uXuTdXkB9ANT7GCxSHAfUZQd7Ytdw3BraFneyEbjZa
Bu9X9Vlqsyykh2f9siBkcPBxMd7DAs8xzSFbtBtCBcEiKjGFn7GXA/Tf+QgMTDRV
pvN3DWOkvz3R6d4LY8AMb5FbJCNoCo5rjRKqLS6/vCJSNBxvBZSlDZexzZcqL9nm
ODiCOsk0g6DKhX6+sz7WliFeoWdgbwDyO3/Igs6k34pB+BwQjyL78pP9XrP0QW32
+A2spSr3jz16Mqw6Hm7glrb3fXP+awoRll92+8uKEP5VGt4qEUzWwEq49L4HgZp0
uu68GdgQKG8A8ItfWSczPT3RcE6r8ZvZ5+DsNX9XLrKHXdkHaCJRnHdP5euCWzck
ZMI+7OUtMRDXFrM2oT4zWqn96AKB8tiBKB2JlYHhSSk12aeAVYWUuDVmd1FuknRu
gPO1/L1M/BP99fVdaBB5bFbi636h29ozEnnaEOdL3zws1VRiIGmDr7qEjfoA0nNl
h1D8kGu9Ni6Ka/zaDpBLwpBjmmAl6MblIZ73j4I0T5CwhQYh3kUp9W9uj5C9rGhT
MFOj5gMakRo6o7d69Qo21aQv+GA2LsJ3aMnq23VAGdPYQnlwg56cCNnmc7CwOhAc
WPS6/9GsGCIQdYeutGF8YJuphDvwaPCo+TPM3Ed0xE2l/pPz0Llb5yITdXaDn/OF
ptPOKwICxHz+HPossycU9EP03IZ4+uhkUKWwdHDkOOcxcu5JUbO1XBr744kGDh85
hgbCbTb79F3ZW7Wgtr2Lhazpskb2Y7++EnoifmMmsWAQOsDVfwmQQPvfgVJ4wAI7
VDivt1WXFazVwQGy5emYGH2YWHxznwdUYEEShurDUb1Bk7ID2G8635tVw3cnQJhM
2pAjOCl9jIwaQhTAytLgm02fS0fla3OEZ8KVwSEybb+APtMHG7NXRIF2l3x/LCT0
bTCqyFeT6NiZ76mC5GMJay3B2GUXVLP24H1rZBiM8SFcrtMm9h4Lcwnk5mzbUig4
4dKuNp36bM26XAAuzKHhkUCkdBNAu45RKcoZarkY1mIPLCLLVe568FdIbGHHSQ5f
d3CI789FtsHrUUTfCXBnM6ramDtIP6LYyltX14nxE+d0Wyts8LZnXvjrFowgEsTJ
J2JjLbR2BpF7uPD1gWsF1dUFRuFh9/vsriMl8JnExG7d+fAMwFUto3dokgwadbl8
i8kOpS3RZJOMyBndR++5DPERqJaTygHxZdgcGG/LLDcWMFVWjTRV29CcMmxnQqKh
esh0wpaYHdq4mr5H9KwfwVbg4xFOpPa+fM3ExDTrxwDRIowRy3amCwWRAh5UC00G
UzSWJm7JMZEeiJ3C+ZX5n/mpzcjVhGvdIiqJe1gTPKPWmEEItbw+IxWWc28pSbx0
pT2hMK9nFzcvEMium1Phoriou6sKyuaiZQWrtZrEtK+VveDQg8cXbufR4UFX2uW6
NFkz33mH+YYf21kZ85SX4iMp7sLLTnCeioZotYMJSgtl9v3QFdSAJFVw2rUw9RvB
3B0NCsEnvoN/ZjzVZYB5oY1tebSnMHv59NGEHfHSC2g7a3YTDzjzjVW9hpMTHOFM
Lh4Ois5jX4F4CdShTImcfIpT8Img5dUzwqSV21CMXfa4gkmcJIxB0GTE+rNtCDTI
S40i176pCEpne07Uvl7nJmIXsxf3fSNXrE7zuPzisnzJSWKQKA1NoWtKAFh6UKIp
CnunaKttbTsmkq19LX3tiqlYnjVlR7slEYvuVkr5TjOtY7ZG9oFXaiOXQT0R8F49
eRQwm1GlpTEb6p9lvconzqVHlDDrG/gNvIuCU474vXVYAH2QlI2ozm3EEbBFTX0u
vDuvqfK4SmewrpJcA2tiGLzjEyqT2GXIjvrKbIuAZAkJL7GA4wD9zK6MZi06qtCw
bhQurZJVJmRzNiGgFifQJdhWK/m8XHgj0rJG+qo5quT7oUsAxUgKtDKPZLRRSxyJ
oplbA0E0nJWOqGWdRLzfNymxTur3y42BtrbYLjn0V85dD3/+hZwAjWjLC7NDgKL1
/jrGW74pvtm+52CgoxcvES8CfbWDrQugNt8dTVrk9+4PNO0xuvgdsXWl3gyow7dm
39bY+1PbdIGFTLvoFK62fWREhErQgpqiku39xZzhfxlYrMHsqwvKZBQ13BMuTuRl
wkzLzlfVFRM5yCzWqDfvN7isn/WaCpEtIKQm1yh5DuHdWgT9GEHzqn/ZuioR/Nhy
haNGmFE0ofrofM/mqSgkfWhuhNYGzhJ4cigJDW28yRqj5jDkQQDV41tqmtvkNy7N
66xsWjfRi9boRFZ5lDbQ74oz2fl7/edbj5lW23PXkvasu/fbZnxGB87KxLTqjca1
+i0FLERzw1jRrE/JbZwMdBoCJs5KJ/OBFsZXeG8SDzVWHiPnOrqyLOsxMacSDrR0
Yc23cralnK1h1fDVWg74/E17rRj3+5xnI82288YqwDQW3AYw5+LCZOyQvE/jm0Fp
z1790NbBMXkZy5/8IE5xYc2YuJHCmLqRIlQ0/7Njujary8N24BHgzNcuoB9diaM7
Rj5xlbo7nyFln+ciViouJDoYWc9tE2R9qI+jC3jgejToKbmBqHtBaPqnGALrqi9V
dpnhwYM+owkFKkuf65pYES7nlTs0D4nIL3Y9+FMuCIAcJwqwKaIZwvfFadIOWV/3
Er9IhOR8WhUOJNclz8Su6WOMudTbzXjqQIY+Vl1P6CFPoq5HS1gHqp73/b/qrGbo
ct2H6b7clkOGjKHwgEIs2ZXg/oFEGEmWXwSFOrRXoe+Z6gO77TkXaqili+mgdosQ
UGrM98UB+bGfxlwfwyKcncw8EqjbehYQPecFWRJe0OBU3kg5OwOnCqeY4bcCpcoh
NZBanv5quF9UiUkGsHJk0eLuU34x/3C/cp1p5KWudFVSm27M/ymJX2ZCYwldBBtW
kk5OqrkS0JKxYj1QRFJV2qNHyAPrBc7r0BMcE1B2ykE7xnwud+R1rU9uDMh/EAbm
bG+X266WSJf2pTNw5dq82sheHVb+0tKg+KWPwlDd5cV25vdopXmemMTVRzyMrSLw
rpxm1kSCu29LPoFg6MM8vj6GkhRGNo9k3lTFSmoGcxP5s492DOGHiPE2io4jYCDn
SGL8ckSxod8ZeHbkRJY6nyC7tTKox0/MoOdANuycp8Q18Vcz9vMZWBvzQGbwv2kC
+btdikJCxUrwX3I7+CZlPIB+zLulLmzK9qgfoGQpstyQyeb5MFZ0/MkYBWfJQz7P
paNvQKvy8kJstjAreSmLxATAgaBeb6+F9C1/72r9pUSpXqj1eciJxo6LEdNyuWdg
OcP+rBqF7rPLA3Fvro99pLAGo5PvDnzxWOgAFTJIkxhzZXKkTExaFMUrD//0kw8L
n3m0S3jQ83m/O+tVnVPXQ6lY39wiEmO/Dylki4JhwPXUDJaTsFTntvsvWj4QLPlT
uTRWVCcBAt2jKaznxmb2SDFVX6QV+C44RKjEIVUHIzp7EATMg4kxdnLgdbbo5j50
9u5lD0leKTicsmE2b0GuT5++7zJguQITfEjd1r0akIREVzn0st0070wJ9SGSeXSf
3O1YxHkfhFwbBWd6CkYv9fvgF9FrA1yuWNgvSRQCipgvyxnHTWkqVERqN6fCrUOo
zvCYRcxm0QzjjXWCoy/x39w9N/ss1iM1XgjtdrBCgZ+lo4nIyZFKn9TW9THe513K
yi+9hbjhYNsNctvhJxOWI1lk369q1t3/b7edMruNgCqriEAhyuFufRWXxSYpFLLL
avn1XYabOil9n9Te8xkeDAaKx6axVDGQ2R16oKevBb4eQGI2RHJPNhSuB7JM6qGN
E47FRit3gre607LHEihdsVekIUOxytcF1TReJCHImI84zAKnOuqRQVjVXLyOGBFu
ftkF5HfnthJb++J+mESpB/faTWwe9LTw0NSNNaR9W+poXsGcHeMo2l2LEG0VdH2I
sG4XtNGrlsph2az1qavKQGHfYas3upuZw6g+EEShSI2l9xMAlzSH3N//iwTrGYcC
oGluviyhk2FpkhA0TTrJbsH70nyaO/K8m2G8y6b7nnbv16V+xgaUJRQ54vbspHx5
yH4zLKIwN8oxKELZUb1vssa4/jZiz82HTQnTTilSJaLgvvv9BuI/60lOZ4lghtz0
bH0a20H2z1E9pBVwHQCn2X63ignhcnF/+T7ov/Lzbqqpz4DGysX5qHSUOkayeYf9
is1h7dyAm59U5KfY27/3ouqqHevXyFR1nuJs/m3+LlRQEXG/yQOwpv79VcJGzjMA
Wg9hTAcEYBRNS2Y3R5L/4VWOWBAgHcKHeMf1/ukKgwZ/fRTZXKWvVxSYop2QuiLd
QJv0TbxHcToSchp1SQedERUiPbzMfGAHPI1utB/+Nax/0tCVWiLJdsnyLwjuhY4R
Ia+8a4//ef1tUZ1ct2Tv2jn0uat3jLQFVnOAMJtVS4oAAXbnAgdQlQWSJujLG0aj
2MririuvCa6fvsTUFK0tCL3/H3dV/931D40xFY+W+ZnC9UVs5xznnU4emqs7x98V
kIFIfwKSprouaWdBEds1TkeLDupVGOc6sFsG9aUB7RGQMbueo8EGV50cgp4JvudS
Ktwhg9tZVE1hreQ2wbHWozSlww3CRuf8yflnODQKGDU8GqWFjekRr1UPnp/zpk3w
lUDKO3NT/ya2vwUZoovjIadL9MUFHzIHTc8JcGkqtLfzOWA0HLJIsyA3fBNeUl4a
guxxFRf2IScJwiOeDX9y7/m9LjmUTTY7zUB3vm9dAR9Evz2EY4z6M6cn50KBuQgh
wF6kRo1d16LOhdFFtl8EHnuDvYpKboehFZO1Blus69LKYslf8sQ/qfM+ez6U4ZLQ
mbLJsP7NqxjgmoVC0qOEdXfWe29yUIZwBRrNysrXJmM/qgH731eFi6xzesSIFG/l
ybe3nISNicfiSiRj+n8tg0fkBcqIpO7Thl8Ba/dLLkalQ1UE6VAPHPfBFlIUAKTp
ZYtqKJW4Bbf3VQUtuaSTIzrTVsehglk94OMqmdb2AtFS17PLhEUpmoCN+t8i47QF
6BZ8vaZpNLzB/OjCvGZVG2GLmyYOXhDCQxKthluvVqOfr5kFYF/QuGd3u3giBrBO
yJEgpKO0qaXdl8mKDQOXQNG7nK3XRwqEioiNtQCW0INiHONCEryEBNI30WpjKp8y
rF28KNy6oyz2ootTdSJ8sVRPPjHR2dhD3D4hv3+2LI/rJzp20P9RWyCcjsFtFjPP
PshZ/jxTwTeqUvqSsTfmtwcegtvY3qIDsYdpnQn4C/7bd6qNW7vDdYfn43i73lID
X9Hf1wqlqH+Zis0MzP7wr/Y+9HnzFsSh3edoZiBXfAswuvUG6pap6CALjVy+Zsb1
iz/go0na77J8W713CpBVgEe5BTqUoTcW5HQyrOsg/KCiIzF/dOCrHdkk1rrTNlxD
25yUubc8rO4+b6ECowaqw5FxZXl+lB/au80J3naGMiXB0gPm4+71ArRnBvQR6W6B
Y75DcgoGh+jHoP9t6lGmPHK9G0nXDz+5xa2jsrHdwYWqKmS99sRArMLrazqtLEwu
qk4FjcAn+1VsQRXk41jcnoHcX7uH8VWC9BhJKTtGjYZBR2etl2xwWwzVHBFLkO69
Jr2NVA+kGomEVuAb+tig2mCUdl+QDrJoV22Mr6Uyipk3FZq681HmCifH1G3FCjDA
IQZHOpFoLEFLLmnYJQZJFwzd6MQx2AgCNlgmY0V3eeJhcw1H3wIhKVZRA8lbmxBk
nQqpJMKHnocgDLiwzgL/LQKJYnJdqw9VUyjRfsARCHZLpryLRmltjZeCRMyq7LPa
WGAiLq7u56U/iVmC4Xb9fbXUQc3KA7d0Ol9u+BZk4xjkMOfMji0Zf9wczmuk0dVn
khXgMt6B9hCmUc4lud+38EZ56vQDaMKNHVyjp36BK2s1pelXKMGLMq3hs78aaO7N
9uIRfC0bOOhcuShDz3G+H1jRnruvZFniQ71ux2fGKlMULsYyyMd5e5w8y63D72Sa
w2hZAMTwdG0sZX76IjyRESgx0aOIxNkSMJOP4afZ3/avomvdaBFj9q1dLqx21xHH
9AKfFODMyWvyoVRsNHFvGIX3jyQz4ClV1QpPbugJjN0TU2JVCuIK0oiJEzX0vQ9q
mMMX5XgTs7bvVsmKntpr5+MTJ57J8U4EsO4F3wQazkPiZSHtVM/aNVilJ2kY1d5H
6dV9XEHKl+XF5ZVfs8xXue3rqoc/OhJNYFzFg5NWo65eiVuJPELqzMjHqZIfeVym
c7aan4VShAjiQtvxCJ7Ekvx7C7T/XsCoyEcOvMNroE8DMQAXML0iT9Zqwch4aC9a
JRxbOcxnmxRoDYHxHyvAV7t97xgO/PusXn0ObqQGvADQT8kaUi9giiZt503zZ5Um
f4R+mfX87vk+ShTlVEszEMqMChtTI6EaAaeo7XQD5qMd/PIsySSX+nqLIeNsmN6X
CJhY31exsZeYBwN5/O64VEcrtzzm27maJaQWiupR9oa0jU4k3J56Hb+9gfcTkdJz
A7yWjLXxH4X+vGc4XJVBIhUf6LOErmOik/fQ6+ZaC9zJ1xmFFSsU4uNbml8Fc9a5
ebhIwMOhEj94D8XEbHpTgWUByPNRBIqE4lR/99glMcsZ2K77jA7TH1eKXJrSjsdG
RT5VQ+hVxQ9hc9YThU7mGMwNoi7OxAjrdgeDr50C5ztuqRBDTwzT54GW7gufXFaR
KTR7J6b9xsxJEmVOH9DoSfp19iyrxCIANY3bPvInr0bruTd8lwzR0+HccMKVgY1C
pWQZEf3vzfkDMqoAEzKesnZE4sRdyqK+m7xwJ5Tox5ibXnyipqeAHPUd5gc8Kp7j
7AQvTuxD0MWn2V7e8AmT4+qg77hRySbV7I1d0BB3xTjKe75J6DrV/lXv2Gig1lNh
Ybh3zvGuW3LelWG2RSHczSyGckpPmkjsrrQ97Eatnrz3LJd8I5x+Tds0Db5Qu52O
axjoJx/z/rU1JtZew/QSOW6Hrg4/O//c/OklNiSyfOBkd5wjP2Aq/48m4M0b2uzE
GWXtARQM3vFq6sSw8Di1TAPO48xyalGpek3fj3nbj27oEmMFwf4Njxt7pNwnKibH
PAJUAiqJziJc9DMXL1qn67DddR3dpmAt4IY46iK2SXnJdrIEUpeu4SWCGlbsf4qM
EiMii8f62D+87Osi7AGJAF0Ck1mal84acyZrcEImVabqt2PMAbmBqr/rdUbp3YpS
RP8+OlrNXrcngEl+3Hg9TMm7aObo9s2ZfF5IVPkw+Ag5OyPb3XLg/FEg2xlZgz1x
Vs/oXdKqX994AS/EUnQ6Iqw3UEt0u9ak2kALE7AWmwpFPtEhfAmw2CRbbd5OqiaH
oBw4iZvlwgeQFq3PRtO9uW3JYNWe01OlZUVc0/mCcU88wmeratrNM83btDatjD3S
+JJm+Q3SoEz3j8BPx8H7KbB8et6/n1beAeCC8dbo+LWpugO9y9+d2wJSjdg5azhe
rFFQRFPHbTW2GqHpwieKvSmMZ0EUceWTcyK9VIgYKwRRk/8GUgAiyNCYkfbe3nlI
V35Y6qROUMpjAiESgZqzhEMbSjatsKfLUQscXDAVV5VsdbekZw7b238rRDGi2+vb
WYv6wec6sw8It9bl+OjhC+lrPAMKLqU5FKac7W3ewFuUY/n3BzVajlGu4moWXjaj
1+u9IBQ8fWsiGHIrJFM/xPYATCm6Oaop/EZ8uA4/5w1p6ymIBszYrGshEToH0Pao
qyfANRRu9GCPeZpulep62e4DV23A382faKW3YrW0b9V6f20rWphE/gPCbpAC057W
RL2w7bnSQz7/r1URPSsVmp6fB0xU1d+yq+FFOcBDgu77EA/ud/zAHKwUJ3dLtlMB
g1MC0DgPcAradzfUzZDvupX+g/oCraiMi1j1RHwoc3BJzIUrAbH7O+k/QHzT2XdX
JJt6LSGEovFQcwx1+e1e1obQq3G3UvzaEbhJcmYNG1NQ4VvPoSnVbWRYDLhmE+Dt
a8V5+6VIPdfEx3f9lYCdQmozkPO+i6Ev1whMYcS2bnKZBFdz04RZr4XiVb46dt+W
yJvus8PL7ncQfgAZo/ERHAJNt5Dh5nKYROD4OVzLBuHbZnpkos6V0WV7YchgFK5Q
0P2f0wi7l3ew3l/JUMOEbGnS6qgytWwEDw2F3DJfhTAtYka/+7y+or6B1dDAuYLH
oSW0rU1gVqK+piDBzPN37t6SHJaASwI32kYOqdJ4AlO31DmCWDqlCxDh36z27HIK
q0Y2RTTy7YDxM0/E8c+I67fs2YfeNNAe19YXbj4b06Nchz6NZD7LcI9G/yTn9i6R
Mhlr6EleAaCHdOAEkXyq7m0wDrLFPKH4/UY11Og6SPTWdYqgoM2qt4PLHkGBNnX9
THDq2idUsI9zevJQuiThyJLxVPvsQR2fo/eSRnHU+jT32Bg+UAtOsgby0vzmQ5tC
5pyLPcmcrjLqvOyu7nToE69s/QMu7mBYjoJGxDJQvFH7bvpd5qFrXXpd87xzwsqy
asCFhgNGwwLNO0wWCY5voXmeaqr6+hiPGLC/Tudv3Wq9YD78g1JthP+pe5HAkMGV
yrW7cwmqowLubvSBTZ8Y537/Xjo+3AY47wUZ48ouGDrGsn2Z3kofiP4WwycsT/Y5
8wQ4SKrqs1B6/RfVTWaQrwUK4o1jdP1Y4esOby5Go3YZn1F+qDZLRTe7ksMkeeLD
j3FrkvqW99KCtWNcG5+k41hMKtSynk6zZelQ24njFmswUyRj6uwBJaQCpgcMHOGm
FcpDNa10UU9wJeeMwSPXyyWMH45KNQUp4U1R8l4FFNUqoWIWEYNG6w78WGoogjHR
8U6vzYz606ti0E+1lPo/GF78WYeSznVmkrdPGuc3Rv/jPZrTKuZPnrqeqaXnkKp7
+eANBjOhwBc8KUYmHUOwTpZ2GSATugzseaPSj20utfO78ScKO+/KembxJOOp4CCy
+pGBmWjemcBmB79G5nwpWhoXg/FPx8LDFa/KMpU9sgIqIOah03L145L+xz6RvYBZ
oqBsTKUueWjHweZmideZgd3K91KR5HM0b6UL1tQyz7XHJ5DNbwkQDPhTZM0FiKmL
Tyz4kAyAjb0CbNxywUI6goA/a4yJ71wlRPvW23IAtykwQMjHQxSWUwIagp+vEUSY
zzT91k7tMtHBz+mNqfXfZg+yBsLvcBWne2rLFMWTTSHqnWztNBq96CXj5OIEkCgm
7Ze2jf1rApBY4EJ1vftJYxEsNAqTmLDfkceU+/U5gfvhqoviNjgrirH9BI/B7aJ2
U4Umub7clWMy/b8tDvDwJQQgfmUwlIMs41RNrC4Eoi8RV+AXwtKWu07yKNoJGe7Y
TtKm3JJiY3JZdU19Kc4wGeKGJlTGM2A37m1SWXz3yDhVU5B7BrBEDsQaY0kl6ktD
BVZrXzSp70TXuiS0J++xZct2INYFfEIE8Da7Aq6Ap8iGimF6VGOpTTuo1HuBfpUA
k1kMTzqYMNg8/iGac36Nbd96g5Hr8aU4+VMcvwGzl18vcYKPvBKZlerDy9JXsPqe
qgr9pxQTiy543vtkGqUCDsP4HHkn6OKgJzLJ59eLYR491rbeRZh9wMfIra6Cgdcq
Jy4ObhsHGcdctMLD57wTv7JMM0Th3JclyR/Jc37zq9pg5vF/QIA3gjtbcE2TssgE
EDEZ+jOT37SPca2MZsC1KiI1vl9bWxCmmzSnQmF+nXF+q7uwCKA5vD48yBbIAsE+
cy9XfQ7MoypwwFyk+tngn48U6m1n7ADKcLsARGYJ1lHYlc/c2kt+7EF8lsaUayJu
aa2yPkm62pwoYqvhfzJv8zloFET+8FBnveReUhw6O4k6OtHPio6ERD6mLOZO/57W
ZrPqFM6hiST5MKawrSTrnfq1FdB4uTzL+fG22LPLOjUXk1IbSD9YCquqsxK0OMbi
uc9LTCH4on/vZ6ubCz63wW8041KbFxXqJnVfiZns/HPm3Ci6RrtbADLddN4wjmdx
GVTQ97oxbqcdpWyJz3Tv5xhQ94KHlqvKzAw/vuQ7quK/rsliJPyzR5MxLS7Ib1vh
W/u2YvwDozfvtk2M+w3Nn1FgcGP0UWQZh6cCUqpbtrudzAnyZchNx9lNgICs+fsH
DA1LdhdNcsUjwfYv9XPmKXlSZj6YKi9AlJbeonaWWxRZUZiHRfzz5dz+NC+3kMx/
vvOeX1bv/hjjZi4X+/lqmoYR5RxR0oYZqhYey0tV3Rcffw11NO9Te7vM0smrKZT+
cTiF7GLqSk3VN8RTP5w/tq5syCnueueGFapSHpP8UtOEDV7STF7H/4TDxuELaxo1
UxfmL8nUAWch5htwtP7QcGRO4s5PZYASClGPM0X1FgL1SnFLscbm1BRYrmTnznI/
GmCmlXvXbkitX8r3oAlLPzksgUHf7qK4xrsEV/jhIMdK6jb4DXubB0vZM0MX0uvu
dT/eODIgD4ysAe5Y++QQt3FC4N5ogI2HQ9+dAV0wn/qr+U34orCFf9KBZmPd6ywU
se7S1JxskB99RFkgDYU/IXkEvI7qpLTqdfcqI7tYdrt2Xc1btK3WAkq7drYHMSUN
0gNmzMOMClkzyESJ1YEz69dOutbzsvi8WpCSERGoDbVpl57H6X3HjmGmucnXmLEP
Kvkr/qF+e4N/wRZZY6WFiOvpR7kDkbTEPSgKAheiYzr82Gp6pO/9o47OVgnSl2UP
IKVLIQG9+zx+HqsiaKkYqBBsdnDdxCERn5T782DAyhgNq1CYHpKoqiHVy5fD9jkj
M8wqlOYbfiAy4HyBiA8ymIWIxdgWD5jU/FKUVTRZfwHcFx/F1saVLdoNo9WpXXQt
H33MvDGhfe2KOFCdYvAQuGK1N90gQgfpaiBGGrIs98/GPl6edYi5O8ftRhuEqTRU
q9uFDdQ/0anm7dVYv1UWX0wLsHhr85Lv2TNmnKxhmAJNmfTag0zox/Y+Gu7bCxyV
M57pU20Ia1vOzdR2ucbOILOBt5zS3OowRhDlfiOM/3vqJicjLLgXvGkvANwmF0+I
ExxHvNh1au6n6aO57CwPQxVqgrF8scaPXkKr8wjBoUUbRJsvb58EhX7WRAzUwVGj
qdl5eiETrrb5n3P3oCfdJLQSslZrfOKy3kb2beIAoP1l/gypqVaovkkB2k+yCCx+
A4fHxfvpKFYszhpBSRWDpRgnbFEXxxQMMrUFc8H0cpluPMi/Dhh5xkST1XKtB8+Y
qqQjGMoZ8yFr4i1HnhOxlYixxzfQSXZQCGACKSj/wrQrXYPGqCx+VALNEKpcWZRR
AjrlLk18fXljHPGKbq5Iz0eLF4hAo3lsvN7TTK6WZraRIZ4mJQ0RmaLE0UZoe35r
6d9gIFM2o3pYIc+gu4fCE3T1OY8p/b8HMoU+7ziBNpqhChiv7nWaI/xduN/YQgfc
DE5N5hpSKzuKdWhF0YryZhaqv44NHWOpm+LKrqNg1S+VjtEXF36z+2RgXWq1legS
Lnn3YbQ+fU3XJ0eJyv+rFOMJRGXDE2UIsuoYO/geGsPSrJOl7wPNKYG71o6HZjMB
GemyjlZkXwERqZ00Pi1dU5BJ5qutsJKpgXfXyn5HahqLu6PPThWV9X+myb0tWMm/
rfG4NejGXypi9MIcoj8BmT595upVPGhX72GZAsN3NzW70CaQDTmWRVjArfXyMvEF
c8xAnyiEVBZ8sTBDLHnq9V5w9GrmlF7w/XZLzgeU1qSmoCz6g3D4IXl0fViV868C
piJGPzGkV0d1+Isj5Tsvei/NqgWmMIostd2XDr0iPSDcpv7LK0tdXSr0iFqXvX/z
qboNCg7IG04HNX6H2zHle5in5vML1NmUTHjdPFLf4AIL6UMjqYHZhLATm1xxtvlM
tMyPFI2BtVU87pb/9xQZ8xvGGR0LpnkigfWnjxHj3ZGg6Q7Otp1soFeDcLp0QFca
NKFZW4NS9K7/lCqFaOhOt1HZZn3KFpXzifmzbzmc5XvK0+La6xqM6/r8mGx2h+U1
ju0dy9pmz/QlUQyrO2SXojJircxusnP3OclOW2rfv11AA3a4gO1V1d5P+vFfcusD
x9qMaGtvdNs6Imxj2POHCI4qZCKcmc5s9k092vII+V85DLHrBrdmSbsnZG5D4+Pm
GxuJJFSFBLuAjDihKU1PO04X5VPrT9ehvQlleELZDX2/yuep5caMXE7c0rlxTH+C
IhTLRC23OampoFAXZqlgWoeiAZ9wTvBS/ZarV1HdsfkUqtzyIsrM3SKtoOb26Mjn
Xx+wKDa7MhqXClqbJYWSyhkDOS2VL1aJo5XgcKRWvX0QoBxp3yZmtPQ0fGcAzxxW
F5xsRyjbuxhVFNNQ2BPjFb2UX3k5K14zohrh0WhyrdK4X87h8Q0TdhYKzMzFGkhW
2CtCOEuanddn1wxREHOJihpAtV/jsSxlieI22JmPrMrT2aUKEhZtotalwLNBuLzo
fOSLZTAMSRTKmmyS5sv3SkOMxTO7JqLshfnsdjprstsYpXhFiMcQuVttMhliH/EP
0Nu56WYdPbz5o1yFuBOJOt3VOSVfROorzv+CUlIjMjtym9KI/K/L/IDdhTBfDTsU
a8SieAAd1lQ39blKdPmrN34iRDbK7zosEAxeHDpA0N+WPK6beyzB/wZ/HNc1rqLR
+hxYlGzR/d3JhAtHyxL5RI8p5Py8oin7vuKrLvN3RFGFTZ20OiZf6Q2aJcXWRP4l
+mlmtShIGZXQ5IKUlRFc3wyleKvaVAXfpfnmttvNWiKrLO64wL8QKFqfQwje0g1Y
w7iEvHdHdhEHAzEwVozF8hEHNtqXXt4o/fX6YNQdHRjxpIPU4sGov1znPf0We19T
AoMezGgyQyoBxouWfzEwiTGxb70P6BxMPXW2/BtwqYLdy1SgrI6KeBtumpFUefQ1
0pEPoA2E/fqDLj6IpPUE2ss4OHY4i+AhclVVwNZCnEXQCmm7mOVRKSkfbs2NK32q
EOpISk/fsR2ire0t5Rp6caz+HCekutgMktOZ4q1ezR4rJD+in+DkiecNbvlhcRHp
z8KrPS4N/TWkqBol6HgPcEnMZdrPs595qeETvzJ9loF8eQ/jfXnd8sglYwQuW9pS
vXpkdLBCbWiMh/3g8PWwyKNtQQSFR3nxLPmOC9gljhXKv8RtAODKnkWrUJSzUafj
jwCWoOF1diqVsA5SFTojW4D1u+wSTowIXEk/UnYHTKMKJI4YrpLrqjb4c1VgZUxb
axqcEa3nebRZVHt5scSR0lJRYVV4jXSqf55BiaaKBrq0tLPJyEJX/eufj2M9nSzn
4gxGKrjs35PGcKt9GcP8o/hXr28huHhClpK9gdNeJ+tNXRujyKxKmwyFu+oUAKa9
y+ccEbvnvAqd7CrlPR3Tngysm+VMZwKpceoqXwFqa7u/llIDNs/S+XTZ4dLTksW1
1a6mp0EAoEqvgzkbDkoghzTer4OImJsderRGeRtErFwZKIh//Ih1Sj6BC7ozMHV/
bL44t86sMh6YbMJGBsBHyPMQIgemO+tP7h+B1NBJWEI7AWAL01YhY8+csrIdSdt6
YPRYOsBdoj+E2ak+X2XDRS7zf5KztjdwVDHbFJ88ddV2OB1wITCGtpAYKUwuzrcm
vF9unOIgEfkN+DJoXP+xvlj/AARJad7I3r0EV1zkuZpgyrEZyxulLv+eft6M2MSy
2h71+6NmB4JpvOCyWuVNg4EvoUt9sSX7LpMCdrx+hbreXjRpfz6DpUY2LnxhQxaz
9KTC2t+IPBHka7+LMGiTG/jy/4KwfucTehWz4BXDiidFVEAzqfhT7y28Dl0/0UUe
0EGL8lP1UW5XmQ5/xIV9nR3RuiN1dd3YRd1i87n/2CPyhwPyBHxRLuBXM/KJ00Nc
0gLamsmpUjDmpspDglG3GhFIjZ2oe2o2a7tC4UeTyWaYh8dm3v2cjOzWXrlq/bPR
peBJIGAWGVwxZFizuIn6VQF+TqocNQ0kX+zSRuxD0knygRXTMa1/3SjcWEwOaOVl
UsjhPZf+cleix0rfAD9nHdDJKDXnTEzOSD4eRbOmimgpW+5NWnG1AenSLHsUZDfw
tL43kTl3JaKuRSSw5y8Sj1OmmWZYnCCOD27XNdwjk98sA9k+aUvAOK8HgIGM9oq2
g9r9+Id2mX7mSydZCCGaKqlCNo713Hdyrg4OjBvQy2qVnCnOqT/q9Xks389Sh51Y
iJwtdQ5hlRQWuPLlSERylXhkwPpmwDtrxXhs3u5SHMrbBmmRzMqD1L3fZpa3oexI
WdbebSsCm8zEf5niSUiqo0qAR5y0qK0ZY3yIck7/j2VwKHSh+q2UUmyjOLQa9ME4
AKT6VYrKb3NrmZL4XWEGNz7hby8EqtMwjMW4qNqUfqqzcHLWyeApArGXmzweIzwN
xFmYu81h8rYnK7Dh1X97P50zRK8ube5SjkE032dJLfCNizq7iSZox9zl1AvEqTkM
2MQlgx5b5HqOU6u1xT1Qmpe5fkT98aYe9F11fz5bWwa7gG034z/pg7eLDemxE9Fy
xG5OgHc01QM48iEiifYBjSj/o1q8DT45X5b9IgoaeRICBubCYj0S7MWHrARIadfb
K6aj/P/PwOgYQWwqwt74pVmbs9F1wxkuviKT49kf2QOjCBC6SPfAm1ejYvWoud7X
VVUelEYaEUHAAutdliDmQDnP+2xPSyyD/rgRmra2/y/1tk//zCJZNsfawYAzUDYF
4Tmctkinr5WsYLacQMVUWVgz6dZb6qRt8IaUyg2TrFJ59Ccr2Sx0bCeqKOei4+is
CdXZ04UjJm059VW2KQ8vq4mkPqkks0rNCqwODaCSRTR/e1rX5yd3i5JM0XWU2R5m
5jLOiPVoayOrSOmfB63u1vj2bs8OswWQ+WhaC2Lnm0n9G4NPq1hKF0He5T1eLWzZ
J04TC7zxUpSBbBYWFS0QskU9+2Nv6/L+nQqOCnt6ApOplaEt4y28inqlD1ezWXh2
UGaWLdq+/YJiwzelAznE1kudkpokg9J2mXeqJNznZvur+/CGTSKKGm0l75PjYpRK
XoLJ9s+7HfNp/IbwsLxoJ2xKbkbqOaFeQUieNceg/NglX4kk2anp6mAAk7gExcOV
+upNTDKZJzm+gG9edJtmtIK6Wdn/FYsU7FNJubO1rDtyXHYAMHzBsx4TbelCZM1b
15ZA0o6SnStHC7o6+N3HfC4OFuh7J3fJv3mPwbU33WVM32S20EQZwg13W+A2+HKL
bmC4Y6NpyF3knlxis6nYr2mGSYTCffAMWf1PAb9sMWB3cnYZ68+q6VPF1GrzI6h8
aBOMvpDDKVr6oDOgrw35CNvu85Ez2M0zoZbNivmhIUuk/0Hab6u9LoiK+lAUmj/Y
VwMSoy64Y3dOnMDk2dX/aVyxEunCwqmXhc8NZQOSejrA5QDqvGCVmUu2Xj5mKZdY
dtYEYvrGTmW8v7BV7AQYAJbpAuArar25dCLXDI8kRXmfsysGo3wceZEX7u4epf3E
1KwCY5ULnkkK4RPHJK/HocJF3UoFTgTGhlPJcnm/HEkAQsITc2EGe24aCVHozcIV
muox/zgLb5ORU15akzhGosWN9eC0HUTOXQFXu9eH83thq4q+Ng9/8bjByWuRIo6I
lflVftnn2V9jkcucS7h/wCpYADaP7NCmJQ7P34UrOEstMxrlyqWVZc8Pzyzf//qV
PXU2ZSbRd+u0t5hC0gVSmcNcOfD3SfEbcPWPPV5AVGVpfbkORh3X4eI/Pw7J8ULK
b0jwn9cIYzkD9k3MXHcKr6xc9UI+lEesq7+xQM8tSdHwoVUl1Bw3PgiRxQtYt4jA
ReK4cfBNuTmR0TsVB1YeHvkF9Tdsj9POKGumtF244GwaJtPLweNr5NfrKu03TMYS
ed3l1qAvV/BSoUPAMlP5elyoy2KtrzcfNjP2TNnfDzoulQAZHBJxC4U2K3CDYI8f
PSmUFIRo4xic//CFoEniaJsDEqjWIPNHSPx8wOAi9ASGF+x63/S97Ibox7Ch/BMA
ls9v+IZ/qwAKAeK60M4XZ5HP7gXS6FVX8bmR/SceOww3+T6qqfT2bHkDAIdJ/6h1
2Ks4S9JTssGq8UgToUpJloefKkhmk+WmxO10pJ3k6y1Qu0Ce5oVD4l8A+w3rFPga
P0cst74rybUL5Ki2kyhY0vDRGZvBrags6L0aB/EQGezLclg0AM38wrmqoNSS3x53
wiPpRp/OY8QlsDXzFRq8Ch1pPLRUaSHFHX5b7jY2lnWc0AL9feQ9OI0QKUVundZo
e9snoDz9E/G1aFHk1AQBdwJFR5imLbmyWdLjFc7+i1+sxqO8BH6lfUNWOSHJYitt
9szuKo3GDdH3dPhD54Amp6puEWPIZFwDXpClliOaMTBKlz7/Jqg0aVRxrIkkPG9W
5DtiPiGK0kWr3cHgeLrfXWrIXo1EeAIa0OKVuQSBhlVX6QC4oEvJzwrMazRb/SJ+
Nm3GTWLkSBSuFq5ScazV/PlyH3YfTaQZ7PJWZy+d0xyBSWnXVWxA5r/g1yp39iLz
gFZIBpr5ZkgQmRH9vPTqfVhE3gTcUBH4nzIR2c0hGOfkUKSmLAD1BCGc6/q85GOj
6q2Jqlr7KZQos318kDWIqAJE+uoIf4EwErlBbHnosF3N7pK7W/JLpn8e9do8p6xB
2XNaMa4aVF4/3wWYWSL63RR++bIvJzwZ/gGy/vI8XvRoYd27sYFvLyxB3I3gr3Jd
f9N2S7Ec05Rj1/w2g/b4FGhYSA41KA07gCOi9iMh4ONPjyEz6zp6jBh4VADDKw9L
W74ipuPF3dl21rmpqeATBbm5C6RkebdHuQ3uOwPMS7yx7N17A9h9BaGITKmHoDbL
inoxCDxXG/Y/0l6pXtWfdIRML2QDAhfE9BGPwKcXbXq1MmemXCbstY8JtF2Jkyng
mYOyIvYrDTsJi+2fEsy7c+5nq/yHup80eTHcD2GkFJLAkdyoSK4TJ36k2CnGDFMy
Y4tMrtcf4DsavPQUuAy6s8mxPkxzMCBFukz/kcF8TQOMU3lU8OWqrJEtNXYPrCwb
yqSyPpgFgd82BtobG2LzbH7En9NBn2j1L+Gpq6F1MOKBPVeyWQ9DJ3PMYi05GFLO
SErbQjiRtEI1P71FosW4I/ZSFcMFD4Xp3dJzX6II01KZvXDogxZ0EyKgJtQX3pRz
Dp+Pwqc5qre2gCUB+hszMRAC0aGwfhNHjOsv5xExxonviE0e+wc/tfrI4KkZAfmt
uhqZ+cwIskNP5d0YLJWbuq4fxhiLB1af9BakJ5hqAuk5uk3nmmk2hkJvVYyWraE1
8yM53n8njFbiC5x2wuKtlGgRH0otw89WKj9pug/3NCCanSuyy2iPXpGxTmG7+LC+
8WyZpLKQOvMICUCGA+PtdEtSJ3FFAon6z4ZjJaQBTOqXm7qd1+K7mDhpoYebsADk
tKg5FyfZ5mmvGjpr5YBdLqDJH8sJP3waeVXsvFx84ldzO26ypXCpXoZUFM/UQ/O+
S5B3NFcoi6ZcUokW8+5yHshio5vZFXFTXN+zMNbyitgx0Isf72VBQa3kkDSRDa/U
+t9dKz1MexQDp+lRIsAwcntxWG4Wnp52WInGP2R8pFfUl26bF4PvbrBqm+qnFBaz
QGefFhn5S3a39hBQS4Qb+OBgmTU0gXxNxOWRyZrURkYrAZuFlxnvk/djeoa6s6WJ
FMx9qLLrUeqI3ElWJBEhW/hPHq1k6cIR9N3AUGVig26ssmys0j2hqToTZnaDBalU
FUBjYf/hK4MZ7OoqeIJDYhMqX0+SZ5hzCS9k65eZf8boxrhuXOnOcJ8tS/7z0ROu
KkDxO1QsvY1IsyIky2bKLyTM95dTMu5XM+rBMtYGYqodTESgAclG9iPZvK43yTDd
23sV1NcC1BXh6qPzUxljjnRpc3tzIEildc9JmLMPiedNLaYXc1fyX+iXumLw8WGk
kaZWChl5BMo6GQz8COWcekybIe6Gvy+Jpejc/XrGb4a+PCmq/KvXt4P7Pi6PE5ME
EQz7RtYdKnmytMyOSuf0t3SvRkb6uiuM0TReHgrJ4zTHAFp/Wf3QT6mxcs26N0uG
A3skDUajc6cB1iSReHhomqo255XsupJmDjrXHIXrJPvr8xv58aKK1TlxmO8uCOpu
tWz0gc3Ggq3QRGESajpSWS99jdgdLasWr1LakBCGE4PTRMtdUCUezdSRwbslJxUO
LFTWX1/WFAC7A9xK+kvNf2U2Vm4Om9URwUL3OblJaWNQZHe3Qz0jUV329WdIyu+7
YdGpB2QT2XvSqF3olsp/ehRaQMaRPhNBrey9ir7rcVicf/30uUapOlgoViuidiYw
p5T9lwDjQVvzv+EAcmVgCSg/Q51wv10J/R8hXxdwfO4d87nHbIqQzlT1GPjNyvdL
Il4kUyOWJD5Nr+TOhGwq/4l5ajFkJMyIlvaxJrfK16SBY90laZcREHPvuRcOg0QD
afz0mrQhn7bsw4wnzmmyiPpWdDQYt0FpnhhBDtXGauduSml1x6C9CdhlK736NfN3
+zL72UJfJCQpHQOJCxHfp4g4srk3mZeqQBW3fRphi/49mfwGG5wMqpRI22AZvuAj
FtkYPlWxybvaLiudNLafx3r6l9s2orza04pRLaxpFcZZNKp07lSuRFBJPBEKF72Y
S1qCGMxcXsShQT3Dpi8LEYqkK95ge3m0krWOwM3rdLAxInHRPYIu/kM6uGiSQkt3
NWtAG+odBx1nph6580WkMFcI38jEcsYdrJOcqkPBg0RVQK5KULReDupl7r4aqrmB
QL6Mo+USttFCub07jp1SVTQjtEKsLxpoxbo5yfNactHUG8dByiMvOpORNRaJhpx9
nao8kFzhD1b9y23tahtxy1N23kiTVA0qW05jkIVL7NXobxNwQ4Ys2T2nlEdQf/Ue
GBue68DoHpVMwqqwIXzcbAV5ssmQ7SKBJ1/AcZGNieID7cec48H4eTF/emFB+cxx
MmNEBfD33VUAOpscf5m18ammGO2UEDfdeEfAiQ+fXCVm4FQ001kpDAR0NOBpB29B
hVHnN/FVMsGfZhMjCRu846n7xi7w+iAT1WFLvgY8Ovqy4Bqw67PL5lj3fU45dqd1
w/SfN1nl+y8Hsfopi8iR3TjGlFrEbVESXyvv5/sjAQZ3kYXFVwBh3WcD3tUpky10
uUns7L/Dxs2yNE8+asM9luCVBV9pjmsR7HYOb5vevjfi8jHGqUb3CTKo/KAPb8/y
Jvf30prJq6jtFzPfw2vzn3Uddtu7s4/oKDGD6+HNGxRgiig5S2kLbjxqFDmXIHzY
OBwntiphBYDtowkk4H84WsmZVYoJIlcqSg9nGbl0LUGGR3QV3MQqc7bywYt/pC5N
09zFa4bS4uf5W5HnSQNok6NLPO4ACIQ7avwWoXV4w43/SpfreE9qVKlzCNd3mNRW
7/47Mec3Ayq3LBxDqkz9112DHU0sUprtmSykIR+oy4HPc43BFiGbRemlL1iVW9Vo
FrcrlENz+z+ohlW9rdIX3VgPa6dw5Kik1EuRO5ZT1hr0vI6NSzDPHkEfjG+mlXfP
gOioGZ3MnaP+7NnIbl9csZavi4N5k0IRuiaS7ehs7RtsGRoJWFLILptDLesJl/Vo
0FqN/C6NWWvcfqn2fcC02pyRiX/vKJOG60qAZoUHiArG4BGU2rK7DQmQINkveVRn
oFqafwrzexa734clZq+yIYPxsP1McsMa/sycYts1lx5gvaYH4fXdDvHSxwkAzWWM
35Loa+KrngIPMyEGlsBl43ehCJz6VHae/WuSpTChGuMOhEVa5PrCqgIinM2Tzn4N
h0ZS0m5MrIJoYqUgD2gbd9NOavFnHIgqNnjqpsjy+rHMf8hik4nsDYN63ZL3e3R1
m46Zj664JCH/FOtZZlFLQ0/51gvM7vyHVFucQ3aIfQmmkjHqhbebdfH7B5LMgukg
l1JGdkJvmsWTM+2wtG4vFjyT2v8xiCJWUvoUOChnag8cBBDPhJRAZ7BKyCzVM68E
tGyPhk7rv2wMKW5+dMIua39HIbKohPs+EhnaMg0WvYE19VbYGp87S0BQEFBC/VFS
M9+IlP8xPqF1EX+vPtIaga/8rzidmAUN1Qbb5z0vxf3VtO6TeLde/mGTiITWTv0y
2UGhDwo0cSinfF3USHX+orIKf8eBMo2Tokru6hYtG1l/2sR48PMwSfeaUM0fht4H
aAr+bzy6fpLSunzzq8/aGvWzlvHFUGs1sX/d7XvwUYkoI6UxLSRKGYweqBbDY/XU
oBpGNlW5wFC53PupQI3HY1MXCSrH6KO0BOlURhmu++/pVS03+ktwE3BVJkjj1mkv
cC12hjvvDjD+RjTHd9NE63QyfABPRhzxZsYLAxxlyIMTFFb/pu5awAbzAfC8TzKw
zN2E606YpPi+4OaMm6pcJpPfuGBbmF1ZgUA0WMP2TzV2mvQDoMMBbiI+btsx5+Uy
5arWmx3jrAXRqBywNqfkrIiBzumZNIeO5f7uldu5R1R0PXgq2HsiKYfmTTFzFNZX
qMg8r9RzitRphJMrgiQ5fx8nEpz4iBTds4+hvsql2JiJ0dn4sVXcPF7J+himk8qO
kP5uz51tgzreF/KsYZwqMgebwb7ENRYwAYZP638nMszms0xMBL2F1FkD7P/BXFt4
kfZ/7MMS2ausRYFrlFvedvpwvqSbsCpWwU6DWsY7U4wYWqNNSBqw5SdlbjVlPg7W
ZrpG13+b/BP6mhQsvUe8VoTca6ZckRLoxO3OIkM30zzfEpDjp0RWzqz4aVis4I+4
0vf0HUSeeWbtiyP+rUo+v5bDFhlu4XGujYLBLqdhoB5BUNn7OvukO/zpxrkyKE82
4mUo0DAxMZJrUXah8Cys1W2O/mp6RB6K7VnzrDLMHwEj/Ft56Zn5ymFt9KduIOmK
RfFf/xU0J96l5Fn+2qkl3cRudTT1mat5VC3Qfc+A0JkqGwolaRxx5zjNehCVdqB2
RwTIENT2qwfNjngmi3YLJxBiv/Zl5yrL9c3VLxL5V7mK2F102FzWu0No76sQEta/
XXfeUE9zt/Ggo4OBmvzUqKMWxyGRu+8heH+/b6Msb/NdSmSUfZcHzkc307aAMLO/
8qVQzrRNyhAONsUXfjpoEzMYVX1tT5KBX7Qf5bAgYKJ/CFLksEC9MMaSFw/o3Oq2
BuWap/J3B8qlFdOnUn08bpbfim68WRLK3GXjN23Mdzn2EH56uaxJXbFFTpaW9Gr9
aM3rCqQB38YT3IxpZVcEvs6hBXtzt5Cc4iqsUWZMzfX/xKyD3iMQL0ZrBl+MXtNV
H9cziuTa4Cj3sR7fsE3sRbFIGsbd5Bb1tojtFmlh+IHi4sYKlHP4xhOObK6YzNeL
0HscJrX4kdpPjy9yrUdI07x3chvECPSyxAzUm4PboqhiTUbj8OpbkXaobumhOqNy
HMf31O1fhCgk0GMj/rrgbQHaHk1NsHNLQoWdUMGbkqmNk9s4hItX08B6eLtug7ik
i/4sn4LFA0w8l59N2x7dJY/vEE0ViDnFWfR21g69kuRxADVhpq1sXDlrR4kRf2N7
CdQD3NyjubLeEOyf1jDn8HBPZfXD7bikbmteOcWDWTjjKWowbDUXqIOHIXIvMCDs
MWf59Ma6hND1ksq7pXOQbfzVwjA/pkENTebOplvJJeEfJK7Cl1F+5q8yTMXl1nTg
rxFs0lXTSD/bMxrvAmlh4z4ZjPONwWV6GxPC0ELYbQP71BNbYdfegmge+ZyJbK9K
E/H8zImKT2ZH5wav1377mXHNZjCquz6JIxsvJ8SkKgHoE6icjMVmEcyWyObtEHMC
n9kMcsBoLVV048TVH2Uqwe4X0QSMKMQ7n/dL1nsjUMxLUagOxk6B9qLxuRQCPjXB
qgWmPwg/saeRj5H0fnG2VXcPvLjp01MHiozREmBFXuhDPSO64b7vy4Jqr+WkO/vo
Poqr/LwGtDH2usl3mNLuynRVE3jLjbRHvRIWljlOs9CLk6oh0TNVMuxSOXvMAFaF
ZqKk51LZwKwCQA4ONghQGl1vgHvXuIk62fvY3Q8SUfEcY0TiHtM4QFP/PQ5/gJeE
n6mcRqnY+gF0n3Oz4/ZVOOZm1lG0XZlT80ipdUNzT+Peyfwfi9wLTrryuiyl4Kxm
rygdQxnPnvGMrf066pLjfsBFODSW5Z6QQMQvb5mnpgDT/GahTriVYXiT47npVmsO
b3L8lxhxeEg+M8IhYCEFhhknQQfvLqOAqiGcYzbqPf9Uu6mpe/1OR4noGAdWAJvZ
V6/W+o53HzrCfWp9O+Q/CSSWhMOCWS1girjpKC98zvwZw6IBZdyEvS83TGrhIOeG
wlFKPWqBFFt2WUqB0XrwFgg5InrxqZdxravgxUIWAS0UGwVUToQAyOsNV5h1WZX+
syQxgSjjjrGSg7hp8eF0LKtMU8ww9Ld8ISLFE6U8mr9D0lHheJIGvzGd2PVr71hX
8BL+PurggMh/3EEhv54+W+4ryVJ0x37TSYuYB1VQQfPlZiGmpXcIHBNmVQbMVvYs
nI4tATxdeBVKUnbgCRRt5jCUg/7U4B78AlOTqRLoqQFJuyITwBqFsDtpzSqoONO2
372OzCqcCVGwQB6ZU2YspAJGnOEXiCjoNIc/OtfaQShz9Qjh2D/s9J/wg3X1tJfg
YfNKnc/N38YY5NPYw11/6EMsKHqjOxary70m6cUzlUcosWPQS+QG77OIgejhyH/B
1pZjXpfaMqoOif+NJtXiJGUG3GpdlLi7zOnpq254KeGQ8l2C+LhRUXYQEiT+uvyZ
Ss11QV+yXketoNyEXRjRPAY8o1JU3tq8ZzaRAq5pXakEx3T5s+exz+0rYw/e3us5
OCovH9nB59/QIKfV5j7S3hf8EYFvN8eqzZFW5ylfLBoQiGNo2SxsMnZKh6Jwz5ZT
vEHfuuRlVX+fzeMiwEkba8vQS+mcO3BywXzdRj0+9wo7kUTgJzOJujgx7YpwYA+A
J7/SLyMGehvhTZsUF+Q510Y6rMHratjcm5PH11hPR/J7zMduyYep4EoeX0ZMEEW4
6RhFQdKp2+wNsAFD5K987fMJVZY+jrIGhlaRVEZFo39MRzQQ9sa23WY1lvRD6MdO
hl4shwPIf4riBtzULENEH16ts5Z1Dnh12S0TfazYd66G9D0/BF6LPEdcPnuW+zmj
w1RRQqpux19uu3CWVk+EaHnLEjMvtiACuFv7QEmCgkD1Lxc7aPsBGIDSVHe3s6Gl
/ZyMfoPaOiBQk/fBQa/3ttCBGws1EBE1LtRetXNNJR/Qo4SXYa2UnRs0YghgUvTZ
ovEyOE36w1+bX3jx3KkoAaQWBhpfaaiALsTbncYOez2MyzJLXGWV081HfGYGQvUg
XLxd+S9MZD93Ub2DeUgABLDjJCq1M1I0bT/Sdvt92v5JoDOjxFsVEmWkwgj4Aq35
t0+XygcOh9BCmEZa5D+dT0tU6MEXjxG9znonjYehByxelC+Qs6UWQi3B3aiui1cr
vCYb8I2I+348DZb31KtL7ZAwFn3N8Vjb50DIi9MYLC19fxVD4Bhe0rWOXBx8jLYx
qjbeoIdAy39ZaiY8eXEDWI1D5FSs8FPB2p7h6HB6qGrRM6+r4vQnKTFfJBbwspck
sS+wGvFYsrW7cwZaHcj0by7zQNMoxQnRQ4PfJyvxBVNv4tZ6iFqAMOYMr8eBRgFr
5rpT/0oY81ndmXWBbt11EnnnOhZZPwgNBK6itv0XaRcmeZkq+au9halwW9iVh5A4
JhNksPDWezdAqJ8e/SmUxmJf2Zho9m6+NtAUgp4CNu90yI3rYvcuL1n0VdsZ9kfh
o18Qm4lVxwAcm16CHsl8NR1s78CNN47QUtn6rLEanCskTP/NRabq6UhhSiiokglL
7JzrGCkxzp8hTrDadbT0vzStFAleqXCJs9TuiPjB1JobePeqwpOa8Wspr3fRB8Ij
sAOnNd7hUiaQIkm4BKmIQwo6va1w6Ihg49rHbbAKBJNMd1a/DXVG/+SQ51s259A3
2v8dbXkpGQuGIR5BpMstPI3Tj0SBEpHiWn+3cK0EOM1UC0a+PVurwSyKtNasOMFR
TQ2ogmgHiqurdpU6y5aunrbCpbfiMMGgLkl4ot6yxGBaw6SJQa2V7hR56iKRr3so
qj5ngD1zOMg5pRY23R/4OvBIYmda6bTAlOBAKQWpuRDR+562lXLsewWvlFv/XjG9
Wr4SdFyrMXs2u6ub2IvMlb2Ueb6aUY3wyWQKaqvDY2zwQNc4jkKq6pxhED6FLWgw
c5zyUFo3RcXlsxprJZ0heQNdn0X7smZH2UXub/UCHRSFknRlCD4UAlw7pLntUjsb
xAyEZKEQAoKkEzN/rYzZ/YBm+oKP0ciEzgtCCpk6oWX8LwQbPcJn2gRXZZXynQNU
uJQkO0ShIxOw0TAbm6ims5vxWLfWYQQsgYUWujT6eHM3/FvV4oxdfSuwlhxObif8
s6TGITTVkFRbra9urcXgcLkStWrWZNuQqksqM7BSv76vS7Xwf3/ihHhN3syVr9c/
rcImzclUyyspf80yTBKSLF6v3b5+/hsGBzGe9StsNJDZAusJ3iLrNIyQyTmQcn9E
UXO4C7Tg+Hn/hm9g7LueiH78Uq0BIs5MtKzU2LrXP0UsKC7KatbNwYU81iXYPjcY
P3q0vqFMlR36CXTbtCvlrVfzb+bYWleiDJ+CaxYEoXOJ5TLLLvYXuHA1+atYSOGa
DjzlzqP58iL7LDQ2sX8ehVrZjSKSMfQDnM1jSZLjjWFHp+02Jh0aa0tKI4rB5Rre
AQQ7ex4g5MqNQvuZ7ctBcaKOQw5f6puDHQJfNGFU7dCr2gqjGGREXSpEIHc3w4O0
wk567dCIM6L2MzUYwdE7xxv/skux5aOq78p4RR9gT6VT9VOoSKgdXXJSEfkDEJcD
5KYo13GwgdFTn0jgMY/pD6S5YB/bUjU7FOl1QIspy2jTRylJ1rnXA2a+Qv3eWPo9
BCXf++kS/g2UiDmW8xYKzOssW+FQRoyJ2XRtDkr5JKQvNpktac203/cuLvMK7/80
vW9N+csdxuIbRAiRDJOmocJZn7uxGZohvlxam+W+b5soR/Z4bWLRQl85uNddxoTY
WSoPzbZhLu86q0FLoNZGvbCqAFXRF384kwguu/0e0Cf2oV51miKYBfFQwe19KRtX
0cnK24efVVnjom9BfDqY0HjY/2Rgjpo1ml6/euIbF42VL7AIp8OFOqjrU0x6lUPx
FMfBkqlMP8mATWQHFXfhriVtNKqJR4jittKWNpeSJYU9Ynu+BsMVKdbOOmFSj89T
IKjErSJgvqVsW9pMJJv0xMhzyD+fH9VFzBevxWd9wD/BsRovNe3bNUlJm6m+/LYa
BZsQvwpccRgBJ/pUWFYuXWt7afwOWdSz83dvK41yEaIyxNnIqZmOeQfVRAHLXKPx
TKq3FmN33SEuyMH+0XwSUt6xWA18m5RC8lXZ+H9vRTmQVA9JggkpmwQn4o6vkqMB
HpNZTLHz4qOHdxMJ9vF/xjhxrsXeUfdNI3c+2wi7x7VT5ec4c2h/HEJhNVGKCemM
T9rJ2zUl6q7QXMAAFNwDtfOaXZLpJXGoOTEmfWY1X4FKgY7B4fPbP8i5rst2qSse
2WsmJwPCZ4aEoB7qoafr7izC6VvndPiZpKuXBDHER3lu0oHUvaaPLXvKhc49EZJ3
pGNSWGs0OhRExmyhauuyXdIjZ9SGMZHfwk4YguBx8/whX1jq5y6AMhmSum2Kes5f
3jpy98f7LOdXd73Q0nqHHeZ9ZEN0DQFKhu6wk9IVzgzyL5xHfFtHah5MRNogFe0G
3Qaz4SEztIKTzQ6A7+CRPVowritdjgWrtvcZVnpAlrpLtvVFVDaL661KNHXTtAo4
2gbpMjjwEoUflkChkIhlHUfV889KEI0/R+gFP7VIKa6XkgHL1en6UzuhBw77dwXh
FDAvRLTzDR+fqdDgdMLreHk5/V2kD3eEuJmgHahKie5ktijWoDtmwNYHGPRPrS21
dT4uhAukLz96VFy2EY+1CDnjBKAVHBfNYwWUMc7V9YV/W3zvCJPVD1IbC+UyC3oL
PwJH59htMtfColipk8DeejsrXjf8dAeXZygymrsjFh5AsatolfU4Lynv2TbTPtLe
O+P173jpVgw9YfaJtS6qTc5eetaj8iSlMWFZj4cr2XsoWkWtSz+8n9W61Q+iTQew
DaYwmUk990JoCa/3a0xD8uTHd21d6UIQbhaSnAoYTpeJzqeMziaPhrj/i+CL+/GM
c9CSiwNOq38oD5bjDiBFXU31NmMt3cPl6iO4euIxktichFrR8iQdLL4rRv1mhbwb
vEl9ntRAcGqudhEYxbcUfGE4ogOPLkN8e4ucHTJP+BWMItz/SG/PQHRajLAMUm7J
SPpC+aIuA4kCjJc6sNJkvSRrLV4lLl3NfYWGyDA1yEMWCv81FaQqn7Sfotn4J4HT
dbQpnRCuNbL9hm4Os2iYMRYa2Mo6iSiETw6b1l5dIzqGC13LVnC+NEq2tidypFei
Jv3UBeGYfqYb/GN0K+ltgBmeRoeoy8MlVDK0kbVK4uSChaJwQBHyYJVmMv70Qn8t
7eeUX8qfSKciZ3dj1QnQ/rX67I+qX63r1/DiwtME2WDe3o97FxbdQcKY5vUwwf3a
TQRPQnqxJBz+iYN0gztNipE5Od0Bw94iuQNKgMH+7V0+y4x+t3O92+WsWiPk8J40
RZJTXjuUnTazkwne9AQHlMHfXpNRLK/U5zC/FqsDXr4AVWIXwavi8SMn4EzPADmz
6T+StzOlYziZ2cLK3TQr2z5IVT7ZvH7H04dy9lrJESLFHplq/whElDTwJf2gIja2
sRHUls1cxoeh4b1fmzAc3lKQZa2JQod1uMgPSOje43772YzFSBInr2nOCgkrdf3y
IYDgYrj1O97w+cK6YckDtXZCzQlskKMq3Z7goiOvqCNFOvNNt070Q0AjLhUmNwek
bKSmhkSG2V6RkbPHAuG5A1X6Oobt8vmATgs4z+3vnB5v5VKaUWEJ98wvwc9vII+G
W5npUb+Wl6F+WfoGNsaBZxo3rD3duDOUkEONB908Ct0uidFmEJiQ4CConSWOnvEQ
bY+QBIc6kzUp29coEfxIeC/nq4YLOuivgHnYqWnQnLd43RnCXdNyqaWT4T+2qAfu
jYT1+XzCT5YhGcXxwDT5HpKjEdHjV93HNMqtl8xI4lQie+8fzRGYqgSDdLBckRwK
am2dol30sh6c633TGl6OvfQnwTrMjfz3T0r0y5nvPe4JcoGVJ3kPsdwCkdm1yUV/
djS2Rn3y7tU4YdnRwjTW+wE4xGhB5c/mbuI/bkfZAoVqVSgw0yfayL9roHoLFd6l
0vBOd4GLk475vjdUF2xUkMzfbYWkvKvXUzLeHajUvS56k+c+hPszs1oP8bCkgfne
s6N2jPwW+ws65TzyU86AegVEQmFGmITR2emP6eqboKyr47ZBTtFbhz1URTgR+oga
im4MfNtI1nePYkeXAm+u6t4vJDVdU2SnT7q3VS+L1//2bphD0wAs1HbQmtWjUwfz
euxJYQujQcK8ZQxaxzRiC07hWQpziynmZj+d51r3IhxlZ8JlA2c4h949YuwlvRIt
d2UU1Uw9xnS3w6dLQLNjPrdR+ZPCirMjK8QEMaDWcBDgCwPMM4NztNmGDn/BJsRl
DqqHotDdfjsqsCbNswpAqTRpZJGaFSWKp4aqwRdu7H0TPJW7bJq+9RKSCRzRlW9Y
98Zf9Ut1Gqnx54HUebTWBNOHfZeGGhhY2Xtc378EZmphb5GedWop+YEJVBZGb+rq
S13dbH5+dMBudfSqNAU7WQA+zh1TpEiYvQebhDPvDCYJGPZD+dVnvd/m6TKlzx4M
4RT+6yh3SCiuEwINTzEu6/5bKav30A0ojulaBp/VVuK8BsSZJ2L+X3i+0cctdGT9
3LBPsUbOdbVqiU7P55z98O5W3Nv4aiNEjYRfT0p4eyBBGI5fsFmR3pWlk3YC5J1H
Vjm7r8Yf1E9qJ1ekExg+vS0hKIWQKCjgu4NzHKLDFoSSxh5fvn25L3q458dlFyXH
gI6i9gOhheVKNc9LFeaoNuvELYqaYdBUpJT4e7fPmPezvLz/XeLRMiADWkuh7YVO
KAkd2u1AOs++7AR20xIQVIgdzjaTpiv0fRa9XGGGGvDVu7M3we7sLae/llhmobd0
ytl0FaIUjXxjYeR3q7B8R1H1Bc33Fl2LtsstTg+Mm0mlvQ+ckNqcxLzEPOfvxIUG
Dx2D0rm3/s8LDW7soWZK2ZZMURjAiM9u2M8Na4KRFsoLOIL7u+noR1M2vWO8Ltul
SCC8m6Rbzs5lBq/I5sQTNlbbNE3InAaNn5zh1sjNPed3+Jn+Uk8VyyJEzl64NAKA
LZ2SA6KBIjglpoE+eda/+EnRepmEgkvzA0/pFzafDUcT+VJgzKhzyypCeNpE0BTo
z/vsXx5jC4mSJSKZoORmnXD4u4n8ZXwhBEbs6ScHWIgF1IcyGQ82cy3P6LP0M6+S
o7nVrQ0jJDp2hBSKr6YzhAL6tWr2+d4o8BsBRUDDZr+vS3vVEvIPVSaTkBMgEFNf
g0WY2PNR4cOMan6BigM5FKUWppQkoY90AUZUsYL+x/qaU0Jmukfo9u/3d6OH/NbQ
qXOq2gzGgglbkZfOVJs7VUumVqt1VEAAsgScQunwjVE+C7fd7Ukct+iHQ+NJASYR
NHtzycqouil/n+677hImrLTb/Q2dWGcCsWSw5byVT9obFoFKuZTeA4HNJULex6sK
6lSFMd0RicOMtdTLdSwZluiecRMWCo6tNtmY9UTUERByGrGbgkq8p3haecZ6kgaN
iu5uUfD3dnuMLMSAo24d+lEXxWB9cGTFGmCdgNJyXoMxll4XZ7OyUCJEyoLTPqD1
ZNLL2+7gPNa3ZAie/i1iNnKCXN+SpGE9MqsOh4shR4ZzOuAUH5gbLzTrAd4/9QfF
dDMR5old2jZ1XK8QB0UAJtOT85GQWK31m43VHT5sUhIjrHZAWOSHEwTWjnvtGe8n
pX8/Bv+34TzpsPCtqp2ZTBXXzIUomnP499xSCRYz7na9UKdUQKmSdsGcx3U9FeRQ
c2kjL/n+LPqRffc/r+9V441EF6mumXiHzdb5meC/W4XyUOES+HHwCmhZbKmI5gxM
P2h8Yn8qtVAOMY/sDFyrMD47QloIoJrh12AoF530muN684rg0LcY47Is4nTNnK58
bXUuRRv1GR0kdx3I3vrarNNoDmOJp66YwSy4qPPKqPqrppZshIpeClNDxFVpXqf8
Z4KdtU/EG6HUoMEbDqc/1ddgBbm2WvNAUV0jcx/pbHEKTI2HyVPSLIDIOKYIUs6l
wD0+KkM1x36zyn7i6LZUm4/aefSoqCjfPYLYqwT9dVF9X1v8JYL6MPghuvySCUcd
NscV2N2NcqlceCIQOdiA8+O6ukhjAPhBE3Pb/JfEJP1Altmm2NAf3fkZDvJqwbaI
iKeuO/D88siYJNwapwLQCKxuCWHMIxyusyW5TGxvxYKt2qsNKssJy2+lIIuxcrYx
inJ5TEIs9zi8XiFtsZKNtiVFDLrRsqjGEpCNup7SgANnq16Ev3jAcuY3Il7+MgiD
wSh36Ep54GxeoxnjRgGts+tUSZ4ubfqMKE+n1r68oZiUgjiFrPE2osCJsZuBFLyw
Be5kY8XloEg1BTkS8IfVEr4yQBnlsQkUcdylDGXDzgYjDXmtahTxkNjL2k/ezsm0
+8CRAFQ6etP8P0D5QPN0qYBY0FVRApXmRy1sg+tXQRxe1Mo7zck4d+wb6P+dtnhO
/ezEK/6+bfC0Wy8qVv7/rh5UkoOZ5YkrAS73VPhcmqoG/9qezLE3ETd3I5kNRdaw
2K1xHrWOZ2Vgkoc6z9FbHySMIo8Mil/DolZR8iOvEAKCvhhdS6aYT6e55flTzi/s
ie2VGMNCuA6nICp3R0Csu64kAAfa4Ymret/eKxlPSW4VkYa9EO2kzohuk9egT0iI
gS4JiFYs5GAwErYLrsX+LAjup343sNmR9k7m0Z5kI41ha40/erPaTQDBj02tVgBC
OfU7V7j+QxCgXzKNjsxsIi9Q05G3KEluR5hfNuHaYkVTlPc/Q3or6zpXbiKdzf1W
pBUAFHuhOJHunenn5UHx2wpyClbVxduLT3/uj4eP7S1cbEzAn7qj1/JssPneBudd
cUzIAJW4S71eX6UgGjbHIHEzIIkyFQzewXvbInlMF1EQm7T6ovXeAmE6UH079iox
/Mp/5qaFkceV/sK9C8VawsKeSaY12WHOoKEnoIJi+wRbpyc5BEwfgtZFZrUGysbl
SIh8vzuBV7lPZb9GC7kOlP7Usw9gRsIugYxKIUDzYrA/i1CBjdR5ihdwK1srd9cO
K5nt7yrJhz9xmzlSdQl71LPdw6/IoAzby+bD+D317vvpktkHjHd3kYtAGvdbGdc2
FxCWp3mmqSNylwDqF+ZDGCtsxa1ZmPXsYHR0VNlxEr5KRDnhYSRoYq/dGGozcAWI
t/Xar4u8T9EgWOZD/0ZbBnGcGRCy8aLsaPpR92lzDkJhh/uegYHFE4tXapdNirXa
0QTuyt+FXbr9ocy3Lzvwq2LBnfoId/cefy3wy9de5ZpiGeIJLn4LpP9OWEbZnaRz
xb+6gifYhCRuzRA7yF6y0QgzvbBJ1KsBEVPwqW0t92u7GVm6wYg6lwYTAYHJlN2A
z/LHulraoCz8u7Clqkx24Box3t6wFdkD9JBYK/EgUi5Vr5iodab4Y+waWVp2fQ8d
tbVJbq/bLBf3YWzHRDAgdDRWGqlQyxDQJB7XDWKwWVoNVBPJuqSvpzXhYufN+lhI
TWbhTP5VGqsvwvJqNj9Xy3mZU+0yu78k8NS28BEApU56bSDEuNdRVg3ncEOUwLjP
H2mdmlIqQCbc0r0TCqsmNuSLYM6/lRNX8QTJX62repFYqm7+UlGAnInTbUN/F0MX
XMNDJjgdfm2mwsXzOLBj91zgngYfc8uem5DxdjpTn7duWkYXAV1bGkmMqdgXpYkZ
QmBE5y9OTAuP4MH8V5tFstsUCewEzW8oCtcWjB10uqJnH3RJVpqEZWylx/7whAhA
K7f/74RoM5oPPzN3uTzXUCUsiurTNYfvM6370HlckqkbvGNe2SsAbkXzD1boxF4B
XLhAa9jABed8h9mmQeuQuqReMidO/uR/h0366ZqSCYtKjSKgBAC+nWayypqOmO8O
HrT18NE73gAGrN8tB8Xu472DtuukxgcUiIZZZSsAHLwSDLEMDy1yl5sG0diuafqx
xMU8/VwqHEntZ/CUObauuw2UzkYpMWHMs9Stl7XFBShJpE5eK6DK/cKLaRH6uNPo
bGMlBEQjxVSx4lEF1qIO0z99YM2N6BX9keGwzKDKwHNTM1NxIiegy7Ih8hOjV6U9
rAuimrPWUVaoaL4wULIacf/oz87P258uGi0iCwQMw9nm+lYvTAntQ25vnTJPS+GE
havbLOxhPqeKWdxjtX3U8Lx22JTwlB0o1dh8hpQfLg+AWhTgA/QVVMhdCKJnKJiG
wzScYQ8ue/4NoquUdBt1Uw7KAsdiKuRiHZLpwPMd5vP53CE4xckkQancevqxrpCR
A8XQVpGzSbakWo6RCZE8jI6eM/CZVdbNWbrLXz/mw7SRcSzHnhLoP7JtO5e0EC0d
IPJcklwy6fKsWhCvKoRuh/7Y9vOsCT1diTFfCPv6HgVScKWleestNMbHUZTexSnk
VSqh8n4/rqiazXV2dcbqCky9SWyxhRfkIC9/1mdjQXdJIW1b9sykDj09xpxlgAvt
QZW+ufTVSjAjcT4HXw50ps/MwuFpi+uHi9yRhIsJmiufm1xCXicPofIB2WcyU+YN
/y5CPgxBygNqNnsUNaRrf8Ca/9DSqebtYgSuzNxyfrm/U/wmpdtKaCgGyjBS0Xuq
XkaiYhatns4ftgvuO+gmYsWDyZNnZU9ZYt9ygno1gZE4WQH9x1pgLolN0UJJ6KO4
w/6xMbt82Zy6xPz9/DVZeEGLscm0HZhwaH7mIDnudMlwNL9aomZEfwTxoppNlr7B
XkqhZo8ganmW14qN4krCZtiYf6lEBti56wrEwVpd8Vl3Z3uL6BpDzoWDZkSspCyR
GZYKsbqp3u7CjKXQusL9rKCc8g0GZ5tmmqYHxNaYxEQlupqxzVL123Zj5EX3eVF4
J6lNYJ61wuT+rDK43zjq817osrSKxMlIUawQUAl+z6HOkcW39DhsuCMbV5Qh/Ix6
n8ZF1aZJXgQPFvp2mkXKiXETDU29vRhRdPcRSmQTIL+AAKA23SAisEUNcxhXBsRY
cuWIuPbjYEaLt3F9o01CTS9y2E8jtrOvIJA27l7J51rAWZbhApygPw7faX0xLPnb
hRs7XCcAGB7fKxQh/rTXEhUzetMY3X6W2Q5cDsFOKo2y30UOrHII9hCTlTSanBlj
2lXR0bD3bz+NcaWFdu5jhbyz4Kea5Ry4ED5XfYIap/h3nU4jJKclZYPlThSo+drA
IekY8XmO1oK7f6VySrwvCmeM7blODUinGU+R+kLGZnhmf/NjCe5bwuLmz2By3Rza
WBk+CdgOyH+tf5YfGhVFiZyP2jg7K5mtPVJS3fAFfhDNStBqYr+D0/N8njFYuqmm
9JmGLhkxM80me42aG22CV75Jxk/vFwqCDYvC5EfsqaWu8/URilcOynUYJuXuCO2c
MJrIBbk0/vvyqi6no3ztkvHVwKAKAS/No2xwjYCiYpuEGvF+Cq7+oAcCcSDrc+WO
Jxrik2VKtoorAM85bL3OjtjE9wH1Qb1ppb5W2s0Ddyy2vaOywM25nTQGrXxgQ7yg
vKtVM1I5BQjsqgife2/HnuGFEAzBqOzguPobcr/pgKd6dPkqb738bsK5euI/oOqX
UT1uWmmwLK2JFHuJUfJQD34ZQ6Y4FhUWS6STs5XDlcWEhMlGQP082YemIPoXb16Z
1u7t9lP2a3RyXlBIApnJ5yrbsb7uBeW44djghZ14wrYFFBv56qm56zYAWY6l1+7A
HrqZZRN8Xa53/a/ZEW3EVzsTaBzJ4AIopSwXQgpFRMnYAT/zpXyaclio6D8CbpZO
o1Szj+fnI70FzIwwsmZ1j4bmvSVzR0wmQWyZ/7NY2cKsRoi//m4e5mtoGlQTnPk7
qQgIllCs8xZOLFT9gyIj+F2pAGPC9NQPPltOHeN00k0yG5FzAOpoj5Xi9BxVb1j3
igNh4M/aUE2Y+Gl6TuCgD717bnOSiSbyS12GzeunYvyLBN3EK7BmkdOsliv0cN4e
R5jWHzEPhx8tUarXVse+Gai9R/9V6jHvbrfUSR3mCewo0j8q1DC1VYguFopEwpNm
UCtfnF+wxjuowlVr2o3MT+/awpnfQ1ZV1nc43cqe64XmazTA8tKmDCh83HVQJ/ju
isRDw7WqMgEytvK+zOtoV7TqUZVWOZTWYE9SdWfhsq+Z5QLS5NTaan16ODTaK6aB
zKI/KypG/hmkAakuEH58R7ukkI6tLRFQMAUu2uaCpzN2thYyS2uoOOLlp6NnKJZF
M2drhpxX23JKl4BBeUSgMFjWOvUwN1xY8BX9Nh9SGR4RKc/TJH8usDn3od7mI5Lz
5jP4+Jouu8U0xNzg5Om+TLo1KieuX+jgvlMhpM8Cqe2H2dhooiIzH6iU6/Il1e4d
F095RXGD96hmIirvaGLrmAYtmwphWMLoErCFJ9VeXISGC0i4nviO8ZScZ+fmUVMU
5+v/e5aBspulFhsNirtRJs2WRriogPuaRdWacEx1wwoxdHstZdqijctbRAEw3v0+
VPbk3vSnmbTc/7Zhh5BpA7iLKsflxj0Nf3E60aQg+uNMW2h7t/7xcaExNgbnV+lD
eztzhW3GJn2n+6mlCFW6iKttW5zOoJFKuO74glX9Fe7Uh/bQDhECvq29fdviv9v1
cdOWEVAVkvXw2qvlnqtEs1euRufxKICmc0aA0C25uUAA+gpQFTQNhUMTvpiQOl6P
OZurg6DEfxDOiiZCwoq6VBguIu+lb4tcnWW7+lOxx9XTKHnlIuo2i+2pRZkpvvzf
XWcruov5xPDGq09aunjgv3s15XF5GeO6r/cSOMy543P4FTYms/PuR0OdaF8feWkL
Zy4rGG094R0ocikPLY8L8OAZaI1t4d9iDR3KR1ZOT9EXj//6ZAe+IRa8OTaxNzy0
8U0zkB2pKnDsApK6hg6DdbxdlhWWQuFfPosM6bwF8pd2XQ2KSZTg2U0zh1p8/wpC
1600wyRcExHYgr64fMJ0zxwOkOU8iei1wONuenUkOUqEz1Sj0P3A2AVk1WYvoPIs
tcENm6xXsk9VmnncJcQpISdKHCC5m/Ey6a2Ypi2PsilzwAXvKW8SoFRyWtDZD+Nb
IcIxqkFQQCpX1N8lhD6UkRYSwUco5LkqFL+gA0txOVq1Y56bA7jqyDxGiV254B4U
1YRzNUHn5D6Rph73NhhnOXngrK147muf6/J8HHaqyGtbNRUOOfSnUdPaG4vkrN0I
MZev9CPPKAFBFL3Rrf85FlxPRNY/q+vNJ5arLQ277q68dW2xrtqan1v/8bxwBOOr
m8ELocwYEY1zNWRaGYFer4+SvnAYdcEXE7mRxnneUBxR4Cxv5iw0oOovNppMiIhL
nKJRljSqEMAbtHqqPxUxm5xMumHzOnRyUUvihmT6AJZK1xeuIKiNnwqmhg9MBicL
MWaJ7IZXiJlgtFd6SituVxx18pkUw/P1pC/YqpPtQp69Xxy92TmfJZxqCCw9fyhP
/tmLABLDakOPoH1CRRlbl4hIa3lTWX0yZ1B2SEbnrLcAjQBafS1BSGDe4wLNNrpb
OPZo54b5OxiMpX55K6W280Pb2Uhf2mmSsiMWD6PFVDBTRP3Cftf6thDCHraoq5zQ
rz8lDaERe8aIP6QcgVQeHIivcQjM2oC6ajS1dslsQCfPWzgn/D0IkHUoJmxmsIFd
uUOV8l6R+bAf1YsEkE7oAwUzxJYwoW6pjFzFQO5bAlquFyniGYNolWGV6coYlYXH
cbI6BqK0iHc2gHT6ks98wD4MDr8DSwvPL3qTO3dIDHr+IJ3WDTqgGLD99IO8tkFP
cywhRCHVZ35hXYY/cqek1gfT0DSld50Negj6u4PNB91tX3wYNeD9fmRQ6H/GfAsY
ZpVnDj/mwa0jDkIvzp9KQV5FS0OjG/ujxbQdjP3o0JEPKT5joAEOYHUjZVKiM50y
hF4Gzjnl/Lz4QGy4w270/o5947p2ugMkl/XZo9/DPpvQeVe8u3D01I3rS1TtW7Zl
w3Fsmz/Qp49wNQARzwIFrY4aTUwZ2IqpoNQ9nHQ239zleNke7bQOZjfz8gGrdXiz
j33f5YMFkF4bS4PgAb7cvsOIrqAL8d3Vxo81pgi96TY+//jgcWOvFbFbHkzJyRWh
DsCT9VSbxR+Ln6aBDH4qf4cj+JFRFvL3z8g3rgtMmBVCfTsEy2IFTEMKn3DNG1TL
sWDzXlmMYSx55PodntBOlP+dYma27EQTco4TYM27VuKCMdSjmpHHOhg2zhEaHav4
n55b+g3+dqEu2WYmWoSz4WNGdvF93Xq/VK5xoQtyTbH7nSoRlZvA7KXV8Xss5lmA
P/VySF8M1cZ3xZuTAE1xBEyCrABolriKH1mqGMtfX4c7o33qCnmwYeERdxr4xazQ
C2mO4e5ehANVMbvjOmz5IR9tnx5H9OxImPKjR7kjLd+p63IWOPCNq8qCus1JELa9
e6GvHaROapI3JmiIukGLNKrZ0NWPEraH5swYEMSbvuAOhPxLbQgpOl0PqFARRoBI
WMh9bdIcoJrpN6p/8b8UllWaOmVfKBeAMRaWt1pVUb0BpR8HVtNqQbJbqPE5Vt7W
bDP9kOezd0eIVZ3/MnHo35GLpDrdN+XAp1xAIHPH8akp51nNAM59a8rlMpCmigo9
IR/CcpzQIt9SN7jS3LhkCUk4MLSaz4wSj+WI24uVCKP1ZgUHLqboGShTSObZ9aSl
73XUJtGQdKKUUooWLPlA78OLlYyc419zVZrhZ1K2ZbuCaQ0wtcrO7fOie84R9UpQ
UtPkvfa4O2s0dpC9DTye9eTgrP8Y24yKBtfZdFL3bRS4gMeDu1zXKQJIPwcxHfZl
BwNdbiD4e7KmnGkJZ/7eAcWcSSWlL3IoNKQnvZLeSmRpIM2VsrMaMhRtTrc/s9ci
hv4239inGqZjvYJsf7cpY7X+jU4vXDR7E2Uq7rYW8ylkyCvvZf0M1emLwimjgOKk
Wbr+yrYXLeiSophdcF/qz2jXjQHfc85k47y4ky1HouqeqWFUVW77MntAUtZBcQim
YMwXKLUw18rfAVtyRKZYPkRtYFnqBTXRp0wgDcG+UAq5uPThZaPCUzRAgZgLOXTH
ATerfTtHL9Bg+av4XH10ignRNFchCLALEUNdkWyF/qxmJdl3l1pIrO7WpQAvY8nV
eo8WNYjz67zAGHlNGY95AOdp5dWwRxp92Dgni/KgN5+u6WI4AqPWdaCJL2P8A6qx
yBeEOyrtVIhrWPQ7PpKqsUDF71DgLlMByZ+CEbwUBijlmLBrzDWtBZq6sWofSX+V
2+1ocJYO97+FG/XfiY+tWH8Ctpa+m8T40VgbyFf7ZVm5h2uiF0VE7QZNt8huX3y8
0Q2GYbsqH6gMgb18LKj0PIjsliJ0CqbXbrf4RdX9NlBXGa2XFukbsWsBZs9VBrO7
suKm/iDLPhmWZhLlRplfzthIY/fKZRLP06zzRI10eDebbewGJFa6vLwkCegNCOJp
71pRMCzh7xQ/e7fXZ7FAvT7MqSQa5uR/RRaXgBiFKX7JTuAwVgLAMg4bnPUB9keH
uKTcl+1iwF/EqCgIw2ynlXeodxntuLd1g0BxXWX+J8GlWTW62VC1z22FeWM+sw0X
X1EDlF9FVTEU5D6CoRNjgAv8/aXb2MUrEj8MNGgu1KqeiNFB/4+1rqlrg2Cmsdzb
oiSrXB4sP+MnI4UUrnVOGde4pVJ7FLovTL+he0AKW8jUqO3cypyZuKMhqY49+IEO
ElbEMTiBybh9ASbPElsIdpvVM0KOz1gR/UZ+Pg5VlFUbp4k9Q7pLmkmrggyb9cZj
4iVhnRiexTdQ6lmsMs/des5/dU9x5w7xSjBUX+wcwGtJpYeVxrp7FA63c72IGCOV
PnZ66Mqd9EbjdwLEFAySfHfhwE3gGWEGujuGVSMfWTI5Q8M0HxS909sRND01K8c/
J230W5UPA1EVfbYKyf5hr5CwFztwaPLdksrWujdFDzsB2yA8+aReImGLyBxOeqYl
axXwBpbl/udauroxzDHu2JyxdjlyxUsyD4f8Qwo1QuqH5b2tJI8bhTkcvBeu/iSR
O69uWwl3Ap92nvdIFzim1/N1Ww2OyPBgsmtudx30trDmTn8KHCMCGI5xLSVV38AB
VrfiVL5QfyLBR8a0UWjydIeftvLm8biLGv9oRS9lJdZZB1yRgtkaPFUIrIi7OocE
ly9IxunMzFiZneN5TJ8L9aSL9BNGpxlPdptlb5ESp+NihytH31LqA0/o3v+C1+ad
kc1HQMx+qQw9os2tx5AJ6Tm1Pyie1SOyOLfz4r/SkoNVFsUg63+uuexS53Kzzaun
Qx8E3FdjsH7/1nnpbHbehEobz5i4xL67o9UlL/ZgjOSu1D+t+s6QKvx6G33KRNJp
dBGeYaePc/j7iU/lsLNaq+KrLa+RAsV7FVYqbTEGMA697tm2xwQShKhdDXvUi3Uh
oddM+x7s34A8VdUFs+G00ndo2VORP+cem/zTSPtO/C3rAkiurvcF6sDZxb29YaDN
2+UoiWlpf7N+v8JTzbUviCrhnMWMhP1SPCJSN6SJtgHgjvCy8f89OdlXG75ohkvp
1tsMQBCJQGAnmHX9VWipC5vek4iJ3q5YmuyHqrgQfpF0oFxWMC/mGaZJrgKaI98D
kISLjDc6FuGR62ncKKIdE04gahtDVYNiJO2lnxmDj4Kyi6QFTxvCU/PUr24nAcT9
208/I4RRadMhQzce7DdpkyjWSJr8c+kuBvvbVWL04nPzLFKuTXJLZQV8j+FQyGbc
Jbrhb7K0j+mhinuFEv8tR2tKku9LEVx7y+qsQJyxsdqO3pDl4+8ObqXR4B5Dpj1X
RGfQ/3AFYTCWL1C0+c3V+39r5mT3VXwpwMoCN6RBM4mP90lupvIdx2uoYSa5xcjP
/zlG+BX6g9KDsnHTshpsDTnFFmj+8umzdKVUBfQgSXYy89QjS5HPBL/mUx1q9mVy
1dkiCAs8l4iOSQEheO2owwSgM+bY5jt3i5rc2pUGWj225FxaE6kuUaUlBVSrUK6V
Wwp16+q9o2meJFNjziWDlcnE4FCyp47vp1cOKyE9ImhAGUfYzh22PgEVPeH+5OQx
HM4S2zzEuw/FHg/7NA/uZwJAXZ9YEw9w99zj8Dnub8QhRK8URwl0vy/9XD+44iJl
Cb7QT5p9ehF2yfvHowioFcHoHp3DI8V3qxhFX3fNQYrQUPxZGxLzArqDX4Iv7QJZ
Olp3b+iIJ2qq60VwCK5934PYiqf/z8J+jxca65g4SpzkK6itTJGCfdFLRXltAIYY
bSC5dsOzx/m/UG9BZ/h6tcLBMhlKrrzp0vEz0UAte5UDTCywg6cSw4GG++qPW5xN
57ZQIo4qv59rcfqpGVY3ucKBOcw9zb6f3Y7pHIC8I9hKqzPvCxNNaWbduplUte96
Xw99FOP4oCPRi0NMPW+Y0yfUuhx/HFhnrXos9KjmwofPmkb9mmVu8YdZYoWa4O6K
UpTUWY+czB/H4dZdZrRry7kbdpPpDFO0Q1OeIFxBcGI01KKsyKZDvyxCGMnd4/wu
VOtLITTnjM4m/GPmH9QUskVZm1W9jo1qI5nFjYCRJpQHKgL+cGeiSd4tOMgjDyO4
jVscLJQLkLarsssPJAh1w8av0qfRBIVBiM0RIuTa3vhWW3mJwm23m+R5YP3i5iRo
6kWOLFD4SHkYzDkxru0lp5zDkziepe0lkP1geavcNxe3R3bJryPSiV4WETWsolEu
grJQLq+97Wm3hFYjRqAWGBinS2NwoTRQIccCU0xQaABXEfL5W9bIIMsqQFYHI6FM
3dq4GmnWgAlnE9vyvjeLcMPGpBFa0fMFGhOnrh5KJ3SGoitdIpoxLgb00FJ1HVyY
DwPWanN/Ok2tO9B2wepUoRacRn2lE/YkH+hb9GaXKApLYgshCr8OsyXWuN+Wk3Bc
ttaAnNsqGJeTDIhHqlU6tmtYNfp/vk1aBUcyNQIueNHxlNbgrE0ZENKlq/925OHn
QOzAICVSArsdi8X+iVllelqN3eEEdjPyQtQmntblrq4L2/TE8e4LQKPXxlmF/dC4
oXldXWB6G14CPOOyXFdi8/rcZPpVDV4TL/JKi9ksYYqrK5W2tJBV1ViXWqLzfl6b
vg9AcT3fBkk+ushHfu22mgPGTNCXMun1MQPv27aCgwRvxhL4jPa5ofcEyHudYEaB
NOChkcQFS8x19D5t0jFUXs6Hp0BotsbMfTG05Kz4TBWhJBtlC4B3EyFQX1W2ue5w
TO3FR/L7hfv+8XEoscLNigS2ghaZsrqb3zGf+iEGDukUBlrfFEkss0ltY23RHqR5
nQGdnYRl+bn5d7tseFXdrhO2WD07hQ27KX4Gy3TqDkVvU34hXFk5Fl9lv6lbO60c
6b4VRPOSVxUrpWWajiPFwc8pXBdrkL9GSA+SjTiiCSTQaIllRZt4x3A4sdDTtFOq
0XSTKiqXtwBXmjxMTkgDl7+66YXLcOst0kcTtwZQwASe+93mnW+uTq3wKlYYfami
rjft7WbPKrTZkMez2Bh08uPZpcXS/p0PldXJ3EP+6253lRYDgpFJH0AvQtmFlBwH
TMICW4RcRVVBGBEiQktCws4SPH+7O3FGSXu1IHYLROohq5OYVT8AoMzEJhkzU8By
LjVWofxvMR4FVPdhqxTbugGD4Y4UsjF9GD4mYDGY9cIBwCsBbN3a78wvfSip9x9g
5NL8o5GYgAJnKmHovmYOqwtPai8nULJJkSeRxGScEEO6O4an23RnoF8osY+OEDlS
s7Mhl8OHAWFJuYbjpmEpXC4JgsiEWw2YmZF4UvH3gIA6VP1DniNQz4u35Z678HQi
o2tR+a+Znmr9YO4lONvcgbwl4Wxui8RDMPDgf30UfhODcjeRWDjEoVN/SqKfMyv9
/W7StgrWUwfwOFplD34npRqRkVodRSUDtI4mfEbVGKSB4soJz49A5uygURhjYNco
RMg4fab7vLbd2waC/1nI1KaT5a1bgn6GAtwy/oKUMa0ovdwJ/2Pt7wIN4TSbd7H3
bPiJQVNkzeD960RfPMRAjBt2hHXrWMtW1Y0NMAvUiY6LyRB7ZDF7lVxWuSIuTH/2
u2r5ogtX7bOrsN/U2XsORu4doFT0JsPYkBzk3N8/11CshgTcLh+YUPgekyavTmJ0
MFLt7BRKOImlo6e5SgCc9NIIC2X0L3TaWcth/2O9p+ra1kDs0hQ/0kc5U1AQFxa2
hGGqKHBGjJqCgdJofQVGw2OvtIYu0kw0KIGcwQORqcaMVs57u3UrfEbWa4L/MzFa
jHSw9VmkSlQC2rbldppGVh3Fdyo49wdILmNN99JXq0ud5PbUg3hDqV1AdWW5W20p
3JmgMFaww8TEvleipDNkbfMXRt6AvM0XbmescZHb6dQZkz1vAhaOKmJia17PlV13
jChRDb0fDQeTPG9eaIBGn0vzEtMuVeCnQPw6kgVN0OLczyjBVlzbkQGiwKLuB74c
APBPMMIn3YJjOIi4tK7Nka4ju0vbRI6v14wwhN9hNNigqECmBuZBiw74wqINVVka
0ASqyNsmEHXWR4rKO2H3F00hHSx/22QbwTNAQOO7YnWCwDTJf96Ali5yGH4Qq5LA
jRahSNgEuGSFieY1sDjA6pwkKnZlpBleuMzHfWnJaRC46hoRj3esh4huR+/+IW1n
CRxOikGOM7W/RVW3tyEEfymiv0xnNa3FPsoed/o8ljEc/nlZqYDEqUKur4JtUckf
anm/OThpApFHxWinOiHaUcpug9Qvms79KPX8hz6O5RthrVTjQhp8Amz/+qCUafrv
fn+268b8gfEIh8yKBGT4Ey5lplfOM9Z2sxHlHazD+abu9b5wa72MSJmDGh9o+rtB
6z7+ZG+NdMuzsVqJoLceMJMRgQoGwv6q3B9czj2wfohy6CJccDUC+IHduWiXQe5S
4ewWzZMB0zmxx6oxPeLMbSoVoFpH8Da5EFd3vQB3TncQTyh30DsFvESwsASFCG+J
wJSKBLvH9QgecTK7wPWo44j5BjIQww9CusELq7IySYW4Vl35oVRxf4GM76+IIOBe
xpEUoigCy/kg/BHFrto6pgg2U9OiLI8gkxeXxyGiclkmlT+U7ecc+Ddzn69uIjpE
m1m1tUHWPyuxdbgcbeHrxLpUBfJU+mI3YGg/KDDHN5xk9/TqfljW9zh6yO0Rsy2U
IE9MmIX5J/FLomudZPgbS1uuzjZ9JbMn6Ta/FIUYYQ4xCy883vTJVVpXmPwnWohY
QPUSALTdVm4nDoumNC8o40eD7TzgQdZ1RXlu1Q/W4HTPXnnxxZuCADwdxw+mcCju
+0rGoXTlkq8UJisIqQ3Y1QKc1n6oAscExbUWYSbiiD15mD8H58iAfiX9Uk2U6Fl7
WxxugMElwXdqvb0emdJsy4k45Je6NSKMo9Zk8AVSH/649wDBAatMZpKiw4pTWoor
QUEuCvE5OsC57k5XUm5uV0ueon5nNryyT1zsXPjDrQvhXSjwTANjY14VFFmcYMQk
0dFKE9sO1/TGrUKRHe6CIYYQXKcBgYDPEQ7wMsQwGoLH5PPKTe7AwOZ5VZQut40/
ZcLtvnbEBE2/SIe7ZBVBTuAu+xUHkDcJThsn8TXv3SZ3ur3kH3L+ttzAijLyt6Nu
bbHSbbnRwPn5G2pB0hMfCTK6LZTkfaidqXBHCosel9TbnIQa6zN/FNqTInypSu5l
WI84IMyh++RM6ia763SFah7xBwdbm9DgXAs6lQHKOvx/lVtTabGN04RJTtZzla/B
L0Xdasucz8viaLtSiNwPQ+YkOpCCb76eu+jCrHFC2RQJYBfG8Hzq/f2Fx2JhrSWM
BoyNPayBpyyVaVvkW8SRM/XI+J9wItYSI5OmxHVz4gcXXhiSIB4daJEV9Sve/vQr
/eF7MYT8hlEdsUh2dxn4eKGT5MYQL8rMn2HVYHRzheUNDCunPLTOkAMNWIHWxDwb
pLY53UHvTtO6No0kAoaoLbJphAIMvoSwXl3nq9HQKKenTLE09uwkplet9aAqvdoa
SiVKqOpstNycYnOyVb4/f1385yIBlKJ89cUWdt90rPeFi/yzJZGM9T2LD3KVK988
xeMuCrStbQ9g4+t1UGPeuwJf8ZmW6CKLu84ibMnW338ZH/bVp2U7eNt2KEi0IE0Z
LH8sNRV6HJncfHpT9LlSvxtHg15j7HZDf9vmf2Z4KKfdkG3N+Q9Ov2elt4qSD8y1
mwmZH8l8HoWG4ZxBVwmPRq6wG5I6yzDTBEyFdyu4xEdg8VAYkCS3g0U510eypRDs
bJmHvP0unn/dUqRSEUxzUABEB207uWMEzzuZMDgENP6r+dg13Ofxw91CwLnLONG1
C/9M1BpO5By+XsH+iAkVBxFqziw5tQmtxkU6CGRiOcra7ZNGaxNAeM3HrM+6PavY
/7EPfv0Z+EoGWJ816kv+Jxetq1Hfs5hZ0efbnFJMnqKp6wEPg+sjpJEOiycXhXZV
X1HegwurBVAdDHd1XIScYQd0zLH8jRJkqvMRStU8uLvIeK+gY1sUu85JpzR3BIzE
HhQ0Gla2/dhp/JdL3XuwKHCDTVyHdeZqFAZCL9yAGOLLGF+wz0eNAStK3TcxPGWd
OMywEvlUMbPcJBQyLbibQJtZhCrVTVvql/ET/eljEr3q8P+PdqRYwCoqQaTkgY5j
6jX8AVlo7hQe1GTm2U48vm4NkkD/H5VBYEboRVIE4LnZECxbBSFCTAWD9dDxWkxD
KLNngiUeckg44+P7hGaCyPz5Yk0l/HvV+vh1b8kjsGblJJRmDBPWl6rNCO9DlYA7
dHWVkyN7fesL++xZ2Qshqxomh5qOXCIQgNG3yegwt2F2WmDGDxcUgA7Omyl7Fo4w
y1E6j0itDDAmlJCYEb8yy5da6N0aMoGplnhoySGL91wu+Ia2gfczaCtJxD4glq3o
/iUIhC+sA+c1uaHPgxW9KQT81QYacART4glpwxmEj9yC4bDXc13u8fPB3YqJpcfA
ZBQ1P8OiZiLSVwZ+rHLW+U8susMpqjWkchj3h7ukzDeaFyEEmVQlM4zQrmTck/rO
14uQCF4315wiOzZB2aDYq1x/+dVJ079Vu/ZKpySPUis+Cla+9ZwWxYvYtuMCSjIR
9edeN+TVbIi2mAfr9Sfxux1IJxZHM9x91DMUXkoX1ppMbpIMYhsaoWh/a+ApuiP3
K94Ud0bPp6+/StH7ICNOGuBcrW42K30yY8DpK2WT+Nsd3igbJD1RMsvBiMc0pHU/
K5HXq+EZ87c6oIxWB0BSzLFQNGczwY5hVI+BdBqXILSxWnAoObP4UHueIyVpXs9W
bK7FuhR9S4dn7nUHSD7B6Zh1NQUijBeir8ywMTkJPon7A/KyKwWx767wDIS6bh9M
b9B60FSGcK/0iPZ+z70x120eoYu2NVWqV19veRYYRh60X8kU6QzE0hScmsaCNoSf
1Z79xUCmTVFpZNfSr1cgnwudwvXkNGxNvBOG0PPs7c1L5mVmAqcrkcM7fQB4a/2f
PalK9P1B2LAS9SQogtxtaOzz5fRHwEEl887QMUhCQi3g8dpStnnDjUywtfx1GcmD
WqR9AJugLTUoyT0mfBAgBGx1UIa6LlEsaSO0MXlUzP/vKfc0OunNC+CVzC++HMh+
0wB9YOfY4GTeLNnPTjFkB4FPXVjwRY8DPkOU5oxpGWqydfX18VO2MSMf0qaJtEl3
iCfKct1C+urw7eqDEgRFigzEcm9ulmcSdGIYR/pvdDVTiJDaMx7PNmKxRM5wrCaO
xqXvgYnJXYO4nHmS+ZZw04sXRtyw7s8fV0XFtcDBxWm895tKgdQR25MvxiOrprJq
qwnlVRfasIsGuNZHBIhztBI1PbtOxNSq7iZBdunTvUY1gIDeHbUjVNNrzCAlLqCn
RJPWNGAuqpPdEDaG2PlsRFZSKdsvfSiHSgT3fSsvVOGZdTVxvLZAFsX7rvjoIlKB
Lcl3rT7pz1e66Trxn+EnWBJY8wj9eHWX1hEJ5UkpLM/tjrx/P3T49TlgHCWeHIcm
+tgmFl9uwDhrDDiv8k8skoZ15/xpUvjEiMLg7I48mkmMfzRUdOJkDvIcta92xXia
6qiJVd7Uz6X5ykrLhnNPtGwatoqL69OLzElkJ+IrUFVgQlBcCamWN43Tisu9RnJe
qJ+OBFlmypz4dE7JvwNjc7zLNwoUkgbUxTAiDSG0eWP+dDH2cMd62ECjW5jl3gCw
8waSgu8j54Rp9ctY1tf1hRk1QjAxUcL4JT1ZrNg5k/sUanYco93RAvBy3HUdsZKz
81hdoBArMFSZgBLhB9dJ9+ln9VIWY1rYsV9d5JalkXrP3x9TJfPJ1RtCNjKUPw2k
cKBF8iM08HZD4uyxT+knttgAyp1Adj4ZnyBEpRw74v7/3w27HfMBkwwl+ovl1h1v
Fn81hgCcVucaDlBO6o+CYGqJf9mjBcY/FuH4Zb5t5JLGPxTyv3kFDkKI+EFKS0oR
Is467cV+IfsI9vporaTZCwGSc2SBjsQ3aCpQu/YRuTsbK9aQ/Pi1LZ5CPv2Nsop/
xlyuy5ohp3Hc5HRbLWskAm7a3YXkUQG9ZeOiMwsIhEabKfH7qdt1ChTfUQn9Kjsy
uK1XCciJI3kterbJneEx0nakW26ejzCxOqceMOfiTLiOfn6lWEbb9fNpQc50Dlj/
X3djPNZkvJRgj+JCRYM5apO0Rj7L76Ct5CMnsDhbrAwC7etkEj/GOSi3buIrhcAF
O9liRtNt/h3+CY05KvZCZn7PtYu30vP/s542gYdG32QSGHcWd2pqK9IGYS6MfTTd
NxK/OreVk+d2OPjX4TPL8xhVG9AIlgzvbdQoAx5ylc5ZSMGDLhq5gKTXto3bmspC
PNU5mY99FnGnIA9XZ82RpjQWrVZPe304gv6AeW//9cppfH7TeYhYG9LCrgaYS0W+
sDFfY5z843hh5jXZz0t0SVsxwJppAGLf+3GUZoD6+ZWk6V/3ZKA+XLbhODm3t0pO
bkH9tKBRytigPu8AWfWwYXCGa+H3DkXTZVfryM4yUpyoZmCjldhxYJyU1ux1Ftc0
yWSK+bLkotoHp4dyJXtZ7rDI1pWvggI+wTECsYN8hivYDGnotHXX9Pz7ogLZXJKL
mW3pz4yb41Z0Ymzfqjf1RlRjlanRurtnvDxzYcR391ShobOW3OueL3UibIn+AhHU
cHpKXUEWThPjZdrgeudQsuPc7f+o5W/fpQG9UkT/dqbzqFm/mUorYCwfjGX4P2PZ
gyBs74BcDOG8fghn9P4OPvgSDLLaV/zVEFypqE0MVEmMG5o7YKxVOCK29fEDuVh2
a2qY+Nre/UHSTvUUHft/TfWW8JwUgtCUjhxhVGhRIS/x/BCZIwlRBEoAOwdmQyNe
2cQRCw97ynpQHKmCEqlz2Pgn5NRMZlnkcZ5f7EYQpJLVhGHS/rbc/mqkB9y4SpqS
aVDKyz9Jno1EF+7zWtFVFInzU3R5oaCe2c8aHiYaGPGZX/hSoUd6yBTYHZBCJ47V
4vOKBUcv6AWBllTx0Gt29JYtYX0rpg6jTM7UcOfSDGMEOAw/fFxQM2UO/e+BAk1r
RAAkjLh7biIuA7hrgm5o/GwR/OrJd/USBS0PBYfZ5neq02TdG9legybrgonebjth
+ysZ4w2mG2e3abZN3JhYqba2Nz70mgXhebksQU9nLzrqqZAqoFT9MIs6ArD5MDJP
NSHt3mzM6YXW8MScT/kYaDAa8mDyGAxcecgHIzdxCW4SXThFzVIoduXPq3waWs7s
vOooBPngJ9wl2CTZfBhJpJdSGi9nHxJfjfforFKWqr+E6gpJViZ/iDO6tMU0Q/Vb
0moWRaNw8CrLZpfUVwMmJlByM1beadQ88qjlcGIxnxKRmpQlGfVvCwHNMGQ0rKS7
mS93fbq0SI7LMHsX0IdMYUwuMzbng6KwTDpEcT+zN46d8OnVd76D2teTmF21LvaA
fZX6745SV18ywxkJe1FZRlTVpbkjmxaDb60m1M8xAKsdohkuZpG4+t1VqlXJdEBx
F3EK1pznePY+1tKtd1BrisdL6TuKLxwVXnCwgKfkN/2uhbDQNBivhDKnvZ41jzCM
NFRihVhOdwsLYgXK9wxSVT0tw3pqZjfg0y6ME7FGmN/HqTMwM/v9kaa6PhOXj/Ek
dXZlO1I3bjG9Fj3I+t5SMs7/LeQ/ZX9Q1qdoANTYlaYftu+oPPZRdYog6wrYM2TZ
5qLg4XxSmg2MqI7sIPvR+bW5yoIFTiJgk6AV0cJPPoxmukVtwwFeFSaqz+VovR82
eknQ0hCT3sF6aNy/dAkuqQgPd/y3+EbfMTxtPmupzZS72qSZQz5uXCt4ydRs/BLO
TvPyBHV2/AAzzbDFnKSHqsLai98EjQFTBB5Zz6N8/a9NEAZAn25cQEcWhINPZ6Tc
Fo/rJLcs2JfLYkuCu/4beuoQJ9V4h1eFwOMIBe4EE6qiKn81pqXIkpHqm5GrVdoE
XRuyeh4xify5uuskE/ZyTloBk+JLOMbjpSYDLu7+cb6L1pEeMGAJCDp8vtbJP1dp
WCZnyQ9mR4862tsKt9HHAF/OLBe4WTXjOHk9+GU4hxWG2kCqQb2nhlFcd2gpZAmd
fywIuAF0tI+wpslBft1Z5L2LnYLKHQsxdSIZmRK29L4vEqpUulgpRO193ROK/EtV
263Ym98LLQJmaLadaSmBPrHjbqGXPLuUFDU5PIH57GRqqxZQA+N+iJ6z0EfofAyJ
wSnZ8dQWavYY082SYALiqcv2Wuraea2KRcLtkiBSlLtwzNAptNQSgbhjeJsub+fw
kliXlEOoV0dbhTW4Pu27KlAU/xALVRq3A5LNQCquX7mZrA8eBzD0mFzSBstj7+jw
8dYlmcHfT3OOvJOWl5ua9fQ68kLaMJRBE+cCCw8RiV3VZMtFxZAPNnZK4cvoaq2R
7+lHBF3ZKChYFrbdJSOEZ5IgJqW5+MQfXUajdmWVhtICvPin/gO3F2d56K8N/O3B
65sRTBtVDfDI+1KfHjY2poL5Os8lg5FP4gkOwC9OShTVSZfmk4+JE4LkG51gcCMI
JENLUjF0YZtNvIrN84rESxjqBqIPGqzy6FqG2vWlJ8kWkV4e65rNwjQfTsm3LgVh
iDGerzVQZEimSqsMPLyDeo7RKAQJcqtlVlLPVxfavuau4phhABvKJtD2B/HBbpJf
SSMB6L4Qh+V9gqiYeUwjvACAD1NPWuoN0Os0vE5UmlQHCe3QoWijjY6r0YkRkecW
rMoDzEhpREIRZ24KuvR5AANKkbrxdvcE/x5KxGYAfeaeQnOH7HdpA9T8hDLOTp9X
aTxoMrItkQS/FH4lPaOPdoGLDWYZar//DaEl/hI0TuqP5Ncm6O0C8TeNls4TKAIC
ApA1HU/gId/ECATZGJDQBSWlCtHCsmudHVrWGp7O3CEN+BWNPcp0xQl94jDEF15x
uuElOuhJoslCWjcu9g9IpmVJ18226KvJ+Csqi8gh2LxXHbuCtwmADuyAu58Wwe9O
pPZ7T9bo8O3qCcOFQYWFxx7gfvwkT7XqSZjEj3pyPIAZH99jtdgSweQ8FSZDAGOD
7cGs6gS1ClrAQiuBEednJH7gw511y/1dyKya24eudeza6vRuu3+ov+xNVgndoAX4
ha7fDnrGtbBSYvwdezJybqjuLcP2dqqwPMoKXLevP/gXmo+dvR3IhF9ybgE7/PGb
eUo/tEjPO3QNybANhMUZA09LbnF5GPQcsgpHg5fzseG5oQHUPR4ObxIzl+SUj7TF
EVUEh2u3Y4951JoEklMN7ZoyM7jtLwQalnoEN/eFyixB4JT7bIN+ZNR3Mms/nwJJ
BswoY7H7T3F874Wqe/F0Kin4gYrfqk/rHW3c080qx+55aWJ3ulcCXKLu2R2AXWHV
Rmoro9pb65sY+MwQd1kKCvaxNRDhqdTBzOPDD0XzB6qsqcvSG8B1Feyy+oJXNGnb
+yANsiUVC2SMQ3PVWBQ2hs3mH1WZse5WNhh9uKECdfMmmI5qKRH5phxdHp33rVYX
U+vsViNgBsynBdhSx+B3HTMDHJCt3jumP/RyFZyXIedj4a3DMr/lgH5egerF8nJl
fien2gX3qdOnTdM7ug8aLL/wZHNesspNE5kfp8o20hJGffRo5Vi6FHNb5ZbBXTd0
u2HfZIT+z827tMRWO4H2ZeaXEGJZH3ZtLf8+FD6voW/2LnaQzglVpVlcSzDBnAho
Ujy1hEKvHyigRTqPubgKXmqpqjVPdaPqymd1nwEAfkS4j91kBaTpliyQ/QvCVPzC
psAqpUzf9HMUeVvxtAJpPa+Bossw2KK7V0rd8PMtbT4VWutH9UHhlBIJXj+YKUcW
5EU7aF4vrpBTK6vS9pa1LToky2MznOQELAtE2eCzuCFilXSreaRt5If23cREaPKJ
nF+nqrtffMvOnKTyFXs2nLF0nhOGCFSCau9eFYt3Myo1pcHGiVlwwnZo70efb1Dw
QSg9XVNb5uUo08zahGvccaMdH/+0QCqfAzvJJqPlCJKjV7uEK2Ulf4Q7OB+dr72c
8OvSrSFbBmLUhzZcNi/YG7lwdFIHeS4cMtZUCqigkfoAMoqpMGrsvgv0vpieZC9i
Tl2yXH28u1xw2ut2AVXmk1qe1xCD71GvMj0wIqxbKhjS3yanfVtfjm9mo5XbTEh/
eAHQhQMNvWG1zcsjSrvPmKIU3kVHfSFVOvjdB3FLV4K0ddNGkNZDD9gZMxINPlSY
2IxtEvHi9W5WJvWp3/hR597YX5Uda+pkGceIPs9LwaS3N6CHL56/LONx9pt4FW0J
cI9RXqDv8HMkZKfAbpa2dcgooja8ML2ctru22ieDthNNaX+PVfGPpTcw4/9pe+hl
CHF/ViqvJNMOuDSUW5TcXTm/sNEZh7p3/lgneq9HviBJcaFtbmc6JiY8jionss+Q
C9zYZdd+rd/42Tf9irx08RnAtu2BVcn3cEFMpqFBFKkEtU/NEmrPG4EPKigCEi5j
OI9KdD5lujN7PTfTBElBfebLeVVpHFpTc//S2oTx2EmxobosvYptilVuvhjc0RG0
wO4lrxldCmC7jhSO/b1zJ9l2ETf+S4x2S6o+Z+Guyl/sgB4Q0dNbx2jr5S3QWVtt
k7kWvKrtLG1HQD3bDLFxwqBhTjun8/4jKuXwSqU/9wdKFPC2h2/Ut0gpGApHy//+
COticmWEhS3eQNp3A5iTTEn4Vw/zkIKy6MegveJNDKeo4TlUFcf9wAb0Vu/Fn3At
P+Ril76JqwTYBTNApDUW+0fsesLgTepwo955EWaqyHGrwU/rvu+wyq54xTsn+iSb
VFFA5XaGduEwUo9JDEauQINdtg8oXxmoJ9RPpjFTj/lBadrT8xTaDGCxTiilCcAm
JG34KvrwJ9FnnESDtdPCItN5UndCzF3csf4wJuLfGJTJ981JQTl2Iamr3NOzPZFU
YnLm5MlzXsoiUXD51zrDWwUw311RLIENimZ24/LIVlAikhor5CRjpecMf4H4ccaI
K9c21QNihiSUhaWFSkFK/qG5ctnFeSsTroJb++W4qSje1LVG81FlsI2UYFetXQ47
Lc0k0wAt+90ZDIALNpEfcU9jPFvlArCusz/vlPC52i8zZYHGutsQFKB5ekrkBpDs
JceZJA0GihkLd+EwxgVpxqfxN5GY5xFhZAmvcRGteRfrMInpesXWmyjnIIliDAnR
C28rgpwoLrIwYFjBhMxf2NLXrFYp706TbS6Q9FyAAkOaeVPgmJz1cb6R9H2pf0AJ
Feuy+ufXN4hKzuUYoXYZRweujs0JIkW+Dwo+9imYzq1pEZ06crbjXIEgwpIrDdlc
qUg/tX5P1JiU5vsCzWvXAgBTqxIvr2023nyo4pyA6wHMbJ6nbWtJi1B74jpGc5IF
nish3ErDcv7t9yDMP02FmcuyS01VE90OzwTQypzMtvh798TTC/w2DsBERg2q0Js6
MZ+zjTg7oErxqrCW1G36binKkPwslpucrvzNOWY4VcyXi6PxSy45UtQ+OPfP4Ob1
QO1y7+NKTpdtV3l1pjDB5VBdthcz8ic1lLSyPtlzL80Qm9oROz4QBGbUlNe3IYSl
bgvr8ymknmh1yk2+QoAMjOHdRbJ2TVTZGwPo86WOfV7DdS9UinYNn0IUK/ZAJNRy
hs1QDp4Nq6JhrsqNfRqt+tkGQP/gcQlc9jfspl8UssGCPUboiN6v4gUkAfKuHe58
AQB8nLeXwEpr8DkMW9bjfhv7/M1Dzbs4VD68IcuTmAmLGHPkaOXGWpJnEO7b3YpO
hqPXXBJOhchSMaE2QhN9KMHsUCf9HSabHfNDI4+hXc+RgVF5d4M3lFrzkCUT4hyg
LLL2A8n8Lg2Z1BXvXJoliG9iD5vy5aIX1UqbNwpOsRzxjczy3OQBnY50uXnrhhVY
EDe3Fo8GnGzBLtbyxpWJ+4C/t6o1sOMEmjdYOrd1k8w/xmOROoA053DWKAyjAw6e
km6lc4nFcyScms+mX7G+yElIqaazQr9nBWN2fN5nXsaV0WMchy11rF3Xa+DvBNw3
h/9uoCrSQbrEuI9nkESJkoalT8o23UNMrFZ3fUICaxRcPuL/H7Qq+HhkEDpK3qP0
VQ2uztVMryAEEp6n3ekjZg3uPNQGNWRJxNLILtmua5hXBEw92RYk0Zw2vc7Q+STD
ocl3geoDxscvlZmikT0yP+PlF1b/znsX3tzjMVlD5reIiFZxX+u2XbP1nZ04V6aP
h4hCZOiPIS2zVOSJjm+7z3AoYFEmq9mFfNo5UI98Z+UveKAQ/y1/0v3ExM7xhX64
2Ldtjyv38P3CHpjXy2Lf0ug3N4h4HjssJUAE0TdvGYUOGOZb/U4O/fgdA14xk35y
jsDxMID8K92Nnbcm0jYs4ofb98qezvnKLYrbiA6qguwaEUXjWHEKDUU3jZ0CT0Ve
rJJVS+tvlTSgra+lotfK0bqYPzvrT6AAU/m7d/RW+z68RsX1VoWYQdevUUKrQSE9
yZ270q/SFW2SJYbiXZYe1VtP3Tqn9hdaGJ3PEb9ijpcbCVuTqTBV2eNG9AlOPODV
z/JazAMV97bGD/hpKb25gu42JGd3C63hdjDWur0YygoWlH/bZzHeXvssBKco3K3u
tNlS5EqxlSTgIzQ+pCAXJ1G/DlzTKATzjL1zxRMCqZhxiJxIN2CeifiNfEq7jfES
3V55WNKw9Ki6Usu2T2tgGyK3HalXGhEIwlqG1Zf10YSAfoEw18etYCiFtz49luE2
yL+RylJWWhvzgQc64HJUb5AbEBkuECvt3nP14NDJcWZoGOP+k3bHTAt30WViTEUK
gZDsImBQIv+b1e0MZJCrikdXmwN6J3LMk+qfgN7i1HICe24P78X8KqUHC64X6EYF
R36Z9r4WdaJOCnvunkRkRAV0/ym2wgaB0nBI4EUtgfzN8R+Q80qrnFg1cuUUGv19
lVDRBE/YIhFBh8FC/MtkqsywTSZm0d1OBKHZ5fe+LmSfXkfcjzbPMpIBbiLl+2HA
+2MGXkYxBOkjqzAxF5pCSGyLa0dMLnI/SMdjtmFav6XDNMyccJfdlqLRdrFcDjMy
6osr8Vx1ZcH/2L9K42snMYounmxcT/sc4ZYDKMq5NFDb5oxmSg4RNi+F01kAKgaQ
UuFkvC0afD9UszbXNqRXSJPjPZXuIqLtUcCes7T03f7CZgHo0rzH+wFRjg9VWFli
tLqzrqCS37ajpfeCZt7tsQoIQ9cepe/LHUJjjI6xYzaEaquCiK4xOjOSEHORdjWn
oFAvDGloj5JdtA4tSMTd7ii4ypIwG/JjedF0uGRJyF2hthsDfBbQ1exMruuBVNkQ
O12hHCPFoX2L/+bybWvb5Lk/4v+xwnfz2V9dHchoOX50ARZosmRLuBfiUp6rXIsF
6vhfyX4wP1mZ6Xpe2YlzvKdgbJ29XJ3M8ip9iWy8NDfI/pHOx9k4j1wTb4L82bqy
fwvC15bYL4CQNdhwe27URlKJ/b4DCOojz2iqwDiopf9xsKPMoVJOFin4GUk+HORm
3JGqOgRISGaY3nBi9A7b3YxDkw0061eyBq0eqA0Zppg9RkC4xJ2JCQG93oyykLhr
7kxUl4b/sPnI4dLfcEAIdbQpEp7/awxlA36HowMCT2oB6YwfqjxX8ANoUSRgSM0K
tKgXvl9QB1rzfHn32tFCc17kw7ArKxfC5YqGy/LPOuOBPkAHwROQNnP9xrFrQQ4v
cqVVZAmKaHmL7JgWHPtNvZ4+IvLH8VvlAtbLmXRfqGLtjCKZS2oaDx0vMxbiyoat
wgjcNC8bavfzd+8L4mO4vdnJSnHl5HwLKrYx5fzmT7JOO+by1HCJ12tVDSbe+cqB
OAZRGHhCbJG6qAe15QslQMz+GCEi+yts+9o/DZDY/IMAixGInjPBiJVKq20yZdYn
5RMpE7wEoglUt5ikkS1wSzyX035Bgdo7lXR0uM0oZsS/vJix8+k3SZvwh26y62sQ
Vpx5icgkjbKFnQvHPgtLQmhxfCXwKE5boY/zm3I0B1ZWpleqGU3Ku71vtcWCuqY4
eD8s8RPwIsqb+O8ah18wyxUJxRG7ecqG2AWA13ia9CcDFOVCPGivLsMY+HMfY9RO
AppOCkMNIt8mK7FhIzkMoZG/q3I9uehEeMB2dEAsnB0VFO/59L4O0AIUBhNjV5ok
aG3OjDOh7ZJsDncO27zdrVT1AvVC7EOKsjav5qidnrTAc3j3+9O2MTk1viv+1KkZ
2EKxSTnnleOF5Ldo/OSGyPcdHRmuGyIC2AcFZ5C9Qf4+4SoMTlNQ2pIX9IM4lYfK
JC/WrSXhXNBn2XbAvCWKMVjIBYvey2IgstNnVAfCzFNH/e12MVSIFfjY6q1pHbz/
Qw1fH1X0jjVWpR+sD+dnh/rtiok7WJrdPyYjjp6xP4FpVmztG3tgGmHUEPSAucLx
TniyS4MCqf8THi9IgBlUxtl2paD89HdEwBnjkl8wXtO6NFci04UAVWD72FdYK5qB
HXWRdJWreH5oTwWjhKg5o2MALDhYFlQYRwkodvE/0v+5ePaabHXoxlV7OY7KZXj9
EiCWDBxMnmMYIcs92vzilB3neP0ZxABIQ2LX85QYmnTxWyu4PHMzahsgdlMqrWJ7
JTaxpkwMDkOaKAtH3UAGIRhqRsb2TcFjRzp7fMNYkfOpxMGaKAnV6TUZ8v9Fli2C
b4uX4znaRnRK9l/oyrtbsw8r1Q2oeb+/PdO0BnuTd45fWuobGLrIpWPdISZQ+V42
2j8HZt/8ewKVWtVLhdGIZpz4xJv9KMQ/gcCHtPHHCSXP5cJabW38G45kq/nZySuE
N03Q7CHfRg85o+sM8QIoExnOO50S6UjGNzMykduR+HjpobrPw8Ww95FteVE0UQ1E
LmKVmlM8dbyj6l4UGA2W7zAQjXJ03/BrXNr9QLfXhGCJHwE6z+06qNCXRkuP1uip
1D/yXsf88J+8PEazvzD3BeOWtY8g0WHyvsK8Js7Ehe7jde1jBh4s+4Bk1bqBZU8r
Mk4kP1yz3TLo/tWG1i0JqVBo0T2KGYXFUseBzzqxjYP8ZAXUwNeoqmv2NxFY6B6V
nydpgBnC8b5VShN8H9OhBKElHfHwhhxdis4xQH2HgI6Ccgpfdkr/gzJYIDv0jeKB
Ig3rWqHdpS+fvioRUfvzUxDU/6ZOe7/tilkmsRgOGdu7aWqQCrNO5O6WxyB1yGav
k8xKPVqNrflO7TyeM+a+ECRna0elFAkQ0FMLFnisnjW1J0uisJ4+I2GZ0o1dr8CE
I7nqgK+BXN7JXP4yX5jpplaxHgE2zIY2Fdz1zN44DlRfBpDZGja0OXguWsyGwBkW
cl4rF4yeZJ/iD6vp0o9NfEdukMvJgtxGHx9giicK5QFw4krL/diZr5O6l+u8mBjA
qZUCnCk5IaWvnpgbo2UfV+nEXzKlHfX1XUwpFZgeZTj0gXPoS7vdpP6AoUjCZyzz
SsQzv3+Jv0cqKvM9ULJthwIiOwjA/iyyziSBAdX65q4vP/tJgR7wqD/telbSXGg/
FBBLNK61RsjQeTgtXgaCAz5bb2orS/VElrHJt8vj2tmEC/ZNq7uIxEPtFm4eCwAK
zwYgLcyWYpt89Qg96n5gRKgSh76o+HNkuG6LcwDl/S0PSPlTun+AR0YyV2tJPkCL
lUCFPsTeP3gXIaxa//fySKg7cCmqLRpMsCwcH8S0PG3SA2tx4L68IM94+yUTnd7x
WqyBN2t7vtrO5jGPbzee9EYqO1IlO4q54pYxNf+f9uubBv3XnlNGxU3abOVZ4LO3
DJCq8NHPS9s+29S78KfyDu9C0ihbI57bU6P7zdVi2Ags/6/5xkqOSO53optDNc5r
C1qqznOkORJECbHoahPbWVOGJU4Sj47/0+WhB92qUJKrDFGz3xOvvP4Nyemd5oCM
Dns1wPLPCza5ePztWCxPF+MnXKrcoUQkGGB+YUN8MDOTRoU7YAb6/XCK++r+fcmp
Ocwfz1GGDErFf229FeEOur4eRKOEcQVu6a0cpiOYB5WWdnbrxdIkfsjAqVrQVNF+
7y1V8hSAhFBYFL7F9RsMJ4tKZ+eaF3CxyRWpOkV3KOTNPmIdNpoaJvrQP/c57WRo
qpQ5SEXEUp7QtzDrIvL46uG1+7pE256NX1bJpRgGsGQZp17mELxJTLow191SgKwk
gO7uhk475NKbzc1FaY7ydq2CuMblFZFrwlY0EgP6p+7+3shd0U5oWoskHU9Lou6H
TF+8Ef8YHQAUQmcOdCitl5gcGDzizpgIE/c4Je5XP5FdyDTqArC4YnP3ClS4mCYT
J38nY2oE/f8bAALoo4Hi3o6z6DU05p1Z6/QSfhtdk1aAkS1hrxST7RCvb0ECcauL
5ohOtsKjWvIm0jTltl4AzulQqN3G4UnAaoG5RL96/Zg48BxrtVRUyEUgCCD+2x4w
osndyf7U3MyuYF5EXnaQd/d5GHFAUK2YYzzG3iL50nSZEVCePyDWvaaQvzfedUyS
2v3U2lH2wrIr1vgs5VqWmqlvJvWLK/k+qWweWF9GIt8h41jbx3HHSn3b+/X+viy6
KPrJSEnaVLjfd8lMWB4ugRha3oEv24hcbe3Hf1BRMTeykJgqsSZdD8536Acy4jH4
636ofATd7Puf3WbenmyiAx0csAqFaTqLo0bJm4IxQyL6OSxONfCiCDDFSF/kf9ru
5KR3xdV63b3yCoIgBZhXPng1dUDw//GLW3ccFJHiE7kUZtJMkvcts/l73ftA5Qg9
4g9Hhos276gHnjUSkwv4/adu9MXTUnMAF+J8G4rdmPu8QuU9h2aFR77fTGzJv/eW
p6CDS4S75gXVC8POyqpIWaxn4EwVWH9Y1e/LwRMYpT88yIobJ4+bP2gGA+No7ae5
r+yXWQJWQU+swd6kSBlkJ60dDuEDpLjippjI6fajeko6wfVbbfB3Lhd57j0jktxW
JE9xekVJzbyCG/rko0Du5AsQrDJF3zwxeyIYg5adpOqz0pYK5ChTlE0UABx0D6P0
t1kP5ZPhKElZY5QBV6AbT1WeHSEfINq5BY5LDx6CQkxxAOfpjZCAH+jvkVMN9Ih6
cUCj9snJzHveJzUzhSp+0/z+mTfq/6IeVRvUAweX+Qo6frANmd1YT6jrWclWDbf7
VXT6OnU0jzvMMQR11JlaFpnaCEnWeK1W/fDh055oB89fiK9HLCLfMGVMtkknJI4J
D3m5PPhLZqjyNXqrXuCUJA9HjpXQzTKDpwrtwHM3k8CxDcwcdW384C7xNoTY8jPA
7bmUx87mfDZiAtveEpuokYLACNGo4nfNlmFIghFpnq6gbImC35up1DD7dWSVDI5E
xZA0eUx0sLD7EHji7x+Y70rUJt1AKY98+7ZS8TwdYAKdKYLR5brVDJjZ8t6jdwKW
iu9vIGuWTFn6565ES3WSop67CnE39v/2T2GjWUnTrc7FPEu4ciVfxwO9AFXkIR+J
AEb1LdS4A4S4k2zx3k5U0DUUfbq6sJKfvvR9CTDvTZNcUZXG/naYDzQLedZV3a0Y
DyOe6y+Jqu5tf+l1jW74C+lZUZKrJSJqfHa18THI6RcQmLYrvHxF0ZW9UvRmo4/Y
Py19TdpkRgWSGeZZMTUZ3SnuyYqtFXqaUD2HEPlbYeqOzmTJW6CGJIlO0rk3TBD2
uX5F2UYaVSgvPiActRVEKw4V6GymVtvLIPmQfsih06JZxZUGnVQmipUmsSqh2H9k
IUnOXLNV22K8jeyyS2185oMQ7CPgZe4zoEOFMG68GXjFvXrfttGT4u+K3oQ3b7BK
W7J8wwZj7mMcufUvugFoxmcbnX1BKmgNgDUj3j+aEYa2LMkGfKS06LGbQZSDDjbi
Mbe4zxH0X7lqm+skY1/mrZ6VygqSEUT8yOcRX4GMm5GxKKuapuPqqsoldWeZvGAA
/1iM9dCkn0nwopdb1s430Z1QxiQD1LVUKUcmhdYDrFQ5EsB1g4T5sfvN1D+KDG3m
+pdEJWR34H0MEjNFrMm7kC0WonlqIY57+skZcogTKF8ORXTzyfNuB9AlLS6CBraQ
fZ20f6WmEJDRVJ0JOXvO6E7P0Q8YDYCRnyoIJmrTiskJYQW/e+M0pW5DH19O35g3
lUN6n+MRS4F/DOH3A00v2d1o9/furvHA7T5geVDsTGbMSjnVe0nYSNG03jYhuQAr
sZY0+izxc99zDQ2OV4+mqTG35IRf080oW2mQLz0lAT2VwID4nc4WqpuNiZ04hOlq
Vz1ftvK+EBuF6vjFXA51TIXCKSsYxMgWOVefyWHLNU5axlI6G80GzNTziAk7xCqV
KKSMh5mOjOCzEjdz3TkUctpV4cG4Qma6Utl6CTBSstg/8QagOZN/J2bxlNyLYRbT
chwjDx6HjDCmuEQ8I7TkQFGpbpYkFBSDJZiVGQwMXzwP9IYfE746swD7lVp9GH2G
X85XjFrBM6Fa/D7p13FthDwgNqY+4ZaspUYVqpNjZ/QcSIHeB55dnY/rri6z6udg
IFnn8R49+cfUFaX+fgcUcY2PiSy36biEkFGivz+jg4FLXZwrXthnc2WiESQXv8K9
OeM9qpPAAZKTFoF15UxVhu4ASGGZz+U5dc1GPbNbG5EVahLiGMRm3Fa3oSunBgQP
RCfwkj+wSR/1+or00S/IAv4h9aohvVCjPoMnV6HqCZei134tGjSORZfLIlpWBdyb
bgRkquTdKOZqCcEdUv9EQWEnTujl8Pyi9uwNRPTUrjCvg4bH3t4xKgmxJeecR/VU
LkMYNoexVBKrBNNWjr/SYPOw6XkFMnlgkGYIlLFOeH4jyHrlwcvB3phm91UYrONp
nsWgRFVscDn7/yr9TxCMNf4wGh16DUr9008CkMYLkTumOOHCpjyFeRQSyVURjG2n
OCVHRZlE5eYPPdZUz++UT6cWLOhK0ugR6+zhIiP004HQOTur9ebRIsZWRBA0y2OY
6WMGpfcKAXneCu4K5lg0rCu/SmDZZej0ScC2nYuv8lvNswyp+DGggDeKZEs2nKCT
06MVu4flU75GkSSokXZnPFUP/a6YOBOQtSQX2KRsKjF0zZSYcL9Ekr9Sc9M3oWXc
BjB9CG9Ha9UNyzDSN+guR1tw0BA6eKc8R+buF0EOnDtrW/oeOA+0q4v9u12vhYj+
NDFqUj20d9zPcfs4kJ+c6Zeim9mjBn/Xrb9cihDRlddRbUm29iyzLK9P9Iaog+Vf
IuI0K6FsHSWnBWs+gulWJYwe6VhQqcU5atbYme6oVx2shj7wghyNEP51tCwq1xlp
71MhIoBHQUXUc+LdY25CyNBNK7DgFa4hV3lp74elvcyrUkce7QBVW57ReuQIVBoW
nxfQSY60FhRxq2TyLHM4CQcj7H5FbHBfLTvrTOJXCrQLhKWfmBtJiYU1OAWSwjjq
oYuSBWgqS08N6IjvQW1s5jb7YFUtwxf4LcVUk3zx91NE4f/s05RJoPeK0nUD277z
HtcUV9v8tOf0sAJGbUhSs6K0mJTQY+ZbPGtWlGVFZPvRwfyhmR2vbLd2QuXMDZRH
eLuoPjrJ8pxmE/PJr/4shNWI/y+loyGUVrooSYp0z7PR/abX9WICfZ03ROC3LrCE
Qf3dqrU6k5b7hQtNJKdeGxLmk+eHYYG5H46A7tEWR8//fxB/5oewXjlXJWVia0WO
bDhXNbeW6+iIbyJzXRdL2k/MSsikPHE3e8moCCu3gSzKH4hzUhGjIm8dvrl1rELv
shfw31D2Blfwid5AK4izivBVzIylFfojjsu6xHWgY3ohWpHrOQkr32BYOZ3iBCvO
Tzdy2EgM2+J1c3Gvti+Vef90lyAjrHc7tLXBrU3rhueolDQptLhMJN0AAhrsa3yd
YRWMlJNeerH8DKo53lm1hnTPyMk8YEwGe3Tm8Apb+P6+wagD5lDRmce2rGFRVjqb
+hs1K7fYxYHncLRCwRGr5SnZIdHY8ER/hdzbnq8TQ0njSVcjN2h47iMQKcbKAYDz
1oQYqJwAjKA29+Y4a/o3zff2LTkNcAJSAvuzWTsJyMkzyR6rbSgXf1C0UZm+U1Tf
t9AotjmXFXhOS7UuUvmcNR0PXvHw4lF7ZfZm35LP3UUgHBZeI8tDSHH8WUyKxX//
1S/q5hWyGCO/2UTj6eJwGe7nJOI9fFjeG/gZEcysFKyfD1uVnD3DIXJ39RE7jx58
RmFuhKuVYEfs1xIaD03ulNi81A2O6XWlE/FcLOntpI/BhjlAsKsYHEYhpSr3kZJq
kJeZfG9p9s3pMvPxciK8Q7Ryi+g5LwL/tjO0oQs9sQYBLs+QvVnYPJRo3YvJ9W+X
+nyUoMCLakAHuvayoOKrvbs/SP50Y4jyWG0eu/jrloF68v9ObvEKSdLPMfkKmEMO
DJVumk7DcziwXoUv3xc+nK5QNcKrVKroy16A1pIrZ4KGk8THHnFwLrzsmX0IZJZv
6jyaMFhBGBdEpPBgxI7/I+yMn+KxftnOElse0fODl11Lcw8ZI7kg+7WUhIhbgTCJ
ErL9WFyXOvGoI0HGm30BQYubBoH2yFL/GGYQaVkAOd/JuUu4Agou/Es4pHLoB70i
BU4vt99meFz1PhZooDT3murYUxlOom0a5arf++Dn2YRlCXLi0myaT8MUY5fJmoRY
QyqwAYZW8D2/mn+M6UR+46pBAPggsAhOnbyxTsYgE28R3PUXCBHOF0fMXjDLuS5d
zVojo8EuJL881K38i5NbEK61BFWjL288UaWKjygJD0SJfwMvv/ZYdE794iuANXE4
OUjTMtE94YMjG0uLFDW+1CPAeQknIZBLj9+C38/GFvyttHeVpfzEeHMTaHfBrqRj
bckPnrU35opUoE/oPzWKv9UtwMDlp/aTOXunWGg5PQRTR9JvfBKQga1MzgS2RDa5
WKUd8/OM7laQIspDADhOl+zSSh8iFBSOvrjHFtlmIb73m/VlCbr14RHLYzfMNFEm
rShgEXSQhcO2YA0LR//iL6MnC/ZrY1VFQBtcOE6g/0os3A4gh7bYc1GyBpaZmUKL
Y4BzD7z7Bq4nm1e2Qf8tTF0mUxwKFTuxRzuptkAAu53EU6eeEVAidC4/mGz84M/j
M8AZjFIeqE8b05fZGAqbPS8tH3nCsEELDws01gdzWUmmQuEuoekam15xIvwMgbzo
7YspDwQcIG0ARAc1kzLltoEAnmqpklyoGpYPvPTrVVz0J6y3r47OZvrhQnEhY9Ib
wJr5s6QgLsA7eSol9dxd26g7SxA4KAx0bcb4BJqqlJi4jrvgKDWk35X0XGREDNE1
mRpEEbE4gVoktdeBMYiYR8QsMfwy/iv7+EM86xKwxGUNZewOUwnh/xyFcPytAufG
4UBsTFoTIXgxoAJ9zC8ueOTSQUHuxN/wF6v+aaDoQ3+IcgYKXIuYfpJEYS79JegK
BotgFiiSZzqsqU6cqJwD4OGmIzo6AUA2NbhwgtpvYCThpxbRTI5Dq0jnIrckOWQn
lBUYAnPKSG/jS2YOTV1uByliOI6Zc0/2HgnJE2NHWYuyNqRbaLAo5+XaMFird8cV
/rKHPvT2yiEcQGj7cPs6OrMzu4+wVF7OD4MM3tmq18B0kJv9HqiNtj7QSTnkFoLx
5odgJ9wiezrVCyqRSReV68uFnUosOunu2tAjJ1SoMd6gnOI+2wkHy83mKNk352DC
wLni9uIqy0NAkyYv2TeeTktFBXK3AZhpQgSkcdK4XPYLbd2oFPKOzdKaNWki++uK
UB0mBOhwhxJi4lHpnBDefGNNq95OCqseNUNSr42ImP0vDi6iGePTh1GTVu3r0oYL
Eto8L6CIQWUyH1CeS2kiSJ2bZ0DsjohXNRDmJMky762vRUi3T3SI7Z2W3Amto+zK
hJL1HS65rnCuE1PZAfamqaG4vtmuhbj1yN79Ipt0/9An7myp8+HlVUdfwT6WpYQl
oCNA4jMZXt3tWUNw0d+731ZG2eSx5l2KOv3C6eUYHvxzQjH7isYoC4Czwhka4D+P
Zd2ol/65DvajJMzRP62BX74CWBX0rXtk5zldfxfXzR1ixWQHKTfHf8BKj/YE+JBn
mupF1EL8gjHbexq+ENKGGS6tm51uXYN4rWrAyJ3DBfu8Y6QDBTqdDYcBD4ZjmUI0
iXHwEVRhYhidklcZrEA6DtC3f8IJblNKk/n5Xpx6hTHRuzMA3gFjVO8HF8s/7jpL
yBiajEVlEeA7jy8uOtW0giE0qTR90EMoBQYwda+JzA2ZnxRRrgESexYJy3LsTVoy
sPFJV1vaUoR6tIyFyleNw+Hq53tk9jfh6gJftRSfuscaqNjuj3RzewsyRT70ZT+W
07XMyooFz+7HpptaDpgZKIwSWFt9jrjatOjlc3DsYzFCaw3+JUDLsUaYUoYQjdyI
aEJDq5MkAQ2qb+4Od2VmrhQi3bt37BIgz2yrbFW0RoLZ90y7ULHjT2KnF6YJMDRH
ExFf8f9edNqLgEhobAxms+5vv7LfdouXh+E4V8YqCc7fpX4ml5ENmwSSOYs1Rpsy
CgSwwzlBbDAdcCkJUJwV/YQLjKUQMtbomO5/xgPEJh+hJ/eSWC3PTr2MicViASqH
vK5HLGehafu09V6ivZi8xQRQBe1XB00FoxzPRTLiVurE4a8k/Zn7rUABNwEHK8JT
8ikE8iwfAQdaaCMl5lnQr12MeFUTJu3D0nVereorO1d2Gbqkg/zOYrJJ4bMkH9ag
8uewqDJvcOFu06J+UZ8rMvzWx6F81iiESa7sU33dDRaQrCfHS/Wife5hnWYFs+nR
jPKS27ErRAw1aV5ii/DQgY8t3oA2297VGJUaRts2bvjcWmqnnu3GBE9g8qXms2Vu
Y3Qa6WXUcRwgxR0GxWAY/JKZYtZF8+fC4cpUiFNpAf3iax9MFTQuKA/ZPMUcKBw7
69jh6QQWBQO6WQVx4bvx9/4c+b/LwjvxhisOOMqLFkUtvGqOJogwfXUl0oNEm39j
XDZfuYF25T4DDECN1b3gBgRNqp++rDfyE4KhgYQAxGwsH1xygxvRF3pLhOMn9GH1
FlCU8SjK4v8jWGQX0bocGn0aObBbGqx8qlHaZ/F6Rhs49GlnvDqUAg5/106mzEsL
oxd5jXj+IawqIwmSdKRhoIYsumMtKG8nHpNDYdXmTxliRf8narZSD4xwDt/NwOew
1DraF8QqY2G70IPY6/uGQRBKR9fr5/1qcr7YVRxygOs6iUe3PNXU5TFGH+IcNJXI
MJtWj7wn7ymBgoQHYVaKbuV6rBSqyp9q0w8hJPHsQlkK8ge2Lmz5+zN/hVhhRAvK
YSj/JJbMMww5aCVKR5jgBCvANEnWv8q+lWnpKDWr358N1KL6I0DyRuOxTMn3H8Y9
diJsLcPrhbI7zv2F5T92aT7t02UAvHOH7DI1i8WduGmALicO8Uq7OvM2aVzYhCdo
h9XKT53YLC/Xqsz5qB2XSzX5lXL+AOzrJW2/QyIRNjQyvC4Xr5rYLieLAdj4czoI
Qb0SG257lJYtfANNjxjuARkPZzxaHjXWC0t7Wj8q+ITvK1xC8pXPeGfbaPm5GhTx
gq+8LQZUmuNv6s1DO5Z72XLEPuVU5KxvBHH3kRzMAFVnrpBmzZwNBYj0w6t+OYcA
6DT/YQupGmybCBzaMrPhtaoNvwkGBQvGagXUQQAsOQiyh52EpkerHEqNWkEQFM+2
i33mtV/YGFGN4BvyqDn8Yar8uCPDtQQjxlC/MppRLaYmuQ6/s8m+vyIkk9Ul53Z6
pftS5peqPHXqPlkNFJoZPrPs0s7jH3h/9lrYdbunu/sadCsMDbj+QQxy7dVD102Y
kciKs9w2hjkHMfZTh3phmR2VWoo/psl9y9FtWVKLvPlOak20KEH1jUd6iaTZfXeE
R8l0zFtGzriBufDTesRRR+CCJZelm9X1ry9Gvy7TQmH/0J6z9gzgNcCdMBZOtJqg
LhgbcfrpQ/usvgzK1W5WmBcfD8keJB2bXXGPieSvwuFBIXMQ8CWmwuAjIjNlvgiS
Kh0lRgW88pHAAQlJ6ZbxkQyEvuwACxSgr0eftEIpGWg3HrWebu6zr325bvlkn1pF
i9ATA/8jmLgBtkSw4kLBKNQCbuak+ykA+QZ9hv0Ajd6vvqMu3jBR9f1ZbHSmkk3S
D7UxRAIPs9bfZnYbgRdkezL8/vIaSazPn14k/TdzGVXsbXmg1NT/4x4UOijQmeoI
BtthgXVcixbC/xuzLVizjtcWT2pcua83d/n8In+ehQkCxq7xwwBG6FFbiDKtkfY6
VVXjMuTnTFc9/ArP5pG+ZQLTO3BarSt3wqyv4eqRJlYQv7TtI7gt/jw9KAEHprZs
MK1+CIy1IEv4pPwjabbe+aSeWJYZiR2UnJl7KGWsfOTWzn+JIKiLFijdw3DmIvrV
4bfmDAUl8sqweH5d3Yn3hEUBAocREq9aXLG3ZoQ19JeCbpR84hHCohhUKV4XAghw
tnfKEuNNO44NvImTl/DDb1jNaAcWK85ojT7MW64+fS2gjVEqKN+W8g8T2VaHzDQn
amWxy83K85kCwYEXp0azKSx0tdM1/Zwm6/aVEcY11UB2d3DvX06OizmurVL5Qs2f
TYZrL14oQ5mNp7jWRWA8WfqLP3aDJL+mT9Y4rS3hxlt9CpJQGyd3hKmmyLHWff19
kfs4sY0yyF4coaEDjKeh3kGW0hTamPu11vlBHJhGuSFmYtICqIvnw44kIQjztXc9
V6/8SmG1Z726XBMlDJI+4hL1G91ZZlxd/FVmVGMMK6RERdbX/GZvg2a2w84av9kn
CuyJHtEajCED1w4ttSbd8QVW0Xhpk5tiLGzHkXkDbfjzab2WZ+iWoVzoNLe09gw5
XBIvya9CcVMR5/P+bRSRGD9IbIXOsFc/iTQeGtwTG9hgk9eML7/CfwPboLDs7/EL
VaZmDaenethp7broZU+ayHM7aUzb7lIQ4q4B/jNa6B6WHL+Hlc3ia2OwDvPrOecM
Clw6l/KIuD/AMdlNPnUOM38qX5dFj2kgMHXbrKNTQswpfHaGiwyT/bKRx9Lge24g
R5BV31C+m5WdpDfcg8aHv0D7LRz2OaH7ExfgnxEm1gw6PjNWYIcMfyLM6m7dsd+b
rOa/4wHFq61IgN4JUP3yZcWJ+mWYaAaL7xKNjoCxzxcMO7r7lCFxNl6xLWmNZdOo
179lEFP7sAdaKxNXD2EXD8CTuAk/RoAwNAtDLbNGrOp3fMFakdnlXCLaiHrG+12W
Bgc9nJFcXEz4yXMUSqAusa39Gneg1qv0lTpwuAqUSj34KAy+Z16196bl0PM7eY4d
GhYN0uABJlXrURqXDznaKlCdQWOTt2bjsVSgZ69tUq3I4/2xx6aXkMxYbd/cKetl
rgegGy7X6ep1dJkMWRGhms1l1IfrDTJ86GgTsr2htzv/ZLMlnvnZ4ZTPnHvNYRYl
ZcZn5QS6a285GlsLG/SHZ1guAr001Fx+sv5emJkJU+V+OfHY1uLWDor6DsBp/nQq
Y4j0Ur6GqYg5oob7P9FoqOTR2f3+gRQqbf39SGmtsi/asuBJW2J4/GIehSXa+q4m
TtajpTtosAx7YG5b+Jaw1NwWMeXifM4B81999jPjUlbcOge+QuJrLtqgIfALFW56
xX8cOlz3pqAgNzEKdd9JUM4CqaJ6mPtj8XpxBoZ4H1n03mmtdz92gCOZImjNlr9q
64NotSxB2SVdrrxRh/sUOyQ/GAR9h11R/gt5QqlHsx7Jk5/hdTs3riWIaDbTs/Zx
1ZBbl/O12OsUpDWkb2/w88KlRcztgc1zKTlVvMxOUv5GLJRKSGNiyzryLNDlBAjU
3MdVY5OBBvVl59P7fO6wGtnRwvVpE8yYpHZNq2xwyfO9LOVYq6TI/nNd4RWwH576
gibKQ9DIg10bqFnM+8KwDMCn/XH5JRxqZc0JSwpfJ3bY2TTGx86iFThWaZkOgmEa
jCET2kb8f0e30wn7HbQmXLFuq5TNVSkJUd0T2p4C0pc8Jvj8CwEob8eRmdVtrNKx
zMy+ohZ7WrNTsDwfYO1bNwMoRFHPZ19Ud8Vxei13kk7mSgI3yVHUH00wfDcGwYaa
pNq7lAGCxOMYdYTStbNlig47m3gde84S3uGF8xznfC9o8fyHiuz3umq2ssXUJWyE
xL2+H+IHhqPvkapjkjUeqMxoVAigTPCUIhH2Ao16P2HXLKbgUKxobz9jtWFTSRoV
sONWIjGBi1aBCjj9Ind9w1NhztBuOj1m+0HjHJwOlnfvy19bepY9kB8JLHqm/8Ol
uBVzUq2qGCwEWQYZTj86LgSCadkMiCH8A802u5fPj2D0Aoa2JVt6pXCRXvXj7JUu
IYCPVE0NnMCMu1cjDhPoE5BE+xPhy06ONU+GlAYeNbeCMJft70g/6euHuBO9xRDF
26qj1uiw+Zrypi4wDdcHWfMtBAfbbbct+ff06f1w7aMO+SVq5fsGQXoOrGU/8/Tz
BUZ8L8Nii8bye2aJ0jPy5E0W1f7PioONbTGsOwfHDQSpXELVCkeVGKkhAZOdlcae
YsOABn72JRaKVDcJ0zb/+DXAz3kfzfy/XS5XUGGgD5ab7v/fNIPMCcz0Rr94hFNE
9h+qU2RCC3KPCvUC2I1/YN9e5BH9kvJVYTYKNYoJgcRVy3XNJNhhFiYb0kqot/sK
tRQHbRl6RndQFRXqhCrlnjV7kVmSWC3dA5E/X5GBMMOk7gnlDvRNx7OxuYbkqG/d
RE/3lBCJhGpuSmb/hEWKr5YNXY+LJoz+quRUGH4FbCZWdXPcy15st1ITjHeALRjk
ZlyNrjaJdwjFmQsiX1R7AmuHmr8luTVdK5YHU71ru/NodyfvtpiJLS6KFRwG3qi9
4NS5OO0BsOVHcnbmR8mYDYs5/7zKoCNF5BZCv2+gt1xMfnIoILNoKLI41eWmR9p+
4ElElkw3Xp6RWWR7vdnLS3ZFEvEaFVaIxqEtafyUGi/aa34C93MEtfE7G3k3udJ7
+WEUoMpGHpdXDTL3/09Ta8iiAadomegVoH7pe9U5SX8AkMcAaT+5K+vNKuwIb3x7
VP3bkSa/9aaPK46/P+UiI2LhbktBRb/u/UVj+/KdXR/YgIYkMQcJjab/yBanMIz/
QQxGQ4XDfOvx5kPygkrhkYwqk6w18/zc8UNVIhxTxG1HCiCMv9tiSP57m6ess2uE
hnpbp4oyWVpHyr2np3lHFEd+v3vgmsUoMvsFMeOEd2Hi0hV/bCp7BQ1C82hwZ+DY
mv8wo2Ihdqwljmd65eiBvIuI/neYxZbu0Eh6Iyk/SJhHGHge8nAq+h984aWcz/y+
OR5LSWR49/T8Pjoya4Dwjuj4+8xoeV9SihGctWtPKHDFfwbWRcu8zTjzLqTrqk3L
Z58ljPAqOmFTrnRX7X3lehQ37wSBbuwkxomEqqJJjLl6sobmKZ0lyKW4RxUkj43+
Hey7cQ7OC20tOH6MR4S6FQCIwmKDN8Tet3jLcOHjwHc5qmgnCgr3kJzyPY0276Ds
5r6s8gMI0QZBBZr2CajBqnNErTO4xOIf6BjKO3UWlFsk/J1qSPhAJ8hqFxSX5Vws
QZ4CH7DWu+u7u8tq6VVyIJwSPxRkFYtsiugT1RmPCaBazmjolYWL+HvGSLALghqY
FuBKmWNbpPmlGaS0tFtLwiQPQPZ/PrGIOqapVWOQWV+MeHj3O1WTBcpE5fSuOKMO
vS73zVtNaFQTF5B5SuuBcJSJAOHHWZYlJxf5OJsZcL3WZTYYNvog45QHQ2DmcmuD
wPnKUiFrmn/WTYZeAKhIHmoKKQZ0WI0VAW7lGdJysgaKS8eQbrZALguyqIPJnwN3
8mXZ5qlfrsgS6Yh3ujGh3A+zzT/uJgPVehjieA2SYYd/ZXEXCkUVCJV2w9g6QHzb
U/mrnjXb4d/Fw9nx6dBsOSeRculc5D30mGiNAIB/G1aXhqsy4VJFX7QgKJ42NR0d
3EtdOjL2jKfk70qBiWdAMBuSk4T5pqQpOO1y248x5XEVJlg/CXAd9y3P3bqsJ3fb
MhxAxGrZ2hA7plY9X6OUoW6g6u47ppBOfbUL8ed+tbc9clGhEwUL7re4a9pumK7r
tXZ3i1sHZ3YDKoW4SMMbjpDHYtcchIJUrjyOT5koqyManzKi0OGhLhPPJ2iv2xrY
a3SqGUDnmFY/S1Qm9JcLeiqnyabdGKPpL2GIoawR5pNi4tTlhbcFSjXo78TTVdJL
RKGvpvlVFGtlz6TfwEjC31t+guLS3xkoP7P0TBLALzZUjpeDmW8+ArAydPwilL+y
hY2XT6z1ppo+uVl5OYC/mlB+j1/vLsprEZzBE7RxQMiKP6BTVc7dAa1CReRW15Kt
pSMeVa3MJ6fRS73M79f8+YOQMKHqSKq2WkVjnjN/xSVI1Q3+ZCOdM35bLygMvZrT
u9jj2GBefuhJqs7WrLi/A2HhQ8vHcLVjh8kOJO1j0ElLgcWW1d+tAPmyWBkrE+xc
he+qxx7bn0nJNRH34+yDVJWodrdSbBPjOQxyynqIN+cfPSsym9SVbHjU/8WK/5KJ
NVofibfWfHBubmK/VRZBwgMQ3/cjQKjj7xy733QSK0+gIMagzSKdUWo0uq1LoIAE
0RDFC4wnnuoAShOPn2TdM3vQj2yWj5DMKLP3BCKhbLvQK3/Ty9IJSVYipe9pRy10
U9h0cK9O5Xjx/eBIWcFn+FQ0TLWJblHsAhXhztGkAR77vxWf9PSz3SDGrdJzrObo
ojcOQkb6OHB3NyjkwjQBygD8vaAGpAz9OkHAGQn8OjJPatvTw+K5nazgM63swKeE
CLJp2Ox2Gmjla61mRvqRJXI8jO8EEGEm+wfk4mA3u/t2U9v92UfpD/WPEOtDMomM
4mUbhFS/Oilty6drgC0GvldmNeDMZm+JAXqdEtUJGN/guir5JvtTcyky/X5qUsAP
/CCfkJVi3Me2V1/thTydDTdz9Cvc9nwJgKs+kPdQjG/sX6/BI+2azvTcktmoEd7E
EZi+XisXpE/xFSgCT5Eot79KzdH5p9wz8boHritmtPCirmKK3R2WSXB32OOk9tsA
ItEimZ7f9buMXpo2hn7//9UwdY92Z0lXk2gI02d46ttfrw/dhKuuQNG11/VnyXQG
c0zqF/IaPxkntRr8RQcV1NfH/pCPxX9E7i8SBRVKJqkLwX+3+mejEePz1uUT8966
gjJNlS/rBE3uUHUOl1jOQiudRGUswzg3TtMUhrs/kSs/B2p8TQBgN3eWMXfXmABg
Lh0uabKlgTLVRkAbXZkb/7I707d92WuVWmlmlVce5KxzROPuFXTt25iOn92WqZjU
pItXuHloLeP7LmA1JEwQNHUFCWwbcDd1cz0SgJM+zLe1tGQ8i6+BLqy23cXl5ZZL
DodyZdSYwxitkmOZR8ns+QTJXh+FoMZD+j2DuiZ6Z5d3bNekqaS4neziN8xzMEFs
Msu4OScslFROAtqOCjvwUOrUwyby//h4X1mp2MM56Oiv2csOTa/mPGwXr7EKgelB
3l7SIW/ucjIMqtzZy42G5anyMmxtPpHUbFVQoDoWXd97SCm/HeHD22XObqrihsCW
ilwZvqXLiIvdbt+ZPKEptV5FmN1xrRdJ1IhuNf+R6C6nQaf7jlKnKob6qdUf7dzn
NsmLTFjI7ORYrtPxgtrSZgC16hbU4B9dtul80Gur0bg8tbjPy2HNwMFvEzrMBmvo
m65lJUEkEjUEq/fYdx38c2BlGLZixUbPs+Q9X5fIurjq5HcNwGx97MbH0JNvxfJn
kahTLu/2PDgaQLRne60CUm2eddh9mAumh9gFoBhO00ZFibeeaU0lzbsforU7ALcT
40if8J83rlNIl5Zd7CT/+YN5yxfvvL8ZRWByzxuPk8McEDKW+no1CsXdaJDOQL2a
R9HREwG0zX4GO48Qt5ni8+0AZWYjT3Q1+sYbSvLLFVH8AWDGoynWF7pF+NeeeT/B
AfsRt/BNH+/Cg2wHXgNMutgk748iJaKn4zL9FXX0SHmO6M99vequIgxhhi50YWxH
VUXzMWaNm8b3cfWGg8mqxD/nM1sOorMJkuK8BfLQILUzTZooD4GZp9K3g4dE85kl
FOQRpMllgGeMWXd6bFUjMOtonITE0KOm2hkPRQ2Bq7/diqKY5LE7IV+LJyrew6t9
5hgif5sqpd238CvJfUcZSwpXqNTQ+2nBdh6NvT62G9PU8LCq1SEegACTQGJcB8Ww
rLb5freHTClBrHXCEO4Zbt4ukHUjl2frZj6DKfHggRcJ4qhHniy0/c4xA6IbMELK
nzi0GcCHaOAAgsJFSMRHv2dmV0ByTUliPOmik/LcpZMZ97oCWz8R8saI1L1VCjNZ
vshXKmFMlw21B5yZTvcf1e/QxbiD3qycuSfH4RvAFXwfwh2KtNJXmvUbO9sYvyiI
VneTaTVUYTC2zkByCG0HzlWc3Fi6cNjaE7ilRuAI0CYuO2Y23ixSI9THiSYZKWNE
UgWrmInYhXOA2+h9YdmL4OPn8mXdWHEYod+MIAdcnwofdpM+j3eUvsd9J6CM25Vo
KYmbbzUok6RecAcYMzhVtUhZb+autiUz7NqnEYkJ0ZC26Wq/QjjdCU9UWhNRrv5x
1mU8T/gMuMt5mO6qi2bdYVprq6LtO6jJk/YYFZBJ/zDFHhdUqEZprYUEt5RoFNrI
y9+qOQ1xEMYDHa/o3EWB6YTwkPO1CZ/wZYi4qjvLFmgxLz1n9ONoK15svWc664CD
DU6TOt0lC60t1CIMoYYTDEwYQ9Lw3+ODAnwNshUD78/5LiHsAkOQxpLJgcvxx99p
8rdc9/WFHFsA9RQQcx67YBtgHwHXcRmLbWsY4y8OM/zpqGQaoANoZNVww2MER9Dq
4Dx5eYaNAusYNkI+4sJyNsgXd0lfUhfgaiqcbWFm+nzrp4tiftZ+GB8HQWJLfMLb
/weD4EA9CpsXQY2qBM1IdwS9CLv0+czxORWeLsXRi03DLDsVcI9+rk59niMMZrXa
X2iwx/S7NnIJmK2BdmZLWSf4caSHAYv/1h+WBtCmEvmQpuW/c3ITMG9ndWJaOag4
46x/IhxFeFJe/gNI7rWWbtTkyKckIGfhuYbFcuK3/nQpd1WgdFb1HMUAhCd7j//8
Y4G5FT0HVdn8xi0RMifjQoYs4d16MMPcguYCtUj+mph16X7gRpzThRt2CKpg/pi2
TWhNHoyyFwwmUDQUeM3lQOD0oNqk5VUWRWDhVHhZ3guSmGz4EbwV15uBmHKCurYJ
dLrn/VTSqGcGEvwGSz1+1BHBPikrWY7m4BqEzLGzwzo5+GKbUI+LXZTkSxQY46wQ
ZcmQvbeFhkwbwt34RZ8pQVwZMnJMCnE46GCUQciZuIdBjRjySOppFdQj9BTjpMQ3
rh7VVO2MOQr6vLuS12UHijXe6tMCaUKbxG0OMXfGEo4ApPB/LtBIcS6X4Qodaf16
JWmvs8vQ6P+P9c6hJ1ecSAagribj+1YTIZx1iGXxgIlk5L0u2WcNGy3wWPV6wH42
56uFZISBYN++5mUDoje7yr0GyupJN1nvdBSIzZTO05QZ9RE+o6Zk/AQMVWNiK10V
5wOYk2LAfd4w9vDPPZ7LVzhQVVilLx6w2uZxIpAWnykH850ZEbdLHp7f17eF6zWO
lzNflv8g/cALw2D0xfNseZbQ4TVRtquyvaPLzXLf7INyZTElDjAGrCoDTtCgv6mA
nGq7vUeAD9pnxz9i8kimiT/7YL6bxwcCnbK/DYNL+smvjIS+q9QQ/TDOoJnixhhn
ebyzGq3DghbVsF8zjllbg2hByGDcYjCkazTQK9LcWhfmjL3IlFgYreqNTkUuju4s
lPOgThiWXoVYS0GBno5fSEnMpoFzf9AOp+NePtYvfAO2b9F6X81cLaURWXfVtQVL
G9N5RVzDSvE7pP+DUy72gb1N3BGYxJY8bfoQPj9NjA1mWymMyeDsSy7fe3eN26eb
VHkLocTBoKbO+ese/K08LD4ykSTu8SrORhkaLoKpHoMbXs9OXSIFdcDemUaGeu4z
sSdewFQ712H1tctLfkRDVnogYmJ2+5AhkcnTbBukYMmvUXY5QYcl5M1/o4B1pi1V
RszBV5Rt6fcE3lXTNunGFjxHE5BwXzflyDrLNe4Zp42VjoucAdu1qiEiOf62nKgZ
E9mQclFmls+k9KLCNTB3WzQORFbM8Hppb4q4zTVFknY2Om81ODjd1x2pRgBklnlj
ZB82QBMEVNQJNjWaesW45TcujrEAV5lNkyl9j7ROQDQi6/a7CAakTdxagPgaaeoO
aqXWDqWv5OP0KB/4q+0+fCVfL23bqdIwaUfy+TB+/SQuhzZ5uZryqaaBXoy4+3R8
HCToNKl3gFm8ElzMy9z5lrhd8zPWEmOlG6fhOz+8qZrvR56RCdvqs+lkuKDuAwau
TSQziHvRK6H025Gxb9/7u3y9HeVOwtwp/we7xptgknkAO6Vgz/i7mJxc5xSiW5gb
+Q2XsHkBjmT8DHGJ6eMjA9uK5WToJ1t6rLuQOyzp+v+tMrhEvmM4ZzImK3E4r3n/
kU6nkIEq4yrs7+ZsPKR+fftiq6Km7YBNrAT+4nO80y5i/LXvAP4AJhWhqx7Qsw9z
yNy1zFGsRx1WGTGj1ZLljXz/qoG2PrbWBfWnIRcoWa6xeZKULzPhtntbq1URK1Le
RfKzUc8fW6Y5JIip5Wk7jPxoNiTKi5kVTRScZwXLfHIQHDCxc65c6mPbfwgLflkd
zhg5L6GX83McUchoi4s4OXA7QU+/yvFRKjprmR+e4A08PxcT7oJmDH+pz8pa10vz
5gOT/kwTHyfX/49epLCjkPG9OVeknj9wqynmRV7S1zYzCZZIeOCU8PO7fxHSuzfx
eRDFmYsyrclb54YZUOpL4efCyOdXqMmQoaxmUVTFiZK3aSRjF6fRR7GzFiS7pqN4
in2u3R7hb9ZfVD1OidVvyaUsg9M+kWes+4ZStVvN/CpKgD1i6sf4HqbwjS1SDbIe
E6MJ0XbIT89gbISiwWgehCwHbaOIXzTBen0m1+iN7e6beewsA9LbbaBc3mUdDqk4
Gfn/PCwLwXQbOlO0e4YNJHzAxGi3h5qcoPmcJ+qkGB6wPKHscddgsK4YxkW1/Ev8
nvGjzC+uWvWa3TMlJ48eoWKMJM53JYvqFJr+zcvaoFG/TP9SFNcXDQuJM8YaMyjy
3YQRpi5JsSPix4f2W5Cnxa/GhyACu2u4NyiUTHkIYTkt9F51bqfphzZedErh0xCv
P48kB2ieRMyg4GZzKVeOU8t3JhkcHtww6EACOvu0aTpZS8Qo/TMO74TGpJF1J9CW
jg/PN2rmwBgvIP/qWi9hUcK46iSg/qmIRlZysk4sqJ60eXv+7BdSgb+8rnR6LddK
j8NZ73JmUrO7oRTvnHxuKAvZVxpRACUdPdEqX+86ujdqTA8vDZbPSY+niDQaZXyG
bfxxBirP/7loXBbCROYQWLQ4s2Jh96tjao0u3lI/7H4YenFLTCfGdQRz2EtVpjeJ
9QxTF8jiNtHPXqwOL/j95IADLV+Hnpb5W4+RBntoxscjo7pPWtms90DupeuUEK6O
1QsNqHL4KOlIZZ8KDSk8rGC7uBelJoPPlpeoBqPKyZIO6jM9aPkfwwznW9XrC7Ty
034zrBL/QiR/fkfqx80HdEEPzrRdtO3a+Z7nkcxyW5TfeD5UuiMiZGpAga0UdB5q
aC8ehuhYerK2+50j/T6EooMg6yv5nBgS1DNE8uCTlYyIMPVDWduKpx78dPWVGJH/
h3Ht4tBapvpLnsv53WrshH2iGl4CxqhhrrRhzc1yTnhHiQyAl5oZfLYi7sPbhBeb
fjgfGqbiWxMbLC6R0SlivxxKsrW3pbDGcXPBYnLXOKqCejncbJWq9HEZ7N4u2OYD
WCx2vce8ngcV9lsnLCKYQusBArpjJfnUkcUG3RfPp+O1T5CqfVDqj9wPlNdrLk/U
T3WiUYDCKzEtD6eN8ibsmZwxLq4cKOuPQvRaHMoiqTng+xjD7EVk8yZGKp78xghu
clPZ68sNTVTPSY5CwZj3mdj6C252y74kM02J5m4FMDKWP0INF7oxsMDxxXL7yvA0
6ajMQ/ckmk1wchyfEAuMY/N3e4qsznc4Zy1yORyupMz52bJCMfwV6qHmvJDm5ByF
VNeN7YQexmQbq2i+8cbN8Np95eHvneY1WsJ8iCyVtAVBid64jCaAm/0wkyOTRraq
WUEdvraI2lHdF5pnZu0JQcymAEMoCptiiBl5zFEKRbFjZgwVfQa16us8vtQrupgz
fdMuiaphSUUozk3R+Pko0ZeCO2JLM5J2ucuVugabwJ1XQLVB/tZvTuV1hkXaW+18
Wl80VILrc2CMGdK4WT09xBTGekhN0gT0zcwE/KFP8qBMbAH1Y6p/szC+UHlb0t/E
m4C8zAxq4/Lqn2GBoK+RpgxfxkLR9DPEilF4L4zNquQT+TMHb6ASZ0w7SECD4nKk
lNkl4XU1O1BEfKHbni+WZaPqFHAuljlL7geuRnitp/J0CtevjZtVwJxPkqYFGYNB
84si5zdXQumPgknfJBkn5q7BRpALkedrGfqmg/3qmtTlnQ6MdyZtP7H5k4b7I75P
q+CHIWb63FE9xvum5AN5C9yMW1+UQjPUvuAeR8SvLeH3/FQKvpDofrAz6JCJPuQ+
/Brc8D0IhCgIki3JNTaRkiQs1/fHSTJvsAlqehZ186oMgR4VJQe7GarkAc38syfK
yxiLJjWaOqRxxk4C5KlVcFfJ0/FW6UeMOhu66Ik/d2Xn96MakAHj7hsqCLDWt+Ez
D/wSCn3PbV74TQcCEoZTrvXQNRyqFDZxGTsWPAZsOLSyIbDz6v+XtbLHb2PUR5Tu
9l0L6apleyDpl2zG+L55jxwEGnNww7k+tDZ2udu7Gbd1QrWEcXZ1aUA7mzgbtBcM
d3ScWKxaNUFKmeqGhCTcZj4DKCItV8p8Xdj6bHTCGSiYML0sULSB3nNo68t7wQ8q
FlRJbOIt0cAdM/3oTr4jJ6DTzt5Td59xCDpRb27r9pXeBG4Sc8koSZH9stsEiiXs
ao6npKKzjNObpxgwAf8KLgDbb6KRzmxINL4BI8/IWtaSr9BVNijelTmSIhDlS6lf
KmpgWnpj/Xr5m6BKBLFC8N0BGCjRhJ250kr0jlfULGvgoNEKhpa0pruHoXWRyI08
bdYaxx2dDRppJwwO9dmi9qK864TUH9CwMTiNMD66wzfqB7NhtRcdyg9pFlsLY+lK
oWEI0BYcMnIxv39KLbnzC6aw49Kw3s7jRjp6RrwA2usReFiDW5BHpwnDEJAi6BDZ
Jt5iijBEVKiv70r2pnuF0gk5fCONcVMb725CRWCbbV3E6WkxLBZ7q9LtviiQIzqL
bg1b57eD6vqx82IE72UmBwmZu/8oVO29pJ5R+v6cPqQQmhAyu55DCdZ2oSLJzAqo
TiCOBL0J/9kwVjT6gmhHf35USRDBrKoFz8CUzef/zyqxzOZzXA2KzJDAflowj9G2
Wl9CHkc+pwJk90el7ZbwtsE7tV2C0MgWMQC49hFvCJw1iZS+DkglKeiyQA+y3xr0
WosTHufbmzYiLfB91ERE/vVpQPwXSpaecX8yJCACedzBm3X3UU3S+W54lqiWfwll
qFTcdQ1fkwkqiFeAHjlIONuyY81qELVRhbxs6/LUja87h1E8H9z1OY72LREBqwwQ
ct2STNh1FzQLrK+kVw5RPPMlKV2yClpJm94CPGQLj0afOrkHlIJddZk9M2WlZE5c
ejxg8oTlOMGpKzpM2dfCXOoVSaxIy3ZyV6x7HXIKFIyDAQBwTi59inFSrlMgqD0J
SSvTHIbuct/HfFM9bN84igXowAyjzBGcyY9cnjkmANIvARzjivYIyoOhCOM8vq29
E9fx4NAylmRCPfU6l6+J8JcOEQqJ1QLN/tyjHuqREwCgBHeiQ46O3+ldjoWiXPAu
MUH5ENsUFxGkOVgAlvXbYGWeld7nd+d4RpSRugss2yGJH06EnFCHL/39ACB57J4A
NDoOnIAyvSwbQ6z7pzqxlfWX14ZtSIQ4wUdWM5Es7kLR51HvXcsiRyNZaMaXj0Pf
tVVKGbTiAla+QoixBs5TeBczvu/dWN6c+gMNuk974kMLXScLqd+NyKKbHpBdXkWq
/HYYcTZXRpZH7DJDeo88xDstkC8vNlPanPjRkQB/eFK/q5U13kxAoSw34p+6Y+x/
hcqMw15TOZyMJCJp5/EJiHVU1Cqq1AZ3UiCZZoqUriM0BLILyPNqQDKq3wK48PVr
9V0fV1mw1oMBRumJHBKeP5QPsp28pIYSM6vS3iUG7Kx93sVFCPx8HLL3r8x2Qfnb
rwx66jkaU+w8i+lGonUClTbG2RiO4gd3Up69FSIG6/omqDkz+rGUkyMKYX+CDnNs
v33BjudiEg/RmzTMaN0EUMuIzEO039ADjOkwW8Y7SC0wGck6szpoU/7joUoUhi+F
F11UanMdSUqyuYUY41adW5P5RRf5nVw97BP6ZD7Mp2yiMIS72Lgj1OVjzZvduxyk
sW5IalK+OInWSL3NGPI13lluz9FHxREFcytbJlTHlr0Gk0cuTaj2brxfiIsJ+kwX
EXorrcuNXsGoJDjT58x7XTC7UlSgotJznG2+b5Pp0VUTXlndvthlMW/nwPiANnnZ
x0EzD9bHz7M0SBrjfU92y8JKdaM3SG/5XoL48HU4BiCOt5C8KbAY/AVAX18vQDyJ
BPCUguDpvZejpMrnho4IaaPlCKpUMfCigYfVydqTP4VJ7CiICs9bwlqoWkTN/NrI
X+6tPZ8JFun/YJZFvc1WYtAqcIfNcyha+055/qhnkNVB2Muly9eJGdKBRAyh7hme
ijsh1kHD4Iq2EacZLkZmshKyONgMZNVI/tsAchbuaSE4mLnHnoNbUApQxEDmAefY
s7grHQvspVKyaKo9ptR+owFT2l/k2SR5pOh3tAhw8JfpUxbBGZUs0npTUfhzoHA4
Zl1Z18hKfe5rk5X4V9NmsjQxi8NgfVQZut8KRR7QWhVa82Sm6oFCLMeaWcx8r+ZC
0vkNMATRtMBqF7cg+g0qJN5iv2J6WMV0QUHuBU9u9n4reVGMUhbzqyg0/73BYwwM
v6kd1ux8xSIKJMPbg55+kss/YbPZn9csxm6QDyS5GAZcqjxtiPR4pmWZ+r6Fvg78
6XAqG1pfw99greSITMpGIRUkr9G0O2c3FBhm/dSOkL9tR7526UZFS5O05kEzH7b4
SuIdWY+zZ/snlcM79NW+QQxw+yxKjZA6JUuJj4v8C4PAu8/gifj1SHenm+66bn+C
H1pySID9fqCFUhYWn0EI5QclrZllln7FCDMcV/p9np3NCS01vLVSGgbZiJ9OODHE
J1SG8C029QLKNKbeIyiB57Rzu5FRsNZN+DJ+90Ldh5DUQ+rFX4c+arOp/VJhnaMt
mzqP90/C7ysvMXX/cKaa09HWTBYzJ/7SzV8lYFtWLZlmfYroi/fKWkbI3izVpysC
50gfYA7tHmc0RUoIaP09mwVWqEEZtTF83C9skD68zAmK7/Ab5sVg18Zm6ryAdLKk
QHoUC6rUrwv+Yc8AQIEG7xR97Mhv37EvTgmogCbWdcLNh1+2aNXNEZ99pgHDJNbr
GPNN2uQJ3nmCBOFUohsJrC/WgGDFP+TBBKiBhrtx0Ia2x5QtqgAUo1c2Yd/0cXWI
MtBC7ixb1VPrJsXaGdFJA4nTKLHvCtPKeRKGW04G0mRt4DeCUz4/WpALHNGaRGeY
lv1/hdAlzZbbAHsaLsOrmOmxPieQPa1H4dIy5HwSv16JKW1dJr7GuPkyoOSbZlFZ
v/vsVwAeGiFHXAXw0PcjF3r4MnuBB+uK/WdEFmGtD8LcfioJEwXRmu+6/lJBDbq5
5MKe2/fYUS3GXuSBuvHAGYilEBP2B7RO6YXYkyEXzzU0Q00ueavHmty6qfkUVau2
OELsiGLhe4QzKuzyeQ6vGFbI0+JoBVPxz2Qq8iY8uNLRllkNaNiHPEyQm9F917Yq
lNiCASGOEbrSgX8dSPOKJwNH/dQusO1rHfRR9lQFwroEd+Q7Nm+CVDBRzKt4ykAT
1einyJbSJqcQE9CRdLVxQLhWU9+/5obfBIOluUFTv4MuL8JIOiOxh+aR8r4E3k1Y
FbRoNB6qxdwEHpR0WKYgUMkibJzd9NnwmltXHGk2adm+L/O07DogGxrWZAeGLVqi
6Lti93lJk7SijwRyaVnO00QtBR7xg6h9ETq86R8oo8dmDDU+iC2f8SYAX8At5daL
xL9HXxD1c6JHmbvGEteywtVODupPJPZcuhNIPoY8YiZKxFFkVOJPjeH8/aSpzOi7
gcYxubgL2SNUr8DM5XZQpActG3D+qNP6DWRfzVe69DX1Gai1PaBjFh0yd3wyYHmf
lrwbqNaGwxImxlcik94I+JKN443ZslylOSYMTQ5y47dgFFhdz1Lxi0dXNKRvNhCc
KOhzDGGHEyCiwLWfVcgl+xLugQ4K9pVOEkwAowCIH/v/SZomAQtaqFpsvY+nU5zt
yEZbELbRXvfwkSdEcx5myeKzIN9uVa/EgwLaxoM9phjDFmPWCqwJrCpyeRiZIZu4
YDohuZ8CIqVB/mhisEZdD9GHPueYq6Enu5VaDpYn6G4gUvzFU5q08BtEXYh5RO80
6CC+URgWUQKnuVgj1gD+49Yu9JArdRAx3reyhqUbBM++o46GptlrMCsE9vnygjyG
EaANwiz0+tiKF2VeqVnUHjRzwqvxwJIb/13atirQDjnfZlT/P+9of7pDDhhF2PHQ
uZEYr1HrGTYrTW8anpskzEr6npZA0CTGnQmXY5YJMrAK5Lr09tiJk02ADg8JyRve
QM6/v+02ReQViLsfNrEJ9hLhBf1/JbGB+PIhCEOgNz7hE5mZA3QR6ifuQ87u/mZB
bqjK8Vkw3E6fsJdvqLnNo6wANav744bH7FnMnsE0Ajfwz39HH9LTpZ2Jm3B0ErbA
BxMwv8uq9Wp7TIU1tFYQB56uuIf6hlZcii8m/APfJ2s1CuZpklgYAx1XGS4R3HFr
ezQ8BERBbAHM0g4c6FSNx92LfKMud0C4lJNIoas3UnbbuojDixLTrynBFHobXYk2
AaumZ39cH9hGdBw5a6tY+ULk/MjLHDXSkp4N7H1m9JyyO31NogXPPlDIPxT0YLZt
QCuz9bNS92BDKoEYzPDm4jpMmqWQNPc/I6PDd3HmzbPylShVPX1zwHeVD2cQRvkk
c9WHijVbMF7Xdiv6yrB+kYGyoVYI48bZ3dmLLs4wC033fKwwWPkC9Rap93Jd6cLh
4N/kFISRLMfRWKcjMQpMv4GXkc12W/eOnx0REqo2Ykq3x4iekgOyg8i8dZDrkWoC
AY9P9dYJ749MVatc/6Abdah0JVXt2YjCJSFnvB5ynb1OyFqEZOPvj/uueocCzEwx
zx8uvSzyuLr2oFPmSOKlKJm/y6/g+98friKsGw0Szq9bdURf/Ds13ygN5NqLRE+7
fHXbqOmdZobf6wcKm61ROYMr1l6w5xlv3OsKuRmNKADMHZWs2Q/egbwdOKgKQSfd
kDpuO+v9Th63earih7wDAkJvZi65GZ3ZyDkJZys0buvqILge6fJy0TJ94QuSbw1i
kZDAQwSUUfw5XE4NMKEjKT6m9vBMgYSr84WRATrrTNZ8ZNhgBnLThZt14F7t1jkd
XamGJ9RBrwEhy6+ka8j2CdlaRShtCjG5do5Q+1/eZ+p7cpzTrc5egcdwnlFElugX
j3FrgcUMGa1vXIrwoFjbYty/q7vazKIxBtQq6cDTnotju0wWiEnFc1Dzh6nyodvP
eAuzetQE8V5BCPk7wJDM4P2qHragJOuDIz6gB/zTi+l4o2LJR9tke4WL8bpBrwJO
TQhASub1HH+aKiA5VLBuR6HfShwSzFm//Nl+G8npkDxO5zoyapgwEYhGnXefUjuS
Nr0jOkgYMNH4PRUpjDlP3w9vph+GBjNdlql4/22OwivOZRNzhm91UVWndaUOZN/8
TA2h4t0zRclbWWg2RXD+mDuB/6U4R+kETpFGK4XdR8IWEgaG/ezctl7j8Om/oNB/
oFrPfwbTlqc1r0MdIuaiNYmZY++ZiTuRTcQyc+x320/ymnFPQ7mDyzHUXOvrVTT1
F1VwctuybjwiUi5ht3l/ipvszrqItcEb2O6JZDUtmgZSr0+vsyOaHgDLJjhBtfAg
6dwADX6I1bFg/vMzx1HqIxKkc2KaLF/riIz1ezLbKsOsjP/MomiEXK+/C11f/Zvb
dOvNanm4LPFNGXhuiM17W59XH03jF4vQyYZb7YndtNtchrjz45CgNgYAb9hY1GDb
LzlVfnc785Gs4jh+fmTsXmt4tREk8PWCZXs9LAxW0m/6rrWcgz7QtpNOA90yEBWy
XNGGVskQfUnBT+IS7H3M4olCQB8lu+dns4TcVeAIrN3jnQlmkAEsEbz/RXQN9Dld
/e/WCjwWCdQK3D+7UAPUrhs4uYxcZRxSsdbfuZp87NCT6169bUt+o7mM+D7Qx+rl
hJ/l7zfi/YNOqsf5WUf28I5fz0Quzg37/7I5wX7o4PgLGCD7+hVmNuXevYWu2ixr
Krt8ZPEUMTuxVbkptT4qMrShRl8QhdEkpoP4hsBtuosJyUA6baWceVJESsTQPkRD
TzFu/CEYt/OOFw8xXXFVWsgRUOe3RTda5Al2DXTna6NmQ4nHD4UdchTrDIlw+iDH
RT4D4xyH4+txdBEVC0mVcL5pXfy7ZI28xsRo4a+fZX2U9uOtQHyWslA5WOuuV/Ca
QdRntMl3cv55xJP/cL63cvrm21T3IFYSVL8d4kgqM2Ga08kw/LMK9rwhBSba4tLz
AfDb6xJutERfYJ8hDalrti7HcCXhZd459y777vN9jStl8NkkdcHWj/7uvPtKQwav
YjwO80lxJ0FnMBrTciJ55nRM4YPj+aMitHA+GDT4icmIKGDvgNJT2hG/SrdBk9Xx
wROWWPUVF5GVG2zfPwC+O4qY2sfL1AewGgDs916wQ9DI5S2eWi1nEuMsrn0pQ0a9
46mnSV1f2PbMmEH+7TYHkUtzhwMMxEUbaeBZx+OzhWfAZQupvMdzdwQikgTJl1Cl
+9rVuND/j3bgBSNOVrXxE/n7LLpWbPZUv098+9U3x8E9Vy3I9L77qAQ3J59x1UQu
p+qk2B/7p6kTQboRFYdWMsfLyUmGa9GTWUVcLad4XGnlSEjQlJoyNVr3WHH8ALrt
WEvyAkEW5EvUxH3LqVj7Yxdk+DlznA0f5YsE5THTw5F19p5TiITsCLTxLBKXihGX
koPelMkBgEztKaoIDVbAcP+7dZK3AcNHcHp7CYv76V+Ur00l4EBWqGRBEog2OH97
qupJSmLayqjcNF+WPNENPCi6ep9ImQSTNtEgid68K/y3oAtxekuCYRx6ZexL/Tua
0OfyhfvWsXuiLNW4kwqSD5jwsI9lcdIrePEQ94HjsKvP/PhOfYYlb008GwO9Nqc7
slddtIfmQm3ekYUlmNdMQth6P7zkfrbGw28THN8vD4pN/2sQil0HrIMQi3Nwvz94
ozNgAZOa8NbECGF13OJOK7mvct4MdqV7E6P9J1Q7upblt1I5phDJ9xn4PTicpGGz
uKWr0ludJcBbGXLbLKUCBQqBsynyRiwE1PBSp0KkHFVticCVisn7egmaauJkuvzM
izXLzdUi9vNSBVUTBOOo0V6+iHwIwyyS/SsomZt0+YEoGn7aE8I+PPxEo/TLxNS0
XFAc9qQINAjIzzrIA9kiSNhsgHnVs80rpxLpY2Lflxv4lcEb1KA2EC/dVcZ5b525
90dezbZGU/kpFBPQNXs7UElKMM5YpxmymyNYw6g2RWlZdKLkD3Mb+dW51jWw0NHP
7rwp7TH/tkNZ3ay4nQOvNcousMdPAaBZBWpXr2sipJnIVofcJYasBrc1YvSueVlG
9rVPgjous/kFN2M+LHD/SxVPb3a7kWhTZrHMwDLbrW4BVjYlTryr9znBc3NkgTUU
iuGa3vUIp6l8Y046MmNIc3B34K4/mS/Kw4T0TXt8Mw0cQy168RvbWmi/L6d0uwA9
8LCwS+2dKOuxY1uelZJcUxdP5VfBi2KwxTbSL8un2mtRIXjDttV4u5tNi7zmrfqi
PT3C8LfiEs5TF9VNG5waYa81+n7GcoT81t0n2M64MlSQa90QgAx7X190FOqXhiba
fmR27fBu116WlhJo3e4hAuOwnUUvJmOSJiTDg2F61r37kiacXYAYb6rje6GvxYRH
N6HsmZ/8RGr9MZz1a/gFSheSCMvqSg1S3mN0Y8Qy2knjNOPZXnZCPCIS/0m8Jh54
7B4Ov1QipI4XAeCua+L83TGSEdvrA0q5OU4BHM96sYatzvtUzPZxUiJRJD2Elgtq
1QymMrTc+XZ4+GrpqxiULTeCbuI7uO7v2qIUQcWqeSZ6jQailoQgmGacGcz5rcNY
tFiZB3nQrZJW3Tma5k9bReP5GdPujydsmiqJbHLtpOWK7YNfZZQU7Cgkaa00fSh0
sgNmhwhP6PVc2ctRrvJg+fT8suqX1NHt44kc1LGW44IvrZLVfdqpgYaUdUX1xFW0
ghVbC161xjylFsQkUECt7UrHe1RyY6515g1rZ0IaXzvnOMH/fLR62cVjmISQfpbp
h2R+cmkQVJEUySyAFB6sRWWHL8j6CU65m9U29MWpRr2H08RKuo06dCJRslEE6evt
63DLxvPmfG+FxlD1/8gcNB32eWBLJZp20xZGt+j75oZG69SIp3HilXmRpqyNtUkl
xVNoZkPUXIHOdvd8PKCc66kCHEs2aoaGYwsvZ8PMTwqJu/tMQYkpkXwZhIWkrCt1
W5CKEsHTg1wAv/SV0sfow9wlGhwnjf9J8bU3l8zJ7ncXtKXJCtJIKe5Kpi+69ARK
Gk1Qga6bZo74PE2xm8JKlX5HvAbO1igiiFARE37kUt/QbF8owCriFC9SVqvpfRLE
VpChVGVPs+ranCS9XpAmosy1HrlRC/9O4858Gs70tuj0XdMUaEp7ySa424qQWbHP
N/xLUmPx6OgZd2mdTE2QcJqt82v23TjRwslTZC0G0W+Lzmy0Smg09dVPfBGO7Uqm
cHJ8cg+Y9vCuUunB/Q4/U7FgiqJcxZAGhoYmdy0m8QtFLvXJHNQy3zy0V649++Jw
Dr0Py+JNukQLTXMDJ/ox7jujJ9zZAC6Gfex9HPa4ewHsWJi4ZB876I+0LXGzZJ9E
z0EyBmf+qJXNyT5T9RRO0LOFr0UUzahjFviL0nUYyT1RxvovJGRN7esEJHVpyZ1z
mV1Xi03K7DSr7gEy48Vquov3Rj6AEuNTBqvUwWl9SSFgAAiBhNGtSRhoQHbXKx62
OTHG4RHXYPH5QSdadRQDZoGSM5c8jpmR9LZcL94wyBoE2RiCWRR8iZJJ0k5nWXrb
8rBsPQqb42mBmVzoErpz7FpUAQlePoBressXS7acRDyjwM2rIjtB1dz9ALiYKkve
QyoepoGm/OTePQuzBfdz5mFWF8FfUhfvqWeJIdTqiSzWp2lfIu2Qsb2bQJaLEotu
o+j1JCHezkPtiiUeozt9bnr75jiE67LQlwPJemFcBNqNlgYhcktAlqSI/oUK50W9
quW87aDy8X3jyR8VRqjS/CiLM7Ptrou20IfUjrulQDoIFd9LHw8N/uDAoTLWl3c+
WJYpVNvcwBoaqkbafG1vLAD1SqNXT4FBkPwBEXFZZM3nnrvs3HwL/8PWqKowEtut
/VkC02+jmnqWhjcMtJkz8wAIcXP3dl/nuVYXxc6J/3841/MxFu2ike9GY1Jdyq1V
qlWoyubgXuN5o6ZNuDvFIZqXg6IWHkxtAMwxDSCaV8S6Wb+B334wsdl+jDcwuwfU
QqlfMygOjJW0HOX8+1HRJz/ro2Xi7CNZTaj7mlaY42eQ4NyFnBDrAwPGB0I5Qn0A
nUAiYTUOIDmlCraXtIJMxSLjKtiXag1fm6ooTNBL2aS99ynsIpJE6XzU8vRjmIDZ
9D91gSnjwTChMOONhf4W0G3ie4H7qkLxp9vSO66iV/4/aODrlbAVnwngG2axZ+Qm
nEcVvaZQNbj0Igf0FGsB18dalCMt9hXC99T8TocR6v1p0cA+pYjcUiw9qTr7Phzv
fXRJdHMs7nCcDGavlc1aAvwN/AoxSdHEiH87N7ZRryFT/3uHIVTuxwwaRATX6sQv
TdkMD4ecwIS7avQuAUEspmMz44y6/9bmnlvJcTQxfcrWKs6PJgILT+mbJE6T7ZuX
z4IksKigJ92xdcMFswyBDO4WtR+3oPv44IFPbJVua3TakzsgDjT2KLBLYE7Zu4hZ
sfpERiHaTj8lUEt5rL8V/CKaFY+YDByUpsWImnQg/m6+1pSrzEtrL4XcrGRj/hpJ
QpCKv1MeNkIdiIMukLIIAggRqIezELxytG27VR6lraN0ycNql02AxR+bstH/rdz6
x20/GjmsY4G0WZ7KikmHj1fQqJxAkjK4YOt+gG/TfsAFjfkLetBS8wjxU1ld5q/G
4SK3j9XbfnQ0MSjsF4eHQrwTwSDaoMFovNkQMApSJaC5Rtt9SaC3l5jwKmMJXsfS
lRSa7pO+3q96tE0AH8IcE2pQDsumYnkVtnlWTNirGooHmhjdehUcSxlbi8cUBPi/
Ew3JBqkoiVKQhzk2qxcOTKxuQevOWJXzKhzDos+KiBC9Xh+TDuL7vAwqm0PzmzTy
RI9zFsPB64wJsRM9KpYxyr8sxBUQ0rVHHwI/ClXuAIDzZB9zN+xuURggyywPK9Pu
A8CPf71ZsxIeSpVBatrNgjIE4w/MGhKVYIKbWUuBdFpBCG76rbKb/Kzx3GGDXhWk
raVORAP125XMTkDinNL2iThvIOz0j+abRPfW3XBlUY5ssF8Zl3jnqEcFvDM7M7M4
2gBHunCzlxhh8V8UWEkRP6rCEZa7xJqYTFadqZJ9JYVvNRnWmmxjy+xfRF1TGixH
9fCo20kkg75VrfPrP5QSTICh/ZJYFszkIFEyNZ31Em8giyAw694rlAoXgB89s+Kw
9C/U9GKfjFBONR6C9dZPmwAda++gVJ0a6e7NloEh5d3lBJ2mycELtTVXelsLIR3L
mXONgyDPQ1RgVm/G6XALEwKcn8/CuoDf0LDoFxv2NSFJnYd2Z8m6Tbl+BLcHybu6
jW8BnplY5TjTs90U0HS4y27R1mkKQk7YjY2NwNkK4q1Pc8Tm/CTHQ+T93n9+iOIr
BJonTIIysssjOOAUgVhjPKrfSE1f4j0PfcntuQkcr97LSCGfpUZ7adA9cfz137vg
cEDQ4Y0hreUOXUIZBaXfsIGOdDbHFS2OAQxe8dror06SSxz/HMr9Ist3VW0nlHok
2Wi3mGPifMLLewL3ZrSTgeIsJIFQKQ3nF39CDV4BsPeSkd7sxaSYeuGagguR3BVr
rimOi9t9zc8tCTFwWPKcdj9RCfxTSrePx4MfjvgTogP3OQoOF1SsYN8k61rW6Xls
BazyzT0eFMLpvGd0sozJTWJSaFLtr0IuczlWqwTPFIQUiC81nikSZcfg6NTktwRY
znqfY0lsJf1VqSPxOWGpimBejbpgMM2RIzpwSQ7lapqD9IxHyxNKzb4vHoFYpIQO
M4nNvegYwmlTg9V4lK1rR5uP7fnVEVlkFrNpxtS1JPsEYAmzn364JKG8Gx2tODpu
S6rG6Rg8XYfOnzBLzsjgae0DznqtXKOCqv/OeYQA9XSR2Crrw6kbNsqDpB0t2iOx
lTDKtJz6t4Kgb7kuABZC6lIDkYiDpeoNrT2YJJu+ZDsScTRTJJ0engXMKAo+hteA
G0M7lZkhVVt6l789YtnM9Yy5q60AgpPDZt+IoZxcJBImEFrHn1/f0C5Z/eb33u+0
yOHNSz+McoIfah5Ci1P/L/bk//hnQhpsCTvllWBPL4qW8qVs2/t9XwEtHxLjN9tk
axO1uv5PRs+EGQtAfrFXWYSQ14qaY7oHIQY8CtELNJUc+V9zDH8LShFx0yYaOeBM
xBNgjVbBmOHp2+bFj8pbnQu48inoIJahG3viCyjX6ol4Br/cvN4Ex6H6FYjOOvBo
FNL24cTevgGBqLtqOqI0aEQxOEv6dGv7hyrvKDsvUSf+6AYL2pZz9aFiM51bjpc2
hfiHkDCh6mMkGGSMTPzBEZdhy+zSY3H/QdKXF1QtyOO5+7SBhPyi0gz2ajSr8FKM
znZBiody69TzBvEPSxKqscrjWitT15BfbvydCPT8DzsUJACC4bjZTHugyr3iWbwc
U9212eLUuIcSDKZAyOopCPFY5F4DlIdxXLhNCfv8WK2a7DsOuNPHdSfUVX14XCvi
TC6zpPTFxkws7YObLgW4lc2rD8lCUp4FKqFzZ4fVqyeNPNKbx9hBHdIwyXZQfkNH
FnmNolEEAw3qeY/ZsF1a2OoZvYWgfmb1/lJnwAUa4o6lWHBQCRLGrNLrzLpgxip3
e6Tw/XRVxE/7l5eherCeU+rb98Y8EGoxb1YuuENDp45+mqPagbXyAFwr4LOxrbAM
cB2083XROT29+/U25rHbEeW5SN95z+Vu6yBHyAIk7RwwhtdwdfEf4b9x6NdlHjsp
epPFi/GlMIKeDasocadS9Rd+OjMy8qHKjr058v6G9jJb1Vo4tW8pWTaNS8JsUZEb
6jHgbUGxZrh6TlnLVLXIoRLJTEVixu3Zfjlnk4NKGFiJVlZ2o/8XScLWtf7EcT1c
XA3BjHkeHuxT5HnbpW3qT1VKVS7YNdZ7W5UGcxp1J8peFKikapf5wysCcozRs4rr
x1czpUf43nhSlfZwvOZbJDT3WMFxj3uiRMqLiHQuUVoDFhZIBB/KveRMkLNA3VUS
KAWkoRFA8G89QmcZEYXPTCvkddcViVsjpQnIBxW5QQqIp/TD4l8f/e26CnQLK4Nx
9WHeuqMN7W0fJP9rDZECgwW+hZk7k2S+zPH5J3z3ml+Bhvafd9ss17PcvkygHhqY
nAWHkBMKrZHQ9JNGjyJq/E2nWl0rki/qxlfF8L8RZqSWaIsQXofNxDuSZpU2gR1H
rVqhvgAVatigAux3jfiAZ4PUBpiZYXVo2LllCcr+WDq467NtkbQKgSzTyaISCpP0
3fNOn0PM49uJc/tTyrIdWhfPnM6d+uC4zehnRoxXB/C3+n5oDX+URy8raLtl3ao8
X8oyE2TH00dxJZH2XmhJl0oQnNQvKzYJ/sWLcMGBtzIRunZ2tbsGK2q5zOkLzb5Q
YNNA0VKR8cxqh6kV5W4przh3iblGrek0o07+cFFYiBy3k3kHxS1CyqsC2/cQWMg3
dfz8fmeCj23x5UK5uxKCsRTXKo0PCEWb5SB5X82BEv68DWs9eDm8oc3nXjbqPuvB
UxJ23PnjlCOC6BXvm018t2H1g+CWz3H7fXLNmRNyzjSK68NCFv+p3GE6+JYSdlS0
sUHJ/lINju3emVR7dF8erGCMoNPCRKHq81lr9nI6GNoz1UGxR0jrNntPGiPFIEUR
vC4TYcAoWOJjlVk/b+CnKM+SRSuxMuE3leWdy9KSVJmIZ7fgDwklyVhinN3ttieC
Du894NmDlFN05LTNBhV9kzqSoLxRzz8tilJT2U79rjQK2quaXW10Wnq8W11NoKx6
stPOyTXjogHyoLOwCa0CIryF3vIO0GWmOIixQp0qEaL/yvDe+EYA5qFGrIKftJ2F
uAajbb6vH8BcyCkFq+ffZ7FHSzQjj8S0dj6IsUSop/nt/GRO4PiOVUX7T/oM8ScZ
2yMTdwD+PbdyXMKanUaNfsJWxzptcTDwcOdLQ321yfWsD3yWXh2WgRrcHlvbPZEC
iDWrn5AE9lS4api9JZI4MDWcatMyfhjUzb9DTk/nckWmN5uK6b6zsjjl+PIZiaZl
/4dzxwssIEwMpPEjGJyt52cvy83list2SKUL2nqYgtjXlEPHPr3jstDuD32AhoAW
DBzXYcte425mAFRsE9yG9ZHa5LPKHCIl6XQzYaKdOaa9kaN+c4qmncK2eOW45/Yn
DRl7do0nr2iWCvu0ANne2JvBcqu2UEjk61tnoTIkACxQgsT0LCVKpRMws86KQgFu
BiSQrmFTCLlU7p3YlwvMTj1jXP0+BD/PZNlhAAQ9e5j4z+6eC3K5UtaCuzS8xTa6
JxEClalaNDXzmXpNtHjWdslIyH1txfYmzcyUEXXRo+wa8C0EdSfMHsJexuIlBehk
nZ01eYfz+72JFM1IAEtR9Metx6ZR6ZhOnOhnSd4mJN7olqAeeqdQMud9CUM+6cKg
CepJ4XvyRSq4hOCCytfNOR/+6Mo50jd9CgcORMKgvRiFKBKoGeVPs0lZuM0T2HYx
DDL4JFxO6tVTsrH/cbuBtJW83kluqRIHtVoc6j3tcycjPHmMjQ3OWLl5ek8xGBWD
xrD+UOVhPXTVTRaIe0FQY0FvGA+k2lgqF/72z+diHhO97AkDjzSDvjh7Ru2uGcwP
Puxi267A5PgiDxcdeldXvCQEVU687/iAB6Dy4FgWTkzeoPTi0vVBR9s69YO5co8H
oKobUfR269DMEXpdeHDOWKzo1gE7sgHLvKf535gIQZLVZ22GkddAVki21quwTZmI
Bygz2gmm7pj55ijXQj/ulb2s0zVApv7OQU0o94xesnJxjhvxI5SAOq0BLgFyLLSV
YR3yC+ji3sfX2MDTDna6nbfKJP39NTUTk1bYSkXIK94pPOJkWBa7gO3g2ruTg/Nf
ApADFWZ+5aiKInwXb0aGGS7tUN5SdMc1lGSCSvhgHrtnFbzkHShYApdaDlWxFHTE
xIDZRzC/MkTY3ZZur0aUHwZ4cse6RAUO8grQUWr8qxK4NkRW7Wv9o9kblMNfl+sV
hQ/ICAra3uks+7V7/pc1LkjywET+ey7U9EiLqg4sZxYVGcDQER76MRl2ry0YHhUF
aE5JI85wyb27H8gyWZMzA8YGkJ21c5Bazv/JstCzEOI2tndAN5URrhQ1e8EPclxP
oaGWIORt6Xo5lSh1xGzw+ZP31h9BUU4GdcAn4+ZDWAZK2lQfABCb6QZ0NnhdMsx2
1tB8YNK0UwFcedSirDdOeDpIkCqDpJ9lqoT93NWt/GeOAdKlpSXVfQuhps6S5DzK
wNzPECejaDlUJvnoyF6B9b7qaGkpmdP41XcdmtMoE40fkXrpln3jrdYzi3mQMGBp
9f3gpry94NdSv8MqbRokLSZ0ZuDDkEk7HLxxmEvM1IH4QsHySSi4/KNeNv1qzDOT
mAW1qAIQAMhDZT8K1QQ8MIA/u4Azc96kC98RFkASUHADCs39YFGwqV+aWZUhASWA
3a9rg/MO6/yXiTn3hmzH5KYQFGnG54jXLnKmfFF9I09hzK8y9oT3ZC1vHc/vLwms
Ad3QndyQ/nBUblETcq8iE3J84axbZB188+Hims6TqtLy+qqmELTaSPRbUGrFsKLV
BpUpWv+tlpTqNOO+yEg+Tj4L4npBWSNAli/YeYRQskq28RKtmGEMWp5+VW/CL6bV
1dUiFa6iEvNugJcM2GgOes/2Ff9XNDzz+qkLQ6THdu8sd253jb+4/Yh0FKtppUQi
xLa9/LhyFcpokJPhXEeX9JYfMW75ikw09OgPNccu930GBvY1VzCCkve8+xuSOQa4
kc8GRsVkiALRpMmya5Sm2DzpvZ7c/1Vek8GhP0+80oi5DEUdJ2LLcKPI5A7RVRbP
Jwd24wr99Qx+mStu0K6K4mXkHCHLo5dzUpgZ7tbu+I7yI2AEzr4BlyRUyjVoD7q8
bkr/QNvkBvk69yPq/+YcRPJT5v7jq0V0WtnEIm/PYPtI4nEdGa8unFGTs4XpbTbY
Lzf9z4t+radvSJec+rUjlanMTL+swA4jmV9XT9A72C7mIvxryWvXfidWLQ8yrueu
VhMhkNC4VwSsofhVnAIEOICkBfHmxGar3+wpA4lX74kpfmpsvdfuIth7MT2y6Xj+
sQy3STPhbmemzxoHwz3U/aOkCQX3JIoHplCcHy9j4tovjJFLebLvLxnOqvKSyVEF
g79CPUlnxH+jc5LE7VEd5JcO2PibT2b3wcqB8fKR66Yv9BRIdEXFqa/f/xP+f/zb
iKdg96GsqfIVOvaxVqNtb4F5ows3I43gM75+OU33YPflNtGO4Ty6bcEYKSx7+wrC
1S83xcEw5yU3FZ9jcvenvBEhswUy1/hV3dHPaHY/n81W9AW2aSl54N/IGK58VAtR
uHYD4O2rNo/wM1l3JcSWIIZ0Uj+RTXW/qm7Y8y0BDsAFXlgjrsF6U0kmH1b4c2Y3
n+wuYzYUWP78Uu0CX49PVCoWiKyt7CL/NjHBAtVwcLXgQqMLjVT0S9coltYKHamM
R+2oTY613QVWG+oBrjlDL0IYjWaqN2UxFJg0f0ighVc2ikcQharqVobPb3+6lkpx
giuSpGZKnegWcD23c5uNorTbNcqPXbB4jMPHiDukxCVc5CILsUUaezXIrldwgdqi
gi8EbDuW6elkOLM9hCmbbE3PLOBnbh9aSqVAuWmtqLBABeiofMsxoeC0tUqCzQ9h
XCeJ0bppXZ7mr8FVBZ5gFYn4Bi8Qt/+V1x8SD+givf16qYD+kdYfsMn+sGIAy1WG
ZMLUeFOENZSNxU3MYfjrpjIAJ3w/9pBXO7lj1I1+UFQCnUDit/ymrG4YMZbON/QQ
Ct/dAHoyGTWmIQx6suzXP5Z6R1Szzw6a+mCODaDg919SRlhVsU0LcPbBJnq4PsB0
i8Q3N13RGmEka/w1t3IWA9azVeqLthocH+clLO8FhWW9PEwZT85NJri7KCmn2vBt
Vd26vmYfWW4PkVYXKsYt9Ot2Vxdu/3Av3u/Xthe1bRHvrPyqXVzV2ilmUg3AqCo5
kvphf0+QoYtjV76dFcqG2rFCWqZvgUyGVMS+mqBAarp2E+L24CZj+KHLHmZwDs4C
7aCdlTHeYBDVa6m2Kp9lVAeKRVZtbGiYHC/iPdkbabmMOt0KjvoGBhAOy/TOuzCn
qkpIY1BYgNvSXcRoMeVdUnDcMulTRpxuobHf0pLmKFpn9RKcS1FYvLmjI1g1Xekn
SLe494Qs0i4uUCAgIJjf1BmpvynXgCf7uOgjkKommf2WL4zF2bRSgjNf6hTVaJOG
NaUPOUMdQUFxTcH9Np4g26VYG3n+8eLH6GVXn8EOr6ADkVovQj5tSesyUqGVKMGL
1IDnwsIGR3haKXd5gs9GGYKSSadVfcmbcbWVdi0VqkHFCelGb6X9TntUuwdwRPYk
ojOAjTCht7rBQv7n3r4Y5rICspSYA/48ejxfnCQpwfJdALE3WkQb96UugynE3dkB
7DRlO8oq+few6A5V5zZYOHuDVJ+mmc+ZPVVdwYMhHpIlBh9sO3VfpUupyobV0FA7
fSCxTUDu/VQlQ28su9f1y2d2p3j86ckqIF87nACeg/cwQB0USDuUhRN5P5VJfDeO
urxgkACUxby5p9sHbRsxE2KRAM/sXPPK5230NxcpccpHP37xzZ1h+yddrpsBd7Vw
byHhhATplhmc9yeifao7kMhMohLIixvkQxeztGw5qaJ62QGgGF6sAD7uwq6rGbeC
7ukCB+Qt+iCSF+Hsh3VSHNBDgR+zIhflDLqXJa/Ilu6H7YLnWuyrHYCRUbPLDrd4
HH6o6RTzPu28v/91u9C3gFB1txp9Yr6gpIMj1VWbZ/Ee13YPLhLRzZc/+8V/7pfz
JJClHwn1vbZW0uN3WfmRzaJF8t8FXEr27V0ldUsOnfzMazrE59GpHY/lTcHoIMkE
/N+kpyLkegtixu2ZFLe1KvzQzg1jIVQ5K8xbIRaJ/OZTHauPqjjPGS00r5MX6les
gdAdhM09yy3v7EhQsOfeHCs+56gMBgCukZSvgpobIK5HpRfYkZea23KAi6NFUUF1
J/gA65oC+q647MbxeFrFaRM3cOXCK+O9w9cEOGGLMSD9Om+qojdO44okf2fvWHN8
Hvhf3bo+yXSrayWeqGe/eSmfZBDPwq0f6tKXPK5XOPU1LuTm66lT9EEnKT9weLJD
2i8jYyX25mQBcCJZ6X1Ww0gn0xfOEl9n1i+uY/UDcmQnkaD0K+/6flzzCVpZK6os
JYFyWsb8dDsm9dOvyD8RkyLKX56sIW/k17WmCnJtjxZt8XyNsI7VlxYvrGzWnDzY
5qdBBYwxWdLnxkcMtUlcZIK43kIPkfmZUgeYOUq+JZ6JRqAhJl2Rm/DWQAZgKbGv
WkgV3wu2TByfHJ7WXaGQ0T75JpF/Tiv0s8x5UW5X0i3JL47OTImcux0F6qa+ny3n
lvLUlEhrQY8g5TANumQnZKJ16QhSUagR1H3WVnI3iO3A5yI7+cUdbDITywja7ITe
J+G9z4dZCcl00I/FGuEVvdWKOgrtE8XL9R9KA7lFy96cQIpjt75eKNBLfv+qPKhJ
tETqq6NQvsOcLaQLvPqEyExG4lYyG1TYYdZQp6YkuAjQeOkujRCFzI2iPQaNtqzt
h0j4sTcV2R+s0imHFedRb2UxSHEg3iENdBei2xA3BjDbpYLWJZDi20IPu6HBAoc1
P+tzDVMjPH0KMmNT5yjUzOcI66Psr7lmOywLEqXdQduaUiW1+VwZzSEXss7CxrSx
2y4MsrhUFuPVpo5ZBDWeQrFiGJWe1TyyFiG5hHKQ2/4F6LbXnvO6eGCQAKbWfR1C
HzJ4k+whG3rF9xyfKLTucHc0MnOq+rMJB9G/ngW1TwgRzGRkwGlU4tjWKKFFDhMb
kmlUt2cd8HExk2PuM0h8a9ZcqJN8AAZUWgfyCH3Xw6YkUqTWyWjxHGZC9EWSKSQy
u265fQFaSX+FOML9hb+MU0fEfRMg9hvnZoCjAdyCA1hUQaV/3R40RR/54lcyJQLG
EOcz4ms9gWTRP6SjQ9EFMOuUn8QIakbRmOv6CdFlyufZymRwiM1B4viCLnpdeGMs
+U9Ers1MNPj3SPl+O8bx6S7GSghW69nV8EBLXy8c4ocJAwXoqjwZ/XbsEjmSTl2w
xDI7rEUV43dagZ7AztEl5iJtpdHC0/+j0nSKmOtacSeXgMwQAYtjB9h2p39pwpUF
PkjseoIFLhhSIS8hnyMYgyhAJJhZ0FYGZ78z7H7PEUfOeM5prDrgyQ0EZRl+gng0
jebQ1yJWTH80ub+AyjyIWEqtWt+Ed0vOkKjH41HPi7pZUtX1kmnXI91pZcs7BA1M
Ov+3Xuf3eqxDt5oXZdu9ybaRz/TrRVo+JcmKELr4X/bv9xYmc7qVsfsRlflOxZ1y
cY455nNfCrKv9vbksYxf0K0eYPCHh13fj8OwzjkztkCfbPojCmtqSjeoVGL9CXcZ
ITR1HwgYSTAUxL0jDlVeLJu/teHSbgeFNIyftNYG907BrsCpX9/8cop2GugBcjcv
cfbhyua2P+yWG8VX5IR+XrbFBNNd9Q/ksUJL2a1FMn06YMVtnO5cI7Px1qyy97dD
yYeoImHa8v7rhi0FO69laBcczS7ItiLUAd7BNQyKvBwqtpcx+XWSLMblRLU8UGhf
z2+YMrax8ABYRd3NdS/COl81gfEFp6oaZtLxxSPEl6I+NTX+BPdNhJjYLlHXhGXZ
KyYV2YVu73PWz/uvk49o18Zr8vH0HLyGQ1ANA4Ud27to2kMeMboPEANah2W4ytIb
CrCBoD6MTUC/gFk5GM2+X6BD+swZ47p945rQQj3sxYJaGotffBRNCorwdykKbz9/
YSHt7EiKljo2HcN2DbQ4x+b7+kmX/FmCklFAj86TSH3rlbDVS8dOV/ycoUuNcNa6
+Kj0XyleRXeR+hG7311XESJo7yBFE2CzjK+G6+z3MNMZe3wX+GEJKfSx8h/6p/Aw
ruNeXLWQsT2RDFU0+mBbbZT0cL1QQLLjFwfWnt8wyrS8fIz77HXpCyud5v0ozK6n
ZgCilig0PcuuUJ8qlRRO0eCoBrBFzbl4kmK8+n7njmnyJEcWGAYErZq1gd3ekr2F
01SSnsjViHbm/0uCf+KDH3bfLUpF9kWkTlESP781niecJojj9PgNQlBx67aqy3Af
O6lcZRetoGc/NE17738klL2x0peM7bd1ITvgvmvQntzuzoG2dGYJhAuqelBt9eqR
ptYawnGy0/W10LNeHR6TMXn2ID5GwH8Ox5qP63SL8JtAzV4g20JKGP4WZa05ccpQ
1UWqHjA/rOCN0ayWGw7kOhfCFhbCwT8QduyKyNsp78xg+oShp8MzWnX4nTyVsSHI
XPHCvWFjHGuAV67qDQZJA1lPrlxSAZ2fEb81O0E63yliuGtiPsaZDCY0OFsvDKPA
pyEwVbjO8BHDJ7U54tEw/L0tktaDR9x+/ZUVJI2OP7YKvIVrB/fYiCdNxx7zLFfK
jzAzx5y708pgh6w4iIQapaB68bwSkj2MUgyRqttLHAyJkG2B9YELc3zl+P2SVISv
ufx4BESB+2LtF2zDAAmoqpx2330WcLnI/gcYEsRaaoejLX+D9hqqz59XxyPVNBtD
IJZW8nr4XErqO4z1hcuGYnjsKrKnThxgHOwNs6UZc5Fe5/zGeF2LM1/SzbXBQVTB
ao8Aaso/+g0r3f9QqEPcpZpqB0fqi/t8PpIX/tR2ARqFHNqB204RYy8tag9h1oWS
hdW08xSO1MkmrA5c2hTmdHaWpKHZWy2RfS01WpJcpCbxaku5px6sB8515YiIJlsL
9Zy/RlVnG4l+66LPBv2IXb18jK5WF7hUgoBL+ZmqkWCJkg9bf5v+MnQEWKKTPlTP
qwu6Wtcm4nkfqdk4ohBhQNljAQrt97yLfhzvrXWo9sBKQoU7bKU8uakfoMEgDl80
HOcKgGl3aGAZVgvuXwKcC74nltHRCcf7Qh0Ab2AdSc7MCnfCDxFzWlFwT/e1AfXW
358dVTV6x3AalyOvMKGOlw+zPEuIFaVHXmERDL1gjww1QrU2Rk+Ucamdee9zPxcS
2lLHLy6GTLjyIkyKSjFw7mOLTKV0geFxV49mbXMjjIs0nq6El7OX3apyQ0XTbUOk
yBVmSdzvnXmGgbELwCzLzbwK8JjwmKC4FM68PfaCP1nXn5BvG1X64E0bAGpwuFxO
BbZqVqnY6btF5zBvTypOYkd+o+OH3vdKFjv0mTIJaskcRamgkapFr+sBC3E4PGmL
mtdxiga7fFY5D7XYPKgycRlIyZPH5sQ6ZCWgKjTosRhra9q/gikD3CPrO2ZaeIRd
wG4ekVuSubYCZfeu9gUluEsJYHyzDrJj7to2fOOlzpIYB7YDRtoxWBJBpYLcAqg2
RXBeEhhU/E8i8sfhDnQdSx+KfdMEodJ2TKwLQADhdIQQJr//cNWh9cs+dzCONF/k
JQjgwgtPY4rQO6Kk0KH9iU9Pk6kEF6+JLoTa0SdS44sTaFcleBJQH4VjM1Tvxm5q
8yPPSsLUcARZFLcFuCWmy2OZmFxv3Of42QX4+HaPmZU/iWr4zGwmzyU2QaA1BcT7
YVqoZVtkmJFGvlZQuPgj73QFN/pFjzyPC2MA/BNhxpdcxTZUlBhEdhvJX8jq7HyB
6ibAQZVE9/Z0nVSAPJmq5DXhuVfLMu5xH3l6uZG5iFX3V9Lp4vUfEhWySYfIKDr2
snWJGE7OrU2El/yBwEsnYezPkwT30HsnHUUgBGbK6LbbJNSnjttix3Y6Oc4NfuoU
mZvx6UkDUQ65W4MMCTJW/dyTHZ3lGIZdQtAztFmNO2CJNPifyn/v8L93kbp/JO/F
bgMW/j7Xk9+uG/e2ZgL1hu1FthtMVNNkWpg3bcRn3jig5PlTmv06gFadfLe1CZ0M
porJGn+mW5ShH7JuNiJDnudYCfajGau1MHLZ2HZ81FLwLdOMA6genlrs1pbhPEIb
ogGR5IZrhCL6547GwolbhZfAeeAwhXIIMNoWmw+zEBcoQZQB5aOIppwTRN7hPClP
r75dtvIAiM0xCwymTQtA8EFs/UwFPiRHoK9cmtrsmvQwGi+UYSC5dvuKNGzvLCnA
gfOMtHc8kYlEnrysrc+BaoIdOO4K7Yny/kXJHlnmA9Iuo2k8d+8u8hL+bdpgP+FN
lZQR2dcFD0237pskwDBCbCBqGgUKkLWezX3b44rAIRl25i7Gd1TPPFXYRFkLCMbn
1NJwrTPME1ZxPMdigsdNZ3POZF+bmpo6PqI+NmOPMlpWS2AC83vlf7XEINhBnvbU
TBy5+p4zLe8sHTBtxzIEOddOYiRr8b06IoE7jYRLBmRJyNnyxSSPi13KFRovCWc2
TtKpZGl0jQ2Q9ic3OMBNwEkD+qtXJjTXZoJU4yNcrNciX+mGR/R6JUoMHCEvizjd
fOsJpBQpzbjpjVtVymOt+IBqXRRq059wvIGU2v8lbEpwBn5CQkO7d61H/iaX2+m9
pOteTPikgTvFWKPMg2sqkKzAXz9Y64frVZK22UJ4DnoqsCB4GScfqDSHaUEovIkd
BpPKhiQ4KrcHbd4GuEeoYAl2pcylN8Rh0un7kimQradHuBsoahPnOed0bvn3gBMx
dF43230sBCdo9+qLcYivv7Yul1XYSd+WeCXRSrEs5z3DISdSlPoiGKctfNj+Prup
BK7sY9jnlk4V5w1PKCMA1xyAumCqqG78ilF9KFxUMcyzQIErF8Poc9XYn2m0hHBl
qG4M2alK8lJ1Pa8jDQz+kRJVIdQfbw4XTtI4VyPjGFqQ4EGvEzppI14VAdPT+ImO
TvVvdQ4BHrL3g7RuW/8PhqtqEhaDwoCGjl+0lz9gbnZMOH2a1iddXE10AVg3jj6d
4/S6NjGJgo0Kh4qxuK2x6k2oo0bRvz6NJrDSYAlfWJ4ykAgJ62+ZOc1Z6XCpNW4l
dsan0frPAKS2rbPrTBE6NQsgzfKI+jBBob1DZjKtLcLRM+sv/HkYfLMgjJyXmPtp
K64lPK+5NMUFwzYBRJhvmzsr1gjsI8vHHDkHnvwNBp7KCt0jc0SdaSLq+uPyPf5a
pzAtHK09GIBXEkKB6G1wpFoo4eVbYGs5yZZrmw4ueM4G8VLBL7grUj8z6p7zR67v
anuLvtVKjlWKNwbksVyf/sOgduvZA3fr8TYoz0IcJ+q7qT1hHgSbWwZokUrCq3pG
/QJJd3oaIBdUsyrefHLC+TnHzp0Ju8+LKXYCAbmNmx8UCNYeygkvsWOq0tLrI0eh
RyTtyWPDpM728L1z/jLQxPn9QOKJ1CJm38uXmsf7T/a08QUDFQfLV+qAyKesdpMK
F2a0HskIYqSXXsDSUVw8u88YiJwipESk0f11V+EvFiAZToczuTv/bg8WsSsIAbCl
V3EcNbjNL/mmoUQkTMauqoFq6ldUaZA3uZh4F8UG27INybCdEAbGD0DjeEzCVo8c
Z9hKSciSbk983uBlvxOXYlzhIk+7zlxQ2cf/gSQC+UhRJ7V0AhPp70cihCaaZlWh
3sXjgNzyswazRXOmOs623ZjEnni+RrGmfP/wkx80PvXkKgyfL/rLzwFd9YavcncH
NUe/HN8UQRsK+qxY3Rfd+mLu7j8nIn35g9MVPPsAa9zmH2/Ktb1mpIzkYBWmPKph
h/BUr26e2Pg44e6oGPATfLaPIRrsteOcJrGOHdQOGkfwSTknY6t+iCIME1/IS1xO
Kmv5o/r/9SsMpi3vOyknnh9/4LMXRiV+rX8g7TBuz9x/8ep4JuD4pLBe0tljEoLI
wMWDOZeziSNev7V4sInwB8TgMKVQtoGIh8E4OlKXwhgU/ZZFMJx8scmefHuWbAkB
U0syatjtpXnbxrbQZwO5LMTpRqILqDOiRxYOwUJzrHv+R2HIZ/xNaDnGTIpiLimK
yzhnfJvkjCUkVSMZCQ9LKLFz7PJJYy/ABxsgFNjCyhsNlWp4Q4qCk+EY4TBG/EjF
H5+vK6FGkK4P6xZFW8hE0uo38As4ze8ALdrk1tui0YqdBnYSODNEZUbjtRbxCs1Z
w4+sf3k8KUjlW/QK4IFnKbWtPFndT09xGRCQKmXcPHLlogXQcY52WjwxRN/3Z3Og
S6kePhs3ypUbhjzzqADH7HJUE1C5CGX8njSaCP7n8dLVMxIYATE1fvmHSjfWkedz
lp9/ugL2BhA30242wZFcdMmjlz2I4Zynmw8WpDkzm6XFHv3cyavgF3i7aiwWc3KA
i/adCcjJn7M2e5piAl/2bNulftgu2Bm4WsI5kBqE5tEFl2GRbfeyx/caVVerfUdW
4eZPRd2S+N9hi4eQ8n/4jXPlnaDq7bv05eZ3XEuooEUHWh1aQTOUyPwCGhql2z6p
mWbFeS09PHatAueUuxc6BQ+tVCSANgfUiSSdPDLvhTv3qeFZzvJSeiiJ8/7JcVku
6C1t5avSs7xH9c0YWErqo4wS7NnJO1lk5Mpwj44T8rbqDgWrO6Xb9GdgKRL/TD7x
Y+yCE5Stq+Dx23dcaAYumYHR25qDzoPfEZ/sh76TkzEUFNdXakjUJPBZDjn43ymm
ANDKA8BOr7Wh1N3p8x4SHsl1JNltwsmb/SCdpWlJdSS5qengPnf6/P00RxVdb2r4
m0E3QnbKb6t9i+ASpQP44SRCz7WAVjk+ltnLjFCbNnt6zsZYTrB0chAUnw2yOMXr
GBrCIzGBuUf631NNQJn30Zhad/oU0YHV1OBnjJNdZvVyB7rcp+XsHWTkAGWBQnqh
eR9aVkp2cCgrDe28JpHh33K9aOs93ZiWrSIjoT58Y16uPvDjkS1U3mwZlmYwvzdd
CzJOIafD13yIPbKVbLrSKfVgaR5+rP+puR1QnVIKrL2fV0br/D2484fPHVyr6XTP
Qp7sFKaZBuvdOlup/B31UAn1glYR0BBVmUVxSs+u3Xbfs9r+mVV3HWdWGwpPQd8b
AOm/CgBMCVHcYgDNqEQOZTaiRzmLy6B1xkMwKAOc+U7eahOXZzkZpHW+cd0IspH9
73QP/oScnxtp7rHuzGxQBQkC20bP6k7fpVns7c+/12uMY0eThO5qASIOMvzIq5MT
3CfWsZtWVEbnGGeVsP/InfgSYricd4enCvYSCG6EwLWmxZijJDadLAXwIs9ASHUM
TLrbSw6I64EWN7sPtXIwb3knXVjVorS9EVPn0kLI5qPZeU1sa5LcqF+lGyYwzkSQ
RtvF0quVNiAtj/0Kyh9+4+aM9Cfl/flmNCcwXeKDXBbnt3Fj7Bz7DUUUvPyEedVi
mG2M7rfzC8EAPuSNEuSJ2DakujbFIDeSyATKWsd8l3tO1p6p3X4jvq9EWvY/btgh
PhR0aWM1ljPdS+FuUB/u4FB2DMlSgfv4RMkPDnp3hud/53lhE0F16oy4AZPHz//u
47e2syP+J/v+FLhHWc19uun55RK9e1QP5ZRBok7EkKObWA310q81WRJHbGf6qufe
NjoGjZi46UT/qCWH1ELNVs0a/aGIdPNveBGOXx7BBUbA39Sp5dT6pbltb31EcylO
fsfa/4RhaQawj/a38rw8f19TRB8af84Xvm77065rsn+Eg3mUPOSI41ziiWe67vsd
8O9dHwDTMKn4I+nV1wqjLHNpa9GLPN3VzqlBTV+FBN3Dzma3K983Mt/T7+UHsGxT
FEe7evEsXxVONrPjtjTxb0b2RwQTBIChCk+bcyul0LlSFT++6/R8VMsgAxHG83+J
JWREXuJN+TGQ9u4NpmGUOBl8jkmCrMr1PTXhK2FC6wESL+t0ZCUYRxzPo8LhSl3n
eJPWb4/oWvjekRNT78Klv0cIE2K5djSMhInBbPGLEKXW4+R2mnfwogd0KnmGLl4F
26mBGJZNqBvL3QWWkNefsbth4EpqW6zUAd8ePI9M+UPsRdXQgpfwOSkNiiBIXF1h
dK9lW0l2b2/J9i05hdatxb74V6LrJj6C9nLNM2FZN5z9rL+C55xxwP47klGwtmFR
Nk7NZOLSVKe70UQi90nbY7r2Jps6UfQMXzYA+HZe9eIKs5Ap5JpLJFcpFpalSmft
cpjnqGmSPdUolsBIJNUjNoBec54YJqMEooldzI3PyrHONqR5H6eT4b5zK4csMMLg
u7tRiPS92wUN2jHrk/lG7gMvWpa0VttZ+VNwQ81sMeDRqqLnIJxgrT5WEf1i7MHO
j+FKrYKg1I0FDBII5fVJyq14HQ8tOZu6tMBsjlprlKU7R/xN5N5BRmDCgaOlf4E+
4Jtk4yY/v9S3YfHBIrIQrs4CHdPnMy8ezeenUMzQhJTWJ+RAHF2K6MfGBt4G8x9i
uXmBbBVoLo9+eke8rxfdJ1rCWmZ9uePzZ4x5P5hnvSuc7ALHfVSebny7bMzu2kqh
Nq/d+yJ7Ssb4FPs6JDvBMmC4qjZgqcH7pLjAZ4DBWVIPBqdMrlvobC/gESw6a4Nr
C4UpBehYzDJWbZ55fPf3YA+phsKcPskYE7Q9+jZCh+EALbU/ZAaxeZrehlC+HfRd
husiiCE+VUXn7cLYUEe9W9OMKpJ68sDBH/7FgQTZD6RucZC+O7imzkTW0a4ivELb
6BB3HCWoJiaKZHxHl/VRdlm4wav7NtfHFxO6ZXgWKBzYrNqhI7uoVxjx4rWsJ2In
O7gTTrkBUk7tcPnEP8avi68hYoijqrEU6Dyxq5hX5AI3Xt5PYFz4gj8ntymz9wDn
E/ZRoqsFOSM0LNYm0nu4Gxw8ZbTq/wAOG4YCzAtURhGcreWKrgTuyn/e+0ojI5rt
9LUbpYrtNEKkE3TRgBdfV31cqJGsGTBGOpZRhHnHgQaMKrkGCo7zinu1Igca+Hzn
1Vz+u46t7SDdh2ibTZ3NLN009SqsIdZCM9YSQAbdGx31WkRAnrqp0EMdIPGIdo4z
429GAp6cIvkzAn9qgHldJSNA6RVtema+SSoAn/HCvs0E5aOgsGwbFPWhPAYlC54M
sytQCmfdDL+tTEBSZH3KFXhK2l/DCJAoHNUatMHLHV8UagT1rWno882p6GkdgIID
qJocjqLzoI2Ba/blzC4wpyY904B4PyztUkXbkChr+lzn1HmCeYA0dMsIfQ20bInd
C5cjcAYM7goDhu1HLSqqfGZWt/abugEppeUWlJPbNEM8YVdG6QT6v9zsLS5dFcRJ
G/319PwanUCMgd+Urj5PefKWd4Qww+I4a+ot9vOg411hBrPYVaTWHyZ3FuPWMQp6
ZvTqLVLx2QgOmZI1ywUUa96Cm67FWSpy2yZdH9Ck2NpOcDpUJ8eLRTuymGwWl4hC
U1vZCiIyZGcUOPUtzlqS2VOODyUvhXTagPUSrNkfbL0q9gSHSFWTe+Hw+uk2j4Q2
kfsZQfR4kBF+bQdjOiolLGaAmjxUL7EyJNAzUE7U3rqzFV0BB30Cf6/NcjChU1f9
uJUg5PNuyX/LD5+Gg8IGbeQ22N2eqN/3uMNaRjFlCTdr0oIKZYs3gkb/5CXMCPLa
/FTee1FwIs9asdXXMNo5KBy6YQvnQgIwIo8siRf+mn0CDxzXV6nTKX6qgRUfweJF
dlJ0d4dUwBcAupaH/Bf1HxwIOcjiN+8rWVvShwtJJZqJGHcJdhaFoLP41ZS3QWt3
0di9BeoKMTH3zmBO8By4v3sO4lqHv+qLUiLeTmV5SbSV2tPI5KNVZTyMBcHjeblw
4by52aP9DFg+QVkGogc7qUSZpuKwf15ksQf0QniX6KlLtjGe/1cWbRCokcJct78V
ZNRaT3Ay6whqgdTKD8JC1qCeyDhazniJ7UO/k+sHPFyxOw6yI4/pg39avUlQ/mTK
U801E1KfDhxG+NaCBAQwR5499TYQF89EbJasnfmZqIEujA/hyhfngJH80zm/oEsl
RQGcGWVvyNus3GOBFF6uI8ShqrY5suUcTEvElJ4vPmri7EyaL4Yt9M65mB/lWWuP
6XjMeN1twPwXa/04PYyONc4ZdNa8oO5lTkj3Go2EhWBPYZzhc2W8c1jd2uUuthSB
1lsrIunAcfCu4F8C9KqWiMHXxeMviezsReRnHLLnT8rHWJQbU+wdheVMuoEMSXSl
tcq+a6r+hV41XFQqYKqka/sDGrr5MSMU8sidE2gFXBwPIttFGARVlKKWYNlNQhZ7
kr+B/8reiB1/aQwhjZwlBG3U3np/02TLPmWQhVgR8i9aU5x1tk+6hC22FBY93tHg
eio0NzhpL7O1EwdN/IYcJCq/1jhWFQYa/nYsuZXslOIfc9suqLkCBNYJzJJzfJ1G
53D2yh3lh2rkfFORnZmsTjs8mHrUCYg7NWN1rIkjkykF1qpphKLArfVvFKSX6k0J
R/qATiE4DEMkZ2utZv/xBVu1BSnDwLTcgYpntFgPgp7vYzAk+9pIfcB67Mqexpxo
6Z+cimIyrFWjVikqcNZ65X1DQNLkBsrYdBkCqB7Z2c/7qj6XsLiUhESZBzyKF4t9
aWE3lvMx2Cu0XG05skVD9GxMWbcquCsPq+lwqNoegqYR2jwUEd8rCJo5VsbkH+B6
xwsmUQWViR425NjhproRrFG4pw/owomXZAo8HdZblr8rL+KvUQ6LtNXynAB9+/cs
rE1MZmVRZ8KcuBORKBGTGwJ5cNwRv1ZITC2PcLMoGG1UamyPNQfThcF8pGBuRRa4
zkNXYnVMYxXqYp8w6k5IioLKTCbYlSgllbCqau3GIuH9z/i9OzDxPNM9PE8Uk6iz
4ACU92f6G1K+k0MFDgLK6oSqUeCd+u3Gkqvgt5eirVv2Oe0zInMozhlkEZkcq1it
91cLnyVY0WgMfy5KHDz6G5ayapMdPo6cby4BorVzoHxqScTbyN45UnsaD2avkIkQ
bFjrmUHE/azFpgELLujDpfBO6Fmxj7qq/+vygq3T12YUnIVDTjhfl5CQYCJ/ZKnc
Wu3qGP1BxjhCQV/v1u6i1/3JN7mpK9BtCqrjXJOuFLNapyF1xzt2zwEjBHta+a5D
gnKgF/XGcy8JReS26o6ss0tFpEv9t7qGVP81hP8rmPzo0k1Bh9UlK4AX3kDlAiKl
eSMj+wTrqiPIBqK3PsHeWfcctR3zG9VyTESam9B9RtCv/xI0hB84DhqkDpPWVDmG
JfB4fe+3kmwsDeZTGlSDitzRVyw4LFiY6L67BoXve08oKvylIBMgK4PYQPD4kAsF
ZwuP3n75EB6dqSPi/zzwxNHb4uDrlt04RS0hfAGYdGfvj19ZjRgxMc7lAzpK/b1d
2Q6oQec21xTUI8X70paiLTKuh9l5q5mUFu5H4rY/QipsjzmZ23RStrqWfDCwJ0Ds
fdJ89VJEETBr3RwHqmLT9yRmHEWGtkZzgMSB9SvPgkZraZHXdaFBeQ720gp3HI76
4M/5v4rhH7DSUTPGA/thZG54mCaxJWAj2WbaRLcysjmn3Mlc78sKIDruZUCT5CF/
tC3/QQsUVJEU+bVvf4AVGEGJz5hjtxWYBbwkHLhBaMVJ5q+ppBj7k4ancZXW6x6N
WrYH/QYkNNl6fl4dHNhqncrjvAxeYV2QF/j2/RshpHcBOXgI8Lj9NfDDRH6Iu8rC
q7KHoiJik1yURq+uqnUs2QwRnFif/z00UYOtQe66wmywBYY6KuNKlFjdfkpic0UU
BXQxsz2WiGOyOgrdA5J88mC9A+pWIQTJpzMYoQwRVXkbIK+N+JeLFScU2izHvJcu
nlKHdtd2s3wINGXPQJiJz4x6tV4z4uHkH2ZmI/x8pm86nwqo16+pc3y40UItFTF0
0NmU0kcVjwnjdKKfX6banU8lradA1z0lmNcIsLo52P7Ty2L/edQuh3XCx8Do5vlE
0gZXLMETfpbYrXRNz+9FyS8qfazo3oboSpXfUq9TYGhOlKcmr+mKlHjbXIIz4PuA
NaJTaswgxhPez0XeyH/ikki+b7rGwG1hSTxah43PFpF/PtWbCOdSua57l5aRyApq
p/8WyTIY6Sq2IdA1Z8h7+NM/oqfZJdoCy+SGK0lbBxscrzwRVfyCsRHcuV3LpNNv
642Y/cPO6I/gIcqXtUBF1geLdUgUVjMj0hCm/HeeWXyrRqyMswYlN/+/6hdWf8bV
8m/xi6jYzWUqvuFgryuw/+SytploXnwlmTBRW2yg11TnipjjydXSqkZvnOgkDQGq
MiJH92Mm1U3y1a8OD2VejG8FvjaM//IVx8uPZTNA+BAAHVDQp0E/5WTOGoqy2DvV
9VqonJJUNn1bYKMm6CY8LTZDo4G6O7/mYI10/d4NqgxQodfyyqJFnXTM5gYDbcak
bs3ChcqDiwZn99YSj//GOb2up6fGswiK/7YcsTWvRHauL/tt5wEVW5izU20nH53Y
EzU0H53A4EStDwR2Bam9OYkiRnzCcGC8SQR7IzrBUXYeIMmeFUk4sNAgIgN0Sh6k
HgL40IlIBglsYyw8LZy7FWlkXTme/pKIqBvW0o25KqllhrUpO4nBGM5ncvyRxDuu
c4dgiMLgEovGG6uaG99fUAr835V5ZQ6Tflr8oLNb+X+YZ5G/VDpkGmV4+utwFl5F
/RPuqqQA5xSpW2OwderviDQPdINMSYZQYpgovGQr8XJSfGZmMvl5sli4vjm3aRgi
+ag2pLiQdCavvCXV7v4oldJdz7UidVwTelSE1dgt0d/EexIbb3WCS1WpJC4L0Vt5
XtJPchLSGggX25StXtadOxIy9lzdLDbp4fqV4xk5M/9qd8ZNjxCvQF9eQDWPjS5I
vJqIFgewjZSJmhq6RNW4+TifTnlfkM0lLsxuQ8AqSY5AmDAOUBtro3ZF9BKLdVQj
ktHTWrJb2ZLr2plweqZoFQJPN91z8tO+eJJMnkLGxx7gg4FChx21vkCRlmoqC9cy
1kBTABBMr97TuFsRfKOiHxz8PsPcjnXHKUrk3dW2h2n+3dcC2LLAH5LSe/gqboET
4Xbi8cntSrRanT/UI0B5rM6Ac7EsQRygmv0hisqsz5GHYDOc5ye4FbIFAI7Rd0NE
zGdtHRaDqAiSQ3m0G8z9F81AqKDzeyjqV1liJuHSOl/kPkJp+Nul8ZzD6OI/n/hw
c1gkzuH+d2Vk3ecnN5512E69HmcoPf2W9U82iOyplx/dpslXi04FnNO5hM1GV/fu
qKEzT9omYgsNY8Z91JGEL8ZHcvmJiht8pxLmFYqsK5EePOxI7gqXWVm3BgJrJoA7
F3ro3u1TrPxBbgcVsXqKTSTn97zuAp/DLvs6KW3V2tQuvyUfCORMsJ3Z6bMmRi4m
0qQI2gQ/yMVVaApJULQvrnrptGANQYYD5IVFFw+dYO3CCtkLFfntDVu3pfGSpCcH
lR2dnTpoJG4D87posmoAEfeZvQKn+1nFR2va665pNtNu/tpOewt55Lal33mUnK/y
UXbxDeSOJG2VKdE7wssTbEPze7n9feviu+dzI+qqL8N4Q/iWBfnhx8FBbYtEKK1Q
wG7mPEFywuRPApblJMQ54ZJVs4VsqRE2h2VLAAxWFP0c32eztu/mNv63ymluBQG3
tzxusqncMKx9rTh3gs9kvMT6MW7A1NvgYtDhxKqAmw/5Goak9Uhv4RTQjm6AozD9
6iQuAhDLkr9M2L8VTIlhdiwwmlpsO0tC7p/16DSXihacUvtWisBnzuVBfn/ZwcV2
2lHAAsIm7Gjho4bPw5ujwmHt8fan43Rfxz6Q35whG9QYUoHgfImPJQ+kzCooF+AT
fF6tLc/zzzTE1hBBbTZ6k16t/tCoP6gDukEUt9Fn7SUv5adb5A3WOWe0Obfl9g2u
iDOogILBCtEB8pz+OZTsFHogwY/EkfI1HIVDR4tS5rhQkRF5iWBkqclVA8tb/jES
t+oTVeHgHTMQT2N8lj+quGjY61jh8VbexeZSqo4fu7i8Yx+bz8cuhnqoF3ZwA3Og
ozsGMrh4VbJ/nTg5t2sLX0EBYiavKY2GAzlc7Q5MOIJTWLtgFJgTo9BkBPckeDVu
v/b+E/1kwfm4gHQliHiepNusq4SkBL3PW02PS9ow47AbSeWhfxDwMwjLB+J23icU
m2xSnvf05ogNmPnXnItCtJFBPUTkoKt+X3sKDPPn7vBsZ31M1g7snOhKMCwmJ83x
eWSPp+0ffGtWPH2OBINFGue3BRhyvjm9/AUuq03N8ncaqcIUUHBjSQ7SXzWyE169
j6HrfqSx8Dp0WISlUCAJ2MMpqNkxbA3CR7xNU4NiI1dIUCW1yrbYav1HRU/1uGj8
ABJNrjle6Jj3tB6oXUCPuUoaAhdBAGAUlEYRAXnPRhwktWVhDdanz+5VOsEZd5dd
1BdZWETbXjqygKRSAEikkm+AX8aKHcUr+J74b00eJ3PEXV/yhq55+Umw2uOJcKd7
MOC+PknygLxboOZCEFfSmbOs1G0ijyuXse6E997rnByKLxN6S2DvBPgLAfMq9R7g
VG8mWtTbjL1L6PEc5YqkFJKo1/+QzWu4IClRgTua48n96xrMqdyYpmC9q326kRYM
5NO5+pHpvTaJRgVXgIsDe9NiAS6/HLIg+9kGAjqIT3FZlhwZhUhyw28qIk1yCJKB
kdFoKqiqInvN4gFzhs3Ro6BwJujAuhzRux9vvOxpjkEwejPDahltmQ99MVZZcjML
mPNZtQp5a5z8ipcM9Jr8FX0P77dnPQEc0h4kzm6R784Umpz4h0KFYGQWifCOT4b5
sVxe9i1VDRETsZK3tNRt/AlWjusRzHP6iT0un6BoTNvc1mcuMbQj7YjTGEKFgTjv
RWB40dfGvVHkVphPDtPiYNEzE62a0wbQ1dzp156hXverBbW9N/coHrGwvSQjoQNp
cTJTdmvGxw1qMESUCFCFx1jLwLkrNngm4103y3ka11HOHpM7FngoTtg8koLu81o1
SCDWCunpVTHbF/RCsj68lg0lPf8YofAj17G5QbXD1bPeoMnH6bg1GyZa2tp4MpGT
2RPZ58zAM+c0FAQ5iMaMtxfGz6ewd0bEn5nRnZ9CJKI3sr0pAzebUDf5/E2srdnt
tMU058TBjN/jvtVApw8AsF7DY/qg6jTdydawLUf49xlWB/ViFbkJsE2ZP7+Ab2Vf
IQ/AfcgebXaa7qfeIxziP6AL8u5jT8DRe8W+M7gBOoKYMsufjlHyeCUD8yQ/PFcW
RnFfUjTcn9e5kJ4Q4DZ8SY7+8bVEjdAvFlPKZ23wYbjFxOGsYUxvlFy+n5Si2jA1
EulYOsGxVD7oDAZYVkdeLYvqHCw42UnO66EkrtZF3If2IVDI/YhX5+WioW8njIjD
lCukwTbqFSg0RSGBU+5yiJRjaWbYQsPywbL3JeMfmuMj2cmfZ6IvRntJovRi6qS/
wI4e+qc5IoVLPC5LQZRHQqLh60OlVXNpNI+/SVcqIh0QxKaeC3CC/JDGesh5HhBX
gT/8WWEWb2vpgcubA5VcTQ5e30qtDq2upyQ1T7NAK5f9JeXCyC9I/O20szw6ChQw
v3rgp4ab+QlNh2aE2ym1Im6216ZvUh3dLcnokVYuavYaepgM5KPR/cGXHEwuOKqN
+OLGoq6gn3ttNwsQW77dwljY4mBGveGX/tSB/eE2ea1iFNPomk7y7p2ZzUlD7p+i
qn94SrUjLBiVPIKlM1F8jBtYCsV4AGVya2nSvAJOpxOwPZ3uZcRtyhAgooRhaFqi
fyCHNo3HVCQW+kd2TJ+TlOsGyT1cQrgFzYCzqs8+q2n4yb27Lhc4gu6qmUatEX9f
RH/M5gPNTHI2nzvi71Za+Pvf3A4wvbT2ABoSi1+th5bcsiLUbxm6hDTF0I6VIeET
6aH6uf4Q46YrDFlOOp2swE5E4elxzDuerELcZ0S8j1dd60w2DZrQFUw4bLBNO4hO
tkJzcyNhsg/VyCQRX5+QR3JSm569HHhiNafgGkeg86BTU8van59Mc3vlVoudWoEl
iexmiQg7yfPeNfOeaBaGXz89jIJlXNp/ZwXfiAxB+B6YwbyBJhuukbLplwcimGSX
tar9x1pyDcQ3knOfHn4gxsNrb54kYI+DYY245Bh0aqDQplB0zXQep2W3MRyPD3SD
xX90OIJ6nw2rUE4EQ9J2n/5XxwJISO5SlXwLBe4MPK5x03VVpilCTu4lkvDJYM18
dxz4SBtJRvJohFOX/Nk9gSGAVuXY8Nj41qjOskqK7v1fw2asWUatDGTK10UWEHhe
jz57oY0PrtN7ZV54NOVC0IdOPftByILngQmskNeqolQ+ItaBFQ1PfH8JMD0URPKW
hB8E9oksd7M/Wk/hMIMbcMli0Jf5egxwtig9k8nzXY5RoDtrUli9Y4/PXkok/rGm
iZSqZNu2xC3wCV0g7sdN+e9t0DMdXgm0JO/5ec5KXfVeFkY8xM3z+2IRcKk0ir+r
lb9joqrGW1yRMi0buQDgn+R9+klYNcXIK3uqIbcwr0MNwMwNLBY3ejqxZQdQo4tw
2e6fTaNi66GZ1sYT3hYfyyZsvqUicOQWL2Wx5BVLVhfIy7xeLgnn/ad8nrPevgMZ
nLQJMCTz+MF8godItWbayK3oPfHxL/Hec7jj4R5bOqx+JlXG0X7n5s+zUchiI6+j
mGoFujIJoK1bYeuLZ8RRkVO0TbgGxqyB2DQ7+oncNJvZa3y4Y03hGNBw6sJOG7fz
TuYvK/9VTVUFhJcKOsrd2pxaRH2NHvfqv6HvNgn/E3/jivAu9C30LCtD2nctTxqO
bOLrdqezRjxyZlRn8ZCxSbcGgn5rMMQNqeQ+SGdxjQm5AaceZJAGJFqZHfT5CIzs
yqxrSI7XFHD+JijdhhoFuH3ip/SkYVCt9wAiFJwUHiB11yVLM4wSMNNDzpgznjMB
WC1sv0vNqROKHf8AF69TahzTOOYmyFNwCE+wnT6oY8llhmZchp1ttjbc4S5Mp29W
LQQDD2/ScEBwbWJH5YAqOrzhopPMWkyfhI5jNA1+QEYXYpBrtkBNvfrIt+/G35rq
Y66my7kLOp+aVE/Vo08Rc5UIMYvSgkexzItbwDCEcnB/enJpFSSzbXdGvunT7FSz
AZYJ2NjNDQ6UAxqbISGvhxD6v3R2cYb69lmWhzq+/kDpkPRUOOsJFS6hbAeK6Y6C
1wYQfEyBBvQrLQe9PIRkG+Xi0VMeahS4qErVYYIhLqu2mO8kUrkQhnvjYDK+doIp
WpH4Ca76M8nF31oL72yyibodCYzMx9SfP3c/ZcHIpviVOxGpll3oSEGp/aDKu2ej
RJQ9KdIEP2JmAjfWwU2fHAAUeVHMC5IWgLasP2yKnPBHbsWO9WXtfFLH+EB5/L3O
GdlMq8mI1ZmvYyZ6yMNmavWr1qFrrCVJ9hCGoZzPjv9GjyHKkSOvxErV99P6Jhgq
Ttzk26v9Z5npCNDxNgMhP0oRMkThPFoj/60MtI0gL84iNoaY07xypvTtADjuSawj
kDAHPxzFDDX9Ne3MoNpMU2pPRjgDV7kJmvSuunRRPcDntZODxszCQCAkzA6tHfRo
p+paXmKrisAbmr11b3BygI7PNPSdnJJihwb2aVq54e/BmsrJkKmhvGkVtxRYJn9J
6zuguor6MuHsayoIp5Jk1ffWuUmEdGHkWKPVvu6aji5nDMaJ8vqG8CkbOr5DssJj
Fxs0fJzZYbWZ0P686uetDz5tKnDJhq/Cna9YZb3TK49wJ804WIeJxQ7eUABrWAgy
D1MP2eVTmKbHO1V4fbnOGLeLfhvvNCSoK9lKLtuz+0+9MnpVVCPSLsY1TRcGvPCD
GZiWe6MckSdPpI+mr+RokseaG5Qp1mRQkrNVKrJPtUwtLg05Q4dvVVPYwMgm1Gup
FXaMQ82NlQhdS19G7HILnB7UInVSlrOudgywe/kTUfA4Y56xKtLHkCJDhvUz5lW0
Q3EAmuI7BKuAz7kOONSQ1K70YWtJ1bLrkGRLYBq2l2NtccgKHSIw7Wep4A70BSr7
upkfb31sgbyvtvTxjs3HkOikpnY3iAVoFpJR/miHsNS/ERmsiKiZdsJ5YBwo8haR
sQ5Gy1RHx9EvKKZ5ojqDsaX2/i0htDRHpNZX69Bux7dopVrvzP160IsWu6B5Xo2x
5mFu4iNm2gk/2NopMwfvDOsjhi9jpGz12t4UBuYcRtj3l3iE0eVUFflwVZyZTpsj
ClzZZQT242NUiBVUDe3nGL0wVQwoaCKACd5jDvGirBKGUsUYJdGFY0NO8rZwRFo1
euBDRwbNMoMS2aAx7+lcJ0tbyChacNEhLgoMYwaa1c1Yo0rnl8y/eNLTCLwNMuB/
QpF8rVN6e2EGqDslGR2jEDW6FQlUCOBaXn840JH5r4iLWbNoYE/wTCHcwEnqLbVX
RVRKF3O/rZ4cDhuCS15yvqwTTxGltFyBiFXcWzq41sq/RFSWSXexrncv27VeKYfx
cl/0k0IUn/MgINMihrV4C/vyJwTI2079jleX4/34hB2X3L77lJMu95VhJ6hDHITJ
2q0/t5j3AMkbCx8FemGymCCBXShi8Pm2nraoFlllwNCqIsaVQorQUBPFv6bW9vLQ
5WHJNl720a7+GQAOcBt3wknsr3B0BuZlhb3I0Vrt46sGLZsgeL6v+OAYQ49CP5SI
EMamB2mquhKjAcItt5hvJZbpEiGmVSopJnVjYB3wUIr5+T1kf7EOfHcWeusI6fTA
RCyk0a1jMNV4d1ZRAfzTM9uyKmHQBCCCbPkHreAxDArQGOpQZngJGSCrMQoXy0H7
KPo7Prq7v6WZC21gaxyvrIFwCc7xwRhcu4pabiz8XDavO2L23c2uA4z28fpqC65B
4AZlk8CJyXmEZs/lfQbehNicgaTJzFYf5jqoU4f8k332aN8lGkoPy1A9zns2llcu
qaULvUheIP8iuVDkJO4iQ4YYWi6ZXQLuiRAmpoIR1B/lywDmLjLajzs2ezy+eXD+
Xo3SHKSZMh2PwNNvs0WB9uMzIqqNiuLJJbiGBUaplOdRue24iRFX4EOiiyEgiTuF
73kp6h4DEk0bSdlrYN65IRqV/1yriD8H/I36haXbkIN0f20YBXFbjEis73z03Vjh
AHRM+HjK7b0cTgf/gjS81+M1EjxB5uBT2oo07YzX7CQXoNB4HQG20cSqTUrPbwvV
jisckLtWcz+LPakzBRuj6W7vVjehI/+fjSthZRgAyBkBStKNBXEULhbANB3810St
4FWiiSFRQhYX6EAL5MM7ollAgonaoyFdaT0FzkmtmWKVsCzin9cWatHJC5BSiOZE
+P+g43cquOBHB1L3S63h18CRbvNMioD6k7CluwxXVhEhyTXShapZ3tQrU8Lne/mr
woQ9o/SDh1Df/Vqe/X/1oC4gGp2cfWtbh9e1cDtZ+AZGGE9nmmNX4w6VTiODPpUF
AEJDrqwJtmFD27IpsQTlQsOLSNAOMYKyduhfWc/PmkAZAHUstEKXqicWcCUq+wgQ
e8EMg6VURyPpl4kr8CdVpxJrF5vCbcqEUM3N7ogoXoEPkrG8R+1b6y6R8CI05w4u
+OdO0NsRmywqXXEqMe+4KDFVw3F6p5ku69HQAgboF5Z7gjBEnGHY9nxqHmAEuEpU
LfAXBWohpIL7NKBMOffpQuU/KpXwRN2Q6I4mfzQXgoEGhLns7aD+3wijJMCig7wy
5rmN+LhH2lvgHAQY4h+gaGKSt+ahwB0zR2zp9L0eT+PpJ7NZOyamPFCz1X0sS92F
An1I3gDjozD9ZDotl0BBr/hnAEcOJ9LP3jU/2Cx6VVeD0XuUjmEfv83a0Ykb0Uhl
PG+qGuByjZF73RVDYI2+n+7dQ2TZcu5Y/gdBIax1/zbjX9hEKP0x2SHOGUyQf6+w
OLkPQm8TaL0Pp2mdJP30pF/jLsCCN98ug4K2A2B/TETpEvUV7/CxyI4zvsRnJDkJ
0bXmnWLqrFB6hA6/BNWICh236ctXtAuCZwagxRvFtYF6S/7cKttLm1EM1YrIRk5j
mBUMGmd/ncXgkmXQ9nWo/1RRPpbkWCoxBUwdicFnsfKH0lgjbzNrF4LWjkV5sjxd
eGL+P6Ee2EIrPdPONyV4u5FMz5KJlZSJ8WghHeijYw8IOH2Auz2KeWNv/8C6RI99
OBxttHOtniuCFKYgOS3++RLB7yezN8vr3/2SprMxuw5SHAOGxwo8cqiKtOyptbTC
374RIQ94QbLF3LS3UySp4u2n3BYHWAnE0MsLZgtT3lFxAI4KwhVew8EzKSfr5MKa
9YAxtfL6e8JtVO5EROt33XK0TNM0fqBt0rmyFLCcCypp+fZYuWI5XmLn3qcAXr8n
rTc4aYTci1GNmqZ4H9SI7U8F2wSTfaacChx4U7SAX7UYiNMWYkh6kmjVNWNvins0
a4+DpuOEorkz2FY3PVCUcynYHO+QOgqBHAZHfbI11owPsOvDj9WTFwqLet+lI+un
7Lsi4C6GL1tAM20QZApfmnABvMWKBzyJufSZUgpz0nlqN54XpH87ih8thwrpC0oY
XVYZNF7mFd3xodpLdDGOMp6IU2RS+CPt3n8rMgLhDZHhBPfAMfb6nUdxbZUuFCx/
d7F5BUhS2FhQ89lwvRY9ZTyQjDCDR/wUZSJ9HL/2QVgbteucRT4WDAZ8/HpN1Ttu
yocM7KLLNPgf+IEQfo9ReBwjawpl5BIqsxFe+6nBsJ9JrDeR0uQBT2LVBMl1Ks6t
+RKc7/CF21MwoHoIlyUmpPoi43z0o6BNAcsQ1TFAimPHBiBd0zpFU4tcUPDmfrHV
r1kiHYZtFeuxwXypv+lf3ADkrYnHj4BIr1ngmSh8/2ilBYqNBYk3RSZboVYbL7ls
O/mOkILCa0GsdVbI4RFb5WEPdigH0XXKVAxlu4UP8JHxUcGmHTmyTwkTSqf6zMwu
qz+SZO1txM8Wqzqpolxkgb4qnvJZyDTvAM0lOUMWlvaB5hrDHsXB5PLZnbdf55fj
W1DB/tNEllJ2JfrNQouO2OfhucYQWfVCpOvBff10sKdChHzYmDV1BtcGWdxaqO49
MU4JUwTf/rG5gWFEO+3Rw19kK4jZsF31JOaxfjqmctr7jtFPfBjOnLaVUZ7d7MoM
aomILrNCen1Qa4Q/lkzJ+VrXtv79A8DL8B8DlNhL/pml+eySjwhAYfmZ/5TvUgzy
6tbDclozoxH+k/FfsJAjo8+I2rcdAQ9VfoNxA+ksYci7hrtxLO8HtxAhfU1CGau1
9hPY2q8XgXAZk98B1edl6ClUAh+Z8WvzwWC7146fJ8pIiXP+wlAAylzsPSLzSOg5
XD2qbphsmAt20SdOtnA1o6x8gayEj6cSziA218gre0t+kRuLwMc9dIHF8SXAIXWP
QgB/Zad90+Nq1T2Cyo4FmLbmra4K56MTmwYeiOtCQaVs4Wk/6b5SaY+KkUCwa79o
Wjx9WJ/LPpmslUFlGYPgOPHkk1zOLtDX89aENDQPmhWRjJslV5uo3KPXPzJGJvzw
LSZj3NP+1ObxuQ6fpHXuIwRtVYTsEQLeGRfp+1rqRgDptQf9w00o8EocNpe+ayUq
Dt26h66RoVj4tiEo9w/PoM7McdH1nTW10U2TX+wWP6+bpD9z6HJ56H1WK6u+jnJK
eNdQVzsWW9LurDPE5EhffMXC6oHUYG+BKvrJUZdRljuGXLLcE9ExBCWdIR+moZJ7
WoZsQ864GzE6ynr6PzI/I1yfefyVyfQu7aW09XHAiIgje6jEJX29eh3UhA8iSZoK
U96Wj8ThDiLpcb9CnVNv0IQ1soMPp9LOEtTqWVk4X453b5PIMZWmWVp3AZMvFB/L
wtd00gXme/oGmNhATbC7CUmSqDPw8l8kCktMog44NApcf6iJnaJp1/T923XBKpXI
Z7FNIa6KyuzdRhQqbk0ouryAAyzX29HW4oyJf9jTgkIRywv3ctZ+mZEryTC2nhAU
OVWxCM5imqX6OWl6dxE6yx9MQMSFG5AS09e9GLaPQm3IKtDPu60t/TmLExHOKOM4
5nU41oEXVi4LOr2sn24nR76/2VemqtI9IHVq7vNWwre0hq3aNyYPygJ6aGYY5KSn
U1mdImIOXeJKT9UrBuChSI37wNmGdC/d4KuS2FqRjkZgoFeQ1aJfD4tjQK4oRccH
2zU4LfAdkz9ASiTi3xbZ/uEUmxCCfUBrB+alJkr3LfzawJnzVuXzvkU1AIQAKHeL
1Awjij5da636tVTZXOMTPSjxZS2t240JbVx5Z9+wRNfTeXnAqIUs1Il+VuKxybPS
Kga+LYbyNI9rQHqu7epQaZi2insXnBe4vGpTGLI8Sz/OwWz/IRFhP1+InyNcAtm6
q+PKRyrDd1GSFnidGo51oUf9qw9NaqChdHrNeJvOYWpcRRu0BXzD8+cefzDxG/AY
f/9nE2CYyPnbDEsENyV4UNj3oVPDE6g44PE8fvQRHJefEKY92NQNgG3GCbM6v2Pq
n4Y8R/+XqtrnwQVsogA9C+cgfrAYM/noSm7DD8qciC0FgBZOAvVJ/vHguk9IZDyi
fvhM0W7OoVLMGPJk9qtvB8CLGIrCN3qyCPR8/6jswR6JO6+8Zk6/YgpkqQwiFfYk
Zyl+XVUdfX349Hqw7wvrpF4/uwEnPR8ufpjb+5g68BicfmuDN6GfpJOltil5pu38
RUxzEu2iw8qKn2dwWotWkf97tVoviVO9XufcoBfEuSejlcvCJByWJZCGHtVhKi1o
XNh+t3rOQ1SZ7aFd3V3b3YbKLZlEIjMFLenG7/4p2gAhHiDDAPfQlmWkk18VO0Ls
2woLRnp0PXMOmuDwSOmZ8NDWr6hZmKdOFw4yYmpfCzC/YAWzSH6JkU+6+YpAoXUv
brt4ifR7PQSsF6qHlAYZbQ57Sgnuqpqk1KEq6tjFJFSKc3/UUanfJ4/kGGt+AbEN
7kHnI2k2CL7vBE9PMYj9EoxpmFpqKlHsugAm3IwQMqWGJVzOP/9ZAWlMwu/uxaW7
/GK8M1aah1OG3gmr5gFaw4GM3OXlcaE6cuJZK+184Pqn/frB3RKwqWL4ioUQU6aA
y2P9ZmNLR8onWcVkGhux9wTKWQcYB6O5UT/cX+fMzmN4D38vc9U+elcuHUL8L0fn
jAovjojg/6LnfJDfFH9BVkuhq4D9+VKKoaS3JnaV3QgXKZ2uBpUYOLaXJjfZeagq
5ahM9f3z5rt5dOTQ4FoJ2wHrRs9feYJAaBb5/RFC+UZWE61yoYJ0ugsvR1eKG2Wi
Udg1FSbbmyEXQk3AHr8C/ed9h9HxqTqPem9oPwwKfDqHoN/03nlX9PpzaSSQpJWg
xYs0MHYRU8LzHNS+Tzbfxjb09cZuMhXZt7wsGz2ZCJm8ApHseAPtzXZMEmJznmfx
yYniCTQ4OSpSWgVfOrmNdDx2px82ASUXigrgdKsNi6aqo81Ps8mnzRRb4ccojB0C
wXh5seySwCJfmUTtXFK5hQlz+Sl0PdG6HWELN+Dzkd4EAzqGVmGprgZdTuw11YGi
jkwA8oGaNOXSizRx+/iVSqGsZv29DlLbq2viaPp+WI5fwscbxoBax+suy6t4IasQ
rI7JnsWx/GHjji8D0VITHQiUDtpyyZnppXFy6me0cHzwE3vDhJSWJlC4jpH+CbYV
SFBByUCI4hykIHs9W2tUe0fDJbAWZO+pu9UrtWEu3WBbmpcakPWfJTlP3LAT7qov
O6i7u5nA0CocV7d7mdxjbArX7FPvhNEZu2wmtEeMjDVakE6asdO6e0ooA16TUkdP
KUDS/eOqQwXcNL0hI5AuXHuF/jc7PJt02On7kgRXu61UzsEMbZprNxlWEalxxgxg
hM1/WWGgvQQxOmex7H/VAZJ/gnZ450PXlNH/Z6Hn6pny2WrMW7pZNqKH0n5fodbi
qF0EbQ8DCQb2HIc3PPpGzMYddchtgEFUVcNCmMkcr0bp+cgMI8zi1QhM2cZTmlnr
tR0DOYqqRXvuoFhfQ67/qfN+SaxSrz8AEF69KsciZl1KC4yUfSELkcB1ajlOksnp
FdG319sy0nTwotH56pK0zivFnAscX2tlo1Qiycq3I0YrX8eAa0CQN8+NvOIY3Qe8
0MsMLJ6wDKpRYwu4r2TzA+l40/5P4YEOR9v2lWETI07+m5JOYHes2X1FTTawow2c
vyfsztKRntnXY0ZmOM6jRsy9uKJB5GjyIiNbJyyB4FxVWa7q/DCdSFkkFa3KS9h1
mIy5vtHbil8kqMR7ps5LURFDq7FziaRdQSwjsYGiKNHFoTQLvAJFebePBs0kV6ex
yJMKgcvtSELsJTEJAKan8fcDDdJhbEbPVmN1RQ++6ksNzHTMFAF/wvp74IJR5fjy
CJ5BpgRdP/dcawk/fHwyXe8Gl6Ln3ZOFO5xVdQZLLCeM6m4N53maPbQbV3KsulAa
svEThIpf3y6Pzx61DheIvWyVaH2fjWA/myMzjX+afrPmkWaIbnj0pXn6I6nVgGWF
L/JuSnyLU/O+6kOCJMjTAOZlEpr2mvctKjVE4CVz03KyivO5q8DW3jMEDVGuczy9
YbM19yBZt5X6p4JQ/5X/R35BBb4nvC9z8+kdzSkajwZ+9aDJuYek0gZ4gHu0OLvl
7mEj4AfbqazkxT51qoIyJGd4HGFJt5rsMtDpEUw/JURIV/5lSdYr7kiMoYD+Uzci
VJLystrDBgNPo7i+YswBl0CnZS2hcc+SQRboJm5eXMslHhAJajBnqB0nMvJ1UJZo
C3foTAjUqVIoYIrrikgOAHmpdSqn8O+N6VvXb2Q8sRE5UC9lLJQ54GFbWmD1n/yh
O9sH7h09pnqt53HWraWBt09IqrKFu5OrFVRTdi8Fcg8ikfLEzC48igYl6zNo0A2G
nLKGFtXAjUmiP+TgEb5PcD2clZeJD8gnywIJSjsafU1E/U/sva4T+fxr2Fcw5lgi
tYHZpRyA6F5cdEQmJOEWfliLhJBwLKOtcRzTlxv9SUJFD0u8n4HtiIvyR6i2g1mF
Xa4hrQo9Ji3T2vPF6b3BuIibv8wthDrZptIaPKUmvOCV5bY/Yd/vvD+0tEcnZK2H
7abZnk61A6S5UN60vnwstzBEN7JfYuz2SYRXzMZ4rAiKfMQGFxMwQWuu4RNQwTDG
ypeFciXRTv7SR9AwViVaC7jPIod1LTp1eC5AFP1XnioW8uTN5EBIoVZ80/KNKlvV
j5uF5oWTxC8ljZNUuLwm4Q9Rf7bObMPMt1L96rmVMyB9K1BACo+LonjULj7xHSa9
IcqM8J8jZCsK7RSQB4mIau20WpHV1dvSaic71ZTX5cvmR6xFl8/MU3a6R39aXNC2
/Wm8FDKD9Mq4r6L+gXAkqFEqxBoGwIyrtXwSAxcTZe3bS/T2aJDrQpZuiEa2lD3D
BWIDlEyMU8xF7wIzYLn/ft+WIU2EXpjvWcXoD34QmB2v6R9ZmNv5U4cqeFUqlXtP
Qhhpg1Fms1Ygj1/su8ty82mNDeFzN5on7KtmqmPNaohZcCX2ABJKcRF76Lv/5I7p
r1gMsTNIrabVhi0ylm2g6ZiEJMktvXHmG+5nEMlDBwUVs27NxbPfU7jMBZoB6aLB
OkE+7UJuOrVaA0nP35r1BoREUsD5aqJjPDQSGO/Kfi0aUrGohY0zwLdS6OrNrfBg
7kOgS6x5FvI51AZP/+HWiU+NTJg7JzNbmwN/HHg4jVtwEpaJxU16Ueo8+HOS3XtK
ovtj7eaTJz/7m5lPww1W197q/4me5IrF5WOjjUySlmtG564qHCcayFHBr6O/Bwqk
X6Tw8ybg8BvbI+SKnf+HmDmZJ7gZYQ8ELRTkqTP3qQqHjCasye6YZlEjJesViNIH
ZMYp8gBPVRuJhX2pdP//fhCWOb300t2MguBuHeU2FjkitnMOQvkvrtAd4WoFPu83
0j6AN/HJt36BCA6Dj3jNUVTX6dmG30StQ5JwmmaYmo3weQPLpzckCUx3OzBB433z
iboSBzmU1po5McahbB52qAhJO+tpgP+LLXc7BbnQ3MkOVjGt8RyrG7ngdHStA2wB
BfL60U5fLVtbYQMyirGXYXAQHxHNNimH16M/QiymLzo3P7K4zQufEy0RSrOCBWvV
OUQYVPRnkMRjMGK15xSBMJ3HZNB1zhkeZhSHJIOVJH0obuLA9F0WXnF0o3+tA1wy
Xk9aPUpbUelflwA6k5liZO49wjh71sR7kaqNCAdeTV49wwXfCkFdI8MapIdKmaCY
1irWAQu7tLNXsaQgY1bP4KNwNGDYEelKnkacBqEk0480yAWDVWkBat5hwex13GLc
p6pZeIXsLdOLMKFhFRBNnP9Mmp+ribzIYle4+CZA+kgMY1GvzcZlatgg299YTcgl
xtZSr/H0KFpTTpkA2153731li4mudkKDV8wPi2MnK2RX96SUX/B9oJZKbW13NNWi
8fVlhXHH2PO3A6xA5hMCvsiB0y4BCUfKHHchZ9A+adAh0acC4dRGurNZsTG4oeWV
k3NnO/ofvr+wcrWPYo2D23KJAKJFcNLDLHSOv9Bf52PhJ7lmATIm5ytUSjPjb6rp
tlWnoKSeP701kNPBsSl16nYVsGkqbOQNMuClm8aJDEgmPf82OHhisyTU0JQjpAT3
thMdZdwMymVObRmcyjjb9+b1YCSDxKnJV7Zs8Zo8ib3qr1T3/ijZ1RhoyYTpln2B
ery7IVFCzVcSQCD+w4JcR12LgDYrpvc3UqyGcp6MkRQXxfKLCCFVjHSd4CrKcIdI
GbpI+b8CKj1IKaJ/1PKy6bIVRi2RtPn/LhadvXFj7XAcnaxYIR/aQNP8yMysxx5V
KA1CPngelUFxz7VSBr3SFOqKUsi+zVpQPkKEYdey7TXWf2LweM8BqounDFSAW/rN
/OztD9IIUJ+KkneGt3koq2p17KYxhx3eY/gATDa4rFV3TGDsh1OZDuud2cljSfB1
pXrfTVI1k7Xf/oYdD+pxAb/4qMqUCmWtOm9R8g4x5bF0kK6xD8+4nu4toW7cA5F8
e4TnzNsKmp3dab/ZtH+IqOd1ssgpz6bHWfpVR6A3I7xp8/toVNZ31hsQ3BC7uufJ
dK1+M/emIoJ6GIRSb0gSFFCdCA/8bYfomo6IKSaYdbScUfO6VJyTkCyxtQZxV349
EwDpM7913edYkQFfSQE5aq2uFRNZK6kTqF+Bu6vVdly5xcLp4pIuw45/8vfRlC86
1s7mak7uq1qaU+IGmvHN6Q4D5QArgxoLIEAwru93v+froTmZ7GoH4G2GTJfpKrN5
IukfVB8pk6afUuAiNSV8V/p/ipBOMLJBTr8sBjY6/uPX2kMlBZHaSEfa21CuV5j7
9Teb0eqBGOMQaPDAwCwD+kL5u0nc/gFyUo8es9xUgvA4FF/3XlCVuTZ8l0/YqeRa
KBrCLvHE2iMkjqPCuDu3utjjlKHkVov8Zob/C74Egp7yBkBgyIsTXi/ziuHdkwM1
QGzFluGowhKrrl7nYY5I2Oam23kg3/bKBzu/0pHikOVH0fB+jZWbXIyXuBxi8Eh5
QIDnwNHtqyuU2HalJTcynUj8YJxNYNzFCw49Jhdv6qEqoNfLBmU+9D3iIL/71kM4
kvLfvOYaO8TY+DTJhTVOknEhjqEioHPlXEmTtKCHW9eHf02avryiA1wRtrChHeRi
7F++IGQZOK59kCrtH6aOkm0bhTxo/XMwLOaf/r1VTwYQirGDcF78SGMdVloKDcCM
2mMS3f77inH+3MhU4/+EI0gVI5TU8xK+fOxw/a9ML/GOViktx52qOypraWVAPf92
Xxue1A7PALdLeX2rLDczaHRLIFk5ki9WFVH8ClfuLMJl5jGvow6D/4KOgO3go+eU
xNhLL2+0u1wYMNtGprJTrjKSvY/hfeJJ06mjF4UuB6zhXi6RtR+CUbL1nuYmX+Tp
nqxfo5LaVQGaXn2EH0/9iP2i+DY3rNIlG0FpNcYjKavqZWJ6Qx+YgZAYuneJv7mE
7gUN4OHgFLShPrDDf4slEG5Jsl7wozKm1w5hkOew39fiIKkz/TVwNbFSS03DXNtA
dBChQsr5UpwEPUMEz6u7AShNIEYqywBBmNY/rzynFLecM96Soep99KtJlNgrq1bf
bNTNAvuqlwkAbUU/lb+EBHfWr1Z9OqUaSJxAf49jjbqRf1oD10uZz/swFWQ5gr6v
hXkDoVgn14CbD2AsTYdpd99z9QVMnc8rudjq1R04ZIElYcYddK3YAp3WHUEbNwX9
f7PgbPufg9ivFIvAbAeWFljqF1JeUDN7P8H1OK48o4vMSwpPT2dhgCsjjyXRXgkD
m8My+/1MgHqd/i/nIdiescdRPNeNtO4nb7fuHkYso5Mspzkzgpul3w72A74TiY5e
wO1Hrh4mlZJA/v/pl/MwgtV6z9dorxhjd18GWaTUv6BeruOv2jzxdpVKx4Svm5oB
zE4wYzWODA3JlxAv+rN+zXEkPgNyzF7SrGCVmlELDnb+oF9FvpP74MKpeO8nLRMu
O6EXRnYRX/BTIMXvKZgsLdHm3TDvc/7ptB+7ymbRQboXuVm5blCp7QWczspIJzQs
tdNEWURuig0mZkf/su3uWgQLO/xA7ZXex3xFbfJcp0QEraYpoAIJAaPwCYnY3lmB
LuMcGXWWi8nFpIdo2z6HwIAxsHvbFyF/WHDyXKLLN+erufCS6LCNh7zPEweJNUtj
3TGvw1dq3FBtR2H7zO3GGw8qyK3zoMGb5QKA6K9fSy/dmfOJXxH8FgNN+olXVCVZ
pjxbw3p2HcI8E1i23UbweUOi18DgGmCvNyuSqNewbNy0JbU8u9BjSbMYBfIbMAg7
aj/9c0eu5UEk4GsfHIXa/+hj+K7xlO3gPTRXUSYFXox4MkrRDCrQMiGHSh8xy7s0
9OhVmt5y5J0bab3wXL4FW8GhLyupX3lm8nTgB7A29L0xTK5+SNA8elhaEi3fM1Ik
YJ8Ey2ha0zgEwmfomElu1XytZzawOrkmBeCRgjT2iyP/6+6oH9guU+rsl/RLmWEv
KCB6y22g1XEtfN+MYTX66vWGhAHPMgWNpcJ4TW2tMrDaVsFhjhDsDseI8STuOkEk
k80GFke4TKDFAFdyg68+3pY2PTSouX4IEsXrNSpq05ILK7xqGupClVOqUAgtDiAv
SxEzVKttv7C7B1jST8msnGP8w3a4S4RZQyuO/n1+WWncPVZAgSyb+JLqlVYme+fg
gchhSkLosLzzZnx2BkL5eAhlQWJcEQRuMpgZOsxP9c2ttPNMnDbig3TZu/kKU3x8
9Xws1V56qwkY9ekmMj+K2TTssOX3MD/aS0Ul8dmdaGvp6tZiyf/zZ/U+sEAvpmNy
XX3NLMbTOmAyECgxRRGFNWbpxTbYR5DeMuTzqbupmzF/5Jij/omqZYJ6ob0arCg0
dXPYuuZQS4UiCfirxsEK7PR3Eq7uVhCbU4ElvhL7DCWOE8Fs2IW1gaslfgxuqERD
uuDRAPlVsoE0Y69ZaCYQ2ttHBgXMez/uj7LCS1zfR4sYteFiqMDTmhvxGymfDP2y
GS12cO6vJWxiDX71GdUZkRQQ2vXowrzGAijmVixARqO+3LBJgeX0gHTRdsZpti+0
1EvtWLx4co/2/PQufdvdFgCDJMxgMIwC3JxQOtV0bMAKkGoenacZeXIEVNE50PTn
kzNjNqtKIs00Ko0i67W9p7wTfwFLu87MqxL60Fij8JS+rfJPWJTtX/9TuJZ82Yhz
zTyUnIcSdr/16jEu4fDXIJB0DyC3HZ2kkplTSsbLQTY9w+aAIjWbVXlEX5KnyB+e
q62+32BmCc2N9stExuycC8PN5Rc0ePJdvRTqljDyvbwglXBNQYnOEo6TTAaZ76CU
OTt8o2cBlAUlAS0SZ/zPxcYSdsOJqgwScArcPFObgl6BrSnRsAp8phzD+v0mb4Va
umVcJ/L8Hqs4VYOHxLygOXSXI61x+F8TQxN8mktZKnyPuAL3Xi+Pz9Vn6bNJzg9o
vMnP6IqfOePcu8K+ZsP+7uXYSafPS8aEMUon4UwGV8tqbYtC9f0QM1Ky95PhBHBB
GZ5A7wW4U1cnWlr8fz+zwqZxTZM99AmVBhzXC1TKG+KG7gbobdUJ4gY1zlnG2ck7
Um4PeTetdyk1Jly1+zDnY2Kjv6HPxBooKTa/pUymTzD5JbdNevW/aZ6gl88f2WOZ
m8k90RN7ZdDT4o92l16xjkhwyckz+fQ499N/Z08dKQ1Nxb5BHlMzaE95aY1XXPer
i2HaUrwIk6O5WQMTb1BgrwmKXi9z4DPgPXwMP9/CREdtyUOThkeuREDm2NEQmiGa
zMzJQE+7O1+a9nMSApOaXZ/qzxEtfxoQpZIXAQEvN40yYz/A6KBT0QNu9OxbQzjb
ctgXn6nE0yzPboyBBFZ1lPK6huFF4k08PtWZEnYxJE9Kck5T/GW0jLs/7LgIOhrh
Ix4ypjUCnk+FAnpqAomQ38tz2KVQX5fL8pqrDuGxMmsqYiGHzqz5I5gg8NXFr/Rd
eBVR6Toz3BkHo9CYoK7bI9nbn2pE/4bScgxaA1X9RVA2Bed5YN8Jp/Tcu7wFgr5c
DBsE+EJQHo1HwJdrZC92vr8ZuuoiUjO4x8dkB9rRD1TYOcGZeK5tJV0UPNUu802U
EZm0HAQLlAdqXCEyAkADLI7OkLhwfSvn30F05Ta2GgpDwJP/eeielOeNTwKWD2q/
qTSGcdbsfTqOLxGxChW7hjEElVHJudA1V3LyRso0gWDUm8ZJsF0EmNqjBTZo5uDb
ttJ6HEyaAWLVuKxk//Lds84ayrz44Xr1dfSGDP80qdfR0ujZKsfR5Ah3VPZNUOZe
XQjCtu7AlPKa/6VvVk+c9ElFVy2hb9j6ESLiq6oJ4U2ZzK9qF7BZUo9WyjX8Mml0
iSG+FILPLkd0O8qs2mnm+e35vfQIjYKYeeXvV9hncypsTKhTG+ITioDGyLDvRz6i
Wsxz65TNs2r3wCrsDOZ82nlGnnQ4V7MQyrN+8Hzg6v8RPdDGZ03NsgmJm7alPISH
/Ecyqx7fpHChPuli6IJ4L5MomoQ3fHOH+dxWJSZUNeUnEkHEalkhanlj8J/GlMkE
Gzb6bUsHwRdMRh3It9bB1fXKg8j3lSLCBhjpfvrAWLrl/BM1krnquGHKwmo9C/dc
hr69kNfEd+zECwOeZquwtdNLovf3cbPPKMVudATMH50YQTio31JZiiM0arPgHHTb
nNYSwqy5b4C7hjwfNKKH2uiNZ7GPtNecKwoLCSpjmlrJ4upCDUjUDFMeqGtW4iyK
Fk58NuwLOyWrGZILmnIIWSA0rruUtPk5idZutKAd/2QzVX3z7XpN4xklhbqDgzAZ
dXMVsh7tR571wDNMSCa6ivX45axq2TtGbkjWzSFUzTj58ltVTUalaX+AmoeDe/Im
UKiTxb4ICN/eGqWRUi1v8q6656y+47Uyak/oI2va94afxZdx6IjhN+c2MLW7s/ad
lb7XAckl77K5dsFtDrltb4U7qCRCKXiY0vbFu9R9Uj+NsOyd/6tARi4spA5DOSXB
552NmUy/znu7fd6GYRCYHHeZHpt9tskkKoXT6hk43etvg7YOCVgBS+/VZzKN5RrH
xdq+BQfbu7VV/wF462ZDQacjScy/V/vcpkOf+2XTGEWj2AdTqfkT2nvrp7UjzpOH
SSd6HB71Iny3SOWUqvo44UQfXEAZjevcl8X17vGIyIOZtv9MDj25znp5dnKiv9e9
ckmqti+ghiz1j0Pq6fQxNOz499/6Ap0oHMVYUJaJ5BkjUh28hx8I/b4ArAFK6wqe
+F25v9I0p1baGlRyngnMaJlHlCLDsrSgJysvxsbarFOrK8qBpNWK5I/I3NvI6ibM
BOsgNYyIsEVgZHYYDoIJaDyDy430yXHJPWGXGRCiceeV33tpWgDZZzN4Blnqz1xL
QuXQ1B/3aHeT6w+7Fs3x7AOAiKJJJmZe81U258/JsPepY1SsTQRLROiM/eRJedjE
V5lm+ac6LvjULYC6J0eZ8ls6gDbQjecrlZoBY54m9maCGD0uCWF2EoF91CcTiJm2
upQsKriGGAz3/6+sf0NfKQpmVC9/yOCej+sOp1rkouIerSzs9zt0/jpBXrar5Y1l
QAVv+ftu7KJbZOiOz7HMvbopkruEyNpjSmjZ69D/Ke9ZUfRw1aWntLn5r81fce2S
dMb30cYdge88R7qqoYB+Ls9lTFXD0V52RKRB7tp7uUZUgaLsCfJMri4GLjOh7yHG
wkwFvJb5VK53rJfoRRpbuxSuWiAlIP6ehi9xVLu70FRgIjmm6CqoXE0SXBgEdAPI
5lNbAVoE79j/Daie7Y3HLaUKS73ha51orQDWVfNJ5XjHlwehYbk+1Cb/z7g4Jcly
KiMALP9EeW62/SRWuZ+YpLko5Lv84eNlt2Lqr+qvHRw9MPyim32Zkr8B9mgZkY7G
FYQx+egHa9H2Td27mh8IVJ/7rt/iaES0YwX8ThDA2CfARRrRR1YzfwBeGVvYGpRh
zuZCjHyvh/O2YoRZZrXqE0PVlExaNjQk7t4TQ6hPXMbOeKJnlU4gWiZ7ZThtatFT
0O/nVYTfYxw9KzAs4vOWXJ0qtjtJSa0f1z719Gzp9Pums9bvAHtUWS7Ho1+fUFI7
umSUkK2mKo66N4HBLIebN0h8yu7rzitc8j8jRQFoGA2nsze1sYZS9Ho3TjsCmZT6
O6byUffcCB6I1c/2zMpcIj/v/HBDTfbT2A/fZoQD37jsjU9g0kKN5ycXLrPm2QfU
p5m0Ohwt3gzZ8wUnj5ctLCnD2hPQAnUINjQPJo9C8khC8Cu3Zkx/QwW2iwAvcCFw
NrC8BG0+I6xCf6++4CZmIBsbK+cmUeiZoQtkKTh5VMBb414KTMYYDGyHWykTGmLM
6a4QIBOx0IvxvRTqWqFuWGBYM1nRA03HV5I4q7ItNp7pLfneDrPOThuCuG50fpU6
u1G6bnuMdVTjROvv52HIIW70dE//dtxJdGELbUGv3C+tTT+8wxf2zn9BFJzVeUGc
muet/a17XbonxKH6XfaZ3Zq3Nxth1a4j4nFftSlPHkNXPj04TRbLOKRkn+/7IFWs
1HShEY0VL8COlKUAshoIIy/xhV0t0bk7NS+cPEToVLieAdCKtSpI1obSPqNLua3k
WoGzuybv0w8s+MGHrKQFfdD6yDDMkVVlzKPchPVJqK6ZHWxRlrSmWAoCIENjgQiG
aovIB6sJVaWbHa8IXln5hYzi3az8BhslWZ//lZeUozyID78j+o6RH+73upebTGCS
n6He3CMuhx6gMgah+jFpZdCRaf+e3CIPeEx3qex1lvQesXPtrGW5vWn018d/wGGr
clRChlEO0hnCr+xlOuDKDzbZfP1H7pqZO6w/boZZZvp4kvl/e08hfEIQKGe0xrL3
lSCfPU8DGbIOzNgLzp+gR+DT0RufvdReEdKhUKt8jodhywAmsMv5IUmoaB6MwiyF
lCKhj4RinM56dLeTO030agzCF8QMYIfpit0HzSo6ym9Tx8APXHjXy5zNGNVtsYuY
v3yE2cNNVYcF+ZhtD7+98WonVOc0hTYe5cudrEsxh7t/1Ww5xiwycNTGkCVwlK/G
u/jE5hTc1cN8vMIvbSlPB1XxbtU2m+1+uzwIT7DGMO2FHJhV2DP2Y+ZefePjig/v
ZgNEaq521VL0wlkJfqDrW9rKV6DMtOEtTnzVSFw4hDqsszlbDPBwgOjQbQ4CR0u/
UN5Iv9VjCzaqSPlJ+DtyLnIHRBesJ3QNg3jk5C0ZDICrhNso/QRHi836c2CRiujG
4pSvopdMxmqf8asYzDn4BIOoENtU9IuuW8HpyPaSZ94zayD76n0+43HTcIuz7Vqk
qWp60zPPWvovAaIZ0NJ5PUimUl5tur3RqtuTpA+5Zvm1G1lghQI6JV1NfPBt+1P9
PViBPBK0OeU3tVhVkIefDws0Reg6/52lvL9bpPAR9CFhqeAJuwoV4nqiFqVAiHmM
N3CzXgScCfb/2DF+XMDMkPfLJY3AYyXd/a3qAkJW+QhD78GNNZuRWqnDvmukeiAs
HZAY1BZrKIMI4+c+F3INA8Q+836lZI2HWp4OGvCCn1FnUX9K3FlbQfcbUazdBRmb
a0vtzuolwVk58j7I0ZRL5W45wobNFAlw6F8nqfilaWH1OB0U7Zr7px1ZkKt71d3o
RJ5cVnlVTeBqiFBiA+BXY2hofChTmfz0hB+4ekNAYwpnoYG/AYD47RooPAXLNbet
N43Qf0a1HXTqhiQAQx8RMBd5+ni1fCUa5C8f0AB0v16/OxCfosBEvcsiBYyhDLCP
pLiY8DhwSsvqdle2WuVfQIIpeWgfFfcIvklIs4itLWb2iNhRP3QKKh5TEvpfCZWX
5RzNvM+uWHDcOfVtuDiUf0jmwZrnmvv9yUdtDzJjInBvExM9l7eYCqmsS4gY2INC
RXayhNqDHZD1abaZWhqpWKuPESiz68MtND/ONOqn1oglakTskEG5AXaBIE2ipx4s
Lhul8LxAg6yXta6k5LA3uoIp1hBn09rd8igFQQnygAH69+YvyT+BPE6SvaXFuh2l
rQnuSftxkZTYR/qRuu2ALrRjRKjtM/z7OP14YMtQK5RNQDooQjU/2TlFujZZZJYj
JDJMVj5ZsXVMkTdwPbGq7Kd2CCIw1aFik7007/lvC35vlSQSXTPGEpg5705Rn4mF
z4zT4OkNePf9luEXQgGl5/XpvcXic04yG/eCN030CItgewjxMEDJYMdyROoJWiIf
9AYoXhnnBbYgRffvZQpvfxSaU+EoZQ50bjiCCBMpjHEHyHJXrBE6UhswP+bcX1Vs
xtHNQrtOr1GNg0+KjqHUHxCsA62yHl2IYalGlReyZuq3fja2cxBS4VCKVUBhBzwY
xb9H+leUcqYtUpuuougrlC7eOafEXjyEaCAsUerika+9JklZUetyO1Yfp+X2eEgM
kIUOaZd2u36No7hhCy+PfHmQSrBDphsj2MohMDiitgUNsbahAwo0PEvDXmH7vZnL
LNle/CBAjYEmCigm7aTsSjA7Ou+hlEEbnHehIGRgx+/yj4QD8/vYSgXbd7otr/9k
p/PB+k+DXBgb43c+bfOzluXWBdHWwSyImkH+K9Fwfru1NO56pQ70JUCvyxA2HdIl
QE7TpvoOrhMdAKqZRgf3sN+1fmy46rM5lrdkFvVfFf5Jp+PgssYQdidskPEp2PAT
HCzab4/YrbvcEM8BW0Koy/23mSOxWZQ77NaKF3IiKvPQv6sYZvwy0rX3lF/CRNhz
tQc+UCyYaweCU0wEF53V+BbY9Vg+fqAWHKUy0NHPh35mf/Ciu6GKUbP12NUPvdjq
Fmia3cbipHxmkPpmsCA+9YeZlc1R1FNnqBNtkhRVjg4NAG3ZD1wZhmaCz6xezahq
gv3SR/Y+Zubg33euYhaQecZLGrTB9OQs8xTInQqZdq5le/Tit2tqmL9JR/an70g4
rgE3QxIFmu5aooYOxkpcp4fii1EeJDeRF5o1FG0dLs6OlBfF6lLHWpugdRH+5MC2
jOhM3MdFu/E+0dzgD+x5Asg8RJtbxUbwpxFspTUZArdp9DC5jqbefLkwBb608fmh
1D4Jgfq2rWKIx8UNXBrnSWj9I4u/n14EpMvqMn0d4h6FDUM+UPbktCRthx/gT5FU
UkoZ0d/YRlMbSB7wcbQNKWYsz83UxxraZiHvsvtXR3OABXO1fZ5/WlZkR6y9eIZ+
VEgDeq8k7GhsD+2uxycvcs/FjWwk93UrChv33rsfsbFKBu5OEmjbXlHsrratNPN9
vRjrDv+eBxFS+PfdQzH79/4b7/FqoWQT2YqX0W0X3AiqNzYOGZ2Yn13Rbnvml7sE
gTieff1BVX6cAf/R9eaiWDWsbbmIYH/yt+xwjzS/4NMUgnIoavDhCwEuBu30n04B
wrxb+lXHlwVoGbDR7flvAqV83xP18C6YaTCwTNCOG58G2EK/PUAEbiEuRIamgOht
g81h+FpMFfXctuDOekZB9cd5+e/ROgfc7DO8Ux80KrLlmXpnEsuEJXJXs5/U9b/I
KhHUBa7uQMHJV++K2TO01sv7Mt+Fo6Ss2ZtQs8V1xgS4WXAlNOkV9OVL+ly1dIyZ
40bDl8R5troyBqHuwsQzMClohA5DUTZjEUeu2odZT+BrbZ8Zv8zy+0BTlY9RXq08
1UlQEo3mbQ6MO1qi3/TDm572q845eA3rkcnZHzlin6ZFiIh2QwOv+twk8193t+bP
J3ofd4sZAwJ9ldW8xRknlwyq++PEY2NNLfal7xHjfKKDf2QgJi0I3QwxDG045AZN
KIN3sumpX50FYfIE094gVcwcw+Uuy6GrpiBHct4OwdSZEQrPuk8VQooqeCxzS0V+
+7X8PXMryZTDyT7JIDam5oxB28kRUi1TBY9/PSI80d2Dx3NIygZe7HTmDPj/RiYc
PVeKxzzjEg/5dUOodV8yPm+DChpjpeSydPcm1xWdaTpVWJr9TjG9jrN1qI4qXWcM
uziDrn3kaA0KIZ1Q8hJtSKRRXNhiWELL7zqTF2x1OO0Rlbsg0WRTpA1cT8/8TSIj
qHd5ZreYJjryJyEMckR2l1wBcSSL05tLxp5W4jrYRZX23WXSCItUn8cnHeKcesvY
uhiz7pHrvBLuVSwTf7S4r75DpZ2V0aMMEqGeUkGbSoLKzwiOHBq3Vfo9BUnbH0ih
hVTKPQ5vGwgc0u8P4f6DHoWELkdQJ1YlA+PH3giM3NjUwJPnZJHAFjA01saKTmRs
2/fzdsImrd3q/oSjql+kdlZNIqRHp/736pcce/qqjfL7fJnx062ZcNldppsBhG4Z
VbDPzwLIk4NQVfDKrfopT1zkf5kuaZk9AnU9gKTyZolABuXE3a5WoOhF8uAwOlmD
oHQbrPjfB1QkI3/YxdKxvHQfa1arBSB2Vf7arlRfzU4S93HlEkXtZKxDoeDUskzP
/YH+Xhg7LxKHydoW3SCbpC0kNcJf8U3TqsHa5AjD/WxgBblkKYka2jLNQeas3Of7
DzB4Yp06y3uMlS4175ISCe23Bvu9nC3wjYKpQJoCuk912SrezQH+7d8bYNWBedga
zDZkCobwl1F/2FTFZ/pU1Ls7zZjGDEIifrwtcf2TWSLLnwsDLcxEA94AvX7Wmd6w
kimcmTgwHYXrhPCre0aljyQuSReNBYsXzTvXTEKg5hHdAZORdt7x3OeK3DjqU4vn
7arBOB7O7BCPJAyXDFlueB+DzRyZ4GSS6MphrO2JNFit+kG+pF6Dk3MO3stq6ol/
nHDNM+xUnY4Ibnk6YbHyxXRzx6OglqpgpWnXBWB+XEIFNlVoMrrZD1RIfakHhLdU
THM33UARFHM1+dmoRdFaQ08z1dOc2zVK4ih24SyoUxDdxVH388OfR/7Fqc5HIIs4
UaxjZ2lEqU0+afPfOnagBgfdvyfq3P4wgyoybuzEtf71W6m1ZKjBqY98xyG/breZ
+49yimQoFipdCgTnNKj0iTv3avXSonsLkE79gwrg3gFMNPil/kCX1dwT1v7d35CK
sIRb6OEuxXgKk37AkJdQVKDyYdIJyn8pgi7X+XBIwG2SuQWaxhlpcyW1vE4akw/R
x1R+vzT1FNoLgip01kW+vxmrQHUasm13t86LJG0M5gnPHOYvuAsVnnvuZO/6P1Fn
SqVQhD1smC9I5jaPRcXhozWHMIOv1EWHrmXq7XmAJlRIWstqY6ktPzuLHoQvBP0J
AAcn59QcXAy7sx6q7fUJfKUbX8DyS/leaUtBVK/sWjWN0CvDt+J1fit1psI5MhGU
R7Sdof6CLZUv9IdGx6wiN2cmW3DlNQRBJzofr0SlCp0mggs6M5RSVmpUqrQAENJt
bnRVCu/QQtdx1zEFG3nQxUMWBZMUvFj2Nr5dIy6zpwNuO99aIK2b8aVERtkLqiiN
Z0UTU1G6ZwJ1aiFrCiExMc9QryhKxtK8VaiaXhRQwEOoROKoURNjfIs3LP1Z06Om
x0p28wW80aCvWyRTCKZ8lEW4YVQTbkgt+CUhD6IG6q812KQxtzOIQvv/yvdQqLdI
oi0n/4JeRPgC/YRK96uqAZdkwPtHLLNAzbqbtsoKh9tZdgtKyDfTgeRDl7FnZZdl
erSBZDoabLM6II7fqwoI6u0KIHTHRCIR1TrA+43zahDhdsZS1iF9UuL2ghOhLzqb
bvhcqRGCWyQ6epGA7k2aa27+SbxqbLykX5mEazanbNZuhRY+kuLQgZ/tcNug6xxg
BVbm43RlQsklcruAP04M7pAe91Hqv2S+EamrUMdK5agQ5/l2RbygMUUaZJoeSqk2
vU6SMKX20zige7UT+rRV30kc4pXoArAuBK3V0uyxvoDoUGkY/es5jFcfvNPybwL1
7l0CagF0IEuHmYj0ghvbfn6spYsEOAYHN+kzelIrZWOwa2zBMPMvjUHSN78G41JV
yyVXrLf3jZD6/Xc00WjZJoeVSJ0L3IoV2eDWbTV5gIgP3wMZZPYD+IqxqUYJD3t2
r5E5xpm4IqAU6KFeghv0g4IKrBpgQnUcWWXBE6LqQytxCM0eIiRc3OoQxaPDi+b8
eKdiw3VQbJzjBkvQgm4u20DRv/hRFzf36ZNxqCqlsP4a9CG7scl8l0M6rFR5fR32
fEonQiBHBOwBjeW5lrORiLbpjpL4GDiOfyc5e4YAC1qKmvlLd8pPPr/HlXlJ2nfr
phveIzsJm8up+swr8ZleFkoZABObFGvvvVNOEw8cltLLYKGDUPpqM1yvBGmIImYE
PaTeNusp1OZlJ7oh+iGXJufty0VOZgl7iw+KhYREJ4qDYa9Z9BL2IjIqv75a9MBA
eQLOTC3OwwWTxzgU4A7747vtDDflSU5RdG7fbGWMi4MpX7H8oEMhF5OsFTWflfuA
/60QVMHsVjSQISoj5m8jhGQX5Kqqu9k33pZy2I2jHYhm/TMbASaB8rSC7QoT9ONw
0+LGW/K2HB0P15VZoc25Mk8+cvqjEZt+nDZOZl4ke5wgoNacNECuOKU75aYcCAWj
fNOnFJKY+rZj3Ke8O80wFW/ix+QPHjwGzfLwCNUYo/egB19dWaKkH5/dhwTB0PRE
io5HweHyIVbc5p55UOg7Cesd3lkWlHSStfVwssgc51ijKIx1XNhBpzAYvnY+fp55
Dl33ZfRfpEQtaWpNrVrEkfe0GTkVuZk7qIIdzGkHhvf/bUO6NYmYg5sFdTFePQHR
V/Y+dltD/etH6vzQAy21iMbIHVFuA5/Y4PeK3uW6eWN8VUQzclc450gVOY3wc4Qr
M797Uz3advCawwy8ti/OxLbPJHgd8dETUADZmeKtvEZPeHSWqo8Txe1Rqq+eY+9d
9dLolMGZaKW5DLY9TfxGc2/E2x2eb2EP3JxvqcDpKhQLL3TgUhMC1TP/etR9RabC
cR6HWEUZ77mm2yPevC8+D8/n9Y+dKnbV9VWCUKjJtK4O7KKj9saVH/7zM87kp3z4
O3anAdIEGuT7bhty7b+rMAYH3OigMcCtxVNAvPpOyncQg2eUTj9h/kn+IuFSlS4K
lXpct6sbVATwTzpmGdCNm5VqYG/1z92+PMonBF4l/3G77DQonU/z6Nc2TjNhBYzI
vRAIyIy3HmG+7NsgZV6km9+yhQ+tUkwu4ZM5FmLA9PR2EdaXZ95WkaerpMA60ZEx
vqxv86Q8+SEeJROkQT7sWuFm0nI5z9wWp8F57vwUpVtXhOMzxzN2XBOPnpoVdvTw
fTeY3HUfvRmmNtUQ8PQhYRdfdBFGRLOh9oHjWG2RayRkCSlUJ1I69S6LiOMIbYHf
NY3HMh8smHBLB2dKUn3s3Xz0mWmBXVQjuwufKbJ41FJ0mfhCGV0m1vrZyUPedkm2
i/Bvfvnl+FQOhwBRJ9cQb2J6u5YjJWhkIGed+F+adE4UdbRmc4Txd8HyzbHq63g5
oFtKNrqvVhRGuEYonEPtS/GFI8F7/DfQqS0vMFGt1FyuBHAQhL3PcEKhRrt+hd2+
V6TIshz1UzJ3OlKsgOTaDDqhlIRjoMOXnPr9CZCGPxwDpBrm2FI7p4NrN+f/7Jqh
07o5P21aQwvoqO5GsvkCmH8zPbOp+Xzac9VLnIYvXZoGBQHWyAQxCrJRTBDIZ2X+
718eyQINCJBTL7v/RwDAthNviTPIVxSFvls0YNvOp/nhoMSD2MT9f1N7Kp/WVuoZ
X8DnDfHtG4hrdvRtdpu0RVl5HAYlmzK7SQ4VQwsDVi+LaXfqQyeuASsGXQLDYhGZ
zxy9mcaGIvY9rR3UWc1ArRI3GgsdXET98JmfSnkwuBMeXVQmG/1zEuph33OgXOVD
xo4UM/4et35bc+VXgS9H8t9Ul1ZPqSYpSNDZ1pv+0uHWYIAqOu215C9ilKZ6OwSR
sOHGlj5U1ILH14A6X+K51dZKfMU+dEeoCtP8e8fJj3iRPJI6lcNmz/18NuXVrUUD
U69xtd85OwDCljwT1E90DF9qUh9Wv2kbcdyxBDh86csB9ZF+naVayF7NjI4dDeHU
OxzW36jefPolehqb7aLAQuVFyFdcydZZFFKLEJvsAAPCGCa0d6lqrH38L1qnuV0n
0I9YK9ihQBCgGVedbj1RiB/RCGSw44+HB03kd7H0JJ6uITNVV88TA6zHSXTzMP3+
2XxNQokV1kfp7WjBcgaTr2kRez+3DALh6Q2MqiRm5Ob1Glsg8/LzbxzISCz8O7Wd
WG46rh1pfdAedjqqivaehBiautj7PaPvPoQ7bw27gqbcbrhnjJ0fGfffurgmK7ui
AqfJ2n2vsgWexNrULpQ+1zPGz4s6px3D/tqdCGr6gIvZAnTJHErlhxf7nESvdCTG
9nwDlFKZA5OH50La6BF4S0iMRMFiP6oSOQ/3OuRFRxZdpLIUxnUDQleW9pVj0lRj
jZ5mMUWNWk8ThiBLwhWQJ60n3nr7JIbNfweT942JEhrQzBMX3c0EHqDa99XXsO4X
Ow3HxygGjSKdwr78u6HxeNg1DyZ/6nj4k+icorIdUHqS00TkBKKsVSc3+inWLnNI
NKsEhpRhbHxBzSl++xeV8dRnKffWhPAF9qvf2/Fu9DabnImCp+xuFUpaZVJ7uU8/
vzLxWWnDA80XhPRVR4Icy6WAUrf7A+zn0sfJ8bhW096cENbo2BLuF39ZfKNj1yeh
YbqqUTAzSX4PKNfWhCWQdFsfAu6bDs9piQ3FU1+kE+bpRxC2OniyV8fmie+3RYvz
arvZbQCm9Qkf4rLgZcqddV8uFWicXjmzsprNHF1kMccVULpZXzfmbKff/VK3VTpe
8Az7hplOB8V3475kIruOfzF0qY7Q3YA55rXSXcSz5qoK7hXldR+wVzesQmG8VufV
CG9aBUH2U6rRLPsoIpT9wJbtynOz2nkQDEO3hUaWTLOi0bqUAgaysfwEkBtjHiUR
EXKcVFnlxOnqj2RMQZHiu4IaCZBz7wwP6uToj8a8tq28o00EWmQsVkqMZ0QE0PDz
mFyjc5LbOp0NOOn9kcVvk3bzRnHo4rZ6wqymnNysUga4ThYEQAUlLKoANWSXsJhi
S8GUEJ8aDqLm4QamvNuwPCLuWoGCy2SVyvp7w6vOOkK0Xm3rrL3VniA0pyE3DSgu
PxOKgzuRZx7WBEjVleoIbblhhceP53se4N1S0VOKWwsLQ2hRWzb3RWVRNgxkpFyH
UBbya6VGmbpIkwVRlZDzEtXGz6k1hglieS91/KnHIQ/B4VsP74sLoOGR/7vJfSOE
nzts/L5P6TJN18X0hphRnAFZVomriUiAFq7t62uIzBsKDkEW/ld++vp5rU3EHiJf
PBhCROlvq1xQfo5W/UzAqxnQCPaaefd9uwtQKYCWm5yYD1T+ekYl5auHL4nw3mPu
avs1fYCb2Y4qoeqCHmx+hQ+dKgMVOPD0rEhXYYNTqN5AWjjea4I5eTfI7JVTSyL+
IPmBn9tA3S4xiDZmJtC9BLPX2M325R9r/+XIv4YfYxiFcwzqfzbbWkxNq5Mp1Kne
Zhn3NKPeVDxTzS6h08Tsjz8uBAwOGgG2rKkkOmSDy0U5yY5Xbw1514zo6Fd81CEU
Jji2yKx1snn/JVvKuRQa+m5Sj4xd3MKCGJMzdZdwID+YV6L7eFlOoL7MWF1z6D7t
Jau+ue5xFfky9ihRSNAnrBhGzU6Tqw9QK53StmKuUl9O3u/YmCnoLAu/2ywp1XZc
RzQuJzpQx4GktEUvV+SbZiEQAh2K74GErY18DKKtaHrs4EOfK6xON9+Z9N68EKkd
Yn/tKXFiFKDiLKim4AUPYmZC5b0ECeZy/xNNV50c9UCFcSzPB7HSFpWDVjpxTq99
U74n1SSbb6oFKokQ4B+ZYvyOvFW46GxxNSb6i7zgxBbJO+SxphQ0zFAyJc+p5Bby
w7h3VL+QMjUKqMnUsPkJ7ghuraVgouQXInHBV1cSVoMirA5GWi47n5ODIznp9b2o
ZIkqq2BcmTG0AbGdBa5sjZLipz9WdIY2Enm3CUPH6EffRFxujgjdA2OtjgTu1aEK
Pax9NqElWe29pr1m7mVLNZXAbgNNMnEhMuCCzrMvBi7nGribt58HdyIE8r/AD6Ih
Bwu1+ef4hRnrpupXG43P2lTn569Eoj+z7HzpjDwoCddXjYz//UoN1JDIzRfPXHOl
XlKcaW0BnDbjCXv3IBW9HDEHuhfyg2aMyALptVywNwz9/7d1emhfYR570kGBaQPz
iEPKkn7jyg2vhvmVqBihmj1P3VY6giCpIrpwmJ/189i1EogDK2qYVHhko62WmgFQ
zsGzDoeT+EZZeOIBEftuwmu52Xl1qJrIVNsIVcbWq6knF9oFpT701gqxhgTzNRFQ
0cHO8mB0Q9C3IbICd8kd4IUUjJ1WAoJJAMWqXwJkCzjyZFIKO6Tth9chdLPhau7y
IVAsoU7OuV16Ns2j2RrkPhoDd03yDycHfD3skhoMaoEOmaUFy54zKW/U1Rz13Y/h
hCnUSTYbtQztG3QDLE3AXsxRTDEs9EFsz7GW65utBzYH3qtKgj3fQj34VBIqCw4P
sdAWD+K1J1/Uc4+GlOcOOiOZ7mtNqQPbpzZsNzas1aHvX3ourE8WRa3kEI7jTr4v
VaeqvsypTOwmnHx9uRCBeHg4bQD47t6XB8NQNsUKAneZrovPMld+JB33GcQXpT2p
R0BrV7lN+vjrWvyqIzwahJnhu7vAAROdClMsuMIubhrelgsGYe0uL1K52tkk2nJz
NxQuX/c4XKv1O4wMDS+TefRIfHcfEQESYmVZFYloMBLmtngLtSA4w8iI159cBs8z
wvIeKEfaoOULMF/0gqmQD1v1Nak9kJs/GHFVYwEaN8ed4X8sxfrMvo63qfwSkJQo
Hl9uT7ICuFPOoc7XfNmOlo7cWMwXZgMn9B2uY5PNa0zVc18TToOJwlC81XnWUmNJ
ncMVtKDQDutPLStLoJVnzDwq6k51u9kvqt5g6zTJpynRDzuBin/vWcP7/N1019I7
D3CUjqwdwGy5OVV/NMJ6pHW5J2kSA84OQN3QfMG19vM1a41ii3xmrapfrJVjn0FG
6ib1dqCVphAHIAa33wCoR4GUCBd6EeP8D2g5yFGnpvIL7fuz9FG8CKap1tbqMRrG
evnGZCEA2Y6MAnGk3Hgsqq3nXH4vR7g7cRWfMI1V08AIiUZeBtrG3IR/hfbtWzIX
G0Djfzn8iW5oQZ3iSj0S2eGHEWsRg/Ieax7GzntwVLO8fRy2kmTRjo7go19sNe7s
cSIX6E5tOtemwvZjCVHcMO8PxR4hMUz7OPjlcrXvmX5fOTssrUCuxUBzduRy7NVr
sc3Song5blpIYv/K5l0qG0Fuwe/dOIfa8u1UZuCioaKF9lUUCTGE/WEOcteLLx1f
oPTvGcBybzNHwU3dDz4wruv+TN4y35YnxMU3rbSrDJ0BEHM47nkG/4qXYzKu7G2k
oVEOQruMvPrUJBHYCvA/0t+RU5ddcvAoc5zonWN8Y0lMgu9QSLbcYXAFqLTx4PWI
NSjopUuhdfOrz0anxVUXrO5DeCTD+Uq5p7TkC+vNDxOc+xU4SZslVtm5NazvNyJa
LqyYUHvpOHAaO5Z5I1JWBdk6jE7TWsAIj5CQENb8W/TPxnjmzc67vcr5cJhh8uH1
FX5vew4VVQNfcmex9vCqjEdfg2f6gKtj6exsFqiTkLPzO99wF1NC+lg7RL6c+Mzc
vD2OzHTSDM1bvBO/4jLm6VCJEO+3zjrzXT/JJeSNIPpb5oF9SiXWU0zSed6dAOql
b1B7wPmqmIcIUf2yWXdIg5R2wCuskYzDsptsRLFI2eAL9skihk2fr/djdy0t3rU9
DyzIF5Rq/YgkUzRBRUMCt6ZzbOjmDZU1YIRNSq/hNj8haLy6SsjK3B4/ot7IvJSH
Jk27i6SkAG8bVY6YCe3aoXdv9sof4LMWSi3HvzJn7oaAhL6dEXvTh6DlPHFCS9D1
kdVDF9BVQySS6FPxnS13v/GBf5ULtwCmfHSzPHtqpiq7HPnVD7vkHrg9U4UOgL45
9VWLaYdX5oXQJPT7hs1NzY9FMGfo+MbexAbVXtPhyoYUnUqNepHr8mucBHDBmfxG
81MZw4gjqeUF2dbNlFB1WYdeYmoAPc8FkHzycOkfW3zNRcPV6MASW2XGiMc8ah9g
XuNs32Qe2gA2Da8ihKtGXEIgCpQm0egI+HiPNBpDaGAZm2zYavD8AjPvDGPXHAYQ
9eKbN/Uqgz0S/4Y0xzJ/DoDS1kjoua0pN3ZMLvDwdbYesjZAdfgxD0pnYtOCbeNT
kdTSVBvAOhH0GPUl1s/l6nny3EdMf0uo4++5ZlpESE/bMP+Cqa4OSfexz9wzLgEV
xtIEPjg2uTEHu2xO2FvuCm8anZ8V9eU4ku9fejj8ptN+vdn52BJZe6KxBHda6f0w
uBCEdDjQp/0rYxbdduA+cdFWb5RnOygf02WtOFLmFjGBMq6fQye9+42PC0Aqf62E
VnBfkWbB3JrwDSv26rVaghmgZ5LHtVQc9o6P5W8RPPLXUaxgMHhtkcPhoxzJUbz2
keitGbhLzB5GX8kXqdOr+NXOuAMC0jrp9+7AqLU4mQFfvzrs4b7tXrpiGTYxptD2
ICUZw3goU9S5SQmaFoYChpNHhLN9wGFivLsSdWS1AV3c5na6dCzkg11pgYg9DFRY
XaVXCFq/nITsMqpnkiPMUIfElWcwKpzm9bP+QAlY6vdaOAXRhxV8saR+3Kc4Fh6F
qaDtmGLf38s8QXeByqDaNQ5zQE0FRFAAXTztvg1wk4HxYyGeTEXD9GdtAjAkJH7E
F7irxVBJy5ntpF6L4i+96PeHDDyi7cspedhDgOPO3c3Vn6LDpYbwyPQ9CkrPvsQI
dZz37dpu/WPJvMzgyvNLGbZTKPqkiUmaSOmsPeYDeoT6/ALrrVapxcHyJ63ALIBm
k4PPobr6E4IySdFKFkXXfzzYqVrUY9Y1/QAWOIe9AP4Z6bVegfwYxRdcPeE/sGzU
I3m2vVVEHUl1eknyFyk8orA+aLvq62F9mZJ76satQmWQq+Ox8bUSCsEacfO0XFoD
UDdPCYjejbS3/EAVexPnyOdk83S69Sgep8P6Vc195NDhgfP7x8k5z+cVCLwrJZRx
rf98P7gV0sy02MKY1HHUbaDLtHRtcDdjzoqNd03NjRe487QtW7rGKU8Rf88yUIDp
r1b/QHirXP7YN9la/3rV3dvXLIb0837Q5ASsHAYBgHQ1B6//QO4mm9kIqHJ3N/CX
afpuuoGJhnbUh3TFAWwzVIyBsBkAndAVhnH/ZPOMWYpyRZp7FE0A+sIN+6CwsWtW
OLmro+1w0ozgPJMipSd4XkSBY2sgy4AZMVsZ3lRIWdx7OvIQirjSEFlOjUKJc4sp
Zv4ctqylXKXRQ3qDeN2RI8LAhmb4kSxlngJKigX5mzAvmDaF5CyaI5/J25ea4YDL
Xx/QC0UQKvbbOQA5l+IcTX3Z478EgqeMHcy8cT6PBjCyolB3QOADf+jqMLKjMHDD
PV1lfGd4RS3ctJsHAA3gMZuZCgaxTflpKoTAyhOW945n3hhRo4etAxKMh93jUlPt
Nb0n+dQf0sy7+x4k4EsIV9LrBfw0ybiCE42obHD2N7Uiz2+uWARjOFSl6ewb10fv
lxKxy1OPGBRAzoxAgQjR1PlMpnHEBG8Uzf+0+M0e0Yh8ozNPJxv4fZGGMHEaeA9R
EYYa30NgNP7kac/1eGzEqlqBH80L5b7e3FJlX+N7omoeKzBY25Ro29E7t9P9Nrgq
UL+3i+rYMSInzubwQcn96n+uH89cT+Qu36/+mHwTkqIRZcaXTHLJGpyHX3XGeYIz
7qUuiNtXf/h7sxoexFzNpIKxE5mMnu7oZ53ApyhxT9SwiYTO8una3LGfjsc0V/zA
TbwdK1dItxZRCUVladuQf8/E/t0xlUI7UCayN/yLUNyd5yV07EnD8TcocjP2Jlfy
jmurgkN8P8bpBP3cSmm2YyK0rKly+ubbtmwkGDGsjldiYxAtK+rLSNgGJi3Jq9wa
WeJjNiDGNhK7RqTw3o2AI8C19Srr8OnA3vNeA8KHOa3ISM0aq+xc5IOitCrMlmtW
10IMuxXEbrfHygCxzSZUPqPBl21dMbXnlzTQsjmzyP8X9bGnP/hWScrf9OSJ0TpS
WbMjN/WuhuVfC2aEKpl/l6b9d7/ujIna87xw2NJNqu1M/JBGat6vRyceqhMS2/ge
n6MiKF2Wfxfak8Se8PkLSqBZ9QryxS/du5mCJJTispWAuEKg5OMcfwpb2MsVDuXl
viX8k+3juqlLdxfbyENi6qjlatgvCG8iUeGOPZlb2yN+dylIOvKpAC1chnKijXIp
ULtwI2INDT9b42h6/naY68lWhpNeURKmmih0TH3LWN2Md4cNaxiWwKld3LSqyfjA
uz0YF9TUblkCDgG41OJpxuIK71rpRQWsa6W05WgD52nmnaQeb6Xk/ltyTNNr9AYT
409xDudZLm3L6k2yapvxt4P0kICq2XIzi4mNsnJBw4X8UDPQGPz4AMekS0HMnbgu
LmOhZBdQ9cIBXRsWmKPUyr4n6dMQQeUrSjy90ekOUcsKH/dZXSP71oaJE47mW6b7
Hd5+lpbNrPrshobEHJY6UyBlEEXk1T49YYfCReD2S/uq684rOVGzleq+xrQVFKQo
9jY/N9HgohFUmLqnDyrCtdZ/QEM4uUR74eZWlNdWl02hhquDZaJ+27yMqr3DXTmm
gPLlUvXmfaHzr0lWr5ZZ/m6reh39rJuVOku9Y1bzS3oDQNmu7EIucn9YYs37sDgq
EIwoU6kzs3CquHY4XurFebOzQIqCRYvbGDgA72usGiQDm2pcjLhvhAw+ocL5T5xt
SSmn5CMY5R1OyM+fa1BJVW7vVHtctK5Ntfpk7S4zSkRXgXy/9tjdmd7f08fRHTZH
K2ZNj2PnJL7bWQ5VfRGg9GzLClqBbl3PurMlABU+e1rr5EE3smgPF67eEBLmg5oY
Fe/GGjY1SGm7a7Zd1/kbz1SxatMaNihoSHKksN7iXdnJyAOEUKTumiaDHvxdDlqr
QqdH0jJDMs1/1Fd6h2XelpEBcYalWwHkZ8r2RzjPzpgfT4bCTW91caB17dzATJ/X
GfGYRYLjXUkjSSSzNciiwFaZv9i/OLfJryi/qHRv3PbiklpbLS6lYPHVaxwZ09nB
IsDa05qUzUPi2WWdSMTuSke6dNH1Mzvg+J97JcXxYnU1Q70SER5cQ5Z1IrRbfbkp
myACYrOv/7oULEytwn7IqmUekJYzy2N1vo3DcnxZXi3ZO6f61DHp0H+ETuVzlJrC
eSOKrCSTl8eArtyMJBPLK4lW3rOAY6VxFlMXGGa8X99WARcLpLR17/pW1I+SSU5p
SARoJYcmG+MrFZd4K2oBxoQkLglycNdaVf5bMAD/E0c6JzurJW7mp6vErvPxPkrJ
pyrcdZvqXMqLRIJGkueN4Qvu+vApLRPn+pa51xKl5LZtyzhl7dh8rbFDeM0pMcGW
1hwmwAa8o0E1nepneMLwAa93jlCDEuoRn7WEpKQHWeupl6hEf5DV/vG0ucJE0lit
WvvORUfJln4iCAs2jyKNf0AyYoNTfTGCm9uNQ21hW7P7q5XFONQ6AxSQIZb4L24m
R95DYbMc8vWcRTVs91GGHhV+kJHL6fLIqx7+0UNnQfCxC+8DqJKKbPwiETQDQH4s
vZVc2r7eiYgNZp6XgnaCEmvgWcZZXHN0QE/M6CcxWc4f+HzdfYNrD9BwzyMKQ4BG
fTshaAUTB30WXbB3h+FhwCfQLOVaEeaJ+QrPsd1KGBilCg/EqvKhTNwBpW9zQKNv
dc69HQO7VzYrcAeMxGwTCFGTDGa3w0e5fNvPtfd21zSYSDBm4WVGs0Msl4mGKZ/a
fAXN/I5HrC+1LimiY4pU4p3eyxLk1g+ae1APMzVY9yu81fhGfzsjaCVsKYKD8CM0
bMyHDTlh4IiSlqq8LXMbADIu2IXxT9hmPONuzkieaRxsjU5kWCGNde91AKWOiXpy
QH6ofGGanXv5gUp7AvBEAS2KRDzIoiyArYaW4/BquNqAkUocSFRiMB6FvOtLQ11G
JFzRIAcyYcI14psZX1Elbys18PKeTkd4H0QbWb37V0RFwmer6+hW1YdtIwLvJ5D8
suOnAfqMThRvVenE9fQSiyiMRWUDpj+m/0Tz7ufrlDOsV96YFhwrKD1ESVKRF7Rf
lFYzE3sT1vRrSTYZHpIJGdkJjrf9GWvjKlO5eS+ETg0BTBPns7j78p5cYL4vJee7
Jqhtp3Bh22szJNTN3RaqMGNygMNgcxzUlemVZ4ni3mJYMsIQUKJBrPRuTm6cWIMO
stfwFP48KNpxlvWcLpf8/Oc4aKWOLLorRMLZVR3fljQ+9XFrZnXRU+fff5MipH15
MU4pKcLRX+7ipG9vTsoROIw8e7/cgHrYFCXM3s+NVEWWghaV22LULBYxTAj9sP4m
53A1pHXE2OvJ+x3WdK04VZug/ZO0QDLJhffQvXHG86qWy8TcASQgP+hvfBabuQqE
aukVW6CMdxp2EgShZIILz9jHqSUQxQQn+d5X85v1tLL/cJ9ZOZuBFOPs3CcqOSWU
jaEuBvagnRap/h1Fu6WR0P2NmDZgFLBfK53WfoStAQsh3YXuKZhfw2SS3QmKrewA
ChTRYO5BVp6V9GjXSL5ykihZIlNWXuDTF/k780VLayjJZ6Q5PDIn/5MexPbgN5Qt
wBksTw9zYIr3nqoDspyt1E/WPSKLZXjNF1fasfmX7TvHi8EyQafDwVswvWTC5UJY
nl2ppPk1lHkWBz45FI7fuWdZvVrLX3cKv2m4ANccE3hQajSMBZzU4env3tH81+DZ
GJEZZXPYReo6kVzdeuHxpeqhuqZ9Ws8lA+lKoXy7CxvppIz5xWhhcwwOxkwLyGT+
51RNhepBwMpppqeWvOcHo4RA6f/Ja8rMm00HB5iRnjtruMuwGjb1kug2dMnvem8d
vq/NA52huOyxFxygTL7NzeWzs15859RVhM1U3ORipTmnRj1bVfpO3PrllNOOiLaJ
ZGEkUwvxNbu1714lW8Bc1snalBjyNfDM8yD14FlyoWocpMiDdS3aitz7gqjg0szQ
sHXMc2CuWq3KKBXndQghSQwkM1aJcd5jfH/KwThemVJTSrwdSWf5bK7ctC4VYoCM
q6HxKrlMFQ8VWSgAGKdtgVeL/vP6jsYPbzd06kRphJnIjyJK0QdD2B/DehcfVXdN
vUUz1H73pVyczY0v1WViZ/4t4V2QBJOoPHfzpReQyFixjOQ2/YuNWD6ztaw9AQpA
GYaVlTsNmFhfjW16vCYJMD6rmkOh9ZzpB2ydtLhO40gPiv/ISLK8Whay4XQRVvFN
GiomHL8b3RexjOdrjBxI6/EgEqNNVrdmg6RBMoFt0OYqRl1eYb8mM42lrj8jBIHw
vvh1H6uxl3gIx9h9SA3ooebNHat0WgNsvglWYSVHP7UhIJaraMIBOEz5mCp+G/Aw
itI5bvnCzakamn7Z7p9SEQuLpYfg0LCK8xWejPLHqLxeAx9SN9XDdU0eYtGC92Lk
zfASEzlmSqYJO3Ao2/Msm4hGmuEqNZs6qM0ALxUezIGe5bIqaZHsoIiSA4XSE3Za
TrAdIyGXe+dqdzO8C3JiuDGG1dkX/N3EF5/KwNA9gmkcrQ8Et+f8CM45KRvjErJp
3DQHX4/KE9qgszwVXYelJtu3j+EGNhKNhM1qiBBc4kRkEsocoFQ/9fD9o45Xk5Lc
s0yJkLNHfHT1kt3KF+AE0dR1cJyHq7+MKcSogTSHOBulkNz5N+BdU7nyEUtc1Ha7
zhzhBd5vpSk2RtnJRwzeqb3y03A8i2XZNAD+G3pQAb1KsYmY9g7ZkxSu7LfnZXvz
YYgKbj3I/tc6Sn8r8YhSeniKDuHgnJsciv6drpYwkaVLicahBm/2Iu296QqRR5lm
SlNUIRPmu9zXb9z7uDDXhjh2mHaR1A2+Z5Q0z+NiGqJiXq1wK18t5cTm/69dLoSs
R6xg9HJ8vFNooQnGrf8qFDcpFdsRb6h1IhL6RQX7tCy/snsTm9cIbFoUeVzYxnwL
sZ9k3DOPoySKqw31v6+6cDG/+EheOcGHF/V9a1xsrpX1ya/PZIqVSvvV/b8/CTOK
XC597Dc2tYK1gDTMXOj7cV3KvQJaty7IlgCo0VSXgv9LmfZnw1/zU8Q/H9prDD8K
y/a9cl4gdVGESIHPHYiCreqSvfyerNReIQ1ujCAYsCJZW54E9dTbrPwWBef8h2C2
WKGF17n5k/M40ZxLO38Ojn3IYkHwpZKAND2IILB1lcHoXLGWAi8d2GFfWFJSHu2Z
Yt562QD0KczDnctahGPVv3N7zn20wjJrbgeTy21Qwj9ySNBizb5CXPdhf8xkX7Uf
yMDb5DA1btq55KzTBkVNA5Q+F9mPsOrmJKxDvNfCjcXD+xwM5w27mwkWpAd0TQDU
KqtbayfVAdxyGHth1TuizAkI6jRo0v+9FcPXq0k73UUrmWsfYR5fomds1d+7tsJe
04tMxaVHCDRgf6bJnggWbJRc+SbwwAjgVaJzrjav1/Tvl3A79976Yjb3UHW/AZom
23qPZxy41UIEqdKpIXMAgY2R4oUW0zBkl5m6podq1U9HtB/RHpzoF+8uXL4npSy7
mtqCJ/Ju5hTWpKBLpNjyhwwMdAh9h3zI517zZ3BibGI8bCjfSD++9rl8p7Wi1L3u
HfvS+QiU1FEjmf1zMGUFjIkZm8djCpPN5sgN5m7X2NKAcKDSlN8Q5xXD4uBLn+QF
gGv7r/37y9a6KdWq8VGQvJGBBSNJLeUBsqLTURQskkF3Ydxv1W7dw39LQ1qtymHI
Llh1I9uqRRfAoCd4EF1JWDZXXvgtdEV3o2QEOvkdEa2r/SDG/VzfLWYuOaOLDMys
OXXfruQbnZHhCyqGQSx8XLBQ2bLlrblYwYY/fCBTw6R/SIVgxvQV3NQU1vQ1MZ7w
6NEEw09A/9VanNsQXDKkais1tVcXwXL8VFtDkR9JAdaCOzwi5H627cQ7SDoDcrQ9
6Hw1ZGYZwP5jAGI6nLrIJRXrniJ/+8+0HGLFAgNzviJB8rrtEYiy92quD4qs057l
pEy1A2b+k87xEJZ4NB6S4CM2tjzJK9erOTzlOixByo1RPiJ2nyZ2bxqnexiCXPqR
G/umyhn1GJNigmmRw9CUZUIRG6nfWL6B6Nu7xYSd39hUe1vjOmBJswVGwHDIsyZu
2RG9jafSa+e7pxAizDxIBPdOnKHHVsPUQL5eaL9+qWSYfD9XxhKs9nz/eEVUSvA5
fC9UmlXYorVRBEDxHS9WP8l3fB7tKmvaz1zNrDLHjcBJ2K1KqE3V//nC8Ok/Cu1V
F2TU9ZvbvON+tTNatokYI9NoJvXjJUFN00BIC3scjZhH409HUD1nAjVc/hz9C3aD
YfBrI45fwOuwE4137wmDwICrTuAy1H3R5d2cW/4UGtbDJHmjJWqCvwoRkSMOTe9X
vqxX8fCtO2pWmCF42MSU92AeeRT1HtFxEZKRvG232XfrWWHXCBz3HFcwxu9yNO7F
7b1bf9rMFRZ9jQQ63r+L5kR8VhTQe7TopO7its5k7Uf4YBvPnMGaQ76TgAPldNMI
6sgV8yjBs6KAJu25QyWM7RbbDrM0TuxZSSXJcXFJlhk/gMhviHUTxHhggUBUQzYO
y8JhG+20PE5SOaOiW+D/LTJ90W5BUdSCXnyppnwn0cAukD7ftcsDKzN9ORPR8zvC
1KCwFykLbLYFm8KypGshByQzZB/zl/451wj6hDx4gF307M9VQvP+vNkQth1O2vL+
pFVr597oDqWzjsFEcH4suNWz8BXls3oWXGSXDWfUXk0LmRTjE8GsZu0h8QlvM4/c
VOpWwM8HzdFONacl+6irBY22oNZ2ze+mXidxP0wc229uXbhZwO+F2gYJ8P6TqbK8
1lOC1sbsqFUEYP5GKKzTo6BC2R6kegKHBdU1bCHqUTqxRDkZz5ZEmGZIZ9EqfdP6
YN4bsHEYnZuGDZf5l0SSY+F64+F37H/KMyk00MBZeiZNJmlwrDMb6o7z8LzTTLGm
I9/IXGDf1HG+wXqxS3e1mo+4XLzwDrDibrCZxQ+SWRdOKRQC6T2Did68vXwgJhfG
NtSdCB7vtXxycPC9L2P5+i+oMpvQhJcTY0jlsZmjX0OEEhziyva+/PXJ8CeUxCPv
e17eN+vlCr6DAE3P1InRMBVE7D1if1872ev7IE3QFnqHTR+3qU2f7zu+Qwqz531J
08qyso4U2qmoFoiabNz/pdWVMkuBkYLQuo3xF7KP/iCxOEWKx6mPP62oE/NZvLOo
rpZ7gOFIlbZ6n4Ze015VARmBZHoF6p77yFqAFPPvLltbbf/EfPyZrJr3c94VVpTA
ZZQygYR6ohWg9Z4jiCqOHFoHl74+ugTQ9gJ6szrpvcn+aSZO5apzNsByDKMQZIPg
QQ9hQ7YfaadQQkrQR8b+61sWDhCaGwOYjbU7DAwPJljFE+Gk2zsD9M0UmZ8ahxcN
6+S00JX/4A149wGNZP+R0Qny5SC1FdUgWGicusmNpq2qWna8dyvDTiLP3nwkNJkm
pClJ4wVJygJhapeCcF/RX2EJgOhVYK+aI4qgsEeOTvrIYajB9fus43LlYaLarOz1
UBuNldYa/E0m48RI36e+vusjkGp4vO3J4x9LLxs8CsbbZkHjivnenlPrvPKPx8wA
6lkx4TzL6bsxhkkDV59ydK+QLIaMtouNdm4STnkrrDv+VR0r0DWTwreAjW8SgwQt
OO9Puo8OFi6zmijfSsNHuzw6tA0Js8pbAAzibIeP9ie3CsX35whLS+rWYdLHZ+8M
LuVqXF+kCj1djRiru7UjlsUyqy9OCmRs3BQ72oRvWsfyB3183jtQUY9C58rcJm9Y
JzL7Za83sFPnyBS6YXSG/q4cKuM6zfXklCF2SVE8NIeEjwfzGpKMxQBsSMvDBFvG
nicd9qpoHyU8hjZQzCVU+Tzcqo7SkjuJilJVXh7oXU9K8Nl557VrjXxHwplSPKTK
hQE/4Ny5I+/ZAO5e4bWTF7BcyxA83viAfE5lLg8azFVZ8ITDSTiAbWo4KJLAc5Na
BJvqeTKHrJEBeMJfFUpSlWxf7L+M6uenwOsujmcBac+nfQYfrcEE8l2Hwc58a82U
X4HpW2SfWiF7psYD8RF8LbzcVMm8nRoVNHxwFRloTyJn41Sy73LG2cM42VZr8NDN
10aJ+szp38VFPkIglg0oQN6c9Lwkhz7OJj2F8jVx4HuTuy5cJ/LnA1ysZtb+zjSD
n6VaZHjw7U60x0xCwQOO/CJgwiOCwPMT/kDeP8dLzqL2sCMuTLeKbkuFSZQVI+5p
sYY317o+Sl+GLu2tIsBEXv2eE6p1CF8L55Th5oPdPSYA4V5FdVDfq/+mt4BrG+WS
qkY+MIH1Vzu/6E7cPEVEaFWJtzrPk8MlIBMddsGEpA5dDkmbC8f78xyb8UFva93W
n/xSUyLR6hexZSlDFl97BqyCO4UO1M9iWDJ7oG9l88cVq5bl8RZiJ62asze9oxWL
gaUlvKICn66C1TTzN5Vc8hVR6oV4ks1Jf/9q9TlupkNGRnzqoA2UJmvEcJNrODEU
sLPALRrNG1M6ufNq+XywhQspCJH4lWj6ocePncha4ZtlTjE6POqGcLsiGg8GgqOw
9dsoknELYJl9qlnI6tjWtIoNuxORTqWOX3mOnVmgca7rPhWvK0cTSxHPjYDO4Wcm
bdtbI6eTQVDlsbAf4GokHavDvehRmsoLfJWz0oVkAuv/Lwx8yGsAh4pg/WBIlejk
DPb7tzNCl5KxXx6/7jbg6UUVYCwc6Y+RhJnGKQf+42BnvnTjjrj0ngNiNDQV7Kqf
ng2tgXqU8ELC30iTPVTHcP62LR7BaiZ2e0oggnLGXT/m95LEinquy7SB5UAa6dtI
Jqnr6cTlkCFNGbtqDx6JH/Dxqs/UNCwzkjgcWQnfHwAScszCpLgQXzZWW42uZujO
gbbgPnzdumMVEHFb6nHWFsV7XtgJZwO1IBpxfVCBs7B4L0EAT/vm1u27UOAl5IC5
35rNi6NRxKY6oxPsm7OKDLmUUviVS6aFLlvRujXijfjLbNNvZ9nWhkB2TwZdPEL/
Wv/Rpn+Vt7LjKzr5r2uoNL8J5FeIbRVldjKCnAXWJOfAWo3cTuNJLNXkzx68zrYW
Kkb16ZXAN2sj1VfJ95NNAAPELwfkp+Kh+JPsP0a7UQ8VcIgFQMwfcBpbHAoqCqKG
GredpXcE5YWURAmEE2H9JJWO4U+gCnNSJuK1YWtWfa2gcmj6SrIztwPyWB3wiHMn
PVUzRUErBioW778VZDDUg1xC1lDVtQEelPzGpmuo0aY5Uv152tp/b6noIrpW70YN
IzlkoPZjtMUrQVl/QzK7Vu3uHWAEdU5tYQWCXay3ZniiReEuTLGC8hwMTCdLo6v6
kfCo1Pg0ww/ZquXb6JPjPNLBBi0/TR68LUW9wgP9WMBZyla4NoHfTGHGpsbApGAT
IjoIUf3hBMJH5f76pbWsqzZPnfInXBQ5iV5bmQapBYUmlO1sGleQOiPHr+t2eZUu
SYUDcFK7CCe9I85GYrLy7joy7JYjGh9iHjSi+s1SPBAyKBt8XTCzaqHpBTBpYapS
PqmbQfctKmiETouISyRxskPfEqtnGudoQaw5Ubjql7uxyTIQM3J7fxawO0mnUlE+
i7uDDiPDIGmSegho02z4klHPnhpXB+niqYNcikj3BNPAhVEsHRhXc3WGK8S5l+os
C3vPEChwJlzSSDN4Yo5CW2zNe6PAwdNqPB/ilZyexzihRBnZ3GG3/u8Xq3u6gCGW
Gmed4nVlNN/MqkGfmoLQkKXlSGMj7YdHny7PhldW2M4qKvd3JsBCxeOfg+6y2XmR
ZGcxZy/e7bnL9rZxyTHM4yUqIDG8KeW0Vp+iJEQftVO6NuhorivHoobU7F5aMJuF
fdDYZQ3mQWaG208/NgW7ILCeNPZvcTQMPJ5g5Taif/YtRUTvN5jKWVzVSUrKlSqs
z8m0F2DcP+IqlYO1vwpU0QaXRqoeSQCoDVnbN6hl12Pv7HRfUyfRgO5b8rY8+BtF
LrutI8o7wgTm72FdP4Wtea6LLc9UyiM7XRGHfL07HNQ3fvu8xeFreXEVD/dqf2+Q
A+iclsi7KMtzFy2jEQWuCxFIalBGMtwiSIxRjjZcQF+aC1G6Oqsqoq6F6EiHi1oP
sFOz9pTB+SBuTX8NoceBWt9y/FQIX67N8s4hVtXvytkGceadulSKY5QO1ASAAuWQ
zz6517a3nOlJBY2SnXDRyc04qvIW3m9AVQciMaHEdrk6GbPLIWU0o9NXsGpPUF9l
0kdXb0/enZ/lBK97xMJNVLwyUw5qxnAklcVM+mim+phOZxUGOcABuxKW4PCNJaXe
srZkQsu8bz+ltSqcFnAquGHHTN4FOF0PUULZg0CwPs7QUaEh5Oi0DU8dCbJMA+DT
IzW9fyu0y7V93IQnYK/ZfQ5W5XIP0W8Sq9moRjcDpwIy2feVXrMPmu/vfe/7vjAj
cV0EGQAdAyD2iQOlE4f0fQREMOD5WFikYcfQk/s4GzDoYqUWDfGDnOFQ9LhX1S4R
fXFxeo7TnAa/Vs+c7F7gNyopqqTaZZ/DtrLIEc5ZUmBe/oJOdU7fjl4TptIhz4ln
uMzdp7wh7pUWh8If/3/ZMyojLG/r7OdaJzwY0SBPbnsIq6W/J4mc/zEwSx697w4l
5cr2AuDWay7gTSiTzStuPs7N0/OROHdBDRJ5P1CPNorESmZ1k/EbldZZZRYX1q/L
c79CO2kCFtP57+UqAWOUqeRfUzgfW0j9uIEFTiF8SpodPVwLf3aLFm3QhgpVFYJh
xBYoLA1KByGYrreDn3Uz1vahWWeiBMwf0Ys1hYvFKpUxe+ssOVowvV7dc6WeOGKx
pRPFcko+Qt3yIg5V0zCFI2HKFacgywoeWZMuvi1lWfuQKxCPF+Cv2LFfNxnLFaQm
DxmXnF8eoxZvO1HQh2VudNzBphiAExsyVxctfX7Lp752UftsDRW+vGX8b+s9UiaA
Uf+eAcK9iC0kpNeJ8CJQ2TgOuTFuJwphJ/I1tpgLLTha8oRucWE7hi/5RKuEE/QG
TFHF4F7Y2wmjlEhC+Z+e2UMpshCjKIw4w6ZoXENyAsS2SKazjb1CJF1EUGJ87RZ5
Va9s95z3r5cDyQ70rMw+woRUuewfmHFo+GCi8M8qXU0jDtKBUitDL3RzoB1rV5L7
ObxNJGk4m+Q0F80xycwXjfB7CNq8OsrA8b8Lz6dFU2FYlPa9wnbO7vtX6ycA1rvm
MoI0CungvdJDojFdSQJzsJzbLdeg25AYbdw10qid1pRtVNoTH3VWhEUijqSQEMsf
UzjwQSSRm/0G8uC0JkaqUnOS+IfyPrhxCNvpDxSz9cirtEV7vkhK9aJPCP23VB3f
tUV+wQl0PRGZId/sKH11qYCBvt80Q+an0se+k+q/RdyGhrsyna+a5oucnsbZz5iw
AX40RjQHGrAKSC0OLlHSnbfTiTKSZrO/HQSAVVxLkv2RJgAUcAdxLVh/pVlsW5Ti
gHJwzgrtlACF2iNtp2pq+EQ3swkY/GbHujNXgfWN/+wdsPGlCTWJ8y6wYbrnlaoz
vXyvaabP2nbRtIrityw+PE/FN02dMFf1QJk13QhNlVPCvj7aJUQnHESy0sZyQ3tO
AP/yhEMpocCIT1u8ubGGCoWQe7hSIRmLoduEue7/6A/lSibsmImaD4E0RiEU0hMk
3exZHDV+xqEJI473JbBRjb0WUHuCP7q8WtjG9X02ODAGnOLNUwnLozRhsOjFaqiQ
8/e8WRuzGOcG9skzrmBBppd0v1qaE/RyQY2IR5VeQD50nHadeoCmKx8MXDDJIFjz
TQpukePZ0/mDplqqeGpFzWD6sET+Qvc+V/FT8DS5zxGYQ5vry8KyvA/vqK2t1FW3
Wyj3M+ByGRKx7EA/HRGZrUvCoczk8fFEST2n+3RBIfbxfnmiFZf5zG2HlS45wByj
bDDvKPkip8VArWlNp0c1R+PlptT5TTQbxUYMnFyhBcTrfp/Ouc0D2KFUUr0Pcw92
HDDgbNcmsJ2qKcIZgNM2V9GAoOL2ws9DcUX1ernGj85B9iIMnqwEl3XBZNYSesDw
7BzeGrQVG9yrYHEnwtIBLiiUe+8CF90PUmEkqxIxRJ7hHvdcjg/Hojr41fp2DZco
9kN+67K4Iv4VTCLK3nPFM/foOWpMw3T2XH7F1w1nyvNiVujzWx1POYDrjwepy0/b
+dvwykzsu+qrvwEcdisGln5VIebxulYL+9J7FxSe18YmLdkZdXUwxfAXixODX9Dn
jrv6RRwlL4qywTnscA+tZo96xRBnQDuq4f3ouHHPpp/O7IXMBnhPONrdKAh/VY9F
jSDTTPY4mFWpHlzLR+zIe20nqfiboAeNAIQgQXArbEJ4Kqq7GW65psMLTqDYL6oh
mDwmfPcEw96Iw3+RRbQeD7B4g1vgDB73lO5+9Yz2FldmE35vuhgfzA7QrZkkIvuH
meKnw8Ok0lW0c01S9t1yCL8UxFgorxr9CV/onCUG+WBz3+EDeyLa3pFXfaauPLe8
MFznXvyPqSWoPU+y6TUkZt0WN6h+H6v6xlJrMPjZ7fCgDeYvpFPmLetVMj4k36hr
lpVaNmJtH/pgJF73BwXRp/hNoKgFYyWzuBRvUCcL4LQnmzbikpmtIpNJpoVplYI5
CUc72qRr+YL7s0R89xq/LV7zwkXnHWGqD0dlBhwHJaKys4n90+E/4w/Q7CbGa9gK
d1H59Xhim2LarNbRsJuYF74yNDSJx8A0t/cjPMfSxyo5K1UvNyZXg10yrfwlieKv
EH05bRzSmjV2sI0Tz7/gc26ofd+P0veB5aOw4hm99dOxqhzJcQm98OJdIEf30xd/
jIrIcp+7GCIYsiECM8m+lDWFpDi3dDsVHZiNb6t9vkxFFuiYDzd3Pq4OfI0GQtXh
Q8A7CihgqJ1ix08AkqVHfkiZ7P6D6yS8WYYrKE/7Oq6RrcuuIlEDtGZMhTTpxAHU
zhcIhDDUJ4m5SStfC8dKasYjuwNMW9kwFrM1CEZyYZSomRVWiywd1dD4v1C83/Y1
6W008mFmqGbG6NXTDR2c1AKWyDrUTmVnogL+0kRYetWyUiF6794kFwOAOndyJ9JB
fRLnoCgnpPxQ1FcYMWDjsCxwCzCRXi8EfZ7rh8+2WCgQEhXEpJQOqYFm5MSO4VPM
xOy9WqzGorkWbtmabwAgSGbpLRYCwrjyquVtNcB7XIeTu/M8iFYec388111CeVrq
RY2Rh6CSdUPtbl2TzdJdcrV2Pi5xU5KN1jOQFmQEGhywWjEyam1obvBUpJ1ILb7R
joY8rl5vo3q9yEP2qR5ZDr7SIZaWg6rjNF3XZk01LWRMUa0WrpN+gYXXNaEyIsou
PcfYVAO1vYNuYcMOYsmOqdNmnaER2YUe3ga63YkO2uv5Jbi6xvFGE2ILrGT8gV7O
HZSiIGIsGK6iqS6lgA0iI/OFzkY6uwQKDxkIxqNgVnhAZO9lI8IsNlPYD7EameQ0
vdTBfJfg8GVPawI1SmkBBe8jmX3qFNEXK3IS3UXOkKQzdlagYsv1ccu9SwAOfPMt
AtA20YMYYINh3HxKVfnLNMOMJeARupCh4fI717XvqGtYFh3veYaRbaHpT1w85KBv
HZYmP3FQmLYuMzkvEJZGOcGiZ8OBTdcG17sQpnyE0kt63d85izlGqRp4gWFWGjDV
ZIZZx/Y73S4PGpMWlcqRII6CPe3ipEV4pUj2QqEWx7rgYrpj4B9pq0YIRK205Zbj
UkrLuMOZ3uSxhNypHHIqybWc3UZ7nA/2OId89nOFjiRX9oSr716mwHrkF9Eh5Miu
q+eZRF9J4X35YZ5v/ZYsJbKKfdml5hfoASb+MI9P+fuMUKzAwrKJKU8cR1UV3vOd
qaWDNEeiDw67ry2hYKKFIHpQjZsypJzMidh/ed0g5ydPBHfO3NaKs+7bqm1+wwDC
alY1W27mqrdr/IqnaO9jKNGZJ19zYJ2Ntv4HJP9T4hb49Hcn4Cv+aJh4uFQgWx9I
xVmkNu8dTm509Hwepte9Iu4+Z++ah7Ye2HfGBqA+vsZRdOQ13fkH5P4qy/y2dagO
Mudq2Ka416JbfResO2LPv8vc5e2vE6JQIYoi56JXZan/heSoegD/+/ueGcv1XeKp
LO93eOf52xnxZgbT167Xe9MEFi7C/9ab9d/2BQmqjt2ClqzSCWTc0lNZ6INoK2QV
/RJtlTnpF2oOBe7woC/ZCeBStVtYMIZcA9kENCKB/xhyBrwLmXHHUCaE4/5vRb9F
r+qBbq0VlA3X4+dfrF0uL1eBMzIr4nF4XV9jwJDTzOorQSC21wLrAKt5Mv+HyJ7z
aow8LYfYSQbyXgl9y64ViAq6wCiBgP/DAMVFjwHALkyCQretyap/pNYgxj73lIwS
L6O8y6rVqLiqaSWk78nQjBY5rsGl1LcJyj74iP2E+Mv9CPfeaTV9aW/DQlnG6U7o
ZQP1f0JtyB6WhoRTO5ROgBpni7O16nxJtidIHvzClegLWgsgLrpw79elwTWiO3Ef
5ViNij6ChfSY1bwlkUq2uQrgCBgZwwvDYJ1IqHWVXQoqlTUDbfQlQo2oIirzUU/B
G1oVFith2MLXPPH5eXhFSEG5+Wk6v2GfTuQWhn40zG0nTKvcfyHhkX0Ds5uk9dYo
GfMdvGbzAY+5Se4SaEHibvSEWnZz0qPnbmAA2iNRNoWEK0MFkfNhGn13kTt1vsN0
HKM6hwkyc7DQZ/OOZu82TmEH3g/NjTsWEXAsEqnq8N4FAfrnr5qfI0IF4l8OOHof
ZQmiTDzE/6p8+p1CvEGuzZPaFOgb2LGp+UCGjd9B0/W5ehe0ouazGHLlIVQ+MDVz
7TTSaw89oP+6tgydUOnkGv04QLmW2jWuqrbK82a+J/Ixp0cc/UVKX5jwQSLV5rt8
yGfwa4qyC/P7qtGjkkJTo51nPYbt9OP5qEggVSc05Ex5swtaNObM9/0yA2mQDMYW
qVThIkqsJ59jGZNgrDniW0OeEtMvIhftHM72+hqUxZxVvs8/Tf/ppeP1xisWJ5lP
d1/3pSDuBxDLpSipkhM342xiipf2sZMxM4yRndiYTBw1uDUnnJL5WEV6eHTeODbD
QQO5XcUzw6YKXw667Alkmu2RTT1JpcyxHioLQYJlyEppfr4zUPLVvYwVaX+Kak/z
4ulY6AF+S8IyjiFsovgCJMW7aB4nzuE391+sHypSrSPRtRfWv42moxfNniVN9GL5
OCZc9/LhshcM7d4msSxLGQW2iD9ezsALLSj0eUMR780KqMZMAqPYvip8XPhd1RhR
b6BLO564VelP8ftTVugmXx7M0t3PaGmZljZzQucKMMwyeZ0KJ/TsZ5J+CDs6KRdZ
PMG2QnCQzcO5YRdEMYVcw5MAoqWBH7h2w7cVagXET2nM8dAla2uimy9V8IrwvNeX
cYKVVSuy1axk4NlCy2HqdACrPn9yCHzIl+MayYtnUNhNulQXa7vrfpg502OYxwvr
ipTWOPXfXSC+6zGbXWFI7+lmM0k/yZp8LHKauEhngT2PN/Rj/n/J8HLI/2IBsFC7
vMmgtjIXHnwAGGbHdB5QtsAzvSPNJpavhtpvtSuREfAiANCYhuYOd716YNivu40r
wLZwWE4804nhUqnKrGxCrPzB6eTmkMlNhyjvXHOD+Dp/aH7r27d8Y1Le26zM6gHG
RxDv0mkhEw3IEH8VjDLnasG4BmE6zqrN4R+8ReDPri++V3c+GE10xmAIlIqSe3c6
34escRNdL9MMTbUUjmo7K0bH/hD7Lw38hEfdcteawL/q07X51vQ5MGDp7g5fjQbf
GjvzcTm72vexCIqAgziXIXB8jn26f3GcaJ+MhCgqpG3t9+aYs8cNZ0/tOePB8uNf
15Uk7IzDkDZ7YRCQlTPtRhApQ0zNXZCnbYkfRtauZyi6d3p0gsfFpsdTA5gdHME7
f53eiaceFuU0NT3QcElXdlsXpNvrmpin9ThTPI0h5qqroxEzWj4e04HlCK+KLZVR
63dB3CgI+ImyENe2dCkbZ2LZ6To2zEcNjVmb9qWAI98Q5p3wFFJFkiSgQ7e9hYpj
9RRdfYOv2hqF9E5SntFmrCmFbsGieiPbGLR0e3DAV3+v/yXkH7QCcxeFJTpiFqNZ
pBs4YEgcYk5gilTqieW2Y/p9rdZfTK3SGQL74pfAr1gw+/8iIVSrvJ7jVSLXDeM6
W2y7XadLZwu6aq1LNhZoFFZERUxUfqoyaciSlP/254Y0gKzsXJY2IzknmDX07Lp5
tWTa7rkEIlx327Wntl9GhQ7cqwODNbb1aZByXEa8x/O+2XF4PgSfe0LkUsj0XIVe
kNhyAoGE4hzg/tPq9ty6sFnNOxnVkDlxvTK82ln8jpU0RbGPX5B5iN2DcJUx8643
jW1X/tW1RF4NxpMD9Wu3i83yXiBoRpvuN5glMIkC08EwxlSOaA8YaZjZXtGVAif0
45np8mUm6d3W9GjxBTfQR2A4rQuX6MtntoJ2X23NWVWLHBHyEc17Lbwhw3D23TBM
LCZMUnR6OT+a6902NBHHmjYn9nhgid/+tMZNyp7STw3FeabvbPMPdG5TbA/J5a6X
ptEPe+OP1SK7MM9y6LQcd6URm4c5IQ7IEvIKSamQSL/23O+bQg+o0VrDe1piT/tA
AVQ4rRC+5Ady9KsLqvcJM5CVqRdIwg63Z11wGpQn2dRmHiNJ4lmVcODNppuyekf1
n+hLG+de1DB3Ovac8BOYdQD4CpIHigjZCB+w7M1d1ZjhcjukFuM95KaWCU/8TgXn
bTYL+MNBbQdAZCO4hsBNz43SEM8TllOFqNIAcX9e+3FzXM8iPpSeiyPpiSeLY01H
szB1N4FI1kpQVeMs/K4dEJp+5WgafwvBQJdXKVULhX4uzS58gd9eBMKKX82rDylw
DbTiC65cEpOfCc4OQ9qvPBcxVSKfuFyHzD2MICTWCvOrAbS2/NhjZOF5UpBitpLJ
3F2uQFxKKPmjSEBUSKluQwQH6+QwNb609xkfrlwswJqQ1R3RGdkKsAiW6KgmTJgP
9GkQZkTdX5bgY38tFkVkNoTycSHS3At4rkp+8QvmTuR67QCqmAO0WwQUke4pkjbO
2jv92DU2cq7qLHMUcn1DtGsG+VOVcZGIvfA6WzRqNMkEv33fJVYB5Mfoz+MJ7osO
tIVKENUEX6PXTmY11KRplNVRtXvuPH9s5xuyX/aZykzcpiDJMZXfU4oft9YNj/ZY
dkUJgcWbPpslUipK/ZM4Sv8x2VvlHk1RAyvUPIxp9HyozaMrBqZ0J8vpJx4g7trn
9qnksX3/ZKaXmlS7VX6x3PYgToItPQpnzTOvK+Ayx86SedMVnALBxvKvT2JXUzP6
WURxlTE4i5JVMOxxwXOvj3hjavt25WY9oJeHgRBBB95bAGmVmimCIY0Q0hLlsAd0
1JhwXMnLg8tAk+xmQphOtEBf8P3zTPp5ga59Fc9TtpRec7H5CHqLm6eqGz2E9KSS
AcIWqAt5KeVXQULpFDzqXybcU8f+KLCG7+l+gk/YxenhWMkfKZ3Ui8YSQYrD3Fqg
Pa2lo7QOYFHyGsl6kukEsOBljR1FkZmrvvXdmtHnwFnTTNuBO8R7KftUg01GdRDV
FP6v+STM5aKldkpORdtzIWncuHv0spy8dTWs9Fnr7iBgA/F7rpz5Akjy7dRvI0Zk
cZh3TNGslG+viKuuJhHdilYTUQ0EHxfA2zz7IOfPikGo0rl3uQuYut9Mq7TPcJGH
01SxakPrJWnh3cZ+p0Zjn9xMVJ/KaxeHqJDD4vr8D7Igrym5WGndwXF4IAV4W7hy
9HzkAqTvLm2t8vlujdybtxYH4d8Hasz5UY5zHvvLH6lyI4tbu40rBLi0DWWIZMWU
K9tbFN5ADnRstgmaTrGk1DEw185GibFTSbIDu1VNr5mZLGXEXbNaX6cbdeYV92/2
S+6RySwwldbDeddZpHK1miW1byk4tazDioLHORt/s53Gv+GmKE4LL9KQOMXz7YRT
etqDGm/vZ5q6J4CSvyvcTMPCfu8Jv7ZWVAwnSa0iiQ74x+AfBmEwYA3gMwcNbSgN
04rnTmMtmlRZr8bCw9VZNv27/udpPVFYFKugHjJoKSkkr3OzG1cKWoaHiW2F6XuH
C1+fRIE2ptQb3923Vf9aG5HQZmN8t/oTIRiStpQPk5pvC5CXHZS05P7tbWB99z/c
05CXlBT4mweVIPEMpwHfoVkit6Uyf3ZUtJ81WrGmwVz5Z5Lm98GFilX00uXFukgS
MsnXKCOSexK0O8g4OHU/cr9A9qOo/N5HbTgm9T6xGRITPb+CH0R+FWUF0SbbdBpN
F0ZpQafh2X0w6ON0xfcbXyOVzwuc4e0A/QrsULAEz6GotDR0x1KNTpdsdM5+xco4
NLnjTSHfpeDJW2VdJVGWs8dIUho0ebuiLppuKgBPVc8NWUvIgGQAcakbjE1Q3L87
KGlyGskaG6qd0bQesHanWsPGwez46+6YujXQJyvuahs8QyfDNebZc67y4pHb4AgC
F7myP8Z0yjFYnpPMxQ9yT1RLuGRiX7BPWD06D+DJy8Jw6e2y2XbRKAHCDEPYYT6b
EIbe9BMisn7HW1kvNrHs7dD9bljk4ZpbeJDGz5LiD4xt5hSidCFaHnfoYka/fn1Q
pO6nFALEE+c3elCqUIPqrhBoV43NKMlakbh7ZLUMtEW+GBEyjJ9dIi+803/F2lTM
o3OKSuq4ijiBT0IJbUgoadYgp9YTU6YM4TJvi5K+2ee5VJ78pwbAcJSFgx5mI8V+
6teEsU/Fhrf1RCRA3JdWWCQvrJ7jwo4X2v23u5zOf38cMZhrO+uUsgf4foPxaI41
NZ38OLgel2HCZkeHJ1syqnSX5DFHvvpO+1vHaFQ3W5/MQDPNWHzk5VxUapTBXqo8
NgESyK0YChe8VJr20VbiUmUYxMRJ7hCy1bApNScypH86EO6/ffIvnspN751J+2a9
ndVJq9/m1+2ArqWifX+n41/Z7AANIvvBczQGV3S82jc5qMxXRuNAaacnkmr1QJ3f
wbOcZg8pxoeIbhPaWcbuuTURDafuo5RfcYIY+oec9//ubra/6AO4wzWCwI23l+ON
rC7j+nf+WPR5Xbm96rgxEgpJeCp+XcnZIJGKG8fPMJshhQEPlbXG5y9I7F067iHc
OE12PRz2Y8/8O5eqIEu6Ek2rqeAG/xoJ4FCq3ZAOA4W6T4JmxHRNSw7cGXo3vEt1
1X+Tq0mIj666UjO8EAAA9veLp/OXn8RBxKc4Apo1tCiUOfbe6bey54Ke6Y99sAag
uXdHdm9QcvuxM0zDX7UOluoJXRmtn2kLZFEYJm9utdq3nOJH6eJA9THvT9uGRXGY
1uMZrQgsD1hD5lB0fmhwsBA9Gt3dajqThnvJD4OkQq97PqXb4RHP4DTfuqFdo7/t
dRhDfFtHHhd0xcuJd7Aw6CXRPn9fW4PqqMdBD2mHrY2TvsMfbs5/+E6VzmElwIF6
sU5BixF6u0ETkTL0cjY0DVDShtwhet92jPc1sLz4WJuL165cCICi3Xsn8yOJXU6u
gNtm0CDvC7Lm5ck5tMSvArEw3In02vsx0iH+Vb2h29JvaqmBuRxkvf+AwDdJn9eE
9ogNHtMI6T8wS8AtjwK+owpPNOoUAdfx2KFQH5zPfkn4Q5m2+1MHTCa0MXdGE9RG
pWtLsJDQbZUastMsUQ0/Ewm1VYkfOWkW1Z08BYePoxC6iq2dvz637Y131aOa0aaC
3VuCJsE5RD3HhiJuIqALcbdC22JDDNTYCkYB+e9Urh2UjJO/8bH1heZ3JRNOBrK7
FwlGIpIo21AOSyNZGdfWJ6Ci49pdw09cYIgwXv1H/lMDwqoV6pFnJGGCSHmcnzwZ
sP9HAJOwAGdRDcfYcHx+B8AE+vHwITyp6tBgjqOws8BHEQbckXtOujHMoNcamQmQ
M1phY1hSImyv3MXnhYAUhSFloQVfa7Xi6pVVNwXSohqHp72s2Zxh1hYH1VZnSYMP
AECnrvRmLN8G8v5l7KFkQmlFMSUo+th7nOtE/3G/gTxO6Z3asCXM8NABO8K+Dxgp
f9r64TE74Z3+hO61KT6dfjHc+eRMVidSInoFt+JFLWmvDEzYWFhs2Skrw5Ydg/6K
M3PkaXGVq2+ZQ7LL9oiWP2XrdbOYifXan0uadnlAyqKnOf0T2IMJWs5YPr9PcnQS
mojFipRRnGRNU1W8v6+K6rKPDR1c+TrQURnu4d99Motw/AAx1Qs4sXs3OxYqpcSc
aUa0KaqjAHCO4o7/kpMnKFPRD/XhdV3W5SiOi7BKYrODU/SRVaD2Bj3cudIlohP/
H3jXfVK7AVq8bW9orB2EotuM+fiGbbEkPDyM+ANjvX9yJUj4Rf75iQwdVhjp/W19
1MLLeLAVgsvGOCWWpifo3hQZ15KaWY0COvTaBLwH5h0nEhSndPvamKu3lDYFLEMu
KG7b0N+EEPtZpKHHa7Dc3MmRhvdYjKppWjWsCbO1k6dufezht0YRa7aX770ReYSl
FavxQM0LIFbmL9nGtqzbYKg5IWFTIWe1ecghe6wJ7tU40draG/HPlZZdz22voAgH
A8RNOTxYqkeOAfTsgkRNkjrypcnL6j7/JIy8+2mOmFZD3ZZRdeMow2wDF1C2e2rL
oyYh4ZohRhPPqcM/iEnYL9BrvJ6wKgQ9lvfdAu8TE6LQuqhURiWmL/8zh02XrwPC
JiAneEC8J/mh9F17bqd7rhHFS4K8OdePyebDEbBaReZXqLw1KmDuE4taG3JlJbz2
YqOyeHABM5uRMc0fTe7zyGYpn2U84zWzRe5cREjQmG7R0jdz1JWB60nZC+jT2VDt
fu3cfOLXEcrpa0zV/Z/YMOc+rKHu8XcomNtkBQd1HXjO7XJ88fueeGMJ69wLDzTW
fv6yq1fl4VF6ms8Y/slwp6+qfF+4Ve1YXICHBTKspl72a1hiTVv8AUsM8HUCvcs8
iM9V4iADZg/tj4zXZvoQ7d+quxo25cNjFtbqyAhn2HxbBSxB/8My/WLtZgL7+nLg
uYZIPZCyiR4Zu7e/03Hl4b28OZQ8wl1EbSoLmuLZeRwedxmPek1xUIsVnwqSMC8j
sJzToTYNjWxJ7pQtSWrDskvz7t7fceCCM6Na5xhOjygjxUDmupbhlMtfoIUkR2Zw
mbQhpI5XY4AQBsp9/Z8HcK3IWcPuFzdlIJPARqwAOwT2SKrNKZ3l2veJ4yoyRr7g
ntRkOycE5fNGbNDu+8MlNMuPDpIOprJzzoDwrEcjlPWQQ8B0LXIFlGxho2ohwjGY
mciCryJkIelj9kg5Y5UVR/yTQNyA3LCaX8eZsXIF3dTN51N7MCCXHePJRdUw25NO
Gd91JfyDPIRUmPoay5U3ZV2Kn/DyyF9H/bRrQJ5HZ0G5GDed4zKd2Xe6u230IZXe
0IQgxdiyyR7EVKNbKB+m2SdIkw0dTd4Y4S9J0LHDU1O2cxBLaPNV2UrswT2oYPbw
RqE++phMBs8++y7l/3jxQwzV7SqH03+z/isQQ6KWJnpsMAsUp/JO/osYOWtV+Xz2
Ycoyd8xDqfsj7OrW8ZXRM4AWrpGXJpF1IFV7SUhX8F4tZwwoiR4QEuH92EQ+B+/v
6CzjoYWMDssmtRmBK2HBjONLFOK84N8lIBnsjPXmFhTgyJg0aEeE2Kx5zVDjlP3B
pr/M/YxBvnbTCrLzGn3WIRYG95JaVS396MP6XdwG+4pYfIfjn3qBRtG0ulanHn+u
BqaFuHgd5IY93MKBLcC9Pf2Y611MpyqqeCCu0jeIIhmOJNH7qpfab9TMXN19PayP
7OQ92OZZlIKmVBMtq8nsN/zF/QUkE/QJYGWRbZ/KwR46l9cbRWBgBB1SzGZqAky/
RZqrHw1Fl3XvP8x9Mv24b++lkDrOxw2RnMjm7FzNMzW0xHYd6WIKM9aElXw65M9L
iozGTyfgiB/M8MtxbfazodR8S6Ro/tp/1hoBvZk1dIRDt0vc21RUupzloessyMX3
0KUWtjgCuad8tAhqPqlRUxEqPeFrl5s9/4R8BElO+j08Ql0/ZI9lmbmf76r8N0lm
d116kbN5hqi85em9pkrq8iRIuES7GYakaz2FpMW/nNTAXYjqyB0ynCc6OXNTi2Y/
bW2Sivxdghx0Qle8TiqnWR2qSSOUGGWVFYO3VdD7EwE1ZpN0srtXWc14pJ/mdaro
5J9+qOqBSocXF93LwrpEyhusbdh60lFOioB8tXOxePlMYrYFWvjQlEJ1TlhuuPyz
4mljBANr8IcSIJEoxnx+LC0eGps/biQdhUcHzQUS/apFgz/udywn3lPxlrRhMZOG
w06yfQYVwmIxt5JBd2CQGB3Kk0LmWN9+0zqXRRyuwmVM9OrH1j//jtoQeBtTpqg8
TcPkXXy5ZZ59OCyAxiGaBAcVAUEjdQVz5SbywfVRHv49QOM05ScWrvYa0XCffal2
STQUy3RgNEiNfcqEReAl6H/DmHc41nKfqaPwrRVasRYqKrwgEwOK2eT9QM9zeIMC
bfnzfdWbu0g5O6F35CZNp8ayY3YQz1z5jJoVaCl7xOlXMXaDzyY00qqG60V5D5wS
6L3wEV3JFMazOAYcQvccBnAq3U5MknhiSGkdFXcgFYUr+mHriAWvm/F6asTfP6OM
NXWjfEgzT7A6jYY4PejjiMj1itciY4MzqSIs3ENJijjw1I++nsMlXqyPFy+uIfUV
HCK0x/PPLhDn0iMaZctha/yluPmUN++gFu756pRtfHPfmDWvOZo1B+0A7JRzyZnc
/wdxeh3XZGZwi4cce5VCVm65CL1UgNUL6OSjQl38pbbm6gwMASmBBil9CH1LIhgc
JJlCEpfxlr/Bl/Ysg/GxpHewgSDUSP4kceJSCPbmi3NxO6mJzalbWZPq517+Q+sG
GYlOvUpyW5esn9PlLY0xPvmwph9ajARlnjV0jN0J3ssDwhHTw1UNB/timP+mMqxL
FuVD+L/e8Qoc9kaBE/oM+kRTSlB9G0GFI5EmNlZ9tuj5NnsCKA/+UmogTlJ192bw
+VCXQpokKq6nj+lG1QnqaPMxV1GTHULZEhFv3+HAVnQnmFRYbscqLza1VRjEQy1N
9IdQB5HQEId/8QpsSSIdbAM90yBW3Grt6K1qPebcOzgLBMNa/C1JBh4exkhU2VCC
eUdW7Psd0xxaCxRwyZiiKsX4DXfbQEBy/5QwZZ0wH+zTYn5s9Brh4Yc+3nEtkq1E
iF/TwMH7GR6fGsknWc10KjvXeOCDYaqm7a+rJN2LpwjdkxpqhPiWqgCqsCfbo6mC
wKfItRm1egnC/lmP4RXd0DXaLVaONJheEgWpAXxvZE1SO+sCBoO2IQ7/X+hXcCfS
9i/PDwP2dflmOPjQTJhsYHR6VS/z7rxYxkYJZV1O4QhyeILNEQlPAbyxYaVXJcUm
THaoiC7ngT1GrHdVFDYKMPOU1nuuehNN8v0zYCpbNNcGn0q9VJR+INykKmVRmzPu
E1RNUx1UE4XPET7rUPlH+ogihxEz4+KXK0WKV05mRul1Tq5/AWt7bC7Ap7p2lLcU
VoFFuqk2ZzfTQt0ncxE6/gJMnbxig9OBMXjQ8dYlmxdnhE+ZXLyqFH3/p1zIMVvr
iwLfQ1tsPii6i+R5/7X+8xBBqjh6c4duzrffptT9renGZMJ2CZSLmuZBAwqfUVNP
qfOTOReP7R4f0cqveXq7vQoyH83oyVIEmwqKXaQU4ii79LDp7WiczWkayGuDRQON
cIwUZ9I0Rh0clOKTqZvq5sPwxaufk04x6V57cH8MlutqEBfiBPzB48AAfT4oo1/b
KNEz/gQZ/PPvzp+cSBoMDwYaqZ+c87PGVEQ8fYd27Tw8yEtSuVHsvBkWe1jYz6yf
yn4Vn4nw+MHVvENZ+rWa0dw4VSGcKYfs9fsX9YpsPbui2NMcriX2qQvc25bruNkD
16S2V7B1itHYyaQwPb+UpWcer+HlQ7ccaLCCFBXXVbfumtR6NcTrb6Nucp+BWc5W
wfT6ZAK/oNFZDONocJ3t2M48ljdSgR0gTtp4mT2TL8V+enxNhhz5vH1ljvaRa6Ac
5ehvrizV5nQJ5r1410ocYgqdWFk/G5fapgK0da/Zf0XQ/9W+OCxH57m2GAXyFrK4
vM/yvVho4/6bzoIFFK6DdwnV63A7dju/CTLH6AUEgXJc2pz1sxpmVqwdhc0eudjP
5DB5y9aixDZiWasQ3bjU7my5utiH+W0z+gRLfk9tpyr9CMqF+KwHdV1YOQNFs5Ra
AYXjiyOIuQbqWUnCp/IvmLdPFCHU9qB2tkb4lLkbNvJUbK5MAlb07LLToprIfkQ4
z5nYJtERKN/eKN0riRB8Q/QGE85cofGPwktrfH8F8gkFdy4IthsGZCuv+5s3xHDi
4O/0/A73eWdYZHRQogyldM2gD1z6tQsg1ZJJwmicr89YjET/frklAjOYDZADl3LE
eF54xFAj8fO81BX82N1b8te5K5uKeiDQP53alEdg9E4/nA2N/ni4kFIb0Fc40nUj
8Uzz89pnqpwb5JHAazPtxrywiCltc2G67R7ctb71ORBX7vuIHWA5kKoSHUBSOzjR
JUd504eEDbW1BF82HmsslDw0yqHgGyjKNiMJonIN3AN1CjLM4dXYHmW0BX3jfmTY
l+EyFneE/+TxSIIGLMaxV0OHpIPw+/QepTHDl32aBKVs4zduv8lMtza8qxY5UOvE
YRg8geN9hq+WiEMIIHbLrkKc2WkB/yyCu321Dhy1Vxw5eHHcUbpTfO8PAKOywvey
fQxiJZTO3KI5fEx16dZ8PAzfBzFgwL9LXmt9wV8ef819jE0eTapvgYqL5HmiUMVf
FXUn0wKIwhB6zzLyMSPX2Zc9mYxYh6pQcLYk0Eh5OkV92S1qtU1Qkug9vqLVnC1Z
l0b2FJcDZX3Nnr+TOT4yXTdtwLCryj/wfBUKicnyUlXNhoKGfKRLG5dSTQsJo/WW
bPYnkF4XMIbHX5+p0Re4VDqXxiG3OFVtrOb3ouYdJPcU6gAhDQPOz0UB9iukPlPR
+rWyvTBCQ66rWUyXbohwkdrcE8UAQGpOXjl4trNjx0H4MepRS7O3tqyA/TJCbMYB
nZQ6y6CsAoiBhdBKJTMLMQPi+FrCQ47k76Ss/8FRVQPu5zE7WJ+CCflHZzL3OT83
Tqv3WOd0WAlKyd9CC7iW8pOYzXuIcBk8wlyX7M14auGV1/HG5TdpAhrRmoqOGiYQ
0GMs6FK3urQEIiTw8MyRyWXFNE7p4aFrudYfqd2/jSCqI0k0PR8fp5UNt+K8OoqP
JowZ9eDE2CzfU0letMVsSgRg+g9MfShlQZY4yJt5x/aW6l143Rkrv0or4EAfZ5wG
qk82HRDWk+7dpo9ViOM1avTaKGBJy1efT9memvJtcGh9yJOt8gyAa8WJsjsyGRf+
mVskj4xp1NkIGY3blBwxBUD7FEgetontsuI0ODcLj8CODPgXed6FROwOYZSn2B4w
rBSAPync6NBLKhd0uBXb2AebBW9uwkiKIAS5nhPRqiuQzeAi6epK4yx3MFFDA+iU
D0eCTW57Wc/xAzZeaaSp/9hmwVTuqQg3Ta1zT5AgR6qCYH1QNrQkTKXM75+R76GH
tLJB8szKKqeoUtvGJxCzeaWiJ9ljz8dOQlZSF8n5NW8UIsqIFTFv9Z4FT6wvn3T8
pLMYgxom/Br451RcN6m9m9ZEtHUucZjwy+Xot8OLViexHu6C+BXO4NV1uslTFciE
VeY7FulK2jIb8Wp9y/d1990IPRqQdzRAWSHDD7UQzYzjRpfAQAr/rt6a8xhdvK5P
ayLSWcx47QdhDzmFDRVVg/DZcPJQltwEd4f8hiW1TaMU2X8n3FpJVKXk/dnItOXD
uTEJ24aUbbxBI6MoMxCw8XxOcBop1HAxjLQn/O/nGGFgZTW/reCQH+HsJaltCp2H
eBpigcb3O1adlBXYjMguY1Ar0E4q7q7qrRDzcHK0+Y/GtXOT/ODpKnhBwjdEOYfq
R0wYS/A7uXq4BRD957K9ZShUq6kaYHpFvqj6l3EkmqW0+a9s+ysP3UVoTB9DroB3
0CRQ8v18Jj6aXlNDbpFIUfRZ2UkwxSII7ytjMs22MZT13tsi4Fj67c7b3zVsftW8
tksNzPPZl6YRBMGzbgmXL/qo0Pv1jOv++WTehtkAuuSzryBvpmH9rfz6EGAMAGbT
k1j8yYitj/nB4hWk3c2ObWq1/r+ienwvfXpKVOdkhfGS6/50LeqxflDa+z8vm6fR
vl55Uf+Z9X1AI9ez5J6gaK5AQIwn0eAFDI4K/KW5IRpHVQwhuEE93UDwZlYLXwP7
z53BsnE2CFjuJkheTiJsKujEQMy/HagrYp3h4APLve6UoB8/PQa2k7N/oJEJ/9oC
Ke3rwkDiOVGrkJmIQwfUwCDQFQSQ6grjlqmlJMzyDMTzVX5U9RgkFOPU4mhPI5Gs
/OfQ9nHVLsOirMUaTPlCpzpe7Z3zlqBpdhrmycRxaunTaAxPe9PVtxuUt3hO49Wf
3DtEe4S/2lO0uKe0EMS4sMXVy8UOS9ewEaalJk5mrCPrcfH773A9dlfv1NewMLFY
tfpn2CqyJzpP6w/9xsLgwcvQh0MvqL7c3VeDTAn8jKNw+0PGnALYIPUUDiN1PCFp
q5W3tPxr7kfFgb4GTxePL0ZvziuBbuRL2or8v6qOPqb0b8XvWskfwUKsHiRRiTnU
/vVQFjSqXVHvbpnQBI7wo/AZmp9gY/RAusFvZOf8V29Koo8j0+d+L6m++g5yP3/w
Z2OpiSdjNLPUMDp0qvwMAc1KhwjHLUJ78gpSCB9EdjqSDLQuJsazL7w8C25HF5SN
XplajgFHKG3IC/3LxV+aXudAvjGLShjIWV+sk2F0UZO1YoBKTfUMNCZmBarWdYjX
T0cPxY5nAVwMTn4ibojQjk9eDS4J8IxINK+66gyAMV5/1Z+Vl1DP+1Gcbu/71wiM
IkDlScWx5ad5maDqEuyajWZ+4IXjaWUlPkrNgA9clpopScLNDeeE/TDUMnDYsqBk
RLrTkWyDT2XdLvAIq6smBm6XMmksZ7R8n9pwshY2xM1G/4B9sWxHlEdLQ3F96CTd
8XvvcNKdELog2HbJ3Xd0hfpefkPElx6x/4etFfh0BHwH3c2TwPicDqNb4eAax44y
USULt/zsWeskjMkY6ZhIxx6A5YrMHRhB67I9sCpeLy3WqC9mU83oK/5GmwBsi15z
mV7P55xtpjYrd0J1JUOtlN3Rkx8Otato1rXrjdAqbS8eMwfXE3AkBL+NbAKPIVPW
yaNNiU7S5RJYP3GHDS6mqAmLvhZINJDmBlvzY4JsU+HZaruX86zG4L3mmR4MwPYd
5ueTCcSgQEJ/EdEP2f8WYPMwRMB68ZyT06Z8N9N1GQrFvMG1WFISgyKNHZ236YlJ
UtI+BOtyOkB7XOyyUx0vgH4IynZIMEFLUVV6L+oC4eLwkFZmnRlAhaRwe/UAvAOK
Z0x1ZfK1IyQ4wg0jdkhovqonZkmYVsXfdp7wxmQ1un3nRe0J3KXJcgNVSt1Lmoyb
k2495K8f5XIJRhH+2F1e9SPCxQlnHC5w+mlBkjCo61s+fyXk+qr4nr5iyfXypP8O
2ardA1EXP/ze57elH0hk2jabB0K1yVXu73OiiScDvLmdJ8Km9BcTzVqIldXgLu8s
NjqVegNCbIZSYec6IM6VkXzrfzacLWmaWn8r05YTmpgVvebjrspyuoJFjJk4KtHf
cxns7RhX5NxqWjMs9nvkOZtsTdE5R+9A1IZ09Qxf331bTxkU3ob5h5Y33Zl4hOvG
/ZFuO1TfoVTTtw5ki1asuh3/F448k2frc66Ah+jN3Bl6KzulsRLZaLU2NJvWYiXN
bxKylx+DipEdou2W/iT/aV8DOZDTwFyz4ZEe3FNIeeNxhh4lBB9tH99T7V/UXNIv
P8XvCbZR8QvrgObXzqrD5sKnwWZqY4cfCoC6bQBVnO4MLkVGKxDNYjw7rc/CV4mi
YUifderz24KxqsXmtDIHX7+/k973281waGLznmmDZeUu49jmMXgJCT35BvhBDI2R
UVXJT8ujCDePaUxnc6q2ScRE0lhu9Zfq6wQeM4oYSzQiAqcco49g6heSXUTXgBUN
2n+Ly/LOz+Aqruo+Rq2RumXBSLd0BeNBUFKwXyFEBDmjsLEPwsyPwwgjWEG22zx5
TGzopj7yvLlKRgl/PrttokMa29bzBREimoz4CtvjqDx8wE2USby6TytGkV2khGdW
FQPDbxoqqkQfm+EHCzOwLTHEl2KlDdXDR1Og27vqn5LMLBCik5qQ3Z5BKTg5zLDr
SxfqEwc0pzEFctXOGBy8XZ6dDNi0bTAUyzKcVWZ2KtBd4jkPJUVSfgQjwijAuSbG
wRw3fVH6BNU6d+cC4RN+uKHmiBmgdcXdHkHPbWbEFWxKkpIuuldhfDn3UehufDI3
Ax36jS63DX0DxGLxG5zAROKt5Msy5ygoN2E80yJdwmO686ZiF+ME1lFD5p8lcC2y
s1wNFCA3KafO7wo/TaJ3n4Ct2AmVJnq1LPjtyvqVZgniWXU9cvjW2wjQCdP22aoa
f2iykCJM8jyP9NbxHFSAVj0zABabpEJMghuic+76uEXyeOLbaRxXEm+ztiTwnOc4
fwbaMeP8yJg4Nqobvkm/Jw2K9LQWpWrOg7JLBqBLfQzi4RZzFZ7pP7+Sp33pahGO
FlGeHaLUyiA+JQi68YnFnxVIDoX88IHTs2klzlXLeKk9Hq4DfIjskVI5cIYYhyyi
iVaakrI8b9wguO0bpxVUroaN0d9ubYykLPwdO5uWVNBfcIGiXSNFPsvXZYSmxLs2
rXGVaGdOTZt6Gx30ytTHMwezaxvARSlagTLoUI/6nxYrh7BXOBc3NoBVWzej+rLW
eCwmqsfvK3nW+0CQ+RtPsrmjKyg9z5uM33w+jhwKazK9wRPS5XrCUUn2kUBq1S2n
VfPGgNjN/pqAh1QBPD1BArsysLS3F0RvlaZU6ZK3MZiYTiu/cjrKh20wUTIIG5ux
OWVUUU65Ism25rePr5iHwQkypmBv0Fp78UgY2PLPc35DX16eDfL5rY6XAdrpwipW
Pa8q7isXjRe1fzOIOxLSYd84tZfUyh8N0SXynnvU3eggnhxWlmWicVIwpG7KgFz+
T5W/1OrpUzdJDnBd+T+CPeJ3xTwvaNOepCW0PB0/1ymgtIKFukwahYFuIohJxf3r
T7+Ua4pTYwfZRF6GLprWiDpQ4sk+MgCViFQynq/kXkpk7UCVYIGhzIW2C5Pk+jSA
CX5muP1BVv2NfY2llXsOsXTDUQ1hMBhnAhRHOu4s06C6PeoRZ3GFokRun5FWJpZ6
ftcUPL5fiLpSwsbsYfGJSeQV79KldxcG5YldMRFYT6OIry0qEw7cnTfOOND8yD3D
MNSOGZ3jHuVqtTtHrOjfGCaz+ti7qL3FmuCqRMm9+Xkbh2Ur6FTij5xx6Iu/3+Jv
TOfHEzqLkrb8oMWuIYACFDed8k+xARQeW9tJ1Y1cjJYY8wlxuvQ2qk1Y9J7/onHS
dsgFjm2bcveLZFqcBipMAPT7Dh+cIi42xPYSW/BP5AnKL0PSfJidHTJT1T3QKWql
mbZI6vJM+mUI6UPTi2AeGsUPI2gOVM9/jobmRofpgtRXnblfuTBRgU+8gBm+/NIK
HG32Exi8Z3VtwlaL+lr6mnIMn4bW/oFGYTsXWSdq4RXGhlJpeHZtYClNHVs0rEn2
8FpTKrqTgbu0sVvD0b5f3ckCirkYMOeXEOjz95qtGhm3BgJOE11OgEzagmumtUuC
/icRU8UXoY0GLpcxe9am0Zhf9k6CZDSwNf6f9rN1M481sR4HHOh54GBFtHNrpn3/
SnzgOv1cAs30zASDIW/treDxP9fyxRxJwxNy1OkQTdl9IIOrKdl/pcGDFjhubYNo
852x7BpJhQJXkzeq5ekZFxShNjM1EW0denpnHFKHMyoYLXhMyz0fGZQ/LuxWcnwi
Q/PiRSvTOeLpcKmGbnalmL8hwKYAMi3t/NsIV6waoDxcGBOqWkq4DNMFkBQpEjMW
sgaFFTQs1K9tCZ1K3IMkKj5z3stloF4orUZaDcwr6leZUaiR68OWpUnKFdWPTsmh
7ntdwhpy917I5LCnTJ3Oa792P+MMrNCrhN8rBOb7XHp5d71L0VRfc31io+UYXrXK
i8Ba8c2vKueJLxOh13RF8Luuv6LcVHIV8AOQ0eiZ6WEY59F2RhJcWfNdYDLEaenR
FBMFYafNxKVeLlXDSAHKXw7N6TvkwjNrf8W4YQWlfno3g3MhLIcLnqv7G48n6V6L
YHScgyXbr6rzV8gBATmw8CS2XKnQSbOd71j0WYF0ZC8Hx9prEh6ahzygBALbd7ZC
uLF/Jmq3MaAptpKwx5pVs6G1VMMgQcDAIe1wI7BrHehiEqmAl4IUg/L21L5OVkQj
83ZKqS0LmOOkars20HVlph63k9BktrVbamw2d9bnb3i7wI58Nc9WeS6LRQvlgeIu
W2UGRjroMI6fbHIM89BHKRcylDeYRMDnLLG1eqPXmWXjk6CHTMZQUZMeXWqICRrE
58xHfrjyoZeGPa/GWvBjR2Bm+Io7kTSoY6GydEp8gppLq57J5rGtQOr4QMxLKmTB
f+SLWiPVrRFipi+G0OnmTsq7mcZFrYFOuIhswtf5aLLr0gD5yGNlgsrB5IZ0kKaX
nQ8gB3NkN8JVWLHbPs1o+EBOQH6CQlZKIytkINIK1U2VJxf69gDO9djXUitogENk
y+mIcp8byHGIkKa7FGDDWTad8vLzhixMrjnTblIvv8e6skh+EWqQ3J2kMLyY5VLg
sdNCvQIP8o3ZX1ocyvjdCKEawBwnXyo3W6nbAJW0zQbN1oBBSnx6q7Jh5H0n5Qz0
3ZDihceAdsBqOso/Gc5vlWIOfA4CX0lOMqOYC/YeGKT6JTJGpTSclC5oC/yl7jzy
afBdtuA0WZddHj3uKL6NFjM1Zw/6yt/8uAL4gzjneLH68gLHwY869nmIS5i8w0b7
nfma88vmTLbiSVpnraR4TjEnJHrmKv+EpuiJBvYQwxmBG7+yzTJNY//yUnhfcuTY
b0wqZcHFeBKhcl6G1iC+RenDHbcHkK8gke+jcesxiNe4ilAnBH48UxzmAQf4TaKD
QFbuGA8CC5rjXM81cudLawlDO1jbDrKKr0hWHZG1gh+nhXvZjZkGOTfMLqAkP8+e
UepF8Y5wgvcEfgDl3UTv8WVaGqSX6JTIxP9PIQk5f3E5tuxOjrLDlaeitER31Iof
u5R5m1/gNcuZNjkc5iiAZeyor92BvbN+U0fVUv/kn5fjP1a89SHM31wHGbl/uLyL
s73wKbyb+WR63cYLp5049ORg7iEiRn4rBLm8Gx4zROTotZia+an8gpKX0UxBwqXW
U3HXVirX783ccf2yDO7PrZV/y4sy8QpjfLaCzoQaVjV3NAma8s8wgCHGprsWP9nW
fi2klTPriKdJP02nO85kngHHGeThbJaWoWKSdVFTGDu3NpSKzTg8A/3YKzxwMq/V
+vHbdG5VceAAlEYovOnItmfW84iJcpIKnZBrWr4pqIXA000AIN6KxT/Di4/+ehqb
GRwfMLfYqWVQWiF9gYX40s8EtgONMzFxJht0B2FK0JE5Skl73EFvXNz/HvYXUPTu
O7H5sd2YeGwyy3K8XrOn0XQmC7EGdleA9jirE1y4Np1yWFx7GL6MXElUXysch6Gj
t6lLnSVoWVfnkYnHONA0ll39jK8hh5HV8O0GYUOOV8KiGWM08boqWq5BVck1RA7u
lLxEt08rlUCi0Qqn3JTzgWhWvCte1CrC3xVHOnpYAA1vIZlYXYL6Z4pVEXlFM4h3
dx0haixOILKoS/D9cjo94BIA86T/yfSqwbVhqV9R4bYQA8u05w/yZowu6NYzIDrc
atkmV//CkK9pdu/gZwuuiMBLx+IMz0UUJXcKwnNHCZtr9oMhRsf3t9Y9dk5l9Y1h
Odh8+vvbXrSXF9rarGb7N7FfaZ/I1JSM320AvHhp6o3BHEdFoQov00bUqZPJIaJJ
YPWBUSF9BI+DvvJc51ZSIzpN6OiABGRiu4DzHMPW2TCPzPirh03U557T/FGGAjYf
yLNp30+SCNrUUct9tEJyzQG+NYw+12+vDBcrWc49hCdVPAGfUliK9ZTXS5o0BvgH
ji1gdlm6zwNEAPAi8vYyBzhPQ5Ep6Jd0sZ+1QhqKnfGWCrLaaxtk0/G7vVBK2JN2
09g1mNmBQRo73udUZT3nMvclQIZGJCK79vcXDZBgnHY6GWDyqAuiHysNHMlps1Kz
d+aIvO/b+HJZ9va/A24c9ovLlEGewnXUn8VVqDsEzkYaSGyO0TzYRZouziG3oQ3Z
4fpAAlcickYXSB8Ssu+oH6utWvSSFwR1hpRilWREUj5s989FA0+/SAH+i5QNYUXI
1XEUaBQEk8zK3XY17GSTkcVk2yK9oWeI6x31CGajhx3cmq7pJ9P2+fW+Me7jdAGp
sCFOt/js7DRXQ+V9ul/wP7gicYQX8HnBwDxtqi2ysg0HV3eu2JgVmB+bZPmVVUwj
fFGLdtdtztnnIhpQjhFW0ZoZRon/7J6CkNV//IMBv+2Gxqnu5kElyCf7ZbypfEQc
kEIEBuliyFeHMlM78mMrr6YbFl5TOuxvJfDATLxXvMbFecmOPszNTY51XnWlYU97
K9cpO+7hMx0i2V1lo1aU1UbZGdUnp1ps3ud3MLO5VlmYMmvENXsXRyuESRN5LuJV
NPU/aqlmq9XQMTtw1BvSBwcKAMpkULe5dgRzyhJ5w7wI5jAWC5Y+23bPRKsoeEGv
NX6DxBAVEQqWnvYBDkE9SCJlj6/A/XoTRmi9kiiIOaxlCk1a7JcGLbOza1PQC8yP
hR9az9Y42hQk2/UsPxMqGFAaEsBT7y11OSnRUWEvhfa4ncwPYxicu7XS31j7OTlW
Q02NbZKRft/xuc3RCHkzB6Dk1cMem7cMe6PhfLDajY7VFJgcZGl13ULOVUI1zX6i
fsy4h1FI2dOlFpjB13F2UitZN+sHhC6MW0e8m5wYo7nXY74OwGZgUvgyT0Lt999i
7iNu18zak4sy3/ZCJC1NhLZiCSS+l5bmP4tDN6XZX8uMypL6k1nEOmnpEs7pH91T
QU3LGJHiZgMEMRVbQmjSdXC5xkBT/91y9YJrGc88Gg0XNiwi7dMaAIDWBvD/rzeB
zjzzbGChDMc1I+NqIJr1hFya1HMBPg1TGNHLgcaXcYM4+KCnWQUbSj/CURR3adrv
oS4miGmhCNCZKT6s0I5XLBT/+W6dtsLCCMVGmpBhuQICHgF1Ehda4VfDQkNSmmNj
PBN7SX7ge/7kCIgzGJtGrp/ID2oKymyUQfyMYZ/q8GM2vNduJXeymHO6tLcQT0zF
3U44lQDCs5373/OKXg+43rT+21h5e2L41w0Bj5K/TQJNBYUl5V/2/UQXg0jMKwMr
/xf4xwQMiy+OKYFsPRzbLvR/nDma3HiaMVTwhV43B5cKbpQpbdHHldvU0LdxwBwA
0Si4wNOc6KBPzHUdeOFNjLGIuNyS6Wo1Izewc1sPHPp7vahAS8xsuo4wXwtGl839
PVb7/sBQV2N6V3Sf0yDegkB1T/XF/r8iHmFOUUOzmdlgmyxSPY+HThsOk8UBGcem
RXvdUkzR95ArIeNNLhT6IYp5M1/ad6MQVHX+2R6iYGZj26rxiG8PlsSFoL6k+1Gw
rdHpGk7kP1v104VZYTQRW2sox3FYfRF8eIK7tcIcqh3FeGiGoWydmLpZxs7oPHAP
I2ZboYyueuhJKA0q9fg7ekilmzkWo5uopvZYGJutpeaXXrrteQqkJdh7gOZlIsaW
/Guzr9K3CFjQZrC/yjcLGRs0nKTSodcaSOoQwEB0pN07PDKOB0qXoEu8qteGEumO
RhWn0CLNDoyZceJPt6FOgmWHC4pwDpLay5AiBwkZk9xKfcO7218run42jfwkRQRD
COespff0xcXcnxPwsyQUyNOWum2cmPZzPQny/3U1XV9m5ul9F7kuE8FWi+eHzqEq
r0xVT+umS5k9Z2CTOBY9fAKzJ+VkafV2Sd3PEf9pc3YMKZ4QrMC3XPguSuQRiUN9
Mn6FdQHQVz5uxFUE/WlO+vl5X7ebosIksYwa/p1Ay+8xDHuCU5aT+yb8gXhy/IOA
ZeiIJXrU2aDn1voknMkF7EVVi2WRKSsiSSTzfiXEJJ2X3KgZsM7QBPQLOR9+2cfX
4xNmxNcRGOUB5SKjVizk2Olqq2+YRHRuvhdoJYTLVmWlCerJaAL6LWTSEF1B7O8e
buHCeWwOnYMnQOOeuS7uKFALaWVYJd72AisYoj5XXLl2IxYClVzyoMmAcFdSQsaU
yM7sV6dcbyBupBT293kEruLaqQMEK3SCKTBGIWXaei9yi7z7e59vanGnVB5kDNLN
RBW8A//8PMJZmS6k7FLwwWYoH4UwF1TLVSgQUoY6ksB/NyFiO3PhxI0PmqsgrZAj
FpuOuYMJ+wHHpamA6XAERqHyumodo+9zRD0TMW404H46FvXf680PTJQ/apbT4xko
kRgknIiqqxh0uK15lqtghn6aVhfrc5+6EKsEhhRt4IjtbipGR/kqpoKwGh8ek3fx
b3uPjjkzFHClDaO0BBXjxYekWUMb2jWrmZp+RMq789yuK1Cw+Zitv4ve2SePtJNs
BwDjsrvOnFMzUP9EEsWj7l4boToWsvS3tmU6eiQuM0qDeYYgFRY/hnNMMrjJjj2h
/au+H0kqiAIb43YGXAnBjviGWHVGjX55HQ2xYo5cnK5m8y33SKWPi7judjQ30AJY
oOS3pP4hAYzfGjYsJrYA9n6JZ9zvCcWoD1qHNJgPCA747nJ4x1gwdc6gPYVRi47P
NXjiouH4EGGnTju0dbxV6tNQ2A6bmBbrV1e+5RDZR9PACny6Hp43MbYqkdRYVarT
TMarZkTBe4FC//n//ZBupK+tOqIKptndAuBCUIZNa169OAhTRMJRqTh9gBQeblWd
Xc1DbRvw/5VpdX8wRRv5vMUB3saqEQdr2c+0HzWT4fMTllIKhdDrZY1d23lYh/Jj
QrH0RKP9cCseBotcvDyHzdIdT8rLmir90/9nO7Hlr004Hl7i65+I2k4uQY3WrCV0
ZwZ85WSWl+C6nE5mv4zonZcZr+dcmOFmqZbbZ7Og+6/TF+/LKydiLWKxXr40EnFu
XvkPCjG2J6EgndsJwA+bJG5DMzyiOy+R03fuhxSGX6bMqpIaQmmz5Je+tNvP+ULW
Yjr4F83yxY9+dCmQ/C7ztw70DbWlwEykirpBK+3rbTigwZuZDXEQWopBESIw/URB
q///u2sQWWc6rb/A2M3ZKsJlFW3lILUM0PcSFGr+YeIj67b2CUBASVvMMB/QTyME
ERyiMM0Jq7kR9lI5WOVb1yjt4KmNIELgh5awMWFR0pLmkWMo5n9/C+vZNWamaa/F
8ayh9WPujw3T0E0OLQVpK8X39FE9iPDdSjnSQqyYuu6oB/7/VqiB4O5AllWgfyEg
W80Qdo1VXERlDUcgn/tf3NQH+QE4HtwBf0JbS1rSZplR+MzMXngpvMx81nOl1Ltt
LF/fIY8mElSPwiPUBR79F7wZTHy1Phc0TdB4DfsHxLXvkzmgH6D5/JeKKr09Lvm5
u8qIrG+YIrAff6+4lm9c4dIGad4qlMb2pxCNQN9L5qqMm/RLyS6+gM35dPXCvZ51
GE7op4JL9nvJLKHSeFqCx04AvPV4FU4txpsfTLd+kaKKJZd5FI/Y79V4UWHlY7cg
TRwrsiAxUqVVegR2egtwxrCZOAzKb+ZMEACxi3+EV2fo1UAW4wlol4LCg0X29b5d
wY/3ddZzQbHfatoJe4RV9l5Zgim9CcJfar/sFJz5e8DWXF055/GYaspf+30DhxbD
Sv+eWXlzKLL+zF0/MQ/VLqH8F4b+1v6jhiAmn/jGgCbmZP+0P2PYWio89b/jGVE4
l9oBg0EiAlYHj6GRjunjFv834VM8gx1YLpAgVvx7qD0+nxBR2KPX+l+DC4wzpHbP
uHaHwcumQJWvGNUDCdNNzEIARcPlKsBVGfYrOVgjBagYGEuJzWEbh3wCqeNHwjSH
7pcLoAsAQrgkUrj5ybsP95/9wgmDos9LagSu99kJMVPKvhsm6C2Y3AB/zF5uolkN
0U9jpUCw5SWEbUUc+agS5nsCBPDrHwZlVGGTrdzzedmoIUFQlRsXTUpdg4uzHn8r
8S+bPP1wfZ9EgYLZFs8H7TEbETM3NRBUcBtAAuANlvCO/3q7aC9iX+PCjkK1yrS1
GFgIW5byggjjSV+dTuV53jvvbWJ4FDaraI3A2UdhdK3NhlJbrA1WSgzMQTbmRmZQ
Selc1lf05erb5GCOkpkTH01aY3MBb7ylNHOl6PTXAgpXz3lJJg/hc7o/S13KM20v
CmVHOmYYEVx0eXtOSZdtFLGYLcdhsGkUtltADH7AkGdEnxatBHtXiEFZtxyD7tZ7
ydMS52ATQkr/fDyqDoO/FwJ7nc0pyH5L5o+nyjsqQa3hM6ZuQmC64bMSneEoUJpu
W0GM+hPMlnTqt+OH1/QLB71dMRbRc94Qnj1ZzKmR2NEucq31BdAXUbn/wudMvnBb
6WLK4QwahCIHvyTM/Qlo9yOCDCHZtgKWdQzGwu2rhZzI22Cj+tTTGbIwUS0z2Otu
g0sPhMVW/zh+j1YgvF4eEx2x7NbNpHfHVlnd0Ma5WzcQGYPgismHte/rghJ4PoLt
X9E5hXBY4x5du6WlC3vy8ywdg16sWzHOgZI8nKew0kcfUs0vOmLe7YCrzT1hM/L7
fGPw48h1V2GP6PWdgX2VqxD6t9F3/zE4/KMf0YeXOfdOLpZcBq+y+zeuo4Vt62zb
ePQYf+yQG1Ota4V9GRtrUmf4gtDaixvbWbJJS1dDQEnY994MsltgKxQI45WzaVFu
Aczd/7xbxNYVEmaAuDrMpkDfrAUJ4PYVsN5o2enWkGLti9utX7rQBeiUJqxznh5r
rlXwsqtWu8MFOd7BoiRnHIU+o76c8RFeM54/hrJe23h49/D9z0zmbb41MFJyrlyM
9CrVPVFoAmPpLOSQjaz4xthOKtIW32DCUPx2THQOdfBvN1Iw49TYQKRN3dqCFPke
XPOwPihoIR5zNZ3h77PHvUDJ5ex+C5C3vt7k2OImy1bHA1WoJNSTJkOAUKKUYwAH
5otDjipTh5qkA7/XuzTRDQAE5uXtvYxaYwAp0tv5wyHu1duNcI4yUhfBPZALvoUd
k38/iTOvxHJgKdNkP/wrhx7UsmfzLoQin3g9BpTvcYQN8CFCQLMXE/w6KWD5ybjy
3Yx0e//HEJsCIrCH4dt5mmX1lZFEtjqQcLwwbI71xMTmiMrl3QkBRJhckeSGyc2Z
fdSk3fMYLNaXVaiZaeWscTXFMJunGsu+bERmiLtq4ckvEjPLGsygE6u9I7QzB9TA
5KcyNz5sa5st4K+mdffwYgaIsGFsjZvI8586YlbT7g7QxLqA0FAZm6B4PeyMJOUj
kDi+75Y9+s2dc4jAQNhaaxiY8wGueUCGqT6otI9JJQWzDb+VXmufn2d0gxBjyCo8
69ppkNMRfS7fcDRLxw2waaPve5p6rL3l/T2cVD2kiy4jpyMmXVQ7p316Kz+hXaQg
QbPv1JHF562PKMGyIITD2RxuGMm6naEyQI4sG4+Dt3gRm24gdIswJSWeQLSfjZmU
ygpyCKPpaRqLJFVZ4HLkeNTTp3kEMxEQJGNBQyKvrEO2Yp42fUMGhuYuuw/AHBVz
nmw/bWTwoI7001rxi4whkjvTXgIXsLzYxyPHA6vdpu+b+PmHoV8uf2E5n6xIs9sz
BZyDn1ozk47Krkc/LnXVUlg2b+0zY423bTbujyuvEh8KBH1KK7lh0KB6FlYLbNgp
QcOSUxkvav752YHzprRXbtkQ/um5CFtl7kUobxGXhebZLBu/3sTx3YbDyLTwPv6v
EK4vcEMS7rS+ys10HYTEhbyRzAY7TR2FrlMK3ivDq20TME5ZjB42edf9MW4f+CF3
WPuCBhEUVUEJj+/6C/fESCBOOcj4oVvAjniLD2Zp2Lvn9YmJWnI5ewT+iu3xJEy2
Z9s9VqdZx5AeQMQGkXKUycVN3rCt2+eOTYm70ngsfHiabb+AmiJvasfBcDrMqkw7
OMNxAyvlJlXSNfSLWIvHvSzOqXxgoOjrpDjBzPjo2fk5wR7wf7Jva/a5yfAePVn5
D8eit0sh5UE8a8gZdIUNOVcoG1UeEGLAen4Jdf3FRD7xiCtNMwfxCWXcKhE+BEO4
8hvfrLpnGqcEUzuAZvSSoY7z1otjFtZD3mKzko9ijU1OEzxdoIz/eRemaBvyBIXe
tQD16hRD4GvP80Ky42VpUvd9Fw69rI0m/v8Yg2ayt4Q05eraZ6Aod0I0qbtqFMjC
q3we6gm+4l0Sql19xv5+uWTIWorb6b3nAYGpHxWoYQbzahfMfTVGb1R1aQj+Dt8j
ESFJT6bSdjFCKVWIGcs3AOX+PSddj++e/YS7GR3lF+rbKHzODtseVB7OM9++WU1F
KBt9qbaibZvJHwTOmuODBhmkmCEPQO2JCXOKAg/Z7tmaFxIGGBNejVwQxG2Di+kp
rm45KBrLSD/wpKq0rOK5TnciDHJXIWZu60enHTd2msiZm0pUcjw4v3eB7Ewy4+5x
/R24i/ukp893cwS7g2IkgjfBN+GZkVtbqF6yIXhBZ+6cIWLXcx++qqp1aDs2HpIa
jfgZOlcmKv1grYKtjoSdEkCIABz75Zoi7nsEH7Lxf28eNeAlRAOh5qY6QI8Eyyvo
h+MGhv7K8uCf4bK865qRDeTJ79MG/U38U1yGEAbaB1QGUIKJkZHXjwe/ctnS67e/
MBIdOjR4gRR1/jL2NU4mtREnPN78trUELxyucclvigi7Lvgu0Mw7twogWn/coH3c
WWy7FKa/ey9YDYKohq6/nhbaKCT9pm7+rdSGHuYQLL+eKSRDxV492qrOQBbbC56w
09hy/Om1nQUNeSymMvVWkC7qV1lslcShxMgvP2FGDZsLK4jWzet/ZDnw0ps5kBwM
fjsEDr2trCrZxX8qtNkh3cbq9Z72YN3iTSrykoFlhm5xcgrLZb6JSYmKo4Dj88un
xVhaRBeI07Najr3vlDjY6JJyqGXM6QfbmDSVGFp8yezUNZmHFq4IEHCRDi77etUE
GFyDVG3pLmod5cakVOI8ZMEmDm+zoR8xhHsNwRPnrNNKY9cWTN7ZJvoZZaX+J1Os
NLUDrry7lZ3mkiQZvo1uV5AZqFcb8ZZwcAxVJCz+oMkzHAkc/5Wi5oiV0o7gO21R
MO7XVHMvnNoSDwomRTvQuRCYvk8RSSLTwKYieeQkLAszNynbH28WgL1wiTR13xXE
Rdmq83NmhIS8bb0peqO2pTQfPHLKdul7OZvG+9Me/Kf8W2dYUdgiDS/xQL4BfffI
N211nGOQ4RjCyVugmNcF1ZvgJa7flc/NZFzqjt8PKENtYKKh8Hgx6Dq4P1bqc34f
TwGxsurN460Lj6xHa7OLQfaEcO3PbywK2yBdTiRSChjVwFxDthgofKhLcsoxuWQd
ysAmu6PRCfDmI8lTJJ2f8Rr56mwC2mz1IA0GNfmFQVnqHhgeBSRW8NWaLBd+x1Bx
zeMnXp+3D4nbda2EBlt+KznLnu8SK/2jU5Pq6J8j4U1R//FUHT7PL/4Fq5DlX7En
JwXgSpwcfMRpp2cUx1NBkeb+TFD2eE/0b49zFu47Ahi3BMln5s2EEzsw4pV+sYGm
tgpxA9J112uAnXZ2RSeD/DtYh993xZadDxgtyWB5VuUXjKAR9KpGRPnbz2TBU5re
7LJ8Dq7/seE9THe5haG1pQpZQkJjVvRAX2gld4DtcvbzNh97oGPq7Unmv8DG/VKW
b3eVHFjicV+6OJRyrL5CoRPnNwJaV/pbWyuLXXkWwgqvSkMa+u1dxz8WiemY4/Kk
am9TLtSc8FJvqPL9eI591aj1M/zJUqPOJ0WaLLj1P5IAVVkhx7kqf+3vaDdFu9Rd
F4vUTmmLp0pF1x8CH9YrMiPih/iba/ARqXQ03zwfhYId1VGaAmrgH3s9o6MUxD4E
JJbRde7/PHZGOfmCDnHNCOVOYs7e/DVkuOF0/l9ZIeejih+B+n6FtjQZ+oYysqGM
jntPXKhDMAaHPQNRPpsnR6aFB8gwSTWqcyuAoxxDQO1yXn+HgXgXq40ow6/INp0J
wd0aKDiw7ug7ybKLDM5oFjiQiJRr57+ErMi69nAS703QFMj5dv1nXO/xUHJVzl7o
yCANxzlSQ1ewZyPJDYLvxFtSCJGR33cWcrjJ1Xa3uTjPRHqFOfPQdEaSTsLetzEp
FyAfgE4F7V7q3qoZ+S23UafXtmWa8R5uY42KqEw/TiYst+nYoJHnzqjmqm2g1jJv
3w4vnidO+Fx/wNTjDWOKIxlcS93mQyJtrk9FMhNV9WC6FnEve+KNxsLOtZlsQmcz
0+FcgHUEAtQZBbxkaqFSFo73HVzQxW1J580/ZkUMOl0dP/aVJvlt28YXFRgN54Cu
38lgP04OSKuSZQfrEOmobHC/dxh/y9mm1gKjCg7LmsMpDiH0tdG7Y8oked+wMOiw
bkQ+yXlsD08NhDswJ7Z280ckoq/Mzlquu4utK7sdvH4Jwh/7KfXCw5CCsq5AK02m
cfb5YS0Mj1Z9TAJiKzG4tSezT+MelC+HvXyxI7PA445H+mRfJKhHaN5gVsq/PfoO
JJ098AR2JRZwe6+eSTNlL6c0b/60pCvlfkUQU8RSoO6c4WUH+mKfya4QesDlrs92
BlQKnQF8h7Ar6J20WIgHD8c0vB2xqjweWVb2QafeZ42nscWhaPqzLB1tGiBA/H2U
PDLgLnCgnLuotwZO6pvDTWwnuEJrWjegplfhKNpSjOLj2eanfXsmHnV79JI1Jtdf
ne8I+XQMgwhkZfwPb5PtkEV09ZacULP+zivgmvbBLeUEtC1QBgWFeTkgYoD1N3Qj
LofkAtzqVmPa9tCb3RgxphlU+O8MD6hkfx5bexq7ZDDAmMo4rxdmIJplyEy0ZD12
R9ec6bB4IlPQ2f2wgOUpWIJCwjmrCVP2PsW+lfO68oI5IMEx2S+WK6ynXQf5jPgK
tTvi7J0KsCfCCxb9EDX0+1MGOwSYesBRXrHaJrPEy23JGKvt5D21azdN9Z84xuw9
h+EBAUPv45rdjLFGhPAE3swrRVeKNOywLPB7O3hau3/K8enfwkvL5GYVaJdifLWK
Zuoqhe54Kosb9jSF1OMy5LQt4GfNRV9o9+HCofmu/SyzEYxrUGaEWVDC/GTSxAf0
z2c71c+2+4vOBEWW7mqZpErcRzgXg7nT+8lG73TGYWXZVkbcDbXN9D7UKLp8Cuqt
qBDsMGITSx7maDj9G1ck0Rlranv8jkdneRsDP0AOO4OCl0/mXIN09qkDSVtybu00
1/lmIWWgRc8GF/txwRLqcuL7jXZgtSJU63RxqJyopgI+KEW6MJBtXbJB4IO3lL62
V6t7TbpNjqAr50om0wKoE5d8UYaqKLfAEuQsaLJT2lxpUQaAPUHxWxhwSWJ+rHXP
WKRKPz70B1Nt5eBUVuUbxsIyKx8GhNrNd8VQQnVFGqkIMkj73hPZHNyfcYZkeYg3
leOzn9gCd6ExLSwe35BJOgcJG+V9CZOXz5sT+wDelHSYGQ3xxPJKcgDtBzhRoTtl
Q8lHmPR/EOmpW+ac8rX86oIJYJfe8T05caBPTUG1RSu5KkkobleUwX7wnXsOZyTm
stAtV4TnJ2wsjk35VOSCKrBoGv73PZpvkWHETHzoJ3MMrSqVoqNnW/0c5cUc1Oef
55h5WPkPNXGcwpvGTE9SLbEZwAMFG0z7/oSmwr+xLhl0qjKcTRuSUEh8v2132j9D
FPshf98v3B+YFoEoGnVLgT+haCh0pRHYiHQlyCwMLp7CmteS4j0YZnq8k7XSILds
sQU7L3nq738SfOJPlZkmSbUvPzmzJ1BvZ8TBUQ3xvQ7/aAizDtZqUY3QG79bx9X9
Hma5UlV4h7hehXtqJs3ISqzfaD+Oxrb4LjIkqFvXldLGtup7EracN0khNhtR1HeW
vWjzpgFbwpFZELdJEf17DZ0o+pWFOHEqyFgRS1jwvBwx6ihmIaEavuVPwJ4J+1ug
3skLcaefUfROilTB2C/myCEClS5wD+jGtSfNDycdAdSu+TUtsWfb/mHaPl0WwxZY
7QSDVns0qjVzGWBWYLCPaGCan0GauOQnf5c9ITMCTro45Uaec+n4BP66286hVxR5
0BohLyEECBiLZ1l4lnRyQ0/0ixty0K7qcGdGCM0amks+74QNDWtdFjfIbux5QIKI
ZWuLtBQyasAY0jIW4Ir3dPPBFkweihtbgSwMJ1bGvEZWcm9ECcSnZ0uC/3EbhvhL
+pAQuyHqGKgGSEiI8BfO3184/qAxL57YMgeyU2s3dFi6LFgAZnm4Q5H1c/B8mDh/
t52n7hGRQcUAWHT+ue4b3Ub5jjYVjoVgacEBH8DZQvTtkxTg/ZFiOXptOUhQjC4A
TmAWCIy+rT09+yfKGU8810T62rtBLaxLd9Joy/lssAzM+PW6g2lgrKaCn8h0Sy1x
6g9qyT8u9jGmyGXEldarCyV2t5qH38KZh1+5mG3apP+TnIcZGfRy/rd97Jn3Urps
b41H06aydpKR2eGHWyZESdzzEmpx+ox28qSix7fNzo4voHGYewUoKux5hycO94uj
PcEecyTdgWyuaqqZ3lOpATPQfi+R/Gd5zVTG86dZnB/ajULS235akzRPKlMZbCvX
vsz2c7jgsgLl/xKAy8k3zXvafNvKyJ0fj4ic/392mjX+woBEiBCwwTkTcLAWP4UO
+rXN4sH1m+i6yDxE2K1Sa0WqVmwE9CIIOAfQGMANjfRzMLn44P0DHmzpGDakUoF/
HiQ5jRF1SDFJO2ievbe++t3C23gY366OWrNg4Kf+Na+WQnkQN9pH2sWuwtOPGB51
jCPTgJj2orWUMWHp2Qq4AiAZo11john7nBTnrGe5KwKkqL6ZPVL0J6kbW0L8Lb1y
9ONkfxHsPkQ/f6GyAD01sTJbfA5eGst+2ErfZ7hFCyvxKOhvUK21KYp7lhfkNThG
M3BX2u5cG8iV9rgmpxBXc+E0kG01BelKbdryqhduKsNjNvV9CIYvjA9+7oOzXjfu
j5wPeH1zZCpb1TKa2O46zlegYMuO+IyYt7X/qQ89eKtA+UrcVbG1dqT2jsLMtziU
95lD9awlKt4lYT0CpK1FRYzIDJj1B8Vio+nDxZRiV1JmDA/KipWHeZ+S2XxwzaR6
yOb0+PvW3I0hs4BqfTxvP4Bf1n3kqP7hhc+sgUonqyBX4/yiKc1PnLT/a59vRysm
VGmNHJ4YkFgFFWXDqON3oGUh3ExM0QbIv7GFeKlnhYIDgR73YpfbhK9lNF4swNzY
eaZEXAmWsUzGWqsvN7NLYa88+QvDPig13Am6f+1iWX8aqIb+tdAQmHJk9eradr//
PMa1iRY0kMKjHeZqNh8+GcECxs7pw/ZIVbZmb4NUVbPXlYb5eL5/BjgCwByN//zp
HmcrFY0ZGWZZBzx14FxWfHKBI2Nn94q/+a8BsprRRc8+1RHC7A7lJ3dmX+m6u3xI
TmPTElfRgbgw3oZ7ls2SX1QQxsm1TEQvO6rEcCaat0yGz2wOy2+hZ6IKmtS8K50d
W39S7XWRO5RUyd7G2FmbZl4I69fMUKU7aa7O15o68wBRlZtIYP6mF0l2ONy0WMOF
6jjdLRDppxiFZEqxyvRDUDCOzAfCl4sqzTjJ6n1jIHpgm0vG6rjdmrDWy2+6duyh
UwntjWr1EKeRcIg5xfAIvRODnOLjyMVqk533dJV3CEtMULgKV4LluL0uaMVkv7Ce
bGX8Vq6V5ucgIEjVmioBJXjeS3e29cbu4RbYtkWcSmsq7WH3qOZV+KrZnZq98SVJ
L7nUvSBU5y2jlF1a3upsK6Zdi0ruk05aZSvZ27Hy7qFkSIejB80n4TdTaJm557pI
EU2FrMwalipc4x2ucRohp3/jk9hXM2h0s0RYX0RkvLKu32MRwuEfVDr5R/fmQz5C
HVlaT2Z9R55OSW0EstoV9dlbceU8786NQteVgeKmBOD3w9TU6N1GKy+xZcFKTfpo
MGyLMEBUC8gO6cLR4jNmfCluuDOLQKLKyN6Co7Ydj4bFezH5V7BDjBJI+dyY9NKd
XUm8TGwZ0IMOVQYt1KkCQMLK+ykR2eFnGKghTgr8DzjO5mHPPTfyzSZ8/eCd9Vfm
Fz2FQjPW7DTKpg2qU+hfX87Z/ztAk2/1+PaszN/3GBsxbge/WnYvciPzcOqqT2Lz
UG8lgtAgpYyyPQkPqRkoC42WJSuL1JjY51pRfefHoo65E5yykyA0pCmnqkUcVrUW
94gKKnmPu2WZtcgl7sOhdER+9C5cFwMZ/LERNC9BSVWflr+OJzqf9yIZULrabpir
iLOVF7UqFSR8L+HOeGqVfcotlPRMXvjUQZYXNlMoQ3m5kZ0C9yReV3/g/LjoUe2p
pOLdMkESIxlyXwLsX8wCz3VcASQtBY7IjNJfykPm7k2Tlcf+cohdxbhoPKjOuFxS
1eNYl62BX8qiLpVkeYjVlceuzyCIjZifzdlV7UMZ/1hjOu+nigeL8pKLor1jPXGC
sNfnUCZF7B1ckwK4zk6DKXOWp7smRSQBe3FCZ9FXHT0wM1h1nSXX4uIjLZhNinwm
MsVe0X9GxtJK7j1lAAd5rONiXV+2YDxDK+4R3fGK/hpd6LlGI9L1Zn9qOkaNxtLc
RZfnTOl8NAi3Dxt5n5DM6ELfyYk6qXoth+JhjaeeKkgoS9fCImP1ONy+zQCgZ3Nj
s0X7dm9sEya+KVgp/NUx5eU259eZmw6U7mJTKZP8Ev559kitsHgVM7nrkWmp2PmA
heBN7B1zSDoKC4GRs5is8WbP+eZfya4Bw9hzni78pQHgbSgp7srsJI9lwvTPZJXX
Mf1o0XCn5qpU7Qb+u89r/WumPKla33UFkReunulhoKBxLyaarpgEoNtyT4t8KJ/0
JMDxQQ01Vzg2K44I4uZQdZ+TOmGeycD3lsyj3NYc0pgWUlmjFEBNQnV6BtX0YdPX
VAN1cFDljSBqfxAJhY4d9FumTg/QOvHjNcyejuuA0beJNW+JE5LcxqPG4UqR0R0u
BNjgSc2bq2SFfgsTjZgISKAl0kL+JXyhtjDHRnhaS9ukMfS2lXtpicLaADZzw/ab
SD0gasCiNPq7+fv20B3o4IW81VIDyj6qNr8QYU4iSv8wu9lMtQud/uNKGNUTu/Sy
gC4JkutIGTC2CxgMkIVzRY17ayQvr9+xotfvux4M3c1Fg3Vbh/Ei+IXvoGfeUVSQ
CX/hT91cTQg3ST08WrxdLCEUdDO9dYV1CLKnhSZsm2z4HQKYYwz4m6ZByqJ+Punb
WhO+7ha7b1jH1Ssg+CSSf+Wp4YYqItIKWA2s1iLCtapeNOcQLT3u3yy5GfQL57w0
3Mr8CMCYOT96tj05LA9k7qytsHOB9/cKXMaiNHp+mxhyKCYaR85KAJUpB7sDvz07
4oJz+zq7BQEft50ychNyEdmMOSvGLY9IH0KsTp7EHzjE4VBWPdcG7cftQiHVFZrW
gQ+ucEwX1fMVAX4RI622EkOEBzKvetmdeAabCKfY6VwuudlRnXVXAfpr9xTP2lI6
2d48ctYJySsTX/mtRnEN98kaT4MLQczLCUbNUfbVfJ/699SN/yONJydlbbkUi4UA
A2J8Pge3mhqn6aoMuet6AT8GGd2gXvydRt0EzfQFHUhQFJXz8aIKoTrFEsq9ATUT
6qRO+1ikEAq0Y67HTIVXp/iLYfdZQAdyT3l7qDTfrTrdbY5wOY6W+Afm4a0WsuLL
zKU38xmNNqwsA0X7wsQW/DaOHOFgTYO5qF7Bw6d4GNOxC4ysvSO4CRtUhPlRDVJc
M/Zk3rWnN0zF3e0q1Xl2gtSqF/sGiTwPLcPfZsOugzJrF2hfieyxJcShDVsfLTvj
VYpNwH2J6Okz+NmtEtPWLSowiPUqCA/KxWZGW/BoEwBlDsyoPt8q/ZLn6Nb7Q2xY
vu2ruWDaYgTuSxswG+dUZBJ+UsMzLXVkNHONhBo+8DAbrbId86QdIl6Wu4Wz122A
s9VYdL5XFfEFq9rJErmoNK8JXWxgTse9SbsftdIHDxoMb/PgBX4CSS2n7SB0/Y2C
dtNyDdmaeULrGTzUmks6N7HIYWhYYpINcaJg5pt1T+nNAueEJ2oEAZy2Nn/LBcyg
+ay2OFnB1LtL9qhVED139Mndu1XjuXalwMIMMQI/30BAHaygwFkjSTA1NTPC691J
ExndhF00ZG2iLQukLSbMgWbe2ZFj9xo4X0sU07DbIf/t0YuAi9zcShEhM+j5dBrQ
RvAQEsGi0sN8pyVFl41fmdQtwuMnlpDGjeEpZKtKv26fTU+NKpjANxETDTHjc7Nq
ThxWIImvb0PLD0+olvXGh0YT8cqVQNQ7+QB/PPEYymsbUTWatbjwYaUS/WJdi893
KizJ50yyMiq0oZeLUXtv0NYWdzBFs5rdF1z6cOyTSMkQZcbYCNYNcNkh4Vg1kTLU
DqBv/9iDYDYtgamDpEeFitN69vkjBhQTU9CzkZTKA9ITJC7ZBYVUXzv0p60OLb6j
WPQ3f96M8uWkvRFqeRsK+hSZ5OJCy+i/NtVetP/8dZBqRaMcfnJ+r+7YSR98WLFd
ttZ6GUYvAymWekHprpZR2eBDJDSdtBjeoIkD3n3JtHBn+ATVl3OEJLwxVp4pkWrb
uQSNeCt9syMEZn8GFcEGEjFnqf0Jh8GkUTZVbHaTl4v8lKzKo9vmFgJ2nlavPdVQ
nqwYHDX2LjCccNdnwOtaPp01yZpiyMon29rs1n1ZRZIjioXQDC34EqhakPNVuPg+
NnClOeA2VxMOIcdx+VYjN2vgFDeumecf1CLZyDi+oU6AZi8z11CzFCnaq19X8mUC
VeZ4xBCJmJr+V7Yq1A4AAYg7KSq3+DkAizhL65cboXKlJ9jG/fIhyi1FoDeVWksx
3HLDEUlyrr+YHC9nlhnXBW5TmdXbLuJEbmSLMuezTORjR2RVH5b0r3nSclkRqv+W
i2cBKMS5E4HdNg0ZPjPq2zO8MPCukuXz9NR4CX8pAYeL0b/tOLtniIm2HYamZp40
UNvLzdkIHoKXo/jd0ofSnNELWIPvccXzQknguzjQD9yFGG6e4Mlkgoz3WrVbLwzs
a/NB8uKneQHE9LhP3RNFjqifgonEATHdPpPBZX4qhLEeqysctdzR8nUskpgzy8q4
9My+/GaFOQOl4Gv4JmWHC+JQXS7gsLb11rntOfhoOpCAR4t/wgB8r/O2j8SfiZbt
Z+SAns9D79OEeHOoyuImRQ77fY0fsJ9kCOP2HG/TEaPqS9YhDRHbvegXE8BUC8BW
uTEOHM2aAzUJ7a2HKnHsWEyQukdSUPc5wJz736etrS7Omo2L4Ha0rYtN+JNpFbAe
Fo0QYMK07/H6CZPKaoY4ymFCHSlZ0BJ6W2lDVxl5mdZzvH3UfzbADAZuOf7B4S0c
jCyE/CJIJoUWOUuixz2NGKtHm/WP/p+P0O7BgHS4TWOKfprq64a0fSSC4SGwhWCf
j7oMW0Q+6fPnMXb+sC/EHchYVVJXCUWiYTUMVyEF+cKqt09PRBTfvot7pTx8shgS
PKCQf6ssQwhnnGuKRX19n/AgPbi91aKefP1k/mBCp3xLrWFOJHfsnobx9wt+gNTO
9cw451ELy9huGqrvcHeShp/PMxqsT+DH35o2AuGGqkUjiVyuvzxkmT5HWt+mu8pA
D3SrekMWbzLSvlGny+3hg2N2zWqHG2NL7UKqjYu9riZHuvDWPUdKEa8RETi41Pau
Alvqk+zkUxr9n8E4clJbCIHkhwBS51HrzAsASKzD7XNnSU1/db1IgqJ3aH9sYCjD
nBrN7NP2eWUOAE38fga9tpLQZoYNeeK7Qt7pDFldL9T2bPgszGNYO/BPW5yUW5ng
8TL0Gmf9bSt6IyRbISM8tqF0hcRg5R5eitv4iDm2F+weKM+oGbxBhoNC/z1Ywkl8
8B9W2UwXH3SOXCsp4LKT3C0ZgS4UhbIiGOdn/e2OZw56BlIHPLv09FJ1D2Ntau50
4n1MWgbTsuy7EV6Y8fohbF/pVTlkF8dd/W9Pl3XPsangp1Y8MPoCofNL+wfq+cVC
IAMp5ZtYQ/nsG8QQCDT+IqP+fEYl8zrCRJgzQ4mMBnANy96f41NJSnudl1ZdyZVL
0tki2uxX/CO+Ow8YyWHyTzjYOC+D24ONVb0pKDOq8utFBuwrLXZq2gAYezcGL+pK
HelRnY4uNZT69yBpACcaMzgphfce0Ovg0BmIxiQo74hnF5uWzp/xgZpYz7PlT8LW
6Vpn8sFtcSBvBlru+Nnu7DLO2PfBkrZ/sMsfanpKHNgNvQik/jn2yJ3NzrsDD1DU
GxzwRELzpQkQmvFC3gEZqdMs5QjT2Jdcnhkz9DRDokIdJXhmbxs1cKQCxaJ6FDKW
2IlcQx7GxZU6gP8G6r2JV6GxUxoyGt8A9TbZl1Kn0nTBgO32GgCBCRAxJoU4qHkt
sKmQXmSjFc9MCIoXTP2a8mxf0kRrJYlUqOH3LzKFa1vIOd84BAFN2bgWcy6539NK
MB6Y962fBvU/lnez833IdBk28nx3QTkdKxqxHfoFILo454WATE3od6wwYNwxMlRI
PoKrMWqDP01VaQA25UcUo0MmRO0u/ROWpCo5XcM0J+tfdrgOO3gEWJB7qDQMGAz5
qlj3CghTmAoGYYf+NARO0sAmI4P1DIS+/+tCCMcbJvuUs14193WZ53uKVYIb5sCE
hhyvb7CBe0VW7udLOhFElEIMjeyqZxz9N3uHDwfj2Mq0jFfrHdSgbgm0yJm1vAKo
eGBlNj2HgJjNVKgzXxfJ56BevIntrvBnAtWKHcQFF8GTYN0Pt5Fijr/lcCzb4ttE
q2SUoR45VYlwiDHarBDv3WwOzHaDa6rqt5xj4LW45Tr64v/wX/9chzjGus1mw/2/
jJRvK2/gw6F3VP0yHHFwNPTBvhZvuRxUhOpNXb2O9wAaNJlbdlBQVZnaRPBzPOws
ioBO/chnSRx8TZOYAS7U5ELL5Y429pq2NQm9LWGFaetnNRpzFFxN3SKItutMJ8/c
HMWGPcDzml3taWvpve9Y576wFCWOgheV3bvDCDz3ZaY3aAJYilKnyCoHl6ls9cAF
5/L9U68fAQUQc9DSJT3FO0vzl0AQn/GDcsDw/OFrIPPJr5XTxxichUnHicZJc2bw
dTKkcI9D7KkByZa2PxbEHgxSDgG2GGIWdj5i2WziAjbistUveQquce6OOIgz2oD+
oyFINVbaQ1FCQOznYW4kwK3oBF6WsoJC1ZhaYPDrwwCKS9m/AO8YqtErU8bwYNGb
GqQ7+C0DGC06syXVCAHKFegI3g9+Y0Tu79UEtik2A9wcAxsIGqVA4ZbeI+bRoPFd
goyG7t1yl6TUfn/Lih5Tc/TFrmbvU3zRCdWG8RmBvuIpOnHjrcVU5H55KT+SZ0JT
RuL7Kfpkb51oOF989PwqfY1GcEd72eh2aQZpHHm0Rm261JiJdKBqE/GawdANQaSe
Vgq/36VSx3J3N4PmMyfD7e9p1f39BI0Jkn2TF0fFp6Q4ju7QLJmOwX4kfs2f+1Na
/uP0uXgDfg35cp9zVAUjqahNxTfIvqNSK36mUHGBbIEumqnTQGLXS1uLOWVxm5Av
50LOHPcp3Md7iEydA2xzAwBcfCDUYCkWD+04+lANymBYVJ4DtqlTyRX/iVzVFwY4
bgfAj65g8y6bGFNIsAwe4DPS444BO/e0TxLczV/W3/G4STe6zPT7/M/Y2J4Umibn
nnp8iCOYV57huCb7JGJR93F5al7RGRjwWWU6TioDNhsa9rQkiCOAHDxPclYQoVFe
J5Q5dMVHV4BLoqebLJmxZdGY1W3vWKmwiU6ZCv3Sot1VbeCDyeK3ufpF4m7YrlsK
VLc/bYcJT5kKfX85Ps/Bf300bPhtb6+jDN6l8kll0CoCJLE5cTbxefMNLlTAKljR
eVmoqO3r6V7d5j93T6LwZgd8GXPz2VjkYP4mKr43rkPdf2YN4vgzEilUlvdqoqW9
OFa0ZPCqPckxMElRNPL7j734YzwZwg7kIUClcoct0nijcDiobp9YS9uxLTDGcsgY
x3XhWF06KIXl5IdnVvJQSaHeN9/Iwmlyp8pOvcM5Vurat2+Q83za1mhrBuyIl7P9
dDOWNYgChC4p5iNJme9UlP9t7kNvLPfoHsmbKLVhqwCuXZvEloCJ2oEWvnccRGEG
iVqdV8XjJE1PHKB3K4o/l8dYgvRx2LASdxs0CqyEra9dgfTNdlJsx//rpCQBiAn/
DmBc9QzHZnXMhyl9TwuBAnFpHfCrHIqexo4fNfvbboCuolyKbMX34cy0p8L9S1gU
xBLf/Spb3peEUA7xXeR3/jFNhsQnVRZp4qjv+LfgzCWsUnoeTyYm6d9LypCfxcVf
R/YP4Ex8l9AuChJBALeXpV2dAVAqukiAmqzG2OlhofoxU8W5YpdaaVzuLCjomtP4
fTyEvSm3lguAyyYHK6GPvP2et7jzwP4WqfriqeyAhq3As5tZNtQNX3J5ZUV2Uami
EqCup0khpb3ifkJz2QIsbncONaVb+cZgbQv1UtLfnt2Uc/RGWUTMSeW3Z4KtBx24
uBDkQOAQZSVpwfvX/dlbdLKCxcR5l8FUjzl5Ww0G0IF6twcQax6baSP7L80KFs4x
1jqZMwSmhAvEt2VtWbOEQYiEwuwCNESdxwM9QVY21b/QuCT5pWnfgycaYBvTnBpI
+hi69gZ+Rjo8pBJlRXw8kIeXGICrzjqr1W/w/3IaWKJOsyL8iYU+e1wbrWZTO4PH
1HzhR/7xvaXAzvss3pEROYUSzorWya4pMrl0jh+maVUrDVOJEOfftatFrmd+sql8
B0V6NDP3Q4tOJenevCER7Ah7oSWq8nZubrf4WLQK8GP7T7NkAkL7FJ9GIkuH40Ij
HOV9eZTsoF1JYD1WDnqeooayFPk+J8eRX3m3nqP9sTSvUB9h7pms6+bZ/rEhZpG3
XGLpQuZFOKiYBJ5DEutPDf4wJAoJpE7y81l18Dwr5+qS6V3EDlX7nX31Y8RFKKNH
vWBOUT5E4oLv//OZyDxbClWYEySO21+Rl+mTDO+q98bkZ5b8cQgZSy+rNQ07Fqj3
6OxomWGgJZ/G+hHULobyHkXzR91hCcKtaSaK4se1TjBYsg1mk19pSuLvVWMT3PwB
ic+cek6HHHBQdrMYWA3qUjimp+w523OOPpUw1oM2/V/QWTU6JPVEEmWEty4B4PrQ
T8J4/WaN1RJUsLkz/3g2+w4blGf7MNUG9L+KhoanBqLOh4n9kFkidKs0fNaSPDma
2ot0miXxfpG0nUjBxEFx7NtluAtgkSQDeOHuIlQab5UeRpaCNQAoJagXW2H5PkXz
En5keP2sUOGeei2unylDp1pupKF8S2795lLBxPpCwhaHJElF+GHsZ54flXQNhYTc
2/Z8uFrJg5WuI+GoPAbp/Pi2R2I0Yz/lNfVkRtvhSLddO5V2CEXRkT9tlPNjqjsH
N8Yg+H7o1Lkw1bFcH/U+M1r8mrYpVkkRNWV+5SRohmc9Tt6NGjdqPCrTKx2dQIzw
IUDGtxIVWZtMd6mhx8Q6gXY+cVaWl12g0tIMe3T+P6EpunDqhh1uX+B8TJ/pNTdO
qEJskkiQvPxYHdXuSTRq/LoEl3O7XATImiwziQnBBmdVcSUSqpiujHV9wl+wE14K
R2ZVbwDmHDD2bXDxpVWCzeU9/nDRcE22Qlc8j/S9CW0UlY4nB7q2kRmGoko1h1+T
QkuvsIab23aCozw5FULf5lPW902lXag29C77YgJDOE4Gj/nSsuzVcVQAQiRPLSiP
wJ9hFwlZjlo8hKiHO3Zs+MQ1pLlYP41pkNc2KUUd3NNr5F5k5yg2Dzq03a3ofJnW
n7tSYvit9DpAy21hoIz8S3IWbdpP38Siw554PEfwnsxPUlVzkCZEU88FqQbLbqiC
AZDmDfO4cPXeHAEsGO04VEgIkM25eQ/pJ1go7uFmTeXjgQxI/zV44FXrIl1+SN08
bLAmA+N/2K5xy0sNh28J1uy+afhy5vxS+tdK6XJYVqafeHWoSfjNjLoVrzYqFLBc
ar3CXQrWEGpjCVxkV3QO/2FDST3iUZqeF527H94kpRg1W441iyHD4vLalvVGCxxZ
4aF7NsryAXYFkpFdF6N4ZvCUU0GSIttrQkxviPSr7zOMDFjKu3U4fLlkBtugeIrp
POA+9hhgxEctmV+kvh/mlC14YZ7aNU8xO2L6vEtw0gY42R8SJ0kausaGhnJZRABu
Cw29uHm0040tmNTmAvZOchSjSJ0IZcKQskuBGGDjJq5OdDWJiXWxccG+kgrhgyzT
PqejrZ3OoJmWH/9nC8mMf8MnI8IfUTrEWBmCLT6pgKOdA4bmTTB1wsTqoMYbn94S
ftswOtWzjtK1Mk1PWChXxFhEr0VgB7yQlAtehF6TgAEXBBpi0Zktqm3IER3XrmOo
N7DZkhwCABaR10TgOe34qVdw17gk/C1THpXesks0QF8pUUWaRR9abwohqA+wyyaS
1Bn7gqzUrLmMJOWWbO/OL96+jFNAydOmuYzuinU+GJNvVn0Izu1IyrigHeEig8HT
1u9GKPMLijgGJ8lCzHjAyUAh7DCUDHoMdSvunciZiMWuUKwxGN6T1sKYE9KGp4QU
4L+tcwXE5bnmyCXffgruglmZBFdSGwAggoRfJ2oNYKaO+lPsHeynNEnSs4hr7USz
3k89hRxNLt7Hjs1PA9SeufWDsNMeYSpTf+0yihTsovjsh6ZfyQL7geSDsJVnHFYD
UYhMUB7P53kXhiyrKENJLtylPPOXJY5dZ9QewjLXANA8PGO/a674OYjHKcRlPNyC
exgrJuWmkINUryeD7FjHb1aLc0qRErWy0QB1Ey+Dzzz0JkHjCZlSr+SxbKq3vy94
dRqT+RO7brWKz0xrtubN8LUCBNCukzgtGtYCpYyi5c5ejaN00Ku4dYWyjBj2StdA
2RmWcvyNoXTpIMTz1o608yhoY3s0OKsIQDRFgUWe540CM0sMTaT9sRPA+xFNJJuR
6sEXex1dX7uKizznibtftDwhzW97Kms/UkW/Z28aO9a51zEBIvJY4lGJXa2zzGvW
A0Ch9seOLcCfQuMRzCRmAskebly+/maPeC0i4HrkfZqv8bbJ23Ts4DwANB6z37Bt
q2zjehTASYDGetu/2pw/LoP/I+MGMTbPV6O1qeqFjkOdPIOqWF5Ft9zoL0TF+1YO
EHQZ3qWHLNlgbL5NCyMN24wzUzePrxxU7i6L8JYC4+xHNTFifQLFbr6wj+QABO5A
dDhKAHW5jGKfEuIPmhbIDzfWI1DMKYbSu3S6K+nQg4pp+KswtrGlJQDsDdWQ4sBR
kUB0tdhUqNqn28+ilGUPZyDqpaz5uS8udxu9gThDHJjIM0QM/dI8v/6yOfvWn4gL
U6ekcdjvt4OB6Tr4v0/R9ut+rmjgPP/LiqEVmWWg3DrsLyGLXn38iXDUe8j7+J8z
Vb3Un5lgtyN9+RUorThNMGk0EeHEhn+6FU+JGrs5znMZWMSMr45Hx4bnS+2ovlo6
jip//kw6VUq65JWJkD9POQJXqZEeVcKfwizzCor87SbrsfUSec6fYJKkaUZSwbi9
H1wlNRjr7l39BdC3dVrat4/lxKxBC2CytzBeqTmHw8NJrBpLvqeudr9c9KSHa8tU
F5/6J+ZapKmib6tWMmmXnR5ZzNYckEUQ/2HiJ2J5V0jVDMAX9wwenLf8U7Nfiirx
wuvUZefTfQyVgwJ5dHFO7CpuYzsFDOACei+Drk1ngusZMtu1v9ciZVR8D7Bs21e4
d14Qb1PrnUeCJaUGnuVrmTX4W1agF39afNE4/Hmrxd3eeeT9X4GWM6h/SivIXYPK
xZSDCXneRkbd3xacS+59BjOJKX7djTF4yubrMhAXMjZvS13R/9LxhVGnwbeWp6M0
0FNzIM0CeKcZdwDPSoa238LUq7RmRl/VocQ8PoiM/dI36J72NAMgsrkjb1nvaiDb
xrAmHvPEZTRjD+3GGTTu1K5vYNr7/xSSM5rfBBzvMv52H/d27LAsX5SpgTB6K2Xu
UmEuaH1mPT5uITS7a5s+0dIioqW59OssqdwcdWGo4RVLCweNcFrVDA68dokpNL2y
YAldmppwTDJYXmxtpPbxdptAs6eGDs0GHJZZNonqgMN2kOFwKKhFV+iUJTay05nA
E1pnbvtPrAVIlaz5UTsxo1eX+z7JGlvtGOoiXMdy4SL2LDhXTptl3MiBbqaXGKtN
XDpyZRyJ2sNo+mo4PQDOzvm18rrS/X3QbvNFSSFk6NIXQ64DRSCFO+ycjANjHS2E
PP1RAwW6SSPUldc1borAs0FE1QTGmki5h4bE9Ex5Ev96sqUK3ki9PjNjKVlE7Olw
Xo2XB+Er6hItzG0WaFqwsXcgvYqjFSM2otCmY6QmzGH3+drljkhr8XOFjiq1imY9
HTgrCu3CerDdBp3gySvAWZbA8QIbDJ/Jq9fPXIx2CDXQ+jpfCXe9MpV9QQ4NV6+l
4YdJsZ6MCzI901g6zE2RtbL8W29H2bveDZiYZ+L6j3dfVN+9Vnakt6mO7ys2dYo2
DZu0xojfZhfAPmDS0RgX7lUnrxlkiDqXYssAOlFb9ZV4nk6BvxhThxsv6f4HVluF
kE4vV1XU83il9v5Yqr50Ss4zMfMMhN/JZuZUDOsc9fLYI6jLfep+hvlmhpDiOGAc
gUhiMbUkAq1E7aupoTmviQdVbH4tTKbHaVpeoCDZ+FY32aAQVgxmHEnWwhHtdgmd
TOUaPgVKEDjST59ipeRFKObuKfNGUC28i4KGwjxM/9A69QepLtvtIsejv3kJ4LWY
aw/WJ7aDpI2U/RSSWK9DbQffS8P//tjzfei+Wiv82uHaJ/5hcL8lH0QuFw7Pkx9B
x3AHfE9DoDtk+I3uRpOhMe58k9o6zMVAy+O0C2fMU0crBfqE5mcWN8kouc2DdMuG
KEr3PUhOaSE6zY2anbE3abGBzFHK4iBbQWJ/w/id6vR3quFoRAMyu2ZicNDTaU/b
QF+vkoM8S/DbYWXQn7g8nd10W7KDBAM0Z9n1T+hq2Vv+ggaHV1gmtIypgC+gpqnI
Q/1IkQ3AbdsYgWCV4lESO908/HAQ7NcS+wXftfLPhoq9sBxU6r/rxtaO0DMJWJz8
PFYruvHKvr75SlZgj6xFFo6VrgPfWXN1cAJrlHY/mWT/KQMgDmXMu3mDtOaZGWkD
TluCh8rPunuoRpLXsFqolLTXalyMTNec0NxeweYMqov+Xx+8Mdv2p9r/0UdQStZH
iHYNQqhvgUVWA8YV2yRFOvePSV0UAdo+TRK6d7kqRxco8DITNn0wT8ADjS1i014M
9PJUfjoA0DkkDvM/JQeNwdDX8ikOtyeMzpgWE9m9TORPbTZ3GrwmVsKdNCRdgEAz
sBrI3OufS9pUOywAIAJygegN/mBTwRik3DZa1PSfjq4bxa2ReK6mMDDS19vcKUIK
33KxHcEipY/zjCM5+I4Y/ai9QfL5zHzF/Ol4FvhywDy+pXJ3S2yZV/J/rM/QDfcx
FEGUsqbk6AojB17jICS8LunP5kLQIMLEJFWWE7xLGd220a4YRAPNSq5KztybLeGO
00a8oz/COceW3hP39WsbFiYfcgnueqS9eEd8zwbl6YXGXaO3iFSQk5Nc1gQ0qTx8
7B0VnawInhKy/KpcNgOPFZeHmsotusvXx7E6bWVxAy8f5O9cYGSkNkLU/hmK3MNC
L6IdtV2aM3l1EaSq70un5G2q2oPf4a1YWZIIOAi2iDc25S2L9OgFp2dMlLs8/s4k
RLtXcvAD1VIDtSQrCJ4ubh7q0nWM42qq8hkcOdhCAVPt3qlpR3KEqjZqLtL0xxhR
xshKSdHMuJQKNSIEUA1N18BHGRab+7uiKkOUnV4AA/FS1JzPtyjf8V2hmEzIfatK
GAPYd9lCs0Dtp7b/lFwOtaCFJjjkL+sYeOeFgAp8RGopDZfMsH6qLHf6NO5A4/ov
d9dRI0tnJqUHbyXvsVJQgSKRUDcSqX9Ajk9wCmoApZ9CFhtfQTzZoAWqvqk5D9Xb
AUQaUyZ4ByB+g88MfMSvUE5d89tdkXRuKsvDhp4oAKqfKTsMOseAzQQIy7IqPqna
1PdN4L5I3nX+i9Yy5lcvV47zIrw9y1Vw5Zzg0pJ6tm2tDUO39Kfsk22Dqbi4xuJk
1Jk0QcOJOlGetLmCohvTY0lsAAvNNzuTEYVc49jVNBDFF4OShb8CMPDKXuv1sUsk
W+eI0ZSQyZRAJKHwGZCVGhnUc46KE+f3+I3tIfigNooLvAZ3IsU73cb1OhaFdnMs
SZypkISaNoeP0rRF7uOJNGQGYj3uCGJRZu4vyw9wUoujpj+SnFE89rR6LlTW/h9H
1k213vMb/d3++/wF/5ZOAwmOs13h6oABdmOokXnW0Hdl3fP4y5yni8a6OpSWUVGq
FnRTtRHagdsEDrqgd94/HhCFBvsv3Pj/WlMGU6/rtKHWBaPYKo2Jjszy5feouSXa
gSaUBLBDHGki11Fb7rfx4g6G4H5mv8lnz0E5/db/Tub32xjLBEmb5c6AGsGoXR6l
Jo+LS2Q3iW7fWlKi7IV49+38sCv3qOxi2JLrVWLzuvogKKFdCOB5YMB4eiIgL/i2
uwOHTQlvA45DuYhvE/27McbBj4Qd0e4uKymJ8N9IFm/8lofXoffqKRWvyFdsyUQm
2aVeE0mBYtLhm97jDfy9M+NZZM3fKON+JcMmPP51UUXesB7CHCJ6Ou4Hy81dgQt3
xxwi3kcdbSV3g1DBc1pTu7EzIPHssbK6orND2pCTekm8+RaJYFtU5toLwunqo1Wo
GvyddzA6Yk9uV/nkOQ90o6utgy5ctZ6mMXO+L50VWNqmx+n8te4SFTK3NAIgIPnS
gfK5BKaL5P6NAPULThi3bNSB6m4VQrJvQVauDahi9JoFmwbl7IJX5ASLiTihT5Mi
i8qoPzKo6i3A/4xZcRfX6TC48irrvqjawuFoxrvQYp0b3z6A63xvcZcVy6iIERbN
xmQQG6icSI+YjKOiTvjI1IYXsXV0eqmAOR900NBb45UzYTIKPoAjl5h8UttnXyQD
0tnimtezxJLT2hUf2ChKowpVAVHTQwbiV4lwBwTp/MXQNoiVTjOGZI2+GFRXttg7
HjpN6Bo8FxgvWVuj4ZLT7pwF5UfwoB5qHEFLbSMUTsRYuFDoKb1rT2fhHx/ZpV3c
NQGgCKs1m80U9W6RXsDMWIhSUY8uuNXA4chTK2SxK7TUKNjkB6fYHk5TLxnu8Ok1
sQ/icO8+/AIZ8vsaUHJgf51uRoSCaBvq88TWPjN7Sx47rOEhYcm6XDh7RdtsTvEc
lganmKJYrTNThM3MmnsGsPGNmehHZDBH5VxxjFelOwaacPWY7tygPpTHm+H15B0S
DKSHhRHUrTj5vx+Ax4lokDRPx+OvmFqCFcL22WJjHW7o6WzuUOgZkY7ZitU9e7X6
v23yLf+6nxihX+9A2DUYNqKue6pc1SBOc4bBvdXwyg96hiO2F1NK5JYALPvI+kh8
2NyIyuVzZHtYuVFcSZllQvtq0FrFy6h80e2D7RALByYmL8QA+DM8ERHsksANcKj8
qANmemSf59U+T0CZLdPkbIVJFXQJfJoJXSyrZBQYjaRKQGhMzCRCapwkrDpPLT1v
3atgY3Jke7rzyeu/WWOzGKEOipkvf0TEc2xScthpATdf61Zg/6887779Fb2PPKQU
H1EdHyXi56Badw5NyFO4csVDLQ5bLqJvpW15FWtgmhBNGpP3YO8nQMQRrnK0qjKU
H0Cp+StNTeIbXaBRsnsYPYpYsHcxH5sK4OHna740ulCvz56G4lw3QtCtvy8k7pUd
VxnKIalsnqu/IcUAvQK7aYZU1YXbxdzB50U18fObZMOWtki0sC8Pdzk1MAC7QV49
Z/ciL67phPn9b90PKRDPywe8eDlD2u58QBKe8EKQPx4TUzwQXazKA2ssd5q6MoLf
cxMuam/AaOWcPwcIP9eeVFyJVteQ9yD91IRkWiiWyfdZphknJvz79xMJInqNUAox
CNk5ooEip7+Zv6b6a1vezhrvd71k0+3V0zHUNvK7+xJkjq0OO+RLBsAoyaXlAQon
E9WhqsA/knk8oBygSztlgQiUsMQ5H7OtEkukxtwl1QjjYleFyHJntrXpqScGJTTh
1qHENFkf/nmNoZDf4duC34s9xJ8aUeDobygLr7ZpnY3k7Dg7WMzcTw/smF8KxTLW
lb0JmF0DVDIYPX9OmCt/awN1OD0bivF139akchcsm1IdDA1YE7ypvLr9Ox/7ntdJ
g5VVkVjcwuu/V/c/LhkrRC88gTn1mfaOUQzcXIh2NuVXfU+P+gUhl7+SE41tfByh
APOE0rfIZDliMokNcgQdrZlfLaQJjI+G4Gw/Srf7feokoWzVdmGOcilOlSHhHuup
1yLIz8CDwnDW5aZ2MjYAvA9dhuqtLDj6A4dxvLxfCLv5nAwUUckP1SiLJ0nkuL22
P1uwlykI7dTTB4Zid+4sKNRfnKOuXJTJut82ILj8eEYzZidqPo66MrWYFnmtUE+x
fjc4ViwmOREViASvjSIbiglNtlrbtHLMpRrytxWxlSxUwHzKKmdZHnSSRhWkKR9A
pHYa9eIKvKFyRJg5ddsPQR/0oEM68Csq2Ej3dUylTLWdJcIpSu4/kW4LZvFxhw12
q8SoEo5Hhb5ev73bUFCylQScQimJoNpF+pjCHfUNqbFILEcZXCikQkoJM89ajsfM
FzUcjm8tAFLximnzoIm5Eo5h8+mdQ0OntD+xEwC6fV8ysKhrLPQMiNkBhxHGuwuX
DNEVzcc/x0oxCPZYbn28P/VkAzBAazJJO1l1H2wYfG6ktK/zTnvngMszQ3TLZh1I
RiUX4wOXfMMS9p/gIiKYfbOyKBhzXH/ZqiqZa38cf1IzhFfBjy3ZF3UCc3RCE154
MuA7qUd1C5s5QIAtv3OHivm79TLGxLRoRD+MVYfDzqUI9hjYb2Tiz5BH9UwRAK/P
jze4gGM84gKwPMjbF6t8Y2hlezvDsbauGowbwc/f+YNW18nIf7ycc8mYnZ5hvlKb
P8EIXgQ25aD4ijeIcjIIXx6ATrrZa6MfdBi/oi7zEsM1XRM8n5EsoPjmgG6rDBFp
6tW7sM8ujFE4TvmZVZq/mnby8HovsyVWorVFmm+5nOOVGJYBoWSRmN45UcxdT7Rt
RekA2QXPdpDF8ROSl6FqZKwA+rTB2ccyZxVxtkxbJ/1k8Uia4vywM1vtyj+M86nF
+zDmsOZGEbX8E5CpE2mh7otRTDi68ct7TVpdb4MDBoUVMx592OP7dW9oNqjtMtQp
MiJEwqWu3L0SbqBsG8JB2oyBlp01oQRaOuNJnL0eTFvwrnCikr8FdBR5TBDaXm1h
NU7NirCf9mIyWIN6N+gxpvVhZc9uT8tCVrbJ2vI1mfzS8o7Sl2NrGfwSf7kixm/F
ji4Uhd0ML+7QsOXIg+kFDhT+1R3J8o0pkG2dq6GTnGkI1ZA3z05Grw+cNcrrBqiv
knZIu7WsOrW1c39dNnK2R3nkVM2/fSzozBdz/YZw/ygYe+F6oDWQNkOJ5JKMmwGO
KWb8gk48F+Ce4/1WlaYK+a++CoDTrb+dbC4eYoriJ+MrhlHef2qgMQ1w9kpLAd63
YNoWxsuzRB/uK1Bv1FLHj0NFhe1wg9qMArd0l3lsa7vsPWbyUH8YP0hCq2KBtYm7
0PoQfYwG4N8ap73JWSXC4M0DQCjl9Bcn3IYls7Icpbo+d+8830xyEerzAglx+o56
PafloN44BS3qRhfC0Ui2xCNxRrQ2Kx8VIDfQ6FYpmSvimP5pP0W7aE3knq3Dt33L
ihnGn1a+etjGL+BJEufHCco32yrYwnYUUF7SBIxHQ6sOTyNOr+EWrtVwUHukHPbH
q6KY8JDtRBjbhctsGoWd07RDRlwCHFrFpq5KkzZtZVVOo/tn2rsySgVd1z37f8FB
KM/mJMtKm+oSCH4aUFQs6MssOxj5Wp7UzIAASoHo6mKjUbEWQugwhGu59Z/ZgQ5b
N2VOvPqzWBXqNQbbMThzoc8Xlw61YD4P3tXelFvB+SRSdXDDCbboGh3R9RiqXNm0
wooTs3bHTFXB4mXnwdfIZD/xRl7qiUMKQg9CycWSQzz5dqtwkphPQOTlwaqvH2u5
o+WcOFNJtwE3nlBFY3NT6JF1gx5Ne3SBUu70tmI4egNVis4ZNTkeRVhr7mck8XCW
qguVnUhljSncRFL9aax48Ka3cRSoc22ZFdHXWIHJ3F+UL7bobUKm+z4bBwqdBB+W
RjmicPQY5hSxEBw9pb7LooLhJupxdokaefKJ3al0jqeglPTpwASetU2cjlpvOU4L
XCkwDPcRDpt9EHi8LR4DxgMtU5QywrqeTW5a6w9wFQrCy7QMsn8vsYa9Vt0kxrC3
M/3x0NLZbJnAmS1k4EVoxV6nKBNYSWhUpZW9wK4NAri4jwHHm8zoXRJCSG//JYwK
MENxJg6+4v/YKr5Slf+502HCQOdsEdn8kQ9RIt9q60/lgiEnRCjPDs2P8UwrPPCa
h7wHG5yfL88xyxmK22jRW6mrdDo97anO4+Ds5ZCr3yFlf4K9d1wTRSYYmzVWFn+Y
V101BcEOn+XVVo/FXfrvdrg+bZ94nRAJBcnsDiA+E5Sk9hp23UutFklWp9MTIyaG
cWeacQeXJvMFi+MqwXQZt4HTxbwuKMQ1kw9aAEjxLrbtDts1On4laaenl7Ao2ZDB
Ub9SQEYfTrmzw5ljxIQAf31TjXE5dNDvYjUFgpPVB+UfeTUJ/sv3MZXVsUS3JILJ
NMTf7uY5aCNpBcy4b8a09NDnj42H9QmbwnNofioeHpmny583OOGYExnilU/qQAPM
2mcDUPGLU382gor/3wPruCbTAojoSMh4ahTQqiEUq451HEjiCKn6G2E1PhdGK110
BQGdZfX11EWYsaAnCogTMH/ItnxKvfJ2S62AJXw+D5g52IPktHre8AvgwKhwa6eI
IN7Eevhj74nBlQf7bG3rC3Y5V6V0EICpDGiHhaD2Sj+7h77Fryqzrq1FCj92k5Ei
YeZSMQGAEUkBTSsVQuxQYiBgg9NaMxkCySQbjnGvrsKDNFUMMfihKuiPnhsiVv5r
27WHLaB163AB/4uKNA2VN9jdwSjTQoXVX3aUZz0cp1eu+kqsnwnDlNaT4R6JNr3f
9wCS28jDWkFu0KrZ5yLAKyW2EVJOT/ASWoBpxaEy5HAkw9MNkGDfjWPP4UhUkPA5
PCnnO3C0dQ3blhbbfHVBC4cPkZcxfxCWu4WAdAUZKzo6H8u2B7AGY2mHONzVn2gt
3v7ym87w8k0Qkz1153rgMaECBTvu0fTuCy+gLVjITzr31smp3D+7RQXMn+T+dzah
gY24ef8yNanuoXTDjXITLFYNPoC97ZlPO0yTKOdBgP52KPFrMfTSKz6ttHbq2mH2
ImHU0BPwFzhy4QMqm4m3nqa6XtwBLjZqw2s6bCkm1+T+k/XGq08HjFfGIyLat9jo
Mcnd5iRIS7lJQxv0FKPn4cIqux79sLe6SOBCU6mGh8a3MCYkeaxICqu4VwTNxbOR
BNErtf5Pl6RKNfsflWXnzmva6KeJLdV7uvRrmcEAqGvXyicLX5fxMEG05xZGepXY
LRrM6sK6+DoZ/rwqS3ENX9T35C7b2kX931BsjNaeI9dulc1IfMryBRFBe+uoED36
GhL2kc1Z0IVF3wKp9JrmPCwTGJXA0iCgE7thBL4OFkoSlj2pcfmav+ndHHUvBYl+
G+PEc72eJ154bxIq821/nx2pRQ1spZksCbJiX9+La+S9Uv/Bf+/d240Ozb/9g6rk
H9kjvG4bT1xMK37wJD0AoKdJoZg4aMckSR0IgR7CFKpRaazhL9lXA0pwxLjQcaK/
ZMI5y/ZCvPHI4FeLPezlzSzEOC+papNYVqI5rshIeel0Zvdda1pSGepIRkkIdLfl
LANSK1c9iq7/KT5ZNPm80qI6vHXxU5/z8KNgJihKQPzCM67dKCLPdfEZ4q89l8GF
oVeaPEI5yuHTmU8dDDEx6OjVC8M+uoeAuRQtSIBr2hIDkTUc04Vm4jEla6Crxlx5
R04bscqRVSOEEn+6I9KcY89k22VWGms6dxxHKROns9eM7H6aojgHrQTP+2fApC3U
iTb4E4hMS/Mkj4QVfA4XGvs7zeJ7T/E2otaWTYrxN+BPpPT185u1dnNaZx7V/ewX
UdgvIHIgWLKiwmDDceJyDspiyoWHQgERTCOHRBxbL4gdrxNguR9mQMdKSnm/CE5F
rfYT2J8KqJiArbrySr2TuJCxhlNYhBvnmlTva6R9GuJ65x9hhhUJ98ojBL3quFXX
mSMB+QD4HQd88wWQDLBBLgfQyTF9DgEFVcZEYMzUTBgtUjjXBKGtDrGLnnxRS4Bo
ykCVN7zEl9jhuGwCBFNcYzbmMI6y4WpPPfGFwpCnlk8JRuE9r4Y4622s68EnGHZ9
KRjps5NunDsugUHL1OZ/hrlm9qs3W2DC/F/+P1psC6uDJcR2zdFMmdGBESLPeb1E
rU7EieqG3Ipt7KsqzrfnLJ91vvPxdwORfJBBQ3V3gdrR1aaqNNnt7Z/UW+fIRz4L
X5A9tpD28rKW13LD5X7RFGFEOj+SSRnUFUgzoPWuynTe94PJ13NvuK7LkccHhB1D
3lEDx3UJvqjiDkdCtoKNSVCGIUvIuP8OR0aaRV7hE75rcuC3UdShAPmKpQ1YF+vt
dotvj+64nE08N3RsEHC7VgDRDzUc7Zq4OJGxm1i8kvJOh90Qe4rkod1a3MeAntFq
Bk4cc4cUgD3j2sF/GAawFtQc/ELKzIzubfr6vlVl0CreX7d/ri3Qw+/wjoSfHvUG
kwYOOmbzFnONM04dW4ubh7ClIZJ86YJlhtAh6ZvBvdviB7n13mTkY8XiFLlozDoN
8mvJqLToF5NcPNLz1uTxhUz3kN/Z57Zu7cpI0N7v7NvaDfqaDbU1D7pkhOI5HLaq
4Y5L8L5/PyrhC9SirwoThgiPzxgk//PSso7lg/voWKeR71oCPfAtZOIyUqyw5tJd
yop3VKGRwVFJ1ld9mug/X6SVDHo37UDb+UF7tVGOTpRZ0LQP73SGpkeyZWS5bv3/
IWCK/KVc3gdKtmKRnnpxZx4kjzKsU7fQDEK3kYrZjfy9byXNSzzhEOTPFmoQeQDb
de2Jg4b5X9P5GzeR1V2baWYsPqrPxR9Jx/z362P6bcLoOXz9FllYOhqeRBPJw0sE
lZo7RQMLiIMrO5OpwX9bo6AZWdbSeQWJs7A/gBLjIrGxnHO0HJnD3JkinRTHr26U
vXSqbdU9/JGxkHS3Ps0hOluC/G6j0jkvAS8MS+5LOjGPEFKbchMHWD2Ygn89q7jy
3MMDsUy7ivvDBl9iee0HtwflLyIQk6vP4BbEJuO787zeCDcpNa5yQs5bvdV+sOle
DdFaOcjQuQ02qzJ1V5q0EgMF+zSyOFwtuDywKNlZPuZIuO6kseNpvkL2Es27kbtH
n/uoHwMo/1UPY+4w1DAPUrhN2AdIS8y7RDCDBflPxD5SfYaKw6rlmu5iPo+pSXhU
KK6PakEe6yqy9OHroAzinXCOHiQWO3EfRb/XP3WQa8flhhO0DCuxU3XQycJOfsT2
Qtaec8CSOJWSXn+5R03bfCWZXg/uhpjfbh2+DwY3kykhiYzkM4/S1QJjtvNnjMr1
a9L1qDCAkWHgv55XnbRPSiSQQBB6bQSnsesjt1IU6AmjtVeUD6p+ySb+5BqSyAwX
i4VJaqtIX8Hhx1n7Sdw/nsitWCxA8b9xxrzGnlsNAEkU7sHvx8oWj5IEsxpMMTJU
8/Dm2jQROT2BgO8IAjLPTdyT8au0dffBdtwUIXfbT5HPsfUEVlYThbMetaEtuqKl
P16qY2/bocqUaBkUU+HXLahSTLX0K8/QqLeZVKhSSzz9o4WFQ+6aMNWKDW4GQWPf
vubPiWYvytQpGgx3ZWTkNQfSNvwb6PziQ7f5mnZ7+4Rn83ulGp7VBUkytd0i2qAy
g8uJAPGYa4YZcsuS4fCKhxw9pB3m+VAuHwHh5T1bAI8oK2CtdMV0q7RBKoBJfUwi
ILE6mbnMcEdY01njacGq9RZMfn7S1sMiC5vDvXyckmLlOx1xXFo84xO9MCpUMGPT
7YJ2ubVhhFOWF1gZ3LQdrRqrFjnbZIwnR5kDC09E2eiIMw3H6fplWQYie1tLv1Dn
TGHLP9ilvI0PePAzQXwD1bMES2weMQoXlV6gwo9pZi1m2O72tY8Ju0X+kN8SDRGU
V5+wJ37H6gnD1yETHHUGZSrHcRkhbAbAyPFZdmCq+YXzW7ZWejPUfy5JTgnKKJ4G
fotqRoP+sgBiYwYsZN04HpAvGSNAFAhw6OsTYEvzmT4pwcPqtwvdAmQpi2tZVR4c
6mbfhmBnNpw5SJhrOUZGUxvQDUDd5I7nc0I6IrBOvWVv7JI8Ica534YsR2AvWuiJ
sU+tqMd0ECJeFgAYC30vQ6yg7Ra42VIPYiPTrCoUxEiIGcRmWN07aFAbiqxCTHYT
TGS+sC7YrAML3ayDDxfyNVReVHIej7ViE3QH/H55GYVx0Kp7Q9558i653ppp15bK
gxk+m4mZkh3/BRfSieJ3Yz6QI7s9A1AT/IF8MPFF1PM4OtN0awILNtMmeZwl9dUN
fnW9vs5WRILWwwfzPzaU7VZuN9Y6k2MKSJffa7v0OBqV3/mu+YdtG+Cjle3owqkX
Qi7mWfBKQzcNSNLxXh85wMMd8H7CDDUDkQz4BRrEkXrGW+RlG9khc9KIUJpCuAQ0
xoJ4rCfWnvtqAX7PDClEr/GYQ47A+kV3Mazn7rYDN5IkMfLwiGZBSYPvF0xLZMdw
iKNksLhX0kF+w4qZiqVdfkaQBl2Ww579k8FZ57vyUYcMG8qWQEgqGmRALq7T9M0U
p5X0aS0H49FUVPxwIXa8nZg2CdRcslqcTI102GFKKpF/6lWT3qdhmlLkpzHXRUsz
+UuT1sPbEUW4h+V36NHcE/97pTVSL9PXnfGnUu4h+Fqx85SB4dY8IAfZPzRw2SKb
EwkY0qRUIIfLJ5MGytcMCj1ImtvgINxPsCzxRwAN1vwOAwYqDaSeH+IflXGxFxvi
wwoQGWP9HiSPav0LDoNgNWYtTjizywDz17yBm4qAyRG2Yb118IKwdqHz0G0qW2vb
xjBT1hUb9EOO+29iHzSun+wuhJGKZKxnk1pC8jY9xtLd0DWLkfI4YajXbA3FRjJ/
NliHpesO2yJsVcHBySaj8OTRN/Wwo8rfLR3Th347NxWB7sjJ0QRIaHv1fCq6IDpz
MNM+9L/MVjvyP4bJpu27tZQ4a/g4d+ogpsM2vcnbkRPdvGJ5jRgqQvOWBtxGEAUW
kM+odsM6pKTcOlfOjK7y0eW87AtQVkWtLxpvoOR+etC6X+BfOIc7iiuPMcNpGV0A
qx7vNVOije4kOZmUAL+D921eLEnH6rxKo9dtcb67bLBklhD5lD5bfcxzM3x3gkjt
SWr/WYVdj0hjqoZEhihZWqbs6OwAcEI6eRlTa+hs2Y1lL7QafS+ycsAOSGmWZzC7
Vq2p0c16EoUQy+O11H1jmHQvHSRT8qE9FXapQ/4+K0vPIiiWWsLlKK3rh+3S+GUr
qL4hsWOvK/qRnPoU8oa+8TZQknpOCCoUxY4K40cuapJt564UFz/b/Ym9yCpeDKFg
ZcPcHqLqwZ+HGYuFDfjj6F19BEyGOTuN8zZUWv6E4vUJA/C/IIPvmPoZrP2NDTyh
uEf531nGKXkaI7cVY+7EeVsCmtTp4DXFHHLaDBC1UJd60BzTgi/iELYukw+5mcxD
BXtgGcaKRA5h3Tg7EfVMsUACHJBoJ8Q84X0+N7B1a/m31YLsunur4ufrcN6CDUZ3
niWLT91EBOTOR3Y97CQI2LKl01JZ6XopoPWYr+dIFmde9xhU/K9cRS658rinqpaV
qxd59FAVIj1FAKFkpDLuPfj61ZzlHBv9yRN9SjAlCRNN4KBVvdQ0DPHvh0ckkI9A
QraSJoTwKcV55gEWCAyn03MNzo59ON2oj+CbhDUf15v7cEaq/76ot+q1HmEpks5i
U/5zDqVFJcAigtBIc8bIUk2ETMtrhrThOMzeKt+K3zoXbN4eU9tWKxyXcN+kQ+zQ
Bui+xkUynAtlcdS6Ou8euvjlNT6qFJhPbpTcJwrqeIJTeTz6mZaLbU3ibSIV2Kob
6ibeRJ0tAHIIIWWnao2ucY3oc40gUKk/9nnp5IuR8BmyoA87oeK10IaJZNmQrlJx
Tz+gecRhcxfHh5GzxiabDw1kMinsVSNQJ3KeCysdTV6IhGrPRMceClurs5LvFAqM
yxTpkYOXfhe4DJi3v1PEQIfDlMXOBpajjKMcPlxAcBsk7ThUCHL38uEETHlfDTWy
UWaF5SakHamGzEJ7T5tYTEPoLNvdWqfenjNgmh0ux1t1gtv2hTTb1BHYKb6HxBMD
dRtblqeUypARNwSgAcNf2d+WTmi279dZCLw+g5tJTyt+4Am3q5piyuKDwaZ2py5L
5c/2POLN16eAYpCdA4dtNvxmgv8uiHz2tvRwmGEoknw9Ac/NGlSV1EfllEF23kQV
e9CvGmd2jYt41FzvCeYHO9l5tEsNqRFET77Wqf0XUTG5OavvSj85M/HMHOkEyHg2
2FnnILkBksKXzJAISgorUZ74Z3w8Vg3JN8GPl9JJhJlxq6m0I/GhJ6JHBoj/hKc/
9ZSRH0nsJT6px45TCxHNB9SZ55IQ+dI0LkQZobT0jvzs50fNkptiCDC3aQqhFWLH
5u5g2GhdcsvSOBdAYkGiOPDwJnTYVdS0Gap28ttei9w24Klht6Gb+FFIzDsDqNln
6SUoalRlUNqjBxB4qXkhmIQvKUd14EDnwz5fSRzi+qFwHK1sgcpiSZqXvSrNPEKz
tleFfrqhfsZQDDV7IfpV0NuZx9kWZfL/znbu1ek01+kkDh+9UHLplMiWBMwivkVH
v9UOefJc5Ng0p9MiHVfWWASLyamq0a6aMvBoz5XhH7P7KDMrGh6r2JqXFULOVjBR
plCHIpHhBy10e+KC12VhklgrynWze4fVGlXtlGknzSn6kp8vIaqcUzln4IQSJj9P
LikHlLkylcdSgYgid4bzU4k5VpwXzr6SOlN4fCA1PIKrI5vsl4GC6E5IKVwjuqFH
Iv+A4P77JEdHUNqyc+TE6F4t1T+VJNbKqTbwT2reVFv9IuIqKKrjoZcz9X9AvtAd
MhOeWqfmxV63pIbX13QOL+Od9fVIGXQJWCnCBmdsd2DLhp9WTxddprFCa4fZDAyf
MfyyjJ78VusuLxtj0FGQTSwA/KrwcdK9QUCcOYnRPYk6DrTjp9J1zMnxhfLUBvnF
xaTd+Obk6Zp5zSem5p23aKE9DtqJhuiCdAEHC4PE+rqmcvfF/UpwiUQ/m0+vAzHO
AjyNRJmdQcVSKjh7CQv5Q10uFU1+B0jkTMYcL4oXPSh2C/edQwq6RXnoBuFLWQr+
iPDFw+lTxQOCFDafcEpQ26bsUFlnVjqjitJYSmFRaZ/WYtUfb1TjFfpvQhAOGVWU
3SXMBQjdHnE2kZvJJZW3W4Q6bZJYm4xcNbSgiDf5bZgnvdIdTKWV8ggf9dBf7Wcq
oHExAdKrfIJa6p1BCk23DpPfFqt1UY6wL/24Kz+3lGpgbG/15njyiCWjB4+AX4rq
1CQQvSIaSctQk7Zw++bgFsHEeJqycYXv9J13Qf/dt06/iEizna/P3wN+72BtsFBT
J/zq1s+LH7S2JJYxe/qdhHPKFQS/F+Bt8kNQAJmmyo59vuoV1OJVno1DZ+hk25gQ
S3i69nxag4H9GddWacgVjfCQuAJNE3SxBDiU+QqgQZpkoqsQMBD/dsLZNV3tURMt
Cr4SZy48CLXppBwsCCW6DegypiCZLKSO4EmuxuFmN+1/JzTudgwo5iZfSkqlTEe+
Wym0EDGDMRyq1TCYhz1UOkHKU6XVnlyYgk3zSMCIT5XHtkncxDfqd/OHc7nioRzq
izG3PoWRk5wokMJEiKQBIloPK0UswGq38YfUunntqeM+oAeF1005S9mYR1g1+eOm
M2gYXsEp+LFMo14ELxBYacVgIdeMR3zn3VV2H+O8qqIS3zjJi1bmfG6PyqTJIZDv
aR8t3E1Y0O9OrBeE1OgJj+nWei2sUOpy7gA1JVfIq3S77i8Ckhv00UOFJUvuBYeT
3ClcNx8xCwRl8Xc0Q/wGEzhdJHhGzqiYUv/fibg4nuE6cj4QQ0gQBh0bGPCDGqNr
d+OGGAVD5TxUOY+o089v435WRY918BtIjSyk8828vQCuzkeW/M/IBIn17UZHiwEM
HVklxbLLUVMdNLul/H04TpT6ABMS4O6EEVJ255lHzs5TkGZKaVPZ+R0RdCIfTQDU
noioLeJaKSxFIdI+KaJ0gQTC4ALwE6z5Pw1OP+33nflqUILZFqGOu/q+/x6VyeH/
7mcqrXdvqRPOmZtn3MUrPwNKc2fXVGBDSA/CUu5qi51QVAGPUkKtlE13SYa225Li
b7no2jKwnqGOLb4jBmEwLXyRwhFQWq8d6Be8X9LAN5ZNTjDJVc+dFHJxNjZVwOhy
f9lXj9FR3wTuPLYi/8mMbQIJoTrIfXO3BZ8RcM8Noyj3XEscEAnuEOBYjhfnwoeI
a+xZBsfqXDPB3claZOrAJ49xYs3CWIiIZJLvp0OfRSKTBMQ/sPJfONwMgzO+K4Sk
1jEYGzV51OKRVWVrs3PM0YLrcsGTQUDcYLb8rJbcLA89RD2AA/gQ2PgTliTt+5C5
I1T3ZAiXvGfpOsYW42Of3uOpf82Qt76mAMWv/cGrm06SMOSlz73/fX+o4oPi+nHk
5P5uwZXnFFAfue6J0Psi04fRJ7iu1Y1WeB4VqaFttJz/G3t7UFqRhNfINAsYkFBC
tL+KZxysKH/aGgV/PJHz4COMypzh39We5BiYzv3ntT5jWCRN4PEwS466TF3pYYZN
AsM/vcUaUjc2E0E1z7MMw8gHPsMxYwGHbX6dMxT59OJ3akt36sGRwX1/oY8SXbiw
BwQFvst4rSyiRRGDrTRr8WhlqLnRPv61om49flhHRUwh5ZhBVpwkXlTy5+3LSQ1O
fagOJDKMhjcLddPXFiaPw1bUGAic73Pa1o8RaBai36sHaXr9B37H8A+8bG5zNSt6
UlA8vJJyxJldA9nLUFRqVkY7WXK7pG96vwIenZgUU4p/Kpg1+g2bHPHrKUNoTgNa
VeS+IWSfyO3708wKTE/OBRonLZpeYgdH9zA6x33gw+hRcCJ7SvtAqigl5A+Qu6lY
m6W/rQt6JTDG2CSSySokDX5rcR3kveWd2Oux994o+L4wk9/XK/T3H0+XzZeEJSrL
eT+EickWF6sxaefeAHYJmjV5DdEeLqtuied6cBHloqTAwj0NWkb81QrxH4mAl3yW
AekHELSOOgVKegJT8qXeAbhh92/tDZxQU0BpeI8ML40du4CVqH2ONHp0cuRNCwHl
A/WG54ooigCLW9z6o78bN+dQ+yvzwfQU7KFtJvSKL9ryriwGFaLQmGBi96tDwtxz
amL/cmcdgaLBxQTA5ap5+t9xiSoN7inlv8a6KJTiGD9Nbl9vV5bDhaquYra2ctOB
o1wqsPSYFg1cVPD5Cozt2nfSikA1bDR7TweQeczaFPsssSEaBQMwApSt5a++39KB
kzHRsNfYKaMAy67m+SOOsemkYMSBfKuAYB6GHEwAIep3D+f76B5U1ltU0DCxE/Fm
zjtPIuaTT3zCRod84iK6Be1QBaEhuMnLnHihYBbikl2LffuBzfcdQuYNFWBt6EGp
seEMDuSBHtHbYTskkmG/ZY7LnYqADRq7i1DjBYZ7pkB02c9aLNgZ3MlhrBrrEB9o
Nt5E6vH8X9KCV/wYnluuYMVynuk5PKxh7O2YEJVgUumYqVLUdsLaEmNfGXRpOLdz
QByo7EpTy737ho83FoBkLVFXniV2zrKrkzBrVGshZA6QNN75vts1Nh4tZfeD0vJh
k9dCVsGraKPKBJok7aCzCtjF1yys831jALnoTXZyyQUHXLcUnPmMONw6NkxT3tvB
9NABf3A3pEyqxEV5LgDSbeEDHth/vb8clIdke/dS9AJHgq0CvzXuKAPrHMytWS+/
6RStKyVgi3/HnRPJf0PhEaoicP/stnl0fLnq0Xjr2tKOn8CGp3ainQ1CzjOIuhE3
1sqD8YVATuGToLJmAwOrGx+4RUuJywxpYhjrnFH+SrjkmJOwpLCgVEOwiqsisA3Q
U3oJGb8aWSUK5t1e9V+RiOi819PNmJCZ+w0JTpIrevTUK5x2j4AiiCy3QEe7scXN
EpCrOhzCbclhctzUy8xadsgvHgn0Yfvj1m1qoXLTGYsjRFShyIM43mWLO2obHK2Q
SZSxHNMFv+Rlz0B7qlpmk6QwDInS5j7ocPN+Ppc0FA3iwyEz8vWZGnGcXK0GTLah
QRv0b9CewBLb27fTRzeqv0yMtHv6wG6oCWpc/uAXySh//DGxMRX4FXMEaSB7RQej
XBKLd9oYVJaVdHWzc8mJoBB9OHxFhInJc8qCXwpVTv3qTSpDagUE6gsGMnyM5Ysb
AEU+hi0AtuqHgBTfDi56/ODqJRf4oFYL2eI8XN6l85RDnoss8YQMNTavX41/mCFJ
aDoFmJQwDyJamHLWM+Cd5gwBAp8ZVdnTAj+gz965DfWi9yggT/lTYwb58vlZ23g6
/5zv7hIypMef7mHM9CnNiiCIUUD9mNLM7KKT3RGGHrmnWQtfDb3JCt40ipq1JjWN
CaEUNgfJ3maD3hmxQ/YYDZm2216uFINxihVGTQ4/WRzBpvkPVbQtBf2H/UYpu9ZZ
7UOY3stOb97GVb92vL5oDoQaY3vhFtLCoD4oI71UR5FZKJMAzZWUErlVFPmntkod
XzBG81GAyRVV7f8USUfDno2PdjdYTmaigP5Z/62kA/ARDbA7h2H2o62g6JvCrojO
NpcPOqSZDAB8fksK/Tir0eMfPY7jPKl4d20nDdexFx7TOloZD3NWGKanV5tKsPtf
GN11x26McOl/bEmKKYwMgF+27RjR5e1LywNQ4CkgCUBBKWcbW8ErvVfLu/zf91me
pSSwXbBL5GNiBIq5PFc8hSwC3hcjiUZe//Vhf9ZGO206V4TLlOn2j2HZ8jbKWZXD
eLH4pKdIjLfkj+TEAyujzYWJ4h/BAn56cGGRzQvs8bp+PrMsJ9jYQdLFM/1+Snlg
8K5x1VKWzIrp8YinrDnitpf1hpQn2wYzZJ3wDVQrKc2cwcR2RfsdLdIL2kJ8AzrT
PYO5jSq6v+QS0Zp9dSseyYqoy/vRgNrpIofmf54fDMMpBMvF2H037xwdUIyl6r9t
hDzxeSMlKjK1b3/ewq5u7wxs2radvFh7VzSBbuMMfHmedPSn+qw8A6P84GcHQjOO
aOf9uzrSasg98OVYJlL0JEM3vaIHaT51hdvpnUVLDDFZ4DRGGVgfuJHw/e4431Sl
r6ynFv7z/o+QQxX5QcBT+a02vhz5ZfYkhL1HkGVkIaUUB4lQdgsYPdM8/oJZRzuk
xOJsOW4Xf7QRjkea5NsLkwUpY11FJHu2SxLWfGfXN4Wdj7y0oS98l1nSlwcsSDv2
8LaVk4A9Cg4NOPN99KFUh3FEu4RvaefJw8XsFyzVZipudoBurbhwiGLPy02y+pa+
p9A9FXLhDuY3viPwXhoJ+v/V9JrQqScPkI7fEti1fx3pfwIZ6DFDo9rYGI4w110t
Hjmn77AEC3aL3PBQ2nrWe2v73iWryoHqQzhnMgFXatb0pVnw5HmgC8NFFKmywkUk
bbY2c8W4d38TiZu1mPrR4iAC/5W4itiDSDz+zaqrqnovZ6yZ8jhgxp8hcq33cNgz
LIi3n4a40io/qDJK3pJhojnTSUinojxO5xPRQfqB6vocUd+DFjHw+bTzNIi2SNlW
AlFicqEBzdfaFtdqJXZGXgVygLowzs9QT0qdSUXlmi41N39DgGKU7FWua5ZNFLa+
V201vl984ac9m/RWzE4JvwQnJDiaaxnSFxZYtrPCdei9QQIvNsRtDNvORc224twx
0fsD0j1KZIcNvqp0ofoVsZXoh10bqm0ekdsRe2FSKs3u8Xjwcve1b4yLOcEvGRSv
HMQ9v0bi8ezKWNQgUCyDRZ7TTM2n1QZIGUhPH3BG1rFdCXaSHpQUYeYBRZXGSFbV
pHIk2PQ8bEB08BpNECBVuRWHYWotdJWh5SQSkPRPcIooAwDFcglTDDTWPatqPERi
By3szrvviDDmBS5F2/pYRDFJwCdG1SLKOoYPpSIPWYUDSjqiUro/KKPaaGtkXbp/
gXCkVA5yWbSbOYZEe8TXOl9jOm2fZZe970fdDNqHlxRBFCIdvfpe6bx5PlYqZuGS
5EYFJ2pYf3Sf+qWsKru6H/8r7xZTy/lfaCNUebDtsBI0bbX2y8eNE8B/b8gsfJzf
0UTBeoafYyyW81kTwI3mthwwJtPwt6qOz8wRNWhXnKpIgW7OHwJyTPki6DyjRpWD
96Zy8NN/KExflDvYrdrDWXyS4E4ipJBWtrfu5xEuBVrs3nebPQSd3nmhfh3tN9kx
1n0lHfUkMgG6bjWcSZnkKgyIr/zSoQjF1qzwL0JEK8Sbv8K+z3YEyG+KiB9R5Eww
KHuA69p5k9UtqLWnzzP/9yd91MCgRC9K9WuHvuCATN80u4iV29RpKquISFMdMK9O
ysKD+a7tRTNtFAx7TMBqwdbsm2pJ7H0ugR80nTQhkx87UspBynGNTCUU7OKSU6DX
+IRZYbsXH2CeUpdIcB6bYLP2nhu5OZH7iNDnUkZILdloVFhYavH/4n/gRCGv0nKx
Q+xfKpzPdlPrZjeI+/YdKPfrutgE2uGWY1GFrVUIOYhvueBuWFRp0jLTW4Rc8s7t
BEsPwXSrb21Qgf9DokeEFN13j6kxXOsXEBtrJgeCFKYPGavd5KP/NhqF2jvAtvVP
H6RVdtymSSx53z+XxmUvPT8fpEUw9Z0joALxBLhUTr9WZkFs7kcb73pQ8ev6JH8z
VgQXofN0LL0/oAxT8oR77JSJV3fe1kwxZhMzr5ZSD49ukIswQAe7tYGjJ3RSVyA5
Ge8WAUir5bNbh1GGfAAc2kivs4/mS36/VNuw9qXfvJYuhwMlyHI8nRCrLIJT8kPW
xPY+hstRy5dz7QxOUmEit+gzvqiBb4too4duAeV6iezcHC/VvnPz/EI0bNmnoUB7
/8ok/76ZFR4LKXC5iUzYNbq/0HgUf5fIp22siNqJHlKo3n63JRpl/ttK6KfLfPqk
NTwwLA3Du3yVLG+rzNG/6stqvCXqWpd0mVxVKb+saR3XUT4y4ftxUY7D5XS0bOkn
FrwYKcemCBMdqOvb173g4veVijfFCW59JlqF/4vWW17oQwONB+lVk0nK5h6twx+F
30hZsMlqUe/C23rKhAv9FfSPsL86uIE2cm59KXlF8CwOfOBQGHtui0a1+jmcrM4C
1Xd9MQGYEoe0r8YTcjn3YcrrLpfDU3c52yatsJFXDYHGigaXw352IBDRog6xRiQf
7eq5SNHnIezOxPqbBnQHgYBLJh3OVQcY699It43swGCFznHlpribY9mU/Dj54xPR
kAznsL1sW6ite4CCHBa0m4N+dCY6LR4HBas6iX0XnHNW3p/u0WvRsaILZoLc9DXt
WJBe4w0LaW9gTc9h2c4eJXINXJelQhpdi+g9+X+C5W2VpvE23oxhzsptP4AHLOih
OGDD5TwAzTJ9FJ0k6of7O0gY0z76lfqmFylwlL55gtsnGzwU/XWtYdiggTdK5qw+
mJXvRFEwXLJr12vVrr+Czn9xgQU7NjoHye1452Zid9hMU3tgtu3Jn+GfvTcVA1hm
jSr90V64AryVGx+NrxGjU01ayOoqi5xYdIjZzwjjLc0B3WxtG7qLRD+2gQ+il3jy
7Z0mM9OxBPyHlXmwRBaHW/bqDuiVtcP5s+NEMN8frnMFLe0zQQMfkvKl0dhBUVo4
bFuiU6s5v1JHjGfMcjM61zPvBy5BoB1tXB8kcz4IBa+toizIEJLiA4unPT+qi1dA
ZvF+iviyy+6yPmi30iI/9CTclD4b3cAtTBRDiAqJlO5QzD8V8JGiztGrP3UzSxAY
KddJvyxLw6y8Qe1WJFVSWFYeD4YBwi919tTF7fm/9vSq3vOIcmT9Up99wDo953UG
VVPKVQeVmKNk5wl0s2GJcKriWHrpC/Z/QDpnwLg5LY3Mf1uMLBhl42c4j9E/ZzbP
Mnq85AU3zZwNpvS8Gw86Q5zit79H4XLbjYsScWc1Mv2vLSDIXNakVmmMjKk/aY9D
pw4qEvjtUzNbY8ZmTJKJCYSnEPKLW/IR904WeMDBgEO+J5hXwiiFbXQXvJCixRC+
j8sA5b9Dq6gdsseZd9+nzoi+fXl0NsTXaxcP6UprxdCqlTQrXAVTErHq336+fYGq
BlymxMOM3BPM7Iw5XlD7ZPKj5qGrnFE/Y++PuOuyxNmsV8aLhEKF0PWU8gNj56rw
7O2iJ+5uBECqHEKpXPtbYdb7UHFF+BR0Hwu2wlMNXmptvcbYKn3bnjk3tJQlBFIv
evCPMfZJJET3txOySLheCgPDmqnf686bVfaO9MZ5bqEOulCLCG05nMCztbSD3gBx
bsXnSj0ffXkH3tuLBTP2RoCXlVz9lF+TPbqxBj9SGli8hNhn9Z3ImSiQG3JKkDEu
n1Tdn7tQCVzmo7txlftyQCCDUDPcjNYR9m+X2gLUQMEjbTvuX50JUzqNKQq6cgC3
iUmD140BgEFVvNhgmNWeRw+Vr2MvsCuTi5HA6v69dF8j9c+xR47rNM4iwYo7N/TJ
j3ilQVxb7/A57JQz0TaTZAzItBp+gujJt7AYvkx9cSjj+u0VnU9toIBCVZaJxHqL
l2t34fOMhrnp6FZgxIlffzXErHkPv5xjPg1oGC3O6C002LmlrlA+xPKXtdX8Dvmk
JMb1wo+WpEVWZwWzpF5j/uDUx2etrUbC/hAFq98vc8h2O2qRubieO8loH0Kh7X4s
drKcf4rZVjgRftx8vpCLMbEG2lb8h/dYQZLNq8t+zhJAIe7vtf2wL6LO4qBv38Ib
tTfGF4YspWAZ4Y3j85NyQ3sK3Mx8Aabqk8qZTE1LdtoF7Tjx8CSgVe/G/CXdjsRj
N0fT9bPa3ficmCyZbTzIfoKD81yjfpReseuk6amrlcHnbV7vXBnWDL3GFWtOlBz1
G2FSJIpSApKGMJpeh9kKk6cZv69pHNqYuTlU3WYZeKVYvgElC2HdCVh5RLSzjhOw
9WLZvZ+lar2ncVNvMUoXq3P6jVoL3SYwa4Ikxr4j7vuB7rTn20QrA8ogXKz285ko
X9jAQzKjaD9ReFMco/jUHzJ52PZLj4qaLwO/ATJE5lufIBk/nexDDF/JV6savNN1
fkMWgJFkCb/G0CBFYoPBLu8AkOUSLEehfbT8C0ZbZcX9F+M6P95toShCRNVuUDx+
ZDQXnoRu5leGJHbfh0+6foGbcPrHyTkV9HUufhhSs/U3+M5HRIs2i64XKZhWSgcL
LD8teYQ1tEiMY1D+Z5yMVQ4Cy6tpRAgJvhGUTnWbvAEX/MoWA8AHuxke1jpEUOFz
l1EdDWaLat4OwuSHPHU9Z9cahJelW0ZN4gFOWFhhLGvvYk/Akf0e76Ws6N0F62Sx
W8FbnToc7zB+b37JFN5ZsnsddoaejACdvK7T7WxnHxlrtBoHjjg+/8ETbLjufD5e
o/Wjlax0zgZMcoCsc8yfAZe/0xeocelN1NMtMbxhrkJnTI/RnSZ7/VvmbCMXrrYv
SmF/5KWEdy4ZBHzaj2KJ+tVfC9BQNjUzj9xre3I0Yi2aIZlkw0+ZqG+ot99nQSdR
PjZwEvcif5ySaoDW7EUcM+8k2aw1ho/xOq6g3mygMsONA4susD16QzKrvipzd0+d
o4sHGTHk/UGTLmlDz/SbDW0MI1iX1CUYo+1lWe3mAoXQWAIcMUFYyWEHV2EY0i/I
JTIryKmsk6byAaeiOF95THBboWDgxdKvNaonsrEg7HwiOG918lH/HDeGgyDOT4tk
P9IPQEbkBu2jeDE1t8rbq7X6JuOIvQIpnaI3PkErTqYrK500PrSZjOkpy/dv8DOF
oW2kJWFeiJITROjNahno0SwJTJsMv0oeY6wvrC9HmSpfknER14mL3SnGQR7I9ZcI
6vOD5RNayM7PI5VyY4EFVbNtmlVdoksroEe4gzjIz7A73Vkl0UFDUKd729uSX5Dc
MF+ezLiH4FELncbG9kYXlNp32w96Mr9LIlnqtsVDNBcXBAslzE2XZOsLPNmZL7ck
5hlE0Hz8ZmwwNI9s1omp5X/I9xBPjrzWdgKufIm2tDjwi2/GYX8cVaPcvQ5Preqw
3Lpexa0ypxYCZYZLdXp/XxwGvWtAjNRCXlFWj5V1PcEXeOWrtAn8lVEPfpR/+892
SPBca5hsFHHLwNX2PHYfjRiu329uRj0Opb7R6TgTrV066kIQ/G4Jms8mXLUu0107
TFdJ0b2T6NvgNyvoZnoKwbja4OGfD8ft3Wletnm70nPaWetq0VP6AHbuJvG+oqqD
6cxCrwqNTQLAc47avuqEFE+bflIWd3k0CyFNCaSIdKituTyEuiPRDIvytZe+Vh3X
v7xbIxJ2uUG60zZxsoe7/CQusLIi6/i1eZrpGHqovQ+A169nhy1idHEsTRjPkrJR
zpVUCErJwuhVVEIiAdZ2jSzYWy2o+6HMYlMpqgLLSjIl13Wju8jGShT8fPe0xNOR
2zWkCWUKh7c+Z7Il+6pEV2WxJMFa33St203Xo0gbofYZW9GA0Xyqi+YYibDXPQvP
S3uABBhK9yBa8s7W6iXjvmypcofya2kFak5NzzBr3Nei1lGqE2Q7QahKHiGLrrIe
pkSwqqcRgiEvVfUE2BeUF7OsdT1qhHDw4CWx480+SmLqT0EAeIc6j/qttO0BGrDI
sQQ/wePZfochNmagTHyb6/iOw4/IsSVRxjT2PnZ0Irua733CKVy/7uo3fJJKgSnt
cg/g2liYU73FQeHiD9LzPoP7Op+/LlP1/1UMUD/+mN7P4HMczvVPouiOHn03gBdS
oDxuYEhsHV5wveQSc5NFClIsNy1k1SCKt1E8l7/eKXmUmrFSVCEfvDpFKaOb8Qyf
OjmaAcvCozEMusThDdFRMQauWWfhi7Re7KGcDexAibv2cZZJfvPzoyIw8/qlfHWI
LSvMiufxJTF3nP8DSKUcUBLxw3CvG9z73UdC7OMSOLepWIjuZtfgQrwYP3j9TtNH
//kZl9YZUA6g2PQejaEyuAGA7zljrsCRNlDphmr/YMpb+gFb9tLqWH23OjtdsUSb
z3Mo0qmShT9GqHobtwTWjZYJGoLeYupYNoEcSOwOpJO1MgFaPnwgmZx/eeuxW2qW
LYgP0b8ebqffGqGJ5Mwcl1tD/7PGiY5Piwn/Gwr6QPVzMcvsVnRlg7M8rOG/7bzJ
PFXuFVc8bGDOR/0i4QARdjH4a+Vrf8x0sZJcrKzUWEaSlVAQXSgaA2whGw/z9DyS
KEgzsjC8utkajmJmxjDpBd9MoUqH6mMAeZ593a2NZ53Ji85fwQ8cTrQzkQ6+J7n6
3j6+8zOAmntpUqQANxc68Me5A8yhHMlZAEvAVw6TjHnmP8pX40vUiuxRs93EWoWz
wB65DOp8aJnZKyuJB5brX47UNd3af1IRyfYAeP0Y+8OIktVLCNeOla5/AjCex67b
ORwrbGORI3bv6QXNt6B+JQh3N0NfLge2cHoRheHd0FkCgzoQubaQ+HwbmuQrac5O
WuDV7OOmr0WrCBJKQPhSzIgnNFoHm54bXzoqYfCb8lLlTFAJxdtLipVXNTg2qY5y
tdaU0b1WHR82qgQaJniTCyUIHo4PURvn2RTkiMX3QO6PBFy9tcurmIiEPhhGuubw
FBvipv9obqGgA7oayn7XQiNoe13SpHS4e5GcUo308ZvXxTwDTM47Se8F9B+f/ojc
0xcB3CQxUilnhl0kOiv07dbNxEp+kEKEAlN8xitYAWRuneYe3jmKv42pPtCsg0g/
Rd6TmbVw+QdlbP3fvC9OoVDxVSPCQ2VmQPWNF2nJnC/+t5n3XG98NnlYi3oVsAdd
lNPkY9Humrwg71QGI83ikouV9pnBHuAS776dxyZQ8gr7J3nyEXDsoSGkqOpSvuxg
8pA1qyezlU+MAgSoild+Z+uSt5XSCTO2HI6xpLV/t558rQRoNXl1BYnlggCPvVD8
chXVDgdvrZ3GwRjwkebJRCU1PJ+j0CfwexFceTJTkkIWaYdqj10U1eTLw+7V83Lh
91vCf0echVEZHxkgCf0BdDuLf0ggOSFD1BRznXH/a3h4FHaitsFinyhypI8wdsuV
wYKm/AZ7TuXABoGTk8AHmrrZhnOUKht0+R1OYjiyeTgHqbUoAhjSGMxN2V2QaM1s
afeoSdETqamHioAO3w51I6E4qeKQNPAlW6fR9I4xQaVMcpA2tqmtJM78gKDuhUpy
Lg0CB+HUuE+lmU0vDVVdVgTOZ7IMTOh8ZLY8strErSe0ln0oG87EzzHsSeLd6OZM
DyeVZHW6T7buuMUkJIqGrbemqjc0FJ9oNCtm0hoAhpNqNuDQNkZ9PSFLsbZNPORX
kE0xZgY/D6yeaihZ2Mjay6V0wThVb4BlocUYartHnzYl6vLdAJOIBNZHZDLys18i
fVO6i9vZTt5nR+dzlRqtLf3I/8aTXyco638mToBGSggYnHHdmGgCTnIGasn0B8vb
Cn0yl7O10pCfEQL4a4X4JJKpqQVLGRX/toqWqNhGsSpBbT+oveeAgItJhnyKKRe0
jIALgaqbiHw7cVcywlLYNTtKVwyMM9ZrS9OrJRpiNZMcXI5iaNZrpVBdWtkF0fch
3KZI1E41BK7/YxTufz9DjOasPLkXCqWEhlIsDWPYOSEJhvIUXihD0drE9OspeqTc
q74i2SnAE9wFYY5/DQS8EkNGdPI/52JyLwux6pNVSm2WKRB0pDVzkrykQ7qzI6vV
0LQRJf5iB9I+v02XecT5x2B6TFpWp9+nSj3kFv17I/UYMtOMga5h5K6vWEMjqhVQ
2iPlfm6UaSyrZ7sPccHai0FXkXCL6dP7v6mCQX/QSkj8UA4HQGmSzDcd+7HJBAtO
32k2Jm+eHIpzfiP0eGElat2OARUFA1xsZjLazrVDIuyW/jcbZgW55xEyfopTUeUq
qM5vh8m0Th41EQWO6/vpERfWox26KQ2iwgch/AdG+IoH4Z/ENPTznB4TBVBQ2Jsz
ZEX5yk3rgxaPToQN+5TERItmuHA6QfeVTIazdVC/5pMesL0xF5yxZrbkeNVeRbnM
/bLCSTlcr4RYovUx2Y5tLbfwVB8d8Wd4MGl13itPv3yIo1rLgFdMetUCWCWdxJWK
Oz0m2VzJmeDQHpQ6lXR4Gf5QUgiehhjmSW4KpGvJawTH3M4nKdClLIQIEgbwRR50
8A+V6V4UyHfcIkyhiT+4bTAssx2QQygbCb+vL0fb/QWd5aIggupq9LnEBNhTioKT
XJrRHPBuWnjBTS9Xq0B7ZUg3vNCCf5b1ZZ8H6vvp6DabneGkHfb2jtPiwDiH7zrq
m1RYVAkdm/Vf4R4/PStbiORznBqCExbHWoWaGDCKrKdHOFKoTXX6UDNn5cM5OXQU
q9gsSlcY29LSgw5d6NWj0xFnJ/LfI0e1ss4YMRFR/fVOherUvB69qV4q9uF+HXSG
EDh6WZHRWfHZ6kdnavAn1YF1yc+/wBtDh89yAbK1jc1sm0E0X4gzU99HR46qqbot
IFsaU7iSBOG1ytDZaRtzjWRfoL7LL8cHMK6rvsCgSXc0F7MhJrxF3iz8D3Dtht2L
A2b9LO+VE519pQU1TBaSQb88qAlhSOAOyIzafSDHiBksd49H69tccObPEaRb84YZ
cH3J5ZLvVwS1qSjxnnO96sy/S+j9lPh89Yj4lJX+/dnjzejCh8G9VlGNziNvXC17
nDeAkbvcOP6qjy6pqiUu86OxCNyyqCYxJxH8o5WYgeU5dfgA3TWWaCCJXV3OPlJ5
KvjFAuNAu2LZvfwgyiAQ5zChw6BIp87jQcHAgBKj9Rmb2JJ9MlDnG9UM3zBPyC3W
rfMIIdD+jcNh7XAtl3fAdsFv8N0/FzXvP2g9luSVDSKtbi76d2flVA98rC/UTzC1
vo1B243C1YsoX1rD9drpsZ+iiF2j9j9JkhAxqj5fE8iS7PFkKWcSGNxGVWmGS7zM
zFrbiCU4lAui5pilhcb6thPxCnBkfhmXFIoMzwbA6JKHjuxDHxFAi4GQBPmk9Bqh
mQbtB4vg0528RDzWKNQdoFD2Zu/aXr4wQapJV7GUd8N5ZLB3zul8IQCie96AhUN4
1Cp0E8nuyNnY1WGT2Mq8biyHkA4jaMcgLE+h/qigHStEm+sWiHpLufdSoEiCw3GO
nvRBh0qZfQms4LH/87Cp5HLUK/JlcTlE2OsYzREDnax9WflKUg5O3WFHt0m3+6yS
g/PJGT1v5lkO84Kd2bsLlMFSKuHgItDDuRaE8mAxtTvgcxZo6scQae1frx4QCwyM
pRrtA9ZcBzdbc/+YML+IcX4S+c/bgEihv9bcIkcENbOq2qGXTnteAK/mlKJj8Cds
v8deVFtsb2sETlZdu/ppULGYy1fVoTS4oWgotH0eP0ZIiPR/s55hfcA2z3m0KrA7
Zq20v/MQAsRUt6l+ZpYKUFEk2xX78OGTss8Gr64rjS2CEac/emtnLl1XpF2vpQkD
XMt9oJg/HBExQgM5brz96BogIpPb86ONu3aJKfB1hN0bSOOQJFG6vQW8WOzStQhS
eAsYd4YhIyESfsQVXQVUVUGmHD73wQibqYEusuB1dKruiFPO7nTGIRnzCffLcDYm
nyC29w210bFdbETmfTQ/gGoEBJeTtQR24+mdIypBd3HpynPWNKwAE9l4aP+//KqH
rulhsdJ6ARsjBQ/OiAayNjQ4Ir3zcv71WcvpAUy/3Z9RewKFa/MKCiYoMUOLMDw4
lS2lFYzAo7iksMpZv4heVpwtAp+18WvleGQFA07ss85UpLD9vjukz04ruN7Hq8Ii
GTR6UKadwIE8kXLfLbKzyYHyMrgY/PRUWFzTPsn2/VXxQ8yQsdPVJtZ5O4qj3Jji
RxoZ5YpOCbU9wce1Kzw2gmTFO8s02jWON5ANE2dro6HoBXAid8yyeLZokCrG8Sue
UT4raQ0bu94NrZOCo/OBr7HaGuU53PS9xFdXUbVnu99UT/u/22V5LbthoRaeie/5
4EVEdImT6dKbi0J5Dc547i89UNxMQTx1nizeFn4XobqV+LgkdChVH+oAlpuukqpT
Yg1i+nQB514J9iRh9C6TEd/SE79EDiG7l07gUp2gqwJgHlf2JIFlB8ce2jsvY/2t
YWOFUvDKnoIFUMOsLlfMj3DPrhHKqSBsNSHD+jVpEY0q3OQSHv4yjENOU5200qds
7BuV9G0Q6ghkTzyq3xbOZ3/jX1m9QV8kO+453uilOzukWSFZAi8/x3QDnhOLNQ/+
d+uuBHOO8EIHnXgpU/QY9qP8pNoTpbk7egCHWAcMvSO8XCEQ6y2IJgIX+qdDab5M
EbT/9nxwJVjcpHNvdSqOMfBas1hEzdniZVcJijvYkIzzn96vvJoX97U0dlErI8V5
VnMIWqvqci1ICQe7Bj17kZjN4+ANv+mV+gEMWcBXBnaVCzlag5KdYn9gRrTnWXMq
zXE3RV2DaGxSjsjOBe/dS5Bl2fIo+0ndhahj2NgJe70RPP8ggmof0lIQPulkVatX
cLd5YVpETKIZNYYLvtatzAHctRqzHItCFyJMmjjvShmpE8KKM5Dpv/s08j9F5OdP
b4WAiaFkUeyXiTJrU+b4QLMO6CBrKUChH8ffj5BJOOoO3dJAa68COqRBIkF2R51u
1KZu1Hyg+DOpWQsRt5SGvwBUgtz9s33+ZfV+yRnLYAXJVY5RG9tyPRgqv1MjqgQf
dF3ObPYBUciFgAv0tBMLsLN934e7qv6AKAaFwOvu0xo2AP9fz7jww4XX+aBnLDP/
byBFEOewAIEvDwOoBhxKmULEu+aMTpmFjM/1bQsZl5/lB/Aeul4PodApeQXpFDX/
aTkSP5XXMPDgbcqGhzfUbU2zGgXvkktatv+UOF0J+LDN8jlL6EJqJrPJBzWPyZVY
s1K4hROwM4gzga8zV2w4y9fN4gNU44MPQHakahkPJh7Hy9jDl5MUpPbXZC6sQbuY
7lK7kIU1CxVsYK4ZZ6qoxjzv1xZyRhdOpY5GexVVNZdCCehCtzdFYd4RXHQkfe/Y
pBGRc/lqZ0ofcrkdDm31iRJuASoGnzQ7+HM5aNjvO2fBTT5i4ZLnASk8Xvb+Ig7I
1DYYHlY+6AxbPKEVexkIRlSwfz2jWwrn10fU7/rt24DEertrZdR7xjK/HsZLLHz3
IkD6JdhzFyhnrWzrN7dV89Iiwx4/OtAUEzCBU8FgdiroaRsJn0KQLS9J0czrYlqU
LolKakN4NGFqPIhM+ZUmm1FvKlv9OyIIWMTLjxS8LxhJOVrt2eSv0hkD6EKQG8hO
L1hFaEGtvPjo5CDG57bwOlH/4UfTxte5xVlQutlBky91pY7HupPBTBoWXIufqTnY
LDfi13mCDEwombXP0+5el3msRDlett0rxZ90HniZpHBJ+XbvTx4NJzhnYway6Acj
HLvNwSE+qiGWyUCAXHVCPbvPoO4SN/OVmWq+6zrmVkg46He4hlXSqEmvIF1/iw35
GgF29AIhbbOpj3ZmN5pgEvp36+pCHiNnmrnWfLnzwEFYCpnOtuBVg8cBwdZ99wPu
68od2H3IV+byuwoRS7RxCDxpiEu+K7MN/dhknvKBEBgZrUrY619IM+sEu/um30GN
DrUQdeb+W3itrNN/EPv8B3BnRu78u60RI2h1JghE5ikyevKKqpVGJ0VkOnPlooOY
qM79yntcC9Tu8qeeEy87pcvOY4BU1axVq+9KPxdwHsODMFlHNSF8kVWmCgSKxJ4v
u8ixusoXiVH7nwCwZCSHGRhgLd3N9UfsSP/nH1+82BpqagiEZvaOecMxsT53glpP
uWW/h8y1d5eJVeskUtF7NRU2gWgRE++GcYURWWwtjCrCBm/1Dyys5wLJfhoqH426
5RjMX2yXThuuMEphqceUN0w/H4Mkk0LX7X4k6yjPKz5DxvoWVOMH1mmtPJpJwQi5
1a4sUYituM4InNM6Lvv72vYdSg3MNDObu9bveCE8PtFPmVbmlGaY4A3JgCDNxehW
/ENQqU44OWHzGk9nEEjpTvBboOttop05oyIm51XdjaEmZQ0PGjdMsBDyT/QfMRdx
YzLEUhiWz2fpfcRMvDoUXhIAA9OPrzqOFunL5z6UhKXvqDEl6HfkDKKHltlDFZZI
eEQQsLBCDX7OpVK4fv1wDuBYXMZGrr7nBf/1GottvSahQRkBCV74162+1Lgs8+fB
6lJ5v9oRtMTLFNku2LCmSVrUuDTrCZPbcsZC66L8Rfo/k20265iaYQePadKg6x8d
Vu7ra4OrApyvg0lFiJg5RfcmUZ3lqlvlFPRI2u94RnUMgK32AfVtm6oRwHNcZsnz
IjFJCNXnUpbxbwLWJFGRLCTKHQsvJRE9WimQg+0qc11Loqij5d0NFhygS/vY6qP7
f3MjdVQSzG9U4UhrW2MUcu7pF4Fn1WyJzkvV4DevceL1A1WTBTdEHOHcvbKj5Dlk
zvSMmzASidAS9EK4t4zr5Bm9arBkMj6ieEBFYrcobAiKsdC4lxpGtw9MID0jqAfP
mCBQbpV4/0CHlN9xHI35Bhe841pVCpMISiTuqH6hxAEoxLXEoa6R/vQRJGwXeeTt
0ZDL06okOAbhZPPb+TIqvFuNAKBpYCRXvXeodWoB858n0v3ibxiIc33p27RH9sWY
Vuu7TyVeBvXBGeuv9UFELix127mRhkUoOp9PqOHqDP44iuBX05V/HZxT99IlzQdG
YLjb55wqokYbjYwtQDmb2t6h1gDg0sd0LmtvnsfOFOOFTCtUQvLG7IHpnNyxkGUP
NJgg3yXnMC55vvuHyb8Yu0SJDlw/9+X8f3h7Q9mzJ6ogPpzH4bejtmEfHuxw476L
z+WZsEyF1sE9ZW9vDCe+EWhPxZaNXm/eOw5u8nPNrMN9lOLYSJVGEyQ3wjBz6kPi
FyWQBU/TftFCffSaMAKOgZMIAUC3L2YcJ+7hkPiENl0mFTiGBjpPTGPJy36Qpjs8
h8bF4OpIswcLguaqYeyYNN9FrodpuSo+Vkm4cPRwRBGuHtD8vBUwB+gJMB+ctD7+
9ex/oLHuTEdatLjlrAr0CT0nweCb/sNvs4hRtw5caynp9eDPr6N1eGQWF6a9O0SE
Lc2k6s0EP8E44HKYA1Wvnsrnu4g8ueXGKvo4A1uZnJnCM4mvXGHDtLYlcp2bl9tX
5kuiLz+EmvlSdYHg7fsNIFmxy0gQAho4BGYby1v2o8Davy/H0nKOWa6fDBdBWcrN
d8orSAex4YtfNYVvz4A6ecfrNpcNPDLHqGk0C/n1vw7MdxWdmV1+dXUiPMl+GQLV
1lOBg7+QUc/OEHtS1ZQfFy7Ps34ouywxSp9zm2y8GIOGizgC8xJ09CWkdF9NOODp
ivyX3OiYbV8FTQtIEHXYOQ86YszhVaWsfj/Gnp85cEDWns6ZPGiTJLWRr/hC0d3r
83kE7iOTKgi0GdBgdWp2xYQznR1JYM4f5owEM+mqiwnfgAUocgwzxIfdYvRxg7BA
znPx8S1aJHCVtJdOv18a9IhtltrMHaZl7UU2bhLgTIRc+V3aF1zNYT8ky8LYZMko
vzC73GLHQShVtn9u5mFm4hEWqB/dxe0QR0PhJRCTUfz3mpV6EVnDjGZtrEyjQgAD
YRXCe/JJjBqT/B0eRg5VdfUPwNvaStq94l5t1aj3ZnuxeJRD7RutZlji8xQiV/P3
eFZ/8zmwVcbY8ESor57S2Zf11fyU3Vyq11cUtuRb81hgMd0y/gOecfqgrIC813g8
am/owYw29YkcygMGq1bIwQM/4B3VlxAHh1iJ35H2e3HCcTur5d0smUaQZbj8/3U2
kEm2P8InOlIGyp2Kya2lIt7CwTR+2QGsMM17PRKsmVgOIHG4pZMbciDiCCrqqDrE
QQDu9C5dBgOKU7zSeYL5iDBoL1kfPyQ2B07Q37kxVnVHlaPEPipxNVpTX6sTpXwh
BIRyc6hFPlNu+mAfJcgCSo2z4ZeDsBUaIownJKqDueIehN9Pu8dhVD+SCyD71D3J
bi3jDZ4lUZ3i/3XFVT4H6huE5oK6yqF8mbNB96z0b/HVExV0F9D8+X1iYZ58bLkX
5d7ATS+1O1vUBVBcE4jPqRZzBpEnPG3kOY5q5uzMucA3u/XPscEs5xU/ThSswqCO
+J6+Tfv5IrfTUcrLmztsJ9TFDiirCDHFKofz6/YOp4PcD2/uIwZzkdm0FGR0bhIj
CIEXAPeiIYIcp3X26YkChkvXbxlOgFiT1javDVO9dWRU1ywbXeu2Ezr/6+s31EsK
h0bw4Tb+VI9vUCNFDFaqDOEOvp3PGucfbIq8mQLHn43ZgsJFG6A5RJNVyBEvgy1o
xSpDoo5wGP+trEUaYTDcXakI3LwjhG/hDVOQ/zIYllviIaDlRach9/6WPWxxoZOQ
qpuYYopwihFWBjUV+Rbxq3VpdBFQ++VPc4ShTowBP72XclVMdl3Sa4+OkR0XXc+S
LgiCpeIiDOQpnaxTn1BfGqoU5NHmgc0K4R2xefKoKfnQc8D9oGWgQgpA+La7BfsP
f8yH2xgiOQiqyB+8wuI8+updsHa2uwPDazph49eRiDL8FPoOqDFW6SYI6Nj9DRFg
SM111riMNHCc44++lABY5SVF0eL5WiL7dTtn1W5DRSpVaTOnXsbnPskWPGCocjIz
it5rZJ0KHX4uMKPHo2KmJlUpXTlbo4NZDxp9bY1KhLyZ4F/SXmvfXIMQ7pKqmn7K
ptxnKdRJnBKItKGqPJjqyFoxe6bf4p92A7qOfOYdzbrMpVbKIfySFsejbBlPNGqQ
4RBj3hcam7pFY/3vsd/kagr5uR+PaSnoNznVLqqdUcBUrI0XiXErPgWjyA3XA8hR
y1360jvKwWMGNdfR7bu1u2TLL7ummKX3hNVlLeJ/Rdop91MrHDJ635pRvChtuIsD
w4e6J3DGhSNpkLCqZF5eQ8g84arrYrOlu0QGXKgj9nwsZ1N1Wh5RIb9O5QygCvVJ
fpUe74m9swbcf3P9hcXa0T933ZkZP9uTBIslLBKL/h75kOC6oOMAo51MPVQYYxYo
KGMqLCqvSrNQMO7n9bMa8X2Ax4RrK8/uGlGD4iRx3+94emREiNr+MVZcBoCgWjFg
44pLI+qxn/MsDTOm8u+nv0V52xoToSso7p8/3cNrFzJBaNS1sFATMWI3HFx0qBeG
czEqUxTKjL511AvrqJLjEN+zaXBmcrLVCCAERCQviiuvgfx0GId9Ewli47YyiurU
dO5a6zf/uXIcT4fqesVOs/9bK68/SK2GG1pnlbjPdWAEYe1MZ/F++lIkG7c9vR4G
X9+bjEJJJfr23XiDsSaCCZuptRv+L+heOIV/v5lRHJifZgB09rqhM5B4cL4zytjL
Nwi9uTEFllZk1z/8+2JjOK8rz6GIuWfWu5yDj/gru9YHmuoHNuMGqXz8BvW+CjNo
6SJXAJU/4phe/2aSEI6aZgp4BHZKgeZLmne0zQ/tOBgAbiVUeglE0ztVKTTwMVfu
PiqcNc6fmxWn+I++fQIjoW75sqPrDrtV+PMbxpcGekDN5jX77Ta3hmrsqJa2QKGU
KhOrivvqOF2ijrx4QVy8N2gH32ZBy7fEys387Ymg8Vd3By/gSRFlWLyx0advaEfT
QC5Mu7Vvn0KQENVoBuhukmh8d3C50Wdm6dGlM/ozfPew9vC9aOS2VmJxR/8hyXD9
4bEiu8js6kxABQq/lUVys5VqEDYBXNwgH+xnZI8pM/1Kcfr4rs8vRPz6ZR826TF5
P8SLNao9NKVY4MBYV1NL1JlIVEj32vaSIL+qViOUJLGJLweNrlsHOc4gfR9isyo2
3KIQTfYfClYu19IXu0U1V76M6CKKdTYOHOYR5oeHJmpXREoQxh/0NpwEYeEq3g5v
np4V4xiE2XKpyJPIu3n+8ubpadaoM4GCwB37QQX3icO1Z0Atltivt2NXwiUI+A5E
xZ/ZnnsXohP6CRSBDUGq4B6TvSy96y25G9qFNVe+1e2EtGlopFKgi/9X0YAwKTE3
ldTGxKWtUu20W1PN/49/WD0tr+c9/eEVUdYssZSWsrNyu7uUYpYYubGjTsts2CRO
K8USpzGWui3oAEzyt9LoE9rqvDCoVOoLUt4PI8KSf0Oi8vWoMYDj5uiyrZeh+edI
LjZwEm3yTMN1wPsqPwcnBy+j/4qNAuYrfvBPBnP+oMV6pOnRiIrLj5/WMLCXLUhk
5DLZKnFcCPPMwExfGhwmG473QQO9YRZenVeJWhzDh/meylpGqVABAvFACcEWuloA
Jqqhbr3lb3hFQ2xgqqfKLkcsorEl3UMJAnwl3vOk/QzsEwlFH7sC0qmICD7oLeVH
bOUvbx4T6ygG+hKEQHyvIHHnt6TwE1/T/s7TQ24HLjNccTDVrCKhF4BbKzkNbHgF
QLV9rdx8ayI8yxJbYZLUDZ/6uDb2XEESto6yOm9H19OGNhbbzB3cLrbLg4ZsdkN4
HxlEN+CAmXQmuG71UA2GnVlIRxXbAXALcSvPsCoAZecNNvKAdo/PxhdKubr+3LOf
McIG8xd72J+kCp1TPYSlriD+xFp60WXXz/13KjQE3uBM27PEU01YN+V2o92cBlqn
z7ksdyv9BEkiloIxG2OCer7htTz6E7HCuLPKDPXfqJg70DCk/nt/pqZnmGBf8rVa
p3xMd47t2TIdThHSXt3UcMcxxEHwDkhno4ow2POV2FXTSWaZd2XFqih8zZ1xgOnq
AiUXvUiBi26wIil2y7XlB7e321sUgN5PWcUNVyN1g3/+VvTJwXmu9q6G/lf4Mvp6
157J429Q1PMavzHku6hXcBzFV3H5hBi9vB08QGwEUtGJp87FnXRiELMOvo2E/11F
ttgc90P7zaFnlXJ5wmO7HgHGWqQ00VSSH47tA74H7rI40IOkQ7csw/TP5WaA/lsP
J6gUFkDtpQQP93X6Jdkv6Y3dEcnsSdMQ1Wmgfb8DOXF+YG2sFBuCAYzkTU1wHE2P
W31M/2d5SXOa4jyGST51GV+sy4aANQcXCn30FlxEXTcZJVhFl2HiwJ7MnB4fjULO
kD385PLmKx9jVVbw1P/2fgGQcGI93fj60RELBL3blcDLJsFk68jPU2hYRxI0UOax
mi/hjSNlqFQlSyrWOy8Bw+xYqaJn4k5JAzeYCTnLIZIe6OwpfFI+KcFu2WfZTdat
49EfIoCBwziEhJTwkfkJrcGNJCSxFRgJzoGaU7fyH27Oaz1UfOsqp6TFgv8quVSx
f4sOlru5P4TvWKaJWlFcoX4Hy5mvu9ROjocTGirFPSApbA/fGkcQ0+H1bsNY7QCd
f1LZ5qU4U94Z8p7MqdIkeG5FSlcLmbLHO82vVBLm/2Wgq9Ve4UPB8C/ZZiBGfgYl
miuSCjWgP0RTOoplk9MnZBDIHAsrgIF0ZoDehGl00ypCumXxFzGtjHm6FS6kx7yD
j21Vp/yhAsEX8jD38hOHnzoApd0xgtHfdidf87oiXDadeZYEuKhpSulgnscJK4Sl
k3oTmZZ7g59cJw/e9DzFWuiF7rljYS/NzzjoBovslMpmj5qymGiiKfo1p+Wb1Bx0
1WzpwZ4GCrMqNbSUZFg8x9c+T8R1JnBgQoLCm22BMEyXnT1g45/JFZFMkYEmwKmq
7s4wWtRwg0NG99S7MJhz3MAU6p6WUPe2tdO3VApqkeQzyAvuAzcEHpLILoZzLz1L
OH98UEwDB1SnxE8N9E/NqAdhoNW8RlgcL3GNGLAI9ur54785ro4mVkiXT9WXfgzw
lnpUqyFOZFktjJNpMxkDqDDQdJkgzgRPFCdhk891yM/jyaBqJ+4x/QcsWFSAzPJM
0bO9yAOa6k1UeiIcq5kCfoHE9mbnQwser8jZllZ0MRGex6a4qZfV3xoORxCXlIIJ
kFWdT9PZHVG+77N7PYv7c/Ht0T/3iYw0srhyI294LUCLY1kdnXKDZFVjeMPHAVPc
jW31GQLAe7jx3Fl2DrWvHo+EY4xJ6w6gbYfJFBC3PT9laOXa/MekBC8/ukEa8Q0m
s96h7X6h3v9xEp84UhlPw9S44YngnJ4NhVHEwt81crhXIWZEyZQH1dQWQXesZX26
KzSg4O1hY3POM5trivlgtk9eJqT2jfoJoPiaK5aTxJSH0xLgBBns2bpWAjXaDIb4
fX+YI5tSbX4MCdUkDdJs+urDCv4dM7QPYfqQ0XqNAw/cld0uVkkD+COiz5FhSsHw
aJnbAQitkLIlJAtUraGtclgsgfT5+/ue/7HR3QJE6RwgYcPI4q1FE+UBqm9tOjlB
fBchDDQkUe0tUBSbT5uld1gcv2qjf9arG2TDDTbgzk/IwcEL/137QkFyqNdqT3Fx
WQ3yhoH4T6chBicLvQDox7xp96xWKj61hESM0USLLAcKMMXYqkhF7/NG4fpTF/FN
H+/cW0J9aqFIFwVgKYA39Rx5p5NVayD/S2eL0h7qYCLs7VgFTQbM9qsxZTw9Ovdp
vnINcQAvkIsSV8w5mPjTRH7ua3bizxdBdnQQktTuGdoMeBCmupd6EnjUoGJArSX+
D7IDwoj7Qv32FZpBwMCNo2PsE/BCDKjdhHetYbZAN3fzvi1Fqa28nlLio4ITTvd4
L2Nv7fi1X/4CSh4VAcYGvqZacKmf28aSbGj/H+yBkD4o0aG6KgPpN+RXEsCuk6SQ
hpXCm7PFUKGgQeCbs5QuhFgV23fDagHjk6J5FkL4qS/M86MASrg5uGm/kvsMuiMF
vSoGB+fF0A712u2gaVo49xcOiilDc/B8guD8hlclW/JGrtzOLpyuieSq5jprViRA
WpaOMmjfrBp2MDGh3eEjkvIt2csjhEp99DK57tlkc8YMEyi6r19sUnG96lTCBi3/
8t9L76bcxRu6rTfcBg/3vY/qYrO4Nl+u6uKJpIGLnfz7rKTbzDXrgQ5NNDsfHchR
7xJyaQhPougzaFNrxmk7ENlbEe+v/+0+Kxi5WyfVWm/hRupu7Jl1YRroFbIfOJse
wvDofZIcwoDAPdh9kto6/a8IvNuzexAuKgrMCd35BRKOLP/4Vl/R+VNyu6w0eWn6
KZvPIjrSpgG065xgiIRk8FeajgUEAxqJ3P5vARGTsUjUKPkYOBiCEt4061EqTaUF
YnyCabLNxNU3CwX4BZMCD5YcHDR/eyJyCapCBq6hqe5QxC7elkZKYll65GwUy8ib
E6p7XoS+z/WFn0VQpJ1/nVihVxFYFS+RVuRL1044Ut3HwMqyFXgKAY9a4hLUAONo
lENxQgjZ6tC+rPr1ahGIizp84oA6ZOR31YrUpPyTBoD6a0zng/X0bow/hux3NSsm
4R8CeCwcyjzoKNlLmlXoraotQABm/PErroSqlVKJfA8CdmS+TKnyxtO0uc8w8cAo
Eprj6X6pcuAJx4qJmNhdMoQ5Hk/i3BXpOc/7lRtyu8FN2nYglwSev7q3MyLf30bK
xZDSPhb4W6yxsy1bB04jL8ceF7kX6i6kpfRToJJKdac/EG8RHmJiHk2ua20jdonu
0XpYvIT2Dhp2X0RNpt1p0dcBSakV5sgsgSam8DhLDGpxcgl7QSXFshc1SZawq8AD
17CNbtXdODVhXvpm5rvTGOSOf2Yk1TgeN8F9Wxr3tQaunYC/BveBti4lH9X7wQN6
pKJzIAxPHVsLA5PtxmEqXVqQp6PylqYanH7o2fC7tGvyF8hNQ+uOBoU1BRDkV0t4
hO5gt+LEMOhID3tVWm4H+WMIVY+rt0dq15OcUJ1vNl9C5u4SbXqNCu2F5r4G1ybZ
JR1EoSL46E73oJBpgBkaZ/BFfDn29lFmYDv3+DC1VWdWjBRg50jI4vxMbxXYE0mp
5D8Z+mCUjrRxiij/NgmFkrWtWEP2RDNlxDZp8tN2MiYiLtUDkGR6Vf/xYBCKo5kQ
KF8xwcYecoSH8CPFQFlbRlPnQG7M0j3ZTtgxbILrddQYYS/iixRg/Z1hwe+PJC+F
a6q7zmiovKbVs1Z2jdB9c4BePkDe3cwyHmwy689ytWVOnYduUHGmT4uwM11PQ3Eq
kxcsATZXMtf1cP6lyHIkt8pyichtI0O7NoWD32R0GIFjg8oRJHnosXOGzvNyvc+U
2j3OG9OT5GCfdidml61sb9lhBqLrmZIW0JkXkcDlS3ICNGXsTeHI5KCwRyM17WEE
vBFjM4emssoz6v+Oyy+FxcTZuReEqaJAoCl6wAJTJ3x6HxWXL8DJ3t6BBElmMwRi
q9SzbxA4Eefah+OYsr7sRudWAiCOUV/tT08HCUByGhajExyd/sTkThj2JT1WElHR
uSQDog2cJ1he6BvhHB3SilTOWXDTXRXnduwCKvKwcQ3UtOsppNWOlSe3Jv40Bnh3
fcxqKWePqd77XmKTUiI36SHKgnwfbwyVUWVhi7cesX8Eg7GyGGZSYi63LBjko1O0
UnqJNP9KE/k0HOC7ULzyKtcbx3pEiOxfOjxNYm58o/o6rbVuOSvdLApIdj8VNTk7
PloI8/GGC9WMAnv6ph5UDBDP4WduDmLIu1IykzLE1VuZ6jReULZvbyX2/6PvbSBj
tks7vMPe89plCbXVKO8OsCooWwHxHW0Wh+vzeOoyFQKobWn0UHbNVmg10LD5Rfxn
R5UKFufkjqn53uweifUUcZR4m+Ha0OAO3j9hB2ABauM9vTvm22DxVVBAfeuuKyJZ
GcXuUsL9YruJSNXPXojgNUIdyJTPEyqTXpvoa0Gm/pDk3fXkRdQdh29tXL2A27Pn
XSVdpoK/b7vr8EQ1tvHMdmoVxF4whHQov0ch80IX2AEHtyQCtJh1jjK3BLzLkhKa
uw++qszHA7nv7LOAyI5TIDojO7IE67dACx95aK6EwMkUX/vV6dMURb02jQtzGnj9
WZSKdy7nWl3IWo9raOSicqV2nflsxZysvNBbpbg3PpykDOPwUU8cpreFOcwCwam9
1P8ayKJ/2Y22xcxF7zgsLNRbHs1jXDeDBFV3milwMhGCATVv8TffgN7JLMjKOpCO
7dOJQKrNer/tPYwcwWSGYOqszJwgMIdTXv3Lj7G75YC47hZyCYNlgumNG+4+5raZ
+Ba/IcfMzbJbulGfA4iAMHsMRjFCpHXISujUN9AkblInRd+ky9fbakxDar+fxITr
pWxqbb9AUMr+gbzBryCxl0BvOO6zRdVMqGgUL7RTMjZW9aPGz7CN29IX67ciU9rr
siBboVPVHE0mhPo4VvSlGB517K6S0sgo+5+6+rInepDMFd36KRDBnekdF4Ikzsic
UC89RMC0EUL1zYkuZIqqYDucr/Egk3UmHG9av9i64HgUfbZIhmu63wL5L+H+OtLk
wC1Qm9KBg9eEHLimGBxY5u2Ps74laNL5LZ718SJGHO99Nhr1vkkY9ccWbbYdbR8a
YFIbgPLzte+Oczwz9p28jYpXk6MwBSfYEKTls08Go029YRF63HkXAjFz+ENX1Fg9
0Dp2W5ajDCl6GQKGswQ9HTNmbXa6mKP0XTeTeqLjWeNxImQGJwyXDxy2fI4lDKqT
kool/MKut3Hrvlu4vjwVmFHr3K9POKfQ6LUeZBoeUraDlhuBqgDHyiUpfm/fmLVh
5XkyQbB55556yLsmo5NMu41zlpCaW/nsROF5FjPO/d2NUuIwED2xJh+pM41UyYnr
E2XRUf1ZXFHe9wbL85PYbEVFDjcnObOgSnB4P+PVUixIxHTdNeoGd1jOSydBleVW
fsM/yF9KpNfXuCpzeA5IhlFPAkgFN4yFVQL760HfJk7OfmmMZpK3UleL5p+7gtSF
Z+/XASG3+nb+3WdLvLBfepSFjaukLVnTob/gNXu2WQwsF40h2M1RIC/pCQAp3+xG
YQi+7IJlkIIYDWeIfKC2CfOHHi4RvsD2uGX4lYcJlU13uEJmqd3YiogJ7jvTExeX
dqpsyRTOILo0p2DODcZ/fGzUBv38HTe2Yt+ZGhfXBMkcyVhEZkOgrawneGfyIXQo
xIfW4sEAxu9A61iGs7bDokXQyuTHdRwLJ2GUpxyNUBtxr1VBcVp6kNcsX2XU/QgJ
oKsRDJKNZDCcjwcTwMp5rUq9qZ6RJdP0UP0lhU+DZQ6cAxXTB/WvnGgVjAi27xDP
KPLiV/Ycxh3gl9ZYkoPFNqBlWlcj7aa2OZLDQU7vyGFB4jNlFiNVJzJj3AN6fcAk
PC1flyxOmW8KNkJ6ihPYREsLSFiI3KiWsxE20eUx+moA6jCnzHqjBJ4Ey0mZ28Kv
AkitK3IPRV8nA9+OLCDL3enlKWbuIrDsDTmaJTxl6iMrKJZmHTDhWTmTo2aIOj1e
wPujDah35d6+7I5fUBH2BPNP93hhClP4B597Sxo+1+s/fZ6IjK3UxqHthYw434DF
bfflhTGDcBneWYhyi9PORAfQm69trE8ufTIa245Ql36Kr/AftOgHeRBXarIrBu7V
s4jY7j94+iD+CDGri47LDdSJj2c4haCPuvX1Z2QHHN+Yz1sQ9lKnS12gI3J1bTo1
ATbKl0Rj+nOwX9hahBuAT8QOd+PrGKecpIM/+YVDWV/OiVKc4JKh8hNREA4ixBZ3
Lb3V5dSfm/pmimjVsJIM8vpqjcUl9vaYDPSgB8cUCRArSbOojNeBcTsRydLrtoM8
k2S8aK3ofkpnV8eQyWjtjY2wWNatDGuPDsj97m0m08/oKjnJin4n1PImVSvaiMlq
N0Ftq7PRhykMxSO1OLyi6JEuE3Aq+L5lFyUqxH2mxGeV5QXw+nxQ4VN2hqhY6OvP
tgie+vmdOobGy24EgRweLE1PK18TFNXGbevChPAUW+yKF5w09aQMyocGs6VgSL2s
xeVtSzx4z8OCC8qL48ajGDnwIPTAMMI7tkJvgqhNwwGyo/ZZYuPMOuU3p3qpvmYd
BjOJKONvE+VbOscyGQKDtN9dlXdVk5/Fz16Yl/iax+hdzzOybLk54F8W37ip6rHP
IExb4p1JFQ1yZ4+9KcCBe1Xc0BoG0E2s55xzGWCWdPrfjuyBeoT5Ly0XStpPsyis
YyWCxtbsrlTtXA7IRiGGpGm9X8Emy6Sx8i8h2lcuqvycihzWbAa4yE7ZcFmd4BxB
BUOsUfJnPbk67Ns9V5BnSIIETJkQLmQRWMMITQpgVqD5kzGpm5jFd6EcqSN1e7lq
rHfxr63yrifKCobWvQD4MVLGRvp1q85jFGJu7diH6FjRPU+CC+l3CQwoSVqBCZ6k
ruWrQyXQskO0D+LPHktnDx+MjllmslXqgUsWs//RDhYiIsugDXdDyVkKKUktrjFA
USdzZXfP0ugUUxbWKWTwF55CgVcYJRqzzGuXkLTJ8pVKqKCK5ZyQSui+QiDcUL4Q
k/OhElV9zMcUXIhRG7x6ziqzWUGcTEF26C5DzqjOYY6AqXwWoQ/V4yJjiVfBiNhX
HzgPO9s2VUPirWDAq9SVRTlWMenmg0pALHrjGveb78vypnPkdpCJCd4t+ssD7Jl+
aEB3MwGqICgHtALGDwZYRfyr1YYX0qTk72+b9z2y/zdnz06UvlXBLn5fn3GPpoSp
dbNEHCBDE19m7k4a2Sf/I4wl4DMhN9+gHEoptC7RvNiC6t2w7otHzmtDhXreusjr
OZgtkbJ+ZbKSVfDCSMEUn2MsbFpwxY3nNPyAOHahDVb8qhUiDKOP26k0LHSgPUsX
/g6BDl2hFZ/s6z7/ztX9GyYqhf7f0LIUFfjTXhAjBgTF5a4/3hhbHmtQw38fU6OB
3iqIBk7AeDGi3e55xYhqXoZT09kCbV8+LT+JwsMmMOs6Rj4rYwgmIoABNI2Dswju
1yAWwZlPMDkwLRfx2vbKm9EIn6G0ZJ6L+T74PdRDscbEYO2H+fyyodsF9/P7Wtu8
eJbClgQuF+l8HKZB1UvSD0g/0ooQAouoInCRnMvwmgUlhKJK/eKDJO4Q6mYRJBWb
/RahPlNs6P4fO8PP1DQ2LKl2L7Sb20OI899XhUOTWSvlrdBXlpnyRFhAAH+rYDv5
tqn4xicGxtM6dXdMP0X0JwveU2qlWt7bJjSOZL86McXbDWJDhbWVHWgX7xLPAVGw
lv/LY/mo//bux0wY/S4X0mCZMpOc/k+risP4vhaGqibQOcQ7zhi1tO4ivUHV4ytW
VZaYr5viX69pxtN6CxsKOVYU4l3Ya3xGxYvlrHUp/TY5Rx5d8YiNA9JeUiOOfkz1
3OKkDoKdOhzoLVvoeMiuTjAG1o9ADyxy18maqPPWDf8pbOvmdwBYvurYJMAqWj31
so+f/TDIzg3qQEgk4I7dvt7zDi8aQl3HxiXL52g4TOow7DTTzvf61pkMaiOofICp
jmapM9EKrwsLEne2N0cZQXTiv05T8/FCRviKIA1ZxocmGOvKPr8EH3gDKHmw+582
qNW48uJynAZks+21T49kFORfFvg6WiYciT8bMkxwq9jf+gFNzoZrEnjmBBbndFM/
rX1fRQYt4vEzk4XG7lJbl2JvHlOU9e1wxLw1kjnGw0/qhDTKna4ixDhRdeIKPcI0
tADu+S6qQ102vuN54ANgWfrZiIsZnSv/jK8UxHmvoyIbD9elm2F3K1axI65QWWVm
VVlKR704Ya8xRNuurGM/KlnfTW7KVeDmqpuYzd9f5M3oEtll6pgTikFCG91WxyKt
FkAAkBwQNOjRwifOOpmIZk5ujKDTkCfQn6VBx/JjIZAbwpIOODfWeo6IniOKI6Eo
ywTGDQUxx8t18pPz856djdv2y+qmvq9t+lwwojEv3eVaQIZnTlqBQZIwC0FbyYqD
JaTSg/pV9qhq5jyXVE98Lk1IlvkPUk4Tnidc/ADcF8jPrtUILG0a0oiXlpb3cdme
Vp0MNFbwbWWJoKtVAVDozq5ywsbqKUAH7XibmjRmR6bSyga4/1SEtqBhTrye0I7N
UgUcqaMzNijPkTCj9RfJ04K0i80lZy7TShgd+ry2o+X0/0Fxx4by7WUb8kn6tWTD
HsombcUKetWFswcSBhT2ar8ICAUx7XzWDlWx8iUoFGOI7gig6h5lNw45nHn1ncGG
HNFJHSGr6+yRPyEZa1abMY89IwroIvdakdhmgdkDoE/awzpmGWFO52J8yNq4CNau
0E0e0XsBoQKBwCgC9ZwUVclnm5JQV8snjD8gO/4PORNxU6stLMP5JCgoMAQR8+m+
Vs1uenBjlG0JyAqmn79AaOJn+b3WlYfglMI6uwq+FXyqkIuzBNZlXAADHTMd5xBD
xsQF6PGlfQSPom/DvWN9n4FQX0QZK1iJZKgcQd+F34GJ/DZSAoP14LLhjs4kSGT2
XjYdw+eZODqGAhclhMO/2L+fyZG1jG/mzpTg8t/GFGIM/8lVKUYOHD0VIHweLSHP
XK6JLu9gW8CWhh/B02h50HVQWQ1uGucoSshyoX8oO13jYNYI+stM9cDx0efT5k6d
+kWIsycovjnOe74+/B26tkD8dnDykIlqh/LCTVCNAQCXLWgdbb+peDKHDS0a764J
SU0kSWnyIKyz+mfEnsFBMfqikafh5KCtHC7TPxujTXm8TPcxM9L0G+zJuM9AypY+
8ZxNJlaoDVNbgCgGsl7CiZKYtMU6lAFXg6k6JebneY9wEDwpsgEHbHCXqv1lK4jM
i/6eeAoJNN1Rb1dBGxNUVg2A8tA6Lium3SYzNMZuNxusFrpsWqxnRRIV2XcCsNE8
czTfn/kXw2iZlFamlNBT5DwsdYMgAfDPhZedjaosQoxflaDqHyfwcDPcZWHD9+ke
GwUm+0HCuiFvKH9dYMfOa6OoIK/TZ+I9qDLwPm8eFnG8ufKQg8+i/GObnkA85Mg8
JTf5zbSm/n+qrk8SgfQ0fILU1P33sOdktsDtSbFWxqagm6OCIY8rAJ0p0O4S2M9b
LL2MLPxtaEGFOjuytDvzcs/EOuulo6q9hx5oV7ybAUhP/C5IhbyJmI112bQa2Hp4
KQmzIDGl7PzqoSGyr6JmOUP3d3OgBxfs4LSPePsyLH2EFwf3peBy463Ae42VJy07
dDdDS7t3IsNCLMkX6JPz6Z+g6FguIYvGqzROQ+XSiddGTazdQ4CDxTAHwLrRX2Or
y2Us0E+5PewEMsVb0/KvYZ8Lu0Q+0EOz+mGJ/OKEoxE9ejILaS7mZ2EcVBeFtkuv
OVQgorX7qDkZDo127tPClpSIVi4e0ALilpoHbkE0pif6Ym2z/zk1fjAVEdHEfHT8
HeSbXKICYuUQXehOszXdNUmCDJA2YOIpLLTZGbLAU6aCtJFZ85tycG6yVhoWx38z
0pC50JqELQa4JiHTv7wR7EhJ2duc5g4tNrQWwNvN+mvZc1Vd2vSjc2sOY1h5Awst
Hr93rQhXMIi3hbHyeWcjwQVRrzypw6EoKxltzPHdgZvWqDoIQZiBm23hUaqmuYgy
Lfkht1fw2OTPakQVYiZmF7JPwUj/gZ1Sena5zwwxTtVhk7l31I3r3owrzB3OQAQS
nusgLCnG21rtDx805HQrncZ5Z4qhHx5+Cb2r+j45oBRZ9MmfWwJJeuD4qGJl37i3
2luobNj4Cjh3vK1UVdEdkT1UuhjQRFtBQvGS/7asQSBkrhIdTHcTnxdUNuSVrs3J
mUJzcgQIsLsxwPnqSGnDF8FLVWKx4wx7vYc1kGKoSl6MwtuL9jjdLN0u6D8GvbVr
nCjcbvVqNavjR2XC1cNr4kVJqHGKS3Z5NDFgZ47HK301nk+5YwwWO2xg4qZwNpZe
49+AFiCdzAnM2HGaSceqltOeR7mZg4dfIkIJE07Wzi3VSJa3+tvNFB71x1Lm7BlO
oG2+yc2JrQYDqyIblHuJBo580bac/z3BPtprzGuHm12vWqXUhYNXEafiMn4q4e6R
gAFYhr6gdzCEIH/ERCJIpF9NukeKQsA+977X7OqIM4jds8O+rk/4unMOiQx5o+Z1
+3au0RC3k2SZV2Iaswj0Qzbqkhw6sPGBVObbeuDepcmwjdA6UXgt/OcXDHbda8dK
7MEtG9wE5i8eQfUuUKERSXYlqoy9VoCMRjKkZLWvWGQwNZlHjvhAJnFYd69222Q6
WVD4Q96W1Npdj0IUaTsgPHNXqk103SV8kjbKwpkg3I18iA9U0A9Nc5f3LTW8c9sR
G9at7RSg/FSqdsDP2UwHmDyu3jhFNV9COFVdgB1TeOBuo8P2EulC4BNifrzIcjHG
lIq1ja8cnWETOqPdFqHRia/gBFfaILymQZ1b4piWkovH0c5pL8UceS6nVlaiO8Cv
TZEnVWbFnKPtn53ltaG2eo8RXEDebHnfyBkfmxkwqbr9ObQLghtjC1J6deADl0ES
yA7qMn1mbQuGBt97bR7I05DaES/fLWmlpgGN4+IzSivwHF/M327Q9s3TZDYEXjwu
8LTGkuWmYp6+iG7+gbsTkihwTne1HRBKGF1MaiknvSfsehlENUPQKo9V4DclZhN+
KfwgP688ZNuC133D7IVx+tgB+uUZN72+QvxalSC45bdXvVlbepCJaneNPI3y/wt8
u84244tr6LcHVtkIN9VgARECLOLpGnyVaoJVa5bswsf6QaOuimfX+LBUJO/hNMb4
fqGdTNX/oSJT97xBQtYo7GLj4axcDQCD+XePGHct1EqGudywxnNAAP1t+xN5Dzmh
jVzgOTphcZYcnv4Jwq1a4/pnPdXpupwKnvG+V5FBN+x4yNaH4nRxevWwXIBUIAF+
2ojElbqxiKM07W0gG/2hB6G9jyNHOZ6UFj5rSHqVi9nHWM8xZvZDnjyUPhTWwWt/
kpQ5sIu/Zka3uo6RAe3KEo2k6t3s9wj2rb/THc2Dr3MHyuzRjcVYWhSJtBAM2qF3
hgFW0+Q1BvNyOiY2VBE0eArgvhpE86SqvlYiQ9yrcnhEDls2V75OphN9+0ADOc5g
Jss3P8eH/MBcJSYpzDzQTLwAhfzg2EWcm6784jJRM9azdE3anuHmE3WftLW0yr0v
xw3tEt7DlRLV/QwqI09csrq9RDvTxp70oSu5CKpBbC6W7L6G0sqkS7P0C2Q87cmU
N09iW60agDR0+6MY+NamC+Bc4h8EAw1LVOFONXb81nGg780P7r03n/92TPrY2hYB
ZYEphHLL2KVRKSCxHnDHiDoX3lzHhNPCMCYuKZw3ha7nr7hZfY/L0zDzMikprEdd
95UAUU9i+S92GOB8/XsbusENhWBd0BbkAH6TVjaKf5aRhxPXSPOeAdNm/gYihJJE
BpOqjTEqB67xbzVuoH0rgS8AhnWDkesVpMBEO50zCkKJLWKxq4OndkzvgmB5HEoU
smbSWhyMmVZmBTNYXnTPaRc2wpP958rD9BpO2mB0GIOLyKWfwOJnPIgFNYjXeoBC
sPXqFPPHrp+4jWMJZGWl3fe/YRY+CehBxJmhRb0WwV7r9CJWG40oS6VfRAOvlXcK
IukBuyV1RvaWNyelTpW+ZqkUrllZb8VlM/qj47E74wPdLKfEs0QtTWKv2eOoxAwd
8AfsJan8Z+eeQ6046SQEYZaX9p0ztCvyRKEjqmajqjP52qHdz9rqoa0GcYZWL9u7
B2AF+IgMTk7FziDeQUYQ80ZmkNqRlmr0Z1wBHokU4cJmmTyog47OSWyEXF4D7YB8
YPbZbS/RO4HV4tGlAIdXy1N2cWM8Qos8myXpe9wuY9SGpyEtpyuFGrVciy5dnzK4
7TiuidUl0wYXFFasZ9cM0NPEegqKngUbnJaIm4J+OOkD7+V4i29On8Z/Sp3Dxl4r
fSVWE7dbn/Rr1McpEaldofKo/Gd0mNAFisO1gQ5B7s+1q/EQhpbTuBYGOK9Z6YtZ
ybuW/ul3/o17Njrvz2ii485rzb/2ianvDG3VeLFW4gwcSCuxbb9ElW8c+g0ZIiA1
Z1wD8nKhCN73La61DS/rvyj3Oj77ZarQvB+zt2h+Q2KDQ8eKE33qQA1YOd1XRd0V
gIyiwV0SukYqMVsfO4c+RtcZqNKqCzh4E4J7MmXggj4uCMFkYeZ7jc+5NEuPsrhl
5l3QsV5S7JZjZLpT+RYkvuAvY2pu9JkAzHVFLTwNZCgv9PUMjRUc43RqSEdtSGgm
J1ooXP0fRNp3AisrMSEXjzmEOQ+wvTTVcmkrLRtdM6dfnS276rJySrSVo5v0mcmh
igfLxVTYczs8gqvhJ2G9rgHTcXcOs04TuxRYoOrK+PJ9+rOQtY+OqMP+y9pMhRBI
ZEPNHhpia6BjlrGfzjztIxi3SJlBnqJm1AGbv3fRwF7BfdfuSNHBPH7b8zvey7HV
8rJrRr6BN+uKKglyoxOVZxVv6/k7yJ51V15deq9AV/ySkBOUnuUXuiPb6xr526Og
VdgymI8uAuMrZCXWcI6f7hxcqCSsQkAate7AplEUFdpAX+Isu7LeCuHeUBI13Hv8
rOGzLbD1K1W8+/omLdqtk4krM9MLg8qRf/6tDqSrjKbMhtK/pkYrg/WrQ2WerI4J
hqpYT/SJ61Itb36NBdArmjRcR36hSKtxv/guKfs3MMUnbPvSm9J/k6vu3eYg1ELf
VuOS0X1+r6MVWuXL8aVBIvG2tB8DLRYKaEK54vmzN3IuVJok/6pcTIcfDAfDiWW9
rq+r+e8wbRnsPJZ3mZDgzr01LdTRpSCQ69OBqdaTSoTzBMjc9JRaRProLxY2kEJR
PNAk+6Vt+ReKq7/cdnXqnVpNAWsCbMoRSOLNTAh4XgaULgnWsGO2vrSOHPE7wlxo
ZyBCJUZp6QKrPOyDghn3VOc2M1NghJDxpz+3mZauFHee7Iq2o+3vGRmWU/oR3omJ
zKsuWCB0G1SAUjG6fx9fFGnQsvXVi8Xij//fxgWvWRdIKmFrxjAOmlFJOicQreW6
Fc0DnVPRmBkOL5S529O4yrMv41Nh1/KDG5cHZYIjhdYzfDCgA6CLReZ51QVhMj2M
84mL6fILZVugepoASafz6LoIHreTq5E0c4A1EJ80WJ6efoKDeZ3PHez/0VSy5s4j
zzrj7NJdxR3Q4s0+5iUet7VJWQqS8HHThS8iHlmY+j8/hGhXCwSHWXyAN1NhUb1X
n0VmVuTOf/5Vnr+OJJyb4D2nNRjljZYVzQyVB8AINUX9pBE2KTsIN2xXDiFM6uo4
mjPfYhT2QZ7JP2RWZ7wdXCdFLRk95Qoss324opsnLOsOQHu+y76JW/D1JiKFxOik
oFqDjbAV83tPUUOfa6vXNsiB+ZyD0a8H79r7UKmlN26td2EW/xTPgAi3+DqlqwaE
ixzE+OMVqnRBGohQL6wUFdsGlo0k2goI8DZtZ3w/CeKs5W2hfWhDQyTFIWEkYLhx
f+qBs9uJXR57vmzNhYc9RPpOgXnr1qny0cFLuJw220exEC21SA6Wj2cpraH9eBIg
xjm1XzwFbWXdS9VJBkGlSnylx9aVFLqa90ag+OlelGGf+tfFJ4TRLBEosUly8lKp
kQuoXx9GX8LjEt+QWJ0G60h+LRSqbq6T90oqJgXOh00BJFZKuOVr4rD4ET/Ui5tg
t4eeyESwXV/XfCEP73H8HSMKkn+z7DK8cHZuuD+9CzzHUgnOLUKBdf/Hs1nsUq/O
5+R2KLvBH1R35kU3TkDW2U2dMKNeT4ljjta26MeQ9BiyrofAmTGZJNGDv0Tz+xNs
k0pb+ZyORvPyM6g9kiW4rRFr1MFrOfmFopjSUL1GDfD+LiP+AbZseAhRX/wqqJDh
K/y+xT5HYf+u/m0NHQ9fqUIoNp/B91V29Lmj6ztygWytAJ1wJINQfgafU+/O2tMw
jW/H8Za4IQ5tNVy10w6N84P2lKr9wUjvbyjvyhV5HkPsMCkWR6xSNsxw5m/jCLVx
c2A9vwEuaA/OwHm0q8iqHJaYhXH9jERNAGRPP2CYB6tuHdmttiusfRLvio97Fe2L
IWHVcVg9pRFKpn14ZTRHUAhNPzsHCF4OPPB5SJZY4Zb9r6LKU6WidRoC39Uo5KFx
WrPt+oru5EZbxOaKPErpwPWParzF3sHhGAvA2yrn2GAGaU2SQQccFI06T8rTyhfg
G2jC+pv3ReKPIaQnw/xMQMMSYTutfXiybWrxzKwuRwPBBPsh4hN6MKe9BKDCLe4S
lRHlQz3JKR+0a4s1kRoR4ow9CC1owsHPayNYmf1kb/7V3Gv0dAI/Gzt3Sz3O1Ko9
M+jDg+Jrct/qQRRhLaA1zRud2keziwEVWgUxpKgOoQogkNfG4cCg//qIePEf6lny
4li9joyNGL4C82akCqtuK5MEAbXNvddsqb9AtnvsqJpry+J3HpIaB4DOEuG57rXX
5n+tq0DYFYRICqsDuhqrqu1SqZJKZ8M+ooSTVxvLnYVDeTeCOuMgu4xMXkLu6MPP
XI9IWKXt88ljIwVXQPBKumA0qhr+0qEiE4oN3SBPnFRCbFgDtTE9oslrQo80kBKn
KNpTWodssqm2GjEBF/bwP4cVbIyj3kXSBSd5Bpk/0u7xAdmrLPyQLUlr+MQpe9Il
yUcME+slTdPJ0/0/h6s7RDzPZG4s2Ay1eB212ihu+UcJlMiC2w42/uX+e9eBRrZM
Qc1OaMWE6CMotD3iC8f6bioAlskmAfyxqewZsBiSu4DD+7iH+9t8gxE9SsxZBz8h
+dvNg0vT1egClUhuQrq0seQO/FsSt53P4KMedMX/ro4zhqQ/UWTSbP9BqEUChSTC
2YmMkfnuQrAwDpDWJpvsjTrwlff0VxgykTY5AYQ5Ys49jDWCCKVOYDYuQZSbBDk+
+LFsGf5lH4bMKcnyaW0SYz6HM8fI/spRV4XZ0AReZmq7jihus05iDNZi+50XNSBI
nCk+7pH/0gJAz7vie/ICkQ/VBP9WlECu92kB0zH6rpJMxNBORJOaQOl7TK/LXBjs
hyh4A6jqjUL4jfbtLV0La5vHh5Kgn8FQrI8h/nQtrT8+s6+0hSg0AvQpuap/Iew3
npmUTEZJ7CIJroIbRA7K4P39LVwal+QTkTEAtVzcugH5BfKBuQ+2EtBVLVCdXCar
RWtfCGgHwDK2aVEH/yqCLl1mdT3Odqykv7IqdhMjs+ttzbu+uZfCcOp0PfCNEkYy
1huKZGvZHcFn6Jrch9w/87HG8r5O4xf07n82yqkkcmBAqQ8ZqZFwI+MessPj3jLV
El+8hAcV9KDz+qPkBms3h0aYrvrJ5ekpRDD7lc3J1vjv6Z7WEOoh3Pntpn/zlBIL
tumswjB99lmqyOrYQRa2x4ysKHdm9C1AqUmW1CU6vbY3VAM438KJMP0EtrXAASy6
TZ2vYjJRnFgOAM+DbOeM4DIgM7JwTadxWrpL102PdVKWunsHb295u6SseObddcU3
k8PzTPWiPktBi3qtV4MbPHuODsu+t8rYiKDqi6jDQLkW753DRhTYHNyW1JWUxmam
R41Z1QR6vxG7Jc4qvvzMadGrI4BwIQrABDkTY6DtenPVG3y8Q5hnYszYNQsBdRqI
geCBhcw4PhA4+yv+JVMrYV1Naxxbgz0egnzKb9bjL6AhZE0dy2yI9VAPvpVvdAxt
9v5DWdE2qX+/CcghGS/7A1ZtWxeseu7TIUHYF+Daxiuzdz1ZqZCoFNTnglSvafta
bC3xSvJVfoHZBta++AYBnCPHMLFUZyizexbAFBvSmsPttmsvf4fdlxhNpUWpo1Tf
HZxURWN4XplGEN4DtmrkhYAodfC1xIXsbXGVL3btJh7DZQYR3kUaZXCI+zilpiD+
HbWHWsVpW9vjGNg1ULJEqpdBcJvIJURNg7iiVsAgw47BJbwMvwDnHz3IUQ4/17ia
jfExF5Cqd8qrIjXpXXALUPoDJI4O5UR1Gw85fwvfQPbEUXGPHv+o0rukSY2ExJuA
EhF36TtX5aSy8e1wcuI9587uVNzkQjhNLgmuxa6KRdLK2YxBu2I5/Aj15Ns8RqWh
J0XJzZ+0O1FyOgzLUOOrO7zSuKAqGQ7zgK7/wy5FhQS6LKbunXniEK84u7Wb5YW+
x5lWZyigWpTc5k/yxXkpRTfYL3Y6YeGBc3hPmKa8hEs2EZH/Mj9ac3xYXj2ZX5uU
d1S843A+PHxIk3ZUiTKZpskZ68qiWiRqcMitxeuDn2EjzaK9APzyJs56FcVavlM8
/B1yBffNcAVmD5Q/0EtalD5f0yJhOlwQcWU2OONTMfai/ZiTNypAo2ILbwDaeXFq
cHSMpzhA3pSQQM+HZ1EcD0IeqJilOi7keuQsxaRe2rUvPjzjoxNhROWvxlyZQxvV
AW5k9huiBbdVMfnPiJAOMCQ5WHY5IR87ZMZuMfIXjCy/FiNOXclXDWMGWOuqDff8
fEe8NbAex87YTZpEG0+Pn6b0bEV0WMgQArc9jiqjl1MwJRHagsixCo6gEaMmwygG
uCYkagEZ82YNKEoKXlH5l1pdRzmcSaJqdUYTQodup8YKLy7rH4B8JZidy0zDUIh2
0Yv/4nFe0rgRG5TLOAIl4F4EdfEgroSrBcFZlN2ZC96g5EJMDTGAru7xFVpVbcnQ
ryItwqQdLe0I89q1BAFrGS8M7z8M3POvdvnq98s46edAeiCxiu2Qf0i/MtQhSyqw
rlNgBJWguyEIPvKwapXsH/lddoKA7clklVMg5vkNmaqu0CDgL3gSbG0GvsA9lyHl
7oqTPTnjV+yDPmpyD+BppweRafWU01OdfNCyZ6rqdpncSIsoaGS6hA2cGFP+Y/Gl
+uZhPdiKioQa6TIANVQFyWOkF/RDNe3F1SyhmhYh01+WZA8G87gQoNvlbeCFWRnh
G6xHKJdrQYfbysI4fOleUweljd56Z1cCep9DbYfKaOR1LZMtAGinfMYRKyOfWSQx
1PSOGXMarNlXjw/dlDrDem12veDI2ah3SJRLTUeG+N+DGTzHaPPudDTzeomZ7EP6
eKwYQlKlUtUKBEA716CrqX0KxfgLZU0BHQ2YZZqPbp9cJvReS/ajMP5PY/X9YbJE
Xn5fiSevS3lY0FDRUgcAbXteM/24wtYxBFwKiqJ1zep2IP3Y2GuhRI9SF3Zxx7MN
eg64qYQ+fCxoLOgw7OsDKI7QSH28qlBe2+U/us5sS+SHivbIghTjIVa9kDsdHZg8
vfDcnL63VvK3aLsoNTRSmf6hk6pjOoQ/vq4NcSYyDlZC8hJDgdzywmWymkANjtPG
6hpJQX0NArgs2Z3r6RxijikiQbyJF0qyigqSO/JAkjmywp2gmHt+/0u4z5R24bwk
F+c/BI5a1CsP8X5VdH493cN1bAVw73WN701h+Q5QhsdcWkc5+3tNHkKKBJFF3rUj
hFsgfWag4l7M6lGYeYSFVyC9v3bZ2pxGItVTm7l0IXXnD8r3mSEWVTfOWWg3XaeO
oRKZP7JEtAEV3JzJAYGic8WCfZuE+XPzCjaQ1hcVNnEoRtiUf3XefakPep89TvSo
xlRYqEzSFdIFKN3Kd0IQ4uYi67jwoN6z5TYHkHMG5/+SQifD4//txJj6uP8z/gqn
Lu3AQ9vcKGey6iXtiSd4SPvaHtdD7bgDv1r7yIfQvlPlhsoFJWcn7bj4eACShzey
RJDgQlV1+sn/upCa/6qI5lJPiwwVq1RrRPglPxbfXpRyM0iS9aevvClzMbQ94UIM
JklWujMDjac/wf4FmVo65AJ2oIPeh0HRKGlXqC55B7vY+UoQ0evD8OqHrW1CNeOh
tvL92/Fm+80iWsoYYTd84DO9E0nc01Y2LaK4LJWpC//7+6zjmxvXU21BEtMx91/Z
8oGrxTZq+tFnyRNOVwAA38NRN1et/i+6fCb5Z8HHko+RrsJ8UCsUjRzBT0CnlRrn
hCaCAMenMVv2ZLUxAetFb8RW+8yWsboDEC4sto/xzk+6k+xBIWWWEQtkOw8xkxAl
k1u+sIxKU2fOiKXlkjYmJwuueVeMdC1Vyp07NW+tPdq0t6NJW9Xip3oeWl4T1ONx
DWdtaUaAPv/Qeqag0zB8y1TVPu1g2RkmNH2nsIAXkviSt5G7Z5Rmc5GMl8+7fCDy
Zifyn1cTbmsly+8bqciRWzSNU4m2X3wDhCnpJ8y399bl3rANeLD2b3MNKP9SPpjy
HnihmJo7TlW00hZKog467sHzs48rPJ3OlcH/+WjjLoYnzEU25X6DMEzgu3knhCVy
qDZZlOP+QOOu4N6xyu/9GLM56d4I9qFEZld5+iJB8Q2Sz2tXqoxHhYrGRv1Zv2aw
fMm0fwkKm/rjnF7gJKYhs+8L+hTKrN3m/9FyRVhuNRX51YVZYaoJ9LzkBYxrPWgS
A7/CdKjxjqAZgx22Rk7RWfqYcdmrxBLpJ+bXyT3Z1xXOYBpuv1FAkobozahHygAD
hu1kTmSrJgX2Bq5xYQlD1REZ2CcEKHcJj3ksJHkfSb61cwJai+U/rLCiclX9hK6u
2rPrhluoqA8ojoZZgBXIe6CwsQOmbDFqr06jU7lIXOawpJ3wlSIR15PdYvg1SrMv
YclXL09YA6ov6yKxnMl0lj+89HddZbJ2OR1tLWIiaI5rPnhv1TKl7M2lZz8yG1lG
DOxD5VZb3S0B4SlzJhLrcgXe1Ka+M7Z+6dpZnB2CAWjGkBUM1z4b8HaLzcluzwwX
TV4U7VNOMT2FqJBKDvQ85I7mlftOOERX2vynbScnzyS7HEUuzK1xV/9AIH11/0Fg
9MmfMlB689eb1JtVLNNAH0/1Aukwi9GEcXuKQU948LP/Dimr4weyUpG4d0wr06bB
A04/M0/62i/aCb2ctisBYS8kAZi54jc7qYrA7iWLtTwyqVtCdCMNDdSXyuR9ngMW
GoM5fBmM2JJN5C+VhkEsDm+yBq3U1UGr5EnL8qkB7YmmLHf0t4H7l5Bn0vD9JKOe
g4VdGAJ9yoYN+O8FOeOEUEDfsN+SaJb/zK2IMROirMNbwQOfsyzEoG9xIIIK6US6
E8DV0xgHf8conu/Yoyp3KJGamcz2eLdUErsefKbT6gwGAuif0w+k0vHM6HXl+/PK
EoVOcdwI6vmJlVRUtXV1VB/vZ+TEN18bxvjE/2rPqtUb76XQX2RxL5JHf4HVlLj/
tPZ7nK3W+XKlm59atUQhgFbDLW2MO1bT9pL8NfIEm7qUOi56coDp0thauA2TAV0d
lmfU6BwXEvWiVPpbuRYFww791Nr8/dMT2sd4x2VRgay92uYipufJVvp+DISxnz86
rz7n4bA0TcX0FEx2VcB88DCm5zFhf8vFGPTSJ87nWuiNSwbQP01tTH7gT2C8eZnx
SX/rbA3of1RETNGVSVMdDzqqOPY99M4Iz2BqdWy3lDgFm4CqbQ9eW4HXx7aDzt6t
/ErDYJy8plxubHguEas0n4nYgHdDhaYaPmtoB+ZL9z5gnRMY9JV8AVp8juVULCJv
VJwvsz9KSYZupQjLMYpTU9fcqH/FTjBqitA9UYPFqOpStxLB0Blutqd0YpaSuv6a
8qmgEAbpaJ1etfBCJY9e+wC3YBainAsv7ilcjqWMIB6XIXUWtsii+kTbXXvvMVRK
tMKsbLGHiAUCORRbDFDZtdxtCDEDHqJCSrUDYcErepllQHLbTPUH/zrluwTFmMby
1mypjlYFpDJUB9PoHXgsM7S40Wb084AHdfzloJJsCn6ySLUznVH4I1yXsAW9569p
uUPQ7eoXaHLnDFJ5UbSDwcq+WIHv9eAK681U91alfCfve6Ng7F1MDMGx2XbaRlWi
2x9Gs9WujvexBhfMM60riygBF7+LrCm+mUghw6HAvux9zYpzEBHQgs9aScqO83/N
LGCtHRJAWLskVHoN5bGX2hOx97cl2jYwRYHDryJ+OUbizJjbbsyKpw2A5dOf3Ct9
Kp5fb1oB0rras9a25BT+zZIK0F/5Cw6uBkg82nYf0f6dgoSGTdChuaElR6AnLAfz
KDiZ7WlpEkcG39cbWwA4R8El2If4Kk+XKvGYr6MFabdxQ99esFQBmlJI2XqEmllX
CqIulQas4ZCRXY1blXlGEoq0KJQNvTSSrW/frYad2uINZ0npxiTUhK1AXFdjRI4H
WFfk9TtSW0JbpEL9FqczVw/qQboFkWqn9Et3CBWqZpVVIPrntDz0ey5uTkNzRNCE
KpsP1SmM9TO2JNG8NNKmj2EGkooGG8iu8glNKgVY6+TWr/EnWmZB43HmsJyNu7P6
6uEh5402D5NzDw39OgEiHhGJwPGDnkF+7dscXR7KcmfV8dR88yB83dwVLmxUR7WZ
UrdRnZgJidPjcRmL6NTWWYpJLkTdq2dQEsNZCQO3UFjl/1jXwoJP9oBhekdfS4bu
S2y3aM8FVSsYdFuZ/Lrl2vG7p+RaC9mP6Q7kljoARp3FZ0T1D7lsIr69d3uI5Hl2
d1nP0qqEz/ILktXKkAj5j4wdotl3NUKjhgzUVib0WxW1lVaRKiFFv54MCAGbLICv
r+ukqc42cLwudTsHv+OK31lbI6tSMJVPKLNtrfVKFMZyZwWq1ISRMJ3thWOAPbhx
oWMdhjqtrIOYKqAu95W1ay14GflNCxlCq3c9LZlYV6iqcM7/3sh7qPogAb6/DESQ
6nW5xDz8A5lZp7NDROobJyGldMfhkfgGaM/FHj6IJvqV5czE5P+uMIIsq8RTm1aE
kXHo13W0nLpQc08EipJeMN2Fw8saN5isQmAPObbHX5sePG0dbE1aaXbHgn7jvewh
YaMufzkOmYFoVnqY8neV3MaVvxQLyJ50HjdoJH4c/dNYrNyfhZU52PzuZhysIsj1
LGhbgq4f9Z6Zg7/mf/r0wyEJZsDLJ93y/vKXFZhiWDu6Iry5J7S5zCRe094/FFnc
VcbMLv9k/xzZ3jBZGULja9sURdsJUxEHDeUCU0RqHnyz1a7EfaNvkbfKSJMRx1+C
AFOHAvYLCQ0RrAhcOVuSbynH/zgZZpe9XKUu8ScmhMIflORf45PImdO6a1qpLU8k
/m/i2ByxBBar/Wf7WZJ5SBbWW8e/V0YJj9T3UMokhvR2jI2R083+mmeJQkA1He8n
EabrFe3i4U4hphex5tvQlNo6JOheWbct+Js1cfdysoS4oRDUfQPVn5FIKZK0uI/Y
Wo6dND2tBG+sElYlxPjrLePQdL29jOVx/8TwX/SBf0ZlUH230A+eOijHH+EHw59X
LDkqimcDTqAxoCAByHLpUJusChP90lzIBxzrsLGXvTb4aX5IJKAkSO3XP4INefsa
aTNKuBie/ltZSS5R5HlGR28VCbYlI8Y/GRH0ylW9sKUQQKN4QaUAMoPaPWYe1n3B
ivWjiyT+KEsCeurxfeW3wYXijepw3Ruy3yRX0IFKJcw7Ksvp+JSMWXNkpIB6HZ3p
VBqTsZ1Zl1KDiQT0jkTJMkX8EoMMfkDKqJ5RZetCXK9Z1VL6BmWKJa8C9ZbP5mjU
6IkmZvHG8NIkqG4mOR4SWXfXv3JAZEOMTV0LwxnMbc/E0+Xhe2PHuJ+dsxUuM9mN
KxdoMxZ/T83Mmwx6+wEuxN0+B6+tr0UN/coPSBJlce1iZtwYwX4DQQLggKeXCLlP
cpuqgsZc7HoMSFFvHEpAIxkQ6ibzchmLxQd5AvKyXk+BsRDmqnaGdcLqV3BHubK3
/klxR4kgQnmhw32gqot7Q7tPMkR++nKXhpjbQ9d28QK0Yz5M/HJpxG3vhFEMPBak
t9+V/h/YACf3taiqn2l6lZ9IguOIo+g0Qf3jqTQSFZtsZcXBCt5imMZTF4cduczv
I8PbdPDVtPry7rAujJZwbtPSgSs0MhKVQ5BMSHuwZewc/7vTSZKd+Nud9rEMWGFg
JXsrmqjLprOs1Ov4/c4KzkAwPP9adRro++Hfi0i6cGQfvs0QkJRBp+IxGRcHXfwt
bZURmKLp4UjiH6FEtfkn7YGwT5NzwBco8XrPk7NLbO28grIyIa/44mL894h2wvOs
e8oy2XUB43PlWzr6yBJsjEH6J64zpSUjM9N6kIsCmafW0CYitx/jtGrbcRxoBvY1
qUt+z3KlmP3PLeGICdJ5CLmRnmpDlH2vvP9CRMgcbNXngDpw/zqcE0b2KJmmzUR1
vmwjInba6UGM6d7ZXHRvaCCUm+TcAk41hp7ZErwDFCUyANFW6955f549nlJQcJLI
sqmvBWIQamGVZo/KXUdIyeKH26Ok+gZPESYEujZO/CrGpRU/GdNLcDNsBTHkGiOm
Fin3x1oP2nSlSECe0Rcb/R0ki2mVc03Lh5PWMMjB/LoDpDWKnBciXROrfTBxZoqo
HtEeMDEcZzoJR0qrMfjdK2JMPyVvKxhiEPI7pAFq7fjqRFBX4eb2EnM9WibNad3p
fi/n2wAvudXLnKvOgR6wnT1x/L5baSffzLQhdAZQ7CI9XgsM6RcTz+aai79zYZGZ
Ada84IXTu3zyESTR71rwJfwjsHXaQQxokKE43aJX3ept7K8+EmcrXANTVUY5L09z
P+Q+QaLiuX3QMp/0YJ0AnUoV+CyH5TTFHKQqlpn8XW3e3SZuCUESkAT0FYNnGnDu
R7LWgJgzHDW5DYN9ARR8apb2z8AJYjubsvs7p3nXHga1dgz9q7E6MIid+8PvOz4l
hZTLV1So9oogJpiCMmvasFvkrt7llgWSPnlFy6wvv6TRjv7Gw05U92p+yPEjcfcl
4QFd8vbgAHR4JEG50l0qjtql7+pSTwQ4yqeihfbFZL9lCl1y02y+74aEV1DOPsvu
fd/BC0WBUlixgw8wMjUJ+HOgaent69uwzkaPnK9+vo78Ym0nSrKal1ILUziW0a/d
oSxvcYIv9NFTxgppHjp4VtmcDnN4I8yBOwdVb+yu9bcyqz2V/44pb4TqCZbMB5n7
IIrJ6o1vTwkEUzH/vKu/8rgbxBM6vb7lqXbpKM8RRrS90ao/fl2WsVC56yTT6gD+
crbrsalr/CLwVmOckcbNJpjz380HCBDUA95F9XeQoeJGRAutwq7TODfzqYc41acL
E9Ew+rngCISqE94/X+iUrtFYc1gP97WNrBNTs9AH4suFiLWfw9f+gw8jDFnrksGG
ROfxksNKmIodLE8Scc2CQkEJe2Nb+R4TYskCBCwm4DPSUbilOEaOPnSrY5GLBNMp
M70ZRE8R+pbb9fujBJ+TUfGbYoprQdYJeNmVGEMJZuXVsVjisJXrg/vbvwO7ZUOx
82732iV85+4ALNQB2y2JzQpOGj4jD3uFD5FmcS2Rexs7FM3E6Vh7X2xhWzYPDWOT
OXDUyV3IQeoStrLSDgdioEFUuNZbL8xxQQw8LZHB+eBhpjL43CPVkbOk0/qR2XXC
NWP5IKV8WHXq/HZGyUHn+0r4QX02azHB92BQrb58PsC8xJawTF19Wbc6t6YJd/+q
GYivSimLqv6PQZmonDQq6F+rIHLJcEzxDwcW9ECGM/xbvDDGivxbzBtzZlKtb0Ss
qo63kqljt3zS7zOq9ft+lsw/9+ASYrRrn49tbX4ijaGvwnou/22lbe2unFNkmZm9
HVP3nEfe2jx12vLUR4Stl3mFaG4kBQfVwJaigXj8dM2opVd6Q2WXsozTpMjy5OG3
3bo3yEKoet5LuHbfX3TbcepuQe9lKr+kPQzC/eMtQBd92XQF1rrBPkxCsChQeQ6K
6PX9L1Ys+ibIoT08DY5e7/QK7A6ObOTlfQigyx7KNmk0rOJ6I0WNua49TbWYgZJG
nC8H4pdj97qCnGyzv6iQJKu/KicsLguZzfCnZ8peEwk6HSlQgrbVg264ayPiazKv
Aa8W7EQim+LBLBA88+JF6rPBPtL8yObHoaLM7j4Veraag8cDNWKXY/YanZZejIJ6
J/Te+/4oVuM0zQoGOh4e1kXF2DDXZKVoc41FB/lxhvUVfPspETKvx0gaMltvMLff
VxCtJ7tc+2MLEz3wyteJpzTqkJ9BgW/daOUr2okZtYw/M2y5YTZPA5lhWFHHGpGK
s16oW1ALVOhmcKVcO/zM+M8AxXBmT+8iRR8vHXIgbcudwuOy+vA2hx+hFMmQan54
uzHJbDxXBdP7bEAopH0umwIJPZ7IP7xAJJVx0+CU+3b+033EPKiR3CTpqekQarBz
zG4ixESLeTWbBIUh7/09CMrV3b7puiVLLqqkYgAr0QJlRJj/aPFYHn3GYpdf9rDu
2OIfZXAWbnLoMcXyUHulKp7ljXOwazSNYZqir5VJ4td10zMIYPKyvJ76PZ9XzGOo
2l6BHMCOGDVJdaE472m4vEDbBcrMpJlSagpgnzELqfNe+A2ZRkElfZKpfDKOs0I0
mQNx4uPq29KAETDqI/iNTr2wWMsMpWbCnwpKu3zJmIwIb5GZC98fEI2xhylezzSU
v5GdKG605WRfVyCnvaMLOOksjts0lBG67IRtcKlBR1jIKzVdNS7qH5frM87kYUsL
cn8IEmDIHJqa+y4rKhWrk7WD/cKs9z0383n+XwzcF/DyNa7w1MsLUJYobM7r+FD+
vRlYf7QpJRZ5eNluEtjOfOfUZXobIT5cui46EXa9qizp4DYlWiE2Z1gxzZxMLiTT
QL6Ad2iLfplWsrldc+Y1R43W/l3cszkKy0MEtBtdr7BJGP009mMDrwwUYuVRrfq5
+0hJB7ui+v6tlBmVVoObyg6wYiSHQaOmBENcqVLFzVH/iXkp/RYY1oYpv76a+TGD
c3s8cdbNWBx4cWCoRRu5rnkEbgz6OsC5uyVUAxL4ZmjhEu0AzOlTa7jeMIXSW2Uq
BoNl6NyU2GqCdYuISMt6o8VkdgTJPqGlbulfNIuFEmPG8U65QkatUV/0JY+KDzbQ
FBLbhBy1JdzCNY/CcK7aDv4gVh2rS/ZiXrGjV3INhbUMLNNswIGP8dH1VIJCero+
YBgNxZ6gfyrbnOogEqw9Ha0ckZLTkdm6ICe4h3aJ5MUwvi4hGnn04D2FPFHvdEhS
mx4Suy5Qu/shcoQaQFcFe5L/mE6CZKbJy+b+fH0xN8sGT2PXKh1JgWIVMWAdDl+q
uj+0ETCjf9XIroDEt+4JRQ/9/yXRS31gLYfZ0kI4YsRjqLCsqB3yF6LEkF/vJOEl
6uCI6JJot/srLGFkc4mzwspKfvU9UdjsO/weajcf+Vicu+rIlrbFbBj0yun4Ow11
AAWXwjyzQJu6a2/344QvIg2Z3Va1gmREU0HtaXTZ3J1KCGiqFLw5b7JIqaXgn8fg
HR/j41luApypQXHSdVcNiKRQsAuBrq1tQml9RgbXkH2dzPipeARZjfE/FpmuS8XM
Vk6cdQpbn5R/hhIgvbU7emqKk8Jrj3U2MV6S3iHs8SIeAPQMlU3mngPMuvupxG2z
cBtNPFQodv/m7hpKZHNxNvyHlivWHueFK4aVcbU2hTQDRRYc4+bxuvLFIq00aLjD
RAh3W5nAcjwbRmJwNFim3VohbLaPNrLyh/40xbf8/ZovViXtVrrmegayVGDCQCWm
UskkfR/sUtsOjvKHAzRiiOf534x/d3dbiYe25na7C/A86yTeofsJYZtReZq2r3GR
sUP86evugh1xV6ktwuIRpcYdOJh9YI4mMchZ1HPVKeiqgwez5gtD0h5Zz+FAtSf1
GBQ8oxXi3T7UIExz08mlCx7e+poXm4GqNtyJKF5mLZdmeYlAbCcWqyN9SeEsfnhi
NtbI7upZ67xJgkYEZeJhz/L1Qa0P0QT4vYz2MMPi8Alrf8bdFMtJ66JrjYV3BUUl
A8FyM7AfAYiKZ5z0OjalZeifWCNACd6Jkiq0GcS+EnqeZI9QJijpRcuUMQdBZh+P
QXyxWIDXT1GClKSzPsq2QtGO38a9wjsIQSQZTxQm4iBpab6BtQV1si4Se9vmwH0D
ghBsQYSDX4k29VSpPqLDqzQEdJOxWfWqC11swRs2Nwy6i95KI84UJVmK8FszghzA
LGD0LHy8vOsybSisweTmKAaFd88GFDxz3c6P3avoXCHcWH3sLYNOGTqpVDms2w0V
nhRO+nL3yx0NccoZ4Ktix8XHNtmKJX+4IGlEEwbDKY/Yd9kqX8fLrN5IbcvbU35a
G3vDTJSFFyMz496lCG2GvLypp61eXjgtiZAsDW5toJtP7kW+li8YgY/LN32nXIOw
v0Om0bxb+azfKhp9vTTdZtaJGsgtvwF4XWhib2NQWt0Mjxhp5MD2cySJo/Dqamj9
6YoVpDfcZJEFY4quZ5RAU+2L2y5aVCUN/lDtxDuFsSA38h87i/FH/PXwOoIV8n1o
8cEcI6oiw44TErF0pbZHUz9qI0CeZNsq8AqtojoJ5juBpDd1dFZBW4OUj1G2EwDt
lvK8dkRLiKNf1Oq+xap+/3vgRRZtj1mjQbpZGpUDbPaHTqoqFowDsuMuAUvEt0Ux
qeHdqk8CNlnyuKhQh33BjpgkwByONIpDtQesJZ0R5q6bKlsfd5rH/13qFSZ8uWcN
ry55fqGfzs0zFNL5D8yjnQuIk5F+lulbmQv4rSrpAr1+Pgthkm7OoT6LiHLlEWzQ
awbIyQUdPMFYFTi/T2u/g7hsDIavsy3I2rSzwUAmINY3AktzGCNMCe0xKsf9p0mU
ShqbDdWrWM+hXtaGdvK4iJM6c1KvQuTd8nh4VbFGGsOF9Sn6euQ29H35n9kvmq/n
uB/d2MhHp3evC06USSL6XX+Gx+DsTwB2TRRwHyUAZE09/vGxQtqG2FtQncm9NBWm
xubJ4H6DK3bqtvwY0NDS+S0sgpODFGHQe7YhB70pe/iaMU2eM6FRibknCZJl9fJq
KJCqJuDddwteww7Kb+tnz0UdOOc/uZXOEgHBKMde8rvS6U2SNYO7kLjnKlnOD5cZ
rq6K/J9Uxh9ZkU39OmOkvfrAEdpbIcl9Q9aXdgFu2KE9VoTYDDu86nv6NierbEw0
XRnA3EAiuWPDMuX2HrL+w/mvCOgEZ9ud4lIpRVGesE8Wg00+/l0wWziPIdWMSdRi
4EyDsQZLdlOsaNaV5y7LUQvkYRL0Qsa0NR53JOtcETiLUPxuI0pjv/up+hwBex/g
qMNCr1Za7EiLt3v742za4r2gRNUWnKZuTZOc1NBU0U1kw0Kt22zbq26cuaJMylav
aj12+07O117P6aYlRWg1xJvSW8T3UEY+2J0l4nCNijDgS90wi2T7cf7O73d4jzaS
2wSX/vXHFkflBONA3F/oLEkSg+ghlG+YMVSK2a/t5eFzEsrF67YH6x7w/rm/M379
H4Y2Ag/BhIwwfAjLDaotDtuGpOkM9NW9+21ItX5ci20fsOoW5xwZhb4zxVKGzX3/
MxYTIk9Xxm6jFvmLncbfqnA/DQ5PjIbztWt13/3fRtT1FVK3DPrF2ZiDqzUr2S3r
gVCYxiDFnQcVZlqFiEWh24Xyne6aMt0LQUhL29IoMvt/AzzZMh73HKhu+O8sW1fh
dxm8C+tqj2wnmd9O59JsTKaHaUVavLIKVIngLsgv6u8ZX8qK5jAdQFI1Y0DgkW7q
yXO3zzJ1QnujEGrmC0aZk3O5QSL9P16voGGapJZq4T7T3nOM7lXIWKBsjW3WNJQm
BYQmIojW1ztVyCPDxbS+spaDgYJkZGRQtkaWT6i1kuMUnKUlUayDgbM3vK2ydSVC
exVN6B/IgegtYehwZr4Pnewbz7VMAlTz+C3G1wK6wTTDyBXpZ7qylWrNSI7zfTpD
fnCu16+7Ecggn+ezRPdtUchnNXCx6gEGh8PIuYOgbaUkNmXsGsIdLBVfyR9SllZ4
/6J7WCzERygFzLicByBbPsRXeKcJf3XIcoMfiBXcHbdZQIICXzvnMlCdp+uaCVzz
4SuI8/tOs2UZt1e3dXQEx6/SWEXkdvYQwYpOPpnnBsaFUdcnIXURoKSXFUnk/orx
C8KgKHhnYJvW3NoLxCvovN56K9uE4tdto4koQ8/7tn+ZlpIVa92lsh4lBt/8WJcL
USxKNJOeDMeAnNcFoXcD+16nB0PW+K+nsZkBCdF7AkWaTw72iNn5GGq/BgDaMKBN
L5pWC22J6V+fWygGMpAOFEE/ixDKTiODaFyXRelmtS/vwxvQtrIhJ/VHe1ehvIxl
NZPGD4gFGrv4VUEmQj34gX3Cyqjb4ckvafJMeX9bySDnqrLTXc6mvvz2BgI55aZg
b/1vyJlYUksIDy4BcNMm3kRjvo+s79njHFhse0cJEnGIx21VCjAYjo1nuHeCg2h1
HY+30+mqACHwvURUrgd2SwARhwoC8WWgzeVADyxNO3IlVK3pdvCr25OXRM2FT8cq
jP6Y3hJBVv0h7Md6SUB/GqH5zdahjBQBQlIs46MQyAHnv3IlsQwdk5X7q5yGK0dX
2ynL793n1QpTPVY/pJAPgGr3Phul7LzpKB6Tw7YnHUUHWAZ8fspeiOm4yv3kI6fm
TiPb7K2dC22cMmkjljYE4UK6IJXdenoQqtAPe+nK/CiGwixI0sfS0MkO3TFow0Al
Wzm8YI37T64nAu2NfxKQ+eruKvbzFfhyD0gqHZdNBbwo7CgRYMptUfmg/PUa1jAx
DiDb9h9KZ61mlYdk2uTeUgguIlNIAUETPJE+khDHVkk5fYMQm/kt8MfzUw0UoYr9
57CqQtIXpyROrMotJr+Kk+iVFfW6SI40IZqIQ+eyo+ajRmhh/EkzDzIgxlAf0bgc
1kAakbrkehQcLlmhL1a+2+2oDzCrU3Xg6LFIzWEz4zNgHZAtP6V1KbAKQbGw+nuc
uBOAzUnd4aFCwDiDOEb7r/y4Kh355A7/cZuARbtf51Uu0V+8ybK26AuEeRAK4Vhl
5cIc/Q61q1rjEToA3GpfBXoOJ9f8AdVRqe+uX6xUPwfDNGJSeAVk0JoHLNBKtClL
aiL8Zr1SntE3Qih78rnQyz9KW4GomogdQ0fo+iat7ckkR8wzlSntE24LGiJj8+zc
X7uThivY6l918nR4a2M+yWdZYoTWGuLkWqwlthdnNqZ1psuMGuDLDTIcGdM2Sgt3
7io905HbjcKm3tIWd1D2UgIXWeG/c/At/SoUfLZn6z5emIERQgYPxprJTfvS0mD5
nulIMrdQFv2wH9QvmLIK4WclfHIQi7yVmbiSVDB9hzhjFVfKChz7NSU5HzKh00u3
hQ7d+bX13BCs300Q1HjuLdZG93eL5sgCDj7AR/UXg6rfxXpyTdcn4yLZ/2ugbzT4
kxsU2ZWg5v/IfEAbsrpj9zZR+HGehGbfSTpin2fkjMPdVZbFl1M963wfFNReV8FN
OMHrDJWNPgIupqw3iq4qxBsFZea6BzHjdCuNoiaJhg15cwxM0YhT76Vp2nHJMiF5
7e6NG2NGDXI/HEmmno8dExpdxfEZIs0cXHVxrEtFE25Lvdwh6CQTdkdsn3bn2SqN
CiE62amecWAijQDUIJwtrN4s6//pBWKxnAF15Q9+/Y9K3xvDVzWz/viGE8haFnpP
tBGV1Ty+FVhnX6hI7AcR3HK74BcdKnQnr69Tt5jNeQ6fsA9Aj9cAN1j0Df5T8P0P
TC8imc4fYp+RMfbJmiGRWmgKASxnFhSj8lnH28hVlPnjhdDVS2aoCv2dC0YKHBI/
cl/chm/ja46PpCfvdzlnJOeXCYqXS3GOv3nB8iFcLg33LotzILch1TbHMQfUbFYw
YyI9RHdeLbGp7a+uVrqCB8VyuNUcImdJMkP6vi/oXdiCF30tVE6189/1D+m6muIS
Skw9CXGW7Rw5ur951CDEpDld50fsDrD0k3GeTrs/tWJFSrx35qcorrsLkJp74i7j
XrfkV7YGqU5pQforJG+NwaLElZxoibkgmX1tun9M7qtbIP7cvipf23QAkPq3IPh8
4n1UIuMBAMK4uX2vyUR26anagPlISmk1Te+Pr1Qr8XbgYc2yIeSIgLpxGJmom5HE
JPOifKUXaO8dLJcQPtoWaUPxf3x7SIQWtkKa27u6iWl+RM/EG2o3CoZJe7qi8ydS
MUxETfPnE6FZkT9gch6P64b6e56rozUOdkH3WRXYxiHF23Ergp+5fe2cZV3HUj+0
7946J9rIhHMPP1YVT+cQFmFuIW8FvI0pvXZsNqA98DSEvRGXKcOC3agi2khlppHu
FstrniwakxwbYuouAcQpOgErFHQhfINULW2Okb2n4T4uRT7MYzyVPipgFXHGlvs9
o3K8E2+tAf4gaK3MggMrrpR6Pw3hC+2fnEbR6OmOjgczURHnn2mbfYMUoLikge+L
7RLTFtRPDiE0dkHybji/8NLzEGa/7SeVheCrUuQvKyMcIr2ZxRxGaNiIrMAVcCRH
bIxxSIDfYEH3Zp33KmkgiBwOuEDvzXmk69mzwLOx1sFhxOpgUVroQKq+Xe1Rx7bh
pKG7C8a9RQabgbbTpjmEu6TB13ENF+G4/8eIyPPfm6CNh6Xg1VaMQLUhgtDDob8E
n5XvXkOXPiC0/5ZXk2JauZhsWRAaDqdORkLXzJ+2sYLkNU/W9/OiNKSuLPD/gwMq
ajhg/LLzyMVrCcckZGVJSDpa0KfZikeaJ0fpVisNI5ex1T/jr4p6VbKysiQGZc+w
EQBwg+03a/l7q9QmFj/T8gUKuBLju+z1L3Wddpi2reOgGNwgWIdpjFSKs0PsrDcx
s7gcr/oLDXCx34SaDqY8CgsNnIppb5Aeeea1qEskTSDcf8dRmAWKJbaPEHseVKkm
dGTXbSYV8MshR0jSbwDFbC4Buu77SMWDQZH+MDh4Bh60CF8tkhPsMR3mi+do6gfS
GeDVkJNgXTMTgVJek1bQbrzz+HV1646TpYWa15iMBais4EQjfXAwPJqQY215a73s
ScyF5s5vHiN4tNaBR2P7Ej0iF6wFtE8lN9ITtSHh7DAaSF3aM4ZQJB5q6zcJMcWb
2c08qMLxtAoHlN86V1kPZf7HpycK2jBVt3UOPe+7Ua3keYLYeM8cNSzbhbFggg16
cCXbGWL9Fry4ysicUYOIcEXa9yFGIhmVG0ATD8zrTN5p7aphrbZ8JUgMOvDuW9t1
wDL3Egd+P+RXsGHWJAFAFmyjPZeOZUBcEHYxziWH39BgfJQbqKGAskscPCng48m8
2xHp5zjlLAHtRAeueaZyj7byQxvEmdKL3dstAlROwKsbFJzJXmG12uL5HHLGnXsY
wOYmbfnPDggi1k1J8hVpIhqaJUnLPGsPa3FUdaSG+5dNe5mK3KNKV8m9rDgNQKAf
mBUnRgeAQ3V/p1voOrS1IqGJMTeigyhgbitvcWwYVGK5VCVrmEvgNenFwLqlikMU
RO86rQBXhbSHU+Yfu/3UKToueyulszgl3Aj03I0gTy0TVrxpO4P+AGXrsU9Aybz8
ovVqIDHT+hxNzKGpEoQme1wss6kR96r7ylokaI6jdRqx6+uX7B9oWnRRq79bYUDV
LVz2eqYO6S4DaU1WUMZ8hcnd64897SF27rMJWSmqPFB5Gd9Ti433nRNrHuAuIQpS
CmfN4My+j76SZPSyDvokIUb+Y+ZDHepOEPp97c8WILLCSdpXHXyEXX7WkQo+upDh
hKRhBdpZ+hfkEZVkS+H5CZnSMHK0cWfzI2O4Tq/q/zH3g26lA7cFZ/Y8nuSfnGDW
y+X9AznlyUJr8Lt+IULvUAK2SdEvH1U1eN4zo53e8dSddMr8eMwtgnzikmg2LvUN
ND2kfb/8nX9cowOmt+CUvwAAlQj0xNq6HMbpaqI3qR2alY887/sgPasn1ai2Uq3u
rP9wVimFEgDIZKMTUoj7tdXuUcUORzaU87x5s7omhIhf5gfoj81gz7OdE6NDD1++
LrIjtblkMt7m+FjTRBygVQjD9xRT/0qg24ApwZE6MCCUFSL2GkEoeHioM2fa9ufQ
uuKUf5glwZdY2UPbqx7C6d22EHyZIne9wAH2tFs7y/M0j5IkRDhULqUs6FWCR/1R
SNznMJzHRgYOFPvL849o81trlAh5wSksxmRyVqV+wLY6bSSL6O6yfCW+h+XRsSEF
5mk1v/nsTpDiL1DgxY4I3f0OHr1eK2RNwKIAPYEcjNn3Q388EfiMm74yZUPSlo2i
mAL59z14lR2IuGaknOYCGO3SQDDYySrG/F6vJxGP6mdq22mAEjpzgWwDOAcoa69j
JB1we8fzekgEfin0vWnzSePiFBAngAt9+fqZBd31vasmR2lgP1/J0ryaXbfVVHRn
fs05UaunwVhCawyunCVhM3iaT2Fn1QMLESRK5zadsSM3Dj0aHJHZh6yCSTLbjs6K
auLDvdbmQkkf/CUIF3L2rktYwGi6ZLNBdqS8fJRJg8zqGrXQS8nBalExYyOneREv
xV+ueT1YkBhpWSAIHOj8hj++LqeVQS2uX7cPKi/eHmcrt6IgC6vChbgCGxy8j9OB
sFDCoSIp0uy+dYj8dQ/gXwgIcX3WXMlr2pNiqKbZGxNnCUOWE30lN/VIiRbhC3mm
w4o7FQvkpaWtKzdLrfxlVDVNvNiokU/fy7s1W+Pg4Yr5Wi01ThTskyvBf4depTZY
+qAnd7OAcMw3voh0N7c82go6he8eyFovfov/E5jBsvGC+mLymHrLFICjcyEupAeh
xbtEB0s2udJxBpbrSr516XL5IVyOv+SAWFw7EcCO5p+W3lyVO0MtZdkRGWaRBIZP
zdO37nVQogQvp5YOR15J+5C0IMOPyFdQ/WOD7eCEKEhbJwwcsrZZZzzItEFolkv8
icw4s6wfZLybvhf4r5ZilieaMMXel6zMk9HNrirIMYqjrl48nfhOJhVLqcrf6MJF
vVpAkhjpgbjMhrw7rG/uCFzmy/J21tKCWRfe4nzPba63vm2T0iNClB/Odkqk9XFk
VnW5bjnnCIorbJ2D3RFcT5G664s/s4SRkU/W2PfoioV42DKvvtnRoJ/WDzeDXUfu
jXrMw8qpe4PrnFc5OTDi7pIrfNovcgaqJizYAvzyB/nkO52dvln6eehI4AaL3EbZ
bcvMXvAp/+nC9xcTvbvRq5nc3BL1Z6sygKWLPitcZQaRseKN812/cdQxonEVqbwA
fJf0h8J1XIKhha4de8IoVSApEVaiROvCo/7MG6xmC1AqE3FXfKf0ay+a8I54AUe6
VGMY9ibeP+Yvd0AdMy21aV5nq2O51bglXN822uwsYh6PIXAt0FYsGuPMsW0iG410
r7HwLsZvTEs28MyzO6XS++Pg1y9j5UlPnfIe2SSgUrmdzDQfGBP31gP0AFGgN9S7
F+Xn36pf5rTvAdX+aXLD0/Hcy7SPap0gOH3CzEBOwSC7RpMr0bTd2kiOXLAPurwF
Ke5j/uDiNGB+q+cT4qwCw6e51neeHB++YWE0b6fv6KBm67IOIj7tmON+GOdJIEqg
ccOiKzj6u/2SqKnB4qBemPakFyazRcasjp0aHlPihbSOaUQhkW8cUX3EXtnPfEd3
HRreOADn7klqcZFJ0jSh0fPjK484uqVkH6UoUdcwe0n2HEY2Zewys6zNI9T8HvCQ
eXFqrk8vyElCvKs084mZkg4of6Hk6dtsGI+iUaGpEIL6JTXaxEsvsv+aSTXPcyiC
81zGQfVb8gATI7yDkwzX436NdArwZw6R1ClFEXVGX1b9SqjVsHDiGZINNcjzCqxP
8EpOBCEiZyLYXJfcGYzNXj7K/7azY8mHw/y4h1TVdquf1qAZJXEjvNPYvyUzcbBL
bHMLae5pqm1jwfR//GxxMa6lRi4aut/t7nYv+/k5ZPoDl4OAEK4GqNEjOOdedVbQ
qPTGctO+XM7ix8MTP1XKhhccXel4QTX7S1/QATLgP6k1ZpzvTRX5yt7VEFkliNLb
cvTzMn+V2LbE+/3vUKCB/h0EMn1+sEIgPihb1qLIpqz9n+uN0nucPtVguu5+CGfG
XKLd4b6g60N/8gEU9t9IXPBJ3tYVp+orYpVrGqLRwVeaD6+5PJ6/Tm8iP+yaCSd+
6LTV7e7O5P+EhFrheY6nJsXKst6BKm9lGnbh+TcD1bNOkXXLnxAWXU1SxWPErqIU
y0AOzgldnEgOL6+VZ7Be3M8hyux2e82CkosWbp7id1YfCbPl/6WX/px4dOCGW8IM
2gZvddZA6vFo4vs/Cbm+Wx18oEGPhpLNYrTY0Wob3qSZV7wG1NQ+Ed4EsOqBI2B5
TbCq2HjFLcUZK6IQIvDb0x0iyuh9hZ5RUtvssvhGqjKH6gGRsrSlWV93hD/HYmsV
mOnL5Cars+R4WeEzOmWJDNhyzZg/Ho7+X692tHqWwRWSo09tb1aImXjXsMfeCfxh
oB9th6b97/qiB6Qz/LsxVGI2GifnTc7BUaFwlKW54FWR6vfrG+yKLnUtI8tK6PRs
ooUgf5ylPHF2FaVaL6bu47akFQWsD4us9dGaFaSrJ8I+9UQqouSZOht2c227VhJT
tZ74+LmCQkVSD+cCYy7+sGMZTUCOI4hOFVD9AKIymPG4UZ1FlvZvTOALBr8gDyG8
uzPJ+igcEIkBkizvcAE7p+ScaFwYbmb63vT1tJc+SkMkO0rgGUnCgq8N51+k2oVd
YxSC8nA+zHmN9MPViV8cSQIe3CDL/T0YfYAXiQId1IFNmBbSp8yCuHWgXmrpVjTC
v4+CyP4UY6XPmBO0T9c707gY9XIgneEZ+o5S3E6RBdHoXQN46WD3zpyxdj+AkQYc
sfRcGGIrf1/w61k5kIpqbL2pbqIunYjX6smmumjWLaKeunVhs8rskbz99wlcZlrD
bzW7/aMLFcL+sQxrgMcc0etJpVDJfEELkPcP9KUaLiNNkiV1HWy03OTP7tkJIMBy
5V2OD8Uj1t1Vp3P3ZyrLj3dIysxImfb9APKEnkjrJiJCQhGZ5MinlTvLPccJx/ss
6vY2EVvdsEjs7f/1o5Zze7lBPRBax0KaOYLRX0qrZHrXgKYFssAJidW7IIku3VoA
7inVbOJG4B7r6GKy7yRIPoH3YKVAoNVK94mQztonSMiUavkAoFNy79iqX7Uf/ZGU
7/zGZYdm/3kKlYigZJDTLylZBZJZCEMrIgjMoILDXIYZeGFquadqzx1QOYMelYo+
HuZPNjT0wC4ZHe4neB+++ZSt7+lW94nYANq0OTJm90H7A0Qigl1eyTwxoQim20sm
CaCrYQxrr/1h2JeD5UQplmBT9iPa2Owh3Sz1bSm+VKI07MPxNQ1PwqTE4oWRYrdB
NazwVyf/YB3UXS/oUGT/vvLb483BPZskGyUsflR+KiDxjuBlQ8LL5goLq2IVgtD1
heEgtuoUIFrpGD+r1luOYWPfdtbnDghQuQz1/lZwdyQDMiFs8GZN4WdBdq9ix1F5
mSvQYLyeU14etpTPhZZMSI3jhVLFJ+QO2dfNwz0dYEi5q0c4GpHH69N71zH1hO5c
GuPhVMQ8H9GAoJBdAb6PNBLjergbhYEso+Xz6Ym1sA70PtzI8RFSYursh9bY+Nm6
88oke2pm7TiBe837dOv4R/ChZz26kj1bmYnPbOfkgW2O7WVSqfml44mzbigntzey
2BlW24AXUBGN4Mtk1XtDSMwwfWOTBRN1Gi1s99wDGE69sYbsTlzCeXUnq191Xf+v
5NIcGwi2iQxExOEDdRkdLB887tlVGfLwhozttMholrhpwkhg/KsLdw+x0DPt8g6A
9JNhUgD/UVjD/bJQYuzczHaTGfhUskAQqbdnLxSVOsy0a/BLQD18CCcooNesd73M
wBY7lQkkAjv/S+3X3WoVwKnh7SpfVZcoBLTo8jib7LWpMnsYGnBTzOqL0r9p25HT
xOpQqGzLOcLwOiRI5yyNOo24zOs9aDPCoDfn4rPbRnxKeMq3uBPRfcSnHBeR8Wvv
lg2AhfMnewSdEDa0Kkdo8FH1FoKbr9nZ43gmV1Hjl2Xf7Y3vBd0ZOhZz11riK+3w
77PpDaX4hhSwA+l+0le0NRrdoz6oQuEGrexxfZdZQTcYVOs09lFs3LxuTfNdDy1Z
ItZav9tBxkozk/SpVbXKri1ns/WLhWZhwC/CtXgJ0A/m9zO4bHgJtbXJPeRhTbab
kgS5vE0bU97NnKdF80+MxdfcNyhmndLbN20nY+v54DTY4YXNHKoKW7Krth5yDmeY
ecGWFn6VPptX8X/53RujExBkAFKhH5i29UAJ1lyiqOPhVIYM4JHIIZ6OSkl0fQnJ
6E3ShZjkTJVqIfRl79OmkrdDMeBE4GOvEfG2gYtQqRfaTvAM7rKsu361JcMVetCB
6zHjbMNPf75+rjE76amR5nzZkMAywCqgVB/BHuKW+D6tXtdbhU198PbXhICxSP7a
LhACp0pSO+3aJ7RsxXeemcwNFG2JneaA6t8uqQ2MDVgQaaaO0iHOz6/tnz+TBxWm
/FPUvgqgdj10w9yw6ENQE+Fh1baM5c1TrAad3nwi4SdXzaXSzhaVi9MYxVExSjJK
nfKhdX3Zr7rVM3v2aata82Z9OlrxmbwDrkG8msB15/U/Tn3UGP7amxXk4uZZS/DJ
ypc7zMmiA8kskm6afqE12rkUArWwbmAQFlkjCN4NpABIxK9WudCK/6G/S9pV14kM
y4YZZQmfpoa6MblfjyOG4RehNgoRqrdSRTdqG3d1+i0ryPtEOuiibjPzTYqTMnyj
XiR7TriPWCru2xGBOJANhHzDF5ZybfA+NScQKctv4m/PHx22D/nngH5bNKfOFLZU
nQsU0/3rre0KFw7EzQHP71N5k4mWBpoltVfxaMMyu0T8WiakSaB1uL1rczSf5F4F
9VPs+GsX+yxw2I/QCNdv2IXcVxHOtFTIlXn8VEIngQi2/MbuD8NVmnCFwbxQ/tgu
Md2EJyyKOtw+6LoqdtNozRn6cVeKAnLHKnbtZZ8H2p6ZSDxK/wWMR/3CUAlHkE1J
18dH6hhzR7IUBry1oBwwDPXdnk1vEEGayvD1R1XhvNzPVvRCcsHAPeABKljHUUm5
QTwjJ6rbMhEb36isjl6h+kebL2hK/C0uSICDCLvHmSdnOuB7w4wyvrKrjucrqaZ9
iNdJiQjswKlV1E/P9WtWrl9HujOQcpulgKFlwifKp1KrIaDbWjZjaixNVXFhKPy3
yNODXDFx10pDjkDgaTNANMdIx6hHWIXy3Xw01aSj3cIFslXd3chI+QiYJxtMnLB6
BksbDS8VtKXJM2r4WKwNdvqQMd8pglMMIS+DO4MKnQ2jEdUiCmxOS3yhmDtzXoxA
VIhTWtQ2kC4/HJPYtb76fKg9UMWTT8nWjmQvK+ZymfetlHBJ/8Xxzvw+0STAVi8F
pn5IroZfDzqar9LJPErf0ZfjS8jfVPM+icEGCSccAB1gZH8xQmdp4pfdg99xfwbM
EhbSLjcgYEdIXNF6PogTn/Hc0rtmbO+N8p4Dr0nh4+fG3QOBPxQG5m5K/pJaY+Xg
BewOIzIVg9TidJv2965xkwbcHyiEwF/vTIPlJsd60nrdNx+0mtAuyhGvSovhzOu1
0EIOYYpLKfZ3FqIw6c/ec759oSysktoNb+RtjeWNxtKQdfQKLTtikeDo+wvm/mh/
XS9suxzKYzt8ZaJRYVUGzPTsaiZ9rWOugm3agkb5TNpO28LRdpVxzOv3XcMzyUCQ
N9C4qLF8dRWLGjaArAx8kvs3YnItBranjEa1liXwnGSYgIV193dR5mdV4thRlpY0
J5ufQnm13CKOtRJo1pzhg+sfXspzMsvJbn2IYlmiW9KIRACQNEKigHlZ00WhCypp
Ni73yQJNs8HcfbR/cztD9/sRJ7LHYUT1QbxhXkXcF/QdluAZKuVDxHwGBzASg4Fb
CektvjX+npsmmPABkFX8KnG6F/lCAenQzviArl8VBptiZ4jfqjk9uGQiRrlA00MZ
5n89QBPF+LFN/5Q5/E+YDYocCeKnXKs66gRi6Js7uUObw7q0DmeKqzwItCunrNCq
pY1CFmCks9G0B9o/pGOjtLthD89FqxBrVk6M4RZKPZsMmw+8yTezNlgAme6Ti/Y4
/UkXhYSVAqN8psAfieaoxe4RFGjuOaDma2Bz8/sh/hkg2z9r+klxocFrg6eyBiF8
5soz4AQvGKqEcMoJ2iiHD3rApmkqF9PpKu9s9aX+525JDn4vAxLbb4uOhXIxZLAW
b2d+OPViLuluQgl1FjE6Zo/Cw/r9QAxdnNCwZvOdRfFYB+mr+/7dZvNLleGuXyPw
3KtEO4dp7KpGRO6YQhtG8WU6rUGeP+nKBkvwSNh7x+alm7R3j2M40m+upFFATfY8
wzMygbIzH0D+u0ExFf2WqJ9V4zDPTIjemBF7x1u3rgTEeU/Y65vLUSu8tuIuPssa
vivACBmohIy75jHgEvnOADjGDkDPrhu59+8hVdIvvgwoB4C2hifDJVbHBr27uP/J
Y25ihq0LZhe6R0qk09/wZ3BqQFQAuPSOZlThD/Uvsb3RV+GLcKzVWTm6Sbn8GCcP
Oza4eTXDkfGYFW/Se4QgNFrnwcgV7Agq5+jA9lQGIwvIzRrMdEfWPrJ3cIQ9FVYa
/TPAXKNAwBeir08zizO126RcfA0C6PNQ6nn1gW3LowgVTrnkXsYAbk3e2NRR3O4M
SrU6F8dPwFAiVOfNEOT7LpCTmclukuzJqfT2dHeVcd6l3XndxzVn5q6w7gIbKleK
H/65QPo/VDnx7AjPRpqy22A44LFJGJEbz8yhXCYJVsVxTAhLnCyrE9ZgjH66tyCs
GUXSf4FIOtUPuwPJuhjS7WjKf4P5WOFtac4iVbulKYXwzU8GaMryx1oezxxc6pFR
4cqca9H/IA1Dsa+3brIvJ9E+C6WQKAQu7RFqQVj1+2IJYwyHs2ty9+wOQ+DasONS
6Qv3J/3i7EtGvHbKIUseLZKHFU6A7JiE3KYZWQ3bYFBNoEA7LnY7BJU0DXmqEBkt
lB1flkNliRtOPmeQuWc+yqgOQyg2fC2i4uuslEUA6QpYvqWbmzfTeNp0wAGApw2f
rTNyqSSzOVFz1kHEj2cAl3MCrTmRdUfqM35L/AaN2gGzDEdev1vScYzipVl8iQwX
4QtrBfxMpPorqMfE5LLcQo+841lzuEfqeb7GzOKn9tPTzkSSHzZ6xLhnYm3lS3AW
taDxNXehQkLK12k5syxJiWzWd5i66Gr3oPq3QR6T/0zdjB9r48AAJGUcoSeIZPx/
MB9jP5vkaDfx2S4fFl0VFFP9x3KN7RU997qzxpytVyS+/mwTiRRPY2t0KuxS78Bu
7D5t+WInP0IPXNMLc5ICU/cMTAYRSXH9Vk90f+es5H60681w+z/7Dy3pVaNql4f+
OCKb2E+21XSys5/j+3ldkVpiJgdPK0K0FmGd2BlB/EjzZPa30q3AiWfMmAOjSQhB
ev9/AdzVUd/IZOLUuii+ONUNsdVrCbr3M7Bzv5ms+uV717T5SHOryAKVhQJNmwOF
mgibz0hO5qxoIyxNudshV/LZlevxH0JqsINYYx/0JeM/JvLVGtfsiYb8FaJVjBwC
wL4WlZe8loWy1Ea4vVXjFkhmOSfM4EeOrGyn8FpzGBSeP5M8B5Ohf4jHelQ8xctK
LstexdR9Ih8DERaBhp0iAmrYirREL8RCEGl/vLijGRPblSaBqc9E2PLcWkucVC4v
GqDjyhh/wjpWSnAzwtKtHlGCPiNHQ6NegCUKzWsv1VObieYLpNxWOGMCcJTBd9BA
JQnNrOFRPtJeA5n33s0s/celMO07ylGMRVYXSjj1yCM1e7P9K8y3qI2QJXt5mdQJ
xSl4OC0Hj7Da6fP/it+Af6X7vftsyDIQ2QLoK5tvdRegCBWkGZINXmVQ6VEquDTd
7kFXHm/VbMceXtARC9Qg6aLJPJUbF2iCB61m9ucreYmPOrU+3D6JscNJN5gaHAEf
3LOiJFlf+0zLRVBXnfq+WlhXOd57U+S8UDFfHP9+AX7Ge6Fa23m8rypImbhSnpmm
U586YeOVQrDHZOdyYzvlyXu2avtdNRMZA7IJXHkG+6sZ1VvpO056698l06kvKWxs
ib7ISwpQiGWXb05xP9Ke6fwBwe/hBkTpVqWDcXOnLd36awT20Bkgfiz6IZviLWid
eckKT7j6U5MEk+kkNc5RAsbg+4dxCe5zXUk8Y8gpfp0TB3KP4C7zPL8Oz00wnt0Y
v9JJnr+n38K5jltwSMp0clSXzG5qM1XjYATGOIZc3H/vQKBTU6Jf1szmNlMqzuA/
U11odHY/ix2qtGFzeVZ06tYF3daImAYNDYw6BlYEJ9CkkVFhZNFkFRakZqxMZ7vJ
lyWhCdud6DSekCXsaFT1AbcKjzwX3BTSlq40DYsMqDn5kfLA0SzmDL1MweuwLgOa
YMKyOFF8yqduJqDNGk8F7C+Nte24U4sKIEUOwlcwFkiqcTQ5C6f9eF0KRK0GyhHA
j83MIi89HjrvqQBvN9nr64uiljrId/2k6U7NSJLNMXxFE8p4P13dsCthWX9O0rM0
QkDyaLreQrZGujqGaMAWmyWQziOcq2wkYWL1fnQi/e6/bGSY7+wjb6dp/PXH0eLv
AG2yVsgFh0BiZ0qlc5EvE8LexPBmiz4dgR758EOwQ4ACXX8GBfCGnlIsdZBZNNWk
E1EtdVx839NPG6/gHJswtsiZu7d8O1+/gGDz9ddJmK5YIXelflypX54+vv7HdHSm
75IuyDI8WrZNWDpOWFb8Wf+GCrt6DK6cAorlrgjA+td8RpmfFlfF5gAKcVmO6yTz
R/ZAZzbYY6/6kg1DDJqSKxuRE9r+NDHshjRymOdHueCVgX2Gep9P8M9HKutG3BBX
qwJ4l3atPsqQt70hfnTUgcMjUqKiPLmvhY4gKtCxmo6HhLgiAiDOJNH58dGd/mMK
9QQB+npT3BmvoyMvynehWWxHHQXIdw4qvIb3R+bu3fgoYadt+VVJ4ItrcU9FqGL/
vmcqIId5or9Ooq6JAHUCbQ8taPRa2Lnn7qoFLYE7JwT7ZzicKnUE8xBi/hJVqJgZ
ey9uW8neP3D8/3uF80ze3i58VbFrkDrgUJEUrpQD7E98JMUEcj3quwXg5l6qwjEn
YMIv6NOe3cnV8tw8dU2H5WwbYKRiYPp5TBlUrQpv8iaLMRXC398vK3jXltiYJgH0
iwSnTULRniMtv0f2oKLFmfolq8s609yuhfLxsJuu6z83AD37WowtlFMomr1wglOo
Dsw8Q1Xrka4ljrJ2R/iwAQFuBb+f2CcQbvmIHCs2lwWBftnyPpJobntAorXlg9FK
bIvhmCBA9CVngEbcyg/M9sWrBW4Sdju5RIiesKvonyUDbQfWAo+JSKiAbXFz1QRb
BIcD0MjXOY72XLz1lzb2KSJA1K4drPlHMuqne36sxG6OBqAUq7dhAP951pcGGVN3
IE4ML8+ACXBoK7DlIR49GsZdX0zdMTu9sTWr2LJ3bvYnIQsG6IVYo1dHuAfs7nqr
hwiyHc4pvpaZILJxZgUxUcpiRFxJ/x1a9sEhtKg640z6gBeQKjBnFemtZFeEU27b
Ma1oO9uwP90w1Y0PbqDYfkLIxqMZ7XYx1xddPzR1cbharwO/CGwwBhypgTA9t7Pb
jJ3eXjgmhh5KVsml733fnP7yRLF6yOLCmeeKT+e6SL0pcHQELI2MyEzeylebyo1+
Tz4AgThg9W0Agntg14+OSbP4fwY1+ObGjKfvA+lCLXDUWeiXphN3a3Hn9dibzt4V
gD70A8brjDA209+qMrsPlMhR2d0Qy2NSNC/b2K85NbZavWc1Qe6ckMfupr3U7/3V
ES6Nv8xUunQeTU6AR5kgZcSOSTkioiztY8hYT6LKY+2Oleduhs2uXjpxuiagjrpe
RksWUrOxSgvxAjpsgFP/HdnBzOuQfzYgZv4OzLfNPZrDgzCpxb3vB78Shg9ylaH0
F0urmPDlEbXQqawuiv/GlOUGADGSQhEF3DAweZGLV4D+W29AwnxNyIWqMkBu4OI1
PqThMoBu/i4D7EYQuKuvOWZEm5TGyneYkSmE3ImWjSwDtC9VuFq44SLo+W64nKGR
nDVXSB07QJzMIfhwTVHMR4D4qBJ4eBvt8slRVL+xTxM1lQQxwsjdDR1dJ3iI34Hf
7B5ovdV2evUi7306STQapgE444fqUI1zuAXaIdqInc4dR+UFDQmx3/zMBBtLt4qh
7KEs8O/x2WG4qGMf6HpYsmEHuRgzl/UZMXyN4pLn3JJAQ0PfVE/yg9KzZHee/8Hh
/kT7NYFJAiKxCxNuCrg7nU/uHRLuFNfVkT+ZSlq2bNcbJ+k09fSxjS4S/tCC5Kyj
ooMkLPnPpjO1KE+8+CcB43vyixlPIpvOrD/Dy2lyYK33RWwI54842NKSRE2j/iZZ
t1yj2Fi8jFecktuepVNXiUa9NJtRpls+pq0ASCKfuhE+p7XVtXkRzGDTL2B3ZFrd
eKylGXd5wFmuGLBgqqZi4Bhb7CPNFhrC/rzYG15ILfpVjER70fFY3enB8fNPImNF
8UHU7crSLQxhNgIe1fBvHf2uQ1D8snUpvhH84YBulP73h5i2lnOap9hdeW1gZMSV
FzbId6A0haoWPN+5lQRhQGOvtI5v/uDjiEHnrW0lYTcIFyEL4iYwYcz/Jw4AZ1kT
l0qVHdr5OJ9W6QYhI7qsD8ecvlOGpTF2AuLrB7hW6VbiK5GLiDsiiMQtmfirUREu
+Zu+tnPoziaN2IpeWDC9Hszp0+uvwhxsMv4ncwPva35wq/l7Av8559Ng75Zzl/Vs
rqz9p7AhXFqHWN/DdYlxHl0LQZTOoSeRZmM4rEK3Nn2Rd4tOA98ksIvHLtewXh/k
9gy0zWvyejxvlJDWLwj6TMLf7EYzistEYxOYwRCus7ClSGJZ2Q8HZC7WronintoV
bq9K2iHAssAVYfsAbbmyQIpH8o0iYD5tT4REICKpFjTtC8nSr+kNvTrJDC5u9fUB
6shdhGYmcnm4ieonAAWw2gPAgBNqfmEYTtQGKlthMQxqViWfN0krn2nykpNFJjO3
JFiS8rcgrKW94TQC9seGGcR+s2bh17uE1ylXEqAj1UmsIMNEegaFE7INDMj9P5kQ
FvO37UlF3s0L3y4R9RQgFiiY2QAE2yNYt2DXo8FIxQ7F6yPpcib1cbXQ0Heao8/z
aNGjAQBEQ7bO1IV3BLTNKouSmpFXFNI60rPG5yLnezA49loZpR0Oqde7bIk26PR8
4NZZl/ZBVR0r85ZG+y0PiJsLOdCQCK32nU9tj84TZrE3v0kpW7432vZhIsYQW+wY
Z9As3ZfI7tjAPIGBvuuZuj9ciiYqt0JUEzH5HQ45PEHpqpNcCPG0Dk0KmQVo87bZ
IML6bXPA3enLncn/On5RhHWKwmEibUxNiUWPhlCvupR7H3rdSOLe1xRtQCYD/ecO
qxJUVqoMFAnZqvSyBcj5sMUqY/Vf3gColsYapiVWFtRqboPtCb9XWfhtXPMGqr1k
BGnbPOrNUvhvJFB5KdTbvObBs1bHoFnx4JpQfng+wSo3Uz/U2ikc2EHI7Cr8h9JR
yu0NLIMVe+MZ84kfgT4nLVcQRJU/y5FQ7pw5zCPYWh0CcPW1YtCKsHdKwOiGeuaN
v1YYFonfLMGkoMbVbzyXOhqlExd7GhxaJDHo5sLE6ERQJeImVQYatu0sCWdluCDp
oiIw09rQAdE6t4GkbSlZcaVXopSzq+fTty5jJ6cfgmP9XYAjwLkYtk7wjORPy8BH
QljQnmLXNLQXql9D0L1uDKPLUSZy3OkDnQLPWUqkODBu4gBve/8avjgrcFussECb
UGys3t/hnTPNJf9GNxoSLwZgP6BtRtoxfJ7c9YoAE3aNDVE4db4brrKg7cxUGybQ
3AWknz2u4ZX+B8RXHQmTtSrTlfVbU7tfT6nRhVi+qEb5mxavsOGaU7V6Kwv9zwtc
pRVn1iyxHF8La3R8p6j6vTyInWQUTxPLaVPYEJCHy5+jiRFgT+esOH4ZOLmiZICM
oCx1yi25VfU7GGazmIdO4t06X1pVshIcWxsMCelvejiOrwsECMCANptECff9IDjE
E7bjDYeUg/siLyVqZeJgOMsQz3mGUEuOb2FSoTlRUwrHTopMEWqK/kst8JdmbKj5
TVNW7bsSJX4DjR2bymUy8zWG7j0uxtv2s3+xv09YSIMLzGDDTfS7braHxmFe37FO
j15qldO9OuyMnXUwZTSCER49qaZsWEurIUvywLPr57YHQb83gU3L/XDruSfH7j0K
7Ni67cNxldPHMYvS9y9vVG+SiQyxb5TpJuESGLVVFX+laIWMNW+MrlihAHtk1qYi
TVcWApYe5m5ezuhnO7v3CTtkoPOOCXuhUFTlxKitADDhrlwJfDFPPKV06aLAPiTV
4AcxMC1+qeiWuaypameYFUv5vOhSMJ6/0d2Cvvv6dh+ya3IpXTlsuOxfyig/EQxY
vTGVqZZXzH26QELOHoGtKg+6IxdjQfux/4qp2lsOTudiRdHBnVKdNIznBGWrHB5S
QoIEEcVtGSivL2Es/6rIvN3b9hX+4xJdNgkdjDkad0Bgw6YMA4X5YonoAiQkovNb
dT+HxMbXXKdpEiYMzJaTI9eC89RcIFmP3kDb9KH5ISU9x4A1NBhgCg8rqS+Qe+xw
snEClO3MNvzs2UZgyKgtQrvfwmfqSBS8kkhEyQz+ddfJeRwTxty6xmpy8Wm3jjVx
RyZRmjwsoNDf4R+wBoN23WJwwxS0/1eYIOsRa0xgfaxVMnm+EInNwDRthdgnEP9t
wKtWFREByERLOBjqZC0ylcE5C7fXbwEaYfBFJTkqts+8tQ7lqsFHj/M0aSLqFdd6
dyK2AADRyiagLgMnmvggMVX8wUU6XV4yVJx4fPQmw6Orw4zoYqumDJqz5Y4h5zYQ
8R4D2gP96zoWnP+FM/gur2Qy+tWmkuQ0YzZ24FZqH5Cd3cqC210yQxTs/xb7cADP
jqHhQF7o3yta140jr5BH7GZSvyMoj2B9r9BAfzr9/gSFDhBftvxkgHfDOIMddgZQ
uPtUSICplj+jxpebMuw5jZGHn5wGllX5YJvHn9XUfC4V+Tn3Zwij3PTuUEvjVlGY
DOkBrDZdwk6Mk891UhpuIG6NHU8Y1hqCdRYpabAT8R3np+AQrgfNZ7nKVbaP6o3e
5X83n04I/o1FadkU2nF2vxFHJpk4NuZXncbt6VSFih07b9//9aN729+tdkMhXUPm
kjG3fCE2eWH+/RAK7mHJE9HgyBIWkY+TQwpOyCZFKplwZmHH8fMMHUuFlCB4JfA6
nz83hvETOyETPG/dk1k8qfoocuGQ3voKnE7v9h0+k1Rh6A4iMLPkzWfo/4i2G0F7
DyUHtSJ6CzVRB9ccDnYw7vZsod3vpi/lFunrOFZM1PjDKvijc/HhASAHM16kUyxZ
oGYBIYHRVdnljA+J/q87hG/rWuD2FlWE8YQ/AySaIBa0lTFusImmv1zv622XP0tb
HwUMLobAi9eH8Zcz66ZVOc3GKK1o0DY++e1I5cFhNyKQJpb81xE7Xox7r+KxXsh2
QZhVKCASQMJWNmQezIyw+eNpdfQFEno/wH+We4h+yV3aYmwmIg/oY8GImZcPwti9
BqWoR9kGyoVjayewm5WtFaBXcJIxduws9eKme4dKMtzz8KZdQhegZdpMxb6KJOQj
ZcqQtnKQ8kruzSR6toBXsaI/4sK5p7EQYVqF2ZsuIxkAiuH6+uh89129liPv0DNo
y3DqAI3a+VnDiD25fUEQknQP05PKJzbw0JXQCkboqh5Xe0aXIk/QoVoPhoiZyHof
R3nr7/6cwBt5Rx4QOyJvbdzx+ZB0aasDRIAAURSoQi5t0u2rnI5Yi0cTX0uwQJHY
0j5Xx1XO+jHP2Lz2mAk1+7OSElB+NF/A4U9gf4XONa/uMzb/hA1zUFv0BOW+pas7
hd2yWBmWZMpoeLOtiCwVZ36cvqj+48b4KHPURCRF7q6pag4XDMxRjyLHKIUzbeYV
s/X3IIZOm5bVv1LvkmbJkQNt2YwC9Vf5WlqpNg6c3BE6GdXnhNkRanWTd+6HsWQv
Ea40A0V7ERosPyilfpJF8SBG/8GB4kiX0/bXvi7piwCMwmR1TPtyDmOg22lww275
dknqe2jtNr1nOtO8T4hqeKGq/XNtQNenXT5rs+Ho0ZAezJfQRUw/PDz7c4lqczo2
1XMOTsF4dZ1oyPGd5CFF93IAvV0qUCiENwbxjHtBFNWQLL36Unx9GNh4gyk+DlsX
XcH0fFyXowL1Fvdsedwly9GZibhYbN9+lzX8JQaO2Bhc4FICvdyUAnxsx81uk6bl
P0n+XqQEdRsXapwJrthK1RTWZ14r2T94aSaAie9nqeBP05ejjUl7Y/NaJeTJdOqi
2nLIKmZ7PrPgQbPnncPM/qN/y8Gm3k2rdQD9kGnCA5ZFKaeaxwZNt4+Ijl4Me41V
owXRsNAjJUHMaebOqXQirHd2UdsNAEfempeqE63QraXz43IiFyLZTRApBeJGvldl
MBdUELaHf91eAeuJiC2Z9Aloh2uRiYwc5PoMIlQXyaMIoctC6fREbEeUwC7o0knP
sI+9L1lEeQjXW2fVnbU4a5IwLRWpFWGyJKxU+/UwJ2WqJmhutsqZmq8Zp4aytpak
BJRe+1R9uJnKrXBToQXTQGQuynhIdYe+w8buyuOLWVfntv1V5BCY8drU/AATb/dj
LUxXRZAaIZHVE5h3+9gl2t9bZrH3rkgy1uC473dr1kLKLbVjJU9c2dEmltwyXxhk
HP/inKM1Dz2g3SfHso1OC7KOP2lDDILk/vtJVisIkDfxA/S+woAq4uTxaikF0Wuv
Gqrbq+nPgqMgu4gVnT1TsXgmiSyLnfiJw6jKXDtfNROQSKzHMlIzbTcUWYRtoQa+
aKnnwtdbovvsOQGmVnjCsoyasCJmm52fnFyCdOuo0dp7ASsfLKrbwuOJFdEnVjlb
MkYwZkvhFIsuliHFCf1hlqiLKM1M7NkoZ/9U4iy1OiolrSyBz4sFgQfNrmvEL5g8
fKuPtNgSWI6C4kDcDJz2Dz1IvDkRq5RVPqnmnqmbra29OLnKpFtevJihFx6cdbS2
CnHwTVwdaiBw5MDfgClge09/Phge71v4hI7A+S5tS/GF7phxLQq3X2nV4nK3ekdK
wTvFUEteNkheXaea0jr/SNyu0GW6hskYgexcondSPpumPItAhlTXfeiHl7SfjWeA
1eI3ZOOddxxMabH4K9NcsmdO5ud9n96sb22gmZF28ptFLY6glvjF/E3mAvNlyVgV
KduIkteh80GxZnwiNNmEjhpCePC1LgXD1N5r054UbT93RbNxSBU1BLM5SnNs1yvd
SlhcuQQFn0VtCojV0oOCEs6IxiAa1dcGGfWe3ML5PQaawBqISvAsnnyk7AVI85fU
hVesnuh6TBGBM9xmeOnfgMik5e+M+6PWds9lg8gqsn2+hkAOR9SdBkHttCeiGILO
yIbVKRPSCNABTx+iAKmkEoIoSo7DhwHvU4bJ/dok5uVMxODV8PIxmZHqaATZ2npz
mJU0QUF/zvHyt/AkbFLqvT4lu3U+eoOsX9Q70U74hSVNIgIcUBubFqjJ3L56nx7a
9hiizsq1LPuWzPDaZdpQBUVaya46iGQej3CATA/1bC426QB8Njk3xPyVijXTEq8o
pa+BslKg+S15kt1Tdxx0dTOa/JOLwWviOzmI/M1oU8dV+9F+uKcH8FwHgjqCml7r
R1qMgvsiEEEkMmBTUUXdXw3hsTEPdsJNfaKV/XqOO6Be76J2ZKIriGZwAClre04s
rTUf7SJAOEHt8URH/itvrFfJ5hGh9IMp31jCS4jpr9V0oe9G4/eivdkCFP5HUtKn
kRXd2iqADnKP6/d3vQ1VeOK7Mm6CgyNfRH52fUaHkoPLWHvo45hSvBmr9ZHU6Ut2
3H93sNMgojml9qdTgm4hq0Cd18JnKyqobGE+Z656AQMucels3nPa5mGrgUZp7xRO
xJ73VZ8bgpd+PhMsknKVbo9IvQTjgKVDVS4xEmFZOz7mymafhEJxjAwxqxVp9FLu
Fl30hX76cHwJl0evPZcG9iJt3C0MH0wFHovRJF3aeSVUZpg4lCo/bzsrJAbf3BSH
x6OBsDwKaaJcL5lVeDpibVmeB4E9T4/gx6J23dMpnJZhMiVXy4+fmafqV2Fr1VCD
saQ7nawKpMNSZZDHnfS4oWy+BLH2n14n32AsR3y2S+fZWRy1bM5pPrPH/G1cfmFC
bjoskltnevYGVtJZlJyO0a2UXTNJMegAp4FlZKMZjHmC6BwbMfBqabaoyE5Fl8om
mLa3KUbMPERa1K7O0ffSI1VGZwNx7olNoAVF/PP8ETRtQqMwiS73drLGm3AWLk7z
uW0lIMKeMBx5F8q3aVlgzv3/b8WGrJZQwe/FgUGDPt38El+04SRNvAvZfCLcQfJf
VLCZKtRQHVuJxcluS+QfIJefVcBQmwvtsnZ43cixBV41cx5kJG8rf/zcmpT3lKi+
s2RZO0X9hCzRg5t6PnIsuaPZ8dAHY8bjM9XflRiY6R5H9wP7DXVravDtCquXWdts
7ypvb8OUu/rpAQsetLWGGbhjcOXl/QNUlrkF+9PxqyTmBXMpVRgbs82DoQCY5OGs
x/isCDdSA3vthlXYegTzEVJFC8Mo9EGJ4lbXwDlAX2oU7+hLcaflNve0Cxodm7XG
tJCR7K35aIYOZzQ7xMWtkOTcJjERB0i5JY3YPbUT/6IStvB3LMnyP12Jj9OZyIeV
foCSZIY5ieL6n7ChsdgaDZC1lBxTe46NlNdwDO3SFBL0xst2qyohUKmuJ381DIen
hJk7PMTKYT5L5aitV36JOKrr3aDISTqVA7UzxzWnnNi8hkroDmuwq9qIp/d/B6e3
nfKtYd6wMuSlyuISEPe2eJa8cKFBIv9CjImVLaUOJuy1kzM3gv1rc518gQJIXCVi
kbDDxZoT3TjitvRk8au01jwXorufd8U0cyHHGIDcXbK1JvwYQ4JdBYgM+el5MXuS
62uN0TTnfoVTWcN4w8nMd8zsJMmYJfuGNXfItd5AbeJfluHSSrRfil3mRGSrjAux
SPtvQB9xNhxOlY7fGFDZLetfAfQssAVtY91d1CKu+hsKXpFilvAVSvI6C4IA8FqY
LEXfATlyF+Y8azTzfEFcHv6NdHPwFvVfE8pNcKHQpU+HikhvkC/qBD5fjrFY0ber
K3+6Yxw9w58dF9HCG9A89ZQ36aoSX2JBhLgi6IiC9ev94ozpJpx0saIsLLx1FFxG
sLN+YGz1F0pYGHGStUa3eM2m/isPLeAabjGtQOqo222ho7vdUmk3FIu3LVbWYUvS
vYok7EaXVisNELZQ5I7BsiBBkfMWxo92H1f8b467OfVCTpp8WkHrIABN9/Wa5/HZ
uG4tR6pwnnqNNd59h6pWnEOdOy3k8Vlo70FeaPU0SihimhQttWbrrWOXBzn9W4HW
w5au5sbSje8ADYPE8M5/aCrviFMkMbrF0gac6f4NeIh5YCAV4cLfNs+1xgarx5Qj
TM664ViRSrYlwbKyVqzDAZWJTMMEFI6maimSwu0ppsFm4dPlf1qfrqjWy58Sw7jx
45Fq9bDTvIcdN6bIVmhpxQ2r2u/s6tD8+6K2nITotMUvheFywbUNOUyeFCofTxbj
q0e0NuzTwI6LLgR5J1BPEvDx8ELB7sJiTcTaFJWlKgtIQ3XIcZtMNisPfvtEtwEs
njFSSCLJhiI8ShmTkkTOot5Nu0si5sZvAaO1H5IyM/kA8xR7TL1pd5q204fezWD0
R0DcltUmoZmw0HqkbGn4cOuK2yu46MZjCtqjon09nWGUCz5/I6+29QcoZZLOQA6M
f4aHGUmAh7o2qs0Mmz4sMNWMeZLW3q+pWnUzUX0Rp6YaglYzsBY8KruAylhsHXUS
spf0ISN7O7TvkKjO43k4aJIIL11Q5+oLZ0c0FJ5Ibt9CX2pIpqyeH7/BAVMIfwX0
ArJCqy+IXd5+HyW8zl2MdJ/z2vqeOn31VfPUldhLbI1NbQCj1SHzPObXTGALydOZ
EMlCwheM4n2z02IxisPKsBvjZ3/JnsrlOsWBzF577G28qKBqsMtcaLOJq91zi8cA
QZdApNz5pyhCO/TtGp7/TEEOUYJvDEemhm16Q+0dlZSuy2ZSfsl67M6+8whLo0NE
Ey/wxoTuuWLYryIqNWmKBtlCBKDRjmy3ZEkM3UX09Cfo8ixtZeQQymzBHuBP5Tm3
2JMvnvSScy3C1blAw7DDEQGBykRYz1wuqNSmqPIkK1hODwGV4rzlZMHHJ6u1Th2e
n4KhKq6iyvLWxXCilD1mk3LGWNQax0zCEuv1UINevDAmpglxTSFLJ6VIqbfPAGMN
PnTkqOYfcTb1ni4qPA6Q6GJejD27vLoey4rV7BN4fhbDMwWEsFPx6yXPZJtK4FYL
NmV/q8UCs1W1zzugB+gPzxvTSoohFZHdbliMwO8urDAXr0ct8RitK3idYC4EME7k
R1sw2evBAwd8+M4+WKotKGjKEw4zbs1zP5ZA+5vvXcf3KZyc10e4ZjNJnb76eaPq
SjdtSN2mI0dDf8byOP81OnMABN8FaFMvB4IVdN9Zf1VMdLBlZU/o9Q2R5QzZJnMS
AXtUkBakyjDCBw0sJ3e/YTZXe2Fq5Da+oQRULmvVu3yPS5HcxjyCUClz0GDLzckh
f3GI8doOC13ADGmBGEJc03bZ6RM7UTQP4TUM/2jxOL9Do1VZQB7OHjI58AWCmt9e
opQLd3S/Vr3nKvuVxqzPgp2JEHx6s4CPmlqtquKLuWtJdcK/7VG2Gh8hVRKuIEss
D4g18cVM8cTjinJ7BLUh47iwqYZbEgwQiOSfjI2R+R/+0hCApssMUjpH9BsrYynb
K7M4tvxrMWofSmHyYwkmHNm2HTjD6IErGICCwc3bKkz8LDiq/+KO9uhPCj8OWjU1
v+LOo9BErlNtmYo9nAg3H1csrI9mVGBWlYOA9oWW29p9jPE6LELUG0TZy4WOrrHQ
BtG58BMDgO3oU108f4m45pI3vXvDQ2QIql/ooj2yzpjUbDJTHiN9Eb86GGGqW/9r
dw8vQA/XMYsqcEXXTTFoqdzwq0xghZp9rQVI4/ukkBkVtRSqFtDxyk91krDGc2kJ
3qWXEfvsp2nKnkmIx9B57df0gBY0fAgua9MejYcoCtl7vE/sSqlGHO9SVf8/CnWA
/y3Lin6ew5pw9NYjmwCZBvxvEQQjfz2/eWvoxw94F+2+/NvI/IToyRLV4rxowpxo
iJWm0P9hXgtGhqFj2h1SmjRqB/YUUl6pDUoNlrzxL9Xo2Q6K1eejg5cgYj++t0Xx
dK8/vH/jps5vEuAKDPY1DwC/pU7E4M8dztIsdKcfcBAz9NzJA9ZMulP3/5oOMfED
u0KPAuQtEZSqQM7QVXWcr7IiHNXZZ43Gsf9EKfrU8h8iTBms73uOPUlz8BzvTVjW
LipaAvlzZUim0GACYX+H2JDen+Mam2dRZSYsliv9fuf4uV4tHtKHcBeks6uOuN7J
k8OU6q0LPNgKMVEcjLdRccqCzPFPmA40U32xf6pbWC5Xs8bCczCfDHnIErOhaKgR
xAjOWsBoZh8D3q+m+ely+EJMfEPGDtDnUMGs4XsLYF4gzm+OFK2VaW9mzuqNcff0
/nfitVuF6YJU4zH+18jSv93Tn03delbMHPjUEbrfKsvuejlf9wYv138eRoD1RrY7
lNTXljrI/1e6uauugAaqaAx5LqC03DQsFnb1nH20wbkSiAY1kW9VxqqYTCL8e3FK
zrzjXFCmPSTQJhpBakpYiQrzQpoVzQo55oIvADcoBpwYalKXOKHw0plNBZFGbTd9
inRnfvn2zvXtJ0GFydozkyVxeLDxN2SRuPPtpW5poEahzAnsCW2n8bYY0UBZdQ+S
sUP72VBsJhNk7Ufe/UjQA02xfAXm3lSe74+V9NdHOzQBONTwDXBAAtfVc6M3XWMP
umERs631UvXIb7JJg587Hd7ZRZnFb0dLb5jK1Bi9azsTdZeio0p/3fj1eOha2hiE
4b6Df8bBDKUnLtYdVd/7z7pCY/L7hcfVlwzb84TBeQ4CWNum981NfqA4N/0TxWe2
BF/8w1APFOopv84GqxVZOHrMP7Ni3RTyeg2xzccrpk2e96k7z5daU8Ihnayn41F2
cYO48TbDmvQ5W1/g0/idevdq7SxCyoJ5cZS5JYsF8GiIKLJeBxaGJp3NG7TiX7+b
kqYoaZBkkbKeyp0HSCx18D9ApuOiFuzPz4w9ZyA2P2DFxP4c879AHMcRa6v+Suz0
h9tMvDCM/7UiynFNEoVO/NE9ptim0WwT1c0DHRh3dMGiUS3qIel5NAi1TnAotIHS
3UI4jkWunxqXWg+h+AxbJvFXojbW9XroUtnB+/C2Cr24LfIm4m5Ffti4D+04ZDkS
aGFGnS4+0l2+Wa+iJ7pRFGyHli/ppB+UmEYPc/v2W/NOxiGpqYmq1YVP3ztX0Vbj
VcREPTh+pZCJE6GN0kmijVZLRgUnCFVxhYGhTJN7dS6YJ7Il9qLBFCD/5PQQnxoi
EB7p7wMbvwvH8KsTud4iLR/3u1hNfr3tr7ekj9HGwfwgpyIgCBHwQolRlR064ddX
ZgJinohWuL4bfbJ+0CQctk+LPl2dK91f37SpoSNo9Val17eU9KVWj+CrSZOM+igv
ALH9ulQlFRNmD4eU7Rs3RNc1dbAr2Tz7x6HJtXE6l7RItOTD6QUnebFcC99KZjTp
MP6gDTHbu8Al5fCMUfEr6nkzrvdJTgy9/SXUfrZavPSLGEuYcYJL2rR7bBUNPN45
OC2QEqzVx+Lqhqvx309UxjbK8EFFyz4QSguTuSwod8SWwmdVHKnZ2gcmjMq3E/lD
6UnDPus9rQtYh4s90LzskLvGikFt9bZKkFIrpg/9fprI/NgeUphNN8loy3BYqdMn
dJ/UU1Pc+uYCkrBBUKyeQ4M5t9NQ73V8hJH1tIkrX0nLpM76qxxBcipV3pqe6sOC
IO9GT9vdg3Uhml6vNs0jrUeeMrakPt/dWvtxGWnCojoB54E5pySNdKrnPobKqZPZ
+VPw8SDhJg1HJU2g29WKMo7CMdJLU2d02MpXjj2PA34FJ8/ncF0i8MbAvqmcqU9c
ODuJ7QGVGg5ovzGt0gE0xjzm95c9Vdm+T46COyRp/CuH0DsGNheBjWCsfbygC4P0
Nz5MC2Z5Tq9uKwL3aLEPCzGaxOr43QhnJb31ZtqrvqC6dSBiiUhOA6cSRkFA7Soq
44U6JShiNFoHsipmjyw8bGDu8jJHvkllDxiCTNE6jSd5ABjrQ8cJNnxjw4f4nQKN
zHCLOJV/Iz0q00xTd+NTD+DcIZpw8WNoPiBkgWMg2d7RqAPj+7Tq2MSzbn9NvFzh
WB6DUCVnK7eXl9xXz49c+3KjhePwC0Vl6Sx8kN6MyfjjCdWNOYaLcXmBgRnjB6g3
VqzofcexKl4rRFzJr/JYU21yMkGKJ3+FevCqVaile6MDAFnLnn255eSSapOf1Lqj
8xVtM1uMVMXHY0QLOpRGUgJa+CKV6SKKZKZOdNfXdnbiI0URD7xscQoe8f5ObBtd
JcFkJn7vb1tzgROlT9xxn+8lLI6nB0xghOqvWEuMW9vaXqVY4oO+PtJ72KhC/g3Z
74oVTShkof0yvDRw5SC0wZ2d6Fp/815CllmHCeJhaFngfQzwz6PemMOgqnVMeAQc
xFvZ9uB76PBT5q9M/QfQpT+unYjE198356664b+i9+jdxBQgf1Uv93sK1ODgs8AV
ng+eicZ/aCahUqTr4ZELnYUPcl3RvFrOi9KN2hH/jZN9rool78hKmgIny6F6Q0Vw
54JoyFT8vp7SZW3vr8BIcP+LyT3XmBdKgN9EBIyDv77n+BDPNWiZVeY9HWGNnwQp
Mmoj8x7StuU63QCF8qxdwea6UORzJJ5SvcHvgmUMSiMmPX5VyAZP+cbuEZ7V7xR0
l/Vw8o5fvtt2nKj9my8f/qCquXmA58eTBEvpN0s4Ljy4Z6BwICqQSNygP1NKqdwm
ysOvWQFQf/8LjwrXRylI7w/3vj3Swg9uSq9Y6S1gbL9wTR+U5Lh2g2AmTFlojIu7
EwF6lEqmeJVu1PMfI6zwO3VOduQkfGSsryfQgdY46lnL3VvL6kRl1YiYjX1Z9it7
7TLWbo/9fTPdJ15vB02RqlvsNiaqSNdOpc2k2I7IvmEc6M7UaI3kNSOH7yhpSqJU
8DCeVZF1+pOJMq6W6f+jJTf2ghKjZjdmZhO0nKWxC4xKqIMaZzcbShG1Xl5NGECU
UPVmK8ZyiqnOeKZztQNzuwIPmdXX2sAyJhYLIeUKgojXhL0oMKv0Np1g6xToVwIS
UgsNVDuRHEOpQNhBnhSjCbw+tmKu3oNkFCKzEmav8KhzCA8WfDFRfHqW31TX8mJd
cxzukyHHkhv9CWcesqybkYJx/2EAt/7rhXmeMUHUMAM/zDcG37MjO/Zx+uqDa958
/QGg9rZT7W7o9Pt05v1zo60Dca7v+Bwwlmi7WjT+Vk1Xz5dUnWBx2TIncAgWnbRH
bkEuY+SwNkM23BTUb1Bgj0KtMLHAdJUV077JV4mAtIW25gIXN33O/gCLwROBqMtJ
kvbTQwq67MOFH4t3tmur/Wy/rOUVWErmwuGmQnb3VfbmoUKQsPVPY9eN+muK+GLh
CMicnEd77xdUjiVkLs+UPd1/jiS2B9EPYmSkmNZqoJo+b5VpEMVcXZgsHQ3Gkgb7
6XPqaRWSi0mg1JHj52A1VHl1sO+99HAPXUKJLhDUKHKaULaaPfu9HmH4opWCmpvf
qiId3gh9ajo2VNROnoXpbQUJaBTX2IqNNrjOfbXE5FAaTX4G3WM0nWY7+xdbeTHX
wjzYhyz+zPEHklUA1vACA68opqZxn+fmLhwQLSWym5db6EqK1jeouNEdyATOzr2J
E3uWDVC+PeskxYjtgg3bYq2FSXPzUYg1EzjuVQffUYR45ujY41o54xn3D3X5rlC7
8w0xJPiihL4cSNw0Cl4x6cdCOAOQDWqRK1YyVCb8iaNVonvR9h52AmLrOvrSIGAa
Ln04rTQ80UDHz4NlM4VEIs3IRnc4MPBgSBNIfOdA0cItNQwSsGIGiMLjqu3rwBnc
Rrcv0T3VjQBOGubfsuRykRs/yjouhS7u+Mhm/XR+prdelg3G9X8MrwmpzgNeFAd4
Q2TyziZNRd+MLNgP00GkKKxmGUH1pqfw1ib8WizxrAkyPQk7zaRuTOgyXqxEvDLj
4w/lKZGfl7vpCEjW1+Osw8r5Nzl4pz3IJL8UdO//qN0nvdvy9UEBGnFdcZwIxSjo
T9zBCgCfQHGn2Mk3Jvz4q2M2kDrRS2hXrwKR7pyHFdG7ZNVFo62D02o5/GVWjJZi
a53vkpNDKTx7ZifbVMCiShZLfpSs/Bq6QHykHvix5pvcPDIsj8D2MoBzOFoj8hAR
sNh5akj05sNNi/Gb9yDiHusOejdvLHDaXBiBKpU02tt/Ws794FnHsGg1jBRRVDcU
kzMIyO0PtZFi1Icl9sy2IwuVie7EEbLZsDOsqutUmAK37qoWc9UL40yCPg/nhanD
lV1sf01lLqtFTXCLzluVBQohXRCthI/lKP7i0DNg+9VSxiQgEnBhMIqOgV7yc5xj
N8Lk3US9ZlVZY43E5U9ZQgnAnTIyZUh0CuNQOperroCqrGQCda88QE8wjvgMTbFy
CIaRP6CFNYMWyMRUEqM1bE98okO8wzWJzh5XK4fZExL0O8ex0bK0Eq7Xs+FAhCpj
IxfHY2cBzeI1CGqY+6Gqw96au7uVNnqyE4wE7ieBYMGVtw9vq9fbHQTfyZZehNBJ
PGC7vvcRpVGC3N8zLoiGa499vdIKYruzZ5fMciFZpnc9qM2TQ/aWA+eJ2DrEPtOg
Vm9xafeMXhmY5eE/Bp84pTIbEOGBmLoFNIY/rUP2j/e4XTcor0eeYn0aBlW+MJlN
OLNqmVrnZkE+IfxHfw7k5NSI3lK0/xlDdX76q9ixIXVCbuPB0mJ/yE+LwoZ/qSK2
y9TGCGI8hYRXC9kEsiTbzm381HXd+IhIppHIucHPe1SemD2G+enoV0Rb5NhgUumG
vb42Mg9m8XnIVVZzY0Br3DOR1/WXWdLLBWDyK/8cwNbJe9XtNtP/fKY3u1h7eelh
qFpqoI33ftKFvdPjmC6X99V913QqtJ0/ZEQ/XnzFqAMR0R6LDg0GJyRo5GgL2a+6
WfEt3s6CMutsnyqAMoIJ8CFACpuUZoR5htsJNUHmc7QzJTd1pve6yULGsryTtdtj
o247Y7ENAYJ+wSfL1mDfQcLhNRi4Sp3adnlOXtRzz0qDRva1zo3QIwVC29M726eo
CCLRjUY8E3DOHFwri2gPuyDL2YTMHCm9rZ7tIqHDw/xFtBJUhbgqi7q2bkYSiOhr
6T9nNtOtGWcyVgAheTe+6OsUx99+YhsEGvlBlv8tcTKT/Mv5l5ajSvwotDxY/xqj
p6925C3/oooP5myCAQ+aNb7dh6Mb0Y35YiSB60CWILH0dEnSMJVFOEHxgMryJ6H+
F3TRKZ5amrnt3Yez1nISp1KNbitmnpK6EsmZqwyv9LMV6xgwHLHi18Qa5eCgjYvQ
pzPPqJNIcqPLiAQG3OwWcEHfM4x0ZQag34wmmzhz+uFCWgMBxX7oUm8KdQQsRMPl
+ae44kd/bEVPU+8vYleKF7XZHGNBIsYB82EG4FO6f2TK82FrVLEWZ7/KGiIS8bzb
hdDR/nIdqMhFy6VNOtdPzbuPYKlesLKHQdDVeNlCVAQRJgHFIi10O9aNL9GG1FaL
7Au3l4m3oNHTFmd6w6THWbzoQC37QoGle2SHJxBq4LfEo8z/TbKL51V9rG44rOvo
MM8ACTI2FI9WeidnH9VmQGjGrVNEZvceAK8sUIRqcfw0sHLbIh1L2c6H8j4OFtSo
DqFjQXiXmlie+62GAxdsxl52m24Stkeghz4B3wtfvc1kN05OgReAjsEcV85lzYHe
adEs694gjf/0fvO2FFdoUZWNStZM2vsjwg6NOVZOyP4TPLoxFjzEBN90ghK/m3D7
SNKJ/SHwxFFILo8Xhp++hdbGAAxjRuSOfykDtE0tjhMfX2jaZZadgTFXilA/kB8K
xK2jyICH369KDWmjuD76fPDmo8G4SqYNuWOwDD3uvZUOdqhw/n5GcNGGmwvm7g0X
hescIMYvZrSfmPMDKcmC2G/DAReNWFhEWHsSF+tG1YGgOMmnL+g8KnuvHSF7jk4t
W3q7gD2ST6sSZua/NdLmo5x7kgkJLHpkNbj5hSqBi6GxFyBfQc9AlIyW2uo5JGIQ
5uLoKUaQwVto7ImtjXoxpHrMkK4aBsqy9iw9KkRBalmM9/1lsQAXlrjufOCN08ZO
MNNWAQPrFPYYUu8j2VEpynZ9blBWhbHFaMLh01011mOhD8+CE004l77K/QCe7xzV
Gzg3wl/mpuo6hKwJn5TDZq7qh+wkRsQbXFbYNOaUgR08vod/sQ3BowH+ugFwbJ86
L+AQ0a/sIdZkDMHZpi7bHCG9xb8RPTZR6+QC1ZHgbdNE/rXb/i3gAHqnFQAMLs/s
UrpnaUOklcjlyeQIGdLOoRyfxEfPIpLyRUQKIHhwdzs4RX+JzOKKOgb+APILAIqO
164v2clup0wtHm4JIPd25kIuN6BiAYP+DIS2eAcHq/DU/NMy3XloNTxs4XrN0SRg
9c+hTjwJk2jZ+vsd2RQeC7BbRzbRZkL4wnlIYn++64eQXyCFbhAsrgtbvW1pZ/iX
OdsUcNxWkbIKy2k7rKLcAjDcCyfzW8PT/Mcf7AaYXyk/yUa6SzgN9fAlMZgzEFTq
Cq2HRy7fZsM8rm1dn5yb2wooKDmrt7/G9QEgwkzrHFF31ztly/eq/oAls6sKa5HT
ciVP/cX11z8WJh8cRLiUWSIBbeBR5UQ/I3uxV5L7OYLX4gMHd0FSavOIUpXnYsuS
vR59/d7afYCbWPZuR3nyWXM6prNazhE+fv3ZZancOCTPYi+s3kmSTlOK0wNDJbOC
WhNmea9EawStCi8ll7Wyu++dZG0h8JqH2wJJmaKwv1grX7jF2It7o/7a2ELPqX4R
aw6jWVRSqzCcYm817DOStnEg6J1hKAVqy8n9FN0N/LLWXghyv6JVlHJsei5pQX3d
/ulQOE6RwJbi6wMSgXygggZ6u6QEpRnOL47ZdJ3224/wCkVJ7fX8sdZrV6jgGizg
H7z+Ulh1RUP70qM1kgjtUDXPcDi1d/q06NnhE8161LzULfqi0mad53E4DdNV7Msi
idVPZ92H5r3h6D9PEqI6eJsIT38gZK522JAGgNk6BKqSV+urscoMNd2Si0dXYsfo
F5znKMJN9RY7YncLIKXBoziDdttpDapsh4n1cD2fN/bVQ15Sue7yUN3orOb3pFcw
367CddXg/MwfsphFY6x8YyGdg6vDnxlSfihW5nU34mjPyz1NUYGkbNFFX5ws0Biu
NF+ZdxWs2ojGbaHXtJMLsPDGE8YFyjvBw0XpexOKPAdT+8LvTTxmQa6NsSs8bKax
3un6m2m9SdFPFzCjLnoDOZSJjgiWfNF2xKITKbViei41SL0/rFnEQ7tNAph7kavW
VVqIN6S/BmVLjkSj2wX0BOMT0xX8w6Y8VGFR1oWnK8KF8nHowUAp42VfllMp9xmA
miN+l0V/jtNnmlG52VZ+AodF6UCuLlCIHMuCzi3ZY+nLTlHiNKbKBWwm8gDd0fq0
5dlbRkvhrnwPGUa0D8DSlI0wGNFJtGhS1dtgZSirEQWZmwyQxMRUS+wWVstjaoja
fH9EIdfEulj8qw6JzVIpxMXL4E9TG45P1eOzBaf3jt38jppB6XzFHcMPMgXRBgo+
G9U3HNw0Q2qPIsRoxATfQw8hTyloO+EHSLMQppyncAfDdXbbXTSqM3GwzGQOfPxH
vpIx9N/EjPoQZpeOJv6uUcTwvKXRoWbD7pVRLDAX5GDO38k08BQ+85u+YHFBHSaw
mMupeuZp+V+F4tfJah+ULoNk/YjI2H3W50sXbPc0gMrK0UDnWRXH/iXsUeo6zxOx
unLrhLxb+Hc3ZOPWcgtI4P2YHC+tKw2YW/WdGFyVcQ/0BOQPjpE5y3JHTqeZVsUd
VuVTG2+t/VitlNLXyF3t8ZMBMxAe/kD0PGq8xWhc6wJ/KwHNX8rD36SoKMv7FCgU
+VdBiSiOG2xIzXfdwK/MUQSu4aSDjrGpQ6pLEVHa3XAEX8l0IM8UkhGFJe+KFeXX
j36Ya/8OYwCd/m2/rXLmeLGhY4o7szkV9XlNmpzi+BLnNgLUH+JWCVWoxenMGFQo
Y2pGVRQzQkLr68sxI1SBTGulaHihevCUsgXXVN/Q9nMBNIztCE7WHedV90CUqdQc
8XXm63/N0U4i6x9qe34MbyS5VcOiDIesygzyP+IQ1dKHstONKEPo0lb+XWJfqvA7
QmOY9YzRQN0DqPpYG5FOti5tY4SnqQJlbYA6+xzk8COkwRidfUX3KOOiQlvAxxIg
CvkGFr1ss2A7NIg16O94nFHzGIi874v+tbqJjk0T1C4ZwouMtXwGKXDyBVTS+LMm
3vCvC5yegpqIr05pdsh40G4PfJ9KR0tF/m4hWaICKhK58+nCgaORMcQEmNKUI08S
rHM6v0fdZmCcb9UHulnV8ytz+wLrlHsHpZ8QOPSNgORue5RxyHpcEZhrtMdjxHLP
vBfXIKtQx0iIRg0jeZ27anSDYP8tkjBMNkHMxGvuz+ZNZF9GMTpPHK8q17895wMm
zohrUM/Qsk+0QHoupKhBcEQUiqN07NAjo98UA3ghPSBrX8YcJiXvwFm9hMPJfOpF
7tIUrXvyJ6mc/g7S3Pcom1FolDPaIlz1Xq5O+Hh/vk+VillyY5ZX66cwR4BMRfKH
Iyh0CE47mF+XFaLPRlprVEsRCk3DiJVOImWC7Vr9bVuWioot9KcFuOSO2aigzWim
nFhK9l0yFh3MAtuOGB+xJTwpK74TcIoWi8c3EH81hVzb1dB4ysoj+np7cvK0Blji
XgzgqaDn7t8C3nd2so6ba3p8OMCmeQEFW+R1wL4IrkSz7MUC/k9Dn4Fah1eFKAaw
2TstQJaOADasZ7Tc2yCscip02AGWq5I8P62aKUHM5L1qa/2gMiuwJopPSrkhxG4f
DQE9BAS6Dj1WfwPVb5KOFT2GOrIqRGRTrvRe0OKJkJJdoT2ZG1DnlmchMHSm/9A0
6OOM8pvjykCj+rvFtvbUGkC0BdGR/eB8/erX9ntr/zfkWBUviZxk0NRNnZnEWas4
WolY2vO1aSoxQ7lHs4zARY9BtNavbn5SJxKbEo3A7KRY/ISpHPND9+sRi7bjXE7w
jrC456IyjlRwzyBPUgQX2em78v71YdUglwMjTV4J7UUi9UDTObvpKa1zaE5FCzNo
OGZBfCdDXktXZOHVEN0yrHN5Fx16005lp6e8SiUTrOSRftTFT9nKvRdtzJnNTFBE
XTmjCYhDdOfEmLq3PBB2lDFgDhK79Qmk0GI3QY7SzCgquhCxCkuoHRekM3O9U/uT
//XwRf1xB/qg893riljZJID8+eFlwO8Mn3TxfoVRX3j+k6D+i3TfC3sXasJAHHxX
0DcrooA2Q5b3GZ61Ie2Nyo7EBKKVDxjdOuVDbu5LyohYy5oftldJJNrzssPMKLRo
n4poWAlqZhgYm6DMq7ZiYgjykLTdTBSc/zbnn0dNMJFnkEjZBEOH72P9KsEQKPAd
CFJE5H5ZO6vi3eJXxwJbgdjR1u3vq7OKw5ZbS30SF6xkPPdPMbwJE1iJa9dChtf1
QvyLHnth+A+JlgeXToNWCFmTUF2ZM2I6Q/unwBxmnOJARKid3pekoglsSwALQOtV
8YfBaavBLDJZRlq+06oiRTC7gn9q6skbckbIcMut83OJNfroMqv78tYMd0/M5YI+
jn2fY+BUjfw00jz6yHl1KamwauqYfcGUU7DUZCL0KXCxpl2WNdQSwj2+Rlp5UXJj
i4uojDNDx0uYnYNk5Oa25jv9EgR71b/69BGa6is5UsVmG8sDx1Xmoy3d8jFqWj8w
Cu1zySWZDE+L0ELIVJif2/chiAanJY6IInqGM9wcHI7JfSFggG7iD2ZdNf8Spkzy
OpnIjpCzkxMlp6cuExPzJyNhAxiHydsVqmXVTf+R6w7uND97LJTggd2EC8m987WQ
1VlM7Jp27YOuzBkdqTo5xKAFmbUew1eu02rddi+hUkdv7SjjTT7HkyYXm1F+/SR8
rEbAqQpjvyJJT4fPwvA9zPHylnQKIF2nMGacgKAN3p8/z/kGyZ6SbHsVe4HpSKvu
f/RKQ+L+oVK/nJo7uecXKfzLEQGG8Doeu2gtbebaSCOrwkkQSyu7G68wucV7p0Xe
7X/3DIO7qsf5fzXt/yjnUTE3R/GazAI78+SZHcq52SXbUddTAowkCUhexxOv3dfV
YLdwj3FCx34UdsKZPUQkIKll80o4GDccphbg0gmeODkgHpRntGoafl0t2nGemznN
MFWmp2mjieih1oFmGgjBFJAnFBrcvI+UQcVk3Qk5BJVWmRdfXkXBuCIlJCt4/Cqp
6bfcCtwGp5hwG12TwlAc5fwDP5n41T7aE5bUJFzHeU1Q6EK9/iVwO/THwqQ3Jlos
WCU4p54pSH+Lg35f2mVS5mDROJzM3z4gaFFRyv8zyzk7RODMrTPRCGajK1OsS6TQ
RP8MyXUFJxhfLm+98IX7mCvhLrZy6B8aldmXcrYDSsOg4WLGbRQnDmwPz71ogiVm
eWVmDmfnsmeEJRIyrD3Grp1/4Wkln5B9+NQzzOyii+BIBgEtsgn3cRqkkyrvac+Q
cAuoFhFyYUCPgz4I1pBaLc3VWqusCvIpcrWkb721Ef31aCilOc9wriPCPFe7dz2P
z7PaMZNsuOFpZ77tSE+zvAoWYLxhA/SdOh8LlG6Oz3n5EeV3w9/mkYHxzr5AjF0r
OejSMQVq1y349jLEo1T5U0endKl+FzaSeY+flC1tQLwEXVvzqaZ2Oh3aJDf6AgTV
lhMBCpkYWMKhI1e87+7YJcKwiLEOqKqz4TVAii5CWmsoorP/G+8+0hNkpVsFsf4V
FCgk3J99lGEfg/lsRN2W+z54+/ZgRci+0iwxikIBPRCI/RcLNoFKKfVhVezGBy68
02cM1c8uTWZLECYEjfM/Y9+6QVxYlxVVM+2clOS6HnQOZi9u88TYxRbwM2TKg9KN
OAzhUgL/m7D2cA4Vp4IiKSz4e9x+wVM9tSjv4Prtg21e0OMUxctyNTNvgVVP6KzR
sYHkYie8mwQ26eOVP6L3pEA8WyVIhrR/zqQ8tdjOwfNMzWQa4NjS3LpPAlbPgs2a
vU2rjOFiglCSlLGhG8CiLlu9z9gxSclqIOipX4avUaT2UYjzT15bQwawtpCECwS+
2oGgp4jSEGaxdRjXrpDXw6WN7aBAFkv4vz9J2U3ySyFtgJDwTlCWjwUttao9rXff
B9nUmR3ztOWlLEuL6FL8qbBUXaIlEsnSxOdLSENiTH4IX+46raMOXwSuUgSbD47G
+y7qfMqzKpAPz4jRp0970rJD09quQZrmlWvN0qIP83I7M/Lxkpb0WXvjl8e0lY7b
WJJWrBLFRDOk29wCGKFi0aOFdiqeV6k/UkWqUn70BTdvaMVEJ39VeIQQZzmg8fmN
EDHb1eebyNAswIwd6KDfFEgaK61SsBFGFWLdCM5KbAgtElKKWKMqY/zzEcYInyx5
8dj5mA8VEutT3h6bWh9Wsu7yd3HPCifDgJ393Y+6e5icJhdkRfeGNWDfEi1fdcS3
NPLuY13uLyr9qwES289+mbROUVwMcytsou06vLcavvw7sZypkoamnxI4JZnHsSiK
M2wQ2aOS3fDtz/wEzLt0K5k1aiSo5SzB23BCs7ACJNU6N+XT1FHmT0uIxT3Exphx
rBZC3w/8hyTAWG01QxSemY6RO4a0MkKkLHeSvgL48b+Ol3RkiUKSbaq8XRLo/h8d
I7dVV2yvPJN67oSWCrEb1ReXJwK+DYoVTgWC5fFQbN1HfYH/iN3UZpp68ETQQ79O
RqXHlfBZjZBKqUc1KOmVHhqH5Mxu1LZ3SqslHh3yMOqo4Rr/NAhmjF/neGx5NonZ
zDcipVfZVl/54sC3nlz+R2diuM0no3DsjE+PmIZnG+1oHr1h9uu2i1IY3k8oMGKc
zZnA/aIHfOYFQm37sdICKnNEAVnltPWF2rnHlQd1JDRL4Q7q0qdie6jgK7JUwCaJ
qLnmTGbwG5bdSCgDz6T9aRwTVN5VdlTyM1c6g7N50CwMiX2WOeATefzCpuaiF2yj
N+dJ0NxQJ8fFfdC5K3wPj7W1okQzi3k+0lAWLQtirHDRLOXcZWNcCSVSSKxONa7f
qpii1KowVxnI8y2Aq/3IwA3cICrZXRxWifeC5maD0mNO2YDGjaIWhA9YafEu6abq
sL9Z8pP3bYdTJgfph5yVAUDq4APd/6DJh416NzRKh81yicuFxASFdwNBMAoAjX3P
4Ri1zVO6DCbowbJKUFbCOpaggU4BgDmH/L56vYZ7Hcn1Buy5B0SMuwdDLLIkE2Fs
JQ5hHinCiJOVXhO6g2nKfLRb5tk7/DagLi3a8OVtVWO72PoHMrM4RY9TKqJevRS0
dEpPn1SDIJcyQMrbVvEifDewTuCAnRKQOyXDrjkvku8I1MQImh6AwzvmilCxxBPD
q5yrrzIe1f3BXaEc6cotM011OochBpnNB1CWcDdK4mMdKkGQIJZeGaotzzkwsNls
W3K6SVq6LlN2D8pmKiJfUNZqFJ5bizgYn1V9DswINVlooeQImlVmB538o2YBMVUX
okol1py4kdvJyPcZ/BVEiUXyQRB4utjs2TVWsT5wN0HbSCjJgZ2XB5DJEHCUacRa
coXy0Flz/8jdvKnFAGmpN2462yT0WwD+hPnfc6lyjsky3He+i3wu2wWZkXhh7193
GM7uP2ha8Bt4okO8O2ORg6zxSr/Dcsdg2XWCiJAIwojpe+j81oItUn5hAD74m+yK
7nL6X6VbQB4QK3BZNBpu9FTntW3MLE7L06t46PyZ2T22RRaD5U3rdbFXpT1iCsiN
YLJ6QRGMcB60+xfdJE6aV7TxMWEBeEP9jVii7EhBfhZRhY19+3wj8BZ0iaTkIN1Z
bq3r/V0hgSOVo/mUSM+wnTZRfVGykvDTKUfohp00HJalsjVQlV1L9JuIXZNPwMfT
BHnonDq0sDl+CHq9eke/bFjFDKHSLPO9NnR+1MalEaHzJYoQYxKUbozhJvMu+OfD
5QVOF4n7gGkVS40WyCxJj8IInIVR8moryjZ7L/TRdFAqlB/KMjwFkIrfDw1N03K6
Sse03R1eEyNf1hqJfTA5CamuuWG2PrghHeW+8iZpesrSjEe+T6IHqppr/i9mvJnL
a5d1bAgZcPRxOBnb+dJag0ge+7l+erQNB/qMjriDKBF92ql5eAJd/qyCw5Ul7POr
/RfFYWpcLAgM2NXbvhY5IhxP/dn+mbUmJnIA4ACzctStB/vlUtBzrIqHF2XRv1vy
FE4l1kTG78+v1/szvoPs3pfUElK7IGzI2pJ5Vog6rMMsPPMJIkW4wG11b4TRTPpQ
iSWC1lCmm4B1h9OzW3CIQ08+dMqK5Sj6+8z+Jg/PqJz+QSxC7KGhVqWUxkKAkNoV
mMRbnenbQsI7q6s4xZRzSwaNuRdYS/2GqlH+p58AXJYgQyvG5r4QXHO54ci0SZ37
EnfIPnnZNVXegfGvbPLpxWnwJz8skPK0Q1fWXS3aZPRcF2fnrZTXsxeIYYbH7sjY
PLGw+34f8FqfTFR9sRsLghYMG++F2DW1L8vo5BC5FhZQ6vXRW+lV3/aLbBhH+vqs
WvZQCG9VoSinsYmlOP97j82yT2rKAq/d/yUjULYSTcLYldO9aLSMVOxLy3u9uCEZ
aFA2bqyhntVmlx9QYCSZN1HU+2HTO+FExPz3VPnjyvL435MtDXv3PFeI87nXdA3e
qLP5XSQo6vc6Rm0aebUzf7W3txN7VgwoUX62A76+wWgc3hCc6eTd5NcNIgKvDk2j
nBCRsnHemNFcMzWDt6FeqEspY1uqisszLa+BmuzgwzrvsD5yiq4z39fpcIFFmDKS
QiB1XCVrVtWmtJNjxZLSr4vO4soUS2f9KXH3uIB8vMT8rFcGAkDUPhZODHINqPAu
O5BNHDU+r8NYpG6NBHLVfudcfjag3iz913g/f1AFFh3kgY6C78Kt3hAvgqZMG3oC
dDtbcu3wKjdXv0fIWo7apPeEy+81PdvnXXBLruBTwqMjERD7r6L0Ht2V8HBpcP5y
R/vfIJ8zsneBc1RBjwN2u/rTki0YhKnPcaOMsgbgYmnF4Ej/JsSuFNArMpLitOX3
gU3fwUy6766eQOatGLNsGQ8NhLyDL6Ia/I1v0xXqiY85eKQ67SB9GYuOwdl0Cp1v
FNXwjGjM3nS5tPgAwsZ4Fon6wKFM7Hp79mm/vRKNAgiwSfFfnpMG//XcyMnNNro0
GsZItH1itXmlgz+jWT+6R1GqQwj7X4tnJWwodbsmy7/od0y6O7i2J/70KtYhWyFN
6B67+woITFg8klwfEwZZ2YYrcx3wbaDhRzPOTvJb1B/72YUGFBkk0mskF6FvjMNw
47MbO+xfWYGDN/yFwqtokCI51Kga1nw1oNyQcPHvTpvvPAHINrMBxpMzjvRU0EZk
XiUAM622kNGA/e8FZclp/2pgDYssWBOAUgwivxjUCVN4vJQzI+jFQfFcARUjVKYh
a6OYY1elcX5TxuLBMp4y5sbMMYba5cT9NCSKouQQZcgB95y6S78/3FDZf7Sra2ea
XvapdIyOaIrobO7kU9xolRVqSpmA8lvzpMdykwJELnTVWBcd1DgjjGrYpRo1G2Hc
Wol2m+pATUf66b3B3G0Wf19m3UJ71beBQeiLw8X/BOzfnfI+DRhehyl02/x/DEwt
vT8KtRijKQzGnb0blDeZoko4IENQzjzMuQqKmRFcNZPE3WclcUQrUdCM0lbSp1YX
XwxZZhXNcDvB0TAlMjAA97zUDwiM3/uUlUK/RlHectu6/xgM9DRARo7I9bhiloTd
yPu0i9OjHXimZy+Iz7MAaY/otFYW0Mt4KIvYzRhis3iM0fiNBiKMJVi9mIbh1tLW
LYe75C6q0agWxI4v9rYYVJAo7t6fzRlGMkIO2F80E3wm4oBv7dLof4tkcvwRM6t9
CHQRRm3DhQYkA5rmXIviAy/UT9/jfjBuSWYj6xxw9G64yBvJilk13zPJuCiejzZ1
WjH+7JpCmAEpoldb6c8GsTDDXdB6WyOvuXir975iO54ldOy4we5suBfGDtcpdm9I
eSqeay2VTEfJQL9Mj0CUgVdtnAbu/F0zSmf80+N4sZrieRDaAzf+Ivbaawuyn4Yr
IixLan2srMtPC/55IZN/Tx8pi5Z3XTMAM6NNf5bVPGe6M45KAdRpKxtySQdIVuKB
iUN7hH9ZarFv4cg2EU1plaTpOLGnkUpOPHfeT+9IHq1S3Tmss0npEgQWwlTY89LK
4tkCJLlQrYHHzrDJV9G08s/yGxX/Ga2rJQXOVmX1yrimFSFLEUeD53zePaXRw2LK
MvVf7m3Rb3KVEPpZbd3YZqIVmAim4c8a7LgJ8nfQIYtSBCrwzpxSSzGYyDVyOdTp
cB1Ir1vIzp6fVDW57TAq8EcWTL/4NU6JnuCfilMH4CEa3gKLWVjc9aABFxWJwwmA
z15+ByG15YcT2kojJ67ZzskkEJis9yOzkz6oX9jgIfQenY7rx+VZcxk4h+7DteuJ
DJtsN54deMJMbrpE/cjIdc0OdrQMH/1+mCcc+k4rLON+NzSmdwjuoOYFSyTikoiO
h2A0gqNKMEmg0QmmlOk9xDXlODVol48fiaOYgGxGwztgSTGWxCjEiA7GwHKJXnt9
BrZcc7qqL0flUZYqwt+zu85yJcGWEovk66VXiY7/m8irrtkQLQUQ/zOLJ1atu+kc
Ki1AfIiDuckeMenM5ZKfChhHdZFCadY/+aYUnnhNzY9DhKpcesNDaTVkbUoi1/YK
nUp13eZkt8wX8G5bRSKHDY9izWHAS55JkGQqIzQTFNiGjJyYzvZJErDpEd2CL3kh
Jxrvoo/GcXyxAWuKkSnO+vXdaOFqYkhvWrme2x2JZiLUX2JTR2Mz/0s2V2c3SSfo
dUuBUQC4UqerMZS9vDzhtZcm+d6nIAT6miXrgk+2J+Zn/XxD0EeWZSGdk6PIEmto
7r+pmo3t+Z656XdPmRf/M4vpAnuvpRId3dnhUntVJ5gMoZ4600IX2MX3P9i8jnYc
wNCIA7ldU8VYteD0nuW/obF+HU390xktYwZjJoIZHztAvG4+T/jPk9QeRkiIO+zX
ot33gGBl36CsERoyVwyUdaXmjL1gw534ginWgnkhb6cmevGBgwFl7aQKShOKvI6j
rQahR0wiVQ9YKEcU/ea85dVR3OOc72nlz3tBStS+ypmiRr57iMmOLd3qECLR3Jx8
kfhM8zrllNRpx/e8UUhsFIPybKQq84uCmGXaVEBD/vuROpj9ct1EPm0wHXFOz2KA
UujqqHJd1566zAzKENEHhiuTpDUB/dszl2kxnUsIijy8Y9bT6lQaxu3tn8VlbsBu
1IttmN+ZxXwKpJKTrdBjAyY0w1+PfWrRLueWeDDzkRDtLQEq0465bVH4ZB+kDw76
NfJUaD/pjr2IBhFD1qqi95s26IyJ7IFIX5YahPOBeQReyu/WYlMYPqekD4myN68E
RbQVpbqVhO9dfnfhgo0u4MKY/fxp0Bun5SzHBInNWmPZSdyQ30dlfV29nh7yYRYo
ZV+f5tOOJS2CfnFaiDCViJRrDIfPGkmXgoM5UPuaxpZ8XG7p5Ko2eXv73wOE5M23
JWjXPQo3MTH0HQNV6FbxK8e7YyknaPMZShQ8tpflztKPtKaIXeFSSmLE6mDftRfH
WecXIBdUNMfgpJIXest9T0CfSBTuaTipgoZtBr/4hetzoBfpUvbweDAijJNQEtJs
om03IuGlUb+722LDqPxfSXSloPwXNJIf0h0rsMUdDmYgcUy+tTMitN9d2tk6AJTz
8psLjPeEkTa/YZz3uZG+JDw2YfezarAhPighkOe38P1bTLcJ0sLjdPxv0zbiTYpP
sPkhHdfZ7I50MLaU3s8o2zgWhliwSw6IC3s57+WXwme7C5QbG45oBSMiuyUaryFu
RIpL3UcKGDrQOVDbos3ofwB1ru8BmQ6+C3WNUMdL8ZkDM8Jse/UG0MNQ7kbrFnIy
UvE2vAsn1lLXoYQ5k23QSw/OQCDbkNEuBmH3q9Snqd0CCTgwdfCdeh+3v6WbPuBu
KGgfXEKpp5NsIkIcTc4dvfvBvHKyWLc2EmEQLXqaGkU+TeQRA9FP9bJ0YYyRS4Vr
U4BLQuv+ZPPV+UZe/4RKh/uCD/ndGEgpqOCGrfOdJmAAeqK4A231awP8lKyatc3e
PRsjYPnCKBAKtk5i/h9hmkUq0hM0/PgOBpJSUn6Pn3pWdwIZbizpVrh2T891js1E
eVnxWWfoVjeMvJmsRGeKFTt5r0A8lH/SVNS6qNVWNV1cAQUpIZHhfvnviwDHp+r3
Jfh6wrKflHtWdGyWKuNpDXxBDgFbOHLCsou7QwCI53LqeoMaUP2by8PbpKhuE99P
ZaqeFCE4bkZ1n5yP33AO0qVq2Kkna7rRtagEawPUxsWVT03+gXw6PQmiVc7PFXco
1bFaDb0W+ylwVqJVBwnG2zK7rIOBEaHdZeb6IrFnKHtYjd1BS3zHDrO5g5dcpaMg
+ez2LbnQzNokS1GxErHe3Rum9ItDueDEI3SpyWcZaUjlVKD9sJbVor5g3uToxGWj
f8F4oByZ2AbaEY8wHuu+SB0zGaQ7GBhA4SWvFXhhaPAjo9GPf/momkostNGggiVr
8wsusrIM5uJzWSwLNrkdHZfk+C5chhHWcWzA2f9lPS4zHaEQHVzfWMNFCDm6MIFw
+dsp1tIrJXLaqoFm4PVt3mPe7smonjgiq+olMsdbXifJxFOCbbnuk5SDWHIv2k6h
KArN/wTRXMHxli7FigXB+ljxSj9S9PF2ODInS9uc4L1RCfw8bu2me7x58AkwWOSX
AqciuaznG+/J/Ca810DVW6m9JM0akg6EZ3an4mg/fY5JosfA+Q0wMt8FTiWkJ6fx
x5kYRFOMIO9C/zndxhDm46qZLbsYvTDYQ9kSW4/U7EYnR0aKzwOqZ9G7rd02r/52
mVniRuy2/dQPLT7GzuTzCDAc7HN+wkBu/SA7dbDGnVpAMLx1MU0YTBhsaH/xJKFN
RzEzfBD3Wo/N6q8XHQi7h5IhImloMAMU+IlAdIBQ07vN40MiXp99JZHfKq7IcF2X
Ad3cnpiiQ3WQEulg3oD6Kma4kBV0/+Z4wPG6o19laMRXm+sVOv9ziDR7MMlH4W6z
6COFdw91GjcHHCtlSE1aZ8klFpafGuoDwF7wR06WbCivcz385ma4TZqxL3O20dBD
zsbRs2FNz/hq4Q3njyqbcW9wEQ4kHFChQAKMDD4A9PXvwVnEx2R1+KJKL14PuYnU
y3b2ExyLx6rQBjrQx0dRbGv2f92LaH1ua23fUiIGK8UDeVXadJgYn9H+KVC9sBaq
cX0wgNIP3jsVs+fHIBi6Pnp+2kXYb40AdAsqRi1eTJAC2Ibg/m9RznBSl3ZdE9rR
WY6SUMkdCU8DQ0dKRdMHWFeaA0XyfGxyMVIpYyGwm2ZchHd5XXKOjadBDxcYOhBu
N01cpALJAxs4MhvgvIGvRy5MICT6hI8KEq87TOoo02aI697C60GRg2KNqlvxZyAs
iVOu26NW0Mhz3hg0MfZYNk97d9d66ZpJHrwkqPS4gRyaC+pGcLCVBcA2Cy28X6wp
fcZRjgXapIlOsdX4gDVdtiYafDZqhC9bjzyxyNYMQgQ8J0kcb3+tzPw6JH81Q9Hi
C2oHpA6yJJsRQKtRF2X0O2/HB+w0o4KmLUS1QKgx/J0P/mrSP9ImPwkduLZACMc1
pOzYXfMz9I8f/X+yWmhN1K6G3pIIF6fn6glE3LHnfoZ3g+oj9kdpPBjh85ZUoKDi
/C2jcgVBFG5CI9ELJgNEKZLbdng2IK8zoh01cqmFLy0YqeRcipBS13M7mfH6XNdB
VJv7CBCggdTwDjdCSLQsfxkgxmYyPcFtbQDgK0E3JRsNdbU79ZDir5UolyF+qfNs
VgS9sXE0YTW/HCp8sORRqvdjwB+yuyhEjuwfvBb0Z+fA6RqLOD3iik+UnJGDTLFs
OsI0/HMPuS9vioEYRBgBWMHZQEpzTNqFBzz0C+lQiy4L7101hto6kZwTvutQ66FE
jnzDcHFRDI0992cI7EWNm04C3KMC/3p18ncR8eJODcjdwIfMX+oNMLxFfGOUy5am
jhlXUJUIOPDFQpAYVeia+yEuREU7Mcb9h/m9N74nXSk7/QqE9X7Va5ksL4za51S/
fSffskQmwH/PQIu5i1LxIiwns32sYGUVPjYxtqgKXrh0dcREsRgpidzWO5iySWu/
DKjUCl4zaKJR+0GP6o+UgrCBVZG7tjdrLzIrGUypEOAhqlotM3OXm3Nd1oU9kEJv
vrd6+g1QQ07D75HIZIufXtPvX519FDEbyBF29ExyCv8cye23/apxkcIsTYUGVzWo
so8nEUj/l1ETVSUZ9AUGt0Un2hlWeSoULMsmqw/I+PH4Nej1t568I+T0XmgxT/MI
LbOH4wquP68smq/Q9gZaSH/CwIH3DQztvCqv4HNf46DTNN/vwqGuVToMW89Lc4UD
YRLYMRRyZTq09KzPpKMd3KlYL6y3p5SV7LUCL+pQmMNv6Ujb/ireMZqmeow34Y/i
WMkf10gZN1DxXYbD067yMe1rpgXXA3056tg5N2xWUEaz7n4VJlExIK2nboEY/lop
tRyErPwnzIF19w0uGOkqdpwu34ai0vChNanIfrdL4hhs2WAQMGribFBs8V4+IK/S
aTT5Aa0JJtzd0MRoy54KPXMbQ7siG1Wr5YjlVocMRtHbn0TctCW4/ZNmM587FN3F
Ljp32M+fYi/XSyYPa1qIivO9JRW8kIxns8bF+xiISxpKjqklqM4DtFHRWAw2YWZ3
WPPKfQzAYOQ9sF2Z5ToBxmRoZ3VVZWHSCEm7gkwegp08F2DirsKBBYVzP5TJcyHK
Wisvuk4nQBNHluETV2gyIZeEA0mOjsWjOjcIM7GMe91Q+7y7qCHaLYtIJm0ZyZFD
VTTM2rhEoP39qzgcTl1uNhL+P/LKsZc7GUneObB5HHf5ckFsJIubZcxVZNbMo5Av
XJSozJgSTfrDYERkQCXeNNV7mHx846AFb0ShjEUf8TolWNrp84A12HMPIGW+eD7u
GKaaJ8967j8JQwiiW8DCFst+G4VBzalIKIpTdaHXFnmJJT0/Bn4Lb5QlVP8FGz4a
q6vUK3aMMWYs6IOyyBkbGK9Hj3nZGnKy8Jd3OmI2TIyWN5yT/nyjuoN0gbsOirST
AEAby6zEEop2c9hfbyyNq90eZbYXcdnwR3g/Tyqe+iCJr4FIkQJDu5dAtR4e4/pF
/AydZXRnPxYpanrLHQJ0Ej9CdOeRzhb7gvAu0VPxcAJpaYNehFwvwz4K1zM5B29L
0IzoXG5LDdmHpGr/91A5R5hoGUUmv45aUgVWvp99wFM8ei/xh0vgpc1y/jHtQvtS
nQpkp6ygypsCLn6X9bJkqq1jqAKcmsZyPO9FrqRbvstTsPVZ3JOHyr1Y0TpsQKme
G0227pQ8k6t2XXga2xj7KeEHWojnIWUGj2CIz0xbRk+OAxyty/o+g0xBMlGllYiz
itTUHepdMuTlOXNXL0/J1DhjBiSbBUQ+bqECfgdXSLhz0tZdOV/fZSo1XIKCqSF/
BSmulIvA3HLLc32EUkYFLg27wzqQ0zzyk+NxumBaPKskItGqOxeK7Jd7lKOyH5Wo
rz8NuYPH2fXmfAJz5xSua73jOZ4Vzmz9RjV41i6C/XEhVmUs6uwyGoCIjq3PMElM
sZsIvz8OIXPY/nxgGglQgjUemdfWBpGQ01Gldq4UkifBm2KtA7RzDtLknZsdM8cA
smAYqrcF3P2c9YiI0BNP4FxmfuSBMFO1WNHNT1Wp0pXbYWulQewEDXNPWnzGJtxh
rsyJrMbAkKPzmqDZnf71ggPHDMLV7cGGc5NVIOn1UlNdrkbJMvKf7FjHZbuJ4vgX
slbXfvEFAC2c6vfbcK1g/3/e0LdUYUXOIsdCXdhWq2Uui6P85CkJyeM63YX0MzIh
JyDoNTEa0cjvsJMc0rYvxY2mKljHjIoaHkWiYFyX1pTyOaI35Xgo4yF54wql1YLp
YWKb+wH/fcrIcM63iUOCQ2JEUE5N7SOGW3eEYquPuHdWtdb7bgj7JUk38lKt1KGU
5uYABgmAUd9oPc5JPAkwxWQPH3etTggOJg6HjkwUtnFT/FzMh0UMZoRkZHQMHid9
JsNb6yP2X6XI2oFEcX+M3CgBBSLry9LyFhmf/qaPU+B0Dj2Sk0/xcBgkbZa/w/hb
lKl8ww3CCD/UyFfVY1LG9O+moB8Ep8G87HSpUFvFmRysq4LyIRJkwgaJeG/kso+v
450/uOFzmuY5CY43h8wCTRhvyVGvOshae0aslHfwxFz0SESaQ/OGOX9G6/MwobgJ
eof1274JChHk/KJtluvllPrkJC4atGoutpQ5q0AIctrP9wPJPubBdOUfvndzGScY
Bn/9GnOOjuTbPVcgfKx1VcOBHigXf4441pqib/ELemDLYcQiySHW2iy4JxkTrcat
qY6qPjPUi3yRQJ1mX7aQnZXV9D4TfHbgsEBxOK508G0aCayobq/FVGGtgQeDOYan
iS0/PyNEpglFqCeuRY9NUo97nYffj3EdSzzpiQVjovaXeMZiknMRL5uWwJio2WS5
Vni2Qq3eKP9yy5wstJYNgjCXxkslhFvbfkTWHnSTYhvmlF/yVm6DC0zKymjW0fd6
/mWkaCbrGQjOeFb4aSo2aQM7n6F+VQM68a/0JwWbaCWLJ/GcPdcBBBPB2j8nqN9h
wLAfU2Ae4H8kK7A7Xxb3JHYuFZymol3YxownqMU+YKo6UfbHE/pWDptluHQ1o2jt
I0gSnkcZLnMZZLO+jSApH1ce/0yqUJS4H9lia4HvH2yqmHUKnnbtU1k6fN/76qGV
qDncBCWQ2xZSK1Fn2Nxvq9BPAvQS1G25PNhhS8R1E/gd2qaBk/DTXVI3HFs7O+QU
l8T7FQhEzbohFpdsxl9JvIzT051rCtRKEWs/qgi+RtZ+bQ7Gyz0gY6TolPvXI9Ai
ms+HWrIZzFXsMma5QJU5BodVnBKgEG5qAwf1tawjJ2k1pcANUjNPW5pK0Q6KlHxd
z3tYwBYc/WdM+C+NW8dQKdV4BY5XLF7t4GQ/TBb/8pRsqPk4Cgu4w1jO3usk5/Gs
EuEqV49Nk4CN8DlmQHD3C6O7rdKqBdvnSbyn+I9TV5+CBBe0HvaWngQQFDOMDA2g
BpLaSpVlRqQM7ljF6yG/7yneFpvAmmKc/hFSrDiOzRHLLhrEstylbI2U08ucOMsR
qaZs5OoY7F9KaewXidhOfV8Etpiki7vOHSl9CWq2a47cAkxvxQIFlGMZi5hXWv+S
gNrl6oRFF1p162wsMPDQeY2jQlcPAuXEY8FJvxMyykJCrIWh52HzsYiUNwI2JgDR
XD5+lqGLxbqHLkHFpac5ZnuwPc59+u4q8f8wKXYZQJ8dG1MZZ/D8CIKaCNCKlC9x
U0YLLie3azIbdUhwZcGVpHKoLUoFWCLfTtSRqXac/3xMBwjHCVD35n6PTjSFBntW
6vD0Xj7uTNEtDWj636yzBtdenz+o4G/V0j5bmC90HPEFznOHJKnRzgUg7yIBZutq
KIhraI11JVnGmFeRYmSpkWAQ2mIwUk2ROq/JWQ1ILxaGq8rvllwOJAbmvEFp36/1
1vwjExN0/fSj938wNKnTlwstFEyoFLkadlZPcS266T0vFnE5lCCcsgcPbaJswM4F
0b1Qpxsxw6GvYM5DFCtjg4iFBHfbFM+tUNVxu9kYzvoR4XTtuftGNJzmLre24tDj
zNDSWYfbkFi1JzGpllyScRMQ+hG3ltu71gBJoh534WK/2kAaRjUZ8JUYSvJsyeA+
vKHIA7U+KPQDGkOLBy5WqTPqlqCfUqUL97RyH9+l+iL1KDZ2zt/mkijkJqYXJO6v
ybHguHs60AvFsh3YWuOQRudpV9vqWd7CEY1uNUzrlmVFHxCsfvL0nxooo1Xh4jZV
s7OCdpqXbHH9Mc1u22O4emuMOh2pohtu/cmpiYyATWWZBl+hL9y17WgT6mhTJZXB
aYQHeyTPJMaJE6lq+Fj/DtRUXVMgwkMmahJlhnQ+tWjQh7TXamYYaL5d9oqoE9DE
aUsqtylmGJlK6QWomRbgLn+/IziojhuukiCfIPEzdh0r6gPPxOZCjS/bSFYxoRks
fD44mjs/HFt2ypirzH+Lnnz8k+dSmYwoNYwbeAZBiRgoDmwSSn38+VcVXEyyPgtD
psaLGuedQuYbX0kVMqk+sNznj671KJzMz4PCJdT0JxcLhpt8q0efAqIt0ykSTBA2
XAC0wLm9v0zF7MCvXRnTcK4zE4ksYdzyXGciaCirHmJjsZvKzzodOK6ewASyCEq7
krs4+y258jz8gY2e/aLqiF0FDbjF5iqhn0dhmbiGn2th7SIY4Tw0D3FPADoVwBTA
3Ju5JQdxct2uMvHx3zAqf+CisNEMsIddEmF5nzUxh7XvGCD9S9/OCLrjnt9IgnFa
g5VREUjSM1pRtj/6a4scovt8sF3sJUZq7b1812y9Dgzbub/cvSDfOpLSxCWNK52W
Atm22vEp42pcrhJCfGKRvMoKmnLwgTwTo9VVwDBIFYi/HUeupWXWfSSYLNl0Qqlz
XumKIYXZA+kHHRjvowzYV8Uj+6k36lHAE3zOuKnSShribNWm2gtJLKokv+4o/TOG
bO+Gf6BG3bsHGmhqDCFTTemxk4bxBC8mPFXWzkIFVjOlq5LYMozzP6h3N6Vrw3ix
181mNtMBw24hbzrV2/2bQHiZboP+yN4SBxWQnhscUYjuNa/gT5H8WmDMVVgIpDFR
lhQ66lTs6l6Oyt2X6FVwqVF6YyefnxeQpvBotbQf8L7O/Y66kqNgUbS9Qa4Y3yiz
BSm2AU+GLazJ8gJn40yjcPj0l1Y2RrBJA/rY33sFSrj39nxeNp6smEIHZiQhg8nz
tvgOr+NqI7E7AJdsp1QTIU4/swdybLnIbWdj7da9Hj243AvP/lWAQWRo3aefG3YA
G2PYRNM99/kgmONLFvI3AxBUwf5DOV1fe/hWX7/p0Jf/7479/g+7+b0ab/byFs3s
d20douqpNV8YyZhh8vbybQ/zT7wUoBUSm8jXId9OiHxm/obMV653YDjkYuAqt//v
9WNoQK0wQ4Tr2U6ZTqGwTfFQiiL/UaobjNKjI5zyCJtKjO/qjpluzseF26iY2uJu
ROhYnEonEB9QVDwjnXnm8OEu/bjFF2cDWe2JLecga3fN/EzCdb801WHcefdbXTYT
z/dwG1JfIYL7uSmxmk6nYOydiChNrbNApkN0OrUaYpv66O47k9HxthsdoaYqgJ4L
xwxmSIk65o9T8j4kAUebCf6fCguw6MubzA3TWUuCUe5KO7yWo8eOLwPJqSeXxi5W
MEMVx0jln0mjaR3t9PJuP1vyNMYdu94DXGACLfdUgOgaIoUMXwZHbLf3RuCzR333
WdrhrlTxj+zAcgmY7uI3S7xlIyj185CCdJ14PD2x+t3Mih8SdPnH/l7wPIwjQwCl
RkIgAy58wbCKqOaB/IZUeLo4iQyENZb5Sh1i3F12HHaJWGQSEHMLY3Ml5zpcAoOE
OSjgbw9wCa3ko9YSwxkLkhdSMDsjdTG1X1q7Vgwb7vT5LRyOSBEVYZQnRo8cWEb4
NEk5qxVI+yneOunLiijxsaq2vij0nSr5IFlw82DROYSrKwm3G/znbXERiuVYa5kI
NCGpEJ0S1gTC9Un1yZBX9zucwWFYUyaMD3u1KTIfPf0MNdNiAgD/i+WuHNcF2NzH
sI5ifbub7Y1sWkbwG2Q6h05tJL2pqJrpuAJqeIV9UGfv+uEriPxSNVkSufloB/uv
DPzS+hVLx8AFlx76NEvsyiIrI1xlS9B3oE923xJ1RF8S7Z+riQNj5iYdOvjqWQRY
ROm8wtYhTfGyTDGEAa7Ybjz382ntyqSCgmR9kcphvr2VYCecs3hXb12z1Zh7Uvnj
NY5uCbM0Yp/1bHV3VTh/AO2tMxUJglel0NbF1vmnMD/dotUmyuskuGeCXDSIOkl3
fKfcukFJvlUPWE4dx3jXUsFNpWtGZunHSODxFlbtO9eMIMbh86jv7nO1R/kir4b+
g2uNWHJlWuanN4lIsl1G7rgjys+6WRFLtBB+8GVYsvyobIaApw1uOewqFoh1cM5H
X+T7c3zp23Ll+rgtS0ZlejqPnrs64qGBzWnwbY2gV8bYM657ljmSvv9P6r2b23+Q
pDwF6qv/DalH7NwpGolN243wal1tREayGLDbRyUB9qccYrOK4MPLYfFBi84EiC5+
jdSDpykPnbgof1pHBTV2Uk3YMXFTzX6wv2JcikB5WuFJST0WrfH9mpOgdIxHHreQ
mRwjUdJ9Y0AlKU87xzCUjLcYpLMIqtYz6hKHJrQkUNizeqxdyUI3eaA8OORQDgoR
yNNex/Bx0LwznO04QI4oCsfQx8jEclZG2RK9DfJauJP2oRtM4Gwiw4JMBzY9ygf7
bGwDkqMAVACkaNmUD/x9+2Ti0PmSGIiAWWD2l0sNjkUibtb4GfKUbenfQn/GYO+5
OAfNTZxw5VyO2QWtFlX4v44lx/1RNCSV516rSkYh8z+hC7RT2kzRnykJHephZezV
6lJ1og8sIfmYaSL4M/rajIpbKRscCVMaEemdSqD4NP2cCDo6AjR0/QnJuE3qPRMz
hU9Hb85JsUjBQi+nRat9TSfL+MQqqEQf/dTUHuA4DEmOWo00ksrWtHeKzMI0J8Ot
oLuJ2jVDFOu9nbMHiUbrDOMKt8udo3/a8LmLfoRjSsaUlWSqtwPCfg0RBZZ9oXRz
m9dMDX84R4fMVAUS/7SuJrmYXI6kAuYavirDXnQ7vz/6MbDE5VXP+kMs51QQqoS+
F9baQJsbw/RYBYbZQNF+trObXjAVKFYkH2jluBt5SJLAlj5E9xhYyBY7WJeFvBx8
709Tn2cfj3fs3BvLqCHsXO+RSGTMQR8EaFHEpft4VU7m1ls0ZWz2jYwbog9FjLeP
5q3edDAL7DpHu5t6ci4pqCo8Jjd3DwrnMmNhtGsPqSGS6mzOetLvRcgcaN7RdrZv
opq0vl0ZSqnMG4ylk79nrvAu80St1jE4eXo7yuDpSjj2C0ttUU6+S/B310DY4OuP
CN4ZJ1WmLZyhPgKcdrzUSdWgQm6CVr8FVFt9MYvON9v/lmQtiTfy860e67g7YHnu
ZReC3acDp5ue+2Qn0SA+2WsUy+kfmUPzCYNjPhyC3lYss/4SlZisXyxtGASTmeBe
KLMH8rEFdCsmD+4XAf6mtYb5Sh//3m4hczCDoh0HHbbvl755QJPYhcVqHz+jpMUu
8i+9hZ4fkRxsdGsCcAe9A25bBNF2/P01HSneinfcQ3Drejxtt1moqRHH4zRRVg98
NLh4ua4941oK/PEbKWlFxtm/J+W3Ppty3tbep4NnmpvAFd0gy5kVC+IefOX36sm1
ZGp7lOEjUNUbnYzlkILoFel/GUTqCPSQAuM/UxKzBTL3ZthM/XIRo7bR6Ki8o+Ql
lJunvxHOEf9FzOrj0hc3rS8WcL+8gb8N/JpqmOJZUOFUHFZOokXSDxXFdcgLKflw
O+eUnmhBYEZmMkMK82n7ZwZ1/W4IthfPhhlautxwAp8WaHocjWyC7RzI9DlxNPOt
l8zn3ZXEbwQUMys0S61XyJ597IoPkwlfoAEZ9CG5KH7I/y2/MDPZd8HpMu1jfTmp
k1E54yQop8B87IGt1B2g+p3gExgAfFGbeRhbLSdEFt6YZZLOoC1p9eHn5gzEtUfk
6CF335kJgxERLBdM1GFQYxFGgDjZLO4phVvxRP3qT/Pw/F4/m2ZmUnsZRn2Scjoc
DJRA7MgXuH4IVPpfqM8OeLH3LXfgi8qXs5Tqtv0cne+f3//HiPWS23TxtrKjFhzi
agC0AafsrKbKqHr9ZN0dGUolxvOdBBirv6fdf/chPVO9pM8EXm0X1tcEb7pI9288
l0h5jiw36gz8t/3OFHq+Jf1ytDLJet4j4mMLii+8QOsS1z5loL4WtAt74s0FOfJe
KhXvRxhgaNI3k92EteWh5LpmVfQEy/HSytr10E88C/Jk073HV6yEDbcgLtfT1DwE
U5YJr6uADzZ+LRrXBatH3eLxAMX8Pxp5sXklZwUP5Rob/oM+r26MA1FH6TiLal8H
Rk2a3TOdh2vri1Ig7jAMBWJMu5ICnlwmyZGj8KntJtWj67MPGAiC22VCfIMz3iNO
I+tU6m3dOZt1A6rpKCrscv3pfIhF9daw349elb+sgAxiwQ4S33kIk9uyra/yMam/
ch7FWAtWSG//FMbLj8P0sOtNMgycSY4YjVf3395gxo8CSlGOD2cs+wsvIOSjnFGr
QubB9L0tZxhAv4BUbamvfGpCw4yrDmJ5+RC4HFKD3A7LZlamKvy6X1wDev66518B
egZKZ9u581uA8oxOoZwdJgeBYT0nDZuw35nKRg4mDxGV+YgKyJhP+EoJYTbsh/Jb
ED3QNuU3fU1CABbqU599umQpmFLdN/6rZ1I/5m55dX12jyPLy4VvEOfM++PhBwL7
josUP5Joe40EIvTRXuHmM0eMwcVLQGK4aubumoWi1euCG+NjT0xY8JGt72DEyTUJ
04mr8JPRt0TopAUX0yCV3vAGG97Fpb862EA+/2n5oFYumtR/BXKQGZMGy6PTIqBl
RRT1SKA1GEfCeOmtyuO91yz5sXYRID5a0aVpJTfJ/SvuXDhnbTs/A9ABTYuRCn5k
bZaW7/cNm7HNGATkGrrJfBpNgtVpKBqm/nd45VtiQ2VoNlFnwELQpBvX/QCTeRwh
7PgnJcINBS7Ybu01viSko6fNYRAZFyQoW5SOTHpAJkiaGtIv4WIpUwKIEto108VI
HWC3r8tThYvygrQkWQg3r8vmZz8O8YzV1Qkakac7PD9sVUjkxvlRYWLI/gUt7wAv
y97Ah1Z1MvkIooyjcgNsutPofT2HAXOKZrPoJG5UAKl9e8T6bEqXPFvJu+f6nk+l
QuC9kAt48U3T5KV6skRCHUN0ciUl7FrsmJ9PO6TCkO2vu267xUPx8UC8nMd8nWLQ
9VyLNl3mFxN26sVDtUm7XhnR4UyOuz2ChbUv1XsBeu4qYr7+1NuUUBwTL7KmyjC7
PRub3XL68SP1cxyib2c4MgXqBzcRpLem7Axyv6pyJs5ZEVFr3i4Cc5PQUnSO8x4G
owL/JbgI8OFLgcVoC2YRQoIavnxM9XTJ+8djwJPE9v6a5/Vy06EdkuTu2TEdLnYM
LwYUZIHi3YSU7kw6+j703SZOxZGG9genxooPeya46rywt2fKENA9KxV9srF+BpVs
7jdg5To/S0aSGr7SAr9sP+10EuqeYz6dh1cJd4kznMB7F07Y3eth8Qt3htU67NjK
/LSn67vB6Iw5OBLt+IR3Pn6av6ZRsIUiKh3T2juatEWUEWotQgVNe6Tdbsvm2r3X
Nj8zlY3DE/oaswNTB6ITcd8vEMkXXILWG2FysTleH6nmBzjvshs3HWOu73rdSKZC
l5c5SFrNh8H2d83skFvIAzyE5fVLRuLbrBqmHt5ICnms5/86Rc6Se4MakEYitYut
ybCaLo163PKgFUkQSpMkwvMXmArbPJEZ8y0SCPf3G4B9DS4LE3YwsOwJodqc0Zfq
T6b5iaUl1oE6JFRWHcZtHQA/sB350XfMiIKJnA1gS1QpFvzsTAxiioUFky/MTKi0
YjbuJHSyx7e7bNvRLg46k/6duh+AYEZXbZsJ3Q1Vt+CocOJvAAZYg43dvyokD5Zi
51z29ROQpijPXfVzmu2ns5VfdgrPnKZ5pORFzStT5ueGxasapN64Li8I1fkCVs1h
FRzWFK7qlkvvcTUJd1NuBfCwHu7oCzr2H85VMmVzS9Ma1PdZuzIafyHBX+78BtIc
bGOVd27DhlSgXTBmDsGspknv3WuCBCiSHcaDvVuqRpPbLuQdn7WYz5mTn+8L0a9v
i6n90+8sxbIYM0ix9A+zarniPUpqerGdqychIQj5yLZ2GYVlq9/wxtQUKb9MC3GP
/hddThWBattIfgHEnB7Mg/rHO97T8gvRbnhXXJJaWrgSGNENMYW87Tstiolk9OWC
u07DzmbyWv3e0wjWySID5u/CRawKzjswSfnPLUU4sN7zbSHwcGsc/4+Kov8xwtJE
WZrJG+C2I/tzcgvPVQyQebtJ1NMqt21C1TDBjgKJhpiqr9s8THWc0O9ZdUw7oIcR
gRN/3XKFNxIes1xh6dSWOO1MlY5ZVs2mb8MIdt75d34rpu2kSlM8mzVHmxbwuZtE
iYvSNZ+Wq0fq6UWBUREnnAtXQNyyfEUijeNqbLxCOkFDxjTeh8wxcOfnR1OTthb1
7KKsqdH+b4WbZk8tkZVq/uWMR9WPyle7WXF6ZjPBp9ajdVVFRdbRYLXVG35HPyjz
enS1vDQtHtOc7yYSSnYD8s9I1a6Oty6r36IXLYfZWEaiUF/IIcebj/KZktzFRHod
I36qKSFfu4KmXskCYRqPMYFJv4iLJsm8BkwFDPcj6/2s5Tu9/4X6jZ3X6ciE8CWY
fmpG8Bl08toBRJcc1hKGmNKG1Tn7R16Xf0G+MpVZmfEjJSP1pr0nUoQcDN2ArxbT
ThuoL4x57GSppL2zjwbI40PFpfb4bvtkuUvEqd79SROk4VS+01q09G78OeWLnU+a
OaKFC8lb97U8NmqM98UqfUVeQh3HVHlQod3i5sLe89Qs3zrzgNaN2ixpI4Ts+ahV
Q7hAZ63/lO5zdQPOsWc/OI4yUTVOOm0rp+insDbi9QdOJ8hm2tAoRsUb9Mk/gYkt
NkSfud+7etnHn1Hac2M6k2/KRpwOP50g41heV1shLcB0HA/e4efA9QJtM3+AuTgb
YfdY4pj6sUgohFlZh8BG0GEsTh+oe+PPn8/9PJFgKC1qRUIz4J0b3AkoA6mg0R3j
r/0forEBM90UiwtV25d8UvTkd1daDSCWDCpLfp2mXG9slV/8XV88vuC9T2Vvz/eQ
8J61GgLXun/yc2SUS8KS7kzcx/MHS2/MXA61AdhJ9+xZa5oIBc9ytXRS1ZHC2Lo6
z2s/yM9s/HB4vdCmaF7GmbDFkBgVyg+YDMitcVjsKMCS4iB7BaqEuA4WlzMwQQgp
6ky0Kota4Pus131JnLmNc3LwE5NJFb7Jd19WEjCWuRV/0m6fV1hCbgZwrA9n3/KT
R6vC1gcAkXAJu59NI7bdRYdhItsogaNGLiRLfm8hIpcjEsaNG4GnQalr53ewXTB0
Q9DpI+uwuv8T1DWBqK6v823wy0Sj0mYFt1+gfWMG+ZG86k/VVNZ6+YF2khxgDca3
TJVr96XjjPZ97ft2G1X+NVO+tPHfrj3k0NXcKFQFs3KuDqP2In4e6M9+PAdvIbEV
h6oyxRhFPcXmgoM1FDtM9ZApP8UeZN8KPTMrw131+yVQrLtpMj/8KLN0noB9pSev
IaUXDqaJmXCX6GIhextoB1z9HIgnBdI+M5qeQpZOmheCtB/pYUwWhKBTUxoD16vW
zx1orkFxL0/Qz22CfakZbfpDbCoflNa/sIRESIDyFITDDdh5H4sp7sCkRZ84C6Jb
Ljc8607O8o0ZsLSviXyxC0hGFGshAfmDN7TxDlJFYEEgCnl58rXQCJI6xVHGdVGe
8hz+dUe/c+UstJKqBzfNXYoTEoktEURM2g4MttBo1hru4EC9FN1wUTB/I9lTgljc
mqtn11tYPbSDEWl9/n5SBe4M3HlVSBZcJ4PmEnf/Bbcd2vVbyk+2vkULyf/v3CTT
xoQxJ6TRQxi+EgWoOH+/WHpT9L5Ow9xQVrWlb7Xu2WZi1ZhU3xyLaegXbc2cSK20
kyIIzGQb0fvpNpJHxQ/GeF5WVhAxBYRAnSysGayiD9ZOmNnDqFQTYDW7rEmDp2BC
Sd7mhYvI6oxe+OwPTaqjZOju4KYckmZ+dgOi6UonILSWWMV8OlKdUh1CmHZ+SJlw
1SvbfNQJhaD00OCluvVsj8M2kQMoVNkCDDtEqLbmgbW3FI33nEC7qS65xSB+hLn9
zlHbwKNfp1hhoqJGyXWH/Rb3OIBVbVrD8/QeiMXruXXEKRCIw0XFr9MJxUMP5JEL
pQhDL7UymxT1G/t2QgL4tGCI5a5/ZwGZq1itxQn6hRJe1Oh+jUltHatHUJ0rbU5G
4ufQzOz1kkefL5LEYM2y2Y8OqO9aQpBdpmKAytEPyBN+EP77RfdRSzpqRxqgibkZ
W24PTbq1f+lLiBXLRTxneO9pPjOvTVmfTY+Y6+1wOKSaTKAGsNPkNOwbilOPWGBW
mH74YIV99WVoG0l6JLpEhv0r4zuj0SN6h1GvsxMQc5Uk3U/6XGbjZIRx50tajrmM
C0eG+P9tu8xNSk6/G7u3AxxNr5eXRS7OcXRQiXeh2RcChk/0ZuRALegBs9gGevnv
CBCwryPDxnQiuM+gVOHsw2AWDg0Efc+NxK3IcakLr1F7z9754F/Zfc3NCwcp5lZ4
VAt9KeLvzXDnX74cjb5DbaB1kc8nPL+iEL6Dsix0YVxf2p86qjcSw1kbjRkQyR2H
jw5Hm3zwG+LYrjCOqCXdjCFeMuuamx88YOR7vGjmj87XVD8s7dAzbbH42yUh3sEF
H7sRoIwRWisuA8DTVcYqcNiiXLO7/ve1huPF3n3hoA2aVj4oyEDs5FctnsPnOIa5
YEUBAnMxZUgdBj2G8mYZ1OlwbGD5IO7lsQ4uGo8XvzkVEV/VdSEoiYaPWT9bnMec
XfKhIFs1H0Dz6b045zYBZAFKAoDulWCQqlWs+UqTEoRlTQK+gynEfLj7VeAPWukn
v2g/akBeNTnvRncInsnXNdSL6JxsbTuQ+WIZrQTm6lCGoy62b9QFpOnH5LI6Axv9
2X3hsSsrelGgI1uDuS1n61ejR9dvPm31yAqdinzL8SzAU/7r7gxCy3KvVTKhxGwj
F3DKEIgBuLk+ZdpDnGXzW8uJy6giJ/FuscNDyG46DWYcDb42PzneLiT9kObxYPJ3
RXsmNzOT7sx/RoGciG+QckpqtVIxodXmAsvncNC1A4p1eiXl/B/hVvTMHlMPScPP
/05BethPUkDuKTmKVrz1VMb3raNsCdpIrtUes2N5huV7xFbLz4leKmIDxQG/yMWF
JFngO8XUSyiOCXrD3tvH1TIEZAb0EYWq4JYbUNRfuqTqrhRmbQW4krZIAdAYpGVb
3IEH+QpAChRinhM1HbYgQiZYeK3B+m4PJP6i/GiW2dFS9VkYlZWnv2Fo63FjxDLK
LUbWGqPhjQbwiipG2DgNNyjmCDtWL2JdsbILYol1A6rMrvsgoh0bMz6cqp0dU1z0
H0DCzRAeFlulptQxSAAVuw8zlzbKb8BlJoQWnKmgdRiQg8xItaRIQKUo80o0iTHf
WTfEKHD2WWCAkc5m8Egb2iCpWaet7oGM4Mi+gRJWd+gKWrUnGaPMTFwXNMWVeHi2
onjQXQWfv865rNkGNdeUmoBy6hTXHgHpkuMcikWp/skh52E4OEnbBnGvmK3o63R6
WW9O/7TDAC+vZKYiHV3KVuDphaD+wvxMBz6hFgYSRu5K5DsZDPKEEkkqiti9CEWg
FGMMtDnA99g0DQWLKY5DqwOZ0Algzr01Ny3QYH1lfyi/HTVUrVpXkDirMAEuUrkk
zDJiLIEKIL7+gNnOrPebQ47Eycz7T38HJV9fZweLmkNc41Q752LJ/phVgcNmU4HD
ub7UdAh7MqNw4TlfWwH8K5E9kSJQX6yLjwRFa+d4JTjx9A/hhFj5qwks4kcR5CKt
OWXXXTDQoMGz9rPgKDRsjEan1jMLda7+B2fkY/15IgdTB/gMER57neeg27o6l6lB
0fG/aXcxkhvJ9/y8Gk4YuYVP9CJstLFCTHiKdFmHOh02x1v40O5DqU2jaXJxfh7d
a5SL+PgUUqfHCGHTQybtWjK+A2f4evu6OHyhP93Q3T/PO8NYVwg8aho9+TCFN+OV
jzOTOo+w7FgNRTbQAssPP9SC6ucJqcE7B0D4FgUOu2I1eL24Z9zodXXEgzhzr8iU
kzoz6+dd8UYAVJzVhXr3SvMf8GZMuyI4eImcxlseM9cuhml0zPyhXJ+y3YPsxwxd
QKA81gsJYYh2+X/TtnrnE7SzWAp6ub9gFKL4ML/idbUDQgjIPaDzF0j25KU0lOeK
5HQrbIUcyJxkWrgIrgMRwJDbKzzay+r2ZCtKZ0tPnRGCybUM6BegIsVgzMeWKo1B
dDyX6SaqEyZNayt/x8phZgVskHoyRxplxc2yMrTrGK7TzsdRGCOi+a8mAbUIWVmK
36E1Czfip57Xkx+/QImyYHTkp4YShjhE0WE/4oE5LGa3a3oQuJSBfq1bw0T32V8a
we/GdV9fhU3SNkmbsTcEgopXWSln8Zs9hLns+Ah8MZJdIV/Bkw8NFsn+df6ofdHo
GGLrUxcjdENUhnUDtPey/pWNlfUZx89tPVvANa4VLcn6AQjGajgLRY/L21GKpiKQ
myg3ExDpE6K9VfKtzu+JC7PNmgwtowbwE5VGY/1bPlj6EnT2DMzyx1D7BPaBs85F
jt/Hhax0XWVctXQ5EhIKhFKdpD00l/VCQvPkShkXFEdh+FvwptBJDXDNEb3UX1Wq
ONrzx/zAUMlNoWi3Sv7b2C624mKZozmdONienAHP/Hr3strG+M9i9OrXyv/mZOOn
F5MHqUXPbyirFJEYVma26maBm12lw9+Vjd2OIv3eqjOeCU6Ri21sPx3UwBCypwqV
HQbcsB8eeoF9y8+K6b/LH/im8WqHDGvlrDyHm19yBP6BSnc6gmanwdMXo6/rdRUS
uz5qVf3OMxp5149lf/9EYD/VYOPGp/3kYbx31y2xTx3ck+Bay7xkKfMArCBsKJSf
+26C7SZ4J2ydVaqr8pNddXVnT7X+5+cIS8K0JMn6ipRTYqFeRf8MrdE2kJIflIaj
hbuVsYfU3W9q5GUbJg38wxM/yXr6Hu2KCnxwXRADqoaSLC8aqBE2HtbL3fk48zKx
1u8tWbvOA4X2c07AYHCENDG+1Gc04a0ZaPBXO9cEs6I84nqu/5VzstKoPWdyJDv9
tBJw0gIdUKTXOdfVYwyeG4ZLqRzNVNKx+kXaGv6bOT0VHcKZwYWy3O32NJB7ZCyP
8oQqJu259kWANlZiT0RbjSWLjMHXrTbimL58ortawSBGyKGjs/o4kYQlG8HFRmvJ
PRH5AVy76kVfsEOXh8cvRgupx5mAblnp/DIXoHntFLYw7k2i0bpEo/kt8TOksMDs
AAHN3+xB6AytU/NX+AaBzLK40/0VTMJxczs8lUWUw+PSo59r3QTBnbBP0QB8FzG6
+uHXg7vdwS7+ynCce7Ko9jZMAyCYvCOvLd7AFsStGUsbLRV+HyIYrJHNCQjsC1RI
2cUo17nILDA6r5x8MLJj8X+9gAcPlulDGG7vQHiTHlI6fnXFx0ZyGXCGvlHbLYHN
870mv3YegotlybSG6F3UuyO3EMkBZd+3qCD4PhnlPheRvxnZh4ph1a+duSN8GLh7
49VhUMRUKcd2U84xXBoqm637tq0mlHdIIOV/A2N4ng4728vrO6UJ35t61vOlpllb
bSgpPqI78ReNMrzRVyPWGGq/Y3nhfFEQX7ZlwV1Gc9HDZHqkki812jeMEGO7xT3m
938seBypKhUwEq684sfCIM0aq/7lwKJeA+QVOmzzTF5vTS7QuJhM0/HNStx6gl2/
5mNhvZC1H2FGkHqugkXn5uftp21eDYu3Ysa6yo6T2GTtE1j/PiTPlvpbtQiYFZ3/
TrXD17iZkwQiuq3EgdemS6Wknwj44vQeIS33uDf5SAWblQs7pm5yY3ZEFaGdgeQ5
kholfLLUEq5R+7p6zlh9zCnEjhmELP+73+LabQMXHAk2OkLSg+AIBRBqI8agcoPM
3SNRv1YnSug53EiBdadJOvfvSPckqS5CEPQkl1XvCsQkYCR+Xy20xNEMVJ6p+ABu
sJvoXNiH6sHK23HngyjYz6Mk4M4rCdqWawbIgvzpPeFmpQZDO9YwskuE3S4j93aP
W7nTolRz5zVl8k5iRNjz1ArRq7N020p8UsMwYO8rtwX6XZ+3KmWhS61NymLlHt+s
81/820HROg+v9tW1FWzp+WIjUfOuoUWVu3YSJrBo20qhsoYahGMG0Zfym2+9mirS
Syffs9KiKPaFH1zTJsuLvdz6lNWQ/vA2x0PTdr/unBJB7Q9ABLluNgIkHAdueETc
8nj5CnJwbTFYzJ2jdpKqvJf8fWTE0lAP8RlGVGDz6QdcaeATkG3TWyiQpV+gN1hl
WoMT/jui3ZzpWXZ0diNcbAmVBJtn7qcryQ2791rrKWKddlJ3leQ2H956FwLdDTAS
Vqs0maooF5+HRQuo8aMWntOvn9+uptrJ9WloPQeG6WoXB8SHPBP3vrXXAGVJwIph
2R7vdKZUyS4GdZ1wrn8rf9WDynExYVqaq2e8gsWOMPCmrUakXzZWdWlYmWKqG1CS
mZQokcBvZKBqe4/+ano/0W8QFJLh68+jttjnYMkdnbWsQnApY2gfH+j5KhnfAI6a
m0C9RM2yVXuc5E+p/w9o9J57rArGUXN+qBes8wnP/8qCMAYpov3rtgvOQKJZzkXV
yhYbJy+h8igD598dVk4KpiWjrLhHLNMrwstL3buJUFoWBhiNoiChhVXlYgAypHed
F3FAwFssVnuiXdksW7iIMMGTgpvxpv5YJ9DK9VU4Fsqpb23cYUQvwTfc2FbUsCc+
nYzcJhj0KphYs6lX6F6viqGxCJBd2IEud9cqYP7ocoOJbKZQubrPJiBt3kxx3EZa
sUr/gemM1AaTDkj8y/JC3TdSOOu0JfkTr48nyJw6p26evfA5mi7OYNu9K4u6K2g5
Lp6SbbiZ+VcEHGTyMuHzQfKWKmMRDLIuWZQM1sWRMQOlWjKLO7hOVLatONiCQlYK
PCdHaDHiDXoyGqxkpqSmjIndRVdb6x+SBq5h2iN7mN8nAHZs2G7ZHhYWKLjIltuB
wUJsYfUW8D6925a+wUfokylLBChkuR/AyFklDoH4TdJ+bYhuRdZZ4l8UGh2O56FV
r1S4KV1/kRbFVquKgC/XJGX5X6ymAEB2NcXRzBcpngDGa/G1fdQkYZjPJ1xPik/1
u8r1tV17jIMvHmtfvojFUioFLYT+J3mswXgT7sNdoR/xSYQuPrq8+b/LSGR6UXxp
x9ffrpoaVv7a7aCEBBGOWK2/TL+E2REJvlsbx0+QpDhuPbKpQMUgatQMnzJxQqUr
lOlRuRKDhCO+splzq5JrHNpt/ezOx0NGXRKF9reWOsdI2E+pfMV4MqzOQ7ALJ5d3
pGsfNZk8ZypvixyWfEB3Q3Qz/QghXz06IkhAIgyJjeHlzMjKetU/7o647LqR1yxO
gTfe4Jba7NlkCkU2hPDI2Yf/jhxrddtLoIqymsKarGiPZZpvmTkx1gdfyAQv55gH
J91YMq+Cp7fPGNyw7TU1kMq4AvCa7Xl3oIVNk4y/ui3ikoNE3zNJEcMl/u+kau4Z
FVkCocS/gSspGMctszAaE204GZN9WaSsEqHy+QJvDbHTVFNdPjk5pCgr13x9WY6x
g38Bad65z0hvhH+N7m8r8ruH/WRPk4LOCHN+A7IS/21CqU/8GLHaQYicylYWS2/w
sht/Xbbt80iPzUNYBMSlh3RDB5rODjY2Wdzfv1WXP6avEy0wp74OVxcu6wOUwZOg
xy710HIe3WdNbFFeiYznQPwE+qulLLGsJ0lLyBoJx56EjfdLx05tjTOd4kgCpvag
rWCC5KecUCb7AI/lUeGBZRNfSWh4T0NVWFSPkE6rZicPaK7v/jfYjRuWqkBmB51u
g+B15PEaZCO3/iGdpl15f9oUPrBdtRbo8tXMh36g1+/g5F2TR4+L66koMTIu/CeJ
s7zfSOFD+17JleQg7b6aPK4ES8VEdFqkzw8rvERtNIvDAB2FUdj3Pin6j/1hxmb7
fOLOdZ9rEY30Dxzx7DleqkXyXnWMrbujomJhl1Dzqhew8QQAh+bRmO/Z/je/eOJV
rzW/04gi7do9xhlCSz/ORR6nbzpbSWH+RRiow8g9UFn3KaGV+g7gDd8sP93llG1H
p38LuLSsav+Np7wnMOLVsrUP8RuxPR4QNTK7v+8Rkkl4/o+fSiqpbm5yhv+COJKQ
CW7qmp3+Ye0MFhre9JmYBjzQK+5ZUjIp9CA+4Wnt/wX6H2IbCBfBjbWtFZNiznBf
fax5WIDPcW75hiQ10fLE4CqAKs9fWqEl9sLbtg4fChwLjCvKQOG993xLseZNYcM/
hGXCgWHSgVwan4Mlzixupq5A9vnhZF+vCaUYnVz8zUhWwD9yLNQUOvY0LoWkPrH2
mr5svHagSYwFJZVpOCYmtjl8kMmmnLFmv/k4KG+SICSQHystsFFxxS87c7joqm50
ATdpem7VhATfOX+ZrLdktiZhRm/4JiybRSwfWcrCprG8qZQYqtRzfqok9XyuJqO8
hVAwreZ7AjFTw9t2bsgPMnzl6hYNfFqvl2lyZnCdvN+fd69VcpMv3rcH08BoaS0w
R8dQA7TGerwk5NxonHZlGqTqFvtghzfbeSyoyEuhE1D2d3T1JNrwIzXG/kJZIN0l
Z6BN/88UyE3E24LeSfGAAnfnxvKVQZO99g9Ip1qJNMnhyAEMwctbFIUESda1C7iY
Hs62b81ouqxAcnhb9XDstCtm/2R+yYA7Wb3jYunK4lJZvsYofrZeJT4pqjphrn6O
1mJISK9ThS0xzDGXooRgDuWOEAZ9axk0Xcsyfm5v+jsNELJWoJaJ9p3F5I5wd1mG
t/ejX94jo8mABrCO+g6guUahizDA5hMHALQ/aHx4D36czxbXt4NzytPKPgaJx44a
3x6FonhLVNFtMqoQQ4KaCqYdN5OLmZAHgViUvNaOM8jDCUyl7pbhtC6jHPLidbFf
7XAeGmp0XcYhFB87Kyq0sukTTjyentFC42sU56TaFlAOIbKNmniqf+2Twrz0xDze
9S4EBpCg6dUPx6Xd3yom0iiXG33I93sdVAB0FUyjNapYvpb+WhcnsVTxdHmffEOE
Tna/rLy+lR++OV4/yPncQyoauJZ0E6ByIwYhgSMwHe8uspSc2EbOD5oB9sU35fUs
A6CLaeuxXxGoKq49ILkE6YxNckSRcXi16tq8TEpFWAUuWGtfzgyWZml0GiqPWCYw
vjcxzqFAyiy53QD0geDpt2C3Mqz3YQQtv2M0wmlYcRmdIT3nlnNiJVxKjpJ9fKS6
rqm/8+3GvnZ5cHmUTvauIVPN/IXeFEw79LuYlLg8TVigrDNbxQB1m6byP9sd+tTy
odl7Pk6TTLHTLGyaID2v3Gki0lmLlTGwsgPokrBl/KxCUbZQbydnR3BiTsRxIZc3
txD83o7exUMYUxcV4ZFRHlM0I347liRA6BP8YuDWIKojwkKrjUw1i8eB69d/eRkS
hSEn80/GidESF93wZpqFTiHru9b8rY6WGxE419fksEGQhRTm+6I7eVo/2sMgnu91
8YpPZSlW+j7gHxkJySYGXaDLQMctpUvDDTdPUgJZrnpzchodeAr1iX6FNLujQStl
2R/ckzvueo7dCYMKfiA5WzP1E39dOCc3HRDhDk6HiG09rf7SGnD/ppzz2fSBmX2M
spka6PIkXo2x2CmaS/+49h6iwhMarX8p/0UuVMIJdz16SwNMK0FZBPRNK5J41M8M
2x3cgY160Wg0C3n75L741P7uk7x4q6Jxj4Nb/uAEugjG+TogmqRLIbonczedPOYM
hJVT+RjXPQESgoz/iX+LkxwlaXF0qk4ePOpe5MO8vMXZx/Qj27R2lEsxMn3SL+2O
0qi/0BLwCtiKKqbVhMNBoZwC9scGS3aHWjnw2IKRbu2FOlqOq5UyHFH2odg60VjZ
qN10U0EKhKf34Rq7GTozpvJoVD3fFyobDwfv32QQUo3u/1ULLkBzdoiMYgv+dytn
nOQ4b7xzUcosI9bshVmTvXNO5TIpyQeHFb+CiZ6KZP96H0Fn4QOeELYtMp/steuz
5h0sSfd/LXqnoN3RrjzvO7fU2CzZ0WBr+IxsCuETR/KoWx41diSPiB48TyNkPta9
QR7olV/i0YfwH1C4EDAkEdqqsuRK4OiAqkfOUVlOH86pQXDw48y2ezmyYB5IN9Ix
/h0YqV9udEJiPwYU/Wdsx72TOAjdk+CrYCKUV6k861zX5qLmBAGVbU68/KgGeA8L
8MPizPC9gHJeqUkOd/fAfO0AjCf8mQ31lr6Pyl0ObGu06+skVNyTV0QFEhB+cp1s
4+X7JgFTV3599sDlSlofJUSGnT9OxtpyUfP6+xzizyf87KTxtZ5NYELVXF1a7RIn
b5xgZYe/XWrZmrJMAilIqRJFkfIFAXUEPD+cxKqS6APXJF/A3PAfc5zc6V9bNxkz
B4d0OG7i/MhOMb6Fbcy7oaGEvhdLhbbdkIwLhGEtLJZEgbs7+MsLoGTlqrWyfJ6k
+Ou2k+77voyclkSlWEiAZ7UYdAbaspKu8iGnCY47xzOyV00yFvOQu9bFf73NLAGB
FWDGcTMOG+d0Kqd0THa9/kHod3JJbXQpzu2DKnvqYmKX3FrqgDrd+C21BlvdrjPC
Pn2lHdsqAmqLGP/H45MpQuxY+/fQXP9n/tSLIKq44lqY8plN+sA48g/UzL7A/9Ir
mhKz90C9huiCpyqOyEyIW30ClE2el4KV0S31SG5WFqaCgKFV74emMXw1OvLuEFoT
FDBXLuVOKS8tCVzpiKo+HXK3KaA9F5g5L5cS5FVQfZ3BG2PD1Q/7/w2m9IhH+CqQ
V3GPAiRBA+YYM5x4FN3SQOjEKjQMnrWCzbQwCziLdpdclp+Q3P3deQ3YTP//5FuL
7jU/nsIqZ5OeQCwnQQYFzWwN6lDHHKXUqukQ2j5yemXJ80oGczpMdk5b04zOrEHZ
vhdehe0q7Uh9P4jnL3nRinqFaMIYpzQa/P/8pGnQHkso6oIjm/JEFBBXCddggnwW
6kd9ozKW8tznoRfnlbJlqLXUc48uR+UPD5JH4ZIQePemrz46mJi20Sz9MkK4d6Ju
ZvcaAdiDLRf8qSCNokPeA8C0YWYyWyL7i+I6zZrHBhlqFxHOrXn/Prq5rPB/y8lk
b7tGkeCxVrZstOI2AyqGlezcLGNyVKvfZ98sHKKl8/osoc3MMqhjdu6tc4lKtIgS
usLUnpXoGzKRqy6pyusXNxuERNEcXtL9RERBjhLA0mOaAnr1g46Xerl/Ik7TAjHp
ruqjtzUixdv3Ee0LXaB4QUeMdAE2zyxFvFMZh8bStZpdGrO/ShCeM8F6SscuLsT7
hjy+QTuozWgeWxnj0dOd5QcX8QzjvpyGjqB6m2Ynl55NDoIq034kGAkGA5wJUfgV
3ln0kVflc63QNpXEyFUHSoUdgvORVvplxka5Or5elt1bfviSNn5Y/Rv2IEt7S0RD
PgdW4848l+k4vlaKAaLt1liPLGE+174AeCtNV9ECxFb3luPnaQ191Sl7iKKoymyu
o47vebV7qXUJps5PbSsHS3CT6fBNtAF6ljjxpyulDdlQ/gb+V0EgtV+RVjabERYr
oB/Ha/iPPYQF+T4cGL4hrqdb5xscQdIplMsBZIqGGpgisNVxluq3XvmAI4hDft7f
kUntKfRTu/3tvX6xQPG/rGMHILmGUtSAnRubQ1DPGIxbIzrwBL6TA8CgiyhJGljw
5oK88PfnMjLXoI51CPOEhQmR06FzmMGljoHCi4CcV6nYjppaGeHJ57xoWXeFM0xG
+D1eRkkoXDiz/dQPQmMHeLYsPhyHfdrSkEKJb87VjKnkZYP4BHk8gmBf+hn1vHVt
eDDB/9gDVvfxpCBIqgFylVZkYmfn0PLTc0WOkJrwefRh31imsxWva8lXw2A5VUWF
F0SZDhKT5cV5rMl3GNTzNPMHWBAKBPEHA587af/9MVJF4XukhPe7fDHlOGECVMir
jb6Hlome79NCy94DdkyMgUkEsW34QJlvmK28iGeq8xB+1pRt7VDnHQvJCAqFpynN
9QhgzBBsljoPvXFbWtXmVTYbEgbo/VtyBsITs5q8iuzL+iw5iMXgscXngPjO6y5T
SYBv8SbY4PNrB5FqDGml4W/VV/wb6CDs6JxK/h24K/2W6LhJjnbmBmksOkoeoSEW
D5R4dE2gNls4ro3vfhCy0hhzveAkhAsPZz/MawvWDLtdCLp+9aH2hRTweGJtVaWr
lurgJpi3jI62VCjs7DI/Pbz9DELj2q78bQZRrd2G6REPAefzWyncjloyXtymTzrX
P4KDCHfSPsXQ/PYMmGDLo+oiyAD8Qg58CIBlNS05PGW5lW6r90iSdnduqJnMosac
E5wP8JtFhULQ/RVKCM74cQk6m1Siz0+epxuFBCYQc3i10J48YVsLPyzTG6y9VDji
yDwa6f13uxVcHpiACEmNuVh1xkojgXiEmvOJ3KoCoRmMpXoakLZt/W1PeYXSiXfC
eMj8UaTWatp9PEooeJNZlA5cll76R0/Bs5QniFRAJR/HlxSjmU1v2hZZ2R+O8qzF
Bs6vuIWb14gBYFPdaTPFq/DGEHf+30oVhAEscPY424kWdiPe9Sl6jVnGIAuPLH4x
pGYpTLaZRIcET+S62gQnP7rhOSDBuxeRPeNgvYQ4HPOSPJSiNsh5qHhDKI5zQqxo
k61Qe/cqTs3aaf2OVD9oTY14fmhxHKw8/spFWC0RDOKk2kvHskkB4j1IrvrqrO2S
myllcQp1kUT6RFU7mx8CzzMmlM/F4jzEd3M1F4wxV9PY2Jknj9zjbVshhdPL0hra
cToeZ1/Op7Ch7Vic7+lM00HXzjBoQ3naMso+xWuiaYzspNT16BRTnYVhwczZ0d7E
l+kJaYtmRw1gu/uUfT8XF0ryzgV/zVAaSqgLK0BEdcHX2cLPRDOp2NnX1rEH7G1R
eph8ox7WxPbaQ6Dq6FCCHV4x5J7R2SWR7KVtjMc2mK1zUMlcc2JtSHlfnS0huGxS
mRRqzoR8mXe4ngGC6R7ChdlgTcJrMDdeZ3yhUkpQdlfX9J0CKodJBYB4uuNpp5nh
1Arnkc1jYjooMAu1K3/qXsD/+173rmbHecAJkiAnaElxJc2XWXnV3Zv+ezGQfnQL
rmXsi64CrQ9n+3NG348UD3T8GYQFO5F23n/D85ZJL0vgnZ4DBBzg/NyrI9AvLavX
4cZpKkIioXK6QjFcXzsyurym0De6Lkp2YhJX6c8342w51nFALTOB9eRneWcWjFTQ
IR5j6Md5fHjICUQYd6ObwbmAWcTGg+zGM6lr302NTzn6U9IKaC12SYwPiQRaqSOp
JAqtuQvW/XcN5x8b1TvWrHvmvOOQ5R9OoIODiZ3h6uzRpmHhyuAv5eL2KRYIvUJN
LwtvDGr7m4lBT9JToMzLgc8TN4ukWuqpvMk+Z9WpBB1EC8KBVKGq+EuNFBDq/cC8
74oSoJ+0K55V1w/cLBU3l4TUZgyrEn5MVcxheUa5KoD1Pwc1jt9DAjGGZsAz3iTt
SF8cD5OHnslMlEdaFi2A3cfo92HyOa4pi4p+zx6/VIRn2PsljOwjffYLYKzm9B9O
Ic+edDrrYNwlgQqkeUPjGgePUOlrzL7qyjpR//nAQC2ykj6eqCpWxvSV7Nym6nw6
AO1PrL2v7qDFZZxg2PdOCzHuOQUGMys2fh9/+oRoq54YFsDT7GWP0OL0p4D9VI0H
oH9eQSh81Ra4mHAUI8tqkyTgkQku2BmZFInu9vozgJUckAuHsScpXpbM5exkJfIM
5h6Q2+zDSEY2g6r+Npsop+1Ip1Q1wQPPIwCK0vls+vJsdKpNcwaPPKMza5JLotgl
KhpWPHqVZqKZNwCSSxTeeJPcED5Sf3pkBDTQYMQJ+Z4ck8EkaubXYSRMpF3UxsSg
HKNnFieTplRVVBqZzXa1NtSSwc2OrGnbkjvvmg5dXREUE2SYeQOhl57Vcs1Io0zc
QqBFobW7QpGhfD18zO4oDEOXQAaLGT2rO7mVVqvljUIxR6KurWSTBw4M/fqXbzEc
PGJvmRlln+dM4f2c/utLiwQ+Ou6KuamCX2HGQDGpW7AwbURJnGIg9tQ549QFbyNv
sGH3zg7JyaYSLFlZQcHIISngMNdV2dcE1HDvMiVNizA1kHDv0sczVIwBIwy2thZA
kGApN7XArA3lWdlQ91eFchk+DJDvHIo7lzGJFfOtMh31qx863lwZUs+vtVdWXocc
ws18wT+rol0RhXQ/1VBrlnht46HLcqmPqDxbgohlnNj3LPtNLjwg0FuGyqZG/9lM
jpwaseHJfODlksjIv7SJUZdtktzewIsxFZNs4Pyypgd4Jd43c01RfCvkCV6T3UM/
zCgbpLNmU9r4NIbBjfQxEMSgdGiZLCeDf2NIgH0kNIaBe7r7nvcFiHsMfo2UZH9H
pUcYcLrx6hhN1s/bdbWLw2E1yAL0iz6i/xd6Cjk1aSM0nv/edMJOWsjFVTRWSr7v
Jk8HQTdJph2fqbGD+0bl8xAovIdg5P5KLuQuROcyg9rHup1KQRnvv/isVJx94ggC
F6ZVdBhzHymLPkTjKCiOlPI+zIDs1Jy7n8N6H0O3ecS97uQqq/G3MlW/3imfcSC4
mzSWd50p9HddbhMLXg9u0IW8Ay1SVgJ9yXPFjE/e+E27UHY3JXwAC8QBXqNfPL23
nB99nfqxASnRdH2wm5DeclI6agkD1GpPEWX7vyO+2AeBDf2hgqBVirvnnpAyRFh+
p6QFEWtd5kxgAUpvFUT8NxOBVIAj/Rg+TVAENoC/fkCMWg/6/1b1oPjDT1py2zdI
gkP2Vl+IrXziuE/Nbjba+9ViO046noLs42zUPbRskJvcD5EmH9ZWSVXdV1UPwWr+
x+JiZG48LQVgUbl/oeG3Y+jIE3USfAloUGIVsujG3o2Wo7TUk/xRyjtm1ZllAYCX
Sgf/mPr22pUmPzSrcdJFXBE4Y1GTdXyrWTez79SneJq6LaUfUGoqwTqeWUBlsfim
UKWRQ069Va9mxOAHdwwwbw6enPBnuo0quPQUPDeTiJMDMVVZHAjFiC8L/ewvVFUD
qjrEoatTiuuHJY0GjVRLdrBGIbPqxTHvTMEsXoBKiNdRb2MytNquK+cuYlXUs6X/
qFWeBEWGjrBntElrVvFKJEx8+OPhWJhFPv9xQNAIsJElaeceK6gOrhqbDeOfYyPr
5SYmRkX5l6g2ScG1eX+11YbcNzKOnvJFPB/hdBqYhiJsaYmIT2Y1Xcny9+2AWtKB
fy9tnVhGp159aQgMxhZzXNPJOjeEsj22JkAfdi/vMgtDQ5RunUbRu07a5QmpuwSv
bzVs0ygFoMBMN/68uPsAKzgJjgDGkqfau/3T+Z+Ndv3pKugznEsWEFjNDrhrgcf9
M+m5AihGrwvUSjSuVOmk/wm1skXHcFI6nsiG2rW3PiY+Z3oR5RMwp7uOGNABagQu
XPb0Bh9ruOdZ7JyYHAocJXCwJeGnTlK4dVPwYowdC4fn9PRxuZ3SRWsDxPmsl+nR
aJ4ODk1NbSW8G39THqWhv2HiXEjyeHt+crhPtBSOQpn3C2pcBFVyU63GfVzfziNp
9HYpaG25RqqVAUR9x67KurpV3O3NKUkEpJ6cf/CfkWXBuu0BwmvTeE0bAz/WfC4t
WC7+WX584FUgnHG+Ijzzz8tPNi2u+9VSnI+jXoM19As7MiHWaTeCKugugW0wwbYZ
w/9BMIR62mI9W4L8W3tfT4Q1lY5w/crxj82nOzWGiAD6KXSzk+2920zTqa9V/soU
jH/Tw8a5ql97bAhMKDjenToIRF+ihoOZqAiPWAF/OonKgSFBxZn/kG/koe0b8XJs
V6kHJn19ev5kFYRKnVEoGTX2apwThlOy+mQ4UznSeIqJa6zTl3HRXh5Hnk/eM3es
H886U4m5b9eEVkxub37JXd9UD6mCeMlxs8aAzHN4tfnrl7ZC+xF48GiEdHppB1KI
MtGNkiQh9HecMuv4CUad33huVUksokrDn6MU9GEtpGvwdnzFV/UNAQQv29dDvnej
IvXUyxZW8OQBpZKmwjPX7cguRFrCJ2gKOs0WjQTeDh0lrdg7dmqa0jdeGa1UcGTw
qPNfRp7C5qUNo/vt4vBOyWn1TiZ0Uu3jRb9SSAggYMNX3uMK9U4SYz/wWIwVlFEW
8f4s2uoXfeDNFj7+E4/WYLOY5pRE7e3miVdipjA7lQLWBZj2qDqWEiNtG3f11vno
s/v5FESiEXQDgh+UHLZI2ySeQ7IAWXXnHHh+f8LTQ2f5o63kDimYhp/DPn9+jqfT
TYDRXstrHBFLK+LJDSZP5/ivTYP32MDQtdVK48+kgfGrByfxR9uWVMBd11kCfu36
VPKui47OcbqdK8bptibcVLdq/5/U06XiQ663BdxGbt1eDBUT1R2oDo8oXjLjfLrC
03XIIyci+Mypn9GKO99MvMd0rJVR8r0EPzV2lFEbLUhWoFg/ZLrxEnYkek9Gi5UX
y47lpO8VWnwZXcnEn0EtcxAEhqxDdAZNt59MZRGnctcqGWqZ+FFZ9Fw/Wu9qHsc7
BpsvxdCpSgzEhctguK9IcGYJgy3Jyh7KaJaEjPO3rnjZMVXksT8neqJRACeLeqOi
2JeKBV3PRjL7T8280Vj7gEjwdBb6PZfMG+3yvyEqiyY62vxVhF5SoEtxYFpatSek
yavh1s1XbieETOHH/w/aKsZBG2NEh4060WL+qVkR0gUgodUu5s1iDrhHTJ/M4Qu1
OgK+9zCfPWaYm780xkotSS6vVV0vKDRD+9jKaQE/dSbVtQOUT9vmxM/7sy8yGXI4
xLMp2s+egrFlAvuKzao2lYpmA8nvAn9mPkdR5jjQ5ZjZDlutqHalSAPIKjqNzseJ
seaxrwYkN1Dhu1mQrhIk8OKPr/zCYYzXIxr0B8wk+V5JZgfxl714s5Y2vAr8jfTp
d3FsF0BjkwSjoc2j01ai7cQelgJ+HqpUVMppMZM4Otn0TMffYHTkpEi+CPNWjMYa
/KoAOcEgPSf1U8KL4kAbChhbBt3xVdkoIuTIc6poTS/OI+Xewmxs4vOnACkj4Y9C
cCWmFn9vaVKZBnzikFuGmx4RHczuQ1HmzCk6q1cA1BEjqQZgpD/6e8qkuQBvJXpZ
c9/P8KeAlWa1GciZJkg3e7fHwJje2FHrkalbHBek1pGwbilcSnwkmTFpn4yFlXNS
fhS6oDFirMg/14snZ8fv/S9GWl6ujRNTYxadRX9651BdlQFX9oQ2QVWReQ/1Mx7z
niQI1APnLrkisi6URtyXEEBHM6x9PLfc8HBNWKuW5yzuQX2FM/V4wQIrBBp7V9eX
H5YdF4j9MHuiGWRu1UJd5583K6mL5LHZAncWRWHHrvt9brcw5erkWONToXPgxyiH
HjnmB973IeeK+E7pQhbYCIm+Nj30bgBR5J8aeFowiYyns88j0gY7EYjMQyDB/g9w
+JFDsgAuh3NVQcyJBK4jPpJstNcJlX5j4cF+rF95NRZbyaRGkpZObmVOFTJjOQoh
0kRZmAHxSuGhCWNEaQQEeSPbOK6Twfo5ZyT6tfKNv0TakKjysMb7hMIGcl4fWNnD
EQSh75+OPHg7xu9EvIVnw8nMeyGSj5p8NAa5vsTwKfvlSPOC4rcgjuxcTLLvhPZO
odJhOfghlWQTvndNnl7Ttk2vXWRqwlk7fWbSUU2KYvrGiE97Cpm5AxcTfDp3jC9J
Mwr23jk5caHduGYQLiWJAHWdZtVC0VfG4heQuNhj+zTifDyOdkPN0I00IhcM4qqE
0qbns3ZuzpMJonhQoj0M70jhbqeuy08VE/hTKVpPq966YwWrpCbVK+9Qx9bXbwwa
hSHp/WQZku4wLt0VTO9F9tzIuhQsoMITos+iuFltzB6dkoJwD58gKU3Bqt9pmhs+
sjQD35MLGL2ZPX59bHlI8zrCS99x/fj2DT0ZpMzlj74y3TvupnOH4xTl9Gu7huy7
UsNEcsDhiKQrl3Qr/JTf9xY6ZJ3vyrvBIqWmH0SOyLIgTn/8AwMm7Sqrh7+vpc+T
0inrcUynxaa3NRbxslZs7fXBE6X4auaObbgvAdMF/hg/IlHZgfLxHDSbX4Ibx1ve
HwGD4Sq0i/bUkh0AQ+GDboq/ikTUVZnQLJei3nveJ3SYKiPTO+FMK21D2FhpSEPZ
ILFW9BxGKJHrCHMmNxt7eWI2iaTigHKffJapdRahuKrPasOpXOlwkHNmDxRoO3Mw
MmerWNzRBHjyD1mDYVAe2m79sbDIxPc9eO62dKA2b0VpYptOV2xZdljkIMNgoVz0
FiFCd2slFzmVLHP69NEKZe9yMZAUchWmHOe5JBIg4b7E83cKZg888yrqt9eDEU15
ZMSdgmJB1YAgO3g0Q/pGdclC9CAmiYXciZ9vn5qWM27vZ/f2u33fHiP0MBvjEWSx
wxSw34YAVlVrsQFuL1nQCOyoPblM/Qfz+0NtSWTeeCjCRjSYfFeM+vY9yJvzw/3p
lCMxCjFxW3S/6sewn/GX+WyLnCAoTSMXTptv0V1SNHUFgO1pYpI+aXVfSBk/UL77
1mD1sakW6FsGpq0bTQSXgopYr0iejS2NYM61rez9R4NmsueK9ZpQWR0GtvAWU+Dv
WyfDsuRpIQUsI8YZJ0/MNJ2wc6eAK37lY5RFd+M7nxnsx8vIpNbmrWi8BQxqWScB
O1qVU+4RKYAqlHkUhAldHDdoVgmjCga1Z35rPFs3ZIXzKgkGWTO2yybveIyaDHYT
6IIVvYhebOeC+xTad9PeHSv5mFu+fEiwpzgnCdi9B5hysvIQSaclYZ/qs1dAAshQ
3C1vuf/pfLSiXF42Fi4xHbR9IexETDybs56fm0pWje6eSriutnB5f+eAcHPCwV06
KhVamhuznQSJsyusOj/ctKqhbWoBiAYrgdKj1rN2cBWrN5jlvcKef6DX3Y4mA4HH
Hna1ju4gM3oRfTdVpqmEnP5vPag1iVIxeOtxbZ1g9wClUiDzAZ55nbmOv4FSQrAv
atNIfLb4kgGLILqTWi0Y2i9ygyQ/sVxoZi/OWwnybgT/HDULBhVQlb9L260VgJTb
1czYd7rPlPGZXUjf1d6sY/Duh6oJzKwRaSAVk9fTzUWoQZlMFc7KDyqBIS0qw7L+
o6I+v60kwMBODVC8DtmF6lnLpl7cfbxcHoXJKQK+sFy5DJ8ca9/rC1lEWdZvnh3a
v9GT9JZTEwybyXA2RH51nOCQ/HwOZxeIL21yiKpSd3PAXib1AgCOcg8S4iHe8ksU
VA4FbAsojLwm9msFtcFLIy+FzHZD9ZbT6dQbNbYo0YPKbRQXlDu7pBoTBa0fX95k
Lwoz4fDwBkpsw0aXid/xK9lvrXYiRMoKzdUsLYxR2Ctzddx90nMv3DOrW1hq8ZIE
oB5yaEoxaw6hac65jWrv9FkM0BYFRr5Cm8YWP0fAw2vzW/gDdXZRfV9lD/oviwe7
R9PyUIpiDwyGPhrd4T5MBIYfDg8NW3qMIUwBT+oiDSoJecNqEZhQd84iD6UXeFcn
FaeIreBr/0UhICF3W6kf0IjMCSq7WUPDGkUh8SWI6uUHG27csVwjpYDBfKrjyqrN
w1cePW7ozAwhotTkU+w6pESpodMLsXhrdmVjI0AEOUUmyHldpWJUSWER8k4uHGtH
KbLgvG8oFfEsLTgQ1q8vO03Z4VhsDY9IWLr8gIlNYfMo4Im2NkrjzFKwre/jSyFi
MKKtMxHou3eq7oFfrFcaaZ+y0TESbE4vNrlyt4FuyNS8FPWJivvYp2O3qyzIvQBL
zUEa2vcKSy3U+GNXwyuCk9G/kpiVhaIwd1WL96I/BNxp4+Jm2b1K/jDzKeAiN0K7
1RDWJRBMlvd2iwYM0x4bBLC7p0xcL9Z9UrnysP4kVN4mDacMcZxdkxDSTZ9eiRHm
rZOjvecf651v91cDegQgmBrvkoI+J6sBqxVVRM3B+YwxWvwuuXmO9H7K9Hb9ox8q
2mWVwy9oYbdplq0tIBtV4Y534jadxfetbgksTi57lMYRKo9kP0dmuTWjvXgKyfZk
MFOckZCArNXObCyVS71aAkljtK+Cb1p96427IB0+dLXkWLOVp2giSsqhn96VLk86
CwJMVsujjvsXnePzv5j6L30Asfe/Up6yMALIOkQaKZTHBsVNSy+ndiu006N/ompk
j1O6/07IgE0Q839F1jsx/8NWAsX9H+URlQRkaa8T2UScJdV8JlRHsLNzjs1+2G2Q
UBsKHdORBNQwZIqR2VG7L1XPki69OKGaOZNwQaRN2NY3Zb2I0bkG58F/2MLo6ZEL
JzOqOKtu2HN5evdjy08fnbU7/uhZTJFMc7Ol/Q18zh+zX8P3CFbK9S4sM8gIRs0F
4n5vdlc9JDKi6jyZEvAO5ihc0717WmMwG+rYnpozSCnnsZCoWjuCtmFaHf5IP5l4
0UtHL7wgad9Qx32btoXGfv8Mj8pQoj5tx2wcOwdGKkEiEJCimRopRYv5O8Wuvp3D
WKPe4dFXv6S3RgzedXZbzEmteQbREMWldqO8tpU945ugvc6dnj+rOKo+WsTZKfc3
Zs9DbGdQNkdmhatSZs4K9kpTG16p6fxtfK7GFni0f/pKy3FoljLN0FgIrIVHugNK
ZB/FK16VGehNmBBXuVsNGIDiovRzNJy3tVINBT1sLolJeYxVECUFMgWaFzZW8KO9
noX7kA6IeFGqiPZW7WsSLKOHo1rs3As2Ad2d27uATSyJvmCjyI5L6u1Nc5FqSPKf
1nV8v90/+AgKBqhh4zpoPgHDBX6EdESmk2tRhXq0jldhgj2w1CFJLujR5trYDmmJ
S4K5W/rZBajF2Mn6mALhywXRgqB4roKXcv0VglQWs3rOKOmL8bU0xIqsPmMglS2/
zfV+09V2NEkw9a2JiLTNlUVtcbS/rOeOrN5sGyD9GvQY1y0Ca9xi6lnDOAY137f4
omX24V5Ac9dHgpYex4RrIAsrRMAwnBqNgYYcXp8DwvgDchxPAPtPWe23hoAvWbPa
JMVIK8j9MWdGF0IARZ35rYhhVYXULOuC99jDLFsGkEIM1Dx3gX8wBKMcJSF1Hiaf
GzFC2wr+9KuGGaBKBJdPchyXWwjd7Y4bZ+Wa02AFqHaTrOx0YLmN0PBXN3nhON+b
E0BV0NNmWVTqswrfcuhk5vNjaCIglcMJSE453nwdBEKBfqTK01z92BVPdC2Hh7Tj
0pyLAAS7StNgnW0+9vjBG06oReTY5L0Q5MafB7ic0FWA/KSX+K3phK1Vvi93RkiS
7aLSILYQxQsUqIzmxuqQ9Vm1ludD5+0ZW3lTn9QpNnUywaOYgb9qpeAfIU+w91hg
A00l5f9o6xLzgPOcZr1YiHG+Kyc2VpofkFGqOzZXlOLUi+9u7wR7DrFNQq6FpedD
yDG1BLIdNx6aqtnSrRgp4oiaWQWZW/9Hrfj+wGL7d+Psp04CmoKCDUPXiT8OdbHS
AQYidVvit8yEnnqF48fXIo5ssXbeDyoPFTO0+9GngR5CT2OV2i4GJeO8eJL8y5Od
4duNHUY0gzTRCqnVjb3S9QJ4xQEG94tXIJW+oxXqPEH17e8I7B5c6S9xxPLrVgoR
ZlJxCRDjzty0RhK1YYuP2Vp988ZHcgi0H1VOfhgTZ1MnqdpOeYF5wnV1JQGZfbhf
qMryoY9Xb/x8201x2idfyXki8Q2dWgXpoUCoyNv1HPLFaM+XVCCrFSd44gNurWoU
9NmF0SRLtNiRD44CANDqmpnl4RlGN8fFrGAQBRk/7S9y6ho4g1Oz7PdMe2qoqb9P
JTbnEV4a5SX2nIopoQxLqB6HCI9bMB6qdyuaAbsE3f4GnPAmSqwgjLDKh6T7T3Mr
JgeNoUh0NePnco80ntfI7tC9+Lynmry70FDQCgVt8BRbcyws9saLX9iYo6DLS2xD
e7UTSA4yT5ZKMzMEaM68AoBRu3z2PuNNda7ZTYUlqVDmuBmHSZXnGPP0/ppi0R+c
andkdWofACdcFKbxPvFzJqywUpcksgFh826p/ahfljUbOYCJ6GKBgK6+elbiJ69i
0hOEjzzTCwMdmdikGKwfOgx8apJFXT+LusJuwRngkp5a6fx7s3V1pERpJbdS4duW
esiZtqF+aMc3CkNfniTmyBpayHo3snmyYU4X4oO9vZktPtWFDL5BXCDMnCE127gn
XS8vZ5ay/Tr5SojBgcf2S6sVqHYwB63Ja4K9fFQ96nWSvysciahqJd3V10OBj6R7
OrIJSBIdbuJmLpmhoyLUZOdkbWCERGf152vefRuDmEUaNCmeoPlqK1Lgn88gogFd
/fKq8YHuiJzA+KAol33N6rZi8vZ/QWdkvR+q+fhqmImtRLTG/rffr8GHGfu/LAYF
zC14pZUUpFxjX6ueDcnVp1/7dJaDTLBZLF/vSYmP+KiKHPKTjLg/dgFS5Bd8MKCt
QCrhMO+MgrK3KaPb8StsqCK3hp4yC8DDf2VU5Iiwege9JYIJk8thIM0cb1BjUZtO
VyQh4m44N69U7u0BlIuR0YzGJACUUUUl6SFRxe9sqvld529Qx3kd8FSMaVxh/FRy
OyYVvt7NemuDJrhYmXmYfVc7sTyCq6BK+UvSdPkvGZQ2VSZVSdUOXAMczYRTo4mD
uuPFN/SphsqCmoBBLR0ZWfDgjcx8QkbJjmL2flQhTODbvCMkP3LrNku87lsgfJqr
8nURixks5vic1Z0IpcKvtAG3CKrRV5NNKk1JT6ii7CGWPPbzptjlbjGeUO9tYnwo
sMaxfzdxYmUUNIC4c7phfMj3gR+mkqXqKX5zkLSs9gVxts+kbJyyXtgFzZUexVDx
E6qqSgPFJNnjMSLURJ/RR1yBOXtIV5E5p8IsDuGBpVWQYt7Vt8qSIHGDkme5n0dD
8/9hyij89v78psC87KrUmBVz+9aPp8d24EsEPPzs/LT7Zxe/hc4plp1xoH2wvhrz
XepV6sIg0OaK7n6gOPyAio9rSXO4UIw8iBj55v0gaGsVWeBe9XyDt9r7EbsD36lg
irvjWTbphN/BXGq/mrO6NUvqUN3jIBKFdunL+0/6G9MVnqSD8H7dU+vCQEwgsvaA
3iPubNT0y+4duBG0uhSsOE0eolQe/VkutIi/nZUhC49P8UUp4P8qM/7B0QA6FCFX
2I8iUETh9LLrlqbF/3fUAB0ck9ZDkzv2YwJgEHHOSnDJz79jFVm54VtqwbIUhZds
iDipI6sSBK+3mZY8hTHnC1vhOTWNBJk2Jg1ulM9pK7d68Gqyd0bL+NVpMS1JakOh
/l2C+B3VplRe5oHydvhCAb9PRiH/WmWXpyt8+U7lwP/6x22qTvoeOGxNMUuuf/Fo
ULtH6Bx/+2uAwL8JRvbYTeUke9JBNlaiYqLTQfBM7R5lgj861j9FPjBrYb2myn+s
YMoH58seziuUgH8jfEhjqgb3Roeu4WSptA6A5tXHo1skMJee8GA4Zzfcih87GrU1
jeTynUW1WtEQm7WPAv3T7GAWMf1LvM6/5Gw5bToDFtVfuga9XVRK5OPIFPJSZcdz
U7/2rn21fsU1ktyY2WLb3NiS7/6xhAZqFTJksumkZqDZHqyp+HA/1W1+x1ZmL2a0
lPjqf1eI6+SIVm2yKVBupeB4qiq2sl/C8ZYj8PB2VvtWP6yda4+nJip5K2nZUGdy
MwkjWtHkTjy1cUajKoBw7D1a69yvv+2nFRtno4BAv4cwVxtl3aInOMnpHoVMtRJ9
gSVW3AZAqjpHtzt/ajj35Mx2pahUvRklG90QeXE8uNgHXDfKWTA9LDS6QyfXq34w
bNIR67yx2KF+PH4CXm6Ld0H5k8IDBTC7mfnZ4bFw+r1I1bYOqVI2OZhPG+srVWEU
D8Xh8mw25+vDQ7CCQJmwtnO4gEU0e/kAv8K/gk5Qfn542GtV13oERwJCoGQkbQcJ
iFQFNi1gByb+0ApqwMvK/RiWLPs/cPCSMqh/Zd8XeQ4v61HR/VHhOUAihvXMzUbl
upzhMTwzD+r57XybYMTibKG6ZNUnwyTWtNwAhn8wVyYxzeUZruZn+oh6TuGA7xjj
Vj5xHkvG2ai0xInd/+uk/cnas18gY3hVrFipyQunt8X9sUUlV3pWzGWh0+xsFruk
4UyoCUZLwB9MY7XZV2AdXvEqA7OVDjI67aXq94UWTQShUcceuxiwHsN4pd5ZxLlv
YIt1waDPbs3Njx+QqovXNn8ZsnXU2rYmZLJ+D+NMFWLVdpqPcY+WblGz6ZCJXKa3
DQMrYnb5b9J0zSV70gWE9ffervvke9BkpkVV3Luf77eCODaB394ajkUyM7VU2OEW
rLSO9G8QyFxDudot5mWpY+UmTsJhgRxlH+LDlI6gp4BAJATsDPu2wES31TyYX3Ui
wyiMxmQ07iAUooreG7RE0AKmNIpKERw0NohZjghkOW9z0JRuShgiO7wMySb/SOXS
Ssl98La9WhBqOcprr4AlxMQjRcqTYIaRXNI4PXOfi3CF9ysM25QWeTUvxqfxhSgu
+LMemJD+kMrz0dH6I2TDydNF5FV6W6LfUcxCbc5AtFjN3V2asAlb7YnAcQK6ueVC
NcrgUzc+P7BPt6WtaniT3W3K7D8YYLhC8v6gUeLRYwNdvvan0IRaj+QjEFCdT5cP
XT7zxaFMhNChhLEU6yTBgQuumlmEYnAIfRlLu8DSZovER7MYrtRMXRG8XWCPsodk
R60HjVaBiq9KfZNd8B+zkMq2YziCzTs0BG2+JVSDXAjk1HHeKbfOm3QxjOObG27I
/ZqEgUmQoUGij6fDnDFyV//1umHs3rml9Q39tGadEf5sNkgTJiIS17jndD9pNpbP
QYOm0GSdpim5wrpiMCxiic/QcBT0zydYrxsJusgtGgi+xBv09D0qzSQTmsZawW1F
C+oKk/CCAHMghaSdwOtaz2G3MC+5FJgw9uT69/v+GswW5B/oiZr/3RD5sHCOv/4z
k5A8OxQsLxl60IMFgBFhAmW3m+n9N9l8nsNvu/yPrOwDpUsCBGM03FcqHXQTr/99
0TRWiUYdv4GMwALBhFLnQdNMpeHkj+En5bHJP+TnwCIyoSRYDKioH2CSCennCemS
q+oC0NrerbD4fNYLg4D/xaZGBB3UyUB9YMiLYLcqk3atSYUUAaksskG/Wi1CTkVP
JJuAp8UrhaHTeLsqIy2QbrnE5ciFwX9JD1DhpOMM/SbjkEda4srfCbs+3v0wXT4p
JfoRYUCMQeIn7jXI+/moMUWtTxF58/G3wd0U9gtiOVqYmcaqMTJwfGmXK28VceKm
7s+6y6ilRP/wS8P7Qe0Zh2ivM87n79DIErH/8A6tOBOOcOWErzuyB0ogN1s/I2aI
woCSzcm+JzbVsC+cyyCd4D4OFk1O19xUcip5pEicL1oyGQ4e79dCQFd8pkFscgRE
nzgC/CTvMkRliKVwUB/jopGjUl+rhL6MOw+OmKoKlrgHHsinmJqMxPlljadT6y1F
pXUsKJwMKlxL6qAayoaeRZZQai9/p4mwp5XMN7iHdZEzxT0BAd2p4c+dJRCYZtTs
06NjAno+aweogAN44hNABF/0Mn4FzQsK8um7HdsQd5ZPPkoYZB86VUmK5wl9CffO
gLVLMn6wnUpFKV/ATvjGIA8qywZJKrop1kTMbFq/IoRdwCs76nbvHvQ9YbpZWieJ
DUHiEwaR63hmnYIOeaqZ7Cj4hpZtjtDVaQwaIgw4UIQvQwTwbe9UqXod6b+9kjZT
cluuf1qiOuCMNyPsRcvPeV/A0N8bof9BOFEec0M5gGPP+a7E9plOrQSotELms/+R
UW5bzsh8JzsMs9C3zp9PS9rav4HJz+Rjo1ze/TsX91IPdLKoWbIuktV1b6613qj+
wtlx4r9YN3xaPmTqFeiW7CuA0nDuZsqQNZP2xOyoVEdTbbre9RqQ63P72YjnW66C
V3K5ZfUwSeTx2lU0KsvhyNNXB6eDyoIA/3eobcJoNoanRcMUimZcaeBhvjZNMWtq
W1yNw4KbtxhxMDy6Vur449FzGPj5gJ0dtgLlpmcO3nGhz4Ij2AUFM58zdMtwWp7o
rRLupsz6p5w23oEGBaJcGygng2a22hjCej3mfDqCyQzultFlNL57v36MU4vL84P/
XA5kJHB4MHMQ2IUd3OBcpr9EajVRhnZk/zz0swwVhFbX/CbMtY/9lO/ukj2X+vl2
k3F873SBDkeAcvaKP4Js7YryLuSo+XhhtTNRbY5Wz++Etwm7wpAwCtCJc9sQX8Y7
FvgoR9rGjgrBDtGf/fDsJzyJuOCM4/MCFNrlrk9MLRugVWaYKR8tCu+gjxStvuRE
EPBEQx56Bfp8pU690CsfxC5tWZuNldGi7EinEMYo8O3/FjUa0p/LRPr7Q3yMzKLj
AoBGwiWAXIkfSeTb3/fYltibiRb7w/+1krAgNRkr5wJ5DC/oMt2OaEyp2rodtzXR
hWGJ8+UHB+FsXyp4O4rt9owCRdUgg+Dcj9XZcLpalNEyEGvef83W9G3bOvzluQLL
z4AaHMajGsHQ7yQd1yItADEiZBwb3d8sa7eOgAd5JHt5aG+oGMCnfu9rXsIuq0XH
dvZh8RlgdCzmViTFLreDiubuQn2yyIUeIkBB2y2E8OHbWKelLzb9UfV4cxqQjhCv
D5Dlg5sAx4hfKZA4+fMC49x4g3ke7T/TbVRytBj6BEuKrWTpVHTbmP1y3GX2SOVv
/Q5nnKEucpev5nkJNAbkyj29ndl3NoOe0JjP07WncxkLlkNTcr6lMu1rXKm6vh99
tf+3PQccSFwRsCa89FwmlMPl5Gtr7R3jwaPCqRMZlrvcG+KqqusgUOND41El4NuL
BfzTOoUXXusrOa5FtdD3WQbasN05o9nlRKbI4CjMNFd06vFpICgbDsGLTbDvLkKH
6BmjVuJKsaSTNGi0noVBXdwm2uJYhtImO61yMQVqKjcG9pm6UhAJu1uI2c/NXRiF
n3TRtJB6nBDkbqIWBgQ4nnowf5uNkCDRaplWY5JQMa7WTZui/VN3L8yAxrAKLAsO
A97mqaNKPq00qgYWWTIeuK+BPRLsZsHFc7DDY9f+rQSCm+8EpNl+O06XGaorxCS9
tXziJCdLcUlAwwJTknMkUMJheMDvKxEi2MPgyT0499uzZriPK/GIBxwfY9HmIziX
f0HWx6ptyZiWOq1cSpFQsP3WokgL2wwFdJQ8JQFgXrWJROrqniYMTjl0dHeIaI1C
c1/n6ITKiDqg/6kr6XPDsz/lYw/IvOLoeqpVbAOz+Sa4N8C7Lemjo+Jy5o5P+4tN
4CnUyRXN3T4A5deyvpD/ra2TD0QObhzSr6Fo13TJ/dfTw4epae7wyKpyQ79y6Lwt
OmxK6Ktg9rPguvWFZz70zhtbNdSOwKyjOhWx3UdD5a+RweLwczinanIiLr9cdK4J
Hi+eIc5h+2AkabvWLtfg4zjhlBYcLAXa1t9q//tXAto0xL5Pgs5mrX/DzRj3yHFk
yKF3e+5JV+s3+fnAcqmXfj5I6BuLZxLrkIqjbpWxSKtL9J5nlw6OoGbCKOl2aRUB
/VrXGlxfxBlfF2KI2hQ2cimg9mzh9E0BWwZb4xPctH4eTH0C6zLeT6DLOVS1tKP9
qM/3DXXN7ieEK4RBtN0y6ziiFahX+VZtK9NJGiClL3usduiiFVg5SmP1q8X8Mf+T
3dXuGLeShUHyrNP7gslUX7GpPzoQL7YRw3tE8Uy3boaY3EuzvUlOYzeZvMNmo5e2
u5FIyDfX4aIzNx/ho9s5WHwrpzewu008uqzAvwFqFiWMZYW94avsw+XAi/mFNPhP
Mhp7uJ+GRvT6Om9XBaelQX0vqjJoNHuQihBaqRUi4WaaFuflFuJ4OLL2EZP2q1ib
1vzUPrR6qGKQfsIqbqgwNviWfxP5NlALM19B12Qes5eUt1Iu5xlXSgeNtLtTCa9w
r+JvUSCWWlUEMZyUq02aBHggnI9W8oD2vrIx5I1IdEFKFwkiUTDLBi/F5Wc6V1AI
JjQeO46AVCGoYWK+1Llr0sDkHX3yzpIHpJsq6cS1G4CUtV6RVA95Rq/UcpveVH+d
46wzltlCpVfKSidgZ0PTBbrOkaSJYk46Osrdebccc0fKyWcMDSG/8QiRlrp8veLW
0jU8uekgrp+bAkxpeNsyU1viKIGd9EZ3LRrPNcYEVQ6DoYkMBdAb1nnpPTFw8+0E
4CpHyOPguZhSZ6BMRiVDoyq/KwKK0aZpS2dwDrPURjFsV+zd7MFRjJTPiwT2qkcl
wh5Whfpzr3OEo9jHEzO/lb8g+um/+ugelAOVTPI4tTzjpfwxl00Qv/tLwG1rJ5m+
N/zlzduqM2D6XrbZNyQ1fRlbR/h+Ge89C0c9FMDb0xIAHfsSafiTVoMob50p41PH
zGrPfJRBJbpnWRs01DTrJyaiOHz9k2NjYDmc4OikA9AZzTmfb2MJ/1J8tuO74Ujl
3BYPTL1aPDqq6vukfhDoxK0E9Qd7KrXQ1skaAij3LmkDLbmxV2NzebEh0wQqo41j
kpnES3HNZfZRFtremNcL02MPy4VekZxhGNDllhbX/K/WZv/vxz0jQvxfkILGVtiT
ipXX/zkGwVQ0b6vG2PA+6acFdjJ3HDVeu/w9cZ2trW8Rf0MNCCI6IbjG7X6pSfCz
dRnBWUi20REgcQNUkcx0gcIHxv2J955AgdapZ8bO2HtTy4aEBPDee6fvybJzZWyn
y9vdh5WH4dKMfMvPBnqduQq1Hsw4RhPABdE82tqDI+mRe5QvqX7YL2+g//IiplqB
9/db5OJlq+nv+x66DaqWPBQkKjVOMk2NdYIC9GOOVFDmCmSzC411InI07vtWs7yd
zgAzfeq08BF7lsW5Fdi/XJFvH9JNh0OnfwLCkEdm6oCZIjqHnabXK4i0vG8UNiEk
NDT+42bwqHAalEKqb+kt/jw6awT1iR8AXqJZZmPbOfjJcOW6nyBswT76/uboZN4Z
lW1fQO5wBkjeGnOrGbS3/Y05eGRe4VS+DxlMxDSztJr+2tg68vDGXhnxcdcIsHRb
We/h3vbDB/yNP2iIRQUTjPZ0NVy/u+4qN2vuOhK2uA2lWdvB72UUs2UYD9zf1AZm
VGQZ9AA4G367c+aOdaDJUWSk5CDArvud1U/C0Mw9zECOPvh52oDv5dby3B/Z+oLr
jRhQp7VpqJQhGaFExRp/PGQ/jRQGdBGcxBXc+Hsx84fqGkxHZj+dQO0a+cbwDw4u
n5ea7TkhmllOd6+KHqIz+oaO7ALWwwN3CbzGaCUK+5Qb7sAC9IXGdYLSSApmNOki
/CXvW420g0jJYIWxomMF5scGRjuMk2igBqX+FyLyr0iD5ZIOb6KEuYcKJJLg8tx8
7rdClpGqtYcCF65ia882/D49rBth1C3CEe/PijiiyhDvIPh0u1G+rjcdcovkOjfa
eehOKXN8GJk2OCC/omBApXII/PPQ5TMDuIipTCov+Eu/Zw4iyjJJb6xsO2EIw8qA
pdVzSEpPOGfpiBcvDdPkuItCBLc7nWhtTmisi1laxKBTYPNPiPhvwVyC//u8ekbb
um1JorZfT85ScFcVBLP1niWzx7rqgU9P5dVr1lEPBrV5KrkwL5wWOusVfqBNhSbm
VeeqjpvQ6nqw75pdcJxLj2n7GibjdDOCFFRou0Rxc5+Vo7QchqZ58DHlc29nyzuM
vJYI7bVCqmvrhFLh652yhncDJjwwaKg5U6Ozi1Mx5zwEbJbj5/yCULQGQ/4vuvKE
R/7N31o/e6O/SMvTsv+dZo3MZTiWFmSmvMgw4CK7hVubvYZRzFYNqk+Agqs3QdBZ
rrAGWadOyBIqXTJqsThT33siny1O/GzE1hupcDLK2oLNSdPqH33PvV9i20TksK54
ekY80k3XnhQakslh20ZSjvTFQDsVtPVJl5gXZFIMrgs9c8Q8PcVIzr2S4kyGIX8I
oxxX1eNqVXvpk34nwvpIFQ1ctW6NGYri5C9ZQMO8DuNY0Zq+ucGBsndyBML31p1s
QjxKwBDU+0ipA3UJaaazeSnZsMj3OtIZ82l0bznJvBM27a+gxXMi5V1J2Bf0RiFU
15cPKrzbgU9z/v+pLYHnu1oA3wCGz+Npy6dn0USAWl/14TsXImjF5pJeh3QxAVaf
zgaPz8XGaw4REuKl8ZWdF4ZFBfF4ph3gdCc3at/IitgFP65TTsT3PYXqofzkl+pM
FBcmUXj1TaqbzsDAoc/lTA1YSd/8R9op0gOUr4DNeccL/ya+K+Qs1HI6aL7uwD7U
XRoHp7RMw/AkPgfqlki5F8wKT5JFcmvmE3c/W+QrRtArhC1H7heRssP5sGEnWb3r
XDibCdpwja6nAjDvXiwWc5vZfj14X14ne9l8WTVHdyWgB9R9jLlSdZpSdvYPEDB0
iV/kV8lhs55mILy1NB8Pe50j8bKVNy3xhL5KAPuoxSOVcX3FnvH10lvB35IdTFyz
C9UTm9Hk7BwmDjCAYZ8czkz5rGWZ6dUOWSHlqJ+sZfs6K56mJxYwW0xN1Kca6rel
oOkt4TbUdhLiJQVkgi/UCShG+Z3/9FXveQ8ClIUB/xJnGe/TyKHYNCckjmHAIB/E
fyoF6aTv+P26LZlDlHlbB25jT5S7Tkox1ZQuZhpgnxUUYh2rWz8XUBzP7pX1rxww
51YXjZDg86SV2Dxy96X9Uv6C6BgesvoNRoBuAnK6TNeFxGQ8B4z60bOcMHCyL0ub
zTfSMWB29bqNelRKphL7p8t7CrE9mXaZmzrNCb8ZlBGxkPduVl2b/59K/kVoEHye
+rs90XPwfquShFpLm3iPbYbE/kbEIDkYEdThYUwcKTwOvjZK8hamW7Ac4Yx66NB2
0k8fviYzxri274vZJukB9nBKQBrt3XfOazu0YxkzfIhJEnB5XSIYSrojg5bE2xjy
EJik6WLSK+0L13LaHbV4UYavnyLG2B0e1HdFmVWhir1m+fDhTyKYW9moT4iyDQj0
6He10dV3sJM0tBUqcs+dKIbR+awftc6x9AP6bFOj1qQhWuslhtw7p6MraTzTny3H
BciJ2ERyEUtJcQ9R6HvaUW2npU9NtJxs3wyXdC+uMz0z6nt1ExnpWm9X23Zlt18Q
loEOm5usoHw7710yrqjLmdRAB5/7fTjuCCWGV7Tl+bJ4xezUmBjbMrtNpq7fjggC
zqA+Hl5AauazYL83OjSJMsCiG5UY2i0fsyZhFsT9Jx5h94X9t6TAlNe6ZxURN/9S
wwfEpBqnxTnvXgCtWiqtON+atgXUuOqLPdWzxUuq3+68r6ygaCHxtUjhpEOKQiu5
bPECn9PLgGc9eNrJXkVcI95axa0VQDW4vxKwBySj4s6l7P1oV62QcS6JIlMc4Ww1
aKnjz0D3PaFEj1beDA/l470ThIwBqBATaCdJSneocJqAuBU9U/1RoM05G+FIDehn
+G+rO6Ynqs5sJZmSsreV4dOYyQyq4Zi20KLVnu52ZSnXTAZV3/I08VcEiwnKpPUt
30bqiu69Yu5E/k2+27ErezkyigQ25dW9JYLsjJaSaUN425BmP/DvnSsynFI5b2FD
+fAdyhVugzCEF8Em5Z4B9A3TMF5A46haWx7eLeWlXvpD4xam8n8k7wPRTz481EsS
u7hZuTJiYiMCNGZthABEc3L3Xx7+CT0HEOAuW1SAZIig2gw6/yIAjbGuzEdAfKus
JJ3A0NJxJf0RISGLPbeWOqoA9vVLPKnaLnJsI+KywM+8V+0cd5LeJMym8+yuts/D
q8VD2siQRd8u+XUBd+PIzOJiDU4uJdJDcN+7e7S7oiOlrwBxtTgocNmvaHK7zsFr
4UUNqr75wmoe2p3oV0yqlXvwIaU8lFwSmN4yuuBU/tdkQgZw+nK58de8LcY/bSAQ
sJ6meGl3canMgXnV9IDghQyCLSeqYy2OXw4o7xqQYziBiUGQShXuGDV1JcYfCOzA
wGssxKxSCQKmMqivF4MS6DSR2EZd8zUuZ6DRKMS+e73tLLjbLcxGAoY1N6vWcx2J
A2qxZpaw95Z7g+FhLyGPygs06kK66LdArYZyNwPP4q9sF/jcHKmlO10EKjWV4cj6
e7+ILXt45slc+S5ihmvB/0uKYWk/brc8PhN+ojwtZN7y6Wr3SFMzydtUvLTqJuHP
+TeMEketxppVbdYCp9TlkyVQZEqiEKgRFClYynjVK/CXpA3C03LLkCty4Pmd2rt/
i6bkkQkt6vP/mUMqcpniuhuBYFNGj6mLvDFijj4mwPLDi2VjKyDK2+zDT7w8Ux2Q
SmV6NHgpldpZ08ISsdnXflU03RsybZvePKfjc+8bSM8qH77FPZgwbCWLmC4JlFY2
ZwYonOv3CNVQwGxaqbBlDHaykvy+VxsDgf65KltSUTT7AnZFnzu4Dpn0lgzXaxso
ma1WT84epw19otF08ctN5j/Fr2AA0KfybhKSbY1z9QMGmzDstPE5SuxUCIcHq6by
y9Ywyj2z9LxwphAderoTgMUbTjBZogeLL9B7K648RYOcB1ipp5JqZYfDtFN3FDLT
VeR5xjx5jDkgi/vtBd+U+dI+WRZGLrHKuVCVaAuYHqH0ZNre+fQdKLlkPeRTfjvJ
ANNfZny1Ejdex7BTwQtGFFDkXIBZXsFssc3ZQ84/kWR4Q9SseED0hCf0ac46cI3j
3Yh7qY5KyrRy7V6SkrXiyBQr4jC0Otfrpk334Z18dBHKp34AVq8IXe+ENnmZ/9dN
IcvXDV5Ke5Rl8dwHt57r7Tv7FIgmhmDjPQ3zEWlCl/nW2amhLtr4ZvoE1JHwm2m9
tU4FnHEjOK/gIcIEbPcH3H1YiBOXea9hr/4ca1EPwIsvcPG5sKaysboGvFlE/OUD
Kb3n13Zcd5m902+ANCVdnTW54O5ip1gHKc37yG1QGSXV+7TKvRH/RWqLK/JOyHCo
gxLNAaKYgGS/QV5uRzEV6FDxXUC31askaQ+IzCicuJftjlAav3PiMkba/13GebTq
y9T9xKYif9VQ5oJMDr27MvJ2vNi3KxPjqaZfjY0i/WpUjsekYILLnPHEOqHAcfoM
CWGuBcOWSkJyE2p8OnDjpoUJqh9Dcp0LhTazXyVTzNW+Q4ysRjTVg8bafu8j/BZp
HKFjWlFe2fH2m3wyah4AbUk0bR+GIdUz3RH4V6q73c4E4IklNhPGQICsyEpckDxj
fp52JIFFstB3B/9QDrVXEqYtlZClwbJ4XhkFwZW74rPwijrsPigJ4cdS6g2EinLL
macYPav9USayKfxQhZXImSq3qEpVX1hCdVZD2VKXH2BEiT8rs7c7ht1W0Sx7jt8N
c2JpzrkRUkesrlee1LGK2pKwZOuB8lce9zCL8m4f31wAn3h0i098sE8xDU8Njcwq
iCJh3bQYk5fxPHfYJVCvbuJ+equi0Ju7D+26KNbz/3qjl8wxyWAaJP2f39QNyGON
L8L/usKiHuBsaxmNH3JXg1CnO5vbDNuNa774dUodmRssmT8MTQSelMXwgw3DjT1b
SG05Z4J+Pa4SUcRRwxsN7NeBsxozBUguBUGnUzVOwaXyxGQqll80kHSQ2eqvGslj
M6z/j5izTKSwvRj2gwwcXU3rlgYjYAIeU3NmlhU0L4/YXCYONUy8GXNTjAY9HYvY
uep8XtT7tCxGcEVdjDPD96xmPKxwjKt04HV6v0KgZDA83/ZUk9BsEZpx5T4vYdRN
XYsUhZGo65+vKVEpmTgnhQQBR0guWxhcC2+e6iByeKgjE3C2yLaR8NLwxA1A9teL
NkMy+LdB9RKYccTDaY//rJUNMqxe+lkwK8GpepOQxi6orBu9kj/mB5MFxVwrEAaN
+CNGOmr/rCz9M04c9WHeYXwLWkAo0KZa9DF8/4Zn6/7/CIQlSyizffY/+U//roGI
P2afJPornwCXYvq041hNTFCuMISdLb4lyR/Ff61uPglk67do7qgYeQbVhYov55+8
pbwLvNwuycLR+A12Bk6QSWtO74jmewaWy64TibiBuyZ06yEq0MYJaJvpPnbAl/Wx
o6h87XXlBrn5OeNcWGPELq9dpXox0qd0VARCwKls2HhX9fre6hGg+B6sHHBrMtvh
gIBPZpzBEcCBlbH4bGpw4V5nXGi8VOxfgUdEax/6yMeFJ6Sm5w9zh09V/RJNS4ZD
HfYv1ONq8lpkQ/bAIQUJSKc5SxDCXHOccpc5QDHmOlnxL4uhnGjz/oAAJRqcJqeE
BP8jcMXtREhRJY7LPevT3fy3d8viktbZw2Ll65Q3zy9s7L/bVjfu8WMXbb90P1UY
KQyDl9FGXEUPT3nbpMvtsdOhykOV6aLS3rvQM846/sJW1h4t/ZDQXv+90cp0ohLG
6hVIeISXslyDfEb6i25LKbUp/uey+1I4IxcWHRGk8VgzE4p7+8dJN4WVDEHWLsXI
cZk0lbl8zKfGoO0QezAeJp7kB7zHwfiXmA8hXX51cGd18ALfeajavIAcb8ZaEjSq
TdrBnwXSj0McCIscSj+344UAcO3DFxkeQisMniYiGeRUoVm1S5TbglY/kKygxhb4
LZaO9niY5FPX1QjLk71yWOZNJ/hYQRcyAsBCHUFkEKh2fsOdpirPnawkQjmixU61
9fCMyE8mAFAliM45UXUA++84OoESnDmu3UYdFZ8cCNtgmB3YVfAOSFTn0i+M7VFw
7RTMAbmMkXePuu4Q2kohIGNRwGE3V5dE/wgAgu2jtJePf1dnf/AA/b3zQ5HUhorH
NGcwEI0JwFKTHe2dzgOL79TAOY1q3+g1NUJmuWM2EdeG0ow4uYq3GLLq0om3F+WB
ujlbEabBw1POOp3i10gQJj/oRcST/xMnAMqhsft+G42r1hboLljCs4j+EHTP5LPm
xj7IyElrALxrfqhYMvQef5jADSW6iT/OOlIcmIme7N9UjGxCzPNuAG1oxHUM/yQN
1FSaQCJQroACPSBmsELOe61mA2o72HUaBiU/JHb1bJSQ8sJA09vN6oP9vR44U5ps
vUII3ETRBen4nWLeObXwwv2VAhaHRdOpzFVtWjj4Kb7HwiisB+BOH/hMzF2XNRF0
vE3epKDM+ceJC6vbD479QWgeupCAasjTnmCvQyI03a1sys3+/eN1KO2dbe47OQIx
0NdeY3blsN2ctcN9kYOFFAtl7d/zvcrtaFu+zwr+sV507ucTcCDsTSO2+kkxneHu
V3ZauO3cYbcoWKXyOTm7OrmeRWR7qcrfn01CO/TM6eIwc/wHlDLmjACjLUeqHclt
5IUbY2xqqv8AcAn78uFaQyX69lxlzLXgjx6TSQ/0Z2VWfCVg5eYSlObsdTub/wa7
9W/WUjUD7D9nwzrBGCXWJ/JDtdFDyOilpih/pEZjCuY2N5uxKlzHEGy74WQlDHzf
HnTmBRPZ2Y9WpvJrisg95SEZTKby0Juup+Cs+6Sr3Mnj+CzsUqDN+hi6ByL50WMp
guXC68mFPhv+CNIlbTxVmh9kLdH7tzojnPplzaQ2NqKJIBtslhDnk6WbrtAPWXII
lnXilc4g4RBtoTeuBltAsy/Z+7V7eQAHsT4FEOaTQtVCcBJ+lAaoLx1xolTW7FTG
xifRVjLwmOfE6BsjlwGafm+UzapW4NYdexajxWtLwwQkCOF/Z7YUeRZ3FUBXydJq
iokFLSyzbQ3yUoxhr6eOWK54WRpjCYs0MrwIaPk92AIlfekDRCaCEfgRPODw3IkB
RaWk0/C6W1KT4GsA6F47h/u0VS59OS2ocTocv8z9Xd/EONF5oxqrRPgi7vfEPaW/
6yANS3cnVHy/1ckNQvf/zvdQ9fYKWZe61IVWhS9gYF2zJH+XqOiYDcG6++wa7W7C
Ly0L/QLc0EeXUWG2JHXUc9JBKWrdKWXOX8gYLZSAaB47cFyhDqp5OOEHWZQm9PqW
Y7taOWz7/4B8cdSaIdQf9GdJ/18BrnbJOhjTDh3+vmMpRG6QtlsrHOmfwLCsf1yL
Bt0lekxi/X+7MNNf8RLUu5AzhwGtlXz62wih5ugBJv3m7hJLQtEvTJpJ54ew4aJ4
GEwX8yVMMSRyLk54OVqXj3vO6TMghg/AKO8Z1S3Csx+bMOgB23XIhdvO5WrFQuGP
4WcO6Hg5PhTM//1VoO9MwbUuIzMkQhqtQ7+SGiHplcPxRS7xRWRDrvd8SnpOe28S
uKqf/HX4uy3/ChK5kKuSWvtYVfkQnHu8jHLB3TOb1fIma6+1V6rHHSuK8/Y1prz/
DBkkNbBQ2xySBkA5CKbCPuH4GQxzbNDvd2y/E9U/JxAUhrIbnvFMNWmlfZbwTgJ6
Pg20WQ9Fc33qIfGVpW1Ylo8JEDe+PUooOV4Sn56o93EV6pJCdi05spfaAAjR5Yxv
zf3SS4xNd5VO+6oFUd3wpybl3cizNKgzwKHla+GMFKIeZqfL20PDG87RtPUec1b0
E/DW3AyvbysmtcOEgCHIm8vLqksG+108vTj1EgMS7RCknffsEaI3DhLRC90PUjEM
yhjXIM33ub+ctb9ZkD5SDni5CIiQBL9VQXud9yOfWUroRIjVeg3H/m09DGrIDzLA
mIzLfywUjwvcRAKMBSiKeVq9Ec17FMGjA7JGmiQA0RmQemmbi7VHcMp1TXtsk4xq
hvjF+GL3m9TMh1wwSmwi3CZr8a5F7F/E9JOiHvzWHiUcO2NxWqZwCAMC/xp26RJ4
pyBhEOJ1PjhMoYR0/mBSDV3FAt8SwDsaKjGnQVLP4TVMMC/F9KbjimQ3sdyuSAA5
k4bCdzCqeydj3cv2ZAPJ/ekOS2ghETdILedGOW3f7GNzo2E+LMrt6sFMr1W6Ppja
eKQwbjVI0zX9utWjPwi+doNY2N2H/yEL6/A5ywww0fb4SJZ3qhuAiCKaCMq/iGGq
66dWhE2cEkgHtFZyXdcUko/I29iolqWsWGIiaLAXKX+vgJUSvmGj+sxnd22rywjz
J3jJTBmsdQOq9a8YfZpSycILBeqzm9OZGMxrTuTUxgEdtRcmfiPYK7ykGKO1Boxs
Vojmx9cTiaqdFOHUeh+Shbd0vWp6KSgQgQGugWaU1N1FUcxSoTrZk3aaedM8jQlJ
frrecp3uHSC1n0Am+qiwLs9KpqT5NxDp6wBzVwqFBWx4yfTvVQ2gPu6jXlgBe3qr
/dUjClOkTqTjNmaya64xEQeJty/L0JjAICtSbHmPDPND9ySEXjrIu5JG2QQKogZI
FLmFURN9UhKtgF6arGspgFqA/BbkPP8QCJi9/ImrfzR7vaSxdV4ZfBGWaBqpluoE
o7mdZ89MTWGQT9EQ3Zsn1jOiJOOZCuupYHXOPv4zWAFzWxbQV0EhBKuPxr9+iZGy
UHF0H7XPLz//oXlAG0EZ3HDJvwLDsatOxcQVpGvJAO+cVxlQhNJ4l1ed4WneZXbz
0a3buENQI8MtSFD0D9t4KZ/8EcAIDmte8e1L5pnhKcdUIauPhKu7HzsKzOf8jjb6
bAs3Hf11+IEis8KFdXoYc9aWOmd/3GQk58TBm6Uks9NF5f7QNR/EXgkVmOwat0rO
kwgW80DN0vQBPQ189IQmt+GEAZN2xRN3ESdQsrjTydb4vfleSdcFY//Cf+obzQ21
pp1MGOymPrQ8PfBgpjwjEvCg3CSZrkEwpYuQE3nKHkWtlHf7Aq5SQgpTzIV8yVcs
7TRzxKtFlglfrjgN5y/Yq2aZYzAvVavyIBE3KQheGMORd1k/DXC4sU3M7SCamee6
ksqcYfxcZ56+h6AFryrJY3TIT6p7WD2oXjgsJNB/zn5xBW22bqaFEkB0g5lFcCSy
bb3e51k66QBaa+zfIDU6QeARpfyA/fSGJgM3ZKDG+NuVyZ1/t6XTVAT11i9YGW6J
8wGCwKlGP18LXa+NvnoBHz0meHUZk+6RpRTZ0CKxA4dS9QxG/3lgT0vlUJSlsSRF
eGgRIIipHz2JEJp+mPRBQpIASSFCj3pL99kXG66MwqQO3HbaKEIW71aH9z0/azLC
UgbQxdhxuQ8WS0hZXiup8cHJ6erw7vksMRPjvjKy9wnXm7W9osr4Uc645Ax0lkI0
G0KKqGGDu6XrzEfeuGqJiwn5El5zc2FsO20iQXgJlzMhJd4vMyvrj9I1n2bSPgWR
s+E5jez3Oz1oD9xDxSCktbw/2ofzMRgUoZGcSKTgJZnq0c9iDTnrcCy3//we/KOt
IsSEmJeSlz4QfZdw8bLxbOJAkdDXoj2///WMlk/3UCyT+Wnd3Dpa+3C75f+eE2G0
0ytOdvFmcQh/lJrRk7NlJ8U93e1RgdhbW3X2kJHLtwF/94XH7SHs5cVsdpBlRYMw
0M9HsL4EDsSQTElIBv+f5328eP+GJSysPNzczKjS5Btf1k+le9X1tzyurMTou4UJ
zNPvDnz50dYQdoZWPC1kZ25AiDNBJk6N8MXf73lVG0fHxRjYyFX8V/UCNS0xjSMt
ktu5CyihaKT8YonyB8/CGcFSR+NgJ+ftOjBhT6ODHYlcd1VsxXGmSYdWVeCi9qJT
jWKJjWXk+MtqtZ2T7fAO+YIHRyw5wtUnCnWjn7QeHiYEEkLkVKNKLCaOwUBWm8fs
WX/Ijbkjty/GvVWpAzdJw0n+NtqR9zBc1gtRmYMGKSAAYyHkK4IyvLEN/65w8UKl
aGlJsni0I3GukUC9AX6OCZ3xHPhYaI4w5+3qjO7VyTIHgiC7vNFIwLC2y2j9+Cy2
KCSgap+9ucCTmpifKAVk+jOqiMl1Et7dBst+/VztxHEvABav9N1h31UAuSxB4FEx
cI9fnv0Zq3xBNOZBdIFeVlMW/d3TgBgSYV9WZCNp6gMrU1SY6bpjGAuTi1i4dTv3
5J1h0WlH/BTn3Q/C+g+b9p9yntZbpMGNfhhcOHwbS+P7iDxpn+AQCsFxdiSJhpBw
C9IUZyaDzxCTpD70lzm3ylBY0jUYNyC+Kc+b5cAxugahn5bAkmLJ+tSYE9Swm1nS
NORH0xyfedP1NtagJUHiy1SGU9bVsm3RCVX57PZ5q6+donYk4ZPw34iH6sZ76bXy
3KndmLHLbRbfpavrtroVBx2+2UHExdJH89IWuwzcErafta5M15EOMH5mTBDjgTTX
dRHaqN4Vzgta96Az+wE7GDiz+lbxba9g2UdyRuzC+rJduooCOrcysdaS9dNZzk7+
uc8QSOouJUN8ifL4pxH6wLX3Sg/1AdsrHuQg59UR8FBigFACBtiPc0TEmZZwTTze
cCIlXErOJ1OFwEYn104uZbYQlw3Gl8VMv9yUJVyVd29PMiPGS/1qIdnGvCWUN/0j
ph1odGPLCqCMP0vS2vfZ5RRWxlZay49VFDcWcdR3Bw6IjrwQuqBF/ihRpHwaHqsh
bIQCP4lg/Ab4gqAStOCp9Vb3oKtn92msMUJIamvzx+1dE3N1b0iVgsvM3xZs4N/4
qJXLw0TQ8Ci6uPCB0SZYHzzU/rutRtdz1fK1oH2MyGAnOssE5wTv9lhuPWjfDBPa
8R/yivr2Tn942VFAw9F9ENudgFSBs1PJ+sZO/v2nYP3LXIRn9FX50sh/ygZLvzKU
MXcPqD+TLtpf6y/D8AbzQt6KZdrk2Wj21HHNxXBHE6zr0pkjCyHx1keu05BcMqdn
b+wOoXKILtfMVZVFnB5ItobbNBhRQL0LsdZ5Fhq1DkLTqCBzsEZpk9+xxq1N+n5U
W2LNsjdNZyj6sYFh9knXsgTZOpWkVy+6/o5ajv2C50o1Q0j0DI3t8rlWOmXBkyHF
flt2F1XOQXL9bKjTIVDVGf9VeIJkgzQLW5ce+0/6FLPDIMqatyeC7PFvbzI1utFm
o8UqijYECmvYlEVkGy7q6KKl1/vdHl2xD5Mm7grLEw1Z4zJ2QtV1eFzUMUMzxq2A
r73RJk4lUYZBewDzU/Fd1+Om3QabAuvLKS18XMa5NamhdnF9U9invo7R3dSTgMfn
/eQolfY7SVSgoNDkznxctAAMhUke6sVbTDKYzjGghH+/Jt8ebXB0mMdtgSwcmnvi
QZXzPHwrg0B53YPPnNP5duWdsf7QAfx3v2yC80irclNwUEWUwmYu/tyWtyFHZpr2
5MzUKKUpW/j5/4Rebw8+GfuFeOzrKVZKaZ/VGVDLUkgBexuKiY3/YB9jiIk0kF9a
xsZjH+RfFCL8G+yVioD2gbkZyEIY6FUBPc7B2W8rMMPrEDOA8+2M2nvh/a6io73X
LJTDkughGi1E7sMpHdHzRTJ1maUZaFgTcvOpiOLKcW9QOmhBuj89OfUa/K9IXtHz
eeF9jGnC9cT6WhVg6l4WCoh9NFBNQpsK6Ge8Wg+C45oCj31RTuhrZasdj7n/EEiQ
VwZkEfPhGc0YgIT0nwycLclMZeVRvjqn6dB8YFPGEAd8EIPysVF0KtEbPV03Vrb2
+Gz+xwp+2ddOQMVBTZilpvAW6E9neppOx61xlZhZDrHPB5m9K177grYK62xCp8Xj
AZ9bxk/jqWnziO1bHn/O7J5Am/tSMuiCksTu5MNlv9t1DHL8kxT6kJdyK22yuGxh
4pX9quDnahIobRupT1zqxshbVIhXPAYMnXpAYHEVy3u74VlH9CrpVqGJccrQBjcT
qDlF/jzUKXrY4c9KV4tKYkmaS06St9TfanM01kpWCDRflHJOpMwaXamjszaxGcF4
AnDmreYczuMYJpPhV8TA1t8Ij8uUGXq9BahjpcthH7miP3gRgvvGSiDrphVkLSXv
U/R7XL0+l5DzpdcWaxLSMFS5wn49h14747lZk/gw5G6AGUeuHXd70FRH421LjPX0
DFb49buRprdOWmRqzQKQVXw8GHKigcWnLh4uBi6p69mgOvClNTjMYzBsFn+1Rem+
SnNJCEO6Q4duyBqU4sQnbyPRYtGo6F4v5Vdv3QDacdQq4W9saQ/Y2jwHzuS26ApB
pvQyUI/0/30psHlvbOk3MPL/G6uOYEuZzy+8O23XmcDCw93+D9F6AWTYirnkkNUT
S96Sqlp7cyE0cJZw3YlXAty/cCOcIJYOVWQbzeVj9qV16rs+FyT4e31GfeEVgf/L
eJ7pb2udkjPTZ97Ul4DmXFJP5WmCIh2o1yTcCRxG4w8spxUpv/h9NoXY46jIV877
weFShZf7pm6MJrmosQuKqLInpu4YKgBMyFIU8rHXuGaGazvJwwTzGAcqZU66592L
aEwX/61g4CxMKtGiyY0LIFDdzPuhNylQPizadKLRwyLBOv8r0DryHEEmG+ekmWV3
0qnF3qcxB8GAKGWJPYWiHddkpnx4pabVyX8/Hm1t2fd7klkR6YG32bx8WWM5e8XJ
POyI1+9uSs8XSFnx1qSqYgDc1psnzxBtj8kxyud4lnjWjurXNI69XQONWJcYTv+s
v77Hb3NyVQzk+/J47cv8NHuFSNdxeD7amuMWbMu+uE5MxdbbM9cbKyuX1V6JkMPg
yHkubnTquBL5wta18Ss6LReCGJ1XuHpW5YOeeuCp1YbL/3q87GTn0gBmyo1ULKqK
CjTsvywyLS0heZd7XR/q47801BJvyYwHJ5gyamlf8EUu6LTfD4LuuSMN9Lj+b8QA
mfAc+MkfOzH5cw/NdrZFXtkuFIOuCtN3Ba68JbvFmOZ0BcTa19PApeegYwCFkwnH
ErLHiOFCc4MMjI4DjDzOl4wxop7xQrc3MJI/LCeD5wrMq/jQFPvYRpoJycLNRPPn
MIhxqWAh/FmYKVZMPPexGscxbSit4OF2suNsPYkTxJPgMMZ9PhCm8ICEQEVGHSPB
XeXzHaXEpo/omc8yia6BVzSNbNDiPG2p61YNuwunH3zctTo3GkqnKcnsF6NEv6rA
R6NWMUuw3CpolvUpxYSBF5DzgleC69z8qvkjKb13aoovYkEQLFWW9Kwge4MuRW7z
N7HQNiu2K4G/wGngha6A8TAXHiYq2KPDw/F4Wf76C2sCmgtT5GOe8rOZZfc+aGTm
qdNlepAU+09bdm9C+MG8leQoQM0tiK3l8mV8evymKOy2Rr+ui7r1TgmZCKp7QdTT
9i2TavHZDUXV4uugtvOG+2Zi89ZDfSHwMeqMmb/fqTpoCyx/alW9t5UZvn3efKYw
wbegDzytSz4YC7xeBzJ4Hy7tIlKRQb/V+YOUHh0EgxyR/b6vQ3zAuWhN2OLP/jD6
SHTQLss2bErFOuinI8f3Xk8u1vOxcO0IPep11ekxXMnwPmywzM5xoPE0e3t1sqis
6MeAEH1XAZeuFMbHlLsl76Ol+XrMqorRpyXrxMaXeij4B3l6xtInRHHVDUEwm1P7
RChRcIUuNUadnwAyGKKOs9BceQ3bymPnSGOW1P5b4LEKp2vJHJSD46sG/fHDwthg
Kal1vJ+LXE1EFFZ6SJdfgeiAOPh/EiUpOAKJKqoeFnPWQOm/LfZT6YGcyjoqG/is
NfvFKKepcm0GJP6BnNYOxN0IWS9X7kPcT5ejmR8oqPtZffFxmC+pWWnwVhOga+v3
2fuYyEK0Wfp3bJvaNDoqrOmUGoYrJLt0AboWg3a3p2Nb/4vgTTgN2T3TVS7HaEBm
WlgjN16+nKao1l8uvbybNRKGnpgQVP4rc1zlTDaG7/LWgFb/ofiAeyJ4QtSyQfCe
NLLi0jYTSB+tyPc5vqTJQc3ee+ZzI+9wsY1rxDTHg+ITDgPEqVN1ywIDf7guFOk4
4oXDy2DwVwFN3KUclLSp3WboRwxpDtKYXgmSKqDbaIGO6O8RC5C3EQjLq169AUtu
S6vXpDsEahBZ3MYgVtwhytnZpshsMOqWaXHW7pqTCL3Ir8AuKxAu4EBSifwEKJHY
OzuFz2aP1SMiZI7zyBwVzUv8eB1pjA+/9lD2s9HLhXhZJs6qLiF17gVl29zS1bJu
duzPBNNg7/OAmhYump8j4tLaTzwt4XqJUI28u8zf+d1BlyLIwdq+euHZHH9FcSPB
6zsbnRvvxAI6bSrwWy8mZgDHa37GC5lDFMBRtbsFnlrFZI9vdnMqOzwJma7hDv11
/tolhCL1vRZYq2lfruNOQSW90TXbmfmLZjfIVAI7FjJQ1P/BJv1pmKpAqJimYWv5
pilU1SZ88mWyjtl1X7/kQ6ryOdI1lYLavW3ijpmK03Px/pDwfeU2WM/OcsGq7icB
JKJyOMFKgOVxW6YaPgroGxkMSktuU2kr+kMIUiHaxBhOlVrplnl1fMIRl6bVaHyM
KSrZpJowkS5rzqmlaG2tiWd3BXLOLHWpIX793Vuj8AtGBUBGe6ja0GRKtcYzqKcB
6mI4VdqpbVmTDRPjtgoEJbAlyhMrPPbU8jstW7ZwkZRXTmJdTBzto7bkRzcA3d21
SYZa9K2u7rL+6RA2L/RafT3aU6e91vdaZesBUtP+qa8BQ9A1e3TG11xWZGJrdZgW
F3SscDzjFsAp1tFtnpM3ss8cCk06j8udePq6ApZidgXgKMf1oWFo/Bv2OgHK4eu0
1EepZMZs9fAGQSCz4LTLopR34c4KF3wil0wDzYJMRjVfaGET0IxLDW4hvXphrJSW
vDzqVCXZNp0e6fZP5ByJCl3rH/YLViqK3312L5v5CR3+ElQ6PtKuXSPoKSy1wXeB
bEOBntoxX7OgsdIlTul7hABrejjIo8IqkmXCnz/xZ/JcoFZWnjYnzZuC9qLhSDoG
i4nXL4vDrUWy/23x3Trdpl5fApIt0hODF3M+CGJbF17D8B7BpFWLtboCPtLdwvM1
7qZML15pde9wUVBb+lL4UjABHY1/o3eUoYDKnYZAyKxTKfOe3+JcUuTpaqSnMkEJ
eAvkQSGBi0XyR/MRKkuVen1iaqTUYLtd9ZdUzWpJ1pyynnibbIkqmlT5SaLO1Ymr
ZpGceOz5P80bZsBaSLsUF1bcp65q/bVQkOJDiR5g1hPLT3/bhWji7LEJ/5V+kiY+
AT/sTuT1FOHqKQc3klLS4TkmQZmED8Y7mHmdqp1PDJhbxZSv6ds2hjjR2DWuhLVU
YwHdNl5/tGa01rhn34CbPuZk+f07qmWYRP8UNX8MwT82egtt2xNWJGYjRsCOTgDj
Sg5x0O5+jxtzRgGfd8ryILqg/5I7Q6vMEbYWqR03Z8xGvx36vQ7Q3CeZNE2lj4Gm
hkDJAJYf/WqmvbYdezPpb9aj80sVi6buNstmFFrlRBAOMZTpxR3pszCy3fGwvcKq
PwtkW8IQ1j96TsuYFPGU0SQKTImKNTEgZr0u+kp5JiNjS/HTGn82DvgFKQEA5AHE
8q2ORibwTAeIq01PQ2S9tcPDyMMCVcBzD81LtMqJzqVno7LJ5bPqDtt7K6Pt8hH5
KL9yB7vtCvdNkbL1dClyynpPyHnxcJXAP9gyHsrCsScn/CzfKpyudYxHcWr2tFCs
xH+/BRl4XNK2uA2ccP9XXFcvFfRm+uvr1g6UhYfDVTlMi1ZE+KRj17Q0yKH9Rq4K
v19LOMvVbUXw0aw05wwPotUJgDUc5FJkyZBV4K5VLq5CJ3KNk8qSRLAoDFX5eHIY
v0dCUS3kF/GJ8v5IrLI8Z/tc6OOJuQWbvww5oCUAa+YU7jy8oD5tcktShLcrZ29r
v20pLQf2qGbxYJ5Yze22PuH/akBLAh8X5DiooXcvpL3nS0LdN629YzsDvDPCe/8g
q8C6Q90rFxD1eoUEhBzGNPltX4ExOXm0Sfvk/eCHTW08iH00bntz3mIzVP/qpK8g
mjGj3TIBNR7ch5C1WjunDI2P1h+QCh5vjHrdXqNKlfTRpJEv6Ig+Vjej1+oVX14B
Kp4AS1QwQ8E62ZhheDrOYLFH4d5TG1GiS+wvFELjBlNZKo8YeI5nrgOLJdQW/SdR
x+sWUv2V+wzfOr0qRtt1GgC//1soohuuAw7V4m/xQDGOqQWQyxRMWuCVVSHk9qq9
JMrmixdkUw1oMbF+PG1MWMvg+84Z3fiC/u3awITa7WH6SzQM3dPzUufAi7YaB+nw
9Ex0+EPcMcwBkql5XI6BCth7b1N4SGYMTaGbIc2Mi8lO2+fUk3WtpA+LH5Khy62v
Fmv/JWaS2N6yPpDtyrXzMOp81Q2AgApconcIfUoIjnKgLG5QXvAQw+z7Slfu7tOw
mZbuvLIV0pJ/0OfI7KerNtfxyEEyTPFy9P9dfT3/Dt+MZyVZ8g/F7qeunXwI8B+e
7BZx/qrWjBkzJK7gEO9ZaMvQ5Pc/ofDsFutXWuPlJIU2SRLtj0xr08spximRn2oD
R7hW1BIRLAAmrY+c15uKaXnHUn5eRxVPa8uT3n9BibjMsdcKL68r+QP8gl7ES6uA
zdchJb3Wn++mUFvUKpU0chQs/a4JDrrTVtT+FxCkwCNDqzr2XkGM346Fw+C+79Uj
7i5KInJs58F+irXoKVdYp7xRgdfVK6MeqMFkgB1T4nfzrmkCzWvPI2+P69YKPCGy
dM9tw4kLjD0ch6js8igDJAujHpOKjCPnpPM2jQUbherzneuWtescPRPAQcEMHPar
wZuP4aSXeQz/b7JkHDLhVScgU5ZXDBUNNUxGAZvLwhl2jBpm0SekinxD7qj355Cy
MP3rniKbYdDX1iRjQ2yOk+8zXMJit5eNR4m2OluygIlWobBL5cgzu4PHXyymcQCB
1EiUV9X/hrfvG9iJj543uZieZvsoUND8v0dAUNyqWm6FCPbS+yMS6P23eDwO7IRA
+c8RxmdqsDiHVt5sNWLcPXkXCiN35MrOn5Jssxn84cLbAyF9j2xYkt02DeuZACwT
JWBdBQI+RhtTI5tF7EKpLdOr7eZf/U6P713bvAH7TliUx+mHZJ11L96XL/LGCEj4
RCJkddYZc5xFj1XVczUUCsT11MpQfitCAn57vO9CjSDuvcGHbVLCEbQGFboO1SUV
fZMQGwp5xmrVpJF1+gHGLS/ljfNfxgdI84206Bpk5SsTaNsPFuX7EAjvki7aazkm
JLVle3YUPqHg6IHk971cRE14VxDK06Ot3oxOPfosJDCsWix9hBchZIV22a6a9QTB
u76iiJ0WcQGPaFMJ/Lc5WqHm5+oZBLdLnl8z6tRydXGzfqWSqspuuRCvk3oojiem
L236OQerqR42u3cm5p0ReN3SfYAOlM6+lWV+3o/z2gaaOfZzlx2VDp+Agves640E
LTr/3+coX4E08fAC51aAKZ6H4Vnz1YdVHvggH87uPeFzVpJKrMNIYuKV8T1Q5eVA
ruvMqm0De4jRWRJgAbNM/i/rJ60KaIFMZMrx0zV8aa5iWZ44SAAkmrlv3qtTjVNS
1xVPTaRkEPWb3sM2BW0bn+RBkvI3IATferWsrPxky0eqXxCaVDa0DUmb47kOghwx
o2mmKdTn7DD22O9sRRaCjZKkQlacS7k60giLS7QtvScmXomz5Y1euWLCG1uzO/kE
Ph5kY/OTon6IapSYwtBdNaWW4C3720X4eUsQyi9hu+eFBa+XkxYgy7n3wVsVuAe8
qnyCa1LjUO2ES2opR/yiOh43m06r5Sz/E6KM6qnW17IV58sUnQzmMyU60kwHV9Vn
Jxrqk29u3DXWEl7YbQdZoyASyz+AqGniC9AP6LBzhyKqDoEc+mcGPZQgP2M1O5uA
pqNuqh6zBfjYTYPnLP89G7eGeEjcnbvaX302oOxlEgThEKbORxWDEgcDGD5hLd9a
1e+9EQCUc4LYm8ilra1AQ/czKiVpnCgan/E/rhHTKIQMz5KQsCfgbfTlEhwJRs4b
fVfXOQAhtEYIFJnKmZHDLGoNZdyoDHT0nz8S8MfQb1Q6JUUau/sPGqzuDNecuUz3
MN8wDB7KeyeVJeqvOy4FO8uRjtUqgorPKrO9WfShOHdzVIAbzqrc8dnRmqhqjuli
nEU5kSDoo/whXNhFOrqXOWA3RliGZBgBUSqYhmypZ1kunNJWvl5P2NAyFaMQ+CdY
YfinLc0IOt2hTe5cj677U8BJEDmlYalurfJGOIi+n0wtTKuzKrwf38DyyrxykKiq
nqKi9ZGIuUrUevefK6sh/EX4HehmlY9+c9iWpBZWPud6HLUAOHVjlENzNtni2itt
wGJnKt5Qyz9Kvyn+nVQ+NBrzT8d5+IyESqt59ZjZ31rofoOKNlZpPgRh7oCdGugP
2/uAFBILbTZ3ggRri3TbwYV66fxDamwdw1FNWJdAJtrKGoazKIzEUYwxkhnqxuld
FZcl7Z8Zv5gio22ngyVJbGpMAsIvKTHEaMWFHnkAPjg0UuZFa+2QwhUIOkzWFEoX
27K7wQaDg8yJaGutDdBKIdfVq1tu2kPtpYrG3Ke5k7l81q9uJUV0bdwS+Bf7rBQE
Erfa8AvlilaDnNT61381g3G8JDcDMQtQtYIH9VmNbsaiKQzw1aJY+XxYdjaxC3sc
b8dVaYDLLohuFfG8s4oz7EGpjZJp06r1bdQr03ltQoC4+isntrjs+MAvAYKdFMTp
bpHgyl+VrH4VObNc8H4l3c6V1B0OgJpB26lyUHxgUXVAeTKjMNZ7ho2B4tShDM87
evslB1cnzwpupkUPrdrSbLFji0cXmcTYgDAhYy0aKP1COZFTjfDX5mj8ncGl/Jj2
cXuDiYFd6OZfXkBn4kq0PiVjs5LgsMl33OCHP2MBQnuMToOckwVWar2Yo9Xe7q9I
S9xPSXGaOgXDoBU0/v5vRz6R/pjT3IvMq3vEgPT4pC/VxrwA8ySeolTRuO2VIXyZ
bK+NejIOTW8rMlVSPuZeAMMLgrZ4nfDN8fE1S60/rEwgLdnc/Ayc8ogZn65phRPs
Fo6pyV2xDf7DtTjwZ7C6wM0GQDccrhNwTA95gp1wWiRaIJwjhpGidxAScBEyNoNl
ddMw0nq8p80oCSOzi8vLfWxaP36kZAQ+fmal5y7eMz2QjgI9ACZewIJbbWvk5E9z
jXxN9bX/ddyKWkpjMQX3ON+x7r0grgTca0Xi7ycDMEQnqVPAKzvzr/1S3JgX0eXK
AnTC9h0o5uto6rC8goiwNAw8Ob2VEhw1ZmdE8kUF5wW/mO1VbhUUIXKurfIGpBn5
7dvC9lP9BT3KjJ7UNAG6gL10JPMwb6rUTlLhHxx24kPWbCv1ZyvZGFZaQ5Acg1Gj
Fc8Zunh5uwL+vb9hMTluokCSvT5CliVBgEHNhFGITY9EF8RSIcXPRxFaJPj2VeoK
llzs38klWjSYmV7wlqGYndfCwcBmKYv3/29yGWX3/h9u8VlHcvH3CJes2cbroZVV
86M3ZiGryd0tR+af9oMdn92YlBJig2YniZ6EypClxk5W6iQIYzqsed23u4qMtu1l
bQ5id/uq8YmAz2We3mrZWVEdjF6fAAswp5/m7tTsMl044mhZgZLUQluSNjBG1wAM
bUzP3FsyioR8PNwICmUL+hzuQ3GCznCAO0J5nCQ6vucrHiJ52UfTzCNQNsUYfLG3
h2CTa4mUOkKgCZl7VhsQ9GEUO5+k7ih8NfIelp+SKuoebsB6wWLmzyv6FmT+f/MX
pGF8O9QXOuJMWAn6mPlydHwlBAuuM3PPdRHAskgIbirUKl9sU4t2f7/JexyhbFOa
xewNZoJBYbNFZ3pn16ghbk3ifRpvMZff+IM8r4U6XnkjE7YAmxZwjTpo+6+qNJfh
R9WbzWjtOrZILcRXGGbIuNy7PA3BEd/kzH6O0FSm7uMbaj8MJpiuz0cEqxsz/Nbf
URdRiX4ifrk8wVr7XqnbBwrRu4dbGhkUgBJsMMrs/1qeypEdipupcQERlcmYNO+S
u0G4ebuDpNNfijHeglv+sL+PSn/UXESL+GEzib+wcy6zra3Y6i6GWLXDotRzyu1H
6Nt5JFZ7oKuzC47kAJzSWtIeE+4d5b7LUPAwLrLxgMK+JzGelOSqlaxqDRHr6fSx
HqHjXnfEpV00njR/EhF0pVTepPn4fxVuod6ykYdqM+3jyM43jSxNe8YQMdSYMJLb
QOuGEkUGgFItLBV7Wk1f8mzKbV+Kh+8YbU+sWK7jKsMfYxHAJesmv/APMf9gRgBy
tiZ/h5qCY0IpRnpYXBzqmR7/w55XnETI2YmA10RBFqCMnIbynSCr/kpdjArfiWAy
9se5R52AHupePNkXtRUB1ZvHCWqvs4+lQ1kJI36YIOjH74Ak/Il/eDBeSnmL4+Em
7RLXBaDWTpD5og/Z5tKbVBsg77N/HSYYqWi3HZkaLdzlXkynGVAaAfRD96xQ9ctj
sp49ztvqvDQ0mPoSh7QSC0fs9xPt9SrNjhgZSBwQWHhyc0I1nyFgHWUr/YQ7l/y8
QglbAVoanOCUJQOCrO6Qo0untOXIEZWoIoXNgvGI9VMGaB2EIazRVd2lNq8Ptyf8
fMcOUisKLwOOH2s0ltL7j/Jc5DjPtOAwtp365eSTRnxt4y5ieNNt6tPHORypm9xI
83qFkSzTlu12w5fGoRTJLLrkGNchjSAAqIM3vXBsFOoFIF61wvws4VaU/0ARO0Wk
QscWj7JEIjGd6V+mlB26FchXIak8ugF7slbd4H5BOwYH7mzFDzasdNh8mVY58TLX
lXvh+Ct0qcwJukLd5zmPkj3iNZpWfvpwHE+63NrVpEgtY/HAKoTSOoDjsXZng1V7
oIy2Qkibd6zKyeROwLUdWkkbiUuTGSWKwtWIwcda61sZhc9UQXgjg6/CPmzpromh
JhUfyIF20zf8Wn1Tat6MRLxa6TRAuv5vrbd9vgH2iHbfny+le+qMR1oDUAHjN1zP
4M2NqNP5oZkzhVhCla6X1rYfrnq9yQfMo44TzUkn3HPAi2vZ9bXT9ipjXLeS6XqB
0C3kxLLwcr2K5pjCfgXXPOLUf6bJUh9wDVq2UTrSV2Udc+PvO1sl6Ts3WJQobgK4
LU0TLXKZk+FEek02+QjBGillr2VQawrCmPscKhbicbH+mDF/nge4c3nYT8ZfndSL
S5gWAvDV1sEoXLwU8RWhBz8auQBrkXEueU9TRypForozT2a23y5gjp40Y/1s6OQV
kMaJJltUO6ZdzGIdUALFw49BxtiAaeyddMkLz44tmD5WQ8ErlL6gzrbnMoYl1t4t
XxY8HeqneGYk92LmdjVhgiOTU/4oUcKg/5CPLtyhuPROQ5QGkF0X9XgsvJi+YUk6
t2qGddgnYAGmJXFKUrUO8MDvCV21HYBVhz+ybIoIuxfPpeTNB/fJda3BTAstw4oH
3IPEsli0jwxK8If1luSB2deBJxeMUXx4foE+r/RcsaU7CTo0MqzI3OZvHPvylNW+
3n3b4d0Z9RVd1aT2Xoax26D2M7LL6HypYn768oVrYLCa/C2F/l5oOWv+MCaZmibV
7gWK4uH2sy+XGLdehTHvQktjcXCMuxBt7kaZxEXVXwGgEUrkN1zm59LHwAh50gnH
l0QRkrBWH9YrzizRxV1ZyrZmmSsANWCfcf4WV1bFO6XEMKZTrdo9JO2u7LWHVAoH
e5OFs7RDVpGSAx2XtLpVRzdDo8CiTt1YkMK+tweX/YqQQ+8h/F0zi5y5IWd+3Z2W
PQt2KfdLFNIli8g7q13mMFkCenwg/IZWPbNZ3NCd8zmjlzU6JQwKQ14+8tFb9b0J
53VrwrpusKELnhR8knNMR+GlpJhR4dxMDl24IxdSF6eCS/MXgXzbIT5maEsAQKZT
DAWcNs1l8CuHWjrCOfZWS30+tq7HO/V5f5mynFwolf46eBSWI/fBZFBTSG5C0yQp
GrnRAE6PuLMhI1Xha2iKg4SqRIEwm3H7U0LDuQD5dVpuYYJAEOSvodiaJhCe7SZ7
hOxjYkcCrALMS9+IHCVCp7vzPpgwBThNLgWq41cVcC12wnNlkKFauq1UgGggQRsS
Z1HQs4JQrDdZLBEZXOOsxKPoUcgY4PbOggUr5sGt20XD7toxXMblYILMxGUZuTB7
fb8CSBO83Qk4yHx5h0NlmNcpnWNJO7qR2ti9mmZAG7nbyKtKVxbx+916gsVI1OAB
ZzRXFB6S35v2AcBJlYo5cb5AIQdix+fzTjpjsbf1k1NkKAbT9840ZDJ9Yh6wgqUa
3Qsj0lHz9XlVyXQ7Z3GWjxh59Xm1vhUqxfCr1opyoof3OTr5EanXQtQYAA9mf2fA
j5zhuHVXuZO5ZLt3UTbMRAL9I99Jrnkxju/nDMvulfL+7zJjMW3W7a3eX0aRoEj2
ifWrmO/ftX5JMcGK0f/+7eKK5itS+Tg8iQnkW6YTPgY+Uk7HS6HtdXziqrwv3dHF
wECVgPVeBsHRXJpcl5Oha9vdiwuXXZAN3PpQa1xn0wAOlywWRKHq6/FP8Jp9Xsgz
NfaFAtsvFE4jXigJS3pgVqmJ5Rp92jB+OzHnvBoP3/qv9GvT9ofdgMjFOjedcTaZ
P35tgob5AWkFXeOv3/vfBJNvFIUKU0HR6y4tsdoZpuhIsNc8TXtSQUxaGanBnyqo
bEIi+q3YPfRGjnFUImwQwNv60buMIxWgucmzaJ1gDniUehi1Vd/UATFxGf3HtmIO
oOUN9iLogzJSaMQUxeAjTsEHaeHAnH094CMJkHtsIzMnulh02QcgHrsxrle9bGhE
Q1N982fxRacViK9yucBIrd/qtb3TqaNpRAYARg9RF80zSm3D62yyqixbEE+0iYRx
CjZ3XqxNENhRd0exCGQ1Fbw7NMRNwX3gYAQzLhjWmAJJrELhDGWZoGosRCBhTuba
sNWGV/c/MdrgR1x2zkEEQniGb08WDhyyZq5xWCdoiOEAFUVfI1gLRygRQ3c0DKqq
6dIxlUIvuAFYaUtsI2S47dmZk05vUH9ufjtaBExqHN2DHroJ57sd3c7iQor2I8Zj
gAZakIMoFzlRjF9SdqP77kehRyJ1Fy1xcscVqD6LiOgNCQU17OoR02nHeBpU2MVg
9cEzt30dc3O+i8LvpcWWSpC+qGm88cgXfLBntBTvbIDXQ0cwDUN2aRkihwdhUo0B
trqEtQWNguG5OaIUBS1at7lG5Q9Je4DxEQ0t8Ln290WqpuvWNeOczhqqxYoSyhX+
nmkMOKyztWLL0qpZXtuhzCjYgWue3gg/RfhXhinsgFuhepQ9TzGnSGVRv91Mi+yI
hg/TPwTCiNtSLKjLBPiUrlpmdcPqmpuWzvDVve06NSBRSQZ8qZLfSFb4qVDl8Vzl
R0jXOUjXOZL6ddfsJDgfrM14bx6LW5tJ6M2/62JHOT2BOWIvbeJ+0Iyep0wa1KpZ
/Y2nGY4KBTPrnlEs9NDJqRo/lV7TWRuxIgK2VtAhBjOxdqhmfoTbSSBNVVlgjQkW
09shn5m7vD7Qf6qWEAnwGicPgPzdo50jvwxduKqmTH9dhjQ4zgMYQycauoswk21U
pNU+3en0jbIn+1j3k8jKVKcf32FUWhxDeO3/ngm4NTMnW1OJZxkE1oGTD6x5bRq+
BZRoUjoo/L9YjeKjEg+1Qt8ZN1Z1GAW7PcKCJevQnrmtuIdctIeiMb/aPXcEpmcE
rAze6RKOk35vTspi5Nu7/iJN7tXzXRPQXaJ2BQ6iFJO55QwrBOW+4x8oIFcupC9a
duz4R7TsBrqwOEfsZOTx95+ZfM4b56m3l0P5vQ9lFtD8RyKesty1oWpxsg3fwDUr
ZsazJ9lmYdc7o44+z/kDmVtw2O2VsX23AVFpGe0gm9ZoOm5gwM1YvTxzppdvDQsK
FnoFu/pwwqVZLoU7kb8JVn6eHnlhDd3+pbfij4mmU9W4auVXJTQQ3dv+7ZArAyHT
ta6PgJyxEDuXxqRonl+ghEZp642fKRoEWq6GQyYriXQMH1/MznXPrNgIsb/wP+8E
wv9z8Kfw5qmdQ447X2VYsfFjz3DW16Itm+VwJLXccBSH3E2GIqIpivnz+7qV/okC
xpv0AQYUfQvM6n/Syp4O9Sc0Ro+Qp2KsjrWwqRbOQ5bnFTWIZx+pglckcxqIkSXm
y8wIl3z86GmYZDV5wOIYYiek7JfWaqSM8LJXVT03J9WgjENS3yzBATEWQg3V6XrB
mFNA2eBloeF8sHpFeQvrDQHY91ayOuPyDlkZFGpsJGvmFiEqDrcKbdZc1ccRW+Ag
ZGgWoTXSHse/fpkhZPIoYcaJkXGC2k6mcGcI/+AIPc+f6+J3gJMrYdAzHsg3CmlV
rwHy87kMWF8R2rina+dNoznv/XBLYYiDFTsVw1+79w7oWecey26btmj4o/q8EbJi
9Q2uVhLKtRCCqxePAvmNNxYo+Ef5WEU9ANpMbib5SFaqCg0tvqPl58yhSTbqj/qD
ZuRlgNGEYEmAaXHxWM7UH5WwcWXETpagNZT65v/57Lnh1DHnF82AUbkMqM5Q4USv
Z5e6I8IiSXjt3K9yO+3D5L+5D0YVXMI++jEQ26h/kGbxzwmq7NMN4Tz0tgBzbl46
OoeEtPUpDOKO4kxuIgDCnGVBpw02tDajLy0JHm0UW29RiJNDVPBYYdYKq7v+M20N
PNTj2XuDSnPT+hkIe/CTTzeHkvV+j3b3IIVlmzx7I50K+U8f6LF/kh7uzrkiwGXe
B1IUSimWNq15f3G3swPcvFDtklIWoKO70mkewlawaI2xeE4j21UfQ06D/WLbC5Dr
pNebKGRRfAySv8CzJUyN7vQaM9Eup2zn2MkWCdwuevovHiLbTenpToOWlvVNkrLa
cROjkYReP6dF5WXXJLLyclMpl1HUr/bt4VbCdD9J9EQ4bYg3mVBsFl+I5QqIdvlo
7u4gRo6LP1EDvUV8pLA/UKFqTisGPpnvw+PhURQo8FJMM4oVoGa3i86gRzZBGrzZ
X5lL81h0dI38pjWBcvFZhSIGUlOq6ylTsvrrsyW/ExefCNpdwGPubP3TO0ed5B6s
lOzc1py5dg37dUrtBMT9c0fa9tS4aDk11cIPQMQGj9bbhUqF70rC2KlfES3dRqkc
WTDuCz74KhN/xjMNpjUrz9Sv3r4s2PF+Goyg7EbA0WDZ4zelcHVfb3h3+fs/7sFl
PJvWaPJ8trifViHvyQFzdcigHFJE8hNRX/NKzqjeup/jLhAWIZCqm9Ty+nR70W40
mQMutAieMyY5FPQnwW0EgFPz2vGUthhrwS1jnEQqmJRJIX/QS74YzYBp7Ij3hMBa
uQVIZ50K+/vjY/gHz5yRGic2HJd5ofGaie12e7y1/XYFsoxXX4JKXv0Bwm4m8do9
1K+m1GDU9EQrZwRAeaHKFNWzwcAhbdW3SW6qLBLPZ3NVCrH2utTdRAyI1BLMzWUS
MHyGaXrx6vPlJ1Xv6oEmar20aN9CNZTBDN0gYZ6r9XdTovZFiR8MqPD4fMSZ2CkB
kkK8MMLOh8On9F5PZoEXhOkMqEPPbIdgA3GmliNtmSsVnaYf5oDMk75USaNFhVq4
6DGmhrVVvZLnRwU9bTBl/oehYF5HGYFnQ5Ev7z6FyWFV634XlLqkCE0U9jhL2OYk
t9PW/xm+0Ctu4+oLwHSMUICNSPDOQNC0/4IE6g4fbNLR2cMJvIon1mudYI0tlX5E
3NzlZDQYLTyV+nDf1Tc73bll+7oesrr7YlSAiq+im3cq+H9jPugRdRpE35zQzMaJ
SlG5TUJjWyif8aedlqVLWxmmpNztwQLUO0Uu/e4S8JXWhfTzeTVVsmY8cq1935Zu
ObfEhkDzbmCe2p+rO0GKhrFoAn6fIS/FOZpxW0XDBJR68fq1SHxYx7CKa8HSZH35
9ezL7ES0FmGxOfn9pKAMzp5YjvXqkzswXzb0uVMNNsKYmD7VkjHtsNmhJpdkW4TE
Ema2W4dtJKz6K28U3A7AcpVZ2WnI207qPf9KRTFH6D39ZoRPQlqjgZN2XfHz9EWW
27DlQi2WngL8aFlbJRE8v4X5YVWt6NceAXROoLwUZv6ohlI1vu4UHamhh0iiIyCI
CeXpINIyWzSCUgtcWpqE95gbTQmgvRb81Aj8nmVzbtuK65jSP1GbMMea9bU2eXGA
gmBlo6F6hFeAhz680UPEj3NKKUMHvmnyG4OyLxgT7OFUxXuDHkJr/4al5w7uf7rZ
OAwNMUOJhMgF3WJ707Y5sV2S65e/y2Vp9/qCH2enJvdlVm2ZdkUF+AcPdliqJsBj
OA5j8Hz698RsGlD143iwg2Zv58tItrgv8H44JY9p63tjhtCU+hzNVCbSvSUvcu3v
pAJzFl4cL2Yw0infUjPol2qFDhslTm7UXjLLwj6F07h/7MGBkGYAR4U48lzypHUR
avRIo6/VeNle1Q4qLVwwc9oluEvbB8hkOqLLhc5CjjrnfU9fftDyfOg+1vOoa6as
v7hK1DZMR3YUig7MeE/dSsF89613b9Hu7A1dYguWeNHbEIwQKNmhQQtpe/vZNV+C
1jUJk4o4cb6HM9fmWo7UNW7TgUeoVeNsHAmNiLXsnvi04ygF0ZvJ+ZsxaRZdE5Dr
34ntARi6Q1kQ9nLJi2dYs8stiYO+pSk3sEPpBFqkQr+XqYHvk2lWQ1nQJFPQ98gI
i3pBrkl4d/D0Ifp0bw/YnvTNmr2WYJb16mK4Gf6JXoLVKQnOn9j+6SQtxZMN5SLg
BIjFcSmhj0+gb70x+qZ1XW6v+kQgJHvjZ2Kga/9AlSprsfhlD8QjXWbm7p6yeWeS
3zoZ2NkC4JIUqbVLNQrnHRM5aLxcaJrpjAnMmDLPbYG208fMEUtuHjxrRzKMpuRr
lTH9yqm5DsbiCm4Rm7NcYyDIWHE6rAp2AEF7IWREngVodPkLCpZGBVC7dTznySBF
ZALmrhem95Z+Z+KozHMRirJNJyTi1hZqJtYTpTh12NO2TYaXClajj+HnKcQUqcS5
Aw4AlN6AuUkHrJsMPbayrYUeq60Tgkh8f71EwiHi+KYb2ZI7Df1/BgFcK4Rw/l1K
asOTBjsNgyG/k1mkKKYdGZkQbHrWPZ/nFMYZKenQvtm7AqAdNd5eyxio5Jd6or6Z
EFPQwfnKVaFdmv5oxSor4REn5yu3zDoV89eSzVSS9zyJcMUQnlUaeDnDyYvHnlGX
gDvWJ3wWDrNfeZF9nqkOhiQO376syIdopCQyfBkR3bAY5NnBykoYzGIu1+fTxopp
i0C5UYFw9GHPLiE5wc6ELISkXAezgeOjl7JiXFPOCbr1ezxZf33wv8KUcw1dAZ1s
m4ho2XjxE/1XTpyc2UKw5s7Trru8dxBHti2sFJ7KGRWGWtRzxqn7GQ/G8xEGGxJl
QM7XTljiLxyYg8YRbicWitIS1KvUjf9YdW3575HHr0xy/bGFlF8v1SEfZ4z88EQa
HulYzsMWVbmbfCrvxPck4dubDxd3B5Rvk0OipoN2YzM3nv3f25QwuEOjyzfdyXwr
D5o5i7l8bL9SJJJsTPjTXX4Ucnl911vrZYRWJWDXeoqVfdy3zAsgU82ALmVh4PPX
CJyJWwGGBSQhlBtPH/qzDeEDcXu2iaDefaYneul48jIvBJaDiIccbR4oG17buJNb
mA3hcDvb3184Wbq3m6Am2ZCgyufpDtGjhXsF5EH/Kx6AYJvc4LkEVGcm7d0tb9jc
4PczqE6YqstldMFaX5hHzMeWf+me3dBVttrHe2XCZVE1nLtP7A+PbpIvCkUfbLk3
4wsuaCZEkIIhSWjbitlzj6/4aP3Lq5o7dvB+0GMZVkFUxhgKdNBY/e15u3pFp4RJ
4PzTFkXuEMVcXMsrYHA67KnS0j5jvH046eckhkcJDd52ufW8BwCvYMssjldSMrUC
43kJPZdidg6aDSOF50bdkOrX9/rYo9u51T65ClpjPR1GPJnqQlk2EqUmXNlo0Fc6
7q0jCeKcqRI/dJc/nX8TonSJI5hrS9cz/C0Ubn2JxDe7Xhm6c3i4uxxrK5yHW6l8
C7Cqm98rAqwazbwBN0+YF50hYorW6XSTflNKcUTwxwcy0iwZkTvAwul73HMoAqGy
koDYbhWHcr5vw1uULhddb1tApSLD6MDZnC/5c/T9SK1cjp84cURYtNEes9BHI84T
Uo9mYwLTgNzdTLQbt88z2FiyG9TKzYap6uhiMbyBOPPJxLD5eOEhtNoMp5uc7LV8
SzMFk1cj14bxhYu0hbN6fchCQnvtKRh0cyJH9n81LEh/cVEC/0TdgOmqktxwx7T4
Rn8vyTH5AZfo6SFIPTRMg96XE2+HH/+qVtfNMFek22RRATmJ2etCVCjZCkR55z3b
vxFI2D2tb8dWrPnvCGpT6BBoxdnb4RMCbNZ7xEI1rpq4tRLR4onHiVZOvcr2qrd6
3Mjps88DOP6cC3nJN3PmjSw4hF32q6Gz6Mz/4WFdexw8BjMxXG1Q7KtwymkalDzT
GQvY1sJBoRqXXUow0W3ZqygNUC0wuWXTKrObmU6vaKsuqvgSv+Hbo0jja5d/siL0
kpI41kA1iZkmIf9rLC1F82S880Ej5oQiXQPkHT8z+UxtcHZkHcWa8j9Vn/7jYmI/
pxNGz1ENHSXkptNNVPWD7rwrHf9ZTx8N+VLyy3wR240kRNYbgvpfYpAZ93cbKfUt
8qHf7Ra/XbJ/HI/n8KF9HWMsQnbdW+bRb3T57oGhVmOfJFCErVBFi9aXzVQbRc01
hYiwbprOomoxxNBg3zdj4dRen2/kFT5xv1t/0ec5igd7jZCqwVWjLyppiTnQGC2O
RSL0g7KjFV0xXIKDj/ZVZvuKzNkHOsZ+GbaUROH3mp+62+z/8mFE+naN4LnjnRR9
mBGS6p52G196i7Om9/cUFGV399GklsOTPGPvYSQQ8deTRs09AjH7Cdc3QSxPNswq
g6H0uQbH2Yry39bARB9lD6iJMoTlyYHNzXdncBTgYPGK00UXBHk8Zw2tfkcXb/Ov
vLIgLhc4uQG6JIy9kg+Ahpsa2dMBEyjON9L0zqlGw5ynyETEdkmn+KwE7rfKih6n
i/0h1o9OXBqlR281AW+3U20jbbzexcdq+I4S9dkFN9eUkyAYjcDSZDluuaJq+R3H
oJf+csWNRC6V4Lc8rmPJ2FZ1OhHRA8abP5NGVWT2ib1CruB1R5SA37Ded/x+tQgo
CIploDT6gkhgB2OjmkOLf63ukHjISGvZ27KCYtECOKv86PFaq43kSu/31v+kP8GR
ktzbWH0Zy6hKAaWbHdTEG6RvCdtZlebPD8Sn9V3UojJMcWDCnGQLRN9vckYOizSf
ibKZx6i8pgyKFShf3FboLwM6CmZOEsctYs0ldPg+1a9GhR9uVjJr9dymZs04rusN
L0tHkP2Uy5RuduInXlzpiLZAlmiso/jGpZ2d2ZaKEN81okLckfNerbDPokgV5cxk
6PFVdyCAUbvdSiX6hGUIqY2NCqD3bwZN1WmGZANPD4LRKh6IUrbPQus4g8ElgK/E
+nMDiAhdM1KOjr63PUHluGNsIpc0wJnm/XmOudqAcgz+pcbHvHnnCAj/JZWLFfxL
Xt1vy6VXnZfe1VVVFHnGiKIrbAXOAZNyLBPzUZqDc71TteRxymYIpcS2rVirvUUY
OVIbA2yiZzNeOv7yDtb0TuVwsI8bD5qLRf9mcho5IB52tOCBX75Fm3Hnq2glSEz2
oQa0pgEPoj/5+7u/wY7BUeeASQpSXm9ClrMKxYHOVFd295gZLY5pPI6dx5AH7YdM
DUQ9RcZTEOOZzP6ZnCAabATKNK3IpbUuZVM3oDjT+dmhgOjLmB8bGHclVQaOnVDJ
YlfdWnE6pGU+xfxyd4ddaGKnkLSq7JsGmBifZx8/UkS/0924V4+5NkUnrUnpoRQs
nESolrbA7co4rKH+lSfkI0cutpOMGYcLO5C/cBU2kRuB3663+Rt+DPhW+gwjMNeH
GksM3GaRbofwL7/ZeuFOW//jsEUxDP/SeL/EvMpu2cM+3p+f0WI0kd0VbLdUJD2a
dCTh83KXGfHQeanuwoKE/okjme4NFKovdqVXhsjrK2LBsagDHk58I3T0GkQ6fpS/
JMakUyIvHs43wDEQ51bga00lK0541JU1YKZR1HOdIuaCvIgXwPBdsacmxJJQfkkJ
u3V0QN9MV+D994Nbc2AvXP/Oh8pmp4u1dBcvUI58Z1h164C/EJZ0MpEHlZ97EOmJ
vYFnuWV5aFfQwPP7PCFjgTIdZJ1U2dFgBg/JVyQHaKJmWxwJGDH0AMyjSJD3r0vh
JlAfO6pF4G7dCr5bNUK99EMtr7Onoi7zWNZpCw7qiJep41qyVPhPspTPYuo/VnmI
9/Te7ry5GSZbqTbCS3klqdzccLzjP7uKDwdDAh/Qsar+HWhDV3aXmzh83NDmt9Ai
vv+5dryCLzMrxrkzwlfmRXWf5yQuDzx0Ntt2XehG7ryN21487Cn7iAm1kEA7GK/m
CEnOeUmPNj4ybXRRR11PSdO4qq+13x3SIQfSJnoaA3gQk9QxeBEUZy8V02QxApqv
2kU21HhKeZGZ2H3OUXQbuX0DxghGObxx6LUw73zmqof1Kesi8foyLoqw8MvDTVlh
PUJToERe6l0u5X3rlFch80jMSfye53q4w7IgGSeIyg+7L2e+AyYkwm0W6XriNgjA
TpnfmDST6eJryClYGLYS4mSSTklEtiUSkoKDYBsxaiv0KIhiKdDy4r71KOFXN7k0
22pmYOuF+Q2A28RttqN5lGZhD9xb/hgl8c70zC1pBw1frLbWaFXbYE750Scqudzh
wWJ2XyL3I8aNnsiceE+6qZJKt0IDoIoVjTt97xZ9L4VMruW492ao2fDfmkSpaSIc
vLF0gKotoASYQJXQDXHJ34gWDNIa1afwLm1fMmDxDBNJ6bO70bszwt1g5c0dMgu1
2NAUeWlYmbbjZ4bFlHBcW4mbe27kwioRF1pzWgE9vJyVd6YIvRwK+RRO5ehrGD+w
XHTxhSG9zqvmplI7ExxE79h56v1NX8kIT2vOiIF8LYRF7fExGeGcj0A+a5TWPkch
dyYIOqVpvw4GS8Dxr7b09iYO1812w7u24YuynKiPx6idJgzFSCn36a96lyxf5CXh
2l6xYzl6JKCOrl3ASfE9/MTjSObMTwt8uW1s6FIFMYN6X0XF33T7+AndguvJCqMi
oS6uLhTYdfxzcZxgHEL9tLKELG57mX8lYuRxQJFzv9B/4txbncO3o+x5Ytu53Voc
uJ6LGBbRlIF5SIVWW6dzD4zR1dsZYOIbKAtqfDO3KImXzvIKX1spGxE2C6OSeF3a
2XZU/qwtJlPDZ2kiRLdz/MJi+cdTb51o4EdKt0uKX7AwBAlu1QbHYLe+d5Mu8gD/
bwnZpTzGKy/ygXVurb1qSAxDx4k5yjwAnMA3cyUa/MJb7N5VLfWxjD0sDLBaIZr4
Fo0U8X0GBQRST6q+Z5fyZBUsBcbDsyF8XY7bamaC1e8QV4IgVJWQX2ZiAbVPnFAD
ud3eaCUn49puRSXFL7pSRXAw5Zy91Cjo69nZhLyP9/Os2Rir/yRAcvZvsDZhUthQ
sVSjZUNowVmXECeokyJCcR12R91xOEtEOMPJMJkxW8Y+R+KEaDCr0EKIAEL9Lv8U
ss/txVwZv73zGtL/aI9zjEewAR/L+GR6Pah44L/Q0aMzOrOEQ8F3M7sug4W8hdlD
hde3L4vsOJkQMNyItcrCPKpK7Ck95a46OatRjxbUxBuPUiKeyvRhgVqTssT9WWNZ
BaAkjpcoRMc/XhM4ZMt+1NkT1aUi0pIMN5N1WbJR9o7+s6bpYrzwZoY5O8TVz8EB
5Lv1ojPyPIsx5ArRH+HHKTthrT04WX86VNU/Tm723dgFkuFOYv0UMNxegPemWYM8
UbqdYb7xfwpdTACZRJnsFZph69pFvGIVAvfJJuOqojBCTKR85wwVqkwVQ7xaslLl
uiYDR+lDuLY1sHDgfLpTn1SqCewvdPiotY2tuzfFSzz2XXf1XspPOw/UK9ugFRMj
RhDmkheMkhfE9vAlS/WoQayLmXKpARnq/Wp4GaZ2lzSIT26wI++lT9jeQcRyl3zk
JF3ZH/A03F0j28V9+Ct2fP7DVCzPoSo99Ccr44AKSxu777KEGnQkT0Mi1zvF5mYM
PqsbyXfD51tKQiNFGkk3tuTHoOphgUA5jZMmSdKhygVM7voIoApTqCGJomdDZS5u
RoiDnQc0juIDK2nun98EbW1/atHHzU8oPTowiteG2SZu1PLG9cNPvnn0RNtNcw8X
fAT2UHNRHU+34hkg7UWhGn5DUzs/VL4dN/hhhbyhSiOiPzwU72oDnjkr86WmWabX
PgXAGEWATzvxzTyh8OF+btgQDIbTSU7ZC9RXW8QdvSOvSm8OJd/nOyXne7eYyXcw
73vBB6wBV5pLXLnte0VIOeTRBDpmQqfolP9Jhnpo10aEfBA2htLk7a8JUa6Bkvfa
IgYCJwHE6bq9g0QClXJfzWbWNYCEocxSDWzBDVqt/BnM7GCfpmXFFoCR0eqGBazM
PzkTZFMVeTz0/OzPPHEToU9KXtO8t6Fbr/VNEVI0MUPGAfmVD5t7+5qmPxFaNeCZ
BusIcKrfpNhmHFgjHfDVEzI9l14ojTb4GBBGB+TlrLZZ4+2+dN/QzSrO8sv6n0AH
XblK0kmkrqR4pr2tFJM9U/DBX6Zdj94acH03VSvxrUOlXYYKQPsJW+WSL5m3kGCZ
8twCPlpLJQd/tvFdb+j4jrtjSNtZnZ0Z3knvHeSaill1hbh8Ce1htDJtKodT2ipV
BVMABdFZxlaountHMR3MYs9xMZ9QOcHzxb1mvRqHvqYPElc4HwUuTcDvnZcd6ddb
3EuW5K7y8s7ogLVfGYEqCraOm23sE2CLaJdICZ0kQiFyocOHBcgLwOsND3xjFg8M
xJE6YiWjfdL1wysBttWMvDsFqWcGylVpMX0vB+v2C10cRLOKiLCJbH0n2AXUN/PF
bst8LGofHnChMtO0vYuHtVGUtTxMaDpUoNt6qZLovC3iogu2kSJmtfXihaReqcxz
bQml0IaCNbARa6+KH+QQva7QdEDfoKQh31rZQyE9iWkuf0yc8i0kyERc7DoZitU/
CYCfxWhVVHYEkJBtUXSF6MoWmErWXNH8X60N5s2NPZODsBnAv2CQiKDasIkTn0VZ
rv//yN8pv8c4H5O4NP0e+EgW/y7zIFTBmJrx1Ys7kzYCtuEtrU9sPEDxiBtTIGlU
iSUD3haQ0/d+COhm4tTduabePsfaAQx8zajnnWTLQC9hWTFYCiqiWJVb/C8pPUXq
4zRfPYvuhjFdwMvtqW6FxrvHe/uVQbdA2FYVQ2RhYAc1TELE2Ty7d7K6ex9EPGVD
9mc/jUJV1J4Mb1hOX/dwRKlT4SC9mu/XiNbQGLnV97hir1rAb74CndzJPM62RbmY
UMYU7fr2D4Mz0zldFuuV9aHXE16+mtVdPdC9bEO145ZQkAleG2f1UgaZn7Yfi9xb
/jDQmoFDIa/q5t/zRpvOSxFvn5tEte8b1LUnqw6+p2SvK+WGvzFttCthFD1BM6xt
PuYJ1fDVKshSTBRwb3fuLCPtTIwXopJLTQWsCTGhYRnbsLsvrEYCu1qV7kzrVzco
EeVsFrKt66LmD8mQdLOmVyUK8QH8SF4btPjnxhBgqMeueD6DUW+6Q4RTanqawOKT
JqcWkoJ77+E7ntB2ztrIBylMRi2t0hxxvBYobM8tHQkLkgDEwgVClsLcGdfTybES
q5RCGWsSL+fDVBvNIWOD4rlY6NN1659FyYF9/5njmXNfII7Kh2YgobTQFSCwkz8D
mGhgM7ZTJEcFboHeluR/NFuQ2QaopL1zE354+jsqZ+7nq6zKrT1HVJD7D1yNfiNE
W3Q/C64F3ezA/jCNdh1SLumzbMxx7pVNZ0NiCGsgOglN4ZD4IR99dgX6JS4HWM8J
D/kMQL7mEkPv3QioY/QthI5Bg8NQQKPaTuKUtT+N68lOTNtueRxXu+DJG1ZPQ3qQ
ss8OAReMPLDAtvdFq5ed5a5mzF82sqWiw3ULz2cwn3tPxCTmYfG0EaipXMjA4wL1
C2FvRbf7zaLFXck/w9x2Tyur2S9zCWGuh4DkG7wfhzI06xo/fkNDfVfEcBnEEosy
Xpyo4JYDVmklUIUjwP5wkWc8I957KXJnaNxMWGNdmJCnhpUhNiR5VFRluo1eE0m4
EtOEoqivBFgSsbvzGTSAk+Hc7d5HCLrBXknA8teV4VIutLYIZgvqJhxYVugFPJTY
K/jpx87t2Kcw2mFjD+glTmkA8Sm00Xr/phymFVQC4xaQ3zc24KjNxKJnXnraknZl
TsKmAGriv4HeLwGOsWFavKk1HsAHoBKfWmd2ODlhFmisZRtCfgmtNi7ZfIKexAoD
01UtRfkmFbmgBAY0ZkpYMX4qEOrQsBRREOxNaysqo2u3IvKYVi+eSLULW4QPYTMd
Nc2PccjfV8wZa+bMFFpsZl1TQodphfDW/fLBbApoyd9P61ZGP9VLGSwtTohW4MeO
HsCXXZAlsjK9bHNObsyVipaLjb+9eIZjOsn2AQBiVGwUPLg7l+jB2DfWI+RD5D/M
fCSafmXrW9vW8h+1opSdSh/eklFtcEDLhGurhTvBogw/+493ArdUnWndMku0r6tm
4pJXLvgd9iI5OTicCzfYlASgyS3gDxQnvzSvlnrKvIjGioZpoXRvKVCVsuNSuqA2
ld4MJWbXhLPNntecSmFBbY5LLs8svsTjD3NRgpzl55qdGk2N2MTbNquu6H8mdqrs
PqOsX1F6QkBm9NN65eGKHj9bzNYJ9VTF82AYE2zuwmm5oT30cy8nVv8lcQ8ZGeoP
5Ab3ZdgRI+FlUmniHY/cpZSW/G4kBSEaV+vXRkxAuoq9Qz/cltixvHRJ3SFse1cL
eKrhxOYLa9h61/2zlun5cNrNeDUosvBvK7Cl32lcxka9IJQjZhVZcH54di9f9RJh
4ZHPG2gp1KniLO9LczKrmRs0/cRm7+ia3BZ/KpfY7VQfuWpkbAeQmqdCmJ/c0v5/
MJLsvXFZsX6qf0VLDwnAWqQWXnkbR9N7E5pTNhGrLBg8oRVr6SrmjjFiJWml/us+
zmVLi/C+osPlXKwKQV/zgo0q09tjaUUXM5vAzw8OTKTYrpG5+uXC6THrfqiZZMyC
GrWkUNhDBaZT6IaKeckiUZXT0wFOQCxQcCbNU9066J32qETfVK2rJOU0BquI8g7q
Y45dR2e08n7MzfKOzT+ovsud7XExW87+jl/LBs7TVjVb+YY42llxyfh3EBm7ao8f
Q8QWhiV9zXooNlNXjYCAJDxTveyB0m1y6hIVoaiNQ9f9Oow1ceJCk1g6BAnulVAR
gnYeP5G2G7GzZ1i6HbyZOpOmM5sJJVycDcko+DmgSPMm/W/qMTrkat3alUNWWO/K
sVeaUAII2Pl1xedPy0mkIRLrJIQ/zJjDf8RMan1pVnq0D58gySbgCQ3o14Xi1EUY
OuzyJ/UjcdpogCljEeN9A03xyMzWCZx2xmxM3BXouaK3ifd0neiKqkNmSsX+NvYJ
C1RWxuZj5Ke3QFyUth2lilHaj/+mBkdjn0QrwuGmN0WwpXWvhb4iZ+gNF3ls8CHu
VXCD8B8Ru84bAasH6vLOJR4e2QrGZV0UXD7rTZ5nkOPNJrhfMvXpogCQ0Xoft88t
8RBF5fcLiZxuXMXZ40l3oKVRMqYUXDgfy+iBU5M+J62iE+xKxRyKpn0c+/okLjhY
aH7meIwZEJ1jL/hqw5UjX3i/SVgUCbpHfIJOxdXgo6nHAjKZtP2yeacBTv89tjik
fp6hDqWMrIYIOPXWaPEG/3r9AguO9TrCuKeeTexPOvemJmQMBHMVsQliNsZ08n4y
cIkrjIywOzVDHnzrxWvlPDsgMXE+VddbmkprQKBtQ6xLxxlRrfEah9NWonfLLjqo
Jo95MXK4OExQdkKfO+aNfuAKPW8Nv0LfXxMy8mFiC9tEocsqvaefi3fZitAh1TVx
mxxbaHcBYxObAX7kIiexvMmxFI5QosArnxQU32kF+DuXQhzirHHr5nM0MDLPefKT
F9uajvtv2Md+ufXOpy2lojwEHaDAROvr9T0rEZuOMCYmGK1ic0Xd6z311uD4sM35
6jYotZzCLMhTZRPmnCuohYctI7JWtDQheSMmfhlfqJ7j4sOXh/rlvlkos4GuOdNc
HV8exeZ+rspg7Cq4CS+/8FfakkRlB60dFMk/reEHSRNMCKs7hfwHz3dkW+kcFFdK
P47bHj2Ehg7DEzT7ynmg+iWtIRzmsrzjFJGZHv+XXbW7L5o42f6TSG5sembHaO0y
WWi9ux+Cv0cOj+wiyLGC/y3gqS9SrpofMBN87WazDCa+9ve879ICNU/CAvqKbGhp
39bsA4bo6pzI6g3SMD7Ysz4LirhYc+js7uMkeFCQAUnsGdUD/EPi4PXO9s4ZncxX
aFNzgQW8z4gMQtSd8TxPxKbcFml7pYq7HwIWtXtMj0YXCeReamgqcPpdd4wuFQ3b
HqiatmhExuK/cwu4W+kvI0e3/5rBRyF5+2maZSFYtJLG456gbYaZHQFD6Sz5U2ql
xnKmdg+yX/PSyi9NGtp+/acra8jHEVJGl8KR3YSWAAzqdW5DU0BT8xAMBIWzuJV5
ZbMOw3AUR4m4CVGX0pLMkPEhXIQmi4iilNFP8fmWQRiFFdqOQm2lRgl1O0v3/KwE
KcXIfsyPX8GCZyxb5adv3Nuu652EzYHqtzbo+Sz/clKcIvv+3qkJQVwrGu+6Gnov
0RkNynDNDtE181UTLThIeKOBcYYb7zKe/rZ5C1A769/jgWiga7vvpycozeGdOy2p
s97D7lzVllLEu5pJRZSTruQ/8N+yqGl54olSVc1ZlQARNWwGa+Ooz8aNuhUEGz9P
uWq09AIvCLz5P8vhjbvq0HDteo4m5SPP/YeKhTC5evalKAxbCtACsaA8lwk+qXZK
aCWA49ryShmUtHzFiLgGBFKV35dF/U7fbhM3lqM+SoxQs+wE5hG3AWZ5mOAHc9c8
zRrIkQU0X8pIXGTm1OWnTPUQjEDmxEOku8QNkUvRBqLBc7LwjeP7Cict5m/h+6pM
aB7+IdJFH1qcS0hWOPkOLMDr1YsUq9XALPwwnp5uB5uvOJhEnCyCAfJONcwzJcXk
51dfiHSQb60zPtj7nixc3uDCHsptfu5nc3wF/FplFMe73San8P5te6At8hUui2UR
VsxQ1pmZeVzzopvdYbRcgzFC3vaUsxSu/1oZ55gEmfVr4aGLUjzzXr/YiFBSNyCf
X60X0cMKbqT47tthlRKnenqLsQbjIVwUdqjK0iOZa6EHw2UkmPUuZj4i0NeZNcZ2
TtZLx6oTHvWSvchpzg0xyuvLjJKlbP4yG3LL37/XyVo+rPl0PQRNVwRsOyxlqIfy
JRFQZFOr0sGsF9218CUOFwmqZM8FztifOw46T9A/Upzw30Fz0VM9fo585jphvXR4
9quGXpJP1VBQ2f4WG1a+4j43E7qn1TTGbfxXRz44YlCpKJIMCQ+XpMgogT25Y5aL
/XRrmgG7jNzHBs2+PN7YiH2ntBfHDsNPnEKli/R/PK8hdQho6y4qWjzHKNjz3/td
2oTnWR5yFrsT/n+vNrFWuDbJeL8oH6EUCWGgbBUS/U+ndj7kfZyC4Ey0o8Fr67NQ
gesLvmEEgG7nfTiDO31sZgWaO2PU9aXdPIJUxfqAiOYyE7l5DW/AyebX9mxj7YM6
NtsArL16wkHM3yIN6kE0sYPGhwsSbPwjzg0447ajYhhgZ2NFiRxLoloFITLQHLJe
M91xKudyp5jBTDN3pIFzVUg67SEeMIVm56GPJdRJ8wna3feqS56kDKgvPgm3RzhV
TmbJGm37TjlnFiVAvP2RqkdSuDLglMEQxbm8gbELQSAD4UZl1yRFUnd2MizZp7R4
eDjCetssBiG8uTc7JFp/oCX8/GHTw6kMi/2eAOmyhX0kCgqlc56MF4QPOuMHw4pO
mnYj86PJE6F/14YyV+PD8AP6SDBuTcU3SOtkcKJIgI2k3/4b8fqHJ1X7rXzjwlKD
a51+etlxA/PGYhnlVevf0rAu0RcgA3wNZmpPmG2YFoEIEK0D8ROkBgGXE3oP6Qf6
0TGZDuWBQCHtvrTKlPkdu9QmHY+dCcvfm8YmRkVCPq4fw5g1QcLugzkeGMF5zFBn
4pVWbdA4GzuBjj54bT5mtJel7GGsd4uLjIp5Q6rsvBTRa8DljQO3wRLiqW8kI5pp
sjSHhsEQp5y9LJNHed73gdZNqUoasUF8O1RaJcdKA3CZFIjdqLmWuKiBJ6nuGV4c
MkRr381Doq8NfYU9U0UCXD1XI04Eahj6ObYdPzp2aTpLbyLOJWb705fCy8QbQM9h
agola91uP9tFDvmE4V9SDTb1NKVFsy5gjp/4+J3PD/uZAWsrysrjdoX26To8gc6M
HFCpzSJfDGCxWO2/unCJTqpa4nMBXve1UtWoMvac+WjwyoXFNMUyKogEdrVO0uGo
Ik9+eiNVBmxE/vI2HbK9JMUZGHozcPkbYgqll5RCFYRyKf+49B9JyvLac1FUqmpn
/usEJHPNFAldf9Z/1PfMzJKpOz4GU3yDrAfbJ6acXATS2GX/IA8ZMKyVt32rqB1M
cdtQ3dCQdLPXePdSKzgR/dhvGlcHxZPPNvBqJ25JDc70S8vUw75YDDuRtrVfZTEE
5xdvDz/NH/tZBUbDSEGrIxiCGhY1mK0rsjLrvNgPu6oiQetPVzMJtdgte6i9hhSR
S+hfYRNBzcO1J011CmL1NolRnKsc4f3ajH/zJbcBFqW+SHsw/tnmdEvtvz+5Gbvm
tBR29uU5aEeQsTumCzkMq2BZ5jeFRjkKRTcvmWAQLexOCu7yhtPuX5DuVHldItMg
xkNG3TRbl+GP+mEEqeTQOlFvPfND0CY2GwooJBNp5w2Gg3+2kr/V3VHOANm+Kn3V
I91FEbI8mvWTrD9GI/ne/PkfT28efquBDE9fXu2gSn7+8DX3+VSHUhYBGC5mxmJN
sKd237hVdUdibObdtxhuH+waOAs2ZpWURRF+ftABY1jcgbPCe0DgfI24AdFKUYYD
Aeg54K0Co/dzhtJympIhvLJnGZF5b969/HR4Eg1NP/WuX4trXPJg9poqXXaKUbFP
DkgssiQv6KnQzON/N0i8JYw1+BGVrr6agJyK9LS6YmGz8KSSiBSxjE2OXw27Jj+6
6Q3MR0wN+8KR+d1XZWPlE1hPAGBZ0QTtmiJlz0eQD8GfgKLhIulkBrZHNCxMa8ka
L4xAQBJd4/WoXHH5xUsemb32mxiksrO0FMH89BDUlUb/1qxU91CMMN3iqDha6ky5
IcYtaQ1VQ4xGX/xtE03YfZuEiyqM+Zy7cpSaimqeA+vtAMjk6a76PMXX7KGXEO+Z
aylMFjvv2o05hcucbiPmgY5vprC9HpVLLcFHYOkr8I5xUFCNb2+P7sBVWJcetfhK
Wo651hfh3KzIqC3ADNFwRMPzLqknQ1oY/AN5ETEw7PGt/ysDuR7glt7ke2nBBb2v
SPLxnOVUB8O1dXrutbEXTmKIytrkQVK41yCqyS1kKmRlGj5C2nT7olbsaA8xq7w1
GntwgYqq00UH4LcbZ51M/m+d6gooVpLq4mOlDwWHBhvZ754N70YwNJT5+LvrXxd+
GmyAXi7TNBjMvdHb8IDYkTwS6pM+BGKLMmoDqWowO+17l46z1U3il8ppIAh7ZU/1
e9s8bSaDW8cWO+iltl2BnYcmVurOnQd0aaws+sz5VpYjvX2J5TWbUF3TYeW98ALp
FuQ3sre4tN1u3Z6rpTUHr0L/Uu0vXK7pw5nirQ6hjb6KYg013pkZ+Kj6bYZN4kHK
h7UDThFfnDYu0Qutln7tDsdqsdDW+KrkDazmKHocG0jKTsT3pO8uHX1GZ8nSGGt4
P6JsfTP9zsRZdkctdxFcrCMwUIX+xDKJURachCmaiy4QgCPBEkyLMOUzyK+geIHj
ubT5fHlhjpuCg54n700QAzczpenUYe62j4vJgILESvQMVaGOtEsK6hTMBbdTnvgo
Vy60EpRhbuPTVZzC6dhFfWu8UMIDhzZ0vbwkfQHvdbXCfu68fwH0BMHaXOqgiMWE
Q2wDq44u8bPb8hotYxBJhlfJCRrZ2BvbGq/TDJ3XDLuKPDx0z7eRZQbKUSq6meRh
gO2JxYPLgjdLGbCvFd0m6w6m1vjOBif5fLHP/0dx/HAyMNrESR/OGGeRn/HZG9lW
T8agldE+lzUMT+QrmGfj/GethFTA/bGeJpQMuKdOszzzpPNh2b40uU4mldJaByNc
tyxLjyiLbq2as0IZHiB4pbmfWO0M+m6hR6E5rKs4KYuX/OjvAqF9zalY20C6rE6r
TGJyKmh9LtRLscwBhAzaPMNmCYxEyMGhIN0RkXOp+7XxDNZ0SbnR2sNpLs/RWQye
fLxdVX9ja2zi0F4lPhL6aMuDLo1nW2SAc+LcFqpbZoK4KGk8cri0WjxVHX3IF8jM
f4evmp8WKvuh6TJXNtDV4FGwjEfLdxxjtsyGAkQZZHbSviY78IEPdxO/cmy+/X1/
oVDQuTW+FFCJGpREFjCmrnEhWBD+RMfKV4yCaWt6r5oT4gmOS3sh3kz4Fv9MUG0Q
8pOhRwCeX0khGBtZylfuy7Fu6N/2Lw2BMXy+Tx6Y+SwDQZ6moixhSvNnAMyLWvzD
eWjrEbLlP3EbzjF1vxTRFBHcQJRm7SiCAfiWwh9f0D19aK1snY+HLApWpeWur3/j
unSrVOXmTaZDdb640Nj7gVkcClhNPSnYhfix1JSp3JfiCbfwsukFBfKtlbAKvbkG
vvUsZShXlrotljQowjQ0MAr/rM+Ir9to7tqnKb2DA9Yg+e7uJCiKE3A+cgO8ttX/
xIU1uyHke5SexmoGBjAUW2/TzYGKn+DvhKCLqSMZKzV0w4o1uKcq1jql7e6ZdoMT
xyBiJGudfSJ8moeDKam9dBJFqViVLcp2NHdoTGY0bgWOdvAHblcQDfYzfjNP8O9a
QJO8ExsCfKU+sVQ53dVYmYMzorQKVHpa+VZXPPwPU5xekiVurhJDGe19UaBplW/2
z6PmNy2VcXmJQdujgzJQUmEdUKxXvObcUStdrpw3ZRRUVnD/LknEQTlamSfOsoTn
0TQnhjhLDODStOs0zEwVkrNzsBRIGQCqtGgZa1cSEvg8j3YnIsb++Jyy3ztUHwNY
Gedl32bxFKpFznLSoKLIRseEUPNZ432JpQ3J8+gd8AE1F56vtz319Gh0XnrsGGFD
eM1e2VB0l4BxW+YZTt3UR+7iwPSEYaAB5qGneNGbYqW3VmNKu2v8atoGRFdVuuii
Dmedeqy4cypVTkbE5w0EJexT/Ny3QHax0+2E/th6GPazrus44ffM+YeNWE4Rqx1/
krWl66LUVzJI9qb5X2zyq5oSTmOfqMZxM49InayCJPcy2vm8rexqaKA+sYvqIrwQ
HuJzX7ZjOnQAdqMyHgv6vwmWwPWTwiOJpp7d6dKVkoErq/5nVnosvlHQ8B7wVlEK
/jvaHfsVffEza10LwH5ndyE8mhrmFbOtcTxPXBuZ8x2pF5T+Uh/rrWhpyxNhiyMs
Ti83v8ujMYeUat5MmXMq21jnKd9WefWg6E27aAHUvLT+04E4g76jmAI2DLHP+yRB
tQ+dszw3wpYtBy0buDc/KDUCzalMqFx7ViO85NuCf+6s/akEGf+9LNFf6nBopn0i
phv+ViQQ9E2QEG+Pf0S1cd+0UwCxuUbGRqDauVVCCPptUDRV1kG4X/hT9megt5uU
CnyE1ylVQAEBnGL7PnPY6pFs7px9d3WfryJe5J68Vxv6odZ1drouR9vt1PrGBJKY
bwJsKT4O27WQxb9vBmWJDut0Xm5MW3XmpZUV07F55V51ZnKgbj0ZCN7kWYou2tDf
bCEM6eqg68tfCaugql2QxU8gxKgxo6WgWSRGVuxMpit4gHxnMk94TmR/P6ra0tRf
PIbVGV1eimHblaDYlQhkMfeI4We0Dri6JGnrH3QPfHWtGSfOmMJRQ6UbBrsfWRkk
lXkIm9/Nsc5uQlEBx3uMl1WwWXoknENO+MNkHN1UNmuuMr6vY+fcJqbUtH6ykfEp
gikYxIoBDTtCxa4iUAuxViWaw9CTCmLIwuKx5uCNRevlF9BhdyuTllnzvuQAung0
LFSBMxdmeb18czHMXk1PiwDjvZjTbckTB9jOrI9uabd/HfJc5JbTsj6ejQINaLJP
efSJLK2BJjOXu7a3pKAUomjJERy7C6Zw1IvXR9GAecONdpo4btABxn9R1N+KN8Q8
C6+DFfHl+CUyh4+eff9ufcwkgoezQ44xingt/dmD+CzocbSu7Yt0r7G8d7c1YxbU
MX6z/zXCG68MZSPvOB01T0KE4+FQsRJb2adbusrXQjhs5GYzu0XpNelnK7dvvocX
SmDA82LPTMXYSq8fsOvl2Wa+sdYEPZH7rERTpkfFTavL0ko/5iXkaF2QE9lxee2X
6FKtUaZSkDyyZ5HvjhyAkQ0sUqPi3nZ0OWR95JlOqbYcnTow1PnM/qsSuaI3DCqC
iWJrs6uV63WOeM11vHsl/J4sBT70TvgvRKu8VIZf85+JgHXSyNfp0Zs8NAzoKHRD
TCkBIEdDjedyUQy5MRu3EUqHP3L2nUJ1/bnNz3FIustSyhI4fdATTeNkprkli+Fy
FpYf8UTHvMCIKtAfQaVZXrM69DvlFfg6QGT/e81jGlntYXg4bKHsDdUjx7hwEHet
Y8duSL8LfiBP4JGzCvb8YGcIaow23BlBBUnRAlYvJfdgsRg/3mcI3TOSVDCmhfM9
rkcXBW/x4NQnz8wm+MAJeog+ti8W0MfeV56K70dr3T0FoqUbV8dfBw/QHyy3lJJc
k37FSkNsb85G6zIaS7uInpIgqHQKyN6BQAll7p+zhnPqPBR4xbdyIsMrbUMn28n0
EIhJ+W/HBMl23uwn8M8X62sxezPcakISOVrp+bMxob8P5EdiGcCSmDFcsMnp6oG+
Vod7V/Zu2DlwwNA/o9IHmjEeAv56/VLFF8PaDTleBeIfE0IY2P3lPg8nUFW4AwHe
j3GbGcGwVVx9QVeefpmHfyKiY4VUEnMlYaapDFv4ndc+3PtxHQ2fVZUesXjENYAW
aWhvOkcSbpAGjoVG9RoE2Hb1mBsIBNKh5JAc0mdgJW9UgaMOM+hmL7ezxL/cMuUG
yyhJLvS6mRNDMGfAAKpnx3xCqbA73E58TdF2OPxRG3jIjn3zzKV1GAdSCHOzrwOw
FEUkoIAeIv1Oo9PtWKU+Pkjbe1Cmberpw/xaZSztyR5DEDiQG+rZuM1N5pLtLigK
SvH7e45iCrBWecpxAYs2UU6BvTdK9kaaKJ0j3Rc6pGrLHJaMmjSP9ttrfXaxSFOI
/FXZalY1tHc95c0aF8JBoJz/Z67+AOTRmWxv1JRiHUHA6B3JqIFAEn4/X70Ck5y7
WsLpZtAGdNgayqFgPvMTWMbZ98OY4WX9wrp62y7/O6icOFqdQcVklaaJxDsWAMt6
gNA0R6cCh+3DmcX9N6tQWfGNeUl2hxN6Uj7IjHtzCZRmwkWKZTsUcxdDQyWyO62Y
FpyPM7Y47GibW94XuGFIzZlHRngYjRoInzDO3tW6nQhkxJSihox1S1uYpITuOOav
hDRBjlFVJlEZ6mn12XI2OOY5O2zGrrMYppSlpU/vwRpI8sCQyXtN2vvx7z65sge2
0Yr6uC8sRFAzJ7ITN5GxSdaHJzQBQCS7SwzhpwlG6eU2f4h1eWmwMXd0y4Cyb/Ba
XsG4c+8DiVPhjP/l66soE3iEiqeMYS3Ju+nGlyamM8YSOBjtrJQYIWsuopwUOZqV
MbfFkMMuNPwncRuf+GdTTpuVvf3qDqcNL9MIndvE2ezGacah6xawYl9vVNY4o+nt
P5hP0K3gqbgxCTE8s14xnyRHdPlQe+SzQzvYtuE38yAAjktHPBP7zdfEjcJJ5i1X
DS0p6uYzCk3RNKfhCvnljlKDyNX855dEfAo1MkyEzpTAh7lnnRIZjaOOuJfuk6To
3QAKiMu/9PY1sBOAHxKn8bGrKgwYKIh7ETNiLVd5Vhsjn/4euPV3i56oDwpu7u+L
rIu4wxa0UyvdLDpZmFCY07mL+IvFIjaA2R2iM1lxcnhkSJ+scFp+udqQu9Ey0IkS
ZL58FGBDqVBdmiLPsEkmtZOYi7siDWyg6drixpCISllWLJBGYWgSgjgDtDsfMnOf
SPJqqhfuiBSaiAu7T6Id1qUTMsH8DV68/mTGjFZXJnRiZshjaDnaBNQeOOeBdmb/
mkH8Wl6ZesGB63ZGCn4foZJf0qSbAWYLZi2zHCDFUnhSH3O1xCyAui/WyDhFIrYi
pVN49pbs8kszbt8LzC1WaFi8PvC9dR0okbfXxLn7KmS+JyRyeqihwQEgltkD3Otc
8hekfxV99dq/HbIX1suvt5gdzBnpH8xtJ4HllIhPvrKgmKHEDkJMrcXYJaqyJdig
1oEMjBnh+5uGIdm5NRmX3OqC+52bXCUtUenLOIDzswkkSNN/80lUduMPXhdgHBCz
2XMva24G1PpZW4HGA85EKLEGvRKr32tRxKkPS8mojLLH9LtWYIWDyMcqCr+Xg/vO
2BLBd5G8CLphIwl8aC6zJDVRU+0MMRFP9LEdqDP0Ne81pwvFGMQzgeYQM9rtXxtz
GsqE+Nk1/2uw1JbfKfEveAUHDATTbtZlUzOXKkCjE0g/S88LzduH6mjodVuVxkrE
KJ6p7JCq6PBhMvOVkrWQL/1dBpED+CWwar70uawP66MmR/P3maWrxIF3ulS2NJJA
fpnCZtM5vCvYVKgFyKrBzufy3bkxE7deap1uDNjEP0QEsdJYTu6OkmbsP2TSf8VA
j3NGozfD8QFY4iQuMEyk5/BIZU1oscHLLYm/Vpx2OduCnN/un608n2aCsykIn4zb
aYLi8UMfFmFEYmQOXTcNB84cge0BblJ2r8wlg4WuWMKuLR9ATV2zzzdoE7KwDQba
oM5XkDpTr4HY/5Azka1ZG9I5bRsgG9wdlGLU0ZL7wdB5ap7KiigmAUh3KnV6Ac35
3MJLP4jSjWPghOGMcEHxo3MXjgaTE+8T1j1RZH9HlbLkDWCK+AIjhl5MO8obsfwF
K+VhzNtg85GrMQQ6rsQLUNgMKLNU8Iv1Kx7zdNq3vaOBgRqbXGRqmn9bkWNr8nz1
LX6b9YrAjvm96bHj1S2PIyCSZQa8GFv240JrD1SS3j1DtLJ4Eg9T6/FNA9V6lyyu
kT+Z+6MP4GsyqIOcftnUXI87mB7OTYHrFPz0zDBIRUFNVdzGwuTN3MYoxc06Cw57
HFcAS+vixLH11xsBYrD5EH8g/RISw4iuzR0ZNSOcKgyD/TjFDwHsQiykAyWAT9FC
pUEQUMfMCFaiVoo8zcajQPzzbVSyjhboIxK1ZS910kFfUoB20WhPk8paVE9mLo6n
JLaKdrRFqBIzjlVeYnpUvJSL7B3nyZjNp+zRcJj4wXGgml9WOZbe2PcyP78rsiy6
eLPn8pGxWbpGH+dqEUmg/LGFO4TWD6x+btL8tHFw4HdoaQi1d7inCansagpMr42r
6Zd+LJTW+N02MDwwmb7VIwSsnNqCPIT+/4o+hS4SBZSdTp8SaUj9pH8ULkY3FHP+
lrfkSK7r1359HlsLfyDngryOdOx5UuDa7/jHHH3rn+aYWy+4hkr0xsNm0KcWz5Ai
bLyaL6djPRA71C5mkZ4GIZtO+OEKzSfymj/fGS2CQvquJkc8iJsb0CVsON1qVqqX
FfHkgTmwZWuJ5gpa1iJu9Q60um1Xab7e/nVp3nnTv62mh2T9e5XunL0Nf/gyqo2n
3Or2oWxXKWH3sJC9JWgEXJq8srPYbM791cwyfZIKnd1cmgo+v9uz66+KAii7d4JL
TTnk9hh5ba1yRjcaydF/93N/Sv54pXNudQVo73v1xLq29Ga+ZcrDPUn84BMk4/BU
hEOgtndj1fzo6knPJQv411yhRbfaqTm/waaQIT4cGUi81UmIU2NTQ0+n5ob1bqHV
7HZ7Cj4Vn1k1GSK26lbM78TF3Wks8/PK2sQ90pm7cIty1q2ttdhBmEY+4Nh8apI1
QRmUtYZHNMH/o2KlxnQEg9Cbq+8RrqpG+AsObkq1eqf7AZz+9l+TMNj8zFJ5JvqO
cn7CITRjebzx0GTzO3xk32kVAwiwS9B+iN6fJa7q6dfGXO1+64PakVAfpOFsX54b
A070gNMmwMADh/fBxx6qX0W/hlaDOobPPBeRI0CRN1o3raHJUrvx1Vue18/ujvNG
QTixk2Z1fROrq20qoqJZv4p53cfRDjHFpQvZBVBAvmoOorfPHfgq/cZPJg7ra3/T
L0Fk9ya7vaNFqDITfBf1DvWxGTaOwWHChK43tpBBP7dKNLVizCNLNaLQ0G4iVTfK
UAjiwS30A0PCqG+ogwFP3BHPiTqG2bOHaPxKAqwrIZAVvpqV0nHQABF3Rn8qbKUk
Mk44X4xU11GnGpfTTEpcbgQQFOa6Yt28N5GkAETKaseB4YPvS3LJxbEZTKSu5GvT
3UPuas0Y6wAD5tsdNcIe0UvCEXaAnBhqEdprZOukD22ojF6RWXj3n/P1aGSGotjq
33dMqRuZXOCSn5R+I1tbGHObvIBRT9yRCWrXpyg1r8JHVM+5nlZ4EMD/YvgnkRHK
+16dqHfUvB8/KCdCbnNWzM29lJOO26NlOhVULkd6VUBgoWAXR8YZiDWeSYwu/PFZ
MifX1Y0IvNc/hMScod6K5/RqACrOuk4iPM0ZmCNj/Sc3mVBct+RZIq9txMJM2Pvv
sSEMkRB6UZOJYu1ECBC7mqPh0zeM7QuycquR98sLUfoOVwbFv275XhKy0AWE/jUw
G6T/j3S3HaVDpBlgC4vdqjwoYziLetwaCE4QZ5pnMHubHWduTFUrsoqHq4w7O8OF
POl6h9T4Ca0hJqbNRAocEk3I2wvTIUw2suzGRVit/OtD/mwPDbsc14KWvC3iwft2
DZ5pgC7pehkaFcDeP26HyjuY0NsTFMdjMYgPe9BogR8qITbojIkF6TizNjljO8HA
To+j+uLMLde1n9NrA4k9XC2QQk5CyZUH038onYgP+SLWrahw+Vs42L2xMEO8A0vo
c4ujergVxg1dSUb8JHitOuJdem/Jgdx04i+bfIUPMWrF5JGexmwJNV4cWcBd0maI
Bz6JpQII8Vo/VNuOgdtqou6OU20oXUpzWqWAIvskssiXvoYEvFef65j6bdw5fyxI
ANJI6uEBjlw7JP/tpDhxn1a8/NRk7ruRDqyDVOWaVq73HNp9Z5n5JzihmdJzIyP1
dqw7sbfpD5YyhZXoIXriNZoYpe39ipJbkvjyjuKk2IZbWQvfpzCCByCNyh5B0aN2
1Sw8a3+GwOsvE7I7qmnucw+I0jrZkmEZfHeEoibnZDKDrKKdRxo4C5BVb0DJINkL
GxUXtxSr7xdHPoWahPtkWkbsQna84FY0dnR/WapINOhY/Auley17qc2g+2X3VuQL
8TO+scZccaUt+r/dCUkfdXjSwkbD3qazBiFxKKFmAfysPiRaQFsW3SGLtB+bi7Wd
HoCuNfS3FRLIWG3AsSDvG1WX4LKwm78UdKlfW8e3MGkPw0nIE1CHa+HQ6kP7FcwG
nD5oUNZe4dCOwanrC3E+dPfnhmTmueqpJ4cG+wCzXbr/Iw064ifsWFK06YzP1Zgs
rHA4iBP6s5aZfYfPCfbDwKZFHtqRlngVL91mCICWJyqmcYcPwMu5xCEWn41n9aKi
B9SRIZSv48jIYtU55V1n0uRn3IUtLOsgbYEilGCmAgnmeb33Hmi2DtDYup7W5Cmy
PdT0iA0TqBGZK442iJ/smX/iD1oJDvHlEMvOWPsGufWNCBOVbkYXud27CTUoK6ul
YaI+YptME0Wl2ZoEO7We5ZnD/C1/JUWvYIwdnaQXpZSi1mRew5lNbMqllI3M1ZoM
/pPkZaGM0dyGStc9iHlCWgV/hkajFaxLrigdSXtMnyci2B5Ap/a8JRuNPZ1k/Ws7
sjaDxnhXnO23YPsmlMpWBm2sZe8aJJ8a4qJOAOHh/CBgZdzfup94RROWXK3xyj+Y
bGkxEUYcC+HtO+hKY8aGyLiYHolhmZggE+CvKO5OOY9fTq0R/hGDd/WtLhQoJ5Cy
sZV+V49qNb464oqzJ0pELXxNhNiVeAaL1mm5i/exgdSB3+mO2h5DM8k6XSHS7Xfd
pLSaNFRPUI0jIEhCJwjgphnAfW/2+FHbmCmVNt793FIHpiRQWmDPMJMuu+umWRBB
4Q67h9QcPZWCxN8Z9IlRXLpyo//PMj8U/7A/mWcItgV4SorpwF6CAt42e2jOvHnO
4JbzQqB3AoEcmsUOWs6K1C1mzLGM+TuHNGfUc81sR13/KaBPB9WSgr4nzmPqIYWL
bLrrlXcXLG8XiIRu2+c+CX/OJimbG1/9GVRlC9KnHKj5FVHsHR9w124yO2+Wz7v6
fJr7K5FhwQPItp+N75TjkIoQpLI69aIBu+JnIFnMY83zZEn7q+m5xWPn6Ry/s+9W
U9949MGy5NU1tdtQUHEBw7EO9cLs+TL1vx36uTg5P1WpCAorHt3Vv6CGdPhPnkAv
kbCyB0vr+ISy0siHKpj2x9+ACJ/KMzDIrSprBkc8uCZjELPAD45Jn5nLrD1RDXV/
pJGMEFa8otc7owaFVdtSc2VlwzltwHT4NSj50Jtw6Dn03QUuSOc2Fvb08e8YFTg3
drxP4VsB5s6R+ofzn4lgCrC6RlrnCnnHEG0m9hdErYpXxTrRuvbbxtH7cmvLGn8L
MN0VYxwF8+HBmU6oZzMabOJVmxoeocbB/gnOPNsb3eDeYsNLGhubWPkXGe4I6Xhk
PZYwpmKp5SR8tbDFrSU4coLE0TxZfmNZBjWBVjHVXFj9uBhut7aBrUcyzbBd+EBV
5DhsvnDoB0G4HhvyIxvtWwx43QbzE3+fGvtW5OzHP8gfL9ZuOWC1OAJN+0k6aRbs
ippIE/p41pnUBbfH2StTEc7+4gDn58xR/B2Egm6JzR+JPotAn5kFOrbT1Uh7oGB1
UcIZgkdUPJciPW4ynuHURVJ+crUDg4NooxYQ8Ips3DYDzjXHxeIm4OcANcHzFTkR
CeZ1jagIH4O0zB0WPlSMjw5RIE7mzODwSxKH6awx4ekimR0NHRsErYaY9YeciL7L
SDLMt8sbwK9qbSX+bPIo3q6idDryaBr96cDUKH/fRQvzP85HV/I2GEFMe3B6W7GE
YxJkVXphZ3w0n1QPcaoXaGeVhf/rhbm9IRnQXzcUJhUWaFeM4v5Wh7LwpGBZ5TOH
x1HDYcQlUdTmwk5DVNbV/b7MvCo875+I/6AszDR1Nwg54NruzLmbWsGezWiZXBlU
XaDHXMjr8ngBvDHPu69mhn1stBrwL8+8+yT5jaBM6Nc54eTcF4IjaieC0wmu/CUZ
YzBqKHfhncg0fUpATXPaBFdIjfsKuB/F5yFLVZ0/irTWIvF+7Nn3sCZ7/tqpfNgw
RTQe9gizzI6rbS231hyTa8kZj4Nu/oimXIg19zWh2I3KqqWp49eqEqL0DRCGnJpc
CHsPfv7N2rLczebg4RJ1qeKoKedIYl0mZBCOa71v3s9Rj+ChSpEhj9l9qq3jXBRu
f2VQ2mL7kZAIZrBHMDncpyufEFVnNJw2IlX5zIWZcgm4npSyo3mBbezVHw/ebUP0
9VMYSjy/Idp1ontKAawrfm/oYXX4Zvyh/WcO/VAU11KZjKx3bYRUlMW9zDHm0Tks
YSqHkJLpjUAQuHyZHViPkwK/JQ1/QqHb7+V/F7CdcgdCHYxH2l1SZmSGLYZsjyWr
Nu/2o8bjy9tLc4DAmWOsNJ/zHBp7XLd3w7beHkO7XetqQJoH3lcxGttN8HWIXnd/
FaIVTsQcTNOWXeX3c7pNf7xCOJzVqtMO7T3ZDKY/HmJ7sitC2u1y2PGlPaxw+Y3Q
MLIua2key44NlgFOt/x0n1DpeBGAIa4iX4VER15FD7szqq9/i44H+sXbWsKoMBkn
oBrDHj4YpmZO/oiKD7r/NQ6wp6Vpxk/JpWJSIOji1QG8gJpFBdxsyebTIW0hCUew
6lmaq56ZwaoaKxFOFdgLgxsFuGobaDltow4f66sTx4pmmB80QLhZaIQSD2LTDR1q
+U9PnSThnFLX497viOA6cZkawgj/noGilYP3gavdmJngIowUOACegqRTIBJcQDGw
SeivV00ptvGkFuN0JeGCX/MTUBDlN73N2837REkxT2b7X+QUDntRT1/s6phSON/i
khjbAbAnd+n34Dnp7Q2khTpEhyDldRHim8a4faWaX+NBAa5A5fwnAKq5yXkcaez8
CRODrswxMgvCXS5FiZbbZpoomoZiHubmFcqUyhzq+rXgazcUo4o97RCOEAKCgxWF
pwryZ9rlDwk1u29KTA+IblZb0J/jlsHh3twsU6X+lijeYKrXGLzG+xfRk4tKBFqp
jwYqFjcaHqiMgWyhk0pHIEUlYRXBfKQ4ekYNkuEUjzLdWI7ksEi7N3Xql/eirvPa
F+dx0/+PSVw1/RKYkrnqqolxa3Nh7uKuOR9XDsSrsGJXTkafSFlZrjxyBClvQvJl
/ZbM2qVDx33hvjhJX/mFd5NZmtsq8bKnWi1oIw9tjmoI9N/YndX+SBKluiKuPX3m
hYFCNcEfolKJCr1T2Usy3eFgOojycdB/GZwGU3qEsFokk0b7sxuadaxD6aF+ANWe
Os1vHrd+JsVhfG9aNRND4hsmACQRyfQ9oBFCR0gIrb1eDQhdrfNzKBOs71qiieTR
RThZq/UcgfX6kP4iOoxA92uUmreYQpUoq1is8p2TEeJqBti2sxjViFZd/RUy4lpD
XFdtyBzb6qMxKxqnW3JkaYfBFKaM6nl0TCZ65u7s0CBH7KDeAfQffdMXyt/y0rU8
kvPadwH2G0AUUjcmJchNvWoUX/j4tYgqmcgTf9vd0hjnccHJW6hSqGd1LmiUSWW3
UIPrZX4IAoYuN6PxdrDYQftctZw5UJQC3hvHwgLLrUB+1XfkfEuzpY29PjkT6G3C
OKsWHBuC+UYw9BDGoEy+TYj7vrZmvJG/lOsuDQmPM11dVMgYqseIjLueaOhbgzCJ
9OpKGLdNM1rKwMNIV7n/fEExqr7E4eKHmSLGhj8XXlH64ZVaS+V85/ypjSVleU5n
JWQL3WhS/dLcIwdFLaufHtswKLVabemECAA+7j6OSrSYSlmnpNgaWXlVX5ScWxig
/brNfQ26ohnWhXPkPBqh7Z2brXSxgR4RXB5GcDTLEoEm2QEGvn1TsT8pBiEkvmgd
aYnlycu3kQdEi00vR8wa1evEhAzbn6WW5mD2An+Q+SHplsYijEAU2X19vGs48UZy
O4XQpljJVU1WsrDzv8WwVal0VeN7S57rOpdmqOO+bQMS8I6XiB1DikSZK00hR+yC
Ds+dYTGRNU0Ct6s9zire1R9xACZ+5f3LbfP6R4ARKzFE82hRI6b+Xuuo+CN/JJIT
HDZO9ZeDoAtP1At69lYuD6MexIai+zARys2v/V3TXYB5HWcWLaVTt1wOaut+ZZUi
0gpBZNCmWqvXZ3pbQ99zt5Z9UMpCAT/DbQXRpgMtD/ngs6vWLbGefP0WP90g/sbS
OHEFfHWuQF/NHAAJrZxrtY9wHYEU9Bz+u09ExtAxYoj9aaSGE7qrCTJbkz3KNkeg
l34pp2MsYuSDxbs6OaSxqifBQPHeBll46rKepmWzDrkuoVVHSyaT4CL4Rq0K3wRt
d2lxpxK+/lc4EYepUFcgBFkd98USXIz4ZAsg3hfsClrcpF7XCQGzXv3itB2pFe7G
KxPI/b+L7RYcqTLyTaOMuLC14rta9qofkwondmmm0vkiqVhxGP90P7CKBaHHzmeE
js/ECBZtepZJkehg38ZI2AoMb8/AbpsEbe07psDn4p3BlgofdPvVgPQpCpo0I7T6
mESSaWqPxQ3WLfQxRdyGNvQERPnaW3lqnI92nvRVkaq5m3vtt4KzOiWng9PApoqO
ORw6KOYLIlzprFTD4SHftdpC87uwPCPWIHmF31iU2LPNWC1N+t+aZ7XTpAhgGQ87
juoe+SIqulknVhZ9VnQvHrlbG3edavuNMRu8Ta1uuki2hrcVdzZWuSGIb6UEf8Y4
HH5BbmajpnE5LoqSDrbnoyPRZvhovT2wtA05wUHAbsS44D71+rjncAuDdkiQAtAI
R5VA4noIoG8I780n+JmR7wzfLHS6QOLl8s0m0T9Wm3Qgbra2AegbMWgkoCLdqnrM
c33UIS/GDcqUq8MHDbZ3L/HiLofWeq2rQ2eymXu/IKDnt/00Z5uh6VjtDCYXs5dr
vIcL+WN62i0N7WOXE7XWT4YuJe+p4jYC0ivuNUM71xPNv2iBYLICoqQ3HU3qqYqo
vUNkaKzDR7dAadyasIr6fLY3qKuoIdh50vOgPqxNA/3xAlJ6IiX0WiAIz9qDYfTR
2Cqwk734maleHo3b0iyvGhu3cOtoPxVv+0453L7tc7VTGHYzu9QfE7+Xc/m+ANXl
2KXzs4V0dUz5xHQKsFPbi8BDjBbrbBM8FGIaGriBXgW6UwJbhxY46Zlm3M0wLclv
r7HSXkwDG8rj+Zl7ZRBMkYz8VyvHCSId9xDpEAd158ahuw8NB9jst7EwAbHdrQKn
H1iHfLD2L6+B/+uJH9ffXw++pZzcL2TDKJIHOfM0rsMp0ZEeqiBwJtw4HKTgbM1i
MwWxBgWKqInqT649uRQQg41r1JbjOpChRyMcWK1bGBYRBo+Q3petEW93+B4WkI+G
cFO5UKFqhVENPpEH5zZazvtySvF/Gz68diJjAaLcwAUj2OjaSYA9WF799Q8w+L8K
jsyW0EtojMc7TH+DnmKnBVkYE7XFqscLj/vJGLrTG6qx30G+l0AjyP3MeLyiz79q
E7wDveemZW7637CJiuUfaqMdN3opM/Ax0AnNpo6MhGaeV+PeJvdsVXnrz8VRQgVL
DrS/T+WoFC+E4B7Xr8U4As0i1oHdSqjXHtnA7O/aw9B9TEFz12ne83J7fDAjhqGE
+Ves4BffcBMT4t3ExGV0+TjcdT0/o0Vj3uW08RGutVv2u0+9NaFGyAkI8HbBUQ54
INXel9vemXYNtVen1MuM+Lnd0HCp55dNblDTnCiX60Qy0v6rX1+6N9cjDYPOaWiQ
bPd+H8JjrUetT13QNjj4mlSgVoC46V4otM6yVVq+lAnpjvme+/cvV1JPUgizqQt/
x5G8sjYVfVUBtzAWYr2QDr1d8DCNDGVWsdlSW4T/5hnOHm2Mw8nUJ/PxZlfeFLH5
lswc271OP4o0+E/TpXiXwrtPrt1u0o9QHo/udphUIFkJC/uIB7L10vhoJ6dVlzKG
MoZ5+tHrBiZvv+6L0PwLV90DsckgVyPxShuLbOXnpzDkRlTK7yrSoEawZm3yGj3Y
CECVoLmHk6tSlSUU5zzj8v3WzZtKZOOoyW8nDneWh2rOU5UCxrAEqqm8c+GjKOX9
mqvSNxIZYnjkPDeldIYL62bcopGR2mhRc+T2YyBdWfNnY8j7m8kuMV3QskZ2IZih
2C9dVPedLrBid2HoOCWxOT0ICnQ6l30EXNisVr7JMK4iSoY/OqJYJiSQZPd9IJPM
2/IeVo22m4f+dBdhlRgKf58D+nJBHRhuz+xD+2HPn/awk3EFJ3hdtTMCS+ZZkKqG
3NUvb6mPYc8/BZzMM0KWZmJGfhFNw0VYNkebDOKhRmG8Su4ncVegy8g29n7iADxu
sC66QFi1zEZnBEoVxORtZzGkTEhv5Dh7pN6hmQyPU9lOJDruZ3TbOPFp/qwXGYFF
zZa1IIs4DE4Pi909OIeEqSkYtwTdl+QHo6aVZpqAAtxI7VgfgoSHhCKu+PwYrX9i
AGMp20kqv7p+uv1q2nylw9Aq3CCAzPgssobD6crhiNyyGwyQxVC6VwFTEIzBb9ax
Ytcx4EDs4f2VjPox3KBKdjA7/BpxuapxfbRwa6o4fRyyl2RRAPHW//zUdwFmU3Mc
vBUeuj06dhaFtxwKQM7cP7ytSldVDHg7uZqJadyYHF7jlZ8tjrXpmiC9eUtrbKF5
GqFck5GllHbVbllf24WyIR1Bkpq17f6Phx7cQIJmIDxOtVrL7joPzBDKV1qxz/ma
TwCOFFRXEq9l0varlfZbniJkfjeZxhdxVXRVDYut/rawbt6L8xyMobPxE4rRiYZT
qyIQBNAMSkH1wxdXy0SnKu5uKZ6f9AoCQdb19mN1PFeetNlPZzv469ZHSQ/bpBqR
Vm1pPreOSTo2W5gZoruGtL2T9jPEMjWw/j1E1ozmwGDzgCjDhgSua+M3wb8GAY11
D2lcovKz5MHcDCoLXzYbXMugGBCUBH4C48MWo/1dAU35P9T61E/zcqGeW7ifrk9K
REGZK4RfOx6AMsicSGCIQtruCLBh+fjCfs5L16C/HxtCYSCaKjcwpQ/21Orwjdmh
qCTnFFa4r913c4iBX1KP36u5r/iNw16/eEeYt1gEeDLZY27LkNUmlZEbh23QQX6z
2Vb32GWlTdGRuggts+EMPSrzdlXuev0h8IbG+9E6eg/UD2XDE13Gs2x23yMSq2j1
CwERGWyGV5nOrhYyo7C3sAh08welwbSEAr9nR10SB7b/2feFRv+/EvzFYUfagKDZ
MS3g6rc9xqHCrSDWkNN4xYPYyzKXL9rRzNwLMPdzu91Sosr2ZK8Xs//pq0WBNfdQ
ION5xFkt3MsJ4lwy6OWags8T7/7qryAyjK545vHvzdA6qR4K28AwgijPcaMQiibt
7xYi31cEx+2JsljItdcYXsbvLGcfdY5+cGOhGxsjg8/AvPxmsP2P40c/j0jgKJmK
o+rsc4m7ysopLGSEgXqec3LNZRWxKnXuR008Avv918685jzbajhTIyk22bLrKkt2
YjInRPL4GrCLjU5aoWoHUSBpb2e55X5M6FhKxsc/t4bLeQWxG5UeQfFZ128H9kGk
33D5+P/pNolp/xC03m6RFvbGcPuPerKcD2aGsqeTbKuh30fpruhdKpiKSS907E6j
ImbtHTi06sK3+5yTKJHtgJaa+fOOmM58Bp0SanSxVLv5B42XQKKizvD2bcQaY81q
BlIOEr8KALBZ81MygMDjLTnpMO3DMuEghMjqqVHffXFHnzoXzHQfmaE6PjamtEjD
1MJghFSAnt0Q0mArYRhYPVBDyX7lmFy6kxoFLPpL7N2EzoIyDuPCmTeNoEc8H7Js
9kYbx1Crja3skfiHg2uHJC+8Dh0B7b80koxyYJ6s3Nd4DK3L+Pts46aa/uDeUIKB
9ZOHhD37TVHtMRrCnMb1fMxdjX749m66mI8LqH7ovg0DqYunNswVjBp4KlsPOwMZ
3fxQkSzwptarzQgBDUdIk7e7kd/aLQVa/hD+PVxeXuzdXzd6PQscxMzb3yyvzQ9w
UcA6JsjdM6v9lbNL0rtLeKlGZbwvxjj0K0xwaH369dT2nWSfkW7YOxOzXBmrri8o
z/8wHnqMKk+jla5U4tssxOKvL2sRytkrVuet7LVuLhAkXhU6TLZDN/dzFT1Kyx0L
7ArRCddHchbVsuRuSV/x6PjnBSyDIfi4yO7rn0U5bpeX8G2hvVBJ0JJC+ZZNMRup
ehOezI7k0tlN3MMkTfwAhtWjje4viRbmyKA/3S4eW3Vmhvi9aflV1AXZb/iP6wzT
9wX9BhrpPaGRtaFy5asFqWw3d8BHoqgSuo0Bhm62pTF+POTiE8T4CtpP6TQvAErb
OAdo3gVeGTlD0M7Pjd5NieREMEBpP65FdO3GesPXejpub3vb2zOuktO7eK8J/ZOT
5e9i3NtjFgYIYeJSSlJ6zHODBkrHpA1ytVy55S98noQsENk6pdwvaigqEkH3Cwm8
8h7mfTna3lMpqFu9mXLZlqpTRSJTvoGm8k/jRD9AUuCBLd/F+BpJjmzT3CXF/CDj
M6nY/j7hvbq22gPpsVQVfcMA0sSj7/5+pDlbEMwZqKiI2N6VK+AwYYMWA29onrLa
42qe5/5/XL6qE9trpuFqz7rvd/PSbB/2icTwlswjK59AshBq57eJgM7Q7HMXNHbY
TV+ntB40L+0ByZCsAbA28uWbUE34iBt2e8DSKu/ETWC+tqkaevFE1M3djRsOJ3Ej
rW/1nNED81hXGBnP7xHVB2a3DJpZWRACFtOv0WD9Y+I9sNzii2ZMLNQyDi84Altt
4CwstsVPFX3bEQ13ik1EWv6BPWXUJ92tc8RMyduqKeKA+omUTMV9A1HZH35En12U
SJ+YoeGImuh9gsbn2ybspra8OMLBq8SLIc+K6/5zvZ1LN2iIZzyVj0crA3zL4UYU
Uf57+AIg3K9QTwDZGdJrT3WQtXr+85F41pJCkZqnlpk/nzjT6S+zBDGUKUinGqkC
xQwLlwH3EwSXN+n2WgzyZaqJgOSsGAvjFMgRFb3jBdUfVoVu9pVy6aVYTW6VKfxe
JzBAncPBt+qPG/hyaHtptOBaS0CqwXfmyHTa6IV4t0ChjHoAFWJbBzu+WL6DS/jz
N6aiQk2WJJBSWqGKBQcpgizxpbx7k/kvismajPFj36I3gQwjoW6nmswv4TnEWOFR
4rLRjKSlRLRmnQrUJsTFUGWzv3QiPILmVOFV93sz5lqJEJRR0AReCAOCEABGTriJ
9GclhoiXfW4/eUAqo/kvJxrTrVH2dZyf8/Ilbz+TfKAcitkolS65jV2CiCyXRDpz
0nhcMkOWwbPprnA4YmJGFWLG6sS8a6mo4rgvETMJQnN4KSsWUZOnNgy+NScFw74U
1hKE9s8EzVHjrz8Ad9p4bU2b8tl2gnZe39Fn/bcC3ilzWqzxTZe168Fqj5O1SHBc
nMQEEmpis2yISG+YOjn8WH9FggOim3vFiFGT4xmOLV/QEJ3xXU2mkJKevOefK7rJ
eOoBWn6bgd8oDGs0Koguk0FtMsla+esqH4LNKjAW/kgViXSZCNX7our7tklmlE6E
Qlo79K3UiRZxxGlxYmSuAaK3oBhTx2BdA9KcH67zd+T0Lqn3PQ+G1Dcu/VionRg+
quOt3OTcda62H1TwC22kNLIx8VE9Er999cz0vr2UwixHMsV5GB85x1jgwijMcZ7d
7rINBkoQ5kQH6txy3P8oLzKunBmSgwQE+g3DDWnSf+2t6jMBGm+RTHqVCKIpsf1C
a/WyA6pTAmBFhuBSutgrh1r1fdtP4u3ifhQN7GKR+iKeFtgKpLV65iz3K6pqymm7
qVF3nibrZMiGwx50UGHeuRcXLtCqcy/4OigU4nQlYtl3SeylOGq3Em1zofP6/p3A
AQH92p7zsuVykS2p475WLwwvRZu071h5S9Ij9Gfioltf2uryI4nViaet+9NhJa9b
tSt+7xC1ZPAvCCytJPXN6y8O29aOmsrcAqnQ0RZM6K7w2CLr2zGtTGJOSLJydIxU
CIs2GWueivUq0HMqpMd5tZ9wHMB7DZw2Nire8EI+Wu2EziM33uhOH5haxphKdMJ2
ZqdQzypaxeHMcshNdz3njFz6qRA2j9Qb27OAzWwKpP+YmfGVvNDhpftD1pgh91hE
XcPX8jnSH958l4xOfcQvWxjkzVOHLOtEYVXx5Bxi0il1LVFbDoHCQlfeodfbDXkC
vZuRR+Udsa884BM0SlqhwJIY9eDw+5k/5cIOUabxZn9BRF7UykxpFSTAtpSjEIba
U62unoDRhK23WaomBF1SN46i/k6SaGG5n6CKPP5xKamuZhw9joqumCiP0czu9Vms
YRQ1o1+vIKfVk0gDN/yiUu4/iKwiiqpU9v371adrcr1/75v6GZnH4MxKqEAAI7M2
fUU861nVBvldD6B4W9GNy8AgVIO73+j7Sx4ie9goad9PbdhdvvYD9KAaXR8/gamc
GWn87QzxyUXIH6Cb1q7W1O8GwwGmUoHCwKLhxrOeCcXcaYmVEtyGKX3LlscnNwwA
ldJLxaCshBvLMSj9NKFMbP1R0c+//d5z/v6IIXFcdHzj9PA9QqbLguxVV4fALVT0
JFwle/J2KEYSPZBwAm8S9Bogy5XCRJAdKIEBgR6UwTdsjwvhfgdOrUmizIGD5koO
k6u39ksJphtnn5JzUJdML3MGdVd4iV5OdZ/KjIV/u5tmcCYyyTIpR4aDJiZwUPgo
bvcnTwaNVY0sd5vhogSeOO1kLzZhGziwmodmPZ277ujaW1VCPiPg9OrRD4Q8IlyF
lg3rWhMs7rXC9T3w+pCnXsiGcko0H8oTtIqAkFD5h1I2XIgFNz4mvBpiocNXT6sW
5v58xRWSM6kuwSahLK763N69GASdeYuMV3JKiSiAC8BHNJ8BRFulxwPM37+C8bG2
LdvCDTtTWhuF3/Vwabb10hzysEmUoUDhKIx4NyeVmTIPiqNy7fOhJgte5xCLHD80
zoZtolGtd+d1OQvW/gsGdYhH5fcUnt0qT1vFm5wfMElSWpqX1s/l8UpRr/fyuCf/
TQ+Q30lk3QIReg+ekSIJ6WNnv1XYSU0H0S5Pv2DqnSUqP4iAd0kjbfLEOeJ1NUms
GQoyiPastGF3pRdRxeaFhQnnmp0wEF1tRf6Nb7S3D/gJ9nHZbWZEiS1XLwSCi6TW
UN4oleONvhmM8WBoebigaepggPuX3dHfV9GcLUZlz3u8tIuH2FkPGHQ+U5BoWs8G
w9B9pcOfIEUWLRhV59QUc3KYLyPZ0pwhPQ8Z3K6jVm60tGzrw4MM8vkTJ3AueB0D
Sv2Oa/ny1QXVkNJ861hBAHR4QSzerJre+vGR6/agfK8K6x5/EhfWyBuqlZoFTyrR
2IGWZkwuzm1754MA9NeTG9rnxvJk6vkP0FzgtIr/zNZ6RRIWfFi+RS215lJW5oFk
E9kOa774uK1bwif6bD9UkgUWhmxgK0UcSlKcqyGkM8CD49jPPzEIyJzodHancm5P
2I4G8Xz7Mh7hw7zjUDtg448J7bBR8A4MHWc4F+CQAzDKDjDtuh6BRsYa6frHs9eQ
IPSrwcx601h2Aja19fcC+GkmKQ6f/FU+MMg7IIt/Dw7E/0VFbaOZqRzzCV+h+XIf
wuDIOXvdCPukXE5eHoMhudIwf89U+YUUZC/5FV6OzArkmEPuEKTGvwMThRG7KT9p
7nju1mGZbMs8ONI+FTrY5YYGUcnXSA3UeYBAP7hcgQThU+yszWdYMUi933U6uVKB
D4qd+iFhmdMusbsk9wmf16Jv3njzt7kBJNHxidmDZlYX/g9kK7TVlTPb/LVMdhpw
xXCdo5DaRf2G8fBDVhwwpnNxZAIpIkCDaQ0msFjEuD/wh4Kfj3TDEx0vdjS45Aov
dqdwIsWH1zfY/gMgs2NK8oCCQtIpIgWXmK2GN/3Ru5yte1Zcp82iDQOs87LaPTF5
iNDyxyOAf0PGha4icHgyQ8qHb9RdM0gaHMVPNiRVLJzBs5FPsdXdSJ0J/uck5FZg
tdf3LEFBQRlF3M0hfH9LhIZ+luf8bOr13y2h+jmH/GuoSuVsPsitty5WXjMRgNGO
r1KzI4JX6kffhzoSu8bqt0CVVd7tXOFE4YvGGiFOlClPst/9JZXp6xqXVodkXD+C
L8LICmpUE0HJAv2uZsGKIs5p4QQ7ckO0UvCq+Csl0mwvC48SGErUhjnpLXKE/VEQ
Ok/eQ15xSKpQy694/cMiZdfeZn5x7RgzOzxVtJZLspGj+ABXWY0QEHYD57D6397V
rWWhgoQSBe8CjkImYH/A7aoUJkbQZ08PjCbQ+tA0tRAUIM7kqVyBJhslGLeU8IYP
CAQZ2wzO+pbKv/ZvWp7N6eWXTzbJPgf/D/dRcKkU0x2WJhpBL5jBRtrL1Wl1nE94
EE3Z5V0CE9LaWkdEREQGl+rLlw5boJP0QG3AjQ2h0jUmUtVbVxej9RigZ1J6F8qN
JtGs7BR2hdveuQZBJRkGQ2Tout5CSZh6bm/B9V5lqZNE3mse5aUhMT2J1qasm5iq
dScJnZ529UgVk3wpfCBqb3QL4td6LuTD5TFT18VD1kFC68WZtTJaOPni1TIQaHDt
4u64Bom5IJFPTVFDpfLdvO+Imr4Xsi430trp30wayTwbXqEBubE9q+EAxZh0axI3
0smL8sBEU2TLQf6Ll/84PE3BNLkZlhOFy5Inmq4fDzmPZlVOccwEKW0XlpEjvxJf
st0havq/aAUUTrBqHMaTKDhcBx6IyzpmrZBOMZH95G2cP4QoCRo2EdyUIsjYYM5+
AHdvFdNAOp8kGSS6AT42mhBHuyHbX03YQ9d4xivwFwkfKrMyl6iZPxD6dG6dlL8d
iV0F7nDmA3c4czn1yonL99ZpxDnTQB71QAkL3P7eRbJKGrLOCocFxNVWOjPPy5qY
cUrV8DQ8jc/T6XUMvMmraN+0taDKtGWNO12+2bkqeTKrko6VCxOk/mq/kfDfndoK
v0SNo96NYL878nkHTT/yryzNrWpDoZ9aDezOitoBuPGYVhpVDRlZASzcuUZZ2Kcw
QvMCPOx5oMd+MR+GHjHxeJvjvaQL7UWnM3Vc3JG+a0E1+Z7RT4NiKqc3vBKmR1D5
LNyf5263mTxS5DTLKAfOs+oV1kz9C6wjHfjS9Hl8e0USvcFId8YPlFydKaOTIb/n
3s0NjNANAiV96EWuTaVkef11ceeIJwGVtLOLNcuieqKs0d9YLThQqrnQCNRvP0fY
3Om3hiRV3hQQx25LXPHckMYmnocDeN8NR+kI792YpZA8yGqk5h0YXCA2bYL4T98P
x533yCSRfZUNEbXYNWChlo2xodI5D9sjkhN2kVVAeefbCaz124X+H9BNjJuj1K+i
5NdyhC/ZWDYg/u2JBqUQ6mjWzG5aNv+FIEfhIBceLDvpWBiNwL5J4InmDuKTkAay
yv5kJmp278glLFE1SNZeMpiKllzTnZuK/zCN8QJ8xy/k151Br8hlRK+dVWI+SbiR
2q3CZI5sxUnPNN+vRe13UDY144iqG+Vd6ohjYxk1+vOMazPRUl/cm6OLglrsS8fE
/ITJk/gbZd4jnPjVpavtMWTkdEmQHMuOVFpo+g4Op63G3Qo6tVo7j0xFqoJ+7o5u
8ovs673tqk6sLU83Dt59wM5gyRl0S4ZS6Lr0TgRpxNlmYkGoP6Gdx+VIklUqXbZd
odCFDpKn2L56HL47vnReFDkNa0+YTwvAWMO3FOj7Wjaz0/x0IAVkkpyg6kG9X7A0
KThmYlCQFaV7jgOJ6O2CR06F7WuY0HPwdIV6XNh7h9qb8w+mQP8xA5UDB79WIPYM
doef8PCz+fJDUSQg9nshEUwKDVrIepgVVsSNw+dtzChvAgkb0BURtvWBqQ0fEXR7
0i3M4iQ1CQq3bEzrNYP2mnYXyalnYKBgrbKaGbdJMi2RG/GukGJR49sByTQPjn3R
J91VkZY1BDGtmbKnb9A1hzeZpCav5OMnz9ja2DvE5PffQdVkrm7cUbiK8Tw4A3jk
3BeK/wUUhYdA62eCTZ3zp6tdjB0lxpEggKnAWIZOXi/6rENB2i3H01tgK7eGIQS2
NbKkCLs7C8qzo0OmcF9vNpQb/7aylFe27BsG7LsHczWk7q6vGXLX0syjOKkQ1XmU
H+g3PJvUFyOf9i/vuOnjWQ/JSLsgt3s6C5QV49OiG+iJopVZ+WVyDjE0YkTuPkKU
qpgkBNSlK1U5ZyUDn5X35McAuDOclIDy3CYui7q2g8mBPiwRYu9CmBduGQBdfPFB
XbT4dcloNGgbuUN49wQJ6YpvaKuITtXjoddBoiSa88eGD5bggH93YlTzD/2MZ/MV
hjb7HXeb7UElkxkzBHCgztIA4lu280qoGhDM2SVSXCXE6ZLZYHPgN1dr0zRHelQ5
//yePTEym3tS3ihMxEeeIrUN0I4WWslozRg+Vi4UNjg4wjm1FQV25WMAdNEjsEpE
Ei/P+4qdjblxp5TXoN7jJLSYyH2r84cC85IaYV2VfJhCLSu1tBomR68UX98dQWQk
Z058IAuRtjbKHfop9S6wmPVwB02t6nZL7ESbrYNoYm49l7CkaB0uqwRDsMTsOEoA
rWU6ImvfHRtS7dxiWKkDXepwg6B5JZfk4FMvvMFTBrfalPKVNbtaGBrdBQM+hpcR
wVc9FBqtfjR2e3TLfNIUHJhrAuCcCjtZASRQVKWfgeUf8Z+ocCz+tA3ZmorwP7T0
3NKGOIdYQ6GGvlTpt8P3dFVfahgtEH7jeWIG9oNef+1Pq313bx/0YgZZ/Rpn91jl
HKbGxd05OycWwSTMNsYDqEBkhYZZS7HcR2fIY62GZJpUZB4g0pY4XXkSbKAfy16p
Me24x40OHvW18DHQwXw/TBYn3eSEdG5KY+jY+inPSCZ8csrbcfavd10BNqA5qtsu
STdhCpVxtOYW/iwSqRHXO4DsWx4uyxsS51hD6ozg0pkKNzXd8+9gdvZryZHnw74T
ExDGcsTaOs4BxyMbswuD4M2uaXVKqfD25LDKs/SZIhNWSfzw5QoN4Je4M1Pf7qCe
ENqvXmfzrmHBRrapWJ3jhdjnj4246P7ivj4CH+WarStcFXE+JUx9Ge1j8UIrBVvz
2Ika5xFc1nj7iyYw8WCvBH6DqAGy6w0ZMVLtvF0rwOA2BxSwtAX6D2AhYM99NVh0
i4jwk3v5pRxjQ0rh3uQbYCMPURBzlwuAdSYBo1NZUIc9o2Ngt0NfLrtKFDoMVB6k
6ukd1xBASg6Cefdwlu4KWwO/UOMMxu9BGOQLC7TIPKJ1PwAlpOPY4hHBrP5S5iC/
Ep/T4GAbrJ35c0yVW0pNb3OPKNeVmGlSQavEExTeIaNINMzIPyYjgn5g5/MIO3FT
5VRDnupeu2avI9Ff+3DOAAWoTRfzPV26fi5nHQJkBDZ4dXCQ9fPmJamKqSkpLjBN
LOP6RMMo/Y2prtQ55BDdQXvRJykEc0339djSZQla7cJ36oKU/dVbjDNH7Iyjo9LF
KSiAPpSaDsnovspTOFtt3Vo5dihsGB5w/osTiYey9vbAdWBeDTR/BbxfxZoJ1OJq
mRkbyVNLQBayN2IyUm5aio/T/dZsZos0H19CAsxuLMDegtPD6Yyouk/3nKTkBajt
3DLpF6OkKaEGumJAOuGi7XxyyD/vHHva2ojOrugrtTDw/AnmwL8cVk/IDKJrC44J
o84YIAZ/syFzqpN5YRp0ruZr2S2vbQZi9KBdAD0l/5W1VpNiD9DjSN1dLwHCxym+
v/qVqwQTQnb5DBeiKLRQvFmxeCV2+0bw0hWhe4CL7waebLpxIN6xoFqiMz4b3NfL
5Nlivu+nDmWGP+cIrNtNHI4Kpukvie1D78xjalZda1WC8SHRnVYnpgMGlXRgKM4M
/Wn2KBVCJvVf193/i9KktbOm6OSBtR5fGrt7nksR4tC4KZul8LnCm9tw3r+422GJ
kAE2Gt4l98FORtIgvEffv6SOairbqofrQheXziNN7sXZfMRdU+tKaBrrLt1zWZZF
hMM/gp1lfPgtpJZ+EH/VziiooVlOwjjI85NJwdovydKaFNZfgw2DPkU8AUiLzEI0
h/vfTQNY1Zn5RmWo3NxqAijBA8+832Xf/IOIlFXOepccQH+kJ7mIxvbI9EPuH26r
qrkjpCvHkHcypFe8xp7Eso2ZukI14uosoHHT//BFURrg6TGNigwAEr1fYb5dJJo1
FJD5QinHZKDnoTOj2Og6r55HZLCeYdwiIuTIpooMVBPxvXV4kqTiOEBRVCCyuRji
roA+7/R+qAMM5mpDfuj0IULu3Tw94IONXsqldXX+Nd4rqJ33dKpq+2us7OtLf/eP
6hLf+HKQBpNvqLdn+b95dQCJcMg4/0wggoOfMyHePez1sZ/HDZ8o5kHaE2NkEtqx
aHa7HJLw2sdHOxQTJE0ed7nnlPn5TuhuEM9grZWDm/ZYqBN3g2nlfmqsV2Lau/Gx
xr869IYRbYe35c2GT6f3kNUJpKAAsJihSjmZ+H/NJmP3eE0W5774ZG2TRaLVgI+V
1wiM0xs6zN3ZWHYZYS5VXGIYZ0tDRji8Wl3CTnfTrZ/e/PFznBn9JeKiIhuRJh/t
0+qIrHagR6HQ4RISNKn6uWwvXmI0MHG39ACcA+aGZOB4sJ+W0iC5FvACW0jVII+T
yqBJ2FV7kdKHPzaAgXZn+dCJAPnbirsKNgweYQnygclGiAOs8MY61NmrNq7GWVKD
pnJwXakWGv4n8TT1MjQq0Q+xEjK6f2ZTHS61EGUO8Gcl32p6e2aDTwPTybaX0Nqs
S7CHem1PHKqsqhqlhHRUkdW2SjycuqXEU6NProNpsEs6rKeATEF/uyqDtI+hzhr8
wM5Bo6lm9Z2M62WNSJZzaix8Ob/FLmfp/5Fmk0Tyj0aikxC6lPYRTC+wvGmK/VKC
9cGaRgWM79e1QVoJLCsHwA7oe/ySWhhEo0NcEY6PJk5vfdwwo+BfMfsvadw2efNG
u6gLutYxkpqlg964dqh82cXrTYBoeugDrc0hHEf9y/1sTTdGdFO5boqvAK7p0pBc
wO3nE5I+mxQ8eATXvX8nUkpjElpO1Cz9G0mc39TiBk561fA7ZSFWZ+Az433Cob56
IMOgYFbZbk9suFV5j8QA1E0JfPahXrCzJwq3tKd1clRTgZ2jVxvqcFrAxRbRVGym
Q9Oq++h9KiQC2R0zKK2Wz5qvg5BNT3twInKfFa6sf70YJ/PE7kLBiKO6/zfun2gH
kLtCAsX1C0J868PshEPO3fwJELfhhWa6M9UOaidiXhcSNcJrdheQUvSf7TCCP112
0KcYPUhyZuo0HhoeRBmDfR1w68YA5diisNSonbpP7pi7updtgeSaA08WHiadAKXR
4m7piRJ9ENbVMK+fqy8XwdZrNRwQZ2it57zPT8CEOVWHjZ/A5QwXonK5Rm8Ba6l1
E4rXYoPOWCWkkTHc3ng/HdFjjp5eMCCsefaI4pYVd5Wm/dms6xp16Tt7pg4yGXJi
Tawy1rEoYmTs/kH/6trUzgSw3CVKcT2Rn7g9S6QpTQH4ZT3wVrFK2OXljptBfGmj
Z2Yjo41e34FItDNOBdl2r9+G/2RoXXL+yteoumSl4cM/MJc6IW8FaPvpJLvD442l
KfnvullUg4FlPqRSrSeCoPT9Cltdi+m3p8yoKb3dqctzmLW8pLc+bPQGTwr7Uiuj
FS1Rnckt5DUG4tT8cFKIX9Kp/+uR3JAXuXia/wcyzGjPrVimO+oVT0pp+RANQdbw
EbM6km0yBLzzcvBXdhN6mVeOewtDk3D5XLqyWeHEvMgN3tAUP8A+rufZgfAZgE17
KdbYbXhWYGFcQ22u4wn0hNfPla5lLUYrvWGTIyfFiFvHsPZgdSbIzTALVNpQ/So/
Qq8+ZUySxntL6Ogt6qxp1kyrj5fDtxc597YbFenIuaRXdVJRBWQRTRMv+hyI25+w
5TrT5pslxsSRNtnrFWHC7uqbrvTOvl4+H71HBb6OFqVWzGZR/yaKTreEISfrZSd8
VPWcMNllmtW+mrLBY3rxbNY9QE6uvZkkwf+MrcMxJ3jDr67D2/6odunEl3j/RGiS
6/938azQQ2BEzkLH8ynCDV+aAxcxhTNvDLMTZkyycOpQTm6Yr4Yzb4pyulRBdotC
TjQpu2QC/QVGGwBUWmv4cJT0ghngcEd9q5LyJag1UiAmj+KpezpXkeI3+A13FM/D
idn2knhUGMzQuK2Z6f2gcz5NnN6Gy3KeJaZXslihe8+eWblSvCmorLIqEqZZYif3
xkz0rh232KrhPvo00yVK8ELBnsqLZeHhasdaxLEO9ZwNimHMotwjWyAGjOx4l7ts
VJLSZg/Bq+FLLbPg8J2mZ8q7PIv73xWy7190PhoXtnIyDb+Ku2Z+TdK08CV5ApGj
nsfPj9XVsxCSfbVQXNlrtGiHB6kbKZK8UN1SoapejrVr4j1uI+V4xIXzeQjA7Hwt
TaX0ez/1YaXi9aHIOD79b39VvlnHGDZu4BpfV9eDTehQzL1cyMCgFF0kkshTItQk
oERUnHP50iiHyDesh11OMgxzEPSAGFjPd1n5XfoSOQKhduqdfQ/zfzlstr9JAIsR
uVP5qRJAGOpwJmbaaLnXVTMCRkWepB0Rzm9LMD/4CWtNI7XKgIZzt92lGN7X30TC
oI1lBfqhm9s75hIc1+wYqP0E28aZ2u9TZMMWXy84BhtJhKKpMemcXE+jSoUf/RcB
+XtnWo3qWMcVjb5BKn/M8ilHu0N9dk58ll/wkOGDf1ktNSnwNzIIavYJTlkD0n3C
6znzqdfETopAC1wJC2B7t7wNYnRdpWgTblIOLVHwoBrlRcSzXSfxbdu3UmBk8pzk
5/YAho89jI7IFIQVera+9IcJSsbsb0LKYeYnoLL18018RZSIKVIJfpOQDAnqBFy5
u1XEnPrXAmnkOSzlgPxOxfT3BrKnTTWJAipUlGwr47NtsCZF3An1NQmJqaXKtihm
1cHO0bovSafRBwhe4QdsbEMoWhv+xS33nHwgSJ1eFoUF0dKimp9cAwzOdz5EHhju
oo/xbUl9jPz7k9qu0vhSvQwRKBwfszWMkbLI66/246/yjF/Jctxi67Kg0IA7bhG+
fuis6XYt1pCHTE/Nhc33X4gwzsF5Jx1xpPz/CJ6lIFS10UoA+9mNDifr6/lV9nnU
p6yYyWtmik1Vq8PvYCN9Aq9o1FMNLosxK+FI8tVYxXFT0BhWGK9+ZHpGEEteN3tl
q+QL232wzLbZ7gan5R5JLg4gw9roxgrI4vdIQorih0iR/fXEtAWzhKdEbsP7FxI/
orLsi44Gi1+Zy40MT7USr7zF0t/MyinGn7H89vGXT2zfjPSJaCQmyFVWBlXA4QWg
Kb1BDhoUWNf65znucKasLJktTFvsDhEpd7SkYo3hnDOn5JNd4QYqXeNaQwrH9hHs
lI0eMH2Ehd/7ivq6zDOFDmwHCgeJNwdURTETSdcMMtAVyD3hAWqQqbehFMIR7FdM
PECuawWZ+uGhL88v8YxU7zT/H2Gb0dxwsFtvxfaKc9y+RBfD2MQ2jH/YX3KqEG51
c9VFNmLklfnZOdkQEjfybjVxj7sJ1MVY/j8g9AA+zjQFqgbvZmdeaTzlFHxlqmfB
NurrKMB9A1/3B1OEb8LZ4k55adPuLl/ClQssrLihbY0dBNoHcCNPok7zXXzfrptV
sy58S7i7Jh6tg2ddynezjjSbiSw1gnhQSdMSpXEcppfuq1QsHtW6zqGuMQ1a7CCk
MFM+ikkKsLlYfI3fDBVqSJsP8XByYG7oIl3Hk+Aavj0LXa+bEJLhMwYzQ+tY5Gng
s7ldUBR0tJ9q6hD4wzfVrLHWi+81IoBj12fEhHaez/MjGao/fii0k8tvJR1OWcHA
+JXe41HycMUkNWTToY9BdLJPDZrCT3O0prho6CJOA+htSZ96toxy7Q0khfT+tVe2
4Ug1+1stmrX75EI6gIiSpSRq1PSFuNnHuv+QgEriz1KQN7Yq4ipd96OZfNwsPLCi
p8ugwJroBwmV5BoiNk3ryb1JXlhUeoi9/N6BDBH/YomOQGRTBYPKw8NvaguEnkdA
ufk91aaDAlHRs+9fc1YVEkQWFwSu0hesa8FSSFGQAZEqISHz4VrnhXpqPBcXbhTM
u9K2atQQVAnDgJux9TKbDzCDJp7HJW5zCpzp1bnYUvoP4hjp+Bn5IKodI5kKnv/X
a9PSa4zXYhOoYea3JLj1hiqf1LyqbQTk60OZ4tw3AM+pXqNpjiYUh6sWhK92hRu6
1n0WelTwA1+9ytTZQcAdk95H38Cs9B1bBNXDXDPMff6o1deWtYbmWLdiRpC4vDb7
aCV9plZ5SwU46dWmsrZ4CwhStS7l5NfU65YEpKe3yBcmhaobwhm38nizZNi7+5oT
BPFfLQCh2PH5yUyNrnWKY2Jd5gxk6vgqVqaki8C8HDyz+Ut6VN2T7mKgKQgp943W
X2OrnOE5Nbzqm4vHfql94b2MjN5A/sCqfBbVLi2rWWCXH0ZL6lHVjulHictArg91
hSChdaNJzNOyhVKCnMvQ2utXkGpqKK2rjiSdMwq+SP3asNd1PQVXQPKfRJG6rU27
Gf7MZ+32K4BQwqyAInu257d4kdXneURAwk8wkD8v/6Sr80GLL7VP16qTD6xp+va0
il1A342Z5Sdr6yAot+Y0n/YhsWIY3vi3BE3d4ONVIyO/ycM0WEB4gDYERpmFA0NC
0G8sCkwOn0927h60edQIKtuFEuh9Z7OUVSonxnv3DeXSyv3Yn4/YcCc9ojcZVQwU
DGSRI5RFzrFSkKSi+XnzYShopwvtzAy2zoUiDvevL6wWH7wGOaYj1fzg9Cv2s04s
m0rGR8PiRhxgk4jJ7dihnVtQsypBfDAQ01Q5mB96O+q1FNbf2HjZo+CstgPFMKnR
X+s+IADEXNrUFJtp4SX+wuqsv7HgdUCB3etIBeenwRfGckShFrG1YaVRt4EZ3fsi
Mg5L0m3OEEKYj7DYvM2nkbMQwv97t7orGrTbBA/bvacdfmmgsw71h+5UoyGI9np1
eXfeLhb1+KRHsibK4Xn+ZYelXUorO1SluOHq3m5aWciYVSu1UwQXstV413Ih+hte
fWYEvRF+M84PDNoOlh9LtayPH+jKhBLLbad2eUgDlv4kRKVPibZhLzPAq2V7qfCq
ypktv+Lxs77wTea8en4d/TbTgHR/P3fYXf/oYScO/395/JIg9S1vNXRoWTJbe9mV
YZOyutDuc/1e5qmExLJasFRl0Lcfwe66l1IZax3oo+Pa1QhGTl4sKW9TNn9MMav5
JtqkJKJRiecofjPeR9uhMI+KnIvkcB7ZfjxclhOlaQtLb9BoZreM576+xiTcdzmY
h1LKRLO5yrHGBELLdypfy3CNpXUu3Uka96vQ3H2E799cV1C1GezJ15esKfs7PbyX
jrcfAgoJpK1xiQUxkQ8QewIGRwOKek9OyRDCim76Civx5oAOjQ2eSnEyYmy7PUwR
CYEhc6A7ZkqbGhRilUddnu+blxmuupLhobfm7e5/qcboVAYutgR5IRvDL0yAT2+g
DplohxAim1Ya4KVpBnMzjcoCL0GVwHVqitwME85QaeWaIUnWi/yYXbD/yP1glodW
UGWLdJdvkl0U+ihJGuoGPWE7M1y1R9snVfH72oCQFxyZk2l9iPOWxNIty/WVdJuM
Dys3qCp+myMvgaCfHdVQ5AMiq65F6fBsieZ4WZrzAkeH+y6GMrlrg2lP2co6tL0E
9EPr7LCkr2bhg+e6jRnPZj7or447viEVN/rYhOQIhJqruUWLfD2JsPwAhJkH8Tda
idIyjehaIj+Kmp3SZgJEwRpEQ7Lqm0ik6JmIEX5+HLa7TnX6sf2xPpjEDytHABBJ
0OHD77GWAiHe/yjFvPHtcL2YcrHXOThSJTiNjWTX6ipuUKif38Uoh340HNd8KZhw
nXNSCFdcFb656esuQP96L5zhzoYAg09pXQj1WhdCQIqVoyCjFaSKT6krb2Bu0lHg
27gx0vYVcuNSfV9jFt1eoxYBJBGMVxucQaaXzwRxkACGrGfcWMai+KUtERqJVGhH
Q+8Kk31SCg4BjKOURoISz/SK0F+TJLXRHhe8zzWaDstl6iZUWpmHiAAdh//4nPhG
Jx7ygj1V7Q+by0papNX+KECsmQRGpT2J7jkpIdTxNpZksw/sIL0q+8ZWaRf8pHBz
ymZV0yx/AWPkzzwSzUAQyKQw5D/ZDziRuBxrl5d4EU9iDGfXKLJRiU9rV1eI4bKJ
qfFNeHp4ae6hZuhDNbRtrGL+MG1vVjOZDeYUS43SPG8nKWoEcqLzzEK/KbJpgr6G
vvNty0vAdXCKaTnNTCNhzTi7lg6KFQ/RoLmift2eHAQtuL7/kevOlvkjvkr9cd/i
mpfEA0pAYWNO89mcuSXX5RLZrlcLAv+DsZIbm7Lqm+jzDKZUiUMF7amjGNr/toxu
zhXJqvNLCtN0gCkWeZjEQzQ1263tMM5XvDkZIuuFLxYwHWfpqhvmDeIWaNC8ScCJ
xRJOLbBi+wzm+abDk0RmmTbroks+TztZ2uLSRO2Oh1RhTB5di29xXPYDQHpEgZYL
4a7sz5V5n/mIOku+EAYHpyXkZlGJhrb/+7JrMiZMvw1g+umQNVOgY5Z8CN9bkQsX
U3LN8f9Nt0nqS+enTjh2u8o6XQJCyucv1h86m+uR1wpvaGP8ekJFrzu4DOqxXezm
REhfhi+r0/78NrGyQbzQvii11wOWcc5/pc7CD5fNHLb3v6E4mjGh05Y4V0YxDqvs
e92AA3Tcx0kKCOgG/kjJVABVDUbqCuc2VrXflRdHYHXfnacik4OtBELZ6diARjS3
HIfo9pr8AVJqqRMopcoB7j4v4V9zAa3WA5Wy5yIGhjRyE/FtfKUeTHGuKQ83S4CI
yU0r7qZ+tV00V0q7iGM/jGBjcqKDJZBwlFlsxgM6xmDe1B9LVvwmY51HJU7+IM2a
6yS1kSmhsX7NuxD77D194qe9aadl7DVQW7ZbGWmJGpIYhIOHyO34VON1N8/6e4SN
/Q7yYJaEqtNON1VXnCiBYwc6W2mUxQgFIKUSqOzFqp/h8caSsiQisnmyLuKlLPcP
Ie3oykP0TaDLUIBRfCtrgbeZQ+5wyXXlSmZsBEtE/5R/UHEJwkAg82Kg8FZzrhy+
1nNVuaUy3RO0DAkHxFLwb0CPC1CG7DY66CTnFefsNfs89N4x2zjlrKYPzGVZIR3Y
ro67V7LcfTB57Cv1iF7/Zx+a2gjYHMeLvRnfeuV0ssDqCJWA+8ebtReM0JAbtkuJ
sKyvca0PmGqjY8i0mIf/muKsarg0R8mk2u9YSe2Qoxagl+Q+/DJAFpgcYuXNgLE2
ccmGSJSdYKl3SI/WUUMI0zUkwIaigIHogWjq9eNNEibKoJmc6fwGSXNFD1U5YiN1
1N0SV/EDk05gBGatRC9JLbdRZxcnsu/jXu/SZWeJnv3e/gqkNAPvr+M4mHJjSCJ2
ZV1tOCTuUSq5uNDV3KAzpmJ1jZWbapAZhIRxfxTbYfCNI/Jr4h5ucXzzY4QVHXhN
EMHQNJvh6pGq3upar+5mTLi/hUW599//O2P5HA3tlnvvGrHV7sY36VncBTZtxB24
f4snldMknO6EpstLd6PVXrqMnPgC2V5zHZAG4SIaoqLQUp0GY/7a2eyofCFkJrX8
ZlgDAh55wTxHZ3IdY0JmQyLKfULwK0yGtwAuRHShCFvI1WLJQppDqI1xI+Pdp30y
aoJeoIaDeT05girfH1ARBAFP47G8t3oj4tR9SqVl8UcoWQsIs6aI1ik7NSn5dDB+
Wtdlc0kTpU/0Ht1pyzLNLFwHoHHSc4cOf7ziJeQ69XEe7D/SXwfe/0ctmw3bHks4
39TIZycs51dbaWqj8AVVMBzGrdDvIIa2yjxrlUCCmU1loZqXPwxNrj7KaY1KzP4l
31YfN+71lqeoK7iWFYXD3I0L4Q50jRTJBtBPb5dip3K50HkXnkEh7iZoruCXx4pt
3EZLeMdEuOCGbgErItRUAG7S1z2Fck3FQOaoAIbpBnDWEYotNeWGsZcm+aPailIl
r3tIhGmn1icJJodDSKzQiIoJHJKf2IJpsS7kn874gkLQ0H3U36Ab9UzcDLrUJYQJ
adaa22QCymcoLIMrVm/fwQAAA4FZ+3VBnlmjCKyHEJanf2BBVxfU1w1dipUWy6gn
r+Dk9POm1mtk8ydCoOXJrPWrUABhJpcQg0rmIOwlQvQtvA4mQ+2NoD26PNMViWYe
JroZWdymhyLV16ZOxbdGtiR5AbnxzUcz3Z7QnIyWMZC8vqz1/Sj6cWDCPRpB1uxx
ZerVT8XkiLQHaICQ48/qDp97zvU/RK6WVzh45Wof8G02WMNtzC8vX5QhmPWNFbkn
A0B4x9I1f6Rd6ybvWQgLJitqqrsyuScPHvXWF9df7kR8CF71iNtLfPFeC6dQo8Yl
2cdNl0REHBzHpga1TfIUg1P96M+23qbRj7GUp3uATXiN9/D4P5MwNG3G/Cy1wagy
MfEe94/bMrteNSpWRPxuL5H5MsPX1DgVjJI5Wu7BACRjbP1xM6gL85w9bAC3sSUe
xOmZOgCIXuIks+trqwGomPbECANrjn3/d+xm3/8ANedarmfbCFkvwCyc/BPX4Bzi
R1xj7936a0NPUZl2vAlpLeT3W5uONbrUkl7WBoJsnWNWAEq132cqtnmrXMQzacPc
RAI+9p+f9GQdqe7j9swE2RI5CSXJ7k7RqmEgvt0htA9e6yn2vyEXwGjaHBhAtE7X
pXCCAcXiNHY+no4oy3AZgfzikSeJAZ9GpgZbmYzUCWvvUIUPY9ocJZW8e8uT9icC
LsBGO40EXIeVCZc7lwq1FWjYo/XGebg4JrCUCNX3Kjt+qzC01nNM2/i4EFA4Se3J
ZGdgsLokEnuWdpBxa7Mbcj7lQQ/rO1BbxWfHdm6aWxSOSdBfM3TaeMRyLl2Fw+EP
4PSOrH8Mgl5bV1gFadDyXQVrUxz6m66DzOcNfqXt5tl1XGYHdGBGW6norUnik1Mg
hX87Vi1mMPiWBaQiIjQJeTr6qb475b9bMCfquoP6cwGZ++4wzG3K9I1z3u9iGwzn
8PCgveoJ9p0HM+C0vp3imEajVOyfgkf1dwEdbpOhAAjn8DmAZRYG010TC5JQEASR
KS4AgCiT6SLIcZVbmIhbJ1n962IS2q6WZ3sGdzq18nzG2RPIsgeGocpEt2xY3TLF
cAmeHlR8dTG8F2aWInTdOnlisR99EIPtROSINyBNdq7sGy1IMtfR480ABvQMrOO4
A3Ku3Qydhw0y3GafNux+IkqLJy4rNmcHJcRHRcCX5ox4nJR9nfggRYbL1E6b6QFo
jCogRQB5EiELw9ab3hjMLMFskydpGaS49O0jY6AFvRHBZxOrYg2T6+eawxVPsGBQ
OaV0TVN8xIIzvaYWLyiqvIup+mkSw1el9nHk7cyQXl1sBVDg3NM64GAosmqVY5ns
MrZBygGzNEQWWPyAO2T6z2088gBtXD5BzqwSVIcyDKnfJ1Y5Rs+C3kKc3zPqCGhf
fiRHUc1U4WDnYnB9EqSJTpn9WVXRd62LocGM2yMClhKgUh1W8JEXfVeKczkjyC2n
QGZV3PRzF9QF9pUxS5tlKnoRU+IG6NfF9OdQu4LES2WaZ/YqI10GfSmkqHkSQpOV
dnzPOzr29yUIbPqz+hNXSmAhwfpaZpEQvqMwOeB1E/2pYYupVLe/dT1m3ta3iKjX
Pganihc8KqHjYCPFkTLzjVmBDG94s7/n1WEnprrXGsh0gbQK02WizeX+v9qs/T9e
82VaMR4TLzqfCt7CwiIgjjYBqgXY416iJsuEMiqbchiYUysa9uw5luPvq7+qSLXH
BTIhLFmRVnlZwmleav4y3OkQlqNYtXU1lp1U2+ngZzgsVEAsX2GSbBzybKGXnaVN
SN93YSlTyDerv31cmMlFEqwp4gWSepyL/IUyvuT1CB7zjaH5xMr1IgFyid4RIYd7
HdvTXvxkJR+e10f9eOi0Ew0oNutXbgax6bL16g0CeHRQ2EJBEP4RiFzTxCC3oK7+
lrRi5BVUyTxw7XQb0vmj2yIOr74iXnYrWgo9C3pIMKASmUi5AqMGidQxv7g7ILWs
5btHlHNZwvw+uVlK1giQyfMnKL7ffUqOmK+IL6NzKKUjswxNTM5k/1WRAIhKEnnx
Lsjus4SCECT18koEfH9MXFoce9jLTq8dRI7Q38JjYs8hik9lD/lz8Z1hvzVSx5xF
b3vAh3NbQQp0AsNdOOEDAOv16RnKkyS3kdcqgKo0Exj8/PlUM2WY7ERfZ1JPmHlk
9TOPxL9hTqWLv02zS7TupDxGNmUMYc+V2YzJE9/dlz9xOQr26vUIJsdpfsR+rEtQ
Dng9loq5yrqRFPcluSvbj54/7tsmR5Vec4leebszHyTUOC/mQtfvv6eu7I9qaD9d
vZKiYR+FMWh5gDfdzuKGYDhcL51fJPFr1B2xfH1zS1FAbFOhWKAGQQQgoPnvlXNA
SAjv/mqiEhv+36AOxvWaXKM1acCi0xU1mp4/QfbzuwHhPwkT2bFmU3csef4os9DV
0OjZ+tIKycc4AGoZcZjDLSQyp9dbKsC4Bb1Ln71zQb2tSEQZ4aHkWslnea5LA26Q
xG7Xn/MWjiFWUbuuTzOlCHoTptGGgzdwKvNsv+Bj0EWjiYuDk9qvuZ0MkvYA7zvn
FItGRTXh9raJki6L/aOCXj/PqRN1jPUXrR9KyNqacq4i6GjHBLSVGDYOs+7QYtJZ
RYrQrOaPPj0A/sGx8Y/gP0//dMWVpRLqkST7Wq+57ENESmf9dscF9G0MNlss2tCN
RcD4OfHxJ4MReARHwFoTCjWVQ6DKmaK/Kb2nAAr0oLJtpNWzHb/fKCmuV81B0eM1
QC6mtdn5jVBTac/vyEI4mvejIOoHGb71zdD4fk2J1FbDqvkDohS95MRY9FduIzxq
BIGMxj11n5wwDKq8ek1GGqq063Kb/uqKtozsK8AkMEajbeMwHIbuB8UOoTpTO53s
zLlTMaBEjNjxtXf953kG1dZ5OEhg6JTBPpj8UGw5gN/m9UeFlXANG0hBqxPHV2Li
F/rRQSxuIX+JT3Zd4uBaYNWIqbdd/iDKUSCSfOGoFwPdiwBe4cA0A/B1m+Jd+4U4
4MA8ORY8g3TMB+EollC6LpjcIwkIL5BgwNHkc8OgrxHWs5alK294rMf7z83zOCVM
lWytRI5LTwMr8/e2iSos3R8GEzF5wP8AEq0gvNaPrUr3x+kunVfN7Xn3P8juCMeq
m6AIPCuqFwxrM3qX53HJXGb7y0uVxnm4z3eviM6T5F2bbuNTU9iyAeOfW1z1DmTg
Vf5mgcIovOa4+nu51/+AZbY/oksRqtXEuJcPrTt75KdF6ptA6/Ti6WskKWZhUMLN
5SeI8myocw7R7Qj1p+sD7OhbrxPw2wHRfeTBfRH9o2w5e7iJ/Vz1hl3cIsDnKmQ0
2dW86eFq2NdF8x7m7Yc4cNy/GJeiztVRs5UokjGB3DUWaTE+O6TgRQhPtApCCA+g
Ope5vxngevpXjbAFCnCDKnHJDkAE1gy3AB1BDhdoc7WZ/8v/FrpVR0xvbdMsyBUn
eOwjwOZCWHqcpCRkBuxD4ZeH/MUSRqSeA0Eit/1snbsu/Jx4tccE4Cfygjsf381x
HEr/t2rQz+sqpDZx2pXiCsjPhjBcqaq9lM7YYzBPD2ilt7+92gXWSg9eskqhfPXF
uDbhybl4pbOcvGNCqLCxWhiv46lLB/OZBC5olzwdrdH5uRPR5fAKnHlbzpKTD5xW
97R+gIjxSxWLQQv0SDknNgY+b+p6xPpm1pTOAOz9YpjfZAgTP5jJIBRlWA3atJDT
RHUN4tMqlTAg17RuunK56IyNLxnD3R9RRLsEAKxwKrS7vMgALEsnpC52NCKsOIAD
iuw34UVCinjYBvKv+yEx7Ehu5TlGE7Syz4x8KSIv5kkGgzeKmTu74CzqjPHsOXIh
uIWBaO7tZXWPzK1nEzN9WrRaqcOG2mlHjK4K8DpOBHTaQv67k+ukWbU1ZNxlyJW+
cB2Y044t9c4dNeg1QKgxaKeALypn2cOdnuShamsMvrBn5+DqV4XGMKRONuFht1Ae
zIgWrTeqomMQdeWcXVn6yaqGCh4GI2aLlYncSPQR91kslEfLC8LTdUKmG7xF+lyO
LWa9u/Fe9SNSAB0C92XiGheaeMCeiMbJy+G2PQqn9WP8PrVoANf2FOOTO3757uiw
K9o8wnE21fSgDaZX+F1TQbPqrIbrzfqARRJPZdxqCgqYtcd7E4CtWYYFgSxOrL9R
wwNDKSNGLGLgUlV1uaFF0brsAfkfsfbX0/2Zch3lDVDgM5cDsUA/UbA/7uvctM9N
AcFc/SDX1x+oSIgNgmQBAn/KSPnFgCWyNpLuWEjwXhsME2qWgGMW7vlPCvoFc5x2
iN3gBjrc/+FwfQRrCIUaPBQw20fYmSzK5ZS4zFKuIvHlrW8ZhS0Gv3JlW9NPXGJX
mxfXY/6crP6P/YN2AZ+RZ/QmoJNKMrbwdL5B/6n3BNq+IQnvsOMSGMr71rjz4fEs
67BrEg2J9qIlOERJbnQhYQov3xlBHE0fg8dTNvMWk684a1wvR+UNn1DP70yg0B8k
drj5F1X7oL1cjXczjcn3rPGd9/Q9RgeLT7P6kbJIkQBiaLuKMfomCflLxmOXRgMh
3BfIcMjF6Pdoh6AMUYa02wJuHZDddnO01kEyifclEInMeMLyLJ8kLWO+A8d18W5F
niig7rTLOvszwdJTDnqCJD9e8gVFghg1AkFSwqZj+m5zJBICLSO6uSIZmMEVK0Nb
LVB3fyvvSV6NAgA6iXIG0jT50remWLn6P1ZVOAsvsv6ien+7isGCdgFDlytFknrf
bVFvMFQ1CsGlqx5r+iCUO07wmIMGUlNwIVekbfZocHZvyGryIJnQWE0WzMgS+bt8
7ZVe2UMl3xDBtt2lL37SLz/VIghXR5Xyts8vNPZOkIDuqZClOUBHJ0UvQ1FT9FIc
woY8D1TZbjvRVf3lmDAszONwsY/I02NkvqRYK6jLojwlc+FI3XB1rjKG9ybtxWog
Fq0KdEuR84w9fpGz5gX+ijXvvLeKflPnr69jr36TeuOEbN3Za58lqDHX8XiEh0PU
k5r/Rt3Tb5P0DYFuMidlAeYUV4Tz1CaF5krunSalxrgtXcikoClrIkctXO6HfDe7
hOsSXnU1lpvOOMcT7ZX5fGe4xVVhdlepsSoG8s6ctLj540knxh2qdJVxgJKFahpx
kCZYBDnuTMTjoGcjOF1wLKZSfmGAgNKCw/Aug+e9G/ATy/6RVYOxUDruclNZkjBd
IVJEwZtFvcI0W7fUhmKVKEuHaTQomjdESDYTTh+s2L8/bfuGe6oBJH8BV1QPzRWM
YaiYgN2nhm8bnBHj2QHEdFfjZ/SylUhoEm3SmKM/pndIcuRIyHGFtMvQLlN+nCaE
uu3gblPj/sVMJiPHQeCbnbuhydBIpaxaM7zIWjGolC960OXyIeA/xsxS6on9EBTn
sF7aQvlxK+Hz9P2vdv9xOxMSAXsA7kuz1N5wpwrz5gvlSa3kQAgSaL1iKSkRUVR2
BBChTJlkfIexz1A+zomffSn6nkzL04ViZnojAb6y2lrcuph8e9sAo1Y+umMrwzL4
ElUH/URXr4eBi5v2RF37QHzqJwtMWbRqzz6+ODdNTpXnDMv8Vab5xouaDxGq+i6E
e5AUFkCAuVCcz414XyB/XH716hVMF1BJv2A3JHUAQoE2DqQrB52XE+gCzBzC8wxO
Ds7suCWfZ/AbwmCJMuOEPvuLUkHHmIP0vFO4Jl2Xdsej7T/WtaOr0Wj5bwzbZRxR
f1qgeswkeQ9LKTqTLC6uyA6SCN+O+MJ/8pq1jbwIsTKYxtWrlF8N/HpV5whA/mhZ
84FQLzI3P5KIBOrBMvvSt2Wr2CtDn2tdaPyRPVKvZtEh2hubRn/0Y3w2AKgMnPIb
F7YKLodatUIkSvzcop/Fi7TPZYR0OnHWjAd0nBbrn6fobHTsZbFNI5lj8JEdb40q
EQ25RAL7h+IRZWnoJ7RKrdFCtDCRPihh2eFWv5fFC1elCX+wTUwYtRO/Iq+C3l5o
mpVjTwiO38CoDH4R/C/1rwQH935YY3RPhOWorybDP/0AqioytLDEZJWr2YLJC+4g
XQvbHjtAdi0WQpd5TGpVIotD1F+negdFlXRPcUFjIYKO/OO7nWa91OMmC2I7AQJE
PqndvEdTAc7jQtIlhXqilqmqm3hFAy5yplhLrXnBgwaKiSUaeCudllvg/NaCGUg7
Y/im2kiVOv9TO5oipCgvCM+5wWSN0LhRnUP6s4zV8iJbkevsAC7ZV2bnnD9uWFa2
Bs6tMM+AYyG5Fg/z1COLKJGtePpWVjvWDqVZZCeXtN6U5sq8NwCopzA6TDHuQch0
CyYWU83OnakTT6nfLkF2fL3Wxz5ZWa+Tl9GkZGiGBZkZsxj7mFNPzsAg8PtE9SAV
28lynkCJ3ioIBLz7LUdO+U49Jb1eT9p/wFsRlfuyLLncZBKE9OhBRKX/w2ClFRnM
v0RBlrEN16nP7D3jd00zYXWwBxAu0prO+hWHbNjxw0H9uNrYL42VRy0mNVeLZ2dT
6V+sZ0ONs8pi/+e4wVcZJ+RSqHr4R2MeEWHyCkXI6a2XPMYLA0JGrCRDnzHAtpTN
ulpVOjCxxRiAt+kee1cjgiA42lWAWn1wtwQfgjgaQe0NIC+dG/GC/q09fsykeBW7
gAQzEVUXEItM7hlx3AaoOPdSRnEWbxe2I4UhczNVqQhjhf8+Wmpy90u0KhnVKPXA
8AGDkF3ygiN0y/cdiRdDXRquDpJHGD5H40TNsWp/pwNgYTdIYHxhLX4ZAJBYgOr7
QYBUft7bh4SrDFNskHXOwVaT35e/iViDi+AVRTNqEy6hWMWDdp4dQfo0P4QuVDaO
sT+3idYAIkkPSrHF59hHsebxXA1ocoHY4AgQRtuBdUUqvMslvjPNdUZltrrSMwAM
hw6Dw21qHroLFB11Uch6Vg0NvvoXfd22ZbqWUmY6Tbrm4kEbW7AdJ1Wwq9AsPt3D
TyWeuH1uXOTBzGwuucaYRtGkjRwrxqneMXFTrVBt/ith45WFk7XPmltgpzhnj9Dx
YFmQR4O/KWIqqH/DfYvzCPGPbmqlOwgeAEFSKJ7kx02rS7MArhXGxzWLlPmigPXT
Y5T64mb6YOHX2MmiHi4nqnHrRz1LiqsjVijdBiBGoOytFipRkpPpBjcX9qD8Xkyi
lS/ybDdbQPGuGMWjdjAhGmtQe01tJMvt2JA+ejOFkoVLXV0nXk9FB4fo8BhBRJ+x
VBg6EMuSRV0VgfP7EGB/HBkypkZ1dlj5iL2FrMuR25wjOrIoQif0gKSW2Ya4x2IO
FZoGXmqeIZpn5OVYGiAdQZi4KaPb5W7n6TqwT8RUeZ6fZTbKVzUTaYvcn4WgB73R
LthR7hEyKWT1xkAnWFrYCOsjW6K+BnH8phVAXIktBo7UF6lxcO/9jpk5rdV4/AE6
AT03RgLt+up7Q3NTVS1JL0NPzQQm1baV5IsnkU/lHcbwvcd+twmTjSdAYQj5Cjzj
pHYwf0HhXfHJ7squLORQlt1t8AK4liPgQJG+UW2KA7unoaDgQk/fJhH546vZIcM8
2p48utJj5G7Ohiu22G3cWGL2ALYZn+A9EgtkAVW9L0hOnwQje31AtE0MW8tc70yq
JD/ZsBzV5ZPdItY/8sekLoCq76fqT4vQh2Yva2/pu57U/rT9sYZxRHtavAkT7wr2
7qSHbZ89urz+NZcRhQr4yXmTz7E74ZS0XrdV/r5PbJQdhKSHFFEMvso8dqCnVg0i
oJwvrmnNZQGNzpY3pyoQs5KSHYLCr83Z+ghVPQg45RPoxRf83AZ6wZlgDA0bMAaE
t8/4elgsLz+nL4B7tFTqLamsmBSk/K5348Bk1BpF4brRkIxEhyBzo1eWTqjJ8Pay
YoxaYziEHSjDugka/tGp6hQtLPI9l4yIfvp2dnFdwIrGSIJvCdcAji78+AC/FqTb
zusFkFPGdCk9/FAFq7bFhxC2UD3760x22mWschdrOz2MjDIQ8vxSlwuoUgsyUtdi
d5WpIzwvzrOZQmdA9NmI55cjQLFu/53rh9c7iXpasGWr4zEOZe2wWpLfVceY4IEC
TOfTJIYzPVGAHl4v4inJseSx1DJzYHfZ/jXoomdWGtrEVEam5sEZb6ppEiClNEBF
v6FswrF7jgt+FxjLDTYiybAtnmGa00cLqPV2lDgjzV3IdELxvbfBlAE/3swhnsrg
esMLkpLbgZgSs+BjLYczsnmEfOU/rNjFR2RpWEfkCwiz6jbTydixiEIWi7q0T58X
603MRrC+p36/0R6Gm27sMYazNe5BYR9kPkP7eBMSYks6zdFWnTQmmAYNI7db6z3q
ozSND26Yhk4Bkl1C1alnD9sZ5IgoFcv//WoCQbUvgdUsU+b0NEai3Hek+K1XzD38
tmCitPKQTgmsffV1HQ2mUEjcAJ9OEaqLxNHpTS2cTj91WPlBpVirhJyTvT0xR0Zo
3LKBpMB0zgGbbUYudzrUz9x3tIus5pdYkzfFrMEVIc5qUwLxqL7evscQN2nl/Gjb
5wBB8R1cdfThOmSMM88jdTXoIu+TEt38ug+MDXeaLCEmKVIkCxt7Kq60CtrFVf/m
Lf/fDbsK8Uh0/NtKyUAlf5yZNzXeJf5698Ktf7pgGl4WOa8jL6UMckTXP2EsQOie
x51UFdki8NE+Utm2aH6PQiQgVE9QOvoaJCvVy4+57QpkXmC8y1I7FWjLjLcivhLD
jWJheSj86/QkzcufHT2lII6a2Wp1fIc52NvdSII1z+Fen01S4BJ5zsMc2bnIWcXE
pIAEjnBfWoMs4AWXDdyUqu97w2ce+UUdEl6VzEfM1JGsv8ivR7Hws1/aHswYV07+
15Gf5Da45gySjYgBjXG3siBc5SuOMKIdgDFH22Rr0GNP7ttqOWjLQvkJe3aep8bZ
1wgeq0beuZWvjBSVJ7duZpXjGoN0NLTAzdlt77w5Cm0rxKUOuHRcrtdny7wsvn8C
O1BHGcrYT94i7vlhG5Lhqskl5PFO7/s38OHhR3S/WqWrM6Zf1qp3gzA2EqCQ3w8x
bKFw1EXmR2T1TiYBcSUmLPjb2UavQaRQ/3UOFdvZ6cIsT0Y0T9j/qw/ckPKpM5cz
BBPgJ0O3qrhSTBlhCWMihX48vKQQayjzrAjeGcrv7zvjcMueGWi/1fZ7o2oksMrO
WiFaruitWQy29RatPc+dNDtEd68UPsFOhqUUB66hvM1R2DbY3EQMe6k1HFbCN+9L
2Ke4CwmcoxgOZhH5F8laLOuSTlX5THzaI/6Vqa0BGTphg0F2A0EHygpW3Dd3016F
47OKXXnHESSbcqdAA1Cvo5hmStl6vJ31QSlvNhPPHTNTu3vj++Yl70Ti/I3YQyvh
e/HmJmYwyT9xXOjz5LdemEE/UHsW4WyTVFqvAIte4YDA39lqXNpMUxG+7TgFksoG
cBJwToiDSoSoGguvDvtZdAE23ZLOSWKzWIzYVfsO/66IKeShnpkmKblfjdXp7mK3
V8k/g3MxBBsn0oN5pKMdZrDyeLrDvXZqTeZafLD17RS5kI6IFQXFlkngB8DxlKHU
8emRN5IfIqvPCQZiQNEMaZ6aNzjRWMx/oyKRuE7slYFacgTGigBmY+qx2ehxos1r
I+NjCXBtrPLbpwe66c8WTe7yuk19k61i4K8TFRjiVvu3e7V4eZQEj5yUrBXxNYp7
V4RQfEn3IfNAvca9/ylLPoD1eFDfsFCKeF1arDNbCWgq19yt5uapy1IFgahdK0tt
UEKVqCGuWTEN5J9SaSYGh1Ab67y9v3Nkp93r14BVdRUEqidgoGv7qK7pYY/Jc/SJ
L+Up0JXGuY/bhNErDTCf1VJu1oAr1PWSrN81v3dn5QzoF+svJVFc0OwFV6REN+v9
RZlTyxcd6GVvihevXGNOMNQClPqUokEiWfrbVnZxSWFaBxDELa7hW9xy7SpeMXS0
HqN3cf70CiZIwSuWGmW6CoukWR2fb6lnViT5kM75j7jOttDeMut4B0kPqTfbc5Yn
cywmoB70MzVx6s+fUCKGG4FCo/Q/PWNvOspux3BO30MEC9q6wh2Q1FtdtD8zlmvu
t2Qcg6GoB+afGWHwJH12rQ15NxAjUZMk77a9CirlZnqWzArCQpSrraH8QpCSSNdd
uU3Eg8DMNJCajOIW/x/j14JBX0l/WecT2RWXFaXukcG17hdFk9gZVUQW+IWsm9Rb
ZC5vjzYdsmXbbXWjUiSwJdSB9j/F8g7bm7U9K1nGo3+tIsHDjxpal2RuurIOBsMo
4INYf/uz+/KevmrMYKmo7+c6j763gmp+obdINOKtJ2tGlY2lA6RxGRG0L6e9lFTU
xZZZ1nHH9ToGLcLay3lXMUh3HnJSDs21SqOLnJ/uKynh18pIBpDHnIEY20WolHXH
e5wpf5AEkO7Rrj5zOlK4izkypHCApahiBUFeoqexrselJXz7XVPE8DegVb3xio+D
4SuBtDBaTqDs1cCL9YJectQ3MDAbJOJnfAr67kUBGfwFMIQYJxsnOjSKeoEgYiYo
w04TcOJuubRPA7hCl/6kbqs5HqOK4WmQoZgiDLAMpVWkLr9xkbuW0Z29KcptOuVp
GzeRxnYi49nBrtyuE3fpQAfmWVs1WiXE2E0Tyz66c4kY4SQq3/fip/rbygEz+4Tt
xyegpSBMuugq9PMbIW/e2yqYBLk67WHx1ujC6F0C7ApoMjzmQTud6tFp2i6Xs1fD
Sik5T7rfneOpgx3p65XfpQR3IZN+ZeLetPmLZ3Gh9u8YvqVyAmj/krWSXaAi4zLs
7QNZZpASkeHMNW7A/ESxj3K8eL2OIYsG168qHmeQLcYJlJsVrny/7dDPoknp95ab
rEA2Ly1F5b7XC00WuWod2Az+DAEpiEkIB6+C385Ycuun1mpE4Ib5rxuFkPPYsfa/
GoQxFfrdZgpuVOA64/a3jAOTU9O6n/NpQ494fGFqOp3L/xcsEMl3r8caGAsbuacZ
5Sy3Ussh6Fx0/SGFy4/mfnXmfa8QPRS1aUbfQFtahtqrxvaFBm9aWgFjVdIHMMpT
Zh9sRu7Fu+LmUITwONs/higG0ECQFnNRICd1qT4n3+TotcPBKNUiaoZs1AhfFQYG
RbA+RqqVj0C9rZPxSeeI0zSyXlDCGVyBGp7xGxv7358RB8Mb+fb99Lkj8mIdNI0W
yfh9GVLJa0Pr1XVhiynuMoLOT/MsefBylbcwmFU4P4NlrpE2oBbIKGoCyM7rsvOq
L5kQL6q1JRTYctwR1nYUw69SOcJtK+WdsOijjFp5kgUxzDWRXTmUEPr9jQinYwEY
HacdJ45XlOWIaujfkoi1L09NyxivHMnXE6Zb6JkuU43vmYyRm0XVNa0vJN/2ImkQ
nE5+naSrwMBCZ0Mfgw6rzVdPn6g7dUrcM0R5LrajdRvZCzg4aGcRo34kE5Y6kqGY
IzilxmjNmshyBzsWQcCsffkkS5DXHR30sOpYeL7DnSPLffY2W2ZJMMidjmuhCkyN
NrCuW70RClEgMIyHiFgLJlITW1FEmfUzdHpoiEqhwPLzvdDfOJC7aNbUhvE1woIx
CI0x0uq08qQN0040L9ohzZlehEbsRapC/NpcIrr1eGE/Dk+a/SGtRR69wZ/oB/Ym
hGB8TVwQ+b7sq8tUjc4kG+6eARD8LSfAEMC6JoNc67FLbZJSCgaftDjH9j6hGL1u
nBzlTI8J/fN+H5HczC7He39scy5nbFCpIDLhg2dChpaCakuisW6aDJOUED7K/pvN
SLMhk8SLbc3aE/HeMMrCRRZjFN3VtC2LGGcSsNbFtwuLgeUHUB8QXuaE35xXWfu2
MTWDFO/rQDA31vxVR/TWrL90zhn4gv6rVP9AaJFZ2Dm0c452LLA3KI2fFayFtpJC
WFto3hB3p8TXyAa89ZROZBgZ7HYK6BguZbR0OLZ9qsCXpBlKsDaqUGyvfreC7QSA
Ig/tVUGLIQQXJaJSFm2nNSj6G+AEXh1cOacD/Z+I9IwDVSo+XfaIIZPE8crjgWO7
aTU7cO0sGl/MkdMi/NrSAjf2gLPsGDZl57pNRVUZGHvCGIvekLtnm79ZKY+b6zm1
sBNIWXEffv2Ka+e86GNgyS9MoVCH7fO44IHwzfDu+m/FZrzYusiOGapXN+mlyeiA
5yyM6ZJTBX5XY33KPvO558Q9ig5JP/3wuRRjh3M0SuWp9sUaswFtzQNgkDCpgkml
Rot5VIGb1GmvY64Wb4aNm3PwUb5AJbxDmcV88IvpBoS1Vp3KFyddwHkQGmplAUD2
FQmCfpLEDSX+U0/dBA7twixsH7ZaPOBxqi6ghPpq0Y/mdeNKJ82cls3jgcMA4UU1
HDuXOXEMk+WUudF9bvop4RyH9d8T6wOqJikwiQeNSDkRJzM+/DZFOMdZAZdBpPWQ
rVqW9m0+9JQz+qlcDSofybDLzX4KulXsfRu9Owm9NyEnxgdMrWcT/Gv6KpCWNA81
MwgFf2lyTrNnbZPkf9Q+zhoKDVdmmrxTIhfjF3rJoPiQUM6DboyNGaR5bfjG664F
wgF257pcrzNKkzl/A3k+Aw7xoAbZZd5pl6ZMfwdYPDpCGeaUHnRffacaW6mwMSd+
ThlR0cE9HhoG5W4m3w0zNu3or2gwdpG9Hted6aomlvfKOq9SxyqoJW1u9bYV+SR9
+pRH6cgMoBBPJCCwpNCq01Ohq5LEFC2Cpv8VsdumcVkWymMy4XrdWgmk6ixsOGWs
YXFU7mY1/Q6xp1RT8xZ0YTj6qG99VT3snMZr0uJaPadsElO7cc34M92SFCZfc4CT
bTm//R+SdUhcjfueI14we6CTpXXyQb4VZt9fkQ4ZSXU+iAoeLUipk2bEkHClEwX1
MNgOVjklQP1GB02WMCG9p3hBKZj1dvlmLYKiftCte7ZrXME3FbBDvETNotJQUEur
imG1Hf/DoPzEpFReKIU9BaywvshvPqb8+844Gjl3N76LWLBDqeOrmDgeF5uuMOic
XYPDV9gquJMnrhe+HbR3wNr5WzprmhooFwweh5yl/PbvWfOdWg4LX8SHCnBlUMnQ
yawXlzO8m1KpAldp0CPqZ9fce2fo3O/tDPEMh1Gl9rDVCHx1HDkA+o3dyPKgGxbK
K2n98Us2bGWbj6aiIltUXj430W5Nx/bRwrPqBuoCAyESz0vTghZNpgC0c7UPJZS9
ZyY6CCgdBceBCb7HjN+QBilSei16Rk8OTVdkhqmpK8hvMIRwPJt5Rsfc1M2gFGvK
uI5sma4335D3i3E+KfvxZRdnaifJZFsSL+TOLq88Tr+5zgbvuMdJ3tRmpS7GasoS
m18kKyoFqKGhzfbr7iPESMHKwyfxvcHJxJtm2rrcgAzCb9eGaqbmdl9K6YCJAo4l
7286DHV0Qhdwz4MZnvA5id6174No+RCKteGAflr7NMGWZbe4tQpJum7ZYC0QpiwV
CREseCYx+WhXevGl41XShb3ZF5mhEicUh0BarZrlc1Kn2h+r5KpmsdMppZ1ys7gt
26QFj/JLsSKaPsNBhFa7LsHLhtn/vlFTUht4FBE/2Z6oydCW3mvLC632n/zjXqFE
C6l4HOzliiuC5moC0S9xF8umQS8sHg1ldA1dED+p5z2LbVYfZErJ5sD8kyZW2PeM
d9GVzHz8X6mXZWwAOHecwHEmbWvnRXbZjLCIIoIRtf1bY0/m4HxWFwbSRTb/pEn5
u0qGKxpJ9m+ebr4jEtJS+C/z+9o2QPUqJetRArO88gKDIMoVoc42S/zLX3JtHeIe
NhO0vExCVpNnrlFMU/3VQ40jSRArEpMJehQYQ5C+2nnqDtBc7SZKoWrHy7b2A86r
UkRu3BPakh20DpRNgOng4MrS4BHkO2cVsUx1oRXKzJ9vT0OJTB6b05TGU5vdSfsB
9ZePbc6iHRucm8FcRM35K1l1POD3llAbod6OofIoXu6LwKMDZHhFfSdeHck6vDA4
ss716bukltAnQYnxJQUke2rMp6ZOaoCL9SS/oJmAnI9lr1R8NDm2J5WzB4HBa9J+
jeP5lFc6+/54AC1U175wi8NuUMP5YmkkzV+jySx1969iWCV0mJfcYn0fR6BTKeiW
XZ8EArfGeO12vO8msTLhaUxB2aAjg/wbqRtiMN42JWhXisftor66jl4rEiDxoBkR
cdpBZ1FeFCLnIO88WZHWXSWad8WhlBel3gFDTue52rNneY+ylPKMg7HH8WdUtcjp
57tj60eSKL93MBBVRH9GL9l5+9LtOXwQeDtfsU26ct7pIDZZbvMcq7cURZa/2Sfp
g8PuYDxEHOuA0V36AMMEl/Jq6DSj+OpxXdi/61XaKnaMOrxndcYPM6oV5YQ5XG/o
i2OrzTud2eJhqhcRsXJA/LTtsQCFQYLCoR6b0W3+bb7wrCW4AuK9sp3ysHMUwxjA
zDtaf7QHsB6W5w4Z7BVSF7RS5vN4cGBmOVoSUpbNP1H3L2FS0QduQvHqtHQXhM51
SQKRel1UwpqF9tRTljxYvbrqMzpKUJX/3btP2AF2jIWGr7OISA46w1/6nT5Z1FO9
XH/kCxsySEjaCivp2gNDaoAacm5ul6MRcsR2sQCuWccJ0qxCIhnr1NNriAPpURb2
wucI/aKGYZiBBRoWrznNfL6iHx/wMz8CM57mPOuNbevFpaNjks3iGHNXfAokcMrx
Hsk6FF1YJt5HQ3lYafSJDyxND3E+NyU3Q0FmpoLMXfbEUIAMTLxqoIco3Ao+kfAO
Ar4YOhRS3C6R9iWVzAZZoJ8Ob3olytpPyGcZBGFGVCBwKQPBCv8ZQ0C5kmObwvcj
Rl9t51+uT9BYsvdqxhW5kklgK8bLWdPR21n2fBIT0Fogrz7biJr3eyMJjLSMVovJ
g2JRmtFhsbs8EYQSH5KlVnL12eBcHpwS+/q5ZRyhrRY8du0ZfDe6phqbSJVEnD7q
Enksj0R5diIzyTatCRgr6R0vUKMineoid5C5y+aa1Fuwxj1xznQGWD5vC6LdI3dP
/b/UEgo4U6HuwWFRnzbX3qhNpy2XoqOsP36LOLo2Fl0oNihIoFyLYCWUF+8wrDRj
mvqxvj5QxwsJWGxfQE3iTJRwYHEAvMe3MFEsfmaskscLmlnYLWf4N6h7esPvccj1
9BEVeADe26STczqwjWZpeI4gSCsVQ7me3WN//nG//TC3WmWVfOuxMkmczL58Pon2
dOGMBQ5DUjlL+atuz0OsTTsVQUbCyJM6IogFrwYyHQH7oViYZah1/ctKi4SbBohx
ahC2Btq8prqW9ri0bhbBgvRbMrSZAB8ytzjKVXMNqAhqElfN+twzSw4/BIQJbpt2
B613wYoBOxlKuvyM1zUbQIWPr4L9zb85pgzrsWwn0Ca/oBc3k8yEn50S0IY5TytN
qEvZiytto7aLd4fY5kfwYoZCQEHgDxVCEQG0JNvcc6D5dHL1+7twXuWFzDW0ic1j
fZOyAh1St3ATPrQfshMElE6GxV018NOrnKAnRnv+PP02tl7h0LMzx6u9fx0hOYOJ
Eq7meV/d2jOE7t6U5DMqn8vriVuJrrV6ooUx3f/CCgg/ajjQS469YvoDoHkbG9ZK
sD/vpTGhhpNpH17CsRLFeMQYmytNZmzPwMu04A5NvXUjtspjXYX8NDFQOuwItnLT
tWxE1KCeQkiaMT4BKvIRnNVHEjWBysok76vxdlRiKDHEbe63ZCIZtNG+z1bek4Bn
r+F51d9gtipulhqus3m48LK9v9GcCzzf3RgPbN87yYK1UruZ/UeNVcS0wqkl8Xb4
HQmiaDqBkEX0t0cn/iKxdKTuP0fiG2mSiRnPI3YzRgtpDNMM2nYEsSZPLL3CkiGM
cF1GiOXNZEe6byGr9tKUf5B6S3O8+GWi6srgwgWpYVn37+9L+wH+vBXjuxCbN+pp
/q3FVSBxzNkTvZ16d0E0K3AA3IZaYPvgxILbyp3ghtUu354l9T3VxFyJCuPhxLx/
Wt6JE04jMOeqbM7eJ6bMh1GwtUCVaXhdud0S3QfnXZzp3CQHsVebTILpMaakp//E
0AEmzbtohAy4jmjrQIqnLq0Mv0bDpq794dPXZ1wxtWOahtosJ4qoASmeGKNBT4Jr
ojaMSQ6oQuyGtc5PZwBkzzmVeYjbJzgFjwOr7hN7yVxdL+mNt2wx65/yXRnXqR8k
GHBGqxHhZu1m9TU5i/X762A6iTqOyLtbn4ZIioQY2aVYiKNnyiAwMfQW3Ph21mTU
0dIi+MiHB3WSDsHgLfk0lzxLtuMn/M7zj0o9qWZDSL4BB3lQD8pYEPaXc/K/R9KI
fpQlj7B4pRgCJQ4QAjg85t0zF2tcPItOtsPtYYNdxU70s5f5IrMBYAbPLPBwvneh
jKNmKAEWjkp5hVQ3jfDpOhxD2Pg3zFpPCqeWDUCabK4B6IJzowC7lGLCH/JuJ0eL
eTmPgz+8rExzoox/4VK8/xxGid29fIdgoPIrybHPURYK8jFJCs3p9lnDCtAeTkrn
vjDrJe3iAeNnGX4vbATRAJI3+jK2YZSPPgMC8teQ4OlcihkUZhpMJnhPSFnq1RMW
dTScVnr3WsYd4YWlCzz+1FwnqOvoTO51rfaiXeuMuv4UmVF4NIi+qfSVD9jFlabX
uoWmoA0rH2f26KKBh4pjjUcdhFvYxMaFUK0FGO2M3sO0WNAT1BCc70dqD7Uh2TMS
/SuAJ93gZG1EBKiyDtivBuhBMjd9JvDDVezwSXnzKCIf3bV9gGta1vl//oBNWrdF
yhlrn94CJDdyMnW0BN/8dgjEotXQ2kUhNShrVCr1ZUA3kKDNttQ5vsdZdv0bbO+v
uPBh6LTY9raLJ/tOSn8o6l+6eUg2BD7HSWOKkYH0ajm5cizUlEiilp8e2WtdP43d
lAeVKM/qYwNuAeBz+WL0m/Vyz5KxpEFqTvSVr+pgyHwAsdl1vbSrTe019XzxNEtI
YmB/LPFlbug3YuY/VrFehOGjug06wuozVouTL2JGeTVJaKG8X9v3sRZDVkOKTj0I
xL7OeEGLN3tfqifgV5GrdmNEBbbrY7TATh5SZrvh8rruwCNbddOLwR9mgKxbbetz
84r9H225FH8LlveNFImkVrWVPPu9kohoxYzjQsiYgjfrWhyjjnbXnBZDKq/Q+5YP
qmtu3+3zlcX60eIXXtYdfEAVKIoaOYaH/RYXTcYImNbcfF+gQ8mX+LPvT3TsPksQ
4GlKAgm9mE2qkE1Qvqdx7MN/A0KSKBb5AhQ4tg8nEH0cuH8o5joBEuOHPWBb9XPd
OQEBMmqfABgGVoXGSfs1s3/YZGEmxIkHSjUoLnYkUd0gmpuj80J9maVlJmKuCsFA
unpGaou5YKuX0znBp0taL0j/jrB6KlYk3WOCUoJKxWK1m4+BVh2b4J5Ukx0LGjdd
VWi/D6Kjpehy3q8XuC1hQceS/gMAMslBmRFVJCBdKvBzQ1Vca3FiQGmkVs1J/8la
m8ScyL6VBiwleRb4s/StrX7O5iYyPe0nFIfJ7MECzExndemJqSdt2arbw1AKAel1
Db3qGUvI0P3Qhbr3uQiiiVc3jE7FkjVq5OThF0YbxpvWBCllAcsLnWy343T0TGpX
hlzxwDDudSl5Cu34GYLbExBq4KD6JQVlnItCTjt6PNLjQjW1v/J6ay01xYy4Hsv3
VDd12ffTSC0Csyny1xEY+XOHl/Bmkc74B7VSk2gNhLzxBfAgffbwVZqT6/quyp59
be08RefGVcMG7gpEOZo9R5KuOJ2h1AEH/BPCAmAJYR8PpvaXE2jRf//LpmycCO1V
S9hbysZ4Vl9MTwFwNRpU4h/P9LlE8brVdHbySce/97N+oquXZCc3qd1menVKuEp3
7BClh/Q/x6kZ/OIBxhuMh/9t0jJ3sWXHOoUOZrdw2oQHLCW1oDuzBVlDHo6ALstf
S2MJVbOeLCsT8pSEUo+zDsvDbGxvTqeGK4AWE263L9+W96ZE74BrtrMH2RpEpdl8
VCN/GlTin32A5dODIQGuJzeaBU/oOB1YQXK4cSwgYOX9g9dNCGJjFZHxFump5btx
VdnDRbQ0LxolKE9AeDuCCbLO4bAi5oEcIfaV2EtBdApjP9YYMOqpq/VPNa6VbSQF
0Hnr5j+m7oSzEDEXoTD/HYB0cFkAaE2XE+67JCEdimQSCEn05gzU/9pYiBFDGvzf
nBc2EwORt0dA7xMYnLxiLrKVlty//nKrve5yOKzI93tlkNasBvmVrOYSmzFNJuma
hlPbyUX850WIOj56o2WnJW1DgaR0cITIhQr07TKq9LzO9fRaaQY4h8xiiM5qAHAu
804ezkQLABv/EBzbMTJYU0mu6DtKZwKUz9xRIMdvH3nXfoncfmsEyDXc+RCuPHD0
Oood9uwrWsNco5jttDGnCUqGHRKeJq9c3m1qVZoskXp3TlRCf0dPoBU/LhELBDqS
0LvbYXjFXbleRgVmaYUlQRyasPUaMQQduRftgbMONxrUnuEg2Y2hAie4Vr+DkR8l
x6NyxtSnPsvV54p22xc5jUwKKNTuDn1JJ2pxL0JTQpMucc4XCFMkLcvGrx3BLWgM
VZ+1qz98ZYUHc2Z+jodKuoGebWT/mtzqsbzdiDnSIFBnSYpBrTX2udDP+eUPJfU5
Yd11GrpDLVxBnwcwenwvonO8K/yqRy9YljynvB/5Ju95NoS519lvGBv8nEqzNgRU
lV420sPTlPjzNmIsRZbkPCD3We7zWNjCYNo3rDjqFDIfnc5/k8QZF/2gqv8qJGwG
CQy7/fRiGrrxEJD6SHZ9kUT5Qd1eyjajyhg4EL7o0ObvrzpWezaJmvJNDEKXWyBi
TOKWOJmpAqDF5Wq2tH+065wBIh1ltiA/7VYW0qolW9cVQnd1WLsuA3UuChs5yP3U
AAumwaAI651nra0q/Ldd0o1xPeu6kr47QHcGiWBstjvvVmPxu2P64JpeYCXlff1C
vdea35+ISW2vmgGoyL09Z6r6tvPaJsvH6+5xCWLU60zeMGARxV5Q7e8qTgdrBERP
rJbNKbsSel/CSyDz5rHNjRH/u2q8J06jcFuJI2WQYykHA5MlS+x4LeW3876fFrxr
soiL+DMxB1AodKKtV7EmZ/rHPQnlGra5/tO/ILqO+3Q8L8fmMI+k9x+TPMyeL78q
eU3b11zg6E4XJISTfVdvqcktxNvc7CYUix2aM4TdcrlkEXxmJLC4LgPILYsNiF1l
rb1YDWaPsMDpDEO6EA3H0IzzdMjmGzo3qVnfN1npqV823q/BTtzWqLKBypEFZnwH
nXtbWrUT0iIWqq/b5fqWKEZAfdpAvKSkjK4x+SJikYtQO7fyQSodQ2+SV3OaofjF
kH0urBJXfBk1DqC094wH34Y2QcWChsIOAzWsesEEm/vxOEzT/iE0J/mJVS9Pt/Vd
TZ9sZbBSfuB2JG/J3W9znJRqD3mfWtw5j5oCgSLGm/zmb5ZgJzzUNsBWm8RtsqgM
a2oBpOwe6DwkzTKZgnk1DDEAaIIkIvEvtKcUZ9Xr22FVUhboamIx1kVOz+tZtI4B
1GAP6gBkmA/nyplhnuZ/g2hfqxMCOGK/UOysAefWr9Ok95r2bUoyYerxaH+KF0Pa
13H9zOye0A9m7Pu+gHu9zJf+2DUh0SkfnQR45i8594BfrD1TkMNSW92KVdsx5gCF
8v7k6tLUXviOonkfPbR2Xbc1pVNh+KlCahAfUmNFFa1j1grZV2at35054WcYCR8U
AE6Z+jwyCFSzo7Qa2iMZZZHvKcBKyMWUvkFY5BRd1oUAAItjGBnoZkJdRJZOc2DH
3AUYUwX3Q3+EG6f1Bi6N7PH4Q6Syd620HhdtMkY0CL/SHul3HYkX0BhMub9GC5O8
8Jy9208Eg5BA110I3te+52TkY4KATalMwFhQwN8WSKouYhtxxYPTUVKPY2yGESVe
BveGdrsg3h2q1iYmTI1tgg319LRFiqFIhkNqTxWD/71sEnVqUK3T61I0F3BgUY5E
igjzr7KUT3HNlosj+Wrv6+nHOe8ve7TVbe1XrnUELBNl/Pq3jaPiZZ+M4coNOpsF
wtaIqFgJGLU4LLltPI6NtqiEDPEz3j8wdDDs563jnloij8CCG65ef5HtIFKJixcp
sx6tG3nxzRDjbNigj3ushGPpqsygr+XeMGKPsvMJ9Nbo/qXGKzVrzooEddE82agh
1J5XD+X04NA2G0mNp1ciWg6RaARr4GQhAoNmu7Frj0PNDZwg7a0BHtF2SV2G9h6p
5k5cQuB10OQ3GL+1EcpoX2czNnzaS8J98erdAyend8atZKR9NGgK5a19Ss8HDAT2
Mjrd/GLirGJ9tSa7wzSB2FSMwhR6522pCEvdvVoUbooDRaEwJrPaD+lfc1aVChJu
Gdk3OOKk5J0v04FS5NToqSD77cdZ7YYlm381m/6CcbIBcdah4xcKYy8M4DRMHOtW
VQVRVkEB9z7lv2BW8xm2wcl0qdPPY5x+Tn4bYjEeCTLzgpmHw+b0tkRliRrGUYVh
YfFXqXdtmD5ASevyqY0s35FbY3H7wEbY8iayc/NZFsjFabLbYlwV7UY+UVg+TdsW
hTJNc+DMllGVEJ8IlAMItMkfFDM88Q1LdESxKDstU+W7jWxGACFE1PcDMA2vAEpG
v3RrPjJxN/DsYgcoM+Ce73yr5k5iB/AQxboV0R9TD6MQ2kaU67NSGzRAnaikUob8
6A3j+yzlH39pCCr4sdDJg8/tU4/8S80hQm4OtyHMA4wYH1LFG0ymxRtF2c5fhVQH
VOmnq6wi+Jd6S1VbZ4bHLMcWj9qfZbKx2AahzsL8WUfhQkfoAcon5Wh2aKHnOPvw
VuZeS/JBf/+qu5XW6L/QGbjJDYmHZdzE/u4TPukUwEG0+8LbslxIZQ3ucQCraspk
qI0UzqUVqh0samWxrdy395iDLUXL42TNqjHJKV+SumFECDqtqHeVSjc6iZQsosBX
PZFs/EXZvqo78cOiIa+n1mvhfNscFH5tsQPU3c305hXR6LqtZXXt/L9ZLWxpC5OS
tn3ML9/bEFKBsDtEt5znJkDzCr3/NOX4qrusEoQII0zloaNL9XapbQvx7Zp8RqqH
FxP45zjzokm3xVP4yt4DIkDUEOh9LDVL1PEZL6172LTaWxs6j+25co6Q7SytaMNC
H6sFb8cJOH9oqaNWpSG6MDRCf6/0rnn3OJUHbuQBAePGqB9oNLsZqyNJeMfDzxqG
gWhC25/BFBl7soktAbl4wT1CvX7Z98yEFeLob0sefQYG7QM8U+Kp1zkxN2XIdG6+
xQYgQsGLB2GJzScNnHEV9wjBGGIodZlL5KE45Kzv/HqqFT6nI7pTAUNSi4hjc+hV
YwIJyrtgU/nnN8kSXMUAk6Gl/DSxsqhGT8dokgFqrgt1XE5MVvGMYqo3yy26lRH/
xNIZz4XAsE2KvIJnwb3mgBxtl/p5A0q9CEEDDam9eBnLH5T3dIXJePLX4zn/eqqS
yRDZ5d5YHMsngJ3y02Ry0PzlPyxaJu+N0ZR6FYABfrF09Yaa4V1v3cWw4wFqVl6F
6yqiSUda1ejHPyYt+DwbTnYpbOgcC9VX1Kin87cXG7jNoWnpb+cyvCtziOM0Romh
Piad/Fr+VgjvJDCV3Xhq1Smm0rvGuOgcaCxs9kNf3FydNYncP0tI+T+IRGUWnCti
dAxf/QjCgSkPvEjAZnd0OsUaxIcLJJpUa4Vay1WUd7Xmlz1J7BtX76oQcMiYMWE0
2cQk/cUfiuXbpqoe7BSO4cDe96UmoGUw13uAgTERfFYgAvgdKJRui5Y2Ugl0RH61
w4xRoKIOZyD+qTEKWgKRGeiCwkHF5dX2eci+HU2jgC+qrwA/Gco85mFddRfpeMh9
Q3x5ZeBf2zuZAEiP8cp/H71AjdHywwKy5A4QhxRJ4uFCu01+3qdhVmufTxThLkjP
8IZHG01vrc0KKVldO9VbJ7u58Q4x7ZVVePaBQoPQQGXxNCsno0lkfdrmUlx3dnCR
AuqYzHm8LJyqJhh7gp8kIg4T95DFjwEWChLPJwtj38/Oy6iCs66gvy2Qgp3me6C4
v+KHYsOjNgYMRv1NK2KrIg+p4pZvJ8pv7/6+pk5BpU2+a6M6XPubdRtVNYSt2wir
eTDGX61FV3aaR73HmKBSaSuizMCw6QSTSstZ11UX/UXvWlkDsn/MeyXQfz3Dxgx9
vMtz0fZRFcqW4WINBVArzZV2ZlYDmp7c2G3tNpJmP1GhaPrPL8ZogoOQy5L3KCLc
jwCj9gQDGLaEAxd6SMvrmYHSUWxbmhM1VQIdhh2hJ8FMjdMWrnp04A2n6AQbl5aq
Lmpg5HBUB8YtZtZAQLQQSOCnypwkqcMKHgv1GJwZhu2yZSkCtDqno3yoXPZZgCPi
jw99VHZqG1MlMRd5LLyVk3nNP1PYIB4LmfVLCQadPK7mmHQE7Iwpi6BaeV2XWb5C
uuuQkopLB/lPh8CXlxqRD9kO94rBGkaTr9JoPvfVNe0vJCAbQNXAX+Bc2YMvZPMh
VLlwbcipdyOks0dw3XRhOS0s9k2sGG8KWrP5GtGJybw6nhcQ9AuZn3VRZ4VaPubw
8TJgqF69JaAPS1Ayb3AMz5IqNGX7QwGKodku66kYjpcL0EEIThQOvqfB1NZrwwK9
CjN9eQQ6goye8gs6TDvGCnSqr2qANp9N7Xy303HcNDfiMsK3j0hx3rp6pVNNpld9
xpjj2JfwZUV3lYjGL/r3/TgxZcCbaPhk7WlVTEpBsUc7+obwYtPoKuBrj46QOnFt
b/uziovRJpAdghvfx73wnCJ71zGXI6cLjjcLAlBcu3xLwFfmjpPCw9VlQcZ9OxfA
sQ8m1IyUX7IaAMTsgkelM+ucCHEzRpg1NYAWKanKbGXMkO3UKY/OH7oYTSap3p6D
ZOYc121ZVcS6K6O+UON8AvZEBT5piVJulAEXrAbIAUnJqX1enQON51w4YQiALzLL
V0YAa3s2bENRaNU2SltQoOrCk+uFHbnQh/liCGOD8DHv7MXfYUJCvYjNVctzRiSd
1o69BBoxLpG3ofDTu216wnPYG5BKDYp6fLUVOlsHaryILKQgHwNEsscRnOTcgXzF
S74IyPEoz1Dc+UgK34uMTJLFxo8+nL4mUfofDLFPqblfx214UvNZGbnF9UTzLgr+
DbaMD6wOzv3QoQNVHjhNh5PN+UwBTvEzx5Gwgahg2+URaOZYIMn6W/0D4x2M+HsB
Q5f6o1HkoXAb6b6vnn2nkktem2LK6xoH4/qFiy4f88sHG1i7uhbidCI6rprnDrFf
8H3p/ovh2QnorgDQO3uJl7j8lxhhIyK5yfPoKw0WrSoOeMNL0b6p0BrVqZ8G3V4j
eIjk0rwV0I0/DjDoo/y0jPVlufzteaQvVciUrCj5XIGbanrqMeNICj2rrXIq2PpH
Rls3E360GQUhPmtslpATdrkll7dH53cn5uU5yK6tnsrMcRXDkjX7l7EaNz8GP9DN
e+969q5FfwL43ozjviHnICNH1JENdHPpBzAZrqCBFzi86scITylPcx8fho529HZx
Q0u+LFjOy7q5e1PcF0P2FzaQUSfHQ5CGKa62PW9CVjdPkMOOyz8RDsjzyaMU6Y00
/k3mPD4RsUSL3qYu1xCVpb9sw+328WdEdeC8zPOCkO030SUKea3OrUckPA0/6vkb
+HeVANyX1hKLts6ZK+KfG3IlAgFbIp33eYQ8EYhwIZIlg40xfTYlqTCbwytw6nkS
9HzP3nqxH/NBQZZeKMyi5CaHhk04kcDxmK7RdeOs2dvbfwZeMtuD7ozKb62Qkf8/
3e/Xupx0YGOYLcED3/JHMUawH7a0JdQ2KSrL3aTuWdlS5w9yYEavLIpubZj+p0j7
fVFlqb7sqgttZ7VjSQAxNXWywMbX8dTByLUrgZYdTmAzaCAk8PiJPN9dB7T6BVcO
Ptw2ADDj5WPUFwI9edsnTmCw7b9VUwbq5uExSkYnHWHP6EnPtKZ2NLvMX98Y7fgL
ijpkX5Rh2h6uGAPnUOejlPhcEByEvvJ6pSKP0+oUviQM3f4nYRRbnev6TimTT7Re
cvTtb761HpnBHcuXVCh4ef9oc8o9O+lEHNkiVBvTtxMrWRl0C+Qg1XlY/HAWdA0h
AXmlO4Zsb9+vxTGcxTANOfzcdwTccRSQ89xXsY5KHeNLx/lbpohaWaJRHbgaRqv1
6lqwwVD+gU8p5IMpPffY77qP+G7U3rGy2InV/9BsiwyGRuqpq72FQJnmrRA31ZSb
vel0zAWzGmRsi/9vD7/UZSd86UMXfEKbaPATrQia/na37LW0PCKdjbZcv7rYiJ2a
5BceI5D5AX/FgwmcNhz6/U9Gglqsm+sG0Elhoyw6WLIB3EAgKPQE6BOdJrtXdDEs
ReqOtHF/yyWyLshDhc7Cg6J9WmBkTFMpz3hwno5Bc3Dy3hMJJcvT3HktrJXFo0HO
erhGiqmfaaRmw40e+F9BASjfoskDTMLRn4RA36XWMyMoAc4OJ6fFsgmqhDrsiMsl
gVJR1yc9nKwiO1RVeL1ojbD1HlB7tQsNI2yHo22F86K04KfIWSDz+hlN3kgiMx0C
opEDsLQhtiWj+VvL2H4+aElx6Cs7TWmbH7nZimuQUCMMnvB9zWfMt7wAzMviuLWY
+yiWrhQUVXVjy26iIUqudZSWEaOgn/rSLotzI9yirvGAjhK0U/uf9ZQthqpAQvU9
BClP53VbKPfDtQ1uACoQpPUxogNvlyx7BftuZI6QhWA/xdV4UIdw7iEeopq7mG6S
DpDxKhi4y1gdjHeODwa5A4Fx1xxRpT8edMKBHXQ8P6Fwc999vC0QlAYWMR5zl/eF
bfVP/N0N1etvl27w15hxYBhfc2OdybcOW9HMnV0rNUQxvFbyv08POfy3yp7YClfp
6ZmeXTDYsG+KlgQDbxIHE+gxSlyfBb4SDxEiuT0XNjPrc5nOO+to2+H0StUKEJlK
pSSLli1BZi30hpsfQ3ngM0JVhht8LprrUUWhUmh4FdjOkO8NqGG4kP7aK4SieQug
EBM1vo+wlFpOcM9TEU57xGLFrKXwathxKfE/MiVLF0a8L/XiAG3+RTA9t6ggGD2V
Qiz6DoqA8oFVNeQcMaOCa08cmGiagfJ1djdP1dt6sbIhqQ7Z//Ug7V2WVirO8a16
5irU+VNJzsS2E5w23hexJk7dGLMm3wkcmE8WXeD36+9a1Jls2/KYTTEaJQ2+5L55
FJ/7bbndxER3mRqlfP76m+boDsDNRgo7rZPagRioga5a2fQhgR4TjWxWW7KZTgQg
CmPFx8YRzW81acl+5cmQkTBxSEoPvF7pA1HJF/VF9nLP7aWXXnZR6uUK9ww/YVvy
csjRRuvSN1XPhNTl5J/Q81CQ9gjg5bYtjre36i/zj/+UAr/O5aUokibyjiLvLztc
88ytVosvbXJMhQOTugWpECX9lJVUsXXJp0QoKjy7q+18LZm+DHfIBtFJeOSQfI61
GI1b60SCFULmyH2NrBNzEZYcNgw0ngNCXth7knwSHVKENc6WpGHusY0tNZP8Mrwo
/EKPdKpXqOwpI7HiXHNH5uzpi45cYi/y+MwYGKPQ4P4FX3eOtIJ7+fGP9qkwYYGe
TCho0rOV0hWu4h8YIYxSrlwYweVA+i7MJT1ZoWkuS6Ibn9AnDXpdlrMy+u+ga84P
o4VaGOXdkrw9im3Nn4lcJbAyzjNATh3jmv/UXWcncNbLsIF58pAdShXZoJP5ZUEi
I2+aCzsmlzlSizjMuZpI/DAOD8cV/PcUM4NUCJMkFQ0usj1mvWys+nvvesKova1v
4DmWPNFIpP12ziWC1i7+ZvJfWrG294h1rCpHwXFsU2u9cnk9Y/dk4bSLBsUHStQr
WrRc7+QWlqIEE+xLCxkrwq9K0CqRj2FFMOc5rkie45wooqsqmUIElweoHG6vri+A
ADOfia6NEl4vJJLWxj02EAAGLyCwhZbf2h5glSXN1WIFwmWwbjFil6wHPZpywlw0
N0sVC1hrKD1zFtGgqQJGQJPmCRxJKV6GvxaZ1VZQmdqr87MGamC88XGMposGZKtg
ERHeVlMJ7ukJu+DiiT9h261b+ARLPQXXueGNHtpWM40zfX+k/6UU73uLkdVYPXfX
N6pfExOrWr2+ZsXXNxZif4KIscBaKjxCOjzFOjM1Um9JrfwzrU/oF03bL+ylwwRR
9ZJpY7Am+yQCNLie+eqstvVZmXwMkyJSjnRBB2EOGgEWnarJq+Bqu1WawLSjXx8o
C4sCvHVEl3442iROiY7SOOsj+iQ9HGak2dcmRHJrDKPcuO6kGFQtKEW/GwYjXdxL
zXrf5TzVI3HqYVy3Lw9gkMyro55olzDXNTFyje46Ii1gK8SSuTK9IqoYalbK2EjZ
zpGqVUeGCDbD+0CqKlBUbn62EoRXZL+dSg/K98u+rAACfNZ1l2h3Iegdpd/VVuK3
lrqx2q33OWJurzscIrwmy8IWmsXhkccFQ5edKkuIH2SgGINbN8czdutmArS1xK2P
ObZ+Rvs2vXKIaC8jcmfsoU8xL3z4kQw8aVPLPIfTK2Kk+Sovw7G3wvPDXrWkvV3+
Bf+iuNx7i2Aesa3PYaMbIhePFJMgE6IErAroyEGw5hQE/HQY/F1XRqY1HRdHeYSb
Rmlz24ctkUzD6nY6ExwjEFnSFi2E/Rz4UpYkUVdLzj/33JJwkAJTJme+0+WRwM9t
6cEHMHC4tasRCroZCWXvznfk3n45lFqG1bd6TCK3CfIVauQX3tLftc9aKhvr6Zh9
cG/xoTTUr4fl6y3g90IsSYQsodv9Q74Aii2CdeGiq5DQz5mm1naMtUp0B8Md/BPS
XJd8oBwFJR5r4KliYYz/HLkainMDiQ/J9PgrX7atZ8n4znQKFaP12f9Kmygq7/VV
E8JSudtMXu85kt8SsFvzEnOm5Looe7PKirLHWqbcA4IGQ1qObtBfJKZ6hcuDNhmy
aeHRR2b8Z8NV50zgsSi1YdJq3XwKz9YqzkkrCvctT2h7vIi9IO+NiX8lAj0nFHnN
GI7YluG9TMuMzMXdgMf0T6axe7ybDspuUFJRx3p8wAVMRC4eN7fJBI/IUrziVDHB
CFgJC/JGhQRwjrn+PHDE8DKEIXH+eq6T0xtcUsTDrSWytk4nGSR2Z/jZElBaEwO8
cu0b4F7bU4bXu+WAYygdSqDwUOJUsxQymgB3AORU1558Gie4U3vimdjo7/DOyjCY
UhwFyLnJYr5Oekagcjzz/R+4AkP04km/BHTPKZBKfqeQPAuatJaTJ7ob0eHlIpAv
igZvet3BtmDvd8hti8DNLkr9dxCDJhTWsdtTxR6buN9+sss0+6hK7yZcjBZRJd9H
GH6couc4WRAZUeMJt3fTSsL5QhwRialD1yZFjYjmfV3HfkXMC+XVQpsOWHmvpiQx
YUeZNjloXfxGk9qROldwb5aWX4afGQq053/ZqyrX9nGADO13YscEYfxatkpBx6aa
h4x01uTglNmR46XWA7CQKRlSJOpnmTBoVCb9Bu+auzedSCSMz3NG6Yf9Ll/6kAAb
RssMue6f1kqLVU82Fk2I+bPPgNpPsvhWxNfrssHRpZvnzez4XKOURZVQIxVGHWq7
ByfetqCmNFqEgLIdkJcs/8ieDdqKFzkGHD7Ir2YKMd82E/UJw+jJffQhdjqe6XiI
fZa0UVaTGTAG/mEGtiS5FScouJ5d+jVOg3mTq7LWsvP0eLu+r8cZ+bdZDHqz+NPN
Fn1tG/HyyZxv3JTO+HJFK+VMV5Y9G8wrNGvof9ZiR8TM98JriwEB+q4CJu5moUk8
qgDdXmYei1j7vJVMU/XNWB85yCuw5+E/7P0FiqWj8oKmesAT/UGMyULO/FP1tZrI
2h78ocxJf7Av4rY8mewqT+giMEP5e7wan4aOPYlZo78fHMU/FE7+VUGr6BkPsGoc
5Pyxptfn4VEr/53MUqmvYA/knoYK3KdN+Hg4Gcnqdm/OnSaYMSrcq4OzSaFkm3DW
i+Cdx6m+k2ee8IumY/VceFJKBED00sNibutzFelKojCnwgm1iguT51zPFXIVyxmM
JyySNfhzobhHBcxGBFnQFOqHDWRee70sIRz09z4qgB1kE5qtOQf36WXTtYgq9ueR
r8TAlap9k0vhaNy+tYNE0Pjro2FdPwwiUr/0DzCten7fGwlQehAHrvJTj6eZoFFO
8x0MBymdr468pmZVATC+uPM2ctkbq6Bg8cFCEiesDgwn2Dwt8FFzvdFUK2JnCgLf
l+OolC8sKAhuODwxqMLlF0i0QwrwSgk8ZWWUj6GkLcrnkdpn8q4qzfHVKeF1K02N
3KYPqug3EJSwSlrf2EovNCBAP6NW5AhdWBOaWtBqU2JwsN3iilukPhhHuFBRV5of
QmgbzyAbEJZrvNYob9FZkkbWvh/3o8P89KtpFAT9XU/Bz8E0Wp9qRXqngs7TvOOk
jjGccAQajFDYXaZ0WwfZ6pDb/18apJVa/651sDbEmFaUYlfBcg02kq4TsNYXnnJn
zMO+WN5KRugp0w1lfxpYNGfSjps9H8QtiRlAEFXG1kDmMP83pp8tIoElxGuid7H4
XteEluibthgdRvBFSaHs/O7zZchNHt3mWoPt5wQHAci4dXy4wX4si7Ny7UVgLOZ/
kOk5rwckj3QA8FxH9kzG3jHKJq4H2jkickazu/xImTdC3tl6oUqeZZP2aNHx+aHv
sHT/kyF78fEJLfR0M51LUWytiDrlp12XGwjsV2loDA0PsLljtaAd7Udr72Cqr+s8
8oWo1nwaR6SBjzGqmrqWnLwY8fLSmaX6OuO782aSnPFKm6R1ZWQkQt2MLEusb/KC
FuhQmPAG/7fQQLcenL0W3VbbqDcVPmP289neNBRAlceU2KFTqostdcmdf+QlarAf
0J6fXmlwNbg7ak/KYRH0aP4uxrqePW02YcpWKN7lJJVW9q484zG7O9VlEXZDOASM
koF/zav0Ftu0JChOFD35lKmwAq45JS78Zg4aXqQYMEHPBrGDv9POqCO745NmZXXw
ZV2JRTJDMdiEPUfvM4xuE+CLTrxz7Z4nkB7Da8hAtDireOcBcPwHRbjU8xtfkQxF
Lp8fOBMubhX2wSWbAMmGq54BUyP5HLkcTBEYDqDqPUDvDhrunhZjRjfjuzKpNevj
c+X4irz0bw2VUaM91TzRmGBcyNtgXLU7NdPfGlIKjoIVas5bEOUMcVYbLvxkCV24
tCJu3hdPWh1tS8+sFZHyPaqRWGm3McpM9XpvH5gvD/pSSQ8NdAJzd6u51kNyY6KV
oLT3/qj1WOq0pJuustHm8UvenXZPe+356g65DNBlvPDzKHQbrQcQRhZyV9mmanuY
x0OuF7KoAnSHAhGqeWmMKpwKRxwkqvyaIYA3OGprW3QsTX+qaLJAbl2Bzd5byewS
I8XlXku+DQP81jFYtpMuZTnOjoRjzu3zJ0VpzyQvOBNBCeBlWO7PrYl3XbNrjUCp
avOEITIvrkrxUABXhb7da3mqpJD2bsHSL9mvoPbBHmpZ+3gnaZwiNx2Tp5YnNkHG
jnlBnWVmIZbag1hyRbHyOeWyWUA44eJjc+dUJMgTbEWBRBzbh2Pli4IRA+2MYsE6
ennenCCcPD3TlxflbxJisyxkHKIje5S645ifUj7cFYDQ0/IBi1P+n27SebDA8GXh
9FC7tzw2XHHkCiXU+5lvBf1vu/QcT/vz7wz2E1zpfjnSGXFnAzLL7dju6MvL++ZZ
fSmmCoMzl1tW0Yvat6zSxuK7bDzEJmz6W6+2O9fi22Gj91q75I1RN8JXzR3oN2mW
ZfoYXy4QD9aTn7SWj3gwuW8vvJKGhBWSmjuuHOTqrL99QE66raBnqH/6ud3l9Blc
sqR7xt3lUR1lcU/l2EbBYcKbNpcXJDDx8iOdBJzo8HlUIF5MbGbUIE1fAUfqh++d
CxrZAjsHMwARMlpv+7P5JzOXVPhFYz5f3Td87QY8HO0L++D3NKuU118Vucu+vgb6
dPyAERNaOGRDdbi+FHpjniB+Px72o0QguHhzr4LZGuqn3w79gtv+KXxlQpK0ICGO
quiSXkr2JayyA742rJ6QTDn3DMTfg/p7zBzC6fIg6nCuryVlAGM/o8hqYAD8on2G
HvmqiIQt1/8fqDrCSgEL2k2pE+YuZxaAf4lZrHQgipZDZbLblDkpFW0h6X+QVWuW
C8XLYTPGULYsVY3IA9MDX3f3RvYQh04XIUr8w/ZtyJxCNgQ4n3OneJSRcuZ2uHuz
/v9QTTzIHYSV0aMiVb0nKh5P2iXSZ6FKEUAFYAPk3UWnQRLOhNp/qllNN7kKawLa
hWpLFI6Pl2tSyf596wpRlGn+qj4pM1z3HrH5Y57GBns/6hg5HCcBg8KmHjC2CvxH
NS38bG6WSp1Xs/eLEXLuqmuCkWMDOQTW52BSIH/TAqhqW+RVTUTsT5udZIah5TV5
nw529KnqFVQjB7IcvcYaIiYXgEWqI7TA1zilyxl1lrkoEV6xG+CQ7D2UiW4YOFKn
IV41NSaEtpVCMvILFjREl7Uuj7+vHjXokaCRRyxQ7Nuvt3aVPmSAdyyMxRhND4nc
KUwH/w1LzVwZX5AYViZWHdJmOTvdQkUTNt4n1ltbcPAVbgYTDtE87a65tqYcRxAm
cfx/RZbzyFBRe09NEs7pc5aQUkyIMdBpUXeetemeW1dSLTPC0P8rHFni0gCbVItJ
GVgTxfrzXobhN1zXwQ2mRSu0NvObkeVCzBfku8jAh9yhOXTIb/u8u3gQiY7Eeqy+
05hovdVEp/4DufSGnHhV/smkzdVzmshE3Va8ZZeG4V9h8Bz1b4X3oYZd2yGxGMJj
nODnMKgTpMXbvurETD3BdBepaPZDmkBXp4sOKpaVSZTvOayjCDoWsArxkujAQ4IE
PHeNoP7QHVsTN+RT1tjBZDRvL0EMzeaeAaX+H0SGHeXRiiA4Qlgbr/tieSZcd3Z6
BTH0Jy2PBvUpmLdr2uVtjXIwIk/JnxmDmGiILWH3bbpPn/P4ebXwRpJ73egHuIoq
MGxJ2ba8nlT9A8FtCmfnoty70WadjvfGZsm4m3FAItfxt2zrYYDzMHHQ1HVyTm61
cZM485BerhtGbxQ5uN7OT2r2eH5eAlr6EgZPabIQp4HkbMmCy4Q9MlIDgMFtbb5h
eIHPpFeA0zkrPKtTFNwp78UJygiw8z5iCRwujoO8lGnSL4HJnyofk6vlZkUEdGMM
U8XA92t6yHu6gE4tQRjBc3j3YUjRE5XekSGiF8FtHBtt1mhdPpO2UHz/mZOsvRDO
gTrivRyfkGV/JyvB70kKpUwtkU28igRcYMakG2/z/TJXbF0fR/eLYpUu9mXImRy9
u8RVNd/Ao1bV3kvmXEVPXmzBvOfM8fcHUQbRK5hA0q3WgDGpQhKCvZKULtBJAxHn
VUAJEpWbudjN8qhXzmtTiIWkWba640Zimbve1zL1PKiBbVjjxaBmqDLGJwBR1mO4
rGzhC1uPQAE06pJf/A0IxXwKSUfqqSVSUVtnSuNCwK9D+qaI5b98lQGkGRQRZiOH
Cb5XCpOy2OdJNvHQoRDl9cdyVEu/og0yz+0u/4q6cEnlYC3o2j+yhlYRuZ0ev97B
x6ArH43Ixeny+2xx22dTeDsfBbeTB3aqqWoGNPp3qT0yPGfWoxxMJeFRYAeeqJxu
B7e/v6oWjKb0Qu3nHIUsCgEn2yIXXisfUfyh3xnIXeXSspFQPqrJR6CU9Uy6Mt/B
ETe8w4+bTcV9dqqQhLU0Vlk99za51l1hZTRbs187Mqz2hIn70Ntu3wT0PCYXLd5c
sIrchdasYORExJalTA+0s48rjpZ7vhGRS+cCjbDbeqxnCuuBjdJ9qTP1a+qvAGnH
eHgg9WuTajGrWRTrjmSx+gDEewpsDIdQX6VHKz9oJ+Z5aVO18HYKhkeSo8Uh5auD
vNC9tieRCncX80ymhS8Rgmmchw6xmsFQxN9loT+g8ZUEzsjyGxhw460xaslCa7eO
jS18LthdnTpD9/FuFbE3GzS4iGPpbmOACGMxB77Dtg2Ge2nEIzs6g4m23mk8750M
V9QTZUMitD5p96do2OGpd62o1RZKADWF/wPLnKep5nfBMHaQQVvYbMMAYWqalR50
XUfIIVtfX7V0GyuuwltwwFZPCctroz+PpsDOfFUwnP7qlr57nbjk07veB+vWEHJ7
BCTxKW0imzZZCoJay5Jp5/Vp/KiOTCZ7H0NCmg+UKhykL76H+wyC9HBmo6JJivqh
mGxd4JTJ6R22L+1JOMJaxQNGsjsHU9ujAwxtrsZwlN5Gu7Flmn6SHKrYfdYZXLQ0
PcypejTm2hEUXy1ONbrcLk9BdrN6tggmtIGDbtPCDZs+VcADAGCA2+pjhOEdLpab
7l5Je9fBcVCyarSI/wNkB2yHcPbBDIO5s6jlIi3729oLBHSjOXAkodJvaL1eYDxr
2XL5tvNGs0pvEkspfB9iZdMbJVCGs9TAV2Z6LPkPw91wxkEcE4bqAzdkgTTIrena
y7IQM9U/bu9zcYOE4GOV2IcR9imJHyws0i+/1XjjZubYvKjzEyZ57PW6C1tL+koU
saLulXJvz4jSeryvBBcah6A8dMI7M+UTYIKy/uyyenIxcLak9bPu/DZl8EXiXe45
TyUyTurhZMUmq8rO88mWz+gd1I9PY4dXI+1a/g/KvOVuV/CD0f7UuMhp1YDFQ7OU
pme1WqwF41w/FxhFoS1MWAK7mg+1H4Ke04B1b19fxQsXvA/+5E5aXhc8SE4Rni58
hvSswJdc+gYAR8Mim42Yq/xtGgOwmzkLIJrKfjferBlToMm02pW6DycqvqekJYqa
jk0GICgt5iHJAQZlwGOlAJSaUjeBoTBJHO8hqhN+/cfylS4iHst9O6ylE3bZeky1
Lfklo9rQcfjR8zGxiEVE+zlPcH8Z6E7h9fh2OtIqX5UwyC2bcUCmf1zGtEaO5FiT
AtZFagoIsNDYrPPeRi1tgSAmrTFc7uqaAkCUoAFaK/J7gMH9TArVKF7BXgEj3oKa
SiPgB094Z8BmyE1aHXuSTUYwiBqmsjKt77nhCFUYQNjajfxwOCUl0wtXuPB6L/Wr
ctEsdSSV4YXVRTvSgmeAie78aTN2lNa1pfVjyxCwSpip3cNYemcUxs0Pp0s99w9G
HN2PZPxfV1n984YuMWYBRN1uEEOlT53zcaH0UuNsodxN/hdxZ13OniA/26HcaGfl
EZShkjV8fuNitzqI1E2csCCkZ99C85K3fN8ZykwK5wByW3+0U1qXtX/O3fXzNmrV
YrDOCwr5RHBzbRtJtQJFODjMgIrUgED+LIeBlq3BsRVduGx2Fm2JFngm0pYWkv2U
1P2dDmneoHG2t/nZGGIsF/6NEUVZJFoM0Odq0Yoiv1lzur1wfCaJgiYEEpttHnTO
R2REbgz5xaoNXz3D4BxUSOcIhIXKo24CxUbZHu3I/RcXfWYqGpD3UTQLjDUuiupo
drXjcZ+BZQbNWs1/oVdvKd0ZDW2ohseeoqdbB781+lrpGHwmfJxNl7z9AlHkG3/s
jvnJF2i0fBqa93vBckCU0HaVt633unD6dzBCqsethpb03pJPWHSpHfk3z7YuaJVC
yo3ObX2r07uONx64cbdmMZBt48OrTR2Zc+wWF41a1sL17kRKJxT9K5jGy00ySOmv
o+vuPD0tnj5Qb3Dv+1uV1OnHL9wcK0SapeOlaG1iNT5UGGQovu6pzc8BI+mxc5Md
/HAMF8ugqu2FdrkCiq8MjK9uXzHX5kj+8/addBtmpk/wzmG1Uffi6WJglhTLKTB1
mAUP3mdLLCiNGtF1PZCnbBUQWsk8mzZpxfMNtbv8c90cUJP5JdHN2D0X8mdfUnly
D3qJ1ViysOjPfFhEKO7EG2cGfSXOg9Y0OFiaPsP9h6k4YNse0kW1bb4XPHlI4X43
Wf7dQUUlzY95amCt27FDXZ4+mE+tbyRSt7J6ThefI1H+XAdf/86VA5pyq1GRpPsQ
3KNHLiJT2e6cY7Xuj9D2weWJwqIzRnS0IjnWIKeBg/hIMvNb/kWgreGqUndsCfP8
BDitAxzZJBsMIl99qs494Z64w2AWwc8QpGX5sQsO6F1V7mCOmjd8RmCTjP56Vhel
DlASrgpFTL3ImRzpapMeMiETKbnVOtb++4idFqIRRxOgLsmWowooJcy/mNOPcTJD
rtlOXdkkdSK0Qxy40OCN1hgiT4dppwXoFsHZh5fUmFzI9k7FzMBT3ReFSiQT523W
Eiup9O/PQOY2NzhElJ1loQwBmnvrjMKqjjqosHgWML4x9gPBanxraubDmDiwhsMB
+2SWiP7o/qO7ilPk9vLED6BbvwnlPYCfltiLvVy8taveLTSEawZ/2c7w/0MWYzEA
9xNSKK530ZDEFFOy0uAT/Y5K7gd6ZSwCf/0Gwt071zi5UrZBR7j6q69Kom/z0zXu
Q7fH5H2HHlaXU0FbRe89LB3pgKB07IwvjkleiykvqiOCobYuGP7LpqKzmRtFrtRt
oHrwVsg21WtIgb22s9b/JRa6zTZ8cPcgiHYiCWYfQoPCezwmvm5FhQiCXXeAriwQ
A+S+fpwPAITt2SNWhQO7kLw+h2zpwFphGH5vS3MKBmtZOFPg6MBZIechbBpsGM7R
eB4Mox+Yr4gfjqE5A63Dm/UML6BkaZiU7wbb5bf96Yoz5aNVmTIzcw7VPPTnov4v
0cI6MxzEviXYTNhDIwkstQxz7t9VoZqkkqxIokC2NN1pUZDsJ0TVYx0/mbrHI6ht
21nI+d8BQutfBopXybLARpzhMPDzz/yAFBfqTjyw8bOHkc8/8k+JyoDVMienaILx
OY7q9Afjr7kwV/CgwtzmTw7n6wq/lLNHLuvZS+WLFz0NUnxZq3oQVjDiRChj8iJl
ShbPTLt5Xjr8oluQy2xGAr3E48wdlc+GbEv8e1zy4sPohz3TT8OgerHGdX4bAeLs
tEFC6c7EBepnCzkCdUB9RYl1+v6E0s7pkJIJS4D+pSUzZtTVC6qbxtQ6EPIqIpsa
Go2EI0aqpAMlxSrlGaOML20eAjEi+DXTFLmq6U8XeHQQO+L5HJ5dPCxrvDX//ZLQ
UVdYwiC9P//22sg6AhKeFqqiq0gUXZYF+fgbw+R8CUN1BVs/n3hLcZhVrkMVFj7y
7V1ZwbhzH03NSGhSuvSgGWR78sZHx8Lx8zCN6AsnCenllsYr3cESIwF3OV3yAGk+
6IwcKUIbHqLbzyQBx+vaZQFUvISKXG1N7k+iMR04iVJWK2ITzf37w0TscBJo8Gok
5QwuiH3Zhbd3cBXDVC9Vl4x6k1+j2JVQHkUL2cvVzhOGNgLImub8eMQwuFhzJas3
TgQugJqNv4t5tFwZDMedQdfeAdRu3S1Re72kNtfDHIloXqIJjKLQV1kN7YQOeUcG
fOpVsHaL8aOEJKygHExToYRg+sZXXdwee0iFwcIb2Xbvow27Bd/MJ4QFDN6GsHBe
ZSSVDSD8l7Pkv5KOg12SyOfu5LBRumHKfmaqEM33As0PWALSXcejYANKqzHEQZbj
SZLKHxT+71seonGDEf3ZaQhYIyzWOmkRUjOWgYTkb0oKIoZ2PY8AGwGjr1x6KiBi
w0EYGzG6BsfecXhFEPTTjPl/NDN2cHB9cT0Gj3xhkTnbcVVnBpaH2VWy1jgHcrzO
sDWCcRXztOMWrJ7RKSpqIEGI6SDZ3JlNSXkfUJdohu/LLlpBbdAwS2Txshz41d9F
PDFyztTd086ciKBEHO2AQ2q2QtMONEX7pmdaL3rIDvCsDiTxMyD2RNIg7vi2XTru
W0gF5vk0NjdPbqgkRLhr2XdTAxMP4swokEESgsllJDhOEcNm4aOMa5VWjkOZwg6e
LGP5MisEP2YaN4KbOPup8ZgOFtniKVun4sg8BsmvilAY/RT1zde30LtHeL0R60iA
dsGn+AplSN26BGlQssIGEcfwl2FMK8ZnQtH5QH4+ayGebo4SFCK8eMd5TJ00aGBf
8UYUbtsYdtW5RXYr9p11hmY9qANOarN5XTUXQhmybTgz7yr3AxTTPGZ6CnIbbs14
L9qI5gvcl3l2pe8XHOdCYrQX1Y9WbawpolJZGoMTb64sLcmyRT3/VOwkz6qtsCRL
dEDYdxr0GvmUWYD7ROTnksjz7u+vSO2npgbtPjAN0wsnyBbc+QHDAZmAZkfyQgMq
85rBMBAkEhKgOc9uSHRwMf/SzewEw6Gpz0Og2a0AzzsF664uj3/GOeLJNKdnIZkq
k7cRaQqGePvG2yZSoFvZdpob8lIwkcJpvBcIQ6Q+w+yjzRnuT06dyzhcYV3/TElZ
jD6QI47i0aEfN0bwuYeAhD2dHr5QaXt49vT0hTUf5fposshomjl4n0aQzE2ijqV1
zhRY1Uk6duRwnxVUdE54FICleMFp82PanxBbwM5wMnTw/sHf0PyLq6vFwfG8ErYs
RG34R3UDcXgSqCwjEVIHrAUuxi/r0/hlJhl7f67V3h+gG4kzzRK2k13MsausY9NU
Fr/hjrrdGmwIMudjou3q3wKbZ3rhTZy1n2PrkQqqU3BiEdgRY1DbIuJ2GKaOl9cQ
px6hlx2Wkl1EGta8mIJZpsxBtdAFt1okDPdupwag/r2lqxNrHFJD1BHlAqt8bP83
PxLbFp9r1E84aF/1N/0X8WIXTFgv1bD5GXQlGQY7b6On8/1ba404c/0tvwrYoGgM
T/dqdhQFzOBFpirSsoziQf85g9Lb6lR2HzOMUPzbhdY9qW2ShqyKlYuT379sLBzq
aOTeSWs19SxHJel/ZntHR56F7/45YWdNeAWDtSNxGIVaxMhfiKGiYaUYLoIiEvbA
+9mx3i/cRbRunUe/MFqSZtWD+KHrHU5tQ56hXSpSXSpf+bYAuy95dWKD4VKujapq
o2sXpmJMGhq+wXAOJcebWEHq690ya3ePRzwr3og8L/+2tNXwcZYU1fb8huJ2NpR8
VwtPuMt9W3MqJGGyyBYc4xQ9t5YmojBMzdedrU0y37mgvdZ27n7YhRpriF0yEzMh
IhLar/YhhpCKuPezyc4s5rb2O5Fv5fpfVZcBS3JLApISSpSjW65EImWbFGeb6fMQ
dJRmjB4JFfHS/ZXPaCmjR8gZufDqd8UvENxTtOJ2n/o0EmF3PgzPJXgFZubaqDxq
KLPfateRABzyMbL5MuZyl56/SFA24Uvbpc8HCypcZLQtwEHTa7CqSyQ7UrxbfWZK
uuxo6G9CZ3jPXmQTEtNoeCCWHQf+Wq8zxiU7Hl/dMSSjykLegucLT+pMNz8ql3Si
cnMIq9aq+2yDozVmUy6X1pBSp1ABqoTEFVTfI4uvBpkXh2kzr3uN4leqCUfTDU3E
yjFp789C1QyJb2vcXsrGKSf1WXkpYcLximlgEUcCnUgR+gsB6Bsnsd1yOSuZAH/1
Ko7u54sqT7ubQ8Xa2cQur0/wVrKrdyVPttUoPk3nVAjEXqhYP0UHE8ACPzV2fWZE
lhtxHhhj6Au3KHFYHkTOmctCx/k5xMioQBXrlPPyrKsvZx+GPznsks3KEzdqZaoJ
uzlDx1xjeD2WXYtqVUInED04PGjwIxsdh9F+PU31cVWa1n2/Z1+wKId4VDbAtd4q
6HYYbanlcxsZ484xCLFe9ouwoltB/oqP3TGfamG+c3CxDF8DPEiHa20GfHNAZ3Go
tAtgpvfHIx1Ub9YlwLhVMskn+tkqInb/VGf9Hu39IlPfl1NHPaT4jXvRm/Gt743a
AsdTgZ42Tjk7rzml6ftCB63iW130b7IvidK59PLHgQHrViieS1IbJ7KKofg1UOf+
C7IhbnpQREgKSdvRYUFLC8MC/NvudcC1bHaZja+PRZwTfQ/n9l/2iuCcZuWabXm5
b7gvhoJusHU/RlYniaEFbEWhD7IDUmMcMJy8wPQ6kuMB28FtkR5h3wcyfT5iM9JN
cagrlvkw0zWgciiiPvl60q2ihwGBbUCpkAybfp1lfDkl+hjdHZ33VzJItGj9C3+4
Am5Xu+zMGMKlBRIio/D9g9zTv5bH27j8PSZgKX2JPnpQlCx9T4fn8PyCdSpLqcEN
hIoJLsuLie5452GUg/5QS9c89jEYDl6FZ2SNFULzHMm10RjGuKRj4P04NRFdMr++
SYaQ4eIlz9fB1D8lehTaBku5CNwjzID1v3mVDavUobxkBSeIc+4kRpi12lz5WW2P
QxpnsEbR2W2rE1ulNQVnqN2MWPU0LPjk0iSO8a0AZMskfaO/XJgIp3RtNHdiv5pu
xOYfbsAbqSopI9wPVoprNv8guTi2JyQbABcXYAHmBd8+dJ1yD9YK7dnFJS1Z6cLT
ELp9B6C20of9o+MZvE3UHiiRL5aQ6qoGW4Sj/vxoZrwPK2wsF/ReD3FXGJyyt74R
ekg5l6lFDM137JvXefVbd2NPhCZzWkV3MuYAinmAbrEBZlt7IC+0KRL15lCyD3Uz
ek+BQT7rVWht2bDQNUDLAH5/pueKTYCG6xobNF2O1egxSqK6odOLOxTTOW7xXRiF
8h8te/UBUn7Y8JljSAtafCqyhsvzzzckP/rzQ5tYE0An6CLGwZlrOEIUtwz2Efd4
sSv2VxuxFdV9uXhJWer1M3rbJDBulPtJ7313bYZ7/jltUDmi4QMZ4R2NwiaA2cgB
S2sxvtOqm8VrggMuIJWx6ccC87qMmuno6RRRFCbGVqcZgwFdg1Bu8UISkJKdMsQ0
Yoh0mEdgv+8fMzx8bvzUVJEcpUhWTGodNA/VQBbdxoUC3MPDQTrRre0OgrInmyru
1ZrS5BlZxswv3I+3LF24wDOFhuUsILpBRYSGYDCwO1eHM1heGVsSRTz0OvI9o3/p
JUZuZvNC1185ime/bcqX/thSD9X7SzQqbF9vozO7lj7czHuFizCGB9dHevL4du0Q
rW9StFHVnzLK2fqQLvY51Nvro7nvTuFQb4D+XTOHX2fJXfhSj+esRdHjYS5CDLgC
cBGosO70xLxPzPqVSCZKf83i1GzZIQ5dFnjkxGIdbrX3y5pdLDlDVpPb2t97k13z
Tryjiyq6q28JHbqMKuMn1TZWAb4V21Gt81qTjTEuQqepFK3fULyODHMFuUDxbN+x
i6oUTQJTm2PwZJc5TMbSxjtP7/Sy2gpL/8TuYpjvtEXVPo5hi52xOxTwxtNXG60R
4NYMG7m4mkuLQeCKzb9BK685FLsVdgPm2VlJlksM+Wdh2u58zJEF/DvqhblUytfq
MyqJSdsvpdkCqQcKgKl0eY6omyhDNL8juLDDDaAjedX6ZJkWNfNzHq6SNFAkEAta
ponE186PckqUrqYPW420SfgacWvSGvbBhRS62BqENmwddlFPdpN2U2pohI4fQivu
RkLpu8/OHGrditT086Cgh91qHO890aE9jdqv7y1Sljrax+bAEVvQOKsPoX/dGpNS
4rvyVt3Q4DW1/pC6wMoRMsRi3BMvrRaQ5YtEWxLAwkdPM4nunkvTr9R+vocVDUnR
NlJmBhnP84Z20rCJDoZQxJdmxKoI89amGSK9GJ4ee3GvUPl2a8z+ug3XrActNToW
uYwyW6W6tMHATojIgomujCDhJADk7F+SEF4KDbHxw4Iw08YUqB7E+mH3ojkRajkn
yI60O9HcPmVWII7SJ/q/W/nJUo+HTS1D8fcuHVUj5c9ITX82qRl2fklGKv4tNxHl
xSU0ephgWJKECcRs++dJbf2dawMevZy16oNmCgrTbqN4XZJemZAzcFL6/WQ3g9za
kh1KGtZn6MT1aw5vUSqFcWentWUgFOvr1AM/V9eynkzi+HOvE9ofVRdX/2Aeyygu
jfvG9rQ2UHPQ+rURuWt5ggOAV0ZEsKRpb+KQGtPu5h9mYWOIIkcXvdeNwyivMNvg
VqDJgNjO82UnNnwXumH6nxHiqWxkIabHQhUN+3N8TdkOK0SS+6yF4yyQOgQ3Jmaz
CmWETP9zsQY9rB2nZT1JszvA962JOQ0cEkthCEX7cSlL+yIc2i28i1UlPxT1khUV
I171osxXxQvOtN6rxh2JsLwVN11ImN9/JrVQpVVpvfdIP4CwfkUDcdBnS2phlVVk
t2+HkdQwseQ3sXovwVzKfdGcFdB9rzscUP9Gs4wsB+v/wEBwHSWzSJ5wB62MOF6C
juMi7t8bQIG8VB2xHymZ614OlHxxMMSabbKWz0COgCLzRUiGrlfID3DGebp2tYsj
gpPeGIDo6NpOpdUif3FC1DB8jVfKdFbm/0bgD8jGdvNWQagrgP0YO+5OX4PeVbKM
37c/6ZDnA4f3ael7Nad5rF7VtsgWBStTDNfj7kQv9MhMkoQ54KWJz0cRrcsaPVhH
ciCKJGWVwL/15jzQa+Ej8IyfJlShRwptbugnWxQzPqmkm6frL6im53cEjvgTf7VY
72pMKa/dhw8LyG4AW0J+P11FviC2Rhi5CDPvslpMXJTQ8/RVrlWgoB67YrbJ0o/8
lqA9kXZtf5W3VStixpcTrPpV7iql2gsCx7u0mdZ3FpMx1+8r07irY8s2nn2+jGFj
PSIpFUk5Y/niXFIDw1i0acIdjrH4jgb9WOtIIb8Y1pS+9MSVUHX4XIy04RCH0Yxw
3dAdydQlcuXxnoY8SiQhmLjWYacvEsopERavd3DmMHiDTeI5Vk58Fzcu826oP/hQ
c4epZmGp5k6Q24ySH5SbfwY0vZKGxoqwQvLtAIg0r081Weby+TXAi2Utwp6TPEeN
cUfgg+uBz98ekNdhJ+V7OoJcZNR6dr/9TNhy9qvu443rhntYjzHHUomFTbihx/0t
XYrJfpKTrLSMBsi85d6w4lUBqNOzaBccWL8MLBzNrwGMevzjK52QoIIHVXHjkvms
CcNhLpib49kYStXz8EkUP9DXSpkxPUz1R/sJ4FontsrKpbqmJoUZD6F66Sq+UrX/
i/6WU9zshnBsDdMJlnkkrLw+2t/aJAogwS6F32bw4Ao+10uVOH4fv3336f5to69k
JSfJbK8LLtmtgl6s8p/d8BdD/2fSqrtYGL5pG7NChiEplfxAdmKlG4OzSwDp8SQi
TEYoQpCfaXdJKkyCch33N6Y7QuyunT82Iwwf0qJM6Bt4bZ5KMjzDArYjuLMRm+cL
q897yH/LZts4fGCVv0Oq6qOS6q/GiAxumGEzsXrhI+OlAdyqzFDCTwJocJEKeE50
9f+oG9ZBVW6q0VYZ7hNNjAz2mD0sXy0gbV+NrIY8KcAYnL4Gf+xbdmRS47GgySI3
LD3Q1lDHulrSWpefBuevk0H+Yr7NJd3LPOPrFYXOd0FyFZSi2927X4Ivhz932Gwd
/LzVn74JglbfwVAyjWQYVW/j9AhuagiPuPpYTkrk67frJFsowfbHx8SC9C9vnMi7
bpypcr7hrXXB5yjOaUrJ4366RszNFL9MIr0j1leU+i+eSqA4bUh6xw/y0rPBOWcQ
rmJgYjUFxrkwTVrzdJynNFxjlI0/GsHHcaHm4OQnF3OtT7mpJ/r7U6uBjCvD7k3V
ZN6CXxeRd2QApRFXzNRhWeLHSgW+eIkFpjbfWuBekbp6RlVpxMC5ZUglLtb0wR3x
gOtBPFbAYxnQOTAUfPw5+eQ+rrYsJ05urAf+c2vS168PEO823jmSGhMXroqQMWh2
Bxrm0KgarbYVXn/6d4cOhXYe+/jOu1aYhHB6ti/0c0IdtM3lqYcBllQ2e1PnqAq7
I4lVXkQUKG4lkrt5K7DmR+5RAVIWNSVTFVG4ff/4G7ueG/CnnExUXwGnUeG4OzUz
Zt5j7RWkYK0l3AUdI3eTUF+2tWTAkST3sQNx5DHgvmIwiOGyGVxDXmaqbLpXW6IB
RfvNU80MsmSrHFid5Fk1ML3ICzzXUjh/C/hZBwUauJW/Mz6Oo3NVEF6HGHw3CzXt
LlydORHp/fncR6zlzrSUixTBKihckh+vpUwDaY1i8pGBhV0KYgZZIz3q8xZ6w8Qw
c2OS9iBvsGCw1Ya5pHsm/fGJkx2zOWnF0KBx9l40hvBToG9j33mrTiW3uyhuDbKI
HVPLtUVucoP+BRl5bAgxW56ofKqQ4ry4Gd+haRvPEG0UCahBxxCWMymnyi7oNHBe
+MPQq6nlSDxZRhvI4VgwmfrIciycaTNnlv0mh8Sq8kopOErtnedQcw5f231ML7dH
JIuJpSjJLImVHsGkcTMXg63VCEp1ZCWZXUKfpQRNuOIqNPz0T9MdO0iIu7zI2F+C
ET/FMN1hBnmuahu3vO0pqbiZdYxfdZ9/9irS5pAfLzkI3XRuVzU22Moi8TkgZGBK
hv1oQATW+3axTe+i8C5911RDXcLC6Cn5TvbP9uPrWgu+Ggqj6dkdsyIstTwrHfzL
mxGp3yLIQoKUhGRt3i9IsI9VxkxZFtPaXeHmhev+YqXDhFgvEOkZx/0LbMW/TYbx
CiioLhpkLxjzD4l6EmDjr4rtl0e2sRJkXwChuiBoF8XtR+mYnR+cbewE4eaj77X5
s1elCk88+cZTiBJufJJzr1lqdGew4DgKg4+YZcCj+FhLkw8s+5U8DRj5XS+fuLro
bEx7Uzuy87hTrWzwMbfM4JzYhRqK/xrMmXVdnCBvcotLjjiEBY7cw+PxlfaMsCF4
CMNf7FnbyqqqmO9h0D+XOM3WyTvd2nj9RauE8P+7VRD6Eq5kuhOdSBJpqAQ25CTA
8vbnV61Y6PTf2dqxg0iRXYAicfretHszc5Y+ycLUiuAkvTz1QlEx8+KQ8gTabUhx
PR/z9syOEnf5dctNaHp3mNIhibPE0TYzY4D5rOnRLodaX9Ca3nXqR1rFCvkIvboM
VGqfmsQGy2SU26Kq5tzLlof2AvH4OhHT795f3E/6lk2dHZaJoKU083dUAs8lUth0
Hr7uPlIoQtJTrX3Kqientk656y2zONTLNmNsaG/lfV4/XpM4/1ogMe/iDE3NPuqR
6XcZNeXldLpsxfETU5ulkScpxlTyjtNiGioFdJEaWEy2nY1DjTZ6h91sLnd+7Ltx
xFBlfi425c0UGAIAzSQ/xr2mL4DIs+dCroYwaIhaxF30UmnRMclBViYQTuBeIH50
SzNMOh4MsaMJMlXHyR+c956kMURiuQBEXRjNAaw1tKt6y4xxmPywATC08XRUz2bq
ZGLi70AX3HpK/eTzyfLR9F8VusNvpDoGWWU3bkv6to3ihAllR/2sCWeVfqEkGaKI
5Ix83x7nFqYd10xNZDUZH0Vq2dozuKpu7T8SbKBaG0nSymz8oPol6zU1TdTNg04Z
GRnm4F/qpK3z/StDdRW0i32BLm+A3ksxDIOrtqbP7AYbTRVkOsyLTECPm4gWYDyc
hz0XEWp0fDvMHNMZYwTCDDwA1i13Z3DLoBa2HnDY4lMdnZoZ8BQnpUF2jJwrzj+Q
U/nLmYCvQrK6ITM4qXbnT4tTPC7Lk8zOXd5/8L2xIHdK9tuXFoCaL03vNpqqe6P+
dXhQasqjPWnG6kia3ROPliBD/w3efEtwMdI+uirdv7URRNklZaDxgBcTCmbj00mr
wFzWm9h/Sb+b5A0H+UeyAKxT/EimLVlJMnRdevUZM0SYa/urqZitR5NR8wSYni2z
AnlMBcFyTip4w/dlWbcCbaYeDwkrVrabIbLqGjDj2WY8XafzFVog8M69sn+E8ikm
1lM5vIH3AIWbuAEMPTZxTGZyqupWz9BbH1BC8GG86PU3U9FbaHCdfEMb47lUDTTa
fYqReh8Dyrwh11Yv6G1xboOCK4pNBq/iLz1UAnd1HD63HnvnnJyIXsVPHdP5yB8p
BEXUK57Pp6tMcAV9T3l5c7cWUWr2YCdNi0jmumFWOntjO3K3K7nn+/G8RuA6YWAV
c9djfxxbRRCDqLFfRSln9xbl8kkcg8igR5wSanbVyXYSEK5m53rwhJVzv/zbeBew
Dc4JoegH3sN6jlu+0Ild8uHi0kIjFy6EziHdJD5f+Ev5GSjL02xI2/WNo2UoOvg5
lLMeVq71xA6GU4QMieggIX57yfedpmZPKAu7Hfku6FWz84a3iwYp0Gmm4/wH2cCK
UxHeBy1vz9sAFEEuipiHl2x/9j/ju4n0GHNKKunjBHqih/Ohoc4W1In1+KYxxZXD
sVQpntCzpvTIcezrGknjuzNSX3sORtX4oIJSN5txR3gW8V64QAY5ASPwxQ+jD2ES
pqmHb12oWcm2kQnLEMvUSKz4AY6y793AS5xacv1FCvXkSsvRg0PIFxB92L/bOwOe
MaXJ31FJwT4vhiVTq4Z+bIkNPR8bpQUGo/xPKoqK8Wlbz5BKZPHhyNZ35aWlECEY
oOdyREjrxhlHZs8IamnKlpsmNnqEA4RJtO2wGGkewaB62ZH//rir2logaJvuhzFP
n9/zSVppVv3BYOiCJAu60Cf3px25EILlceNXcr/XGYl1RSVGwC7SBV7HaGJiIP//
3ktIZsMBUsa1MF0sJ2jf5HgLSpUGUEo1pu41keEgcxbvf2HfsguksKW/+G0E2Yig
Eh3s1+F2+y4q/NIsgjZDzTt03yu4X3CpdmBX2SUN9Bz8kVm+50Pw8Fewm9/Ev2bF
kjQ9ifxwEuLFlbdpUZQd4rHN+cL3gi1MQP0hPBrjkIvRl6ZpIRtuzr+lkJeGVTix
6AXGDczJ9HIvZgWftqiO9WTHjyZa5Lle54EM6gF/R7bP9m3czYpn/+D+iWpMm1jl
7P/LF7zVc2ekReFCM4FAcSIZ7PJHwtlA+j9xoozTAs9SftNChTWkROWnw4V7HxRO
aThBkZo9HqOc2/iq9Jdfi1b94ER25gbOiaPQeGh7vAKVumTIgtoh7KYX4ox7EpLD
uFmFfroh0ur/znif4JyYDCPalQzSoSuytRR4SM9CGowNkCKTASo52YrzT4EXKVrW
3McDdm3prS65WrL/kLG8PgVjCd8lJZozgOwBO7pghXiqn49YWi5eQKq8/SksGoUa
+UromnLkyJmMqkZARzt0QNo42mE9IExR0iaVs7Zlg0pzSsZihBBGMhJ2aGp+u1D7
HcsWKJikEcSJnPkIE0Bk6Nr1Xz5tPc6SrdXogW03TViHJvoJsO623EEP7oLJVjn2
KWVwvuTAVGWZtYTTnSMjFder88yNQX1MeUmrVcw51aQVTtQ47MJlRAzVBmw5XLsp
6gKNgZcRAd9agLmYSNfjuEcCDeuF+liG8D/i4/7PLxnsiKi8bm4vAdPP3a4daQUF
j/LKt3LNBgU7tjUyWx0VMDflvsUe3yobat0RBHAbYlqGbQ88vTWBWQlRofssDdi/
QoUm7HNYsJR1NI4wSeGy/QjC4W6/WSEJB8P528BRme9va/PzeQDebEbUe0ZileK8
6YilfVRyvd9GkhmCkA/REppS9HACo3GhYjiFc6kk9cdYX17ltCDJ2l5T4SRi3766
KedZEMNHN/5/F37qjivUgeuJQxSZ6h1E15iYo+SJ8e6M5C1Gc0/fcbw9gECfftK4
VDzDtDANzyw4ahVKckKyWNSprRu8hp/Z2NxnvSr2ji/OfPLOvYjt8zvpzKquEXUI
t4naCyycdaaZLXUamqcdSaPsdhhSphiKQ7cZVUqGiaMGDcfxiia5yD/+InLrii1W
3j9lwqG9WcPZexDIMlXYRqjeWAIixeiyV5bAfg3l0+gQGI86Nzdj22iMWY5BsRsI
BT1Dpug5GNCBTOIxp0I6sD44iGsdpo8OroiEp+WtyzBqVSenDwZjA68sVOBW+hY+
t5+5dsYc/mVyjRRBGwsWAYBtD3dApR2uIDjr6A+Ix4+rgFn7Jah9TMeTaKqwe0Ou
J+YNgVtQuHPo5CM8C4tqeL02E5OEpNKDjmxLrH08fODUWmjw0yV7rlm5J2V5g/cM
3HhoKNG0a7it8sBS/3yBIwpBzzdnIhn2u3L+MAqklQ6tqwtFFVDrs7Qst6cDPFkC
pcliCGbYNVC5sxitUVJWB+5J56yrEjaMErFklV413DRtfYEYoWjAk1N6luhtSqY9
rKG9Ywmq/DAu1+AIDLuF5j2H/fyD/OB+xfjlxDZvo2VrVdsGD9zcHG0BOpHkj4GO
1bJNzUd/0fi40VMA+8+OXf+nJ+A/ioH9clTj+OyzGh5QI6+VjkB2oCoxiCc+FIb8
sUEbiAdWdNQQA5zE7mqrXOrjrKsN+gQi9/Y2201Rl5aqcYZWtw73UzwVoeJS692d
1Zn3rX172QevPOdXUguE5h9bSSHZMGRnhrhnqCgLcIe96uBAQFlaeQ2xX0xlFyDC
nxjLZjGjGGbMpGQ3f5nV+jLYZIB8imVzzlXsmQX5OFw+icBOuX06FDVwruB+NRNA
evuB0aY6px/zIhbcKH/K03/uzgHy93eQ/XVy6u3ZGL6Z8fcthSRks12EmucDdaDp
ZJJtOzdVEdZ+Ww8JGSpycHXfX6qNRF7muu1QMaiZHkCtUZliUyds+7DjloFxMQjr
zLjTt6A8+4cnX4hdl/VBApO3HBYIjPdGEyyxVPq+eJDB34eyb0i0apRw6YW0i3sn
bpRzVct/M9FXHdAv+FLNafdJQ9fvt5dtrRn4AA4VsCOxlNEB2Ch7dN0/4tPDvMdu
e2rCnBfTUD7Kn0AY5e9lBaGcYg6d162fPtKtv2W8vMhdiHuP8724l1NINaeQfI+q
qbMO1AQC7fEA6qzaIDZtqVAkp+dFWhcl8e765+EqYx+F3hZKg0r+fNFOg67kFGWg
HzZLCDKpjAY+tdOAF5Oi7wfsecgd+TDUh8Rp7/ke4NDXmArB7P2VWI6+V+jYZhO0
EjpvkpLct3YImqQlXQIAWP34Q40AcGufZvtyh7MmsfD9J6apCF65oX3Ki/h2h0T2
yvmK9bTNqYvWxHS6CLwv8G9YNG6W0wtxMapA7ylnV65kTlrCXsWhXRM7fAAA2uH4
HRpl87KQWyPeh6/y/k1UXBBLzW+RUS0WlmBE2nIcT2Xv8Pwa7CAhkDrc8qPfjHRS
whMWs4suIhPS4iRwZdWTZZ0Azw2WdjN9Kzlm7tY7vWcQXurioLkoV0MSChyKz6kS
qxm1fu96ETDZrvRgCgzzAKUXP9utW6WcuyfceV/0CUUhcuHfTMEpZJUA3qmSzKCr
xeAmOgEHPpIubJhdDZAbXbIzxitaRUMasj4kUFseSEnaKu7WisLu0e27g2rL7fBB
rPAQ8g4zT/JI6RS4yChhfg9LZ+2B1bptVR9by6dz9ToeQPyB1cd/RoZ2LPWX+fc4
xnCvFxHTYBUr4k71MyHZa6NJVvE93+WxaxQeMXhZ3eOJzPUbQo6DqB0h5dhzVryv
Pm9u+32KWi7ix+yLIQzcyXd9zzA38Zy4DXzEjqdJHIImAiAb+iz6LzNkzhp1ioJM
cQ/bRU/KmnYwVztf1/4YIbfglz3mAKZFPxYEklrEF7ADB7wTg55BawHXwLbR9pQX
LnMV/7hORpvfvLn9MnQfSbe/6QG6mk/nJId2N2q8WPVn+SssiaB3S2lz40HGnm8j
k9MiQqlXReFUL3Dy/Ki/pQ8WVLgUW64h3WDIx6xd6vBERLbm9MXtHLi4uUKTVk9L
YaAzGBI9NK8O5+qiZfgPwirRggRosOGxskEluujjhMgdhT3+ximY5OYJ1W1ejYzK
ixibweODhwZJOHKoWnEI0JqW+m0e/Q9ToIgFULFaE0ERMY77a8zFuMTHwfP/EqJn
v6hltCDeJFn279zlfoj+flbCjUTZLegAvs9bFv6J10fpU56FX3/YDs9Xa6Ke+GSb
TXZVHTtycwjxJ6W3x3wYtBpfhLSncXt9/jBk6OUS5JUn0QknWdqMqc1IUO3Zk4ym
X9YIzjY02xRIQPcST/Q3yQKYwrBDtXDSMTnbJ0DSHMFiBPybHaYOhkdqsKMA+ffs
e9nqo5ZJlgLxzQsBp9nF7GmqNCB4MY/x7ILdIvr8HnFLrKO470RsA9Kd1fpqgyVx
epo4faqhevTRZBW93xBsESBLSFmwkXVshLjzccF7XGtDB8p/0yQdRp1Vs5ob6CiC
r6mOUCgrRrinYfDpXPNpkYkCCxI5g98Arit43uGmAPEz56NVVFKd9HVGQrlFk0vT
sTn5HAKtPsnVsqQxdxBhFre1GrL3a1/twOb3Ja7ZnSn5JXPFrwHDhlUCjJjLFfkJ
XVV07j3yg/GTwuB40BamPCVVGZhI1xdJz0CE2WiKXDQzmg8oZ/o/7/S12FkmVAl8
hlCXKDqOV2UFM6FEv+8ec7m1q9ne52HfP3pCUF86hOms1THIJIy3Qozv7D5sCFif
xI/QVZzdu21YcB7MbnBBlZTvLHwoaiJwUIchPD3YbJ9PYoUE0IUtErJOFgWh2G7i
xr5HjFJmZGTgnh8tqQu3cZTZMKfC2OatFqkOgLWHpymKpYpCG+jqWKxuf92+8xhQ
/vigZT6xKEDcJfqlh2czsi+E3bEAWuGJO9vA/p+fi5PyW+cC53orXaQXGbnjs9kd
hDwmlrUfGnMGjkGg7OGy7T4h6llxA1KTHdU7WxcB5UDq7QrJOex045pY2vVtREPN
T+UUbM5ewMN/vNJwqJZ+S1f+tcj67l0vhGxkJdd2NWqp5SMKdmCqc34eBEy8nqcb
l4h0686NOhgbfOeOnwmDQjRIjubHHNW/wBDbg3MxSrYDn69IAKnvoKbTVMHy3vH0
o66K/MT7li/5j9BUbsmGKdLArafSpttV+yKsvf/NzkodY5DROtYwiCUVLRbOG3eA
FtqqJj7H8rS3ITVWpDzlSEiPw8rLveEgxUoa7EwqgtefTI8SfvcHPnd74djmOD4Y
E/0pcZF9wFZG/ipsWIrPvwN9M5amPjTf4dld9MwffdiFdJECSpftUesEoXyhrhra
1FJmLuAJxN216sRP2ic9X/DqInW/v/6CMDj/gaNraaoL5Fxs1hijQOHvE4l1Y8kp
m6R8QwxWYJXtmK5861q3r/Zj4vix4+MHXVr7p3KZfck97NU6Uyae9ndpB8HXoCyD
RSo7195DRkIDTGpMAKnuYyXB72VyF3DuB7Z83E57IhyK8OLKUm7Vdm8wkqj4neyb
9/W5TTSfFWFlOmS4RkcvUwPTb8AlcGveSLACzDNx++HGig21xpUG/4/U0WCmRhCT
DSWblrc1W6x0tfKjGm3JgS7MmOhzBit1KM7rjcFWLvFGv4TM8CIqzV/gsrLjM/gs
MltfZ4B5Yv0VEtdZBgy7IsqMM2k9JrWikpfknNBYjp7c2TLSfH4C+WOuJjmn4L1N
wNH/F47rdTUouSoF46LdKhwrIhfwMyzWzjrep2Q2o//IzoJMjYGrKptkUyqAg4fK
aJYJWO4m9iPftBsw0htKZbJwxHmi+SyS6k4NKVqNYAyUnyThKTns721R2C8PGPka
moVkQKBJOpDDTLY3T8z5JhTaqVsnkAjQCHwZ89iyNMVqahxo5R4IU04nSQGadPwh
/hBksyqSwEG0LaLUyLWT/PxPaZCsLbjD6SMmtny20jsLCSTpyqJTbsOL137ZPFPb
tMp8ee8z3esUaNdWXNn8ha43nfD+fRXI4mfAMeMlUi/s/obzoK+4opgLcRl3UbTk
Qb9o6DTdgSOVMHdPVQGP0ozjIlA+oUk/ppFQbd6RhmL07g6Uy2zv2yfUHfEtt3kb
/O5qIoV42UkpGcScaBe+eaVMXKNwOA7vISGJJGly30qnWnMDkuhu56oFxrpEbgyE
VK3AxUdOQJmYqwTDO5ioPn4LvugLrJm8vKU1GtAPgl+XOhUsrWEgRjzE9lICjcl9
oriHe2sKAnMgFhlyGS0mTvxPiYfjtYJJ2Ig3GjJb6i/OkbT+UItwedLBSUha7ENI
Rervq4FPRufkJfPoDlg/Zy9K7qISuIhCiadJTf0gyGZGAOQufJDxTeLDaPuvuj4g
KOpree0nFfFhZf3HWd+Nm7BlfP0YvEwWLo+ALfUyoB+DXOWn2YEAabQRRjbGKdW9
ne+Evy/4bE1P3I3C76pvsAvSv8J4LQdtc9FtF4SsehRc3SK8OcI883rA1zVAiwq4
2SCnXoiHJ1ARTJtWHc2AzusrFRRqJVA4IIZDzPsqIXGKWvD7KFt1ha1EBsaD+tsd
bWoXoGDZGhrUvkF9q3t758EdD9sWg5wpR2+yUszo8Su/hIumIiiXnL6YhE9lOElN
2opkM5KZo9oaV53YfAmewCrVKXAzcMTlOjkaomF3jlYOc7VZY8XgsSeLVAq1xMPp
LrJNdKf6sTSu9xPdiZFPu70T+VTNGeBHs4SGvESIoDqk+rgIZsXOnwPYtwAQJeTt
wsGwU5wWZu7RtpIM345xKXvS+YQ/4f36/7MoSAuEz+2hcfQtmtUoYXbHkyohKztE
FOOGbXscH7/Sx18vqjfLE/NDJRHoBMEVAMRzMJHCO6LyB89kHV5fZhG6J8GudJuw
5y8s7C/kCnxYh/TdAL5zrSYKCZ57VkcKzg9cCquWzBSeuv5P8hoOF52CnKJZu/aM
nenx6VwEvvox/AZJyoK0kRYjVKmT91ZoRpMg5/KNbNRrjVW4bqz3Ss+rkqFtWoLm
XJLHkNXFiu6fZ336mdqevW1o1wykdEJx3pVXtTpuUcZoxcTNZiRRY0E+B/qBNIAm
LkibLu/TTRB7jSYUl8CNMvd93yxhJYqx0ph6UnGIx278f1PC01iiaWAXTsNDCpc/
aK9+iwA7pGrB5nWJAl6l9BjFXtQI9JyiCUC4lBigNCovkhI7c9WMOjyhOaNscG5x
hUtRfc1T5iVmyOLM8fOWPiHivAf288IZqn7LdCgfw9b5DNoOIY9YSkJ6jcIty4rm
UCG9jAK86zwbATmeG1DN50HU7/QkvgIUdNtUz7l6SHKV/Db0uNZthjlyGiRDQoxX
VjUKa8otgf2QIxP1rMy+MsK7ay60174wV2i8znH3VNftY0BZIO5UkO0QSNA2u+FY
67t9naZ07g9VcjDg1wZmKKg4ZsxnnlxRrgViT+LBubqcho7tBX1VjMxPbvQeOz83
nVMPM8j4tdxLPyB/SVUsV8bd/irinz6+5umNmOTodml0lDES5l8VQEYd4T8scCSj
IRu/HjgrLVIu788oUbjp/69otdfLRj+ehT5QUGN/YGVV3KrdO3dDIpp2xqdTjvP3
cpJEz7Fg6i9SpcUKPQWM/coroKHWzOX6T+CrfF7CZknZkJBaDPhfRxw3j8Nz0XOv
ytd2FFc03ehyYB0swhlxSB6DGC6QGzw0p6q5y0ZYK5QRnhsRkw7nNdgRtjD1mTLp
JAwf6yQ+zcf1B/D6WkEFDXjzFCvnlIOESqWccVWAnu5ua/W9ovnuMyvGlKTR680Z
Q1kUwl1CzRC1eaOPR1xbtZLm4gmOh5a/o+emkVoqJZG+dA9AalWIY762729mjeC8
cXxGEN5Jo2tJqq6EznivxOq05TGZcJ2YeAC9WNgEk8ed4hKvLycx9ziMvW5MiuTe
k4YIFcWEIF6464OntM5dGB1IUNgDxQQ30vstJV6ipBc7cs5C9Ck7r4qN4Neb++Yi
BtcaR2vT+zWfb4R3ztAaqjDIiX6GiyZ0vqiS0q761dLOl5hOAMvfhid+YNlQZrxx
sVdUCjXyeYT4ylzf/tMdAuFd+f6kth/sAaxlpu2UZ31vZ33BFxhL7USDTFqthGXH
ppql8WuLbrvPd2oeTVUkWhCyx5qTwivZetEBFBP8rH406A7h7ZUzNhGQaCfkbHKv
uyaEHdfyPe3zAysjcLIdWp5N1N4h1Pi6h8I5vjA8L7zRukrrnGaIO0TSDzXtzSWm
VU1NlpT+OFZf7Ea+KnGbg/Jr4vBR7wSVzwPhsIfb9XK2an4kS0QBBR4m0ZtxgTh6
/m4KtXZdMzPt5L9pYkhqt0CloniWxj3l8bu42q+uP/y52Vbwr0LuUepCJw1EZ36Z
LSLJARiF0b8mjI/GNT8pEjPki1aBPZO6GEGKyek/0jOyFBwn3+RYZInQh1EdpjO9
C0pYHaLKcOJfU7doPubOz3Fsrg2uOql9rvGArAZclAX6fUeLZXdGogVmXJG+1Pi4
Rq01XfNVuRkZ/RUXIDmb9HmfZ0CAmmC+MoDMb4DLV07YIo0zOj7MJKqhTGGQHaqc
/cBRYg64tXyzuihurvcggla0Z5E8sJeqwKIxOF77+mTc7JiR7PnsfNIHuNlECFja
e4DgarDkr3fXGg9wRNj5veeTkWTwXZsjBPXbWBSJ387csaKQrbmrVXMhvHXXD+OR
rRLZTS/CM/LugoumPKQXcJJg/hFriQ2xEEwtKL5EfHddICgO8s8n50p6icejiIdu
BNwZkj3m4xeuKu4tTVF8Kr2ycWUm1SFQwrVbSgxpKYDyKxSVSfr/xaskNxK4kheR
0cQKVIoSBrmIc5h7xpKMIPB8rkWND1Vr23Lv4zGZNwG2ZPdqyBfnYgnKCLoNm8rJ
p7oZTwjidjHg+Kmon/3RQ9f26B95Mvs2EZwkwrWUQ1EBKHHnbAP592FvemPIY9UD
4J2J3tQ8vR69PrtCeHxprfz8k2uJPDwZHReLpDteFEKVdhVonRMDDhpC5KjM2l+0
zZnW0beKGqqbNEuSDSVPQlPGmgYFfDP3raXeo+jfHHxdY6conz22n2/MNHlyn9+O
NrvcbeaJT5I6+nyaGea8WNUgo6DKC6RDeB9CocJh9Or103au5F9flqI9+eAS+d8I
v1OM2f3o2yxadU+oqLgg6RuiGZbARY6Sqf7N+Alc7jbhEEcjinD6sCoiPnpihlr/
GtMJAtSlbTQ8YWc1UGOWMHPnQ5koJdhVzeNXoAe51SQ2UaFhJb3iIBhxXuXogQKc
sQWvXzk97tSBwiTD1EGxMgkBzY7LRsm8mxuzDZwlODRP3KyT3KT+AIqpjpgeveyt
2rbsKSyaM3cj6bENLRqCtpTofOZylalmWvyM2yopyZW5fpzZQ+aWGiWteqxubevy
wu7BrNgAxnWGZs6rosFo/xrB4fQe3IRPLHWQJ5tCLi+y1P6TciQWtM9au6tLvLTq
rDiqwUtCevcssNjfuwWtLq5k8VmpNYvXDTaI46oqP6+nUcB+9NYwm2T8ge2Ax8rF
rGY8TzqtgpqvMpcn2BCDlYsGWy/cZMm0eSi5A/q2HqXA+yiZvr/l3FZMPqYkNP+S
jD/ms0aNGG1qpZrpyzTTEsZ34LynkEXtZBDvFKdOFMzYGuxtTXJWr27T9m4KLdCF
10zRa6sq7WW7FBSWeeoKEilwKv0ZAfUxFhdP7nL/dmosyQsM4/msqM2EhcwGJgKC
xjB+3mJH9OdPvFuDUkVgDZTj3Lgq5xx5rfanzv8OozagNdybLYrOeHodeY2Y0aUV
jzFW1ERv8lUgpd19uORISfHMAgMw2Nm3kqPfU6/WIbPXsv6G/tvR1CwZGusaDE1Q
/uLCojpqN4A3jdQj531Y1yfe5IlVojhJ/Vk+3z+ve6sV/H4hweF6xY7auFAYvvJx
mZSdVDj/m3ZuuhO5KTkEEkbv+PPe5tY+s5jFosW8hGNj/ee4Ge8VWs7GfrHV7qHJ
7L1QjLlb9JbWYV9bhfdS/Q2GgY9WQxs2lPKESSVUnbCxo4KovvjfminYRjrhHkY5
hskNAcgENM7GOnpk/htIdQwInk8NtXXAHCsu/vfMtuNf1AhZ+X2dIwbE4WlNvRg9
mWMgDB1Srypg//QvdNen92LX/qvvfRa7ba1iWXSEbxrimBhwokScVrRM+DJ9rRw6
7NfIevRtDXZBh+8au568EDTzpPIdvvhX1CXFAVfCMGZMpPeArB8PcENpUt7/30WC
NqZWBtegzsiDV4yPbWq2bDaeCMrC3YviDR8mrJkQAduYpOXrx8hh2plm6m5/PvAe
QA7gsR8mKKdFGqsOaAOk7EWk//5IAAPgjlsTwuCwo5SKb06YUbriiS5C93TJEgCF
KmP9XNsYxRU/Y5ib31jrH25uHAo+9W4PyN+2ZbP0lpCUB5tkBxgq0OqjoURoZNXm
JQzxR5Cw/Y5AXCjuyDLIOeEeslmaeCDpTsDXNf84GUzJQKVortWBrgKAbwU2RiEQ
EKEnP/TsDxIP7RPEaaxAzWieFKM8+x0gKTbGo5PmW7y7Tgv081iiPg+ej99CIJuo
wHmZDALtURfp8QQD3/ZWBoDDrhgNIPAKjHITTMLd3qnjXs5nC2g3APAmjF75SnVU
WjVlXNICOZCLomd2b/OUEsU+MVlbgTUenu4thBFHEOtPbp21RlP2miz4hVY9Lz8x
8RepJ6wHzmRH6ejj5WkYCV6z+gvZ6turnk3MRSuy2QLf7MA3SGSw+0prKC8rhLzE
wOd8ywH7R0JqYfROag9HLI8Uc2N+AxklrpzKLf9Phy85smdshuUyTUcnJ8FqKYzj
iDkkD4K81sAQA7QqyN/AZ4BdGc8GVNjNoZxwr3vLhFq62uALI3d47EVAnOOrex5Z
gq4qFmufXjfwH0h1ZiOnOp8d0NKzw/sAEqtkZ7kNvdhSYN+J2W2ty+EcMw9oDmwc
kzTq/NU8dUx8uqv2XzOBnXGKFXbyiF5IzjBo9ZRmKS3uOd3/+WVCvZIiaydiUM3u
SWT2ATLqLnY8VYtgZf5sJDlRP6X4ezER+6dRQhqTbjS/hb60H6fgs1gqtZUHAAhp
7P8pufswSiTUCAixFlE4kL2vyK2l9slL/WXlP9RMGUdZUuMh25LeUd1XK9r0R18A
CSeonD3alZCm5/g4QTONNx2liSfVPkhyYHyZAWR8jEwdTwu591u6FlvXtQpS6e5e
R7zrZJuN4nj6kotw5d5R0V1SXBC+oc3zUGLwPhFJ+suoHK0dtSQjqYwAhrgVxrSS
qLLkxmRxvpoiZR2BBTIz/WGtNbrFry7E3YtlkpqNSODw1Ikx2/pD1yvEoS27Bgul
mjQWpJD2FxKh/JMhCmXcPfY5G06KojBXgNy9FftqzvxXCo7FZh5ElCLmLJ74iais
5glqGHZcWqP2OhtnddeCzOveQBGPSDOB3Y6MmdW3vK0KCZ8PROUWUCaK0RgDloAv
1yG2Vi8WLGwhipds/DpUzFwzaIqzhycR91eHgZnVzHlgyUdII2NiLYGux82LVUwI
etbbEpTZnVrqDIBCKSEF7jSK/b4fF3Nb1YNLyvipFa5GNDaYJhSMCVT2PLBjY3ed
zyc9EreGhM58Nvw1oaGtwFMHbOZVDzSsPmhIX/JVfl6sTkLh3ziQU8XUq5/WTfjC
l2iVGd0ErYXpIqx3ask4i9yUsDQwUn35IlmTe3sfQTEmabADkk5wkYPouUwZHOv5
mmzu1HglXueRduE+8ocUeWRZQQT34L0TBMbIre0BGwBdQhccKXIyM9vzCZ7u0eo9
WCIbs9lMd441aAqA7ITPvp4BaOUcZy8KzSJZV7mDZsWZVf1s7cveuw/mWjWGY/Pv
eklZMRGC+zAVLYmftCPhYNgbL12bbuup7ts0UEgEqI3vzo/CZPuYq1jC042J2wjh
krrL6x1rIihMEgAm321ju6bhayB7J29ckmo28PDRZaFa4C9nUtqKnpbLv9CjFUIr
3zR5tN38L0Xs4yR46KFz/cacf5qY7Pxp7ZBWMbxegKbWmtinTIv74T227T5TXlCD
fH1hLheWH1U/GVIepASfeLLnu4l5O2SSz6CsazaGLbuV3iEaoRydDHo+clESwxtF
9sNyBeMcN715cqbmvEy3DLFTT201NbhLiqzweysMg575arznp8fQTTlReqiV/F4s
UoU1urZvBD3A28X+V+z3ZC6Q6qXEb794UZZQatvsiubwoPnLQ64R1k4OWxzQnnpC
TQvckmd15tItNa04gDg0myNmXSg86arxvqKuMgZyZ7tSBUW5L2vXhCzNZJQGYDDG
WCZXwN0oOWaLroIzVcaQd11r9QpfynmIscKhxtBdXk/zUTlyfliVCw/xnUjKO3zM
8iNQgbTB2DQhMDNKSiMV/J3rZTnii0Da8TT3MUhNjVXyrVx8XOZ+z/xbMYqQhzT/
Q2Exevls2g1dPNhblP/tJfjOr3cVWNWB92xo4f7Rt6gGqcbQx8LFhU0Y/J69aNvQ
4wDGzAc/SunaSue27APOkWHLUtzBf91VDg6ve77jBhpHeKFITeL+ILoyZI4kDvlV
pK4ix1YcXClIToh8YpEtTNChZ4bkIE/MRGkcslA9MYfgTRqcfv1JZ1oo2kjtirbl
VReZoKiVh2JEtJabvh28P3c7JGvBqD0QwqkdoOCbSTEoQ3GhCoqHI6w8FPfNI4WE
7v4MV2JXniP9Q5A1JTCd6G8Lclu0olGwuxptZzE7hogj+MYfxldMKaaUE45Ov4t5
LnEeJ3ZVjcmwF9A0lfofgCdvc3P0OLhtulMiy3l0sY6x2ANqGo23zwkiePXYEHeg
NsehUV1JBaFUyAjXB2wvqZ/UZjXLgcMCxPIX3d5imFcjsR9mD1ojanbEstrp0Q6R
5YM8ttzT2FbUMqf+MCfDDFSZUsjitpH5QfAxbnWMKFnyhblwam7SJarUrKZ9YaOq
FYd5S/q/TRkIOIF69ED8C+UJ1m/Vrjpvmm2VzTWf/FC0OXB1UYlrkiNoopqSTXXh
53MygwsY5wrZ1JzhiYA3dahZo9HEU7KCdMwvwJOQwjyBJodGVj5aEl34DnWAVXQK
feADIqrfxSeV0qtcn/M0lfVqqktTBVJ4pHz1WrcoZvCBPZ6jm9IwQqRx2Xc9FRas
4fPpJJCoeD8qXxZoqfIk6TnAjYV6wDKkXhqO8I24O7x4IO3JyBKhksVq/XyPRN5/
CIeqPUwMLmGTgOd8sro1Go7YF/MjmSVAOfBnZlgxR1ka1QlZ6mMA67aA8qDuokP5
nLc9xfkdYOMwsv8Au97Yw6oUl4hBb1wdme5is+rIL8S6YIEM1xQ0CzQ/7P4QESKU
xKR7KWgeKaBr8gkgcWQXVziJ9i/kOd0xg167/WtERMbMB+sPgiqtMPmpfT+Ai7Sh
C1P38i2CLQvbaoKN05Y7FEjhKx0wkaUb4+ZOQp9KKwZNaZxLivISujEYgAND9TGR
SU426DQOifvgYgwztgLsSArAOc36VZAH/kvcnEPpukwtuOBSFaN7cAswPXUlnv9D
xGY3PaKnUzaNWDkWrd1JzJGVqftnzJmSVrP3vA2830lyYv5hQwe8Kje8/z4wA9ES
9QzQucfZ57OUSC20sx8mLM4/CTvMC5fviDQ1bQJY4vI2ULbXVkNzzNTGQLemo1vB
UFv0aOUhooRWNDKbYhSJYQOx1nxtjdpZdz9bYQ06+gTVY1YUiSsQiDPC1ZDvQXlJ
ozMI7uZxJ7OgxTPYeBIGeQG+kYqppU0i+dV0aF0agIkYDcp1qdqtV4r7nDTA1VgX
gJM5r8OcMrdKT9HH2ekSexUIUMjRlyHsuSXhRw0gmjXIEU75JE5QFp4tppPYVbDL
UaeH59pLFyCDUnltThonop0wc47MIskCbF2tOq/B9ZuaRJXYsggYOlV/bwKuNQ9i
GVcAr/wbHiXk3gNKhYrHaWm1fOPbspQEP0+RdILTsbUzmSdfcK92ELrNMnKCHINX
ot5lGmRE3wqTpGbFu+6vZmRtuRgcBcwuJw7mY37j0ya/iuOBp/shid4nKJmTzDcM
UdgEvHOo0AxaxibN+v5TKgRV54Ulv2aB9vo6nzGzeL2pYRHF5baCtQd0CcF6cpGf
egjU0Yet7z4CrY8gboa0C5chLXHqLDE93Zy190hNlzHH84MXSTrXM1kKgO0kWwFZ
z7oJS5hIJ/nBKIvsqc06AJrD2shGCLMCkqpstU82pr/GWYfiYdUphQNGoRjCiu8o
6NFkh/nbUwLR/fYei5AshwCqu+XlufrQBhaU3TjOgAUIO4wazX7NukCOIqw2nhZW
ym0f91M/39El6YLb1PW6kQKiIDdJSvTjx7pdFwNazN5daMxa4UUWHNQorGrHt8qg
t8ZRnCx8EPVckEVtMDun5ACCGhzjm2FqXzNDW59+2L77zpSqtlfnwjDIJ/LEcOIV
z0+5kEKpgi0wciYtzqRML6zj9c2rFP94edFg3b2J2068iXZR7SgFZdkNYypkvtQL
8l52HUu+w04ZOWVxDb1NahotUG6UZFNl7uSfbrtubq2VQqvhTr1p38x+AybPSCaK
rqlvmqPaJnsRRoIom5Hjom3WbhI5HYWU/jGSq66GuuggjMiNmIjcchmWF9RnSWvi
KxnKrgqvZH88g+jVqaOoEo8xRkU3XMuSgQmHOJL9mhcu+UcfSOGN4IHU/eESJXOm
hKSZ7lWz53NfdtvtWUO4gPRsIOoMeOO8xEOxrACw6KKGt1mcT+lPfPfiwVkwFyJ5
WDPkkw2h6j58hRTs+AyvN7Og5BNH7BTaTwnhjMd8uuXMDUz/KWU1diXHHM/VqgLl
7ingfdKFjilbBq7WwDLbrTUu5yNq3c3Xx1BggCq9YBOrsGgTq69mF1pVlqb+UhP0
I0VwPb/8yKNFHNBG2JhXSEWcPQS4g8HQS6PUzO7z3fwSJkdjHJ1epHstHm8R0757
ZtEYNFJGlk5QsugBjeAAl0J1QH6jRpmJNYdpxb9xErg2Cu3c3xekmZF1Z/zElws+
IQPZhMqHZxzEqhyTZNhuMG3XT0sT2Y13pMW/PYoDWO3omzAykGPtecBWC7Jrn5x8
spgIEP3B0TloYkqHAmV4E+tnwQv7vcX9NP8Vbp3rnZVTXSOfw3t6/nTxJXbO9FXI
Jrb3x9j98e4pgRQBrgXrKqbwdXkostVSPv0iDvg5wQa18lQSo6SH4fvBHzVHiyya
mYScPrjMLOLx0r6gbR+swUiZGJIHDTkc97iFKwrJ3lqk+TNJPrXSYfyGOeHX/kPe
6lhtP3SAdqmW1nOzHktTwxVe3DEnOFhSMCj/2+ArssBqa8BjK8hdTl4LA1CXF7Qw
eruGoi6XjprH/cv31mYjaGfbzZmE9ASOaDpSTxE3b79+9jDQZMqARQax3mbGBoNq
K80OIZjLmlAhOJLge4Ab9qJ5XnUTsNxHAAnEIea+xf4q5ADQ6GcuC1vfmzpSzz2B
d4484efeuQQ9ifQkqYzuxtgVSVbCby0eDUQ61fSYyIIexNdCMZsXEKxMIryT5ERM
lShDNp/QN8UAZXp2S0F9k8V2ryQc3Am4eXQYkALTYfIQbPF+LAuIhn9TwUu3znCo
LB4xSq6lNzc0BUzcEpRO0ZaQEwOmqJZkxK7fLr96xTAk3f2/ee/WcwsvB0djyWCQ
TRTrKHxOEaWZzHZO0QOz904H6CN1e4k+/53WPT+Mh46DHhW26OHlEyQ0DV0c3E34
tX5lVsmeNlnl01aIxmgbEBEp0bWivMOzI3sqOYqryjX18dYh9eulozmiu8coX1+g
z9Y2PGgRBYzc2162Ji3cInLhbiWwzIzvJTKXWDI+m+JY6frXVEMDKbKKFRmg5fdt
G2lFJkpdTrhU8vrvmSMHsUPwZEsn/kjMwIMEB4mW0CnwKyKUoapbwcvwB/ADIMfQ
gCMnrnCxhuaEsDPO6VI286er3QkE8hEmzLuZcDqh39wRzsRF7unHWJCSpRWbbeY2
B8CHTWkHwsSD73NeY/qeQ/TzGJFK39bMyMS0uwI+aCssL4Cl/mpofwPMiUPSmYQJ
TOR8VH/Qw1Ti1uT2BFpMJjKVTRBVh8Rnpv72Xqu49HHrnk47ih3cKJD6lqTdYZp2
PnlwhYd9jJ6abvpPkJTRs74tYpi24qMaC8gxW7L7PKaKHfncqbb9zw93prgNLtgM
Ll3nR28VZt4qMZ5L2q+nRqX1tj/wxneEgcvTON1JTUMLhOGDUBuHxIHSGZ9/fXRv
BJUS5PuLRvDiPmWJ8KWu5pMulCctGRLAfDf36afbk13876Qi8aTmUyDHwgaQUFUm
Q3g6ZEa0MHSw0bPMiXMGSyHH5a5JHOi4qW9FTr/dBTkfuTioF4m4bNqSVU0UKqUq
f4Mj5q+UxVwuUYVRVpGT91uSZ8ai/0Wrb557qxvkrkW0eDGYHpWkocyJAAj8Q1kB
TK68oU9sU9Jcs29d0g3PNZ/LCMEmCkRfx1Cyvds+Uhm7Qsk7OOkb2UVEM09o87W1
Ru/yc5vY8nKrCoLMhENGZ7ExP3CFYNK+oqFSuQX9SUkzPWn8/bTbqKZJ5cEosj+p
vra8U/aBsnDSmiwbVzE7emNyUXpQE4gnAFBXDkc0scq1nQ206KtMkDwtN89UqwGL
4DGAnVF1Za1ArbVkwOSjyrwSqGu7ogITU6r4JIBhciQlZiwlFQWnnPB3kTeLLzkZ
1mR77kPkaNooAWD8jXU+LwRxQ87zms6DJ4e2pg9qlY3rMnXCYlf6HNfUBt1jgkeY
ou5h/6V90SvaLf2bviAYAnEVS87aP73wwtQR4GPXRJ6WK7gB8JorkaQ/q8HplJK6
OTE9z2WP5pXkW7ary1/sG4WxprEWQONExJLPjZuh3SpnGzFUOXNoFWzrBvFcPDjY
+jRcD4sxhrtJGNQ9fl+4gUvpkeWM3V6Bb5N/e+0Ydyjw+AVJ1zZ9SwMN8Y7iY2XH
Cbmu3enVZJ0p6T9WZB/uxqcVib3yf7sani6sdALWHtJmVQL9f/n11UQD/6oG3sux
CWfrSrhEKIHIXWC8uSZha6Z+aqEWP/ZGove2FByBxRkRjjDmRj6Cypd6uzg4A3/r
2hZM3mcfr+9ImBpzQYQ+cAauyrxzdSXBZH8Xl4vWar01oMsO9N0yn7ICb+A/f5/Y
7CrESZelw6vvm5I3tvXukwv9Lt4hgjh2IDtljZVQUtcw6r9iQs/C3gw7JN1KChMP
tfydvr/3SUmkoQ+d2KHB9nIF5vHryzc4Iid7jPbJpR7VzrqKGNaEsbY9IZft2FiK
u2hM9MOxWiWikZfx0PXg+kwzKDv+YOGKf9kqM2QE5oT/W0rFBI02pWlu3X0J3z1X
KO+DdedcfQCEE0roZyrkaysVX646P4o9NE+73s/4xlGFhfpDH11guSU7VbGuNHTz
7vOEozmILJwIFs70s5AD4oaxA6wkcLJNLybLH098UPzgCjxMEkgEJ15OCAH91uV4
xXs7zJhETU4bqE5qM6X4iMpixB2S4M4PBQfcxRkEH/pdyclmmUY3GHLBXJWVC18V
woZU+BvFnqoNNXPSgKmWTgJBiJfkZyswmx2dGBEhlP/ldlgRMZc+7tpnJYLoxh8B
c5igOxKWijU6CRf79zSA+aQ8hc/mbxDdImGB02w5/5FUFK+aqbQERHWzzUo4mD3n
mfWSGue4D0EC+i20kzbILvD+7y6KDtyTDigOSpKP3vTbbxRd01FMtRn+atW0JzrC
xzIaRA2NqhzEXTJHr/Abz6Pevz131ubese7hc5Ux8ScAK8da6v5oeRysr9QMV3kf
sK2wtYuU1bR6emFCroJufSEERpNZk4Ysz1wuFgHDDxkejYZO3PpTwwIpCbez1yG0
6cyWdRg4zo4FhWENlNe4vsmyBb496TNcb5Bc9zZ7rSi7F6dI6IIPtC2ed3nJ3PlI
2BRsX7Ro8bv4mYoC1igLc7xSmclZBSSS4x9j/KJ7oykzzOHU0lkDwyq61jKh53PJ
cbQasK1W0oEZF6L8fbSmt9huCCDs2MWWbna2+4tre493m+1cSXjP1Gj35Mi1mVEK
pprleR74zjY4TCuE27e+kOfoOHExhBeDqQtLYhYuUv8A0kaeV+N4OWMGyIojz1j8
jMNujkV96p8TZbrIIUBdlXe/jdoI8B0TD3vCq5fiijObeIyhMXejl7uWqhePGkYs
kzymg6LGY1nb0inAnT2bk7yKjB1TKcRgeUfmlRVP0kHkbgWfUF3TpE2MFzUVX3Ix
NWhZRZHrYForIEScFYTm5Sc/4S84uy+A2SsN9vT2nFbNFNozEdmmyT0X8k9Ez/z3
Xa0rfzMBLjH+lEC/n1p/zOxApd1QVBCE+orF8BIlQCwTYqhjEa0CdZ5wuwU+AaA7
JmHX0DCCRtYNZB20juPJzdXH7leI3+rvmdCsT4koUh12qPVBCapM+LN+ZvHR7/3p
AZ9v6QO9EteCJj8euEhMecK7t11Iv28q0g2Yu6U9LjdffP/kRYjPM5Sa8h/Sp60I
mA/ei83O2ppIRorR1q0+kwnJVFWk9SY4TIDKbD94exwYoWb8Uty0hABSCYGKHQXH
jfeDrxpoo9rxJa7s8dix+kvAExREjhVG/Pn1nniS0JrIDY6tEuEJYZdw/0ojIcKO
NbgyBvFkszSIjIytxFSmzdVZEHFEeqR/nc6aL9zvOaO3bzuihWGkt90j2VE706xs
Ll7NltrffzwxvHuiEsKIEK+jJmVYrkRY2azoBCjL5OrFLqCBbgrh1Ign6q0jrile
nP1K0LGbq6fPvVDqwvzW9eYMojujCSPZM8ZtraA05DQNG5fhaIeYr8JR5GEGvjI9
5sIiYpUcXs3KNbbHFiUfqu5JMklFAib3ITAxyuC7tMFopuvn/c+fLnI9bwevcK4I
O0kRC3eVx/ikEAsccexlaG1Z9wBZLYPO6Us/hRPlOgrb9yYFQLsy+QQ7Kx1B2189
NHxXTj11ij+sfm9UEJrSn9InIK57PmQU7li668DknrSLA8ElRbwkbjclGQsxEnmq
IiZjKCTLFRuMsZ8gavi35RAep4w6rtPWvjHYmqUgewmTU9mrI1Ei4SYY0q/SRqAX
3yPfCF65jmljGNQcWq5cFvIzhwX2p/AG/smQt1ifMVP4onM5090T21sVsuSZc6aa
TUW7ddxVo9oLJhf8ab1I2vsiSb4k+tZbwi7TBtJsvbi9OCFgDzNxBoxFwakoF9CH
jFJO1TmFyX6y6WfimX0LDsxtOktQeJASAOqCUhJYuExd4WcT362sXR8fcfqtkfDz
+mc3nIqwkQhZLMaxHJGp7sXrlBhzOXBnTz6NzFsMkxZ94284qmS3S5BkMLZ0Ftha
gMUBudB4isn7+8zo/RuckguKrbBcc1fXG/0U81S6/+LeP2OVejkIhfbYbF9jLL0K
7M4N7jngeLnXqJKkwe2z2vGSaj1Q0a/ZFjiV0r/0eCoG2TH1pjxIUkuNZBNVQlIH
8D7UakjQE88/0tGFKn341R9r/meoU37zSZ4YV8ayh8cNtR13aqOibUGehvqAuc75
xDjfIjgPXPnqEYYMfwfJcuy1rXzmpvQYLMdb+M4yCwbFYOq6QDhgL2JW0SstzPLM
d6ROvlfkbWKtBmxA8ieCdUNPuLsAQVPeNkivjzLepVnE1eIhP/83Sz5PuQ52coWe
8ZUXBtJorCBp1/gZouKo/670uUd53p43wrNXNoVGDY2SosKwe3/lafEhPBUqbDxa
ZzRqOSwyPCWLY8GKC9SfJLgfJSwLoL79fxQ9TqH8N/gXNJfTrPGnhCWUimfusYFx
IGByJtvhvYzOsdYVw4UTOJCRcERhLPTP7AvIY2iN1kkCyEVl/IdwA5Tu1MwG5jDY
MkhOwu9IKOpNnJzxv0q2hSemRvAf4hC1RuEKqtifEEIkaDx+KZEPmBbXw12nRmrF
31cUQ6aioEvSCMVPlQkmXWSr8xfGzVRkKH313oHYmRcrJNTi1xOKso+kQqofQDpU
DQ5QateGovIS/Hion/oKIyPAmkoRsh0HRh7pAAyPyQfYk8KIFupBN989L9m2DtZ1
qWjKP1QQnnRYYTsH88rT5cUxHiOcthy5s5RFwAjEgqLabQT27tNfVLKH2GG3rHX4
yU3cQpBxxsKPKpR81BLCPDlO7xJViXTocyKg5YyspTpcEiuPuy+d6aIvrlPWq+j0
271BOgH3RUMPr72HkBXlKmb2bzO7DEybsV6ytCoff4mj5lJM4pz8hrOpGPMLmP2o
LEfu7FU7UOD7Sn2ydtddYDfxgKmlIKt7WEEMUjCN33nc12fxlEGKD1xWD8Ot3blQ
uUmHwKuxuRctVsFaGGIHIiAwoB8FQdB1A8cf7JwCKvFCdCj8OTLv/VMlD+WyOm4/
ZsgLahKnrNtBnjrizWxkSDIIf39g2u7ppCCcnc3TJ13ZTLAa34ZPKDJGGgXuELNE
D0l/HdffqKEZIMXOeu4r7YW6IO/PZhl/hl2nbIPPY/3WVzEMTXL3g81g/o1T4Yj6
QcLJrKbyYmhC6dAXmaivOdfSpnUduUWbfS6dAZZIJ+5Syx7w2gqzVBTz1fJcVj18
toxtZ1JlM9oq+ttRfNMUSug1sUb5RZEY6Qp7cDqntmt6SqppzMcwkYLxMirsGU4V
DdaWNhtDJCb4v5InWJ1E58OUSU8eDXl81XzF+0xilw5x+6ch56bDR43JhsjhKNZf
dxyV5ljbjn8H29vYjlqTIT4tJVqzHs8KaBwiyMFU5CAgqfys73Jw6131/8QCgrQo
XHNHBUw6U6w4DgEjZRojDdSiqwtLZD0m2bHLB9osCRFMhr0h/1Bdd7QI0Loi1iy1
7cgirqqZvk7l81O45zxIfq56G3TsyHfSCAbXhktiZOqnNB+el7pKDLzx6dMEtTII
+OHo9W2yuCKNVH8PpgrrIrbtHJu6LUAIBCCopi2Gm+tOIsGmDA7ATOjtweeY2RNP
CY7fIuJYbfxeX3tqGVXkGYgJEON8QyddacHLmgKu5E4WePFvBL78J6m9uPtJQ3iX
Tn9k8Tq6wJ+V30hPXISFT11gldLoEQtRZCEtVJ6Yyh0kjnoHXMTdzzqwpHU2yqmR
gpGt71uudpoUmA7K6NqAquXCQ0+UnWu28HeC3aMzyzf3P+c3bvmU36iRndlgzBX0
9DyF7/Ec/NbLWhMV6AP3aSn28oq0RYsT8mrYqNlGUHpA/vSD4X6jjR9X6Ms4d3ny
D9liUpr7i4H+iv4TnqHiKpvWGpQpUnKlltowy6MPtv/d4Mob+d4mibmnYjbPPmGS
e3xuEVuwFGY4ylMd93v6K33ptyhysaqgevhUd0PQwpLQJdakWBndDB1E6KYZ7xk7
Ru4Iw/+dPk7HcPMpdhhqd0SIk40UXo/kahh0fUKlo138Qsku8B2+dSgvUb22pGSf
11zH2dAi34f2sMiYDubqfvojjoRfsHpC+6gm7s8QSAdYblNM3Kz3+V2HfguWn/AE
hZxh0cZ+oP/k+pM0Cl52endv08lMUMKsTzGpxlo9k8ZgEXNe2GzKxFdOF96iMAWF
rFBeywyuae94Gd4APvPUrtjxARiyja3IwldvFf4FO+SpYgTblbp8R93RI79d+TXw
uDPyh3Umm55Xe0dfmKomTpCl+W419m7XQYgqSeerBidCIrfVvdp5vmFR72s5lJsU
KJZVJC9TiSpX3qyOABQhfYnjVtygC74ODjyVa7ob5CYPmyS7u1wzgcSWO1+q9tIl
RNMWClVaY4qO5/v/+PKTor1i75NZQTWPJ6CuU/dKVlTjUky10XwLLo8BfkD468lS
gGo3aSqzBOj1LotL82yUqdOnDbL0sSfXgcVFXHywTJ/NJosyAjqU3j0lGkt0epgJ
xcrtrJasGRYjFF7XNfGAtmY2t4XS8K48/E8MwI1rkIJOxX5CGc8Z+qXdnmmudlf+
+TgPbtIhHBIu59znfZB+n51Xsw6l/mvn1g+G5fD6owdeGwQUc2HdYVxQY/y2ADKR
yVZZjVkU6klF6SwK0E2iz5fyyB4v53A8cwDouwoagHKjp+qTLxYlZaGngGgnArGV
/nwb6iRJDUSCNyQvz6/ggJIgplxIq5r6IcXf9mqHf1rrzupepRYdD7xwaFlMqE3v
A1SpJkkgVEU37NzdlUYBXAHdUgeS3FH3//0Id9P/GagGzknGatok00PoVD58iqXs
wCnRhlrmBxLuLUBJZ5TaAfoA5MuPwuwxCQWX8QC5PTn9zxXvIVm+IysqwKuC7JFq
Yg1bOE0FTR0iu9Aj5pbSC1nkhKOWW9+zuIDlCV6OJvB2ljZXIxMfyUqqjpeX++r/
wQifuXP3/NbtJsSU4lDo7npno1qKnSXN6D9aBogIvTTKdD78Z+Sxmj+FBhbW7sbA
FMfPT7XTLyX7MMylTCOpYeXFZjYe6RTOYM2kzoN6fzqBxgBFbEBLvIkSD+3q4LoH
FBbKqyHpg1OG8zx23R497GWmjxU+Gt2f1GTumlhjfwyEaqb68ELgAmCJAclQGVLw
icVr8w5JUYnNVRM5MFGzs2mcTDNMBOK1uwiuEQ2qwlGH6JvGcf06014fkjIvHRl8
9rG74IFEUgbvT7/vtfaEXTQNPWsxmOWucIFeFR4W1rR1xS8Y4vVqtIiBkAZFKSNH
qR+r6TKc4P9yRTwhx8ZwbENf3VmQhuxVuwT185AA4LA5xEhkPbn/i+zfVEvJy9sF
as/bMQomEert/AkSA+UxhZiOnXPsyZEb+VnOHHrreIDrddcagvKD9T8l8BVgjwUC
WwKPaHHryhJmhA1LRwklxtUjIMvmoIKjjgVT1JqsaZo+Moc/dR1uGcoBwZwQo2H7
Vz82QAbxTUH6sf27i7VC85YyC7POBqTNUuPR629kvqoyDfBJIg+UxCRIYGXRWHdF
g+tMZO7BE9BkY/wPhnqGcmF90pgNTl/Fy1w7qPZ3ooCNttLlEnYXZbWOg4ZddD0I
/uPzdaF6pTgl20JArr6Y+XMwSp/S4NCBqkldwFiWYjd1kakmO5SRsEJh3wc15aDm
Xvt22MnR8vjNphCZWemD2OopiFakn6Uy7T/dZ/r7eq/Xir8pt1j0YifqMrfpnV6s
ljhPzkQDFQKizK4jjXFtrP8qnflLo2wVusfc4ejxr97cXLmt/W9Mzr6qOvue34jR
xOdLtKf97WkB8KGqvPhPIJulZ6vR528zzgaZ71g928J7qjDa9gnCBnJoPQcf1Pfn
e5G0xlU1FBkMF9hc+r0R+4RqcyiRV9j7ZzAomgbSV9Ya3RzuJZvAhUetwUwXZnTK
XT8ABmcaVBRA6wXyvGjquKVaOeL/wDpgic66PG/vxTVGokj+joXeuGO0CJXDkQ4K
f8mGVYgHIN/eb2lDO2ylMaaHJumWs8Ehe0y3Kf59T4UE3bKOJ4s2vptbPQoCiX/P
UwDLb1IS2bgwRi+vl+/T6jvHhXdTpscO3jXPX34rvKqD8v7mNLnPFEDpgnGDb8rS
ZUHm5yzBKVZ4FtlRXnB5vvgSTcCP2wW+Z3D3goIr/ValYDnkxULjyesL0NTKvzHC
y7wyOqQrpRw7M+Pmv4H7O4KD/pIMp3wVmxd7iv4jJ5eadjYuT8dbaoDX3dmPPIHS
1voLXU95z6H2eeHQqvxxJA27lOT8BZwbDYR7s38RgDGFWe10Yj3BAg24DOzWD7GC
+6Bi9kQB0DulIewMHid0oIXZC3c7D4ZpkrnKy2KIZODxgBhmkBAOcDVCxC/u3asQ
gzufppWBWHhQ3hx72uIwQPQZm7JIFOBwZgNetI4jJoqsBqW7TG46EJjThXnL+jiA
Dco1gUk2Le8YoijfxrcGqy4aHYzg6AKKGeyZL1P4s3nAn1Laj5kFWTV/uzCHS7NM
RyY95J+VfN9a++QOMcPGQmugbuY4McCb9haVRQkBZ7mTbasVVDaWfLfzILoq15Um
821ltkxz1LL69c9SjbTA8Ds8EKEqYiw9Ce89+jZFGJmc+dn3Npd69NWFGTLUSeW4
gb//c0YLVsyivA4p4sohpzSpAGXz5aiDJ+nheZjA1a1t2FWraYKrY5MaGqASptYa
DZN6zxx4vbX8KKTX4+SPeNOeRsgyXA9CuW3U9nTGvOcHadnATvbmdngsoV0XT7+x
fq9oseByh5TKUC57GQuY7y40aqYW770/YpcwFnPD/M3euvTmYQ1qRwR3scEkoO62
31MsvwOlXM1uFpJKJh13HkcjqS5m7LWP57DeOAi0LMvG2Jh433qZ44Qc56Q5Wl8L
hXsWh8Pz8klWkVpLh3ZGw2sa4G2+XmigQDzDuywnL1RrqEyECrebMbs67otqIdE3
cq45IWqvct83eyUI8fz7edd6VUgDDozKg4MX/eNFPYMIPnRoPp2jl+VhZp4kHSMB
/BAOpfdFFYIhKr5/hm1FKwL/OK+TxqKZa90K5D6i29cXUqtcE9SKeDMaxYeYV7mq
3thf47fR6YCBw/HhI7t6EJOBbJXv4skK0gPWvXhsSAM6eZxYfuHvdXfAu3ED7iKi
/5biv4hX2722oGnw5+T3DsJ/HNFO2oxMez21bd+bJbPoPPHPcqVmp2G3qkYdIMr0
uPmMdnF88YkPFrU9dD3D89urw06apHO0MlU8q1dHUJRlthxiU/GM2P8TFSnF8BMK
A2cAP0K/czb6k8Kqgc7Aq8je5HQRfxC0VCwr559yev9XptM+dIUQ5J/EaqlSnpT8
8VG3ZU8zcLY8Lf6vX1px46ieC0m0BHIrPbGIK0Zg7qI1hmk6V1XKUrW9Jli9yaCY
PLNUmTWHBgQJjabJir/J7twO/9m4E4EaW8cVz9dVj7eO5S8srqvUiiWhNfxOt1cs
BY4MvNXJvuNwfY+yZElrnZlK06aLpg66mZFLehEz65zspaCfEIVS6ZItLGBabmaT
su8gpDrn5fe6z283Y1O+0wbvc0azidNRrgMSHb5hTYIYs81984umQVuoOJL94kK8
fP+etsGhHQG+SVESinCzO/wVjR910l7+QMaY0RqQ9oNFmoZOfluOwMOcFZkoAg2/
FWydIljJXiXukhQZg3bcjklatRMr/FU6FTZYqxXKSDRqwXwJ1+4GwE3/Tcur00Wb
gbw+QdD14Ta7qZGYfHGD99UBQsZnIDj5SKi1BLEK2T6HIZzQ9pmcvpu/sthOBHbO
9jF7ecKuj2/rzl/p3LhrumaTUG9dmbAvU6SjnVLgxglmgyHrGTYkSLpRfkoJ5jZp
5oN5UWtVsUqf8KyCfhjtDXpvo22mA1HFABKW2faXm6wbL70oGKLy+hR0n8iwurEU
Smv5knQhjrJsmAwiorhyFcRuczw8QgogTkWRCXViIlRXmeSyI61VHNSXXtDc8lva
3C3CvqDWx0lQl+vtSJroUl1qYc25ov/hR4WScvvc3yVmOSsLsPBR2efC43BfcnB7
D1bojIMmIEq47+D6U+1zISiYzErYlD3uZWcglQwkWdZyPKzJ6Ywh5FkTzC9wFCtK
4tsrUAoS7A3/bihvGKpLQJZ+e/F6apCzIIa/wIuhTY7T3ntkUk4kt1zG/kny2ydA
morUrtMWw7LxCEG4qR4SmKChQgadkcYcl7dKRnS7btXgfJ+8jVFsn2LjumiD4uHk
CzqRMJkm8skxWbQpaF2cJJ1NWllTRIwJwSs2/IZVAHTDkyrPafY55Lztz/4ymVvl
oAY+OclQNZNCpLl/WE1qxhnpm0WLaz7wvxZSKk9BwmFkmCAxguGk28+mk+Sm7rsS
SvmjMJ7CnI0xNVCuel+v93CtZNfkNZ9+Kgo3SjkCIA+V4ZXy9zwGPAdD3JGTs6el
heX/XSbQ3KgG075BxR1mgDRfWpleUIO8tD1zt0gtIBCJwWrOozbrCAEKJtrO27wh
FpMPw+acq4X8ofq8sY+N9OGOR5DnfgiQf3Yti3DeuO8fXQwnPsSg9W/IC9VP3KxZ
BZOxwyRV4SjccZZLKJT/YsvGQqvEMtk1naDkHW+tqSU1asjE5l+27disCb1Z58m2
4vjYlJ+/cetxDy57+RiBSk8ACMnAESPsLw+i12tCfMIs41KCY8nfk5U2Mo0nOiIc
A95/QRS988wXL4POvk0JIkUCY9YOcbbVL5TmOWaifDzl/Koj1irz11VhW1Y4Tr9G
6NWFxJnFHjNMixLnW7sQ+XiCDJCZw27dPpI0NXUa62imRuivX8q8SljcwmDWa4A8
3/x/Yr2TWDnQZVXhAerXxVRnlR5Q417RmSmRmmIF8Krretkr97DEluWU8sqZ7yen
Bw6JEI87sFV4HaPWjoMU0T8Qo1rmv83sSuYLSO4mTRJTEHjAtJsG9Se1rvKA1QCY
Gu2MuZ1rBGqih9D696QVY1QcBAxVzTTl05OuZvFy4BbBYhUAhnW4O4kb2/2wmQ8Z
sQU23TmMYY3T8zl3f+TH9w2ILjuxMz1oMTiVrpabT+SLzoxTs2IbcGNNyQ+yxvZg
PAqtS5sfkoW75Qp7LGk0Uc7u0PnYRSjvknMWoLwMHq4vEVQ3nRkWZ83RcoishxEt
a3ToUJ6dp5y1tw6w5n+4c+1gwJ+umCBswZXVaulsdz5MiGIZmdzHhJ6ziYzR9iEB
PawEv5C9s0rUSiODZxO0sruVelMVmTNhuxHFZxFkt42CmMI12htdgpxAmd04dqlL
j6VN4/Q+qdDBY3u30/k7gYIx0GXYp/oSc8gFfOB8oEHXj+3I9WVp8fhNhxjTtI04
P7SxskSthhcTvCJk3OsxFdKIjAVVzrJn90/N1yk27OKu/VEEIq82HDiztCdyP6cx
SgOROcypGfgvHGDAECj4fIuqU2+mT/ganJhVtpjGL82vda9TYUWw68HtycAVm+VO
VNLjid6esBNWmhNPl6D47yv+HszT6uTTbSixBNqZNpwodv7pb6wsVWgy6xQq8F34
Bk0axkyzhASFEBTMQ+pq4d1wMM3+XwdXLHxXo5jQWF3a+AXKWx6OgqwWqHENB1WH
kRrh3J5HOfLbJ2jaLvWZk10XxU3+twaRlQuMdwz53GdZHb1em37vLN9i8NJedvhf
DeG+bcc/qmIndmno2dohM2ujIpFOAssIyKWKotOZUMmSQQOlP6h2LIdiGkB4BBeg
zReMATqbufs2Q7TO2y7sCgFMrzwRGw5Mgtjw4vH3xAzhM0lq7oqRGDt0MM3AwNmq
4XXHbqt/5M1rgWhr3rHfa4Upugo+bGmJOkuL3ArdzBJewJzaBIpHSCV68znrlAg0
j8D5MDwcwlMYmrk4kZL2ZoAgfyA9DECbV9ZYucXFje6rZ/lDUXXI5yHophyuICXZ
AGgakT/UGWEuVFodqAeBuq7my1Jq0QvL4r0QDrXKb1eDHaAjuK9jbgnClirrwF7S
gVWYvUetqG3V3ixFdzWGbMUEPipDxLUhQT6LUdYXKDB5zT0SocpybeD+cxTdPPVw
5Vv3qosjCKyPiMWd3A4cHQeOTL4JAGoH1vyjAsLB2cpIlO2MsZv3FyD+Cqbyud04
EQj331wr6OHMxBfFUbgaXGKbv8VP170YlhPrqZb96cBIfor0+O/M65MBCL7cxwQV
iWcDL0RclxQnG7K2Xkfg/EdIGxQ0bJoSUjXgFxL967sJR8uMf06xFV+MNDub69Jr
P0R+/VYqHZvu4noWh6x+DKjQaustwEPgwb1YJLDF+ew1+qeCWub8K6OsmFxy8mtT
yLFEEXqeAK+IGvQXY4UYqTho1Hf7dOaJQxMSJr04oZL0TfpHlYvJfP8vEHzJGOPk
SNMBs7VcbuUdjH6UFihZcj4D/bzaBJiobx2Jyny6T9Gl8CtiVu2QXa0nml1aFSRb
t6oMvex9rNENCu4nrK+dTrtcUk+iQxAltYM7Qiox9R4vAevHV4+s6PlAKiTmGBeO
SAJe4hEODgKVvKOsOciYCHg+wOaY/G3eE8QLRliwtkyqsrZZAbAffpoYFAHo8owh
ZIlqi2UkO3qjFozPnELTOAz4G3IJoZWML8SNVgpczBEASM0tKUZHcbSZjjc9N9HA
6k0f9gXCK5lrSPum2XhqhRTK/M9NnnWi1ACO0888LalrKcakgxeDlKhWSLzFzSui
J6oZI5nl9mG3sbDlk0eXwC1WW7NbjVES77hPYEf/DKdgLGDUGq9e25f10saOEhu7
Y3poxfc/HamwnxZ9ALYowpJk2k0akNJHtQmH5ftKZVJ12OeDO4Vhs+wqvdKVZyXe
gat3H7kgz04HPz9DzbNJvw+Omr7UhWHgsHjBiQD3O3KencSZoxaz7yotYCcRcP3k
lGm9gnymxQpA9NHvWNM0uK12M7oAt6FVwoPNDvTgpBUbY1J9MJVETiv3g3IiI11d
hmC3HX4LoA7LfHM/LNIN3OkhXbnun/vu34dy51Bvyi5hdOYjy+LyLbB4QNGiU1vR
wXQOUH8nhHu2sREDNIvc3y7drDxQF7R47v3Ggx+o3yWpPcYWVErfsBKdbLLSQKnB
PO52vby4d1gGOshSQUK26XaHQUxJIFPSK8L9S1bRQdmOWzCaAI1zgz+SbcaPv30W
wDJ8XAaRwpw6H9+D2AABhpEKOzx5PM0nN4/z4ZN4j9+HpV0bF+noNjnddTPnSrli
8aEKlAZIJgCf+0Bc3mT8TOajOkGcTI+6AYeCZFMZEmh/mywQOefuzwTTFyaHn9Wf
CjFQDBXjxv1IxJkYT2pNdsoN7eomz/ZhHbF6uSXQ/mAPRLYDcR4+8gdsJ/QJfQ6z
wN1byolQfSb9Q93AZGoeob+apoC0fZOdSOBjPz0CqKGGvF2NTlPiFZJTee/WplXg
0h+ljyai7EXvcJqHKMrTFGIHnAaawtRAZajnXprdnxEB4AeaX54wsH4+n9FbUsn5
3oIGzpcCkUfYMuvH2kibH/4ToJv06q4HS7T0JpXBhBHuj5ccBIUP+qYhGlEAGSj5
k4Yl80kq/y3nJDPynYlNQZDv1j65g7jBAEwhVtb6r7+XCgmptmVGj9UX/LmfjlTT
K+djdQxQaseoyyEdwk9O11Q0SiK8L2TgGkEdVKkoCqslkx88YM7sZy3TqMV5BB9w
BwwRLF05Xilf6qMYaciM8UQbX4HHYxtVomebXEKsKgEgL1+5GMBWB0/7vcuf3K+g
SO/vJkpKsoG1MT+hsVhAR8S28/8GzKpd7yJUhoPT5YgFj87wM9aE/3TEDmKCuQoE
QGOnpWLIrEKcLtsU0hDX6UJLdNledM+B4YsG2z3L0ByaSx9zAIfDaDZIkZ1LKZmM
oI8YwANdJ42bxJO1qVm1GaSDtlTjXDS63O+Wn08vTFWe7yRdxn7PCcmSaPiUOMb1
YPY+4m/lUEigMgJcZIqs8yQh70SUZs7FnAbWRquW9NLEHqwFKZU9PzIzbvPaI0I/
PP7wFBf3kudbRAW1Ss4LiNp2//zjSX2o7ZBIpBK2T2NCqwyYOjqvyBuhhASpYUhX
CN6A6aUL4zIMy8FS8Zv4LicRRU4KZCWYJNFa38tNoEpg/RYnSwx6upgsQ3SDvS0l
x1e42nbN2Knt7JSO0/JXAhTCrbnSKqINIPRVEZprbH4gcZsvyOOFRwxKgWdi2/Wb
/oD3/DzulD5vfgiRt8YtLu97Ft2RhqJ2biSIg0aQPfjCU0tshBgGOAwuyMG+somA
UY9JvdAi8nTVz1neWF3vgsoBs6XuTWwKOTolf/H1oTyZewGVq6pYweHlEAZoAr6d
gx/pGQRRacMtJxsFxFVcY3jTkKBRwwryY25UdEqng8FKce9xi9WMUXx619o07E/3
DjrmyOv0recWRB6QBoubzgAbKh6c5DehZ93rr00RZliz7bg5njDSXhN+8Ythv4Is
yVvV+iiJJSa/NhppKjyzo7EDXDys1wu1JvTZ+0jbxoiI2eGAmE9ZGyync8P4BXx/
9yLhy3qPIhUezSmM6hLKs6IIRSOsg2SWHaNFvM4wZeTScUfXlmy8jHNNGOYyJkFA
Hu/5vW9mxnzUSYpSxqGHN8O6P0jStW/YrBrXLkO5kc1dhZ+z8rlcwaxF9ei6wc98
Im+phY7KW2K+WZBMl6dkswtYEMmKCf4pYH6a1aum5snUDdz9608AXCF/JFNGbM7F
YbSPtXs7xdAL/jNSY1mXNzUPEacJ5o2Z/vfTmFruN4lM88/2TSe1Z0udsdi4zqRz
c/d6CXD49TUL+tBYpESvxhuIaBWLofTOg4l4EL9OKTwGEc48w6UwoFbyennuatRm
y0imfq61msxOGUHoj/D9TqM5aWPrAafRIrtWxvzaX1KtZHwRNF97WNOl1F5OpC4e
TXyyc8Cdmu9UfLTiZoJxi2C3oxs9sK29dkhNdhpUMeDNKghoOrzkX346SjKetvYy
la8Yp4NGW0Ri0uavUrfLMrYmi6SlWpHbYDGCvPMSb78qJV8Bmor5P5SzViksMEiI
Sv4j44kuhcGHJYcFftxiUq/5Fc93rzNAj4s7LW1Mh9QVRK/vHq66oxnE4Y3DX3uZ
bBYxbXvwt+tgwSw/2NzrPycIp3O+OESdbFnk2j66evDOenrsc8ucyWb5CPIutrW5
chUuvCr38+1wwqN73cODZA4ZRFAbiDk1emkjlI8FgmVu7tAM7zMXgU8bV4+Yb09m
c5HJB5SNUOeTaNSE6dBFk+du9p/8RtqIuBZ+c+Q50uHHuG7a9vWIVm0Xj7G0sFXN
vG3WAYGasSjDv7dnkjLbpNeRaQ8KnHLmNEbNXYUsMVXE2pMN+PI3vKjPOdKlDZpd
cm6cDzHTHkQUTKP3vSWy72mK8wYIQuSPtD1JV+dyJ/6PHf4cyd7aY6kNuJ2uEHO7
upsGF57vOM2l6pr6POKph385mAKQ9YjVeN+yaOKkLqtDQEMvEBrgqsaoXyGWxaRL
6NESOOTCiYl2hHs4yAhNPjtrsknb+j4+CMJTeyrolMgC6TyzdnpciVxdOvsM2+66
MEH+Lu/K8sUYhiafMBrF2NP7SatERkL/pRMO4bk0FoQrwvr0+AC0B6LbmeoMOlyH
ohBR+z+WRwwL4v7iAM1cfB9rH3MCcCz+jLEv0rMsD1nofXj6Iat29Ae3q4zJu37z
QIkB4As8gjLA6j5YZy/tWZwSeXEEtW8sDH63e/qB4jnU8ghdom0ag7YV1CxVxe3M
x/8gRNLs+1WDmwH+LXdiXjU1H3ZyfSCIZ7YkSy/SPlb2n5OAEjZhmxBvvTWH/cyZ
aVkH+CuvoLYvFdY4n44RWHkZJP/fxaG94lcTWmSYVWrkALkspJkIkTqPV7HQSnzY
/EC2/u5HDQa/siLwgbCo19c3AxzYxmaeSPEOfH1ISH4dBtIk5aD8YjgDb8LYN3BO
ivPBFLaVDwehMFHck86MZOaems3FU4t4drVqG6ZnG41qP3kU2+nv6AQy+eLOMKqr
sNHc7evVqXE7FeJeUJ0bjqYIXq2Zz/qTlKjvPerSmFYc9ee1UHQYnPOqXxgZzjfr
RXJpJWRGxXIlyc68UNVucGeLQtNekUNBZrJ6eNybr0Yyhz9Xod7e+P6AKOPJIuqN
KZkQPw8dZxPwyNKIDq+Cm+wddbKUuI3BTlIvXpOosUmKQRUgUgyBzReq7lzRtq1F
XPmefiQ37HEXvL6kHq/BITV8qjqVqDlZ/cSNjoTrpgtC3aYkBxkk9fUtzz07wq4q
jhoTApIFefnl/X5DWc+Kcg4MEP0wO5neZ149MvY1IVo07ZXNRBF3V2LM1XPlK8BO
yIm916bhEGv8PVSxo/JdFrOHIvccST3VQ0SW4I469XFRNKkW5QI6lKVW9fd7P6vI
rh4cjZ/cpLXgo3NgrPfSykBGWP661+Za4BsGORcPtrTLPokO51GTucz+7NuSjJLU
xfrd9WGpYJzLV/4DppRCkmiWKcgoSOVgrZSJol2pDlEcfUAeS9yMlsyB6Af4t5oP
KbrB7xCeMMEQgaSE5tc+YiFxDtURSzEsIViZBgkYzqTfVfWt60Tye+cBPCPaCB4W
QjMaBaLhZr4tVCLdsNr+c1Vo67Fqosze91PiYIf1FCGVhxDkq500OK005GESe2+2
sX/voWiVWIIrPbUeKb1S7wd7odJBnbc4olKX5t2MS4Fjk98iEu0Y9AKK/G+2BWcN
dVhiTi0Du1GsbHvm5rwTdRhLpL05mdvVC3fsMRn3H54PhQxWlcex3/W5s87DHHEo
qAqiPkcQ79L819fi27hcb8r3xs7ghrQxCuRNrHjBbI/1MayJXC/mFmdpdr5cemIs
3MvvkGyKm5YkQAN0OOwY6qJGP0MScY7J4zdvQnYHmt7HifR1dcqVx5SNh3WUA7Xn
nQB61jdoi9ZRAbMq5aI+vRT0ORCXUEvbyHBYBgBTxORtiaSJwKGWpJzhQtnobszX
ZvtPZQ1+5KHOwYWb5nEG1Z5APX0N1h1jtfbC9K1VVR7H78dwN6J30tfePvalBLOA
yk+8ZQODtGQs+pzndMLpmqatIz2jE5Jlt/ZDbtFfXj66w3riSTpLt3I4u8YOK9fF
D6NqkSvH+6fx2GKcyq7YQEEM4ar3aCueTvzRAO40unY57GWQP/rn2Fm+SecQzPxO
HBGymrART1JJ+EmXfg19m9PjYzJCqNv+os4W8R5XYa5kiMSlnRuFbiEb6Sjqv+MK
sZWf6unE6gEjND1qBtC4XJ82QTESGxg6kEzkVYeh3XlhNxkoEHYbIOdrqiU2FkSA
Svx3tU+2IPRrtFUDxRWqSiAI2e/sWtFGed5Nk33Epv9S29sAlrPsexh4720h2Ue6
JKYWCJxLCrLbE6SMqmDyAY54wZE5p+RmNgK9JRM8JCLUJ+ry6te/FNlT2pcmQQTf
hSLgqPCevaaNmMutC0FRsnojBNNh06pbDPrcoxaLCBE9X2KLPM0VBKVOaQs9ZbHs
RAueT8MYm9vp5epNkzb2nXLyWF+Pr86QbGDOkaI8OqMUC+CViIRpdtwblU/ysQRg
HATa804YA55WgaJuPjitjnplD7e9QJifdWD5RySfbIju4E3zCEwM58yJTWaN5m+F
62iz2nkdu5xGj/hLzRgLXpkty4V02hBy1a+ph3Hu8YJ+YZMd9dipZoma8iIIXXmH
7QFLva2xtukc0/WiQg74OGSNwQDQCGqCgaFJHWhI5ZoDhW+nJT7Oe0VaZDkMHSwj
qPtpexCOSTiyfcxtx5dQCcviF+7zY++hS0lwZMOAyiPiQuCRpzp6GOzKy6k+A6SM
I/E0H8GgEDR/WtvWf9Bt9boBJKMDUmIS72uoEHj6lZhUVSXA3FD/F0QCSdR30UMK
06RREbC5+cw6LZvrjctfH6b899LJqCz5rE3odNc/5HVpVuoiAG7IzImN4Nc07/zk
1LwkYDY9eXUXaqxGYAhbk0o02ti+td8KNrH5L5RVYGsxird8UhXsaqp6aXsZIScj
tsPI/7J21IO5dsL8JxlBLSqUdpTOAvSHzenLOLOnI7pUUGjFJthDbWmzTYooXifp
dI4/kHn3vyxhq+4yBWkK8/vFmAMzqFI54Pe9yjlTCXst7gi3AxZxCmdkVkbYgVmb
Bgk2lDnyTW8zYphLMZcXraB/lRvxs9L5MBEHlv59xP0q+eK7TCVos49DBi7P5pi7
9q9O7cZWTq/b26cTp+vQYsvcjqx2JYLA+4FfhwbClRo8wuKagqKNMydme5W3tRx9
fZznIG2YRVrIw6SEMJVpNeWBF8JkGY6Le5vmyHGzIYveDJfXAjE86w2d02gUSHDV
aKSdK40pDD2n3wf7T3aZRhF4i6wbCYstXgSOFG3vseambNrUhI9Om9kc5WSQ9EoL
9AVc//DG2Rh250fhCyM/Mlxu4NaQgAiQIhUOTucxhri3vprrRkrSngshh2/XL6Y2
LTbKsFa28vB1wjjdQz9ji9C74GMNwAYor4AcoBlb1ls0OrXId65pd4hjSwQ99xNS
PzM1+YEOJboNJrRi6UAp36bohagyheO0N5h2AO2arVhrrcnNUruqDBvLxmvo8BgD
HuhX4rGJOdbtPKyEeh7+F+k4q7rv8YcdBfMH6UhyQ+avRjsZMGrWuWwrtfBTrKU6
R2D+QcusXAtbifFZXW5R1WVLUQeA72fcLSjVh10Nkx7EY/bPIdvt5I3hF0gzxt5r
0mk1gYSxnKhmUPoKX5OOW4XQGMiukOCYCMTxxtGqkbicBVH7bzgDC7B0yQabgyqC
pEXDq65ST9bPJHk4vZJhYqGJwzPY7PxNzNVSDG9VQGtXW+8IlqivfpoZ6lJZABMU
iXhlLWwcjR2Yy6jsemMuC7bqCXUwNAg+iJ4zCdcJbRm2MDwMycsbJGXGTHKJ9vw3
H4dx7yQlWKABlTzfOYF2Zv+OvZgFBbY7Yw7Doa2b3nDrfRnsPpI4gcKnDHljE2gz
736ff/K4RSgbjM2Ip6/tpYCyxY81rVu1LWw2ku6kiRwThydjTq6uKJoQna3VekEq
ayshndp3cEJX4ceEE/n/fAUjYzaHExIuN9tpjP6V7ngFSO6l/ZBE1r+7LTHSTU3e
ePmqhfYeUQ+vJgHY5KsKLggd17e94fPNItu8lOZn29K/w4BwphG5fqZ/1glBCFaE
qbYj5vYrIyeva7YfnJ9xz2um8mYvx8YsACWG56r9Q64+WKFeifq148U23+N+jDBY
iGGa+rc9tBz+b42Wv95zhOpW06C2b9BVilpFYE7g+Of41OUNSC1HYftPDGbetA2+
RzvGDwgaZgvMsK0I5LsgXbn6+le6a1UC7wklL161ncOuIoqU6JExtXixiY5b1781
pqgHOoZ+l9HxjuDnT7+0BKQqBq7j6ms/92KlfMT5BxYCnD2IlTOpv81WdY/vzYqy
jhDKVu7WlSfuNyonc2qS+T/zr4s5r5A7z9RfT6U2kq+1FyZBOV9FLQf4FruH+tpf
MJkKLEASUY4SsvNJkaSdUd9iHjgQDwEe3WCJqbbnj3re317XlAC4khZt3NMD4x6k
yrMzXKDiOSeQ5NOHNx7iI7GdV4KhAHfXUU5rRkHNdR3Df3Oi+6VVpp3nSd63LEkh
vUmfwQ61jH2Lh9TZ5IBhYCNerQC7eE9aGE/Au+1OQo1WutU3/bSfjDSCohPmvOYh
mjcPh8y3Kme8X2HRL+CQwocFNJv5ZoWyMsooY2dBrqQcda+LHBkqb6CPk+1MR84T
hsKy6bJzxMkAqE9jTArocSqgrex/Osg7oktDuFx3oJDAtApku5JwN9O0iK+LCGzd
ueursuvMiDOauH+dEGtzWv3riV3x6pDP2xrDEzdVkr/9gfv9mvgNfU2duCAr5Aut
nvLjG93pCGyak/8UcaL4HxudkzgMkLuURgUQy2WZUEyYNCZuokVdNK23BJ0Rnl5C
X2YANscs0t/s9giKjGb1C8gh2GBt202zc2WPMvwpwgXSk96UNfWfU+goTF5+rYzT
dpim2lrLosGZIvibUwxeKu9dpNTDmo4xhwRlz4luoCv3Z0YkPxSGnrVniIGzkU75
e+XRha2bdnYuZAcrtrMjvkS6KSkHozEK2DJ2WO55Dss/OthXYlpGU/NIUxZiWDxw
5C8tJ9nlN/LEwV4Me3HgMqilk5fG7yWkSQgkwWJXA2p8IMUNombdPrwkCa5pd6+n
MBstr5ALEns611mzg0aqa9rA+SbTenR8jg9PmjUuzePNzYZg+FvhWE7rANYsWfn6
qPh69GIS4+ewwO9arqcr70fCAwu1y4kl71W08rdnA6KiF9DhuzDmeN0KgUJvx5TW
XBqB0qMsM2Nnv45MpemO1ZUC8K1szw8tPsQCsJlPU3PaNTmOyElTbgHFv/MaaHq3
/jbclICyc64t3aL58MzvWS/qmCxvU0S9bPfLzrfOe4w4b+zZO/VN2cg5mLvUMRhz
aqb+6AyuCjPRFY/b6t1spkSlgHv/2FHHUmgjiT6XuLh+SQsSoWUdixi/PvXoY1WS
jiQcVdTcBDUFTHxiulF2NMKkCBWrTEWmRNoALRgQtXkE142DEuiSW62MG6V2Tgq2
vJkyxk7NY1P4tTOy4Zh/rSILXdV5G824x/cto2JXDifwaSYqCBn8tD0To0QOwfep
795HcTszpi+izilaNqBJKdp8/wlz3QR9fRzAB/08OtQqrs+ql0LMgXpl2VL+b/LV
LTawEJPB056AfuOIe/xR4HpZ9z00wcWOEeKcQNkspFAzYi30JxLeRzSgDDZ//aK/
niS2PNyzGBsnjjKmfBYC8MRqUjAHY0QPZoPbbW3kY4O5syCu35yHt9exHIGtXfx5
MCTT1ERLiNYMECa/4H8CCK2uK3j9er9InhElrSwNys0jpRYRSYnf8NSatWmvGLBJ
r6vhze3cmaWt/ZlQJAWN85WEcVgTfZGwDPgfmj2SuXbJLsIVESXDySEOqZGqdevo
TB6AQSuXslUASawXk5CCCMR3BsCHv1eWZIallXApJPxWw3UOP5+sL+Lyg5TuOJYx
YDiTOiYUCKuMuNmfwY0Cld3O1nSDPs4IM45aRJNxPKinfIP7J3IuiplY8Z3F96Ml
GJXLGlfiQz1CvDyC3F8hF6TilOPGCfpDAnE9DHe+yHD1TyqT06mm614FnCw4HzYa
3FXnGSQ0a84H8pIThynxcuzMaoOhqP0iBMNDbKn+LLuvUNbonruJzg/8eeTqDo55
ewzrSWA4U00lUdcPqlkbZi9Hk7kUrSRPnJW8kLp+HnQkAy/5NHTghlIp9KkvLcV6
ZUKf3LZbkp1lqd/r/5FiEC3wCefic1VWNZ2tKkTei5vGwiFBOz4kC4hbi5iXhToj
jMmA3tYfKTc+99OecrS/yFM800ZjL0fwi//WBtgz4pYNI/ZMQYm9Bnxa4i2Hb5pz
AB/b2KK8vHW4g7Ew79zF8IlLcvZHqtV8AjMyzu97fGI5dV0v4dMDfR20WMey4eh2
OZhGPc2jWi5cUL8y8tbxQ/52ezyE8JMz2zzT5xlU/g89FMI6DVX57mvvFuS3HpUx
g81EgNATRFnbzqpJBylfUcupmxa4Yiui3/y9GrTOCD3ssOCnJ+xpy7w30bgxU8EA
bHFkP+AoKQ3A4iCA3nCOhTeIYTe4o3+cnDGnLq9xu4fsVWoLViqCfSto9YXVaNzE
I+K13GcCJiPG3t1zsKJksv+ghsyb4RsL6BD4JZBLttF7DMrqjMA2OVoscbXW67B8
xHYP6Xh7MDDQqrTkc8+P3XoEoj+Wp7JjScwb4F8swNnzKKVNqLJYrAdNMCbvzsF6
4+cAjK7HC4ihFmmn7UMwtinmR+eM23NLehcj+iR0zUIOshgD6/G+PnK5rhLVNUHW
p9/OsaQBBgPqUg3T5tuDYFP8UV62jW2OvQCBiHb+++73GFjVUVRdNfIcSRsbuo2i
mUrdHyXC7FWORGoPVpNBjoefLn9Onqn1NkO1ZFYpdx9NC72MrDPjl4VSoaXxdFqq
bL5hZSYVtGTATNEBAhOzqe2D7yfacbpbZ2XGDb7hBQPQ8pnChdOylZc5lJ2N6o1g
7Bl4IP2GTMMcreRf9KPxoUGmYENindoSUPc5lhnptb6HB6vbb2Nqng36Y39gnICP
3OMYRFObUUODdYFTkQOgf8i1sThigPcisIZg0tXgfcdrC4wlvtjksE7kZdKxlqxm
u9mYEtJ1EY4X4KDLXBlDizNn8oUjS/kdlu1NV/7yxyJW1ZaegBgul/+3DQJ/K7bR
FvG/mI0wiCz2XrJsO66sVylLrBrTpSA8cxhxjJBZxbbVCJYWsaeoBKo5w11v53bU
eAXbsXfurdN+5QdEzfIyJyo8EM2Lmky+SJL1CRt15TsdFEPAnIX0qJDgo2jneEQ+
tqzO81Jv4vYKE/OtKQ78x+zcrssB2AJFNpozJ7XMjOKjjhKYZI9O9tq82jc61Kuf
9pOhBT0dqDCz8NwEZWb2ApYfeRkzeeFLk1TvladtVC1prphBUSqR1A8+NIfjFWMI
zSk3WnMejyqdlgCWyRoDMM12W1U8WKIhvnmXQhespg4q0Q4stH4V0UJynelZ7ei4
HwAYKtgq4yacSwNF/nUZSQEB0yPnLsCdq6JU71mA8y6i2gountY1oETUHN0HNCjA
cTBXgaZD+Ftm+V+RqdrUbnZhSmtOOqsSBGgjoK7yP/5GdsJ9TSgdGK/1bcEIxOoz
V3q8zeqSyPHH9cR1PDxD40y8qiFGUmulFlVWF9IYPk4g6FuuzKGMtK2d+LbdK5mH
oNpN2bPZf6YXr6+o9c4k1EvIyEkYmXHOWPKJDKE1kb72xBa81tUt54JQ+xGwt1pu
0nfDR9EoTCSV5cBZhf1ov8T/GA3UepsYMOv3ZzXH4J1AHqnhSsgRPQu3RDx1/ssN
ftNxvVaUHwqOKq8KZU7+zsnVnUn5UTnkMZP0rTtKc5pB9xaq9juT8cPz8rrAddfH
3wOQV2mqUvBNCkQ/eXy3I0y1a16J8JMh8FQ6AgcGTP7RSGvdKzIBv1bFOIpWu3bf
PNuuRhNaUE0goRk7iBx7G9kD1Rvc/0SAP8FpshBQ2q+hF9tgwIPoRNNqU2Z2wboW
EJUxV5pL0oUM6femQXFMQU5xH6GxM1skNhbP6PW6TeK3PkJhVacmTxDPnMJVlYPs
8sKuSy0mK9AejApJTcc8oyNQOPPjeFSTIYOPGum1rTtMsbsuJAMnezrDhntyffi1
2ZKSSA+YXSbV0eIlq5B1/d5Tig02QLM+PKfYU2mdGLfblBzTTiReYgr4+OaggDnp
ZIF2/jSDyShqQ+U9pbB9tGtThJjYw+NHND1rrcqETH4gAXcnVs7Tvb970GhlK0K0
A2Fti8VjLxc4U5MsDwTY4JBbiKxuOXVO+ZSwYhgDwqlYCpaQ+43OJlI6xp/uHx2R
bop3WFH7fvvq2RHw1OkAw8A2ZbcCUmEYxtP3ebTbPP1SrBtDuvrsdqeeFSObA4k5
g4A2vDrxCk1HAxROEZ7Rhc0HEWa02PHDvQk0IxrYpdWVMchnxk+fJ2JiibZCkD4a
K4lxtWc5eem4F4s1iC+3XAx6KmOBtwtedhgW5Mjb2U0R7Y0SwWinx9W33k9RrB+d
xahXPuv749mrSUs4zTZw5DEG8nwJC/QGB96yn1Bzxskiru/vtTtABz8yxRQWGh5F
HrhfeIWppm+CrBClKv4/6OkfUmDld5eVZnXM+pZJINcZtJ3fDvYCh+nhPYIvkjeE
w+0U6IL+AJ2u5RzuzsLzdrWwOeVyah2jPKQb2jNm68mB/sWXGHuCR1gD/XNegMzW
t2xq1K/7Ls3IoM+94EIIAHMqG6DgTq8jgSqCjUphyap0sCB1+AXY6OisQP2/621R
VWu7UgO7v+uCVbK8/2fARITaSPnAcGqMkY9JEvXYY/rQttIN9CMbp7apm3XFSRZl
4KJqN561bIore9Rb1Q5yk32Rv3f9jkMSWvgg3eqkTWEd//FDkyY9hXKY2Fody02T
Rq0EyBIn0SJqmn4PJPSYjrocQgugv3qDo1cpio9crGPa9C7I4SmbbUi/fLou64kg
2lYc/Q87u2jgt2IDzbreB9I8rAWbgxInplaj6RP5IALXyvXdszVgiY+Aa82gGtXB
TAG3rg/ajsTyGfs5woBjy9snUUiOD27fh0fck9WMJG4YmGyYlilqMnC3PyY2wrN1
1c+W6j4aJOVGYBzW4pg5JAB4rxOz01ik+1Iuo7PfttbBm6P6NbDhvxKolUCuaGRS
+vlgEeDhtrbLvQ218AGs+Fuo372HVVelyth9BNfN0iIlKcNIYU+2QM0wzjE9vJE3
IPkx5Q3cm9wKS/Phl1IuOtIE9tKjhetpSMnBkGA2PF1voDbgfu7g+z4EqSR5wWxj
ZsBrOaRldQsLfap58JnQJe6IHkXDu8Asl294IW5tgMmidwma3hvq0473jImNU0jO
/ama9XIy18jNYHTqvx8yG91Vo7EaZvmfgb5vm4m50daIRMLGxrloFiS3jvrgnJO3
58s2OWsSJU73Fn97nW42Q4uxzX3+NoLI/ZGCG/8qu8359y5guqhNBKKRBl+J3VWa
tIPytWsqUvb+JmKFcJnuGOq4K1FS6axXO6iUqgqENgbpOyFUznc0bePwVA2E+yJs
FvVAvooz+FC2uEu2pxJr5z2p7YwbwqoVRfdit1hICud5TjiXc2A31+bCFWMJo2rf
JiOSfkFRv+fBwzPTqpSr8tKrd+eGwPA9wV4cE27aYIEB9IExQ7Ju9MMhcyOCp97o
WH+E4TgoJ2f7PNKbLyxMGNeqPCxpBT8j8tMbt/+qk3Vs/bGVIHgOx3EnlBo79zIf
bhaSlMxLn3lnwO+Xt9sWqKy5sCw9wuzSCCkSfb/O8ttYhB7TbSVJyO7QtuGmhtlq
GjuN+I9LqkXRaTkqHw6/SWocjdBtFR7NRCOaU/zFKl5PIFp055Y/nPTGzQ8bhYgU
0PavokvPE+S7+8O8AnlCpQ9DXomeHO0CuaWpYKEQXWYPSs9H+axYVwwOKJQcjc4S
sob1K0poWsIY61j58rb72eAFg22vfgJDioQCcuptLbskPJ7Gpg01bjMcfBvqXF98
X6Ww37n36Fk0Ixu+N1is6OQmHawfFMZlvpF8yWlVvi/c6aGUPJd70H6kI8eNI32l
fr31neAJiHy7IxmOofc84oUNRTPfH6WLfhj66ENLFdtBBOvP3d4HPv1kZHXnq31g
WwQlwDIECylHCVlT8KzOtraHRcKCsz2Sf3vU9HIwqhwtelN0bXI/EIrmQ+TDoGJv
oXEfpBWTh8aNyLciIxU1+xUgHQfyppu1YOJJu60Wc2wsuhW3ZO1UO7+A0O48m919
HPGATgSOaaShO62h5wesn6eCP4FTcc+WY8mHRP54qYNygZyoSkU1qk/HkjkgAgJJ
rmkAIWLUnpP6w9P77GopT0XXG5mmUwSwS9QxmUl0AdQVEEMBYi2gLoVd4Sb1+fiQ
wBSrpy/psO7JEy83qePp+VdZNYN3TiTo7Jivvx+CmdI2SbjjTFeLHMtn0mf3met1
XIR/u+04h0Ol2jYKGLrSwAQT9aSLymHvgMTcq6LbwNN1hNi3R+KTuhHY68EAsWcR
s/QsaaLCxTrGkW/dPhBKgwYHkt2faIOirNozlQ3SL8xQQlnue819RQ+Zd6zw2c7v
5YeqxuGkZT4IJLBWqeiHrc6Qihd11oZSeQkEWLB0IcAAv3X0ztaU9CaHDCiGXZSw
dGUeV2h5cqeDIDQVK+UXyzvAdf55pr9C5okfOTq/i7dOKCasCVpgoXD0t3FM6eLd
z1c5ieTtkdzkRefi3x7GKhVPvdlyvxMfOfjL6jSbEvCri4zJJMvnAQ1LQWkKf/P5
S3l6NpaqmIAaQiMa11YePFs2LDtmIvR2NJDDsmaUAb6DRu4FM/m9thv8awzEWjLr
L9acIUp/lhIowy0IsQ5ZAZZR0kSvT1TrPa0Z6ylTr/QDj83KQqOxXN0/Zv8Blx+k
iIn/ryK4PZk581VIQMRdN0MDvsWxbIQIhw74n9Wblsh3XroRw5kZWmPvPRXAu5Tm
KPi3CEdruWN3sYvdfyM/3i4rESHRqe3/4x1XfwgK9mvJCSxjArkFV6U5N0kd/wvP
HsvOZcP5jpd4Vu23EprIzraRwS9WuAqX9WqWFPZxI6bmf5jpmZF0kxvzkD+0IGYQ
/W++w+H1mjlHhazjkdV7jtI+6zfnxlXzNL281XSm444yUHYAeTWevWJvVF1CL5D9
zDU167Red+LtP+pvHidZIrd4Y+FBruDW07UkDtzP+sqpD3rcIos6pjKkRXhi/5E2
2RwGuRTARe7CDq5ta146eOw+UfKham1k/bCbhDjFcxYP+njKOLhhtF2m7+vrE5bG
/v7SByeAMOqOja4Xg+8Ve0GOFmH3r9m/gLxupfe6n4u4hg3eJkM0Twexr5yyuDUO
8FqXJWM2uJs2oXwzYM3aZDt1HPvPTc1QjgA9cQvCcFXkccYlXxPfpKcgnSCOqDfW
L+o/U9vVqFqgU/uN0+CdZ5W86PbvktgamingichvXtywC28eZk1ohWTprUGhNDzI
9ytPEe5R4tDXz+zmbsefZ6JA2lDztFyCXa4oQ+KA+i9rUxOTjk6RJNys4lw/xzWt
av6eqd7cXQFniPDdP+AEZbYFqOtdArlPbotazzSmJWSKfamxDZ3uPjpeizh0dcf3
3co287lFzYS8J0Hxrhs2SA+Hpjwn8sijHYTuVQVzpizB23DRWxFDSuP+f3SlBUm4
upweObJycH1U33Qao5Ny+gkO9kCXjAxz34iOLm1TORNgNDnwHI8Oa7nUfOfuAtyF
9l0nfO7qKnPQiTaGmw40CPE00ECEmBF9qAvD13txKPjBsU73XETQI252lnIBfhrG
6mSBUwgBzgD0ov4c+1ubPQNqbrE1SZ+qDzz8IXBe3ii4A5xpNvzf4weKqAhfGqhj
YMu2rrxl4o0caNQXffelPQmf0TqIqTCNYXh9IOSdjovOvM9iGsUgQ8q9qiSeP4Ii
5rYB7tNspV3VybnuBssZT60Oa7C9j9mrWn5doNVlB2/a26vAfo3jD0ts5e+vTUFB
9AtHHWeIdrWkCWUFX3RaL33opa2vSLe6l34beeZBieAt5duErK+3PxyRUtQ+ZLwB
Q+R3gQ+MI0LF6iiZSplJC7tPMVeDQnmHMnCU8KpnNAt9Y14B6RONOQIovMaVpNnQ
VA2WhnZrcCKqDveXnT+52mlsHiCYGmnN5+Poz9fk2H8DYUVJcRHfGPntFV/3NroR
pyjXMaDj61Wd4/N3AYEvcFsqDoAvxys8VeZj4nekm1k9nqC4LzV2pidbaoEccpVf
05da1k31EV09P6ANTHPe1hFnLZFyPi9rZV741DXyjLuiXb0S2zsfRF53HzHBjw53
8X5drHAewpUJT5h/Bywc3JuYlf0AP7SZPoReWfMiGsLLTxjTfx8IDOVKcr+RTaVi
bPoYc6t1W9UVzfPvTezxoZoNzraE4KdsMt7QvMUG1262IX7M4RpCKL8dB1dPzwOV
2AZAgh/DVL+pZXFdI8K4lP0CD5ujdYV1n4lOBApG22Zmfbzr8yRsrznwcYQfXKTF
yek9V5QHyhUAvA3Xa7fsDGuSO8sBgmixYdnDgQMj7QEARSoCwKUSoHOSVVibJavN
6pwJBxv0zz+qkbnYSSacTq4ta2rgqsdpYquTJrIR8trWs6wMw+wZZMObVqty7/xm
OkZr6cNUsThbgXVQlLaHM2HNX6WwTII+v6vNDfO13qwx/hY3xwYn5oyZU9/N/Pva
pb/sYCVmSwpzxLy69M98aUgnxKg/srx+b3nxvzsHcCDJ4iWlys7GtUN6ULepRqsO
r67+lKhYbb3gnbiCnpuEhL/Vi1FadYY4vzYRs4LocyYLvFE13apXgLNGRG5hgR+i
D8Ok7ERqqFx2FWBf5d8HZ8K61LwoZ5sxZxaNUEwGTItJsQ3TzLDNj4PGcJk5O0h3
L8GsHkUT8ijhm5pa9xxbAw6CxVCp4t+W4zYa2ji7CkfEKQd3l0e/vMsDGO4sG+hA
gkfAIJlxQ8LBvSsIlMjNQZGXBr9z+rTWXDjpWrWHBNK0W8a9pLL92V9BNC4RwFyP
9MTpkxszcp2M5BzNlcHpu2sVdZF4GlRqEXFY9aQcSLg3Liy1sdD6fvm3o23vVRcR
1Xau4TaEt315Zq2+P6ziPRKo0ToRLHf86qxjvWKmBseA964UiLChykZ5v3D75pSO
ddnSlKmQ/t2NsZxViphQdcZrfqDLHy0zLQryBAdNGW4CF0PkDsAzN3bXanISF8HA
aln9lRDlYTtZyEicW/8ulx5x2NUocGF9EGj3KtD4yLjx+DV9mtcnUaEV0umQvnqH
TDbVIhkp3QF1tAMJqJ6zaGrsw6i6zHG14dnoBoQR4ABq3vbmeXZpplpiB95zMGcp
t9zp2bD1t2XfCrMSdsYYmyuG1GEF1vHVfa/9vhm2wSQaH+r9oJFpuZv3IAX1SZFJ
IDFHVJJHlzrXr53uFwXiMJw8VXWda02mdY4SOitUu7yTFz9R4eYlf4raBqJrzRJs
FlKCHvN6pbDUca5/imDyzpxSPTfg0a/5vbyHNRTL+ouc7Lg4IzMuCurl5DA88uEa
BV5DDFubS+lRAUHXq/siLjM2mr+whndV0zLxbI7KjKxefRXzfwFgrAA4ZuIl+Aq3
C0ujQAXxt2J78uWGrib7MIcFF9cScvuMOjfov+y6h4hnfIjWG13XnBY62PI4jIuh
4scNYeG0eKOATzMPhi+GMyb9zljPrSSDEqtL8ge3gnjMVrhcxxMe34eaVjWg+iQj
pCthd3vfZrEoxDolTcasYd3PupsX48ciCjnd1ucCZokbPZpFbUdsinVJn8bXFDzU
OIG5G0GheWCwhaXVxJ9cy0dTsM6iGBL5XmyDluAOCRzadAlwy+8FAdF3dpkN+ODh
IWCerZM3B6MQPnSAyDXTvmRx6tEUf43FrLucRLTxHaUL13S08TRP7XcKZemH5VnO
8A/gPZBqBHvuiK65j0Qg5NMX+ttftFL7/Tf00cwSrsVYgPo0z49yM2vKKEx9H5OM
V5olCJonxD6Qdk3asQS6cXIF5orFDV2XREGPpD7mkAyfHg1X+rFYY7iSiLjUw7m9
1ChD1EJThaOzXlT5qPLK0iVkpK7rb+soeIFaVEF9zzRM3w+f8YQDV34LcMxcBNRB
5VsyBj+gzdN1CiWjD3vmua12xwIjLuXxy5zSLqus2bVrRpP5EyHPcJcSCr+5IpO5
0Zq0HlKaGikPjxauZHkYTXVHUc2xTyYcn7ha1arA1fa5ql9XcphcHwrzZRBGF5Kn
NU6+VEWVK4ahPzLyXDKYsQp7JufI/tQ1+ejSOn43Qxs0sabMlBdHaLQZXJNviNHp
I+O1WeJGj9q5S+FXH4m7OaAcnOf96eEAzN5RLyY2vsGRUUMVBPK+xOaIg0h1JCtC
CZPSlytsSMIuL5m+tWzMYNka1803y/JM0U4cUyO9K0Eb3jpLQlqVXw7GplMRdEgi
l+LG6gOuop/yz6pIcT+UKUsnAg//x1OOSu3rFQIkbo7ShRaWAP0xE6cHIkOB1JjD
8U8iWHRlwL/EDTQVe8p0UP8zK0p63V8SaQFMqzfvLtVtCe5ZytbGsyD6CitjefZA
WxSebEWxCeYxYRpPW9k3r8LnAnlJtTKxxWzGk34sKwhIE3ClM/L4dUt10MoG5l+/
i+7jPk94aT4Arj1i65wzff0W1bHFpEXiz6nFMonrrj2zx8yvJExV73lELCSlw4m8
huij5jUfwl16El+UHqxL/qrbMk8WADtflvfRvGbs5gkNlLnl7EevuStAht4PsZr8
UcTLe7Ir6NU043IT19ZLiDbqbBmNWC1wMov20/fuMoQYo9QrX4iQ85jnY+e/LDiz
rk29nSZpXO9J9C2hNROqdmmvY8mon7dauRExdP0gZVY2JGF8I5jcqSB+jbVFu4MF
NK9Nx5RmWR0Yz+IPThHIAC0tTuFR/pthVWq9iNWBC+YTQR6+SLb7hDzo+/GVy48v
C/jSdJXY95myuMXmgKZO5XKHH1hNIb3WjEJfRUCz/BjR4wyerEzmXyoUVq3V34bH
nvAOwuEXZvIGILUKScePo9kzcdN8IjpX6zECoLx9+RJt0MMmt+ppC8tMgOjkeN6f
C+9IoLH2a/gU38NOtjPTdKx0iGEXXU4EJU1UHz7PO4z6/1mfD6U7ZZWGVzYWxszN
paIXIMwR0PvlNA+GCgQGvKKIyDGgIXiwmJL8QlnI95esqRzYnwYzvX9IIxaeRrQE
quCRA4KGEpi5g9Hj1t/5ksZF2aNXKpdOkTea9MQExoNTa8mOM/kjBV1cWZmyA60q
sqMo+R6UorByMwukjCGlp6QIVocUP4pKre4iH9697VgrHt3kXBB7ToIvNiYhOtoy
lYrRlYdWKMP1W6VLBZ/sc+dtfFqZ0ryAB/SqGboTyYWm9pgp2FLJTVN1yo+m4zco
Zv62qybtmqUXS58XaRTirJADDf18VziGeUSCaZ7SeK/CxcKh4dH8L+oT/nxG9msH
OBezybVd4TktxPlKiTFEskUt+scNafhB4cqE3b2189bvmOJBn9QucWItlL8nzCgh
Rv+SSVKUAhJvB2bMFXAs8KnyTNcIZNnyFxTf9QA0Tqf7hJSYnLzEMeCAOj5ac08Q
HR48+TTmTAhuuKatXNOOqDsQh53WnoYEcP+sBvsOW6d6hMl/k3MMgGy61+38HUWn
yoalqlA8yyDqxdN99JCE0L+LcED4k/yxpj6s+KMGN7iYxauVUeZ8LVe/iSnmO1E6
pEQ4QLMA0IMjf4nLaF7Vmg7u5OC+h77+HA6v8nWMilYWh7gpGY7IRrsPPeCnTY4y
pzSKUKJ6heBHojOvqxwykOemDbX63QtVHx9lNas3azHKIE6ycHGw5PuHLsflBUy7
+GpdwaFprFq4lsFHPOdU7bVpncFlMkDsXgIK7ZmH23tY1BZr9v5/jrBLqwLKArJk
6373PCfCIvTwMH+S2lkC4MCGXHUARPdPamb+JfWGzRGjK6BTuMlYimctCcszxDIC
YpVYpLxjqUzRu8FxrJuHUs2SeioyM1KfDw7GV8FLHT/fFt0gcSxot3IryvB8OcRx
STx+vUgGjy8kqm8hMx3GmnEHib6lN8q9dPtg3qX7b/dtxbZWGyGdo63BYgTAgNZx
8a/8QwARmq/XWTFO2Pb1Czi0PsHa9I2e3KF1j6OmTEcG7BvPoaYyTV7/4FObz6A4
jrnoBf1nbSgJGlJNfDBT/zTmyiTQ3oN8Oug9m/w+wHFE0L3dNAEi8AdSgAMQqHmQ
QFdtZYc1R7hh+FogO2BmVm1Fq0u+/atpdotTRsxxk15BtAX/vGxmvvMTiLIoTgqF
EfBkEkK4R3wpdDoAuh9Sx+xHpLM6BgsplQKeKXWdpGoK8eOryUIquWybPtd9rZZG
IqBnjX0KmcvJCvrruQ956vkmiXbUig4hNQjfhusriXIbmPiX7Mi8egxGt1MMevW0
/Ay/nwLuk7ZzzWTv8ECEjyzGK6RbeEKi1bM1HN6Or/mW66J2R+tiCt0KOM2IzB2T
Y3/ltHLY+0bjUEGvak4Wsa8dwrbpGA/ok9Aw8DC5rdvzkV3VBAA7Ji9uVShOV+Cx
f7kxLDkbow5/7OTuTeO04eLGi1p1EIo0XteLo6/vaE1zTKnshG0V3+kslxJHQnp7
5MsoeY7lbT7464T1Ly/0SuL0jiC+0aPUHTYGb6OaevXHeZgme5Zwqz5jYBOBzZ96
UzAYlbnDWF0zcFcJiC2AYPTK4FfrD00Fj8dR8FY7e+VfRgXc8HnqfFaX9ca06adP
SsK5N+rQ2FLXJ2Zbhuhdq5sHn7/XkLPR2s8FVgfW+szilEKHWgl5EcWEZtG4Ap0U
EwJXJgXyQ/qHxiq3/fR1lBk4eIbSDT/S2V5WaWH1yy0SVpu6G2EKh+a5u6Obva52
Z/0PfxEplbEhbRIeo6TK8Q8I0rcU8UD53h8nFxLlt9Mu5KmBx4DLV3PKer4wCz7d
LJYufbl1npJ6h64TM4Z0DA/IMIS/ZJpkKtKQimKB0tWaqYfs6Z3kJ0X69qqqMjur
yl/R5Dk1y1zagZVf+WxNtKMi1AHemegsS4tYSDoDQYqcK7AY+Us75k53Z3aNXBo8
kElK63LiEtq/p7YoA9VYDGu6n9iY9VEo2ZXTcykLL2aZ4l6Lire/7s7vTXN1JIpi
yvUGqIfFFJEkWJRNTh0SEKm0cPOiKZCG8FWBRPijOcxKFzv0qjXjuXv8tn+IkEY5
d1G48IY1bpHVQVEeewZuO31dNARhtiAblebl2N307vbNJqS6HQRB2dX0IV9OkDkr
WWVhTabFA9ekj5wVFVpS2GhEjsKXPdH28Yd983/cb3i13WSWhjrP8jooRNSiPpKe
EVoSn9DxWqVr9g4mrSK7EMZpufxMe42sLPzJV4ik4A4eUWCrpHvQqhIr880bqb6T
PQDmucXSolfwzLN1HN5kVbOW3LrHSytYUbAEYdWwwg0HeCmp41vL9wkKkVSIo6wR
YkmOZ8caM8QcgoFTZaz+mXA6r0Oca9jKnrsI83w14TyLwXa7xn6ifwuE76C2YQGC
0mjX2C9Db5OogYKSXZCRvvwEUWdCF4uvpQiboarc4Pgyfk0dl04DpXi/qmFPKnC6
FD6PE7/nDbyZr7qcEXxzVeAZbXiJHHKGwmdYQRUOt1N1TUXE8asDIxh9s9K12tQm
bK2o7VeD47WTlodCWlLarJw6JmojaEbdFrdmmGrX9hWm3MU2n47GoYcdpk4Sz3Ct
7nNCYofNXwhA67ntDY++/niVfsi/UtoQsk9yldSRokXRgMQa/zYaP6Inwjj//nUH
WfwMRtV8Cyab8MlmwqXqpxAzn6oIj+sqDiyTu8fPqX5LnNa8W70yDDVeq60Bvf8s
VujR4czvYLr+0RLH5TnzHoKaqQ72+wKZ6J7W6VmToztC7OmVW9lZwoTzhic6MtxA
W2URSrFRo7Ek7UaauPWraYRVTSuSCryl4tYSbkcCpHBJWmDhuBiIy6TfVimMRSWJ
xyQqf6DxzvKtpn/5FqvnnaEyv2FpjRJLdYxaZ/vPl9z8CvrUV9PNG9BdQqZHgJr0
eeZsSz/IwCRX1MISySUrPphq4zDC+PjZzmN7oGUxM+K5TddM+VL+vshvRvDucVKt
Bqfua+s7FI07b9dGoq73FpPd+CHlUkjrrCsdsQf/TJePSwWLSnJwu7h6UstaU0Qt
P565xgZK/HTguUmtta/yPLePjV9Wm9+yKRhd7WYOpcbvvjfXvWMDNEtDHT8irkUe
SoF18riATRsDk0oCCx+/L8agHM1nLgedy7GL3iqHCpBzqQfD1KsWWn6m4TQf38Ij
3kHCRn2LiztR7jjkvN764TYr1OGQ914veG5SsB5z5kTYVQrpRtedsWmfBWdjqGmP
Sp5wCb14BRtZN1R7W/E8nlXGd1yPuA3CHMmsTb9CX27gNcafNdhV57GbISJKtGvn
jutppdCSzS/oeFMf+ApjxnjANEuvZrakJsy4DIzB20Sk81qbQLzXgzSBVfRpdPos
K8gdXniex+JJ1mxPI7fwzgHQSwSybPPo0bEAV+5xrn5HzA/HyVVBWr/N9fU2eV38
5fG0LqkvubUb3VTKRlpADC7NM+7wOLt9C8lc2J7M9ypsRL/zEPacofO8T8wbb5Jf
VKxrUqfL80XH0AjKQMzj3Y6JRhRgFC/j/i3dRA9e0LLnBLnb0s68bYkxBXv117mR
OaYcl//NWjsK4qoLrLs7+ZALLus6clgx/0X3FoGakTmFxEx0Y7CZkkjsq7t5IWlP
0txdRlz17CG5z/aBhdWGaHw6iyksHOA+L9XmsG+uKqm+kEns23dpVyW//eLVz772
RJ23sU2tSBIg7kL6SiiPOOaLWhxspvqbm8N3Ig5Kwnm4uB3GMu9EldYSwhCa8wv0
baNXXpW7kje1ayq3Ip/7M5SCGZo5odXgx/ssMevIhHD49DrVHVRIBqvYbEcIopJk
XawdziLlKwpMjdLK/6WUnENEKlCeJ+YLQRakdFl5LviHtxwxRnFXrNmLajVvYk/9
23TMVn669oLL3FGFygAzYkTq3w3V1ZyaAExrtYg2Oh66drTEXhpRAWV6YPr7uoas
89XCwHI6LRD8MUlC3xz9WspRUvWItyrJHcyVjQO+wtIy5IbQXYQsxlqhBnLBfm5r
yRp8c4FDZZFFZN6ppYdF8JYgq3jkIff8FfHBgIeBPWvcWXAtsHnNXeAowmdteb8W
MW7cyGsM/rC1JDQ7PpiSy33IP6BUiNnmHGSJH7w4nGnoI+VaAPhEuLhTbeQWcl/k
z9LrHmS36nj9UM27PdAqN/+R5QLr2wDTH8vosnEMSJRAuGLF1YwA0FshTgIIem9l
s5ZPMknRcDjQOS0wfKjxpPsob9hKjmjArGSgvFd1XDogZ1lJsyv8pLB0lanlUjMh
Ye7BnFXLN1kk4AThuNveiI8ENJ1zRalzdt6tLwMCnJKoHPlFDC9Bw4ip4yJb3ODy
fZ0YrZTBkv9sE0o0oufKcbvjlyroTBj0ug93P+8HyBb6lrnuQO/i45yKIODqzM40
peKB/CHLEqu/Ivth3Y/gmsPDMxlJeYLabxLcWccjHp3Mrp8fI0M/C1YFV2aFelKi
yQ4Hg0u/2MGhdSolCDJMVJYVnbHGotpctbtN8K6bGruc2JplT/uPYZOin2c7MWrh
W1zjZ0yEmmN2H7cBvk/li8ImQyarayKkc3xPtdxK9GH2tZtQHDKpdCW5Z+/cginc
h0D+dCboSFBhBBupjt4dD3gkl2D8L2tiftAOUVpGjQTtBoXGVGWXF8PQ8MrxvYX7
muDvDuGjL4FgcMNIoWlWrB64p+PTI85smV2awdyTZdjjC4Xm/dXqny7rTYiUXGSF
L3HJEQQzyTEPJknee9ZlT84DlYe7kATOXrBQ7KuyDOlBznRbVFyr2k/8DYQo5WqS
UyWtLFisgSO2NJmVtriQs+i48DcN4mhaEyjF6/aG+ICyCzl+KlbmrxbiuK7QxdRi
RLN5L/1QGzZfhHbG0Q9FEWYnuyw3ETSTdxoUspKoaYkImaiemSs1+UcM6389d+tk
oh2uHeM6Hj5MqBRpl/Af5fQoJM/ZfN4gScuhUaNAVdQdRU8VH+T3CuM4EygfI0ns
UsEJeiKj3sfdSILBrZwk0U06MSuEfsNYGNoVn10XAXhWKD8uGUm7UmzTKbUDDO/N
j3t9TmpFOibGOkkZ4VFzDNub+G44O0uCx6OzV8eQfIzjnx5cBDt8lFcZJtmkFWtj
Igwj31ZjqpuBbHA9XNOQRMLBCMc1n4amP2kSfCb/cRIJkCsIMnDu1HvvZgXTScew
+jBUOig493qfExigi+7aMllINFaJKE+g86q+chxrEbyZgNJxwY5IP2UhAJZgtihu
YEF4xYmsOF8Q3lI+/ntM9NyKEUuNZEUIx80iWJWgVL9i5fOBSqAi4EkdBdjg1Do1
RXkFTiC+6mmEb7GEl6lJY0gp0wTVkxCdzGtTfsE1TllB00WNDano950nGy0rc5nm
jkszmsVWR/rXwUP4Y8oFuiFa84kjV6wHtCYhJ9Q8IhWUE/ATJBq7eIut8GntjeIY
kzoUAeGSYl2kfFAxZ8TUVmbYT9I074QUN1HD+hRGB8AFxqcQCxQrTlpfcWGGYw0O
TbznKV/gGN+PgOmU7kem7XNiWyCTdhrGfsZema3ytr580AYQzeEkZjXV6/bGR2qr
4OsbiQRjvj7E0nt5cXCgiWODHgPICP0a6BHas0WLoNQ0DuVOEt+ZFOwL53F6qGXx
NMhF9pwmq//+ivNKM/10r0PinWJdDea9pkYeP/vd3pVAbEdRprkB+WFixdrdE+Jo
/xRWfidVC896ZFcx9Zcv5QNT82I5+vZG211MlD3DgMMveKQlhv1jwhxXQJb8lVPM
MYZyIjhP045ax5E69sBxvavgEy10Y5MugW/rGg1xTRW7Wf3g15h/tF7aK+73Ab+S
+OosurL4uYXcUTHMS8y/nJlevwtZbqar0hAYJlDe5k8CkKcv/x9tjzq/UcX98wY4
QIk8PoKD2ejlFdsIM6TBFuaWw0rW70YNJkVlDcftEjNh33PJaqEOWUW8iyzy9yUk
FfiTVjUQ59CqvAi4esDxSeFmBxUUJgHHruJkmws2mFw1JC/oS0Y23fs/IkbkHCmj
HwnAis0T/aRujzgjKQIfj06grALLXsJ5ALw/Tqkzy5fQrelow98TCFNzNb96fXsO
I0849AEJXUhxsv0CG4By3lZvMq3LokQotCjryOv1g8swYVA1DvG7sQ6tuoDHmOYB
BBE2x0IoeOLg6LdwtsAdy98A9YXIHayi0SI8LiSmFrXjUsT/8It2TZleCKCFHlRK
sEC0e7sfyL76jBqkUd3wA+kTsx0xw714jjOUNXW6L9HmLnzTMc+/Bc7j+4D4kcYU
g44JvHseFUtGcYQ6tQ/l5bSZI7nEjUswyg7509CTzKquxOstG/XSiQo8rQaq1Uil
SC5K5nxLSb6v6f7ewQC5nO+pUQ1J6LoZ1Rwo5UWvQ5IZuUPo0HV2Ush5P5fAZn/Q
Fim21ga7/4Tybi0SqNbhuWOgcRYgv8wiaXz/DkoKvYogxN6BxsYA40OsgDCEwcNi
B3lCwWuplJKssZXJcdhZ6jFyMjn48A28B8XbmzzQa9fCJiAXEgztmXxornZPem4F
/KbqooB0z0Xjx/NALWsQIiHzK3C13HYjV9q4dUUJdQY0Mico3Jye+61V60ku3iX1
I9m2rKMj8C+3JShYu6M8jspfszoxS7ba1drNmT+hl8JiZuv4ZirzTf/3/59mZiOb
OvhxqfCRwtoAOAqjcqjjtwVmOQHmaZzpxmQFIeW/b7dvQUr8HNkgCsgbaaCfSUNe
L8Poz0ZMBx7F+rFtA0t03x+I5x7r6z2gk+Kx9ME1xzBIXm9rt7JObbUZFDh+xYnP
RPqicotk6Xnko2PyRayV/WkvM5twnIlqN9bFXxm/bBY3dJzWd4W3AfWQUqmeAuof
kDW+JdoOrcxCEiCnuoUhJNeGgRp+XocUw+i6N/sKa97R/KH/jVGg/pyuUINbpSg9
CUdt2/2CZ7jn5oEb76/hnHla63UsmS27pEe8b5gMV1vc0OQ9sSXw2G+5JYEao3U8
8C4mGCf/jaItfuu7xHdgkkqbza5M8nA/7ePQLRE6os10jFwz+/MBSOLkYDPxTbcg
RI1XuJdMNEpFjJ60pLXEmA1vG3ckIcrKIHC65CMZlzVcf1KflHwtHqjKq/SqdzMT
UISNRMNHtUsN+qfI+D2Ho1CfuXeJdvTBotGU06TNL28SB9RlfhBJAioSzaEbakYl
VvIOJmf+MnXDe6NDdztjC9iGPKxH1XuVYaM7mkt4Xit85h3SubMO15dFBbds7nEB
nrHeDVF3ydCwhmvkQw31IraUnJeOFySulLOWM73avAayjjuWouOq/SEBPbcHEjGS
AywydIArXDZ8XFMtWwsBd+iiafeMKAbcbCOWtIwKwXSD1yqJuU03KT3lZmCRjwdy
01AVgBpPgVD9XnKQgUey77Qq6GJvxNUJoNqChwOBl/E3iCFQ6vI9eiKuSxboCaM3
xvlhucpvkUtFE7qOGTO+LmLBUWA2ReCYiVG83+e3QUvaEdgLlnMMosAap8+z49/N
Hxwh6Nz1OUPEisscitQx3n5u5OO75u56ZGZ5gdKn5uDVaxxKsmpcVuhSuf5n+bOu
bz7wbYixMJ6y2EMTC9PGNp3OwKRNdUYCxupqBvNfTk6wFAXwhC8mPrz6S7CO8yqb
G8hi33oZgZ3DnT9Ub9hSnAIaJDRzNKRs4VhdMU6up4hDaNkC8Pq/xW/OlSjPTWI1
NpN2S2HYkRm/i6Vp0Y7RlqxREMa6U6A/wgiglJMp65xk3dEjjqgEaH1ZgVTdj7KI
1/RXu1n+cXqe8mVrcSBALKW1qFGGLEsYuOLPx6QwLSk2E4RVuLKpg59xCbEBe3+u
mFo484EaKvGMp369zEkRenTTu87QkQZi1h54n6eezxGi4BBTtgtmAxVf/ew1SYrG
BHKc6FmreWNY9IW/KPWaH2lTjCJamb84BXJOGdKo0ckNDgnFmLZ8TBMWz4mS5fhM
20cVMDwp3dsqwsYuxx+rZ76PEYOQzRSpLMiS9QrUX8yuMwAbHi3F+oVgkHQvszcg
XyrkFXf8W0ZW1XVw+L0T0ZYHD3kUL2lie3ffMErIyz+nwlxQ8rs5GqSDJ6W1eR9s
ITO0KtBFwZSJiFoLbUSXwZyz35jWrsHiIIeaD0EB6Nqh3zSSI5AA65NdKhafcBJE
HFWAcpyKFreI24FUIDNRRvSM9tCwhYybig377GxqRT1mLRsgqFdySD4v6Jz3xPix
g5eFkAdylfXwfosC6/5fX9yIS1ZrbUJnCmQDlBi58104tjk0GPF9FDcWGjKGUSKM
81JOW7ByPnJmYOa04fUufsAvBxhDf8+mF4ijKWCeGHNjdLs6r3qJ0JKQjh/N3131
yOhaI1DAF1/H5paui4uTQcdOX1EB42fL0P5P1sLiD5C0cJDAN3MZngTbmkUqXVuf
JzPrWEIz6jaHYmwVvJrsf3BxLDjzTg5mBUxLSeeCtEmh5Y7ownXvv13m10wR2X0Z
y+6X/rt/V5e2tVoniVbjPmD+rOGCzYQDPmlfqHHwJz7E+oZMo2oO543nbiSCUuKU
5XmQWmnhKGFq+1H47+/01WsmH9mYAgcA6e0gthdbPb0MI35wABLUJMjZWA/gKHNd
nJQn+/v+1k6RAwNLWKABQwSjeyFLydwhV/jLxM5RWzoHzuPmmULoaUUMIhP92yrb
YofV7Gb8NeTr8+ALW56EOcgCkWExCVGBj1GDbCEiSPbqj9dqSHGAu1Et7w4QCNHJ
jVWl0qz4CeArQ86DFGN0tGDLUt0UO9UeqMQl6hslM0L3Z+/9uJJmfQ7Xj046vPzh
Xb5oH/l8vq23r1sJdDq7GFHkTH/MHgOJX96sueYz3uAV5aDOd3rf5dpN/aa8b8ji
6qYMYP67L7nTD90FM6QYR3o2jonQHsc9W+Dn2TBlg3FFurpen6/ZrOmqQuG0TE+8
1WS4/30MZjNe6BmKOP1KsGAxVk2IbsUhd53LosejqkL+fQkNLagibMXVYzapf32k
vRFyOwJEd6YVDeSuplUlOtOl2IUHCdEWRelebhJHV+hOt7mGQifriTlEQlLnVRfy
DUzRp37CXedQ3tMqrQWQbfnu4uKq7QLnODJok90ua5gENPSdL4FJuevdCvUZkijs
VyJobJQ8vp060LVbg3jecIvGcsQBoCn5PZCr0eo2IU7999+ygSyOiPKznpFHVI7+
T0zy3XueJFYMYKuo8dTKcIjlGmdpAX5N6kyDsKB02ty8UD/2yuGEJ2cuTWNniidD
0AU/AKX8Y9c/qb02vEEtG8puxU/4PsGw59J3NkkP9swR3dUE7c1zLT4e9+NUDHOO
oC21CxZzNQ1AfiWPZ1BqYt0/+Dh0Z1LCq307j8FEPUC1jL3bIrTkYQD8mHlnLIG2
kjmzzvioUB45o+MGDnAjnrs1+T1Hhfavh3K7CtZuGMmi4AFjMqrWQeGYcqoiidJh
u4qhTDZRrLM2cCwaj1i+DQ6aMf7ovhfMb0zJBRAvS5OE0AzMXtOWrtdHRYOQJvmJ
TBTsfPGdatGU5MBZDCrFTeViF2YmkzQ0yWVcB5SDmPey+XRP6VdrYUCXaDgK9lzV
p5xMHseX5gQU5jWxLmuQsa50pqaP3dbCCkUf8xaJM99KBLMjAk6BkungGJNJM7UE
EUqc0yM87Ya4JRMARTZuTazTcmQ96nnSfU1JB4Tjoyf1HV4rQ6Rwq5uUjIkT7pAj
xFSA+UKB6Za5lzKNv4A1jnl54Qme07fbywjlAe9a2JVLKXNVQzVLDixtaQdkkDU4
X4m+jllMp1wkQYdbNV0jxeXI0BVJT/Jop7CSyYW+BBFytTZDgsKtD4kjuaV6Hdc8
0R4J9a+4nYVm+7G6hq4cdIerSh7ci1BCE9A/Zqkqt6HWCsmlNofsJfKwqJEbBi7d
VfdeOFLLq/BSETBQfMHClVw/55Z+6j8aSZPycA2Ji1VrFCKsNoRbj+Xn4oTJxGQX
h5UGUZcHq6LxjNFV42G+/I2UpI28mDPxGTWHwpN9ZzuFKvw0BceYraT+hLUw/eD0
t6zm527a/dFWhfyz2QL6rhCicw7Q9QXvECOgcDsTdEHZ5D/ZrwsSZUlyXGrfbNha
gT/zkXDVt0Me6YnC7ULQCfmnjw0DdPHLooUyHVVAPcVIw2HW9uiJoBke7B0AfDdJ
He2aJ4AzHp/10Y6hxUZHzLblo1J+CLSbDZdM+ZpVRnyxPmBf6ioyw2GDK+RWkiuP
MP42JBmsBfGliuel7SOQsRXps3Ldrj5ZBG0+Rp4TAY2HQl/f/pZEpj5LQ8B5pu2d
ooKKzONByTQQ1SMfrggHVUsQcwA3GvZcRtMNH+/4qAoISn6SBUiZTBwc8JTh9pUu
wVHC43YJCLUv725WTWpi2CXEfT1qor2HWE4DsEJH81yiwerkgBOayQrjW//B0YIL
7+GV8y0eXjyq7TjBrDAeZChgvSmBKGVYNKDoDK6nZfZBVdTqq0kyvvSBLXx7FsBC
26z1SmO5u9H7Vm8xHTJQLydjITd5HWde2TlpuDP0o06yzTm45oQ8nj9bI8A4o4fI
hgf5VIFJz8KmcN0kVQrR7Kq1C9VfJY2LUuoL4L5yNHxwxM0w5E/8iDWoZ3EtNe6r
SwWEJxecCw5uN6HZ358CtKiILHkF07NY6NiIY9b/FTFf2LlpfmHkui84V5ld8rUp
Qyb4Rd8x0KnVaQAo3MFuTef44Mh9j5JH8FBv3NIBEixkmDYFLWqktrS+lzu+1Tpm
aaDvHebQM/Dn5zy6jZAc6H7C76eX2si7MJXuibozBhnuLY0TFZGmLv879btc0uBW
K+pILx13VKuavxhL1R5UzW61HvwpG1tW+DAkE7m263f8krQgNhRSOyTni3LSDYA9
gn4wbLhQlyvYi+rGQ1SfHHDrEVZz8QnrTMfCEVS9PlFwU/uOdxlo8AUlBRoHBcvR
0nzGqGrx9bLK4bv5Nc1LHtKLe+wjZEGP/+tmh7FOmPHwlkAXk6rJAC9cAIl5ajbz
ovdXmjel1LRPrkay1ElTe6tE4j3ZRuFGhatLPCtuTxs55Rrq4NqBjZT2g0+lZa9i
L8BomwRBZ3XPbvA7nW2fEN7DOOiuY8deP1T3VMB+VXVcK7VYm0pvhDxLTAPIYfy4
ZDfVeRUvk02ArXjWxwY+dKuGVSjjKQZ80HjEEviRf7kyp4Rj2jUvC05h2O0EPGh5
iYATH6bCpayscsYCSIsUzpgBtJ/y0wcnOVCSm4t6ZnqdNtChfXjurE3wH21e4Msg
eJTISzOF/yGfuduSKYnRwFXPGnGDRUh3k18kfo2R04SWQE9UppsexzPNob7wifgW
E6D1phf3bPWCaol3K2PfzFZgXa+ehwJLnqqp63HtAud7cFtsuTJGn6VDGRL1KB29
38rr5bNclTL8bmHLQQL1fHUb/8ObXadu8qycZm3p+Db75I1QicU4vSVtemjITcLs
j5an9kdet7y7OlNsjBRTT+pUNuRty0ebJFZQyGWk4dINLpzpGnEJIngB1FA2D77z
FThSkLQoxfbt4PutI7PLZdRDdQjsmqz+iim3punDuYJMS9YR9uAynr2Yl+bk/YlF
PMSZe2JVII+npBb0783OEmV2e47NkBYgOX9DINpr2/Hr5R97Vi1F8+jAsGuwr8Sn
ai8oXHPwQd8vln03tWjfENKrsdaKrWzuIPO5EDzRnRsnGLyEn7JQDCkPHhqKQ+lu
esD2ULUaG/PDYnpLCIvagGhy+lzAcj5ZyWKfyzjXyGhzaki+ym9HLnC22L0KMmfS
NxZyRzYL7zD7GdsBThGbuZUxB95PNX6HSCZrkaGAMwMdWc/DGdKAHGI4ezFh6/mx
rmckPOoIhKmUbULJV2DQscI7gxd8MbHg7KSQM81AqpGG+zVcjFr1Q7Sndk/sHtVP
64gh3EoPf5WTptVRFIYcZ7q0hh8AfmQs5Zy9dNGqIGSzdorS7olONaNf9Ng2uV5n
W+/Fs6WhT2GxQ/XPDsTCLcJvMlU4ZQt0lFV2RfwviMN8SnWUc+FCM2nJwmZABmZH
L+t8N4vNNu0YI6v68R+p4qASOaV6mOwnrbAM1IrPpcllwWKtDxJB8bV9KFZ6VlPq
Xhz555joTE8Fez9oacqwbVySQtPyRfxF7jInwc/2QUaLkM/s8KJd24d58id1g/zL
+R2/imNNXUyWTHw+bpqW22D034cqums6qjkWGNp/hcg/CYTvj6RetUOBYIwyFs76
CLAywpkX+lyPnhTxhF/9C9LZ3kVfEi5+WZvJtQq3QkSrlmqn6WLS0j/+VwM03uVb
2qJV9VMqNTmLtYeq1Jbzct3RrZHmYtxcufkpDjPbeDZd8mKrgmeRAiT/Tc35WqU5
25YombQ2Qb3IYvlMzgAysPu97FFjTYz+c9yZcl0MtHUJYRYjBbGAHQ/20McWxRwk
gh5HHYV3JwTW4299Mt7oxrj7EsI4NcsmZAkytEa+s5R3nsvXHoFw+bqW8uldb66h
aW5aL+sJbXrmUmVFbfRi3QW8LGOEcNLfRinVJ3QJXG0LjQ/D2/mdXeoDmJrw85Ge
cKQJqEZWpLQC8+ZJAcUmuRt4QSdOKXvIzO3JsvmUq/SrXTH2VymfORJ1bHC1TB0K
ubdsZOtdqVpcdVU+wRRpmyx+wJO9D8iuXC9ipGPweDz6ksdf49qnZLOg0z52kSzV
l+r0JSIu3eZ/PMMMcZoDIRv50xFoc76W5yaQD35upwt5ztLK3bJZadWBrHJtzXyS
cCsXWcJPUQ8aO82QIQUq/257ebbaglLdyYBIYdCBtdwL8EQr+pZHVvbBjpXQ6hvE
AXI/NTc7J7wrJfsHw/XU5S3pdnMdr/35s02j7UOte16hWEX8TrIDn3Ll2kc6HVd7
+CWPV4XAdf1agpf5qJDwqqS/bdC4IlHGfgJmjjevHK2Z+V5KI8eBlVERGvxhbhEh
iMaTe5MxosIa4Mj8lMivkXy9FSL76UKVN5p0t6TAYLs279FZyf93rq4Zz57DCSkL
q53CpW/LM+BcsQwyp9vDgFd/iap8a0ZWM2+GZjLyJu1tkJBA9Y1SvfkZGePWYdiY
2z8fIjLFabrqc5mx2HaSb+vQDyX9c4tv67NvzIeTeOBPtBgqzphJWkG2TQPUToW+
ym6OuTSDc2aLZorWkLNW3Z3OvYN+PXnOclt9eFWndGT4xqVPaCYzGyum7IdQDvqJ
rTarzOZb5MaiBal7jWmsJEY6Ktf4CExZQ50IKhBbJX6V1R6nrWqmN9iDngBxZhbm
LimYIpI8kdHkVYZqfUuBd+GskKIFStrspdeh1xW/kapv701bz9pA7BWJD4QP3Sy0
RDMlIY4H7+QBbVlwqAmYEitYFGxJ1F3fYzhjgkz0CwdnsOPLaC7I+DCgqA2WeVzQ
8+bpKuFTU3V3WA3MRWjP3oq/fEpB5duqoxw2kS6cQETgFct8whnDRXgWq2CGY/Wy
TV/fC9y5PTv7UzpYwJWLVCTi6my4GpMLsCwTO8UnXuQMS2J9HR59a8yqNUrgxiPy
N7D+Whb6D90IMm9OnPY90tCg7xDM2NPkj/8B/SYyGcvAdzGzqO1FyAXUK7zIPWek
8T13SqAVrduo92IJdiSm3pdB+pCpxnr/IJf+KbjHKLIC9qYp5HjnAHjnPaZh50dJ
eMxs61MBRLXAt/ETWTZSskyRJs102DPbZj2QfdskWiYFGIRfgGpxJfJaTjxAYbVv
ysMIET4ZS31E0h0TQKIsIpBsnU+oHD8QrFYFKV/KRT6cbMYYfOFKdOZMGb0H4d/p
gimS+pElUKWaf9qsF+AfS92C6F4AFRG6WRu3PHGIWucAUOww4rd9XKn5L4c0c5em
hZGvPfjJM/d+94VZYBA7Q/76yD/SQmxf8uLcwuy7WJx8w2L6mmqjQOoHuPOB6mYR
lsnuQ7gx8rs2Legwi+p5VTF8St9CbLbnZbs+yukUQrcl1XH2OUzWe2VZGLeWGHLB
LHo89HKF0Y2b+moUq+iIgB8VQEKiPLcsudDIXbYTeht/BoYO2mzsDq/E/Fq3yxDr
48aRVyuHWBK4GA8LGqV9SbZ/GNWZgDVbkF3QteIMY/6fcHTS0faKtu5gK3Jzv1vD
38Kt/Q7ocPd1FHtNge4zl334QeN9XQrpSEFLZFD+dnxVs6ZqUB8IY+8W8qJuAwbs
kE7BXqcFx/F/eg3eQH+Drme2fPu6fu9/pPRcv3rP/Zl3VUdVnz4LQCIxHnA10n3T
zvcYFPY94cW5V3LMtZYPlTjIGnzjRHYV665ImdPZksAH4mZMEMexvIBta+t1Xij4
RAe0KzeJxyU9C+bgOGTl7Gqc8cbKpJbGJhRYbUOEK3KVxEKzc5GZwe+8ee3lvyDw
A3TY78zQ3zRYP3W/+eE4ocPJDLhLHHJJk86eg0B+yQD3/nHNyl0Ce0Iq2lPeT19z
L7semzOhg+ts2FEZ4mbz8MAZw24D8mhsDzQcapK2aXhsMTmUGoaTJpD5ZiePVoNN
OLxEJWqUbDg7HSTiYB2nt+BPJU9BYZ+Vz9Qf8Ft2MUsBRnjh08wsMIlmsin2Dssa
7+ngsdrhJt+km25n7wB+nP01V7gy5dnHF5jpF7V/+qJ3/59PuO4Zn4xDRmkLL2VM
oC3+WpGhLIo4qvywiyZP26oRNRpn5ublkcCMRHcXklXojgZ25kuyhUIohXsm7Cpe
pD3B4TDo/ZuMPjfNXOtd3ELvZVHslVD3gUuxYp9Iv9iThW8TpUxc9fIZqNf+MTLK
mlZL70HbdeH9sviTXfRSXeSjCxiDlm66aMnRe4mAr60QMrkDX87rqn0ioxfWMMtt
NrUKNYuifjjnwSM02sf5xq7umAmaiYbkK69KO0d6B3B5oxYecBMH+BtyajYt3rWF
MhR7VevlacIUTG7I8xsxp6wgGPSnPMXM4hXEZsn/9p6Nk6+R0AfMLRfa/fqhWr+2
4OpKpagrBvp7K39tur1AjeHgzPmi5r2g1DzlH6vGVvRkntjzZFgVTSf3WuIlztPC
bRYDC357TIU8mcST3+ci+BacQ2mm40LfvhkF5fuvgxBGZ3GOtP63k8i/p9TtkMHz
sdo8bdwXYLDcx9bpH4e4nxMDSvyY3u4eOU27bMDXZFogLVhlCTy1J0kf9A/pPcL+
4G6oiFzof/4RGWBRV6ceAmQILoh+Jl/ZTPmg7tdfkLn0/PZ5Jm1Q1XpC0wJP924h
DAMy1ogcopYCWlNyxPNAOFHBnD/54TsQToQhzpeLrvCkmcR3DPBH4lpsvR092wUa
LDT7FO7VOm/Z14jMHOnIKl3qKVdCMNSftbsRxCsby30ozRldpomOtD92ca6Y/fHn
kN6uBmm4KnnopDcptb6NjhSxbWPdkQul//Gh8/VMtSvMrhgxnmT7ZVlbedFVB4ES
SMdHUxFqoOnx7AN6jPucewf5EfvswreJ1PXeGoHnrfL6PLugNKaKX78dkQb8tizK
xktkgJtEQuu2eziEGnn3Cn8J5+McVydruxcRnlcvkgQOtNThxrzxynEpdfykv8gW
vbdXbtDLkRy2sNAIQhREPM5uQXW63ycG5XZNLakf6UPTH1oj+JBkey1O9CHRDyJ1
74gluNK8Bthj587yRiN813G0PnA47ibkBGuva/dFP8Hyf+xbehHk7HVoqmfg/hwt
9agZkOiQ41VEEAjx/r2eM/pMJ0l80hDnEY/JFXfaeuUAU4Ma70KQwf7FSjdNe+ZT
++VTYsJt33uERnLJNbplJJ9PxjNw5uYihPASsRiN4WfPN71Wqwg6Heizh8XN2ZQF
vcfu2nUHfFy5WUuaFVpMM3BkbnfFNiHMh5RiDVzmT9VAeRcpgrDfOvWMNGhyDh9l
3CgyF7x1ZnOwYSphbYfx9Rky4KjazM7ryK0pCPM+G3/XjHbq19+S0mHY3m6oNr24
nQ5wPPU8E9pOgm/OavUj2jPm+rwNqivYqw5X4T2JyrRcYC0lY53iyv3GY/cZz3wU
jgTSEkZt88BJEgnv1gAjbIrYVdfoYQAmuZ5HjRFtP0nvhBDzmJgr/wf16eTvXDn6
X0HJLDaW846IJ1L/uIf1Z4dPH4KbpWpUKcpluQprtXMZ7Z9bfMK0b10IdUiGeLAH
Dor+Fm3znhip3YNmQ4C0X8szPbIw7hoSzgX7kvzmdElfxNHeTtr0qs2wBaS2O37M
vPd34tCNtSsQkkqQIoOZ1s7lDhY9Us/31APQc/hmToozgst6Ls7sCrSRBytrkkZe
oyPY2RyM2uMoCg9ntloJreRvYO6UYZuP5AoGEPAFuDSjbBswoISJlAy2ImSR+PoG
cJWrXT+f1Bdbpu4BZi/AcjMfr4mZ63Ev7/Fko2WWKVK0FXymwZvXPpYeMFF+66jJ
35bDf3GKB12KWqlTEJ5IoKBnEReCjxUxsXpJSl+IpP6D8gB1mBBujn9s/CRQT/tk
8KFi4680bcEETQ8OaMxEjYex5S7PZ8aSaSuf1CDPWqNQdqRAzT3eIp+5MkKCUYzK
BwXsBppxtN+Q7DXSopHKP8IwKONWaiTRDVSn96XUEwARf1aDE5os6Ic0d1gcMGbS
IbkSxIy1QnV//H6RfG+1WLyXDlMCMBY8110Eb24eJ6QH/ZZTgccQsO73ncKlxciw
hiE2IYXnuGKeoIFKvEbGtv8D5ZsVK483g4m3gRNV1xu8pRIHNsH7R5K0FCZ1glDl
aXX3oM8tQU/efGms0GGcT9qy9zP8p3BcUe0d69wbkUN6S4Z8t8T0odNc5KRprzxJ
XgP9dRt3UTdtB3Ibp8jgNoK2qjDaucj8OtDO52K97GbkEZEGZueVVno9rmtD0dIu
TIyY6tovnzejhNPuiB9IJixKwxIIH2U01Mu0fkiO+gv4NGk9O5WMpFoGAfYw6per
h7A6nZ5SYmomO+6KRQ+WA8L5YnlM9GLtqAjxdbAfwPACr3ZCCH8dwbBorcGhhjtO
ykVXlpy8KV7boDvnslZ394CNvBkWegfa8wupWXmmgunfO3a2Z1r6VrU57ocowc4D
PVOeY1oHKFzW4pUSLXPEHWrstzGIT3JqlB6CQuxlXo30HhkixE3buxGRRkZk++QW
8/L21uYfcxKRLTPPAXg49yd7o73FBHQ2iC3pgqhOMs91zBNd9Y/ei8hp2K1tjqHz
PtTUoOANka02HG0vhp1wKGU6YpnYp2l6AEpt2WdexCkiFAnnwtXqLVaEiz1OysT/
x4PfiF4MIaWzCcyY60SxhcbiXfFJKFivr0EMVoRMzwIfTcezxK3KldtfyyGgZkT3
d9wvNe2HN03wZksLNKHedzHkOthlJ1jLjie6lL9JpjelWcezzSeG4Gy9PKwhF41h
ukY03rEDzRdRehkHqSR3HpPIQI07UPAcYilthYxb5sECNYgLqWYYACEBVbE0d9Af
lh+QojRTH85S5NHMfFGSYEKsfgPtQIIi9VCA64csWyWwnbWUlPuARoOArkv6JHQe
kMKC5oVYjnJYBeZpJqW3WmP7HbTpghl6S2N8ACWWQVpZLDWVB2YdFNprffyxZUc6
hWRSFzoiKSst2RaUOP+IX/CdBSMzHK3yQt4zLuQnsYU62F1HQhUzLaPvWdR099AT
u0AAe404hGdGtzTTnuATaj9cZCMoqvZihOoqSlZ79J8vsF17GcBEv+GiaKTgxKvq
oxom7GANoS7O2oJzGeWZ6Ys34pUTo9SWGbFcbSdPR6Qj7uImybJPl8PVgWbFd84X
ejpJVm4aKmUYdc8o4Se54QXXgaQc2ZWxWJJ3RZ3i9TO/SD2kMpD5im8lNRXl+chZ
Qv6FFkl/l4kx5NPLHaLNlJtTMxkB+ERvRLDsYPlp6Ddf4rTxcDsbAHTj1bNra9oh
sIvFMYt7v5M/Il/Kt7HOi846NbpGTVGDPUl24AcrA/BdwHe5lJYtbDmfi9kLr+em
TI1vYj3X+mIQ8g1LO7o7Nx16sWcOFfO1p03UhkZybRrN8tO9LSwlWm/3ZylGiTVA
Rwsm2TTb9kAP2J+ahR59Bj0adGX0b3DBVmUcE8drsS2EYJmsEZ5+wwcjIGtGvmCk
pewUeWt2R2+GQMjVu3UOdzMJqATXhAgyw8lO6RBY9pcaJo6Y90Vikfm5v3EeZV1C
KBkguNW89Al3FgnM6Afo/oIueA4rxZKdGqNlfNnncdX96MJP6kt60wlfgKazSCaa
f8TY4r9cVu9s0l5p0uhxyQO593Up5bDnSLANCPYJU7EiydU6wC077ldNhANkIbxQ
PvnKQWWlzDJJUHl4Ni89FGtU3pAA1O6OS/Jy/0PwFHgHUSHEXv9PqPZMR0GPcLmF
5TM4kjJCPTh6IAJPz5i9jcjesALkIwtE1CZwK2Mqotf85xgUP4Riv9kvFpYYAXa0
dKMrChQWMmOK2TdrTrGlCHT6SueUy+QX/wL2x5U578xSlFYig7Z1pDUwEJ9yL+6z
3xkVe1W/hOdEYqrvtspj2GAP6ofzU4Zy1jVFoNt9E/Ew8bHLwjXViUDb371Gp8QV
UaGXJEieFrLwu8AzSoSCHTC27i+kh9+4hunjpWbp0loBqsEke+mUxUUlmgwVONXj
Tc0o3hpwhXLs+gDpMeyEB4rRSFOgb/bDSKo4l2NYMhp49WzqAhFDgyC72TxhlaPx
zbBDwCgFhylcPCskE8tpjI2wAJ6KbCwM7h90LPR1CaiDgODPB57NcxOfc0DvgQwf
of5hKIDhIQBk19kMP+oFQAweFak8EcFEs5csVAko+tR8/TvAhE2NCZrnpOIe7aLh
4Eb6A5QEJ0G0gBoMdBkf/0sClRxibGG+dSr5PUCGYWtywxIbRTtfJxgVyMGPORAZ
Mf9rabmjxbL4eu1I/gv76G4nC3jEhTmt6UJVA7EH/f9jqyQ6PIT+iptZZUONd4NR
6RkmQIc8IJVt9p2J7V1fOY7qh4pi7J/jkkodynGQKrbLb1U8tp3Adj3fs6B81bcw
mXSR8j8+/CS8IhRATE/8b+xyp43AmfQoq7IUBUVrIlMLOfJyptnMOmYJIY5ibvsu
MMtQZdWi71Vgh+7Yz4R+vVbcjiitk0r80V375B6FKRcLCKSvyab7qQBAMN5ixiJn
+mY/BWS/vge1yDM6MIibvn01dFW827GYaZyRUoviVyWrtAon75wy9uY06LH4gFui
sDjIaTxyy+7GIhvCHo0qvVY3OuzxSj8vefe8dW7NN/iZJMIapGUablPArgjjhS0a
60Q00dE3GQSIecrrstajUMMofBRVVBen7FcPndYRfHwTSim0nleZpokn9Gf5Sh8h
7DLJwsNNqPwhfnCMSVrjoPa0zW38+zKHYg2M5e7kLbziuUaXzKa/5BxKL3AK+WnW
PdpmC8hxnyO/hfpAVJKWGrHxMiawvdlA8Gh76kU6PDuekNHxSNsr6poo+DYY7R66
tfmQVNv/AwPxP31fAu28kuxFKE6177TUmKOXnI+G2V6L8AFcyRBx71eN6ihrLw5X
r1H7Rk5xpj1F9xFuvkSh/0qpFYO6PpxvjHN3VKjokBDnY3cCfke0L7YHsrm6tUi/
u8AwTYNWS0e2VJLfArGlDhTY3yXXi5BhhRyuP2piVJukda6VGKV7AdQdFvneqFsl
3hcwiJfQwiEJn12pry+vO8YvrgrpJYQwm3geKK3nMf7Yhzo4OlTa8sXS6xy5iVmd
VfvKM7X1m19di8ekMXQLQPbsTQ3N/X2t91hVh702b35XV9Yw6U+u+QNDqnYMZBmI
dT3X7+iDEnENwi+uXYetGt/IPLbIuIvW1NQMHT5W2PfYLMZmmnw1zLLcWemngvsn
Be3z/JueJ1NAcfNlQoCTqjnu6CL+SaAjR+YdtYqLPsJnlDVtoqeLNLRgzpUnDv+j
K/oo88QX6xK6Sn6oq5u6CA2pqx1kq4jpDAk9ToRFbo8GJZs7w42J5DOwpfLcVrGG
Lr5p2Fahx3Y5YuYVWgU4QhWwYXJML/8aW6B2KqhKAbR+sPLiWjsXF1YggRuX92BS
1Y1YL6d1x/ZVnrBK5c84IFbr6TolHhCaB/C1H45QCtxPJO7Mj0Mzs8OrxARTSj9Q
RRwK/U4iKR4pM3ijJEMVEuSC1uEXFKVbhlW7l1QHbT/HvG3as+iLEXx4W0GfPTaF
eidEaGn7SVOV+MdOCXXChf52EmZ5qhhoUOhslhlc7vBNNEA7k1Q5IadURvPwgHjJ
0jOUCfa7wyUvVY4iGwTKTvKNr7jbM2ZQhsy9NDM89rYjkPTE/S/WK7FOeO9ShC8C
de2R91PZroBmfWdiG+etvj5keSQ0xGKRW5TN6EvB4g0pmojwMTYavI3kVen0Dsh7
REOMiDP/TtITlsN4U28jzQv841OCUsXn5LmE7z/Ji3AmFJhSvRF6eMmlKeS4GKkS
kt3BJhDMpmso6FcDXXkFyGLCMW/E3AOlLFeyQC0f5la8qsX7gFIz6Ng0ui6/otCi
7O16q+D9tkn+jVlG3UAgCxvfiMixzUamTe/1o6ATtUJZ3DCeUQ88BM7m8ThMaF91
d4Udbc7fqmhjPXMd+x5NJSOMoF1kVOM2ahlc70WghIXG2a/zwi0DBnmaPJM7fTM3
e0omKgfkbnxumAzLB+IsxrQsqIaqKgGMx/31XNkUx5Jl0GvlEEpx4bY2TwVHNg6z
F+NmZ82TEIJYaqnuGE1AZMM9bMMStAeI+Eaw6SmZbylyZkPXvVNGDALrWG6ElXXV
0vUylIYSKJx8Nes58g2fp1umrcSzKw+f5dP+jEoJLHNZU0p+q3+bzngiAWPpidLe
YaaCAZdSNnQHTMyhmM9hdF4ttl5NEBtrKGZuCllQkC7icY0DhiNamMBrJsq0pCq7
jYX12eFtvUTiam/aVrvoVjHtG28V9lJF9ebw88EDQZsddvYoTlv8sezCbC5LkT4m
oLeMy45Kk8wacnFZ3VucXhfRYEEqKu3wCpVdOClBzxey67fLKkkKDMi9SWh4Dh16
T9NS8LaFINKV3WqLfcvtuzKS3cOTXCRd8UMM4zAQMGNk9jh3ROh/d4xTtETV0W3t
Y+HAWI4qYmGBkA8uSEVNJYkt9XpFIj5mMSSLjPHov585Usnk1zyNze5Tz1NAdoGN
arhVrG52qczrxesmAPKlDZEMg2j01JTMHa/hsFAKyKsg2hn6lAS4WkC5KrHLWcgV
40Bpxsp1p9YIUBXtqJaMzpDXij1BA5Dawv+EDbYvUEOlStONbHqDj8i10Ce9OV5O
+dssbOaeGogz0YlwF8FmA3leDP7fwqpJPJs3nfLHiK2z57X3n0yQv0lA0ziMR38r
phmO1TQMNH3ahypUCsOteoLE9RXy/TZgGr6j+aZjJp/8V75V86+ZO3b80h3Qede3
rA0hKCZiJBey8edpXEOBkAOvY+JFtfrUIacXTZAkl8b5vvQsyhEGDDxZORYUGRNS
OB3XXRk4woHSor4I5F/QSAbBPfmOlM4WPZzpJo0NCvjAQluXF83bARV9HvlEaqDN
PiO3/ocNSfm7Qki8GTlWB2Kuh47540TNllZqdnNHn948uFxw7VmZn34fkk9HXm1T
3pAmZFIl4uDbj3ChqXoiTVXxSk+c0Ih9UrggP1thFe5zJ2a9wv8SnKVVR5mi1ItV
p6zladTFwikhFILHpgVl7CCgUHk8yyqOD5ET4/VyFyiN96DsXweJeiJzodE30XDS
QI2mAN890YIUjTKa1SJM55cCn3pVIcV7pYJFdc3rISmI+nMth0ln77gdcRxStz39
yVONaL6ZAq7sSwkd8MGcwN+USxF2XCLQn4y5rCuAW+notIS3ZTr/HRmB6SkpxA3K
Mhr0+vJWVxWEFZE2XVsF1rdSGDkEG5XrEecHAvmgEcEISI3uPUJTa/jMn1inJGdH
3tz9G0gTeL7UIrtSy7unby4GKOhFI6hlSL1hR0MuzJEGS3g5VED25aA298JbPICj
ogH+j79Li83LcA6/ZjEnnDt46WQ3kVchyrzh2kJ51JNSChR1ZvqV+iuwiMDfu4UP
KBtf0t+TbvDW03MdaIWIAixmSrT7ehOWxpWNDPHZ3UxPIP/qlXxsDUAvZW3TUZAf
5aPVDc5JN19zdUoS+cPF0/YULFyLnX97GNipWex0BlIhMK9dcFRpXYnXLLnINpyU
2aY5aW9PviSTjPt8m48EzvM7kN+oPDFR6t/Kv+/zBV5shi1Sfd3FKY92Y9MJdowT
/4U/1L04c8F5k40NUSIswQgeynLRnL/pTRgn+wL3QgutqNlKQ5iCqNulOCYGrJVu
P/1KKKf20JainkE9+PFGKBsupZZX4bL7HH4mkO3+rfvzbYLjqadkCLzCMrD35ggv
KPDr2AXXEn5EpfO9M5NqgWb2matg/frWp6BDueTjKskVpxY8W/HHoFI59hgdT7Pj
qFCTT3zNVBNRd7EStyk5J/JlzcHa2nHecOWJwH62zfx3b/0xPXiJUQlyJteHmExT
7AIuugDCbToahZ+eLiVDkXVqeY4jpl034PMTwOyiYjU9tVFXfZOZVN/lgFFtNPUc
2+nFcYh7sW0m3cu4SSN9YXjzpBkt/3JK5ULRRKlvj+DVEe9Ux/vZ2RaCJg+M0Eza
V5YE0q5kvebsgdGrRCfJDRsouIpoCZOqDfm6LYxTkwXf9WpLuc/22W8z3gqFsnbS
+DFz0aqk5QNvltO713KwyfiNcjBWa9Xzx/FVmIiwlXWnd6/WVSRPRSdBYvV4wX8+
h0lsW91uvqpNfISFP7nX//j8S3DiQ4qJLCGzr/qNZ0evHu2jhltfH2RMN5uY7KST
ueG+4A5qIYOQsaQmqA/bV8BW8xfSfbWx/j/oax2wdvt7e62QWFuVA/73EhrYF0Vs
FSpxceTOJBRtU8D05xDlkangC1pO2xJbQ1gv1d7kPi4JJOLCyTY3f6julwC+Scwd
Is5TFxdEVkLmcN0Rjp8wVkgEJSmnmVOL6RxpMLjqDGn4w7yF1hc6Tlq9s74OwFGg
MfxkOb8oVG0tJZ9ixCRmLzXvVZ4KI19HA29eTER+Kptx1ORbwxDL7mz/eShSRG2G
5uH+eTaJU9GUyZhVociyGE6mOtSz4jUdnNs7ItI2YXpGwn/bWFps8WunZbOZfKKy
1am2w7CwSkvZy0CSwtkMYRdn1SKTwXcEJWHca4mHv0i7bUm6YVSXVh+goNP0Q2cC
n9iWmJk1jWC67xcVQTJsAE9uUX9fwELBZ6FQGC/ElUmcANZvnbpMrSg3OX3Xlmdc
4u3J0hhPBoOewAhJkC3ljEfOqqjGK7ApJVThqF6BZMuG/6DeBJHgfXL04LpEbHdf
gTMrtZV3VYxuHPErX1unldULaPeGMwK/gpIke3Iu8mYt+ED+OoQ4bt7e5O6v4F6T
KKjYPtLnik8zV0WXzdnWB7VcA92kJZpnO3MHWH8VZgy2RRZHJCR83o9BxxSccVLN
lawvwSdNJcR2P6PHURJeZxSnJph+mAGQBA5nC8P23Yw2IlAkRlGvlAWA7zeKck7R
f6jrdCUqR1SvaGs2qI+OgKk72Bu2t4B/gubqP94a2IB8sG9mbp/DiU1j6UoBRgAC
myyLSxp4YQ5G9v4+pKPxdwMBBT5EM707G3v1d/U2vzfHdBSvwbY+eNIVbUWLPWQM
7Pfw33CWTh0NwNEsqpnLyb9QcPMh7Y8CZRlGSGs/YExRQnZyadxI+lk9Yrgl86Mk
Pz9P4sN0Yuv7rEWoS/XaEJDxUlNeGrJ+zUVxmJ4qRAKfqHFkLUZtAMVEGmDJLX/5
t8qNkio1hlMpluJZ6CXLjwrhnyeAm5lpFq1j7ljhna6vTZbF3e+Y/Yyj+mbtzHVi
DmAtCqGjJg7mb552zh7OZ8XiEVtrUHtzgUiTOWBPd9+fsol2PqdhS01qRzfQOLp4
WRT4QiLIuQ8XEkE5UsE4iY6yzMagSKr3DpP26Q3qbs9OS6mlj4hU3EUQ1cps7j0+
2rZBSM4ax5yT++ZudCeotE//UkPNDFI8LDXpsxByzmDBKJVbTccDI58TQONgHcuA
tJ5LFSwbrECTevDIASWNdV177MvEcYQi6/FVWCdaHZq6w1yBVzXpGP27cC9scP2h
/obbcSlaDMvaggEFEnIgw90kv6XvAkn/+adHS1Agsb0KsL8udbAYcZr8JYZF6SDB
vxoJjUQvlyZ8xZuxTC8ASEx2Zwja1Cf0k4FZm4f7Iph8cUKLGAUM0SzfjZS2hNP/
fUWQ7Hh9Hcw11QrMrEp+v5RYyiIPCtmcTEeeDYU2um2rUQ2eB26HTJcEFhnpfZrt
zHlddKAOBRqtA4ZWajNlvVq9AaWvrlLxneclrIydMbKtiDyTn41kEezmZfKYB7Ug
Mp542kZDrbyxUox2YybU3rHJ5WAA/pb0TrBcrwCYVB4Atm6Ojz7SxHjw4/K+xP44
JgKt3P4376qUwd6NLHeJbmYXckEQr5KT42zF+a/uZNq3DHvokW3fIkIsTKaLxYyI
sxBzx8plc+TTWZ2LNoytNP/jinSRQpfM3v+YmjHeCiIZ4bFSpA9suNT/Vy/YyZZD
Uii/7VIX91oYs8o4wtEmlenAqB0EVqLc0UYs3znMvJI9g10GDGtoC9axJocaB82N
54RIJm7exL0rSZBXyXp9TBeCUN//VNDL+7SGDywLXyTFk8cxKuKmYD7jVZxQ5nmp
QxHu4omUTx8lIn/N54NO9UbiKft23YgMRctuSwYTdl6fhI5+osFGuWLYB8383Aqd
72qD0cKlZvv7sObEDvlYOZ5Q+OewB/D86tzhObQmdTV5xNsqSX8+ig/uiA/yJ0p6
2v7Yj4t4lXvzPysbH4BKuz/BcKHXu6mNvq0Y8nB+PeL0u3XrmLrVoxFmi5o998XD
tsRsaWefhkVezEjn59z3My1QfD6i19MDP/NbYJlKIOhrxXT+GzBSw0TUvLoxzAe5
m4HyiJKt4EPJv2AjsW7bm+7wCYvgTRULFmmrOngIqwby5o3dQmKHiLCXU0Ri7yET
AmvvJPKUR46tabcMlZfqRBwL9YWKRdaI8ZSYRFHKAMaCXMplkRQtRMz2E6h25Hus
WL0R4kdg0iJ7xq437d8yrdLT/H2WOa6kbdIcc4Rw/kKVnpEUjvqDnfdeU2imfvoG
DwiZ8tA5atdpWW4BgTioGcJoSnF7SPDogqqA9lXd2C5EtK7MvKVYDnzNF7SjY4sj
cc5iS6UBoCkg8bejZECYkJZ2fWk44gWDHXw4SCuakg7S0rZAhGS78pATOAQwAdXg
QU3WqFL58P4fRZQmE7gDjH1n8RPYYIag3J8W0kn0yxZ1OP9MM8SWu8IJTVhR9TrJ
YZE278UKBTTtMVNncMvPOJb2SLAqwAmYMECdE5+vOKOJoiMlJAzFitxUBOEzSPmw
AMeEwd/CGijgyMx8+6ahamJ+QXZlt+UQSuKfr57qXvlHWukWHMS6xFo4kkkwi/Qv
arNUTgPBs3v+cLROV5iNoTnPq6omsblzHMCxHHJER6J/6LAgcfUbTnkysLceFBvz
lLFCALZ49M2kidOxlZK6EWUiwPsGJjvSKfdwlF2J5UZwuvLMw9A8tAvCZQ3tKt6H
lVetD7akJ46cLHJTslxNqz2TAOXezmXnPsQOSA9rkuii2ApCiU2HYgGN/VdgTOIr
GXkv81NnakTEzjDKLIxJ7RnPPbdiI79uYauDtQUOcvOs/O3hdmx3U2NgfrrySots
wq43/lLpqdCgaRzg0LI50Urqgp1RTC6BUKnw9hOMfAzb14dKfmMGtAyHtn3917lr
Z8kzunPKUll2p9/1DZKsRwwVRKRboR/yhafJdIhWQraSC1mL8vxbERmScYextWK5
D3t13oAEAgCOmVg7RkJ+FN3dVty/gMC/ArmIUChY6CpxJxL9VTYHXng/xQRe9WdJ
kVxlybeMA2iRh0SH0qN5rAk+W3X4JM0QkFZrAN9MJwi/aUbHRC9uCBDNEDulx1bc
7a05yQwKANHj2xu9h9NP3UGA37pqu0mwr94OSqfaE6ulWQrhuIBoH9Elo8QRKiN6
EZ+bg5y+lQ6E5xlYQyJJyZDIcykbJ8XtyxL8WTJLNpt+Rls2ophPYkFDXKX021WX
PzhsoYSKfsB/9NBfNGdgXrvmOHkICAYohMhUSC9CqHYxTR7WkAUfRYHPtfOBvLqc
KVouxuC147LomoPmCcXa4QGFZl2sp6glvC9XkMdTv7pD+7/frNpOwyxnxn5PVQUx
3b44u1dsEVYJzYofTFfk0g7sDSaWQM0oWWp17zvYqu7rCcVeeYhqjl90bIedeqyn
6iL3CGtiNe+kBQn28KUvwJvuulz4zt1KK+DB6bIUublTd3WWKsj1kegodOSOSD/I
wmnQHA7gcHWs2aoDZESreu+KPeJbthdJwLPFgZRwOP1mRzhR4THM6NUmX5S9Qmk6
sFX71ueWw5OizhSF9XtVq4ghemSudmGy88o2DNrmPfOAStaYAREMRFFKoFCTVQq+
Mbbi044GsR6wF7qUtRPhBVFHpNu+EmhZxBRN7reM4RG2B8OWm3bxiAeL8b023V8F
WelneBO7U4NZq878yeMpPIuxWZrUYt/4ljwEyCi+n9VNfjMIts7gn1oc6fJ1fqXe
ecFt8x8kaNY3CsKsYbRnqiqliEcxNRLkb9PoeKU7ZB3ZI8On1MJuxpN0zChdBeQL
FIKcJ1FjZN4ybObUCT1mZs3hrBrRUb2OHCoAbdioTDfhHTHILapSFw0RVYDMGke+
1opb/Nh26xm1oxRJEwl5sbG/njvLL6lQC5O8GpnFh+mPwnbxZz2LkR8vNKg1eZJX
lOsljgi4CKgDzTFGWZwL10BW+fMu/FNFXTht1Jo8Yo68jNs1YM/zeajrurZg6OME
NM4/dRjJ5qgVV48G7b/YmuQXP8FaeMRNAAUO9kqDh7CPpAFUHZg1A6c0OyiKpguh
UbWP0NBPkItzUqDUwM7DCDSV1a8d5Zd5NS4yRJCvj/iUswmTypaeRXEAEuP5+ryL
P48crSJZrLQ4a2BSrhXvdeojhkAdIyXenxJIWe2PUAIwgqjl5aTkYejpQgKXiQb0
z54oY1CcpoTZLKMRAEHXadoPuDsO9kcK7Pr9eKmoRaKjc7cm0y+RRJYLJsQkEim8
T2q7K05XXKmSt4niHlHW0DfUv2/EWMgIWcprHTcVCqgjhD9anuZAgujAYW8Fm/6G
alxQDsMjqoqIzqb7T2vqg9ERrKNpjO/v8v6TyfwfXulcjc1+APQdTgJ+c6pfrT2V
y2E8H37C8Zksz/JTI4fbte1eiFt1Yo8RZX5D1em4roQqzI6RSmcQHCPWsEbYNyYx
bbB+XhSFKRwvCZuxvs1CpQXTWLvq6HxDnFvzT0CQtjjLfPUIupkoHS/6t0K4Jgdx
7ElOprHggYdAPQ0WQ5OG7IgD5LJ3NgCkPqWND5xC0Gx6Qw1MgVebRrB5hkL2DGP/
4vn/yh1AQKHk4w+XxVJyUpc4gohLEtw3rpPiWpkYT2qWBhyUF8UQ2hOWUlyu+mjY
yS4eycEjCP27vmhgBuFIbBvRXWqF1ePEPUop3gdYRCn+vLeGcYFdOq4qRHJUkfIf
EQKJLKWt191/GNVlHKauu3WJXD6e8I2B0X/67TU2uK0sNZdCYBl/HPzuHy+djqLN
/8u8EVUi8NNQUvE9x5kcurmfC4hX0GXbMKTdIMFRhTjTzS46277Xp+f/n/nDn23v
a1iQjGoxQUTTLs8OblYVfjnHJnvI2A9iAFSezY8LKMuDGZTuS9sKMBTxiPP5N9Ri
RwS0MA9Qe5CvDJcBNnEvw0ikqSudvHq6JLtXZbj5SBOP5H9qD12vR9doPPAv8RjZ
L+Cbd9rxtwTsx3uxhVkShQmTmcF97fh92Y3XP0RsPYlV3ztjaaCX8FFZJQN0Cpuq
VDqTTXYwu+NaIbGglvmm++XNmyyPUv4VwRSP4QdIfGp4W5+2K4iLKaGcHaO3EeB2
rS98aNHD9NS9jieTuBkO2K56ERCq+0lUwdF5ZoShNo5VkQm9XYwACgoio8GZw5br
U91N670pBg1gHaquO/pEUznx7RujKKDnB0+ZJMwWiRZq0/v6G6tXhQSdIGR+PApA
nSCHdMJgGNTMIrQNSs+OW68XA0b74p9YjeX3hq1yf6sB2UodVUkeo8pDWUPXITay
GCHRxMS+t8rqsR9bjkFV7UfMmr15KXOKt/p3yqbX6xGu7oDfpxXpKATYtWnPaydW
uaCaAzA9gSICqdgDjCnJoBZFEofKomoBcTecPhjnBb5OW3Y/LKaxbhh4jx8xnyuA
0/0drJWv3xU41VSlMkIZhLk6ZKyBpeeIUYo/csh6PERN6KTIGcDWxFz5X06VUGVH
A+3eWjyVcelCEamJ9tdUB3hLNoZ1u+Zy9HJAyXj2G9e8cRc575Ktk2sYgx0q/rc7
dwnVhY2oX3trnfMl0ykYb8yK2L4MGJCaMzlnxw9QGlxb65ePuVuqYNF2NX96ahnM
gsVAKupROiWpBRvnTKqgyg2IzAt9us7hlApSswTMo29H9itWZc6IY3btbwptX2bV
qumO98pzocCyCrxZP4yjC3Vyqa3Fu0Vjgr5KihuSIbcmU5V36yK8AZOHYaT2IDjo
CMC+FB0j4Pj487E5gvXGQS/v7wDpYoXMAwHrEB8QH1wF3cgMOsITehwoptSt6w1l
mShNWjViVUpYFOU5rMeSTuBYXzfVdWHVZNwGipt9drxygBKX7kyil6qvU+Uys7hc
t3W+3ZNWIZkJ1tA6mmVp3LZoPrIA7vAzSUPpwSmzEn5rN6wPJHpjkU/9n2juIH8q
SZgo5P9XugQzg4MlGkdXz1uow1ZzYFP3P3hGK9+kt2igfDXJKqlViOG5wGmAVi9j
jR3fFbjW+B7u05JVyf7ZkbaktUlqiqrQLjWjezXzGuc0M3zpcUCadDAKz1JNgT6U
glCH/BLr1rmsLr1OipyTGMfWHKl+tGztEf7HlGju5l4u6QeKAYp9OpkQ8d6eZyT0
2hAzP5hNggIReP2wgCkYBDfjxlDsPWq5rdq+SdUKQoGH/Zfv90fyoyexBv2eTALv
G38/M9wQFAuoYyCRAsG6YXBm6qhF/CULxqfp4Iws67x2s/gwMcC5I3fKqSGpBBkp
CuWfC8uBTOFtyfVGZ2YHWF4gFSKrLgw1fkHaCRUIPIk8/RUm1zS+XQ4rHBPGliEq
QGeE/O0wJ3G4fKLStlqt08sqY9tHJHX12heLgtUbBV7ApAKQaCM/cqUPHzMEF+su
jvG+BV7iqaZh45h/jRCaX6jHCvHiOXWQ5u/xHO0t3wOQvjy6OMZdkrKuyzSw7E1P
rG+3xPk4JxaC+eBHJEb1PPFpoFH6SAFZ71PZgb1iFpGQ2Goat/9vPuuvmXjaQJTb
luZzRkb1nWgyTOdiUqx4XrctVvAsNcuPjY58cKIstHurgQAbb5xyuSIvvDhCrhi8
xi2JdrmEoDACpuHWCHa3aWGntPEocw+4Ffu0Bh5ah++0dXoWuAARBx9QapsqTP1k
hFW+gh5v2AZy8InMhVubf2hMRIZmqSzlP9n9+WoiPeiS0hUnmbnmEcnsqwzVhCW6
8rFiZiMJ5f+MOTVzSsZ0GvaG/ZlEqTtRZoidbW3J6CLQUsQBObiJzHrY3kGF813S
1wzSrVo8lHjj0HETO6/7aNOAA/jnGtkwSkOt5tjmeZ1jLgPBlH8QQWYHteJ3783n
c3DHmf+de1kC3LxzzCH6zWZsgCaJrq8KNE5Es2FeZjr8OpVp9+dULMkA6ho+4pdd
0Y3rz+aUV3qGb/zNeCqOrGZsduAnSeu90uGKBZmg+gDl+xg7wVGZFSoousaxBUK0
CoCY2dbwBl7cLisbjoywQWJowxq1yeRQSxq6mYmZbbPThPh9tFvi2qxK87hQDATH
zS15iU/215K22+cCtXHzbb5oZ65IoZvPwayU/EnxSpxsa3svtk8I33UKF24PmQj0
AMLWaP7MdOkWp2MlyGvmTJOgzaZPeJxlQuX1c9UYBTh/Yachos6Vz244g/cpm69J
C0C0kq/qj9bnidMObXwz/gsk7A/r1BDv64avrthNXBRsGnsSMRO77YhNl5qOE3l2
C470OU07AfoBvYDsv4ncP7hs92oDIuWBEQSnG4ClbgrG9LbxqrQHGPb7EW55Tg/f
3SwmrzUHZeEcQvFNxFL1JvLU4t5qNsv/kklXiUwyFOOntRMVfebQeIH5k9lZ4aVr
QJk0kIjTfxmMKaA7MGq1WFYyF/bAmQNl/4xAB7LpDlVRvINNWfw9CGWwJpfGo90b
7Ey/AVWuuJFHsglA4OC9qq6UOZG28By6kzaEGix3U4euM+1Zg4wjWqHcWaRj31Xz
ReFYzpGRjENtfCZTLkh6fwYZ/xQl5uz0ROnTHL/DXmLPJ0yyuqcMC/8GVfKoi/1h
J5LWXTDA7EU8tWOgQADrldthSIhZd858P1GsNfCEVQ3Yrv+gP0nl133VCUAoDnPb
zf3FM/GVUMUtbrU8xslXduMubWaaqgPXGmivGCrxIAiqi2ES4CSy5x/AegPeDwqn
kMm/BDfufrwmD5B85XDdFhoxTq1Y5j81IlrQI47VaCdByZyCeeBk/dVgAVdC1bki
vnP3BXrZZPxZpUde6rkh3AGBy/w3FOExpT6LUWl7639wyFuVi+x3UmNk4mvlvS/p
XEXRDnbx5x/0X0XZ9D7EU5WmxA2XJCGVC3QmMP3yRCw4KNxvAptFZMr0prn7t6uR
yL1V2W0syLLFVHCMgqp2xavpc8s99OsXTZfDQCzJ6S0E789II4aaotK28Ke7V03k
1Ho9RKNLJF4Zpjbw45BkNbbGSXWSIxoK2r/zdxDQ0lSD3+vO7so2OWcxjSTVIh5w
7drS7MnEZ763jhQfIU+z7FBjsGN35iwbeiNSHhjn8MEIrdFMEuwM4ANj191udHCk
FQDypb/AX/n99EGFih8H2io8eQXwonQq5gOb8H/VCRbfCnMrHEDiTUZEqWm5Vo7i
8qW9vl+m0JRFPwFo499GVP18LOBCR76zqbb6xLtnrOm1cmGaMV/IWaMLrSo3k7bH
lsjDmymg0mxuPczua2FncUd4UkmXnRcUq4z+OKbM96TTYDDaW2A1DGKwSY7/QlTC
wkIT6ianxPHCI9+nMKOeO2c4gsEdhBboqBT6DqB8iuMf+1ALgaaAyzgleBF2E7Q4
7LHaQQRB6TdFLs/6W5jiqFQ+3q4xNZpYvjfwRA/l/J0pMG3X2XPniwsH+SrWHNc7
5FQIYg3mwOYvjiYF+K+W23kqtUXUb9QpkUecPCdwkFhCMsfd59PRMJnzQN6/x5Bm
3W0PQfkrF87Cb1R+dFeFAWUuPfMTwXH0eSDJO5gNTLMgm82H77BMlMqSgWJXK/v4
vUaoNVk7I8xa0pxLUDeI88WzZCQtRKadYHbLoHyqe0flbS4qQ5FC+fQCp0cEFcCu
KBunAe2r05uahDhJdJcuEoBdmnGWt6McO22rKIq3TbW5JW/eWJuTIJKymHXMCLRi
ttyCcwBabFPCU+Lwf5ZYpulU32KG2m1wmvvjiQUyjArERvGPRKz72Ugvn+8QBDV6
T6SnPAagbzlTl4+L0SzlkbN7DCYbX98WXViil6bfayspBFHtsfGtk2nomQFYeMK9
UMRBjiHn+PmJI7Z5ZRWYK3gMsWtjvReLm5LVqawkTEQg8a3TpxTzGdt+gzu5QTTM
Z4PNXsiggAr6qlDO+ZkUyZjk0I8dPYkTMteyeIDn6isn4hvvt0a8J5Bx6msuPG8J
bdpybGm2hE9Vf+FlT0QZQ37aPXHb+pfECPv3+FRdhp5g/w5r9/4N4M3R6if2Ue8g
2FVgEb+4Eayyc1m0rGlQCNC3RaEYDQlsHuXrzPGk/QgP89F2wAeOCzXqwaLKEihC
pAMuOIDN16TGQYeueT/cAfzQVOI1KsIKfhhjLSW2Kn32K6h1JLq7VVaZwA8fFre/
kTIeaLp0k4f7L26l2KiHWaH2Ud0/0g+h0ytZW013JK5JBtrJGmYvE9UDUn+5QhQ8
KmnxqXCPf48JVs8QARbcNwO+ayyCz7lbHZI/xl1zLh3EdoBF5IFjRDAFuXsVKDsZ
oki1i3czKCLcWpoHIdeNCErEmmPJw1xtRPWMtQ4LKHbx/Y+DTT9kUt88N4Y1BDP7
la/ntrWvbiJX96Qw+61xljv9Qgnm9Bucsr4ZUOEeJSkrqUArdThY+xxnPNciNlc8
9tDzUlXxn+xlynNhbL+IbaN6XP7WgoGr9RL5RbnDgbAzk73a9NV2sgNNwgKtyHP4
VWvFGg9RW7Pp28zt1YGnRf8qRS9AKqej7N4pMpFmWKXooJPUPauX+1MtmOQYNg8q
M4MdPdI1AyLdPIWM2EYEWPXmnoZ6nlKrP72WtTYTHQl5q2JUlSclMiQAElHwB2gj
IhhBRtBI6XOHnDDP9AYJ1cSX1BLwOC4vFK3NvR64kHJiOrDMzPRY8kz+m8GfO3Ji
TvnMF3QbGD7X3Ic/qx5ePK2q+noBD+/wtT0g5ZZeUE8Y23PsyQauO5U3gb6+3Rx9
SKWny89DHhIdhozTVQctJH28+V3953SzEVyMV0fYfrAw44NOJucnBWgMr+321eoo
7JiS1Fq6vcXlbZC5qWbrxHAbgH9Z10AeEp447FKV+ELGWaM5qaRe7pXswRlbvcyA
TjTFKqA36eTsxZTkEBbMMW2ttIwCV31jv8QiEE038Z5wPsaSi70RhMYvukIAw6ld
HaNELgPjx2w3IEqf+ZBOp6cW1/auct1JgiZMDm1K2pdneMJYeOqSkLuLwUiFeXUQ
Qi07NW1ph4ac9YcVAVHUwLwSsUQIw1Ype4lWZ8cMuTam7doT87Hnfhxs5npPO3wx
KyMQOgcrPKLtI9Vrn3JNlF1UEDjX3rlpVel+17e6NQiBS7vSN6DecK60gY35ddR7
+reGwEbBRlAPG2Xl4dF4octKPVjhBDJAHy07P1p0pS4iv0zsxOlqgvlyepcy5STd
2XTzoaMIc6IWuI8iGjhdSoxVoSKuK066qoXXr+dem/XTuirwTyaExwh8O00xpWSy
ez2PdZdPTbh9ce8i/ALA+xUhjQrybsyQhI7rKz6Tu/l2CLcLIoAXChnnP3312izW
nEwtP2UgTPLg0p73TVYqsLrtbymX2b9h+K4jKl+3uWmIP/Yy7ftPs6gYQzjOHuG+
ufgZflwyX6UAGfRV1IBvm8+2GtIlvX/yg79fMpcl5wpILolbh1rr1U/jyLYPXL+V
LCzOfk51SiIJPK/CGsE3ymGctI83ExPyco373T4pt+u+kzyvsuselwwh5FQhUIs1
qGazvYdQjIMl4epOX8ueJOiR6GvnFyrN7yJRR7Y3KN/jpBJKS3oYEE5RgacvwaAE
egGF9LolTVY3Xqm2BLxdVmbECRmOHoplD4QUbGwsEL2nzs4t81wxiY3qGVM2H01D
zilrQzdK0mSR0x2/oV+clk9+JK7/OxW2wByuLLGm7l8uCiXBYx00sHhHzsc39emq
mu++KXw5VdcA4uRrX4bci4v1AKe8Ia6CAXf0x3OmJX17x21F5WDfqTP8KzHdw8nq
zFX0P9mkg/9ZkzvgdA+zgGVIGci5uAAgmAmBTutpGuTmQbKNIWRwt8rCTeM6IFnt
aN05AsbHSx2QFvLiJkJEUWN4GAv4wDc8X2NFo3zq9KWAUsXu/teVFl+PsP/HZBs0
ZHrhmiTqHRXiPqNWL4/nTKHTYuZhfrrKQsLpHYOzOssBzhjGBsahLkokuHWxZ5lO
KCLdBilUfa5NQ+Ol07pziZ8ykNjSiPHreUXt7vqYWGR0Obh9c5Z+gQjane+Be+ka
P9KWEDa7XHCVRieSaTd0zpl8bYwGeH7807ohGQ1wdAN68Vy3C4v6CBvXtKaj8dkF
3DrvxA82A3K/FolCQ1C5ECuZyUwcjkvFCcvDVXO0t4j12XVAlHTvecFnW/JnhyP7
Gbpz84+uX6uJyf+jHm5ZD3V/Mon5QDx+JPfFfRKgqTOfHJ+GYzpG0Tvg++ik/i2m
6SzJOQVpIBejfK0iWLCIhwjmkLfbJZ/DtFryW/NdeBB8Jx4w4tATMv/NbvlHTj6n
X5pebJ16lKvtOiNX5z7JlFGOQQ+YLNSCm9XRfSDGXJLG77ytqYCri+h3qltXAU15
iOT0VpoEqdWSfGvx4UQ+LVzToLr7yccSY29CKug57EhES6i6MvvQf3sOBiImqMjx
O70j0ckWXoqpUizj5nAmqo/YEPmQk6S/7XBN2MF26hjaOGbjWadoYJQrugd8eqZF
5Odjj59mR6+6yy1hzogZjK3YjBfqZSxCQ9ip/fkvbMVAYfXUgcNcIYisPpu0tK0b
2ZaZ2PiFq2CiRWsPdg7itLf72/kIicqKpoPYe5XdKeFha51OTQEH73hg3o4aroRm
oBz1dVVGKKgpB8gMAJXX3idaVty25HVvVXaUk3PPb13m28zE+vDuGkXa/7zxyGzp
uLqEv+fbMFJ6SpT2A3UptljgFutG3/SV/SVq9In2oSRX1ab7q1RonDQsxx8/tvd3
aa5nj0UJ6r4H7FHtHD/esxQwqkUS/pC1DO4LwYUaNjZazKW12kHJ3RvsNcgzjB55
JsbCn4yaeRBH8ESbDigfBVLfJ7sQwiBRM7qiwBKqagwBQ4FEmnuwdmVk2FNFC5Gz
WMP5NVCc8w9I6oNqJnDDcEJ3l3qr3IO2CJ9KcmbKq6n9wwecEDEm8AKCFgSeoCke
26gZ7ncVOXYEIC7Q4e2i13UyTvU5DaeS674IlOa0EUl5iIjgLGMI+T3DkYQK8Vlk
CvZTOjBku2tK6eMeVKzYqhRmu6+FdB07cnuEOiWCu6OsvbO69eHOHRqQd+gM7ast
LfMMWq/9/lvvGkBH8H21+DCNtvEHmplTykl8aaSEcX6t2nPtiaQ7RKa64mOaFzwP
DqXtRHq58BHep69VCd3jShSUa+XIdtW5IJgJzCsnYesefu4gRBfeojiqyh7BskeU
qmlZ5g1LVJsOp0OkjBBAahD1eX3KpT5WAoXnV5MMU3KrGPJbLnaT74wMDxQjrKDz
5/M5DTTeAZUfoPlEQBdKB9Ks8LKMY6SqnsFRxaRkGQMtvlR0yYVx4rMBlXyR7WQY
qerPhwzhQEjHMQnEYVczBw4W6n1xFiSoSstUxRe1wmi47NvkC8r5HvFgF4QXvaPG
urP9j2FCt66KdvG2jrGkmLkmDiBIHF8xNXxl+vy7X1ENcDm3qFrXiBgCDSEluBM5
T4TYdRMuCsg7L/hAQ/4BiX3KhhLjkH/h+F/vYFmHC/6k7pja2D4F0mVrgSRLdTXs
0vEUHN35lMqlQzapzmebZkXcolc8bMra603ltIJOECQDCFrX5M9xS4U0VsjE4TVw
x0aqx/YsXx9+Is5vqehEU9MTjD/d8utKVMZ1AdXkC6VnvTuBq+9WwgBeC7tE/WmF
x5E224s+yaqehzrFnFlG10tZ/O0ZTOy0XnMStagv3XJu1JijDT+3vHYmosCpfz+Y
vT2MiyRTVoyIHOUXcFrFbALPm3b93typGIBwFvHxo355lKpAM/YBorftnqyqVv2V
iMSr4m0P1C0z8W5UNfPD5q6EbpcZABltcvKBRhTQ7eHOlBRh2CvxCPITW07PZTbh
bvLtwzph5tzzuzeWXsS9MPJ43VZAat6+bEoDtzC95b0UC45VbdNmRi6DHiYu5Gw3
hEku7UY4ZETHCIpAHzOkYoZ0ADSZUgV2svKvmZzR+uSbS0gkJywiKDdUogLUIP1B
C1aHSYBB5pAJ7dXjTLJ1za5oilvTmlmqUhDkoKnb8kW9WFCdLbeQgNKaSmO5FPXM
nzeGIN8lcUUgxrP+pjZYcSHes5Iu27cxryTtWQvUCtIXm6ZnwwdrjwHMFAi0OzZ2
sHUBSylDDIK9p4dIEZHWPql+WI32CwpDrDkbL8bm3lzPPBJbYkZ3kd0y1CV38Rs9
thJLgKAWbJ4SE7GIpHFVOMrmuz3hZv9qiAVQOhhnn6OoeW/hUDWMSgyGblL2WbcJ
Fs+BDvKz51A1izvh5uKtKShVBEHFMoWkWxEvbJgNsEYVDynruutYLSZRfEX3maDi
Mc+/TDJ5g2N8G58vod2W5H6JMPgT51rxbjb5M9XlRhlT8EcXfZe8BOBsmQRpy2oK
/dp3+Jg6/+YcpoIxO8TBFMNDZGoxNhIz6X6957Ing16X8hTTpIW6lT/763Ltpwsx
rzDdNxcYm6WstkcvOt/9HZNLhoB+8rXQtjihTMWjnhtjkexpwPpEQF47YFeSSGlH
dh4CBcYlNS0xuVJDZDlo/pis75QsajHuLA++cgMFRUwSXUMCRiA5XUNkARvfLd2q
W+2CoDnkJB9OaA9IysexQvtDMO7f8r8OwxrYqsJx697fA+bsiPQbRATH+vFj8c0u
FBsuB4IgHDco8oEuitXauqsVo20i8a4c8Ffy5OTpB58bCfFmKsSaen2XAzB9zlQZ
PWh4slFsQxrv0rvSUtei9Aenk9eD3cgGrAoQ9mFhqNhJ8Hu0Ym4+nqUeJbYozu4A
ioFQZMFGCb1Y3lVj2TcwJIYu0P6+27hYepH7tNHRy95IFiKoFWIslMgC6ZkeVv6M
6huXcIOJQ8POGoTNLmzx6uctyE1Sj7zpsg9mn2wWOYdOh8eUjYVz8EF0RGK6rinH
HL0i7GzFnK18MVzdkQet6dxPjBTWKN49snM83hr0+PoMaCmYRBaDGZmrWTAeGLR2
C9Ep4VF2aK/cm2f8JZ7YUr2Y6tSCGvMLBXNQIeTqTj5lZ5O7NRnJIfyCuYyxcAco
hkS3seYH0PnOk/dn+F36rPRjNlAusWZ0UjjThMcGNzmdGbs5WDm03D464YcisR/0
7s+OyL8RdobdMdBoKQSUAL9Sbd41LR7VhFodFRO0h4iuhGbMp7DD7gHLg5IWzTHQ
a/RKlKo82DFZ4byjX5FfqZkMPJkf1VLQPZnBBjW5dxR5sdsrckwdTszdB25AWaMG
1htUPOHyVZ6Q9SazMsklkzSVsHe6+cvv70gTZ5T8xTe5IEB7+bNZFg2F2sybGb8u
/+EJM35UV9K+8j94qQIcHFb/iOIYusf/hSChcA97lmjfDG9zbPWpYtjnRbyBKNKz
3Lw5d/244P05uafwMB2F2+RWXg8aVoZniDSB05A8EunISa2mR1Pcvx5m41EZs7ge
o92X0PcnELV+GGCK2FVB1orZro1iUnkaiOsV0IercupwI2/7xNQ82/3dsIRKX+bh
gqJQolXCeEyoUO1BacKSwkexQPhd5y7SDPHzEl4bysuWc5F1CvJej3dMSB9Nxcln
FPfTHP4T+meQcRqU09zYItiWiCmwiQZfKsOI1I4TzPfJ8rU++oSXNUjCSqinLexS
gfvWqKKQiqt77C8TbIqhxb20GAyVNQQ16r8vhWhNyWeaGK2Vd7MeLC8bUEgsVG9A
Iui0lc97iU/AtukVqncxXqCRZYBG5Y4RSOWORjpCGUTcUGCbCxTm9/dE0FVhCxHu
IQfGVYzextSJ4KTD9QTyYUVt2hgP4OomHFxWGjNwckeRJHe1Hxu7NWYEQHpOAxiK
i6tmad31Jn6HsryXEs7OIF+6PZ9Ucr2A177u57ZI4mIvlr0Z5MihEIEr4emWuGss
uwW9b4BOoBLyE70FZcc0E0ccLW3Mtkeh1gwEWf87C1orazp29a7Y0GRb4k1AOQid
+V9DQrYcacTn1Y2L0UhLaarM+9DEX2KYxJu0QofLVuo7ccV/HsT8cHU861cV5+jX
7YN3yh2EkUpCUMS2c7FVBWcs9WeQaBpqPrULyNjZm9ZCKzGo6ZUInf7ACP4V59p5
ExPXsxQEMdnVqbvQE+EvSD/nvkdNgmjejzwyTIID6PxSok1488tJ8kzO2+WDfhvo
rmidX7H8GK8LN2uU2LRCj4Y5sYyJ5dNEPCQblU81YSug/zUQuxPpg86YbJHKmlfX
OwCcAC3CSzQaMFz1DEag1HZHsxrKsTRhrnHjiu23t33vRq6NYs8c7VoFI2MoJVj4
T7a6aMlmsHelPUox8Rrp3R0AXHzA/lj4qcggi9SLDVbqxV5ORY4wMib9UAfCSxd8
4sEv7bAplLlk919odZ1NHvUtIUd+0CJfbNnw1MagDVEyDqXwHDRjcSpYA4IV/0eQ
N5/hWiCLdKrvPgiXZyTBqmUC0Lru3OkVIDnxtnp270Rzf5fjg4K2x9W5SpzjfBEW
UXS+0wsWVl9cbKseszuJZjpaZqf0P4nnzc0We2SbsHvy2KGDV8ooZ+i8PjpfhZsY
RgCMjvsXz56wnedSAEmpWcJaF4eN8PAYPZSfgcrwV3LhW389X2zZhmVCQW0xrawt
vHJCLxtH1oDp2o4ELtkJXsgGWtS5G65Z5gXIzKB7VdBc8uKhY9ckH8ZBeQ8aJ5Rk
lmZnppf4ybuRzPlDrfuo8U3kpZHogZJagzC3Wuh9vLjSUzwrAbMqZrpj+uKurIeu
hmsUsPPRFv3t88yXpM1dwyBRhe5q0sXzvBeXJBFOY9AQ0fQ/Mm6a5SFugCnSDK/v
x0Udri+JPOSmp35oScqjK2MzxUDwQBQoGidYKXy6yHbiRdm+htuxfSKa4/uoTsgz
R0PMEdV/2ctUVlncuEWJnQWrdCYZk1OWKLvOVwodZHwLiuskhcE9TgiVsxyrmdeR
ePDGzppd77emJ6TIWEzLCOovApNHJmPw66Ctx3u8b1kOQxqrdBqwXaueBJPBobT9
toDbMaTyOqS+g8O9mpYzpjooZmYxwULu5oeXiDeZGbrwm+FhUE7G0jc4Ldm6NF7k
Yy0InLkY12nLhYaBBIJ/0ovfKh7kRguHdWvESHaerRjGbgkAIyW4XHjCfTWy7fQS
rsShpjBzVWgsqwYb0C8dy3gLfUAXqpvp0htQi3OH36pQ7o2nMmjibutaFXr632qw
Gixa8VEpAfMxiD2oU+q/ouyqlLpeq6ExMhR6qWS0IkqL9wMNbC70qP2JR/9m6T0M
9b+3UxBYAiGxnRx7Za0Q0tkgpFeMsxeccm9DrXkExs4XBIqYZNygkGwG1P2J1OoN
XFLb215mUkLJ4uKzQ5/9ql5QKub/DVFx5kYdnf6Y7KNm7gWw6CnaZw0DNd2KkCBN
6q54wf6HKbqC4Vg8I/2smEnxlehI9jAsZa81EtGcUCFL/254XDRM3WmQFZx1D8yS
Zmao42JFU3DJplxTNlB5C4uQytR3DsLR1buVbhCW9bXtuAyKNPBKzYk0MLW6x4I/
iEUPotqjY75/MZxR7TIHZJtoNHCnuWOTfoTYZpAuoQ7FJyhZufvVrjwsTXnYQOaz
ey74AMsmaAm5qhHn4BSKg89GzZ9722myuFKuXgoFuO+dkqcoKbXOqhQ8Hdvs+Edh
3Zb0ML0CwLQs+lcpcDjBObaqBye3YgQbjgjcHEjmW57tVXCQdM1X+J2kJt1aT2Gt
HsxBJX8h9jFGgJnnwuOD+1L3xJ0LmA7L1auGg8PTQZciJ7FymbnlkEJ+DinHAPfI
6JwCtF8GqOJBA6KQMpwQ/ZNbhjPYY6q8mgPCl9R0uz6fQ1Eqt8Ylndz5tmTHSvak
hrwUtakfUZrXjV3fe+Gft1iFMV1PhoGN3RCVqkbcRElPsVA3GxGTJGN6r67OV6Xu
OD8Js6TvuLvUFGrKTouSM1R6sFPdIrCbwsSti5Hy1HNpFCm+FBQKEjG26cLHLEZB
Yx0NHFZ3pr2baftnWDV2Po/avPh5CfJsAGeSxUxkfhvW0PoOUwUI/WbuJK8+kUTN
i1zobDO0mOLvzA6AX3uIgpSntPGLvQopgRzhGX2h7UQV0zAQcL6vUH2R83HdN8+C
3dYkSL82sJEDiDJlsS74w4hk0KUWmOEwBb6TVrc03ICcIaEgSrXWUdsbr5iV+l1N
ErI5k8WRPrF1MYGxDhzSBtCfFkMYupMxJN65+qQ41OtJTi0AaFHK6AGW3OuFsdk4
4tPvB5RzybZgWjsT7keJBtbET6suMiGLz5CV1R/UMT3dIQdzRvRPr2YmX+v/1U4i
4uYkcBtdXx9fLVy8IQWHrA89fN2QKpcYQ2dMbLVhvAPY59q3GjP1Sv+HFbhso4vL
TT4/eybs5mXtBzOZL9QfQLsAoFwC3A3MG+LD3QBg4H4VNAoCbCH0gLLplp8tOCbW
q+E+fzC+lC4Eb55upcx+0UiblejM0ar98nRnyetP+960eI3KBZUxgtyzmmQzqwb7
1FE9L05/TxN7EAQEHccPVUnLlff0SjcLpkkSyFkjZFecTp9/pTza/5XQM/DYT12K
ed7p3z/Dzbr3HS1wINcYVMLgh6kPTVz70APu6LvLIKHReQDY9A72WhhzfbCK1sAc
CC434W/KzzNsU6dg4zWinmM5OwErJB5arKBaeIDBw/QVjLnkaiMkI/QhV2hWXgLH
hHPvVpt7G7WvjW6tJdglEo5St/V1W14nnzpiBiZ1x4GwD9+BXXSXlB2UxCiDa87y
0vVB5mhRa1HvpOey++wwgQFsbAGekTFDtemnKESoZOdAD1qnmFUH/R1D2znUX5CV
jTiuBeWGo2+pGGxdCOpGDZFk18nfWfloRzVFUJIEwwgfzGbJyiKJGb5XOx5llRSS
krvCjJSmhFsvvxL6MnQqHXxlLUbS0sq2gnTx5gnl4RLPby9uzYTsh//1j4F2rZDI
aobs4sEFlhLJxX78CvdBZNgiWFmT6EObmu3/N99FDMPeDpFD+/j2/WSjrsICkH7W
uaFHThvCktUlXaUncR+9z/RaQsF0lY/8vpCsmU1bODS0v3iFyNdxlLikyZKK3Pni
STrRXA6FbYaz915s2xV2NhMbVfzFS0VMUaMVBlZKJX+22OUecteoAlCpV41rIYNe
TdrWlyRu7yOaC6sl3L26aG/+UKJeKaTvYmI919uC3OiR7Z8KOUiNY9X0LaEEpC2b
5fXbkBR45BlGwQRQ3PzE3m8eYZrZ05hTRk8kJIgJxgnSvtNhE3wY8NYw/g82fW+j
lboYDEuu9F34JSXgqCTM87AS2jjWkU+OoM5u35Ay95R/cHyNqEGjpSCplzSK1EN/
bcVYt0EA9zijkP50L6Adok6ISZ9J59VqqFIeaOsgdoK3UBl/9hDb4sZFz43LdaEK
Pw0Qp+s9nIuzkJVnZM928lj+G/EgYoJ8YUWoxwK4w/JRGcGgcHVigXs9LXgAftA9
MDRdQA6deiXPE9JbD0mlbHIgtW441xGgRwEAC1KSJ56S1fEBIm49IZqkLQlp15yI
zlVFZriUilAvAxR/BUFY8v1UNu9zlLnOU16fqd16af+sESW4fm8RI6MyI3r44/Tk
EdG25u2+hVc7AGm3YqYTAGWHzvzg5b9rLiWNrhkh7KbABGtoAmRI+oT6vkx7FyZL
bDbJ7eh1RREYcs7toeNcZxPhh3RzO+c++o+xJ+QbpdVGclJxgi5xkpDzhFlmxsUG
RAYhQk+2mkn9spk/u3yyxxUfIVPFETJS+Ih9DwRwLf2NU/p3htYIg8yWWSYGmqix
T6bmSpi+j8MM9vEl//W5id1zuwU9sHVR8bfbcGMEgkMx+OBju4hOzIStNgHErYjb
/GZzaHe7s1xFoJ7hygZnNsAXbBGM5d0YNjeTaByUiPtd4DYHmzM5IpZt5mQfSVXq
9ucoIkXVrzuUj8dtV5ulzHkRG1RdzZFAdv3v3ZxhhoW7iYnhBWtqhBPukNo86H6K
EHERxnP1GO1aHJCaW0D+ttSXwYXW8LEnaBsPiJ7oCQamfzDNFVHt8GhYA7Oh4G0k
Zj8wqYTZ2zxvgAAZ5uNnfC8JRHUqcwAYVucSSTjMRnoUkA2yBtuRFLywLDg/guQd
Su2D1Bvw81ZiIe7cJqmYVscc9R89ZKyWMgLODpuzc+ran2OwWnwaUMBlT/BaWied
X15rmpGowKuDwnFvRprrTwXzuW/dE0gSpwdu41+1CVD3E6aG2LJZxkux8UkyJEA+
aZva3wl9L5XNC8KWhsOVh0BGDX3I4/Gbs5PDC+sJISFySQqC+7/myHcZb/aXHPvK
B7ilkkAtp5YqdYU7lLvOroM8u33wMKFRDJ215+3xQsLOzXozqc72Zowho6hYBEZI
SfQHqYVxYsH87yRL8aENL+2yUtYZ+R6B5gWzMeDEk3YKq5uYwpEAwCpHW5TNTlAO
e1Lbw35sKhs9QTPfbN/w0cS1HnxVs2oyKaNvxdrrvh/blJeHhUwjWgh1K9ZQoqNh
u9BBmq4jok6a+dYHRPONzD0VZqwCUI99QkSnvfY7wUb5dj4W6MPvtrCrU/zswc9h
4+mvzUBER+FCsAWZyyDZ7uKeaTjVpYpfPJnalXsO5F9sP4hlwVGJXOFyHGIvVTfo
TUQEjkkCBUy4ULwd5urpdtHZvxOcKh5Gh9qT41HMgxNA76BjiVs2LaQDmXSdFufk
2p3vKEjDzPZKLs26p5K8USMGpyDtvZINmz62jzTzJYMmrJ8M0cGdvIx2SWAyeJZ/
cWOkzYYdgLVt+2cpjw+w41x1fWQqyO03FDgaCLPD2b/EOI/N6rRDApW23FPQudKa
JiFYisvjhViaIVyEQ/cX9vq95qWRIYDUrhcVVlkzYNGZSRM95aGa8yMWWwKz3t2P
0mFYnbk/f+2AEBPCxRu1VywJUa6jAYeZgVQPzWNH7WHyCxcL9W4TG/jYZrxvO0Ra
oA+pK/83qmA/7ZG/wh+2KoRlSNCCz21AulT73aLGLtqLiuA3N1CiILXIHBa1E5hq
uvmVFVCpLjNnyVsQNxI3nRokkpxOrmx6K7GXqmBQqh1nCTEUA1L5KRVo2PRuvFzo
UMJIpAZCvNXhq51OdqdKpUKjAVbyEptZiCktH/Tp7nnVMfpMNyzICCYcYH3LOVUZ
quMCkVXKsHJh3uxM709D+dK0HHITd81jAz6Ow2KcY/9OnH2SCoI6Cl14wCrlNpdu
o0uqBbodhXhu9XGi3yl/DNqemy7OSuko2LTg4KdvIDutC3y29buYUi22lN2a1NEQ
UsMLLzrG1pj3bl4/JbizJ0h95nLQzL+26RTUXvYiqM/UkPNZhPNJKAFsnFh74+wn
Y/VbeJKD1FMt61Jh4enmhg765e69oUwMbiyWGatgyB1a1rubz1VSYVj0grK2KXjj
RYKEcDWgQgwRtRiS2t9qlYhU9Gxm+RQ6Rqqc00IR188UpIe29XIpp+vRz5xlvTjO
o/m4SmJVMqP/qPfA1ig3eHxOFGzVPYO/e+Q6P6pC+HYlZWIUqYce7fEh9ehGGkZ4
EUgFNYJbLxKU1xhG1TggTuL/CaYuy3Y25c06SQbERLLJHYgmevuSjZlFuj26q1l8
tv3DZXXmfH4lbeuQLa/Es8xADWbQ7nO3zg1h88Vc0W4oZ/vrdnewconypLrsb7h7
S6bFzQXZnn9/+JyTd02/3ieWqFISMdvxewFN2aJR0BdOQJXFJaWY85MrLhcjSsZq
PjFMQUajemN9E6Osep7XLhFT8S1RBJwz/Jn0crdBovj8hdFzXNggqQFdlBsqElkK
yqoLM9LBk9NjoJl5Q6Nt9pkLrOTgY2GFU1YpUyLRkJP6wvgUSfZkml9vvcNTfOtJ
/j/Irwu72HbOwXAMWqjIEoJOTIxcitfL6GHKY1OhqaodLy1/bkSsk/maXO3BcsGu
KECyI0jO4d+82lDjPILaH0l78ozw4j2vAw2jGYYAkJhmc069FfSUYNGuV2Yzr1Lh
FeA122/8Rs/7rnYjDSgUKOVCf4ZZGjwIwlaS4o4KWNtp4QGUax4os1D7FJY46Qp0
EbJsmIwrcTw4yxCx7AKGZy8Sf+tLw3tHNBh55yOSfu9gxD+ALFuziwrWbNKdh/nB
xZoL4Ktcb4psRhQk6K9EWtO769vhC+dpocIxNmCeda8JMn3Q3S60K780uIvj7HpB
v6aAJeNgKzqO0b6pEncapnnz2t4PF6SCuZhxzxBeh8gy3U3GuB5w653vsME9NAOd
ZD5CZgXATIpjcaqSacE07q+bJBtcqwKriIjUjGxbumgWE4v9fwtQTL9+5KfABMp3
uXVYYMpBiFq6gip8vUyLeOcDUVFkDIb0TWiKpnm0NREcg8J0x1NXfROqQw7qE8K0
deFSIFje7TmoDA3dFOkYmFaFMGP5ZD0U4S/8EdSiDpv/OQdVe7mW7rUuv0jmFFfj
xz8++8H0n+o6KSSD7Eg7ABl2Pw0ARnLQj7jp/7Bm53XdmJGLdjKjeeZPbtF8OUro
uzMuwIOsMLO8Rtm+h/cFZf8aKpa+A9AsA6wEqALQ3dKaCn42j3hvxZyLFO/cOymX
RNAa4lEyTWlVw29IgPL/op9tA7W5zqUy28fJ/6F/2AEe7eSA7+QjT0Z9SucV1Kv0
JIOjclej4MNk+oioNDTvtXi+Vnii1O8I4+Fmoy/3U/jfbedP6yuln7Exj7uGyKSx
yYJlHUKfuDov+QxRu/sqxr9oo+s54U63VVZJSuRXphk+pTuXIpDPrvrCRSgbiKzm
G08bJ1vKq+GoIOffzyeC18zAle4aWCLk4fn68NH8lwx4ZyrSUyM+T9GMpX+Q/9eF
v5GOJifJeaoTZ/W6g/IqfQPFKrOq7+eMeJ9cQg5gPFogCOg5KFwo2IUwvYLIKywi
5O4PxPKVABZjr+N2l6zFgSrsiKhtH0qCiN6edQBxjMDeZ8VRaeLatcfP7rmg8E4U
4CLd2+2fB/wnretcO+u1IbccZZ2Pd+9EltV99i7HATTxtj7i1lcFwXbd9mOyR8Ar
y7/zZ54VNkJEYmRIO6Tp3JXig8Tav1n2gs+kz2AeZuKoRMMlpYnIDvGifgL8HnCV
mx24DZCDAXMFAFYMZIDXlveycoHD/v6r8DfIFcOp4LyY2SdqHqeAwnY7DuczLoAx
Mz1mC69TRVci2RofM70eojQc/PFJWuTtHPRtLOJaljh1qYvkcKxIWEr3Pc+5bVYq
37TNSM1KKmNhXj0kfiN2erkbTpNln0L8Y5FXYqEvFQhcUG36mB2xskVW66YWO2W8
KWcbJWHV5/c6gf+gQRdCi1vLXIImiLKwGBbKM2FWus7gLE0WtKS/u0PQLaW2un04
D976isFW0c1Oe70RfXbdJzcAChkqd1RdqELau8gfL1wLL8GXxjuz9CIaCqCkqhkg
gjZXlI7W66HD0EnsjJKQzVR/FrRrWkgQ1nosDBb0OYXVUpjPtKh3z9d5vDAAQxcI
zcfwAog0X1HP92GhNkM81ScObZj3Abc4pn8iqWVxbdIB54y8NW0+ZsMFSIJTPF3x
f6PJqlnPZ9a83k9WGC3LCqWUMLixuUC3x9Ky5WiazSCySQNM0SIXzurJzB06VHg3
Ny199SEBXLHyiCfpdq/LmfqXXEEpro/TptLK1c47PyRzrlAyZ4tFZ7PQOfjgDfaD
S9T7wLUYP+lueOpTphfjt+eIIs2AFmYaZqWPb25e9UHhUYNJ/EjSMrc3vScQDQbp
9XC7obRmgFIW2YLmOnu/YTUW4dnl9PVypnQzkJC8cnMCqai8Z3bvdcqKoOSkv7S/
K0TLhp5OWCmN2hi4JeupDYnyXUBbiAYobFAcwJRCxiFj5UooD+1GA/xUDpsfqTsz
EuGacoxZs2obKBy8xK5KEvPyzTu6XnXjbjuKmyS0M7qPEtoJFUJOhWUDdI5R1GWL
2Dakv/oULYcN8ucjX0gYEBzhsmf0a0vc61AP4MQvAWjqlnJScST9F2BixV6vutBP
4eSNcDuFVyS156Sj2GyWuFQF3K6RmQontzW+Ai8eGFPRzQbjZTAmHRGhY6xwlFRk
ZXw07dORn4N0GKfnyqWYYiURweG62UNmz9vhoQ+TNuQ16sv6TRIHVDSjndrdsi9z
7ZbN9LQwII72VrDZHckn4LcWqn5fPg6s5LnIw+9/Fszw/wN2IMok+1vFi1CEisqd
ate4OzajAD9U0LHlDyt6l03+mKXjJw5YynoZfwVuEyoCnQZqT+F9yGFXGU69fORu
NJ0eZW1dTDOyDfyrHLo7UtQW1NYUGMKhix4YPxswCX1BxHwhmaj6kqnOXGysC79R
SHuxilAxSNBQNXSCrL/JyufyO75SDnBJpZX/I6jTEqTTLJXkOzOHxaHLf0HkNq/O
ISLxSo/owO0WJSgHQ2I1xUNMbbOceVy6TEQrMsvmHAR4AXmh5hWmuBoHxp7qiyq5
Xw7zob44ppCGmTgNn+ebOMunoX1IxFnEzuPdCIW2//ZT7h8rGsL5uU23VAKl3In1
mbTAMwdkIKH30GaXsjBVJw6YXejXv2+mAldB4nODLV/s/kutA8rYo+fYIFC/EhUT
hWETFPtqOYanbg7maZDVdLy5oEm0uP1aFF/jgV9lGOUluyqGoSXkJJ898DbMCuj+
N5O0fS0DiZWiptCzFA0+WZ217rd0plqO6s/ez/gLYXZgjD7zfz1z5gw/8xYezz0m
ArYBCoKw5XENQq84qlXYrshPxZif3c/6oXV3PYaLANHV8pGl+yClGccj7wbf02/l
aj0M2B8pAMB1Q8GssUtxWFlt/NIDXFqEL8BBEiFEt/Jru+mG3Na+KTGIknxVsL2F
5C1MfEfxYz71cKTp0gp6naSYioHT0CvB/ZlmS3z/i0etcm1cWC3RwX0L0/1Eqirr
sBjlQuTCA48KoEEFnse4oz/VbEz9Rtru24wPM25UolrGHklmQP31CLdZOhHnovmY
bS/TMZQ9t8QdgRlJ3KnFnIDZgW7mjxlqJeL30zsIaFYFa+t40dUNxE/1XKtjtAG6
JcGGmLbR8D1Mp5k+6djHL4qGr9lai8hlQC09LhidNb+HlXNCXdeDXKT6cU5UiNuI
xmwd1+xEHH1fhTY0jlU0BT+2CKZ/BhDWI4fKOZizj5Nk9gPMeCB7NwHo+J0Ud4+r
cyprM2Nr9WWUUGm9ocdtLYwkwLTNxOswFHg9dy32+FS7nmVK41QPuKziSE1Drq7l
2g7QVXPETsH8ogBMg56Q3dFjqGMJcQWcVZIEHmsKJS/kuY92ZYIO975yErUzffzF
aH00cJeZXVKjeRuT5Wj8s+K6EnAIGNR+zZ1yGAypzlp1n4Mk7WchZVROp+Uj4GlK
TENqJ5XqS1ypGsgSgn09qcaUANN0Zn4z6mHndQslweJT+oKSbExO4jTOxFOs0pFP
oDqGQqeRoW7ikLs1kbLNA/nFeodvTqgumpUP4Oz66LcBJogOM2e4lfQ/5BFPWFuH
Hp6+x578K1zbg/hf7Ie0TuW1XCPItGMoEoBZGBREY6apPYf39OM5uLPVqUHHfPB3
7dnFeqk/KbF9Z3wbxn99seFwt7AHym+XWNEKNqy9hP1fBJFBAXAnFex0JRnzR8L9
8TS9v/xyy7z/+InJOWiHGRSmyn01b8vKnshwqzS3Dfm/AYPvulz+UmhUZOPyCWHz
ru6j/PCu6CZ3LCmV5R2rVZtmAObHS/QpmuDNFJUb8KkNlo1HYCroJg7F2GTfQKPM
Uf0gywfDof9Fg25CyoWIzpePkFIB07ULh1V1eQWjo01Gkx0/SCKsYd1KG9FUpvwC
jeEcD/WrQvPAwQS1jvJKszABrdyq5bn3xoYn5QavO96pDk4m3n/bqQADc2rb1gXs
hWEm3Q7z0CJJRmiNj8ZaxFumKhcIQCa2oAYAbfNg2z+3zGV8mavM1WYVdreIuba/
rlkGZhMdN3fhXXIUavvUbIRA8jsyJ/KZscw0ejTmvQjdr0e7R14o8E5+DXlGnjEP
ltDFxzTQTYSq+Q+HWoW6PxMRLdvu8AwlLPXVWhTwhT8hiOjVIuTB+tROulV/MPNc
f6YkjG09O+BqJ85exAbsMUjU+DusRnM3hSP00QTG8MJr3SpW67eM5V5GEu7lrq1L
v8CORVPIMicBbpUpreURFwIWeGyMX4zFRrq7kdqdApbTnLafNk314XMg6Kj/35D9
T7B4xTQw8kl5mpERJZ2181jHdr6oc66AW9HvnjjilWAlFyowCOUndXYvPFcJLG7F
7bKnFdoKutLbfmn/ptkeEzqkja+zaaxRst+U7331l6lZSqjUYSIbIq2eH+u/MhNP
/sIP7Re1Gq0xtpUn+gahEpKSvcEnklQAld3NBNL82EwIQoWWTm/l5FPFXI6pa0uK
SldHLw7anE2gDhfj9SgVKGtmBBhqY3n/GwAzavRLHQMiaEMjT+wn81830XPg8EDU
FE18NJSn1zU7jufK878pfTEAWcYbKZH0Bo3NSFUdnqt+zTaeQ4nOnSfw+ry3AXUI
tP3U5X1RBsUlRgekbeVdJEs1FQBnhWCqEMDVj+XbTK7g5h3uXA7aEk4c+92tHWIU
IthOp8FaJHdH3/900I/Ym51+v9WX5jqzxvqYwaogs+cZDN1D653utjTRC7ncMh81
QkEdVu83slzOkwnbXN8e62PXdNRvIfKlRrQpuzaTSrdj4YzxkT1hhYVEqRcE46lq
bVXcUbBS/kpqO8IqdA34Xnp1V5Ve+4SGDQ4YbCZSoLnc1Hu+L/Zb8McBYp4qBn+7
H83hP6YsPXfXhw2JyCnWe38PXZm10wYyd6aqlWHa8QaGKBqKzZcFEBL0FYKeMiAB
GuuLNioB6/AoWrKpLjo2AiVsLuQyysHdKk5dRErj/tbkwE5qQkk7QopRbatOAuRJ
Tgzw0YCF0uziVfJ82hVhb/xjs82ZGRqnrE6iHbpbfhmJsqNcc1XQ1nm6nEDtpEE8
QtiuhRwdeYT2z7xM4p6YNPXSc+PfzPUMYw+yyGaJ9NILaXHSh5zmF7VxAuxQ/1jU
ZdqwLvLhqkqgs6ud06Uhy8eFlUjaNksjfyY2gmrCxx1MkWLFCnm4xMCVAi9Gh6jF
XGfc1a1o09YuymMPOY8e0yVXm9W9a0EUTp5KLwZVVLKPodtW+ACwGmr3Mlb+uuSS
0xY/KdNyaqoDyZdzDd7nUqM4/jIdjCZ2PmvffbsNXTFR5teYx/iCFkrau6tf/Ih3
t9gi8Ola7Yj5lxzdEEhWszsPFmZjjbssuwQBV54jsZdLPOtGUKhn0jyrhQ1vLl80
ejqph5mXeN0suORkadIAemrbD6WSyogPgm3UvfOvUyykHRCnmlCn2Si6HgeBWwKW
9cr11jPoun1arflUI969jpG2254YK09b4ghTxgiB7hmZVvUr1mc+4yK0tlF1flEL
IzoBuMmSnTxRzo/4xKMdBq+YWy2c2sHkJZxW6L7UGA94bnpkSLGMgiV4FphONhF/
M1oEO8owgnLCOvVZywjfuS3gx+kWaUMXZJ0Lg6mTs4R6UBfPHc0HwPx5gjMgSDeX
EZ20IZVYI/h+3DrgoSCRb5dtVbEfStFjNlfHdWJdY9arnMiUyGD29Hnrzp70ZkGJ
hWNiQPsVhAn7v2Ly2ikm+EQmfjBweVBz1GYBV0UeimI40XNm4A6FVuGnfys8+uJm
ysmFFXjZqBoHNw7ZbScTgOwURW4bO5PCDeM1Td2yrDGwCIy2sbB1iplrewt/hfXm
eF+DhX3bp2nIwbs+G3Kl5RZNFcsex6MyV3YiIAZlZAxy2F24sdgrknv9yEvh3H8T
Ar4sSVYL4lSo91ZAYor/fPHcEHfpeenrUQwLPJBoQjspmaBVBjfZuIa8aRrNng13
orSDHoPH86hNz0XCtwx2Y0lgv571L8Ajai+E9t6IW2fFrJvmVWdFPGZX8hL3nHF5
h9K0QiAG87+OBf4ABJbltR9IhbAfN+NY2n5hb4yEMXck1C5m5OTyJDa5WLokEl+l
aFu+WzAh6v4Jqj8xEi/GLswvhBTNaFCs003ljNKplpfPv/bzG+qsKbDhcUE/6imx
gzjEqZ/fd2YAlyYHZ71977Nv+AkYLag3IHyiDrrU1dIHD3gFDNs0/ary3Q/bGIUh
BMgAlIYwNA/ksRCGmjtnAUeIZgWIETCQtaI/jVWH70nTp27MS3PcEngpgKxMYl0d
FUQ+3AoVRO/x0Mg3PmuiH2mKFXaljWc5YFYcn14gu/LL6Rx5q4CzfTluk0L/69aq
050SZUzCh+KN6PDSnkuAqo+kUCL1OeJdQUEBkTBbjkpDixOdaQ4edJTi2Q+DpEfI
fXTAWtl1pIIyPktWo3+fVEBqqIxFUoWOHeM+HcR+OsNUYHVoE63F4rGxbErcNi9V
RuGV9vPIr/yVyk18pi8PMv7JFsxDcYf68XLABkx3PDKoXBxQ41IFZ18XDd7UTSYo
+qQCIHIYH9oHfkqFWyWLPxrfv+K06wiO0u9N7E2uGTCGUwXhsUsUVql4GiUZ5TDC
/qoJCP0dUmds0Zxu2V1MGOZWmvgV19A3jiP07LwZPg30vD9XpfynmRCwDQyqmN9w
ix6WwFjwk7p/1tqaPazgUH4V25fPXVpUhk18wQl+UJNA3szKd7HG78I38EqlNeMm
+XgyaIX4dlegp1+F1LVzOBBOq2SD+SErFflyBaDENUUe2ffmSXSiS7hjmJkdhHmZ
J1DGkeDMoABHp/ZpXbpPxr6yCSHsgt6WizKViMia8NGsliwVE/sr2vFhSRAPZPGN
VeMzlDbTaA9YijvcsDqNKsDmhR7O9a83s+qkbQNDuYgE3VeEcJEPQMccQ8FOKFDU
PAa6COjICl8zl5nB6GHeY+d9tidcvbgUEip220LMmr0FOLIp2lsrpQUUfbNQNuEL
fwTnH8PxQXWBVFMhaEeLi/RrdCnEiR3ZXQqqieDnW8FIjV4kMopGWfQmjgBoF18t
9T7OpE9BS1qJ64uWOZ0z5jIKQyFIVMI3N8seVgBCXSYxPKiTyySu3fsi22E9Irl0
+R9r97hKon2Zh7j2jlvJ7VdL4fm7qiWWOfPZjN6ONtZCkpZ9guvMCJnpjghcRI15
vaSsaFLgR/lJzRLag9EdElIR20d63k0xxPu8xs9RceAjOMopt526kVOA8uuiasHR
a7tzdygq1MlZtz60nrOlXFZE9gqsnrYyDmCzWTK6LwmZkbWC1aU9tkjHkZi8Q24i
vXk0mMecbvyEty8Eu6w0JbdTPhcq2kOYNbPYLJlbFNbA+/QBIy4vVQgtaDhE1d3N
6NFnIm8SL6Iu/dnpy1JuBp8lJEhLhpi2tI0tD4PYvwqExUDfrTb9ek5FCMdAN2Ky
tY/HvrOs3EYTSfN1pFdE97/jG+LvQYvh/3rGRFjpZRRn+tYFkW1vuSb/iOdlJ9Ey
G2s09s4c9kkLfx9NbQaFzJogEXXqH70QBLNl9JagcZ55Gm61MvLSl0a3ATjHfL9W
qR7DLD41iDW0VMhF2CfNGp0LWQ3GqrRzQgYf4Qg4yLYCgrqOcmfgqU70F5IWlqNJ
NIC3jvVRxsa8mZpYxqMY7RKk3JL79MRq0bgah2ziw1SPwlYZWd3ojBzhnPUlCfQw
zA4ke/KNVirQ0b1bv+C3R+eARZ0fYooqi/lCYYngBiQaWb9wVbZJ92n3c62ECssl
bddLTb1sFKxhKxyHoGf175+jXcLxcMiAd3yWXP6t7miT+Ct98xQYUWdsaHCcJYG5
gcqYuDFpJlrTxl0vjttCzmxX5dH5sLRYM5N2g6lO9wPI4ZpAT5we5DbyoM8xxlBx
81gO0/k/dpd2RNNw+TVWjcZAcOf2EShOC3on7npr35Iud6H8jnKOX1r2E9KT4JWk
wFUbM4CziK1smmzRcMfSzE4aSBhKTUvuzLm9/5EHVLjKnXn0I1ERXM+wpKgMrG6N
Ndp8Cs5TSL4PmedhcdekjTMpDvHKpOOsvcaG0OboA4GjCeevUgEJp1EsLyEFLQbu
u9ZeGf4c1nAfRR33H9mDXOAo5RGXMHDyDKB8NeJ+yvz30S5prFFO0moiqEKRkoVp
kHYLXtIi/KKxF367WGoR5qJ1itFBQwXU1IJdJFNYjZsEzhYVOL0eQ2dyPoQGqID2
EGRCfxF6z01teGhyASJC0gNWSIhmAqdhOUdqSGy0aVTb/XP8jPRWGqTLF9HWSZ3K
A/oLygtMixSmVgJu4OS031hGGnRVWrFe1zsNKrJhaXreQEeqQnRMsqvPYkICzbt1
fy0M2osY5t5wTjdHpyJWtUTJ8aMUTE9+3icsTTT0MdBOkPh3FP/6Q9vK5wsP9Bil
WrRDgJcO5KHKkH5XwZ/qQzxW6XUMvNxuAhFWISRePwrxoIWw1+/Rw5pFqFdh/34k
g/VxupKM1D+A3wgvk4KIQdDjw9nEfoXOR1G7AM658ZKWYOXS8mhlcM/Knh+VXo/r
kfgc8wqpLQs6SxTwqAlDxR1rkF1diGhI6Ief7ul4cWfotFhMNvPQv2lLKMRvVvjW
GGFJ5pDniBTC6hcZ+LDIwLrADxeGwxcj3K6rsYQNYFOWxM16K1aOX1kn3XYH8Z67
oTr9BraVC6PxvvP4XLWOUkyuC3JdB5DW4Www8DBgMjiX24FdcRQXDyqWwpkHj/Rh
DbjPHgY9hwXtXUZEqd0aujupRHkHOxx4Y7dWHx/hPrY81XexclBayzyKb6rd/7FJ
dTts7hQCHsrraD0Lbp9/Zxu1bAlBYTzzAC+vZituBRLmVbQ2F2wmZ5q7q/K34IsH
G3zYbGbVcRoKSDJVYMyQ9SH5j2ofoJsOuIY3gu4bImxusSCT0yeuE2unjpmeaAxg
X7kKYaeVWSSV4X+sbJ1ZO2I0L7/h7BzzoWJO9AtbcVIyQoZvl5vSRmJEZFeag5c7
AwDg89fkltJVkylSwpsE8gXfvwOdsAyEnZ+F4+J0CoLduOS/6x/bECbeiIqCWOKp
MgblMKWoqYqG0J0lVc4CawOhqbqXqKD3/3/25bzC/Xft3ztCIh3FYlYH/FGmz30b
LCpCx4gMGTX7w0mGpoDpSkClnJzXNZl0hegtX+WNVr99SUKoewZAYis4ulkKFoXQ
UUkVlVyKGVNhHSCW0YMVu2TIOGf0cIWeSEnK0AmRqnhuj25jt5c9bpLLSK9WaACc
lKqeHQWPONufpnv6t7gzVAkXH6Vd3lKYBBIe9ickRbPFD0pJhGrxBuJf2GvG8gnT
+kY06hAxeoToTI84RSjM0IeBxHXIDQALPNHbHvIkDBCn5YapHDb2J5wKjJyb/U1/
oxGh9Tp/23PRwhV4yweWe5e81Y3nlDR1Ow48eLHCVAdo3G8t/NPm/xSaRpcZSsdN
UdXpXkv6qiSGRzowuFPuuo/K1+sbSjDwfFjs/G00TEiNar4I8mcuDNFRP9cT1Twk
Undeb22gvuXmalTpKdixIK5Lhy3Lv5TCthxUsbgofXGf+pTRVT902Al2N24k3ucI
ma4MWvyyx/Z7bA0iOr8pXvLe3Si6mJJ0TIEq+Gj+7rt0hCqtA43eoADkjEHRp2Qw
ZODdiaaCGYCbv2h/MJQvhIRzej+9qza8i2gHs+jB6h8Qpwk6W/ULVozRhlyLWAon
HwW3faAdqAbs/SPI9u5sB4CZxCaEAEsEL5Fejo0NB/jFsLXen6eO8CY3vRtsxIjR
1bHcuM8FYHfCdYenRUilwY+xCgpIyiVPWwyhzK3b4xW7i/GtSpSHzVsfBOO6MTx/
rO/BTW43bCGSfkhzIG8XBKbROc40b8X82sho3tjTp7IpiP0gCZSY352lfhnbHubx
N6+8+DRqgPdzQMSdmjlFvvWJwwVpan+o2A2YaXtfmflSKjXSbeC8KGqRNrteUd76
3c3ZhPdBkMs2MmztaiehmuAo4uS2PzOYbYdJOcZwRm0wNIU2FUg8N9WS4cW9k/8h
ZE27rrGthZ9VnetZaYsHufEh3gCDJEFatGIUaG85OoYmjzGMEVrE7oFsDyNc3pda
xJ+jIHZLdqBypVc6NsCS6yofsh0jD4bJxi+GbE5BCio4FWYSLigRIa3T1zcPXjLT
KNqzEjZ/jb6P3x0viQ/TGIoBz9u6TQNxPM6nJviidhY91stNsnW/6SANy287OAmB
gi5QN1sPifE2YMKQwu5Ya5JAo+ssfheQw6ep/01q7s3mmdhGcdDvfZXvU355oKq7
z+2Ac1FFmWVe6H9bQwOxFXhi1HhqRYbamNkuiHQ6frdTODQwbRYcRRRCaFW7WBu4
ZKHOqTdxZBfdOozqyJO4RwumtGNjczV7z8NQzid/PZQOcitnyfq4nGXUlryxjRQP
IQuR1fSJBqYUHEMSvFKGHN+MFa9RxoJGs6Hx52m+CSKsdTIz/alM86cmEZtDz+ME
HD/uahxwKMeZQ2DZiJWcFZlu9GTidbb87qSRxB0hKtmrRSOyRVwboEzAbCfjQXQC
DMm9hE2Q5UhkRqV9VBJBv/OopyEZgtKkwcnW0ItEdJGhElhRFtCUpBcspPHoGK1b
jMrnvrFUyo6WzbmFEezCaferC1etDWAc1BI+8fe9kcMSPF0bRpdwFC80XoUJCgbJ
HVzjaRjMLduybPRxp9psTk/HnKAlKX3KhKQ4eu0OUQNCNywSr3k+oMET4eQwG8dL
sQ3ooTVZQtirm31fRYg1Ca87b3B7VwmsS1yPvoJ6dWgueueYFL9+lgguBzOzDVcc
I/cwuce/xmsZAzTz1PUfTWOmoyFQI+LYLCOczZB0205SUJ4t/WC3XGvKkuJKnD2I
epWS/Y60x600BPqPyTS1oLI+izjqQBNvDyLm0mqRgVr3kDEk7SOkDLcDbMpEbf7S
a8mOESE/7CTV93ZqDqfqqVH8cgZ0JSmSK3EF7asUyfjVHxnZNF9Zx0yRIB9Nj6pX
oNVsiB41+XCikJ3GvrJiEuqlwjN+mm/KsUfnGY4M0/pvT3u2hlba/3NWBxIpXJWI
yYsBcoI8iVhbFjDOh/N98t69KGxH9wA6LiMnfN/HJ8i57d+1nvUHVGCpV75wmrKw
7bvcHUqb+Y8n3waCK6GiTN27Lz9Bsh4OdMioSaYw+1VnlunyKeVAPZwMgwmPQGe3
xW9rFCvo7K4017MVHNj4EyQ2gykH+LQs856Jv5PJmH+iWXwQESihFzVF03bmLQZj
vr8rtZigrtd6n4y+xlzxvk/ucx9ldQc/0OtxMtIBJbz6gPUn29Q1WNbA1wzqF/C+
QI+LISKJfUbiM0mKiTUemayGnJAuyNRSIocBj0jqlw6R4nUbqn+xHJOoFdqQNSSt
5jwCOyke2ccW4dBoWZ0kc5L9/MddGRv5nlX9ShW9Z+rec9eS6XQjaXSsPFxuy2DD
x21lBnyPQoSaOySvST9IlB9MYzd84xvfFhU+qb2s4hLPtdFpKRDpXF25rjB/hbfI
5zO0ZMEXd0JXbpQrQMy/0o90JT7GrcrYgEmdIVglM5M5qzAeVbdCRscQwTYApC//
90ldPxARy9JfV2MO97qde/cIpaViIqWHXSBAo+Rcql56ox4eKzVmH07+vSFYGLKE
pKLQnJQzCWhYrDXGFt+d5a3IR4Aua2DwRUkLimr+OzzyNkMCUybQMFz7eiIDRgA1
iAsxFNd2Q2Xjy964Lb4OMQC2spQFxViunZgim/XJSnT8F1RPokzHYnBX+kvMSUGs
r2gMeTBc53AqcuLL4Edk7E4WzBC6nhySR8xsZez24sw01PUAtRzJJnh/X01bvTLm
lHMGnrnUqh1+Vabrgb/3uK2tCInpC8gnGzLM4jDhg9HbCVIV0am35kuePTyG3ADi
m6XfPbSghTT+QXTNqA20ylVKKEVPGOWPuxWjEal3J13EArsixU7UroeqKfP4/Ai1
JXkFokF3ICbLwrq6eSVTTbgF16dIOdM4atXI96MIqYUhRxqOubvriGC3UZTdbu+m
84YXGYASqEB5UP1JqswA9zW1A7t3FZyoJlL0iBLBlstdHvj+XQ0n2Spj4Tdn28gi
Ae1fc1gRxwbavyz7arv3Wb6Zpwlz2pLN9kaK7zNgQ7JZFJudsj7DNW/ptX7YUOa0
iggXG2mSkYU/SibXCm//3LdLouiKND3pyYccy94iWtK3NkskUO7kSFZnRn9y9mZh
GRenZeOQmR45WgCwK+WTbCQK0AKUUxemdaF/cjp0okKUoEdPJYejHRpOaJijeeHi
ou7Tssbea/NW1LaxJ+nwPIhw9Zde0cj0McW59KZjGnXxByy1IPkQ49qdOufsITBa
aATiSxOnSTZC1Kg9DZkuibuefMIu/ekUGjJ/9/RJ7UbTf+pJFGxUWkIJWomTCE4X
yi66uDk5ZZ4I7kbAdx48AG3xiD8OWQalAPoVx5h3Kd8lrLSQ8kYAnEbAGX1oNCzD
8n3k3tijQ1ahMd4SYnuyzqrO22XPyhcHPkefvzYpR0B5tugi1HCdwA4K5+G1yR6F
Mi5bK34UnoQgrr5Fc8dB1RaSvfzMlyWnZDlbv7rKH6xs5Q7d3FQM6sF9zvXJljpX
BrkrQD8OLpmC396OCkTA4rJVExQgieAQgOG4dWIcgoz33YOLR8n/DLNMdq457quo
wBo0BRjIBW0B3Pnmrgup3WG4zlP0X4AJT2Vfyn7RhtymPCXWJ6mknt4CYCQc0WKO
Ys2hq3sh+zqnFAPNNtsTZ0AvPGGJ3Axg2WqbaxbR8sqYYNoAvfbV7hN87tfgxrlv
XYTicQI+bG4mRDktgTQSF/Z/Ymlve/Rw6+VxxTz2tnMLilXSruPXsDs7jXYY0bgz
/UkI5ezOrpIWqPmfO1Y3p3H3SlYYFwL+Id1mb8OVyjWHqNwwbxZ4S4wcQ66PgpP1
FQZXW462VvzgdOLFTr6jukdGevYHsQDEaV/gBJ1imMVbBLToKzITqo7rtmh/oc4L
QeRygdfe/YxGbInFE60At8NvQYLIsxNP4sVQ5A3UgioQjtPXe2Jc1Uo7ZapoGm7S
b4totL3NgvijNtKLq0hBEDYH6TQaoBeRYGpddazoqEaYGVwCn/wVumZa4KdwbnQf
Ge5g7PjlSpkunoGsnJuqwDj2ziLSxsIQUhN8RWPqYB8KLkUpbzdVeySYhp0YHAKX
Ewy/MpVFM8ActBl0IP9olZ9FXd5nWTwrXTw02VFbHkmHQySwPBT6XVz/GCIH6x1x
CIxlO/BU6EEgxw8sVX8Bqto+PfP6NVdd9saGFDbLkMNKzd0LKXl8vQox0NIWdcVl
gYY7pDYLqm0A6q3097ymWRLclXjh6y8bd+qilSk2FDJwREHNjysAkgIZObi5lVXX
NfoZZZg00tW4s5nwvXQMTB93lHXs37cK8E6LqJoc548lZFEfpZYNG91t7YrBnVOS
aekiGTG8KnD8fWe8nu4vifI2QupkDslV3wzD75OaMhHGK+gJvkQ5BckgJOMUM+Ax
UmxK3KgFYpBG739ZKYGNvzUHo4VOPf9yXhjDhOkiOZm3WZtih81xOjr+HktKiv71
yuZ05oNKlAqFUz9+23aes8kzRkc0IJ665LvszWfAk4PTsdgUBEDSXQ728xcPI4FI
jzm96ArXmw5RSnLz9oLlMfdOgfET51XPynVupWvhptlpjpm5F3L7ZSwtFrI/iOKt
Umq7rWgEHM1yedA7aDocyASl+guSUjRKxpTxyuzgb1ugOEGUqhCA1g1nX86deyjW
jVlrVk8mJMRjkJdD/nVAszzfWdeeGxIBAKi0fLgT2xEK3W5x6N+EiqB8TulDJiNw
cezWA2mpDaoYQpFIMvIXYBy8cKR23xH5h/jvICa138OawOMC3QAZoBgylbgrP3lN
E0XDNl+UXgr9gqXqibNmhDx0elL9cDFcMyqkVsxWxURlsC308+1KNC0DHemGrcFh
bGpd5E5ZyUsf5In0pmzkHe3n+LwqE48Kd/3RxefPKvXiSJdVNyair7GtMsxuyrMd
JEf7c4osmfJCb1sgHKOSiuZ6Oc6BQFwVfnQCV3MDHTkhPuJg2VW3BEunVoDRcx7h
SANHZ38Dm466cuMffYDXFUXpR0Xgriyxd4WOI85SoZ8KCWk/6+VffwUXGUIWAKNg
qaBOr7qSZ/tN/qEhC1yqyw1wIFJZfJBFpQQZ8uuiRrs0SSUfsSX2U6xAWIHZ3VIw
pLniPAf36UoErokJPKhxFkz61S2RLcaNhyvDoOBTcR7RHVq70xqwDfueM1GpObDk
ynhSGwvNJ5yxiRIDlagNjvcGquSYZgLHJuDJjhCj1ApMDGVdgFogVjIkFEKIvIyz
3P+11OVldA5o6mZmgR4Ff+VLxHVNY8QqbdP+oSK9feY/r6qycG9ow4Irv+uGR0G9
HdcRWf63b+tBhZ+kotZK+17D1NO7mp2/7+lUlDGBt3c8eIUHjkQtBH3pDdwNJ/mK
jaNTNMGGvsLajNIE0Ks5Dtq4qDYxbY96AhZ4gZzB9Jt169aAlXpAeRCAqUvTpilT
6N7Qx4L5tqy0UCsnKfSbyOjxPlcVgfI5C1/onCWAslbtF7AUeKmpCZ6E5sQ3M4ey
pHAtofc4Lr7pPrs6qfWu2RW4vMv80OqxH/qcEaiKBSVs/JUqVB3a2TC+RznqzdNN
17vwHXnW3o9oyLPmVvQfWi8lWXLyaW8rCeyRR01l9ppJFDRJLAKi3JFyMrfYi3FN
w+a0fVLtnywX6IzcKlvAN4BBPSFBBMpW2UTwD8vkh4FuwT3lv9xtbd8cYfTMLqOr
7KjgUZKw3rolnEHTvUdj9Dt3kAJRo9CrdCk6tq9nfHfqU5aYD7AyTvMp/Nkfu5Mp
B/ByoEYkuLknG3/kYEZ5SJNRQ4Ylg83nFXftkYEeosSJQBUt28RZm67LV2PX5vG4
IlsE91r6IIEcrb+r0KEt55VTqc1Df6kSNYMloO+a7+tZvzHo/8pb3rJdZK+67HM5
u6+oL5mBBX9Rpn0QklxN+/iRbxMI3+LSe0AceiTRcoZ7cpVgO85zSV6qMd2zzkgE
28q+wzUmJXS/VofOAfJuaBFdm3g6nKpVD0dUjyh55VcbDBHVcAY1Qy4aB9Pe4pdd
+zEp+8fRnLG0MIFLy+aDy8xmrmI0c8MVsWia2GSOABxxFD2BUPaQ+bGcDz6Wirkt
oe5wv57mVGNfXUncoBWg2c4JvWEjOglAEIcAV8IPCFUfgwmsJ0oV9wLF3hw3Mals
9A8aUXt06Jpx6KSfNbaEsboMECi20vAI48Lt01cdUzSz472ZXaZeUJlJzJHhUJnH
w+E//99xIc+yYggommyjbw9ZHRlPV4xgxLdyvsPLLJodjMzgVJvvO3g/lwqKUBPL
8CP2eI3euVm33pORdRF+KOFvW4YIql460puaIJc1rjIaX0qh4nyuL+SbB72varpW
gA710AtJyJWFLNYjxTJ6NCuVADLuTju0z+Zad31dlay7g4mVceegmvlgTpeScISR
GAqin0K3b2dNGsfLwWiRO1E+LuRDLZNoTZg7ddCKGG7X7FDrSSKOAgMbi1wAS2Z6
Cvl6oTPpeWBpPcWm5MrxfXPePy1mB2737kfT6zkk2pgOofgEdewJ8a96PCg1LrQG
nLtP+qQSlC3mQnicW7RKO3ClUwWKBxJ8WvdUeDuVa2IhfvPHjTb1x4OdO4HNNxGH
QNgbvxJy3VZeXfZgMSeMmifVSUwnq+LQObYtAt8VG92GHzGkSt+tq8Eeh2evEs9C
NrxhQHV2JMAgdz3yE0lC2V+dszL6oPBlRT8W9hrjn2lsOfO4vgGA4f2gc/ogQaeg
GcpdS52nPhimi3bH96rPc8Ew0GfpfZqwh8O85n6fDm+I29sM1/aSsIioVvFUm01b
uN9Enb6U05YDLhOzLziDSOARWQtNq2g065+p4ppG+LVdIWZ89+tGQCf5RaFf+zmp
YcEr9pU0pgtbr5yCubzMDHriC9qPoju0VH9mXzmDZX2ldk12BM7XX20BnclOxADc
fcQZDjGdcAfW0srEQsd9IftLFqFl5e2E1nyVQfrhFGqwuSu+25AyM7VXgiitgAde
UMkFzlwLzil6HJ62/W4MyXoiXh1WqqbvaGSRQAiF7ef2G8jNXmg9F0dZWNdepaHa
kJkvyOfQSlhz1oJsDt3gsq5gCkHjFSPif+4aLdG4EGTdLa3NT9g/auqATiNpFD7S
QsKRXVCTXG8o1rYXswrbbaTp3PJhdlBEEZIKt6GYv5BOgha9zQK3YSKJzODhKMvp
chuV1whE5//NRxdWCD9ufX64fN/OLs+kUWQDjHhbX7KPzwmFFZe5oNhYBOHwb54E
pgg9X5lYnwJ0TCeMiyy1Z0W/pH7AWCfXOiAmoh7WEHFPSkNAkigvJjCcf6ouw71h
HruHKfnaOPtPz7ngo3ETTkzcMPeiJZWWZI4tNKMFqDhSK9T+HCZ7YszcJAAX1xMe
fwicylSEqJcUgkvp5A5q/1w8IePTKvnBvNuPsUo85dJn6dQCwRpHriQZJ5lH4MPW
H2puBfl/RUcVTUyr/8Hw4/fRj7uGp/aG20LSmp2TK2UCjMY05Fqg2qduGcILKv6V
puuVzwiEBiVUGyMMVgORJVZfs3nZT4QilA9vmbuzysVkabimu2s+TNdzftSOlCvz
boDdcpKpogvyWfjwKiLjChvHYq18/8gJrKYsILG2Y3IvfTGJqnQ/pAkLETWE/HhH
S3P38FnNTStOWAWL92UgAy13/0DFVFtU5QfiYC8uZLyo4K1tPlBoKIEWGXNPoL8E
12ZgK/VD4MzEO8/uZ+JXoAXvBygoFmuvrfJt8b6AqiDntILS4kxqOjlZdphBpTJK
AU3mV1bfvcL22kmTXAAdvJg5gnYhZCIa0nW+j+L/rPwIFUnAJ+mZDl6zpY+C69ff
ky5vQ+9RD3XExL9vZrKJ2oa/RIjnJM+dPPJgmg0IPbQZ3c0TXBVKqT5lNewgsZYA
EkgG+TVOZaYMv6VafbSHctWWc3APMncZESLB3kLAP6/YlbTqamYZiKNiXV82sUGY
52F7U0y+itVAxf/PTqXHbbwrTBh2u0tJr1tbpL5Khi6TVeURNK/wK+KInHQ1Qqt+
nvKyVr0Jy010bCgFWlX9MH/SznYsUUwN6i3ApATQdNpsqDwqbStUB1pfM816wqTi
Evhq/bPUEc7i4XzUZvmGCGbih5uS5hAuA0L0Ez90nK3LgsYlFdSo5uYMtcuCvC/Y
o43p/UuhId6QslHIFaRevC8dwvB5RGa61+HS7WlR3cHpiBtpULcevqHIl8QTmqtp
+gInY6+HbzXSeKihCwJU4mPG12hZQiS9W2LUL2MtIuyX4EBMJ+68ScndCgq4oc9n
clqZ/B5gW6ng0tGLuKY2yJZashplUw38KS5v2+M58SPJRZLrqMTUmXwcgSUr9NND
wZPpi7/hAa5dk8ZvuTo9S7fw+xR7802Y6xXBIljunK7oUKb0OsYR5uJSMdMPi81D
ioXEZrgjvQo+rYqn4UkXNxLv7mMX3z5SGlcymPa/+mdybPXmfbfbAXgV10MD2ULL
cDGEbBs7a9xXqbaBeAraS4rsxmK9TfHolpA6qLvgVm9OxNVnpMM0r1pgY4DzKbpg
Zt/FCn2HYcErMPGYQIvLamf1qcCjbk3Tu9uXh2tdrDG3oQY+3ZxJ22yT+lkj1Hte
t7XsdecATJHMEYkucmXKSKgnecO3FkLNebcqeJB18O78DbrNMtK1Wo0lCYWWxzMl
KGq7ldLua84O5yvYYUxF3LsdHWjYOvdld6Y9ySx3xwoo+GCqnlOzw+jEoynU/uVT
fD8gSb/853POXLnm+HD9QZiMB7ukxf0ETcpbj4F6oO0bnZObld1Zr+VITsl5Y+y2
XpYhZk9lfk8t3FD6OmuCRiYkqfJZxWzDvbgus9oUUlkoR8fPFc4INSWamDO/85YW
D88vb1I4HhvU1hHdmyc/MVWvc18OrQJw9ySM4cEIUJ2rvyMGWdluyB17qswXnDK9
fl9aRIY8re9EIcofidqjveTzSSBL+gtkX4EVKHwUjIhtSByG9G94W8iT7LLucRt9
N5GV1FQ1ZK2qpUF7MWu41oV5hYq8r9VtTy4mdME99O6mODFrzYM/j7599nff6+Hg
T6dZ5yK18/bsHSDe+rh5hMjV2y4AQVGcVeHzcTsue1TFrdkcHh/kQ/Ri9zCkIvEa
MPE5J/PEii+tGaqwSiauy/S63mZoLqXD60hxeNbwlh08oDuf+YQjLgdl2PxG1boV
tsAk5o7cMBsjt8sljB42daRcRfdkAIgL8hNera/CIQXuy6rbk/CjvUmQcUVImqHO
r50URlfM6PhKOyLDvP3Eaba1Uemil/N9PpY9fH/dkqhuifPnRR7oPlgqa4CMubBx
s5jZEWGHJBw2FSHYFdqRhpyID8eQU53wv1X/INZ9v560z++CjPDHt1E8jA9LmL52
1n/7h8Q2GOteYlUMF9w8/a0Hy8DiooDcpgl9B1e/UckE5d2szL/alGHJ7RxrKu33
5D+Er+v1LGlcur2SmeGr5W1MLX3prcgRmwLfu8JCrT/Yj+KmWpSDsDU9NxDX6jBF
C12NZSnh3m9hgMAad5rL2wDdKAByRr3zZ3xrnJZpkrUY4Q3pBlgIsw9vD9iX288C
6WnKU+djvCjsVyyFfoJzr4nzikn46xAiQTrlYtrfXRdhNVIqHLGNERcNQSNxyS2N
1BXpW3Tch5hZ+xvo4PmCnm0t5wa2JjPJGzW/DYcuctdf6fW4ghIatuABUXjZYSNx
gpaeKNX+Xn5c4FiV5XfY3NVK41/EUJ3Cg67I763XclfPX0ogrJak0VI6bJlKiEb9
CD0XK35qosL4ykIevz+Gs0O2RsvDPGMl22DFzW+jBhxQWuKtcj9GikZk4M5RPh4P
3ZzsFXqO/mM/cwRd6oJCK4ykNgI8u2aLyY4+4DAaNwHtKnuFTBzy1UGwqSiPlbL7
V9w3QvmUpmTziKOS/I5fxJbYY+0bMZx2djVM/joWtfJtscRyh82Dt/7tOGCtVALj
s7i2GKXS+mdbL+kqX/xRaSTzZPWboCHHZiqAxfSEOwZnnaNg+/wh3vWpit1KCpPQ
AVKdTDhI2/6Oy9hciMX4MAr+Af7WhJ37zKT7SFysugDpO8gCbCbPQWcogOxT6Kbd
pQnednAauxLIqrhLHp9W8rIkSVVm/m6QpLQfr8QyojQqqk/uw0XkdPd7iPoMcASb
5wlHXKFrg1uVxVEN54s/gTITpTzHLCCN+cHaCGVx6X9qwIbU6letsaDj/J6gjqlM
Pd/3YAUzZEHAB8YT8g55I7K0VdVAGO/xK7YgCNpTQSJ3G2eRMtMj4B6kKpppmhxw
zrssv14dsEflXEOwDGLBORZr8Hb+nwsKs2kvyEXv4glHCFSc4J+8bZAFDnIAOxMW
+sxTy0kQ+90gzUamXu2qpeQw628oHF5T1p8ViM2/0ud8d1pPwRbQxUe2MiiMcZQW
A88yvZRYL7H57gmtR+971jMwma7TDgvGCRhRXSHtpmfYuT9ux00rtmGvCa1w48IN
bqMlRAMONf606D/FZOlMmv07m5XM82efswsJKQMyyrcrMjpDrAKcSdYlPA81hVy2
H99e084DtItjyupN7L6TQl3uxNx8QvEh9JWDMPxPGmIFqZeFD0PyLXOS0vqxc/hb
UHZWsLkchVEKig1fQSiqKl1n6PZk5Bnr6hUTuwDr/wL9Z9YSebxX0dY8mkOQM5I6
KfUXn9iIGrFYAbEnEzZePjlPj9FwsbvG1RL0g4NHAKqsfbUKYIIuC+vYANUJEs5d
fWy7CkaaVbbzW7sTIX8e14N1A5/R/QvdGlvBJXxbfzmTqU52zwYsIj8eWR07iQN1
vsuJC0FcmV9qyp4vE5qTs0754FQ4lwB20SuIfdKQX/AQL5gsMd4JyL56SU2zbXHB
EgVA5keIjes1PoqOlGav12IkJi+jTw/r0cxMXThVY34r4Zum38irf52uv6S/U/yS
xLFkcRYmNzvTrWxE8K/MsLpIRz1hrBibuCMxgwVfgj1cwaJMThGg20egNh2PXxiK
mM5FhBN9a1nGC77VuOt2UnufAga3T2mH0RdIw0KN6G/fxMFy/VWQUpwRBHC10Eps
DAk3Ky8ZU1hSKBUqDhJZitZiPXX2Ut3bmlptFw9kLBmSNPziqZuvpSirWb0M0hke
3MtVEWxoYAymdeESaC3rBjVmC/c/gk8XCv+q0IT/Z3BMac05JWUWfZ/9gRLXV4u+
P5oKeSPWxvAL5COg1wNrEzy+lxIZPfYJB0vMRsuV8U+iJQGz8m+R0308VFr6/LC0
3sj0IvxWTvyxFTvDZxuK6MttiYlk5pT0f4Qeftg2T7xNiiyTUV0FEeqkwZ+gv51T
YALreDrmF30VU/sMICzIood41TzhOUoTHTbG3qiq6Grof2B22+a4+Sqb4WwTIl2b
2lORCTe7MzUJMaExESvH3k3r/KKO31+Z1TrfSZTyBmOWJJOG0Urkdu3gMrmSD+Pz
09WDPaOl/lqz7fBis1xiDJhDUYXbRp1fcsv9PTLFK+TV3FQwQMMNU9ydFV5LQx5N
pRvyq3DC0gNjgQuxJ7t5cBLCkUJdwzFCXPzPFYx6KasqJFYx9MRVm2Ue8SVkgelS
WIEqJqi/hb6HQ/8GVR/73DZOxgGNujzVHiCjwszygD2Yt/XmLhfuO0HO17xZOetI
EOXgac+5obSg3k3Ky+zQJLcmX2oCatX+Fdo85cXbQRatcs/fJqct0WhzRnaOzanZ
5y/FZHgMHLmv9upZOE6BvcFNLup+tg58uFzktJgpCPnOKsD8wePVuEeTItZUra8p
J978cPIACjSMlAvIozfuGvLX/C4ajAdvfK1iI/HQJLYyHqa9FvbovecQH/uQGUMz
OtQoWxetrF2IEghcfR13G4Uk1GIDMLDYbQLwcWiYIM/wq0jE/YKGpNJOhI3rp1K7
7LPj0vjeH9/K1h1p8c0yS3eiBxTY8ClQUA5O7OAVubLCbSXf/PuoFHCLLm9Ikver
zMtNpX0/KbDWrfJQqu3oFi9bits/8oafOgXX0hPRazJPPPSFHCcegQDUy5FWrRcj
m+ASj+hcpDAmMOH9s+mNBNrbCnWuDRqNfVihJj8xugV36Dm9BxfUWKSURr3f50w/
TN4ZKiBi0t/cesd1vIMm1Hf14uSHSHdOQJ8yQ/GzzlloPHCxsHQahq0GDHce+MAe
OZzAmordr+5MFDk7UacQRnBcFh0PxZ5OqUbWIq+g08AK838NpfpAkXDaB7vFS2qN
TxpYgw8i3hfK/siXOTZSgqmhhXeH3tpV+rhr8Hj9cNhFIz05zxSU/szFn99hpUWw
5QGO9/vQYoJQqflTiad+CQQoXAGI/U+FK3pye7cdUfYlxXyqkybA77GuwotYoUFR
zs5fAG7u3DGMKaOZ99ZEkWQnWbsA2y2npmmGFZmCflNsjGt5+kwgo83A+pdO/SCJ
2ob2X1MsBjxU7LvhvS6TitLjhxk1pxfL2r/Sd25VshV2/idEMFVle+5pMs/YK5FH
gRjCfhu1EmaFBDj2nO6xgWdgcXIZyeDoo+yrjpwLbt/JMao2gxPTZC9S59Igah7H
GSchDgGCq3k0PkMm6wUVUH+b+bLMaVo4OnSgDOpvzsf8JujcvjctcmA0kdMwhcAq
XJdCyNUQcZq1cbhy9ZtwUNk8F8c3JVq0rNDdxIEuPHfP5Bg8lKLULmcmWfLttq4h
TPI2lu+NaYE2S1ZviEQhtyO0rhwE/nQYqtGKa0iA7DFq8aOte5a4I2tlHwKenHBJ
7Xi4NT/2vpNXmt01vhwcsGVyy6+rjuWN1HIuGRulYMY90TlPmOQpYWnvBT8kMHee
8pKHeauAO09SRLGJeRI7M+u6c8d7f0G7i8V2pvuq+EYUUM/2BzO365i2ZUNJua4l
cmBmuHknDDANEZ4e4Cn5G8iZORCPsNYaoXtJcjRr4U9d1Ln0LODFJ7au/jvoS1tz
nI4g5Q+csprdXe2hm4ORxcOvzBlURJj6W1AIIfZOsHdNrvrIzq+ASAWqEEI/gKr6
nWrcclWPH7FKrvSa0tIsokYftJFNHJg1pF4R1IGfdus0RImPXi8MDngiTkSPbDGR
VPukpvvR+BDU4caA6CT8jK7IkoHAl9Zh1GsBY5Q1RBgJdXWxu1CL5DUZHbn99cj0
+QWeKZpcaDBoJOit+/tMP0tdsw0X4FM34tvqtO09eRuOkcVtCil6xEyGlqy1lxU8
zH3WBSwHthV522WIVD/F/kSuCE7vPpsHG/24olJ6hWMyFitSUjf9MSlIlGW5gHQk
nA5KoGYkXQtD0hhnEl+AGbsdhL9JKT673edWpYIvnDf3ONKXVHumYuljsisXIlvj
1FjOp5r52IUAwzIWsmLujPOHvTgZMuvK5OelX3wYWEua9j/EqQ7i36Ub21OqEu2L
2YGh6Ab1et9/W6TY/usA2z08z5uK1fpiDbNRa8RKPpuBKMXrchE0wzveAcvUByiM
Um9CWtByeuBxn/G2gLg7zwkTG0g0rVOAsvnBc2Kec0xcB2suR6mSae11sCJlUONa
9+4aZZ9yPGDyIMs6vVVZy+6Kj3kYsld1OtCUdiKS1juqxLB6E5WPmrq3p2A+fxV+
57HSnN2jsB701OapjVRlbSN+txTKnfjWwLp8Mb4ZIQz2tVPHg/cTCDskYXxjKIi4
cQKojcSaCdUC/EuKbBNBOPZYlZ04DOlA+/CDSirW9s0vlnn2vObizT3mfTq6WikZ
zpuw7i5AvdGlZFDDXmno6GvxBBuyfs/F4f2J5tOB+WDbLkk9EJs4mQCVkcKF+u0c
9qPS8DfIQBnHqjROE4vLAM8NtBB2g61imYjnt8tiDEMIvFNm+/CnlUUMNGiATKQq
rBR4MnH5NUyEWvYPdVLlNqOlfFWNVmGoux2lBAswo/qNJL7gGwxdP9leCThRjS+/
7wBCKAjgrVOQ9FLoceVSqP0tVMdnYmSFclgdHx75YQLJ+FT5YgOkLCiQeFgqaOov
ojvo2RJ5QdTUFuuMUZFQ8IHSdov5Qifph1aG4o/+xPRuIy61JNKdg3k/7O9lG1/U
2+uD0YDu9Gv3334doPaBdXabAIbvcEatfflSrqwlaboZNPjeDJbxMkH2GzWwH7Zg
C1eS4Owlmh92BZ5Y9NhH85wUlGTgNRYk2jJfxgHjBBOmAf560x0ok6I9Cnm4cM/h
h4rQXmTPSW2r2bxGLRKlCabd45UtmS2eJ5qM9GkZLutVUXmv10g0LSDw6VYDOAi6
Qoll0QeWScAxTMQ3eRdqAbNQmrRxew9WTsE5dJuwnaZrICuLjWutBeTAN7dy9PLe
dTjDJ9DNAbVnZC2T5wUetuFlmZ5SU57mpmFRP+TLLnAYbIFMdsTJOVIfDrvdqE7q
U1XFyVgMER17XaR5Xlq2+dDzkXz4Q+LfdQugPhOVmrUZPDkpuvh2wbwJoC9N/+d4
+ks8S0FtuTPRXqtJjnraIyVWOxmXFy04b0J/fSBVTvdF89c35U370zns0/fIxA6E
Xdyp7hKrTcmFxBS55TM0fbSq++vD4k6TnDf76nGW/f5Z84ibHeZ/FvCTMp0Razgf
wGRSsC6vhZlOK4BbFsdQ982fDE5lOxHh+fEDXICtzXEFHj5wnHBx9mV5WXefO6k5
gfxNL/H7MO1P8pz08b/dmd+jVEmldAa3NGhPkFqfKKE7wtseHKycrSxYZQiWNtvL
EH1JIyoQl2fIoJ3qQoxOvt+BBKQFFqJVZgwQftt5+Ru9c4V1TftvhAZuomJ/ZOuj
0Mfx4iQLz9Vg4LpDo1Qv1AdtuNzr/b9QUezYlMDuqr0PSjUsTMXvPu8B7J9noOb5
AFM0BPKbYxcFabqTq+0RgUoQkxqrj+dmdEtucQvnwA1RwamXw3LGiUH/3w/xjo0u
HRR0tjCP0iG9ZbSFCqUiN39tmFsjXUZPTSooUtgEpXWHOeuDU8ip2yBGPbA/JsOg
BOWQUlvWeYFICxtmT/u2HKxioUBx3sNTt60I7IKfcL58pxMY7TCnhIHRXnUNf60y
IhYYFiU5WC64hU8UK7xd3OK5iGo7craBbyCvIpXFpyCFhk1HplwKfCscFNfDDvio
XhQwJiht91EHSQVl/mRrfICBfGBHgEY2HNYbrMxB3+Hwmq3ZeZTaN+mdg+EchgYy
hzCJtBme9tP6CnLp+RPx/FwhsoaGuvvFaeyxA+yqcg0aL6AwoR+wqHqrSbcFXkoR
hB/2G/FJrXY4CN02C2yTVobZ+7/yH8Tzygssxi6W9dbdCLx9yUXdJHvGk1eNheon
4Z6ljjEt3lZT41bUm51fji4dDDRjtLD0nT4Z13TEjBE39VQtTSyBQnNcvo4Js5VG
mowLgnVrZ5LllG5uOVDWfKaUOObmcS/8A5JYA1/Zpgo6aC+qTN0OQ6psza6W0vzw
IIOjP4hrdgeDzKa4w0YEiMo+84X8P7b4qF8Vezizkek/yVXCplj4OXMup+36sZSj
/Q7MU1CMhWFacJXrwFaaMl16vALlHNmeIkPnEk9PO9OiSCQ/Shen+KHXgqdLRG/n
mH/2I8P5oObfP/TZquonH+q5YnmPGWhQvgsoC0SIDAHYfrRmHNiMAsKeWa2gd4X8
InBUTcn1txoPRdKaQ3CWNYIAkOEb63+ijNZwrvhZYJE0CV/zF7de4AxuOi57bIhP
lezCu69MB0DZiWtxV4apoIflHpUrHU4rBl06P/ARFDDBluN0YT4umWWsxLRfDDMQ
tEmTLC57x0qkKDtRBCL5pO2qp+AkcB3lO047FBHG7yKOlHjlRfetlxq+W6kJQSP6
WRWS6sDuTmxpMNHKbgGNALSdDj+mKQZsmrhSQ+3my2Xmz5jwHdZZ3QfYHCe9bF1N
X4NpCk2VukuQEYGTA9mKKqVOqW6JMuBJOK5MegP+TI/XZhNCGcjN/oABzxmMcXrD
q0BoOovlF4UmZG0Sm0qTbTe5n7Wv3k10/6v6fm2eZ2MaojK4uV+OoegtU9croC9X
nMsELjjgF8bEMkxipJXt61Hh8qGUKvEpCMH7/MbBHjQzZxnAVmG28c3KjFgp9hgs
p1zO6ZJXQl/PJmxiqtva4Q4+Am+m0pHDTTaR0pSayTht/ChU1XK9mc5FWcGgyRMg
Gc9Z6zBh0fHEVQ7SF2LEciuiZFL//HXIEaOIWu++XoQpg6mXNfCI/bUvPTKOtyC4
KuM2JjB4VA/hhvFkSnnY8hrj+GIWTUlN6OyVp7Dm2mox9WwC41LC6/h572zvU29s
NzZXVmwyM7jmX0BDPUB1nja1xCEa8Vbp5oQY4hGHSTB3LewYPgj7WQRombKKAM4Q
vIUz1HbkDSI9aMMEIlTHqIMZx2/r/Vesq2meBpHxE/a5paGu148uTWAtLeCo5Wth
T6FsZOwUzsdpK5NwwgF85LYVkC+sTNaGm5fQfEpaW8DKOPBzuAd/hsrT3E6DZTth
8gf5QOx0jco6KzZNdAaxe7M4CAERCrcglOKj4HNswvKf+TdLLVqI1AReqCnKjGGZ
bXR3Zoqhmn3KX5oAOG/15Uap8WKoSJQvcXKqB6hm1Je8UeFMe8Q1fDSoVKA61sV2
Ds4+HkAu/uN242wy6mR8UhFQkEehSt6VpqjTuLPQAr4ufcdeHKGC8k/0eGo1P+z1
WbgVlNAC+UhL7MDg5SygedYhNkIh/P0rqxIdauYMqCXM6Kgfy8lodKa8IszJ7nRD
Al3bMDG5YHgQlz8K7niOTQ8xEpnNzraTdkWLtexrcPAMf5xLO3wEVHC+edeWhVQl
+laa3wLCRBahfYGghN/F/Xxg/6KaUK1xwcfyhPyM61nh7jXF8+QvQS6I6oe2VdXY
MSMdCEV8XvNr9yJF5s+4FGiyDPWPn3rZMZ/g9LnbFYQh3g7+sVzxmY0Kqa7KGR3J
QWyn7y1WA7JtI6bdJwASeE3joelz7/iOtbLwLSWz4YIJQmuPdf2pULhKxU7JOcqT
OZdyGW2xb/qWqPQLDrwVDuuGIju+l2XV4I1Fe5sA4kZQceu5W3IsV1aC57evANm+
zT+nNKmjNYYFbn0UQd3CqeaOC9JHkzdHlG0B5Eb8Ao9E6c2rpXmfXLo9L+YIWdrM
xszp2jzrvC9bpEgfxO5k2P/0gFTp85p7D47dXbY3baTRCRAgA3nCzC2HeMOr7LE6
wRPTJjFvVybou2kpBXEgD2D3quuOynbEF1vb4vV6ESe+tI0fxJrJ67svVcXyzCy8
kCGXapA8Ql6fLVV4UOeTkmoftcRE/YuvP08jB/O7EAO1vYxENwi1CdDqiZ2YdiA/
lGYMMiX7r4fXmHIblPCia0bN64aiX/c/ksYNjoCvaOcc+dNRorP+VrHyC0hpRQKy
FsZZBy2sVGTO6qaa0JUQWM1pUtNuaqwLUeNYHHDZL091c9o4zKIbg0vllbimW4Sw
lwPa6xHM3vOzVQdTgDaSCnmIFhRi42qdyPOgVOl6uijRQvRMf6V/fO8pKAnG/E7k
YRSVmvfJJcoPURVAubJ7Vj8ODH1mE72LOzu2u9Mm8zzhMPaCHPLJQfPxnUjtHF83
A10ihXhYxJ7la+eA90Ns57+0IBE5Z3FUdlict1LsNY4J53wOeBAL/iBMeFVu0YIj
6c6oiZUE2d9DDkotjIwcUQTVfKzq+Qk/pglaPx/YUORKte5XQSapz7bweFC5AGkw
BAwYQtPEHfPG/zw8uVWrzcAxwmQzoS/XPu0ADm5RMhoSrLb3lt6PORwae54dyd2f
2Ky6v6bC4FKNLrx/DCUdqayi9o+Ki1SiA5AFtPylQQzSHBtXVcyu0bcxOhNN82Uv
re+h3I9CAFkQt34Tpsk+/QI0F70tO5LIH9pz1hUJXifSi9SFKt6ZibB3CoKAZabg
tG66Dnvf5799eliAn42miJbE2/2qV/4aii6aitDFmJ4Jnx/Df4So6vCvlpjJzVfX
xnzk42cU2IYZdw5VKova99USiauubPkYcVmrvNPLbhqq3DfLfOKHsZ0+BoEBOAgi
z511iXid49Ztn0fX4T47INDGAQzi340QcWKnpzu8VJyLSTu/YB0xmxPkxF5jy4gs
34b229HT2ZtOgTunV+gY1CF8y6uqVslP57e+7YCxdb3tglXetOcmMJ71qc/Mj3tb
c7CnJ7oDXMdcOw0kGtcPlSH32Gd0s6BA6zttkL/rgUw6rWQvgewh3DzYIDGb8QHl
CGjNiSyPGeeagIRlRDZDLKWLQj54JiquvtttUabJTtgFtYPuiiz/VN5nUcSsvLm/
1unO3A6+d0p3/rHbuzrnJ4J5fUIqNgvkEt/Hci9wmfGQprEbeaeKM6lCSmNj1MsW
xYqXoVr3NcEs8zHcpDaakC6ZiEdqtpAeEi1hv1wqQUW6MeRYlmFyU15GmUznO/Gw
70hl+QtaQiUSFbQZvRrxhRwFBQr450V1l0/eKDvHwnTb1Cod98bUucfeAfS8FRGf
6ZwfReqPo9gl3hTkeuYhfZIq7m0xi6lK/lHzZTkGrpz+p71057rRAIJ+Xek1LkYl
hqkztIqAWUnJKQH0k8d+V6QqPc6zYXJBZemLjSnoQ/tatuD7Pk5yEK8waJc0kwsr
0i8NBtrj2gGTgdbEt8pur1Rbo94KHqI+2hrHkyqxmBpGdDzzpIfXu+RpNfPtCH2j
5z61K00yNwKGFCL31XTRpDFf/ytC2y6nnhghTG+2DIJKuNTiLrJq/cGTsr65sTgv
ZQAQ7dEw7j+1SmjgcpNCdr5YO1iExWnMwC90xKK6fXm4hcEPRi4UAPNSqoI6NQwe
FEls0q5tEBh+umHt29UnUMiqzev1W4MkRaLLOZ7ZGA/ChclWOWB41z+3qm7EDZSe
lTHWMKYI4k/Zqfyw7AUUQI0myvtBxyjVGjaZHYFrGYWTV1iQU53JCkSJvI/sT9ee
bKo0ACvy+N9n87iw+OrOBXWQ/7Fzbx0lpdo3KgsXPbj1wp77dP4+ZqjmS2nf5EBV
iCAxaAGLYQ0ua8BB3lLcKC5s7tB9PtS60Y842Ukb9T7j6k9L93Fsr7KpZPsfc/ZO
7aFM+m74BfrNONeG0e+7cf7fIhd7P8vwrgHvxvS3RzVYHueE6OFM1KxYtMHO5w3/
NEYiFIhWC0y5xKsLzFdLWL96wrNYuJvIEAv74FaKJPxhI8Q8Je8lnbp/t0zMoTr4
me5EOjKEMhvTfF9fR27IrBmSb6Y8Au11R7sRN8Xta+gM/KQkKTejrNN9dORneUoV
wP4XU0akAYehKRehRkq99eYhM01Hi9i+NsJ+5oQ9jCg/zc1stlvK3qiV5T0X32vD
rN7fpyndoSYqlUT/lkevEH2bvwqLKpPmDCOakJ/zeB17C8cnwiyQSzg2bNwficFs
TGNCMqiXFsYRTYzGZvK8mREAv3alxxyrqcjdovoxL9FeH+/xlAQOidebPCOyZPWl
Rgjx1gpOUTBnDtAmdZhlijX2H0xkVZgo8TBVND5XuhNTbSRuRErVvMycmjCoty00
/ackBZY5HEPsO2X9oFD/vvStvPzMhvZ5/bhajsXEraciFd1U3brF4JE6qZ0ROodq
4gDW207RPQH7mvFjSAVrLa3f6xYk9tTzvESpRGkECZL0QGcf+g2IhfQVvLGKI+2S
zAKFLlX7fuJd0yTdqi3b97vJ/YOLiFLWaR7DR5CZMvF7zzMctmntbIytfVBolBpK
b9mfHPWU3FvuOJkKwDAFb42biE9FIoyY0sL++5L2YZuCLCWMg5yAlIb9ofvTqqM6
5DhiwxoJ40E1nIg4yFDWJoWKDp9B87oOnJVZtwwMiurZME6kIKJsc9Q/Tb6H2V8f
3h6MPcjJQGTXIiZlvgFvv0wTfp4XMHeQDbgw+wvqcP2U8EGfbtjSkNNlPJWR3t8y
IJd6EKNHCmYzTu6udU0gbaoSJQ8IqhtUJmWM+f/Hs5P8lB5vrWTLwEiKTMF6D1KF
9lbAHeR5EMbGUqNfI8APjzTXxkQkRmAMReQUCrYWObw643GQllbYhKBJheiSvBAK
NpPQAg9DT0MabJzp0sQOe732f1cbIuvJYbPhz0vuUgwI4SWfA1KeMBIJCG/+SdTs
YM0618VNQ6ZtFGtCDBRRjYvXH4j69/8v7YBfwOMqddpbnm/kRhLmDMc08ngCknRP
E1VEdCQ07rhc+CGQM2ZSBj5tXYxphid0lkzZ9jAaPrfSLCQgG+xk2Wqt4utyaPqw
Mh/jMcQGTn8xHd/XKMt7UntDbsjTC3lPN37zaopW6wl9R/G/Fcm6XgYMoEFE46M+
oYSZFU1AKuId8kAk/z7k/c5iRgflCMonA7S64ggqZl2KdB/GeDJGf+dL4aPdbA7Z
cLavlAHtT0R+Lu2lLECthF97fOJiIB1iuWZO51hLXu9ZSGgp4LU2aEfED6Hq2evc
cistvo737wOVExIvhUXYPMur6i8o/MSWZvkx6DGkfLODlI70IpsRYSJzYQDEgHiC
QghtjjyUMc+4PjS3G6cBEhyJm9WeIShYhgbR6JQUbHEkJCkp5fNhUTzESq+Tkr7p
2LnKlryi5PLHQXN7rBV7YCW+1vWrkQbmFicd+01QMdn9TBqyrs0WPFIaxcAzZR3l
NTAxvJL7bDSmM8NWsK617K4RtJBImIibHAd9QfUdIn+pwgnZbmvy2WBj5DTsggpP
QXz1gorhcgUY9zugRK5wB0gCmUtDIMQhE/IACcd5E6VhqfLT3AjNQRfeCZsoKQzb
9anMOovHNMckH3wtwxbtxpsNi4ekCn4YXrhDUWjrVHIWyyP1DUmnQ1/6Nxewa3Xj
7pf+t9wJ19qF83pAOb+D1HVtTHJr5QFNb7r++i8do0cRmwaS7FFFwQOs3GcL/SVz
7TD2eQyTjp+ay/S+vr8B2sx+is6euZ8woF6o4BZjTwsypTimbqAHO+u3Ra9+wUpR
DyRzhe0SHNlTmNjd52X3CYt/5ElTww/EvFRr3LDD7zlpuAPsoj8zLM7NETWVFTDm
F6s/JIRBQYuMX9f7QijxwPmjOnJZZadxhMyVHwo9kPkuuylvjzqxQsCROrYAPyCw
ZxvY/Aalu88gPQm+C8PkTogY0Z5cx9IA+MBHIXT8iRuJ7EGxP2O6Hj/ZXH8wXDKY
XORr2ZlvLkmo96hfqsC/vohl5PCHufHVGDBfR+HXDuIrBS5cPaHXRZDd1bRPof1S
QrqERUhsYDVn2lSyBAuWSrWkfqpq8rvXOozDvorp5tYOTncs5r4URZV11yYeob6o
7cTEvmuTNV6a8ZiibXpULolYUqchk6464SufnAzPwQzijxUNbsqOk1Ik5tZGcxyZ
4kkQSv+QTTb9cqaF4m7ZynjZfMBBPi0+O93BtLJFy2ttKr4rMIVpccDDZ48Rr7hp
1xFYNjIlvdlpzDdqTtsapfWaQVfYPxzGKdqsJz+14G9cvQ/16Y0lcqzBuwfGVjHN
v0Hykj3vqhbnvyt0351YJPSghIhd2/s7NpMQMsDJeyae9DBluJKl/m3hkqunzX8X
A2cogu6HO81IenMKTcIKulq8sTrOzOoKTY0ltpu+B4BQ0UEQkYJjBn7K4B25yU3j
ivBRwe3cgk5nbVBAyKIRPVqxxIonB86obo3cBbE1U1vAIU6GBmS9sg2Rc9Y0JcMm
Y75KHHS2LB/70khUjUqNCQxLBKpGWVWUBCY00nTsd8j8b+7laYg0UD3Cp5jjf9+M
qEZVp5KTgZuW5iMn9g2VnTp5NgKa7IhpTTVODUSk1ghxBBAgWt74JfKzkY8a8XBX
Nl1DwxMrSBAF1wGs0emDGmb1AyolnBV/iousFId8JASZJSxBWj7G1ZYbQEcIWvBU
E1fHr1WA7SKZgHvbvevk9Kdp+2vwGFbZWWKC2SfDmUKsKAfgbNa6rxNtWT0QXrXE
PcVUCLq9HR5ah/lbuLYpxGCJgXOIOtTOXKVA98uZi+ewvUl3bwY2FYoDeRoYp8Np
fRjhL3zzFu6Qvmj8ju42nEC1px0vBO+bKnsAtw21brzuj7Bi9GAC+1VhXfqpoOT9
rKQe4dA2SsqL5b4FAIfrKZFCR3IWpwzspKqUwgmgMZhHa00fafznbNsfeYJSRDir
W2iok12bMBcyavxjzicygg4JyXhOkeTdMQHbX/dtzQpHERf09jecVNyl5v7bBO7N
A2dl1s/6t1pwV78jrfDdaww0NkeFsaGh+xepSI2xI4A8sdhuYjYI0BB6pcRtBysk
Z0qu+3TKi1LSm033d3/+y49/XWUs6AiNq4mWyFEWOBn5Y+2pHvy0/8VgyGm5IBBs
slA865I81Y/Gv0vB7gMch8kfDEvYb3tfsCu5qzhr4btN2fJKVR9G5ipsfprSUYqM
HfFkOhRFZBZ1mQjGN2XitZYPVUey9vDLheX8vXyDKJaWkh+15dl5gncxJ9pH5ciq
tup68Ym0K189Fqox3J5iopbROgNcYFwotze2OukYihAoRqmD87XC4IArgF/czIhl
JgIaM9h4SvltSTxcFMqNPWhLmgrFCy9w1ADtY8j8NpdYhgEFiXIYoBU0i4oL1Odn
APbEDKHAVqs7UutdkDE0m+xN2lIyq8Bonm1qNY5TXQwmwN4t9qZygzPm7WwXJGzx
Rt60AysIZH/MblJ2JLV9eyKp2eQ8LmoAclv+snrHgA+2x6E7qQdTQ1KjgACqF/Jy
onoYGOviWpQE5mXFlf/opf3H+ZstEMbVKpS8Bth6vMv7Q6O6WW7OTV1IdM6N8rUF
ojJtxnCGa585w2YfBxbeHeP5PZAnrMbMlZiEF8kLfLZX62wCet3WHzzEBY6miMHd
auFwjcFIr0yzH1Th2Z174HJl/EPvl22F1M1uaqr8fQ3teSbMESlNJ63daGn3fNGx
c78Z6yp85YV2FRqaUME++YA6AiU4qH0fv/XLAXLGFkvUVEaxJPCj2zeFb0XDQy8z
Fb3pjlFqux1yTLW7kiBLYww6p3nfto1InxNp/uv7y4ZOTP7UbRlf9cUUzSIy2Aq9
BzovbPkq9VHTxISG4275d7OURbDO+5LAVWWxxFzvDIA1SXtlAViA+MfBIvcfP+Kj
E/rhUk68FAHVdtRcZLmclPg3pyP1xgOv6E5QHqwWL2p/pG5AKA9QdSqomx80JLe/
pwkq8SyyhV+pfGhd8y+3FnhnaSyiruNYUFsABk96LX21Cm/NBMo+qX6yRbEMxUMY
dtEItBY5IJiW/gy0f5Rw2lKzfZ85dft51VNZDFn+kMIHCnuK/MvXucL64oSFkQdY
rHXuHM/qEm+2mY876mFjo1bv63IRfZWHi3cTGZDg0bR6QPLUTPVVP3sBLdEF2igV
sc/Ti06+YE+UcUyWFXGMv/FYh2zhjQqFiTQYXd25FpkDu0aVCu6iE5x6cSWoXm5p
odfpHi30vaLSZs4K+ro2mxLrm1iMQ9H2jm7U+t0VAKqFt1hich3A4849cNviBX4l
QehCGVMOADdgxJHVUO5yR16GpR5cTFxzfY4CPuqLNlOx3kq6aQsbO/0pe24X6gQp
mgz2YWUgiNP6pMCiwmxYRhVMgIDeMMkpTZD2A2tNrUAiYWL3r/pchfe6PXOs9GvI
TA/cvTMF7CXebx6L2wT1CytdO38tjmBuvighWqDCREws0i3uVhvj4/2fXUxmj5sb
fCV4eIcIno1az3PkRUOmnVwnHbvxjBYMu0q52oQTZkdRJvhnD+oONdE1EavMVT5P
6NaOZ5J78BvI0KPXBLxFC4WANrPn0kgOmYuqwaU+5+IJK11GoZTsM+evhixaQRfd
Ms95+cPYbG/sCQYYHPCdjUYZUgrpqCtFpJUHlD3hSaZmoHlR+lI7OmR7CtN5z5xY
NsqvQFUqTiz38gYsM7j/ExhWVood1po9m3TDNAm9crYoYmgkQfSR4v+58rPdZvL0
vUs7iaVQ71EE2KmSPnCtT9mwqwiFAyeofH9AS81ENJRnR2sklsulqakAvoY5t7Ez
Qn//iCPiB9iKMYobuB1G8pC8Y0D1wk53+3cYRbAUB6NQPkvH4McbrgNUCTy8xZbp
Yc2YJKgf4gC3pbbOqnP3B1tVFK90waHNPSny5wmr/kln1e/jeH/nAulAQJJwreRt
AdN6NVvQIL6RJQ9jipxlHIEsuKwVv6I4wskpZSPCFpjwZGucA5Bo76E0aETQi+l1
fgcPWggCuqDKLL56m69fIP1z91/rOsPnA3w0aKmE1gLT7atzCoYqt1NpISl91KeO
HzSPXmnIftutxzM7HNDdy0JrzDeDnpW6NlJ9FCqUypIqJwbl9/WZO4Wd2w58rviD
P19gsepwYQJ/ttmlbivF7ZBsHaP8afwpMVbeUQS2Iih3B/em58dd67pR1Lfa5Y2R
ZpCaHsfjgJ+Jm7U3aFa1UsOB38eTPlZ1rhjzOU+sUkf6kegbBu5Eb4+1mtIzlhzE
YpjkWo81O+mUq7Os7VSkHiefqfVGwUKnorPCiFb1QBWRKCAGQto2BBp2n5N5T8CN
f+/6+1xwKYV7ofDFEzgDfClxPBS00jvbCrX6vx3UUPux1vHQulPNvK6/JpVwnWvy
tSF/LYwJJ88iFfWGVr98GkZmfaPP/DiY1mGvCTptuRE3FxNc9LUAb/T8CVEKg5dj
w2yFWOlQlyjvyxRTrnohjApGoB9kvmXGirkdZdsZmVymu+BFJXy/vCiEu4ViNEcX
1uDr67YvL2VVYUDlDDAHzVGQ1BObzdbYddur/vohXJja39AzGJzOFS2X0fV7+Tig
C18x4WXEsBPW6etHR5ZIVDQ2AbUP92xQNHTps/kHVqNdwz1shMiuMGHAlW5JL23m
c4W5dJf7QFAErymewig5NWsKBlR1dCyh88VAJxRJtcQ8bRm2ayXMa+jziCKwtuoB
wpp1xz+HZcG016nFxL2kuOJb501FPtioRwsfKUBo9pLaJwMelk0YSio9kYZFiA3y
7BVV698/fEcD51a31DoOMMLIg1D7X7/goou8hr2mhwy93PGI1m3fs32eTDqxsKfn
3TO9QRGVufPlM+qoGclOAjnllHya9+P68WLNnBgPyZPZe86xRW28Y7L2jHnJ1AAg
0e8XF1GmQiZbcuZVu2cEjavByBh+qI6/5yYj9Qc5C8J+Ikam37G6jR0lxNUsyQOq
kTu+AaRg1TNZXguV0GbqoCAR7ZIGwopghkHWTR89DSYboFtnaxIOX4NvccRTaFDN
rjbgkfT27rREuObzZvuCU1Gl6D4I365p8fFnLLMK5SOTLq0X0YMRrh5XmpJh2EcW
RSQC2SBIxLqEi/3aG9+qQf622IlkCxn4uImpnQgiwDx8+yoMHi0/G8OPGxDnb8US
O455zUuinTAU4wJMl3LlUFPHSeJTnR/AyxEoY4sY2szCOfretzXBS5igkYCTcs9U
kilOu7E0bX/trz3YAAuSvWmrGLqeR38yobk2NXC8lwjxKUeH7cNK0LWUYYJCsIaF
qTHvdtOWWVCuHNVLnnFG8wiT+nLJaRs8X/MaAOUC0S2K0cLOFZZMTki4gC/ORCrs
Jqt3Z//Dk0ckJHx0XiMBmgLdKkcteEYhlAJi+32+Z6Ml+rUCb1CdrJ1Hs8K4oXAo
69RTdGPHcfqizZIGfysp0TshWcmxD12hU7ZdpIo76/y6S6vxQfXRJdjaI65/BzCQ
tDcx8QlPQFjdUgAls7IED+raV1EuGBUHEOHG/aZE23YLvl/Cb9Jztmbw6Ut7y5Pk
ex4+MAn0AL6uR5Uy2TWmnaC/ce7U0MZjNxCfi5Jh4PTLn4dQdQvdIHjcOpe3JO2S
QZkLFK1RoMb611fn+k+/EO42FsdA2u7qN42fJG7KCC40eJmS7Q25rbFcmw8dqkcy
PilAPZlqcubaIMq1AMWW0b57izonryidfW/m5sBEYgUFNNj5Lh5nl5/2QYqIFNKa
2bjkeBXZqabi97A4TXHT5RMTMU5nj6g0o5j2US1rkWibj1y+6bz5rZhX4qh1DVCV
M1l+3FTY+cL4Cbn0RDGTbbqlg9lS11BT+3NCwjCUBjyADg7wdu2g7S2x4S65lxt7
RGwj4HdwDhPCO/ByYMbsJkCSssjwjuq7PwIHNlMnnnGBFR0iaVAmWuW3WWX8RW81
X+7fPXlPdrVRbm5iIREhdZZFu1vxdEuAcdLZsLgBlD/nrGWWLExmKFIu3T6qriu3
LD9Dw7/pmTXcK6Kf2TIpbyQDtUfcVK9b+DG7+wshHXF3eon0rdObFISpe7XeGnvO
ouDoCrnLwuDj/54jRmJglOKUL5UxGWgemwXJPpSn3hXHhDTVM8tvdzj7gnDZ0mXU
oLKggazK9nb8Nf8HMq6GwcfI3hPnudUZxt0cZoKxI6gRCgX5BQA8uzUhwEbPDQUu
xKmjsQCvgGlwWmdNTcVsNIEhXxRzJ0gjhnQ++w95w0runRugliYDWnon8MQgEhm9
hWXuWfO6GndD7Q69FZ5wFDO5Rf1JNSEaY29I4/zSCkeRtNlL+GqR6S2W16aeYr4g
jNc+gmLIjsZytfi+VEfhN2tLxlJrBY7S2W9LYIUcqrVqlGrUrQrzdoTqWrnzNcwE
SeHKBXrMInoSpip63ivLExDEeABo4tITd96rTIsrbvcCoCp+nr9y4G1DdIvaGJOZ
ZJoZso3qQaeqzH3/iaWfOB3xxYfTCWrUgYkqCw+U1BkjDc933LbBIyMBTnwsYrmk
xMFRbDiht/UW5XRA4KnfsS5xgpU9j35CFD+/LW63wxsO68ar9oBeNWfeVgmQ4qA+
RzQKZINYgHeO80NowN9zHnRAj7RS8suFnl39CAkGU0RubCTYXM3iiF8QYoo6Y+gL
IXXiLxzXuLBW8mOifDuQ2GrUNxjqK6OCtCg6tlF3vs3ESYGX6T36iAESYCADVsaZ
7KVZ4jY3oL5hiUVQfsLPWmoE7+Ki90KcZZXk2bJgsqL0hqVK16Tn4XFG1jF3iCuo
OUaGDiqT07fhN2K4IrJFQLLwJrigIbVaMUwE9Wj9X8n1knJmwxNiPlOJpBZFFDFY
n0zYgo/34bhHfgCgQJsHgqT7GrsSXDdRJVkOYY9p5sRBbXtZNTMI2+7D1A7n2RkC
v+9Hh+5Qks7/flXwx9BUEJ5YbgXs6H7JMU9J1OjZ3S6z7inzDh1aSMczkt+mZQrS
Hanb/Q+EXHLenJnxWbiltSgx9A73Y+7oyMLvmI3li3m1IhtadVnJWvK65Xc6RX/u
6jzMc7kegJ1w70g1Odj+E5AN3sxFk6lGCEEwIPQMHwkB5ntg4QkSYSD8KxV/uQ2p
n9RX0e7Tw4HTevIdgFyUS3v6vCmK4bZUWhTBr7ojAUNecKzeLpAMoxWC64f6A7G7
38y9QSLK6tbLiC+BTfQVOUrQSP6eaBfdk4id9LGvXIuZMA5ysbauRhKYINaoUZAV
yTr5IB89v4cm6wjplD5V1ptGSKOrsoo6BIwipm/8Qq7Nty4UY8bIMpAd3uL+WsIZ
2PAo1Ppejsv6nhI2cgxx6mkYtfSd2biwr6j3Gg8evvIATqHGTwRcDZnayMcszn64
vDsarufb6qUWJvtFiAWN+OyqCHiBfwPThcwVhDpfoqSoYmv/pcqO/mB88JpKP7XG
zXxrQdqoz+YO0zSGaUM6t7xab89rgYorHHjrEECWNvKgBLZ5TmRdWngkyqGHE4/8
lLHyAeYcCGRx8FcqDPwRSHVXuCkMc1xQDxoeotvIa/zio0xgRGZMD/EDEUz7jjLg
3z5u37YA9qqmRWssw9hQ8BafvFJA6hWUvOfw1ViAZKvVn5SX+CS6e8WGPa4xw5xw
IxZ132oFX0otVRIBHiUx9MEiykSa/eAzP7OW6tDyNTRss7ZFghN0ns7D1emKArhE
Rd1X8Dexgz6N5RAvG6OrV5wTksMBifWpUGHiQiEZjOCVfNqagmyCYRsiBJTSesEP
UF6EGGuy7HYOSAgVH6kLPRblRVQ1Qy1zQmePhQWQEGeD+nE3PYSPkWtml10efMLx
kJIWekqwJCmbtnxVgklf1yoKo2HoXSrwNk14ocUXTnI/gXvCaxcpEXxq1F12LLUs
X0zVzkQuyvpcguGY2V0GftkXwOXPRXTvPj6341f4YjVI3SZ4RTAxK3SFyZiwDvab
Stu4cHYifqtowdC0vM6pZicPr7J/2kqQDkR07WhXDrns/H4U1d4o4umM9LaCH8oE
g85NoA9pE0kZ4lxU0mbuP2EppbNLt7YM9NLrK57RlmBArf7vt1cIXu03YSGOAJuy
RAhezFXDMd3EQMQ7kjh7H92JQFHHen/R3DnuT1v4mIlGBiWcYvCB+GnwD3eQoATs
SRFKcea/LEtHYU/EYgwzwCUtrUqwJj5cfJPjwpFdXdnUctQX/Iw/UI1lyY9xB1VG
LO9ZOLEGAZwSLifkTQGSmMPMzu6Gz5XsC4zo1oMpTZPFhkQJjSnYH86LAcWiFnxL
Y9oQgp+E8JnoWs9Ls5UZOO9/al1N7d5+GXToYiV1bf2qMVZyo9jCgrrsW+llRSV+
GcmPjaeROGiq/5vXtd1fqMUCycHocNYREVMGbq8VOySrg2Mg6zawuCGr5nakaxi6
KC28a+ELvRKFlcEvbFZeCPP9nVZ7d9taPgIbm5K1WZx4Ez9iHjvx6Pl3Vjh4F/WK
ayo34YWON2lnNl4hAfHh0iVCOiWyheFlTcCQTAQbjyLKdxoELii/hxyxvbMtfBid
aTPsbnRKJ4khxftZM4owzpE2JL2SxLaLq05AFQ8nd7tFIHUd2nuXijSLRuRbQFVp
yKBQ8PdLA0fh0FKFMxK0WDoQlfzFD7VKW/Ihk5VL6w/KfcKsQcqEqVAm+k2fkSjm
O7KYEDPQqi84BWBeAF/MAkgqMYERq3KLaqEJzWCSiJyXmBDbeH6tAdeIBsrWdZ1j
q5nDuEPni61ZQjVLCA9XW99rlUUJBg0+lotB44sFOHhSV8vsVV26hDTnPjo3ECaO
8I4SoUwMYaG4faBn9XoUewjIjFr3+VpmlDRKSv8WXbbJv6N9XkmfKJCn5hvpZsfS
2vOmJeBMLHdhDx/liQH7LhctEcwNP6mWMePrSPLar2Pnx8BWSiS3mFhLSodrC6Rv
96fZ2xLqgb7v6VS4N5Fo+Al1b6hufyLmdyY3xTzf3HQFFt1BmbiHoMDP86vjOFVG
WIn4c968c9Jx9wobe17Zl3iTLV2Kq4X4fxr6jIKTJYbTu66IOuYNCAjYh2I2Gi/E
jJQ0n2/T/VGCaFWc7xnaq0spZvG6dXjmKnM02BlzQMBvi48P6Zx7w4UlGiWia7cq
ihr9HWTg3W8J2/AZWhQrTqUPwHtdVnR0A75fiQURuSYKoHupe9Ibc/V+eXFRbXAJ
PPUBRGh0Iyu6UUzEnefIxeXQ02rGLgYeu+70yB6wdRDh9xfxOwNLI2ep3E8ZvIDU
z2uTguLUlKI/iIg1IB8Z423RYAL+OvCxASzVDjtZny58G9rIal1gzh/Ba9Agevj0
kGwuYwJLQUDCCMuCmyosVzg7A6qJ0QbsgySpwV8n6WHSZdv1Rc4ZdpRmvfeIA6WY
3jxIjAHYV+dkXuGhxgqr3TR0ZpeIbFhUgZ7JCMPKHmAvBB7pE/ScQTU2V/iesHVk
NKB0sc7W6dchfSszaSieuioNhuMDxpN5vRSBi2YIHaEfeGBUoOF/ofwzJDnovF0m
jh0GNor26gEAjRy5epLautP56Z6hWregXot8CatRdEiMl57Q48Xb0tRSwu9plUF7
9yaKKWUgYnEeQiuvojmmVdxG4Bu4oTD22J23GhBVqfNnyfPnV2Yary32joSkoP+M
Zo01wZgJrgaLUI69oYLSsfB9HO2c0Sk4A1CTaWT9zY9CZpIxVw1cF91TnHlD/k/E
/Pz6VsF+CGXew5IQ8JWB7GSACEPrzkdGHvZ08HH+SSamVaqrJQC3F11G26AJwO93
nTqSeW+4oSnsACqxvfU2FazorKOP3qLOq4JIY4kg1eyG/2hrYtRji09KdboStQB8
E/MkHxRsOvchhjQjPlPyelpmb4q5KWbCXDi+c/46LJYysmowOeTonev4lg8mJ6ev
//wORLtqwRHfQBwZvrfQLjARWq5e71NMKlSTHd8b1LaXs/x1E4fhywaMjRHp+KoW
uw1NPEIgr02frmZBCPtyqL4jaBQNA0oksuYYwB61Lm/ulXOJjXsuN88iN9ROgFcl
bTltXaoMAqKs/px9rk/EOgLCM4BBJa752KnUv/IzfQQJJddkFRlZdxea0sKPeDhG
sOkpbUzMnvXrm6f1ntbAWTRdnMpCe0sVtnJeF0+c6syiLWUmp1O0Ey4Kmyq+W7fs
tq+EEt9OZ8nEzQdlr621cnE+ACSmDXpSTZoNWDtVx+Hz6nF4y2qd3XN1RhwSPRb8
pWp2nYUikkWTPos2mIqdVCzuUh2QqdKfyQHkkZjPrq+XXhBkg8UvQXQ+RiDehQY6
pnAx8eoKVCR7Y9+o1fM8kAfJMNcQCLsVyc/YTukiTVBeHwhW7QiIQSMc/krN4MxB
4v37rp/1xsk/HCOuzvm/f19hCL62OA4FterV40ttf/1VyhJd3YrTxytCAm6J29kl
EVSiIvhec87+PoyIChFaBsAv1PkcZ2HTTwuzUdKZ1pp9z9KtbfGHnFTwq2+h0867
xj19Kf8mDBpyrPAWQ7NqAzspCE/SGoxO/s8QJbl86/sAilmju1ApMmWTkHrIWB+D
frP/NycajK3ZU74vy8V1tuzSxd8tUP7wlL1c62v/9uBpUnJcSt924nh/urGyongw
B+iiCWRGjF237iIU8sTm33eCJagYvqiiJI2lbkb/j3qsHE5KzvTxTTOYRzCZha5x
ByqAOMN0qKUIUqMf450nfR9x5Kc1pR9ADz3ppI+fjgVJA20NP0qh6hZmbonFDVdY
ACj6lNiu9TFcW2D9OlgXBD4X4OYTbn+TC0vqhGETgAfcFYSXVR5c3GmHKT7oBWiu
bCrvXfjcTrlHX+nJngnTNRjOGFv279OZLx08UtdKIaZA++lKP/zpBLD47BQz0L/U
lhC7HQVD0JDsZ1HyDCuHqH6Ntg8sB4OhkpEJkYj5pgAJmTFS5kJftLgELpRIKUS2
tfpt1z/lDd456gBoXh4prOEkiDo8xcnRVaAih3XlaZ/+BQ5pywmqIO6VAj0vqTn7
2EXTlSBuLJtFC3Uy5t5ZgrO77pcqUkF7Ypib4GLtTW51H8aoG3NpcsC3Z1Iz2wt9
wgU7olpzLNu8z1Zi3FGhVV0x707mMcsjemZz90XzKwTc4rqrDcJtLfc6XjTTBddn
CNordLvJV3WeTWXFKHu6rIh0GxdvNMD5kzL6nmBPJwvXV5ouuOqtzbcQVfWPy9CP
RxUqnevLtvNdSZ2fCMia/onhWvbcpe+jN+3FFAmeJD7aUFdZ5E7h3oGjJba5Q2H6
50dQZJJZKEiSLr9qWOFzUaUXZGvZxKXIUly77gsonvfjRINQrP/dXJz161YYTKqO
w3Fq28mkB1u09qeeYb7/z2hrzh8bMY+6UT6/7mdoRvdHnwO2VMF5hWL4yZR2eFXH
2JAuoVlUwwJCgqmQnOyNlwfyfagNK4P9TmNPEdemOj6vSPVUWHJrh04Pj9LbXF/R
cgRvMp+z9jZ6jMDlHYZdqzjp+QfXtODxheCmx1o2QF+hrF5sT7fXNgsQU1rBDexE
UTny/jQT9qquw5zvfDr4PtyMtLCADdV22TKbbUWiabJlmxhme5bWAjN2+Wmq9jMk
GZ93Nzh3arKQ4LZnY56HtzBkOCfeuuMI7CxCPyfeJ0FuG9+34XTDYXKALw4B+iWI
kMfllStE+6aQjriD3qR3kkYOrfGrJMcJiAAdsuVSPsKDgRl5vX/3DbiOgSxpEaOW
rllPiKxjqpH5nRB6solRA2OIzz+j8wMGN7AIZ4f5yDZ/UOK23xpWhCR4DbXBhOxr
IQXZG2itOiHLQKu3lTaIGhJtAV3yllnJhsqAvnSFDx3dyO/PeFJbnTXjDDyB12ZN
53qCISA9YdgKv8KM/l9EKODi5TRyf0DjOdvqFl1GRoTc2doTRJCFuT8L08Xoso/5
tJjz4eM5HSqEiPdxOPedn9hegy/ObTcxiFlZsekAq0VFk0tJz1Rtb0emUql/rJNL
jPxgqUukaCvGB8BgJh7P75/tsjg1Uaggy7F1JIiRn5XB3Jynheypyw8IInyvMgFS
ND1CqUrbBXUZ5Okk912fpGfYXoKSly0zpmYP1F5IoJOWP/pHVuuX3x0rxdG6lEwD
Jjd/1e5lAuJ+GfY7AEn1JANcM+CY/6Z0CLDr6VTp3j3NL3SYr5gMY0mXXPCFEBiY
fVyHYbKgtC5eWGxKMH8sMhh+A4qWlWbXE6cJdyaAKeyeQczjvdI5B3JLWDgKPP1q
T89u23mtm+eS67Mjkza4mcLIH5aXlFOPWSt5uJTbrT8o3xXZ1DdToOA03YwdyuHs
DH7A+A42BthzQyrPD3LP10XMJIhoNoD4UONSWFbti+C2YBH3MNNojUUfA8z0bPMY
APgezAXV7TGhtTUYlThlatI81F4Wlc00dBrQFeaXiZ25VKbVRlIX4n5H0T1vx7np
ptvLrjt2eWS61jTFQRWVSRseLtL74gclKpm/fkbL14linMj3/D9HWiwaDVSvmEEo
eF2HLn+/wb2FGGKXEL8si/y1l+QzpHiiOZ6yw7+B3QI1AvHNHgk2Uyf1VJQb6Mre
1wTifSwJy1ePuRGuAlixZ32jwX8t2gyHo0a2RDICyLqXTNYnJdjZQ7eWa0eh5vrO
vCrUYdZ/mI3To4kqutfT82WK80rUpDnMJAigxuwMeqbdNtaqTgnvDwVxlltlebZI
MjVH7seX6pp7wY6E8pu00bqG7L/cVbox4l7xGYOA0ZcTqv13yYHvv/akHYTG2ieR
C4nciKPLFlOn62pBuf7WWtMH3kS28TZ6Q6nI6PxyQWkFBXQr9dLcDdgbZRcDzqGx
4pk6Jp0Y5ezmyF2j6URC2rlyQTdbSpGN3NAaqwlL2MYuo+aYE4/uYmc8xF3t/kon
NsRturXcGWQjzfLhd1Dg+jtQHYFoFF1HUHsmFTGZ6hKgtX/uPTr9g0fDH+3r+j7g
+GQSps1epQSk7Jcp2TPjp+qNBwpkzIzUsCPGq6g7cmpioghYuSe5++pmRsQOXQt3
O60/ylOoDAyNDTwKR/nyc7xalzly9IbNu8Dw8zPYlu46d4RvSc0/eY3ZcLEcoJCl
vdWLc+rjwLdL4TBDnOG98rJMJdr/t7fTRg/fkkWRtLtmWNx4JYqR9X7FDM44p9ze
+NxFMRHuW8Xco55ek8oQBmCrWgD2Kv4ytre0TuKF+1qyDAlhFsPL4/3w2ELLgaxs
DR+hedmgt84rJ7oR7Rmw12Wk6KmFpuvpkeC9bW6R/EJITACCSw1EQM7j5X91UoKL
JnYkO1ddy0azLbxsSxC9buK3ccB4OMK/mkkPoH0FCcqdsXlA0jtRaadK0xS4OG7G
GnQB22PkhwBGtHeZebWI0mIa9XlKPEnwzv/1PTWayaTHLuWuoDSpXTmUe35SOYZB
BOHnSSPh+rySVYMUghlPKs0oBHIdaonZkbmRN7fRrexjQoX3I+HdnCLdEacmJrpw
ht6HwQXnSVlbtiWsFl0/gzD252m2WrKpxZNARYL5T3sz9QzLkM8AAtOcLAi94jZO
qwiDwxSdRGtdoWP76+ACMApsuuUK8lP0s0gFql8V1uGlK6r2UpkhpESktT/W2zRY
b90FkBJ6sCzvMSoxLpBIR9Pdc5MRH2t5a6Z47b+h3VLH7lAspTCZHgY0OUC6W54l
emeQnO0fEzDIsI0EbL6VBWfKAMHtR+Xck9ZGW73UZSd3+2/Om5eeG8Ey+TX3dyq3
XnWlq4Z4/nQUYdihuwpvbFCkC/3pimW0PARZntNF0ksgEGluBiULObFqTf7c9sgD
u1GN1b4FKy6O8zkvzs+qemai4YsSO7fAVHlO0N3TPysY/qrhUZy3MRe5YmaejpRE
rgDaQBEfyYSi2Cn60Rgiy3XsHlPYjdO12Ll32VmC2TEAhFzxH9ljAmxC5fk7ZOkj
B8tLTsNgGZNg03UQSlMfIKgEKe1dnfCiTKBMUYhld2abWdHCEQSrI077EZ49KkJO
p5IR/AfN1iXMS8AxvbBv32cXFRhe0roCdzlCBclcHwlbfpw26gXDinWeqyFEbaXt
gnDCTYWitUXjUkc0xhrkPbQFNvOQmMH328mpDFdaWVlR64CFfYJXJlHQ5c11yMvG
D/x7+O9oYYOGGzrgBLs6RLaUOcLzldrhjSfmm0jwpljEiG0Uhq+2Rc3/xzxj9n0K
s+Sscqp20hOpVTIXOb6cnTZ31zoOUCf2hLJrgHM3t5bMF53heCL8zfhvbKA6/JZu
Y/fjRCeI8XlAEW5DS1BHzcX3QPkfopuvCOXqp6v/fYfiYuyxcCZGkZNkWXY+0aE5
QKCEhB4oYV93fmbpFSUHCqWfaLOzUVhGuyW3mE0NMIiJSWXxqAs+COQ2MM1z6nz2
21/EiF3P5V6pK7CijiNRyg97ogpd1f/h0/iPtTazQwmEuwJq97pp5DSaSUCK1zyN
t4c7r/PqX5Gl4kbUxXBth4qknhEfb6DkrZeqzLCkdX+KyLcvFkYr/Vjmwoo5FueP
gHSZqwGP4WbEd5Ew58PqEjOyhnVUXKuu3knyCpOIBo/8Y1NWhYR+jAo3cgrxRVFL
NNJ9FimCzgyhDwgAWqf2CinzgXGkc/H18/iZuETOuBjffYESFA49iwAsjAVyWkDQ
6+BWhZjUiWkB3t4Y8Vy0WPABtvJvHIWD9BlA8r4cRPVCbdptBhXVnhYd7x6m3uiZ
o2s9zhMNLSDW0aP/BdMeP9TkMLdazqtHoIS8JSWzyKBImPE1zk68d1aMM9RZd/sR
6OA9M8F2uGa//XxFb/dr394rNvWTilxT+E2Q9Kc09QdOBCQphVQ9Pm1JJfc27T0i
oYcxVv8UI2TdwulC8by6LcWjijc+UTUS5E+QyJy/y9WuIf4Uujy+542nXIzOCb+y
EIsV0nqEMEh/KdWHqdrDC1z/YHbnB0MFsYTb2XhVmWSfLRZb3yVf+eSlqNWZqELQ
aNeVBYgPgHQk9d3QN8H+kGmpfZifF9ODZwW3JnTeAtf504BPO6J+NdglzY4ffDJR
9H/sISlqejVgrENT1iW1GG4zm+zg/LekuM+XsbPN1WHzzReo//ou4PmcKcDM+yVD
Z4UW8KrUhVYhCdokfxwG1HdNAiN+74NU+vSIwXPIfwE/SQ8puOYURVhxs4hhtnVU
iESAenowZ5e8jk8BaZ3HRte0aQh8BHLgF72JsHdrdLIOy5HxZzu2w+aI/mA7Er1m
+hYONX3sjPfQSvQ6njs1kLUSO6Der4PsEeQE8w/3tL1E5LbfvTPFJ08nCanICsLt
j7xKEAIiqwg8DmDGYxMS4Uytg4zyI5030ty0itV5Je7cy+WHH48HonyivUYOLqNW
+vyv+zdpBHmSeNU+4hunyJ6Sste6daiGE8FGLf0BbQii9MkWGResN4QeGEMbFbKT
dJUl1FQgQH+AFOBBZ5FZYQHNX8J484Q2fiitLj+53nN3UfAO6S7eNzZfNIVPXncO
kWOgNGQJRrhdudbo9RuBnDz9NAT2IL2Rzt1rjiKpWdhGa/7q9Me0j5aGE28byYGa
q76HfhE/yMT9/nT8H6zgEddv5bDBB2/9e2aJ17aQyrh7f+seh+AJuiZ2BPtB3maF
C6Tux14Vl+2QH/xT/uS0IiGHlXmnGr+lND+2wq+k8YKcNZDp7Oo80VH733JgUSs7
ZQuhDzvAS6enxM+94KapADLZ0+G1YwcipEDHW2JS5IhArxPnU4uT1denC9EVIL/d
Ubvb5hFB7aLPQLkm7+3MGhr9ddbYq77XNbmgi+6qnhG/QqC0sUxiC20zRZX5DmRE
/BrhKkStWUcp/lDe4oDNe5cLPwlGWU+D4M0yOjb52vgozQ9lduFsff00RbdepGc1
v8FzGgbDR5XzdZqkYpl3Hh6hFyTP/EXyy+0Mw8rGOak6V14UhLqaWv6RK4lwjWAF
PFNk7E4HowfzLD7skzDUnHEUhk1As8EChUSg5wQ5/3jv/lwYGttrgHrqA4V/xGFP
2q3+TnJLJXhSa9JHTBOSbBkJwBPdKnHfdcBkZTmU3CHGDLUvHZ6Iw1/p51Q6kyT5
EVloVlpdQMuQP3jV8ZbYAYqFDdDUCDPMk/zgXQ8V5e8y9+Mp7eusgftYsy+qgt6F
hwvPXWgJMxUUC92zB7UY3s2DGWIbbpK3CuG2Bc4/iSQfATHfDzj/ZclXfXHBcjFD
pt3VPgBV9E8iL6+gdI7Z1bYFeXUrY4Ir2nbZerJWVJ6Qz8rhWTpGC00z+DQ+X5ZJ
E1PXqGx3F00UqVy8UmtT/eSK/eX+EvomWrEWFRjP39HLnsjHWKrs+2ETM0IDJ+iV
7BQrd0pM+caGqPFEzOsQaMlM7HfMIpekFR/SBmAtPng+N1im8rKsFh0ZlIq2aRZR
H8JAXOlwwJ7brKV4z1TQVKLnSadPErgfojwUtOljvY9HkBezwgHTmBwAHMNlySiT
LZjM49MimY6w3rtQYcQmcfp3RcCiD+/7AW3amdL5Cf/xfopOJ/E9PdSWh3KfSLKW
oKkeqgPPRTGKp95/TLbo7b6LclL5Z5SvyqIP/9l7NjiueKvFpZ4KZJx++omTBGGK
qCn3WqV9HnHYy/OErQMmZmCaCYjv0aLtUtRDGmqTQtydv3rs16Vs/jcBFwufHguF
r+rxouTX4MeOaCuAyJb54rilUJd2L2gt7pceVqqf/GYENSNG9VkQ351p/rZdDKe9
6tBGSNtYF639FtXKPBC/45x9RzOB01yH7ypJZgjWOuKlGqAfdnd77C/wDQae0J9o
T7PYEnpoaxr4IfMcNyBuuMikML3zJ/p+Di7ehre7hFQZbrAfFpT3glbI7lisYR3C
Xj3nkWWHQW9T4WCLvgajT2kizoEDHtm241Lp85ypfGElZh4ymJzGqcGkJe5rWu5D
KSj89q/a7lk8/kI1UaH5VBWi913S+5lpds5vzlXIe3mL0CslQvga9ZibHRbUqter
0JSzkgPniOJaC8vW9AjTLF3dz02KlhUGlEkEmWknehO67TxlBGBF1E8khGmm8s1U
ZPr7ju+5zwP0aTB8r8dXu7zjUUmqQ1ayH2GDhs4bwR7cgI6MdKw6MGXlhTbMqOKn
CjaCcM9ZJA+1a0y9pWPJEemD24pD4QswD92mFIWZA89jPL4VUE64yWSI+2CmOHA0
4OOQvMj18Lpnzs1P21NF3qMG2REIIHqUpZ5OcPfcsVtxDICxtrexqc0QMhR67R7V
BxG2jRBjTqTq+XIO479zxxS2kqz76TuwNNLorhLaWn4GSMvpD6nMQcJ5SpABrObB
tbVSAofGYqjHv+IJZKbruco5CEfnCxnUGn1puAH4lkT6Zp+81QdWhG9FtsgngS+O
OgiDOz0HD8efx+//fy0duesymMaxJ7tbMh9e5DWa6Jqn2WH4Z52lDgG0ep1Frz70
0Qm9kB+E8yvvhMu11C+jY1+sacqJ83fvrUnN9q6xt4X2fm4ftsV6E9VcQPQDud+P
jz0SLY7aKjmnKgLMqY+cCBrqGjOVc/LXmOM28VfMZOk9RIaIrDof9lmS6jgOwb+4
1xPvIN682qXWSdS5T2PipdcwJsaOKmmSUNk1+S3pPPej8Loeh0/PppUanGvpJHUL
+80rPq/iIfCN8vRiCrffOJWs/CE281MhoPJM0VUcYz1b1u4wTKLb47mKDIhs+aHT
U4CpeIRyjTn2QSaHuIZO2jklS/jiQ9cjNBMXoHSvVBjCZ+ajhGQDvLU5yki7eajj
rvy8nr+YiRFVjBf9rZYhfLNWCgOjQsTRW8VtFowCu9a3o/36SCb2M8C+nAgL5lOO
sdrGTzsauSNcuTgyYGNtGqZFzjtHj9IDIsPKeoYs/yelA+nhtywTGui5984ikuxu
PLJLJPBt4cG7mITq+MXfChr0AoYeceeMd7vstX+jHB57IiQfUVRz2bMjK9nxMxOv
C+yBkAmmaSZ6DktY66GjlgWpMIwxkF/DGMHTzRhfO7EVHjTLK7UoegM7jtK1M+Oz
Ay2th0/mJzPctE3n898zPKAhoRbJJ4+mppWDK5v0g0hnh7ueNIrgjahZDhSkI3J4
Tevsq1D8pDOWXq20sUTJ7GTrWbVJPjt2ENtWopA/VdLLfAPV7uCmIE69Tt1CMvAi
ZqElbeaCtYHIIgn6WGXeG+CnoXCp9LSGh8y4/fotkc7bAL1pdeZNxta+ArOBAbJE
AWaJxxNHYcuYTVGWzuFv2JWT4xfozdahjrRfMF5Edat2QIfugdG3Nd7QTlVMzTQj
RvO0g6HJRY4KgJ1VNNZ5d7BDpmEsKMIbnM9KJ9fg+mhalAe2TWg9IxywJsrVDct5
MpBUutzcQUTYhh9e5whVDcenx0TuBkXbOVuuL70qTbdoSHV7VcfwFwuQYAk0TXq0
BrLHP/C9kqkPCU3UAW5jgdjwCNt6GtT+7YJ5Tmqpw1hlepzyR203dLb/zbXu0kBF
yH7mig4foM4HD2IIj3xvQJKWeH0Tevp9/k1o5EFyeKHI7w6g1NEwtTC6Zy6JlBb2
gbYZTg8UNWwsoU/dy1DNRekdkECiM2nx/RAAh8GRrQRjeQz1I9f/UakwX015slX0
8rEjxg8UlmtZ+dIVx10WE2LOEka+iFdrRHwJMeNu9ScQhThKSz3L4DJE9SvuEC6j
JM+xAh4SaPaGy2g2gtiDWXo9mHjOWPQFADV+YUTUI77nCVPd8ZHZxAyxNv5dH3fQ
Ym0NCXmmeWXRi95MJsYIAJIhMvBa2etr1Vpn5C+Uq/Oe8dT1IQ4TMfVNoKsySgbp
2cwkeQ17M1y6sx7WDjLOgzNOEbrHgYco1j8d3apl+ghYrWb0xR42/eTrqE3oLnfq
452b2KRuoZeQpD2gwv14qYlUJBq8jZs0sH2zzkoN+NZn4JdbEZYDL4Z7NGsXOADU
hbzP+rjNBLsz75u1RR6e6qLL/5/NXmc58xRdrejQfJvgiv2mjrE3ila7bA560POv
q82tzZfLoSneai2kgB1SxO3BU3JUzEsS0kournNNJEIe15Pq0ttut5gNlibmoBSZ
NcN1+qQZWqaj+BUkKQ9+4++jRI2HWYBXqNo8fNWEJy1nQ4zFJWLzBM0f16PqkPI/
3Mr4Kwt45+TI4PJDNJviL3eV6T091oRguPmJXIu1FcLOzSPRcGegdRGd4CPXnM/i
DTYzHRh1jw2bsZKpMCzShU3CyGL8gkk9gdGC8M/6mv136CKSXX1/kRg9EWXAGKgN
uARlUkLpzdq1NU/GbeWQo2rTgmX2oY3IQ4Ry+V/Za5hHK6X82/C+iwI1StHp01A+
L+plNVRZn4GdUBtw0dpga0UI0gMLcA0vshbPBrUrwZ3Tz5qHuIdLAtGc0i/FL5Xc
gOy0AaHZ9VGK58xURGM8fK1JUwaVXEhgFIMJ2+VBPHA/nzK5QZzhddorrSd0xu4+
FywLrfChq30bf9I0QnZLMePqTXjiLP10+hYyK2iHWn3NyYvmiuyIwGbBALuQSZuG
ekS869ne6ACpsElwQt02iQpbh3A4yYttYdYHITIqruzKnVfbHnm6K+4Uq6nW+FLO
WjBQotEUE53JKg9sFtLkVpWu2Tsrmospt053Bri5fmaQI4zaN909IL6e/8ygD1Wk
+WoIuroKD+Ly1yHDgL/e7DYp/QY4PNnm4QGmJ6wJK4U+Sf+qSRp3/oQ5xX1tMxPY
LVJ/mUfxd1uP7AYjXK8cIJp3p5LTzId2m9yD17Yu3WfPrfOMyxBDnO6itjP2NwJM
iAP1mrYMQtPa1AsCv980mrTwaP86GVytDJxlf/j/WQakRwnDqMNhhhmEcCqCOAKB
UWWVI4yCYAv6jpscSrn38z8YKFoSEkct7Sa/AntL/AkubKsKyvBcC3rAkFQQ5EC2
y2QbIy5uwQK17Z3C56X+j/ZqMF76NYkVppbynXEeur8DZX/fk00yPueZSDMp8U8R
yp2sB3U9K9nSLq1xxXbCXrKOn5jFOT9wRBHuAX9fuoCeEL5Pco1f+BWbH3qaiGqW
eclAqEWx6BRaWuyfREhydnXL7MGySeGpgXENVLoCy/e7ueUFHu/+L82GtyRnRs6i
EQokc79UPanavG5c3Cc6o8vfm3NujnYfg1kyHEO41w+w6NshZBxWMS8yiOimbIHX
lE4L3lmDaoULn4tYYGQOYqYji0ks2/T/UNPajNFyJ/s57bYXB8Lb0k6lpuDa8tvs
tq8cNiZqOiatz3mZ8tIVL6Dj72kgk0BWmUjTaXmx9spaCgOzJBQStS1o3TB/L7Nd
9ywD68BBAEGpW5dyqbE/ZE2xIxO+CJ3h2VMkNhDzwWZHpAL7aJc1oyFVpP17sBQi
sCvqP1Xc80o6pFogk0Qy71lxINAJiduUMCJbUtlZtsbHy4xU2Q8OOAteP4oAYJhj
X1BT71sDAzObqeq8w6XBZsLOF6Kvv+bKWLB2wdGwZ9m76SD7rQ6n/6NleReI6BIH
KSJIMW9QdEttSdKX4a4XPfFalDP5GcNnBEqfAx8PJmMCmT9yVN++MqqJRV1w1jjz
Wt4e+IZZH/MgTWnBHHJQtlwDZTa0GMRbRoF2+tT1wUMx4eWplL7EuOP0IvD1XQBA
/VA4u+DguQSWIVHKmiOLB3RinBSbDq7WdfDhwUFFYj3d9XrAdUSMD5WL20mhdzHC
h3wEj4ihUJVGMcVUtNtzd86HV9rFSl2XQzM7MlHSUIzmQw3D9dGY6TFnLSaZMoIq
DCbriCck8d+fvnRCbfZOMNDRFKELs3lBD5aoaNM8RNC9sJE2e8sawUQRxduLs8od
aOAHc+IPRpbeMQq63MkRYMjRNFV4FexWEOmrfOtzQmo9MM1UPg3LQgH0DJnq9cLM
YkoA8PW8+Y20nbtLwg7291zZK7Z/ZBHCzM1pqImOy8VTdKBHEWQ0/1NoMueciQzW
/nWSlZis3dRjosRZ00u7G6X01idEkLcZlshGwEkFppJlKPK+p8v5/+zVb4HyeX51
dMlsGPGFO8Ql8jdxEWPtuMRM3vPL5S9Tq2hhgvkm+PQ514MNDEUmutUz6dO4Nx+T
8bN69sXZTbDXtqwBino29NqQLMwT6A7y1RNIfPUqr3oUhv5X2H3KsoKgWo3OzRxU
91L628m1pLpd4ryhI67a/qjii7z5kznI6ld/wuykVEnTfFNOs1KtABM7BvoS85S0
6bqPx8e95PycxyChZil5cKGU8QN2rttsPQBy7guI3jxGfFgKMpGjyMo4z4i9zHAo
AWBeAXVQWT8ysvJ9l2QPRPXa0CipuJF765nlyo31cEx42XxBxwGMtY6hIp9F4YFl
718A6GqODY1wbCY8Ht4VHPDJgZMQe8jkpuG3Udk83W/PJQYLFo0HAgbop9oAZU+b
XwfLusQcTAhRquzUvNUVoDo9Ydzaw/UO+z93WSrjdgVmmHy4FXAR4kXpMSxAtBMO
YSvz+tq2epIa8hud9pmb9+ZbE7IK59W5lTblz1SomXt6tjFFIDn9R4NOs1OvLcPm
uMvbcFChvdwVunGVPDzlG9lKwyKBZK6xp16GuJ2jtL/xOnOZ3Wq5GLQRII5K9nVB
c2SuTsMpuyUyDMrz8i1lIWNG1Pd8/a1hnjEQW9dHWJMSaxpK20vH//PzFXL1IvKv
edhSKJGmORs97ZjVXUkfPwLLZzUiS2SBXdTf48c3ZApnHmzTGjj77PxPt/cRn7th
iyP2/hPxDh33T/NmcQ4xi4gkakr1fk3K9uJe8ndkgZL6A+O6nW8ql6oARUm/3FmV
qZ1soGGtAk3MoqZU+hhKfmCSoyMUvs4zRz8YiUTNDR3rJz2Kipn91sftFjb0mJEJ
g3wxw62voB/PxANoTphi+zqHh4uacIVBjcrf2PBfhlKs+jwtMUTrjKaMc+hoqZpt
NfqF8cw4+RYD/gmoEkHPEgugiTrmsHMuDUOTRCH3HqzNlZCQojKT6eh2NnEUwgC0
gCj8pFZoYemWQlygPv6AAUqA2v2OeeRHgKEmijvQUvHhnbNfLU4vZltH+K6eXbOq
Kfo67RpWFd97YzRzSdxULyedtdD9/USs9cps6Dd2QScCVJANqbRjwsY7Irv+sKG8
SpCMS96zn8q/SZa0VJxWCDCJdYqhCHmoviUMItX2dFGXDzxtPF6wujumSiUg/NLM
LShbCFLwT1pkPwibEvONqONxkH+or7NwdFksTNjnpj+6ZnDybMRMg5R8dub0kEmF
KHWt+EpuuBgLb0OSSzFa+gvUS2okYskVlNA5gfwvyhD8a0IZEbdfrI4U4KgxuDb8
aZgi2k8YQfq/NGoVpB4eSosjbjULo8qBOj/GY5rD32eU4MHakcdFo/+bL7SQpc0K
oD3wgarRZ/dqsNoEjE+w9TBdMoc0WFmoKwwnElb3BPc4iZry9VVvpYIoW5kMK10R
QISgBUI6JRlN+JPXccK8E7l1m4AzpaLA32IvZnMC+4ogYFRVKML+yj9gPiiiym/S
JNH/Xn19Gtw+rYxSq5gfPC+oYVwuvnBX9YXhB0NTfPkl0wr92mrHxeEhcJ1RRaB4
TZvTmuktlXbH15YwmM1EJVaF2NNq2shlA562qWYpSgabW0QgCRONHcpJU4+kXWgu
Xl1AZwAA8GmTC6Sz0mJNgfyg98VS/969qkGZezofcCI2nSGQVIDaiNA/z1SJs8G8
GyAzKHcYYT9Oau9WnJ8hcRed21OkDyDh/DB8BHDMIoOfwT2AVCW1rfIAVjPnrDSk
JXwLWoSY0gX2PM0x7zfeXcFI7y+7hd3NAmowEhbaZnd91M6Y/B+wpokmtqrcApos
oP4W6QZ4O1YdGuV31IQ+V97/wBhfDtR42bVlfC1RjWP6tdPbcsY+6ExzDkAy8bMx
O1hDm473IYNjNKG1e7OlPVGnXYD3N980cjDH0tKgD68IL2tG2/ztqriKDjbVO5zI
5evUdrXNIRE1lZxSVHmvswrpC4wVZri8hu9+Gw6VNhUIVZjinqV55b+bDpK9GpWy
98whBX4+mOaMedfUqmYcQqW6SUB4vH1tPpdEzruB5RF64myHqHnvdO3CNWuzYZy9
i6zgw1EYYfDriKo4QzduHiOrxjBtDwxpZtiFv7Zf+Z037ZWDLRpJ78sYA6Qzi9Xy
8Zso0yjHwdXqBXM0T06HmIOGJXZT0FrWznCJW2fbO3ufeFXwUNLWcooKoGoJ11CY
icyflUIGcs0bRTOoQ7WAfb30onJHAxFQP+dihIQ+dLzqLJ153tavPlkgcWd51Hv2
xT2GrZgzAwsH3X20DWJefTkItENE4Rt/1ElcCNVehiQqKjLar30imIJxqnuy+5Dy
jZawLZwQfLtubZ0bkc17p+U4fBoGjmBR6Zwp5w7PPv6BaH6BP+u/svrvYhOEAnO3
PpeEj6i5h4KpiEquEATtZc+6mK2MS0bvLP+FGM5StrZV4KIM6bnheKP0VJyu0xrm
dT+KBAUf9OWqrHD9lNKlRUyeUghIrfj+XUKPA9UhTybLKmCbfC/Fimar9KyuwwBy
xjTlX6pb+IO4Xaow3TfUScc1+c01vuJJjZHg+Cd+WlINU+sm0jzTFGvNE9vQfHij
GBrJ1EXVChP1/9Sb3RtaGhd5gC0w0VH67zq61QiETuXru+BXx0rT3tLMjNXaE9sy
6AtII7g7hF9Axs8aBShUBedljZ07OVkca5Bob98zjUxF0Ht1w+6K4TIG8BmuQRRf
fkWFNraaYbKIx+OU8e7q3SaDV0W4ZPPmXXpS0hv2H6V+NvNbiKi/fs+iwYRHl1pH
rOMUDDGiLMGN0sjXM3eTnnM5b08ieTNMfIhAQsXw+eOen30BA7nWBtzl0/Ldjy2+
qF9K2D9TI/bctr8BEMnWa6TfjIUwp7QwnCt5LF5b6PfwwZttsi63Tfvcgl5tUyfn
Vn1qlZEGPLbJ2Cd7yKLFc0673cpofrU7BmfZYHfv6Z75mtYN9orlC7UAlANfRVSI
1kKSvpCqayL4BKtex6mwRIxcN7d6PRwUeSWlOz6qr5um+bPHSQsEhVvRk6Ln99ri
q0gWxv0w22tZXhZshPimA/LqgD8SiN32W0lukFOusKwI8lijtO/+7YK1oVBJ1Soh
gqSa6oEypga/f1ubu7ihyBmaF9muVcaTYR5CWWI0McFcA5AkaWKOP5WJszB7dhLO
qSqnQDBGDYaLPks7RwktohJhM+U0Bm0m6JkrAvFtXrLcR6TMHlCdJ1zEsdSoBfZD
GXFsNykNfktHnywEykUwVM6FW+Xb0phRUngc0YUH00hKRuO5E36KRY8u6qtK6Cjl
q2nbtcJbfD6efF6yrJpYTHYqFiZ8/+O1PhAgDgTUm3ZY3VkjvLEd2rZNHcncvotO
QLq39u0aRtWSJXc/lllq1/nvYS2qsWLgVQLABCQNaCbszIZ3e9OwReM0Z24ImrhJ
jzvi6vAWxffoS7t2pQU/DN5ftK30942qYG14hXi2AM3KY2INu5Myakn7dtLplJ4C
DWF4YfLVoWkXhdXkyIL2ADuhQ8D9ieVNjn6S18bghalaxHGSYM9in1xnW4e+BrVA
UdUpi2T+fjVGtEXHI8h/9yTShyQa5cb6Y7U6GluZXCOdg5cb3pe0tYASuUX7uK3z
fjuqy43K6FeT2LWkxIfpMZu9fsbA/q6a52KNsNQMKNLM6Vn++aDvTR6P4HrGFKRh
GIudpLKOr875AZ/FdWyKRJtJnRNqXCGMtn1NOD2O7+xauPifRIBka0McbUnyc1Fb
1t7u4eDZjT1hUYgBXG/XUXLzLv28V8hrS6vhl6Iba85I7LHa6uXIbfxrkn49Tips
872BqAOyEFafl/pvO1FrF2pKM2KXgE4plq3AKpUzCyM7+AcgNhhPyVlH1EBc798E
ykPC3xrvTcAG3OLtdcpUuRO/BJtxOLG3f1IEJHMBtG3sNMb6tN9rB9PmUwHYIbEN
KeRV3jY5Hzs5F+DTIlheiMR5Io+KA58Q9S9g0vvypj7fmnBC+aM+VVcI9dAVT6hu
NXUlmjK8eYF7z4OqthfYhu7foys2aIpDjVilAqSOJoTYJEL0twbzVPnxW6r0GsHO
JrbbQiPjGqcHhkWr9hcdUJOMmX+tLLCTiIl1kfJuktwNkH/5Mp3BgYjjlN8gYrQ1
rtssNdq4/EC1OvWivzDtc9upgTpPqNQ9oHXsIDSUTFT8CzGoF97ppO+fojZDucgy
pqjSvp+u2BEJxKOL7Fn/zuZGgod1VItmdUcMSolKiWBZCkH/uvqFl9H3d1G1G6QD
P06ClmD4mgMhyITlem0vgWGFShGF6qsnCZVQyubT0W6/vQUdqT/rjoiM7OoxTf7F
DIehahWXWFxV8mA2VkISK5mjMD9m/+a9OP4rE3PiVNBMFSI6+zilpj9ubDd9fO0o
rTAusVnq51akmnED3G92d6isM+QhnXpqHAusyrkv+OOVjnKOKISlOkpFTxojsX54
nOU8ECwH8GOIntF2bjfkVkwnFkGsrY3OA820c0jspewm159hsWx3SrDEVkHO9VCI
8QBp7Krkxz0BxoyiSVLHHmpFlgYz9Bp9sHamjlwncAk6WZgZVlJiIMqw0105S29Q
A6/b/oXK8JSni8ciguxhAfYMKpE7Wlcn/bt9Nhr9sfSRejXziMdplhs4XafreQwP
I5uYzQzFQk+zjUiY7NvCln6gjv0YeKTnPdScs8Kr77VNZ1qhHDO/c9DhIh75XAAD
wxa4jLkIykZ1d2eWUzCNw1fPgkEDhM+RXyr+sLBVGGTUEWW84FyJa6qXiOzcsGN5
McUZDL1GWsf2ga3va/xzHgWs1T/asfCWmOk1VoL1CP0K0UeSVB5yUxkRW6MSKFEa
OXQ1AJpHcZYOVThf7iVcB8Oat5u5MgDy0GiBF9I1rWNnNesCehXGH/ecNgpxZXAk
yG8Ex0Bq6sTAkCvqQ2u5JTBTRVCLJNmQGjLDVtH3Bf0xNoBQk2EtH7OTzNytXhEX
tDg9E2549X/10wqtDo4OBtd61c0YRdWMwRzUb86BNuWFZEYY2eeos/Bc9rtrJpWw
4CT7hOQvfQg7hUYUnxuXLXcg4Me0+g2g+VUUNKjqfjsmSTPFlHiKGdNx4sd8itJm
/+ov1l7mpulQCbhwNZErZN7KnRWJ8HQb9eAdva6xFKiQmU3SWwX2uQOgeLJ+q9Qn
I5w9Qxr14XYyS6ugv3yjFTY0v9kCs29uGjmaPgc4bYiYl8T6rvZmvFNWTJeX2fz6
Q7W0rv1dWadxlwmn3+EblvWBy+nEpshuEDRkCUwI1hhpdH8YjmOBJ6Ekbr7nUGt8
e1d7LsCVry643kqKeIEDwczCaCb3vr4nJF8VQ63o4PG2Q9fyRMVcq6fgt48yV+Xw
5wqxChG5GhmmX6BLHn/dUNs3SXeil6c3POcQEwgNulpy08Qrw8fqAE8OcEPUhfcz
SZMr8Znb8mJ58a3PegNkCfplPGYQ/NmstKsmtpRm80GsrosdY3eyrWyau/uBeX0Y
AWyNIKU1sFTflkUqKqstoStk4fzyRGUjfCfHJUkZS6pZlUapq60BWYufhD9ukRBy
Pk9KoM0SMtVJvi0tYX+kgOXvhFAuXz0EgGnt1pn9JGcaecqFkAgNX3L8un3bvYfd
iCChBXP7/enfPRVQ7Ue4uN2m9SYNwI7dxWwvKP07SlN1VFyorYg9Ac6VjVUbUeZV
x1M+BlOrM7BOnY4oJ7G5WlvNVMix42q9v9EmyfrRny7XymhhFpu77uQMGbr8RB/S
DDXgSM3FHGeU6Mtb9UvKXSK9l4wtBEDrch7n2N7khKEE4hyGOvgVbjuB1D/w3+bP
M4MJ73KQosxYydfSb4Ehd5XbC0nptJt1PfYDpyTP51ourDN3C2vaZxGtJFVYP/Up
vb/LE30g9Qp6rxBgKEFmPPhVzqw2zHy061C/BrDrO6TXPaD/dwBHUhFUv3zIjEMl
aOzJFJd1255VcD+qGBzTtx738XvXX3l8IUCLhGQr22qR4EtjcSFjB1l5pj+ZGhno
vYyxTOUUC8SWtS++wsYUQQ2bNlPhx7eHG0MA/a98Zb3SadnoF5cNW5+Jn2OoJzIJ
Z1oIeSe3pDHq5cuHvUsikY6MqES6RZQ0PYIaPKihXv8Z9VCHcwwrrR+YhAiLrk3j
jJgTdUr655KbLqMnJO23gxuWQdgCZSzYYGKMir7TTNBjU9LDVJ6qoE10zM1Wm6QO
YriYZ3F/cwukK5aG8eMYkHq7jSMI4eSghdtGXNDZtSwlq7HFc2FkBs/+fW56Ow+f
OUYp04/MF5KXxWAJ8nt2uHgVR3O3RjfJL52SB/w1MZwL9jhAcz1ygBzwT7kQv678
u1Bm2ulqvySkZ6S/1P8iAbjQasSrEHaYw6idPZk44DUkMk1c91enYYNhnH1hWgL9
Ed3PULmWyZB1QmCmKqvJKu6MhWAGVPPbsPQa0ohd5vAzHl7Kvs3lEfinTvyQ34Ht
rGx7NqCcieNBiwEw0B94MzZjtnGl0EHIZnKA25AOw01i764ddoQYKSqlenIzZpNs
8r7VMv153tI9ykvj4wSeHBAPO7xOG21zLwp3l0gN+DnGQtgFvjPEfz9296L3cxtX
If7r+hDBD1zdcYv3RxF1joRVcW/DvVmO/QhVKZ1SN/xAynpRtr8GI/Ajauf2CZ7S
5MfmbrP9MNCBWjI2VIt87RBJ1EpnKi15G3ZLt3t1ub4woxOXT5mOzRYDGDoFAirr
naSddYD3DGq2Jp1sXgTOhm9+sqOxfauldm1iJ1LOd/pAl/Sgqi7HSXCbWRcpsO0r
Z7T1mMa0x6m5WpNnHzQ66p3XhWwspTzpKS3/+6fV674FyHdwGUfkLGRrSaM3HWG2
BtnLUsZpYJaCul/+rz7EMGAGXDnyXSBgLOSpoe0b9xEbUQF4xbZTJ84jCs/JWB5w
tXFX5B5+ejDZIShQ5LhSQKPQa3jTNP57nopgWf+wyjLWeHMDL7y2cr9GDmnXsywU
nTaJ9Qv3kNlFxDwWv6tvvofZvR1iCVYD6RSqIgIOAYJ5Br633ziZ93G2Tenru5I1
9S5SJIWXP5cNCOU1GPWHieCvvM2AXICshOmLYWc1xtUnZYwDAjDzRHeCf8tUed+5
FiFp80iH86wNqp6l6PPO1KY0Z9mpsk3T0Vbqxc3pmCDaG5juFYBjkliXhHBzuSKk
vDq3CaaDR7kqyDBax3wPvpUqu3q+A+bap+elx0CB+6noZR3PPAvLzUH3PTiSwug9
SeRqA1f21sLgddk6dDnYyVrMc6OQ+k71gmRbiOljSgyM2N9YTCuYTW+fu7W5sLiY
eRviF6Trsjsl5zxM44vAL+dtZN+7YyguejOfyutuobnSEtWJo2e2MuqjOGBeGM2x
esFiZVX2jo3BVV8XRAuK7bCY5AhZSVNq0XQNXK8+a+eie32HoG4/6GffLBT6Q516
kvMM+khO56seYhdHXOWuS3ftNaTXPUfi3Wvh4TARCtITvddo/mZ4HvKwRvLHy9Tt
kdpdCluifPTrI7scYFdB4AOAOgomCL38lDQRQvltK5eazgv4T/mFAKi0ymD0096y
Lq+eJ6D8JRaKC9Sy44Zu2CZpY1j/bQ8JJI5EX23xt0S2UgM2AZ6jrx2lTFEqEG75
QetHiSGRUEwh/fNdhREvHbjKdNNlhKDZdz+J75iZJ61karbwbJi2rZTHhbQCqVBB
f/Q8psYWWcXF1fRzYEHcXcdT5FjxSlN6A5GgDdpsi6V+y14F4uiHQqplH193JiDZ
ag/64klZZtZ+IYJfXHuMzbc/qS3HlngJb5MLZzXxaFWmVi8Bxfi5An1DX9QfZtKM
eMh7MnDzdnCWPqJHYpUMcZv+utRNg4loBwI1BWpD9E9hSahWccQV8zOYbrbzi1Wr
OpBkwnfjIwOHvUYg9rKMNN9EU8OuXMDD6sF/auzbflJidv+7MzFAgYqy9ee52hEf
gRVoebDZSP+VbcveGKvmmSI/fLMiHbtBBQRMPuCE1xymk4fedILPe9TYja26Xqoo
PpeJwKud95UJvpyAK6vD1tHRwSdfupnMK0XUFFSq+0fLXT9OpIHS6d5CsIBSIqAl
+/S1L/E80DhcwxoDmKgoFvU8CsuH8V43+KpF9cCwkED4Jbt1wLwFbKTKleJ0fmYs
fMcA7ofWKDNEm4/kqYjFpHKV/If+ova+n8L7qU24zulScYoCAZWpMyl94/kgGKi1
48My3bBkyrncosfOjB2pIiPgiuk74ChJbJoWcNO5DxNr6mlBYeDm9gSgp0unkSGg
M5w4Yr+H23gNseZND2QsMRWha+TKdkaFcnzoHCKDMnB/ZqGTTiA4b0uRglUx4ylo
FQRbWHdI+WXX0av2eTOxCb68HDeutyx9LsAEQpTSjLt/KWbGg+deMvrd79CWi/gm
NqgnaaIriXWrxeClw9wL89N4f20S3DLrIorGawhNcDvz9SjbJPJ9265DdrUV28nD
b4E84XmT67tQ9xchPmttUXsBzwTZqxJCXNGVyBVvAsvYtf1F7tz8fHp+dvJA+lAG
YRefpBnvW/6z6tOgbCadBPKDoFDEqWO5nE9CbYUUbBK79/HppQAv18WPG6BX3l6i
yUfAHmts5oBJ0NivoX+wHmzRsge7DcQ+P79/dpEhn6wUPfAytLRsy4C3Z8CsgUNs
jbb0XFdgT3VVr9qC2uZmazwMPNm6aOYegLdctUwFj4taDApDqcp724vFJyoPPAx1
5HV/Ib21BZnYVfjXzz/elfoW0dImJ/RlCeo6sQt9Jjf6blTuXQrdbZiAeFeImJFJ
/OrTsPz5J8PXQ/Jd9Dk/vpRT1G5bTZd8NO6VezwnnttgU53RChwPecDhVCdm83hv
P0OVf0/vOjvlwz9kaK9WzGWHTDSeyiiRn86nUmxG9kHtQhlrfdhq7JTnq+wBEx+N
yf5A5SkBfNdg35oqFoOz+eO8SbUXs+OI+AxU2rGOA/CLt0wOwfqtgnZtnXJMrxLV
sx/lk4mPsS8IhEXnv8gPWlgeAxLzY/vS4bEwtd2fwI7hs2F4V+yw7rlmxBMgixA/
qx/Vyj2KDP4Y9cpYHocER530fFC4OJyiTtrtbnm2ln0/camUVwOjK7v4IK/22Kw4
TlpaL0Z2oV1ktiTS4daqJwFOnPexUdvpUW01EZs3quS+4H48BI3WL8mGYYcah80C
11EV4Db1NrCmu3q6YaPzjwDRKmD2MDdBdsegA+AAju/k+A+gv9Y3JHubbi0mXqp8
psuMEPISE+pXscoSso3AzxEqghbhWRpqbHmyDzpzGtw5PEkvoIsVRpUYGqb8nhU3
Rrn0dgpW51MzkMAXqlI2bnWp9AjMOV3vlF/cj1sE9wsmHEyumnQ5Xcr0t2ixew3+
wHxMP8ZYUhiI5CkJM7vcON7omjvWrouaii1mO09D+MHGzpg9rB3ljjbMOQXQLme7
iI1bq7YWy6Emq6SU/Dv5djsKffz23PQWySqfYmPmESgAx37KrZ1r+rNdSE6kaoRj
5UpDH51a3wpbj4b6QLtjDoyNlHtw5o9YACH4VCaWeQmD28f3b/c6DbemvsgvCUto
jcKeCC22AaA5W8ER/RhOZLz3IROjqkwOXnpdSEw2V8TH6yrFhXBegkMLqSj/Vtep
IuN7oxClM3ZnJ4irCQ9X/HkGLr6lUKFGSP3s8tET5k/WH66+OVXTM0iku8W0rfWD
8jkqB7TeGagkE0AHQSOYcUqz86APkL8OGacj1oot+koorXKQBj7tEIgTw5K6O61X
dsSxW6QrjRNsMMZ+Xr7pN9PgDcEfPp6ZJeH0XH9sUdLkb49mYSLMVK4KPttg7NAP
iXqAE0UODhy+VDnAZwQZGil0EnZQ8af/MJ+C63QzGgte701ByyQMh35cs3zQWZHQ
EEiNtA/pUr8Vb33LhDidLZ6ZgkwRUtQ66LPTZ9LX2New9LKKELbOCIJpPaLqv7JW
b1NZcFf4egZEqv4TRN38mslANbZc6SIDvDF3DRF7cge1UEeWLR8MZwF9v3ScCUZH
wLobvCPXRnviGWC3p1Q9PUuh2xa0pICfMZiApZRpUt58O5TyFqLpQTd7qFR+tgR6
hZ7vFn0PUnbsg7AsFGT8YkseouOuc23Zn+zwlz0OxSOb8tu4CCaXEjlxykk346ps
6cu4RTNZcab+P30lho4kNsA34Yp3z9o9LSoo4y4s7K/wT9vuW2iy0OL9kEUE8wpY
e4iIIlVxrS3840RQb3kgu0u1I1PF4a6WLLVX5rEjFGGM66rJvg13l/u3iQPbbW4+
LCdaxuEj/UQL7wXLIVL32HFbPVnWaxGI4Ls0nlgIlG/bgyGbfRF77pHTr88dfpKf
1KPXkzsA3zjrKtGro9vw22K5KbKAVJiIfKJDWjLmCqR4NK+mLuExp4j5xXxnpv0o
FNoWJDSd99QA4OPHivMcKfSdqKAnQDIQqEgON1KE5JuK/xo1ySBDozg1/rrTofox
ineKh9fgGn2r3g9iH1ZPZku36zFa66/vMVWIx3t2iExSDmRnrs0MIKlJa+/kUSnY
VdTULiIh58cGjorTKtms28+PqfwvLVVwVHSaJKYUsxran1qKE/imVU96R3AGgzBo
pVQ1ZHEXVMA04U5pSXU4sv8KcRVH/3ykEC4rB+n9rg/F4gjnztkNc2wjNnR/44Ax
vnwAfaAFM64IiYiTJGv62yTSec6Y716MoJkJZkdGU9DtFuwKKmCMb0pXCAhN3Iyb
sxOIE5U7K3nH5AeseRllGfOOgf5nALbJr2PEuzU9n4ztuh4S+uVTmtPLHGtRjb+w
mPZrvDTIw4MgWstq81PWbzoLdTvMeTF2XrI72iGMAzSmyW20TZlgIz2tIxfA4Vzs
CKTJhRqXFSh8A7NAZgNyCted/OWL83BQiydu8bsUaLNbrJwW2asoZU1OsNq3Q+do
ovmA/CNhXoifas8n6jtbeqnHHxeJVQ2Dk7qQk5q2OlFCeAocGeryLJY82XFt667D
GR05k0ljKBwU69GqEpTKa4/Q6URbRUyVWrd2iGwEEaxYqwGaqZqsFtwyYtib3FFk
niFQWVf2sLx9VcggH1s4XPMgfeQ6fZzo5iKOM/YUGKH2+LYFG5SuBYS4a7axo+Xv
fmOMDaBfSnjczVqeu5KNtEoZBpH0yU+3ePe0/HbvkDgLJ9/EstZ2fUqrUPc1cC42
DCFmbyVQT1klgO+u6njuF4SEoVFpoKRDcRtl+KeIJDKiZcqO71auYNi3J+O415fD
Pt4x3pKS+6PaTLUEsfrueH4k4qZhhB/WpcwggnhYw1nf8o8lNoHejieNc6YkxIvW
I4xAhX3y4cR6Z0JA+0aQH5EM0TumFB81xFXjMZ/nqRLsbIGVs9HQ5CFdW606RR4k
1/NtAsDGv53WDSBQx3eAbDR0Cb4qaJqvMDA/VfU4sRfLe3nlND/kb7ujVtWzUz/P
22OIN0IfbEiEBxu9kD6AOh5ySvDpOLkkXS1xRHq9kLSnsWOBPtU3zl1Jej3QgjtO
N+bKogHfSDJoOjrKLYW1rxA6KyjMMFtAIki6VrVGRy+SEub6YIPgj+8BXnSf6gaM
b1IwHY4Mt0aoZdDG572YIya8UGFJ0kqxn8Xu5DfdS3ExeYWhi3ksC9/vk3JiAIvI
JaQzKDCh+obJ8kyu18J6oNJjv/RziVCBAmNYX+6PwjAVrgGBnGlT49HpWK2EDMDy
TmyqUXGkJTvVHrgVFroy16eaxkG0shuFa9JNJ0WaxwTdFJ/iIC6vFkjz4jDBfYs/
55Nh2mMrEaN6HUKMJEt6A4FV09Azchg5hv6j+v/Gxj3ZtDxmwa4TBPo3Hx5ovSSk
obvKaEAen82zUWw4K0hd3qnvxbVS0HRjkR66fskD+3mu0+BCMKeHBjYCdddY7LE/
cbkjFf11rpwJw6yUBVholyq4ybAxDW73h94rggHR4R+r7jLl0gfDjgTAaPy6Ravr
ijYKACuEsGU2LXSp/77+NZ1S5b1xMkklZEStYd8WhRmO3fpSuGR+rn/L60ptIZdV
MJ0WqOh/5i3skI50rP5kuqv8CRe+e+7aEgwDnhAtZmhsJf5zNg8Oglv9fYaW4C4m
mVtunmQZ6DPnog060vcyGrRI6VifjU9VaAe6HyjYlUihLJP8SLsUmdbDjOIgb02O
Yh6gk9AKOcue8kcO/6LpWBlfWnpjydedA5Di69NhvqIeoHxTHKy7Xoba7MJIinhN
SuqGc0e8o1hMc40GMg4e/WKCIP0+pXi//pKIlNLoweIPFCTr7G2BkUI8OiQ2MI0i
bfSs3P+LJYKSTiOWId+P+i2FFjnuu1IrWtIza1+eiXud6PjeNxKAMN7rfb2GuPNy
bNPb0CNdk/JuIv5mANo+UhI5e7qPu9Ar694+vSYB7wyL9fQRnKQSEp4WhnggfnW5
rviK+RhJ/G50+J0JGuJivK8fFupY0xXrxmB96/xHp6CZe0G15OkHQSNcRTHKt86k
nqIen5+/y6bnhh7x/Uj/x3FCAdrxRv9xVwjU/oc/7osBqJN14wO8mxI+HSwigWbd
lfuqdwmyTtH7s0872AlSOOJIvn1wGnyWFZ6dYrG5nbpAHn1NM7iCfFCsBn8QOjzI
raVCilxlnJx2EcvDTmeEVqtfQElDODkhlNALffFChK9W57L8q+WtOgSgs01eIqbP
kChxFw6Pu2R3WiTogNcgAibFNQw+ZOPQRk1GKLhtEwGL7rw02vDP7LLt9urVngjW
1SRee0WPDkGTLDi9V0E4U22UFyK+ePTTtkP7Lu/wrXbaAzGWc5CXtl78cghYUeRQ
1PFw3jrN1Nt+BYhsRfxLQ4z2hA4pjhGxA1p51bdC2JZlDdvo089Qn1xDzlsQgksY
L0kZsXYyTt3DW8CbW+yA1NA9BSn7Etk+tZDNd7TvoqNnasXlxDIKlALMxZo/LVut
3GqD0s74DkmVFbruPuXZCnQffhVXzZtAhQl/JgUdkFDKPQ9oUyQXuHW7JoAN+VIO
E7QGQMMUx0ANeg8TH7E1NGTYR7ICxKCzmbWLe8nTB0aA++nb7vrH1yejiKYbphXj
69Z784VrQnVgSQcqbkhsSJUJ9MVYsVy6dEKiNqlFiCR43Bpl4AR9fEJh13iPr8lb
056wjl6eoPiqKZFuqWzAOEoLi+SGmr2+n/1Xk59nRO98tHSJ1coth9Nq3l2y68RY
ZOwVTo3jlKAL/gbC2PHtkvAvjA5v81H8xPbnMZUJ2UMo5l95YloNWbMvvfpznyZ6
nc9+upez5JFOPncacws+C/cR7OR5YkyZ4eOdcidejaPbUFpjW0/vgykcxdcHiKTZ
nPSA+b5vshACVi3oQdQnquqXyvuyeeXotAg41wYeUDJqPa9FnMSk4SgIcq0uhvg6
8d/JShSwpN1meE1CbdDxi1HNZQAuVghoB9XLT3buOQNEfy1q69yFiA63jcLej9Lk
8dS/ULZa6c82MJ0w6ZWrBOSkZkF+3ynfDsOAeym/V76B9UcTSEv6TEz6mlqF142l
jlrf20h1GCoV0VmJVx4bIbVHohhw9rJl8703XFj95WkrfOWiJzE0AT7hXOrh/g3/
IwDsxjHTRPhFMDrg77JaN8a4Y4+NksACvT14329EANAMgc3orXJHQfZI9CfREpeB
uyl7PU4JM0mc/O5Wne2XiYZmvHMaRw1tVjqD8ip140B8+ctX7BKfipXZxioMhpvD
ITYhVyTpMNgYgjWRKZcvrgqdM4m14zqFKweteqhi/8KvAFlqjvZGtM1XHz1JvZJV
//tY17gLrjoSCEcd2o/Hoq9Dx4u/nOkuQdpXau3I1UEIgj9UrZWC9Awn2XL4dJUo
U8PyjproEDVcFWvDM8jPUgg486+sAWB3Qd/Hfwmm48w9kvD8nsQ+33wTZ/+GT8BS
LmsC0sKMfOSrImWF7omNqfAjli54kYipeMGTMlIzTD05hZEAuByPcJvm1Iauw6gH
TsW3HkFl/PmkxxF6Yog84j1PHoRDB8GqZKuNKbGYNYI/8IFYBegzbGNqi/lrfdwO
fM2ugazwEMWP7W0nIylho4nFhjjtzw2sPl3VDancFbKWSw87UOWehLqRx37xfglh
eeLMue0QtJPaWFSAxxpkUlw2Qt9PSlZYjGkfYidKr/pth0OpPkwLHelOzPzdi0IB
tAeT1BedYCMr3WCmmFbbverRM6s+GMxKA/+zAHZVQtz0k1AG3katixKRlg8jiZkx
Nn3znzPg1Cb0+EeiABWCjyXGGM4BfUWYwrD1cTnEe2nLUOcyUjIPHqSDTFHpuuLe
OhF7acuuYAUUH6zNcYIaE9b/jDVqUzi3rG0zVVfdia6sW3+jqJF3CmvySI5kkpbQ
w6epDwCQ36CJ9tzb2wPpXtkdiBk/Slhaq2tZM8P3tWHvJgHuD5m3LaQRM+26wWrO
UG9wCRO9RFpCO9+t2t0Ieg4bhH5SjkBioS5Pg8fUcZUlxh3yU3qeYUzgdfFjeANu
2PniL486K0eFypK75fVZXHQ3UVbaaIzx3MKwHHssy1347Cew0TncKNDzK739Bcd3
BGME11MQIidLDDaMoZHfVUtOfe2S38amSqFBE920meUveVnpB0P59itGNo0QmNH5
oFP4eKbkYS7mklyiqoExomDgr40WOIk5+/ZgsNINt6Wv0QetmMh6VrNikj+fF/sB
bfRMUxCTxx/Y8D0TRMhMIM04oVd0NmT+08IPNyO9MTJu0BO2Vbk8mCDe6u0yn8gP
iF/2NfB3mQru3TkchuW7G2GYilpJOMrvrNJzxFfLxc2w4JYV1re/air8NONoPKKj
LDC4xKVbB1UO3D9jVJaF9rml7rmz0tFF8nzzLOQOCs+l+zTKx+PXeg9yCO23n4Lr
/SQh98MoFwewuXMLRYOZRKrjxIQsW6UNOgbfIv9cz0GpkogIaes4TztakMAqc2cF
s1660saVivJ72VwEB2+Qg+vdAgYJy590CkUP9jE3m2jUki374UR+EMd5SDuw9n2S
7RBnFXbh7MDIZ8K4ZCTvM1L3HVAYyioUugx/baykN+F4vjg2rQyZkeh5R8cv7Zfk
jG8zXyvHcK7Se7QgWIE8IU+tT6b/w7FvoK8XQtOleqE5Iu1xhpy9XQK89y0Uf3re
Oj4Lu3KDEAoMZVH28tdkNfiV+IV7dWBIrE2ICA0cSzXIf5Hj0sTEumu6c9qJ7Ky/
xq3nEnEXUQ5qLhxxdxxLl1qCKq1jZhqSKtdJf9Sh2rwvTdDcAorKxeQbhIv2ufPh
4HNOLcbVZx9jec6tpiPV6OlckgZh32efHhLfdeTSNdd7L0AV79/FSEsVmQyDiW+Y
WOvrnEMHdb1GQ+Hy80CtKuz4wOUusVl1dFNPT4UB8w7xy7NKJNRENWEv6kfB4Q1M
rA8I+mifBIyGyYh5kMvBDHSS05lWqoBeTpbIGXW4CI2Eb/04W/Y8F+jLRkVWipoB
TOZQwmxBArtP7VWWa9tOzwpTEo5d7HQRfxxmGduq4TkRAMKt2qfAJVUN8rP+AZf4
gAWQQrB2gE9W1CJr73TycIO8nGyI6LtpMJcoGeDqSWlGcSAp35Mdy0VC1QRTcify
qgLFarVAj+l2xcnp6eakvoCx9/6ZTsEDf9gZCWca8c9C7NMCUprVFM0k8ZfcvLHw
Y0miDOPLsuBzN0iATCylIZtmUbhoqS/HVotXvX2XUFU0Sf9MshLo8jFfSsRsIoNM
UW6qTgBCQzGvV4O4PIXfRwWmIwUU6BsuD4qONMScBnbjj9TWt2DiSa1w6uRepOg5
fywwuubjY1ELl4aWyhE+RwUJUCBWgkqViPUlW0RGJE4uB1jRJsiEBlpj6n3vVbnU
XEa3KMSt8hjdmVqQCC7Ewkyh7/caxmjoY84e3lclgs8isb0LYjUYnHFkZcHFqHs8
J6Zk7DQZAZdXocz4JJv7qEhPEVz77WlP0LgKJ/P3rxjJxBsd4lGQi8TCzyuc98Sc
0DIuZccFJB0l7FG0MEX+N2aASU/SJ+3g2PUT0isAWd9z3w+gJc9GrNDGx4y8t69h
/lvi0CNRKpDBbjHFK8OCfxqiuJRRnersP8nnzAchj367RkEPlPcbWbl+EhhTE6Wy
5gdgglNCKDNozuYyUImOnkG7qFGtGFzA29tezYGILdBE47s9twVYHBMjnMR6sqBl
uvDO0HWpfCnHHLqwVRCEzgFfDkQc50mM3dRhEvR/5jMkm/VV9mXtY1WZkUCsj8ue
ccaT+f2BZ1ypZGqExQr8YXb+1TZPlBn0kHwnxUTib6XPh7REobk86OGnQu8QTEvq
TORclMBKO6zaacMGOP311Uk1GgUh4HbrD/4P00k1ozNBe7s5dZhEeqPC0gUisfTg
G4G0WcUlpVt8EhIVxK+3R8q3ujylqB6cr/ddrFSWJRVSnAHzAomD9IxMRcGN+cOB
RN7E3NptnEpLjsFCWLRpQq49sOZiduH6Q3o5hZ+CmT7kjcWs7X/8bNHLmPoL56DT
Y71MLL8LZE9YAjPMklKyps3nSDdfpUpS0DZZjlSApmydMZ337NdlajuPSzZU3dgB
K5SrFKSMA9Ly4PJ28VdA8SE6J8eXEb4t8ej1jNXcu4/XE4z93B1uqSbBZbOQl76F
84+iBVqRNXNnv835ukUWQ4LMbACSIHnp8MP2vFZPBJX19zet67SVShgjuLJTIWXp
ZR7y3XA9rSm/pcXlOTOxDhaMnlXFsRzKI6rQTfObEN5GuyTZ3jK3j1IJDFMOyGFU
yiaJUrOrKqRmwuNW9Dvhc+veqUfXDXKztgNz2Ho+ceUb6j8tAoh5621PD1c7sicw
uG4EamIcce1N0EFiBzl0/WEMC/Oev0m6/tSIYBN36TdGpQWP1Hclif1y/v3Tdml+
llIrtgVvt0Ra5KHAEWkoXNR37h00crBGbrDV3N/7SFs5F8nmpMomQsT+NSaQDc2o
Lqncwliz/nZ+XaqQhIT0BFiBHyjLxOVdI86SUdRMmioLxS4jXCHe9KRIFHk51Q7g
1MRpRuMny+zcwqpapbRwCirorXdmPbfOpRc1Ce5Kc48VZnkr0o+xMy3S7OgBoKwt
Zy6At1XbAo+DVAIgYQOUXeTwahkByRKCsGhSeeKsP7x/B3RQknt6bsnxiysltsgZ
2IL02510FFOlLeJweyE5ZPeto2tqQ4uW2MZHctesoUIEA/clAVyANpLPXsC9VPOV
LnnyggSfnaU7hkbIeZktcrhJ8mdpKO/LsgVRiE0fBMphSQPj397rLE/nNCkMU3za
bXjfLmgOGAaM9AQ33JnhSJdrtQYIJhdgoVh1i54QEDT1xZRPtCoTRzuJ6wdWOxU/
pUJulEjUqMazp+GpklMK+NXk7a95PptQiPzLF9h9/VlDi5oBEt2PxMTaHzrdNGzY
VpMx1cd7Iuu2SAGZzlY3WYIrp96V8Lv2kRJ8nOd0cR4NON44rEAtsqtmhhZuUMh+
sebmp2bwf6oTyllCrvnQX7q9lSRW9KZpiY5M9/IaOQa3NNOLT4tSDEVRR9/yASM0
GXcB8KmZAbkkRIE97pg0HVzOvNLFmuS/ZaHi1NUaCVgRBAhKZtTBPb2T7xZ7N5lY
FrKzXigkCOLKSL5ihRlavyoqUgsw70HVrFofCpHiDRkYGDQaNlzdc9+IclNTFNwG
AlLVe7r0k8gbq9mugcBJ5Q7+Fo7rB03bVDr4ad5FFDC5GlgFO4wHVEzqsjWQIuGI
5+/eG67JdKdU8jVsoHzzSBZDstHAv4hY2Wgy0H2IBVSJ5w2SD9sKYHKT70PVj9Cn
WT1BWdra6FxEjmgTKnnIvC/3gDwXxobsiH+pi/HeRyZGapyLj1q8wkqnnNlX3dk3
eiS85BvV5Os13ur6V8lEi6Fc6aJrD7G/nNreybWrJGKf3ptCvSt/cdtSMe0V41l0
jUcJE7ks+0p3aXgg1SM9FFr5Cslv27nOW0UujdV3iQ6UyuNh3lMdBlQCnNGl3Pvx
M4nWeTn/ruZKUEtOcQwtH3ZJLzxYum8ydEY81UzWUPO5u9C9kPaPZ//4BDPLg4fu
Y+HdXik61hTeXqOdJVJo2jevy0EtwsVb+ay23TMzI8bPMXjyUXEVFFNvHp5+tH8R
KW639cqnU6jwod4zLEBQ2KIYUK1kx7H0+Is80J6yHXiaDnYgHcIqGm00aCZlZPJ9
djVR+2VO7SADIejpxQ7N+N9Lh/YuEc9XSYvWf13f4qZ9ZWQV6l4Cu4Z5OT2VHMCT
dfP1VCDwNJGJEvJvr9r+JwxsyugrWUpzB9dASNjJZWI0DeS1+2JGU+DwIfGUV4RV
eXAqihcG7lBfx3TF9j8EHvrn8MS9faMqnhStSqqg2OIaL09dFYnXXc0hxPz+m5hh
i7oL80nEzbmsnY6XpiNKmfn5cHy9aL0Lmxu8rwIFcqM4RyiifOOYmgP7kY/BeRip
xI60+iih155qw4lD9164TOTaGbWCIF7H0/oGloRrCjJp5SPXFsT22LWupc3aI2Oi
LlQQNa8zr8kWxas+wnkfs9ke1TSmQ9wphYcAhm94S56t+NVqvNWpephn/6ZSARzY
FGMrAYQjBzZt8UlzpLdMG3e6nIcA/NDJfauY3C3fZUtgwjnUKg9h5KoKGVgh/NPP
e76pMBWEOuS/HZPtaQqqXPX0Ke8oks9wPXghpdffB5WqJvusb+hhNrh1OZBQpk7D
yQaRcYiVbwtW1CeLKiMplDCxnMOEtwSwpkQqsDydYyp7tqlJgjlpf9H6cxuWRpFZ
Mv/UdSwMVtEp4FefKrB8if0f5wAxpsDZUOxOqGxhBSE+ZgglPhXWq1U7x1cYep4+
PEFPhnwsKN0sIujVtvNAdcejz3/38GjV/6K84ZK5cO1m9hO6j0jvhO1UYQPf1aSk
jJK07B9n0KKh840pdoH2hOwky5xcyp1QdMk0Hg4nYd14nAgyMIrHnsy0Dqoywm9x
SJWbXlJa1koSds+caHfFSQPw0XATZNXmqUpWDl7s6qrHGOpb1irZa862Kb79wcXU
7pg4lud/UdY40s0myFW6lvnvSxKHPW3qEll1kkbamxnAtqNpHj3LKoybNfCHFzUv
Df9cQjD2ttNK7ZrKxtQ1+G00QBoCndwfFZ7wpzx5Sn1KHslSSImiZSTW74eYaAmo
YNoZUVbDxg9GubexOg18LFsTz2aBHnf3D9M3wVpc7E0njCZ8bYr/evIK0cFZzWuQ
buhVz2tt68BfY+ZkMDyY3GGBYKtp9VJb+fB8tXmkBt+XvZQzYEd4tDmNmqBvcOpN
3dpai6MTETon+oZVAPNsCYlElyQGBSSOvI2Htk/JP1lHXuXOAGDftv5Lr9sQnWjs
jXO8fWDiHGWv+aw2Opxd0qcxAgCcfmEXsNGiLrXirPEE1y7NCOmNbI8ZCeZKq8F5
fl3kg6iz3aaCzbKYpgjmbpb5LDQDCun6dVBbgZgLZVFhc5HCWrZyjHo8px4h94N4
46LzNnOpHyC6lbPzOhJcvr45QyviMtrzK6uPBpF8iViQSPylNUJLwLYAr7g1lMs/
9IUdWx6JCfzgt2P8nuuRqtoBQj/FlE9gAT6yvu2YeVtOWB3Z2obNqwKTTaQpcIEF
Zv5pGc1rpJi42y5qh190hGL+KVFjHzlCyGix1xLFtpD8IEhu6idsFItGr3L3vhZi
o9eNYULeuwOI9w8yJgvBUzMmvH7M1vnd421JvELQR1XBBf47pq6wY38xvEPf+z7e
SzV37Uwo+3jkP/DECcw649RQaxemIYT07Vsuas35fz/S4uoV5NYGHb1FsaWmbnsO
LA+tQIpz40utR1ju0b4+O0Pkxbd/HFybca8Jfhdrlt5eyfbvR6MDHqYNPaWUD7Rd
zAc3RcrgsiOtFqOcOqAaaJmuLxXPazRJDVM2kGgi9LyQFdmgR1CCJfxPPwdeYpVa
DqnHmd/54zeeERCvPmf+zM+trzOrzZ0pgFU7jMTAwD11Wz9sVauRd6N3ZRQz1Dk/
AxxlPxUFqFuv+l2hKkeVq2yWyHBFaivf5KeRkca8RvmAmDxzvlXR1J40zA8lpbgJ
icq0ZGBBvkvUf2yae7RqYhJP4SbPTVOmhdF+Z1sqpJTs8dYAYDE0fdNjL/vYXZfV
3LOCMO5kTVPZWaNpMjhPxc45kIdWOwVbjBfA8VXByNkdh963uQqz2potyg9WkKYD
jmDjEhauT4HwDEWFchd5LWRF58bfqgQ7gf2sQgDh3mpcZbO6w367/Z0lUNifa1ZU
BB41iZl9AgonG+NUDjCTUROEmtVfH9aQTaFFtsrEto6eDiU/rNE6uwVpJxWDLMGr
TPmzwgSgRhCTWRFadgTYyn1WSHcEHvAhtJxyKVDO2TyIUCMTmjy6GpTwBWqYfpCp
ecZudQmE5lX5NsEhRxavCdVGKXEgtNYDY62eq1GZDi3gJaTGqjfcYYGskk+yVI5d
png+XCG92rZJ873g4sHHhdhn+NRSYTlMgEf4dcrl56MyVRRWj06n7wBTxWuDbG9r
lJRAeIocr+kI4RrDjuxCsTDgX6hUs5rmZg+FdGhvLvrF/Qw+spJezqhPhDb5JSiq
YZOKY6zBNj+MZG67jYXQmyHrZtmN7xqkRxxmuln+XYK0eVRneXIofUkMtW3IOE+A
QuGHo9Oop0GN62We2C6vcl8zIwweQr4pEh9iEMqV4pOUaGbFPCz9W944xWnzjPD2
1VXgrwfmdlmGXJwN08cB0gK3xrgz/2LwuBhaBNr2Nk1AVdv/MT5815G/m9kkv0wP
RAoaGhmQ2Nym3CKkCtl0jKseemOyMIAakUIFD7Uw8zoeUX5MSTCzpkHLqSxNaijL
ELWf9TzStZg76BVgUVeG9KdCO6vvLgZ+Qs5hwnQzN3XKHLtT2y8C4s3jisSdX0cV
1/OK1CG7AUmr8E6Vk5JDXkv9KyaypERdbfIGMqddiBRevf7hLHqqYi2DQ7NrC4uH
sOf4uHp8hm1X9+wWWML3wT2urTWWOE1FIgvgSBrU0TECs+JRbp7q65UrGRI1C58W
3Mtc8mMx8bfz+ph93GmtowPZd65zzA9JLj84iqKqNagznUN+P/rV4CJdKl6mFt9+
3dHJfw1QxZQetKPTASPtaW8CuDbBUZMfRfTaK4p/y/IPP2FTwVroGOlCKzLGME9p
D1eDOp37O637MD3VzKl5/2FPD61K6YeCLIppVYHcJeHK2f1qNY8rYdFUx1Hb5MeZ
nxS7cUU2N7mcgrvXTy7oJM2Wk6UB/K44P0fmlY9QtAIEDGfYkV55Tr+eLJBg/QdD
InzIXj54SH79v8B8U6zqc6ZzivpcilGDEunABhsqYn3tpCEigwwsv+Lx/Iq6JlhH
0du/rJhnC51BBKJ/w9T5tMQzXyVUpjkpPAzZDqpaM671taz05U0jfv1Uxh7VBvfT
3YrUNay7XL2C4NzdYwc8NHMB9LTrmXd66JxM+LEmheFVpyFcz0eLoeJbPKhNZdSB
m16mWQWt86456m4hRJPLFOla/wOOj6BD4coV+1WTBZAzuZtlvm/N0ycoxw/pkihr
avwAPsuvzv3hv+dnctNL5ll7ZGP8TFwQCGIfw+bfnwcAroGA1a8H5iI/5Ir8uSLG
SuIZaNV1iBJB4Wjlc6hdojLzN+DUQMoB9RO1JhhsC28Uv7nl/CuOjwrTiJCW8Nra
q/pz0txr/xYBYJfodXeoKBtxZc7VK7m5gL/FfzLRQAzMXCf3xbp47n8M4eC6pRtg
qO6SeTgUXyf97g6Fy2nDUOzbb2PhBYZlKvMPh0Zfude1r28qqzzDfgh06yNB0JHV
mSQdZScMmbXlRg0V93oBsswF0g8oHxQJkp8jo3BDLmB+WaqrRHGm/QczGgqaYMHG
J1ElA/8bbAevreQz3pp8MxKo0Gw2xwWYp7UlAe2R1MNzj/UCysYpFlyDV7gLulIA
KMJ/rlghD06S35RmKDQ/nqSWZ5RvV26bedQdJg8JexSIqCHSKqMNgB0xP23aEhzx
Bhz2wpzMDLHUIxkgu4hvLhzE7v7nnmNGO4SIGVHjK5UlmAFtm7P7rksoPvd0z/vv
KnzX7Oo8PcKo3Z5eSWc/GYyK9lae0kl8bWF6rQA9akL7vgMcd/wEncs6wsWLFNdw
m7lx1fgAuP/ZKzNq57ZtrYXsfysAb161xGb6tWlt6OWZCtIo4Faor5XctjyTX4zn
m2Yn6+Pg4AfsPfx+aOEIxr4S+sgPVerDPOUhKmXRFKv1CkNLFSLgsbiSpJSgdZ7r
s+BPx0+keUsdbDEXAmM+TY8e8TamoqFS03SHaIZY8Ir8oit6Drsdo+NILUaWtyFU
0R5kw5kQtk8OoSxvmlxK6Ent5Y9e4OL9cXI+M/nLMz7I331ITelK8q3Z030kYIfV
tWUNzkzIVjhJNpbO58DLq0gHpcwPqmQAiW9NmcSZZrnqW8kQtxdnjY1eqggit99L
PFVoayPYQDfvpQg+DBwhocY/95adV/EWVTcFxhML2qNNLyuVC12dHk57z5YRdIEz
NeZJZqsA4fNZgYATD0f5QJcQo/KrdOeHnmGhuUPxBN+XyxpnVUMEo/i65/iqlMfr
dkcMSKfrsN/I22wjSVoFPj4s35z3Z4kt1tsU6CChGcY3e5oW/qbuE/TmZuzy4Qwk
drNNdmuQcsCZOzXfeR/8h7YQSTBUt8VIwJTFIAw59B8hu3iUz/LzO5edxjZhkQBC
CR5doPFBfSy16jARBeWevfmpNGSDGEbiTOK1IePggxDbGdmH9Ob8qalNvl3JGscp
AZrTF/5sOeaKJFHvr36vj/NNrxWZyyrgD6Mkr4seUQV93b57apAqnf1aMD+NgTHd
QtWL4kMANp6mX55v6e3sbKk2MR+j+IMKlfy0tGu3JiyuPeldPrKwtZD4AMTtFksL
JNQz676hFPMLce1xRr9+Gnelqnhzcan6W7FE4q4mwjc+Tfv773NbKTHi1wgTzG+H
arKD3F+rTjPiRwYAFUwq7S2ddmpKh+AOpTJcj01CGSi817vV5SNdL0/Tu8t8pSLT
i05us2hY+bh+E6a03TlwNosqAU7PN8ZYjTUaiLtBGuNzSv7guvtjTOMePoTS0PLx
ydnaYYwuU+sa6BqSCd5Gk/X5Z2LQKNV6nQS/lZQDMbEnx5siAecjR/AhMWgjvxbG
6G8vZso8LdSyCCPt4maD9MN/ojmDxwLQrxEC8UoeAzC+DU97Y+ARha7VvaDl5Fyh
hpJq14t91GUHBGB/L9dEVRpSGPa/WPQOFB4HkHMSUXLA/uUsunc7sd+yeAbf1zpT
duPWGtP+YDqR6lVoQ0BUqOVPgouoKBCJQ/X6QwS130CnOE7eEtkJ6mp64fTNXF2y
vDlrqb1Avp08cEZdIZGPxF7uat1OSgBs1JHPGaHQ0wvwVZ6z+6ndLrl1nvScraaa
xfPEBAJXk4+dzoRlUlYFChN/mPJdScR/yeQypWaSsodKBGXio2quHRXYU0EMsTBD
oA3rOX67Acc07/pYvXW5rp325Fc6VxAMYqf1kUMQPuNJb1mq6SUGdph71nTGwjAZ
bJVZUOu/Wf83G/6X6xjHqIrU46Kp2m5YONumzgns4tmWqkQHcg7qwYBO4PPxbgSk
7LM+nhdebpOwFs8MApMKtHmxW0k0WCIBJYuzpQfJD/dYdCcBO2jryixZM2pP3f8s
rdsYxexuO3Iv9HsEUz+CElrXN+0046bb3GWks8gyZ3XK0+xCzvVfDLaqw9t3iGDx
+gDERq57WfySk5vwnOVZFnQ8BVZPfs+HImhqAt83jGEg2Sma7PmicIzOw1JI5qv3
dNbWdoib49fwVvgF/e1Z0hHU6yv4Tk0ZG9+ImHPerdEuEAQ9M9oG82PxXTGG5bFd
Pk9ZxEwKcL55ISaAkyGHPqwkM5ecqhDImYvNpgTFdQeGuIoYL3Xw5Lj/o9Mf7T6s
aUk3HyFgPIKpmJwnWSOOhW0J7oELNZNjqYH201ATxSx8IaEHXQqP0nDSInbWgwp4
qbwaWgQbYJ76jFxjRsy+VxXKUJ+ATyKrJE5E/rVxejECxAbLfJL3wFnN+bCxDbbX
5pQFepbRCrBIpQrJNqQbqu164fq3WWLg1hX/oWKi16LYGc4uPjoLxWnGEclhgyZj
XunjTKGnPNF5ytlDXKBR2WHtw0ave4IbeI9jmcsnvrlAjaxPf1cusyIroklKQj/i
7PQc5iImz2Wa154MrdVLeqOdlPsDiiSAwNioAYnFwoAY28xnEf4YsftT3f0Wx5O/
n85qI/k2bNSTXg7l5F80THMk1HF2bc3E6FO0blGhcSLkHm/Lqx4Mg68T5Q6N4df5
jvLE1n8rtD3hPdHvud+mcW/+v6i7Uhc10q5liP6NZONB7rR3qnC49oBjI40Ri+MH
LpVBCFXM0RG3sZ6Gl8B4WUpnDVkUY+bFOBLB2xsZVc8l/ab8K+7h/T4DsVFQi0PP
ZzkqasybJih8fzFUYQJoe4kZcnVWBJjrJbERKW9iEi8oixAosoE4OKYAFIPB4SGa
BKRkB19ApE9is7MZGBYIwyZwVt1RP6wq/j2tKg1TBuIdCqT0oyGlTKkm3gCtt+ie
25MMrc/E4qGfP/mLCpJDk5B8qdHpPuBviG9MLLGNZOOUBQ9S0vfosO0RD1D4AuOv
sDUDNNpOFPyhJP1CId994LKJ86TpIbvSPzjBA1G5QUkaovV8gnFiQ/oi8VA7PZT7
4niHJxZMqHDb3c/fZ+PUih1La3V0CGO8NZZBE1HJmxmSQwImP5MvoaUv9QkQyfpq
c9dJfVGxGHpklaZYnFpdmmLrs8kb4UqCuiF5srUhAVV+6yM6C0xpCWVseQVsjexC
8B1BC8sd5V2eT90VOkToHY6uahbbq/ayX8T3o2/C0tQNypw0KNf+4/55gD4ur+Ya
HHRA0oTf7zo/1B69Moyh9yrAGRR+kz5FTyaCSOMxi+Z7/6IWnXELWJR0TMP3WCXX
H63yrsKZJwgrdnUDQ6C4JhX6QNCANUEOq4ws9669T3D8ZOkSt1DqmaandepR48wF
i85jzs2Me/akASxfKDEszzUo8ROYWWj35au6Y9fZlgllLNmOWakRTgmizMUyf5ZR
a/J5GidB6ghH2Yr/88JG3P7MrlQHJtrDim43X4s46d27Y+gX7Z0pm0bTAKhzu99x
tdj/LuEvCymjzavfF5TH5LHUJbL0qpsJJOk8P6JkHkrMLcgSLYACRExTX1Msax8T
bg1djx8iluD80e68sUg5UPR5OKIs+5QN2yPdYawg2zP7UiTCLZlNwUunUgF9bk2m
cgxzmU7ywOEMBOCy0Xu8YTwpwqAk9szRkENmkpEPwawZptTA6RokKudQErZCJppJ
k12uaXAjfMZGruBqHrkj9vTZLjpjkbpn2oXQKUyfRQojBsMWAxV1NQlmRJvZrVzm
RT3LM8+GiMMp2urEq8vb9dKG5NvYD15minewryrjGhzMfY/9xYNJUA8lLFPv2dku
WGGm5ZmTIdm868Lktvxaqnv6s3dqNgjj3CljFq5o48Z0px7Lg9OMLkHpFSpsGbPj
sfros3XlUxhadqEU4Xx6Q+oiEvLjmV5VHBNvj7EQLC4ciG5JCnASuO+Ne669ZHEU
pC8qjxEkxoN9tRqT/j8LZHkjtjP+8TCH3E1mcLMvfKLnMIJrLTrlb7wty7g4cPVB
fuQpoOU4qiFDtqONpsf2zOK28af/ekiK4WxKnd1WGQOMuHgp2nBmIryAe8i9MRMa
yVdaKejxoNvTT9waVKRqJDnqib5yi4SJOjBw35t9NcR7RN7ybIpqFS1aNC+S/EjH
gaN/DWG/2cT8vWnF0p93sJHsG82Jgxz/CKAWGJpf623qL1tGXM8PB/Wxj2yCFCsk
W6N/HI/ieOUgk0Ge6ElIGJ5NnviYtqp48PUxdBkwPv8MifYERMCpQ0u4omXZuO/8
CKHjRxzhKwPegu78YhKcNb2VGhrm2wa5wyBwu1arZOCmUNITtRA0sS/bzIS5NIFV
JhOE85HjTs/RpDEKP7mw1ugBo1eESDDUsuwDqfU+W9UjSFWBkMehNdH4mFkXpuRd
Iisjds4qi8wCEdEssT/4sjIA1WeocobHEjRMslfRtrkpg8vvHMJlfQFMKsulwWG/
qU8AVLwiYc2sB2VOy5X4xDRQ0Vx+/j4ZTiaEYDV89CAY8q7zhQNtiATzTwcIn0y9
ds/sRMXzlCH+Lc5II8ciZPWnlOYGuiWweNGnMY+QMjfn/mwH3KgLhvjd3UoePdKz
bfsg0HzAGFrfPytRAy6uDS3X49LA0hCcOlt0xQ+zoL2uDM50mqBCMWSvVGxsPT7r
E2VQFCF4Tu7gwEUExwG46kDviNThnHjjD6K+7AOhUi9Y5LjkWw6w8eVOT8PhivWf
y5Ahy8euninqVRyFB78RE7+CNuAJFToVF2Oq2F4XKH8UtS3eUscqQh4oZVXdwd2T
ZcHIMGn3d4uoYMx0eHCE93kjlaOR7j/RQDhWIUuL5cT3m/G/y57lbAPUEArOSLx/
mo53kVE9TC4OudkM5gOn67IBG3VHK7QeWo3b0FyavOWSqLlNkNjpjTdz8+G7JFCX
lkQDayW9ipGepZa96BVHGYnJRd3GNypY2pwvIuWx6jVem7ecxDVl4O9uQ9C7mqL7
QlxxiIAfBQcQNz+VaIa6uGj0ZI0NBAdegyqYxJvUGqVVf8tvw+Wpu/qxqieMQX9t
rkbrIjrXtSDFb0sctCKFAlsJdvEPVJ+l6q9iDQydT4GPoXMlEFaWIDAHcjHQs1A7
tKNqvP0nG6fSw1HxSa9/XiqXILXuZM4ge4KQGhnNSau0SPUKH2mQt84jbbxkTrTp
gWSh+Y9+K496SNYQrua16E2hekZMKzKzcbW3ZP/mb7onrXMo5TEFH++Pc7dCKq/m
ODxRr77g45nR06+hvfKUg1kxa3Pl4vfKT58nr8G0UIgMX3yiw0k2z5Sm8PNDJtTg
erQO7mvHY126QdzZX6LwgIs4BEqOlqGYT/IvF8oSO18nQ2KvDvnqSjn26QEQpSVK
Sf0NtYh3c8mHk2qnKoC8GvMbEPi1FBeyFcDW7fNwipDhz73RQkag55gt3SMq6GnV
Uf2x9M3Ty109LNU42i6e/RCOiT6qMwHwSqhi08+WweabRJPvz1VWqSzZoBBeyofX
JzTENa95oC5cEm4mUiU6Ag+UUlB/rHJ4bvSwNuKvlpWOsqGor5DKmd3i3+XkI4kV
/FEbO0z9hQ1MRx7BDIHvI1BoAyKoi/PH+lKeERWJBZBrPx1zGD3MyjqHKxQf7Rhi
FVPQnGyEmiOYpUZl3BG3dpt9NsO7CLKwXDEx+zMmBWCmzf5DfmnVaAtIK5+sVN/h
mrcuMSvMxbBjInDnnx6vfaKsXLePjr7r4JWeVeMvmqR/s1duPpl8/EGhJX/l7Mgt
rID1TJHNaCEGDc8+XKsl5N1CN+h+26DqfEvg7l+/cNtRjJ8Ms1R5YoVIgsLE91YM
vmD5CRXkp+JlHzrj9AAUb02wUsPb5fcM8jJoiwDyr90KN3SdNIsUJJl3QVQP3zb+
t+hgEkSZQgq2t28iMZ6//xN9v/JYHTv6hnhhckYJJD/s6NbKu8GXwG6ryyWYZKI4
JtKWRkQiTEepypufyavavNQay6m37OMqwGiLz5+4aCN8ZeAQunm9W0ZUMdKXsEb0
iPhcCs8pqrLB2zrgpUabMiQHZeEI39G3ZNvUKuGXb0AZ+p8IsE64j1YzbsNSzqkv
0Z9sEyOsaVPY4BJnhB+tYbrH3NygDdMvzUO6buS7gISWeEMMNW4vU5JmZCQlZowd
9X6y0BzWc2O26oCcdJ1+TVQCXEvxt8bYnmeEKU5xn/bM0wnrgeUBYMj6gvSLjyqy
68LxmD2Fq0G69iSv7/v7mI1YBi8kpOsAFLxc1DVoj5cEgLo90qPzwES22N6d9eva
y1cIXIBbMn1ItjxxIG9hWl0GgG0NQpIEWRlq2pM2WzKuoCciI06O+3miMSZUrbRz
Y23/zIJ3F+lHvXZ1tk7jcppKX6cv5KacFYqlHjuI1cI/c9miSwDZ5Q9AT/axB3yL
2a5woxH7OKUvu9i95vTr2ZteYMqNt+7L+R/SicE25h3uvZe1D1k1Ls0aUnXUVTy5
MCf1Ej7zo2fqxkIgngPpQZYiWeeshdeqcdV92xlMomSzsXXE5h/zCvxFL9aQwXaH
PeNGI+GL2VW0eOJtSk/NzkE/+tYTSD5MPoRYag5IjhxAX/KWz09QbOHYignCApCc
ykq3Ab5Wdv8D0qTI7G6BFQ1LQE+YKmiP2JLFDKAfOYvOA+0Ta2l2YrNAigI4ZrM5
YwUFo7B9GKomScRgJ0ZRb0JMTBZWwdy55KubyuNSPwaTNqay9nhvBSBydlxLw/j2
DKsezQ5bL/6it8uWglxqhpPv0vok805qEgyxn/6ZpccmxS/z0zGftef6uU8aKCvc
QpdXfM3RoWrcYjJtn4xyYzRGCVjtPPd1BXbsDLLlKRjaw4Yb1p0fU440+B4eR3zK
R6GauuChJ/I+9Udvl8nbliLaZW6F6xplYjoAQKJMGAZUeNfWsR/8aRs0k2mwnmPi
JCJF0lqkBP4kAuh6XSchGOq3VUr7/kuvwgwy1k5pJj6Ft1tITPyAX8jU1G/lDwlK
pLqbXqQllY392qCa4CYZHMWapWxIFRgH9kj0EmKGzKclZB6eZdyTuEKE8iLLMuhb
Id8yWZeHj0ecNGts70t9Vy7iLUam0Qij2dGBsJ5kx/578yW1rIYEMsvufZDj5old
asdsm3yaKxDdPRpyqwFrVkLOd5gyBHKWezZ72ibaDnYUaignJjmlF0HqsxL1gGoq
6BNakGf7Fi8FAP5QIL7fQfC4uVCRBVsOy78grXBc6qIBXWIcumZRpR2dYkd+IZhq
hqroGPxgAoLLUv662brFQ8jgssKUFHD7qyAI9OT4hKMs6jIn6nsWhbBGUJQh7ccp
akEXmOxobxyn1kQ+BcGi9xkoxST2kufbotTXiaCKkdG7X/2toph+uh3HCQtOMAXj
UDavcAsYazgzLzFRbxrVVHyqAZBzWn9mD05b9SXh9eVBK+5HE54+LzEFeq+LWhRE
KB0SNaKFmoT9qrutW4LTJ0KkWcXttqxt+GBpwDPAA1jt7+iAnswksRBh2E+jtuyM
Q46XfhOLBA7pR5fZtXkcvkV74CHzyeJOviCyhr1lYdQDPQbHt6qvmgdY33tQ1lRw
st93+6YJ+QYw0eY3vXaTOj5DzXAbDz+rcplJvff5AP8556btpFayCbvp8fdkjyjE
5TBbCq9f/EWP2MW24Bx79YHfMbRupsvxSIvbrRBOGm1rqssDVP5MYOYw24Ywmh+T
2POD2sWT1y5WKxishVxi6b/32fsT6wvdiB3T+7KqANWomhaSMFyaXldbTpT7A79C
XltEGu2gnv2HHP7Hgliati+uWkCWd4Fi1o+T83NynHDmEQTK5hyqIYHJ4dKvinOM
2E6YEtLk0SGlPlvviyjaCPxjW6cBa2LTEf4Ws7i4g/VdNAUtBfn69QJK810WRmJj
7XcV/vd7NXhXBO7Mesx97Gmo2IFZiWjP8uNDRJWwt8ysR0V2/kCDVireY8ZDmP6Z
AJNKzU/+CeJn3DHmJ4bMnmwKWWmeYuBtEwx3fHPQZgKTww1m0erFwm1MPGVMwLGD
pEcBah05tUNvvRxlcbMyXpMSXtFfJ/NMmfrL/V2s7dxtkX+yIAIIQlZgDCLOQUiQ
wycb4ZoI/9wE2vkoD3odiAKKwQZaoi/ay9OLCio5nyWTNUxoaKerHxsBfD2Ane+q
1xH7Au7ryNANCVzY700M5E3vQgh7zabNm5O0iu/8iXGVREexqQET1mG8UXHCWYjI
mPWhumN1QYt0swUKjNUSzmLhe4fE3A49XvF/MRKToeLryHAGbSog4d4j0KaCKwlc
OqEWwcH0vkYZ7bTybBW+3l9ByI0Ojzt93ZKaoFTQzPz3GvwHMk+QeKJBLy4xUuXC
qXox7fLGIUKq/hHWdhwFsJM4CIs9PFABSXvXMrKfxdLw0kvkI0uhKqjKOsmkLrWw
OY5iYnn2b4yhVW+3VQImsy51egyj5SuIcBQ204wz/RccE/i7v+RXJvfY6eS99bzM
a0+8VeaFUlfzdSzQiw94spwZdBaANzbwQp3MzH/dPaTJ1wfDBnNiO6xoYmwrrV2i
hLXWug5c5NgnNPXOHgD1Fduqmf6LK/s/mq28Z29lTF40t5TMKYiWxRCqHgWZl7rC
qCZEpM2PtuBU6hSuCYlDrVIzNrxtNKFfs+y/cZtVbKxoj3+TfQ7chN8mk0WudSXE
oEZl8RD1GWSmgtxAMfMZG+DfoAAxY2aqWTXg9aFmg0WZK+Z7z1gd5LDVjgzBz2hY
mJsgOFgsX64YzbWNdElw8sxMGBqk3atosZi8IHJbrOXIEmJmyVAZAm53nfwXLP8l
Oc9ZS3Y8qIgW7R74x/ttGE1RZYcVF8nR0szUT3NMf+rmSObmm0cz/07NNGiLHUFL
DeWJ2HIu04nG4s7kKkTlvM9tMqADypeyVQQt4gIcmwbyfr2OVsNdiXxRJnFw1OSk
rwAX6Z0ZnIWDoFN+9a9Mw84MOMzHqet288m1FX3VwMpB2juITTnUWTLe3BXKunIY
+jD9+OrAYhAcnaGmFIDhiz/7mqQTR7RCTSaYQ4zV59C3qq/PE1tez8oNuWdt7gJJ
VzJnCpIU4NojZz1OlVEIzSMeeuFKcpYaIXVPSPfCIJkXjS2SqXZTn9xePpuqSl7i
V5A7+nFm2yRoIQhkLVo622a0z5vV4kjVHGLTZQTeaJU6T3SVnetGi2bQ3nNrs64j
XKC/0na1D9Xfv7NbUZ58rxEvDQ613rRGH9gM/wwC3wQK2hcJS0dAcnuIkML2Ooue
YtR2qDdx6b0/LiHiXy+2f0+MAlJz9XKDRIRTTSDw6jhTf2mUSipj2+dO29+qymxK
4lTJl0pSMonCzwRLkLokBNpsG7DF+WEoQEPQTbGc7w0jaVZ7+S/rfkozP0PVuYy3
cmI9fg8Sb4zPHeqGt2cBmuUStZyDEbzegNrbU8+6MzS5JmBroEH+ookGYpaiu7kH
dEIUSSOvRDs/FaQ1My0lXMGFSfX75a/4gy9WRqxShXv/XITYeeKErvqLtqPG7WAx
nNL0YTaU0mmfl/NOhjaOjZnlnIJvWfmefETSafdoKRyJBNV3/zjtITfFyd230pKe
7wEbpRQZwe+QA8nOEbc/EaJij9qE8a5gH0dF6SubNLQYhXHsh3d5bp+P8spRGM8t
ZZLKZzEhbjQc3SgWcua6HYLyJD5SVEUX6CLov2EJ6J0NzHGUnLz0rYXlH+pY5G7n
nx8Nc3hq+hb5y+iLNFpvOtyMkLwrgaBRsRwcyOWsK1d9/Yk9xC57RdWCiJELN08U
pBI0cCo3Yh+cUyYF3V+uaNfFDX7MdB3nfzwuVL7nN/dJVTvrvlprLI5BP2x7EHtG
d7CGLS26xUg4SMg+ce7WpsK+mulRxmTpfGJEMz7CsmIIUS6a94Y3kXyl0iZMRU/n
w+5eNZUFP3ssP47/NL1TqvF1k7z1+WvEzJkZDwASnUooEaFNljc04OZ5yR8aZIRN
S+Nkswwq/SsYz9N7vnguLj2eP/YdoiczHOq8rG2C/rzWsYn7m9ssz380JAvO6ros
p/Q+amq+SQcyzZv5dPokcnE4fMSHae7RaomINanGz1KbWVFAFaVlWZvNDvDt68Ko
aEQZwbkcWpfxbMnG5D/0scCxyE5WEpZfLLyejeDDZhCqq3SsXbvs2qjASEX5Uqe6
paFHFhpcRAEfIkplpZZ55dbFdE3umI//wTBRnOSUz//RF9tKyWJuIhKl8doXr41R
TQEOgKnNfFkGfoPigfPZhl3pbQy4hYoIaZWyjdkJxqa2qlObb1eiEKN9QsXRb5AN
HYoLn+ChXFViFf0KHxZG7WMHhXvo+PUpcDYMsnZw4MuElCgzY2oiZKBmwPQN+k4B
b8nPnxMa/kIOz7zjjDYA4M6jdUUaIHjzuGKjxUNvv7DFKp+0bGh+uMwmNpoyQ8au
cX7cZMyuv7R3DNTs15+ReyMbvLacigy/H/hl4H4MelBRrMGsKdeRwar59XL4QdOl
IH3LDIxzuJf0Sw6ADoUp1hGWk86ePI1nbWcb747Ajq3qaO3RfLutSqrES1vyg+Q1
cVpsJXB6R3Vnz+vbU4TS7jwRi2o0vMAMtdbt/PEMlBgFORqG/6Yo2di78oDlCfji
QhmezX/ThenvKnvG/wohIZaP5+D6iiuPfs5zZvMToMe1zfycX53PZaH+xFDqBjij
rLDHyys2J9JBzn1q0CTO00lLu/AHDHoXk+1ad39np4ZmyBYjBTlagtQTB7OUF997
s5RxVnztCIlIqooGn9lC2PSSZfipBWT1CnuUXBrZ+yJrRFAPQaD3q/7KlTN6MmjF
v40NrQNuRvk2BJK/YLr/9LfM9CmbrEENZpWS3ueAr7+iBv78WnbFJh7XB1GlZNFg
pOHXPydcMNduHl8H/snag98YR+/x85P65gC76PHB3bBedzYyytREAIw+0ugdtWnf
hzHw763KB5WqY/hUY1lj4UKXNqNkIDXVmKg9QQUm3o1rWvAlVokEdmgEsvgvJsWJ
zDGClgslm00XyFYZKLJnb6sF7E+U71xJT00aZ3ur69WmMq2zyVhfGdOZmEHsvFfp
A3fXC0y6V3F4QLlT2KVGJuvpdx1roEmgl1+O4lI1XyoZm84/m+a4O7ddLhppWwQh
fhEskd0l/U5SzLN7tnxEf6rpxKUDzARGGFFO8gbJfcPanApP0aCr+YpwWu70DE8/
2Lj/7n7AWQscrPXL7TSzg7RRKHwUv8TFlEuG4tI7SfwyRB+rv7V6NYsvbkdWkhyW
XyS3EkgrsXvodT+uAVaGoSm5QXG37xA13/S7PkAnke8aobH/sRQQmci4/El6k7Lx
D13uHLCn1tvWquEd2s8z8geu5b9ykhEPNww4DJHucEoHvbAb7ZfRWG+0riKJ7qT7
o1zq9eW7M6pRCypIKWhEa0kx+ah7LMFwcp0Ntaeh5KnHkWg+QGUWYXu8IWuyi2QO
LG17HmrFnztoWzN8TTDKE8wMRpTSnpYhXmgGcyvlI17r6FAeoh98+2aTt9MGCXOd
XA5BAj22g7NBQDykV9K6srzEdbOORoNkR8nlY4mBzPqlAJbTr68LjDR+NR6Wu2NT
BsabNcPcFACS0nTQ3ZJHswxKb4L5F4nrN0AyecHpAWEJfCvwZL7ECLV5dtkr3nm+
r2RYqZLiQJuBDgbNV8PDV5cd303C+5seeXkHjyv4LogTkcU6CMmWQCe7YdrQCBxI
r/f3IT/mVN29txvUeE7oLr5KMNsF73UU708FbEC2dlv8ohfFyV/n4p1nQXIZbpZ/
lAB0/5xM+RDEq19jseikNDAenNWZNHZZzNmDC5X6nUG/LioUUOBetjF+it3u8nX7
du4MSdALuEzbA17DbgLCp2D4lY+XHK5Cq2D1sVuPFHlryk/qo2UlxRmLjgYG6KsH
1s59ARKMn5rlQGbBuh1CQiseLyI+fjEu3fusiizjcGdNZL/IecMO8t0tWgYvE4ig
3hNO8ZaccKi13y6qm9J2nDmo3Ij4Lb9Jv6GjoEb+fjP2cki7V57QPcutC3KtfdSJ
PSsfiRA3ODAtQC1bQs2f+ylzphnQd6IBoKLEn4AmI8Vmfow1KgKd5NutsuqOcR10
9SrI1sWop052BP4dYbJVOrLturek/O68mSP3KlohSZfpZUentflRtYywnskH7G/i
8LdisqwLnUIjVNtDq6R84SGjWBtnQvxsCjky+CNsDtPBH9vcpHcLCHkpsB71ZwVc
MkPMd69rDt+d03dG8mEbAnLE0q5Ng13a5FgLipbNanBY15JLsq2c8ZQ4RVvYvemm
x9NLmDL2ZTBnGM8C2+TUy3i0I/W44HJ4K1YJbZKeRKAqUVjL1V1JIKTfJTdRcCgL
rgrk0BK1siuBl3LWtp47Ke5RQfJxtxvNMpBkGxE48vslZXiYjYxk2GEptETZ8Bzo
O2i6FSlaHmihQHHCd27gky3PuU3TJaghqWKvq+ho5CkbE/3N3HAxzwP2/DL7A0kF
hll8W8RHnCqVYUeW9Hp4rAlZMyR9lm5n60hlCt11k7R4uJ7m51YSaTGqQwsOiqYq
c28xcf0U/FL5jIEM3AwR+Ogb1s4yqMiEJOP9bDP1Kh/oTVLailHyGGe/Qex9UxMT
CErDamROJDfnowYvnomdeMgsZ1MIUg/r8vXS2xmGzAKR0KMTRnFTe+Jki/CLUYHs
qVPZHUDsxP0cDIGcLTCaq+S2qNI/iofBoLjtbtGdPYCy3D/q03PlQiPLdwkBP8KE
WTKzm0338vmTZeQpyDMrHLBYoanLdFoteEXItyJMR3jY183tE0JooYVYVEvPtahM
i2G/WA56HIfkQTXwvkv+4bXBPeg7uqIWTCR/l3HhabIaLZ0pBRctAm8rthd+kgF7
gB2i4qO+rl8t/bLbFDWSPlGj8pH5PG6wWBnzXJydwPQ48/YNUZ+RcmOuOmtPiDtL
pdA1awkzwwWxBV8vcxQNc7sqZLE7A+J1ZkfuUMzIKEEec1QPijmaqjQUMgmXYwRc
8cI/hXWR3xoYfavFJopZOcUy61+QlmeTMA6vj941TmigyvY8s6LCQdJzUrKvTZvA
bEYf7wgDBqLINQT/afy/Py2uDH8aA+ybX46XeGem1gEN4fLe+wpNqrJ+oFVCcQyR
539CwPOYd8VW4FS/9xsLxRnfDAeYVYM/tzUB+qENZfyRTfbNiDjRdlet9k9XKPlo
3RQ7wWwuk4Ap9fgQvzWk8Un2mY4qln81S5KijuA3ksbT3f2PMBTLszDRafoq5GpG
nvcdjuSdu1McMInWyXPxpGVXJeRXcE+ax/7BS1tOGuOBmvBOFjaG23kWYKM3BArw
OKylntJl9lllOgkKPn3aVI2o7+ToyQnyUqL4TWmYOZxbz1OanlEhFq14vVO9Lmn4
zRYW6zDZ6iafnxKUlQsin4qwN9hPb2b2tr1vox+NFlEofDIh3PdrpbxaEvsT4W44
pAy1pok/ZOCX5+gn4o+X0G8DT9KboL6yPTMqDIjv/xb0yxtmwEOZ+c3aOZPjbpbV
WVwJJOwV06ljdUd8Wo4JbesIJxfj5GSMUK+TGUxmnV1vN+nMulTxs8YwkLn0z+UB
g1xhcXs/T8GTNGeE7icXXV059mDhxsw497rg47PO28+Yqt4lua+MUMux+Dfh8rQ1
oV7PL43KPCwVqq9lLfCqlvoyfoFX1tO45iqi62K3zYu+3+c5vB9WrqRgoEo8fuJi
NDgKccXg4qFgLukRjrYvjxvuAkReLlvmJ9hJtnUkYtd3N7ZBhJeBzcI4GJ88Zbn3
rmuHT7+VQTxNh4outVrHAaxvGzNVp718g7bklMrZuF3nGqwNyzdGYXZg0QIyWaA2
vsiqj+pr39TQj2SqU9cjQ9cTrVNmaUxyjX4Ch5dFkSEo7Hy2aFq1BrKPB9Epn/6l
s762tsYRv5th9HTf/J/iYve2+dTIMWJrZlU5Y7qPojkMRyrq6VXFaAD/EcEgzpSr
DFDC5LfHAdJ+F9d413Hg/YNJsQtWH9HPmsYm7PLZbUpsKl3DVOj3AYIgx/4C9Aqb
hJqYYz3zeB7fkfnShK7wsj+HjOjBo9fp3+WvNs4wJKlRq03eUKi0pxVEx9nPDWyO
4rrCLmu2/ZnEyW5UW0hCHZshy79bx3uYhZDZ4b8LfChjeHVOeecP88RnsnUIYyk2
b4wlPmFwKlts6NBkBpKRp8z8967Fcpi4QXBCZ5ZqXkeUPft9eFLwlrvsu+eZZhqT
WHe3519Ld9F/DATXax9cGbiCuCbKa5py1CsQJrB/nXlBi/QQRvy67JlWAQ1qCDHX
Ccul3fDSBrdbAD6KMluB4OIxfoOQZeTkG36RQ/AU1ac+c/gb81w2ncRx3BNcs+eF
G4YJ9q+6LZEWOPLVfjoCwkhN4+wK7Tde5XgOIOibAzCIpboxmmGsLPYL6Q+dgcyE
dQ4MvoDt1AX2pZXCCdS3T0XGQNNRVi29UqL0x8LVykUj/ZHlIr/9kfo/tIRO8Jbx
MoFObVbuj3r5kRiFYjT74WEg2hfQ15Cru2hDcW0XLsvxqQ9KQ4jnjJSnEtrcvGXi
PhxyIGJ19hxvvokRQE/uYMxGDujtB/IucBUvRB23CQLOZYHry5DSqj396//AZICe
lFlSii6JdlCei9rgXWUXaGBQLbcjYIpmitlVUMDY/xvHPKTb/WsSM0ytUPQTkLER
O5AF1OZaesH1Xms2BXoOYYoQ+WXqIgcfP9SQQeiaWFyX7kpgKdni6XuKx51oJ0Lz
Jl5RN2NgtjZgbSaL8t+JEk+DDvUADOv3PEDdNWpnukfkpl4WzQ0DK9wahVs+/HOx
J+X+y+GtYGmeEpm1WVTDqjldVtJbQ9vLJrJj56dZdlKD6pMTojEgBlIvIEvkTm4G
G2oNmnTXn8iShw7Vp5uGop09P72nQoSqJbsbm6fXWJ9h/nxhbeSqrsQmodo+ij3U
VhojptTy32BlHiJJOuuHWZXAM48zlJhJDgcpp3zhqcK+yCr+KwWALFx+qOVEaUGP
GHsX4UG8kayonVf8Z0LNOGmPkRhv2ofoKDCUtnM9kA4ZMJ0h+q2QzZtt8i4kUpK4
8+Rc8rEDRZbiY/cP8FyrRNFYxjkSr3r0s1piR11KDm7swI0AvPOSU9mD8lEKGJ2u
ly6YnEhaZ/oV7qnjQED+/JcDjTS3YhCSU/VpY6961Gk+qJAcjrOifBPkBkKJjFAM
PYyc12wGTkRsDauStrOV76lylUicEbgymzf20GwC3GXa4qR11RK7tvT/D6Pbxnzs
xGYPNPBCOSMj/dldYbMSkEO6XFsPpzqHckkxHcl1OKpJUMsNh97wPx8f2fAByQ5v
CsEF48f2nZfEvkhDhdXaoDB2azQ+L5ioNuqehheHZLdjutbKv0iXx86x/2AB4nyj
Resj7VRk5RnaXqbU+RMnRJ1pDIxzEhrpyOkZV4UTZpEv4JvKWycEcgOYGREqA42k
BLaS2FiR19Wkg/Os+t4im4/Algwkt/PG3oJ76ZErIjI2eI5BcS7BRwFfGxmhD+iY
9LLJMpPGp9y3rhsRZ3a518Wjh0XwkNAMyDwfj10vgJF9lEph9RpE+XwMip9Q0AQo
EzIoXV+AJXjQvrHlJHQPpmiXGszr6Ugb2/Kp3B8AKXPxWVfQ0YEYDOtu6377RvyR
2l+2Q7YFDKV0efqd4KQjpDgInXrY2pPat8pY/tkEzMF6juZLYOvGK/67f0cP2OBZ
wbyzXr4sP+9neesbAOPnU0Q8pupwQP6jss9tnM+XsHilyHfNPuLkBXik/t4hunJL
cy2548WXlpCSwXBO8X9aU55iqxkV6eR5J1LuYda5VfIGu90tcab/hj7n2bm8Hy65
GRqnBVIolWGsc1zrj3P2lpMgvj+93+Axup6502XLzBIjkXKeoqrSR/r4s2BfHeNW
BbgraAd+wK8BGCUwA5sXwx3/zhpzdMWLIXCIhn2Yp4TME6p6LVnUv2a9bKTTDPip
EakGQAQoPJz1AKRh7KUZ+aZiYgxxwp7u9atYuDc0NPBld80+lK7BWHb338Jh5b4Z
9PLO+m48THcdVDPTJoy8x/PeCHSaWb5Wl+O9WoacJ4IVhfKl57wt6PX0lXZxVR2o
LVuweP65cUwsxoEO+e2YNlYPcLPDNDHefD6eFqqTO09Qq2jmr1oSziUHQ6vECkQF
N1KtcfgW+UzVT1NepAwJ2pCKKdTakUmhz74+Il1EK3KQKeGqfFiqcDXz0VoqYlNe
+GubgJS+Fb3y4jmUbctJv1SrXHgyOAgchTjJ9Mlr6nxnICnD0vb3tC6wcQgx9+NK
trgPycwsqBMi+eDzcNTtkhzxVkX1s9yvv/dAjrq3GCE4L/Mt6OK7gRFktkD6GQ/9
koBe+R0GqntrCkROxM96L4wpSh+v0StddnQooFD82HyKAmHcw6CLAT1/73umtPt9
Th9qV0Pl9DWJwBbjK6n1dq/5/ejxhoiVSatC61D1ICvEYS4uJwdXwwdr9iQIVI6m
qlT7MMJbO9n03xJ5lNSLyXjn1Fqzp+vxgJ/UBWEq5UjwmEV28M+0Ft6O6ssRz1mx
zZAzFnbYcj4/kPlNanMzNeZ67KY3huaKeknBr4xSQuRmXvgb1XpVGNjG9RpefkxG
zkgKGY4MDkv1XVDEICIsoFGGsHCJFij30ewmTx6IhNOoNnY418ArnFxVRvPMY/T3
yPdEQS+w+jsm3E+GGaaC7e9NRPq1czMcHM524+ROvvGP+X61NVEfhETzUGzU5W3c
ItjnWBEPrvvy5Ky/VD1ozaF//w+vDK90CFJD+Ar4QxJSUagMMSFf9Z7O9qdVlCWx
eDZZ6Xk8qL4tbrsGeib9JNTFuIsQYK1Yif7Pr9vh9wzImgpxCNmAu2Q+uD3BLfCK
1xchYKRo6grRUgSgMgNSXlk/jwkDvtBi/nLG/3D4WXhdggUyqo+SzhbWMAJCx7cM
BhXZkyAnVggMNekGI4AxEanJLXV4Q5uAPkow/R8uxmuaRiQ8dZ++R0BnBX7QN3tm
hSy1+wAtO4K/V//fNPkYKQLPoRphiNU/+TiwuLw8ZIQaQOFHaqQ2tVgKdjlU3mPP
4wYemwMcd/nX9YdW/zlQFWJjH9pLVSxb0UIKexPUEvHtugU1bKiTr6ST5YRjghDj
9IHlklds+p+VnfXX11Zk6yG2qeGVLI7ygzz2mshnSFvlfyD7j5wtUaCyV3ygLLxP
NApl3xczAReP8CPnMwkYBDqmFo1cL4YrV/FFeQJm4cwZ20C5GEM4ZCD6Omr755y+
b6j476fwwN876v5MScy/hiw/7TfrHZ/5WJUa5u/0ueqnAAyWE8HFkRFKJZlgo178
W3qxQSfKH/dbnuv/P5HHFu6ab1++6DJBoVnHGzoHiUwz/CX4orFHtHb5YvV+pva/
cVrrL5Zyx/KU0hErZSECHA29Csx6KahKYYxghEoUnPCpZ1rUKKPLE+ujqZpYEHwa
2QozPaeSBvM5Kh9pNiaNYwhTFMY2uyLohv17wX4MST+Erq2A9a0rQ8+kMUjavzs+
bZlCYONcXNfwUgwpvqAHaoK4//GJiVk0u5kBUuP1rYtwNuaFeaqpbPHuVXCEB+E5
v6EksOPU9tFWG5QYzWcFkWx155QApQwJfjHXT+W/B18302Z+tuSna9JNMs8TAOwc
b/xJ+GUkAWEuVw5g3NnoDywVjn7X1N7tzZtTsiHY1UlvuE5lgdfqCkfdsn8JGtTs
AcpPQhe0lLaiWGbnKqiLCnBorNs/UgIAtBem5g9lVqa3xstq/Ho8c9HiswbnJsCT
hCdGt9SKtWhPwIxE1XYEJgWzW2NLwsaF/Nlof9r9qbILSkY2tpMjlVPz6BhFCSGn
JUd6sTXX3+T+LTUNqdwCsfXLxD0TNO93R6vkpHxL27bx0uUShxNs8Gg8B0F8Kv5M
pZuuZf+uDTVpYDW/vAQ3XRCWSd4282x1YlN66X6CfCQY6PyFv37N6qcUrmRgIZHE
/dRh3g7/b+5LRGVQedN54Rco6ACgltpRL7XmZv0K1SmPfRlufNP2MH2qCupVqbdM
M+YO+aeOj0uPPIWd9RqgzbFQ4vC7iSj/9DcR5D2Nt3Bz4GXhXm/2mnBb6jV/+2j/
LeaWOfaE47Qut4pQnsjgCQ5CTxx7Wt2i2a75g3mP6TysCoTZZph7+xSx252MLiLl
hD6Pv9rJK3ArWGifvOGZuvnpHvZZxo2brU4rMLdRXRknrsgNOPMXBBJuUVh2i2n0
j69X4z3zAUsrl6KokcU06T2F8ES6Wo4iRrLpkrma3PUiyOxlDn+lOV9blNPA5SKO
RDkK2h76yRy9Xu9WLmnHYdEXrwPlEMWSdOW1k1VmFSkMXUP8b8uq1rMZwHbbR0ZO
M0h0gpWSD7sfr7L59OpXipWTlttz0KvroPrWgsOhbmeq7v1Mu6ypnjyOBgovZJpe
tqRz3X6EqWOHgQjeAiWVv8aoem2n0LYYkaX0OWP1r4gVJSah5B1S9VDXduYEKC4b
IYrzSgOXVeXYOxoJzgo4SktMoYFw65rU+MPYzW7VCZ8JwPqwAnySwbwJh8UBipO1
P60jVlXZQVnXvxQ1jEXoyVFlpND8ggMhsjjl7Tetysqy6X6BTGaJXRFgStoL5mld
JgtPx6NlbPVZj/SFMjQwG57juOQxrDUoLxZGc2WruEXhO2Aub86qK5q6OqQ7fXO9
XsglvWCMsmEtPYXcMllEv8EHOOJb0JDbHVx+5BxG7ZRoyJM2q882FGT09Q0G5Evy
R3L8Gsqodh8eNPKRynvDhNXob/nj478dJ2D+4mEqjsAQTSjFZaCORUDHDtMpNp/G
hCyAZh5aDRk9EQ2A6j2FgCpN4SYJIQXItjQ8dpK8gdiPs9ksuMieA6k5NhYTJWRy
2KtZxRfAh+lxcIjDYtG5d68PfkFpoGDvSEvFx3i12b/6Crp8hDTIcUpefnVJtprJ
BFZ/3L19iGGnOgGjkH1AyU4gQ50A7UVq+tXKtImeVWC0iCwYgKiUhgMuS/22oFqD
uFvfOSgaIKUpLdPbWL3PMzv+DJl4A+4crRTY2A/UG6uatd70LfK1FvPZwU50JAEo
uD4oRuw0eWSlGywgV/FT57qcUty6DZzL+zCZGalMRFc+EGGruEWGFfZuQ/IGXhUS
1VrwC08M3fgEEadrbLemWlK7sA1EGoYANNvJYfRHg6Lo1VndhtKJgJ5xJTcZpg8i
hP5WH0WaX5Yjttur7tYyan26fwHkd3PFenvRMAsp9bohKuGHsLLb3jMPbOnp2R5E
aYJigD9MD/cuy1pecjVhOSxp1zX8hwJqMNtfLZdicx+2n39tPAvws7GU+6sdmNFp
ZapqXDnjYOMfvxfw79mgSruKRj3LQ86c6zVLaywzGa+qJwBHLlzfFuZH/nl5fhGJ
aFS9kw6JcDneKnybvLVD0pUDa5zlvG6D1B9t3DSkib+p1uUpZkznIJRsZGV+mvm9
8LqNTTgWbhWoLtpZQOr8RmkPZaM3fRLVzs0w9HYUfLhD0eNELW4rOHL02NTSOrJK
xk9pg4HMMl+nijOKXTNMVPjVf1ac4sDqWTE1KwzOc9GQy0fA3WZhGZ97hGePWwIe
4p7ElENVXnU9+J79fPd+r7t3RyIu+gRdy34QPc8C4qS/WPpgRLMRXfeihwQK/bqR
EUqBZmqo/BQOia8Vwalx8fNvT16aFEhAuRup+1FHzC0G2Qu0OYdb6GOUZZD/yamy
KaqYwtV6WFzx1BBzNYbZCgWf6c5ikz1e7mLZt+p/vw8oUro2S9y4+QxI8RQV24gq
LXHVszEVI04uXex+wgnguDqIOERwXTrs8TB+jJpmPWg33GKq5F9KtNvGCyy9QKjW
zpdzoCw0AE3DzcHhnJ/czj2hpBcRQx3w6CVBhr11y+EjcCr2RWw455GOrBhwM4do
2Ziq4VXLBRqQU/0cl9ObCE/AjCeAvleap9l8wqL0iAawieVIwTV8MuMMEqbfvNIl
0AXV0AKbw35+EIgdOgQ1KFyAawc6TkNxXVk4yChHnaPYsQg04T+DPmWN+gVazoY8
tNqgiu3wVvDdkaDXfNJVRF8xbhAn8S7wybYgzXmLpkR1n3R2CJb4vbNl5NjRYl8J
j1lEw0PatWwIzQYAHZUM+i2EPZCZRC7dXCphCbhRwZ1CTmXlV25duYUKN//dGXrN
A3881CdxnCSN5sBb8g17c/4xpKoT4xSXaW/iphU+xXvKvM60o31R37rjO3g3P64m
BVZeqeCH0PbNCmio3sotOgOM+kruTBpm5wwFPq8801huzrEV52ovL37h6bu7PmCg
GiTWALCHGg58ypqG5QgqWeiZwmoGLRL83hb0SfVAU4hPvT8wol65uJOw+GGcGMSg
HikJJiHT9u6Diiniqsof7OiSYIy8Zro3OmnItF/9CBvL6V3Ix1hrdWSUJXJbak5s
Evkkw4TJNVN02RVo2DYAfb9kGepyHSslBd2uSHcZf6snG5RKFluO5KujNyEQbaHx
4d53I3p/p1ITC+YmzcqVUAdj/UcEdygfUY/SIq+9P5yE+A8WxqXkB98n1sz2//C/
8IiI0nwshIz9S/+Ml7XW93Q6TcsuYMBNBIT134Vfs/qWUypmWQnIwFjvciLq+Mpz
ENBxw5yKf+Pf5WdgbqPlqU8IhMbC5L4pIvd16DO3iYZ1AKX0wvJq5gc19cT/wSIA
ktwCnSRE5XKUVnscrQRnbnAgOO7aHspQK2KrOd+yR7x3OBBHlq/F7u9JpPT05EMM
qLbi3dCiULSqpQyakU52AwkHuqjghRvrDZNvyGKUqwPI/imGlvfknhw5795QrMqv
Lwj4FNu7e/0QENsGix35jIXjij5S+jSXsQamnm8AXximYOlYJx+5U3yTs3lXYIK4
aQ2TkTjUlHuGnNI4AbjrFInlkhlH82/6O1XKGRJugCSSL1rKq8Yofo961Lww1mxk
cVI6RIv2XXeP9Hm/uuAORYazsZ2Gqy6XLvB5mXExkZdMGjbtH7Wh3gisEfjmY6ph
tWaAiklrxkawnY/8WVP1OY1jO3GLVFkw2pFf318exYdiHKxU2uQAXqEo6p3SZ7Wx
+Oie2NCHbiIRml9kEofky6kWE/meNnt7Rry/rdHCDR6ipXcI9Xm7fSCRUOPURt+r
2A6dNWpK90On4ZBL2/Va1nQQIVxTBghqdA3Qkg9x0S5EOgmdvDx6VwiHzql1DQg8
39lF46jJNFGsfCmmnFZnmPkxbpE2VDi9ZtJH+cD6xQsXJkxfFiKuKFUknmvgQ0kT
2oWB4mJDSFPBdr9AuYWuq+6+mAOEXt/qx/AOaDof6QQ3je2zT/Nfj2wtbN6tVJ1f
RdwGMLF/Zd0tGUlBw6fJZsYQq9xgvBj4zMbWgiXbuclim1TXvUKhpoTjvw4o4ieT
tzczAyVb7cgun25QjYbn9gnIVZUWFNMdpJc8lOeDVUWKcgGmKa7mLjihxtmVZ5RL
AZhk+MLEFhI0aAIEQUpAZBAzWtkxKG7fCFlPeadl1f+6hTqvD1yFiCd7rUHdEdtY
Nkj0M5g6rxzaHzh5ZR42mJq+A8dcvgsHvaACf9fv5wjLfE3hRMjApX4jDKl2DkjG
tIxZu7iifEP3IpO1fVbQ6gmco2Li06XoYXu1BcJULRgyyUJVYzs0X5alsTvstalG
cZ+yEd5blE5P09K8Kspe8uNLdv60ecOnDBGBep/OiZ+PS9DoNfQJP8XoNCV71H3A
s1nbU9YnnPVa39a4o+7W88bzSZNPdzhyS7jYtgFrM69nL+0xyFOoPzoa4j41RTis
dnQVbBFzWzCn0ITdovJbBnMz6FxkDreb69CD9RgLiXRYiKaQlfUzfcux38xVcIU9
HvISFACR1CmhQ87YbtLLbqMY9Fk2BjY+18hWizr3U6pRhq0xq4XlJN/HR5vyb5S5
IzWG41kVdAINxPT3pgRiKXZ72WtxYsbGBEHhysMYjZtl+cXDl3AX7drDkvxxZwmd
UfA2+elB4W5DmNCUKeF42Xw8vQe/vhQRwdoJ9BhMtGRaKqEjcDR2Z7mkWP53wNPf
wUjMEeWK/ocki+zobYXteD41ENxnJ4lg/HNhS2WjSupBFBCSazTH4rg/Qf0H0L21
2iGWpr3oqnz4baWsr/gaoct0ZBALmuTYKMLnxwDscztNIk5D1lzpL7nGBjGSexHE
KagG8bgS5MGh3Ko5bJkZz3dMyqOSrb+cnWHVhmgtegDRPE4wawn4+hW2nKbF4IUi
j9VTSLhao9cug+Ym4GSt2FJbLpXtpnIvIGWjPadf57i7KUruRimX98ru2ZSB0pwz
xY0r4LQue91Hr0PoeKvomkW3LtxNvYq59v69ayU7P13Zp04PwYBvlig3ijaJ0ihk
BYB3e1gI+Gj93ULH7cWOdrQAa0Y8ssrG/kHvwCcsxucgcYnJm5fMNm0zmKYDzh23
eshTsCiaYIwTe37MAh8c+1FrwIXY0HVmP+BQUSBCs1JVWXOXy6vLRCqa5US1vLuv
iowcq2bCXoF3f23sKoXvgtOEeLBy6Ia1BnO/pKJGz63PVeXjjDZALLZZw8VGouKJ
mcHpPJsmhgLzhsw9CMouJ9vUttqB+frXRU8OTz6+M18o2V7sBJM1j4A7tb3d/5Wv
4MXSK1vmrNP85Wp3Hpyg7o14LMGu8+q4DydjDdpl8uwvgT/cayM+xONZrYVLQahZ
JUXmwK5P9DPTks3446KMsbGNSpxaYMA5UZAyS9qWU75AwoNw+lCM+P/Y79ljZrVe
dHL+r8i726kZwCEvfAxnltPoDI6rxOP3DTuKGa0UaOswH/gbbntZYagUvcPYoRwk
+Jd3iqEqoWkpdTmYfICoRFyvAXLs1GTJb7ahwSffh+v2/fNwWTaA3ATxPn3TW4PF
b2qxF4I98gmN7Mm+sHLfLXPDFrL5fklbOMBiOJplKA0H0rkR++ZEfMlqsdJbbzvN
7HA/oBKTxBziarjWcVm2Wlyl6v+ZH1OJZ+AAHnMxJxnJXsPExBEXMioHfAjKHyG1
GUIPDpRzUHytekMW5LM8Bbt62f8E9QIKRrqyU2woMDgIH0EgD7dbT48/5uEacN/y
HIlML3Vh7BWzWY+r4DhVi/M7PGohAk+24BIPlb6MX3FisPafskpMWTfNqoeC0cez
Msa90rAV62bhTU85xekt2KKtiwk+d75e7wzFPl5mnD0VNLeGzC4uIchc6v5pGkUl
G1Mhoc35D7Hk/7vsEDTR/v8GB5VXVEMxGZD5oChpkISNfTDyGkIRM2Lbsgh8Xkgo
KqRSK5c6cfigMh00ckXCumJrzhqPhOfeywi+0vqGjc7TOw1KWDQdHqdqKmGpaEhs
bpI+LWRUEGMi51zpTgOqzOxsdVLjqmMEozS781EHTymDh9V37EFw2k6dtVAQBCxu
PV1NKNKyXNcfLNb5BnRV8oof9qvvTT/ChLX44TgGjWhO8KnC1gVMaMDTAFqWt6pg
8XwXGqWTI8DI1Hr+V53kGeeeR36QkiupkO7lpXp3esjHNp3e0+4uW5UBeGoyxXEg
XwM2xZjKOhcHoFAY9I+UQvyazBnwHVNNH6xeMRo4mIXIK8Yb01r73tc7Hhdgm0hB
4yrHb5OCcqvPaSWPGwiEl86MfiBMJKtJURrdKRebqJDaPg/FbnojcFT0voce8eu2
MpjEm5m0gWPL7sws0DPrYaKJh8lx9IvTYJrVv7Wehxsh0xurk0iQUKGIKZ/9yzfo
ohNt//hno44mlwInSYHG5WVanXi/WtpN7keJ/oosyweEzdSzesaNt+uMom5nJ5XS
4eLdFOSYIk8/zgDjUJYHXp0RbO7yS5HnmsqpynWUbYVwPNjufZHb9wuvUlxUuXB8
C5yCXY1yEzivwQcX8icR/8jurZjvL96hL0nI7Y6PTOhhju3u7jGb2It1k/aXN2b+
6mh6s+G0Rc4egG0FQBrHHy1Asr591D9QBBOTpT1nZ+HKTwjMKA7JltHbtBh31d6L
g9DLdf+2te0eCQZFe3MRynkh7aIT0vtYoXpxhn9ouhLiR3BaWXNlN3OmlJiTOjaI
cSDW2JISRJSa1J16XZcAvH6gxXvP7bFwm3AnELwVUzWagfHUgBKWV5MZ0TRR6Wkj
XB1SI4x0irxoEe2irdv9LO0OpG/JVTE/+MQGDHpi1eRjsE3mIXvh90A/+5iG7y2K
5b5YYFk+FcNcnI/w3+3WWO56yWcNrNP9tyKWsiuYEFSYNA5kKVJl9INeOX6zz2Te
Ck1Q5AYN26+E59yR2gb/xGlIjcZW3iALVGjcLBqKiGad7KGaY/aAgzVIPdHEwMhp
rn6B7SE9E9+5+gzt0ZKD0bIRRDauHWgdzmMmbIUlIV7PC3zBCX6AJ1t5EWCnI9g5
dr6gZBJxwO5Qb+4l0CyY2iBNYwElVNJ95Nn/ekgYpR84Ucp7RtClkYcmgNwatvMa
8nNNv9FaG9covKFDuJLWfdpa30q77VVkITEmrkJDC8fmlrUV0qeRdQ2fv7ScHFzX
FL25ncMm3wowenW6bX4gXvSz3fhA62AhwWtAIW6JMgqNByOPAsBTbindtmzVwag5
0COytoH70Onfemknjn7m1WRLN9xVbKrT244AknOxrdTwahrSTasicldGTvJQ0ApQ
3IbKJiUvey68bMJeq1olFwR1NDrElB+MiP5oGLNFCc01Q8TlHwtlZWuD6VatTkX2
xAUB2SY6VI5SI0S7kAKA8/8VihYlt5Km0Fu8XAKMs6EK3bzsnl108GDyTJymv+Ff
cACQky18BcXfdE2KSEcwS6v4jBz0iJRcrArmKDd/3o2Yh8BpcPpYuE4oKB80hYTX
gYJ0EBW4+CCmKEsD/s1Gr1k4anu8vB8NcFAHXVZEC5+O/ofAe4ahHYogfX3Bs/Ch
7ppueEmGnjc42Dsb5nZgl9hhDX2WImTiXTQ5z93oahJWpZMKYb8KQToqkysD3k89
OKEwNOLYqUHqmqeZ3PBukdnuKKPLlk3ZSIc0ap8cRMPHE1W7+lJNnw5DfdNSeWnq
q0k2I6C7tmsonyCQ5gV6JmSeFtHSZL0Qd4q21TUprHxw1n8rMlI3YFMM4VSuxAAd
vkB0jtoziIgMethr3TDHcLBt6PpaoaVz0sIK7lCJ8OqE6tZp1oj+blfahyrP+/7s
kcFkxvntAZZirW1qatwju2b26FtMoN793XUpgDR7wKob7zNV+Tms5SAfUl22yrfH
HhxqTK5/a9QySJsP+QHsirig95GAFGsbAnlnztIF5fYCWilLpuPmX2U4q2wuKotp
4BPJr8kxtCsuNwLh6mBWKNjSECfrjXY69kT8g9QJ2ZWRJJxpEw2pAhWex4WsO9IS
yUdNcGM7G+6i6a4mJZNeyet30Ubw4qfSEpxc+SoTPWDu6BLuyg7tUx2n2dGoiWwl
uvp8S7rutRzKA4M/lNx3dWx4zBBB4DtTmA1oOHWF5gTM54umt+fBWuxx33VB9jQh
7/09U+kh0T/hgEv2WLiIYjhUDW8R8PQ40GvD0ranSugJCf/+Ow+Dq7jaPo0vVo0Q
j4XFNBadyN0R51Nr6b3pR5AuY9WeQj0pqFCed80+wYIs5txBI6VD7fqrcZYwPLq4
z2Rv0SDpcAlznZJ0XkIWH52XcXSEmK3Vnl+LAdILgbAPkT+u/ndoMC97yCyxRinp
PV3qbfdHGT5bbWokJ1PhoNDk+7A6KJ9LcGz5urmyY+vxU2VMTazn5lB/c/ZXpY30
paR0Oba6IKO+nVXfCC81kaUa+SvanP85GRxejK70Z3WcaMnaPPerw3bxfJpX1Yke
O4cL455LZu0Tb5PLKx3pkMj7SS2rp/RCG/qf4rdivyqr39V/K1dXF+8PHtyKZybu
zTI1q/NHmuDK4o2dCpn6ni0SgaDEyN3hJHDCQC+cUBhDtlDSXIEa96RnQdY2REn0
1Atmhl1YTiA9wPzaMN/CkdpNUa+P/pNM97AKMXjpsS+AVrriNFqor0G+m53MqrRi
I+UzSZg5DHdXBOXMsZJGDic8zNRaLnSDmbs4jAA4QqJRQcv7mMiEzedW0AXu0Mj1
B9y0AFgSrIYb9SRwraCLLRZxBQoKsAPGoFb8qxnH1CWkB1lVPSN9UEx21JBLtEKG
HN2QSd+hAJIXzbokAIiLMfF1ihICb4kejxQ2WFrjju7EeS3pKQ+sAzNHfaAnhv+2
jMF+76Gsr/AETqnCUG/DSMWZDvbKvZojTo7LpgJI3SyDXUE80aoHFKy05cWVGMjM
iwWSt8cZt7Qh5K6qAmY8GLQewTl+9UJKSTaGKe2nYrEjpc9r1EpknyZeUsY5+fcW
6e7xcHhQW0o1ltl8l+ttdhPKzPeqjj+GEbxmZefL7V0/osdgoaG5+VHjUmPjcRPy
uohuWw3xjBHuqWPqJmw7bzMBfq1UG4LuyitLpKUudW8p2zXqv9/POqUReaYiLgIX
qob9R/HUBBSmLveRp5jucq9qOktunfSC+kgnN/PFWsruxl6a1wSSWNSz44OWxSKW
vna8Dgbg6Vf79lbbAFXD8rqPzSbHR1KRhSu1QEERrtej9b447iQms9Oy5eXWinVV
qqSWLzMY1/Yfr9vtX6wf6ozfnBZvFLZOHcP3QxwQfW6J4hqBJtRfLzeE3CVLlQZQ
G8k3Yf3a+uxoL0ZzN2YlnHVeNNhkDGcxbz/LAilavOC82ngWsDZoyLgnVx4E/2iK
KUfIeZu0Ii6NagOipvwhCXtlRbLIe38hmr3TEuPk0gUcuyUmy8cgk0I0JoSpmyMm
SOB8myAR3SG+Y9K+ADCUgd30PWJC+a9aF5UCcmlEBlTROjlFCSzUJJ75v20a2T6k
ihHSH29vaTIPWCIZ9sb+ix9HWEEXkKFEZJOylrfByc7OSeqN21FJQYGhMIZnfnlt
kZOJ9I5vsKSF6554C1Pi8ZYnjtOB5rNZbOHcDFGg3socLy9MaGqTjIJCF2p6o6nl
Vz75RQ4c4CFw24tamXumPozenISrknb36MoFluMztvDj9VD6EAd4+hTj1Vge2kBp
13hUYIWj3pM6uIMnexh/w2MWL7qg/WbVAEfmTojsRhW8PaOA4alEgey2dOwLoyUs
OIupQGQL+wKiRjTU9GbEsbj7y8OlOZBgeTOH3ltNRwx42Ze7sCT8c5vbruHHXflA
UropVQEhDfbvrcSxmU6/zFC7vwLN5vhnvAFVZKD7JTVrVoHQbPyDK9alD8j4N13j
AknOjqhs7D6Je6LNB6eYZ+F/rNbRUsTT/P4zXnS+csnHfo4OyA3/1FhjLw74UMqI
ZG+HGmUaTYcd/B851EROgPycJCy/qoaQm1SzwEwfPn1vRzAPdstfVT6cJNuVvL2+
yyBxzBdhy6RKBLinqfAZWkPKS7srih4wDtY6nbZbucyO3DvkoZf0Y6EfiRkOqdBD
Oa1BfXVgBaGMp8oQPPpw7PtSzsMTt78dZd5spCDLlESjBVefRBIGXPvEHFC4BsDn
SPilXOED2wqD+EfohE0oCaU0O9Bnqwl39YqmPLOVKAmDR131FxKggSLK8QB69J1z
KaNehAnB6HX1SK6mQAqomyjOUUPsOGkKgoxNo7jIgkhzKFN627jrDj5hmfhEdE/K
9U8jd8T8fwz/+q/hkc0/L+MOXGW0L7c3H+IsXm2GNZnVA8vTSCmJNqEFqiQD9TJ0
oNDj73Zen3mCrbWsths2wRpjWax2eLVr1iA4zz790AJayGVdGFNSSpZq8J959+MN
ef516RrbK+yZ4YRhhS9KB9WFKVvHrtFJS4goFxMVEnRZzVy4KYmtiVCr0Oy2P2iA
Ibe5NHyiv1TFnB1KIHEgek4lYLRi5aTUpWBA2Ug2NBZdcNdWRxXNNjzjZq2gAUMt
/hqQufBu+dxJDzZ6poNTrOtQfIyoEGDcGfJ7O8y4Cjp5ifhCj7s1iaq18RkF5WEs
qA3k1pDJGDsfpUNYGvqLCKFk77CJsWsTpEzMsl0n5LVCG7qd+AArkeCmD5XySmso
ALK2muduV6KQt7rGmYOpRb+Lsx3KHaEgXNsFwi3I3whQmUQNu5wQJB64m9v3c6ll
Q0h1alTDE97RZtZZmulquJFNDV1JSZgvdUq91PIPQrO/EvevXNeLRe6dI+bk40eu
sKdQLjJWhFFs6ZNpn19qdKEE8AJQpBIxi0hNJxFR4bhuMWZP87tKg6QH/VpvVMr0
ET5Mr7ggkNoJwb0O6MvRc2UXyRICxoZ4+MHQ9q8m2AKodp8jXLqKrQbpDVtbG442
UMz1doIJo5J1zs1T4Eb3N23919/SX9yNYALVNzabvnBxuKusCVXx3stAS1ASYPEd
IbPrSV3AXiCnZqcYfpFkE/+nc7pqQSJ3nr7bc657D9WwPWis5Mm8OyPUJD7zJQa4
vCwE+eYmk6Ap1kV0Sk7SG1MlFXLPnsKjL0RyF3dRcuz6C7xwvMOX/PLwYsezjAfh
aABSUaS5zPOf6wt1uVdshVWJcgwVhgYhA8syZRHyb8nHZrK2FQxdav1NdkMtgHc6
TzOBfkVK6I9rtgZ6t1q0zyRRRfMKUapTWhh/CWEMrDwSzTv+9j3ZYbTBt1rs31Sn
I6g37x4JbZSGvVpI9f4nIAat4/+J9BPRLXLfeBiqCNwh1y0H/7eZuNi1uJp+0I65
fxwUvBFK/EIdGtflfdBPV1Eon1H6B1AZ6/xtBVgjmqwRLphM5iFORN6wRx2N+vaS
ITtwuA3+ZMkEZ1+GFXVrqNE4va2cRvFAnxXHdQOV5QIUL8ROh90501iGs4WCwcOY
MSEcdjtj5wgUFNsDEXTRYbqmYfVLb6tGx2n1snR0VKx9OZoYV63ot+whiYg46Rpe
boVhrEgR8nw2Wr59GfiGSGC272R2lW673598I6tTfrrqg/8xM96dMLLB1YV7b0JV
shB0NPqxVQcUGTxl3A2b/35OkUdujCXuCU/LepTaIvnjqO61eJTTdjovi16wDrhz
XI3IGBZR+ocnD8z5/ro1DB9r7j6wtuv1kIqxF+VB5GIN4Fcnl8pswesX3lwudnrZ
x+nT7/V/VFz2X/3cVWedcQf/ISi7Ib6UhOpzHxQf3ywBDnCRvx7eF8TXN8T2MI84
p8SLJy5NtLZu71a/kUGHQDTtZ2uefTvnIXF4kuREm1nCXEEfPZbFqw1gKqBkNKza
c+A6JtzFRggiYwfQ0YMJg8b3U9g892SLJeOMjx+BjKKdWYzYpdHwBTMXL9i6ZHIj
FCzVTQ6HXUqMHa4DKK+eVasLQ1EOylKur/8sQ0Bq0yn8pGhomELEIWx0khnRDkn5
6+bcILdHyYvau8MApkIbPD6703H9o1/xsyi75nJGy9ZqvnWeXt/BE26MBmdELMBr
YitHL/5OnTziWh46PbZGa0F67UNB/FHuWBODLklJ2HHxkZWHuiI7Q+immeEuHfOZ
I9b1NQ1f5g29SzBEr9GSThqCm5pwqz74pREQ/exfzZsGUh5UmgCdnoo3b2yIz8o0
Pp20RonPPZ9fTssVQ+VRJnIIUTJC3xbAvcNVhb2Ahlv+YPB+SEV4y3uptiiTek9R
VomCYbbgUZ2H/iO4J0b4gMyouRoW3p3hXzvd3xoIwjI0Vqu9jRly+LTL3b56vw+M
bUN7HDyO8WzMrI5rsc3PiYK7M62E3Z6sShO3/JKCyGBLbcwofoidGP0UL+4v+5LW
pR942AsELRYyI4WNmvA1Zo4hsTeykN0iuZ7KlrFeLE3wAQFD8JnsrGoJ7v2EOsXD
thB92skEn3qSmw+dRJtbGJKRyF2SkBalJNx8b3znAX0mMsG0cFxLGWf0+PUc5t9M
CeJDe7NN28HZBtLXhAHSDyp6KFgFc+LTpk+oZCezaADbO6a8RTJr6z4EjDO+8DgN
yBM2hyuVQBFX4UOdCPqcwC/Dx+XhbQuzXfO/BdsD6ESCDrW+zWjCQG/UGvp09hmP
YHUgKuH5X96HGBgCpjLhIex+YOKOT5vv4yLzk7Bt4YB9kZfhBwWO0FTTvMn+AXpX
JVyZ++kJLkll9JOS0o1AuwG6CHhMIsx7ZO1pmVba9fU3WFvQnDE/YKdtY8L1FPeV
gJVuxU9dHYSrerxdkRytypiywNlNDs+imySXC0SEdjl0lhHVXY7xjYqAPQLCIidC
olv8/T1w7o4t4DKcHBkmF9KQjpmfHoKeDduEpcCX+tEizfRlMM2vVKJleJKRzuky
aCo5VnndxVmz7coqhGo982JNxR1/LMMGqQLObv5Cx4bqQZIsUICODpVTr2v1krDL
uDCe1CWqO5rNALSgKA02Y1AqkkDnkGDzZfAaEHFMoKCROjh0YYs0GgyKpgvwrhgm
IN7DMXZRrw4e03EQi/ivgUwT3tyHZUKZwLYE4j+g5fUMHpx0lh8GEVYysaOxOftx
woX3IqKlN1uWyPbgGKOOEThj7nnl7scrB0APrWJi6qXHWlaDRSpDT4EHLZc6hLEP
JzwYLBOBWmqHFNeqUQJUJlVXU8cjBvekt1sUGB0m/ACVf+rYwi6hEAQrMucTbtZr
3xl0/yXyd1erpPGYjDNDHwtn5oG+VNWLFf9PAvaobHacOJie0lisiMFeueQMM/Zy
nLo1WyVbUWIDGmyxEesi+RVLAuCAffUeF6mw111E8PisYrc5ST8nIhc+bxcLmiBG
4x97R5M2ATUQJVZZyd++odp+i8kPRvnA9+dKhhxgCFnkTx12dmrZ5jiJPRUOWs16
LUJEZb53uIyGTB+ltTAzkRqady+ZWa1Z6lWjrGjTpdVjWwn8tsxyl7DD1Exdsoxn
BBLTZCRatSyI5PzuPbSt9zzZ7Ez9BcCAJV7P7cRDZvm9Rutf3dVy1d7nyHayITbb
kWkKgXte8CUcoUgRfuYinktKUgXZbSrD4lsxXoZ6KETWFeHqsCKDJiGCzgB5m3Ww
PjtRjlQ1pUkMS5CTVqcJkih15kUHIdQgo0LVkmtKwE0Xmyy5SVvvj6gmuYEeuft1
6o3qO07dmwvBK0rZ8RTXHk2cH/fWRLg4RwPF5xdcJ218eMiZqGunjEkITXc9fkMG
rBURL47Po0sWK9+xv1QIo2DwmRBtsZj51rB0UEtB8+ucMzBIH5+quFOgE76EQFVO
glJmi4fekyi4SLQsl6W6NflJ2H9KlUnKjTTaEZ3YyU3wiaDn02C4LELjTw8Ll/9I
4Bjm9ohfGzWRK09tA/I9Rbri8/Y2epq5REEoGzHSbrl1B3xE650RQzbUT8FODnwH
jrwqEbCdQ5l9t9jgpOYrCGaKj9oBF9NqYOa6VFeTLAEcr4PfzPg4sdO18Ffcdlvl
eaBKQNvGjeULyzCVOwsxJE66m8aZJ0nQSaFjOH4osLIsHkAxelcaxpXZuHPHc/VA
Ldfv4Ie3NYvQLuWcnipWxmyrplHwK8QIxVrKniSKJhEtt6sl+dE7kDQpLWf3KanL
Z8coOtr6xBCJRRYo+kt0Btyr3B8nrYoNqh1hrVyZOzqt+PeCz6W9/mKef9eIx/mA
jYop/VhHslStqhr49IHMNyO1zXzfbDt8cFv6oYvXB/hQ3MniaAXHdioz8zd0anx8
xRborM6Q9V9C7aWz/vUkGH5hQJMqM6wlPwU+srJgL2jsImP4C1BzCebGjabDOYX1
1k8YmSU4ozcWq8dqkQb6Nc1cPRYi88p/0o002C9zC8hb6lVHR5XIkIRxwkCQY2Y+
XM/dVu8xSwbKZY8P7XDO4PguVNQzEA2HP9jMuOzETrqFmUOUX0tiOcFumgWWfYHf
h0htBLN2cQu6M3JS8sP22tb16XtZyhLHbEEpRmEZ4qiyNSMMDF9FJ8j6VXj2g/82
TsE1XZ1T3yoBOGYepp0kCIf/cmebkrGV+zU/X4IQj4lN2JRNcA4zM7FWGEYNL4tv
nKa9dI3z80gpmxT6S9PHFXs5Wg0pTadryZZdGyKhES8lt5DGM9gghyl1FddX1g7j
jDnJw4FLn46Dtiju3xhsAhMIfelD4kDtbQZ6zCbz4KLKjdTKPmBuRbKM5ABuVSc9
Z/FwDnkI10V9hKCFUzuPWLhueUV+0mMDace1QPU8sJ4HL1WwG4OFYDBJNYHhln/I
bWT6oM9W4pkFdhPwmsvVvoG9IPTPCaZvZCuBZVKw9zPOKlZGnzvozeWgJAgLAV1p
E9kSGIMAYSTP0ar7T0kK8B/9HrUM9JUQ/v4fA4ixA5ZFR29S8KerICTGah4++1iq
RPyhKNJqF5BUb9sMH3tihl+HzrkI7eQOJsB3VItk+PhEX9XkGCF9B4UzZHm791l1
P5cJZRwH8q/2LBMeCZURZdjwDy+SENn8ZX17mYH8pc5fASdSo0M8gqEIqJ/MY7K8
mB7sy9i7V43TBGSJwNx0UrT/e8aOdOSw3QQLAo9T+3hto37y2jxMaWj5MPY7adDD
pYjNmuFYjZpzzsZeGtyEhNEKt0eEVfuocdnPsQqJGFz44XkKPQTXOIB1xktuYtVI
8eaz4zvsBWihKzjyLxKSj19tg4xL99/5YAM8q6jK675DqlB8m9KV1bRtdbg8PP4A
fNkmrrXtBRcUZBfVQUWSftOxTfhDYMCrwhDei2mqqzLDz2hW1BOse6aMoNTM9qob
BtvyLmycqo1HI3YSJmICHaUd96Cx0jqhOpE4X1+p9LgDHhRwPDBpIwlz6gblzoEZ
Xi2c+vT/CsU+IdoOo0JQkDwKsZaTRgAqBkCNiJUAhvCWMgANWzLStdmAc9/mHGlD
uHNctDknn+hU+jJT85Z59q4mbyKwZMZhv+3uDGAofCxGZiS5akAiAj9YCppPorAc
o5hRPwaP/IpXC5u8QXbephgEYMjYL7bBWgFSSKlv7ANyVhdDNZ3/7z7KM71Co94u
7MdP2K8/vmKedHVezUuEr44qUh1I4FItIdQ3gkaatUDcmKttSmoUhRJmRWaC/9ce
CvmKA3+2AikjEfTEKmRTj5oxBH9SbS+LX2UlbPPffwtRTYfpLeEzqT414nC0YGBw
0jAMsCB1cyHPNE1Hmg13BOYSPOwViyTiSUndreMRT063Bp0zTIh6jeIbkStcqotc
Vt0J+TPLhbaAHMGR3jkKpKEXAynew9SPWov7SUxsWpin5lNiNblP+EoClLMV3ijy
pitRq05r4NDZgIGhxSGvA0o4X/vDTCi7UMq6tu0EZ+gDOmPkmPpwXlPJQaK9mOo4
7w/H6D8MiGJqW8k56rqBvoPVA5Apiu380JrNLGvwSjP1hNBJRR6IqCIgM/1F2WWb
qK6/r55EWprfWp/84ITZr2nvYckAgDGl4/BXQUrshoupmOATPRY6a5vbo98xl0HM
oT2bsYqQYozoLOlHkYco2FAV6aNZULyWnSrPb7PsZR0FIamNgBVnKQ/bt/bNqxzu
xAR/eDVVBqIKudf6Vsum8iNYLRPETPjsgZfQGbcJ+99Ji55IhV8yZMT7ss3M9rlb
7AJRyqAwC3+Tn5mBIcOB3TkjBb/abSHVG1Q/WeWYbjgIWHHyJZmstHXJWGP2gM9B
O57TrRfkoh85AQ6liuqziu8+rkukfRdmSPijo4SNHR14eJRgx3yc+nbSZ5twntJN
CVKyXFncsLiSXASHOUQ5a6x0uuHosVEAm5NHT5Fyi3i3OTc6zHMYO+1Fked93+WB
x2FGtmCmgfFZU4FDbHV1xSdrTi+8GPM02iRz44yOR4CnsZSb1dJrWQL55OKqTcbf
cGuTY1cUT+uQFCjEeN4W1d+DQUK9O9ZclvwZja2Sjaa4CvqoRwKQQzuWjIxNxHia
Svqx7Cafrfd//PyzA2OfCrB+JnVw3GfhV4Q/Z00Bt3rKwcKyf+BKHKz33RQ1cE2k
F/c8rcyB41voOEAXPdFeB2dVARhe6WHF3cCzhBjDRHZEnkUuFKqEZqJSUGEPVWwE
bVMbOMH/aj9F031xn+HrW23eAEl/4GzGVDh6JEOOVUS+LJ8DupCv03r92P0uIQ4r
JErVNOM+o9XonvGBOv6y5oi5recEwADtqvt2DYOgmEkmP8OFJ03uLuIpdv7N5WYb
NejYj9Uj+XAyfWX7U/Ldamfy/BmBGpZ8EgdC/MzpsG3qWAdihChPgHNdJO4jrna4
gDWNvXV7rq0wq3WI6ci7DmROgamS4RjNM/mlhsFNPjk9TN86PAbnzZBAuNTG73gq
TSomMlk9GZJb1PpXNP9+GNptQDSYJAEHDQPQZoyjqFtOV08Edn6aSjbGCt7zTnXP
O6gVJKSuZVpSd6UTOSjDqH/sTAq3FiwgEv/1cOFcANjML3PGv0iyBwMVrulOdy50
nmERhDsBlPv8mMl+Fc5GXArA9uL4dTOlvFokTVQzN2e1Iv4+K9ZUs+fE7/C0VZxA
IhMBoiPdLmuJ2R0IJl9LS+rvruOrfCv80oD+r3MfDz1GVUwuwAmwLn3ed6uRMRwq
y9fLCYF8CDegZCvkUXUQkwGk5QJx2ZGSTOr3+Z7ZJiLalW9POr355YqwfzY8V0yi
FIpm3nFZLd/jOJVSsHPdptTqgmiIPz1xbeCjRPgDGAmqkSW41XAF/FN+UbqrSRqR
fCXeF8wsHrBSmJ3co40bCb2zLOTGtKKfiBhHKb96P+yl63QQNlQ2J8U5ilbEs6qK
3udHv6KFBpsuJGSZfonYo9DzzkYa6vxqzIMrK+OwWEAbkObN0vQvQjoWQ+Oa5zpK
ypdHGs+4MvJZG9C/Eq6JzvfmNZw5oRwCXDFEhcyq2VyPpfp5jkn9z95Co/V6CVD8
Af3qvIWRmtmc4iaNkTJW7djk8lrq+r3Y04gBWWc4nxufhF/GcIeorfRSoQ++q1MW
ooafoXsl9/xAHGGXddGvdN2WOOlctzuoOHw8Rs1CU9odW22SXAMFEBXiBW/oADW8
HG9R9jpcdmMa63MkClAO+kQOauSBTgB8g22m1fgqoHlrtMA4q9YuZV9IIVWzNJRy
ojtuu6i9wlv+hJIx6MIesthGgEW4VSBON8gTpPThMlZDGivkQIVUbeCdjInTvd50
SrzHbCyjCLfUQq7ico8f1IeaUR6iVDcmtrGk/p20xAxAkCAEIiHtcz2gtTh6/Dat
5qv5VLix2+cf9jZ+ZNmEIele2/sVgsVj6bapkz7Etyeq7AL5c5P5cS3519pE/bte
WKteJKiPYeJ7zwygthaFLBosn/1F7qpIqB2w20Ppebp9AKCpopi7VxNqteAoBAoy
wHMNhpuZ82icK0KZAiioeafeQJdZP5343Bb2NroPckgEqH3/yIbn5Nc8VQYSonBn
/hSuKDATBF9xTNBVHNF42gdpykbMBCJ9mW8CskX1YgHhNnYdLBXVFWLdeD7+Wkaj
zTN/ZEOjLFGWkW+WkchHBUPQoGFI2OlVkGhyayqcrjNcERZOyQZmmQRW/aglY9Gf
eRi0Da/549nZ22KS/TrwgdibheUaaWG9YYJePo7e6jdWvoFwWHeoe8TAePNoJukM
dmX4b6j2vRTcIicOHDoJJV2eMb3NIsvGEfCtb9Ujf4bQaxrA7nhL1aCwpIrru8hv
8qiAHGnhaH/uecaXeqU+NKdn2d0WYbWaImBOs9zAFwQCo2GHHhwI26gDqMVGzwBO
u5LFP05APc2LZBrLdGZD0aitO1IBYEAmgkvxqx793Rnjlpp7tqOp/Re/oNA+6+dG
JPIDRXF3LVgpX0qr9NaMYQ+BVvqOFw1sEODjMJb3g/jXSRlVHUL6tEDJ84kYyJbW
nRfqWW+dPcWhPfv7UawdgZ0B44OahGtviwMfvv3K/H5ReVTNumfshjc9+2QcF03y
V5cnddh/z/S6wf9Kr06l0g+gescHDWVuII3X/zAAqkEU3cNdUM3CgD0T+5ymStb1
EN2U4ea7JwLRlpFlUpEZA1boxRvF5zSkDr7PW2BqCjslZrLD/1mIFI1TsnbeSUh7
1W/lSAY9G5CuiiXgILryRjNoZ3BmkOVz6X4JM+jhFoOQjln4TXJ638vf//9iAOVe
0MBVOl8CXAud62TLrfaCjU3k3Pgl3MnBiR0U7urOyEfUFOHlRZjXfWbQUYiT9yp6
3In/sz+UGGLIDWV4A1WjyV55VmznayJRl1z/mP6uzpt9KL1nGnBlXz2lLltgvVMZ
jJv6Xaa75W1OVxcg828Tc7+LjlpVefAQCxbVd9o62qGojv9kBRn1vG5RpyPGapSu
sag6qNlUAukTqXBz+j2ZhnOmq7wosbI1mC70yIuMB89HmaVdERREFWFf4Hr3GNDX
KyZdpY8JIXmr0/PQ5S45poNs0Qt0yFvnnXP5HEVHxRsrUhE67CNKszAlSCeoSebQ
B29Cz2ik4B+Dfn7/yWeZoYwtTjZjijy9OfQoBAJyyOvIHIBTXvQd5LS+OyKO2sc3
YXtAHhi8iWoi9iCZ9GImURgnmCMX1/JJUtY4z1uUFl9+cG5CXcHIvteCS5iz6NrE
RUm5Hu951GmcIelu07XCTXl3SI9hHxBVOVF0PcOMUmo4I8PrleX3wAWy+IDKMr6u
bwV6xM4xCe2m4MwY6liEYAgK4HK87M+9EEJrBVYFOdfeKQdNVVChZxZ5qtANUafN
1LhhDR5Z2ppjRBymVtBhkmbFM+jik4BcM4Z7h53sj17sHQnaWoFynNXktBabcAC+
wWRasmihlO4UTBRg4RCPLBessSVymGdhb+AXQ2dOQOHT2nGsw41Nf4V8AJLMYNWt
TcQP3lVZM1EgMaLV/XJECHDT0Gd/wQMLDqNFXvBruxx+13pyYDlBsxcgm1SrqLDi
NDOF8t69lVDThvyLid6xEnySH6EATBy8YayyDxYHeOZDb0SgfFxebzlq3T7sKklp
ugzEmh34xiGDIwjDEKchWVIGBlauMn188+MaihfzKeDguFM2VG0wMRP8v9gPSmu0
gtAP/WcFQrgjRholiZjnYE5zoDcm2nV4cqDHItOCSgBpBtSunnple5bwpOUb5tAU
QUIcw+XJfvAnMPECcB2QNpw6VDQDFG9lw3ufZh+Gqg357TmD07OhGSUE5NtW1acZ
c4ClyuTjhMXwfY209PWJDal6vhnoGpCYoHbfIZFkBcVOwOl06RLCHodyhm2hbvyU
SosMvb/jQsJY78cjVjNAMYZ9eKye/5TCkrGbOjUTtn9dSsvIyrrZxlnMpMB0Bkus
4m6VRXSpb1uxvKesq8sOnbKabR0xnnbVYH3yyJASdeyuse6hBttXo2YmKXYwBPtp
OIZZHuOwbngypjlIEf3jVnakugmPzAkGXuU0sPUPTiMZtRUFxGIijPDUKvFJEWeS
PJUYV0O1JmaieojkYY+H+abAo+Av1yW7clomaLobBX226/ZsXkmmOcqMaoqsMU1M
w98kPdXUn5Vo6e42DOyqVz8P+iKUSDhrFKw8C+gqzfPfa1MRMRJqGZEcI5CHc4fc
rJT3PlGUghBFyhANvfD85+8AkwoiJC9GvQBxFs0K2n9Oh7yHM9QoowKM4hVRv/HQ
XNPjkSeSd6fo4D4M6bETIttYHd5i3cm1hhteBZVf7M36O/W+ONGV+Bcz77QKviTo
27+gaxQ8Y4ViDYnZiwhHYsMK7wthIlUoJb4t9+nUkpxR19bWyWDpZ60SUoDX3Iub
9GoAZ6KUY0se9QoHPnNWEezSDIamz4ZzYadRL8uDVgW0Oz1B3gFyrfUJc64ODm7B
gEFROzAJLSPYfRM3Qmf1Pdl0rk5xpjmvHsSyeywV0Peuf47ow/7r2cDcnwl10GID
OrGBylT4IOCciTyGNeNick1kPNyUlpJtx6s4iuk/gmzKwkq7gkR9pSf+arof3fYW
6uEReJ/uJWxNvE1CoSUoQDjkj1H7+kAEY2wYpmf2hUZIeiRzC3HjpxeYawhhAYyK
mvrTAPUv3wTF8dWa58UItNvCKPwf6Xqpo5yJZC/4DdogAwNShf8sAY/0pmYHZgwH
BClghbkojsr82apX/roT/BGX5LfzMeSGUqi+PKhKFJQrS4FOv3SQKvBehV86tG6F
0Dx8YpWn8IgmQQlI5owL6jkM+3Ne0SNANHsptb08qui0TIhkGVq781aw9GiJfJsn
2uzBaVJfFbKq9Ct/n/MsDc1R7PGQ3tjJl1LUZW4C5rr9FTTd4LT3OlzN5X2E4eTu
0zlcDGuA7JSCjMhsTcO8F2VoYLhOUeKL/EhN18OD/W9i9Jsfx7PUHE5wOe4N33g/
+rkw3IaPnzGjUVJq8oxH9fnaA48wLquGYo9boIapuHggaByRZU/CuCAp5s5oQQHf
pHb14d3scnpc2qnbV0NlHfr/WLyS+Ng1MLEzVpZm8MmfvY8xBK9fRfaKz/JBqo8z
sJhmTzkknftLHacLfJR44+3/8rEQn7VXWSPNo52MqqwsHTM2hUyanYj3PKSvP6Gz
V/4FvfCr6lpo7k385kpRQVKhIBt+UEQ1RhQv+WQI/D3OmYMpaIE32lbRrfBGqpq3
trgphaBFLl9OEH2jY9TAqSr0ND/do0fY9F8j+gICaAbWN6tbU3i3nm6RpF4iiSJ6
3eiPVFSnXjJLneYV2kzqAGFQKyf3TwrwPrpsUreQUkyhyctsWYTbdm9/AdljslOn
JyW9flijccGlA4ZF5oPN3ut29yRzdhNj6wWR7ctPCYyLvtErWaB+D98WCQFlrRUx
Q1t8QK0z25Kg6+UsaNscl5IEJzz0G/QKBjeUraz7xxqu4Ms4leRv/wOVBTiogg4Z
YMnht1TS9yWFiRTPneMS8uxKSWMiTHwUnS9iDF4owiCIh6vx5Fg5+y1n64id+DiN
HpP4empsclhS+sbsNdr9kLSORpL2jwWPNi2SlDskZk3ILBuxzamfDLWo2KFa1wiZ
uxxsiZnWYn9UCABZthISvdJd7YBd4+nfHChZgFAyS4Xqc3wwD50U1lNXvrtnxult
n+ImP3eZPAMobGPqDKZ5Gi12mB4gVw/eyAz7BcpQ4ywzLFzfaxn1/Dd5h8v+pVvW
7m9QdAyjWRn/eVbE/bhqVag5VArBgwDcw8J6jcQZcJ+LBll7QlvMHLVaZMIoKvu4
Q81l2Il+Yi63nd0GtUM8cb+6IHwXo2VdmW77m2pl+T6PyEP22YSZSsViI9frh+9P
e7/PpLMbV8tnw9QVur3bJ/UcdplwEpW74iLqTUHS+dRNc9H63gD4bteNLJbl6dga
Fu7MQk2AtnEyvKMqXReH5LI4ddrIj9s4LtX8Ro7gwu1t8nDyA/XguTaGN+hg1aRa
nHkp6cv+BIIIi2rNAw2YG+1BdRw/DQpVMG32ZKyfQbjyYnbBHOAIHsLzyeZGSOWF
eE74oq7qq3mHVQWDTRYhRabeMkaoE5hKoTyq+5JEKdCJz4JTRNz11IlTYCE7wGJa
mbfeHHpuYM5gw3LmA/dWrmQGuNlGzl0z4aeHBCAMdIl2jcCUCsPnkMbJcRdeykle
ZEpB3Sl/LiaVhITgUE4iKYhevIwGkaA97cF5O9pCgAFmHL/A45/T91D3vU5HpCrn
3Fo0uCXgu7D3YxsALF43//fYJyCXAyOUF4PE0nfMXetFcTSvse20Mn9J8foZAz7U
BYRT9I4dGm9HmqNCYgLHhu6pDJkmRJ0KEHE4eLb7dprBmNf3+M1d8BGddrX3afiR
xLC0JGREGE25Fy5S/6jHitwBtRZIpMjPYhxdVsrs3Trs3S4jNSFrLvu/nQS+j3Hs
vzivZ6bmx2a8Z7wgWTQ3XbqYFbjHMYPFsfzK5Y/xt2FB3esXeSFwt+Ws3LaIZoBX
V/Tn6P/chAOEIrogcPOwdZn+IesWIKPahDiFQTWB0be6nLFsfbGJCNR1zBamI6uM
XJjlGc+sAngDLFKRUV3R71zKyK7CtzVpNpsd79ws+TZAhi0369URk9chzrpJ8cnq
Q9E8d47u0+ZxKLoAPJufzChpGzY1ULzLlll1dcnsKdKioKiSnyTlrIoEdOtXGbl8
NUMgIo3kXpSa9LLNZ9rtAuoz0YLmyOVO/uTeO6Hb8co7DWq1uNuTkA8Dm8PlTimm
KnZjTqXnk6Wjg12MTIPvE89wH3ODR1vOCqGYFPnuHqpZoluCZQEWewnFzsBCc3lR
4T7oDs9xGtMmXj+MyYayXESR1pgx7u3zWWXA8gJaNashMSVt7O8nJfFhabBM5mlf
DMl68lVUmsvB7463Q2NApXJuwmxXWqLcVQkbmjtT0h1oTdIj+42XDqIDGpPm9CVp
FSzX69taA3R8YNXvIZga9cjiWB7ZXyQ+u5YPi00v6jb9EObvOZSGBkIbrUYTZMu7
UJcpVG7Ar1Ze+AMmTfzncAB2DmhRPgR3J4nAxIu05xH2hV0a2wurNcpP1uEXX0hX
8vGUSG3k3Q/s737N3GLkNWWpwXykpDpVk5A7DrKKcMSFntT2xVGn7aaRkbXr/dmq
ODJOOpSHFZdepEDWdgrQ+BDvrnJ+2Oe0gpQBATnzDSm6TJl49YXasRhMqPrd0w0H
1oc0fdDMLzodlIGpXDGd4K+aZymtjxH5sbfopeCE+vBoAzDcNEVn3/w2PaGLZhE5
U3fuAhbjydvxVtc0IJRwPDUd5Ji0CGpTCJVGuaMyaRiGfyJ3fwa4ZzdYiRU2vTta
pl0paBUQ/oA6RwlHt/BfUGIfja7a80H5xXrNX0NlFr9+Q621pKN6FvW0piHfuu45
ZYNidnNvEZGS0gdjLlFp5DJ6z1UUn9QgclhwfioipOlukqVSovCRHDzXQQVd+ZJ5
o38ro0DEcKFk0h8cRkz+kBoz4Zp5FE6YbsVymj78Y0c6k6TPlUk4Ge/ETTUiTO17
QJf/LNy/GHBBkTMAVnD0OEZEjAXjxrFesyompudn7iOsLIbyq9M9yzWU6r99bj/X
eCgEBBa74oppcq/8O7jZDulUjr7t7s7xRkdFSeSxNX9HFRTwYIN+to9EJVqqFPYw
9g+zL71+iOXJZMsM/JRA3MLyzcd9vnT94dfDNJe77t+JteHCfhX1Yzxt0uzcSqTC
sDO+EKtky+H+9RGPXxXwtpsllRrgXg4Hik3oEu991fclqoyxfXN/k28fhEyklAdu
Obc3fsJkOJ3nclV9Kf5GKtlmVdK724ea/7edwEBbzBoaeCdNEWuLHE2Lltk2NTOU
ly8narV1k+Q4baywiNCV0N7mKAwPVpSrZdVCKCmPHH64r25UdZbCwxDhiNwmfO/Y
MjNAu2HAUtwfK9BrcmMqNbfr4vr+foZ3LqjG2kVQSN9qmL2dhBBgrYWQWL+kgvQz
YPGd0X51/5k6CYhRKOvOX2ZirAG3ip3y5zauC1GWge3rQrRUW7Wo8en8PNyKmXe/
4VLj0YgBU3dXhNsafSK5tI4AzeO3wb3MCNw4hmEKG/Lpe1badVyB8Wx1iDEoHYm4
/NMcaAGX9xs1nB5Ps2OLc/OpENcrXF3HUpBl2PCPet/Cxa5QKKxSKrnqxtv26BJZ
KAMRHZj6BXNjfYjqOMtg6XsB5jGktd3EDBNEhggLS+cfNOd0CWXh01cv4NEMOai8
SL6PceXHTEXkDKY+7c76p3Zz+RUSVfUjrT2gc++Y19MPDy0ldi7hlVHInedcZ2ky
PC4CkrcFLFoJGH1EhEQJA0DWiO4McheEE+tJoOfNGeAQ1mlG4K+SsTb6t4HZaet+
G2H5QvnKUZuDWGo0y9VNsUPv0itJ7G53F7aNk/U7cdKdVNVzgqAVJQZ76voUoEsw
e6Gs6Yxs6l9BzVzio+sm5PrVkUM+nFpuHcFNz/JJW5udsrLHAz9cabWLvWdtqIZY
IEqbKXuiMpDlblkH0ND5aDy22QqXJ69GEVJEYYTpArGvM/cPWqIweVKtZvTacFAg
2k6Bu2HhwkkXLobmG6/ceghbAsWTraHu7t6R96FxM0nO47wnEsX5Au1/YCbGCwOY
4TVwGr0M9CEg9GV+Mfo/XjTkkDag7lWslaHXPzfiuhPDaTsrRYOvCu3x7cqdWFoY
6UMwJlcZMAPFDG1mCq0FsmipVUnVJWUmnwS2QybBxC7EeGnlPMjwERNzkpLwIIFU
JKzHcHFMYHB45ZYF/sxeLb4vLq0L7sxY49nyek27MgC+Jy9iYqpnuA0TYlrSFT9k
JfW+YFAKx8SG06jny25go7PFBczdY30LXB6pNeAY4hDPeDSY0vp7xChnTawVp1aT
QxH238zi230SglEyl9io8pTV6Yf+F0cBA4gwjJC/zYQSc9ESW5eEX4k3cpUe0GiL
k01Yus6HA4CtmGd3MVgOj/nTAeGQL/pb+3YSempugt1ZB8DevvJr6ciC2KJD2n70
TjRhX9VJyKyx7B6QHxp/An2VI04TdhtToP2lUCoLbVx2MZUDVEEThQXX/TTYOdL4
YARqNAOPtWY+O09UZoOHZNQS2ErFgBxM5VZT2XaBhzTtZV7fEMmj59xSWn39I3U1
vOkqQ4ISG81Nrnq+SfZD6jI+OHmGwwuuRj547xkMunFJ4lI5sxJdpceEmL2vunn7
JKZq33feUPhLVYZGnnt/zcYVD9k18r8reM1qyywYAAf3chYHYOmivTU57s4ySN+9
T0J1DMwg5VjNbVBbYCCY1vE+fROnvwX6SN7RqK/rl1jQWKa35wk2BdrTS5C9FTQG
hWsDLLPnDNQ3XaqIQ6A0cvN5cnepB6dAiSPMCVMX185kJ/LLKELvxm4PhkgVRD+v
rPo10g4YuMHT4FS67HSfJP7OgfVz4v1UKXCT8SJQuwYN6VrhRMd5KT/oDluChyva
KtOryUpqbmIo1potY1qSFXtUK054GV5zB+eI9BVw6a39qnST+9gI1tzG3cNH8m2m
OtU5E40ECw9lBrR0umqZ5fgngCSOmE5BevxkwASi46I3ggcdYdlzLpf81CfoMz0D
0ZJMAGPVjd8UcXxltEilMydY6pogYyYOjGw7/0N1R6+wq8nxvO+iirhh8qcM/4vi
9lNzRanMMJm+R8is6vLdm3fLeqLELT7qWCjw368/JVeReFuHp9P47tnJPN/2fbOR
dxttciK4dn228c8OWOcZbBebQKlWbdBaYi2GjGZWCqSdq82U9QeaRCA6cLjnCuej
0BoKr0ncB+jEftYtrUiA80rZWUPOYkDGy7UvR5HvkfLUz/fzNVYHVYv7kngeq0+i
uRWGo0pPUPqNvL8pQHRj77bfDYuukjAp9JuCuZuR5/lV0BnOq+qzHoJxo+eiMdNl
Y7InZntxPEto8Qk4ve4HIywQJzcDtLtYizj0wD/m9v8C/Mvimik14Zl87pKaPGAj
epn2p9UuM+DMV0TL6aCX7wGkYkgSujJWHZ6SidkZ4O56dgM7gebGP1Md2hLQcN1b
DxH+g6UMsTLSqVNin2H4gB25hlcFEa1apVud0c7isOxeC2dk6N0DdkyB1mZnR4xV
UQJ2nWp7fnvuZYliH+QT3L93f7dSp5e27j4gQj0tBkog/4M1s5xAF/wgLbWu9QpM
cUJE2dm0+H4oCawk2d8Qn44ixQl+VRKncaoR/fs4AsV0QAhz31FBny8yls8mZTve
GEG1nRvHqCCbGW+8VqdlBJ0rgGL/TMbJ2vYOwB49wtYUNzs8BiMHfzQHJuGHAEVH
glfKjt4IdbTs4sDzeJnY7N+3taowXDCRtlusifnEPrc1WgWoA+NuRq5XfstQRSC8
UQdHVXiThcGoS07CLSPgHa1QOvomMazrdXXcOn8Em0I1Un1AVOf0YEfYn4dkNT49
yHEVW9cdT+LYh2sr7MJJRNQt0zHVTonwuiesxjVelI88S/qIJ/NOQzyerQEIBFRi
q9vsFsR0plnbWXoThQuVlGi1LhDubvzwJaremrwYSnSBDCIr+W9IMie91qAfQ5H2
JXGfeciDX9LLLfRE3/J74+tcpYpjOwHCCUHgOGL+dVw8fJg72O4HszvGEqVSUNjJ
5794Clt8IhgQXq3gBY6wVFhJfTnapiRNQknfbfcHMwa+DfkEk/hvuw8u3HWFjDtX
nou9xIDMTctllFNb+sOSzhOap7oThx/wvaMizUowPJHCvmhWghn8+1daQTX+Rshg
W9KaZS7YssyhNh9mcUAjvisG8oapXvq+rfsRmKUSS1C8/r0zSZhClmsQltzEbcsG
mMDcRhlKvGKG+buZi8E8XY7KuB4w+Wx2ymJG5HFukxi6HzEBXmzHH+hDfKOhTD93
DmRzODhaclDvR92tLtmaTGDx9Qs74sjZ/00u/WB6xacCUX1J+nkiZGtsuGTuG/Dd
9zihXW/crs1Y/ZL9+jH4Y4wtFeCg2Ske0Swuh2bCEJDBAbEC6och92lMHx2RUdrt
RY8AMeBIweE//EhHz4QDzdAf0bRCxHvSt9qEzZ/9WKyy5Hrhn1KAfa7lktqkS5Fp
P54kQszlcsfKbU4ogejPcHbL90WCWibztR6CmS3NNrVt+VISG2upaN74i8k5s78Y
hq5gQ9p6LbYMi8qrcmmE+AnV6ztlJJA3k8941OlrLLtdnuAGiwV9wpkEzHPy59un
NaHbxttXf5FgSdUfOiTklMgH+L9ckY0bO8aKSG/Rq++4eTq7NJnRx83RY4wWx+q/
WXuuMvcLD6Y8E+24F8ibSOrdF+ky5BXfCiVYOeVFSTzsVMrNJQ1jHSleckq/8L5N
wjOMBhQTsYzd3IJPQ69cb6ppeZsJK5+Ctki7pVeAaXuKccMbelI1lsmgHkQ4CWvr
WjrXVq2s0luBjxC4hCz+8vBAPEkmuSayEXfiVdAT9fN666vFdEA3E0syYfwI3QTI
/R2K86fIB20/T+HWmAyW22m9xkHc4nTdbTI7xklOqDN5GfgMDq6f8vvpyTyH7L5D
sSCX6+bl3bAXT68IXxXxmBK0x44DYv5JJV0Z7ojdCEZu5OeMuh1Do45f7fg7kA4r
S3HH0SVWlDDvB3AIJZqhHIyRDNKiW+FltBBV2anZruajkA3clhMkji9pFh4EaZfI
noXA8rPMsvSk1I+TOWSMaY4OCU901ZKUgjo8WJdW7BqXJeVkuMYefPaEonjAtWVd
1sQjOVC4kWDouhN2leyRUCL3MJXH0AzLJ8FwZCyT3Dm4Qgv0oCuvNf3g0rLuTTTd
cFb3OkQQKZiRGUsEaf/AlDs/737NYrsT8a0PwGOayfk7Z/sX+5YZ78QTqsPuWWDF
B62WBKbT79HjeuR5WrOKp65hGHrFtYf9SJMCBpIJCydBn2W8PCD2+yVMhfNRVDFI
vG9OYY+e56TkrMa9UKb77mCFWze8Qi6RRKIbL/pEodhKkAjaskAPYhN3C9MNS9WF
6Ax+Zsp4nOn08sLs0CcP9IFo3YU7LUfD4Av7G+tWmAjY7l1G+D88Qlm4q+OTVry+
EPCCgLCoyAaRQ8QORjyb3/HUWbt98bRTWRmK0U8p9WWp9/mJ7LuA+6q0f/gfwV9P
2Hi4FTglbCTsqGKTTqfrNScRzYYBuU1lav0aXVkZDUUM40H7enf9E0+LB/cT1wEP
7UgBbKTwMXgjpqupHJoMpQc77pHbevdkXYiZwRDt7P/44V+P6S85ikRXNRZy482U
GtuNhaBjeJahkx4Y7erLaG1n01dToWYqzC+E7ukRZOAWc4M4fi+u6onaVCt1sfJO
qtQKILx3j0+MwYE85C0Zp3N1OkjqLqLhLCvCJi32O7Hpy08HXrxYc7+q7C0142tN
BM77W5KvvWYocupcez9PPHdHOx7YKQsqXGPCpf/FyeqY68/4KbX7y/PLnN6IW6VU
+7arcJJB+Cbw6jGxn0RwE9PnAiDkDS0sDP4QQKxT+jxFujl3E3hJDyNqpFsuKgfq
T2u/aWWr2msqHI8SLP/nTLsxe7vegPb8S6WpS/sUwrQVzA3OaooOCQltMTYSHCmU
t6GfqcNBoNLdxX4lBfabccgU4wiq0KyPjTzEyntMvhYbrDGf937Br8YN5AZ2ZeN0
uqV6huz+jJNL8LpYqQOWPc0omQMaFey8l/bPChJX7YI8rRkaSWWTWRorVHOOzjuP
6USjfQ1/6jNw9CPt+PRZTSVm3QRgKVYhhndx12Neah7EFzLTqdJTRRiNxZ+cVr6H
Xnp8GSWaOfBN3mai5pw0JXxaU2kSLwKGJ79Dg5TxkCyj3xAQ7HQ13ZNzOyUV/aOh
X5hnRUNumsYr7rOEj0MIq56Fqxv6uUBh8fICtdyZQr9GLVEsT0RfIPIeCCD6MsMX
F2OqzyXSQTsZq7/V0Gq2yiBFrAT0WT+Ser9VJZWCcy2GSD4zESgBcU+W+m3xon87
68nzf/vypvSF4isOxcgVnoxrOq9ZLMOeb1F04L6qYUZ9wy0yC75sqv8wGZ4A7u0a
yZyQwrBGDPvgTcCVs/cWZi7ey3S60BItj7Zj40JyzA47KOnFuC/3XZWs8Gep5Fiq
diuCQvI1pKrFy4iYlYrSURfiGCSsT9UakhiNy3gNJ3ktTdXIv63LV6ZBzrqkqbrP
Ji9OhFI4UVJtuzj4/IFUJaX/t6HPh8haxKuHGtXtNVXMpVltR93JhAfsFRSckoMU
MlYm9/vaZylZnGhoAgy85CJpWQbM9cM0SjNOK05GmfqlVSPOvS87hY7dlnwpbwNh
8fsv0nSZLJMSoChm7Kv8ylIYTSCQFemQD4o8/xawfClZ2YMaTNRbPiQFA/4DeJPV
wHz1VgBgMnHwUPueL8L/7H+PHenKEbmrIt1GMsZ0AwarJu0o8c9Wr9RvLiomD/fB
+/wHtHASaVTkJmIpOHpR5GR+9kWUiOwDf0FGZ/Pcd4WB+TqWGJUyie3t3QhcWBOZ
wCvXQ8RGrJfn17iES9e4n+yImgoB6Is3hPpwqV2ArkVJplnmIJS4V4WfzAP7zKWE
6/EGhfcRvj9Tz7VXc4ut2OiFHPcCVnjjXuBAH6nbeSZC7LBCI0s2Cm6e8gz3oUz3
V0+VV+pKwT+WlgyRKpyaRbH1iUym0rNiggHjaK3+amXA1te6ftlzZhLkPEmRkB/j
atyOA76CnNTs8AHlBC6A2K84Q0uuuNX/PgCznAU2QMktXRLqloQss05yiQjw2sQC
X94BtpgblOpiMsvn4uPlbZqJgDg1dfITHYo0jCWkhbPMwDc0sfZHShm3ZlXJDenS
9dfz9zYGy/fHLCQ9BXEVXWZ2W2U3jWdp2JMt91kg7J7/HQ1PriQruI+2DVhXk3DO
eUQ/kcnzf3ZzeaxtczSaYS6SjUd+7LKXh1rgtENygNpdipmopW9WOUpP2ePGuUtU
7kHZQra3c0lJ1+AOwWltBdrcRrA/XTq7Bfu8RjRAbAKD3yQxQnt4ejN2aP66LYSP
c8wI4Qvm6IWRriA9ncxHuxwxcj+cJL/ei2pNwg6w0PmLqV90rk5wchqSC6uoogjK
SyWIeyZDhzhvY6I7kVg/oCKfUA5WLMGe6fjgGPdsRPCirf2gWzPfyBg/vN7tQbfz
Ym0yF4CPGHEqLu6m8GzkXqSvXFfLnJXa8WAS6XN5Z8qkC+bPuELj3K+QMbcYEjfQ
2m1fgkDbcmVoltp22KH6cq+8wWXU+mMd8Ot+t5Q0Ww0aL4oILP3aN3YsJizpLgEn
FiCNwvvmp7TznJ8wzIVGjstz0ewAmLF9eOXG/EjkfnxMaJMo8P2rbRNdEyPDqC0+
mrKkYgpnC53Oj+y6dvTznCaoD14fYOTloOLzyrr2ll48b8q7n69vUfJjDT4TTQZ9
SKj0FdESW+pFn8K/9OWki6n9mYDkS0a79cc5yYIGICgjaQpJmWkir5kBgcM78mlX
ybIWY2CChBDISiqXeDfguylH8qAd9qahsz+CZGoo7aK8eIXlPM8bkzGUOxKUBi5X
bQWJ5WuQ3yJgaaL74OUVyETUKGV+SsGd/nNo9iUFc2P4URnoSCRS1I7QhVSSFwIi
Elq7IRlUZwFWtb+wU7/8MzKFeNerac23vW6LtgWkm+Sy9udh+eIRM1aKKT8LTPXv
6Pj/jf+11WRebOOMbdYSz9qkeVfuT3KQyj4aEpMzSrDvy/UmG79BYe4C9O+XiH0X
FWy6+iJx18GCu2n6rzXl8MjhE436SkBwOiG2XZLEu0SK/JP8oF41iXAI6gF749MG
M9si5pUenAfVxk2NxD6mWzf/IovMZ3qwj5hx1Uw8IqPb+90jsjaT+TWpbwhivQAm
MKVIP6gzAUdbL0spfFvo3ZCKXHpwSv/2u28Sdth0du7C50OJiov+WC0cqjeO8zjj
zo6Y869FpseWj0/9mQuviNHufKZQnelIiP8b4OCNBNdodZQ56PCnhLLiAwsONQZK
xjqWSwhvntJPqtj3WAD0lXwYTi9Tsc8G7lFTZN3TZ15gOgapw9f24q82NHjJlJ/U
fc0oAGg7ZFyzsvLxNqGNHs4+qIXqDBWJqscaEoaRpPri4rs8nVhi2RL+oq14IRvk
7VzADyFOfAyTttDWH7iqfl35MrLQCV7ALUeThQQjS+3aSmw9HDOUTneLAfOrEFWn
NjCRI8fXNq4mngDjyL0VNrwUm6ORk6a5dk9IIlp/cNP5+g23M479dYBbJafTOWMH
yp1TWbHT3eb0c+eT7qdLr1u1D51gEBmarKP+0wcECKNIQaOOqnI2ZHf+pKOznP//
rtiRJjRnyHvyQiILT2azlcWspS2S3iHoKMFpnKEDSCRs7ZHhvqXm1Ye3LwN9HcOr
bePE9BLPEiGWyNhoCsF57DidUPb1CE6CltZTx2mOVVlf3szwVoTwKZucilARDrYv
ZaFHCD0YEFBF+2UFVm2hE24sdRhu/GOnmQzRAp4Oj9r1j8Mjrt+40afD6NvjXHUK
GTOBG2JF8pospwF2a3T6UeD2R+AhzGemRRgJtmXpFviEUWTQ5Jer7x9JV4gRcGTQ
AUNIUD7KoB2AEnw96ZLcV/VqczkuwhKVKr5yuutwGLmbKMhvhTd4iFpaGRWhnGYb
aRFak6UM8UuhPYM3VCU1l3MTYHOl/5fNXzI07veaPj3nYQk8d59bZR6yUDKl6NIM
nHqRy+c9JIIeAnqW1dJ1ZNRl9vjSCLISAuJRPdsr8fZktZ1EPaNiXZNsOXDzVIcc
TKkmCeP+xuCYKZxfpQ8L4LYgj+ZLv1GXlyzIUFNsHpl055s70QHKT31zGH1UFLSP
OQWG6QxKoubTEXhaON83+9NjYEDDAW9Zrq9ki/tw15MvDwpHuFtpYBScZzP6FS7g
h6COm1xcSmqzizYm3kqS3oUId2qJC7BKqpc/wMb1UoUh9QsEMJcO+Lc20v0pQOs8
kZZPPJH3zXdqD+XDmiKr7aq62FM9OQfy5YUtRZg0WMLh33Nn8E3xKOgONwSYPzC+
mBKMMgjWvaBxwnrDldZ6l/DDK4hVzB57CQ/h/LRm9NO5+Ramuas90iPJcOeqe1NU
8xvwzxQVnHl8dT3x/eDQjHaHo9kK3zuu8RVJIbsqejZyTHsSO6m1bwNEnQEvnR+l
cqpoQbZbWnKy2MDZfFsLRQtjSAciwSj+mOFKL3CTVf7gWVkR+YEENWPNiANyR5fq
dbWf+qjMrII1EtzhO2WtH/aRCaIabJDpgXWP38UJVgidyIDRQpagK932uQn87J8j
QE00u8b5CI/2/86sYFAzfBdwN3cc2BaPWhjRmxpAq3MVBV6GVjt95NMvtnHF2qs6
8hTKWf1lvZMAXhbMTbSKmEJcr9qbmwPTGGaHl0BUtUID2HG0/x0uYKCKRso2yiro
cywOQLKH+gxjItKUopCGbsQ1D0344LIGGNq713zGjAB4tlsGxBTshRm7nXrf+Ri2
pgrTMPSVkTpIXJ3bUUc5ooETV/fHc4rw01YvDGg5S4ihIG5zvour3wareCl/T24Q
rNQtuSqi3jIssQHVIMwSj8yoFdVtJLPBQcdUYhPHh8DqcteWaUvMrzv1bMf8nLIW
jTqKrqzWtHSg5ETBd0ih2KLSbgxItKgsKtZsuUu7hAT09KoJN/oBdxYlADU6nBHz
+XpokVzg2Bfgphc97NWwZItDG56t4nHTnyAmPw0qL7lxWLCiW3jABQE5+/Thqtu8
By5pSc9IDdOwCk8K6+Yp8Lw4nRfVnJJabw+0kh8mPaJwXFT07Vg4PjAPIPPfya1n
1XVeQeJr60+4oB3ivrXMGSZSnUkKiY/pdcdGP+IDSzYhxE3AZ3gyBnG6ZzhhU98f
T8uv5Ed+FA/x5if+iH+HNMEMFkMhcjZNiyphN+xH5LVhcFQnxEvIksgifQzchCqU
Y00qiNORYO34D3Zhs6IKdPK6CLfPGsHJdeJEJP1kX99is3pwIgvjGs316ttL9ey/
c++5cQsmKrkpSbtKZEBTeSnbh/QiTOZOdEktLGG5Gl015GIMV0Qxv+VT6uvM7oJw
AGoR0KQZpJ8vo+RUnTiT1h6JRjoQ3f9lng4JladH1K/U8w5s/xgRzAXK2ho8qBqc
HHba61TEoJEe3RAnZTBLY1xCwqf9HbZctv5VgHtpjDiWH563KtC/Jcw8l747u+98
K2G0TWg+GSRHk6ZceLU4RdYl8fiBI6TkPmvDCnSpG/13QofARA9Sw2YDNODcj0Fu
HpvbVeXiiDs3HHmu0lfMGWzZfgNVY8x4W010rv5H8bT+jwpwf1BoxRM/HDKyNgUo
Wem/H9312hech8SpfsTXnWoGNMhg/wCB3P9LhnzeSw+G4jlPQIuozz0H0ZRRw3RJ
x/YnZ2P6amrKhuoBkaOAmDCpdlvd5oAzFZkod7cyJlb4cOol1bfIWxTPL0ebty8U
oWS1gmFlYFQGNsdBOIIwPyl9PSHqNDM1aMYo8m+oOGi2pjlkIG8F/uMt+v/wkKIn
GDoe/Gp0CH6MP/sSS61ICpeofefVR3G9IhqhKczPzy5SmhBIxDGaM5Hxbtq9Qqv4
EtfahnpQ/4hAcbE/edawz6MzRSfAk6SZlf1X6NZu7YRIO9TScLn57QIVFPTqyY0l
ogBQMyi2136ADpEv3YqRwG0ZPsqwQEQiJtLkZa1OmCSH6D+h9jLKBqOxP7zMaWI8
gDDwSP4NWtARAGXZfKS6MYXwkbq1LBrlNjoG4oxwsH8SxmPsk0WWdlPf2GpV4DdC
KK9aAseZblxvploLXOk32iDb9t90I9RFSdpcXr234i8/yFg8R3MiJLRaZgiM1J79
uXnVY615LxdUqcGs3EN5wkZ+8n+LbwMdRktZ9012eLLqhIuDGo2WrVuDoMrZq198
YRunyl0sG2N5PPYPOQbm0Q3miQbb9urWRIlnBNtMEBruYTLVkFNA7sAnlW3Da0DC
pcU8vA0Km4G6ec6yQL/LN+W6EByNFCVQWI5lCXCgr3+LkiwOT8UAEMGKidbMnDLA
o/dMmW/zpDeQMNSb9YXZ6247M8VcHmARybOBbmhrz6XKSHTxEpPygCrgChfBRV1g
0Y5f1vzX5i2zAZLB6ygIy3rQtWJVyGIigC8lMZE2bCko7CPZVA88LfpLLJgDE6Be
NBfCIIRXFrRW0QiJSa8/fRFz5QpSghNMFTr6uWVIGi0qjg4Vhs73k831tXXWckJx
v2cuo9Ag9QL1KINmJvgVOnXck1g10UoEMvAxKo/pohqW8sNanKoeDk39Dj6Fnis9
LyepOPq+p0vCyMc1hraUmxwwnwx9oEMndMHkVMDHfpJF9pkGbqm12AKjjVIUG5ZE
P8ei2RxMfnsBR7SJRokX9AaWVjnpG9+gMwwEHHSkhZ2SvAXoVgrat8whQcjZL7FT
DhERiXUQhxgOc/Ejv8dRxTdvH87o4ThMBfFzLPfTrQcA/wPywzcTRW79beEHpXqm
K5ekcoSbYDHVxEZpwmEWLn2SyP17oY/nfbIeUNlrRSo9BvIbGnYTFKdDM/ExTDvU
TB16Bk5qo9d/nVa+GICWYZzp8sWH9BGmupPWdDHwH1pqJV26HysBc1Mlj95Bur3F
YkeU+aldACEA9RR12Cgs5iYRx1/tv81v6E+/KrFc/G6Rvpt8fujdloV+5CHd0Sx1
akZNDU/zbbwvxE4G9k7IUb7+YhExiLgNUPMurOyyuGewM2QdRg4L5QvcUrRNkFq6
KiTSMpQj4kuVFAKQoos+e+/fhrYV08hmcJcQUMgLQKRI4UZd4IUMGx6SCdPNcYoI
XAwItzfdEmB9hZs3L7E2gPud7aM87PhIWcReT9wjTzFHAK2tPva9zw27YjDH8ngd
zrJz2wAYX+iVMU1nAfYM8pKGtPh+Rq6U0tF/7lUueT/h2WfPlnUqBkch1YrsPfrc
W9uAdM/UomR9QylfIOG6RvOxBr1pY3LlwrTNOeIrD5Hz2GceUjSKB7Athg2JCNdD
/sbEvaSySGTVtWBdq2ZkGQLiFd8Zop2LzM4EYdmDklaSQ+URE0EXsfc1vymeN46l
VxEiz9kqTVnrl4j7CEwCB5aXKdeByik40wX6F+lfGPjMWtwJdo6FxfUxygMAlrV/
gIoEV8n5Bdrugd4jK6o3CgkTitxTNojy+9g4DHVaAdsezAgFGH5MTCrT5MexrukN
XIRwtr5/wcn0axlxcjEiYRP518RuUyCo4AQBqrXveSiGY5q8ifGyrarpqGPWficq
erJ3mqe63maIKxS6HJVK2HRC9tIeo8Gh3AH6VLpHiM85Xm1a0/ohyxNeBxNMDx0a
Q52lzoNvit/Vlsid1OqNAfId39/9dAxrf/2qPQQZ2FSEfh1VXT027cthIWQIle79
u33yRNpjKuec8hBZORsXtep+7CCQz/Hx4hjApaccLMaPZ6u1e6twpyRSxsVXICgf
Vij868zaOZOPqp2xvBHgZ/uly3bHBnFckB8eF2FzU8hnhVnDl7r6TfcEADSHdYv4
9v7iYBSUP/3pIGTyJI9RhPR0vX3JWfnVAEB6n+e+2OvdDbSMvVDi5NyKzClUAR2w
Xqr4dCCQ9KCfsTw1kOR3To7esD/RivZNBLrXOJdNAv5YLfo2shd5FYpUtELpc3V0
Xbep5dWmos4m+AHVwt6XWzvBi8Eoq7uWqgvXG5pFnA1edKZPsgeuwaFmAHry8lgQ
pnk1V3eq0z2vEx54S/HmnVd+3kgIEULSjST+ZqAw+9v0aaT38Gqj4P15+FjUUW5E
KQxLbBbHgekOSTt1yoCfj+KqVj4DHkdpZWCCB82djYVxYmwH/uamKQGmp09x2pal
ymGGlb1dYpi5/dEUwvkKpRppVdf/mL+Alqhng2uzVVyeGwCyXgJJUR5jjqNxKX/K
djzK+QLu0++/R+QnvZYwmBHoMEd4cRAhShHtWm3lJ+PeER5WLLlhjsL/fzKFtS/z
+kLANMnFw/9UnVM2yl8wiqlhRxecDDv6uEJgN5pyYmmqeFHa+/RvDfavLDo8ZepP
WjQijaFUrfJx3yFGDtgP7G/VOf3tjVNDeAH6pOvFOrabn1BaaQftOltXS60cUgD6
Fo6xougb6+898HOVDfREO7fTSvCt9NfxJBp2YdHa/O6drl1Eou0+zXnoytGkRxi8
u4kP7WBYUKnjGAV1qXiXM1ElioF6BfrEIt7GnZ+JbGJpP+Ph8Sfz7DHW8BORuMn1
Xu21AJPpNiJq+chfILkU/SZRDSCLYBZgRSTQ8bxykvv4RyfHM6TFF+Fga8HKcau4
i9ygLiX/HRmS1kOkTYxDQ5DWdk2WI4KsD7s7tYXfWbGJU+rRWfsKgSskGW9iecXu
Fca9grkHAcjNo2NWejwWM+XC6vlYt6LsFC+bZM9xIXINMrHCKcanJTmwdHr/2j7G
FfDqmqnL0mn41gRhcB2mfUGT3b6gr4FrU28iuri/cnQ12y0Bx4j578xqP7rjCf/e
aCgvmtPKI4iz1Boqq6GEpx357M6b8KY24j55KmfClsOLeBAdLKbTfYs36FWbJCdU
sq4RY4mAHnduG6tunSrXxREZBZioPLzQjFd+VbW/R7HHz6emfr/KBlGtpJWlZcv5
YOB2CeyqcBSQzT8JWXrljiyMRCwE/mWzYRBM780WB7Q+1lo4d9NMXiXVXSo94dQU
4yJQSfeQBWRltYoZkJ7tzTWtWAJ2rxkQ28k4xTQBPnTjZmWxeJ0RLhjiAe49b7nr
RUZm50ggfArvbrYRFN5vh5hi3yzXMJO6vOQQ6gNKDPU3aPxKoWhDtn2S9sL4oTo1
OJP/JmvIN/KPXKqf7wYW8d9YPWKyV02sRQs5GjjAXqlXVWyHcJoO/ARPq2kkAeui
YRAdouk8gnq7dJyR8s/kg6ovK6lG6lRnrlqa0CcYe0V7RbklwcnA/xygR3qw4L0M
2VVynCkzOVvNqjg4zLdfhfXL5yGjs0WRtrehiYuD8nidXxW6rgG8I+6ILEIrztPW
ae9pwjY6iKiIiio3KKBm/1jLNsHqeIi89thwNVbOvWlgnkhVH4TmWIqLmQsM81rf
9I/jMQ44W2UcTXga4XwbORXurS1pfyZ+eeflivE8wEGeXew1+tGyzTkbb0lthAvZ
xyiCpiIPdMtpiAZPPTHyo2aKplVKks1mz0C4LRZ2K2oevKNQtra/OpQJeP9D7Dtr
9KDS3iVe328rib65dA/0wpRgobFcgXdWHvAxBISfEy7P+oLwFNmjidaMUdvoyV9E
ICfy4XWu/DFI8luxwZTVqJGzsssP+O3/v8PlpP0w9GV6iC9ZiNAHXSL5nG/sIydf
tUVey8EJ3R0zkUuiUCA+hk8VfMI8MAVTkbrKRjOWZFSKYpF5ZDXgTT6za/D2MGVy
rBOE0NAwEUxy5Eu0FjSJHav/uO2Xg+yxHmrU69SQcxc6R9pCW9iFUM+UawvaUcMY
ukhRp3h2/KlFRVcVw5v09Hf/4mDkgi63BvjJvjlhZglcYOfyQktQVT651cnOVzj9
qq8KVpv94C8g7oDaK68ylzrwkZ9igX2dySjHl9HmIQ/NEZ4a35b4oRJiSqj6sWyX
qVhBW58ZQYmB//i1Xvw1hQ5GG1z7Xok5wqb2m9MgDB7fnFeYmG4zTin466aTuKQx
ihVZHgKA2OyTxh+q4V823kVzQ3f6oeoMiYyaminzzEC0HrC6A6iZHJJbywsrxgp3
A9p05y6KUa+xUUcCCNgwTeoiUNxSZufTUjdwkY2bUc+4YWoTC7es7J8YjOZW7sLe
NdAhsJ6AtCQLpje0+VMKZK2da2N2Z1hqKNteYY3zURQqyjcBu5bYxjPR8LXYkuDF
65IsI9PHuTpVTZlU1FyGulvKNNT+Xav+tDWCLqY9zInZzrj8+epaRWM+bGL0kHOh
8l6x1bYck/bV8Ij2yV1XEdAXzEVah04h7xw2kp8QIMxfryX3lxiOnuE3QduzYEXT
lMX/Yt2Q3X49fzGPLYJAd95S7R2f51nsccLUuQwFgFfisBLc86AVq5tVbRF2fvaF
f56ZgJliJSDqoovWPmT5rP8RjQycxsY53PDJAfDfoQj6nakEf8+3HnkGQlerrsJ1
PGA00B2L805PiFRCgzlsJ7ufk5KH2La9VsIQppCqORyDbmnz37ZZze69QE12/GRp
VoUZ/db7Gqc8jCUQnAEYPe8SUmgblsLASX1qiGH9gvNVQQtHqyUgaGYYXvevTMOx
sDSALOknOFMA3YavOLGsCKFdKuSk1yDLq/69HWxX2y9Czm+haU+Q7KuMLBeEKSe7
K+Iuvz0YRW6D/XRwFq2Kcm1nm1B5R6HrQcrQnaKEgKCJj52IV3PbYUCCuPQBf9yG
nV6FNUWp2GBfBY+0hiQkLGxAXbAo1stsYH24+7o2T4EOnXsqy4JJsM+JhWIt+JoF
P2CulJZmVeead0KXnL7cJdWkgYVTdJErM/uUIsfywAy1HwzIegmZrrF9/QviCmBp
fIp0RIdmWXaMB3DTUEHw2tshuWHliZfF8Omm8aF2CuXsSFrYhhVwQpznVubWTNOc
C1th6tYaQgYDBvxITZt8mk2DHBEmT4aMhktU5kboYviIx9/erm35Pcfd/yjHdvpE
3QzxrZtl26z7FhH4hFLJbjsnoZEmlTBef83YtrudqohZ/mf0FrmAn6Vap3/WK/uC
aR1I5+6b4uyHgBL6XbwHXOnwr1dqODRVjQYnT4CDbrM+L71ulmEwpqzd5NG2aGqh
s+y3/GPLF5ChJywJvPgybLT/w0wxIQD4noA2tEv7b1Hm43yj2Hlp4fpi5LisAPnG
MsZKUsGye5i4YQCxeAiFVZMIo+tn362X/v6ZGaM1pyv+YSE2EEfwFd9pweejXF4r
N1foXb33bGDtg9mOEvGPT7/BUIqYtXF/4PQHkveYemAqCoWi2T86X+SJSO9AQXUd
r+8x+qDexDOJtBNFRFZjeJKXh85U1aZeWUtx5dGjPP/8h3kQvp0kPIDgm8nljRTw
J4TMjI6TrAp/7LDXYwtMUfpZLH0+age4YaJ6w1hjoQasC6MLIgi1BbjjgeUDwDSS
Kn17/DyP8MiIAs9VQL/O9m9qP6RXYme8agoQ3v7F3k2ZhNAFZN4fjjqRlbKYBGcD
R20kCTq48pw6xtykDjU0fwIgI3QzPuiVTrGRnYMtqvia00/h7YnnScVSKm4QpwGl
0oph1dvwg6t07AbdUKPQiXq09+ArjMPtloYnsKzBv06I6k+m34h8oviSgY0IFYI7
KRsy9N617mq8tqYmi4NzeFHsQptv0N2dzPMUXMC8K2fBxgHzV4eCutX4RQsuOUbZ
E9tPpb0g4QIz4W/gcRNigsgwa3cPJoeQcEHu7Gw3X5gUP2P8Cp/IT0Afo0m20oI5
LPdIo5FBapZFZrqpo439CEPny0z18aq4axy9+VlScYxE2abs508eNW3XP7ewhGwd
ov33SpAy/L2jdsw7CnW6Tw7PS1+bW6nqpb4oepfOd6MENAUSiqAppJHfeIzLO9K6
O/wnRTAMmDDHCQSxgexg0w7RP/Z0FKPU5SQ2WbR5VLrlUYZ/9ahh+FGJgjeGU6c/
S9qX2wL4NH5KEXOuRdF4+xBz6Aw47e5sS2y91wIco1v/f/X/wuUYik60mHunzsdP
3y8IsQ82Vmr4dDpqJ7V6t2wLYgsWGk8pQxR56GSfvXfSRV9h88RxL2h/KcNmfmhy
w/LNnP20k1NnNvdowR+mHjOHLug1CIRp5fDDSAkDDVkJUsR/F2ifSSYal4PWm4+x
FIahHcrnaK/RYX5GHUmCc52YHAhJ62RmPzADtd+jPHZ0mDlf3+PGencIGBojwrto
Edq0BUCgntdiNTrdoLf1NhrU8JxfX6fREz1AcFEAvOY2kcqtjQXdZud8N1HvZN0g
r6SGqmGksy0fUdnNqWYYgjSk0sAkvtqiXo5m+WzloXa1ap0EE4CZKL43Bj0QNkZh
m53ai8vsZxnnqK6aoeC8x/CNFCPySjYBROY+berXBtgSguo3rQUc5+g9nRYqxIug
xwBYrlbQhA1njiy/Z7zHLgeciICke7ZxDuAQQPCogMugYIRF5Nh45Y7LT1eHXxZV
i07rw/t9kRww/vN+pBNAOjUOhv02Y6/BbnQ/mepLlfbfjyIck5uSZFHDsoYkzE0S
+t7kfK4agCUnxous8bpUh4tpn3/7FqNYdGRwsWnCH3/LGSRYmUYgtCIiMlIEgVSw
RUKmdq0xDWJD572/EXVV2peukAhf8HVzqqyQle57lN51nKKUoB71Oo7+je16WD2/
xtHc04rplbdS9aGeIMsVI2ckXCo6DWlbL5OowN7yxqyMUanBcsjTaqVFf2Vx/2+4
VKDzoZGKJ0zAq6Eotz4suhi4ztaOV/YMt0K0MWnahJWMguRSSdjZhIcE/VniCPZs
nF3JiXFx99Mi0HKwmgvr4au2SROrqwtPGdQ2GRPbJlFMoRyXsva8rZRygaWe+k23
K+ZUtCll7aHxG3lVaw3XFHjCdgM2Pr+i68QCCkP4a4VdLbNBchII6AeKkC59xDwb
SqlT5ntmBEZFeqIPwKBIeawOItG5iCWXJUgCSTIeIQ9RFjY95L6CPjxkQQ7w8eOw
yvWfpX4ISBeE5ns//6dJd9K+8TFgpk3jWjrCFRkgb0Br0e1JI/vXVYpFwYFveeaI
EsJWZpj3rQahm7F4Jr9gIoUrsm6CZVQ2bsmcdE8L7bh9zQAHlW9cxEiZwdB2hfIk
Lqu5vmQ78Pf+XXAbODvJINI14vA9CStRnMQ4VmzvWQpKUFGJ0bqJtuQueXO6OoLc
oWpNBGCIEZEH3UUNWG1KXPYHFVmmZp4N8LJ63BViTKuLi0hhcjhAdSuqIUQ2wYCj
+ugRZx1++inFDeBK0xg89xSO8ckmM4cl+KfWBm6aGpYwfKBJrBWGur3YYH9HKYtI
wkT5s5Dn8fXaGZ4RJz3P+/49+WYpoiT3RkbpbHshYJZsc8DWyepAVdNYVFusV9fi
VPt4uA18QWSr1BPFUqSgVKo/jD7wLh9kUyRsDRIzRVF/ZkON6K2hgUH03qkVO6sz
eyspIYVFGDpxERF4juLmRF7rN0+ymLQywDOy0A6OXVCTWlWdb2GGl8DkrxlVWhuR
amnpQV3fdz41g+DNVk3Ws5bymIUqk+q3CzOAzxakvYgrDcZbIsXx6T7Gv7QUaP4q
9/kiBPNtleDcM84/j8WtAFsslhfgmdL0/41FR6I4uLR+qUzuOhfhDs91Lf7o7wOc
sXLhUtkqVPhAgYsiiRbmx5319la0vjb7FKIcmcrbnv9XoohP8mF8PolvjJEUVcAt
3j/D+pRyzOtjpazg/j9kxV/O2NORsoRkSI1s8Ourh6ndvktUouihxBKVbZ2AGe4+
EhVD0myh74Tu7I/GkSpgY2gEI7muBmUNYU3BiZ52nDVJ6b+YytBbs2dM+6AqRr8l
OK/gUTFu57lJcReTMtB1YlzQjz6rhrOuuQkBWaJWuUYll/Kndep0QFgn4jlqkS4Q
WcaLiC/1IT7xCjX/ROfN7JM/yReTppV4H853KBW/zh78cclSZjUjHXcRe3g2HEoF
jCUHWWaBKHp/mtdFhGzAahtGKYgJTG2AWsLFBGKcXJGB1nyBLscUTyLtAk1r14q8
eJJNpn6xLlzikAmCAsk24xLZDfngRpL98zx/lX7IercEECLt8kQvu9/+iOU7Z+Ep
TxfF1g6w084gUKr4U722M9tpZjAq/7CZwSt2KWDAqKUXG48ROJ9QmXr0qZ1oJuHH
QLJ8xs2VzEUjxY7/n4+lXLsd/m+UXxtMp/9Ft0l9A2/O6W6AjdRdo87iDIQNfHM/
MG4qSJC4bkD67JroDMc8Ru8oiHWBVW+gYP0Vyo+0HDv6x+goKfWhUbaPNauvc2YQ
so8z5+B9SpLIniZ0XLfVzkP1V9+t5p2BGZaf2xTLbZjNpggZ4weyqJ4MTF/4mhYg
gGDsyU+kulPFznDJ8qdsrt+nnbGoFgKVawn/oH/QXV0p33nWc5ov4YZcWGz0EQwU
EDfhX5NVEx+TFaN7WvaV+xIpB43JJkUo4fKk7kkU/vnqxK4+nIW7cmTSjPn2Anb4
fJnmb9RnPRa1/elBw8ZW5tlO44FTe8/+ryhjwsX3qh2xo4W625nu1Rg6GHjHFPCh
dlZ4yy7nGy0UELeYjZgeAj4COgbDuoj8Cj24+DIlVPWnxcncoXLRTV2tOTrTB4vQ
mB+kgGB2VulRJxBYJmJbHVD3syE5sEnFgA2fBEUI/J2BradGu6lRNsIOzKRV4URe
0qjETP51GDhY/V3NPvXsk7uFvTXQXfZmcl6yfJvDo8tLNYH66CL993L905LnfK0p
IL5VsYsDf/cKxvz/4L3JuJ6SqyHLJTxRnvqZFdgrK+y+kKNXH7YjigTPisIDGPlZ
xCVlXSqrdgMJWVAQ0uJeHD/H4t4Ymo9qArzjZO8WFNs3Chyfy8MTLhUIB4ybReMN
QXQVpKz7Ie6VRu+ca8fQ+KnSMzqlnuZ8p8P8dBEcTfo3klAXi3wNPTY5jGk/d5Nb
KdSSACnBKZ/bY8n/t1FwIf5aYGt9b90jjbS5yiceQP+mpAmxjZ6BX98/6cDHQcQj
lVzUIxkIT7726HyS5uzA1OTbzwzqA9Y4EPpcTYx/qwYs6xO4d0U7RancDobTF6bU
oev4L/SOc8ZcIc6/H84ej6pAdlANhevLS2sMqGUyn7n/099QTmEJNykCAYjptqcn
3KV9SgSaiEGFfKkpWwzZhlMT6Cnj1gxscWxkrkPWErBUP97LInwMeFjSUx7VcssG
0jrnOQU4eM0EaUk0eUqeeA+82+3vBj5/8Gp6D4hvRUCu2pyagZJzXI16IVUCV1ev
FxqZG/J6AFpQYPtpZ2XpQ8wD/2ykk+kKP/7n+UF/8++FLc8nDvTtKFsYo8aPyP4Y
vUnJ47frlDtHoELcd5B5CXhbjNNb/S4wOA6zsey1m0jk0FUjQHChMvbG+QyB5pVt
GT31mpCqP9kNpF6DzrGZIutw1FWmrMLD7fAYB67LR4CjFqI+dU375bfsXjbaDiUZ
7XewMlzXQVR/IUIjBYIvBLXOhmEAQGgvigLQvYKLwnAeop4iIp5ieC/EcFwHWTbH
Lvka/J9ith501OgO9i8u5buJTt3O7PG+E7qzawed8iOXgUZTAmWgF5vy5l7l8Ejz
2OCwBOEpF+fL/y+ig6FYk3dyQU4rlCNXr8r0DAQD2HpM9lmlxpSfHof3CEFQED+T
hef9wnW2x+oNGVIC8po/T4bfTU/SZtaJWIuu+npCh3f7GuRWUDYnZuNGGKCEAwBk
Fzan5AXvOwFVcI9muv518oeA750GVSFfmtCIXrLqMax6PI4yhMK+Owe4hM1bgQyR
HT2mdgO1Qw4K0oBxO0mJlnP6wAh5XqBU/puRtgqCK0L/DM6ExHOfQyaFNSuFI2/r
AoMnnBwIpndfFZKDoqLfAIfVG4a4DOIJZ2Xl2IW7iBRvI0JOlcpOPWgS8jN60tzt
tJl32Jup0k22PCn5y1ZVG08Kn7ArAokqj6/FY/WkL4lDWt3to2gEDRYTe0H7ozeG
907fD/XIPkTFrxtGN6OBelGTb0rzr7W0kiq4/NEs0o+j/qY04fdAS5+nENJttwX1
XqugbODjUy638XqBBi3AhdqxQfVaIw/dpH0bkk/ycGd88Mz/Dhe6Qp1+mHuXzK5W
fgVamZXdAwywJDMq7PjF2boJzk0VLtf02v5DjBWccWl2ab5gf0joKX7sTm8i/hIg
8KML77ofIZAOv8WUBzgLZB7tr9uZT2+oPNxh9ISQscvHLlsqJJQtLa/NTGT41pLv
cnnTygDPl78BspaDCWjPB1vPtOIx05K/J81weO9YMMYWpHWzQ6NDlS3GscJfc1UE
HHwlR68bYyuSQ8EOnkjvFZN0SOrYThw6kybfUNmlAi/SFjeOv4tXv0nZJ7rVceZy
I9xP9h7lRVdM5pJtcGb82r4JfTOJmRiDEZTH3hbgikMrQu7RitiGtS08hjCZATSu
eAI10Gg26632MFPAzR2I+7MT4VZ1Wybfd8Zex4LrzgbducT8VyolMlA7X2zrDYSf
FFW1d81h93xhLIf/fh1X4GBlbGN3jEJowgp0/zMJSP08VoTgH+WjJ3iR8mjqHULn
9/FXGjvtRhES71zirWWIqlOoHBWfZr3unICqdyoFgdyyVZyTl1FaJ4Nz9oiSxHVI
BHtMZC2MAVsS/Zy2WpSHVtnRAgf/QDgZZSkffMtyLkQC0pA4lstPMg/rZ/TT9sMj
P2BA6LH5Nsci/TmSMgUZiBRKSiexT7nlk83Nj/47VdAG19rhxu/Uisg8gvifQh+i
u0giqgndAxv91mD5B/9IapkakgMvLdTiNeybt80QwlY2OTCHqKQyiaxycVxxX9zp
RZ5c9jog5DGnwo04PnhppT8sDTI28OGGOTeLX2MZKHK/JPW6+JcCdlGRO7JfGXCP
IXx9k/LwwDvQtauljJGiLywo8EI9FPYrTCrneZfWj8nuo10lxMyEYW0wDIJTiqcH
nVGmuiCPI+HuaouPhAZxrT9QrvksSfPPHQj4sxVwL96VVS0Z4h2rk9Hy0924pj0/
SCUyPLZmvTvdI5p6QbesOnknsQeG8vJRkwMoIGHX2CFVyiiSmUfbdkI4sxlfHqUi
B1l78iifxnqUPtRwo6WSUdnephJeYWzJCZd+JloYcXhv11uhqcHX5Oe52TY1EdfM
VzJZWZ93cqkYKX5emhz1ffYKXTfWNnA9jnEekS8urvVJe2DoZlbCKi2bdqbQtjKM
MULRd1PNRXv4s8H0sP/03Hfpc+taU7GHx4zHWf8rLEF16S1WGorKOaAhDDl11BGG
nXXF/HRteUVnSQWWr+sWdsWhvk3mm9mVgRF8lgWT+6V0WpSLeEQxDVGeHFJuz0Hi
nk+8s5IcERw3RM/8GvW2ET/TjK7uy9C0RebC3+KlqXPWHoQGFu0gt078aBo5B4fR
HbWiubT+dfBeNw+Mj3qKjvVk78H/bD8rBF+0yBcUtf+KA1E83bznomnC6RteWV0P
ApPLrgXvrRp3fzhci8QWMZx7O+vuLUo/SiDLwvpxKCkMd67DIApCp/qAfzwQyk+E
CRRpXFzRj+Zn7ESM7ofGtoqzKCR3Wa/zCTwisnL7VpYRYIhHCu5ay3YXZLO3wO6f
u5r/FoYytLCoUhu7H7wXLV1oVrEm1L0oNM8jqhF7HGyN8aTL8+8xNJt93gAm7laD
m0lanpra3Xo+2we2gw25kRcG4RwAhPlhHBc+nuOrGAXqaCRKsl7mZhFTHOZwa3IW
K+bYScm4pp6/rCaoZ5wcZa632ujx6v21+pLcOjokxTk8vaLSPTYhl7FP4xfvdFb9
4GKGcb4vNafNS4xuO3TMqO5x/p7BrJzCDI9A4bv+SfohODy6TB5gC0JRAmOMYNZG
DYWl1fSJ9wSQUM3+R9RfMTIKsu94iSVZGUrFAgoQC1qSJPwsk4FcHuBdLXz0Stvf
VfVBaRfJKFXqrn1KMQdCMob4n+P1eqVWOJnOn5N4QesoBPLqCpK44uR6hZi9/wrJ
Y4gwY8qSqFFjRrxMtbYAuAdBSF6sFbkSNNquAzJAFwDupepUj1sboExlI8NSfJHp
QOSBZ/SvgvsmVR/cU370e6C2FgUm/aa2XOtVYZrtMkUijQi+qdcfcEhDlNAyN8Q1
xbhpLB2k5yhaPW1A+3/MrSPfK0n5i0Ir6ohhDfQ+Spm3+kczZpk0wm/Vk4mA1aD4
Fi5Vgj1mAx8dYMvz/cDDLUKPwNYJZ4WSEVOHmfcxHRQftphyYtOmQv0UkozVb++d
SL80NEacSQfJpfmZDuwf9vTwc3EhJDVyT9hpI2qhLmDkxVfw/20xAbLVPugkt07T
y1RiTBXNB1om29tszm/4YbiR/grqubAIz0mOOgxx45XiavQtnMCLco9+0QpSDjXq
mZDLhJJBLSWU0JELsslwc/V4D/WAPQkPPR1LfMnVehN50WetzztVj/H9loBhvst1
PsnGlGJbjg4ddtATlmkyQ6dXJ62Gj63gD3MRgGzl23es3Pocdhw5DSq0qF8U7hNI
h/VM3QKbgvRLFRpHmMnGrUw0lFY+Lc+tOsbkBZMW+IfeNUnGmnGzPX3H8sueDHUM
0u6mWfObi9IIw6wp10RDxr76LaIhuxrci12gHrJypuMreX/mCH+Rb9fR3ohG6w5+
jAQzMtqyYnOgs2fDcnizZHBdorJzYeuVOtPnVjbChVfDAsXIpMOWvSr3mKKEdv6i
G7sqHTCEVkOP9mC4PoAi1ZW9GeDwYvdGf1Stx3N1Yh06RrYw9dT/y3JKCO2H+3/l
VajI/lG6tWMRAmkQs02PE/hkc48WRAac0j6xs3D7gseT9qWoX3R5AMMKgTRzoemm
sbFKH3SeKPr4IHXxx8Ty63cc8p+0bCjPepQZ7aHsW/ncGAeG+hEvGfT8XyKH7S4E
VTPj3X8RsJRz5dGXR45YJ6HzRt/sbtSky/AcVPrIOwrc3o5yZssIqZxPDLHn3uV7
8zbk4iWvtOG46eXEa1FHN0kqy2fh3zCEfgCEdN2VEzbF8BNwlTsuGlrv76HYMSV4
EZzJZ43nxLGlINRurz1oEJxeCGhj+64skP6cimT7sn87INInr1xQcA64xUVkzzk4
2zh0uH2NELKg2llEWZyyzIwCXxyIQsgTr6JNcYO7y+Mv8nUbxBlpvbB3ziL3Ht8z
9vrFew2dmeEGGM1hUfcPSTQdD8yYDy2OkAvBxX63nCMqHnY8kFrHpRqwv7GLPRVh
2ymcKk/M+fUVBZrS0IV/bpQ6OiDMtpjiIbcsK90n0/RZV3GtUmfcA7utQ/FtikIX
tznRfbb0ZIIFSuw66arHDajtGOljs6tiHnGR4zEdtkmeMFPt0RbCA8kA2/5ynO02
+XUU9ENBvJ0FFKmHSvEQZIxdPyp4vSfff7jzS78bWS0UcSwqoMRYWVkY2bB96P/o
Aaqf27opVn+a6LhO6yjOMqg1c5GhK+6DJDwG3iMDW3lDqQGGHvNoVECwbezM0Ntj
3Sk5HfNltKHUtwSgNc52ZK+yHS4un5RS6YIWecr8hF3ETivYHEDvXKzCYOopTdHJ
dG48yrYzz46W7RFqP8LrRvScRxD6Tq2hOjuwPpD7C33gCV+bFGLoZ6GGNoxNH5u3
KjYWc09MRhIsIbgRrWx896qbS8RINuaehvIzxUUrMcmuwS51K6+Ig98OfKR+YCUM
sufkyxt3u2iBTJtwsmM4nng6lPtkFOVZu9n+sQO9pitTFbb6g+xEuqcaJ4zpNPCt
FroLZCiazTjpW2H4IZbkbXXcrVi1bqb7vspYFPir+vxzMrF/cQIvhY3Mc05L6pK8
I7Inv4xHBEvOusH+j0MpabZHlGn+C3rcp674kCmdb5mIhJ26FeUPSdo0uQHw5bO1
rw8Jv+gV57NmXPlGBYbtjpC9blN/ubTNsZHiPGl2lQStwWVZH182eCtmNiyAHFN8
AJIpUqe92MzdqDVcVIShmhB/jB1z9FhD2bEQFBUBZ9j3grb8xVtlGq2YZ98xGCvE
9AwdWXRlOJmevONjIUWtXqUGRO8VoYQL7ZS7HAAPphk+1r+QAUVDlal/IAmgSpkX
8xDuE7b68aBPorLrUkxY+Pi5yleqMpjRyFyqY/76IpF+q8J6eTQI9pUPOb56VCaQ
Cwsyym7rLTjmHSJmpYryE9WXYKZjzCTOSXs7mmc1OpODaHQIYkLZAbdWG8GWH+QV
vtvGznWdLcWu+7jsXZJlNCax0VaRrEd+jxP/Er7LW8bulidFnWF2Fjn6UEfQ7AjS
tZ1AbtrsJZ6TSNpVGUMnsZeLKoGe1GwowEQ9bX2Y+qeMSMVtdkXPk/A9lZoxjVng
IFLqWRtcDeOabz2T3/25cHXm/Il44iN5JQHLkTn1c/IYDLdNews68XX1pkAjNu4O
5IGXdRXvEz/CdP/8lwUCwANuytUCvpytQDasFBxMTBny6vwWd+Gp65YoJFnJg830
9LaYl25Ao5mWn0e3HAZUhJAj1fZ1nDh3WQi8FrEUpD4dXPMl4RPrWOUZwSl/M686
WRUvfnVpqCntjOxUmmSdVgkNKyiorQtjztb2lNrijcdarLKYDK1+YZNSWdAW1E1A
I2wMD87ivhxndCvHlsoJskMwHdPwX0DNUfmR1r+Qty3h+LWWoogeC03wtXfJil4l
Kay60FTISY1aqmR8BLsSpM97393Z5gSZbdj2D4vVE9CrCvIyz/G0rR09UBYSuEVn
omEGpB4efbg8rwefeksd5ZdFgg5i/KZjdPtInTIfrWSDa693usCQtW+di+5B5cjz
H5BJoHzsXt342hm9a161Pa06WyKOTmuIdOYMFQv/A12ZWEqTXtTsXhYLE3wqB7/i
GSN7ROyPDFArRH0oDnMn3DFpk7euH7Gs8GIImqjediT98Hj1Cm+67h+jKJBGhyUA
wpn6/g/ltQAYDIfq8AdJ8FhdN1NadmIgIaUQEzGnkF52NpHZc48kecx9/qrxVDHU
jd5CfKrHGobGpI7dGyxiQfOdz4tQsxKBb0emJh9jxb9Iw79CX9zdFf9792N4eXOM
E7JC6k2Al5zcMNXjYDmjK6I225DOS9ZXBcnx4Ou8gr9HtkSGo3zWB1iQj2LZsG4U
zeBqJksOG8gcDqpBDXLeB1FxQ6LzG7ZRsuiIYEuoYGyjzTOa3QC1apY4abO0bpWz
z15TMA+9hNVLW4kOsSlK5/tre5RyNDMB0YOuz4EBOGi+SmurXOmHuhTtQjy3Gdi4
Ll6glVja0MKZfcMbvrGJ9aKU1Qqt/5o56Wy/iz3IX9ove2Wol4Uz9Z6uUsBJhdwW
KTa5h9/mTkR7cPS6kgTDc5tD0PkqTBUjOtsraxzRyw1GelwX3l5L5ho0zc2I4tgd
LcYk6d48SyvJ5Ti8KVnXmOVvHAeZIruHFAKz6/1y1Qwb4eN/nSZBv7W+jmftCdG0
RtZMwNDFZHWC8fPDHolAs7lj8xOqMdgO+1T181p3wNMJQ36feQuo450Lr4cr1Iz/
4Xj48eGa3xkW6LKKC/QMU+li1Qx+jP3X3JROdvrm5Y79tZ0rp0qykO7fXQyV5hDo
wJPa3DyYLFDz55+Ce52LtLq6Yl9sO6/MIiPU5QkA1cXLlQXQkpDBsemtycOakRkQ
0GVzm3yeWD0rj9cz9y7syC+LQZakB3kOlpWQJdVReLoR6yuc4dreWcGzsjERAN/U
buxGTcTVyJI6tMbslV9H4dlQncYHAjBjY5zmQbi8WRPJP1zw2tiMpgOtTBZLbI6W
gk5wjW9rPqvag/0Z1AH7zJ3K1ptE/qoUtbt2d3Epo2l2qR6tM6WcNJsWX+tZnZ8i
xVqTmmglY6+4bYsP3Tjsc1X2TJcHegWqzuNoCAXfjA3yZ9rE1m/d6WO+ug8l0MOz
84AyC7phzeOPPhp0n4cTdhUM8RVIAUTCdlalC5J3XjAhoOuTN/m7Gf/3e5lfS/V0
kdLkFJzAI1WzMoWOxNT4hJFPfX3ywF7KNk16Gyhks+LIayc2q7PtLq98K01ISalK
deIFxOw2EMwwP7dmcWdAdeKHREt8QfW0S7pZ1shw93/RqvYKUP9lDT2MAtIVETIo
2vxhoY3xxve01N6CRNrsWGKkxfdypnDN4BgCUOl61munTSleO+o2EbpTN7HSXEHu
qQ/oPLLVtQg3Wn3xKlL6ScmRRfyOhjIeGMJSFNFDPYmcTc05NV1DwH5EhT/CBZEo
3Nq8AWVZmi+f/nVzaTbcVAtNFESKuTzgvIer5grBgtt6JJsfFWlifvGlUWLjgiSM
FkWkh2h1t0w9WKAZyUYTP4JLp3dSQQ+6/DJx3juwr0LMigGhkTu1+D9EX7mUO6rU
Ygon7LecRej/25SNiFK+5lKxQpTz4XwsyP9zioq+J68Q1jSRudA9mjLZoR3AchuU
Lp4c2mcRQK8mtdm7ldjQR8G+Ua1V6T8S0Mi+3ruYrDuveDjLaYkXMGZ5D5LJZkv1
uKmIxVxgPvBtUHueVOa1D4R15yeqMolBADndI8ZgXKT3WpX4eHjTLPLVuq1ip274
BTVY/7X3c3qvNv6DOnXqFoUP9GcrKHZ7uDwdPYdVylOJdopDluuOR+qiA5iF0UXo
L+xTvJtS0660fNqIG9CEngHCeRbhmYm3IJDLFlNZyB9vzjc9LKwqKti50pnBqaJS
Ej4Lm8M9G1uVtXrvqxz3+mgh7ua7/Cek69i1cQRjV3cw714LmLJzOTiW+IskFwML
D41aff+SIt8n7L48vmvHBV5XoT1EU+zQw+7TuSMsiny3W3e1FOuf73W2Hw9vR/X8
cCFxhqs46ckkV7usm3MfHc5z4SKGutYQt3xcs9Eg7IjcR/0O98zBz1dfP7CeISFm
0Lkf6OYMpGoBY4+3FTBIauEE+j2fcVXCd0IUKEXFhJ9RZ6vrLbrPe+edXuXvgS+f
Vok+mWq6JruKoMZly38IT5nckag4EzGtgTsavnk7X3efMWXTg+j+hPRiuJDMl4FN
8Zuau2psJamK4gyuHselnCdnB3aA38FVyVAfUKbGqLsaN3oYhUi7qkHSq9WK4zoU
G28S5rn5A6lb0iKfMRXHv2N2dVoHgG1/umW9K5ONkigVgS9+13RsiexprdvTM3st
UqU52SJRj0BGPECDYsS6VyaLYhwxWx/y7RYOFGrj8XRKNj7WJcIIU05uapRWzZgg
b4qLpgSLKY3L3IPn4vFZ9+IJkN0Zl1njWxomUY6WRT6FIonLbjhMpTLi0xAR48LE
hLVNZ67wTYpjfgsE6VsaeeXQoI2xU6QeLJ0SN1nzmCg2TnihXL53+mX6ItMG4t+k
UBCS3fJwpJ5NAsXQZkG0UXoxz5C02vWLpZJbtC70WQTdvNhY16Q9SG3mxvGFxQZ4
MOa7P4W8oUwQjG1rcZzsdEKQqF6/Ho9hGujNyhMSsSwXJBkD4xA8SxCc8tiNutGV
gZUaks6V+VAU+HjZpHhIy8fvoJ4/1QQIkPSeaA5lQxdaTTMb/ccN4bcu+Y2VT3Cz
bgdONVs15/G1d1mD/j5I96UF1ueAHlsnEjZbLP1mnJytLk0tkx5v4UCPeRanH1/n
cVtfFEY9lHRuvj87tdaQOHc2sBIrtcy4u4xevSwuolcjVCS57RksGssxg7VkpIsi
4qihKvjt1sC5Pod5+wevo0yoNZLvp2MxOAqoQYAJGXMLcvLuZcqsskfJI8/yilN2
ozwxxJEcJiqgs6r2KIZBOOU9zTIADNF+IplpzhDuQRgBAAWHuwA4jY6yk9qfjYeL
gmglh6962f6Dd8BOIDomVmscWoCZpdadDrI1D2i26f6bMvmZ6HsQ+EsuYkUD2F7/
jCicq+3Z8YPCylhfh+9CTvk2oIWNkGxxb4ACNj+ns+UaoeHMcyD39/UK+vQEqXes
Vuszd1DSLC7hDBGUiz1OlaBmE/9Bddxuhq8UvcvRRmXod1wRugprV5J9ay5/yws9
MAAJb2zPq3Iytk9Kxcy16LJvmtbzLn0op9oygXCh1mdSrQkOKcXnsKWNLc5G4qBm
TauolpK3zYaC9nfYuHD6Eze8yXF4OsCCnKpt1VaJKbIT2VG1BkbekEMxH+q/xQwl
sxnQ2/F6C6Po9PM8lt4pR+E7oDLREg6PeELKBTO1SYfPALqM9rtqM0cYM9oTaRnR
zWeAPtx9uBuvpANXGSrkeidA+ziSTKRZhuv37Fd3znQxcmY5TicY6vGHpiFn4EJX
wPEedMGDGQzg3TInM6RHjnWfJ7jZU3NWyC3Th18J/O9xjG3DKWzTyaPhq/f8XhJ2
+SVnMPl2tZlG5j1RJ72YBht87yqAkZedLa4EXP7Qzbbs+fyTYI79B9aYjv6bqgg5
i8Gih/UL5aqFnYhu9y0IllyOJf3A5+Tx4tfS58SAdnZryiuXVBplLhsoIZupFfj/
h0Y8u/aMVlqt/I01gJ0nrr7YlHVf+nsnDy+I7quCe1VJZeMoxFVPHhbdyzZbh/eF
Zi7I3+9EnyBDOAVJfO7juF6rkSJQw+cTd8/GrOCXn5GVKXQ83y6WEeMqY+8U7+1D
FA1Vp8iVNiOnIAKJ9QXieZFuJsYrG7L4U/NOi6PddZn85bsRPOl56r1I8LgO/p1l
DIUq4OBoHsNG+T1gysYbfhPun9eJgyVVS9Vu2FSartDYG7m5NDKzk74ypWmftO7d
+GzerK710uN51AbfuqEuCQZBdJifzuOskMD9Yy7ZJIcMHO3iQTC/Fw6/Pl3m2KzF
I7QSw3eFfSxHwFo1xf6JJJgQI5WqPPPMUxxzE1WokHXTnCvdT+eOai4qJnFVURUe
nxH+vG5VWHk+P+Nq+HEOs5K4Giyt+Pqn0x+8ZVnH75lZvnydWzpmC13TznCYb8ds
scOSv7+ky91QZ4n7gV2BHRwPY+wJ8k77yI6H9gwCPKskjj6aJxdb462b43gxvUNE
T22tdyWWIsT3nxNUMuR0B2aYL7F6gz6/oIHb6YdWtFri6gqPzITjhCUkjl6trRm+
GFKaT5aDPVXjSntByXFsF5IqlMR2ZYHzAtnK56ENG705ftWSzKnQasBc+rptLoO0
IriIp18oFscUmk8/folbBgRyXDBdc1AK5cJOBK2VlTEQbQBXWoaDjpL+u1rUj0aB
H88aQ5kvgvM/4+UWrKCQKnNca5JGRQ4FBL5GD5BcCgcKIwSNPiP1L/n5O1iQtGF8
YSUGgPwZflXMFSV1gqUBrXuMRydkvZf9H90LeBpEZ7hj3TRLzebxZEboGgsmcrh4
IdeRHuAdoDk19rBHX33oYIgRknsffLciv1zcnpTog859yj0DoCeefdM8yKrioVNZ
jsR8PpO1+XQo2GZ8WyEG6PVUh5qL2TGukgq2K5/jEqH9ELQuWw++QP7zBu84IO/5
ThEVp+C/1cFQ3mf1dhunUZGXhQ6KRN6CrJwJ2cUXvkD8BEwENcox4GgJ7SumlifS
qMAkCpiEs3DVWxDjcBI8IIoXYZAHAeGNTrviIwkAAZvGxhlS4D5S1qmSS+iwMwnT
XTQZ2dzZ9gbElWJYf8qgnNpg4Wzwp89fawRZN80+SczTdhXF8RHv8eO5ppa1ryA7
vWZTfPR9IbL0fNNWyVUGyJNmf9hauV305ONpOAktpmy3NnukfawaHN67zkp9LVAw
PraQ9P+pbM8Czr8KQqTBLKBusJBkur1spuZhbYnGsSNqHnmdO7WlVf+poO+F43sI
0JUIszjs0JeLh4Dhcov/22lFMtIAkUaHLuPggVt/Vj8BGZ03+bohQev9aogSx6UA
04ksd7/gjuZ+21WmdnKbE+Qbq2OOiawKVF9/b1x/U3NHlPQO1pF6zWSu25+3VmVf
tRJJXL7FOtlDHU6NlXieODuWPVL0EyJJWpeArgDrqcnEEgF4N/iJw9JNL/P3LZdk
lPU09Phsz3+JzbBTvLZTsg+xi87fBth+jWIkyo91V5zTHDz/lQ5rDNZ7BAAm2RtO
gHtiMfQaDh5QmeQlboXyEF+0GjsPOm4uTayBwCa3OO89lD3M/KhclEbje1p/Xd+/
oBTo3UXhfiPsAGaOCQWg+inep7kSj2YL0QdilwWddTwpv/2D3nMfVmsUpmmZnxN/
/puOG+NoAfhZ2RLRf+wrR9vWr0VRBHGB+exwXjSrPZQxNezQ+hxnTQghVmzTYYng
Uje+DnCu7+aNGSJdHK8EKJ0sFVD0tw6Yc69/61Ay0dAPV8+gBL2AL8iMxoyI4Hth
ae6LKhXFtgFbF9WyZHNFQletMqpuSjDxr4WG1LPWIAFH3x4k6H+n6p1pK+IPuYVf
ruzJH7LkxJRHaudXTm8VQYRnU4pnkG6sk7ikSwmJqQkYw6e/2Hgyl+mX0jIT/yQt
+8KVzVXmD7PPmOGM83OLsxkE1BDW1pQbNFazU8gU/db1pawaC86LqOMEHjpQ2sVU
wvm5TEDy2PXCp5IRdy+mjO7TcEeVQD5FvlpbdlDHUZ/TiSsEXyUqrcxztuFRc2w0
yd8MyaXlFJD8ybRGiCF08yPKPznhebGcaxH4vYC54Zz9B66Ga9BWrNyD2u/sd5bQ
ocJw3YFeD/hjKUDi4MRdzqBZD0fjVRroO/8HshSPHdqhm8fsBbVyEnloBYp1xGQi
X88dGtQuTVaT2xSY09FLZqjdXLFaZ78MiWUF6oIt9JOX8lhMw42TJOPoBvzQL2dg
leZez3pr/HrPNRuEfv/XKBcLZdoXCp0vL0xJ9sTS8VNmeLRUBD5DM8L5eDJgU436
im0n3YuOZtSjWv6j0ZLHqm/daMWZYIZcZrXBRgT6TJsXTOabTFx06ICRMp40JWzj
RxmAyFZl9cKexYsouU+b77OXkzoNJbjS/pYS5mQgSq3UfYRr/uNI+ngKyYbw4VCq
4aBveKcwU3yRWYkhzzxVkZqWdK37KI39Thy2ItiObNm4c4GjQOdtNKHdA9LyB8U2
IdemJf5VWdIENLL+0t3Pd1IFCDc6eNdr6H3yLj9p9fqXVctfvSwRnFTB9zT+5VKV
SoWtmArt9zLKPmEIHGlaDaFls804n2QCe8hrROzcOlbAsUxb61EwJfDcZbHHeNZC
rkmMazB+hHncA2zpgwPfanV9eBmwBUk3tADh/9/NZxTX8WfUUM/HS8WriE+fs5mP
eKvExWKQI7UON2qr0zSkBNNRU+q45HBhcOeyk1KcvBUKjAuJ/Vw+8xuRZo/WW7RI
vrM6+v4RHkOwYiGUdh8Y2soX1LVBD8kKUgvpMZ9z5nCxCYWk9bjlJAfLKOS9+F1G
xjQ0OXEldyDMi8/C2nKdbnvYXZGOsMqWRVqkp35bvSS4NRm7SLXxlFcIFcgTCO7R
j9okGu0iqOwM6CCqphc6eJOwZeE/BQ5KbTlIwGiWxtYrij9+XNkIyGRQM5lwIq2e
PMYEcgTdX++4cTusrnedAn4wV+u0rEr1+ZeZv243HubxekH1C1y34eC04tmn5C0Q
doqvvkR5GByAjBlJ584tayoREQ0Ib6OfAhil1Tiuvq+l/Ta8Q8x8riD+cY8eBLX8
XWZo0fOy31g+GJoSh0YUId4F8FFC8NRb2BE7g8dVvtBcT8B5d5d7luLslQFK/hRT
o39wrK/Ex+6QmZxavOjJgB2hKNl8djx818RCZLMxm/7MOn5Hx6GxPfYQVrJO5z2l
Tt2A9L5KGBtf9JqeDi6nhfVgAeSPpkyrhHSRkVPn4VniDhGJL9dOpBBsG9EkNmM1
TnJVFy4tGcaP5hVY/sdhTNV11lzZ/GOeF4JxHbpA2Tp5VC6rcPdDiCOlmJCflmcZ
p0MPD1JFsX90ALyycMg1Q2YFZzMNTImEP/pNggLqgwAMr/4QuUTCgsO5vUFIe8tQ
vAWRHyWCui9cDkuiCz3bqSV6YtnFu94z7Qz5cItOdLWTT67RThRzSttYdj5kbaVn
m3YPnTeRF8Moa54dzaWbiLLRWx0/QFHIzroGF2NMnBxSFhQVKLPSLlSqSI8d4zNV
5blgg0ZWR/xrGp9r3vrKZRiI7Ks6kbPG5/GSFmFm6aWbA/sHPGQogI49+pKwQ0Ar
dU/msg6xA20gV3cJIpGKBTI72uaVzSskf1EnLQ1hxxLgIvKlACUOC92KIGnd+/xE
PIpCkGsr+zTCfrBUjS/td7loVNOxmD4uweXAotyCN0BUN96tK5BMdsbvf+UHrLWR
e2nmbYb2tb4//dVhIZdBwmPMjU6g/ClSMMR96OjvTC6jwioMCUykZEtNdVQWvxQh
sCVK7juwBRZQsJyZAjj7iQL5jEBEEEjk5ANavqLG1C0pGcSfh5a03Gq0lcJwigpE
O44v7i/JcWOO/WR7bJiOP79OlcTdYaJGvXAhDRSlZezgAgpl4nSK2+r2MqZlihCT
l/paFoyNJuEIvoSANlTg6OECTcefcoEHkIy+YTnGXUcVqXdHUfK1GIDvJEoK8EfN
XUc8PLXNrb6extpyqhoYfBoK3KkZ9jBrm7UgYESwJNezNOYhXRJFQLGk1oIuefxU
UyoDutcin3NPRZ3yMFAJLL2hX4wFXRadR+TX4v/zkA7a9j5VpPUJ4390gNC1CMiC
Q8l+rY2HrcODZRAQBu1rgpnOd29Sb/nE/tP/bT+GPUyPw1jqQ/DbYR34E5bU7sLC
/QG4eT2fJlFAoNjiMnbQu1hROtUCkxNvEKnLPGaAs9/p7cYdvmTVZN1CrA9eLxem
GthwRHEEQExZUYP307gdyFMIb8cKvKjt7nVsw63SznTuJsSSvxokat9vbTmRTAKG
WRSMceW/+B3KQxLgizLHIFthSBajpANJ6I+vvQjgycBMGhmPLF93M2aaAr1ly5KQ
nIpLSv0k3H5GVgu2F1MQwg3x/QoXhMMOSRKGPRhTwVaPRig8UrsaPCDxvSqYs8iO
X7Jjfu+RU6qSuYTSBpe9knX0Os83oaW/Z+MD6o610VB+KdTSh86OrtV5tzY5XBzK
ZcFpGUAE57hF1DmOrVTURI/hBO9/6CzoHz9LP2SjjXEYHxQI2IVpUG4pGrSgd4gZ
QnhfCfPgQBQwqFXuJtUeHrINnB++0+EjB4ObFuxCeaxSswUasUY/nSWm8FlCZuQZ
79iRzDjmXOltSWWmJHfpMwQtqBbBYzoaYLKLP1RwUjh82ODhwbdt2U864VODaYjX
uOx8kL15UOxlljo+LgafyhBiK6HCWFLLcUdTOBgA4SEwhduN5dYf1rrZMF+7e5kY
3a3f0DIHYZ2hm5ZO6Hs3KKfBrE6urU7ICR0NG5hI8VVcv2dWDgomRthluh7+mmCK
/+DoMQU3qk73z7kKCkslFsIQpTamZFvTTSRDQ2MiutfENKVheENGPeHAfQUplWWN
4g6e2kjVQvRTluhtuLhwgf2uRQgV/N8j1tx6B3Iha+AYHkkTWohVO1+eHVgz7MoN
PJuoksOrsPutwKSG5GcJNTsgmxUeO0Fp4eea+Ij/giyrw23rksWZqOz6xgq9aBiI
4f0ani098gqGbPPTAOzndWLpi+aw97EWTZWtnW1rfRH/mYzsD54iabFKhFxmgq6a
6oA8LUW51MAxDvtKtPA/7hKOVj7AK0RS1wtUt0f87j2eCcUjHYe+Oh3NcLfXGpFP
wKZ5BaWMU5dLx3VyYWjgNDvN6nD/LF1Qb1b20iQYxIqucmuhBz2d7lTvmzjyvY+D
t9ERLQujWT1uHWnXKU3FGpmya1T6d/b1sLCLUYvUBBuw31nBES8/nbotXY8t77xK
ElvfHYRnd4KwRkYHxUtEI/N21icCuemlpNcxfjhsEL2FPN6W87NJO0kNvMD3OO/j
kFPxVbdkViQ/GpFy8yQi4DnvdOcdcTCO7xWGwn/qBS4aMkYsjgnNNkH1t4xy/ll1
gZLZjxvy0dDKWBXmNDa+Yts5pPlsNZfdahLjLPnQwpGVZEg0u/eI9aUbfjXhrAiP
pDA71K+Eyl+aeEfE5kTyHW2q2hUYJ+B7/tgcBjRKGRGepvGRb9sFB7rffxTsuI5Q
Kx8qes44jGwLzZktXSQMXxPs9fsCG/Y/0pA9p6T1mewirfFMPIAL1ib9hh/q2lKZ
FQK0F5p0wOvHVd+Oq8YD8A2BJvQOl/+blzghneKxVwVKYE/j87TA9CNxcopowwdA
dNfrgTVTxJANeidFzXJazTCYLs7+7PeFEzctK+Q/xQBD0VhsF00sOkXiuVsgFfwy
cJQuh6CLTweFRLMovSoz4zVHfoC5tzF5M8yIAu4AzaepU3j8SdFq/WvxUUvWSVBV
9hd8ZB9pTwm+WATP/gL9CyzR9J0nAUXRK/cH4rTw5+HGq8uzSdPq0iuJuwY7R2DJ
55JDKN05oTS1dvt6BTFX/fx4ZtfQfrm1Bhymk+g3XP1sN4+e/LAdFHybabmgXxam
5CZVpj2aak4cFydqt4ulXAoF18nYP0sWi5iVq10xyy1Yu/Uczxhsz9MTeWYxxhLs
RwtTvyOeAJEsypVtMlG9VsB+p74dAu4EwzmjvyanpyNvsgBPrQ561YXes6hjkCEY
j0JVaY8CznNQfgF8FcO/BPJBiU1UU6P6AZQ/i8wSyhk4uf9avu+vzItihrk2/IZ9
wWVrZS7YL5z97ecsJpdIB6otv7/Op0urN5DRhA32PQEOEXgJ/168b4nqh0sSD1HX
jOqJ+n34Kmfi3CYbH2oFNkMXh0ogM21oHf09TQuCfXAd/MveTQy8p2FnhCha4Meh
0wdjP29VZuX8oBnkUSVXHHYj4dCVdpPtcqXo2e9oAX9htttkhGftLgnJvzPi32gv
nQK7nKJqONAtJJi6GBdJ8Nb/v0/GIgCVHTinf+t+7DUS1jq1ZYZxRZqj8odTVAzP
pXEDQOv07BdwS89HczEB0ytCHFziVXW+sC081bT86Wp/USA9fCJpBSH5+Ia9WMh/
E2P2EdTm2brK10vFXVkMUZFJNDtXsC7FN/vLC/6WjW56iyxnrAmSraUi8dT2lgRM
ohHTaRTOLzWKgb9os+ABb0mRPgq/4ZfNA+tmoc2ait17s2dtpgvnp+mkRMVY8/UR
H/Ss4dB6v/1M0Lh2mwawXmvOD1kqOEFxKsoO6P11gwExROpqb//lQSI7uEE8jvTm
z3cfA0s5nHySB3/CbbVcDTemiG8weCm8s7RqPL0S1TgvIq2vMwTnc3A4MPkPXgoM
oJUhkaglZ0BXL4wZhaoWpww84qwbBMdI1W8mEHHzH/7z7i0F48vadDRkuT/xVPxS
WDowuSEjZDDwwrHeNDVDYQGrK8QzJavVm9ZdRkfU2rTJ0gBjmB/U+xevRkIWgsWY
mYiOCcjBDLcFryk7AstCRlw2HdgkxnxpSehP6Cgahkoy/c/SVW1smyKi+XOhW+D8
HuXMOJTqJ4FUnX9vYV746vKXPrPuHetCrDYgBdATb/owHcbUo8Sfq9BU6poCtpUE
PsuTe2rz92Wb+1yzDZUgS1os/rwwxKZXtcxMjCTAMMSrWhhnowv3w0tfYhfkPr5u
NC2YmQuCGIvK7p0Wf5G5jZHAdQtD+RRWfd/Vri0DJhJ+8LBCvOXOQjyrWNkqx72V
lLVlSh47ch5LtpYEnvsIBWB2W3v7mTgzZ0KjjXF0qSYbd3xN1K0NSO6CscYo4ozB
ZkzHC+8V1P52eb0pp+F7zoTOBeX9NCGpXlhLe2SXeGWoTeevJO40m0AO+hn96Npf
BRldfTHP9XMzSYwMMBs243FDPtsMEJFXwkwN5b8n6rZcJUL6A1ezgV/+WK3SXSy2
Atd+imaLS3WJOI8MJKEJ9FlQRu2Fi9DGhpRMrodFuHmNKjQqk3kit5hxyLqGtiJt
LtjTsaLxa+izWvghOW+3ZilZYIthDeQjlU4hyR3EnQ313rscN6hySRpQ0ppvALlC
NDNMXPxNeOu/TmiEejDnsOdBdPw71kQG+l9CjuUoTiNegzb8VEAPQ7joHO6Kp4PY
kxdqm0QSNe78EQgFXm+SX5ApnSC7mJsxAKq7mryHBT4uIHipapMQ1OGTcdMcQIy9
FjND5Z3vkbyB0Ihu+OCFL63ctUp8larFD6itOmzmG2kKNyHtR3NUdRtwZlAKjzhB
VxCLHLcBgVEERO000zM0Xvo653yq87vU5XpdRtW2+0EUOc+sXvHRj8B+HyyjV+lH
XSn/3GNFKZfThzss2PZaRgdfHEn8fukW/bZ2YyTzaPlJu67xExBWTTuzcwifymii
dOUMhwD0oobfuFYMlawdpbraUc1wKhwQ7dWaZrIoHhj6YNGDU1WBJA9UDZBnTfF5
urvUkWPHjP34rw4eClF51apxck1BhTrUT9W6pT35EsAql1Ldcvk5edHBQRzTSLTD
D/s9tEWej3WhFBhdcBGvV0hl5zbT0H7y8b7MjgWNJBChHw4UbJWcYvf4pZdVhorL
6d8KaOlOBTXqTimaNtA3G4dV4uEbkvmlnePundpfHdcdmJ9KJ1AL14jggSP/tRGz
VX6gnW2t09Q0Q0TnrOwxiwDGL78MZYFZSQqMWvRlcTQPOHLYQiw9iFe9lH9iCiAK
X0le6BK20UJGJ436yXtwQCoB4hALx0n5O52f7+gNizXGuE2waa+yIUiz+bjvy3IZ
4UgGwEeSab/jYnvHJEfOoay8QxWmUT2ia9svCpqQMtZ48H6BPdz1m2lVpu0kHqcz
os2sTe0GjyTDXs3IfdoH10AzygH/ZyvX38zuVshl+vZshTHbYy244dgStTRG7lKJ
O6lfsHkaeyPRaVqPQ0kMcf+dfDBolpgZiaO3l7Gjy/Ufg5V7DSvjfC3E34a5syPh
PwRKOroz2C6wTytxoVdIuVNtVDlI7XvmyZGCaLJLoH29Rqk4ARUm9V/jp6Av5XqE
Ag6Izn6oL6eTgpkuoT8eSvj29xDuo6nPclK37JV2FT7yb8s89OMdeNODpyNp+e+f
IhVr5txSeQr/DEDqQYGHCeWiOhcU+2+s3bEGU/gSOyp972QDwbxyZp4CJ4YNp3HR
KXi2WOp5PM1d2TGXa8K254A4Bt5gQhu25FjKrjYNZk5RgcTXZf0rM7GTcKMiYwns
h1HKzWTZjv+sc7QNyhMLEC2LuB1NgtVLNAwLgSdIhaTAYFzh6EzCmd3w4mKE5zIH
fxK52ZMXxIcs16x5/v8OPky1OKQsfR5W97rMPYIJKNNA70i0lUiROz2C9uj/PGjm
I+QVDItwcEY9pRIXojTpP0N8Ux2spshk+P3pz7gkc1IbCfLHbdmBsuEIMxIRBnYG
oCjaWAo6SPiGskGxNl+gPVB7q2eKRdA/41GfLBpHkNBHsn2xGaNjBO5C0vZphQFi
cXWjwy3icel97MsPWVFPdAgNUoLuttFHVG/yzfg9UTe8zwG0rv4vVxjcpsTc/Mec
+DugKxKM4IIhRlWcFYADS2EpYXuyKKOsTB9Pvv6aH+BX9euBbCLlsnAH2IILAE80
4No8yPJWurYo+kI4/b2QS+btHEW+KU60ML4f6p+VaV9BA7o6xHJ6W7h0cjv9SikP
tdXjFPiQe4QvMrLsBw8iVCDIhsQkbvJ3bnSswd63IzA7NoVzUoJKSwxqhSWLpS3o
vGqMlYk7pxR/UXqwZVh9XBqfVOPX9dtrf9xag7DO53eoh4w0Veygrpqi82z/3J4h
+dkoD9KAwOTNKS5tpMK57uVndSQYxaAPUoqXWWNvBsDAsuxUFG7O9G4XqKWbZYNK
YUD/o5wGXXFB3adsjlevlv9vT8AxR8X5+kYjJO9K6fIOpXYhErR9nGXZZBdNIMQN
UptwCC/JMvdJmEQdvymLIUakoC7aHy+4j4KB9vDyyraLBexEc1H8v7taovbrpmXZ
524ywtc/SkXbH9O8OnaFLH65QxwxCDjUSMSZNb1nHHumqyf/cZclXkSjB1AUs5h8
IB2WETWuONMO2aNGhPBuxtcNKarxmAW19a+pUq4vztOC3983UI70BSS1yHY6Q57z
1/uPGtS+LPWgEMZwotQ5Djq6+UjA8amVZ+coMrO1Zj3YygMRWFdizLpA27Ivt4mm
6CPAMekp6SDn4ygwAVPENs2g9iFFEaGl5ccdal/1AVZBwyUfXNe9Xn4l8Yd/CLEb
SmooZzQ36MqrbV8F6pYYejFHobzyles9qRHu/fUcEDsYMiiP6qJpj/HGXhHSfRiM
4KxIsuN/N1qrRbEVkfmbeGX9HnO3aGa5aKOU5WYzAkLTunFtM5gp9+KQ+XyK7mJo
g4mFy8ZInJD9EzhozsUhrw8LxSol89Wz405lR7/nN8DhZv8vkodOh+zqBEWqUUD3
NPIYF58s04K1OaftsMnhZ9MFdsxkVJ7u9uC4h/kajyqm3UryCwb/BH3bRGQQ/9bI
t+mS+f0Di5KG0N6F3gCrmmmj5YoJnxpquJpdfSoJ6jIAafI92H8Lx9ncIIOc8/Rz
qBxubfN2rFyagv5cDQuuOzHlI0t9luBFm8DRA1TXHJXgOvVBuCHOahQfcLLQNJNK
kvTZjMK3g+JFjdwdSTq9QCCqKMYliV0mhGsBou8C2s85T4w8PBohqB8H0AjmC0ez
1xkgAfXso36nd8WWmvGlPyCzyIBked1Az1Kc1kIdUrXlbJQ0Ari9DrPreGebu7Ku
NoYVfDTZOrwwytd8XfwT3qqeX6Q2SrLR6IqenzQffSBdM2w3dTmSA+wHdTFVGmVk
mQ4bDkx5vypLfdIeybGL2v6CDFz/o9hp3mumANK15aqpO1nnYFNxp9AQLzRLWTCO
cwh8SiZlPrbauMAPGvCz2QYX16TSO8ub+4i/AjEqgV/gHeOj4NpYVd2e8UlMXZ+/
tNVzbw6FwywMqJNubM/hzDUA6ERBKCwRIxDL/mn3aus4EEp+LvvVj9oOHD/OBLa0
MqzUAoQ3X80qC+hynVFLuwwBzhVTzCmOBzXOt1E3ONFw64heTDYaMqw4u5RVZ9P2
w6PoOjz8fECHs2OgagSL9S7f8a+rz1dFDte7K6MbkrcZiQUSoldzi4PMyrsVw1qW
GBQoGHKsvXAbpqYQaxzDkxQjOPse3K+Fbsq/dZFI0urTN8gcYs/8bdU0cjvloEo8
QD+WbIq8HHmJX8lE0ZmKW/ZK3CU4qE75w5QVExBZ7N02uznaD7CkiqwGUZW7et36
w4lqQFM19cl/M7dyMrrRvbEp4S7JJE/Fe56AFsKRN6Z+/r/+E4WMK6HnwVupKAoo
pl4ZHnQwZ6gzuqazWRuOIpzT+fGeIQ4I+8QW1KRKjnnLHTDTDTiMBcNpv8pao4TK
u8PlZMfjnD8tcnBHlNHrSWUFp7dCIS3aJ+1/vPFOy9PxBMEPgYuUskM6gKhpnhcj
3vDNCRsEc/8+KoTj9Z8/IwhmETMBU50U0K+HqbK0furCdFvGQ0AXxLDUScl+z9bM
yuB0e/a9l0wrJBDv1iHHp/NB7+Gb9V67yySEsnDkh/T+rzqiI7tOLM6VHfsFjFdv
hDX/WdlMdnZoYBxciqRnjf7xRhf5VKZP+0q/BxOgZP5F+ZJWqD41ZOLL+ACsvQul
e95Eny3EZ+7et7AXMsQGgUcydUKAP3/arxl2b47/aVwxw6Zj+Tfj38WATsfKyMsT
UsCTtf2B7Kir3dNf1aj7EDt78pFrlWAgU2YytuvAhpBQN8C1xMftDhxwmQ0iwtcB
kUAGLQ32M/06jKqFP/PHCNqcS6udMZbumnZytw/YAUtDz4hr0Dp9rR/JQbJ/TPwh
Ij45SMPgpZj8slsEKVmhlaF0H41EQXZ2errIfw+gU9OLYBMw0HaEGelhyE6cwIB9
zBQC9m+bR37S/XACfLeR2Ol+J9KaEZGpVaI142empvbev3F7TDIQ+YLD1r1fCpSo
rGUoHibNL/Ncf+drYaQbZ3zzSvMIGDu/gprlhZrt4e1fBhpbMlEWRwywmyoBb3u5
sJTWqqMx0gcmnF7dmTA6HL8tldkM7wYEripsU4dEfFUCQC4W4vj1cpkHJ3u3tNkJ
4E7Tc9gPTmN2MHnQwbKq28ycpwspYzXV/EH8PIbFsyiMiWwHUbJee04NOgMGGbaJ
9kd6bM9Hln44UEFGocM4zmxVaRp2cWfdtY5pBXiwKy+R3zLkrjW4n751W2gKntuc
/hNLooUv9qnSB9n1Kgv9zfrL0RjmoThlKjjemClIqHb4WcsqfqP88GYhFVGvr4Qs
auCuJ3lJLDtqhuUqZZcZl7H+hGZUHhcYkUPaEATnIMk4VU3a8krsQcJo5op/bPKJ
qNKlH3rZlWQ94RQl460H2Bc3FITptqphQTqMJWgA7VKvA0WfOcsoxpiklP5BrLSw
soF2+a8Yky+sHdIeF8k/Kkq6C0yZl3wbyZ48gIudlvEOEEKV0aiNLA5Y3eks+kPD
uRDdSHaKGEYg5pXGEzf7p08U7/5wdOou27hzJ3xRLTH3nqiv4a9em5oaIbk3+ZJl
APlIWHg87jW6QbuVNL21vy+0KprfNNP3VRno1IYJblVmBCi5RuSb3QRSNhHPuvIZ
MN11rES2LZdnu1T4JyUDe5zJ3geUUug6kCa26l0WUEe9F+MLfWQ7ARPM9Li7E2tn
2dOMmZRi9oC8keU4dKgLWs/4e4fW8onElUrOsxO6awYRABmjGKxgozSLtrUlrM2h
TyFj9X92swaYPo7xph0gMxw7MXiVuEUAh4qFeN1y5rJDH+wQNtFNSfXctWRo1Wz+
+pwxpYggm4bWifiMTQTxx0nq34fLV1Wz1kBLVArV0A7+BTwyzELdF2BdTYN5g2Fv
TWapuQ3b98JLjpv9a96Z7u4TJQlz4LihSbhJMfj6hX+VI7A6pdONixIeDFLnu0zM
RTzrmczwEE5vMG8DCBl0mdO2b1p0UfyYvc5zknr0q26WcFD6o03qSleUZTNuLcfs
s4rsGENaUAO2Ljo0enCtDAlg76DsexmxI4eTqhwf7xNAXoTDOr2+QViitFCWOjda
kF7KQvFicjhbBHlpg36NWQCvXg9g2U7g+b2aLscyLfqYjTlIDkZ5xZf9isANLiUF
YBYQRNmrPy6XEgBhU7OJVPU5GcHpuiSP+sbSjivdUN2Hd5aLFEGfB0794a6BBErt
w1Xyl0PnakJKJnCpb9iQ3tA63TYA/k8hFF1ZYsqNKTBwIw73n5ZkUIubZCK9FAU/
I+QYA6ODky/3h/yWpVSr0xGZU8yQ3M0BuhFWEuGQzeJOnN5qZRtkShQseLrLmLP9
D2vZkZrewFzpCRigWxFZJ4gxWjUFBSNVrpG6E+foLC6HvvkxcvzFr2oifbY4CHzv
9a1yzNqhRR2EkSrhof5q/JS4swDW2KxsPFpUEADPz2aOG07Q4Fy7ejbmcSzEbovo
2ffsAQi2B6FmQKUy3anjmLvuiEaOKoAaKKOXFAXZUihqRYls43kKazu1yAHwgn/s
QkXxYyKPjQAFVVp2E56tXmYUu5J6gEEvpRvfE5V0e+ky5HyZBMN+/bepg52FnMSD
n1w3LMCsS0BKmZW8Lcw4vTONBq+rPB08I4wwkXNkA0BvTCwVr7nfqRx4Gw/g28HM
5xXFHvoW1xgeziUwou9pJHqNiWE4rufbX3KASvayLQLgoiLdGWlHwl3Dh1Z+8z1q
V14j9w8Qc1BEMnbLFBFfffhVXxlRNmzqd6wryN3FJT248bmxoRItQ2ee6vYPntTN
Yid14t4t+o83CBnD34JUZ4UbD+fcia70i5Lnh21rQYDt2JmzkiR8m1klsl76TG5h
1NODQbK1NzCq1fTaBkrdiFpItqSTWEwu/VAd7Y2XX8xdu7+bW6sb3uXIg7caQAGc
HrzYkigCr+AYaO+5Iq5SugE/kFBPyFH0vvcdsgit4elJYi0Sg/+ExdrsvhQBFEqN
HHx0mynT7iNTYMvrwuCUwvKHnpNPYLchamsYAyBTPastE9aBSGwIS1SQsSi9Qa3G
4DyVRgFYOorRrtE23yG5f/K56hmiPm6Pr6vuVvHcSiCmUybvS2/37g7lKxdAI5Li
Ie6tZz/lXA4VLGzxPeet5Uwp6ALw+gosSvPTlk6il3mPLbGVKI4PoMgAB9sHGRDx
frgF5wxlVHeFdwU5ZCazLom0rpgUDTCnxHjbyZ58s601tXe0hafleUCBi3Kx5VC0
6MTMXfqHXiWz4XTDrH+SpeVFO3Qfe+zIM6DURGuqlYkuvGJeWnCwLKAmXprv32vU
k1YGO/BgJhRGy6L9Hajsxk2ze7cTu7Y+1Qfuk0UVsLNe4un50D2ZgUcJ6iG7wN3y
K1Joiz1XItz68u/cqY6cZDGwLGb9ytx7Dc4ZOtCgRxMiDiiBmoyI+vl6n9Ci3zsU
+ymKAFKK2S96tw09PPOd60msLGkgZrL2zFE3QZQTuj8YvDJ5MKJztMSp9DnmQGb6
RZ1rl6XwEXdV8ZfkDpwomUsViglbXq00mWFbA4S7LWuFQLHS7XmU17RZufZr0MzN
BpVz0YVaLx4aClshNWq0oKCstWNrH5Ii1yfLpRtVfB5UFypiK9kCY1VR0b39xyK5
zUsoryUGHpDH2S/H3ipVgE0msPyEWUWlop0PvUBz2itmHPK6zCHi1HlwMhU7y3Fb
emr2qNbXBVW0eW2yUu8VnkZhgpYrOJYLiq2fj2JRao+z6NLDHCLmcxMMK79zh2eX
P+KnCJuxAEDDII6pwqwFviOWtiqPyq6iWOn19OpsArD7OtImNWO2pSwbq+BsJNkm
emxK1/ggnVJ0t1aeZiTkru48JNfXAgkZBXoZJa3tP52hl7HFxGBDEVLxRKnHU5fE
lmz4qoX9t7f48YIQBfuLttJJDqCmho9riqRAFPO1FpyD8WNOfpyICjHwWygA5yMP
LXk90yRtFw9reZ5q1nzWzrNY5uXnEH1R3hsS70w2m/JyUym6QAE6FZzgJBZa+X8p
Srr9SIm73mXhkaqfT4hNKFvYxj2EEnq2gac1KVbOPmXlHx/zbH4JY9T6qooGUDtm
Il15ohxCHrXq2AwDEMBv5IIKoTS1wKd5hUoSlVBdpvIP2p33/ZL4/CN8kAQI3xhf
e1U9+ZkofVp8hWivKcLAy+5vBqBgetwsCppT1//cmUngC1va9q16NrOWoBpyk507
9zBK9okXwLT12Si1kMipDfnJOwERtnytxgnXw58+yzOe2b1epxI82XMiGMNVmabb
ftp4rNkPgGG7zMaN80Rkdulpt6Hb6mVGP3tAY4r7Jc3A+qF6Re7oKvbMWa3MVC3C
qtjGaMuySiXU7dHu5qa3duLu7wGSRKIWV2aE9MdIoHCUzQN0np1S3Z4ep0wJ3BLu
tbc/bw3hAblTICnrQkZWpIo+OSM9MNvvALcyF1AaVbEwkQupJRW1MjI0Stna8uB2
pDw5X0vLcpVakB4fooavDQQqdI4GTnmYaRsNoQvDyRA0jMmBKxpK11jrBTTInCtn
LVAEgiDFeCYO8j5I4rF3Yk4+79y97Bv8OqzX5NV+LtqAODEMyqwP94dS3HZo/cvo
S8thSH2UvAz40CJVdWZII+YlQQ12m0GlomkDRXlEzSs4Qu4AY1K8LlTu36ATmeTl
/V8YG6SN+8291ygCLu8IQrJmlHIG1bRMKO+KY3e3LulxpLe6/NnJZVVBrZ+aUq54
suFjFwckl70Knw7QbkI0TZ+wJ0iBgl9rcA0aJBghJcK8HPFtxtKWbyEbTKeI3q6C
sojjyIXKP1mwWL8x5fuMI/WaO7Eqadfc4X6lx86PFAzpta464TKV2vUxj47GOGyV
5aoOwurzH3cZsisVMp4nwNtMjQAkLDJKxJZaAxbPY6UhtMW9mo5IKi5svNmmxl6u
VeTZ7CcD6daXjCup63jz67IdGracVTihyMTMroT4c62X1lUwMrD7s+Q4fc+0yzWa
ewF8+pTyB1LTYxgnqmVK7EFVpL8lV/qta0T3IjGKMqADX0XofHH7K9hpZs8KSVB/
w9VoJDTq264TgiipHk2480UYKRSbC5cxVfvT8Xm2UiF4WT+X9dPNB7RQ61ehxJFD
XnA6oZujJ9GwMntcY0D8tLIOt9KFgP1rOS2rvxA5OLODjpoLZaCRyDJp3wl0SdfY
q6FvO2Bzcs022g9A9jz4HIIG2JvlmQq8H7ZKiYJCdTrvBKaXJs+n7f/RL5CkdV12
Zqh459Zz4sKXnfDRS6c1paNMBeXD6W3y8Zz7J8pZvGK36n+jM+Q6hAZzLkHa5CE5
LCRSg02VqeeIQmULTCWwunqvmYf6e0ULMR+Qlz5rC5Mn2zPHuiJW0tocFdYT5vfH
q2nSQZzz3ZSb2FLX/JPGIXFw6Yyu/pEZLxguigTYyKeRoRFqawrYkRt/disAxXlt
XvM6CNMSJwPVFPpa1nvNxbEHuAqlPLbhwM+XWtW28gYC27Zg6iUzFGJ1hsvlGUoz
8VelGywlutjsl9vMyO2/V6t7PpYTmvR3h/Ww/RZNFxG0/AWcb8CoUlyVbAMjJnIV
okppPnvBPZITQOouQXcv9eAZJU6Ry4APaT00KprVOCtGxPH8IhVjyMEtAMmSx6oe
A0XTYxr5pWMDM8sFvgF8/9R3kM8n4cJNc2NnwWiuwQ09sSrNvSVgptUXlwReG6gh
NmdU2BeegrYpWoKhYO+JEwQnuqsMLu/Gsf/Xy6Tr8yOt+BkNpIebGVkH3hybG4Yi
mIkC0l6J6gDJ4Mb7qrmZax4Z2asxnRPWeTi50UWFpzqNQV0XqFrAMzW/6K1BYjPK
qzi0OgjJVP3cF2xn1ja21iPPkejZAyI27KEXWqYu5goqbBHQyF3OOetlGG6NEWLH
ABcmnu2vIorwAwz9G0miAIttYQLSap/o2cVC8UEVOZkNLs4YcMF/dbjWNHKPIoHV
oumzT+x4CEchg2vEriTnIH5hohdyim9QbZfrgRbCbJE0HUKZ7Ma7JpADZQVpVI4t
a8pfvWqbKMMKrcOJiAWuy0zGdbhpdSHN4Q3MYJcNTvolYxvuTvNJfnSL4JKuIO1I
iDQhKN8AQPnrhWaVbTlJ7b6SuM62OHs+5pfQ9XUEi9eEBphwJc0FFM9gSvOH+TtW
kfq6jstZ7PcMPoVoIimGkdYCnWtencHujAJzl192pAg4XUsQr9QCpoq7kPc/MDFI
PjAsKkJmv/sAYea/TkSEQOIFsdRcpSRE/ERodVlPjutsuc1bxrwdA57KIWPaQtUL
LGDqMrOwROCgpO64JbzJmuQh+9OQ9+EM611mjw2XREo+UOHkqfLokCyS2/7b7gVt
mwYZfwLeKdjSXgqtlWtPl4tn0T1sfgsHBoavWuEazuHoFLr6rpi8tCeHjSSuExU7
DS1QhzuDaqOCu/mW0JxI2UOS2loaDZmucmX08rfDGCMMps2fdDOA+pYnMyh+/nZv
k0vplNENg26LtWi7Fo5fYccaHPo82ZszSgCWJcAiLVSYsh2ZD4va7lunknphWLiX
PA8+rIzFuozPdYvIzLtsPx+Jp/8LshMQdkI/q1SalxO0CyOLX0HFtRU2AAFW7jOM
5zbzwQu1qC57h3lmsofAt3on0Kgu0JFtyfEnWeRAoG8JS2TIk9G+9/YXmGQrpERn
nPAMIbXF2EB4p5N0n4MOw/AGIqAbwad/NszHjOjMQUo2X0XKS/afTd2Gja3CLPna
OnUrdhH3BIrlgdBIpRNS0lYhBG260wsYYKk+V3lBAMF6RtQ/b67hWbGpXiUuXWiL
2T//8Kj3MpIqEmdxcCjwihZG6VTb32I7ogyRPkDpWYAqIa3G8LYICmZ9kjNT1OHP
x6j8ageiVGevIcBkRbFRKtriIBV7IU/IUE6dtWfEyryzNTNHR1e00cRxoDuL9hND
qguBIraQv2Ssi2EFa2htHv50B3bT+gJq0VEduFqP6XlU52ksXioaLTcy0p6DFxtL
W30OsYw7UvkKAbYdA237p/XnJnuPtr/Ll8Pgd86HK+wXODn+IEstoj20+vGqDPuA
TNa8n/LGkes95wvUEkqP6dNtsHuDGo42Exa0qModNEs0waG009rMEI6rpvehq4WL
yKywseSjlG4Li+lTS8tB5W9XS3zDPywcjNFZ4McSbi+8HYzosMa+DlQCwF9sajoe
WNQBVDF7sLY+GeaSu/4o4YIfiypkS+3gbJbUVYd5lIRs/AcYUFruXhl4jpLWUN+b
n0TaVjqXguZBJRj61s/zJ5KOUoBLx8m6/FOG9Upjwy1fZGCwkqTyzSeB/9a0hD0N
MuO5UzZ9Jas4hqHnWGmOoh1D30erXv8Sv/vXkwe0iLX+jydIipl0OilA80CqeVBl
tUjaT3DQkxz/B7qyvxx7daMP9cwPoRXnlAe5tKNIZ9jEviE+EmTK4RUrXTdsl2Mk
kjJw/uVvJY1DUl6ZToaeupdePh76AwPVHnM6RzLhuQB6A+nVWbEqSslUD76H8mis
a2uJZvQxU11cuDkYpq7OPvcvu5LoCGEKjzsVQAWEvi4WOfEnyzQXjHDYkh2IdwJk
4LxWjLNyowFM9V+bcdruI4EVH6shZIafoEAvXMwm1shihWSThpzSoVZFlNdmtF5n
SVJbRkZlIS4HdPEo3QNcPRYuZF830g3+mLQeqcPZHpunY5ZN8F1txzIkf8vxmqMB
OXz+FJqjWRlc5YKorLDS/GOR1hUTpAzz44WRQI6svd9RWyRyoOU82Llbp9/ulD7j
rZAUeUR6x2UT7rk4kgoTFEq4KGfrwrgB8TQ8Y2ETEHpO6qH+xo0MmYhtZGKlLzbO
8NGNMNJltDKq1c9r/2kQmL0B/BohUs25qbqFLLyN15/JNxucPWNn2VWfn0v3A0rO
rk30RXCIylNlYUQwFI2jEyUK0gMrWn4gtjlxMG78A+0nAdtLCD4YJc4dU1agcF2b
6pr6kGXdCI5tU1ChmxLHBjv772Y3NFLNeCUZQj6qPSLDWwvs6ivzfO/dTZ6kQiBQ
csOm3WhPxjC4HufKfvBZhD6ZuwVVOITtElDlwbTHOXiODQagbvA18dQcmdHYMzZ3
t6MLmvV/gpeJv7XjiHgl1hQxMyuDNN7KFLT4LRCf2/xwi657s7zhzuIVWdIewHHB
eubz9GC7D2RRtqX9Y0o00HDKQYDxoY9hrjItKxWJBRCV7HonC7EhjC+DGhGjToNO
YSviFRRGEI7uFdWiwDFryF7k7aR10iRjbsmYzQAjEpesepw/CwPqHjIrWdJLDFlG
VystLADimN8j/LEqvc0PP2rll9yfmqNOPdsJSwVrYEYKlIu8skkTeLEX/yRG8Evj
+paUMzO1mcaTFEKqvwjSO8zzFr8nYrHVqfGBkxHRlr23EdeWi+wrHNzSUqUA8QE1
aQ/p8NcWvHPGa046po9xXT5u1qdmGqS5pA9XppoL4+VhDDAgZpmEHoBLtWF0KHRe
YSl7TG9Kxmbg/c048yrjHxK7Kz782gNw/jFNZ2LUMu5Yx+d7FONhIpjgQQ5WOvbg
phdhz1agd5PBZphjJRZNmAWf2xyOhfb94qyvrBQstcUOglsUb6Ljpw7kN79Jx8Zp
vBfRFv57fC1eHOuA01ycszV21A0NvZQ5lcqLjlzV20Qep4wKYvTvTtOmjHy4skoW
42/iVZ229GCiXsV7cgGuQ0AXtVLmV3Da8uNeMqWBQbj8o/j9xnhW4WbA2SWCxZml
oRHzwp9F/Qs+RjqIZYvh5EMD2kvFJCnssFPJsYzjhhleisaVYPSMq2sPgUur+lsC
0RiGFwjr6suIRbddEBdO4acW86huB68LvWj7S+dAWYk9SUn959UD9X/p5Tg/+JdM
xt6FkwHqwrEkBkHtHCgeNmzyBIpAAocpLhCyabvPxlN1OadD72b1zDJKQHs96FoO
OlauVRqeUmUDTjIztR/L2zmexJMNomRx2Dh4UHX8ojalfQkO2bCjz6uFCEPcxwVy
g0j4mj6CB6bjuIEwIqDpsNU0HRpDqdKUrP/dh/ldrCx62W0Q/hSlb0YujdTBUsq9
FWWYJEPDGYh6M+TC1smvNRc0MMCbdvXC+24VVxOsfKNG72iBoOyYiaZhoygDcb0r
EtMhoeDxn55CS+To4Loo40bZ0FkYklOkwqB9HU+GnW9KIUoGt47nU8j9+tx8vGJ8
+bk9mII7sjUkGvA/NOL3soFFm851/kHHnna9F8B3C445otKMvOXmxcr5Yz2pctNl
ZAViKD9UgPRwgFM/94FRCe/0Y49QhqcZ1d05sMu3HGvDTbcN6zGAkzrC2E8VBR9S
UlXPmbyYlcYzNAoQBHd1y5kLvDCAI3DYBEyEGX2KeWzk9r4cogEPPKGPxnPqPKv9
mH+hawe47qTfunaXcPNom4fXbX2+D0GNRt9tQeobZWQ5lJIEzzH0MUtUuhOJynsS
i4CCk+r+ZB3qBYnBnTlERTg6NruGOqFgYXX3pJCYSw78WP22ssQF5puAaKWmDHrO
NXOH0AI/dXEP8N/UKbTpVRO45TXVAmyV5/77gnCF/IFViEOFKkB3FaJA5eI8q7+o
u1ES89lu7qpX7mM0cq6PCqv/lSBRvYhglivW3dNN0sG0W+B+hGqbiEmQDjDvg8E3
STc5gBZT29g/K0mYjLCqg0rKgO7vjqi+PuHOOXhugmiebX2nyTjGgoFDzG3m6BeG
ffF2Mu0CRMm/rblm/AzDzgAtv41Eu/9t/YoMrmfpzmChCFZbELTTKudwhhwQJMgK
1zBRbw/HbfyCzULLqknQWio6JqAxtj8QztbT95j++H91FCl939XveDcBEOA+PM0H
lLo3fgMA9Kf5LNN4f6zyhYZ1SkJMtXk76Znszu2HpHviK7CZC/mcnvmGdxBZbdjJ
PFbD09j60zMDuXPHRoC9JkTM6ThKGVjFNwcDz7IXF1++d8GTzqdmBJ5KMlh1ihZ0
8oRt5T1Ies5JUdjMiIY3SayUvoq1sE7tTW+yRsCaYeD4EE2pVWPo/O/btF9GvPc+
5iC2gMYVrh7pzZXiLkAtdJYghIF9PMWLUDvP8sJobIKQtMtKK0JP19cKJFMp1ZQ7
IeuGFl79BlfsnDM+dTGyScWfRRRe9nDBR0vvektTLLaUYsrXZE/foK5AVgefuEUi
Isz1pGTVtQrbO8/gMCrnNs7XsRQl/B1nS0EXRYMoyJKZjJsGV7J1jHi1iKp2QVwx
PHFvXKG3PXmAvOXI07BFYpPDaibKs7BnIda5Vp52T2o2+8K71hassb20EJFKEVEW
7hl0PnUgyPKWqm3RZbRtB2TKGUReJCVs5VN0UbM+rw5dgSdxw1KS+6A+DXB/rDhO
ejtBhcEtzlthzuuooSCSTCVmZBgYx7EN4oAQTUsMRdH0ot5lP35aXUCCD1K5XWTI
xCqWWhchzCsGJ6nYgnfWKVm41f6XWhxK615OrXOByEAvjElrV9iLCX3npjusKrnr
lJZLyb43Hr8GAPM9VkBmrqvm3SI72m/qbQ+CHmVOLdeiT2HdMRBTp+M8ITmKwYdp
AO+7HdlCmK10KwSAeSz4+SJbg2Z5IPIuKHQv6FAUld2UaDzl6bkEPl+yTTLeDALT
1jysFXnIgU9Ry1ZtTkN8xunL9yv2MIVtQKT0mM98G11fJsSgREuACJGSIGIPBMPr
PODCiPODygJk8sNVQM+k2q3YzWFgrDim6+inuBt/J3DPdM7GOA4WghozDfQGoQPb
KcndBCW/ruEmc1LG0c/MLxxGlXIPJJ7Z2poOqOSHof54KvCycUW1bwXE8CpxwTwm
kwSMTgQ5z+b4Yc2KPVqN4Ge/SnCQgNgpKnUiG7QRFqNSoGPjp0UH7Z6ioAKCJRKm
TUaq5Y7SrtggwcSRm9pItvE7/BcuzuxuKts2/4TlsjEPhOHulQFhhqWASLSGmR4M
4QcOLxtifBeyG+3l2xuC/mF85Hb7eDQNWr++nEj21+8TbBgrRf8u2E9kknimTaHF
ZFVZd9a/ST18Xgp5ZJOJ6EsnTGGnP5hKGaNb3b8lantMKQ3JBGgk2lDOq7qmp3sG
Zf4d6llX46+xEge8F+/q/4/GgZ895+Js+7ZfeeyUykVZT4LWT4FeNikvqchHescV
/7+OL32KaZoaagkPDN5ULNr7+0yRglmAimc2TF6KDcmiq737REDuk687EY7DeKs1
tRup2YzoBR1GiWL7NnnNU4V2XNZv3D+3uFuR7R7VR6D7msq00L6cRAIbfw50ExCU
NIuYuhj4LJlxZV1JEFszNpC/Q+E/NuiulxyJxR9ETh0887ZVDFRBfn0VhJT/OWcj
KQQImT9p/69sVJ2dJ3Bn1ZpIMsYG9taSwL9o842rDFowjlkerfGPCfJaLdS7ryir
iH57Dk76GpzVLCw/Wy39qxd7IgW5U3elGF4+M2dXchNjzbsuRUVWndL83tyuarJr
wmSmJ2aVgCGD4F0er4c+8yuK4oewqdENZC3b87R4dGKyMShv2jLEV1qWo4TC3nNy
ll1C2/ldJ5FEs611p/x/jDzVpZt4otBvgxvyJ5rkJXs7mbBcx25hXZ8KRLLOO74A
+X78/k4N/hzEhGKE8bCXRn+9bCZDXWID1N8unRwZrPfgsnw2iBR0skxKCI27ARbV
/V6gXh33kYnkzqnK+juL1CnDtw6qzbSnBBFUefjwKLLn6tpTUnA/0VvVsbTGkX9g
/5is0FDbESTskMxiCiiB/vpBIkwVSin2HjGRYdSzR7dLoBpfcrCGnHj78hAvyXRD
6cCLK+G2iWaImtmYv3syKp9h4rT9PgE+PlJ+S/XT1+V8EU5SiRutu4clEztyRpRF
YZm88j1JvuVv9ZFp1jVQWUg635Mj5pBaeDK9PRfxukTf7RyVrFDlKZE7gC8WJXSV
8nQeduSg/ePoEhcGQTOfLIAHz+BeYRSGNO9aLuYLeRFgIr25tUGzD6I2dV/hkNSw
1uNS8GjK059WUOKFGLeHJK2vyCFqkueUZvD4GV0B+NaX/msULJziQm5YzGjwaZdd
v84q9tY4PMLC3D2gUFasbpbM+LhKc26kAjWW9tGWSkwiAHe8UWWVNWerynSrHFma
deCSuPgCo/0Z1p1Z4LRm4I3wsMn8K9/oKnqJ8jRqy1i9lFTmi7DUQheJ39WfXUJo
0CLdIvSYU3PyyRidi5AEIB4cuZxykBdrdfbG946CbAL+EUomB8idTaxk5HTIF4ah
4kHuWy2d8/km8vNC/ZOOpJtPLUcx/TyLV/JLuW13tVHvJGXyDSscNzY9Jg5vM3ir
8rP4pBf0na6CvmqVmUrkdQNWHH7252fh76zMXaHykMug4mhDHBtVqz4BsyiZz5j7
N/UTCRqbBaR/Hv3+czbO1B0y1DcjewzrkYkUMQ73qqP6K5KQLuQeN5vbJO9J2Sjr
QKjczLhoMn+1JJCaQmu8ziF5aa8xu3+gdJBPMpVw6QDVPTlnYQ67zGQW8VHS+paG
WlrNI5HIFvKYpd/7guPskoWLYqjKsvhu2nYemNFk1s/XbbhuFu3yViXw1koSfTIs
drlk0mUjNfB9NMSkh9VPGTGGBoaDffR6cyijzZ+UHLl0/jIkTNvxRTfNYE+yt6Kh
UXP1xFmAcYIJQ63al7n07YFA3/8vTHsDEHWFC3As5LiAqDySWoKDOt53Z5X+tXlO
oBM2KbT5SRsbwNJ1tVwguv1ZyTmCeBjDd4tuT4ilIQdk9cXOplcvERePO3tu7NJZ
vJ6a4BvuyuxfcGWtgbNrCUylTf2hjdOYUZiqFd4ogBvsSxnjcXyqF9PgI7qtlshu
22VFUh8kIxk3VY0+BRZHkifrfi/nADxIafV0I4lfa7MSSzyMyJqtWnuCk54vJQTx
ivNiiSAL6VcikOSPiCcRwtO465C+tlCn0m5F106InsWDp7A8HTsMoslDXpRJkzmx
dh52JwZmbyeuyO30fNxGAIz+DlSrmkkkNawBwCXGaIp7JaHokIfEz5ipWShCcvXO
wDd5HHCLWg+Sbujo2S6xggMZj+a4AxMhdgSbve+Pik+CkpLKZzWNmQltbh4fpQVI
i3s0KGAZ6mA61Q8Kmv8KAy4G4Oh15Hs6WLAgHKz92XlS+C9xU4wmwELdDnRz/Omf
lYl0KtxG1njfSnDQfrLfVl/xijkPa+bOqGN+D3aQaceYbx4BQrdY3FP/9YULleye
Su5ITr7TPXW5l5YNOIxe+3I4nCxNz0PwSoWODWY5991wi8ZmzzPu7gqb2CSQLDYO
jlKICxgPr6JwCf+yF6crbd7ZYYbQ3LZ1R+e2CLpQPOMumojJtAF29Rp72Hb4bLAj
8mPRkzZJJ/fWXTjZRGvfgcb2WwpoELlr1NX2m1t8NttedTJAvrQhS4TRcgCu96BL
rJFTvt5mSyyM82e5RlfSc3cEu6xxyz77EGkLsqnInvGfDB79JuWpfcGwNEg/JQFF
eg9HQuRI7+8eVThBAA28MH6VMu2oOYrfo+pMzySXPitb9I6pNrbYIUVd37QK7byE
ghjvt2+TM0EPOkCGzdbYceS423LMM5vFXqJZMSxnzlU7yDL488otMAarTT91BYoS
kTwHyITtv7BzqkWOIBXCASd0P2LQkzeeaG/afT/hoAGR5Lv8Nt9WA0Z7qWvGaZe3
xCr+lPbwkxZfpcFyv2RTxi6+mCFaI/O4sNh2fKbh8cCQKgrfHXZ27ajsuoivuopt
L+HzHOIeq9i/IBKdp4pEiPwnG/6+JcBuI9+oxmm56urlHG8QOnNMWc1Oj4x4cOs+
Z9Jtu5c+Oy5jCvPUS+rSqRz/SjAM+OV338M3ciqYJ2L2iaTnQjt8V5VExG/uce6U
tEXIoe+mmt44sKaWIrtvP1hdneYY5s7eJQvkTflwJjSDJUMsxy7d4FSfYH/caG3Z
z8CDrrY+sUNKDTkDKwv05ZJtKStSvysqY2adU7dxn+mDHoGM8Z7iAFIWWVFrRhja
ox0B+ZtWuplWvZkCGeSHdHPvEzNrKTkrZaTpkxzr+WUUCn9fHJjVISaYglN/fLm+
MGKiE0MSP9hoQpv/t5+Y1ISrfHuKVvKIqUsGDL0ZuUgIFzgQn6rEHfdZKzFxWiN5
HXNyPfFSuLIti1yxagisMUiSXywea7yN+uorIDhbqQ+o7mA+qeskO5hPGu7hdBOx
s3fAhtgaTlDbLjZMgmRtXQMUcSno78GcYSNcNu6+6mX+G+vq1I2wHWVfHqzSqfZ8
HeSBf4LaGU/JGG+U3FKaHTx7oL4NPY4OuwNNSt4OXXhsLb9XfmPxzSV30dKLILBB
bB3Cl3Sxo5HJCPAYGFKnYrZ9PKEOvA8cU1jNXNSe9/ZXhBbHG4ecvIx4cH36J/xl
9joIzQeiUnFcRuHnWfXodxRyE0+68iV7QwuUp0ixf1bqZ9L6/xIbmT2HeyEPcGxT
zHey7qReg63BPEZyC7N1acVD4Eij0Ou7qTVVxjtNkU3LsUsl39RFfp2rZ36r0t4y
iUhdFWeESKlp7KLa67RnlHwKutVMq3iAja8rRiIHvqliBYRlOlbIVgvFrdsjekGq
9EsiUoKbom80m3toBgYHVQBs1N3HAaN6CPeYnWaQoICu/k5cVzgUhdRgsV230Rt6
YL5omfg6HBsfgGd3j8AZVEh4nQVGzmXfXt1T4iB5a2+hhO8hmXK0whE6J6HO2woW
aAg3G6ry0oSDwaDVTnBIOyuRUgfbxoyKw8LB8dFAQiQx1/lRM7jKn2xV8Sl9cm0B
9x7ez0GKwa3vlgXE/Sx87H/FpLQvJbUi267owkDgvgsM8ZjQnEZzb5YCqZtueUwg
6L+v8hSDYusAjeitjLDSUcX9GV7afyNHKoDEAdPAbeiDMK+Jf7q4RWkA1ndy3dse
7g18AYDtY0YVmRHF8tM385e0gOhjrAb5fKk8BApI6EWVr99KAPOqV5Cvs277vt7T
VXgNtGV42gunh6KPdRjw/stq4HwqOjKCIFxmPUD1XiofYwgFNmrqVynX3jqOWqVd
GShLf+NfoVK9auUORyi2Zpih0bUC2z3ZGPyC0X0UqtW5HBiqXHjJfmMLPGvwolfH
73M5ekvig0OK/ep+CF/0IOlvVzEeYlwl8UqP9MuB+PkdYR6CMeCi7N7t/19bBLHC
+EmfdNIqRUpcmfgzgBVo4wbRJdxCPRsm/zvCohc0/6+tB/nznjAAnAUHrVpT0bns
diehDvmBjdxtou+zXx6ixwwSoBQPY/kL6urHwnoibKE0Kdyr8vop5rUN+QuuVlxD
19qESAWzhPJ29MF50jkPR709rWiuqSPtOXdvXyqRx0GE2ZNs7IgqtGkOCeVhwTZI
RisH0KC/KYGrt/4F+gelRUhz/iiEoDKqyTiAwZSUrGZBSPWNtZkBQmyglLMIY/Tp
PKAXl+4XQ1xcyMNaB0B2RFQBYwvo5kRADEGPD13MZnrXM+uOT0y/tlD/ul2kb86y
zWeDiHLsZdw4d5LBV6wdGevdmEtYnCCifaQKYjbpXgVSt+h5HZoq3c6S5D1VWXIz
5kaFzXn+6IYvGUEF+s4DISEU5XpffQDFku3FLHAD0j/NbuG9K4TWGwF7Qe/jLCGU
o8GBqMrgGuJTLo29FeGlFoZ7Wv45IIq/v8W5hNVj1jq+YWR5kbOt8K+v6mLoAuOF
+7cCcf/YNeWPYSryCFW+e0tYHBeaipBlqQCqrNvHk50bupR0oA4KlzcwM9QAlXp7
B0APuyOBzS7qo2a32kIgKuQYgc/VUZd68DAYnDcq2vl9vu3Zwm+/fb+phpPXEloe
SG1NcbeVcPKLl4bbn1avpiPfFMm/Rl7qeT+OprgoeyQA7cA7EPN1l2U7WE9a7mxK
/aa6vK39q+OsVrOF7FISX6VCnNKNal3fCSLuzw65/sv3Ngr6vg57vfy5a6UTWTQc
Amo8AMbxkGl19jtYzZKdoOosEU4Fg1maSD9o41A1nN8fZMXiGK4tbYBJrs6lxaiU
SxXlfBZEwo/6qMUU6sJuXHA5sosJMsdWCuvY90RKZx6jBwpEUlQ8dKqaXxfCmyo0
kL69Njht5YEhuimH519CI6fA+6G//TeSZBPbga4x0jQAxmOjmjFohuhI9wkvqv60
LC9+0h5X5wpW1j2luuOFpPUmPYMgGwQ1UZQYNCswup5/OJxpV5lWHcJE4G1MbCvT
FaaLujHAWPj9TM7N0dzp2Z9vXpKseLsQU4FX6T+1KcoMc0Jvn6vqEVCrQjTZ6Jql
H4EgTC4pLOLE6fPS+9WdU21Vp+CteGIZXPZ26+nByp3v/j83tOOkZL3mI3W/5i+f
f2HDyZrD0SJO4oIaj34cfhJpDMn9vbl+pyu6xC56FmDkRmTZa9A0DQBrfrDYnaMB
XsjSgqYCqZRAaNSqwkQJrl6UPD3OQgKimFktmAs2HipD4JWy7gbHHdVtpsVT4EMA
xseUf+XZDgtqXoZk8RGUGkPmP6FcELqBRU/dRvdBD8JwtdPX+B1yF+0pyYreJXtr
Q9tDB73piY/+f0ePAGN1HUeUShu0ETdESEIfMFwafZJAkiprLaPWFTHzWbvFmD7r
NH3EGWWKK1CCwBx5W+N5JtBNlMHQrjm3AbMj2KBBMOYG05QJ37PC1VAn9fUOnxle
f/s1XpxjU9rNIxrq/nVNJcGCEOtXT0e69kZYS9TJcQ/BAkiLvQ32yA9PY+UN0bz/
V881BWNdOH8oCOI3UtaOjjAttPEzQOn43mpChYKb55S+k0ko5AIC3+z2l7rF9cW6
CWxGye7uR8xmEnGapqBeSlKjhiDXnLT7pbo94a+v/j2p9UHp8lsiklrcH7q+0ueb
ckhaGd87tC0g3tQJqM4f0ByZ4tqm0cSc++PxO+P31XMTyLFYpAl95nJDcar57Ilu
Vl4O49aO00lMxEe8hfgCQiiRHBRPWlCfIMo74diKFRSu23iv5fmbRlf6w5N1KgMg
i+0NysplBCbF8YcAyeFSzkl8hU3Nv4g1RATxTwJ5QfuaIFTYMyNsEWN5fqJhJ0Q0
NBpKWyPw7fN4jPYvbh0mlGjjB6Dl62xI5hoIgU6obz9OIRDZsDeQyfyJezdqDsyI
/PiAFuzpzfflUiZHMeUaUtuV1WXbMVoS93msLaANA5N1uXCP7iCofgd96lgiIKWQ
pFBcBQvT0jr8A8s1ygLeEWos4miBFz5NlSAaJSPlvZk/+HDnPYO4+UwT4PjEKJq/
BOfMgP6EETfUUmADKRJ+8AIS14jPHQ3rPuhfErnZocflI5jaCFaTA8FjJqjbPiWq
2hFBiDVnJmmcw5XGNM4yj4Hcq8P5DF9s3etB+2MTlCmLFkkysg7oynFjlK15Zdwz
esH+T7Z9cegFE4SZCgCoLtiWJitlWptQHLkk7pR2C4ZpRFYzeh6xer1VdrEC2grp
6OK90q5cMa4iukI/0noEoXiapLRte9rUv0t8bY/D4OYXfqG6nWPfYrm7PqkNrbK+
E2Z5/pcMPhboZ9UVUrPJAjaqFI21mKMJA9IKqQrLarCa4akbLqN2+qKBnm0JQhQU
8szlvEo934p+GHeUMkrmnUGd0UIKynvOEYkCq+HRUxBVMCSjjLAl9Otyj2VUgWZi
zEMQ1EFT6aqOj1pch8p3Wq146FmFkJNXIt4phySopfeHwAug9SPdZImtj5uzLQ8H
WpF3Aq3FLw+KCYx8WmWzyROYCJ4IJKOkDwsm/a9b4x2RwnffJmE7/JgOjaFT9167
S5NiYGBkM9WLsDIonzD4FZWw1jVzZdkwI3g0yLTULUc3qU3956RF0QVnaacpxpJ4
5IpSH6GTHqvKDFceVBiY9zRkh2VfzfKb2CamXD81Isuaih5sfVovQK0Em5KbnEA2
bEP8Ez6G+/2meXEX/Jrx0PfOr0wwY9MvCakDYZKIu72BxMVhiZpj7fYuLlPG4KqH
6nQRykv/RI9CyAmonPNEygCRN5dNX/fyCj9uV1/oS2nVGOE7gjn/72ivhZ0EpIKJ
Wi2TUPpJswSZJGPsvKNCy2TcbSJ/4Afn1P07mnYgxjkRZZBBr2rLTjv/VXk/OX5O
DFZcDRp82iip6GXXC9hi/VHsab4Vc5phIsRmMRWxuGQXJYQXhU9Y18yMNOeT9+GN
s0h9NMYfjiaWNSWKckm7V7UdXIDPVHLiPe8e79+xgYFzbecDC7Jk/cYEgd4ju1Rc
qpwfh6dWTTOytrv4a3JU6zhq1ADNlkt0lDE0pwp6HcrZ/q7sX/EZlzev5W+h1kqW
NbrB78+1d3NvpBznZgkZlpImNlHAhvoASmmHcZCkids6APsmW+/to7KOLzYU+QHe
WrTqDLm5MSIPeDjLVICJNhmmCIVmxEN2yX426rRDhFFKyjlAQjkT39UANh0yhcSF
jLND7QQf+fi82UNhB43Gq1Dt+XSYxaemsqRZE59NTDNLoDvdwfkXRCVpGajRkAxf
1y17ECgPSA4C+qcwqgoMw6857ZsMy6Si4zxkV+yoIxDmtZaQEgZbxG5KLR32VgHI
EeHtpCGLyIZkkpwr05nZzSXgIjYkrJpO4cxRiSV78r/CugwsCWYRbE6dGirlsrH6
qp0+SmFwKtDlzlOPts6BfuOIw3nT0A8bjvr6noTzycNbMwmzlAvjSX6jVCEYGJ7G
JwtAfYu4PtLI3seKz9mimRreLMwGi5wXpScSPtvijVYzCUHDAtAvMQoD83ESkD4/
VstEcr5zF04xEp9VAL1tYp/tfcQsiknH3ECcprpyABOa29mkJixzRUh/zBRbGuc0
A7xv7eLEttvbHICUIfgQTDYU0tmLCbujAN7mIbVSPsEUsPBQEJXfGskb8BHYcTQx
s5/rDVOz61mNWaIUkBU8QzV67rhQHDPU7+37+w06eUWyNix62SrOB6a114t9PN01
TKHNmT/ZE3FszZXGZ4+TlA5TKvTxS/oS1KnLcUKEownL66bK9WeGBUYR67XjZr5v
FDpdL7Ofar416M6Tw7/jV6gpU+f59nIFUxKMkQdxLqO4j3ZRH6cHF/MffH46m+zk
1UG5XWWqBO8BX4YG/EwQ6nU3/sYzY+mDVPmLuDUXbOE19K3XEeK2UVPFMryZnO82
iatZiViNwFSAjnkIXGxWBtLJPsUtfQDnbdATYoPCDnydYLSaSRiZPhWlNwBasvLE
KkiGKuj/RUrVDzebjkLqri6juFOl3Q8oLm/O5O5fvrQoouuKeDXuGfmEh0XKbOw7
eW59x8u7BK7GHKchFlJE8HrxzZQWv2tg6L8Aut68Da1J3GzhIke1VKBP+9yOKwhx
AUynUJg7uidwM0oI1WZk1TqACoYeNYYv/ZLnN4gheEJO3C0X8UczA6bFsv7aAW/3
4Dghz9cZUib2E4H50p0bBUh201jp62FAffFgJjt5xi+YIwB7GvYkkVZZR8BIAKEh
Xd++l+On+EhF0sZilCAHZk8vxz6I8ABOQz695VOmmmXPAyhBm7GlKHf5nijCIg68
QnG3L7laq0foglr58p7n4VfDnTrmLLTeeyJ/Rtp8qUrHw7UzJUdlcSFyJYEz5jZl
VBNaqhJuzom7ltjFYd/dvabst3C4p57dN49FCvFSBTE2qsy7HZ1Y3ZaPtcb1Vu4x
RMZgZUP5obtZPUQ1D2+cxn/S3AxqeJVQA32tqdEBo6N+3dn31++PEGndOQSbtGCM
r4Jl+5464L9do9cZEm9MaLMk0aWGF4Ig4DI74lwnci9PDzKFLcHgHIzvxiVXYHD7
YNZkhhXjB0hESGXrkujNvZgWLuw8sWRzYbE2t6xF3y0JR1/vt+mMvodhmUL0E7cv
Sq+l+WFywd/No333BUOLXa2lelRn2W4IAK0RVH9ZyAz+l+vlSJm3wRyo4ZlzMgt5
KxBmQS+CtL0RFDiKdDDBM7ZGAYBWPzwpdVHFEmCnU4Dwvg++pbb0bcgFDrK/Q9/o
29DFhE1Qc1OUujWm4KjtUPm3YqLTbgC4w0BYEd07qStLmKr6iuTCMjQHWJrx/gAs
2tRcKla4wTfXetKidhzoRBhep9Nfd2e1uG2MtZ9b+klDqxd15EznDQqrCRBSrNwS
1qdAwg3fxGcWYZC/QpyGJfDLdXBjI2/4F98Zg6pmdhz5edcoC9kzgDMdH88kwhA5
La+AeoBcsEja3PwN4jgxTymZYUrzZCafWyUJPRlo7gEE+sSIIvps19gs5cU5u+12
5GzLHQdBfG7n4dfSenDuARBxMu0e4ATi4D2HFw12hOjdlSQVtc1LMih0Kp/fcV7t
fenvC/4IAWUa6h9OylNprwj/0hpq0sa0vRjSWVermRNsJRhc0OubCv+h7GpF0gBB
Wn+ltYKJOYWCmNRZ4BUaGy1ytLx1m9zN73L+u9PQnHL4OLs55vcOuHsJkAT3qa/A
iyYfyrr1ChgP12KAC24p1DLdNGaBkndu1FrLyXYa6ubyCKatnbATws96y/9Vgb6g
CELTb/gnxZ0FNUFepSOxNFQpqIzA7jPi9AqC/o05275vF7QBTqCvYIgHhe8AXgLg
50WGc/KcEYQk8Zn0+HzieNhCDoS6mg+Q6Ol42aPUwEq873oeRQ8RNm6kvDqzHVcl
raGH21FYqjxR1YkmSZhKvmxn5z/ol4IBqzxtvIEu57pud2uDJhytLWgBB16rcQtf
sK73QfXFJzOl1tJOVsNmjgIYVEG/G//biohIJjg10tH6xE8uIZV+5ImxxFjzneLO
f+hyuCvPzfm0p3bpWSRHTYrKR6DptMLztXaMqqI4FbzITtHRzNCEvVfbsCd6nQ+p
t9K8xAVSb/E57V3qubUGHlnPvFcyfInmZ7AcqJXFmi1QzCv9J0T4n72bcbfOgUnH
XgHdHOrwER/P6OYI6FcReOwIG2w/8zgcv0gaVPvJirUglMCiqdaW1Fpw4vT8q5a4
TZG/oheB3K1u/7C3cNkIq7Xp/fPOSkR8eL1N69tZlofB1LUVE0888aFzqYCm8KFr
9+EVRcNwn85XkvzY2JYRgGDFkdFQNGsbtawkXUAV5oUt/qY/H4L3jum4DQD4cQzi
e3w1xwEy93N8UIURQeXkWxLkqUSI7Nm01x8x/Ke9X67QgiQ9osn1kJeo+6fbpBIR
90HsMINQoLZvlbb5rrXikrwW9oLKv4w/12nktk2EZw0nYGoPDynNc0MQsAHx3F5N
q7f8ak3zG+US840D/StmQyDoYTSYdN5bbhOjtYKPi2yVrahgtj+YHp4aWM8BISAE
dhE31ZoG4VSGCcrAYG3c7ZnLWuM6WTeE3WklrmBEFq2ukvIGuf+q6DHa1etrX+XF
VGbf+kcuCU+mrHimF3DcnseQpfGch1REJmKmob5FK4eR/YRjkQXAFE9xw+8xwdT9
wEWowmuAXXfQGAU5MhaE46wLgvOa46VLYWIJSSzyG+GpGjHN3uSKB2qz6MbmYozA
ClH8/JJj6Xc6DSQfL2g8oEBB37ijqw3Of0S0jC5cMcvIbpF6Xbmr60PmTRrw2Jiq
YDtt8ZazuHy58yg3Z4iW2lUyRtEdixexA1DZMQHYJiYAtt+UYBokqyRhHA3OG/2g
j82ry00OXTt9pTv2g931kiGYgzvILoTXhsdNm03tMECWYZYu8HrcS//s7S5f+f/s
VaXlORGbnl+0w7JUab29S38xquhV3I5RVi0DIYodnrvBOk5MHTVUl9DhElzFDcPu
wq6desRtMFHfnEq7LVqklcAKgFYgucImAmUGjxgh0JYYXoD9C3KAO/dCJm00maF8
45U9VvzoxcXafV8Ux/F62+OhdiPbapW7BWpVvvGi89azc5XyvcRrFmR8OzCkI7lU
pfcuiyvIzHQMfLWvkmCQt9xVks+FC0ay+n9rRSJLycjh4BKQdYJtVfXKLrYSyDvE
R8TG0Ocl+wYioEL4/nIYpdDgD1e/6Nzb0DxVralHR1LlGi5Z3S8EpVJRkin5ws55
/4putN5L8rk/mFZ0Oxhf+gwz/psnytslJvrb67GQZp0vOUrZLxTyg5KS3v9cIvZZ
Hvj2Z3AqGzX1Gn1b6/zi5ElsJQqY0W7l+XGICIHYVMdvffNSVWVUI0TficEZT7uV
0093J6U0Mn/W9RewD3BGOsKRp5Y9WglgK+s0PTeP1OR1Q60yIK1YfXrKR9Gb4Cdq
ihUPrPP8zSknLCMShibSPvgcM2xv/HncXqBuiUTouIz5rHA9a2Az5EovV6nmhY3W
wam2zZzHx9vqLSjzYnHERkPQ3Zfq7tzoUS3/O7IDKDEjZvHK6SRUhOQXnalSqBb/
uTzXe3H8PA/WcJ7mWKDalktoczVRaBqgjZlWQY4jQnaDwo2LAaaSE+Y0ejYrhd/l
V1sjQhnxSgK0e5UL0G0HSgZWS56GLDB7DoHMJUw/v07U2kIA2OLfNaQq5g3vPH/Z
P5ghA+AU6U+X/q8FFAiF9RvP0XZPJBXzFgRABrtAKFmn4gEOV9cWmKC94NBsJvQE
4mHwseaffw7w+7IzUnLS2o2Sbcs1My95RTOBIT5TJTodRi7NQCwHcjl5hGEeQMxW
iGK/jQ/it/abXcKRcG4fBOVRGzKarxXdS4en0oyhT0tw9hNzwjhNeFriZOUI4ttm
ZoJ5+XuYnI/VMUEtsWvh52gJy4oCJyffds1EHOpBsSABn/PmSkwtT7sx7bqCNYFK
wxyXT9xiIjfIiSZqsgu/+QU7TAR3MH5FCNAfRRmMSBNSXtIH/bHKJMIVAz3nPSdg
O024KYOjKLPep3805lXc/0f/HbDguqfDesjkzc5l77UxsKiTN9TVjo0hlQQe/gwX
eFTmk6hRMb16Eb498WbkoQCrrX+0hhyzMkjNmvpPpYsHns55NCgwCFHnTB37CoGr
zTtgDlyEa09r4CxjNFg1NUfgC+UpmcWBpyDYNRxz16nVzknViKYJIrx7twgG/uoo
iM9PZD1GFj7gfdkyNWZmt2tEA45TRYBXlAnJPv5rQdNyHGk8I3USP8jXm8kyv+JS
ET5EQRtU4+3K79uHNxfqk2+WDOMoKc9dTpP1NXaPJVMJQjHHfHwmFTKL4oJVmk5p
Owp1ZMLcbUYdfUFNcp9iZlSEf2HVozTGcEKUrkiWiA6Z7AoELNYx3c5jpvycQMRq
SkrtLjKdjWHqdMbtmIhEQMdDn8rD/9jHGCsoGUr8slbVRZQbDXzwmrDa0gNClwF3
ciSx3k498wCTCoKzS7t5/tzRBGS74+ZrGzIPCGZ3edpX6NKuqS1Yo66SsYvT8UZx
Ng63wDdSVrRwoGSTt460e/CHWWALXoEw7SATj/Baua0McxNZO3oQHpDekLij/jM7
1xCqDhtYaaatPVnB+1s2IYy/I8Lp6ZfGvZMmEx2OfAGJN+CBg/mMV9vgW41a6eD/
q9Cr2TLvikG3Z8fTy9S1T04DzY2Md5/A+bGxTjHwURp16L5+3deIfY4FZYEzaEDw
yQA2Z5LDrqzQNWJhIt9+QDeIxMBuB994pZshK1SJs9kyh7GyK+pG/humuXOGoPuN
BlFMfd1QOKPe4GE1RyN3KOFWO/CscAoiyVY4qGiKmSd1ik9dCrJTdrAUY5Lu7KcT
zu6Z6hng45gKFhV9rgTdMRoUWqFsfJ+MwkON7LFxV1KmsNbAoAo2xh5TlUJ0LvaS
BLl9E9WM6jdiCSUlYX44FZy4BFqG2HvyDZjsu9zHOvn0w2hr5Os1lIlSp34heUxN
U/GbxNkrULMRr3nGEICB0OTLnuhfPv2PYRxVwN9BuPVc2XX78Rm+0rL+W9fjxomu
fZAfyAJN8W5BhL+fzvq7iiZRVtVRhwg8gBowP5Kf+XcN6e+1nnPGUD61Ib6asvQy
vn/gL+1Rhm6W73ODi1lIVjrUeuTbOhEKx6PMPknfjBkyFI5BVhc3cgsbJx3hVUzM
1aO1910g/IDczJq/6IgfxnqQLtBzIfhZkFU14tIBd6nLfEeFsBg9x2tzUI4pq1Fl
oN2pm6lZv+XQb5I5lix9RISevBeaGxzUE7DxFUcC9hqah/F307MRfCNphQIw5L5r
6NtmPVwatY4e8mXM8uiP4fBH4jF2M36KoGKWsN+v0Tfj966natWowSF1nn4ARkbc
0gXQJkMtZ2Eal7A/W4fY0DuRAHKcbqVrygLqcWqKItrJORp/jeWE//ItaTFBvVbc
ELdfduwhZCQ1lonvF1p9xheoc8aKWfj1dI0F3vVVtLVDVHhx9ePeqQFgNWC8+J1E
HQyjPKz8RXd+pDn9enTXmZZxKmXkZHCgxNr6p8c7RIJrYRoEFpwjPXOZ1x9eaWjk
K/u8Iv9V2706wQM4DZlC27kcGWMJa3K/+6vpa5R9cBjZWqfNN5bWfO6hn/yDbIet
5+WlmCPMGUCO/sLGGrpm0kbffNCh1SQp+SVGJzttuKb6GZy6heKUQgbagf1WaWw7
yo3yLv5HJ1gzQx8jy1x/FRdkumpoeFY2wKWCc8XsdSz7Yw1YjB9Pmf6AUX6FOoF4
i1Hxo3zP4id6OyPiJHlCKjsN82gRgHqqcZ/lvUi+HBrSXPX9B08fjeINJmKk2U/y
kch1Vc0sCJTX4DZ6t45nq2bHB/JQFB8NjbWy0vtZQL+EtM4B1AB4bBJCsHWlmSsH
h7H7hYdQ0K3+yJ+w7WFT8ZBBtA5zMb0RFjA9BmHDU9agsA1s4x7VSKRUGyJSnjKa
84iH/HIK5HGp5x/V+6jJ6+ZIbGHKFxLZ86H3Yym3ccZuyRveWAcTAFWzAFKYqf6G
WXh7ioZpbJgdVOv8zemt3pbBlHjkl//Zy2tTCL2A8ajFpwbFuEJM+aBHtJqr9qX5
h6Pw1cXixmm2ltGP04bNSSk7eoYW0g610o0c8Heowd1w6aVGJwCNQ0NWBYAV1rCr
xpDmYefyTzG81jmOmkse2KlJ/B9sDScGbCBu+ERZ7N4jtm+3sbh3ldvrRSYWBsDr
SSXO25Sk/Y+HfmcyKFLaYCJIhk5JDjTOVwXIWx69gn4jj79yYMS+p9o0fn90BO5E
0VFWrp0BPyy5ojSu6EnZ228UBLxVULKENZMuwUNQMDe8KrcKAPBeKo9CxVP56HW2
NdM155gMpu/xTMALd8H05+v46IXqU9Bhe8DaRVfSv5ldZ+0VChJv45VGvTzkxDYh
A1FqgmJN/QYpqvMF272ouiAnVDSg7MnKkl3e2Ev7Z7k0Dv4CDfldbsTKomQyhA5L
2SRwX4uNcRy9sJ4VMrdLhJSYZQH1DYu2bdw+m1l9HjZFk4WFdL0YZopwdIIDAvWW
O0X6sj55u8lfLVpQWVaPuiNir8zAUep48tt3RT0UT1wZTfYNdtGNADZyd6E4hYAU
FoxCCDlCusCT3GsQ4AQh0+zxRRGYOu8AZX5t2bO8ygajEAaYioFCcyefsWuZjs/l
WFElOr2U8IarUMWJ2KXLX3xCebkk2SliUIrNBJTwfkyf76gmbI/tHwzHmkAxkgqN
hO0iyqBaSzt+riW59iG9xtnD/mL3LxiV4v4D2I3JX0TcInrtjSi+hGpTmlVrVJXS
prNC5VD89ZNqyqcoiFfMfvzxyzEhVHkEeKRR9XDlNHqDdZriA9uf+/ygDYzC3f3l
ZazUPS1bb+jcVlqEeSz+ScnLVfkVK/pe2IDcUWQmZvSd0HYrA3LnnLXy0gRjPZjn
VUI6B64NFe15q8cK4uESnv3WxTp6geeyqgGr+U+9IQ34H5rYt1g5BHxpOjaT0qBj
pbsKX8wj4PVCNzcnQ08ojvDEdxEosYgRp1fwfXBdSvSVYzPPkXIFJ1dye4o+AGCc
L6rjH5ak0vfborAP6B/cGL3ZdQ47Pml28OQtXxzL0cZryU+feDg+BxEYx+ULkqTy
/NCNPbYiueIYErtFpxV39pnCswIZjCtKRjo7LtYQ7+QtEFv8D6gZ9wyfQDyHSrB4
7vfwuA4jDDtEbs0Egqi1TuHsJnBf0hAOjjNJ8ASiHhHH0nKSFwuzDHSfjgLO2r/I
tfy9c7N+6HRnPH0lr0XRt/o/IwCYgTBCv+I4V6bpznqRqad2bZdULl7/P2gkGZAh
hjaZZn67BlGL6RQDzj179kDzzx/GPvlk3EKft4ixakHxBwjcgk/0fpbT1eeeCE0i
M0wyFGwRg+x3QaPaefPO7JQ9/khZaokDgisBay6pLMbJmfJvKgdTE4mjCwWbU7tX
e3t0aGO+cULAnZm4BsaskEJV0LwHw+EV7Hlxqi9HBkN/1PhX5+TOWu908k0rYkrw
pjPoSbfsYT6ujltFlRwQaPedgsNSdZaZyqjjtgVeIo6K7U5j+vgwoHTRhjtAQQwv
NUZvD3nOr0sAcWYrr60BbbEdByPVGvp7u+hPDaZFH/zpvDhySNZz22g8IobogpfK
V9UJ+6ApnKO4xX6QuCK4KwRH+7EcJX+p4sDrMEpZdipfc7wwPI+Cu0Q09a0DZeot
FfIk61HgScU+fR9jcpLrZWEPDQse3wZoY3ewviicKR4liEvSsQXNr/WeDGU/kQO/
mmnZZ51PPaAEPgdnWTLoWLVK6UwJI3D8Q7LX6JFB6xTsuzkj9mEa89PxX6QEMZ2f
qW/tLcglGazCATxOIG//02YXKz59VNyp8mYFeTpSFxjLTI0mNvT/9HqZ1HNduDlz
AuMUqIAlyRzB1P6fDp46DvRHZgxtW70bL586c9VMxTYAzkpGXIyTKJSL17Bnna/s
VM7UtS3bpOXTbNdn6QwFWlN29oh5EDmYhWCLiiIyazXo88BcxlOT8yrfnjwzkAdu
Yvy3enmqjoFh8Nr2hI/Vc5r+Q2vannmMYNmQ5ENy5f9jNq0lltDsg7NNarkS10I+
k5Hys10yRbx8xmexUuVHb6eMpTeSeGaHRlI4FVtnHMUnufDMLMM9juPNOzKBXLrw
LwD6m9G9ifFjs5LIkSB7WkXa55lOmT4m8wtrwXtB7VXqvRLlBvdPL7uWq7V6mSbk
h6iea1BS6G8cMPuP9ua9EvCGeK1BgHb9y7G4c5S7rTBb1qsMiqtysWPy+paSosEA
aJa3A3huawE9rskIfG20L4W9m/q37mJLQSv9hFBA1Ya+7m8TKYrYQJrzAqzID/Iy
zOHPdjbaHXMx6bDsujSta6/gQlzGOLZVa8SHAL8SMhIIaZOyqSZF5xRAajZ812QD
TG0cjz/Ar1pdXIhQgh9LgUHnOsNGEGnqTXqguHoiPuyJJQ49IcjObs8cWVwOs2LV
+09Zl8JXiuiUyC58eHxbI+NI9NpbXURi5CDgEP0qX1zkj2JW2v6Rpet1fRsLhEQW
t4yehKKSUmTMohulbTUCdf6zj0R5yASnWkXO77S7iicFRcRZkiKBb7cbyxfnhUxr
yinPviDUxUkJsPgLPqXyQ2i85dghnXB9gKg9CjVBFYvwe+5LXr71hAILs1d2FQz2
2T3OMJ3JYdQX31gv6SU52+TzjLsNgCrIW2nTk6kAYnG0g+L1nQDm1gnD6I0mNuNT
ZafgDFC0tbS1KAeiLBlbhfG3jcahFQgBF2Tyruc+0NIbwN9Inm64wXedsW6zQJXf
KjYyKkzn7AqbySoMXCJEDiLlPsDs/+fbE2ElOIuouzY8xMkznoRddhQBBxMFW/xT
H6X6WS875lGLeVtb2rOKzVj9JH742K0230b0vj0Wx8LCqvKo5BlgdHtIsdnUw9Jt
1CdXR6gs29JBcclzmKMtp5emKmFPD2VtL/HV63mziTwtCZe+dVlE3ddra8DPD9uk
rcIToJ5i1X0PDfX7Q4WmHlqPEo9OY+XFkXQhK2U25MzW4cITqLUMIFe8AHVz5H6L
YcVYHrMmSlhTgd/yf8Yuh82lrRDU/ojuiKVpSwKGxfCDB3LMmwyJQU72B4C+vdmw
ovi6RYI7JrwN2Srj3LyqDynlo81TldSqBuED1q+VSXLVM3b5iwzb5Vob4Rwvwrky
US3sipiON3w2Zxy2XD1PwjxpXLGeAZaDympjdpzeL7JRGrDnVfXooXORDG3HICqP
kNVWYKjROhKBVfZFfjupGDdl7gogSEc598zPDbESP8Woc2WrmHu/6tFkhPTO2zOg
vatM0RRi0N5ZY4B5pqYwgshEgpg9iSqTeh6esHA0l2fZnpochE3iU5GQ92jxUVou
tQkbiGf2AX23j4oTbIyBovlRLm/nriozz8M8qlm6l+UsqryZUTLqHaBDF0Q44BBo
IaLUNnIRetQV/Ln2l5YYnPp84+aaXF2JPtQrYPQ66w4/kXM5BTx43HmN4THY+mA9
4PLKteGG2C/BxgOUo1qoT50V9fPt2+Ac3oE/yQO+KAM0p8eZTemvNbAbfF5Hw19L
VDjrQncx6inIWIeH7ymIt0T9W4byv1zSVwV0HWZKipTOQx/M3edSrhRAmWLLmgiL
sRXkRcbyKofEZcauZllbMYjbWb1RPI22JBCZySeOmeGP8a+6qiWbtbUHy8whRVlz
+TIIDQTejerdwF+R9VNWbsuna0XRBHeF5osfb1onafkRNywgNJUPEAU+i/RFVEoo
U3dHqcukUWD1672FNHEFibgO1PDJ2glyol3fg6ptvMCiAoJkDk3TNx1z5KhvsUp5
BM904E4/X1AoadzDLBZUuTu/VrnK9V+5k/aAvFhBYzX3lmaoZVdcG7CJIZvKCeEy
glLCcyXCLO+FgPhdUbAdqjIsoX93Xn1f5iGYCFoQDyAnSAmsrBhFNYfKJ6v2De7y
hU59HEH/u+3Y0bOzcGUkyAR+QYCMIRghF3m0teEDI1qvxthtzqUMz07O7KAIc4te
WVtUAfyczPb3JGrStK7gVCKwwtnZAgeCbCQyus+rmuinEhJEACKqMV0q0UrPXATf
Y3dC3K36yPUVWnIXYT5LEGQz4VUbR+KIcAyn/9HmLMBCCxlqxvNNPdo4guFc2XgC
bLEScCY64uBNlvELMZraoN55eQkuA4MTwD/k/fnxxJuCEPQLH4tshMvR6Io9UJJW
xdHmk8kru8uidjX7G9uucpOD7Cy/aZ2+LEW+eLR1i2vwePTqPvpWMFVE8ZMMwmph
dTdHJq3d37fVdGWQjW/5Rabia0MPEJK3o0SoEkBzJJM8dnt3HpeinbQowF79RyKh
Q19RZEoizIHWQMt/PXlX4cnfaMWjtZrxmpTM/QcXtQNWfsYaQ/ZNxqt/pSB4/9u7
eJA6ObZhqGQe+LXwJH/1ta8us655a0AphmVdpjABmgTVaslNtPEabsqkCYYiG8fc
e3wJpICOntCU6miz9SapkuVbyAPZKRb1HsLZ58lkfluJVQ0ZhnCXZmpI9CFtGwZz
Q1q8ZBwG49CeJYJgyN6uF5MAdICi32ELl5YiH9O6sjENgbl0DdLnhc+QsB+7WPsj
yZoFMjbghsiDts/sy7Kw6hgvrw+nueROfoO5YvK1POdGGt1XsX4gopGq48Hm5VCb
7ctgKwkvU91sJo4FlLm2xv29wBgzLpm+mhHjFrk9UO88B9+7moAqZ4BpFSZ34jSy
WuQ+oabPGHcLY2cxlq+rhPnal/Lg0JBWOzQzsBZCo78eVQNxS9hms1GwwH2E10J8
s5+z5VtuwqQkpey8rutJbBX/N/Q68QGc6HW1mvw+1Z9y1aU6bitjsenQ5sAO/EeL
Lhd9LJ5V54VaiUjKn3SU1Kk4QPS0qtSSRelYbr9kA1+nci/q0JU6oIYgLTDDAoBW
6ydK8ktPEg2bYPZCBUc1mGbY24f9TYXf2C7Rs3GDk1Mztbobx2eEiFEHKl9GR4ZD
0RIz20p+zZlOeuWcoE0HzXiEPqnhUucyH6Mlhj9RJMIu/a3IaG9dyVXzmXzcUZPP
R/3Pp/rxs5syh44e9AzHjGDqQcISWOTuo0+k6MVXY4DkhpOnkC0ncNvD9Uzx0612
a99Cu2p61cfMt1n1aZ8dYdgw6EVm0kuHdV1OgOPH6mUIl00lbwruqnFI0N/N/WaZ
bB0eo1CHxwx0Y9jDaX4SDPLSlZkpV+aKGuNpCOpJ3txDqwbgMKDQUsYbM/U5R5xq
XAMWceDd3WZcrccR8LV3UI0Nh4sSRe+O2ZtMCDjRr01pGd4x/SnfFA4bGPQ/T7it
5W8WYqT+g5gFIJxmk8LBuFV8TDwTBmudUxbRj//17xgNTrqhdnN16YhLFUt2u01p
eKdR5Jg3DGFg8ktD9pG07VwwbqTqMjuiYUEZy5WeyGv/HN3lnowJIhYAyfFh/aGE
mxAOBEAXHmPcDzdVxyQpbk0pZuOsKF8OqzSQnOUKvShKlTmba+ciHc2OTytQedS9
GMHBsgu1gx6jt9DEn2YX4Vg2FhMy7gUvGXKNGLA58QyX0CW+o+U81fIS4v+EYLrf
GTo950Z01IzbiKr4pyAPxLowF2ZVO/YXb4DNhwfocqliQfEpIq1MmlHVh3QGY5r5
I8a+zejaaSK2fz4Dfeoxix53yZE5+nI1jzYhnevr0efQFI/q5GLDmsHSTstydI1P
KJhDUV5C1TZQYlTRjulmwv3xA6M20LLEmDDuopaWhbLli/wUbZmRlouVRA2qIlbe
QXCX/dNU068KX9ApQTBJMsRmh+gMARVFKax1fdJlGR8UoPL5LsdcayAK5Yhf1Ke5
eybMwTTV/GbW5KFxuCbdRSG40j12DpZX8QGFk4uX+2EqvhgAmdLoi/IS02UqYY33
IK9yNsNimwzJ/2kE78Nw1AzT9hg8aBdPgw4LDqaHWE6lAG2vtstyBq8f4PIcaE81
35ukUSGa+aqVQbploIf5nP2fWVABY50lXqNDjFnXWnqz6LQjusYcxtfG+0QSkHJC
mSfox9EA3ZKi5wbc1x9aRn2j/2f4ZrOqd/7OWSQlMbIyNRFmcegNsqgrTASHT8Vg
8Q+CqN6HByeANNzUZCKNNT0ZVu4Kjo8jjPPs1rl3Y93m1mscSvQdwo+2sRuLKG+k
gW1vshndkExIJXFl7lTo73C3jngrtSd4TyugUe8VQc8y4Sd5h6cz3dAaaK+w5RXr
zjTHxf5SM+eqKBAu5rL0K9Py1byEvP7bXU1qBLvCPzHupdSNqjNtekS/vG9EnvMW
m6vIGYzrjEJlx/dWyxu8X7paFSB90lGq6yN13O3xZ0qaY5CXi+53R8qp5AJgB9Vo
108s+QZk1ayngMxzSDgrheKmM/DKkZb/kXIb4iq6JL8Dhhkc7onWchlklllJlaEI
RX6lHT4U8FOcxNGwcIxM55XUQnP0FKDQvrvRy894Rd9xw6l/mLeJI2/rJR3hag0t
g87qBwb4//P3AI6VGuTQO1HuwHw8TF7xsQel7R8T+PI0aDdNbz8Fury4cneG7XIP
VypUKfuVNb9r7z70v6svU1dvXv8kPq306HP34UCEfi+NFsfqY2O3JVzxWXQGQCPN
oTLowfhV4P7bApCkJqk69ODF/R2ssJpJjcxHT9Gzw7X8D2ZTsAc18ts1daCRZfhO
cSshBWnWj2S6db6cVbsWTogjrk5q3CCDls/xaiqxGKDkZcng1gvrQq+jvwcZBYfF
PY4zWVz1iYt/UNszw+pNcs06VfJNGir+GkkjVjkx8WV9FSGl+gpI81phhrx+V8PK
i6JMMEUJJO2gXJqDHg0eSByoHTcKAmyu5gir03VgpBIXuGAliUpGj4+C2RaZsMuS
6xJLUgta2eLe6xQfGTbdK9cVCKLTIB5IPyBJd0OHGbatDNmq/69L5UiSQQO7ePty
RW3EX99h48UcRuP1a1tXrbdgmEed5ZeZF1ngI/NUXgpVhgkx0pSHvL2F7pyg+w5x
9952V9FnsbrngSEe6RCyaVdV4t+kWM+wyT/+hLyqOvIVHOUwTOhKKDmby7TgWr9n
aQs+Boiz4pMTwbF1ifMq8ItZm5a7zx/VcxhraMt4LO2B9GjweUQCkSyD1OKKDT1C
4/s6ZZjhQGPn7uzEuWV2ZD/NxIgxIYnpK1SMSgDWQrafB8Rcg/PimM1dbJrihFM+
BRRs8cXqfhYo6aDXlaKJfkFZe8G4n1jILCBz+N2UskRkelCEU9PTEgKLgl5UHGrh
Za/F/MCiXFq79a/5I/sOqAXKOCL9PoPjVqWgryq3mimASAaktpRh5mgbUI1l7xfk
+LlCaP56h3GWp0/ZOhE85Vsq5KI76qj9rzKsHWdJ+4hsJiMT7bqBVm3nvXUQaHnG
eJ8U3AKWxK+XSnRFTNQ1TUPEICdFyHBnMBKrw/vpsqRa10sZ6ke7BZjW9IlCZCwl
mcuFWwYTK5Jbtx9al+zMlYEHDERRoyUbov57zVVp1JB0FiN+ckeUMfx7yq7A96rz
VZjkdRAqq6d6KvT6/yVRonAduzsd2ASoasr0Jqg1VqcH5jSqwr800SKv8gN/4Xzm
13MAmqvI0JinYUy9wVOck9p4rWDkCvzGxkEFZnAXrFbBCqgbNr1+TcQhsyzEE0Ui
85KlCiy5NCrWbUzIGtxOHvrmrEkqPlyXJqKy2awdnilVM0MIZqEeqRQ2Cy1Qn6jF
OiAkHWbypahhr31OLvcJg6vSd/8kpF8eM7kLzUR6ZtveC3TcVNSdduQj5zTkUP+S
/NQ8F2VjSkWW4EKYNueCQPQOr+aekV2/ig8aUQy1k+s356A6Rz6MqgMCssHcd3eP
0ZMj/0JoNwDSgZdfv4tOIs4d51Ov1RbqkvfBdYLtlmaapB4f5EvOXi4DJghYqvw2
7sFOtpauZLoue04TnF6WuxeVXa4UzXWxHVKoy+SzkF+Cp1hScv1eJ89pDqFhLtRc
w2j/BSRSNw5DNQcaR9fcc/uk9kcp1IIqd0ciuqxm3F+wCcOV7O9cQCHiFBWGmEnu
MSi3nhQs+kJRiNAP7aNWESjrdFKd+sTIRQun1V/ZoFl0npmhaNQEsELXQIB75itx
P2bnSidjulG2/KNoQa01MDrTiK0qvNmWgDsj47nkw9WkhJKYnXSZ0lE3oh5l7mTg
0ePw7PWAy5JprMin82yLmw+JZ5+amzKM62z4PKvAvvfyrMNIqBZAfZCr0UQszisE
GTo/4xHW6zYybQAz0JVJjqKd1bynJbpJWj+JY15urfrAwyv0HoFPeDiG8tvVLRrg
z0C8L3Fr0fImWtNKTiVMPvWga+urjt4v25wnEvlAEdAVWHnddKJnB5iC9VBul/m7
oiKIiqSJbScoGQYRdUQZgERgHis3wVbq1F37pdWTjQO4jalVwa5yqGlr3II4/rsH
al7xm0dhuPmqcDefWvIdO8QV1usxNgk6WEHBYUUu+U0iMwKUTccljPQqJdQt6AXk
bcNkXYcpBb0oKTWy0HHQ2ykqjIHVqo4WTolupayR3terpl8V5EW1WO7TJZOnvwPP
MEgG+7lZxvaNe35QYIaCVi9t5uK5z6bbw+GY6BJUzWYWd6eh84fJlV6/GO8PTbJ6
3NTYeMwM/dqhY+GfJ6xIyDb29N7CFidJGzYcnNwd8U9o6vyyr918f9xTxWn/ZRsF
ga0wUYiBfQ3Jk7fjYkbDDdN/4lSnHL0bUrSlqGtQL3P8hpBf7slIxkrPe1cESe9r
gDPdI+cGE6n3IWJy9rgzk1ORchPnnwDCsbbAcXUuE3sF3DoKuExXKqzmXGZcOVXF
doxyoHj/0KJo5iEYoD691nyDxR0S9bSVCTjo1BAqew/UVeGdbZqv3XC3R1PNUywZ
0zAdRZcPSwdZAMnoP8McoQec1fKOxYjgBIKE48DpU/DRoZv+dBz0QLUKvkDT4A5m
hzrk/tqZEWb1s3OI0iBGyd66IQchLAXL9lTsMDJfTkhzQtU99AzirOinF5e2KFJn
GnxXdu3IeRTcpfXPrxRL4wmCJisVyjuvqQhAJSkgzkr3vLgwgeumUm95yMtsvtMd
3nDcqezTnJlXZpHWxiv2AZxM0dy4pwkKhWhDYzk0L+BBsBEUWG5aft6FtIFUClp8
W7zhwotZlQDYGFUrUAgdAzlDuxBqngIVyJYc9jlyhMcQxEg7yjhgkhNQgYLcsJMq
jDoz+erw5RxaPo4uq7nMp6yd3xNShBUh/DdqU6AlqNZHCyn8MAuxsk3jVuGW7cM+
Xoig0FteeJqsonRE6jgTI3a9tegmYqXeH7hf8wO3X2vz5KsvXqb+nFaIo/e2drOD
YWfv+9nlvKaGevl/toEajvAET4Pf86U+ABV582BVoXSg4/Y7rKUWWCNiu+pri+gr
8n0ayIY4KbhyAGvjb9qxBZxUlPKiYLbIbIgOlXzbyyj3J3dlF7TMJpbqp5cXVI2v
01FnmktNNcZH5GWLW4v8CRGvCAGjBUM0p4Dub/XFbLgOc9Oyl76+PHf0msJYxdAR
s0Lhu47wElW9wJB/k8ioSw7A/LZJMK+RaviEESCdZHTEsjNj+ZtmAUFkpoLfISpV
t4+UHxrsBxJLiP2b+JaRi1qLSphCwa2FAyP8HFKf72NYV4h8/IrIuXogZT4n3VLl
gZN/7hS1WmM/9rNa0wZ6xctd2z4r2lQZZR+79x02XyCm9AjT3exwBJKF36Ls1Zuc
zMb6SjcE3AihmsWkfwtfA7eWp2PrLJiBbSVVA5axYJIiTPAi6lX5ow68lqbCYXmz
FUIVs2a9rlAp3px0X1GDGCgNPRQrjZOOYFe9eKqMJn4AqBqoRsDt8f2a8/WwdPUc
cdJVQuNcg6RY8BidtDi8J1T0RGSfg8gI5o6veDobTJkRS/RaxGss3a3AFb/AaqIe
OuF4pQ8krtV9ccudCoogRvWscrtBljUUtXPid76pNFmfU/dxIp+8tq6ExrK0dqUN
3TbKE5av+mj+cvQ0xY+lCwXGVSi2MqW5s4U/VpTtVgaoo6sp1Yd4fXjG9us6dQ34
j+OyUY+irIJlcIyWJloSZjcsdrGDzTFRbWPOes7UM9u/x+NJna2KSeeLvgJ304jr
WS2kHSbsuZygPbdwkVq9zCbSe4YU+eK22UJ6RyznPuwPs7mgthVgZY/XIqcBHhfE
vy2ADydqkK2HX/f5NHLaIURTtkpXsFk8zAn8FCbS1yVE3a7NWTydY/Wc2b8s+e4+
CB/kwAsx5YgRO92radWIbRNaV7Q0FtQtZTstlSr6Jus/ikTt+evFbPBMx10+Fqyz
sj9wbxZpxIWeGfE0ox4w/RCXTnRFCpTpBoUDcmn0kmgvj/BIvkeJ0NDf2DIAaGdh
r87w7RzhBfe8EcgmatpMnCmFxnERrGPsZk/2Yhk8UjNOKaqdwxlh3CeK1RN6kZ93
Tvoqi/9ROKHKR9hd7OCW0Me8MvV9+Fau9KtQOpnaGe8DxSI4ouairqTOsrtG8Hsv
bdTXIPNNm6CS5X60exmNO7ddsIHCVRBNTYTTVkz83uAyMBSjtPmts/2xQXE29v8Q
U1y3S6qF9lj9v/IOnlybRbZrFu5aHvIXRzJV5oMFyYqQvDEFcEiFpsFomYOrXuT+
CzM6CkkoZ6ZcrAZ08xk96V27/nBJxTdMpM5PVVNz5yVa/jaV3ThJ+vAOjcmM/u7y
XbiTqcWZP/cCY8iKufwtfosrDz7tMRD5Uv3wsuOabDWNaSkZO+y/ZHd04l/j9mSC
qv6NY6AK2Wq8Gd9ix2zqBvg+3SzoDf37V+CNR+jrqQKWkZ37V866jAOs+QCZtHNJ
LplrTrog04gydVVUlUTOZK1bwC564IhwGRv89xRwYljImDOIRXih8PIiozyP/2rI
fDrLQp0ZwQeFNQMfED1mbfMDqs3TRaeeNV7+txAye0q9o78zc95ZMbSC47qGaxV9
7qTCrk6Tc0We9fIIH7K/wNdo9X3o6NLZlTuxmroru3a/rdpQ9ofwYkO2OCnkzAE0
XVacIRR1XY+pURdxYp/tHK7xNJ9otaQ9xXi89YgCPTDZD/F1fYm2/RsWp50NXkU8
OdXjNZXQTTe7UGEFHFcxQSVSnbcxAuqVPxQo1gcZsE4jTQ0Xr6f/WIpSSOncx20+
mZjd1FJVvTpNMCHS46417ewpk1JCaP1/zNJpjJrYBvdtSsfaORPaohwOgH0xL/GS
DSQnZVr6CBUUuB0GEB7OpPJgUxHnBk3NjZyRjpBeU/rWQUFb1KWmeCs/T2nW0e1/
aKNMS5FL2qtnPCe4MrCuKlBmYhQ8TQ/ZvApjQrjJ42yPODltlUvqezLjggwY8BFs
Ei5DCnI/V+NsBVUhnv9UYWmDT0iEogu+XGUBlwQYpDhhmyOzDU/IlLVOTcDwB7V+
gkTEgrNrjp6YRraScJtkxjbzQRok+112cjRoVIS2XgoN7zjWQ80AObSRolyRKvLm
dOMSrJDMprhs1/CdAHmYZrfdx/muAdmBgk8APwFeYF2jt/HSZxLMh1rCUyVJnmf9
eJJM9TEFpOHE7Y47SQrc/MfgMkK8AIZAWZufoH1KzblNpatSot3zbuNAbtmkagB6
QZ5NpA09/g9DtMp69JvDDTYewoAJ5wNPX9HtyGzpUkDkRuEbWtdiz14dnwGmJ3+4
8QXrHL9gTtMxq+NjYAK2q8onXVCVHqlaKcCr1s3evZujltDt28AYArO8rEwLsBt1
hVfuk3dwy8u2TLHj43HKdIXFHsSuNH+Vc8bh9GzhwGev7stVXBw3/s4aHuO1yJCQ
ZHoDlNPa3/BC0BbNmrbp8F4lOCaLy49RCBcXc8kqYNgsECmCQo06ZcJh4BTkJYQz
fJyYTueHmFpoFsUI6cscHx+a/z2MCM9n0LQ3SxredkG/6HJEMcogBqpMuHtZQzNM
Ovy8JkVTV6No/fxGcebtDFLGAMOMsq843G65gYe+dXWM/ZKbpbFioqou2aTgDgi9
TTJTZsagjh61OSiH8B/4o8aiexFbjl/iHM6TgwaTeIeHtqMg9AxBViW0jLFYwwA6
URb20rfPkGRQeKN7Qql79Oc5njhq1p4oIRErba+cVp+EhZDVlkAz2S6F3F+v1fyx
BwyDUtaDqzw2oVs3xV1Izwkrd6/03hLYs3CDTj/k/KMyTfLVFVsHPKfih/NOg3Z+
cW0PjOO5RQ+7z9YGQh9Ueava5aGyHyYouRCgLaW/IqhhLMO6lXCxsHwWuJIIir7C
kteQ14yjVbN5x0ElGc8910kPMsTEVw4i5KeC9MaYH7z0YW5ZfhMymZ1GbUeyiXfv
DhpRreCcSWkf++UTN0J0xxEePcE2Gbpq8LZi8/sZhKHAwiG+j0lVNva04JgJ3e+R
qVaIDgk1cs3r6q+Eajlmj0DLb5lORTXuxACOjhsacu+N/JrbqWE1cKNtEi6o0drL
b2SF6ywVn/Ra62VhvGDXAKGscI534kVxy91mp6oEQaejMpQxIaf2yX1zVyslyCX7
r5vwzUT4pv2TpSNTZol8GcssRx30l/NM+qnsMi27q1KM2Aow5FPLsLiwgChqEOWf
4ES9LVDH8pYB+S44h8Y9oBFbu2GIBUO8b6M/zk1N7lp8BqzgbG8AqPNHvXxZ2Hn0
bvkzOIfxfwyYRjwYQWo/Cnk39GkNcDlhnjBz5H5EMskfbcxPlBbbWdIJGDjH2I4x
08WFmKbDZnmJMPDIXrl2JlVFLFTpxWqA1wKGm/7IxRfkPY93PrkacF7fy6J7EtC0
KZhCOhBJyHSwv+vruYLUoon3bOsVdH3lSJ176JBsAX6asf7qhG4+cWNXmyNgpjxv
2wMV10BpS1Ljys+O6my2XCbkgJtHwJtxyzJsH1z3vdD3A5EHlnV647e7/1Qc+99v
BNoo0GJF6eplD+Iql58ZySBuPBo/gj4jdpPd2293g1/G5AzrVowVdzr2p67eQqzz
tPU0gFZfcdrsl5H5G7I0JSfVu0Q0JDnsvBQcRWbxsuZpVc2Cs3LetCX74psHlfJW
+MupYQP5d8AXnoqaj2f0r+fS2K5lo7Fj9iTBpDTd/oUGliUrf8TD9NH5zKYatalq
l4gFh8SEnZEB++W6FYF05UDsSk52B45OSWyf7WzTorRw94B8pklGvwcMe6vz+VzW
pG/ToLysPbRSWAoxJz5ide1RNZb+3gyn4XhypJoIhrT1sVQbE2dl1TOtnS7tpAX6
FA7nde8O4l9jk1VcV/V8fjw28IA3aX+Yg3MggM3gU0bKBKETvXzyOZ5AUImYNJkx
MihFd13Xp7iXrqrFqb3FHWBZsLREPGUgmSQekipUPzAwgtT4rsyI0kujjDG8mY+U
B/n5REVbjsp+mSRN0IcUf8s2oXwkuz/6QfU+t3Hep9lz4e3YI4Sy0qiFMh/1Vzta
jcXejuRj1fBklqJEZq4pmUcOWdN52KsOYdnPtWn7x8xBWZzcvrH9ar9jOSykIExy
dDYaPVR1GqslR8WFrOOH+EYKQkBDT0kKW6A8FEy7GfcZYDO3p9Sj8gnaipuP9w4I
dEQNSZAbkJGQfja6jK5RdpVCfmSTkLKtQCq/vbE+AQhPTYe4r4DgNnJ3hFtNwreB
/I8da1vMJySUBCvtIicurwJZQHVNULRonWf4Eu2YGOnRTU9IDfi6dVezRnLE47Sk
+duOZwhJludeOh9pLwHS9v7DzDalnOw5fApCqL6V9l87kE16xpFOskcAySSQufK1
8ujW+YEM3BgCOlRy+7O/+uk0d2MndUL+hG/70/9OiEIuH/qaSBICCgUqvwnoNqW2
qLffgMz0Bw/OoDFdoa0taqRty/dfPUfM8GC7AZtPixC413d36WmOFoStXEeoXMO2
VMZOSB1OTArh/5I4cUhqIpkruwG/GXzQ64zBS39cr4060ogIf24XSl5XlU0uyWsx
28QavEHdHmn5p8iX4JzcmQmOBEFRA790fSZA1ge8YK1FhezJTPkDbIPq13siddZh
4gzPdLMTdWEiegIHNSaaaCwNzSgotqviyROi+iTLujZFfjVjMaXc48de5hfh9yaI
UG89omMiSkUqOIFC9IRri9XPZWpkk4cIT7x6xg0Wvm2SH/aKJhnKLTKNeuqpLSK+
MIqYdSIIMQYANSz2Xc7hdQizYZzexBt8Y7d3xdoiINexGRZEAdaDPtf+XG58eYE3
HZVqWdGNddLf/GR0rSjyasOUhX8TY+at8//WIYdVfaak1djzbxrbB9KNj+YKSOT2
xYnM9UHX7GmeM7c21BWsHsWV54Rb1kg4UOIVK4TR5GXPulMUdKxjdKZfSHUs0JCq
xIOEHOEjnhXfbqXbez+TGYGA0FOzmCtIS9GPxUlHCyUnUPrL0Sqp+CUcXIJWq4fi
Du+NTmxZsolZLfT9CmIZpJ1lRlv/ikQ7v68KH2Hffuh09UtTJ4U57CZASvVbeLt9
zEqG7DYmXXzSPo0cULgg8dT2jJq7VdIsjf3eDbwYLSdAeoRTwisQ/UnMwE4cqGzc
eWLPUghVG9SjyGkPF/JteaYhMQ8M7bp8XAjUfsbJFtu42QEOfS1wctdmkaQwSvfR
JSWmwd6hERrLhqel2BIIjBcTBD5J8MejTDoQkY49dchSncxb+4QrRB+hL7XmBQRN
RAYalta3eZe4VWEjKGXLx2VDqFGa13wUpXNMNdvs2WlnJm63FZVgpYwAIdd56VYj
yrQwvfqjUyM9Pss0okYHJIh03m/+hkBEnELFGAwnGOUj4NnARYK63TKBN4rrvMoc
Nzww8ikXdxTas07mF42EAm+ur9HDI739/wGq/qVszd59z0S2OLV71+hsFlp+mnoP
9X/jAwPMUb6/MPFFMTtAv7cklDi1TmXkN5tAty4waeJ+/Z7dCrQdPWtv04Thb9MF
tQTnrlMvAYKWnTAoaLY83qzNv4XwM1lyvrH5n30yoRezta4gpiReZpZQLe5cdjpT
VcKB3PlDw981tdwscXLPGt7QmvpuwyxiDUm/37HwtYoWwG9FUUDJ/JurupWvvji0
u3qyNqjJFwM5sAllMvS8mJtZzSz6LQh5/S5E8+ygwCn5FvWKUw4IY0Yy1pFMnwxt
f6h7i+V4hwcQfN+lOf9b2frLjDa8WuIg8lkO+qr+WEmeR3sav0hGPksthFLVr03a
HYbGr2hzAvmW5bO/Otc/f7A2s9wddPNKjKI6Eb4I3XA2nHC20uy2LXGiggloUojW
C93JPHA5O9DKBAutC+3BkhcywsIGylDjr/O/mwMG1AR2VDLX5llorFXA4p8QI6dP
YoGNxS2CZBEANDGjrgxw0EZ8TWlJuyH4+DLiIkvoYZPgHbP6qHxdRyFCEOBHUAsX
dnTFoyQUVO0xmC3TX0d34h4P7SUqfQ/On2VOUFEjyp6SeIOXVqRuTw1GOGlTGVD9
a+xD8uAM1W/fKZn9UvBh5D/qsD+sUVMOzMKBx6KNPFwd4+8JjfSBcYgXhT8GxUkn
V/oGiPuoT9EdFH10Avg52SrJ5LgrAwfwXNigrgye5zMPdX1mhTpPqvKAn64hppcb
WKMX97bpp6G7VBDpPGZg6Xsh+qTyxZcwEvSNxhd+LgRUfsfoLw7Chwqk2aXRLn4J
/Wt/Jm2hbiHMP/W9kx6r8pY5l5E3qS+K68kGbgK4X5rllUi4Je5wKc/sVjAeB7/m
jVu07sRWd3GwnRP9LQ+T7JB6UoMI3zoneThhrGHXmK5r1DHf3HcYeK1zYvlYEVXy
zipSqh1jTjic+cI1othjbRE9SZ9uOmndsd3dgza39W80PJeS/GZbaPaiq+5uftMU
J0OwZtRq1cB9uo2XO/Pp/SdoJ81WvnvNJv7Ype+EpguYI3f/oi1qB5pCgx5oFrOO
ByiaDtXlK6lmouTQYdT8nT9n6G0QBBQ8hW85XP9K14O7Gz0edAbBoz8k2SezHA+S
4uc6prMzJReqAl32uHnP8Jn7GiH33taw37BXEjMRuJvXHMKocNgD6LSH48AjnYI+
S+AFOApLrTqniMB8onc/71mYe7QP27yVHDg4fSbbpSzQ3/JWWoKhGeTFPEkK+VKi
pv6jFhnvySmg2SkdtbkGrpak7km+D3DFmgqyLxkL0HRacJXCbtvchg7U1bT1ax+0
HOiuCefcEBUC1ZVF9Sowo2siWGEkz6Htu+pxw9x4itIWqKdeZlp3Veqz5GSg/LHS
Lf0+d4H8UMze1YMQjfqmDVeQ7NKKk9YnyMK46QhbfmZppSG2/lxnwt7d3ZN0NaK+
ZxibV8O41oP/BmWlZhGtf0v3SgnBJkA2w68Jkk7e2oGnqq4LBOpJCaHp/C6EJybJ
NiWbcSfhMsx7WABl3eFb2JJmmoI7aL4f3JFCU73W8XnLvsOVvx+YxJh5wMACDfkZ
SQUDlRjseThfxQXyO7pksGHuRSf/TkCIyXWyIwm12/A84wgaoghM+rn0rZNybTWx
G7Zk2dFzVZCAHU6aFOmkiBOChJQI1NAMNpo8P0Mmmoa/lbZjyu6hDDD1cN5LETR8
M/eMhytehveiqsiv1U+Aj+ZFh1ywfbh1Y3m0XrHoh8Y34YYYQ47+dRIET9l7htT4
RP2JTWIfI5eHw8PD+hBEY4jDo0YBWlsAEW8gN5ISqav2ttbdfWsTfw7+gWSTAbHp
GdRUuYV2mik2AeRUeB4jUHb2XDAltVws0hylt8ca6BJs0GClqhXL1P7Z8Q0O9+15
6J+7xKGPM4wWt0CtY0m8A+ZnVZqeUAx1T+F1RXcMmPiTJhLHTflMVxkdGh7M6ESC
5c5Na2QB4xRDrvl/dziSo7rrvPmlsE0DVoJt9FbwbnWPoVKcPvhHbyO8gkE3aa4C
DaDGoP+juV714AjZqSJDetkYSVRNk+5KZVFGox+kWWTL/i2CG5b5tcpdxSezz4DV
VQ2sMbOuj/PCKkQ2GeQZ+ks8c2Om+ZxFEqqwKdCHYjh2VmJsd1wtVMY7gfSbq114
0t2IvlCVgdA+EpFHTKHQxOKlHHA5mE55S5ox2RQEbET1LfeTETzek8ZFMgczSfwW
uJFlJhC0tP5hI6g0lKuem4IidGfsE6UyVmhINuAZcXIqn0vC3m58hvQ8ccR8fGM9
u4m+GE97Tk41KMjKQfg0Tcj1SLsaSGOZvfQszgjj1HOukAWNape4sImQpOmIJf4V
5iP5H07tx9lO8R8QXybuTV3uVWPFc3i4lUb80Tj4UvOLCcEtEgqaHnCR8uejSSsw
q7otQEb5LlOmHxpRvtTdILjed9iJbOtB7j5ugsKZAGZ1EsI8Hs9xLTSofgYk1m6m
Tp7Coi8gh5r7CY733h0jy8avciD7zTJrvfDnUhuyAKVfMDW73B9gVSYhTjW+igN7
4wHp9iLGT6YrdLYbhur9U7THdOGa68VZhEPUKyMyfAwxfZYXANW1N9eSGJXtbnD0
wiUZqxxeTcJ3d+OOhyXlDQDrRlMMzI6nzgtCWeIyKU4SbLttxYFHyz8KA+0sgA3j
euz8e+8bz7DCka6Y+CIGqwae/U8xvQMMwOB8sAy9HbMUVnzcwnIw+DwGvSkPrvmD
xyEHFVrKbCJojLfE2YcRRJusQmb0NyjumeDotHc/4B9VIMaIpXos9VdONvX3fF9P
ALJ8SKngI0lHxpfOPCUeDPVZjK0+GaivUlDbljtHjVLDjqtlhOVOC0Mhf9gcvTby
0y8IrsTp2Udak/I65atPIh1GfPQlfPTeJn6BgoMJWbsmOO/kDxjUMsYJZdg6wjc1
F00Q0pzuuBBmpibbK2GREY/qP4twpD/novi0mPQmXYfKNv3WhmCNbvcDqR4GQ/Bu
xkmvJ+slIj8ylkqqUhKrajofOjoELt6yfpQtWBprjXOp1uNKIO9/WNcAX/1cFRuh
jW5neaK7roqsaT3F7R3mZFjEddBGfFlT0hikXEFXC58Y6kWk+qlYOQpqpMa+adnd
+Np7h/m8w29letSAZ8FTyVVDD2B3LC4JHTWncYP9bZUAkmkk1KXmS9jvo523VPA9
pYns/AHrtj+s6lVHiIoFzx5GaTh5pU+TJ8VjXqtZQtDzPXwg8uTKkZQf104S3pye
TVEpbBEhe3NOkYEAF6ZIi+nHYZCZJyASMX554xP3f2cI4oiwehTfJ34Jxuxb7wwA
xIifoVNszPyStOxfaI4FgQDRDRofj7yB+L2o3G5syNpcy12GiDPhnZ9K/M5eqpXL
YeUp0LUAtS0otIiSxix5imQAX5xzdRxjdE4Jy4vhwPJ5APFmP3Z0zIlAVbtxwDRV
QKOZZ6+dyc0bi+HKICQRfCBnT8VZwHZrl8z6iGuZNOW5VynnHzrbXF7KfwH7mHTJ
xGN4d/CP3oTqWdVNGRXV/avsmlE0vPdWoqB0L7Cl5aIMZ58F9R72pLKvRqiszfUi
Wls/6XNLPePGGPllQBD8U0eQyWNhHE/Vww94OlyN+ZbCVdZI1CdxwGPY8zas2UXy
hf8qrk1BGcy1DpBATtGAoH4QcOZIS/YPtzMsi74WtFFhO2iC0CYbckq+Pu6qPtHG
vFQMfeCEMRi0AUdj0XG7JtJCgYHN0dozh+pf8vw7zFa8KxfuXf8pntkQXlqAPcVb
koegR7wJ29db6Xjmb/h4blj5Sv1h4VAOAEcs5o1owsNJrkHO7lJjVHGR5EzqBHaP
X25PHqV465ModndOV/TvLBt6TJPMrfzdtaY7hrlxvhMP4QSTmM7iP5CSIvGreKQ5
5ROs9ru/5xaS6xFuVRdckd6CBFS8L/rVGUd1OmQqczw3mJirpN+vW2CDoxlEnwWH
OjEQyClFAniS2LKAAXzCHTrdn3WZcs90Z7eihBWLG31s2coDKWXNHd22n1GCGoB0
oZNLK5qkdy2Ps+HnNKHGv7zU+RueSSWVtxa4WsmN+sRZSs3HC5D9WWtwamuT6IO7
XZKT4nCqfpARcjANZXDm8hTaR8EbH8LSSooln57+yVrLE11M48EVyJc/90t+Q5ko
S39/QLQm7JRdaUMAaQhzVT9lyXRrxFgbsVjnS9Y90kF04YSB05PHw5yx5jR6dY4F
ofIxkCVpvYxyTKdag3uUGACtBhGCbBE/GMXTXAP3EokZTlV776NSVG3eAec+ti9k
D/O+Kt6p0QUVP3FZCkejJuzqO1xmwb8R1jrfRbcT7WWo2hh8zmWGRd46g9ANWKnX
huyvZywE3w1iB3UT4H8ao79s9nOthArtNtjAIgeBOzuRx4IpY7InmgnO4yHe04S/
Tgun5NU4rOuTGoxiDRUAanRwO36ivCxWyAkGTiw704P/p0nIqWlEgBqIBF0Jt8TG
27l4SNIE0ZtppPEAdihqe3xCsKEKehEH0DxHqzPEvmAs34AyrzlY2xWYqdG14qMs
QLATngMxT1zXifRSJ0DStIFJh5weANHcFZD1PAcc0vCwma0nzBVMR2oyVo+oa6Zh
Mr5222qog16dp5g12WnhcPjp8tmir5dzKV6xiPweDd4kU8KlVxA+dN8qQHU5RDSM
VIS5IJtGMKKBWNxsZe+3V+3AuPxnMeMIsET5liQViHnOcOBMNtf+dTU3a11DMrxv
ms+ZJBilK0UdHFJ6N+6+1BA3r5/YtgDFTHb7m3ogOD49Mrrw5tvrNvOX0unxjjD5
auS/DundpbgR8no4omTWA1IeVxVEkTl9PxOUnq4LP4gRfPYRQ7Fkq8VA8rfq7t+N
SaFBGSAj3bOgWKqFXygPyOvCDyNVLMrNiq+0raUK38j+a8ZcB/q6OksEMa/QFG2H
ZLS3flQdJ7AUKdXWWrhymjK2ls6vdHx8/beECG1sXLi1vc23pbozAleNHkbYXFe0
OfnKGmPoQZkH++uJ3FltTeSFZ6uB/X2WmJaznecvUkEY2B5XyiUsfIdZlBuoGNGF
JM4wD8KQqOYYJfcbcwU3k84ANzEy/DPuvt82w56JSC7LRmqEJKIHLQ5KSAato0YW
03QGgOstINcR2KcXFu426frjophk6g3yJY8p5jum3QLzZiOiX2+CRAIwtxaRH2w5
FDJ7/QaEBdj/X30vYvKWNMdmamJJY+kSIpuOPF9xXMna3Ix9aLff8qUCTb0MkE3c
SgEKU+GSluY99L4zfRGJ09QVbzMTAX9rP2HgDn89sFHmY5oET3fHXznT17S0ePWT
C1pK0wNha7LKGtOyzSlwlVwsgR0mZZY9tNyQKoMC/OHXv47eank9aPIA1tc5Eh/8
ZP/IbfVj/wGhSOGSAqe1mkL7KNt0M7QI4fNU/sXw+GSnUeYN8U60D+R2W6cceFEb
md29ZFjjpiYjfRE3NYSObxPLHA9BCQ5alqEJpSyNFWopjLd+aynmiagPHnvMYMe5
M/fs9lJR9bOh+pMvqPrTvy8cJBfUUfHscshWfRUOEQ8yrLNyh6nq7Xs/dQa7lSeJ
AeQwPeVFBD9fhqct/idga+r15StOhjr4eZEkrPe80ijAT6HTVkYoL8nKjMejxQGw
UdSgjpGhgfE8a2PZlgmI6eQRhrLkXagr3KncKMb3fD48qmVd51Le3Aw9OPvk0EbL
cUIBBA2cId6oMdCN+lzOijBU8qXzVTv4uWNPdltavG2Uq5yYOOo1vtKqspZMUkgh
ZFZAOA6Gx5l5niHDF60+aDImgn1P6gvzIFV2ZZ3JWJpvf7iove1twI2emfw+WBJw
kW7kwlmQ42hQxkRWLqw9N3+L6jXWAYFe+WjLsEdIUiPb9qUPm52JmeqZvXDBq6/j
ag2HJYTul8H8Z0i8XaTjSinAHqW2WrD6AXClqmiYr1CMWZouxIl1od4yUHwTru2y
fbQCxkESfmXoPF8gsPJDt4PJTMLt7larRu7MCDGcQGfDCBmI+U5ZGzdMrtLA8M8s
ShnM9g3M8ISUpXOQH5sluBMEFDMpcOXo1UPXj2sfHtfVLftWy/Y1lojEoL6HT9Y9
VuDLBIVwJC0wOO8QPuGfMLvwKKUm1FSCJbyHSxiBRTZlmUuKUn6L5Fi5jc5jcC95
cz+LrmyD36uFXNAZ1jomZ7kWETgu0ePL2JX8VLkZBL3Xte11ZmTkUF/d7TBt5CMG
RnP1vug4toKBzFu3mG2mk9t5Fidae/8IdBajflBAau7mlDDDqcrn+WPlHZaMQ5jM
/bdbpHs2MkERujHqZ2WdMiTh4GgdukwFAUdUQFAQNqgHdOGSmqrVyqsDHqXix9Jo
HJp5OtZvYWwjN4j1/Kx/FnbRcO42LlUMgcEUBO15kS785qWE3owfwYcZexPB88Wx
gHxGOhKVUXPc7IftZc1JdyQgcTLzYCfab785c9fmIK15TSabSVOV7hnIRzBclah1
+7eeMZO+fycMZP47lijeYlXUeRLOGV9PXLdhtWRWllxdD87Qgb4M2U3FKrv+GFrf
JX3miJn88IVZAF+O1ykTxtppg5ALkAdq8o8EG+OAM2dqeltDyA5Xtyf4Msa1Z3nM
btslW12D8qniFqB1PidzKgdto3igZEhHTTEdxN+7kciGT1Vr8DYAxGOttyzVRsxV
I1fwUZZim4ichO7xjrj8sjOoW4z2NOOPHLbnHM9SRxurc8eO5LABDa6Cyy9EX6jy
1qPq/pJ+afOSVYW3qSdnT1JjB4GksMHNyPwN64PPsxojIrQDcqnLOHTQuzMulr2B
A+FpoLpl0I8GsKrewvyJ79dXyHVtfXc0EyPJwpV5DtRQRvC/rJcWEM+s9YIkCLll
qkARkjsXmjVEhyV/jxpeluubVwjdqDWKhcO1NlQSMMzq2xkXslzi18BUVrWnaUR+
k1Ug19FJBrud8TOnIW9pOQWjCCMcXxOUp3k2Pi175ir9SwTibGfFKIUQ2/OtJYmT
xqqp1WZCjdiDuRWGUypSygbPGMKWpfiNWSxcW/EJh9s63Lg4oT6rVVNXnqdQqodD
XFD218OXZjtFW6Ffin6OCFCSXiINSMoO4/HmExpZnrB6pUzUXcoXIFeHNEk2SQBd
A+6LNA0c6jHzubOtMJUblZ6moN/jTx6tKXRU6aKIbHREIxoLhf9EDaQlKVrYaTCT
Tbs5BUmcaztbtiYmn4iHNumMBtYELRbd+UdaVN+/LdPQPVdYax4gN5ErDT3gH+10
wFA1MH/RZqabJjDdrXUG7PJPMmLGtsw6s+MA84AeQc6X59oLd9tQJ59XV5XkLFlE
olhtOZLAcKARrPKJfuq/hacI3vF56OViFXQTrh4sH5vkukirn4pGf+2Vg2tVZj32
d93B9/4jMlzZ6Tu8xVPSkj8NXIoFf5bTdcfTRDFilT5grXBg1vVHQWLROpeXKSmv
RaGkLP12dq+dN55DU6rF+Hgv+yFzHF6gyzYVRDGWL4s4i/0JBYpz4vRhCH6p4x+2
PvQaI2vzLPf0DTCBF0jlAt2oW0z/Jo6Y3cfNGiqbURf0+zA6P4drHw6XsMyjHZA4
xEpd+0XsUrCVjkLYLC6dkV14InTbgLCVgtd/iWRQDqmIomlmPy9b/uXA2uVfWmYB
BlgNXbgPN5YS6hQca+i7AEmKFHrgpoCwFjfszbZNPgOdAGr14h0v6ngOAWZoHrXi
UU0+O6XO6zgK3SLngTTr54YSJ/XRwUvp/4f3yKdkjr0jvLIqPRAmWA/H1/7qx7xb
6VanX5ULhEu8bzlTGJPXZ7QCS1/utMLVdGqc0/r8GoBApuDUkJ48wonGQoRHpsPu
S2c5P1gLalH967oECBAg904zBBU2lfZLcAHYOnyYkaNazTwnj0H2O6tlAuMfra2X
FNpiF+ukP6+9J7NuUIiqczY6jbmZqoOBjjq0XJ0L4PGhsMScK+DzUrLfMYsoAMyo
eMmzDqnPcxlRDE0MFUVAcmu4uv44OBtNg3vZsjc9/724ltQ+5/Dtszvtqe6bJt5w
ouquD0VHHm57l95J4j3b0a1uAE+C8ra8BbWxYE/nEgTOiE1KJYhu5/ROrgi1K6Ac
efBp1g5otyJlq+kaLZUFQYhG4hCVDi0GdKRU8CRJI5csNHsH0ne20jRGTvK4HeD/
AgaDBIEtbATDl1HRKYvHyk1b+YKmFA1+JvSfspzT/U3fyhJomz2T2+Ab32MWu5ib
uGOSU9Z8jstXyDaDVBFLFjSfRI3nbHkGvcNot5dIJGHvWD+RIzFFWDio1XMl/4RL
pXaGS7h+ZxDxCom004cK/yGQNXNULG0w1auypajs9aV4v0zqhAu1k0WlyRXb/1So
bRssEUSnm1m/NO0IxlwN+8btesiMIxvq8uFAqgj6edW9JmNSVhdM1O2x9LWPtRRw
6RKs0HgyfyGbJZUjynWkz3B1n9J3HU28ZMQIbpU3GvBlPHP2a2V6fizn/717qlmN
cQr7z65klN4la+PpHt4bhtZEy0trLdcowZ/5BG6JSO/1AOcQ7sObFWneR/xoKcFF
7ro47rTmBxCD01eXOhGsO0qkHdpW543GndshultqzKW0z9VMC+QfJrpVdUOMw02D
LUd233DvZ93lvlOxhLcC8AU4rs8P0jtpj3alaAo3cRwhZk8MBhSnebz71E2AcPHo
5cvMDl/Ib9CNztie50S92Gt1wseIfhYH1MWtJLkHomqI9V2ZrfCCHsGv1k1ZuD/P
XhnEjXClr/3SueO1MbGc/blcKY9EHXL2fEPVaN5qDmUh0BSaqN7jEVTjVNk9xuG7
t4NJt9zpBHLVLuDnfieVKHTGj/ebpfMTg8Hybhp515Ov0OFCuiloI4nS8fi1Fu+x
lVDvoj98wL7sMVyWn0K2+ARI4lxJps4Yd/kaqP9z4dXa0Fl9WR44t9Y7pULWKmhP
hoOBHx6zaEIZe4XXKC7Os6ZkfQpoXOF7RJT1V9SX807PAwmY2NksqNZqG6Iu8VEU
Oum2EQytHkTBjNWVuxS3vC3Stc1pIzyqO/7I9KlyrCwR7Ujm4keVvLZcGshyAYA0
aWOCudhuf4eVX+sbrBuLTAVv/QU/evGGKpcTAcChYDNM587m3eovGeF8mK55YKne
dGv/cPxbqLhIBhkgSbdLkuCH5//zDvb+AcRtiot5nUeSy8VWeMlu8R4p7yklHm+X
sOw6DymkiHpPAtWoXf5WZjehQb0pUX8bEid9wrcQYz917TMopxpfBU7l/8w3GBz0
Abq4c1GksJkFJmAazObD2ViBIFoV6L0kqJi70uC/+k8Xew3AHe64G8giJxnnP8MG
abCoS+ZpGHCKg56R6XD38eEG5OOvkLDNULi+ZWr9PcvLi+FUDRZxYET8TX+SZHhc
8dFYvKMgbTo20fa5WaHQ+qWlFbnnCbt3tLmqDUTglq5XBUP8/HOreW0hWYCIwI63
b6k/VchceMPaw3f7etmpwQcE05nY6U+sHAnOvLXYf9zuxWqfQP+HigeWTvVvs5IP
ZUedEciPudo06VYuEldaFXCGCZohM3+DVYgU1TuE0WiKDZqTm+9vrdg0I79PlcIB
/uUwaBGQbzYcMOmtiRWraiEzetgV4AQ8v+2OisZRthwU3p+5/z5oq+xRPa74M2Bt
XFy30DjRZPg1pw4dC/P5yIMhPogHRgaygdGGEG2EVkV5MH/XqmjWYpe0+AMEoGDv
rD6tuL/c1tUaWW/IzJNYdMtRjNy+ZCOGDUl4wxKCnpOuAvq7BOlMQvvw12vlueuJ
wlNWP2EzfeV2V5h56+VpR2ijTR07bj/dTS0dK3Cu6xv6BOeSM+ChbkPqa9De9F16
omyxUDqXzlkZMBuwUjbXXmXMRecxGQaqj4ZZFCEMP8u81LfjK8hD6Gm3aVGu9Do8
BAoqwUSczeNm+0zPZAhvmI7gLWrRw8pnMLRhKuKrG29qmVk2qzvIICPX7E5OJcVL
o30+o8Xvw8OkCnF6xjoEuh3X55/EptYqvrR7H9HNDXf7BuF8BWHb1si/Mh9/ShH9
6BeJrgFHRnuy3QNqimGEpgjJjPbKHvixAv1EtsuJ8iV77uHuLTkJcaPZzP4ImlXi
AFh2UjvbHu73wSw8dLVYv6r4ei5aSHnLoehuMTelKF6cLQgIhpBtNAe3Z7zzP4hb
Wp0/TGo+ETMHVFGhjPuiICXlX4PClH/uvkkpCGhW5qqTYudnAx6uinvw7mKnqN98
OTufZNbjbLb4ZgJ77+7My/pQtKmO/HurzXHef6oAYxLg5SsNiPfjM3S427ZM5NXe
39OUCyG3McrDtjCGqfA/Pm43ogSHlllZgwLcPDkqliH/PNilGRDap8MVFtOS0xQd
O1D+9GRFLlHd9m+IkVgVhFOKdm6JvKUxaDmiCeqxRM5b0cJuzKJR9+sy1gRwqsX5
r2GMEmKugd0StCfV6WVepz8ibuNCPfI3Kl1smE8Bt3/7IntAoWEpoSDWr0KLz+mG
LohKOGmXn5x8aW5TE6vcbPT4rMy1PafvQk2SoKxGQCFzkbTpcADNBIzKqerMXowu
fqwkzKWDEzSEcEeLLv3+2EP0qx3e1N1LIxrEGJ9l1xxCZBh2boXcoJfhzo1nATqF
3J4wBfG06ZJvbEM4s9wAo3hAhjUa1hC1Kwc0Rw0vpaMhUTH438hrzDT6YRSixxf4
oPFmX4RP6k83C3sF5kp/PXOv61kB3BkpH9jxv6F2HehhIb1qA7FLY3F2QZVcCXln
VjmBR+/YqnGYDyV3r4uzojFv0GDvVFEiSxiTPIA74QAfoapteej8PXAt7WzrzLsC
6e5didIuHF6XnQ12V5VDajInlWW5EO+PHWS/7LK1m1FdyzNwQaEDKhounHPhHJai
u4FTyuAQ0YpmscrQ/uVdUtQ+okZEkkc5btdnjPS2v1JT66LU4KQPehp9MJPcNmFN
Pk7FiFCuAVhnZH6hnxmEI9B3zszoULXQrFTjbq+bIuXN+fjspY2P5siDHMQWAadA
sBUjwTuQp8sdavCFH/dMQZBVYieeWT04B32QHQZZxwupqnDAT5a/wYmfQbVUpdnx
/zUOhF8IkvukUNUqkIhZrJYrxazQ78/ZzV49L0UfN4LCkD2xPZzwVw3poAKzZImC
Zv60xLhJg3n6AagLfvS+w81OasfC0B7xpPZoLWTzkj1KuGg4HATMAzaj17AFNZQ6
Uafc1UVedKitExY9Jcsp9+wDkDp/qmF/XUSMUeV95yJXv7QviatjzDmQi2kAhV+K
BZ71wU5SZQ07DhhG6T7L4wv7RqY1401+au3i9MEormKSEi1PkN9B7javRRXPy0N0
BosW/FIOg6Z5KE86eTK2dSPgS3WrGKQrEtq3e1vA+AM37b/g3hCz8VAzYcmPjRSj
aoSqbJVmm0vSXoFoEjLj//j/KlloqNKOR5aQik2Ms3JC7XD7hAhdOzVvllOHpCL9
tT2t7gSzGatykuYpvhyKnMevcASTjZsu45HsEF74Nv7rjqgNZ2qN4txLDhlw1Oja
qrx/xN4aMZLBb4LAOGItIOLRFlFJTpimGRVMf6Vmr+Z/4c99SPaH0jBqHUyXHWVA
o3/d+xbz2k7CSdbQsN9snkXCQ0ZHqakb0pdT1gYIuipp5Yibl0jGDT1XsXsPci/o
r7VWwCH5fOP0Tk7rIuvk3aO8+l/08iJicMj9NqvfpFezxeoHt9KTtv0yoXUqS1OP
F+XxPpWOQWaWFe9RxATFH/U3+I9dH/XJqLxiNo6Kqh/mokTCu5W+wn8Ht5KFHFCa
J7qqzIJmmB65jdefjnJ5H+VZBTFLrKM9nGDkQj2XiWsrr6uYALuvKyR/pq6YNOa8
zzlH7e92V2iTJnfOo3+OVu6Km1invvIIAcnWmG05hbXHzU3H2FkgvDDiXaL7lHXz
tLltuwUyFtiEC6DbA2GKvZJ1KSduatQ6SOIDEDVwJwr3tFLY2LEmIk11j+00v+1d
RXcFwQu3NOOpKSn7i9CNacess4fjYYPD0ZsCP9O0Aufu6+fXHlUJrC6ZfodHvLtz
nGUPsBrlQqr9C7Icf5iNvuatLGJjtV8Pycn+1htlq7exVppL2GNzwDh+3E9/nOba
NObjd/QjpBfpnzLENFU5Iz6iJ5BjMI8lGl/m+qMy0fSTVupotwWaumajF1bbQTe2
IyFYcmM/9KBV1IYqcTC0GdGK/Gij1uqQWUlGgX5Ow9kGvfHwFrXvwWxZPN06inEW
2kMKKb2y2U3tS0ol3+1tLFpqVFgXd8nOn1QbIj7Fr4kfQT+xKTfhjlZO3Dhk23yB
WELAxKVIByk1oa7hjdYIqIbJjzayLNj3I6eZvEfteYA6uaqPO1SLicFdUYlev+68
CfvNBpTNkVDv/cxB7F2JsJ/iW1/sxz07jksGo8c0yZsmgZ9l7KzHvqzUG5sMyLYv
bk3BFH6nNjpqORxRu4Az9BD+IKv3xeS89JttkV61Cge6657tnF+zT74/GPf/Hs9/
O9hiCymJ6S5VFUrSUsHwbc5Cx2CcfMYk0pfZZ64evQBfVu8B6fy1cDdNXvbjjGwd
tbIYCvp6vd5JWtosjTWscebDBqo+dKaY+iim8Yj83LqPRpG0e64wBHkdnw04Wmxn
FxLpriY3IZb4NDHQw54d5dQA57Kjyrx4LLV+38efT3KH4XsiY4vGEtp4wJxBxQyy
HBKypoYbzFPDnMzOQYf6EA0RgX5PDYvQr5y9lViTXoIs8NsY4WRVnaWlH9pRKdjo
u4p2eaMDt/G12ImYMknx48qngPjg658tBdbjdhIRPDV130Xl6cHZcbgtnXadI+tr
yvDEipZtRDVWL3n2sJQWaNrYuKiYDsE92DErk5bEu8pFpPVMan5cZ8W8iRselyfj
w0XQah+EpBK9N1S7HDztLF9zPlSaWj7MFN733GWb07+Lm9wAMnAxEYR5tNOhG0vV
TRAfDakvMxBd4w7XXFhX2S9eIZNsJTMr+6z3oP3XAPS24MmQ6TBsANU+HqMxuPLV
vRpCWNG/MpJDB6s26fX4xEbdQ7cU8PFBvvb7yveR2T5gyJz3FsfUBkS3s3Jx+Npe
i5iu3MoRL9M8yD1jHae5VGy4TAgllIH6LH67t6QFHhEpoyOIy9C4QfuwKPIEw5wU
xUbOzC/479Eka/14bWs/BpWWi0iflepSO2NnK9oId2UqDCA/TQS11bAqSxjcVIzE
lyNy6NtPkWGU1wcg8hUTAbXkq57ZXoXm2Gp2cBQnXoKvGuGapD0Z9uVNEI/T5uxx
evYkVdFGj8t48ehjocc8b+39OVhDjSitSAn+ROfbGdkuUEuectC7kx/lpcu43VHh
On7EZ5zoekjWlcy/Zqjx7DiZU+f84HBBAySCKueIIRTkYMxmETHLi06o8n/LxSd0
HYgGYNFQxbcUQzAsx5FWRRLQQlefvDhjI8+t6i0fiERn+QXGNQtVJZd0LOpklx11
/H8Tne0IWraUCJZ9hZtwo82IarDP0NAziL+qhCY4FG7tBOIOeLU9kc9jP85+2oP6
i31VxWc+sR9+XRzfvtP/mlRXOk1n7xYOSkRWl6iUQ1GWiADceEnSyZhCJde0Xzxv
XCEfZKxJr/ijbwA7kpDqsRTUFC1Sp085kbKYUETBtspIq/shDPJMZoo5ILei8Tqv
CXVIkgxdvBbSn4YfHRcDVEi3uJxWPxFQZkbuS9CD6toqI0QO8RqJS9SDuusUtLRm
/O5VNJbciEAi6nG1kDuA9sRYycVyGNnHh5/o0sWYPbb+61RFNly0ZjnvuUacvgWY
OdId7mh5dvw0j/VF555pUljdKQ/qfC/gffhbVQEKsDP3QgAngJ8zzdJqHyFmH2ZC
bC2QVGsuKC7ThI9JfI2r0VoPQItlrshvr8ulxmkzHuM/k7T6LQPbMZYBfmoptxQ6
KUGfYLy6TCcjAorVBx4FT/Y4Bpg1aetQdPuwq8PkpIEit5GU1q423C0fARu9Qmw3
+D3bC2MgebjK7If6plL6XgAKPGna5lXIZ2dv2AXGSrI24ZDW2DGMw3Caqz7wP+kq
9IusV6gaio2UiMoGvyWqa/UEPLZTuuMJD7yFJJ1nKeFjN3A8BZ6/DDihcWW2n3US
+eDGvKkqEBUzPeP3YDqYW7fmTt99ZkNoab+Z9vWhTFyXH2kP1nzbRfQb2w39s0Ln
pGc26DJiFc5QXw7Gl7NfTbscib8yu6OP1P+h/8yaqsQlGhNHGFxkFs9QsSK/U9pQ
T+FzheT5RZ9DSEOmlxRGj0lXM45yiqEr0UN5ttNXAIMCFWONtkYV/yZVS+HpSOkK
w8TIhfZJ7LpNpYelIrA8tk9Ll9LJzGVLZ9QIXoFhvrWT10zj42YZoNCydjJPvLuO
DGQ0+d9yCYtwPSfAD8cTVc41XJVVfNWCI1TSWHjehfyzZxinuOiKTFQsg4h1s2QC
YurxoBn7yL5e0NB8cRVgda6Eef0pI9Fz7W/f/ud2Tl6euEmBHFX/MeboURT/Sfyd
X4eyQi4snrUy7I50L7NhOaDcwsciyYjWBYAVztc6pyak6Qve5uzadITYlFOH7ii1
WL3FTu08IpPFSWh9qN28nXG+Eol2Ez1pHKwZ8i/oNGjYouo3lHwV1VZSq/9KlauD
HWIeI8KFQrSBgDK4l5f1OPt/E0ryq0jm72adG6dUOy1zmogGTgsdC3kZfR+wtO8d
HFinbLbLsdM2U9ZArHHaMHLSH7Y2A94dpcAUdAGtAKluOFmCNv2wTFsvnMiByxDX
TPYqnGP9wHYM8C/MgSJM7rpjhPVTiyjyYpC6+pGRMdp7cfO2hRoFwEtkWnpiJRBR
xCpp7RjHASZm6jQ8ddYmeEOxMaviZdSBhisTN6KPqlJ34PMHBU4ItwBS9oTKuJEh
OLdtZxBbio1Wq3j+lPdVrso+HJUeeLOkARYzvFJDalHmOUxbI2AaADdlw0jB5QQ4
uuAOezA3Jh9Hw2w4+Qm2xeofuum+aS63af7EVNNHLj8zOl3dOZQYZ8Jcl1HHa6FD
ksBD9WCID8+MBDU2svR7bov0cF5FmaU0ubEcz+uCv/VKWqxJhpIzHF8FQKLpPdaT
YEruS0oMil2qKJ70vsoCIW5mRcN8Ayse+GXxgnZI7Oy4kCRY6XY2z+HkiJlhNdAa
CD8+NeozHrgklrM7UTHZnb1RayJn24OAR7hg5tEucCx3j+sHn9BQuWGrhp2+/6x/
vgMBS+6IWCL7vDbs2yjRsMH1ISWnEHB7bj6qs5+kULqbhQC/ZPbUzfwcLEuWF66K
e6XVT/aFTGms9N/by5MzVj62g4HlEmLhglYBVtMn2xh+ZKZMnrvg+u/D9Ri+9PyP
7TTR8+WfGFPg8bBMTnQva9w/4FaVnvuyl/Tt77OP9uWwMlvfq4sy8cKWYsxb1gDK
p9qZRb59xy578Y+7l3dW9cPsjy3dngxR8Lcj7OMUGIdkfzSEfmm5rEq7EEL4J1kz
wmQGjwnAdCMqHPs25R1D0M31CPGHRC2gI4um/fKipZFufFyZwqC9CjuN0I0J7UfQ
3UED1RLZPYTT0/aS+L3Q/B5gfZxBvuzrI9TRqmGbWK1kKQo2Cr2hIX1UwKQjMnVC
2VN657PaJllyOECEP2CQe2g9s9jg/PMggVBu2hy7pdumTJOKcOjNwvpuOfQvf5oe
4CEkkPokS/k8YhLYoodKYApbfrpI3OquKSwqODi/et+X9BVUKavgKuyAhV5yvwke
mcdiarGGJ9a0LjNysidY2rrKhdYotzRDoBhOr3VGG/oZSmwTYer0M5azWQEUgelS
h/brBC+UL/fuYm1yzj8S44gbSMXFlSk52O5O3DGGZkh3EzKEZLw9DRPajoqKRRy1
40x6W8ejvQ6Zziio8WkjjOZ7EDrKQwbBTekACzd26CjMmGt/z5U7v59YdXGq1ptP
1UXNf51WH4dNUXBh8HD9wHHS0hX7TIZWpFqhen/dm8dN2q9VWbV7CBRk87WduMVe
s2hzV7XhonB338E1J3nR+vc37mW+m6L0EGtoN6FggydulZjtahw2uJ+cszo/V6aN
PIEqjTv5Na2s1aw+q3IWXjS+vPICFtjan6Q0omv1gjXEKFhpb406hB4fscKLGq/4
tvEavUcB76guBryoesYODikTwUTyxynLf5m5/xszJDINh2ftUWDjw9XPrStuwOwH
IHc6vSROLdtt0hLGnRte1zzI3dMmyUkteZ3azCz+MpBFTt6iFQBMNr7cpkIEmaII
undDaBz8Ua3izoRuLvjAd2Q4PI86z0yDCuPsd4NbdqJy0KKh9tC0EjvdpMD8fNMl
6cNWzcfJ31Ugg1h6BjGYirObI49Sn23JQ9zOME9U+gXIb9ZLI7AFyElHPgqMvstW
CcinHBvuwd6AhOxVITi/ggMrM228yzU3wqTr7+cqkOzeDB5ZbSGApd0DzZw1iMAn
snmlX/21JFr/Bnqfr7zIWWUF5Ohe5DjCfdoqvkOmi8sWuIAxUpvJdkejrnIPHla/
3vASdoak6/iofS4bzrktFgfTiTnVfn1d9flf+fZXYiFssReJKRnALKBI4QuHN8Hy
UlTNgPXDoX5GE8LUOTocjA7Y2eWzspS5wLB9lUUWhxDGHV/Kd8DUjgJORLThymtr
5e/TOl1cR06C3/ROvDNIDNduPiYYXVzUVZWGtek/MhFbik7D0qmzt45gf4pokChm
EQNcy0KdvDLcf1UDPFt4M4GOpNmTwivQSceb0wFrLqrSW16e66azKgPsJpao5WIM
xVywoZCrDTaTlvEvjMJrBvYK798CjA2x0aYeoAhdFccNJoh9O/W7N6puxi30PdD3
i/wFIJGQ2OzLwLMZnk0Ixhes/jy4JiidgAMGxEAt8hWYyIug7y80sOmeKZ2J0D+e
yxo9A2IkaS+pyFC+e917Xz1tPMTzZTPLywPzqawOfVlnrUwejq1XRtc/oT8wuqLZ
KOA47b6jB4p6LcaW1d4ex7oSAUrfDoOAUIEjLlW5KhGlcMU23TWJlVBMJMHjC5lX
xud4JVSxCkls2sBStW2apKSW1FuFz1JhMV/0XEmES03ML6xW6dYSbG20VtomZFEU
GoYjGjiskYXTYxCze9Y56EQufR64i11a8xeSlPoi9sqEIgirbS8r5pR29Qg9kFUM
DaNqJSHTV+iSidT18FOgxhGLONkjZzGwYqdHWWiJu5rCSzSUfa2hwk9p/y4DJM32
WVWXmuFv3Liak8/25L+KEZqxDhPCgmYdbMgK85j9fgOQwxmrxXO5iLpe0lfRIwM5
neeFg5lDHxphEVKC5U7siND7TwT45V6GBg58uA50mdIvOc2V6YAeDGrnbmCk4WTx
Uz6UuRLQmOSjelxs+7XQuYWdNz9hA1bpABoYDxMiojMqHKdUQ0StFujazDuzDnz5
dJYslkhph2cGsudDg3BGS/66P7zpOATzdQeS8UGXWfza25hIfVsY9MYvvKCjFelp
9u6Vn4IYbT3hj0OhE7mOuKqFvvQtznCu5zIJSLGAOShOkOxWJhLx4gMCSyYh15iB
Zess0qpwO0dmkOB1iw5DRnUdpjoDzgPH9E/vRKd5P889awgUTIg9GWBdOiakZ8we
72uOZ5liupsPz0EQ3uQXBBzhnDLpBG3jJS/4XfIR8nwCr6Glsf1VeeJ+TZBqLPo2
rEIrAWwHk6oTQqs6RYoZXl+JRrmfswxCq/FjNNMjJC1Zn/3csjPQliIqR5vc0bZe
HXg9H+5+Dv0G/+QCTtPfan0Q3p44dkwTXQxg1VxLmKoRmnhra03Uc/zQvrTY4xiG
l3/x+Q70sFGVNDP1OfhWzDwHBpIpKc7ibYnII2hDgBj+DHVWXVU60FCqm8MReS5q
roM2HCKKf3cDXvMUowFAIXiUbXi/keLGS+3HzWsP7ReUn9zc2H2Zh+x3a0p1MACi
CCdFSCC096+6HppbEuZ2h1ujYt7wd05A6/55OGR01v4BuR8lT4+8I8DSK4N+ufY6
W+S4SkxZSp71IzCg0E0IT12lWVoj/rKkOkyGejrFfmiOar8hSZj3VReoAinxv5rY
9lYHLKRU1GZTu+BFrISjJlfwsJbILEekAKoQbPEG3rOyPqbrWtzpinwOC1VRuemb
JcEqHZKCPt90VjNcJPc0xExuDm8lIAudVTcorCQLdhTmQHkK/sqz/PACqhVyr4ah
FiEgneowpXyUupVKOHxAUsmDD+96qU5qOfxEPFngYAqr7HbPRj84TEziwaMFr8rY
yrQuLFscvbdwWawh/kUyaBCCyFIFnyGnBRBkD11n3PzEKE7oCYPxf6GVzj07JkO5
tugxvTnXY61BYzKJ/cYWM2UCnJ0hzjyb+dRu3fZ7RIEqBCiTdUKEhTvI53tN7TpL
pAojtktaxXtR0wtyABwx1aOH9yXFhYpjDUqWlYbuhC5H8jHkjUxtBZ4neyqdNEjp
vOjRi5USwxB6UKbYe57g5/5i4+O/zkJ+S7Gz+rir8MuYjZcwGwy+SRWV1WXgdfeh
TbxkORcNw/TTE8dkT0rHLaDvcjxC56mFWjckI3x0kln3v4XRgOe1ZCnPj8tPrSDq
e9wRlnd6Q2QUkP841Dcm8aINoOGcofqzfaWZlGaqhT1cPPD4UF4xs/NuA+NWniQL
iK1AtWeNVR6za8i+OCQ1kBKFV5rApdHMTkZ69O1kM95RWF0miwz49KSVmbej2duq
Y+sUPfJzvLQGNDgSRjnjGwQp8YQo5Gnw6V2RNv8u7nKpOu8MPdchueliAPlsGmFu
qBGKl3S39KsilCRT4r2j1YA1TOShduTkZK7Cw+g7yTM42ELQmpAMz6by2XyCPAL9
Ma5Bc3FnMi25cIvMQv0hluSqbi4mxqpE9uHvliJGRugysRIvTwekBlm+S0/g0ETr
cBu+VqJ0Ug2CH3Mu9JHsNyDIAGZ70Q6kI6SfXWVDv/sMIbfRylvVQJJnNCIQqIE5
v+NBYTVDHDJFe0pycePs6dtcth6V5RL/bSVhIPj5jHWYvboU1xIJyv367QpahSpI
LVZpqDGrYefCrlt5oMR594LoXYb5Ko4kYLOJLMwuFJ+u1g4tt5RMhBXX0ECJmfeU
TSI5brJS8AXLQj+ln35ey5dNcOOiaxLJTfRiQIfWbPUwnOU+XLJk+rxm0EeaQC45
F4/WxIueas9By5DhZ3xfZNylcDalT8tqdK+5C7RBrbnt6HLegWwY4fRM8q9PcViU
yUO8u/MFV5q3Mhh5KqOKa9dqIXEHjBf1/btofVPep8lJPCyJZ+cqUWu3saIZIRhE
I7InRGrvHdrtdbhzZm+wvLLV1VFDEHmcgltevD1wePrCKW2YmI6xE0aXS6xmNm1M
K0Vu8h6DuJIZU4L4C2fJQ/rRGoYx2jt/ljL6z60Uqw6Bg2myKwBxJ1fW0OdJ3sQT
f328qALV7GJFtioa6l+xi16QoeH+cM8KzDS97V6hJYhkNL1RaNTzhjz7b7ltb86M
BDfETq+53PJdLBoVRzt7sP2GosdGsAYmdcuKsumWsJmgu6+Y9buGwElAmYF9lWp8
MsPOtUiIN1Is6JdgfZxdl8dDxA9OvujBV4DBc0PkRjMq+mzngAACvbmOcbLF7s/i
jXxkMKtYrll+2wowIDiArFfEc5NhVx1y1a7/n6/EN95VfEPql26qRLv2QRSc0ffd
9EZRsaXcFCDWa82z0UrxBk/u1tLf7Lqs5BbnYI/xORIiz6Lsbz0zZL4J+TeKtGLP
rMs01OC8Gm5CFS1S7z+C9FDzLckmT5nZbsFgV56LbzS0hvtK5qctZEa+bo4hwoIQ
LvRMwehMbop0DxXucqPs+sXnLxI88R1vdbkhC47eYfoC+YgnxPc4+3jZmWOz6Ki2
IWYFna1o5+QnfCAHYNo9tqs6va+zQQa6TCH8Em/J2/1p/BUrDINorHoWxGK1FBHP
arSr6y3YGI4IanNhkNo3vAXGmDr3xsc1xjm42LpvAv9AG9gr1ak/lM3HFeQOfxd0
9fZKSbplkKqROJsIn0dYsavWs087eWOER36tg78yrBSvx6xkvSPuJhkUaMKS9h0i
A6w5vs5QcGjKgVRFY7somdDz4XNPGCWWMRphZPwGZyBS5wj8OpBYzft1jIhea38Z
TEvMseNa8u/WEGeHBC70z5sFmQoA2HX5vaJE/1bu1RdBo6TqPohDhwxtPt2ECVqJ
QRKYY1R8egUzHW4E2Wuyzk+WEBCDB1aejlCDYoWYO2J7MVdM5qMYKA+bPBAk59VR
mor66Cm4Ujk2lewoii89Mv1HFrxuxkjhHc4MMMKAhDFOeFKJY9qgoVdklt/EmUcl
KhKmDhMb95uTKXpWr7aTPe7gdK7YiOQPvC7ac39dGxUtl7RvF6F+jy+d6hRX0znB
FHmzFfi5TuVxlsaFqBCyREi5SaZZMcAFvFqvHyX2r+tOHQ3Lw+Vj/rpwMdhHFTrb
q48327OiAmNBBf/eWXVvrBhnatNOTLvKi713g4kd1WJO3xt+7cX/EM2rcFsiKhgY
WpzdgT4yg6jiRdZwEUS00LN0L46rW88QtEkqIXYQFKD8Siopnoir46Ioo/FwpfpY
78IdntpPzXgkHX2zxFjwggnU5sSEowSrIYGcelspfey8TlEeEVYK1B0TP2mWCk6P
40X0ui4km8XyGP+kQvLNVgpjXfeoGt1tVrmLcoU2XcSm5Aj9o69o/dGSIb+9ZTBf
Z7Tc/zMuxc8U7mJ6zD3wgE3G5gyQw8yzFoL+CT2Wk9dPWhFF8g5xgqop4ZMOWZqN
n3dsDUBGvGJZzNx6gKuO+sprLK7uyxX66rZAxQEURtnlvG8ufoP3Ly73j1ZlzfRT
sWjcJjHxmSpw2OGsO2x/LCQegwEKxewr1VB9NAgmJcvI94vV+SkzbnIVWQPpDXgA
Urty+AXshbw6lKImsZlzhcyThDg6vUPV6FqmCjO3xYE+4Bu80TAc9R5cfZXRZ5cU
uGVXcsv3DL6McG0U65CKB/D/IQbnoRR/gvLS3xS9tHJUbMnAHhTHKayhx3ZPnZJW
leorR5hLFmEb1EvuBj/LX8zKVT9x1XmlzG5t/7RCrfcbjXGIbuEEjerIWhbTFSxW
o5I7tEObRzmZgOSX+axaQK7oGH1qkvIcvz9mmIMOWe1LlQ5C5hlTcMgOsoxtGzzg
Tx2nr8ABQPPRxMnerus2NWjc4gJ5EH9ORsdLEdnvlzVOvr7xaGhkrf6GqDzhIh0k
kSHHP+OOBw96QY72nQPQCWOwGO35VYL30P6irVQ2+rZNQXk/TZrXH2G5JLuRaVVb
08W2s8sfK37RNodyRHD+xxq4yCqCKuAAUHJl/ve1SBkR6rRYZo7nt9Czg5uBS1gM
fKCsoC64sW25L0XsFYWLQRcv6LkjkwIBeY0V/AdhTTwxq9pt9mFFkgicIbuIhE1K
uPuR0loUH2OwcNJsggAqkEztr2YcSzYJVU1D7YH3tzYU/5GW/i4NAuI8FXd8YT/d
nRuSk4RZOnSeYQyxfY1sZIzM1hHyYrBQ/HMzSrzW9d+4TMpGbr1Cq3ppdsKvpd2T
PF/l4Lsi2Wnm6yDaxB/b9mUmAkGgXPuQv0LmP9MUSd4N59hG2XMK4NlYpa5ywQw2
sHRN8dS9iPqxpU0KYliRHATmEIapJRi3GISflD4XrFVl5UePE8WBoJtA83KNY0Yb
PK6ryDMSsm3cFf5VY0mbq9ATXgjc2W9ZDDFCrDc5f1wTTp1IzYr8y0S5ixalpZaq
dsf9v1DaRFnOtosURS9UwdxKgZCR37UMlBlXc/9IY4ft901k7PulS1qfSnj04jF9
EPZeoDYcu3TDPRNAtNPU7IH3yYoVC30ENNoKxxa/3pWrVmW9IK6uGbGDQpRNJFmb
U9mK6AVjevdWOARk0F4zXhtFHGlI2wP2HxzFAvWuOUv9Q4a9CT3Vi4txT8KeXCX8
vP0N/d0ncD+BySLQqWY3BVKsXEDh/j8W1OUMvSO4WoMBjetlxca2Z//Jb2aUypcw
fiArH4aNskCsLai9sovM0+mva479DnN7aKHyTPIhTmEr/DsTCvtAWN8mC0AG5QXI
FfFVthaeGRnYAR/JZHOFqS4RffQdJIEOyxJltRjsDMy7cNUpCvIzOjthyFpqJhqZ
lE+pyRAxtY40gSxJRJuMfykbMLj3M3wGNfMCzvkeNcpqp1aw1ByO2EAwkDNjScJa
U++/DfGa6Evaimw5tLvgYtrIRqkOpFZaEG6eOS2YkpBVxtXRFf/iHBq7H555lxH3
1OIR2G7v2z5PE+KDgJxTeNr2yXCP8oG74vHqpkxXlC7MmxpFxjQ2Uom+j8VRyNg4
Zc0chB0EsQ0yrb8v9gR9k04Ck9zvo17vLKiFgSOaLFdJ9cmYNRXi5F/Hqfg+SLIi
EyHM/Gxw6sNAhleGHP8Bq4/6xTdSg4tgczhXYbjrMVs+tU1pq2ZwSOViP2fVuUYc
awGlKH8JDuItk7Zwm4QuJUitTXqwEkKyPClxLm5/CcLbrwhlihny11X7w4dU/CPm
1jbEbTa2ClmCTxrOxdrJHaHgLVQQ/eULsuvBSaaE3vNZVrU3K1yL8ltBiHwpQ0WW
ShrUfeyPguWWmESFkHijgB6+Q7NX2Izm043+LvBvt0rCYdEAicHq1tXcBP+8hS5t
5fyItom+SWikw4sCVPwF9HYIhO4arD4NHjbJaHS6mKI/2KlrSTcGvGLIAzqhrL6F
Gxn/kxtj96DBOrHRiKmsOBCx8xOZ8MOeqZQZeDQnOEr7qPggGjn5C6Vm5/THkAa1
qVd4eI/3MpFeaxDv1oMRcbWay5ti642FfR6ecjW9iO8W4mwZYnHBPqhahAFmtOjq
4bHJL/yOZJq0mZKPJRz56ELY6NOb9spD5Pafhog9fJKo1vnCGaBz7x1ivHcN3wHt
A2fMfs2Txt5O32zzSjmMNnhD7gLrMGKwkzcVy68TJ7M0MW7LBbEcPy7vuLVkYxT2
OUHURvSyrDfK08KVevQJbfEe1e9qLVxyGBgxbRYvlKYWunMRD18mhdT9mvUD3QVl
wu59fK/OrircZgL8eKscpJzLNE5RCqJVfOjvUD1FXCw5PQgPMww78IW+n2KccUM5
+/22cc5Dp6yRMqptcRi9PJznQcEnqK9AW6kaI0LLE/7Py6DHP4stud/iQgGvv3Ii
xg015GQUJFndW/grVHaFFY9+P/ZiluLlH7z50WdLuFv/46qhtzmFzq+GAIxtA/cN
tp2IEJ7MyMp/8lExGmackAAQW1cdRTizCA8j7YRJB8BZTiZiUQ+yRuzNYokX9YWz
q8gyKWSPXsD8JWcdwVJBkfNTgjr6ZIP6xAgoyqYSkkQ2YypbKGrdeuKwNALVs+9I
hcGnCUqCcOD4tt0syTaLlqeiy285mKBQQLPpBY9k6EcfOynWPtxf8pxEqdmzsbbn
0gr15sbtFYNWSPhhDk1F6Ha8/Y8bDFG7vVnO7JmUb6QH3rQxju6fBp2S2cHWv0K7
HYcN8NHmSvlA9hqJjvR39qresejU7rVN3S2+y76MXGaQaGwb1GSfm5xOe6AHwKjP
zvjcsnjhPhb1hubc4LQIuTopxotrpvIE7NkcSUaJvBmx5nIyCobfvhJ+quT9AE/i
Sg0Tx0tgekRAwQhnmCMNNhxtWiIp5DwGoRaPYf4YFmSxs552jH/w9g/Ps40KaJJT
AA+MMcwymrVOXDLaFJM0pgpis+fAwU2ZUtrmgZK2Uxykqw0uHwK8DtnpAXbW1gdn
M2Wa1cdgblbJdixHwLQpodte2P84P0IEIGIfmMN8TYIocAQH0YjKObPUbmIIa2Fp
fToFG+yCcb3QjRKID0m+elvc4uLT9mtV5tToqdsxX7+b+ISZn7Ht/wHyq90qe7i/
D85Y4v/8heM/0Cc16HjaNUkwQVLBe/bI/ABlFxqCjTkFpTzvc7KWhXBiB1LsjLKO
wIGGlzP5crJv8LZ1jQFYiuyaqukW0Il7bmFUNONqCLYE+tHX6w6NPzDs1HbhiK3p
fgCUL8tvbLRNcqluzMIpoK2lLgA+v/yIBD1wHnJcocSDzLC1CXfaKocEgENRKW6e
MwoRU0vBSBRbsmfZURUbNmNX4fP/2pYog+T4KEUPWUzYEwXzPZoe9uBE6p1rtt6B
xBODsUi6uT/RB4ncYg+N0Tgx6rshpy1fPPdAzddPhfdxpnTvUoT1JbLEidoWLTji
EHt3t21EfaOvLgnLi391O0SYXd1SQfdOy0oa6CHD2K6GlU4KyUcJpr6YHw+8XccF
LpvJwfqQ2XekpVniEqcmgHuymheeZ+zwOomSTuveGM9f40MPWxgf17XSkfrKkjG1
JyjEtykkIsUN6y177oCPxqYrH1J+9/F2cgY7sEsl4uJJnlZD9r8LgXwYH38jnVmN
x7z59xhHEnFeAKkszlozVCAUv43xjS6RpVsmifV5PRM8fooXBXNI78n9oW1kF/t5
jp0f0QV9NeVlVC2TsAwhsgnZ7zNEgUmzBt5EN3CBXJpbLr6Pn9MliCANWGxa+eoK
h08nh+0vLzNqx/ObY4v3699oF1eHnax9SSr79I/lYzOxCQOkS1HOUuNwnymjLsjc
KFMm3hOJ/n6Yek2zb6Se5OrbYktouAwp2pujjI/UFqF3fxlLem5sm2Fdvt+VVrzg
Gr/wf8yIwgJ0zWk+8qCrdUlMM3HUhxX3cNrz+eni3b4dT27tpkzeOXO+9Yi4wkoT
gpRhkoQyvyGQ1Db1UhlYBRvnO2vAOyBNkF86LQKsqgRLKMvB1SkZ2HlCDctEKhmn
k/RPww4ABvN99/lMEvPiheAaHiRLkJEzAdLJGecfr3RgTrg5xEoH9/fq/LTseTEh
S1M/aLUicQnpse6mjn/tVZev+iv2vrKViaN4gp/OpijSdOFvRFwHZwPFu1Ey8Vog
T6loaOPvf7OmmlQPOAKYz/R5z4kvBugFrpcpj3m9drvUC+ADSrPJP6Ad6CEgVrF/
DtOIqDY+qJ4tENC223l9Kj7uvzC2/6OiBytkF8/go8lnq8/SNeDAD6ePz1tiuX7/
XRF9Ta7jIeLqlP+miuvMkXSxT8cNepZy4W/OnueJh9Gy36FWFIvxyfUQc4hMdjbZ
ndyZUHWFtzctUT36t4dQliNQJgwwmplDtwyV0IBMrZYzuW8P6AKY4XbT4OSAjla3
u8hhQCsdUegqZOQ6TTNoQ/urE8eHiXVJOxPYy5FI/afowJaI5C5Q+e/FS363OMFE
SOlaJeeo1nGIsYE2npDdxpTcIIWZ0c1tKFdEGnIBK/YzQTwIVhFtqf51TvNUuPdn
iV0SMoTBGSTGkdQICXBOuwDGTuoE9IHKxKjDYUlGzPjzRRDzV94YyVJHlLzdha+s
gDK5SPUfMO1vVLS1S/+2QaWuFJSzySNwypu0xJfR7JpZn2twxIOD6mKkiLACaQUV
iANxqpOzjl9DfOyTRN09QQy9Ex3xG50VfRlBlCKMWG/RmJXY/CnzqxDV8cZnHmWU
17UGgnXFiJtnqeNLUTGb/aajVqAVWgZUT9mWrXDS8EWzxBg+bAyEwy1xgnTSkwJD
+Vc8cr3LaV86BjPYQD5EZ+qdlSMLYJDr0pFrH+HgqqEeHIZUhcjM6UB7tajMvO2P
3uHBQ2X//lqKR2YrkdzAg86WiqazGHwdTY94qAg1NttjDgTKUGT1Cy0cnIX9JXfJ
fBFx/Fx/NslTu+YFsUocvmKcBd9FXRHI+eP906hlSmJWzRoxKja9Gxa61/AlyM8U
VjoQ1jYVkwrQVibdVfgtuaXVqP2ChA9Qq2ZK4hr+Q0F8gCXWZNUKBQtGlSV4yrNq
QeAzTLGj0ys90TTHh3lHzyWLzBzVnqS9FFcTKilVghTQbWQ7y5YLLn+g/EImWfZ3
hr9x5LZMcNeZjuWIR/4Zq5J2yK6XCpW+wYB0/jiQcb6t1W5o9SbN9yzBOFArsLRM
c7LCa79sNmwf1/JC0qXjOKB7nRTkZQE+6J2adU1LEbB/3xalAo3vNuYFwyXnWrbQ
FeoNUh+dHQQA+RmMNtSdpsjqw4V3yJQYU54wnuUxHOvI/0wZXwpGvIjCnx44rmHI
MOD/vaJDgthUYUNwuOb5eZJ375rCPaQI/K9HQPz7UhkaVqYMauA9446S+njHNOdo
VxlzWGocME8RDQtUhDnGRuw7/fuGSMdJ2lUasJeSYbDENxc5ihbOWb9ugmm/MkUd
Mjm67bnHYFPqlC2JjUw1zEc+huInZ1Mh491h7DG9OI1y341Zgy+gkjpUGAlsvHjU
jQOVHHc/Jg2RjFa828oYgvJ7KzbRHlGR+guB5U9UzlKRfG6TsN7Hns88sii4pWXe
8NSs67ltsIyQbAKsLj8lN5ZU2oXtCcxvbnIqeAjuu9ix+OxTbgsyOqf4e23rwRNg
f0B+R6XSdr53S+m8h+N/HpsSjk90n27HnHE+qf9wIoPfNzPyruvED70zUd9NPXv4
P6WBDCIFTtqksiBEsHHUWIsXfEM4VBPbNcUunhqq4Hr9yzfTEQILrXsrW/bHI/QO
XM7n6M3NMnAuWmV+XRnEUTMx0RB7VrtmYD0x7RDfivoDAi9aPUwYF5f0rokaBPWT
N21ZPEvHDY5XDd0VWKfeV+NiQjSw9I+ik9a65rmK5Xd7/oY/eNwKntUVuGfOuwMY
Y30txlTt6vHuxQUKD2e2nXGYXO9sHjzTX5HlFeTA11OeLq/NMtjYDd5WkngqNuL0
nPoeZAZUbWUkHCFwx7mdWYI3qK8PlRE/xJwIFGYqs8SpgsxB3wc5glDqwljfPxX8
gQG94xeVnyo0TPyrPdnQMFAWti/a2nUNLYAL9IOv6v3MZ2UKAmXJPt1ZCv/X+M18
ooKHIHNC9P+ZIPC25yfaHb3HxUZQX+1pPdE/aLY/Iw9JM6ZLHzTbN1L3nxdB+/xj
htVSU5wXc1wfZVacb5998zwQrr5BQYj8SpUJceDRCRTZqwFAV/JVFJPxT3nD+g6w
ZPAbhko78Op4bYTSpawOF4H57vznBH/9V0GaFgt5rSAnC5mjMzLTBEBW2SztsZzU
7LBV0cb8eJsi4JYsD6A/cVa1KBFWxsnaNsG0GqkBKuda1QX0PquBGa00ePBc3WxB
UIRT+zCWmxj9h9RngzuBPc3s6xdTeMvGmki4jK+R3WwsU3e5S6ogN7BK8QWcGee5
M+itpzqkKxMLKRvdStlKia7qKwM1PE8+8ZkvdN9iblG6xr7V6c/EuQF3CkE4PoDt
sglntuByqOIafkC6XHlpgBkalpl/in2pPv2M2cA70jzs0s3YM9yoTyxlbkl8qrXm
XyjLmNDL6ZEn6M5ukmpPHkLlL/qIQLuAhsjPwlVKx8sHZyQJ8hzXFAJ8Tn4+RFys
muKfegrua3Uwp9OqXlfhUZ//N8txsAMqtncXMMBttygWM8gbcuu7tDfc25LTTRng
JY0CSpGikjeITlXWdsZIoVi+vRKKbxpEAW6R3xgq8ypzs5QeFiLaXW63pebuOIhO
E0EesdrVjXBH1FyLnPe/dOYi0EbGXawhrIQYASWGKMvzf1K6n0tXk4vbMJTNi9Jv
/fhiPcQcACiSmieXzj/akNxb1dDkVMzr8GnGID7feiPxW0SWREXlepBhnSZF7/Ks
aFtGEgrMXabr2GQwEShFczVid1lAVA5Q5Dde7pWQWao0pc+xku0c4VB83mWkCEgF
lgaTaCOQNktoK6l7FOL8hUVm4C5UmGQFkcoZWB9RZFA5kPGNUIOi4a55R+Hwhe6w
Z3z+Zkp7PFJtu6re01J+JB9eeRuppiB8TXcsBwtX63JCLCvxe+tI2TxoK5sgkuJb
8DIkfPBu4sbyg5Z/K6A64Qbmejq87gscunGi3m/MJ4zfrG7vNRPNqIzZfUWxZECH
Fjlx7axpM6PG/xMLk6gOd2VCCPMWSDKipcbO+dnGLs0FWEMwSqjYGw+TePhxA08k
ImrMfh3cVy/rY5CJ2ECLUiEntCoxGbFxTRZknwNnqrkG4KRYLPxJFRB1qf0gz/11
Fil0sRnqhuRNlwwiPwxthTFr/vs+UzqpLb4O79IPhWArEDwK3oE17cpGU7qknUl9
yxeb4i2qCTEZ7kctfL40d5JFNcDC2ECSCHr+tCukyE5p08r7ylNV44Ra4PxD+dyq
vwFC7hV1ZzwxOouWVIQFoEXUwPxuytYAeXEWV8byrahIS/5jDuGBmBDJlPNtimLU
RbEA+LDQJynH4OSgtN/sdFFU2D+RWIAKIGYZWluT2DJqM+fsmsFTFXo0LXILgQwz
zQZ08i3z1GT+CPtVhwEM1NZOEvbRquW6ll4J6Vp8LnhbX1/+OmLnMbnngdoxgYci
FBiHyHLFT/65TEhqqiEKf+FJl7o/SYbLx1fwhJBbdVctJ2w2emUECzk6J4Fv2ppH
lbXY9T4ptWJTsPHiB5Z4nkP5gE1qYbGqfAYEC4+F9T0YwYCvymZIWD87K0SqgMvj
ov8qe/b8TpC6YykRwzAa95PH3DIUf7KBKeQkMF3H0NRTkRYWLeI4SGSxR27IFgFN
Bj89QdJLspgOsqW3orb9K5AFP68UM02kidy6MkCp47WgWDL1XDlO2+PNOHoFTnxX
tWmMFr3ERrmtx7WWLq6WUTjIziye7GlEAw2GNNI3GPY3w93hF7e4crVuPk3RAxvM
U8NMP+NfkKrFpK2a54ArueQRnbaaMZpT7T1ddGZWvHWeN2rjtr0252ve3sbtJqo/
wk9vK5urlqSpD9OLqlFbqG+b9uy8oXPDesS1LFIrjOKLJi8uDIKhigd5BC5EBGEE
ZJtjOJ9oDnoDLohu2TSRH+8kPoW6ojWX9ljqxwbld2hjP6ofChl++1zfdWOyBNfI
4k3DFnM9KrAE5djQjkUeHc98SUd+TSO9Hof/PFUFHxELIC4gK0Nz6+PHsoTKgP5L
vcBWWvltkujFaJkxtrVGHD2gGHdBYzAYzFUU80NL84wngajXnTYL9sgAizvRKkCM
bc1RcX2NqfX051X56R+47f8NT5Kc1MulDIPawh3zuwQ+l6JPJxyoJiSGTwdWnomq
nwUyjjSriZTGavu0HjvH7b95Zx+92FHKsqBApByKZMPXyWDUa4Q14LkEBew9lZ60
hy+hrimJOAKEmLDzudmn2iT4NMIyz1SGDPn+XPTpId5ruh6a8aXLgKHjsNbM6L9j
dUbYW6omQjMbImQl9vRZE11S487/zTWQUl2QFyIIO7yS/iJSKlpRfF6iuxxPXezo
z/H6ZAIM+nKbvBZhmyEdODAHXpWKJ8obarHln/aAU0aqSwvM6lKYDTB8HcIg3uXV
0nl5Hb0CjnqWjFuRME0LKolCpsaOlkPC+E8NH5NAPb+Mm4zFfnPa1e0gCwnDQjTF
ZHij7B9q7ziKceJRsu/N9dqM3XDLXy+wPCX9zxhcBrG2MJhoJrD8KP43a/WM0o1F
Lio66w94hC1wva07HopTbPQNGm9phsodxG1gPDcPM790JmyOp48A3OjpP2LTvRup
mZAzxnBL+JlOTkmk8l57/N41e67jMIzih7D28I2nlll9DFST6ktWt9r4PrR7sWPq
OSE3KI63D/XMx3zMcZAofYp3VeTczEHS6gSNfDS3bHmT4fZ3dGiEQjSISbWQTree
ixtb8889KGWC/B38E/KZEXAKTyo7yxtXJ2Hc6m1Mr+NWGfpiWcOgoeKWUk1mm84u
JqvLfkyAewwGdr2cwi6VuQSnfdSgdxd9LR73X4AF5fDUjpVc3aoFrQLdAhSiDqSO
rBrcCQIt8AtU60xsS7taW2UTHC9fKTGJ2TvzrWImcbk2yJiRZOA/RNLZR4trQdUG
4uPn6Y0w+13FnB95hE2/DnmvyOX3KE2W3swItJPZvCsJosmElyarWZCnbKjPPgkd
+4moPxn3mZYsM6HJAOkBQsMcB2iGEFBV/EAlQBvxKZnmIXpCICq+nwOynp/k8PLT
831IBFABn3Kd50EdG6bLu4HkgxnOD66asLTK0ySGbV99fZmQp8yBCaumots1WfZr
3nm8FaIbiGOnNBwl/bLQFOhGI2DOdFBUE9/1+Kw5kvFxajDW/aj2hYnosgJssFBX
0McR6fn3u8uk8CaOdjCdOzGTN+ZYRWyVpTN1DbVdMT3lD0i01UT9j9lCPvD6NFte
mF8t9AnLmEU2oMrUveAuhhRwZT/gE9cmVvX+Vdp34TRmzEU1nht9TAfi3lnjYHnD
quvu4hgKQmAlgpnHOx0J9XE3NBj2zM180+pWNLtJ8AdTT8FwDLcweSG6bbqD6H4n
D7xCcxUgaC5vKBbFt9ykLiIlXaST2xjgvh70+72Psp/h+3xALUul/Y/6zO20ICWI
nZOtSXW4me76qKrO30KCLbRv/NgkrJp5C37+FWQ8ddW63UypdNvTcIIxfcXremlc
km5csJUquC7IM6uORon6EtAK+lxw+kPKPFZYs0YCXmYXYbzmT4wBr6zjWxqVaY4t
H5b+sjOCHrB+NqH9LG5nha587Y/Dai5jvPjwvlqkiJyvdB0tfsQQygUDOdxfjgqf
ocVbQI858n6QB93lMtQuBMA9XRctE8MXa9izjaNZhtseA8CULfvYVRZnSYlgm+U2
vQ6R+b3/gOdcbmzd9rxRj2zroiCuwVPQFj1y9y71I7fJ+PUX1MWCU0NU1QkpcBsg
g4HOScfDm8aCG0BvB85RLSVcm/XCN/PSB86yWfKFOhfVK6UTsKwC7jOxt+cMbrmV
AOkbLRKOOhv3+KpZZC927qiWW8SiD+BTPAsmDNaAanKPcxRi/b5KqJCW8KO5p8w3
y6a426mTs8++M6rDiOt/UHf6Wkr5bVwO5xiP0QysaCmWiS5UHB2XlDEKUkDK5tUF
ENa+1OeHY7pXKFV//cmPlr9c4JyjbJVrDulKCi9AfhyVTCn0sv2QmIZI1GdNG8tR
hFpofXlRMBKXdEtdmdl1zriP3UWl+pacGyEEwC2GnYisY2xuU62kyoXbsDnZJXQ/
LqLExOYJeXO3K1yRiV113GFjbzOSisxVF2OGBZrr6mD5pX+42pxmKOkQYLKOSVus
2qpzTdN7HpfUTm3jG+vSVT8P2iBPS53Yl7uyWkttUl9g3ElAeE/i8GZNRh4eA9PO
ADFIO+2qhENnSaUCh/rsXKMIjsfg9GJu+m5jkLg2MndhAb32NEeKnJp5ESLJVnF5
76s20G5lcHl2xfwas35Bj4VBpe+Egp3Na7VB4tPS16tCWk443kYvn1vUfwY3E2zw
oxOy344reE8GURO4NrJqduW0V7UH1SrNvEEKugBbdW5gywSNnSFDV9uI/6pnfU+d
oBoMmq/FIwWBHFbmQBxoFr5GnEeeQI22IqSBI7eUkfn7R/cBPpqrO4yRyHbwZ88T
54sHDA1yu2PqPS9+snZ6XCXoIU4WpQm2TBR7OMurTnL9xmYaSw7lUZkIaVg/be3U
B5PjdU7Fv9pvWb9WMl3UDd0ITBxCvvc7IuUsHP3ZY5uf51TSH6r81X+X/ZOo0Ahc
JA5HNqHmTK+kGd9d+e6oFfHD5pH1NCY4zKrcNOeCH7Iorybj+5rGJgN+YfMnZlGM
2v1mJvTB0sE/u552dYPxxMxLLqySf9HXWXTa4E0b1SfewLBwf0N/X3JKAfMLznUE
aa1w5LNoSqyUK5Yu6CZCKUuiDHmA7FnZjLluUfBFxRSxCVlhogxnR5Ja4uxSTlRo
3v9d48Qid+Z3dFN45zsnrSFfPElUq1LvKJm1GzE2j8Ze1mxU0AjYx9/q/0oXmQRw
GbnlCE5ZboH7ZyUzO6EkjyOJ8QJ5kwh6o8UQEdmm+IPX/QVt3HTGjv0TPzDVeKmT
zFTdoH+2Ed+sbqVfBaG74I59ssShCK5hsOJ3D9hEcyPZi0zGFn/eu0ExPLuMd5Yf
U4BJzzR4TfsDS8JJ51cP6oQ1ev2kfQ3rWwXzNYIL/NHrVMCa0yNmMXAJnSiGEo2m
94dtoImgKqhEPTKuu/3/FXYE6C6mLD5/T5JUMqhH53xhIC2lQEnwIe8W7/Le8m/7
Fesg15gh9ez/JDGeSMq4daeI7EFnOpiprIKKiQ8xoGksOxSbwVxlyEiX6pwLU52a
9Gg5P3xIVDFH9JgxpB1vFerp6RM4/PB8ZbMknc62pJ/2I4+06m+7f0JQxwH2WNQi
NHVKd7bHmD6O4UfvRKoMZmzrW3FxpwlLKi6KdZv+B9Kb/T8YfwvegFOAgXBOm6Zd
0vl30IeKOFmb+1fCkFqM9GOZB7ntUG2BaxgDbbv83ZFjYs1RLmlaAin/Mr6lnkhg
hnJI2vN5MtP6qcUH+qk3g+EgCEXd8DrP/6fddhBAkw9Mj2+5L2EH93/aS81Pk1n8
uLyIRdlpu1HwoQrNErED/g80kJEaMZL4Klkw/aRjODHNixpFVSN41AokpTwCQYf8
2BN02N0WCV2obU48nwb6kY4c/dxFWHooe3p/ep+1A2GMYtV/EGzEPy/hgDOGt4G9
m/DjY/PHwlS+g72+80+P4Fka873amGwnoDjgdsdS9lsxnDwaTwDxGGbHRxn3W5bO
KVN1OwqRMbYoshZzUmWZSNsZWt+b8BG3wC5oKvkb2lT4YmOqc6NHtR6d6dwDPekQ
xjE8WpyAdknfUZGh58Q8PS84dcsaGnoxUustOBUY8A6qcaoHD+eSAjuLMKwbuJLV
9nDuPHHZV7ZSwz6zrPOYcoSv5mubayDmJEsdt9vzUfzJl8yCZdREmaV272neAZEq
Mge1q2GECeLt4SCcduEl61OdNY9DAfklAIjFIZR5QOfilSkFOH3bWBtv6SxM0KxU
vvUPMyHd4fL/JhNnmvSuBG8lh9V7i00r722S3ev9g2mgXgJzaGA3BZd44FgZm70X
J60JKtRvRtfXHBjz6BZmRfyGXTJU8QURajC0eZwu/qOBWxIzwTJyk8q9Q7VVJMWk
Hy/G142hRjLPzxPUFmIDNNyRBUQLBwRibjX3m9MrukFg8dS9WcNY0gQvZpb/Q2vj
kIAxzv5c0qeq93BX/9S7aP8IpMW/Ya/YCy5+zQ9uORcTmuuSxcdW5UEN91BOyO49
WFfhZXWJvmWPnX18RN4urdccG712GVvQbfkcijLXEP/CMwHFeDvfbFwsSDVEOvSc
K7l5jHXNnjJq7p2hnwF9rYog++DZGlUQHb9KaTnj0jif3ZXtm2CgnIO8osHXmwOx
Dv6oafZotJRD9W9oJvFU8M9hsIeKHMwJvO0ZHbXt4napXfa8x2OdHhAkGzojywce
L4dJZ72CMVsWX8t2VKLxDdc2tImUB6cIBEOBfCCkq9ks+F19cg478ZsQSPzQuG5c
8z/Y779sJ3CPESktLjN3dIkoNkKGnguHZL1J3YABxiJG6TM6xwS/h1lbNiih2LJH
Y67cbAgC7zWfppwpgecpytHQQIXe1OMGQgRjGp23dS2Aud4eVnpz3WxHUTwe+x+4
SoH3tBFeZDfeDUY0Ap6MY0tojN9Qm4gn9vKnFJ8Giad2JDSaoDYWRmUOsiLRJHk9
RaoAG4At2RtV7lzuZGzPn18m+4rC3ivEOc3pnY16cwom18ZRhpfcFPAFctjdW7s7
yJwLtePxIFQwWxAGT6O/xbj08j5kOnTbidq8sKgTojYKhLPsW5M7K5jK8uNUqPmf
u3OHzmgjZroQQsGdF8fTrVbgXbNipFD+T1NcbZwFfnt/2dImTJxENa/8YJIQPyTK
QqnsNuSXLpjoyf2ij1CxvuxnaatGsKzPkRFQSnccK6poxMWXDpbnQSOwHKY6GLFl
RbVRT80XaeRn/yEYmOpbecUtYaUqSBiCOLkMivCG6yY1maOroZA/qvGrfahO4asx
3wnAi78kpuWJEGvVpfGHQdmOak87uK/TPFztoIoY/LI1qRhfh7w2UqNgRbIC8JMx
0VgARIeoJdYB2YOKlPP1x62M/yIPRiwyuGV4APq8ThKfYTyXEBySk1zBtURkRFb6
WpU+PtP5BSDPT/zCqQfQbaXnWySeL+D03RvkUROh4pVD9lNBVulNkliM5Zl9ypG1
7Qp5vUbE3jA7u81+sebs5wOKvZ3jdsLTwr8Z4VfF6hSvFZhA9amuTiJgQQsHgErz
Vnk/i083hx+ynaXB8/81IET4Qvf5C47IE/ZCR3RPioUmUJyIjutxwyASw6HELq7a
GTAWp/xQKAtHTqEN8Y/Of9WGlBjCAa9W6splzP/u6pQwpW0i72TH6v+RENyBmqO6
XJcvMylB4w/5iWOuH4oKP1g7ck3dSc0GupAMN+yxc3vEl2gMX8PSK+O6uAJ7SgMA
VI2iaept2CenXqFh50pnI4qID4SLW8WS0s0myXDd2n+0DbJVbKXskkIGbDeQuXQv
fnRc61yvfMme5qxpcUm5KdpTqAhC6FyIhzaz95w3YV5DTfXVLfZNN+7Uv0lECi9M
yDO0a79Gvwsn0aomJmpQf1q7XU5vyEgYOA7MTHfi+Q+k4Z7PD+rzYzRvWZtE1nfP
0mYjjkwtRhUkSiav1e4BijIFBVAgzVhhCHT0C6UDnIPn937MJROAMgp50QV1Lplm
ZnzPLzVV21YzyQ4L8ZBpqF2pN55JcdFnxCWEjmt2ZJuWmQhQZ0d3j8VStGBl70cF
Lof16t4mfujijKn1jihNeefj//L3RueHCE7t+BbkBBKVmKV8X9yiwmLmIqmDvumY
0kzaArrIyJRG9AbjeWdw7kPtsCzAQXasXzELQ95w+1/XW1Wsji9jaFMIwuZo8Z5L
euv1uLHJgGh7mpRZ9EfQTRi4DcevCNSfoojYkQiItfdfPPNt1gO484p6DlT7nR0A
ijNTJC+vnEu1YLj5iZcKEPqBAIsZktEdMeHgXWMl1FuCwAYJXwDdXNBJvGFTdVzZ
ybpobgdrKYhcOwvco1rflPfzytF6V40EQbp8bo046QKb2dmZfzJoHXNEciiBX8EY
jeybKkyctuVcMfVrmQDzkdFWFenuUOnoEjveEtGPt2ZBEe9RcM7jEKQdxdb6/Dy4
bt4JDSr0P7qLXM2UpsIFv85iBa9dztbNlMUcPeMUB8AvCZjhfb+GFUs7WNJlJ0i2
Jd/JUD5sTMidi+buKN7ypGS2YTM8HaKKwdxJKTfIUZkpgmow29JYcgbXJu0RBKGh
kYzfbpNaQnxvB+3s9Pb9VPNnqeWWzq/FDPwWplOAnEbcWVmwt7Wuj3zEbfJ5iwaO
Qa+GWMLNNTHFL8PrAeWHAKIJcgGfUQ8H1E5dk9wdTlj4iF3o6hxmh7eQO+fg/V7d
zWKgqG/seekEw/Kz4yrXmrjLNaiKeXxZI3U75rYS9Vp19walfWCCUuGnHY+z+YKs
Gf0sgUKAryqBVG3T+qLGdSezgtonYfb2ufvf+ADZ934rZq33rx51gb77ukKlu5i2
jdmKpcEZ4GHh5MdkXXVafKfKwq4+Oam0/oIdw5JPr59xMqVat6pzIoaoqa9wPvc3
KHkBetBW6gKPK7wzGj0uDIMB6TGfDxZyJ5E3Ah04O7HWbEGUD+OyR8nbuARNuwA3
YeESFCA9gHwj2tQB9TmSGKrsDusKGHlhz6QUXk+4Gk5W2Y6sX/02dnebZXiuCXVB
t2urjq6gaMscdpg20AAPnwK7CRr5CqFb8HNjAzClOf08XGQ+7lHwAygZQ7+LPBeD
1hhuygFMtZOLv5HupeM8LJyYNHR5EQnVazcaD+lxkSGZ8NhVDs0O5mGuBekiSUPP
EZG1P++o5fb6h2GgYd1XXQML/JIgrdIRy6D91ApbLPQ6ZG22u1tVpieTF1EEWrCl
HqD361hTpBBJo8bXndX7rkCIJcMDu4q9PON30EHq72Za2O8VPRwEXL5Yc0il2iOW
BQaPSlr4N6h5ytxwq5yzhqIURASz7vRyYmcKn4rw9GquXAc3Mp1+yXAJb05jnlzY
IOgEGg5kvn6IRwfNJVQ6PdNQnRiycZs2oUVn4PWMTF1XIp4mlchOfIFa7S0zEnq1
13hQFpGwM7RvIBom4X5KQrgqZmzQnkUpsPYRwSTdDb4n8XqTWzmrgqRNhwKNAB6m
t6iZBWmoSsAH8BrYTll/DpeRizsTPhxzRB7yYTPaFMDSVTb2vrCYtRjsrAYC04Eo
PfGcTyHJRiJSCWg4WqD7k3CVlQKNQBlmjLb/5LRH77OeV5txbBoQGjVtK+sAe+xZ
duzapojeU6A5Cf4CTIDeqJiFRiAHkpw0CxuaizWA24AZojeLqBzU9xsOWiVlRH4L
DlY0UcdbRoW1Aden9lA4oB+sGYMZRkZTPebsK6tOZfeo/Uu9KcpDEH7IMcCglLJ1
baLrAq0sMK90zn7b3qw8Io1rwcsxm1dccz3bcIbTSIMvdhnhNKe95ieYyLLghC/f
hsghahU/dNkgeMjZMo2XN5G8/+Uz1cTH7C1kIwztWy4ad+y2/qCcO0SCQjNpWoxt
8/Wp2z6MmHGEc3EZ5ojXDR1QgiEQGrUkZEFBb2eKwUMnCe+P88pZGgLKCGRXat9X
3imQSdGWYhlN92oHKD9qi6Oi0tbSIX8fGK3O+UG5o61pakKOu1OIobpqzVYgxVAT
ml8mYyP6FlhUmqo8Z38AX1Kieyu9eNFacMV4k0rlDUorDD/E9+RLOEpG90PXH18T
ADJehznsz4/30GWiyjBLg7iq/UDOwT38NgTjmmvpVrxG2SV+eKRNtS/z8Z1M3msD
cJHYc+NyR5fauqYParBLPRJ+20euiN8Cqh2FLdmfPxm2pLhrC2f/6wOWfdOedEmp
/cdgJVXu+7i+JlfdjXbQDe47F8ohvqGEMmiMlxpbZlLXJWAkJZmRfQz6J4DvG1Lh
yYTEiTg90pzfs/XraAY69iSu0L4kpkTr3g1Ippp0e5vx19ioRAsV06qleHfpGnWt
/nj3llEnBV3Ug2SLxwfXmGkO52d+jJitOM4HowH+topZbZLLzEE73+i4zz2BURke
Rx0e5WkPnW74RITdF5zL7src+4gGGBJr+I8YVauw98C4NqSZRUaFcw3CXwyjEBax
Lp733COg2kvdsbYfo1D8YfpzzIL3XY6apSZ8Jp1zQe23dtYr4jd5FY3kIH+v32wv
ObVIBFYnyA5csMtwmZRnSLE4pJ6jitnwYeVW6BHtUtp2LzOVzQhtyuD9mwH55r7+
n82vy8WpySt5xDzehRTTkx9irv7LZqQgHZdJ/4FQC/Yf1DpcWnVYkSkuwU+kWwqo
+PMXEo53fvbZM+ojKmWMjgdPLlhvTF5Bro5LAKhq7E6NbGy1eKiODAWQUB/lw0Sw
SbNbkjdkWrwNqfzQPuGzauWd0nfKWX9ZhQObImuQU4b+BDolP7FLC2RQ0uzieYFR
CponHkq7BSbZEx3eGaop47K5rv4hxO08ZBxY8toKa7igmyKyt+NlOgdsnxVSls5f
Vzz9MDejnnIvJhylYa2/9mVYy7h2qcvxhd6yFVJk9Lwac3+TxzoXqUDyJmEoNA3q
h+94XHBs47rr/eZsRLwvyh6wfLRisSE/yhrrtRcOvsEeAz6Wtuud6EwVZkfznak5
YbvtRsU1Vam7OwYgFZ941ZdVDYi1vpowbIw4Yndlxa5IaUYM8kK2cpSr4uDGl9de
IEiXKHPBRs8ozOLnJht1ZWNMsh+9tEUh6+183RqW864SzDlOligwm9fqNYe136f7
uj3JNCAwGihBlQEQ7PWwOoYEyzma0YKgFSovO/3pLFpHHsC6+aNrQoSw5Js+LhsF
PjtjEmwdEU3VYLemh3aBniPthwujrb0W6SKjZBoVXSI3v1GjJJ2sA+v6BjXsqBnb
mL+QMOJZ4qdtspnRNko1BrtpXoBRGYyZUB12NNmxuZ+wGVOtpcg2CxDENgMAyCfA
QP8Bcq9Q9tgmUCEApaUPrE3uVatEOGs2GBe1OsdudiqvUtKTImjsvQQlBZBmLW/1
zv+ZRYw2jrxFmuG3z88vD65/gqW7wqN9PedtX3lBuZBmyy3V2xXeMdj5e7DCVa8y
vmXbkOEuvP7KiNeEALHuWOWPOy0+nPflElzGMX0TB09JyEa3pwQz481gg6ofbt+Z
RbVtyQamjLAtcVUGb/9adcNckxAYN26VMyOR/HGQ3hXqwlT0xxNP3IkUi9PevWRO
q2IMcxGcfA+orncMiSGTW6Sx2zFzZNDiElyUFsefASOa8XSr4mjVY0kcY1Dj4VKV
SWHk/XYmKfvFHUq9r/4dexThGw+tegub6j5uD0nH4/kKQyalNVZiFnkxDdIsI7K3
DczWk/KLYrgqr0/p941A/LjgtUKRQLk895epLPnukqZ+m3CJGbv3u45nc3IvNddj
c65P2ROPPshMpSsTHjozqDiKMAA6zH2g5VDwWyCIJYRumpHYhM9lDVGcuIstvlCp
/hoNKBjJxFwRnUVfYSYufQwhelNn4NpqDNCFcT/uGCfqvSfvN+S8DzmGOrho/1qY
v3AwlKQ/S0/+LIpQcjdW63EASXrWyP7qdIcBjv/7h3ynG60HSOM0tiQjo+KmLvFk
D4j/4B6mbDEaLWh/dtdLSErOP/4j1ecpqgtV5uXek7VVwTUvPfzQSCJz12hXkxRN
IQBPovGU5Q0RMuMtF4I5nvig+r3/UUp0rOHMqonQ6TqTxv1Xy8FDfldMC8UXj65u
c0habwHBCghT/gxdezwKkrKAIoff852oVTFGCwl1J/vapNOuRfAnWR/KX2p2KD6c
8j4Dh9tJehaTvI8vHeofOszF4cZDt22F6MW27kduM4iP12+b2a2zsQuARhE/xJET
/lxFu9C1HKB9sLeNe8/MhxGrHUZzLbefMN/zLue4VcYL5y3hfnNLhpALNYBdbXgh
KGqnn7EkIqWhEfc3No8AhLlHwczUWF0W6jXG9mYm5AAjP5+6gzBpcC/dedLlg6Bb
rb27+3Uw05+kJpimdpjCM3VebCjEVpPwcAFCmH0wbTLQI79c4D+tCL8D3JGtUHGU
IfppKsMUQpydjF28QFYpsvFnYAmactlSW8W6Cm/EpH5y977DOIge3O1fQWBJnT0k
JKlw1JR8PMaMNlIQBJrpUFKMXtRTndgRsOXnGsh4WhhZIjzGwZQYKGRG/53A9ltU
2pVrJVOSodPg+02RKWxpPEQd6d3g5Rj5WKYLa0Sih5Hynpl1+58cM34fpvjddMkT
Icjcwgy2lTo4YsqLGR35UCx5mzofALi+Iyz4eZhbZmuS1AB78KTG333+sby44Oad
lAph3USfFkX3jf8uQZgwPZyUbrQx1BFguxX4zZiRJf0OSBJVxi1y8uA2gTEHzxh+
OFpRc19O4vVwdpzyoUmupUthZ6LCDBpZv5K2GSLea7uY6z3NwepvfTMpjWYXofy6
MBhGSMSj9Nl8rXg9na/rNTdO3sFRokuIoXiRJH3zGQ3dn8gtvLMwSjXn7O9vJO4+
jeQf773vGSMKCYSZ/amBEOGLe7w3s/PbZHnn6Ha+W5L0ussUMWOkXxHSH6/IWdsE
C/r0zNukOwZDf/9Araq+zkGFzFhsr1rrAUc8t2+OmvM1U+/p6sAJlkOimiYq0A1y
W482/i3QDj09C89mpBNmo4ySuGpc6W/XVZ2ASOUK94+v7vMyaj0FC/YpdhYbT48/
wq1uOKd73SbuU5jucNjIe+IK3qQmRRCQ+uFp6kOySOAbJNMNtGXS34eM9BgRHaim
OO6XMbDHEGlByroZa30PpbAh10mkVcwxy6eVCiC4Omo0b7YinvYEFr/CUgE/hG26
QgXoFy6k6Ie3Z03WTGruF7aAsJIo7/EJacVMfz01yxTtr1pFRX4kkzK98GHsZHcw
BwSG7S8++HBipVWzl75eYTgUoV2c7ovT7rEwiurBSi+6sBpSjeT8adWtK0jQtp5m
c+Ku1LTeN5qFpecXXq+kZIFBl27GKQ8E1KVbq5mDOu4Qo17LXhMdPhxnxvuVq9Wa
4kofm59B3hRVOhiovBTcMt55WQw4KqUNRjN/qdh7DzMAiy6lsTQH0aICz7MXJZmy
KBdDZgvEEbrZbmBjcMv3DcKnSrPxh4OFeBwAx37lY2exWb7QUxGjx5IjvD2m7daE
UGkFXq0wl8O7j7MCYbVBaIZ604Q+5zs/7q94tQOyZ9dXcquMkv+XWamSVmlztJLP
80b16SrRFNUbGn9/dyjTGQLEarddlwE2yMsEgwvkEIoTf3NSlSMhj/68aLa5A6ad
y4GsmniWfGKdoOl4cO32dpbj1tcV89H7uXzKmLKT5GVmTgYmksGU0NPmruhZ43Cq
BdFdQ3LAYwP+jZ51WYsLH2sbbkabNpLQ27Dkn1Ks/E/AIJwOgKe4dWUVt5uz/+Mk
mtwmRCJN8ZCDcnl/ZVnE/kg8HmN2NZyoO52DUYCPQGZgRVS6WMUL96dNqPxkRf/a
1ZQN36yqhI6+4xieN/9Ki67M0Yz0MIc/c55QfWrxKgDV6TE0DEwY8z+EOUv+cvC6
ci+Ygu2ZDBKW5dpQMjdAJbpibZBoI8ND0KwNxj8mpzibgP4T9CI7q2ugP0sTn/jw
HQRsXT2C4YT3x6cJXceexfLBtLujY0To6uYduQnn915rPb/8r6BGNtLVkNwXPz6M
wOzYF1J5vOzyKpg0//pzc2HqZ5Hux21/jeYdpZDMcarHI+Jje6LIFvSMr0eCKuTa
6We+rYBqYj3KZC2I3Kyb/t/kFkLQAUBK4k8wpRLqhSv5BGutgKqQ4MWBHpajx8Ob
VLvGNwbUBvQRLuHUBpYYkmh7mldBRYTlg15Sg6BaJRewj5y2gw6vBhmwHuainHZn
zPKBVMsWgXNnFvslgQectixvxXFy2B6lkVEe5gBE4l5SiSOZc5nsUmUWAj242nb6
rZTqVtqkwz7Y9wPD4THch4/jpSV1BngOiO8qsqBKbeFbeflPSRARu0byjFsWwuNE
0kjU2+c2eSnwxUGQf73vVsPevlxk+gw9JHExUtbH6ZD3t3WMNmXgEO98fsn8BqSd
Yr5ndz+iMlmc0SGkJuu3xchQdankWxncfpHGRLhdBgyG4bIV0g2qqE9Rd3KZF0VT
FLjLNS71hWHU1b52pEAstFSytBZJxOcS+YWiwNOL4ppg9FUhUd4sxjMTLlKiTCy8
Nd2djN5PuJ3O+9p78zWbLRkO7wFffaUzwG6CFJ3B3eHa5j1n44SG9Su6snydRdzd
QrjlGosdmNXWiZ2dMZO+GNJzK0QxhuG2FZ4pH/xw3um0QJkwW7+7eto1lbJ8NBn7
s0HF1WYl0hzHJhMLvpitSuSsB8yU2flMAfvPoDWl1ghVDAvJ3nTZKKKAnhsTQMoW
DO20eUcfA1FCRH053iL5Vce6C+M75+VG2CZ30u394KevMMcR18q+8u200UWQC6wl
1V6qdzEDXvm2wM0schlp/QVy77xj0zAPnht88sH/4eW3RWpRDo0YcWzEj+yxKOfe
VDiqzI6/4KBCyieP0blAjzQUzityK+TxVFdvJfd2NlSfw0b8MF5CZCMRrYVyRNnI
bb+B190gjVvSKLDdHaBbTgAC9iiBscfTzwbwvKS0+/kN1tCfHnu8CsETEterhCGD
1IcsNKerdJ4+AvGNT2gerxT0aqopKM8cIEfwQXmUrad3wOUVR7nNr5OxmFQnqiyc
AyAswqyEoUdbPmxHvip/vezOK9xqUUQvU055dG7DcrsttsdalvzR5XGxQJ/oQv0N
CXNDKOXe7q1ZK0b+lVo1ql5HkSBRSoo/ng70YuZlF4vxtW1BXVlGIMExWzT5cup1
PEuuJetxeYqmelh2VzTLjAFojmg+vI5qgE4xxfGaRfqkukX0sdb+ZfWWqOdnd77A
iQUyEDrM9KITZ+8aV8Lpp97GzQE9RdWhUHjxr0vAcjkrjkJd98oj+yISjEEh2Rk2
66UgaSbcq1l9pMtCwK0Y0YEj5Aa/HTpMoMDfuCECtVkMm2I7XYFWh7ibGlHJ72uW
73QhoWlSfyv9/wYUvGsVXrCDiqCN3ubl+KAug2lSnC61lGaZ0nFaQMmUrZajAM00
mSiw9aIFmt0F3t4kG8R1muDejShEPdKTHJ0tY6r80kgCLateRCMrTYwPuXFhD1mq
eNshOMUP5LmxU5GOoHFeyu0B/tvnAprWKiFSO1VRpBZk6aZz0qRJ/tjiFPIDXzx7
Hf6Vdhx98qMfrTIPc4W8yGgkjEbaQgDtXprpEz4JVtfdq4NuH6uNfhlSbZ0Byy4z
chAcjldQdoEoH5/NGlVTQQU9dDnVBHG1ecCTkHOhuVyFbVRNEygO9jksAJbUshJA
MTAh7I9QTP2/TrUOF95tKkFsjnS7YyDb2EfB6SA3Lg/1x79vKLGqu9IhQW39211I
QOvBc7leo8DTiFflUwvTbA6oM7M4mpXEn4vVpt+2gjc6hQANZFvgfTSl5SbAW1Xl
Xu5ZkbTi/mTliMEqfgpNlkYrz1Bs7XsLqVAL8jEsfdA5eGeBR/UxFx3cw6jXTc2G
UTIGimOwcHGH7mgpGKiuk+49FKVzIbm1eSkGzACY8lXGdq7p8LZVg0HFSMgAORN3
Pe/XwouG8eBuWzfPFKU7GDFd1LLV31Prtyn0fSlIyze3DNAKxxUuhK4N49l3Xm0R
8/Xfa8cZQDXK4nPKzcXazqtrw1Ui8HVAZQNTBabihpH2Seulfk6sbh8wnIXiisEI
EbPDGc/nW81ut4W6eGxlDf8tWt3T4XjIF06cfvFqJSgOGk4VlpEzoE3VcHgEQPzj
xIIRZJNmcg7KK/45ivA3Euf3QroZb29WWV076QZLRI78eJRYXogK/DKGQK9HziTf
s40etAagf2sE/dmIxTOXfXS+pWo2SyTkMTcd88Iw1QQWeFvbTXNJ0Nd6gv5r+peQ
A00spaP79cdo4/ykpWUNnLaqVpy3JHY5M8TC8AxxOMPMoF5NwQZ4sAbw81LFrSRF
NdU6km/NDFpZfMvKPPOnEApcNLmLRCV3XPfWmwUlHOKd4QEYpMticq+HdE68SdoM
OBUNSDnLWQDHes8KEQh0DmlhTEL0WvLGCVPE2tVFQHmtcopx/6w8RsV9Y1Bh4dA6
RXZmaAXMNlM8P5aoS08X9cMDEE0bqD1vXB3fwII50Ct/FQ+a9TXBNDMaEGYrLHWx
e9LqPlxxB3kZql4KPslmCaKVHEl2qH3idAKehXxhOoVUkDAZASX94LviQmS3UMk+
WDJwY9a17DI/PcdwPU3HYn4IzTShgru5XdPP99nnhub/mU/o8fdfFutbkSg4P4O0
D2hC0Gr07WjI7Tgdd5PHg7OcDXqKcvnAU7RaCAnqdsDndk+cKSJyp7eB5KefZM6I
fa6Ke1eAbUMzlBbIB25o6UdZJUEFZrQln/hMwFAsIAyditSNEmMwbaeKY4GHGxiU
giipYs3G20s2w/i6Hd5QzufByhss8uLbsBI7+Ghy7Gniv0LsAoaMKk8lFLlhMY3d
67Rh2urETcTvUPD2v3/vno2OB3g2mw46WHQ7DN00+k4nwnina2RcwBp9JqYueRSG
gioG2UsT7YeJppWNIXFzHX7gK9eyzcuDUxChE1OQN/kF0/vYXnKtPGGgUq5F4mA0
zORq9KXJqsB7863fvK8nEEj3RwYq67XSi87iFx7wnf405w3vkcv1hyNfh5sgiJGD
YoXDu/xwb3peEfrcaoCFRXu2f9JXk0lLiDK3dOIQgCoHqWHOpK+MgJi07lZgLXiL
fFJjWYbUQHkp1irpw3V+BiFXw5pfAMQLNLLWLvm4f8efZeZz8sn3VRZ0uN6u87Je
PJJ8wRjVeAsybmj2ZELOhhKxnCc0UKkeHeuJLpuobJo18X+gsds0FNXciRvmsiG4
aY6EFZ2VyzQhFfHjZc3cTD1DkRPPFyQG2Eu/08XFFxbNFWVoUeyMVIivqxXkqu9E
w3l3XsVrDJlE7E2F/bp2X4tgS/vZlu6P5n0eVsteY34dDz+CBTAfU1SYVgAkr6ZS
04/VwJR0kxlUcJ05XSb8sXLDhS7KgH7rBoOmxsz9CrCrxUmW+4SnC1OAF14jUAEJ
NTXnkzmA8FNPclF9LcvDLz9jY7Di/jjtqHGAjolOmpFp26tarwH3/PwZAdQGalbR
Xq5WFKHOKTuAFRhioOMsAfc2Xm+itDZy0+2aUQRrRtUZw1Hpwdoh1t6aD+sayIz1
ETrks8dQ25K/4kLTB7e1aLoB0L6O8vaYOKk5TZlHXT1KU0qopeh0FMMbDKc9j2DY
H6eU0oX/XhgM15YoYOs5+54znK3bq0BdkmhiJ566ODyilyjXYIxhNrG9w4uyG5Iz
xMv1t9hBaGTlNd39gT/VNLwFdXGlTBAVgtyHrxFuMpkBG2ZvGLjOEvVOJuE9lcc+
6BPBJImCRBQoFfjVytiFWNBEA0oN22uZg8o8aKsdL59p7UJ2sm5Sye+bJG5IOa7e
+mtC61qypB5pNzuKc++Avgt3P8NgGU708nGCq4HhfsMFFK38rbj26FSvrSaUQZv3
ju+u8zPG8fCdN+1VL/q9YvQv5yQEKONLB6iqPDtny2A02pDDD1mqNzhm9JLAj3V5
wrsAywoquytu+ghFPS15tk00BHEYaf92mfnoJ0kYKVp7821ozx+DhT4aGgzgLZVV
j2aSkR2aZwk8byY9C3hQtwTyqp0130p6HMoi/GV38plxCuBhCEzEWljyrOWbKhL1
i62Z/iw5m/9ddS20PvvpUOsjG1bRqu+9N5UgnVBZLLwsBTWiiGyh9BV7rlKw0xu8
o1JhSntSMW0JRjpb90lIqRIEDv03WrcgdOudvmPjzdX6+uDxFWxatB0Azy8mdD+s
6beZTznl1UmIDlff6sxOxfdcVVSCfXyRoBjAAmGNOtyb1RmzY0iVdatZROhVdbiT
fpJLqVeqQhPLgxagY0/J+TTCQlrpDQoxB5RlBlVdTg0lFnQywtJpcz/BhJet4uQj
CY9B0Vdv48K5+iLKMkMbvbp6ErfSBpu121Dzg4wgisz1xlWW0mHGADK9nrNgcm/m
I720LyZ/X1mEL564rIxKKKFyeo9a4a58T7ZAn3BLtY1GYldXziI4scZAleTI+7ff
wkpSxFqaZAFEqw0Emk3k/dXCokR3r+Jk5FlaISSSRZ/cDUFvJxcdQFv9bA6mUZJy
3GS9IMr3gHK5WfSO5GhmYxyvUGoCkjk1/DDESKi4qs06Ky4hro8SnykYHdQ+SSd2
XCdHcqas+Wrlkd9H5Mmupr4lcuNxyCQmb/NY6+SVO6ey3uk062KP7l/uQ6r8dkLK
NVUEKLDiImp93jUGdZA5RnMHoV5osXW0nvYugsAfX0/VhS9apvvBDsyV22aBJ9Ti
SkMjYhXEKkinkes+AtmqUMpwBhod+BbxEvjE4CYNWwMnm6vELaDVedjxwFUpoNQ5
C+0mwf0/o0Z8CGr5xjyAwQNi1qxt0/1mXc4bL4DmqlV5dBQyLYMvu7dio9Iw+F3h
QaW2HkLc611Cl3twvbDLbmDsrtPa7GA2k4axJs6L/OugwOLq/oMseqonj0jxpotG
h7WN2aa99bkpO8b1s3B++l7vXhWKohzimFmvFaoEQFAeR9HRHHwHla/C2gwC8fLk
MpIPGVBNkgTZk9psvY0+PYFzce3HlEGVrzcUEkZQLhMzVHpB46iODnQMcQEk6Vbx
NgN12M9UImsGpzC3kMH8nJvPyPDO1NRBszyxZFC9zXOFt2NDYU1lXvAE9DliSrwI
px9XucDfuoa+LgsXxlwXArhw7WHl/5sCRh4zErxQGsjLta56WtYFBq/Yj8G+RBBc
HhnYn+6b/N3J0jRas/Q+DvsqNXK7FUNBKA6v13M3Ams2ntXzsAAC2BZdNZCBABvB
YcpXPd/3o3N+g+z0EajQq4f2rAEj1dnivKKlm8nScxZBA9OnznaprPqxdQnsHke4
na566N/WdnSJvvuIWfpSvCY8CaSSjauGKuh0cq5H4/YQdW93yKoBrlajAowi2v62
calQ4xAYdgJeSlmT3GTGeYORiX9vrP6EqC2VzmImON8y48TLEkqHGI2DzzwbVCes
D2VaNNDNbTrUylB0+4EzJfZmFR7+gxVetTsqcuoyi/7tbkNQGaeInJvpON18YuQd
YohIxfKCORBnzMqcCPrNIcyhxgKG9utZPjyicUHmxh4pBjLn4sX5/d7PGHsDYnAA
dbIH0mCbkttOs8G/pBt/ZxgsjME2HZ/pL30Q1423VMaRpAjI/i/XYiBpnpaGdGyJ
q33u0CDsRysO/JtGCMcmqnCMqCf7NeBmhjstFaxB27GYPO01nf/U92rBAF68+xNT
GDLyppL1eqLjer8qFL89hsYEal7UVaaSzj5cRIQHxrldTT1dyJmrCPvzhdXWO30d
knw6OEoRzlRdtI65FglpJxTcJr7V2TS0G9CzHc44rq3H5gFW2EQ5qhCaf/hdL3O6
lQDefZbLDII02zxdNdBvtMtRnEkcarZV9QvolYnXBXCV6TqIHEenjKu+NvpPRs7q
2WUOork34fX68pc9VE/oC0XvoIy7PCh/thT96qkq9FXCVczN038bu8kj2eQDUHbf
JcVMpMRMXNB2LxE0SwUgq82zCK8ZJV1lPx7Jb4JsSNw/6p1yPNpyhNMMp5xF2FjW
safrMw5tbH9OBwG0M3n+lXLoNznFqHb5Zq9hDpxtuuwLG/0/AL/edKrZe1tBNS9x
Lq4gnuTXv8vtHUIm9faXvYEYrS7ylpW02lHzCEbWc3IkcurR9WlrHEsohQl5LSc/
50SntpjxsbL1ORuPzX9QsYYDUFupIWYogRWi1PhIeDXKiDBQJWbK31prkO2mt+vl
50ES1II+1fafDHgdzKYMrv9qxNBze2LfraTXDoPzvaxM/MSWWp6tnj4cxc2KJskC
nUnWWkp5NtUMXxvDCjCw5PKkTKngMRmeec1owBUBfUPbzgNn5g0vLZRYLhBjPqlD
EtK6MHwsQ4+f3Hmxi8VmMA1Y1xZxOv/ru/Q+LPfkTcWmbF7JmUdxZZ76NQPe8x88
7zxy2XSvujCNXLRIvXhWB5+lQxNPNc20na695wpcbsL8CtY0+TntSMBodF9FcyoT
C8EjVWRxAcfzZHx1pZuUyHxB6FBL//eGgXTXVEvbAaU1xa06yO5jMNABkL14Gyye
k8R7AOy/zeW0tAvmJt7aIUrefo42j7+QWYzbYoFiZ6E19hXR3SvfIchXPc1LRpoY
TfQOhkEohOTEpzrT3Xm6AZ93ivOXPe4kRKofuY/0VQEXJ5yzNKDdLgGYC3z+VloG
bxP3fxjvBe5LX5kxlFqlWyVBwM+/MmMEq2U+ywrhFTXekBinjtQ/xZJFCXGPIhKM
9t2iPhiR0o+MPFB/cD4WkS5RLHseIrvoH3J3EjNn7UOthQ2hPEF7a7AQTQxIXrtd
0PmnHWGiJvdm6fbJnu2APn1/DygdPdwc37GDCCSe1h35kNfBBkhwTomW0Xzd+pVD
ckGzyT8cxknORPvZVIE8u38ngZZdWY/aWU8gHlTRQ48QxqI7c3vk4M2faWeUW+4/
rPHjh4wX23RKEWP3UAgHv2kkzcJUOUyVUfnohAncqnSHfoAxiZlH5DTBsvUdNZoW
gIzIF/5WonirZeYgEqFZ+4g95HQIrq3PS5PXaxhkDMNv4VfQlODVqLUBI0F2KhTb
NwKD5uCs2nFBKeSJRMju4J6MC90PqYbQrs9hOsb1SIdlVvGwTG8dH4h2DvFM69EU
5JAVC6u3/3xekPl/d1sQxDuZLEpUaC856FFpjNsFRYivkM2QSMoXcgmz7u1XIzRD
eQDZ97MoPfZw9lGaanzSoAn0F6RwKhTrFHWR5RvczhHQZewcCM5k7vO/qEBIE+Gy
Ym/0+ZaXlmXYixi5pUDIupzW8V6MTMTiMmB68ocF3QRnzZEOcx/QEV0xh6kCT8hi
+EqGnioh+cOe43J3X4EXN4sZCrDuXxhJHcI+rJDSLQ2lJH2jrjnLkYMgxCfAWmbb
e1rku8TgqEykJyGkQ4JzcVbhmbWFeJi9VCbGTJx5VWaejUXwsKF6RgdR4vnz1G7b
nz/qXd6A7QbIiU5O1EoID0LOMuU2wzEPQc5YFSG0XFd1+/S26b/1gHV4ANdprd72
lYrcwWXLb0HN3UiUf4S6lfXdvALXLx1Txv3EMt0oCLp/rurDFRiGcbnEpTbszF4u
zO1khucyfeMAIpDgj08NkxBEj56EdbdztkalXMjEM2AUbMonb6NaNFu9Sg7quAJb
zXa9hrm6dDgU0Z5w32Irxy0fFjceWzO9pA9o49KCvM9ImvTQCFM9MZ/98Y8jFxt1
uUxDHAdOM5l20SQVkALDvXn1AQeUZ4cC8Mg+Fi6KKYKRNR/bDPL4lk4yRG9np9Pe
CCNJWYhlszJ/36wJS+yP+mb2lp+Zu9LExxn1+ZyyT/vCIL0SvHmQDD3d5Kr6WlKF
FBKH4iVyJsQ1ym1UuEPZ9lN5+ePRjqLi5rZIeWwKCgzfHdFjnykettbnAC8ZR1rN
7CCYhnANF7GQ0tpugos4kpx31WAYc67ARp2THZ/Ak7lYOzIFjhydqqgXx0hQvwfE
KcVi53eBqJA7y8cvdb0HbIsPbFNhjmNs9gszrC/ruhUdAJ9/erIFbKM43t59FPRY
K3KsiDTmd8hgGDe5foqtQ/C/GFZOwFos+P2bYyqRWnm5BVUH3Sgyuw6uz8NdhHtV
hlloDF9Fvt18qCNWtMjBGXwZ8f3sT0lv+lGkJ2L7KcgMidYKzWUSF/69L1O5P8xl
30DQVS+6oSc22TUlL6N0lceHG+eHUgO7QPUxJqCkYi6PPIPEFUXUfaLduwBjq3Xi
wKYTOalDy11/oAvudp8TQuJd2SMMp8ynz5rA+S8njJMr8C+JsKHJmr/XAxb1GBAm
/ENH3DOZj6xtHElBj3XWDNYYI9eqr1CxJ2FVn9LuNyRbUAjyWtpBV4rp3nVz1QA8
OO1T6CMc/ENHlYrkr7B57vFqaaZ1XWF1Eth3mKdNdFQ3jZ7DY8mPBXmfztuW5yeu
ggRzZkWLt8q61741A4cdnGyviBKYRp0qsXp+YY4i7lSmtQjXDocPaiCxeOPwHgEw
keKt/lnD9+4UP93R25hke8jLBDxpW8kIr7gVOSHME9Fs8e4/rob8A2bNIxLU5jwA
LE0T2eQZUcAZKldhdmNFve9H5RpFcj5Nwp9bRgfIcM2HTc43nFSIR6OPkpVARPAt
mYaDSHdicUHK9by0NIukpVvYocTmMsiGNZsxIvoqIkC2ewkblZOAea8m4sei3dBB
PZhFwUyqdRiRY5ovdExS+eFyFEWMq7qm8jAQXXtFUqg24R8N2Tr+9Rc43HePtTxY
yQtf2ZLh1B9aLmBJECete1vhayPC3MYEJwFQAY90fPTkiHGX1x6K0qmnrX8pI1wI
z+7Eybgdyh7MAuO2AhRpHHApk8Q0DMBnxYIhRRylvHhKpgpn+X1PqfYB1kT9NsIA
ofNeCzOSSREls39P2AAb7VukE7H+dsdZzxy/HUoWDdzpX3ELU29CffXeAbzrAMri
G9D/YgC1nEFWXwqE9dbw9G1gwX1R+Au/mUiHqb3ClsqWLe1SwTuzdX6+aSVBU3Xc
Q5Ycf1tW9MSgunTd/5AuGQf/vt2TMHZxpOPlz2btLQbm6HlGGxedYYm21fczFu/f
Qhm6LOB3QD7EtSHT4idyObD0Jc4boX6HeiExoj2iPoKgQEApLlO8kf3RkMdpmFLA
UKHVx3nlst9Lg/V+z0Tfk9fkLsSuPgBK57EG71GPFaxvTcpNMWhLXPsfiFM56bFn
O4jRfc+t5e87XlGpcaPsV1tqcAQYY/BaLPfvrvpXePCHmq/voo4E0J/4ChErC+wf
+XaIHVhf0ZodaHn1gVIoKIgb6zN0lh5PhakBO2UpQ1JS6lkLAk2qzSXsNu3BQWb1
kdQ7i4QXh1usR/yvtXgrBPLjBwl//8b456mOUjK2WOo7iSiFrh4gy0ucXrAPtsDU
tvml7PTByKCUTsZenMfi67JCZknr9s85Aa56OhRPgnO5ItftvEZBIOUMbdngG335
ly1vK1HMKS+uxyONK517cZfpN0oP/ZlqUiEap3asmQxZz5YK+OL6XGQ+rPZbH6hZ
BH5cxglnGr6E0gDOSlrWKWW7Y7KyFdUVmX+cvzLwLtO+J8Z/rXrQfHzA4X0I8Pur
hOqG2leIbnyzMEAfK2QRYxzrKdrwOxvEWh0VI/lnB4mBMl7txmOFo/nrcPgGJzkY
RbDdNvKuLunXljrR0sbXZxvi7zDSK+sFu9BcGWJLWYZ0+hOB8cAECyazLoebbKk4
yD6+pfgh3RiVkYEOWHG47+2u05woI1hAjpw2zDvFS/s9atbV5L2V+e0Dfbqi3ftZ
HRsbx3j2yYDr0REyLqCPbRRoyNSka2z6aU6cIdjXGqOp5edvdOmCJBCfzzE7PSDL
UqIMElUEhVxXkek2PRT6Gnol7ZDHlVQ1N94nfYzOH7MkWNnlAPzESwDVlzpxPTow
loshZE5vwOZt2S1fw0+mT8NFk6zWG0XOwFh/68Id7Dd6QDPc3bvjUULkkFZK8ofe
I1E7J94K4VVcF3BWitjsLxCWEPMQp8I2co9807dO10pXsCR8UyzjvFypmdNFEZuR
J6VJFtLBw+D+RBfADt0Ir3voHA8poMLatGqNTYN3a9Mg18DCMRC+FO0A+ieTWwMv
DxBK/2SVSiozjWqQOPXYESEv8FCrDsFwDQchyb6LSypb+sVBf8Vuszta8oGmzxuf
UooQRmHUa9ZcjTgt1adviOnq2quJb3pWGiA4GWgpAlSX6HCnz0xoeMsaNn36GNVl
bUm8mAYs+ficwEFr1O0bALtdHs5gCdf6uZblNSc/sSUF4p4LEQxRP81G+7IoWuEy
GO1ygL7U2QTQzUMBY/EMH6gKj7PZJ4RWHKnHFvNEtq6nqEm7D4r7DwEq9+UXjmYj
AkCbqv/a9snwUEd2oHpmn+NcLcov2Y3a3ahEpf7cyAY7hM5K5FOGnjtp+An3BnjL
TJFDJZb+f3mHE+LFoHu1gnN6YhLZtnSrMZBzpNXkseRyPsKCRwu/AaGLvMgi0DhY
NIdQNeiSM7+3ja5+sRdljHFEoD0mo4OH1FvN0TBqLbWgp2AOeDfpAGoEhMRp5/qN
pjFEjeXVJkiG41Lx26pxzqDQr1NfVMk9RPb4Vs3rsXMl3U4dRabX9z1RLoYT01cK
veSq29SuFW19g6RUTxYFBOdJOz8Wyj0M/Eia6WcDztpWI/e6YpPEK9ExhSJOzprl
i5pb4zKY9TFdvJYdub9wJ3ovncxDF7xY6Rm+skWmpDGOjIv13lxICwIOQx8dET8U
pGGqRkBpcDynx1FIc+xNVyTJzG7jMJsKh6ks3JkAmfS68PfRSeFqfUQUfMw7uqJ+
iQ0qTCKpzP+z//TyMa1+yJLnGjHFgAjy+to16JWjp91DB4Ff9gxjrvHO5k2X40pj
abSTiQXA4Bz3iiWVR6cNS+q1iZZ/D7q+VL/iVCzJffdoINJMpYbWf/u3fgjia3Hn
bq4umnF2qI2c7aQnc27o4qZOX+tyzkvZYikFUQXOujrXINZngxZTSGa1QNJqdMro
A3TDmShJJioJwkl22hGfX5+JJbzxmi3WgsHZwipZKjeKa5mQii5enlD8pA9vn3ap
r/3rhlr9uPaylzEreUQPTBzDnO82b6zKwnb8ktudSBTtuUaLQbmUn6VoUsYUCg/S
b070bsncxK9doO+39XcmAMU5zc+meJ46nwXD5h0EasvrvfFK4pu+b6d8Gey0hHkR
DUCYy6sIdZXAzY54xCm8dnmtr0lFIL8qIlsPzoRCVrpNPQV9Gcn78vC0f2GYXhId
DkvOBiAouGnetzFkTG3bxqOqFttoXKFo1dEOpnv87Lj/x2D26Azo/N+vAMO749Pq
oOjIs/WjL0DTx5gFjJJUfnmq43ySdCUKWCLa5/Ggc7+JViauvWK8ure4F7AR/1xP
QVz4OO0a5lgBlFTv+KBs4h2Nbk2/in5JQ+nironBGIc9N5iEBFqjTxXwO4ACFz8K
ynAu+4isE9w8dRVT2OeP/KAVx2ffYYC+4u+cbr7QH0q1NXZV8f3ypCvzCL9IRGOE
zkKb8urjcixV2XrYQWYQ2Rrf7pkLUk7K7xo3QsVuUCsoMhYqAY3syXCPEeI9JP+r
2LgQAnJHcJd9/sqKLJUQokrFd7VjxKiS+xRcYrXrSN8K3C/bdvPFF8zAnoZeQuUI
bIM2ak6+yJj8jjE+jwQZYm9wgAjVDmTRJanaCwMcYBKdeL33OueaUvPdoOOzciW3
5DHG1C6wM6esH/ZI7wVjiEU765V99chtH5kBp2YjQPeVPOc2MzKsR2AybXbMctnI
NabVfNu3LLdVsYAua1mWrWGJhydPDCp8Zxy8AjTm5NA+LCfFcIsayeEnfPKOgTML
rxw892EFV8Q+dnzAuVPDq1aEiUVOKs+IHTjXfM4q5qIQ3dNKW1Sy9/jJi5pTQY36
L6ZzsDJug/SjRs7d0Dmb4IFaA99ETQiK2PI4uJ/Qn5k6bFFLC58oxRXmwUv45hrZ
0K41nWuqe5K+9XkCWF0IzqWcC8DYH79CBwWb0IFVSAWMXJ06MBvQBNA7c8CcuRbs
oBlo7YpoSAV5yvQ1ji3cBO8EqY2x2lQlGEGQBeMoC9x9kj2vHM38cinWg/vUqrTk
IrB5MFXAt/9LV0EyJcTRu1Yp7fbpqgyiy2A5v1800w4biNAvv7tTGSvEsh7QYMJz
COhQAHrybLeecRI6Sa8R/4krdGztXztdrlqjzYKFmDDpC2H8NtrWh4quGYyFQLz2
ckkuHot+FiWLklhVhMsdOOlKmAugpz/S/9qasbHO1wp6FGd2g+AjgNNAROfd2QCv
Og9SAoz3ZXqTW/8Lu0fMFgD2crK+QhGdbfRNYoDStvufKqbY+7YucPp6nQtRSrJO
qzkmuXbOiAbxL2c7XujbxxJ0z5EJIheBw2os08APW9qG1T6+7g/f2OYN7vjpTV3W
MjC/djJLjB1sWAwNNtUrOSTrnJm/bVfFtcsVsXPO0g8vdu7rtDPYqqACzTuqAdtR
d/Wbh1/hGwiZj5qNvkoaCVRY0obIGcSvZ5pFGUFJUtJ32Ra7cUSYiPfYnCPrH9fB
rvW5F+XD2OJwkXrZNq78fL2h3TVwAFDx57g4hFnKaa4/LtJb7P2Pr4LDL7Tf4Y/N
xhxmpxhHViYGcF/h2OhuUpt3RBph+RMDbYVqAz1gXQpOcq73OH5ZYiXuT/iJk8eK
vHKqfT9W3hgDKkfill4YkzAVyYBGaRjU6eUIwdtEIcC13q2g7qQax/Nr0Cj4EnQO
40I29wrvJtcURsdi3r4Q6xrX1xhU95lw+MyqvxqQUoMKQ46D/bXolBHLSSNUHQEd
bdpyaOJ7CASy3e38AE6O/xz1hY6OrrpVOrIvgnPjJGmw43r7epLFldbY2jdEoO3f
yiXOuSdKACDTRwHroJeNr31SAZ85MXGPyQnD3rDHZsmtQVLY4tC+XdXwN9LoV4c8
SB6hLqk6q+JoLtwcxwKNB9xc8+VoAsCdSmJfpgnXrwVpesblidt11ZEWHjFWepJD
vW1MA+92JSXmVJTxRxMfJRbEf5a2n3EpsI1A/SUOVRNUSI/HxI+DR+v7XA3vPnZd
CK7Or8biUfYMKaIWmOEJ6y9y3AXdWCLGZaKATE8SvutpKdg/FQM3S38EPhdR1OSr
JPRsRh/FrxbSu/nI9evbgREvD7ZIQogJwDPUNo6JbfYzEo6msenOBPWiadCfN6l+
w+u/A3a4vde0tFXDKjOFMyUIziogIqqQgHkCAG26pOXToNV6xYrATFDCRh8w7UB2
ffsTvCYy5/TceXvNgGgYpj+jpX1rCcj8HwVqHsVbL9TPqQnR8tWHWdOG/WWhHwx/
5pptppWYis7FVLHqvwR2xb09XOnS+gTgd3CW07JO+8PsMvNMtup/rboz7uWiUWDW
A3qn8SKP0aa2lvERBydQydEu7Ku30rtl3i8jA84eRjNz/k5mToEcRvMeh/TonkbT
NtM/QnjPsQmdJwYsQzNjri1qbf85cH/NoCUH2mayngFLUgIgiLRsTrja5mnkfjfk
PWc5nor7VDG2K7aHTW+yBvdt7yQbtNH3HfZAMJFDl+TFEBvE47Q+3z0W9HwfodZ1
dd49f7QoE2IbDpjvCqC+WM409DxZJf5Frcc00l9peINfSMR9yJd9NZGxSodI12iI
5IG6KevGZi5nDp2hypljFRYxOwAAVZ3sQpMaAHnfa5IHC/vXBSS1i5MOUSPF4LoH
PuGde3Cvo84jI8KB3V7XDmzLShZhh5BKZbe6TEaeArs2lmvkUgWEh7BtvfKXIIa8
OVzT5RuYILsR3lwL4IgAS53OMoGGYf4CbikUAXt6j7Mys+Fqe1ArOmc4eFfiLwg0
WoLnvjQ2SmMqingf+LXue+EzsTyifTgiJ1LuoQs8vr0nsrbHx6ybGOjEDwO3d1VY
PKv4oTzCvIzEeI3zejum8YnEmKdFUpxPNxwaWQM3+VKw/AabtZppJ4kbv0HPTNBQ
gxT/tfGEl9/tUVZlXcvFx4P8j7w+oTIVbSt47LQFGyAXueu+UDMZXys39va0ywtc
NdojnnVXc+7UDmUiuUTMe+wjmzD9ihAFtVJVT6y6jfkhqJ8RBl4CeennLTqMuHWj
XKZMu13b/Ik3I8K+Sv0QGKPwhrpy+6N5jPkJ+wPyHA3dpCoudq11GlL9i7Glu7AU
87SQaN9bLplNqlDPgquIwuLpsZjvhAlI9uqan61xkPpKHeqF/3Kha+ngwqxEDapo
190eTmlYG+E6Gwsh0EF/hC3WhPB9qLvbekSl7a1q9gqculmnk+haq7WhlRIhZLgn
zuSsCmwr8yltBOwrmLVYRDhTxnSOw6bm5yxbY16O5DCMHGnh0BOpJ4A9M4v9EvSx
hEFuiwyc5G46ALmXyZKGjI2twSF5jPWbC2h2WB0dHkmJwg0sBBLUTx/Je+HDAKia
kl856y9hk5dvKM3WQIbUKqUzQvKKxaE9hBTNvPT+EykwuAUvl6EtwFIQgRp0b48a
j88xquffLAXQpyDWsyM+5MbgLRwAg4Hj1cZs4tl5tP3956sGc828hq1rhpFG9uni
01WgRPkLXMllZxwaKevKNVvno86WAzfvKiNq5shDQZf+mm+XY1jjSDVurXdvobOz
s9AFB5SD1wi3/M4hL+5oTXqE8OtibkGxi1ZUHw+K9F5RhfUss7Iu6CCAAXwWZL84
Sle2l4gdwDg00iBkGYdLjKjPByIlQVF+cacYTxb1cmtuXN6V9vReNXhHKEh2ifpG
21woSI1tsNzZjFAcyKHjQtT1fpUrgDhfjhluuebKop3WHF9j6joOcqgBW8Pdc0mn
9DGNvy7927p/vGj9jThsGI6XgI96ezcxfyzjjHSUFkaWDZLZOk6/l48Lv9xndSCR
5nv2VVIYS7lsAnG7Kw5KYyTF1wdsYs+TRcRYmubsN5Ikx02oIOyqjnM2ICG4KiNf
cFpbMm07S3+EPad0Q8Cy2CxCbQpTkKS8QGySzGOTP/l4HwrcbjfYlM31Qn4M6dto
oYOdTTffMZl/51sWwckTTBpD84Blo7DHgLXLebcitp/Muo65sjn3Swvda7kT3Ibj
eCMBKNkqe0S4lMh9Gvx5AcxvJf+PMFnRy0flLhJFqVr7r/GYPli/56cXCMIaH++A
hYIo8QINEoHoadgNiFRUjcxK2tXevUm+4MZdWs/07yJkM1cbeZ3rDdrQCdMuayjr
LSuPTC3mR8dPRtdKXM5J4WAg7vrQCwHYWX4m/zd1fZPIH6ko5gOcgA3cpMLexlDy
Wod7LSl4X0cngEyzC2JSFrnm6SxglWgrhQ6bITz18xQrQYUmiy0neZV2Z6f6JCJ+
/YPs3BQS8fNegvwPX3mtcmqjygxu9EEQ2zNoeYwd4PjkTwTDk7xuSNWUJdGTgev6
2cJzdV0YGMOiDHt0o7SmUlMpQitwO7FTNTwN63o+eQEAkcxIbe7C7CxbUg94ZhXF
H+KCwGGMOgkmy16pMb+oyPcmHYVQr8Tt7M+Br4Hssy6uSpcZ9FFOU9U1/ZTAp4zj
PvLsDpempT2HiMIfm/dFEG6VWKAdizG8EexsJw3ATjpdS7I2ASM64tejnaUeg/Zb
+da83MEjwBJ+ydHEphb1mi/bDbrWgBYyEp7C+v1y+MhlWs2wpKCxEX5K0WJjk8XY
nVKEjfxBgyun3htMOfv7n8GtqMiv6bKK9uOgUAi220+RFiXBIaZnzI4aoOfRrs9F
hmAo/ZtR8vnTjWpP+Vb8wnvW1t2CgzfgFflR3tnJSbhjosCDL82LUicfY7uvLA4h
0U5p/77BpU8wkk7ZTETDak5mkibAyn2Oa/mMc1t/WRos/Q3lQnOi6T2nKwdkg09o
fU+N3tQ4Mu2v6o7K3HBBJMUbCG4/SIWz5NR8sCZ2W42Ds0I04roXc1svZBbJfsf4
oHHRiidu+UIS/gF30Tz5Osbhmbd1S7Atte52pXPNUh1e05OyQoDac8gTiBubMpAu
k+T0odPEetsqy4xKSfJKyIGWDmQo+TBoYVZKHU4ZxlksFbO3Mt+UaCb8YZBXrDny
TrnfXT0FEqHB/pmBYnTjHKIKC6ULQXGStjC6g7TvdkWqL1Dd4uXXh8IYzt84MzUe
XFBR9enc3HzdyBe3epBZeUYbGKlntc0icAZPDgIYoHQzywmvl6vGz50FzNBK4f8n
gNS3Ft+sYpQ10ZjL2YVTcOxPRv5brGP69L1Mf9/gabUVH3UGonfmhAPdNf8kmw5C
GJ8y1f4CN+ynTsFmQiSN8nIjk9jUNh/2URIAK8CtR67GxNIU5zRdo3/fTniaFn/4
BalArxxJ0r8EGP4w0p8XklVYBnAh4WN3ZZI3YZB2IH0JgoRz0gn6GodOzLXtMcdj
AJ9WlU1Tu/v/SYKu8YSXKXPSTYOaqN3PoJk/0zItfyomOh/jmQimGomNCKVR/CJt
oKr8r+1ULJ1nMwGlFRJk4FB/9CD3zdV0D2S1LWokx/abv5V22Z8S3XS03Tp6uLbe
3skIwlxENHWKAK19abJyFXA1p71Kwwonu5tyoEcfjHJkjJOMr3YIkHxpcrKCgihX
0qC5rqKgltgA/kCsH0oPd1Kz7tXimwqeOGycPkU7qF2t50OU4/bFipF8dEwrXvp9
hqBZla+USWLW9CvDoA9urAjNpP7ejqzLmSkG/Er0ihvrVA+X5MZQinU1T/zG9FkK
zKTNwyL1ykLYCE8y+1jQ7P5zyVMEVpgmY/cuYkjfm8179c0DvxrHz44ONDdxOOFc
8g9iT4vdTK5ESbSsW8xxHUQeKgGz7sbeQTeeY8gR6BSmYwohxm6tru7iJeRI9tp6
5iPQa7HKQVr3VhFX1iueogQBquFmmGh+pFY2wdnrH1dYJwny4HUtpSPNI6wqIkpE
VDUcD4mldO8IR8+Ns2UAgXMDd3mKnh+XoYpWVZOb2fHSTCXoDwJYr6wNFgOqdqjN
yfZWJz6M1lHYqV+8l0ZRyhPU+MyvTCFFSb5lH2JvnLDDTY6FPvro4eKSww0NjGkV
F3k166mIKCRGgYNeWuB1DbYH/Xb9Onjqel4+KXYcIrHQoSnQaV+FJL4MSL4QprQw
vQlhlUL7J5Guwk7+opLoOkNS8KDesYZEkjv5go3B9OZi+VEXCg9hrivYCGmfC7tY
P0kZknIFjW/sSSM+6QTq+L+Hp1h2qr3hAyDA8Mulff5+mkceZw1K5VONYAIo8zdk
RyIeb7QvtZ7aET/MiXSwAOP8Ex585S1hV8jY3ZveWdce6TateoO1lEgmPX96XHjd
IXOWTuPdxQZRCGFZAETifrzV93I3FXL/+w/IaRbaLNxiCh+Y+tE+0LVvAkPgxp+D
eYWmjb9KKWnJfZMvL36DE21BpWoGDcOFhe6vb/NbDWE0a4tkdJZDgR7yOA+lvYRI
nnj3bi8sVUZsuzwtKE+7ReNQXlnpP4MNUwc8mcRiljl8n8esqOcqmbxvf97dvqjD
HPI/cJHcoJ1fW7mJNMfieAJauN3p7p5TgMxGtEdrNT/wdja5P4/q/4nSiMNKDdoj
UbaWnMsqBDJloCXqy0QHCxCYPlnwj2Tgg63g6DbNHGHJvWA9acF8KMu/XOXyJ3BL
2XD8h8bKAI++8NVqfnAtQVMatcdbyxiDyvIGhaH3ro8sBmOkFkgBcj2eKMHgXxax
ilpOCnOsC4AeVoUspMgVeqq1Jm2dM7W42EUqys+DrodOznP6Wzr6BIxe/Yz+H84C
xD+FYu0MI5G45OR5dhwcglzkRBs2XXBedUlZTdURLyjpwnOHHc/a4jxMyrsnrk3n
NEpDfich+7pFylfANcQMEHLfXCC74VLlBbYJ7BARPxSUKefaSWv6INN0NhkkFSDK
e1Tl1lWvFS/K+W/5UB9rsYL/dq69DrmvzXSqmOwbnv9mcOJ0kn2+41t7TZbCww1W
ax4kekciMbZLjzmyFCfFZWOW0AsZcereDWEv48PhYeJ5ODQ425LAhV/slG5gIdZ/
zeMA2PAe8NwRwOrIaAhfgVLxeHpEvlMKK9l75SHz7yQxbuP9aWwlJY6IzdrMjr72
Dd6LLAexdehWFpvZS24PNL4f1Nr9ei2POmepeXhiUf7/CUj2uHvK5IUhScQnoMhA
FKbQ+NhYvHDFRGDs5VDNSnPrUxaC6uTszc04To0eGmDAid5Ry7B76kN6+/X1oQgx
eDMuRdF4KGPg4Sl7jLGkK1s5DpoAtGRKLOjoYxTOAB07mL4RRXU8EaJjLZLBwzsb
RjukygxjiOZOFDtbmPbHC/3CZ81lzvJq8i4KGuxQbwXVJbKWyHZ4SuPKVEPlJFfi
Ign5qimbjC0K9LyOapzJ4JSKEKqb24XL/maOelwhPYlF/E7RbDkfkdWvb2Z9h0qt
rNNo8oXmruw7rMaXy+lRCPP4pC8fDvpHM29cTnIE17LsVmYv2rg4Djf4mP+Hf2+D
3VgDCwjxJBVC2l4TRRfcAJposVVocvbkPxmvk/tpPhzxldzzkCyY8a0p1F3s8eRr
x/AX106NL0bYFmFbqfjqb0Nzbj1VAqs3ImvIBOyIHxOOzBo8k2NEcVnF9wDzwpvN
4Ygm2QU6LHk4X7W3LgHdA4Ls9HRZ5Wan8JasGvP0pOoHBZxHDjyK7uahLGWqZSha
Le2IZn98whofnCYJ/lu6wutPj0jrsyAq8vTmEIvkdcQBd8in0u+nFcqJBj/0wr/b
/QJJ2C5FLWbqZHulA/S8Scm3SpHRy5RVpzz6YGsCDfxSvin15nQBfqjNwK7N2zIc
up0qccwg29xUm6qDUAmdmGbc5jrAkSaslCPeuJzMkvPQCnXdaOK4k4bOKTe0CI/4
voKUBCAFRY+TQWOSTREfC1oclH8fNJXWRKusq1cMMCRe6w96ZNXHLoO+VVovGr9y
9MySuCrVMSPf//XK2Fz/rXDsu7OKHUkVnjxNBHnob7rktRupdJBtzDaS0+oyG47V
EBzxsZG0eM5sCrBNwQB4t6KaQJvU7/QTYPsihhmr6Tn6c2sM7h5XWW5+OyQqvpUN
6u2fFPU7WgR26YAeo/Gq+T+z6G4TBR7YuRjCT4/JWBKzx6f9C+Go/2f6mSmwBs85
aImr7jzkYP43m4gayFx7QwgqB1FzxU2kYRlaE6Kl2Oh2Z4Ff83c926sGYajneAlx
i4csZV43Zi97Y7jpmHuppwJ555xUKx6deHSDgqAoTu2KoGlsfMdDcr8qL+A3RScv
sOKyNyfsism2P+pV3b4SaCksn+QiJ1C4I0Ar0jCADtDgvlqvFkZEArKP59XS+YEb
Z16ELtUV+Ar+4JbzcBC2hiigiDwHaYNDvXSCQ0ZuxP0gxauujmbfGY25RWZm+sbZ
MEmUaqUstrbDRbs5i2PiTBAdbD9vBs1zOh6Hr+qRkuj7j4itqCoXknDEyGsXdgJr
3qVGGaTY1icea8u4rEA2RJnUpBNbmsVVZQ0uOZC14jzHbtadABVpNyIjVFZ1mkbV
ehQwaEZPMqvnWv5xCpm+2PZGqofdiz/qMc2Rv/Zvq2/+jG1yun788wIMRJ3msWZA
Fs7o0DLZMuNyFnjetZ/HwwsunqKPo2g/6XdM/8k+xfGAxF1eAh7QoNUzCFSLTKAj
6CqCl2MfY0JQkKSDmS7sh0dp/za5REYLLkEKXqH2Qy7rflciUioA7dTuVNvU+BHb
yV+ORtNPrj4ejfWb343/yNmmsF8/sDx3XGBCBXmMjA+iFw+Rw4S84RQ5BKVHQlx9
pPfZD1BLme0m+nnHj5QhXRSsmRLwkUhrNcUWSYfLQZuPEJQpafxTTH5r7V6Ud48l
lWZRe6nBMegCZb8FjlclHyE8whQd6qWD6lm+HPjMDpTLs8HwkTN1vhr4GK8UEGBW
sVF9neq4xrOjE2F6yiolAh0WuunYZUTPmADb+3K0i8fcKJKA8lqK2Sb9o45EwlHr
nyH0TI0eWp49bkCBUTFVvrQRP8aVIApRMQCViTxMKWH2wH3sLMwYKGo7Cj//MgnA
b9LFswiBNtHBWq/jd84otaZtmAHpkm4Wv5PJdLEFD0j3HhxKiBC0NbwyQaimXkws
L0tZW0QAUMA+Rns8OLVRBiSgdvO5TVbsKJxxMv/LNCjEH/3GGklB104LUyIDDOR5
COo+99d8PPRfefv7DCtxfDubjB7/U67dMZTHlMilOuErl5CMIpY4NcgPZiX4TfLT
2blyzf1Vncav8WT5I5GkxCBgZrC6S5SqeZiNyXz1hBdc8dZ5nj3VEd7MqzXMr6Md
zJ1ICHd7LcK+lUwmiHOlhdEn/Cc/bCdJ+kO6fKBwSuSRahoMIbdOpBmD3zQKEqac
DXmQN7gkfX5IYOomyS+jA2+jOo2u+GfB7ISvyke8Hk3seX1pF1sUhDRBkNAETQwO
IE0sshKDgixFMVTbE9g/aTV4cOIOSqeiJ7Q9BEi1otGONa8cgjyC4CLi6/IOxXLF
XF/qbH9FVxaM3mJS4tUQ/7VvXfL1e6tJ9d6dzeI4jMRlSMTevpCmc141PPqDhwyB
LFmw63XRwzNgGhB25du5F0RaY8PGKGIklE+pQTUHuxWXCuA3FO2paG645NRi3jlZ
wdKG6Mo+EmD+UWyssRQvyUF+/vS1OqMHCD//s+59y4S+BaY6YHaqqPsQgUdu2C4q
ojFwYFAQRIe69mxPPx7SERdCGss5p188tZuDH3Hp9NA0fNHrRoUfUrjn/zklfxtR
saqhEUIccLwQO6qJH8hhxbzsl6agM6XbHk/g4ywMAdzzcR32iMEoAWARTTq0oNVB
fFjRmBVHJEIjKPxqjX7oQKavDCAGuUaARsFS5Oy4aokarDlze8lPzhrTSEJxAKVZ
/S+uuKxCY4yODw7Uqi/eeJO098mlQsWf5HiOB68oa8DqNSrwUAlxyug0DHfOB5vG
deEJ/Rtz3zDwMm72Lm1CuKTADPz5Jem4r+wJAS5EtOixRp3umpzljmy5ak4njPEV
3nYNZddgajXpdp46QCRZoJeuHAipSPyGiu23L78eCaXUkUP+I5MQ+HW5nL9O1HGe
kqYjgrSTKQ55asNIlKWFZYzTEqEep03yI3aG0F1p5pgeLj1OdKr3X1twEc63mkb9
VWCsx8eoWi0C4vkyu10oJ7Jopt03SwxkTH2/ct4rLduZQPl56PiW+LT4sy1lt43i
OLjkuHdhNvcbk3Zb8vDo22hd3SnkZ6E1/FnsVZZPpKcEiGmH8r1DTxBRUsCYQ78M
EBpDBb+dSsrEsvbI3EsHEwat2zEp99f8BqiwXq+t1X6Uvkq8cLIb35o1v82UU3L+
Vvu9g3fncS9HhtMNzYe4f4b9t8cHB7I5hll2uNOUvxxeWpvv0HkXrl0VNO/XHfz/
f3Rrgei4elWQyGleQBVJxgwnbHGSg4VlQrVQNmyhj+Hr2NRtUdwNtkvV7CoqW7Pl
VojecWK1z2MkWYPaMfxaBs30dOFhDMFpD7Fz/MVNtZaBZ+bdWwJEVbuCy3x+jLmf
oMv9aSiqlG4oZLTv2dxkyEh7wsK5tLz9lhj+uCP6SeCTgYXOH8b8Z1cYn/J6HjsT
T8r0XMcDE0/rPOqviFnPzup3SrNBxikGbJWHzw0IuJc73/qzRP0m2rjWqjt7GBNs
uOIJnH1sQKTr/uY0sWYJjIKIwU2A2rI9YxJCJdqhHBt5FsMUE51e8PqVHlRLBfpc
eJf/60Pm39iSRzhYlpL+m8R5G7xfb+t0BURpuBumfHQJK/FJq2Zm2Nr+UGVjZjaI
1Pzsq0NuLDdUBl0avuM6juZDUEQrmE56C9bJFM6ZBt6wKda5lt7mMnAIDeczg3EL
3kChElOhQDGWezZ+VV7l0+5HamzavFgm3qWLBqUTXl1wDp/CL0+MoNut670h70j9
g4/o9i7IBiRVwNIH2VZrJEV3T8To3XwHa+tjKgrFmj8J26+nKAXTqAiJCAALBcp9
6fTFyjUgurFWaKXO7GLqJik5eZ91l4gjRC0bJe9QactSNSntGstKzvyFfC00Fgzr
gdV0lrcvGMONYvPQx9a+IgVH1ylPe9P6yorCqxQw41AqMw0OJhxdrib1BenZqjuZ
Xu9vX5aXDNm4mJ964Yl3OwH44BXA/2AujGNY7J+yQKR/v709d6NHZG7Vu1ZYvc90
u07zxyOal72BASpvHqW9gVCKJGH0SJeEGaqhq9j94MRqnz/2d6mOJuDWV31QRIyI
swMRcCOaWVH8k5cq0IhgfJsrDlvtWC4PmJQrUnUM+44fEG7KYoq/VpKmo3biyss3
C7vEPimbM/z51xbo29+7OrTA5CPrHxiRZGKRlVctClnVu4K1rgIH4g4rdFfI0j7D
stDODeYc1vjXsr0T3HQ1wwJIl7/Q1G2O7EYENK8/WO7oiTt4hmwsmJnWZbhQ0Lzs
b2kk6aJP/UxKjC3Fq885q/M1CuYD8G08aHlW1QeDP3Yp5uPPXY4c20ECh/oermbV
tzgOrbI2IGKxs86nNgm+ZFV8mCMaWYDRSUzzrn41EACKz1FMvw2ZUVfsR2FTibSc
/p0GY/W/nS7m/FRsqkYyHknBSYqfoxbb+5T/dziYrhZlN6p1w1p6rrhZ8LA2h5Pw
0L/KW1EhsfUi9iz2mOFCn1aM88ZDUp4duNxwFcY4S9EBpHjXD/HJpfPQGPl23mB7
xfsPlHyZyfS4Nm2rwzaHYduP7qeHG9qzjF3QYn218akaSrqWgyFKeDZP1xkxo9Ru
YXUiM/HkEeqqqOcW6o76Ok92qfzGRK+q4K70VH+2V0cdNhadLmjXzsJLqaZfMt4G
lIJE0kly0JPRaUipW6JYuh+tjNAR4kFcHit13RZ3xFo99YjwTgvfOjmDH2la8keh
vhpbmid+/ozCTyjS9X9XtGcbQYVNXURJa+VlFjiogMi7mByOvf2K0UdIEca35kZ1
e2FZUVkXK2t1izVVSjoYgZlQciHyl8fPjpEtZjlUemwp+e3FJy6ai/HnjBx5Q4lx
/rpk5yfEN0uMrKqHx8neBmDBZEpBTan/VAwiRjA5iOXA5jKJ6V4RRty0H3cljat0
oK6rk3gyKePcuUS9KSiy33v2BmBnTaqrwtFUHCX877zIPo17V/SqPPsFtPAhTwa2
aOYau65JXHTs1PZ0PrmTqu0HNc21I2czBWQFbbP4LluW32silTAPRVwCG6pdyQql
UJF169siTC3K5AYehjdlBIAOgCqi/BtQ4Rth50U+ZelqmjmxsRfTvy5BFygFIjO+
tHfqV3lwx5jBEF8bPoFh5NeBlJookRw95456pd8Ngzg8FgeH5DCnVQ3pFL3ZxPlI
bA8zq6TdObx7Hlm0i6cPEJ2aGgTQKu9m8Xw/d1I4tdD3QWxmrdewh7eulYb5LlnC
fci2knp2y6F8f6pixYHIja9BnDUNy1ySGOnKm8L+R2gLQ88/noG3OKUjIHma7hBe
LgzKS15VROlwUXbdS1J3zoGM+56LlR2fohVKVpHGiH8vVq/VKKtt2l5knOr2+sLt
zMqAA1nAn7Vgz3o+99lRA3aCMhfRexKJFBgQ7j4Jzegsj6b7fGglwgVXL9ug6ACu
ARLrEv8rIntYIytMq9wlz8Gno4i4oDJkV+pOmsYOfhAwpZ1/SLzKhj4A3iEyvxQr
SoEB7mX4ad023CGE4gcVng+telZt3ZFoXrALshGMq2ZCXah1F4MlyHqJfCKZcYm0
NLUzGXfwc0HJyoTipeeckJBq5XscFZ2HCyEpogH+rk5+WWXfQHfRTSqy0bv7GGyJ
Ul7vECKyhlqDufdYvFRBXN6fBijqTMNPIPMU2Bo91vIFWF7Ir8WcjWzlnJJaHHwT
tGDfKffYR2g055UciqNcyY8Ot6Jdc668/EMPQVKGbf+o+GueF/tcTOUcxeqEQNj/
MtlwmL1O8G9GdDGoRMWpiUkWsBdO8fuCEFQ6U/1YXdzQd6i5AamrNL1Jd8ZjgQNS
nq2PQN516cGCYRP+TW3CbuPJo4E54iXWqZUvSdUc4bAJn0Mc9AbwnAK9YTG5d0Lp
ukfEBGoHlUV8s3pVQubm/CL99qy/N424ES70E73PUjrCB82Fm5BLGPGMSgtA8RT/
GYSnmZ99Fv8glDvKWrvkvNylc3KgYX+qSV2F+OjSqJG2n6O0HJ8mWuqnEtAKIhiJ
lRgMotwTrl1FtF0h0pYQA7xWhO5CE3gq7bqO1zCtlEO/WM9ltE4PDr2IWhJLGcp8
dXkKlbj6oEL3XVTlmrJzXeNJQxE8zyMEWq7JtDq1g9Gb1crcwOgQ1hUnpW4iQl3P
m7J09jVZoSVi8kPZ26o/iRxVioiY3olXq31QWV0Kddrve8vCwQiIYt9JdVxwm+nk
hCAISEYspcnQNqSGLCLcyTm9RaRoLvHnM6s1lJ7RT+LZMOhMR6+bXREnnMTDXIqg
Y/ARJ1HbtfSnebaEbo2pKzVSUP+8W2jvlzP4pfYicuUlJnEJPR2tjKaa/iO/UtlW
h2e0+JjBID7OUOCSIY6R4aY5P5Jgfj0ZRn3y3uZkqpEa7vAaiNMYKkdrHclchnxJ
/vGSCfrUBMG2I8oW+xkhDOx8Rm7AFEuV1qQnGecbHm52RZVlQCwltzDgP2y+UiYQ
lVzFO/z5JzkKayo3vdoyKIgkC0h7GtvyJokRuEb45c7lQvRDRVYOmMOtE+CgKse9
m7gJYbYoHyghWiXSq4PIAI8rgKImFW3UGwA4GexWwGshzn43pjznzZxSLvM02yLe
zbMklF5ES7w+fgCMhB0XE3SpM+dNsC3o+YVWKyiWCXLn4dLG2SfrOlSVnSbtKORi
JY5Ic5M/9LaiFo4xAH5Mqoy8/PaS3xda9Am7Hgsz9TtMCi5raac8LLiE1XpQHgSh
IJ/47zo6AnDiEUngcOPDtSl99qA8yBOzR3QKtTjtJmiElSmzfBw7w07Sn5UnTRSY
MWOhEJUbx41Tl7gaXJvOQBr2hAN6mzCaeLxM8W4kBiAw4sS6i7hlJMM4GP2NpmxO
flB/TI9kAiygLL3AZEx7OAjqXiNMFkafJ1YxZKD89oR/tBIxax2/whmweiwa0Eyg
69/dikHijRHk336WsJ5I2IJ5E7NIdtlvi3ey13zU79xrJ1GTddsyqGRhUU8tjB3K
fW1fODwVOdVwoD1/9KCIhT3tBRMD35q7rYkASDqp14cv7MQpUz4pGKbiAQZ/Af+X
MoB1wuU/oBCXbw7kbCaAObyHfO6wfeHBW/tpPWy4HDItvnn8LnTUkQM+abTkQjwd
piOsnsdFyLv8rqxVuY4PP8yMab8aQmAMZHAWRvaxswhqdq0MHGaQWvnYKnGJUSct
Hi6R7LS+hdXfEg8dfo9AfctM4tlSEh1g8mla7l804CFS7edUOA/YZ9MwdUSmpxiF
6aJ1R58dOmJH0pg29wSq99Z2FGKLQ8xVvxfzpjajBjONFKKTNs3jibauWEJ3dj7X
H25VcICrTaJ3d2feTYrjWWd1OWPSYViOk2gbUIDldpzguTCN7guv3k6mLwwDNzkb
Ev3J7X7B1eY6Yz1/2mRQ2d3fW1Co+XjieGGA9WheSKTTQPpIFg6fuFG3tihKScol
1XDnn8FRxmv2IbYKjJqvQhevdKCS+RLQqZS9rElMuZT3Aj/njVcpildhSgCwCAO7
Xhq1DWZLO3rTMowszTSLJzWBNPNXNNg5l15bsX2g1LWffzYzDvIpgIB7w32RRMpO
KZ44AuLUaj0JbQNUETXySGPuQbK1h2sCkn3w62mXfe2mMIU2fEEouyuKyFQEdx1H
azCAtfoTOBFaP2PD5A7zH/SqzcHmS46G4m/SfcERCxWjICvxztHQSy1xewESgGMK
zeERK5g/pCrjsF6HpylNFxRBdAbPAif6CMK3db2hScSUR6mbmEKytpJ7/h/P7g1M
z8Led2d1L5UCn5aRRwe7U63Bfz9FRt1paWU+p1nVfOkHHZOXKHJ9HzTGP2Gcnycs
XKV/2/8FdWwDdrORRxI9AoZ1t/qureJNC3FEQ9Iw4yGUODo9ppeW+6CVIPAsVpYl
jQKdL/wc8HJXHYCrq+WgCVtpIQVOoJ6CR7dj8g/1MAgvyzcGWsXeFw6ynISUDdr2
LaayySWtYlGU88HKWjbS5VLh663HdnsEVX5VVTpdjnjT8Fl0XKYIznvRuux5ouOQ
tGSDWMyemO0/ygWdCh6e+qjm6KzpLrsE81IlHoSwib7ycI+YoERmxxsCBktL0HYg
Vx+N9WaR6q06a4byrm2QAvxbJ9qE9ppB/tuEWLMN3S3p4AAuXkUJZZQkraq3/0OF
wqJ3uxaRy/ONpXJW8BTJDcEBgfAPPMVK0x3wVKDUTwyYfU1wW6IuosDL77iOnI5E
L7uzyIM2nLE0NEZvLw9EXFhe5RabXNkqSEJI+q91tIri4ktuN+SDre9h0VqqlYsb
P/iyENHeEA2sPGd3kmUVU/6zPaEmwWb12oZhU3wMAkmH9Fi68zfQZYHveYsIWkTF
zr8RtgaZjJvj102O1+k1v0xUd8yKx2t5r4LvQk+EviZp860Y//q2Bt8Uob51Q6k0
+RdliPvPc3y3KJhpuBTgH5Uoa/Glg0So+DN3ks0A1wGOCQYaiPhY8xf9UgmUGXtV
Uu3nJVuW5W6RDwuOkXk+KUj8kENW6t/1I9A1rQrKRLPLZGfWFHh/X/gs4lVEn0xo
uB9XkuUy55MFJxs3lvBnAYHgMo0phrrfpgWOvBzSGvmSU06mELVJseHZBuAF28om
CS1cuG2EGAEFJ/UrFH8Qktqya4WXzoymp6FutdtH1B0EniUC+utztW0hZbuPsNFR
cuN7IkH+s/PxhLThYAQ11XG/4xVrn0PjfWsmBJzVYS/b0pMBZeHc3gM1U7DgM3kz
I71buNX6jDtBLX/56f+VLm5mUdSuM8LAX8mTOVxC3o8heXHwi8+EMfO4rpeu22vl
fZ5YrAh+LIvt/CBX8IDqcRJDvj67gkKMUi/eG3xjU6i6IldjMIIjKDtlX1CXFChe
TUvQWEW7inWZM/AgZfpFymmOe9pw+0AQhIhefJs/xUZr9t/oYB311qIOIWhSGD25
haRCEXcQIm7xzk/9plRqpj58iLOGcBfswzVCjUqxxxboV1/AB+Pdu6Mw94yOhZgA
5qH3s5CmL6iqE0sHWnac6Uui6zQxhlXUoZ33+7s5QwXfY/nspY/1reFROGxamb4X
b3KYOCz+ry1zHLQmqPW2AyAXGlNo+nxlaifOjDz/dUrpKZNMaze2w51fHOV0w3aC
QzlwEt8gZU2Zyb2AAiYK8+lo2QvjoheHDF7S3jEn4ZJrTmtqfje8nSvilnxcuo22
977Ea2hmi4MK1tD+gS37uVgTCcmA3UY9Zy+bVyn1CK2RiLxTGcVxfQHwLVAIjnLH
onRpqe/D1oNUnQMN2pyh/5B8QRbeFnzDbQJ5e1fyuQP6t+KMsCGvN2+Ryn5yy16R
65rjMYohSyMOQuRxMEumsV3zYk4SOi9jzvkIOBCuajj+ZrgNQeVWTeyHv01yyGLk
MIC4mvcNFH9L9GRrFCmXHq80OcKU3olV1a8j2oX6UEWrWPbOfiLM0pNDkl7vzNro
J4gXCjlPyL3XyvTYLubwZT/fyMW2EQRb+IWZHrV+F9xkVpdh9ZSoCdw4vw8/J+Lt
iWsqmR1IpP/m5rz37tySRXpT8hjy6Vvpn78IqoWt30jxgO1l1Eci4SV1d/YzaBfh
UrCbRd7Z1pVci3OUgbODmygxW8e77+O4gEYfX6mk/XTgwOhDcdoV+fUWDOw2FdvG
md9LCgK3HXKszegnNewCUAWeG2rS8qYQFkv0506IwHnNhmDDqpmHEU+N1u9T71Ql
CQS4OgFaePt25A+nBfd4BQnJP6ZX3goQ7bR18wrroNqKed8jivveXtSFspDxDWGT
qXsQP5aJ7m8Q4NK13wJgVvOcfkCc0fT3e7MuaLRpSKkd22wTRke/7DzZFW6sN6R9
ZaTDRee3cyDIFV4wL1XaiF2fvj+DjdWWws1+yMoziMlI3Qw8bF+LInpMEeDPAkG5
yYUr7YVLCUWpQNqn9ZN7SRbgKgzlSdxBmRZY7/OBBLBBvUAUgWTusyV6lsqvLl14
IOUipZMh6Kth6Ak2BYvRIftFmMk/IGvkzn30BIy+JZMZ/e+tKerXNYIhKRcRGuHH
GPNlRsCNX/8GkHuepfh6YD8C62DsFMIfIMlwvnzrvfr/fG0ZTmF89RZkmWVx6SRS
PqeUWadE89y/qXgztFalcKh4SObc+UJNA3vNMzXFv69Z87zgqYvvHrJk0z3dZGv1
E20sHpCwI7CPKhlMqTa9kNXyRNwNdUezA32+XW4uodXqrQkd3P2t1IIw0uVFPSWd
8vCSfMf6X6YmEGI5kDaIRsG/t4OjEufqq1EXyljRaVCjF0QVe7IYzSHPHlwKMdij
sWIrA9KbDK02gQzDUkuLEVxLUUSuhaDKQSypKx6OCxW2oraKXB2bfsp2G5e9lH6l
E54WFuxw6F4mGX7cOgo9s5ArtFeVD1uJk1BYtOBeDRZXhevzRpNi1tbxMcDVd00i
1OZ1IzaqsAgC+Lrt4Fw0xXlJ8tdaiv1xUExT3OUti84eBZQ0BmI4MZWx3PXVRDrt
VCuaFQTQ7W426U31H7dhd2rnvyyi8v+x+mZVxfKV1h19khWmRouEIbYoFJxGnEOz
Rgvh4cQzJUD/18zP/KNNVJSfLEI7m/xsHL5U24PpKY+ig16KK/ZOHQkLujMjWCux
ciLkrDycOLZx3ibCXVuNK2v9HifxbK3ZZCs2kUJ2XWhYZlrZGHG7nbAVFIXE4PgQ
NVJhB3Ke1gE2COhq/NSpv22olZ2mmL0QjU5O3cTI4U48lFskmXSCroswJLCcz8cj
W5nfsm2lFxOXpomVBC+mKhuAF6ooiOEbJvU/PTi2zvXV8quO9G1l+NivqmhT2XyX
oauL/M1+awlznGKHkc9CP/tbWEM4NQiLTqoLv2xVrARKVDH/YJyd4uYd8yxyXAa2
XaNvB6IpmDGZi9rXq/21bR+inc8/bD+lFJlqgapiHjaDw0EOuVekF9R/8uknvvu7
g/w97OB+HYX5aqjHA2+kqlhBoWZxXI73YSYk1qyhsDUxkRcdVSWdz9qpqnhSWgd0
Eiq9ytFFTSh6C2uNzn/qgAi1cU80zkSwSmDZ5WvbHeyZt36MCHrxBJtt5+Kgj+Fx
idqs2o+TB+gtpjFgJxHt6JuV+ykYYVpra/6nleJdIvnTNvkIyl9SR/I3w04KF/DK
rcWPBXsXXSuuW7PeIlvTE6AZc0uTF40p6kNGyHDb5Yfec+uWxr5sqD5Nx0CExIGZ
f2RomvWiIVnJRvdehCkuUa56CD9PkgGy33Q8lK1RRN6xZ9RpLoEXSoEK/CnUF35l
hVhKJzNzYWwslPOC8ygYjk5FC4ghkpvHm0RqlQK1Twzbhitjpc4QhFZsHdv9hZw9
PPYhwGOYCXfOSrslq6DyvVIvfwX8Tbc1saUSLHFG0sG40NMi5P+2YtyvL0V2lqqW
PjeqfSm8YnDsgSEVuyqaL9anI1Lbg/tT3OFCRQ2Yn34D7I3yzfrAFWTdCYCE4MeE
Zl7D2qum16Gf8v0uUSGOGosoRST1G9jvxItYZcpePWo/y0cIvsU2RcUs+TRAXcDG
Pqz/WCsqRRNrdC1P3XAKuM8SOi/tjb0HDy/yzO0vzqwBAJrw7RP1N9yYFI8c2L0G
Q14Uzh5MOz7WCgEBP/4lGbxoueeQSVgt94dN9tQ70FTRekmYWF+kdiCalfpYAK1E
ODSC2ii6g1muiu8SgqA4IqADjgSDxmTWh86UKWcVns7XSrbI501OWmECz9CbWGRm
SxruaiDs/TXSteyGU5mZOmOIm5u66KICZtycDNxLbajDmfnpDoVgvojzYw88vOcy
JuEsytma6+JlmlF1WNp7nFh+UuV6nbJcG3bgPrqcA6TNzHYA5dAfCKM85hH6sX1F
LOW4dU+mZeow7faluvnjIQhjKEVdaeIiRShju8yEkvKNc4iXNpJkpd5gKQIepyPl
Vkb/gRfJXfU1oEKYOpjOpGD8iANkmKRo9stjpxmUpSu49/4wz+UYvT87730T6RG6
yd6ivNpPYI9uv1w8sKZ6RrD895+KUqY7shMGjk03EmdoDT3fMshpNg4WlDUi1+d+
zdxigCvyPfQQ5hwjF4FzLjePQdAlFGsyi8VRFP7qDYyN2ccrTVs/Xkaa/W9w75tt
p+FCwD+V0oqeypaGOhccol3We8W3zyGqCbNSRex0zT8xm6uWDasR4eXjDJO4MRIc
4mA7oZqtRBMPSTB86G+bfBwBgZm5ZovUbYCzgJR6ruR8mwo092ZYMWfmRADYP0oF
/1CILvPWUjpEetcFjEJbJb50xeuYsBrWNLweyh3k5czKqmm6tTb/YKDdDgxmQwsu
B5RV90kQQhiRAvlq0cQ0hekTUjaoEnZMYiSqt+4csjBgIUWySXuBOkXw7AwNuGU2
bo8dUoiSCeTpsR7+cDDMXYpIWjDvWgyq6ze6hcKVCHl0yxmVtXGoq5JE/rYB0tGa
IiX2d99AnkqwqxkalhVn5PiCxTcrrZkTvEqYOYZWaHu8shfC5D9frx0ULzteQRjK
C8GnINzlYC8Dt9SedRqLOpzHc1zeTe3+97XBBIqYkHO2jaSJ1YoY6SPVZL6l6TBC
vG6fVMd8bPNZzy59mv8zmHkRR+PhT7opZoecFgF8qakIVNyaxUGI2sftyriLvrJZ
ioGtSAe3rSukThYJxY8T3Ml45rmwkMicvL7qYZcLhq3Wbs1J7MnMhIjsWCiHBdLu
1B6Xy8QTP5w2UTEvqhfDGeFVwPWagzoPEJFyzIoSbTD7v4HgSBdRXjvynwHj2HDD
YggEbLxlC1Uupkx+zlbY6hZn18JBfRWQ+tUwEegbtzuJj6DT5l2qtIzyD2Q/PDrM
Ito2hAeqgzn3x+E7lZ7zVYy29aFYGOnETRUjyBp3KqgTMVrEZBGLYurB+3vzNZa1
I1XpxA+rXumdndoUZAObLLsicsCvghNHs2nHdH0TxCcdkk2BWw+arGPkXgIc+6my
vBbfxr5P/AcXrOn7lzFCrdlBWFBvsC20FZpdJs37pm38V8vYvj+EiONoQJhp087b
RdP2xWNBMNwBkqWvTY7HkPDXtlbx2+I3PcFqBQjNcVBYq+hao94kNP/6qH36ZHk+
RHzONDExWBHRhq5AFKqATlHEKDn4OMtX/ga1dSidPkKSfLH0WtytQZZPWha9iedm
/spFinG/rQTAJ+8iH/dUmov88dSdmoDOUNMJb1/7X3JVkF2h+FItDi1uczN+WYt6
Ie/PPOWPXog8i38EDmPRKJrftfpN/fMUeGKoJNoEy4kX9hm6zYe8zQqtURld/E6p
2//waNLdyYT3SUmSpMPp9vmeamAaRuhP3GyCdBNZj8GV3Il1l64vkmlo6gS7Xc6r
X6RnjGCsz/TubGfPixU6zl9rDAtLJrUPk1iK5LvV1VZ3IVTTQB5bh+odb+exOnvk
KmnDAKzSnIwfRhRZBZbbV7n6W4r8bNXk7e84aMkGafKf7MyiaEHDJ7KTCBsFoONA
U8ZXpH3dMb052hE1X0I5yBDTN83NsCCzxrugqPGQiNohw2uRGIHxQa/nBRtBC1eL
+lNgvuQpLaFQ+ODW0BsBoSm7yFRSyEYo2rNcLRLrJVWM4pldREzc93oDWHYJ46Ts
z4waCB5ymRn48ejTey9x+b6OJ31dU/ErwBfHKIFFRIUlqAvYQp8//iA8U4ENYgm4
NEWaSDvq/LdyexwzWkAz6dFw3ErU8/iesnM/WGbhkgPIBK+ynifVS20od2ApTJ87
d4tegXZsL6Is94EWEVRCS2HoAiIh+Qh+UmZwcAz93mYXHnfMxEOfzyEjaTohmeOR
U60Uvh+kPYhguuc1kRyASJFgTrfXzzrNqeu2LgcPH+qgN5gUhPaSmrKTrPPnilTI
9mh3jK+olWi5LVA2E1MtLED1ynmlOyHp18fXVMzIR6KK8vM+YSc4Kte7/4eeSB8w
+JN5is0FGLN2khSmt0PltEHWLicdh49bSuVErZHCn4KV9avTdezPI/Ergtp/Wh/6
pDbqIL2XXg0wlGTP9CK/UOGVXb5G6b5xGM2qqXaGR955mU7Dr39d7gZEuMFWFT0a
p/FP29fZ2zXTLzYgmvuaJ6TbWR5/bDvxm+lFqoqpbt2E6pHrVVwL1U0hBDQffvBK
mXXhQYkqq8seVgzV1Nn2uOE2dcNBIqCYtWZQJp9NkTtUIMwlKACjVfcnmv21Tlfn
ONEEiJRAumLDkvbFwDvlrF2TzcliDHw4c+Wx9P6Y/d8+R9wY9oloGEholEjJNnwp
cGYt/+aEAiYdothWYhx+JzdUPt1EOIQPmS6mEl41WiRjm+ncdOcc4rDqgLQmGg7V
198Bst5Hg7d3pvDmHpQupvpiFzRN3W5oVvW4bTxV+XjcM/LG0iOxMyZAO059LJu0
SMZFPOY1eIPyiEq+s5fr2GSWXWOY51ZJGTY5fBs/N7QmikhzrLZp/tGzEVx2QzQJ
W+CR3iYBB4ucG9GAI6asIqLcC7M3k3TChLx4DG9iVsVynCFxlMTDFJ1e4bBpCKi9
Y6uUDuK17FnHLZmpFTdyaV+O+BMErBRSy1jMR9HpI2hYu9si6SO+V1qE3iY57KLq
kVuY2L6vWcepRSwOM71swEU663k5mtvaivmbeXmpcGrFBp6AHcVCWgDpxy89lVHD
73Zz68+QIxGOqFD/ZKQV12kQEbONvNLQd6ieLTPcCvUzTgiQxXNG6vPyGVXkIRoT
cFbnSyHkIbzcjVH28qezxVps3haUm/I8qGEKT/wV2sCuwRTORrvNJDq2gpjEyvT+
CiBU3PKUKV5PkgsH6kWU/WCGBHTUu3cS4443Yap/c0W/1ypUTO+5yV0HPmromxoL
W7lyKl8VK+T+dQp3P0FYnlYPAP6KGwO99c1Lr06eqPxjc7Pg2n+uI4xPsFNAaGwx
SKZbtUGmneLrXTIj34VnVlzeznb978QG4iZyFhWV9UaStSv69j1RGIEKpqp3YP+m
vhrTkWAFjhUhqaScXoWaiaRJh+ZTinnIygTCocMJ5zWvJeqmSqE0b7yYBapXRNTP
0jWQStvLeGoUt0Mp7TP9Qj2ae+AH0G0ihY8lOANxMyMSqxu78F5VdJaK7bPQGSip
wFOGxVZtheAZ/fnmdokP4a0XJzeoN+kM5cyd0mVPXK2/ZQO/xe0gCtF7mMmy54Pa
ibNBb0Rn9OOyqlNYd5JDWTg1/u2imr8jSJIKcMJymvU230LTtrJ8enAakD54B7VZ
Es58ZplnXQQrNhlPrDNd6asoW8lrcdobQ5QJxKzIQYdqf7brWeTM/+ypD8qdUtU0
I6/Seqh8llPz5Y2F26WZc1Bg/Hn03vyto9QRKi5/J/cQ98hUd6FY/sTdoSwlLTYS
gUf6r2K8tu/ixT9Jp0gn+i4zc2oaBc93OTXQV5tbrhslX6ePmJCLvJwDmQwT+BdJ
ZSmPsBuborSTEkdrBLEaCtE05O78YPhI/HI7Rht3uwkxRyCrkrFb+EERfPSVV/1A
genJ80tLcWJCJDAufbLV5bn3NHm2N6Cagjc9OTi9dJf/ktdVQIOd330XnvSdmBnx
WBE75h4HkD1tomSo1cC83uChTsMwnLyuvFJVy2fVsx4ttd0w+Wwg9fQuBO963fjr
f758/pFSDZrOZKGI6SwtPS3mePvmF80QSjjJT6TWTSIloRrwAJyOBjAYkW5RTJn4
pXAIiEW9Stl53IgjxwvU/G+gZFgxqldXBMw9RfRLFqJXBewQnnYTtA3pL1FP8Inv
XAJQsAKvRYY/vn/uZZ1ghqPTZapI31ODZjW/EMjSGa9wtf7nwRee5NT1hd9d3Msn
h94T81lK7f+qkY8ZwoQHu31GciqdxgVnQ76fVgl90+JExZmz2sWUkNrXa87WoUnk
M2E5DjoLEXceAT1Lla5GLWLHRbgFLMh//rbeRAbQuEWTGniGKky4IeI73p8JqcCk
fg+iGeH5EFPkfa4UyQ2xpNUQVtz6w2nuvFaADc3l/ZRZFLedlwXg2G7LFr9ryL4z
+MxBpgSXk/dJ9Kc049P8EbmsDjOuJuklnqV+9tDXdYoJd9mKppBS6FbClScI9wKN
WujMoTwryyoLF6cUSdOwhWaEmuscUz9czV+Br4SBTYB9w27ccJWa2N1a5eIoG89l
Yoh1IkZ55OfzG+7jdI9YgxZdMxt4F7QI748S2nDvngi+cKMaP3iKW6nr3AjAyKlO
+U9n2+KJQIaCcIvask8f0TTN5oPa1b0bqOttCWVve4q/7j/LY+SFhkwJUVZYtAuk
hSoh+SD0FKevSEB1FFpa5q+nE66g7Btnu4YJsM4mKxLmUtoT1gcOfd7YLrJ04Thf
HGn/ojUb5Zpmu8KfouZDSIyzxcDHHsBef/xEN/r+JRiCOHXs7LjZCncNvXAjduv1
8AuyFIQWGPso8rLX9hdJvm7gSeEmx8caUR0EoDEAnh+2CdvuZNxpRam471Wz0CEo
NLNCXSG/ddfzhF7I9N00eaQ9gLF5DuhtlADWiQI9lyYfSey7xDyVDlr6xykZSNwN
1BwKIKI5XTekJyxhs1hCguX3JiDmFYS/8IN4j1LOgCmJjYEAfg+x44gxF08wes5L
Ge9gAc0LZxbzepBghap8zvujPaPPEhzdaMDtrdTvHa1FM0fSCtHFxyG7M9Uc6Dgw
eljToqffnk7oGUsNDlq3iNRqx5h2j33XHtcGWng9W8pOnOjvDrAz5EJN+OjNhFFl
bbgKCSbv3XwiMlIhrgrMK8iP/pnw2zOlkhmZ9ogmLWKunZirrlJYHSK4jGO1Cmhg
4NGtnFCAsXPwQfZpGinEYiBUFHarbfUc7Qe9oiWvoRpSfTM5T+DsgceJ1U4IRYaQ
4TDcEMmkQbumtIQKRcQEjuwsarx1H81ecGCSuQpO8Kfw5CGTbvtckYfMxBrXkj0N
J+T2liA8+rD8UyVrHpaGRkgVeYWvrA8qZS4jlLCkDe6jhTMNdcK9of7nUsP/1hlS
kGhQe5J9TTxIsKY4NAbVcRfw42/ACNYh3rWRVCDYFdpryuuac9DyHMLGYAz/2AIL
fCBMxE1R0ollmHjiORyQjbAWMGp5hOeM22hxxgLpUz4OYN6OzEDRwOFYq9bWFijq
6Oir1OY15d/8NMOPwiZUElXeshlKfn1RcZDucECXNieZJ8Mk3+1JFhzzCdBOUZ8o
eYFK2cCHum+m+uFVIOuSSpd/Ki2yETZlfzXbL14HajF4XGYwFZWN+9BCuNMvmtj1
JtAL/Vd65VNXPLVDTntxW7xMyhCgzDXp/VBtMQ8CY7Hu9aUoQPnhyHMZLeQ3gXi2
1J/QqYKUmpjqsgobfk5lK2tRcFjwOoW2MTp7fMd6rXNwIl7JtWXneGhIs/N87AKr
ghTKw7nDt0Jg8VS6JLqws3TVVtSxZjsrdVbyL3FEgKOSSmpT1oJMvw2FFbhU+LhC
lKZQzj/lqXD8nkTaIuH6RJbGjhJPnAb38lv1gzTnlq21fp9QxBsVnWR0T01nLzrc
KorwestRk5P9WBNKJjBwzPMrcfM1TG68osyvrkZMq5r5QtJTMPLlaOqPX1XrJq32
UQ9WUzVtbj/ndSoiAMppmYAd0KjUMNem0IC0MTefVLXOVLXqI29TZjSUu0aGLS+E
cx0UQ1h6eaN7sWEEKFNm9QUmL56OoCIR3PV96/KGcQFV1/TJiSqDF5qje0xj+VQJ
qQmbUO9O7NjwEeRpddoZGKKyU5/JIL7gPqd8hcMnNRllHVr2To6JSOEXosHOnyi3
Es1NukGakGEmt3xKVdSIPqlg5Ui0zyGgUAruljhAe2RTShjHC0DLBl58gTCBBYD5
7ob0gNab9QkKVcbM77p/Nde+5s3tztsgJRqJfNhgucj1kZezOnwMTUBP8zK7DY0R
iSLFFJN11wQZhGYnj6py3x8GkuVlT8kDEiLZdsMCDOlQLm2+Kmp+0Ae3NnoiaNZw
aZ00gRjei5npx9Y7Zs8XQx2X/abVF+l9cnDXi7pmtyjvhrCzlwKuvaC7cMNdHUqn
Uv6v6sSK4j/eEofWk8fV2ttSFCH2MU56G2Dx6RhkN+2ZlZDXulupVvFTTswoQUAy
U2d6hJ5ImXCzvPummV6jiR/Sf+4+6LswzgFMuq6n65wp9DXRL8SaUJMTqOxpZWJZ
u0vyaj6LXGzWYcQGNJiMC4b3AiBQtd7bcZI9YiP+0/NGjqNERtXYzcldGkybZb8m
ZIFuD/hJ1u1+JyEThlfxcKZMjKux7ENemIQCsP8HyOzBNEu9qTl6KuR73LynizZJ
HqSuZ4Z5TB/stnFGQsJEJEW8Yh8wC2KtLwgNtf9wvA+OK+EvzdPJaQo96ls6387V
mYOu7DHmACWOZOW1s47koYIBfRG+IYGYomcTPTZ15B/jvY0f3rGU1zkH+PCZRsBi
9ArCxRyydvanWuldVXEi2O1ieRSAxYKBGUhFp6Yv1tYlyFzwsVPJVN5N+fos7o/k
ypgIlJNnzbMVcr0j87Ej4jj3frPxNWPJml/BzkiBPGi+Br9HqxX64Jan60nck516
7kXjRqTlZ6VynMkHX5n4YQinxFub0hVsV8ZEmPEWepSvDdj7LsFOzayx/4MUrvRp
PC6e/NUweRPZFv6Kn3eW5j2adg6fiY0NneIWlwZa+HooN73FNWZGKj1wPnHljZ1E
v5EdNu38OoGx5mguw2ZQQlJmAex4qCG+3dkw7aPg4rpdXTI121YvenO9RyRioMuw
38XBQs3K/rnRA9heuuRpQDeaVdty871V99cyqNQWWl29HJVlT1ldXjQw8++WU9bF
HkAipozGwIaZJBaUENRFzu/Xb/VkX7mwbXL4GTBholz949NJR/vO/L4hCa48oNg9
9FdiacBJuDpo0pfMqQ29vfqjzCwKpw1HkU8op7S9PI3h4Dbvr/9/aaXq2P33ccoE
20PEXi1jeBz61JAOx5mvaB6s4VWPzOGsJtGo4yGMsrQIjA+RpK0S6CSV6RcqqSMO
rve2fitkAqZKl3TmJvmo3sQb8KGUkRtb9AhZlxq6a17NxPW3Hf5jg4e1vZj9m2r3
j9iLQ9621bWiP5e1BTeyft1oSSgHH0IjL+vEhNFNqFjDVp1DV7WbkB6VnqrQ+1XK
fwrP6UqamLq6afvnAFm1MoCo/3mYM4e++5IduThSeJ1FWZ4UotB6TWmKWPRAVd2C
rlj6Mwb1/oBrXVCCPeEmr/pZS7enAYD04Xy0SQ3mWnD8RPSrs6AoE6AuJPzYhpA1
Ho8Git/nwepUU9lzJPl8/nEHi7icB387ti/8n9jPfg7sPNqSBHJBG5KZoijyshc0
h7ZYJhf90qaoSOVh3skoK+jLjNYXywumKKqd61Rgd43dX+PH1ciWoDha/bYlm7I1
buTTCXcL0rtigxgcXwePIoOZ5KqXMNAqlgCUmBIY/wAuaFiGs8jRWpx8uo2eGjQv
583hnMjkql1DTD1uTIqyOQDsxul+x3TWlsGvmJ4Ig9sAxH4pu71w8KZEFT+Eg0Iv
5zN+a7yDXeA/+vQH4zmOi6FHS2J6Vm38sNtkN8V2Fs8Zs9tOlgKFsNhh4iQozS/m
bGAMnrJHeaqsjxNx0qmm0Ya5d8nHTsqQfsFDJZP76q+Vi8C/eZ3E7rtk0CMqAHOm
iHmefmer1r1z93bz8o5kxHU8Gftaj/L5O4sURfHK/MitECmZNtDbttPztlARmINN
/CMWlp26c41y7eyL3DukBLDkt0SNxum71rGtvk8RZg4h5xhhmL9HIJ/1pRdYVKK0
RWqdFzuZ5V2x7S6tJUxS2ueJia8J9hC+l8dA20MjRxmotrRkXLeUXP9nhW9Ak+Rr
5iswf9m2bskcKY06UAEHkmnD50pNwUkv4ZhbOBkgaU39OodSMluH1QqgqcFiFOXn
NLnWa5iSsEtenDeDs4qh2qE7Xg2C8dcAlNhRbJlMuPIDxCfJW7r+Vhj4Mmy7tMUC
G8daF+I/KaN9XPzjDf/3lgfbeRC8n20LvdjVL042nFPgAMt17q6aSHFaxCMnBvv9
OF2SsCe4LwkjPTtuA9qQXqUQbmAVVkh6OXlFlcGyw3eEep0f3tLXgEoLHSaMXocg
uRAOnzJMMKd1hvJCgsEvsKZzyFdRFu14tFJAhCMbFsIVffSXoNfIrrLc9r/HHoBq
ULnEPPbA/JvbBOpdcQ2J3zQKXsESY+dm8kgPdrLb3Oeh3RUFzLIMwkX7DmY8+WDL
zIzy+WOymlPQM8g8DSe2AXMcN0si3dSKRiHhhehb4ypWbRA0e45dV8hASFHOo/7e
miB/6YrwJr/QdZsrUcUvRSWWzjUU0+964wQmeRsdvl95W/WoXVjkqv420WfJfabQ
Ku5akwa+09V40u+Di/qraPspnBaFJCh2dwT/gKlxulu5MA/86uxzZl/jeLvRMTqk
zSeBTg/DvNh6xXIopfhYmmUWrgRKhANzRzCWqoYU1SX+6kAqNnRRwG+bTU4yEB57
2bHKmlxeRXcwh16UvCps5f3z8fGc7/ZQpmu9BtKpLuKF/I0S6s5/mLqZmdv0naKx
/o8PwV6z8qWp5pWDDC/RjPPFzPl2JGG4gZ4GJz0rq9jagYqNmRvgJTkdez3sTEwU
99yV7oZrbK/9hxG0DE+2G4qgcNnKSoXNB5wK2NwbYoPYgfSTdHZ43yaNVuOXk7uZ
gp0rZB2qu8UerbglSfWIBRhF2IkXbZuWBEhNzxraR6eg95d8rMem/DineV8Arz8M
FRZmYUeWEwObOJoEy9HelGNt12oOXX8H3F4R4gNuusYdBhC+XHxq2ZaRFhjCuQzA
v4O0leYZSML+jcThcynNA0JfczbVfV96xrwKBFEXqAUao7VWfuTR8S2lSqKw9EBb
VaXrvX7zf5Xx0ZCehiQOw45oU6DdkzJhjI4Y4Gh2Y8FOrJewD+ZMXVnTxipqGJ2d
Vvrg6K/AmFWosEcVoVwtwMS9RBH8cujJzUnTd3uF3OkC6gNkm3I9+RobuA3xoZuD
w8r/Pn1RfuZiYEWCminNydjLfwGl801whYpyYa7sEZKlPMSd5//C03hz9YUtda0u
f2ijLCu18YyoVkY8x6/Xw2RpJ2oviZ1KHxFjV7eTNE9GsImkUP5bqrA4QpERbx2J
P3m8FXXc72KzzoUMdNOn7O2jj3QI4g8AEbN9DuiCvTNG6s0gdD/cwdAHzgb87fDO
+7qeIHkUyTsV1l7ND5Inz0QBCK26cVdmvWYFSlIZUEhBtr//dkucwRB0oqDJd0tn
LyneACXai+NSMDwYaGT1ZYuDu3ny9mjyiEPeogc4Hj8pIfIYiOO0qVJHzC9+kxCr
y+IKwexI4HtsnTXBO2qiyV50xG9NW22qGfiezEwgeoU4RgdN5M8aMqL9HB9QeeZ8
qn8Jwx0ZO6hjANRPxH4KEASun1yKS1uMOyJ+ie2StYPaub0xkgMhjKwUZ8FQL9qq
9joiDYKd5rMrgFMqQIG0duVaEQKmAITG/PO6eRe5ljMxNj5THuG16ufpNqN07nIE
ZFEFOrhSuVEEJzdGb4RONnXJ0EBUHGn26x2kfA3XSj+GImdG+G9QUpAkquGDF2WT
1atH1GwvhqRfNv2xI2a+FNczpyESZ8WnOmBMkB4nV7AfK1As1OSqZMSII+gZkok0
SrzWmkooSRqywVw5A7wB+iV389BqMpqMPjZWeVCwaU0ExykzEdUMiwafEqGsAOKT
1TYvIUAyonjWEJEAV7KJii5EtRatEN/gEG/IvXkr0xPtoF9F91orYvFxJ8si48aI
bp6ZmGwLlxTESyvnWTJISuqdkFdI/khpGvMUGT0abfwgcFnMaCAkZ+NtrQ6u/mgx
L8BzxNMjmGkxX9uJhGV+nC1AGH6/21F1H+QlJ6h4B/PcGSWm5FJKNfHAHMD4cBw7
Ddkxa7bX833BlvcGjfjA/1vPSIZ614dtq5+1tVpdk6nQJBGdPaH+TLQqu9h3J83O
agaZJUIi5bhFqOpCamodGeipN7ZJbpLkzYoyvBGLxBp0T+qaybclcoSe4v0Lo0M4
HPppANNnah6A3amO81j6jmyDveCSebaWKh8FKqcylB92BMPkz0Vd5msNcO1wYpZ+
WEqTYrZX2vC8wxgK/kpuMTcJ3Q2rG76B54HFNiFr0siM0+uhiyjdOgw8vKwdcevf
mwNUIQxSpM14wz4BoPAfn+bZhsHXuCQo3MxavS2mdu00z35sUbnXNfCIGuQ44+rn
+0miAwcXohBaPoJI6DDoa30TGhE7KRhtcopwNlbg8Ip1VVF2lDI5KXAeeN27iGiD
yd6xBXh3QFsnhpcYgMB87oLkdfkv+9sIPVAyqYqEpgRFfirjNbjVgBEFbzvgvDhq
y+uSiFwKbiFRWB7kqYsW5qCNxQ6OcUlLe7X/IgTLqVn+cjkHDuFGgSMjtEwfOrzd
/iVWoV/fZa/bti+PF3evp/hV+INE+RoxJKgpe0JG7yC6vN7mKXVXbunVSlKWHisZ
1mkWbfrJ3YwpZ/6aBBaIPn/kwu1wTXaCeK1zRByq4LlRz2xtfHelvgnbbvc1Eypo
leL/eBK+wnB9/RjPkipjjJ/fRwluijsR802wffqgAZsuTORrYhCuBzSxEztT9Pm3
juZ2JywgxyAuuMPymk9MCm/XKPvYOV98dhpO39qpTFORuTtp6ILYBdzJL0yBDgfx
300pwINLVfAJci6863YBY7ZHX0vAgDiNQrMEf8DMMbuRHQ4uC4Q2Z1bxtoUl2ba1
Fw+knnhOWHQYEyBGidH8Yc1zM6CYEPX1hmpDrygiVzhIgyUV8XKlUCeceWH6s2Jk
NJ5Z+IsJXspPP+fl9ABwDOjTk6s2egCjMntJDgnv0xYgK2EyzBEmZEJ1KLNfZvDy
cnY+hXaudd0T2qjMrYDD2Dp+4ROLX7btJ1CGrb/q1UGpI39eqVmtG2rYb1eNjqX2
udqrd14be9Un20SK5HnkccmW/b+q79JJKyMHhNnwvq61Bjp830qHlTWEa/zSMpA6
hcV0elXC+QUs7ZasFmdR4u+3bWpuDAeh7pCAzFkP+V1ckWHNDOYy9b1GzwzQSLHL
7A1mYAukY5iMUodfldXvAEdFYAKx7lCxIXa0XmlNPVgpb9kGgjIJH71roDgELZbk
44TYdRqYMU4oMEVmQXVerH9qVozHWufCRXZkPgIOKoeHug43+KRuyXXj1iPRSeGs
66tqsa6F5erKLIg+ZH66/9zmfoHs4hM29xgeym34y3ijmaNuIulKriTfoJN2vOdA
tOyp2zgIr71ldiJtL6td63WyyWh3dxi4Vj8b/HvYohRKLY6yA49k4BC8qNTAaa0u
cOKPoWhB3blQ/u4KfEOuaZXsUsDyFX9qFD66Q1u7ZeHKMVgU+ZoZmyZAHHSSYtSK
HMe45YdMS11AvOo1BOQ7pJczhif2RKRVul7gdf4FsG0LMEm06xNoJbAPoQ3tGvM4
3G9/ZrL0AUWjVn9ecSMSYTq/QWkS/eDmGA8Ux3BHrm/0waK3ncPWYF30BxyU7zqE
LbF4My4THip57LQt+CKCo+0fB+SDLA5iv8EOhgRHGNqn+HLVQPMi3XD9FKRNMEoM
B0CMV9vBUw79jxFaI594f5lZc0cl6+VtpJBMU0WOM0iMMVw7jZCvnEOKZPhuhy2L
GaxIimB7Y93VMHIxJ+X2L6lqHsGjUtSMxlFuNWD4a1gvYxZvG1w9Ms7nG3nxR4Su
BKdLpSR0QOfWWzUHrb+wX/Xabovr7zyWEWtfoU8EEv/RrahoRUDjPOdop/Jjyv3w
Mtpe+tfAF83p6Cic7AcwUqaHIvR0TPSyZqY52WemYRUZK3p9dY1jDHBsBaCoH/95
q6zPUVKHptZcrv/eiybv5hXCWkIdpZCY2vDPj1ovMcpaEIq7mEA3HQty8vaI603r
MvfXI5dFcZ7rv7fhmRNpvZV5yYJPzyt4LTj77wlPyM9p5azN738OyA1TuAQIAwmf
hc7LKkQma27It5jzIyEpjloq35avhEQPRrRQggR6W9Bcm/ZMSCPjxeteT1Fyq1RA
AXSg10cCrbnA8BoL+itfYl/wu9c+/r1zwIy62leCzrfZvGyzNxfCX1UMWkt1oqEF
oAZMgCDfARxu6ChqAo3vPCE1LDsqJpuu7KxC0rnyaoBVskZkOwuraWJ4sKTA0f/H
0/21h7Bnz/x4EoDYIAN0UxgWN5AM//dQSHQPJBzIa64zd26cSc3klzJoJZ4dHbnb
cN8DCqWZtmNLxDUuQX6V/Ao9SNdqJ6c4bJXlzaIEidFsikwaPSIL0b8V7WA+/axg
uHD+onL3O8ZvzmfNDXl/jwp5kGFj+yfNJNVoBFFYiw8ABO8iM7siG0XY3MGwEPiP
GMCuplQ+1paHuitNve+76QwIxhAU1hsuREM34n+zimOfWHMiqVIQcXkpeLZUHF8x
SfNtcbKLqJTUCgCHJH8HMe1j6wE+jpTA0J48Mr8jXqcBFk+FLKehIdW/efMaiwYx
N9uofjdngymuwR2KnGL8EoM7Cm+JX207JAXDYXN0Ze5wmZ6ta73ij97pxPRttJMV
7fnCkBMslYqBbul7wEfqCLCMkQCFjwhFXl662AvjZphHhueb7r5n9Xy0j1fNgHyx
qBTZywdEeU0jupdmjEd7R4HTaiyt7cqy++nZ+tjcudXq+s18osiHhL2osPcN/Wd8
MWLmBdUSDchUVhJ4fdnOO6cKKraFJHH53BBDTpdSTSHxE9d2U89NhYHEmrpRNiJZ
JZ7tB7xxhVQXEh9wqN8u/Fvv0D9/OYIQy5Vr6M3hKdS1QxOZGNxOkOnU5j/8FAe2
KV5wMPxD7FNtyx+QFknzslIwjc8c01xR/b82EOB+kZ01+7vJyWdKgRPzBbA0J4Km
dQgVJ+YFvghj1NtW1u0JZRJUbncJx08uassTL2EAfuz34Z1Jf+UpzM60dADP/4pw
MImnySw2Ss+Hg8W6AhALvjZG0aGwCY1tPsSjKy39f6NtQ4AeFErONdRcQstMXFOi
S9Yf8JgUQxqXr2gCmlrjZnvqHUzbo4lqNiYBmBFvMsJrWKVTAeomsK+LYLGjQVvs
/1dP65xngJri4D5ryfjXW9VZZPXOmiIwtSV6QJ3qcU1UmypLPd9oSQc+ubnX001/
YsyA+513qLw1uqXNmaYAQNppu2HudnL21+sO/69ESOCAwNEVoxCR9FYb+izhFqGs
UAfRprz3F0YOKpoMkgJs+hMCNbF5vhTuPETnBJ7heDENQIN4DAhphYtvk+lxKyy+
1JqAY6Q40tzCsz1T5KW48cUTr4tNYRNiUzohENe2xoULYWwyawvcUiuTyWNVoCbA
iO+nzFAgSM1KM6igJtephgQzw14w1bLyPd355ctOdxzEjhKk70dZR94LXdtq6SHC
02Ar/HNUXtvFLV/E3kogjEh5oXZ5rC650Z5nNIg4gr8OVlxN3gYdbmbT7KL+hu3b
3hcTqt+g3He41/lDFZNTsyLqjrbx6I6qof5hD/yktcnixmPJ8zZ8aqLQce27gPMj
ZqFQCu61f6my+v1U7olZ4KZUHuH7+3mTrX9aMXhokz1n8wSMryxD0EDvJgkDEFWj
4zhOC0v+wQce7oa8AyedKy+R8NqreEa+PybMI1vuzHVsXqw4XldtSwZqsg7L+jHc
Pz7Tqj5Xg52RwTCwnHhANNnF9P5uNjWsf7/Uq8xfc0CBOLhNQv5Ie8qizQ1r8QxS
iTC03hKOi5MKJAD7vOSvA2bVoOCQhnOy4c8ZepPNqUtgTkKsocfwmA1wM0IcgeWR
xf986cy0aXq8IPki9axKJWHds1eCf53QAIJW7VrvHgL1NKIjquJCES2Zxn9bj7nI
3bpvNHTKTbxfByUwj3p+cydIiB3UCjLjMYA3B7z+ykZ8rfN4PS/yMHDOn6GcLXUd
fzN/w1ol23eNkNYIe81VEQjnjimbUu3whTOlIOy4l9zIF/iUUrjW8k4eqUBcfOwY
KyeTGsMcBVn+SyzCicqN1M9Vrc1VMSlkLP5TUL6CaeibvqGbxOgECZhXauXO/so0
71WperFIy7BwCA/BWWantgI1xhzof6yznoVvwZ8oxFS6VXqjJitoazayiLIv6/rc
gNxkyAN0Q/UMUXmxnQPzq8ED/6Pu5PPbip/ikCfaArm7mr4Avfk2y7fUTqS8aAie
jPIhlPWTME3cUpZFcPK0SYjLKdEj8Ew1fs6QiDJGdAX/C6UEYOXCUY9DE/B3MKj4
i3wxaYtj+7EOB7E0IStu9O/YWa41sWdlCfUoRub7ToxiWS1ATTpjFOT0KkB08ROy
X4mHqWmxjLurpPCn6R9dUG6L4DcXq9DOz4FncRSVVXb4KGyNgmJd+eGl5sOHUqfo
FPtK50hQf47K2oR9RExsn2a0bSwQQEAvvIfaOuSJL6uhYnZ1SWj9pD5ZpfAsaUaN
Gw/mBqQfWl+mN97sSlunxCReKMpOd/U6MBwwL64YPrvUU6AcznFrIXa249LPHDqo
YnlMtLZq3Iac3otSZTbyKXUac5byuEr0wGvDaTj/N0Y5kc19KtLh+1MBxPK47ASp
vIIy0MOkRpwUXxZ2gj8v0VXr14FxixE2P64BEgsx4XYuDJfdjU6SJVti/cCPig9F
ELVs/PVEs+w2aaHOh67nYJgiQTcuOFa30JIxom8eNNBjY0PDoA69Jix1MY46XCX3
W3jMMUywIhpvTYfYjbCJ6YGShU/PRCgCQeH6u7cDxSDL5Qjx+0wlNwgzgJRnDv5E
PD2XDN6T4SvspBN2TDrcKrQ8+qpSREHxY1+9a/w6sBB0iceixhtw1QHgCmk6tFNV
VgtpysLo93oCXcjKmBVOj5c+KVqwStG+pEhPNn+UCU87iajIOvUmflrXi6HXYUEt
fmC689V/NedJzBZ8jeQMDnhXKTM27fl7KwsuF7yEs/dVlBIcPp0z1qLMyfrIyDuM
2UlKlebnoHxa7HDW+yP89HGALtHyY0seSl/DBmaqOwah2pf4d/Xtu21BGcNv4cVU
Qq+2syBe1pclnvMHbPBxn1OrYiBKCa3X+K+Bg+z/RAq7VVpk9i34/sHf/8u+WBJf
G0fxmjQlxTyTNHhxJ57cHr1l//SCyM4o0QTNbGMZxz4P5AAfZLcilaHnKQw6ChQ3
EG+aMSikZouNhhJxuFsHOEIWuwJl5CcQeYu2DSburqB6YTh46ob+fvuzvQGNAZ6C
7bIT7py0kON8BQEATVulpNNp79XN3162zinXxC4zGiJMJS8gUyeiBNxfZW7cs2rr
nKMo3bz1D7VFZQzDGwnCwI/O/CQm17xQurTJErGuZ+IjKdoaCEMRaRKWUFAItPlp
GJDa2D54KRQmugMSYS1W+qP5BRY9uFf+auOpQOegX6oMRWw7gblerW794dhzWSTg
kLTxzmI9hhTxPj0yEtEH+lo7VTTi59Zeg629ko3pP5BvMoMi/TfSh8G8sojS4JrL
2xIQDRGgRKMNr/piS60LToTrDhs/AJcBmU9kjT+/MkuYGTrCDhlIDhWFB8CxC5c7
MmcWw1+XPbnyCmAyGfC7NdtopOpsN2KQyQHHUNx7RCR5IUYRsRwEjfR0i2NS+dvS
nDjQ8f9QsyE+RY4c/X2y8XbpUw9o7tJXkLg5H8LXn2EdpmyQfUAaXA7wEG2Piwai
fh4nSLrr8rAp6cBF2tLhfFcU+exi2fs6bRb5difxwIb/1r/zE3GtnFjxB+udQTaF
yjHPQp6oOOt4wWFmZzE9VSgrcznD6HNlQbSQVurbG4T4BPAG73Dk1YkJ/w8WuqiT
bci1k+WBFt4xFpyUsJnhu2q1LALHa0NeclxETMwvRGXqxh9GW9zdFKK9TqCr6PYx
eRg9GT3c2Ek3QuJdS6RUHP6ThnFWmoDX7e6jBm9Svncs6aslC8jRxFDhvlv23w5u
8GakKBLUhTUPJZFzSADhpHUof69yhvvpGs8vljZ12l/dQ1KzVGyv60Req6C+93It
f6AzUV90XtdWm99/dO7BGweHTB1+bSPoPaAm1d25lCGqq4vEZr7b+TvYOIb3/VPg
BAR4Lg0i1axheqQpy4F6QmtPNDzFtWJ6cX2iwhR4Vd6ELSpKTQ7AZ+8ytLo+4if8
ynsIhdivBZY1JthNgkzJpFJPeqDVZABfSJnyVKcJspaUUfToeV343Pre3lnCeKQ/
ZSCNzhqzdLPIQPJ7JBvcGzNTkE5o003U5sWxMo/0HHqP/cygJXJzdhAmj1uKdNmM
J0NT3B6QrW7v/+7BGkTmwZr3onNU5EPWfc+dyA0Dxrxzj3Xc99w2ThKmoElS+sfJ
9i38p38+IVCSLWBSgiM6e1a6YMHBJOQpGzCmfoZutCaj7AYaHFSKPunzL8/G77fQ
YnCbZpJ8/1knFyiPZa0dxbLKvs5kuSwTataUjdXTRHXgbKpGi27JqudPyIVs6zgs
rzen2nkWYhTrIgKHHs9E48+AP5Ou52BrcVIhumtqqygW3zeCAfkxIacZqgf6pCJG
N0FfPXrpo65UqXqlJgdJpUbdzoaYeQHeI0cmNfpCFSqwHbsKn+E/KbeCzhZCgU9w
7s0dgpHqjd3koQimDoSV3jMIC+E6J8lrKTGXcYkv11jNE5vj3HNmIMlcY838uWYq
HtLPP0lX+sCbB4KbJxCUi1G0Ur1hFhpaMRNLWr4M9TTvTT5VKTSOv7kiqW5H2Qyj
duwjrsUCvB6SL0cTE+5oRkbZgr0TZGa8chuafmUTDJEPmXH5YrmOMfZApWgoFmuI
eCI6XV7OCR5k1c05BUG3cDuoJoMeEPCCr/47r+GyRtnrhF5fUble9GDb8i8QO8UB
9ScGQ3YOZty+5/rWYp6ZHP2RF7TYzPbOaKI6fgSwJRhss/6A9z//vQgubngf7FeP
fnH0WvEFQBoGJYu2sSckgIK3Ao4A4Mnu/5kWwBkVhpHOdCHtdtdYbCzz6OIxHTzX
98lkBvF3oZXWBQf4Onh19/QtWSwSrSpjPyluJ+lY4dmQVU1Iod7OPC2JOgfJ8nMS
pvb9c6iWGITvVGdkO67XOJI44czQ+nEelXq/qVBOXCqYhM8UnFY0pgJ8TzXkGytV
gf/ZzI1lcDasvkjKNzp92eDueeJuqk+eoOcnzitLgOymHr5KUSy6G2luQ5i8Ro2R
zJHwJfYiWVOSseL7OUxBnOQgCjSV+IxZx3CM0QYNFtgcJEL2xFdx2I6i0PQf5Sjb
yZ0yc7u63lGStn1wK0ZzTVzny5gI43oiPpPgrT5p1Ydr33UVoP0hCSjTiZVG/yJZ
hWRKRLsfmNNkFNBJUqrktb5eV/A6pIjPvUKumqBgYoClc6rc9mAPPWEbSg2VnYrY
1ah9vibVh4tzsuhlbifSswmBnPuAUZOfNO795BVI1WnEPTv48xwUDOOGwjcH8AU8
HBSLSwbEi3j1Ojo+bbIv4zUeXPL+jz3f9WsKRKIhNCbFLSsEYbn9m6zI+aE2W9xq
C2Y6hfdsFb93wGcv2NOR0NUpT1CsBL+Bly6iyzEILm3n2qhwsnJY6HibLRxX9Y2E
v0Utw7L6wnvyJkKX4IgcvgPAxEArdTQ0NPlR26CsZCGp/FvNf1ohwpBK9AcxGirK
mF1B+xQNjrOgjJdryLC4nJy1SppmIHaMTmz88LVuGhaoXTqkEk42rGwsZyx5Xcy0
4iV8/Z1LjEtNShlDznGAQMFdZIoD0tbCX7726ELU+Bzp/+EMzcax8OyTL6otcF6U
SpCAPr2kAYadP6gbV58SnYCF1W7bUlKlFId2rlKncYrXB0tmKIGm4z+AjSQLNwkR
EJ1pY5i4JJEkMh7OihsaTJOwctX0641OjFeLYHKQsMvO2Xbtz1aJRAai8Sh2KLNq
/GYI9q3GawyQnu4LpAD8OCeqwRJ/oQRd8AIzLQRAc87NP3eisc/XnqUVMropjyQq
XmOLRndFqpIuVu9+Nffb/MbZf6V7SKF4/2WaOFG+pyRVM+rGWkU56oTM9YaoQgL6
wk4WvL66lgwJ/SoeWmghiMMKBnuFwOKzYWODDZmPmNRzycHZ7eHP3zESzfQFDPuL
+FMqhK+xdvPaPyPah4WVR0+P3iQPdYpZyKjASYgM7ae+MPh26d7LlfthGpvO72uL
Lds28sDUywzIGC3Si73qNFhlqD4iVERaM96jmdFiehzIE4s0kNsN7/8OMELPHFiJ
dUQSIP/5OSAm2I/4OXPsqH4cttRx+H7NJKyhNpD/sNIK85fdycLPadTo5LhNLm/t
7X/mvVgCKNQ8GerSQqNpB+oEup2lqg5NVpvPP6c0O5KYdn8aLAz51rF8OP3SYcU1
d9220EIGNAegI5q+A1OwK1z+pRL/oG58dYmDcD3ITEG94dOkHgsNHdBNbrYoMTIs
SPV7f5yOVEDmlxMbEcj35Ce5dGP8mWETqJ8Uq5iekrXh2851La9K0VuwaZCK5taV
Lk/tERVJBVEcdtHUfhrUVBo4k9JQbHxYbIuez6h/NZYZresJqcw/daigm5urROnb
K/myARICwUWBpF5byuO5QNOkIQZuuAzhAobjqEh2f0foTlyWTJb3/X4D/7+a8K9R
igd5qjqiw6YpPEjg/U5MVGTpPPWAYQVmGAhWd0EDM6XjboeHf8wE9OMrYJJbM243
UINhjd2FcznV4I8bmSErEmSUrem1SKDL4CZZDUBp8LMRQT9WBM1k00eMZRiJCqb1
wk184oU4HA4pushSURuCiL0bKPiO78NRykVG8cC5o/QoRhbKCsfTXcr63/my12FY
UBPYFUeiVz9Wv/fp8OQOodF/MP9J6vOPABmS1vn5L0EXXpVeeujr8L08/Wsd9V5s
Unn5ifjWWZfuwxsXyBVNpUO1RJ084VO/BpPVhdbkTLO2FbkQM8F58Eyr1OYkpnn0
nWvZVHc6HuEY7vjPlohGj4aiZvibHbbes+mKVLnTe3UhGi6KpRSjnHFoDR5SQgay
MflYMX3AkUdz+SPAvpcudyRc4reSG9OiOaExK1dnv0g49acbbof0+3y4AVosMOua
1ukwYt8RIv1wcrm+EC7E2wK7k/kltZb2h1I5Gnycebg//dW4Am2Q0dJrqxi8rf2B
mSO8Nnztjz1b7NLTEQze4M1OoBJWcofDaGr0y9h4kGvL2MRABzlFBQeE3Ocjk1x9
tu90T1AoeMtvG8e1nU1LgSvjMI52ETc1aRKMaaMpaaQwEeFOmrReylR2tNdaOYSn
fb07AIZKc9BMYBrbDHzQWXfn41c21WyQDkzNUgAug22nHCsUdQNSpwIS04l+T6rP
QmQT4XajMH3hnEwGeKOkWK9HKUJ6WM18jXE3/TlWHvXc9SAIRWQ0woqzmdkw+9aV
sjOdYMBJx+BpYhuAYtCWBBpaYsGgjphUCZXCQ98OowpBPdebMHHWGUYleZUwTmDs
Fx2rcBC8grm1hHU7FKGhBMDR/cFqjGiMHkGEsp6lIOxMeGoZSJa6ZKb7AcPNZF3H
8n9mKO+wym0Z/JiVeAZAwST7ZhUR5QcaHe/q4P2W9ZM3z8/NfbLQ5WLvY10wxkDh
tUIkzWB/nUXazRVwkLDizgLB8BJwNZk11OreTN9bkODrjCVGwtXhrjb9qdZYnQcg
gorDDGyMdYjOLDjm+IohyTIMak3jAra3wVoLJBEqA0bHqTq07uxDwVygdU7UBmtP
NOyOfbuto+jz2KD+syYKEgPZ3PdvWvMhK9fcmvAU2E5fp5I6HjjB7gKA0RO77s6i
5BIEd/2qvzC3c/cVLYOdNPumetqkHy4ieOKzZWfDwmNNIFIrb7+RFFkCrjlRTlvm
/52KfJM0IB1fdcLWRIDuPuyWYlPF1FNrxCm8oKxJXElnj1UiO5QQq8qkWq3UI5jd
UPf3w02MrB0RXjdYjArozm5GnZTIGtpWNp0VBNAUunnNcgWTsuyBCHEBHjc7cVsx
gezamt55hCogmqOH/eXVnGdSURnT1rxvoJUaaWIhufck2nD2v7QNZxyGO93y/kiQ
Hvn+wjNdyAfSQbHAKUaY8gI8c90GfHBkJKeFAm1+29edRRPVtJfd+8ULe5daMyM3
8w6lTRyJ1ZveeJeoOT3Gym8gZiSCxZNasH8F1ljiwUf0GNqplZlj6HSvxju6W60s
zFQ2VWbWtFRqTpBHCAbOILmUSpsZmA37+QOlt+iVfXHEge9pDkEEwNGYkWSLyCCb
B9ZvxQtNXtaSLBJTzPZC/6RCOwCdvqIJVG7ZtZnI1F+pprU2MSRBYBRGD/3S6fF5
D3h3i8QN8LKK+dwLk8tH4lN74tmOtr2HjssbqGhEzt/XI0o4/x3iIeKZS84kMsB+
bCAVUiCzWEO5jZ5PXoVsQQ+BFyEhdszQy1Jr8Tg/CwYVIVtZD/vfJ4Xc/rZLV9Kp
rkvSlFwS0p665Cg/BeOMCmAcF2mKjTiIsdRgKZC1FhsVUIsDVgnXWTS1Q8AxwPXh
S+g18PKRx5/jRz7c4urcO17tZkm5BuD6d37iTMWy8GiP/rCNzMUzblasEmsCtMbv
9Mon1LuSCFe7KBVlH3BzYJ5NGicn0g7SYb1csEK/yQDJgdze59GC6Xcg7j4Eq86o
N6dNdUnxR81MOR0C6lOnYaTTh95EXsLISKidid1LqAgMXRPZRIFWXhCGjN4AaH1u
yJU5J6W0f9/jw90Gzbv0Gk845BuN0hj2Y7QcTiRMF6W7vf30Tjn+sYTnAKwusi9e
gYFcI8qEkIhAKHi4UL6QIrGDcnNRGKjBzDPYJhGxkPQ9BBL+0pgbHREYMokRVVot
GjkuUxdEWME8CU7q0gjZjtbvA+QN9vMZxCfePpi6BIaMXX0XBH2VnBm/uLts8rFs
QUuMM01D/jri00hbsyNhUVevHdExA/IwK6QTEj40lZ+BeMPRZ2OEOUfkPIlv5yKc
1QDO/cbn0zHq9Yrbwu3K46Pyh6ac3j4w5/nbeYUORiYSGWQfoONoFhq3WWjtavnU
MbvYM/zaH8mpQIpPA97QWOIiXRtPTjoCdIOTwvbTm+WJU+869pEgA1ALj7dtOh6g
s6m6dDW1MAOR72wobONInWR8Wps0jA8m+nB/tzh4HhiX1sB/TjPu2mM/eSqTmUu1
NPL+/PcOTBKuFGgrPiBX6FcvvOnTswFmyxVUp1ybJgJaBUcLME/CQ2MZSgK1dktx
wToWzMZfcQjZI87W6LjJobFujEFlE2ekXvppPsjI0m95NFwF3gLI9+2OgQGBYnyj
rbgPFdlPWU3sG1fRpNO9QZ2ZXvPo6zRQX6gwS/iJscFSyZTPjKj5d2chKkYeSHVd
IiNRbRwdZMsfz8J9D0DlAd04m3AoDxq/7HpgGfdlMJiLcBmebNbPMuEuKs5vlaIF
mNJD26pRVdXbNjHFTmgXIoxKN0qDERLlTOS5uvQfH9HkJFhwVVi3P3hSMcd6Qitm
dTo6hKJOFdmchM8jxD5kszxbwGlw33LliGK2RbNfKNv+NJIg+O5q5EIXwSCBAhj7
zwxo09Sb56+hRoJzRF9X9+wcRqSWOrzO2Qhq7DubqUt1pco0Q1TcmOEpqhgm2DKv
Ml17u07r3ER1AkehTphoJLxXJQF8Ht7yBg1lQw3fi2l8Udt1y0i0imU+lnVwuU2+
kKx87xwE22cbcyGu2gegt060oIWB5VLkc6NJB5aN7u5+hzwchzID/e61vZnZfSdF
aHBKacd+LtBrKY5vKDdP0FIxuS+74SVzFrBGD2JuJHntx83I4J1vT48HH0u3RYrr
ljuwj6A4SDH7TFLObKfdbub4Gzhx7kmxh2C6ggnRZfUXSZ5cL18ojLjXIUZzrPyT
T/VqSXRzrKEwPm47IjV+xEbxsVDmiEbYuWEY6rxW3dB3qjYBqk1TFcyTIzeayf5Z
JKLoJPKRLC8flby9apl8ZQdQ9KXm1Qs/1T+8tzMMcFEs/llPZfxYpO8pHVe6jL0X
8oHluEisVIA1kwvVcS+M34zEAYSDN4p6aUCSK27WUipyqjO8M54ozKekxQtBtoxo
59RMEWUcUUKVP6Hv2FWDlOQxh7D5FN1yhwPJYqRUb+bAOOAyvtFcGDt+DzLO5GVD
pxlfeB9xXDXvjMw+JbKK1FJKZh+3EHoe83/xzioH8+po3AY5pUW69qG7Ie22D5v1
ThQFjWJsgNYHk04qkHRrcvQR/4/AZhgWnJp2SJ+hUZubiGbHzRTZttmpplgLR1tE
XCENZOcRS7Q6BePowOF9RVov/m7PTF8Bo8JB1IZudxvCYmoxJLY6JDNUOf2tG0Qe
2GuEr8ZmzSbx13iyMLC40RVsXe9Wwt6EsbH7e8lN9+S5jWQICYjioQrEw2GalmcB
8l6CrkpQr8D4ON+1twkQuXdIgI+RpRgNIBkMuY+MftUJj4S/TsuRnT9vKA2TOIjd
ICPW31hgvHo4LMuqSEn/uatxWhDwkus1cA9gSAael8QbEqNGgPwMr8B54D/e9I9e
MgbpFHMu8mJ8gMqvFNLt+schV0MKMnRyGEjHdmMLKLmdUqCOVdpVRkgKiEzgnz2K
6EdEoJ8IPG0FSFNVNHsCQP+FPCss1d1u5SFfseZyEF8t9PWR5wq/roV4UIibbeRv
kaJe5X1LoqosrAzB6opCYWVlMJqKCI+h4QHVWuqbh2qMuA0cKeq4uO7m5nNozElG
SpdpF8DwMi/R2np10ajEL2+o4dRiCLE5diT7kYS0jQ0BQMo5jS8xq28fypwK9wgv
xHbo7oAl4wv/6aIppWwodq0/bQTM9aSw2f5bs1oFsnAm0GbUnlW7+wQYbU0DumjH
c/xJZTJ7ZhL5kdd35IAso3CSjEHJ1VziE/h5Icyc/0Pe/7tBYwfLM3kxLU3nTF/6
mhnH8acs0s9oeeKzN3pOKxrFOb2xO1LxIb3ap4YMuFOaqOK9O/sIYG4so3PTPtQE
Tus6KByKE2JAb0332Mv0gsQa6pqx8hvCmmb3EvLwBqZlFfHx6hropErR/3MoA9hb
GutHirTepvN6HN779EIOf+p0mPH5Znjctzl/ZYg5f+ZXBIXZvdJQQ+AnxTxczvbE
oDbBP40PQEpGMx95r2sTpPjjgiL2LWVUizuFivWM3qKQ/5JJQy6y/n+HjbNVgU3G
uZt4GlggPRZCaqDwe/VlUkNayBzkNUiprwmfwHW4kDnlfIQFAJkRnq+c0Lm606Sj
xHm3MLlLIBXXRvJ1VoNlED+bRpG+x1gTVzsvcUxtTUvunzaRf5Bm+101jDCAX4uM
8ynLCtUG9Bt2wCpHiVIJJFVWRcJt8wQDIkkH9GsRz27O6hqE+TDi7b5CGwmLNWL1
0VH/8C3YD3ENTX8po63CTDvEgGW4vK0NhTCkiE9QwN/OaEijbEzYb5inl2gi1tzc
C78RjP+eEkSUveQokx3DhEPIxeIaP1KGZ/WinUBVRAMnx8U7owntAfsdVx/jfp8P
2+PLjHWNLqnXjZSjWm2Ga16zf+lcFu4cLSCfju98IPH0LgR8+LSDAxSXUMPBDDux
vetYmzSzZldiMKqQjSRDkZ3EIXRepk7q8J0yP6pS/ZzkZQwM9IWBNDXvp46TGtFg
/xGl1+ih5HnD7P0Uh0KdDSAvswmitTBgh2wj9BgvPjdJzJ/UYMxecTatNErv0Shm
EIk89cDaxiqGvPtKXBuWxewBtujbHHlu5McWbVb5XSp8fFtI/SXY0iX18MqvKpOb
ZqCCA3EJ+4AFC2xg+inKBCPlER+TTxH98tKWvdfpFw8Q+O070s4tyqfVIIM2yfRs
aKh0yz5OpzFk0cbqyXTYa7vOfK1qQHf/F2zNacyCGU07Yhs/NcVQeDWy2qEOJzjP
KtlKgJMgLHNt34v0kEJ+lblDo9aBEup8ojnC3Ml+8A+nP8m6C0IiWnG6VtzxSqsi
pWcVfZWV9ktJLHykHBva9qRsc3PR/fzAgmNFldKT94n9r/XKe325PwFgaWsfVzKb
a4DjPrtrdKlzT92Ks2FKQ3ezLJX6XRKPllwucpai4jYT+GnDUmHu6DIyB6D3ZmDs
UEvfCwLYJ37SzqZ9rJCUGlqri/qb3DG4tmtLi4ocWpht0h7NHhdx7kkHBYeOAvbQ
/4vH2Gt7MvNgTUrhGtQGdPaaUOHLRAe0kvVTKYXREKXDBWx+CkkH45y80sNnOG+6
VFeTPAg0sSsQ8OsqCsYw3h0kpE9o4r9/XO0xz5EJzOV4Zh88z7HJKjJheW2T8hjT
YEYPVV2mWMGJzAbczUUJ8LpqEJgOGrynPiV7d77GeegM21HRe8lXmMRfWPAiYVHS
Mt3m4UgnVbt3tEfNgMrUaxsRgNK/SN5fbmbKwE9Q+MGGverbiecQ1x1BPj3ly82M
6sBgCqUAbBRNCOgj9YGwIpTOfp1OYoOGM1LfC9y6Pu7BmAvTvKNnWIxvVduvhGIW
gg/47t03wzqNSgNCGtZk5Y5r53pNdzoR1kZJE54+YcXnRm68J24JYwSmZOG8nggZ
dOmiSRWvny09JDjjjtSspFcEPRpe45QLoOfRheFyOTn9maHfSvuHzv0KTdOlm9uS
I5QZ7KLB3gkxyJKa8Y0ipLUjvJR3heUup9fa3d6LOFXfhZcwDeqXopN5/EyINjYE
S0mnFTgS3Wduq1Rob7cwOxKTYS0vVKc8Y/b09Qctt6b/94ucG9IhMVsKkwFb098y
yF3jKuTfFAepi6CMde+YOr0zjSaZwK9wupV9QKJtR3aNrw5F7/tkaeXAiOQWMDUf
yKqLXZE8//RFbiBUseOzKYsBPaM4buXi6jtsHW93qpgkLtb3G3/eb7mDJAWOwUOC
AjiU5+aUL8d4HjTM/hWAp1lGRKL/mCrwICF7AiWTRbYiM8N2xaxfOqKa/Mmm2bbN
bMB2tglHmDG0ewqCx/TtHEDpcWIG3sx20P79nHNDBe1BqiH+3MYu7aF6NZdksC3A
9bFxW3twnTBPU4WMFC7GQc8sY6J96Dsi2OwHPUypBuqp+aDskf9YKCmppCGYb+Yl
f/3gnxBN87c9368ajCJ9kuFZgyhDGkiRoXC+RTzZdkrqlzfsHyen8Gvll7wb1yg4
xATG2m3vRwKICKlw9EQBcBQSViX0g6WZSfShW6KKDdH3uM8fuBFz/31+yqNopTOb
2fb6x2JRTaZmrflFPcmNTaumZPdxKgX104Iw72a9L+kh2P92bIommq0UGhUZ9YYH
qie6m7uL2yEg36LsM7/MLFZCzoh7Xbakd9qGeU9biEyIsD0G8PlXr88yVzZpjE7A
56Y/DBbKXEq1eKYLYpC96bFOGGeztAzd17jxAl5VNfjG4mOJ6k2gY8y0xZXRnNsL
MAelgmi+dMKuLWWOtqkzLRLnUV2P6PAbQy7hCjhS/J8c/h7PMG0DfnvnnHdgNXsq
Mz8K0lHbwl6hZ4kplPI7NSnf2icSYWBAekik3S33uMaVBlkepxyPw8cCpJCljZ7u
rPMoJykvGECzdi4tB8K7a8jkeZ/Bsz4YhnpFmXSrlXS7rZljS4/X2oz8XZ9w8Le1
VnNnLNMh93YiuS5Bo07X3K3BzLUL7yPztIXb52kK7Iax7v/Lc0BGyuz+8s1pHQpD
nwGoc/2rsVR9ltqHwdd3BgnA6/YVinNmXDvWJaPGouj0XJSppzlMQvdRNQ3kfX+W
pAFVD9B34TtBIwg+RlpRAazX91GGW+4bXLH7WREjCLtG07z+TMhbvoIzfhNzua3j
+fORReNvdzar0VtZO0kgoC2BlQnCRToW+0z0NkOnd0rsh4J9KOv4SOFiHpp3Yu3L
sb79YOatHPuL8qG6fhPSNY0j8aGbwX0Y+O8a+WN2EvSCLIR8Kpp32Kx1eB52hodt
Txy37Fhp76LAmwPSWWvpZo3TubIBS5410j+/bqQK0blCQbdLjYm5CPNCelY8sg7X
QIkp6shdcWEY5uJHacqGBEWoDgLFEcWNGF1MHtRto6D9aBFpVR8VwGvAQ14OlQDz
tsS8jGKHmkoD5BHUX1gh7StFlKSW4aLDHd0wlNuUsTyVCTJjxX8qplxbqnLflpps
clZ2RegFbI3513noJ7d7G601MbPR/XzUyBNE0tYOILvcYDu1tF0xpn2B7ItyFPeH
lk+kEY4RhqQ/Fww74OHNzDp+0pakRNYVTlzOw2fpd21Kkcjc7p1zPKt3kuLsVrFf
ViJ9razgkZC5OhxQc/FpEiH+ZnXKE7/mrYa2GuiOt4tvk/Y56vu19/9JHqC5GN2y
QFuPEqVZSnFEOYlv6hUNQYupRQqL1RBKFPtQHfScrfiHUO52y+8VJrC/zk5a0UaT
CzJPo1G8Y5J7VbPthYpGmzRJ3GhjHpsHPCjkAQzmpfm+8AJMN7byUGHjo5TcI0zx
Ss5e/T3dh/8T4T27dBMVrk6bq3MWoAD91xuP0OiY223yO4QbEwCkZlG8t2oT8Ut/
2MQUmKWAzdHJTR+dG0p9vbb2qYeNDHEh3EXDUJ7dq5U5gfh9wAFd8kw1Q3eVXSC1
shLo/x4aYAoof5EJcqMniHjYDLMpSp0UrcOmVn0pWFJvwWFipMnboMlt1/wvl6RB
FerQEPQfW5wNwT9fzm/J6knOntn0nKmann7S5YplHtnmO+upPXWhzqaegemTX8xV
KP4D4CshmxRA8RCI3d38Hygy6vgmRBEz5U8jeh/9jhGSoATJWMIeXnOvkIvra2E3
k+XLNILVWOybTog3AedqRdhINQUVTxqxaWOAknH8ha70+yKNMt61W298BqsvdatG
xrLoS86pY5sy5ZQoNF/v4ZnsJhwIbxCH1qqsUqDylHMfZM6yc6AxxpY/sEwKTx/T
tjx5svMNhbP1hD1xxsMlcoPplKMjXpFO1qgmGoeh1/CcZxmXwy8saE0jc09LlkWl
NZLEe+uMBiceMKvkVQrQrbCDil+F89e2FnpwYdyHUaBMNIlPh+TsDvFDblur4qh6
U2wqXn7jS05lLUcDgxq5hpd+47aDN1jma0dFXk5G9nq4NZFaIlQqVXL1EoaEdJ1u
PaB0DFKEanyy3+QvLYkvQSGAeIOiU5MoiPO95mSFUtfGxcHpQsFQVxfAoNgZ8zEZ
g69bvaXQL7Hej8HC2bh9m9cSYF0tuVnxYQoykt3X1OZwtiZxThHyWfpxbYxD0Ed1
JVeQRnA6q3EIKkIvznTYse/gbidDhjGTFaxtuJcWHS9h2wbt9kVsZ1Y4P1pX2B9r
trvhTM4CHC6yNpAnP07p0E2PSsDIPTMKS9H0/jtU29ww1QGXkL32ptrX3p2loEra
abdUISyLRM20SaX7/N5P8vRxFhs7n7uL5xX0ilhfIOJhbBoTaRYsiMFVnKfZKDlT
G6FkI9o5cwp3ZyzFD0fdnytPbTm8jsN3ay+OcUuW/nLRJwdTka2wnyAfOmK4/9Yg
EhVNJNGrddWE0fuluG9bsBqWh0uun70Bor0m6NbuZ+s2QQxl61YNP6QO3GqINqjy
lLsaY8DWOt71Exls3QbCr/SF/+lqBlPcsEz3/3+YU05CT1BGtKFmaOa+o/1/rY/K
mndQw1emk9JarKfoIFsCgX+PRuZMtlQmiWSJV4sGWb7UIccsgfJVMioE+ng8mZTO
qgXMWZjuhDvLK77Ur4cunDn+u7UKVmcxV/OmqvB4FYmnD1OdUFh6Kj6j8z1Wn735
7vBlOa1Ec27xhvSobLN4mw6LgZKeUsRpfzT5B2S/m4SK4I3JYmCJKLpV1tSfrHI5
cDyqZg1/3STCkymLVBTVTcqm2ZrYV89aZrcwT1HEOiDB+UnMmRbh++wYRrHE2tLH
MqmlOOJnzp6It+W0nhl9rs405gNzHikMdkq1ucCbpgDRthfg/J/bSBMdjDvjeqAy
79eaKNTLpV9AkWWcT3T7U8JDaFcsvaaeCscsI9D7PDOxVFqBcO05fRvb+Ax97qtR
WONeJ/G7rwLPME9Yj3xSmcE7Q2lnJVHi73endZ6BhnMqbiS8sh2xbxbH5SvaXKxS
t1KfWSxrY4DTOr4iM88kXWfHAQc2o+oRHfn+S6XKU+Ntgm9t/S0tTPw3/t28SnP8
ohFWuGwqUOe7eRUBx3d9FFwWIcFGxMs6ZdfpySpLL6fnX6xzcCQNs6xj8YD9+yd5
XaCZd1WE2FYCbqcPMdohMtiHFk/vDIjkHAFSuPEkmhvXCz6y35/pBp8scJWziT4y
I9WGoOx9Sp1GY5OQU6ZATuweXboChnN8mPcpiy9s1PQg/50I2n/OTRdsfE6xV0pH
OZ/lMtbFOT0xTznCFaXlD9ElscfwquLv5kQO4+dNwYQZ+kVyMHWE8iPhRZZ7/tql
aQYXadk0UE46FNjmiQ8wfWyzAZG08GSO3FZ+EdpSglxM963+NyITIqbRBet5j0+0
q/NyDfv8//NN6U1zbA1aBHjvNQiodWpPfppWUlQuG6pAnN5qxKlLMheKvyK0Blyr
IDv2JnPB5yS1EW3yE545423DAXLy/rpoKupMnnGNMPDAamhX2sxmsRpHmPKJfSqb
C81KiyEsOaTeApRtxq54Oes6UobOqVTy9J+6Mpnj9UeruLYBdw2qNT0Za8HlC4nR
YMOgGQZ+CmJhhM43tjJgTtKD1vz6l823bc5QIO05JT2jMS/hZbH1DSMueGmSXgfI
Xr8P421j632p8HoE5lTZJ0IpjH13iS+ZRmYVwuQD+hNfo8MHhSIe58/F73CRUVcx
f3PhNc3SS1z8ZO3djd6hPuKY/R0y6EbmMxqzLGbYGRdwBVG0m+jgEBFuKlFwwi9/
bsZAzjSzh/LJ2tbgt2me8EnrO4qmE6/Z7ZwKX6iwVgIVfJwSxvkIIZ/wVdvUebzt
1O6de4ASSSVutkv12OmsAuy8meAxlcAcQvozd67TmWgdciI0sDYZamcYTSdaphEl
wONwbW6N/Uy2Xu7jP342Ws6X0rkycCNGxNWLfAJ4F89Mn3XE87uwf8YuHUqNzsKM
39uR9XYXbsECL28gPymvfoWC2yL0thAPddGY+vv56APr6CD3CkuzOTFH//iTSYyA
jsxmjtxBEqTg9hEa7LZR4vjvBTLy3l4jhLSUAqVIcq7LPLLx7Vfk6WJi9LQSCTBc
NvxFM1J1kfQvvfzuo857RjNwypauLfuoSgulPkx8piVExWz9HP2bbMhG/gAjv15Z
hag7beWzhoPWf9b0U4Cryn+tiXesdqGxEQViL7yS/npErL5FzIODKZuFPJIQ/2/v
TIsng6b/Jl9DJZWR55FmA+w1c6l+3XGMT2mgyYx/RCWRmyBueJSBWGWzTECpPfwd
GaDLtW0o1WiB/lkeh/KDopsPnmkvi8sJerbGSEejYeSxvCFaP3pI2aLoW4bdeSPd
NdKNvxI8Ob+VqDZW3nhGV4X58+Mnc4OK4F+ReMQIqkiCEi10T5ozKlQHXWBNYGkw
UYC5Hixw6GNoaHhNiv5ayQCJDqcR+H9vJRVAtjr/skm5oJ94Rr3uRohBurnbFKXn
ts6naZPlo+QGsUfw8RvcIaa9/JZPQaLEflBdm+cm8gJVyPmhrWjU6JFcSn7VtBXH
2lJbJTcDFu/8g1MaTf9+YyqjrdNODhpfIthLDhntR5b+O32dXwFSmu7BrKNlb0TQ
4dL0wtcL63GI4ZxaSfiltuRCY8FAUIB7pP3J6hLjdJrVWQiwjGYhYIBaeIQqnLjd
ztrpQzdnNuprfq0/tZHFzR5KD1HQaukkD96Qumv7LFgmoOknyVP2yx0yJXc846f4
gPQJp7E1xrM3q2/+JCZPtyCUXzNTyqbsAQhR5RGKPqYmfvC98+4MLp0qQeSDjU3Z
VtuBmHImX/HcG3Uvne+C0VsyXKRw2QLUMAqoSg29UIF9xqif1ge7lpQoij1Nd3v1
zj3C35txfmJqlv3QnuVheoaGX0qjyNjCg7bo1+8oC++DzHHJn5ZeqKezs6I3lTah
SCbIrN69uAKqaOv865gF8NoSAlBiH8RQf5cW2Gt9V837VMrymvuUTxLIjhW1SDu8
lida26rxuiZDgPBF6XLRBWb+cWvWm/NqsiqH1ekc5IChgAhE2MPmlctuPtoAy540
X2WdhAeuM+HTMFHNavAKra5X+isfX5HxJxVSUj8HBC/As6is2XaZr/KTU7FIfLan
JSXMhi9vozPB5PZJI/Kg3E29dC2bySW0FVa7id/eqAWFQLwbsUgmmpVjf8X4jWTa
qL59KPH9nDprFref8Liwd8gXaIRFSrnvi5xWrJC0bwuiFyf3wyZfY+TFJzJ5GItu
Ue6LUbTeXkAjt9aNz91hOZRGcdXqls+KFyqSQ8CiHVMaCloJYfx5nKISakFe4tlz
mBYxZgw8jwsF/x1ib67iAy5o+zCNP1O6wYzzbaQcsRXa45aCKl5CFDm+fojPsTwG
sM/Kf+67QDWsLRu2WlqE5nYLwWy3GffhHYI7eBAOWAbceFOt0b7xPg9Z/lKDpgpB
IGldCUdP7RVEbBgbp4Xi0I/G5JypENKkk19rNIQWeDxnY2qPZxurD4ubBVMxMTMA
Mhh8BlhIYRsTgLsEtuBY4DqMR1CYpHUL+VrML+yvYFGvEeRH8abI4t0eSJnmk1kJ
T/VtrGm4RDq+N/crL3RmwIARpJM1TRZpaUQ473sPZ1wFHeLmUZafe9DIDCz7UX/M
yBoP/EqZ4mdvQ2eohIrq1r+hQmItL4trw1eTSN0/fQ4KxH0zYC5PafALbEt9Q/rq
BEOaFH8tRHPUxd6XswA/QviwmdFF8ll3pUeXu68OpuN/1sznu0pg89U+Bpo/kJ7S
7L1hX6dbMQApb+/y0PsFrLp2tocZejRd6yaBCQDgf3QY+U6QFBQS36Ao2/9nilbm
rPEByFXwl319VaRi8A55es7P7aOhMDqqlmqteOk8FqWC7Xjs4VtxeYo4WKmh1Bxv
clS68qkxGkaVpOBvVLlLShXlyKKOGIzRRSPEYRuTCCu2sgceLniOD5uSToxe5t4a
bt24xQbJMIze/YGKX1rCHY9o/A4SUsMdOzyXGPUV9QS43KjJVyHW0wc/hLTuRRU/
RfvYgmCZ7F78FlsJNVaZy3pbi8mbJGVJUxLxl6n4dZEBUjsCBG8Nx0sh8ekYdg07
y1YzKDodWGPLh/FrHMOoJeFTZmD/9Kl4Gr5c/yUS/gU0ZVKAq5dDcKNDnRhTA7xc
tpdbliz2HIO4q4NOKP/fBhJc0KaEGuBF4vh3J3bbOcofXRaO8ShrGjIVfm1W4PqM
nL7LrtHtNXTniZRMyobTUzpXN8nYDNWYAi0W65AlHalhcgpxEorz/bfsEKuZ1aAQ
VgJqyRlFyruU/mH+eimjfmCVvcLMhzu5tcb+Km9kWkQkUGTt+nHghBeFLbZBSlA1
D20EQn9LjX08sCYzfYmUaZ3XyktlamGIC0FcbMv9HxE3ws8wmx2jZsbpOKm6xc3A
Lj10GFMFa4y4yu7AsjOT8mErEsE+I9779ZvHbAyZEaNHnux5oe25876sVOOGXhJO
cptZUrUa8SuPk4UZ+KmhI5xlIFwrNwh2x3z0xADvMBAPKKMd+XjCNB2gm1YIt3Uu
sCabTeFDbXQPQePM2mNA0hMZo8dZyArt65t993vJnJwc685XZeJzoHyKcUwwD500
z8kEBICrgRprCSeVYqdNmi3REV9ZVpXa21XVPPpUmDyRmYhoj8oxD1MtDkF+bdED
s+L0+oKntoS+TQXKVwyumuPIifnPXN5oaa8SmEP9oceVYs1n7215lNjMKO2mJOJ4
b0EOAzqJ+WSGwdWWP2PaV6d5hzzS6lLca04zorm7+82h6qnmroL+qf4h1rsw3akV
g2QSS+z5QIdG5F0nKwUYP3tdmObRrLxMTXRYxUoT/PBmXBhpbAFjQjdZKTm6glHz
kmKHOkr3liMR+7bGn65Y++1D6c3O11p4se7mbcupEpvfCNw20Feo4StVdUBhL3bm
fgDtQjtXBAHzfCefEX/5VMPtC2qswVQTsTI4K/RTYjbD1+NPUNoN3FeOfABi1004
QuHsK/Pc6h4HMX2y+q7xDxuX2DGbKQit9iHG/DraOvU+ZaC1HuO38NAd/P98z9Za
LE7diQ3nH9QtQtakKaTfu9NNB/yVUuFuaCYYcFuFOeGRXWau+QnNYdAg67FgXf2p
nosjK8bDtmM17Z5iWsel9JCucAAuoC9Gx9nf/Ib2G+BlisrXlsK1/wYw9YmNiAx5
FzBUC/8pBp0rK1jYv7vCh+U3Cq2ZYEmJAbvJeLvKKHysSweQ0Vjfh2jrAnknHlJd
5Q1Rllr8b61yIBI6paVxHJpWLdq3xc9gk6agffC7kVL6f6yOHKizYEjrrqCDv7y5
AvT21cU/W9Db+BnybcSZsEoWJKxGmZABNkFnsGXEhYj2STMDiAlbldMnTEw+9sUZ
jZNZeMRWhh7iYUIOlf4X4nPb7XJC+IBFBXaEsrUbVDdV5XaaonfNRzFT0DKdouW7
vG7ROPT2Hg+S1XAiKjNanM4T3AMmdeQWHNUCGpx5r5EV4oB8wemd7008XvFErH3+
qY4TCzcRMjvxWubWqUlTh0cY7x85uZ6giVlDt1eL1BcfhF/indbtAlYCN0n08+rd
4FMPibZIFSePM7DPS/WH9yEMntbmg02gP3iWrxaQEyj9TQmS/GuLnPYXzTUM05F8
AWuEoS+OoIsAWt2u5Wr2MQU//MpyZ719jvlsls+YK6Dqqq2gnKFgP5w71dDHIklh
VilUxIjlYHEEZ4fOWYpYK+5O73wL4JXnoxmfA7wG0YwcWduQ1ROD5zOpqywmAdZj
efEqcp2+Q/U+z0y/EauePKuleG//qxU0EPEPJTrFCVuDZ1+9BQZaeL048AVIj08+
kmMQ49ONyix5zMm1icQFFHuuQwzzd67BHxroimg3oUAOBLL6QHACX88UmfiaKcFR
kviXfn2dcXQLvO7WmAoLY43IV7pj4BeqgSw8qCpsslGBwqSckQYLwXg2UKruJ9wh
C63M3WZkn3Ku40evWfd8fto26D+UYkOhaXVi35Pt9gdbPVdNS/pfB1EgxhUUjwhd
NgCsUCkHUfkM2ceANLBsrCa6roMoh7S98yFxq5K/lZHk5WycchrFvNPjPXfoeyDI
H2opYenlBypiNfLxWhhPvr7WWgMRc3km9wE1zLiqqp60mGEe1Z5ot7o8Li8PF9k8
x14Co7bkyP7VXt4t2sUA7hZkwmv+3azuPhvEnSCjClRYW0wSrtnUOebcW00yt68T
CT7DbqoN1wxdzvFPbjXFvigt8F1mAPu5LGhMLGxmrx+OeIh9tIP4dwCfVvzArMQI
1xjFwnlHTQgC66RnfdA7OnHcwyk15FbgBKKoMZrfS5lldy3kenoKMkA9HeHDRCEL
rgJegzkkVMEaUlkggHOg1d9SbSJAX4+aHNTV0zFQx2Y+KfJtQNxYWfwm6eBEkloB
yipywaT5/fpDKCm9zUqWW858sfgcDfvGJH9+1ZS7QLxt2wRx/51JeT/RMdK0gtBa
iPulj6QsBHkoRW/lUZ41JGve4v6QQg1+Vi7mwINQgr/YUS+WNDoLnZw+t+6Q8nY1
ODHV57V3G58SPThLxEpWxxwxYyz+6xm7n+TX2kPUit81Koi4LGSZTrXlrbHtbrp8
pBUDOiX38U1sGZVld+spkg20d9mD1etv2DPBkSbaXyTs+OLTC35otT1MVcL9Brzj
iUY1w9ZvHD0bOJIBK7n6DY5ZxvpoeWnlikew23AJBFNTGEyQHy1ZCJI4RsUjqlQO
xSodyf1wnJqLhlACxvHO3oM7EU2e/LfU5W1/UPh2DG4ZGfM+xvunE7utVzjA5C4w
2LIJcXI4D7AS4IHdf5WV5qEodCupxUKkptpZOIxFZRMPtKOwL0zSadfYywkjhKdP
BN+pktVeMK1ZAL5rjibReFkPrdxqJhydwm1QylZWFzCjNsKrMNvHrXLTZg1LD3CG
P+OzZMl2CcAUwvre1TEzL6yEYA26GjFX6VrcUWXJDptpInPmf5CXyvJA06p1xTkn
avYtFJfnU85xjx31cIvxaHnwur6T89Q4l6n3hrgnOXIZLASW5ZixpxNQ/JNO1oiL
huC5tKmoGejb09Gu3A3GbDYlMgO1y/Qaj2WG+VYKsm7KCON5QPc3iPEH2wVLiHQR
LE0D3OLhm3HlV+DE8cq3jjW83KltcK8ZVTu9+/xp7REoA3s3Tiu7NztTOFL+2fFb
eh52Ow+aehSM7j3BsWTl7ylGL+dWhnHtwS3mqHJPpX1rI2OxK7lHemTWJVeAIrE4
SUzSrNfVDpza/cuS3nzPgYKvtR3TZFs57YHH2U0v6otjy+bEKDyAFwY+MVIQAX30
8Ab7SwF5b4LpKqIm3jhlXFSWwK/f7+tv0U8YyC5uYUA/54UoHZSxVVni4JZLstlV
LOEyUXrYXBKAJmL4cu8N6Q5yDJKE/QJO2/TwfmfLnyWPFepAww4vKyusCnJX0PH+
r2y7V7UJRj/o/mUUwJxCFYWQmAr7pr3Ra0k55CW8jaWjnh6YsHibH3zPffWLHmJu
ts1fPunhURhEGY+DEk2HVW+nseVZLp2jocGVTEdUdC1+MdXEBcNdV8+Q05v8omCU
RSJGxbyPkvAdyQBsuwJpToGmW4gmLQWWxFD2pC2LPna/0Ly73c+etyRFScBh1ZIk
xbY9/mnNwCvbc7/2dAprNHI0KY6wouHduBLuo+QtiO8dguF8j5UqM2VGT+hCbjF6
SNH6+SsWY4TUE2XugEsGP/byCyQgXynkspPDyBctUYoH5l5egEv5c5Fuudvvxw1w
/lq4WWsvWUJjVxE65EexKXjssNzXsGktlni/+GP2jQQrj50bYGc0UD9rYLsDENR9
nPya3t8dRsYSn4O5vimOJeWh8yL4n5Z8FxiQirSPE8mNwRFEavcA8X7OOAs1L9w7
RmcSasBZk3Cn0IS8J7FUSvt0Yr+1Pc5XHa3t9urEgu8GIrv7va0T2DGQoJgED1UJ
Qx/O1IZ6WpSRFPsEzaqsdEF5r1io7SJSARuKHf6kz23oIcpp1ya0rKOaEmiSqDLI
HuAp2pNJii84IGCED1WCEkSA05kIX1Y5MbUX27W8PVSQUF2OgtaPGP+xbO72vnB0
LhzkoU1PYKu2rrRcXVCLploC+R/jbqOyJkMbgx9sG1ObcdaLuDrpcIIhHKs4iQin
B0fenXrxGyHYhKvSYck65V9Uwu010zAESEpNBiKGnHmfqlxy7Opl53ImE0skrB0r
qDHSpPJ98x0lm4Ef+SQVCacmM8op55L+fR76Vx95godLgG0ZestLAQoZ8KEtaRqM
aon7jRFfKZ9IHTo/oqKNg5Lwjfz7H/8oFP/4sfTP24yphj12kJxbM437pjTb1XYS
PyEuT5oIESaL6wQZweoIxHudIvrECj/26a49ZsA1S2+I6BHoUQ9ZnbSPLCxJVi1e
vtPbrEEeJ1wdumpk2OGAQNJF/ui3k8EAFA80FFWQt+/VrQTvZy0YxK+tNylFb6uD
4TVrN95/GHKvfur/12kHMPcGaBHEAEzctKumFNYqmmTRNuS/MwnBaQNkL3HQRGc7
8bVs7VIyvxmYbOr3+i0RwF6alGD8tr9te7ik9HDU4hemYtv+QLyxP0+ySl//87dm
cz1QgKr60Qkky/5Tl8A22ktk8QRzqM+eizlxIZMmW+vOymn3N+kPigvfAwVixxO6
viOIQ3496LFwmjT5pl9/5hIQqDZ/XbcsBHWuEsXzIHSxHAhsd/w+/H6QD172954s
XKse2TVBg/wDISxNLVp93s9r4EjlvQTvvW5RxZw8gpCEFPitfdz0K06MASlil+LX
/LouKmbMjE7+HsoZi5BW9GKCWFrCNyN9vR5VRvg+Ez6XWBzjy74JN+LleO1JkofD
Ze0n8v7daB37i0aIcTadb1ljht/SO2uujcIEkRKYtxra02+YQEuHo9VMaqDQLIEG
Q59DYA0oLLjY+n4lmJWoEHw3oW2lAOJOV55lBLwVsARDzCkRHqLtVJ9ciuAVtAJ8
PVMrVFh+ZAGHgHXu4aUv8cCrG9SgtlwCTR2MWyej1avHQrU1EgPcc+am11ijJlwM
g/daN/CXG3AXlKHIfUT2BZ/QbAk1LuNEzFkO+8SxLFoK5++m4TCJ7TKkBHaUNvkx
SWr3DtDGCfyE7i1vMTUUrCZWxZ0u1qWv2ZJqqWvCxBLqPda+6xZsNDBWnVAglNJk
JyAnD/kCo8XjCoWjWcerp1JIMLAw3R8wZsAxx+ycSNCpTowDhSmwNpBPUmMNMIEz
oEXBhIb6M5oftgG5aWMkwnIvOHhNWk5dFHH+RVgUplROl5oEfkuLz2XiCeV17DfZ
vKSxjqPqvfsVnS3GxAcpRMCfHptFi9VrdoMA6mh38bPi1cPITKRO8HLZ8MmX6UNj
El5h3U6EP54wQkomDfgolRAeSSrhz1ui5zJ3Aflse5otn357CUJ5H8ZnjsTTRY/l
TCio78IQHBPjxX1v05rki074R4IS2rOxta0p4MH/vCyZqKT8Iocyg/J5tZcCnWss
w1WZh4QxbU+oS00iiMX0o4rr4ZfkkgL6cAdTrA6GhEYsoPjsXP+gZZMynmZZ1xqA
unhRTb410kYtm62ulxfTFBWw/zCtDPQJ9e4tvIM2KKOO67AntvstaPetYRDfiwOh
hZIkIlr/MvgG24urRRTQs9hOGc9EEk3rQa+ns6PYtyA7reZfpmDSTV5/BQIqizfV
vLMobkz/PAS3sH+eGvB+dVOpJPcfD2J+hdLNk6BpRcdO3e+6JKcFd/WWd0bVMMWo
R0lNk5423i5uNUfR6io0wkciC5esSn9E07eiChofAM/g+oochnbaCLHykrAOgRDi
Iz0QtVmHIeQe74r6eY4RbKvWnx+/nNyFQ06RvysnA7OhuJh0JGA3lGkx5nvb86/a
kdQdIl3LHElOOwTOV1jNJYSoTzpihMKIfiglrrt4YxW0qie9k9Vl8qisq8wKURfF
dlDil7j9DaIXsDVryUrS0rA4B/cyi+ZzCJ+Ti0ta5+iDCIqVMqlubnb87QZWTo5V
JP/OxkOsbTf81Uxk6VwfLKG8wxN7frXHhyXFzfqgQjHi2Wr+ZQbcJ92kS5BMGwX2
SpMG/4wmPrai5FAeqNwpkvatQC2UsEFarhgpJZeqPaw3lWea2b80ILL06KT2yfai
Cybf/FasrC6BN2feL+4AlNrjFK1/8nEqFLSKI2+EgfbKHrV3wD11ooxIfZyCtbUt
q2HtlVQVBd5VhC4C3/Y4ojsbh8vG7ZKr0ckN66Gmh4Kws/Ldsx7b1ORx3a8sJztD
DJ/jSD57344iCM4M13L/dEj3cXdvLmwTJNsC29MK36wuSlOaaB+VJNBKROGgthFJ
rl3+WWBCl62DOP80B9wpduie2AUdQzcC4jZrq9Avugdf0aCib78irE5XottwsUv7
6L6X6kaaR9DlUyxzrap5XWZNxtg2qLBHlcrnQgTbLjftshq5MOuscbVA9GmRsQZf
0soHw6oj8KP3mdG1LllOEXg7nWqJQHz0kRvdU0HIvOfWKe84pC57s5zPJnO3Qd0T
0tl1eFibFONquD+wZqUTU0N2Q9AX8rA0iy2FiHOdS7d+PdzM0CWUcHLRB38r7yDD
1Ah2a6Vbz94CwiliTnY4YnPbcQa2q0Gp2nerrriZNSMlxFVAYApYU3kRQXWpeyDe
peY/5ZPQ7hkCpTcDitbpG/jb0P99JeVsF+faiOs00ZDHnDttHcCzzqQpURzvlFbF
BaiCW6sbtGkmxuoVEjXp4cXncIVWA1L8rDALc08Xilpg9rZ9cvKvT8pQlZeQakc0
UywysTJCderbd2Y1kNYzNjmvznFExZMOsdq9xtdOI5/5/dtdT4PKto4JJ3DGvgpl
1rz4kYiCOTy5AXIB8daz11bTF+n1gU+9f9if5ONRw6TDkeQtadtwSivfrmq8Unm2
WWsdrHqgTOJ8BVdiNw+XXr9/H5fiTbQoobymiTaIZNB9vNPxrOa7425qTyJ/8bib
9RWGb3YUzS6gX3WC07avwE2d5mCMIXtp0oO9yOk2gYoFdK/KlWlwLFfKNn+Rn5Fs
tpaJeU6yML+Z28XpKRtDZQo/9njMnn6Uwm03XBnAcxz9I4na+YI4tbAGnJEgph27
9C/SyT4rFfdL6b/mR9AvUQ6KSygdoCJBCL8hMDsg0etjueKdaktJ3ciHsmEWXd5o
0VGXz5EqoVq3ARzKxJpp+A32+W0uiAF2wwEzcfqOsH7rASOSxH3fqn0uemNKyZp4
kyurHtJX3DfRpH1mh5d2WV+X26Z+czMXDoQOmypdQZ7PGyTOlFkthRiqSKMc/LAw
yXWuH/Sk4+7AaS70Dkb/j46viURLG4CyOxO1rjW81vfhwexpP3ec/VIB+HUoGmKD
WI8qMYtFyilwH6bJGt2U99Vu0IzYVWtE3FrXqdFaMZLQSF6OzSBo06acryTOTD7z
BMb2kF5hvI1h7ChdqemuIrsgaI0hMj8dbCkZqKWTJdWygrmSmk8pEY6S1ms3lbeH
Gv/dvGk+/sIM/KWSi8tZN2VR20Pda/fiCFI+FZ/rX0mh6ZeDDgL32UDgVxeyEQoA
mW9EOWNQbGG7ODTmebN8lBRqJG6XlfFDGyzW6E+4qgOb7kuaAO0zz+b26xLHJbTX
NaIuJdXAaNYm0uvBcsjRbTLMn7c957ZfQxGJH5tyVHM9nQBFKQrKgxkNds3aWRrU
cuo5Sj9r3vKGkRT6tVI3Z1aP3FCjhbm4V/DxVMNFHXMTWD4rgcX0rmOwItOPOM5W
Xn9SJ2tDZ5gbolSFzZitWcs564isqf0Wr3nZqWBvmYU7i6OgVZniwCvSvkXci9Y1
MJEM1VP6L7JWC1a5YikZg+t/A3Dw9D/Vpd1DDshMPiBIs1sv+Vd8GUR7OCq+iwAe
92egVYRrA+98xtxtMFTkcdavKaB2q5lSZWFVjmehYq7/NEE8FnG8kxCh4S6Wl1Ox
DsizaEQVwbgmrrkD8uspIkXKtMnw1aHRCWvNK/qY0lEJCBQn62Pw86fTLT3fXmMH
RVL8HRtUnRvIc+fpyXSqehF6H3YfeDbCi1S0SyOxil+ndZ0YYz46qlMYd1JEfDvb
hEEe3+B3toIvSJP5OTmVkHEekkSyFMQZ2E4PYjyGhwn0cz5ccD9fhgupAGZeAPYP
O6QDRS6kISgxW0FygDoJKfa41hxenE5U129HccOlPj8aFTMiMr0ffQZSlRRhkn3j
AmviYTjMsTSzEkQadFwkHUwBeteTjSF85KD+JEhjj45idNuEp6Cd6X95N2Iy1xbZ
h+rGT2Qtp/sav7ltVV/OHAUMfDR6jr0/5UZXkPlF4BNHYalxA475gMjxxTmYkAqw
Y+lo3fsZTTD+xa5AT40AWATqwK3napfhks0OZ9QUcvOqVfKjDmiWDFfHY4SBPwTs
0BHEEiH7mmzPhsd2Jpr8761CTtDzbuZpY4N9KnFyepGF7AW/T6QOwRmleZ7VBQPD
66JZ4OL5dVIceV1srLa5o6ppxs6oSlckVnyk8NU+AZ1fV2ErLlHmWU1mj7VrHQgu
w2YMDGhQtLm+b1QIcP6G9zi3EwIWJdVHAgl1Pgz52ILp6CpQHMKFLzosRIUslLT9
gBfJXGxMoNzHPgMOWJPqnAd2hq/y0vTguluCm7TIc14C0JIdODTyNITymnrTTuf/
iSvVUaJdrTUcuv6Y0DYghYMTq0oqForJMbqwjgPmQxB4HHzPOUvVq7Qv4XZAqLaT
byBLu8lmZLmNtDx8c6n6q8ZOWzpXvISUgTDLcMJYbi19U5YDZxzyRKg/9r0CFRrd
rGZ5KK++opYR8dOTEW29L5GefXaZU5DN1R8rIdCba6ocCqx10NNI4dgzUoxBrxnX
+Zvc+x6PTppCCWTQ2v7WKkXLMtHHygEGpFyQSr1meuYmE/X6X3bGtYksQ0p7WPG2
1IirwPiP8wZuvHEC/79nQuxaB2dTP4mZAJU59CXYb8hCnJUbrGjYTW0H82gWwhBd
21gqxntZqtg9WdpKA70HBw9NvkQPyd13FgodZi58lpQFoNGFBFkieqCMsrONlRmV
F+o4E62hqtXtxrQHoA01ZSo9M3qSHmP1ylg3CmR+XhenNK3J55cGACoVtfyO/8p9
rLZRD5WJULMUKDyw4ybM2BbFaIM4v+Y1/xpoJ+s/1kl915EcXTDk5bCErkli34UJ
I2MOobFLmpbR15PkzCd6Qcah+qo/n0L8w+DxyO21e5snZfBbdn/ec3ygjid30klf
fgTI8drkkLZI7IbXsO4Dy8jA/FMiTvtvrpeGbmW42ot33Xm5mJ8IQQbi6FuZI4WC
Ir8TKcWvSmM4cSqGIa8FoEKDlQQLBerSbcFmHIcnOxXcJ0PSfNd2gVUzdi5hYxaU
0WrQ5xu8gagZ05fyPj+NfPWBihzuY3n5B87kZaBhBzJLSTRCIw0O1837+3aCGb2z
hGeXzwFh/sQmw2+bud8QebVa364gdodNvCPbftomeKxJyPocPiDETMaNmGLF9e3l
F0ykwOa9NLe748THdVs5c/hiBjKGY0pKZB3tg6chMIhvyBBk0n8Qke4AsTqXdoU0
aaCDVxZXnCwa7jlC4HsrIye0vlAS11Bv8Dwcc7DATGkUK4V2zmVXBDAX5jAphzv9
hihEMxXCK6ntNXwFsJI4LxjA5Nsmsjk4NU8JCS/rlMc7WXJz7W6gY+vIwDAuRl5I
oyd0sdZ38MWdSY1S1ftm8dRiG9MtjafR+r9LGhcLpFJoiBl6KW6Xw9HtCnuBH2rL
8LY63wQ1o1r+Aphn+33s1bPEHTzNRyqzB6pdV1gJsh5ZBKcAeqFZWZXMY0m50A48
kj4XPCF58y7YUDNKb5Mk0E0yosa4tMfdALwkNYkVB2OxIYNm0/WXHJ6ikw4u+Asr
eBv3tG2PPGJmW+IOYtWx39O5w8k9Bxi5ddZoQt+Ats8cVpHlJGtGUcFDLNqfQC6p
JlzqdePehj4xszxtpNFB7vlSTrcGH+/j7DH9OcrrJtmS08itdgAovP+tIOMFkcQ6
wfgK75zREfBRlZD/bwXgbG7aKRtNkVOvyFdi3BoM6OmLFfHNXMUIvy00eXLZQfmL
4ymp7TJGsLDy2z6ebh2Nllo5O2spompMVKFoOYewgtVVVqLIaEtKFZ1gMDpE21YX
0QQwX7Xs6SAYlY6x4Fnq9ebDkswlqRsHhPjGejN3UvacWLW94HW2V/vIR6wzi6wk
qVXs4Ytgin/+GW/gO/aDk4GfuGRsmXamQNL3pJ5EJqF2/vuoOznZ6hvWJhPvG/Fa
dn+8Gm3MWiGLA9KW8oTMoxeFMqQQkoWqenEhHz1KOGMzLWMlcU79iJaeOCC4DkH+
1hW5I0V7F+KGOWRCOr8K0cCYA7+ZbA4oUH530crPRT5fVWfDR1XOXNCQ+G8Yd5ES
Vs3P/zRDkTvr7AA+eOPpwGBpoXuL/2ggUzMPZtJXE0ZeYrNsydoscz6ao0ifgvrw
T/5gUOwTDgZoh6FKUeMyWXcO/YD7seIF03Dmynr8/LaQVqOoIrmiMXIeZe8QMHPt
x05R2TP1Yhp4bd2YmeCkyEzJIrDjBBbsNyh2fDnLQf4pgMW9Uts6RCuo187mxvca
7tI3L9GH6qOKF5M96KJdv/hv5HO9jC94532ZBpmj+bH3g5q7CgAiF+ezxY6Upusk
a26Wcnu19TfpCbIJYYlK8SryJ9FOIsvbYadhJasOLP4EI7JPN4pNDcgvZmpiNhRZ
CmV2zEF47CUkqYjjOyHBe1diAmCsrC43WrAzDgOHokoqXJH6a4c/lgx5v2jvI+Nh
Rb/CxkPAtqyhbBdjYDj1QSkpYBNkIKLCtCuywoSIYo5D+mgyxmix3IGGlrkcAQ/f
0IMnjtZnawKhCDyyAOaA6Y7tIF0VqArjFxU2xBizXlyIJiGNlf9FinHKrAO+h9X+
IYuvekedqEx3J+ok268OYOd5lXNodmazlH9SQLlcOP/2HnUdzDthbhTrQqgfgnQh
ViwoAhG60nkjc5cy95J4ohsDTGxduts3xavc0HL1C0BwUxzjzMyVkZ4Pz3UE1teL
3r28ivXpjG2cR/TzEajuf2jNRdAeSHnx1h7a4SqsBnB0tm/2Pds4KM3+ZCvMLRGk
Wf1kZG+IXH9kRwTIv6g9ksTceL/z7dRQRBLuVv/P1ybD2MeSNy7sB8aP0HIL6BRo
FT3MCuVmIZxuKis1uwIc8XaegyWBtOpoGEowFOsggDz0G8FW+F237O2bfHyO5CON
GIGzqC73cAVaQRrmdRRkZsHyFDRNn2gTfZIWhmLQJbBCV4/jrVnbNqW0ZqELOMIy
CkskDLxKL1caOmo+08YAv+L0mD+g5pgXNBfkbASIFXOFQlbEUClIjdUU1agDYMgB
9HzrPt/c5XEsqnisRCsZCC2NmuCcJ80mAMdMu8dzA191k8LSGpgxbL+qJf0Pwbli
PBqbofJ9Sf+l24oFl6rWu7LhvV5gpDqKMg0jz/Vn6p/b9LzrTe5f0w+WMxZDael8
6yQuLveMayMJKJVeeGspaaMvs4/r9o2hA+dDE6bhnJXQ6JgLjPkyYgplqT8xHKnj
qDAG5mThEYRULXCBL/38yT4LaV6+KBDRaNHKlfw5KUqbrT4nMVFm6MPIfj17y5+O
+JciRHU0bLmV11sDpPChqBXD8Xx6UycPGecySYDJBUOLk3EXSG9A+w1uh/C47lQ9
ZY1uzQG1lGFMOjBB5W8o4vcn+OkWiGSH1P6/bumuVakHyL7oNBeFm+21UBOzoWzU
V7cSiu8XrjG9ugIm8P0B92l/iiuaTSeGg0JDGALovgVfsWpvz1yuwxfHHP64CfhZ
FRwlbP/pDrXrB1GmHO4fg3z4OKhabes4dzsaUk4iBOHiNAANuLmi59XkuGv6x2aS
lG4Knji2Er4VffCvkOV4lrlRIKqgwR10kwEjReTie8MGbRP30uNMlnb1AaEVbQ1j
irMqD9a2Qfx9jpFsjbPyEHj7OtLFIqTfBO4BUI5mO5Ubp38UsrUnd6/duiuxafCu
8Xg6hlYsu1nnNfMbNr4GBlHYLwUHO0kl7eQxR4CVtb24fekibgFR3GyQB/yVCXvX
fU9bKzuw1//EZSHLFRwmCs/OOaS/HBez8W+2/MY5H0spyRZ/swkNV4b3tREePIIt
xoOqomHzIWh+IS+C1KoBYJm5NG/AfAoz8YdGz6fT+py36hH70d86dEwPVTYegvg/
XlH/EiCwe5zWKMQyoD15W1HIT7dbqIxtJA3p/zjaskSCSP8+JRKjEy49gQ8DYsEP
fs+wLHX+zFGVNHOWn87IQsAg4VjR/6aAYv2XodfVxBup3T+dMF565lXhyN/Hh/7e
KcPdnqDyI9opiclf3lSQNRJ3Fuu2XxOVF0QY7shJ55lbdqBTDAz+1zsga+z1We2R
iYlH21nql7xZIjSLAOWpyd91U7hxg7K7z7rvvVBCr0g14/HDMeC0DKK7NaicYkvs
DAkDj0ZN3tlM39Y5ZXVgTXOEUnFEiLDdGE+vnALW4TvqvOqYX23fSuPx1SAdck+O
tOYlTgKf0SqPJkizAOL6uuHhnvmairoc9VPbH7n+vxCuvSmw6qeCrg9FKNX1wxCc
dgOR1yCwo0Ofg7F+3XojnjrWE9fQwr5NbkrE44kHPP+CdGVWfEIBAO1nyuOJprfW
4pzK9zdPEB6sZHI8M3tqM+dQinzc0L7ekbGT1RG845Kk3f+heNgWkN3mZkFXb5sT
+jj79dU9WDPhPkidLSfqYJHgeIgneBklKBEX//fs3SxBf3mzvGxI/zu8ebgSSdhK
r2P5m3YxgWrRzZ9wPZZR2YI5wN2Z2YBzXZPkXE7tzDdUl/rjA9LIsnyXQcMWFDxb
ArbVE9Quk2YHbMR61ZTu2OhFMQSmNmQ3i/KDhKnZM4klWxPxH/TO5ZtyIQ1x8+9A
/cRRBpEHD2hnIAwrEkgHTq9VW0TZFb+fP0l0f0ZS35Sy/IIAHyRjIBmyjRiMZ5mk
aCcqgwNk2tV2sB18yKM8Wzin/h9V2XZGHASBofdJNTq8YFj/Ng8GdZFyeYHAv0KZ
YbIyo5H16SwPRZgpImIIaDltkCnVy/Q/hMCEDp3FGLrdAwpZDd6cEj/mFixrj6w2
/Eadggw7inLTNK7unNKpGPupbjPAgxUHbcfjS12EnYTkHOZLpzF0KZIe8Rfph+6P
GixVjz9vhEnE/6eQv2hDVtkSUIQGOoQwBk8K9DC087r7kI8uNAxIaAxLK8Z5cK17
OtHQJTIr97DBN/bXge3vunYFwy6L2HstP1wkGQvMgDsbvIG4fCI6eSA6wrMwvEdg
s2uaYdglBZQBwHPkiwPrTZIEYT1bpwTkjC/WB9XI5RjNbu5fAQvCPq5DMM6MC7ZT
55GHRUcixiOJRITq9EG8z545oPxYQuBCc8x9pUx6u+mmcmd9iMM+gBIMReQVAAs6
jNXmREoWjfQHQmHhCmuBP7+hoY41vYn2HJd2juGrPvo4hxfnB+zOdsV6aPLhHVY3
QPW8TvnEWTP3+aVzvvTzPvGjd3C8FJ16ls5V73YZ33dYHZKapxLYzqdW2CBqFwTQ
Ygj06OaMipNGwj6BIUV5wA/FMafDb7Y9HqWN07cHworhADak1og1YIJiTxszyOAL
kqFKEPcWF5R4bYiStlDoaSpRBiz/tzlR0PVRY2xvv1QOJ/xldKHc1t9TJQmwXYEG
pQnkXf46sXydxlQa9XxM+QTy7GViVOUfNy6hSRIoRi590rwlvYqH4ForgzzbWhCC
yzlo/oKrPxEhUb4NJviUWie9wZlm9+9U1QLqxAPJBHtqjztLPD5phv9/7nvYdAZU
8fkQEdBhmZXtFaiu7NgM+m2s4AQJWUdpqsTZi3LEuzIk+icgLLQbauhWjmpQXJKi
+1hEZQCIdo1R3bPf74zogNaEweSy+HsS6QRVU44GB+Q9yttP7Dcl827pphxFS7k3
vdEGBrQud3GRYssi5LGpj1KJRs2bUzeX9Z5bdXc8tIhSGZx29wsfvdM3XuSGQvSk
vZEoiUyYRl/E0Rek0E0hDjYwXSVi669o4DgJh8G9zywgbVFXLxkE6bBumZ6v1CPi
joYwUFZvqGI9DJYfpFF3exSyeO/qdNbluEQkmNrJR/dNhbSksm1r/liEILLamo9c
6ynjmbC0WUau0WDIrqditTqmiW+BCmzM9oeXRZmGuCoJAYPR8c4FqOBxYabMNav8
BocpkAN7fBO62wcNwKPoCWPAVc4eE+3Po/xTcGMJ5cFDKeyJoVG7ESlxVqrrI0Jt
Kv5UxTFdFSArzr5HrFxykfDMdf1tui5T2wSkOukfnDOXSdbjixUt276Lq4CHpXEB
0/6LCwS2p5vnCQ/IzaoLUG5AtDsGd5qUYsytz2JgRwjqXF2iarYTBzSDV7yIA6zn
ph3xp8li6fgChH0g4kn4dszKiKMps05spFp/JRujGGSkjOpYMJJGyQ75r4Tvvg7L
JuH39JvGHXM3qxjoWJ7lSs6PpcSU701kdXQOs48qKPBKPS4rgR91KQyr6tm5rk6g
R7Ow3lryAx2F0aUZZY1gcKlEA9L/H4qbKXNspI0WepdQcQYK2V4KC2G8qgohGVPb
maTsLSWpLGvVCbndInANeXl9kiN+1qtEak7SIS7KaSGzG3clhCcxUnLrlfEdPvgF
sS2FpIEkhAY4yr6x/YEETaMMexM5BIvVg2EtJ2zbv+oG8yidy2tuzfXlKikbMCDn
r+W9R4Mke7uffLlLTfWJSAegw4aPmWtmn1nStRMN0vQDGHTrd7kaBrUyvml2fnn8
oLBEVIAfckyrkGnGyZBgCwLydqEK+qNebXWFcQr2FvXD+IoO1gE9TQw/gtI6vUtD
cmjBTsWcUTJ96rze5LO0qnpeoIHCG7d4v7SWhjGdaPKoR5pSfg5J3t/+P1uMAtd1
6YDuLjoKCYctCCG49XAceOyzlCyUqMKfpuOU66wbG7wbARwMP0GrWF+jOR6CWyZv
WByjIw7zApbAjsH2nX5u7Xej/aG1QBKY+FhGWNPqvSqv9UPlMOwZO7n43nFJtd+G
+MZMb9hubptd34HuYfTfoo/WuE8CsztL0/4hQgFfyvkTNjdGVZfIV67xYpmGE3Dz
q1zY6BCBo0iQ9R8xuSxSH4JVy2+aXrptWZ4J7C9BNzoYe1ONiqNmcMFUDV85u3rC
54NaUR6ndMwzkCtYGoPdl7fwvR4IsiqYSty3hbJbjl/z37cgIuxXFJvKADPIfiwL
Tjx153tmHupymBwys11RPyNPZy4K+OR70gZmj9zKtvEojTBeV1928Ux14r5SoUa5
6ZE+12WmcIXbskTu/L9CmGcCcwaNDB1aPTfEzceD8FPzVjBru9r+U2tPYMEr0aJf
PbE9fB3OpSYPZ7iXx2eaMpbSgDHz0nZV2p/8I5tLBoifPrpP3mbAKAcLXTeHphUv
0ZkKKIxR8wM+fk5EWV/oIRtwHpfiAfzUY9vDVVLGcaZQ9PuLth5oA/98v9Et6Qis
Jb4K/KEaJe655Xawl3+NE1SRBJEmGBtOCBSvuoOOJ2szK+M9Om71sDyp8znFNMOO
dlJMDtNgBZ4ctELgTap1BtAIQgXJWdE7OtWuMOBC+YF/YhvZHmv761et7Fnw7zpJ
x0l7+KCZJDhKQON9zPK1mgPPQs18BfnH5c5u1sA5VCPVfFYghwP/dQoVL7J6ojkW
KR1/J9YkLJ3vMX7mZ10OBwa2oukIeuleeLaW6P/Dd2h4BXtQbz/aadxAXrGVTh9l
Cqt7s/Ow3FZfOMJTfqwdHFO9Zr/OlFpxdK185HscWVsiUbYTTQIIvBSeSVsttoVY
hKcpOofCT042D3lDM5858fQAiqWPxD5DUHVABTHAA7Ljf2awKJQcj2lf4zPsv4yh
7eiulou3qvf2mX678k5yH1yM0JWCfuYgPwze2qoIKYq4j+WaxSE/llW6+cvlL2z/
a3e2e831SEydKF6gpk4CTSM9BzyVTKP6ENQdrZYD3qPu5M2eHcd8LlQ9y+d1XdQ0
1TUxZTP4hAter6Y6wq73JhljsMvtMnMZQ/hdz0e3UefPln/bgNdVpd/EvTeKPtIS
zVNi9DXCw3peAyVUZWSMyls0It/TjHBY71TImK3DP1jqaFAJpW7NTHKJJuUjXaOT
wdqwapTw80xQE1X3WdRm/sqfMnvTUNp56yBRNMQE0JVwQGNsVGBjudtYLLlM+DZt
FAA/OqR1ElLnCmE1dgx45V4LhIyxcn7Pitg0Kem3I4egxTg4Wvn6N3XwYzC1rSPY
hMR0d7Isa2fssVu/rWLRD2AyusuMkC+wqbGYBsYFlyLdTFisEZ64ld6fKim/SLpM
I/xREe5C4LUvQYjy5W4tA7i90l5sY+P0wZDUFjAxAkmkVgu8/3Rje2OA+LC/lwhp
w538bFCmWQW0G56qskWtKj7uGl2fgVPiH11bacapueRogljBnnXRSxOyrpd+UMO3
5R2V00rXWK4LMlvPXsPm5XiIXn9mViioNk1uhN+jbnsoq1ZtWroyGrYAa42fQN1S
ZYJrkvQwJW6et2xjbLjTDGJDEz+l96i92spvKSsmN5nQvViASRF3O1D22ZOl7u2x
LuK0tR65pbsb0H2JQLTBsaSAWYNceMbcU3iAfGeHSMWAvpKrlG/0ArTbK4FH/SxH
e9R/bvEh9pHCIq9SRPwA7q7NaqsqX6/d0smX9/Zat5DyF8zU08mBlkUEK22t4jCX
HojCHBSDjjTUlIIaLgv4hAMDLk/Tb6qTo5e7xtUkB63zlHFdvizeN8YMaFS7HxPX
BICyolRPvwn6Xrjw6aQNGVnsts0jnrXnkdMZEOjk17xFxqKo7ds5rSdk2iYFNoEN
AA0JQIvGUct9/zDG1sSHRfIPyGcfDsfgVgyGd5JyZ3cFOeioJipfRw3CYNvNKXbV
PbBBQKIffIR+fu1bBQThwnaxenn10YEXCqsfb8UuZzA0KlI1DHq3aI23/kudMs1U
lspoK08FTl7WOBV3cYv6dYJ4lBrxW1OvmQsln3bdQfBFvsdkZvDznea7RckoTQ0Q
lvKDCCPdR4n5znoYpWLCQq/m0nF3uuiNQnsCSL/R3xbxh/ntFNZDfJpykjySjDpE
trK+7PtV0SnJ3pQRNgilpgLS/fmPu4LMqVzdyq47GNu1HVRvn0zoPTEM6Vj3kg9R
xyZAuej6jGDZiOYUezLuV8f5bwoPQ3LFtWIL8ZHtDMM16z8ri2+hKckvNPHezjP0
iBVOX2B/xXNhQuckwjl5GwM1yawWiG7y0vjErhl+vG92XdO2BfPzLFwqhsgQVjvr
TvUoIYLYuO1gK6QmZvojhm44RETQC93/B0YQC5ioy1LUuxVgHjxTpjoiA8dd2rcT
28M2wxHUmqfxAQTglWoQFyfmHjeybiYmRN0hh6UQ5A3abir0siZVoZhRNzZOvc5t
5qMnp3iGMKNoPJlSx1BUv2pN3vVgB3Y1AnmHwba80EJGpxd9+j0bNwoMh4Q7XCOc
afeT5rpWaU0TS2BoyZPEXRNLeNsDe9CqHASut/ngjUw6aJOuXxZhsw2N3PD0Yb8p
MlXqa6NIa/mjxddqX4LuZyzD31cvh3n87pNe4ip7s6oB/5N3TnxQluz4KpSd1L9n
nHHeIshBvi37ohB9e6jCs1aJfYOc7nEoS8ANtyRv1A9LmkwXgyogVWIZYMXxBfWz
YDq8pgz3Qni1pQ4XEZtUxd9BuOyUpaKsPYUgHOOABbw4gcy3FAysj640OmlR4m4R
sZR5Y1VRVOj9DZOt6n/RTqDO+qlSNJ4iDmggiuoPZN+JdBZUufiWT+nlkceFCBIq
ESPVE8HIggkd+bJYLwYMQBfphIikZR7H1C+e/A3c7u4wpDvf/jNeJfceAfvyxFuH
ESEw0sBm3gn/DzQ5Dk8Rc1SEhza6dbNCY8T3V+TTIQpH9UoHjP9gj6kI8KKSEsCX
gGAYuQ5MlwRjHRsW2Ey6qUUApIExSiSeiDumXPexffJENUh039OeSIwjKH24h01e
X8DMVAHxrIR95mCViK6pte5YetCY90+OU6X36Ko9C3HeMXHL0ZbEgMy0do3ql4hn
5Gw6k4QVtMOV6oh7BAoMCjQa+BO1GpVSFQnSPefJwGRqeHXPuHQRMpgeQnLr9X3S
zvlWGygMg+egWGuhswmdTHx8sAOTuzgkT6vZ7LSP5fjbOZU1/ydD9iLlmX7jp7rj
PByOJDRHccLWNGqU2dkX/XsYA7Olo3t5oDPF5Kqdboa3lNWKCBpvFav+Yl+H8HKo
XNht2iV11/7fF9KDY7DXREnl2rdHrZqipxxKNv1wcbqhDfnnuWy2PX6hacN6ovnH
mzWXKBdDp7KHRzp0R4Us1/BjVYj8DS1p9ppmz578Ch0OuYN9mwO/bZKCINYdrPKm
uTYKrT3ua4uZZTTgxf4DnsAeN+Yk5JC/ZOhg7vdp5ltcR/alp8gWKZEngZvFYvtY
Z/MvPpDUKh3PJEEOhPfnGZGoworhvubYzi2kSzBPv5hyCiOWPZ9+NkPqgxBLmEbP
XhCyCmbQXBxBxNw0ncHjr4mhNXUg/K2SO/yci4Vo9Byl3lRtTTeGvR3i1cqyGDNh
gRJeUtgHr0JjIzk6R4dA3ZNO3d9JP5agsN2qNpmjvD57FCKns2N5jf/BaxvnyqaA
ryB13UJLD3mdzklkl4WnnNAJj36talZTpDgZvlfywtfYuBNw0OLTBhAqb900aVFt
mFzvQQvKfeS/uoaI19hKf9A88A8+xQbFmfWoxsJ2uUzZXZ4iNiF3NE2GQncBWyHQ
/Dbjz+wy3Yuv2HAZcyeVG+KE74fxwKpMGzhcxmrexjP3/+Epf655CbPWMoLjBE3o
Q7smVnalb6L9BKQO1E/OY6/dNpbQLITc6VdPaZ2lUvgEulWiLlUr+LqYEXwJ9TII
F4Y8SHRcqOZFyqt3lnYRhjBYiQNofcyj97hMskENyJEZVufQLym9BGuiVHfTEJPF
XRPOKxupUNw3kWifUNuU6dYYKczVNsHSN8odH6zAfkTnpihukn+/muEpTSBfIiMt
tPXTRUmpmAk5yCLeammScN5wP8H22ZSlYbvd4+YPnRF0FE9ODyn+zzmOlRFIkBiD
qFKBY9J9X60ikGXHbjTXftNFqG6VDgli2HZB98cR+m272QYKDGMFeC9D39XN6WfB
gmHEQIVZ0Ffp3nPBZrSU2DYoyRET73eMBb5VS8Jex6ApSq67GcitdMuwUusJ26lu
fgirZrPHed7zhDJ+0l9yEZ5olaRyrZbX3Lt45dkJfENIa7TFwE9/zjL73x8oQAsr
HzvVAvts/07Hgn65JClNOb8XHqUFf3Royqt7Ah1ty98P6l9upg/dnkHtSzg4Msz9
W2UK7HH5g7GzLlrzQ82hXOoN+mqnc4LeIHrONuAy8XxArS//Bf4kSAq5PvRKjH7b
yY3L7GyqHZkZuCJP1GW1zcBltKsudVwJedCD+pfLC74jn/NMS9n2S7cw6+sGBpPb
lE6e98iFtCHToJic5KrFsPQyGcCUWCayn/yvliHVwGzr2L24B/KHyq1aYWlFIZDF
0hC10GH7ZbGIkRmYc3IAZyHjRWdc3IU2yM0TvQKnij+TZ9I2qFN04MbdZa6F07th
UgRB9Kyv2BMkFyzjVvJbxtMVvN62RugDRE5Sib5OxxVxh2Qg6k9uTFntAXbYM51X
W2iqUtcVxvSrGQEJYMcC6dL3fXypR0JJf7aOg0EEzHhm8iINsqecdAYs0fW9pHRt
e9iTBdP+50FsRnqsvOSxmZuOJkb+zpZHg6ESm2DnMGwbGhNavhY+l5IFe4zJWsZ1
2XxfhuZtp7ddOl8Vuq0ztxA3wEaMAb+u6K5AcGzudNqZI9bTdBIorlgrP7roZEMU
5AbXTulXMAn2Yj2ksAyFdd2khK7Rt9mnzYGTWAWeVwWSL1+br17t2T77Tslnld6x
vD6UOSkAAjZg69UeoTOVnYxgXl+NLehqhr7BFnlav7ChkV1YREEPMwQy09ihiXTv
m3lzfpobB9gIutbBYmnRxyRyWlRsdzVk3ujUMxUCbiBi1piD3iZp/LvGuKlaXL0L
POF1HV+RHVtOuORPwUxLa9EhI9fVXswmjQzb5izyd903ksgO8fNP1vQWvECUyW4A
cdv0J1/NuxPFKqC1g1RC7D2+j4zP4aUppr5KkafjW32BXaPFtUhDrimD/1wHhhYL
7GoeTkzBLZRDyaaMSesO+zrs+HePdsPYOy8A1QvpD5OhNwj73Y2UwRTnyemTb/DT
6uT5Sut2hLAeN0TXVZ3OMbmiJH6dBsEWyUgt6FzfNjCbz7k8BN/ICfYowaqv+h5R
x/QHCvdbDXBWlZYnqfSHm8UUzIOccDT3vaLCXvpEz3p0WK4jG2ks99SXnOyMHPD+
u6lPymLq72vM5ivAUZCESKk84YpBgIgXQMIJyn3ZCKr+Fx+BkSQ5LW5I3JVW1vQY
YZuPDxLADVjQHLzOHqoo0yFPFgGgG/Uc8y12S2TbQJPlb4/zgfkc5IbvO2vMQFML
0xNSV5hBiVl7igeMYRLpI+5chZl+4eArEgQko/XbFauWyp6AJufuO1wLj3nEFGsX
OupaA0jB9jRChuFzho89TGezyEBFBHfNZawsK7rrXcbTQC3yGk0FOZlNNmN8wnll
Atdh5FyNSLtg/g9a7PUJmJ5IDKr9Shxzx+sPAO8BXf0jLPH2jRdv2i91JHReyXou
CatcfqKM5ui4e29Jn0/fQ4kFCQw9WVy5cbCnwbBC+i/IgmItGRb14+QicmxpF4+G
pwgWf5X9Bq5eaLQZnsumwO9AQ6Gc8nFxLVp+pefcM94qEKewaYtD9HJd+yakoZs3
RJSNBiHnQo94LRuf+DX5ojNG425vYGmrn8pkX5vVEidR9yJlvD2KsvaCeVytYLL3
vWY3i1lKJ9Yg1bLn7cqb1x2pURsiL9JjGz0oHznZRAA+2pwdsehV0b3EpNqFyrYn
kbOeEv4Uxrbd/8jV5yk6Krp+BVMBFVIZRjgrJhmW/32v6uxhTHH5HvJddXkAy/Bx
GlUVvJLhXx0MSoIPs/ugFc5RXWfZvKWlTNJ9P2p/s17snuIdo7KlejAaAxk+QxZg
36LzrtnquOxg+pRZpC2EcwqTuIsmz8lAIHt7oHuik13PgWyg6rTD/S2jB+TQHse6
dS46aQM2fRX4Y5UdYueFRV7fMDjtviuiaNuipIRpRJ4ne2kjjmYFdVRKJPYRiiDV
IxAvV8mbAoZE5vo0sVtqVt74SPxhEkM5UMEEgZzYS0weESqm043lUDJVx207cmz9
Q0xU2PCvllP9RvF58Trfle37u+Rqo9V0mD1XiOFh7Ztteh14feXICzLKlK20p9YX
wOxcyxHFhePZURVEh0sir91n5yXMHAXSbwnaLMobyYt0alhI5nj2kEQAfKxu5p+I
o8NoIJLeswu8rr3b9RVEt+F3MxwTvtyZQ0cBBKe5JsR7QCmnLVjqK4PfKhjlDcah
Ss7If0GhiDMzpclg0XhfBbt/5YQAhR8t7ACxBg9ybvvIslO9ETq9m7RwfYrvOud7
ULKDuAxHcOEQKe2x9Y8mN3h4eKzIuTBi+/zvUaWBoUklG0d8YV+067MA642KD51q
uaQccHkBmb91smDfUwlTdDHJriBu4MEGw8ZBWqR6KOJAyOv273ys5W0/cv1Ucvt/
HEGu9k0pf05u69Gc//okz7QG472RMXeJV3AvHYyPCpLKlTxX2NqIHcqzd1kX0KlI
Xwo98b1hZ4tzzTe/v35OCOm67DgO3AtAyjuiEXw61xUEbam20ZvMkpK/YjCtpVrG
NXrr5ewGZ7FExYcCkj3EFatj3G6QjHcr+vUbEFdwUVBNxVlBK4vnCmhkcn16sLPb
mm+ifNeI5Zd+GrqGnXalKe/XneIJ9h35VzL+3PcjxN5RACeO8GRFxtdR4lVHENu3
8NW85XppkOXQktJHAGKWOJfA4exn7tju5RzsKd63XOWmqRVDo0Ap/RiFgYs+m54x
L1kD7ryVuTXXf6N1Jv2sAVN6uQym3NFzOAqWWkcGg83ar7SiEnCVlIYxwIEJSVjY
gZbiM11SwoEqf4MXDRgP588YHt3CKeNjX3+SyXC+V3UB3BgtnDYeolU9l7ABQ0Sp
mYfwZcmaNbXTQpO9O1U96GgwTbNKiJQKXGnn+6kQctFE16xuABQlUFCUn7o7ITPM
/zjs0uKSaHpaFYGFmTMbuQR7qgQowc0XAWxG2Lrx8AnlEfr84JyjpdnjJC4Z2Fuj
n+/5oZ49qPix721I52ge+p245mqG9Mmq83xleolDlUo9m568W7LNaZxbYLdl4ypE
BeMtgwhNbT+5FGzQaRG7Sh2nYSccIxRVSuJXHP/XgBmMvVyl9O3XyfvDzrEkjS21
xnszAH7w+c3cPeWIFhXSKTt+f4795y4bQYWpQ5t7Vkeq0g4kGVGpvjkZLybmEMLO
qbxpKFVZZy3PrO4vkGG4MI7Hbl8acIdExrLc0w0lP2R5ykL2VeLklpyc+EYwLnZa
TuVZ5IcMlBY9J3Zs3ZaafCIxsA+BBQXgPZwrsa3XhHA41tuDgTpqP3uLDUzETTHl
XYbF/s7fGnYwgaagJvOekjxetNB/IHW5Wn1cX0qrW/P24LqSy0leMlSg3zb8TrwM
OgE8cEJOFocPZ20YvGK9uU52I1xj0HgRfEAH0A8W8Wd4NBiKudJNXGgJ71utkxMr
/6/5oA4hb35HjCodIS4v5LabE/up3rmDmgHWWCW+SU+0NhYSN61IwxavhfPcJ+Lb
A8biC+6vImpZQTbPahdBMxcJDaXYsKjBZS/yWHxhhvGsn9MY7qFCO/JFZ1/i3rDA
WfpKoOPvcxhGy4jBdSQWSHS/NOAdjnqXISHkorUItwImzqF0UzB4mofk/P9ixF4i
0u2wUApeWqZSPxrHyDDngA+TgOrF5QlHgIlncjAL68ptuWMAXA9VRZv2mjqIidYu
sFFKr1p4gvvAwJQkGxcDq48U9jreMkFV6c/++zlbvN1Ge1r0xQXBhDmuSAZh3Ckf
8fiGhEsiARpuVD/YudINp8LjPnpZ3CAQaKnba7bCt3y3ES14MIoJ5lmivuXYFt/M
QT8WD2LzJBf7DfyXKyRG//sf1WbWXWDgPYkTN6SDqEXYQhhw3bfim+8WRJYoa+ZF
Wm7tLmAcAijLDYWnoIlfHxZPz+I35vzkaWHFRHZvINRs8tB28lAhViVrGars/NB5
xd3yBopINY53abKsA+oIgXYzR2a5Z+UR5bCfUgZ7xFMyYqjSoe/wUBlZfuM7+VqB
Eth30q1Mr+CEMBznCUBI0np3/rkBN8RlexqT7IHqmqAXuBpbYOkEVhK/GiiWFI9f
esgXV2atvY0AmxcDRLcOMzSRjpOlfQkSWuAECzTkFbPq9nkVndQW63ZC6phaoK4w
KUg5Dv7VkMmKbAPX2dFsHIMPUGtKIxRcJvkOiCMXyK7QvSLPCn3ZOeUFJYyAyAjX
Xf055jh+T9jmoYolJ5MPRV+DUx/HKLJsu38hmkkqVrsq6XNvxBkOJe0FpG3JHpr2
o48cMoWiG7dz9ZVuzN4VwsghYj6wC5X7CqDr78UrwJS77Q1BpVhLhRn9Hu6KOWe0
jYz1V4xCdmM627JyR0PHESq3aBv9Nz4HWWatKLIcXgG50Cv2euiGSHkhgnlBWn6q
fZhzs7WVZjpSWpdC3ghpdHtujY6OOuVTA0fFF7qgJYl0BtTZCiVTGwM+diIx0UgU
/1iNSrqlCOmnRYZCnFVWj6uPhZAu7APH+ZATofBJpkeaB+cKKpp6lYQmkSKi8aJP
wavnQf4OdpbQyJ8eIEH0Qs+9VgjoRnXz/6uPd64yHO1qzQ3EFrNlHGCkBbDcHskw
BU55f1KWhRsEmY28G9ojLwjVHUDhiGMsv8i3dNJfb8orTXN9LgBb65D+6jso1Ik0
HycnsKUkr4pWFbIXyzeLWjKzz675xXhgsJPbKa+H7QQzslyUh5kxFhKzXi7TJqmA
vyMODVLnHE/+dTW/5vtaeV6Fu2Y8BJry5y8nB/OzuTVYdkaidQDVN+b9C0VErZdw
TrhiETg0imJLxgstN19Q2x0yFcVU3h+XayS7l7TbOoucBm5Cd7vQCPhVrZws2YgW
yYb/hIMogMMcEmKpy26xAjQD6xxkCj93smemKjfEVHN921Iu8jVdKW4mq/YewjPb
aGYqo7ldlL/j+axX/e82ddUr3ATQIOy5jUd7BL3k+Ssv5KqNnhgg0rNTnkM8uwp6
ricp5aExfRxjPmobZtLlxi/ryodhWiQ5zTEm/QsUHEUoBUE6fgTaxMrjrzaDVr+9
RT4xsCIOMIg8JoDucDQdVISM6k/VmimGsy3Hv/Y54tsyBqHQXI1aZpIPZw4iKzSR
jsrvYj9d6w0F3DJ5Q7voMoQn0wbQo3c4fvGSISar9TnldSJlu8XMwDDw6juNjMkv
9lftTGrphDkNFJjR/VcfR3XgLGcuqG4jBpcJrW68uuJM+UnSNaCSBvdfb0VhHnaD
EA1q5kzZRpWlGOyu5S9QUsSYr7yl2rAGcYCv3bHzR5bndsgvJI0QW393GThMwusQ
FLeMgu3n1duhRd6ymC9HO3k6Pg0SPutr6Cva/HWQBrmSHs0Be1O57srz/w2QZUxa
n3/m0gqDp2QzFYFjCT/ORSufG/7hM7Eqctxz+1ltIKoxe2+i/SwmVwyOdCLDW0Zw
GPyr9uoQlkalvTuDjPeueroorbP77PKg41WDvkLnsc9nqpDXwIrhiMvpDNiqR6vy
+1mD/Rc9bK5tnDJzo3DRT0ALTzF3XQgPyB1y60xnZVkcDIbsSKNz0alga9Dqcn55
P6vwf9+/o+l6+oKiFMNObtvfNy9EGQBh3IpTXKu9CCteZ8jueGbaK4G73A9wgLlg
H64tS+3jDPIWyKqRCcaZJeLDKD1hcZFaYQk2U7ZoFg1g/LbManTNxcvz2gj7ml8R
+QerZZSbf/9r/EjvFFuAPq7ABBm84y/up19O+gCSq2waxwRg5sTVeFDoIdKb6Adc
UIugNTdERqxLlwCCLsDKGA+3O+nc+DYPYhZF4vU+Yoknsg6YSBPD9hZUVbsRrX/7
eyKgHD30zygNwLUGHcGJVJy7WzSl+sb9RUizlHMc6Y3dn8a3AiPfj3Yq4Jgwcs1b
P8mTQFbKN+pZDDw4EPJi3lfygUYk9577VD7QUB/J+Hd0GxtAPbRmhmSoh3Xd+E19
bP4BNZqIGD0uDnW2PTO9cwxCfKzbhRHQn5l5xPd3fv3TAYNiexvWnU2WLc599xUe
UHb+MBdIoYSd5/BiDPuLgwhvwJJVune0UVwmXzi0sdCnLNk2Qdhw+vrTd/zuBWYg
OV3gKK3eLZGn+Q3mZGdFag5RFF166jweoOXy+yQX0A9FqPdXivvnHoZMBU6hd1sT
z7c4AD15GIWsMdvJgfXOGm6oMpBZ2vZe0mFm6ZOGi9RirlTnLMqEzoNqDbOMmFt6
x0jzimAZ0v25wnGyT//sb7qxC2r5BcoPkti/dxT9XZWKBDJ5ivhLTLgHJgyjceKg
Oggt3T78/XayXHKJ/qMjAq+frtvm2CtU3Fq6dziJhsECg0yzc2Vj1sTr7whIQZKf
7ad5EnNoT/+mXyqdAma28y5+zEk0yMTBRunO8N/LIIMwC+lAaqgSOBp/nG+fJK3g
LlmcW4QMc2jkICY40GcqZG7+B9dIbSwFWPhgF6cWwwSmfzH1B+8JnBLsxxbN6DSj
OBeC1MgUw65GhqN3Cuz5NNAUMDkXEKwQNcN5L1j7G+g8s3GXLXOjvfBDe2JYVdnD
VrFEB274WJqVG+p3dAfgh0Yx++jgoxH7AhJU4r41zep0Tk0RQJdhtbkMGfmcQvgP
ny6NUk1FC3MFE7MsP8yFCBPRknzz0pon23x98PAsgtvLrXG9vnIkrfg5KGTVA4dp
26/NNLMhjAdoJ4aK+uPFErgzhjYXufhN2UMQifWpw6MGl9SJXz0Yba1/53iatCtv
ijb8sQyzEqKnWj6cpV0bV3IZI/Q9bJWvNyqdTfu39ailSNTc+fAJN3f9IT9SGa22
uO1GdNhgW1Oo+LxGZYNZeIIBm0gulEM/ZNI9rsQYP/5RjbE/7xvi2TcuWF78V3tm
J+nu1RBOX2JDLAWb2EiO0FyPGjn3tLYGH52b9BOrbs45+p/Uj3HivbTP78t2luGZ
Pb90vtQ84k1Nt/col8nnkBJuo2vD32NmkeVvsIBdRJmhChHysDk3A+ng1LyRYPhc
qrLCapYT68tBM/XSQrZJh6EoEtwWM5ijQnMu+p1l4fX3mps8C+GQCjURyEwHYe7I
zc1hy6AbhLPbTPUBiE/krcItPhsg78FsGWhyDB8NFGDtqpu1HVM/LFjC0UV0SQ8R
73Bwpna/L4MuO6N4c3SrUKUd7zHoL68lHRYRCtOdU/Q7B8HcTmKty78lnH89qDnB
bNlwgzyAhBeWjT6QSZQmCBdDBPwB8A0lO2jkHN2XfuOi2pTPwECXooSp/5zmOy/P
oB/4UGlb+cSnqw68WPtN2oeLrZ/GORIFPvIc5hz64IpWhP90A+3+LaKZXCUAgoxV
KoFq0lZQ5mVNOpDL2jSwsTuXyBn/syJQ4iDBL/eq6pQv9ipAbwqwLMUUA3bnV0qN
soHSAPEWCSAlXxo5fclE4xS66+xT5oyK1IiC+XrGunbuX6uDcDGKs1PC/EGGDIX+
RUq2ZF4NLrTmdA8XOASnG+xMX+FHOt9gFXM8X2YLJmrpF6pwKt5Dwgue28dytiKI
CyRnnKaSMHSCSdhEDSd4C5CHPzKIdW+muMJx4uEKsM/uXe2bNCpUNpK4npzU6s7r
4rHF/pyr6ZrgufShDzqtdcqWjgtGZn0aaxE/aYHc+rf5TW03DcEoiaKbUcnMJvGa
LdNyeY7Smb1PHjKMPr9bbeGVLl6ik0KAW+eIGB0tKl0B4Xcndd/XEsVxGvQOK+xj
0/IpEdwa6FAoijY3TqT2PnYaG7wdrqf7ftS8xsWpyb8M6+UnZgv10el8b48eZ0lg
27IR2XuwCdgkvNNnqdQJOt7k8VvgKU9l0UUWCDCBCxrhGnH3Y+Zfun5zVHbbDJz9
qSwzjYxV35LSFAG3tQflJzFQz3XzRynSc7PLDwT5xdKz9Y/I0/P3/ax/DK8ufzcn
+P1eg/U92QrpoDIChG5eqYPBEJbRXTDHl420JR0gOh1fPlZPYX0pwrAuYSpiQ+XH
/axiaJrjbVW0sKTVhTvRRXTKwNmjhU17gFUZSzFjrMfsfkdtG3R3wQilSzvZaYXM
b45XIUhM90WJ3R8/fS5zzXRXQmGg6h5oLeotLjDMdxKIQUc+AjLjNBsANuCbal1A
dJzf6CCEzAsfZqo0DLRmjvpIQ2TvHapZkcGGzO8LVU7scjZfYQFsdn7k2BE0uMB9
TdwE0VSC0FQWqX7OJhuWV/iMQwTMTnNjanfAuqCbwHl895IcnPoBvulZLAaMPs10
Nri1brVLw6NHuumb7iAnNR9jWKfurfbGY/1LWVEOTJI5X6lY7hS0OMeDWVAXOlcl
XBilrVfKPkSiT3RaZ3z0Bes2DdV6Ru/up7qpKoypFO0HbonxEpTMP/1MEEGlMmoA
WDCdAMpyapmLvhzGfRE1fGqZ44lLYWCP45Hcrx7JOCa1Z8xHFjo0OdYSAzIAM8NC
zAuoe1T2pLjjsVhPlrT8YMQVpTR61iMZOyYPqMM4DRqX1Rs6AJcEIPg5rSU+ojVv
ImKhlae181kaFEdNEdJWn1ESgjL15zi7QvAM8FrpwSTjAhFtBo49oVeuzg91AO/J
TCSyCsMMufa4ZJvUsJsmieDuavhFJThLBANVQTwSlnouTgpEqiTXZ+yei/v0DYTg
IuuU+pWoXFwoL1lPCesS8WhIKUfsi585XK6fAGDsag5gTmlFYmh1OpqLSQi9jFCL
s4KO7Ab6faHOUio+pH0SJXHrcacNQoUJU6cqB+flRLubTSxV1APkPhdqwtHa96w4
TkPQHK1iE/Gc/4voc3AIpEjMEsSrkZTb9U6LPeDP/pBt4ddlZk50khFOxLDCaE84
eflSdeVLFtv22+sAMtlynOhzbfHo5//xd2Ehhqc6nByMbmpc58Y6+muBQPmI4zG6
rfFXfsllRJtjoJPU6/McQfevd+gtnfdn089Nmq6d6ZrGMObKsKJxxjisgV544IxT
UCNR+XYtDTNP6wQAsKAEPd5HjSbzFoEAqo65BRtsMIhLRpV8gpcWZY2vcv7roWPH
h1wF5pDgHySv9gCGPoPie2YxmYQiZiogmxvS+Z4fLR+gt1uTkuU9EWCEiBKmPWPy
zdVO5FuWFwHex+4TFajQNgfnlsZ7hrW/zUJGzGTLlvelyT3PFQ0APNEDXeEDAJZg
rGfYDc6DkroUJn8i8LgaC5aDzAQGivW+W4+rQiATe1OEj1LrEpsqKwUW3C8yhJ/0
yyMADGpyKyY+e0hbYFekpiPO+kifDwnW5JaNHmPQQ6tK2WePzlkGaU27VI2i/4E3
lMy78JTBT5jfENg1cOZKPNtOOExdl6/nobjj86ndje/pEhGuVlwW6NPTybFtMWmo
+BY7BHKUpSHRJ2UDcd2uyKKaiWmM2KsSJf3yhqZ2gPuLhVpvO5Y/OfSMEfzwcSZ9
+J77iO4wcllP02uMU+4lf9wsy4tIncJ0RXE9Ypg4hbnCSM7RZEAs5AbV/CE4x/wX
2ObVEc8jbxvFFONYhFx4sI49YJCfDq8V67uZb24W3SLPyKA7FSB44iNIIKDdXRV3
LxAsFWcbzAHEjGIonaEzQcpb4lNvB8Brf7za2Au7uvlJuvGUTBw8KBnmRUEgckEP
2Fz93WCfrEOVReWEClkY7NTDngI36uBb/rA9pqeKxAFD6S6sAzTFlBSDl5hJv4lS
SOvh5kSB+xEDUwQfpB40pvr0MyXU3yJKb97r96L7J0jQZdaQK3vAIhOvh7YwMJdd
6dhhDkc1jMVYzjbrGhKcKY67B4eIf3hxPA5Q6UXstH7A0Pr5lwvU8oaDqtbjC9ef
LYiKYbk1sQhia35d7birwU7UIkS5IOIVXNliMs5nlsgsQ/6xMBH6jYi1vOOwZl0y
DH1SipYQKyEMZFTxvMgAYmFHPb3UI+/Swg5Mxyu2gumSMw7YWcwEh8940mZmpSOC
7Dz7nLrsy1F0k4ZrQ/KVxv3tA+N8q+HHF4qqRA4SBKvgaT8gsmeqlfJe2fU6O624
Mk/OjWT4IxS3u0VnGPH6uMzDXt9AEVmIkl8Sn8+9VJzg0WpBZu22FzENrYLCOnIQ
4+5b7tiSuYQOvgHx+ki7yghJlMZaWSfcYD3cPdvnR4BCRmwFYVd9Bpn8G9X8sRHa
DwJYFlsoAdlPWupSxynf2veqmI/vihKF5DoMYo1F/XoF06ns+3zCvAM7V489agwd
oIbCiadMj3Qp73Oj2UB3n+5zRWfFSxmLbQ40OKLGEomBdpXATrXGsryVGxtkaeL1
G0D2nxaCIJbmsa8jOITLu2pxzBAZduKT0DKcqsJlPddNaO9N4zrLKvLZr3gs3a19
eY62vSXLIA0I1e2eetVmZjY7Oxe1Sb13VBv/s0P6PfwbNidah1v7dAekW3x69wu3
AHBNCToA9g/jhJjXaJ3GmI0vhh1ba+Nqc5zC2afq4d96BDHl0Qh1gnpurwl6F297
GGAxhoPT5+bjJ+Ta2Jt4QHI4CJteRKVSjGDXpUcofvkZB2cHqS9SdIaCjdCdgRN2
1BWz7rKJLMSUxnEJCFr6YsVU6M5AxzzKwC9Wv6Nb5ANJ565C8DixGV+Rg4N8+tma
PRSgNfut6O5f8nB3SmVRQoXYPytm5s77VsT9Z8w4vAHLVIE+PH9a4hTzUF+v/iJp
GdDXRuVCsGoP1UYLtuvpNx9uvmD5e9qDcHoFDY5GJ2sx0eX3l7gm/ccwBceDaeKF
8reZvudsyJOpzJWMxs9v1JYg9scirW7lXjiDTiI8War2n0g16Uouiguu9Iij7sJp
yNWyAfuF52lOIqZkL+f0aS47pbQDskE/P/BakGaNJs/jZ6Ej3mh4De6GRHpjgP5x
AtHEIQHZG3BOx1aiw1Ij/CIIeHKp6j9BOXYHFezU0TSPKuOPZeTIijLforYpbtkN
VoswCXiYrryT1NOmEFp7ZrZGuje6YLXjbjQSyDzexxI47+WyPsCxFhC+hrvOeOzE
7Bfkh+2ksr19lvquVx2wyzqq7RIFJm4+2l8wcSCQha8ncS5O9O0GgQaweZTJCQJb
8yd4/7ciTLddgah+i6kez8c9XQUaR6JWCfeLPrOWHGgo+5JhdqVaDAKqotQBJ1jO
/KWoFKDFnOSGWGyiM06uwWZxCLU2xZqakINXlDtbeSivImmVxGESy+QlY4EnMsI9
r5r6X9YDDH4Wmjd0ngP4XaB0F2lTYdSyq+mXh8FcFaE+wVuaYqbuarV55VSRwmO9
vii2OMe8hnY6YdOjnDt85yWNevJU8pgRGneyrbEmn16I170SbsCsLXh7CVpuM0CO
5qSqOOxO74uME9f6gMJu3YtbhVGN4cem2dl5AYUwd3W4WaZtxVUexAjl4OPiMcpg
Ry3L85eOjt8gHJP5zR2JLe/SE/w9d19B2zn+wLI1NLtagms2JRHtPgLMwZGHLnOg
i9wLjzmUQXspZG7uoj/7RO26SOW5X/dV0WyrLx1vt7R6cQa4ROIAV0+oF0yPD4CK
nrXj27hyEptd+BBK1SrWYFsLF8fGbVhrMTC0ykbJUPy8CypcieNaYej2tM7fGFvd
3PlK/ufG6i3e6H5QzqGYfmY+cL72CEK2CJCZeowzPHpTYhvCjvAu18Lq4Kquuh3m
ODsj8LEgZjzRkwAbvAEDkxDrrICTR8MragJgZn8GzzQfrXKpx3KTyf/RbW+9RNOH
sSnHiG2JKvHY1m60NJTR9YZE5JkfDhSfqj7wXu7jg6VSs7T3y4G9Pywgm3if9iZw
1yNo9d/aCuoSMRgX8cgrJf5EUcQvFaBskhBmmCksTdyqc8kc06hUa+7v6IgqGWFm
tjDRpOG0E+n+sMFh3HPfXbIcrI4uvS0jWn9dTbCHH6EcSJ/RzdfCmVFS26yfgR6i
B0xBFkBMymS+tRmZ9NJkC6umJT6Exh16sZEQxuvHeqjRnxHYiLTArJiwlwaLAD2h
oc6Z2yAziIxSoFNZw8OOrhatWfe/+Qex/OTwDhiz87iz1zBL2Qm8QPHevZU1x15Q
FnV3PLHAXgIKIKUgnp7YypitQ2TRIv17qHqVtUoGKED51R7JIYbpSjD/ou7K43mF
3zTL+CPSrffyn7xReS7Vo3l5a/FR04g+3wJFdNVBjDsbVFsN+WQ8p6U7QctScfuf
3JJgz2GdiIQEeU74mpotMxdUCHIaV1n99PnilKi2/yZTUCOir+A6QNQo8yIuR9ki
mVBWMrqYhVY8vScCf8zVNCDYHqhCh8ezsZQgMSaEoBWphKL/IRADM4DQqhPYEy7G
oGUS3Ga8mBzK46HLcXqUqEbYh7J5xsMe+kfncPRnYBejCxCgRow0JeuQ59aZMHd2
+CiqZTfBAmU4om9yEzc7+v8EEYW8RlHAjXFbYxY5o6C3u5hKGaaWuVpl+PlI3eJt
Qn0TAWVSls3GDz7ZDZVzpqFOse6fDt4/qM2rJmrEfshGa3kD5Pi+zKKXFWXdFSrj
5tbfPzo6AC4pAdYv4Etq61iwKIwlAzatVNqY9X5fLnrBJYPK6yqHVCnu2e7tKt2y
W68AK2feNbuZRIxiIQ4zEfsw+0oaY2lKl7rCXFMQ077lHDWPoaek7fzjNe3p7hiB
QgCMdqoyZUo+WP+0Hw33/TTghffWWUvwgKtlxYRkAXpS4qMyFfQRcOIcUpNzODZb
oyLdvrV/pOuFpKTokOVGH29iu4RphipE3Xa1Qz2438IbDJPl97ci6+V3S9TKciX5
cc30BpGrchDMuRLoox8NqJMbv6nCCBke/Vbwc/EyQ9AQ/wDhA6CKSAZtkFn7Fc/k
e9oiMsR1m5Ra8tERK2bxPQPRNSdSB7pI+jL3+BiueW2GwuROIf590EWOd2Qc/9T5
tcqZgkTVslOThPczpUjRdWCMKNhiApDW/ndXO+AQFZOX8Y+z/wLFUH8I45gdWVh0
p2GAQfy0NnhuBbSrEdcG66VzzW8mcW6HnxBWXmI+z7IQs94zrDuQNzaYvQ51ReND
542MhOagQRbkzGXU8kmEMU/rQZZnGU+X95FYoOVkXMWB3uOqOLhdSrDUOlhBiDXo
KM4m4LrCGg73dNSirsad7yLHFieZ/4I/qRUMPLuH2cMwvphvQoSJAbRpXb8ttOcW
uITO1C5HleIc01cxpjroNRQ0qSRoKYbpA/M2NVyqWqkkzyTPhzi3gWjsIVscfA1+
6sLKAlgyOboU/fI5B0xM4mxHmtoNsEgkCr71P8eku1++Ufkh4b14kFFjejEGolwz
4b7Yuie5fMaYxg9Y1+YVXluibPSk3YbaSSYrivvt6IGi1ApM3mH+GzeupBl7NfPs
jvv2YU3PTn+/KyGSV8wudlADMBuejAGdjuZstsxK6uY2RQU972UmV6hTIoN67arP
ZLRXfZNb2Tg+ukQcHi7Xl9VS/lDI4rv0FFN1k2yTamZU8BCxRkPxoy17zf7DpB0W
kL+1i4JG8NaeVvOZBEIhRCUax7ZxJFV9cniC8UFCxrev4byy9+7iY1DbjxBFV3t8
qjUc/7D+NS4nUAmNumVag+vhqG1xsWI+P0jtO98COTdS2U2Ww0ZyfOQE2AWKb80q
odoVyRbIOjs67Zgv5pPpfPcz+IGsCMKEsfu+wlrMT5Wk6XgomrHG6zr+ZpXwGpMm
ovGKaiNuRFq9uZXyOCayIsHKNt3nwXo63s4xGngFPxwBVEPTz1nOCGHpP664fEC5
jwAyvUk37AT54OeR4QB1Dx8grkKVTz80zUy2JmIwRyyl1v4y6zPVkNpJ7xx9YgG6
1spXxo+7fQgR71xf0AwyaCPIlhX0vrJp4pV1j1RVW/j3rz4xy6wbWxg9UFTY1fCz
66SNbfEiVfxGjAL+0Llr3kcvXA9A7ycpecOhH2K4mIgHxN68cDa8AgUqZd6IZQaL
J9KnqNkYAAeLiDzaJOzWBHSDwXtCkRZBSqTYGMnVU8GudBOi2yAIEViwIZS08C36
BgLJbFlHdLISsflMgLcuKyKs4XtSXuVVjmRkqoq6vQ9IrjFVzbhKNdCJ2Xah1PgT
NxOBzrD8DbjXF/+wTqt1GBGT37uGutEO4e0oLMcWIFeBTnVwFUb4lEkfkt3nuVNv
x4EWE4gScSbhlf+x8gdhIidwBzsXM+japkdFZRXj5bCyARxaF5hnXvtO8D6amv2x
syi7cYMPhsltCQ/8NcTt3WAnclcpxWun7PH0gdAkslIkpg+Ny9jJf/uN4sq4AKFp
AWDhe5b9M7asflabEvfWSYzisM1iActX0eocQ/O3+PmB3Qk5t8dQzan5tRj07Ipe
LuOf3fJtHsS5Bry6tIgFpgaVsqCg4Y28RWASreSdiL9k879Uk/Iu3dtX91Nx/fsb
8gK+BI0KT2QgOFYj7l2dkr0x2eAYO4xsDjZP2yYUxb8yOoFJlomxILQZhrFeSkp5
7YX2hqapOemy/ZaiqnEtcWGjZsanetlDrEBAGp/ImmLKiXkAjTwD+y/ZxwePE+Ij
DM7VXK5fd55zzxqeR3c9ckxgVREW6/b17iD770c3s4ddTzp60NnicuXvxysURfr4
ju/frZVTBqys2ttS0pd4Yp6MSaMAyPNpr3U7XglrK/dWQhga7/gSSW7QHzSYLzS0
kgY22G6f1T/dA7z1B5l7JArCjrmkutTfszsmi9otgTnFWLpLyNCjV2yrzlVD90ej
lXlBnPpNgYlF0lzYsrv/CgdjEycSdWFeMwv/ViD/2qF1nx23o57zszjeaMK3Ykvg
OFl+YdDqSgAHbX9S23IPqju74+52fmq3lLE+qExMX/9snf6X4zj7zQ5kww6IekhL
EPevdIMVwD1J+6yAshlveUm23BnRoyED4No3Y4d9rieXDTAYpFJfEvLuid6HvnUx
CZwpbdNhqSXrsVgRhM2Rsx/NXbctPEAKA8uddWrWmqxXgxOojWidcjKbvkGfHckN
suVREd07KjbHntN+cMPWX+3MfXnHRZzT+irr5lve3esNHRNdxbKIWPyVy8p/C4LD
R7JWSISjIE2aBx9LF58LlfAbLXOZ3Bgyez+rK0q1REnor48BmhUKMjfjm4L/GcFD
629t1XpmnIzISZuBoDRETBVjQWWXFewpFSZDMz1rE7Moz7FtyUYGV3R6yfcLYA56
WtIsn2IejYg1ZdT+bE9pj9OwDf5euKYm34DWnx3bRmBe6j844U4rYZ61pA5biBAB
ER09xqklIF1Vvh44ndvGrW9pwPvTNuSHOOabsgybXVnIe5j5guVp6XLlhVaifMNj
0oxTo5uY5gYaGGvu3M/Shz8kyBHDSplzrvATBWdCJHhVPJuoU5p/HNMejkiCeF3S
A8tf7CoyAYunzQJIVnbbDC6Yjrhl1Z2KUhfKd9dZpOD4GPLiyEbIAb1B0MzwnXgO
5hw/7hNPmF8MHRdCwcYS+9Gh//7dhxOVtSIhdfj4C44GhfctMP6SUHxqCr0DKiSK
2Tjxl+NaxFF0/TfAOiu7y4Kq9GJKOVeiRFLZOtsi0p8rWU9HnqdmwiPDewGH6Il4
Pua9hzhfZJkdgAxmoJgW/9xlKK+Z9fr54YxfiOfBT54pm7jfLn/mIVwnXneRAt4u
63p9cr8x/HktInayTXLb+i84JkIfV4WeIFUXdi+2R/HpC6Q2yOeuHbm8/CTqiUDi
wvIaX41nQ5PYWSkWpJpJqj6gZH0xlvl1LtWZZ0Lw/n4PeIs0iNzGeG+cIW+y4HrF
CcwhmZFRKos+rbMIjUhyZG+e38V9W3osazEaC1F6jLe5aJwQcmjYYLhnJiNYytFn
SdNGuGWghW9QQrsfONMcvzKhf8ya27ECnm9mYjXUt0yiLzGVE1FMyEUkSOn8HDDw
qhQpfl/tRKOuBE1q7Uz4YMs00nakn0H3d4iIS0PUXF4d/VuJt231CAvEkDzqV/hA
nhpqLICLkwjxnGciO5NZ0QL3jH6u4sQWb+S06mW3iaBgHETjd0nJu6vsfqqaUkpt
9ijC7ObO584c2su4RnyaUq5vgwO8kJXe9I5145XYT+OXawwaJRS/Gf/kskqSQPtX
Y0dIDeL9d+pbrnbKamd+CmMHN0AkdJLNjk433CbzdKE2rU0MqSE5TWPSSO4YuTgu
eUd3XiW++rQkogfZn9GBvipGXX7az4jvmyvpuMhqS3+vjHckx3QidYPmlEF3F6Zo
Z97c49Fdd8h7KgYGCvCmUZKvyiBs36pUanIWDa/FCJDqm3mCn8XXtA5WoPp232s3
WXCiia+0QnNFiM3dJfGtV2yirNwqxqLRn1Y9Z6mX5PVlqdzFWOS7gK/3sw9UiEoJ
fla9w+W/FE2nbgGAwqexY1DeEQTnSW9jr9Yjxn0DqnLMgFkLQlWoK9tAT+kOyC0A
ZGnaYtUH01ARY1dqmavbGKkfAdSDCNzfcLt3ZcsX1HvC6DbDB/sERttWlDjSRkBn
kc7Rxz9k5D1FHSXr+42l5+nYIlIGVemfNSjNyPVRWMtttj4RmVpp8VX0i008CHdq
cwsgMAQ7KdBwr3b+HEYSduBlDptcJ5/8kNlA0Zz54tl1z6DRWfFFudcc00LYY9Vc
QeQYjgg7fb5IMVqGgF+F5vDdcOcaRFvqzGrTG1+NOFKoZVxBUVEZOeugl9+CvmUL
0OyPDymRSeZdYxnej6A6JPjtGJLFl6wfyQwU8PrnlJiKSkFhQUVgVkNXNKpEqVru
ZF28C+9kxz7CKG1WaVSuEY0y8l+7RKpOwPTAKN3HIU126UtRF1hMcZur4KpxxV14
sp1lNKwH3G6jCnhJG+grql0LM940kAm3XX/jpTn8CE0G3uGvHjhAc0UYhZICw+By
xSCXEL3i4WJvkKOClvRxmtvV2ST7pc0oK2dSdzpXnNYDIkpJFcuJ/Ay0hKqj2TpT
+X8hvSQuAyrM05o+qE3wmN0FRka6WKgZCIeVTasWEu6L0sbEKHJbvBHaeyeTvHGt
lRTU0ljjwNKUormY4NNMpIAmwFQyxshJGnnfLx4t/xJ3fNucaqYeozLcRz8nFRMm
Nb+cvL0yiBOctaTyEgMoNxCETi3Dbr0/PqpIgQEiwLUpS1wi+sO61m4TKGSt8Utv
GCUggIiLzv8cToygkRFg4psfAe1ooaPJ+JS78v+UYzQT5dsqkfrgsYPdGwC8c5LT
TJk29bQDphdqkdAmmTWMiRY/eC0GTHSGjhaS9bHM8M8QGvolbOOsv6AO7ORZcoro
IrI/tFDNwCQ2wsQjjS0724OLPEqZ6slZdPzWEcR+HHLmbIuTvhi+oqDHr5knAZbR
c0kpb8AMOeO524t+gOdETirBAxRTuC1hJT44+WVdr82kwi1M8oRPQfAfRp/3A4r9
jLo1KB4UU01aBDbSyTVO/RNm++fvDXfS/wYdhzGo2PvfyektPLCvJqA+oX+n/oG2
V7zFk01wqadMj+yZQv617qRIgPtCnNMgTrOOB6Es5gna9QZxVyvGH1XoADQQOcdS
XMQSYLgPdtTTTEHUNmWnleFl6dSsoK90md1itGWocdFpbUc9WsioJLdoDI3oLiY5
NAaPC1x3ah9DJqiTYERtFH1vBklBM+ftyU/Gesbb4gN5+wq96KzbMiTMKKMDXiUx
VUlZ0OLtFKrW4KdGi8qvlfYcIfoAeVN6/o0Wtq0TleUO8e1xT/BDGz3kcJzgju0z
iZgtvVXHqh00Q26RZQ4yPWGA/x9cbf46GPE5cb35inSpaW5rMggwCr7MU4NQNvs7
lZqUcWndhg0gUW+VCmi78XyggXS9b4kBDHLxRxAFW3CtF7mYntdO2m7oBG0yD3BU
vs532bjtcmbuGYDKzJ0VWx+sFMtYDs4ZFCLJ/o44KQa5AzG34x/GMRwRKMspeQWF
kj2Zr6pRZHmrqymutGdMdOYUSu5IZaYq+TdN3jnMvnycZu+369Kv8sYInzp1rNxX
9+g8bMDcNAFcEiZ+lwo9jfZSjZKbD/tzgca5mipYJWndX6aeR/SJiv/nFS0yDVUK
9GFH5Cue+/cs+rs1g9/R8PmV6Jot7yav6Ackhdm0FZ3zfF2hqbO8DbMfaAJ3PJgO
P7vV4KPdq8noTptOicU7Qp9T/PRhHpClOwt9M5R6BZSjQDnmSn/PO3fPFS0s3Lpy
Dys9kFgRYb4WufyR03Wc6PMMIskZFiTqRrKgfP3+ZYCHAhyb9KVKP1CM9NZHBSY7
mZYG6cjo0SF27K4hovjJ5n4WhRJ40Kn46vzm5M1gtpv+YIaAekeXN29DhKudex2M
ZXOmcQcqg8YpScqoHPvD+G1x1ORuYMdxI6qEH0i2cd/32SVhSMdOP9TsURsxmpjZ
AdW781d2LdRlkXX3Kq6IShZq+w29G5w2DGQwVV/FS6SB5kuTGcRTwyZTY4qWBond
8g4KhDkjOHnHXjZm/FT82/Xvkpg8L0YiMQggr8lL+0F4/EEnAB+dtarpHdjZMUTd
YTWWQ8rmO9pwoGmUtkduraNp6Gs4wj/g847KiTzYqap08YFK1H62Sm4Dk+/R3lGk
ctKlUMvHKNWKrZnOc44Wczea5z15VLfDQbKjH3rEwVky0/A+YEK47Eg+whTNsJly
oZ96OODE9HuSGAj7rLQSvDPKpIDW/q3DAGP9Q+3PE/nZfGx9BMUrUB+SWiRimYVy
Woman8OGowx7fnISrBBJhAwDIsInh7An8BrHW3b4WwtA5P8hSR1oXxHrBY9Nfh3Z
9AYk+Nipt8MaW0Oj7rQapWBSq3W2z5roW8p+TMh79FmJi5tC/hBdyWN4SvZgHboy
+KIGPzR4ye3rw25Otcya5sll7K97tKdIf0Ns5uAzCUPvREX+jvDIVPFPXNKZ90b3
3tUs/EbeMvr0M3nrH8OhkEgEHs7OTmo9W7cPIrA/xgoyd0Bk9Izqch1RO3nd1mxZ
WP82yPtMOmcTNJ1KnhUysRiAxnT1E5w3/1iOgQgC/8JvlNIb9OhX3x85i+N39KrW
hw5pAfgHKKCKAQWbAxGs4ohp1JMrzNW87zN6Y5SZdRwSwcE/34TA0yy3uYtYqMe8
V93DSv4qZDxekkkCWmBCawQxhap5tNS+zFpR2qae9pC7PD7ad/K0Qh0NMjcD1XI8
n0WcYBqMvxHgttGbVE1mJM5+CF/KAlRS24ixR20NvAq19DOzOl1QjqDWhp/9TeVf
3gCRVv5293l/TyzInLndQZQ2jAKCDrHO/qk98ZS/z3Wks6RgF5erPialazpoqvSi
CiOUHJmLKJLafsC0ar4jh3d/cQvLFZSHxlwecn2bL7ygRE1f5YxS6Y5UN0aRi42C
W1BDiiB9j4yMKfa35oA99QMviBg2K+x8zSCe5akYqEwki3FpVItgJLHZKfAnIa03
MfiVbGeocDRn5rbWOL7xlr1uh8PG3Wrx6tmKiTz9DM1t4t2ujGl/7yFivxdanPHq
mP88XBcNOvfzwyZYydrgENKGTRMCskjXLgKSvPgm4AYhwIHiPBFtjbSUKmJV7N9+
Rw1YcEnlm1Q5u9lEWaAWwHMCwP+OXjg8FVsNQHAD2+K3a1Qga8y+D5XBS7aEVfPH
8PQr5Uqhd/rHouOcNpQnLwUA8irHHPAaPw1X/O2iwi5hsjkTznwOSFylW31AGf1W
m2UhhvJK5VePj4IxHMptmSFbvOI4Lzdxbw+0rYNK6RnHByGrQIlmHkWyu0cKgeS1
GGyTifNF7K735ITzata/M/qK10Dgfuwk9ds4P99mamCY/432zKG5ZnfBwJtiVT+g
tmVnHRaPthKEx+xVghsXtOzdn7Zfcjyx6w4dE0AkuQXwqa07TTYntqIThk/MChWM
TRgQWGojABdw+AR/3vHJAq0zG9LOV9QuFtmd713In5Ramr7CRWWlBOLcSQkg31YJ
dRiBthTx4muq7Q7XgxLMr0zsdbMWLFz0eZEUIAAAPCRDCYGF3WCyGbB+mWPjXD3i
s9ZX86z/a+sXwbsGI6AHroCgX15SVCKqMhmiHchhI4jhVwK86R4E1r+M6pldoD90
L778NliNvysPKBbuaxGc+9OfCa7WOoJPuAp7Uu67E5D6lqe6xXjNPMPkSH0foETO
kCJro3NhWbn8FJAB9E5lJxSR5Nw2Z0fRC8VS9NsCcCYt88trAkV6qd3CmmG5twKY
g0OY2FhJGWDI6bA/bJtiO20ywd4Qr23a8cDUhYOSsQaCD+Bl8RVg1dUoqNP9mLua
tRDjbAC992+v9ZkcXgOUXIBD+8i+1/UNlSn5aR7PVKVTRxOHXS2zaTySSW1Cri9V
1LEKV6LWufK1khtdyUArC95TrGnsBXT+NKP8NvThOV4Vr2W11Sdqw1S/c3LxOnPo
RrqIpzQMZFny8Kxj4GDxgyRBenvQQodEUEn0rqn6trpYbenXyguVwq3QX3v2tdvG
6kPvF8vlAHRu2Md+RxKgVQ0N4kUrKpKwPsWupgM6C9FjHza3v998awiYuluuEurz
6mRCb0bWoay1EOynjX6PtKTWlKSB9Al778DXVvTm36qgF3xtvUtbhvsL7q7/PmFm
2Z8fMUB18ohAV7K/KsU9bwNwOWvd/i+3IiozEMjgljQfaxz1kNddfjRlfHnfVUTR
eW5ve+/+p6fPve2YaEFS7GwyTepvZTjtXep2SP1q9bQBQXXYsOQ51FPLZX7uQWna
uc+Db/ZbiGIyB70BXcN1yY5u4JYhdu8eKnzajFvuOKhTiCAcAFhpfFtiHTcc8ddj
vtBKLyHm1wzkSjzJhbgnMDhfvNSIpJT3hoUi749OxwQ1MQ4/1K9qSJg050076oDD
65Q/K4Q8Un6fk/aB/5bdaATlctYF3jrrZ7fFCcCkJ7Y3aoWDOeGteWLidQGFNB8W
T8fhz8bL1hwDg4lbH+6cKrfB/UQkxzLyRvWiMd/9619GcnbZSNgBHOz3/NT/dNeT
l3GDum1WaKhVQ4irkvLjjjPO1pvqArBCGv4wlTjmpwFWObX11+ug1JHfRuzuhclX
fIsIaWw2bCYRupGgDVepWbkYeG6N4aAcOD7JaOkap1/h02Xprifp40JgO/lTtd9L
c5qJrtQiJHh9MO867lOnRm6uF4qefEr1Zeg9pYvZn19t0HN5eBOUxhcpujHNKBDo
XeMxL/EwX9+xDaBmD07C5zrSoul8MHI3eBQl0kRGSioThakUVhOkKw7uDowRWGxU
AXXg1RzR3eFiX3E7VCks7U7IrAN24HEP9IdpK/dus/OszzH2pNNgOfvysSh1/SMy
+s2/8f+vZBJK7VHFk4lmRKkEBBbjSekti6/yEJFtZBPKVF1+cJCJ83B+p3m4pJum
cWulvKEaoNXm5wdSa1OiytD4EtL/gMMWfy2wQ6JVMPygJ5grji/6mTPMYCKKdOun
2VEPcA2YVEoQNSOkA7Td120v5e4lQBYoldNT2D/3QCY7dAy1T2o/0a8W7bLtAOiA
8LqOEZJJgUsX6rDbQvlxdRuRZFEOix8GhzGrx5Y3Uw6nA4DAdJWx32ut4z4z90qw
4Gc3Z+xH0FCNl5pGsOkOzLZZGkyglxgwJRNcaCMfeh4Oy31fAf9Qg84eVq3SOFXQ
BR+HEySovaYM/M+5jupXYSNyfLSpszPCYuyxmPo6kD95qvg+OApicTve/rCuyBP3
HJhMR7MozWegoNga0gbAtJh+ADGspdpoTKxQ9D7wBEDtx8CPj1uN6M6i97B+i55M
wSNHXDt36L3XHw4PHRKcy1EMRJctK/+a7bvQEIvzUjwQufEp31Lp4AEk7mpY6Vvr
sA9XdSO8jqoae/c348BIUbyJIzidoIRKqqAYHAgNQonD0VjDaxH4nsomkcWeqFyy
FxOWfAV9+SOk0I9eAhno18c0obr68xSxG07V9dD1q3N9gRaWF8qyyshUi3WxJpYQ
KEpMMnradHTC+lXhHFxOne+56zBwaya1SKcKDTqCwVuG7AZ3kww2+Qg1VrkUg0lb
sASNUv8sKvxxnZ+EhEKGt+y2Q5bS4D5mK2GeFIak5KJSxJibYt+IBemBfOm+hL4x
2TWhancQZt7Dr2eIS9txx7HBzu5xhtT6U7wrZMJ39XVnKQbckjgS14v+sH9lecSN
r/4Bz9FfCd8QrR/3JOkEeb4VKAF2t/r+AramwlaeLvPuhBgYAygUBydpCG/w4mf2
h++Fa/mODW4LYyGvket+yS1EJGgfF+kBQ1WZQLnqNpxMR1MFXL7bC2x6S/L5JILX
nMztcS9Irbc2Us7o7MVNP6hg9PYRRU7VVo6Of93GEzuL/CQr/XvOmbo50Hi7EGNb
7OvLBSbHu4+00Bxi9oHy1Q56wTbgtBkS5AjHWmmUg/st6uJQuMLMaHF2AZiF3mhC
946BP4Ialb1BBZn7TBYUTBd55UK9081rxSVRrSI15UYjsFdhffCLY9GBUHLBJ/t2
CG8/XLL4VcRwp7JzGejAv3nUEUmk+IVIwpIYXmlH9xiJ+4NKapiw0M6lfY0gOZcJ
0uRhQdiWj7KFCgvu4QUx13++nsKNRP8qlOJd1PNyD25mSC27gW5UMNloapuSaQt6
RXC/8FuF+g9ZBMVFgX2ERdxDzBgHxkH/oVhw/D8jZdsSS+fqEkaNZ+ApRdeM7oEx
Iz/X5bEswqPhkoH4I10RKYl3qjqsxZtMxSua05ILGkrhQhZ1kwwrdC+xd5CvkZ2r
2LScMzMUcNVTGe+VsOcAQlG/7GfQFEdtnm41vKitrnWnb44H0wicBy/dqViMhGCW
Mz66gWd/o0iFv9z1VbNb/3ADYagGn6sFpSPnDVmZgKgOU9jpZpdeXx0KkR8Su3UT
udC/slBOoYn6bOqtbUDAmrT0Lb/8WcKKV3wtVeeTm9RiE+DbfkvES5AYaahZiIyM
gUrCFUa691iS3RkqDxFNyHYmnYhhd3dBaEnjMcfQ8a2tlLfB9UTMHVNgRVpK0Ws5
JAdgmOpwly28KIiavXhMLeWMz1+kgcabiAFz6+2LMXHEyuWo3dGGyNhbV9/MN0Aj
+By7kbQi5CyNKk68o3WCBmn6Lrx5ypn0dvrFGtumuhqguHuZK7UmQT5KsgNe1prl
zNiNujzmuDJjBCz52tRFcA+qu1ohUnqHKfoVv49/Y8NRgXC0HeW4XGcWbcwqybVe
b8bKtLCykHnonBf7Tx7rJAoiOU+xnfoX4oHQOOX5RbObCeTcjXhCc6DdJQKaQC5S
7cc8n62j9GOTvhVPquSfcvdEZZUR243JMeW4it+/QyONECl+02dEkDdojbGXgSq3
fN97E4nYui9ISSRooLlWvNqm0UJoSvzWZGMN9tGcG3ZR9EKnPu/9bpNkYerPsd6w
+4TU0Q6EMCR6U9gsT0vr023fFZgy7PQBbGsCmAp6sa9j64BOqfRWgIZ5uNUROzWY
ZTvvbGcQ0kJwlzCCKgxAtVKafOFbzSwLwtQUmKHvnk9auoRGcU2QdOaDL9hxZnwl
Fu7QtBEpJQmqUKqCWuKiNJSFlIvtRsrmhEE7ir9styqw57uzGOqNUsjbnbAjZB4+
6ecsO09W/XGsNi8PkprGQR05kelizFkfJJ3v6gH+JJojEYF78muDBuMttZMIags8
ozegP2TDFiRVR2uH4x8HD8Dgi0avOtGxhA44wdmXdsM8UzH9UiKL/3mYg0aBoIFP
95UGtC0DKn+nj3Ad6zVLJZmyNdepyrDO5eabK5B6FdYP9n9hR8ojWyYBgZz727x+
AGjiVeNM006YFA6z+VfNm3iXauxMGqtfLS3RBZRhD1ErCPHdQzoWnb5au20L+1jr
hUxOrf7+zeRIZTJSl4N0WffpieWD9L2NPOwziGjzJepPFX+gqcCmk4vb8Lsv+u+a
8YCpMcjfmi5clmwhvi+fYu1+ABk8aX3O65nf7vTAgPLbgrG3PSgbHEBkl/ZjNs9Y
BSPLDG717wRDd841qoFOd+l9MDMKslD+4uQhpkgHcahjiMjrExITYJpBUUyNFMxG
fHkNtYQmJmllJmKkH4ASr1fO6Xk51LNP9BaExb0AES12Jia0PDZyoMi5E+lep/1T
wQCnthjuZKA5dQyYQMa2rAEZ9+0zP7F6hZDS3QQtVXh0Ln51ll9KW+3B95hRUiMz
TC8V7tuRoqVV8Yg1sHrBXi+XkuIIaMnUrKG9ZFovxmW0cLSg0Fe4UWBOIpKedG+N
GNJh5UvhS5OoBT4kyaKeK68DnI5nj+gxVL0+mVxfTYp5zAgEGMkQR3MNyKciKv9P
05F17lQxBZLcmBJ8P64WuXlv+rG/WnLfdw8Z2p1CWs2jqGEEOtHNNNar10my8iFy
H9mwwr5oK+TVXUtMJzLGra2naShO/ndYiY4NNChZNCMEKmmaBWTABusE2GwNLIMk
5ytNFvD4uAQprSEwGDKiWDizm6ikME+aJIfPFqDuyiFoW1lLnXpEqK4N6lUEGn7y
8rd3/Rq+kQqh8LNVZmNJf/UXEBE33+HGV7YDMJvGzvdPwnKYfiSc40HB3emkdEqM
KFQ+JA6JprcI+M3LkWdFS6SxIqrzYeUhFIqvSpH2PbCz+XWnUa0yhbpsOLWoCtBA
BqzbDTcuJ7OY8lnudvMHmQGHZistKhJGLXnpX7GEV4F06wUnW13X6bRxUMRKTkMZ
SKQeN3qKXKVz0+geoGwdul56lxEoprZawnyCTYnduydevsl/em23GEBmioaeVxRb
GrJ/xraaHsomFl9XwCkZpfm2ivWSYGjUv3sceywx64mtnfTiJoDF/Rwif66+cibu
f8dMfJ077tGN36RjOkL6Kmwqg53BX+qCUkZxktimueu7uGUCj/4kWoxh10WpUDSK
Fhy1punXOlVCemMRGpHQLuiBvE5E1CCrFyY0Km86QTMxzqWP7s+KWS0ExpQHnWBI
CawGGceJ087talKLiYZfvhXAaNLpeI5LGa0OBn9vzOQKSqhyLIWj5+NT2k74lVht
w7otNfRf0XnuU3Ge479bOgXN2VMlnxMEEjiP0WbFmbEvhmW4dWUbVZ9FZlSwpKlS
BwlC4t1i+9n5TP7MhSjPu1mn+9MljFhdfXk5AhcwXfQM+xPezABfJc94rkfIatcI
HCvFVD8A0HzJJb/pBYrhb2MwxtzE0I75hyMXZitfbOD6QT/WSxsiQ65zYvhDMZkU
sCJOc7lTWipodRcWzGzkcPNsvxNXmUYHwtL1m5hvSLfpoUOXcIyPbgcSKEfwfpJb
yuOA5wlO9EY/Ti3zRRTqNrmaudc5R4oZzX0Pg0hUZ1xbHrq3jgN6NpbWFtnIRlaQ
mMWPyNa3kydEWUDiiAe33rNgpTgACq66ZS1aVv3sqXpVz2PaC8fNQ4SjNP6W+t8J
6BiPVlbF+ELbWZal1Cm6Tw7JgW1l/re1Knvg0HgOdkLdZmFKYgw+WsqMEkcdAeC7
C/h+8s5PLDWsCm0rWTZGiAWHg8AG+kez3eiueyOHj0Hmr3iSXvalLoeVd4mLKW4V
LEybsSZ3x61giuo9bdMZMuK1v8HMEaGlwnN9nSTkPNy532HxGfrAlsviIz6DpVxJ
LObPgDjXWlBmrDOaJ+DvIO9KFn3jJdJ7ZSFQsnZq7Ki1Wg9OGZZxvKeQ79ovrInB
n9h9Jm97P4jEtKY0zbQZwt2/JdKClgD9F8hHFxZDlPv3+S6oCOt8/ssc64JxSTeH
ilOudcoaqip794g1JtVTeUeyDn12xgKhUeZU4apyRouTkTMTA2dZlOZqbhj4cxb3
HTPLkKlWlmrMQwgfda6YZInGoXd5nTgTWrHyinwPUKVhNEjAULYFZGqRSoNIxg+Y
jMW5fQhAMdeuCY96+8DNtI4d/g7e8Gw1GF4PEY6Lv225I7GXs2KGdS7E2aUZEpwz
+eEMgy7D1q/Egmn1kqXB+otLCBG2OF2aWASt/inPkR6yFD90zd1J6pOw5ncYlTqp
957D+92TogN9FXG23QZUxRO51PD1NT1ABHF1KLUs1JwKM8VMAwjPd+ttHrXZk+1L
/b4Ki+hjqyj7D0mCNb6AVrit+7QSxIH3Uoueb+Tl6spfhpFMj0v91CHu7ufYqig2
q5DZKn18WXOaS5LV6JCKocVC6qOwu06opuQ4mTENTEv1vH5Lh5SRrvd6ejE4TLdp
8/Ijks1E63G6bfNMIM+VshC1hcKtcqZ+rRyOgJ5n0hQPJxbpmv8tHpq9q9ioOlPv
svzLBs7AuLIqMiaJKqs9yBseoghDRbQlpdS/66b3oIG/6TcN953exlvtiYCzVx99
DiHnvIe+iIO2ov0FPiwAIEmc2noFTM4mH+ybsEg5MELZOGZOj8XCWyVbh8G/XpV5
pD6WlQ3Zi3umFN7LE1KQ8rNq/3P5I+u1yyswH2fINwQtgiA4lBB5QsCwzDbVDusM
5GJrI+jnR1PAbXReSMid/CjXBkJbfhxhHZeopDi+1znwDUHeWoJo9+6rcO1s7tB7
dKRClMBGYO9dGmvvg3Pf57G+cMU1SpBeZPIfOT9J7a7+NoOJuUgdRIO9R4iNGHEz
U4Cdb36+T7TYUJPtdjSv7xNzP3BXq2ULHvtCKkzF1ohZNsKWimmDc8JOmlBjklL2
XIVK6+k/bKuo64pXcHsc+5qhuMzbKcsHFMmwOg47dRYlsvpgCxu8Ae/b6ve4tNbQ
Socj0fMeJnjjQ5RdFLSD2zqFZfYtL1l4pUpOL0BodI/ioq3NySC9ekrlXqjFJBWt
J1lI581ssw1K55VZ0AJS59766Ufti2MPebzG1VVseSVZSSR29R+k2vfItUBkxP0a
x7OdRjhFO4BJP+Uj/C+5e0pQlPMZb/7hkYQQsmSY1YYTCD3B7GfgvLjkXCXvOx7Q
LEiiGmqM//ltI53/n40BqTcNOB211e6dSzPmJOH09nRgNbHbgMbQLXPKmBNfLFpF
HxtpCzGNF1JiRvHDygwLOnuFodraH6u7f+Mq0wXFT9DEMytJZfPAra6XyP8aXXM4
zPTrY1sNKWvRVB77zsFB6PKfRS09UEW1t+WfulCyP8bQIdMfvTwVLfeJJkpriOVC
B6YAXBUilwCUNCGsaFuzFcriPTXHnfwVl7vfkZaNB8K6/IKsLBwSdRh/xyfZDBlE
152lPS0U0k4VLyguoZXVXGfIdLJ+tFHxCUZ1r45fBvnkXUSbT+syWgSnYvHnUxJj
odR3xuUPd0qAL9mMRyhyQb5NeAJb9uXmswsEHBZn/r13EBPNjVji1Vv81mQsgsqw
QIYxFPHQcaAGzoiczHtcL6oDEGuK7EgKAbeF6DJ+/7lRiHChmRc/I+ad+H7X/pNX
6/W74jcT8T7rrNHUit3rn/BGtPu/CtfGNOZyu5bRBQaIPiyWWVIllW2ulgAqDXpK
1BYGC+OVPa9CjC6RYC97gKKNHL7GvQgEVFr61QXPW0QpfIdd++CZzy7SH2nuqFAc
Mq294XrqhRF0pT3zSWPE3jtfuwXGiuNoKoEVQq8/A+mx1j0fyy/EWpcAyErwKbbp
KKlyZ+opRJICa8hbfrbRDxZjz4E35RkL1HQSvya+3UIZaeikzEGzuAN6zbTW/vBR
qZxiwuXIIi16N5pBW/OeykTJUDoTEWcJpDhpAFpqwL/rwkhq3pw+srkJshK++yDh
0S8QzkzHTh+GOSs7bW4LtXVwWnO3b7c8FN5m1+zveULiE3bGjvg/VQtJxMCGiFqZ
lqtYBFggvmT2xyOQnCyqiWTg3tAomn/Y2K7ewDmPFlLQlLVE3Hevh7ATaFKXrkJy
LFQQ56yo6+8kqZmtDVEwPGFiyVFqWZLS1IZ2DrEImV0RxK2fkJ4V1O5awt2F/1uS
ELSe7ieBZp0LRWEd0gl49L8aq5khtMSsmLdVi+ssmmDGnBVmygwoDVTjDl80ET1Z
v/jgUEsnAF3IWCLPwaVkBAE/4uDNKqluWtNc2BVJFh7iE7DITO1X9WPmcFrQp0FE
XlPir8j6Aee3ixD47pFmYDkargKDi/f3JvxH4CwNuBEjcEfnDMia2jQ9S8e9w5y2
YakR4+1NScE/QpCU13cNaXr4zHsSzalT0axxr6KZer8LniPhOpXosC8yh0S40uSr
t6q+wm5c7F2c2wEoXmlZQ4ihsGjm6gMPVsPUWIbrVcDeh4mA/9GS6P98RUtIqrug
al9k/7eF8OFSw/83SUX1CJvotqVYbwfaftPCmOi6dD1uoye3o0u6S3PgW3XEu0xx
v5SUrG1nawUIeC/5WVX5Qcukob5tlWWHHf1pXYXA6IbvG4wpZHNC2ttsjfdZCZ/3
Z1Uq2rwJZgzuq8ztiDWRt1i7ODQpvYHWPwIuWlD/AqnWUJcf33mOnbG2Sq+dShuy
7KJXB4rSDqvtphONPwKHXN6lEn5E8qJUHmlgWwpbMLCIThekbKfSauW6WCdNuAyn
WLNhjmdEjc1hrAZPGfCXa8E3bSZtt8SVoypq0iSpRRXakGn0ozuMGBjKAv26YaKo
Vv98wN5y2AeJ114V1rAui4PBLQRbQygxLRjtVPabhGGeEpB0VnUPSqgn7HxuIdX8
l/xRVPwy0MFzu1prg23qDdc9crtp/r9OuGr1nfwwn1SOmOdZGpwgjv8PFQqqdYGQ
EQq2qoPMx0e/TGgXigNfDBkeWczoKlopaRlDUCYpbQpuyZ8J5YaQpsTRm5NS+kUu
ogI3sJp1AhucF31bApC0I+UrEcY/4rhJo6rW3ho+O0kPGyRUKZ8Ffo3hr2z02LBc
mY3HGXfQhEslHP6ogbCUYRYKyD/zYCWX1E151nLI+CYCYVzMqdJZTulQFP9QJwsR
aG3Dk+GEIUC4Qgsb8N8sT7b3T40iMvMBPx6WklqWhfU/q4sMBat+/kGPcwzDSy7r
A7GREmdAR4cQCwu26rDLsMIjLliPvPalYRIJPici5NJWmqh1wOBkL7O8g4/r9sTb
Z9boUjDsrxtMHMZz0K5VRXyFKxZkPaSIu7GEL6wKLMLqnyuic4+Z5UfJtYotUQ7g
/g3Z8Jz2CM/5gCCsCM/uecGibfpSrN8RPFiIIC+x7eRFsBp1sHgHrWFBVARYF3RJ
Kh91fYpUvKDbtKuewQbxd8+HEUmYq09cAaUSkAxA/N7GdAeSGbFxBAVIy6XGkuLn
DzX1vMVPJkhr9/0+QjEWUjgVEs53HS3Toac72dEtjp3TaJjVLICp59ozMroObLur
cekRfS5Pw+KaFggM9bZj0z0PaxVWbdaJ5oF4027NXnTvOyLc1nJvZ64eK9XlDvpA
R6aZZxaUcWem8Q1N+QGXAqT9e8SDemfzWStJQ+8CG/p8phWE8skdRqXEmktH2kj+
lTJAxSiK2RInYqBH7EiMVL8jnDUIoxKIUJFFjC8moYOucSK32y6Q+xFNGfB4PJT3
YfCEcAYgDKh5JX5P0PaYWxC5uudeXT725G3gr3hH/o/aAYM/M6kmJgNHx6K3MOt0
5SeyMipHaMTZRGfUsv+VMl+vxAVJAz3UdrP+VsOpCwoHIv8XgemU9I2gsbWPAtty
4PPehB9pTj6Bp7kvZBS2/tu+ZVWM/IgHyToXI0TxO9g+egkEc0m5FgnkqhK5wujp
M7D1gzV3Zf9ygar+qb5kenUs116LCszOrKCksNSenC8CadcRY963BMWKLHE5mXVa
UI5Wg4f1Uput+inx2qqXZXSevMst0a3WmUXjTHtQ3waMV1Yh47CObsDJ0IB/IwX4
soQ3yY6ExoYQbWve1BBT69NcOVtHAS43VwS45yAnCu+hPGV6FFt4MRU+YIlL+KSY
pcRVVZXJiwgsXVBiA0tFTKrFXo2VIGVeEYyt2l3t4SQvLNavjFVSbT5vUW5yFS0z
5hGPMRdjGOPbT6gKj7qkukh/qyFkmT1kNnlXUsU/1GlHeavdtg/Bzze2lvjG8Lsy
nmqW87T7yEY5lzAGBaaAU/rVjWaM1zjFtIUQxE5HoLn5asQoo54yQH27BZh0W8EZ
f5xXDHE5jL19xiVmv+IIK8GyinCo2lOKVSf7ClT2NqeEeM9zj4hlCRqy7PgSE9Np
R1Qa+7MTR2BCBa9rglPfif9RlrHipA0E4fRyXQKzqDG8h7NjjunqvGisKLfBm+CG
jn4GZn9/7JAD3BL0KWbizvehzSTMUORIHEAdeLPtUePDGHHpYVwwOqESIcF43+gw
+bsNq6aOHvn7eP5mZWn2sruIzFfViq5VceJTx3CgajPxPHH0Qswyv1qTFZAggm1r
aLUQflMW+d7xpSE6HfxSZYKLUJ6sQ7n8FH9i49Qe3XMMYp5ZI2JrXR1o2sEPd7yN
DSMGOSE94cSjPsdK63h7z5/jAy6pz9tVirX5g9Z/2pRBFxI4Erff/erjFef4GeS/
dPLl/rrwTlClJ3Cyu98acWooADtOWEwietb9hkWdo+AtPQuUK1lgc15WCMkg58L6
bVIcnQS9WXw0HRqL1cJgSI9lLHLTLyLJeW7RcYsgf+dh95nIhv1LZEr0/V5ieTPQ
k3p2x70Rjdp28i9488MLk5kXORujw3Lnj+iAKLS9pXWtlWTKXvXPEUqSPFuXV+28
CHWq3mXDs0U7XbTWdlswwiqiduAZWyClYFCkjowUKVWkFiCtrKnHK0ivE7C0HqIu
eBwbT0uNKHP+unSyUICqYOUAP5b3Eo9dbK5rIf49A8W8xdiNHOQXbg6emrJuDD03
A4u/PhA6aUyEX+zbxxIDWnXjkr7IXwGN7YKWSBzEN6tE6kkHIQqNLyqcmaV12FKK
V69TLnZLP7rfPilmhPDab/ENIlLjG0EVFWFq0PduJ7fzYxGkx6rctaiGwFSBCayL
wMKA1A1euEby9/XwUiyTEjqUs1lmYD5xu/lQo/6mCiZaPUjdEhKEEyQB/oFv3LV2
ji9ukMpnnFFCvlIdJW7f2KbofRqtBtx4aJTFcFflnqxavxbM07fko7KmWOlOC+3T
IuuX4PqQhYw7+vMRZVDJ/J2xSVThpHFLV/+gcOcSchvE2yEFf3sV+xeHuohQBtMI
mCM2C6JOpb641eMOj0dlffO2/DfKx66oXkuP7XLifE/PEPSngz48/U89nUOLVs8N
II6k9NYDddDQG75ft5JmEwTST9g/0+8rRtOHPDr5y4fFbAnjYxLLSovqgNiHy0UX
my+444zPWAODw+zyteYEmh+4ObvsRGdX09KqUwC2isWf/fahMvnRyKYm7BzN1jol
dF0EdaaMwwyvZPrCQCSnHM1xGOaksCJUYF9DzrlyFoZP+0Pbn10XEQawNNW9boNi
rWtI7oyeJgreDz7nBGR1Zp0EJhxfCBznIgnacoN7QirzByr9mw9J5CKAHjWKRTKz
eWBGWJkSWBJWEBqZ4tHmFHl6X1LJjpnmwcNY6q45z4CCPMJwRfUl9hNuYdKtM2gH
laMMl2LZv4pSWgFkLlLa4sNlWMGtWrRpjUVPtixdh33TwzQSTliN0LXl4kFW7imC
d34JC82mSA0wH3QnG/5XEgA5jdCagm3okZmFBGCGrMzkFSlucw+hkHzPMIRaHEEZ
y86Mf9/BJ0LpTNs9QpBHH/WdvyoA5FURGV6S0i7Mv3K0sGVocohkAZuRUuDO1ao8
nx1cPqusZdqgFm6RPy+uvwKwvC7HkZFDqGlWA9l5+ZuFviMiAt+CnC/zeWq4A8vv
ZcxuD7MXq6X9zpkBCa2AkCz/maVh+yLXduU33UTuiGRxGrFmQHPm/zXWPNV7W+A1
/rE+Gz733aKFFnfXzJu/RnevlX50/mLBKwyjliZLjZZrowSrwu5AFXrUQPOlx+VT
1FJctGzevK/J4qoGrzmjqSzCgmkhUOcz1+1BLDYZqEDVUMMtEDj1sNZ3P11ckzP9
bFWjCKWBLQOrWDCKqMbTsuYZrt9dGLpApD4Ag4PJ0n6DhTopkK17jL83BweGX6ll
cFuruDiabhFF7GioA6EX6UjtnI3OnDoRLE2Urz/cdl0mZwg/fXYOl6nrZJtlfo6h
i+xYsWGpJXVQ6WfaW+6Jkif3A1udXFRmvs5fResLYdd96dUrhsCW07713nOvFmTJ
adDTQbGSA1ElM14r9dBiY9D4vohNJY+nJjbxEPDbBpFdnO5YJxGgRe83KnUcJTlQ
7NCLGc/6mfcw9Cvrteiy+hdG6kGHIqq2AdOIi42LWNQlld0iaLGq39piUi4ePxvW
84mraRen18qIZ6fA2iZFVfS7ogYl2Ef7DfXKmI9Qb6cvTzUTeiLhZOMZbL+dlp+V
x1NMrZGEe5wPd5oAJi0LSFpz3qEUdq80AlFh9pjx9fgf9pTPoJuiUHZy3aB6l8NA
tq2rh4BxBob0ZG2gHKH4WAIIHhNx3PkD+9XJLiA55oC+bs8/ffmm+JGuZgpJM2Qn
ILucRvjw83ZIJr9YU/kKmewkCsvlCMahMJ60uYuCM1HbEGGMSDCVgeTL0f07ah+j
7/kaIWADZZBaztv0TAda/j77K1kCjb5keZSpQXrv/jVjZQpzoyRuqtcDL6zMTG8b
fCihxy/t8K/AZclgrPWXLuu/EsTp0SpUtn/f2mHbQ+HWZjnpPcj59W/+zYNi8CUa
A5Yo1oTaJjXe/KvZKvXQqCxKCP81qfNzVKzGVMHDY/4aNV1QV+MvxB5td4bc/+YG
MCV2i5yD64X+ZcPNOVoZIsRr8bmBPUThG9k8KAZaP8C1ANNIAWCzoqR3zsdK5v4M
IHCyfCON060HjN7ZADI1MQSv/5IR+fruK7sK2nJfCkZuM0MCXcfMr9fRHOfz5KPC
0MYKKj0V5xNV6KTUK3IMR4FZq4aGDGYYTCNVG5RhhElO81IXdz/jnXQh/aSU6DcM
OWhYGjBx2YghK5cQJ8BkDeac342OQbUJm7xJWYYXNhGEfwtMo6NhNzkMqn2dklL0
vUbY0iBShOUTix/ZadQjMzVwD/etGVHMaqSR4604nwu3cxnCQG4XKgu0FmQXWux1
vy8IFwiLptmQApbTwQlzykXqXP2c7rhs61P7Ko8bWxn9p+AaTvlJMjxwsKmNLwQj
liHGk0V5Wjxn3tlZMNh8g7oRpFRUxFD0CfkoMu82oQnyxbi+cauA3YsVVA/6vcXr
LBF0nKoEvWFN2Tsg7E8kfff+tM3CqufUFxIj6YEDgcK4YNGFOXioz99MkNES7MH3
yGFh3KhQzVF86nX4UgrWY/g6lyF7mc1VvRPvLln0/xdWXHGKXIWgW4Vc7OBmaePT
0OdiwnlF7xz+I5VR58Wj+sVdIosjYYNuuW1qxV50CBTueo95OyCzPcJe/PPysTiU
5IPiyEOVeG0QfsKY2taHU49clmHrxxjiwUpNvWDVf0dQ6sSxtMDWhgmYOyuV2IrY
1tIAsZyUD08EuWDMigdsvksdA+AHbrKM6HdK3DZJcteE/Y9DHGKHdodwd6L2lbNo
Fvw2GOpeRCBfL2JbOp0NlZqnS+QnJ6cyKsxVbEtPMAVuL1vHAbW57d1nOeI1Ncqf
nCSNI6jJ35LR1c4OzollmlbVfSmFOe1rYWAa96n1HOGIdoZhW1kSH8NVq5vNsFYx
SynpBYYqVo7xRoS3umWRiMKTQ/ztYHrrk2VXhqeDga85LPNRliWJKI5yK4jhkF7Y
rIDShACY7l76J/y3JobBmmj53IU/j3RMZVUI80nQRfbHccaByROXoQZdXTB5PWmb
k9kKH6xNxmtpy9MhH3WqenVAd0IJdWEXkod9MoeTW38pTO0KqGQwGYhERZqhp8sU
kusrsWT9iEe6sYS0Bc18lxkhGPO6POtJoblaDN1imTLULap4TEVHSLRt182Y75Dh
x8g7vk+jcLYA1GMf0yjH6sEOv5ovbVLab/MagI0PxtLnr/n2JGcomm47mOcVbZV+
cDes078vzfLz31EdLZCGjD8WyqJTRegs+lCzcumuYmGN06lX/GdT7QjGzz8I9uZK
YLLbbPRKY8OJrNSDOOv2TyTR6liMvTXqb+r9+QWrxXf1Cd3IFoL/u3Q32fq7d5qQ
IYVOuGH+ppFgNL6kGNrMx83Wllk85FsG2N/XaIszqIz857V/ZpgT/9wBC44RdUs5
ypFoWZc/oG0mIny1g7dZDmUUlnI0v00vjP+2BXaoF5KTpf2yZCn03hqlUaGC5qBh
jiwI3qWAb6WekVb8QwnQrpcKzkxocS/UVEuBE7kzv6knArVW8KlP67mVnKHgghVz
X07tfksVgrddKbzf7+C3q1vudz4Khot7xdJ8lQgf+G0Hp0jFmoqjSa+A+xsuZTCU
4bRmbnnqN1AEleS751NPpAnlszLV+I7IpoGHxabp5UixYuWU9OSlUvw4Ys8gmL9/
vJ0ZVKJ+HczbcANXpPMIgS6oLtcjaftAc1TIEisiu0FVC566DieNrvmangI2jkQq
TFS4Zf/BNzEZxcCkJZQoE/Qk1ReTlkJ19DMVymF/i5myZiP9NGb9O2rT4xYVefNw
hOKDtlG7OhK1W4k646rkUpesUTlorTHWL15FM0Y7ERn9lsXgyc2X7d1pNaWXaw7r
X2/tW1QF1unyCMIxMcy6waYu2iRga5qnOXy8ywk3dfFVv5Tq5uX/54GM2rGGHpu/
4vsDqXOJhCxRlqwF230ymO7IuwOM45HCbb4Ve/mXi4k8JMHm5Z84NhOCOyjrE0QT
guI3MsQaSxnkzKV6UWNKnf7tkUEW/n1jYZS6lZUUuQcBQjYgDNCbl92TIfNzHIKO
+INNUlrPXbSw3Wk3M/cKvZT4aaBo9fHZUcF9RY0C/37ZR+pHPt74ionFaMFBRh+U
74EJqKcLc/HcRDEfm2u4dhKAR51DMfvz/lPi7dhTqXgsB7Wp9x++rCOwbR/3V7pV
Ft10jJIZ91ooUKk5g8Pd4ksSE9ukWPChszbzO8+WdF5Mi6+8VHWtb9X+Ru86BvnG
JKUJBgymwFqfnfYII9YtEY7Pc/QP2fihD95UDz+UCqefaRAfr+JfaRY0FORz47gi
cEmymsdu+oQ8SgLW0K4P8JAv6EpezcRYxtpVUc1Eer5Svnn51aydXczKGczwdcCu
lArLkAOMeuDYFRXR/KJFGpq3e1nN94XpZ0wZsbQlrcvCx++h7728pQGaptqy/TUh
s/YIDA3p5klH+XPHnyK0yGl62nrcxnj7of60q7cyJ4yN+Gsx+F+UkzEcUwQJXVQA
f/P0NzePEh3Gu4aPhCQ7Y+tF7RWvmu0VjBpevKYJqw/rKlXsRigoiHMZPJBDxq9z
sJHVUhIp+Wzn2H/31D1zdDmPzhz4MNL6DL7W/KzjmJ+bvPLRyZ5sVnvbRUKOtRhv
JERcuAmFN1BZ0zYYz1VhtCq+B1+hLYBQUdr50qCV5mU/a4spcbuFbO2U7LqsnNEU
x1P1NwnzdN0xzEqaeYMABtvIBtpA201QU+a9sGErPoMqcONF7WwT+MRmnJPr9YPJ
VTOfx8djF2J7V86OmkAyHZ94LqkKvSS7U6PyqcxTQ2TXVM+AbrYB1Xjmz8RwWX84
J2qEz/DkKzgUhnWaTOEZaF6A+6VJcuxU0WSXFo5IP15y5xGl2N9V0lC4A0r7ghtb
FkheIlk+Qa9P0FK6L1W3QZfl6ugbmAaiAbvcDQsCgjnSDFu+OniG/dctC/Iqvpas
MJO0cMRXDBSGmBF0qTsFWK6f6+kUagHjHnkw+PH8LmgMmzxiFfDtDBbKNub1tpKV
2174JXKbR+YoSouSLIKqRzYMD864mclvvTiiwgyClckS9uGruufjrkNY2pkbiuaQ
W8mFGpHkc+WPU3HppWIQkZEQt5YFW0yrs0Onr0qLP3eOUrutDjOw7jh2LGOBM92P
EPtv3mXgLC3uEhXV3eUMIXxnp6thSXO/wk9QD/xKJSlrI8HvzLprsY2GurpdGWk8
1EZL8nfL9Zp8NVjv8Iqryp3InozRs2Pg6QWZV6GvoC1ertDBTyEh7TkQLXwaa2UW
k3vHiqWfPYi8sygkzc+8CvJH+PBGg5kMHkdRyzERwx5oN0jHxJWKLT9g2sCMbt34
KejfAW77HYtBP8vIdVqKKyeCzvz1KxYPkuoTeIahdzi9eF975pQ4gi/QUuxFo+xx
xGBQkk/K9sniNKDcM5xLPV2+JRJ9c4I5uEh0I/L8LOOYWm8aCV2uIuY25+iQnYLV
RlLE3NoXl3M2NH1oYyBeG0lPyWoUgF5mRK3QJAt3bi9xGtlPxSLl5FjLOgiEfSQw
kigF6AnP37Qlj0k6M9nzq82iLnj9fdMO+nKJNj+Mo9O8pjHNkowjt7wOFt5Gs7Q5
0/ukLxQoangibK7IOLt7boHnPxicSxcF1gaVrulwke8ogsrjgUhdpLR8AaP6TrNK
d3hOPQDXv3BRHEUdfAcLw5EBsD6k/KO+SOrhxxmRkIDxeaLsxj6uP8rFCcIzWvQ9
hYmKhPzhAYA10w5Pz7z0AIDZHbYP6BI/+5qGEm99/VmL2FS+T23vuJQY5FXgaPb0
/Hfv+UQdEyhbnWnWPoZYOiw1umF9fSWm+0RNRFEZoknujlm//BmpYzfV4ZN6gHSk
+LC3w+j02fd8mgE65GxILfxZTIGYzhz7wci8AxYPJW5RDSu7RyN4ZwxlA7kle1eW
NN9yOdTSIiT6zvZgtISVdL1W62B72fobUAjX92Tv/8lJrzc/utxlz3a1eb9FCnwU
mpK98Hmpry7AkvFevGE8OKGiWCJ39GSIpuhsK8V5OxptDQY13VvHH55epI+bUvQO
Nceng+x9mT5D2aUr74nn4WBnkBh3Qp8bFcayC9CA2s5i443JWrFFY2XXy6X6C4lR
RyeBFs9jbgcIkWZ2z56w5ABAsenRRNOKxJU39m+Z9Su9SFne6PEtdN8UdeJiWt1o
3oryoUv8aKMvCxqRGOyD0ldSJrrd4exEzCrbzt6f5LSTFoUMLqUTsiBx8Jn1MfdI
A0IRzwb650UngQxIMg2cso1T8BlCMVBGVotkgonKkrm4L12/GMvMI9fOUiUmU6GI
4lBvPuE5E5TORT5NDBCIwX2cJUXrYej3JQ3y5DlEHfhfXPyCALBLVbPH+zBiuh0b
ZanSi8gyV7v0BJA/cMhE/7a3t6wsfrx//yOJ9lvjHgLDXNhc5dqfKz68F4+MMvpe
YYf/vET8lfr49qvbOhF4cxw7i49tMSV1X7uiwmmJyHHWBvrt3ajK24by+Chthbe9
RIhEFXba0YAZmrSHbXJn7EeuvvkUn47+ECeybY8paeehcerhIoqLQR5fHkZd6t2J
0Aktne8+Bw7tHX3rgnUXQso61RVH1lzqaVF0+xYEkSADcJv2TdzoUBD0zZ8ARlvX
Vk5R4lBA4+py4U73MdIrJLJvzAwgeCr5Q8ObsH6XSWiPM21kaiaUFEzxi53WzEel
Q5bJBYMgHd5xPhxbWbbDt038fQX9ePVGQ3qQJ8puUMZHOsTOooR5auCCdqosJAZE
59Lz8RUAZYYIGkEXxuXPBFl/acyx+ItF7s2D0qMqaMcZIJ9+i+6zcgpFL4M2CQFq
YMqJOfMbYhZ1bHPXXRl8I75zTFZWwx3VH35MLvkoo0o3nf/ISXZVR0XzNI111QZh
7tVojK1hT3FpkRfcEndwJ6hRGr4AryyEQ6aGgKJMp9ecf/pI7NaxHe+J/CMXHdMK
BM0P+dE5n07c+uPIw8uMS+l20kDSoue8TXV/Pb5zAcmMIGSyGMykn8+FUGnfU9Qb
j3ajWBGTfmxRaOkaVTxThfRuifnWaWyEw6p1VjuFn/vOUVnY5HLa5aaQ5aJsfanz
KpTNyKiHzSh6+tNCEoBzXw3wjkYjue9XOEfkaPEj2ToHoOf3dPplw47MaD453sRT
sfNAmxWOKuCgYpO0YNGYSozkA44iF+ObM7VwRDdHjfCywSIGSEVdvI0oENpExZpT
M7erGELaLzVjJgQnMxv2QpgEJowh2T9OGJAuyLFsWnSX8XhsQslEO4l5ls9HLar8
+Ul+utg7Zc+m0yI3UIzT0D7L9JZ6sWpkxNZ8CmrMDHNZ/9KAoZvXa13RA1au0wPS
vcFTca8zxj0zj4+cFkVBXntb5PydRVw9xvinM+El2y/bGSLavt+Eocp9h4WjGLdM
7oj+xusGpbO1DlmEZlkcv//w2qy0kTD3oqbWVGS2i7VYssUHW48or4chTS9Lmbfu
l9P50JLM4Ar1tVRZtvMUY7TnovaKUX21gpTUujUDDfh9JmDafL1sr4fRymeIMTC3
nkp3PcOO4ocOljNR/ltg9JP5r8mEIZNLnJPzLP8ose35P05VgGMGCwvc/jDeMVe7
iAw5h0ItN1zNibm73IO0oUgl2iTxXUvtQi7/fhuBrY2yFJSMP3+t2Dk11m1ph3i6
OEYrYuuFI+HfrbMFWOXrVM2r7JKBlTvZ34yZjHWgYPa1mVmxPBn8LsFJvacOZ515
2U1pqXr3nCmdODUmceitck6n9Z5iPvxrhH19d7H1puPEqwtPAevZTMu2YZPtDT1T
S9zumUeU8fL0bSPAAA6mPIoUMUMvkbuCDpRPK8mn6kE+nGuIwMAVlI+tE/7O72sk
WPTws0WLxnGob63xb0iFWMbPEVRAfvaofUoNw6XrTtd5H3MVx+zPc646rihcAvEY
NIRbuNBuZPP99J19IiyNJH3zYFwDqMS+MqDLiFLl/OLP1bM6TLDWEUyM3hOykf+l
rqTN89lVu0+bhWlxyOgotTD/xlanZ4RC0kgg68Cq4hR1e3Yev+y3Z2IC6TAYxJh+
40YgaQZzEoKYs+Lh+S1fwoaPdG7LIG6GBMz1Ah/PiDcMt9xVEEUtkv2SLcwoPKc6
MU3sbz+s6Aq9I8tZDsSL8Mk0kmGHs5Jx7ypDswgy0LMxOGAGcZfwKnXCHNRfyluj
CdU+BmP/5uE8SlKrVLrZI+YsD+0L3PHptQgqqGx4dWDylUzodhrT/zgKVKrsrpNY
2/biE6Gq4+y0ePg+oHzL0twBkhnxDWzNybUTp9lsLdtrpVU2aUbAXvrxkY5voWtI
Mkt0aZNenva71by1+xzkiHZHcxeE3C1g/qwJdfFfmu9VvhgTbHxh1HpjeHf79yAM
VI5sY0jtT2g7a00XMPtkgejYykYySBuH5VkL8iP9SjeUL+CJo1q2n+QC5cSv9hwD
aJzlhSFPoH2YVPxuqwdr99S4mJ1XU6eCOgdsREW5tc0ZnzfuiCHjSRtVOVTpu4aS
+zx3wvff6MwyVNayYVHnGd6QoWLAG6H943I7yMqInPfu8Y/+ZM+BlBm/JuOKxwvK
9kqxm7lIB95HRF9tUWX5fn7/jYYqiuOq3kLNeLQcfd5pmuwv7edLUSpnFn2sKnZJ
3C/UKmuRAdaMh1ZtjzJfiGuIprlQn/GOfhdajQ/QNhG3JgQ3ZWvY8Tavs+DpHJMh
5Ge78S2QaWLwbuVCmCeFXnz2ilSYZmIaNb0/73DgN1ebx6OkIcMQpCqKANUQ3LCT
qpDII+xUQAUqVQzQ4apSS7j788xRET29IpTSobB/sLiISrl7y58MuPUqaiohvVQ7
pC+1rPsvEcKQjh4IMn6pD4DV99QXJb1l020ctt0T5iT78SAJCHXMDrQQM1I0i+Dn
13E5z1D2p77wk0+G1ORkEuiRI82DZ6qYeGzMVVKHaOsdbzxIEcOzS8mmN/bTmjlo
WKYxrQ1rons+RyS4SMBcjc+5zEV4VnIa3Ilf2Or2V6lXt+3PhAQmoFGrJVnfCNpX
tMkYN11EHrS+DM55COLy7w3XXQPPppqikReoS0pqs3A4ZN7YEqviql9tS/D5TT3g
SrSZG+8eFB0eC8ak+ncYRAvQE9EADFV45kQ008wD1GB1YIP2zZJ753FFW3ZAWlTt
tNUJ6S0XWUy5Lhja6j6f9Td3TfmYd7thuMiWBOuPwT6KFyL6lTHMZuas4dS9SNMJ
aRfIpraPPnPK2oKz9dnA3ynPf/QK8iWC3lWw2JddZVOtdZs4IhsbtNMmrlUqQ0Gi
rnM7otyVjYql3xk6SpW2igemRFSQ/21rT63OWicz07MuINYhh8eJa2Hs3bHuNyUg
7EC2RAOiYl/2AlA7pS3zVjUnmnixV6HNHQi7wvaQGk3/oqDl1P+eOBKN6u4Wr3Ws
1JX96iIr605VFlLXorQHMjTxoRN7VTWn8SKxKROUaIauqJGLMsM9P8q5XfDTFnJj
6BxX4LdclLrh7nO/J1YSifl4s5tAEC/lvWOZgHtFtk8F8Fyo1EjXzOd0odLPlaAu
wjX5nl4MfbOaO1ZGLKb81fACXTGry+D300puHdVaVXbhSgIWOR1H3yirpkUNh+s8
4VIGCjIqTD1DS77p27L2e+ZtVqRlm65rhd15NFXP4FJcLMfbWJL7K7YXPYHXGg3V
NK7sHc7In3dxzxkrd342PPWAz6hi06tKs0gPI/wabIQbp2lSs8jGRBIod8CsdWUl
ViRSJoK+F916Y3iuP0hpJwBitv/NP2zuZdOTtCquxG2XEmX4uAJx6NaJ/BiYzq79
6A8o2CviUEN96C7L54iT/9wnCZUZ3ps4T7DtQLMqZspkQepIBRb0NPsgX0tuRGVi
Cb61o31kqDCmTfzaVdjcCbWDzE3koh4nBodM4WiYf/LzUnrirGc9RWC54EEl8gQs
4I2qL2Xosq9WhzbhM2pGt/zMnxqsmqe4lnG+QYPaiTkTMaxpnfac0fbD6mZAu8pw
M3Ki7GjKf1OyXIj/LHgmilC0t5WNhjC1WBCWCDgp3t+fHNS/q4kA0c5EP/wxTU37
DbUH8SvrDRMhsCiEXletsmiy4ZLWyIfwbtldB47UfDUTTmS9xXySFa43omFZDBuV
2fzT4djTpLkLDyUajATptcWMmZxich3XhXd93gBGxxhZTv8T+cEalfaZmPPeLCA8
jdh01CXU/V4uCATTQaFs+VaoaYmNeB9+q2BqeAFJ18yFq7vr217AMYGBEo283gc/
2nCw1lDjM04abYV4iodLXKWYn+O+TTv5PDGp+bbWztaZcR0fpNrsrngqgwGiSFLn
FGWlZkcbrQan9kV15340vfTMj7nDG43aRBdZbXKD65lZVBAddCTHpFJSoGPTsbqp
XyksdzfpjIcmzLi8oOasaeY6m2+y9bh/V1+VXuvYdD7MU4m4rEyjG9ujqamAYvkc
nY7aXulY6WkNSkNRJLbA7rDVP+rs0e0coGvZ2BfmjHKRoEktqTsiS2hIYdb4xkpY
GXHIP7KW4wc9RCpr1WgEtKbZ35rr47s9wllluhWpciheVLVt2ljeyRIjWC+ZQNVS
CSbz927Kca/gqRO9Q+9iJMC7pn588k/cauKV/lTGzpXLG5DZXrf4rQAT1paWdeoF
yNanrVDnI/YeqhjRcZuGiTc6CITysHa/qBJSJJSXLkgBVtnuEm5z1PftW5gkAFhg
ufjN7eEF5fsN1Dqqn2VbgbIDR+gL2WYJoYU/tFg5v50yFvXxsjSchhb0GsIYoeHA
D+lmy3mTD38NIS+F9jTq7z65ZOFR7iIHFu2aSBElNMNOphMf1tCuuqArVim3eWPu
1B/29z5FBumPNVY3lYS5gyzUAJ/e8B3075vFo7F33VYuaZaiQj1SgI/X/Zuiz5A7
dyc1v3lSZ+AXOtDPGhbCJXYdMk+K/S112SrIrhRozS1pmgPz3AP3fHPAiLxkAKqq
A1fjQQOkKwu0Vujo1W+YB2qRYIJceShCw4NEg5sWpjGK7QuP1cciHvNdSn4h5AzE
Hy4txOXd2kTdNWYDse/5iwbYPxpx9j4QzCSirTklSiENq7RQDIqdPxqLlvT2JmHW
UT0/QOX5YD3PQ4tfY7pTx1OLT4a28uJnsEcruR5z2JOjsTAQDNXJrDuxjzn0QToc
89++o9Hr2O4MeNL8F6sbvmVu64+ev3l5KSuNLe6jXsh0+lXWrxdz2/2WdSklZbK5
NSrdncEb/U8vNgnpjqO7SFk1LrAmJoUF5lixkROLd8uuVfWbxvmh5otCrrRhfB6W
WLdtsLI6DmcmLyuaGGhPvc+d6wOmbWq43pXBM5YnLv2IqI9567zTG8lys4oc29/w
d/XJyOuWqd1/Uuff4gOH7pE1RDIHMGNSunMWccvPoSoN9XuIACmlZ+zBc82eUQic
v17tzd6hZzPvCCqpXW0e28GhqkPNDz8xT2ulzvvnS70TudSQaWney8UXa3BTjyUl
y399K3ziYON6BhSujNVnI1EDDbWWHi7runbuPWcKpunPrffI6b7qV3AUj2K+FbM1
ijxJqmlEy7K0RT2XfSGiI/WupmSlh3kDYw5g5c+qIatJozjwY5V0CI/sWRG7NFGX
MD8e/qyHHsSETQ4krtBZZE5e26xRxNyL1BJd92gwDbmkrv2jijcw1DOVby6x0HwH
8oCedV83ObBs1c/tr0xCF17mDGo7eJgRMJN53vgR5I+qCXHsAV3WKPOXde8ryKcO
bjgR54PWPb6GTfNqL4HvU1gUAmusfj46VxQXvpcqe3ukFvDDfHioko6NGZbRtaCz
EWBiFP2SGoNzTUlfn1TLmvT/JFgMCv0XeHyxZE6jRw302x4RxPM+gEHa5lh4sXkZ
imrw2Q1D1KQ5hUxqAHSfTKxqMiK/4kWxyzLuHBA3XK0HttpMi4Gh/b2AuKx6fP08
BNx/UMhuxEazh7bdvrG9oKRbD7QLf7Xb4TtKOqsuUDS/Rrz+6KxpCxeQH7K3pLM0
bnL10YfL7grMSaDeZ06+CxzWSbJJZ87ABmcGhK6RuOgstVBJG2kMiyelWa9n5Pp2
3e+ti7G/Wn+guE0dDslBnvroYfzoKnMN4YI0stt46uY4hkijXMU/RuFEOASPXKU7
jn2WrcXm39qPtqw1esy3o9I8OFaOYYwdnxQ0KHuTJ1WYN7MHX4wZY2Qh7Wu2VEzc
4oDHkCrw2B0nC/0PiDHSWsHFdbrKBIeEW5qh5+pvxx6+cOLYSfbDFFQdOQhyx1NY
S9XA0whG5dOfu4/FdLMnoUQXo/775azRTQnF5HviPaSC1itX6KY8aCRJ9+SJwFRr
4Nq65leTWrfWCH3EhxfXGyzHJFjLxaUrvKDxxH1rGiAiyOF+xXaJfO9lMVPIsHjO
ST+DymHuPJ0/rlI8Zf276/7qgT1Uld0NcAbw45e31ajrnRslVmR6xc+PcBG1HqNz
yEy5KbiBQFWi3hQyftd7YEnm5cpn9sFJYtM9ehZ3qawvLj/nIGEg9cnIYFLoaqyf
UoiVbaOgSPvsHyXyW1Q30m7x5LwiTg3mkXt9DOvdgZyP/QTKPJwuOCULz/oGg4RP
QfNjT/Y/LsQ0pXRsmfJRsYYQDkqSdraF0CxqTQY2dJwKSuCpAEljtvIa0zInZlj0
ANHu/LJNxBBCu/NST74ZN9dfr8zpeG/kmXwdgrdl5j/Ab5BIyXGWNxDgbxoUmyTw
0v60toamQEfGXLkv/6RkCKcUmeapIpzW25q1k4aNf9PEKagTBX8qyEtwVOaT8Z0D
NMH2DNGSpWWkIM0hsQ5ifLr66c3ZSS54JK+fZLFzedNy5jT01zbqolnBPwVQ++wE
0x8yl5IzHxFqFAZaqDKD6i8D7ypLO6KK+XVs7JbAnWGl/Qzj7wtlg9Ebrpu9pEpp
l38c7dQcLe1QtMFtuhhAeDgKB9UcljXucauQGkyt5Wj/PxjIj14VEvA+ZFY9jKtU
uy0Q6nRkrg8yVg6FiXjs/R/1ZTFLlXXByiprHzql7pVI34xL8ThphVaRM7vuS1d9
ZrMzlxZ9FsLXd8xrscNB9s2U+pwpsdzFubJX6XCLHLVraVYRgiuF/aDc6mE2mE25
nA6xVjHohZoy/gxZhkEf8LWfNr1WbniMpUUgCym1HHDYPvlxoScT3CKPv2I4MNRI
Rebjv5qxD9zZkKR/78aI+F4rD4RZCDQrLPGpEVmEunmE6c1MJxlXPOzKj3q/AfgN
qK+Yf9liF/XuKVYSdWdXwdppql3YWQAqWd5T8Z3lhKeNARtFGo+SwBQeJud0qS/P
snGfkZ2OGG4KxEBYn6qsWzgy+3FEd3i+tadWleQj6WnjAQ+A+PWznpWnrJbIA37f
LYejsRiWOP3Zl8EANiBmoqKvK0JEiSmMuzbo9yQmCmhrrKRIr1eKD+I/3i+wVLyM
73dfWRsrOwOUE01Hqb+qj9mvlOf8UNPctldYqeVmmuskR2kzD53Zrmimg9kMnfnu
uZTj/iiiXjzp5a8yHks4oyYvbO/GejUaVRBqRwIPk7pfX4i2MMPP8zsqeJUcnJIh
J9NU9av9sXYv903tkSk8zXSUa1ML4PmpduBzikjmnkncjW8UakQfbSLXk4wybe+e
CyLVdZ7UdrNcKK7fVGVE9B36CIMW6dwxuLeAO+qiPvlhDHH9O8wufpsXcb+/1DBo
QeG4/t/heyeUKG9UJJNT670LrvNXfHgcE05Rf3Usi4UCN1Bck+Nza2g9VWyabRXj
MPZas2Qoc+P7+JoaH0HfDjHbH/sdbj5jR/JrLYy5sov2kzOoda2uQGhH7HU7eSk7
TrbEvz7UNNCA7yLTBikh6+YXgpSfEeJ+7Y4MWlvtN9LYGzJ3p7g+rAS4jP7ieuqv
FN9I+EkM68EPdyA3m+8/8+MrE/Dg9e09zjVLPocstM3BFVSx20pZAEHSASCkzaad
tdiKYx4ReeLJw8fynJFLZc67igPjdO3RDzPbpBpoBLWUI2dGW7onjOidOZNukU0J
T1ZYaB1NUrTKlA46Qn3ykgD3FRIr3E0gZy0yI47qs52F+6udkyqbBeqUfx/HQ5LD
lwnptc0Ey2GXuY3X7R9Ol0RoEWtusiAZtPU+D42FTgJPUOcqflC0GAkE7pjMnQPz
TLaDc4rpG20D1FcP0BYLZjnQswwHq0LbPb5288ZnLTAcTAVs9Le65P19PajJSiiI
XrpoaQSVO328R5gK9rKBPAu7nDTtzJ0R+Y4vMKxcaTaitNtjols2HB7O5FaYTSgq
8Oqe7oZI660DNLKHBYonjgTmQ7lF4cQUY9jnQonTQklXWM1Cp6d/aKket0K5uui4
/tU6yuET/LlIp6sD3sZ9jQ8N4brGbVxFC1lXDfCQcbSe+x5QUpG29GAZlQK5On9X
oMJU+G7H3ecNnYhBsXbHJ5sWV3j/i7H4zbB+QQMVOSrBJasjEGuW9Ri0g7l2coOu
UX2mjUOr55cDq0gAZNXlvUHijYoJQ8zi26F76Eynsm/P4RwBJu7x/UhUtVf9LKtO
v8SmpIjAt/+gEfZCvCtxLvR9dp1zWt+N77yM+37MgDDYpcqo6nzjQeCzwGmzJ82K
+TkivtrMdbwD9Mg+1LkBo5dzcKP4k+RYZRNx7Mgd6riGYjgHWhv581f1a66PL4D5
xZjRPWmSv9RUk9s/1cWShjSxdWcVvdHlChqcqSSVHgKYUMyfQEAa3a+hKxDDBKKv
hoURavR8seMASHCauf0FpK7W9KE7QbPQFc+nINSdKDCQsxwr7DWmwq557iHvRbe+
BTrfvHgvkUI5nvcUC8/CtmUQ2V3FuD0FlIUxhoC0KL2T7bV+xBs3J2kH8G19vH6P
yZ+1kCsa1tyFF8NIVZNaUYMHNAsF5VgXnhdTXA9q7xJDAfRpMvnZ5yysLw+unudV
MB6b8e2TG6LL3jIbm3wUA+81Gdh0FiXPLiJ/NDdNrVsZa6qfevr7iCVBnw8FInD4
1TvDPqNW+UcVmjAXgS7mqN0E4ntwnOBKwiOhKCQgQQXhhFlzp2qh8usiY0MV44Wc
0gx0gxtwik26/LRY97Jn5+sU5DTaB/3tFExih9dVNqlt2behUnim7o+Yo0mSK8GH
IsGtyaEpIV9xPTik1x4Om8TAwJR1k32xIB5orC+W/hp63vvhMM/RMAEVfd9ONpc7
g2gyi28fMDJ8+H2hFBflR3WXf5SFw24+OUJPeeoq8t1eWiqcx1p1pWR0Q8rYidbT
RDael/m8LUodx3D6frGC5Zbr/B94sUHz8+cgTMyxBqQTa1JGqWbKotnfciUXKKDt
JAQMjwQ691c+HlX9p/k86uUoTWgFT4BFzIs8uhaNUbwrSeynwXIk+HYSQL8vJUwd
S4lyAb/u2MlXtOenfpYRs6yiKcELNvW6jYvZ14rczmG6Sw9BGMOE5TsY/QGxvF+s
zWOSWtqodjxZYj/qIFcjWxNjFoC7eWDpKACTYXnMIF+QOSW53LJHez6snGc61VdH
tH9pZzguFiaETXK7+mjJrXuE2E2w9PQcYpZHfZZL0Q9rc+gF4aQsImhcEVWFxDaT
M6mGOkYcBSxz3C73KoRpqmegnvDCO68t8PePkXn33DWkh4jHcdSvtiKNFCUhtMcg
VZjvKo6DwgPDQBX/4HWTDXVO6NUC+VuyorkWzkkLgtXTErMsI9EGK1qbtVmy0ZSJ
7qhqYApJ63pO8skbXYciZejA6V7nJHcX9p2MGJeyorC+NF/AcMCMpeKPxKY0h+ZF
x4exTewWrypMpc07bc4UQ265LIUxp1Qr8ov8VqW+X6X0Cxd8gr7D/sMPJit6z7Xb
A1z6SShjAZCsag95WnLwhOVivRs66Fov38qtmiICDf8p6OpXJ1AyJn/ih55RV4vH
VbjhMTNpWpTX+IYZH3jp6rwt2FM4cOl4u/aJkMPk/CyjDLpaQeHeVeVKuPhPZGP3
bYUTcVtrIhZVhsA60r5lQueLxBFzO31yrq2tpJkVkCwHkkPOpgSold3nsTRDQrFC
F38BaxvoIWrRCQV6wOMhgkW2Li3VF83qEmafauXeSj/Uuy2xOp+wDkwsarhCH9lU
KYZA6fYgk4le5t1cExRiuxjI5LGjdrmB7ZI9ES31JJMUt1xJmJ6LSbi1awRUcntt
4vGp8EhNatmUDF2shIb3VlUSWWnc2i+3T9jD6IC7rgWCrGbgPQLDjG407tQaxY2u
hKwCZrQkvG/cecwtj2yNSjDEa+zsz8sTCCtBHTN1DyCwBnC3JfsgQlhYIoIfl5xD
BVNGwv9MFPqPVUtJdpaQKvR5YSFbvIMFoNDFd2Kmxz2uX9ekirRSO5m6SR2yiqT9
6D3IutlbQMc7FoSmnW0AswpZEheubge968mXZJBAqrBZtwy/IzNV7xRpe94izcqE
JWCjcWor3qUm/PeYAYtxH9Q7t7vPDFfJFUzCZQZM4ufuVGcuAjRaEUlEdMIFHSQK
KfIybyPxAlbivW6VRKPnnXETAT5lzvpJs60A2cVtrkpJ4tC/EwADrKzY9tXcBGJN
OpnJdtH6uWxteii7Gs6zVnT623j3yrOMDgeuz6CubuJYQOHNOTaB+W209wbRKO/U
gqhSVXa4XbP4CQd68a8LRWWRytmaLutJYNeu3dOlFNpAuON3pcnTLPtHZseAc0JZ
MYDph56PGeiWvcN50SYB1N2hJ0uvq1bUuQ/HhIhNEPq85AGFUMQmYzz8WR7SLs3v
YzkqGnQyAELKfvtSnbcsHZWPGGlAgQam7aQfkoW6WIpp+VfPqjcGnumpU/dKtTmA
5r/Xb4JP7ww+yb0TCgC38WZHrwyaw9tlAUCwjKGT98K18vkZDxbtYvq2QqWuuiNT
l8jA7BJI73sfG/QgD7cX7NkF7WPCJyS/fSOGRujgsobDzPqmosTILJWC3dZooE1+
i/VwMGDon/1bWdw8tJ2PQuT0MTNtLRkDKTEa2Pqab9WXJq50X+qWdO2r5KgwHTDW
x3N119MF67aSIS7zhNHto96dJ2jf4AMyHf3xzRWDCyybveYFCSj8hlmFMzpZ+n9F
0RtcKG2hE8xlGkndGr0ov0M1xf6OUtxM7wurX4JNR668K1czBgGbapj8f46MP78b
1bw8KzeVd/pLCGYbEKkLMMFEGstObW1q48wYRMpu4qne/YXEKKpXQtsKYCbyGAzh
x9qLWk/7Fwx1nfiG3RbmM+1UMLqm0h4Y4qODkZBUlCdel3m5hFkw0mPNlNf+HIlp
MMBDJGVxCUETeSyGTABggNBKKIC1ctK9LsklUi4CdgI5FYDFWi6XatWpocEF1JZS
TIi8jPuDnkdGFZhEsyzXMf8e1ZtkPUtPKMFpKfl5aribw/38WaEuYaD7vhJWaS2t
IVTf3ncB+7T0g338VFNw/QWsuh+bzThBsOFw1a7dH0Exnwf5F62PhH+XcV9486dq
OiF/5tJsClpAx2RSdhBuTPcH2Ss99axhBWmqBIUI4L2Z1udVICWHSi6ae2eTzcwU
JeV5LdrCCzSeWVSMXCwVrnRk5WooT5tgXn3F82uFtwGsfM3VOqrUpT9iZ/xnjY7x
CnRPVcUotHkGW4XiIHrGc1YjO7HkAmeuVRRxLDEJJkGnpccy1xeTrzwzm4QZ0LXG
TOUlvP9NTWo1wW95zdBQ3u510CtQiZ84P0dxug/6F2bY3+vaBgRue0hgF1B+eri8
eXPMN4+8wIya/3MXvJJImySXRw8vnARj2WBiCsUbooJZec+G/lAsbMAOO+4d4fpn
IkFmQMIqOPQ+3IEjcefWYQc6t4Y2hn8v4H5mRhdc5Y3Y8UtgQpcTQw6Xtrz9qoeE
5EHLJ2wj4DnjJgz6EWvt//RFPEBCESO0yyiiv1br5RAvxtI4ZDxk8m4AgWo6f3AS
D0AUhJnhf/ZdPZj38LbhMpNC88/guE9LbIeOrR7Pulv+YrXnnMQsHiOXaKCgKWcz
DibiBxQInOXZcj8ciehO4+BA59kWcztyMvD5uVqZeQAGd3nCR7rM/Qi+loK6XwcG
t/4VKQ2BxQhwjSgcFsMPGeTf19jJSngKR3Oie1HT0UgKlB8DX4VUEfSUrmFjL4oP
7yjN6W6aJjr9QwGk37K2DUPyecCmg2Bnaj3LZVksQUR/DXFCgBUb0AODd3AuEHNi
euJpXql8NbrSgXWZRoOUDQE6nSoLuDhmS95F+AHCXrMQGJebWG11DT+KH6fyK5nr
JcoQS2CTK8inOQWWPpYXOCTnhuxdlQnU0q/OFPwTigINU2Der4IJFGPUpDUiyyq3
tHUE8GCK6saIRUJdQRAGoYJ9xl0avggdNNKD70LDGEH0dAOTyLgd1ObHYR18GrK6
s5XNsc5lsuaKVwAH90W/HDzjjnXnpJm1AhFfmUt8TwHUbHZIIENX234tt0tklLvw
uNhe6A6HRPfx8ruejQlRJeX+dYFQlBKI3heumjbpJ8kAFxiyxv8+jOUnLsDKAbPO
A8JBoQJ0mhcdSxAsdmGYoZ9w1MVPCdcftzVy6mCQe1LW6OzzyfM1L0wfB4n+mnKq
3pGy4EjNQavwf6sF0DTgsvyjam8cQm4n07k4iiJmlrVgHWaWX2KUEjUJuHNsnavy
bspd0accvAsKGlWvS9jNk8MlhMSW7cso8iNtXUl4ZgTtQTdRsZTdR5db13sZf/SC
L3P15UQL1s7rQjC1NYU3zFVNDIahKzfud3ACwlpnaig2itfJjkrtLAwtgyfgktJi
i0TRrDoPicI9+dvtM2FJ8lmf2JgW+imtNl9LXRGj3WrXZUkyrkgtM1wWbNiPYdCG
nLlAoFuyRKGpXOV+Syz4oPlbp7zSnqlDcIUANSwGr7t4xea04dmoxG4I60GfzXMe
yN52zcQFY6yrLV4tOM4TMTg3rb4r4mHCRBWwFGp8v2LSy2K0Ac3m7BWAwT++pfxK
5RmO/5azJwxzhcxFDnvV5t8HUcELqn78gaDuH8hgwloRvuPkAaUHOw9qkyGQoPNK
DzP90982nAqKQ5P1F9TCfhq2TD8FyS5Bk19I9J0FizmxgsQm0ZheOQ1dXvmq5gd6
91r4H3Zv110VM1yO3ch/hX3kYgJm6mKuS6dzNRi46jahH6Iz+lrK0kXWzalLjG31
ezAQTmk0nCeGtzyohEFmmg/XkTcBgL5SpOE6cZA+m4qK+bBV8alK1fVoL540Wuza
oJ2j8FqY0vXJYQZ7aQdgZxgHVGUJfHsS8+E2t36FuA2ZR+HLXPnTs7rePWmntUa4
ii4eEkA5eOHYqGdEp9Q93jAfo0l1NwV7hO1bLtuxxTtOVZIR4wRpqgAGmo2rc9CP
jQIwhpFbUAg+vAxWdTuaVQWYnycTpspghHU+xXQbAgCGF6i2AXzMud21lBjui2+T
BFYmQLZM3yEyFjH8dWKW28HbtJ16OctkBdFUExL8CCT35O1iToWMNe4t0Uqgy9nw
b/poiNJUL/PTNsGeaBQROnXVBqKYHiCy22JC7WDX4/unbB3SslfkeVTI0eSat+0d
4lIFPoXW0I/oaocHpTP5lVoYaEYeTPVdohKzVWsls5sOrgOrhV0YbmxPEtF3eWrg
IQsZYHJQdKzMv/jd8AbnEps8iGyIcJUz52MNfOQnqqWXpyC6gNPxrLKkQWL1r64U
nZzvxSlnYkVZMJ+CearYvZd4TaKr9fVIXazn/Zgc4nNk8aDSdp10hoXYsAWENHXN
E1ZFm3EjJhlAuDuVFEHmtVVdRIHvfP3l7aaizvS6+95O7cG4DZvJnyERWr5Z1lLV
hIA9m27PAhJOj9ZSzs4iULdCfy6iKvDkEAE4n9kytdn7gz7yLicSTRLbQAB0OYRx
oVW/tKZ5Hpl6t2C8sDV/VP8++GP2PIKeGA0MCB0qVe6hk1B85tbNuoYTK/MDjjcZ
++6R460FRNLhv8ZhapBFPe2RxDLz2PYQack9Wr//OWRPY+6uhiFZtFDN5aqBXxR/
kpJSW7qBkSndTfz0wnxvzyCXGMwU5OHKF7+zQOWUKaoVORlejPJ5Hh3kDWw92ULc
kbvhNSwZ+lYMKMP3wa9mPf/GS2qjqs8V4m1AsChs79Q+Sd4p/6V3Vwd7VzKuqX4z
3YF1YNz6bGty3fxgzruITHPG1HEPh4CDzlAmMdvZchz+0EriWivkmvI73NoSa16o
Q3G4zpRvlX1lG3vWHTwXBlVNxerKtWsaUffuOXQ10YAZwdElUApkhhKFVSndwRT7
1IG/4JfwuT5jYlcrQU7Xn88tROYI3cZ5p+jqY0UIjOVe9A5AIdFI2+xCm4kUUYUM
2VeRoG+t5J5QjUPqjfWOK6lGVx+NTKVoDyHtAsRf3tNNs4Xuj6Nakma0swjC5WBN
qeiCvV73ffngklucja5kFXYvky25TrnkASVnPJUsVnAdHeFYwAQSRMnurblq3dw9
yuQn3QhEbVUcBfnJZxaBmVuwpzuiOgHvdjMiqof3P/tle7sY//thm4Dh43xz/D6n
HoaryXQU/SBAlQarqc5fBxEW1Ru9bObSMpBXHCJ19IhjgeFTCtnskWruFZaYHocW
lkb1+rTNxE/k3SElJULlN8hvU55tUWo32ZSFiljpbs44bDwe1eWfC5iZCt+zyYHD
P6uc2HAemgVfRw0mc7BPO5t3EfJjr1dy4qFrOolqRZEGQ+nNc4JpV7SjzEFRD6Fk
EMkX+lW2LTFlglNVbOsPKmdIBkz4wGK+DNoYQ7NRWFrphBkl6+Qy3krWCJrupnlC
/4J7eptKJwolHlqOp7/lGGiI2Af/PdsLXy9Rlky5gtH6SgRcG9MosIt9Uu/LxHEn
cmgv66faPAMpxW+bJNGNX5WM6KxK8L5T3Bm8o6jNISs4SW4kjSfxKJR1Ikgl0BfD
H191Lsd8YMsvn25EN0B53QL6kFfWKwBgl2QugEhhmsJLQ615Jv/bhCe93WC+iRmS
ZKRapRGIVZOFTbOrR7rw+Ynv7RaR06SHqfGoD+rEf4KD4MHq0LweUYQe6S8Kv/Gm
uMZbuHs8+0gIw6ETgRnEA3/LdUvScFBWsXDja5OfNc0ufbh+0TBAllkcW6Ji65Wr
6V20GwqSz0LX583hAfvJlSB5P7T1G88dsvvFRZW/ugClHftErgAW6uCPzmP1DLLZ
I5QtrnnCKvMRxuhpP9tLNljJuqNA9UzKIA/wy0+DO7e80/34XeCoviRjlXTm+21f
BZwABOLAXFJNgP71nV2+Csv2/iMlsZIXFH97KDSv26PgxczC4GLHLBHv2884wEih
yLNgGk3FWbo680rRqt5h7vNXjiAjM3GR92qV4FSpQQiD9E7aWuU0w6bujHqdT9PL
l5cvB6yKocyCykCntn4ZEljFnBak/CvuLxOFey0AGagrs5kpiec32MFDzP3dZGUU
pN18sZGNouy1E/NNgmsi+2ZS/EGH3qrElyyDCNUkoMFLr2VUj3Y35NCLx795QKt3
2EvWXzCoB3oyZFL06J6lMRYvckkgFLUF4+f/wO7XzmW2x1jfcWxd8CH9T1cvNAu0
k6g6xx90Yfms1gZ02ui2IAqQWGckjL4AfLemNYSsTdaAPswz5QBACgYux+IUVNn+
n2UOKRGMbNeJTXrPt4gGxLtU3kTQ4NuI4WMR3A4ywXy9vrETrwc0HkABBFCAOt+d
cIt1Y3P8KmMTTKdXEHYX96YR64e9yGNz59EnT24ybRHTEa9xOx1HGpazL/uSjpJX
+c+HduSFfVIwyRVb8XiomHpcrmGpMNJ+BpbJfbkJUee7xSA2hey10yf0Kd0R8YY3
rTOCuuNStod7UaHPNyJxd5RU7wDJZ+K3IBbXM+nz/WsnOzVBMJEUpx451N5fQV4N
noZW1vaU1Rmgd1ZkkG3Y88UCyRcq78f6c7sQUTfY3EG7GTqbYafj+rz1gWWkk/vl
OUeb7GBYRr8v1RXz3JCaPHlaxpZzWFLTzuu9EHzH/c+4p7D31X7c3MnTBg+uiAFc
kQUNOtc9uiN0epTVMfzYIzyCnwZRngIYvM0H5btshEC0QAni8xgv5+o83fHthbNx
LwOEgnzdnkdl7eMOAObOpMan6YeR+4mPqyg9nYtU+aRySC42cqC5CJ7Z34ewtoT7
iL4qU1AwlYAQYB4lcRTeWzXQ30qp5FXWu8TnzPD/WvuLXBUZN2kBKhhJYQUlITNj
+Bks+tVDvyiRrzxQTu618s2gkvf+LHQ7v8ioLoxd7eMdTcbvCyyJU/K44myD7GDk
BNJB3P/wTd2KZ2otTv81KiVMySK0XF8D0eMfuZQBdwYHqCR/u5HOzH5B7/sXTfFS
vjmaf88Q0yuqywZpVCsq1wTw9dct8iC1PVtcwpwZiyA/3i1hJBsEJXyDaDDGnE44
m+QAupgRIjHIwTWRIInupZXR1ZgOd/h+H1jbG9gal6p905yXlPCgAPsn2nS+ULux
XqWSEtGl4CqmNSClTKwhgnkz8e6larg7K5EI6Zd6D+EBxoc/Y2dVkrmR23EeMdhz
VoIGyqAvKpid6XiVK8WoPNvGHFcWPQOQzOw71iKFy685pkQYjpNjNbZnJhWZX/cd
k+pAaQppWsXG5Ew9zH29cPWxf2GwokdKhDarrRYeI5Z2SbjGwlb+32G0pIBTw99P
eBayAVGFzaSGr33pruhqv9E3h3uIR7dSoA4XdW3MBG5J7DDBUuHvCZHk+0hSFAFu
rs3+LAriY4Qf8nlwA1uaSUUMTfXR+VDmLh7/3MWVIzTVkEb/9MLmFZ89T5qNuc+a
1gp9sX3cyMisjUh0g3JMSljBMkcuDSVBxDBflgGc4gw07td4Os0AZORbZNtVuenR
CxvUe+fbpZR2SdJ2WQo+cI21zwrGHtAM1APXwKf3yoWZURfpuXUYj/jf6ue2X80N
QnFVI/H+cdbioFRHnJVpVy1CQl8mzl1Ze5UrN4MPG0uEC0hRwN3jhg1yuUKo0lgB
GRrYYWVTxHf9U5R8OgZdZbILbRIGg8QR2H4U3P3gioH6Cki1JBHlubkUVeWC9mgY
74f8a841xCXi1aFxEWksBzUfrXk4S32gZAKN+hKOyuLR7CCfL4eIC+nVWjTJH6QV
crC31Oh62EAjf24s1zgsgBNrrzanTgaRpqwY9xNnx9blfnmPgt7Hvmqle0//r6OL
h/e7dIH0J6Yd6eXASCTT+wdao//moNkF2bKM9mvugojiT+bz7L9aYeunt6PEAiIL
jIIDBWZpeFL5w015FAqMH0GN1vkSx1AJUbMNJg9923SuWBPUc7oRu+VtHYn9EAAq
Ehewd91PBZcdHuap7Uut2HGfCcqTIjxOoAHRbNlXZlBzwVKef0S66VuyfPCAHO5E
8OWkJG4+NSKOwjna4vY/k1WPV/XU4qxiE5pezQWM18vDDVpckaYtcuiCGMcfH7tS
tfug5hYCwXnG3CKDPImPTFyC4XVHSWSwvq0KrJo1Ie/pEDrkCeYOezPevkiVA270
VA5EtUmnnwBiZ2NpBNB1VXvZ+8yhJUMWr+/wNnwXjZ8/K8kXE3i6LB+TiXiq3XXb
b78KyuLsHao/wDvW6wj3qI7g7fdeSzPzWR7Vs1TC8rP3qO+fwt6B+WG9GrO4D42h
XrREJuRZPDI0N7jhliAxMvWJXkXlVeXwU4eYYAlN458Vu6HCcSspOQ2+njKzr9+n
Eh0uzhoCR/2VP4pcuab4hpj/kWFPWbSV/MFFcxW/hF3kvBlZsQhIc/vtkvbLKrw6
NQROeCYN2iWHLZraJHUhTg/0ER/WbuOZ2naJEZIJzQuudnhBZG4VyQ3vY/xH8Joj
IoiILSvTIgSgqKlwBOSOnH9MuvPoAA84fuW5B32SzvAoTFDOhAP4FTA8FmVecvy+
AbxdCAuqp5OCLMaFuP+rUUCsZ3dsydlEIUnUBwcLYWFTiqUgUqKFQObIUfQZtrfu
jw6T9ImENm2OJU7K/0mwYUMUhTp4vrKR8EeqHwj7C1qHPANtPVTSLcsdLgVyWnq0
XISvnSeJ6zahwspJctGPtIVGIpa6+URDzD17Q0loFuS/EDqKRnzcMcZKu5aoY5ml
1D2oodydPd8r5YaMIdJ82Wmk04Vb7srWyIobh0nRCsZWXQe3kD7oxNnjdBJnjrft
4DTHuL1tiprZTiNl1fKJ64E88pu5qvH12TTekkQOUk+v+Lrv1yEu1tc3sPn+BLfQ
Z+e/q8MsxBXm6EeecLrnrOb2MGp5DP59+JLuRiGXd+/a49Wf9QAoKvtWHjiC8fhL
k5iMtEP3qqGFDOMQktTtcB3bpB7epLGJE7nqjSs29gQXJzJtNZXoHhwlqi4q5PRv
UU1GkjhZmb7DXlKa5bzmWS6k8RamUv7shM6+yNUnondbxO2sEdR33nPFeoXWK80c
ymxWTlwpow+8CkLGoH9UtcLUdhTE68GKGPB1mnPzbgvqzX39b2lByIPRG8mBEx/f
bwKw//GZ+Q+D/IMBdKSnLpLobjBfzu3yiesJnMAV6sDRs7mKyPk4k3xb3qY2/SDT
lirWT2BSzKmm1wSzYAT5IDiT3+xuvPgRmK727WBsxGIXOkvWWOl0t53mf6OLJGyG
Lei9ZdGgzMXyyfoajjdOjEZM5Zv4ToNWCsHwBUYmhjI0hX/ak03N935RiOyNcEwP
YfVVw/sMdoqBNKKX4Db8LfvaJ7Etz/q0YPT0V4o6p1BrVt1G1bqGSGUamaj831dp
cuNURruo3mFZdObUYIMX5g6uRfcF+Jbwzm/j0BS4XRLwyulPjlRIyB0mgzNrNjGf
Fc8phCc5KFPHFR8Nn/7OQXkjm+mWrNVtOfBfH+DrLDuykBtH2ps5ZwMEOOGTxpuI
u6yhXqCY254XjFK+sJhBL1UDyk6NJ44Lw/d7JmzSuScnI59XSvwqWRv2pwGMT+/x
UkK+Z4bSlucJByFU/1BgetjHDiNn4X6yjYCEUMUy1cMD3QkqiaPMMQcbZ9dNLHGB
LbkHDePBW2gLmHZ2hF8iidGudU6xAdIXBy8C9I5Lm9U7osqbzVsIGiB/ZIl0xgtT
sZ/ruvVs6nJDJnKbv1IXCf2hDSxttKjQQmmjNoj5bqET0awm0nJFjixQVGJrvXdO
7q64Ph/o0qjkZ6g9Jd+Uq7ewE6/PFpJI6fjAwu5Xbj5ti2XQgFNJW4mr2ymzkS8B
7ZNQrpYlkbokUjpy6OZwhLhZXUYsQmQgkNSAP247zu+fOxeCdf1lJZRd6Gc6MGMi
Brk3Ey9WMXkcU1IjXe0jMhCQMiOTUSKLWVNWpYWHzjBNpMQJm3yxZEPstSGoZ7Gp
t9xeH5MCgUpjh6zKfbmUQcooLu02h9x5DFgC9VlF33eJQ0hxJ+iE+oCra/i4AwY2
xDdGOIkFRaeh4x34OzdJ7SkQ199GRV+jmvxx90hb0xqZ5zoNBUK+Vxx9JPYK9BW6
YZRem3jCqThU7/uMBc54/BLmZjVOh5ELmvWWKX9sAMYys6P/U9u9hpbGe6deWZEb
C3CHIlLsO8rV7Opjo8NTXrlDb8sZwiRRkBnoJ8DXRS4f9/D3/cZmi/qAVtseQf08
MbQJ5rFqSmbyiJ5x78WaqLhkLqk4MtwKpxq+/0ipA81H7i5g2TLV8OlgYlOkcId6
XbVQOCXCXrJyQ9jHG74YcRJT/s+grIvGG+jPdjoPLOCdTCWJ6D1DqU1e650qAQRi
XjO/ZZK7g18VztlQNRFDNkNbnyvry6PvgdJZ8cN3d8Hzp0vIzteO1e6c8lTUX+a1
6HdkkDRRImJ58SsJM3gDvqmxK78zj/X53P1tQvggSFm4wJO+3D4gCso2MmDC1gb4
UjHFR2LysnIcEhtS3N6Ss9HHrDmzcHVjQ/mDTiNZFLTcB2btMUqvedjTxp9N0SKO
eem5YFHoHfuAN2odya3A59nHWDIc1C9K/CLa03QhGuMqLgzZF9PuUFS9jpDSjQC0
2TH7TliO4dC7247bXNVfF47ScXUgxKDYjA2ixQm67Fqdo5CF3l7j6nAjgFdPyD+3
en62PQlcaxCPSzdbgXAaWlXOWSJ6YJ5Hxp41slNmTwZJhsha9N+m/ux51Tbq6OPK
mLlJHAWhbOhUx8ZN7QG6CXBUZ13NwvNAHGYOaeBzm6aKfGmZGD6HdG4UcawaF0d/
m8CQYjlouvpJktpi8hAsFoCXtaIP7f/Z8mgA0cOE3jpx/TW7f22AhtFRPRlle4Bv
k7MxgTENR+i3oTSO64V0za394CvCCcE1LCqcJJkLc3hWftmBxuBh7ye2yFicJwKw
Vk5fConA142OJryE5B8X4RcBLTY7ruNbi3MJRYsHwwG8mdkhpbyY0C32lkZJMvpF
YOsbsXOjyuBCJ62Q5bBJLKZUQp5s6mlU/HCgwwYEFKnwlq1ZzgrL/usNQgo/2vh3
c6o+oqGfv/XcgGlaezu4nvEtiwmIv04FiCbrxdT5U8RTMtzWAXbp4wkTrNM3SjKB
+5TC/hRI91pqpePjmjP5UCJt2QJW+ein/5alEBYh5hVKfIghT68Su1NORrDOvUqI
bpyqQ9BVRpZL9PeeCpRKmXFnztZkM+944Ku2lYhI8kDqCNeJZae0UZHs23mn91e8
YYj/9KtAbwwRibrPoqq5i1yeSIxpEpoqBi8q0vA/JgRV3/0ex2VD3d3tHVwCFw98
+6uqf1ABc6Fp7644L6g1smbfDvk9F4hOm5ZlFXkduhSx7aEW8PSzve/xnQyxuhB8
XqdV4/re+bZqDDjLtZifyPAKt1B6J+8JI1o1GUJSqerIng83Y32qf9SNcjjK/BbV
UpnSItezayWBXgX0vF2tlLEt/qEsOT3rNffkq5wy2rXFpLMkRnP2byiJmeA9uJim
zDalAqJ2kdz+dhfbzGwJAUrHKtzkQ+G98rLCkF1KqjRqDbdM+Nta14IsPuDhMulM
YmbD4ztqWUJesOXdHlWefv+0bs7q7mefOOrh0S9EQJefBqPRfEBEiD59phTlz3vB
0cPByl564uQ5EN/9L6/n8ICfGt6KEBrzA8jGZrel9QF+eL8gv0NHlGI+K6PcpQRs
OWyNrWYgShOlIqQ4TX7JgGsXzjV6pM+hGPU2p469qDFVe43K8LYRYbMptW2V6zmv
omLadlSUDXscKRAo4ZIhCkifdIMLgh3As1299bgRU66/2xjKXKz7DlX7fZLuuZWZ
kkbEjsWtgbUIHVYYdxpZJZjAE5Oz38gmgmEqMKhGtpLL6Kn53IPOmEfgIQD09WG1
/BJ/4wf0KCqKpc0qbzSzh9dCXmcWvqbhobX39ISKhgqzbL+R8H/Y8wIP00dXvbHP
pgQmpcAaYKiurGzzNzMlmkwzTxChAI6/D7ynPcUruGBWDAVpznW+CljdHe4qOXWt
x+fqX/MEKLkalep9eiU+EIRyHPX6okhy8H5DLryK8jxXMPgp8AHoVsGC4arpwm2t
UydU6VnHM63Hytr8IjJ0Hgu6Vu/jRHOjiZSkWkRHczyPg4ze/4DjOsDcUk5DvyL2
kwvNIU7vREIBSaAN1PFJvLkbe54qIsDkDbsrvclKp70PuIH+EDVBigzmQ8XAzcy/
Tb/P1EBzRc3REpWW453o1/T99756S8Ptc/0ks0i3xUiRmMqMIyW4NpbbV5RTQkd4
2/kA/Xva3j339FextMzukhaZ2ZCNvFXOuNIlISNr5yygFEApF9eOSXvrdYko2Px9
kpmronp4TkH6fQtbJZPthdV1ix/menhN4zemufBrJZTGWge3F+CI5AdAJSuTOcqg
3gaboZfJEO8XBPeXxmh639TsB8eFGkyXuJRBLYuNv9qRsQ9IO4V9m4Q2AxHS51VN
hCYctSQuOG6e/bWD9YcPhhmcElXlas+zn21gx4kH264ItBmo0sPs3pR3pz5JaN/D
89KLJXzWTw27D2WNyx6zAl1lkxJDu1stZiZQFbCrVRzmWQmktExCzbZqbEamkxTW
bOo0gttOj5V+JU+StdiI65tLLvQvvycm3UdkeZx/9x6lda34lE1CM/513K1jO62b
4GH4Pq1LOnCH/5o0upThp8OnLJmNJfUfer/iD/Ekx+E7rA9VZ/cetES+iOKaxFJ4
MdSHOH2JknNRTXJPyho0+VyfJ4JOgMlhmk09o0bQ1k6Ik+/wiKvdgGIw6aneBcUC
TojOjuP9aNyU3V+imeA9haq2c5DgnFHmpWBKornknjI/DgytMtIiD5e4QeVPEAA8
6gXO29OKUAQthNHERTvSIZF7RjM+MqtLbOoeWwTvv3NUzho6m+Bt+gibgbBDJitf
WuA572u0duHhyih0s8H3CVSdH7CuGQ5ms50U4eAXQixLB8pSQGpwUVxtJBxwL6Bc
ml59PQ+fmrnU+qWVIIbu7qJooKa1pCS5oAXDgtZtXEhhrbzTLzh3RRxqPFdJlUp8
4PpaHCDRGke0bpdvQLd6k3EaLBecNJEp8qW25lp7iZklekVvCmI3nYq/sLE7lTyH
t6mSoCWB6dyO6EijNIRYZRiN9kDgE1ZmzZudkC6uJvZ6fVsVQ5N8Nv7c3VNeS4d8
XYmry6kgldh+R34K0GLnoMBhvptcX1gajXVKgGbrWlEPoV8Jl4I/20WDXVD3xypL
wSpSCBPh6mi0Bw72h5kCLFVDYbsq5EYjbWrCp3z6pI55MRDGPgd67v6qGhLv/YX3
fbE/P5R5uZT476AO5LYeePLSvLA/n84JHzgmgZzKe3uP8fJEzDjZRn/qZbKyczIa
su8B83esSh5kUu4rLpZCtSXjtoIZVn/Tl0zZbOJUGTWWucyFVAsGM9FLbJkDfZQJ
/NSyZsoPtkPmNrvW+G0bfyipFNl53q00XeQNom6GECqGhn3A2FMEtkZe1C85IFT7
3YO1efiICHtnk/SfOLHrhegA+I3L9jei1tO+RGAcGBYSjKY3Ev2oGMRaH0Qr0l0h
3Qu73QUSgaXmf1l7Gmi/IS5/7++TU0OhvOsBbX9j8cUPHVd7im64PV34QsOCsaj1
s4r2UZ2TrzRs4Yhq1WMJquZx4cUT7flRB5woAYX+TDPLxrr0uIGTr3J0W/sf8ua2
civPhYmeQ+T20OlKup2iloB9y9PYbm5LNoo/6WjQ4Efkou7OPhjcvow2DqPJUbPm
HCya1OuRZPxCQ43Ii1m9xA045WW0uYHTYlEVTY4M0w7xhv7aFUmW/WUJLI7L94rN
tm7C5Td3SWRK6r4HHqcCU/xyJ1p9q5r85ufkDQX4rycWBuYzjVhqooB7Tvpt4esb
qgsIC6bktEi0quX1YX2jDxyyYTlRsxWLqIRZhQVvn5roC086Fkpg1FYOmkI2EHja
teiNUC5txSE8xEfEZaFTMxpS46rrpj46r7IK2Z2vPaZaTaSWEJG4e307iWdZL+0S
c4KOa7hXgRv1SicvSUeg9Et7lNKuYEbb7hZorZXCuTGBKeGbRHNcoofLwE2hmszu
JgNnSZTvyQaXJU4djMHLW9igsA3iRNGQEnf2joXT1j1c2lYrEVLPD63kMdnq0BMy
r8XhkNvDFn650WczFozALxul2ACQXC+F7kQZSljGAAoJ2bheEAhvwEZZyLSoahxj
/FoiyEnA6/y+c5fzjqk+h3FeKvkAqphiwvAFrskaswNnBwqlVsgb/NiTuJZLaX8s
hs9FQtp+7EMwYtPC6+NYPmwRSC695ffU1BN2KW3X1mIpTukl6y0cCpCbOxkLT/1E
z4kgmAq2Tr8nHqnaIAuOvlZgaaALQhb2ach1ochL452TIWljR83+PQl4ebF9L0cA
KpE2orEFzf7wQvXr25XUzHFmgD50szuLNr2fTBLkueOzuIq80qzrZ4DGk5SZjJT9
sHHhhlhI+bRv2Rnhn0rToTIGX2sdbERBQUGKe85C60m6XVZP11YtlBVYe6OW2KrS
To3qCCy0AqU0RjvO9ho/QFP7fqtAU3AtLokB5ndVTXe59LxM2Ek2yX68poqLba4b
2Y4RDHllS9bbGdyBrHyJEgQnWMv1t5Qn9i4sa7t57klTOKx+6MYT73jAeDra7gD2
JaeubDsd1lryLfuOGLvx/HN5Ol+V07F/4s6NalH0g2aRnoSEITD8thKSQFoj0bJq
f+FMgGffDwDot8ViX3kDGnJbqBBAgDFtkx89Pa+F28uCo8FK1ffj5hNxqEOv5vVs
eUtkih0HDAdYpJgCKoaLarj5wDUrzvfL8pwAsX+wgCNGYQNXHHeeUavJhVc448AJ
+U+vUdYUyoPHu8Dbcdw8HS3Sk3bKkhnndZr3MgqOnLT7v/k3723UFpFvfIZJdXv/
i+vkvFERxmsYIgOMP5st59fDG2zjYGtSST3z5Qwv327Je+HooSBhGxY1T6EeQYHv
bQKFNAxCtrdm+vTSkUA+s65kqdGy38a+ZF74yDi+tE/hfs5bwtVXVHFmGPxLbcPK
9nBGROH7rtYufTqWz9n5e1ZW/z0yfFwWqGQGet9IpBq0+8soctyEpB7IMZZ5lw1Y
/uR/UOmu2DpTVXoa1UW/VuTHGvqjRsaOJjeKR3J9hfqJt5cx6WAWQntVVHYTowbW
z3/3v6m2IwK8QxtPleFYGbpgjdyuuLOgIB3DyknB7cd9lQ0fmYRJ2TfC7/kN+UCz
Lec+ZAci5Xo8XobE5vXA9ccTPmp6hTIIDq8jwnmDWslCFPo/S/OVe8wOnAd8Mbrf
VN1cxBYxAsTfN8kxteSgr4NAHQCAZM6P2cgceVLZvbacZZZUA+uZhtaVT2MBcwE4
5bMC5a+1CtjH5bEF7mmOiJezseIHa6D3Q62iJ4zlegI/gxTKd5T5g8s7zx8THLKh
ZWftoQwVPtxhmfzl9nAcF7FctN24P7p34/eW7TIJiPoZSuR3TwEt9LIGF4mEEhke
OgG2xsnihZg3oJN6ygF4ccBmmE/8cGuAh9BHPy25uTI1S8a9bgZgUcPL7zsg1wBk
a750o2zOsoj7pg97L0T+E5VT9H9U9Q9myXALB04E5YjgpvSq+46IF2l/DamZD40i
XeZgT4gS5+8xgT/o+EktJzKZI2nqDI/KiRJZfERdQkji5hJ7JwBJspfLMOlSknf8
acBHF1WlZKEPh5TaUAlrZqiigIRMnGA0iDMa4TVA9+xNjGjBO8ICccjNHNnO73zV
HXKhy3zuxAgYDnzKyAlUTrANX92Wc4e6hhL/ZZICFx+i6UE5woYWRhp+H6Asb/4F
9/SUSWNOA/uHhsHvdZO97U+8CkZ4MmXllDHwdDMh6CGG16lZaxdpxvfkyiNalUeh
CoDNqPj0fm+KElZKNkS1HNQkMMMbY75T+GUjTe0K6lXsKTU5qFV4wXtV53jtGFz8
1K4F/S8QqXbM+Ohstd4zDw+piI/Rcz7JbdRLhld8Y6P5cMWecRKaLhuO4r2mDWpy
BcWib+v5MJr4b6SUB5QLtY4/RSnqeTQ9uJ3i06PdedtQJsSrYbQ2vy4cTzNL0EZq
pshkxyG/jbOYc14LoEKXDzibqET0bUjXXcFmI6t7xvqPmqLxCrWdzDA1LsN4cWf8
n6VpJbQFoRYv7bynqYP0k3Rlwoqqgs6ylkxWkpBtXqGdE21ivINP+ooieYvMDS1S
mK+V6Rw01BoVARLUA5Z5c08j8JcK4kr14PfbtrgBZLq9VC09vEFps9DXe38ZHJNT
LMHgBKKM23vl2XZh6iz/78XbHYssuAS4bA/EAtoDPVDL+rmuxiuPTVoKiiKp7OFY
7jD0mt4K7gXdTPrjtJEUs0/fKXGkphwHTbYk3RxjWZhmyt6foxWjSfWCmsKpUuSu
vUhXk7/bpBiIA8tH6GtuklgIWSBAPRtvemY1WiJ1O4sUiiqDMNpWjkQlgHvcG81j
PR8zFjsh75+9jcfJomiIfrDDXCq1kNWFUySEkyfJekJbTc0fiVgQd0ZY/uwZPfwZ
rlIj0y695hAyMejvwNLiFGTWtCjANRWaDDijzJI8skoFBib0sZscTJAt2ODh/Oer
T5hseVE34GCDCt3QcrSX8C+1MKnGjJqa1UnvH1YhPUz/PeK30O4cbbzh5R/yIQUt
LkCD+wXSx8kAooIvH5CWpdS9nTcO8kNeDOq26QlniJJnhB6aJAqCKYEUpc1arNvz
/0DphTor9EX4haXyhrXOF9/7XQtmVZOdFLmhEmgVLC4ahBXYmnXluVRlcRYQJIXm
iJ7nsWim7fKIw7KKB6xitbEOYqrVqOTWcnHHUuMmtKn/IW46FgxVUwFrZaecDDt+
xrA12Qjpup+97yABtboIca3UcRhctf4YZqZhQuJgX8sjn9bHA4CE5LqY2V7/6fqO
CAH7B0UvEdFvrND2PVS3Gj5HWhPZpZnEWkJ9W/u847DZ7tEufIPEP8iwjYjaynNg
FLOAPqBVeelvaKc8btQ7xHKIlscY66Gwr8t+K3QNc5AH9jznxOcNXp4lYE6jqOvz
lbKoai4YZext56EIsFoGUOvTirg7ZZzooqQbr7lHjEPMGvc3Tqp+yb/oDbnWpgzY
6csn144oPjY2ck/0MR2pSfeo9mRnqPVfgiWeH2/8DJSEEqKlGjfjvxXw6fDTzEDA
mpnL5jkwE0of/tezK9T+crISewY54fxZE0pHz3MSDpvGo/3QjHGF+ls39pgM34s8
jYy0CgdD0TFc+7avTZQNXWTxVVzduyGvbVEdx28f/Mb8E46VXaMT/fs5Bm/VZ30q
SWKjCt7LBE5mb8kOUXHR9ZzSEmamHsZYjF3Mz2TUz6s+3STEjCQ3XU2I4rbIO+p6
VDf5EZZGjDoMSmZd5BjzC8AK1YgddDRlUhmkaoWJNyqE2x3R+jisoprSjVUC4HDj
r4SUOgkHbAYvXTkeXi4ivETIjG86GMrNMHMtIDAhWZCZbLchox90Sl6z8C9qoPIv
0osMGGBsfT8qHnVUEZSm1hiCnHGOL9Xfy8ck0Ojbtm9Yx6Qa020QoMflcdmt7gC5
T/n8n19d6db76MsRgsZJXmdcdBstBiHW4FDPlfzCCklChXwAofPOa5dD0h8aChSr
q+LfgbxO5h3RSBYsmrGn7Rub9aMyVHt5R8lkVQezxXyhyffppfV6HFE6ZE3Go/8m
j5j1r2Z9IwIAhduncIrnH5bFCn2hpLFogXtdTSGH40/wZfu6fGgLwZKb+VVTDQZG
c/1SI7Q6zpbNRlk1YqwNwd849eCsTwU4a3DUmEnC/A3AwgWj/vuZn+UcyBQjBYNA
A2Hs9uuNS+qfvZ5yhA+dpMBFIzXLHUAx+KLP8wK+aReuKyWYlCTQM2x6+4g/umEB
MnOceHawByNgJcLs39VcpFCd/z2q2qy5mlAhPFo+fCSBpyptQpxI8URoIwZnAGhn
ZZ8P414UzjS7/P+xZTg+N06XyDnkQ6Hevb/WZPt80JBOEmiXpfpbTvN/kOxIamZ8
8wr+c0JR37ynWSBzLm0okkDFx7uPbJlRe10B53qqJJQukxRwut7bKgRtybC6NGJe
a2db3YYYPwdiYmvKslkgDib5L4dTY7gAmuGbrnVTpfUSxnsnf/QhaFptXuhPl2s4
/nq9wZcKk2ds56WjzAisgZJyP+isBuUROGrYCIvI1Y1IrbIV/eQZ6JmDxoSE82t7
6wDqYzl4uggX24NZvV6+BMkSm5L10zMnSyCd4IDTQH+1Ai/OyUFt7SGTlMIP32+p
XO/95yFvJGSvyNe2WRC8iUpx9gTATLqQ0oplYelSfQ+GBfygInBJ3QVHKRueDEEG
/kgUhrOYieOog4ylf+fnqF3KYofZ/LrJtTPfPs+G/yYGrAqJxui7WlwWn5AmO8d9
K5QreIheEzP1s9gEsybYVkbNru95I9R/Ijb6plvb0IiLz5ggkUn7nqYUHyI90KVC
MXnde4qN1uXSGCEJVD5xjHVhOMYr1K/jWk0g8Qf5v7oyap4YUt/oEtePnR2Ya/3e
wzQCrPj5ix7h60O3Z2hJMUgXJWAGeX30lDIbD3yWcFdzRIzCzphqMstuvRPtv3RI
CAsJ1Eo99NJ8I3nNMa9873UieYOMV/Baddx7nv7a9TudsoLCxkTMZqdzgUjV9IOp
svT+NJKx3wymgVvCh4fwZNcsLilNaqoqHSTpCLdYZUPW5WWeyavng98BLxwYXlxL
nBn4FlHUIUDeve0DqH0wtHRswpp7EyE9xHZdOH2dOWrkKW3AJqlEfRxRw3iR2OKI
nvgu53Dj2KHA+8LkAqxvMPO+ej9vWlOlZD0q8d7z/Rp6I2xNoD+qs8TZ3BVWjhyY
TuIJgE+wgB2EtGDeQ9V5zU+JmuRuJcC6uH9098xHTR3xWBnpDnL/zcVKH1yH6fuX
Kera/PKkepCSI+dH3Geffv8zxTtl1qmOOfGbd0ZUdIhGLmr092FpNstJOQj4PqBy
HCR718RtCIhFxtqiLERTcQt4thV6cq0OusfWEEBWfuG8wmyPdIFzFKWNJVWVAzPP
LCEs4cXTwjkp1wanrEsd9pN9QteUwfGh0Ahch01TZMJrtaWRfk35B5s9+fhrhZEK
MXLEsaKFT64+D/pXy0LnazTi+lNLXhbGb5RilXgyho7a8sHDCYfq3dNwQxCzWAWx
ZqVWNl1D53T6F7OFftjs+LYRXO8SvQzSQbr1u2/ekxUS69rYOHDy97BgvK17nrd/
WVsrFun0WurdPaS1txkUO8+bCAN2d9V3CG8ttv+q9p4rpUFqUdGD+FynwgwNeI0/
QjsmtCc87EU55bTf+oid2xVSvrAfkYUbFKutC2D+ZImz+jsjPh7gUVBuy8+Mgy4k
QgonJc9XJaeBP9PV4kIpPXlo9snfie7hk2p35mXWVpyCzCenORmbu2dIOQ7UQXtJ
RLmieBTv7VPG7LOuJfbnaWJjZerlUCTYID+I5FxOdeFg5+kvMPXgeclBXwp9LD+1
cUBgFcw/4Vo2Sp0BRyQ2lFooK1gQkWx7WxHQkwtpYdJicGNquHy+rMTJKlu7YdEw
3DmbLJtipUcpcVvBURBpQEDgoX/FHbRttex1M9yvepAZBHD3Ua9m4C19QOQKHp0y
a5ltCjJe/Sq0ipvCHB78dBwD28QzgU0K96lF8IK7nHjFtlKhOueNQ4ylb3b64Ctd
GJxAW4sLrfEw/E9xUBg5GYuTFHLUWMMHEpvDHienINIeyc9RxiCRkl2VxijMr9f2
aoUYwvGbo1xVMmP6/qkQNWGqAoKzPzmRVn9DRRSUTW6C+cM8ey15tsSvaiKzwOuu
IsvOVOUuLnOQT3MakYPnVPI/+3Fq1brelNGJVYbf89KGuzakTw4bO62gMVehdZnF
UJTeRmIZ5DtsEYYbXjWqffzrDcjXCyC7vwhTYVc9iSPKNp60titw46u8LUkpY7RZ
vjH2QlqVBVvbgxnFnNKyxhCsnUfkYDm+gYbCUetl7o8Xx/yvnTuDpeFF56lpkn06
Oow8xyp+sqPMFiYFk6cdGi5eVtHwMu6Y6qErxQGjxjD+DSoRs7JKM5VXeO5WK9+9
F5c0w3I/5VrBrLCgAk2ub+ld22xDB5gVfSTq7p7g6pKaSEIZz0e9Q7VsppZnSOeh
Tdz32iR6NiG2UfDFG8eS7/5YBDFoP2tA5ZXILNxBGxUQZMuoNybaYPi/m1FjI+0X
4+vnJ91hiV5WDexZf8y9SY2P4mOqqdmCPevBZxUH/iRovVK1GhvQrFf+bEbeCknR
AmrnWLNGe1ifIBYgMo9GAyWZ2auBxPWC4XwI8FKSjpYd9Y9SrkTtsrlJ/gBmtQ/1
bGYdrZ2HVBOtJYJU+xU+kRKXcmdE0UCoqF/OnZ4XDVO4MU1cJa4K69HF7ne++Nrb
0AuTZz9+R+t86igi+L65pQq7gB/wtgKW+VtveiZN0+TVVZq+pD2vXrHjFMzhywoC
iuOcOlgK3dEq2YhTzLmIdxH7/oLcW0msYjbRzbkMD1ERGo0emj284gpxrluLliTu
t3J/WfZihLILj1BiR35TiCZciRPzue1jMQsib2j82TKKNTIILd/bEBmTnqZMUx1r
St7Ibso9LIKblV+w4gXbHHazLdqr5DpDVzpzSDmIjRRJfcRTU88hfhKZxFAv4wZl
w2CZFePcBsKLcjEreTmuTQ8Wq/lqLgnIkGK5a7ISsArpyHWGYNNH4VjjGBTl05qM
4ROoh7PYfsTTd5Cu2FrYmpwi7kmpNUn5UjlF23FcB3/q9QsxX6yBR5sHf3QNiUdb
Ncl2fkJ2dAIX+e7RrTA/IqIyrb3vuXhFoZubhVsBi3wrasyjvcLzIjIcvwlCiB13
fctgf/FQHfieBLCGPY6sbKwc1152Bq4vrvmHg9nEi/KT1qHVXhedTQORSTwT+CP1
ZasFn5A/n6m21lhJ31HtT2k5SZApFmruB4L1VfOryyNZuxbSTrW1AiktxuFBE4YM
YZAc5CFwwWnm+LEEeUVBcDM6tTXukWfKKXAl912sb6acmTRoQcje8bJ+swOQNirC
1HfFXh0+nF4l/Uq3rQVdXjwGng77hKLS4vM6yKYyFeppFCGZj/ML/dUJ2anPJlii
d0Z9iwSdoJSD9AoYBg/RGECWrFG+Vx4oqOFLHRLVsm5RXCKvT+qfHsjv7WEJb9DK
jx/d9Ni/iebsbdmBeAnRsE6Tm5wpXqM1Ktryn0SDQk2j7FeKUiLzMYupDU6Ujpvv
/j2hEM5KCAcVQUxTgmxJ3zV64nU2/91T034OYwyLcxEfN9T3UrdHqxOqnPzNw7cU
PNBdyr3Ftg0/WYCXaxB/TgSv8knxA2e1UDIG41Xffa2qLKAHrakmTom2HEGVIRsD
N2BXkZL4oFMICwieglI0xpUFs6XCpSgEDFAEjKqWySkUmWgNwns7wEr+/C+/JE8N
Co1zYlo/fbdzMPZUTe9Kvtd5bwzOKqnq2p3Iv82fGlmk192Tn1JbvPe3GvCLLx46
ARIOTraPld25O5QIgwN5UHn16fd135SC/SZWCnS8eRc5uFit4qLOcMf1wncoEHDQ
AlrPjoWHWZjBgag26s3ms8/FpcY7v9wcU/N6jbQ+YphDSFm/rMU2YQF1/5hQ4lfL
EejbLXrxuXSvS/uP0SLuaEEYu3riP/2jfGSJnRYAvAk2TW9JXs7LsQtXUEz7vQvt
gzYqE/UN56gyeQby6HWmKcamhFdlls8Fb6OkHmzRT2tjp/h/MPI+YTHMO8/2wDtH
0tHwOfttUefOMfCIB0Hpq65hoveR1iGjr1zWpfKQz+Swj3UeTnBFHFgXW/ykXAU5
J206UVBQ+OEdae1bFP7uspAx9iBNKGd/n4SCL9GCe4xexBkqNSx3Damh4NZ34zgV
QmEDgLFqUM0JhT7Q6Nw4aJohK1bLo5aqvcNkH6Sy0U6d1qdxKwXeY7BZoRflnx2b
nGMht3SXaQM346oL60OZujZSrnFtVmUWMRcfrJYgU9f9rpf+sc17YYojHMVHz93V
9Iquv/UthFGwIVpZUuNtDWlCpsMftg1QrzoXVYUFD0gzple0PV8E1PVDC1O4+aoX
IM9SSiaOENM2ufZ8AfyS2n4iPkU5GXFJ9XFWtD4jtsZ4EIl4kmNEFgHsBZb7hXx5
6BUr6xzVLaP5G2D09FpPp36lCPAUk0Rklhd54gw8JRg8SrROollogrk8l7DEQADI
zOM9oFvLL4i43AiynXZHrV2P+SzZ0K6Clwmk8NDEMKkBskO55sos4fxgSg60IAKt
0pAFWeX8YyGjlY9fZK+GEb2xGUlRAfffeaje/kF54vnNEWfqnIKZnQAMU5yfB3P5
z92jfaVl0RBkDxMQ1Guh2vw/euYRN/YUEenVOIAzkQGww7V0rF5DeGcxopnYVojy
iAw2HXZANpSm/QchgKiRGUfZE2CXndoHKfE+YalF5duNReWCE+faqVMsFlItxH0j
svt3nBjdWQQmoZVu1o5cLWDt7fbTLlZjQ4Igmd+ibXAfsrLPH4NpD2B04Kc9uiuI
fUqpyeTMJ8L2yWK6X9cy5G/UitcNbUZeXzP7mhvJXQT27bLwngTc3HQnEzXcRxRq
ZcWkJlSsna76r0LZT1mNIGkyEsiX1oPChAD+H1maXPmbVwBwB7Ab9mC9yKwOmFV2
CRjTjqM1pDxDvZx+gQmwSjkZfVBjbw7+cVttGqd02MrNbwIQ9PSSmzmfQZi52pSO
SZTTgGZwj/njDlef82HVajMtnNiF7aQGiSpJUy2WXqSWShe6U6KGfPTLTPzVL9dq
9THqHQJJLojZrtZggjmPXH647Dxv4l2fYL8hasVdYAeW1GAtdqLWu9X4hn+8QvBB
ds09fguG7MDtKVAdC6KpH1KqBMWz/RxK5h/ZpGgv4xZtDkhcBKd6j/tTap4zU1Gf
dW7cgLCiwDbgWNojjJRP1BXJx2iMDQuztm8NslYoMyMA/XUxf7SLxGSXeXk+fK6S
gV05iotqKE7CBKPqcYGseXPZw73hjt68KXjLzXTj0v2Gt5jNmbFP27XvTEFKZRyU
DxIEMWjWuXtHCO3Hu4AG9AwjCss/MQKWO6hGqrNrPejAE9lfk9pfvCRGpAK04gEd
dUdDMeEXjb9KWy9tLYUUca7HhifvprJ3eI5ZgWW1ag+Hfni7BV0eK+r14sQj+DH3
+rHwzLzY4WCC9IrnfiqZ+YcnkuTG0AaWn+Mnafyh7N19FvQBMsO3+u0Libmuz+PF
Ic7Y0O34V86Tv7lgxf5ho/ndVnVJBNOws8SjpzCGS+eVy37XksAX6qmef5SraeQn
Q8Bp4Z+QPKYaiwjeUZRUOWJO4k8wWQKNalI8sGvogYytu8sRda7MyasIf6ZQhSCb
x4zs0rkxUsCMJl/V9DjpHiKhkj1igLL5Q/QSXVaK3x+tWRfoC/gM14h5sdTsKZtc
YKtS8fj9xv6RigWybSFSF/+EWB2HH6/HvAVAEhHiG2Ai51iQsvI/t7k9lj/8rdBE
VDRvYx6GegP6G4B2ik9skTVBeK9kijBhc1TmLnwV5BgtbhAPqTjX2fairXeRE8TQ
aNPanXqV5M1wDpTHNgfqtdAQH1lRSCMYOozt9Svohu6y8+n16AIYLs0TiZTVPN83
qSlaNynKN4I1hodZSkpxQiIO8fiOejbeu/gHcMSGEbXeK8SdsfzyjXcFvg2vR3cr
9a3AxZIBLN1oo4j7MW2dATr0LdsOJ/NP7YpOUX1swQqQbJ+3GaH2xWKqe79N2kO3
m+lSqSQujTAHoFMc3hu0rhVtUmBMI7izbbUk+q4DxZu3vLSVWvcqNFizrhRL02BK
1lH+02zCdvNrz0WYNs9M/grscFPlpu04wjBqWpQp2jww4U8npEibal4/9dvtIk/S
DQk+eQd/yJlZZKuII68LSxxef2RvhBON0AElblvG4P6Gt36ruvsBLe49D5Ydz//C
FFENJPolWonuULYYcnwyyFYd143rWs/jRMLWZUcadh2CWvYzivnihi6xQhyan/SH
8i6e5/zruOmltBmrUauCnLeehXie1lhzd5FIX/AJ7LKnt3uvgL+YowEId3Op0MPt
Y1VCLiAO5Q5aIIMjxu2ZeDnkuSVwQsyt/e19d+TzOOyGW0bVEdT01V6xTbFfuu/S
4LvzEV1a0aNLvV2l+bLlrpXgMI2YTUXWU8+UXs3rvSweO7XZqieJ9bgC760sSieg
r0nEzPGLGxJnIlFlKucAJZnfXeYT1mzHmBDn0pR8WDBhyLkHdLxfX18qf1JzbyD0
dxLO8h+PpnyyWG1rLXItsLQaIUD/eJWhYxJI7pTMwzt7atTMdy2cmqvEXalKmQRK
n6cg7P9pO8ITxV1fzC87PXKQraZOlWPH/vlTUw3vLujJCV1JiVJs8KBIlVK0y27b
dwBg6/Ov6oEkMMPQpa+nP3wPs7DHykYIIRjAckX/99BGB3L0g3Ak//qB/U8xzMz8
WLXQRbQ0CnDp/LhqbTsgysnFU1MJOEC4x87kYdiw3h+o8Y9ZKlqhcGYTzoN4ES51
B0r6rIfxXEhNfVSXRMuxN6eVcUvXMgQ4HZ+kwC0ordHlng7Ml14Bp8gN1N8Yi4Cd
ssrwsWTQUQ9N7sQGUls1VVsQe4gP872NJpfq7cuK/ZZFpdDOMRyMQSo3dEfMm+sw
+IsZql4dR+TU3JCWrGkmkyN3vwSFjiLZdaMgcZa1Jog55F03IJTKpo7K8OHUMqcc
rncMezMFlN85mzjywokYJf/jngJFkUcqEwXzsWMAQ23OEJIvSNzHCUCgrFrde0aK
pUjOC/8Amg5hBzHV26GIYDeGaDKko5LCnS16NE6MEMe2+xAcc32N6sm/G/pcmHGo
D4GxCdNVmE2FAm1YGD9vyx5auK5uSALfvV4GR+50BE64Mo8lyImsGz0R/iZ+fVbL
Px62QFSDUJcrHbdhjWJmLeoCPBkHYF5cQ9tclC5o8YGYhfKcD1IObSnO9fG8eCx0
WFe7k5Qame0XYEyfr9Mh376ovzHtR9k/tSAhEWlg/IYA26ABnDXuqeX+SJf4QHIQ
mt2ZpetUG8/XbDbxkVsHSnwdlGGE1ar3psuv3WWCvUwJJTtBqPsNaIrDE+5fmFbS
cVx+ykHfItLqYvG+P74Xpd/4Lkx/bWlDzzsnFvltUX+6QOjal/TD5zAeXDhsX/zT
sgQ9lI16LbLqGNpKGx9Ka0r9ZdzXWMiKhr1q0mPLZ+E0BqSKgH/tUz3Mov12i1bK
b0cUg6LCSgai+usX35obDTdK8H0fduTT+eefdhkGw04I9shOaDP4FLRu16J7Hv3u
l3+WOXoyds0Ou2uykPuSt57hLUuLImrCGjwe2Qleni3qC7uJTlRKBNPczd/9Pc/L
k8LLxrU+x5Dif3dBUUjnfgOmSeSJLTJEh8upoZHlxv6G+y8XnkqXTUi6KHD9hnUz
iG+5s1O4I2RHx8PNpUL73HIq7G8ZKIjYu8YI+2yEj28gG08M316QQWZw4/4qxzuO
YZR5BNRPmxtW203HSVRAwsIgNIRcHBMBsrRhOqudOWzrvL+p1Htwnmsn2fo5XfeT
QAa6TGWkj+ZD6oXf7n6wjL9QYEcC36SV9IiYjBaeBQlHJUj3t4HgyxJ94r0/G7OR
vfeS/CMs6azRVK61ZVBhGs8cl58d8iI6uJqNSrcgTjKKugDed9StQwGr1KiWxFZK
Py63Fv4b9KEb851GI2q4s/c2uOCHgn/Yy8bwRb7roy3N71fFAX1MVvZyBqX/yDPq
QEWeqXGkxRrhZ7giTM1F2Km6E3RccI/pSiMYjk/IZ/VTIS5Tknd1TjFy5+4jSZNF
s9+J5Q4s735V9LmJGcyMVtqGUehVfUxur97ApIgVaWi/j/wq/0mNaG+PQUQqEh5t
TOvrAJyYasgMtRsMt6/1bvAYR2YAETgv7PNFROC3XZOoHkkkh9WZspxuChtHIVPK
bKT+/VnjORu/RJWsguJ1+kSLuG0wgLW2yeIp5NKy2RicPxW2vBbMLsKzVg73tho2
gjdTrE/hqqpFCzQsayNVkaAFZTPKn5RsD47NiAnLm57AzKlFy1gIJzgQufVp3j5s
WHmQTkbDEzF6N4sq8lZK7Gbv8E1j6bLmqBTAaBDvtd1a+QRVFuQdM8CM0YnTYOwB
BZulLqM0wmDCuTlEgXmSOW0TI4xqAyh3cq9LtW+l4aZhiway6rYEosue2AfcwsV+
RjAe0O1oYVlonb/nSaSNRmfhvbo9e/UhLS3QVIUZXZeFuWeQuk1yu0qWF1HuKgXb
Is9ywDH4CGtIwHcORUAVPz35ENqQC07UdkPQ/L1Ou9yKjs07Df8lUq8xtTtdmiLg
vp2Dy13MLW4w65iL6LnpKFQHzH72fyp2nRrsvzf2CBuOKJDRwvmfE4IWtKwmHo06
DKjen20Pbcze/MQyfhrJ3afNhzNz+BjfMkeJ3oA7AhKklhfIhXe4cMzZD38BW/58
KvpFa7q5O+WJVPqnB4hwmZmsCo/uv44yAEjY/Y4BnjPjZfXYZBKpIvPFZ/ApriEO
SDDe5hx7AVCgMjjRDpmQC1r3fTvE84PusFfhG+YkYsdSAaoWO7ydsOe8ZOJeKrqS
IppixfVAbFY+vA+6pZE6shtPi5YTa9cyKCI+G6pRzg4wIjXoiJqmdh5qpsBA+8VQ
SRJiX1qgnKkmKoN0mdk1IhDQ/a6eo/zknq6nOhxPWh/AClZaUU4RPi3ghGIyfXvP
tllHRrXU0v1rVkwts8AUfHpbf8PGXtvdx8gCTSXbzx5XwWLNyWaT7dDivrDtQGaC
/3WtSAv/BtAEExBlrHCo6//FomPKiZAnqPfYUxISSuugFoRPqB0iiloloyKMRTyP
h3zlBUBrP/8/yEmuk6Si1diUovTQoIhyFlnL8q68r125njM8jRFODf3SySeDqaoH
FqDNozqVqKr0ZsMeWW3uaXb1nC1/2OMwAG2rjxfBcy9eYibvRUWfZFjSAvM/JCS9
d2hCDFh2FSj+V5XXYaU9YfdkrY7TqoyLwE8ACpYiMaakW1R6nD3kIOVJ7d2sKEx4
c/swnRnH73ATUPTX3NTNod+44RgRUQYbbJeF2NlNNBM7cIMCrBq/BlW6J7YyXL9U
B2F6xlxL5YrlcQCE+kK7xtpPFFiXDAGEPxSuC3Wv3SAv+i5DmAC/nthVsrid1N3W
2IssxghjkpVuxEaSZcm+QJJxsN7kG4al1QNn/4c+KbbZ9JrNCd2+VkMujMj8ZNd+
SLhr7/kvvdJUnXOX7wS6684k9OYDpaZ1fIynRyTqzeRUiCnCdaikeFO+DBbqwUQW
cDca0bxa42qFOR6zSXjPL4WGH7I2QmMbqcYNz5V+ClEqGqwyKZ2AKSgubuuJVySz
OikB5VHj/07VXoegPlus4FKsnbgpqLT+8mEcdCpJyG+PHuEDFqYNZTe1qdTS9s3A
KYZ/g4TAq/iNhFyAuTjDxCMqmZfwaIjg/JS1h2jrSWZF7xkWXVl4H0asgRJvL4Kd
XJmuM3XKiImQ0NtpJY5InNLK7JICvQzNrU9N7Kqt405RCta7RytjH1APF4kTAmS6
9yW7FSoHDAjAOTHIUtN2FfOBehsGB0jTjanksb0kZRyi62UDGWeNpP4wAOHoo8Gh
w5WcUboJtQ6rjeCTPlgKMWaC1T+J4Uo8yPcbOvoerOmlsqU8ziZ9Ea7I6gPIcFYI
7IPi5HNRNHYWvpaapyII32qZAUE/JJND3ImxbqyYhzmQEGZ/7LjJ00lPqXxNFW7c
dR+8XA2ID+M4T6ISvsiLbaeVbJDHyXsqpNtn9t1vCv0Uxnnj8ZEESTJ1o4mL8+sG
BkjICCDUWWbeW25JaoDvlMxtJB0UkBZT4wUlmfLgYhDvJ6gDdeOAUN1WiWYhC9x7
hX3viTuiWJrHX67896nS9k2D/q0upuSaDJ1Gw484d1C6XT7+/NxfeCX2qNC6ygse
/WIeBrNNHjnhtsjYS7vwKXH9pDfe0gkLzA15D69YLhGpY55SiEHsYmWTDM3fbXCa
hjZifrmfC15J+9VAt4jcs9NFlxaPosI9ahw8UwBzh77JJPhv73fZ/8A+kkYv8HqI
91unddRhxE/8v/yrj5IFNAUo7mE60r70sBfTrT65Pu6v4j+NNliu6VDIBLdkWJgy
WzsYgVWkpF3HSq0HGjtdPog9bO6td668mj/gO1yzGUote8rIvTpPase539G501tQ
F3dHdwfGTmDO/ixt5jmJavPrPlRufUz3NdahMEe6wPZrGI1Lv3YVffwZAV6Uvze/
7c7ACXn7MJVQVdzraEQjmjOz0aWAf+ebP0yTJWCK1Ow3OdGs9iRmoAEiiPejgBxX
4sdpfC+dF+7UzspL9zATtW12WcdUQUPph5R5Y2RVYhChNH8ziHO0Ci1fI1JUkPeZ
rZ39UNQnqi6msvSrJTtWF9sLbhpIvt/M5SmEBzOsxHXcGopRfRuBp8UFFBsmWoQq
6Oz1FlYc5+zJTGWI8QWm4NcWPY0yITNVm+geN+TvJe8JR4CkqO8xRE1U/KJF+cTV
Q1ZGmWTT/EuG1ECQ/r4eWBR0So3cl49edPLMJItsm8TY9euFurKzYIb1R1dHgwjU
+Clo0o5bCsW0OZ5tsR3dxjFJ2f/hikUf2jMdbsWOpUpFCzqyqCbI1s5sYoOVvXep
aJasufq2M1puBx7vk4j3SA9Lv4z2zLhOPlCwnSDA6KBeE8p19gRCIz+/aUPY6dK1
e3swgAijE8NHpS/pl9/4x2bwABF1cnkCOnmCwnCoTpR0PYRahntBFMnNGK+4jYF/
Xr/jDgZ5O+dV8Liww++82UPNANdmGe+Tkq3GHVS6+r2eBgTD0r1k/nce295gM6A5
/P57suQJ+xj/aJxsrt/fK1zIAgGy8/kdTay4mHB++yIJ7jCOzYEc0UGBdRARh+qM
RRxc2u2ky3BKXs7xdJtf8P3k0KZvm4AscfOriog2ccqXy2Dzh6fpO9QZ+DdqS1yQ
8uX3eDJadpFhbXlSjHBvg6p7ksjtx1EqAH/cmiAIKioiq7G2N0r2oyFFtOSdYkJ7
WVyPqAlixB3y6/osv8WlRpP4JzCSeRImJQKWCldsbB3RANKmkZB+snfNp9dho3cX
Nhs4a1UYqosvotvmPVqAknHXUD9PvT3IfFf7JjyACTosyMCR45AjkBcEE3otA5hD
9vki/8G0nDF56O1dnWHSgoXxBlcNNB0g5CTNVJzrglC9C3/7dHzJ52LTBej7w6i0
oEKh6oQ3ZFl0oIjCDwywZ31tJ5yPHN844ZMSgFrnO1uJXMY77U0Ec8MSfhO/SEaT
d623zB7/Ksg8+pUHmePvTMAE3lR+7lerygzl9KKS8VJsF66cqAB2/XpIzrZa5ZCU
TrfhYgTSD65xlIuJBj0ZuuJ8NoYRf16ArGfI0rcXv9HkejH72RDt+J4pxIWze7vq
InDrw/qf7tQv3k4krmhwPj2g+n0VgO5/tGu0kdynx8NqYJm88ApEINfIVolVDl+d
V2m/dh6Tzqlo/syCQNj5CuZyxyKAl6HwcxNcfjNOIJJMgC3hNgfOR8whTjOVns4E
D/gMTcv7/5cYefvqmrj3cxL/NXKXyRFJEVjn6WdKy++pbd4fMdMqrOUGsMjCV/Yu
iFMI3qZgwetHWTVyOn4RyelpWm5Jcir7nle7uArjVpvA0dqSQEz9Jjd9caA4SiVg
eWCX8TnnoXVxwVEz+YRfi6vBDZdgSBcXz8JQzZ3uvn5vcWEiW6glvnmPO7VEdvcP
1fBA49OIwlDHOLI6F669lwhVostLoPo853RH8A4JiHcOBOVIRpDpe5FoZHc9dHZS
qvqcQ5h+9Vvx6qll6BYsHftemyOkdDJYq+jatlBTX1UguC7Y2PBNJ/N8pLnRRwGk
imS5fYV9Ah5+7/CBcP8o/glaknI2lkUKIp0ma9kgV0cZJFwMdJOzoqwpAzd4num7
I0ebQpfBqiJvWdEyze0ZCCL6YSyjkr10e6v9jIxCyldxl+smv9WAyZX81qBYsq+b
w4n3bi/4XEr9caS7d14OFeQqhuQwxtC5p+bRVt742l/o4ur4iwiXi7BfgOd6b9G8
gPMiV4+ghv7RiocZoQw1jmS8GTRo+Pvjb8mwMaphO2WcADTEkzn9cTMPBLXfWwYw
XjBDprVub5KvoMSqzlD4EHJndwTi6nPdSO6mW9LG8IPEuHB73gCWEKhyuK0PBWDI
w/d0MkGT8KGXKpDXIEnd53Y2DvRFvmZDEXgmvi72s44EKn9KFNew7YTMYlKzXEi0
bU5VCkXM4GZ09w/ajX8REL6EiEhXlkF40Z8vvhjyxj4SOtXhbcpuKtzFNTu8bt/+
HkEcocuuV5/t1qPrheSW0c9hIX/CwQZZ2+9xHSF4G99uOaq1GC/YUNpTBsu3DpBn
tu30VZBnklKh1G1BQJAuj/egW915j/aETsS1AEEmC8d9jN4N9DDYbMqDosT51wSt
gCWlv9cHmL7pm12tlFeeqDzdmFhm/+nuBgcVeC+f1isWQkWZqgyhLbaAg1f6iugc
oDxDdKa/7Q8/0gpcET+QZoM12nSPd61o5qJq9T4UgHELpfLrC4d2CoEGcrLIR2CC
YUwGxDPmSE7iywf8GooNQ3HZS8TOUFZLgfHO4OrR8tp1orUTwcPJJdN4szOPQwPe
PqVn6wcNAtZxL9bHtJvqqUYprbAIdRJUAYflXqY65HY3nHOOpAjybRkY8D6hNzuh
nbbgLhgCnQDSNvmzEUtFXo3xQ2MXISorIo0mp8QDbJDHcOGFB2I5utdd9YZTcCDk
zsciuZjFv4pFknMKiZryoE+L9t2z7aVCxDNm+5xjuTvILRPnkndGj2mOZ91VMK7u
wtMWHkUO9WCbBitSSUI2aNaahqsdH/dFIxuxak5hMcWmAL9XCnt7jRWChbuKPHbv
UDFmqa7Zvv+t9mvPWuwrGdx/BS8+ZuygsMHEk8uwcIIiTEY7bH6ZB+OpB8pdn4U0
uOSVqFx4noXaLgBar3scvUkJVZZlYwVBfX2MoFWBkUODlsSkmw0wZ0/C8EygIZEO
Y20gfZ7j7yNvJT3MiS/VSNwoAUviORSNzQc6mhBGrzZLeWjqFXwYzWmy34oS11dH
LzdgZ7f4KdeUxkr7hFKKkR/o1zP/J9q5eok72H4h5WngP7Nc32jyrJeoqd7bKHNv
8gFswKo6pV5IBv1h0MeSDmfHpjx16XWCPHd5CkMfcXGWkaQTmZeJlI+v7/xL6V5Z
s5d5vfO2IoVVU4IJVIoJH1Z8k/aQYth05vnHhMya4YT7eLYMh0umjMKsBRQj8SVZ
4wCNXLvZM/MY2GEp/q9w2N6OrgvW/P8pREVbPgo07JnbRoFD1y6VWUM8FfMKa8vc
QCDPMwkjbErrKD2278P/gSf+fEWvsal9kOJvlYaEjUtxmvJ4q4Njra4hTGko6ThW
SUKn+vxj7FtJ6BFNi79Vg0o1jmfOyQet78PFmpuSpYxDdlBDMPpTIex3rM0YAN5E
2cXUZbMpeOsrYqahmO4xbHa7vO7PoClxZ86MSnrILn+oh10tIy9IUPl29o5HM0kD
wfMElfgNVgiOhLW40weQfoBEri8buI6EwNqDr4vueXYYWY4p61KilZqFZXixfAhe
7vasqms4Wbyt5bPMNELO6LTMYCKC1GMiQDjcqdYxcy3BNoPmoeIvPVdtSEpnUPZt
TFZEsTsHhOCpM+KE/RWrhe2Qgrc5RtO3Q7JpISr06V481TC4+sMhtTyxEuW7En3i
9Z/ubEgwyldnOdG51iPWwi6vcZws9ql1o7w5pg1gAKralmF5aVmp89ROBeJKnO7t
psNGWhIXVSUglEiXBYGMfNf8YXBQIjajYVM0ntHJmzJ7tPFI9ycS5rC3MhIlj+dw
S2jePxfxYkA9Qp6AYQHGN7qKRmJvNlq5ocwlAPT8LKZIzRyNN/8YdRbKz4y80NT7
V1FRZT+keegOMk3cr3yDLI7q0sNP2hdUrmRR1MEsmNccpqcyXXWKxgKT6+vkbUY7
dBNl0tAZGZfKQhskT86k+694HpG8Ia+CFbPqpQ4NdxcwhLrrSWBZ+hpZr9zIpchU
dqEPMCJi5YPpk4RSuoX16LEMmo+4ZyrFEtSpcjWSqMpJvcPf5UId8dnlFHmZXmy5
apgEDPAcEEvyMQzBqWFHLJn6rAqOc+EPAjN2pbkf2QlODUjWT4uOpMcEvCx4Y9Kb
ykccRCdfVKF+e85rQ+aZb8PzDPpE6fO+YuaioMaPFJzjj0ajAwsL38K1urOSeLLy
ZpcxLIEAaGXwnIYNPRtlA+OiUS4iNjiEZMjplizFK+IFA/d0DjYANhSaNFA4lexf
i68499YdIl6cC6f+KUOWMMiv/8QBm6/lChNvMEGIQlTfTCwztwAuCibiFvVJku4Y
AK9c3Mn4m4dAE+rsXdbrVuEdru0eMO5NF2MjsCV6elaIYiGH/s/rLBp/r52Tm8Wz
jy4/PfZWqrzA4mh58vvFbyyB/Z1zU+f6+I5aap+fy9cl+NbNwUmHg424ZliibrOf
/0pSSzNd+53HQbPMDJN3WQzXkyc4NbBZcNsvFcsjMEczzUUHIN7U/MBaw4bfh7cJ
mFiQFaHHtiGBmtSeoKz550TVQuYf3rhPabagjImGXSZm1yI81+HJbZ23mQrpaMcE
yO2gC2Oe/J0xx3Twpf1gy3807rXEA3WyKSRCCFdn7nqIbH4pUnSYwjwOU7xnajoW
3hX4Zvb1pJ+NoYg7IsrlNPlcW/0JhnnuAMxlYxc/1rHRZZk0Sz+9OObkg7QARZ1t
YzBMtoGvR3bFgQ+wRYIlYgBMpB47GbUZyi38wwSCE0zxaU2upSTcXEK2u+jgUz92
X87N9WYqFL0rgWfyBX8Uw7SuzHfIvo+MPHSNJq0Dlt+1dJfKGrT+0Jf4BWdXQylJ
3wCIYlvX+zeBTyf0qoGfPEASYjQ2wcFH5HnzXr2Wm3QnYTqtDcoWI8CZMYqGIG1N
kbJzwq++jwzWVbXPQr95FNEeBuXvdoMZCYq4EknUgGMlmS6K23DNK0gy9HiLEBcP
w2NhpT/qGn0tBiL12h3GTMP8G7UqOC7kmYeiYi+HXl4CtXkA3as+H1/JQShnXPnj
dfz29pn+tUoMtYaMPXAKEkag1ohu2TDCDoJ8maSd7zu6BNzRx0BqYIvvoHWf06BP
bGvpZvhpNwoCII93re6TUeNyA5PCg7YDz0/wqLEkfdknFNdbeupJMaevV5UQ8fr+
xpG0pqBosq7MPLRmswqIkHfPn0Ny6t689PLZ5EaiTTo0g4Q/bGpld70lm9HGKAyq
uhu8qSYigMeM8JU1GUf2B8TNcqiXiIq9vZk64R1mBg3x1fgbO2JYlDfsPxObPxbw
Nma2A7Kg7gds2jhua1y1jv3FBfb9b47K94InERZb5sCfQop80XceoAqCzpZtCifZ
t8WTl+Bv2gLE55nrZwhb4rTaqsTvlTFGsreYvDSdDiKDrPtPHTIcbO5zeBste8HI
oYJoom0Yh4fny1S03YEfbOTvdWB8qE22n73XJ2Vs8CDLWhKQ+0DNDGbZZkbwltnf
KTcwOLEBmcR6QbsEedOUnVEvAy2GVuGfyBMUsxD4fW8pJRlho5GAgyLax3mw/PXo
65+49kNG0wM6JJ03RMSijWa2+dcgEZiWC+EpWdDq6/Uk63AAn4DNbMEWyYZACWr4
CYCT+txERUZs1sik/0pCuxZgJ2oSlpWoBj7l0SHjzT71b4cYKIoIrw/pFS8aeiSn
/VTC99QnrnTAUxq+skxlvf5CsLjnd/6RGkZPfDYnPBg7V+DblC81zbePw305ax2M
iAusTPfcOEGTSwduDt54lfNnmMG7yEtYQoNZNE2bpq4+y/xxqiG8ta+oOx1ik1gc
PjI9cG9xN/Lsg/CYtEhYcNl7zjepkPW7lBS80Kovi4+Q/Ps39M1UdxRcz9DdgUwG
NV+ySBXt4ptEsvWQqBvHcNU4g3Hla31NGwCX1HAkqxwICh1msqjJjMuk0s9griaV
CkGKVrCJTVuAnBIh55SKgSZivnfMEiJE9ZbE/ZFWIqs2pwr5p4XAwHZDHBJDART3
CZskE4Zgz35vvJSmWKvX8gXLTigAbe5720ic4N4i986Mgg1hgrGcZickdFcuSAp6
bwB7cGpAwLz1ArD5i93xiVZKfZCSGhlCMZQOaTTMVdjLHwbW1d3wP6xVpyWcCpic
+52l3mKF8jd09oAhAuY4TKkGKbqWan5OAsRc7BcH74SJU3tDtbH5SJX67VESG9lj
CNRdW8+8mesCOoaDo27MAl4rU2FnLgwERysRdspyXOGXX+nhk1qZvHbmuPpRvm4E
CS4TTzDwYqzxf5JUw0hjvSDZLLmv8KgFYPjg1K6kUQITRBmwYyvy6NDLCGXmdDSx
lGtyhSGMMQL2plLnqgxlPkl0K1I1pHD4IdqL4+zGRWSE1VF9R9HnMnM2SEkaVZGY
PmPcUhc6Rtv3hL/FaC4SmAR3TkzsVTD7CwFi8Qp1AfAl+SHVUb3/h5hID+KmGrNx
8B1f7OlRPVL0vtHbuyOXtFacqXL+9oJRVt2qLV3LJ4AtCQBk8Sj9dOEN/OBZU9WX
LHkgRwpjI61KxkRnHOGGxqqZbDYukzHqLIBjFQJQByfI4t9wSMhgZmswCEYFtHQe
hu0YXwD+83uBkQIPY0aZY2IVtR7okGIO5+/Sc/OprGvxtqhCu4Zq+iWOrq23Ov7u
tuWC1eKXiWMWxZkEXD5cAGxkYWQHG4ZY7swTR2h5T6OGYLG9K5hT1omSE/+3yD9I
rlKW+v1MivBTilOndja8so9LZFUnWmiSmO2GkSc8adUlTd0zJOueyxWJY/DO9Bxb
Ccf92o7EF/Yo4ieUrC+aQ9MrxR0xbatMC9QRCi5QlYKNtkkXaxfnJSm1fVs4xqyn
19P3rDK11THQvXlxxQ07Fv7CxrJnTe401K7Z1WjsfRhy9NnEPyPtXTbkmELrW3sS
EXIuBcS+ttfJ9URM7osQNeGissN7eBTSFEjWH0gA2CPUPWasDQ2e5SlhuYN1VQOj
kyhOe9oQoDqqRdkDFEL0w81cQ95b4SBM+Wy3PgSBz0aAFOEP8t16pBTkumBEbsl9
B/EAYKF03/2dGoDY/u4iwEkjIQGW/l2p3fgNe7jnKtQZQfbzrSxaBEA7Xa2DSYyc
4FLoNt/0vjwblRnTMdvfiW0lVZxXSqlh1F9HlVeAnaMycChoQNpV39bWRotLkz22
2KSK74q0QQ2ZwbsbYlnj/EYx6TKK9BRHk8NRFpR2mG5RvS5M6nYKDi78Nr4gcpTm
SsAxFlvV/3LVgzQZq+0lVrwwA2roWmZF8tOgi8BL/7+PFCahHewXswIzqghIz02W
4voJ8c6LhlLKpVOVs++pJsAtH22VSuYauFtH7Pq44RdwYW3fgbabFSIarXbJsbQc
kjmNbmHzOiPtY7t7vkaM95A1cSAB4ulDXdynFFRBYg5I4Dibxb9cUnc4TG0s4w+8
3ZIdzeVvA4/LTPwkud/GZTg3Creg3m+ZSc9/or++ABkFvnSvJdsOePpcGbfKePNl
VaGTmnbVJ5BvyIj+HV+2bNZfQUxTO9Qa6IJYcgD3PaJ6eZZ5pzGQWL0yVWiOyb7q
eDsAwa7cxyA47WpQ3NxXRClblVnoFIqjNCYcT9F/gK9QI0kB8+XNe1K4lhcksGSa
03t5cvjuEO8m8e1EiCckCCH1ZuYdtuP8TgHJYPNB9FC2iWHA93pjzzy8n7fhuX3M
BAcsTwDLsfOyk1B0445uYVuJWFtrMo2/ppLZjjzmaNIf5UhMNPe1sYGnT2wFk8qJ
QeEK84t8VUqLRN6KdhcgiJ/ASTMbJzXVFQAaPiNqmls6YmLZdSO5JGm25qLS7/++
7wuZxy67olhCzcdCpuLLnTXturxF3w5rL+bup+zzXGWu4CJonOZOPlXNraG5o9Xv
jdkTefJPPEqSaHXQd1bp13AACEcumsuDSttIeVAyl4IHkh5NycMx5o0RAYherSc2
th7NrWZxgnYFYW/O354ZnhIhs4XQYnkcHdPuRr4xJSDraZuQtwuawL0my1oqCKV9
K5JYDJKpmqAKw0XbPw2Q4CPS997X5D2w/AIrakp4YKoyQtADUddqPv7+8CXK9EgF
l47lySCrJjRSsBZoLGzyN22iE4FQEYvhqfkfahMIIX/AzZmCjj+SU7K+Pf1cT72p
BrAKocrVSqFdyXItzfs1UlKGZrNmoqBvw45ZOpTxOH+yxrMleJCHWD6Zf0UvJYTC
ktftPUqelYWAZt3FfapPPsRENTC12SKkPU9irVdENNSOKaZRrZP+ssRZUBsnNicX
+8YWE4OLP9LS7Yn7LScGBTMzpycwezAQCg1e9bhH6EZzXcosXkHurrq7WLVKv+yj
XKGmiHaD4ZGJdgG+pBoDpKsbrp1TAZC+NGcyXPKyERp3NpUjaGGa6dWZuX+Fhm1P
22K0bnHfWhJN0B00r891MNEw1tsQGFiYLbDQ7uS3Qt0sOvMZGWIkCndLgoO9qIVt
qNESGW9Oe3675m8lqP7PecNIF07GjXRC4Nzv2xn6jHb+41Y+yBeYj5a5UUYULUJ0
WnCd1Z3VIX8G+FWh4LmGu45iZeOyT5IBq8f+oBGz/Yx1WxOFvfzkwclc4hzMp35n
l/vOwo2Euj11QcqAMiZRxYyr14C5IC/QpH42+0vqpryrQxAaFkZ8aUKMk+noR8vk
i8FitBcYTcruopzlUqUJnZVxNMBMVRHtI+hTUCptnIEgOesj6QlvMJfYuZbcVPkI
uBJSkDyUGYRwdc0J5N05PsOjIrIOs9m0AAAKN/hucbcERDyqaVVfKacI4oyURRA/
jva7gFU4lX+Ia8i1tPhBBpbXD9kySQNMJgOlLzDb/4sgS7q4t55vmo3ZP0fJ0H0k
W2Weu9ePWLtr7ZrIxRKxN52rACppa0XFRh3ztBlRVp//Kg7QlWpZ7nthXz+Sfdkj
WmrPh1ui+DlN8/MMB14/OmNf9c+A4qby+qyiRDubc3MxZhwAkpGnB3RB6t1ZyHy8
L67tMFCZWnfyszKlJzSUgoU9oQLJ/3GQZ8Tb4MFu9LMo1bnUjgCkfVoGYHkTqGvt
VJMsDljkkM/49EoKF4zYfGRVB1aSG3C727g90QihFvJNm7b9PgOwzJjrCjz6X2pc
6RjEh5sEM20vkbXlrhmS9aDQMR6hI1XH/ytyExko6CY3BEkGLbxsm0PA5PcYrsGw
ouRHqtTPqlIKWGRb9iLrvlJ5SNgeQwpi8k+b7NWIKvUV49E1vsNaHR/IoLSYuRKY
7RamaB9cuVFtG3qNBU7h/LC+HMim2KPiETwMQX0NKyEyjZLNzA88Ak9wszbCNORh
0RorKjRT1uxtA0bRHJpZn3WjkFawG2kTNG3d76OFmfcIihVeG3OSSqgDKIN4LhH4
Jv/T5tdNvD5xlRK42uur1HwDtH9wL/0cvpo0ZCdLWGEMgJhWUfTJXxXOmGkD9WLd
Zm63FHEfj+E8jitH1QbX/qCS0AdKOF/irl1OgNQz43Q5SAhMDmw4LG9xOqhhfcCW
OYr3GLCX2d3p3BpDffkFY81ig+jc6eTiCzp9oM4u2EUvE7RLrit5cm42mjlPlFP2
zE5Kt6X16PD57E3EcrexYBBZ2+nm4FiLrAcAQyl61OW1kyuHcz6bkoH79l5C/IgO
rpbJagAJKkp1whm9r4ddH4PYx2gabaKfUgbGebB+gtsZkPWJtw0oiDiT6364dkS2
0F9MJ+NU8PkLorZB4bXe2U9ZzTpA5IOKpmOOeT1WLTaLW+F3+bmwwGGpzUoxvdwF
mGZyo9tZyA8NA9zkBBs4lR3nbO/+GDXYgCqZrhyHWiv8vQXVXEEBBNQM8xsEr8pA
+v2uYJvD3xNgpZjG1lwcKIuDDEOOD1oOSrzXKDsmekO6blknKtl9XWg7HaCTKIHg
CKfd1y7BmxjKRKGJ+K7lFMaWX69ujQrChtvg0kRpC9a2ZploPDqKKZhzx1gtYpKZ
mDBvC1V+V6ciE9F2jI3w8ijL1/9luD6fJxs/bZhKw80WTok/kFscnuFdP+fw4Qbe
qBlOrErTvx/8w5s68CbLFy+I9UZyu0MnnJZ831P++I2KkKOPeEp7ENqNa9Ob2bgi
Z7vSPDF9/O2y+5Nc2p4aAJwMka0fVR+XIY3VIKPOgjHsjB9g0VF+zDe8STHDhMqI
1pj39RqNrCWLWWKMqo73Y0vYSxeCe4ob2ElzF9+u2QSWjLkA2AJiXqAqAsN3KXtO
lva7nBTJO9UY++nQLYnMpSFoH8mHJREFO00yNQLUvRuQYY0PyDsErgkLjuURv98C
ZbZgJwpdw4zVO5w8wppYyYhsFsNw1yspFMGhikGH9Aa0qZ7R03SPXRlTadebZDvR
JVJshVvVw6OaKXBfu+CqzCKkR2IBbbT/uoX9AfjSbyjWZGXyMvmr5i6ipJLPykIi
Mj6yEkYL1v4YlaZTGHxoiwWO/Zs9uXz+QRdGpZSrj9ZA0z/YdJwaVurNy/96+RoW
i31sbw1Mb3OGGnF9Yjdu4lMg/y/RzRG/A7vMcw7+rufWKk3Ez3meHobAOF8kgeGl
lEy7BQ5WO5h5BJ6zsF2vrdZw8ztCItyIB0flronlps8widouNMyAlb6dFexU1Pc5
IrW92n7i7l/YAvfwJn/Pk4l/acSrYFyZwi/LeJXiG8U1lFSi0IEbpefNdSv8CIPF
T22sPguqht6qygJfDhzXZlZk5V5QRP59BOFyLafsQpJFY3x9PWaBCPOJWO9At/8B
WwO4hrwGCdOQ2ybHnHklj8V0UAeK/vcwXXsbYBScz5VFFieocUon9dAoY7KiCJdU
+LdNckmI4I2U0NR+SkJwjDIQzxlMABAoxBm7v0iRq2zFLLYCiZ3maNVV1TYhjBiD
Co3+D/rZv3kqqafqjBR2cl5Js9dIb0Fn7/MGFNOAflKBRViMmbIEhnWwhf+nHRsI
j18PPJSfxqnaNqbdBhrbi5u+zkVwpMIlUOYUfynUdhwzTNklDRsHzp2DHvAJIx8v
hvtT6iIaqe8+hP+murFkGE4UzVRqPDbExaQ+ONyaqIt55KOPRiOCq/GxcqayX8Wp
qJqifrfVc0qR5lONPDRM5xI1ggJ8zj0i8Ff/JAssBvKZzOk48GiZAL8J1VAOy9dN
yTGo1wXdIl/Hn7rWNXkc2eICbnL4jIWnedjYJ4qlF7glga0d3bnRx7wS4rhC6ayB
EYT0XtGsa5WUb3p357dbScTU/8D4ytjOz8OIh1SX+rcPY7ctGzN/q5Wy56HtGey5
qiSR0N3QEjBJJc9W7gsbJSgNcxGBao9u1Cs89ufHyFHPUIq8j2JgZe367rXFcCYX
bAJPp38XqCHtrfPcVUVW4gUjk2kZPXfeY5rJNvMVSW//qOqmTXZyax2QlwRbyeA/
SI1N+iwNfZIVfDtJr17HhhFlmnpfGJ2sfuIOS+tFOEq1rXDwMZgeYLbhTAQU62wH
NK3oni2doe6TvdBJ79kSyz3c5sB0abDkcZOZg5VgfLyVZV81cVpGzIP92H4LsAjJ
VRHkxCMnyrTC0z+kzal98aaQbkXRC9Mwd5gpOkx4oehYyHdZ/wdY+953YS9Ebtob
6/TEapqSLqWfMUM7T5Q3LeVKndBb73sc9gxrEb9XL9xop2niqGhRyzWY8a0mCvAb
TCnga9JpiaxkztWvYUhpJmiP0n//JY8ktdhdyx8TmQlKHxhE1TTG7euTH2XPGcCA
iiLsWy78NgK4Tj8yhsTJXG/JJimUgu5IVBCC9UFqGshuUWkJk3fyqxsUDK1DdRoZ
Jlye/wGVG6cszuIDDVcVteSEij6j8i4KGcIgNt8kcOeorqlCTqsOTviggg5nPvF6
QB87ulUH1zRGYrY6fC8m7L5j3QPo9oiio699+cZvv5xrH1zhcLz0429GlSoIRg37
ydecwTYArF6eHYdO+6CJEPJT5sK2xzBXJ2su4QTeo+cyMqmgWemVM5P4kwJ6RMHc
nJEOMWy09ZIY/uvDfPrl8pECKty/QdB7uU9F8ZrNEV7pkcH6dh8iSi6z1v3drFnb
Jpb3hXArAHkfQfHlTh8/FwBL0gC/ZdBtbUQbDbNNzYkMID4iowPX9e8kuQtXzu/7
Hg8KI55uGnvGKoYxEugW0e0p8Q62YWaCpRVxBwz0L3gFDQ2PsOJ/bY6oHaJP52hK
/t31dKtMn3y/kf3xLy/mLrVKFyY7O8Q7h37R+SOd1rZsRcUCRCod4QHNSzcmBTtR
IZgVPocHyunSU3MdqJZwEP8YPuVoK8b0wlyTldvUZATtqrSzxzuxThbiBlxmE4B4
Y10u4bOY7PpWczfl/cHvq3n9Nydu7yskR3byVm7S2A1Ti6IowjTTIt4RICK/t0um
SA0g8wIYS52ZbNEi3wLk62X//SjITgibLIJXvMftimwu7DxJSg+Fad2L3lKYioiG
PqfHzhNBMO4yymIEu6ObXKqe6uWjTS7TjFdRW1QJeDBjdTEi7gupfP2j/dfbRkrJ
OjCCtWdHSOvJIhqyHGC+O4JONemkQuGHWxglKysfvhW97kQ1aE20o+wb+9SojcYC
llKcI0M99WHnvD1GYZrAOqx7Q7T778FYSt/ar25gwYBLh1/p4WgsVaI0Q6DgPPIu
NmbYqPpG0KRRdQVj9yTq6QGAbjD52l9GKwMTXQbaWwA1stSy65KrraH+857jrtqZ
VF5ZauH+Z8L0qv3/dMKTihSgbR9ynxilTyvc9gzUZDakYXVMJqPDwJ68g7BRp4gR
y1Y+XsPIvt7nW9e9N/u6dbauA3gzhZGNXOW/78umM/SkZwq2CguseYyMy1V5/Vqn
Ezv5nCVDAvgy+sfQUMXfkGGB/hlK0HqhZ9QcL2CDKbq17QxiioGPo398VMPVi/3f
JwYNs6JiDDMDfJ+r9DKcfR9BpsMiHR9IK+6FlumehOtxTnf872eqhJSg2c+lvSe5
Ydlce221stcnAkkDBl9vNAl97v3V1CHyj2EvkAVf0KMnOOjEce5uldpX87l2jvpl
5RjgXZByrI0LJ7DHMitIYV6lTqRrI6qm2/xTn3MoQfxS8qOiYsHlx7YILh1hj+U3
Xbq79xL9lIbasBKJCAaTJRY6OA/VWkWEFN3jhdCOxeRlOWtG1VsYqX5msYZcZJwE
MGpO3ioPJKn/6JjRGDbPq3Lv6PNmEePTxxocDL3t6NEsdp7WX+QzVWJV5G82Y3E0
eIeu6TVQ5XVNQSt05EPcCOVCV4MCoKFGzcafVjx0ejycKcziftg1oeyB/7cJHsgD
3PpQVYKGmYPfVBfjeIWwFOK2ncb6BZqxo98H2b9v13bP0dLL0kee4USljvm1xGKU
Y8kxOEKnomuCE8HiJ/ve4DZvGo0IN5Jeifb9YZ2xGlDn4SPWJ1dgaky2mEMsz38j
XCsNpDf1Nr5VYWneWKmGM9ieiVwBEERtp8VsmEMGfwcHvOuLe/TUCbMxgOwdS6xj
j9ROqryT0KJwrbgSFoblj7+5XoBt653PW1i7hoYDaDXwlGTrVSyNrFdO7tTuBP2P
MB4kRIO+pjQFkzLgf3hRA9JGbeR85wHahPZKSca47P8ebUJVimu63C1USbRz9QQz
juJB2YBCYnCmbTLjdvt8+M46b506Ufv+aVF9q1rouQDteuHpw7w3wlYaoqnNvsvc
kNnILeOzFHAJykxPtzsliVaKYW3kVR//TjJoCqS40W3Fyux03N3izFzfFTFc/bEo
cw9Io0bwAjLc1tP+vBTNMP0KVeJkrdP/3I/2een/7K4K9GYXNQ/EAjZScUApPMwH
YME9l7Z+MXkumkTOZh4wHKTY/mXE8dK+o+ZVRnrvYM9YG2e7j+HQuw/NxpC/5sp9
KWFXX9JmqJTCINGkJuFhHtJrBFA9qTRnYND16MiYYkyd6qak3uUfmUJrjbcu1YPY
ghRlM5cylhzf0W81PGz8dUsVSRBezjquQZ44/szlGyeMZgP9wMEIi27Q2eMraI4u
BZM1TCS166Iq4fPHfHRVMS+PjAp/04xAJe3X2iYPt3kcUWM7J2F1x4vKBU+yydOj
0iPnYUfBrC+OLrhVoLlZVBhu3/Qa/FPbJ18YAoTWQeXYplOs1wwU1muH8NV/OIVh
huJVYsszlTt2Y9tllDUOJbqbPhTaOJMoCc3z7UpioJjc4DfDUQ8pGR4i9rskaDhK
VJ+pGvcuZdhWygxkLrGxac4zAaA0y85pYG7m+9toaeoG0viTfASLHLEI/ySbMUQn
ZqCSC4AZPSBtNSx/sXHL2DCVE2Np60KQfu4Kx29nJGODWeqJJfiehik1NylsX4NQ
iObk0E2UEL4eq9PWFnXyBR1uVtY6eBQA7tF90jwnm1lkK2sPI/7/hVWlhumUCPU6
3A13ndjg4AeHytBfYmei7qk4HOOeHTA8x47J+bV4yXydVQ8BuPIIYS1Lpbgi8F02
BoRiRZm1SgvnMScixAZfpi7osEKb1mnt92A+0awuN8hEldCLpNrxAM395+r5wAQ4
/YsBEkb94/AZcN5jVRl0SWYMxvlDdFugX9kLH+d8i6TQse7hlUp5mDwVon0lct6k
XQg98fhwmeRsADE/ZLFWDTPQxSTkzcnWrc7iILzxQdAfG3lbLgg6pEGifpFmmScI
3tu/KzULCssFMn+dwr/azIEKsq0l/4GG9E1bPQtiaZo6kt2SMZrbT+60wcp+2HmB
egudby2pfkadWq9t9nKTolLywSfJXrHx35Na9grwTaucqScwlgElY6kef42dD+Wa
wqLfleYp9GNgb0FnBOB208DxxlCsogki5dSebRsqmWMnNosc2ZEPLtoIapIEEHQf
3CRNGBqbDBN6cCbL8Z/VqpoSfqzTKgd6UNV4Tbj3P2xSHAd/YGM6CQw8V6Aw+VAB
3623JX22mUdR+WIB8uO3JpWc1sN9efV/MybPFdn4O/rysTkJ+sXY2sSGlyXXwIog
sKD7Zi+Bu7FdfKpugVkHFJcx40usKUnTzwMWEsf7FQ1bFLMZ2AoX0jaweDGiU6Mf
YikCIiojmzekN2kMYCL7eo7XOYecg6q2v+pJEy9QCYxcuRBjXrrQXcH0lk8Y0mJa
SzR2GEd7nomTSBsHjvwGSi+jtakpI2AWsx8Px6Zkt8k7eRC5gj0w1uu8F8NYi4hg
wsjcrIsbKo9XM4VO4rg6b7a+EnwjwYwxPJkbcLGouIkW18FBoz6KkNGBmGXD7aOC
8ngRmQAFTZ0zvvUuKHlgj51t3197VZNNMfxMSHoUMkzLvnxCw3Eg7xCVMyaB+ql6
yQwN4yDKaDNd+TeU5EctAFDXkJ71ti0c8tlo0SqCu2P+/TMla/BEt3IzZY9VEHS6
eMQw089lp51zR9IatiSOo9S3uJKjMtLY23vd4I3CXQWLPdalp6x41e7zqbh8HD9o
NOHgP7+rKqRor/K3p5sDC4KQbmye9SpsMPhzV2lQ6C7l2hW4ObNYXx1smEIdVQaS
Nm520Neddy5rt3wW1znI5SZkil9ZDvVBxPBfqZSnFUUvYSMCfZwdWX9gvDabegT4
MO3E7fQMHVJA66gLs/e3smO0tUZsII3CSOswbzGVpvILrdbHb1h6SWk9tNuSo51d
HVFFuC7Kn/XlsRUJnthKzhyjlv6i7X1cb8VJTf0N+XfeYDRFLaTMSQoAirJEl4MH
r/rZoJHfMXcMp+Ltkp6ZC3pCIxdpxcnQ1oGuGI+yQDNMp3qqwEiN4pGwAISMT65Q
fS2y8gbKyYqfhEv7e4NPrB/ttUaxxVL3cfo50hBp1GIWrUJR0P6mCwUHlU7T7/fh
wz7mvH3UWFtV+Th7NUAPt42AirwFifwRPjWvEAMlNbWaJHcW58iIGOK5omz97Cwv
/zq6x0QOyVyhawGu8SW6dBWBLYZYHUJ+1554qSogjbW7P2jFa5ZVUx+o6mE5laE3
3e70s3D1jFCSOjGS572+uAvZsvFlL6+/crAnWirlHANyUaRVKj440YYiSylPM2F6
+GwksqU2odKAqNNuvuEFlbLegLl9pMutZXFUAXxC6+MrFwFUeYKeF7gsRWAsrNLn
SvSDK8intSZ6isyL7+ivN/MDKJWqOz70KrIdnaqVgsGXkH2DkrZEZ9KvzM/nqeQA
O5Fc7/D/2joBvIPchLAxBjsgOUQGpi1rojWDDu76/4gqKNrIRhsY+bDKC7UeoXlg
oVdOoac7VfKatS/w2rVT1/gJK9Mvwz3ysP5xuhE0bRIPUQya2X7YWyllW2/39xaw
2OJgx0rbpZVltbxqfbsa+2MIHN3p9vO8QZVWcghyd/CsNXzQAhT/rmWJNzMZWn14
maV/hv7rCjQepF6HfTxsKmXZJgr2+iaz+YFMDd5o6z4BLr8pNF6g9B5SqwNpBfAP
LNljDKEz11RwgL4DLzGVR3oxJHMXq8ozzOvla0oKHR9aQYe1FysJroeyaBzxHe8z
yIGYiwS8TSgEFW4IGGKB0rXYJcqbi8NZlKZs2uWLmxlUJ6ljFp1Di3loRFOiDegw
g+TcZc8hpUvdIRt7mec61YdVL6QULqVU1WRbyy1KHA3nqrC4s9G2414dR6V45iqM
R0HNCu4tK97N1TWOePnYS+8YoCLhCtWCEjGuCTUYV26ponmthqClXIM345fvadTB
GF+B46XVlPWI7Bmqgq0uMa3DGwqrUf4jMGYagaxGR4Y719Vni7CwSnCwlKjnLdR7
Zw72yXFqXHRKjuoQ9tv2m72dycFRtDpmJ/CgOtMzdFWusF7eQ5h3MF6YTBh0KkdK
zlhpC5gaE9mzmK4yKd1QlDur+vttsoooTM1O2fneDmHLammdDYAJ5p6j88H4Iie1
1KRxR1DXDHiwRajrNjYPLA0L+tTyJdY2WdJAYUofqSLDUihuFb+gWn/7cK9e5YJE
+WCT0oi5uSpLTegMFSJ33KFVsOs9SMqpzk6B2ATc2ueHA+c61aJvY41ebEI4Ry9+
mE1dvGhDD36boeKOhdxsmV+TNKz6sz0d6fX/aNoRsKf6SJm8eurdSfRdMuSkTtyJ
EqxvSOpkjm/SJppLzJyzOP6R5kmsg18dHBup/JotasIeVyXAt15tIoqBB1iDNmqg
g3A5d7V/iUpXQDaNCTz2tTHnnVa0XkU9nBMECIhTwDmUc9Ld6v2m3iTAu/9h1OTX
FlXA0uw6LgZJjcb7zWZB2tc3jDtlqz8I3KRQrbfPrTsE2MRE+IdxQDltZoxkvmQs
DX90Msw9JogDXZtcbFw3ryo7PlS08rmuxbKORcQqjGo6YszsPUE1ngCI9ULebuWH
tikBnweVegte3J+y3zSTfC/vFpQ/B+rxMcEg4eFksjSttlESqZqdHno8OqGjFMpL
0sx+a5oyz3mVy8RC+4KEz7/y5EjZsba8B8bxAPYDdIjBkNe7uTtzdtLQLO1voANf
Uub+pilbkaxFU+zBBF6HDrOYP/iLI/ayV3VwU8/0gZxZv0+r0aZOd8mjU5fhzBXv
jyc0LmC+YdWPgDR9P6SFfvZsW5RJdVksSyOa7pdBZh8iek/FpaAWZ4Xik/0kn4+H
X2gF+qrb/cEomBnBzOR+FuJ6pEYo2Jidk7Nl3uPadgGyhiMmnqavp5sWMhCvDF/b
8XYolM/0FrAYonmSJcHbjKAl8I5ylHwz0MJCv1Vh6X18AIy/S6cPANhKdyAzrsUv
r+ce95XfQwwOOjeZ7T2MbOOSpyEKMwrcT+kPfDS+pV12SM3j/S6uq2Zf2A4Gdhct
f+hGUF0MckPH8LCpkoVpIxFHTmmLKMH2MhP0/A3IAOZ1ZEbQj7hahEjWfSpolNRs
gyHWfcFFaqUCb4FY7hs6IALGyyF1sivvWiNuilNBaqixPilbL0ccIlUyE4+71MP7
O19pMuZ8PKWoQmnZxFcVGKbhgGdwV7YuJvDlsbnYUWVn7oWVTwcbfSRTHkZdw2Sm
Nma0JVJ1fnFhC0Cjqmq1u7HtUbSzdrntuD1CiI/yePROOfk1te361Fat+TD6+L3j
aqwpkvbtG0OkXZvHrLQEytJd2qGpGzk62cP8a/k33tLu1heC4TlplPzsJaOkBnTO
zsMGp8Igcw2U8FN/kjiud8FyITzkxBKUIy//u8kZQfYX7vIuHuKGcEOY92+6aEB4
WUDyqQE70ShKXuwPwgiNbxVrrXtybG+vlSPIGKaf3HdC4R9Ch7gif/m7wyoxcDDZ
zNrWZoQYNfdb9mMG3gpfmErbLKOUBupo5V+javEg3WTdl9tm9bbHaORXDZqbcHaa
JTPj0xYt9/IoPtDtf6X5DjoGZICIyjgD+/pDMq4ZwhHSRfqULrpdBSHzMK/EARV8
OQ7KLtVfewvF7PluX7VyswItmyzm7eMu//33xddL5Kd8QClbOoEE01v8traII0MG
mbfp6PFvvgbtH2vc/i/2ZBj1H275Oa1viKhTW4MnUtl63GtcXHHZS6/aAUR2hoDI
RQQglyTHUV89uaSe1X+Uq4aghGokpwWYM9ReSnRgnC/OXXUZ4eOQ/VNX9Nmb+m5R
JmXbFyO08NS3ufJEG2Fqvr28pylaxQmAdaGaLUVnBxd+G7/ClyNaeqaoFWaaDosj
Y1Y6zrOPntlDuFZx5sjLgd75jMkycul+edtHn9S9R0SR9CNoqf6yBi0WqbmuRDJx
cuf1szAEFNLqEXlURJf0Atm6AkcapzTKKwYcp24w3O1IlC/KJY2CXRaw58dtBe1g
rYmuaJVAT0qwjRLEQDiCfZ00hQ+i8mtiQOU9I6yBh42u/dCcB4/qPV4xc/7ThmM1
zY0VDWuX6Dte+aYqfP1K4Yvd2of1EBaSolbf/2NPrj14H25HaKMg6vVwT09Gq49e
RnBB0x/yEWv34cwJlOxWzYdh5osJ/oPnPX2VC/wYIjt+1U2nRMOBQ04d8va5ghCs
EvcHxQtv/yhj0OR+HcxI8vT7O8KvisR9xDJIG7HQMNpZpy6qDAkdktUltt8ZiSBP
RVJDfoK/CZxCefUQ9EDZAMcMe7y5jiBpSWosvIp5c6/YJwSk7G41puW4kvzAAIX1
4pdvIckzvq4DrCb4d2maz52H+25Gfop/QzJBcbPCIUoI/69DZldvnGx7cYP5g0N9
hbEDVbhPV+PeyUvDMWEDqsgG7k3C+ayG0UH6O90cTf0kInZbvjeHWA03rL8gbnDM
1CloAqpXasx3/8+l1lB6248r6hB5Ron4TKeYKBULM9K/7usvvcsfLBV39V/1E8vt
iy2GWvI4NqBHJp6GMWydJEZ9cMTm+bYfKKVzjKiblaW2ria0Px/hdNNhwxMzvU8y
vj+6Pi3f7+55TPAzT307HVnTpIrT0WbWoBAERGUBxOczXoBZPSv28vmks4ixc+jy
FBK059i1wmZMQX351DxRpPSLJBtJJGnl34EevjT0Jej+1q/JUjjKRWGVFFcERHqk
X4u/YppyROg+LBcgs6/tn02STKRiTk/Bhv6gzv4AuwC4bp7Bbg1EetKBYV0xwvc9
9vXP0cWUSJEl1nKNlDpP+bTQFg2hDi7tNQ2vh95I1Wg4Eiy8W39vxkVHtX8nY99B
XYdrqxtnU3AbsQg8INc0hWOOF/WA7K35wn5Qqe4SwwMYa+oAGDp7xKLFgid6/s2o
e6dASo+aemvuDESeWHPrx2RXGWz759LQl6SwXQxDtKshpiHy2oIqciaHPtBFfb1a
cCS6oXlWe+63aEKeB7qBiMmdj17JtpQGx9TiBBt4RJ/Hzgk8Q1Pyk/QJ5SgDbDvX
OBQoDivKhLQMjA5t6BXK2sf3MTarjwCsHAeMG1P4B3Bjxjyqikn5V4ygOV7wNjRH
cCDSSfC+0rLIaN6qnOD7TJGwEbqhJvFuYfx+wr3vh/WoHgxn+eTx/r/cRxQiD305
+VJHluw4E3aEKov7CtLLJbI9VvHVaorPt0duxZjEKXv02tSPZbNI1Ylaq7f+o1Dm
gWv2/9eiQul6ko66OvzDcE/VoLO8ubRYudC9SmCmhCZqc/wH2yKXsBrt53pmRi/0
tABHOKmlWFwXuVRVKhvzvE6mK7I3Lt9zVlBb76qxrF/YDn30xH6kxTQdP+EoXSSF
A47qSF+J2aQmtBYm9ejDppTA1sxTMHzrlGKcmbTBnBgHXpt2pJEpTEw0KTQjjWWa
YLEyPj4dOXIcDoOgyPXV1Go/PVoQkylXOqkqQ+MB+66ww5DhTlT97thW3Q8dFz89
26nbM2VhCqMrQIVb26GUJ6+8znPmqZC9EzCh/U7ZvY06mCxcWEeSKJxbZHHzD1rw
JBlnopHujsvQdFdL5z3N6gdjeZENE+AjrPeO8+EYlS37xFSLeCLer26EfX3J78+V
jFKJSGhIrmSAtWBE3vAHrKHYk/viHJ32PbecAs3XCQFtlsAsThT5edFvfnwKveB7
kIny5yU5iAbPYs2/XKSECUn0pC9YogPEsbAUCgH+AsvGUEW1moUIWsahOb4geE75
irQE29HZQi1VVpBpNI2Rr2F9IHb8sHB6o4DOwvuuAo5e0hV42ewsUfbuAmX7phVM
MYG9p7WVhZ9005fhwnQR8D2B8TVtQxxxLF14/qNoxPvcpS3EcgNPpg2VbeMmkkAs
3J4tUuUBZXVXojFHhxszgyR2nSGa7cIZDd0h2ljDv8Jy7iXN64IyMM5peJUi2AbR
egMdJtejYBAxOqvwo3pmveXfS9HMGBhsSg40zwQbDl07/7wNFS8XLlz/2dm/Gjnp
4H2ehZR5u4/+5Q9bpHQOfZKx3fWhtCyyoWnxxgumEwcoyDB5O+dvNZd6bGqP0rxZ
omccUgCV0OizYFz7xtEZ8/Gvd7MiTIG1D69WQnrgfqNH67ENTAw2W6I30/TlJj74
iNKUFZleiFHlRrDmiu/j0OGrP74tdlD6Cv+h7stHeGccffbkFVwA8DUIcWCqaaNp
fz1m0wThoBxaQ5QO+3lOYPioCttWTFRv34zE37PB0b2DPT93WjmVHegT3dmrLyxK
IgZFAhR/onwf8LOEtHuGYK5iyVoe5zV+qVDCPLl4mAyE2pTfMg33CR5Y8vgo/jbm
qUo7Wl0sZ1C3lZZ3DgyeaMNDZu0A11ECwpVSeo3pGTEcijZPlqhxpOGL1TJEzpyW
Q6xLrakHv7LCfAQjwNhXVqnWSAdskOUupNz3kWyG6fGtcPwXzB3n4sX3nM2UBD/I
Xl3k/JshNsmVViWnLzjJdgoTJb71ksNCdx/i4ULz0v7ExAFUUj5h1pzf16sKXTDP
1yXkmJTjpRPHcCWgO98DbKdrriuV1Z2+9DpQOwitchyy1Ws4OBVnysXa7csw3eDd
TGqPSqbt26l1qLuPagoX4VGblpTDLYRUc9xbvkS2vfAX72MzixTJ7gLQNMcqxxO8
5qSj8LN3D7o3gK/1Bet4z5MGgje7Kj3s3wFpsxyEAV5QG4JTK2QY20r3Jr+yNi4r
hGyIErxSoXz9vJ4YpLzolXhwclSR0PYeuC7EmRGdEL5Bf1NANT1w/qgx2noYIK6X
TM9zaG41ShE6mNJ99jlbvFqlLv5KOxSVs4xc4N8MNcFxnbiaZqAdruSrYRgMQX1N
lTehI9PF0zgElomZ9n+AQHEFHsLkG88zKXoblggeq7ANeMSgUUJsgomyaCbcJSol
93Ag8uOA4EBJ5wzRzYjIxj32iHoKn+bpMQxiQ/JGZ2kM07jN5RfLNURyOahhqrm7
gfzc92F+3NOK1Yqa/aNwQsNRfKk4VoOxZq1/n5MGB7UWDqJzGybP1GxVE5Mx3vgg
o2qfcFQhtayB0vozVPcsFxzXm/+MNER3AHZ13FPd8YITA5hoYujlAlVFpsAZktO7
yqFaFHi0hdZfYJ+itoyb8nSZcqil1nwAdy+nOtCnT/LKnI4sSZJs9TCnRMY248Ck
Ni89r7FWWW0SMbMk9GXwiFr3qQewZFyAkSAg13g4+CVyDnDMBkOloLSjNcv/kylL
zlkFtUsyST5VvxttIWfBulhuV748Cd7BC9vXU/DREDMEEdYdBnNbQbLsPyBT7/+9
GdeD/YZXU9Jv98YVov3JrkBVOym5jS99ZRUUCEaPnYZbfP9GATiF0rQvb9bB5ANi
DkQohq6ACGBjSay5IPqhzL17OW7x7JgZukdYp6VG22Xo2di0eaMMnpYv+U3j1EK7
nRn0a3m9csWMU+uzGSCQp6+SMqw8Y+R4Wm0MCSX8+FFKwGjF0XRMPJ9hBWeheebs
OorALjthnbaPRabSeYaPuqOZMihaVRq3x8Pe9Ny8xfU0tBSr1HFtbN6LPKVkM/IT
RofFM5utE65xOYLKbB/dy0ryBbXpsGcKLxbBDYGQ5PXuL621oUizLcLO5dx77kPC
3Vrj7Tu+wWeyGeH+15RQn0WRtD/elullWpP3aF3kQeGXHMqGwlciZzQNnvAdwhUh
DmB39lRIXhoInxny8kQF9Mn4+f37mUh34V/spfS+FCQf8M/QkNmYcSWRnL6E/c+M
5F7h0yL+wYHqJgCO6i6YUBQ632UIBqc1iKUA13+df7BGQIriBIn06KEYipKZI8GW
PqlkHEK9kbXRGhT77C7HRsMSqNckm29PLyetv/jdBamDYKLFDzVArjjbp73/fDEn
e1ucjDTUZv+HN6+31YTNAkmWYRQVa1FKXzJMVd9zGH2hoIqJF4oPDt/jcCu9PVZx
dT2O8WsfNQc7XRALfGvA0UPyy50+kduuzWcevBYcqZ5VkaHQw66Y9jEqn4GDd9WB
LG8bgrBlAcqnzFfbX85dLeX2kbr4wPFrcKTpPFXrJ1UdETHADQmFC7dlk8IPT6XX
JvwVOWNvDO9rMOIKuVWnIyLysvlsw9vBScQs3EQnWLcsU+26I/u15kX+ecCLNOqK
maToy7jV5B7p0hG6OOMCc6s5O1HEoLqurh0jLBvfjzUEc6+RG55d4GjlukR4tTRM
8gB17z66xmqtf0E/yqbb8dNq8OruRzy7VIgzHepcegWr0YvAsI1KX2tJNgKXzXtK
VRz3IbsnlZsD3FMraJJeTEl7k+LlYHZ93945zUIPgHZOR/uhQoOUvHKA6jHBqdV4
oGyMbkFh4fnrL31oc4W+L4c9M9D+Oh3/DgGdqb2kSfncWhkSwlww/XonoISnDK2R
QLFdACtIguxpriMvqtmzWATs2wxd5bgEt6wV/amOaIHVW555bREy+lRWkDVT9V9N
IF7jISw94PqbZTjkR11wFkUm03fdi84+HcpuhJ6cKSVyXy/8SyetixHkqkEo67bo
GMJpvntkR5WrSfovLuMXEsEvdFgBwf8835/ca/5k5LouRSGkxd5UQopAqcBYfxyX
MLOuycYpix4NS/fOWMxXNwUhspOpF6OB5z85rGDDkmg86MzqxTRH0HoZTqnaCgR/
cBAPRNzzvIVuI7cTxhPT8xYJZNVYAxzmXZ7izJn8Z9t/X8TGk6jTCcmBJwByv+Sr
weQw8A8l+deYMXWMLmrPCXddJzng/L+fLoMOQzH3H5ZVTuJZYNrZI08Lpgpedhpw
WVux7LWIf9ouoDHHkvpu3WozAFXHTOzk407OxEnKYCWlkUXckdpp2HDJnvtmC2sa
xtQC2SNMrqlS2WZX+ePod1N7sD22EA1XD9i0kPO8aJ4hDFFvF9bc6Ap4+vA8jm0f
G5oCA+mgxUHPjUWUbXm2jAlMEqBuM89RIY/4HBG2oeDDlOZmtNluzQIhx1clv+9E
zFZG6fcTIUAu4nC5zu+y6+1ShKZpzI6mlYH3ImWfbia0+kDjFWypm4hlhHcoAJw9
nsrFEVm/lH3uVB0DEGdi9k68gtk3E2spPJaqu7Hi2GRsZIr4+MkWl4v2iRFdV6mR
WnJ1ZzXvjp008sjr+M0au+sUCcQqRLgyKaViIShuCu8oNtbF6yEKv3n7unW1X5F4
GwHyE6fJWMNzvUHYc9mCg6Q5BWS1I48eCOfNIPsU5kfMo1DGb+5ge7m6Dh49Ti97
DO9LSTbV65becKuqoiHSj3UBJWoDk9B4Uvc6CJOpzTIcDxwvnMy+3+yVzdVXC8HQ
ovzAWLuDCIFJQwmK5i1VNnwNo97qeE79zPkukqXbaHOd4q32xiS4GJmsQWzSWpqq
byUv/YZbeJ5LgdSnmYvtV2DcBUzxS4ACbtoIhqNl0u3s+HaQFPfVPEiWw/P+0PRI
p6JWsT+R/7B8wvhGuv8+7GVUGoTsRD6ryrhKhb+huwj64Y7QgsVEWYYnhuGFbJgT
874+6KDY1GEnV5fj9lmxIbFt5Jqd3NwdjPUeRte4v808Tjhau5db4s+QV0y4cp2o
wd4fg5DgVaO/LMGhG0LeLsuVPQXDrCTzZhoSWFkOsuN4pCqdqowRH1b2ocA8DxZD
lb+tzWOxNlvc+xnQ4q5PaR77dn4k4nHIsFw73k25iGxYc7T+ThNMKREvWKOdLpv2
WZMIJnmwQvXfRz/QIWK101JAqN7KiRZWnjtnUxrLk/3Bi+V4Zd5NTw76j8MRpoJ7
eZPsed18lbzll2zkgldOSK1IqSCyq6wss1l8C5fKiAj2+fSodqOd3uAYwWlqZife
XYlScyWDG3znUGjgZujN0BLaiIbUlw4zrzFibGOOWhX+I16neewO1aWOo2cUIDNA
5I2bEswF9a2RZidgqwdNWNSzJA8ScdC6N0Gu69NDeKZY1g7jjLVfSlz5/HemqMtv
wjmQuMQWc/pL03ZyIWoe/tnd9uu2mNwhzaAjgqA6Td5yfJ4vLWlk5MUQiduc1ZlQ
m2++QM8+JKGMxkTIjeEM4BOuXoNYgT5aODiqohudUxUgTi7gB8pdKqTDvI+FXOHE
h6aauAeGl/HTqKj1RFQo1MNnWKYUNxR8niSKqFQYuiLW1DvrES7d2u3xOR7T4gkG
K3Cw3J8OcES6hIg6HkmKNpRsqJVq5m8FNvvZzue9ZTn+hy3/jJXfIcUmC5S88rxT
zhppgwOrhXwruzgh3gfE/9B2rIWBRry3ewnPBbazCYY84phHrqCLZsVGQZw3wEzh
/mtkUs+2Cg8I9d3scWuN53peJmQS2kx3woK6o5CMGvA7Dsxy4IaiS+vSAHPoQdc4
PleIVCZC18wAb0uoLlr4d8QHBkJHcw27NplcJcKOuavnKZFJwUimhzWN1gxXYypx
XXg65LtshC3kzJoTBi8xWOYTMAB3oXwNvkhrToCeJV2lyOFzPP0MULPR2UpM+jiq
RhmubgWHO8ES8QobFfSlmg+ccvxDmCUv04uy9JOL3/OoC5+4r1Cp9DZCL4QHqe6P
0W7Z7Z1HyQGkVWjFP9UDmT67VfRh+nivnKnOk2IPDef2OCA3+uiU/g6RYv1GKccj
TbnIz2ZJuALGtLNhStgHc4Z914suvS6GB9gBWX3Y4N2Z0HrTLXTqtGvDKuTI8t1K
zs2aoSX+IS2PFU/DFUckTIm6yJXUcDbxEZ8xlfUBB5CoNevnnGqpnRrl5gwhSLgz
RZEaPZJ8dwv3vKjopAGWMstrf9kheCF+3da8KaSKtI/eGfneTETXR3DPcpcYweIx
CMHzLSBjn1X26QQyR3AEVY143DIoRnFIEooTYQfWRVAhwMQMRab7GoPIB46dJb3B
zz7lRys3aCcQ94j6ZFnxOwZheZ0B9sxvbqIJnKfub1NJWaj/Xi2CLhKe9morEVLo
ougbF9WrWr1BE6p9qU9Z9ecaPeFpkZ8mmAxFbSou2FnP/B6qMUOgUcugqtaF/FtW
bcV+KL0vsEuxwc5Y4S2IV1DBs79jfLl2dfRTKHawRHdot+0I+XBOKT34Nmz1UKaZ
Eh24wxNNA6Eo5VtBednf1YX1NUNYVAmiWvSiJg5jjrLfb3IlrdVMoQs0k7ozS4ZP
TdQAexihFmN2xGUI1ep7yp3RGn8n0dufQWNFq1VEFo4zxbHO7wy0IbDZVMAfdsZ6
S+S75T+O6hhMyI4kvJy44rtoCGEg+SQKqPlcQgaH86XuqufbNk+eRC+TdNjSdrNk
9RiDHaovqNwRnkLQPUZWVB7P72EXo5yPnN7mLlK4m8Nrviob+Cc5PrxP2kX70xSZ
wIuYMIOjI4jyFg5baAAxr6NTrUlL3wEEoJOelwaBWGfdtZpg42gz8gm5gW04Pboo
p5Hj9G7D929GaDm5y0Qeydq835sjrZzN7J4o+hfuFLsIYgz7//w5IYJFGni1eoBy
GGDM32htk8WaH/4xYNFmV9cljYbvkhMZFeL05l+CBXzNKXKw8Ukc1YUzA40fsoi+
7/l1iU+JOhiuX216rof9qLqs6NZ5AmSp3t5BO2u0mpCrcliBXK+93XJ6ANf7349S
lAzwd0raB/FWiK9CWkB4Nm5yTBPoHlavXaSvJWliRE+uPLOzBZDDuB5nQWtyaxIu
EkkthAF6+PO2DuaevNZwAr5p+VOKRdkn2JxIWxURTYTbCFXK6ZhZRz8fmOiHoR3u
PWqUPzOGUD/ct/dTAZFR9BT6SsNQn8Oe1lIrhy7P2Up1XqYDkxBl37gA5eHetSlg
9rWvTZE5aI/yroakGA5jOmkRHzMOzjn7YAYZb4Xv/FFKnMLJblPCCwJdRcOqDQ+J
nyz+0fcnkVwh0Avvb7mlAt7C+sZ2WyhAWBbyqCMZjr5ksvoCXulqlpxFaKmOXPPo
ONkid5AqohrjU31CGCRUnYqUrMAgcuBnmB3qs0ERjHTa0vhg/K7efpyhBgV1Z/8B
0AOJHLL7ux8FQE8E4KciJmPYebc5cW0G24v9MUJz2nK2rsHx4UOwYYWjZzF5TZdD
Qk+aiv2PBb6Lgrt9XArRxXFk47NUUTrVHWqx3y2c3wc9/a+7KFjXVTA6kySj7MeX
HlGg2AnW025iYYoh8VwmrHZWT/7m1culThiV+y8qu5R3I7fMjGFP0/5Bh/5ZXI/u
vDELNz8TrhDYss+iQFNWZKvkpHozpRJdImCifQe4xUvUUyagUhALp93jwQ3AxqQ4
37MMi+6Uq0iniZhSEw8DYxnqwTrTn3SDXAGe32Q0pFF4dcSBw0nEZnqEkYKNlwiQ
a9JbKjvyrGzbpPSoJHQzFsApDzG89DTqSDK0IRhRFcfec9NSvGKt/q4MTStchDp1
Kji61k9vJpQv84FjMjFu3BtwTEhj0cixApnRHF0qNVnvE6kGjHXOlM4wN6sFJ4/t
RNZN0sCj2viUJVFxnvv+EM19GxUeNgidWiR7XIDVecfMwxbBmfRc25lyj/aKMBo1
mMoPKaivmBYVIUKcguU5YbuN/u0VIcreOuNtHX4zxMXOjFW26jXdBQ9+eggV8eMM
TMGJ6uokxfJVHqJ4apEx6gYMI1W+zd3mi0beoXMvvv6swXrDpDEbEpp6R2nym3Bp
BxGJQkv6Uq4vl6a1nXHPuXNbGscHsf7tPODCyypW4pFaHGOQVPJVOsozy2GH4EMB
dazEm1guJNYB2HrZWca64UMxu0yxEL1ayF8+0c1w9/xMGj/nIJXvpJvxNzl1/nYm
lVmsF3fZcYUW3PgNTuAzmxv3pnuokDlKPfX8F891TJ/I555r+vCA9zQd19kN8ZnM
puyLJ6Vi6M9vtGvf0kNJGWQ1HCIgiWlLAwMg5ikT641xEnlwdsmDadiOHBewKy1A
nUETAc/JG0843ajOuV52F55iGTrQqqrAedltZtwYXHelFT5xuBczbs30LDU2Bd01
3TciZV0mEV1EzT+uga8LGu5Mi+qnEHSiwue89FQIFcq6PfAoR2KActMqifugHyLs
eoCRqiRzY+rt35rB2a632Efr51HExuLZE95j49bdPWh4avnv0Ys/gA//8dTnJQuU
/gEqqe/i1XmGyVPUwpOClDajbRuP3oBkmju62DWGq4ckWGAveAJAKQu3F/9BtZ9o
Pfi+Mm0ouFqgvxRJUL3sIgPw050Ya7P5LzClKmuI1lkTTE7c7krArwLX2G0jBLUm
jwno3glQdjvLDO+5ms4PUjzrEktc6ylpjUreUFhXlDhwbxCR696n5vKV9S8P4Uad
GRFaim0N2Ylbtq5i1czgAegiK6z9pDE0TjQJ9bPS2Q9ibSvI1SeiV2HPiwLVO2Yr
OASRBEhh2YQuuq2BnUi2hHj3kcabTHjjQ9vTNoxGMMGhkHat71ofJJE8FDfVAfri
tiN9vA9+K22wvoyP/hfU9cnRUBZKj/HvlnQzFLrL//ToAnMEvI5ciCjd2X0R7ET/
FTseUZl5z8MIeFAtX1oNux/Ji1rm8a/ewNPsiaom2QW/6gLXKcnQ9BJacB0UYkGT
+1vjgdUtzzaDBvoTztSQATMM5RMt+mJQjt9X0mq1E0aUko3xwq/o4K+XdYFN1OcV
fGWPx1jN1xfvnppmxJH/8CV22S+JICDK8AIKA7Ap2/ONutiGEpzrwl6gxsqkXp91
+P0mLPTJy9aB70fDKUdzF8PRUUoQbekxKwibWYgocFGGLHS7fMLW/5jLMP9BM/Rz
qhwaSQjaNp6q0o49zNNTzNhk9kzFbyOdoHv4wrjYxH6R7qu7V0ghCOPl6fBE7Wo0
mMRhBMRRoP7np0V+JMYWgU0CtShrx7xQ91P+/U8QfK+osBtl9o6wkLOSanPugq65
FQkCHM87aTMHqACa/jRO/FeTkuHQBZ+XKB64/U2lLgpkJPuJ5Ny2OC5+mVkyIDpm
hzkYXlqAP9a+IrnuzOdq23g3uUBu4ZnG4QhVcduq9APB1bKKR1U9RADUC6WfdCHY
rtjb0BckfvUNKRcdKIXEwzJlS5xeVzaJv9uostzHxMUqs7YiPzwGF43x/WMofmg8
eiBRL3bPefCu5bmVZgIXfZ4q/78kJBmNN3Tjt7RIbz3Hj8a9tErwr/ZQKpSWQ3wT
/JBmDGawolqoj2I6kpxBErX9TdEk10HMmzEdWKUylREz8XYhaioL7ml/5P5LKuTW
cEWIXX2IFkx8q1lc+JA3LgpMnzsxtL5cYmxkEbhRJCQofeqOwf53ykdL2L0lq8F/
Ah6hHAbzWsmR4YDMiOEh/58aHinQzh3i1XVfNv54vfFQZkKOBhceJgLhZ8QQAX2H
7Gm2UlwvyJsPCV15GhCFW0RTdI6Fb7KVWYFfosuxCFLfMv89WjUUYN22VzmRrtp3
kxp03FYojh34XpLtj1RXlJokFG19deS2mbTLQuMxDygqWFuuyijYDfGCHbysiaa0
ngumJVBzdObln+4H/YoOr9MY6y9/9Y6NFPA9e+XE3TV0fcsyMHmDgKpOIZ/tjJME
vwaJMGZNazreHVtJ+qCMnR8m1DEN6cT4WK54MjAOD7zj4V+WY7QlPonK4Fyf5d7W
Ysq6f/cwF9km4z0eF2wSwUWeqDaxPySsF2MSQWp+wUjbBHs1BjKpC94m5srYpIFm
Spi+IGYQsNfZbQZnT3xNlyFYguWZPdf5OzHQQU4IKbQjIerIiGcTKd9VLG71w7Gl
/G14Ov1l3ryh0ZO60mCDUfW+htX3wP9B3UrFiUygpGu98y2XrsMMfj7wcs3bU1CT
2dBC+WKPn0wtcoCgNhWm9TVlr4t65rMXLhFNeiRTK/7+1p9oWUXabjP6dq9pscaH
6crWVd8F22I5E3xcSCUDWr1BLIM5HrYH2qMgidjC3C2eLmVzA9JwD2rpG2BRCJTI
3LS2QZH11KibK8wWK88PmopVge9RvAcOGhIPmwf5da+Zfn0DBO9pMWlYGOvTuN+y
Oar0d0a5jixkoK0MlkT13oDNOfjLm5E9LglGraG54uRAOibOlBZ/X4CEomzKRfH0
e6CZLFkuzS16IPzn2uPzKlbuAxO5qaJQ3vtjyaM9ETJnNEDzdgXL/XEyAzHpuOtY
zXcZSIkSIk/yLiRcTSpS6wYO1ebPaB0EI0yAkBn9YbjLCov3ND88PlAnqPnGrHGm
65dS8XZ0dQHHH1QeJYPYbloIDUDUkF7ciAdN6Jg5jenmb87TvmKdfOWQG7rVf//a
mG38mAVvfUH4jfVT6kCKeyrXL1nmGoXGTFrhYApXaEzIEiBYWHCMpTqpC2tmbR/U
L9nrNUEk2bI1OE193HpzzqAMjdQg3N7lhuiYr7La8mzklUQ9J/8Gn+yk0P5Yv+du
QfXGmI8GNsBDDGpVRNLd6r9sVnfhUYk8XxuLAAWKaETqm+nDgX81f9XqGygdXHZW
qDylEUfVpKcM82kBSMbe5Exy8n8Ck8WXE97wNDujF1o5VEzyrGIpwnad8VXkWdlB
uCwr1O8GA+HXtGhn0ZpZBnpsVY4xMSo4E3WyF5t7XzJ4hrIMsDsQKBfrC6xcZwaE
2GvuFK/38XAQIIPSVEeMVhAeawjuBMqlWEdR8CN2U6FmifwuUN7ZnYo3y2no3iAb
uuYp7ab1AM1Pni1NjtZhU6luf/ePUCOvfF7sDV+VvnRhPZ6X+wvh9C97FdrF/TSp
sZuAeoUQa2p2T9xcVr2NFUiUnvje1Qmvl59HUz9YU66+iBxgyFIXFWsP+GjjulMR
8YaeWiTjJD1GWZgmsmagNLCeeLZj+J6rx7mG44jliF0FVTXg8FI1FpO6aNr0eL/P
cJnFri619kkTvpkJm4WEGG3DWqNQogP0EXUDbXb+FkwXzCCFlq0/E2kfh4jiL6u6
h81LrC1xT/tcEPrN/DGc3vZZ0jjpRF6tCInmD92rI7+UH5oRFXPXtuREToahY+4g
oGz0rdMiLkt7TpkS0lMCK28bSkJ1jtuDtjgc/wWy9ZRU0JBs1Mti3f0AOmcO1gW5
l7zSuJBGsU2uu+YI0ttXXUfR+kn7JAJjSJ0TWgvadQjPpBJ44p8CuC/NNgYNIBck
EtP0vB9wc7ky9EeyL1MQ9t0v9WDmqdZoAFi+dd1EeT3tAF9Jo1pvr99SwCWi706z
bCOV6kn/0TivRo51bnPTPV0wv2Oz5fslyEtP4coM+hKK+TiAO46NG8DSX8UNbvLb
PmFTAZVnEgb6aYCuAMhTozeJw6ED+9s6UX4iBHJ0qlDsJ6e2Y+2Xt+BVxXLmEi2+
lCP5pCWassvyLUqIT3xaLfVxUXq7OmDsylQcRzDO7jTcXf2EeqjoRvn/u50QGzuG
f2CGPBqpxNMPTFzxfmm0sFoEV98aaWdObbJhqlyUWpR6Iejnz6uowQr6yNOp7xXr
hlbo4EySMdjPffu8Vv/Fp6qM+JMztVjTvjaAllhY0uWxhbiiQXCRxNhc1uLlMarE
dBFk5GYbNQ/8v+8y/LdvXMcThuRDVsb4K4rU+thAbL0+9LK9XPPVVKh5EkBWb94B
IAATBMHJ8EJlpLfCz9nBTiRBbbPUb0veLWmMsi7E9VWLlkC2zlbmwzU8sHosYJel
3btbAgWttKU/AEuRPxqyDh9VsMtuoT9NMs6IrOSWOv9dWRj2bR1o8eZTpkSDEcY0
5KBsuMWV6bM6rJwypfBx/9SsFS3p+PDmBqOjt3uMWcuop7L5w/34Ydfqtx/R5QMr
Nojv+MVezLGx3vqcqvHzz1AcxOii8QbfvFPHXAwXVhyU8ZACm3/6803SEK72G6kI
VdtHr645rY8t/QxLnVWNhQyBI83+huq0wNPvUzn9NmB/6MVa0djI12M7BG9QEoKR
hiypozXc8eySJZ8j7G07Y5+5ouvrHVlq7mbZP9Ls5qgvJ4KOPnQ4YE5Jxc9sSR8N
Bpd1hXidRQ5qINAmmE8yJ5nJGvuDf0AK+ekx1LsoIQW721ex93p4uRGZjXqZtoBj
u7//Fk6S2/LAElClVfgPEjZDwfITLMGh/VGfrDQe/OeAxGsVYbtbwPudyz4//Fyy
Xiorvtj1kaB2rOE/hPsFTt+pjbFHeyF3e0vBeFEJptvpA+QGLJn9dci1VODhUAZ8
oGZYr4p5BVVV3bNXPgCsU4fSoLj6EhxooJzwy/pFDEyHywfgiFMsa+GxUCUyrxYz
ZrehGbBE43a0RGG9C5IW+iHGFi0XUlpdFsKbsP5CDfZKlCI+5mg3WAzmu++O7V3+
c5YtbfYbrntiMH6NaPVKWlKCvhQETT4tyX9c25osD07AeismrfR7zS8pWGYsPk+A
6T7zi3OZfIFDdve1I6TDfLgJwMpNclJbQf4BBfKLHFMnB2iGDyhYDjtesxq8AU9U
kekd88uPp0KLy/5uV8jV1YJT4IySipOd2uCRME0IWRVTGmBW30x0sLKRKfUQ2KXJ
VeZLxOHl3uk5KKFbBTEcZJ5biO1JynmM1/l2NDO/eTMUbz7JWMKilR97yP7eNg9N
DmmOj4fJnDkVTusydppQ2GWfYtAxZs4q/d1UGqsWNmn9vPWYBUt1aNkHKH+qHjUo
nJeiR1gD3zgvpTg3xPsk5H+af7d0jif+9JrOmEY4seIZsSmk+OEuOOUGOgEp1SG7
hw/0GbQv/TQOAyOr9KInM54XqB1SnqjxkSDBYzxnU3FCARUO5/dM0EVwCzYl8Oo6
ZljIEpEIqiBr8DND4S8Paz972Cl61VlQlmiIki87+/YnT/6NLv1CFPTfSxldYtrz
Dc1JaKfQDQvjoU+bTPeAQ28Qr626onIRXNCHfpq3Zn3SrfhbQq9NzX8HPJnLsAua
C5/tOciy2m96JnskjIl0NdmLKyq+KGovDj8k57XsLuRf4gGNlMxB+6WkBjFR+NmH
j/n/habXLB7IsgC663ZkrV2ZyFvIZesxRjZMopvxbyqmAnh0sEJOvGGmF59vFsgr
36pyV319vaqBb9SwFFfXvW4EjPsPZhNi/ap0Fbv3uiGMntqB3WfkbibH2VJtggPs
sp3gRoRawt2IGEWReIV2XYtrritgTvOdjyR5PbiVH/DMqAqXl5FgY27jhEiVo76b
m7wcI5LRJXv9cHaNRoyPSTd4J8wmaeW9YSnJmjvbN1b5AlZsnY5NYfKDXY+yfTWt
DY1ML/Dg16ou8aBcXaehjPqad1422WTlDsR8kONibEyf1ThwOaF/17FgSNxMUXEF
1ACgo4ASZrkiha/eeZ5TD0e1Q/wgGS2++Wc3+iWqaybXru69R/+pGDnZTuNEP1Ru
hJ7pMAhQI6K6Rb7b1SI7uXFYsjyrlbUNNKpeZ3lsY4S00dxaLPlutQGPZgVPXcNe
5e0mKElRanjmxd82D9VeL3vLKDnaYjTAK/pqkdlMCMWB+lnC025GQ6ucuSxYr9V+
aT45A7X9py235//AsRWZ/4pGwL8xsh/Im/O8HsfdjFdQrX9kfC+NvplZ3me2ByWk
hPrITokZREUupj40lXcyYa4yyzvI08adY3qbC/Pj8G57Lm9FwzTUakBrd03Q7rR4
k9evUSkrP7cJ5St3CyQVVCwddnYIqSkZaB1bPn2dDiZCXI8g65RKT8ZHIQyPrHwh
OsG7K76x1bnkLSZjMfStyRzpgfgyQCYzsN0W1NZ1HjLToVa8mllONDfPAJJhcZ1U
E+vs+oLT3D0Z935pPi+QK/XtCxmfkOPuENgDVxNdrxoHeVRM0ICDqkpLQM8R7ILL
1KXcda9gOnRn7khiWGwZ7wF0+Cd61At6IeRwxf34lxP1ikFsjSey1GlsBTmyJ3WE
TzjYhxw6Pwgm8aJc8YkFl9FEyE9v4JJ81OagiCHTxjVcIAEIngpEaHSwdpHlkVCQ
ttEqJ3FsujKAmIkVAh176rLcmgi0mU8M+Lk7ZlllEu2ldCQNXwa+MdsknqHggiRj
YLjTYok+H0TnTQEZgkYcZom+ftX5BdDv3Ult5opa2QraBpP1w0SG9A+Di3a3u//m
G2TR59PvETJ2n/nX6w+arwqnOtxv4oo7i6Gci9JLkrDI3Ejtx0xGDc1BReDgeB6Y
5Et7N8/Lgy/fOL1NBMKU519tVzgo/XW88/sHFye82ros9CMTgHVNJx2NTmDWVFgs
+cJQ3YcM1d6DRwNTDXwmsF9nQiiy+tmUSPm2xCvBJJt2jHMpdhePorqBBTqU/yPq
Ihek9WoQUkkz4XI4BESiyyvo8DmlVPvyYzAc/4MP1bdwUW90pqwaCCsPcKbGJjrD
JMNm9MzDpMdav//Qd29jGiRPfOlKvxFwrkbePwdydrrRv1GJKvDIxAjXolYmJYZJ
/z1tH6cmRMg6QqNh0xcR4xGJMq17+XJ6AzkhWmDzrb668ptzMneZHfJntCqX4Mz9
gFy2Y5J7DMIAW7u5p+R9Zih5gCCwwMP9HGmT6KSfBO4yNqEpRvTMSxqvGoAl7Pvt
6jLsAlziwMkeN3HhVahJ+KbRcuicXE/hqC1I7Uwl1dvwk7d1RttGz6nHi0cFlqts
tCa7Iitp4H3d7UQ6ag9SMxi5gp9ZJ/orKugVX4vPtIByKbnJqQoPM4seh7m4H40i
4id8GbFlsw4vO+dMKPEpj/QoonhU4X8/yw6XTf328mjUw76yFb/DXT6dMgk8JRIR
dNbYi1rIxGdSU1xQUG1U9Q2ODCnCEj9qa6omAMVIKUij9A7S24+9i1JA3Jfe30EQ
ueAgCkuAP8cYTl1Qof5a5ra6EN21+n3Qo9qpqDeNCclHO//iVdN/XO+okjgpJVn3
8lAGqUh05T0lWIIbYbC6718Yq2Tg4zMTxKaU8QMVAR83X55mf8PI3b3pGI67M8h9
lY4ZWlc9Yw7hRdeNXNEMfiDnAjDKDdShC47jbOVC3arvYYTFv4n+H9qIcqqlijUa
5EH/pQCQ9c+ZDMcRrAFxDekozmEoZUiV9lXnjNphu7mtI6kR1QrReQEfrsq23pvk
zU65eCAAqZQj/NB6kKhepb2Pg8KiD0Nwt18+orpP+bLJDE8CdZa8yGlp8LAiVZoF
+1mEwVn7w2rohzcijUnqiEbP075NvBbd53l71Qnf9nh7Hel8ED3TdaZb9L55yDiN
eIHXtOyzrXP2ds6ldAkNGPNbPzjhlZlOxdAxXdOzqK+mwR3WzQXqbx1y+Ji/87j1
olB3sjHNysK4/8haf8wvNnqxjH2UQsXWfQ/zn9D6/Qh1N8XPBEtz0k35AgJAyRZl
LUG7cC4nTF91A5psF2WXGcxBCPd3WYGNW2S+1e5mo2Y3mDbkyHMTv95ELwauqmjO
amH7xPHNLVS7zDbkMLK/APN7wVIF4f89ci6aLvTjTwQy7RPlFXXYGPl4DlrjB10y
7TbvaV9ITNNTuufqoaZ12ZZ0+iHmTHVkoKG3AAAd6s3FtBRuLnoEF1Nc21urZHgB
r06DLb5Ae2Z88WdaHZRuTN8932tFj6dOVG39H8C/CQmhTtCCAneIjxJ6mnU7aH1J
x/TdvoPNdrKIINwVj0kV3dpgU3FVjAe4/71VbwresFgp3ut9gLloZdcYiWP9dkYB
Q2XLnpMe7cWZVTbYsSVaTs5rCwGf1GVfX8Fpd3dS+hI8WJIkZshJnjGzd+/XJnXH
EfaMbpTVWVOSMYSpq466KHzi/VBZiccWPfpEJAQcrWXudFiHkB5QO/Rin+t86I8p
KYsdv28alMUsQgglqr1So4ck5ywMaKjITfu98zdWSQqDgXkB++ckx2xbqOXWJ5DO
HgrkQEIAn+v1vZ0PuucpLah6AfQqFgfF4pnthxF9S8hl/dMOCl5r5xCaTu5178uk
tndwI4W98EfuaHEFNNy8mHcOPhXkJECCy8YCq6aJ6AWw0SMK5xNJjH2/wDJa8Y+c
sylEayQ/LRgErUnxSexen11GQNDALIFV87mlvdYBE0No/uBudtFJTTSaqN/MiI64
9f1x9OxS68LQupPJp9esWGCLh0e/Cp6CDW/J7Z+6DDmrC7nTGs7eu+eHqM/iFMmH
DPmSgSqNiupKROHSysNuv4QeHWHS7VrAV0XHFKJUdEoqhJxWaMOvuU0Ky2XR//1d
5hE/fGMWiPkxW9imCWoLJ6Qi3eaYk3mQgGd1aeXE1aRImjh16VCZyT2pvM2el8kj
54V81yDHW0osxdvOKz6h+f5j3VByS12RbdpM4hLL4L3N9VCeIwfUPvWm/L/EK7hu
B+VbZu9bhz+0jF9sq9zU8hmdXvrXs/qFSPDF3msbjNIXcHDDTnWh71dGi7FaQWHg
pZFssn0oZJ7DQIoDY3d+BS3+xB6x2MG+/gBMtn1nryaLBOyIxklPuYlMrssVk0X4
G7rBuKHl8d4AOkiTWUYojFuMRqtVEjHMt8gXo7fmEW56bjpdVEmHsQh0AwdryUCg
Tkfb1CL8gjCIN42PFElpOy/+785VG4Ng7iSoddnTEIt00SUi74Yr8mzKLvuoVZy2
xjtVTEln+T41CfA5Ya8wggZ++iKWg0HdIwPXwb9eAsaE/A4/84fo0RHI+1MH3FJH
kg+1GLP6yN+KQ4tQtdYc8KNnKGPGV18MJQrlXZyHOwH2x84Y+vv8Fk6IIq2mVOLe
PVsGNHjDlVAARZaogIWxesBRqlbJpr1hXZ31CtDADMJLnSxme28YarXHWT2oYxKh
8wrq6V5va793h197iEnXwbBGx6qvA3S2phIgNcHvLNiTdr2NTK+h6RBHHEA6JCgR
z3bCH0LHZlioFqDHN8rNMQ5mrENVyzG316lAeVnp0+0JN3LTGRj0h7ts3I4dSHtV
WiWYddU4wEf44Fmn8BOch2DD7Uz4AkfqE9ga/yhNMAFHZevEhFwcF25e+JFiebIk
lrRNN4DHu5WeR/6BVNycU06+rXn0N7eTIhPlcF1wOmuJCqfZjheYIZJxCYyA5msI
vJPK8lPV+6FuQIvftH0Q3tMYiwqjwLWlny7ye/992d+ku8bM0GBeK3BNPLNskXui
7VYSWVDln6VeVsZEoi827PK4T6q5Y02vC1lYXowFcI3083NTxziMvvBwxv4wG5eZ
U/8wWdBrTSJgvF6ftJvOXU5nLJIGgGUqwROahyjSQCTM/OmNN0Y39DCF02yLWmOT
L0En3s0iLkxjXzv9+lp4Se3Gd6bzBIwpysjrMbvkZV9p8Kh7ukcuXufuDAK/tF3X
vJS6oM/9bwmjIIUBJwYth7b73zsnQ0eONyDdWrAHM6lI0iTmH1mDooz3RwGQi7+t
HxYhnkQEGi7mSXdE/ApivBNPucJwu36L5LfcV942GmQGB0ud8izvyC1CuYPjBJfo
7SjHJEdkJKcCgSmbaRoObjyvF7xiGYNmCSU5KldBYcSwaWCLZ3i5yt4ayZLmbnkN
CicpFLish/GytXtv8yVv1q8LeVYvxjk3nD/ckqTqUfUKJH4UqoslsEh1SCkkDwFn
cbsb2V5bXqcLfXjtZ3eZ1NNnOJXHoEUMyUUHNeJnQvNR7YjDBWETksMzNq9+HbV2
kePl/2+duyqJqJJTeoz9jy0YVjyDmXuMosqZ+mVvLUG+o0LtZonNwHBOPb2qK3Wn
2XDe1h5fZquTqNSAM++5571DOnhEXOUmpJFhqDr7ff3WCWwGTDE9rkmjBTV+5esR
K6vyXN71B/bsxEEZsyH7G9++2e9rBVlV8b93KC3O1haVVdJS4RdhbMvpjRwT1v0L
jB0XR6G3jvZO6tBKk1VOfXOfEtuqnBviUSuttRXLaDGoUAMfdK+kZc3lsb2M76kw
xTJhYbzsOaisJZ90H7IV7MqJeXfozxl+i7lxrxh7EdsjfH3P9d0sBQCkXvOVIcTO
LMeQUb+mfxDG94HslTB3yDK8SmsPS/Fj1HMD59LvkMWwehNGIoHzixcHCbeJI10b
+xf69Lo0OyL8YqMv+1fSL7m1SJ+pIdG+xwhcktMuUWgOVtVvNcjE9fwPqg0yNbap
5vT/a8Y5zqKU+3MsbtbVg4m78jKVtadVjhLV5rTmEXdxzSkgcFyhM7WVOh87j5wI
pMQ9pRttkD1m50eoWDwYwbTs0Sa7MgZoysjiucAxOXvEDPTppcGJu/HFx0tiZ9tJ
dUSUUN1sRpo7tG2zBYavrNXH2K1CQImud1t0TexIhTbG8de7QQCN1KEhaEroyrBy
rRIppmQCcV1p9VMvHmmFPjjDrWyBkFtqSmth7APHM7DXBavgTqNzacp9mwvm1hss
PApOVtTCgvDnqfdlb8ntlJvpBSJAe/g2DAp7jpkirnJD06B4zKCCJv0ZG0If0xjb
Z1vtunv0Z7Jxe2FoRFuAEW7gs2grUQrxTlo0VIRLwlIiy/qhpGtSFAtTUnNunIUs
B/wQfS8lA7I4hW9x8LJ0UabhqAXJ/xnUofZdvocfIvhYfKbcYDj6QFZlY5n4rQuZ
4MGXQXdrY+rxGKudPqgEImgGVEC36HxwYZrQwUrMKlytY5mS/U5yKl3FZuxN44vZ
RL2lUaU6UqGSjzrytY7BGxkVvuSRUUvHO64pGPmvuXgba2Zsk8H2+F2g3gxi8Wyd
kms5JxlvPWVkRCfTa+1N8aM8TMtXiQBPg/M7BmLRig/H8Aq0XB7dbPLvfJGpHZOh
LNrx+75mgX9jGZJgy0jzpYlQnNzkHW/FJzn++qbIvcdjew2OoNWGUUvFLk1CAeDv
ONHMxqgjn4UjJLsOyWRHf5+8MvWcuW9vKkSdQ69c+npXTla1B2rpmUgmu1HDcxRQ
akMah02JIJ7PYjMyP2VMqDNl2xEDelogLFRDVaVzio6sUKMUAdzigGaP8L39KMxT
3MdY8bq+Hnb8s6MSp+QanJIhS8CV1gfhVX38KhKUuRfWeRs/w2M6fUIEo/klUTu2
6CwGpQM5hXbPchLYWYqhHIiF/1ZoATkkl0XcotqCFEw0fLFKHvWj6vEhJin/w4zb
B/e74RaL2m+SwZeUs1SUnBUMD6q/muy5G2uOv/Afe9l//fKXfTBpOxdd9Hs1q7KK
IZnVSObUWead5ywysOIwuM7zeTz8qTWO0f8KjPOoWYrnyJz5ZKZHKTv/mSaGHmqs
uiYRhS8eFoFHyeRUcAqOO9/9asc/rqMDxb8l0INBHcYpRpN+B40kiIz4wA/a4ITz
AGBjcfJa00lW+9HNPoaOctYqdHB4HLuAr2Gri7AEadVezqUVmky9O5OLT3C6yaWY
l9OkvX8klciySN1Q3d/tYFGk0HUiS6QDvfvlGwDYzFMK016WNGQvTnsyloO91ata
K0QoLT5CxlFzN9F7grhZTlS3q7iBWuKI2g7J4Kybaqz34kgBmebJuD01hDSqD58Y
gof/YXkebeXl57/6GtJmQNIm8kTJqZkfQvhIrdqT4bD9UJFTDx4tVcJzgAmZaTAU
kOaPaMwL1DSj/XacZaDhIzWtPe4ZVqZfp1I4aT4h+vv38RgkIcJfpTUNWRY2ObKy
kwDt1a3egEDYfRWIxqh76BeQKDm86LY2/+l++1K2ok2M5ub8lLT1ju1ipKsoVLXL
OxB16P4WpXfYFSxB38uPkcPuS66jkbJP1WVOWD4iRoGenQE0IsgWswz34DAHtsQH
2Ju6w8avBqzy3ufdjJssBVCTFely/kEurpQetrmBLP6UFugQO9ay6mqqJ8700HI9
pEtrxbv7KOtu691T3fYAgt8AVKSMI+FsRBy+LzBPN5Rsa7zyAq2OxB30Z5xkhHDq
8dNTq/t5TtQz87dSJ9JIi9hUznSHDjhZd+VI/apxHyfnPmZslQ9ACGtYNgTLaNXG
ofbyqOWj1NW+Rlmo18O6Pk1XoWqU/66M4YJqyCdWz5LVzI43VPxy/d9XRgvkjm4K
qeATY2ej7MXxe8TvIdt6dxTFlm7+X38qkS2QksPUjVOxO8FeRb+LBlqpx1ck1akM
DtCmdYxTxrMaWVlSNAQOlduKrVPw5xthY9mRHkQT0VXyk/6U0NXXAhIRuK28mmN3
RHJPa5gyIsFSx6tOCXoYY850PtW4oydr044fS8ZTaVVdTttieGA76X+VPKSIBNeU
bfkZ511jTbqGGUAirFm0JuBF56wOHhmPECP55wZBwbMcXn0G3P70M7VMn0NxwrWq
TCo1QLG1pphMiVZ6sArYlGHdaGQihvn7hG2kOrXldp9ouxaqGaTVd4PcLt/DDUcl
HrBWFwsTuaQPh2CnTGp9JpBBO0WCL9r+iGtQ8uxp89+PnwNg6aTvQSGBQyklJIHz
hxOtvzhgViMjL/BGcPrceQie7Af2RLwrJNQzNooROnCI55/YYUXMPp62hFCeYgC3
Pa4YZvCUJATomaIgLmK9kcbUqcswMXxn2DvSxlADMdny2PIQyefLVQ4VoBR8azq7
uSapmMGvFafawdjUBR3PtkblpK5QyS1RaKJF877HsHcsl7u2a/VfDpeoCQLNh8Rq
7xEHQgnM7SZ4trVDxoE4rYmxZIta0qD5IxO1KCE84gBmuztmDRD0cXpAPXbiMrIA
fciQo+3EJ4W7e7r3/mVFle5nPbPPcMVHl9I+0InoPnZLYdU0L5yA10JklU+dUHU1
yySNZFls6YMFowNgitJaDypjrKl40o5tVOrz1tv4L1uv1nBvOCcgqU0CgqLPBNcz
uenFIJOgs6Pf5MuWfQZW2yUGlXh2DCZbzDhc6yBfvzBalh5ZM4HXSmzyA1S03jf0
aG4+7UwR0+sVJDnm9T82CKDP7WekJCur9zYqdFDSolQA11CYN5mvQtx8Gb0GzmH2
U6cdw0qTe0WbuLGW0T0/nUXtwPy0ZZR3TEds2UU9ASjpjaS7nYUyRL2ft5k3sJ2K
lZzpP2nfGG8NRYQHt5+4Rs84q/wVUzsT/3FGpukI1pMDHrU+dR9PiN9ZnhwolmRm
5ihC5tQ+ENah9b4rWZvEi7vY6U+7tvsduAXWYge8nZMyDOpupMI6supbnLMI7nZa
2AUkbPSk89E0jKnueIsoazmHw9LEBeVD9dUGraYP7lcyoZPwUtWUtuOkPqe+HHBa
EHs3ACtTiARczxbK6rMl1oq7IDE9sNzrpY9484ukJhD0butfZGDZibuB7Pwd2b0n
5iI0iwW286ib6IDItyoki5rs3+l3EkvdBYg8Ktsqkih90QkOpZ6kvEUK12Ku3Kvf
pPOTtnYsrrbtQz4qT7l1C8Om2yw0TqbRH7kmO4grB85hjIdT9LemkLL2K1lilAGs
MmHxaC5L3b03EUm9W1iZTN/V7/70w1A0RCgb8dEgeELnCZJUtNNkCyxBnqY8AwcL
+0OSlcMTZVGaT65xPSu22Dnm3fSJRSBJfLimuKaM+lmuSJ63PuJ+rk9BR2qnLzZ2
m0AwLGSYpykBFsE1Ua5nP/ISbHxv444+9qWuWM81DvVVJ1Ch70wMvfNE95SFLkHt
DQX51QQ0u+feN0fZSZmDdskI1B8WvMomPpbbGoVTH5RtcgoqsJjmrVqjfn1coYlQ
/gubddmRXuW5HgfWd/wE8/9X+CVB/gEf64DeRxhccgfSL41YOBXWftDcHoIh9U/S
D8lG3E2wh88W3JFP6r6giI/cX/4aO5I123JWjgObyzlZuFqtWV84xX+XFaKrPws8
8axwxYVEkrtq8UumTjDc5Y0DqUvPyI8waAE560dPfSwRMkxzsaDB7wvGeMUVSoY+
ey3aArIdw8J/cvAy5d9arXbx+qMDFvKS9TEwXb3FVSuyy7ZSICwIjTmXunz4Bkne
wa/Fv2MXYWzuxYRe5yFsQE8WeHMnYiu5IyoFzAN27cv7X5RvicUAm3sUQYemGtez
jPCVsz3en0v6RP6xkXSxqNGdkVnAl9rCQZMIdAhoA7TUR1hcnkypKwc6SUjylMJI
WLhMozt7ACgPkgxEg7A5RiqzrrSTibEjpbOmI+Ty9470OFToOhiXF6ajziIYsZHL
RuLuP5MUnKEBmVqQA3nFDNX2yRbeOQt3Mvdta8JoT6xEurgL3WnX48NMEmU9RM2V
ZGlsQvcDQ8ivnNjT7Iav6qF0ywl3Nq2dSjvhplDRMemfbAPxhme1B80CgV/tl9vl
tYTb2ZCyv6g7OWXLRhVqaWBQ6+2MZgzEqOK1MwQl1cxPzehQuDAEB8BdVToEq07x
K3EpPKXrbZ8C6giJclCMhHRLs5XTcFZkZ3tekUkg51i5j35nm6MAQQxEk9AfjanI
xdnjI/68nJFGGnxmKAB9KFSfnWxSh+c+dqi7fuyoHcvu9807d0gqOWMpOrRIlC9l
95Ch5zdBL6r8oMK0LpwNGWnNAWzBr/VWYKAuF3BbToSJlr8ZeoJT79W00rwCOMKC
3MZa3gcyazEuoesN0jIquXVq1GVQ0K1vDtu3cyeCdjoisQ5CNWQDrZW2WKGHk9uw
6V0LEtE5DWCdl6IWkiXsBKRjCKeyNOg3urST0gi7JVGUceEDp6kcJTV4whyZycJf
DXxTvKJ4TDNXbIDyJ0h26gKhPZIFWyTrfs5ymRU7DDyFVG6XjcQi18v4ihtihBFk
Yr+kmFO3glG9JTCqHFP5cDcqbUzQH5INWdVk8EQwmmH30ei/hmiKKoJnjkPH28w0
jdBlMdyMXLovbBpVsK/7zYM3N68N0Ra8y3q/hdNrQsgQg30+lKcK5ksphPlBYIIa
THwey4PsfOc9SENqh8X23qXvNvUbcdL53xhJB8liuhcZcxk3fSo1SkoYqjkNRlht
xYexHGgck5bwwXUlDOi08xhMAG8Qqwt2qEC2nT2PolqvOGkBBQ9gWCM2cwDH9AeN
Ov2g6OiRfyIs37XiEUPrW7vBnVuJX4SQty+7tN4E27M+Sd0vSDigwtgd2SILOyQv
hJYqQiwXu8OeGUDUiz9f0dYpnioiV4Qg5vcBegAFvIAeogyNs+2E8466Rz2+Cxpj
ofrmoqVAbt7/17qiCDiMUu3PBv7KasPNXLXfDD9jaNfgxnymVlN5im8H39t/OUqG
mpoir/qp3o13l6oPxeO0Zrnjpjub7BPWs2ASIJsPWbScpLYwuP+8MVSH/Cl/BWVw
MdNcuc+cPNszyJ86yn/BdTT97jyII0DezTTYp423CiTzieaEbkiOk5OKWICkXW+R
wVXSvZRUYFn5UHVLv0mGoSJsTvfhI6a1nvfe2609czNUie+oVWdKRoPlG1Q83niv
+WRtzqiIyum0AUTBYqA41WkP5kfcb1pRkw8fRLnwuznkZmxpHRwtaPymm8lJCkXh
MZPJMIZJtdjv7/50hmjod3GUgCfzQkiYH1zsuszir/lrI4B3WsoogbQxCV+9UeTc
EojwUO73T3losdOPfpZk2wsBWAVsV++Zl6ZeJNLG8PljomRRoC1t7bPVNGQ+HOgS
BzvvqT32B0eMpucmm6ksjOdJv3vauMfuZgENOdBtSCTV7SbhAHFzSA+K0teYzDH0
rThrRR6KFrMFJvqb8gnqN4WkDd8v3moWQVpEHYMMg5doCamhysDMs3dOF0PAB6bF
ny1SCPs/fnj3kzSqZlVQKpEPAC7SwUW0M+ajHtoDoXolPbfV/OCsKeaIcezOU2Kn
jkExpjAAdCtXhXG7yRo5kJwFVPTDvZxRYLwa7mS+g8yYFaPHfH3Dpht2h0Qm15sq
8WGNYR5qCzWubu+LjU5lcjEwBtMOHaKFcjt634cM4Oh56zZ1P6OgC8tfLKgIjIU6
7giU3IAKs+Cag5w4gaHnuHVl8hX2tUNgsM9m8M0drfDfUFBWzogEJ3t/lGSq6WY7
YbVgJhS84h8jc80VbbOX4mwnDCs31SXmP0/n7O5ph1clxdhf8Qh+W/dvC2a+RNoP
JTHJjAL+h1FcYesR1iBveN6su+VUmQ8lxQDXSsWv7ysNCoT7m2zyJU5QMPb1T6S3
pIyvIDj6hxjXNZ/d6ooBbl9wnhjrrxzRyP7nwOjNjn/noyb9DFuR5q57Lz3o4vJ8
fY36Ijg1bQMCwtFncAvIaMB47lKLHNbO8vLyyIDWGH9qtGrjkCap7BcQ7NfGEi2Z
7HZC4ullSbKf0iO8Ye4LRCUC72KhCRsWffr1IE4/eVhHJZzHwWzzZ4AlxfKz7jsT
38apJBzLoiz7Sy9gggI8liCUww3dPx4MoDWbiJqYNGdlv/uMhXDGTmgEk9IOYrOJ
tXLrpTda1UJ/GVZN5BBv5X2KjFbCIIetIYlOcgbLfkJ04tBZGaMXDPwk627prJu6
3VG5seF4tne7Nqxl0N9FbCgzHZ4HBPzTHMaYlIypqQo4RY+EkHsJ5FxcHeHAsidA
SPh7yE/gmASO3i6uzIKmTPlaECeL7OGvH7RpmVEXV/dhUhN8FDmk6sYbLI2a6B6A
BHbF626Y6fGDKvbRBxJ5CZQGYBdo4gzfWi3HGgyufNPlu+yoIBkxcQoOlyZ5mgNc
zoVIY77uoz5eKYStSdOnEI5uaj5irQQ3yXrwr3oiekAi5g/LhOjDApLc8h7g86RJ
+hEPsI4HCb2wIYHlxR2oBzytYhG5qchVFp6voyanjfvwpjZHSUZObbWl7jdlSpIv
5Bg8In9ofSlzrtiQ+286zkXMCboFK3H2lbR9wTUyYQUIHVROGvzr80nj0t6zTvjm
SQQQ8Uf5XKVsCv8ghrlIFNOAz2jXtz0hd+ci0uN1tDz1Pd8Cjr3Wibhdw9pUBFaR
7rfzOSAI7ldzWsGrghRxWJnCKaylTXA8pTGiS949rPq7tfe+1PzCxdt4szD62v6t
7BwS0y1ABqpolueuy+JOQtRfozLmhjq0X4nfus/k6DsmUspOhXkVTuN90XnLxW2k
jKjvVsNjNvUM6NNOy5cRfHgPZoVL+c2v3KBBDBoO1Yck896hKLzRWyDr9p6F0fhZ
gPOCUS/IMKrgrKJCYOloNSrzL/EeXMealJ7puPkV0VhXd0a1FgYhKDhmmoVkZAxJ
QjXpz6Pc1XqmO29RWYZqQIs/i3qiKt6X5iRjXIkfZTRKHG4vFDH9MehX6B521dkp
Iv5PRD7w5bGb2e8OJZhNME2/k4XwHwYEBNTCmVLp4iQeFDKebkG0FCbPzaXyHJer
GUKTnx1tk6QQ9Tc16jnofCowv8kePOlY7FSRIyVfdhKDkUiQN7K++KpyZ60ExCup
czn5B0tyQsjYSZW+CeccpDKQF1fq1MxX52iJv1Yg9g3ei84gj5JqwbRoT0eOFeDB
Tz/O8nv6pTk85oU9tu3T1eEo8Xf1pmFmxbSgV377J52bmK0AVLb2a2N9vNR6olBE
tpY1joLhhQuGe7x4lKCNDBjpz3tlKOb5Avwt32dxAKb9BNjTGIwmTCHfMGlfRBgt
uTFb4i89uD2crzSsmA/aZ9m7UDUnGakUfQdTgNaOp2HE8IASSFNN+60pc69sTsIA
em+fAp0TBxLKkRgUKn4/bAjd+P8JjAS+vzhJt3VjHNelXB3PEzj/cgDe9e1vOXwr
AEx1r/IbCT1f3xM3+ErsLHbr5ZC0MAVIUDIQP9/PiELzYYQoSv4YtihpSHRtxIS2
CHJYkEyNiQLuNdpgwHepAuANjUbWjBlaYEv1e2LMiG74vLbXIu8mwycHiPZalVLO
N1RsQ/MjtN+iGqAhDN7io066B7YDqmKKmNdK+Lf0e/yVP8OHeLoiGVEJro2lLxSG
gGaA434CJnrMzzHO4rj++7cMgLK4mahV+YxRmabmGqXweayS3ZY5KCXiCD0X2IMy
6W78hBp70JnUZNx50I9NTU+9Nlfg8ABaP3Rl8d5izZ2p3phmvXgt3wHcKAtjA16L
oH6teDjtkj6BvbW2XfFW8kh6Okkd7iRp5dROLTroI3Hugb0lZvlWy6iCo4f3Uobh
0bn5YfQ5lLKM7Zz3mnzOHfPaBf5JybEKZgPR1YkD4mQLfrVK2TXCnqxWvFOBKH5+
Kl1zrPUQBfcH8tNZR6grtZzGy2pvrdsJN5FC7+iktqTQqaqKMrPicsKMvKTy5Hph
aV2Sax9XoORqrMrkPRvGybkPsMPVvzdYieJOVtAteAkD0yk+kl7BbD8dVljQSWeH
4y481CFkgzeVEPDsdb8rkuxJyPqkuTC8UAON5bKewnGls9QNKRn+IC+Wsunkd8a6
OQOocwOXcIdq0FoSRpyryBosZG8xjcpTVgXn5HQ8RpSs2MKP1OfKZ42Zwsrz3NqU
0aRp1+t4EV6ohMXXX7DgAP9bfvUrijPvsmwb04RjL64sYSXSzCK7O19kb0Bl7lzH
g6n8AuCN0vs8hugVZhKa0EbL3FVcypgDIpIYz480QUue58kH1k8KmhUWaBUfM5bH
vbIcPKd0zs0/3Bm9BXxEXcj8lu7CpswOPONwfrz70GFFGTDRrXP702+t+013AQED
jhwnF4e1HFiJE01T2ImWhQtASSBkMnnCemS0v45mUC9jmY3khL3WNiBVnC2hqrqJ
A7mGtn4v/VSXBBivf5ssxPCg09NIerZ2gSlK0hPwk6fjyKCYBZqZYKtj24/SBU8e
CFIMbWvB9Mv3YkCKBlalVIxGoAHZ45dEZKOv879SoNULiXiZLyu9TpI6lQCG7S7O
o5Fg84kFmizD1jANyZFKM5RJ01ouYwIDpNQGGmTiUY1JBT13Ft2XYwU7r+jxPERL
guzq0Iv0FMR7hyfQMDKLPkMzSVuC8lffK6u8nqOEBGwwR21qFpcBpDkyevTNhM2d
osl9paRnz1VRcNWNqDvKuIYYveRUhY+YQbj4Jy2ejIaGou9a+Yc6o1DT8cLuVnAb
p9zPJvaBsyY6Rl0TUrWCqX1AQ+BOIUbOW6aNRvmAzjgksZqSExy2QoxUB4kJXTSV
hw/T22MpCLx3CQJl4rLoN45KHn997x47uZdSV5PyFtYkU8U61QQaQwQasa067bzM
F0qG1pL4Ot3+vkqJLId/PWMXv1vcaZGechRpdcIdGA6ssQyrvmy+Ekq+T6EgKBRT
9I0WXbsv8TEilK4n/vpCEI0rU3C5PUlZ7EIf2IOdr0LdiBKwLgvDmq+tw4TwcJ1v
aCFh7lKckwtHQ6yvxTjoC6FQB/8JG3bUAzsED1etJY28Niu0jsS2TW+4eTFq5E/7
3yauW4Ekw79X7JIEwiTcnRERx5CvoeMbQWJlq36mYNr12UO7hnIJshUXz5YpT7lX
hRUX3SwBMh0n+SmwT/1eYq2FARiKbBd0Lnvl4WSvJ2ibeXWzWZdI85phU4F0WMa6
anLopzzZcSdaYW+jbVb0TguWDx8563EFUwjSEIlK+0L3L3HNMMvS4Ee55jFPu5eS
mJUaR82BcsKzU+2N+cwIEUmQ4SIdSqfUZyUjiporJWLGwGYNvUhnzuunwgyabz/H
XECw5omC37VV5kyVEUm/j4dyoPSH0Lx0f0PXAEAWhHAUkvjXPtXbXtJTzZeZ8OOB
EMItX609S24Hi5L7Ji+AYGD82Y95z3ofQOJlWg7FfI/Wf6abuGLU+1FBaPMGhFG6
uvsESCjtbMOPzI+qmeqqEEUP8h76WKwSTOACQQqO7h7Y4vrg5+ZMbW8yO4rN+vFH
xF6R8szz2wBm5VeuOpxmxxieUPv1xEfxW4UmjTPb/XPUVl8GmgFG5dZooAVy/1gt
PUH1kQNeVIiELt2YBCK178HEbgoCl9JVEpXF5jIp6j1P8cyEOhMWrQbJ3QGg1bWO
7VIB3totcvCs8UpR8JbPjePvK7VPmfCmW0C7+EXy3FVOop0QD3dzvo9fEgRZI8QZ
OR/i8VOcm7ZVHfEO7tQk6JatCPdo9VjAYUy2wLszsPvzFAqzXHDgC1c/BxqTbSFi
GUSQERb3POgjHDr1YobbYlfWxy7yIYqrOnMTKDp+2XyqX51Dn6RxiP8lz/ut2Grh
TAh+hEiqs7pQ62w9DeTIgopP0/9b9tmXySIOBoaMWbbuUgm036aHRYZbXnqmI1DF
GV3RbWfdCtjBF6UY78ONtCXllcGiX/AGeEprpfldRyMPVEDzkNhlXVc/Mu3+acAx
xtbWItH1y9gSIPg+joMIEHSe6WGdJUAGfGcg7vS304kNGsUMYmgxp4ixjqJlKi99
nZExj1TpGue5KWJiP2hBjogzJ0fnRCizmN8YBdXpuffNmgE1bM2TcE6jf3bLWF+q
MO6+dpb8+yWY/DrCcYs4kq8DGFvsQA4eYGEyKSyqliBDKxf5zxeijzSW5Z8wWxp8
1NyMyyuVq9JLWIVjY69UB2lZEe9mCORo7wFOnvFvLMsHNyuIR7mXAxvpZAG1MsFd
dvTLwJ7KDkeuwujqbWcKO9ligakNJkFJeCqvMd/uY+yqgTIAWIgvkqvZvKI9GUwq
SwZIp4fagnpEZBqA6DwxL2MMG6ZJL99LtiF4621EwbOqcWwUyjVpTHC3wBM4cUon
d4dDPTgVhIKGCuD9U8E5R5Ed8h0byoxn/ncn6F7Qt3tlcMs4lzDg6KRs6xQNTga9
pIbG+2H+SDHQy93dTbWsrTWM6K8lCWTeEZNDsY6zbvCcREWHC8EhRJVwIYzvcUy6
NgIlX82nR4ZU4ACXs9pi0jZIyPUs2i0ICwB5eSjcvzM5iAnLs2AEpcLfKAiUX6cx
UOy8b0Y46T5GjvelfJ+L6+rn4FQqf/QmxWw0zXuMl/L29+F+kvRYGAw0QRuRSt25
3CVVCqnRU6nTop6XnyMH+dk/VVZejyP456I/4XLUCNSNdvcHa36szxd0dD51fa0K
wJZ6xroBaE71d1xQShpEUKQ9ECS/6/556pVZILUQ97DEubMjGf+UAvt1vnccN4Zt
BJtwlHv9T2HzhlOWnoh7k7a9Lxz3+xWZzveyq9+iX5tD1ZlgrTvK8AfnGGppyexy
H4SyaTalOjbAQ21Bd5PHuAKJhfBH2E9RqfVo2rJYfFlkTBp32CyZt42ENxx1Jp7y
8b39IN9ySsh6XSMO4uo8bvbwm73SHHarIE6xhYBBdlYcrr2JkqwEkBJPqUaTXNnb
wlGswicTIiEsEF5PTpxH9R9Ms0tZXgZ3tH+KRJ5/hAm0YM3YBra3XLt5v+YCoYph
MWkAzcBbNYkKS+Kkk/fG3RxHJ5+zH6iTZURHvJDUFyKxvTQ8Wpl6RnBjtHnj4EOr
ztSP9MAZb740zeWGXC2P0uniJFEcI+XXSxDs5AwJRvSTPjrLQGHCYDSD4Lwm59Lj
CHAabCoiUNUJNenuWM3kLMF3ODJqqoPiyiUMenrKL+VWRqW98uHlGcPi60aL4NGS
kxH9FYAKFmIiUv2E8A1t5LEcZb+kzXkv2GkjH2TzTP+QnXV9xsHVJ2VmPhgMBHu8
q2x6UcQFYDLpykyDTLcUHLwZgNh3VfVDylZWbFOmBegMrzTKxs3R+njGGq/JnYpu
33uK5LLTBl4iLUfeYCpoKM3Cca6gQbID2PT9M4HP9YT55BdQEelhlnKHSOydmNQy
F0ggf276iIXUketXuwoRZ4VPs49oxZgrnYXCjJ273Sd+vAa/N2h+EaBh10bj52P1
HxMmHEkhQq5hJ1OV8HWrA6TkZKQyx1MOaj241Bk1rcFQWXXog8XPofhVWzZH5hfY
XCU89M/2nWBEBoG5s84j2albBFkQZbAhg90fNB1PurmIX6toBzlwH1gfDdLvvKOi
RIIC+Cke3bP78PZVQMPjcMemPG4aENgPPBZkKsQMcu2kgQ0N65FsHVmjGKeTR8XU
/kdRgS/5im9sCv/oo1rA2vMm4Wh4Lu+mYzs2g85MF0HY0JRQy0RjcrFnZ4pF0Mu1
x+aegAoEYYFe57Ydmhf3prChwFkqX+M05n7ZMTwWHghPFySH/4ameLJuFm/jy0qd
eZJFC2W0QPEwVN0v4InhWu8o0iZFO8vEZ4HCDz4Az6m3ExfrBGZMqg/YH0tlEFcR
d/+P3928YtNXcshpLXuPZ+/l5fgSIJ9iSBJqG0DuWcmyC7lg1EIAHRkfBalp/I9t
tQ07FGYrSQNux1UsDA5dY508v5g3iMuLi/i2mgTPtY6u1VPXtbqvfjW9Xs9XxDai
M1o9s2RqnIaiOLsOyKbIWDz3So+OLnSGea1YwUaf6bI0n+sxGkUIj2fWMv+rkvjw
aGyEfxD1GHzPncXLc/zlceRFhqOSVG+xXtTWMTH9blem0g8NcPNcf/WtWjiDM+6u
HisY/wu0muzAjrbe/W9AahT44/BVG58uJSCwhuMldIfFOqI/tfWnWc6ASnES7gQT
Oi0Xrz0+19QYdQAt9IjMQab15o8QxpVweXseXXVO6pRh94iQNZ7BCAwnJZFI9vyM
d/mP4yFmy7qyYuEKq1h0UGld6mTtyRC/hVBylpoEw6bDn7LEgjbKJwPPUvS5T/IM
z7bpfe5Pgp/Co/1XDTL2YBKxB0hjvTpmz8E/qvC+eQC6190QTB1hTfv4UoKKiuFU
p48zOfrY9HpkAg2Wlc53jWoCM8xMwzPM+yy6EyvzYiN8I2CScBG4AmGQgcCMmvQu
qmQ79cPXRS0ayptQPzg5CysDituqP6mAHogSgjV2OI6nJpt8yjTZZ1tfgAex9sOp
6SjnyIzMy52UYHGZjFwPmhPMn+C4wfqRr8hcWt6lYX8CiSqOnvzImpEJ0E2bxJ6/
Q14aOb47YN8iYbzPNZqvc0sS1bxCUGyzWf+0lq9O7hXUb4MAcq92ES4sR+1upnmN
yaveAoexCKtPGjRsexYeHFvLbz+65zdgi3HkCKC9cE88WgXzGDJicMB4/cFS1LFK
RhcfBHO492oVqNe1WcARhcc/eXkmgdtaOQxW1/w9/UChSmeJMP+CWnOK5YgU3u5V
/dqsgzomxX2d62/zlO/s/admY4xgsi3amN4cUvsXOGYA4hbqFb9/m8lR3rLeftUu
qxOuzvlTp/HJBvTdSsvj1NeFbCOJDF7jqCFslQIL8gRizOW+UjKjLfOyDJfybO2E
xDPjiZOUaDs3qD2JJT3I7GmEHd+JsaOPGN5dgDFV4m2N1etqcL305RmwYrwycCFb
4leVq5sL5IBEjcTnw963X7HfbofMwsPQFBH5LDzWBSw36gSo4/9MZCYn6mqUAomH
PsNaPUpFU2SDTxsqPDVtoOkMeWQEwzr0qNj/VOiC122cKYEr7GhEcPZ/5zpPLt2J
uGuSKRSVOUb7k0MBmbI/Va7/bWFn18NgRzy8Dzeumsr6qjRag08StWpxch11O/9E
YV1fPyAmVHujjz83+QsvI6W+t02Nzy0N5c+B85TwtKQh9753I+GmLpBJz2KRgdM6
vT3vWsLm682XqtejdyraBRYlUNyBDzPbRr/Cve3Zz+O3isiE2G4oXzSUcypY8m7L
DoL27Yp8dmm0GXzf4C394agHF8oDwI5sZJ3+vw2N6CoMm4X3Ejlyc+1bTg7dxdu4
F/cT6dCQhVse12AkN7yOfy/lyIU4kBWwZWX8Jb3Kh0wwgUFQm8nBGGDDW3U2Cu8A
Y+FDr+8Ut3m3YfEZdEf9WAsTmnR0ETw3j1+cS6GCj6o+Up6GKx+FBa+5Mp5+oamW
whA2fr/8ue94Hk+xCYUk4rjv6nnMx5H+aeA0W2KJzpjizBchkcw1x7UPYU01jZiq
cEWldxJNB0iXvC0d75ns0NuQUcb/3KRisSbD/9Bw+bFqvtv3+erilzbowv3BSYAX
DB5yisBy3JeLo6N4jw8UsqdbWx/jeNzD0rnx5XkdjjihPLool4twutcPYtxjC8R+
K1e1g7oQBn7JYAsyK5CTfppWjwY3sIjcePc4Q4AGPzsBif62uFOgo7AEtJ1Qwj1p
2mAMRIWRK5oGBtYrMWTdnb/zRAt5d0q19oB0kAid+qMt7orQH5zywtkhTKcg9jEY
/9AzLzQQmAzkWzIuB0ntySVGAoL0evEnaAzZSHkCBw/8e0QOk53WumvyBTluo5Mj
AZ/NqwP6PP1GJ8dICaPrUabiDe/3TPjz2X/JMB9e5J8j4FEN01MON89xbfSRA7Jk
TO0+J9UXV+CMAiMykcCW4hkc9owhnbqVojgkRVF2l/R0ywqX7yCqxI4vgaUBcRS+
pNy7pZsC2rjowJ3M+mWjPSEVJX+FNGfZxplgY12ZgAcPAhrd7QNhNk/ZchsbpF4z
oK0fCXhC1rDFeQQYfa6qHYCwhUE4XhZ9laxMnN3DW5gyz6HZCeM4WlUuIAdnpvH1
R5INSmYfuxeDsoDeuLGDH1NJ1aruQ7K+VYb+MeW+HmxEKaxrAYFpfq1O1EwiHu/5
B0vNI1HLGp5a4vRIDoejio+VplIMoTxrFroDaFVYnmzMFmcrGKJVDCxSNS1whSLu
apnpYE3DnSbE/vW+VpDU/nxSkYzeLF31Ep/xtcU2Dm2M+CXodpzdn14WCRKKYs2c
GyODwPBGR9tszNFvgUnVHe8II4Td8umF4XTRTQC8COhmsi2NJzPuRteyKTNxNe2h
wAWLznO+AmQH48YlwcnEyRlY2kSGfBck/t7vn2uXXQiRxGRN/N5AiY8K8+mWeBH2
cxZdMq1UsjIN+aLr35laDphSj8SYN3WimPCq0pQBrl7byyqG7MueVNulsS8X0LyY
R0t4GpQ70v+aDv3nkjSy17fQ/KHBjws0vdx1p8eL1MTLPo++yAF1zzP8rf33wm+h
gfU3c+5+uitDrqi8e3gV2cgVK5r63w9duAcSQtc8bdsHzVzxFX8GR11W8nRS45rM
v/gf9CUrBPJ84+2vNMojwLMxquLZdKFj3Y0MJ3AKlA5B2bPgWoEvoBrtOgEjc6bd
RdgH+AwErg/28EJ/KLHkYNl55fkFI8qymCC7Y0e9bWOf7pMVitSpmJO7YnUMj71M
l9P2JWXWJekkiuL5b1SllJJxeu3PowGP1sY25XrmGU3Mjrm67XGDnQfOOUHUX6i2
Sfne0x3+/aZ72s5n64/fdwmBQfj1p/+DuBLqB69TZidMLxLiLJ9zp3A6NSTsYqml
lnC+1ouHmFneEFGEIIe2PoBtVujpowszj6i5ZQviBfpqw7Nq6pZLIQ9KJqj8+Hqj
7pknCsLBeWxQD1vgSl/b7ajDpWR/Ci5oqs9UC8EJQlazxG+esQAPzZrF/nHL5P8+
/wO94md6hmjFcJWVeiikOhz4ABuI8LQ2d9oECgk08HHKKHq7KR2wjas28OxSXZ1l
H0tw6GWFyYPIKYi6QPsDRdqXFMbJ8wqo0Wq5dS0GZSiyOAPxI/WpmOTgP+pqa64J
X9cANFZmOosT8i44HC4gBFD5v2vWU0XoUDwWr5ICTBl3XAr3dooCsLs3l6X2Dt3s
GiIPHA2wI+pwStgFg/ZwG9cOiSyA45nltUffeZL3sXir2Vny4EOO7KR2v7iW9LAv
uw26Nnx0z3RS+Yj0j2beTqfvjIBNv1Dn5tDX0iNoxioejPYO446qBBFnwToZ13OV
SVv+bLoq9gNjlzCFZQEv3ZsFHZ8BPyCWTIkyaAkoa0FTDPP5BBNIyTvan2wCMFeA
VcV2tx3QrjLc0IebIbXLauhhLxPy9H6IBRRQoqmJxavx4y/d0LmBdKD/5cIYycIC
9wpsTc8EwqWoJDAwy9c0JkoqDhNWTCmcdYbqNfKImuydKSoifVhKNs81l91iNAoH
Kyzd1b+CsvxN6FiWvrxVT4rWaR/Sl38HJ24Ju9qM8csXnNMdLTH7ysjDjVw3EFL0
Ms8D0JxiCkfNnUPx/Z3X16xtZhIAdRM2mB4OkWY3zodAC4JEQMHWG5WY7dkZ0nkB
kEKbT+1EOd+iUZaUX54o2Av+bCawdQdoL95Kx0FmaMWegpSpzX/MRBKGjsmXcbzV
G5RYIBah2fKt34tgxoaVLsuGCByS/VJNr7vQO4WvtC6FdB+QuQJ1EHZMKIbMCzY4
m/FiMB1mfGMg7yRwwKcipBrRr1PgSHMKv4G0gFccmMq0BU6WJ9UaKwRkKmYJPaO9
Qj8c9etyiqyX4DHRhRlZErjQ8dZ82ruLEGlbl4lNd3Gk6dC3IcsgUon+ua+zICHv
5/eHAEgVjjxwL0/H3iqYx6ALfZxEGLMYnkXkZGVVrrLCNUv1muO6yjV0By04YjOw
1h2UMwdw8Op5c18itd3L7bZXst2Xig/lEsEBFZyvh+IN51qRiWq3o6x8Nrrn4QMZ
Cb/bTnXpK9n60a37QlRp7xsUM1ulI1ykyuMIATPnwzMt+ap89wm4bD+oxXwfgFug
83iVoUYlh01HKzJoNXqY1yGYMmlJ9nUYYSy1/TjKlEhuWMz6id4+Bov0aYWQre97
ZpDhK7SzbM+cKITfeLS9t1iCbY42vas7ZvDPQWMCD/ydw9e31VDJDwsB+XjEsi8c
dG+lVraHKXtLEDqc4A5kmd4sTbTNeTW9isbG/pW73Vs2kewEPphY+pVOzrNDeTks
Sx4u3KR1B08IYzr5FDYbf1CvJMvYvn9U/wfMXN7+DMTlUyaZyEL99f/YDUueQ+U0
TtHTgb5tVzrwlyJSScUcxpvTJiK/Y3HnOMxoSTzjkgB8CUZGE3W3wyWzzeG6kKG/
J96jUYPeCriJRoayE+HCYuvB5zRltlAYt6znySLeiIpEMYLHN/iClGF5lGAeeWFO
PQDEZHvWEInrYLm1gQ7tCll21oi25JhW76O05T0qxSFCLc8+07hEnhZpt3MBHZ0y
DhXttRoiqtPo19wX/YIRXB5s9DnvwDp/rZu8lBFf4IwoPoCni5nicE0wRYmj3BoG
TFwR7lLC/xOsZ04mM48cQQCeBuvNE9h/Cs1RTqJPbWN4QqRANcWx7rnp2Zl760KJ
lRERT/W8fPAmo0YGcDHEPN145SLdIbf5TfJrIdlFex4IBns5Sn7GfByj3Roho7ZL
Nujq/WMVRfS/UgLCcUeY495T2Vr0bDIod6rcoqkMqAJ3Y+FgLNPKmUjrGbjxvqNq
KyOAnwSgsJ8XMaLM9tHv2ZZEBtjP/6AD9vmf3I6trgyyPil6Hvj//BxlAqAXYlIy
9Jwz2SiVdtko/499NISDbND2dslzv/QFjziJgdqEu35pOPX79hM7s1xkwPOmXkyz
F3c4tDCmHClcdh6rxrHY2cMW5Qyx6cfZyrn8aob1PeRvMYNQvJX4BM2ORDIxJwi1
nc/w7xTDhgI46u9E3G2kmtarrLT6fRa/zlm6mS/lLU69/bcH0zYbm7V6omJdKGWi
FjsnKAITDbl+25aISnht0RsKTmEa07YLrJM3h6hRMTqsihWTXGhV9BiIK0t927OM
b2yDsdUp1vAscxppF2xBEWBRqydYDm8nJEDxiP33g0yUMcwqoWn08ubJsHvG1W4Z
foBw05NacvFXvtHjVy8YCYUDp49hZ0sVpcCkrMr84KGend6n75uGK7T1eIJfnHmF
p4j+OB2F67Hwwy9DPpBfh0CiIKRXPnqLWlh8pOvmt6QtUSYNlis/hG2gmkbAUlEX
E2pFtEsVrebx8JT3k1+qZiWiEjUMpf5NZUWgRTnkfErsRHaHNlRYVeY04S2KCPG8
H2suvWPP9kdBybjNMQKnoYY7JYYI6z9ABOKoENg+KtOA1U1MaZrQT7adCstPpcuZ
3c27Vx7p7bsX+7RdG+Wj4VjOC04puw9vNP2syTi8p5UV2PFDUyxPesaO9Mr32kfo
qQgRj1BhDTVLAiOfr/rg5uKp2QMQwwycs+zthMn7b8sxrnK+vOCGEstT5BDBYqjc
owrp2xWT86q5EyEkyJ0O91d+MLB7TpKsCmlCOr2/3pXS1rkG8P2RENVwGp/kDWFk
oW2SQlEP2MPVS/OrG0xzSdrqhmUinvhqScSoRbSYqiytIy/sweM3iPXxzgIV6eRB
+kmO0QVpuI5c2JoViegO7UGF6rh6u8bbbV0+cLh+bNUMn6GoT+AKUs+H6lM9jUeF
NQpFLpzaHGFp77Zb84BG8Usgpzx8ypaubr+919/r0or7ucBvBhtfh7TfV/Afcymq
c0d3p0mtV2xjg33sibwrHHcmxzkeFDT5bAd+ndDL6pzRxhgrTOiDNLYOPRFBAXyY
0ChchCZPMKrtolSkmjeZHWY1tayQ/n2S77GSbtPUsuPHwMbcRifmT764h96wxlJA
qF00fjwjaMT9YHEzmkUblE9yiWz4Sna8kYVs0DrwKTE38pwOP9QCantJZlQd9/ma
QF9ivAIPAQsDeQqXSre3gfjeqUl4acSfZiWqdnyI6OIr30b4iwHg5EkqIdEsMg4V
exHGmeNPrkzkgUS+Gae9ClXcVc28RsCqJkuiK/pWxyWX5YbjPShAQSHdwElScuHY
zrq+wvMWLDApo9uDn4i1ja1pCfQP7iXHu7pL0PA1a0MkNDP3lVEPsw9SyGq/M/z0
q6wyFN8X9rtq6CcyLP+B2AWKUTvcxxisYUNmUCJExPJOY4m8aiqU1tyCfuNNMzov
2tCy00r0c9DB2akdrGZRdh8ffiu1ibo7XbAZyME+tM8AeNlcw+JjxascjYPJke31
AlZiXoDY5z/Ut2QfpY1Xa8iC18obtHVDhoOoP9HvNDxebAA9WWb/KqKa9zJywfOP
1B1dEz93jcHUK/ouzOEtcZ01l0dwYaFbXf3kTRwgf61NpJL6avJ/wn1W9BwtQrYF
UxIG+AWZ7MaB3Ron0hr5frgPz6jpQxT6Rz62BRALjqwfKMoksJaWMa44glRNQAfs
qF9XGt3/aN80CRj5eC7WYA1Kb0dzPJSEdmsbFUHbJ8FWzXCPsudZalnR2D7cdtcM
mXQFcyM2RvLSVNy//UHDUAuUTOuXt+HoFbRxJdcNxY/EFxTNP9+OqN7eFD2TL8X7
DAAaDMbuuEhmm3gJiXamK+oMM1J1nNK2FMUFPbnVsBxyw7/3ZBT1sFej0rApT+SW
4+ceXfAM/I8liUMIRCP1jw7oONJ17WO3mQfSYNeRMJCIoFV21MqTo+xvzRM6Ld/9
vtzWrWzuR6JzxwAGY8ZuoxhIln9pQ0HxiTzr0K/LB93oAD0DOriVK1k7sKV1fgwE
ta+7FXi3xHuBK6yDDZggQAokmXcpxDC0Tz3ZbNt4a5pciAfRxBFHRbitgp1Ahwz6
rY0EXBhVZbPQQ88f2ZSsZAlekNa3vjfjE8lwagUzPGxFqvSQsix0VxRh18Q015fg
A5SMIrat8nOK+645QhUQEHcJEhhLUmhfboH4qdCuCZHmWpR0pZKOtLatZVCtZI5C
lnvg6S8cdelvMcQgNB1ewyHPiPWVIlb7HgMcjteIPZn8vEnwvgy/RN8WR5g6pvQR
gAW1NsbO3QTqcBBSFBIpFxRKjbP62tNFP/DtiYGmmmK1uYET+8Dw/DT23osq7kWj
YRb1OUrYZcLQxJF7yPBkW5g6FPLn6Ci2iKZUMkMGNbVj1WQ3i9O0wjfI+aC0QmOi
gTZlArjorrGuuzDmSFopnrIo6xd/jvPdAdkfCtz6nzQ9KdZPUL+VbSwC0ajUX8HN
9witIPKTOu6e55o0zC4dTuA2rWlEtBVTwgWyZiDE22FdILLZ51hj6j7Wixgm0wYc
VKhPL93GbkZdKE8tJSsSGeVVvOqbkbNTwSsesSjYhNMfC76Vcp8xFcMceDpcRilf
HyOwDxdsbtdnSI9R3/WImSAJUq0ASDKnJqjzdSFW5OxbVbMwLTyQq1gmGn2V70+X
pds/dfQT32yds6By59UmwPBe61bs301fVS2k/5dWJKdh54GwqAFUXQxEBiRoqlY9
2zUx3IGBwc8OCeTFiocP4d25bj6X03u08ehJWoZzkSRVgHcCnbPZ2q36fbkvG6rA
GLmz0i64l7aBcvejb3wrPhBrCfpFvUMfTufHzFdY5ePfGf38+ALIq/1HXn9x/jlv
/V6bNUxYpVxNHeqOjv6XnmDxjBW6En1I2iUhZe/8GKpN6jFtkiLxhWHx0VtXRurm
3pgOHhY8gLqERLXwh/OowFzimVX5JiE0MoPVlGFHFvV/OZAHWboP6soKzf6spyuo
bPrAhSxDKHS02VRbz2fBmeiFKs1OT8A4KaaZlUqBhIVHvuXL7AvZc5Ggj09jW9+k
DOMow5qgkVhCWmVbqr/4+EeBlXhubErxIBX8hIbTdMsDEFzug0eiqiM/DWD/rgnM
wGLgH9Ea8OzSdB4vDbbGf1nBxdeLlLeS87SPG9snVP4EQgMrAxYIfGfcueG9G5cX
xsAOH6crY1YgTsmHYgc8tSEkX9EIvFksKzk+PAj/nAIDn8dQ71XUVZrN8aWm+z2r
CZ4+n0YAJ2NKwKCxquP7mEgUvg0fb0cpptBtnHjHGYUvc5AvZljaAf2MZgO5M0lS
XiQ6J7j+gzcWwy3OjkrEs2FgIO05enmri530q39sRNk57CyNhIWNiPvzUbQn9/NB
y/fxvrSIckgQ4aQMtTJEOMUMp+uJt+Y6B7w5l3Q9IZXjbFkPfEZ5karFs64cZTFY
J7Dg2T3aCeJWpjIqWWUoqeOj78HX03zpbF1ZvTVrL0S//+HWaDQ8sLGnc7AI3XQO
BtJLgT52vMOuFxcj/1r/62E2Lxup4W/Lu0QYPdj2EEM8uDbfR4aXGWPbd1yVcwlj
9u2F+RW9gMKvXYcepTX9nB8WaB7bNhgT2WLo/vcxb9l/wqND/LRL/JuHcD26bBTF
Ab8KdlZ+WPjRaMnQ60xZZdurZznsAbGs4aW6L7IlTi7AmtL1Pi6+iVoLRJ0ldgqB
m/YAr+tg3sf4OC/aHMfYHfV3bnzGHDYaXIlG14LmUb5YOim7F6ySdHGQwcX7/PcT
VSirRQLkdRuSGYYc3hJ96q2IpIRAaNAwkXg5liCuHaFib6/+hpl4ON+QO8MoT6MY
JedNhzxlsqjungHbeaWdS8giZgcxMhfsRQ6HIPxcywdaVEzSZhdR0Ut06yzEvHoX
1lMkWAq5ermH4/n0cOunKAhWR4ADqjh89aZxWeUcsZJn9uZgywAZf3+IpTO+8yNz
YXiFXCQivgSKFHoaEmnUvS65iCrdMaGf8/Agiz2qVk43yJ+Qx1D1FiBPU7ou/yRq
hw6aMMbpA4bi0FcHK+E9k7FAtj/FhuYueHuKslcmDj2R4WPajZbXYNXtl9ghVg89
8vo+BH83wKKdUxFv1fQQ7oVAVkACKFlnoveQT75iPxzOyFUTdc1heqyrS8lzpKjT
K2CtdtwyWIpJ96MooePM6fGafY78Y0kZVfk4bblXwKqqLHzCx9qy8G5k7dDIRk5x
KWp1ECsF7BeY5dKL/hmXMlPRcQEc49/R/iFV1/d9sIP6fXtW98eUcLK38SsNIS3j
26plFd/L+elZQj+A+P+fzs4yp6lUNbG21mX5SL/n1oeBtymqCQM3Hj55hR0fCHKO
grC3DJ15Od461ja+C0Wf8WCZTlIysEcHiAyn4xgRjBiLPTDLmvWHcdp+lfgHJlu3
g2Z5e5tX/n7pFxZTzuNcqeF/NN3VNBuodRYH3YSqphRdP/aLI9NSpy5i6XPM7j5g
uEXwm2DuWVWPrJXWyvkMabIwjodlr7o2wspjMh+9yUmTnQNTW8vkZoNrCncbX2xR
MpF45E9gHFf+zF8L49BXQHmjkzWnhEWgzedU7Xgos0zOrLfj3zHY4ZmRx90YvYF3
sbnfwHW248johP2e2k9TIKdKnCcdPWF2NIWFkkU2LjRc9K6PLiMhS70h9yFP2awc
z4CYTLquYR9IsP+oIw3lbxWqqhThptWsBuqFk8z1lL5l4AOFqF58oESGMiEoYhri
8ZNBhYvtXd74ePCEWa1VbUZVAzQ/Srj4BL27BLItcjqE+czD8Z3acxvJQ7SDiz+g
L+RT7vFOSqjM4iwP7dNe3cHUwJyO9mQAzzmkRA7w4FpWrT504HyiNtQJmdfROx+I
NpH9iO83HWA1Y0RDvonVohG8toNxl659kTLccS4mK1c3ggky0c3lkhDXYlSuNpx/
StaoLP8UJAzRh4XlzYmWHmK9GvH+RcAqd06/y8VBt/nAfHE4EVpyumFMemSpSxsG
h0e0fQEWbPbKei6venbEbqFfvWUh6lYFFp2YcPBo55cfcMRuR9k9SJeIUNOTpfBl
XQI7pgrTjLU1fFIYI1Oy1R/ma9kjj3DKMqcIPMg/WMSenbsizyywbBxFbXR5pExx
oslt2ntwgNFcXB/bZn/+15d3LphhN6KT8LaPepa8tG27cm5YHIO4c9NqtIFn5h4C
HimysHQAG6EGJN7ppL0p/qaGosAaGKl/Wwrb/fq7ly/H5O+eRj5aC4hL4z7BFepK
VkKPCBCb1qKkrsuHxC9LmyBqynCo7wMhQT9DYBPObR9roX0pwGOLVi/FapR93rO9
lZakrvLHqSvo3kIM20lAi9uhB2/hNAH/I1Ohi2NZjKiHCEkngCn/E8fR2mlbNb/x
I9PML9Opszz2HGbET1+IpuS4JHIznek64gGtswCF4HsCyPQexpuzjj8Bt38PUwGs
6NCg0zwnV0YiYdXGV3oJVG1YqRgd91KDrMm1ONIg/F/UxAzi9HUaTtSiPJP9ueRL
fJUfWac9d2WNH+ZdiLI03kJCh3YglhuBT1obwZK2e7TpJP1hLr6BvBNL9TX3luYb
50NKLb9NrzuAAAqPNd1hpa7dRQjKjcEwTq/3hpDYj77a3G6UMgbvt0VCot5RJdxf
FQbc0i+mPpCgDW66H8IONQ6AvIpx5qnBJqwcEsRZi6nIxSV4ebLnXcqAEixLc0dk
HnOLtbcHFK51fE5kyAdmOBRf9/sH+W9MABNWdQZ2fCZdgdRZGPEsK37riuGYS8Cq
wkwfhBp9/VkrZJ/5PgEYs9NUOXKE9r3aHz1ctg820nlKwpNqRZz32dqaFIzriEM3
zP3NyRk9fpJ12Vz1wjejtd85klQFMwQ3HAfUI4pjW0fm7MvAZxpEU0gYCO4RycXK
Zq87DL0h5etjyOn39l/78dMgf2mXzQPeZWnZAaNdlB/aov4/CKvOClIyWfE2ZyI4
yWqDUsEOIwLUoIFFQB0jgUhAHfBnu934QA3JuOaxFO/XYz7mNh3N58gNJvgskzwN
wwqfsiRu58HYa/jHx76FwBm7qQ+pbLs72pDUD5ktj7W3K7yeACc2ZoFVrnvpIw/m
FpUPMPzw1dTvxyktl+kk28jof6N7tSN/vfbldK80pADqamyr+BUb/xcxSL1INvHH
nO5EE046W1CikXDBt4XihIyo8PB1wCshjfaM9ID6fzOAqaDWzrfoeZZUSBkOYw/9
uMQiJz6lPzkBJReAFRZHXCPz2qdQm9d/14fMOjUQPJnTnq9FLx3lgBFuBWBAG0kI
TCcRud1gmr6oBHX2uP3EK1zzWF+bjQ/FLIapFWj6Dw4kT3ZtsF8Bm3RVLA9nyLJ3
DdU/Ytviq2FP74QAVAFxfxO3whclHT9TgHDrWxYFl+S0QtZmvhczOwNcSJuqVeBp
YL3PHza2h30h1eaUc2g1hOkxcS+ux/wvVX0LCdUIakIRjq+f3eqX7NgT2Lm16B3z
1p4b30uNa2dEXIdX+iFvXo7bHeF70QBtnnyscQoj85wR4U6qOwhSLpfaPCStr4R0
hlSfa9yxiNmYsiI14FtF15/49/Qu6t1nukajWRIkkSD+3EYoIoHMgnB4gOe4jRua
1m9qRXHeQlvwtj01eVk1uf9X4nIgDEYBOC1JVAebXLj4hiEvSANN/TV9UhE+Swwf
PWzxS/rRmLHYru+dqVh0OkMaH0ly6zWSX0/oM89PXarZMPmv4k2Q4kOT3jN6pMsO
mM4ijmJLYyF9YtjhSC/YZMi3EK91idQZoHEu9qmA14D2w7PdgPBv224N2fITMUtE
xWi91EQMhrc6+7jD/bPoBiFg1j6Cm3AtaYtszqRgcvhtLGJks+cVAByVtDIMP+G5
w5BL8zm+S3q5pMRN9GGDxa4K6n+2M41tSOX63Iah6M8RVWvE1WohLrb4t3K3bBXA
AIxgujXVum+w7tW2A1CAVUSbyL25cqewzvN+XpFvXMr0niUPviITfwSd/xSufAYe
VHe/CZPUeOBW0rffRk373TgxcDEN/5Y771COHWGo69ocX0e2ftqTIRRKAE6ozQxY
qoUrfOhhbrwVyGlhfPCsaB+4ZK6yIgfw6HjiXc0x4Q5DFOkTjqPHHv8u6fwJlRYZ
8yt/X0GePsoMsmdAOfyHDMvtRpfkI7L9YAYnPyH9y/dPJocXXX1PQZ24HtvjP21l
dj1kQmwVQWNrv/3ieVrXJt5xNzZQ5VQ3z5aFVFj01I57RBbN/WhoFWPjzXd6wpn1
7vQ2lLX9D5ibyKOSawNY4dl5ST5ppCOFADNkwo3f1Vc/wyK2bB4O2WUm7W6igyo4
qJQkdYVtL6z7sImOBDLTRLfiEBmMnNKg7SxNoQX+YkP8zgKjGzukODUtvYwmAS4a
z738XtxAwHK2yx94tr1/b0+WwRrZNW96eWuWJ8ofYnXruzgkdC0r05WUFDD74sV+
Zptsm5Tfb+BrWc8+9MM6+ZOEIGXc9Hu4npMmCEew0chrju7PT9eyXS4PkEW3yaCs
MooqTkp+QPDfAAYW3231Q8SucJ6KcNXB9wDZxfcCwbPojz+t++zeM3xQULsGazIo
t7vLny95HE1p0vBHZrioLdSahG3E30GZ7SfHJoWlmD7N0A7h1rqhEzUrp02zR1Ea
//kC29TjNN6/SDzbAja0lDcvAoGIXDmfE6H5/cKLBCpjPp4c+nKbctForOkIz3sG
GUzt0UXFnXKXMCdOfHTwcOrKMAxiC+GJKbb7o3WuTa4QcnjFWRjzjbMOuA34EpIR
rBpMKy0RLjO6+YUkv+RfLsymJpn/FKgYDQIfchJnV7dgSFIeGalhwgN64/p/iYK6
wGT7EhU9Z2jHTXgJxvGTFC0VUsQiuqeH7RP4gZBe4pfOYHAnlI9YNhnvZDLs5dYE
RglSUf3x9/lTb6MtpKFND3NgwfNMxARfDPOolaRhT7CQxo+cAiILJDIsslxAdAPZ
VPPaJpkoa5wUqGsM3ktRKUZ9fpOhnZe6IST4TsKciTwZZa5MjDbI9gPtOAfHIdmc
Z5RRdOr5yAp14X7ndl9ZtQTEIkTcb2xTFM9uMLtfUkrxtumYYgvDC79kWSsAOjSo
b1ArTNWW09CKRs8BOQ2sU7Y2zRXvDQNt1WA9fBJZz9xCe6T27ABPP/6pOl9FJtGR
qdhShszT6B6IADZHvGmdkDsITKgfosPKg/JPEUPf7QlNHIrj70lpNm3CQmjfTGRJ
aG/d6LXcXhZKjmFFTXjmzATdXOKX2BCF1TbqMRh91gTeVHpzzav6jFDyhKTdA4Hl
3l9J5Gqz5xLipSRhcLZJ+58wj+ILjgvRzShMqrCrR7cUPIG+egtRhBZC/W+qTopS
IdO8lAoWYFMA7fLI91Jbidr1HU0hwMTZLWtjkFn1dY1Cj5zxCPcWQhW/RO5rQnT2
eXHqwIL6T+3g4mK/ILpqWBreVil4wY0N805RLsn9FjLpvCEI17a1NN0/Iykgxz//
rNVedllzGKTEhXlsMc/13iFcFQR2GraJ/VBO2gu8tYja3JiRC9jf/jAUx8FqW7Q4
q6UvxZiMqzarCdqTLuboe/YsaCjB6u3vApH16qLkM4ihNxs7vBqkMqAyuUgccDse
RM3zNVJNzvzUNFZ8mKMpljupZkC7DmSiCwMutdAc758TgMoEj89W63xh15A3RlHz
mm4imLXouhv3kmOMAxYPO/dYjNgTdYcWcPtAllyOUoPRYMWDSmUKLp6WoFSzFCDa
LtfBKlC1pcAQhsnsYLrhsotSr8Mb0eh+xuyIr/ik/bWUIVoZJLagbBYZxPzOE7ev
Tvz0Xbl8YszqBDogGuAEjrGzdhGvK7nShRBJQV9gMwAQPyNp/ZDB82Aoyk2cjx0Z
LyrTcUEMbrROhpjLnHi3ezE+t8+h2isioZXIn+ngoN94lns5mthIowsnnkslP20h
ZiHOULVVFEkhK0XNT/Gfr27P9fQrwXSmnQFdJ2iJcsCXwDlFH3Sqvt6x+tiCD5md
fzLF44BWmtOyadj/6n15ezU4uA2jRsC++gzjyHzxmDXELUjTlEqF5rV5zqoY7gmd
NcwI+7mNMB6e5XaLdjCFK9CT/ZxUcWuD4ZTsKW/O2RvjY+0nI+ocPIEPjgGBeC+E
E2Tw+YAr5a2t8OrWYx20VvmAEcU7tEnRkipCsBrQFQSBtZtTycV0NnImlcE75v0Z
orPENkjFpshTREXszjJHu3kq/j0s0QJlpAUOCPOHGAhGx8FvzizaVJh2F30tV6Ou
RK1iouFnl68mW6lAMX6gM8lpTdgueNXgUkxZXu8eLwaPYBFogAjdvUz4lfxugzbh
4fvOyK14DA+YSqszjAeNuHYTOCBqJNc7dWQbKWVLIsdLTyQZzc8A3JkhCmTL2wub
wyQ2g3UmvtvHm7kdVp9USUbbzq77OlTbem6SUYZ6IfBoMLPYypUriTE/23v3t01f
e4DjqRue5QmP1rhkVJ9FgNA+JSJeKBtBOAvLlDrWKCU/CJoq3cxLR46y8U4k9tsN
oEC4TfHFBi50GA99DI40E44uoPA8wd7/Okxaj7tu6jF1q8kBy/X28EiMae0t4u+F
tKF7aJqWrNMCpyqQORVQ3/mus+cPpDZO88vvZfxLX7Cf8ttKo4sNE2eEhj6I/4dt
NK9ETRQ1X8KPtmJXRDswUy6Hgo8YTxLwiFBcDUqWk6Waj1O77k+910vF8rohWP61
8FJBBYK8ayvcGntOJCr+MlSTIvxey5tlkUdl2h/2VSNLEqqAF/1IlvR4MjyKz/hS
emher6o4r4WgY9k2XuFK2fyHfQRsrycCoRl/+BWvbLYaAqklco0Iv0LDjDYTS/6g
g/0RmU6flo8JQNa9RSy6sAS+f2CGmOMuNATMhjDNAuzCw0gTEl9JNu4TuLlboJIf
02VaqNrSP4TZV2tpAVFom/Dvpt6a1uVl+lpPs/t9T58bN7PQe7wcMUDf5b8wltC0
Hv7Q+rqaV7awvWltOCsBD8awLYUco+/CnEtAul9dIkTnDStcxy7S5TdMcgM4LX2N
Xx1oSdS3tyHdANRwZP7jQDaje2RYhZ+rkNfTL4QU3ExONOCWWKyfYn0+bg7abSGS
byfm5c1M5svOXM3r913iK21tfbGwKwqB9AkO4uQbe8TsAlRjQ7lDkrPn3bhw5Vf0
nsAlMcwVqGfRuewl26laq6I8X3TJxBOHd6djzejx5kZjzQl+cZABadOO1O9lFTLg
PINFWbrr+GEpzy9S4v3ljvgvPw3cejz3ihG/oT7OjF60ZoffTR/dlgQubF0QT69A
+JBsoKzH23m00cctNOdnfDBQ+toZwnC1YrCUz0o5Oe9Wxv1liQd/p686h1f3cuYR
h16qHYcf8MSbvepRuJBLJz5vKQUP0f06sM1zCnQiUYHNA5zTgHMKNom1F4vOUy0y
L3G4QOL36b5HPH1DpDIQISaBdcKphVdZRr2NCxNa5EQy4VsNBOm6GGSB/yn0yZbN
uh0ccY/LZ/lTRX7DYa/1MjU9dNCBjOXZkU9gHmatGUZVfw7oS2pKPqZQa3hOwoVT
TbDpUirwsk4pGnV3GcZsseKkxVjJLAWoqAx+e0xlZXOgQ0eHn6rJ7+L3sRPG8e9J
6469ZErZwyrqVMj94sUNZZXhb8i6X5VqJbrp5NoKdpIk67H3CMsvQ+iSwmMrv02X
JgKgIVAlGYSfcRvsSbSgED3Vi6ulCM34t4uoAMJtvSPmefwDJlUY1eqfn2qh8E3M
kiGGAin1/3kVQX6mQ5Qtw6xjL4PKO5QpuVer2ozWvXqTFkgRJpiPGyy3/TLp8gDB
F8ODzfIwvGSXL38jlalAIrcyx3XQLLvmtfsn9iipUhmRmrdujMTxOO2jKd61Qfnt
pJybM4f3Q+yKvvtwe3QUWZoWNKY/3VRnVkfCIY1ECR3YVDcMVTOrF7/pIGzsFb+b
BfB/knbrp7J1wzrMnHGWjrKYyp26x7gQwr0uVmbTajw7RMXbq185kJYZULJSQCZD
6mKFR/lyOygXLaAj6CSjAKlZ4Bcmi3QkAOj9Sm76Sqz347B8RWe/q9PYHbNUV2eC
SP/SQRl6xDK3B+q5ois0iKhCYzmjTV1/zdLjn/DpuJSnsM3jHXo3qM/mXwH1IMYh
E9j5LPFr4TLHi/hoJtEaoOzK8AXY8+WK7bWjTS47sK7t1FRnEouVda8IrT394iw6
/iNDeNfnqJEdbKZNZ6/+61S7+DWzeQf3LIn4Xq6idN5n2jVvp+cgNnbvlUL0Ctw2
3VkMKUyq+a9DZqhlyUdGZledEyi3xYv4w8ykvoVpvMdtYmWZcZU4R0VJoYkHXzqq
OosXPt1pFWxmbkG80exh6wXhfa+egOLOlhblebQab1dkDDJovOATn6hmnx1MHgXx
zFYjAG1CEyKp7T+V0XE80QZX0m3G+suT+Zc2OQ21EG5FqM4kPkLeC71UP0mFyqjZ
ShbLcriemEhxJHprlhw+gDgQJDJxVq0SJN7InopgLMVidTN0Ev/Cp3SMthRwLufs
NhhkrfvXqIWyvXJ9Dew2qUqkU0XcHY1SfVK9B3/WXvQZiZA15tkqN9DYMiTtCsC9
6UBJWgkRK8MkXUXuLe0znBudQQY8j2LYSQ0psc4oTTQRm4+05wKcQazo6RNoz/lz
28UcS9ZjLr1Mq2WvgR/85h+6qNR/MZlsptjqH2scycUgI3F3JqyVXmGYUC3CYXaQ
J/Tos14t3OLIt8Pq0+w2VRhD6c+ftPrNXqhR5KmMAtaFEwObmnuhF3ChHlJHj8PT
ozCfZ/eTIV5IEHI5vJaYs1AZKIbOkrgvW0p9wpBccCaXNoXVFVGQl7mbgysVUMGN
g4uOOhSfc5YwC/E51FYAz/HVrurgX65P64INeRf0eMGVOl4XZgdmpkoPrANQeqiY
mC+sM7KoU1nl9RvcNkJrSj+MzB6hviKY8cls3zjjhMBYPGeqleR4RuH0eEQ4aTta
cmki1JUKntBXILUTSWLD5i+ryCvvGB9Es/RBzEja9T4y6VW5Uv2gsihporlk+EbR
/bzB1B1ySqwYnnrf2fvxdIoIIFcCckCgWpneA6U851udrcwyhSqS4LNLwqt4GGnK
rtRzFxo6rNRhiytHEMgS04n1fzj+KMyWOAXsx+WHl7DvRXnHQGWWMjdy759ZKuyL
kmfwOLcNJmLctJbVcyeq+CksIrvfzgMD950UEGlUrBr+cmNS1ztMPnsiqM8WDe79
iX9EdzLvBi4QlIoC5aeEuTk7vf2Jk2BCIubnBVR18pQOSXqScjIiVl6eLDL1UUfq
D79i0k2XFO6l5fLuc6jfaDUR3qVwaDilV3SsGvJn/fBdF4lf/mTsj84qggoVKWL7
WHVrjovmvIeeFCG8nlME8sq0Dt+iYjKgM5DjNh6Rjbr1+cenIFxzIVGqv7mLrya9
g1ZZlUUkL0VTuJS1hYGW14KNmzFwcW5LG2/Q6e1VfwxHSeZGQUzJBmOQRdMX+kjz
0oqLbWwFuWaRr2GxzqRS3FnJYhlHmai9XTLGpQsGp+nTcw+0g96iYN6v2FRn1mw+
F9K4k71i05z3gC7akG3UKjAJKOm/I8LfJZ/D4XI3Dm73xvNMAJWXex3GBSzMSg60
6d4Ct1Qi01kb8VuKnSHBkDkK96eqtxz1JGPfVpZrdsMH6rmhIQQfLNYHEN4nj7EF
PUp0p/RNa+iUjO8iEpbIByhyd+P5TZJMaHxFu2Qs2Si/eyWsaGGO/mv7CL8n7ghs
sadubLhY2skrrD9aoveEIgJgBg+mGdhxjLv4VuC3CJkDiDxkGlF1cSFbAcKlP/Ij
P/ldIb0dC4tm2NaFGhfXjGuT8SwCSuzWq929ugrwGeNne4sG6lPNZbMHDkhfneIL
wV9JvAu0O7is6AKi0EA0XJfFlVn5l/ntQFYBCL3uJPHIY6oCx6cz7NQJRpFSYakr
ZVlysmFfTma10pwUkTcK5Y9xHeNbibsMNi+LGjlOHv4qeNDfYXbC5Oj9CjyE88na
l2fKAqvCDRu5odmt71fXClZz0cJg11dB6boXfcHtIWbySo8/Nd85cIq26xKuAgPz
HUb4ZnQ7DlA53HbUK95iIiBQ6U3CRk/jC5rDRU4bNvctmBznb2OilpML2a4um3EK
bwkyqLRCvva5n2kYJgB+U1kJoUyY9jjvUNdSlnBTcAVWhZ2+K6bd3L8Jn+y+cH9j
cuNCWT4pwCgD8VKJ1cxIXbm4cFtdugl4bc8EnGQQ8akHWka8x8wA8ik7/Fb6PZGm
rdCHl8F6a7ANkWDvIcwu6sKRDqHAotwcs8yQZRVr4/MiwhLRF3pSIY+IjQP9aB5f
U9Z9s9APdjRwIEhONm83in6mVkSZf4/+BsylL1BNfBlVrWcaQsvfzQ2w18PTI72n
mBIqTNOfTbi5sUiYK9x2hzTHcD3GUKfzu+OV7HmwlADZG8fMtoe6H2LV3t+fDBTe
0q05RmXF9vyBpGETXL9eXoQvRQvdzwXn6hLjVPuxFnUyVwrlCFjcYESH1IP7X1NU
hEWLvUWwxcRfP6n2ME5xZUqFCAd7zraQvBlqyAx8aqWhMRAAAUWSCJ1njT61Jq/M
Xcm38WgihaZ8dSBj7a1zyBg9NaLFA/P6YA+AbFF4JHtJgvuh8HpmUAYiVxlzxc2o
6D/vP1mqqqNKVtDv+nB9Xa66z0i0/aJs3oOIY+NSks7eil1G3VvnAh3V+UCUxkQZ
5VSEMVP0YJ9py8oWpYH7ajQFmlQ/HEvR4vFmocqVouL7ZefjAqj55fW1hvxZUymL
584lFQ1NCVJQ5gsR2dxQc+vWQ//C7hb3zTB4w5EmLh67/xaADwM95tIuRYcZnFh4
kMVHOLkGeVX9qUuJOLOl2j1EbgVxEfngxv9XSv/Epwjvy/kqWYwhpGXFIfpGZut5
q6AJm1g1YrbDU9JUw0DUbzBprabGpT6AcJM0dGJusd9Mn2YX1t0ONhaBq2IJW7To
+q0l8odMGmqHVT1VsWn32DKdpMyAVwH/uKMbndv2tZANtGhnYeDGEijG/3YAy35n
G3/I6vyoZXc/JkyX5IDYI2bSD5jwt2IirHjEVQiEaUMSJUSuwHHzAuKbE4Iw7Trt
gqCF8dno6RZEnKhh6REYuNRuC29cfAx6Djioo/s0Z3zr68V2KaM0HdcnOrWMYX64
xWv5gZuAo5/8VDuqWu/yfisHEjGI7yhy1KxjfG3DfT6iiS7AE+IGhMRWQHxSrkMB
CzLH1HD6zRhI70mtHwixW95UKIOHXImK10K1eTCXINu8bdPVacuajzA+i11Kz5qq
pz4/WzVNeO0/g5ta3reSG7q/g367WSSRCM/zpjJTAE7I+sRNWF3+U+k2Sgrh3q9D
DyK30O0wDv60I3ex5zI1Wj3ws1+fn9GHEs3LW88VjVtL+QOLXPLHPbd1RNa/u61Q
CtyHJexhC/LdNb46U+pzEjDqM+wvuBZq1RFZjmjIr5AvdGaMdF0ZP6yLjuWT759D
0T6RaFmOlf8YJIz53MtuvDQPMuC1wcT0A+y2HMfMEJUkPPn04ShO4ZBm2ulGfNLv
FeTDgvxu5U3e3YCA5JxOmPBG3CE5w5gPgvw7vQobt86ZCAYe55d3B2cOpLAWJe6n
6Eu1lnmYr9mPCkmNwAlUV3j3Ukn3YdPWH+GMFghLvzaufotzSfBAMa/+gWh5EJBw
mFRRHBhmZ5hAXNBg7GJXafVC6Wc2CW/8JtC4+FdjjEGehDUopjT2iYaDiUTA7Kz4
2ZfuKjWdAsqf/H7uB2h7JN0GVDvvTngv0tycFYLwZw2tThGDe3DBTwTQZt33XaLx
fM+dtrbYc8awZ2tXIEWf/JzRiaSaF8Ft/PUXSoAN64mLXZm3VtgejQGl+YrP5I/7
7O9o19rmx3+QIQD0Qo33admt3Yd94WrgNowjdEerlLFv62gHB8ItgqY5gO0ws3dj
4awi1B/ZhGa0j0WcVnVKRPJqK/g6+FAmsCZ/XA3fs1W6Ezo0UGYNPRrkza8eE5xv
+QC/BxFtKtjASu5Ie+o9lqrbKwL1olYSgQrAUH+7vhtMlLGl22grK93qhl9jK3LY
dR+fzHHMGg9buVS9U6/P7VcDtMSr6klJ52TyLwkBwCz/Nuw3xnexo8VWkiXbwgli
RlQAZJa1/LvQk0r5GUuvck//gYri76MgI+autqByfxz/tKE8RRO6FZb1xSVIZiYZ
aIlMlRJZtR309ZWqF1JYZDJdHc3wD8MqhBzI359ScABvZVkeSs/MIvHO7CcwLhEQ
mTJRC/eq7vOLjLho4RgGaaWwkqYox6UwAnGeURlljD7vA/0qU3hhEIXRdTEaP0z7
e4Q6bdxvVfXJ5wSjsrESuLUt7EP38VNU6fluWXNms2W3xrl4ElzVV2jLxuqw9VSG
OQmzeC2sLevMCOcwLldMmf8x3KPFOuPTOUqCIr0VVV/qMoIDN0R+wptlS+xntRqk
XML4A6VM5eK3RWIxZg9s5JMfGK2cNcJ95mf4I043XdF3MWaRDEmr2mWQ/Aw9fLMz
RxdbzRtjZ67A2aZIZPuS5nA74LMIyk3DQdeEkB8nn5C8QMmZIps8SCg5TivwzMRK
SwReyNgr7IX6fz/Mr+msZqgl57kkmgI4olv+hbM5avDydZPi8dORhOXk+ZjR35eT
zvroeDYjVNJlmHs1XNY+bnU7b8eK3lzqadSC97wi6ExIgALHjXx3nttNLJFwJ53+
DQ3dCfz4KIgoTWkvqEB+FzO65laov8nhxQzm9VqIz/9ZlN2iJEcIbrSqZO+1XXeQ
wQL4TKKzouB9poudRHbKJY96XYTM7LlWneqCdX8fyG7hpAuSzfVMMOVket8K2Khk
GeXphwuDUaB1yNAI6dAWUpJFAIehd8DK/8WzjFCnK5WeRRr7gvfOxUBDSE1DoEUP
TRehDzV735zCDCOgvPUKzlez8YMcKo8RBvoWBz5TxB1ufjDHCR+bZPmDjO4ZSaq7
99b8p8Xd5Q/bPOMrc7qpLprrL2dYG6D6kcCNfnpBLt7apzEf1WY6+7zR3sdGW3je
W+6/NMUNxmldn4dsmAAvO8d5djboGS+qn/PSk1CAIUpky3iAYNKBVV+uhQW4TYEy
oSeCQMQvspy/31v7Gnpq22xnw0pcY9vGDdn/4N+V4aQEQ8qcOMbJ5/tJ6FAjKIg9
FfNJ8oYjR4rnvS2JmLKK0XR4NGX38xK4Lx4fx4xkz2I71PbKrrnbxpbV0dR0PkYV
rKBW/jFjo3JWW2P/7z0+pY+ra8d53k9drZ9Wd7YZchX1XlekZDk6lChF16/z32tY
eti2exUqnD2ea48KA41eTvMXthfHF+tXO2dvjlkDYSZO9HYNT0euJYMi52KMWY9A
suQejCjlgvVEGaTyAJRBm5PC+5oMKayTz5rv72h+j9hrJTHCKew5OqkdYHbQ2yl+
bgGjT3eDsrlazxai5sDAVgWXnTIHT3p8zfDq4L1p2AVCRzPck9rv9NVnZLn29PF9
D9Fuo47pPKom4d1U265nAm+XxLIeo4Lb8F+cMMPONFRA9dC0Wep6CjF3gvayPhuP
NBLnEylVSOt9o70F5GrqFNjyujYn4Als63RHZZjNj3jtIbZSa21m2B1CTVbC/YEH
ZSKeF7IeP+/16tVkYHgnbMJ1AmhBHCjbTILFH6Suw4Fyy2rnSosS+0LeH1bcg4c4
VlfuB6oDVtZxN3eZsK4tzTK7wL5rqGzUcfSCS317mnLLhdBHbOobSyMnJzdF5uvK
x3YgipHxCkQs1sb4Hm+idQQ5NwajbQp72Zbq/8peO2rVOtDVW//695RjPlFM8ty4
I+NZ3ClZSKxtfMuF+RdnoHLVNzHqeqOy/H/4BrZg+j3PEv2zw6k6oQowLYxvAqqx
O1iKINU0lwE318aTVla8NXC+oeNCkT2OTSiKg/zZE21QUbyOdIeAvDFYhJ/8/CC+
jqEWH1j6V8bHxfxdRrZcU8coPDhxwaehsc/tUlJd2AvO8EocyYbk1OZgeutW3L8r
D45EFQBx/S8fL4khawDRGonb+swJeGB/o46ZFOk/q1k1dyw7+VjgsWcHsTFw3OWe
uMF14089Qxa335YAhwHVJanTegqdmQ3iKyXpWF8awFcnB+CIoxpfven2JLYXA1jf
HUHFUKnsF9Fh61VicDqjJvo9K2GSQ5SM+WL4+PKh1jczwo/iO35hyDDm69K4CJRw
OvhEQC8Nio1KMXD4tznRmPcD10meQsP2p4fPqUkFZ7NJuvJ4cqWIhmiNiOC+gFkH
1Yo2khTFf/mczxrGw4URQizdnQDw+KRNk5YnKS/ULt8EY1rVtf1H2Z9Z/9N+e7Xp
H92ThRcbbct5QgMa8UwPBe/ZH3abAR2XLQSDSgzKlwCbiK0pKISwoK6T9OIF/pZ9
B2YKt2Tky5BTQ1Fk+9ONG5RqhhLwRO6u3cUegfncw2hXx7Wnf+2qHR5TGeVQ47Mr
kmXlF5UuzNJcuppX8qUn35kLJJUbVkdvzK3pp/qFYoDgfRf5c+01HA2OOEJUZsZh
XsfaN4CytOABdEpqLos972/OnEkaXuwGJwOgyar3q0eX5QH7inFSy8S3oo2QxWKH
VbkXsgmCnr2AXsk8WTlanlrR9JEhd94yxlg6v8V7Ml3rl71qlBnEV2ogSie+K1iV
KAbdD9cQ+kPd+ROQgqAZySj0KBrWdeUmCrheRnhHmFcsH9nBrhKOHpBWHbqlLG7o
GA+MqQUQrNMCpG0hO9KqrkaxXCcLS6FMhCJDn+CWpV3feDeHcP0aQyrl9KBHdA6l
VOxop8rpEtOerCJ3/Q7aTham78ZTFwOHbncQF7KRo+piCNJ+4NT+Hb/HBshGt4zV
ZHHnUxVNF8ETMzNAHKkDFhLnBCRUjYCMS6NOjDIM0zfwgoFgurVdxh14WLDXXm7/
7YtfHFDy7YS2WwMMZqqsb086I4CjyHXAK2638XblokNLd7btfIEQ42w9igy5cyAc
gOIGu1P3EaTkRHk1sGVszRcJxw4uQQBIWVrwsO8gh+WWJjrXIWCOxycafOz7gVXE
T4jKdtTYFwl4fvNMGkZx0feJlrWa/nk0oiMb65Qqp7HEmDX9cvBFQ/TBHGdhaXgJ
bo6kxcAD109teAOq7Z+vkyHLP+06bD5HidYqn+C1ujHVYwJ4y6BRSN5ub5XuQfxv
gsgbXzFREqYVDxE7InsdaxL8Nteke8mUZhXrUqh+nX1dHE5M3cnZioPVAYxibuQB
UciZvO79i2s/8k690Iq1uzzxD6fHXEzpH8rWZkN2nFosNFvK4akSV5oUoWhNzrpA
2axRnyrHneM/6qZ/Ps2l1Ajy/xtNUqjLXfNXOsKF2nTe6jToXLUKly7rtlYajX5y
ZYboKw+kH256Bfs8guGrcwOnXbfx22c3lwdGRY/Jykie6WNQi/6yS9JgIXVbh3Ph
+4ycFD8dYhk6sThP4RcQIhACO5BcM7sd3mEUXvTdHdkO11vRjUSfErwHDHHovTb1
/wtfktW7cbLDEuMYYaU9+3Co2m5b+iKAgvNt08ViveuSpAhA2N/wv4WeAykzgGlC
70RiCx5mel6IIWYy8Iuyjm93dheM2+8M1j2s337qEXDlDzMF0Ds8Sz9dnRhhPcxI
PDuAmy3Adj8LVor6CBOPshvVqYFcmAFmWy2HOd6/kjGrSeemyBgeWj73MuJ4CXZ7
Q1NrWpLic/s0mlh6/W8E98d+w6KTfSRrxcc8JHEsi5uYXwun1sXH7sJXLe2K+xje
bNHFDgQPzoodzgG1kK1TBX9eC4VG+ztSZ7b2fjoKbinMfbXfG2+CBhsXmQRmFRVG
GdVsHxZtCl5Dx1gyUYAfsCi3yOjI+QlZyUcL21gtWaGu8ANhxi2eNE3gBU2IWq4/
FaFWj+5FrPxfP0n3nW8agr50vSvV4qjOCsu/Bvy7eW29g3FHBbNuVFqJ5SeyNLxc
gsQg8hsXKMBiqKnI3J66gVQWROAl+GU+tQYocCESRvdoUhqyBp75seNMyFQn5xvQ
WoSIFsX05BSGQbL9OEwoY+ZXFFvrT9ItEDqVCnLyJ+2EgoinYPdsoYRzF+/wmtkc
ZxgCw6CuI6We5VRtsx+Op1QdtbEqgmr16alrnMlhzTDe6adDeYHY5m4WbzVkuoW+
rWze50VrXvl2a41nXsSXCdoDnSc8r5OXeX6HY4OObOCILm2qJaXOCDIzjtyDYJV+
pOIAKIemZu6tcUjIYceupjBoLaa1+o0Ev0vSQbX4L0dpEHNYt7Jy3oRWDrNZGZc0
szdpHP1GdB/ZjLFaf6fOcYf38TkODL3Gga0wf1ljbjnHyYdeSaJHWzkz2WLhKRbs
H44YpEDzwKao7byjdVc8BzfT1n2xrL+PDwPx0ZOgyrXY6mlLp+0Z+pOOMFVBuWvn
t6ixeJEDBHwz9tHQrdZsId5KTdLmrvKpO+Y5PDlN/bGmqmsfmA6ePdnbgdVuS/2P
Y4ZkpJbgu+qs6YbkC3othLNAOQCrytDlxOZnPdnsXIGWzte5z08bg5Q4nCvCU+Nu
aV/pkkdV1aDG3Z9IvbGxVm2DeB/znSgakDAEgS+cs9YSrDgZDcVNQh4OODdd/fBN
iFGmTSh9+8t77+132Ud6gUjpA19lrUoUg5yJcRlokMIgfycibJ+kAm3/oLdjsXwO
bqMs/icokSQPgVM0DNagf7J+9yJ7YJ9OG1xJ8/V4icSU4szetomxSLOT4GkXJZbe
P13r333vZtgUD47kSpw6BQt88Uo/FQS+8YlhHw8rVLXfeQtprXiP825f1Q7QzaQN
t1sEsspGwLF0fo9vccaBTtax8RoUPIoVMjt1IGBCaZHjuw6UVsbbDq06bRBRLMD9
eUmgvHmZXfAPAecEaDPMwwxzTqF9hAVI4lB9zVVb8Ef04fCxRwhRVAbuvmEoVpZQ
ZfbjSSo+2y6FqgRdkO1KPo737xCOfKsC3EaHT9jVYe6WkIxo8SlKLuG2ZC+IM5RY
fWWzYYhr4cJO7tKdUqU6CPmzp1HvSCKv8lCiS/QXwRaQJEiOhHTqnz+GP0Khjz6r
d+78y3mK4adbjqE1smoOSq/69pqkLexvO/rJlMkNANxh0k9hnkXJ8462EompncBM
rWMN+TEj7FzPkKHpS0Ocy8M/6iNq+91tuJba0jozmw9Z5KE5XszZmWHN/PkYrjkn
zaAHLb/xXX18LWPMatYkBlIfabOGpNqJIMcahpHAWOky0AOnIqeCNeLLyUZH/ojo
bwKh9zF/O2VkNY0BgAvOb0WiEUsUG00L+EuQYMhSv7TTQ3+k9I3bgt3OWT8cEDiE
F6MeWaJneNbIpBcGY2MTkCwjDC29xQwrAECYvADuUEf7wqFhZEFDZLI2LyZ+OA8S
d3dOqPtNtvBUNZV9/Kr0SH+xO4+kGdcXjl/sf8GLa5iUvRLjAbVcVH2eM8dblV3h
pjNrc4PUxQJ+Dp00NgvpzVNpEWzhl/3NqGNPnIDBZdi8oknpQd3DVEDJAFM4Z47a
UMyMXUgoyQJQOxMO1c7snrS+jzJqJNkypdfCb9k6pZWZhH0vWWaYuQSefGbolJB2
yWIYqamB7Kzf/dgYgOVbwj7LConiy1BqryZcUHwmMig4fNFpBO5NN8akaiFtP8gQ
fPM9OoKh2/3ab32CpASu6YiL+Acc+RkCUozoYCm4LdPPU399B1fBowFb1LOHEgMP
coFszXP7a+fzFxrSbGeY7VlOeAlMHLh/9Dx1WSKaLZmBF1Lp1Od4a+SU5rhdHV4Z
HX8ibBWTmD3hhp9F/NQnLZ9Vjev0mRD1pCUPRCE5lu2x9ScycTdwvbok5Ce3l27u
OQ9CpRuwr/swL+jvpVln4LsWW96AKmSd0W0QXXmCTyDVUVuJ925uYlnxTGp6oRie
7IHekkiswnZ4b2kTGy/Xp0WUHqAogC0oxgN4yxZIHrrcdy8qGP4jNJKvbMHnYwdY
uIcgdZIyQnOs4cM4hK1TH5Xt2wX9GZyioc3HYFp6Z0dy2RYySj05emE86EOk0HV5
CLqO571CrVl8cmCiRjSdQYa7mqBUVoGWDqpwkHMd52E3Op+16HHdK4FEn8tCG3XE
0+d1uF+697hdpdAzU/zYBK50ZaVUio3kN0SnbpSrpfLrSNvTXrzo+QLP5QemPpNZ
v3sZ5bo7S4sx3LZr6lV6J6afDt6VEEaxiYfFutDxkv9wLyIXp5gCmpnYas7lwqKd
OtUyjePCEY69BaHD3nOimIVGLedpVQLrOdcsNWPpXZtbaRt6Y8gYuc4w5Kl/lstX
8DJhQDW+Nt9P+5t+IwVSPDtMkgEpkxtY1VAl475ufUwv5PNIN67mu5MnCky717b7
bDWF4Wp0vVd581APsDAZanVyWOiGJ5JkvTTPdx6NjY+WMgzS9f5xsrogVttUm0qU
+nEvlf+KM47iasmPwn/41jXro89ekBhgb49jEDofc9wZgjtp5FRxiua84Vnv8D8h
Eykx84ag3AJ2hv+uyxNOg8cbSJwvC4dk76eYpo8hk+0l2M07g5bxkcjMSMdCVn+h
mWYGNeJzG/so256RQTl4mO88EjvB9Gqr6hcaLw+HlIRY0nSbEQjqMbgCDh18O/uk
6ZhSw+DFDXst0mVhVavdozOl2MaTBDqwCYjsSb/nilbBq+LD0eawJe6Pr8uFbZ1T
R/uLXcxzmoqOzZTv4PIXZHLH6nBQjSfXJutQoUG7gNL2GASrFLYvRyw7+euau+js
F2qAp58fVjhb6+shJN5lL3TMu12j38vii+5hkFIZSQ5CPHArWdBgQNQk4n3m7UpM
08lBvcTPwR43mYWM5tBBgplhKNQvllm3r44ZdYeFAGViHJs8njDeTYUUViUXaWDU
+h1pGKjnBYhgaeSHJQnTEysRnTN6eEMVQfTkCoYffRIRv7Rs7aRjqvzwJAFSeSoc
tVPyqCwJ+BBxAQmMUQP7476kp2yRDg36ew8U1E/T8ikPZ6DM3seYx04aPNRmNkYf
rLyaq4YHe51t7hssOGJD7ZcYlV/Q4pKyonLVpFOrBfMSKBG6iYLb3P1DZItI18zv
y1yFyS64qRmLbjehvdlqNFDsSDf0e6vJCK5/WeRhqs4Ste/usbhNtcZEQ6pXx8Tt
QLtlSYx52TqhiPblLxIhN2UHQpHrMmPRWjGNQVbHzjV3jwceCyodMJfXpuXqnHjk
entpLXcG1KFDjM5RqpdkMlmBLRd+W0NmBJuGSqS7v/Dh1pVohxI4xnqfqDeNa907
pBBcmRlx1sW0tDyTpmWRKeCg6/g3+k4mHPbBAUivzrvoh1/0MVUzGYV7tLpEmTlx
hxaeLGwAuLGl1uGiLrnnzwimam3P/iDSapV2/atkrxfiYjod3QJ90ptYwG8y1DFn
puvh8omaEHv5HPmfuxzCGZGp40vT4NbcIUPyyS9d+nlsytet0X2pwHTKUhmMYl0I
Wn0ped9d4nd54uf65GRLalw51tmL88ULZcmyXwa6uegFqJkOF0UwZKTMorc191F6
kbsJsPAWtc4QBBOdYcW8ItlZ6oc5NA0oiQeCI/IFZSd/T/N26NwUIoixJERFwOjy
i8dUWqKUf3sT0Hdn1NZox5owcuJg/z6JA2ZEVrogoAChNpJC3k0UrSTDTNkjpshv
CsZjElcjn288z8DDvR3OWtW2yd8nf8AJmxRR7TX4BruM2NiAgdsFh6o8ijrnbZL9
2UKwwzGhpK19JOYDO+gSiGdAsTwJ7o4t88/7KEFccWTIWzt72EDTHzniHUIRwK3m
r6qJde7fUzet36NNV07v0klDQ6Q+JRvU/ZK9uPvdrP+vwBZSqSqv9HtOtZJ2ja4r
1zUlJIbX0ZDhPkkZl8JzrePyKvkKdGV4w3NR7inpAeHvbQbwqPJGnUdYEPk4OjfQ
68Sy8r2aJCcDx5F+zCpcS5/h+YDrW8XB7HG03mJ7PdU2+xd8IemqpAHqPoOKn8dZ
Dsr62qjn6R/wpkMv0eQNYm5Y89EVHCVxi+23OTt2wSQKxsFutmLsvaF918i/jw6I
XDmnKaMLU2uDCJknQFfYhC99bUfntLXhyldO5qWBUYErCWJ4Y4RaiukWOk+sUrzE
f4d1aumsrPqqx52GnMXeTvNEowbBOlJ/H/MimcS+SbvQh23tekdVaDofziOtSP/g
X22HMlK8o0nLCHhJOsjiOrQuUjmcrOl/90bnDtALdNrqu0D2fV1tpURb3ppr4aWT
XvlPZn7wcq315j0YmYwJsNlFseo2ak+Efd+r3a/oWfTV2s4C0GPNqBhHrKhTkzI5
ZWczV0pJgmjBbW/cXaYeupb/MsgEDocwhCFf4CJ9h1lG/EDP9YDQrpUt0/Va5Ph8
t3E/BcZCLe8+gKUuuQEzg5G2y3M6y3tWe5F+1Q9XHRGXc4rAU/QGc4b243faeQC0
r9obAfFGU0PYn+umCTk0T868+dNptInyKkEd3hNL8o3kWS/mF6ejbk6vm9VF7+o+
ugp3Vsdr6ZshCFeuZXgXYskXhB706d53lh0IchL/eGcizSFg2Yscz6ohQOXB0kiP
cFNlpNhsH4aFlzir/3Ig7AhXmfgMvd4/YfrnyhBEXolBY98NDM8Jj6N8n+vJDnM6
khhR/DWhnGcJQptbczyQY/KGqQ12jTNrAH6Ps3SK+VjIuIc1g6w3aNFGcVsXD+BO
+e1IWKeT/8LaXXNuxYRfiwxM5eLljxSer6pxgt/H/MyBnJJnuxQNw7K40/VubZVl
BDN5RDleVcDnvcgJHc68/qFL5Jc+wH9jr/5D/dZvbHYwRj+AYmH7+sygcatE/Tfb
uj6Y81Y5otZycAH+4NOm9qHf0QXSx7sNddwNnwiPzDtkMbFeClbrYBZFTlG1SvP0
ilDylfcbJTj/XrjF/hlErKH5LNmBTJPb5QtHELU6ruiCGJXR9AxGXanR2fuvf9KC
QZ/cZTPlLUAjwuOYNOLcvAYNhNBUxDvPPZ/3knoxy6olz9T/Ul7DOs0myXp3+nzK
6ErObYy2LFrorCVzKa+jJkFKky0JculeIEkWnvOIVg4xIVUXYkDlnuE6j6nG7/2P
RTgKoQyF+Etu+8wILmehIm+GLMhrN1jlWlEPO9MxEwFmtTyWmUFhQYasd8ZLejkf
yyKthb4NRKKKciMlhB6RPcrMmAd7E/tWc2u1G+z9xzNvu+cv/iyHW49YYzM3SgUg
Gj7KVG/f1vqSQQ7xlgY7rRZiqoQlswmLQ3lH+h5nvOGlFAws3LFsP1ausEEoqQC8
VoIUIciNJsa/BK9D76QsMuSrzn0csj9pY9eeAK0X7qUu7H71VN11tR/coYvREySF
JG/1F+/2vrwR/69r4XZUZTOWmstnF24t8GMc5KdRSjNM2L3zJkcMPlKD0e6PMWg/
fssHougkbcde36gOKBIYdVAI5NE+0gEpSkixdgWWZQCo00TYUfkTNXTbQUM9q15U
BmYrYKr0JsBLfrKMhbYsM/tHEv7hoYlN1Els3C5+1MuD4s1qgdNO/CjkTkYQcIHz
VyOFEOzFUd07WUe2B39dKxMTt6j0hj6KAJyC8Kcdt/eq0YoFFAXB8xQjU3UbL4An
34QFadp5JaHbFDbG4tgDBZaN3Leb6rZUxXvVLwWmS1Bewh1rAvlh+SGn0i5goXe5
zbW3PAivEOKUG3FYZG3ex9WAK9HWEmTE6K6fk/AW93Qo/vYO66tDG0Isd8fffnYU
uAqeXOtKTz6bxVNo5b8hPiGTWlkZS6Pw16g8D03Qkup5ZDpZkMDSFEdvju0jjsiA
oXRTH6EH7zB3ljmtgJuQM5lhE+9AMeCoEVDumGF5psHV+JMcDOk/Sdwo8ePJpXWI
ZfoBrSRgWbkDL8NX0RolDXAQZ9jaKafUSoXcKinKGHEe7R8e4xXu3gb2KzNqr5r/
KqFvnPYjBaVPxRnYaJRn0iktjbHX6aJfz4UTmLjRyZoY9gO871FskTgRvgJBuy1f
1WaHfeasfdWGY7l/db5aduh40EAYbiMYZ56iZ3XVzeL+TPWV7tJI7cFbRYtnWUWK
x7CXtlimOdZdJhwN0t5lOm1uZiBXfoUc6g9YYMYptu1QrYY2LgbeWY5F7siSzSxh
nwevdWnG9dWw8Ak+vnzXPkiGCAqOV2XxXPpmxI+D9oKkwUW4OS57wf6PNi/ZWSTU
kyS4vwfj5g6JvNO+Acd5f0E0NxgPrz5K3j5FOvavKVKEOozB+RvRSYPTQljR75pz
0hGIbrDSoMTv0SmWJXKZNqlu6/eJPYMuGFtlMvqoopwmHbq1PXQlovGxELyuqtXT
d7gCRCtTpCV0YqPOOj8poit8XR1yA7BdnV7NszXFfeep7r9eRjVTr0gusinoW5u8
GNqlFHPk21C1gBvqNIk8Yr7f3dnErQmIRlVQLG0gqMiumuuTDnnSEJBhL0tz1Z/f
ZjMz+seY958XmMhhzSHnwYfrR5a7dOzLRLeKsLn4MjSAmwtUkq954m02SG9GfRhP
6erBSWTmfUCVMV9ybtvfg41Hxo8EDxHWnjeVBQUbVvLPVdk4YkWRRAunP1a1LO41
bRsWqiUKqix13UGAvmWlrsHInLmhQ/a7I2jNE9OH9Dg74+8j/euL5EYqw7pFd0DQ
k4gBjA0qPsTuEoNEuONO5vCkXUVC8JChCf9hWnZU3GXt76XH9RNbiDsZL5+pyMwW
sleZ5sDFRlKapEQ6SEtaKW5KeQsjjIxE8EzXnu8r4UmvBFqWEe7UrsoyxNYq5cz2
ITsE2yqtJxmT1FN4Oq8hIhqrU4RbRoiUGgnbCstSvPezTxkKatQgDNUb9k/TqCbF
Cl88AMfSH+rl48Ht05EC4ZYg+c7seTQY6TPiWzYiSwOLbKamcajLiVL95M8KrPyF
rkjHflmsqLd5oKJEiNDTpgU+nTYJLQcXRRBWZ+S/L/FcUctZQUisEA6gD7tqdtbF
5z4egZVHAd4E0Rlya+kE3BWeeWzw/S4m0u3WopHMNV8rjMcMgmVyUhNbf368/eoZ
2LrEhV/b/ZLrTv0CiJ7xpZ4pi0x7cW3NV+93yC9kmRVLtANnu3yPTNW/HzZCTWbJ
L45WBRc5uqKsH15mWq9AjMSC65/BqciGt9MvEd2JOT71CzhGzvaD6uzNmFsPTSIv
9VUzFaMgx8UPpNnz5w02et5UzcNPQIwWPm3j4vXRMbF/ayT2haZ6Bpn728lElo/z
b15ZKxsCNO1ZEyMuZi4/W60/JQQNLYRC1T0Q0E3W9XYBa+anUOsiRo3f3y619xnT
TiOi6QVqH1oSV2or1zQGFj3cz1zUwPWAJYDrurYuiiFwJEmzC2VuPFD7upPCGOCH
KW2RRNMOEjifWgGEpmYsGCj1tRgRvfHx16DaD6NDLmZ3uYLexmbqgwccANfb2e1k
T+xwN4C34n4VhDwKXYDkAOXW0DX2KxAVP1zfYBisww4MUN1/x+6D7KIwbL1VoPcz
C8FfE8bzjP+xvILjXNL4Fkgtbif6VA9t5pHEujZd1IyHThjg0s5P8ioqhDOQUc/Z
63VEjlYgV5UtMZGhee5ypL5g+NJceZWjX1sC/D8dWBFxdYqiEv3wk0abcJ0o1kS3
G6tqhNBlUnqfqWIGpZfHzztquRy5DEKweTjaBDb9BKpTPW23yFkzMjh98HCw4FD8
BnXJ6Cv2PTzEv31uuPaNr8HUM689+x+W3AyVYF3LrF/J+al/rNqeJitFk2VwOUKq
keF8+FKtw5yOdhZ0m9gpWEw3OXnp/aOzbr/OdHwa9TGqfPiRlxt5W9+M803TM2t3
8WAI+aHLi/xb/0zGqNtyp+DQXs0I/paxdlEIZngTd/F+sO5n5VouMly4o40Hl6DJ
LmP+IP4RLWxvTtYxfU+Icd60JWeNsZeCuvWU5qZkDEkMy7wBUJfvnhmWxoZfQKCd
kEfRurFMEvnbj264p/d+ZDVXMtpKBT9DjTq0dptHbq4zkC5b53zEIRC9QW7HyWm/
8IHIJIW617TltZxgaaAlx9dxc2Leiwl35j7RLsCQBR7wUYi1ukkJrMMkMqTwRZF8
iEfDJVt4GOhQ+wkRl04oMH6Ccwe/85PXsNYcW+h7bGDpgU9kWyjSf+sjw4CteEff
hhPsCz4i0mgRcl9XZlmHd9aZjE0mPptA7V52BoshHPv7p46wkdPZqku34mtlYrbc
LjH8RYFEYiqjcIyE2SQ/9NpEuJYzq8LkQyeCOytpdOCyAOJxBsiPo4IFfiTTp5qu
EEMmAw1lQlzKu8ycBQ11qx8Kf23gAziXkU7gpj5T94buemQBV6oYjc/vq3YMZZEc
Tr9aAXJn6sY6Ng8Dd1fcGBtYFXssElmUTN7CiuWPuONdARqzUEcy/9FLkGk49VJP
wznQGe6tQGCq+0hKW8JDhcsXHgB6d7hdZ6uT5+lIpt/b++fSSbT1doPcPr46xlpI
wIm7pej8vb5k9rL6nQEFzaWJrX+sVrqb8eQDJe034eiy9mED+3G+mB7FETKzOI/s
t7114k6jRcTpILXMLETxONrCZ4IDTzJvAzDFrQ0rHZNvCNyoubw2TQklhT3LwSQE
0U/9PaZDzihs7lE2nFkV2l4oMjgKPBwEJ314m4+PVrevLuAnUgA1SYIV56iKVgg4
BbMbl/pm4jOlKC9Ld60wuWYSxGEHKAxwyOvCMVlgOJFZtDPJWPLX+iHF9PNpx4bD
JZGmbeIxFGL40m37ODIFbL6ilMLroPu06VxEXZVtPNtPfcOhRL2IcfrxjYzzKBpd
ZVfk/rE38M49LIqueetk41AknbTcTuwPbnPsJmj+HbmlY7iK+gZtoSXbtPMc/u3j
eesJ/BfbWRshVlMFZy7Z3tfAR7t+OFWTsFclY6rMIQNGKWgOET6A4nlMI36fkD/5
k4XE5LtUZf97PeioTw3gVa7Sp2RvidqHRucVkyRK3RpbSvD2wy8b8cfcAxVidYsm
QI6HPrcbxx0QTdKAFUxwB1M6SanfqoW0lDHIlL9oJ6DZsUkZyzQ8tjF1qh912BmT
7vft1hEuKIyrJaAOe6856sMtfjevLsLYncRThWq2dw6/uPX/Lvs8gDLvho6ZynvK
TwMfHC++ywr+eJcEBk8DUU2my5yA9aaVJPa8owlgdL1FeT0KtWhFRc2ZJtLDvgKX
qP+ePvupiJ+lrCNUedO3TpY4Ak5U6RYp3dQIhYk1rzPOnaKe+hdVokKGRB5U4PBN
tDn2U4bF7onkB6dmnIWMWoGIyTwvUn561VGxo1WftQZwStMq+xJ9pugPyV3GuSpZ
krZxB4OBpLBxjCIljAMZj2mSzy2gdA1hk50SjwW3x8K0cLmgLM9xlOmD2Gb1ZIio
2xVjnas5Pth8sbfyWNsg4u3Reie6/qdEjg+AMb8c/ZsuBjQwyX2W0Gu94EwMyJVu
3BawelBOeww8fvcAcreJFxV8f3wuDU47KRLmUDW5Rp6z7slQ+Uj9HI8Ngh9UipD7
+h8mmCfufiTm1uUpEmuW8Iv0qhKN62EDvrOvjCd4wYBdIPs7CuFsZUE+WDAAUUKQ
32kBUePV4nW5ad/pkEdVdWMkBL+Nc+0mfpun5I95AFqEGSXi3mARQjr2ekEhPQBJ
f55c9Wy768nDOppsL334Yx1iEvLPO8RoaozfM7iREGBTe/LX3VkbinnoAUoWuyo2
vpZ9j711jMkUzFUgrFNeqPxYJrnGkmD9L5dFP1gG92WPFscw7Cpwv3QsZXgbeQVL
Rkygis0/v2V6vxc1bTr9rY5pFTbspLxBB7lV4uDUAFu9cggGrXEJVgqg6oQ1XVYG
yUh+28UZn2T5+FArBHg5JFFLN2H5WxeacfuVRoCkEv+ij+E9HQd1+CWuRRZ4PoHO
SlFRbUFaR472K1p+uqNC6jwVGo6Nuowzp0B54yIJzmqIClCb73bgb3trhZOWt6mG
0Axg+ZcZAXIa5OBKZcBWvHBBTLhjEb/ceHv2Wyys5P/Xzo8owtEPijQOQmivbq2t
K7Py2I+71IFYKhN1TjcP5F9HlSr2MUbkzAjyjPNc80cLEBLFJOrRjIHDMLLwoXDv
qiM8aULAlstb3Cgqstk+y0dAP6m3fE7pJZCHTaU6LdOj02O1+i//OSTyyA8LMnOg
oheJBkcqRCgQPL5AtEgC+1FnkTtisjrzu1K6TidP8SBsc3CtZBEPYkf35yYm2A/d
tDEEHb3nlpWPBabhQZpsB8TEGXAXHT1TLPxvJ9rpYakv9gkdz+5P+qfHcpA/m77I
HpL4yv9Z0Q7irJENy8yKtCzcZ5bT2rc5iqhdq1oxyBx5hNCm7qA/cGn0HdeZo/7A
rtMCaQ2dd2xyyr56CjGP+vd6Dcn0HdGpTffg7BJ7HaXMejlC2/fc61L+nb+haVXV
5z5qi79fiDKnjvm39dMqWUeJD40BkRiJTGD6FOPF3CZ0BPf9nBtF7iWKYDJ91SAC
ssLTkn8IAJVlDI0vEM+P9P2MNM5xg+aTLMrzSAj60unu/M/aN5DCzC60JOw8P9Z6
WuE9PmUgegD+bZrPZ0tX1kdomlhc3q+aqTdNsPuk8EhOIfzvKRubxUFYPBOL8dEv
yE9tEOPhTgInLvl/FkrZ/ccx2cLESJekT19+P5YT5lmRqd+300DOMPQ5BJo9aaEV
/wjUy6ClzNGtaGOjz7BP+6YizmYjDOZE0ZYZzpIYKahW5t92r+Z9XU5dEZ182FhT
RBwoqZNQagcdpd8ZWhK3+z2JMsPcgmvrr97BXJGekBSG/61S41RpCpQ+JEpe/hZ1
7xdh2Si1TMAyntJRa7qy/A+4ugD7mcQryrxFSrlg9GN/w6y0TCDKKU0BF5tpfuf8
tZAFCqAlKChFb8I7ApZU534t+Tsv5QE1bZajwlW4+ultqOk1xg3rZJdfCm1hGCw5
Rx+GT1Rik82ctYuxE0BYULWzQQVmmS4t1eNPEK8ImfNq3ZBlKslMXMidEh3eRtzU
msXGmEH8ToqTruie9XJgT+9WMVHMOZoMVvecPM0uvzNEr6Fwb9apt/TMPTT4iFhM
axmLP7aGsXz2KUY63YgHvmhfrJjtO1sq/C/e64GrrD8beVek0uAbDkptk9OVmhFi
+PN9sqygursnX0fxhDG4f3tme9I3DI/sOMzSYrWLinT4Iak6SJvOukvbiCRV0cGJ
L6deY9EcDO/aB1XyeD9b8zTZ7nxeYag8r/+XiZg3d4i/CH5kamHkccke8QtlHM7z
cqpnatHlsLAGcclUtp5+PAlVXNq6iFuFwUFvnEj46APhNlSTiULVcwM+i3oqvim1
uSFM/G1WuHpmDioGUcnYCmH27TN+GFyFPVaBSesIr/YClnBmv/SFLxdsl23pGZR3
0vLJoIGtnZyoiSH72J9cP1hH15ir6RIBhSaT8N2O0y3TCe1LjB8HvA9ZHR+xhkFg
fQPaAF+JOO/nbiy79yPj2HHuyn8UlRPU0a3qyldEfMhXrKlQwM5w1HAUaJzrDK3o
X5YdqcleBmaE6/QrUomX6+R8pHR57uRqTpXW2dDzPoZdFE2fvCJpr7Uhcwe2hfVW
DHOZJazvHf6sEySrh6mLIMG/XK5pt928+8a9kAk1gj8X4yIOTUncoRFlcKGTIRjA
283LNfJ/95HwgQ0FBjNEz+ZR2Zvs+AugY6nPiNxWOrAjaG4oQWsfH9xWH7feNUCU
/IwjoQiAQMp/uKBfsU308u9sQjCM9ESw6Us6PtgGM/3mqxW02Fy320UMDQ4l3W+j
7FH2BVy3MnGUwfRtaMsNosB+8cTQKFLE+AqW0IqUxSfk0/Dqw80FyeGWcR0TJkDr
JBkeggbmJQuqtIGJLr0u39l5HEs0rtPBMZrqk+hUo3rf2Glrm+b7jkpq+hHESNta
5gkAV/j4ibPFaDw+aCRldUH8d1CeE0fS8YVSRVc29WE5QkLw+2ZlzX42XK1BUcPV
czdiNqbiG5ckIHrR1GCYZFrx9DufHbt1oHcYjBKQ3PUGiWAKELM7fa7b0PDjKYrG
l9vg6Cg/RJ13W+NVhDLxcrJfzzAwSNagG9kp/2w6jPQf+7pE4Pr8/EY2F3+0EZcW
L9IYO/v+ZYwjRLTn/LliSgKMuCFUI6KKYu12G9CI4+YJcqFSSrmrP2CjjxI7uFnq
GNlsFSpStuRUpWL39jts/qemqfI0ZU0tubRu+MOV21JIrlXSojoBSI2ELdQ3Tmlo
YhHZzmhbyFLmbLLIlfN9wgaqVK8K2X1OF//cKn+DAJpBf5NnLKvg/vMe49N2IU2O
juEZYtuR2oOBIoGAiKO8YHMLog5tKH9RXmz/hqd1sgq/Ug4eakJUfw1SIJqNYCjW
e1skrX1z0Ccpe2Gg0p3H1ZXSXxnjla+TQl335Ljld5lTHqva/mgogdoYe90iDyse
a7CTNhl0gsxRIA3fAP5WnQucLfHZn3KgQL5iCK4xF8c0GsoTahuHBLpVjL3LOa2K
B+CdDiLS+ALS7m/Re1M1nLfEjv2MESb5VhPAW9jMemtIJt+NijtJGKdkK6hc6SSQ
SdMfYdSePS/53ppwwryF+lWayov5UPr4LWsoEhrbrdw42MucflMcqqIi8DJEgwnY
cCVOHZuBpSU1uKX3NlqsLdViD7jCycLOqfqhT2nZlBdUCk5xa3xJZYkspLtZzpDs
Oaryq8bf9zLbwqZNi8H8VsazRSjVxe4HLN2ScOXdV/JWvcvhjvN6EHyYkhyZh5ah
2G2zrM0OyhDfIvGvTmN3wGdXdPftAuXA6kdJW/h+6Fnxiagn+uAKLLB/tSBiBl1F
eg1bKhRoHGSqB6YZSmD2lSNPhiBV99ILTl/gD7OHwdeyQGSuNHNd02WYNhMDgc+H
fhiw1DVmGu0eHkqFw+P7SPpvMAzT8ZJz8vBW31tNZgSQW7kt7eaM9qSzjEFNyYFV
uyvhYK+vdr1D6YAmArfznqlEuxAVP/vU9NP7jD1OabjRhEYvHE2FkLzte2cLFn2M
QUqEWTMQ/hM1O59T9pfQCxdlSkubhKmsQDSC5WVisEACQ+U8TbkYiJpxf5XznAiy
6bRTKSRDgtbXZfG4uauQGt2+p5g4u8sl/nZ5HsNREFXbq3fcC06TSDbufJqPKH1j
OxXcV60lIxihuu2GIXUe/RB+kcgAQ29pMrcoCVA+WVJrtM9qmEg/+H3AdymHoMzV
QNtVXYuQG78r2JPKUQeiVwYnNZFrwV5oX0bex/gQH/TKS2JDWSSc1k2GBcw2n9tx
BZAIRSEp/S0EQAXDlur+tRN4s23fjEWLI/zFvqHQIjApwypzAk2zul3NrTmgF7My
6XcXWaAJLH6NNKwKqX9Dm98Lnarr9F5LX68g/29nSLm5dstL0W9z8qux81ocNlVa
WWBrOsh5HHGbwd3gYA2BX94h9/FukLDNjiiY3ZLXDZnKnVY7rDK6SSDq5uCzdrSX
gsRQSKHpnjoUCJS6H9W3EmtlgICVD+YKPZ8+AbajVnc4/pTLcVkLTED36HgZbunX
7m59c6Dnj4ZcVMfLw1xNDe23tTZdZr3Iz2IDjLes4aS9cRPgIDRIqUbag/HZocJ3
FE7V8iS/kT2ln/Xc9ofy0ISqvxZsutgBL6eg1bAh+SlpPnrtt5EHcmfsBsMVqCEI
SJAu9p1ebmxloR9uKEWKvNu+vJz3R57ZMKKpG0w9Djqvxhfc+qCkljkNIruw8T5N
6LpE4PyOH1rZIjJ+BotONJO2KUgtQ/6EdMMRqPKjIqmJ6Bt3qvCViGpUxdUh80JN
2G3t2p0H4OWg7ja204tmnCKQGgNVo1IQhGW1ynyncmw3CSQ05m6rCAvHyDF2OZji
dbBsqE80Up9ZOpzomnniV+5UYgZOECfzezjBuMpz5gYzGfoGUXF6d8YI51zXFAaT
m9rg0tczdmveiIGFQTJS6BW1ym6Pkemocsv7tbRtK0BRnzd6i1m1OMjkSCJn0zhy
HXbTbZkDJgZPmIOlkMe4VkQlpKrAzTLkW6JMNqDD+mRQBoOg142e80s7e15tncdn
L0ybG/VY7KEY30bXvJCnXBnCu8RtpQLD3nlueQp3NZUsGN2RP6lr5XQe7V7WJNko
66E97C0mIZCI6bSK7qxLtVU63X4Dg08Ja4mSRHvM1SoJFx48N/jnHZoLGoDOFpwY
BBhsdljb5l6nqQqI0OHchtN3Ilh198V9lCuRk4o8k8jW60oHHTnUS02f3bds4paR
4/Qw2IY88NRpQJ1+H3BGLug91HSPMMlp97Y2KTNIzHSc16FDfJ7Bb9t/BMi++bWW
hRjNmdCGIsdPHhS+VHjVS9ibGI07Y5aBvuGY8R/K2FuqozRJjHS8ssg0UbMn1U4s
WYY52f2BoW7XQjK3QWQrgHYdgGy+6/XXEC5qIBLwfTkb3uvm8K99d/CRH6mPq0/9
Ozr9O5f2xhZQgsY2Df46guYyUEqoMMjW7IQiX/1MorWTG3fdOs/wO8S+gsNiQO1c
A7MVBQ2ki3gDC7AP7PnPSE0DdD9zPXr/+20AJ9iTdYNvbhSUl8laUZGWQLqPWJ0Z
WLXrRbFcIvM8W16sQ3RHkHZMsH7Kuk4DsnSnCEY8tcNWk/G3Wozuqvfn67hT43gb
xxLHTspZ3x14iprLogtHWulYVd5W7cJ8A26N/yzdJ0vd8SDfbqzuT1Ngb0aBvE5v
gJPekD97S/vyG70z24QLS5cE1fKXiZwUQ7pmnbiHsLKDAYZcDsTcnChKbL0wxDYM
T8106HKEjqoke+q4EFPPxEOYFqtYdYbPSFOLslAk9ZwIFa/nqAC348Y9498KKfcc
yjr4XxGG1XzKOk3ncJVZ81n5hbxrotgY5A7jDxewkwCm9ToMc1+JXfZyTj6opE2N
KWl0tB9HIOFM+ZR9SbKVkaUxb4TT1Nt30qFDwLkRuuGFseDTvcgUyajKkzw5oHqC
uFcEbaKJgDJ926l7ExjrYhiw1HE6ZMddsTEALXl10NINcq3t5gfloFHqCUbrOlVE
fVcXLv+fICmi8Nd33r5t92S8YgDrkxg4HtblVtUIIOYWxCbX/0KQrIR5p9VgjWje
9EUMUu7qr9Ut/vsMeEyXMMQsMqxq7Wxz0o4uRdfSyPbUUY+1zAi5ZOECnNj/q7kt
5BLKhTb5Xmyx7cfztSQBSNNOQnGx0mN6TjFrp2HQgO3e7fvjjluPbDy+Pz7ST3Ek
pEdlmKSqHbJluc0fdOJz5DQlOS8CP+Bww1J63tUFBrnsYSsLlqjm/elLDbgpaKI4
McY3/oV8zypaVZ6n7m9blgPAPeJM1+3sxiR9Izo0xAClGu2M+ixnJEYwMnZod2X6
t4bJJx6WKl0wuqcTv028o51Om0Gbx+8zQNZmsae5fDSV6/Ae2rOSIs348Qd76A/F
QTnz92j8FSVm9eYIvQsvKHjxK8WxwLTZYcCr++NknQIOJIEBArpRtH/FM9Inyfh4
NC8v+J7l/POuHHbHO8k/Cg+va30I6tlN9Ve0A47HeAk9AnAU8J1f0n+G1B9dOg3R
WymhSZmju+0HNchtjFp/1K4UWb2w12xkBlx8bkXh7qlxj3hgqh9S0Hg/aX+EiR0f
vkozVB+fSnx9Zv6ciKZ9RjW7yjxylPLzGLfilrx4yURbt7bn26B8cUYEixJ2Zb2t
dRIhQKnSoet48CX+LIfhgZVZPJ3lHhxDt1E2MAXcH07MM0gQ71aTM0ZnSjpTT0qf
Oxq6cTjgWMgq/b9jJmlXqzgPkvr93bNf1yrq/6FKOQ33ES5FdymdnwJ24QpEkigW
YqVZcCRxTIdggOirKSRnuehOwyh9GKovF3gFG+G6fooGzMEegD6lKvwrQMatfnPb
sjmSLDNVHZ5oou9Q8y99fzNlsX/ssKBEflyHaIZEQcLBiuCoUPatPazDlr3n27O5
n3l/6RktztIQJEKOT+0WQFkESlKZwXEV/H0oFvghXwmL3KJr/JkuwjwZRysP5mRE
VZo0AkpHkueRoPltn5bqmSxH82+7CItfb3zCuoU9ZdX1CUPjollXXY8Ncz7tfvYA
cDa2/QnologBJ2cp9ZtwaQgq2KC6awq8oa+jv7nanrfOLCXpzufVOcKWTlQACRkk
8m/HVhXoahUNMpfBPvKVhZHs+kRBNaDycQicvg86qbqcHTnkL+87r6F7V/VJkgGU
ZHa++6pyiL1P5onrM3rvaMV3nNy0MMMU5OFWE4BoqO5Kfrexyn6gWUAObLRP4hMW
7EJFRlHWaE7rL545dVWHMOVqrdJzs0QcCbm8BkcOwMrBxugEjyEAQR1AXwlvS02N
SBg8VetuWyupo8DI0HSRGNElS8uMsWSv7ZhcI35+IvhmuUFHz5gMAscyTz2SxKI7
6jhhbpgIENKK0XJS+K6yfEvxZNNS19C4hqPDoG/Ve8oz4GAKIoUDa/Hk1i/JhauE
exqONUKyK4xVqXh1TWyjhfuVPx7CoglKCHhB1OTVmAaki5eOqmFwv+2Lu5pXMkmk
kujUs0q2mQsSH937PN8SDZ1V/QxZMf/SHn6LkZPrrwVl7qNJ6PHSbVcpyjjx59WF
yYRxR1DG7f+7lK15JnJN3qC3JbK/9cgXmIDFrUF4aiZTGbrus+N+V0f6M0HKQ+V2
5vfmuLI18EJE2GWBDdk1W/+IuhVOnGunb23YYFu345Sr1/EWEcGywbcsaRPyqUaK
lyeEch74+wGm+uA6XlbogpA4jz4wMkYosS0nEMB6QjKL6YUYvjXi8R24z1pXBmFp
EsUWW9c3f6GgyIQ10rapxi8EJiUdQKC409i66sCez5J6mSr5Lz1Cr9ETQE+zcaFn
6cDbPPBo2hwn5i7Kd0KwUhiI6O3WJ5v6AwrfHql6o6RdKBb8tOcyWRMfXwLeXdAE
2jXMTLCeo5mYTN+YenV482fjIYgHUCtHq5tjSaXymwAGJFC7kZCCF4h3uBY4KHV5
oIlF+sivsVc0QMaynyneG3OmbyXJN4k2vvwu0H3F37nLQ/oejjblM/XMEPBQyqwx
PmNivjbxwS1kfsGGuqBwIW+Dkxk6/TFPEkMs8chorY/IwIE5kH1bG5+ioriE+ro7
u5XDBYTTunmH6OQIjg59DgqmGdlNCnBft54y/87PurLwVT5DrxVWfwBLXhOo+E75
P9v5sRND/qd+GMI5PsIxYXIe+6KoIfmHSjGY7hGTc4rK1js0Jd5Dxf1JVNPaA0gV
/NlfZJZTwMpEKhjUlApNBqWbdlZqRtsUll+PdNo5s7oEEfEpSpvtZcsDEw0RW8hk
Y2NXBcRoUK0gMqOvEzKiC4O4TTCmQu76iCp7qdpOTDwS0EXs+0MS0dQX8RjJiQKy
TpoxvjD1/Z8X1TMpBKbgmJYKghz3yIU1A7ls2Vf5+WrdrzTwpEeJkRePwq+fwYvv
atM5dmwhQJSxOlaC2D2m4pIKjK3y/TQnhUaRCh5tW2/EARQQehTVBjO/iSmKE+Ne
9vKoQzoEszhfa4moxGV4D4+hBBrOIMZFEAoj37qa7hRmz013dgF8u/l3uDDjglE/
ljXlgNscuyZeY0WYgkXQ4pvmBH+Kxjh6jsUTATbZSbRrgHaKlKg6k3cfhlihmfkg
v1ADIDvBG3gcRWgumvxCU7fSd/TfhXoXGmUzWl4BikLyxlKUlqd2NQfF4AsS3RMj
5c1jM1rL3wmXO930SqU/3GwmZOOf4qh6nuFBrB6YTEahnTERRtwjYS8+oylcjnpL
PCqznyCzEWIIU7Dr+blLZDZa4kYBmVozaEIJ80lJXgDdytS24Ve834TiJM8gooWP
gUvqEG4fQgFu0YjV1tPPwPhOU8vnqqKD7CAkZ4RfK6smN0T0AcNSN+uDMfktINxV
cWDN+PGrlva+0GnLUK5A2++dhB0ixIi2ZPDUDKe37jfxqWxk4rOb1yU46pb4qzdk
IiM13Pu4bOD9HXrSJ0KWkeZk/j1DuNbzlSGUkJ5ATaVsN/WOKvSSsz0lgnhlD1TH
QidF66WP9Dq9kP192/04sqyDTk2zqjlRrhilzMGmbEA1RJWBfd0IxMdtjPcn2dQ8
Dh/WmNry6kw8tcvvQzEBc3FrYhPAnOiWG2JIciJSZ0B+3dn3TDq/xipSRiG8Uqac
b1AVCmQEsG2Rca6WRk4hpLQ4tR0WRjT9doNnruJJA6GB8syy6p1ya1OXYxLffuOQ
GcmFjpDioB4ryH8HaZOpZG4d3+ntrTQv2bEw9+jJ8nSkmzu/M/grKilrS2qZ7Au4
atvS7ai0vYGQRGkfu/GXqF8uF1tPRDgqm/xzBd3FOzCyqk1vTKBSTQGPhgJAsphX
hVYwy/nc9dCIl5RtfLXg5HF+PN3ZsSn4AoPQTQtz/OggGcESUOrUZWQWK/ZyMmOk
EicqPYQeI9umbGRDJ2jmafCJiIlPsOMasNz464hnhfTAKAOW62kkBJFnqf4IGbh7
3XbWSXp857tnHa3tJzUcseUnqXFEJuCo5/CZXA8g0zWEEmccvrPJ12tc+lWpqV/+
v1yTY45N2oHGnnLcZOu3zvGqLQd+OPAG3u9iz26Ie6VhgnUlsuktnuH0W3xCYlva
+WkKKW0Fr8YHFa+0E+iLbGPzSoLRdHxj5O5k8o204hcHlgXkZtNmuqygHp3Rrvam
6JOwcaM/pGishY8s5saI5DDhYO8zBWaA1ftMJlIgOWEZyZ2Yz6Ejv5BlR0+/xPwg
+fzCsx5nMzBVzZyjpS5cLcLy9SIkuWIHB0MT1zgN35WslFCMHfHs3jETl3mncDT5
z1sZOQDwDpVlxCPyyuShpVK+rDtghhvVc8a/lxcs277LQccag5cbsMPr3ZwbvA5D
F4BV78NoP4tIjg3tWj5pgm2MsxH7rd2X++vniP1nesDTFqL94k0VfkodW71lh0gg
3w3TCH5wA7mUhpAkyS9XowWIm2K2yJQX3stp3GPEz7g0upVJe2tQmXS8M4CqUsTB
9tY37R3OI/3M299mTIO/wFIMLD6cPrZK4FJSR3qCmKo3KWdJNaILD0qlG7D6GR/F
xrKcRx3p48/+Qp7z4tReZa5KgES/wM8UU42roDl9LuG9TQVmqx0KdSZXyiF3xr0s
qoVXBxbCiiGKLjeTCTKh/8Kl28fG9BERGst4ogBgAncTzKjHBVRC1EtIBEkJzOPN
m/XUzQR13CrjCF7p5+sYKO8rhNmfA5L4iHjKw+TBhNjnyqN1tPudemeuyuOkaV76
HKL78CF1rFh5y5MGNOniNiTv7xbqNVLvF4ZgUvRqVu3Rnjh20RtkxfyXIXv5+h8n
ZEstPs4w1SSvSB47fjsNiFbG5q2G9mnLU7Qsudvoh1BxUsG7KWlgmuuyr6+gE4aZ
0AS2Zz2Ka1zYB1gweJU6qR296RtENx8uBNFzxdESjYIb6c4suDYs+9MC8IqkJ8yp
KRVM39LOS/rHtOG9H2qntn0eaJDa/98wxk1z4bvOs/Y/swPMC3xTLPli/5vG/f1R
zD2LFDJ3uS5WZdvw9dxYi+1z2c7YkT6IKRjJ6UkJKIETh10uqFmWvWuML9TcjwpT
uuq0QUjWhC+UhIVFcDjd1TiVWx41nLjqM2JA2ALC4xCLZxWKk+4gqBltto3uIlQk
Fj8vh5ufEQcsCnFnMnqm1mSNDzQFDr4mwzME3Gv5MQ4c/ylwogzC5ff4fiEAA/FT
Fey5Z3dsJ+KQbsXGslLbqBTM33R6L4wY7W1gKIQ8lsOUcCWy7w1FW76oU59npny/
VrdywfCqO85EEkcMB/DnRmCM+qU3xT3K2YH9UvVxmyP/ubam8MtubdLfBIzwoOyn
guPsTQKylWpSUJwG0//bm4SBCBINizcNKEa541oV9ac0suE8hEjaqyNZSiQbZ4D7
W3XE6ThS7qzP6HXuyzQ9bqHuHG7hnlfUhMEpLPq3u47c6N/2l4fVi93rfTHkm6qR
10qgg0TB2Sqo+JjZmWwU9+QCIQJ08YDNGTpfby2OkQLCuHTN26hX0d2rrGi/aspJ
XVDwQhu7PWA5+EpCUc645J/KYW8aTMnhH29xVeNYqOvwYaV8QVyWIUAuQ3hIP9No
Guj8iEyOj2+Qapki+1yusj+r7oY9ILPghykiDGtVo8gbbXk8DrP5Wfd/BlqckfGl
wyq3pGggM7Tz+Nr/VR8zXakpXLxRBjmhZP8to89UEOGhpbxZA5Owd/h+yxN0cWx0
exgY1IrlpF8m8JarWpOhUvybMeK5YEmSwCHOagZMWiFIZT1lP7fDIpvVMUf0l+mL
3VzsJka5zAT8EqznvYQphVzQcQTjbZVqEcLpvCrYPQI7XOG6EUVFC9qjt1HHtU8x
xbOPAQyvxERc00hWQPtOpeKLngHS38CymKDWYETBnACs6b6XWp6sQcaKktrTAL47
BWoTnBryWk2xjKHS5P4PtnxQF6sHZF+I3UCsuQu9BGOAArT8tMgPdsjsLefFFy3R
SlNO4A9dBufl90ey1npBfJ/0txEnDYl1pVtXur5FbGHeFpdNfBAJx/3wRNKL75ml
XE2jrN8SWejtqjStQNLMCUThrRJtxwFNW8NSpIA+/ASBu0LcWcDmEcb9pwQoogta
nsVW6GveRkxkiXo8vsukCeJhM0b8RKIaq8vKby3Ka5YqKNYPg8POEMvDBIRcY8pL
KN4CEb2RX23tjK8RmzM/aWth8s80hsqcEvjw2L5u8la2OfOGWjp9IM1R6QHhgufC
SDzlfR5E9YHn58GvzzAhqOw05FHIqhj96W3Bz8yTzZaawIK1tEjcc4We1xNY3qGv
RdOpkFnJ1IKMWp1nRoLJbgdlaB1+ypb3hEF85cuvEekkd3u2BD2DIByVgoEF18Og
zh4BJPLKTafG0iV8bUEEqo6QMhkd84+zDGOuXxKwsQqtLc5rBApLtAEuYtz38OUU
IRRVqGJEXwo0HQXP1fCcIWtVXT8okyW5NkRMUabw2C2rq3D6gypWKm/DHkLAnje9
9jyiJNMHjjXUe3xTg/x3W8Cd9anlCBUBKw8y/Yw2qm1al1HsZVtkTDvfPODugiwa
MQfAuiZur9v3AeuCiahlRIXcfbM66s6951z9OIUqe7YL4GvUV13HKY/TVDiTQYR2
WEKkUOwBspfBqoDiZpVyzNGOJ+YQx8RWqtEevkIJ1ehPiXe3rI3s2TOnhnu3ADNX
W1gluxIm9weaIvWR5tM7830F0VMBdqEMqrMOvJB+b6qMIcx2s9mCzyXi0kcDTDnI
wOtijjg09PrNv+ZiQPnZ80bZmfMQaDTjy2ICd0ysIJHy9vjUVODqRP/8jOPie5/v
GmVC4S8jJfqGcT97H8LH5+0At/z1XFfTH9dpJXgJe3gvK6qdp1o8eDiSBQH6oTyT
PcEKOkk0qmMX/oXSitOkHxJItBgK8lblCY/LTgHmEUooyl6lvockrCybZcfiME8D
HtjO3fd6l9652zWPpQrmbUHd5bj6/JNUaBIDcECnQ9m9JbIhdz2eRxuFRcNexH53
+MquE9sQY7ry5ceJNb+FmzyIk/LqcM+NqIEQe0RhB+AJXJdCMwkeKzTnjD4QnRcn
aWNHAXZ0ZzAKOhNkef+in2GoxD3zHSfpxIr4kzBEmp7JxCCWl4GT5YrH05lBseOC
gFpyBmIb+CTojGR7AhQ24Dk4MQ2niifuLZDNCGUv6BiDQdlbXvkxqKZwv23yPrEV
M3FAZO2sWiLnHla+4u0oUtX9xgHNfohbghUeKJXsgr7ae3PiW8fqkiqTNXNkN4Ph
Wa8BPoIKuxdr2kLLkW0ufBUhcO4XzZWF0Z2a/Ang9h1h8eSOGjOjWxdekc9hLkNL
/v4OQZbMJqfq6l+WMYyQniLLcwvaJIV5i4GknLJrbcLg3zadZdyPKh1U1rvQAYcy
6frN5PzxJOAIeMrzd/+YZc0lgfwidXJGy0tB5REJ4eF/auozcayVZYlYKahCtH9N
iX6hXepxzoJAr5EF2mxf8p+Vw6bG0X5jkQl5j1N2oqhF5t9JpJoKdT+iIlk4WgEJ
OUhGjqSXZNYedcNnLENmDsRbQoUgKcRJQcxcOgN/vcsoqdUGH7B9Y/MfgjVm7R4o
XQKqEJrI/tlifJ4Xc/vNnEj59wGQmZ2Oxxm4S7R2bSH+Ug+LXmSFrclkpT40RaE/
754lcsi71PEAi3SuAJ7druHxm3s/sup7llDmZAjc2Etw03SCjTrHYutN/y/D2CGQ
EM4Nrhm3DjF+biU9hzH8znwt3wZk0/uRV0leQ32XncEOGE+qF6VFkEODRk2ENbfH
IRsiWKu37q/pcDkhT1Eq2zEHLcLPmSwzLWG9R7AkB2DvIvJOfDCYZfpLSFbHbCEq
uHvOeMotuCl8cXtEJAGJ2mncxcld6GpH8fToEJIu9aCcS7/EvT9tBJJJ505K8yIg
6n69ztpBksQIwrpaMjyExv7tLHq1WHLEG/gRY73znS4gkQdtrSTV8cJbSpXl8i6a
JEsGFL+37FgUeysf9h9ZxZ531t0e7UY8/42C1Z0wbYzP2a+GbAWzzUZu4D4odai0
QJU+cz7prtz+yapWnLaP2eUzY6bOHHkjqwMPeiISxIn+br/mDb5n0S2zzGer7o0p
OjCWRJC/wb9FzmWWjedClrkO5M9G9+m/YVmVP7vi2u3Gt6T7VIwFtklGMe6vG4ow
hO/vyUApqaOThLUZa5gBoMwfvsqbDK1OeS2vN7qEEYfhgvF6r/8nGx54lOUmkdPQ
3b2vMOvdPkp0IKREBBIB+44PnC2wjJUqnZlzf8YI43zo6KpYXDuCwvfMzi9qiVyi
Umr3zTehzSnusDB0bgIr1gGdo3QPPun2BPBSOadsSGQmnA17yyvQRZR0xFIaEa+3
2l9UfJXDKxYiuO+4pFIryo0CoW2LWQa5hsbzKcLrW/k0XpeX1sFGXHO16w1d7GBm
9EAQcDpX45TSFh+y2H8gax5zja9K1RWr4mxbx7XXceCSVmZXtPvEQiM6qIhciI+v
bGTHGcNq38ecD4CjS0CBBDPSs7mZdrTJrs2rdriwjbQF7VaM0GftGDfkotfITyRF
K1hIXp/7REJACxNRUrzoCdcwU50SEzpNtX1cWxJkBjBzpSav92qsOebN9rNUj2hG
WBokMqhl4gEginkJ+AQaRYjEX6dcC35Rq9dYYN013zc783d/VezNCTNsmTBOzgu9
MUFI0fNdxuce7srIfzNjcS4b9ywxZZQXVRD/QwJwbwvmsSbL2bn+NFpmf1ISAEYp
hLnSteMDPYRm5tVDq8MFnNzqvZLj7LdjRJJNjCh9j+Gr1hDJ5yf+njUkYf6VAhuP
HQzZRSfrG5Ai8Pxq1wCTfyeLTcHvC1KDA3qeXNYs1nThtpQ16O7TIQIBwnVQU6cX
8OvIkTuk5daiki15V3qU1Jut/kL4geg5yL4usChK7S5Ho3zXasOseCb7ewM3fid1
tozRQ3eaEK6qatiJ1poJUFYv6o3PwBRWDpXwZ3HmyJvpg2sAC8BdBkyfHXkr578q
hROeZkZweAoqpRyW5BdON+ZxL32WebqfYJcF2zUtYN0MLv5JsDJvmp6wxEOggT+I
MUNBA7KT9FNq7OjjApqdmv35lWvvBNkxYHppjUGNnrmZ6le2lbuOUBzxq3fjVb1g
dwNj5WkkaW1t5PIdaB9DxBVSlcv7vdU8ZmJ51z3FRTZL56Mv7iEF/afozNm9Ogt2
54rYpsjDJZZJ2eRjkyDl9sQdTjL/LHtb8xnvvw1Fbh3zi04ZXSn7w57PJ/EFtGnF
2ZXAlAuxA5y2xghx79bJ2JGNXv4K6I6Q+312j19u/+ljXuTfOjND4HU2WXtzFHGf
GdMrw0ry2//BOjmgz3GqLCCKqct+LB2Rxxne4Y+LmK38Mv73eCgTz8f0DK0wWr28
8GPcJKXeEpkjWadrmUNhclk1gruXIpFX4futduUzvZC0QIejtfLWwf1YMOvjJbnW
uULWzd+vf3fmiy3yPEisg/G5jxwUyFdbm9OChHRey/NP+6imMXu9a1XIuFjKNNtP
ok1kfjAaVKtZQ8ZwdFZTEG/pYzKxqzKpoFoP1Sr1JuLx1xiz8jO3JAsiTyADTnlX
jFj8ruvPZvzKns5pBwiSybxE/vwLXCrYqPHFLgjBrNWVB7vm84JURzVb7yzDePsH
oebEDRb93zs+dQQ9mvPTINs4F5tbOUr9ljQdmlNJ/JF6lM3zrmlvlgQ8YN95r6E3
tIiKDGp1Sl7NpwVyqi5HkhBp0fXmi8l+R9LTJuWTRIeCaoghJcI6iaXxdJ2pJrkm
snF3Pa16cK1zB0XA91BGlFpC2zJmX2x2JtubminVwVKAzpuh+MjfrqZDyh3ncJX1
XkwcfpX7QGtSBxxj5pVLIAdXfHsfeBupmw2AoSBVy5OZljsXPVnLK0o4JacEBPLS
xFtKSml/VfFtN+LaUIXd9gSH+sMAC33yCS/Liyes5ox4kSNgJ7trsv8l1zKtJlSp
cElNqo+IIoqhRKBVUQnnNLrpyicCdVUjgQQjkS+nju37fdZTfBWA0lfKc5+2DmLo
CcxYJfCxEBjweACWb9eNw0JFfvn9XIDqAY/EzvcnWtIdE6HA8cQ61Kly6pQi+kYR
teJcpvNeXRJOihW3M/TOH7QdZHxYVuODvG1ykYBlqo50vriUOrD853RfOMQ5mzaH
9OLhtcMImDiOxyPQ1Pr8WidaVF5/eFMA7hFZThXIguJKlmP33JIp5YObwu4W6uuh
V05iYob9Eowsfl/v4bR8Iq8HKvPAsgQY4x+tKnGDquzlNSlWcOOlfdYA76uJXmee
EuRT851KkMIxWNAYeHpSNs+g6+Ttg6tj3MzJT7HYfNW8n98eW+K5RST1fH+PlYJV
NDJxxe6kYRbY2rZmXMpkQK/YklI04Ag6xVOveMAb3Pif8K1NPXtmipoWlydvEe8+
NeGRNuqT782DyhQv9/qrEI3lBVvX37Bwh/fj8J5x4DkHIWW063ItNJdx9caaKx8Y
Q6h/whpo+yHJzS08AxMdSwlvzYcZnHeXlotTtd0R91+gG/Epy+MPdpvHmQK1BbOt
w8T8/XENCX5SH20lXOfy5znTf1QxaU7zLaKhnEIXZc98C5k7fKf4jZqA2oW7AWZt
Tnx+Ym+03XU3Dad+sFElu4k+20cjwT+U5u36OoEt7qFpGy2wzFwiFAGVQmE1oM5W
YMXmL8O5i3Ax9BSzXFYZ24/j2XP+TWCnAd98oDGKmdMvEEnYcrtFAtXWPZc7/98C
TAUXttXeb3tUijgOC/597iGbylOLYuhu7BZF+BzMrY2vd8mf7OWm2l5z0M337QZ6
1ZIdlQps3Gzp08pLamgNzj6XMsAun4UcFubNx073Q7WHrBYn2y5aYxth0Umc9D8x
CQLahKQ7Hhi2g2tdBSxQFychIJG4sD+FurYlG1ksHSTOjKwHFfHXpRuFCDe0XgAY
PaQKAdQGibG0dn7WinUPV0/OABjm+gHDfCY5fmD0viCJsq0n84PXE70u7SGFayQc
ckfZ3PMGdn5meYQkJ7YFx0F34RA18cg5ACSxsQfs5hNlx3JRUd6jkLhrbBidHd3I
ob2yk7h9Du1INUbXxst4JR3t3vh3ecjGuPDRvZt+TNwxlO+So8w3Yi2GqyB1SyIE
oPlFJYLp3csrqLK8r+/UdXm/E9j4sareIBolmoP3wIOTukgGpSeNG9JyNPeV7Swe
Ogm53EWZkqwe4viWCQT68rsSIU6bs+DmozJ8ZBt7TVuAuL6RbGD25G0Vjs5cD1mF
P663EC8KUYqgFpoHBCm0Fvg7UtiXSTCSWnCRvpwVjkpu9BFTbQV3NWXYqH+fsNNT
aRwM5Xc3fQ7Buztb4s0gvLoU8iFMSL5gbLNDRvGe1lN43yUKnErbYdnKbJhrkVM7
jBE/eWUd8/b5+hKMBuyiZIkr1CO0mWsgBwatBsiRTjhOM42Yda8H8ov42Em4p7tQ
/XTTBFDAg5tAglDs9f52v8v4QATz2/get8ouljEOc7b00tAlKjtBbaTkx5UjB9Ck
TsNdt6aqlAruQ90CEH0xd+/rmqcdkx3pSVgdq5xB88OUD/yYo1fSWrJlsYuWZlPM
BU0oNY+EqLD9qPL+uhC298Zt78KkREzRoWj1BBSVaqBbNfXYMG+xnJpRVDAM/gtq
fKSznV55KKRJ3uqKRuj8r84+wqZF3WuvrnrIn0xlfWxju2NgwR/kEiZMsl1T5SQ4
sHkIoh5AbelwWQLmUJR+H3B5eTIYTrI3rVQqBKArRPIxokdt9eGSSvBr5juD1Ilb
Qr5j29E682pqsOGTDKbV5wdwSrlm+MGMGy+jSqFE5jDktKTuSwt5FBXEDTlJLGqg
jv1UtbaGIYLbx6cw0VxyygL8W2x++1CfGMDY7VPfKcldKTuIvqyksfeQ9Nf8k1iq
Jt6hPzYOZj2xpDzDBaA573+AeWZEivsuyJIxbjTQrmeqL6L7RmrmcvWsSW5EHnhk
gkOSXKQztXNLd3qd7SVsvUGXyzpn0l1XfO2oo9qY/HtRnsYohK1eVBUBM2b8Dt3G
0EiJwYMeyVbls3UdBD5w6WUT3/5d6Sn5bkHrmvwcjzMGbwJnsTb0TN8c63d09r6e
I76Yf2ypLsN0YE1s/0rIX3hYp/BVZbGCmXvlHV/H2VG/ZWp0Kap5ezv+n0COWkKV
ZrxKgfcYWcSHfKhpvDmjf5duYaSG4YHCUNKHw68J4v2VNeeDof9+ZZ7I2gZK7UKb
He4k2hG9WjCvpmf6Ypv952L9PnkdEElBXbHtxoQzxCsQbCJ+Wh3nESEYIx9/tcuf
Uui2AwqT02k97b4FcF+FWPkYPR4ein61xlpsMr626MidQwk37IGevmsOxrGGTfX/
VFohVHWvlrIMv3JhyQzEUD9d8AXNY1mzND0NHIGjQle70iL3iDXc3G1chHqlCFN9
GzM2ZZlfbUAH7kJL2tgKVtvXqSHAWBUbB0DAJRB1gEC85ta6rBxP7MiJ5xrG4o0J
VgNftu4dIQDHZ4RWDhY0cucKo52P2azaJmTHApmJucns4mALlWhHVLF91kXFZcTn
EqFzRh9/8LfPja5Mo4KZotilGhoFQk1kbfyknePN/Blv3acZHuj9MDMWb09OFIoN
asFpaKWe9hMv2qO3IYBHlzAPGpJapf16eK26eCXVv9WXc9B0uZLO3OvoRPkrJBN9
KmTFptrWhy8as8U+7Zzx4MSwhf3OxwemX83D7vUPBv+lZN+FAZ+CePGAJcRfXM3t
AUurNmBP47mP4peXeKKdx77q7Gn5CT5W74G0Jahg5Oe5A5h9XEqyMrs8q1N5jQbR
bcfOP7bmYowcOfA3I9dyVwPqC8Rw8ZfVugWnYnf74HpfO3JCHOAj8kR4ywiD9n7o
o+R5wPddX3jYE7nfwEPA+AxNdY7gUWUX5g3Rn0VizfWgW/UKJKEW/LglFEcjC2gt
TS56xu29z6RJkusEZONRB1Ro7FAEzz1+2V/2Kn8ZX0kKRS0/DUF1FbSf+buQuaTX
2Ie2hfKtUcHNknQhiUgwieyJee192PznvNmeRtMRvvt1WR+aLFRVriTr1adbzcfs
cnMGDjn77n2v2ihmuQ6zBOAW4WpB1eQPkO41In03y3A8IKuwh3APR1+1ZqTDY73o
8nSenugrS05yYIq6IaV2P2wrM07QcDbC7EbAz4snKvKvluxlB2s7RtoYmKveNrNO
k4sN28/XYQNfaJ/o2JXohoKXeRd9NdVDKNwTrwU0JaOOkzIqxglPvLIvc4JZJY1/
U+ZZ3Nkdu1YXoo5Q4XwihzDUp+/1rbxotbM9qgeNHK6ajU6cax4yrl2gLglCvS5h
5FWGF+owRat3pcXCEMT14tIpOn4qudPQBIAaFMikQCI8n3wNTNCqpWWpZM24iJLB
/dDRKIiIF2rdZonm4Xg7bVC4a96VOPmdzoEGaTHw0o1O31KsVAIxqBZcxvqJjuI2
9NhBmwrVI/R+UcmAUP/VZ3MZV4qJ0l0BARLEZU40KctveEL/3uWw29hNiU8TNxyN
s0duefQTTuiFMgwIL+X+LEPUVT+wKWr4N0+acD2FvcS4Dq5VAH/knVIYjSHZm2Xn
q5KgXXfWKpNoq60cA77x3RLsWRIY5cf+JgMVPsi6paS7DNhtq8LgLWTB1iBCngJu
y5IrOL4lDQMLygzYYsFf5TWtkBbBGbAmpDOgHopMuodSrnTzz9mTLFbTLbV59rRu
dW1RMxRxdHq5XK3gGBz506C4ZgZthfr2HANGSvV1wOTSfqi+/5GTvpqDdsH9hurg
5e0KfdNpOJLVlcneSVKDMPFiuJGv7cFkZGiNcxxtN2zEEfCfe/y/3o29+u5dG0DX
HfVsH+mAbHg9mTV+o/80Hoq6CFua1JFN7fpk6Rn/zJ1SnHRf/w1H7RYPvfXcQIHr
GklYVyEUENmJO/FwKCOnO9MHtaW6DhDmvAPS2zVrUZYTZIUBvxfL/FKG9lDx8Ggp
GoPlUly5iTSU5GsTiKfnUJlrxvrdx6bs+OA4eaQMi0hOZdoCobS4QaQYNB12T9jS
5YgfbyUvJaPHGsHqNIhFNuC3tv02Gg2mXleJ1lNBIGEtmW+6DATa7B5JXLwCmSkf
f1FtVtps7uf+yO5gewmuk2qwn0z2EnweXY8lC0HtbPrhclRpz393jVAtYszgXuTm
xlXCWZ+1oHwwfW93m2ADKxl68TlLFgFm/gNsa2MEVOUPyXsxlJ5MtACZpfE3SNMv
SZImactNh9cySYUJDjP1uXN6iagOPr3QvQ5XsDwUjM3Nyzf6zi1WcosiPQk0nrU8
jo653vtXorjAuBNyUuBft5pNYFHDM8aafrdpowInaDkLjxxeaMoWdFjnCmRJX2Mu
atpxqRW2oz8XpkIsDv2/X26Xm1d0U5OrQjcTSvCE5cTV6udX89VzoA4mqZv5x0+b
motnRh0FLoo4bGn8iPd6zPYwDUdMfh1RVDb9VkyMjKr7DW6tDK5jD59wOedX1lsX
QVTdgS4lfAU8TWlEDKYaweFma5tOaB7dGNd9hdt1OEYltGY6Tgfqa5xovFxXBFZ9
Jhv4O7CG5qSxsnuvv5DWJi+x1iBbkTo0C55B7jFyOA0C/BXd9ovV/rGOaQ3GlaFI
XJBh/XaCvfsPaXu0dwefoKF8T6st5kvxRnZBt++pZKPnPXgzJuj9R7qV9ez6fpcF
PhzQGJ5PqQeC3AMXKfjMXFEoa642oZRvjPec3G6o0gjzgri+ORMdwAc3bpd/rfxs
hPI7uD0Bk8tlU4ySlXDc7RC+NUCR8Lr5t+0F0n+f6IOAYmFvdQs6CyW1IfXYWZM0
B4j+2vXYzKO+M6QkbzWRfiu9EaLQ400nPnntwmdCvGluzbJvm8CtQmJ7ZFeKgtga
6/dn8rL9Njf3KK0mO49TujgY3KJZyIlzYAAQutZjS2P91yHWUkl4eSbsGG6ztH5Z
+Ii2J8O+N/geWPOt52aYG5484JHsF5pouEy7VUqo9qbBZF+2jw1Toel+KMBgeubD
UZVzg8k2XxjVsvUr+0sZBVoQ5uUv0fLDG23ZZU83oruQ//D0eCmsyFFam4XYYpvm
udAJbjmPxgASiE4DyDvxFicc0L5OMS0XbFmMwBp0jtPjhhu+m0aEc07lbHxUf5zo
ec0ptujijDrVJPYLwhAHRKDDcbHOp2s5vuusK11sg4rv1UExCx5P8HguWxFHRqC0
zcO3WGboyDiofdcOG8/rlarotovmWZ1yuBwsbAXQE0gp3VU8vyWLH2PlzgaE57b3
8Z0MGztxK5t2ezIsz4nH3P7HD3GrI3qXQ3IROTBbfGNYXHFmBgbmseFYjMfhxflM
U7g7gtH1gNzCcUiSndl2K+AmBvOO+AZLNjOw2t7IHfx4X/80c2U0UTLgATitdfz4
jZg2lYQOimhQ3rh2QyRnT487Mqpuzm2EuN2evuw3/9zKUQ9mcjgaWaP+u8ChSRvQ
YRqQN8cuvhCAK/TO0sazpqyqO1490CteMXZQIZdFWjEIQqI+yTHzM+iTFNghCmyR
peC2bDdhME8ameiFqok5+MNIbnplYUX+1jRKSC0JnoHrFHOl709Q3dsJUlWroogk
RXbGV1x4uJ4Zfh+ctXV9SYF2q9fSmLcv8ukH8OuF+VPLWufMZtgor0vQ7rlwp2+4
SMqf5hT92kPg8/ogizULnwz4LAqGb8d3mXiBWD6XRXAD/KF73yx9VxV5dsHzoBKN
okbhwoTCsuH1otnhyPdHNWicUMBLudyxYpcPOsyi8hhr8rZndi/zX4ZOUIagZTQT
I4KzWo0sGrM7xr2mcM/bMAuwgtMQ8IYoNmzmJX41DWAx67QqKdr0ouYa47R/17wn
APzNu6quZwlxLhoXBUtqPmf4QBg9SR8LdYqgFg9gHVT9lDHbGcDYIwnkx/2ejbot
8pmEyUzH/LmQSgEST5bb2zMbGiVrxCaJaKACQD5dMzbzvj2uevh3lkNr14/DYEGO
elxW8jqCtbxbnZXLzENvOFU92/15uOHJYMmJX8VIwFp4QTXoWWAARnFlMLjZY13o
yAua4Vr9gJ5HLw9PREbBTCP9d3KergnqKkxrEljU48kBbbT22PNbf5jcbj1CGj0y
O8tkvdg+fy+oDKxZedDjkXvlPDbV86WNjfjUyCLHIihrFIMa0QrA/9geYDZE21Bm
ni8S9VzjcTsp/B3+PEtgjPgp06FMQith/PvMkei+RuM2pG606Mc1zyOKTnNAAbvt
JNY7Tm3vyECelEZo6lLMGXx21131XcJqxBoBje+HksRtEzZkC0spqR5n95Mntpro
Uh3cIVTXzN0Qyh09YnafjLniOAVhDDOso6c29moMXRvnDe/+XOrFFqFWa0EOc3LV
ttZYWKoOBYvuxBizZ6oIifPlUHDWUZoyPU0ynOTqdRpp2QflWfWIesBFkwo2e03/
R9cNootmaohinW2mRcJ9ybk2AxgSoldWxI1vCvFC2aIP4i+0IotmfJP1Af+eFJ1N
PiGdtNAHF9m2RBZHMBZyeuHqsnbrP8xoAODybIXehjRMdGTwZjVAX7QdwAVLCEb6
nO8Ojz12TTSvYcxdhY786JcCU9UwGe5XwqxnoAayF38xDSzxtjK8bGo6jtJxCUGd
O8vOpFNqKypskOlQrNwaV2Dknp/8hBwM6n4PmdplHq6keTozJk+XkT5otekUxv6k
eeOUB0nqXdv9RDM59Fa/A1fz3l7ATVaeDw5oLuUEnn0fulz6d7ujlQ05RwQ8aJN7
sryzAVUoBlIb36osNJ9MaVhWhFWr03LXJGbAg8sev8oDqDTsDgOB4V/v8NPI3qOj
X7X+hIAGBlJblSXgxb2RbWBkybvkby4Ivsx0g5q1+l+MyCPSdPLia2lruILSeAFX
n4NeB900KGEeMnSRhkAp0uxp/QqIRkQC28AkiP8eijg65eGsYoVJH2vyGOesvmgh
Xzvkfu+yMn2+Svl+dGeaNcHh6q28sAXw/zZsLV69oM3599hWgJHjHowOS+/aRsIx
Omn4XmYOx04tOOVzLCeqi9IKwMGs8ZnspkT7saG9tAfsyviQRyzyTek6lxL/3l0y
5zO7VXLe3cW53hG1jF4/vChTFMhD2Z/l+5jPOmd29DPqUpLV950i3musSIjMPZKc
2PQBTpXIQPP5s+l62j1VmnQjvVuOjpGcv0kWEm4XgWepKjIy2c0UrzDE9Pvwh8ST
yhUcj+ADOzik0J+x2W1trvlchfEmYkBPqNeEIZYCuRGLy4QlX5Ska6mYrHDwo665
MG2hPd3tp5Jqyw0bKrYa6ksD+PsMPXWMryXxLSns5S1wnsA7LI3JCHnv3J3DlWK1
pXqDwyC2jQBRU4xlHDOS7rTmFyZqS316RhEv/T5Zj7WTLvZBH43LgbmWJf0U07ba
AiXkihqus+dY3ZB6vPhES0scw++AFb4Doh9sVjOSeX7OnyDfPwiTUzR7kL6SFv8z
/4qJ+vNt1h4QKbj5PYbwViqzAgU6iE9Y0+TuAAgg1v6pQUY/XqkUUEKGEh6oApqa
l4NwOq5tonSozInSKW8/vSr+Mi63YpivTmUE0y8xttQROyrroIBH1e4/C2dWQ8nI
SguOCEflRGE7WGG3p3TXSnTgCSIM20CSxuSqrVY9R6Nc+DUm1ioPNb+s09r6n1zX
Ma7qIg/leCawIAzHnP6VNiL5hgkD0bh4BQupmByXMzts9L/KEzmDNCtR015MY9lO
XapRC6PuYcxg9o/epggB8RTxGZTwdZRtxXRwkrqsE7X9A6R9/GgDzWn81SlmTGNL
rkh15Ce1tD6FFrwDzslYMtvzBY3Fw/0yB6UxF9UkGiikRWhUapsMfS1Cv1uFqnVK
aL963POYLcld0+i6u9DhVcKoNQzAdhW54N8Bw5c5XUL4548XU41loZMig9ULyeGw
tq3aemCh+e40QxwmoZ5DooyO72pX/UOhucm2Zxli9QJifJGvoW42BW/K0EE9BDeT
3CgIEoLeUApxS4b1Af5ql2+GMDdNs1ixTDVgHDfqLOdeGOgtLMUJBibp+S3y030/
kq3N60t9k2WqlglOoRzWVRA6QI8xqUnJVg+QvFdRMlBi9FYeosRyoeYg/ZPtEAtS
7Z7zeel0XUoYQ1pSkAmnM0kZznmkrWVsVZb4iGtikfGnhxdHRPQnLqXcywhtxqnm
n8Lyfa/TkdBbf1i0AYihlH+qoDCTHuhQ8X+tBdqGJaK0wgnc+Q/MPz2jYTcdp5ph
i8+JD8UaCrpITxsz4cyfNdVpFdSSyhL2A4gQLET2749grFndCW7QsvgDQ71wEtSd
+VbWfqdvucSDctgvxEyE+fIUXXXvPOczbaDZvKvGrSY7AFO4djBbbAjP9uzey1Ny
PxvLjbSQSOi+Gi4gZRy+L4rTjfPJhsdwog6GdVKWcww6fUZnceYPXdleW86mkn89
U5hfH3k76SoQ3QfG2wiEX2wg3QI2mjcxywHPaFD8ad6sg3F78GMFVOmm1Ek8iLI0
i2OvzOzrxHOMUSIKd1BTPLXs//gDHPJxZDMHLFDRvnfO/N4TrloJzo4UAAgaohvo
kQkjVEpT5NqbUAUWtxdpGSwljeYexhciE5R8XsrLKujbiETn5DOmmT1PV9CqSsRe
wYEgKl8OrZMF6eQ4uCO3jZTpq6dDfA5cWzfYx75Cm3zcyG12+YorOdkraFAEAQJ8
gzNvgUsbjLqRIvHttlU9HKztKawG5wPSmzfwHTdKYRs6Tfk/FKdkrXkiD9zhYaEW
y8Mgs36nNiCInbPsewrmFJUbdMfkZz/m3Pg1HFbEEBtgmEYGXpv8xIWBsTbqUOaM
rFNBTyfNsshwnlZE6MLbB4zTrenJOULT7u3wTUTH902foXEm0SlJgis2rlGJI9aV
nean+/+B3Qumbw9r97b1kcvvc9QPSiWCFnuWymBo4iD0C7FomYB1dlrboRahGMDX
GbTp36xW0DNzdYmk4F5kv0efnscetWQCcN+var3F6o/bcdxDwYD9BY/Jsbhr44Tg
4JzZfP/FgA42f8cvkhPxhEMU2GVcZlyXe7dCLurr47ubJUdRJSelC08bAZoZUiBh
TBncc6uASon3aJYVRUiFAYNF9rYA+aq2i5iTt3uqXc5/WkIkxBcYWc/BAsGZ5F9U
0ho71adFur4eGkj/+MOeyUGCGK6f4TvJjaEHzIWMltZJSMwslZ9Zked2o7RZPyEr
YkGu7419qpDGvaFR6tDuqeyLDSb0q1vgBQG/zNQuHR+T6rGAymZy1wxop+/GDDvj
DbPCQxuy5zfrlC0xVmdxgU6BudksBTE5YsngUfM8qX9rFtlKKQ8r+LsNSU7H4hHM
rh25p3CGW4m/aWWaBzhqyyx2ihu5T3AaX6CfE1h3kkgGhpb4YZwKg5JvSJ+CSF2B
2x7sTA5tg668JyD9TtoqrBVfqWrXRGVejAstImfRoP/uAeftW+s8aHja43+W3V3U
DQwKr2yBgul1sGbIOn3PtuoF1Y24nArKJBTN+SY8XDgmLo7yc+REDklo0VhoLZaV
e2KdXYJSkHwOtSQGWc3NCY6/SaDhs4nGUvsdhzwk7jR8sh2lQc1KGzhxQXZPpUY4
U3yRReoVDE+YPJDvOljKWux5qDO8RvNDtu1oIi3bIopTXDXIDf05unpnbjJkGdNr
nRy0+kfwvGW6o9gAy7bEn4grXg0MuRqtTM3d4cElFva8Kln3Gli7cJ5RWJaQBOh/
PbdND0sIsFY4eXS7w8V9ijTREmCRn5K6rzBIGE/lfqWY1KZI1MVF5aoCQKYyoVWf
e1WHD9+A/L0Jc9ebtj7igAIb21qJMHa9sCop72F4SBL+fCzXdAVLk/Guhe6TCSSF
dNlXVYoATQjFUC1SspQmHFpV/eIRgpwEaRiGQOmtOYTTpaeiFKM+IN91k0ZkwOXP
kXn2EnahjDX0opYUs7ApobmQQlUY6Xgs32G8QFCjjEDN+2Fti5AY8uQnIuEtGzY1
pdCahgtrmnbSLWUIVwz5Y/7CssruY7hN4K4DpQ6JD3Vljaq4RePLpPWaliHtlFF+
0dkbJ0t30lZ+a0W8y/RxkJp4OUksNgVOMeZ4aKmyc0MtLoLtsjsyZN95AsCUmiD/
VyILKcnZdod+nUIqX9HqQCTAQajFUu1W/01hEzBx9wMb9lm8rvD9EqHX5BwEn+NI
sHokjOfdU16R80mNAMLRbIUfGmHajm+h50+89ih1Y2tHWByN836+sjog1rRCnvg7
FPlNVMoqsOzaG+c8VS+/xva/wV7yXUfNWbr6GQpVFvMLlO18neeAIkCkxXq+5pS7
R3QS2n9mDXQ7k4GejrR8dRR2TB4fUlA9ur0zUVl9zEvdW91dVq+sDfRsMO9oD/Mq
FSmKAvGwJossagR6Z5iV5ICjugIzyClRHbnUDMLp3MbjYhenoS13UI0oHQnWH4fp
/2hCPkVp4Pl52NPe9GmXLt0/cShBVVLY9t+SrWs/z+vqjSluwj1CsXLhivprHGWB
cFj0kk47+6NrbYjKC8YwfjKaxaJEqT4Ev5wk6BC/W17XkPHlANul9Kn7u5RVh0Q8
yHbRpckMu/vRRarzUzyc/007wpNR1ylAVz3npGJcU0ACl19xEp7CDYVBg5Ax/OTT
nJh8R6oOCa+dbwcpoef5MWbzQtraZ5it8AnT2o2oy0v7Pf3j+QWR48l240ZAXKfk
rADIBVTpMSSE3Zf3VFNbjr/Cmr5w71LE3X+JDmMQmzqmMuMc06i7bF3VD2hc+o5z
B4n6kmbqWCrWv0MzSsTPwLozSl4AxcpQwSHwglqjDSWEDvoIAYa5iZqbBRy3gtJS
F1oTvJCjvuPHagTpXEyykasS504yBjJPLoBHCPgOPd7nYPx/wYpcRNoiRoAQAkXo
2LP3m24iNF1qUAxEUkb6LmRHH9P54YJE7Z6cHCmDDKmb1vz/aDqfMbgy4FDOZFbP
jHUYCd7JZyAXweKZ1t4HVRgQHI1IyaG6w9Nti/PzDIXu9A619G5prDxjwqeApGlp
0QS+dkVJ7cuCmQQ/xLM8olXF59Q1bfXJgqa8VYkyM5Qv148s74sw2PvJAaIn2V1I
8aVfnebImVQp2aCQ1IWLOopENdfRsp2HS2nJ6xEbicQuCLyF+1v8THiBAbDp0rI/
IpbngfsxYjQwruWsA13sTS7GL73dTqRyi79FdE/IU6TZxpUe7vHk6OXZ9Wa1UuAo
elWkZXl/EN3zEsMlniNKhloyNhmqG0VRNvvsVJeChf5dUM6clHpWa82QKt25hTqt
LV72XUd+G5rXU/oazLIEwDMb5lJRcDeOHkCgND8Q1Ndqnl2wu5UvpXTrlRDsWbs7
0g2CqrsxynhmPC7C58k0BJeCftOWBHxr5+lclbDSRWtKoV41+31/7SUZWDzZg+Tl
eo0aB3Gqo3Hy0m4357ur5NZ1fxtRd40o0+CBuNDGYbpuopgCeFoPYeb3cOEo46SC
OrbEsvSh+8H/Xfg1mHKOUpWUQL2O7xCSqbQi/2m/KAH9OyzG3nkQZ5sS/mPaXfyu
608cUt/JmHNA8H1CmihBwbIzV4H8KIW9xUwSfJv9Y4j7pSsfxfpDfcq9Lw2s46WH
29mSKciiIWJnnJPVdm33Ji+GIGlSE5FHwgGFtWTrdKcGJgiOK/7c6GNiLYLOim20
2QZimtCEQfj2+VqG4dRzMxuR85IWDoHRvpUsoQ4zUBvQImo5IW9tcr7dV0LrO8jH
MAlBYXL+JTdvs6DfDNmxJMGITKtCN/57LhhyDX1M2hZQyFm1H90ubZYdb9orDCOR
7hQsnoxvqW6h22qnmU74g+zpmAh+Snr50XUxanxvsP4LGEasQr12MK671DrtCiE+
Xv3Zkqk8L0zTwKXHSwks3ZT3fLsi13aSkQOtocLWHgv1TJrEVJwdgw/7y1EfJSEu
WQZEgS+B3+Xozg38gTBkmQI7Y9jew0HEDD4iRx+ehFPmIXvBgRW51uoRhFRctuhD
UOCviJmbWVDQAZH7g9pmhekQkloCzZdd6cZg817hz461ztKv6vwaIAGjc3hnWgQZ
Ab+VCwdGBSSwd/r7ZS9w7aBpWue5767jj8rCnWrMgL9fGs6/DORTyr6WMfjbalsG
Cg9g0kzCy22GW75agu7GKaBa/IfanvPUbXIc2ljhdLklRwvw/Xc2zs8e/fH0N9iX
gU/y4c1hXnDzQRjKL9w7dh05d4IvY+VUtZl5xUjWWWJollNACObexRujfEweI++X
RniCCWB5bPnnQ7njsikzi1+fVRbOPoS8rfcd3tpMYICoXr325dmNKrdosebSZw0K
76/N+1h/e0Qx2if/lSklVicZbouNWktwEQTv7pCmb3YOW9+4c6hEynQU1p/n442c
OSY21IvNIKHrunyxD22wWfAcBMuNgRv3L+gYaPGoRicnCpMKpcW1YncYdvG5Tc5O
acWiF3lNiwELmQ2o++fg8HQesc+5yXk7oBNQDbIFkjnEjAvPSb7/hn/ZN9eEDyHt
V5kq3koVOAV2TCoVj7gIdfdQB1dG3GPycPjevEna+8KFstFqCl94GWyyYfyGAnFN
caNmLPF0XByBnMHwy/rVqMdm9Pz6bYVmjRoazwT2ejMsBpgCDVcTOk/RR7hyqExI
X1NqQEKvKmI1rGAJaxZr1gPleUtfMHEY6AvgLiXfzBXNBOVu+rr1bM5HRTs/5Myl
B2rQ8rkxQ/iHSxQAnqtY+/zYwpOhKvos+7B0+ZDEMokl3vOxE2TQnZl2buDMQF8d
+SFy1O/3hb17OPYorUodb2pgQ+JkiaHOPqSNDCAttvmE2L/FZhXQwePIVv9A23Lw
1RmI20ZALMRfmKjyjWwOI0ikhKlkDFUZIaNVvj078040lOxLU5hRliB84wFLtlzf
PeS7lKpgLf87ehOrWviynplslWuFMViVcbvIKUAYKWHXDx902Pl4cFHIQlwgwy44
YuB2GiQF4mPIXjVnhGBMDpfmunj+eHlOM6QxHbcv5wFJA2rsgbZg4a9ldgmwbPlG
nBEY6R6HN3AHty4Z9DVS3/dvI0td9k6iuH3HWckLSX3G97/EaF6VCztn1A3Bpgke
MrfnNkGQju+t6c7Qf9/RnsMNWXEwPzLdj4V7H0T80EkxCK0ZCM2csed4L1Vc+C2x
qx2N55env02GxzK2FjFqh3+UX6bwCLvIY8mJpe4Wwg1jdjDujikJV3oCohO51AEM
hrMAtNrf6rkM9pz6lT93iT1VpzjbyxyUIurKGP+kFcdVriOqAYu33qzmoGk3+G4u
81NOpmQ9GhwSB/4fBLSOqN5A/j94pbuuWpWMroGRQkzaHl7UyKz5TqUxnmw0E68B
qtCaamb8+BOgJmSUs6CCPch2a/C0SnHIgnL9gIz/qsSXn/c4oSBovVYLKXsjGsEi
bEVfmi1cHU8ULhrxH1I4wh335E4c/Ujcetl5ttrLJJfqlTQcGT5do2SL7juCKv3Y
1KoCoUltQYLBi/Z/Pe+eTjIOon/Hq11xQls51oDigwO08dmFRgLndODW3Rajo64E
8QWQLq0JLm8gE1S/Iufgxm10+tw+E3mZpK9TlTqlASw2O78M1UeEAwlY0a7SLSvC
lNGQmWzbPVfF5nWZuOTCFjeTzCVSdtDF0EPQHUDL7iQowye8vvv/pfET3Iw1vBbN
JJDJUV4sj8ZVMZZn64P9Ja6EwDxEeoIXczXx16tk6loSBkQstBqX/39dhL4AQdQ6
3UzLm96dot363L+zwxRDaQaBZ48CikPO/MbZDwite5rp2HKbRunkJNemLAF0Jqb2
YCB/2cANXP7llf9iZmnmDU6hQSHoRCL6QMZvC+RhPSjFy9AP7F474nxKFdfFEIyn
3JDHOcWBskIdtczNYrcG1o7DWHcFsD9uT/mMbATjW4+Dg9vp/VoNhd4PAp/N4udT
8lAF+eanUX1TCymQzvmC9Up/JHcAmX6c5hmHG/SmP683IGJNb4HaIvTp8/xu9pNh
wJfqtX1tPigZbVf2x6eAQ85v+ODINnO3XqB7vK+X80JOYzaK8wj2RfO4kcoX0PUJ
wDvl9mAAmbEbN97ppj16GSMaD4CV3m+xfda4q15NSxW9ji0/oPfDIWl/M/V22coO
AwCKFAEoG+oz1/HCGxCrDjmbDTbzDWnUMwwJGQ6GwBH7rAy8eLu2Tm7/5r9ecFmz
BCyvBF7ug2+xVHcRhTcunAkNz7HlO5lyu66BJLbgqZTf0xWekK4VkLMnIhc2+RjD
4s04nTvzC2W3/3HkxpwHbx5HJn9ARFCZgCej2w4aAZvtbFKgAL5zj8GFJZbq9QN6
IQsXtBpWRMaef6oAUxUZdPlG2StjfPzqYkmrSqy/6Yllt536FSpMUGpgZp03/Hnp
Zuo7HsH7AdfTFZ9wUALTmu5UzI2KWkNN6txtEwTMfWHUf/s1tnnVf6Ed9BwLvFBd
OK+MMHEa7Lg9IzcQxspiBwXo9akpzh1RRpeH41ee80rdPhGb6lWyTEHuzWV7AEWQ
GQAR48od230P5SoTuXKXJq6WOhhUOL7FoSmnt5BCnAbkhEKszYJROWhrvAZ+yM70
sjJeEjHMg1Q9N9j0lvZIrqx8tSCjOCmyRL1MYLvPSNx9eLLoiHXfFi/2GS8DZi0S
hOvAWgWY/PjrvIInpu/euGtLSb+kg0YDd0/NXOVkXOleGrSWYDgQOeK+onKxCvSy
vZ9nJt4xSzAcXpqyEHVuKquiLTJgxw6tIQPVanT2qUvtq+yZ8qAtO2G62SQ0PgJX
S02n6nHkZqBFc8G9IC4kn1k/2zV4UMjIObgWmqFeQbS19V8BJ80kSktmODvphAfj
HWkoTFTJ1mqgrsoipkrByioaE8ZpS9K8Me9HyynhosqzOP7/TNod94zd0fGD1Lyl
SdbD/NzxCFzn6KIP51p0bCBXNku/DLogB8hXILkRu8YvCJcgql+6umDHMmzpwO/w
r4+1pUPkM+osU7MlNtyFggQhpsq/b6Ftd+x9XIsgWiSBwjRBvE1Hly3MKHaMDDuV
+mGHJxAA8zvJrtmZ+QMA2+2wIfFuKtpOl6YD7ttyAQg06CuUV+RODtRsrfXWwicC
0qbJpgloL3icjQvSBLj4V8P0xsGOZRgCNh5jKSJWXnN5pk4QJKuxJQLEyZgQY3cW
QTyhOXfhWNSPXPN2wWI/El/RK/ZCn5miwLDpi33qQyXz34Ru9nE0oYGDIMpmbCjj
TSft/2ctaNP7yNC07h9k+pKoJbflf7biAoVz6DyeO6yi/AF01VOk2x4Obck7VdC4
lUNnqrOAcpMQbdwLxXKCW27kPtpxH+Ut4Ta79gHFxU93m8tY35O2a040bC9BB7+F
Oh/Yb1pt3lWn80DqlzikvHpwvgshNCP3q8lpFiWa8yndCLmfRIq+nr3bx9RoOUT4
de+CrWNv+7XU/ECoZr6xqVFtiGQsoBZ1ubZn3x+o359tHYx2lbQUfY2slHvkFCLp
I2CBC5gyMk3vxj0DGwG07t9TLJ1mP/C8fkVa9wLYjPRj52sn/qwOTxuuiOOKXP4K
W3q6Q4n4CWGUyZHrIpWdZqigJr6JSjNbMs307mIBUs9OkNOUBogitslvcWg6AkRP
L4KzE/CwFIAuGcctaF9SgNDE/mgDl0+Rv6R3YhrsB4v9hihWrov/3tSX7DDM1v0/
JiLs9O0oh/dN5SuTL4R0z+WXD7ZUIMSszCiJ+YV53jwRyQEgioEIH29LeIOGv8e2
s7stmUnkZLsTQZN7x/K8Hnx9eqxGWb0F1u375jMLVHFOfxvcWy0T5h9ErK8z8Ldh
Bau4+r55dD3TnOhTYnSBSkS6tk0YxjfEg6gpvW2dd8xA0gfqiOzheJztjXXS4CK8
jNBTlbj2gcKtHQLE7UBHkjSk2qm+TUFoDFrnsAJRMLeCBMRVYf5PtXOxLRtxgkMY
eSGf7VXOy/xw9squyYkJiFWzBNksnQ8jq964bhSTH6rRRcX7ltPn7ekeQyxeDZgx
qEheXH8ogbbXZ8IhWwuIDFtrRiWyJ658ZR9+gINd7Omxle1VwIm4cjBFeftMnJ8/
nSu09eYEv1KmyFVKbtACn2/rp1wiQXW7+95Q40cJL1AytyfrGZdwI7AFBTwUFMgL
PChXLjLf01cwMfllOtNxBkwfABo4s8jzpfgYjsenR7OaO2vvAXJtwVWFiu0kw6q/
ZK0NX1Z00VluL4ZWiHv7OIiO4kruoIRBPRC/oW0p8nVAM5dbW13J8gMOJlt/MVau
X410JUqdHrygJDU3tRUjsDoedjnyiRI9eS9NYahHFiNYDlSvSAgkkQD9gg/5GfYA
3qS7DJvsSu4i22QL1Hugu3loOYJqV7zIjuP2N0ANRo12FNOeu774FrmEbAp2N2rW
4lY3aNTU/qvV36k4Dsd6b4SXzd2Y/eJVliQCAgsUCEOkxmQiiMzDsnVWHkDABhem
Ycg97SZfEv1+0+U6fM1GwRGydWSKGcQrPbMHViFMshucFkduQxayg7hGjGzdMB/Q
CheAwcc2UGWhlA2WwMtnT1wXGeP1VyE3w6foDOSTacsAGufSlc9s4W+qgOz0WyGc
CAc4d7emR6H/6gWiKueThPL7EYKa72moigvz1dsCUyFhPOSZMCBR7ny+FiE4TMsd
AU2zKKJvikEDgilVwdP8zCqhKzrAym0qHxgETVKq00H1Q3mTsD3KhTwNLCGIwppF
7SSqSFbXEztzHNBvjwS8wY6oFf5PwPEMMIHyWWkrNJLaPkGrjr5EFI8BKum9SVwU
pZ+wDPeyM/xfpXorw7isqoFXh2hS7oLwCQ1vpd4o14M86tzuGsHaC9L5FZqwDKrK
Egy/L2FCFZzE4IpvZ1SI6qVAL4utp1KNFFm66NULWOI7+s+AmEKINqW7WWQ5/YcU
a1mkNjye6w8XUkvA3rjEW5oUf0OlPpgjgNTvBnsNqrpWoZIj6utp8v+3Qo18CjJf
4tR/I8faPwadO1nfH2xn5llGi3M1aqdAdEZ1MKfAhKtyxeiwxnRtvL/ahZ81UW09
7o9HQJo1dTyje8W/fhAJ3MghV1T11ArGFwf307P1/0D3JTd20OgiZT48O4gbXWZU
53ZZG6rlO4UqM2uFCm3xeyKyrwM0KRaCuZFcRPQP8FYhwtjZH5S913uuG1Wl6/Ce
wB/uubfoUMFEGXzsEp95EGOzYI7HuWp00QUh7qjUXdVZixW8QRdZjeSXPB+pxHuE
AW4cGz0vudhMkUJlBYzWpQvsHgp90HjHv0rzqEH0jHceNV1ignzrUpuTe+22INdl
pjK1NBdhRZlarRtLLxtEOCSwgqZUdmxcE+nyq8kMePDsQYTASd2t6FRSJNLqW8P7
00amMWILVHdjNUKf0cViQaKZV9VVbWKM4P9K5nLo9lRAMVuaD6jo4mM11H40EC2w
UGMkmQDavO4B2EaluxfjK746OanuWu8z17thjvgWsyJsZCekBRoVpnnfeS3KpFHu
jZ6czSst61ERHujWlrfkXqwA690UvPuuW/ZNsCi44wbmfqZuKNEnMQ49PnvvaW+E
Xokqhu1SdHSWdcWAkoFRr3znV5VLGqO9ili7WvnbNaAn/qYxAx1tbsp5TgTukoXk
mJtC7btAD39ZlKYrt2/ePYB5B0pmGUSnZU050MPBq7Qd2Ik4wArpdrUeY+KJGfJo
JFC+yb6d0E+39xDaZ5S4FipqHhCipEUu0GeUQ+DqAOnUq4D1rqGhh24Vdkotf+r8
PjM0KJquKm/uG2Zyh7tJwDVj4NZi9GQcuwAdzvuIY6nYP9/pal2jloAHlByftBNJ
xm/HILKBxksza00SspjVof5JTgwqX++OZiDO0qgSqw3RUuulXNytFbrlb2i6xUI8
GB4FbtCNmeRssEnoSQUoUrpgjEa7xephmPL0LruFBEx9z/R1Xv9gMyT8eUiEnYWN
4N+MXvnl9HbPVlUrq1ldEmtav1XrmTCr/HRoGZ/bJ22xdB/OmAVVHdIsmursW9h8
crF/rSQO+d/fI5/Cy0fWsi4f1UwTnhw1mTiVkBMpClEyd6hR9RKZ5u+Xcs4IXHyj
8ckL4CAYL0F0fNb4RrfhO/1je6xskwVMGlAe1AbQry76KKTxn14WouWXnCl3Ztkm
l6iVVQ1TXJB2FMMTv/5vYe6M9OEg8SlNQFLEGkgBybtQHKOZfysmZL6NroVw3Jho
wljLqBFy6EamkQWUrs8DlBgmpDVtPtJGlvEhDebxhvGCRLNvD/dxzuCSLx98mpfy
kXDpOmRrm/oq0NqffEWExrW1MYZXm593/anbCq9RWH10nZgzVJXKneBhqmif7K9r
osLRG2WoTLFEGr6OQ78pXdE8DOYshfiHJom+SL3H7NlX1DuQ9cFmf5ltKO0wdZG/
2dsghzcpi4uPs+ep4FxtV9BTL33lsjVrMzg70Z69I/m5M5t5D2WUegoGqnepsdD6
NeP8I29LoM7Utv0Hpjwy6NxALtyutZScSmyJlSEOPLozVDroaXicq7mXw11spmXx
3VGn+Ox4MfP8I5Rs6DIYoUZdiFSWvVgNwK/ImdpPN4969d4fbJfpGiDPQoisxmUl
FXdpsr3f/6PhCojQGUhY5bI2sdNiZsTc3m2G/nKmfWOrA4yCdOQM843JIMOQHDXI
3ttoQACbEqr4paicsvGPZ2+wXo5WmruDZLHIFN41BQiZIVLZXvgxByMwUaR9UKju
0o/80BSd8wMecOfMhhVtQk6YjOas8UHEkX7Y81WS502C/GmDo8tfe6kNtNvzhIMP
/Bmwn2wZlp9Hrp8FhW9xgB+nR9bFypQjIG+GzKxabMCEpp+5FRL2w2ffcy47wHAP
i35Q6cY+t2kFBGDSbwO5awTm7mzGZElRUHOGo9m89sgEgE0VPfgbAfiIKybN80O1
ty2i3BRWUFHulOaE8ZFspVboBvxRtdeh7ex8nqgfGhpfJ0PvaEH9xVYyt7DX+Vt6
c8fCOZFtlJleJoSm/+IoegbOHXDdJ6Fb62PnXHWuF1FFagy32fqTYZbCXnGCiGZ0
I8aqAnFQJmaqwgFUJP9/ZVczlC9/wQyh5piNn/Cc7nI0OOwSdPFYMEi94H9qnpv6
LBNrEVIDn6/0Wx+iKgab4+l6U2e5+IGXKemu4aINmhuSarQ6lDZNFnHeFgPvNTm2
U1YVhVzjq5rfJ2v/mqPiMAPNUUCs56B6yHu9U3uruEckez72F2ClFB+zWw1H7+xA
RWrUc8bxHOXHA6uaVlYDm3rzz8LIomYBM6KEzdcSs8Yux5ms3L7UI7NMSwQj9Ad0
UcgasTyodhAI8LqsbkErr2HTzGWLC4EN8HY/tK512gIAIeIrCg4ltmEWnVb7xe6I
TAIwtmBRpmc2HH2rV+chWrcPMOmfhPixitSaxdFqYk+fqAEeL0oCVghe1NGLB5ZE
MGsQUr4TBOyKGmiCREKX4K6J44GUezv01ZkY5x9pKCFcmXIKJrlmnD9QO3lNA5tZ
2fuAqCufPYMvink6i8tdsxkCmaauUoZE7e/pj0qLW8IZ5JeGbhLW2cWKDEotQbN1
Ilng+grzBlAsvY7qygN92C0QAOCIpU0Pr2Qkg4gDbtOf13K5GhOlmFi2JHTP+aiO
+E3Tz0C6hlCkoFpIH98kYH+62Rxy0yVzMi/5gKUV2P1C7LKhn3jRpTtHOQ3Orsrl
5tptypnUjxB3l/D9iErVshzL9tY8SMRjHotaguQJ/sqd8pkfUlIqOR52iG+EpOz1
kSP4/c6JzZbvD6VOWrfbJRB9sGoVG1PNORhYEjoJ+Cqwm8DA3C/v3kDUBAyyHQG4
Yla7uMqRn7f8fF5Bix+vfeFTNBS/yxNkCmDq0G1zTyBQsUCZi8A9mMGfBGCml2P9
C9eI3TgzYhwRmEI0zct/DGJpJ1ie4pONMw2yPe4eF3YvO1v5OyXFPRtw6oSwCIuq
s4E7CeqEBvnV1PEWho7KdpmeOU8gQHov6nhzxKUd/vo2u8xDTRWcttHvJ1q/98CF
aCYV0BLEoRFVtGpjmOhXs8AD8ocoRu1sRdF3bguILgCsHFclD+IqapypRzR/d6/H
wyq7EKhCpH2ce6dLjzTHBLmei6A5dc05CILvhSIPUWEj91XF6YYK6fOMIDcjtlpz
bR5aQTgkKGbjjfxTpY4zwjiRh6Hxfp1IHPObALyV7z13NUiBjiFDrpvH5f/lHpO7
rhalCvSOQkPnoTZhUgkWpg4Y6Gl5gaoDJVo+GNAbRRDGWgci5uZlHWhPxVHvoW9z
/z4GXCh/KJBEcV1jz7gv4BFkBFRmCxHopeuffyIrfGJZr6nG6XmpFcBSxLtVKwlV
bwdAjbfxxI/+Rw4K5VVJ6LJgk3YLQWbwBKrd8cDOwnQKpB8Q+hsGWi1eWMmdr102
WkE2JygTsBSWkkU2ioPrXucJaZcorah2Z8NABdDBaChQ7P2RbjCoFMf9/Z7Jin0b
ddwenHnwFxJYkw0rB8FeKa8dB/bp697YaWTW0FBwnayGhHEwopkLr26MVSvjg4Gy
JUAhiTdWglREP34/imJ0/l7GYmweR+3R7I1pjtvk+YfHfH8TThVrHSTzZSXQ6Z82
RzNg/2ZxqD2y6LXkdN+o+WSAQ0yb2vqvnYhvTVhPUGRrC4zZmVH9e8I6NInl2f5W
xYvs8Xt5KxIJ/mf+lXDbMKeAnNab/Vz0ESRskOWfzk980hVu8Uxin5PMSUgFxw/Q
s46Nfupzxj+YiHRpYpcoMlisYkEbgtcUHKQvM4C5gfwYA71oMrXHHAE2noCTQj9w
ruUGQgH+4O6cVgleQ8580yLo1VI/+OFFykVu7RKlWYrtl79SglZmCV5RnaomYKvM
shBM3lnzaUXCK6bjALLWWn6yFiJvbXcqHqElsblRSFJN5f3SDUMHVhS83SukI8nC
1cgHI47or7rW0J8un6YngrEFdKRar2XQOkyzDJdicT9TuQRwf9cLnvnS3co7+tFM
yV3dgvEsKAGGbj3JdLr9Ue7QOylKMUDqNCxOhn7fSEQqIulGuw7qfZuGtzbhzPIe
Av8o8SqgDMod4P3YUPKlY49Ni/h9ossba8+2R1v7Fw7rqOcPiuNgvIfLe9sBwPwP
dgJOTsUez8RBDSfa1XATb/ocwRHGqe5s0yHzZVlB0XnA7CukdLA8Si2Zt0DidHQD
5UczZQCtlcdqvi33MSIwikHEvJTam9msLQKDrGbOLVOcd02l8s6dErJjR4eATKaz
Fxh3jc2GI3hJJnKQtKKEdGITm/MQGQoLIIwoicrIqg27EYf5hsHyqtyer4XrdEoN
7Uhv5N1whgyo8haJqVYyDu5Z8Y2D0eZe2K83jKEbQ8WUfulG+x00YCJWHREypRGz
uMODEkwUH+zIeqId4Q3eRYbLiATHNA0QKxcI1lrBxIaD61lmmslDLttaWNVBmKNK
96y/S0GWAjKZy5p7xmW72kmrtv1ztgvFuZm8MfiWtCFW41WUDLeC/MAg/0H0415Q
fN0vkNs7DtTPyL8H5/Csb75NuLSAAyBKJRUC1umbnwsdBPq5l5rkXJXjffuBySbl
TOEDwCfg8U3bfWKm4t7cU5Szd0y9PrgIln0c4CECP1AEoY9lng8CKrnxC98HH6/S
bs5j48AKHrWoEuezqqhtL8cxkQFA1nkJVON+QAX2EqQkhKxEtmXHXGolV0JqB4zj
F4mYfrls+Ils8s49Cxr870wyd5KLeQnN2/itgz1OXOgA8FhsNToSdd+ZJP3+MdCe
iAK7b0CWcd6hDR/Ww/0Lzw6yiIIgKkIEynJPenhGMSanWAr/qD9Gpw2M9w7HSKmw
hh/rJeN9z3sryR3x07nhNN9XCsNLKnjA/G4/pSn9EBMEx1BPvDLvZrLahB6JS0Aq
Zdw9MaekU71T6ogMM+AOiCsfGK8WYbzZoy+UK0Q0kEeNxWt6hz4EYSRwctM7ix6T
cb/Lfv+ff4DYFI8gEa6xWS6hYBSSsaYWS081qHkbpDtAjT8coipK4C+9sPj7tWwd
/5lcuuIetXqYt78CvJHmgs/y7dsJFRet9Kk2FZcwxh1rBAaIVxOzbSINwHuDuJLG
ObxKujgY2//A35ugcWNm7yUuVHmlTh85t6pfeMmIGY/GTFk/OyJPc4bNOgOMVjSL
gxoYKp68pqPUkcwGoEAEBXC0quyewmQYgb6ltTEwp7fasashEaxdC5zaDnH6ZI/g
BQD/XmJjNTqidAIeaUopTgnHz2zckyZJ1dZ6Y1jk+PgItT4I37LpxHrZ7gf23GSG
lBItnxvB/wFN980H4tj4tdC5HxYlhz3HrBtnmfofiUWrQswk/NQtN7XTNxlNBubw
3JFTpl6GvieDJwme2sI71A8omrOrHI6Xvr0AsWPLI8Ly3dU7YsJF8FE6hD95wlm6
93Gb3krC3QgJbikbBbef06O0GATbgL6gjWf+Cby5jfwyqig9eXjFJcZZ4S3ZecKW
TJRJdRmIKY1MjN3Yhv590SMAdac2kFgmQv6vF8/CMP0x8m2LR76P5DYKAO7q8Ge1
vEdQkYWx52OjCY9DHfaTb3NkPUp6PQwi/ybUfTXBN3wEcuzR0Lze6wAtt2G5r8ti
XfFkR6tUFDp/pShdCBqOqlwckPVxsoQQn1EpL1S7N82EElOcxHhgNHDnmLEmfE7E
s2FULvTUb9hxStPSM2ne/xhpOKGkniW89By3A3iX28UJ6aQJxIMW8FQc8NcS6FSU
g4Nt5EkR1Xr42Rbk6S84PwI5QyNsOYECKq9B5RqSQSfc50IHBdGtWv4u4sZ1Rt05
/JhsbC1ghvLPGSyKdUci1MRrA3qxNSEKR6nJBC0tHQLes6CWIrAgsDPcC76/34/v
ru2LPmY4skTVZAJHUKKUa4PHPH+IS6DLg+wvh8qcncCVT+ByCaglg3kiW7lRHPmk
bwjP3lCBgcZMz6IwxqUrrg3aPJl+NrEcl9vNpQef/MDeeu93bS3FaGO3Tp1l7m1l
ilN28zH6j73PWG14UKl14I4Z79bkB6Cu/qVD1kFViv6CZuENAxqGCFs9vQ5gfAgc
863PkY0jPFwmniKBBpKJeZ7grohQ0bxrdS/9GLemiybU8OK4/dWOXOD0BjQHVqHF
vGqOPjbGQt2pM5/Pke43p9QP7zvoH1ko6On2OqBpgX/4x7lWdhqq4srmnGwtNK5u
Py63djbOZSs6Rv7Dwj96BRw09LfB4+9FN7ZzeSkVa2raxt6l59Qd1iOqyz8LqDVT
4kuimBen9HCZhkGElAsZk6WraPS+bY2Kp9o0CNjU5vbAfPUHerfqCPQpXtyWlWEC
aUS3VCBs20gn5AoXLUGaP9gHDFhrqNX5Vd0iHufo3F+WDammFq+qFbJaDwspqOE4
qSdMiXqmIkZAwFVYVokPT3thvWP7ilCzoSaXnSDI5ashPMD322KDhuAYuWu6I5rL
6LSKFocPWd1rBSIWIjaIgl1mN4UsJ+8h+/92RNCQ7Kv02HJln6XIM2SwbU76mP1p
odXMpNRbnrDRKsj7Nn8GY9+3RZOnCKrXgv8c2AHXW/yug/i1TOkZl1K0jMK1Kz9X
CAOaYZsGmncNK6pOqEwqwukDbX62hmqBRMi7y/L29xP7QbKcNoy/d+w4dK5fUOva
VnJjS0quhM1xaX0ovMaGsKOcRVK3WuUgGs8M/e25Lc8xKff7tlzb2cZ9SCYmn/ak
hiCeqUAP+vJkKSaQEXmMxoUus5DufaMj6EuG3LTyrxRRTV8Mt5rohy7EcFl8sxeI
U89wJsanzLiXhTkWhske0Bfx0j8tFBN/5oOKrxR0P3K+dOaMuZ4PWrTuwi7B21od
02Q2aPntG4bEkDFxIOhMLOyoboe5nZrRvgwvb+fH9iFxPhA3Mn3DwLe5GzTlwsz/
DnQlVPCKLs/4TJG7pIdmgvU9B13UnthGCP8V1LEHoQvyFZcpOFCJv12kELISmhxT
leOQKy8lwq7iuzZfIWZsfvoUAn46cvbuRCbmW8nCAywUL/TTy/z0/7NaXHTbZCIu
IIr2VuMSlAjlRgszQISSuwzM/IjwBIu6vvjFqi+F2hiWevsiAo7p5j2a8+dQbaXD
Sj7QkQz29NH+2HCocDvDCKAiyVI7ZEwmRqxePObFHp+eUzlinGzsm/CfiMmbxXdS
AyoAGpEpPT+jTO2rswmveHa7vHdnLHQq57fTsSY476JqGlIBLi7HvrUTU8V8pmRH
iw6kpugzufREi4z9pvrbj08LMGxhCuV4THoVg8ZjqBNSNSQnYu7J9cxEenOAj+nZ
ymTNDNko+fWy2WrCppgTZLOWhZrSwvte/BJdn0i6bY2I5223BXbMpRb381+91I+N
B7rbXA+hJTElK8P84JLZjdeHAPy0955y+kdRXnLVZMd2MEFOOkCLETUqB6bwp7Yn
hE6TrhGeKnyIKxY2j+/3IYz6Dao9MqGby+IK4dwPh8lGinD9hIxZ7hGa2mftmtDD
mF4vwv3qthxeNZAPO655QtjfpnJlW/D/pGJtjlftIaehMD2N/HclneYpuaHBpS2T
sx3uhTdzcW427WQyXC0JTPLez0An6oIwbi+EzxOYAntPJXQHjdb3CIPPJ948JK3j
pnFMlU4TeLSPiyrNiTazsE2RQ5suuOvKvF7jmA4Laj1hNhy6nu65zwaiv3mRayzR
q8Y1SgdEFaqJNwOrsnoDxS1JBhdf37Lb+ld784a/hzC/fUQbFqQWaiCv9JEGr+yc
6yAx2GIJ1TmSpGfEx7U/Pe3kPyBlL5wT+bbc/w3ZJ2Vj391jSQ8q/Bthm8sGoZ54
mrxZgxJY8oDntpZXmcEaRwcqO97gSHcXraDdMxDLTId6DCptdYv+3qw6sLdQgp/4
LrQad1JceC+/mT8iUOWEHBjJoN6S+iIeIKIC0I1Fn/UiYSbQXIQY6HeaFBKUGvNC
lGX4J+ZPbR8I5vw1GfDWBGGrWMmRmcs0eQfARFqoYCnBJqiXPr8/7BPNtjrEGLPc
Fk+uFde7vy/sQH6pdymG7wzQvtXd/oO5PhCObozZDYp06BYR3gjk2yKzdsraGlCs
AweYydvIQ3lkjlqsCehpWsWYNidLnG6hMbc62VVlYT30UEb/wDLU8Av6d1IwnzMl
jF0fKCjJlRJzxS6szBlfYp+aeSM1lPa/MqDarSWzWOVYS7mC3vyFpIVLU2SZBZCu
v8yKOmfZd6F8kSk6YBc8WhfFdDX6xuHx4BDG+azuGv5qq7uWGIjRCWxlhg/brQsJ
/hdKfAhDV5bfu620r8hKQhQuNe6hAkeH9HUAypFt88fRd9zv13bqXa9P9KBE9Vxd
0nIl/GeTdXdb/Kx3rq19sXOkzVuOHlQpa+XQipDojCirS3/vWMfCKH1RDbg3Pd/N
Wdd/IS9C039vvILw44/2fobvWmlvn2uzzci8pgwK43CBuKTsEDe7ZbUq1OiviCRR
PKVJtMo5cqdNV1aj0Zoci8LiPzTYAQX8dYbHEQn2nh7uqsOWfPR4505AddUWlrOR
1Br1wiA0lEvqLOw1MM/S/CFX9CFUowu7op8lmSS8kWXvINZIofjsDqw3ta4YAfxE
RQw8JuGkhlcPwzxagrPZgFGX8NkUAnfW1VSPt6tadwdHFNBVwoDE2nyeUpoYQ8UF
5QjUSEkVdWxV8hrDWnT2eUG/6WCmkGa9ziF71CBt0Fs5f5o5t9K9M8/1ZBZSz0e4
6wwMzbFR7Js99BS92NyPDoDwxdgKkWznozHGeRfUDA9PHT30twokWCceCYEFt/ra
o+J89/0YNGb7e8jaPQAliUDjbxTYVA+NuXbQwBBXEpRNKMuxndPeV0GQ+zgbbQTT
2AFfnUhHagj4Y+ol4ZXMSphns5MvgQEoDMdrmYm0fid3VeaR48Lf93dAEd6ebEee
dY7KLiuKJ2gM+LohJWCg7Jt+swpS4uEXZN7J86gEFeBCzJDo63pSwxK0tmVuRdtz
X2MSb24/Q+Sg8ZyF4uBT07LHK9PZGyIaRlsP3tCInt5moO6VbfoWyv6lM2FlOOPr
gMC/2RgYqwpNElnYqTagb7reUCLHO6Hy7ay0nT0s14JfR/CPEXx8r4hOes2u6kcJ
RA8nzHlqFshJWTutNH+h5nKV14Vv6yLIfG3uwGRm/GkQ/aQvOhsL4/3Xt7ZLfixC
TRsZ6JU70Ltv748KEKGBf2QgjYX4/i3wsAy8E8nKszdvmXHtbJEyaNenpWWKXnSa
k6T5ZCYKVX1w0mzcWN4HMnA2NAgy0YYMWKWVcDyMB1l2Rp7pkReYPaJHDOGAVs4Y
w+aD1i6bFYVBgeq/3QidTRcT3rQ2EtZ2ADohBA5RTX/nMcLPwqsUO8ih2EI8Yjpo
9wHvsyv1fY0gzLkCgpOFbUuPqSYd9PuuCz+vcVlHXjNcQCyoIP/Kb2A+kMWWeYu7
vPXB2DR5yvV9etfVHGp/tiObFcPuldlj+eNwpzODBhPH4NxTkR6gEOka7MWN9TVr
m4ikbbnHLpcrwUXa6CNR9jlGsI5DjL0nB7BPWHih40as13gyZQl+V7yxOLu9IRhF
v/VGuifmF9I1R1+K6cXD40XvSHxBbt/An+ZeSvKxK/M5vZB3aBGc0qc/VBP3JgiG
qDF7siLk9W+2O0mW4+J909lVDExev0c6dfPWV905Da8Mfr/pLWQ9jgQfnEiJsCYf
znl4Yay1DXhomCrZ1PUN/DHdYk5CJ/TMnmbvo8rMQ7I65iPph602W1u9l9Sw8SPF
+VDMmIxKffeKT1lZyvolWUXIo4BYl9YCpxlYhgn6Ht+9S5ReLG0fXhnEfUKeG7gP
ikr0w2Gagn8eYNbz3luVSNOrrDOg8Eah7KOvzFJ7cqAwQyJFKLP7BXadpxqopWl2
+Ryi6uf6WXMP9Ikmg+Rej4zMS39oC/4WQJb6RNdyY039HM2zInEKTEIO66Jg/xaN
X3QvMFAbC2YXiRP4mVpnn+OjJXbuCXhnrocUxtk+trh5NUFo38aehzDqJ16aj03M
clfRz6XVsumv0KXNBEo+qUVbUHcCfPe8G5hH2gmt0ek4Fdqys/aJOZD1ejdhQpgD
HZFPT7Empo1LZgWxX+A2zm5wqiqvbNkXNpwUk1dxijaS9c+l6Ko8Hc/Iqm8QYeNr
VMApVid3QyLOwqiwxB+Itok2psk73Pvjue4Wa1C2S00wep4xviIhEXijBMQrFWa2
Uyv8AUDvlQDSq01xk1ONOv9qgvBq4ln2Nix1vMJoCleN7qXGWitMRtnexX4n3Zbu
eIO7f/HQT4KZHpL4rLjFPr3PZSyY2eRMwEofOXWvEztJ7Fp9AX/uohw5lC3inmHl
SWixXude7+3earkdpOkMnf8oF3kAQ8HTkHLaNy35rYmQfbXk1/4Ot07/VMnjYqGv
67Eln5964n3610hs93VszxfTQ1T9HPdbxteWLGashM0aPvINCNV9vn0IjNpdZeuN
o+WDi5iYTDclvpLWp2YEGsOH4fVMcnpkqSlfZyJ5AV3726dSEn/RHZ2uBLklLHEH
iEPEpnCH2gcaSjmxM88Np0hbmmw/gPzB3wboOShLNt+dVbm6qT8ukm+8YHLJnW29
WU11ws7ASwMdddAQkyAqdSIx/AmwZfyCdCcJnx18ai9LZp70iYL9r98id8zw7+0p
KY5Hpfl8IDNPj27TFIH5r4I2G1q2SZr+0sqagJjP7ecxMr12f11h1WvDZtKGFgkO
HWTcpfy4qF11xgNdYf2s1CVNRhL8XIU6+vvj7b/1LBMs37Bz1u4twmIrL+umzDBq
T0EcZkcyCBnAdj0Q7+UluDFW15nsxYeJnpmL5tupDIxiL9eD/0rGBG0N0/rRc9Lw
5gQfVNH4Rp4C+qzsf1tvuqiY/NiPTQ7HWb29oe13+svouJbb2BiEDHnDaoLVOcIS
Z+3rNjgdJhC6IBGODI0g1AY5Nd1IF7yPNd5V+DSw4x8isMWXxqPQjeMlVYE48faR
My1v0E2ez5QKl52xlU2YNe9Eqlnx/cn5S8Jm1+ESKswPY5ggkVjH/gxBfWd5LWaG
tW6OEsMVBBKPdAmeYHVYG3S1A/oxbG7R3Tu8S1a9hnRzmOCTb5mqCNkGQKbsWcRb
C7+MKRd4a/+NQqLlYS7Kh9vRJQiBk1fAqBNUqZHw2UXp15LPNU77qgs4XWRR7E+C
G8IpgKnVgms0xl23CnxzUcHYQZZ8fqp81CsTPwMte6qVPdhGp1Zdk6lHgL6JWOtv
cwiJohf25XtxoU0cBGyPTvrnQS3gMx3KGbocw2FG5Z23SPt1yYZrtjtb1DAVHG/z
rWx0ydFu+a7OfpsB+o4f0cBF2IdZViAMOfhgLpg7ZU5eY8HOJ9C2NExBGCgHG7bz
4R4GPYc7b9Yg/b7ewAK2MCaoNEE8+N1Xhlp51ELpjuN3AaY83JIPVnJTpEpwP5Lw
ds8Xj6ulJ6of3AnC8KcRJ3SqaP9hfKONS18Po8gl5WVEpopN3mN8KoVMr5WO5++1
VJ6pvH3x32Lbvon5kAgKEyP5rB8pK0e5spnpQHtEZpy/1K3W30Ldr5V8U4x5d+KO
ZiMXz8keu6Q2usohLNLDZgkQaoo01DsWuU/K8oQH2PiX+fIZtXTTD1BDeAUncM8r
bPyKpWwO5efhhtGDzILVV1r+mXcBfvZyXV8xwnCeh38Cdh9u+EWMbXJrPDm2tMBy
eehIQ09v6vz7ogfxPeaqZAWWkdoKlzHSmMpyJA6r5XS6zjAXgdi4V29Q1AV/PPOy
KQlbJydzHtTC+Q1VaK+YZmAHaudTSLLhlvTTthRoSdMsNJPBaalhqei2NiynlWe0
wB/81ApwavYP8rcSqcGboYDfqQg6MzcAJgTECAJvQaC/GFEu2851zeaLe+uGsQ9K
ma2+z6UzNU8hQsLzPsSvPwKe5hEsl208BOVsLI3uc+pS7Xru0xpbFCSjUAt7J1w2
1f2a1N7qGOyRR8FK15ZzCovBbmajDu7d7bT6ScvZLBzInsh4zWesnHpixr381GEj
ttejooCfN7wUc6Y080XqGWnWtvyo3XPleccPHPW/z9YhfnvWt8yeCH4ntpH4A7jG
S5GLzElnPkmWFfsqPXmFl9dbF21gqWDoctVHoUP0KWCVimqVqEbsJj/PxuRDT4iM
OnsPB/DikbxVZK3uqM1tujSIAZsJ5Ze3cKdmwF8kmx1dAcPc8sF0vHlMtGFAxN5i
EQ2/sGcdV354kBuahcffJgBHX08QbzcKSOaq3INSU7MdPNsbUt5kvWHlyh2rCNEO
dgZhAaD8S3e+bJs4El6SO1qcSGSgVMCxgobuNKTklaKXXhtqIGjy6V2eKdvYO2HW
iQ5jjhHa6paZQyN44/XZg6NWY5Teg5P8U1LEcxISAvyji69dGIuF4/rbu+DT45Az
RU6BkmOBNx86XH2ActKaJHP+XO7TSr11lOy0qmtko/GS6aUmWGl06mcHoArs8kQA
IBqDrntPDj7fDdV9CbVtsA25Ca0fIIgGljTOnt6y1n0sUgfL0O61u08bBJ6eyFWj
UsWDS7aF3SDJkTnN4zI/2nq+9WcL8MeoeaidbSxw0Xw5IJiN9NAk280XTlVoXCfq
JQ9ZFgLuA/DcrZAe0TG1sexifwMN1lulp2AsGirtX6UjTF9OyJZkEX0CwgxuvX4A
jSWjxcvn7HRle44Mpo15TZPSgJPngyOVmWxLIgXk7phtnfE7eKUdoVRBCAgshZdv
aSEOnEbQF554Vb5TskkwzMOyUZLsYiset+/wRSz1tA21aRATcYl11+wTrwjX26Ah
Z+bzHueBZdXEfDrTeTBHejmn2OM49z5L4BCvNOZR3KRoURvfF54G6hp+pWn0n5dQ
5bkErsXLTYvCo1DVSsGL2vcaq6cUymAqz0s3I+ikQ3Rm6+uQxx2hPpNQwq8oqVlY
557AWX5wK6B/jDbz1ZbAAapOOZ0aePqDcUEEkm0UsZH1lEOtjkbOBiSNCvo64KAt
aqLrL4xjCZHZHhIlRL2cT/fasiaZlu9sumNUBO69gjbynYIdmKFbuU6zzOZWy698
JlJNLb2Y5d1gdW6snPMEjJNYTDRIKIUJOmSCei/z5cdzuencJklKoJmUK0wpy85B
FAofoOiGSnWjorH5PCpKV2beDVHGQulqwmkgnrQmA30Td3PG8v683Fxmg5l1VhIG
B2JtCyUSwpJz5ykRg8oqN4+7L4vUZhLYxR5cnZvIFSJpK4Plw5+MCAur3fmoKr39
sq/XniPF5Si5W/HnxycP9ZB3CvtclBiMJk5FJDK6FwrZCp01yz11Vs0aGAl7Au+T
WjZ/Sz1J1e1/i6A0+MXTxusUMqUlKmuST0LgWLZhem1Fy3+xli0Bo5MjO+3c5PpN
bayyOcG+GGfB5U2HiGZ+kpPEoLfQKOAvZpJamBnAmlJVfy8DfBhL7BE9kb7P8S5A
GSAU2vU0apYEldngrs6n399Rc6brJkXPjniw1qEIbaJV/FH6e80vVYyM50NlYQxq
2/YWOz64gW75A+NKK6Y3EbFVYC6uPdwNm3nDV1laglrmpVWUqbCLnCmF/Hpt+vYe
jiKbAG3lJxg9apHqkWjU799LJBBheZyZPhvV8SzZI+pRwrqNo/T8nlLDz/XdMe86
IUeI2LUPznUIok1Ky+wbXdUI7Ubh24eg4cU1BjCPQVNoYZkvDa+EWvl0HxGACcPo
RPLFU90TBed4Kp3jc3MSL375yESb26YAtWwSWS+L9MgtGYJswbjl/Ql/XG7hC3/A
bvDtyEOTT151PytGISve+vFezjI4sZS9bBuiqDLDlA8ES8KVB+X8p43LEQT5+eY2
EOATSeKAhkDpcdcZEW6ODpw3yA6FC5j216GT07ERoQsXTisC4YmIAJQTfg7btwak
bDnZ2CPcZ07/tC7Ssf3f5L3ZcFCepJCeya0nEobh3kGJluELUZEULpsIlVc+6v1c
iPezSpLXdYeYmnKaTGWF6gD29A09xzxsa8TkrEAwnnEi5rIejOO7mHf6Bbo1i+KQ
LKVThANXYJseRr/AVFiFYfMIH9nTcbRqbjnxvW/jeWZ4FwHcJOHqNKEXO5Yqgimr
7Eq+oQYntO2D+404OwnZkNOcmq88LwpiVPUiEpyptCDa4afi/z99Crzu7xqta7Dc
NmZEzGuqHJqaYzvpV8tgl6gQm98/2uES32dxpKfxuY7PfylRPCUK1U++V2WFj/5B
puIZ/5orjctqRpWSwqEbdaxabh78sU+nptD+cB7TBvG9G28UzG5TiLxfk6Vf3eII
LQOJPfAXtp5DnpjFpZuASGHAD5ZxfY60EbKHfMkDUaBgVBjoytyEoRxYvV5LRT7Z
uyLfzT6OPfRRwQ1PZANB7oYY2DznAC5jmW5ESLAC1iTXplZYbne5jV5kVoBdS39z
ccgrwEy2Fj3O7FXRS68SmP7tmg2DQoSOnkc3HTcvtFRPfZ4a5CJdouAEuCFXtIzr
NZofoAO2JlwNf5wgdV8wqRuYx4z6srcyXNYaPfbCxTEalJF8E6RsclTwCmNbZgM4
MVUnQ1YuineK5+ZuOcg0qpEK5T0aFTdMEWUK8o2f+jnG3yrc1CkdiRbxdNnJBJ1Z
pgtgki3yJMVxnSmurU9FTf6YM2N22nCafFUNz8e/mzoXNHWquLsMMBZHarDvzAzj
PIeUYwCotZNrku+O9krCoip5f3nSMaUDWcjTe5+TMrt0pQwhUj8/YNAEtEF0Uq0M
cStImrYn0900JEG/E96Oco7xijTwwmKwyf8+eb3HoVMKMbGP0sDG/MSGrsDWde9B
1jFye7k/kBGkhHFEvwWsMrCcqd/+G/6zpWqP5R3zOTWry8Yu7xBnws+feGgXydYU
Z+oqPGCTlaVuevgWQ60PwiioTdQrIT3Z9JuyuD0YbEFxJ6t/VoWqi8j0Ljxj54cd
wesdhymQIRZLZxddbg+J3TlTLcclpk1mBeRe2ArQII7fdXN8FgAot5xZtQ5DapUy
lphwVRYpQKtzihJq4Do7F4FMV8CZhcpLaz0DDxxr7xA1GnLEsxkr8KUukGOzOvD1
cN7TaazpeGeA2wkgVDC9S1Yj7SBJ2Kta8ocILanowRsLkOh3o6hLkbkANHINOER3
2vvlr6UUXb1XNrsy62T3PnWyO7zGw27D0Op57DnB91FyX9QvR08DAybpSv3inCLM
RLdN0TlnrD/K3JmdzW3NIAZfjFXkH4VoKGiibojPaV2nGxj8n1AS2BAmJcI+1H1m
Y1p2pWr/DxmfAFW4wYqS6e+6ike3wZU2mlVd/Bwd5Ixg6uVFXHeSQCRANQF8bdFW
ARuDXY3OJpdZzip0g1bZgjFDnBfWn4ItFUEWf0c11I6B5W4ost0cZia85yZUFTKU
uXZdhqzdK2i6EwH2ySCk4rNv+kxN8s1Alt4cLZHt9aWbLXFXBmaq3r2ARCAhiPhZ
c5eLIQGZIBVpZ0JH1QkubwP/EsDUxXECFJGoxZ9Yh/ycgoyMZIMDoEtrT2Z3frk1
1uIr78b6D0KqYVoUxVNiZ6Qhi+P4fQm/60s3TF7t1xOj4UDMRX1xRNcTRDNMwj2Q
aR4rC6ZQrB0vWDT6URQRc+jUW8wAU3+HFtw06l6jqDHZAlmi66UBUQSOUZCkHtNj
tL5799CExMm6c42EgSgnKfHi2qfVYJX6DF2zzi2oHgFrFdPfRpNVXiJ4tSkuVEOT
nJ32LpZNibcDhU2nEpHocrPEDwzXzWgu5OyMQRotvqQQOff75vgj3Ex2mq+ABaCl
NEKxHIlx5SHnXamOiL8vg5VuO+gMdscfq/1vuy9HyE3po7uYIE+5aemXCITir3kO
58pj3pfx8h/eWI6JMUmCtLG5jDhjzirFMi0CibEGvmbfwapPgXoMb5U7QqrRDp2R
wemZDZqgnCitBFtJMEiVYtV31GjTG5aoQ7Cgnw2QlV010LujTfhA+pwn2ggmE5GT
CZrP0PY31IxFyAfoxWcVelOr+FoG9EuRP8uPdRkDA2EJPuOfjqRTBiXwKJN2tIkd
sTd2lu+1pNs4K2kQMcyN28JnnJTzo8Zl1WuAg7xJ8yDdN63z6KdQ5WRUPqKLIyQO
uJDW3IT4Gg85RfIlldOgjFZ6uajZ/oHcKGDM+7x3+Kzm3zfo46NrnBXe//r983AL
LbIMh56iOxmVuvDzgM1qZ05Hk3f3+CAuMMy0Xx0+9RRZz0an+qwooIvGnrLOpN9R
GhMCXhJPR9znpMLAVWT6s3j91zhm0SGRu1U9x7Vl9DZW0k5mVrE2qYb8MU4lqIhl
sn76bNBPg6ve0FGxLjwJgpdyGK8enXUuwcCUl3iUh1K8iwMi9L7goNPwi2d3cqtZ
EwWAS534Dc0tYnleraW8x8WZul3LV5QF3OkUdUTwL4X2rKt/qehaiav+vP6CIENR
Q45RTNX4PxCe5qD1KQd3z3jxzAZwXebMO2Q/0R+yqrXm7zCzq2bqMSqKGsvvp0Dm
IYHCfvOrRFvWbhNgrVKACBpToVTG7aCPso9yTnztfi1zEvNZWWiQbrzBKmZz6aOI
MPGzTQtz5aXZkfURF+k94Rb2sPVSnZ707lEny7ZTFJ9mDxdjqZpav4mSSKfBY8Dd
pIoMBM2MYanDxTgAORjwVI08AViviZVfbPXczegPHsAYFttSGA9+q3lhVzwDFyiW
XxiBHsaP5Vgtp8NExnwVGXu5GIoyjGsQQ3mnWw6eeyJq72AUfBfADioOR0vdWGYK
dhsKsEaA8pASwEbBK9LRWGTzoWWK/WfxyT17oE+2nGKRKpLwtDGEugXn0O/WG28N
QatOFfIbDlNIUG41ZpKMuSgna4BvNj/187oVvHdCoS0ZPhIyXwOecBx8a5yE7Mgr
+6R446cLKd111O4kNq4Z2RCE9tGwoyzphQK/HPp/US7BVVempxECz7AAdY9mtd1h
4x+qbefAqRnOLspkOtsG4NIkCZk0kdaPfFuXsZ0gw/JuQE8jzqglZ8V1dkwswIs9
foWI1pidK+gvJ9bOWiQ1+BLtJJWgqBvj1ClDelEsU6av4RnQfh4/HouPRZ1EyRPF
pg2/lNUWboSJFoNjfOtey7A06KWduHuVgDcIEzO0En0Z2hqDrvGZXeUpD0jfI359
u6bV9hE9Zb6W+c4SeNZU/8Xk9B0uqH7MptAykmDv0yT3+uY7mEpfAyI9f0B/bTDo
67zvfQtkL723RZuHqnR6jPSi0m2jY61g7+m2jp0Vi6EO7smnTmLUJHU+jgfHt1UF
3KpxGQ6Lt9iMWFnjgtS7uewmNX24biJPVN5D6f3lkCScfmBbWPDSkOenyspP9hXv
2jNHi5mvcaSYeN/FJSqChpjkde1fs+TCg/U9eh/E+HREd5CqdwgYetei7SERZbKK
fwJmc0fyXYEt2X4ykA29ck5yBVlAJLqthNMdzptZZRoVjHL/+uf6sTeFAEoiyKg7
6EbzDR1YGBi0JE6L8j9GutQBPZS0pSRnoWIAAB/g09K2I5x/XnsmuKWW5cTbm45b
9MCcNU7PiO0VO7DanWKQ7pP8m/jmh7Nbw+BT9Y+SfrnULEtDoVuxSCillCZ2nNUV
jBISomX0NVxPjEEWMKDEJSWR2pEyvqZvMzzggMLFMoqhqftEQ4B1G/LDCMSOGEOt
Fqk1N70A70kNvLtOrR7lzBJHKc6s027qaonQMC+x8v2zXQK+nuUuWmKRlur5O36k
QAvPPVhYFcSMjn4TaeOUdKfzlTRXaZIJt3X4jQwDsQ/1O7nn2mdtjAAPTAg7CMIw
5WzNoAdlvCMDJQx2ZjpgOau4zZlUVJgQykgqB4Gu8HN+1w6w3TMQUt3NRKVo2dJl
Zgfuh6Ki3QFSvIUc1lMf8nRoWRK/SYbTbbcgFrgYc7KAhkf52ZLicSRPh//ZoGHs
XxBKPtFmnejxtivMHIu7+RxYZ+lUdWBHMiHt+o9iYOFgcyuaAy8jKUX8GaP4Ur+J
5ITHvIS4wXoMRnm7FM5t6XGCR1wLlAwZTt9A8n+GnH7fWdj/xyT9EYmIAvycN+0x
nvc6jezOs6Vhyr9I9EttFhLdNStEBFz2rN3O79imKpxHoPg9IvHA6/h4HbQrp2YM
iuywhpUi35oIgXY0zZc9Y6snfz4vy7suW3UwaZmfBJsYule0D9pOIfZut2Q15hNy
gxeYNhjgtsCtvBS0O6W9/bkbO5seKyQpATtSV5opwa2+5T9Kdh0ndOyQxpvstEXB
kcaHJ229tlWpu9AE0XbhDPQ8yLXfo7XyFWLTXRDquNrhlXfC9LwS6/mXiWcBkRHt
DhqOKPAZ2MY3Zk+UKtld+8uP9e60HP5fuUhXZAcJqR83LXAkAn8W1PZZZZIcd6NS
jTt5d/NYulGFcvymeit9i99Zt7jLElPDa7AtNFDxhDZrK6pEQ4qSBq6JoPG1uebM
ewg7mwe+fU0h35b8ATXVIhmfADa26qLZ+MOK4Tfcv+LKYGSxuPGbI8WAaSCh+HWj
/PEJ4o2NLCndxXoCfnXvMTeSvyyY3r2/43R2vLyHpyPN/GyowTso6aDkff2h85ye
urqndfeGNoDN/kGvBqZktPHgXAAVZpC8B/P4eOAcLjQTAmfcEk7GvXzY6LLNMQKP
f3HoWip7j205JZizRwReejA59Tw+46xCXFvtCAMchgrEOOJ10cw6gPuBhrfM6Sk6
eitMvdG0cRANcxQZVv+FhS/ojjU6aR9c4UG8X0sFVcQwGlNs77OC2aP0BlnFJ07Y
BRGNW5a2wC6PdD1Rs3C7xmqesN4B5lNekLiZ9KhDnywMLUK/tpBcIyRsMGnUQtbx
8tgEoHoyB3FwOBVOkHJcgogUMP/bKzyn8CXMXZ1vQH0kO7jBRJl+SxPSHPOaJY2U
H2GJCmq6MGPDXWX6CN87VzLjuHda8M+XZd8zId+5/cf5T0hC1/c4hS/e49Bm5LwI
8pTD5pEVwhcWMWz0V39NNwAjnYhhkTUU8eo8YiH38s2Niis692x6zTibesxWMzxk
CxFGiEpOVxY/2cZLOyVnaBZtH1bL+Hb1Yn3H5B/a8lE8G/QTY1TYNG//+TVBJm9T
9qEZ1LR8OZ2lquRzW+TCQuK1CnP7gTUPVkp3fWwp/zT3fDrOxb2c5T02THXur6Zo
bUgIskg5YvEgah9m3RdsZf3D0aInE+a/hAROeqXHTsL2ZEfgEBjFLRBnt8gNb2WU
qSgS39ifIDGh3nE/QREr9teSe/ft7FFbFWXrIgO3QLT3+nB0CzrSi0I6H8g5+Aml
E3XuPU3uuS2psHtK/6wWUjEvJLBH7DvvIvbmcDbAKkg9Dm5Aoj1KsPn3IHKqX89L
2ee5/OIT7OCyZ6RAoFud0gDWISGLRYvGFYMYZ/vBr4NvYNAIMxcf/JZqE3h3BoZj
bCLjM5aueh7C3+X4C/sfluWysRk/+OFM16kvbFjOaOsNDOhqrRS8SBkRerrBjEUj
OhWaT0Z0eY7byz0j492mw7Cb3DDYOkqhw//xZbXsmZwEVgrkxl4nxKGi4kUl5EtN
hwWebgFxGnPdge1h1Gyv6l+huDGtR5KIcrT+tJqlnq5CTuDqWXn1PzNsQyFNFDvJ
tY7MBPVY+6tklsZuuaaFSVcasViSbKrVaDqQZNNM688oTkWTGLojen+16/beXgqa
Q14Ge0OFjypz+XTNdApRgBkilbv2tBXOo0Ez0zkdAeuPovcugpeyTI5OAuX3zx/6
J3Tw37h0dejjmePCivFh6rMV9PVuoXrRgNkm+NEzTO9qj80PY6fy01ezSnfQ7VuU
MSbTPfGODqhEi7VooOELAWYrDdmMuriItv72lnmIqm6dYZy80tJiX500MfJm62B6
37voU2y6+Mv9h1dIIF/oympShBDK8waC/WRkmjJhW2kuwNEzz1GgzsF6ePlD9eGb
9q0NTa009BMBCagwPt2+WSE7zchdxVO5HfG5bWZeWrCav0oXiC1wV/ludlJHSe5Y
kAS+kPTXHSuPqk4TY9NqtzYxsNmtP7/N3GDaAxeWPUFV7MEcZ7bvL/PW7T2l9BdR
+VO4Ajp62DYd9iLIHP6LJeHZW1wYFFTKWnadXnTI1RUC+FbnjFSObVBCCmJ9Fiz9
wBcSq7imNmRpjnuPifrvJayIVvOu5oh+BM8gCOWAWwoxjTv8QYaTj+7Sg+rfuomi
SkBTjWkHJE6rVMS+wxrJndBwa0BB1IkZEHp3gzr6eGlLPRLkvpKh+4ZojWB3SLzX
F4NFRvT6zm/WmmD01UYRT7VG88YdjFtxafY4clHYFKdcIIJ1yKw25oUq8wJAHhfw
JZKTh9zLGFkDtry9jlZmQASwbuud60p4vuCQSzz1KBMKZGKflg8GGyXPDz3UrO6k
zm1gAVxhjF23dGSweoSfCd5Omk0WGf/Tnpe8sYBnnj/hsXYtWJCUbJkY/LqHjn7H
NLDNDiWrL3f6AZbGiBIjCt+c0xiyy8UJDNGy9bbJb+hCPAgV+6/6g2boy1mKCKB5
OkOCEvMtzDG2ieY1gh8F7wAxsehDRuqdqo4SoRktxlNHFbhwf6Cd+L0Ym3XHbx97
P4a/rfESBNAvggmCrdTk80BBJMRHAfWFznTAbO7H2QlNGDbqEXsNC9O5dSN+hi4C
ZzEWVXK9G9iEarlZVagQXA+8ZM+jZIec0VCXcNg/NIKT1BJkzPcX6jsa5oHqFlqt
sHIs7rKKBx0l3Hz8rwRzNgfCKFszZQ2mmz9nLvJJHhfJ/1dwaoRN7E3gonuG48Ut
Ff6pYtimgbRrGmiTAptKt+O1CPUhCwM8SvF1TXhHn8w5rakgFFuOGq9qtrV71Z1+
nVaKO16WSwe9Pc2NCb0NGgwAVd6KXoF9JqCJDiMMqMUElfsYq1mw9DzlICube1JX
dgNH5UozX7XhchracsweNMsTfQeUzw8inv9Er2SY/Uy3pyzJVfNQspYXpViLTVr8
qgf04zpSJCXSY34Wlh88Wcug0eNNVc0cCr0h4lZc5AOTZKuH8znfvEqy496/Ra8J
/wbDbeoce8G0lwj9MJImhyjimCl4jz+bi3RDpqIVsh02Ryaepw5EGwBvR4YR58FJ
EGxi2qFzQs8kMC87WXvGOUvkXsgfvF0FC+zo8mtPCaIONMt8xIlRnJwegJW/gOMI
qUOPJddPsoA7t0A3gOedSmzF4ylDBQJ6YkGzoYR2yQH9YGjXTZ/i5JL1ISMC3eij
yQc08CjpVeTiv3cZLuJyRbB1GXOa+EFJ2Fw6ZSMYYBzTzpCvTE/BddWLrh2DfRbj
eXFFuKympoc0yH/saNYqLlainsjO/uc147J6mGTqxCWcQfcruu37UaeOgDF3gVsu
Q8OEGoXpGxlzr7Txmv9vlNhpv2VSm2vL/jJ2HiOVC62y7TlfYAAPFBJmu7nRms3J
OqWVZMnHueSN5Um6Z3pVvjWGAbAwY1SK3ZEs+rNFfwWfMZeXHsXbK8uVUzy1cVny
THXV+Pvmc3wjG5bHVK2bVHKRFyxo9ui5/rwY+oiWmQtWZdeQW+3xZ4GV14yk2Y1i
+VheqMNZCMTA5mWMSvpqyUMQ3bEVTdzurJIYs4LC9K65Q0TtDkFq+W6iNqNdcDLd
zASte3XYzRsqypB2FIM5F+uZNlkeewcKlfrtBo1k1soiaPkRvNjwGdiWxbiBkQUL
6wAFzPrXf5AjIMayJFS/fCo6mPTBJByq4j3swSAwBOwxmYfIga6Fy6DjCv87UD74
NdW6e04x+HfzJCVYqgaUEQOGnDk/xFRgY/YTSOVr6lryXGql9doxCSiTz7KqCg0m
lj21SYc5Sp+gexUYAbTX+4a3I7GKEtz5H557zywVxFDhM+twwQkE88bBLVZsqx6Z
YJh2IqIGa9u+Z1UIPrUDyf8FB+OqNg50AhWErkjsrOtGEPLkTOZPdh0oq+jDCPuX
RLFaZj7WVub98Ak3PkTMFNpqs/nh00W4DvuuRKeRz40DS8WR6W4IPjE1xynnHjJz
VWOmeGjB9LtkS5m0BQmcR+9fJOOphi4Kx5p8mXse9zYWI0p5VTMMBF0ZPZIZe6zJ
nzevWa1clQn+Z4pILOdcLHE60ziNTn0KfdLkA9mNJa8R5LuPA/6uPve2vvPxJ7+h
1SXhS1Ui6mY9jPADKkfjREdA1blRmTPu1bsMxLX+4ieujRJGfLsNidsPWjPc4rip
Q8XzCOyS1hW2NFx9bbzYJhZ6UQaJIUcP+UNMZ+RFnMYDezvTLnBSt528mbxiP/YS
PrbUAOP/amNpTsfb75397Q+q6dWNjG6pQWHVwisZwCxgDubWlQceIErYfMGMkLWw
jleFJDmMVw3M1U/OUOdvZnjVrK2oyp1HO8Z7fwJ3hHwrf88XQNfdKC+TJwHXb/ob
TuYMSdLM9LAojAZEN8ReLY05dipSpV1sFOUpMW6AivRNWozXUje23ZwOC80oslFF
BKRUaztDkDsNFINfKx7R9clnIZqV5yp+l6J4tqc1RNUN+dCZKAv/DyOizZhkJuvl
rL00OpnSqfMhq5kwBIwXdUwF4gXi2uRS7+fovAmW0qJr3P4F9ZTJrfQEba7nb1qS
3eBUOjh67MWDwuNbyFT4sMro7zHGi2ogn/LDmT9o3EuViUo3VzKX15DDrlPhhkfh
vzD5vMNLTZwIEO//ZNSwiFrYfOEuTNC8qVBxNXyF/bmmAQijqzHPQ8Zn3f9HtoRa
/Dv8WuW/nq3FQOrv3galyKq1UFTZnazDENy5b+dJTaK5mJk4P/DurQh3kUl0YQ7G
AzuCIMHalXIHZ4++Fq//r0qnPFF2TWif+Z0ZFSIeqN/jhGUdLH/7k93zSxkDlMnd
otCBm54tvuPQSEM6Ny43CRFNp7tDM9EwqDDjmOyKf1/027dpzVIY98mnSAEr1/wQ
QXMErHwVhhK+Uy5Ctsm9CZ5JPrzwpkjah6mgxt6v0qvtsddDEb2zc9iVMHuElAWv
z53+UMBw9J0m53Qh9CBldeEYj8hU2p98nxR2oG/GnmlPCee2BnC5Q46KSDsBDEwV
zCzYnaLf3HiCjLyZRohfTzBMycIgc9UpiW7cuXF6iwjLl6jHhmujUHJxqbES/7YO
jEY3DCkdJJJIq2siPbQBxArO2v5NINeQTJh2hNyc8uZq7oIDQl40NCZEiH/+s89N
cDhF+Ztyeks4BAxC+37uQsQ5o46GmPOtedMRDcHITRg8dsKGrYkr6CYR03CPbqPD
/tgndeIuyXbwxQO8i3XcQD2TLEIlFwbR7I5VYOMx+0YvCB3l0/netCTcG0qKylv5
8hojx4NHguhPSVnPWUMIdr32Me+tYPrXLEvS5m51Bfais5gR9+Q/epNGYQGsR7u1
FZOrfJf/HQHO8ZqU4SnC9WtgeUB44Ad91u11+O4DtYV+fAr6VnK+ugvKF0rOzpqX
dU1ZXprkIfDtR0u8YI08Q1QM/1fqS0nYvwMaGptrPIYhxz7sW3F7fgwkJLmAKLzU
RUmzf9DNSs4bbwr/Ygefjs96vB/4ROu+9cxQybwhw8bd/7xLH+d4HRApyFJ6K2A7
i539NU5t4qAYmEfxgd3I6ELFcOjNGj71sCj80g/X71ImmbabYTA3/EM8xif2tbfl
UKdkl720XEM4EUHBq+IwpRssgRMmaVwEqNecVa6NVa2ShXH9cMEqfDErY/O1+9K0
mle+TptHm30kwJimakeLbzHmRANcMe47VSTCsvsGYT3Nuuzz30XHs7hnmLXeksHI
nWQ5I0SRSaihjba+H8P/OkFIxJefNiv0VYNns2kCPBR+K2YLDUfWxF0EB+AJcw3B
uqSHz4BQJoSVuOqLpFn9S9rvjJkj5mju77BMveQKO4zDrewObQc6jPHchEGCOiOP
fXj/oYN4BknH2gPxER5aeFvc6Ctm7RBC5i9oY6F0BKPLkGPMF32LZqI86w72C0nl
w58OCb5PmMs38qI6XLYfP9jYDIqYX/tCY0jtHn38l5sEWAaUErnbxRyk0RusohQv
oHbACsEx53lFeZ2U+44kvP0TtXJScllSv5g17390OLfRUpMyRLFCqyCcBkQzz6BX
gJLlhkkuuKYu7tkYWC5JlPXdClE2gktipe82OUV9XdvadoAm2GUH4Wxkgl0dO6u/
+LEnVUFR7gCKItlPmcard0IhO+gfmUWdE8zPT7Mu/2gcMGWOue1v5gWqKNqXKhU0
lj8RB40P73103KQBPx92bAkrd3uhQtsibgwHU2Moaax9KdocBscxY70QlSIq5BhU
2Gp41KjoFYPIB+SV+CZ1BG4GdR+dhla5loNmfz6EswjcCoQpnttOcgObP2rozDo6
+TTilZRb09ykr7+B7nqgQXxWgksf6bWaFDq+jKqWlHYhky3pJQwOwnOuqboVZEUr
Onl1tv9vrgIx0+WIawMhV5ff6SmqAlOk1m1IP4OaWqxfAPT8gyloH7bFpE8cSv7Z
uB7SUO7Rs2dctUh1tNbTCT/Cn+U598kbuxSrztCgiHkPXZW990SSqWK7amlQWdpq
I37oniNI5hNkCfrgzW/eCAcyLF4DgYER7lxODuxEX68VaX1NSBIYH2Jc4lQ4wUdb
XnC8zvA4fqEAWhJmQXtLYnBTpBn7SanuUBC49eEWg9aZ4yaLBEnMnA5GnibJ1Hhx
JKok9GWvIhqFw2hm0vXbZEGNaCLE5LCmnRy/FMRXb8aV9rLLh7cUe7hehB514GxV
j+20v9mOmwVQMuRZI8gXT6SPkultJ4pWtHPh8fYLNhpHinURnTusD4WlASLabN3V
mifuEaKO1v1XpUQNj6hBgdRAzt7+NWQwwP2oMYxWnr+zOIGQ8t59XkPs6TA3X2mO
b+b5wr///eLpzZoos4jM6bBGv3pEd00O5E6HhDoVR4rZBjQtCkGicQDFfYI+ckKY
ftQ3+FgiTHdjTnKJqRPVfrOmvwJFWvq9G5RYC7szt0i8OO/edL2MeS4M3VgTxafp
gpteNZLtGOdYuJqgkk+pbYvmjBygneEivQFKZC++zZNXS07TgyHEdlj8bqB9bOUG
7nTqn5HXiMEjJd4KEqIzyHajmkgjADnh8Q5lWIzbiuwDFXRGnzmeK5xA6HLAJ1jC
Lq/eCjh4tVrzDw3xrIdhnbI1z3W8xv5jcZIHIP9tXdgUQajGX7EgjeEQicK+YlDR
8cMzwcJZKhhijGQ8BCJOL5xTCwCSmbBpWl2hSUbtFz1b/71y2QWv3DfqKyaTd5XS
vVwoPyA6V8YLEHwDJa3Jkxd7eJEFJzoz7yQbOd4SRfZzrqh5HWXEkPnc439JSuRK
j//5GTBdAQVUsQGGnO8SGUv3qX77K2TDOb3LJ1v+ud0S+J6GD6+f1N8OK3ifEx/A
onlTbtt8BAfd5+yPHr5ZuChKBsJoTl6IXoJiCMfOmwmSs6WHxaZwBylXqlVd7ypl
Z73pW1rji/FK9SJwJtpDckR/uCzYOsZgLfO8iEGOsjsuj8lW2DcnTZ7oh9xdP3/t
vMT/tzRJ/hrVS7iAVJF9zu4tQy0mOjnpzY/tA6MjWH/HAiXlYJb/mwxYAoHxyPYX
YVSCZZJH11SWDMG9hu747fDJ0ETCUrSnsEPW2Z507G+eYJOLW89W4dKxNr178r9s
/gVvm8djSW8kiJR5fZfW8aKAy2THTxgB7QckdYcmdC3spmpx2RDkvJeHZ3Z3XogS
lEdVuF1g5rILBI13Ne/BEH3pSwDfZQETPInKpyK6UdzADQBpNAh28sIvTiA631Ru
zXvKvPyLUXGddwDDBujGPoV9cRtbv55emw6JT67LmcLNzUBEr88nMt9g+jauY59J
A6oeFK2zjAlVFqFzVmVnPErsrnHiN6gnVSa+pBPuO0bHPMCK9r2Rx1NgK1/9UStH
4LbNOe8pxInMBxFt6nf0jKTitTwJ+0j1HAXSmO/P10T8YeHrFVwv6wT6EG26epsw
w+Sogw9qFO/lujg3T5JQhfQfCQ8mvvUpMs3jAzzRfklq/l8ncYScBqVDl0rOsFAW
978wJzOvo2EW9ai3Qi6JCivY+lEd4BftJ5J8BMgMfn7RccHYOZeyFBeab1prJkYv
GPVKutjq8z4NlluCMmQQXxG7ssnPeBhuxOW3DW67eHsbLb4xaAygXIk1M84/hgCK
7BqLN3MfzuYr7cBWX4aF1gvB2p27TR8oIplXMXhn3TzDACc8NvKk1XgqYjx0/pOq
BD+qnyjS3L2kYM18MRzthtiFAkvY+LY7EEDjepAbWBcC1rcp02ACbW0SFAdhF4Wm
uEKhJvKBiuP6Km1/REKK+8yGEvFJdnXws3j3PLnIfZkOwWy3psarh8LGPJSbxx1Q
/lsry2tmcrgc9RKw4raeg7NiI8ayhOkEfIzkmZQIix0VzFYcIsmnTVSydQuUfASX
Q2koPvST9wLAV0Mk/4FK/gceXCvM0XgjsXn6/fjxLzLozJt+qXT7RImkfaAdAACW
fujikMvZxJUGr5fQ8klOVaAHRK40uqsDH9ZL4RDcIcGqnfc63hpd7aJoyU8nsvEp
Z5Rf6GxNf92FYlZIt6iUKFWL8ynNyPImF1FM+W6r0AtpNoXQrcoRScaxbRVWEj6L
17jt/WowPOclvEsmIDThQQskxxq3wo0ll4w49/LoFBFBFKPCaf+Fh5/bDX3XOuGQ
2PTyCypao4fEdBxcc5kOSA7Y+IPQQWMFs4GFnPs54Z9UaORa4o7AwVjOFx5A5rTy
AbAWsYfsBWCAWzzjR+IZzfIUPx0IpEHNdHnNIn32lM0Tj2m8R2GuS5jfLHcM0zjy
iZp8yxLfQb25qr0tiat02ck5LthwUj2HvogT8miuGVPjXYxgQAU5+NVNuy1pKo6z
UjFvac3dCZmcYZ+90zOZw1Yh+K1aa1dED8clhaZWJYS0W4LL4vulfk1N38Y2xakD
lNXntVjqKS3Z+Sioj4iE4WNI1fA4vDRv3K+J1CbipP2P7Qmy/8AmWv6HHh8aYxjl
g/pwkaoWaXv+P1zaQVi1w36PvOyOjGB3x+DSQ0mNt1XN0UID4R4w2EwPSZAOwwFr
6SF4ycphmMruwfoatFi1aOronnR1FG6q/m9KykA4rFnDFJAxOJ7S7RcZdXwrsdKg
R3jdQiBMpLm9HV1FzbWBABPCdbn6tbHnMQ2l/F/R5nRXWhIwRN0+yrQhs1tn6E+7
ZjWlD3z2+hSJVFC+krg1QA3rHERegqeeejED1kHPV7aoCRuhJ8CQA78f+xO5qwKO
Q+En/JwtAveC/Xje+UxmNIRP5lO1z1mBCcswFlZ8fqLvxRAUOj2hYTd+yGWUEn4G
UDkTxNCozU3LC0GsigA/FGdL1yE8eAXSiKzjywZXujT0bMXn3g5g9e1FAK3kEBWA
BtoDHvB8GrVp0Hq7NtG2EN76gTJI6b5q6stBQOTPwXO8pHvq8mtxnPOOWYkAHtTE
n49OWN7E3Z2hmmiUaFbKcri+lqzov/Nzzof7hwQHovL0UFCLpWsejdRpXBSWxRdg
fjskJRuRXEj7ZdsRdGIw9irxgVhSQm3HlDvd+ZGI8EQmG1ivbB9d0ETlD4hb2bBw
PJfO9z2iDGlzwHLGkpPBHrok3clFYnr1jkU649dMccK54bV8x/n36YU5+EG4EbPe
iNZ2j1CLZ6y+XkAlPVXAvNPzGVPyk1VLmlDrZWDaQVsisY+IvPw7FqtZBM6tG4X/
ksJ9x3F25V+veXYpC+CrWR0VLq9RuZLQplpVNBJsfDGriVZCO0WyOwH3LCCQRrEZ
D6zHFabZr+i1A2gmVdGaObJNhjguoBFFKbUhnuEWb1ImPPop2s7+t9WSVzazL+xa
H41Ajb4s/JH1M6sKK8U0aHhf3w8p/vbxldn77H9PziOHJYX+Ssi4+0FjmLPBSiUT
KeA/Rtq92LEyJTHc38/lNlN4UJ3P49Gg1emxicf7j5t+7pa90naTrX7zxEupmjq4
lwxfOxWobS1OdpKV65u+WEp0OlxQBFXkiZOYFWuSJQkDD8/bSqGwiORizIfeNXwC
DOvAtXCbLWxnWV3v5S20Tn20tdzVc/4943DnXG5RmaPBP7/CPXO109uPIU4a1PXl
E2cV36n8ymsaz02LORdmIcGkwv0AoVKJZ1/Qjh4N2UCTptfQjVx1AMExbQSEP+qB
nW6Bir5+bTkz4hLDapKgg13Rwe0/vNbDwIaGFvryzT3WeJmW1cE4vgobL59S0e2+
FaX91i4xlDbmURi6WVegk5sNuBuAlLULUkdtvf2gDalP9EnhqDn+cOgsPQtaOh6z
Uyx3UW/T3pxL8DAc5XWQ+gsGJMtoyhQf8h4sdZVRcigmyjbONISM4ABIjQ1RlCrR
WXgu8MKW3VkKm8vJKbiKvqFRJ6cIQlloB4l+Yhh1/ZEr6itYkLKtAq3F3mAf8Ssc
eXPbFuINmlOarE7tzNMK+Hn3L6OC37E+TkGVMG4PRpPYdWSiFkg5l0rLm0bhc+6Y
vfXScBgoC0nKQ1u48z4IJQwTbyYsHmQ/mSqnjoRHI/Pzik029CwbjTDK/jVqqe/A
20g222BoC0LvNeuRd8ThVDJTx7d+nX4dcLaxDp5MCbrAWfVwXmTnBFkCw1jaQ/d4
kmyCT/3BzqjitrRlCVTNcABBVLFeupjuLAW4fMB+Sb9f2RxO9fVYe9iEckyf/bO3
qCSZGgrmdvW94x9PiiMjK0YIq6NYsu5QiyKuVxbt9lr8/koPqreUtt/WraA8JjIy
6w4GggYsNTF2bheoUzyzekQ9kNBl7P23mEuqVra3BE8ZM4738iB+qE9gQL8VfewV
PxBGMRocg9iGFvhjgIWNe2pIXmkO3Cr54g9jWnAj5mpPxKtYDc7oQIYfIYEhx/EJ
hjIf/NUKOZaJfuxPz1/KPtBgg7iVWy2XU6AOiP/f9rrQA7A3ucNw4BGDvi76z+Hk
pCiH0zbuNs79cXn/7Ts67efWp3upvSPPADlu2qFV4P0Xt0L6BVkchgz2xRzaGZqm
fFRMProO3ANBJu2ijWCG3QbG0rRXDKkz5s/kcx1Ux4W/K4+uJfu986ba8XVVSkq4
vsFnuVAyvqwCqGFJjNH4B0KNx5Te6wgEsHa9BalXTZ2HjFLkeSgAtXL/62CEzRnk
42DxR2nf8g/leIpJDM1amLo9YRrQxC8SCp13rlaGeT+BzGfI+z4NWlZVy8fcKZXn
A1DHK89q7VuQn2BXiyFPoH6RaxYZEBxyjxDD+suaN2xgb4FNpAX81p46i1GZSJPH
qQkEDyiFc+N0IYPbI/a86RyUna9oV7bHn0Y/98JN19drxCQ7KaRbmUz9ER5WQc10
5EeaF0ohdQTpY0qFcLw+OHdaoyte33bW8Jt4u0eKcEkkJsTIDX8hSp6ShkGVSSRr
ZR2viRPktpJxg7B8FILFIIA9KQrPn27cS62Uhl3X15G6JMweRzxaRe/haFB1FwnT
L19PW0Lw/7PNSRSwhSsaY5+i9lVCxqmGlejO9TqrifpeqKGSvJgLlVfwkCyAUn9R
GRdHS7g/pOJfd4JRZuo1m/2iHCdEti7pySPtXGe3kT4YA/fp/nmYGtdrZCcDQA+a
BjiBwN20auYMG6XxmuyPK1QYLv5HQEkXeLfDI5DytGrDVwq29X50vXlkpfxGEnLP
2X+GerHtYZrPSGwlyJ6t6kC7eJaTtTqNIGmtCCnh/UdDgAbftgINfODsbhBTzo6o
pEFwOERfnAjXWCtuNJ5wZd4RknPgVHHFByyUlz3YHgVu4J8Imq3tnXDBRvrbSs9R
zPvp6Uybg7EMJnSi0a1TzS9tl+HyM2gB/f7KGuxLtvo/jAlSw16S9d8hIoycYlp2
c+ErEMmekVmO8iTTbyGLDi8VLRtHycvlPqKiCm+EOgq12iIOzrXS/UFkCkzQytHQ
JiMtnelmfM7OM41wgrt5xcgOnYiQA44vO+UIHyrZiKYMhNRZr8gBOQpW3YjZP6Uh
u8WLyz3T7/PGoM/VyV/XCOzrNlFQ46niHS2PmFG7jqdv8hRrVv+ETowi95XETUYG
fE2FMJ6KVOYiEr0/Ie8cwxxl/zf4czIiMkrPNa5W7mfXvMZEhilaUY/fv4kcX0qz
jLi2XJ/IRM1n7DihDbOk3MXh0fl632LkTctdluVSUjn0C0ykfJgIeHWM0BR8qfIq
o32Nn934oU0wnVJPjB2A9ULz3kZWVCyse/asEZseTKbvfoZGzzy9KQFkARr5W+tX
18YwACQwxNKorm9xd1gB0NG6w+3cq+qKRPN0PwhGT5fXgEI18u04RvRu9pjL3cLt
Q6MfOXuoQSGglYvuqaHLuGWB3X/HX5qsU4EdM/o3ryVizunW6dvgr9UPgKwqKFdB
o0ta2TOC0MXrXfQyZKmYEb+ZChH+yTb+aVWoCbIMo/Msz1omXQzAweAf8abDOn8Y
KgJN6/m4hNV1znyllkSaOO3g2chZmRCFtYxopRHN678hzH8tjNFPgkgG6a6xn66m
oV7iW/eVaEKWpZEHN67RIKy2uG/Enrkn+hPUKNFqM98uw3ciuXeckXEeD+Jr6gFm
hHNhXjhLS6Qb1NvpzhIuC6IgTrI2O07KKtS0KNqaw3BPY36KoF54ye2AOz0Ymanl
W24wjxvNcwl3Nz5X/yNRWVDzF2MJIWo2PDvig3gtEdBAzDTVjDbWXnsmlX5A+hEc
rheD46kSMeAKLs9/C50eFvFtSIQEfKv/xbzPRT04A2wrFjtcx2l47fobqvjBe1hR
wwg231hW+mN9rqQuYi2KOG/kZkTHn0lOI7XkNI/DdKOxO/qIL6ud/w+W34hxWixh
eTk8lMV6ERK3X4IaurTHMAqkPI2GjZKsctXBXO4BHU4eUanbTJpUWCq+rjh6o6nH
eWthTrVUdhqSWLMuLHODfhcCfiWelCqG60U4hDDaJ9p8Modo20KLtFqaZYSUU0SG
xKXZ3LqbntpoY1LkQaFi+XKK2CTUaJ5j9U2s28MrPRD1OgEkyiKxZVZfDVy9wEGh
GTtt7DYzxe2FICWjQUt6ixFuJ/dK7FLousf9FXGouK++rw042ZdLfOp1GD8zEFn+
Yh1oFwGB9LEGgVwFWyjYGxseHutovbaYfEgO1r3m2uyKXRc1pqvj5claPYl30XEF
M2YHbcQf9lD1b5E8PEUiS15pXdpXhUM0Gkmyyr8afnoGuVyapM4hpY4+Xmsi+HHD
QY/irXwtmYkq0nA+acPl+7evXTze2wFmS0xhhSbkAM7yXbgxMJTbe5t8RbYRQtBa
xVh0HJHDLgVpf/i8IJUXUIyEo1K0ScoggSuSy6I6PDuQymXwfvJuWEmNhCkIQia/
ygIwjwfZLyYsD8vN8+nbdq+E8YHDK50gtqR337C3ss4bxs+d9mXVQsHY2VU2QjEV
7Lr/nat4LP5EoNgkZ54TTtqqatEGUcIBZPyDslrbkd9TihBxj5fNCz2vhAKI2cPb
ZkfF05m40mOBqcTwj5J4e61ZUrVnodFg0casEHQKPhn4xKxDBxgv6+SctuN1pkoE
G9aNv7VpV+Ubn3Hkhd7QiC7f4XZ6Id2QplAdOOItyfQTsVckTs9q06FkOF03N5+t
EJ7PTjPebJA9mML4Mjzt8HLv9PxeCW24S9Sv+WYfboxN2Xw2WBTQdUUknc0r0Quo
0pbJIKe3w3TxJTpErVqoTXsxpSaF8jd0/7uxkcUAZHaF281qTulUZcG9a777IzE9
2NT6CTviTbLUcflhaGT+6ifdjPrU9rh6fUNYYhWPhZLlfAE3VmZ/9cLp0McXv1Un
UIwReF4Ajr95FrtPuNDYOcHjK+j1VZmiG6whchM5ZcMmxUUW8yjWQVtj3Cokej8j
jQ0V54MfgqUVMEWOT1WfBKDBhfPVpiAqtXyaWIVtiR3GKLe+6yREkfE4CXNYVfIX
6lJsmhSmgvbITkB6jrOXJoFzTqeFRUjDa4yYPXYUWT+Tvu/rRTCabvHROh1bP7Zi
UIZ9T4yP5W8N26YAKsDl5Pphr2VImiAaqJy2bGicFKv7r3YhXs+Gm1uEhbZWYNuM
zzL2MGhAORDJ+8F/pq4kIa7nsfsoX+b5PPCtWJo2lGRfO+RmJl+7Yax5pb2xZ9WP
48xKjzKCHpHZXyk0NISNaZ4JIWqZa1L0qMhcRbmBR+WLX0u3VIoi3jWqDOjma/10
eCJ7YKppnocyS/FnEFOH9FJswy4bK7FoOs5xfoL7EQfNGYajiAx8CYoYSheP7ap8
FJ34XZQdc8IeTqZ5Npu7ZiuyvuLzfEsr+5n9rlGKcGqngluu0vChcvAKN+qdAbT5
7DzCdqRVqP3WdihYxAg+5B/duisJRd7HbeYPCbGoOfSQ2vs3C3wBh0Vwoqpl9/zn
Vjtj/dKdV1sQe3EubMtkdMN0ONLtPSY0LS5/+EYemmRBpCoomWjUuJxz66X1KKf1
CprDPDxqPoQDbyP3MhmEN1fWaXVPAXkD2ns4PFcDWZU4BdHbaesmjgBDpNVJHDfc
IRlYJY49luCxjN9lLsGw9r8bSi6EpYGPY86lIMMKE1AO8/gOAT6ka7g8atopdrdb
d/mvYotBmpE0zoaMPxjkCx0yr3D/asIFMhXFKDQqv2dWTHhzqk/o4fCCn7BdTRZI
bvlel5Dza6SNXWtIsGkp6esLUJ26Buh//Dee1grl/Fq9UlOc4QIemSe0g+4wB6NF
jTrcymdUkSzMflwy3KPad8nQOlr05tdfhykMCmNOVxvST/sbGwIwltsVARe5+o6c
9lD2GPapSwKY7T0kgBnlvgEgriMK6VA22rIDJQhpZSRexuGYvuQHU+ThxgDcYPDh
LCn5As9767pwu20QMCzPTxdzMzU+KajCu4WK5xA8h8KR1dQVhgXx9uJLBr3MvXa/
fAKNNApdBzPYNvM1Li32jKr5bo3/64Vgk8f83Y4GS8dYpTAKfCknWLUNZZTbiJey
85Kg0BtiY/ZwUBpeAx1ZfocMZe9jvYQSCrooINEiz8y4S0FxZhuynW+T5PbxITBq
PclD1EslbmhqHPy9WUaPhV3A1vv8TQw7NGVvTadCNoKCmYCF8D+82oVLLuaMcn0Y
xgvemHKEEdTaN6mvhTtuLMnlUbibTeOFf6SbmlqSaGUeg9btkLXbsR5nf5sVPqEr
yoYCiWZ6+ZbS8V1ERuePv/blHlklMvjtvoCKn0BPZWEXhuWFzSqmkAlCLgkHYFNa
4YP7I3Klhm7gbbGUaVTrVNKZoi/SSflFfOFq/8rTG3KrfRfNapYnj9KVAa6OhNyz
yGqX25hivQwb5thqFlYi6wlBYx+Gh9Mv9RxS9Q4/OeQPVqVQ4OVAhbiQbhonYSC1
AEZ30OeIsSeCO8dxrZ5cddmpQuQ18Z5HBYuPjQFG+OrorAeozpwYqHxrx0zsDlAW
NJHAeODnbM09pP/oqvoi6e/Gg6AG+P467XmvlnUnjRivcaEmj5cQC2x4QDQfCfwx
pHT62LJ0jtnrD2OTUDcwA5PEgbF+YqucBg4yDXJN9aPDI+PBmApW6CJmshhy3wwa
37JR6YL8+eQQnu2Sssr6a8ibJtyVk7Vi8F0fhL8LraVrRWJXSbAuf4U5a3KIwg+d
JspQeAEQLNUoHI9fkDqQG6J8kDvs5EGoE7rKdpeBbdysvPNss6FBCSXbTDdYM55P
xdT+GmjBMU1S8Tm8by0HqNmL9v/ci8HTbgFzuQWvPc0PT5IALz3chVTKcTsrUwGI
765y2uGCYMft7vqJb2BDzoDf09FCvINPsH+k4gO3lUkwIavby6WuRaZRtdwzl4YP
qdyNP9IAZerkgiPAR9LhCRxieORMTAWM7RNcMrmlxkS54EnT7R9QF8IB8np1WcrX
tQHG+64Rmdcz7shZBK8biP6Skj0jPicIZ90MVQ1IYPPG95PadVtzqRnuKVdZ27Wn
R1IN/cFed2fN7RGnpDoqFQpPlugP9wYJ4hKCWYefGa4XEwHWelxtU/2Nl2WMFP7H
2J+3kQyUTvw5nWLlDZJ6Frtp+AyRJ3iW1Di8NcP6tw+1IIkaE9eggZHXe5wK0O/r
m6IgHdthyE2zlzTW2dW+Iq4+kBFDj70bPP7WaYunZ/tlAGTnfxri1iY1aABrt0nG
gIhqtFl4F+2nlPE5gE6+YX894KGJkLjvgwQ2/ZExY0JxeaYL1Jx9KFTj44Jur0yC
THFcEZBqDfiZLuUmBetpYAweA1H7KCmku1quPVf7j1CcyWV72u59HypTmTyk96qN
GZgsbEceZSLQOVa296dejUxMWcLbJqTf9JA/owgEdZh6kUE95wGyw9lBAf7aUbc9
uDKLMOFKSKz/e/CDezw/phqwZp+lSjEcJoS+k58jiXQzFR0Xs8N3oX5MiVeC+HmR
G67aQVx9F0Qgc++35qiQxakR1Zjwhuc+6ElbuphQmtyxusFxndPaI89BadPJ1QGL
HXpZfl5bfk1frr2DuDVcmHKD91PKvgeqWdBdbzJvgPT+swx2bLdOKbqS8nt39q6u
Co9nTjuitgQdwkdd8AUHyE49HHOtnnPB3jWUji8nTsf19Ch52PLy1y22NrI5iP4+
TAsHkUKWxvBfzPkydEqEkiErbEnope3XmdqW0zHeK/K6zZY8eGpgewjVwRGVROp4
su9qpnIBRG+cNA+YkYrPsMnXEdm8I+Ylbs/DhfGbR8Iao2u3vrHw3cnR5HGA6rCJ
636CyTRyHp+qIQZYnHrzLM6qKDUNPg6R18D5C78cH4J/k1bcF5e2tQz/sgkHLp81
DRaF6F47kWQBBm9iBWDR22Fo/LG2i6w3OxyDVA0cpPdNKbLR1bxCmwbuSclSTX4g
r6E4YxM84DwvrJLNc3eJJTt8bn0Keu1hFcAIO/kEGkBXR+kar5P9NhCmUEW9MdfL
UosG7OGPwKVZHWDoZI4AeKsoSySTPgBdyTQ6jLni+ekDGrtRUEkiDiiN0UjaZquZ
oK1QcvTUbfBOqLw/KHOaMkz5kL3mq5xytE+FmnpEGEGlm9bj5X7DpIpdoRzHjr0a
Pdqbtqc7+bYRiSOM9dNJoAQnp16x7WQYAqcQHTJlH0FDxXNpAKTZ92bFxJSC68MW
53ehe1mB4RXjitbhhsQUkAIp5TAroOHnkeCy5pCTEgmzzlr50394IIEu7jpxLTX6
L8NPAEmcJin3rlX0alQNP+jr8AjUU7c24HyxoN4Z34fT+JsgEG2Z3sCm3sptrnKD
Afa43C6YANUkSYCwPGig4iGZfKZnZhEeBf+5NrvfW3/FtQKUrqMgG3Y9IzIdhTOy
DNc0xi57APntoCzVn+PqCa4bDe+ciKFNkaKZGik+9Tr1tzTWcM6HkkP1lqX8J5Ku
LRZw+9D9OetWh/5jvgzDMvY45Y1nge4X+ISREL0Vegz7UyHE2LA5dTwEaFcwzeB5
ZOa91utOwU0GW747+UyuHl6oMzzSXt3RgAE0OUSTsIYJmXz4ugF+wKNCTIPAAlwa
dUrJ0doIz6no04tC2W7j27/dF8ukOLz4OkcYxXfUm/RAEMkKtcUrxfGLz0c7JeST
5BFVG8Gew5yz01QVtOdkl49DcHhgc9AfOlmqUtDZMJkrIOyVMQ7jgd7Y0cGcWKME
GA8qh/zNqq4ABkJLSbBG3C57rV1unktKgfQNY5SVI4H7UiCbjzHSFNSJ7+xburiU
3dFrjELfYkZ5uuRD2d3fFihPWF65mxvg9mVyGKLib5pDYS7Xt/IgAepbeYWfmfz/
sdBFKk0OCay1BJD3vezHSCTCKwyoVUQWXfbAr1PwJLda4Ftm2ZyrPx6hxmP5Hyx8
2/ClYiuE1Ad96OpPs6zHX06Idxswpdemf3Yw6UsuIvInlTH6DonFTEBVfLtxfY8m
bMAouaseZnuDgRDb9vcd6NKig1HlTQhVfoCxaFVaoddcPoI8yCwE6aInPcGFdQo1
9g/uvIOTNeRJKs8WLPVXvEHpPIYStD+bPqLvzXZrrkxt7Ae1LCR3W9wf1J30Ly9l
uJrJdJ01SIgnEo98WG8oI2gW0yS+OKeKITRzxU+J4/Od6n3ue4iJNRDMUdGWi9Xr
czOwXn9IYeh9y4Ktpo0OtYk8Cj5Hs/G1ly5v5H8nbJpeEALbsMHEJhEhQDbcMJNb
dIsYI1PiKhxcXz48lubMs+c0m+x3vCJ5DJwKw49EZ4lpjXLyxuHLEVqwUX08YO0O
b29Sl1KxLgD7yL///bX/SSxWJsGxt4FeOHttazE358/PkykLFJm8XTujcIOeRxaa
/yjTvTIjsfXIUNic9BLJ51h+cMv6uQOe0bZppQNi+4a5+9beIyt1IfPqkWujaLbC
w6TiI774PrSwWVu2sHWdrUQJdWLJ+W+gOhY0eiwbq5js1YujGIJfSspmvbqzs6zS
gvTIUhN0ghWdbYMHdRV1K913RGiv4EHzCYMH2e5VLwb1j7qiLiHbhFPbMXOn2oIX
Z0mi0lwoB5TBm6ZG91z+BE8kNGphKL4NUANKyGTdX2zAJIDyQOAdhnzDmiEhy15W
9RA4yOZ28zLOJAhAcqm7/tKLswXg6FfY19SAhrcw2Ek8jPUJ2o4d4Jfjry1M6hE2
Lg4uKngODhY558RWFCfE+KQ2ecncJ/dgFAqNJWoZG53jVHVnq/D5I+ez26o+hZxR
y7k/4X3RqnFWtdZ4sVbhlNEfgdhvTxi8pLZYMQSp3a+vOlLAhLBiDhu0xiIZI5wn
v+WIy2M8MEcSMSSpGYR9SjMKTC8D8I9FlzRcvWsbxjdaSv6B7oeQxvMh3zzAEBB4
G5IeKj3hH8+EfoKUY14GINoN/oKvWRF4TyCm17TR+gzQlt9XG5rR2aOAw+hUAq4m
S2wWf7rNw98nMS07vPsVsshHUS+iC75Boo7htAWxH6V+7gM6loC7w7GJBz2lPdzY
30R+nTQmuJGC3WfluSa8z2H/SLIcoEI7DZIuxSVtg6y5+N0BNpbruCKO1IZiqZ92
IpvQ7iazRLZC0MdYtVm9LhUGKImLaZhi8K6HNp4lGKwVRwH/f8RFHSvf76WmPB6a
dqrbXfrZ3mL8wZR7Y1O5JMs/myzOpERvZwZi/8TqFiF876OUTbRub1QmkBZzHh20
xjUmUPSDPMufbdPhDdiRW0uA0Ncd34e0GALOmWmI7HUhR5hNDv/UBlIs+Iwu8mrk
LHlOF9HauMRLwDF2kdYI3Ko+P8xeseKSwnVJXKMVkwEcVkZ+db0Hs0YJaaApENil
qkgVv2hpgmS5jn3/YCjSVMTtrPOESndpXK8jeCHRlXj3kOIUb45ZKsvFc1XGgrFj
HzW13ZjkNzCyEm1euRhcXsYBmNj00BgmQSO4hwe8mSG1gVL5QVyy95zeHXREgHHo
euxmiEcv2Opx/R2Sc+c/8iNnhEyaAoU6+At1vI1hazRZt8AxTFHRXWJ7UX1fRDxr
qbLIvGXCSFcpxBAR63GBxQs1T1MsOrjcw087uCrRxa6EiefYeZbqNZxeZWLw7vzE
oPnL3q0c9tdqay2hMX/XFDV/aIobzt1u0uv8coJxquYzjH8xlQv9bIfd/+aDPxZz
Mz3nUKTp2+AFNRQk2oV1ElbmilgkEAdF/QCaPY4ertkIXwv+8UpZy5nzfJ+esw9a
7sSI16VqkFcNl3f4jgcWApSVYLvDFLlSl7+fCAVdI0ELK1P6YJrfm8KBxlFRgg1t
VVVGw1TzLWhC8ZAuCqU4cigVzGLHGdzd4dvYR7LGssgwvJNIZTOPGiobKl3ieTDJ
A0GhBp8rM6Gg6GTzWIgUtR7sanGMSW3/WBySgNkOonwx71F1s1LGdXKW1+EMKIh0
LfuwKeK5rhusW5N6r8ygPOQyLiSZeSaofekQNNz63kBd6QFnnDFTywDm+DPeLe8r
Uj+0osAziB7NP4IBNgGQYb5Hn50gMj6yebCcZC+5+0aFpOHwnjIKuSDOyxn+m1Jl
YtOZmTmzbBYGUxhXm/FI/dmKKunoz8MPHfhHp2tD2Mi1Drh5Q25V+d//IaITUGnk
ALJA+CSh13OcEmjSD1VgS7YhHadd/e+OXXssfazeL4tVuM/UuAPGUvizcTha2gCF
F3zLdKvsenXHcYpUaO3OKxjmZBEIGO0mkd1rXpSOxaUgekxvgjdJGzw4yutlcYYP
R7T3Fgdd8HOkQx3th1vAl175tMhG0cTyCgfXrV6xeNvUaFes7K5fdgF7O2iGJ68B
qMjfo/fHn6h1Hp18i95xGPdb9gOkCB1Qnf/Xs+X2sLyP5Vm2gnIlI1F/yNuOvand
4zMsEGoPn7Wg0Q5LTWSLcIlkKLCJ58EqEBnXZG4Y6FAV9Vmp5eGoSvYoYMkz/F0T
a5hsdhqL3WQ6tPbwek7ooKIFHRK9bJHOczidst5+sL1MyWCqG7RYbu+43ubbU+w+
RILYo4d/3c9F6at1DR4r/LPC9E4nRxqcqXtthotoPdVdQ7KqJt5sVOLG0+VTDy4V
6PM55I7VXbMFCfq4QCCtGA2xA4B0mnX0UzOGqOK9QJi1pkyV7vYodSyyKNZBgAsz
j3MVzFyCGqsyPM5ETpkWCLv63qjsteZkPh2ISH44Ju1QlFEsvbOuylTD7tf/YBaj
YZvKxjYWyW7sznmESMbkZpwbgGErrxVwhkhpJuzchRBd+C6eUxEV9GtnhsMyGQ3v
EBiJ2EBDd86gir7Ox22r27UgtI+6ApmcqLAoa8yOeu459kvIo2tUZz8oZKDgQ1A2
K0X0bWVVPnhWAc18YZENEl+3aADvnHLpQVo9QBQAnOPwTxLR2MmyGGoqjNTz6EmC
yxUbEPzY6hk89M2NIPDx6SpgvSNR183Ra07M3/QmydsHpWododWEVrGfpDQdpcf7
KQqPZVZMZA+L0+zg82Bg6HZ3I4tNcIAi/xscln4ZMk5nwBs3AM8oAWqST/ZNArfg
lQxZIq7zVTsKX7afUYDACKoxWAUSOaAWnLZErnnWwSSlqhyzheIDetqkHwSrkp9c
mf+GV5aU6n7JuNRnZPcBJcdDL4gp/pZacxoj0tQKW9f8vQCk1JI/ga0KMOWc/fMG
dnBhh+Zn5ptqTBDgspn3g7ne2m+8k0EU9ulZXsviiLhSZltOe/IRlP0VgODBcJeZ
pSvCqtuJAFLvfpCEoCfguYU4UaH3Cl0qgLi5PTItRVBbvfpSlHkEjKg69SMezT3U
MGJIekhAe4y6ju3LSitsli2VmtuDP0VrHNedfADKXR90n7JdMkVhbCScPkx8lRas
F+tlcrLADNd07IaV38Fp40k4crdROIsjrAmCQTCP9r1G2QxlLa+6Wzw7fBrWmREQ
Dulo9o9/bJhu9Xb9sPgos54lAzcCN6MQKFF5TPWlsCGUdTlzq45r+HTt3GKLJoZZ
5lw8/7WvLtf8HfaX568ltdm4tGj/PyPtRoehkZgH+pg4Ar0w7vcnuss+cKfzxTvi
rirRpN4OI9nOBYCdsPRwzdspdXoEs9dT2//Msvy2JwN20PowwHKUb2vLBwAGXaUT
BdWRO2sTywBkHHZYhEQbbBr30Nk4a1cUr3TJjhcZ5HCucq7v7JBp3IUfUoJwYXPe
2Y516MkndTwrVUdet/Op/HTwunzwIxXj95/Ys6XAOrGrlKmY4ZAu9Tu04JW57seW
CWFZDplI0P3vXQoopX0A2eOsxQXxQiQHuTt6fw+QRhFYnlm/atnQSPBVq8AMwhBc
Bsru+akGIjcHWhhuJgDBAkeHfAxCq3Bo2YRVrgTgBJIP5e1Ds2YooBWp5VNIlvEL
AEtwpEIaVwK3XSD9jRkHV1PpzX5mlsLXZViwVmZHosUGGuJPDZhw/BE/odes1EyB
TbxVrSzMzVTs2zldb2eX0bnSGvefjbULZYKKXOMj5OKjCAyuCqJl7/sTKBZd/RLk
QnD+yWm647k+N2A7ZOMziHR/5wyIEE7uRQz02pz7LVnJ7xeI9mc1WTH6ZQDeOdgt
ve3vYQUMwbjGzXi2/3bBRelmap/5EA7/7ytOpg4m/OwGURnK/tDu7Nxx5Q5//KRV
5C/7rRS3y18N3NhVl3Y8on0Eo0JlIXWU/wznT+1SHmRVTGCk8rv7vySTOkpuv/iF
78LauLEg1wCmbNzhnUFTiLcYP6Ugi2zfiSyAc0ggV6vGXotzBS61qQmZIvxBx8/S
UzTxvIwp8esa1pF7F/Jks8v1MNlpYt/EwN5Zt6Icv0tGSZTTDxOshvVKK1/scm6J
d6jBeeYKEUgqkMG4RVVXJCUypXHwjnI61BFTWsolatJZrnHNX/8949GiCd4uhMuR
r2R6Xv4REK95h0645TLnGT0ldALwpcqh1cifmJ5WVISlu4loXvbQ2Mlz/tn+rOyk
TdJ3wg1XOR4TVZsqkCVleXsjccbWJk0PceATgMTxCGEclHEQtOnpvZ+A9XQd8cLO
l71VDwprY73WQhBgXl7ggdm1TKSuNa48eF+yNN2H1GX9PrlB6cmwtgRKBHPivQeP
xtd6ATY/tqa6XfW6HcGtmjbcd9kTimKRIkPqu+JhsOu0NlrogU/b8Gn/n2nnNsTU
ChbSxPzAbvHI8vknhpKJREysPViSseYzme5yrOO8CMk/o35WPBahvWyGGc9s3wla
QPYvgiPuZb5YLEVWW+5F5pvJkP68RDmiToWizDCPF+lu8xd0VhDXufmQEHbUu2q5
wnDhxxJcwZoqm6wmer+mGnAMJVZb+HhB2buhN9FLdyyjamC1uye8AfkrOyTCfAAn
766l0IMnj+2eda8zrQV88QSq68gNn/25aZQ1UkuwnihaCimG2+DNFqlrvgwSP5mX
ywNlKy+znbaJ0v7NJ/WrAj6vwGfaFqXs6CgG4BdIdT8VcqxhH9IZ3CgWEzcrTgzI
LJFjmgGJSIoJJ2Mx2JYgp/C1d9FD2iA6dehRSSU/vfUQ0A0Mpv4hi2pTAtX9AiUV
1tix+Gwd+sG5ZmWN0OUOiCx+WYNhjaozBi4JfO/YjzV+ZF6D1AhHPOmCBrZ1hc+5
Ws4BXh8KzZpZaT+viWQ6obfnEwuimn51QQGbCWOplqCbfdGEezurm71OKpcnBNAb
LGTc67wWKFKgH+MlcZQpjmI4BzdwzaU735SuWobHzVWBJER3XsWXV3a7xDs++O11
u+TnFQLJ1idD2Qgl73S65SGb4nu4OVfkzWZJlJLVm9qPg3oqs5L4vIAK3l0Vx6TE
EIQ0VGRLCxTRFpfBfmo12+zKUBF8DSb3hI9LHntl1d2v9WmZMUylpZnD4D36T6NF
gBu9iX5I0v2i8NBjNbiC9iCyj0aQfZhZVIsAkPtCTfUIP8aoDFZJcyD1vALCc1lW
wxmkK84iNPKlYwmuizpbdNIXBUZwTLsIb+FKwp7KK0dFohrLao2rByGL881uRXyr
xjowmA/L2eYdgh7hZPq87KKLPZs6+8f+4BUv9qubF9C77fjhD52nW7dD7BUe41vv
//x+lG+JPw7knZcPE84bgJ/e5vdx6Ef/J6xBzH85IK/UqpmtHezdnFYYclsSLYSY
ROKwGlhCCBFVmQMREq7aagnw43+DIuZvahqnUp5Q8etTdrBH3hjk0kRmPz+xUmQy
nmPIEI1EKJ44nACCNwPSu0EAVSKRYj761zVgKXW1PWfsMeO882uyayLNq6jTaeLw
uuBmMwrZWw4R54cW9lIiHtIAjLgTRAWheR+wD8wrjR/ddJ5glZaIZ4W3gf12gHSH
xS49CGY0k003osmY9LUw9Cla+VG/JZe6o4yIc4iePHPnsSK/ZlBETMZXkdK5G/ZD
C23UmDFYKa5CJc1hr3Q50OKGDXeQOGoAlE6tZQfn+P6/eeEdyCfqPjlhzS5c1jTO
TRgto7Au3Wwv1FymxCgDDpJh3dMAKSGIsNIGBXtwQDW2XNg+LVULOeP7aQcTyyAK
JwWfmRkiNZ3jz4QBudbfJ0wVW183elbM2KN5W3V3AWKCOluhjGROzTpY7Zg31Y5l
I9SxuRxeet18PCE/p4Lg5uwY19oNwhFt4SDPMcCKM8+2cXj4H2tk7GtRhEwKQ6Jb
k6upBsZeyEXj/mLqt321oDhVuNx193DVguhi+AZsoSs4BGD+wYIXzBt4f9SGAA+8
2FcWoTrt+8Sfgyb4Dz9aoyXCNxEbqQW8nZPwByzp45lGqeKdkoQIbUic9wzQf2Mg
NsK7NEXlGMgl9nWZvQZsT18WCyCmHQDdLSjQiR4SllyhEZdXd8j0NFbpDhv60fI4
BxDaK7FQSPtpbgykP2yNNE3x/x5afOy0WHGFunMIiNsu7zbh2HLpUNhG7lbY5yOU
fnQkzz4CDABeyE+cGg/+2q5jowlyJDixpma8JRevcezMBrHnVXqdP+6EzZdIyrhP
+uOf6z1KoB1WBe1zT97MF1SwoCrUG3l7mV8QCm/anWkeokZCQSTmHt2XJKX6Fqt1
/XxFtuc8lDUpHna3U6NKci901tBuOeH2mRHs9p//A2ljhtmofR8BkFTruqeYUFIL
OX3UFnLV9vyFg/gTohMxhfQCBO61gRKGsPiM2iYnrF6Z0tKkN/JojjJFezYr0VSx
kfwI3aUwXRfK+dbgU9Yj4iJm9wE5eVxwSYOHeyqm3WMA5QWVtuD86KSsg7DYYmt3
KN0zUS7HMzAC0RiA5QR81n/97fEBPPS++cDzh7Oa43zHXJoHlU86ix9Jw+DdogQk
fw8AdFCF60v3bdSFjbtdh4GOJmdC2JNTFncp2oAfZtX/ZYTivwlwNSHgJ1DlSXDI
yXFZX1F9+dB3qUU1vN+hXunFjOrrZeczkIepOcz8Q6LxuH2v1wcfmD/yFgq2NL8C
fd6iuameUHdKlVfyYkY8Y8HOWWiXV1eWpxHMBZP8qvLkWHkJN5dbFbCLKc44+6Pr
CM4lySFiZKUZD3gkNL7ANuugj+PR3q28hNSQy9pnBiLBKzY7eRiu+IRBAMV9tRGo
C5fNhZkUeOLQ+Fpk4/YVkeVs6X9sIy/BjQZm3d1yVsjg0YfrPyqzEHfMwUIJqa23
JgU2Hd83RiyKUrYElQlDFyN5UjIRxx93gACFwGinMaCH5bvSBOA9BK1SvvVYk94f
TKpoQgf+OdZ40s9mReG0MAQUcZ5pcASvnLilLaBmvNdGfqc/MIh6yZEOfGeEnTfj
jtJaLFe3Bbg44ZZw5fy7FQzDcJVJLvGoJOH1mBjGclf2iETfGveMDPK5FpEtCv3A
KZmciKvJk+vTcBxL4KgaL9GhRZVSXXqlXD/tHRYewSfzTK7pyIdkePKAXsaN57HF
qeMuhHBztVr5cQ+wTO2LsQdmpTLxkDCjiIKeqU5Y2+FuGyrsD8JIQVE+8tB2fa0b
xkPEQnQg4MLlvSFxybV/5/EJp6ODvqo+CPspbOVDKB/t1b/8hGzz+mAUy2ewLmV7
bBiXN+9A67MTCbJ8eCFiO1a8W8ddrOoCE9nnjBPeB9IE46XNFps5ZrHdjMspZffU
UxyWT376xvCTMqee6TTOYkUkCaaJo5cv3SYyxLsY2MLJMCHfGV65bSqn/ipCAaWd
C6Ks9lm/HUukj26MV/YmSfdprsxbDrln9vVmoReyGCBtbHt/lw28pdL9f4BP6bwB
Lup7gBx9stnWyxa0VGd14l9phdfNng9jS/oGTbnDm/iSJJidBMXhNdANc9gQIpXM
SduAIMl/7PepVAeGetgoUJ5TuVea0RCxOSR1cUpgQlv6cRhsb4mvAVgYnlGtnhd1
nBPShAPVJ7hxqRL7p5BoIQC8xlAevt6uFwtzrMknhSjborjbR+FnL8xXvfa97KOQ
D7rGnuKc2Wa7yWqKQlnklNdgxiJU/S7H54NAQfX/AnF2Ymv3fXOFTldEp+z788b8
TI581JfdZLCkBR4IL4P07OsXc6PTUvC38OrqbJgbF78viQl2XlEuU/r7od/zX/ZF
vxtA/Ir4yBd+l6fJf/8MCTeDC9bdm9ytuPDw29sS0r+eQJCt+OsBwTYd9XZTpXtT
+t8BljK+B5NWnO5sWh0eBBdmMe511ez/WFe71AHNrRj8Xjockzpigu7EeeZ418c2
jnnr/xUIuxla1TmHnD/gNG89tYxCcHLiIxtBEY44bcTyY1vWmEbFnVsLVAlxVabd
Q5eYsY9w7+032K073u3Xyu5NwK+01aYIMo70BbaZ6xW0MKVg5cJ+CWf2g+Z/SOem
CHuIgdjAYnpZW6866SrK19hmlXF+dv1EGL+Ht0cz+FtAx3WTSJ8A+RVx4YhAjuIW
x2rwvO6V5y47wamzbS8IF1byy8n4ZmBV0X0RA0RRe8FBl409k+jhslQNtKZwp2ug
0S2cHV3YoTsyucHxpisqCabrD2foMTaCtzIuofjQ6MCOYQ6ikaxCVGMxmXFomnj0
sKvTzJhHVP9187TnpRMJfDW0b/a33QvTlo09fQwpEDWyglDP/YSH/p7G7FtTjpjL
oCZx0JicLhXJajLFoJ2s2OX85mGNmsNVdCvWbO+VnTZETK7mFfRCYr8Ktf3GuS/v
Gy7nuSvUzs3URtKetNJJUTb/d3nzCJtUO6P86cQ082xREbEQgnoJkUO/+CED5d6b
DfnsW4M3wL0QAtO4AxTjS+KneoF0sJNqXGsS86VZJrZQRmtj4NS4N92z4dpNl1f3
O2FJYEdARWp5GecgaI2g/1mGViE+9CFgmtoYOIaf3VYmbJrY2pMgH8wSB0irDZ2T
lXsQ5+SiiHXXqnWPrTwMXkd/az2ux4GnrN2JXGEOgHRdv/WvqfjDF7FJbf3qNy1H
CugJXpGBfK9a7ZP4R8ktJ/TjaT9S9j5WOp2vGCo1ggHuHnowjr3WSlTj5VCAsh5R
7UQUbvfZukfjwylBcNTm7vSBrB5KGPdprb2rCyYw/wQu/ZSJkM16uX8uwrEEiPnc
NQjpO00ow374+ak5N0c8ZRXN9vlUO37pjhefZXG0h7jG8eIhJXjXtNw1AcyTQJG+
WX7qmgwIi8RnVyqwuMqody0O0rz26SB+Qt3TTtmmI0qcURcKKEhrNa1orGLDV3+Z
nobvZqMkbYQDS8Pb1HBWKvqmFJll9dKljOVdz3oB7TgTCtMDfFPR98jwnE+ppadP
pLXlHNDKfbN1aNej5+Gx/Rs5s664vxZ+vmVzg80/y4Q0o2c4fqLhWjgc8CSD0FoP
fYQSfp1L7GHyOnL7swCSUpKfwiLrNpQVjdLHNdNpRwSANmxDl8zTjFf1f8/SMfY8
AJqYgiRSj8L00nb0zyTOVmc7kmsyKyweWo1OvU+7/2ZuLsTPKuIiTGajnGmvIRl0
czSMKLGiHV88kmpp5x88ZQnmJllIfHEEKUhcHqLkuu9DchE+u3ZhDJCCcqwidqbR
lzkd0XjCgHD1XXjb79D3J+76GLQ/sB0n5mRRP4zcm/8SiY3jPrRVPaXRy3LJCui0
Qfv9JkoPROJ3GXyt6uKA+nyj/DWyOlwri0w96uAmCoWMFvPy8eoX1Cu2mSj1iUB5
lyAKfkcgb4gcP4J4Pj9XnmOHooMeM/UucAIcYQu5a5pi3OsXwm6Mt3gYxV/p6RQN
D3eRwSOYaCxagPZcHWWU+6OX1dhPuh/jaAhpnh3ZYJjGWcBd0TMSFnlqb5POvfV5
3driW94YniJjiQgZxhcp7UZVId4q/khEp84NLf/WEP25yVO4bCbJiIov0WX356ql
J47Qwj55TDFcQ+CcOYdjrur67Iegaq7LQnb+SC1VyN4u6f2gNaVOpxATPa4Gav/Y
gPu2mILbUfjNPed7RS4Ve+Pg4Xh1j4NTPhFrKAAgEBDQvFEUwXrEyTMeYxVRAYYC
5HWgvcszOqwJCq9fcBWfBi/HOxtr3Z4D1kaaMR/JUvgj3kdYzQPFQqXAtJmcWGSf
hiGXAyXNM7351VFfEzqBP21cc5wtDu/JAxY0rAREFBgopvAOIaaIDNsk7+3JzESe
SZnbL9s4RsGxnugARqEgc/s65vrvFjnyQn+GWI1VW0LOtW9t1ndFLutRiFh+WSSe
X/HL2UreEz24XPwNNCU+iNNJdmYVLuec75b786aPR4/m9ZMYsbeHKzsY/I+y2E3Q
JSbRPiak3PHhXtTs/5nTx+8WzLHAm2bno+iFYTAM1pnj038l5ylzhUX1uxnPJFw1
5qRhmRuSGGeORjaAV9XU8ADOKa0zrwc9bwUyqIxvrnYrzQ8hG4tSh09vKHfxZy/Q
MWZ8V+M4ynpaEzEck09LN6xPW+0qmhQWFQTtjlM48tPPRzxPIklKE0CMktZTZs0g
wTYuIFBf3cGigk4mpxLTk4EOKgzo/rDitWQQ8MpRfsKyJrQ+2IDueipfBNwYMatV
tgJZ4gynBcM1EPrk/sGzExH/mghfoGoaG0WqzDmblBofQpXSBVREgh9QetDh9/zO
RbOwNvsIphO6B/TKBk+tmJXyvJ6g0g86CmAmLmb6+m1gfDQel9RvS2RJ5it7fJEo
mmFnBIUvEDV2ihM3E6qVVanA5+nL4eKjx6F+BMycNS8E876+8joqxKzno6Nk+Cla
h9mKzWn/F3Yf8zlcyJ9Wwj7wyx/KhqGPut3utYBr9HIbspixLs1W9zC1sZy4qcLZ
ek1V0T5mDuvyNl6X5cCacJ+ZfB9cHvV3GscdGekWEZgn4NRAXEof4EYrqRytIJ4v
FbkPQthpT9v7r9SYJ2NDYBcUJHH2CnHePy9XcbhqnL8HWPCNsa6gnG8CUSp/X7Zg
D/CVcXWLLoHVRf4HYf+s/KDaxVGdXlaaOj8V8IXIyv7G/phDiXJZNl2PMiGBuUb0
Cbl4oQ1Uj42Q2TKlB+yYkYoKoH78AUF5/Kmwkg1vs4hAD00aXwrvgniJSeVS0BRc
tx78j52hIFPCY6sNe/t17gX3ifqaDD1Ox0rz8ouyTqSXtFCKY94D7l8WpxRvBsKT
ST3P++aFUkUe6kpoQVUNpeOe2e5g7lvwZJNqbm3BHZ+oBTXJpWQISwK007GQSAaH
K6nCNAuQcoj5qpvBgKHFPRwU8g65FhH5pNnWI5U5gOv3SGGRSxF3wmHF6nVMUPdw
0zqiIAsXTO34yXThglu/9F3pIsS8SMndg65ks8Jq91hQzqMNpKsNIG3xZ7OGOBiW
3Qp1pi1kM0ypSo8cSdCe2tarCiZE1AoaIHAtFVqOVB4qYcnQ+cD6Ln9PobDc1CvC
TcPzCaQ+MjeHAc2WCgnCyXqVyKpZV9L3tMGEa/pmXQ1SrfCOiSN5GAe+eeEFNSn+
HPqjYNkRp2B+owpAMNd/pK6s7N5Hf8lcYjPRyeQQGwrOve7UrAbyhuivPxUS6L6O
Ml5wjY7r/gKlU0A9Vdpa82NaY20ZSL0DXxlVmkQWIofoc+NutwTu2qbkiUUhRFq5
Hpc8IgmLiPMFLviUUMayvTIzS5iTi0K6NpaUDkmUBhAdKr1bRyYfNOj3SIp2JJfe
2fCEmMu+KHtWvygG7zyVX24U5OJZ+cEKaka7nk5ReHLgYmVqzTkdEORS1oDXF409
ysGPJbvadqIQAGrA8RBPBk+bT/sGJFGwZHdcY/A3zot6bwbtmq8+J+nSIcwBTtA+
E2ghTNVrWm8EgDFZu3dGJjPZjwbAP1H0xXweWqDB1xsgjanfd8A5Fi1ThWK+D+o5
q/kWTK93qdjVQKs+YxbNiyn1xbGPJRkp2AjROBnXYIjpO7Om+FHQTuP+lc3eNQEM
BKGwQw37Y98kw8OLSp9FP8UcSLmnjhePX8tZ/M0J1bIDkoDMJs27e6ha4Y4DEmaB
7o1Thga8/eoroSjUssJ03TgQK4e32HQOp+1nuNgfeddR0xjtyPkPyxmyDhPv1lu1
++naehjq1/OZJPrM8jaslUGyJHJKeHxzaAKyLlp+SeIllzV1EyqKCvAD/Bfsz3n/
y1GjvHUpC9AKsX1amZfeam0C+cgghi+Vi9+sF+oIPtjtnTvAUYi23USe4rmFLxv1
TBxilEvFQXaN+WGJfpkUV32vBfVU1Cd59tq8A5MAMr25ZMvZaXfzEeFaFyiAFReC
J8z9iDJzquG/0yKn4Bb6vY9UMTWVqlw49wP27bwHmd6hC2eHqljdP3ryFzJrWl5X
gAtK+IL+5FcyuwfJJJB0Bodpzz9OD4ALCM9VzC3Jx8lueBYVGgIzFKGAVhM3BQYS
ovtGD4qqmMfYjwuhv21uwMYyfSdWktK9Z4lR4lMeOM+j9RFjWL7dDTUd237JE7NK
UwAlDzvw9JiehLfv0RGnYtpoKmRjYYCfFQ/Svjf4gldwqescukz/Cd7dumq06nvT
alGHngQ/pFe0oABXui/RLrGpCmYzOcclagxb/DpHt/fRaUfR9vMKD9OPAbVpdfMX
a8P7/MFomfJ7CDwhWUF1LRNJJCNvDUKPbsO1HsU3V5M9EO3BcyHVnV337AhQuIuB
1VibvXtdwT2A4ewdgHNPnU2h2fcz3gX4qv2ZK7iRRPXfXuyZWbfjHpl7e5/Bzas4
/sQmSxdpO5XMqU9wfFVIghXqeoczrcmiY6tFoVJWbAdNb/5Ij3FiDVapa3Jx2zgF
5gkASRAUiqwMYsdSOXPqoj+ZlGM2O7jzsuY+avWef8YJ2lqOSkKzMeX2XwBqCwW2
cRDWamkqi+VRc8SgQiMnn7I0TlOCzEl5XNTdw3agzHh1NvMiJ2BcDWYRuBVwsKTm
zVkJTKlJh0kMld2CuhGYJ09ydd0kZ+Qh4e0oZnKfFYgDjayCyixUF+XLhcd+ECdn
NqfsNId2o1JAHRTCRNqzqiploG+D8/idapwPn54tYZhmUIDy5atNXumRcIJNB3Kv
zl80PzmbTo5It1b5p4TIWbGytEng+ylJpM59FrVlcAN3V5fHqPWD76o2POgUGLhn
XeeSPPdFEumO1kYTdtA7KDA9IhivuCioO02KZD/mGKvmnv03Z2bnDgNnAkG4OI8N
lbihoAsMQsLt1b5KFM4D/b085WdAOYzm/NS6BT27xc3Daj9irFCEzmzFvj0GvF9V
uzuqycwYeuwkso6gb8NDqa9e5SGZ0jguOJqeJGxwbgtMiRBYiaydeoZtRCm5Gai0
NU8q6d8YDD7dUaFJvlsuJ1Cv7XA/fh+eQdIQ4SpZFUDvRcdukEAVPNSPXFlkHK8q
LYSDMlqoDzO4455l/hm797+shZS7CsUp+w7kP/LKkGNwPUEe3QLZTs9m2fa4NDf9
WLRkTrE4ik+ajwlToWPvoFOxF+k2pRVj4m8s4bD+D91rlg7F9luWLqerrkRXxtyO
/YYUs38WIlGn3I5iwfq61Cz8gxKmMu9tXxP+zZ6p/dz3Acj5gaHWyHXnEqalmlXX
8NMDpUk4/Rygtbf0JtpDiEL8H0CkU+QaI4bq3QqfXBWiUjABRXeMSqny/empCTrQ
KqUT8szirBc355B6iVsLr09i+tWyMaZzSoBuAXrG/pp0lHXjbFWMtTB9mQFChkeO
pvrWi+VImktTePPnE3KHY736pwwgLB4EOUCwVTIsjm7/Lb57yA4ZnF4k0oPizN3v
G64yYlgVAZSEISDjmlX7jAUWEk8OkzlCfVZVNQoMJGFXM5gP1sDGn9vxdcCzPIV5
wQn/RwcyFYbnDC1DICNx+O9PWywssPPC0s7G5lX8EqcKvMiJhZjsTKpLKXfwG4Ug
vQED26H+FLu6rjNEc05kRzoqKNFi21HmX3dxhN9zIKzb9vMsQyxDGlRRplqt3nDj
SGZQBghpXASmgoH/YFesyFg/kR3hSQHntqjrfzZKOtnAk8qP5R6VILC7JtGPiu42
SdpyVAtF8hEE365IZAnLVCcYm/GeNAqRHtz0HyE299MHE3kwV5cz6zvOZszKc1ID
enmVkpNfU5iQPG/Vctv+0R9i0FBWDhparPCBL8yxOTmNpqQB5dIl1Z349oKQkDXs
P8/Vwn2XJ6PtxIf/pe3g+pyBW+3clUWVumL9lV9UBYpaAv0qyUTDuuLlUvRNZ8nQ
CmA9f0A79WZ968+cFw5QJ8hs4RLPiMoRhaNYhYpP1Okd7j4DcQAvKg5lbJ9oELTQ
HAFSwFsvK5cGhefEn6OIYhce4Mwo55Y3W5urSw2L2gGSRF3dCv/ZLGQnU5AWo1l1
lmonNfC20qFNGzzys+nCz9d/z1CzC3ecZFLf0YGbdGoca5YX5EVjym0E7WBY0o51
AfxHGKycnj1K+FYlpXEpUZb6PnKUoq0PeAz4tVZVwGGcZq2mOWBKMu0Ib/v5YsFI
tHMN5m+V87P3DB+7aILoaao0cwd0FF2vUqfxj0Epfnycb7ghlDfhexbLrhhyF8xg
74/upcIoB5avqxDVo7PuZ9W1zYVB3MPzzQyJSVVqypo/6KwEJWWkBwlyIQZcCjlg
2FWns77vjUFpL9Pa8juy+1Iqpk1YRYuhDYsc2IA8xk3HGbFYdXxMccbXmBLX+bfz
YFKmuJPs0ooKKwbzWe98DwedUiz+tRaiNuTghV20NGbSPa00IUxbHfWaQuNXGgon
XMQN4grRNsf6vLxqBfzAle3tUbmdvupWvttCKxVJgJGwYHEJdt6RTFByfvEgFvX2
b67zy8Njzl3kYJm6rGHlPIlpaXwt68ARGK4FXgwEpoFjghwW9o19qGQ3rlBuBRWx
3Il+QqInOeK9VkE88jGkwO6tUVx9QvCx6bpyJHOPP/fqLBJeml0JAuT530R1q0bh
Y42H4SSnk7D5WIoBfjy2nuwi7Y2QCdEB3ZzkPRu+O+8wFLfO6xb4Gvs+R+eVMXDO
poHODzI1vTUbUiKQIA9WuzeLXH7I/nRlnQs8vgvW4HSxauTppQz9LNFu8jGxo7Kr
H7MKTHCcPgUGx0QVP1Rhh6kDyTShq5qQkKsIr5awBNtliCTPzcAA/gHNxEAd/pKN
QkGxhd51gSTZCKoQLHCF4an6plnNrOHyJ4dciApJft2F/qn8hYee/EgDkvsqXJNi
Bkroxff64hrglG26xjDyniH1bt3offVSPbH/6My2mqcpYUcF+1HBfxr4vFK6QgxR
msXRSR0g86hUuDhc95RI7Q2htfT6QRiRY/zFwyd0Ri+6T3YqU2aUsndDVYLY/YHt
5+azAweoM4usyWQfxS2He/pFbVLUfiqefHK5kh1hMLlGBjnfekteN937iy2fp2MI
KD4E/AKeTnk7cZphL8CgN3HqRGBZpSRnNirjhx4BQ7AN0Hda0FuQs72iYo2wKhRu
xgf9qxNGJ1krXhuyYj7ByrkhrPtlDSjgmcAgqj+WDLOTYHAwfsURmbjc59ita+Wf
ZR6cM9+tEZ1kOAkmzsUaW+j0cnZ6XwnOIpfYgBD85c62N2z9GCG7lxeUdLXp+RTJ
wTDWjjQHIFo/1g/u4zfmX81RWmWNCBhVruLaS2SCZnlTPF4NvNBJ4Uiq4cf0EI4Y
jq/E02FoLvolxNidK4M67RtBqQfNx1A3gmcXiqZBet8WH90C224kFA3YooZL/9Z6
DwBzJiLjLfQ8usajYvQ5elxLlG6AQtQegNWv1qwtY4OlOTRO9o8EbU/+1/gmgG4q
PixJuvkehJutQD9E+U3gvdUoP1+jfNGvQbLAXLhVpRwbiS2cNKzaswpktdJf00sG
E1GuCQOAwJJNa8NyzoGIQn4YN0rAu/50/b+5Vmj1PH0ZRUwSIj7lJqSxzh39ge2R
aws7Bna1aUYSpemev3VBzdwRODCKZIdFnIUOHBMS//J36/4OF87/tOgVcFLYH8Ab
HvXRglNMmTv4BKGMsWaJC7OuU3O2p4YOR+enRpg3bK4rr9cvzyjnjCjG6XOFhSvJ
m73SVD8V5IqABoN40ZJNchZCaM/ql3kT9KbJcw9Y1GWRhqYCfpm/Vb7/GbmLQdH/
0fISV3OrlNCjv2PMd9KpAQhqtlfDXcu0/LQ7ZbTm54Guu9OfMqiSKRjzYmJ+CnCM
OOYzWReU07Pksm6sIbY6wyWT2L4aVZEmfYrzWxQNIcnW0b2cUzQAQ3712oOvVA6A
3Z/ZoGmde9VEdQeUjDqG1aHG/Ztbt5Lpd+Ll5J3wdOirFb7UGz+YXBBbz9hYeTeo
aO8/M8VWTPVWww7HYQPNTCKmEsSBgy0s36TNfh++M4kCcmLFtASdYC9BYndMHDbF
MDAqXf+t+/sYMNlhIgAqzDTMgllFPA0JBvcbyVrQ7qdS0x9sm2CjLxr18J6+gXol
FipPzQHrO35jlKVskjWjzi9K4nRDNqwRcY6ED36EWm/Hlf2omP5LI1tIkhry7LyM
xjnlvNEg3dCEduUsymGe6qRsmFxGJpfE+5oD+I896BLn9F6N+dVVM2qNfGI9GOc6
u3N3XtOWc3iGAetLjhqXmhmhAn2aY2LJS2BMbbQqsOMJaJDLu75yhpvOmjA20+5L
izMgmHv4s2hdnvYKLkovEFsAclywg4Owl/341CZ5SEXSSgm6uUaKp4SjRjYqAKfF
FXBnNHhAlVe0klD+6TmJszG2+KDWpkz1E0m0L77QgBw4V1jFW0glmqo7HrDu4G+M
hT08uyzDbR4GpajSF1UN4w+se6+z0yn6tLQyUNFxO7xbtOkfCxHBwRNbbAwVHslW
kVKCwFLWvOCaekLmLDCjilxJmTYX8OY36Acwe1c5FX3rbzEFDEivWovpr7zhstEc
QoDpqiWsh0qFBVe8uXQU/Xp8m3X4xvYoFBFHsfVIkFNtFUhoX4oaXaucL6stSeBE
R30x56gOVcgwL4kbgCsuoMr3uy0hPEj7GpSxpE1SQwSsrNx8UOQ6HjyS6fbHCc0g
aZ3NfGex+36KWgVxaS0Zp4ffau+n6JcAaEKJRmydhiBhQWssylH4aoDUCt19Gbou
86nxi794y5tCxaZH3y/gjeI0nb4y5enbhdD1lWupJGZO/sh8NHs13VLrYxYaChIk
576QdpZU4MdQydAZSc/2T0OoRlyFhRTT7BfT/rYpWi25JlX2dvy8If5/Qrj+h/2y
pfI8mWG5YyKZLtnxmc71RaaQ5IG+0AJosVg9AI+HXuP3Gdb36M0erpT/nNOo3x9f
psBdERgq+4kIVdBkV6TV2s2lEnHrMwZ5XWOp/aDsMzD+k8C/NgA12pBonqIu3WoV
HgHvyjZr17OXvjz2BVr8HhaNJ7FHMo6bOOzdJTk8QCSHNZAecXFwGQ7tRj40MP4p
B7qFxZ4ACRMO2G2WOaFMhxTZuMK0vvj22gWn9hJ15TMyCnQYtzuXEeUBgyeZLK3J
YSY/6M4IfcDgjkz1fas4MeDddIgzajTbfgelFfuw0UhTLOG4UfG9+LyvAc3kv0Mf
rDVQGZ5rEH4Z0/1YjrvEiESyULgsasN5jGK3pwOccBcJRrcet0nl5lS3LcyqXwXq
+YHySVWxQZdj7kp7r5zeNfQlustodZWPXRW6ysfkGLSG+jDjzfkT21W3PbfR3fbM
JH84l3POQ2ostvHhrGoXwpTrBLdUjmlVG0PQMriZLfWth/wXmhJZmVLAcAU50ZkI
tyTPvIt8d5RLSyjGs/mDxggmKp3gipdvPkUPGD+2YTObRP5h6rAo4OUKosaUgMK5
RmSHBLsmxvq5CeyGeol+eUCGlYTZUBfucmYeslxFmcrbOp/fsegbS0ORSZZeZqsA
QhFuTs6lgsoAuHVa2ApnHzbYNy6mf6HmdLXnyl/sZKSxavZSy+69YdLvThkckK+3
0NO036tly6sewXVPAL/Sb3xLty3KkMD1XNUW/zsVp4v1JSRhLTzGK8gJ9xqNCoff
/UBKqgTEEklwQw494zG+MIjhuChVhIlTBQ0TyNRzhPp2n+gvEYdNFS+LgPUkd539
YV2AxC9X23A3hJsWabK8BKgkLS5Al/InKwybfmXEQVGhyHMU0YwU6VNMQyrn38Xs
NoE94sU/FOb4CUJ+h2ArB2hHjHP6h6zyZq/DMSrEhThcwrxmRbWopiQOcRhgpMNf
HnZ4TYWWYpbacFVC6z7k2BxAmYLQ9/mZKpSult339JL2xJdAhLoQ+Le7Dq3i2xZd
99duPOwZuzD9SJxYdDxZXjWvEVdg4j95aBZldrMbgf+qZ3iFiZ7d8DDyhRuK/D4M
Uv2Dxd0WncnMfjMB5Wlo7AT7JsLlFwNJniPb3+WWkq+T2FP34zh1fgwHDva3idOo
2S5QeWIre+MXe2y63ZOVOt1RikjjCpf/KsQvh/SLBS2tLHc797MF8bE7NahWwdbJ
oPX0KT6Ej8T8PN9xoWevZFJqpyuhhwsrj8bDd4KMB3lsptVyLJ6RRT4luOUAZ1Ma
FZt9eNwdt/Vo37d1OKueJyx+cA5rBV5ZIIAjT39btSFgDGPQLmManfVJC+vyQ2nS
DNkOO7qwl0axtrdo96XZSR1jLk7a0VUW3A9/roAcke1fr6z7GKXbFH4SBewryG5a
CE2OzLG1HbyjcVtbzsuDJo1/7inCLo+zyXfk9M3/wwdJgYiMaNA+7heogjQ2cbXh
moIEpTyS+KVxiSXBsd4MukBa9sn+A/XrhKQoebmQCLU58t/qQIPEShZ6mHBdh3rx
+Vwd2BujdyfmTXK2PG8Q9Lc2VJK7jf1YFOY3lFHRxXskK6y+BNEMc3kzkaaTOxz3
k2CGtuETgQ/QX4YRChrDer0k20O+qV6ptrDzz+O5Kl/c7rzC/YHANjST6JKoy4Ib
dvX7794L4kXwxFhseko/OJ8yZVKsvs8jZwJ95ka0UrYOeLq0IWiexqDuKC8ZxpyG
Z7bO4WA/qQDMepKk89VuzhjtIr0daSgf3TRwlK0cRflYATEhnbDxNiSf2Jjujcfo
kSDwaHjO5YHq+1xbi59RGCB0WNMbrAkTYuOxUgI6XBevowekN09HpKbRqXIEO2tg
kBarftzoZACktZdwysV1D8H9l+16exgOAFRD8S7TsaOEL+WW+7MW59FZe3mlI13l
x86eTNvjBJSVpSXFUrQ2ZucbUm1JxFng5M7vzUBGQSVQ9ZZ0A12ab1kQaHlWij3A
pZwKvBbVOcAg2fx3a1WlrOM/zqcY8rAWgf+9PCRmbRh9THyQ4zw+d3gueneCC+OO
k5PvQfqiVmWj/YuTdmImGi3JlhGCHkMYwTXgsZHM+7ox5R9Jk4TABcV1P2BudViW
hFPe0inyUbNZL7ygw/z1yM1vnSgpsHLvO3ZZV5+qkc2PaNy3m70s7yYSdR4phcq3
CT660C7kT50hEH8hqImSYBjRORdrAlX+9KmjNJXdHiBgrzILtnvNQ0TwOUdbo+qo
1W9mF9iXoRQmzwO7lBwstOvn4wKSLgJlfi5W1g4Owrq9sDO0Cz1t/Cw1bhwZdClP
JdDN2W5ZbddiYurd1BI/pdQwEjc08vsaCNqYyanhh+IDbNjWuUDzzQazL2XPs7ZM
+z4slkerwVR+lKJe2GVjtlVcXsSLghQ0iFI9VDfP+buM4AL8bS4OVU/y2rztUTKT
rIGF/9LeirARzF2TMpg9yyLdcWmDjXKoF6iXVZsD8MIweGeCqk9DytiqH/toLO7P
pw4Lnv2IybozHKxjoQJO5BqpR5B+1cyZSHhenLNWCWQl4z8jN/P/EweLtbTiZAUP
Zk1HTsA6+m+O7pDXcahyS9y7vxVLn5fYNPuwlnKMgodsPhIGxNv1seFsWGOayTF1
VNjDKHhgK7q1LtAEFi78OH9RdL4lOxdff/LBYKWakCJyJclMfpYaIyVVZFYzdLvi
KhTMMkBBuITq/67YFzGVhL1qW/yhc+UFJpnL4YvPmvoO1U0pBGH0uumIF8ov2AIK
pqSh6UL5EePmrAkTlryedj/GPXq1S9xLQL6zELEJi98zcQzubtG2l8UGZbP9jsgu
/YyroLAjwlWBJnWx4xnI4MdhDPTVYYcNwbAEFfZVTlQAvTqNrkR7PUR/+mkUAJfy
SMusa4kzn/eqfHyNNmdavoQqzvWEYiUu0QEtbtD0UEQV1QdZxQopurvZDdGCHIpd
qrF3fCWcYhBkb5OCWzF/2R7IZQYbmiMFO8T+8RMMH4xlZ6zcyJM7aAykjHxADEh5
o7i/GMeWyTRvNvbyUHOsA7FY2sJg5YRzqreGIz8rykclMkAxAhI2dfeoKZRhJTAp
46qCLnH05WXoTaSmf9tqgBRq2Tsj+pswOVxx9X6VYpZB7btmxSSDIg51/TtZlv+6
ck5kzwqQqAWbpIpVDNKfDY9xTSWVtKAWTds41K9BxaALPsFXEEVhPtB1vy5OFLpY
Wa9P/l+YbVZb3BASTYrcsJ6JWqmpl0H5m8irczw2kuNTrxFE/OW7nsmgaAHpqYCd
Nu/x6rHQ7LMQPgcMjKhYY1xBt9bszhe8RYQhpprTfvFvq7HaZFVs1eenfbWeKs+L
9NyoxGwWM5pygP8iJeAHJ+pS0V2spxxJUddfbVMOa+WpeW+Fw+6b3XEPzte06Jt8
JAdsT2acfL9A4WKJND+tyS37sRT2HEsNtl9TB2P13H455C57uxb0Skl/EKrjzP0x
o9hS6s/ikbhMwSGGfy7r5P2lLS2XaplB4fUP6LRplBeOKyKcYwvKxkBN2vXUKxHW
jChrH2Dsfiz7GS2cIXWiss55he/o7EaCi1JXXRjRkU0xa5ooVFHuhM+PzfwsVbdR
NiZzzxZZHsfLwr/odCcRK0QYKrx4+4bMkOo4RzSK5VmrKSnmRtdqeHLpdLGoCC7r
NIc+/+Jx2IK7NjaeNg7AQmE2D6C8c1MpviQsjwY7nALJWDH5w9kNqrWEe2UvY41V
q6eoJTSsPYsf/h0yuYC814pVOLoW4I51Vygf1I5N32Ncg7o/XiVkYLP7RMvYpeIG
EODBwIRoMb1833d5kD5TJtZ7ifUFx698OabWd801Gh9WrB+yXFaZK8qOlvUI8d9z
5GSbGGy3kyqBSDIGkLPU2QdxLJr75UBRjEeOZAzTVvLtKi0Nyp+UlOu/eOAExgBW
HAdTlY9lbhJNp0Ij9+uM72WNqXq2hQCDIWISremSoSjTUrrMpF0yT/5Dyie18HNk
Lrj1Tt0z67Icq+nFPLtnOYPU1gGNNQtfe4Osx3XJ6H8W8LVbZ+VV0M5mYtViYDm3
sqylPIPi58JBvfVXRgYAGvRXrX1RBvsQ3vrsuKQP5xS6h03aNonIMiuzRlgJRK6P
QB3K3Dq/OkDbs3NLlgE7iq7HPvsY7r9q3svH7rkuqotTEr46TkdbMinOUTg35B7U
h5stW7+xFyQHcP71R2z8agN9jKN+TwBOo85Pl5NFGgV4cZ0FRkMgfYmmzrC8rB1p
Bzqc+xPEXuzCkCQCwxEoQtQf/T+OwwmMoBr7e5K82fzidMTtpS3yqtE1BhPtjyYK
a5ZTP4cO8JevLKknG7LRxrFu31Wjdf/WguCspmMmCcva10ygdQKWQvvtSIXaSszo
boiNBZv0tMEPpzUvsQ2Gf1pte+H6logLnZN1Ryv8i+b5+ki/BHIoe2ZSrZGltuAs
/CrHgctkwsLmHb2gMvNae1rdgm0kxChagZLaEgaactDoZfcU1M9wfP9M4r9PTvt5
8eSrPjvROscQX9PjS+4aM8Ap78n29ewsGB8ORDmFB4LyvIX4XEnl0vaikyPLk7l5
YmnvOYBlhTnm45c/4SH97/lKcheTea1uI+VqFcFE9+xi49mfn/PB1uNShGgqcTVf
o7g8o50WK9OXrGM1yidsytpdHsl8r+CSrnwT0hhoIBzdP+VpkybVLyIDx/k6t9NV
1VpSEYWazVxDJMYm7G45NIwnye4eUG07T4VZsTuoMzQBu/p8mxh5AAZR0D8YDvN8
2IsT9bjxZMFV9uI3exHVAdOJBTTo598O/1Spgj8Ff6xI+Xes7T12VRb2jVrSl39Z
SrZaHyvLor1HE+qYfbNeU6RxRRMyE9LLkTcGhvMPQBiG/WMYrkXO9vLPj33aziRb
8RcqX+zNOGl6lXFkX1SEjTn5MSgRr89yO/xf6JAu1yTCusZ0o09VTErwcgqKCxUY
ICwNvZk5I5AEBdzSeXD/mIj1xlccnnLJJIScVq5IViqE6spMINfubQLCjmNPTTUp
Lzrp6G6O9A1IVsxnhTT4k36uz7X7p/YRXI2tNP6ZHELkFKsdRPxK49X2akPqcQlo
Mg0RZrSYolf2UTno+/85jBw5MaMvbq/p8VXhhOEG5p80IU6jBtwhRVeN8+mtkfXX
ONKb0AhI+JsatmZ6kZ6h2TkIUX4BIsIRnSrk93YuXJYOuX//7CDzBLhO3Vo22wGw
Bw0kAHyuAhYBNqe1E997G3gSzQ+WXWIAPJ4la0h2UXVOYFYtoI4eUoQeppV7tMG0
lS3b/dO0itnllgiUm+3O+4gS6zdSkFxCs/O6ijCQswWwVn85d8XXvctHF3Azdsol
pATNeeouQcykgoNHLyVbO+qv1FyceeKBY0u8hF7ofGB8Pa0g1gHZtjVndRai5FXN
swxMdAr2jyJWN2kOnIJeDNDtO6XSAgnWndySFxuOU+6e+bKLerOM8xvslmbjptGO
YaenOvePbbe3WU+0t9W/D/AgkkD941gF85PGKXb1JUScqlJcxj0818xOZh+vCiYI
JCLMqUasSS4IEyFyhgEPrwYZPsuQrKACyvwknC41mo9BSgL0MDoRoWLA1gUDr5g9
tLEs3diJ1juaOQPZCA22FJ82eCd77weuqOEpMCQnTEk/a4sSOF9ldiODq+MoiqAi
TNgxy/mheCGVPSCAjRFjT4EHuPxfcLqKpbZDl7nJLu76xmswVbNwAoJO+zn5z5WP
lKKPFLfsW8UUjZ67W7PlBvdJB8ZmwxNlXcz8slV4jmthFOhcuPlyCCNWFUa7sR7Z
KsnbiN64iNKzeqTDczIxE4HnBVEigfhZdbL83fuep7M2pvoP8gRc/8L1zF2K/Bd8
TuJL404/JMS/GHHIfT2Imj/0p52err7K/ddt+N0xUpWF8m2MR21vRRVi9JxLGCnC
OgVOJQJtn25RaE+1qvUBK7pCvvZOsW7Rv8XLxVDx1jVr/aV+w9YXiUaOBOIlZ9wq
iNO+gef16l1yXztE1fxMV/L6ON676QkFXP7xsOfgd3j6kESw3QdMhKPyWuMdgSIF
asuANwatUZBAt6hEm6ttXu4lN3ZahHBASXntLzjifM3iHnrWiDVbsF/YyUAD/at4
bRtzd19xi6QBNlsQ53Lg//r1FEHhKaZga7sbvAypfBdyONWhvU1zZ7fzqju80uv1
G4Hqvbb4lgH1QBxoa3DxeRGmchOFy60QP8hqmWAKRjLEyfC5vxlvpOYA6JrpMU01
/mChyDLWrzDH8uXUx3LuWhRWor4JDIn08I9J0J2rNRtMKpRqvuqtW5i8FK3BBUB9
KI/ncOla8Q7WwjprUGNAzMGOXOntElDGS2/2zryupXvCR9ps5ZexRxiabD/0iVWz
ZByIsO9nVCCQ4PgdQflWqssR51ZMtffoquMxvQ2UBdZBrVTNur/EtDkqjg4XOsma
6q3fAHk+II57aG3xVphqeDOlPutSqkrjKbdJj3RHm3WDSMIt1a6oOWTqTWZpuXVb
V+v8T5p1zCHguqXxl50LDkt8Sa2coQlXh/gtstmNN0+tLIafkLrV2R5BWDuo5szo
fwmbiIbmID0v6+OEe25slNbfgAOJ3j7AFgadB5kk418o7bYkQ18PTipX8vQb4k0u
lxo+NTEQsCrgjVmnn6qPOMIfvwxDtxsirmPxsXaj/WaP6ZHhgW24+Ps7ph6soFDK
yPG/nXPOTPYVfoP86INi7RJ2n5lAKBMFd90tyVoWES8TTv+Y5IfxYaAqhL5SpDi8
oF2Z/WIIEKrOvIMDCRtzBCuEucba6b3F+X4bfe9eIzBkwAcQmdFpx9MQZAB2gPiS
P4CtxTghJON/sePtIj5BLdFEt3Gkd59HQcMdYk9pI70gIRRQ6DC3h2oOm0vZPazg
dMT9UI2zHC9L5eRu3bacbH7FpVFST9pt4Cz0pyk4F8/VfLuAn40UaamPw/bvMjE0
JIgSnT1TaYolpQiA4ZlKHuZIyJiunZJLKgMbKyXAZeP2vCYlvo9/tXjsbEnrJW4P
KM9ESv/ssrwT21rRIAsOAGB41L5O9wh93AOckXzmOukrUF+RzNluzheCLduaa9y4
p8z0a/aD9DHQfnDhXDJVS+2Y5PPJsMFQk+9LynP7JaW3ECf7Yg+FuHJCZxCWDKOS
LOqjqIZsDI++ZhG/dc7cIKjipAGImyAGtNttF7j5jjZwniJXlCWkHWJFaYQ4Gw7T
7+NFjgPcMgH69AYynba1tqUsANU1SrLks8xwPiUnpQRhmyLVMwHdATEKIogdEVuE
jylNHi7rAy7eRDSzlc2kuA0sWFka0ZabD8TMT33ASsNdVw4H16WMAgvKzmzZVxvY
hs0tswgQI5vU9Bne5AtNGYz+CQRQevd+AvBxaVq+F+4FGnyo/CnXAYSueQwvay94
gQ+Zb+riOj5wG8R/JRn+2rZMX52HMtEb3OHEIbD1q9H6/yfpJCDogvCHVrN5Lukw
wR4kFZHUcN4GgCVTeIqcPQOmh/2JYOp8uvwhWa0v+oxA3+i1VugoY/wqYn0gnfA8
XxUut6yJ5687VphY52+BPdNIpPs74TTWqQ79XS64v7wK6/Sjf8R2nOHJ9cH6Aoyc
PBZfwv+hXc0id4SeYWcKTNE2xxj/yL9slBKG1u8D8tMs6rvToRKqLvNl6BaJb/Nh
urXgD7h6kmfQdXmJqUanjFKhmGlpDUeMFXD9YHxdmK8woVJOVbMK2EYbHY/7cVWy
V4aq1lxpxIedsgsVvuBK1/TM3dAZC9Pz/2Q3ryjNmvssPdkC3bCHbQ0Y6cueyDP3
3oK4VerspJL5tWxTQiXYWKEmFL9snza5F3R1jsOfPgQQdgTw4jFvxZkX7vca3cer
aPTMLjJG9MkDhb01DzJzfVUt9d/azqLjTkSIzCFsWhILTcZwcbg7+LZMEeCGqJR3
XDAWryqH9RTHyovhafTNxGVQxpLc9I4tfYYcVboE1o1TJG2YvCLICIyftYWVmNXU
zYfr84sYcRMN9xCN1svk1Q7qTFRLe4Ihx5Lf63pICh570Y1q3KKCTmFaTiK4461u
KzewNOzMD2H/oFlwuHDYELAw69LB6ht44FxSOY9baE6jZqHKfqmwb8i9bgV289lo
I6ih+1zmjy8XtSErZLG2IpNSO2DQFVwXLQmC7AuT1uC2H0xjmE6oj3a17jWpN3pn
Xr/y/39dmTJhwzW+xgpciQ+xS8wgi/9ruPm00J9ioW18zz9WIOFYZITpyfkmoQBe
2taFzIKzG9tsmJ+rf/znhpJtaHPdoVbNM9JeyuHLvnbzb5YODRFwa35GHMIHLnaL
qW/Db4UcY6ilbuyGiX/Aopl0xfG7nr9zhB1LyXGpo64jp4cagpRt2VBJrzFrfRUV
klQcMdvDv0TwzQBkWrt1Kfw5Rb5gr/p0ozWHcUX+6s2yWO4b+b4wbHBHqRkN7OC/
NEwWwrYtCqtd/E+DEK4Rp6TmCMdgc3UF2Ot5hmKQYIirbGdSmiZXveRMiZqueGfV
nwSULsa8F349Hhqluxqur+tI/VgedbF3gXEqmrBAUrfdogxo+/6agSi6iPczFic+
nJmlUZnmla3c2TQVJP1IQDhXEd/H7SBsyafWue0W/LHACCRZMWa50QQ0QZMX7lFA
hkZ8oHprP92+pdplVlxFPiR7aqm/K6Lc44uTXU/cQTpciUuDKEGQ6N0u/wXuVxZM
QXXTjReLuMdDYlLYQJr5GgaZ+U4rbOFrTXvl4y5K6pGUJ0Y4Ycw8KnMZbreqjsNp
k6OpTaoaeIpteOVREZyj7s04N+6HqdggPNVUKNC8FTv7n8NpVz8uAPo2XJc66cw3
5SyRcuorEPdVH/NGAoK1ZPYyM1Ch4A2GhOjtkbO5DE0LN6dN/9QAzAP4GcHkuC3y
jSPzzmnIsfpWTV3lWTZcdIMlycYJ6kStuQpOOwkjVYzu2V8hOeZzEWweQDaeCQVE
NHnSSSe5l53GCzxQoAIih9broNTLkEFNxOyVPUfNRxYIkP3+5JuRBMyxUxGFejfu
V+Mx7BHYVLYdCcD/GFdbTUDFUT1R8BNrjZ5RfpsBYWpCarJWRWumQmVNpRLReaID
Quezl0pfm1JhHD/UMqcO3t7WaDIj7rOHimVhC0tJ282UXyygxpSI3Rjz0JC4Z1HX
RrlbNGekFTgBRJPSatI7MYR1RYOX+1kfvFDYzOun9dic/QcfEvwZPUHjuQxvfDXn
FDfADeyKpaHx5/8BO1SOUQFOmUI8BRvzCXMeLSbBGHyaaETMOWApgwnvJL6PXVrK
cHuwJ0RuYV/v8UfTv6Wyawx4W6IwfBFwf0CbV/NUoDVXDKD7H4qKxzqNoqvup+At
JukrUIy+uuZdJZDKbrEoLpvm70mHwgzXCWIS7G6R0JVkzFxrFhyIFsP0TKmG0JEi
X7KVfXfJTvqAXUa62qLdpI3GZ+mXnxFWBfeEi0k7AeD3oEaWYjyenF81Tc03SrkT
X7W1HiMIgR33aAOLf0L/kO0MmES6UDMerhVWqlF1U8ZDyu6GfP0aX/IUhpB0hHID
X7DfjGzTVSTCKABYQfEk3q7pPss5PCxbaMKoq6CSz3J+ya0//GKkzIzhkqHPdOyY
0e1IBerHXm/I2GgsHbAQSQsOqhxfOXoSQBPVp4AlzT+8k6kE8p+R/hjwR39wfdS9
CWbS6kYi8Ht0/Jc2z+oTeAtjVHQrgLAyOGwXSvhY3J8Ilc5zc3Fe9w9FmQjh7S9O
SfsE10AW//7hUSlgqopjF49S8evAZga97ID3gbiZVvGpl/CMAXrDjxDxuuDSbeYs
DspEESVwWVimkPV7a/v64Ox7J1QxWVkBAAv4h07mYEPaEmoRTC9PA9SXTbnjt8Qq
iHDgSgu2d3tuu/QRkYYzD8joBWdIUHwMoTSlKOT6T+BTwYp0q0goSEAepwS6gjEp
YlzCX/AvDUosayf/ew6CQfVSc0YwD0fPZfrh83xFdW6WOUUXMTHcfCW1aHmtObud
VEzQqbjEgAHzKdWyFCJqJPJzksuUBv+BWb7GmumNPDg9BufqzooLI8cF9MRzsWCw
4Bv+ks6bJowJbkSONOVey6uyQdl1RRIiG6GG6M/TVZsv7DU+aC7NdDOAMnObvGIV
4OnSrOluUtauU6pc9QbVg4MfsFKQ/fKHBes5xa+LgnXnxLnOWap6uePjjXp9KeOj
Fjxgb+qrXF2Mx03wCmVqJw/K/TLAlRfadvM3kMhekouy/DpEBOJRc6Z4+BXfiLc9
aAkeN3d8Yrl14HegHB6THiYSRkulKIu+ziYWItzFQRwJcPAN8nDF8FIX8Q5PNpSH
QCNvA0uL8CN/8HzbEg9RJnEL7MqrrkN6KpKCw72j4sgqU6R41Zjahgnf+6Rjr/ov
ZGzQ9YfeYWv92cvDdcrlBzyvDcZLF+Z+UYRkb/cqu2eVl+n8+4YoWoLEoYREBWN1
X9t6K265WbG/vYbMebt2HOyeDjmcEijJrazFmstMnljkWCVt4R0pTyj5EW5/cJbI
dtJW96CcEYVfmDWGOQ8dDaXLPZCim3CL5qp0xpNlkMlCRjC7tkVRbmB0UDmfgvLa
ZpBRd1dNrlZCHJU+ngFRHHG4CJCDJjgufbpt7p0symSZ6v6VBAoIQeBVA8XWiJog
6KjGdGTv5Xz+AcVDkVeRiYeWSr1Hy8j7ureclAy3LYL2tNO0Yc/A0AKkQirfjxuQ
B3LiXAx0bVt0m7xPJMHMGDD/UCz1zZLgjZdtzktBCQ2R58vJAGOFu8VdY6vqOCeQ
7KJbE2oKkrMhxtMe3gh7TTKw99XXzY2F2Zu0IFIuRhVHDHOb4tkPl5KgFnmnOLkx
tsKbOBpRlkJPFJbc53uXFscXG0NmHv990Y2Yrdv8QxirplHppRm78ebVdxFSBwSu
4QE3TxHqGjfi7hdhUQZoVQWrqpLIGAWXUQzX/BpvHmB5bpzisTm1nZz1Yk/Envae
XLGYjso+dSJuRzhDdkB4DzqUhon9CCPeUoN8DIopXQK/jGKMtxsYuKcTQuZDirfW
uvA0bgFE0P3p8Lke7qbS3JkwOWjW6vh7yuNWVbQCehRdalSx9jIpCNinfR33/Zjq
RzKBX4bXkzdMcQLAw5Ui660QG0GBCp/9gZG+QNVFYajCEoMb0p4KI6s63jcx2xO6
7L79JJsmdYmDfeX7Otd7NeTOEi6m+292e+8aYFP4WsBs5QKMsTrm/gYE6QkhGIMY
SYPdU5gCjkOuTfL9IVvnePBugHBbY2dsBU1YeuELvsBkI6a48o+TcUEOXGfVE/tJ
/DrjGsf9sooSeGCX2me6kPOjXnGSxHxbI7J1b76nHUyH+5rFGdpN7yJZLCWoNSEa
bNSNLUXD4oyH1JbgRaWeQdcGz3nh135eZcJzJ8m9x3YiqHRIgBCPBEQOqjpNgrpk
/JaPucxqFoGlz5rfSbH7dL0+xOKjBjBhDdX217S5ckiKuf/vs+/wm69VLDV1M4NZ
4/6cxr0hmUz5b34ECTTbxrett2h6qfzoQlpTfy8GXELoSR7shbiwInJTdIjPvhEB
WIVwQ095h5i5Sh2o2IQ092ApMzLXMb9Rd+A1WVh+24BfeULnMZ/woWzA9lvmDrKC
0m6RwGh20Lhb72oAvyFAH+vcWi4C7bX7A6qXj+y0JgRioeMREqEoUTRIL8/Y1pJt
EjTcvMYeIPCO9XdWpDIJeeFgR5yYaW3hXSWf8PG8y/snWXXs+9CkqMvFcYOBpJzJ
0o9VQXXHtz7r09qMSCc6G0PTZTKD/PgIXTE+0qT/NDGbbA2SaQeI9c4oGuAxI6dn
YrNEX4yLEEKQnH0bVR6WLsZBGjtYwTd1w7EytK1lECxUoZQy2RWP9BEx4VZEPY1l
cIxyd/51PjZwEf8gya/gqNQOmqdH9S0yHEIHsJB3q1xzSycCD3bY6mo/yW9ITj2p
o+QoCbsV0M/Vk3DKpD8ukHUPurs7mgaoQTF9rxY1ybObgJUZ26Uax6RmvOQKX2n0
AWxB5kvtQYzEVeH5xhgJWU/odUPvf8PkraQjn3oa9x+hx8AwnR9/0PDXEcBROpgx
CMe5dhYrwK+DSXpWvHXOaLTpmtLKBniNy1O6EF0OcW8PDUGCpp6xS8U8XuLOmnc9
QxEF0oUfXWXjAgUX8HCnkQkRPjIcoZIaWOOUhwTUFiZCMIVaaaRRv0MIU962tufl
fTpldsdGF7wUUwa2UdZYkWwXTGbgDuavk9WFUkwF7VRg4XSuwjh/I9KJ4/30l5b6
CBX3vJEI4cE/gIkQgou9zW2RtWVOU8G8H7Mgd81uKE3E9q0MoTbYrS4Fg7bAbBxf
zAR2iX0buNp9nak9daq0L8+t09GzZ6D9CM9Vct2E6LhmJ2gNtk/PkGkj2KOadSbl
6q9Coj0FBKHGUmFlAI66inAD9MNWT5gUpxPddi2an/En0kJUgK3M6LhweMjF3SMF
CzN50f8UajKhs2H7OO4ay8iexbCb5st02aC19cgj1jvOtdGGkYtSkSjize44bkkW
BdSEG3jjbykwz6GSIkaFxwhvqpfiyhYadh+3xD1fALustXpuGtsVr5QD6kVk6OHo
7ms38Eip5KHIOaFhqE8v7nDO9jy7DqelP8ZP90/ekcFGA1MceY95iYYK0f7n3xSk
iF4zHWEGq+vE4uZU6gg+zPxuCKbTBq7PJShb6pfdFMDj+rwK1SosR6HUDbhUfUIw
WtdK58o5sK8G0FiNQO+CGlwJ1fThhbTvr9KRqAWQfgxnQFZ3rRiAEAqWukSQuy+h
q22aiVO7I7ez/EViU+3N1uR2/LysfmBtSS5zbb4eA+AJ9lY5Q/hnI++f3HhsVUvK
nQmPhhIyRJCd4JEVfA4F22D3CK1mmCmNNED7WL84m2LhuWFtuHddVGIcxud3xzyA
zoTq7uknd1JfCWhwVoGf5lqGe10AZGm2gBHDGxewKSPi+FOl/ChJzMy/eBYI8rqN
iYJ7BWheECeipivHYUZBxL7WsUrzx9mJNdifKNr0eQz0y/2YnJfb9ePhc8aO3t5I
BwSszUC8tT9pP3A4J8uHDPfOId3UVPl+cXhaW8uOQkpspFNr0L8zBlYFM40kWZE2
90CMng+XDKnhrpGWk6+0a3R6MJ/90U8vr2lgRx+qBo8QtXuqFQE7omMJLOrehCd+
kgCMmHqc/jEWWIMQZYLPqwOf5PxfywO5cvkj4BQT0ZIpitREROzbgxvfzNCyGDyD
4rJ5u16e16IMkx/NqYk4xX4k12CL+2jb+2E1FhVfrmW4BbcBqhkiRsYsK2v9oYGl
4aKKvkR3zPjn5BiGHaUuLYdfmnVU/2TxfndbmVde5pAsKUnaZ5NZtxJ89rPGCBLU
kqhoVMvTO4T7IqhqaV4rlWTcfsazYtxC7sO2zlk8TR0vmlH8S+XlDTVluk/84Fey
koG/mWUxYLZA2Trxbq9Vai4c9qkH6qYTEstT+XF2fWfDCjiGxQDVNCzvRoz3UBff
8xA7+4TDxXMvc0Wbez8G6GNrxoQvP0uG+h7wBgFvn0lYlOQO+APPjPeBoAXlJpeT
HDXVL/Nsb/bU/tpeCDp67scjqka444k0SlTmIb9JDXSSDg7A3SIzpjnNOpesgztj
689c8ya6APapcRgqqF3QTHPLsJhZUsAl9nOJ9Z7cuN/FAFF0nDgkxCI/yYMYanTB
XwzuNItOi2PTVtUQHtCUsr+OcVhDRr/8eycJL75J+UHBUjmRzqwZS/HSItNRAZJ8
1FdC51AWG9UJOrYxW10rd5bAYC8ozyuPU4/gGvdcBo77iiPtUrxKqWRpNyT46uge
rtvVd//mKHTCU1tojevbZ6zDLXAVeInYOw0fhrXDaYOTW8W4XG2WTpDEI/Rob6jJ
+vGmLGIHVx4F3yzSutLScxJ/ggyy43XJMzzkWPGOTxUv6oZwLI6zCED361+ocDey
G0zvlk71PJ0OAJNBwRXEEpR7ON2Z0Ck8u238M87SuM8vXCZJ1LbQqx1aRU3KCIRe
Dqw3VGJXWC4eu+PqZmSxFV285VYSxZZVpz/SHcBe/ZXNXN990d4BNhROvKs1y/Xw
XNXnAkwxKQHclYFt1pDblv3lao9Q5aKJWtP1a9320pID39LTvourm4ZTZvgOVlr1
JdKveJnnrwPC+sy3I5bDPHj4m0PsnGqkKQYknUogGfyUDRVLwVQIlZl9Zo6nhjh2
0K/XjlKUf8pev5EiKRKMtCtz2SfKKkDyrNcZtbI5P6/YD4400d7eAAUjOkOoHa/M
/fgsnc/58zMoijJjkIrxSnzcZa/MnzFp7UGpHxMJ3boQHd0HIshoVIdiflXEAdtF
9gIqPRBP4eTrfke+YY5oOpScAfSKP2VDpbJ2adjC93/TLRl6muc4DtgBbQ1lCAm9
+DGV+utXyRel+t29yS+h1AcG7BP/8Z1VbozLB0Gmt5SXhtJd8wbsKo2idBaMgsHt
kji+aucGyuWtw4bS0rXQ9XoEycAfZfjaFVpjzdggLzErQVBkaqRO8VC+222dOwUF
gb2fCzUdIYISDoODn9oZG94Qy8+C0NTIzKPVuNoK1Z0epNV6DyjclH0LNeZo2LXE
rXvmQ+/K2h5k1Nuud1QPOyiKaLncsv3/al+Cg/Is71dUAJGu0sAIQifo5Av1kSZN
AXsu2Bu5KMTfuVziY7KSf+0AT1unQLN22AAro8NZwIRqNU9XnwzX+20niD9xFnZ4
oTagp/EoD60cAmgEU8gK/VCX2sIaZqkrOLkUcdD0vSHz3MuC7pHX1Jw18qYgl+3R
2tt1V0HXlJSnKBN+ZxQLmepMuNWGsvXB8YRGrPsvuRZblzVmuNCCEpHfwW6qcoJd
QnFdCH4oSZDSW65msMjwNgpJ5U4DGDZJM9S+L6K4C9V96cZNz4kXxyOlSFV4b2Iy
dxlzQIAgZWq+gS62rr8g6Bw8WnMoVKW3d3d1/2cQy5J3ruIA5BJgHgksVuJODT+L
0ETip6NqIw7ooIQuGbjfDIXLJRTa849KNkZ3Bqh59ZNkwtep02o/cVNGcqbtwOxl
1XCJsak66MlY6P/TphxASw1GvnVoiDdHoX0wPBeCobgX65xql0XYPm4m+dVZG3Qf
nJVj3E6/KNukD+08CfS/vnN5DmQGyVkEMtEfFe+PScWXG6zwzRrvATP4kxJwyO8H
U98DVi+IHQvuWRZ8fAwc8Q2rPDAk3n6Gkwp7uIURmyIWP+l4slKtjufC9l/4d6Mh
D/SzARYpoxvTVjWLc2rrye5tuc3sgicpJXxI9u7LideWCxApoVxOu9DwnhEIAVbd
idEYh70TH9PS8a2rLtInC1YzSOZyAQdh/A+UwBqWKk5W+rAhvVcUS3Z/qvyLkk7x
Nu/sTdFuoVdkKkUh9gv7cF1QyKYa5hrle7QFN3Y91LwK6TqpGeck7zWU8R47+S/y
gDsNGvb5Rhq8J9DtmMyYc0c5Y4dU96gtHby9uVSdIJljVlkZNp846OtA0DrNzSbM
9gYim0MkywA06J0LUaKnwcCwer5PJjhm/XICCh9DgyjFGGmL0XdRJVJi3YEOMSde
KZCSoyDCfcJN7oPj8eV55y0OwQmg41SXhrZ2bHV+I4sN+rC5rCJINMlhE+BQSguU
Eb356pjfuA9+vmwkUEMUOxLkkTH55h/yHe+IPdFv1TOllMbRIo/55yRZuZW2FKa7
Aut4kxMscQUtHCse5kFoiX8Ak5iYczANH+wDVSSdtSLodBaVuaCMbZDl2ccJgio2
y01S4lFL42FdzkKmuDR7/lCVvNyHb02mi94FoTRUhCUogcuhhbxzvt5LvJZbOu6Y
clo+lSZf1MctqeogbkUgv3Ba902vVJZIyRNOhdYgmjlJlhJ+/kFhmDzegNYUJWWC
XDTzSqJ0z/1VtgtHpzCGFhlswyleD9KHNoKSUdOySjjRVOYon8eVubqY6OUuQ+hD
+oi3H5lIWCCXe9vp6iOXN+XUFfNgtT9o4go2VLD+LhHHv8mP6cpy+AsRdE+H2CEq
PsXLCKm3T33w23fssLWr1s+mP7hPgyxSjtNbWgIhwzl8nRDDPfi+BW9DlpOmDOBH
ZpcUce1uwtsdox2oCRGTVOw+KGiLKlQAdSlGmI70afUg3Hspu4FD0HnXrBujNYDn
8GoA2/RzYBhG7cOGlA2o4ruO4gJESAGTrJxJwqEoZjs082GX3z1OYDiE4MmwJsku
uDYo68uiLWy+3Wu91LK+AQXishBMozU7WrQsxpp5y38YFt5PBdH9rImb4xW/P0rR
4j5znctyXhPeA67emGsvQ5nbmnDgDBabn9j3cmaNhgWAGFcy+O/aMAVGN3odGvv5
J2PHvm0kmAVVfsvFWzEGvauPPi/FfX/lgNjh6ZDajpgktVOovOGXA8TAUfw42sdX
YXzYxiVKDOAToUAAUZjkbT2tmjzasH/wwEkS96xpGABJbGZubVZ13rYiPziG51lq
1F343viJRpDeFwG0ulG8L5LuybW3ElPOOuMVLTWU2ABdj8U9NWGNQ1qgK6XBmUNE
4mgJSkkfReh0sSXkSv+1kw36gRJG2ptyD9+aIU0NLRwkykka9zXdvaMDjPXc+szl
FUNlTMQP24LxHeiTCmYCTkTisLO8DrDrCiJHdyMK62/ftjmJBhKxYM7qp6y/3XcA
cZceQGeEb+AvAWRHSRrZYF21j560WVuwv+aZ1eeONIPeiIILUEkRVxby638bX6KU
LMP0spEKncPe2YkT64786hy5L/lVRXdfKFTQQ+knCV6zje0y7Y1srS9GaKRnI+8z
+bWeBiFpDdTJdXkd1SkdoIKyWqijDJTE5zZluk3wKotkeqPVeLCuQF0AZ8IxYiW9
rEig9uhjrBnzDf00fY8ca8Lpb5C648yDOFL0sr+G9Eb3czsvdoyTSxVI+7o8iXO1
VbpNNcuzm9Vi3CvDV69WF5KLfLS+b0TTURXyCqBuAKzuBCqZZVQuR5043HD0u7b8
gEosuRquOI49RlzFEMXCbYfzn61Q7ObPXLhTx8N2iDGFMA2UGPfBIILrDuAby7KM
30DBCD4axIiPnoXk9FXr25CcbNMl1ELdTBWUeGP6V+LZhuSoWfAyBvVq21iMoQYM
IqAEmhQ3AYzUEWxeLuLx8foFimstmU+BUsl/LY32fkS9uUGto421QNjQs0/hZhsy
PvKn+2phTX33WfD3Swv6jsrV1jtpDOFf5J/aD3EUmTwAv5RtPWP5xIOZdFtrscqS
QeTEJHEnyvvMHsf0Opvvx5gAT2qVlCjjKI9KRky8bwBdjyTghGnoc6u0xsNjR2Ce
VcljaFPZWDAONE/ImMMlVxj6vJskXEfTgUQeHVZVn8QuxwLZS45L61OcHaK/z3Hf
LmlTa1IoqmwDCcRqkVGI02AnMBFNtOF+VjeO8/WCuAKydri08LlhdQMHdNMZNC8i
hGjnnt/OM9ywbgMg1j6MPjjsfHysr6n1nr36/P+9JygjdIR6dH1QVlfmI8lXsnDj
KrEODdeTsM3+8jlkg49dzG+UUfoEMHydBrcA7PjC8o8GsE8bZrgeqIAENU7yA2y9
nsp2ay6zgkFYg97QEtia/MgxCaeLCqKx3qtHg27ftq/4L/CvmHtxFL6KNsjBeOZC
0oF8pbbK42y7klxUdHW7umNNgk1XougSbqXZuGKWo8ns1oKPeGssVR7sV4nCZglY
rv8Ng8Urv1yMnIVX9aFFwI3OJR3GqjYJa018iq7YiSaS0/QeZMyNiOyBkg5piD6m
39rcgSOtNhn2E/aXy2FhVrof072jVUcAhybTImlNlvAdvcralIfQwtZLgMdoVjFe
O+VjO0QhPOqMamBEiq4UIAzTdv+Q141GEDHjBKDKud0zfaspSGC6bpla9DClhdNT
GYYs/M1XYnbVKAxeQNfMMYg8ut05Q0GYp/oGhWBtoYCXbEvHVoLvopT57OqSnujh
tqEb9aK2BqAtDDjU/eQMnS57fME+mXVSDWEVsSjZEnuhZjTsQpe+E4+eE1unM2Rk
WVdTy3lI/pXxoKexyXOLMd6YJYYKivsPUzbninROB64ns5pkQUrnTaeexEuUd+sz
VdUQdl0sHVCSdq2K7drfQ5D4R2WnzMUjt8r2XcT/Z8egEFuy3oJsnB9uvSs2Q8o8
z8CD7292zDDWSxQZ/99kkieyLAr7DvyZAxUwZmFWeZGv3yJXciUn9WcnLTWbEjhk
GC+WwANCCSwdjUA9HlXFt1Tmr1ovd/AvPHCbbN4DtJF05THtudQFjZBe2Aw2AJfj
Dw0aMrOAS5YkPhwmFFAh7+oqJ2jdXU8638lJLHawTA/ijX2le2Fqn4LTn8Hhyl4B
u1wumP59CvKzDio8LWFPIGWTCUVNI217foY9hvuPxcHC4nCDDCX9+8LFd47Oemkg
qX3wVlNyuIWUd30yDcpNy5IsJQ8nRpys0F9RrO+wIwLAgB9h1ne266NQB3AoxFYC
Ff8D8ev1mnadp5aoJ1XG2YCSvyRqebnQm9R7ZM6Ado6VR9gzDaZr4ImOZ8QG3Bo/
smCqDjUGNENrWN6gaV1gmMxaq4VyoXeRGw5YpbUqsS0he48DSs4ky+ATIn73cG6+
tvVbKxcQTB3F+7ym36yt6HvZ6kF+a26m44lWhmq7zUm3JZoKQmc0TCu89zCNefV+
GwfuvHMbql9H/hBwE+llQW8cu/7q/SbpymFkL7hiNZG129dRNkdQcK0KNH3FJ63p
5xrxGFldkGaakAaHasKjSf/pFyPH6GhrrZJ05qwMYhF4FOlwD/2EzQH/pxOcHxBB
HeAzye5K4SjRWm4sUEi3iF0fS6HIczvybIRWqFHQ2HYLWSNYa27gaC2N5PTa+WPp
sUeuzB3IeIJ5ku8UPJCS/BEpmpToWBi6nvw0xvrdPrnbGLBWNO5d1BFOdXt0ntNI
WFQ0OzQP0hilgDC5V20LZiTVJ1MesB5FfDrpMJbbo8rFdflSSWZaDwDG8NkbntAV
8bIVVXK4rsmA3oZjNRIpXiplYqRrVQjMLODHkGqzP4rv8tr2pGF7uptEeqyrPJS+
2kfMYyUgAe0Qfobz7ovzIxYIain1oDBqNujbRoqcQBEU+ElK0pkso2E02KYC9Uay
Z1gmhJNSs4frulcuh3q/yk85V9Txyl7LvhP0z3Cp7lHOJLPRwPgyH+rje8HBhZEl
yI2UmmazJ6HFGNBjI6qDpXuQ+WTUwulvT/WL0rLWAFbnlmcFl46Q637UCGiR4TYo
IW9357vRLDuOD+Tfr5IreJFHhF/hYUs27FDFlDgusMube3yl+mfeD5BiR0Rc7H/a
pOxZztgVi/fLHI8iZa2qMLWm7C/dawMlVGY92nsbuWliMjrf2uVIa5jdppd/QpEi
dVh17IVfnW2Yec70wrfV/wKeItcIUL4PlidYIGpj8Tq+8Dcp2sP4tAT1wJAgkVzM
G6XFVl1JoYicUSA9BL15U1OTc1u4e/R/fBxTJO089xvQyvg7F/ysruJUhz/AyFUT
W325bqzaIc3hHcte38CfacqdKzZ+iKu6oGx5kHPhjwu3NpJQLyj7a6wYoOgb+qOH
Kmao3BKafOhvHgH4VcBoYoHthhxZ/HJ4lKZWRglX/FesN4YKk97ZReouEt5k35U8
Yg0eKhaBMkGeqxNp+ethVODynDb780x6yIs7HrRCTSfeyQFmFM4zxi5VpOn0ZePn
kstYC2N5NG2YDYVJBQI7Emlnsn5lHt+C70oBcvjiBtOuRdfc6BkKlqPn91ybxKsh
vXRoUgqsADHT1g93jBrJKq/jSSFKFuD4UWi4JW/l5vtwBebyVUVVsl2MSjdMAZtM
MNNsHMG15QJrqd7Z/hT6KikKl6e6CxtCHG9ukaP6+NFiuLvM9MwdKAtfJ4pUSoAi
t+llByJQaNOL13zdVTJEfH6pCwaYysOiYXe67FIvHltJfqt+hjBr37strzdOBeMo
E5o3IKF97UtisALfzYsq0+1WHfXeIDWfcZpCqJfOYziZmWoILUMhNvcnQfPAzMV7
UfxdNU6A1dsYdIQDXhyInw6hxWHucnd91TxErvDi/JieSldsyVQrzMVVbVgxqxJC
fIDFJ+JARYCscoiLUFXAN0jfn7WkzmMSqub9aRfmyeF/B5WOOVJ0nxktZXz2po14
bpb6vPF4sPshep5gKqrtpxDfHLr47htBb9eBYCH0ad+rACPIz3qAMi/TBRxiq0a8
ywFZnNXICZOKU889D5O80TD9F8H3nNge4no5pL46tI2H0aaWOirTkeKsEOiApxkQ
F9S6BMx66dkwIY9nhhuLwdpozSwQL3E/WlexFFpKcQ27uGUp2f7q/3VirRX41wNY
+Ywf37TgLBPLLuz6qCqPNJuj/Cxn6OcrTVRDMxM9rkZcrJtEzAq5AcOjqrUldkms
rVRuj1RIlxdxE+HNXbqfPj5cBi4pGVECl7p77N0/ViGjjSTH+d/AAXlJ/GyNRb0b
rO9xzV0TL1astZAXM0A/kuA5GLlToee08El2E1BOQAHVV/GvLjEJbfK8w7MK+LHb
vdoSXP/7kykYdtIUEbHqkzeSxem/A5mcycti6xERy83EoGP8Bb8eNfsBLFmqU0HO
Ca9LuKt01rCVPyZsN000S/zfjwgEw/IU8VNwakrnR16mJnAh8lncQ/ALZSnp8F9Z
NUbAdKXUand2h8BJhZ4I5T1QiJgWXBN8fH/6Fr5Gb1skPUPWcMb84/n+g4ng5i58
QmEK3eyb36cok45uo7FAH1XRVbXHwK9DWLSyLlcRpma3YgzQhtJbMmOr0FaiwEKV
63OVEbloli75YwtBdlhtmRwV/9h1yApzvQkRSaGXL4mW8kSNfnfmk0lrwnGF4mGt
awbkfHJiJYV4526ZZ6fP2yq6DubcytB6UJIvC1Fpr9VsIq2SAXrZmSQTOs+6AI7Y
CK3fnYEPpEc7Of8Q1Mvg10xnu7p9foSYUbEF7ZzdvQn3Fj3Lt/ZWgv5nuY8OQrRu
wohhc/GhxfHkyNmJCloJdO2WEMQmQbEARpp6wlop6+MPGMfgPez6ERjcZe8LY90K
GM/Y1FQlmgnss9kyE1pyJrL7ajPPaZGngHHI72Pyhj50iz29fUme2mx5sbu9loBE
3MO8yWuMLlHdjuV4OHEROldqYMsO7Ioofs7ApiAWUvwwfDBfSsmdqa5ZuwHBHcdk
1WdyW4/IrK7FRn5xaJqlUNSv4ej8CWbesCNyW/Coxs5Cll0kS1ObPcrluRS2X2xC
Lid7E+XS9aVMhv36uvPuDJNFX/4TA0PRcWiBkEMo/SrLuQQ3TkOB05pEE8bRxB1o
zzYDzQWboNwWoguk4HN5EQk1qldosGtLTvJU7jMSZP1z1IZddK7rHTWC1iWlOPDI
QJ+/jjHkQ9zJsy+NVj3rl/Z90M5Y1QW7eh/5iY8EzEJXOIV/bqmiuimBegJQfUkG
LDKFccAEVIRK6qG/Wtc0eyi29lXW3XF7bLZZ4mSr3QNEATFnXbex7h8F/4YEYM4W
L2KVyC7yeo/MrXC/YNYKMK6pfS/gkXSaJtMGaEQi3tnlrJBy19vIM/CPUiVAS0rg
Xqh/+h1m+8FjLYtFrE72EgXOXEzIyC8AhRY8vfzC96Qq+LBgrMCW7kegoc2tnNWz
udynD7oeovAn8l62grwpvKuxSW0m8D0VQIvq49duWPGmu9atKo5wIy1ZWUIRgkFv
1Ns26aVmOdlBw7L8Rf8b5Tl0D1SnLsrgdA36Hk1NWzQ0fQLq/fXr3cfpaYhThQDc
vyoIGDnyoPqbUWGcexsPQas15GXjMWTIv2CEaQxAtTUoLu3EtdbTS4Jcc/NpSLT1
16xR7HOrnz4GqpYRRvcEhysc+uRiVf+eDdmgrOpT7mwtd1QfZqz14Pzgg8G/Ec4q
6kML+MxAcTZe94DoqJkucjIA2Dygl6sVH5vniT0G0GTEim2B8BykVHhgecngm5Ae
HADR1x6IhtaDCtiYiaMvgxD1ju7akjAclwWUPOrVKEumwzdakW1SFIQlYWDDSnLc
o4EAryQm1IPeBzue8AbXXTbG+Yj5QQpVIWcpx3yoJveD+lqXjxF9sc3RUw+g1mS3
4RvK5WjPrc9HC1iaB9lseU5rwR7LHqDRvKf+qu4xXD/vTivgnMf3XNLo1u4sn0+Q
9cFY2UFgUG83C59kcVPJHEXnU2XuuxzOsA6/te9tBIbGHCqcqlOTWNHGw4MPQ4oK
KQXY6tz/gtvfEm2ux6BEUOXnkEvZidOmq2+ggTvQ85h297fE66W2gr35sVfG68Mz
yaOHExAd6ZbO2ZpCyT0MKmlsshqB5wVqb7SwH+SnRwvpdRahSMiMXPvaoo749kju
wNdcSJl4slPDjdmt5RcpanV5RKcUIOcE2GhAx5jMt/qkquiGUuej1TTQEqgK9xwU
p/j91LQVkHi/ByynaYhQ/t0wYYk0kUPSPQcgI0wbqP77vinTiLu43DQZf/rXbJwp
uERBuyZUetgni+sAuIHJFpqdNETwOSPN96sv5pB9hLoewR1uWzDcdQ1x413B0l/C
ceM0O9rIokxEUzRtSTjs84frL7q9AvLU2P6gQZSjX8lde7HMdS5vIO3qEeVZzb7J
PG3X0tKo7dCcQYUZbKupV7O3k/JrtFKv8JroBC7o4kpTCqrpN+NRPqLKI3PSCUUj
OmrtG3x3sWq2QxpZdnZIoeRdeAYmtwnX1R/xX3KFc6GcyS7NoVBiwFHz4nCBOzrz
BK9+c1PquBoI2qinzcw3SDqU0h/JBCTzz2hmWrJaZCfkzdRfbPZXDr1YAa+FXEEj
1AqtedEHDNYR5NCCBo6C5C3TdoN4M9crH3MJTO0b3JkXhOO7E6VwqOKbjzbDbgtP
lrIDFSzciLd7kWxwvPpW/dTxr8uZLOTfL/AShP/Pqg2IrsqXjvIK4tNyldnvSXwn
gScoEMfol80U0LZOrmXBtpOHZOIWe364gZvWTvCqSD99QDUHWFTUWhV+R6qLXONe
JRA9C3W8Sz2AZo/xP8G1Ezckvgno1APQJggPeq9NYuVIvn9thKDHwyjNhQbTsGFu
ZBc295ZvxY8ZYgqapDyRWS6R8sdOpbe6dVpVVwkhGYBPUt9rTEnIFCuiDBXDRpZh
y+yKJhCDwQi3deDJU3K8cGw/Fk6/9MyNOk+AHyVotQ+K3Z23r6HO4jwkICz/l6JD
JyAixHejfKZTvjcjP8aSWa3F4jx/MMRAqBDaBO8tsa2IEJOtTAiVqOWG7OIEkR1A
tHenOCCS7ewA+dmDzlBco1KuHHKhS9h4FjDWlWODEM3p97hZlZlO0grJgr9QR4vI
4wAayGAKmnImrJDioqYV9pazDpYeZ9nkEaiWPWL3fu4C8bUhZfmTDLNKyQCvhpQL
XlFmkf+chBSuMOrvNwS6GoT0oanJ3MMnx7zIjvOkg0bpsCakgCueQ8e8Mv23nhY7
H1WFouBvX4cZTWabJ6Io+nJkwFQgEKvIcnHTYFYQGPsvHxUavTNOpFqjhrJFp1ur
oOIi04dqvOJH/SpQjo8om4NIY0hAGYPoqS/F6RUsm6MptDxOs6Zn0BS/zhbMTnjo
kda/tXYh2X76s1zpgu139fpB1ymi3JZn1AgsTpAxXaCGJtcqaH7SYOA2R8hM9p+v
xBVd/ZubnIdkkxt0+bg9q8QavNOAJoZtgh/UYPucd4NFOTKgAbrA1G4bcKtbR0qG
jH7FDheMFnFbAcHQzAuoXVW9eASHdYyG2CUGWxiz2Fgn62pU7VByfOzcrDVPJaM3
rnWBwy0zZVKWJF4Ae/qrs9wE64EOw+EpISLAYLMSXGzOjSZcZcxmqSrgq6+LmQXq
M6y0vk2cSt8R+H9qbkMbAc2x9I6ntgaVuJrTNZwqA1vzP2o9L814nnOPAKNBdeZp
JDGYvanIzSsSngkfZUl6l1tGGakvIbWbqJVbN/JNXSyVZYjn4YrPhToVwVWIoFZx
Vc+UxwWgvdIwa/v3Vf02jTnRqkJmxzlSA+ZiIYfa1oI9W5G6hKxpzH1OJAczd67J
ZKLEwwqkKC0/K5OghSXy5IcAgPuyDTW78B384PCgWlXH01KjM9zJlVc28KxKaiGT
EpOnSjDblymkMnbiU+ZySLlmozztiTCn4pdBX6/8ajN8iXOtwaQ/k1FSpWR976tE
YToX+kSJfo3WWNVPkSVouCSLd1rYMExVCGOvegtYZVQZ+VV54B68K6sM9O4YoeXP
GqShzedqxItbKI225Bag/xfPKBQXMBD96j4Ry2Ig18RUNq1RySBAu8DPoTji3uV+
Y+iVa9Odesaakm8ioR6O8OZn5pWpGueqSQfolc1Bi1wa1gDEpXcdZHrdPdZyxhIN
FcZ7mcdo86f5jCGtlYgnHAQMNGfFD0At6x06GAo+FR2SWa2DwAI9TCnq6WaHNWZe
FRbmBcbLRofcFciA3DRx0o62jI9CjIKZXElwzSzNNbwBQwshbe6sHCV9NakMeAx9
hcfAtEZm/TJ4Ahf2kOsJI8QOe+aBNNfoPLEQEZxlIlYisOvTyBj9qr3oQsj6Ofjk
+MOAHZDcFyEqci6baVP+IiDvMJpXC12iITsDmDbeGZyH8cK4TsyApJE7LxkwPlRZ
Le7EAVJAWAV2wLt3dAWOJe0nAKHc/JZHzHMgH0mKlSVx768mx3PWl2dh8+A4PBEG
ZxARFZt8Y0juXG5qCGGkVGZ4AsPy8wUxC0vPJNNXZCqlt/p43MI0QMY0QPsVSm6a
NosKehf9rkNf28W7OVymnt7lINqFkvvt2AHmheiVr5ephpKZJasfOwN7z/su+HL1
1Ita+HpoU2JYo077vZUHR97TMbCBc0RwtVAWrY+i31KTrY0PQQkZEh8OdOzEzkKB
n42s8dydtiNqJuJ1JWwqAqM0vUF9WY3MfWlMB2GJYCGQ/CWhGI48193CkRcDMxyT
H84zYwEltcEMTDGtpTyPx0uS+86A1X6nFvCCpBezCMjtMGMeU13dUCjIC8V4qy50
ix7tZeu0/kLpYpoxVeAxXcKtqDj7jMzJ5pejgoI2SOSKW89WmDaWmiVNHJh43QLj
g2cuns8HC86ePZt7i1sA9oz4QrGiVKv0Wg5fQL5PLr92Cy1TVxKxNQ6Csp6xnAnS
PCb2lAZ6KCY3XQMFmhlotWcvSvDvZRORr8pcJyNZyAf/MCTe1qGBC9SBJvk8b2XC
38+gGaz9xonJk9A0hda8rQOS6xeXv43cYXgrAJwEN2ggd+obzvJ4coBcs9PPjQUz
RKbTfEZS70ON92BZoE4rUaBxOaV8Bs2neJjeIm/7iuvGRHt8JEL1gKxTQz9YC8xB
OTk9eFK0ncZ79A6D5TWN9pU9zv41azz1D352AFDDD16QwrWAMaBYFxZ3IFXSE7qF
0y65O/gcTJw8U1M/dPSa5tSTC5vnPJ4bCq3TN3LLIx5ysR0L5uiJl0ZuE8XE2pGh
Wc5K7ZqS88Ql+B4D+LNxvrDFCVVqj1cHvViQjk+LBjat7KCI8BPvPowDEOUUKrvY
gxSTMI9DPYqj5RfulNWbptZYuWUHZuK7gFPd7QMa+ghKQw9KfzXmHGo62Sa4a1R8
O5S7+vmPN9C8q+goBpki060MgdXVDpx8zzQdoYLX3L53A812vYaWN0xR0V0OlTtj
/aOWWJpC6JDjUEKvTM9gHtI0aU3v4JKDURZ/UQEh9qKdlEAH/JWw/M/M60Lm+OMC
qoC+ISkYSpW71TFWeK4MsWu6k2vZEnHcXZ9k+PtKGTSBul/bIo81Z8ApXCDCK/VD
DyOD86s8Cd+dFczyS5bNJ/XIR6DjxUIU7z47iIQSKhkYs8fZ4V5ik3DPQyjtHuYO
pgGRzwJbRJkVu74R2ZvQRweGPrutJWzSKLFj8lzhr51gOhQjSChEoBFJpys8QB+K
EDwYSxAJYNHdLxj+4NOmMXsckHgxeY4pj9vOG4W5S+RDLrz9KZqecfgcjdyuc3tq
SxexEJU56xdI5gDSDyutmtUb+QCHiu1ldVCVAVcA6g2q1hKiC2eLouV9Ot3CmbjH
XcPvQ1LTOajMQONMGqLErj8pO36qzv4pVRpQlMdzaT95KDWB+Em1Z7d+am/jRraf
7HfhCdBhYOpdL91jU3KeuP3E9rsdSrNSgaV57a78NM3zEx41l8ghkUs/vWB1iECZ
1qvUlgdJLGX2Za0uM1u/idw4COzSlkYnMtqFDrGdjGJKCkz+2EkW8V62Jb5HuB56
wzpHj4mHmrJusy6Yc1Niqk07ruG8YdAytbc2zsT3KIzKUiQA7qgfyWmBZs+72fnb
Jxh0dt9yuJ3X3Me+HFnLcOI2Ttc31yCFc5SP73axpCyCFcvXpFqC46k4Lbx5f3s4
J/rfTrStcJs+dZsWoI7V5qlOnEx0DyGYkNpYMUhc5EHqFagTJzfP4LnoF160Zp0a
zrthY4ysMOEeecdQrHTlcIX8FZ47x5uTKcNuDi1d2YqC1TP00vXxEFaQtowDGil6
XZhmOAs/l9tYukRuTzF2c/CXnOU4D6VuTfo3loZ3U0VnRhLwOgq/jIpfYTUoCfYj
9mMKAdXcHcSUYLuEuqCvdzyYd+ZkRF8ddL4q2ewQAzXVmUWUYnZFoxbjmVIDqebI
K3kcegKvoxxM03EcjonUwbn3oqXrJ1P+5yQdqG5xAnaqH6I/rbz7JR2Wv2YwEZIB
EcK4lw9aTikM18RzNVHPTGH/pjaIRuv/QPeQkZwZFu7pMeUO4ta8FZcOJBE1WiAS
dG8Xw9OX/Nx+caD1EoeD3rKNNddQH/2Uv8cIr0SDWsvzYdAQHP4a8CDPC10W7jFo
08kzESHUJAIRxLfDQ5drpYxcaPWKqBa5kBftIKGFIBvUaQ0jU+oIW9bkJIxNdGJJ
LMQx11etu3nTHVwLdOQ63bktD8lXVuXACzrk5smiJcVzJMveIjsZPynWI3vve8CA
pp6F+IJKdKAhb+Rp73jS/RJQ8RSMWlwa34d1a8YprmCK/7JwYkFxU3LXSkAygNgt
w5JCZ7ay4cWwIGI8HYyQNPmXVg0jRjKISiGs2B91bpelefOPgMNVj+hPXRlVu7Hj
x+HWuxPY0JcSsmu04y9XdIWEd2ezZ36xvWg9VexcjDIQFRco5R0yOFDQ5s7lUbZ8
5d8NADRggXGSkiYviKLngFWkMNJU0Rr7iHyBLJd/q+Qrz7vZLEdGWXMu3SnANkgt
3TjTsnLP2duqSl8tsbXNmQatjwBmyRc63gE1WXdMudbG2s4XhjU2j7gL8k1wUir+
w/OGpGTY+cBlNI7GwJHMyPgCHRw+Xxgc0GwzoCZuxml5H9pb8fSwk1wOk1iHT7xW
/x4UksjTdiDFLzESyro6Xv/rSzllytjBpXPtbAewsGcR6507yDK5Lodx8+BCN3Mo
JzIxh4tpr3m2RIMZh6L263HAnwn1hPbv3elk+bh8+J9sdLyXc0dHFkcd7XUX7q/N
qgRE8xGJVg4Tcj2iud9VuP2O5Ljpww4NBigiFbs3KpBbGPd3dwKv/ab/ov2iUJ72
x/fWzRrAASso+3/7fhbbQG8/7uqrPbdWUMmhqVuvLQuZtSr5BAswe40g8/ZxJyu1
9Bfcovne7jua3Ov5bpE7/pSWRQaFaWrWf0bnpW6DnynBP+6VeUpTcC2lxi+LxGuc
3xRr2dYpzfC1n4XqroyDqBpAlfmKJdfwdfxAD6fxaZmB/Bp8h30+u/l1XmvRYZja
gJU8zs6jlCY8guexXaorNdKWaZcb+YyF05uLrcs4yVqnvfq2yD4mJDK1BQbn1G9g
T0j700L4XruPvJMQVMMQ94wGzrk2izEcfcIVm8URQBxX914ItmXQzYV3L3C95qhN
KU6DDkNSjCPXa8z4YQy0vG3tJfP3zdP1uCOlIBq8gDOcxzovqkPnIaTaOd9c/vV6
mIKn+PkYA9ieHhZfdeve0DTZ8eu3i0B8gjhIYXT9yPJwv+eH3CbET6zcHUMZ/fWp
SJ4oxe6tuXm4OP11sUxMOC502nVgTBVfN/0g2OYuNy+emOSIPbivAWgHXvJxfumd
olzIES/jolNZkxeQx2Tvp7u1MqzXiZT2vI479s5CmL0YuF/XuVZfn2NfQ0ibhncv
Yu5EqvW+1L+kYzAxtLpEcBto9kVK16QN1ywFDwacGUaR81QGepB5vT1uBaOSl6Ve
NuFqGW3bRtQu9NwvE0yBGtdTN97fRTNE9IuGzMGqKDEtrCj/d6wLzFeTmluPDUJw
9WFYyjvxjbShSdq1ck/v34yInUA2gg986UXq3sCfhR+ExGPOXGQxffqHEa/ffscH
Hx0fGlIiKiH54I+J+HgtMGdb6rwd9H05iSogt3cMgZ68iM1v8yjmU6KOg6gMPZGt
s/s/JRJteYJxz0Mw3oRS35ULtNUc2FWnw+VGW4pybS34eDfbbXRaTycUlvE9gXcF
0LTDk4/1nv8VflmiGLovZaq8UUcqHDeaAVT8TdrFtRZrUPKdIRNZELT0xUbJPJze
Q7SNpU0TGLS+K95aAFk5z9C+lEFIE272XkVe1tkfQS+2Ca/VgTq65vytGrz6oCrO
CSu5YqlgL2eMW45dIpzL90197XIHIs/y8s6TFFCmdHa3Hso7iXSnxzp52xwx/Vos
yVrd5pXOWCSYwWw4QvsM5tVyz+o+IQfS0OLu+TIrA4GIwPDePZUqR6olRhEH6XB2
CaS0BUOcF+RruAGQxygIR5U2Ud1AmtHpTqyTF1vKiXMq48c0HA5aHiPlh2uc34Bh
4rDSn24Rv8f+nZ6DXLrhuBAz6RvsgwmiD+wncnpF1c7ykrh+pkbyU0UcnXkJy3XX
nryLmgFrY9nOAQ/kEspjZlVulkyJaXi9CPigk/Pg6MNSzLIWyjaPV/YevnvEd/4I
H3tr83OHCW6c0KgpYkH+0ab3J54RQcbLtCkii1ic7TJmSbL3oabD7/2BDFyQnGaW
AVL+nnv9xGROw6a6VM+FUSUihRkS0h6S/OFGqpBitxcaggD5edzWm3OHWGa9Kp0j
WE/uvRokgXd6UyPCHqaVwGYhh6sL0JCjZW6/FPfyCHkCqMzreXmuIgHeHP2ozhfv
u9699c4R1JdW/8x4HfBlaSgvlhJSVZPt3ENkhBrPWgfxUPJCCDzo/DV0jxV4PSSu
rP7UjbaSQCrP4x2s+slGwA/L25thewq/xaTxfkYDsTzAzrpzwL01qiG/7Ac8C4cm
0GDSitVphGEXTuYPlbAjYstDaalo60Xe1yYqfDRAqtu4WTeLf5VjxrBHXoQGSxF1
buicbyVNFrtGazR9XRZ6QPdVadxQCQU+SLMvgLbxWlosWPddPfp8G4XxyPCDVLPu
m3/SoUcS2YmEt0+8n6eXAQc97qnOyuw+FoVflgxefVyvgEaIEvPkqoZWc4fB/gUN
wwDvkiI6Z4LwjMyN7CiI7KERUhkvxFVlx2ir+0hdc7JSuzetLUq5NOjfSefyiqOF
sI/HvvgkhNiVGg/i+CW2eO2Q1h45ZfEcG7eR394cbvN6taf/1exkxKwLyFhf5hO/
DxF7WVUcdo6hqjkNRrEblipolM13d7DNqVh4NH16qwAYaTmCx5L50MHuQHG9CBOY
xs8rzPDTel5gs2ygqOlKlH0Tmym6uw1/g/anehxRRno2OKoaP+bs7dIbw4WGC782
RmlnN611kNY4d0q4aVqi5EtKs+kYHCcXTHgKUVHpK64NB2fQJNm2UnKJdEdM+YZP
s537+kV2BXHwpZeVCPWSf7REv1PMUTY4cxXuoOM+ECwA0UMWjySEapuNz0AgZ8yE
MJlnxKKPku16A0DLeB3mCcSidiLJmpQumjOWOIpD/i3MDSa3kIV11l/QBWT9W5+9
1SuN8LemFTtnHO9i/AQalO0adaCjMRMTEVvzy/PCz7XAhcRrAeST4ls7mlZ9W4FQ
Uf5xPGBxq8E8V/NtTs08E4rGcc/OPxTLszRM7RYakEEW0euytHtxe0YVZeSoMtqL
hcRJyRwhZQA+BeWDWLBHN1v73zcUgXE3NKsgWKJGFaXcid2BJnQIihxahK7b9eXu
7KCHHqu/WOZksFdoLRhI8UHUvg5frLh0rRbRzL0/3dfPKvptbgiihiRlkn1WQMNg
4cMC4a1FfjvdpwGbKDSzE37FL1x4SG2cSR6xHmEi2fqtISiTHIByRii35hDvSFww
pN9/daDuVxP6XAmnBIrtApz/tx6QGY3b2f/MxO1HTUDw5hKmaDI+J+sDNqY94ypn
C0eA8qmBCom78Uz2BUqgZ7bkXoLPTwAy+nknBkXo7OCP/p7s0YJ9J/CHv/7uLEMS
rPOfvKVbvc5gKM03NgjsJB/ckzVb928WLRfoeldC/IUtkNxMb9xEDiW08auXXtvH
0FeA+1DnZlMh9dFyoEKvPy4o53qyZ1c2aE4ROO/Hi6nUv9IJTBA6nm2WKoWvOALZ
UqsWujj+3tUHKPUJfU/F+UQ3ofNS5HfT+WhVQuxpZlzaavSpY6ru/6G2mPl3U4Zo
wKslhToz67gw9UVdpLfrR27Wus8Do5tHw0CdC/M5Z7Aefjw9eanKos7RobvOLRq4
D3COwynsBugqxtiGNXuQ2SwzVBsSWbwVRJtoe/U3+M+iMMxaoFH07/LgRbXfaXfC
i49qc1+D6t9Xdiefdt0esN6uKWXHc+R73CNxzWVogrzYd3tj1CLiGVYtODef7pmE
O+KcNen3CVoaTPtlMF8asq85VPId+Cmsac8BUb+SIl1X65/7I3JETgOLVfHeczs1
3a3jItogxgij2P/xYjfKhewOQl1c8CxclduN2UtAKYcEzkqX8F4VQXsQIobYmX/I
kVJOemY0vCGceVRXc6Oc25hEebmU+v0xwX1NCtTcH8oWQhzE8nAZ/GZFC5x9PPEx
QAq7ZaRQtn2unTdQCmYpVqEeDpTrwwYnbjNradm4LGCc8MzD/X8LWmrwGJxf7gFU
U1UemB0hPQveqktA9gmLxgTSKoY7voNneZOerA1PzE6OZYKAZLuCDQYGbdr1zO71
K5cDc8ZB7/OVdQzM1xQsNgqrXJIudIHMTB2MwTEfKYGYQuBBKGaYW8OJ/ePKpcLc
KElrHV/UZpDyoB+tcplJvQEAGu5e1gH8ZZzUIgOPfTdQVcAWIrpYjDWYHqZp/Wbm
bXA3acBFYGNhpehBquQ3/psaxQI81DP5KqKqhV5ZSX+3GaUjxskxAduyPwD4rvn2
NPav7Yn8+MPEZ2JC4lRGHVa+Vzy+eVGCLy1+2ELcX8/W2qbiHHip56ljaCeh9Xa7
ihxqyfIMLK113qzZFmLLF77ctRdzgj62wYfUv+V+EcrncxcquxHhmOQKR2Z1lwpS
gG2OMlGguymRFeqMovj1Z2ytisDtT5bsEhwOP2kVNmdlT6f1BN41YyO3FndQwL1/
vZo5CoLBBVC/sDvx3ufTaeexT/oEjbi4nXfETIlR+4RX5Tkahf2XdsjA6jswC+3l
g/npWezsih86ouAmXHUUQkApw8uX4qZkFSlFBxdhzLFEltH0k7/YLcJvGI65THat
JTUTTF/1FBrrkZxDD5sAKNDagQM0bkm2HcUiWYh5c2tlkXaVV893aZbiqfB9O27L
PPR4OYzrucmWC0rUz/7ROfj3cPZ7aQys2wnPGBABqj58AfCzYmLIu4VfaoUNf6yO
PSvLOa98Ym7NhTnplvnI8XcJwMTddAyEWSxnXUU7Qq/WYbCMG5S/2PCxyQuUhVL7
+zQIFZ+umafTDTzQZ+zKqK0e3un0LNFrRDtOOzTVHaO4oZqAtBe7RvcuJWQuw8dd
eSJ9b/Xk+piWnrrLNw8hVzgyuzHxW7kOZmohLsFx9TJe1nHb2qDbA9A1GnIeBrzw
DscXatFb6lm680LNp/yiHRIjoPzyCD1hznmNLYaXXh/rgpWsZ6MpUHBpdzw3AubD
8QOp6+TMSu7enIEfeql0aTwvZUtEU+X25BCkZVbbHAh7FxwlbM4/KOzxEAKK/AyE
/x7cJEQIr9/bapVrugBAvAUcUbZ5PpWeSReaOTSM1JbAYFLPkiBCzjCEtnGX35kz
CTH9KkIb+cH0oAEtRU+6mLVpKu8fgkZSKVHxLu9CE3ff/+KyZ03Vv62ybmox5ixq
E4PzrynRBM2ibhx6Tn1VJZo55nfWmXDtNF5xHtu5hL7AetKnxQCPG7kx1ggDH4pz
PgHT0TlULFwkcj15eI01OlYHNxy4zBeJkJWYH07SOhN/blp35xzosLnFjWzmlWSy
aMqx8PsnMuRGGhQAxgat8XGxbDut0GOvU1DfZiBJaXmbyorhjf+U5d2t1IQPu97e
lqrp4+uECjRH92Pf9NkN2uxfBBde+JbUiCUgbLXRtYDqU/CA4OcCbuUNFabJz3vT
FMY5hlLaMbUX2hKjFXGDlk9J+NxQ+6H80eyBvJm6+EbmiNsn7nSGy1E3rnJBQYc4
Oe59NpAxvL3nvTBUKJGVRdPxI5QLs5AH6rhCXOXvQTzUDKZPvpHw5/OIfULdd3yA
+c0yxRDDHwY2s9VOiDXW+EnVoB+SlM3mfkBTmWMpcBt6rtsHRbDvkrNhZwsgljjH
gXyw9K9Qq1SWeNyRfGQ2+ItAWptraU8uvlYR9IfzayT0sdf8Eav3wWGLIcSKSqnJ
ACAvxYoylgNPAPytFDOsmxzqwtQ/rYSvV6h95+1H++K1JCsxc6N8de9F6UdEd9ET
ndH5cGHYAaW5xUarbGAwNnAnVKo5TaBYFFpymSENnWLfs3kiOANzdTcBTeiWuQ5h
PWFS+NkuYGyW1GSM62sjmMRESwxV544HmxVYZS0fPzUg7tTNfgYX1MUt9a1mj2nz
vH25KyOP+O0Qk+LF/IMuRfjoha16LapSqzO7I3WMjbH0/s1zNd6j4+QAPY+nDYG1
nWZWyNhfiWzrZ8CnxzYkNSra5/bN+wgQJWt5Y1TTz8cdEHpkGeO31dXxu5wy3bs8
dfsXoZZ5AtLAcsJJ4a+LlA4bsKYgnm/q2RxtvaxMw0OaMKV8LlLGiEMnVfuUH0EB
Cl5l7WZqiOOYR4o3fjX86A9IEhgRSPIVTiSac7bosqjB/sATMylvPSgNX+to3M4N
Q2nCX5Pro1Kpiu9rA75KO9BLD6Qzk6pv65xPEtVvWeAfOhsHX9Eh3i0kLhDBitpn
DHO8J1BCpBsam5FVtRLWRo9QqIj9QMe2/uogmigRrkPJab4S6ZM+yRrsdPic9NNk
CYTtgRPgtJ43wiWwiFEIL86Gx9Xemnr8GwgiyJUGrS2LKWs+4LIR70WSXyX6Qcq2
Zv72rDvNQZJ/PQNk7ddBLrWrUwHX/NJu55yAG08OAbx/ErdCn/u522e1lwuQFDIi
wwr8bmOgct8sfcExLHSO1FESu4nk4X2ySdC+q2vBCAKXwM0Fa3DzeuAiCAXY4fbY
ymX7GS8W+//gxYYR1pboZatohcZaKx3tul8t1IeqkWp/EPS4VRXSegxr3dgHJgyC
vEcL1qwis+KObSTgMujY1AiTVZq69QcVE237TdaN54Oktrq4pCr5F4lPMQppXsoE
2XS1ellUKFjZeQL03yq0QdJDOp6NCNsRzEDM0mXUV1LgevUTnswa0RkDx0m5teJd
ZkRWYwd/JZNbu+cdDv8ofpEQILM0dteHhojpFwQKS6LCwol/z7wg1CZ7LG0YWoiJ
L1/Xgu5Rumi66PFhxc/a4eiJ7HR7EA7N+q0r67ystQuIo5MGI01IPleddNvqL0lO
zVtpm5Wh20roSqgiVhOuCCDG4fdbmkfbIYNo1fJF3jA/O7DkVCUAkrClTiif2Vay
2NfeNZS2i/ZucJq/RUt0I5ZUSuiGXs2IsZAdbNRbcxuOqGZjhQc4ao6+8cXHQkcz
8wizSChDdg1OEfI+W4nKIBPks/85L/hcSqQc/UzNFS9OA3BVVAd9w0IrDvPI0WNz
vFrrGfNMC0MYhKGekjPKlzaer2IYzUVaWRfZeXSHTtZGy0O0FWFBJMgvYZnMaDlN
1DWHhHL+rZslaCfwRmiPxjGd8I/Sx3cLBiOqsh8Sfkk0FbhuJZRYHQuNO92fvrev
Lq9eSbprLqLGhGAt0Trgy5NUJ84XDNtrQdYMlGbY4YizAHjNx3URqAAx3BSHT/zC
D5nD1bA0Acc6UcqrCIkETwanspSVhPsaNVrTAj5fDwDfCFshkMnWJvAasNkUx9yj
O4c3/BgtB3djyu5VusKK25xI2twKQuvnu0v85fbf4eaLMFLip8SM/TwWMjN2Mlxl
whjugCfkczB1y91n16AyOeqlHlUCO8CDx3ERoYL6ihMTy6Y/RVfAikzfsdmG89hL
+MMnQZoTMHi7hzymiifHUSVkxzhBMAIvYPaG0lCPGZTAgpMVmjNTMKgBvCuhogYE
+4tpQDcQ4dwuIAEXaTl0QxkxNpkhVwMrJ2fKWxG5xfyvpzTufSyhrc8Cw3yxl7co
FoLvfKGqI7jwvkNso1mmw2GuQHX0XUCOARNZBAC6LeUk5vyuytBFaYq//HlwenNh
RW2UNX3n7pqO/+/k3gwpibsjdm116Lh1mR0mbfoHHzETn2rTxfF7S3oiwtxJ4icG
OpTLH1feiyFqr+f4y3PBro9TgF1jBRpUt99dXAOXkr3UgcN6eXPw4WWZIAOVieDv
rDZIOCr3wlg77v1tyqf99S6NeicNVJD7F/r0O4ylniWEQkaYuibUOEPFMC8MZj++
zXvUEtriDmzwd9dTrejt/8N1MRZU1x/e25oPZsfofMPiDWREEE8o/a+qM7Jpnuic
lPYT648JeEjHSpTHAuJyj2+9E081yNjiI+TwvHcrRj98JNI01ZA9nxB/5MD2w4K5
VQzLtuzVjqddWtHeS5nJ4lUJeKbw7/M9Gj5HbeJglynbi88QAGjCFzgRcoCZPrnc
jlxs6cyUdOe2P/DJhPF5bCDE9DYnJjjdzTtZdBTv/OMoceYo23n2Vre2beAJMEqv
gArYKE5qGWoD8cqjAPWmXWviR36wBbDfCtyY8t8iC66hosOzNuiMnouwHXxFabDp
JsgaT7AeLpzvPLvzxWaDbhbyu6nxf9L6fyETpJl7EcvUgegSJW0wG/iKuC8aHbPA
dSmZRQVtqKJ6dvJeg05XHp85t2gRDJZ/TzTCQGUPc6e6CkgEjv++3ZHvYQaynlv0
PA2HJYjbICFfUn4736E0DFS4Ideh+rEsWdqr4NJEtP0qvjiSt0vViwsCSQleM7Q3
HdPyavJIkgWsF4IOPGVVhRnrjAlLAR0Lol3ShXvzh3rvE9MZuIkz9dzIviTUWrn9
sbPFQAvYpKLzXt2gtdqeRXMasR4kfkPS31vFUdbRSoPXHRKfyTWI1lbSCPLA0Byp
en1UVOlbeSk9k9gRY19jYoWZRVWi5U1a+i26dr6A7X433rt8hokuCvNOOmW/SqZE
9bD659Wo1vumbyrX151UmuoZFjHnQUUczD1PZNXLRsPLRYQYdICuZ4ncIhS/jcyW
uaPbaHTrVFBkMmnkc8qCnB4n/Hg1BFbFQ0LP24s5rhZ7dr5Uk7OATuU+rC0MXDit
OcGlHQmIupew4LBnTOu7nwH5Qhum3I+Yc2/vfjPXxOO4Ac7AxNDgmyVnQ4mQWtf7
+CkqoYirnoyBjaSmXf8G3evafhnEa1Kxxle8egzZwDO9tvkwIcpMpvAt8xvLuM/L
w89yDjRMizhMPj3Fzv+MnyjqErEqY6yV7QdJBPoYAJus+/0vAG3AGtsa1T5x+ye/
bDMxNOoOQ6w6zU8Sn6NZdHKNADaSaRfux4fmnRVUVQ2JUNefbwwyZMFsUWc6Kl7p
LuW1/FHFtNUNuUbj4aGErwWHnGnKN5DAJ0RdsO/re+G1P+zcFJDHIbwitj4IDWUz
LjyA7rjxRa4+gbh39tiRiGHXqiCETCbCkyWyoZxThliCsmw1gaZeG6M2s2uQtj1f
Oe89607K/GSGEaM515Rkb6kpjhvZ5OVn1QUaH6u+Pn+thKGXWYRA5SBdVShM9KzS
nfcK2eXUFWaV/FJu/xtbJjO2myV4abMjSyLtWPDz/vJEnezOCJrycB7Bk/eBr6bu
2YuelL7grew00k9g/NcfJzIF5bzgBE5Jzk/qTIXecpoqEojpwfBT2lRYfP2u1huv
kgrcSOe09whJyxkmSwhhAH1u26xx//kLi+P6I2TnZv4aDUQXVRPE+Ujfb2JgTbyd
T0OJqmnaStjcuQbvPM10a0Tq2Pls675Z/YqyfBfX86YBquwcMtj+jnvRzgI4yi94
XodjWiqcxiGHzHKPIXve1U4/FbDQkkrGFMeDePqMiCEFHHPdynybovGDJRW6zkp2
6jDEDENbEkLIY88bssV5j3w3YnLN+pAztCGRr+V4PpJ7jqK04anoEGEJRPsyNDnU
hlbk0zWx0TAFHjFYQoM3WfyKqoqM+0tTHZF6YL7vWRM1RE14dxKTFYntHsIKI2VZ
G7JwmR1bxhXQO8qPQEP4q9AU4qjNEQiChLZTKJg8vSdlOseVgNiMKuNlAD/uaoyx
KCrUGM03E8qlUk0dGbKQTcjSMC/BII32B+EeExPVrd21iT+Z4Uln2APrJt5L2DdP
NMgAetIRXOSOM6JYEA59DhFFj71MH03OrQL1RmN3DW/ph6C8XrpcfC636hiMgqG2
wrwajx6ptfVmVnxOB5+5W3bBvZJ1FBPXcZhnlh8JtWcan4Cve3TFcXiMr755XyMP
mNKqBlkTqfXgVM7SXvbHYxiuPqncCr30yMdjGJskYku8gq7ENWQfHvOEUHhPBz+O
r6v5xJ1eF/jZngohENlDTzxeqjMzw7Tenp21mtzrqEcyzAurWYcunHxZe4rYWof2
iDP5/z1B+oad7dXAFSu8d0dlv5U4ftRWsSW6b0cbwuM9i4i+gTondLbCEe1S5WsD
rZYsXl5midzOv+6yT501EgYi0stE6rQxoypNab47wKq4FKJJi7/d3hgbhNthCMPp
nEbt7QjDYhFgYj20AUFmJ6RzukR4kiHSEAYGG+o5fdraqWVp4KHOB4JaLbMBDZqj
k6QltcZwOcUD4uvQKakxkajkZApt5iemBhr4iBHsBh3Bn9HUrgC/Ief5OKrc0bxn
JN9H1wfet2o/5szgShOUPvYh5Txhs96497EfVFRH7vyBAoYWV7aOaa3gAkqVrfY0
BHr476Qbpe4caIEmg0Ae1hcxWI2aSpjYfQPAQk2hdN3u9C8HDoxn8rwaCDneu/05
A68ww2oMSPyKyLHYg1Me5JK6L0WRy5uA7YHUozLGPOx5Wma7+nydRC0j6RS4qyoM
h+C1hDtVWNm81jkD8S/fxB5D7s1oM5Ez0CQHYDjFzLnoywZkHv+NvEtZE4/4QR0n
BS/nsmbG7OgU0ocF4NFPJuwKk7SEL/NWj/C8j+cK5vGvZBgALMYuOBlZbL7ypJM1
IJrIM2DgfA6ryt7aeMp1TYunwEfr0zG5hK1eFZM+vzFp6vY0AE4w7dQ7Y6D9dCd0
cdkCza/bu7WehEkqNKxC/iJXBj8oCsNbN5zY5OzTYFGjZNSSj4cCfmvj0JcNWnk3
KNExzW8wRY4E/G9LORjVycz7wLKMD2SfDsuGbRPQ0en1hI+ZlHe8u2F7olWCPYi4
SL3evkRSNPeWcqWtBEQkST7giOLSSEBgVs8EzD3oVadgE4I3+hE3bigI7Z3OOJwl
50ebgmqs6VfrSQcQnoOx8DWyqcbG4lvCzr9sbSv95/kzp7o79PY2mI8o5B7AbGqV
xy3F3j1AzIVFqc3Bf4U3xarm4tLuSG21ah+tCjKm7LonAyE9g/sHyZzQacMiyAUh
XqSq7xahtLGNy8IZpI+wDmnE6e63Ey4blDKsk3exMPA/n48nrX5EVx5Wu64T8riQ
J3UGwVbVDDZCxA8pT3CbJoDoXlW+kediqObKle1CEUmsxs/c8QOGjcMn3zke8nco
EyuaMs2IL+w0GQsK+PArm8Zbu1NPKZl/w8qdN2av0eZdkfjBOrRBbYpn+uAJ2C5P
BL7d6tkHmsZ+HFSTSBBQjD7us9xFpS4Szr8CM1Vpdhv2adNGFsF/jKXBwYMQJAwJ
8YkPjSzHif8zYJlVUvrkDchPoP04ib2Ov7k/wxwZZRCB6gPMq/kcLR47WO6j8e2l
o/oOcHXulfMyApmcoSjqmEs05wECqoQpBpYHl30gevn63RvTJAhmng2p0kZqr+Es
iSNXkuqvV5VdPbKmkDmgKVAri3CA/HDNT4Aw0WDw1uKVJD/jGLRzc58uy5Prl/Za
fui61yf64uGXwOma7BrnEemXL/VPQtAzXSv+5JQp/wq8iYRUDpUhX02krYdfM0i4
t0ougJthEhz77UIBmWsXTxuq/RfaYz5QWkSvRFTf6d+HdKP4MfeqKySepvBo7OMb
fGdgREHiM0vOpz5Ci2li1D0vD5L3O7XPZii2/5mIoZo9vFZNTMIH8kY9W2XFvs84
J2hIy0Twl284r/QpF7XnHWaf08U97Hx668X3LQW4mNyFpokPPDRn1krZ1ngZpsV0
pRM7PylMyRnsNQ/KDwW8/PIEVylYdWsk8QADvJZm51K6bpkr3cSiPon3OcvxK0aS
p5jLFrFnTmDgzT4rhH5v4ptc3M3dzRogYKMZh21PI02kGT6V06EJRuyjp1LkC/rd
LrFNFNxon8CeOYOgoSXbaQPgXAw6UJnw93DibzFgfVCO8rcWBXc9Iu9BkNgBxJ/o
CK+1/K/aYYa5CikvfCjKAD6HWod6237Mt+7gDuL/nT23lfwO6o+NUGjEL9svUh6a
Wzf72T+1Hv4qvSCxfw5KlGYYg2RkIOY0FVV0u9QKUvhhnbF8Rsa1sJTPm/Ir5z0c
Muhuc0lIQ2qwrPiDyeSx2VXy+nVJV6hTGZP0lcKQ6jX1HNMMevXA5J/iTMUQzagC
T90wMfp93YPH8n8z1dzKq57VMiZCzNd1USi8kbb1XEtxdHrVggcgd5/c1vzfHcw3
Ic5ElXRciLBMBq/bY9egFoLhdHxSYMK8uZ4XfeVZ6IgGKctD8RejHOzCE5kI9pNP
bULJKtXw83vkF1L0OrgKTLWwF2yMtOjE7GdTrwyouzb2Bp0ZToqUKhZc951/QMHK
s4JdDZ45H1lpJjCfiJBglTRwMs6WXLWMeC4JIg3Tl2ScofzvpZDAUkKIlUzwu/ih
4/074Gko2oy5L2tCuvx9SQstYAXvRh0MtrtihD/XK41tDOj+74sIi+bKDqNMcj/A
s+jftMHdmJYYjdZSTNeVI/rrkjIfXa3V/3ed2O9WW0/Jta5MiAIdlyz95RH572DA
R7PRVLg/fUiVR65mXXsJVukO0lWElzCuoejbtopIBmqwbqA5XtmRUrgNEFX5APxu
J5Z4YmmbGPrxTqeWiJcDn/Qi+ojN+AH+RNSv7Vxt8kEgzChstZW/zG0bAkdhg9RX
HKT8/6TS8nGQ6lkz5VsDfTqqJ6OCIBPXUEQlYevHyT29zue/gOGjcUif/KA6R6Ph
5kgQxqq5Cb4j/azUdZoZbwjjLsQTekgm5f+I5CfckdmiQiGRmg6OKonGTIhgZEe1
ho30gWZ0PckdeK+GbhWp2idPe93BNa99wcvUNOLY7/ij0H2dgnct+pMM8z1Nakhz
MvEfzVaYqroDM+2EWk+cANn3ec32pmEKzBX9SN9p1PAlB3dAnhNNbmMIplJeVSp+
743O2u/bKloFAsdyOekxqHJJRLlgkrS4vk2TkRlSI9gruFdy+vh06Fvd28RGwADv
g2vYPY/BfnYmxr4U/tGXIC0ouPJADA2E5eQDlEPzldDIOtHU6X4b9x0dRNLRB75g
YY82uflikyUnSZC3MErjUPJIRSXfAJbZxDqh/tjwQQI636bIJZ+sTyO5YRPkHWMf
aZoUiwwB2+dAfQxYGXq2poLet6bz+mKDpwbIJCO8PsY2pns3elfTvcq5HK+Pa8QO
tXMgDzInHLtoqgf/9VCSmX8JDZtY5bfrmOU2mNFPuCTgczIV5oF/w8+wFLARfJy3
YcVY6MYvshgYYm82VvXnE+50p3mdxcPrXNNY/XlB08GtlUPgJlhlMrQwoCRKSv+B
aJYyxDu3IxjY2QPb5kVyg8DF4J4ew2iBNBR2y4O17E5MjCpW/imf5phV/1863frW
Xt453h62nU+HgI5MZjYVaoqTTe8pU2oQkAGY/T+cH2QBrD9M8xuP42HaK3dQItRP
bsrR3+USQlZD6QGUEO4C0d5AnxsbhJ1Z17GhVmXjiiqCnfVwmf34CPW1bY75vsMn
ikq4zSyMVgIS7MSfX9H5gkw3v9MEKwdD2zyrv9GWkteDx34yFS2KvXV3sVZcs6o4
kGucDeWwS5t8LHUCvpx7iGR7oDFOglFnQkK+kgYNaAq8Lat5+WG61HsZxXs0xfNf
n4j51n90JcMLxDIl/jSFmm3TlPNox/Ka9BHMk46UmK6Nwgv8C7Uf2deYpXCcJvDn
4Kut2AZTnrrf15AYdwjwYfhg9Ow7wFxRLMj51hLceL4XRnVrccATukweLJT3QeDh
3DZcYYn5ZGKxkWBzyZvlb2hs2P5huSJqcr5Int4GV1bd646aBNoYzqggVVE7Vh1P
+cazx4A8M0SOn2joeSOq9SrOBioWQqcYlTBELqS3xD4DolvR5jJ5lbPmttcLSWi/
JDGwN5zWPHtqvc3xUuT2WU2BKA6Fk5rTl7F25inv02aT1NqGOWm7AFszBHw5dsC1
wnn6V+J0Ktknr8A/v9QCdI++RYIRBl+RQJwNsIASBR7bJiIHyyQYJWUG7+FavD9D
D1I8+MTxDlMUyTW2aXvSFoi9lgI13RJ/PBPx/ZE6xY5vyllgEnNljJfnQUevfzRq
a7OaZrKKb99ZDBcttQ1BrawnImrUVXAE1CAvt9EkYmxlh7WSgCWHWhDBGY238BN3
JVIADB4eKl2l7e4KnB3CKOya0VcdNTgYwz8ZCC2SAisoiwlsU8S9sUUcuiy4zMV9
gThTXeP5m8sg9pKaMXAeEpE+RahLm1aPzEqtb+Bor+f/BjZgK5cOp5yFpyGSVB/C
6b6cso79L7isl5iao6g7oAO/WjHuoJB5m7UNoa18ZDcNxR+GEpQhxi906Kc/9+hT
2i4m//g40elZVSMh33aaoJMeImU9MqMCEq5V0IlyX3YFDzA2vhn+8WRlwWaBgBeN
MR5sS1rstYrtuUFYeC4UMSZ8xNqjhqCgW/+Gg+4ybLPXukhoVaMuBh9hdORzYtq5
V9ZbjUEL5ibAekB7DkY2Wc6plR+hpnDZpvxM2Zy4mTaavobj2xYPQeD6d2fqA7fC
X0Qr2xNoh5abJD+HvGCWnNYGPV0HAAP2DWAoWVV04pNazoHmpETJWhfkv443iCR4
BWzxO5l9FQN54heBe9jJwGdI8m4aPtZV9HDFBCw3k8DdzcGQoWbtfDBrQLOZ+rrx
CwBDEX0iUAus88sRMWTArLKCso0W+DzlBgFuQpds6KZOQNmi8wYtG7SN54/4uULU
SyBvb2R2zTH37Aqox4bCB7ndBPnBxmUsjV3biD0/vxEfB3IR8KzDIZeYSArBBk8Y
Km+MM2ixUwjgu7idCOowZAy/L2qeYVE2dY5vQA6abz3S0foNCcob7V7NPZbwvgbx
rE9s796406my1Um59mMATTqIuPK17wiXy/+abxkhFlJvLYP3LDd+aP+7L15Wf11c
LR8hxklElrgkoEnSrFYntZ9R9UP3AYjtlHZjIlM7T5IfpwBKgQLMtC/iHbJA+Oo0
tpzGtA1nDbJ9bY4JajxXBP2t7GIEP/6QkEmgG5tu058OGnxY81e2DqQTCFuUAZ9y
qiaKyTfRN5AYE2PI/hOrk+nibyRw1RpMsYael86o/ENgK0KzKCgVZs+7zFcBHd70
5/oo7b+HeBQTQEA3qni0+Spsa1quNSRWAw4TtGwF9tNPGNikDkS3kEvD+6zEWmaR
OwPywiwvgqELTXcGDwsWTnnjm+e3rNeLfwX0vfWydzp5lpAdfexmRU/1CMh2ZZZL
pDb6OSJdPnziIAGF8wHoD7IGI8nIMIIVPVYzCH9zmvtYZonGfzFJEwAaUN95GvKN
NzI91JLvnpaJdkZzXuk8QEXiX5siCxMQbyln6ktXXGMHfFV8YPMm/1Z4aRZP+OP/
7MHJmBAoO3YSipz5nygJ3HFy96iDK9mqG3NdLrjH50lh8CDUjpkzTDvD5LaZK31C
y3+63UWCjEnI0Mjy85qukqtJXpUE/oA8hrv3iYsaXPu+8CRycSfBMFvXV1jeyLV8
GEXDgoJ+qbeGJi8LHlLE0XCkhG7e+j9LaF01oTtPRNqy+ocaZ1raEWw4GaZW6MAT
1M4dy50D+xpFafAyWvcAgbU8lDcFg1ZjRYBkXdrbXxBcAQ4LoQJFhw4VMXHqMrTZ
Vshfkr9SY6sqbvBzLzVzIor+4bkdYmt5QD783N4MNw7myoSmf5gQOPfU7MWzZiud
bFSVKYqTyfmKicOOSIG3TKmw+kbcR8awmtPprHYSGVvVuZErNXdlDPRTC6t9AVKG
y0k/UMIYbqGsnCbUkQREV0H9+tzVstLjPiD+dJ0Y90zNRwy9C+n2pjCqlZ0nYMxF
ADjJSYYqr5d7hkyYRYZ7RFI6wBeyiaquW7+Xs1gXWLdenj4c3Rsy7a8KusRiXg6q
Xev+cN4yhXrprAtOwBmzuqS7MFX17NVHV/yZYMuMHdlVaixUH3Cu3Q+yBjvZu3xR
tV3E3bGaS2wnNq8tO7w3f0MKxSZVv0o3qy+1dLmEh0nNd3r6Cpz9q3S1PL9X1Wu5
OuR0+/henoI+uGqY/4omsnDoG6kRyHiXig/NHGkHGf2P0BevAqNI+rafo0bwEcty
7K28KYY2JAAlY4OBmSWUUNMAlON+m+QhtrqjFjAks6s/ijpAxeli2isB1XP/LKT6
kOluBESDAbmdvryyi0Xno8R5nzY2b8b027coC1oWbi2Sx8Rscpge5JjPL5ClFcLY
s5SSFdiXH3QPcV4EyQGKRsLdViFAhVYQRfJnD1ULLYF1u3nFpM+wAlGr33B1aJ6p
DtbUtybcgPvicxsmRE0XNTXM5cfqXrqmogomO5HztHW7oI9Irah77XWeAvg43VMv
MMGgWjiARH+dMQXR+QmHd/5tw/ZhYbN71DzkGnEplNlCZzoumoN56eQ7Lhiqq+7t
NRss8KMjSovW+EqHCr3bk9vksfq0MxGa0UKyHduW0lvbiE/esF7l6LHsDtAmqVTd
SnQXqwZRdKKhmKeHYQo4q5PkXb68iroaOJ2iA21ncaPEU/1fNOJSOg9MfwB/ekLU
4r6nrGn2SG/ZVq+cYEvIIXO1ZR2piK0leMeSA/a1AGlk22f4rqSmF+lx769tIVZy
C4aOUkxmKIwduO/uWSNgNTHwwW33rmYiQXU1tuuO8wUNnfSBClaBVInyHxFXekYn
UUHBLGqWVl7LwfanwGDRdSUI0YJpns9a1w+IQ+YxtrbkspBp+siMXHIZgMAmB2YR
3KYLCzEw4ZN/xi8G6QGoq/y5RZ2haXOvNlyNfxD89G8nzplzdZcqLPYvijNEhYaG
gXuFr+iC97TRR1H9+0VDYv/g/9q0YuVE4oP+pYhfVb2eCEHCSgYyATrl/m8IkFm2
0bOiw7NHo4J5+ExR9fNKBh0Rz7K3swhaBXE+tCq/Gj7Mx30A0tkyKrEZ6pKQ0tTw
5+Xg9AUWEZkNP+LptHZeY7vpNiNKLYOWAtOK391jHi7bxgsPo1aY2Fcd6YinwN1d
k0VDsuKM2rjoOWt8D8ckYvuEOzI4Q4AbQI6+XiPDkndvuY4xGQ03yXx1ZVKTP4L2
kmvWVCDoSd1WQbFDC63w5ujwd2/QglPhKdZa3D+wtIT2gOLBAnRE3BAS634niJot
b/LJLgcyDgGYSHMx8vTOE8IDyeW/V5XgfNQ7m6WLeP2q/YObvEp+3YYDuYR5DUKa
dATMVoL40wR7FCxyrJfWRdCvXoqyyKD0a9aKbl7To/3Chz3Abj+tvE0vTlvHP4Ad
wTi3uuqGfX/r8UTmJ4mT2OgYbFrQSjPWJ69b1c03B1n0cvgxmnhndsfb4z1asVz/
c0V8m28+/ly/owNw977SejwGTo5JsosFgAkqZvprddiifRTAF3zGxy5NJlvs6c0v
HzBXhJ/rI2/wHomIng14ULAeNKgsyV1rysmRbvralpMTKU2M1Cn3h6Z8qofVCPMd
B+8q0H/y9myLfbHhFZnpZS3sG8CkLYJ7i39PDXuAnjJBKm4hwkV6/ndWTY++6caM
Ha89+TQfN9bem8WCviexFkGNMX8k+f4ZJe87/ZNxLYXIuvqCHC9/lHVdIE9M0djG
L7BdW//DzBzHxAeY2FdDeUP/z5WzSVs7DphFszaN+wSPCv30noj43Zx1mE1zRhm5
BZsUE23qtCwqhSV7wp7QxRYvINJES1NFMxBGgoamoE9y8kd/SOBYVQvD0faYtPG5
+A8CpZfda601BfdOurOoXbBPd/eMqdD4iRvKrjaKwRkzvwqXeKgK08aikAsjT/wz
vz2om7g3G/+1PeU4a5hFB/yQ22BENCP0qeUqzr/5Ne6SdHb+zg/RqWpqTk0WyKJ7
rddVcKVZXeZS35D8P2tyTKLvnR6WGui5M0OIsqcUsx+xCcJCfMEcY6y0XNDWTqoi
FGSUPwOYWl7KQzgq4pz26uZS+bbkOhRpeNj3WPOQqc47flJttZT72N2KJ+AUoXKJ
e0zT/pYwhBIzTMDpyWD/OehYABBLkZKaM0kVbWNJdDcKUY76nr//FwGqz2IDD/Bk
E0hPCzqqSSgt9tpHSsPEf0lhRVbS/HQu1g7N0MXgRhJR8f8PrifSOy4XNmSqpmm6
5tlWGC46ulKjx38sHB5ltzbDmF9DLgaZOhezFGjkTXUDhu4/w4Jnb575N4d9pS6w
aUYBbdMpX5xEkZ3Bd0+6+GmfAeq53WYr3n2Q4bF1tI3UV+lriV78yMZTYFC8+I3h
uwO33XgGS5oXJ85hRSXg/VMBjUTM+7XrZwHpaLS2JqV9IvdvXpEGKRdMOmpfpoEx
jfxqZQDe2Cy+Z87A7D1iKduZrzjykjvrBhNc1lkm52rHVpYkjXpcbyDWjhcb7mPF
8llFWoNH70b7vQUHDqBcdeVDNe9EbaILVjrvAlbwRp+O5PbE2lEHH/6CpzN5f1iw
6uhq5Cc7VPdOnOp/aEQAq9ixVmkEdiK2y+e2a0Zb66tKegxkAB2ok140j5NKS7zZ
GskS0yM/OqLFvriibAHTq5swaztytx4KcDmPpmV4FVkUlSR4NKJVhml1D+uxsbNA
WRcs53mI8o96vHmaHq4ezR6eE0NZ82ZKm9mYBiJuXN5x7fXxv+kGj8qQULCkkFFx
jHqs5RD8yHJC6rswSL/atLrcbCAjet0nNdnwjBHkd7OkfjI+43eH+hD0fENWL5v1
SaH63Oh/Qo3sPfn7Nc6aUPqoavemM9juW74lqM3hmJb9ZVjAcBV69NI3zzWkVTeO
4mgtSo63gGdlT2MsrTTyToXvE7yiARtyi66+Ekw17TdRAjA262SjkYw35Hb8XLVW
UXUl0B4RTkCewx6zB7+TnU0JuByEfvxq3QeM+bawn0NjhkqW7bO2siTpKvp2HBTw
XBye4wyxyJqFGW1sQl6+IXsHBqkS1YA6f/xh70NZQYngrnbRoB9v1UPO5+epnk3g
neKQt/BmTfHcpQ8qtjusNEoaXNmGK3W98tCQmRumPZoGY44kkAKT1inrHRJJOJjx
X7gmFhUhUHiCZBGvJvL2viGLKRk67cmaBr7fI/0Rh/JrnaYzK7lrbUv7CiWWq19i
c76wOHdZMPWnLly36eIEATqkIv1jZQDpialxMvz671RK4Uv8W9Roh53kT5eRncYQ
jZaBIwJOkgl1VX4/KuzhDqJr/hOCz1Q87xhW8Wtv5NZt9Ifm7fF9G90kxGqtN8Gj
i5fJD5kmLi1W7p6x3shZaU+2A/M01WftJwdezrhi8Sl/N89MGPzEYFIVUy5Vx1u1
9rBi1EDpujZ1meNJ+i9Alddv7tZqKQO3dQP28mO00lRxivJIHfz2l+eAZJeqjehH
PriegP8j3XOlvHjVimza83iP0BXX7Amt4GinmvsNXf92c7T3zz4QnB0Sfsi9witI
hiuczWm7SObzfiEuBWhuk47VokCHGzr7D8aWT2VkfbTfCIh6oNNbY0T1m4xuHD57
dRZURg0RxiVJZgflYHO/cvRtLhtTD660dJE6ZiUoy3BL3O75KzBJsxujyj7V9R6u
4wxLKhQFf/j/4W1yKjnvImGj3s7ivzk8AORBRSx8tgAQxJtr8/c90ZEllkjjJ5ti
erZoHnzN0DAKfNgs9BsHlNCom1kF9kqhc3iCE0X5ZmaayMka+Lqbb6KbwOCU6buv
kaNkR7C6LpejOPHD5lelFHw5MerIZnY/z30dsw7QWjSSvPaweJmCT8mPWtQMEWaW
ru64kpXf5yJ3Ttzq+oR/p3KWgvb/NKuW9iOYbyGcmut/7gWtVLhObLsp4iTpaODp
AV4LBEx7R8kh1Yc8fZEhwr8FXqEPm4ccZMDgjRGPbHyGSKCHYr9o75r5B05Hrxec
yonJtSFMk85dst21S18f2wt8Zx8pIiwmXtVR603jl9OneoJpbx8o3HlExY7NBe6w
UE7xY2P5eZonhxTnkmW41c/mq+vT3bnLpE+ZPHKVlnDEcIQwxcvoF3dN6r/yYuDP
SuWVuRns1EC/EL/I4tfTydWj5S8Ko1lyyW4dzQSZnWzNkLDX7EGQVb5it4dieoTt
SkG+s9AO4JQ3IphDc7MbJZ6xPlbLzGP+KeUDNAuJOLxvYvYm3dXv7op0kenc+NOP
mDlIf/fXzaZ4RO27UD7THDSpg0LdmCDnxQLc+BNiohAoAuCPV/N4GM/IcWBrIT1L
/BlpAJECaXK8sD39JCahTEzuOkDzBh6SXHEm42GZ9HL34pFnH13mFOHjlFGTr/UG
82ci5oOJPSOnQCffi3WHavKo2TUx+yyuR6Kavq6D2v2+ZhqwpOeotXwXPfQ/ZLTB
2QGOBvBPhagHXRQhqwmPiM0JStWhKpaPaCNPHAuwwConauv0lYOv5FurYw0+UoeW
e9/HwM5s973iSeDG3B3E3/LOEiJLMER/PXPUboK2JEW1e94ABJkNWvDi81sqVeWz
IGBBELz/4eTIsH1x1zZySrMMvIQu264e0Gr/vpvpd691dG0L63+UQe9NLFsr2hUw
oVrIGXry/FTATQ/vUthirLrGeRUyyu8ukZTCnCSR9UgmjE8wmoMCCJfGUv8mJcur
awmGlXZj2PJdSGQlSBi0csPryQPMF04HD2hULIC3mmXhZrwzwBBBcvBppb4ats5p
CA/ygvw7M8vLGhPElOoYUDm2KnKo0GMduNNXoeivkXcp7wRf5gPvGt+LSaYYiXkZ
/K+OM0sgvUximXoyQLA24fYNMqdqAGsJo9T8Nlls4cT4Tv1v+gJ/Ue+N96IMpjDv
aRD575pbdPIs68CnKZ1sQkIjD2PuxIhm/1m7coe3sqp3NvBpAhHf5SWd9oG38voW
sMW56WB83CIxCIvWQIyn7KpfUjL7ml3KhSLx+FlXjQrOJ6hOKCHeoTIXlSNgB2Lk
KhoM7ZHI18fMKNpyMuQexogas79m3YHZu8qyeSXU+3UE+fr/kKRXzABtVEs/tDoS
Xu9ShZ7P+5u+9xah8Z+HW4qMkax5tPS6lVMdtRt6m3ASvBB5MsBLdpsbTTmpOPlE
T2hluoASz4O/rzGDRy/XLwqX39DVFkPy8dM/FXmUn5Ow8e63rowMtsWO9bKx6jo1
6oCnEQUVrA/0yIXCRGIJPet1xbAW0oMU3AC5M3CdSx4dcY31fzKE/Q0ky9NJGLlT
gb/p1ukkfTsEEIJDM1dO3aPsNHaLR2V+ABnFK3lU4op3U2prrTOK3+E1ksl5/XdD
M9Zj3hS0pmZ3iT2iW7U1sG0ShnfxFQ3u3uts2aVxPzAZ7HRZLbsSNHchXrE1THCn
nybrC4KF4i8XTLGIPBMJe7x0Aovc5GFIkVZ3ZzR8PTDPbHb2XTYwERnkG89tSb1h
PfDEMcVmOY6WQzIAN7RjBIz5W50D81VpGh5CypXDwqEzOtGl4/MM8LH+dHbWQ1je
Czshh/WvKWUUv7QRjjkz6g97Crxzwe45Mrrxqn13GQueYQEYknrytcGQs1xB/swy
qj2UAgRxeb2G0Cp5xDAAqLVbZP5d/W90V7fPF4FEZedgcJy4KA++ZI4e2uZSlKth
K2hlhD1apDOUc0Nkm09TQTIQBKI6enxjpA1M2crFvbuKyMZRigPSBeueWBKzcuv0
kuqH6Mvs23JJhR4S5b3e+8/BJ6g5AKzGzTySAV+1FIP7sGnoBjWL9VGZvJQwA6on
mgOAe9Zwiza/5Cah+n+DBZfAyJVxGY7yZ3fepkumm6ovbqpd3/jJg5jVKS0QKdpY
Zw4GQkCXqJJKmNODdMYDOv5PDwWQSbJoQzycW4VLapWduFzECpo+DH4rYzWtRkkq
KmBQlK0Av4qU6aS7IJ+m6M7OehknILjmqKjfP1HjnSL+46Gw1migsIu2msxK3Zxm
CjNcLn+BEKszoktwUfj4k7FBvmrgtnDzSRqATaCyhvL2EDhztZaRRbrzyc5mjlr/
DwFOfK0qC0KfTdo1NEOhVlAWxoAszy818uLKdB2baS2vNMM7QJZQpWsnoshPbT8d
YIleGNfb//r1wHtw1Uj6/5OrZRrJsPkY8AGkz3/JoTwxeN/43c8Tv3WBNEM32Bcx
Xtonf4Yr5XGSqtvDtB4hbW+vEIbCtGTIL+a4uFcVRNHoPbeF2P/yKjZNeGslixfn
kgFXAdKADhh+icJFg5nc/fCsJHMWdaSxsA87P1sAqk1LswwLSmFS6dx/mV2XcoDj
mPbRAK+Y+Tsqn0UJXcicIY0pltNbpvWePsc1O0LdV4+tnPVaINwfEBydzMQk6hlj
tHfXlpv/3HWGquzjzM8hX4Kn+oVgBu9Vd+74pe5a4ymqXxbhKrl16FOYy+P7oa/4
xm2IEzEMfbkw0o9Kw18KsvFS8nM7qKKWi0hsUbTbHqagX8B+oQ9GgNwiK0iZZ4Ut
9fI78q7ECIm/m+4YXA7eVH1zYbPseeywFtlFDMBDpWHnKFzAv9u+rXjmeaJ6ATGx
0Bs7gX4i4pfxh/xcq5bpLde5MaqE5gjP/gAqHUGVy4/hT42sblfWQsQJzKp0eMZy
H69lIPU/aTVBg1U45QfQlOgp46+zUlm+hSbAKllqkyStbv7SbWodp8/021xgOwSO
wsAL130rXimEt2FvyVomnAManiQfTntOAysiPheKU3tJ4Wvo8q5Qs+dxh5Uz5GKl
Gy4/mXwVvo12JvbZIJ8gxCHW4muwm2gGfbR3p9O3iYgDdRj4aZOmWKFWJgiq+kAR
0Z/msHQiQv+BlDNi2LZCjNC+SPNkjWkXyBAl4SfyHysslWk8Vhl2yLnadkXKDC4Q
g5Y5ahuNEtxyaIfKRQ8iAMi+8Zfc4BhIxPlCJjWwGGqlaGM6NhEeu0QMbyzbOABT
+h6NBDN6oo02zsyXOcSGRmabuSpSu+UH2ezAFt5XhzPB56KLe5oaQN2NJuXkrEIO
0JWHOOv4jIpI3FcV/Qg6L9iSB5ax0uIRSQ5Prx6PugBJyQXgzZGIwet9tj+zosOF
4J1PDUDCs0Zuh6G6foDeuIuRo3/CbzPIvVCEGC9QMQMjexic7CGW6wrb6WwUAIhI
mrb1cC8RYxqkN7eknu1MhHh8lqtcPwKsjHR1toq/eyzbUtQKvEzOjV8usEjKRm/m
iAsiy7nv7G5eRLO+aWVBON9/zcSJuRDHic/oLQS+86fU7JPn+aYpid+EMbjrv6sf
WoW6qXaqgaPL4gklUdnsn3PwzGQOMD9TSr9ZRuctSG4AZCy0AyGQlxccthnGhsB+
bxBzxzHXHgcqOf5mYncf/S0gJzgdCcVIbQrXadXAbCPNKg76v2HDJCt67ZBGCy19
cKWqkn25eDgoq9enpvKATUqi0hUi3tJrI2xdDsQsVUjX4zGreYekoWJ8yoid1iN1
MPUXJvSKeqVYjAAQ5Pzkja5Q+mHbHhTaMgD+IkZc/9hBvNpIMswRBA6SJ/Kp27Yj
xFSHC/6oq+ueyx8l44SMY8ci4bO3X2G6v/kY1tKsGTdCBlSc5vgf9OcJyNd/HY+k
PXBzbTcRdl7hu8ZbGiGmtcY8tEsWS82FA38WthNjtWGouYR4t/4xEVvXB+1W0OEQ
//PpNIHJWaTX/Hme+b7McvaAhi2U9T21AHeZheCKBzd+sMuO9aGIhf1USpJztLeS
3HIm6kCwb9GnQ6OGWQ0Ecl7Oj6+UG1uLe1W4JkmWGIEmcFVFvcsq5bkUn3q5XJZD
nan9lFytidKJ/+9dI0BL+zWaIrfSEx9f8C6drVYzgh+gHo/HPfCZ4/kWas/kaT8N
yAcnORApOorqAPZKvWEdRHl8XCI98Llg4WFzhyEBvHtb0boGHun6cXdOEzyHogzW
+cT+6gH6c3QPI+K1oQjMtUct5SkozbR2MtrYoMrkh7u7Z5fUyBjSCPgc4IhchCh0
A3eqLQsjCPG9xminhKECPK0NRkJijUSf/5jYchdUU/pvvHMap1b/XFPI/VHTqDje
sC/ug4lQsUhRn1CKLZrkbIMLX/eaux3PMWAtOrGr6NqMpJQEIbO9t1gkd+s6pHO1
QdlJ1781GR2v63JSaOznCAGerkxjFlVA/sWGtJUQH48wGQDTLjtlRxavxCT6zWmD
deqIOZ4a18cJ7ZH8iLlsB31A4PzizTf4+1GusB9Vlj6SwAzgYWDwY9ZxZDrAD2h0
PuLdUugPvxAfpTromaeZpOMYs7Kn5JxUhPcdZOMdlT6Tq52kyCBTELeBWBUHzGFu
s5nRgWSvphQ1B3fXsGLFnXgV7UEOVCM+b3ploM+nCf3OE6XUJOLmFGwwouafCNge
JBkEi+0e/GkbLHNjTZ/WzfEv+8DfX5YhOUA72BDxOWTp8vnjN2wSsMnNF1j7+Ca6
Rqkr0VPVM6ODPwrEUFXw1MoOf4+B+sVO2Csfl83gYdJSxc1A9iirRdlsJUabeN/9
3qE2JjlOwbUxaCPrO2ND1lbmg38CHoHv1anwU9AQ5yEi9MAanNiQ6M8kS74Bgvyg
8etSx9zfizx0YEg5M5jCg/As+MMVAEvV8YouYS8j8Zw7K2IDnZWS13Tv6nepewcy
srC2yFQvK7N/Tf3hy5b1djS7vv8my6Oz+jxv1hYRSQiISZxo3zQH19znTIOZNfRs
A+e5+UWTqZlonhNDM/YM74hZ3TIxOlF3ljeA+PMKWmHz0HrAtUiW312mpMYY0orf
hQC7hF75blbz0+FhAgQzTUTNt8rOMEaSntSP2hvUIgjlHhVrokuSC2ktP4BpAzjw
TKeMQHBOFw06Yk3u1lnwhqhRCB/dnCDFaC46IXw7WfbqkHnK/wQzU0Huxnaki6Nz
GWLpq1og7P+wYUMLXqz98qt9cIP5SEpm87b5rA6phlsO05hOUrYydHEbIbUNnmZ8
GpQtzbFX2psp/RzjHbbfjCE5rYsR4AxRuHUoJxSimbShVbXKyTxHRryDsHekgZEc
kSfyUCIFDRwWFdXdfo6eOcIf4n9RJNyT+ZAkiXXSxTzxquBf4heaJHqKUFGHQnph
gvwoEnBqa6QYBM9rRgRMjpiBeLdgXdkz8k+feEzQpAZyA0I45XZVmE8QPRaBn3kc
qEK0L7i9FQR8Q5RXTealBaeSHPmNwVCTQbnT/jBnuZLBiKbgfaTiUawqYrMnY6Sp
kJpB+BBITz1mv+H/7yBSTB5VIyBkBJSrDouTNlA1yfM1kgVP875uGS+G8LAM2nmQ
CHUEdkytFJSrFQUThXeycCbyvm2ISl1te7YF2tkqPpqc9UFLR1m/S/KIayTixrEO
t+D1ucNInHcG9haZiQaovdnbzKDUsn+uPFpyA6GjhB3pRggr0AbFuH2pG2DCWvWE
Kls5VYq0PFgXInB+4g9Ghvw/5ChkOew26sh1NtmWd1/f6IgPKbmCD5Fw8PLy9hLu
rQ//qe5y0lBZwZ8YazmUBkZJ8V7urwVG5UKdSFpmlp9HDnrCI/REKyqg6WjyXFSh
Khr5uDMuyXqEtcbp7DsfhgYHUTJNP8CGGvea4NdG9d76SowE0mz353jIh69y/+CZ
Y063Gac/wUZXjr91UG8J4HBCVNDNHlPoVWV/2RbfdSSkk+Iqj7duE/Aql0gSidXw
pCMYfB//k8WgDJ+LUGpno4by5OzYdGHIKVzMrAuTQxoA74LqBjyQRPJk6aKOnSUv
JIIu0A25cvN++0BD1zrjBRJfPZmu8UM/4jS0RFrHF3vvEtrcl4qjbwTUUbZ+m1DZ
ngEXVbUxmgDWQoupY21enAhQvNROv+gj060eFAm0/TClIX7u9DILQhQVUrQmpXe/
n2k9kTA2hI4v77uF57X1B/bPF1CTZGf3WIdS3i6BKXmYln6UehJc99GPTJi3Gp1J
6BtzYPREvsFsR1xKM874ALlTcGtRaGymNqFc6Fmbmzg/ucOegDQQe18y/0mFqHcf
QvCyntzyzUdMvgyipMl7H5TwtaIsCowxv3XY3x+6AnV9JNc+l1AJ/CCsQre8RfhP
JjvZapLWuggMwak5i9qKBQd6uPKC4bqzVVsL3X6tvootwyzfuJv9F5OZ88Mm+o08
3TiYk9ULO8g5b6LUefROLXF9yNzJgNpz0iOd9gqIN7XRQXDW9FurdvyvWv091edt
QBhRk+D6NpotN/YqwDpYkXPn7dzFcocZM2c+OK+2DaxPNBE4CjMRbvCw2QTsl5TH
XRmiGwgGU81nAVsjEeSjkDBVEbPVUmk/yN3mOw2JpdxcGoegNnyskCu4ujgPX96m
OnSv3ZkFvRxQjr7/SWj4tYq9kTK8FHTpsNfzqasv5RfN+m8ATVnOO5YFxqAyvjea
eh6U76mM4D+M0hGuN4rv3U110I+jW5JH1zJJsd8PdMvMiXilfCBctMNh1YYORUL2
nkkUdhsYGCJb6uE+94vzJHXCAi1ES/mhWe6v60l+IJlcKOTgEkxN/W8ojB3TQGbC
sMYrxY3ZMfCMyHU9BYI2HGraGag3J2z1sadZ6bPMAvW7qR2IBjsmQ+agXFVE4uYH
O3atOdSZmUeTjMMt/PVp7+5NlGgPF+6XARx6vWPucq1KzE7Y8QW49mmG5BYs4fQ2
1tLhPlqHHz18nUyhnreRhMWloLHma73OGZMPGbqOH98BeSYteORU1NhSeWH5C9m2
dWPJLVMfx1Etq6gkzDenuTOaXrhbZtCNKdRpOf7Vceed8O02geEWJDrLMv1v/rpb
QxPdQ8eRcRL/z5NOKQf9kKtkXw7Y7fGr6WvzejwiACE5stIi4KIJXk99nClZ0E8h
4+/P8iXOM1pyiuqNBVq3PDvp4UuhkSYjGXE4PlXacRATMxXFp9jqqb9TiC+YwSiU
kFqo8em9kOqiNG3tR4lNer4f3yUBExgEBeIXFqWZULXFVBoCa9EtfBpKdThRo9gZ
OHkFlc6Ly1zxDu4A2tzht5q0uEZAFP0qNkYe8WprP0bzxINlVifZpEQHeD3I1cwU
1J1ICUi1CgK2+UuwwWpgKyR1Ywfx4kBjN5xdaHVFt97ftd0UbiA6qHjrW1j6Xdjs
+3MIrtwX8Nv+QJLtK9M/bNi6SuCqeun2b4EhNWVxqFhxANtM39QVFL76LSDN2Bbi
p4AQmw/qIxHH0d/0sy8TlwVLgBKDYud+KYTGkezbKx59/hWHXu+azyLMZnoIVsE7
6fF3d/rt7Qc4N7/UbAkt99PSiKnNNHV1g8wVvncLjt6cWbyoxf+MEJ0x6pFJ/9h7
LjrU3U8lMMaMfXSIP0DWvLUEVX9YBqU930C6KXXvQq7AxSiQW7lEztjeKZZoR/CX
SXTgGj2ltr6Qj66xmfq3rBBEeB110Na1txJ+cntANH+sNTkz5MWvpHv/EDHCPNen
dQKet2jLnH6e2zA/4W4P/qvCqQdtgf1Mn0K6DHIt5I9+rDWixnqby7Pp0uq8N6mX
gXht//CA/a8BLE1JMXWL7XGOARU3ZYp4dh7mVAsKv/4rcapahdTHAvXPxLI7CIHL
4TIiqvEUN/Wzjv8WjyBpylawz2A92uZGPb2T0+MUmOBw25RnejWywUlyeEODLcSG
S9pak11En9KGlWkef09NDPdUiHiIzqAa9jDLhfYrRphANBy7yOm2quEzhrqKuhQa
FzOCXaa/XBsvjTuJHro+7htUg5mHzDsrTYIedpi8oO5tWy9mvfXGgC1QcUxx56qJ
bjXId0kh4Yy/lR21XQFBACFvCq7kH8RYjKPxEV0TOlh3JXdtAIwMHogjGY5mvDTx
bYWmWMqwjbfdk5G4VyIcrJGbZ2hMB5VXIrgY1F+YKb1CV4kAjlWST+6ZdH2upszO
QZiBmgJD3KxJr/SksDrfDr1OeFn8jG9uZBYZLtvj2qZabSU8O+tpRdYf8rB4dKYV
O//Y6lhYbEpyaYMrXgP4eBM7XaWoBNCkn338CXWpXqe9fHrTk66HikOk/1tnigNh
5Fmhj8fBvPXa+BPG4+LG51TjVeuLb6ug+IJWJV+eHFALvOgiGcMlQb6NUwTgvsFT
mGZ5W3XLi1H11ldOtybz+ZI3omG9lWDllD9jhiknQ2ipenfzIk3M89KPRsRFDAZC
La+hV5dbcRMWJjdi1d/HZ2eQ3SlHfSjLeCdvH7+xuW8SLb2XHB4TUBpPX5Gt9qzw
jW0H/iXR1Oou5kMRd+59SUmx5Tvuy+n8xU6e+M0lOWaWEJF72jXShMKvhQ63q0YT
GU5PyyO2M9eax+2szVJQJiASjz3KHp8/UHO5MhdBQJdjOGH+H0hz5sF0sMSf7BPy
5k2Us9xbh9ftLiu8MyaGgzh1Fkp/QkH4ewfjfDqfMGjLlZ6NUQdYPtrPm+C31MsX
Jr1tXGXXwLeKpU5Eeni2seRhHIURy6AYdKOFsJ9TFN47GSDET7YMlo6mwBpABMXz
kFWwkVK+4joaDygRuEo8fIOCZMzf60IWkLJPn2kqIZuQEMfGrrymWdGT/ghRatUr
G/PRYvxUPkge9VMrwKo9SK6k+RhvYeXUAFydzLgPw5+4t5jfLPLbn2mZjfuHOqYg
I364IUR3PY/turfZdGRNfpOkhoKUTrMI2+xugLZIGZblR8mqMf6S1dAagATOYcTc
mIFhisZuoCM5a30YeNr3hB9VssDziHKcOvfYf6MfNmIFkcg1TT7zhrnNPT4Q9fSZ
VSKOO9bHSo8FmhaEXJP6D8JGrrT6H+JBO3l/BoJ3OmCQSYu8njZ0Fw8w65h3IoxX
MMYJXySCAwo/6QGnN+87B+YUCrGx7IStpRi85clSjiJZjA5Y2eRiL5JDL+gM1Vld
EVHwZCYTwjGD6d5saB41NEIHeeAiKZp2U0vwqaLRv6gbXixdMdbrJUz8rYzPEg2K
G4LQaQxgEO/knRUaD3mJ1cLPL3OXcgG0hRjDg2T3Pjk+8UkrM6QsyGHDGq3h1ToR
NXROBKBTqUgMSwsEvD3phADP3F94aC6P2YiEGw67utS1fTnbQnBJtPO1FsUvK8YG
F7m8jKENbbRPDK9zwRyURft/uDeEKyyaVb52Jk5Y30E5e6PhvOMGWF8v9N/KX4Gd
dnixCr138zKj4utDVtVcdaMK+ZMxlb8HKCi8iiOFkRqiubpQgDchRg6/B/4eDAf4
R2qVH2eMYHBTc6LjYrV6ayRvGN/MtfcoyInD79obtF0DxxvgmOD8P28rQ4UpSS3Q
bTjq7BC3dAJthfMvOYx5ulbup5JvIShC+4leXdfFeOLl7QhTO6WZlRCXL3rmYFOP
Gx5Np5HfLrYEMjfeyI6XhS1a4cHMVcWRUNLtYhOrq+nkGsDF/V0Pmnj7ryi4vp1C
KHQC/BvVHMDf4jzPJ+MzMc2ZeIpZAyBlphrBb17yoJ+V8EJ7ceh4gsvHBmZiece4
c8DHbmvP9cxcPNx5jW7jNhg2NlXsv+Yx108uX2Ns7wPEKM/uioPbyGFFfeVS/Ze4
04cW94du1t4V2dYp7KtzRBmB4cEJbHx65y1WsuTMutBsPNNNT1tbvBdB2DE9Jnn7
vmzuNzreL/ulhHZYVx/pBlOg5z6qkaAblZNS6RksvWVN9AfvZTaCJtKcF9NcTcTO
P+9CvbzTOEutf78xIuavpJFvMwtOJtDmzhE5lRMRUZW75LJ7ncXfNBeewVZO8TXc
kS/wNjEENcQZA4oxM+eCEfqO1BnQgaaRvQSKtD/wQ1o7nTn/KYiOfFuyULBQeieu
undAAcn6iws1WmKkXvuZqQJqo7VcuhcUCXiItPtORqRcDhze9JN77iDLA0Dc3QGa
Cp0GqUejmNIDD69PP2Sfm6AVhEdLLis1EY2tSqoXs98dglr9NNZUUNT6kUZ5UCWs
dvMtvhaEu43d44i/3KaJ117UHhnkiIbhNdZ7CntKvLudevTURw8pEKFXANHQo97m
SJUXthgfwNsVyBObSx1M5M+BTBhhnt9KAXp5pYl23GCWaRuIEQ2D3ov+FJIqTJmd
i38nNmUXcI1kGJK6JN24b1sDG1f7VWLM6IljhTXAD3TReTTfkPsy/ZqtLRwr4YYk
crcryR9vZQ4LOXjCIn1I9dDmeXcy7/a94L8mZAOVRBAV2uoH9A8ayfqRwBAoblFn
MUGlyg1pDWBkR5/PZClsfYlyKooP4O3+u52miLR4PM5JF4ZjyxCf/z1elj70R34r
tTfeKimxQdZQxs6aGKR+0+F7cjZKAPMiMVV1iNOog4IrAIv5oceyIO3vD48Qd27B
S7BRONG5Bz6mYCtyQm1Dk9GqmqPGVJpB4uk+BEY/10OPNASMIvuJwSJPoDMV1neQ
WVn5/DfcvAOXutg6RKJGXaRtHjgps35HpRbvAfi/P0RkOhgHsfTx9IA+chRq2bCT
tGGv2NUjSjZtYZqz6bzz1UUvcgTgJMIcIPXVzO4d/cqXMQz0N/KncVPV4bInEDkV
Pm+S+d+ZAPlGOTCMpuG7/PHvLhFDQwj/6DwXMz/7UTJxf8OUpQbfmeyE8FMxNKKA
JpofeKXY5QGjN4c/Ew7oOl1lEi2F7KdooGkUwM1/Wi1x4LtHSO8lxupaO26ubpET
sBgLW1FsuNSBbJ9Kd0gvPJa21xtdAUaE3dFoaLGwL8cHpa8QD7FOtXQ7lKqx8YGK
2hi9RKkmgVSY3z8s3X81TTHPf/gy9zaP6Q4J6UwRUA6vwDjTCmktFQ2psDYhFvVQ
owtBEMpIN7F/fHYp5g4MuhSQSkB6jvchkZV2GDOe9ieopAS7bTJYBLSTRyfotKXc
EHcNAR/RgZLjtZkvmJTph1rTf4j2JE3O6vtOPrrJna7tLCYsrBS01U5kZbPjv5cQ
BVxpUg2rVGoopgxz2XnxzWvWEJx27/yhG1kfPzZIVVHcK3mZW/6gqP8NjyWiMhau
0rcC//Y1Y0bnTJTG04UcfRxdtJly6uzrMFm59bceJcryOdnERgr0GpmJct2soIsS
ITGtW0f5TmtncWt+IRshdjoJyZRnKH5fM1Hleyw8HlzpBawqxqrCDKsOpjxd3IS6
Gj8aLKWtOX/kF6L4BlFRSJbeYIZbH9q+DgKBQVjvAtttKas5jwp8qOpMtql2SfmK
sQFbVB6eu0NDAeiES6YlX+5ngCE8zj1JLR806FzTuTckZ/NgP4/yZUjdkomP02j/
dTu08cIr1cMxHjx5nquUUzxvQz48mnAF4YVyNdpclgWCvmpSZheHfSu6dfU2u4mf
3zUTjCqoVKw07blpErFVfjjz88o68XHPQ8fGZHB8+Q6kL7AC43f6uVHPGU7+DHCd
l/d9i8JbmUc8AYL2Ryo5L6gDTTssCys90veG32YNjSwoBi7cmqoAnJfmFvcazSoP
lpdHHctSiA7iFf7lmSpDHSIGvfxH5d0IxBvDjJP5kIuvCqy/efnUi/mtWlgff8gd
kyBOb4DZ0O9nsa14JU9IGsVJZaIhwzas/9h572ITGJljve6rjkvzUYRApW4XNViu
riM267cbmMLZ3RecJn5qdubLsIWTBeDWqLq9PPTbJYce2eDgPSRymRqqLATGZHa9
cRIfYx2hoBS4K9/uJMZ1eW2/KwmOxbpi6a9oUOPJQZpqt9/GMNaZZqVY9T84yBek
cNAkAU8+UHHyPYNj1XQizBzzGhWs6fc3EOysBfd2L2sdN7CCwl/3BEBa4/XUbELQ
tvMsAu9Qly1306pcW7K8roPAlBVz7ndJiuW1fvu6iYoGCmk/14kbQPtlYJupdi4B
gEpJyIogGi8e8+uM0hiPQ6z792stPWNhlJTAPbETAe8komtYxZ/CMZMTr1gH4ek1
KtGUyQsYcK4WD3S+5L51xadr79qjJWh9jln+cCM4DYQXb4GXVNiiXKrrD+01ebZc
9B1le37G+XlkBRj5gSZBS2zOsDk1dtAsE9r+sgI4jAkWRx+aFl9yRzmNVq2Tcfc4
BLBwl1gPzUyv6Vq9hOXUG75tVF6iOVViQ0qdUeM/5aDoGxvkhEN3CUdMJTC2w39Z
TvJvDM7BFxdmtNX5OMyj6jP82Hl+4V3PzOIRVzZUKnJTGGnzOdITYI8wrJ49gZIv
O00eGmGZeRqg/QrT4Tv9HyFUV9IYD4ZQLY2N7o0BLYjEL9ynHv83sbU1QJ/3TZrt
SbmJUVbUuIJ3Z2qouUZm/9mXTPLdg/il6XBfuLcKj1vLRVgHtkXNT/wwItX7nOXA
Wji6crkZn5IXipVsvdejVMv6j2F7T8znjNPgHqwOINlHA1ZSP5xU+yz05wVr/1Pw
078b+dwuvu7zZEiSxa9AwZncMiDu1g8u0678egcQHdLNxL092ofV9mEO8Od0vN8h
o4uLng0oob8zgb30WDRp2/F+r9EpcJFfzGAho/pcLF1EqVD2DP9VrF3rCVlGcUQ2
/iZM1dQf0CYgDe8XQb3BeDm0+mAuV9szWdC1NSMMDjQjmGI1JB1ceKfIE4pbLUSx
ORIxq6aClo5zA/8QErzREHCxRvi/1Fz4zOkQsGXerkvEq/AxKGn74/82X9wb8lSx
lwM49OQQyTa3/q7L5fVXcJ1uNTkebLmh1LyGHLfUlDkh6GtYQ7bFh9oAZA4m8zrG
5IvY23dGP1hisS4eiK5SN0CWxSh1NYym1Wh/VuZOpacb4C827JxTFrlLFF9E7fqg
qSs2xLIGihcdct3fYF2K70BgyoDd+5uwjbMYK8IGUASkqwM3ipRibohB/N0mexjj
MhRlA1xRK6LSFjQimblOgM1ASci5TV1xoiGTPeMK7P+ow7EvrTaq8W+ySa//69mh
qn0juOV//h6MOSSjhqbRcYnvdmkV/ID8ljFJ8FVacREfWnIqsQFKum9jAF6iQbPz
BnWP9TjMelSSVMRTNW0M41Dw3DkD4cAibOttUSCbgD1+A3kqWTZ7QSKJhcnmOWyv
3NRPjIwJ4owabVUSfkcS6/w4HCZ2p2HN2bozxHqte6rxG8gHtdkME5Wc5URjj4oo
/BwStWY6mmW2KRcXj4nxRDY0Zw7ndLHUe7Eb3vxEqeJbkoREHqTPj1G2x3QeOc+t
4AhBUTmADfGqHGgP7J6z52qUPKvXNSdWSpVVp2G2Dv3cu7vNkmfq+bcOWBMZ8BUK
0qdjC63aCfflnDWkDDB7gINLoyl8E3tqmVrYrYpcVtNTmNzZdoGYd+8QEH0frHqO
NJj31f08u6/Pj46PBMbn6R2r3JNzHyG+DbitWFyCqOpYzb60pdZYpmsBGjI6k2Jd
lFAVOuTNjmkTLDo/uM4p6lz1QoQDOXq6460KTvtidAmwS+8Vd9BsN4/PMy5HCKQd
MXhDmCsJ7BJGJcKhTVYLsb5LEktWIuJNy4nNAPdQt5f5XwLd71xWoOj1rEE6OmCq
rzTLl7BbS2SzNH+XFa406PkxHVWSuLYg7Yyt5/m+d9lACeq6e+m7VYJsX+wnz+C0
iY4uV/t3OV2uVgbcuZyDLRVwhkiAmsLhf25VzojjRw/+AtsaoBYgY2JL75pHDAgF
zupNhvJrrZYrSUUkcEEpfOh0OVb6XZrhofU5lR0LThOOLQ+0zxcn0gfPvHFGbTu2
T3qnnM8JVe7VyVx9tFk/bHzejAr4YUyi//EVjCgMO6IVuvVMhw0AwIqP3ZnTSl55
YlwbKZql9NFZkpaW9cgSp2hJ3N1LjNoFiQGkD+qdJ7H79CSAAVC7plBAaXgVux2L
4+vR4eT+weIHvJtPWEUL0ArMi/YfY+qIsraMYud8q6+hmbk8pOY1rspJCdVplFZu
4pMgiZ0eU9Bm0XZzAbap/eLDyTcOnKKLhrtpKA9N+2wlWQa7x9B98YituIUzO4FC
pyB/d4LFkYKoJRA0Pb3nMIIJ/6rdkmuw8BWrdQpAHhMmUBcB2jikYuwP/jC7r+0L
djfqKRew02P62kbIH9/qn+AwrezLDyZpm5lwGBePlE7iYDC0yfxXqfG2lRjyE5E7
pIDQmubg1DM9FBPk6v84po7vzL6rdFnDeAnp5SW2LLZ05H7OiQD6R/ZSr9r+v+Cj
ctqITxT3Xhncy2gxROOdInJu21vGxKxFvG60pINufKq4qLSSYF67O80er1qTrCkJ
sMRtPO4WLSOPD6zpr19mwDlN1lvM5q9O8xF2e+59KAqrcxvDcLJ0IOXQdrpbpY/Z
gtYzjaif5RzDv2R9HTy6jybC6d/c3kgnos3feGhBBU321mV2dI6bZ25JMu0L0Zqr
xG7k+9fE1RsJJrVg30xPoS5pAC1GKGbBX/9EdnxhXKBXXVV2bm2jGGRnfI0TCw0y
I7ZPYYcZBqBpAitjw1LoooqyDyRMbF830nifWWxHhsv2TRxLdVPvnjhQL3nAaYaE
I6h4ycEWjiRmN9dGccyRRdN2mXOfA+hSUrqwnc7JJOaxxBvBJsQ8PphIP3tbNkFi
c0+cIOrhi65wcJX+/R9kFGTV6z8/lwKPpE4CjevmFgMxOzhxhG97PDAQh9v6aM12
zjuaabkS8iOa8jY6sQZWhbIRKKF+eYSkUXkO7mz2NRWD7ouWAe6jrbp6PjYE2f12
++YrKSvcV7bNPQ0RB89UPkDyiSnVbhrWcEFqnen9JMaLtda27T59IQYSkC4ouAIm
cArMuSlGv/GsNN0x+aTXgZVIa+L0MT95fj+HEesb40CHodFcULU3QXDFVsHuOdWR
ovNchf6RIx0xx4qaOsRpllJG+14Mn2IdDVSjur70MelOkBlacomuJ8BeTgY0WBzT
ndpGriKNhkC8jUZ0ts6YIAh/LKLCPwpv25WrOftDnSssbRV54VLxQHt0c+lUmMlz
55VVbFzQilG1z+Z+l107ruHWQqe+pUzZv1LZbgfw3Unz9ydN3hB6khT26V22iPCD
qwE29YE3WC1nIbD1HA+51FKh3zLpo1Nsr/3G25TQVA8pyZqZnJb3d7UP3HydsFqh
EqI/vDAWpKTQNKBGKN5DzC8uaPTBqvdEhyybZBA7z7oV1R+0QVtq+EdKScetCoyf
Gijbpa+la3tNwXdCO4IdiUdMe+e3eU6eh1wrXnl2U7qsTMMAy97dqSN+zJ5XgRqu
Li6CsOPyHjxfOlybA7fPJcY3eO8YoAkMVdI+BAHuhwFzWFzEAUBrnRL+xE/4EtoY
//X0blkbqYFT2zZ+F4pfBBLit2RLH3SXZjtz4ggf670jwNkSMkZHfDRBGJh9c9Y/
j2uvBVeHqExI6fIzP+m5W5uo1Cr7oMFGIsV3Xcu9LJYFZrwfdQWXHnjV2QAi6n8m
xDm7rLfnDr6laMqcLa166caVqw2oemO072FjHh6FjykSlkcphBuv1Md0+BGz43Uv
z5U+MFuHytW+8aI3Hzm7K/K4Fkn4yZRCIv43bTt7cs5WLjBjQZm8KcCPe4m6MAvV
ZtZmfoyoLd8w0RLH3F9kL1bMeykCm4x1d/1kgtpE7keaFGExvYZXXsLtu99Evkla
cC5YaLwQ88yI/7UQpiBZbClB9t1/SY5VHz6mo2tGp3Yb81Jp9rTDB8h2Ad+H/BtQ
xSUt+MhjkrnSpInU7oQUYaOWZ1wW3/Ml+uNq8VPcR8AfEELRhCpEVujRMvJd0Vef
SGAubTeeMNLzkXgMHUhKBk06p0QGPCuRjb6BWuywApbVKy15zNHivGMvnZU164zn
d0ySZoA2g5JW1lQ41A+/HY1P5JOk1ZVNjKTP++dAoNp0ls8GPfSElgkq4LZTUPKg
1cmoHziqKwVuq+R4NOmBoijvlANFvSTkrWowihy5s2Sxizbd1HREKCdfbPrrvXIT
LL9tsP34KKL6eJH3t3XsnfW0D6ii5UE4MTKQb/CGR3A/4fzRWur7LePRigDBeS28
rYEvK2KXfTwW5sSFPUIzLvljW6lA+09E2afmgqifOdoPtiJ1bne7DtfTVQXhyAsr
Q7y6QxlTnVu4ySsVimC7+dG6L7eQSPwbSem5Hjzu7uExtoYYIVOi46wOSAogiJkE
h0naaNLyE/JyLuzdwvBv08sqXhWS7w4O9ATWUzvZbDZsc9D70aIqXqFX19o+teTh
5293u+kINwvOVrKz11kIAAPGh6Ci2YaoBCwBL9mnS4nmz6DkrUnsciN/IVm/li5B
rF35N/rnVX7j3cokQDkqx16JQ9b2ZAtOKN15Bj7VWd8iUN9lpfRxrvqieymroisN
lYc/az7RYHIvRuGe841aTJz2Z3/EzgFzB4dedRDH4D/1HocwK8V0OcK7l6QJCI39
Xn3cDLHDqZpePI7bzUuuSiUbE/wRLjuz+dVXE+FEMIHEKDh7RbGIvUbJrp1sPw4P
BHpDQ5QVyo4nNll0fJDq8WgVoCPaugpFUx1X1hxSmd3SGUnoG7Hi+qjh/9fd9jy+
asoeV3znb1Uw76a2HMTp3DDCJ3ebgAleyyeHHVKU1cIuksK3y7I6Mvr8NKeSfVGU
StssQWiJi2c6jH8gDLRpf0MTfZFrP4i2r89XFDghIvqKjziyP5QI9XHvYuIPDCD7
O9S4BLxtSUEvkrMRaXfSQC+/Vb1C0oL6VdPyZ+3d1Q7gajzaSEmmMP6GRy+IlyXH
dBqyJRuonZz6H+JdqgY22gDrn1ErrDKfArp8tjBYShBSu3dZmZcbc7o0eL0I0y+p
vAuAwAtP/QVt0Ji6zUbo+Um0s6JFNYLIoyaVFI1HXT2zJPONF60RqFp9JBsWZcPP
gHScrh8gye9bvjRAEdRtArpjbSyyYkMA/rguPDVMyjp/ki/nzwvOnzvhNb4hPfCi
JwJME9/Px0HaUV/2j7HDQ9JD4bENHPgkl5ioyPJxkmFqpRTdCQqomHpRu5vsVI/Q
bljUcOx/U0J2ydySXvNojnGdxBUOUmq6dOGe7sQJVB1U420Haxvr0vB+bGQMKocK
Ponbl+pNT0ryC3uMbK0dcpOEIN6LL6dS4CFjIxrkd+m8Dw1Prm/AtIxLnLZ5l1Q4
xNaPDOVNgiaVvEC3sGvvHELlty5yxcRazd/PPL5ONsNgLg3knNoCYelFDityIeur
mtF6ug55lxoHens2+ic2534RL3SzvUtWGCuOdWrvi37TdS2sMlmnpFcFw1eL9ZsY
UpVrTFiu5yvQKnlo7kc0P+dwvJAOGwFRRHUsX40bOARqKrOB79msuVEa0Qc/G1K8
TLG/MlqjEv5I0Djr46YVRBF0GwbPAflzn+EwJvzecW0A0TrbyzYvMoivhRTyX/Or
ZjX0cJgzsGmXlFK7mygEZ/TrP/lWYcAdpc59T2bdfnRfLQ8ZbijfU4IN06gd+6b+
5nTWSf7CMRno/NOslOAdQI8FcTjwpR72uPVchP4CvXRv/JWvrMYKREeufL0TBZ5S
3yCmYSfmYSdviVOCU/Qca4eJv12unYSqMGTs7e6jEzXk34v5eDpgx35jKx30j/e5
NON1XJAyB4Rkipuzfwv3SpOD5v3iD42Qlz4bXT4+m1U9BwSjZ0JwJ+E0gLU8XtpJ
90UgsKId0N+qwhcPV300wlTtmPrDlsToZvVUxehDUVg+VEGmV8Jr8LqAEbDFPNoO
dhY5GQP9enge7BcqtZ3V/Z1l4/Jtdv3Lg0VvzGBA+5QULEkqsHoVze43dDuMxLQF
yqBrMJPMYjBL9d4iP6MROcqpU68cjpTluheMQ9JxwGTYurnor/Kfnmwmz5pAHdJc
Hsz1Xcbre2WjAVARHDPRtfm1ErsXv+9oXDkcaiZndmglPSGDG8+hdNkUGHmUDbCW
hbMXXgOl2PARZu0ykFU5nzM0Gtz/EvBGWvlgpOpm+8+nOU+9vZicqkfQp46iRXBD
UDGrLQtdDlD+dT1mThpq+akbX/LnmhmMgq+TAMDb1+/h8K0RZJN1TV0c1rPDsbHo
Vrs1PZhtTkmCvYiHBnzu6pfWVz2A3AgptjqZxBdoQkiKQFhA8ysTryT9HJBig3tF
3IVHWg2TGTyhtrggc8lTXmEVj0nfrLicVQ6IhWVIhFm1HLrvyIuCR9abtSrV8w8g
HYsHcQoQ/mfqwEU04qKLyYI9epTZ9+miGZ8nolTWmKIilV53W4O9aAVXm8mwhCHy
lSD+WZHsVs3k0SBrtMHQCUYsUkYfaL0uJ7UsL/qORM1xxRcokaz2QOjRDjq4TSI3
jDoqf+cQxHWtHPwIbne2gultzMG8Yffk5hFyOOnlzDrqtfCR9MtLFq09AGjAnxV/
Upk35zfDgX325uvvqqXinuUouWtAczOTffN6HeZCTrHcWaBa+hq8bmaMgge0WWbR
TP5mIZTE7mTJyORw1d9gcWVTd1hI2dOiolWLSioo5P6EixtKwRj19TMcMhuIeqzp
qWGMVp/eCJxuqotHnfb2VTRKiLsWZOQ2X4uZiCJyOnevNUJsV4eU7dlO9ZygXvdU
5q+MmGl0oR8Ef9MupaEqr5r7SbispuHK+LZ/syS8wXJQ9fSAddfafH9gCGltDLc1
ebGhASCVFem/SXevpnv/IHC4jm/VC69NCsekEzuKeZj7NDyanRCeONhiROy9YKiH
kkjYQkRqZdJffNMoRFI5mzN4W60uEaIccpvJkM+478FAoAOFHkuGYMhw+hASuxOy
Pb/GJgWmDU1uaRSt2mbPilOaLLPm9K/2N/u0/IWfsZJvHsTuv4DsN1v5YqZcchlA
UcT0ZYQEtvri1I4zK5DCOvtpGQQrgvGGI7HP00Ji1q40EYrT96uwQIbxLbkgdXnG
Ce6P9VSVpLGL2h+2KN11lGPPzlDPpabAz0Qq29Qzz3Zyn7E7UTBzm8AAApopxtZq
C1xveWVDk3gB//u1nnrluCGo5FExUT+2DyqxZ56hgSTbmjDAS60f7ygLDg5EWqqm
BFTEcIElCAnP+q4drbA1qdD0SnUa9YGDvJeW0sqaiT0EvV0YOWZCgVWB8AmeuIPt
5z6ab6oSp16JdUMRMlcHS2yLqsRQbPbKEThLWzU1DZD/C3yFqWCA7yiFoVzRiwoq
ULSvUaoW7fGi0w0y2L9EUAfiKkBV8ucO+JRd5pj8KqXNQNea24iNuNrPbD7VjLVz
zc3+ltbzChAZm+PQfVWs2iAiUY5h3Y7vyPEoDOBrtLlho1xk/nJqsd51WkoEiban
8EIdIeIpGt+dv554Cy7bvVI9E6A6/TVE1ShAH3AhEJrdN8kVwBEZNufPx0iswVmj
t4Tftmn19mXhWc9rpoVvOc0i2fcM2hk58FWq+orzsFlaqkEhlVEspM1gBFTeNjPH
At4LmH9/FfDqb6wZilG7h3mgMl+rldsmChR2qT4QuUMG2dwu+ox+gLcEV4K1bdTs
Fg19XQdEvk3A/I0ASSdrrY89ok92Is4c1JCsu2lwTvpfyw1H5QZ337ucq0IooNBM
B3jqZupflGd4uRmafsxUNsS7bJXuKYBvR4TOyYyn6t6ra09f/ua9YJnhWR1eOZxy
yrr3uowJY+73RnUYzH2IqNJ7pY2Ne3fmIvS9OCl/xR+ot9uf9u6XQZtrZhHpa7Tv
RJipXEIbUkWZ2/NtiVHzfpnkPaMW3mS3epoar7hN3yV+V/AM0x45DYhkWP3SvvXC
0zE3Q23NDq9X81FWIhyL7cvXmEbmL3pKkLi9il5qx5mSw45Oua9Rf/uXIJ/eWBny
tGIZnoEcU8dMRn+aNRJ1aDKvqfldIK5smvNZtlqhdwS2RLTAHah76abWfiqpwIt/
Wgj77OWx3GxHIgIyMjdJ0PgALcWVSwBRjZ5/V93XQDOyFoKFcHjkakm429E1+XxH
zYX5QRSS9tKu1IUt51XdsOWrBFubNmAkBkqGYvwtsS0mlUzVdAaHTq8Z8jDefhrX
8nVLFADNhoQUJt3Z3pS6HC958Vtl1jc2lujVR3b/mrR9IYRQjIc0PZrVUgxHlfTZ
IbtN1VOY3iTyxIpa1t+kYekIiLMln61F6iK7BxdGjooGuPwL/PnexYjze6J744i4
cS5LI+oN1yR9+DlEre3gkOe7Jiuo0jmFv8XLmNH4wVjp399Cx1k2wYtWabbECk31
IZG2EFiSQnbBFVpeXfAQ/pqYgwXbRvkSxfCULTGxUUJaG6OsoM2O0nqOKfxmanBn
Vz2HTIfg6GzxLAL9/bQWbC7oOUV8EUMI3NHFrsENcYj+ApfkFHskhZiTmoTX0Sry
ufffOZawq9l9HuUWDrE/syS4vkh7/IZd45IBKvjzXBh18lyHLOHvWYr0tJxj+0Pj
UV0teW6HpUBs8Dunr0ZXtZ/dis+pprXuso339RN+/N0gqCAC83M7FDBSv9XSFV2C
FrdSFPErNo1pq4iffWpJKYhV4Yvb4pEhiZsKfS2aGs7kzXe7w0GAWIB1z9qzfqZG
ryhF8lty2mckgX/MRa9WsyM6Ks8NC7vvOA6xn6egRO8jMbMaehEMdwZFfNSLJPG/
fHwtttoOdQELcO6bVnU14p12xZR4MjsQN/bD2F77PBxkypyZErU1soUGOhAsKNIi
8YASvMByk4oXmkZo+M2hpI8KFDF+2M1bu+jtLxmUmjfLi/8LfrJhKVzoADLD/nJ7
W25qH2v6/1Ymit02j/LreqTKfSFnRPLni22rYkF12m/o/xQuKO33m9vgy0ouUbBK
lObkbB2yz6t7WREKIPsOt9hZ/cLfdLbWwaqFGDNNSeUdvbi2jHFCV6zJyyuiJzwv
FdEsiJFRwSSIJf9EGZWEGvnd9pmEF8oA3iFGf9fku7ZMzH9/aupkyo9H/7gmC7KZ
hHuDMrv1llg5cuCncVWy1ApLjKhm001NtyIqyx7xcSRjkkvOgH8fCLRuc9pgpgR8
1gfR1Id3c6pAkLShnhHvYWaZ8zVTXytPu7VShxL8uJCADcz8EB/saMb8IPpSK7qy
E7hzK4RIUaJlkMvCkCUpvYsoou1oJeVFaVZt7VVDwS7T3maBAkJJ5EPOv0KCQgWI
ReTQBvyc1KT0tUZfk9vaTNDV073mSsg8nzjnDyYTPZWJqWP0Oyb2mTKvn4vCwm4p
/ZAOPihK0UmnA1tiko8T8TXoddw7V7vCHi3MuE3H+UyS1TRPwjge/O3PCS0eF2jR
htV/FF8MgbXwgIXe4e+IE+zwY3+es2RIsWakEj6yE85o+N+vXronjsddMrhNUlLq
WiCkx1hUZYtd3P9WyvmRQ4VT/R01o9XKVr+76VxDgX+Sn5dnPgrwkuLZK7xKG+b+
vgD5APo6HCn3mS3pNWI6E+LWq0zvxXYvElyf+rl4J/Gzjn45mOT0KpZD5XlRfCTs
JP0Kgreb+NnY8ZAZscUt/6PlWChmQ9QX337i+MeyjIWCCaSrqVgJ7tecP9NiJvZ5
JqPtBWIgGPfbgWG31C/Y3btkPnvnOK+LvUny/L8LdDWCRLBgN8prTYJLyDtQ8YDZ
sbtLTrxjWNtGRaLBO9AsJXUg4NAskPCYnMd3g4Oiczf85MlpDWWrU/TBHEM0uMM7
vlK0p3aoOosz4SkN8aYM1C6B0PHZfnqEwUOiVqxwktusiTiCTUTApQmd3jcMI+8e
GFl9xmgQiHBlPY/9cgJcDRkDHtf9dHFoaAm+/8d42zKMa8EIG2DvoUymP2Fo/cm/
bcpeXopOfpdrRexE62ueumZu5GefEiw+rTNUovm0v7ho0de4OheDYKCZwEcYj3OK
l6ehoSHJBHfmAoo1FNcfN7zeCYlqGbUlgqC0YDqBDeSwC/ZLwj0EKOYxkpeud7b5
QO50FSXPSz7DFaU1GLspFY22rl/p/D5Y40q4IUi2pp8aUeAWE77x1WwFxDulyUUB
UrSm33VKwBQdxPuHaKUKv6hYj4cZB33ahJJn3UWWzzf5hoAJri7CvRzvac/IqgMh
LpOqLv8GTSRZCecZWcQhLSXStHfK7dqHtRxTENj3MzUoAmqZdiUJVlSmdbeLLEqP
oZ4DRFIThlciNDaMYdtcyHUXozH2SQrdhER7n7okjMIM6FZiQrnfM71jN00srMDw
drOavBGO8Mf103ouLXW3cisD2i3nnP1ocYjz0N1ZwVXfpSVZFkl5KaUPtOphH4US
9faVZzN267pDX+LK9Vmz6EaR6xUhPKJZb1N+UQ0FjMgctCEU6c2t3bGOLGhqGgEq
5D2clFoz/37+SsrluBdsOOWUSb+73E8vCc0pWVg0ceAbQIU+bzV5+HNu9/bsyWhU
4h/h3frqYQIa/uAbVJrVc+VzuEsxQ/9dqfbSWAhz+ZudUelaVGjMLuZrNVbFLQqT
tJi5PAw3eNFMoHHFfpY85tbu58643T085u2Z5xJf7mnE6HO4w1BDnxTphcAfx2wL
YeOCePW9SJ6X8mJ0ZZ6XA/EoxUtfLV98kKIRRlkOuzNMoZLdPZv7S2vF9f8mda36
HZNjpu9uM4vPrRdcTrQuKc6tvoY/AUwT8BQ7h+W5HgGRFAkbrHhQo/F1/YsTk+Z0
PHv0Y6Ux1B3WQca3fDtaUL9OIs7C8Q+ztZ92BVxcJAKZa8dryUR11udSyTd4LY6M
fzNU6zRSGnHUHdRB5NslN1Hf7ImK/VV+IOUbIw/Zw1R5O+ohjVbz19dS1Tgs3/if
Hi4TdjBGDa6y+wCeuwmoKaJmHtcRNqcL2g/3QO74kzMyY1jQsSfp0anGcdz0B/Kp
mwGrLyOsCwo1GTBWOX9QktJAuPeXpCRXa+g+MN6Rs8vQ3a+jJTg9j2j/nWN4yz3i
e5n+faasGw/+EqhoJ9Ljiitfm3pEcJqVTuwaQRnxSzByCC/YuVU5XT+W2NZUpO++
iTdxra7uRuXXOiviCOdkTBzldOKtlwXQmxRAMyfcL9UuDJ8EuHShxf3qesJ4mZnj
igbptXpaoaYQllSvH4elkscPm3TLYO+cGGjGUPT3bMLAcUzbs5xqC917yx8zLDSQ
akwXdgY9kt8Y5h7f/NBknSn3gkXN/Cmu7/sJVqHiCra5tME3Elb5vNI7hDEna4oj
MZcJyAeGRcLeNj9i8HdbzuiT92snb06s+s8ZlUZ4CscaNen9uHcjI6RsVmqNFSd4
t4CcWZ2MMwTFBGUXhLL5O+SMpIFiSBr0LZW05y7/8ENQFPP4FuvLiWtTodjJ1zQm
VnitzWKlSDwpI2XoLFL2H1STL0OgZycPfzPFyh3boeYYduytgTyLzJkAdkw6wHh5
O1ukcd+oLVK+vL1oONVqOT2sMqnsL43MExzj+6kEg1Hrd26wnNpKPjGO/rZDLezp
kRUGbb4LAwzRuWODN+q+XlWuJEDA43SzIsGuKZZwAazKchaYO/hir4lvNqhyhF3f
Rz6V82VI/i1rHr4M5s0ZrRoZ1recv0ir6+OxcKu4HeRzcuU48DlcMLWpWaxwL30t
G8V3gyIEa1EAyXccmUFKVqAkPFa9SzGhbgxx+GTz5z/ggeMhN8HRm9N/YBOxI79D
rQnOW8Jh+aSpJaMzPKpagho1ey+DPY7MtdvXE6Y1Ga+bq34LeYpSyX+ZzImk3Rds
xb6knHaK+GCFNPYINhqAjVqDsUPt02HYJBoAcaiHOrlKJ60Yaa9rX0tUc7PvKpOY
X5gBLbKIClIzjR1mmhTdf0GlSXf8WONtx+hkPol0n8RDXavgXx+TQi7qnb0gFge5
B26t/5+zjyFrZPRpkLA33NKnGD2tdfyigFIgobq9eZXi9EBfTa02wcuw12A5eElX
TIho4tdvqz0aqyijRLmaS8W9Flvw4f0D5ry5sIBa2Z68gqIGg1cEPnS72rKEnzzI
V38S4rSn7YtWk4xSULtBW2R2fEQZ+vlNJN7VNaXK4NT8HTPw3Rj5Y1YTgUNYxAvz
zV01BVzP+1AgtqVO37FpxFU03owLZbEWVqiKHqR0jft/5hMvoTwwXFSJmR4HwqSs
0ED8BGEa83Kf6K8Tze5IMHrgyOtHhymjtenwk0bvPnFJwuzgz6vbm9NZwBxoxhvm
6cK0+hx39HFeZQ46E1H4BuXxdvRPzHihhqiwN5SeW69kqDnMfm97gVDoI1wRiXcy
Ta8rsEYhqdtDM0Qv2E2Q+YrXK6309WckxwE5hd9dB7wya2ccGcKMyyicnyskp9X0
nbo4RbUHxoLWXjaWoOHFlPiA4owgTNk0kJPAIG6YsO5fW4Hwqv6QX7M9BuXMKFW/
pT3YVW3zAlwxnB+C5E7jU8CwWUx5uH8+a35xpVPKXaYPmmTsTzESl/+mpfbwSXCi
JN6Rn1i+6ltjPJTrkrjrmEGah5hrdBjDcObOrP9MnAXedeWNI/wI1wRTtRy5EAq2
BIWdvSM3G+KocezJ3yhoBuLqA4dcKOK4kCel90K+hZpdL0OiJSFmciYX17ItCF2a
WEdQ89sTpOKBtgkLD2eXp9hVYHZCkKDSm2b7a5gneK5k9EOq4YP+QHFU/zmaDyLS
Txf7zAjk3//ycGCtrrTcMiSiqLIW9IZT6DjwF4Bz65MhbWlzMq6x/EroIdZk4czw
RWLaQAoHZx+BIHhOvSNa/3tx7yplVcHztpDyoBchJtWH1La2J0xKG3QCuJouWFrJ
hvW2zga4e83GVTd9PSzvTpNAuygTkMdVCvUkh9IHDJy2O1rRR6MAhtSirgo5Vk2s
PVYYSKwqpMRGr5Rq+Bn4MYJxmRdN43M/Ps4h+ZIcFF2aEWslCZGt2J4281799FQA
V3KRaNbG3U0M1XKmEGTRdMizlNSCHYfjzu3+BGUJduADlXlnt/TPalKmTdnlfIVY
M146FbLQz8DmHlok/3gGvVI+7l2vrzkNArfuwi/QL+GGqa9au1YGuhTvKWONJvqA
lN60MdKcJDXDsAQbsoLMPXiWK8lkMRXAeqXYkvSUO5vmvyWza8QrQjExMVQVRPjE
U6ZuwaTA8B6lipjd39MUL5/r6oOhg3yUIgTvNReVdI4T8Ro3KgDVmq12cNnuRtJ2
U7O/uXyJWGgGGJk/A5vcdswDSUhf6Ute5NEE3w24gGkEXpgcJiETR8lhBdCMEEqU
pp3UQRvLcG7o/XKwZzzySperedIh/tze3ndyhwkYvgmqhqi5DBmTF1ntdcBeAl+b
FW3+WB3Fnis9tBovCNLW53EbDCSQbq0ITGmmK1BM7RdWN7+XCcs7qgIjpkXpC8fK
DcBscmkoP1S8gU0C4bzFiwkLVQFpVXgUAHsZAts/XUQm9GXdRaBGUK4Z3U+UEs1U
et37yhZO+wMWcoYeAgRSXXMn7QdPdBHnqDhPb05+9b51OgW+DcKgi55LS+pCcBdD
1l1CMYdmAmr9GBnqhmmhkAjNNNUtK2OdcYYIuGgj6Va58atQAU82Api4LgOq9I2/
Xi3og2pBT8fQdMPAzH1mLaXFp9eNj6g6XB+H6KEmhuPhPFgABKdsB1RWO/5LBdRm
nkJUMnhc0ofMo+122BMz907HrJq1HzLXF3jOh5BvRM8iOf710Vp1OKve2phBVFtb
h0DdTbIJB8t7ajZ2AuuhLdfWxrWUfMoE+ctw1+WPKrsxS68cYKmVGE+JUTiILt0Z
VPgyVkOu4pWjP6i+Dbk1KO6jfco091hjUrXQW31fcN8MQgLLOsPJnzx9Xg+tiLCw
xUAa4jDyJbqm4QFJzDdtgULXRHBJ68ynYX0ckBJ1sH/ZZQbNfoHVQXi4QsXvkWr0
/jCEWwUrCpfJbEMaa9C161ULiCVDAW8rjvTzimNFecvFBfgAS9fQR37hw8zF65qB
3VfMwtAov/lXUPJ8z3uiMNbrB7QT/rqnaB2IlWJvHG6fPKGjkO24nh1fLelxzo1L
0ioWTkoaHErHur7p3lAuVWAG0BioThIBDscBoZNfcqMJwOwVzgq5OodpzKIsFcXU
WhjLLCWd8zr6qGQCvy5Ze/N2AnoY5lTwgXpvlATL+xSgmIUKR6oDc4hHf8bgi2hJ
zCjwJRgPOHQ8z9baMML31hjociRK9hje87eqwgtdZFcoBbB8Sx2dzlL9Fkc3rb+0
w5ch5ELqn8VmEbrjVQEv+bFEdonEKC24F3th+pVhcDHDjnxVMjg+rBAz79zU8rlv
5HQ6CNiL2CbJUyEEStnILsShcoTB8fBVEAS4Endc93CtqDwkRQtx6ILRygFlP6+Y
5kxmnj1m4BMmqV/10tTxoTVTIvInzLUEIkJQStGZddwuwzTqlZmHEWmTXdcYGOCG
8E0DCNCaKxH6ydsX2WvPMmSPZWgo3eQEAwFLYwX98xvXlIhG7xn0BCmI1UQG6at7
w3R165IYo+gVOQSpu4Zc5RKeIB8KHrs1pMo2QSYDohmmN66846wSfdetHRhyYffY
B0Ow3C8qHcOXbXTQJHr0FBp7tlPqujZCPaNZvxFEpFqvflz/w4FT+VvWqYyho3WY
ivjdTJ603I9blwx/d4UZbsvZHWsVBtuguJnQ96M2Y4rF8gjsuIFmphYce4QMwW6g
lB9vb2l1YKRKN8d0IuVNNpckOjm9Fd8t8NTKzeD0dAMVp+baSvxENT4uXmxKPYLN
qMaNfrlSieQEoGhAVfpGjBe/96W5LT6KxI+EZCUYeFwZNVYM6gGFHu+LR2STt1j5
NxYUpGarVjQnh1ihimBK6kLYxNIhDPcPNxgbMbOTtfrUcwmaVz+MUaaxu1tOX/Dj
QmcYw28NRnUbYB0B5POYNIlC93ZzARhObynUd+TgkTWWaKUe6m0a+HLtFOKUaM0L
srfoSlw+sJrOfGyqYU3IOa9OSs9VMTiGLugGxn3N0kVOBrsiWJ1mVslg84I3wce0
ZvzcfdIXWYyhB7L7gXR4gqExPI5iRu8di+paWNIx6Lv4S/q8JJuAlAtbw6/+LLcz
/gazVewIynYHO7tXvQPktHQ5uTPy49LFI4VrV4T3aQsWIUqFUBZ/aMolpXI+YNYJ
9EDXF5743VEtJpBmOB0i2frwHLoYV0BW0IJw2UpdfUOazvsGxl+UO20wlT8DufYr
/CvEDqKQcdyJjFzqrvKvq5shi8PreWILzsyUgsjkI8lxhy83in1gWgy4kZDYzV3l
t46s89ObZKpb9Td4vcUW67SFE0wS6oh0VcI44wdcaFlC/Ze5dOL7NfIILzSVFjck
rXiyMvNDdxQMUP+ZS4FPW6hoqnWbpfl4p5SEOLqp3bm7mfDJ3s+KJpqfPMiKIxaL
dBxCjEa4Ii5ku/Zq86diVHedm38Z3B+FPf/q5RL16g1sY5Aa1X+0J+EJQWRI/RxZ
iLwxWaurPjkR3ujF7TOhQLy9KhGYu0Is3jt4nZF45JAYqGJ53l+jaVLaa9ktlDda
kLaRFSrr3mFgfJpPkDluoiliXBrjgonOyJrYIJaf4eqlIfr/Pcr3gyn7qEOGliNP
SKlyE89k+IgIwdgKUfAcEAihI6687zvbsJWn9gMWec4ZfyEqMXr1P1MIFM5G2OD9
50VkLWF7Rh0TmHqPF+QYrWtA/EJd4jhh8Vot2OKuZerT8NrygzNDOdpTRdlYC6Z9
/C8HMplxNfFbIkx+3xXq75bbB+dOYxXAR/NYT9f2wXrgmMPvlVww6stdzl28MFsG
WowrTe4DGWhhoPg8oMlWoJ4wYYqqeln0JGtvXnHldykopYto4CyuNaMntYMo5qpY
OsU/tHmS9k6SY8+DZqyJDPeH9zxN6dxi6+OG4RS3gRiGatCFcw7/b6f8Fc1BD2Kl
SnxAXyZr7mcBsf9/I+xxtniMRdMbBEv1/OMH6/vTtQxNU3UiRpEk6/HvqUbqbpzj
SeSIsh9wFct0RZdIWZbLJEBIdr1HOc05dlkeidGgZWg+OWwS/98BUsoNRZ0+6fUN
5/hHStpti/XJo/zqTL/jOI8RT27350EMP3aWVqq/gFcTm/GX32hAE0L3mZ+OWWYe
G5IvNeL2wBW15GTa4+XTV9obvzE1CodqPV0YVkgYXIQv1SMSVVdDrioupG61qCIx
M4xCHUSCUDFvC/TUx76nuD5fwA4EXV1LnMKAQwjx+dI7C8LHB6qYIDtAwijtjI0Q
oBh8URv/C4ZxmYIM13P2Qgw5TJzsRny1aaNmDbPLpa3XB03VU/kqS0Nxm/S4aLZD
ukqdF+5TsqJAiyup1V43upkdMb01JVES87BXo9E9zp5GwpXyOSZmyZbBde2JY2Qc
NNRK15X/nx+1SJCUCQnoHXGl/b/fkXThmNOkH4WLdSVH2w1snNAiG6aXTyV2bV6Y
FmcTUdbJNk7Q6GU3+lrrXlt81X7XmS8q+qAO35EmEOXA4ulQFrBt+QISGPEaOz/F
BmjbX1vsLoCis5SpWanc7FKm0dnR/RmfIKv3XLFYyBnSvqqjHmfhklM9ZQrdLp5V
MraJycHEWXYeAnJCOhhr8y/qoVCN+SyjAdrYtz/S5m0eNARsuelbTc4jbQOAJZ4X
YDwmXXA6RJOoeG+D7E0D7LxPfHnKNzejO948euOjJ4f6BVfS/w7uq8aBx3V/K0Zq
14B+QdFi1m2E9qOqGTy9aKAiKtzDgUBZHblbcpO5bM/zIlyIeyTvQVLz3+7E+JyA
YO3YJXLshVmfy4ZbE34pfymPdHh+SCpL/iwWT52MhV1u8C7XQvUi+VDkYXPZ4XAH
MaH2z607d0v6Ljf039CbFRr3TnZA1OK/EtmCDNtqDZ6FHmCnwXkb+avQyjj5t9qp
hnNMHTFJSkswW8YjBjBR7XKZiH5F2o2Nk9lA0xUKfqr53EDgA4AGwJRrCJjiQeqa
6DNqVzmNWF7v7uWOrQ4epahjr6DtG09ERFnl0cPq7+PBizYpSoig08UYWoUYJP5y
PLJH5LiagEYAOGzkR3MngJ5gylaREzoUg6ipJlOH/4+xQ92ZXM4jQWp/z/MMmSSo
iDLhbd5lZEzPZgLjrrRvlP/TcymQk0RNWfA7aarO9K3EAYjrvqSeNJlpNBfMvKJ9
CjIw+wtOzjmeoiPp6PW0/FeT8Cn4DyzHRb4RbA6NSPXQTf8G19NrSs1h1ixVtRUP
rXMXLK9XRc0d2Z0y/1Zi7TahDukcG/d0HyPgX9iY3X8tJc9sujaodFlJxKdSOvgb
OSSE9CdUCXHiVM6OQHzS9W9jVrxzU2L1OT04p2uLPnH8wLk4sT+WwEEuv7GTKST9
ivmYQVPL5XiPnfUbloobzCmaJQT1rBifdn5ApxOMVHpSLezDtMfkD6yv9sD5ClmH
6s5QQ26b07DJ+DUGMXwi17Qon5AOy4VW2YrXYYIJL2KPIz0R4oNJVl8CT2+yDFGJ
h6U7WNUe28TYlGXD4DMnFZV9UUBn6YU2HrK3h4Ula8RtjJqpfm004U9qZN1nGD48
nrtDfVpC/BjLI3fY0ocS6kVcyomzaHj4158OwUGKAB+oRtc7HxQo04irCSizXqMf
d9LQrDtRp8mUPlTYp4/hsDEJ092XRDAqAvN8PbsQcrbfzyL0eSqLdUQtBDIHQIMK
nGbKfNqDdFIl38uA9oc7smraO6XAihO7S9PSO9QEy9Nbwy8tmyqnM+Zd8ftyln36
aiNCf6NOSclS/A4YSimp68AdKD5PU2YFDVds981FXSI6N43iPKGcX6O2jmtAlmaq
MceY+EqmdufSQZQLLC+w5QXqcN8K+ONrzWzLWu9/F8UsVBYBDx/A0jQmHXxsLjzC
QOo/Dwx99foggja5xHdUVUqIMCnpdJuPhUn6fy1GED71sj+gTbv4RgWTntIEX8SC
DR4XwSU57Xi103O4nRTw1MfuYZWFZ68Guu9zpf8NLIIGBKJFhIu9KfvWUsBwm8Vy
sRMePSyofW9i39xA5jAmHfirBuLIdHKp83LzssN3NsI1iCec4TNpkoDsfL0b3opk
eFlC3OolRWJlamtK0tshQEiKFO30NW6c5rEOjv67sVuun3un5b9j0oPvSOCDzYn2
opL7Uq7TZmDYDsQ44bMqwbzIGO0UuGdWfJTgnnTmBAvR4rVZJSzNimLSF2/PPFhs
ocjIw33X7cQOy5Ve/yCF953/HvSnPm9cXSOZ436yBorBfx71EQF429kUz3p67HgX
NlX186x/SaiQeXOU4nMCpA7NInSmZn0yAITOl7pU0E1n/2tNFLCURqbO2WKIAy25
Dz/Ysk5vcPL9ph67USKLEBwK6oFWpY8TyyitMOJMO3nRNTc4T6HQwO59YtVlUyY0
WNpK6k7VomGVisNMNsY/silvnYSR8AwJm6U/bov/TfqLa+PKgIxXlOAMcd01l2Mk
GYFtQqTawZ5IdcZNkWcEc9C6mZt25V1ALr8fIxmnrsJBJ3tbWRDu931qoty977Cu
hcBgY9ve0UUN90kJ2tpKGO/h5QNWGyh+l56xTOIMTbko43O6FJjGUwRITgDrHjPl
ebMtFSg5KDWwYezV8A6q3K1Zh+asi0NbPbjwa2YOnZDWFYCggjZSmQnEG5DVaPFo
5sPqAnAVoRlkS4A2tL60UaVvKJCx9pGs4F2hHAPAZ8+n2swQMdyieKrTKJ2O9Qlm
jOce5u5zk+0sGx2T8yOimF4A5B4ciTqWcoa4HKXZJY/AHi8BsBz8giH602H+gfi+
pvNDO0HbOdXOD1oIE6Gahthzr71XJN4m+Bj04JQvyxKPFQTae47wipxeImD2N8tg
FbP2sb1xtiGoVP8SOCLYg4e/c2BHy91IPFuFscEi3brxmGMjE98U2K7xbaHrnWqr
klNbgNPIfNGUCyVu2O5lBPL4GINetfjGeMnPKCghxNwYg+KCDvoU6vZpX92hL2x3
dyDdMrQsxTFq0/H9rS6CNejpJoR3iry+x7EtJ8Z4GsMRxOjAbLP0kv1hnwYtWi+6
sn+q62vPdb7q/OoiDPza+a7hL0m8FuDc2O5XMJGVFF6iT43vPow4qBKOUnyBTH1U
KlAyHkEK4eTCAnD7mZ950G0EPVTkrpyo9ylypyPerROooVhrgnPQOc5v2g7sbtqk
5u9LidWotcziVfk3VxFJDez4IX5A57Hx0LWQwh6BF1U3MYWKEh7JC0buXdEO7t/i
vX6r/r6U1UcjOOdh8OJsfA7871ol10I8vni115usIdjkE0xIcsoXGsGpaAEdhQv6
FmV1V8MjrOgwzPekLVDTvxPtaB4SE6KEz+8Vpqrq8d/6b0qFP2F919u2ddpf00Cl
S1/hGvRmGnQw2ymjh2rGT51E/tEkyWUFJoWasH4KUoGr1SAEvZcCUYGbLccjqE4U
FQ85jsufyDKBakiDnoVFEMJjvj230YQs9fhy0JBzEkkdRdDWXD1CY+3Lz9XTNkmq
Ws/d7XXWeUmCd+X8oNQVsabIN4+WNG4LL0qdDphLL0nFxmSXByLM7PglX/CiZBbo
ztYAg8CGzpvu9e8Kn4mpwQN7CWUXYQFbYKf5mx3KPferuezblhZF8AC5kKWFZZ0B
RHrDuzpkpNYuylUwEB+yISCVH/adCm6YlOcGR3jQIzLKJaELSgx70lMQ2mcHuKh0
0rhm4sGL+pwW+/qf1QgBKygh9xYQsG97DCG4gkWy9jhUOicsrJOtL51OrQu8nTZ6
bdlJ1X2v43T2uD7iO1cOfacJ0s4Rw7Z2ThsVsr8o9wQ+2wGlEsHxeixSa3+rXbq4
IJPh4fAjhri/OMbyU3ykWUvvxgYfz437DDUyyUhFsROCvT6WJRozwoStkwsRhj0r
Zf1Xbfsj3o62OeSXkdNCVwg1+x/k3F/62G5NpaMVo+7I/RjUCkBrHQyzLbOpYurb
M/ISr7I+CKbr6cXBA3I4Tj1uMPU7gUIYuX328zLxRhFeCWjieKHLaPUnmWRPCTaL
JpbKC2zJveB6r/DjxlsgNSuu0gtxkLUfA1gU6d6pn39FimYZwBUw0pkJVgesiToj
GwvRcYZlabsvqXlL2bjXx867Iqs6RtJrjQW+uEXspdfk/jwwNy51Ti1hqst0zsnm
fekpKPpAMrkBeF9HJR8Q8/Js6iJxP1im3Yb8t7rFIDUbl4pFIh+TkH2CokgdtyMf
CKXeuISbugbPAajyB7MZFMaXqZsVUWfmc9rafSWkjr49aqvegq8Jd4UIWJZYNWxq
iC1wcc0OIKKyjKzGKC1uw2FAQxB3tMY7I4Zh+bXg7bzybeu2ufhbKDkI+HCIfZ0k
FllA+CJD3OSSzphLhpQ4kMRiyh1iRq/DTQNff/o31/ecgtHcwmSd+wTKahM54rnH
TU+ToKMzjvdbSdmeEbSK62DeQn/0XHrlAYhLGvpyFcENeeeI7c7Sbq+MxqIDKzzR
g+coLmiplrsloIJlyNVkLpJBYuqPkut2x62LKQchnW4TXijcsLRo+zJuowOktGL+
VInb6Dd8W1BgjrbTdwsVUIIuiYlfcoOHdE77YrJc24ZwRN/9QaXH+LkcB2fnkEfV
KWscHPeliNkZiBaxuA4WpplmpQ26R1yCYln0damjNCcpj27IC74iJ/XDXYN0gz/K
fBtGvqWjDfECabJPZRrWVKV6r67DIWEt7I3Iq9NW3+6EF/PBMxSI7aDjs07/BZrJ
pvfKrUxa+fV2j0WD53ZU6bOytBZTO8KpBlRlYZrKWbc0xIwDXIjjKBHHw7yH95jT
nEeVxprerT2cTS6/GbFJDhF9lhslyWY+IB3wKO608eA9n4zWNw5McrfitkHseR39
85Mtebl8WF9i5msEMkeFTbpBNV1e+OyeqbnOl8ANzbCfJACwZzpaT1NBHCC8tP7O
Wuog5RgdG3S3EWqYtpw1MdG75oqBhxiH1CTx5ieREWltSWvmlblp9wMC4k5VOaXC
BazegoD/g6AqK7GbZeVjKbQaWbrhuZPh39Q5dYNOwWHE27OfIwdBouHu1MPpr9G4
R5bxl7LdXvPbtB0rXUxLjyVqmbf52OTuyftPa9XnwQ2BS00opmfm5C3aC5N0Xw0C
LEjNYZA9sCrA3NcW4EcwpP8732XCv4uE+Yb2dhIm3UDiQDSUDy73VLZHOkiQ1DMV
36d6ZRsyDxAy2s/Z+ew05q7R8FUQWmptg3/6lc3qZEyeUC+Mn+WjdxHQdGSxSo5m
Soir12D9W9xJ5+O2ht+IV69Vhd64yxp4ReE8FT/bSVN8lDJkhNtIl439DxCIQDAj
thLuDmvVDH/9pehWLV5iESIWrakqgJ9m1S/eguDaFKQJwvpK4GzrDB72j/jr0Jzo
egxGo/xlz6Y+oJ1MNaMzOG+xnVzrcP528usrCJpbxXrk9US07wKIFOTI/QLx9yfc
GsdHFlW0IaCdpC4oHTd/wLrSFU4D/V/K/4djLy6Ncz1kjVTRveI2REx2f+13Ulp4
LTzrXhj/8Lg5RwIccUvjy11rMIk1CTC2s65n8u1Ryy/cq/F9EOrlc1IwAL24hR7P
I2aYx78UxTwQkGYAln2H4Z2PmcxNB8fjBc+yLO7odnFW6NISrkFjfA9K/aDSe12d
paafdMc0hGy2oyG/vwEIbgiPXyKAr5quSCfbGugGfE0X0d1nbxqY1i7EEjl95Vyt
nyIX3l/GAU6rgG9ztAlN4N2JQWp/yNO9lk/EYOQ4NYIUktBk5cQKFM43o4pWW7PB
RNRk4QfybCPxL/gHDCYgMM8nD9siLahrMCS9B30Fe0s/iIdVE2/Mkub8gmmKsqwy
C2PW0Id71HPVzlTR78w/Mb1XXhPFENhtvZ9M9lfIjxjs93W/b/eIU9YAZUgYm52A
x9Z7hgghz5+Vjwedw5USLqVycwMpyaf0QPeHQHQ9M3ZtLzha5le5zVAPdOwhykmS
owdxsdTMc8hTlGWsySgJA4NedaVgTygXNQMCHdDdHjSkk9Htp3GI9cLB7cu0bSMr
iBC5nDqivMpatikR0ziWGh3Zj3AlXHyxmR0KjujUm+oxmctMfY51BROkxNB+I+nN
hJODI3feC40GsBRL2poppWs5OGZBvlkHuxahV3XEV6ZoPmltHncbi32VgGBTAKDP
ZMKqXQkTcqDx7KhucDTzamDWJNn2V7NkVIWT9T6kvTl1fiEfcQeHrqJOKlwWnFiy
Ogyuj3xjfKE+XgInJtS1lxtK2YBvpAwjPPeLBY+411HeraTrHdEU34D4XbUCvo6g
eFcPe84XJfyT89hdKgIgSLCgsQJR/yGAsyve56bugtgXaDDnivV9vKUP5+hL83cv
mJQhK9dHvOTTXiDsOzd7wy1DdeKWrgGZHwP83tfshkMy4PMDEIcU6oSw4oQPF5AL
UCGarUkd6uRxasLoN/7evcOYYPk97NkZrrgP993FdGKpMg0znSdMU3mTmRUu1Q2P
NbuucxVNp6Mm8rcJ3bXbhGsoJ4vzVC8CqmL+ChjmoQkX4eYQDuLgMJXv6Sz0Hleb
IuXbcN8cfE97K/kyWe7XYvCQmPkKVlWa52HETfIkIGAqX26yqZjEoi3tueKaXYXl
DL//NfHomzAT2zBoljab28ZO4em89K78rlQWFU+5fIBf2RqDhIAVL6lsHtipbbSo
xaNTZp9ci92BmNd9naptmGSQg9lwKs9Xx8fJGCA6ZqtAkLPh7jgSVfigzSjWeSgE
sVadfhNbGpoulP/rgjGc37xLa8Byuv1vmA1277BNCSmejdNxw5zn9/tRtE/pzHke
x+kMAVuSj4u6Xl3Gw/Ehg6PMRWqw9RpmDtOR8ODpPpCk2y4DYDjAqg2PYVmuExb/
a2j6s8AwbOEKJQXXnq1aqjP++TDycWgNX3LvqQKYbdrliveu9q1qvA9dtVIbY+cM
iVPMmMI+pUESurQKVtl+ow9N/la0xdPl8XCPjXSqQsiWK2p60A0EySKCJjrWo2Yg
7pv6qtFJhkF/yPuA83p+iviSiXLRTiFn3C5awCI/8gr1OFLZLRzw3Z3zky5e8z1f
ltDlKYtcj88lrx1C9RKO40VJaRU1aODQtfVXSxV+FezwIlEJXAu51iCfb6L9qaJo
0tpDxQKdDiJwOvtPv5QV+8cCaddv0uI9mkfwJTLRAlGagsHAtRHp7pT8svxdCLrs
Bf/e2QX6iruhGeXc2K0UXY/saViGkvZs05zTsZjQGtYFTULivjJw4bc5qPV2Uvrz
siM2iexlXk+Rnq5wAymvCIx9Qzj9uiKtH0nTqFl3v9apRZGP3dkQX9zhizwyhAZG
qrsA1RQ66pGkrKAV6v40jrXeUUSvEb1xxuLlOehXhHk0SefO1V9jjSJCpD59LbPx
e6BraHHXVsAT//tBgQKVHIULhF5asoGhETuNzWd7Y+YuhIEgP4B2WxpxAWuguYVZ
C+6HAkfqXBKf8l32GWPkJlaSpFR/Fqq52GlpBixV19WswMk6b+fbcCvU343ta9J+
NnsL0v5VOClTzjEBTWh4T+8cYuftceem/HTSJZcOeiFcUp5CbFQiFcpEEGollgNz
yXW1SjU0svE52H7rj7VzbyknPm5t0ubFHYKhCcQpA3Hn9AtDMUVyD4He/w9B3qfs
nyn+QBVxcmbe7fK+bpANTuMTlg8MKBgbTueOc9WvI8JMI60LejMn4VEv7TyBKT1I
j+x95qnPLnjqOhUkCjUWrp4OVbWEEccGndrmytCSTmiwcC62ub3bvyXSy6ieihv9
pUG06/GC+6CDeT8IxqaWBLVzN7bcQmKsmP+tUqhtPNutx9xoEvMmW0mE2ltlKPhk
A5IIN6jRMRpODjdHqNdPgvcguJgMDv/tyZZfk07K+AMppPr6qjJ8Z6w3L2aCfeRd
bWs5ZhRls5Nos/DEqYSbeqksjmjSuz1HQt+bkXN9AVzQ6mlSoqDKHAQVcW7MjvDb
TVjGZFV9GeFsghpp+t5yo44rxG2JuteVFtTMF6OogPVWKIo/vnyUSSeARX1Avy9T
+7qWDtMVOsCsTQR9wiihd1wk1WJsgXlPhFEx41GsSbG52FohRALnWYpV6/iIvdW9
EsSPskSSjrSd6p1uToH8hjQedlWnUcg5qtdwr+Yteg9JxG3BGDgT5mvYOWJVgBtu
oLwvcjuQP6F+Pwu65c8DJHxCP2oPQceLR+iTXGUg2cDkD82JOL/tfjawF4rUEqyg
jG/m0nD3fGnvNeofcg22/kv+uJUK4pXBQNw3WKPybTnJkrtGQ7xhVHAldBoIyNXw
nkgIIK7+4jl/mkc7UtY+j4rFIFhHXOemduc/JHQ8utiahGhPvjnCXJSH+bxrEGe7
FDnQgyquZ6p93GD5uOlDXEBloa26zsm+qa4l+ZlHtHOCXQIP7ac6XDYsqIOOvY9E
DkJ3P9GTirzh1wRfUKzI4hjOZWK/09/wbTS7GFFse6Qt9nyLIAJh1VeBiA3Q5tAd
FPxNlwhPnod0qkxy4ULgyvBWzGBjyjbDtSK1KSh8KFUodx21jB5CBFWo4nArqDq9
QnmDA2RX0tZnzlL0wpWn7feWeBbVRYxLkmexfbeKYUnm0QNrzIgR4IcTfBkpQ/4u
U7lT7lvjYAkbxwPn2pOOg7GbPkcD41ncLuXQf+MFtG+sbRN7uvOQyo46kY5jEaVE
W/O9BV1HBwiuo38LOQko3g2rJodrUUurb4f0TGj1xmij3WEEzNyVCbAaCdixPTRd
wd+qOJvAJhVYXe0UqDEz+UygMutOZIVIV1/H0tICVdsBw7mplscZMRGkejtOEgW6
JoMjCoB2mvxBu7SYDmFUdZYeyyGl8tBISJ+nYfirMhOC7MgUp/S6kcWeqbC7ziJY
CAZ5weDlMJdZ/4kmTkh4VcGEp0+GVQdV0p9C9Y5XtUap5l+BEeBs8B+eCKELGZGT
ekpxH9zgO5diMpHgn3/F1WQc8pSf4HbHRhiJdD6gmJyk9gqQo36PNPu8EDSoCvVo
hE9YjDuttPuFO8d7IUmaZ9O6tkrDy62WInVzU/ZyH+FvDhIhJ3lgnx0mLs+SDwAA
WWFvc0+nuimAUkU8FRttl3xmNXd9+pMk8Mwm5EUel4znuNGfev7D1aVyu9o1vuSS
/75iO6CROvUzM4qabten1G9x/wi2CNk3Y4IbPC6YAWBLore9fMGVpcM+k4R6XJ/p
njfkv9b9fq+o9vNeS3dXRpwWUt7vwg+MCUBmKf/bZCxXa+Ymb7aP1u0ujOPtBo3h
gNU/MqKfemZKBHhCqJ2tlsZlxSow/el1gmEAesFmQZtfm3/80mCLyYTbr8WesvW3
zKWcbVlWZmE4+xWAHqGg/5b1823mVBZJts6AoXgezkFee/fZAo6arRGJnNyYrmu+
RaSnS9U1QPyzAYFsNpwfHKL4hsMSDo7jUQnn3c/J90l4HdRiAFtua7lgZPQr7UHv
trPCDIhK/8qW/TPNBR/C+D3F7JFUlpId+37j9NLAFih/WUP7GfB0tiNL/n1t3CIc
PnPY/j3n8n/1Nge8fStetIBNcKUURmBS2gi/xuNG8CN3N0vrhDfTLhuISnHzkBzA
HjWGLv6/dvmO1+7JFtb3ydXv64trdacmYCdKvo3L9PlR4yNs38rg9OfYsAmihCkI
+iD45s0lL3pe7ef5SHINVnY8RwUgsLopYV7YSboIrmuWUHds/WeUpNwpuqYEu7hm
j57W3NZoqrkb+bPDnZKF3BUG04qV+oPfdoQ0e2fNu7JEpA3+RQm1FMwJcQ+IQ0u/
P15pSi6H+lF+rBlchLVsQ9R2DklDvVlSxyr4PB87dl5dP03OJnzFa8+bO/xBsuPx
7zGWZBA1S7tQDUx/DLDyr8ABt8fPBO7JmE13J1EBPWrc3HFO5O2IPeviGol5YLtF
Ex0bZ3FC4cMSj6rPHwrWRKsoyk7ODv0Jy54y1L4sCsYI5VqVddr14V7iVs8iA7I4
LNmUtCvmo5r4ium8L2g6YURZrCnRx8zZcO75aPtSQ9h9WdY/88G9C9WPi9p7xxDb
Q89QCgeb3PZ0HrDIsVFVeZ3LkGGk5FFB63kkjnBRKIyJnromr6Ik3nfPPFm5eXQz
lNdNxcdQmicobCuJ8jQV0LWl+Sx6vbgYTwiBQPMWqYvSrOvbAdm0UiJuzz5kfB4T
zoLZj5DayamoTGDwY9j/DYIDMSi7qZMUgxW/DLbVdjIzKGaYaqAXyM+X8DZU4jeT
vLaWuLC+g5j2aWem1Z3dzVVTYilDwt+d5jAHpRlnEjVQg8LymJG3yAYhRs9B/QEs
TvBK7c6Mv2uQc/PWV8JWuRY+jGGNus642KMdIkq28IQkByfUvkbCwbtGa7r6zP5Q
50SIwsbZYCxZJIzchXc0ODFfLOvNu8NCujho5LogD1WDbvJmL70gGU0VaQVKK76Q
IPYnINsscBcdRWRJo+uUbXj8wWDmslHnfAQDdExA/WTvLLyKPmOpNUWqRS/5kLFY
DHzh2OxIPvOs1XgVniaJBoGPJRmXdhhRNWLN1VLrHKgMCky5iF8S5F1ZEgjMkD9R
ImnEy+XLEgVTyoDAsbTetw3ambb8D89l6y2DYxWomPw9AymEUfWWUyKWANWD3wSQ
GU9AckYLgBPHNnkyTIq0eXsdbeAee3o3ZaIuhMJv/mR1o3WUZedWF+3cch6DR5l/
X0oSlLOIVZ/2bz2Dnjfc/IIgeKYoF5xDORHtRdJAEOictK6bCw0hG3TpJqHyK+Ug
BxKQwh3Dc5dUaJfxeT6LBrvvgLikzgy1WlRpL4WNlQeKvt9VlRPkbZacJjuT1/KF
vc34X/xl8IySoMvcV6RD6nfWtegdan3dOwy7Z5Kx3euUttC28xMD+6EqUoOral7D
WqOdbuYoCD8L/NWk8H0eV5n0Q4nRiu9pESKI9Jm4DRHIOUIJp00l2dxUCEctbPj6
0JaDaqoUEbvLTa/Vbd82GtBJmGs/zrjr3HgLYTkfIY6ecpwfI3EPbxuy9XnJl4A1
VKIQmYlHrRF1YuhRdINvmy6xbjJRh0l/fXNir0fQSSXzMJKqw28W5O6aTqNvZKCn
AhBxOUfklQzM24o9bsKzSaQFpVmW7Xb8rWNHmSNnl3g6kxNsgrhgQS9c1410Cay/
zWgB81yWHW+9+4KJ7zn7n3izIQ0g6YlCGqRJGXeiqLJnJ9jNlFX763YFgzZnh2J7
C4wTctKOn7FrUxkuYJ7wjSscG4YkfoP7yCxDTRMUot5i1FpKrr+WjGAJ7U6jkDkG
+MSIqsUaTjQ0v1IimuLNhNPB5m4/haQUgrvoJlR+mcxDgUrJ39aOj9fbM9UcFJGY
8vnbd75qXRnG3MJ1W52l1PosHMxqqmT0ezMT0XfQF/1trlt9vQ0vLNXllOxvSKAa
LTldizDhzqEBRWUqDDNvJi6qeS6e20bnc8RzwEwOp8KGBx5PyvRQcPcAviXOSuJP
4pvMZOLF4Ij2QOor4AUmn+gLGLUgHBuxCNHQEZNdFV5ovmZFshaXu2iJjFti6b9/
15XLv6l76PQCbG7hl9eybgpJw4OsjrJb9CqX1i40OTt3sh1S7kT3rWGa+VcK7bjU
B1DkEgg5mJX5p04QAHJp0jiK+r4m46Q3kMSHKQo3PFeVoGJCAyPw+sB20OR4D0JD
t9OpMwKpMbn4b9qFPAgnMKK70aIGTVMznBwiQvCaWUtmHROsgJB4qr7dwTzer3go
uDpp4T7TdBYOfnkH4tzqMgE2U6bi7Agtt6v1Q3qTnMSz17Pr/1OCQ9+fWZmUGEC/
a8rR5g2tee1eXLIxZaU0Z5NZUG6W45aPb1aAQ58X7bosY5TEGRkLujY6HUAzfP9Z
TarNJXQd8XRjJ9C8mlZwPQr94vkPw41leuK63DANCAB0PFm/WbNGRlz4k0YnXuxl
bFZ6qQVf3/FsviKNIfiYH36ly2OfGN8iLstamsyqpaVHFqMP0qUFSEJZXx7CEulm
5cODwJvGLtIrwVuJJqW33Itp04Rw+foJj61KgqtSbdpXVAuNRjpStp2CzQ0ei76H
t8VA8NTJUfFCZbNdzC7ve441ZTAemzrLOO2yykfDch0cght4bpXmGALZWISXjy6X
m5IvVK8zMfjQv3t1o8UpkXDnJmMQ4RYcPkaZRclpSQj9/dnuLGMCg4UPxRFIoJfW
IbKAHBdWhwI3lgN5EZvWNwOuIiEoTf0tyosHuegF+nuDAjAMT7x/wv5oO5sw9iLD
gGrSkMr9TaY8aqcYEecLqW9CaY15oRYtzJw5yXvoBRRFc9QV7hXivuXR6yAZM9wq
P5H6fgVWQsnA6ILXcJ1rZEambb+hojzCRVep5rlvcz0j0OqMCjUboddKslzzmapG
VFzA5YvXRMHoB5lJcmnC2ofGTy5HgRlflNUeEzx/9c47nX1o2yRIylESSiBFAelP
+npDjJWteOvnzwGPGCbtFxJ3Yl8Z0achpzORWx4pNAUYcWB8k7AIc34AVQ3BTUwU
74sH9G+ACZRbodxBVgwvrbeeF4dkXO3CFDFV98ndg0MzApgpvV+NDXcVNXbU5d60
Ra+zgqhzM+NOWu30/f+0cMiyq0kcbDx83fzSCYLf/AVqLspsJdc5MSTBiVu094tO
tZOv9a3n4VOB1O5y2ufu3uYdTQG03Xs7c/GtSTi1tjePfxVCcKcDEoUjpi9NdH5J
2VnaGsi7Ac7wdhOp1yYpYqvBiNKwhUSddpR+YmmnwPcdfBvp7x2tBB8u/Xg61CYH
eY1o8j5HJuLOhr1MwYblQA3ZGdUCkzN7aN0BO1PrBr5ppABnJzl1bOF8TRVBPhs/
0x+qYzK0McvXFB4bUN6/Uud+jDq7W2heLDymQa5UZdOTbfk7yYGiMNbkgEL/Glex
MKrYQzOnXm42B4+675sYCN9wa9rqF59sm0T037c981s36ImiCJ0F7JoipnxFLgmJ
6T9LifcWQmwBQhGXOFZdKMMhJvF4Q3lnpDMspAbCKkqnQxVKS8wTldRRLDBep8yC
xFOwp/J6A2bS4HU5zY41OUM9bRkMZZYrCIfbxx7tw6quXJ3wy7LKUcA6N3qnuKCr
B3dpRxmzMglrpDC48n7cGQvKLmnxvQLC4q/wK6z550G3FzuV7yLobx8IrCLUbmL3
bdm6nFzlWegja4Jz6ZKppWsCWz7bVX2u43AuzR7yV8u/tSbT0NMtJMLNUocLT0+L
jm5twmuQy+G8g0ORrEIrGdBflgR2qBJePDyquRRgGjfGS2uqT0/CWOsABhRTGb5A
l6gct/GfFWzoySrUK4gl4KOhB0eL9RM6GZHw8NVXVV5QHrqeng8PmM4jWJBF4eaj
CItM2UkwVeznlaxPmT75DrLCrorT31dvJ9GZsijwqKT5CH9Bh4/V7V9YL/rOaPvk
cnPRqxCRu5mqrmA/iVFdRAdtMaNqOpZDuPzVuttdWS7jEeA9NJaOKSw2YTpgrLNl
AA5O5yzHjnCl/gCR1/IMNpjrsI4Zc8s2bVzqfKMrAafTT8xeXQcRtmYJY3Qp66+a
M5O7QQYrMV8l02mMUfFfzJ29Vy0GjQbZH6D4s7wnMN6ESygQePU3UiihD1oKVLsz
E9t2ERlBZm1l/O6zldA+uvOkGw6vfuhImTbutj8+Xme228MH+FkZvO5mwhuDZzM6
EbibmoHtwXqHVYYfH1iU+MuQDy5YfHQESUyiQKcUqg2OLKOw602cCZ+17CKZOIa2
J3ImxWcdoUMcuZv28gEsLoZENd7K91MoNNjK4+4moPcvgCS3z1bVR0COuKHNm9Bq
L0L4ZMJz8TpPa/6PRaZ4076zig3Hg7PeazHxu3nLUzY/JlSGsynyYFFqZ5vP/TlH
rWxl4AaChsFmumR3go2qXRX2WorWEfKLy3/KYlMF30V1nXgPSuqZF84GryEqH2sy
pjuR6NG3hjx5DwE5n8hY51ZxH+ZnEL3nE/86rRezImuh7LP4jxA0LnVR3u8stqcC
zK5nNCWAbU2gJADDgRzj4zmgq1unbSRBRRS8jYEeiCpaBgONux/t0q4tOne6bWfj
pstes/LMmER2eZdKWqwTVMEV7t1YqX0oIoKrxUac/WMaylzjD2hBz3EX5M9Z/eHZ
WtKIvgJoPtKkJJQ5dJqxJZUCjk+nbNJNtqrYJepfqIhaobKwYVlJ/7V+XfVkqVvI
pgUN19ZjtHaMdw6SXd5OlsuByWt6aVVEUTaVDpLPJYURFtPTD81RuVD/kS/YZNo+
v4uilzLdHjDCmQdNUZRdlcq7ljqQWjfe8OFntmUndogxsZGmzJEQs3jHI6FqwJ8f
eHmrL4LVPBZQja5g4V1WUsqaME5uOSNPtrHlczRXgJXhw4yuknysvpS3oQidn+v1
P9tGdJ32wwShtBZgAKiW771RoFdyoDT7V/mktidWdrsNfZmZivgD836sFcCmIv6+
TzCfg0xz57IysOdzzm8JxGzjJubgqOdJ4x0A7yppde3ukcua4hkf0yp0uszrZcsF
hxReQrL99XTuNYrT//sEuQD5BnvVTg0G+iNjdmRXnG6EFSs0gBTbZF3QM+AoV6Ve
Og9g/oYrnG0N51y6dHUap4wOfr1bv3Y9oTXjXczCysMll16SW4ZKqEk7YijmgtDL
Jqkz6qms2WZp8ojCUMFtYzB7c6WZKgB5BlBbLqMdg0F6Z5VX+FF20W6NY3U4w1dh
TnLSWyLVqYdgAoU8RHANCbH2ZqZk38+7osNC6cl1OXGsUaZIjUc3RlIHrAOUiEwX
oimMU7LvLKsajO1WXW691JoqZNS3r9jlh6kiGifDlUJhKecZXJ8PGgv2rhChbP4I
KHGBfRmX5LTSzT8xZE2z07PRuvnZ1wUvVcu9Alg/ldSZwbpBZ8hx0DvtqoUphKWs
iz8h2Ieg+4goqxxs54iMLHBT21yLaLDdZPrfQQbSS5b4QRm040dJ6Uhlfgo3JE2h
MgPkeWbt3wYDeMuo0/1bW5+LR+LF21RFm29dHZ95EHhg1C7+3j/vYk7VNSvvH3cA
45TfbF3c8ErQGaDCsQVl11HC0P2ksjHCv3m2Fbwr0dALl/ZhGreUtUVfgx/j1Amu
2i2z8oq+ZvoaAgVJyyOjh0bpmXtCJOhrg6QP2rd1iiUq7OexwghpQZUQvL8LLNCo
RvBb1j7vJ0rLbNT0lTokOFA+vqMRKHF60TwU9KJYkv5Eu1+WrDKVRl42pnNE+wc6
Qmo0VP5wSBKQ/mTPL+92rbqQHOXS+WwmLm970XzGI37FhdhjNpUtNVveeDNxvG63
AaqA80b0rIn7xLOXQjEaTZMFDhqDLvNyiBkVQD24cwEk+Nyu7lauDzZYiWbgPDjT
bCCpTAtupljvdgn0ypxJruiNvjr4Izv9et0U5CU6+/L4rEqjYS1qa4SRCABEXA/i
5NGdo+vzE5y2YMNipynSiDYiBqlRiD6bAZgmujO9ZYIe9P+MBOmXwPXPVejKAd0D
YSsxwzt6lPPJLYFmkGzkf8ksM4afaTV8ChXCeu44c2SXLtS+WoDFVjuQQrMYHLW6
rS9JRNUwPqHk42R9IL7I06gHgHupq9Ks0+cvwkVUNAlQFBaZnlzTYYW/4iG3tQPG
Ajxx7DVenbbKTRROvEKUDuSK3e04Kvp2/CoicT7Go9N1YIhE2WMYE1B62hQdm2QL
OacaJN5nox8X9KjWM/Dmv57D5CKjpSSbAOEJPQ5DLePtrMPXPCwm/7auaknV0Z0Z
dfTl7LSFK7kVJEJuJ5lB7fBz4A7fgCxDVWqJ9VKj4KcAPbs9WtNQOe7xDvW9RfNh
IvgfN0UADTEO0HpByI8zPkdp++LBXnV9dFvbePiD4ZtmAibpWowZGES35T7/KCJ5
U/w0gWlsWKhQ7v4dAMAfFj/dsnWO9ozuEP6nqwGA8rTCiDoS3QSN++gBwaZdLFgd
/wzv4eJq2Lw4EruQr8Crhg6g5s9klyc/BklAiLKdlHu/QI+Jn6cwXINcqGZQ7z4W
chhWcJjgx/KLLMgKqnvNlJTpiyQdZV/Cg5jEUohv3so07nU3aVIlfytbxetNGqmY
tbvgFFCbLx9YCUUPtjmZ2cBaMYhlL7WmpE3DPflKm+3w8lwHtjQi5+726MQsRZQ1
v23uZK5MKc0FMWHCjfJbLinaKiMMQphyo04IUJxzXblsmwO60GQjtVhpvGDDLaJx
RGUwQHgye+1HdTkl+1EHbQfjIatwc/VnpV1yM6NT8btiim0q4dTEcwlPXcAN23Qc
0vM3GRGD88CEDt9jx13C7bwUACHuEURlBJwZqVtsNyDPbnU+GOBjeVyuux7JbRDj
Q0MBVXTCZLHtYbi/c1JsDVEbR8/ObEMDwueuWL9H/TWESAX55iOQ2cl+EHRYt+XD
bvWnNwJini8GedAOV7wHyK6Rw7PVGNxQwLPR/zPrTZUFiM6eTTwdGAWSYkB7xvb5
ys1lnVIbTxvaTYI2NNy06NNF8z0M1KrQN0WX6nHY6qsiumTREqRbd2gCFEQLTm4d
JsdlspGT5V2jg0LRZ50aBmLa1rM4fX7QCQUfpLwejsclTJpbPklvXbRjAVv3eX1+
09XR+naVGaabIwiC0hf8AeL7wxmXQig32I072jB/fvnAsVIXegVsqFFneeRSHfTJ
O4FmDXiZ6xmDtwusjl3zqTfDXBHUrmOqfvK2KVmiU21X67vGS90eYsec70fYGx9v
WI+1pQalZMnQP2GCfNvkllMzTalyFrZwYYO8ho0WgKTbihtHJQ6BlI419toujiEA
ioHqv6AZLaBZD1wem679LcPHE9S/T7ICnGbUlMGcDQjrod68Bja66AR5Mbazo5Gc
W2/vx7wsdIAnEsUw2y2uMIv65Vucx0ouuY3ms8HooCwdmAV1NknUyEOH1ldG2/cg
Id+JbYxBFBG6JFYxt8a4WPOBKKWWPKhxHaW7N08rQ5BQ0IQMHR9Ja1ZRixJQnjGK
yWAXfUItkQ5mz298C8YwAiZJnSOijDtn1siaIUttQ5nLOJ7zj3EL7CiQX07S8lA+
nOSB/Vh2pn8AAVbIBwhwHfbBMBhuGDMeXdexO+4LnZfItbueHPxKX/eHzH01KzWv
4aYO45HEMaOm16ifUGpvpkmM5AvL0M5ucNNO7NFG7dZ+5QuikDX37ssRA4aV84Db
2C+ExpmLgRZbUo/3An3RgXp72z0etCcVG+jNrfAIQLuzBT3QIqKNMbrcuKhyYyG+
GOivXZry18IwkuXGbOz0kxKrljR3R3xnV08WhdKThirjeb695AYpuQvAZcZ3insA
QBeIS1Rv+t79G0ZuU+0J8nIcp+MeimB1AloOGRnrxQXiTm8u5tz6LpsoXjMuoPXO
uapz5nMfocZRSua3cByCnmvfldQ6fwnoGjRQFeQcQfmNviDoxL2R4fI+EfldHrc2
tvgudeQ2nzK9Oy9S/dyRyQMFvFtz4uDXHT/cStRZ5vDKl8KulBLUdOxdlTlJ0nQS
FjEuKEHlRi5U/aNFqERHaEfDv9y57TZGtwj1i8jdTvJ9yMAmPJ5FBTHnU1Bg6srI
oo258UoKV90G++IwIVULK+Wo0Zk71IZeMBa/x/tufhJj8xx9U0e435a8osdav6q4
eFqn1BEw7cj8Qnw1+6yscNUcPz01S0AMxJuLsvWhzfdp7udz3Lc9hhtA56/bvr+I
RgnaELzyTKGWjrrtBAIZRZVuSrkz2fs4t5fTq4xXyWmPltlkC2hvXebJyi7lvI/b
fxPSZfzoH8tOji35zpagpjChv107l//OuYDQriLgX409GwgNPMU9I1lge3/l8+y7
fKxtXvThwIUMXIojmlbwOSWCWdcAzhYe3/H6LokoDFYqw/E0zbglGhUZSZlXj6DG
tTJYEzEwgbWpD0HnGFPzMiYXsiMinY4MJXDskofcUxOFtPUftB6iDL9S3rFiDWPQ
nGP2iv2nUd9/rrJNIIFtN0lTsGwdnZEaML1+KILCBUZ8IVI0Uk2Mq57d0YjL8DsR
Ao1kJQa0OyAg+4o4PY6lw11IaA+hJ3djZLQzwPTLz+CyZoVE3GcN6GEcnCJ/yrPq
MC0dkXLdbg+PdHS3s/RvRbOJGajZtFE1LF28qnh7+GQEPl4XWUo6tfbPxSKlrxYv
sPi5CfKg67hgiz7Oqc1UFluoMvDo9zpKVqT82WwJ6mMqSIvE3ki4ZBD5DKnsb1Et
EtTwuoVmHdDeI1rhQuZox3T90lsVx2vUe7SGh2KME0wnWiB5OcqM/GcidvF621Vp
CH+CAlh4PheOYXyB6unha7iZJi6TQOe9Z7Fw0tpHI4kER+52+kK/8md8D15ILO4i
gg+Nk9rKUA60JuhbW78ZhESmOT1RPK5ADF2Oyhv9/48H8mAsWUSREIFXz+kAb+qT
XC1VgX+G00hVuCJl7hHTYqEKu483bdi9Mrs7b4w2StqPOOE1wWbbNc0PvuMZ1USs
2odlz2HXKm7Bcrc1CHNhbaBpdkqlqdcwQ5p61eP1hyMRyKFNLNh59jNR7VxyNYus
iFGkqCJKDl1yewxMt2TCpTziTV8jsAoJbwUn57WinyflS5IbgbRl+EAoKtcdNEjd
IOdB/PK85wsf+bhifp6BWgq96aEYDUkahRdYdBG2JBfapZit82IgBteqJvIhTJWG
5+juAJrxQjmbhQxPN8juPTf1hI5W/Fgx9T66ZTr/QxzQTLIY8GaQP5qCzncD977E
+uagMkul9JiPUquooqFoS9S9UY8N6emuQ2vTzSMEirwMso7gDaNgzUiEkbRQ597Y
X2xhKnT7+y7NW5rdlBInk7SijkD5T/Ja7hbgCRbrWi5V3SVlJUMhNZpfEfd0V8sw
nD97CQ96UHma3pdCwdZzu1gq1MfiATJBda6H6COzCkMYaYsoiYApJDHsrIutl0nV
vtDuqOKemhqj3ik5EqAjlfNos7U/7VdtD/guca5Km/Wh1pSzRidErJaFRxvMamJx
NVq3orHTtgB7q8NnOgJ5a+C//gviHGSBxQnU4JoU8jS9NhoZpgs7L81MexMwswUr
tZ2oT4vFpR/PoHDw+CK7xjJOKQn3qcbgb3Yi2c9M0F61aK5ObiN5QBqrl1kedtNs
hlEO2lijKnrx5q08PvX67KcDJ9RWx1J1g5dr6x154Pw3ebozaIy3UjpZjR6z+2sa
HnmY0+zqk6AdFTrgOwAN9aBVxxxWgHk9MV6vxl6BvgsAjWMxQcHWEbPI9OtL7Qhz
crTJQaEuiNGg2P+xv7SLzxf60JZU4jXLOySIVzNnzC7DGhyMgYPVe2zyZPk891wa
MVJ6FuB3mJHRDP+Zy8bIcx7IjwLcsg8aYxWc8hoN2b1eAVoyK3OAmFMAg32CNE3P
xWAEVPXz+6TcoGDoQKcMZFpAH+Ex7x3KIqKIHYdEsku4GSzDOnP9c5VMQWgOpTDD
Xwe64RmoWSwQOYdUB9Vu/0ugK2XEM94+Ji8GC4xog/VhgOWWvv6SYEvrmovf9g0J
vtsp0sHtH8acrN57073FQvnjHkijNogHjP/MZomNDFmx23qNfidC0jXaCcyzzvSJ
x2QeumYOqcd3F3yZFi67IzuaUdhvXNHb9hzWd5o0kJ20+HP6w+0IK4LDMAy2S9mT
niCl8qSvTQ6w3vj309IqVZqVVkt+bikgwCPsB/FKSr5zNMqvtaA+F6wJ0MCrpY7m
VT4Z2jkoQ/PGo0XL7GbMNESEpizfuT+7KRq97NC4HzVKfhtocHmMcXaas2Ri2lrN
uIEfHqvTQvmfrylBPSpit7l1xOLluwCpHHKF/MR5sI8GFoiYd6TLJ6kNaLzJJCpK
USBrDPWxAuJ7+HV1Uv9wVf5dqMQqu7R03xt7uL5pijaZ5bejSDR6HowJoO2Tiiff
X+Lc5eNOW4LkKijLL0wEgfywjBZpYk9+cM77m1EZclv6s6Ed/E8IRy61hUKfRDUk
WMv9oonlBCUPowcpWI3KLFqPOUH/Byk8INCdoEqgXXUXTDoWeqooMVADNKF7cItc
R2Cui+09MSfATfTT4tdVkJlI7/8DJ1rAO4CsTzp81n9bHcxkvSMQ0fBfF6V4G4L+
O53LNV3/+70aYYXWiV2A8PBiBNvQqMQpesxwE9/RAJso8d6REanh1BJkxMFdHmGA
CqN3b+iS7yI+wvPk6XJIzr0TA/MX4XsyiMZnKEW0YkLUkFIcty1NOlVhWqGIs0pZ
dPiBlYxrGoGE+BSYdUggwOkWHW9pvj3gTDMbT0NGbKYIHxC7YuCZhwkAtFALTFey
oHDlkGlbwXkP3e5gsd2/Y5r+ZQOOe8fmx4uK26E+LAczg4DSKPbMPWJDI50SF1bo
NPjgMfWBCv+sXfFBGDqXX0wIM52wJRHoA5ZOmIzG2eC5ZKm4F3POUerGPdt+yWck
YsYSbGWsrC1RyjeGIcBQsmSiGxb2eS74TRefGrv9qQZrcL7xm16/8c9IzCRt91Fd
O2PUfqWEpEk36QmEYytsLxe41LS2vkDtyflJ+rRC3jY/v3OUMoa7dlZ7e8+z/cG+
U7oK75xtbzn1F4uEeavzA0wuOwtgJOA7BWKS6e9Yf/1oaOzLXl786VU4BGmWfHg3
vd6L/OP8SWngw1lLdWMoFB5+rFgScO2aSItew00h5fOjCioi7zIGFHZmfNMO1zYk
9agCV+R8R5ZTODN4kXYVbxLRsXH0pmpmw3iUSjEEHKzqwS7siSQyIvS2+Gnglkg6
U9Fuf1MfsUceeer3AJjTY/hAjtHFAKkFRt01sQevUtAR5rwXjU68KOc2uPK3nHSH
ZpNoH0orvVcZM0v4q3f2PlOud0zUb5yIpl4jtcxi9YcXNjAdG2EjutZf+jbGaE+p
d1z83ESAdzxuUMDguTGorncMCFSABOKFhZnhFn649RPRfgdTF2XEztTi8SGgR7/4
GEDABd7xDRX5nTIi9h0gbn6vd7QnYrCYe0MtLZEzxjQWSAe40VQuip7K0H2iA709
b0xmes1fWuW8+ZjhFdfHt0fFPJ3hfqoLs18ZMJxrNxroHJP2xliHf41dk68W0uGo
KALQ0YB1hhtQpDGM6U+SmlMFWbcw4LjPjw1W2w5M1Wn+vqCjOwAtRXjQiDBTruI+
GOmWYsQJsNclv2C9QjGb1OwI24mbGV94pCS1VSWsdBUIH92eeqxlJCqc6KUCWhQi
tXMhxH6TqjNkSnTUefEOphIaImtdPrYOxoLHp2XjtmrVqUpM6LtIQ+cYksyPzncw
j8I+iaCNgAwfwgjP1iBp81KoML26DclS9QGXWUfaciuv+dvJcYSQjWWqR1GvCEXg
IwWJiGSlJsIGCWwkRj/okqNvW3cJrpr0cawxeftT5z3XF+1TckSGzbl8X8jQuJPP
UWgTVOZNznrQEPAA7LJeq4CbdbfHWrgVOUL53sosfqgqPaG7PglJPTAaxHZXQ0z3
6PbFI+JzVsRFjdY5uq/I9alGG+N3dvjjBSxaSv7lXLmV1qH9fL9ABflIRF39YEtW
dMR3sA+lP/kG5eyQHaqNpV1bCYd6dh0U0VHkY0Ok4S3DIQ+x705uwXuMrgMVKjqP
zmFd2Nnt2Xmlra0AGTbkdP8wnYMFvvjrMZSghy4Nfzuc3QKnX0nFt1XHQS/KV9D9
nLwa3SR7odCX9sr40FhAeNZ2BZE3vKifTmUK2QrZfVKrzAmMhqQ/WjMMIWy30M3k
pL4EnrRgN51yqbNHKJfkCWTimBBt8HIQP0ByE3vZq9tSgYp93roixC0EGpwNbrWi
9vqK39UTjGBsmpn+Y1rzH0DTD7fU0LinxzJLlqUZeBSjmVYvGW3/kamYJj0KDcYD
7rONneE1ottoropVuauh3fXFnF9bUn59C86LcbwBZjLnspAL15mCIPZMht+A1BET
1S+TJJTZDDWUZteZUqUso/Jc+kdTKDNhY3tJJO16gT20LkHLSeSvgF7YTJUMElLf
2bhmLV8v+dR/Ph8YTRS/duu2ZwDBns2MOtcMFgE6o1JGO3+DX25GAtYhiyKMhTcx
s+ValWoAedJ8cKUHe2iQnP0FjejfKFdi1Us8HfXDTq24hM0rOoyqOGNLR0OUb4Ef
2y2uBOYIs1+URqNzeHrkbduVxALuKvMIn7+Pbr0RfEX9UzezzZX3ngXVjHCeOXfm
VZr4r3u9nlVHWQ4a2+jw18+SFGJsW9jrEnKghn0F+Xnx9L9oAw5nnLR2IcPREQY+
hx1+IvNqRuhyJ2DS2/gjounkJ9hALKqC7vXpCpspkziGRtcqSFUrzDlarkd0vhAR
ySd0ygYsLzwIwkOvVrE6RGYPLpCGCVcDJrfgClraq0f0RWPaV/zli1Cf/4uuExM4
gKLjUIWrWTYCk/H+z8VNWo5XmZfZScUiAu0WOX3mNkPQAHinv0cyatYwBrbQzRrw
+zjuPVAcb6NYXV79xC36cA64w2KaXGphMfTbZMyTtuCI3ns4/k3n9TH/1uTFCdj5
Fzv5mdzP0Qf0svPCNSCuCtpRxX7sUNkWWamzQYM6UBYiyhxK7O7eQIvS4XwvdQeg
ianuNDLtc9aS/RxyYOye66tUtduWgETb9xRA8aWJkOjhgtX0ccJr/Q35MZ9DveBH
0UaZxUwqqRy8CAsExtgEVya7nAVX1a5f4x/OioIoU6EEYj6pIYub9XyOtiWUHVSe
vwFjoqHeHRDf8zvJTZjqhvSsKbVWOaZcC/hNLme/TZODl/pb7L9TcgyAPxtFTFg9
JzaXgwQrfOGK3Ie+WM0Gx+56PUfH2OyVQ+YAwtAev/GR9YtpWMjzcAn2xAXPZrJ7
IXFEUPMMhWWJVNLzNw5z/4ZiphyIVfIHGpGls8zwoHTgKxhlxQyeHZa2YVaAm1IZ
aVdx5n5KIaa4DR7IMiIu1J2JvEz9qLpkkIwmHu5HG0lX75BoJaR7VhYZrasGd291
ImJ9dL3/IclQ7N38JdU0Vu793P7zYx+kzREsOozopSrNF10nQhI6uvdTmce+oHBs
2UtrrjGU8/P1nL4tiJ3MOOyfwemWF1igzX68e8UsFgY0MTWvGTs2vfpl/Y34pViK
LjzdX6G4VCsmJ+gMqiQD1CJurt84dSE/3GaFNW4IFBbFm6C65RkUJ5OyYhD99pU0
NKKr6skkrA8nZVSrdzVw//7oBepUsTmRvRu6SORUvQgOfPaq6J+vJevHHa84DEsN
FBPcWwEfSARu6tjT8laXQPcVITs8AZsNiI9vy0cFkAiUQMfT5Fgj4aWOdGPw28YB
UrLU/6+r6x4+loQQr6lQfhgnqc9ISSiw+Fu1xGvFLizjr1m+PBSn0jmOEim/OpOI
ShLyTB8QZkN+UEV8rrL7tZOJ/LfS3VuCcDf2r/dS6yYKqv1QYnCDfnuogNdfi9oX
T9NHs0zNK1k92zJEoPA3Omoft8Xkx8RYkWJ8MmRKAbBJCiOEmwlnTIqytNkEE7AK
9GeZ9jOn5z20mxhfCloCw3nR8cJZKg+JVmnn+Y/2B2NW2leBZz2ohskkNVmU7zJk
8aK1+RUcHpHVLzAisvZLqeHsSRk01o9EmRRwSBeMacQfVrArqMZR9u2NUodG++U6
LSuBNL9tI1LrP2sUhvciW9sdvC+M71XlBeu2jsOo2VAsiAPWd53x5PnNMlq4jR6B
BKgEu4ZnqytP0vkltewQrDnERaNj1DR94H+sNqiyp23UvahXS86u0MVJePT2bkee
mKTWiG8MfRnwkPH2DEEDlT+Xmjv5+e9em85cWoZZ0e/MjWkQnQkM2SJrZOvz6aJ1
MrZovy5PZDC0GpEZ9qLf7z3Qg8+vNb7eZHYGOAnw3x9Os3QL8cQuWSPW8Ax0cwkC
OhRkvHq+P21Ww0pbDDKPJ0KllzulmxLei7GsRfWKzKPZAyq4tPvcZCiMZ2MrYbuI
ASavO+6LJBmNv8CziCRtHexq3dwpR4KcZPpcLZ7xZcUr4KA/g1DbE39D2D9lBsN1
hUsl7OlQLEr3MOmaE0FvZxjtQSTqETHmogIo42ZudWdxjH2rEvtnfhKtGz22Moym
jZpvwlAD9sZabh8IRviwhoJLb40CA70jmWp38KUmPG9B0Pl8vXu+niV3X8AWAEsZ
I6n4RoBkAKjOQFi3QJoN+Nh7FNADOLdTrLVc3Ne9Bv5ib9AivAffsfv460w58ghL
6gcrNNZrOV2TmJD1E6GLVs5jgjCEz2Jpv7qVo8/wnZMxUAyWSlNP4j950Ok0Lsmd
AzMEeECcoLHCAljePdmpX52fgK+0TvDTWADHelH3a6UfzaBR/xN6jfAyMxqWdXSo
QFbQR0vFzep5iZicRBt9XbG1UCrf7BEKn9r99neMCHfmiSZX7hvJLk7tdb1ktRvA
eNkV/9gO46G+x/s5G8yUWm3AxA9Xc2OdDr3AzTeZY4EXpVZg3ve7wUch64d9D3lA
N23ZF3/FcESQ8h+4kOscPuy9vQ1TDHq+xRX30cGIclcVD3BWFLiTzFHAliBMv/lC
/i4veWO8VzwsXTV6RH4iGqapCZmrRH+mb7pBMqXqX6ri3Q5fNxKPue23ME7VOfa0
DS6Ccl4DIg8RydvmoqcNIZxejEM5eWarBQFrnf3lStn+nTehRbHC0iALRTH0nl+p
teR1i90EQSzI0EkoHvEx464hJ+20o+z1nbjwtuHNTY2MMnMsRR/GlJaCr6fYToRj
szswJgtc6Qf7C2EX/CoPaCrol+AKceI+mFsNiAxt7RLlR1AE8vtEEvK6qWKaKYFb
9ceosNh2jHaLwKmcTPDjfS4yqxORRM+DZoGFOI0IVZWOtTQ5NsYQhYvNUTNVLx9Q
IDOhYRZ980eloj60e9lsXz4xSnTv910YJo+EDD21MdrG+kMU1jYriCjaAsTOCoI2
t7I2QRu5AF2bapFullBmatX2dvIdxfFHPlVCDQ1hTK7pOKg1aCjykXkf8PZQ9aQe
lW09v1EzOz6RmsGvXPyvzmGuqHyg6o5awdj1zGOSoQF9BYM82qv6JzVLcG3ubfGg
kdaxstMTiorhqVxoArVmxiZmFPm+NltQ06fphNqTHNekgBb3cdhTmnyg7biIo40e
NgRj6XSCnoFGDLOAdaA/XQ3GIrtbzyx6VhIONUPrnI065ctzZNFQ7qA/mBDce+S8
X0QKeTsvZ+o5FWO+7uU6Hq188VR5ehAat/QAFb3YT1sOAYYBm/gZvaX+bMNgI5/d
5hpBQ6Z26rAdevSppbuhWpbFMyM0AnQVDMpk7T9gta4bEvVY/T2xDQyuEhUT7Bt2
e/5YZK4Mhrnxwd3ID4YApgKCnyHodK0+7QiJSvz+yPDfxen58RdUGbX4RgMcwwap
U/hScij62Uw+XOq5EZhoTM16cXEyqcJySYu0JrIdgeLAlI1OZl47jBV2IHO2C+dr
OXD3fUg10/BGxOy4sLu9zBbzWXNHEvhG7XlP8kMokrOiTS8GHcqJM5MMHeu/c9bA
C/BrQuRTb4KVYd5I+1w4gu3fnuTpxMj9KLqDB3FvNwzmmW6pH/eNDz0FVuwhjMUE
owqvkHzxLIjEWMFwEsHrzip7Pr5Sl1ZLIifPDmuvu9PIH9n8f/aks/GwAL3JM/tp
rHpbImjsx96QqiwW16hno5rk3QT6KH1Men/6BTkkhzQuYIZQ4WViHsyEzHKzDTYP
twhVgt675c4vSlq6t6PVGcLgbOQibW5GlCxFkUZyJot/F5ndtIDerxafZbuJKDxu
HhI04rFOdgLsKHaw9FzBqUbUPGOoU59J4JTSIxg3ieEufQhimSmeFyhGmlTGrMvo
sMJQdLbLwYN79pMWjxhZJkBzEs/IPbHngJtL3Apx7tCuoN2QRFQ7lFPrubJChlK+
OAORZp4a0PZ0+Ds4bps3A67HYZb+3PqrSS2EjkJpZqF6ayygYMpKF1uAoj1CKaJ1
oxh8qtFnmWlP6lxUSMO73VoZHwgJnMfQEk8pqZ7+jj039ARs3SqGfVoBsRzBZOWy
GBXkvMUqYBhSY3Pzs0cFq/II3wJRTm3dR+XJfFY5vw7/mVFnCKISqrFpGXW9FwSW
l6BKKyNJP7+NiFM0AktLnZIdwyEL3wtu3IuwwBTSJ8+PC6Kw2EiD3yWBcOQp4O9H
OL+u/wnA20hJHtNNZq6JtbyzarlVpRJir07/fzsMnNUPEVvC2IbVJS4p8jZ4WbYa
KHRnMLkiz/stpcc11XB/ENEoA5svZ5HzdCctniJzO8ok0HSi4qCJn36cI82JxyBy
9QDOWlcjEukl679SuO50E51vBiwmeEItCNKuDxb41vDDuo62rCnkTVGFGlJBZFfd
OmwCkXUOGzF/qZg+j3pI34f8IHISLh5qc7MaUcqmq7De4kP1vGyiq42nnIWsrvJ7
AxRg+DVG7HYjXKjgYcr2PryeTaF14TaRGhpvwRvHZWwI9+gPJpWVOGWsV+U4LbAC
ZxXPg0NRL1N/o8zhmjsX6b0/1QhHalWzGKWIaOxm7GnImm2ibQwGvt456miuCwXA
FULUVRTwEkhvLS7lXYF82GmKxwP9e5BFolsDAdTi1MAM144CSOgwFSM8vnk/GCQa
w5IEdd8CLXcQaaOEC/YLk0i4qfT7vjnd9a52Tn7wIxZT7bOyayEjUPjUBJCpW7ql
f8Ac4gVrN3Dy8J9sXiAHLRZJDLF36BIps//4At5GMhyR2MC6TuBKxrQ5e1uwdQsH
Xp0rKQAcDMNy1q1CZ12FedzDji3EeDu/iXR/qPhKjbPdmh1OvTe/eggsubynuxIq
6jFC6PPRtoik0hR+i2DQp7SUlhStbNIS7/AnKscJP+gCv8yWPH14nMBmEDcCTHlf
8amB8VyJ/Akx6dRKa2Xx03ZYoN1FnZGR7EfUasIbHgDB3W7baZEN1yDZgelIgY2J
kDYzNAzyzOyu5gNpNmsIttWGVXjLUYcYmidkoIrd5gpXRuYacgvXeiz+Bx4OlorC
17dnRpHxWiWcBC/M1y2OO8OeF5Dum2R2LfmH689DaO2T+cuZkJNMryAEcF+NKfm7
nCAkeaXB3VlGzzn3e1xbb2rX6/2/UYBW3T+UG+en75q82eiaIHjno+gC2s+9hWve
vW3M4BWPFXfw9+BC7beKcvwZQY72bHdVQg7UVPTOFrJvyKQt9AFbu0b5zKOXQxA1
2TeFGQ/OLOCFdRgsjXrs/fDwHNf/WVkHVf74aZhRVebeE820CSdOYKvcmhK1Oiwr
loDPj2X1Md+ZWEUjl4pUiVYlG+owCZ+T2ZxGTl2JWRlXCRWM3rPuOrGlUJW0F+6G
kVswCF9uF4c3K4kloWem7CH48JzjsxwTWripOHwlbBbt5Ol2Abl3fjzicyDFkcVF
5wTjgq6fUP5qo2hAHHMVzXRAfpanOZvwj6avJDS8Srv1jCdpFvWLUgcBKa9WQfX4
xNfXwflEM6cJIGtcFqJv7xaYj+TDZkw3GHaPLgec1vLEalmUOfaLAV1ATtafEBQ8
GJkwwsFd5DsdREoqFeiRCVfWLvZ7pAK/WHMAl+OtLeLWiWtw+Jqead1QesebuOk3
94u6Y1zOwkvfJ0/1WIxzwvyPbgqQ7vtKEiZQu0+Oy1ayTW16R3nwRRTBw3u6s2P8
J2X14xAvQoxdqxYgqcgzew1/D3ZE1gAmsdJ0I6l+SONhDa7/3JHWRYO9Z08q6GSI
zfz55vTDNQgrkRe8oOBW39xddqq+jiyPIWed9za9p9CZxzAouuE+h9udfIWFuIdC
swPndeYzx/6QqPJRkDKXzoVQrXbuZKYpfkLnO6U/umnFZxxhLhvdrHYj5ya+C8X/
cmdEsNfswzvC2hJUVxED8Nucdwa02+LLc0cVMcTEVYxcHZv2sLhnht/S2Q2jCzf2
hQ9khDySMjpiuwgqrIL1hcr8w1dhd9CEf83kD6PC1P3dhuYDx65j1aMFndXbgv3y
l4WShKHsMYUHFI/Cdr1fILfeE4POZvl1LJs8Kzw32veA/2+5mPaY7sRN4KcwKQ7g
dBdGBleLCAiE7A2J0DiEr4Y/f+hITmYMWyoq3kVjlwtipWecAywHBhfSKf0JX63E
KfnNgmxi7ZwGYBzL9Ve78/uyBuec1dT3apevcImy+q19ZboPpWkpgUpcE2jEIPjU
HdsizG7Z3iy42VV89VwvHEi9hdTosr6kTwpwnvT72onQzr7cV7ZyzBt4X3UtFqTM
0r4kTE+cVwn2QJfKDELONk6xGgDVsJdMDEz5FdzLPUwmRAp6aJBcQy775Aqyrh7B
fa41yHCoMyOukPckp6VpxNVlN4c/Zs68l6Y4jQq0s78Gbim/djBuHFJIGCwu9xPD
zZMkK6Gkc4N//Hlpx2nKSVVaSdy3Y0rTB75BqZQLJWiNFtMFnSRGI5nkdXyLwV7w
2BNTLmDV3zO3hSeUiF3fTL7erMMSggJ+7jQF2VxisL4gTrG9LZ+4hhC3x2EN1bKP
qwwPKH2wkQcHkDVuc/o66SW+MaxgmYSRQ8AEqC9/7EIWIl1NqZMujYwKc0Q/Fqcj
NgHWVipG04742cOMJShuZ9TUxmx+Zd2N/zTbvGgMX/oW2pN2zd9mQLN2jS2K8q8r
H1kud7BHvIlurUFcD1cgBXLckL6/LDLC9gI+cV0RarvCgNSzRWgKGB0WaFQoDwPY
xW36aBDPYlPSuIpSsK2LXHLq23cisnVyUXlpTX0JOo3WLbNN7c/TcTfAH6h2G1Sq
Z7q2OVqvNvhNWuLOILtEBu8ThobWirgxewnXW0Urvvq8hodOWaoSXFyyEfnuNTWU
5VHfXlltDCd7lK8J0NIr8f0F+5e5qgYQyeiydpexkRM2HYbB5rO/QAGjgKaZjZtM
LqwRfdAmocImWznvlLNG+uw2XcHz7RyI3LfO5yFHaSp2fDJ9chcMxxzFYXUze7QW
R4LnYJVChy+MfeyqSh/5QAgg90LMXeQZzdwVCQFEM322OLB4IhzhATymTb/00RGt
Fii3kxR0e6nwgzsFDbTJ+gtz0oqIHQb5KGnMRPpeGOTLMsts3SdX13X1DYUsJEYg
KyoPOGQfx9eF/bScGzouXX+lljX4NqQMXA7XN4ReqBOIPeRakq0G0vm95frKD833
ZtbvbzwPFXO1RWaxDeanG5ZrMvvZanMR8ojda8v/8t7On8J8SXidDddGTMn0i5aQ
sCoEiLY2fleHAO9JNMSOPfbqy+FeiDz/l7uGqA3QmfIf8W2m0CO2Cb+y/sFy1w8y
f1IAvTApneW18MZ540XnSeNxFpbML8Ts3leM6KvdHFOEVOD2Px1kPnBJmW1IkSXS
tTuIG0SlDwC34NscycUWXcYJ0IFSUrbfNvcOvCGxdGPNsh4JVjRkmI+j4GWg0o9I
D0GFRN1IJgsILE21EQA/r4cfbOD/Lrfddhg/AlkR3IxpcnaVX7OPq4u67gvQb3Az
IU9Lo3BpXYyqGDb4O0bJCWXbGwuY+j+8M7NsQTqWz/D/QXz0HXXAzBnkmkVyyKSx
5Kpd9r55N7a9tNrATNudvcLdLFsFpldNKllfww4Bf6LEcvsf2S8wG7Yo4dY5x5VN
c3kIj/svhCvio/MM70pNN1hn2Q5Y+eRfuuXS3L7csbwjsg6u7GRpuPwu6rIN7QL/
WYKGab7WN6sZVL/oezPRQR3tivMQG16hC5i4ou0KXMuhmJK5ygUy88UoUfBrdOnW
qf0dY3Bo3IMcUl3tkaFl/SSR7UQUxdD1ROk3UmNjs/zkvUSaEC9kVufVkSROqamx
SfY45CtpZNOO839EFxyJFQG6rEJz3Yxf8oOKoJFakoOG+hsbYUP3XBWMFrv2D1BX
ydluxu8Ur1ubsBOfPRX+AlaAhyUhA7hGDnYtSKAD+nAfuMeN2LaRVzFVWMyf+euK
ziLdZfkDpOdQbfTlITurJ7XCsTPKKSq94s65jVpqRx3Z4A2Xk/VJqk094dyMuUkB
A/bQY/xKDjqHll359WGL411aSSqey4hIClfPwvpVgS07oCSeQzwHazm+3tRN6nd+
maixuHuqrWmGWRT8zdo4YDh7K5sCjLEa7rcDEZMY4UWRBz4hzScXwSnHPr0laB6/
Qt3uWuA56vTT0Yl2aW7aQyZCrXrgPDQXPdb/ORwGpLG1U6kFfwOBOcZjiizIOmF0
sOyHf2zTFRnXU759KYe6L883fkjzZ3fN0ptm4X0lhGNn9werNvs5eIn0dnZ8/FvZ
przaet6TrPCIfUS+pbZ1ZzAwrO/YLIVO/vNFZx+A1ozVurdP+VduOMaM9yxG6OUM
xP2JoXf2MlKnDJWY7Ihr8tczARXjnS5QVnL7vhDA0mPs99swC3PhpWGAVXe25P7X
E8/cR9NKltPeJpWZk2Al+v5oGq/4Vn1Gx+zUZQ+pnryS6UhJeafEVG500e+lYUeQ
gowDOXKtQK4esjcyi3TpgGrJgq2qyW0q+CMzPMuxrILgbj/OJqySGaNKGxAv8AW3
dcZPWJaLXahY4k98XlZPnBEGmrwEAnhA3ld67m1Xg5rLSvOU572EsYmnJyjXlt8a
yDnsOL+gWSjxLuVhUUVx1KqmZUFb6+93gGsuccU5KSRwJK1MmuLVALPDpWxenCeE
v42IHiLgulovoAwurpKtsowMWt/TApzhJ6GHMUi3yNBhLz8Zyin6WrJhD61NjqFV
4z0Qr8XsN3Tll2WWSmdFRaaEhuH3/zbNf0fg1gR8voEOLpB6rvn5YN5fanIMXuC3
AE0XxkBUmOt8OMBAchaMdIm80MLHk5Qt2MI1QN4lqLbqGEgNFsieYrCRL0K7/jMV
7XavNy3G0M4uk0HxAl2PBva9z/bvUnyEeOoYE8jRFFSmJdYSobL8V6/JWeda3Vpc
nBl+5tbG8LNfWvj4RbHYmL7kqY8v0G3DhORwace53itbnIkYnJtyz6Ue+3IXEOlx
ys0P4uqHIi2tl9fl12S457/nEc++xWxsUnBZQhgjwaejJD9RLRbeIpGIrM2kw9E7
l2mMsCQLYZJ2NXgXGA0MiYvNMHw1/XlgEVbT0Kk7a9N2SueYg8bcqAFH1jkjM1FH
bTiNhG5XRIw+0lCH9hhJLHoU6LDQo2UaALlsmu18uLBkVZITWpYDMW3zke4JnxEE
MCd8KU770HdmAJoazxYWiAYQHEzbh3WcNRGYSrOgtDlSYUUCb8VPlyG4JSNnIuhb
52Qc8qj+NW0fokf4r/I+uukv9i3/N8MPqmdsWGlXwJUxkuFr/qOtyUX4LgMEDIP+
fG2YA2zSIs16BHF/n0tEKnpJ/6MryDRcpMhi9myvKojxk3PV8/9J7c+GcT8BnkVr
ggWG60wLPsdAT9C+M11Sj6nqdQAX09DrZwBDhAU3BTWaqVBOnAb3GLA9N4Hvce7f
EMdWa17y24d2Pix2DHx962Qsv14d1fV61ibjUEaaqYeGianSu4w65fTyXtEB4/6x
ltCR15WeggHUXxax/40ufDieREl00jt+OppKtzWWVb0tQJzbhX5ocvqUR9VMVzb8
RLv9kJ3EZTiVTVePpcHVkXLejUUcMmN5UlpXVChWxN/jrOiA+O7yTi+sWXCEzEwF
OJngyUxfcWqpsQyBLf+aXuwj+h5e7DzKiz6d3mZ0hDTh8mFWW+lxMQvBNCz4LIVH
OH75DQS7vKGRXkPX4gYbd4c7TDPCIBlJPpU5eFP4/4rT7Oa/cHsGJo8zMmGqQq2S
W5Vqp19FN2qwMi+CpJ65k05vLLpUdcZslYRVPtscj3UEr/YC4mw31pH0mbTAYPXC
2luAMvrttpv5E7X0t/+SYjya7vD45VM6gwLzKPtoE8z1tbodH4HEeO2gImTpnVsY
CjdoQPOGOxxfdOLLNrG7PggMLiBhEEv4Z2FAuTeMvp0b9PZyLX2CNCNKYGRS29Ym
qLOv/tFBQyqPRShj5g+zmdslGar04dP2XLZBAfKlQu8JLLhGTqPWM/6OY6Sc+OSi
sx8IsLP0isDchPwGwQwFzee2/mw2bH2XmaFvq8bJlCxtYAPeokcSKZCzSflxCfli
BGkYIb5g8AUTA5WSO9l7zkyQw1nb3i9LIki5+O8LmQoZcb0mAX3XcY2qIVDQqinR
TD5+2FEpJZQHF5u9zuiDbowFSrrtcRzYOL2N+COlx9Rn7IScQjjrgCn7rL0FES2g
AWP9qFDXHjiEYn+ubXOdfZFVyz/it1r9FyNicfOyQsYFO2LHf0uqERbW6jY3/myv
47jW2bWyX7dwaTPKgxq4pWH8JUCWl68iNa3PQ/cUIz4WIzjn0UOB4M4aJ6ApbmlT
pNJTHoMz1msbBjVnC6p0Is9EAjahIdYfQI4mVW6X6CqQ9Mr+dRWB6dKreWMlxBoH
Bxflo+181VbQ3x8UYgPPF261DmTQ2CZaMso9sfQGGlkFVj9TwOqvsY8qgh3hWnun
Iz4mhMgZzgd3kyzC2mpbm2IzuxKCUNZr7GDnoGKGyznX1FjuYnJqunBJTvaNFAwr
6xsG+vhiL8YwyGNVYNYRGVEaoC+Qrau3cwLbde4VZPuIUkjXkdmaQJMd1vQwK1i9
8/xWLZO9O5Y6kNMzp293/bmbUazBUFR3H03CNz/jsfyBX33LQZekTSWOxR6C2k4g
tojwl2GMIKL4FNCuhXV02Arn0XoZE0ZH6M873Fyw9Dto7o+CRyOwK8vswZLMkQW4
KsaH6+mJMZ1vA3XWKYMHxQl/FkVyC6p/XpVWfjXpxUCgL167RTFpyiZvMLzsDCwA
F3ebtxqKbSzoycEPj3supZ1MXS1SeR+rILBDFqg+5yzIcHLjFgMb6Rdhnbe1G0bi
gZrY9ecxn3aoiQ2LPi1/IBzr1riSqSrz4mxCH6l4ta0vH+IS+GsW7AtPBr4i7mTR
zobhrNwVv6ZbvwDg+Xs7lq8m7jv9/OpcvzO4i9X8WXq1+ro1Euidm0EEmYL9RsOZ
Vo6MvZKK4+ITpgGBg4uBU0nevEFVuPgkDik7vgDdBNcX5a3ThiUo7R1MFQ6NMsHp
HziBA1/DkkqhO86FoYhaL7wFiTQA22Au7nwV79X4sZVua+L8G7j9uOXo3alSxufB
EbrEMplgsvN8PdSpsLPDlRqLDPzAnkYultxE6Z3ctgkMNVr/qBOgtf0V8ZpeCU5y
rHjY26zqnzWqIc3C63xizEeQ5jrSXL5QwGnt3SVXtoZp3b7dOc7VBbBoPmkZwv4Q
uctOw4tzrpYwwXoeUEf+EwyeV/Njofgw0IR7vbpGxZ6uW9BYXF1/7xqNwhtVtiYS
NdQM4OSx00HaBJc0pnrfSFtQiyz4o0F0WsisiMITA4G4Dy7Cngqlk1JssEORcC9X
QdN/5xJZVeDDqxYO3pBfWU05rzF3gngtvj7aIEsygNUk0vCxsGSnfuU2C7BA9sdM
ZpVgAn/DsyRX2PFWANfDl3FVClJAfNu5QqSsSj04Un/nOfYy1DslIXoxotjmyQxB
q1q/W7noJlnanvas6SlPrToUz+pNAHpZjCG0Zj4s+1FJ7OdF1J7LiRTEdZjKUM66
pEAdVjJ5oW8KbTpG5Nld3pw2pkinshQgsRJXfEEHVeP0daeTLlSEbjb8MWNCQJF+
soClnvAmzolVsszmDBM4Uh5JxiM6MqEapWomQGm7AdQvQlrtpKoEHw31kXxGdTPY
88PoDDVyyXlN1/RTIR+zOZJLl5vXKRCe8sbU6bgCRNbSo0Ku1+/ItnSk3SUYg9bs
95j6+ZPvAShYY6G0Ce69t/2BONPdqLKdrX6vdmUyksToDiyrXCTJIxUFRDnX1YLA
L+Vp/sKOl2dNMTHbsm1idKliSNkXuss/XWPYzQH7qYwcy5lF7jmjArH+OZXYY6Hz
H/VZzD8Zv2UwnDlDeAtIoHZuSHtWJeXQSOjcHSoHZIHICxeBHiq+/XFu+BmaTB6x
gdxcrReO0MiiIvX91Tf/i0VvfBR73X2OcFff2ZR2eTQMDC3bwTqrN45r19ayn6ho
6xy0r49oedHVvIhlIU4SG7YzbV23YolQUcX6nc90mGDkI4puv2VUyeOhnU1I2Hxo
Hy7wJuh4MAw87ogs4ZTNlCx6Njdc0KCC5+E2Zeo66EEs6SAs0tDXoAEBa6rdBBjl
P6lTEppelr5BgohMk7j3nbIlTnXTLg/JEQpQt5wZoUNIV4ke9E4h/aVMEWcyXi+s
w6JnvO9nP12x4nieEfBa6eOtJxZbSC5MGI3+e8xr6+1B068+GAKk+PHncWMGOEio
za96oRr2NBzp48JhPymjPY5whUlA4ftx58T7/qo6qW3zWL4UbSc6LqBZJbUSY880
R1KYGnhryqUZK1ksq/cbglaUu3UbsGHX/pwha0imDSii9nsM5sOXoaEk43VvuUSG
Zw/0A3QcJ9mmkj1EX+imFy0FtVUqzGy7kgfsP19ir/vejoEolg9DIE9xjDit/5tq
ptVF6hj41kShU7cnjNjOmmWfO9bdPDsBDA+nhGpcmluL4Ma9+RvQbWyR9/8HvM7c
KF+xsWcUY3gSM1QcGVD1suLM6iWqWDxel+EIKrVAUiSJGel9x+V24tt1LF0YfiBG
TAHt3rlgW3v0IH7jGAcp+z9y6FxCGBqp4yTxnmK6EEfvhM1CPn7yNZBb5Dj+fivU
Mfns3E7ydL4gCE/cbMUQGtadz99l7fpqPIiZ0kBMqglX47bk/x6uL1ABqNk+z5X2
cw76j7t6978rh7ehzJ+tWG55/Z5uMddsAf0UQww9j8eNxlnoQWlLlXDWR6QdzO1W
DYn+UmTGKwUtmR4siicitVo91WAGAaZaDxcDYEwjo8vrF1Zf74bxWrHEPbPmwuzI
/ggxiaNZHL+cU/fnY7h5nqWaQiw4/qg1RBfUvLhRJBmJk/aL7lMcL0AVTP0qCyff
fbvcNNcIYLNgmi1ATYtvXBFalE+GtchYdHMqkf/t0hqeJDHns3+E9HTYufXMM1ht
25ld0WFC6cRnA8otMVwHHy2gmbjH2PRTa+A1ey8UYLFWUSyDtUp6DHLNbvjfC6+4
yJohrzXTFkzYdsiIAgyQEUwpyMqymBLQ7Krb/ZzKrNmq3taydf7QA7KdgXu1T/Xv
g8BmixG7nEiv9i+zZ3BaLuiH3j0GS2GwxNyeZE0XTC7+583dvN0JIAWZPS4RIR+V
H6NKFOOBqz2EPEqrxZNFhuuuexU0Yr72aNIVrJcS0CFn/4EDEI18fQVw4EWwBwGq
727jE4SYpTNWUzWKimZ3tZ0xPVD0Q0GHzXFWxho2DqbN4MWHqbxk6KpjHKvc6YWk
JEBEStlKwCxCsUGx6cYAlOestAs6e4AQL9Hv8Prq0T9f276ONfRSzIanitatJl88
NQ2gKzt3dDbMTnbj+YJHcMbAAKoIc1LI5GDdYaLBypIKA7+U2Lh810b9rd0Oqc2T
8Pq93nhSX70KcAHk7zbtlK/8pcuPG/eRynGW+mD8HOT2KJCe7XmKdE7nX7vG107R
+I+/vXJ6xKB7QNMrp61OTEIeyFKWniu45WOJtM0bNNhZ3nHh7m+zXlqEBFJLopiq
cdmPabYQhzujnSjEit3OwtXoM4e8DotjtnTBGpaFM24na1ybKr61zt0fptjaj19N
I50re84QKhFPv9XQF4Bi4qNE2nU/49iRI+8+lQ424MG+cQq+82lHNjeC8LC8z2yn
JVvycSJX9IpT5nSORBNp1sWQZ3WCzdpQF8D8QTyRQU1M7y1FwJ9ll2e11O4sKylu
2D+SjQRgcs3PP8dAtA6xxMOCOUWRRoqkIZ3M0NJeS992QIKzrjWSJ8gYHC9GZzcv
hHi4+VRmHyLR+pRIFGxORnNZTb2aGpIXeuLpFAvnuwzRswlZlsuH5kjf35jMfMWI
EZGq0ZH6LgLJcwqRWXsquS2JsIwpQ2toTuLAgBDUnV6EoNQoldZS50GZ0sgHXOw5
NJv4MVdhnFl5876Zm1272zEs5Iyg7n+vO83rFXQtOYjFaBi0of6aKgNBEdb7JoRo
1d7hG7SHRf/B55Awpw+sLFNbsBNNtpc0g8KTSbOshbeZ+1uh/t526hDKGhIdV6LQ
6/n8hQDgDS4CdMwdQ1euAQOGbyN9hPsz12pcuyPi+6MVS5v/ZrKc++BaBjwpQlqE
T1ie2B18BbfVihKHoMahh5Trn7Fy/j70UKayfRKr0nE/BblZ08KnGhLiXJdD0bgN
pl1VpGy3tJdkqXQCkCIhdbYaRd/mQEMyOxrs4W2Qhsk+dFYa1YdCvXyIubMIYzRl
iREqyqTHCTwrPC7mscgp+2BA2cZTCHjJcF1te/TYIwBHloXHRiwfVNenKM+gw5L8
GjgfwCnsuU8yn6HIWyxhacD2oa16lfng+ZQmLMKiICdWZo0JK1lngPc8w1r9P2zl
b68bZWA2uJXrsA+hjtbHcYxrKBmFx/OzR/lklk/27MQD1Ot+WwJsWzuwd5TJJR+3
FDASbvFzvDOMP4rx6koCl9HJA03PE/5N01K9k3pWkFMHwmVw8NQTNTujfm2oe4b6
/L2qstbUwqP/PlG8N3CBb4l6mseCZIGJxwl7PgXronVE63b4N4S8MLz/5XbiMOg9
GfnupGgpaqFnGzc8EiGuaW2otVECA7EZBCClK3hPnz7o4dg2lQaavKpg1xg2eCqC
AqSQYwutMNWbBdxvJ+jeWO0MFAXspGDQfZgbExLbUGhRoOSfQgSgSPBATYx8pLyn
M55pSM90gyI/OMkWLFLVNhqGxLDJ/5vJyBH74mQCKrGH7fuAT8bAHzQCIygCnbCe
f5d/s04I/6mydqGB7hRmwcjsMMGEP01mc/JRVlPusx3kTlozqRyJUkvev6tEd7EP
asFJsNbWNcn+NGiaGXfV7GJa96CXnqyp1QZXUBMa5dChY5/5jgPKgJBmhziaGWEp
cqiXMBLFZuuAJ5WrJzdZGfNXocjd2hCzCKMrlNdm0d89F32IeTM0o0KJARrmyrUp
5vqrgCLuKX8LY5g52A8O/38g6jlhksD65oyG4mTtBnu4THTS1hhcbnravd3NJrk+
MjhNsPZkuX7+rWNOTamMc3vqUthF3/Gx8qnhlJf8sU6zKIruDtj0s2vN5NUYOeJ+
6PUw5By1G5ui6ALm/U4kMejCTflqF9BIaChWLOgrQ3mRKSGQd3QlBXkUgMFczJ3z
0fQ6Jd3+uwDa5ssgiYlaqSB3VnMU9/YIJJDCw6UDXcMSHtb5+fcyI2AGFO9/pADu
PCvVObEEwdibmImTJBKjjKEDZ2r6psVX9OIX9LgTubV01CDUjX8AEOubPtwHnfJZ
t2BKBWcIPUrnKPjz275rS+xi0PYuvJcuDAGNs6qq3/ki4vr46I62oa6eqQMWCzRu
kG+MnC8gU97Y4cjm4eJyznBLpAKy/IAAN7BKyFpSWNQ+pPHtR0RzlMuRBfL7ECjB
D9DM8l5HoDsGly5CHFyOrcTEs7zKZ9bGMxhcm6QXohlHLw/m4nqaaKJe1wyWAWvF
HfvsdThLITmpERhieOAV/AVAuJjKtyAiay1fB3LqkcVHYuOWn9KfDNcXumIXEEuR
kXOyzHeodbk2EWyE0QdY2B3DypHaun7xXQgcgFIbAa4z1x8W5/jfUVqx1rBmR0Ys
j2FUU9HBAW6+c2fDZEJLXxmltxEbPbrRjw1HKemcm2U53FDKeN2qipGlzV+GSQxJ
p805n4oUhXyPijVGMT98QFD61kdmHZHRbActPg6VvuT1b/OYUXGRgSU+DDyJ4+Kf
kMVdQNdtnfyeGz6RrXYfOJ4YfDGApFW4ySmNwd6iAjAMm+hVJ8DEjmoUJjB8MUFX
MPb9IwKH4tR4Qpv6SBSxt2/7TAZFeLXLqazV+NwavcNjWyEAM5PTB/7BqlEjd59H
xIjFgvT7pMJj1MJY023SXhP/aMDNotIRw6XFnUs5wKI+VxL5leAXWdubs4GHVToR
iszDKnKgOmK44j2PcP85t3KrAK7Xs2BexmQ0w9MnbjhA+pG5QlpX2HXSaNZKQM77
x/UYB7EhQIn4lXbU/bf6GLqyiAINIvBuFQvb+xVm82KG1Uen7RGPwd7iEkJL3pnz
HOqBPfuBy/UhlO0fl6m9gcHaB/GUBkkz2KqWgdtgWaKj0EcFqK/LluiaMAKPRIbb
408KcvbiZbUVlo56J5RFtHJgNmsM2L9fBLF4uAJjl3iWgS+cWw+zei4VJNlWhmtX
Q8jqaRMxwt3f5KP12Zu56ss6ihpN9u84yl9Ex5ao1k6rLQjYqJdT4Ee2A+VYL01o
V7HEF9W9HZWVED0Z+H8qwz1RdmT0NSTkQoxZYLTB2qvBpn82PydUEMXQmm9ogFD1
8FrsYlBLQ6m2ZnHXzUS7p2p4trg0aJcFtjtPS0MnigX48ypQY3/h/Fu+hrkcGp9Y
hqxZi0JOMUFl02UoprfEv8InAHZ50QX3eaXRwZq1h+4v6yqY6QHm+sYWV5uduHTb
zTrWTCu/yxwW4evAO8+4AiQpmBlgxWxpYs6MqrEThC8V5mDe4ir0qb28TVPn8aoM
wkSrwi4eyvlrmQ0Z/i4nlV6zfyxkxOiN9/s/hkmzY6ipx9IAdEKKKr1luK5xlJM+
Y3LKMK1mbz1ZQ2yFAlwlYl9J9IdUZM+bot/5tCe2o1oMqGalzibgnhLY0sg3sx5Z
yrt3gX6nCyCaLvDtQMB08yir41HwZHvwAwwAsksU9vnn/xTRxCZmUmFnXMMPzYjj
zMC8z2YLtpX67i5NPaNnoQ2t0C6inFt7itpN9i5x88yeiHoBaFPyriFyDz/q6wMv
1/r0hSYvyWDCJqCkMBnckwvg6O8P1tlk5UkAASLsbdEzNpbjB/gXNjXlzUrBYcm/
inh/T7gVJ93Q6dDhwYZvprx68ICkoLRHDTnZattcZv2MZffVRBkxDAQnQ8qVCHSS
Kf8BnfpmFJaJxDXPcQ11v+9p4j3wlkpFbbTHxLWu5SgybuawlesFJvHapSPUCWts
vFmoIMjf0tVKKQ2i7Q8B6jKMgAxgnzzPa/JEPsSukpdbKT9QwZ50giPirIZX7blF
36jprkBGp4w2avI4pDt4k+Dxy2zDJiVKgpL7Yn8Mq+j+fwhPXgOQYj5clhUtZH42
Y9EwAeGzftGl0ss+sx9exKbcSrqF5r05A+EY/vgCUzi+/a5SYvgUgvLKXPy5BgT9
tZBfrJ0kGi1JI9kGADToDIMm/Gd4LWlCeTW5yJnKn48SQVAa3Olp5kYg0LSnrrMP
7/BIGNTEhykY3Ye/aOF+EVVz1gh1VPms+P9i2xScmyEuXhbKBhkTR4jelU86a4XE
EMC/15uy56F3IRRSjJrRiCM6QQzVgYIDKymxTYJUDDaN81ONbdWDy7CHRmzNHKcT
Tl7JviCUuOfltm8o/zzCDNIAgKFKiRwCG8SoDz0WMtVJ+nTASRnYWDmGB2jQoAe1
EAbGAUIRUGZdR+l3k8nh7Kq9BcCE8Yfa33PMoL8FRupeAB6ljuj7ctgTZYmy7Qqz
wylIWx3iofVx2H45gYEOmtTTrWyQJMjZEgtO4cLrTsrCjMLQa1ke4Zcx/WjJl6dl
S+WxA7rmCOGqL5Ua/3C2O3/f4GzOEMqPtS0amYhBptD//fUJCM2shbYCj8D04VbO
dO1jd6VP7d3MashOfTjJ6vKpHseV43ljRo8Dzde/yDjnc7GfUP+ZfVhi3qx4mAcx
w71/znQ1Rf/V+F7htY1pmzyUUL3nMKP14xB7tQoRRvqOTYsR4n1tPnIpMC1Bb9fl
229SBVxDdWPBs7uXIPYL0FlEBL0/gCwDTBUKXc8ulrryjAM1O6mgaDlmxDHgWI/1
jwiiFBG8lt0HqCHX7q7OK1f6gefw3+FlIxl4DCka8Z3PbmBaXK32J2NoO1w00Ly3
xwUkg8XZd3gQVe+lmKddHl7p9BXMWTwTxqg4e7htrI2bqJsQXWiLHDb6U5HFYaC/
k+T9/VNSugQIwBhdyvm8k0KEmeyBkDn+xlfUcc66OdUSl9lUVGvjdSC6NDYOvEf6
O+9updezcfQ+7atBYEKbu9JafOrDl2RcdYABQpIxh8tuErd9gVPoGM3nvLen4PjS
L3/Vg6icXlJaj42w0c/x4YSaYH9C9BDtfbc+e6mApfpQsn+ZBnuedTn6xjBniqQB
H0j3+KZNiuxlcWqKe8iUd2hWISVSd7s/v1JFAf0RAUrtYWDe4T1zvj/6bYRIeXTQ
cUMpFcLFlxqu609r2KynBDZfolQiQS6F2w64XLY8towH6Hu9ikVcEVXrxd7xytny
sFVVG7kmGfAemm4TBGzLzaia5aMTHPGWnaSYwLdcrODuTO3GvBaQ6al7d5k2M0gn
WhJplxhXjsC9Trbjaxf8OOt1TBGHcOed+SvCLPX2QBOdeNTnxUOIiBkCoDPa0YZU
Pocz1jjum7L6D0Gu/e69dsUajcDyIIq0fodpAYbpGO/wFRWy5iism++dNXid+J2Y
aLx4n1yL9TAYl12I4c3MP7R9U0rzbZP9/v5PftjuSOEVqTJKOgeAWlEk9dUwltiS
H/jWrzocbt1PSxjmT6avYX6q8zctjJSu/Sn/GmcYgAQUJ5nHlufcXbo5DmnSzsIQ
35VEByW0DN1LNacJ3sN52WrZCLykYzMFbPNgCVZ2CDAFzZGmi2hwJe3oHAwYfeBj
BJXU8vZWaw1tXQsKfX1ga9tXRQMY/qfBFriFfaECQ6UMq5WYEPZFvZ8Xca+FMSDc
i9/lgb7uDGX7aCtcdqdWl7Kh57WvgX3BfM4gQCsd1WMN9q2t99EDT9Q2qaYNnQuo
RqaPdd1l+pcjmJhZTFwsa0VP8h27pF1ZRdcDpxrYs1tlmhRaRZO8eWabrQG9CNWf
2pKsYURVF1U7TBhKIfmr24T5TVr8+TnCDRCqDc0BZuATzASCdLZlOCnoMa66Nt3w
fKDJq8byXQDstNkksACLVSEYpGlruSCJ7YfcGMAJXPCgPlS40DFenaPdycdp5q1o
2vWUOsM6/KKw36jcNT62y9wZfTE8n8a07UxNcCyBR5PiY+JRhk5xJhUyR3i5QQCL
m8dVvfL7RJeNmvPAwdhpAN3yqUchTMfXzA+urW1lfl8lY0UaH9qDoTIVcI7czC3m
/Ht1zjm0AV5kw89eF4GzyIcpSEvHmLkGsN98rDk1X8Y4cxMxlwJ5nirP/uzOGbTa
QiqjbUwDj0TXIE0/UCdWO7s6AxcyO37KWC71fsbJ8JRA1Oi6ufGjXRDz1A9gfukr
4Vw2chLtRHMo886o3se62R+KcRupKcoO2jNUCAGUGxcmVclAnHmpJSAlG58svU77
s28OD6rPuQjkiqkxmnWOI7+I7+MP5NqjvNIJzGC3memGJVmB/3XTJUq5emMid1mX
6+Syk3Qvv0+JzxE9olGgKnSvC5l8lu/E7s/MNKVhtL9USpgFVKUInCuAv8UteUMp
y0/sOYi0QFdtxr4thcA7BKvdTPwsoWhczL8me2oOARQ53lClW/aiDehoiTzLPpJq
UWEmqyxZpCn8nRdnFpz2aO0HYwiSjjcSsl8dUpEYjE57Ej+LFIFtQEIOYszMiGX2
P2LC+ry2AvKVBqM/mcIiyMDK+PwEf4F/BQyq/toxHwcgxZ4jqllp2nxJ7tFJqd+g
QtkMZgd7yg0vNun/BGgLS6wWdwFBkc3akRgQ4V+rBNT/1BylCGz6sv+DEEYpRXch
hIm+U4kMMw3toVbWVXNcmZ6pCCfayiSmF8hIdkJPnYNwtqngUEkNybbSe3r5DGY+
yZJJpIEfwz+8Gr2qa0ZL7E4GxeG4PsBR+5Enn9xeJsgJM1LoBYYUAsfysKCMdmON
BMVSisLWh0XtGB0vrWjY8noC6od6QtSkHRxMdhvLV2ZU3KkXTHK1mbHHO/Yll0/1
mJCrKdDkyIFXOHf0M9hc/VS4EEnhuY540AmNI8CY6Q/x+ljv9Z4JQUy6XaBiYveD
AKT+in+98cX2m88PiycGXSPlOXtPa8CwuWWSTlWmwGyingBoQFQYCA66FBt+qQQ0
bYSMebzRnqVQ9S9TX2DMuH9ID31UzrFH8dyUXJQ9hSjhDsA1qFQlyFIgtafF7bt8
tvmIgDpA0zY9YzzKBk1lQRvsUDvnGjXHOpHUN99mnQG+hvsdbL4caFIt/ZVbfa7S
uSS8OfNZRDkRfvP78BOgNdYfdP8Tp3dkE2QD4r2b+6RCKb6arh7YW4zHFfvAAzOX
TReoClkirl8YK7CHtHYQQScyECBIUYukag0ZOnUXXeQDpkdW1OH8YOPhHzoyjuPA
j3LbRcuzjUl93ekGjB4yitkhcnUdnGYPnsxjYJTxUrmtwlLA5OVPgwKdCd1jDKaO
gkCBXfnILvfkA9j7a0Ugome2S0DvD8kJJfzCkofvgRw6rwqBOU/WPNjlx9rdLhMG
aYoEsCf9d30s06mk0Xc3Ix3VzEbXhjrSn0xh1q/8vDhcl+bTPW7bQvQKliOzy9/F
NSdKrLPCJmgnnFtHLwYw7TieBhYL/nzcvFnB3/EkAnjmE7uBprHnmohc5sPNEZrL
ZCEmGkb0SkQC3HR06+ndk01DEJiwz6QgNyBeRE/L79dKb0II/wMMs/P0D9y6JRsN
1vT5sLJYOBveM8ABR3hXiyCjl1PdX9W3fRYFAT7OFnZbG34ASFNU+W91i/uWKSs8
U2fdSmtaImyTNJLaRayt3sqLJVMjnZxR0wayfEQ8hqvjdALDJEZkgm8kEQrfLb2p
pVm51uq81/wdgSoh5j43Yn1OLB6DTfK8NTcVSLYo8tK0Hjkrrex9PJK3xhoucRRo
Z0xfVaTwn1+scB7iSpEkZwrFpLsxNE1+s2x5ONVe8lBX3mqIPm848DErtkAxZYbS
4d8ZMCtG4lm7cYeB7nuMf8H6QIywa8pHdYrycbYeIAA4xEdg/oK2F0UYbNJawIJT
RT9Ww2qqP6bi6vwKGUnYGJqGab/MSKqxpGIra0QuPOh3JLPVlryUmKwL8bAG8+qg
uUx6fBmo0CQ2I7fUWt1xZpi5QeKepVu3f/ApM1i73G98LwjgbxBpaaLwalNn0TaX
fhWVzQ2omFOMknJxuBKwH7L7nKitXGcI9EFziH0HW0NsGxNUNVPRGvpEltBwfCKP
aQqbSj0pQXx8fChCsRxajILHTPOUknXhsGJ9+XGUWN1zNGrw5P0QWcEciKC9A8oK
jKEgQhDnWf6kMWXEKGC0JXacl+4TpVCEcLPiijk9N+TC1pmot3nxN4OsOoBvvTri
1ZHTURlZm+pn0T+3UxU7h6hMEp4p5EeQYT7Ome6ucMk2Q6TgEIEM9mBcta7UII+5
YQoG7mJaO2KmlBNWJ34cFUPhLe4uqq07INhuiHjeIrHm4TnubxwcMduVU601aG+z
vaeyZ9fMduW4F3dcxMMC1kyI8vveubIT0rF/r0CkexNZe7jliL6hK3hpAckHtxPd
7UA3ab5vAkMi/leeTesO3Vz2itCx3h6lM1s0/bo8AWV95c7VYxFMoKqzZ7r+lk/d
ypuMOEUwQFlY2H7X1UaXsKBGc6GjKGFzzDUH95EV+Lgd4rn1Ues1ZtjTFO2fF5UV
u7MrrFwhbzEM8nwtVfl+buv9j5YbSuDZBtZnzttkURYCW1kyv4VwCWMBTEf+Inxr
fKJIlzq5pAHvoyORHA3ekoVHe7P2MtF6fM/5skwcX43gnvzEyqz9/UAOEv/kOnzy
MSSwQbtupjjYmHyEDbp3x2QD2J+2/xWDlj/3wj5DmGaU/QXFU69kq63XiQaYq0lu
nSd9aEbFAak/lcml6wiPNNNY3O+do4OX69POiGCvuxDw4Ke51eNEuknxZYVF6BQ/
DtgjP0G91J68DzdT8ZzJS6gVfa1mafCgqpEve6Y4lns0/77iwA2/ExepQKl6fCMW
haixMv/QLX35Fa4qJb5PJ4hl3K7YtotcUJRy5PDz2l8pAcR0FFTOqGrPWoNSQLBO
8kvcHpQRdFkUxIVwDUvj3GACt36cPzEGru5QqHEVppOmtdQ6PwM3B1Kq0rJImVIE
p4b3NqkjuTq+31THXNYAyUnnfZi1vxljH1s0n16gEJCcoU7i1XscCNc1PN80XN5y
P6fa2Hlkqz548/kgfNN96nEW4JoT0Rzsu92ieUz7ZauaB/puLt6L9tIRwBCxJj7I
7Ieceag5Iy7WY3eAuNuGWQzWW7OT3uQrkkjXlVMAZDIQwWJtFPr9dpDxrmsyOVjR
ws2HO9lvMuRc0Qjm8hw5grskipkGi3nXKmbMaHglROUI7WTIue40dih25yP4uK1+
UbfK8zTxWT7VARztHVgpz6rapVnbdDbVZCL7NM+lOaDga49IDWB2I1MAUkbEYdzb
XO0QUoVgfVxnTizlolcgYt31PtcP/e38/B5NWdPtdNBJUm782DqBPawVP5o3VG0k
i3wMpNbHhch/I1tZJfk9by9wSE4+VW0Rrg5kkOvccvavw91kEfzIXWZaVSsW/GYn
G0WaA6VmDBXdGDb07I51l3uH/eTx2mLBW5nXDpzKXIXVZVjZOvyX/LV1pvu5zogg
9wBx4kzzDk9B5Iv9SitCXw9ctD/KeO86pfqxVy/JhTnQx51FsSFuxV6rhyNqHQo0
hcS66pzD3v798T17B0MNKsP1qUaZJSyE0ajszTyrB+O/515n7MmKjY44Dr49oNe5
iR6W3GEr1VSxBRoRSL4yiQhReuAeR2l71Uc0CgdBWfteTrps2kc3S8/KR6/2vB24
X6rM+srw0AzPyabUJ61mzgsdaPYqVAqLu40dnee4sukuy/N/m0dWT/j+djkGKEve
c2865REmF8Y59Yh7c4tfh1m6vu8fvVWtFXcnHyZsLtOSeAhSP3JSJoRPD0SfGk5Z
+M5rhpenyBxHkmdltLX2Vh977KD9sdZK1j4x/E1mjpGvicjQ466Z7Lagtzgtf32X
WgzGRrTuJg76SNH7/j4elMlv+M/DLuSvbWpCPB3dADkpLbN/7Gw8I5c5aobAi/xj
DCYqGpuxyZ1HuzXX5/WJ7R09Q44YoD2GDc3WBBOzcYhJ1u4L0VwS0kNlRIHFYzxO
dW2kuybHDndLiOfLTcZMLdON1auEWTXfFtq29NDArj0JPu26FF4vLBAo4iK7xMYj
5UCthg7c3ku8SMSppkxL8U4Q7LbxiyD27RUl8Pg1QxFlrVXtbYPmDX+tcSlYkwR6
+O90LK95ASSoILHbMTyHzK470eDw1wbnkaeZmkTdrmpJ4SdQlg3fOyRXLsuq38EI
RE2U2hh9K62EDEU59xk7lYCa6A2f23iQD+101AddmH5U1uR7/9RaBHMOj+C8CDxn
j5hxjdIBT/kw9j3I7WDiZhDfx3PnKCE5c02SkT4DFHN0IZp3fdPUiaKWcghU8Vui
AdH6PLKo+apXfCPFjsdjhLm6Hhrzdkeat3oc12ttcWyHFf6zbq9iE5YrD4VWLqoh
NRc0WRL5EAiLr9WmY01nugclhrJOijG/kCulecMqdtWb9z21Ws5YcntqWQVAE82l
nJ/3m6xdOqAoBmNbTK1Cs7uX3QI+JxF4gPxvpnWXYULQMH6lnVZJOHyjfUtTswnB
NshIIMXlz0r//JjxEXXWrZx4Ze3ZbaqqdF8fDrUGMek5MMRJdJf1sJcAKNIhAk1J
EdHispkbrhd8I5Vhw8YIbSxca3YDhMBSm353cQt/+BUuts7R8dhOO/TvGVX3Vkn6
88rRhRNEZk6zQTnnJ7sLrudCfa7NG4GYs41Ld7A/Q/pLW18ZvL3hm16PMI3ClRU5
7O+S42OWJGJrL0INM/vnT9BGC9XPsRzVTaS6H8O2uAQGy0RbsPMgpwWo60udSzQW
daJ6BqYmBqDzsool1zz35wMV314h3mWFgLeN0vAr0Gw5DzohyrXpN3MTpyg1ADKp
DruHS4hmo9ysnA7jyk8c9iXWti95jDswR4nXqcT5FEJDFExrEa/Cbd/VZSpxCT2Q
srSTCFOChEensRKNxz9MeyFnTro2W4s57jjEKGotbxyqnFZ3PCc7H46k/z2whjA+
kNsGzt87CYX8j1xBGhswYPeIsLLX012zySmxG+v8XLnSVJ+NklBZNbhngqwkEd1t
CBC2zB53ukt9xZZwBMqs+yxu9Atnn0Zlx0xjoVUKXRXhgw+AqAetkCyDj8sWl1+I
Mv/EYx68GzHIbsc2JGOVQ2zxeX+zWrtGhEWCCgILDZvL++QtToq20Z4gIRUa+AIJ
stKL9sJcwYkYihb2Gbw1Ahf3DjNrAKkK44C5DazToUqIueSGJBxEnjHgoKifybeG
mkUcRkoewwguOr8uicPsRWCBvEH5pAm1cWaa/PyzgIQ9TqkGSdV/0Pm3L2SZVloN
b+fOEVQbutYd/io0iq6a26zsQwP2VjIoNCCvIB2iBP+dyuQZ3BWdM/D4NwuhBeuK
7nYbb4+3B5rmmXm2OMeT8rH5yZzhDiewZBJnL0KHdQ3WPr2yPMcUg9lX/nTdpHj3
Hnn85HXg3Rec2hdNZA8oyeyxev5Lx0EKiIXQLOy0b+csCo1FDgFRHfxJwria9RJx
qek9/YBNGob7SfCZV8Ype2ly4rraiShsKcqpO7UQWIyYgs7567ypdEtIDbKGU9Vm
dkkmBNIW/oO//wvYECFx/1oXD01CM9CP9Bfn4U72bGuSyIn5ryL1dOz1wvQEty6Q
axwOvptZpL1CV57FqtY+lMzqSJTjVpkcoGAzBqwb5hTd21rl8ed7WHgp6qDNHDJH
hCRoOQtoVc9KLNymFeJ51qFhzgDnqjLyaC3SMa5VHy1nic4NndOLXdg+u8Fi1r9H
it2lUI8sTVLqxUI2mp8lXzjSh802jXrqVPYnuP4lPYU/E7JQyhgIcW0OXneJPkL3
d01fYf5bof/gP7rXsQtosZZtEB7p2/wm7EIc0FePenfCxHaVCUzKZtPU4B2Nluh2
hOGpOlfR+IEixP7hTG9ACiquzLcZM9wjOi3gGYJvXte8BP9lonw+W50v7C9SJi5E
yQoGXAm3IFvhvSDPNtlbKl2Xj6wuXebN1PzNgs6lGs1R0irPY0eo8LqwnlVVDmQl
wTMqwbdjBiPUFNDA6Bmqz+8NKumJU5SJEPfyYAp+idj8cmS+G+uhR0fdOzLmzb7F
B/PAn5jTqFgwU6ESdqlkLUwIoyEqpFwL2Rxcz+h3XNh+fMQcwEa/kZJdxVeq6Mdx
nveok8Tm4m/4e9R4+q0PrxJzSgNrDb6v0ZiDMOMGVK3pk/adU1lnfA02ZHYyIVKt
FPFCw6mQWFzdnzUCQMIsUeTgqpSBarW6thF3h0HAilc/fBS3PGUVzltHC9QvaKkP
9llh+2FPp1ltuDosrWWRoJODpANM/QLWnAqQVU13pP+1FJEj3UX0C3pNciOTjAiL
tLSlP0PBrqvIk85fhLeNCWrDeu4O38txbooXGJd3Ej0SLlpXFmN7985TXejpo2rw
axB5knM0qAF929PdnKgBXkEnJDWaRGnHLYgUVjmfxeQx6BzCbnmcJw4VtrOgFOKl
sm8n0MFnj7MTsNrNuRzxSvNH0PoMqXFK958NCi9BytxRQKy3aPGUlP3Bc88TLaB6
pYTf0BMopRy1mEIfNDco4M/5vHaeaoVMhWUnoyenGyVV3fsvF+R4+9dC6l/z/A8I
+M4PBS307d8x0kutj/oPXcDDjGLZP8gzyDMQitY+67+GfXWqdbVadDZifhCSqV9q
jLzBEFzw1WGD9QBeLkAeILFkWIkSgNDhA/Zv/DRxyBah+JZqJtXycxcpN37GkYNc
NKqap6U8Zl/FE/Rujv1SnUFPS5n2qaJdJhkR0/nWjl4F/584l+bsh7FCVUUPtOnc
nwAUWnXGIieoazKp4krvdqmLKjb2sOm4lpyykW/fkH0e3i8uOp31vw7A2MXOzQNO
1uiAK1wM7Zkc+MocSl9/0oV0vroITLEGuoHOSSItNonTzoqBSqu3Pn/ibGlCihCZ
Lt7WCddvdVpQ8wyw6PCe5QzhpLIALHRpqOZ5CZRbCv5zfUxwoPgsiRupMFsJ60GQ
gcRkuTllHbeCQgCGWcuPNMculdopIP/tAl6K+8EaE1VpK0Ffx/vH5U3FxDXXnZLD
NkQIdDMcbBcLYLmuumsAyZrxVkITjHsBPlXQZONbUP5DIl0j2bOKBCFP6TllBe1r
NjVf4H1+vqWc2xYDlcy255qNp+wdcy8pKvHejDg98YHzKlKmVt5h63MHwnnk8kne
I5UZ8OE6zD128JjRUz5f6rK16qM2ncovFuU4rCVA5QtBTTdZ2FhaVm/AxeydQFcA
Ez5xN6us4Vudn8qqX0JW12GrAWIT2UeC0uDUIulmg4lIKnt1DjkLMiKJIZWdWKzW
2dnBhyKy9GscL5QUXN1l4uqAKtr5+iPQctuz6ptuHre9/Qdh8RxSkEp6wOoaZTSv
eWYYtu0lSy7TpgBdGtUyCidCSqUOkl9gSUfQ+POCwPe+ZXMX01zuVnNZVby83EDg
7Lv0QzLmso8ewScH7GWmZoEFVLkdQ2+DXce7C++kCv7kmW8v7cAjrkdlJ5M7LcYu
ls9B61MLKAU1pU87hSP7wItj/zt9qPKTiwcECeG9c0/spyZx+LLM0XPH8QAneKAn
mjSMDTJQ1zZZjQwWxNI7gw1Oyxq7MXNMcl3l/pjd5elbjgUvX2yHzasRVWt8doEi
8UPHsyTRgxu1CvRD/sR8LvJtyU1kkbzyouV0hWZqVVOROlQarA4X70AC/7s2UfY9
Vo4SmyvA6TD6YoZ0DTyfxdhpmkfYOaYIcMpMzywWVa5/k0/ZA4WT6Rk7kVQGRhXl
B6Z8RkgweAf5kaqoVPN2v1qshUgiFPBY5nOiwlxyWnlDyG/uHrCABKbRxebiRvK3
ksHDD3nXjfo2Aych2KHa7Pu9rXmyWHpS62sHhrvssjQiY5GS6RdDnl/JioQPba2L
WiZVAEA3J+B/y9O6Mcb6x0PdvNgdlPA2IYCQgtAHKPdDpEpjs9imdl5vxeGOkn8P
a4wHZkCyHjZ44g6oYtPvLR80GUFKjAvhHpGhdblKC4FdmMAw4+OhHdd3AIXWcxA7
pJPa13wYtIgU9ajnuhpZINbk+rjVDesHf1m/PySAaOh0ZEy/9XbD8tUf3pf2j8hk
T0SzYZ/JE6PozkMWXxRTf7+GGOk+WmsoXWxSECGtm7EyNe1zhRpZL/Ft/GInTzvO
pB39UG8/GDqnJaQ4e/5SUMyGl0GYM10y42bsW2KgHAP2N5/S6WuFy/9dvtjfZLQt
2LkmAYPA7hHLVOO5+G157VVJwnOQLd3nhXI9Quc5KMUsgR/tF2YeAOiD/p64dylt
J86kiVvsNLeDHCsi8E6GwP4M4jsClM7QXKGcaDqvDQafm8NEPURKtxVJZyguQE5k
DtMEJbi951VFhXEAjX3zWXSP8gOiuK0z1gN64Y4k3p8f03bFqgfAMKyU1vvpy2ye
+6eNCwll/3oGYU1h9FddCLeO5q6mtG6NTwvoJs+wC074sKvz9KA5MJjkkSHjHRjz
B2Als1gOiBfbQ/ZMOYfUmrrvPZJg7I00Q4AH8wOaThh0UU6IInCIZwrFHp3Yrr4I
3nmHVUYOU+8CO+Cjho9w2xVHfqfNnut7sHjcvSNvPWey3bgIKH5Vul0SQAvoBP1G
beeb1NlKXq98oGshksOIRY+7UC3cJzcenOAlPeiCwZ2EvhIZjIN2LtJHJpEMAHcJ
px0cTc6igahDG2E1q48Rp8lzdo/tmz+MxmRsk4qoDHpaS70TDQftJzNsggnv72Er
RzP+BlKO8jzrxz28Q5fhdfz5txGUWUf73pYf6eT6U2fmoW5tI9LOyUy85zXMLTKF
SJexCh2MbTc2kz+LZ+jIPKCaNSi5eO0Sm/wad2ESeKr2dGHdUgsIjl/5nwmzUUpf
Mad1RzeHdsGJk9rSYr6Okf9Fr6hYxSOahF2bT+IwBgHI5iU6d1xWF+OUTb1NWkrV
11+xVE0bDDfHTNIlN723xM74wztQGiUskC/6g6umR0r96Gf/ssVr8hth30oZdmxs
a90HWrmAXVXD4M07BAqoWm1SO9Qg6d86FUCLtCLLLAkkf0j9qkZ/cuVlyScJWaRa
m/jtvwfwTA3USlbI2q0pSh6IWEeO70ElzKzMTi1CQAVxAztCc1lFrHzMztzTuRQx
fXvefKWtEIWaTJdLRkoMT7/H69F3RhUKkokfxzNxav5db+LjLHWfAG02aamKK3eW
9+ZASGSWl6ML0DDQEmbzFPVlfDXjVKe296Bfuwu50fRKpMJ3E1E7IvpuM7jD6Q0D
44Xb5OEUag5gSGprKzQDxUC0pK7POBZyA0gOTP+ItVXJgjK1gD4CFBbuODkQBXL0
D+LjOVqd/RI0xYLetjA4vGqEUrF7Eo3/01l3/HLaF7CPVTQzk7JRE1JLrh+LOgHo
fNSRoxk7idjWE8q15d3nEuNmUAQ8uUolCuCdADu8ku8qGr4O5VbmW8QDCgc2HN1j
0QsIRuaI2E7HtH3Kb8DtbxWuuhquyBpFQZaonfr1Y35wrUBS2xxN/YpUVqVY2fEx
F2F/NwPBSFlQzAYBO+FUBxBFi/59CnkLg9+M2+ZmjJhAZdpXTCWtpe/AxjTlzrpU
eOgfqgQSyaHLrcUdIxUWP045hkBdckVEQ807U8ocTGLWINDO5DyRRwx5AjUpYMsd
/gdwemYIbWLzN2WW1mEzkmnYcNbkUQCfN5HdzyvCGeFs5wmb+qU1nbcj/DLx5QHP
ifKgqvQgeIzkAWGGZM/yhQjErdyshHVqVQXorcVv2Sa4PPf831t6YHlsPqPZ73vD
mVBxN0h596sZ6bx9QLrLxSTuCEhVoliRBgyg/kBD9Jkg3HoL4eyPtLWdtNF7NDHY
qU1gxFQnkD5+qxicxalmAdAG51wbJ5/5ZbJKvyM/8Q/tfShmVLunlU9EJAU4oQC7
KNkn54aRqMtYMDdv9JIDKfPbsA2DWqnfyXCGXi0PbRAqoNbaCMUdN/zbipORsJ1F
xNvthlgiCrVf3l1zmu7NAkhtJteDwRFNIgDFXZcqo5pOpbbNMsGa961fn2cFKgre
STKVoRF9LwmF/r7DaN28Yo+VrD7HTyHe4cEtmiVPR1RWsuqMYnmzHGcMNWNVdj+g
IXJPS4EhIzf/s1XE1oQQsCtIi63ETvox5YZw69pMov8FSsCU9RZkV2EmpJ7BuoxW
xYTnUC+YO+zqneKoCUhrY2s9mHSyKbRSzGbpPJujhbXtTi1DnrjYtEDBuR7MMtKu
jfzaePcb0auv8x2RQ131yW7wWNGXqovnp2vwnBdKYeEzUyl5xS1/knsg7l2cJsZ6
6dUpQF5kgYTWUJphzCgI/lYDgq/ZeE7jQyLuKpmk1CCpW+w5LCNqeN0ZndzwICf5
+TE1af/4i0UCIl1nJztcl9CS3omqBmJjQFVBQkDzQYOaBsnDidBgeamZ8YO8cfvh
pHnSdY+gvmBohVze2SrEV9i3oTTFv0Xun2Vcju2UQcTJlaTlg+9B41/Qg2taHgVN
YPgvbhKax9OM0Ft+4STH62bzvAruXkOP/mZYCXiaOet0tNOvo0Z/9GMAdXt9//G4
JuYtpqsQPWt3GLAj8j2JTlqwriSjjX8PivkDOydKeFqzQFiGrdkM47AM220PS8Oc
Yr++TSMCYuIoE0gladGRrCcW2Opl49Vln9mR5JupNm41VXvdc1dzyTruagPcvrGr
JblMrKxpTS+V+8Yvi8iD+Q+lZybMXHXBxqgpRwe6w9YyJvpnPZrql33s+Lzactt7
TmmiuoTBVG9luGMOiHjwnLEyl10xk2DUmMEbEhFNzKuLNaQwPihwuH1IPBlbfJoJ
xtWon8ocwbtvtpGW/qv2TDS5v+vB+AkLVs7uWYlGFkOz2p8KakYTuxGzWgdnIFuT
fjQlud9SNbmHp6ymPOUfC2kZGZimfKOaOp6wAkEpHbIaV9PxR4RSNWA9ynOMcPiK
SanLUDBqaoJLflvlWLvEhUk6ViioQr+P2XgMiixnthHPns6llc+3YL7TD7S+8c+M
mlcog+I0VKMDErqwxRw1THrQQ+ilWO09usfW69i0huiQMSmX5d1onhbz42DhShXz
O3ApKXPI3xrMxYT/PYrnyE5rDq4B+Qo802x3zuT6/CAYaBKNrNwuA+nxmzdv9m7g
6bWc63ScCC/iMmkofb71oeapRKbqtaGMQ2sslsnD+FeGOIqKQjtVPIndG+i9k+M8
a1SHv0/XJOPRq80DxBbQkydr5JHYZWaGCZuCuk1FlVSntxewAMDbbHp11Pfke7gC
S6I5OJ7VGGm13xjy9aizii9czLtGKNw8XUsqn2tPhlR8xL5bnp65PE+fcME9EXWw
PvLDzB9NBIxz/o8zl/ujnROngJaq7vP+8tihhS6FJNMo9CDHw0umeGUnZdTRLUpM
EjGixFkDmC2n6UKRN0in0IhGXolLG3uqDH14KZqXKYdl+LJycjdwN31v4djLVY5F
AU95k3OSrHL15b3m2AZwB50InQ6EOfIMo3eGxkjmqf1Ib0Um3w3wSBjtgT3FAd/S
YVsM/jn1JNjwhN0lLe/J/vaWiqKjmLXy+9KqsIaAAFFIGUX7BSiz0Vu6Mss3cq3M
m5BQhJuEXx31g1h7mfnU2z4s9ycls+nu4apUqI62nKMQOfXcUJCDtBOB495+p0tn
2YAd2UWWzedTEP1Xrx3EsJqILjH5DSJTdMBKe80ldIXMEW36OXy+3mHGqIdGQhqb
zooc/S175GflQQRGNuJ3U5hI7PZqH2uHWmLsZ4qMJOsPLeDoh9XkMlktxpLkbVVJ
tzggE81zcjJtua8NFECl0xp7PFz2jIw0L8B2TZgHDRhICCQF3aN+hJUI4N5lSbb+
EUBDj78vN1+MskgQKDoTV4Tyc4LSNJJyxylkrTbVvL4Ubbijjlq6nGkD8Iw84tae
GfvJGU+boeeiwVzksYnv/wVpmej3CJpjDBNmtRrBqUYFxIomkrE3truTYLleOJKO
azmwPrJr1EGy2lViiNsxE4HK2mjXfFV5p9qPRSIZHr/qBIY3r8fVi0BsmS761+nF
+rHlYoU9IpKC21zd5swdxvOSbNYlVmfKavSIuQuIVg6FdZEHAEymFHTwGlFfxbPP
/YfeScxYWbngzIEjG/Vp4in3S2elueWA517moMUqnl1o/UjCD3iCxOgentOFg6V3
5sB513WYf8L5ruvS4jannqhNY8Ebt9pqauslZ3f3nyYlyuzQLRekO40y0HAYIylN
iI6c7eJTnUpKcz7rmUZtubMdpVtQd48chZiL+Ms8d9z6UzPnmyt2tBJhpmegus5U
jbhfU/76XogwhnMiOw1fAZpdr456/IlI+KOK5j7WfoCTsynuIBfDn4ZtnYkExWfp
X/QAEZM8P0qNlU75Q7ZvWhUPPm5VBqeftf9zxkp5wTLjRhm1jxC02gBWs+LSr2xA
DOYo7BlQZCRfJhB/4tvnJOWwKgLCSkJOMTJCYw2j2cHPM9znuqYxcqecOGGI8WKB
faHsR4HZdWHjfMiWWmcbhQ0VaQSx0DZAsRCJ8G+nSfdNDaCJgc5AqaR3K9FP9KsL
41UpLKa/pKCHhUA7SNJUSTZDI/vf2hXc2nAplRFxUxZ8rAY5/7oo2cEcFu11bNaa
ZS/PjrJjnlRnNjrk+ChCYaHWaeijypZBJYPtZDG2pylzFnP5LxMUnqbRfoNHJP2i
zWdTmNxUxC8asKNDSFdtErVXx51SgF6uMhFTq+EfNJJlWAzZdseg8a9i0w+WrrmE
FbBfZxlgtvMC2jEF6zbRJdrY/DC1B705duzuKTfiqS/+xzEXdWUCphT5KYN67Zuh
ddz2oQ+kabAwys4KCqgbjt/Vy7o8hXFc8CymwK3Fz5g0+M1f76AXohJZDZ6mFpMm
XliTGUxw8lVWJzmB5JUZF/mT0hNM/OT4tS+PUgoryAfLIDshmtPgvjJVvG77Wn6B
dRYHClOOwiybn0cNX/0idVoFrlbp9JUXb4lFo1OZcUjx5e7Twq0EE8mTp8MgD5BH
4Ke0frjuowr2ZsHBZLuZHXJNYz5aOBYXYlW6Cj4odvAhrHQcz+WMQr6igqByD0uT
R0aJxX/d6na00PXLRwL0VmAIOOBkocohJKQbQj17gxUPY+VXuZVkTVv4bpURUeGe
8Sshk/wWEsyXDv2LbrlgXbkJIFE8Hiojn63vdZ5u8b1qcJBEO3QeuPyVHTRaDeyM
ECZqIWek4nJPNc7SWC1MpEy/DQxVTycKInQC8eDBefId8Bs/BVHxMlwtC5pSkzgT
HMl5e6udyulFCmPW5vLhzQgFzQA/WYUkwbm8U/nEm+wqQrgU2kUdXuxk3NCH5yMN
sejghtc8WZHmH4DJKEsS4cfDZxJwMefMXhN/UMMZjC1fqKHqzeoPEwNBCXNSNazm
qKUkQBdMgvrZKo1M5kKMrvvP3m+VIE5unrsMh94dBWed2Y6dAp7Z9U/KlPfeEJHh
YGOK/YiIeNp6QkQDQiW+332rq6CgCa5s8jNoJi6gvhJxqISGm+eUnSNr/taCB3gw
LHrMkOkLwEMReaVD8uMAVHA6rEQZER5CKHQ8ofb42YTI7P76CXXa6rAjpSzLr2e/
e2cyouRF98jq65uP/Y/GPWOJXIyqeDCc8Ayfy8QSW75EK2aZFA0SPyG5OCEnmEg1
`pragma protect end_protected
