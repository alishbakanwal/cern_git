// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:02:11 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
U22RcnOHEzwtjdDVkqfhdMZuCssEUFWmqHG0l5jtQ+Qze2B5HlK+WdIhEnq5BVFo
tGnqBzGlouvQpbYtsj3LWz+YeddSwwsJ0bfqwaohIeDEtQxaDMUoSJX/4nKHFUnm
AzbJ21B2L+hht+1s8qrMAMMW71KmQ+/qGxe9MJY6EBE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7712)
2V533222YDfAP0EXNeg7W6F9I0nIc/WYRW5a1XFjxEArW/HgGsNt1Iw2aXyrLrM8
h5AmCHuU2zljsXn3ycnoBAfUOFREtgNduAzr/72HQSGsmXSClPWFbx3/6naUJjas
/sGRP8ztWHZp5ZRCmYrpg20PFyU7JJ1JUgxUVJXzivySutKjHJtyJ6ZjCTcrXXR6
r6sgEdPuPwHHVahDC5Q8m/CX7U/HnQZqedFRaieVugJEMIgOjWsHzgLjvbb7H1u9
O6tTiROVTGe995yxaQ+jv+iSaw1BggnciN6aKJwx0k+d8iNISIuNc1U+tJFV33zF
AQnx1JTOceTU/y01ev11Gg2t5YMgtdsz+oKvA9wLHqi4YhrM08z1qvh6O36ulWdW
unQZp1MLqX+55gGbH+Pw/hFszBu3sidk4yy/xv6/s9MdxhXAsJaTxQpgwdkz5trl
PkZgawEiyX2XY4CpRyYRnYsJZ6Ayf7neGgiUjlM8Y6Z7SbGzvQbYXlyR3A21Wecj
X42gMiOZ/XPdoskEA65wuXGxg+Rp+13g5DtiuTit7LNpuEun7Wwgv/8MlVSIlKtR
rAIwkQqklJ3jPQ3v85MlPzYU3GSKG7udcEfsSQ9w3YENvjJZ9TbtS51S8Rh4HUl/
x0jsilobfCgOwhj8m0NT+l5tbOjtRlTlN44fijZuEdh52/ASB7HEWTyAvIAl3YNY
susT8/cYoHDroKPmjtZS2hx3P1J68LziDHwrJKbEfOqB72SEqyJzt9Tkgx9b9dRx
S1d8yjaQWMnu9OdiHL7whvKGee5V/JBI+NFAkX5BuMeW2HP+nVZjn3+W+7Kj1hj2
KpBXVHRK9FxamNgDxAZiZmRZT6/QFxVXlA6Y1jDfyuzCA+EQ54+yZSh39r3zCyGn
lEF+76b8zq0eWtNjjjKPE99GWT4Sr0SaTfCJKXNdb2VKLMzYHii1bLEPxGYN2aDp
+BweCY6vZS5DPR9kirKbaaoNKNqLV+qI+77f8uLzDr6zszVDzuo0Fh9otPZ99xXC
jWeohFS26aJgwk0GMTuN/oyWLEISChGpVuwEfEeyGKBnFDl+8fis+Zq4DWMnTEZe
Oavoy1z5rwARvkSGLCewp+WohSotXYmrA3UGFMvlynMmZqQeLC1M1ldCdHQjbnq2
j+eqQrunVs5AUfOOmhFhbGhgVa6Xq0RG0w+g2WNR3pI+NOwbfyXBfKp7ot710vSa
XIqcAj/Dn+GIK8Xwg6exf+GBUwP6wNIX44ww68ZerivxD+33GaIRxrGmCapsHG+9
F3nI+qrFGZuyuZcgl0ZZixG5lXvkiKGFRP9F9JJQSHmz+1FjF16q4U0hqcSaB1Cp
0cCkYTWij42eTVBR05VHkBZi1ujPv+TYC93ZPW8wKT5kxLm8qfbZYzRbou44UI0W
Wz1d7J7GegFFPnn9P6aroN5oMpMXF7oNn2roB0ur1sKH6FerGv20Y7BZTBN+YD2j
+VwVbT+4DMQA7t6LsPox253WZDilt3OeEH0yK8Mw1lHdolsqLpaPZgmAl0LATh6p
8RKfbs4F5ux8bsKdjNkckAY0BezPybVuEozkq8yINRe2bfuLoUQzgpNC4qimPl0+
ClewBgTPWJYm6SKQigUSO43WXS/ZhRlrEx+sPeAYd4NGqRk1GL9ne0THSavxdGTS
KnynAI4mdSLr8y1i08nvO/BPLiKGKS9jOfX/1x+Da3eoWzxzDWsZ/dkAh6ghwMWa
MtGn4wmFKqGvlmGM2RrOrB1bteinE3Gyy/xmocokA5Wa0lcQgUCyRPqXeZk3JpIL
2HxLHxjyAqVEYcjzF50dmalJ8YcAkaN7jiuOMwf6QiACBIue9rOj9PvoK2OIbrJJ
rpnm1MxR7kH9kadSe72zjeLkK91bN8xXzrofjWFstFj3gAzchWjsptEIvypbhEDv
D4UNsidgOmxaDWEJrVXdM0YrkfpNnh9Q/QIZ9lYx7uhjqEj40V+h0foUVHupqtvy
+h7lKFrgWCtZBuB8FbZCRXAhDs3WRK32pSV6/xVIiiVBwFPZCO8G/bSMweulLsSP
BwPqg4nQlHAmPGUIlWdKh2m5modbV23AmFGGOcWZFHHxUGoWMbYISDq0JFHR3HOF
GXrd3QiClrr0880LwFKSArrZu34q58kyAe/ApklvvK2Bnjiy6u48cnjrDIPlx3sf
8nn3+QlqrTehvDkjOTe8OR7/Y5O0XUwkU1e+PIxE+BVc13x+jcBV2phUxFT9p8u4
TPSGrzFhZn1q6nJTnXaKd0sZaoosRfC7XesuSTLlcBIJxwIGkholDNXVWXWz2xFc
ZehwlJ38JoLYgC1oeYhhLsVn1JVlZatEVrvtuUVGdJWAFZ+CgTdjLxbGpJ/tCBnk
0iI6U9uGaHCJaMPo/zlPG2ixrjS81934lTRE1Qg3TPEtHEXYUd8kk9jGctnNNZ48
rjAhCE6QJHrc8uCWSURHsNmvd+sDLBW1KHDMtKJKusbxYD243WA76T9tiKxUx0OY
opQ+40wjW+NxurypHtJpM1Ei5u4r8rTVin9DegryJYybiyQU25VSvcgIc4ezj7b1
LT9Tibm0CDqWVDRBHpSrR+PggYZL5O/6NnD9cPtLIEAdgn1u2YaMXNfO2Q6QpRQ5
8nK+0p598H/WBMRb+0cFVJYn2DeTvl6bb1tsKyRdLyJKCH5H6JAfO2bHGpa5aVs9
OJs9wIZWZmvEKfJVnL4mxki47FlF6T2KK4kCk/qKlQbnumRX5VeTQ0CfMgBLbU0E
FVZlIeXWqcmd7WTd3mRWZM63e/vTEXC+jbA7+JD2JXF+FWD+J9AnEatu2wlUI0mD
nB7M95wasg2LaXrEdfa+HTXqRAb3EAiq4o7QFQJYyVdbg+Biwzy2ti9kz0lt//Di
7ld8Qf+yEgYUgiQRWxu+95aQvUxS+2WqXEUNKGBkJl4mORgIy/b+ubRxJ3UfrYEQ
w0kuVlR+2xkpnng6XVNeR7Oh2EBFSErPi2mmInbkzXAPXvO1LfkcAiOe7mIi7KuJ
Pr3FQzcG0U7UqJ6q12jempDNU5+OoH3OOrD/htH5XZfHgiJa64TyofcFzRY46/JA
WsHw2IylxLe6kLZf40HVfJKOsWofDJyFQA4KkbCjHpu75MjweT7fM3hKaVq5TTYH
wOyHKBlgEouRn6R2mP5m8W98O7J/Z7iXZpCYL52alt3dxGCDxpD60mUjZuHS0j8R
QyVeZAP2EOhrpWzawBMmFXcmN+T25TXZ0Yel55b/HblMSaLX3aGU3aptvx54DwT2
AQqK7BJSbys8ExO3eE7wg0/12+5ej+qmSViLKBhjg/q2PROOMjKjf6l8d19UxczK
DkAVj66IndmhE9dTb6hexkeOBDuDaeTgfNo+jRpjU796VKAorB5j2JJgQ4NEjwbi
5uRcNn+RSV4uHNgVqt0bH4TUBr6fr/p6QuEJW+IL4MeNxLJNvZr2lWNZui+EoIyS
ZjGC8MepXCxcRSsap2+ykMGomtIK+WHLrsK1hRKtLcuX8NzSnQ8Cr3qhNnV1x1Qh
FSClmi+iGUvdClHo/H5Ou2F0FuCCttHAsyZAeF0aUyS1n5sbBF6JuIBFUQr6Q1Qr
0ykiIByd/5pD2ZOGc9siG7jsFscNLuTOZftWyaZTjfgyayjiyfHhgsg8kdCAe8Si
RnwsKeBIZ7slNT+jR+h+LT/u7C4z9UoMWQa/AmPw+xcJ10ysrOEUxzv64EkSgm4d
aBgiStM123UO/haxfuKamJOTDP+ecl2jNxE+3IrwOj5BVQj7BphFV2i6infaF+5h
UHE08OUv/XDS0mviiVtQd2wp1cNz27u1BXerNJKXRtkvmwJ9k6uFP5dWq+fVCIZP
z5GLY3S1fRO5dJ6UtngkF6E8X9M26TvtCANQEtgye1Jp92hZfALFCd3z8Dh2fDUn
NiEhGv5e7WY4yUynOJUg2M8ltx7yIrb4CA18aotgYMdSLdys59u6hLTCxv4vhYXW
LKtdDNrbLBvlwILD2H84xhnQRy7SWzsOGhjRp1I+enHI9J9Dj8Zs/bU71tY/WAE5
FoIeZ132TsasywzrOVD/m2pL3o0KPDhNglQX5GJWVIZZjYrx5SI0hGRCzR4dkv/1
mftoFp3hoTbojy1k/ffv5qrxsm3URpK0cGiLUeBx3GQaxoXpf4sxjZIblW9KRzc7
ST7WcJYf/XVTSsClmEE3tgCJ75sl2JQepOFAU93ntyfSnBxNevZiRXDQUnFvnOv4
kHudUI/0v8XfpROArEI0muI2+uZICqzR6Y9WmFOSZn4FKvJCEJ/XzicKfnH/b8sv
TVNbpuHQLqLSJ0v44Qhl8I6feiko0g7y10a1iOSr7Ycm15uEk5RJIyhAa64ORpF3
o8/IsPWmkw0aJrd2ctmKG2JK5oJYJtT8MyQzgxB2FKpDyUOeTk8HNG4sV3uVFhX8
8TkqlW4BF+JGeetzLsDGnjMyCVHha7mh6UsPu0t2pIMXrk/FVUur2ZQE5Oi6+DYx
dBZlq6M5pzeyN9J22LZrB/wD7PX0kHDKnc0Z/eoezWybmutC65vqztCeKC1u43yw
x8dQ0elIYa0vMpJ5qLBVH/VXkslOON8pJ7hS8oeemUgr5jGkNsOdadTm0d6VFoAA
xpovTQGOXBP4qHpKkskGQZFyxkbcQKp8wpTz8RTOpbBkYZo9vf8oX0m6fve9E3Y1
NRYB22gPtw9Yq0cQ6FrwVYgb7dsl/Iok7r1XpFXX/DbfGNj5K3hNauRaZ3yGVVd4
wFH5qa3m8l4l+6l1WEj4YGm/TQ7NvQr16sxz9KUcJ14RDepcHA7Ska7i6NIMqC5u
5eMqcq0i9yqKC2J7UzaejImy0yBVVQa30+fkqt1+0ZQuBptfnW0Sz7+mCd7Um4pw
8h1o4RQzVQRlzJVNaTlz5eS0vwlqZyKS4V7caCsVe7s/De9Dzy5m9qkvfd/JuP0W
zpU54cOQ3lUlxXVUblFq2g330+9pO7oIHUoxHdyOrFy/SJNDMiaPudUb9Eepa/EM
IN9RyZ5Da8UoqpHz7Re0XLJQ9wOiQeqcQdKpnnox5cvQmPJ6ECXzpX4SemPJM8Dg
rfXzYPg3FDrwooMfRc9stDmmw7TQSlF+15HPboPOHtd8ZEabQYO14HYiVeXRMVA/
sO/iqM7W8oT7T+urj8k/GwlDJpZIDTh9DwtWQXuZVMbQ6FjT9oZ45LIo9JxkqqA6
2I2T+3FetEgTNBONr1MbAOG8ZiaKUTuXV2JGa23eClnC1dN0kjx1zY1rT+qhZtGF
L82JfWQVL25IepCxkmt6/tpUf+JQxvuf7utLTWNJCE6YT90trYORbjuzsGTu4gE4
VwU7rGwoOQtBSdk74TCJbXAYNIR2eAwRYJE2d+ATvNsQe0a/Kvp07QOi/n5fGY0A
QM0ZR5MEiFTK2ut+AB2v1J64X66x4HU39tELGL17n7VYq4RtftGVlmbyRvZafaLg
kVYAKvu+NQUmBcJBzkyZbYHKwYW1U/FxV2I5fGSomC+EiRLECtoGsALrBSnJIFQN
ElE868pdAnMJbsTTAZFkKc6KP1jcpuMZf9Yl4ScDdsNgTwfdzGdtl/6U0I6wXGXc
ABjZ/8DI1RG2VXyl7xT+IcXW8JAbMxfR7GZ7SBmUImyhYsRXFxmRw5fLWt8lo3k2
XG7zr7AhMlR27z2fpkFxgdND77wJYDAIKsB5XytBnH/WCCecrm6xKc7SgdSRDcii
TLEs6/3EJ2TYwfmfKgoqA5533zE78IMyCGz6If7a6Or+xpaQ5TX/syYG2cMpHqFn
D5hYj+Ka4Zcb3D3twzl+XczauwWfUoTUKU4jzU4ivmMe6x3nPX6f87On4CtCue7p
UDL+DIeLKGzNnSDsv+mSnGukuYhPUsEJ2vcCYBXOJf/upwQ9w8zk0yg2IJoGWNgz
5iTpfBDsx7Xhv/523IfSrLmB48Gezm5hvjz7SCZRzB91x9zO9zuXMGdydPZtb+Rr
yGE6tyuL9buM2849+elmO9GQveMKteCmLwTN+xeEt73HwUNgmdDLSiuI2mm3ZnWZ
S9pFsC0Sam9Dao+i0S/xa9uAXQbHfTvc2h3xUFyQvDGBlq2svNEz6USK5iPZaf9E
dxFQ86NMWvdUPJ91cLwR/f8QG7qIIMGsCMgPwLX5pDSKdNRm3dWLlD9OZOjnhmwL
YGmFNk2bLbNGUFvhMMDD3mux4/uwa3lF83tb8iQNR/HnAQGtz5FEHHCr69UjQWXA
kzgA0eFcEgo7eznrCYk+KfzwwflH2bMhJH2dNXc8X1UH9/e89WGaflmU5fiXpipe
GklDaj82cOoGX6Z30r8ghmHf0fRqcl+Wl19DxLDZ+eG1+05vm7rFZi5YvQZ7fVrA
6GkJ6cK4NO76waiqWAYHQMPyjtFoYQHTJH9dOqh/hBwjOX1ISbBGQZG7Da01eulv
Fq1wNJyPNcCCdrF7ebh78pTWnWpJVpSjoTAlWDVQKJ8d1F7XGtbUS4U5TW4RqiGN
keLwWJCC2m4LnicKWXoEIXaGi/gV2L6ZaM2LZVPIttMgFMEZcecaxJBgDdV2f+yj
EILPcxpMVpyZSStToUbLoYx2pKYV0zIw9BzRzrldTm9HnYaT//1a1RN9jI350X0O
pCfPV+9lMLTicZeG5amMNyt3Xak2EAHNGHbjL8dna8QMe/BX+VqGPnv93Zvnl028
hdbDNWECdJ8A/A//K+4JZEI2g9cIG94fDKZddU4DghOyU13krMCy/ziPhdslRU/D
cwMXCAqz7UPKEJeuhhIkVYMzYayA4N3jQnhhF6FbPFt0ORFeyuU8nA3xrYh7VYiV
XIf46QBz+Svi/SP4Z7zrD0agGTwTs6AmK2x/2VG6QHJ9Isj8f3q+Y6+EsI/HgqQw
nXxHDF5kwqyxO01EimGDY3l/zD36TwJuVbic+O2Xku+7T2w0uTgwEgd2udxSeUrZ
0UF7cOCTr7ArozBcqmmf61TpMmoiYbi5b3emx1nqjm9pmQ4iLUsF+yTfLGQ4eswE
Op1CqehqjVIuIKwWo2Q2TrSVK4aOjJ+f4W0UMu8gebXzi5CZ3rGL6dFZvNRVeo96
kYtcW8fdeRATm0kl3FK9qgZgyc8iW0PELXx+tHgmfVWqRll6q2ZduNsxX0dPWdVl
z0dTyFuqg3kUtWp/Y+h8hDr9khWVkfTZnlNI7+YqnGlojOuTWHoQe8BVZjXSBl6S
nJmEcA9ndct5XFdYA5A0ka1ig/Ew5ikA0mLk9XFOJiv6gUw5WtI+5Y5EYSxLYQoZ
rzS0UEorPTFpqELODdPU2QRw7tHc99wWEu6YKoITn3CATTboFB58eYuwSqBI0bSr
iCE5g8QePEvgjbdE/9DYSPujZ7MOdVkUD5VR5m5onfUBZQeKSK5EKF6izB1zupZA
c9P9FbZr5mhQhn/1N+W6TZiOxNStY8TiQ+CtYi7bpddQcEQCwZJI4yaAUx45n+ia
7mn9CWekQTNXElK/pkT6iiYLNyNBkpZuP4/a7h1MXvf4vz6Tz9wTlDZV2LX6DYT9
ryJC73lsWARWaPJpTqsZkN6JrJEOf4RcUoCvZj6f0nzMdvtakCMoletjBytsFk6V
FFXXExarqISktsZXyOST4Y6NrU1cjpECfQ1v/pFloRN5Mu7WsAarisSYjdal/0s8
y0lnsxzWcekWh2OUqiedxgNcBeuMot+hpn84anMVjKNVyCBgIUFCr24B/GghuZMh
tmAk9RQ8XqbdWujQfB4dxGDl0dzVCJ4lMUmxFOFAbpgBy72cxurpLTI4AQQaTTe1
+VGTuK9HVTMRZlxcPjo9BT1LDgA+sfcun94U9OzCVrBdf+TEbnWTnWqKgQW8ydFh
9ffekMUC1RinozQ7gweVM6liZY7gcWHB2jJB7YcE2bMRolIzdwurGwjJc9+hCqQA
8t0155NXS2bYcCWBX70GLHFc0IHkBrZFYIeJB3iO9xkd++GvTts7cWiw7fX8MNvF
K4wTitySR+D6vEXSUiTGfpwmDJMcLT2k/mg3sKHEFOZTE3Fji4yGxB8mMjwRu7qX
rQ3UlBcFa7YJEg2/aMe2oTULMmFS+MgBVl9W+iRhwxkM/NIFZwvlt/kPa7IJMrec
PdgzqQ/cdVJz5+6NqRcLQ/Tw9h8xOXFl8c/byGNl3PqpsGbsAFB/k90UjXm46Xxm
eM97oh57P/MiH69VM3ofgv9zK9eyiR80RdmzR2vj0l/sqPU1SfM38Q/ywo6L/Yd3
2stZ/xXgr/pydknTmip17Ya3XzUopRT4D4+qeIEayTyC1j4ydCzbWj87Z0ExjypA
ABZy4RlZPcSJ+LptKon5vuTuXmu8D72d3i711d8AcHk2nV66tozssnkWDngOLTq7
yhHA3KKDFg0agIAS40rXdpKtGw1mO3vyo5LlT1J6mOTmrFuqrCUrYVpFQEkiOxl6
Qb14ZJzZtocdC9VhIh6EKctAZpu5rmCaH1BjpXZPCd1SKQkWR+Bmh23crmdroaSk
bqC3KjnYwNBzOYIfBjaLdB2+Q/A9Le5BWp0tR9aVefAu0wnrWYBUPffK7L4Y4v/f
A+TtMqSZRuUgTCvGB90kKkOfYDx+UizirmQJJnLVhbR6J99sT/G8R96Ay3fq5gVE
us3d4i+lbMKgUV+xuNGbGX3rl3K2H0ia4WqaLEcxlZzGvWto+hto7zDtwNml2t8f
l7aXvhhbgcTYKnsBmp2go4PBaY1/DCg5XvJAnBGdDDSeYVO+awwyTNg+ffifJanl
nqYm2fY/4VCsecxguv08zCMJRTwwP0AkcXq8rqB6WGhpW0ROTrGXYt9XAuFOTMQn
WsxyjI46kAWhdlGVLlsDNnf2+iNViSKFhj5AGTrzV23Sm/of10Wllf92Hz3Dq7Fu
aR50iXqc71l2M9k3psmqZTE5+0SBdVrLj6tLypRU5VKvo0WRvvsRsv5h0sfiawDk
QUVP56S/HuPncfG1NNZc9eRA4lt3uMPgSPrDuNLpGLJLqSY0d9TiFHrDbUWb3TnD
xH+CSeos0IQBnodgPoD8sgW0mvD724S93yEOK3PcmsVqa4vFreZuARG7hJzD1pd8
hjs4HKC3gwAw6pxyMBX3zXHLxSgRqBRC73Pcd5Z9VGVpKYu8bIEXWYphQNW3h0vn
FaRUWw0k/2HtOcp8i3j2qBN3tJyA58CQz1mUU6PTK/NG5CfVieltgXz+4ZZoEQXi
K7um7dzuxhTTlnpwtDR1MJXIK+JE0xtz1HXFfLVfFAmOt02YJfyidLB6kdCOGsP/
Ih0ByBuJV/McbUne2M70eau+K33zKgrO4pjlmuJ0tV6/x4jodZ40vdUhpu2WHRkc
FGSd9CkeqGvUpQQeB1L2IxiotFbg8rZ9moUYTiLfMi/AFmb6kV+qCh4xEoBvxjKS
LZba9fQxSjQKq2JQQgB3QoBUKB8lSt8uwrSPhK4Ufi7K6ip+UPxsUj1G2p4VQ/62
iq2iRXhfmXgbKeDnm4MirySZN9rFV5HjLgQHrPa+J3kPRtlNKJkNsdWv9XnLlAkn
zWcU4Nx2Uq8k0PTi8peLfLH9bYNRf+NSfoNotHNwDW1WUThnWBnL6TB9kgRHt1zH
j8goC3UasSq+DM+GU+dDVlpLMfUElCLYC2cSbyBMP6VHsE9KPPU7V/ofA6swWlP9
qOPRzSBMjPE6wgeHIGz92No/I5QpJXnygU4PyC/s1h52vFEasw4D6icI7IyURdOn
NtRTrIIqaAF8kp/2NO7VzDAZFB+hlR/i+RbI3oKtWINR9m0hWnj38AmXDny9PTZq
70EPm01qu3n8LKo4Msnf2wTXQ9YwGJBbehVYKA1H4CS1RHPzVXcuqv5gIcGI/oXy
rAHVfRoAJb97M5HOPiBHtWKP7KpNZMJrzth9CilDRy/QQUBCIW+gv5gjJccX91b7
/B687JUI3JwqxcObsIAxdJ/dPfhGMuauQ74WcvIsRMi+c4K02Zn2CI11vRv91sKA
PPpvqpSuW3EltnNeAdY5BKSP7dU7AgDxSSDxOayJkSlrV2WUtZ89iuFMkvrP1TRh
K/PkPgPtHaI8R+ZqbY9CAGSfZhGD1MgJzHvAq9fcBNReteSRsNeLR2SoDsLUbuLD
K+USCNKpT5Y6eJoPNc575MyvqVPyxnReCB2Uo/4Z+OilHBBDzRiWbJ9aeSNM9L3E
aKm7Tt5wVo2VTUEHAVYPFPuc4F7jWNoA19gmLVCNwBou/CwfDhauUQfYTGO7OFbC
4tczBZl/gx8vRN4o83C60lYPcll3etn4zQR0BgY85CZuwINXFcT3FS6YJ71UuL+w
oQc3f3/khe7UIMlznvwLNj55l4lPl7KaIi7O9xiJTVw=
`pragma protect end_protected
