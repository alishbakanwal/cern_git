// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:02:08 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
tNWA+ijlDKEGPKVYl5DKQUI3UBD9WZ73UpaJqmmYDCNduy5Vtc9g/EyUYDKH1Hlk
ePV6crWQh5RvgztO/RASW8yZGrYSETK342kdk6zNEJbmHb7leXRdKe2BszYZ0C8l
23WDZZUMjVOicrP/OpS/TUz/VWEVHs/2ckMsbGq2EoE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 35392)
vDuRctJbuxTsWkqWZRf8mND9TbBYF7yA3RHplAHsY1+AIi0j5dC9YhPh10dOtYlU
jT5K6tm6d/VxjNG7tXQOuKpiOGqHibkgeL9C5zTxPf26jik0fk+XJHlvJ4K0NKeP
wKLEvfmJbZkFZqrPd5amLJ+mhisbcHlN8A89UTCSE2dR+VzovtLnlTxDNneL0bqP
9u/N4SdXStpZzDZJYO6WfBB/wVUmhcNMac+2SI6bVC7tBm31/+L7/DEKWT78gX7d
dkAtJm+i9UNpVmIL2exTO5SnNujnsrnj8XRsSAjRh3Lb9giCRANbTkz/1JUQ8Me0
iXOmKHPso6lo7sWdrJ3yAN27d6xDlkwxYBMAQNwio5KcmCYW8PPE2ODTzRAKvcFo
FkSKn5GePwKcn/23MkFiWgryptKrBj5wfLzSossB/J3KF21pk0ska56KoLF+J7zk
NOqE46/C66WiLCw59zTNAP2etr+UYAscwaUa3rsWC5vuh1xr2cnNJ+KBjOak3cQE
V+Rh5Hrr2RJimv4xwuPUlOY5zv5qhBVoUL5HJ/ibSX/rynG1GOo7+QIMRMB2BffT
N1xVUbO2LOkQMf+rcRLry/KedVnsuYjvUn3UuAEe4jmOfb6PbIdt9IGtKFEeEfqT
u0XRVzvXXd7igAeridAiCi6m5vAPaVTN8ihrNyhRMYDKd343yf9Y2aRPLIrzRypD
ByuEt6eBhgYCANo0LaJybqnP3tfTL7t8ptQ/Bpb9e53G1+QkHPnyW9wFQmfAzB4m
5eaNgBRECUWKCt7kqdo0pDnV5i9swpl0ly5pXIHze8DqzTCAiqO70Qx+Z5jVjKD+
brVLEVyw8nYMIk+gaNJBozMQqnlsZVSfuk1mFDei87GdVIWyRiDjzOBBAUl18iyY
mcy4Gyep7e+MeJaqGAc0vonRZm6e434glDqrwwQhNKk36ls3ZQ29FBQYJd11fXNO
OPd+Q1enjwHWJAH6iK0rqXBVouRh1/P+6JAl7JqCtqPFja7mVOBNUfRlRQIojkEc
K2JnM+XaZz/10XLEBzzMvxIi67lDQwm2Xc6HveJdk7bji+BTufgs5o12BC3/e4qw
fOLGiPx3lsWkf6y36rriNnMP88s2kf8J8Tw97oEzbd4vbiq1eAeMg1Ydnekv2Lkf
Jsm6SnX1RPdm50MM9VYaedMtEdWR37Hklya2SX/JU37AkqdhlltoCRD61my/a7ko
M+Ctsb5NT8+T8xgiv/9k9wZqEsR8PznGrvjvEiuH1GbzItKx/VmFPDNXrzCUtV3V
m4N883JSKFJbeAOiwPCHLRxoHN63W46HlEUZRaadDHqDnQHvol1AGtPBK0E/FKvT
HI+MqCU0lAya/RXHsByMEyleR3UrhKqW2RHhVZluJd/Und4S3G6pkBvMDzG7cyJE
thNzL7L9Wf3nWPbKXJKlycGNnT8mUj3nWUy/5a0WUUzX3LYlD2PoROzhaqiVPZ31
o5Z2/LREKQen5s2uoKbcz4POZYVQYCKcCgUHBwGswHuvf2ug97AYr7sjqLrQb5Hw
e/xw95xjFfoCG1bPSXdWOAA4bKwDRkEXWK6efpn+Tycyd1Sf97IXVY2rleNIRBEp
t/1H4q/QDZo2TA6bdEUQD5HpIckrvEFnGTV9iB50bqvzGKHgE5srtaDPDJY3B//W
SfbhIDY6Kx2kJMi836e2DRQs9l571LTw9n9LjYtkiAx8caHw5teCaH+EdiToInM/
bplZpedL5z5IYGOpiHAwdFZxO8a8NfaNqU7Bz9vGP3QjJi03RH70zIGbjLDU8vQP
kgGr+eTki++PinbLEmiO4Jr7IjNQMdtw4hNe/CDboNCG7PrI3PsRBjezZrOqnLTC
q5cWxro06K4Z8hRtfYUrktlM8wew1oJxSJqxUmebFCwY4PNddj/2599nBQ9w9wzJ
xPauQy2PkKUpyn4+UlnEtjXenRVvgbmMiB4bFTUCBePNSbQUPsrIMP2aF4nDkPnI
8IIK8ARG7jASDaseUHzE7UCoJh/sUfN7c1k2c3CH1SFAswFT97cXd/KuR8YCdrkB
yNaN4wbN5KxEp6XIYJ2tLVGGPHVfvcm+VJyoYNUT4mqmOhRcXzAzUj9XZql+2EPr
mBsGcdgh5VT1HVTS3EuD9hcGXLIqXC58NgT+ZqlxeFzc2mMOpEUsncr8wPzoJ0nk
MnDDfTCd4zcomH5/NoXoabzEunCT/OAHP2x0mW1QiFL9Zizv8SlnN41bMrVTCIaC
bfUb2dDl9ZAKNAbEd7SkVmVu/zGIu07gNYVFgED7elIuQSp2HYxLpK/0MMsL2V7P
HNYHuHxrAWt7xmXP/drvx22IMzw6ClCzqkiaubdfx2evl+Ostq7x1LEJZNJnmkjZ
3gkwNE0zRYtyX3DH5SUhm8nUDpYgVw2RISPg29ub+hmhuYyqEZShFc0GgZqQ5AVS
fgegkqiAzKX318wJ+iOndGEJP1NY7CT2pz4WNJdID0RVijgbbuV7OdSqEu90HhE/
RiWZqycXy3ZY8rTW/40xcYIWA+lb5IQvMO4pkvohY4HvtmZplGr2FaOuYVDfWhPh
WmT0wxm7Iq67mE1OK9VHIahUsBaOO2i3JgNurFzP0cW0VK1E2Rwjv7ES/99b6vx6
lp05t2Y2jKg7rdQfdWd3x1L0KSs1yLcEW1eKt8HAFIYJNub8hLomqbsZERb8e/um
C5fDei6q7y7zYgeE/TPrfawU/oApDFfmDwgtn46P/xxejLdRAERAxA/U2kFjaYD/
hVxn0wsql2qgYv3KiFn+w7GjAbx3BexmoVEvswNFHgPo3SB37DYOOdhAcJWPLB5k
b0MA3M5JdwlGy07FY+U5/lDNIW7IgedNQF4dQntRYNLowfRHebGqLAm68F5ADEeB
y40S3RSSfSiiCqCRgpO7EW5rBH/FPQnMtKCMJFHhtGJQWuR5vJbhNUL4QIm8BlOH
i0MetZduP+LXHy5Ll2GCr3Nqym+n735UAfGoi14U1JFXXloibvJnk2/KD6qV1xFR
J1SAKYOabIkSfCow62uyi12y93eNW0/mpDb5sluL32hznkq2VSy4AOUy/zZ/Hk5y
PJWO2A9tc6Y3pEAlFYlmeLT0+7djYRVQvS4ytxtRDDq0zSSSgRJ/YVyK/zA+2k8I
f68ZyyTgUsMRKO/rcuF/oiUsNYzI+QQjbVUZCUaxqOnycvxmSLx7VdCl5eDqHCjI
KsH65RgpuskuyhvM4h3hiT1tW+RCyLMeF37lZ510b7SnumrHLI0UjxiEqLMLfYr0
bl5DAskDd64mitvBAbnhCypt7Wrl4m43iWvHmOwrX/TkEf0wMVXmral63NGnm9nt
voI9h+MccVnDRXtlAUt+iR1+u89Gzl9ouD7mEjth+WsQYP8qnVSFcf1tNf7wW+rl
bvoFGrvWfi1piBhXlY5RArpItGN8PSQcAxIdlWKSOt+FpRofXpmSI23GFSBXhr2l
aRTH+Y6eDBXt1Ie06SAQEMJF+l8D4Q+41N2PJe95jBuOtih0MgQ+d5GhcditxTwI
qHkg/rWxYJWmavEVIqVn9ewdgtaRQnl6aR7qliVXg3FbqRz1SK8yIGaGqfF5DyqB
cDnKr8NeTO7zAJyAmLBOfYzS3rBBLs2nOYjJSWOXkjktAGMemrVyqhGpjuycrn7s
gxgx+zYDYw9/U5sidZzYAUIF8JpxFx6jNRAVAJkUCE5TmkZkNwzLub3/ePhgz3/8
39OSX/rk8gW/COeN5H7pYtaz/X6g9MeSycgArOpSmtLCBH+6vyWjo9HWryuu3B9K
dCqkxDR2n7dtMtXrEiPE5NfOVEcVlwY0H6cYBRimvEA5sBKSASGlJ+smun9Qr+Sg
AAawHXjJiCAMjegR4N/yBb8PvuGpg1uHlA1j2TWwy/9HMWLCLI5BbmWWhLmynXWK
U+pvsCIDmLRQmkh4ZySQwX9BoM31mMoZ9/iD4hygAo1K+WqvwW91N0O08Z7Tf2qj
d6E7M2NMIlCFdOz7TQGuHrxEtVa7mWbgZltjMOHTg6TYgFe3QwUHsCFEYZIeQWk1
cBr4q4KbvdAa/8WTyYcjJnPiSwCObHa/KAsF39hC8bGa5NNyUIUuGvClwGW9sBp2
fx/q/64ZDfREjFo74O/FXh0cGEC708PyDIIRFSOPtnzlcwNwFnOg6IfI9tdQydwT
Mt73seuh45rEBQ0iXhPUP5zYaRz1jud2PYcmChVoQitTQWWV/6poJSyFqHHbb89P
qwBcHzw4yjfm+F71q6pQZbwp2MfJlfeijfhataVQ9/BwnQQJeG3/Om/QFXNSXc6C
p+4volrQFGKYXXm3spCehcc+HTa1/SUO8pIvxMoMwHIq+Gf7sI5RSNjVmv/N8YHY
/iQbrFj/vUn2ogixX9a69yeEdk+Di8mV1mCEJp8tvjmGQW5564NRin2qSj+8anuZ
S9m1eM9gWbq7MUPxr71w3pNqn3X2s0G2pL4gKOGgDd5eCzQhYkXYsHmDL+P63vGy
n4MfhPO0YnFLAraNRlpe7THNjAWwK/lyslKos6TeYgTRCLl1ZYljpQqjI6M62/8k
qdtQfQXOxjTvds5jzNDLF8Y49wSkJ6eOIi+GvrJPOxPq8NZ6NsgckoKW0BNor6X0
px1DCzAB4AogIcsZwkDnzz/6tAnA/T2fH0Do4KBV97vl7x4IuieA5nl+G4yNn1NM
jya9uRyNQtxBQOUOKsjUTSEv30ZC5DwtqzDG597yqIlfWaeV+FniYDTc+suESVvm
J6U56+Wi5CNlkXKXy6l/gVsgKixvgAjhG7qRPm5riBh+XJ34lqPoQoAwXBRQau6c
gWwugj9/bXd6FiCxAjtzfwtZRcwzBPhbDNTlSVR35IhBy90n8wFivpad7ZBe6umD
kVa/1PBmTAn7GTQmATTg0ly0mQ41gIfGJ2Fk+nLQoLPSIN+bW0vbT/bFQ9AxzgDD
Dm2WaIpSuedOflzsBugac7p2xI3tWRLN47QXce43gN7HAIme1ePd08wT+VdoKZqT
3MSiBQfsvUNS7jSnnwZuUfa/MxcmVR2K+DWhrd1Hxet8yXTglaIkkenPFe92jtuz
fHQQS3JnGYhRrmz40R1EmEGi9+FlyFU3d9o6aNEO86h2x3PtQ9bcbgjItUta2kxq
TnQIIMLu/ARVYj1N9X7kR0g5WokH4dUt5nqqiL+iUVw80S5qxqUjSIi3EuGguMTY
bGPG8MYZeMZ0Rq6hjAzfTUErkGUXbk83FqCLZQ90IU5jY6PlD59IerVFdThi9w1U
G0EQz1Ke6NZhC+dXkHEypmNr1bttGQG51y3nnnTNdgwsfhvU5oEvHw7/UOkKN69i
Nd1gP7kfP+ExyTdCsz8FgvK4iLu37M1q6sfBEEHjtQ0Pw7XQVSsHMn0/P4GieDKN
4YFOZCnpr9Q56ZAYcBD1gxo+Wu+3ZB6FFh4JCBaOM9K1vIpDk2FB+yi3JA/UXRDY
zAiQrAPGnAz9Qr/2kV0JGwXYyMIu1HxFyXmYi43tNbGgIZZKZRg5CH6cmlKfpKH9
fb71Zgxn3mNJi8A9+uV/HKEWnE5YIw1DhLCLzNPplijnevZ916PdwA0D1Ml+1iNR
Ci/H31z2/YddOw4z1NoVimFuyWARZE8FsD478MBZVDT75/GmD/XITIR1RamCdImx
HhNYeMTFsjFA9FDYvxluMJJveK7lkT0dsyPLIWMJUKI8m76X07UJnK6xiZlENIqF
z3b9iGRquhXH+JCWtr0vdKTsYAk1VRRQ2+qmh9mkJlXwsA2Inv2vlbffkp3A3eRW
Uzp3WhoSIh1PXPabiliLaOn6L1NQxl3cwCNxysVPi3djwxcPBXjw4q2zz2BEUfhd
zVQ9EPCY3E1kvBMo0NrEoMsJk3skf4p7Xk1yZ2Z0tT6zD3pdCJXIau+CdWdBLWOI
kZW3telv+gVICc+GFykRpPhNJNVhwzGcOpZOF/RyxwJg1cay7Mqs5ZhNC8hVmzMw
5XsR645zQAC2TziET0qc62uiMptw90nLiSBW3OvumBOtp8bF4RxlV2rlBE9LfdWG
OgXartM65UCoKIwoWQc0hFlm5rg9gCaDencjYkijEdfF6vhRbqPb4yUtm8CsAwYi
EXZN9Tg5qMkKo+h3dk8dt7xc9kaXPQOEAmlpVF/EDOyFEKYiR9QMYRZJ5bLf3dP3
hh9k5lnxh0XDWzdBs+xSZg5MnXxBXApMVPRViGimVRjrjedjMeFoEROIk/FZmAZf
gXTvPNy73fZB3nlYMs4CuD67hKSw9R6pkv2ELhnFRcbk3NXJ+pCSgU5u5TJCZWB8
HIlP9LxEdEQHGrwg6e92YhzvJjpHqvEbG93SAAIHq12mdx4LgLDo7KdGtl/kvAPv
TsgK8vWEHClJvyADShnqZk41xDbiVbaV1LSP+YtXIiuSRlvsCsPFUjSE2uxq47yY
f9dGtxHXG/h7KHyFxkcKAzBQAyDa7mJgLNOMsPrmcvbeUmZiJ+pDd2QH/xFaHy+6
UjWa4NGdE5B+nj1ZaLBDhFvvHTIJhz9LGFLz1JGEcSITa5faFOHuJ6LzI0YSl7Pz
g/ZOqXXw15WRX8g2IRFnrYmEaZBJh/ezTjtdtzyOD7t9j3wjpfMnnw588uZo9E3H
9pNYZpURJyyYuYUPuiGg+sNKc4ZS9QaT0t1znfc1/TaRUIt5wLVLxyUPpRXHnxZ+
T1sRwCDF0gG5qxKXMPfMymvxiavfrs8f8ezQfY9iDOGkGNJ9yiXgcBxQQRF2OHFp
IoUz2okHK8+L4x+quXE+PKPskGJSUHEggd/RsaejqlbhUKEClGr+xN/qtQNywqAS
Cqe9HwoWuA6MS4Zytsn4TZxfO7BD+ll5pJodKg4PFYh/c9LpGJ6uHNxLIopRTJn0
veXk+VO8FeO+LytKGRXgk0pFwAoHbmbliJoWm70yALanfROnEV+7A6vrj9az34iW
2A9rmzO9malA6E1EWHHMQEZ06LIsO+hwCv2VZSwI27WmRVWuQVtUsiLBquTgiZfn
4UOTncXo1JEUKbrnTZ88dNVONkq9YYDcyDw39Fa5M2/Am9BG/V2J7eaIEuxVIBRs
xwWiDzfEUkFsJR63lAQHWl24JOuHmJyv/BeUbmNwo60Cw0WF7PAfYgJ4qEBa1OEe
YtptUEpq/xZR9U2jIfld20YjFYsUNqtGurwGUcmNncwN6oEOpLFvd/D+6wo5ArJq
hUg1fKrLeRpv0ZHIYU4zjppE80wd4wxq/qaoIvO5hFWSxMyfs039zy8sm+FhWk8a
N6cWat/zc8jYiPTIcIsC44TR7Xis+CbD0oQBbeUeQo5s8g2Tzm1IFVJkew4/j7FS
WPRbkLpKDrQjqCV2ARCijvL5cuZ+13qnQ7xPCxTyjrU5k19WcDftoKO1zuWtT4Rn
OuAKurPuS757EKOsbAhMSU3rQHRVY6ZfNjzGJlf5hSWx7enjQrFwIGHC1sRcDR3a
AyYRgQ6SLJhsZeqGSb6DLczwbVFS6uJJ+khiJFNk4CiJE4EJOZf+XpUYK6c7oDGx
at31O4tado3KTwlQ52X5rPFWJuhzdbzEHTdXhiZW1gfV5/60xIm4UCf7dcqHwewK
KXdZSV4GxGBZXZgwahjyHz8+5seCGsz+XZR3CMsZFdv5MnIxgGo7A0bFUMe3g61W
XyqSkRkTdQaSh+VmPXzBSj320Ppk7RNF5VVtumyU44/1OErKGYoCOy2zRxizgjU6
i2zCr/El/tH7+AtbUpxe53TOzPkaEiTMy3k8rc5/1oLy2EdtiNr8ZPZIe/8SNcyh
7LJEnf1pWlsBu4vszZI+FGqYkPvD91QgJ1dkZfm60S59g3Xb7/9ZdamkX4oZA/rX
5z1sWvtNBaIl9CeHEyoyXh34gQB8z9+14mcCFtDYbCIXJaGYsxNhg1V0vBzGxEed
ghm+kqezm/YqzjGK7N8oaD2pHD6vldnsAHf0w6h9aQwY9+4c1EwdwheK9dXjDDtk
Mb1+iUxvP56Gy3t2O5ghvP9eUS2spckM2Cu4g7rbfw1IlfpKYuEly5aG0OhujhSk
4SdcWLACRaISJImdtjasntiNSyWZUwZzMemy+hrCJBuBSRKtp2IgqQ0L9OABYM7m
LSXqI924QcohEXpC4OTWrwazK+TSdkjrmF0G03/YF4b5btcK6T8HfkCetxEJLFKS
a4LEfKo/tc6A/7bFZQhNu/4DJkrjmqsaGUV6NGrgxZWHM8QrpMvE594fKiBBm8Cp
3FXiB2+rAQazsyqDr0f4cclJu4/Rh94eVpUA0H9VxYxN8OXV0aLNh8cTWobj8yKo
fIPzp4uBXFBVtsu5QTz2svMduqdgDIYQEqRcIH6WYOdPggXBXq4lQ/Fy+jRnGF4w
GFpj6cWULgwFFC8bJAVIWAS5mL2TBuxEaaXtW0nlpvng/A4zMKXYCiD09s3ArrpX
2hYQQnjEoA+FD8iDoTcQ+RuUQRgfxdCKoFXvBrlBsiz7R92DT1LAITbRI2xHLSby
NiEt97CgqTJ0CFvEh/qQKv5LaIDpSyVeZvihDMGAui3SNsLdVqy5yaGgH+Nkbi7/
jvcMe9ppvyoEDA4wLBlNYqgR+64HXYxMhV1B1i5bEUFxv3zSNABzO2VAC2/OBnRX
9xGKKCnq7xH7raZPkDMriVj3BuQxWuKD56ZKtWly4e/F/x1ioZdpu7kDE9A4+bam
bX5e7jSDJAfPQS7ec1wZL8xOQvXVzPDAcYnXusNexxy0XD6gutq0TiFc+7OXn+lY
l3ZWt2HBDrVCA9YSVWZBQRGQBamaL3NY0xH/Cej7Ks2sh6u7Y9ue6dSKuJe70lix
2ApOM4vKEPPFvfHATYvCV8pgqpXk5wYgnEjVA3+NUPr5b3eKqwUsT4SJyT/blGMe
yXJ0Sx4puRmwVfK+G75Zeu1VffVLqhg6EriA4FV17Upmx/Iown+13CTh0LhdIBFX
5ey5JvPUpFmCSb+V6o68ipWC7ulVNA2DOoW2Q6tHkHHMmbGsYluwxtRYpJxT/u+c
S3g6beZacatlzcbUdi4QGPCYN/Thtu9hCp9PJUs2LuC2YTx82gh8f8alBxJGK8jb
teMV1Bh/KWmK7mj2X258kfK5B8iPXozZ7AgBnrPr+YdPNWpAFL2mU4Zq0pG7hAj7
XhYiezcMPYDHemgcSga+dE30taNwaN2jeVTr6BnjmcJL/v5nqkUndzk3+1210eEZ
nXBQMdUNGaZPFZYhoXpD3RO3KUEU4C2pV8dIb2LVLVa5N+LeSz2eKHtesWf6thXl
R7sew65OqWSfXI0/CbzQu6eA6SXgwENrKb4H8jNj57OrhnVBmDJeNQXfCZzn5lhb
zK6ncg6NP0B3Zf+w5N5JaaojbSX2oeJfUD4Cv5BjZf829nn72ujc3QiWc6arUO3O
YhfSTpxraPD7v1ITK/nw6+9szRKCQvTtNCQQswMosXeUGZJWRVX6ia/eCyYHvAPU
5MWYw/r4cZ8Mo/BK45Q9DDCpIqPu9R/UAD5cgwKnlk2wuET9nX2Kk3SMWpatjI7B
c9gziCFZd1lSQ4IcGoci00EdzV2aY6ny3HF88eY9qTi7bfRj+L8kK4h7z7GLmkzX
Sc17OUjzyl/JTs1HJ+2gsIvaOHCDAvj8k2G8pz3Maq7rjhBXQqjnNKlTINaUMXN0
vCSDg5WZmtn7Gp5Eeyvhh4B1+J3ugJ3+RLQS/uEdL6J6R2nGwzIy1fOMR8XEfwLX
br0uwFJhhKz4/5yPmyOZTrcfx/6HuxTMQr7NtUSo/JJhtj6elsENpB8nF3n/CYDT
AfQYuSL4iV8xPK7JrmgWPecx+o8U4bS7KVzUl+Vsr/CcYmYEcNa2Ib73EUaWz1er
/y0eLlpSzXqLTXb14oHWrowFGntNyeA02ZTd1ewzCP10NxWs6YuXG8xy/+L0oa5g
FP6HuM2USlc2M7rgFElCwthS07Z6KrUnTmnY1TCAQpcwTAFlIHpeQez/qHLeyKl1
pu1QCzOW7eYzi7+6TwKeZkPaz/e4gud1Q1/QeXt2gwKnUfov5a2d2CU99t+7cvsT
YljrgEZuoQIZ7FgLfsBq79e4YUy8jF5BrxyNtqIWurQkuBZegHzndXHyqQUuvcbH
g1BlT8SevdrE+RjyhdYhPac7TnkXCEG4Rghr/Y7fWlaSchr2/xQRXC4Zm+N3EVge
DcIKoAvwP01afB40rRCAe8hSd+viqN1BMKNx4iJbJFx1ESaRID0ZavcGXU8OfEg3
W9x7UQHtpv5pJVZ/Xo3J8WEEKp1RnwamOwGNaQDMutuuXOjqTcVJ5JvDD2HwHaaE
8RygRh3QDxc3a5342orady9deW6QZ54YToKrxXptVVHo2u8Jv04q+a7OZ1ZQLEjn
2MH+SnE+oTM7igFH66T8uF66j393CLfo4V43/69i2XLkqygcKFIwOKem7o7JoV5D
EHXA6HtQe7bJ0xn5WcsnJgGxbzziL+PxLsaTg3jtnc2Y/y37kOq4tVanisIFrSdg
+/dWlXgFoHvTXf1kU9aGpPX7nEzsfemsdagRG5t7/6TMjDsRpGT08uNXby54icUc
gU1Xhg6d2SETO/yYTKXGfYrPC4oae7395/waUUlXYIic1BX8gzyFojm9tsMf/kg7
xRHX3HKGoRAKtUOA09PK2A2eFqFLA9wOwdFrEmorfGNOndGc4gKxEDW/1eTe5byv
hHowdD2yypBEUH5ZXuqeRbUXkIgTx9YSsf/GvxyApHAwmPEcc5wK7NJHnEfP8vm0
r+NVZV5eOabI5JYgNIchZ3NqdPS08GVBJ/10U7pLDQHtT2zlehJpjhsY5ZqkV417
ZF9lTPIJn/73nbtLkpam60QcLx4DjNARriWopTuy8acB5gVj24Y6sE6z3Tqm5wjw
B7aduGXqjGCv4xihWiAKYaWOdKQiNtEUobyrI3jOtohCuTrc6mvoUi3Imq3BKBy5
+hP7qAQEAbUv70aDu8++e0RzbMBk2mhGdYfRaLZ0A/AHZ496ktwwoV8TjsC+0EF0
shhIdUt6OJS33an0/fCtPMNBhPWkFb9ZYRB0ZhZAtE7vuMqC5rIz11viW8/58bHc
d7EcBFvsXMLg8Rf0FsF1S35HiXLFMfOWj3C04NSKO6e0tZfTaPHxaDd18UymvrIF
OYLuzsn+L8kdaNqvSdhA9wka8s1jbgaPr+gfKeeeifaphIsWNPC1lGRxcx6Rfxi8
bHISENjOgVwhOOi77pXBZJy2FGmfOaEj0/YAN6iS5TGsrCyipdz0NOcbp9Ndwmkw
gcoegfh0pi3PmSznJtuZ9C5c6XamuDaQHz+373g173hPjx3ZXbslYfZZIhjPX9lY
MiqXAHrIzym+4QNopYKs09gtIAkt5aNZVWOr96/mg6gD+DIeL9oaHJB3kcRDLq8r
16BqLB3xmIFebcu08AKDO+8XrpSC/nVV7fk2JhyLKkJPTybqcDTRyOxgxoUFhzOv
B9kroXU9Y1inH08SyWFMxc6TUQdZbuJbB8wB6V9IZHnnGStkpEwVbpjUu8On2Rfm
2CXPVmYW7IhLTQRwQ8yPKSiiWmOIVXYFNnam3RZpQGBtwfxNH56LlDijlOex/AG2
A3NpO1Ul6dvHNgZeqMn8+PnliIVkPHHhdiXKRq60lZiLQsDAJKuqpDVF7AawyAse
SD2SwVhl70xdsWmauAzgMuorZtVtGdhgjbOXvuShldyxnsOsOlk+d79ZIBr24/bW
YKqsYhwQM8Jf92rZtihA3aQN0octSGnqC+ypcgTPdKnZ+nUH7DajVh1AVnm2mld7
3tgPFDY+AxmyCDZSaUT2qHbOCXpgExj+z40tWyqR3ttH4qCt+yLJnzvD2rtPEU3J
MkRoTZS+CDlVPIKM4sfE3kQ8woORsSNAYDiCmzgK+gevW6xRew2gB25MekSiih9E
voTOqI398Cv7pkQ5Yxf8ZOeSChw2bs8jL/5dpR7sTUI/fEx74DwpLtyYGRruZerK
gMDaI4yA3Q8Uqq3v59xlHolR/ZzxAJC3zRTpkWQAENBtT5L0FfXRMLxmf0PDLi8f
EbsZ1uicKAIsiBJFXmNCyR232roN6vKj+8Uyg6pJH1T1G8j3qVpKKorVFPtvK7KG
pFMLR/YI/9RNWNJZvLWCrMoQOip9lMgZPOCl1kf7amhdycp0jsdjcS8nWSV0gayG
8ps2uaibyVGHXZk+kkxQDE3BkNgLaY5hu0yYlyjX2mxaJa3cFTMqCkjSXifDmlTL
hGep5HSfhIgWGmoJAxFzOK3Yt2wnDu4ADmh3NHnqDPZCr1wYxEO8B4PsRwwsdfGE
+Ki94LeUIQHy6FrPX3zVzVwZrXv0dEVRkld0bAhCj/6+20vInmsD+DmlFzH5d1e9
hAafuLF+/XfFtpXEoMvthAJWhaYUp9O1/Q5vowimDIexUsekyPLk6/Dn0XrpxfNx
gY6K6MiI9AYWpETkmgwe6PRYBG/Yfg5y5G9QIv8RN5dYwbafHoYrC+SRW5wJZWUc
7W+75/oDXNXOwEV/zyyS1OZ+ufXoxtA1ahpHTeDXe4PqRLnpeaKtKyF+wYkajBlB
xDTUZRvK73wsLREHkTzIZkIo43s5nK6yvv5dsDPWbAmmRamr/+uXYJjJxkUeC872
F0QBbb9chxFDdCuDh+0u65PXWxwJbMEiJzU/loBL7Ri9ja9Ak0XaQMiztbxm/CON
vh1ZYqP6vOaZzaHhnu2lv843hW7kDeJOJnPQYkUr7I9hTS2xd0zO7m9LCl9//Uuc
nh3tJnXWCpzyQsy2C21/fH3BLfEkmcfm/WaFOAhr32oosoZ4QFTvr6s2rbymFa2O
ELWkRVeFU+F21yGozeIroFXs4nAG3ZtfqdepAw/x9GFx/eO+te96SHpoPDAd03Vt
Xia+9R8W0d8964RxV4Gq9mWhgcrQrEOHGyAL7CAHvvMI1zuB7T9SLCYtpOlyezqe
ddTTC0zpImcb/JdDbtv1sZbuOXYshD6HsYH26RuFBDq9MYJvv/hw3kVzhFg4MTTu
fQkSJfgN/CyK3DuJiVnni5rQ8cpN/K3DL0oq36bJB4thznxX2qZesrQhdMlsPmdm
mGkv7MUC9UuFv91lDdnIZ1gYaCNTdyAQJSNPX/utzdqwKtn1+YQ3OvbpAlyFgOdX
9OmSBdqE9wSPEJGcmFY9aHYIPZFqgrJcqnp/ZTCKq3U4QaS/C/M9or/4GgWI6h2O
ChrakH5gvxZXFxtdouM9C8jHxk398INt9e8zg8cscd8+iwKYvdLHPce4sIwP/abO
T7vkeF09I/orSB59nYLQuTe9hpijrtHT4bzERNvfUX/Ky5+dXh42bwARr7vqzgzv
Zjwl2yiuNOTjDjOuZb7lyW4mPnrilgl3/gAKIAuYePd5FCTzo1FMNWIhNbkSGZWA
7gzAJSbW/HaDYcNHZAnilhUZAP9mjYLjbRn1FZLtbunmtWFx+iN7L7RohmZpRf14
MgVuDEbddwJt6ox5Ywp9wdED+G0NLLsqMKNnfshmjccFiEEz5uNeHC3T2bUzIkO+
JwOYXePL0zwhKxAwuK3ZriTzgC0669PJgID5NJxOjAqcMkuUEdehCCH3hIxQ0pKb
4XsO9Dy/K0XLkSbB99xK9yQuIQOQox70hpjY9f+hkAJZOq7IwOQ4mlA7ZJdc3vW1
mvw3Qw9Ju64dhanEgKsG5/ufyrIDzWDxIq9alPQXzR5r9GzNsqZrcoIH6GChaV+d
Gdf3NjZmiXlxp0niaOI/d+3KaEoAJiMZbsp32wVSL03/3MDB6KlK2ZyVWNDWU1kP
hM/OIBpmDN4RmvTSpwUmtCYOVKt95Zla4He6GiTmnfH0gJ+RZakZInp3YRYoaEiv
v4P9teweyTH1OTfXKLkau8A0/z/+CHpsUASCmpIxBQa9ArBXx5f7NQUZsfyKkpin
xCkVFef9nvAmXTp5YzCU52DUU0/fSw0c8JEsaa6Xkmo94n7N9QQ/drvnB69moxiC
O3Drec7/XxAB44fqBqGxv8fLj/cU27t9af2RVO2WZjgs8sKjWOywwxIju/v1RsSI
AK7mBERuBD862QYtH+Y+GllztGBMOmilb3jBxF15bn5UJf12BxR9ZDa0NsZe1bLZ
Jh3nNS4/7U7j98WTmrn9Vn98co/dWNjMow+5iUxCZ1ZqZZsAoN4cL5YgaDPhYpqI
8wIVs3zXF1Le4kWHbV14iEzeRktsAxnVH8ODYZLxsU9jYShS4WV4QvSakElpkEII
MJsUMfIE0l3HEbKQ+RKfRjqTeMZCBClVatvj2MVfDUrEdtkEOdRx+FGSsoqcrRXe
r08fkNDn46Ec3KNQ0V3FCDxUtbZlTax3Sa4Mzl0/ojlFyyX+hO6Vp3F/dTIcX7g8
uxv0/mRfIahMZPFuyHi3v4gatmwit5gQ9FPTYXmm2q4VAW9spSx1QGX1/e3al9qV
8/y6+U/PMKejQnsyLX6+cSPzG8Q/lNYsiRhSayGRDo0xVZ7OOIkFhliVZ0q9yOJb
29xyJXu+0lRStKy+z6xHaEcQff7cGoZFI1MZK3oPx/P73s+fMAf3sGH5HuLKjffo
zO5jGbi/5ydFWUICqysTunJ6QFPRV3RONtzaJSr7+dRNLZ8RiUDL/8MmEpcmyAjn
R0DKJX8XffQwXq6PsRjybDZhmi2DnTXOKo0/jkevaUdn37WjuZjQnMV/z+2hy8rc
26S6Z8oAJGWc4mHmLEgmMOD2yMJCiU+i8Sf8b3kEYlq3sfK6F0K08mMFvIVRG4mH
FMF1CB3JLjvIy2W+FD2L2dZ3QCVulMLeK4SMQ4gOBSy6TOjV+gYf5Ewg7uz5i3FC
d6fdzVlzz2O4dW3Ls4JSWYqwxIghTjkhP2TsyMyePgOSg8eQh3juUXcXmF090h5d
Zkj1LgsnHwDI2Szb2QuRbMIpDSZZV2l5Mp5Tx2jP+LZLIfbxYVZ5lRISjPMcRfwE
E/RBaxqVSQLervqy9QyvHiN4aQkQ/Fom+v6V5lWwiVooSIME0FhxPtwUiOA0eeEt
6YoydkAfRgNQmWWopsJd44D9yqqiTXO32UWyqC225mNz5+00Uc2Rr8FHn3XUXHhe
Un0m6OFbC7g5oEiSWoCZqjcY1peckPCJWYC2ILd/YFc5l0TT2nDeM+SwQaqOCdBF
rBkTYoo5Qq759CIA1E0VlbAQAD08APyC35fj2fa+mdmrEXXHip/CkMj86InrMXYz
zvyHFVBPr4WU336kT1FC1i2D6r14OX5iJnT5xQmhjJ67OlsbM7KQOFoH0koB5hyo
cnHJ87o1h4Z4+V7tItKCIdZBmqq4TzaNoCrluSmgT0h7q+5ksJQ3SF5lOJE2gpDS
k08jbtAtrtSPneoTSuBIY/dUUgEUbFNn1G4rjdHEob7BCSOs9mBO6uNe+DRvIkQf
hALjTTgPHNtHelX2gINsbUuG/UOOG4fdsg8P3sRbmdllBKQYW02eRxAQZuXzkQe2
1wVegdLyJDC187OBAKWXboGX8Sgn//6YeWfNag0x1UDMhXdohziPxJXwSX+LfnXH
ah/qKvWFORCiAXcGutUSfpfE9o+zD87KlaHjWdQZnMlyP7dw0paeWr40FceCq8Jj
PDUGSKmfTzPVtUu9sFEVzp4LIcnOS1Q72fSj4mZEwLrWHXSI/1Ww7MOD/kNRIxQ1
1QakOLc4hmJIKrvkQiIJ6TOddz0Lwn0lNnWYfSz7Nww131CEsgNLqnz9pykzxgq7
b9oVkfr8L5c7TCr+cSZH75lwXMfN3DKlSpq7IjrJmWvti4nK9BfjtJWQMrBE1gAk
qnNHuyJFreNIWrnzeW6IwFNclvVMb4CE4+GWIh771lirMTlB9oBZn117wtUNLTtc
yRDaIVWExP7VzYZr1h7bJgnRurR+ocN5zjr2UYd9GxyMYQVW5uDBh45u20rdSd8Z
diNr5KPJnZAqBLx2BSLIyLmJZ2aqJP3Y/Gof7NcDYJf1vwt3aesxU83M1JMOMSIN
Sf9VmIoc+mDvp26RRjTms50YrA5tzmfTWSsyMra7H6Jv7lB7rSIHE+Y6W6ApQjh2
ZH85rm5ZFRWVHCiKUj+vq+CbfkiwBCXHQALv326ATGFJpkZwW3tcl1vgYDLgHCGD
hHolo4y+/8rvNGaV8gKkwcOLzoYkw1UZQLE3bvBFxEuQlCmbao+hgbwZ2K/w6uPc
CkOddGEZ17Bs7v9xJ27MY8GU5QXZz0ZCobZHY8kx9CIOheIOHiERY2uZlT+1/T6u
CLLdufr/04YnYUmLGZPCDmVb6x8vpFq24LvUbtj1E6s946W6ulFI6Ipkxdbao0Wk
7i23b0oQiZ0bBchUfCqkiuikRvM2zvNx6svvzTI4e9q+LePlE3neUXyZtg1KAhZO
m0AcQ0w3/PuRRMLo7RcPvanZUukG4382PX0EtiOd/lN/b00zIHD5JtBq8S6SzlUk
T/guQlZFj2Yy4cyCayoemqZaarmPEk16tzUXc2C0mTz74KBCUrLTx6xvA+8ZsXg9
eJVCw2CqDhA91ZgCE34XOT4giHa9ZKON/ZOwQSmH1idEoRtZu6aGbko6QZN/GClQ
jVoI8qrjAdMns/61xf1UAGESoB0y3W7+9jJWCyNu5U3xZkVVBFPE7Dr/SEUfyc7A
d54KF/KrA7ivJueooEwfmPuXZqoQSfeaXidKv1ZdAO3kZ9WKHR70Mse4XqOktx2Z
7PiA3bdjHz2hWls5CVtDRpQfIxC5evEZ8oVqbqh6oj32In71ACRykrv70/N9Q3sF
28QP1jA4ldSvyAFkfjprC4jAPbf6Um3uj7ItxZ9Rd+C8My/xHYM33kHQl0MV/GZA
IbJa+w8JPremyGmtFH75XI10rJZMe1aHZ7Yg1pJPj9uQsaSiNRe5RX2uJ74O8JKz
IhH6vJL2QPXjl9+z6MyEU31gFn1yaybhvoxRp/kp5knjWgYFWynPQOAWTDgKn9tt
62uviJCo5xo2aNJ/PfYf7gTiDAtaKlxWWZxX8J+CYkNGVmojJ9S++zPxVit/iG4A
Vpa952W4wZUo+NevPDy1rRIOzr2gGPq/O8HOvA7ul4XK8oX/mgMKkzrBY75jL5I6
yRBFRr7x2/dvlv2DoOWnxILFWTc/6io6ZGXdHIw4ODZ2e4tDbo/BhLHL7hMOs/O5
AsSY0m5+/8poKlnKk6lvZbrlbxs6BmohRVLUvlhPajzZN+ij3vyo7zLvU7xPUYpg
Qg9CZpYjsPnsEEz0Wvuu22JrQmmEN1686svdxfkXO1TwuI8qcneA8V+ZuPbhRY7+
nnVQM9jx1ZU64ngCfX/3swiwENjc1wrvfTcvhAKYaqFGkvBpZFynVSPk/Zs//ieq
5LzcpNCQYmLebjYjCLfBbMm8RyGCPrwf0PbuuO6FG7/YNA/xapyBF3WC1KtAkYLz
/Fmrlvfg4BoLRGdN/73OXin9O4okMgsCEys57iv7KiV8E/9SzAvCQ2if4/nyVfye
A1mOdurCfpCQ4B504/qdFuM/zTTmcd446kbi9wC3xYHwbTVXSkYGm9luBGDEyaZT
VDqzIQhAUKWiq2XRLtB3fZ20v5hQtAxj25hGvdSO39E36xiGH1ZhTON+CLJnXGkH
h8LL+lL/rR6rFfl7qGCotZNw5B7Ub5oHNKLhFPKoElRwfEwn4mxIqwGzL1BnmVlG
m5GYkPgXKu7jOHbJKC9cSDaa9XHFo2pna03UeAYjCDf1FUX6Vs8yzmRNb8RnjxdK
75f/rFl0zMlEbO87ARZo03CyKCf2mDkhb0CZr6U5Rjjc4OTc8Xz3X7SF2dvcZZg9
i2tPDflNXiLftGE7wu0RrcHoojYQuVSDYRxD9lTEH/sGDU0jc5l7kJTI5vIsiWUW
GRacJS6KhPXpm8t71+KPWgNmTRGmQq6hOfc/cbONpv4VZ96gP6D3XY3lPM8nGvLR
BgoDYyCzrfBssmd9icJkArePK51WIy5WutEz8r0TP47QlcXdL3+KUJcoK+CdOnUq
fR1QMC/EUWJ5VZTsSiM+QffVOIOHguX/m+1JrchZ1nur3YwhsqXidJVBJfYTA41S
IATeRMtgo0hteGNz06ybXmjQ9KA+0mYOzh88L7EZIv9fJYP3B0w0YKKr1Hy49Mq2
CNkNB0v9q8RpsD1+Fu5s7sKjDJqFBIrxhvrXFFF+eyyct7QEF8WkCet8LaQ2Tcy2
QxYgg7jOCtET6dAs6AvyFhIKcyuiaF4ohzbQa43YPd1DS4IPrFHD7OYpwwzZ0zZr
fENfDlZ6HxXcjW8nGDesSe1nZr2Gas7KWCxXpbZFCEQxDCq4HdsjKMAF+lPYMC05
sdEhwmOrvDMX1BwimJ3Yb6iiakfbXXrfxpbhuJ0X2jUWo6Amg+I+SRcO/hI9GnUf
QQ1h0IX23Itqh1n4b44+YmSn2dbuA8KOUClgUoUKQkatJDLjs3gkctBWa466yu/I
WoF0r7WIyZ8IedAwxM1Kn+e9AdaEbQ1e0/y2hHX/Z3YS6dSSUR8yeJAW5pPDh5v7
u9pvZUIus6DmSwO79GUB9nZlG4BmPvNmWEDNY8zBHJsWQRcQZyNOnpcih97fXctK
qYXTbJjKep2SGA1A4MyXmIP5zNJXW1yS+pRd06XtYo6ThGohS81RuRhV2AvUvcvk
43KtZsiKmaZspEHgT+j9h4Wu9RgGEQBXb7wQHrS5l39rbzya9sKvMHvZoyTfZjug
x3ZokaoZAsG5EO60sc6/lhBF3AsH/H6qrGQ2ssT8k4VdjGJ27pKbiAublZn0oVAo
9KwehGhy8r7TidgFRnPTs/aVWt3W1MunXiVPN60tGrItIfXda3+uTVCisuV/NxzU
RVjnsnwLDLmPgBwGpb4vd+luTGA85+mqozSGycomjT0yP4Sg57asjM0QZfmmZyd2
HoA12v3OAZGybnLPpNwZcgtsSF9UiCL6RFFT0AjYl/1jEyjFbIM1MgJTm6LVzKTk
BTybfw8Xz65YzvfsVmsOic3Poiz8XNmGqR2OQ1DQAbtlJHE2k5AdHDV6dHPKGamN
AVFacq6KW2QrMH7q9/Sa0oQmyRrARY7qxW1A1zE5LopIHCO22e7s5Zd2vq0zUzE2
km6ADAMfmHtH/rXuCTerhu+sk7qGCcV3jfNKlk299k2lAFNBNVkmGenXIO1aH9M+
wIMiytoFKISnNRdONmA2YWU+YfZbm31RRU9Vpqp6UDzbLbVRfDaOEG5S7SSTGoLn
7M8+0CQPPh2o7OeCWGOPJKQDAnXsF0OjZqdsS0Lvt+P6TB+lHWICVaPph1O7CTUd
/bPdNgU9PXp7eBIkK3mu/kW0Wrb/rJ4Iuj/+QIbJv/3YJDPKrmjVhbd4B8CXImZq
iax2flvFFGUWrMAK04O5YybAymx7vJBlfoquZQ5bBYra0tDLTEmlbIPYkalK8JPH
Q9cKGYm0tJ91kdVhaOf7HH/F10kvu3eACd+X8vX+QJZM4tjcjvnM6/L9U0/Pumch
B5ZMAI4J4jkYnelziSimy81UmnVlhOtvqTRKzWFgkabA/7WaTZjP4+8takdcWqJA
WAM4JeWQlIKDrKbu2yUOUBGvvegMZLikoVq10/rmf0K6seFxTWXcEKA7WcvgGSxM
73tFEuWZVsqrArnDJMG0GRz+KX98qOPcA9Ssugft08P+CTeOXA0VGfVNIqNToBaz
a32v5s4SrYKoCRXA07hFaLW5+d7NwfS/H3PvXWgxlSslg29HU4GWQEwsb677JVnr
ngYTPGs6jQqM1Hv20SNlQ2bkeb1NO39RFC2PNl7Aex7iuOeUPbqgu7OhkSSktE8U
lc32YMmixFzHjwwA11JSUm0zHeDoNHJxAS4O2dUYwps/Npr0Yybb2PrJl+g+ZP07
+i0KoUlbMPEiUuJoke0MdPwM4LYCz7qP6u9QKm2cfl/kOoLN5qDubJA6OhJ87bHg
PRAfHt3FunhejPUpTHK35Iqxg2RxgQhtbxzGiciamQVKh0pFefgRGxi81NYgwgiG
s0I0ZOniMaUNhgjfTs3I7zTTkpGNPIH+HiP/TsgNDpOg9gvH0UodhhLzJUmR9JMl
+N+BibFk3fz8xJwct7JCRKwZNHUcnrGh1FMDXCVJxg/NlWPtLH3Lcxwu1BLJk9r6
QoleHxMwoBrTMEOs/UxhBT9Nrl8wMv9UCxtQjrZw214WiUnNHTOyQKMjMunorRgZ
aKDWN/vD5QiFNSkL1ye182ONsoOFt26zy70YGcJ7kKe5L1YbMsxUlk+YZbqqvBsQ
HNVbE0uo5djQhfnwQ/PNrJLRMbmg2+ZTGrrOShtJwpZsx0zkPDa+1CU7SrVwguq0
2iGswekfBEOgGSGUy1cPvb/rHh0Chu/W1bk8ls8gqSip+DI6YnOMZLBx7nV12lAY
neTsnsTnXGQ0tRjG0i/9ZVzuSBjThiOMvm5G2RgXQAiD2rrTx1O32Y1wutF9TOMn
4dDenL2POQ3IoTuZJFeCLCqreerrtcu1tsLsRGtRbrSMRe5LCTc5IJtYTAJ8XNLO
usQtl48ap6TDH2WfNbjcr4pS1JIRzB+3sToX/uUqYNGyqP7XH2Bj8kCRt2oSOs+O
WsdAf6nAfrz3fCoyddiPXSh6IkRRnax0D/Yjbuk6GY4WMW7F4BoBN4BlY3GFKqfj
A3sVEWCUbfRKEr+4XT0UlRErurW2j/sqQD25auIMt2D7lByJasdHIIHyv3YXTPzp
MsVTIrH8qM27Gy8TVUKx8i7OV0E2OP7Et/HkS/8Y9/bS0oE8CELoicm3LxmbnAj8
fxmHDGLjtqrNS6yHqX1Z4XriSctYX66eBfKVYf5JjcuYIgKv0s80EjIETRHjg8xG
ryBsyXCB7ZvmM7ZPMWCCEZvkRNHhwi4xQ3drJ9XtxPnlaWiW5NA42ayLJDyzU/zd
LlXX2XX6JgZZOKBw12x13NDtAhRuIW4gSe6EzQM0oWgVTm5JdjefI9zQWTCaHs8a
mVkrFp7YXMZlMA/SdbEx5lspyhgIuBnUKLQ14AWkpU4+dsRRtIk2TuIDHW2oS4L7
7CZUmDtdzjZR0JysApn08vsBy7ZNliNaf0dFXQT+SkDLtBivQkgXtw+ASeSX2V/Q
OI+wEbvM9dcVGSkXjn5eXW60NAHFcdMe1WFKD5Yb5TVEGu/dSw7YtH3KjUagApfQ
8rrfQyW+CM6pltsrRhfFJAH/RtyxitXZJGomb4JjqEuf+3o0Dc68KlfbO8ROwBMD
YFZxvzTF13zKLHCkcqNQYH6CXu1vrncEzq59yTMrT4WzpaXXiFdfluvnO6s1hhBv
0AmL1fK4aCQWc3DiUPHmOCMVD8DondiijYktzLONYkOZ4dEJbPzGjYQIclThHI7k
Tebe1RY9JpC3oBJF1buiD3L5FZ6sqb/TLeYBXKzMSkIYLcxSXqNnQMBhkDtAWMHz
3+5E1v4ssTvsKKjzwJbboXuhPOTYj4U2qyERwKRPEN3fYA+ed7JiWOre5n3oLzH8
0MB1t/ZNbsB1Mk+/JK57mFEhY5TEloiQEAbINH3p3Up8ILAcK+IBSnxxQRPCekkp
o7EQqemJDxHvR2SY4lv4dz+e0r+ZnwA26A/+yPtxPu/kKN0IEpejyyti7+MMhUn1
WCZZBUKjaITExlvCltOU6edMANguNY0iUtl7X9aoEY6phyrrD/UNvH6kuSlkQla+
EA1756nK5PcWwWXcjek3R8f3KUr4BtGPICiXRqFUQHcIbmecpOyG0S7CgIsYBOkq
hkx5t1IwgU51jLrGCZtW0dxHlroR2sjp88SAMv9IN0C5Xy2xWQS22PsQehWtqkd8
/W8H1uUpWvfJOlxLEOXP9PY8R+v/aeAcV6m6DeS61zS88Jw6JfhR78BdJsaCw8cX
OLI2ZkFzxglxSZex2J2hkLzZovXwDRDG1NmHFb+fUgVQ1tDV+T9BPU04tlaY8ef2
fJNbyhem9aWcFKpT3iO+7GfSGcwukPe2Xv7q2I0FcA7AER45sepXVOvk4yqj3sjn
BvNBZkygnbzMEclJf6x5snZJw1auadyZWUNRl3EVGToLaacvxu37fspgFJ1bLuWR
rWVD6l6SQFP9Ec8X52f+aTBMGYGq6JPe0i6ZL/yZw8SzWPV4wJbUN7avrYqvTY7I
NRo0rZkSGBUZkfaP3bN3yXF/KOamE3Gbg6/hFo9LXjLkY+8u48A7eDoKIqbqwGb7
dcOWBInvVyAtLCdBLiW6c3EihICOFbmzM9FsNQ4+GvovUMF1j25UUzp/s6ACKpR2
oFy9741YS5P3L6cYUYv6eyzAuqFhUTpzLnvzUfbiVDB8Pxwm6ztjxS24/s+07YyQ
ymKbLS8iT7AVHNrLpRghepC1jtZqJDO9Bb4otBDvWbZs/YrFGFg7A51FhHMJg7p5
6YSuJ5+HPn3tNlMYmo/vJRD0CpKVU56GpjmGlXWQViUktej1fDPqTaf+NguxP1NV
RFU9QxPpbPwYSp2ZPx853DMEgafxUi19afAaQAIlggMkpnPgGQAcxqTNXCXuDS/P
ia6YO4rP535EllNe4GiLrA/dnCRe7abxuAVw29ekMGQdcC/v8iX5B3oSo+ZPgwV+
Y4Z0sVxMAZ089wz8yRYK5jZGPpByOKteg6VNg2rYMN8RrrDnPTlmeIunVCpQ3tH3
n5f+C4MgUlWljNRGZ/bpqpXGWGB31WOgQbIntRocYF2e8LVTyJGFsRWYJDAnr/if
WTjMhePHWFFSpfjFZe3r7GDLDD+XgMjxIsWzaPC2PgHWELaRUphhO8mnHR0Xc5/A
g4DqcsKtItAAlrTej3ZisEMnGE0o8ANNy/Ex8htfbaPVYRy46grBe+TInxtGzQyb
g/w/8qeam/hDT41/YdP0HmWDC8XwuwA9YMS+39+HTRrnxDtmy3Kk7/185uaKnDxJ
9pIriVcuTRZ8wbV4sX/ZEhB45qic71ab7xKnufUkLWX6xgOdyvsv7JVKzn+JFM+f
nOHbVbzwq+/UaRm3aGRgK4XhihQ8+1HV0nx0/heoWfM+YzuHzDIxlu37nURan4WY
6Qnyr8yrrtdBNjJhrRwT3HS4Kn8CJIjOALjGFgnd/kfpOND6M63L7sBvKUlF9NIU
rMhJkcciguE3cRLbINnTJf6Eo8yYBjkJA/Sks7AmT63VcKFGs1jqD7Yit7Dm7BY6
d5H2QYDY1d0/uAvKEWskLKeYACWYPUYyLuaiFgk9FkfRS/bP7qIFV5EQfqjNZ+tD
eq/r6fh/yryW3Wo8pGUh/YLBpKewQOJJhHNMOR1FYcO2vbZD8BBfu806EdOa62FK
wk/GcbKlRqWrppJCRKxzCFKkyVvPeqHPQ8T1b4Y2JCJRNtVGgaD5ut3odIs6DGRH
QRAP/VMniXa/8GFQDZ8aKLX+R8Rr+l6xyqW9QGewwTgWBMHsTenlMc1me1gQyCJl
/gAEOT/DWKWFFxHRDbebvE88eDgH2TRJ8ZXebboV2s/wrB0VZI0TOoBDvma5WKii
JMongEg4wfn0ogVlyMteuceeCy7DE21we2lhQjCsAdKmAqxXkNLCAy5Mkqxl2bO4
SUL/8Am9J19LB7LbSkVhx/Ic7Uc5W4C1W5drHE7IU717YP0/mlipZwOawWmkjYcs
nZNJG3v/b33dChoYUkT7RxLAoahOFQmripMAbM2S4ZUcJXGCHw+p4Ovi2hrVa4NX
lVZxWW6G9SzqgwrdenbPU1TePkfsjqsLqO/wB+QmLYTaiLUQKMV96hXylUKP1t0Z
zUhot82f6hERNv6yPbNVKX3GSjw6i9Z+XEnEMR2h/OxMX60DhvzJHcECOSP6yp9m
YaFxY3Z4Ggj4zJCl150+52zHBhS647NYTUC4QiyqqCV6ezbAsSvqRPleh8tKmJhT
Uc+9oyvDyQm/yv6NXuPjVStHpKdY8YvPox/8LoQ8gKJXG7TxsL6vP6nKsiBRu0mO
mgdPnOOotRqOC8lXbMLgufvAsdhvvWchBYSEeq2u4c2/0VmZclKrtZTlesNkQ7bx
ZQWb7EkhluvsQuJTWXp/lttFg2S2trE9nhpKg2kg5LKX484XGBd3B0hv9X2evrLT
OBPKTmX8Z/krZ6doNG4ev0umgyTW+GsnY+mY1leJOpdmMN3I0XMMeenZpcSgzwL/
HbikIOZzNEmIk6sIicoyIPX7roGCT2gMLsYTslurS1mc2rKNh+QbUfgyrnBO3q5A
kZ6K6eqnwE1d8RhiJvxPYmXHexozCXO7N9o7rqM7+b9TM7OjTOiIlyknatwNSnmw
U8FBGLl/sCV6Fy0W5PjEOgKV28sxviHeOxIzxsic1rF98yonvnALw58P8MU2LFw4
/0044wt4Eoxxpg1iHtaqSoGYCEjxqQVd+07FqrMn6EXFT6GksWCuyUgd/861EEJS
1suyjwogjXWcsifHTcFiht5pLZCjCCsG9O58E3CzsSTvTxwwtKl6Ivnd7yibxNrN
DVCqSuzUkBy1AuJ25oXiEs0TVVnr/ffA3PqSh3KevVWoLeaYTqHZ6FxZgKHcamvi
H9e4QJwhLgwQIEwIQ/+wyyLOtutaWTQ6ymHXf5BeKr4X9F1jZkIgNOZFyhWVD9Ws
kUFVmM2QQKrz1ik6uGrKkBj7YhmBnHnIeX88K5IQOC5NlKDCCEgXfLT+UUNyJuJG
v/3v/r6rNVmLCP+8wXuA9ii7lubI7P8DyBH15xQD4XsQDmpx1PKI5u75WaoktIvJ
FjycsixASZnDZOpQA29i9057r0qMNoXMjgn3cs620okR7bdCalnpkqhsZKAB8/tr
a0WRDn1XanJ3CDLnehjtMNij3K/E0jdVQJcnJw086TEddY2xlQAvEYfxCl2ViVQN
nqf42/M58IRuA1fEuzRxM228rPBEUt0g1+cXwOQqC2G625bbxpEoso1umvJSbZbb
8wH0FUdIbQX7tnVdF+/5UQrj2OWze/NeOOL1XLpPWU0Z3tJKYH0kEumrkE0eDMIt
9s86flsghCi6ssqCUqz+Xo1zHqFLbuMm+Oyfa4+MMQFukhn6sehSYLwdUcO5ZY+2
Beso2eoetLMfB0Y3+60NHgX2ZWc4xXNRGl3JM6pot3VOTeWP01WogWy8qvFwDXuc
J0jpDHOyCc5mxPld+FRY61yGbs9TlaeUpQP2vGjdy2xGdky/TC2HM75EUN4yekph
E67/RthlTn2tVF5UjkNYjC9xFXHxITeMJQ27n6GSamwsxxRTeINIeUS9VXfJocli
juPbb4uzZN4q1AnGRsz9AqjF3O3n9e2axT48B+IQdDObcYPsKW/4MM8/1ZfmTmLS
QrAoUIzu6qsVqwbqQoPpzvkZzWFDxgG1fQk0L60YTTvsiPXPDfVXuke+jsnQdeq+
htLVVUwgn86EyXpcs/u44dl0421OcQCL1QNyzU2GsSIV1RrInNjt6D7LXVv+GImK
JLgXSFykD6oI+zvF2DVqReVUWcFp4rF04d+Pge+TsIVJmmIHTcgQD63GhOEtO06K
Bi+uwcOO4MOHryvH3YwB0YtSXgPETHcpyVtGUL4ldTGu1NBB9fH0t92Hxr6krwhD
X/1xMkUx7EUhJwGsG63GgDQ4Id9GuAXw+bmjp/BVTMdKNYQOaHBb+Scaw4x6/9hR
9VdXmqj3rN3oPfDSbANOIm9bmsY3Pz3APQMJnHflgL0152VB/2MdhLRh7YeurvBF
zxluYO9Bnp3cD/6QRvBMPcs9GHsuacTIqGlXDoB2DE2nE+vwm8FWN1qmIzS3yesF
bNqy1Th7B9EPq4l/87TMCZ0eScRxc02RuO+QwZL9xbEKnFh//1siKKCEa4k3aMGE
JRnPG0BjplWvdGex9RuC7XXkHsD/c4qYR/4+FGZcEqCOVQdiN1xQVQo7k3OGmKXz
p6X+kcsiPSRSpwqdw2NirYWCh4EVpOHeYEfospBQTtv+iXcXdJNlmt0w5foVhRa1
D6pMToZ639kxToipx0vR9O8b6c0asI/+Ev2aKMU3CmU6OriX9Y20OY0UckdyThKY
54jWuR5ptJNJuSK+Cu2h6ZSmTIDRv8JXLs6OiXkmkv8E3I2+5wkKKnbfji60w5op
8+ERFVQLzM2JaKhvHJoQk1PBPsUxu59afJjoR1AnYh7D+XgC3lkTIdp93kzz9l/s
mzC/KxW1fVjaOC/j1tK+dmxx5loWQN5EEBaKmSBliilqQUPnG+xEduwpeeqptPPk
kt08eu4Gk5T/arnsuV6lWzqVtSH2mfygLLlLSRlS4ZA0wbYhO0YlsiAO1rAmAO4+
iquomvjgiovuWKA9kaErncACj8BzvctOI3q90ya3jZAaX92CqtYIXJBJlt01MVdH
DTYr3wjLAsPKtdlzNL7IHNJR5+3e67qitB/l5Un+TWj9Cot3N4NiPSRwHmTzFBP2
Nzfm+gshg5ZOpAxeE9LcjhHIiFTsQy2uFV1K9WLNP46I57wZOFqmqIznsO0jY5rx
wFQu6ylDsAs0/oKJ1KhtBAVmmEs49EnNJBXVjWtk7dGFojn5FZm+qlipiJ766+xE
J9raoRuv6g+i5G8Aiy49Ch34EvX74JCUYuTkDSSgvoRJQDa0d3qcMQBSeXJBG4HW
S4T6lXeDmz2XApzlsveHckA/7wIKexXVY0v34HAL5cjmvIGIAYqnmyzk/88i1odL
Rc4melR4RYBd5245mAs4cch6r8rB5Mpdn6zQy2omY80nsV+SNiOqLqeNqDWQ+MmU
9yMJolVsHgkcoSFarHhE+Jt7gs8hRS4b1R4gxOxfnuxQa5wsJaqBGa0trtB67cel
Yl1RtO7oqODpDBdnpXiPrcv3MLKAxzI/rKpN5eNH70MYGh/BGn9Y/QVKsld2uhB8
+9AiXOVX50j9JzZyt4AD/suwyLHupunK6BtICFQSvN/TkL8Qsxki0nNsk+lgUSkX
jySzgKF3u8Q0ZMr4D1X8C4xKiUmNGAgVzMMmB/Oz++3+RvHZe3IUoDVs3C7jlDxH
o6kJCeNFPd+mTWKH+wuqGdK5YEeYGtvSZv3rBKxXSfaLpxjIhHBNZFXRKHVvES5i
upmwayBXt6lL/eJ0qiuy/jtaTvqYshVdjTm4ql1VchvRQAD4VE/BsIBRhPnY32oF
qruQgdjbE0+bpmc05mt2MHZ88Y7HHv9GO7Ofhjt2W+hpvw8id4fx8BZeS+YA+V5u
X+vh9FZYxxticZOjQhYFoUIcwNSm0HkMUscTmahhm1+sUKXeCtAeFVr0DMzV6/Um
ubcwPQi5Yzjb0mi6p9cneoVRqYAK1ampFZfQDYoqbsFfpInPpe3PQPO3sthrkpdh
4CHM9dMZeQAnSHXQElPg4DAEuAzfJ+AXzKzEVmxP2BcS/zcyO9cZszGiDLPrpF2R
ylRYUeE0VzzSRPzHZnEuBziF9S14jiFjtESpRASZDgyAH9iHklwfq/IYkgVQTAUq
Tlqxw93nxtMmUMpxSWkMdjRC40QC8e7rQgJunIhrDMLTe+yUOTPS1g4wD/buWbIL
27NcdDDF1AVE++QhfYo152r1/zrdNMFMxB4FpPWSTYMjKEb8F8w+ixxDd4zlW9qI
OAs0u4lilqhyL5biPhVVMhkoHn4NGmgttg5w1TlaqG3z3HCcsPwI/1daz2VaEhWR
w9jJtY5B5OMnio42ncE4iN4uz88p/WVoPnlFp5mEwqCV+TQfMbLpEGB8VuSvALab
hAyqRGZwi3jqblhhU3S1FrqXFIUdOXQQqj045WKRdrydygw8zidLE8PYq+twd3tg
1W21NJdPDKbssnQ9v3d2nSialoUELY5zTgvhKgxixk6nk9/lOPzNuSUERn5GNPvI
176ZNknaqLDNZRHOKqrlGAZ/+oemnRnl3CvtztqYvuannEhIAHzob1pTeRc/DFm6
Cnonw0sbOv6W7tOLF1Os2AfEOCsPF47Ic5fkvqVMe0N7NP96bxkaCqe/85z28jbr
FEknqDigyQoaWhDmzMJGp9oAu1JUrlZqfGrS1DX7tihikpcVvF8/+6o5RG8wEppo
/FcmNO41mwr8xA013uu1v5f4H2Ulz/vgxGEGHVG1P6xz0e7rgZCI3gwzRCJiNINu
jI+T6EfdWVfvKeU4/iR4R4v9XBCm7DIjJDYdUWYGNSwZ+yDGXlw5YzWxTmknc6KJ
cIqvo3bypAfMHTY5AmR/A2hEQ71FyArBABsTiTCLJae6dpyVlCPXYvX0zejCvMk2
DfvexeMTgYaN5Wpv8hufI/h8+uEOp58LaN4UTiWW4xu81htgvHyts+Ae/l7NOLUl
5px1q5ZiLch2YYqIhWbiAA3Xa5sE5FLFW6xy19sXX1DBsnO2TuuxWkl0iYBXthGO
rwtbZDuvM14KwJjZuHKCnztRS5YAjbWUfvV+olwjthXIk82ksUTIDh4JW0gBi14g
MKifWPTqC82E9OczsylXLqaDh3ZPqjmEbKOxJRFtBmbPOvxYIYiANeaVyg1QElrj
s0KvxLFw3ESOlSePYq8wDz/wspV3bs/UvnpLfRWs6D1Xmkw124aZBWCDel5t1FQW
GTm/ty+8t6WHum19bo+EZo3iWHV8j2xxGIBGDRRh02ypWxMjLaX+uT23l/dUiA3m
+aPNtNqA6wirLE9lAi/iaEzarw8/uUYzQgoVTqXBAZceR3cAUkHuONAAfQOAoy5m
koQTkGmdtUd3CVCOSkCHBBttNQeldXDDeWbVrQNptsY49VSCExTl1MwPYDLm+ti3
Ddw3Gj9paEFdJZ4wG8dIOupQIV/+xK0b5LQVXO9vPeAXGHeNPw+zQ9eSpR79Ysxr
/9PEv1fo3ZxPN6MoAupEalrZVtZwyIerZy9hgvK9fK29wPnXoOU/GuKrX8yYKWll
dgkA/CkEyk7glX/I/ivy2e0YBHDOwZpmbwNXFR/MWtmBtK8zy8dmbucIODMLANK9
LxFuOOGPKNuHj1D3dkNmLPHP9uMVksXpH+nhvU3IFW+SYqU30ToBNY3wxyfF1Fyx
0jQj9tMQqeQU3QlwhemuQDLUTZcmVFe8MFcTBag5q73TZAPz/ZACESzfWFKOzitW
+YQZCz8zw+a70kB9o4p1VMvWqFJ99zJ7kg+irWqe8puIm1X6awoEa4qmjLHsZJyz
BSBv9snsfeL85qBdVVuChQ1WQlRFaInxNMiPep5jUx1LV0IIDUJjc2T5oSwv4iNK
nOZe3ja2vHqRDKALwt1jIiK7tVsvm+hTcLnVQ+RnI3uze8XqW9mwCk9SKbXsIccX
nohAU68nDdgcUH48YNdSnjHx2pDDeuqz0MDXnM8/RxIEiAlXmbnBp89CpQqyG0Xd
ggPvOytEAgaESnrzjWppMOx+MbScLiLLQprIJcJ6/GlB6ATWQkrxHp35bgv7HiKJ
70oo9GmkqFm3V+f5P5D1qrfTlMyMlJZOiEMH4tporTWqHPPoxwjJOegBg9JeDVeA
MaO5Mds17Qjf/O1SBLJKZ59x1r0usb+Sl5uWxkr9IFYKi1ijSf6BM64Hb1bxOWwe
7+Hp9peJtBGIPr2ZPCfkr1HEta8Q57LF0FCXE9YW84mk8a3w+hnxcDGg1LsNhVqb
NzKipCX2COK/q2oA5qbCoEp7cpYOK0vnPx5nhWIAtGKDCdUIZz9ic53Az9RuIql8
y5t0U+ZtTOrShOFZ44qaH9o42TLAUa7NO/Ozw0RjfRHp46jRiRK5f99cDqCa7esC
XMv6sbo/HljTZRGaQJhtNrxN2up0LVUFpC/tiEP8+6iG+MrqsFfiBTUyBQvq7QUB
dsanYsbfB7pR7EyylS1qakj96fxd0Q/ReF2ZggJ0rpziya2zTSo9OrwrrkCOK1k/
mdtZmzGhU1YkORzkidjY1wUhJQ5NjsHQYCqhLZG9LP07o0YlrlR48WVCLj97yHXx
k1N712q0WLO1SwcSnVp10LgQH92JHgXlK98i1sDN4+qo+Lie8rc+4dyWCvx/xqyR
eZgjsOWdg1PpwunqWxaJJOtm3M8A0LEl8qTnXKTzmobJ73SyB390LmGBStjZltFk
9myyyqAXGI9QKob1im0luyCg/3wJ2OFlq9SZcw8/Fo6SjIiwCl9KGzNv16O0GwDA
uCht7yNAi+bb6QIg8G8y3t96+Vhbdgne0OVHn236yr6UmTBegkgIBg49mWhkL1M6
AKofPrkdkbxbtg+qxhy/nwuc1xLWWxtRWY13q3IfJebrA+moZPQZJTbwRNziQUJ3
Fzaqf7BTR+8oOZZCBdo0/ZAK8pIiFPzNd2SqwhesL1yuj4S1YcDjs/W8MK+85fc1
Z85VKxtwYndsJpiyS4wSJ024ScV6k5szO6NsDAV8RAygl0C8S3V3k9KoXfnDzUp/
ZsJqWqlo9eSz7Is5L516F+/77QOQxr6vPwrjJvSQ0CTBkRiivuD17ny5nO6DP949
jdO1LE+Xj0A+KhtBWU9fsmFBWlnMTH5x92e4dmlbn6F0mkmU/o35cSrSQLQQkrnv
KfOU6tt00FxRlNrkV2rzF2Ezql+v22adTQvTNx8jM+cb4NXEncjCnXsFeywXu3Te
kEe6EXTdXc13IqA5TJT0fCJHKkEk5/URWwUKNP13XzMUMfR39qxqCE1H2DvWH4CD
Hoifkla7SCKCPULfLKr2YQzhBZ8GmscAsLjIvgMG1myCox1lIH8MFAjjcLOJmoeY
4gGKJD8ihgxEECeXOlAlfXJMIgg3Y9KaoHW5eW9lrpDCqq7kRzqws3uYwbwA3hYx
6EN57mslDhhvle88VR1dKdvsLdEuuPw0bHd/o3rTvWg9SzhzlSteNOs0wk3s9TJ6
DsyKEueYa3MmSvMeTMF2N2JvhIDSwR9Eo0oVo9qG2L01eLibHapV1hFh+tdbucDU
1MBBcmcJcTw2zfpXycJpr5Tx2rAmaiXwL7V57UVjtIrT9Cf9zW7t7V2w4j1A6Jla
74oV0XaIIOzA6yajwCt8PCKP0x62ieeUM9yBnUgasuQb4nb+h9mjD17bIkDbQVeF
0ja1i4UoZEH191gWgRZG9eTaL3AXWjGtlZbKAJ8q2aWVJiLtMSmONEG77HmvnQTm
FVedVHp8tF+O5RUW/3uOEZP896WWXTid4i6Il8uMnRYxbDSEuFHgZjB9EkAyCpXE
/duAuH1mjbDG3qBWKicYnveYDQ3sB9cCq3KxLDwp4unfnRJtXMjlHfeLUaMfmpbt
Y5HfHbhZzcO59c5Nf0N982kKXbrgulbrRdewIUEiE9d1phHOj/9ETqvNlvmPUSOZ
wMvwHXlzmXpCnrtb1b2t1xG+5TNzkZOwu5vhQ7PZ5VChyfIMNROhPFVJa3jNYC6+
VkzAFUwvynplagtJVEBi0g4/8bAHFa6n0Cf3AuN7V5PNQ76Fx1bWv8EMFO37GaM2
7aFRqqr0wvWzloBxoJPX20Ip7aYk6fNs8K77qpruSLNljczzwX2INaoo5XekYcMU
TMahCSVjPeeHoHJOPKsZlcvpe9c2/5FHWqW8LxkXSeYlQEAbccIE5OPkWPF77vyr
QcQMrjJi6brvbpgLHpAw7S+8IB9s57PAmUDVhMCjz9aAP/hPemKC9G+Bsj5rx13I
gOoJOf3HODK9hxe1EbIiX2mHTl4CYJkiT+9qRYY8/BXMeZBEeiqJdiJao05UPPsU
wyhKjpDUvfa+Jz5gZnl0s3b2diLuftzD0XyujAucIv8udF5Jq0jgymTu7OpUGr67
jnq82SLvO0n/AQdqNkhK/P/SsmZOW/zsPUfmwK47DxZmy2ZSFu3FrW9rC3tNRXUX
tgaxjI8pn6B6ks8JEepJoSM86IIcW0AZnHmUHLw/aVYOA1oocuyRdpzmrN1+GLP0
5PPf4qvcbFsbCn/54Qom9ElNNWVkxJGmNt1MZ7WjKGVLjVMOXT+2lLnqWe+dU/p2
FeCG6gmpyBzljt9v1MUS25N79E6kjobDugQDDwnCKNClFt1hrmnLRztgUFnfP7+d
irdIrKUK7AzjpP+K3dDq26Xyo/J+d3VxwVYJgMIqANlhuUnBwMcpW0vq9ch6EnPM
leAO+bP6lt35JmOZXaCxVPhbh0ttOgutNoj2kysTQPVBcBtAabt7HBrdynGBBC8Q
1tmdE1cczDW1fUW5bJjaMKUDfLgqmZJO63pQhwcReAiAgqL8JRalYAd98z1/BFAM
lLVZ+KAKF3S2gcqmv/rrppRrCjjWyapP1XLNnDwMleWCdeHZAJX5qF7WynJotvQ8
ZbgbtrSp8p1uAPB3T4dkwC2o63Co+4PpIvWPtMJZgTR14/2Byo3wLDIJQDcLe/cA
b2vzr3hna8jQgmSqo8YYC8fL7OrZ1/hTU8wb+xCpbL6kxTNOtZY8m22x5Xq8xt5r
ZvdsuJFOWyN4dQ+hNRocyWFClVbEbIoCwg7eD6eRmQvv5WKrffbLaS7kEusgm7Ts
HMlIG99CJGa4FSyuXQhstBJ1fyWFWexMB+/2TXANiRwidiCsaP/62HCYUCo1wwfg
RQhnBd4k3kU0850HUr+1p9FrPxeM7nKEDtvTP7KBEGYbWnktSdoXREoVrEjHtWA4
2qt8oPIbQSC1h/CvExLMvqf9tRqKFCuhh9aO3ylgKc+Y+k9jDFKMHwdKWBUzDw75
oY334JC32nCSbepx0ZHdO1BjiKBpT5A/4ELu3guMsWDCrxQAANF8HcZbYbbOnSgK
zEBeH028w1z7W/hzY1gehPqmG7XGDC9xEKcHq018oos6QYwiHPm8BqA7jAKXW4+q
8wgweAtFHJmhGRSxsd+8xIt+dY5EYZlK3my3eb7kQ4vfQDiHBEVR0MPV+QByTQbZ
RTD+E7MI9Ma6PlGt7khRZovWecxLxGkH7cDqOzO16vTwIoL1PS1RnsCytEvmQ+Xs
1QAjlkCKovZBmF8afyPzi1bJNNowGclE4yo7sffSlPhRUbgFpDVRHnWGXPHbBure
tj8w+I08nEUaVCK9/lYcNjWqvQinEouQAasvQRc/jhZHMvOPf3Z9qPMq4ZloY6Ox
Xd67oYCgZwADnmf367AYZYPSuFTLV30iieMsSYNwYyPQJMkxBvnG+SjcqYXBjFPg
B/8Hg0jH1npKnBgrqpUFObZVXgJxG1fwZXsBgGerao0K+npThwaFoNASginXXQRq
4sI7WtLUyj6RHdar+cVmSVHgWsVsGoo9BAt01kCPQUCF78JwOQMi7pjUOIAxVtKF
awaDUoRRfI7JghQyE20uSmjSM3NLECp/lNLv39ybt/6EsxudPCi0Uskaxfxos+y6
5uJmx1CWJCA4O+lQL3tE93DZs9H2Oo3/3IjwgvcsTT3H1aD2XDXNPD+60UmA6tVC
K0u745GbmuhGDDcg5PcWIVYbuOB1dO1ZI2doCIMP8v+8jB5R5wEs4OOblovSDiCr
WQzu09/Byb4IZVOj6RbuGm9HcULaN1kYXgyKlMrFh5DsRoJdPXZx0nUFUNBbZsv/
dfMePdTSmzMPOtM0sr50PdaBWIVJ2vxOyzE3xhoTmJCdmc2HvGtyMyShVCFjK8kZ
zoYcYOLkAqBTrdBAxInQxNUCdb94ZypvRhn21twK9UMO5hSlGzwODabELFq0IiTU
QDZCkS7cU4mr7N8QlX45PluK/IvOwOJtmLPhg20KqCKfnaME2D91ZZ28sIW+KHA9
Dw/iAc5wPUNETkXntYcbl0zxmHZbixdfmWaSqgNOTk2c2nULJLVQ/VU5uF0Z34pL
X2xaL1eJoMCp/bZjtW3kcutbseokoV3sh0V0sHyL3xUheiA0mfckIO9iAjU7Pxg3
cwQsPGFu4jQ8y5U8zJdpP5GZX52Mi9kX3Ye/OuVEUFHZT0LJ8McRndy/35C9IWQf
nqw3yqgJ5Z8wFGrKBhOuao2GJ7+trxsqomhT5XJzqlvzvxqtBt3DuTVISpkwDH40
8nVWzW1PJls13R0VJC88T6sJNjcr6rSg25bnRdwwfhoTfxBHfHE9N/pGNPLMt8yI
HFNlvwSXqfJ1mSE7W/tXniCbkFA/K+XjW0CbOae1uemzsdF2cxy5p9KD6vnxEgQv
9sVs/IBTbKA8T1SdyRa+hiAZa5UcNqYbew4yM8dIJCk7oz3Aq/TuuWnMaaeWdU+t
6FKoomYZXFqfDbneFvADe96WTflHQGrBxv0lJjR11WbeN0xJWgvHmCfaurMID0sv
KguA8t9bUygWunm6PJWfJEhmVcbsgl9BDPdnWcMOvIdK+/6eSIpxgw2LK0r2Ur+d
iC3UUHimnlYc+RVzcmdo5S0rpi9hqYXkdjcDjE3m103UdP0APo104rT/t95KLLxg
aEmalEM/YebTl0LsYC+REQmSSdq7wFGX9hc9cYUlmqi1UIRV3UuzRfMLGx8N9r6g
NrWjqWiBDvY7X3Fo6Ly63ApHsseM6K275d125RyTvgYQT5CdDZGIYV7EXepJAD2c
wwyVLwyhn7fR2Rm8PbCwyGgVWIbtdUEQVpqZ3eFy1SGWd7aAjzvsJ/WTw91YwZyN
ZMxuNEiHBzTOIYkrGdOm5SQgRZH3v0hrK+4NuB91kJwu7hO9LpZL3nb91SzOt40m
A/X2f09zC4ojacE2ca+vz33JbrylpUSmdjR5U3an6dOQz5mFNkntLPUJyoDsqjnt
O659/gNyN2YfD6RU2lPSA3ZXQNitZ98psjVHGzoTDABf5aa5XqG0ngdh1c2RgMEt
nvpBQVv55Vfyqn5frNTaCvSS/pTF9wyI5+sncumxghxlzLQQpUh01tQQjBbgz0wn
ZL3uX3qt4N0KBPLGYkLSw+tLDHa6oCRxdXSkpK2QxXDqk6Bt9WMkrzaYRlMEvR9m
QG3zRU9SzPaFRv5SwJ24Xw0d87vZaAUYvMvZdXCPx4gnQFeE6glSUYBuBDoLY44K
iz/WuEVZVMyjHSeddB7yLSigVewguNtyngy3QcP1YYLIARrheH7QYwXvGH50n+Ma
lZF2wUkrW+23BgQmXrlW0Au97ZBXywgkCTnsJaYFE334PrjHsl3w3E5VJ9CS1EqP
n0jGorR9QUJQc3jMp3QoGhzEIGvw2/5s1PpioP47B7r2SAiUfe2HYY4OvvoQb8Ou
MzagypwEry/oJYyXlOg1VpciBfRu7i5vbEcJqpXWWZkJxPhN8rhfeMecOJNghPt6
y9nlxhu2qIlBehu8ku1X/8sVHYdyQFpLXF8Vl0GYXu6zKIxNTLQGLuYfh2C5GGVM
UzamB0tL4EMx8s78PdY9++jIpVc5lJsBmYlXetS7rGW28wANDwqOHjVhz3QHWwIT
jCZmYdDICfq8BqoF9ZHzoBcOzih2MgUj7jcwrIHK/KzPLqdCwpln3CvrBH4hWiyU
9FNF9P62Ya6XXC5yKecrzrwRzIJ+pPkEre5URftWA1h6OenaJ0gZYmYMsSnuwt8V
CTxFv7NO0Gzj9r15IA1Bskg51kWVTHEGdU8s+XK3VogOZGslYJtk/3ZQ822OyoGn
cxJFmDqQhG4wqkaTiDABOop/K1mDubN2F8Bcfz0644e+dIL7y7d7n21svSIWH5Jd
/lTsBfpg4AmGKN655V1Hn4IzfDXWo9Zie10HIjCOfvX7/b3n43SlYQL8alQdQAdy
32IwaBaJwh9oRsvUhoIkiUagUuQHgTwBsx8StTxZzQRIaKU8tTvg9Zvn6sJBJqER
ZVIO7E6JdHgstbeZ/+c5Zx+TzeLwJjn+VY5aRzdBIaBExMpp9hufsN+IWaZOy4Eh
ayxCGj3KsEnndx8oU9gtBYsoIe/iz+V7BylaOw0i52KG4hUFYdgzwUcrGxc/4IZI
JErEBs8OuflxuQmZtiUfLLysp7qw28uzxv8E4uELoyouZudJ5SgMXOqzfIoSg7Jg
4RznTMAnD7kKwdqvNiqMQFxDPZ1d5Wr+LeYd0dLyv8cRE78rLkhIwH8P4G/Ys0vo
F8pKhq4YZY6rok4I3iDF9qtXuX4cuqF4L6eKKbfyS1KaXVLaw9htv/c/BokjcOUA
uMEQQk/p/oEEeI/j98ZDcUkU/9XFT0r4yFEhun0GeJNqSbdrX5Nv/ih1iwXb8I/R
Uf6W3khyocBZuT1xoPMaYdWE7SdSwOSBprwpb9bX0Vw6xae0ksLMxXFltBArWOhw
iniiU/daZxvZWfyV4ukdM23/ABuPPczD9yJgvlgUgalMsA2fdLHvzE7GeI0vRARs
pQrNTBg/xUMhqJaxCOF9T59ebgEPhG8bYuVWvIjsV0rrZLF5DTSTyQdLDhTJbWNn
/g7cG8b5JzUaomX5/dOPf6r+2LhiFMdwgiKwFnnCNQhVeturEIA8ft+3OEHgbZ25
2UzNZfhZqiM6AAl3JSCAbguUQKjs4dazz3eREOyuh7CMHpy119FmKWedUPzP0RzI
mOqBcWtIBry6MCe6gjJY+HpY8oWOjnZs4gVjt1XkmyQHFN2q/gnvlHNzyEhQa9dO
zzghfGeYPhWE/td7anlIj+nIkZ+EUY/YzOUNcCBK/0GuU5tusGJYruK0YkRhHaYj
7FUkHy0o7lpdDICi03UwvmV+g8WllzZTC+yWWcNHmHkQkh90SWMb8JZu/W02xP2u
ksy80b3JQO0GAa2mNthM6refvjYBYHay68kS/hPfhfSXifE4Zy9m0yb/uT5jK5Om
tgelNgVmBLoEBPmjdzPHlvpD1BME4LDcyPPVOBd6B1L334+eba67dl8B0ZjuscJ6
u8m3Y2j/aeIYDGKfvLlchiITatMgus611076yoUHjNY4W8xOoxnQ5Dt2bLChNJlg
/fQjbc8/YSM2yH1OyVESLXsQc5Z8Fvle6/nKLkkZdqByJNZZeP2RRs21lvf+ZQXa
POs/x/BNUHIRwsLlJG0daRKTZXvyQsQDY+oY2LeWSYGsF3c08T/gO9nAE58x1gVT
naJMOWKlDCAM0R+nvNVvld1AunMzSjXMckAy6hlZLgUq6NCrLy1YQGxRwUPwibBm
BkObsR+XOGFnk5pi8y7L/xi5cBZqsT8sQnN8OPoU5p2k/mVs4RyO58NK+penrbDP
kGehTGnAhItjBsSsaBbPhHISbT5pKRwJ4Y1quP1wSPG5/EevLalIWbhmltDmtJL0
d7dWxMgfqah+zSXBiaWX7+vqe6S4lh4sSvvl1w8/YukA2N9sgreo9eC4Pg5Fnuxt
QbxWGsCqwKb+kxqxyYb9HaaCX5Rjq1IOGPF70YgnE/i9uEiz2MYgFY75xzACyiOr
O18M+ACBXIyiBviedwfwW7TQ8+kJvbeclxiFzCaIB9RMFZ29n3ZYoRr6ZRqFjE+f
HAthgJJ3Vs287YNktMhVddBQ07dnHetXCXtiakWLQRaFwTL5YsNK/07BeYKSkoV6
Ixq7VDnMHnUqGse3dUv2y8Oe3kUXNdO+YrnTdtYnJE5FweIT2qlXjrOmMUZByQVx
L5UI7+MPWrb5Kv+76Pv/nmveDjkS1yylIBLCAZbE8w1c0kgFMNWT6myg6jJcnVOf
ff85GnnEPm9IW2stbGr8QPRjaRK2INvsuvE9YajLsYtaw5vqYgjN5i3r2hKC5s0A
aEOTZh1g7yLRl7oUWNFm9KgumyNWWEkzHdXem+wUDZ+fQe9YQH5gAQb0n5OjeN61
Mukcz58i6/TxfpOG0H3kfhZXl60tsbJusgc1hoaQtQmECcja4n14KUARmjf0xLfr
ZJMnnz0gD75fnjmbbKneCxuoRfJn1e0bUf1oLqMssTVmuV1bKaP0D063XZyZ3c6i
CFM3SdESBpLWYkVOr3BUUg0zP6vovAlMnhtXz6vLFIZrbME0WBJVODNNaIrWrJG1
EvaeVUTcD3zf7cXA0vulaMS7j/HcmLvBCVYcGJhV54TM9NfYF3Utu0NrS77wGS3/
PsPnDW6XmAZ53XdgVpJU7hzXCjg+rQkX064TaA3rl1Zf+9lMV3nZhDlUjTfc594u
rtQE1VJ1/0SZA06gzAkLJ0hDtpvHBNsVPplfto1lpJHeRhxX1Ps50dT97d/g5woa
VJze75ATrygW12BX9BgHPxO0ajLiRe2E+QvA1qnEH0C7SiqjX8tPrRqiTqIqnpoB
RXm915u6nMnVIlas5ohKTnGsq7Ft3THPATnBZbQl1ub5MgL7Vr/mwkIRl3Fmfks/
9CLyVHSfVGpzje0/xFVuaqCHnMH4n1eK72VcLERlCobIqxXA/8e1tJVpf1EyDBdz
j0+SUc5peOSA7PI20z9Q21pckFpuFtTQ+9sv8nC+NIvs6FuAvT9rZq+tVDk4nYS5
6s24qwCE2HAVrpResyRqnOKmMp+fHM1N847rEenQRN4qStq5cwbeYc7WvauF0O/F
JddphK2TlMT0fcpIlOH1ba4+Dip7gkSvx5/MgY9IrwlU3kh3zpnK0K14guLPE2n4
zGUpyRwO1PWvLNIDeC057z5rth7YzFXjASxRLmOaugRQWuBs3cDdCBJjfZRfKU/M
mL/0D2VLUTYggkG7PAkUt+LuKP7pxa6YJ/9r9ldg4rHIFHFm8svZekG7mt3DtwRX
CPy0ht1IQI9V9xi6PFDciKSUptWi/Uhhndw41qxxj4kubvobDhLG1c0qiZm58EUG
vvs/x4JuvV4/PHmRRWWb8MPriyfWKpEmW4JYqMJoeo9N40iIxJ253Fl6wZtr9Zbs
07C96TULoLHNQXmbjvk/QikyeW34HNpB+Sx7tjkEg8UY/Fx/Cgjly3dCMFshPlH4
J55DZO93lPvhN0u/Lfc7yRO3eCNNZtgnsTu4QPA0w5kTYNkNPfKJ9CFxBd46yz39
+7JI8Va0n7MtY6ZGXv98HHoNXpJbanzM3THkRKZjrOsLIqskbrtw9WwRauoVdS0H
DsTvob5QRygy1+n3V6LKPlwnAVPlAmM4hzsgJQsnao7KMMAdFYl7gNxVZC+1B5ls
g65RuzMEcS6IcMmeEioMyIS21OPPrfy1PI+ksuVtedXI577yyFL7xC7vFxtd70OA
LUJGp99KmEtSadxWqLv77lbJxm9qGu7rqS/0MTxQ++cyynuY+aYQaFCs4/hAjTUe
CstLHITP5LZikJEuw+0sg4djlNF2Vbyk63jYvKHzV+FLgMKmx3oEEOe4YleuE2Xa
/mMgyGvThTs/f8viWNqcBZGUHmCRI/X57uFVvCIKLECHyZ5bEg7Gq6OSSZAdbDlV
yZGvllkz7Wv6TBTPlgQZ//ogK23U1VhSjPEujmU63ZcMu3dWcMTi4l7Jrn/Qe+gt
3M4pYzvK6ZF/MHu5dTu7/mNj1hZNNpebxhXjRLaMzPzNEsF07JT7YYXhIkjafZzE
XkBE7pNjJ43gcJsR3TN+s9kSLhhhvSfXpJ7Zu3M57nci6CTEhwZDmUYGFlvwzDdS
rPQP4Lb85wypdShsOI7qcu/LV1rDbPx9Yfn8367+GjO4L6zeDZmm7gysTRoWs+fV
5h/SWzSvk199cjUGqgAFq+0QmORhSdopDb3MC5RabmL59dq1JAyEeBS+U5eUqgAW
9z0u+Tg/uo7UVEIIJ5SsEDGIMffBCri24b1l5SaYq4vOrYccGsRMzO2IbBKEoEq7
PXnKLtMDHF0errXezO942OCKiTAdf2dn1gjUpFd+EiVOQMcSgfWjhJmKugqRVyow
dFxngqsMOkff0KqPz5wJCFMvubzhEZCEFxicKK+P4NeBN7tmULKbiOXgWBz/Jmon
rrYaOybwU8HrX49eaRcqEwLFbE1AZykI0Z6JXfXbF4AyMrKqjX0kKcM6TphqSi32
lSB1pAf5ljlTQRkjddiNU/ZHsgNBs3RzJ9nLkjRV0kmMTyWa+GhmPs/Sq8Mi1Bbc
aeOgcZYV3A9ZxyjFLjRtJlVnXB4U0JCeS+jyAcSNc2ZqaHrnuPbIaRwRJglPT7MU
Ot0491MD8vY41ULEkKj7KxGdUOJvR5YjZ2MjQ+cz7jo6rynLg71aKxvIuTvUTtgi
9qI99hWN5zDNZJbTj6AX08ZiO0KMXTiOVkg4HGqB3SlGiVOSclZI0wevDIjt7ma7
opAwbKPKVTKQGfT07Y5Yb5RbIjHOlg/xcin1DwsMq5zen8VYhkBzh8ymZU2rKwP0
BSiCWYaQzM1n2eHR5CiNEDxjjakE7dNIrK3KuDvTaH8Z8I8t6f7xQancnDoKwWuq
w7e9sG7em1rDWOcthdo6RiuEY1CmpLcB2OevItKgcasWmXLCQjGSns/6q8zTcdhP
UgDXkTuahQYmNpN+v62dn3ts33JWk/q4CJ9Nsl6k6EAUvtF5LpOtkUQP/XNwVnwz
J0UnSGp/WiiHVJBrJmnIf8a0VUCp0zezK9HFlfpODg9Bhl92cOL7f8Pm06LYufRO
gfcZoadme/t7QR8q8O/VAMkTooJfWsylbLeAU1pAgEGE0awCDvu6CBIjcSIhoKKC
WgPUUMQxSRRJ/684g3KMIx/dXoKS2M78pUbKe3sVM+8szLeWAnHRqPtN6qvglB8S
2OJRB+ubrORDxND3RQhDBrIJEDBB3jlxuISqlYWP6SgrwC0nZL56fDqWSS/ZJgNb
GO2S9ouvHC3SAuE8mf4YTAxqU+gbytwd2/WkYiiMFnCkWsVMBDZ+RlaSdP8fjU9g
tKGqB3nueCos1755Ewh3stjaNevv1ho2y+3TekpmGOXR8xOo2VOQpEenoY2CcPOE
GB//puOyX0edlGNw9ArG/c3SHjXRwoPnxZoMOI655XT0ZLM6je09LRezFCfr3pJx
jpMaswVcFXP4CkIVIJFe5eQC6vyBQEXK7S2wJYxdvC55K+B6sHWHzbtFxwqYxGIa
aO1HjNCQTqKuHxRWIZFtvcCEqiuuiJQ5+ywZLxcOStWfm11I2+bUGWqUfKm2lYcB
DhGjZ2QOWfhoVLBeL1MVQvXJXOlZCNGLdsoq6ccGfsDhEX4DmEdHdaLpm4AIw9Fk
aE0TbZ+ZySx2NtoRx/KLRZlJFSF2ssP7uf2dij/qO4jbB7t/ypJ50dCH3tutI9At
AdYvCFaixBuTaC8fcoEUt5HI6UIHvbRl836y39R+oGGDt5P4WvoUPLBgCgKPBbjO
1PfGRz3ix6WWpmC4TeqfLXmsocWMKo5px62FGUSKqqWh1Sf9tr1q/OjZTOTLCUoP
BrVKkzkts7NawjPBEbfdSABknEz1M6vKZz+6rGBTREBqKIA9OJ70MVy2N9sULVq4
q9YFj9DWsAR87xJwv9OZlBpiBoWLgCDJQiVozmKP+TVeXyxtB/emds+MUUytCO+g
FZYu2wNym/4DQo7dridj3nNuPtWSBgqaqBMukGGugHoxii0mqbProm4sMeNXNcS6
yHeOa4WkdAPLbXkoO5egqsgu5qzJMtrPQVAiSF8N82VfI5SjZCdcVG2taJmMkwoO
S+PDgCFhXCQAF+lYZ9g4gWVkKZVY05p+NSJwv0iTjOwVXuaMWEMKRWJW5bY3UbLl
kYt744I6UuhX7h+Aeqnes3WIIe894EOElprZcLDKAnY9G4O7FCMJXXXPgxq60ar0
blc1WpLeIPIcOhOOOEbQy/0TyR4uOb//E3CjUlFC15/WjlXdYp7ffTDF/A0EjBeH
LkcocnGL2rPVWqBd8+g5q09UEWk71vD3mvJ3loAhew5hHSV4w8+jLthvcnJpkWKO
50ki1OCiwJIzC2OYtOesBazu66oSRk0YxeIPuUwj5zFLzerCUZxXaoHuJUC+qmZF
9UzahEabpfNpcBRByk8y3NAjf5k4LYWgrsd7szuv6MKRY2DjhX23X6XBqcqeq3Mo
VikwVu0TvWb5ayIzSKWHQJaNdv+3US3tYc3sLNtMJgt9xDMbRAP0PjtA/MCBzmyw
d1l3jXKNd9Jv7wwfRaYEfTqtXIOrJhrU9opnnUUMDrKbpbVT4G+BJAcwKXzRrHXm
zD/c2EcLdEVzd3xZkE0q/hCDM0Jbekgz6a5PBPHBwAQss4Go6e5NTValK2zzRzT2
fZlRTx7cAnNfynUEbjoDfz/htH7ta0D2w/g5lq81ajC2hr4S9LTEu7KgbXTaRGTP
/GBX4f+9cMFkjPgVr7d/brp/krc0X8eXmrNA3+B+FDG6bK28KIz8UhxU9Cur6IKk
xUPZpiXKJaho0otZqtecdIb1ZLaSRPp42BsdyMrX0RHFGGK5kf25hDlBEhK+Ic4G
aMYhXqng+puhlTn9/ltgPlFbrfHuXSlcp+KjVLlBjIACq5CW/qY1EHkQ/n3BbTIZ
zO290bxAHR/vHq8zeMErTGRWGHAinWslSc2R4dJ9DUt1GOLql8nX/rnVN/TM+S1H
xkq9m6k5tbSmeWwTL5453IIYvjO1Zx0zZ38akxUwsnTPztBX3Jrtre4nE3cXGSmL
6eShJCwHv177gukuPB3X7EitJS/ZOMjnBlLRBALBakE6Z02tkxEGf+HZbpnC9eGh
RWO0DZqT9/Q0sH8vLNz5D444crKnCVHrrQHFIOvwA6SlYALBYWL0XKXLHi5XIfkX
UGqrwanW86KDnzMBuLXDmzjsmRq2GOP4uIQ5hTvkwm+4Y5rYv/2IRribUp6KQihV
slR5rdmw97GNIz+xSNxfbfpicKCtqX4D48m7Jg+ULckp5O53nRIwNCQrwK5eAlcu
bT7x5OnOSjHCOfkr4N/iOkWaY5tdTrsRlPa6pHRl88tNlDw+aWUWso9XK5u4yKb+
KTTlyJ2b7fWBoP7pok8WCIXHF/63XOmHJr+VO6n5e3MCHqCI+FlurgFu59Ry2Wfv
pTDBt84l+qXYf1VmdOWNh3mXfYnjR8bW3YFevwocP2+9943S1drvnBVcVDqCh5eU
HlEfifcQvpeoAVgrscdEMHDH0U90IahxrtWm5eZ6Vss8YUqXpJNkjeE42Wv79DFy
KTPvCwzejO6vOZJwfIUwLzZVkN63Q8fXqQ+WW7ZmMNJ5+MvrIr3EeMB7VqGyoUyo
i4W9hY9THmP5bSxlqJudnrcDV7EPFC1pFxRtwKaSWTkWx1vFmgWhjztp1uZM0T5R
o/8hRDBSVYhqgxawgp8kBOgIYn+D5oI1kKv5/wynFMlP4w4BheB41p6/Y7T1foVZ
XjTKcwzwr8q85M4JJJfqHiK8H+1gEBO704KA2yRQaFA/0hDVqINjj9/+FkxSdf0I
vsIrXvjB7WYUNpbXFJ0yN58jPd7ftxyZSj4ulQuuFvPjPFWuLpYVY7Sym82PH/RB
GmivZUOmQAm0jUnnih4678R7Nf08YuasFCcW+0VdCWZNpZwuWu4SVgBMdNln2Jrs
tJElPopAok/wvao+ljUV6pUx2gpaod81TBwT14RHRp4pWRbqc/4nm4Eo0RZ4NGgf
ddxA/85aFw+SatQvE8vaCntNv+R/HrZyE4+MMz/OLtg8Ds3NcAtcnkgCCuvtIkBQ
YScFc0z/YLkjcOEtstfhWph35l22bCTOAv5fJIevRIQYSYegwI8JRDSE5a3jzLpU
yaaB6BI+4+G9r1AR+sTLn78ZmBkNlzZhBi+i92cAd/mQFCiRgv+CybOXMaXe1qln
bTDUb+tQC2FCgYWrpyhyGCTVBgA/E13m7olRm4kHs/y3WKTEbHfbHOjbhIJ6p+iV
WtcVU1E/uaw3m3BJds9xYIeHPO3x80/iTv29xsGid5qn2BccRLJP0BAeq4ySlzjg
MXrhI6ktEFKOY+dZE3RzKAUjTYdYeqH5D8n9iYzWgEtMlTeABkWYf70+eCTvERJ+
ob+Tl7HcpTLu+6CgD0fls9sD3N15m8NdndRTrdqlgds+469QCPxtluLPN3O1i42d
ogGRKhSaHBvsUh1n17Y0Q9AZBQ3lSeEBfw56LAuFwb8p/BGQ+z0jUSwcg3ZLfTRk
Keivia6WhgTyqfVpiCYmkIQqQ/BEDDozw4AcCM1a1vnt3T8K2psMbKz1BcZ4ZJVr
LxS/I+iwpF9GtUKZK50Pj/AgXGFjv/xE5JTpVSkmk1+skDk2TdcwFyTNJWr+h9Ls
SIEe+6ljbvoL/HKHGqCY64DG+IAM3JkZmmbwJLOaCxUTkxyvqHqw8w8OQUXDk88x
Va6KI3Vcaj992Ve4InqgAIVcL2tgGvIEA4LWuYaW2YU5+dXtXYy+/x1O3ZFIYdUo
6vx/z03tfgcOoiy4h6JL2G3LLEzG+U4Hrsikn1grgWo2asO9BRjG2WeJ2bPPS1QB
o9aeHW54IqJ4zjsOmCiif9OaN3scUhweK+OwiCEHFLLzzeqPb4YgW2fU8SvNktU6
XrQvad72SSgRiPwpO6TD0VgkJtMKaEJs6m4A8fIbmpGhZZApKn7BZX/2eYWtUqnK
U3knLu9WEyHiq0i2jX7L4d6dBJdtsZ9fyn3F+zARBNR5TokJHNaVIQZLcEKo5ifx
14Z68Yc0JuGZWFBh5bCHpm0ib5Akb3jpyPQUbmBCJ2CPMcQmvEVbQMF7wD5HTTwM
9Kc8SZaJ0GxvCkgLUcNqJEpiEdW2PVL/6yJ7Y6ebT/uiZ648SXUzkhoYeInqmk7z
zFaw8dpP+SZsn7F42p388+zZwCzhvF/PB0WBOrzhj05uWIT+W36ibbmi2kaiWaHY
gbqu0AcCL6BFlrqeh6iHARKor3rs5lHISx+51IiCp/bZFqdQC7Yh/4Zz9AyvCqC2
NYcMiTFsyasZneflSYwi/0aQCemdyxrlZ4P1+vY9ju8XqLLWyqLP0/hJTCPZINR7
ylUErjO03aCTAhEt7FSz4YXDEAh79FiCk1baUFlplLTt06dWclmZu00oG5qmCdJe
HBFqb4/EpoDiTyEgqyeHS3y5stltmSUbl+7Rr9V57H5Gz6NB9xmd2sKgDUiopu8m
/4gopdh/LU+N84WOFXUh57cTYOtx4jzWkuIJnO+8Px1f5oo8/jzlX0risoRlWtvr
QljsLkKXkEwcNGng0P9Vhezl74/kttG2uLhtEGXERI33QpgBYFpXSuIy7kvwWQ2e
n6oPx1/f42MfDgtIh1ULetWkfv1lZcRpvvepZ7z3ULTvtiBIHpEkD6Mzef/sGx+n
5vLluj7LJDHrMerI4xsCjHsUeFml5yEc6k/K2gNbIIGZmGiEG3PEMtGUsNCJsdoJ
x10df2dbohNoVaSGzijONi1QmATfEh9C9yITCF8kCxmdEFMl6IOLJkSawhPAJuI6
Y9eNfOryhtfM6yxcqHAObZCWQH/SwYljO6TbpqyIey6viWzdketzTKQv0ev/hM8W
AAYZNVRRZQbmtO9JnrFCyatrRaMOyqpETx+sxui+YGDzEAwDz9Hhc3r+A01yPauH
Y1gkg4B6MopAgj2MreSUsu32vVPwszN57zOlxLBuUINYeDX47M1U5N+M8Mlx59Df
W55NHOs1l5JBg+CNv40a7LRX1ZMYNnfDvYbNTxWzEp8VII2CRKQ8jOlAt22qaI3U
UVoJD0zOOjRTJnDnUszvh+AzZyRbHtoBrUb822xPZKIAb2UI4elM/3zXi5V8smRa
DRd25PSfzNUPgMjfEydB2E63eKu/sfU4QHwnadKYQ+B7QIU9dh+VvMchqcwVUxO6
LaMswnjhl7chVVX/YflCm08Jyb9RpG0toKVfJNt/XmWLuLq0yzhEc1jskcAX2Pk2
zKsfqwf1JHQ2QrBvnKmA/35hATLeLCs2iapQ1UQIqitntBTaxtTx3Gl225EdrPQR
GaqguLUZZUH0sCr6/l6nzAGe4xQ7W4O9PvHKNqxXUiF/GVpIMq5Z2YhcHjDBGZnR
8h1pqKCaVEwemkdxNRM8UQFASVoVNCFXD5INPFKw6duqfoMr9OghJz110x+tHALo
Br2MnPQOqStDojan1CldZgpC8SVNnLBYL9aIAI9sFrMNAhOBiGqWVWvZ5L2/NvjF
J+azhu1CJZYnV6a5h/JFAeEfgw0FXC1JWZZd7s3kaEApoloWN+24aZnl86o7dXaU
4EyDNUG7xlZhFd9LHtnJtETBjYrX/FY6pKUmhL5wLbE00l4+XhX6Qfm4fx971YsU
3Po8f3bVMFzz5K6xCIgTuTbZOFcxM4xuz+YnVvm+wNB4/MtBQ25WdknnBtITd55z
T59yFsk70vY7/dXTTir1kshYnpmOlVz3EusUtWzC/kEWuJYIEBPIUtWgBkdLOBwN
bG6hOiRKC1UMHa+D0M3QtYYCx50xlH65qg1PIXSNTkDNO0itxvcarcIf8HwBlp5r
/3KuUbpPczNocRIMTK/20TEhx0trnd2lpgmEgx7HBGqC0aOWM76wyrbnAaNmNPuo
FLse9Q6XHObZqI9A0CQhbq5a7m17QYmhKHQz2bVz0HVYnFKAukFte4ThjnjckltR
/q4Z+n7jt9wRLscrX2zgbAUFFrMjbgQAgi8HpGCnmuSGMxGCk+9o+I8oO47k+Df6
ycq0ggwcQtRr2VfcbwxBtjpnfqUmq8TB7XIkW+mPn7qi8GPeDdMsc2giZWuGqPWH
N/PB2EYPfaQQCSfn8Grg+OXkulzlIuNzBzRnn2JrIRrJrFrTR6NWPR9AvARzZUaH
kscYbocJvUqdM1R/9N8l8WmeJrVRQRuHUbrCbbHT3fDhUx2j2EzRPgOyL0hNI8aL
GJa8/RF3adZQIsZ666hgvY30GdGDkHqb9VGLMC+qIiQTLnosYiHfd3WSNlODdlv+
yQhEb+u9oFa9xoLsJsJnksfZZ+6jE5MZHuofGz1cXG9uj0wcyz1w26y05LMQFc6+
0EfOOQFHjpAts7dPe0+rTk1ZZ3/v3dh5Ohy+Hl00h6fQtOfgU7mYMSkE50D2G6Mr
Ls2a1n+3SpMKVSw/9oobSTuwZcX8zPd+6umy9WXnNTzQQ7poYoVLYmMceimG1Gag
9kS8dySCTq4lOmzZyrQoxCP9Ym2MvJyRn/8mNbsjLgSh7bL8su4/9PnbQ/Uwvu7o
J4HqkOgK00ZaEH/dXT4xGpU30ziu041Khxj0JB1C9nJtoTnT8fpf0s1iSP1WfYBM
/aVEak9NztRfi3kpKvoNW8jwIwW6Dn7CrqLADy53HkVJwaLLStpIIPw4O9oEtgJm
0+mMw+zWQSo8+VOMhD2CQ3if4Eq+RWedSA2eV70B1WrPqIci+Al/fi45fPH944gn
TTtpVrka0f+qju9NGVIezk0o7X5kM92KyaLfR/resk3eZ7N8+1kj7nbvrOmJ8YJn
Q/zDc6aROXV6q0tw/FxEns/tH4ALlRDWVQo0aQ7PPdsc2MfeGYvSupnRo50Arrbf
BZPY1wlhTN0y3n/W/r4g5SrW6U4smOszUaEmy2mR7G4Jz1kOOtod3Ot4ii7Gejb/
12idOkHmSqAMsq4D0/eXpHlofWrNGRxMlcWKKy7Xa7LMa0x2eMKaEgtu0bvQIi+2
55gOTQZK9iPQnTHF34LoW4y1VE2HddlNjzv7ueiuW0DxDH7Q3ni1ZbKe3kyK0aod
Z+tsytDzvyyy27gKySlrONp9PF8Dri0fAHZzF3HlkjrAB8DrQcdDY3K6O0vTTj3L
CUcJnZ+8Q9+ZNIdX8hGaL/rujn8VgdU1nONDxn6pBPHSowUNx/ZWhRJRpuqAIz0F
p0Hk1248nlsUPJmS7Yrl5fZTXnAj3BofI/t3ihHOVOIqsnI49uN5LWxlClJOqZrf
MdXlhfXLZ6ebN3c1eFkRMG69l1TM7ylJS4JoPjhBsUYOTKADkh5EBkl9gZnN4vOX
SI8018qZd9YMjywPDcH+cA==
`pragma protect end_protected
