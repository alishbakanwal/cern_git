// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:05:28 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
fVb9Ic7fpXpAQSx/v6KaBOvDgFz6j7QYIVlLrnU9ZwTxp/h7t1EcUSa2zZ5BHsKQ
hUqIpOfmxuHlQbp5vktth6kehlfGf8Cyq0ZLJJi49hyjIOCszWf2jbuFilyJHKZx
N0h1hCG7kRafZc0us6Br4W19EvrAFtm8dE4Pg2JVvSI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 36880)
+03sZ6/qYSQpw0VxfIdYJuPTvAihhBjHHS4Oykp/GrQkN2I23yclBifjXK4ODh0G
QufrVu+jdJL0gs64SI6UlJ+Iqy0+CZeMoiKLR5i7Qqsli5qTXmJndkap2JEgiTMm
Ahm2FoHeXMOZCdROll2RuZNAQpOPxvm9SosWZMpBkAUU0aQgRGlSlq0c5XdI0J55
zH4FwBfcw2mZVwb5H9+l7/RcsUDu6QdrxGCtnP1V9IozoWko0SDhYwxANIuM8oTG
H/AXaavxsdxeL/o1gGmAHD0ZBMMAQnLGANfJFSE3FtGvwT96PdgiSkFQeQEHRWAU
ySbtIV2K4jo/V7ZxXmgx6/IBnKDYqCkriH/P4emWE3PtMtyfk7aN9XWJIERngsh1
i7+5o2yT5s7VpNfMgXLh4I9u9NmsJdfZASwIe972DPqGL9YlTE3+rBt3Iig3lNX1
3E7G6/+09c+BEUsrc2yGX2xPtOSzMnqz8RsX0cFBzUrCSuEWK36gNdAPnysNzFuY
cHdYT/iJwrnisSaVLjC5sbSN5IQidOtkpTtih/7ecmQM6K4Ww/WWKf51effn64kP
hJMn09VWsUB9BxLaSFSi5z4QkbgCqts/8rCHa/uPVoSC0sb2d25RSxODg0mDIGdf
T3td6LtuQQ716ykKrenXzxiV0ADg4DZ3v1PietIu3ez5JhtbERDMCMYkBgZvQLXN
TwImMyIgwdXQMrTa01p2bxeF+1garBejaCbCl3IoneqL6hC5tcS+6c3w9A2U++DX
oSzNqM+ikbTdNfmHOyzHk39K0Da6xvbuqOqBD4ddXzlxTGEZ1zRStsqYIH9DwIYf
pQmagLqgpvoNhCneLaJQgSrnOZr8I61w7VReVfmdZz4MTgnuuVTwut0ShV+vWlpv
+8cEF44jVgPj4rKqBgWxcbpb3RYpI89Ht0UNG+F5ZG61lPnErf5AFX2tlCNtFFFb
YVTeSbGGyOmeJb9leFqy7ysek1chHUPeTFJ0o2h+6vEerURfkBWx0ix4lk/Ls3Ag
SakveqZuKJrkzETdetkrseVz4Atd12ESbuT5GGwCBdu0AL203k7835bXmCq6iRcS
6bKMkWnI4Oup24aM5FzPFpwQpufFCmw4psh4MGbFtyaM12bpUJrHgiyQXW50tX+g
pnAJzCm0rfNMWAZ3ROfYDDf03WAHwsfzuI68UiuT0ioGamKhOp7F/hzmbpbOUSNP
9KclkcTcc0cKLEeO9OlwQnU+2b2jkmrxHgqm3EZklG0dwLihuTn5Li53bduiITXG
ECVHRIw+SAZS0iwimNMPWFKzCnWMF+d7GIC4+itf8XpPbvetMa7x/f6Os74PjU8G
fcs0C1EcdykG2SIv9QDwGqeig8raKaOCHmdR6hQQGARm8bwJ6mSJYsk/61yA0BMh
3/NMp+aSCTae1P+S32JZ6Fs61AbNQxLJcQM17zTqUXitDF7ezJ/yWNGzPmBGwaKU
UjR0/G8FAhKG3LV6HggjMVdY+w8DENZzAnxewJbBU+z1gcr7bxG57j9iqouZR1F3
WZp03WD4DTuNuIlDJHU2m7lDYNQFKdq9ue++1OjDclN4NqCWg9VNq9bfwsJqudG6
Y4vN5PIFCChugBcOYuuE7y7y50P25ksuO2AeHq7Jo+7ip8g8eO9XLYY3YXDNqUE9
2oYgxI4krVGa/9p3e9/YX4snomaDD0r+we73MNfD48zs9z3wYvI/bfZKJmapkSDR
E9lk0v8utHmNy0bf7y2sDEASmM1QYiwura5I5W2IP4w0v/BXCqnEaARdwv2S8ydT
iyLOciglNYmDXKkVkYKpEisx7rUokxluiQe8AELPGn7XOKY4LXu6iXnFn1nexawC
cl227ggmw6XgDY5N9N9HNyaPnmjoICYFQ1Tx7aiWdNWo7zkEtQuzI21Aw2Wx/zqH
BBCxHZVvte+f3WEpJDXwgQIrsbXbhQNtwaqNZ5zo1LLTpAj3KJJtEEW4FLItDvN5
rJFBCMfr1Vs9RFgVezDOQxYIM7ADogewioj6Etz0KJtZQIIsKxkWw8pFD6tutzRX
HjvrhPiR5cMdM+aND5XydMle4+t9I/3BOgth6MPDs6uHd/jOaMOIXMGnoEMq5cub
3OI5Lw1lbukS4fWkq2gamFmsl2OwMUoZtE65Oeu1V5KIbBUfPiHh/W1jQswL3YKu
GGBI8Ufg97wleoKuMtok6FYSc2326ynZMws8hrL5rsWlcFYRHmvLYYpBa+f9PvQ/
/gA/7kW1+7bGJiV3gIAdlzEqfrCPkQ4mvVGRALA+jIocxiwLBnpCr9T25aJCoDH3
bgGB+DwL2Xo0KIkTZOJGDrmSEfMQR6m2Q3cb6VGxAN7ZzMy8ETQFDuFLroLoUiMG
TTQ9ehuCjO/SBSXhmgW1PSs9PvqKaP9fulI6/wN520/dhnW5gYzThH1e50MwF+os
pUuj41zjyYOqcWZ5c47puN95B5pFYo63XtYLg/RZTadaY0G0L4JbWUGi6lknbHQP
avGQXu9yIqQkVcTHZQRMZoSBZBV+DN0yVqLjkydOEPh8UUCAGAQ1eisKMnl/IBuh
PBaziG24SdCUdUZKMr3fy+NQxw9FqCqftt3iN6F9rfIrhr6VuKueLNmtOaQSry+5
ejsGXHw9Sc64fIqItx3t0xSXPg3H4GFUhWbTNHJTNlHd5nPOrzUayLmwV+EoV7nR
2xViVTsuVG0QelI1eksTCxd8dp+XZO14zcNRo1Jbm8+v5bK4bEKPeMx01XrG056g
AEmpwhZS4A9Pkvv/e7ryiSymh+UBCyGxHIsRSvAisLO5EY5ZO54v5bGMSCCHY9jp
/JufGALKSqXZWj6D0WxcIdXMkREnzoJ7MctSgqM/hxZPUA7oVyzYI7QV+o5biF3Z
gpvMDJNQlBeL/Z+ATA9C1hfG5uUBmBUcgkpxLKIp5cRg6/rH457wG0GVkJbLfvYb
vjyAcIYBJMcEwDnmbZO/1TWx77jY8E4V5EJ22R3/m12kmBQHhsr711xx5WJQF6sx
3hcSX3ywpMsPFNRSlvU3z6rvCsmRlycuJBUZmbWND4cz24IOKI8tXVnLJvwUGyac
l7VEyCZTeuJV41mfu/60UVzPZljfNJSCfAT/Ij3rmw2lK1y9M1tMU0ugUWf7qcE+
TVYnaexNIomKN1jXmbAB9GczjT5LqjIxY9ZbEelpxloWJZ4yIhJIsFXpIrSg02zz
6qo1nxupcgw8/6pZcjopkA6sDTdCJDRolwHHlyInSbY3OebLYqbwJPEYqswvK2p3
QlqUl+3HrQB1jtJM34e3v0EP89QQGn30yBrujYLJDZ0MBJOk4PSyD4RTmzTj6Mi2
UVvN3Tvz7dh5C+ZrB0cN5+jP9ruskXOdIy7MNJfYSPEG0+Ws0yhykylykZzpyc9L
Ie0NWUa29yxf4z+MNE+SvfL+js+2h7sZ2RM+1UMEwOYfLhvO0/5BCFN3iE8K0nKc
kTcJM7wWzwNubtSYdJwiQKuA60mPXF3gn7XbAzjM5Qeie1DTqVxN/nftd2F8DNb/
loh+BuKCFhY3OB3WShTyW9tsx2DU/mBofHD/simswTU7nGwqmcnwpKoTPjgoKFen
NXhW47Ux6XCOrJOamFNM8ZNsldvmZHp4jM16xCyJCLixpa9wYfvoQG0Lo43OkMCG
JZMEjOaOndyV5aCDcmz3aWq3CvOjWJA84Vw+BwSzjBSRJ+6t0QBK9DSz4f1+vtPZ
JVHQ9ndKZG6LGw18xmJbSqgsMSzd3yDjeJnAO3pW0kbYu6q1W3PHp6LIKNk0ntIK
KUDLJoddmWosSxKTfhYsWDv1sPVdPV4XzK/mrghm7mLV2YeFL3OxPnXewbQ+XFLl
n5MptmHYuj4958ZjYk6Z1+U4iOTk8z0zRJgrXPjAgmIr1z8hXcRwQ8DwImjgxpP6
KwIC+dj5WLymcbcKm3h85O7cNxM7BMIIuvBB7fp8RG1bXBqkjlYh57KNbaen1dYy
kyT8ed2NyC0BGcHrGsTq/8D/G6FCF+sO4iHl3/hk1GKra5yxZtJ+AV/GCjeAUZog
Mpe+LCSnRXr6ZtVokuWTieFutLqCxnUKLEj7tFFzfO+QIN3tUAu5KXkFpOXEA7QF
tsFEd5JoScpNi04Vba/ALyC2LNLnyBiYMPSHaJGfrKRsxT7KcJcx6BT6H6Xwp7yB
NxuEmX683YMZev8Z8nP/WUSYBIs792Fp4Nl8KWYLuZJ1HhuNQHwjyfdZvSFa4nOl
z+185vuaokFsEg0kWJtvLVJr7iV2DBP3kfcYeJAJrrBoWNfdNYAbnMOTf3C5EUZC
b/AbxPmVJfKJU1EwgP+e6vMl6/F8bA63B+k4ZycA6KuUnrH7trB18zB7h9r8pzBe
isp/r1QVSk5njUAIETMjflUAuDSTLAmbqb65f6L3lORZAp5IS5WXNOjbNhU6zYik
EhDXsDDnt4fEZDGRqo3s1GxA3vSxLdJj0ybThX03/rTsPyblNoZPtv3ntqLv8cZx
aU9pNQCju9EQ3dYlFrqT9V1NLOsMiA1h6DOAvd4Y+QU3AU6F9HA/J21Hd9WsF/If
Gm313mrB+YrY/J6z746hycNWitzvD4JU0GmWXml4hjEf8LGps4NcWS1D0VniEnVz
ahTtjzd+9PMyCrx4tl3ZOSBQ5W4S+B4fwcRNcIchnefAgz3UAgCDosSOhOfk0TxX
xtbrc6x5xSvVGwu9MRBMe41NK8XSwKVEoAFToNKRUgZ72QmNKo1Ka1iXIbD5Gbeu
d0VHbSG8J1Xq4cCXIIQ5zZYy/wQcUcvI01c5Glh92oANuolwZyyZEItqxMS9WhEi
yhSYBF0JN5xcT6QJo9jhUqRdv8Ij2a4HXNVwKswCJv7dt5JlR6/Bg6xdA9PhtRlG
y3XcRLI0+JqO44lvlBL4rTADSR9jX6ZWjVbngOq+fH1zjPJvPEQtTFcdRQCbcPPg
VEEOSv9Cnk3eR2x6gk63ymtE5xH9I2E+sW7Hr3N6o6uGUSgCtXdMWRb9nG2Alntx
oPnBcfxCfzaUlfkg9+OhiISo9rf12cJL2pgo46F4h5eWJO6PcqL+Mn12pJTTdML2
BV4YWccn4YwxZZNTl+swPx/5TvqGf4odGSnaV3aJfMR+uy1awis9/7EWF6PTMNVR
dj/jxynbkgKbI4p1nWURZJbFJd0T0I59PgmOXSdEb2FHwwNGqpFlhM4CzMBv2gkE
C7pNjIA+/BHtXdY0gBgpxAh/v7IIHvfSvC2AhozsetsSql4RmxyWhiMbcIYbvQUB
EkBBvKOruX8R4bXAlcindfroMRg/PBilILEnPjxdan9TuoJE74ghE7VMyyNyhl7U
f0srozT/qlSt4FZjjSLak3kC3oTCV5YNur9c43tTHbKHNTpsYxV8tafA6dknmc8o
yBZXODoxv/7sPv9chK2cHcj0vd8sd6j0wA//5nDjW6GBu+H6ct1wLFlWZqqAzRNV
o1zsg/y+LnKtsgWocYFPuwpGS62+ElgsVYcA0GBmqcGr4WNfN4W0aFyZRbRF2KtD
K/QvkltVuhjFHTWr8+tvTBWDjW1pTI9GWrEy9pk8ztePUI8KWjqXzCUKO4VnzJZG
7fHegM4fB7WPUmB8+c24f1KupYIte6UmmDHaMpavAjoMX15OAUDdgGVilR4qdE2w
J7LU8nUMZjW3SX44atPcqef9jhTrsvRExxA32t8js6tHrmOp1aMJ9oUjxntqa4jg
Vjo/5Rm3SWRAaEFP/nRdHvB/Oz3FxWIyrlAjBmeRP8UKGBJNosdmSjFsjDgjbpxE
upSCRBJwW6d01BcKiQ2dY0Iwq7AFIXYaWRTNrZTfIa3pUUsGFZmjhg5WkcIvnFB1
w9HRMv3S62B37YsH9GxpyAjpWvrQciq0X1rSGl52mqgXvqmQMS2+GT/kKffK1ms8
S/j7XjUVCLDwmEBLPzWy/mYyDmIXynsNat0PRkxzLJNp2LQ+veuoj69zRGCyPUw+
fnsro8elY38CFBFsGj5zCZdCw9zk5oIB70iRSboSJMjY8EhJsktib2AHPJAxLsmP
n5cL6iwLQ+c6G1aSdFsyHaQSMlPOVDSwlGkJd6VadPc1pOKEY99f1MqVs9i/6urd
8mrwFPWFumItIXib/BTmTVmAQAq1iZdDa9Tk4sPi4Y5/uagStD6fncKgrjvGfAds
8+D5SyVu1NtuSBshZOFYz4W7sTE0XSpv8uPBLxM+wY2NSbXHew48ei4QEeaoVFw0
zFDudfSE6rNckxWl2OnSGb1E060gYH+39a8Ix8Z0eFbJw+OGHO7KRQifqiHCBPVV
GEqnihCjiyJGPc/zjgiF9xW4t7o9eRuQPZ8bz/+fSKTsQFf/1QwFgMEtfvvEeGci
KLh3rWFj+Kcx7UAVdYIJ3XI23J/KLExKdcDQeZnh2ZLzrZnKmla5X2vAyxaK4QBm
cs1Hzdf6kK/fyjG3IC+rYrVWpebFQVV99Ls3q3o+uESel4lfSyMuzOl/8M4PCRwi
JKh1tDRXHp7IpK7UWEy1NKhE12IYbIzKoRudng8Sxt8ZqlJ38oToE3Bhy/N19nGb
sqKOoiOjjs6yH+eX7ceF6VtAZ8PcStsK60VqEgow4MmYazA0AhrorvR3QyDbgnPG
Cvsjo8CQJXMeSJqlMvPdv2GKFqp72iAHjS3iJtRyFGNGmnphx3zOAuI5CIiyBCUg
1tpXeC+jMtjESVRUJD0KiBk9LLW3BaYbgNnN1RQWEQeCnp9ZUkR0+punJrGn+wYP
qCDf02gCBYL5lmFqDipov1tEJhTCqvISP8lCwpoO+BBeWspdlCSBbjNISR/eMKTw
zl9yKw4qoAgd2oC9F/nH9IS4RtI3Q6qMWlFFLwlLu24AgLS2IrBzvbxqSQOp7jgw
10AwqmrNElzpsFzaPF0sgau/+jcGWwT3L0bL0BFrKcz0yyrQZlACPBS+K4W/PCtf
5wmmSNvIS1IIke3s+m/uO4rqjwv7UNprBEM57YhwRN1sq1q8ECd90m29eI+nySgu
/pdGeAOC7XTfw8Hu+XZMnUBrbqOfbreQeDC1cICxM1ick5YLxUNmruWYPU0JDZ+U
PhTfarqDyxnhOSqppwWm14XTnxWGHZZsoldWXtml5Pwpih4sv+tcCZhGxcSKgD4W
VslTw/llG/Cl4q5WDk/4Yg59cfIE98eRcbnlHGaoZ7wyZoa0IzD3BHcim0ifDuwA
aNTzI1IozUAy5IpqHCm0SY+puDSAtTCWwDePaUsEXj57CUDW4n1BtPCf0Uyq4LqA
IAll225b0zlBNofG3So/fd5msl7GciRx0V4WkgUA1zQLStTsrTocVpxAULYgpMwb
31QKsZtJ7EscyEL7ah4b5p5MRY2l/dKx3wn+Yigjv9EWDLedtE/FLKjaWSz0tA4o
YYTfeqdFfrYTEtflpAiuJsw3jFJgxcJUaeFNsSS+Kc1yYQb7bDWyWMqojMfZfcLR
9A8AqYINe9I2dtPOeHev1SvY6Gipo9Wu4kl4IUY6vGWTEkCeDjDZLz+6uzrJIS+k
Qs00FGq5LgsI9SUC1EelyMlGHpGDhIsahkaJlq/Vhnpvmz5QF9Qv5WCCzy2MhskC
BPA8BRfXVX9wdjScfKUtJWeuqyt8QU13X50b76U2nqYeC10w2Ch4QR85Qj+m9vb6
Yq2KEaESMJQz44kiYtfue1fb7LHpAyx+fA52zd+kPDvMC570HrhF4k6kf8/jQHgE
nmNyhgoFdfd5cxxqPfa+yjP77noiuBorLLvs7EJ09Yo/hREqkkYoYEecsguZ+9Ap
HXBdgk2avO0sNnQ47Vihzd3m3nU5fLaokaNP2nUZuET9o0LwxHYhi37D947suvgG
uPGEDVEf3AFBQE3J+KGlK7npesC0lOKp5S1yaB/KtCG/x9ssvMEYUrhegTZ3osap
WREUYeVpOPFxl7g9PhQF2qYVjKLIybg80ABliPPUnZ17nJU8rcnl/gl23K/kZfKA
LNUTyRRKAGAN9odBURZBuL0yS8OadLpKZB/4Ho+OAgK1bxaA3g/7Cco9qpSm3/+Q
DY3XCtMs+oGJGNxBrhMflZO8AtAsmz1gG48hpmZq1iKsAM5oUgbyB0YMG+InXfUw
/x9OLx+TBUc4J6VKQQIpvmyS95p+Yl76WelVD7ygBFbb1y3mMsFDLgly7vHJMZs3
QJsnNNDVnEa3dVMXkpKYkhjJsZ5F9njXNFi/fdvgV8u3NTlKzmI5T7GUbik56utV
HqF5KhPyNAa0ynjMxFlg5VQmVuhJA55ZWY7G29qGLH4LapHPUuajmfh88jSFOwF5
IDrjwIxmyOX6EFh0403ETyXrBvHFpT4yoB0ruOejnCodAewnm3XMtfwqiR9sgG8D
9HFnQBJkPVMx5ILZEF0wBIqtyS5QMiJM4PWScftUTkWe1wSvTuopIM6GwJJYDOtj
L27X06YXqMVawdJxfOzleYvbwYdx7gHB1SYFPiY92wQh8KE7o1/4sLQH/zLBkUE2
rK7uwDADpS8EML1ODL7tD7/YR1DHDIdzcyypcY6gLyupJOthEHu3WM4TQ1Xkucwt
aetrzyyq0vSRH1ND0vKo71wZPZbmUwmjB954LlZUx5mWtEFoLlPP/JR+D5KFACcY
QwcJmRNQO5JwUM7jB+bWeZSb+JB5++HvreCBDcilB7YxDpa17yt8jUUhWBkCaQfD
xmojWotUbtQUVXKH0pNaElzGqsR0yvxtBN+sRhRFnFSF95XNBiRzdeU2zqe/HNdr
0uEvh1plvucVPCCjBBzWP/oOXr85OyCYtY901BzMrVXsLuwJI9JB+8WWqtgRUi24
pStYsDoh2isyxQcmsKR7aDszN0sOYue/HWt4jDbJUjLUDOMfYsJGcpdi6UiCzxow
Z/v69vMNFb8RudOb8jsvdZcSC2wCLQ2+IM4Ogw2wN2JRJMjazBdi2DFzwcDe1OUm
Po/e0ir//6pOAa3ED0w6vnNVSk/6Cr+RBBTwi/vdoHx+R5Wa5iSg0Bn5EoS/oDYx
bAOC2CrGUQx0WHWBgSYa7advvLIuF+54LhdUoUi7gDHa4DWmNbTqaa8bIdgkenoP
hIUYktH9/PjF5jdFb8qbuFu3iyKd4Sh+fWEDBePSL+Q706QjhR9Eq9fdfSpCmzq3
atBBcKZQaatjk7iTusZU5IM/yWYmyqFsG+5LqVku6kz7o5ybjiagV4EMyRwchBs3
aTI6qJ82CJ8b0zjLnN2uoAYga9SxsUyQ5LerOriREWUgVHp/MBxT2TNxSvwbkRdE
ldhz7iNmcgu1vQFBJfwlv5+4JXoQ+M0hcCZjT9vS3lJSKRqFmiwpkP5IEoouyNvP
xYV4jedvvU6trKPeWpDZ+F4R1HU0tGmjvrKIcM5lngWgryLZaKdoy1p0J3fWMQMS
F5jBiNbIIqD86t1pYJ41k/grR69fJJuYRoUaGWFkTbd3KeOyJMjIIGRrSyMO+kYX
eEpTZ5w2b8t+XIPBKuVlc8GZ/Mrx0HI9bW5qATlpZQd4w7wzcP7zajdlt1Ezeznn
i42Hd7NGow3lnr83NmJagAKhOJjObuhhbD3rYuE4y9va8HZLLDTnoupiMJVpzx1S
WFPcNd4EXCsjjWleH5IpO8oUnSmXBHMgqoj93l9aOJxcSd/oR0v8ONWq+3A3Cg1Y
+b9rqqGuHhvq/kETfbrE4KzjoexLChm5AXcXtJE0cZNsrnV+MYuIqHiX6RgnOw90
P5uvqlf9Qu9xeEy32VX6fslUJEkf8gnMrrlzcBvEVr4rE6oc3eYQ3PAAD0TWZ9pf
0Dn8ds8RUxpnsHoGZcRRyEIfaM5AdvRNdkkhZMUPUY2p1DdIUncIVvdhzTXxjRrZ
eh+NDVBwvpLZ7Khpp9VEgVcvlRRnwVy7LEZm9R/7TVi/l302l0pGSFHID4Ctm7l9
/BOFmZyAxMe2i9M7xmvAFaA/JzfcdPXam+Jn4Ep7x67yCnPXDoSeVMtO8sUq+ErQ
aWi4zbm6p7KYLCDbITIa53kfkQegIC9YqCPf6ejO90Imn988er5nXmLYz0bvJK8Y
whGjtZYMCLxeZkaCEmBYrqF5x7F7DbyuoDszU09WVRGrjYqs3IwFelRVGg0Iqk6L
xosdVTYXWBLg2D9f69b7vdMB/bpO2aGNoR2+29h4g7wjih7MSTXlBEVkJ/x8tGiP
5ZrLUL5wH21hI1IgILXXrcDz0kdmgpjZo5twhO19CGyP0vTlIQdyz5qdlNWj+h6b
nhqhULStJcp1xiPwjHG8Hs6HO7aoqX6xyNXkSaQJCJfuKz0mCAaKndhL9mWWrqPb
bXVMDvVjkRRoPnQTGZIiC3este290bHONMMRpGHozF5s+xDoaWKYnA+XJAoQSWn8
Rp40bC88bXk70vpNBvoCf9VfqCbniQ9ueg442sPahLcUVfaxkgmgaFx0ffEE+flL
WFJGqOu1UV7x+JOKbvGJMYvd8OxrjKyvb5pRIj+R5AR1TstSo5dIwsv88L3rF+2c
8+jOnbyndsowBDtHm9iaa5Mz2jYHjy+Zgtb3t937TBbCGwcU3I7ZTTBTJ2C0BvrM
NGXLvbbvbU8riV1fGrUghx+21NZlb7iaE6my8sTBjkcLy3/BuvpP6ZyRv514fDpY
9jgHHG4MnNv78FB1CVXb935/db91/bPUrZqjA6ye+BQapufq22EGs0w3KzpVObP+
6GZMH9BfirpFuwiWvir6XgrexXnwpLjBaJj4F4237i24PNvL2q9itmrieANQ8Mk+
uf92qC+6RpDrtAF5ehulNKGZLGJdbvBFEBYHcRa6eHbyvOxyWcv/lG3Jd/Si5pWQ
Jfz6H5zOoMzJ26o2yDhl1eglMQybGieV3BzQrS3Q68CrG8Q2XxoVX8aU6PLTXBxW
gfjvXWoznRMstWlfxEc70OvM6N9QSdIIE8gdwdeKwP0HS3UdXBriaHr1pJ+KtKCd
3CJX0Taz1IUJKEW7tMXZTYHc/rmlpOh0IP+HpSmlbWHnHaiIwxcNh9RKW82QUl+p
OLssO6HlbGprt9jPU9sJfFMHKLhw/HgpSO3HlOlrTzXLPK9tVlDc7ghFTawvXskH
Ije5T+vKLABFxgB1SrmqVG7TpVk0tqqDLuf4KH9LOzfA6Qp/J/kNCGb5v9/Xxt7B
p2C/b06Udz0c0sD/Qmy+RXWksjiPeCEaQLUgAL+Zv2IUcnhRwhxNN1zzjwDOAFQT
dL2v6nWuYK2ZYS6J2a+90jQfwnU7cw92rTzboslrPQCEcip5UrfXY6CZsUO404fr
UOKVj7H1lPCL3/3oNl2S1F0sHkYOwAK81UG+9zUvti9yVs8ArYZyddi1zysXwat2
oGGShOyRnzoL/JIcohPSdtYaQZCgUfuMrk/EGRxN0oI+8T2dn/NnE7pdSiAxrw6w
ObG/exQ4YaVMktnpWNR2YwpWtKYR3/Qtba3aWH8S0aBmy7XCDFVRGdFY8hc0V65C
tpLMO2MRtAHCG70Gqci7NcE85ViIwe1CWpT3QTlodqnFm0pY/SGWJjTq9LLVYk3o
9dx5EXGWecLEijRjgSRD7asdFLspzv+rF1lfnRLyxxFQ7hKPpSYaoXj3pXxZIENr
UcyGKWCKBM5njbcwRfdrezqvurTYkyL6HG9zZGfxABzLKaZudJsPB+Ovnhi6iTpR
Qp0VFxA/+11yCJvF4Y25sSCsYbMal1SXTpKNnzlBnm9Qay0N5B3daP4pEOSu0cSs
MaUkWqrUcm97I/NCxePwCKWGpI2cF2DRxLBibtwGsmT/ctpoObpmJkMP8MCn3/jb
gNRSlYIBRenDqe7ARwYSpIgdcHo6SY1yx5Z/HX8jjKATfFraJQnKZVAadnZn1Zsi
ACVNOvw+EgwT1QrlSf1STMiqsoqnpXK0RldW+x3IDP9G3dmufy3MOqu8hU6FydZh
JJHSTL8LcthJGQKYkNOUcv+SrXTYsJkNVlCmUQYS6L/7clNsEnAhX+8vv84g5NZ0
E+mTz5u371exvB+GnKiF2UuBkW8RlRBV9BbLeVJbpZ0K4Od5DGRH2eBCVwr6QLKI
b0bL2jT2N6jv7FRFonAn1xUTwgzIlt/ct5Ok+Bwbo0eE+h/+i0Z453eFO3Z85P+P
0mCjGHiqUcPx999+p2BKMqyIreY3PTIVM7fcK8x2qg58Pvm3HI6ugjFnkfqhX1EY
Q3qBnJ3H3pVgSmRF8Kxv5Wxf5GHJs7q3DFAEcf6KzKh7u2EENDbfQ0joCUrie12R
wDY7yL4/ocjMLNRlWJ+FdR/J+2XkRkLk8jzKwB9tccJnA/55oeKsqDF5rVcai1Ej
lHbmenP3iBCIRtCFDRmljtG21ILQvwBlR+R8P+2bVtHx60HHm+9fbHT0z9hjeqKZ
KSSkR5AK9u9QY149ivF98CsqumXaisGhoH9bfN9gC1eIYU3YozzolAhREKERO/6e
PUQ3uKn381FqFxR0SzHigUvcCLr6vouUjDHICCEYklM4NKxBGe/X6xLdWFAWdK+e
btOQsPNI4Uo4uM/mrQhXsboIi2BJdOC0ipzr/Vzmt5SZpXAEEKGU+u4HFoZbDO+A
CFo7TQKqUEsjTNjt13zio/QtRjXS5k4YBDnI7wqrnyor1yDhPOhIq2WJmZaSVdfT
XFkVsBEAwmhdHaxurE33f7jni2AzDZo7Z3eDsO+0D8bCqsOTmlOZuLcWTb/cKjX7
t6kIGzj8wj9vft7v7Mk+KS9083k6fPPZqx9/44J8OZz4zwtPr1cPKMOy2kuYo/74
OEcInc42tY6MGOeGlKesAAAFaWQzJOFIEyNzcShHpQ/ST0D0z+RURTbJixuHktX+
werx0MaFWNEddFvvBfEb2q94N14PVVE/k1n+gIr6dXn5kn4Doc/D4iSjtVZlQFWx
4527dBmcLjb9NDpZrhpJk76CPM6H0BfMoxwQw5+PJXWbLByJabBuo4/Pyaxt4urp
WkiGybAQR4UKWGEOi2dhWKjH6ZQy78Y9B3EKhZrVfdLLveXvzKei2/cTwfguS+Pq
8K+VzMoykNFdxfz3V+4w1F4go5fF5kY7NLKBPzq8QR/zA4TR5MNGSnUFzMzj5Wbu
kLoccyhPRWCj9O2jRUDDSXGz05ZnFeGx69cgdaqX6+pYlCFMYRIovYfTAFPpW+Vp
3/Z4bgrhUbMbLkCEWVqB9rKvPKODrmWez8TDHVsW+9tRaFVOf/+IWgiM1ZoCCD/Y
+Y/7zLC62YKQky9zUvokk0uhwvzcECDo0woWLN/2cp9fEMLWHFQmONVdbbItVLKY
Tivy8+n9C/qUS22xqvEAVPgpGXGIg43ZPeqiyx2Km6ThcIMVr7MrVOzjzjxBDTOr
bJe2CFpc/15KHt/DmowaSHJKG7TqbHomUweb90uzjS0q/+Ap7lw8DQoNsWjJIwKs
exCeEqvzSFqX7JF5qeJ+MFt4bU5hpKviHqD7nc5cwbDGb4obi6O9LBkZRnIl3Yw8
EPoQTPkBZ1AqBi5m4wGx+nnditHO4nwJi9tTfWNmdJlD77jmPX+By6RH9n9zrhKT
bDwMp6InnztYc2hGiOS1t0sMOe+LgSBK333j1FyMI5J9fQ+5kOsBeL6OxV1NO8QS
QkaR24GNZqTxXoSvK+eEwXB45NYlbTegZH32C5Etq7ywFVUJ0C3ygden6xUW6qP8
4lROtY8FOMaXBrqKCHWzaJyHDbSNOS7ciGqaFd8ARFGh+JTvmM9XESs9JGyAd5Wb
93Qoh6z185YTvKUSS7MwwcEglSGa7p2VH9LUwpyqd3PFuj+OAWXs/vMYEdgzCaef
uOhmfCYzjtVtCMw0J+1MlNKihqZ1D0lKuhwwHflOeK9APqnCKeWCl7KRlIBjPtja
9OkO5FrV1GWxPVsnMna4NL0lxlgHzfzu7PUKe6FaQGm7jGLZsuGgU0VTHNAFhb9o
jEP9zeAIR2jgLuSWlDr3asXRe7F3r6xSSiulFeyL5YdVlCBbjH1t+HuJG0XfYrCL
ubQEcmLWsqIory522Ci8CoqzvB+Z0achvveHkwsrUw+EJV3EnTJCIW5rHICtrMol
oaAH+3YamD1oh35YRizsK0rQvO7YvKlEZvV7siYwNoF2Wl3elWeX+B4ENN55hC7Y
4Y50tkSwKL7RC28UEKBf6ZdCYt5/6FSH19IKM1gARclwhuuOEBLPUuLHW6qn3m3H
65fcCgj1nGgIiFRl8E2B/0V1Elnh0SOlbagh+INS4S9qm4W/sV2R/uj/Z2bOtbgb
C1leqv0PKE5HMjAE3Ks4ONEbDQ4Y8YqzDiexxFmHM0wlEc/y/YFR4/e5zhm+Dwm0
J5DwVRSXcydXrLeCrWxVkI4TLO/IPXmExmoZDnXlCPFwIOcnjvX5W0Ph+xcX8B+r
yo+d9yS/i8np+FSp4+gPU3wiwLov2P89StzCTbo40iAflvEuBBVaeWDVGM1zIgp+
uAvVMooxGI3GJHXDiSuN6/OPErk9ptXOPinav/OYtS8MfvoGL6tDrT++/ZS1vtV5
az/kmHjSYJzffiqRWFkfrppIt/eVpwWx22HboZLY7pIzPdLnCixuoeAgXMsPqEBz
CVecXrmiPjCKGF/eZQk4x6RWBUvqOiJZOWUtYKEnECf0OSrJVAf65SokpiAOJnlE
S6NtQdFyV1nuLk2wLA05ih7cx9aXH+EVrZQHJ81ftBFWxv3ctA3AoJJEnrDaWGAw
62xJL+wo4S66C1dBu6iJOfNU3vZOy9I/15cnJ8Kx6XOBD8zPkIzMm2Y6DnUASraP
DM5YEumfllYh2CUEcaGHy+ojWCXAyT61xLmIvS5P6CvxXHL9DU7an2VeswBnE6bH
aQnfOCDv/ozN1CuFNrph0v3hyy+i3lBM3lxkiUsfR0oipuxqb+ei0rpswCORrRfX
nN4BuBxVubzR6byKejIBHq1iRkljg7jnxiKYY9tBzI98lgLFcfseQZW2evNfhdpd
EWUuNU7Xd5JxMfSRnqHgMCIX6yo8Y94LyYeFDIhWRJ5FK244wQl+W55bxF0y/TVv
3a9QB2492ovmS95UBnJ1S9K+mEdBjLb1wzG+DVxKFRwqxhJ6kAeo6wjaZCT/lYwl
5xnh36wMTwXB1Go6RzJbuQ3Ujow8Ased8z1OdVrZoT0lWnPoNL/AvB1123ugCrM9
KLhL+0EVMBcZIy45yLCvpH6f2VgjwKZh7E0UAF7N4Gk7wHbAiww1v2LNg6iQB7pm
ZmePc4J4y2ntfGUJmkfcHyW1OHXQ3EGpHrnO5w947RHAhomw55sFhMfpFk1lRk8X
WjEO765w2YV39E2Lcb13/MZP4sgaHIj4u24CZd5txEc3Xv/8HUkHxdHXoqOn7CgA
kinCANE8g8rfz0nad4B8bgvxztmCwpejkbvnwq25XsbUABR7lOVfHNKcXcesqe+C
ITpnbk04X1fzXgEghVMsEZu1vELj6d3gytKHKd21LFAw6orvUtehT3Py39qCE6PT
YNx9yBPRIUuLKg0xgGVz1tq2mj69WvBn0dVjUATNZNsTHnsD7Lqj6fRy9V32YPa9
i4RY+EqfdV7xoxV3b4Qkikqep7Fhg3dWdEVIBJ/kUmvynwq1USdHXZ28RVEEPPAa
It9B0wZSQc56uHYs2EhgXgH/rLKIxKI1R9CPWvU+9gOd2E2RgIVQSVYJOkxi3rID
RTnnURAecUh8UqRr4BotZmVZabIkvaO3v7j/M0QBI2983fckH0nAGtZWgXcxnddh
U5Lz3pNfrGQhJi51DI85cHqTAOdgOltrbGZhu6WFt/xg4lrcyQaeUwD7TJT2geAW
uYYDFqDZGS7LH3poe2qzLPOFlLBsNBrBfYgf1H8XFolpYJt0q+169h0nGb917a6j
UzHwo8PDSqLIAYAJ6RZEU6t7AAVyNEZTv7DFvxJNdBEgQBkEcns30LlZMMNx6JBX
nwvsCqvlcJ0RXXexOt6T8VAvfFTgDDIcvYRTkThMUtIE1EZkkEUiteLnHL61foMz
qgnJMf9sd+nXyjdnTJSjY4RMQeWiFhTg/8lxKLYmlzkgZmeXXEIfU80jirBUTGTl
wCfOoqgQsNr+wOP82JbO6/yiX8eof2zvbw6/iBXY9HD62fLfe8J31uWhH/mOnc8k
37GZKHD97KHVDaFMi0/GYVlubMplEbj8sIvQa723/sHZcLYf8DL/D2r8Igjequfk
Xb3fgItepTS5o3+WzgukXyaaTbf+so36JacpdzOgqbm0tHo/T2H66cVFe4WoIR+H
DRA0O+6Xs26wb1XFh6ycmdXBR/bBzhvsX3YjSmaMATPPGu1PPGZlMLTSxiTvbZBU
6RAErnUgSjoUqENo4BoabjSibgErQMBst2T6eQf0Dk0EKUPZE00DZHRRlRbRWYAG
1/+2Ab+qAHvdfputOgBhkqYKICotY7lgAG0yE19xJsVW4GbnDWuJYOw03uea8tsf
G1cZPDLdfW6Ww5DA8wCRswkVwvt5J+oYxdFVJyu/++iI/lHEJDk83AErznDp+fOO
6yUON30oiu2znRFxup5qAJPk2SFZzwd7cYnx1TYI4mZAR2EZrPyaVlCmAThsVXdZ
ssSIqBp2mXCXr4SaEGq8/eFFlOLvMOpUR3hH91RjV7BcCZL953ufiJdX+Dlr+9hS
8cpoIJF6eHrxBGECnZJADr+SYvGdx+2Pl7jlAUll63i6GIuexZvJ8rufiGlRurqJ
gIwcAAMSkWXrNCO13IbWUnwelHrZ/GQwDBqbAPqvuDGqvjvfXJeMwdVOV9Q9pFKA
Wilbgxt/o1aVymekuW+cvUBffSfYDRpzpxIz9KImVp/Ik1yM1yQvOh8s+fJLkYog
/PQWT8Gdb0L6y6vkUfrmCHT9zpRmIXfSS8WE0hN4oJTioQQUqmhs/yUBwMjKpbIV
hgPTk+Y9/uR6m4iIXRfNVnOY4GHFZurvDt+prJzXK88vR80JJzmuMDGLZ4uqF5VR
ZbK6G39G/rnbnIAx3wCxnarm8cox++7dQBvrgfW0IJrkzM7TE3T68IXoipCFoFKr
W1HnvmNT/J0y/p0TahcDBt0Mt0F/whoAf6CUnRtbWKPm2DR4KGhgD2OjbnYc5PKV
EH1KYERsnWrcTNF2wfLWCLg/t6MM2YRc/1X2JAL56Vd52A9SqobKmDKhIZuazoB0
708G1uzxqP6xyJ0DwOa14Ubph8AafQuuKxtcum/WVdQ020LJqrjNHTLgbmn81Fqk
2y3PqKV209//QcQ/Cv7ZdwIvjyP1EWCd6za9h/OPOVNGrUXGj5Rzmsf5bpZ3jEYN
ztr98w7MBWu+c1BUbBQdHbPOR/GrBzumyP+HboCwN8rMEZA05sf+qEiW11unSNwU
kZkr9yEGUcmlzwX0VYV2scnQhAju6ATkrETpSvB/E52oki/tKkqZ5RLKbukY8Vdk
b2NDoNcZYmab4qZ0SVvuF8BXc3vv8cicMInXR4tb33jhQ49OteqyrnjzpwP1zB2n
D4fl7hq0JM9Lam7QEBin5Rs+3srAjQ6dg8cSxH7NGVk6kuVsQKvHMFc0jk1NU9s8
ITcSGqKyiWAhkRUyg27U0WTpuFrI8tTdjEAqAAfxhZ5hNMIdbWbJ0SxUPatl8GjM
PhOj2X3sC5APfpc2DIIABq62NJlNPUNy6QfegA6rkkWrKlro6XpVE5Nt4lknnZUY
YBKayR49oi0ntJYQUr+fzeazak+XDdzxiM1lOSp4YEl9gY92dddr9D4xqDr/g3Dd
fN+0bDZJZHU4ApdwJxK19nh/JG8FRkz+KBd/Cv4RqLb6cO0QDsfXBCa2GOpS1c8I
7rWTj3TOoGBdBsiTPi1c0L8nBQPJnyEJ6ZP9qf6U3GFiOXT+zuBaVjWEzYJDsNO/
HEqB91wpBhcMjl9tnE0AP6ea6wzlIP+VBfVyKqZ+LsgJm3zx9jEI/yrB9oYazAeo
5oPXuU5HpO236nDRWjFsnaNOOs45aoXVbtbygaAi0ZJRlhXDqTtoQRZf4pkotGzQ
vUepDba0zewU/UpwqAdB6ey2dV2NnepFShzqUTrEcWH27+gggeHX0Plz6Ww3Dcwt
7E5UDCK8R7AzT8LmA4L9D+JuxViyZNp74rhHLuNBKGkcyugH1wG94vkx4eiCoo6S
sUshNEicdKf/bVYGRkfiNDMaTv+Btgj/mqct0uPaeluOAogpDut8t4swuj0XGdEI
HvBNXMxNaLVEFWLrFtfXOFoD7WojmsH9Z417IDDeWLanRAydezJRXT1Qj4PP/6Ff
bXOIP7vljNs9KKQgTkUjFH8b8QhrowuPlfbE6hWsHKUgUI29xIJtdIktIxnPCZaz
hPDFSWUO1tKS9mE+F0VS1D2SlZ7PY0K3jSw8LKnmmW2cc+JWu3BRhhZ0M9D/ZcTr
Ytg4Kaa44WMNvi8iC4rcmc/37ObpsRlbynsK+G+n4WJ44Dw/MwsCvw3awv1h7UJT
2taPB7QVOjcvfjHMOe/8c64In7A90cnXLsGbZYUI3jec1noe5eQWmfwfEhEGoluh
w2zJkWyYz/feckTBJx0Qp6+2e0D4YuaIqHQ4WViJot6hCXNw7oXQCaLV3oSfLlrx
OVd+RwiIs9SorxLriqAG2bFhLTDYU1OBCd88TzixW1Gc5cU9hNQSyB7YcuDLOH7I
cM+clc284bnQfznvjz7HhrQOdU+foK9ZEahrZCr+1Ed8xfiDQjSJBGA78WvKunEV
M8f9sDolJ4k841bE0R/zBVbw9s1h44Y4WDv0qXq9onycAfuGIAtOhX/LW4WHyQK9
lvSJUqInXvOc1Cc8WLLMnOk3jiVhl7nNN2h+ciWtLi1D62HdorM3xYVVWrlz1pQf
eW4+hY/3nLWbdIimjiJCHYhfjO54p5NnwixvGdbschl5ppm5d3xZo9SIj/QreilZ
4uS8W2ivJeCnsrOMzpPH5toB3KXw8pTsd+XbDtayj6Y/rkvRPh+9KkqL0lgQgkHA
FApySgHF5WPJhilOuUK9WL364hx0biU6bZn79Z0Ls3YmjmbXt3OjiU4RlPskftfm
nFF0dW5IukolieSXvWgtt1gibHqgxFtV2prIwlv2ObVRYja86OGO4YKp0LpfWMW9
LPE1/oZlSC3tdeWh86XiX4UgomTAAalU9ofQinkTfm+BcoilithX1AuK5DneY7hk
Rv83t+cqjKLRN1dxfkIMErivOLIUJkBhnuFblHmJbeb9wqTc4W2Z7USQsewYhGD2
87a3C7htqMoKz17+v7w0/K3AlSSVBvbj+vlq2fdcsvjdc6HnFbVArbpfeKVqbD9O
mLAE55mQFJGqLY4/owFcxRHWNTXa001d2eGQVzktSDjEf5CVzjdqsR5RXQoZeNy9
wgQ9tGUuAn9m2/IqrPF34NDzx9waicKugHlpJkTzYMbKFR/eZ8gUEGQNvXj4uDlv
NA10WhCLNI/Fl27Pv4Ksks697OBoQAV8S/rBlfvlEe97Ajygblo+zwwUZhrEyA+8
uSYRKRysrBJ6YMq+f1pLlv1gwIR2GWH06BeKWw1zI1Xr8rCWImWbIQnwW1xZZxnC
rg7SOogahOi5ZCP4kxNmH1jRndq/Z+/BCP9aSXYKod271m0igLZGe97Kscbl75WX
vwjpnAZq8bK/kNwkiBZ3ykUjn/nFkKlEKaJWNSRnI4cEfV/urErjv9WkpNB+BMAd
0MT8r61Rm7vsa/1clVoZeZU0dNrTt0GwSiJs9jTscK0qHsRBnvuC0leC8GEjzRDe
ohHzbC2yUyfqO8iRoloCnVw5rGwBRVf7anMGBJ5G7nstBD0XYl+DREnGtbT+vD3Q
eReTDqy1z9qGD0y7GcNRSaevpYkhD26Vx/6bPhAe7+kg+9yIAxOB53omGhqWPpzo
YTvj+OoFBoHgCNwgO8ESMust3j9WVCKZ0vciLyd5pR3WBk46kXH9yl+1fcDFV6J7
oP/V/vPNgW0sd3HO11XEnYJyizP3tQawq6touzydChYjiF6uCATjPi6oGp1nSDBx
avArKvk0ZGRJeQnNyiuJ0Eef5xEfkWpy1oUcfSLk8iUg0OqTOvHXZtx9IPdDMlXR
kbNXGXKM2iea0Mlw/3LY/6cNUcoLyGZadwoS3Wpe6IUqF765V1Pgpi9bKwQRN4Yu
nky5onOR3Pq4St2VyxGHyxIbl9MzQC0L9+UWsBD4lKtbNxBQjKDLzy2hh9QQaNIq
dRe9RTlFjcdXE46qwiLBitXROPeE7Jvh5tHe3WLimVIMwcfTJAtBGSk9dcul5oSj
qAUrpAZ75RFnKa6bmUR1FFyWuXNSXpBeftaHU+Frv/TorWBGteU+IZJqQxCup1Im
FJuIxpdOLqiE7xddK9Vf0gljnwHel3CdzgY6CMQ171406ZBzePa5+OZgBhIx1d+V
OT0JIyAaRTUBy1+U8yuk5iC5wz9U9DKzglHK/zLiSJuDpCMgvrknLFd0guQ9lTvA
1mDNfcrrFZz3/Sezdxyx3cz9Z+LAAqJViS/FTrsQPxPcnch8ixd0G0IlR9qY9AY0
GCf5520+ZwuSpCiFFqn7s5l4RTNw4r6prFYRiMficfz3IdBMuxmVVOCiOuWKMwVb
rnD5BxWeG5/jnSxxYyex61FqlRfOPN4evIheZIs5uadQDJz2nrPHSadujZgQUulw
ZTSu5Pc73fhVCcHYNmRzjVwm9DQI59tx/OJ0OcRCsgF/+7/6XsQ/Uw/380eHO7VN
CCs0Wxb9WhRZjmZudel570Xy6DOAa5h/0Kg5gXCQGGs8k/pVJUYH0ZVNBXRLR+bQ
xtVj1pRF5akswgFbn6a6Vt4+aRd7d8etyYfBZKNdHofLa5P2/9JpYnokWHQO3dPm
DpiAZPh3WlEVv1dlqQfYbrKCO19X8eEOCBO5e3MlhOruuvvUJI8hTDS+m1xdc9Xr
mJL5Kf4RbvQyIkPf9Bylk16bhgp/3AYmyenupOhxZTO4HcFn4BCC09XC7SNP/lFs
uTbKpGeEanPqfIowMtwToQ6tIuTTu/FTplCPiPaGD5Y+icj0GEX27mfwYhWYSlVl
0rvEl7Y/SxhQLCypyPpd6itHrbWNJZSBA/NWd2+Wafq1qlfSxNBtk5QZvrb/lVf6
j6hktYXiHMGkm/W+2J6+6ir1XB5iR0u18IVaJdj/7XoU/SSgP8YfFRNKIqUGcwDa
/V5QUyehXOcJ0PFXLnlvEdtrhhQlWm4XzL5EnMz3qB+LMqUDYuesrqOVEPTewJrL
DcQkjW8RZ3PTARDgSPZW1hvaLaYaLX3A2ZWjuzfggr8Wudbyv+jid3x4LiUkH964
iLE4ACyKGcNOLEkOkFfKysmDdKFnI95gNskjcnVnqeqv3DLW66ycKY+ns788a6MO
p13MFYvDvA1f6m8eR4WJIoI3DnbguKp70tdTdhUN8nmYTO7pUwiUg0DdbeBoDDjv
eQa2Nk6ieNmJJ1Yfg7RnI0RakcUCTE/FOsE6BRoLbzbLVAOYdPXJl0fE7MzpiCZW
67Ob/ACNm+5Eka2isHkVd3vsX7RK0vKKo3/xMxP0svne4V4QcIFjRToLc2rN7iCz
XwE5ndP0cBAuIfj2Jl9TTZ/LJ5RgBx3UPySMZsgywTHid8+vkD2X7I+ix65ZLPvQ
YNERD7c7ObIz1wFtibyp5vw66rpnVV7EX6K46DCcd/bZXJCKv6PGdlvzgBG68R6q
Cg/0QpRhJx3o7YxeDYujE88qBhjGFCbLMIArOTuh13RUbQ5vJWbKv7J69HIMDFNC
HQFoL4hckykk/c1TY510JVAN6UF2GnNZocC6OINgnXs0FLYhO1+mDoihvSv48g4/
tZRLurM6iamgdozK1ThS8nAvaeuZvDMcdt9cdc21eC6KjoZ/BCxwi4SxapgQzl5f
0mSxVfJJxWBGsvegLoZ414d/iUeYbPytBRJ0P66SxPqAA35QN86dCVgp/UMF7Ji/
upIjYaG00Hm3EAgJBzB0z1w9e/A4o8JqA/w0OG7/aPL7Yy5MwTu0LaBVwDFhxTOk
oQN4V8kEfxlgUCGgUHOn1uEA/obgodIMmnZirTop9HtAh7dmsDl8P0AhDZrY4RW7
zcODBfASk8cRBLDMlrmw8d0Qhh7bPgFWn3GD5VdFlvyZ8nHp23OtWSR5ujf9ER7J
5L9luZMH75BJO/j56D+81eKtS5LJYS3AOFd+BoSFcrgQhsX6yBszUj7vrJ5qJOPt
P7KDyIPhXxPwcLtMqfuqZhUAO2CATEc2GbcLOekOGEv1+qLLURDrPXtrmMxzuBBj
qXqHaYs/aPUn7LXldO7qs5fYLhSgy1Rdo9pNPsPDXZ2uLr5HksOuc7S09zQwpzaU
ASSKj5tD9rHHjMn6P5rkyzlLYEr0q7l9Pt2QAIAWWZIWU1hoa0wj/kCXZK0azr1F
IG0xmnlqvgVogF2IPKhdS1650II65l9cd3/LB1XCAmCMMtsIDYria7dpUiK+wGWg
6XUw0yVJUkybQ6vGQOjb3VsRcEUXYQi04EM+Rsc4eeGpfqL7qK2ISQBRaTkCVXqQ
gak80kyWbObeUV97cHS7cNVHadzFcDJOX5tQGZPVLJb4zYpMUOANiKWJY2DQw1sQ
+alE6oHmG6lEj5U98BjWscgQ1I/EYXtPlLpZGapCaNG2AYzQObV1uZxMH13uZs5l
6tIpB8xpQwrP2OGKOGP7OSRhUAXG8AHG0JD6a49CgUWkJScqDVy+Q7AbIq2fDiVh
cCRmca6l0ijG8CwnAfRy0olHyzCk6hvxZbTO2QVW+kLvJuxww1zNVZ5Q/giw+Aou
6A4N27jZpBZDt3iDKUgS7twRwXs5piWwquQJFUWEJKDojorjI0trwZidjBoCRgBq
uCSr5l6dI0/otq72GrZNyoCyn5T+W17IKpp4xXAhIem0ylFVjeExd5Mgh0EKL1lc
Sn9wp6Ed4h9rm0v8jdCyhd9wyqAZZKiCy7WoTbNTDFmkVEf+vMD1oJFJ95YAyH0+
86wD5fNUOveH0JzWgjFrfJdR83POZI8M4NZR5BeRca5kGi42wDLp9Tsm4GgHMZij
RuuG7OKS/VNVrorVe1WubPWC+tNvVjk3k5K7oMPyci8xR5xbagVAvx1e6+E78CTz
KqvrHxACN8Z6FLHzXpYEmgazLNzcomPLfO0wEIQsjjHuVsimNhXPXctOkALqPjms
D9qCQ7ODsAVpzvr/FArdxZ2wh1tU3LaG7K3RjFjrY+Jm1MgdPhsWA4DI3Ik6++nq
7Gsiw9sK9k+bA60mr0yyphAp11z8v/jfhc42KxDTSAnfdwYeNRTUUFx3ZKTVG/Vj
opuYd6STYUp6wsvIznNCwemPRRf96ceFvhQFHsC6PscMXYuv/XbY3xqL6YOhngmW
ZMBbCZcP+Js2M5hkqvhpe/MZIx752N9oMxDNVcg2NdnuWgw8EweHRKeckDgksNnQ
mXQXAQYw1tBkeXzsIe5+BRntk0FLNZdnYUW2pfdc1nXWjcMhjCFKZELQkriRnvqd
hOkDnibR2pj5sAZlq1V/GwDW6dbaLxC20ArrOVkJESbWMblokLYrv1BhRMZ91Odh
8J6/LJHJtoUVo46Ie5p8HlCA7hgrNAA+VSXovih1zLAHLcOciPVg2Q24rVLU6ZND
ng7NF7OV2ux1vSz1glpMv2VNxAoFBcRkzlFB2gfG6G0Z69DuoXZ99MKmJ+PboL43
ACvS7GPOaWcx5uAb7yf3zK7kNlfWVGP7yF67whQMhBSJdPN/9kIv/OKp5CYpFlKM
urm/MyighQSJ0r6CfOCqvUk7drktbqVKVr6q9nq92DFnu2LGCVLEZ5Ckb3PSHQwf
1j4YYmYZo9/CzAu85EhhxxnzJM75UIjU2ugVknPzxTPiZlEF5PNQa3Gdvf++cOHO
xrqxms5l6fhr8Okx8xUtgzZ3ZhP/kKVIZ3AA/supHB5G6vMXZJXodpRmScI2w2Xt
X/MOdK0Chueyvc6ounB3ZfcrvggXleoQyzBVoQRzqoLtfpEEWBAWG+1mVLiXOP9h
0u7Z+Ot8tOrE6FCA2GJatm/vUnSd0fIMOvdLSu4FGAIruxvv1qpkECZqrifZyQcP
ivszMNWypuP1Ua+0ItwP8Fu03DJqApI/PKGUFZ4eSFBEUPJRZpWZrVB7jEen+gZl
jpN9HA7KVwc9KNr9Iq0F7ug+pNxoh18/wdfihea59ekNgYpTeAkUlb+qZAlWxaHY
fPYydbDPYCp72cDLdcAn03iijqkljGWa8ONndzGGg22ynqDyFHe3tLSDmPw2VmlK
C6ed3F68se/IRQEjJEHgJN8x99OuNF7cxvqHwkXYYmWAFJ1ZUBQElNwkITctZ/ea
/d5ChOrt8Ob0On2V8MROB16886k9QF0VkcH3Nft9cpCRqXArv84z86RSwCCl95QV
n6HSEGE2oJQMxoDzpzE3DNDeStxgch4d59XKIaUXXncjf67/4wVoZOnCDE+LJQnx
RdHflqCQ9m2Lyookzt2rHzfXo4qteAevwjKLBbOF6DuDRZvlOH9keMCWDlsmokkY
k1uXYLuB4A2KtccxGvQYENWI55Rqw7YL1PERpD79or87dprwnDSWBLZ3imRc/j6c
IuU27SXxxR7WBEYU+j0WIGjDcsESNIE0L+DU125I/cXPpFE1T37xwgZN4pMkPSMU
FRrqeQNG8ml40tENClPWdxFhEi9M1XKuPqFQ5yIUuxXCRbCDExmzY3MKAYn4mhxL
1vF4W6v8U6tbc/oSa+xg+BwQY0XyYQxXFpSfbc2SjBfoLwBlbb5qYUtpQ0k8DwOr
jpU7mfsGhAA04g3W8GoF2qH8LSiY2/rI9Y1ndFOQ13JtQaqb+KEGIJ215pIIZI0H
DkBJU1Y7IfLMWEvvOsIbaERHteTcORUtpjo6AviW6rhT/LotJOUD4ObSwR1vSwCp
F1VLxTIsDCmQZ1y/QX0E3KA0mxEYQf5mk9+iJ/cPFun8BdjuSl63ZVbITFMwRzt+
+Po4nAX6HfL8p1Wn7jtOki3j6rRCH6b3Dqh7VzJzcJAXbGOAmL88TCrG4PIEwul7
5HEilrUMKu9X/umvzvMTGyxRmPr+fCmTl6GP5VCfTxI+GuXv8z6xUhLQHXVKU5oZ
gsTRhKM2PjNse1bgx1ZoSXrLsIGZrsd2eV8v6BM91F6MdkAnDXNpYfBi5H0kU1pa
Hcf6Lq1ru07i2k60/6blSd4Mmi0Bn++9R56ORhJoUcvS72SUbVlpRtt59CCeroAa
eeVhZLV2skJg77TfTtV1G1gXjqbeQ2N90lx2s3kKBVSDFuiPavzuCsos4UbUA3od
n/eT+9z1uf4q2pEzrUOxwtLbwz0LvVFvx0obxTgEt2SA1D1EcposBdJsfG9kt+Ta
2gF65NZcHCFaNINkSbOpPqRctWe775S0hPNnD2uiFOSxQ8+ZL3kL1j/kwvR2ojv7
Vsqera20zRgAK7yTu2iz99ZND6BO99bouzRzaTd6ZHa6+uvkQdue9md6exsBav6z
5wZtI013y/UqdMGmTnbSNBSs/uDDqH4U1aj7FLpgB8CAfWYc7W2r8v5z8iCL4xYd
2Y0nnNnQ/K56vt20lcdK2l4Tka90IUhPe21DoeS/nZ8yo+t/JfOcgcgRO6zIuNvX
JWuPrmRWf2hLYXlFN3VuJCf9Bohp5k6zakrThuAODjlOmxi605hSqKC7MqUOJRhP
LovtkhRU+vhE42GNIOWZ4E5Ow5RUi9ilJXFeK8NwtgPqSZunj7lYgceRbYTa5CeW
t11JRITeEBIZbArUFx95uGeuW50ynqLytoZZcJYdRbFK6GOPyZqoFK55K0g7KPW4
6ZDUyay8fx3xO0nmVurZniRw+9B3B2MpEX1stGvi/O1JYm+9ZokmKwFqKyMiSk2s
/TRJeaV5HSuJo5itHu2rQGc3pKfOmdltE+zOX/aeOSBOSP0ynIUXMDyJ5SzacOoo
pa2xylJasA+4ZkOumi/89L7cMiHtaKtyghT+R9B/Cx4bhlCzmSrMtOafbYZaQGog
pGUPwlyCv/v3UJ3G5UxzzxPWa77siA/K8lBvqD2RC0a6f7bXxrya0Up/1iI2ALLw
aMDdNe90c4O2Vf2N0gFqj/T/viw9gmN35QAmpHrTqxGqsiRjdgPOthrAkcnovVv5
GnCtmmcYGeb0DEa25x8wZOz2inD/1waSDgEmUv/u4jg7SSzdEdLahz1eY+alTB4u
X7MmENkzlyLOzZAsKXhCdkRBpcSpbuR62z4r52WCBw2kbgjAtMFjHpNdQSeljGZg
TsX1Rsw7XORrPa5FeGHi2CPjf40KyPU58PiqSWSNgbzZFaTG9YqySBSKM6xCiKCH
8eKBw9aW5KJZ8dMDKR0gH0qvwBsJW2BvkRTFzbf8FB5a6R9h9M0G5sJho4JqCvEb
epgs09mexxfYr6VPAJZYIMEnm8UnPuiTl8VpGGaoQadlFruBt2GgAx2kgVua7frk
901lVspCQ3qa6jhj6Z06pRsRpJG8jNCNLaTu+tJ534AsRuxNCewBaOHrysDZ1/ik
bj5rttQkSECF2JfCiCQaXKH4Rg95wuPvSGdZk8fI7sZQ5rBJC/UayP9XZRKlHO0j
xqgTe1Q1jy6V5S4pqo9adGyfAuhzpfrwOUC61tjfzbqlUkKUCbCI8XNVW3dn4SlI
c84KnLCgqtvalrhabYNBNbkCIgcyBBpqiYZeP8MWqNLX4zZfzkQ8lLIWMiW4BmB4
VBzuUm3p9hPIfAodneACEO5FVIM0FtPa7D7R+81sAK7zPETuOQaTtSTQ9yAXACaW
xPPLO01gJJdplPeb0y/eUCjH/2wlop0glUEFjn+KBxuBaH+z+e7gc78w24o/j4nQ
Yf5EqJRGgzLTotdC2zTJJvSevGWu+UOS9f4k4E7Rnjj5dNKsasJaAfxDXLHl1+UX
N2LjhNldiDX9J43mIM0ukfamGFRt1C5JBEXnRlarFy/U9HZkosDnUv6LL33RmkWd
vx2w6dp+qA0jpdGFqBNDtxHutFhJwnPrRpPHjHfL0wXPWf0QTrkgBcMBMhq/4r5E
HY4LGHoO71uCGI+WnRuRVDefVXzRyJUYv3Fn/0u/e/vQUbfrALAEsyQ0YKHGAONA
Zeb3d5JjSrBrReDCL1McbjbDIsSSNohjWtPfQFeYYD7FthnG7AqDop0DdFpLgcYx
gAkNUOHZq8BnoYZxgMPdGkuB9zfNezq0cDWQCa6rTrAAkssAyQkqpnke4OpWiHzy
9S0vtlJ1hMyanjFpeh4PDZZZkR6PVv9L9Ls3diybNfAq5brOStKGM3QlfBnOuh0k
Z+ROnp77w+dyRUeukphzswZKQ+Wpo8CYf8vyPAclSARZe5r67WmIxxkJYb38UIQy
e08eV/kSL/5DDZw+FeWQXphpYis/bbKsbJd1hKNk3BMEYRv9jXaBic44mJgkyjab
CNEwkI6lOqOgdnEpZ0sccWwdWhsScIJncohDTMW+7dWa3Uh5iJBMDZ2cWHpjsq9U
H6O05ELqx5D5ymxoJmnu+gQ6YI7AAnbYGq8CvI1TYQv34Ngp82vBFeDKwkbuxc0T
B2k4BQv7w/3Zsvr1z5cs0bABsu+Gk0rw+dhbS/DY6/b1f4XxMGWQRprmc96/ERsq
su2cYAkL825eAUtaoORujfU53kXmB945OmqSeAr1DzZfJDBQq/BkHwaq8JFIHfqf
82HTrfzbwpx3NbPH2UTZcndjpB+OY5D1ocNKPwM5Q0YHQ8EFrAIDaAJWKjvMSsO4
Na4yn8CCuE1Zxh5QGuGUaaDcu5djWkfe9+aO0krBU8LaZ8nqK0keXKW44xU0z+wy
pYWQgDbRCRtfjNb9+UOwi62w1xSeeYxlXZDHes9OM+i03f+PHmf0ffrI930l61/B
MblVLEOwNBYX8iqlI4ticUirqokA4k3Zqq1lHCqmot7y3jVsox5ES9p4Bl3dIEX6
iBkbFuTneDMfx/nS1SfjM2cYnguwQPwXFnyL1R0SVbvPBBPedvyL3eLVtqKAMDjz
gGkAx0EkbIVSAey9/QBqt2hhohAo/qCjWE9gVqb/pYoqW6AmbzqvonGgZzOxh248
RGdOK47a0vriqSXm5yJNfnT0LdPv0on5aU2e760F88luth/V+qOCXcM/TYO5IRWP
3XB4/fuPvBogBW0DEbbuo1Q5z7XQqoHcd4jnSn6sUZqqkdHzYCbpny+lwnvaYnLv
jbypsJNW3tckeKKm2EhJfdcQlsEXDLnqWqWaaVycVeJrT2KZeJy2Q1vm5/RonKIu
e26jxpkBY/m1J46y8L/ZEnTRrSZSEW/9i+3jRWHqB/8TA9bbskiJdH98sCBc+S9z
k32Zg7xo/0KgPFVoDhiX1GTkpueRIWX2LZVhErJjQXNB0zV88SebV4qX+q9DowC7
dZb7APVpcLyYVtVEsRTOtabiMazbHNld06a19YfgLTt/VzaTbyy86k3KviX+TNah
+5WX8ErwIBjpqJnXhSwMVPY35kLRDtTIVMxOiXj85AnwKbeUBZ0kPR8Q1cM+Hnmq
nbIz7Z3RLXINCG/t3Xk2TOUvy6ZIuSsQrEMMy3mC1JAJYh4kwZwZ6uFoKZPuG/4w
iNNo0/D3L3SL5o8Gb7Len+MZgcAmKC6ljr5HRahrmgk0qxuVjsuFzdKeKyrvLCgK
FWVVrZ4Rf0HB5RPFjcN8Pa0CXfGgYEhSj8LZvivPAyRXqDk7gYugOOss0Crkox8n
CXwJuo+zZf66m6nq+rdbhFw+MzmBs7dDSCYyRbfdCrs6NsKXHvuQ7zJZbtERzRJR
1Qne6vMZu4bfQH7ZuPwOziJLcg9wsdFNMy4S4jmPuhHx8OnRY9gFcX6gay4L8HP9
Sl1P9kGXVoVOJc7Yl7CBKwwwl8XwpeOkqXTOELY2HiMXhyp4BosGr3Zj1wVOr0Vr
BWnCA01WNPMhfh9Twc97HW7iFi9NaasdTVFEg3ko1Yri9ADet9JAt6Ux8nLH5lg3
jttlcj13IjSDWd1+U9XHf4MOiZtqnDvsqEPHPxdDAgvZWmDl1bqGMx5B30x53vJb
PT2MfZJFw2PT/DXvlfVh9pghDCWh4gwZgJ70wZUDWmje6AgzDQbfI33s/VugEIs6
uYIgaskr0HlRez+PjYogx6ko4WgrRQTr9OW8G2lpXRNivcwjWkBPpjt3fZBXVqya
qB58BKnzsUmD0hWmFLs0ae1JIaBTEN46QwWZjZoCirNaZFB0oLXqKkaf1s2hw2K3
zrcQO9233ySaDThYm4bQc5BsXJ9HkH6NjTMpmq4d+ee0RMWCCl29VfjgooAKyCQj
rckh+KAp9/W3Ja5G7HDKwNqllZTSrYSajLQON2G8Vh3JuGPzWhPrsth3D3GJPFfV
iJ4Po2spXZ0yJZM0pmGnTDzuQYKGA7Up79jyTMU+JgT7dinWYmcTVj0SvGVft2tG
gjFvzaduUAiznyppPOGJZcZjKpvKXaohb0AaAcoXf9cu+BqK8hCUR7qlABLuJvsP
N6XYcNYSWOfy8i9C8TFtPSvWlaB/rmutyAUEqmOjzfC7dlU0uosYKvA0S0jhiqmN
zcQWqXiWf2KDuT/03P13T2VfLZaHHws1hFx/goqbhSFnlVrsrABwXmXERunwa6BG
lrruD6ZQHafhiCg7IEBpG8GM6d9xQCP0lMLz0FB6OV2S5H7RI3weMrHDNSHLDb1G
fQh3XdnJb+RjgHZhMLkEcM3XO1r5mSIbYrYi8EDrhifiVuWdZoxUcQfbQE+fDr7f
NU4itTivM33R61oQCI0gy1KCZ8O1rt+Q8425bssAyGsG/A0z1sBC/CjbnBQTMBGn
f5vzIqW0/nVZ+AD0feZPXkUFKtzujQclpfySy5J5lm4qshsAb620JMbLtSqEUtgG
RFKQRLitcA/vMNFmYSvQoXOy9/khVc52GqhTqQI95/epBjZiYSrAyIO1vComHYyC
ohiDsHJzQQElnuPtOUYTjYV0ja21RB2kuJKhwxhlQhwI43fwPTmb9JBxt2v2SiOJ
7360SjfIBaY1EMbhe6WL50TTrsrduXYuff0YwyktMWcZbqbI9VAqt3ViPDWiOVhk
0x0rtFJMj5MvBb+3jr0WtUX8d0vZytppnc7K4VwB9j4R4kHlU2OKxgeLXXONumGr
M7uy+HdPv8D2iM2/s5wJuEfc6EdmRkK4lxxM4LGGi+J9cXp3wkcXZiCBMGuNWfP5
SLtluXYc/CarA3RHVtzT54+JuxnWbUAWM1p4tR2qKdyVm6BmslsetC+VaiCNoPsL
KY0sWXLkGruxGO0l8PQMGhokllLInopln4ydpIvYfm0pB4KWh8OXQosmJ0/dTs8Z
FwsdI6M3AfchQPwMkAXiU+2/uQuM/fcaoKcTiXqT9mGKUhPOtYJTY1nXepFuVUdY
VphmhA3It/gN5FtCsgL/taaLrP8fbl2ctZBTZYAY2S/e0qdc3kbI//9y0qJY8/To
2s5K61ZIlFfYF2ltExF6uV7Ef1Ih8oR2HwL05nqZtiG2vxlcfomPE1vIC18D6Lbi
WeZtE5wf6zlUe7WZ4lbvYcUBlwUKl6Kkzn6pwrEs/b9/bxH0dZUJvlrgy6wLiVf0
6dKVzbMrKA90Qn38vM6ULhNG5VD+jzPWhDATZCAMkRYOG9JxxIHsezl/OOBtpXWu
6l0DLy/5wNnIDujnu2cb60Esds4PUSFGdnF/HblXeo1ZoRPcSFkZHDA538F/irha
UzASQ7iYSp2AUJl7JfnHOMMiEW1oG8UUBY2cHFHzWJawDlu2VSIusFiACV8FWU+8
VHKHtOGkpy6CXtY/V99VticPEZ9wnEvREjfGVwoeC4nzD95I6a9M+AZVytBR26gF
S9FtWY8DPOr3hBVyz6BrKurowb/OoNW2OEmtlBEaAOQm9cBaprdYerOCSBylndWz
xaF0YDO7vsNWdEhmKpqDK0RWBOhqS1FJoYCo6opURP3UagKM3amLSbVqZ96EjJAU
y7Hf65k5dlfj6DgLCWD/r4RrUDUBsfg1DDOJTuquRzE8LtcXeO+zFlXMOYNMsqvZ
6CxbuSK7EG220QuArSUVxD0ygW6YmHVVSuC/OlDp72BHjgACettV8vZmwb4RrcgY
4n4lG2ysQMM/trO6lXSyPfV52AJE3/yGLJyEoiBRdnLUQkc0US34PlA1m6ck4D4v
gX9VP2huP7AYoYt51WdsRkD95Pj2QwV1Idiw2LHQW4oqDhsWz4stbQiw4v3wuT4C
yn0scCi2dBeizx6LWEF9EPX3pgjqh6M6QtITPgiNqvUJrXZOti4CQTmFp5NJmbdG
KoJZu4F+zDaSHGPmnp9NVS/qQxCw+ovAz/4yzB8LPwxflu9i3EROutYhqdQrC4U8
hcb3Ojieea/BClwbIeJUESKqMbYP3GJbMkim2EXSgwedJxoI0rrqdAo5AgIGlb+p
R+tWdmeHWi6Ei8oykS92/Od5vW95gc7HDv8EYv1smvmPftEfhjBnEKLTJxhmSKEi
aRQOtWKnuRf0ypppEFlPjzm8yyF7qa+EUsVpfTmJPy9pAOICUGBRq2aX8Eb6ZEOn
fEPhEKEUzpE7ueZYZp2MJOEvIR2uiT0awHXdbsSc7D/SZ6CXu1OLkf7+bmBmPHoL
QdtDw4REuJSG+rdogm2tV/kefBrasX+ic8medr79g1BAaPL0cvy6DFftfONsbdRs
nG00EV+qEoWhPQK6hD1Q2SbQ3S9XGzT/a7Woj8Kr+h5AtPbh4hilMmDMcbYKiVCf
Q57p7YfYSc85svnpeprAEm3OYgA5IsAkna+U8tAyW3T/iEDLk7+tMZ7Drq6Jb+xi
5gTcGJ1rxato+yUmlOU7So2BThiB+xz8fIydoBuvNE3sWl1vLM1l8KekYnQwB7D7
Tb51yw41iU3fujQzo9kCzJqjbSFrLK182HPiJmntQlNSYweiCuwclCZr9AmXCSjK
UuqRcl0ED1gi/h+Jc3Bg6PRHkkzqwTrNIoki2fffrPZ0IuQS1TyGyRDk2CXEl3fM
I3Dq1upnG3aHbqmd/3p7WPK0wO0HJ4qTQ2ze7ZgRoFUJ4hu55nbRG5Q8WNO32qee
6+bbaSMKrTjbmoireqCXT0EOEMxGPuzJ50B5K8lj9kFDa9a51jLxdJqdsuLaqM74
Wh1rXF0VM9AycD1x7yDgC/AlcTWNXxaJeA/IQxlq7cwN+u2FPlW+PE0mp4z3Zl21
nC+Og9D1KvkiKl1wOCUDDURsA7u4VvHlrbU/ZUzlPPRr3svDyW1cnq6eV2EdFiwW
Cd+LG5Joj0fBxBtgOeiPJCy/xggb6OaEzfdsBJ9ay/jaMfsIDM99mCamsLzVmxOA
NeUrJHR2POAivqFksGgPj7cvTGNYX2OwYXvu4naGIwxtftW4qZ5pvoq+/KdJqa33
Zk7onUkRzrf37A8XTBZg3DC34/u0Lvn6/RsfI3UQoeDpU87VWQ50671F66TfvpP2
26EdieLQTM5uPJNLvZiGqVeiGsvdqOdizOAqHPYKhIymV13h4RTL6mh+74MAwUtj
MZhWh8U6IsiKTU4H3boSp7knCjU192bH6VRW1uzvpP9/+DM98M+g1NaZxEG8waa2
dE/zKdSuY7rsZEFwm6EEjffgmF21s4j2arvJGGin7HJtrLfljEOwuvS1qwN7L62Z
PaxLfzotGSLr5xzbNaRHxTLD8RFDOK3Tqm1q5Ow5qX3Hu8uFM9RsOeuH/BcksbXs
6hGXqRUPnav5E/d5R1N1bPveVqPPzPls8c95+ufiQtySnhwMQDzjQfrV2BsHeOcp
dC3cAXjtDarQiggvkPZnh8G5JAsme0ew2DIxtJF/NfzZoEloNnl6Oiu824C0gzBr
tPdwkHORg/XDwUS5xIc7//R4xeZpk6sioqkcWn6FfTO2TQLkt6/SNopcoQ9WuZD0
vdAXZo5RWwl8Ftchw+DWlf7KgI18wjH8dZHbkJv9rF9Z31sGU3JQ3cgtAVGBFCIG
Bgi6BMeO9U2ZhupsbaXTKWZ/S+Qx211Ehp1fbNe0hqj4gPaV0RRwu6/WtTBzR131
QaKClHrOYsgVWEyW6gvcKqWJdQg6F9OkYE1fWpX2vFMc0v7/LOxv1Mt1lIJ35BH3
GTyDDT/T8OJ+BTOHGBez343eo5elSo9izBN6/61XmFsTZJIHHXjYPW0UrAPD9Fap
mWj+8EuMhI5dkSWonvjtTknbGPIDkpySqQqrvllpApyJjnJ/fD5MZMqHLFeYOqXE
vrtTPQU4sZJHpUV8SrAB8HcwZQklQyBzMfr46V8rdE0sTRYmeD6q1+0ZXn9XNr3D
rgc+JMiVS/4c1Qx4wrtX3ZpIfa0+brKZB2Ei3/8m27ohvqdNLrcOE6l/C8/2w6tI
+9I/F8jYOR1fV+OL3Sdcn6QDCJtxwmCM5vXqMYr+lv7KW27W6XdX8N97ROoO/5Rx
EYfFgKQTaKS2btHgQVCK4NLZD9i7SHoFIUqYQyNvSjLdLEGmiW2/oG8bhlR5lHci
YjVB3tR8n4V19x9snvwNtcuwt1A27cgRF6JsuVEQ/7eb0V+bkNwmyOG84I37a6x5
9eVVtnUkA0hWlK4cTTMPC5aGntkXtGiJtbWhNVuixLgZ/87Y1J4Wwyboc83gZ30Y
9TI1+ytkoIV4kWt2iCBq3WLB3wqauGUYg9VvcPj+h8bIl3zJtHbMqzNGIVHuZ9pP
v0BQ9uhgoplSmDLUB2WkYHpsIXdW2hhEdrRQZz/TC62TrINN4qpyY0j8UBBOD/zb
yUlrE8SZaDyCgDHIVf9O3jAZg31b5SOrViXN96Zv+Hw1pP1gTWD8j3ZRzEilt40q
uZijcS0YES6aTMtR33v0nKAN8gy4UTLyeT9zIzvg/5p61vBlnWPoSA8JRgu/cf1n
AzjZ/IQX0garSkug/kK0DY0q03z/OOp/XX8hlChfQV8RB61dGo/fS8FDwsLiLASj
Ee1XPwQXftsZIXBpnjwPgmmDKJ4onyOCg7kfOGpK1JjqSgzFtq6XyJLgXf4zkE+Z
fIobF7CT6HQjayqxcjhPp54GG2Qtaco/pD22rr5HGyDOY9FeHtXaJS/IGMAy+yuR
Az2fotymsymcpIXgQ3/mfovS3hqPByKBfiZs36yQBf6NRL7slotCHAKHKrBdvzNm
FQYpre6c56i3U9ZOmX8ZC/OwF2d1BEeeSG4rdQO+z3946xCPrsVz2T7V66U827LV
lxVGd9Ci5TrGwZmrHzRpc4OnVbGak6eIbAQ2sf7yEDgmojZGNWpJ1IWdAH2Yit53
dGpcadlFBB3IT8J6e4Om4xDJrDG1Zmj0lsKCGWqSBMVZOPUC2ogIIkcNIRdj7Uy5
EkDPWu4YK6LqUd5RAUAhgA+ILbliWug3OiYuLyfttEcAJHfJmfr4DfMsOx/cSXev
uIpUG8h1Nkl8o/A4La5atMZ3hcBcTufj4xuMUlCePEF+cO5KdfKruavJTp0r4GAS
7UFQE8zTR+eULpQdCD1ldrgLBUenLihfwg0I//BPK7Q8b3dXVq3vcXfZEA86RYd0
C+f+Z6+WLXt4gkzK9lfyLrkIZ9Dl5EjQ4EH0sKGiJl+IEsriHW1RnQDo3GCYd4cT
1lgDqNCfgnH7D9kLHQ2E1Z8WLhSl9Xi6Nxl4oGFCK8zgijFqbUrchdGUkgyhmNN2
l6QE/yvCJV+b+o/mCFTOk0vw61MAOS+zNiCWo0KfOxzc0NwsfrSZ1hOV8ZgD2z68
qFZwjkP//2BdFDMXpzKJ+IRM8QZ31adip0nEu84puXRPy5T8hLnWQd8Uk1JZZA3I
vNZpuMSm64Hcbz5wSF/jZvCHtTPL0a280AalP63Cfl00VbdlndJjJyaAuR3HQimX
6uZztOr5PJ5J1zGE2grjQ2Q51ach4jXFBkrX98/dhFzNezpwAXatUofJ/lx5hpIP
U4rHrb2vzYslLFOhSjkfNJbFZT2oDYMuaG1YVyYBi9oiVjnjPtIGi9hf2JzoDHzW
sFp/Fce38bq693AP1k+b9JdLEdIhH0whMJBw8CppGn2aVvTNtVKe/BKr0guPaeq7
xCUaiVBfy6uD3JKFUVjdM483tnCQZ3HTbNVUnuDZLGm+CHp0s72DD2YWhopsQ1gZ
ghY0iBIINXL+Qv7TPt0FpKtPpkhXEDHUkEW3H2LAXHV7aERCtHUHWxGDRL6wmCtr
JD6cNHq5BWs3fg55ub79hZstQO/ZFYbt/m9OhXxwOyheQ5Sc2AP+R6vvxaE8O/C2
ZgCLQF4gXJIaTjW9jPBnGOYkEz1JC6Lz801Bq0Qa0ZIjx1M6hPuGfWCWAU3JqJNX
iZ9v9zv53765RJ3hVZ9t7dBg08k6qpy+7WOD0LMHMyUKj84dzNif/sKc2lpktJb5
kbbR/QdWNHPED2HT9nFwtFQvyl39uJEr2fS5ZqGRDaSGrOVYK3VmydOXqZfO5rpz
reanng5cm9ibENSaNYK9FeXRLBidqiAIOc4S+JEOgzPyCmfSrnJodzW3lxX9f2sO
WpnhT6SxNMFNtQdjiOP2gvp3C8Sp88kMqsDjS/bVSNruku2mjzrxtafPI3mrxDHH
79SjqkvS8MASypu1k4n5RSd6GHZnkLmhBnw+09j7mmF66WrweWPSj+bKZ4YcFWz5
fAnhfTW/tAX5AWhJmadMLnxkOPl4t1VhB9ChsTCJhMjtsJx+52vw8p7/WrLMRA6P
t9YDczDpO42/7mORZwblK+88wWtMXor2NxZK4yhKtxIb+Ky/l/lg0yxkTqDAoUzK
uU86LTDMLkjw/Wq17Nfrqxbd5Q662RUbB0QpK6X2NGz1jTU92uWmsADuKH+NxFTd
/DVq3yZy0sxB920eNTLVPUcOIFnHfxRl/Uh9WGPVkGGmU8b1i5rkBiGNgPcJF7GX
lHP2v+jKCoKZzR6SqlDesZOz+V6sFeQq7i9dVGMVmwZFXWHQSzJ61DL3vTsoxTk+
0NDFLfbc404k4gg7GzzPiVt1uSGdCyWvkEX/eGJ+4qFnqhkrJJoqS/eyxBLDwQK5
92w5I4ymXr5n3sHp0CQbg8TKRa5V7g3u1o+jy3K/yrzPRemD+xF3WoTJ8Q1pGPA1
hLdTL/uEapmOTx/+ey6gZJFKwFZI33iy1x4rrbfSqN5zYpGfRlAN7rKTME0q4mRG
X6cIlE1/RMfXYtPbLDSuklEXWzL5Al2FpQ7MaVIVf1kyy6LXIrxLxXrD6Ya0hXEZ
jGN9J7MMnta/7tASWPF7XF6RJWE05GcSCSlk58Jssmknflty4T6bmljCS3xkMBGl
Y/47I1AqQBRsnluY2d+5cEpPeuAI0arqw+dsk9Lna76Ph9REs+r097vThgEqV74L
wo74imC60E4guTDebqW2Z/+2CEo/9BLPMbPpxciOIXWXuJm0iLtyjF16rhZcDaAJ
GoIRbmBNeFQmC3DbHh1hMTr7oEwk6Nu9Smn+OHPjpBKLCL61iGKT2cwGu/nWEepw
9PC4g3yD5wQQ39j/IjFerwTZOhTsyWz5IzH1z5c51eWASiGRafG3h8nZvS11jHDa
bEgXjufrUVm91EmDKP6hwlVnpd8E3t1y6aIWk3gYOWCVdl85GSfq+wwRAtyugUuJ
zn/oYaclYj5JGn+IKDr9BqB1Xf5nldiHhwUp1RTzV5pruipUj4b1V9AKxXDDQnr5
hzrVSy3il7lUKT+FUY01pZvU4NEmuxPBTWbJn1fsdpDMNwys4hLFSH6U7OEaoLtq
bZnKErwSoR0RCIm5nmc7e1rLr9D8yxQGDGuuivjfBRnH6uTs2vsrajpFbMQ1cB/2
U4aH9PXNUNNGi55G7FcAajoKYvF9NTCeoeaks0XbD/5NACkMIv/qqmJssJn2agj3
D7Tbij6di3MxUJEVCgCnVvsewtWy+7AQUL8xHREJzTwR1Ps7YG4HvHOvH7gIaSTA
yXJiJI/S2Q+EcVyicddYMHRq0IpCq9WZs6oz/NWk5Ot4NV1nqs0/zpW9Jj95QqcA
uRy3PTX5oF+ZC+rvODc865H8IOw1Z38AQtMuBKWKVCaAmLm9Dgv3hPUg/hXYZiWU
K0Nwr38qrWQPCfVHVmQMET/pRTeoSQC82VH6Tod7HW8GrtyLQWvmMhJegfow1Q+6
KzO+n2fCt2sLQ7uUhrCayq/xwtlj/ZQvL/7pcqTCJSV3WPj7DyKDs7rZPATFCbBm
Mq55J7b3PmS9cimMqs6FxSMqatcBO56wyFFKVZvJYnwr+4dUo+/YyG+t3z35bYbD
9y/q4n6Uame+IywfToJ+iBb39Qvt4L3jOJchcYpNfofkjQY1KTSpTVAMfv3+Fx1e
qYqGlCSvoMO6r4NM+gWVWkLshj/nGXAPMjkPUfVUC2nSmRPXUOLAm7y1d7xqLhm8
fwJD2ZKi2xcbsv8UOEcDcpMuNnQFGXd4WTAsJpCSoPOyZFqo00821v4BcEISIOBc
bPvKbT9iNdX+yuJgeXmoV3bYpv/Y+9YuDrx130hFtjwRnMf3eFir+HY3FX7GUODu
2cKoida+iEF8Bbp1XIypnNxKaDXPXay34jn5F1icvDqi+YwqIvuiSXWDbQEzSmVD
/I7eVOONCswOyn51Av+/sH8wz+BcOS4H4d9a8jch3AI3RJOGCwdIGyqoH8IKfosz
97rT3IMHHLnsyktK6wdF720hsHHBHu5oqqbcynuuT+IP0lrGuecegdzq2voZqwfJ
4QzQvq+oORbjdyS+tDllSog/abEPzYR2g19+HZhS19kKG4R9bzi8lsh1Ax3ZuwxV
9NoG+We9hiNZemeFBhhalT8q8znyJVEU1lSwIo0NJA1VDkxgSNQE89X+Gxr0lI14
U8y+dnZQy/MpBsoMQMxqra2zUzgFuB1OTyyjOynw0X9nZchV1lm77yxnhLYwipY9
L9benfq+t1hE4v2uGG5OQK2ep6H2Ep7D6oChTV0kW6+SPqk1lO9rx0B6BpRyLx6m
OrTM5APH/Pu61x8FQ4FDLfJIXOMvf/p5c1hedW8eZqZcs7keaj87HbZW8ykAcfiy
UB/TbJ8xnOd/8OdJUSt6pxtO+mrNaOeM0/zENawFEyI3JJCdWaJALSF/VCdsEIrO
w140+BMEzti8br2g0O6Q5U4Uy2IpsKo+FNl9u283xvWjNAA5B60Cl99vlW3/VK38
wulhnOxR1iGW8B7Si0cmrEpr5HoZevUO97hltpKlC8EZNVdDyujGLWgQTAf8oN75
PJF3CzP2ABQ4Ee5kystLkEhTa1RM8/fmGxBjniCq/5OnRzj+RZ1PT60xTwxhqtb7
hcYNv6pzN4p7pfxTscvUFRX2conSaI+RJmM435B2cvZEWPrOtP2RhGn556kAcLdB
9bMLPnekT0odpGEuf0JPaPH7K/sUTFXU6MrRsB6kNxfeLbiF7MU9s+hr8jFlWgvZ
j/a3XmeJGAboPQ3A5kjd68Ua7QvkzmpBPr1RIzCDajxEEh6dhENGBNyEuplzIONJ
Poc0AXLEGNvX7VfHEbMyqD8LFG5znQ7Y+MfC3NKnOCvJ8OLz+vghaIcwFNav66kN
KZctLcRug4iCk4a8ZWEm4aqFmZGL9dD09QhQUN/KpYA90GMVkSBcP7vae1FgFIpk
8oHiZl9kzO3V9VxA8aeLa+EyKZe1cXVAW6lEiHaNEmQYsspK3HbdAg4aI8B1BGjW
DN7ojQqat0a6tX35EF//vruy3M2G0joQRIZ/rmRicajt7P+K8XMxIX47LioSB/RK
OreaPk/a3u6El6UnOh+Q0TdnUZDOkWZY5y8w0mSPnBm+pIEhun0lsYMMjpBKAkQI
SF5CsRBFIPB880+Sd77VfqMrLCnWAaMwbX66+8TterzwkcBt0HPV3MfeGkKb5QEf
H3LA3Gcn6s0/njm5RazF3oqHNlKAsIAP0rHaNZphS2Ymyob+CHyJCwD92AHigETW
pI3bluVep6k9q8hkXcMeiVxPRgg3Tl8h1dN0LHv4W5XKLGFuOdCjj96F6nUP1D/N
rYtNCw9zxkgCKYG/L0YywdUr281ao+eVVWZl63eKJvoMQ6tYFgT01INiyRX6WOpr
vIBlszf/UdqU4Kgm7JxjhDAyyrG518hvs6YUWUP1UUfZErh8Hg48Wcq3/sO/Fh07
5lzItqq3d9A8MBb9lYk6gyxne5PuWK9jSJ0TcLx+WONzXr8aXwA2WljUXHjx9rOP
3mkws8NkPaHhSuDvICck82up+BZqt/rZjL6qvR289kn/N42tU/LBx30vml9gnji1
jNUYaB5+jr77aR25TRQr2OUIFndA0G3f5wPXNrqLvJFFFRxciXvcVRO1yJrYYrhU
vzv/lZ8m6pAMbIYccuGdtK217Y0c9V9WiozMW/lapyISAmyfq7AZy74BH3H5EJvG
zX6AneHdoFu+nEmv0vtCZLWvPif0NT81x7L4kJYF5f7EnjxUUgDHDjilBNC1qivl
ZyyHsTCB2Mu6ObcHdG3H98aKVAeGpvcx/rZTPpMj4eNAIb6ZN96gFkLgo10hxePc
PNJ1RoUZA5o4ylb+uXdxjGJtBzKl/x5BQ1WMmWIDnQlJDRxwIXwGf9sc2teDIMC5
kaib0wykQH8OzQiy90xImnac51IeDV/wtuUN67nAaiEnLQR+grJ827A1gzur0E2F
FMZJrfDYAGMXvpRdljT0avP8O0z3VgnRkEralbDecPTimjEfGrc5w/WSdhY/T4eq
vxrv+SR94BORwLEMU/Up99vlvlkGHEhMRuUSDkCA9Zv9SMUXMSDZejR8RZoCL8B8
GiTnblKrKgOuLp3Qm5anu3LMBy5+qF15QuKHgfC/3FUXF+BTTAiVmOpBq0uDm7Yb
4UdEXXascMmA0O0qusgpfrYMcOilwrdP5h0BOp4v390WTAXd94HHJBZpAOpxkTXP
+Lq/UeYFVR2RKihpqOubAF4Zrg1DVM65riuxjYE0X+mBbW8Y8GFYLcEeBB5lEOHj
gHbRQt7Ogxvnbt8Q7l/SFPUHHm3PIZo9M1nHbnuHV34Pc3UhSMP/1QA3J5sgJSZa
b3gW0jFx4YzntiseisKoqpq33hDhdec7zqBFWKjKf8YNU6BVdE6eUV3vtPYMjiiX
XMrM0uJ6ymjcGs5P5xE1XEpUSXgl/zCGlMMt6MEF5rLnAQU9LiFQfXTO6wdLyA7+
FqjL0RPImphcrQkbA1NBWjAdPymn0OKQR9aqs3QAfSTDDGvKQynTYPaVy0woTprb
+f45DcGYUjFP+acqfRqq03RIToz4ixmhcCq43exSz64RPgjPVG88sm8WQiL9PNjB
NnbgEoLgQ8lUgYV0CFiR0Lb2qKmwsRKU8jq823gsd9I3djkkg9yCasH14rcHhWWo
jpisohbRd5Un3V2N/3qrgo45MP6mQ5GGrZED5sq0/YOytafSnnv1LIQafCiidJsQ
nchaKrXiVs4l8iJz+jjLzatYezfRQLYfa+/JAt4gpi/Rw3QNnsU1N/+RBh7Twepp
vpnGveWY1vgnwKVayzvn7S0qgqb10ayAxXAN4p5Q9EEZXxLgQBexajaR1JtW1h3P
OMten7m/rBsbK5VPGxqbxPISLGgpkZNW+7AGHcKP8wZ/FJHT1eptuHgrcrfF4Pdu
a5jZBjF/tMYqet5c5w1H8NRJJ395fPR7kCrmzKltT/kpd7zB0KEWSNXszLwew3As
1kdDOBBmdZH+CoBEQCoFkQ5IcujjZLqspFvO4bHI8VxozmABVpjfBG5yTmzspTCF
jcJBowfu/p1zLhFL6KbXssDgNaklDW6WFBCc8qObBnlZ98rIj3XRj+BAalrksQWo
VC5qBjB7t9DWJf43OdeG9LP73akKd9E11WB6fqwOObxQeqhULp08m1lUCFpEHPHz
4keym/OLPBgdxydXskjW/Rvq2YdTKu/WpKjkLEF4pnsLbEhQOBLuKv6rSQLekJ2P
BCjKPiboN4+C/YgLS59HI0wjmXNu5iLTVPyJKqOyWQ63Ry0tMvvLfqGDtQOlQr1c
K5Roq+bm9Qdutrd22mLxcNWA6LxSSy86A3tq4jTwiN9F3ynyBu2P1fTS+Bk4vB6D
tE3U+PlmXsA1MAvcyWKQiBYRmuAFd9+mEIP07KEThTDqGsdPwue3PjBwjdMFfljJ
2PtTa0INFc//mTFnIY2QwvyZQJ+RszlwFhRpBctUhzK9toT9heYo2fjVHV2VcbMd
yefFBVUylC0s6J6TPO0ivabtEUGvu8TsSrAz0fnYVK26ulPxTH6uDNRuhMAmoFcq
WdXu1Qn1ZVvRzSwMDN9+N5cGJYZwt/+YiL6Q5Iifo7udnnlZw+mnIwcRlAP1sVXn
pZHQS6uLqDDuQ+rOZQf1kIrm1a/zcibQMEiX64GxfNM7shS5AYyyGUklHlgwdcGS
kzTJH+iBrnts8gEbsmB3rrxLds1FIySv/Jt615fTwMcgUDJfOi+959jqYG7ng+5p
6A/3Y5y/mS139/QehWYfOq0zv/HQBPNzRm7ptOI0UuQ80+8eiR6b0ZXBy4BEJ8TO
L30HPI3xez8uBBuGa6cN+vfYgflnxn9HMKLvPiQrP5D+d/MOEDYF2CesfrheBpB5
4kbItvLdtN9jwluam0bXA9/kpd/Lqi7nbDwQRysVBtDxeuSjxH/aywnV9KlWVGYj
F9agk1rJ3T68N9h2yri5RFRcV8Ob0REwJass1HtmC8lufR8M38Wv7/mDqUrika7P
ZMJK4P4sEWr8jS4nASbRXE/4+iweVWqIxeFOC3jV1qAaEjGw9XWdV40BFe6PA0nI
Gg7gtkMZbNwmlYi4u1VhasferzTvjk5plnKT+wDtyeEcJqqDHz6DJ6jSd3DTDNqZ
gMeXn+jzEdZPAfRJEdyXtLNRSACZZG89RZVoltNvEu6CRBsvLq3MUckmuklSR5pl
NqtsF56YFKW2TRD08/cG19Oe/p4fh0/KG1pSf43jd/YEe23YEe77VlNsX8kpktpw
LYjQrE0RhMIak2WW1seFF+f+Mds13JivfkkqZMjmf3tQjviqiaucMkEgV3kTcaqu
pnFYhswV1OpzUmexJSIqE456+L+nBXptOfuTGCzoHDz/XWoYGB+eVQhKQ0h45XaL
fyI3Hy5xfCrpKoaD8gfMvqOAQrHjT1m1zarG3u0+LB96p6HeB+gA/6c2RkYDS0z0
sDYKiD/fhsUOGAoRyZV+EzXPDp74qeD9pUa6iNoIk7Vq8rfZy4sD9rq4rV7FgeLq
46H9U7wtTj4PaCVdB2e3ZGheOeEpii+DgRFudmj4a7e/wGTzfxhvVjs2kSA53K9/
IBoTGInyh8tus9cDIZuWT5C8/GqyUzhk1cI/wCLsIIzShaPg1zaBWHZ0UOkHuCrT
VWdyvmGXamSJkjm1nPQ8LLmudZ3ePfto7yLBB83UIsXoEHFJWgrm9mzjk/kpJz6c
ws3ZCHDCOJFbX8OuQPv4CWWrVqk4U4wlVaCxsHPGbGUA17LKYEQiFOktpqV3kamS
aAo3JL6JJY+Gb6TTeDO1xx/sKqHNjLhQwXCNcGLngRY2SgApmVdZW4YmYKQCix1X
nx5tqrNjkEAIF0TLybU+KtD3459+pIeT5F/MmtHPBHGyLckeuXb82oVQW50vO+0A
U81e96sZBA0DT3GIdZ0kOJb5IFBVvt5kR9HkilMofbbLAkw9Jklr/mm1MEive/M5
17Dsns8UtlrL0M4PANCq7NlGoSpJhSX2FSvDN18XlvK8ZxvxWF8Tgsj3QlbzEzWP
PBF8FodznncZYJGuYGeBEXeBdxQH4+yjy5O7J26OX6tcCSBZgSrSNeuCZg+/U96b
f9Flyj8j9aAS/6edF9WcygYexV8syIy/amgrzAjfaaj1tLbKf5zp/fOS3+91rK0c
VsgaFs8+MBtu9QAds7uRWmyVWMe67tPmGe9MkvTdIqounvn0Kx16zRLJaZ3cK91Y
yMKf/+vE0du2KR+B7KtKrdW2sPw4PXjhDyegytYOuWydg0WZQlY6qhx3mRaDyNoF
ElYP7va+JvXe++vhkTUGJfGKzwlx7HuQG5cLD+nhi9PgXQl9QTrs9f6rV9s4mEda
/Y08p7OofJPpwSJrlcVGNljUOnEmsc3JZeoATAemYQrPvFrmQy8PmOf3ACwvVBTs
AJ8/APSunKZIv9DIWZD0gNxZ/RJwUFHOO6ZTnfN4LCqzMIq6NeN5sMcp5d8fUka8
f6aDgvI0cV0raBcBMuXHkLQ7s46PuoBRlM313Z8rPB+wBCKZ+XiVvfpXFupecvg1
MwzSIOxsXFx9La4TslmfBfICuabSobYGsV+APx+n9682KuLd6FFLXZl2Ea2C3agV
jhCUiUHjZSZg1eY1RqNSjA8NAbfATNG0joVItUwsSk5Nul4xtaa0HZDNpm//mwA2
2RYIFORsGn8gUcIkm+YlATenYxZaOkRO/FfIR8SODcwVEXAHmgru80FP7M2Bih//
ZfZpvfscP8boYEquX3HVBHQq5lQemBzLntOh+Gam5/4kOoNx/S/FJFFzYx6F3iek
RRGNSNGh5+mP/72dKVICQUPWfJhZob8FtdKmvDjMXK/zvGB94pj0wr/K3IJ+yCov
BxnFDbvWkkaPnYxnhUpGwySqaxCN+d1ZaXgO+vBiXysuHOFvy8lUWAhv9dZy+xU3
s6SMfoKDpTHkYZZy2fnaNzTlTAfchXjyl9nk48xDBxeKSOJbdmA5SYTbJQRSZQnK
aPtGXvQreXjiGf5Ro4C87Kn55eE2rGXjthJxZlSTvntXbKCkNpmkguSLDJeg1X8Q
o3TUp5mUnWDkVa0L62dIvIVNTduKA7XdFLDi2Hsd58Dmc2UGyyxyfr74mdU/dpf2
RFTe5b5pe6wrzmdtq/LmzCiWBONCp5EE2MqIUvjiCHytFqsn/h14Gpr/gnefN/OK
xhlYqlchiO0rNI5xkaT/v0ioaqw4pxD+jPMMzka7nrfAOeUjCkMSgP3fI2ARM1ow
cCk2HwwC3LsheQdbvTUDRpR2UTSFf62JQcxN0CO2zm44HydVjrOqmi+573TDH3Qg
PNdKBSK65xCLmwITxl1uzDyzY9zPQMymI2WXIy9fPERB67Al3k+A0xeVl9ONmviW
hRZRZeNcdruSmeQJDea7phaRw86oF5ThLBnUCsSzVl9p1nNzB9aXjSjoyn3p0HBR
GwMG8T5Z0n3FjxPGeJ91RwjaoW1k1SL/8dddqP7So9FM5hLpXReFz5TS0ev9fU1R
/mp0naP6A8gjKY7fw3nwBemGEwoIqF+Urbt/yltDdX7nrVfPpBe9HuRDOSkg07Hn
fjrcrgfh5O8lOcMyCUVNGms+0X6M9IeTpqtgh4RZq18utgcBPJOE7Kt1u0zEM0/6
qT2cVp92jrHo4s9um7ZHQH4d34FnTE1V2d4w5X4knUAfVL7OSTLXrJCk/tbMTP95
0niAkT9M7QS9etAyHDh437SoKVsQiVkJ6CZ2KNI3UwISv4MJP36TQHL8T+xcOjae
/9Vvfzdj42kdz7Ih//RApZlILF0VUPfAlLgnm+fgaMdUKNOezpoM0Dqm2nPC5iMU
L0yU/uuiQ7qILGduem/Sb7HzepsvpcIKFsFDaccCrN95osGjVgjzh5sQ0HpSXDnG
GPrAIpkzvjUY/p2XAv/nZxskvFT5UQfnXIqXtDl0fv568OYFY45nB82C62ucIRBv
GFgXA830nTDGhL+yL3UyDWHeqQXb8D4fUUNu5ERMS6/2k5CX/0zg/Qr3DeFi66Bp
eNrdT/h4ntT7G0LMLMLG5LQEcKeBDbgNqSCUlIVUqUU7LlWUZ2JunzfQndPNAd8r
5QbxW0qrAvbVLcsl59npQUtCucMhyFUWmCAQ7hqT9KTGNFPSwsZAa11MJDeT+CQS
nZrzhhJAtcf8bH3WNoxiSj2XT0RYb17Th7wfMxvG2uJSIgPYXU7rsjgfmEoZ2M2P
T7eiuc/P9qwQIvyO4BQBSmg03Oj7YcSP4ceAP9amjEZzE5Ml4+jB7v0WR7F3Lu6u
Y0KsGkealSS+PcjwAxdxHPXOLmixtafi3dYAg7s9bj+/cy3pvGk19X4teVy9VLJH
U+ppF17Pv6JOIcXjaNR3jwelZ52348g3nkl93WT7WTkKEtjhxdMfWCXaAc8kHH7p
nVB48ZRF1FQyr9xFYe+xRLVoMGJ80blwCsGC2oOgyA5C7Onl7la4cMVFuCDmsQkI
sE8bKQCWnNOPrlHXi3hGP0tam+HDtbWG3dQOirPH/g5tMSiUtmzSuVUxfOAhN9NU
a3f7Rph1ewkfiEIBF3gfbRiNgJ+3DjB1uPpDVES7EOWdCniTNI+caG17gkQOKBm/
54NeEoC69d8K9cxF8Gkg8MAbkRVeN9rzDDZxUtBcHbotEXnfmsvaxjohfW+vWPQz
55Lppkvs3fhhWOZnRMAtyEf3iim2Iqv1JKqAnO9G0Fm9YyPyuvAs3OK8WYZ6Epgu
NloSEQCOPMGzhA2mKXHtjcRX98qTjheepM6SnRvJ28TDg+X+bA2T9LNbSufMjqqs
d/dF/WSuGgYMWRrx3/qAb660P5NmJio1oyzUYzJwmrkHsnh6zXbfPv8c3VSC/3Bt
gTVx+tf2cQQCMSChHp2/aBEctkSw3aTHTS4tN/2DPvaDnO9C5fmkqL/slQcrI0pT
RmbHdqnTvQGBlpm5JKQndPNOW2SLcIKJZa7WEsccHB6bgAObSQFVrrgxsMLVXkGs
F7uZEUPX7e4Y4LCGroUiPVxS/AorQ2MAfVj+3BTzSkiju2y4AjY06HrnK45BBzgn
NIxYX9sVXD/441GLgqu3RRNP44mnAej/Bc0Tp4U4FWPYr19K5Pa8GHc9cVIzzWet
Reci37rf4WKy8Kt+hjZYsJjHNr677J6xwMekJoc5Weupjivrc0VIfw+93FW/tSiM
q/JqvAhwVrsUBfQNiW6Dc7DmSOmhAgGj0hT91g5sh60w7RRsdrWDw70yHZJV5Acz
SyQGcXfAmJgjyZD0x9VKlJYU4uvQmdYpJmsTnDNC3jRZqWdRdihCW1zQ0fe1fWp6
6eX6GGxOaTDHeFTkkWGiDZcIj0tv2mz3SvT6qYg++AF5CFF41yjnm7A8k3lnegzC
AfIT69r00jB9lBbN8V8FsSMBIreUEAabvA9YxAYroDE1EeK2SUV3Ga119mg8cyet
USw83Io+HFyJqDFJcsPUASAwEGCpoSxB/vcj8G1S+huh5/aCAas6lv7DdaJ38si+
oIRA1COJZZ+DtOSgP2PY+cWZ4bUyJyYLrlPLB8HAeJL/8ipF28tQXR6Hw4mzdagn
bHk07/YzSiR1FZ4TIXmJg9DmoT0ZpFTdUmIz3mnPM9B+JZG9WthDQvMzSxA1vzyY
mUuRsXMK/qvQqS16lh3JI0n3NmQXAgiMaKT7rWzBUHmZX7k/mgyzoKVnBjP7dkOW
gIvTD1ZxXvnAB3L25G37XePaLYBwlc5JwHgixVmivOWIvworfhDgMZn5xawKxm6I
b9aYtsBKxTn528/7n5G3RO9Ul8Dn4Gu+CA+lAcGZrGCau09ERXFINiYRbKE3Ds7x
4NMBDZ6aWOMY2Eh8HVLGGJ91JSSrnrjd4OkGwMoGWxYTmHyttwMdGm3UIrN4RwWb
2npx/v3GtxBuvY2V+8euQixgH/RKCQyGQRM2oe7aWT130rdamWNuAO3tGsX/hG2W
5Fz936Cd4KjJlNS4dvxf9j9M08m+eJMn6rQnpkmJNUpGMlatkzndrTMIFXAPsIKD
pbAYSX/dFRnGF43F7p9aBTpEM4E/5spTaJgFv5mpqPZTA1aI21jQKxfVqzNGpS42
KIFWOupjbEXip/oNzE5Yp056BjLPXkoxlxLROklmUuMBkW25GByKijvQcHboI5c8
DQgl2+3l9OvlPmNquJDI8BgIPiiBiKO0gXyWPNaNhcjlasvQ02xH29KXXkDWQV2D
OKkAn3z962ZZEGeDSCcYL+7epQjnD+n03Vm5/OzTUZa0XJ6ICWXHyM/hrNaHsbKG
Ah7+lwXaBtP7rOdbR94hY0DpLu3/sBsAwX9t5LX7Ip1PxNN2bFqnXOXxNEbYNuOq
DXqY9FaR24W7USR3V1u/n3IQo/J60AtmvTKxvJkLw6k98hb5JJmX1YvyqCubCwAq
TM26Y1WWPj2SiQDZ00ZMUFeTLsA0BUg50tXCDqV+V+YB2fMEGfzm0rm+oY17cKza
vMd56fQ9E4uec0KhZTXjkjsNI1V+SbQVZpdiAl3l+P0JzE82H4/8IPvpUYgDwy/y
TIXdU7eC2dvSjMHLIHGDQKPcQ8z9mvAEoUIMIcKuCBbVd5kq4+x+v2VH5BlfhC1H
HyuhjrbE1nmcNpx6xorJ55Id/kJSs2ZeGiywC8yCRaWnFrYva3hKxxFawkI+s1nN
dFubGUggs9zzXip18gy/GZ0KOq8vYMQ/fonfrys3UEnWOgPtMI1Fg8pjzn9SUAkw
OvmZzr0V5UlDGA9LDJ1AzN+3JTtt2XppJVWCt+L7M9b3/3jlZsXYY5ZJ5BnsAXKL
LWbmYZgdB5kapQr+jc+qG3Y5aqx7rtklwdwKXeuUJnwD+HlNfPw5ykefMRh5jt9c
/MqNuw/l4Vrp7RsjX5UQIpho2gOyst8QwTMYS2w4GPleuGj+fS1zf5WgIfnLyH1A
oqOq1ixr5FiUeLBoL70VnHEI9G9luOJDyW6iV01mMDlldBaerXjWOloNwvXT3sk3
F3GJH8bgpvmjSP6zOXjTsLWgazKqWOSi2oEKUcIrIZfg39QtgAIp7eKXurt8gY69
MMR3esKAOH1hoQwVyk+yNebQpcM44PMAhqKrN8PyZVMVx+NWNqJ4QFtLZmmqoiOR
ROryJQsczxzEQd3LVwpMMYUr8W6pCteXQ2xSF96AL/Gs8SOJjPMAU8KHwWqL7pDr
V1KMsUGER3Ad/xHA0XyRud17toFfLqN8yMoe0bRkChNeYnuefDVPRO05GSAAU57c
macydc/x+SmbHYeHNe3YrZiN1iFfYE21/Ii63ghr8oJUFnq7v1+CfFjDO4RKBnzE
l1ZbQTsBuCCWxsfavwjOAhj6LzcOgMpQ3j65RBkPLaBAMau0ZS6y7PsiLsLzzced
9+t05qyAa2v4lD7epSS6bmxPYblCQNaGjur2MAPj9GtAWfCaQh9JTtZBe1qOT7wX
nNVqRt1I3WASBCqteXVUYmjLKQj1L5bNWQIDUOveQZz8JfUnJLWGyusXclIwU+a8
opUpVIEQ9uKCycjthuD5McyU3qZiFaCDunGMtDES4kR0gfjBdBt8wA2hPxNiW/wi
J8nWdRwwfKCy5kHVxn2Hjn+vhtCtR/nfcxIYK9/fKpl7r8SdcfPIt31cPYLUvzZp
nSxUPf1rjzG54GdGnHeswz+QpZwmbAXkCtBGpRilyPwDJuQ4dxrZnHVZRCuCwsOo
ttxBFksX7aoIQp4cdiKFhetH8wmbnrfriYbfeIMQtV16YoNXosNnkHaRc3lufEhw
Nls8FaOVI9KraHhja22oBFh5q74HNZxMEAK3RWyT39fM0JqtpsjyELfY4P+WfseL
6b3Az8Segmt51KlGW8NCVYsQt6/XeqzElt514lLQUENvGdb1njHXYgwjexLmsVg5
aswyngjHMJM25ICh67Z4vrCsbFiv3cAkplTNhu889JuPu+BeSUSfyjIwZIHHB+tP
7Yfe//6D90JzDFlZ7UovsLbUQPKgQ6B1AWWJKEwx7RphjyGgVNuGoPvbkmPfyzFd
nz+T7GlCKXcStTJ92UaF3SRmUI4hxCwUbpYmFt0ACvEVERT/XRSBr6aa9r/g2E7U
Fg2P+O4rvB6kqa2d0FszcGxrq0Ag+BHVdvkXqdPAky2B61K/nRkzz1Ldqc+4+c7W
BdWs4IuuaMGjwHF1tzOlS/PANE4UntVsBiMHzngwIHzqYWVRWb/5GgSsccx92uh5
lIeNfHDyv0bAO0VFSazHwi66PqcTKWvn/jwjtiBx2ky1yoO3LS0NIC4uogUIlepX
3xCePuqBKOOxM6x1WCWSmfrj5t1kt11kNqpVAnzuDXBUnwGpSPRF2pe8fBPmCGZq
J05mppT8CxAV7hNgLQczqGal/qHGq9keVUQNArgpsmlFoVv4sggg6Bs+VkR+xnN/
to1N/jtZszq972qlpuJ74BmwhnCBOgetcXku8jWiK9/+JAnMZ9U/RqXwUJ7wBN3e
gFK6aQJmOVFb/PgPTxfNZW1vo086+0vD1Fdvi45LYmJ9h9fn71wsa5AYFz7YDmNx
XTNFJlyotO3i/RlleTaykPoRyv4UoLG+9m1M2cPGRDKYkDDAK14FqxvMUUimbKda
8pV4dt2o/cNDGvBTBKnBd3/JcvvLHb89qU6i/3ZHAaPGnxj4qIkQ/BRsSOEb9ekq
ezU0wRcN9+X1QU4Aiy6GDRe1fLtYr4RXUJRuX1Q1jxtjR31y+Jt7lIttcbGcoMWR
+WHU0K9lgbR+8fEdVZfQxe7vY9GP2fCEqwrYsGsZbYkjD4am8aB8KHctbYjRVuQF
5TJY47arZXqWjY/hHNmVADeUf4FIbGm+P+FfI2Mlork1Ig0pEVdSJcTxQFi1DwyQ
Iqa48RCdqOwb+oqGuesSIA==
`pragma protect end_protected
