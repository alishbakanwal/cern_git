// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:02:17 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
RIr5DcdiQ5/wVWdaEqI7kSiT7RPRM8iNxdFQK8Xk9hQpVhDh/rBJgzAYFOFJo/6e
qDt0Rh6xChNbiYSqYIf0nKJV3mR8dFGdKPZeRm09Hou5nghckrGi5RQ9GvxcXa3x
4z28isAY8UbF+qZT39IN+UZq/r4iskIzonli3eDcCqY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 32400)
4ZyqD7he1FBtcxP/WNeQn5ATqhzqb/j7V6aCy0g19ngru9COVgDQQgJ9EujQsYVL
aBX1whylRuTKe1kIN4NXE1pysvX7h8TgqFzyaABsgzRsJ4sbTBTZUVG3cEyKwNsq
V2tugzclGN7KUCmITxOEF5V9V6G6eBvIhOsWuV5aY4WXy0jbYl7WcSGqy3YDVW5Y
Smo4BUxGYgG1opKV8/3pagIzfpOjVGxSfzRlJl2suyexEZv+MAYXwpDqdnj5zZC6
TlP9Bg2NYKml1OT3r9Ga5k3mtSA5OcRI7ywYuCE2TXNbX7j5j19jr0nbxPuy987e
e9B19e5PCqtfbsCJd/5T304tt9VjxxYH0djnglKmETZWfRUfUE+3QhgOHrsePO40
5FOXcrlVHn3u5DySiYlngvQOVHL+El54hn4j1ACh3SXfPe0eqAO16ecciLmkNZwe
D02vtSIFuUUG47sPNL61fv1AmQXLlGQ5Wr1pojB6eus12tCCvkbyoBTIP3yUHxem
bWWz3akLpSz3ctM2QKA+rhQa28SHCXNHY1jXzYkKujkLucjC5tLiX+x6dxk7QuNE
ZYVrrBC2JKwcaSDzy3AXuZRlWqtN8i6zgdaSViUMwUP01UuAM4Va03DYz27Rgch1
RBAFUMKDP06ETK6BrEAMblZj/ZtsujioNiYiWXH9VqMLHM5eUEF3V/EIJuSgMKZ2
DJROGcoPXdTzegxeEqJlS1hck7wuTjWxTZPEDmskiFpp72ALZ0yYaSJp7KQ4ETe5
RWinkgXd5CCuuIO41KYC/WAxf+2n+3exk34mLp3TYZos8JYteSIXhTw8AI3lJNOH
+AzJKxCOMoQ6jzLXef2TZeF8dbTzPVxeIFWGkFN4b1rQjO1VhvyWoYkACGxkCyFx
CgIECnKHr1r+oLwQQGrLcMRa06OgiywaQE1aLfHrZ2wg1Qnhlj+3LoXf6Vve8eAF
yVdb9aYgZyvtJVU7VPkISDkJH6NwWp2n+5QXTeW5hF8IXvBxVAkUnKcuCtgly5St
AmdC2ndTlgfjDOghHxRVP8PmhhnQ0xAY/SIJHZ91BqOvdNpvUYuceyyh5aK8pKV2
MNwAZAe5vpVMQohveh1OutbTCNY1L2zpMywm0kzquW2qyg7itnIhTuvr6C9dtoVX
+OioAuOyOg3UyM62I6pmbe+EXF8ZN+XWWuZRjbUBNQJJqD5ME+4p7phf6wPHO38E
nBLt83pkZxJCjK3cHeijKIFJstFGqYR6NOuKJwl54Vo4Oyy1tJ7h58cOsoWAXk39
f+hZ1ZPWl+jZRClXXoT5mbZezyqfGANKWYj1CYui6zWa3icZuD2X2ipS5/fNNO8N
LCDeVhowAo0PXo3wTUc3bLg5BktL0G7Y7YZJSYOhyPi1juI1l3qEiv2oadChWNfg
JYdVoWmAZ81cH26NJdsq2L9Xh86/QyHYHDmPq6nc5LwHQoNlSVfFV+aiF+mQkXts
5nHX1tfs88Vy5Ke5tOpQlm/X9pXx6scDB9qdXga+JplmJzKWS+GP1AI21e1Y2Bce
q4sQ4jq6tc+UkKz4197/wMZ2uUFp+kDyQmS/ZXvLDL8YL86yavt3FXR0v6tz1Qe1
/CffCIYudIdDOxzOtnwqCSng+5nK54iuUAz2pUZWT5deYl2NnSX0wQ3Ei96Msoj9
iXY20eFPbeOnQvdTyg+ETHo+WRlKntuhuLpZ8n1SOQTZa/JH4YpwjYUMlEsA8aPw
hWiDwUmt+l1SBUU8l4Ur1GnjnXWAPX2yE5BlPZ9LzH+0ZnUybZrg8XTZ1xrd4/v3
YRUjq/26/zK2XsRKMskPT517Y5O/6AMu6rLHGlwKOjZ2epvT9DllePHb4BD65eRi
3tk37ZGTCisfCMBUSL6VJjIYum7dSXrsk+UjyKV5FyXYNa8rQJz1lUl0fO5yMwnD
oG43nDICOCKO205fBoHJk7JB0RMgrgw2v9F12SzgbxZ5RUuCn8gs/F+B0lrm69YN
7x7rp4VyqL5gxphToeIh5d5yU/OvxVFF0q+G50bM1F9bL5Ke0/+7dedFmsbMO0rX
phvLpo3rzXCsgH7xsPzJpKlrauki3lNcPO9PTKDFIShMVjSyrVXuGvcnxJsbLe6c
P2KrbZQq7f9jxAGC/r05VhzhPUR6UzgcxzaYnDpoDGKjrsGWdvOLbZb8SeMSdjeu
UdvWt4UerI1rNAb5bOKR5whRJddbtjqSHh+SjECIhdARNU4DTnbN5tPcbjbfpNbC
ZCs/0fITH23IEzBPKa8SBEonSunE5QjF7dWqLHd56iAIb+6QSvxCbzp2muzulwIz
RmNZiRHocMnwnVhLhCY6kStXNgPI7ugGiRWFRkenvm353GSdqfdw/+8zrO+SmDQd
V/0xIWIANlDN5nUoZHlCa++fml9PsCtDCI1X3DZr7PtpztzGopFxIm+dZdkmYI4j
oHXLLVXzJThj/LuF2NcjxsQrpxSimDlf/Cu45Kop0N+EOYhPa4dxC5KGnM1APSXR
inzeY52pap/CrA6N/TS+uQ/tzsbAB+X9PyyxllGkaQl/uiwCDagH5I7nVgFFsXti
D+4z3Gb99M1X4/4sXctgkfmOlCMLCi1DGj/VvjhOL0bMw6oF39KqHheN+8Dl8LSe
4llnmdosgFw00XNo1+wnX+GoLkyAfTaHyGZ6fUddAokwptGOVf5a8l8a9FbBn5Ex
C7FCzL6ZtxeQRUvuxCoANRb/DsOp9oD44KBFF8t2GZnzbviev/287MIvLp6LXXTx
STqs44eyHh3bTHKBVkPIu1kWWjd8H0L1VmoNIlIYr9dsTggSrXuMlYxcVWMsPMEl
1uHlhn1MeOQ4CHenMyaH77sLG9gGBGju12OMITjBonMq4JHfgHBRyiHzmzj/Scoc
5aquXU4TVOIlxrlyd6vVqybAZmUysrOIRlGY8OcH2iiVtnhiT/MW6o9x2n4VKpHI
MNgW5iJ276/B8d78R7o0eeELN1w8yk/4keeVlojEb7UezqF9n+5jktw3Xqmpijfo
e/v90gFlkxF53iqrGf5Yf7J2C27PTYMfKMzpD8zjS66hmQMNt4fQpn8Ev4YdjSJh
cobrhDkW4C6wyat/gS0xcFf3k/+fq4rvO/biU09xSaXmTvv/CBQ06u0SXAMUdW+4
rvWgPbC9VhQiEtaljAyMS7SxjQZdHdE4A55Rwdyi05elEp3H4Da6G4L2lzi1d1Ts
R0MSyQg/uOv2b9MXmnH+QuXB8ZB7MkSpPqqYYulVJDTJ5vKgYS106s8sPLcPZnss
jOOcEuHbbsMVef8eResk/nivWSoyQ2hJVuYQVGu/zfM5CBWAZPJvJ4MiEwAOdVpr
YixB4lc6eVlg56pCauRbVOUr9WeWAAeUqbK4bSRSPfZtIHZYXIvvNohrdojwj7O9
6+0eBL/d1xl+gI0jrs9YPS12h6/cAHI7vWeJrfgJAb4XfOHS1TQNfP9zzmL2cERm
jRlsXb/M/WdAl+u4dJGonq3BBqobpu16v+/nJdyY9SIB//pA42rCOOv9JCbv9/bj
M3O3Vb7t7DCPw0xL6OW+ptsaBu7ghV2cYHXBSxPXeS0A/Qu4068veaP5VAj97IRa
S91I24g6BeK7nchXHljT7g8mXWontmhtJjLeGU8I5kjefGKwwBj0imb0QO/3I0Uy
H1tT9LBOFg0Koydjr1pCjoHvs/MwRjQfcPNHpnC8Noqn5mnqUq0/bLBI1LTcxsIW
UYTzEMxHuEYmsHa+njpkrq3FVupvmVlE+49NtvR0j04JrgUoqedtJtLsVaV8O1z6
iKztgF5gdR8sFcZpZtt7CGaZiUbW4P/go3lmstjaoIu03E6fLdwjPnW00cc6t5yQ
447qLbrDjuFvuAWjS0WNSnVhuj1zBMadj3eQNXC+2TDUMmzIgJgeLpIJl5dKP0AG
a+mdaHvUnwcM9bH5CBeEZnSiOxkNT1j+tquce+eYdWjcVZsNlDMFtMNjnXMhcL/G
wb/6pIiMLdSNhJz7zdQmsmzY9ATU0t1FZ+3Lb6spavGNbZbGt3q+MW0i3lLd6+wr
wEpY6JN+HXMrP9qwCiXaQVt9yjmcmEI6UN/5dM5+cL/L4KnudV5qPnguO6m7cj1+
qUoTqDMwfflB4pYuE4S3M1ga2ZVExNzHSBPglr5qBsLBc8xcifQQ7RsyvvnMh7dx
/2+10+1nAZynmi595gqDBDRfI3n0yWIwCqbUjdAmyZQa4TeSudNaR9LkMZtrQNnj
eAKagscXmtTsUcTRotJAOuC9gfoVSSHLAP7Cw7a7vCADCM0HjbXMfU+13trrJExy
el2HDUPBV7oMBrgS/b945iugxUSGlslI1cbJV/bow/n3kppGpGsqdj6b+UQYkM6+
erD5671Hfuri+r7mLfUVPGvbFZY9LT6mdLmTGPo6ba/A/GT2nP0P9B7Ij/litoeC
T+zDJbKPzGu3Iqwze5Gal50t/Id48e0xyyIbwlZQozRUS7rpJah0qt+qzNsx1u4H
nCUVu7tddCP/v3EL4fDuIHN+rI522MQjtvmhxUVuUku3XsEqppyuEMfdgX1W0Wf0
aX0F4P/qWnJ9MK+ABAxg/EKmrasM3AdKsVsKLI/Nq54fU0HyKHSn0siHZJ5/lAOp
Kun6dHaYOMkiEpzKrjSpqotSk3HAH8dP/Xe7R4kY8lLaiTounGxKnxgkm58Lw5xj
jJjZEPCEzLuRrWSZl0NJzPP8MJUSz7y9J4hDYTkS8jDZrDTrxogaKVvJCv1C6Hzc
P1/QFZg6ECooWKBE3a9Hsd+krePPJTt9O0dOkDcGnbdGBdpjbv7VBQYwsRx9TgqF
lphIxjoy0jx4eB5DC6SnLB6hj5bJTwgY49A5tUL3A/AL4sQAegOZOzrlgw05DO9f
QwI6bNlfzpKsgeKJj0mjO61EPkxRJFcOxcvY/yz7QfD3I/Mf0ZjoueOEeKeaFb9r
pt55v2uJcY2U9rZY/CoJ5ZoP2/cOOrHs57W3ZzM40zgVuDhXGt8wozIMr3rvEXaN
/NWH07YrS3y08Kfjz6GBuqboFo4XSZbIG6q88tVWLqvfItYrQAO40xs0eaJFiHiU
8HmtEw1SsigUh2Hla3odGhCoDbF4HMED5qxBqYWS0LvVXUtKXbjZ3XSzXugSAs6B
luvR0PTA8/5aQ4qpDsMh5i2ApC2j9EjAGUtG7M98rxlNsXsrPRztalgCV7HKphGJ
kaC/AHtUu7D1AHVDkf0gxtwlQhwOU1RKKb1pCtNmST0DAWeVWNTwFOThTXbxZSGe
JoxFdkJiz5kT+L3B7zo2lUauOnMlKLUyDQ3o7MRdEozWduUscgp/B9Kw/dsTAJf2
gRY46dfhDsYjurCm/fyiychpN6qzysDU3hPnlIUiHubpiX6tJ/qCMrYBtDdUDtrK
IThGSS3w+TQRTanr+KaZqFdNopmAXcZLU5lAK1Oc2fTbgPlzalHQN+TkYZYvsEL5
v9mAeWU2Ua7SItqWdW4T6T6QP+flSdZhjTvhxy2vFjois9ZKYwWYZFJ08/YjgROy
1q1oF7HiHNvgv2RjvbZB9AklgWx5OY2YUaeyeNstSpqqq1SPkD2G/JxbsKCe68fR
T9MnSNXwJIuxDRi1DsFZrw6mw5kDxVlViZe9GA9Ft3PXUsXQ/pmFuC2SFc1Tq/Xb
tooeEQlNOWnl2pcZ58tWo2m/9r3P4oU85GxI/yu4vXxAr4lx0iwEVyor7NU0MITn
h5e4EbtuYgCV3gQtWQxorNEmjvkhe5HSjxveIFfVLIMhON7xaz4x+EtVL8jbB2mV
Tnn911Bin6ZsPmFx+cYpz6DXLYMlcwgkiMGAKZ3DpihSzP1R26mwQy2mcpvyFi1H
l/Dbt8BtwWBONkFDvEoWYTtAMzZEcj4VVjplJ+4sBzCw23ZT/OMbbynEtb2ITR8E
8gMuKY/anhRNqgXTVZilf8M8kvV8HvDpvy51Zky4JIsjREXxK1o7IzClRaZ2NA2P
bIbNSypmWfNRennEX7aoOXNx84UpssCKOzL0N+EX0UN8z2GjNKsrxR+jypTBtZmf
a8IqYkc/9EGQWZlKZWi2z4QwZttUOKchFfaZR6a2Ik4b52tION2ZjxwzedRdnRmU
125dvGe0DwefgIYCDJF/3CQzM2rNmPDHnBNLV1kwinODHD/3N7+jI1B0L/qWTADp
kmQsXty7yFkQyoLKSSePQJd3LgZF999KB3T6EKopuyZJy9V5Ri7LYkiDRC77dW9S
+GLnodEkjVCW/tilviLTCGiV/pIFoLuPfQoFLhmaKO0h0Xwxwuvr2a66vCj24Y0h
h60otITqH091SLfpst5aWL3z7wgdYJHARggMVh84UHXOKV2hvOQKOMlh8BSp/N3E
UIktM2AANkN3fO1dbCHAMRepan5OQsQTA3dAIWsxkU4Cy620F5WqimSTb+Nn5LGD
v1pNuBj4Z7E55tJc952mOVS5Et79r13x99e2XO7Aayj1/dqi88Lz2lQsfDVkVG9H
K2KbNiPIJalkoX1WDm4bAEZSgh/66nSEdKibB9Kxl8FlwRvPm1IrTKuUsAl4zw/a
3l8X6owWgM7EP6vQ6ESvAxUOtGaocrENtaPMa2t1FBxlemCPxF9ZAvFXel8s7kGQ
spiHWMBWgtOU1ap6q4c94qmRTIuKT1U3AombT4GKxoCwMDAIa7tK+qj+o6kB/kbk
kdb7vZaW7UrU/yrAB5ccwXUimj6JAS3H3ZkdZaw4uJUZDbxcVzrSVPH7K9wAPKhL
ARBU+u6HfsmBdFdQ+dZHA9BjXxneaY1lVkwyeoalrmNzi/bpAqEGa+cIBZ+ilkGE
NU0+GWYUhpDNjEN2miEV59U75y7CFiIi0Hqhm+GHYub9PYFuEC6Lt38YmeiWuLTR
rCarfHvZQRZY1Q4Xct99HU4+IS7VZJwlKrF9/JCOzWQveW0xKR8cXZvACnHTN5gR
pmydWz41iKrbolVpYjhoVtEfhc2n7cDIfhFPrJF/Q/IohT1U4Rwg1fVSEbHxMc0m
QPrk5zbeKBzZsVvQOtTqaqywplItjsyZiY+nFtOKr6NAi7P4Bv4CSmadGZ7Zho+J
ok6tPw0VeaSptFhOpwlEipGRepFtmKwzwBPn/5/CuC9PdP4NmVswuAKPgFOBzSz6
LYyPCxBlHzp5ZIBnmtfPsqHVX0FpTx/ZaZ7gNsK/UY4S0ZVr8bw0CuKzcL/4VyLO
clBd4/j8HBi3UKS6n9dvsp4s6jpL2bxQ8Cfls8gubtmioh2tVsrCqvZllX0MYr6q
ujacXVxmiFuqM4ebwr3dgnNDy8dubOe2vtbmDasRv5sdgcPoPCGvEpDblROfWN8+
QyOs1E5UBD8gPQ6LemHLdzA+szqxilCBu9cJ3fWiHeCgBlRei066SZNf+zxodGCn
OxWvDuyj/oa3atjSGMDYRa3vkTE7BDRl821H0jpaBlfPGgizE3m5fYUb5cdnE1QZ
18pHyS95fd/yzmluN+NbdI1bb2kCe80fHE01jrMRZz9dO6WPQxBScTL19ziOlhq4
+GVnjc5fu9aVFU4rbCYQk6DAgQk5WLheD7XeAihTw06z7/GE89i8NGD1HaCJoxWF
vZugvkmwM4bxdkKNfljs4vIJffULs72QJ4PBOzQq6SiJOWt4pKIvr3T0NBbPza8E
FUlsh2M1DlEgNP0DRi7hmpxFdA4lAqp3sJtV56J6Q97ML86muzZoG+z4ium1tQye
vQhSwOQcAwWhgEdCNyY0gKHrQbkxJm5QFoYC3cJlE5z/lT6BeXQcfscHRz2Sstax
jRfWsG6t4iVVfeAA1exHj7u0Dexo6k/7HD+UdddcJjOBeF65yyE1VHbB0ngP9Bwd
epklImUAV/+vEgEsx7VB2k4ONOCrZ4AUtus6d5LwdHbwFFmBdQwf8HvwzfVev2Ni
6XFdKBEta9SD4K/Xa277jWt9WAvfqsn0ZdyHxel/Uyi2PexPgiD/6d8LE5LtYq1a
4/21yDA+W26fn8XCLxHhDLEeG11QFsow8FbHWlebvNtqkRIXbKK8xDDQiOltB0nL
h18mnTM+YNfyGiAUjpFFnQICKpcBUxJT1SyOaCtDbSyB792NHJxBoP670ZxtdQTY
sNR0hoRwQgNkjI6B0osG3aOuusd53NNMk5GaYaGv4A/XBowyn/CTl1jr4qOrWGmw
9NpUz5weS5khImKsvf1Wnc0lbRpHmfJaZmidQDbXBONb+RflVCbzHOxsrkU+U5MI
MEfXuLk1egF0oaOcutDLehCTF/SdOeSHVpyXjofiRPMEKCsM3CFJGaUVt5+gkZUU
Fv2Wy5XjbFDZsZKbB8RQkrhyAsark+VQlQrG61t6X5WqujsGL6R7xpDbWi+tW/UB
E5m/rSN+PNGylmgBVubJI1Jycykrgpk4NhLm0zO80MTW3Cyj+jv73p4EH26owSEF
rYC7eMYz8d5hvkK+UlJ1Gb8ux4Yk839UZoqJ6f1zcN7cH1+aFntGdrvXnginuxys
WVh/mCqZ0Ik1Njn5eYTX788MmrV2YFDYI9NHxYYER0YhbeCj1NHR2+/mJ04u1sLW
5npYd5JCvi5cWzeEYZJrXWcGbHYpObefIfnNvtBuleSyrxkeufkpyfRPMyBUAI1x
SFKCjLODa/11dprAFQ269r38eM8STovuWQQcMKDgzg8fldiZzvK73h+GvBAuET27
19GhIHLu9/AV/Wf+w83rjWu4yRb2OGtdEsgqjJqamD4LI/FZ0jFFOkW3XfvbPwi6
TErDhPfihgUZOMJ8K7Vcabx+be7fliKSIT/PLaEQgh25M15A563KuXYhESDSJ5JS
OEdNJw1eOMq9o6HqWTaDdgKmsqapNXRy2DHiq8h19SgLsoQucMnmeiPvnrkKawR2
PMzEWZPPupyS+SFDzTq+dTNg7Mnmlcbqs8g0QitPZ/gCWpdlB1NdQzJ5A7hXQr/F
NNL00ktfQjUI63eF5W9M0RDvxqgeKCDCzDUBwD3guNX/G1OmN6A83/WZQttPTG0s
wHjMsDFCIMoLaKqWs187Dz5gXSTx3JD5b6ygmIWRn3cJiIvch8TiGIqOLsUh1Nia
UDpzGrV8P6OgzaeRsXnBSGEAgA9jnZ+TQaKQHZaMl9g64KwSVOuMF/IyRRV3OFwO
6s8BDmYlS8Dia+m6+toOAhMiZniTpYVN74REc53+jzbVb+WrV/LeaoRpmz0FQDNN
ZtXGpU2o92LVExddEsF96Tr2J7LndmOFpWTwUgIj0k1HdwT8ePjKyMdJFo/MHlVE
+v6MjuIDqTcse7t6tKGmq7my+3qC2hYEPqvgm9CW/59OTozvoo8NzE57RQt9wpup
+ahYRPl136+qzbfkE3aCQ8re4WYyTqtL6byXgooV2LG8CLj2MpDV1rXm6trFbYSE
Hc++2l7XZOL2S84+GZ08b6KDTvJsKFV4PLrQTnWMAR94Gx5fL52UD8xD3nVu95ie
s/izwByeZnRqQxedSYuxsGa+gGESRL40w2qcfadmodJ7WPbXQf1sbrb3ZhK09zFj
stIE+bAC58zKEoxgB4ryfD1Y174XwDeeNntuPnsDxRqEnAY6QVHljUIZWPKou4bs
1ChSxTNhiBp07cw3RTdLxNz3xriFmoJr4fuBFKD2Yxqgj6HRch9TXx2hIM2FJl6p
FUdAsyrrog5CWSe6qDZCh+jx+FVY30Lu5zK8ky60z6fbaObWi+4TOMQdVC4qC0qs
Sok4HvukiJzCwX6A0DTZZBQ3sOXBfTSAAtA+IO7Cln67npWEUqXxqxOuyf2lN49U
Svj0XbDjgfS4ZhHcLYOZcTi+bYW+2yqP7kVjXtPxb+bmPWS+bSJy7/PR663c1E0l
BRXvwmQYQ6VfA+QMZIhOgNaBPwAuNpOd2Xb2I8FXFHHDCnQXuLBpuqanCc+kI3M7
fbzf+4AQqiYlfDQoM6JUS7vMcRqMz8MPBTDGlKGE5HFpGS+PN8YO1V+W4c4q5EgO
s5fwGqTwMWr8XhuVdlW3EDkBAJ7LspSKmUBDf6wLCISAuVOIZXcbtypqZSpQb4pw
JocKwzfdC/XKPvA2pcx6uUE4ldh/Lakev9JXkWYOaR8PPoLeTirZrl970PDAxG/B
jL4LXXV9sd9PQuCrHNZWob/1cNWLaZNLBg5u9Kf7t19NPrO+WjqUK5v55d3sCDLC
GOeSLblt977P4bP0jYSQHjjY35i8nzLwhS1v13AnF4z8AbPV82tgm7jR0QIvrOuN
J5tONkXTmxqI3Otz9txsqjFIhM7acoITZT/XlOezgaCxZl+ZAPVnxn8XMeGAU2op
hJTChjYO0j6wRRvh6JHcnmU01joCbys80N1XnVjXvjgC3S4vPATp9+TygkiFOyLv
AgvlFjKKyQOsK4vvEwX8IxhNMmB6YJWcEuWoWBWXz0ZQZdoVF+ckx7RxGl4LCYn/
Z+rW3ZCHwgC57NdvSCLt+QfwQhjDI1DoiIxa6l6Rs0BS6d1j010su1R4MFY1NAtX
XXqbOjuwqmmzhgTU+T4jls/kCyoo6ujequhQquFM33L8VA1xXny9cMTcHesTmndk
rcWn554BpRwGa6gK/7AnqW1lQPQXUL+x/sjLKdu56tYVdJMJwwC+dJ/NrCfLR46s
fMPcSn4B4i3eLPRtC7Ux94uFr4ruBsba84AkrP/TdW/1m3vM2NggF1lYeYyQbIQ3
BVdn2i7vNX5K3bSB83EE0dhs0ucVfdLU++jeFZqUt/ic3eG2qAfwGzKlsqcoSYvZ
9KM1gp9khGfQL6VcQHmWHbJ3hiBVjoM09IzwDFFBlu+o2vGb/YEviVjhVGU0xsjV
v9RQgPz2tg7eNjEPjC2njECMQ83dbwaHUAvF13ycNZGeBN4nS5I1PSpHqGBIIpkM
+A28IUkau1k85lJwgt3vPvi7FwHXzF1gnkNnAoOcELrm/VcvJkQ/K9hGy3dEdaO5
zLZvdN7wFrQH/TBwu6pgXDWDeaOhSVAOi4G5ev/3f6RNyqIYrgw7u+pAVhGiQBtC
barXWwLs1JXEYzm2OPrg5uNamJjy0QlQNMsT/LuI1PIZ8BqtUw46Vq5jz9FWUslG
/sVFpFBt1oMVbd7Q7JWCC2Ce0p0wnTRM5sfkd8JPws3wUFm5qiCBLWOjIKKEmFT/
vBtfo7zYao6mbDc8eKMMDE2J7f8VGsXVZYTUcZlM8BIJBjaU02ruLhzkX9cBwOPj
hl4HMux8zm2KJAzw2yt6lznwJCeme/00Ipr2mVxAIrimRQmsmWfsWbXDS9LEDe1R
CZKLz5qEjRgyb7O3rYZnAiIlP1FoH4i0CdqCBClIEaM+BFC8kbjBnC/36zWrwVP8
XbyazSEmTYf99Sb1lKneNfRSngn511ep8gc2AX2XMpRgrqv06aorrvn9qklnhsC4
HX3WnPijwUgI+xGyUv8btIM28MQLJ73MG0dvVKQFgr/6wQsVWaoPNaRtTFLo7D0Z
Be7LLOLTkV+Gpdi+2bQoycxKo3DoWBBSWZkMAyzufGxi4MSfnNVpU8cpDgru1Mck
djzKYQGZY/DJTqqkROuzUzILKUfHa50e4GSQf5Y97h0kY7VU4d1SOoAdcI3yTKUF
lqRm3+BWnTaLATYrDjp2Xcdiq3A/IXq2sWJWe4cg5sHSImsuKgQtv8m2byvBqWRR
xUl661i+lSHr1ki3gsEQGOtrENOjqubIx0sRhItSsl8gVv2NiImyg7gWaP6+9i/U
kjxGseGcJIKFCdn+jQAaqPxsjOgLZUI5s9cPJbDrOUX6tio7oy7676BmPUnZIq8r
32SrDLiuDFNuArIqxylfdPV26KUncLTdugM2MVlGMXx+axAyOg6QMJnWb9KDoAwd
7qgY3owIwNGXyr6rNHbidvsphoywN1OYugGgWFJ/Wt4In6fgouoP+qntigisoRID
jazqQB4Qp5XoVtOtdZK2oDCJpcEgWz5S5d9PoQw6JJPbSsBvXMfCAq5Q0K3wgmbe
VIt4hrZ/RxWUX+zojSZHK8IkcTVlyO1WDQJ7voVCy5rxBBzqxYIpxv5RtY9OpwiU
d+MpwFWaLJHol55a43tXnATI10xJ1std6kQetVHQciO0gWW4hcxinL+qO7U6oUpj
14Uch0YDdq7AHbUo7Et/zSKe/AfTcr5bYbIGT9z36l1xUAJUUaMtglItpRM7PYx2
eYIx0/BV+C563fSdfI8+27WKcgoOoEhPS/Zu4Re8hL4j0ZLa1SIP8FGWqLcsH96Q
KeRGP4hV0pKwm+KvwJqMEbLSQEx+KV1Q+I4d9YPkGJ3wq4yAVzCuySUKD47PJAqD
vSSTlvCUk3IFjn33si/pF6CrfFrplNIPtJRSsTsiUXlEMPG6R5UCumydoQK4V9x1
zEbgy6L59HUaM+akvnxnScKOqRIHN45JlYc1VvZhuaRJXG15SbJTy9HA5HDcYoYH
vd7pEWsQiRO9IHoETMDp0Ve9E52rAjAUsq7XGfg6OxpU71go5soxvlhTBh+Ufukc
hRvAIG+RBAC0AYshX+D/AEX6Vkpmx+hjcR+kM3TT4u5IHz7cYiWHW/DQEzD1opxR
MRoJXtVK2pH7nXSzI6eeK3m3t8qgKgEQO4gQVL80DIvTs7s3CJ/3XlBQ4gHVndWY
FTUg6S6eZkBSTKtn/+78tjtnNJp1EnxO6mkMQ/X+Bhx/HqPKHqyI/k+jFUW55vHY
ZGnHCZRux5VtUeRdwf0f6MqQ7r7GR9874UxtMNJ5sbFQMyl3y+s9JcrOZr1SzYjG
R5ahqmWkElGcbuNOyX3llawDh2GkZJ9wlMS9BtSt2RRw+Zo2RAQoAnan0frIv1cW
aWvJiCNRvrclO7i0cBBOCasd+wAUwjlLW3iFikUS85TyydjjL9xwOZLPT/zDeemQ
B/vSfI4PnjyVpG7jmx+rbjXjRG0rhMPrurUJO5zK07dJx2HbPqGPGdl0gepfWReT
0CKNc52cN2JtoWnGTxusc9DOnWaHGNuOQrqPhYMwOC95Tcc9E4EFd4P0zepn5VV0
5wpU/UkTO4pDeRcR6+yt6Us9/ude5HeG0wjkIghpzmcWDfkWZb5Yv3XYjcuvHK/n
Ls/cSHnGiL9FArYB6g8MJ+Kz5Sqy0qdR/7c+wpCk2CwK/eiaqxFRiiBmv9z228wb
9220Gff87gaQYw6sDtNx7NAed/m6xBtxUK8HAsl0Mw4WJdqLuHlyqnAp0YLDLTx+
YcOb1tnOhryMwsmtsYrZDZCodYtf4bNJE6bkjS5DPBv6VHfDNHaqpU2hEkkUktll
TuTcoREpBstLfJHIF3ohxKxON2JdGSKeF700j75Be82y7s3jP984Xb8onYGIAt5K
TVLVEqZdBVdNPrlEq24j1UZNMZzL+6QPZQKtVTTlIuIsVeho96hcpZ8gjXd2jRTo
lLEyqhDLnkbZIzDn96EmFwMHqbO0fRl+Nrx9e9zHc2Pyo2ajJnX5eQxcUfgKbk1h
iuTlIyoHErypb3y8p/IsipJeidhnYzscqkjzv5tJpfSiTqHSu9orRnFmOyIHKQ59
slHWNVhEYE5GlEFTK7gwpvR3l2Rf0ffycCR+tFbwad75KFnpzcrftbPoPcLRPjfl
cXi2lmUHT/7bSWn+4PMC6tvOO7admqD5ll0ECFFucmujAkuIOz04Eyi8tlXiW9Df
qwHNC7u6xZ7jXOAMXtprTVy5I/W3+YReTpKQauNIEmvGhHZoS1k+a8051Ixx+uc2
1J97HCbV/XKGHNfnQGkyRfFapGKA4LTUsFwqj52PsIgGMUVV8+oC39cGnja62MVW
cvUCshP7to95arzq0xDVfFKq8jVhs70IJvnpfbWiYCE5okEMbagk24Vn6yZJGPBE
elFFFEHF+k3Z3qiQ4+y9yF/odj79dUZPVwOeZGlefoxB2TMinFmWvbYZumzjzvfe
iVbukNG0P47aOX6aormYGHb6Rc66m+eTo6ah6EgQKIFW9dP+SMQnk3140F2pBZmv
A7rnKcVYh9oEGD9oYDUZIVFc1BTQns8TWgF3p1MCWaojn6abTf75ob5MoKIKnGH2
HBRJ/5taEYu8bJPRRZh7prRd8rSRdmp+OXyn5oJOJdxM0G10zdhyEPyWlpgSu04H
gCBlchD8Zh1yQ88OIrrl4J15Bf2xtFKnDDQf/FZhhT5sQl9n+OP2N1CNjTrYue3g
P5wtrQCzoLASn2VS62AmHyF6LabpRQJM5Y8+KyWIhX6n+u5OZsgx2Mox/tAqtPtz
aRwN4oWJ6+r+Kurk2P25MMQZUflL7MLW8beKoZ9W/Y8M9MXiLI/Um+RKPsIoirRy
Wp3VT6F40P6WRFcODLmKJinpIuJGWbCP263TdTa3GcIaRsvsbCFpZOGos2SZVwBY
4+dh1RFKgc3vvZD1VrsVC/ddFjzVDILfRQiNkCn6w7nugMEQmYAQPADZ6OpuSPPG
8orLE/2Yk67D1Oa+aG2Krr9XcqMwdbHrSp6vZP73lNRkzSdNzoRsxeLqsKEcr+Zk
R9sV8JMAhHCbtaZhOXFM35kMeCaIO3RmcEjTJIVY34Zz94TvaSR/KUBcpG80JhBs
DodBWA+eGsPckHt3D2M6aj59pMlw1oXr6XKzy5mBcrvUbbrOB+6JMPjp7gbh/eA7
E0Z3Tl2oLNvKHyvjEw+Pise4txRfEPiCaemrBG0s6CqEiCQ93I/1vmyTnNugmmyn
DqNP4XlZw6nyuUWTxu/WFnb0pioRO2hIcpA/NaPmrHTiwLwG9uXJgDeGXmxXZTFd
LZxuVHabQUciLQhPPxWomWxuLsiQfWdBWnGD4cFsiZyloT5S81DmebYlH+9/TpSz
JuxdDntagy2OSxZbRO9H5Mq/8IFS2BkxwjdRSEomqXocY8qPu6EwHm2ih9BuZGeI
FbWrgFNy+Cw8yvHPANzKZN4UYty4JC27CDzcnjSMOKXhM5plUVS1QBZUBv+x81XE
izaSxxOkRmpvEP3a4ieyChtY9Ku4z+WgvzGgIjzd836YJPeIqyk+T6no9sKqT3+6
mnLQe0/sfwW4Nje0o0q4ZZLczNLGos7LpRx6n9iNuBEfYOkOpJRk0uJ6L1puZq3u
0SZ+lHbhuu9m4FDg/fpcvpyNpYt3VyhetI0YCz7AmVFiHkbWkpDhAuOmFYVdlj6N
DA9j5lXLP0ajOPQccqAJ5iyOT/Po+TG86ocT3xoL7eTGEKGaNe4lQqfMePnW2Ny3
JB7oZ8pay6/q9DontDRRfyw0ZmhGYgmw3ik2tgINsNC/Exv4aWwz+bVEV5Uy+8xy
TqFbSQXbgYxTig5/YTzfW4O7GwsbdZ/2X47Htu2VsScbJFBTM/R1letPxJK4GnNT
uXO49ld5KJwUfquLldrdVaESjMsfSFk/C3LQHhuKx7YN7JiWF+KYrtnNjxDT7uI5
ysn8pfaHFGeV35Sm0Q7fmUT1UkD0e82/YxdHVDCwYx0sUljvWryOZuuaSkVyCULC
dAwLeeRb81JPmxGWclNnw4JFsxCPI5fCsobC4o72DRCXFALh5tm1CF9LVwrOPE7a
ozkU1/Y7Vy1ZYowIG+R10i8smKL+KNG4o6iMY39bl/EFZQoDu5RFHH4IFGYpDyjC
nbPKbyl3ViUL4KSO53QJUQcHqOeAZ7rRpU5lbnGeraFadzCBFQ3iD/lHc0yG3Wlg
wXdQbQ3d2oNtqIup8NDQjwT3znEXNY3UhJfkEZC0edeylw5hr2VoWGtfIIC2Hj+M
JeTQPoigR7YyZO6l1W2friV0O0tk7o7UXNmghOXfmj1quqoDX9RZ9FKCDlSM3TeA
wSbdLqT/KKOjOw4bUudhYrM3ayqpqZrGunWIxTfpNSsAkeXJyAjVqh6WjXpul1IP
/NeerEMimAZSWDKd+sFd3JtJSv0L1/aUK7FpgL4heDRuBW2feHsNnmc6qiyAb0m2
k9s/m7TGXYmT/wNBoqOhPiowcvT3GuqAr5Cxb76c7M1DIpLl37vHXebJdM+qgHqk
3s1eCbCzg1kJovzjjoCl6NgGkO7XvCNCmaNL5HvO4UmlqMZSgtzoTh0lNeUUDKO8
rjwpW/DKcipfdrYqo+Il2Orcpp0V7JKbKcGO7vhOhJ9JyZSjadN6lOrWDpmDCurd
H+hEm8VN7ooRhtijzEYsqmrOJi7nu8TEtMdskL2uCQtWEyXXZLniqk+UyLSQsRAd
eVYvoO1SlBpBfpNouD+l6v2Ttu49zYLgBBWLBC9sc3p617IjvhFQJrujvYGhcHMg
BpRiQw3ugskXYWxap09tMq5PAonSeC384lbJ37/VOgmDKtdFD0mQlmrmyqOJGVzX
kbfDqXuz2DYE+8RTOaohRgbKx0D6SumCbUsYObCINqUqaw97eQ6UiwF8r8agw4oL
faweRQKurlaEvENP8A6j2X+GW6irHrEErUfcfCfIFEEVKtf/U2NkYrvVv7Ga/r04
0eQOc2R+loSBY/NqFI9VbbtsgrxckhjU06khnaT0e3cGzV7EG8PpW8Un4+JgJnsx
RU2l97xO4nhStfAntH+tbcC7O/vcD1WzfHIRNbsryvavGbN6lFZzdZsLgRhTgBFX
b5KfePYgNUz9z7p5xEY4RsmoqrTI8YvUCoL29n3QgdFgxq5rZ2bZgGUz7rXkwZYE
Y1n96ql/pXqd78YedwcPMjrJwjaEY/L3qZ2pdgz8SioZ+pGhGs7R8dxITXZk0JEf
EVsXUBA6bCsWjQRtmM+0enNYGNgu9aol+busijufnRupBw2AhGK1nizYqrJeeqva
v6+aA+T8kMziUCs1A5VlKLnVGZvlxpAjJqalg+GUTit4NFIrRFbV1+YtKQxeXHZ6
ij0sxWo0o2nPkBtA0Sf2H2tTmmh7D6iI1qO8EiEN95DuIFEq/Cj0viAg/R/Y5Hqf
O+StQBcTbSvVCQ51wmtYCgLCn0NOvfl48fQiAsCbXWwe4A3c4dpMlRofNDQCZhJU
DyUtde8ZoET5YuohiAf956M3OCifI0y944KutDXKQTS/RHf/zFyUWvhWMQrOdeL3
SM9jcMz8wLd3yMh1wxSOL5U4mdmzdGiPoys8yYZOPhHmdmVK3vf6z6lZlhzoYGjY
mb+KZNRgOtVqyItRM4lnFeTXjf6kmK0NqxG2i9johS/qEPyUrl4qhLuKj7Ccl5qT
pAXVtS2+iaX6cQCwhh2e4DToZ7+l+YDyG5+NG9rD/UESrMa5XOBJjrCrCu0tajTY
esHP94KutY/dF9KIkIEXq4Db99DzeipQxa70qyORiG5+I6QvYiX/Z9BuqEXS09+N
A09U2JQixlAdoQ1beK/W9r9U5tgG07Mppz1dwH9ifr4nVuVpwW1YT50hL+e7lp9p
NjHLhk/SEHoAvP6pAdK40CnLqJA6QXglzOxmvY4zUaLO9eXkptVULa8AHzd62i83
g6Ya4KRGCxMgfYyChRjaa3iBd5yGxFc59GGiMt/Tq7hA0wToR/mYKJe5ViFpkiAx
MNtdL9NyFcqZaLFZDv7nu2RZt5nI+EQpYGKPlU5qio9BMaU4hYeNg67rRqHwJBSo
GgVjAb/be1orfycPHN87CJoR8BuoBvDgpePjfxjEdLW9aNdqgm5qpjTn9Sbug/+w
NW+D//T++F7qLIAnZSjv6uEAtq/h8yc0OuysZjuMDR43NfrvB+JwSwZgTe2XiMpx
2X1/2i9PBTsMoYaqu3b/bIwvLu/ozEIHdibFpWJVdYKjQov8DnwTZunLcomGGWw1
/pwV3pgQVY/+gDrE9BVG5narPOjYtiyv9EKyiNhmyK/Evs2wBX2Geream0PzQvan
RfHhzi4kmvIvUpHCNB/KK8aw/Q7N/KFEhlpq1mFdPZJ4Xeut/Fw760n5XltQeiwD
pKxja1CiBRanvOhyZ16qJBisnr/Klg3W/hqO46AJngLivY2CV8hVS4C6qogkFOF+
cVYdUBST/R4AhsvaAOz+T3UIYO3rnk0wv8PhDeSVFvZqUw+JQbKm9tCcuSdbt0wO
xGN7gRUHq9JmYNZy0JrSe30P2tGwYh9Lnno8jNCtAtTnmHXKo4HkmJkCBxIUZ/Ql
d/vHWe6CBwkrou5W6TeudOisHnzTb53ZidGE++hhKjOW3vC8AcNvfmEV8kYEGz61
ouvVTRxrkP0yKkLYynImYhR+BYILf3PWYeQeQRHSygkjq3/GAkyxenbtccjBkmOY
vlwmUK1ymDPrA00HAbwMZrUN4ZJSPow5rkwBES5u96ZAN9xZFqwvtWJuiL4CFxWR
jwuhl5IYHPnyO2lPbpE/+Gr3PXS651dAwKHolIOhm8fmLKxOfJJftsyyEiMFagwZ
7p345Vle94Vvw9rqjWAW2CuDWWG9zP2m+b2Ou+k69Wnu41o8qHWP0mYVL2oKtM7B
6kUkfxr/edtzhQyfeBhOFtORAjsQ/pkKFAMQKnuDmdhcxpd9Rg20jHUuDrMKjn68
JHvphWrfq0gtqOomPQGrJ8rQtZu62F3Wx5JOR89g0bsBqlte4iShoKt/gqOZdkMT
mp+caIl0eZR+kkj20ndLwSVfsACCwGNwdnMezCG+1i7JCoFVyr4KSR9B5EN6aJrf
sDzC4JXoPhV4Kbbst0Kuf/OHb2G0h+wS1VkCgSwLjT0mlI2H6LxTGdGBpeHiy08u
8ecYUzpB2js4gc4uCqsIhAnKiYzQtvWCYBSkj0QwQhibNOSRBUxlvcrtpxQibOvj
vPJnCX5O8ImMydAV7VPxIrkoIW1axzJy6g+eg+Ri2EuI60u+Zf13pLUtnPUUkFXl
bZ9KfCYOUj2D9eAfHmSZi/mhv3BZMUgfsYapIDo/5on8iyyLfpYRcrdMk6t29zNE
MYsdcJbPl0XNoayMz1zUAwiCtbQwV+pgUaavn4v0aP4i9od1PB+AwxVZjmFpiqpg
4Tq5XZepTy86bkmlDyXTXKEV6yaP4TbI7Y8Y8esmAs0AciPM52ccb6tg27xC/+h2
3QOkYbxkVAKQA0N/50+/FCjuueAtLOIJl6dsl1Py48xOaYtHLe+7lVO1y0B7WDKN
jHgqYQMxgcBwa5mWYlZV+nQPdsCKW3dcZ886Qnjm3AZvVCnsvAavA7e7LlExGc2j
wyLG/I87KAV7Ib2Sx5f4kS4YfD2RoA5VcWZjq9gXUp8xkyNQtAvnVPD9jqG6zE1R
w6b9IA2hRiB/F2uvPL2jvm/lPu9KPhn7cPmFSotOUi2gJmEOYfnx66BbzjGHsclJ
L8bXdypCmX6EOM2fFE8abpJ3E7vDrobSTXVuNF7i8aCwlYnAjJFYFjZBidYOIp24
LuVwSLblXzQFDqlPFLfhhUA8Ll4craS1e0X++YfeJKrZGPYAhtzUYCVhlFEN1WKt
3ebzfT3Wp8PWtJd0QUT4pM9+tpPD+0TGoWyW94jTbIET84zi4+CNt2x+qPOEx6Gn
eEMNC8AZIHGXVLnrjHN8EmvYSqZgGR6YuPKklCAr6pLtFbNP2uzby7YPNabLJZHy
B2BTqMqB/YbIFoObfDEFJBqq6A0beIsVERnLZYPadIPfc8aANyEMRp2Km9vanOka
6ymB+N4DH5v9gHnOd7BVa0kUi5BoYzIJcFkfBPXFJi/NlYijh5D0ouUQ2QbGtz8g
UwHzg3fflXs3OKlz3yhmU50/YrCkxk3gIe4jzPRtxJ3AqHpSXwJCJC8OAFWcyWHm
nGd2gkgroTvrRsrg+LFOZxdTxMESTahvQuXnADrmSaXIIZxQ7jK1THLQwReSR37d
++4fFaXSIcRdkDEqGuHJVdHR4Tu4EX/LHeVGDtK2hCebCvIRsbAA9Fl8J6uZuIq3
O+xPgtOvLrys8vVguKDpJJPzFYSmK0fb3c6TOhxIL6knHXf+8Ray0mlCCdA/Zn4i
WOn7gdCRdoCQTHwZaBAP4EUPQV9gq+lLlu8MyUYlqBSTiFqwadip3p40Xcv+bSyS
TjiKGPJaruHQZRusI29veGYoFynjxndJufzn5kUxydd1m/i8UomujFO6spU7GPJ0
fMHsZ/oSzXraYcm7B/WimUCJ/hdl8KLSamtYi8JM408o5gAZ6e/JAQwzbfgOSwAR
7LeACnTpSpv0UdX+32DOk3cJcMbOTsHpXR7pA+DH38+EpVgjK1hm3Wp7n5QJHUu8
ZsZgQBUvzR8ZcFYcCsO6k5YyHrlNu1v6Phy5D54DUguSM8KLicAvXjWkGyyd2qW0
ABBF6ASAdZWo6f55QGnbHlF5tkZW/YPFcup3RpFbcC1gdD9BQ3Qyaa6fhAqJLKKc
N3LnCPiM2sCMoaPE44BbtDcYXjMOHVa4if0VjLFpKLzHWFAG1SdKhqD5lFkdnFPm
BVJ0ob0yt94EwwXClD/GTNez57rizG93ayhT9MiCZHJmL6J8S+fN0AqFJZMzQ55J
7b9BaMnSCojP3afhRwzaZXKgVtyNbMXvnLFItrYrnSUhCy8kYtA53t2vaDkDjU1K
S5HvZdF5qBh5MmvrITUh75plY0kHzKJ+chWu3TavzpWgAdoxhmObrlga6Ceijcqx
6PXA1Eq6yriM/5IRMl1CyjMLYnKM3Uf9ouGGOLVECbeHQWK2A4d8g+4pBTmu5uJA
1REEci75r7ldGT+P29F2OR4St6CpBgmiepwZxl23LHd2CRxdnPJA3DzA2JWz8VW5
hAiSck+V9+HovEuAeY4ZrROIKEBYOnFWcVWJNeHgLe24lbPta421w6+PmJp4LtuR
V1DVQVnw8kYzrWlgRCB79PMIlv1cNjFfUtcrbRZIIAC4uUoKDeu61W/+oeQRK4wz
0kcQq2g/zHF59WRQohxuAUJqVMEUqoBsvGEd8Cpn8kEsE2Cx9PaZL/qtdgL9Gn0s
sAPsUmuFAI4eJEMVQopZDLUHixR8Yp/Po/ElatbHOxRk2llJO/zIYey83bt2PCJl
T5fo2LuF6q60hifWedtzZ5uj72/8vI9z5lpDYVJJZtBPUVKAQeUgI4ZQNmXgoz3E
WqjC2PbXSOvLHK4QdnpZg1zm2Jim4CR2j8YOk0+9gWmUZL0eDoMPo5bAOxVGN62/
5/xFJfMGSKwyL/kfyFDEDWLPYEW4TaVA1yBxsN2tpSmfG57cvRWq0jZ/rpRWQAK/
j8DwSoN9/+DDJmhNcJHxcp1vUOrviGWdo3umkmss9JBMnxW72IiE9XVGyyPFzgMX
3Vssga/7m/6+juSqRPhDTNowEMFt99cEJCGwG05bgKZwqJhaQ5QfWc+dIC8ES4cp
fNlEoLAHEMHxXrsL4gzIkEgfXEigfJFlPwYpwgOcxdj7bF5QnPmI6eddu2aoIlHv
CTbSmfG6grBDkbw+eSeG/M/WFZl4f1Q+q4/x2ZlXW99paxssKOAbHLa+0hGQKZA5
JqeUEpCZgDlmtAHkogpX/ztpchCL0nHSE7QrIJZHJlmWrX9ZICkUIbjUoSbNtGuC
Xy68XWZRZyPCjcuPXpIWnIA/NYgbsde7cn0wa6cw1zdL0v1Qr7HCizka0oMSqtsM
0EEKWSqp/t7rBAYPm1IS44cRIKxng3BS3Ia+jbe52QZy1BCOB2yIvKEq4VE5My2P
SzfUlxw6KZ1lc310xxAzZdF+nTzN/y9Yc20bg51nfUpffLx6AX68oQq2h4tBLQp8
4JkSMosoIkTx7cecKxgKy19z+LhdMkWZXeEkEyzFxzm+xc0lDu9OTLANjtamTrF1
qaYePfT+oD+oGHV7/ZnJqPwD6UfgkwlAL6cnlWKH2KAXZFxDPAkYzydUk3qWeMaF
Z7yftzMZEnksX5AFLFm9MHe5L3pf+xKpoYRIk3UiBL84sWqOuHDr6dOO2nVUjJnE
3Fwt7inKb63BxqRxpQKCpU+MNplQPDDxouHV9hrec1tx7Kazv3fXW+pFglJsCDO9
oPg8IVlMFvXLcn2YOuuON36yNKAQU2yVvy9MO6wBaBHIJOeguH7i7vNutboZzXQb
2E/e5H6swaar06uFge9B2ZehP86oyuwze8aRAyzM1Mkr+hT6VQMkWxVsIbWsQBSU
ns0GuQ2RWRvdaOrrreE6LiVXJHoeQkh9Exc5IUep7rVwoqZvT7dHoIzIsS0Og4sd
sI+MJDDgz5qXOZ87cZsl1XGSh9YWZDqORnbyX/WEA0tI3hDGhLQ/h0GABB/qXH48
WG36bYiqv16/KCHteoQC1+Xo3KCjAfy3nyfrPtIzEimxnr+jGuAcu7Lb/HEpubtK
RfiAp5GzFAb4lPBhweSTwuA+NSr2qSBeFIwbRG0dW6ELa6PYoAUNPIWHKzY1lI/j
xA1yyyRUyLsi1fe01VFQm/xk2O4a2B4Kezf6GwT97CBdBO3RM0fE4aSs9/Eh6iwZ
2uLc5WEIm0Qoo2I9W0pxXZRVctLQvrzwS29azi/SRYQa7r1UXlAfuVEea+GFCwjy
nhjNxoQ3awWPtiN+zvJ5ZesgiOp9/s2l9FzKTi5Otf+GZuaKygQQwCoq+8KsRT9p
3zvix6K44ff56WBr78zvNsrzmXaZfh0OF2hr/uYOtRuZYadV00q3ELvFzeeC8FSe
9lS6L5wF3uydWja0BjKpDdcm96oExWj65jQvNzdSMGH0lKVfY2wOQQIy7rz2yDiD
NaFcdK93dKVDBW870M9iq5Ib7T+sxk8FN7i54+rJwG40rRHZ3F9OFh/wtnNSav4o
AdVWB7idqktWo24cwdOpu9FI/gXwgkbPvvJv8PP4Cway01s7gdt0d2ZeLoT3ueCT
slgPzZzrZVCcjafSJNFfDeSVVZ7WhzKs8Lkkv21JOLsbB0iCQCFlLoXZpWBuec2E
aL1dpjhWGY/rnD/hC9VGHOBOvjfbmEt4lSAVOWdePyIT5JfJ+DwggQta330h33KJ
tcMp9fpTX1b6z6U9M9OYNEnceDgR9akOlKAyC1gO/KQmALEERdLXTXeqD1SktOeb
QNZHjWZo+LLysey7iq4TvyoE/0PqLE82nh9f1CF904AUnqNneVXRnR6t62tO1j79
kaUCIiBG+y95S6aDuNtZpU46N1jy1eXV3zeqmMP08cM5xhD5+PbMf+l4rfsFO5FO
QtY7IDzrlYN/91Z7huPPrK3I/qTQjVyn9L5t4MglL/oYpMtuOoLH00C+leA4Q0lt
q5wRhyZ7wmEcUtSuTbXhGJnbSpaNp79a5y4/E7CriZ14iiTE4LutnJ5SV3Igo75O
+fyzXmsmMi7gJDww/8ocPfOpaBGBez34jlZiaSY2Bo1CNbAOhNuqg/ieOpDewcaj
r7mcXmvZSWOuzlHtgvjbKIEw/36xGumRQYy9nJ/UcS6y0/L7hsGR/7w97q5qhxU7
XPm2Yw16/N2vMFL4EEIAepgoD38Y3YD5nDSgQxKiYXhFUuglpfuAR9R+s5hvg97O
0yDOhEvmu3/rFE7n44enrWBbYHluG6KOFiWgpvzsZ7jd5Obl6KVWDegfIABJ5AnM
zJo9PvZ/obDcZYiSAjLwxL33RyL1O9zzQVb/u68zrknnaIPGXl96fy9scrDsAMed
d/BNqI2YVZmlxnNp0pz198ahoeIc/1ao0zrISxuk5Gd4ZRYe7kB4PLs7yLEA7tiO
NDu4rg0Caf6YyxEZ57YC4SZ6LJBljPNyyHgMjbIiO9xAiV2A/u64jHsI+oCGP17u
FgG71Q472HLIhvwa9aj/2cxPH0Sk7vlUTZ/S1EqgadgX9lXkFmo9KcN4TA3Ykohm
kaU0//nQ6bHi3OFzYoerlxtADDgslw9dzMY8GDLV9oxpluz4O6zOrls20UbyYnGF
OikvLO6Keu7Id6KkMfTi7pP2+CMJ43hiEjUqSOY9+4/oyqQ2OXJzu7+O19PaQYhH
yHdHJwV8YVdURCmj83SfhGdLi9kB9LCjLmqJGh5dXdV6q7XyRJbJ2/YxHexMxPfJ
I/xeEVZ9WARrvJS5aD/QXkTqfKRpsevYm0h5aKnwzjAImDydE5lkewsKpQvDCi+j
mZwlS38xVmvvVtB03hop0jtTJHvvTN1b/m6nxNa3c/Ud3F+DO711Nr3J9OC+y3bq
BDUroMOdjlRPLrEuSHpPC1pZs7seKQQo6EBFlXSEtjAUU7As7RQXNZ4xBEctxllF
QzEJeRIBXow7eQ+MCWxCBgN9r9pz6n4UIfNXOOyiSpKD6TyP71EYu5tOstuwhysN
6jp/kctbDE7o04KT9zLCfvN7xlGHCf4UkjAYR/ednVdedZfA+YBzSjROJTYIbdBG
vpSA4Sp+icnOgJN6EUg+gkV5E6AZFxPd7HrbUCtk4My6nzOFoMXl79e3IrbIgsb0
XyWcCOP+P+qPYW4lY7vobOjRGBSmOHo7nN9zeD9hEAYahQcxy/t83EtcHUkSH70P
BvTm9c24GbjZr0hUbe8u71n9Xqy3qp/iWoHEURwuAM2uwkatvp6YdjJ1qt3LGo5w
3qV0TKhBeUoS0g0/9d6JaEk/d7R6Y3iu0Tp6e9Ty7ONWe+AQNKgBnFTkemUGSZL6
lNepoGI0nPD/yot0cjF16oaY5JH5WMqW8CrOj8t1IDoDoBaq7Dc/zQS+zwN+zbUZ
GNe7r2jq2cAwgLEVwoEWJ2LrJch5CmPHWTqxee7JZQLQe7zPbbDiVTSwhwsLTeTQ
4gA4ezwR7m8YwajjNY2uy1VOhf3ymYeKOTsEAmBA4Eu9We9eRA5zdOFNePJCogUx
wRxTI5F+57YaXI2g8UB6AyjwGzkxtILs1euiKYelHapU6aux8Rk2eg7OJIsXGDt5
sfMVgZFFjmKrV4iTuRzj1iWKK/i7G9ssMfGgP0FktYzAlLqlqF3OQZ5j6gL9Q8yi
s0xKGjd+fIi9HAavMbKa4windqaLCkmHE/90/8aPKARg2AmOS82ceDhC57CtC4rN
RSbcWwFQByz85+0aEzhEOehi/mz+Igr4MdbPAaA/nc3KIVH3E7zMeNyzWujksjSJ
HNt4Ep6IdZ7sbA7JZZRU8HuSpY7z8D3WyTWz5vYSa0mCR9trIZ5itbO5g7Es4GIU
9XRvhg9te4QcH8TZ2C1A6Ka9oBgrxI1d1Pu74Zi5xqJkMJbKKkqjC4zPxSgHPnq9
8A1S7vUyE6FXJ1VFzmfngtVQUKVBtcilaJxNYI1e1ONpVAXCDN4IB1Pdp3ShuPuS
czAfg7qzHSt+dpuoJSBnHMJL1Y3/UgyNhwWlgGGsNcWup+UUMoAtkPLkBjU9MJe4
4EOpaX7x+wT1rEx+bmsOng0lmoC37K47QyUtHyTfM8pPQ5MistsEiM2JFxNI+Lrg
Q/GAlLzS/rq8VlJ6jsFBa70UoIjt0gP/95iDCIQTf3CaDwweW64JZQ3L/JUAXELG
EpbOo0a9AcXAwpgTOVZT26riEIQW6tZNrdvDtwPpasu8CA2PGrwxsFYFqfANpk2t
oUFxTdiDC9i12/bf1aG2RC+pfuw/A+8cagJuyomOxqQg0joM6XiIb/iuw4RKta6u
BBpmpPo+VQS38IBow7ReuvB59dfowc4D/rEyM1lovzjIwY4ZwBdlS1ieGmYSsoeR
tpSYIhXdmkIr5kcTaicdioLlC8M2ViJgaZWfb+P3IVtqB0qD0Ets2FoJ/Sd2wA34
+Osv+gY4y5eIcdcMM7bM/L8p4+FpcjeZ18FFyhvtk/yZqJXiJxLpCtzp1YaDkr8L
T99uCBVosbyP/xnxU8YKYSi+WVKpXcimfPxylj7eNyZHTr82lLJAfO1z3HPEEcQm
OCuy+/6MZf2vtiuuoDiaAbs2IObIaRrPhAlpNlrkzlQPND6kuYSfTJMUKnbJnoIc
1vMe9xENhTEPFQ7yQ71ZfXqvlgTQTLGxJzH81NqpYz/FCAoL0EbjQzFC//WOxc+y
uebpbIEdsGV1cT9cn05kSigPhlRy3FFTUP/jhF2zsR0GJUMANqWOwB+UTB2nyxja
RdQInvG+fRMVZFISPTbUDtMdSFPIkg+FVCU1dZ5k/IKd6sCysEbXTv5yt7tJzS4F
pDoNi5JdajUQO9JqbygZs2k50ZoKflotl0OaXIoj4a57SUDuYfOE+qrxnOzoDbfH
aKNV0rd/Q8j0GzE/OP94TmoUaI1XwX7CTHKa6onsAERlBSY6g24bywE8jRZnzltE
ZRP4aui67vCkEYfjsrbJZotrSgTaDrl55nH9kAYVz/b5f6THaNPqtX3kwS6H6BTH
BVXXjL8/zhVG9Z5o6zCGycnP5nRqF9ozsTZWisi7VmPQedivrPgFA7xDNqXKsZzu
DY0TMDAMANu5PDqnJbOlQ+wGS3PmV0TridT89l+vdzsVyCP8yCvbDTWa5ZB1hzoZ
g75Cs+zIB4kRvp85Bs6UIbe3eD/qBXFfDNAydc7D+E5EHIFAjzf9e2GFs5gzBQHR
lcVfs4dWA8OCD6j0UY5XAeMp7zVy4O+Nelpc5VRE52pcGJhp9OcXa9TaypRivrCC
zG2sAl4BZipL5rh39FoskXnYZNd0bsi+WEl+4nkB4oMxD8oNvjm/KMm9YUt2s1CW
fwTVdgC0hBx+cKehJDS2JIMvw07Usr0FDjlhf4sDdOm78PT3E6SPIcEsF6pkrmh7
lLq+3pUdsF+x3UTcfuT1FKeUhVA6jP7X/4ZTuAPfiilw8KSGkSoSdlq4O8/X8R4/
uUIo11in5eICrPytOaAKWbAcyy9XG8uVzljBFL+vy2bZIzvfUUcPhktumzCvQOqw
d2lPOfiurCGUD0gICQ8lo5F/HoHG2PuyolVVN2Iux4W+/07a6vi5j+cIBGuJFkhC
Y+3g/7uk84UMT91iwS+g3wYT2dNRtPPePh3T0RNwRQ9LS3iVpMbGZ+ESRvHFVDct
3ybQVBgLtBJyBm30CAFu24kPoD1chBErBOLITj73EQg/tO6OGZc/JHauekhYbHkT
irsuwo0bi8qfrOIBsj+wh/gUEm6M5cRUwKs8lv0X5cR2Zp496CRstS24hCWW+4B7
4cx5UScCwbgIUYEW/eMA1zSy1ygl4DmFZdSE5mtWXsWF69PswIC9B94oBXH/qGN0
RyfrcDQUKOeA5+S2gkxDZRsBQHWxY4bw37bf/QOTKELEgz51vbXnI9rOKCq2qsdA
a0tNm1H4NwU2nlNNTMjdw08GN6Ce/S+A4MGmf4+cfHihHAf4A0ARbNrRpiyj9igK
CtvH3K25JkkfJW8PF9GLxglOZDDnkrniXNJ9T+BfMPVYspLp2FYsMylAhhkucCdb
jwl+hFAGbHM4I0A1oK9gAfJEct0vdhVTnZ/BmQ208jPAxhxFdhX9o7eSQfl/5OWO
um+MbqBdZ3Fp1GhZT1AZa7jijhSHAwo+S5uexMwOYJZq6dOB/UnHZz7E9lDOggKU
tWRjrPiHBDq1ER4GnG+OSmtPOuiNR3GOB0P1ooCplKDqE9m1GKfwSYxxJ5GW1A7h
hDuKfOjeszFr2Xf/USGLrlCBpXDJ4szyDgkilnAi/AmOv56pDhEW4lddqnEwnr6J
YurYDZ3+eBpZZ9/jqbgH4DDliW4JT1PUcxYMU4KzIkWc3BF+wzZS0TGBlSPGxlMK
5PUCkep99W7sey3xs40Gp/cHnsclBVpjagJv1mOraVIAIxDBvTE8lLMlhrjeHHzi
rMUmmNDSKOUTBUz24jKEerw1UQCWPX0mhbLJQo7SVJAWAsL6JxlVG6fWVzhH46KO
SDyH+IX/XDFZSVnQTDA3WihiQgfcxnkGYpzmLzfyX2QPAu5M6SvhG1tO/MDL1K+9
7752Iq4J0Uy9PzIw+E3DGiQ1CehNJRor5/gBJmgQBGhpsmxi7UNP+dgFYdLbggTc
I2jaw2lY9ppG/bmxSMKHrfDtDFj7uXWX0K9mRKVKub5gQwQmVigBHmNINYluxMHm
UrXlZjsEEdTcZFk3rrZL/u0URAmmQwzt2fAYvaixll5m67HxeKOsAkVkdEELkimS
fec85vQLfZO60AU3TRnLdS0ECvlFmTeJHV8MR25/IMtfSCwqQpAJaucBavbiJVY3
vJljGwW1D69beLiK+KxOSw7VcP/o2gLFySMPIXK3gM2NTURleRfAwLiiztQQFePz
jJ4zL7JV4ZLaTvnYWV855ZiyWiKLUEQjeglK2l/k5NTr2QjwWoemBpdNmZMe6yvc
L1s6/+KEmxuCYg9vG80Onvd22bMgYiiP9C61WpY1ZY/le2HoVbj6+1lA/ifSl6eU
P3CktA5j2ZMdyMEkyZQAuqy/9Ce6oawcmM/ruWiTwMEobTwHKU7G0RWgsgF92h11
PRoQmOpdz4qPInK0GOTOg7ohkjEY5VdPWdA6sRoEqI9ZDujA1SGzLnYZcsWcf4mh
ZpkeztHgQXfdGTx32gD1GwF7xKPBb8rVFEbhr5ZQ6YIbfTsBBZ1Amnt775Rpbf9Z
wVvQs6FTVnaMbY4AXf9bWKLVARm7KbxvOXyJlpcoKhcBi36oBjCT3i9SyxIDwkdO
+Y/2FIwuHDwbD3v6NKgW7dwR17k9NrSD3XhCOhnaSIJIR1nnSdXOTIiP2pxQ4CzJ
mzUaqMAqkeGkCS5Vh5pJMrav7FQFNzgZ0ZDIbToDc7AZ/1pWQ1itXOpxpOlXeScE
vmPSrezpvT3viaYTDVDQa3I05V/Np/+Hx8izM+C/94BOmlmQJiP8OoTFB2CNGtJ8
ZS5S8uu7KJH/ru++FoHAxm2pH3PhsIrfCz05DMq/jn6gsYHZiaqjWy75XCeVsxr5
aPRzcmry2BAEXGJkeVwbiDMmWI0rKbxQXE4wiBfSnTeCj1soEiKuNaMCANVvtwoj
2YzCnYYoX0Mn/PCgUX5u2XX2aUgAjXbWkC/N9dt3R8IsJjcct475Tcd5nrEAy52s
7+CsTp629qN9qs2kiBQ8h8zVZlPoTBvCPHVmJmA/CpcFYRkGldlZLqGlHEUd5QCA
HXfbp11AQEKM5NLG8gSi3dAi8cRXvUPGn+i/dwckualeQIXHndpU28sL8GpaG8SV
R/tv/6tvEkim6eAshYtKRfsblkqdKJUN3OnSPJGC4UuG/P9J390MfQvCeJV6CETE
fC6Mlwl05AwIXgd6jIhE4Zi8RRiiyU5pxEWHlFAt5oCpulFkx2dbP2ar+kUe+VDZ
scto6OhnTQupAB53OC+pMzX5JJ9TfIDWDe6NW8nWcx0IPuyg1D/7YeczPd2+3P7L
zreffJxM44yh/ko1uCovufn7uyDaPJwSIMi83HG1/xRA9h9St2ksvQbviybSm99q
1wOh4X31mSlB4rvfbFVRZkCCice5JJREYx044jg6hR7FENVf3ffY5EIlaiz4qrQj
LyV9Dxmmg7rBjPgFpsTCR7OgOaqlol4lzhBueKpi22OwCmHCdo+ik/sKeojOtgYw
IscEdIpJckfzxxwv53ENO8BfRz/Tubucecb3RxuhlSsDzPIV8v8hVXrTGy8/98EU
jGNq3b4dB8uRnO1GNjX6w55bHd4p+AA5zhLzSkUWuN3mqd+M0Blxb3n1lcovYNC5
weJ9brZVM8OC2T7NGRvV/NStf/IZO/hSVfIpNjtiZbmGzH5fC0Ip8DrdfGYmz30U
x6oSrGAWipOL1IkF1KUGC4+bCk+dSKdrkibaMTuybar4lG3iH5H5FwPpitQVjinG
UdkjCiN34IAqZdZU7ZCcwDu3tqemneIvjlKeSWe0IE9h2HXtOlAPGlmUtmRzSieq
liAxxp2oSQH6YhRddOxedyjlzdD9PE8q0GoD58dv3r2DZ1dcBxqbHAemrv400/qW
sP0HjmmkizOmdUWeU0oeZ73WsqWs/Nl82y01bzkTTf+5zQJs8nmwCMZC3JWlKUkI
0shlEI1ucw24le5w5VfX8BQdHhPCK1MZahmV0/nIqDlZBA8X9ZqTMkrGl77izu79
g2ZETkaHG9x/OhH2VWLTB/05j5x02fgJA7un+6DVclx9Xv3rZJ7W4WBcyr5udqNN
dW+T5w3DPWYuIAyyzOM6fsDC1W51XvNM4PDXl5VHzSEbHA8bq/adnX7CuRoQNbV9
oTiYm40C2rNUNblL1CQ5XRpYRTxIB/i5AMrYu5Cm/vXdL/VjN5FfTF0PLwILrB61
7lrIe7RcCftmLXTUlPOaVNV3DhQNE5QqDJSyJ0P/U0Mdn1G4qo/5LSk1TkzQ0aPZ
vqMHga4QtpkFdyOW9Pl6Z37KyvtgRJFIr8A/yK3Gd7ISDa5nXq06E5/YyK38XDr/
cIWO5A5N8r8/P4aDpNIT9cDdVH2/YUDVFgwBB+fy1SRKkxgLY/zizGL1/HuHglet
f2CYl4utj2TS6zE5+kn2Ylt4+7/0zkihV29fKVfMvWMzQoTI/6WJGIX/ZTHSqYXl
6H5qBfcpQj4giVN/3tCWpxQBcME8GUKdY+ltkbdCJ4LvS8IKrJexYU5ssxtlsB1c
czTxMdzPGlPZAfNNCLyaB/5uWdCJpXQh1YxGvwzYpVbnfU/GwtdaCW43TGThFW6z
TmTMy+21xin1vKF3KZbl1ZnEurQR6203ZaCfaI0eAk7464uq1WRBeT07vcJZfjjs
CjubZoRR6kLeeeqOGfNq5iP6OG8Ko0snyrP8o75BaoWg+va19LB5ARyK+fOI68VP
+bUpELP2oArI9v8Ck+42Ecu3u8JBeE2Q+n+YklU+aMFjwn9X2fpZd+IgDR1lwXxj
8tBtiICRtZ+ZBOXyk+A9+9Ql/LBFTv66fKwX88iSnDYSIp2XqPP5ZEs5qq9l0Qza
/NBNQvQXVGuaqVcYAM9xDZOZlp4z+R7garP8dr5kxHTIRrMElrDuwoZ+83DwGNSX
q1TMimnEwt5cLGSwHx0nwRbapEvqKIfp44/URBH7kJu4/F2P8RCBuoL/6WjfbIzA
ei9gu/uW0VqJPG6vd2WH3o2eQYD8JcSSiP24OGf0kcUcpdThwiJ4PNhywIE6N8QZ
s4bm3Gcl9FNVW+AUXVx5+yvctdZL+PxGAqDO/poujXAHAtY6n08Aq4+26dQzCDRu
1KCalnq1E6Y6HujDS5Io/0w6HKWU12XanzM/5dag7QX5Y0mLwR/8KM7WvwL2n0Sj
Z6SHw93ozH9Qcr6P2P5+1PZspE7GoW9mO3HWwVVjPpZ0ETBdRj0pyvoyXGjMhEls
b+rcfkrQS6KCTLX8bNateUW3eyM9zVv5IggX58R0faf3R4AdjOUgYRSrgw4BgBPK
UfL5B975eqRzveoWbV3L0+moPzL2RkVQVmha/8Nrr1jjktqHUI8alj3yhnrXPj33
tbJ8MVlvfSkVrNdU3i+4C44M7VdC3262f2NWGaa6wAThizVKTPE1RW7EMbWvWSYS
bgChnLER6K+i2U5A9NdHtq487UMNNfsTs422LrfaGyyr4C8sLwo6MNfYDV1wIx8h
quJcmFBR3HGQdwY3Fbt+bmP7Gc6UDoMzK1rWBGJa6Rg++EoKXTGjq3ChqYbVxyAJ
puYESh5vLpATm6GN8ujkC8srAtlwXF5cnYKQeNiQk6QEH8vRM3mrdsW72LyVHa0u
8r0SReUFdl0ulgyKvfRAQZz3bHeDZl0Vy2vXaQuOUL/qmewV/7RqqZjdsMKPPUBB
wkEtvPUXuOuXqI1uQRmULOgh/jO/b4KYG1pnDc1pmYDGzQircJAjorYdFkncA6+4
gmUsLraXbzbbfkkqKq5jjFdRgDYNrVoH3WbG7VWHx9Ol0qA/ou0OCCM/Ym7QHc8C
6/tDyGqb23ZRI4CBRREjfjviGE94GY4yhs2MGGmGn8tO4DvpRHIUxdNMJr+J6iCz
V68aSdx+Pg6F61gf7payI21gFB3gWb1vnThUIDRbAA7V4BTw+zBa4SZiJ70pT2oF
fhESajiv7YLm5T50ofk4WltwVQNbE2oayYwpsD2Pska3njcI1jposGor4mGrfG6G
k+P2qEr9u/nND7rV7AVYgXB0RMIg2VuMUDeMKYp3/4j0m9kVXYQ9UPN7htL8QUum
HLFHJpMP4RZ2NJpHaQSYV9qNkbBz12LaZwu8OjlPgB8XC3wdvObXD0Jz7OqBOeC/
oBO+J7jE8Bs3qVDR4/HEljkHQ3qbblf9/IvX6wDzokUDXtH7YXtVxu/yRy0lvlB6
sqSV8BWYfBsiArnptVf3+dLQUD5IeQ2fXA1EHfQZynpj5Wlq38ZeLxoCjdZYKeOq
y/jGsX3gkWqi0eT36I3e8wQSmuy3KHKXC9TNMpisAw5XIoseVXY5OLgKC/ZxcVcu
KhVxQ75ygHoR59Mk1UXFZo5EU8I5LglSO8i3IdEjp/g0IUL0QoXYt3SxOxqJWwRB
gYpjMES9n98dCmmDlaNnkL9Izuj7K1HI2eEfCJhiSM2UMBlJ/Fs7Fm6EB6tzBXRx
8LWLEK1rtmC/WOzE5v2fF7uZR3Ik1Q0Q6VKjy+xTtWjR03PI8yYY9w22LDei0byP
KdRZNlmFv+uu7R4oa1Y7A6RqluBiFDwW6rZEF/cSMmuQRQgVTT+IMYBNnQVrOmiO
trgJip4NMxovp93+Brav7GAnTrwzcioWut3pbthkAx7+TDgq7bO+21OmX7PM3sqU
hWtOX+pMiRr0dPyiIpPn7FR75IeQ+woQv4qFDJHL4HTK6E8dh5Lx+60ANfcb6beU
pCGaIepHOJCzb7h3fiw4Wi07gnej7/St+8j60xCDYBBwlV2VPRMUI9cyEGt29S4v
+rUv/rmIyLlZ4bf9L4mYLnpqIYjo2O3xorESi57Fi7Y2snKyR5p6Ec9ognaSn0pn
Ol3cEL2UwZqrzyG8jcx6mn1aa2QG/HrOw1nspihl7d+pl6CeuvtQ2gGjkCJevWX+
WhZ1av2vKqI+fSTY+ftAkt3fHCZYOJ+0+lN2hTZUVBDbnbB2qZMyHUv5aYQRBgut
16dPLG3qg8Q6eHqbpq1VCqBY6RZ9LQKk6RCqtYl0sVIqGlradYcwttjYCwN4gaqF
XqRjHFbYK0abUDEl9sfeilFCwFkmuhx8xrec8koz9whxukxCdKUHNfDAxVUjGjbt
Lh14AP/3VFPqwQG0oelD1CWPnc7ZTrJhb2tU+/jyT7aCfI4ZTm1Nukxees1fqMi7
d18F1kLmKTiJ9q6iiMrhUBQPT3AKjxRRD4dwa1UDPb7rPJYy4CS047FJhMCq/A8V
ZMclqk3EbaOEl0gS6JpB6NYbVS1v8Rd1vieZYzqUDZ9ZQffYasSC0FIJuIfO9o7D
zFIceYItkIJTLcKxQWl1hieygG5WDhEOAjNwS4TFUaiunyev0WxUcrbvhE2bbhhy
nMq8xEFtbeCiBEc+uD72ToFKXrU7PuqqNFFrJd2xUmwRi16TSuvYrY8voyoeWwp0
3wDVvCvkl1ZeVxohKjbwnMNovjk9xGeB2u/6L1jSHtV+NYjcCFFsrHNIFnlcYATg
za2O6BQPWzA4vRvY8ydBd2ZiXhq1to007QJl8yhylDltH2afKnuEky+BtS1mMDeW
sVsDxuUSwL3Sq2XrtMYDTXpvceK3DKxs/gP8RiNneOKejrPafbhVIjUvVdv2D8G7
eE/3U+30oo1tHME9dXjgjIQZScM6TzgXAc7jisllpadx3X4VjKXbIx34dR3a6FgL
u5zqI8rnriL9FWSImEhANFIn98ymBB6gW+wlWnPBBut5Hmll1wrr1gztDDEDjgzR
r0BlvuwA71fRvq692DZZTRcOYg+8LZwGftE1e9s5LpU7ocPDK29eWSSrJVEqJ8Sc
sGOlnSiD1P/UAm2degncF429w69HGl6IalGqRVKvqHBWoYXFR3PgQpIbvWmEvxRP
R4VUtYsCFXv3pc4o7YVJx7HNpfq7VUs62iqRZMOGq9BqQXlCiqrPEnX27QDfQMr+
Bgn4rVYAtni7iHDDdNimfPobLLGfAlJooufEHhJygi2XRmkKrAqgazQG65UogwlD
h7Us45ZBkm1KLV4IDpsUDfrbqo2fTkdCZstpXTgSSbB0sqgKs/pqPdJUGpFeEkhA
KUj4IMtuFk/jqkaB2ifWWKleoNIlVdi7t3KPA1clPh6IY+ghJZo6w8q4t/dTo+wz
HCNo/bMk1LzwT1r/XQuahXlMRNl/s43AMDd/yivxpY3TNUxMvWIqSaV4EUdkPHtU
tSC+z72iW5/JffqXX5mAYnbxM5ZTvrMZOkBYavI43CObEJekBT3a9d+L1Y17L5Cc
jP7QpJueoApwuj9k38yKGm+T2v2nijuZNRRyJYAuOJq1EQ0i8jj4HHck7YKyjrhf
CXS2VhptGbOnN+qNaj02v79FD3/tIPAkJwi7kyG/AuV+Ed5/TSNfRjdQI2gAef+o
MGxAkCBNHt5xmgAUSkLSF95VcjXEzwzPVA0DUhc73s4qR2j9PI2oNMVue8AqTgx1
kwXEfQ4M2fUqm5iQcKk6TaGe1AqMvY3VTgrfb2M0PP6MCuEMdChR9wnaVGQS9vox
YeyoTVNCYueikBpAiNDakPPV05rCR3OZkZ5iYr9M3Mu88CPwxbsFkrrgY6q0cjVN
cyHFINs5JJU059sCpYLteC6C435+3+NtcpBchSq9gmJ7RoRg/l1yC+MIV7bK2S2H
lpc+WbHzE/QNPLfUN9kgEjYyyPHSp6286exlwwK5lwRrOFtLp9SBWqupsO99eCFU
QOahigvoHVYbdna+nhsRWEHcDkcZ5DH/0WX6MOtefaT5tWJY7jk/0IVR5yt71kX2
hDP+evztmbZ/Ieb7uZzxWe14QVWxa2I64UOtZKaQdQUERONM1mQjne3FZfZycBfV
PHk/IaI3aISYn1lZiaO6BvJ6GmgqiNjYg5pg1OgO03RwMLEOrmR0WsJGFnu/q8IL
fFDCwgvxb0QVCHzUyiXgZYLWaSeCIov7IA6l4ctHwgWTE6iFs0c+aLjFdXSRqMaE
Tr0+IP+0DyWHOMtcXl43L4HhrhzhZEY+kCQfiOXcerNZ2asg0Y1zFd6zGXmLZoIy
YItKUKHr0IB1KUUF0yxd4SlWfJvttucKFZfRZ6rBIGjUYslAjMObFGUb51yXqWDK
DT7xEHBuq3wKreumcKoBR1DwPRsVwJuTSGpzeicywWOjMdOq+cw5hTUpp6ow5kUk
oFavR15h6hpreGbmEVVTfNVrJJrU2Pnr7J3rVg6dMDnJeF3CsU26hMC9utZ7ZABU
9T9Foot6hg1dPChqUwSIgHDGbHfPJR2B2LhV+G1lIH8KQBedWbfBhKtZFr0YvKib
MiFyRmOH81dqYxbYK/oefusv4nQwtp2H6JfDdjgvMcIm1+1ZJihGOZxpKHryKZXk
xdffb22ICU0/RHgZAwH3bxJQhQI2kuQ5bztyK7iOJH24cvfR5gAnZmWQjtrvp4eu
cGbGQnV+lWpfRjMWo2ufipeuObSDX7aRv0bAOp91F1rSNjjP0BMcngWFZxto0cM5
PojfYtXaE5XLPhIdvmwAtHpibuDQqAjzuikQrF47hv9PFeU5He3aetqI/DEstE3J
Fv0BfvCSr4KiQL+zIBa9WA4sG/53fQEP808SleSA3fpCSD0SRaDEh+Ihujrf7KG0
lBJQlFeHEVrBHaFdeiMXH8myVacxApqJWEfkfhfeQZqUIjgXH4cXPicyp5oZciy2
NR0c/YDk4P5EFTJUTeUcqk3whjKqn/14qdYEus4txofes2ZZfef2bspwAzowkvu5
KacqRjXxwA/h4gF2qPypzI5KWQWvu/OTxzbVZtIuuB3vrh4xAjhva6bhQAa2upha
T26gAudtTq5wPYsaPZQsUil0kXcJOTI5lurcZ8krHpa1N4Hjg10WLasHKwmZ7rMS
gTNsrru782ssTS7Grr28dIqEnnSMRYf4AAFhzqI1idYIv1IfTQyxCNQIZKyi2NXC
XzRLl0LmJZCz5FAO9EX83cpm3OM3orUvFjUnJp6sr+hDHZZaW6oEO9cCs9OpuQx6
JijfBzrigXkuVKqBIXQ/goX3YMBwgjVA9wpycaQ8Ra58nwEEUt2S8UmZ3pHmlcLg
ZZIPZbtYS/+vaCUHT4T/Nyqikrpenk+VAsLlpZwo3FmU8ixBB7Q2pTL3g5AAk8B9
48IZrgjR9LN/gYzT1f5X3IGuW4fK39Lv+3mPw/GbOkIabKkvwjPeeZJRadhndYQM
hQXjf798eXA9Y5XzfE2dI2wQlFde82NuWGiZRQ5Dz6ZfFTN+iZz6CUSMBMXdXi1y
I7uA1pZEn1/4hcTuIJ7bgs21Dt52x6P58Yfs9sOVNRdxklLmrIVR/Ej+JVoF+IXp
zb6G7sQd3Y0opVq4EP6WppCv28XMys0J0K/CUNA2G5lVpO62VT3P979DXN5Fzuru
yLySY7alurVIpof9h3G+URENUGwNqVaQyFy0wFdfk+qHGhCeG4ltedY4mX485wWb
zhQo0EJgP+byLwdPL9W4P4oG7pkqak4qEGcmHHdFh8m2/W4yS/zFTLnc0ez598Xi
9aENIb2El28uJIAEL1Nn76Oc+MwlhEfKWI2bXS1o0jrt4BsSe2nXy/nDXPaoiSMb
QrIZBL7q/21+YET5+o5fX3oNZv/A/RthGLYqmyd0BPimfSZvkm9svzhsH9t9URPP
4Jar6L1m34TAsXdXKxlxE9BrAkfpFH0g1S9MGncLQJ6RwpKBpNCDe890+hjpYtLy
Cy/5RkiwSkBM2+dr/GAjt22u3Fvp+HW3kzfqXiYsGTu+swVutAxK+sYNkBjXqPPf
Uxus306mICbwIkRbFIzAw+5Be5gviI2vo/UHdq61bsDz3Amn/GpkJ3Xz9LJJKbn7
K6HAsUuhwLO36foeebZ+q7SOSuIk10bqLml9PUZMZNewrRvKQW3JZKwquERD4pdR
tYHwEhQQ0x7fJ/rhjkueuYXIQ4/2fywvVRRX5xtuLwlMCeaBRjj/Tvc4zXJmZNDZ
yw8RthkWz6iQ7ZEsuhdmJJaD5ozuzW/Qca0j1qMD7zhgz2Tppa5UaZFqtqLu1HEV
CKPETCRHKxevjDZIvzJApzDDWARsGHCsGZ3bj9zTbXJSXdrWEbPAxNePlwyeml39
k+xfelneN9opxq7SJ580pzfuLPB0KPgjT2zD1xjBOQPvokwGoGU/7o1Q7mYPR/mU
QE0ojN4Yq4LvIfIAQGSSEiUVa/1Xv+E7aE7xl0uiHBsM07ouOhh02mYihphPnSo3
UmEl6A+G080eXygqTfq77/9+AjV2b5OtnzgKzd1g3TA6oyL0FSHiqjKdXOFOZsgO
lT7gzSxqj/26yQIVBuHi5rjtCYfk4ccJqid5FHo5vFzM0Q8YMcP09fhdWpFh6cZn
j87Mh6UzSfO6jWlJpqp1R0tA9WNCOkTQjwRAIlOsB/FuIQpAphSGv9RMhyqchRzP
sLg3VlzwHNHrJAvrGx+SMWsNbpnyJFAXHql9tQbSFpjfCDy8xZqGGb6KwCua0smI
QhxROx/3lbzY4mzJzLGdQD3Vm+sRrJi/CdJSktGQhyJzlO2txLRCKOR+xwQTxnNI
mG75PPCkdJcKVqMgHqQs8Sz5Dw7H2Dj8FGcMugdVQK6u3z3CKQlVAE+6MuBVwDcT
4bwWVHEtxnPm6zJs1dBPUrRDYoRkzMxbyPTYVeuU8o/yYcyykU/OUrg1YbVB8mPR
8Zu2j833YYY8K42kdfy0u0nufCotabk8vd4nnPi9IPqpEgJdvsxP+PICyhUNDS3c
f9Jq/Mov2/yLPv+012tDb7PwSKO8ZvmdCtNc/XXV+FnXrrNkGDwvPIuYNynSbzId
HGZUewkc5mu4rK7GIbgjRHmVNBT5tl/CEbQ+aAYpbsPjAFKno3BB0VcBdkjD9cz3
wHbELARZaA1bDhGsxHIFVv6525/ws7Bc+4rhUy5wUyOuscQsBAprYxZuyqt1PHkB
5DcqeSOQMOus/C6/NPNiSkftyANh/ypnKs/437iHYiyJY7ZatVfUE7fZlEdKYAip
i8vSlmZXAJustjdfgzds+gspnIL5mWz3QxnCDCKYk8kH41pOhrj60Z1LHOIC27wK
x0wij+iUnrjK9v0QRxPKP1H7mJ9hJLgTqZhMEFmYSP5yvXuHVRuqqi4e+BUV8Oax
Uqoty0GKY0QS+GBbm1WBcCU+7wRF98vtmLcl1wEzW+9gZY7eN4zuf3t5F4JIZykw
1u88HsOR3gyC3GOeuNKtq5TeBv3fjMc5k5oT5DTnTF55h0Rd1VIT5l9Gxc0fYWkP
p3YwiOwGPvZ5SIU32BDVLMRBInwWr2BGRjNHolg94wr9CJhwaUx1z9JVw21UcKSN
bP2PAdQceGq+sHxC6wURLQGz5L/M4KHAQkAnSCJIleRmXrWta9XRqx4YhJJ7ucov
w6Pk0i4yCvGTGTL5QU9/qp9ocUuBitUNPdHuWPT4yyF0UZH0Cd2WaDt/RXC/s43J
x6C7ykiAAMcl+uAG+XCOJQZA/cOCtZIqYS/czA0kW7mI7sItAiPRC2716hfoa8Lr
43X54RZFTCDkySJ2ZZAPwR7yGv+ihtfwXjKQJ5IeT/n8xzNGlY8rpqzQVf2mndO1
kV+yXK1CRJ3ie4sFHr6Kpqc3eHDxadsfHDVBwlFWHj7y9tnVizPAj1FiTPY3bRc/
HWDnrRajDVWEs48dMXqhVyLTVvaC5UqnSEaBLqcwe9DOjONpQamlQ4vbYJ2XRR1O
WlBxu7j2msMcl0aFIkRbrFai2kb8w2M7myk7bN1UWKSPzQ9V6wDgmgi2qasr7WtN
inZV0IcHYa5F00bWljdLbOmXhaaq7qROeVcdJY/Wj3LPflNQlli5tpthl2eofLaX
rIp8Ym/TOVxO+LF4k/3TXppr2HwU+2SZr8/fTmFuo3gYHX+o1zD2Jv+X+4UWUkd0
hgbRJDrcDoi/rxHjmpJAg0G6MeLrcESOmi3UQtlYBjb1T7ejiF3Njh20Pd1xH13p
B6Lz7YvmgKYOjGsCDyxPeAFkydvooVtEfa3pqXPYUP7xYAXmeTXWdN0+fK6CbS7Z
KTsRr0S3RM3b6CFSLjRJ31CmEqgdOWITHHsiLCsidKEaRhg+D5m5DS/BLErmtwen
t+0OG8zLmjoX/ZUEotFuLsSW3/BB3jkBHNZPZhHTIQQZsehdz4b3XcvFsoZmZk7P
3uEb2IMTqBbpZJ2hUOXPIhIrMpbX2QzwfcBGjLWvt8wxPVB44hFrHco675dT0EA4
tVuDXxQZ+h5O/1SxDpKT0s4K7MrHT35eqJvdxSIYv/C45tbPt41tjOc3/BlctL2F
9cHzJx314xjC92RhWN4gzyh+HOL+V2LgN0KUmcFl+1h03imRBQcfcTta+yu4Er2H
ZJ/7ayiVvfjKo1c/DjABo2TWUJcp54juJC5iErusIr4eVVFCWEcTwSUreFwJccDK
OvtMVbkj96yQ+LlT9jBPw3Oz6+Z/QkxDzhgW5Zs0X1ruW2bJ7287j/MGCN3P4TLa
1OlaK53MkW6+vevg5t2OAVlTCAESAI2X26nBM8EydorKWyDSec7PNnkAL545ydfW
18OFFXlvcNpYI2YH+ZwRDJtJ6ZQSdVnryQJsejQqmmBGrS8DH+QxzdB0vGlPW1vG
QXEO14meBO6S3lGmDaZh5u9wPBBP9DnvSzewBVzlhtPqz4G5h0dSfobteYtKXcrG
/7qwy29rbhYtUbScAbkaPLiPRAAmmzxF9nc1kqrgwBqSG5lKhA6+H5/7ANTRnfW9
d6MBwgI1HTuPlB0FaR2T2tHmtASq1mCkRtH0Yw7wU+FioUji3qmOmcQ8FNnqi7PI
PD/91g0oSkvEf5rTY+BxQBgE7krqatxiWT47sTSMmxehSQwL46ndfIvgS3LYatcJ
lBNzgFMiMg2GB8JhJrH2aameaUsPikSZV886AOy+F83sVbO5IRtRVhJvSwKnukFl
cPb59HfeDRUXtIbv7NyaKW7dYSTIElwW0/58VQO4DQLuMOBnv5ued0zUzxNiP2fk
fAFlttDVbzkUJf6XsiYumdo2j/K0NpCKgqh4zSt8JRz7kfK1dQ43M6xPWjBAVp93
7aCn0hAtN0pkLl0zffC3f2p0WPXFSfnCOua4GEEQ66QvGDYRHual34rgpKneynOq
2eTxRYQY45YCFf7oMPQXPPTfBeZIvYlLd9DutccyphYlTKcBbrvTsZ/0XOJplJ1b
KfmFAqO0liJQV9+URwWIfVLtgNPTQ1UH0WHHMVLR9mIMaCxbx2wqEMZ8q9ATuHuc
qiaR6MbYvQeU1TZBLwMPVNr9m2nKy/rEx2Fq4b/w+FFepc5+RP2SOLpd5b0j1Zwc
mE62U8WJWomz5MRfhb7YbDGEQrNqFKlsYn2psWB3ddXQkh5ZJapPRcG4GEoQQ6WA
vShFWaWWeWd39mqk/5XkLyvhy6+UQKGqgxq0+NViESXw+Ou7LPqm5ROb0uRd/Us7
AY7Hyi0mDJN7LRNXKK+5PDKyVZMVVnEwd0xuVQABdrTIT7nYtf+NPC69mX7GwWma
0IhvLGOeT2puka5CU3k9/CLLgQVip4hOkUgq0RVoKbFPh2YeISft3WvbanJed2fR
GeEGwG0dIJrlbQ/xFzYrmCgvueYWS5CBmoOeJfPIyLp9IBHBs2C8JXx/rdVymU5s
w1wo6D2JZAsNR3QnuyQK1R4wTxo9Se0ut6gQFxX7RJjPFnLTJ1q/z/W5ggcY66k5
U3T8TFI2jGjL4/dL7oWILVXipxlL/KMCQZWGe05OdbllofF6Gu4qW5Xb6mTACPhl
6trInV+/dHAEruycuMMQOVoDlpLGaGPblHADvYifTnyFdVxxD5RimJ/D9iYTkLMj
yTl/i6TBdvd8mMHO6sTVray5BSogbirjKAAfcRVujgFv2l1ua0GNWefbRbo0zPLA
es8JbpgBzrinYJ7lgI2FMra6P+w4qpx6JLK8boUakp04Kr4IN8F8N9x9rVVhHQ9e
Qz+Ir9D6Cc4kADh7jbo64acO2fAjgJYgHQDyZu+sjgRA73/TNFIFDCwxiD5rk0Vm
QrfiHz5jI62HoEgC2FsNOru764Ookil7N447ZEFtvqfiR2XCmM78HM78klk+eWdP
vTk0me/JIsRXEgEaMtIr+1SfeF/DW9x9nWW1owa1L65GLAtQua6Gxfd/7kh6wRfZ
YN7tgGxOIp2Sj9ZdKBlAU6AzZabJ3E9VZCntVDH7pewDXRxlTct0qoSDnLrnos79
nTwntEGYjEwR7LS6R7Nu5iDqAQZfz1HszskOTmYFZqvMJ7rnOYCgxe/vpjnAD95N
y72ik25uUn2slPSrTf80GSNmyLxuhvYsB0A21UGec49FEItpl9M7wtbo/Gm2eEK8
nhGYzKTew7k6ir1SWEkCALHbloFVjvKygbYLuKyr3N4ijYyVq4+EsxLUTd+xy+/V
PeYkaV4cR59XzMvgo1A4zbqTGw1XNQjqm08vWX88KGh3D6Y9yKJburjjikqmQsRo
SdMJY14Lmxa50vdbLOr2TiFRiYL3XMQrfQTnmsN2Z64/qWCkuJdAammBDc8uy2rK
rjAXCdnPnjpKqgLD5cEJEN/dfgBEGsa3sGWFMBg9Fkuz+48tm6Pc9MYDps5WkPm8
RooVirKs90xG4vkVIc8dWeivl+yTVHw9Lfz4xTr/qjZ2d0ZlgUN/4Qk3Fd2Vz5S7
MRDILKXhb8WXi6IlSmAzjeElE2/gfBDUaqYEBD2Marl9a+iyBin2G9aJpFxs2KAr
IGQdWCyDi39joaZpkbWRDKNd0ijZg5T28srgwNs6m2NiRb11pW5cbwx4u50Ud7fh
ZZUTMEdu6olx9CD/MjmZIjURoF8AMHJeF2K199kWnF7GoTpLFL3GXuSgFqJ2nwAv
nk5aNI5oZp7n/ZMYncaDqkheqzLa6aNgQ7BjrRA9ivEfphDW7vDt9xsSGfc7uRmK
Fxg08RYVBp8NqeBUCAnWeKFFvr3TMiU7yKNF5hroSKLgnrYtrJJ6eJoENpgwcGG+
FmPpIAQsY83nndx8CbEauBVagd3jUgW/Z36YEChkwyjPynGdpZjsPzNUOBrhxJ43
NxWqzz0CscZDQYrRssaIUfe3YdNaEPdlpa3HjiWTGIyZYKqNFopgKErWsbn7ivsp
IpriHsBcqDlQsmlpCjIpi2LRKTzS1dBh6ka/7W9Nki6DX0O2vuttyJki9gKQ0iQh
qsEWrK35tR31obKac4xyvseotyRiH2dp2cjrRtkq99EL1/dYCdrqXAPFNAV/irJh
dVwFkzFU/GnnlyBkt3OlJpR2WeGwz51iQU7Zbea/caeAJTuSif6ioEek6rv2LS/p
2smngmSvdrYGqWHl6o08jVmOtDpT1FZqWOmebeb5VKuAOzAcJvbwPQAN5XgAu+T6
PGy1drSmwmNWbUPhc3eEIyIoDJiNroP95TgqpKo/8HAWEG3OB1BLFwjP3kPwH+at
8cl4O/eNng0R/prQIug7lhQAccEmPzzJAR/Y8jTcNOUICqNrFpEJtaCBqEY43z6I
aZ8TazGFXVqVGo+H/ZJffcSsvXOcfvQGGmmwprfa1G12YGvKxSWXwpOgVHNTf9MT
It7tBN9e6//PZkgFrJYavDdUDs7Czh34o5oRLjfoMJQy94mCpGt1gNjmYnOS8G45
gPJYeCEF6VDYhLLXXvRGujzb+PiLsY0HYyXzW2itrhuC6Uzp5rvsUKiTkwwBV2kj
YMyd7genvcFoMESMs4k/8bhG3xyXszYa4Il6X0ZZnMRgKyboFLaR/HVHLtVXZGPn
nq9wJ0dVn4quu1e4qVoK8cN/rXbUuefyL0YsiCewXTRWaziYIU1ABzsMSUD2V6Ji
yjjDIw0cl75EWGtomPP13EuQSxJLTaruCyDnzGMxUfyZecdkzjzZ9/GAADhA24rQ
YVirgcNBOzcQmb9YoqQBBp3P6rstT58W1GNvSFqm4DjyIy97DqppvZuAfpCxM7Eb
gVNKUfXUUd4vIDpf/SYR02aTkqT6HRZRTDN0HLjAJPY+4mUpghnO6WX3dMbSPIfQ
MVxIoR/CL4j3R3EdkDRo4t+kCPUAL+8TjMdf6Iyk8nIIEbsWcT2FsfFEe/5SXjMf
Ro37prLzuebqI33kHJTJjASEc88t2d3OmDFSVS+iZ4ANT4SOsVNGYF9NdldWPxoG
2fm6i3aVvD96ILn+jgmoOUMwRSvG+8e+8ygXVHX7ZfOsziLttfi82a15ZADAzErM
Yeq/mcRhqXHbOd5IevNcVei00RSpFkgRPuA9UxTIU2HJ0s6aC1kEan5nAyeoWswr
jetMBkyPamsZZaX2bWqGX/guueCVXnMTt/N94E4l5Yey6ws3P3pWtUYNqrv/dvAf
aoz5SzboXfnmnbmhRQ8ChvX9GaZoTj5kBy/zoRQYFo0gshDxP4oDe5sQAJrC7BoG
obiV455qLoEGAa2JoJxgZoDPHvKbBjA7IVzybgPfs6LIpA2Xn9Jb1gEJq5l5SbDV
1YOx1Ay/rJCTGpIkVLMq2IxW4UOLDZr8NNTlqSFwpF1i+0DxLoTpUoOLEFNkKUf+
ml771gUQcsUWfj33r9Pvxq2T+Sr2QiiJKA7ng6cchdQIt5IYLb+23h8zUERZ6bWV
6myqmDottZTEz7lsbUfntNfHwzRcZAUSiOYjyQsZGYW9ZrTFz/OuGmfPqhLY4SOb
MxGN6TMyRLTINy/Gwmno2fQtSupf5cyNJqNDFt+95UIhrgeEeEI5i0SCn+4Orm0V
`pragma protect end_protected
