// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:02:17 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
C9tCy0Rp23bNfxpdb0p213i6UaDPU8eHUoRYNssSSCSSxQaTWc56ZfTleGK1MRWB
TOK5kX9pWhRX0ft3qC8gQPIUMOZu4NmrPnX0BL6VEssU1+bLRNWDnVjTPDt8vYR6
+C+cVKiYfY3gSp+20/EoYm6IglaG8JSF1TH8/iHOqmA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 180752)
zPEXyKbm+3+SDCY9EEyVrh+7Za6Si2UwaC+fwgdsIxNpipwyGHK6mvgfnM7bJWqS
b9nvYxxZRERQQUDuaR52aKOJ1NsQJRWlYPzuaRnKGGl44NZIaaADAVyyWaXF5863
qXrAWooZLMk4QI0gRhtHMII+bnMpqSlOuMfbTc/gDSj3vTTb9byN01jL44OmXQ9I
Y81YMyP3Hon7fWfINTvdAPMiKM6NXzbXEr2WktJpE/nxEPR7lHcLszzBDCrqS5PT
KN4SSgvOOhGxGuL9YyR4a9avH3qQ1/mM5iQNjqAWmVNSWLEsH2Wm9xbFyR57kmSw
jVwIPIGcyi61RkcKAGPN7Y08FPrDcGyGeONY6f7RzCwlH5UpAhwGI2XZeUzRk6TD
s4G8dGOmji5tu6MlxPCwA41SXah451odvlTZZW9msHw5wrqGwk9I40xj4E9Se38T
ec5CRSGznrMkJ1YHGkXen0iJtvFTW/P8/dS5GcfbP6uJGxP2Ys64d4gxGXcuNGqk
6Eoa76yE4utz40c8NL5Y5MVBnmCSEc6OxcqKjGzIsa40XikL7cTWkKj2bD3HEy3P
z2gW+qubT1/mdr8ldymhPKY35bgdtXiABHhKcfwH5GsDkyOBGKTP3U+ifvHfUnka
hz/UMPyQpPrjRtzeBQm695scNMMzAzMaD2hBLTZBGfVrRoHZ1z9Al7d+xWB27ChS
HjIoawAX2imBlmM6Upk8C6D9vPje7qSJzYPPyprfzNwigKHW/9hVEC0q9UmKoygP
rC7dUJZpojyAMul+ZcS1IjhfojIj70WQ8KR3wXkyLWMqMHFnG8HWrH9wiIdintbI
YIx+hZ3clWuq+zYMDj8SU2A+mU+i2QAKfm04CSVA2ous3SvhbeZHwmn02+cxKLZL
tMPvNWBoDYO64ILE26toODZvXy0HtcX5tvdODVxr0X3YAm2h71ephf88+fEYmNDu
WG4raCJt00wW3Gg15sSic/UDhJps+J19OEZTb99CFqlipv2KJ/DXevaf9R/4RXMl
ymF23BDL6E/EQs1kKIayL96bEMh7VMOv74A3vD7rm0TVt88ih5kb+biH5qihjTUA
scHIdOtP8WsyPUc1OYJE1orWFbuIu/fGXaVWWaRnvmLQL/HM8WkUDHy2s95iJvkS
De6kf1SDo//D8SQ/kbz3kD01LFWp/fCfFZFbU1lnjEvdNSl+999PKBrkT6Lv86Yv
Bq92DU1wYIFiRoYBNArjbOzm/GMBpTSvtyQluPqJw5uqtbJI9hnQBTzYNzh35op7
glSBSBDgIY1WgWZ7AkqhNxA25dyq4UxvgHpyQcHMefkx6AoANNMc98B264QrwGcg
4VQmIxJKXTyCiDgkQndvjKaLuoWdn+6WLzhuG5mhZZYOSbMm9vuECNxepDX1GFo1
j+mTFG8gZW65PfrbiBGr9Why8i4tXUawpTbG6j7BYHQ0v6o84Rp9xEOZSdS5MfCQ
ToKTRPs0C1Ys2zEJHoVKVGDlgXQTVg5oK46gedDqMLAzkpuRlSPZq7ZodhJLdddq
czM6kkfC53ZCUSu0G9Z6WifAXPeB0YVFMLmkmg1UaVX7VsZ2xxfRerpgV72ZguEz
k7xkga5e9vJxQ4dNY3Lov5BC+VLUlSWnA41OKeV9vRWLxXmqtEURTYwDizWsPlHa
FPAvTBKF/U1qR5EWXkkqqQpllBFO3COQDDqG3oafK4A8X5FFw4g+Nlj5mWxu9UBd
NKYye8wFFK9VuKsMJ88zsHbe3plc9iCqzNwXcIxpQjXdMPxzzctiSxUDzX750Scg
EmJDIl6SzhvlKiYJqVPWb9Kc01LbhHiQWjQZUXIRV2HjVu8KifKhnwCHxW335gnJ
CjrVCPEv7gtiBHZ3RbUyK2oMH8Ye0urIQDNXcqljYprDbp/xXw59QA4jWoSfA5WX
1TyaZvLoyjP6taKUp9t6rXSUWDYmYsuEB7hv6fPULEGuC+9uFvzWRM2Cq47/xweR
y/lOrPH1H+7yPsRMsvFYfHZ5NatuTry5gLmQPlcZxOdMfD+vR08nH2qu7b/iJ1xO
07f5HL/H0plhJETalpAuC5qzWZOCvp1T0ve5CWOPmJRnLet8YXcRBcVFEO0ILj3d
qfxAUUqG6eyqXuopTXfXZS+pLo+NEKuTbsHyKMhoRF5MjjA5Qeq2kAXvOT2qXNef
QuTNddolO299MMPtRm3dOg334DOjZfo+5m/bXUQA01qkJLIpXicbLdwUbgNQM9Et
H2b/KGGrJbaEzc63M55AEBgVvwuZx0oVS+P6aU0K+AKVdELobAMcma7VChxCKtnJ
rif0gepO1JVQ5iQP2AXLCETfkECpr71NoDP6h65T1XJd436G2fF2YTor7smfq5II
sdAV2YPNxXkh3fw6Nk6Kv47V1iUg0dE+Pwq2N153Pt/gnFmQjrjv63GvMlJ48iB4
PMUTTOUIREKef6xqMlRz6506Ztl+FAGKyRaL30mBpzj85wkpBoFKo99IbwEz5OAi
iCJTpdnfCDsX+sXYPbZcCMuZYavWaVvwycPZEyIx7hepwBgrONSexHUJG2kPaI6e
YQV3BGFlP5GlZrXJhG/s4f1Ah5eyZzeu0Il5a2zTlpUMWW/nrnU1TEWhtu0CWt8S
zZBjHz7XvKDaDb/Pp9dONKvCN3C3M1WWUbp0+Ki03PG2uyUJ7T5oeZKnjj1YwTEj
Mc6p5m78oe9EVccBNLp+ZsQxsMUT43NkP6hGb2yZiBKNyhsTaaHg6Rv4nCzLJKuw
LzFA1dCPyQGyNxdJ3tFtZA99jaYfL89xmzxAHGiJEyV7+UNJ51j+wg1O1eVhEkOd
RyFZUvtU5v3r2+WMPtueX/YcCDCKE4sO7+D3/u99lXjTa2NuJRwEXrkfaO1kXbkQ
xwN6d29+Ek03Iw8jRjMtExoaUlaR/wVNxNp9lc6g7epAOwVAUqSAy2B4JImy7YFv
rauMnXhEC2LMkkt8sPpoXnVWvc55VfgP17V0qey//renQ21oVmU2b2/TFJxcu0Me
7ULoeFPMvX8IdE64sxRVAiX3BKESQEzHusgmiIX+8TsSOrcS22PYl3iLRhd91Rrt
3ozmrVgHjKro2tULDvJnCNPxR+v4Y2bIKaStxTaAe9X5hL3x9zdBPQjs7IrXSYoY
bJbFe9vK16J1Va4qzXS3NZ7MKluw5yjLPIBac58c/8Lj2ACk/87choJZQ0upYEoe
37EkVa74gKFmQRxlCsD8OoexOwQfkzgyJuQiTBVZmrYKuTZLkEMq1Kt4HOkMFyoB
8O+0SYcxN6YgGe+HtvtMOqrKaWYv6sTePNueQdxz/HSWz4dTGm93YGWWYbzmOyd2
nVzZ4fpsfFxhI+JheIXWx69oPrauFs98Bl0u1OL52fZ4zc/phYLFTb7nwfmjIpom
PprfZhlp3Czr4qCDEJZ+WV7xMd9PIsVcJYHPa+RTbk9y9ZeUuesbIjI2YJmgChrc
YEbau4U9mDKeu09GdlYP/8mRnmKgKIkydCizvrGBG7+OsLWj+jMzrZlq5nFhyk82
A/2SOGXcj55NDwZH4OvcyW2XYRmRJUcw4cbkL+Vwmc1eskJvLz8vHxy4QFHrIxFH
9akeb/HDr4b8VTVSW0KpJZ5gAO03efukt2NlbnJXC9k1mA4sZxg+3lVQULjTJExO
p2dl549juuL6nLFiO57c+siVQ6zMR28W32xghI9Psw992+I2T7wN+kxGePdA8dIA
Z9dueP8PoYFLY7J9ySp81aHsxEdCsOBfYCy7JH2WUmvDBkeWDYQShRqS22pq7Nli
BWllkW6EdX3dZUbhM/W5p38rqGO1bW14Nq3+osPQHbb/HWY3SaZttLDNem96Veg4
66ifzff1Xh/jR1/lq9YusJfOTOaYUxlXJk9z5VNAigRWYWjNWm3rarkAnA3N+kse
r66jMvDtUT67wx1eYrolgfja2aAACNjpVA87v0pS97qLpPKkTbgP/b2CuXjIKQxa
+AkUQs7L+T9HktYQydyQrOLjhtuGmOC6wj7yn3+O9RgBZIFCkY5yYwqHi9dmw2DX
BabfHR+FhhJxn1yrJN5ksG5ym2Gy+9TKZoihAGx3kDiFEFGiWch25q2Rf4poZLut
BOXvvF86NPYykI5tecfztXwI9UQ8QVClKXYqyegGoaOidigmT0zpDysmFHP0c1RF
Zcuxyt+2AGFE6c7XM1S7LafZm0LD3GoaJunB6nVprkpbukOog3najVYY8ttmJTGT
XCdnpTOtgVHWR5oWLfWR2zBxwgT41XQT5OhtX06i1yPKYNY8+mRdEziERYsqX7V5
AK0WoUE0XfX290qng6pWkNi1a31pIPmeIvyvsEzRu1YVoiGrMmG1ssnicM3aSzM0
Cdh33hWNq4wKmAo7z/pd6VG98y7HlQuuIH4AHwuyu+FKuvjylMbWRyxsiiLh2kyo
ehu3fK3wHTJ6wAs5OwWS6WlBJn7vxXDI0exuDIVfS7FpQTePT+2j+BAmUKrqrcE5
GOfA4sb86rLmMt3zhzLd18paNvv/Uihsx83XI3xGW9u5SP76owogHESN+V9d3kVy
xwjqp38VTZ7+QPOO81p4h4RldlEz2s5N39Sc7UYnuIRyM3Oe7xgAwp4SSb+hM5Dk
ChSP9JvUlqC4GLkx7ZTk6hsJoyW/bI7I3If86N+QbKP+kz7hS1SZPtC3V8yP+EWK
dGICuRxXY8wESX6wkXvhnpVlo77hRLQ8twwIXlYnK6d+mfvb28wqcozvWdyRvjPK
RiPZcdi/3KSFPLPM0uMDehGrIoZ4xZ+41KVWMV0lTklpaRMTEhhdLryGmqIinbzK
zmDMHAGR2ALQjBp7D9PX/jSgcWXrQdYPUuC6v382cMCVkjxJnHbIH0vMOyY+Ykx8
mOOBd4eq3VXlKlEHIyEbSKK+7+vd32HA0+fqfe4BjmxWZi0woxfRob0Ly8v9LjXr
qCyrg2F8HR6CtZ2yxaL8G5MCAbVo5sWSb4Q8yoKRrLpcIGMCWOgb7Vks5+VFIpAW
sx7oCRAWFPcEWTjuWfP5jw8yEHGyhDalfVV2gONhH5XGGjqNRnMs8qWNaz0I1jlQ
SDrVMN/MGtaJuv9VAB/X0bIkNySampi6A5nJL6S6NLzGaglu1W4VPVFC2Ogob1rY
Yv9l8preHQ0wrCbiNgs4w9Jn2CCDEdGerm7crzwwkEC8DdZHLZWPGokScoXbrbOj
mbhECHeOKAkj/zUAGR4nb83A2L4qenvxpNv+vJK6iILP3jCu3UeWxpR+ZrqoVkGs
nMW5KDyCKmajZRKWXW8EVBconyyxT7+wk+x5IFe08gk8LnijTt+5je8n1GEm2m4q
TOxDehG+uB9125MBhUWBmzxS3xaHzA9CAykLJHfDD9D6wcypQVvBx7bAZ8x1tgIf
IwHcP5q6UOFrG/CXKEFVJYAC9mUvJD2vPVEye5Rs7TMMhUpbZo4ChToDWkyeBvN2
1wYtjWVi3Umtya1rwpIArn9HPeqCU5dO4Jh9pDx5RoqlYn0foVTCex7dvjoQ3f58
6GxCcO6om4qwfofxeWORv42cahnOs7ZbKbAS5qKwncsy4w81zUJJWMTwr5BXp+TM
9ywbunYauY/g1MdyDtIQN2+QFfNCHl35tdBjUHLnQU+7wvWqdS0aG1FIHYkfQokM
L+n4YVbyY/X0cwchtFB62M4jPlfQC5NvVmfgxEMA0O54AdJ1Bqf9xlCsiev3F0H/
kQt2LKBJu0elCPnmrSHqbiajDFz/zc0HL3/J99YJCrCPHdnwp46V0v7K7EC2lvDc
d62XtH+rOc2+6HfmNC++OXDJjduJp4KA76nn7oZARq8KK4CBVlaEQSbT/p2UqoqS
+h59ZtFi+gCsncZGD6qk7SJOWO7azRfM/jdma5o1t/1WY0ecdF2EItliXq9TJZoV
aB8+a41BIlxY4S65Lnuj3Yn3PLK09LHHPVzzntvwths+/klNMnRf3gRxh/s++zBZ
MsclYP7ygg/9qM6QpwlVGzi2jQmFsti3U6h12+/FxeWRMVMzNTP3sV7hqkl3QIG/
n7FXIpaCvG4Bp5XCJbXv1WJd3WFAIxKfIzkCHmIh0a0s5Eb0qJ9GWwPbOCjTgB2J
H31qQmFby9B6DurJsa9+hix5bPWi0fphNpPjHgjQmBwekRP22geg3kJDr8Egji36
gsSxy2r95Fz5OLPvz1aT5G3U7egEYJgwZjFZ6TV4dd4OaqXpjHpXG/L0EbxmwagN
hG60EbrQBZqr7Tyafq8aCWghd6UcQrTRN48UDGK5rX0jKVIDfk6i/1dMwYeHDlqA
6Mmn0DxEaRDbH2i/4GqFVMIIzeP5mkYwvh+5LF5YbNAMfUQnFhDplxO12Amm5YPK
WaMnFxdrZKWJKyCcHpUgp/CD3zSczX37hgynKdbIGVE+DbOVd/fTl/NN7wp3Mzkl
KwyfRQf6qJ/HEH12dH11/bJK6ANN2jY6przupRCGcf/E65RFWS3gW4epy6MTaUI3
v7zTI8wh1i8Br+DuGK4Ok0L5+w42FFH4Ix2gfYJCUoNb+TKVZU7jAfepvPro8RyS
RGUCinazzGxEazYJZFhvpXnKepC6EMQy7Ay/1thOx8zuRdP9Az2fRDkgPzgLiHgQ
DAeZjse7YRx8bs+fSYp9nlasbmcIzIeF/f7+XDJGL1rbQRoMJIN82lgK+i8RueN2
EsLISdddl/NnKd3n2BdHaiG3Qz4eOLGpKa7AuIozzct0akuM9BWmDEO8gRBlP+sx
ac1d3gMHwc8i1ctiP+0QyJRVBthHTp8kzfCu3wzt0HwHLBHItrc8NTY2mdTu69gk
H5u6Xp8hoyVcPaVvKrN+0r2eDW97mEp0UIaFcGbk8M0AHEg4uV/8YIsfsiEISg50
Y0+3qKmXmvg30uDC0XYfDtIydEHa3oHY4eNtzv0YdE6D6H3fwFKbBm9HrbsGlOye
K2Nav33L89x7Mf5yu8BNHGMR4bjcN4RatiuTr+Vt0J+7Gjrt7RlPfpJx/BM0L741
4+/yV4TI1sqkSb1rtcu23/SWV+J5i7ABIi2Modvlc6elQgZ+9hM5Di7eGc/djqAB
XZFJ9w1Es1oKYOLN3UJfbQXgjZSfYK/+WHjqGXCwU6gXa/Zo7LlP2zm+qkWMXUkd
r34J+cst91+ABRdcw8eoRTp6M7ywEJ82D2HBEIW6MK6zD6oMwkUdEg2yLUFTsZU1
tL5J4CCU0MIIWJO8M+NMKdJ4P+wtQ+WAddUMTiFK6NEmB/Xu5VNXfutgLWS6O5xO
Gd7eESqIIpoHrnYN+nE26OjHODdkL7KHlo5NJPvbMc0IdcaymA0vpX1ExZvPu/EE
tYlT9Lj9k1E4RtAUvuAO5Qa/4NjLeKQ1RKT3fZ/2f2bfElfBt1mtAzY9MiV4BF8j
6Fww9jtOhYGGubrk0HohHvplgzZQGfVleaKvIsmQOtsB2x492xWCANFrLJ1Co8WJ
t8oSY5RtcYx21jOL8QeC+30c1JHOHwePCwNVpuZA2y7gnvsOPcJN2/aL3qPkziOL
6I7cXrIkkLHRMLAxsQFUvzTxvCi5ltTJpplZ4xM3ECe0p2z3eL56k2p5sZ9SE4Jl
HMGdYxHcFvgDp/xjgV7OTAtOu+iHuVpHga/j7JKFuL3aPt87Byr6E6bTS5Hzak99
aly07Zxe3MZdu3qrXD0Xwd8i0hQAwSIZFaFpRhwJ2Obhtg1rE7XK0MD24JaY6Az6
KkBqg2DvxMyj7OwljNDF8tFb0DudLkTleggHKGEuzby/MGeRec+W3GSPLFoFmiUA
FXP+/Zmr0aXrdVcjCNyV8hv3y7eyLnyk6zEIVJu0W3fWM8STDpsHo7F8h9467Zvf
ipbn95vysNJ9QRqsUVo/1GA1MCjMkX0XhU4KLgNze8kHSOJgtOyFGfV324PCCcft
7HVJH4ZbQFgGAG7bqeNNP881+KQGYOrwAnIV9k0LvM3+GVtf4t7lLUogYMHTrCbZ
6dvMIzyUN83VrbKKfqmrkxAp6JtduuLu874HboEgcv5I88OwF+CxV/0lgr8/j8Q1
3yaiVGzM86f3b/mbxWCfK8nOfvLO9M/XLoExgduUH7zIyqTx+t4coqXNuUX6hIqq
DbXHJ6+VCXtvN1rhNJH6Prlslwuof7pm0Y3V/n6m9o/nZyhCmmKJr+Yeg2pCabzC
+NNrHnkeiGISuYWuUSw6G9Q9EsGygViV/wwcCQljVKvK4dXPfavzJ5rRksFkxjmR
Wu4CDnapr7WNPTbaBy4tE5NarOhkFVgn+rcFM/dFKbK7GsMQBsb94b9MxiVi/JJu
+nFV09TBVzmRdbRqFDnU5Z2DX8G8kQ7jN8bSV1pyc5M8jMQwMDltHcKC+4AQEdb0
XEo///6k7J8LMNjEj+AAhNrXvyZ/RBCuhxDnq9fA2ZVSOU2oj/RytL5wVe9e8f3I
awku/sb+PB7tsZD0NSDuovgTSoARivroqFMmDPDC1KMPxx+GbT8ZJTXrGJ/hgz6Y
80TBzGIALYWjdJFpgWPxgVq52IBgYEKNv5gFjB6r5UJ1wxHNff3CCFHMFgo+bt3w
AcxIYAY8dfdO3qdbe7dMCYPFAFpU8l6xpbiSdePG2KKrNUZpNEirZB+k0dyerXq+
BfBLxs9639/vD6q9+JRj7AAbD6iHqgwhRXG7qk++dmtfSXujqmLot2gEZAWzujSA
j3JKahE/gANSSpnoLe5OzPNE6R+NY75jm9EYMFGcNfmHTWxXAd1UKRi/NxAJchRW
46KAgIMdyq0zDN1JBTBUWFfxZvd1OCG9yE/BYeMX2lrrIvjI9k+QVSATgpn5xhhE
xbvnonZgvB3pylmNQYAOe1JmauYxcL5Gb5RPrmUmWdAuSCgm1EYozHk5u/NfB+l3
vlCdI4uxFjE9/SnYmeHITfAuWbTsyOWiyupA9UBv+selMvEh+r8ExlmAN2xaBD/7
lgiYgyCdvRD0s7V40HyuOH8r83i+n35C4FvR6+yqGAB/abGEUsNxQ/D7W7pF9gcO
hpXHPmA1GxlYFKWYLM68hFxT39yLw4E/3IA+ucwwXZgGwouq3YQjLNGRHUm9/xAE
or7j9hM7vdXu45PQoUJw+ko6fPWIKUsuPKBMO3EJwjX5jHAxYzV5ftbi70Ts6vNA
txoLoxuCpS6OhiZmO07BYcNdFEDuDnzfeAPL9sJfKhvyySgenMyKKAIkwjEQW5Qd
dDuqWLoHWUNfLGb1Gxmvh5fB/qACySuWeKLq905VbwdMS/qfYqHRPwO1x1q3drqC
wZWQSEqQoHiAsdwCurYDEAW7Smg4jjh38qKBmhypQesT2HNf3qTC5EIxI3gj9q0/
F+TTqfwdcR3Npl6abjdQO1a60SFvq3r9Kvw14ZHmRuEx0hsYYtwfA4yeakNj5I8Q
ICQMfTRoG9hzw7Rw6rTD7d2OwSLLjOG4AWsCLMSoY1A2gasATWFnfC3AEVvsED0E
VRYXJOYTE+voo7RNdoZvpqgu8sv045v0uYr53k8NWIYj1ju+p/i9Ue8xtJUN4UE/
Xc08nsbIF79PPYFWtNgNwJHS9VkS1r5QV/FTTJmSeGjIPdaiptVRyt4AYJ77+QKH
dZU/SQT9lKkWnfB86iy1bVyl6fofQOcDRL6Pqir0kzBzmZX1x1AijUKcmPJLZris
gd4L4/wDWx9oD/MfFq3yPpmYju1QdbvViJaVYygef7gLj6yt29ZnqIUTgsC0og9K
uBc/forLHc/brzLaTNfZbG/FNftLgAe01795jfR0RvHHSWM+TFzm7ANc0QAYdu0Z
lHK5UvDC4pQKTpcA1rrppTQifNVjqNbPnHFf/CaZSZW9ozP+fB5GwcfhvHjNS1Vz
WEjHGqb8F0o/LW9+0IJQeNNJ1aedYYjIzPdQYDJFkBgY936LFMluJqS/LmhPtMor
zwpYVNzBA4Nkbr3PwNbcXZlBTRnPzxcY/sUF6WKWiSUzdbL2j1OH8dGFn0UREIe6
BvZMvA/IjVqyUymvhMWu/cCggUdogsBjB4hzQNCAIURmnICA8M4GIhkQc4INE12A
JydUoNvvzduXx5vkEtDoJ0+aPxo8KDfHxat9jIlFC1wlJ1SY/jIt542a0I62FTZH
hNIHfRby744wm6bU7a9v1pEk98ia9LLTnZZeuAqw/XVpHBo3zBfQwK2JsK0OnMrk
Ypnr/pqxyjBBzJe9HLPhr0sSgg1cJj9z1zlFfDXOs6GkMKT3+y5TLGi4lYFdQo2z
xMVJ+2GNCffFdut03koYQBYPwLBsMfv8CuGce6Cq/7df28fnVPaxNDx/EfH7ISoi
KNuMJWaCGGVoIPiNW4S9ZlNsdUlfWKv6F7IeGCytjNal1GBzceWNUprpjh1iKBVb
epwZBDNuFpkTYDE2MPTrCBlEkHiywgcfdkseVFu3o+ineaxFR7Pa8Y2Yl+Q1SBvi
kOazBOGK8i84LZiXU17Erfq2PJfSA2yfKwdWMGQO1BawfC4t1SPZxI6uvaoHVcd5
iGN4Id9GDn8HnxJELojHqYM64pbr2VXrSSq/jLz+X8E/fENkIUUiIWakV2krf85N
pze+UNoenJVR3zhei9LKhANoI+de4jIOWB4qKl9DQ+CPBXG3fKu2lWBq+c4cjsC/
yyq6HpE8+D+rN9RCTfPV6SIssVW01t0QFjCAlZzJoARSBjFBvSwPIfS3vVK1bdw4
1+ZJV5UNko8eIIf/Z5VJgXmMqruj9cD2nc2YbHYFNBzJqWhWW0RDYnnntFMbRlvo
65vjK90sML45lL8AeNsKGFrFFPwwb9vqomwceK0+XVCHIYSz+dOy/hZkr8THHvEH
pe6g/Vb8RbL9u9HBRtIdUJqIDAJkSc/vV1fFjKWzKU93n0UlBhaVjXAsZNO/o7eY
mNOUSb/+RTHxJrRACVvibG2NQABPtyW/21Mhxo1IL0dGp5f2Ay7m9YlrJysYCTP/
aOWPiNZv73Vg8FcwL1738bU/I2b52XEq4wD8PNC5ROldanpJcmT7z6lVNzn7BKCY
B12hfR2AkvMvFygXWWCBBckG66fFvhN44Pph0ICYXB7ohAWRn2mxTVyiFVY/6uDr
BoqFFdrGm2iGXByAWl4MrSx3w3q8i0rmfg7wegPn0g3wSFGy6saBsTOyEL6XkJoK
oAlOtYp5kC5orN+Bg7zUT3KfyiesS4aPJJcQYSArrqpEQOgIaxUFkaAneODfD3h7
K+z/PU1Fpv6yHaAJ9V7ha5kUzzkCxanqiL0jEzw/0oUVhh+3yFDiVHaMKnGqfaI+
OkroGgLNaxqr6cvVgAuIGCfCYhofBH6GO2GkQ6/0hU3EhzVznzPKxSCLPI/bwKim
QUmokerg2IzqeyaKHhgFjR3+QFhaSZjeYtgJTQkrvJB1JaOZvsfsV4cYW84cvb/J
qezxQxE5ijkpP4+I7ecihCKmrSN7H8VjDnwo+W53HBYOZgLmu96Zq4lBE425Ft5q
LOtm0yqhIqpFBsrxwO431xtyffwvRRYmwV0mXDhjIvrSkeRcu6iYoai7d0uC5oHm
Nd3ciFCaNhuY8FSVmUnHXl5hKETQ4AJtGhcwGracEvDOfUDc/Zvjj/nahyB/ZP9Q
TTqW2a9bLFZ7MBT1wX0CjVTc6bYCBswP9WSBKvtDZMu2GqJjtUDb4PfwzNpKTzCi
2qfY54pRj4AtKnlQpysB/6/ZzXvNJtUATkr+BUqZ2GYRG2PsIbcUgQp2DiiJWiF2
CTU7bHc7+V+6QzXVjAvIHiVFMo18nt5aES0QnJuneFyqZGjpBy0/Y2IT3OuHfy+H
ZFBWj0duELuND4OsudJoQNny9BNK4AWmTMY5q32mMwj12FUjSprQZE3IceeizNqC
mvszj2GYPqqNebW5F9OHtczCGmYOQggwDE91XuD/knSuOjrbtbXeS2/6ns2CWg6G
ZAYTgLRJC6U5nMEFm4RwjOZy5aMuv8Lbf5QyDAH3yAzER0kTJdhpykqX1xTNz3lt
b7sMMHbppcN2vskzYtI7IaQI9Y+CaL2ZbyCXfCcySgyXInz9K9LRtIGr1H0bq5yV
saGVab4LdB2sTPGk8dCTI2x5yzqosTjF52RAq7ontFkhUJOF8Bt0VCgbT/3Y1Thu
BEguXaACT4Ly2GoWo4EUeilNan60VDm5Q7hs209COMu7C8eCBWkP6CcVTV1ylCr7
qUlBi7P440J6gjjtpXBti+XRgvyClNfz4e7wwAsGYCNH0IsZOS1tqomU4ew9WC6h
WfkJJ7EgjrmrjFhqXYE8QJ6wZsVi25Ay7v6FQ4+G+iPLYz1y6txZjMRGfk+PA2Jj
1C02GoHaUleuMa4UuJNO+N11gLvKPc5snockUG+kqYICLpTdgqtQtYt69XRWnqAj
x655SzZLWR2mXcvkKn3Gg5B3mETZAmdohnv5O43w9GWgTRmi29YVpbR9lI8KQblf
Az1v0WEnDXGQeL7CtlRn3Vf2fMT2w4dtm6FxIz/bnUgkYwcah/haCjfDXqQnBjkd
TZdVXSEOB37N0B5a9As8pLTXF8T9SpyiSNMdcx6uiUe+7idFhu65O25oNczRZuTB
oWTV294obSgfxcZdJ9Lqx7a2ZmjUY3tIqYte32LRrwwh2ySvarfhjoUb7r85LlSI
gIhBfQE/IrduGGERPwycyzYHtX0fJUNMAbVBs0so6LTm/VsMVziC2q3Kx+I6XgCT
ThR71BNOiWiwttKQy6iL9SE9q4xDmtUujLxRMpNLFbwGjOauvBEyC0qEaSu93GXc
bRNb5wnR9Y6sWhM2nCLwJFOGL2AXkZH144g5iCYvvDmO9HsTQU9jrxadwFZj5jik
OVtqfj7/X0WVssSl8nB65OrreNdCN+h2+tTX42UkRJ1DwdDS1LR91HiQYIARL9ZX
5ad/t/9Lu9tmr6Nnjs3fLqH6TaqfPzBl3ZJ9C4LFrHoRPOgHgteUPyLxbDbDkJsH
z9zP98B/PI9GLFktrRL43icBEG0mYH9Pl/Jg2bqn6SookWAYINHHYZ0K6KnWstZc
dvYWCxBAv6J/7H8IfE8KMubvHz/aj5lwGhZ9BNkfedYbs6VDqjcAHT+dQc3V3eSy
Z/bMl2oHpoTbqyS7fdfUhazHa1fmHRNU/NkKjgvSi9ghW/lKz7DyWoCKQumhjP0f
NSn8hc9yJdXuw2NYah0opAId8/5xy47Yaq7b8EU7Zz0NQsJncUSvaLcUoWEiIGn7
6k6j3wzNC+dy0XiVL8EiEqbjgwCgxdd2cVgoGchYuDFVlGXdONusQN3G5BEvd5kG
F7Cz+ljy6qCi9uzc8tLSlnb7zYDhPaRIHKP/VdALr0T/mEF3xjfzaAbkuPDsufFb
PJYwIQ1L3VaXyb0wmClaQE+bvNWO2GZ53h/38t30OtN7NBnlBAvMESqyU9b0Cmx2
kQwhmUV1EzZvw7jh4x8v6yAJssI+ZDlnsW/7gp8efCV9VU3hV3+fG6ol37ZGI+0A
UFqIdAvbX+a9X+S3NZrYiFItl07+zX1M2u66fLxKpPtU2T1X6fDEbEXtJJDRxgMd
opp+vwkkUt0Ju/Cz95d+MrANvv7Z5ocMAp3BPS/0RECUeJ2+iuXqdgxvgxv2BivH
CDsBzJvfUiT5iBx1IDll4WPMEBbjXGy9GC8b8gL5TmTHkgIZSDSPHb32urXwqouV
FC6dU+1M8IIIi0my5wnjBQNI4fZg8bpbjL9tXj+EUFPs9L0/ycKF4/TY13LsPIK2
U16Ta7BMS+jAY6k3OpHxaw4V/opg5WP0SFrfxRK6zk7HS4bJaDtAL02ZN7O802+D
Rb/1AY6Rqow8MilQtFV170XSrv1C7N0LGfVepVk31DLR4RUbrPy0fjuKxRIBhWZ1
G42UxUzqdtcutvnr8QHPsVdUonvGgTfKC6xQLmbeO48xXqY1TBvtawA4QerHkXCX
JYRnFbSpFbrR4+yPM8KbqoGjWclaRewVuZlG/TW/VWtvUzs5RM4ngQRgDDQPGEsO
TlPkiD788Ji+kF1D8NDwOXaj/JMPcs2do+dbFPbAw3mBu6TuoofVNs/HEaliv6TL
83QFFrsmQV/rqRiD4ivWug7wuxvDhv4XhpOqiTeI855OVsLLK82nA5H/sdPqRUX0
bljmATW9a8mL4o0MdfYP7JIGEjgH1iax+Cf/Dw0LPDYMGlIBRJg0JsmvKNICy7R6
549V+JdqwQhrLxowAfYGL6iku1+fvkMTEsQkEW2TMai9EvSNynlgLl+Cb6WhV54s
doipp4hs17zbUXLweDBt27DAQ9t0FRDo7JEuDL1NhvkAv+TKgjrAIit/X3l8Mx5H
6XJjhw3zn2oJevUUHlNikEc4mM3HZa3GgxNvb1GDXWQdQc0Re49LqXmz/nslBE+i
dUzg2K+WZPXIvqpHR978wHGbYc706tJmEJ77n1ggvqgMEw7pcf4zRWC2vDeYu48S
0IM1gr5YBgOAOtcczc8zP65NROuZWjGHT8y0Uy4M658+avVOZpkWC1CMjkuhMdHa
MYvVfZurSWjToGiZuw+mKjDxIgys6NRnWRIkZ9Es7W71NWrWB+AFFROz7lywuzoC
2SX1qBSu6Fs0zZUr5Yur7jOBl+GojjMExV5umulYwgmGWHm+npsxiJMytohBgj/5
ihxSFgWR1BfvkmRLYfHn3H5u3WhVioCFRN5fJh+c03VguSwPdU+T2YAyFd1LaLQP
HmzMnn8Y32bwsz5R+Jh1z2OF4WhZJes7bYM+6MPr03Kogp6wUOsXg+j1FuLF8V5e
Y43gG6QfJZQwzvD3W0EPNbsmLTqmbHT/jqTS6W0xhZ7ZOt/6XRGSiU4f22w7BpTH
RmA2ckiTENnCxTHmUxEok5R1t236V3bRDGi7BsYAhCAXFgv63PhA/3XR2KLc66Tj
LTP408SLZZ31bYDo1+tzGNjgcPRgjXXSlBPbbfpD7c6grt5VZoGC9D/wcikE75RQ
O9mNjYNGlV9R58LR9fa1hkQorKxuQoQJmK+wKDBFPxQYVT5EVn6EK5sxMZdrbFgr
+CnvTDUT8JiaAG4aLVL3X8DOnljTsLgL2Bjn5E3mNVgQYZ6M6WUo6LfUeLTgZy68
Tgrah/sprKh8z5HqmBDUJq1YPaDLMRB66bZLqLYT3MNAXMCH9NBhB8Ltm3ZqDnCi
z7o2BqrXlVmaP3fbMbPz94R1aWsFp4VuoneaLomHyAh624fTqWWRqWdKEBsqbIzz
0eCzWECx3uGn4zaaB3ELnL7wDa/7C2djxdOj46/ndWb/SyDaANmODq+wEWhBJr9j
W/iqsST1X2H25YV3/439UQOraSRSV2CMtF0CWt0YOX2kZNqPVs1ZnE642IAaBUJ0
SLfsrJlbmaXIY4ePq3rRYx2mTuEE4TszlEmRzDvlsVnQpvLWmrUurjN21jQy3s37
n+APKwcZnyyYASQCbD4Nlh8Fg8z+K2JZuuWZbykLIcfXvX+bXYRDrHNrVhdkTfpg
m3FfPfi9Dux6PRosX7gorhp2kVOdhpeM9PzptsWIPoshMZRxYGeJkOKSzlRtYG1h
AGQj3iek8Hk+yUiWrIfqTD4C9rSuxuKPWc+LCSVJSojtbvMWS2LkXdsMlCBbi10K
94B5jm3jbBTzoHAuhbq2p4UiCr2Ksg6aPgCuFJgWypySaNtwtP1iJRl6faudVHlh
Dk7Usi21h6VT3Mv+wto8x/NQeFQqdPVTQK9eCxIAHpASjHGqBsSeHB0RWEj4yCrG
+ifN3jnkT4Spzh9B1YP12Vx6vpoS5hXw5rA8g0sdZutNtrCIrhvJJVR9IUpjltce
O27d+vUUmJm2bLY0GgDJWWAzXMhbdGFRqMXcHbjCWvDkWogyLcH9Ut/6FXPJBpCr
xJbDeHziUqMcdYH9LgEijwMKok5jpXxtNEuCz5PHVbZ77E3P10d9y4lEnsTvBOeR
aYlm65yMBAhKjHjn7/Ilhe8izUqhPC04LtDX9tjRFmuaUX3QmKbsk++nRQTxT7q5
61osWyXRKLmmRKwovrCKdq34+MoHrf0XRgvVbav6XOB/2g8aJI/5D1cHTfy2Ujzg
cRcTXY+umClrdmJ9MiPsNfmDTPachhgbnEezsert5l7Z88gY9m3p3PZuSxwNLOdL
3hYklRcrdJH3LbNXEtGYihP191wo/ZQjkTBBTJwmrc/bty4zUoVU+eY+cvDu3BCG
oZf6mBn5ATTGo61gjRspB8OQbRLPj0UqebC3ZfA+4BP0WBKObgmpmd2HCyQxK3PM
qFw/0gMlzvZTs+ootXPvuRRbPX8puty4JvpiqsAGQsz68QcxaiUii+283CIdCNCw
LQ6Ka4lh/i08bYaEFQ0cbLYeAcb72EFNG0QpL2PTIzVBie58/yOkeJvkbx3qBAgr
aIkFyvatiFwWOXN8GPjA7HIsuR4SudjuUQB4jJSq9jIPSDNZtMAKVVsLANk6Bo64
bjiT8y7pECLFyU0b+CYnjQziF2TS3VePit5An0bInjFSwjZiDHCCdhW79n+CjVsr
XQE0Drj8s+ma6NVkIyEFuYK8ox6z4cF7XF/3WWmr6jtG6E1QVQ3vl4KIhstHGEc8
SCuwjZH7qmXfFAzG4Ygug9dBUE7H1Xz2gtPk2FagLTC2tkTBUH5y7FRHjpHllN4X
YEXy3N+4xigV7JISEiI+Zyypub5CS+tmL9Zycz10eD6PjZ9nA4MsDnVxdRjd4bZa
bReQk2QB+99+B9vxENO++2ocPuaqWFG1q9TaslU4cz9BVfHec/GV3s0q1n7hmT7K
53o4dwuO2HVWYjBvv0HGc2O2J9Hh+ZYUhFhe3qj3GIaPKbkUo2HFWrd0e4w7TdqK
4rpkeYQ1UG0zziXJdjb4/TXNSiEFtakU0ZLHIRwRIVIF/P5MQn2mneu+YKrkQP/y
qBF4z3xfnvlgBBFx99LmZqLiDmM4t6xbJfS/Ch0ki/zi6AmvFZAglgxWp5xf9OKc
Lk7UySUVAtHo8Os7RKENdEJJktcD3oHnOGw+y13EqBaDoIPmBqhMOh/ks8t4rLAD
GrIn+Ge6+lic5lSVG/SsoWV9EehiJeyNI56J/repyO4ZUD26XQEIxOdTxyRd0Q9g
s9e4lRk9kaGxTABn0mKGjBXTOUg4mVvhZVol26s3rWfqE2fx0G3TFBHaQndi8VxU
wbJfNlYa6qZY4hXvzg7hzNCHBNnp+XNWUZ4ggUFXn2QhRs+pbmcX4wyVIE+P0RRh
b4J9CdkGnHCDwyQG83nKTo909MRXw9erpQP1UBo7GmYtru5wxH7c9sJXTC/1HOwF
awmjluFjw3lU9DMaDq29eHHnum73PNQV7MKcBQNQo4DrnI+DexpW0IlR1KvSYVew
UHfZ60wVkRciFeoe9A54z54+R7A3NiFpMDbNZXDuouVfiyB81+ZIDLlm83J7G9RJ
lMAKa13WVEKg9dgPBcoI96q9fH9kWo5jD6RYeOmY4VxGPD73g8KPUG/sCyOIyc2o
kqXYoD0xZlSkzqXfk6VfufXIvoATGjU4gXcH+l7mmdxmS99U2ndQ9ggPpFDoUO4G
sCudc22YcmGGOfI1v301odJzUqMpMVcQAgIYavezoHCWJgfC/aybTMH4EBUv7Iul
9bvICu90HGXrD6dLwmD02bU1CNlhwR9XnheHcTOzOdUuIdI2MjdxxE8DQ+9vAn/l
YIzbhU7aPu+85PYmISpso+OD+ZAFQ3D31chUnny5p74PVrVxpU+8Hi39tVIBqt8v
7nRurbCh6kvItqTBJWCTYxclaPo3C0GeLjZd9UrpIAWGEbuKpZJqVXTynsC0cIWX
9+WejWTDtoJO33O4z6tQDg1/gdFjXcXMJRysq+wFRQkeDO5jxnFdzCSrukjpJlt8
zWb6qA2GfGDjpq0mPlDwdTa3UhT79p8sWZqMcig65JGZS+0P7B1IvCRNQBpoCGlF
liYy68y+qosyHTiCKaZe2dTFjDfSOlt4qIEQVKawPUwjiRKqG5/ghSs1ltODr3Le
sxJJ8EjBdlNoLoi1spiIofU6hW1NQh/GMhjUCkWmjyj6+gNg3nd6lJZztpKzdW5n
o4nz9NG13/9ZinAosnYVZLlmR4JKbCo0q4FIqkr5PxcQ+NfajI8R9Gc9wIVpiv49
02RU8ZsRDVM71FOcr+0nDKp7kgrUtMwKRl4JUm/F56cOSRtdCyoiEqHEUMLK2spP
R/UIJQkFSEnAXpdldZ51QVfNizjuhx/fGFfE2VmlcvmOpR3iP/AfovsZUvT0baYd
a8edq1IqMImqWrJegc/7Ge+PL38MtbLjTrE94dGSiP9wgNZ4KUZDojwREm1URY1o
/ePxR6mBNNTnrmbIttPGDP96cVDXWo7noJqBOrDgklwKUpYqlM7hroFzWzjMiigy
Q7ZhKGGs+yDADnH6odEeY6yuo9yuRUhPe2jm7PQv/W4N+bgE/bNEAbqJ25+vtvIO
j+irkQMk7M586yb8wjICeJy4RG9GNP8HNpZa27mWMY1S9C2bXLfTh5NvuM+ENCCX
hBOZvDISWpwL9cvvzi9ij/TX1Vf+yHH+0eEER14Up35mHNmz6ZaARZeq4urIh3Ek
nYSJ1GJtv9AzwHXFSGDRWixzVx6jotpBoZGxFwv9/etcgiOQdls5cFB9LTPorn8l
1yAFbc25t4tiAua2/uZAcu++CKoIUIi+LCglWaGJ1fZ8Y4nvNU93rNu6tLMw4ZHy
BK5FxKIzI4FfxASMP/CPHjWWYXA0VqhRW/AnR+6HtiNor2FRXcJFxlkp2cjr297e
cyF333pDbacV1ET9zUlsv7D12rHzCQGVzVMeIbWd3hIF9M6/QuY/rJDD6Pirzrfn
3Ru36Rns5r8WtcWxmcEafyMWHsZXlfJ4WUDgeR3LQpV2mnuaZQn3YDIOlV9uuYDd
AePzh/A90MxClRoWxQ3m3LbOuDlkS/jrNHsiX3pzYm3F9UUH++Q93+n0QXBh2FyG
H+7TvA8rvRcVQPDqucSTYMePk0KsHlXcdVW+JcPVzVA5V/AFS6+x0IL89S4LE3Dm
CSuvDNKgMyfoPBSwVyU9BT08FOxhH9rMIbNlOerM55IjlE29xCEtGtcDNufhNslQ
fFiv0SwB4xWD7hu7phmIqKbuuIUMgu0swEYKcYncEmT+nqVlLrKyqUA9QeHTpF6x
GYODlL3mwiKZ1SzyyXZikmN1pdZ9Gq+48sLLBzkcvTuMgwxD/wHWNZj6OyMeYscD
rsQTzdF4hXyRsePUukdmzjkACxHixuz/s6Lz8dy7iobtP2Qc5w2yIhGlhDCGfITJ
+eIDLXMpBZnUU7IR9xAV1wP2t/5tL599/jeks8rdIDOtk9RXWo/j3zp84bUTFl/i
IaGXRWWno5xjM9jy6ueifosNXrqHpPJu/EWXheSBV+tVMFsubDLcJCv6Q6FnrZbk
WLF+8gEXKBuHrvpJQ+3M5POjqCkHatWw6Owh+vItctJDT2IaWsOOw9jO7YktL4Oy
Kbi29tnvWo0S5JbSLg7d/9O4YHuZuEQNhSbBgLYAybuxD6c/qot5MgbkiEwbybtf
hD7MSlekHR/tiwogG5C9C5dnGe0GD6STfTyV7tBFzqpSkCFt6lnOxRaaDjPtGPmG
MGNlKBMteTUyHR0OLL5SSxwGbuxH6exal+nY3HRtTDs2N4L118g5V0BT71xWDQ70
R3jEMU+iEaCLZ4OXgX77lXYl6ylOgi0cXzCAUlJcycZ+VQqR/7r2qjjC1BPUGGT4
m6aXojA2hX/rj6K7YuLu9UrWmyqy8QX+yD6PrsG+4nGemhs5GEckG2Qm2mNjZ1yk
dF/E8EjvCMLKoB56AjMsF6t0iCeGQHFlsQYr7BJuXX16jtoxm0YlC1F2gqGYuCF2
Kh/sMrMJjF2zW2csRLSRPzvFtW9EmXq6nfZvJfxw9cntUGf06p9hMBaAx3G2vMRb
5xhxqBAYqF4XxQjq1Zr9k6oZYrqDkCYKMMnXwXLXZ5I7ipfe1qStewVMJrsfSyI2
E8r1XHxXzqteEjC5HOm0zzkslx2Fe5fWU2cvaO61ggQWzu/cQLEaKO+Xouma4pgj
MaLgIL9DXkLsMLqZsAdeREWKv0rJOiAHM9JRHMt0//OKvG2oS/fYdU7MAaV1SjwZ
8yKbqfnwWWbyysXGg4DmmAKOn51DfTU19rrLksGj/nSRo+ojjGfVaFDEM+SNlzQi
3z+cEDfkgbNgiuT1kWRHtmeHKrdQxgGuJU4VyqDVwCVwSA4jxhV+rIKh20DqWa5S
YHhCKNqMjnNv+npaOaNXtSpNjF6HUbhT0USRAaktlPImF2Op+MpHojF7sOcgpx5o
k5bCLN2jZ0h0P069h1SEwG8xcCyjAqWeccaLK0z2cgDdYy2dgJ3U590ioHHiqi6i
APvTDzjIPsxd3iTq9CnHyc3Wj4b/8AbsrckpQM3YBJRCzDAjvzKdwdkf837veApj
wiaHXM6CaL3guG8JWHrd8OM3qVm/6InYKypmNBM6zEzBgRSZGJ4x7Nbr2/DSeN1j
KW5JdjycZXPdi6VyKomjh21m6TNh6sgJHvAoLqJjRHTGiLid/uuquwThZKHcKFFk
uXCbEV+lXRhajIGQ0mFyUeS3j0Xzf+HRVSbbtbgETZEZLDqwotE5XOzafWdfHtu0
PFuWo0PwORK+RCZ6w7dqW967vyMOcS3DV1ruDMlkuJzjLRvBsffCH+ZyhN8+M/dY
TXecCNtpDTeLHIwORnQlSpSZutPabBqX3CQL6kCJEltNMKuvV1VM3UYH43xXJ3Wd
du0hhzu/Ew+o14FNWrO1HPzrGkbUMiDW1xJW5b7tbyCWjgdikQzRI8pmX5UxP8Nm
bvwtcrcd9J4y7g3CyL19ovfs3Fy1gtZgUXsw6+2MMdrRtBzJcp2OpGY32V9ZHh1Z
f4c3NDNkORDKPVN0VqtyJIOALfwHm8a1IvJ4uePgDTfH6OGtiK9Wppbp24i7zD81
vKzVtEL/nT2jdl9Y1TZ8kLhaOAzaX+YipgPXvbjKMzboxoBfS1UCsF2vlrNhXFzK
zNjxHdGn96UhjaN/ENp3bnvY+OCwdGSGJ0Bew2IqbzpWBQCwwJsL0hLveop+b8Ds
KTlOkBaZsPv+azTzNFqNg/5fc5RLHuicfzq3LBEh9KxV/XLO9f7bbCWtMZD2Mhm9
O3Dsd06AiWCA1rKSuDsNc2cOC+09Bx6Q/6Vfwh5pfP46PRZtt6UaNcBoqntubKKy
Tmwu48qF23vtZ8Jny4iuFKAAHky4YB8rx8F0AakPyrm3uuoZAMPkq87WLO1T3lqQ
z+tyE/asDztrV3yuprfWhtTyagJPPozpY6sIJ1VcsvkSfa9AUINZx7uvBXI0oEQt
tIaBj9hVJgUZ774shM1E6OKKEcVvBSPiMrCIuV0CaPWFKvKIJb2qpv/gUxvAg///
SY7So/+tgvV5B/YZ9O/6Dq1KI5VPdfYL2PQdTql7SOQRTBmw1z8lpulbKMMtFl8Q
RmU8EluNQ0H3E1vyrFpCg1m9UZjAuiI825npQZlg8P3Qo45TdfZHW2owvmUpOr00
1fJ+0wYGLDaKSDd4jp2rMnL47hi62dXPQn9qhCqYIrm8DGwnS7dp7vbu34UheulY
vqsXw8sD5zlEJRJ12fi0nLWOdLbYXjColkL7x6xcxEZ33UAJMFlGFchiE+mnXEKF
BPGFoowc2AGevoZsl9avouAr0x9LF11bTiwipdcksVM7oB5M/tLIvOuwnOhPhmwR
vnafEjUmwIsdDt8AUUCMDYdkLaKqU7B3xi0LiTNbrDzPz9wwOPg6b2xvMhD90QYJ
PG+621uukwKAq/u6dTOrvMoRQxxSS01XcKdit1JXP3+3664mrj/F014Fv0LcimGd
eEYXbUlccP69IQ7AemZjKKssjc5HltRCFT84EtxLu7EqguRlF12TzX65jOL/Cv9/
QXoMseBvmDXpY0cExvC/xxHw/KMmRwvRNiGcelYtoSK/7wzJEs+TPH4PsuCE6LBn
0s3EMsapnDAKHnFqph3+N8szQkqIfGETk2avxpl7kjZRsCjPEXFWNVCSgAIv/PM6
lxAkP6lY9DHSCaPOL5yyRU0yLCg5M7UD9u0BxERM2GPW8m/4DIrWhz3JtW7/FKvG
Vr9E22BUDTLpsLwcx0T7d/23C5hec915T6fmJcqP8HY3VwRd3TuBmbp5HwBMTpBy
mMuss5WwwvYBJOmjyYGnThamevD0w+sp5fJ8gaw7/0sBfL3r60h0rHCBhfsEIIYU
Y1iEkppbhQfqaRFRPCbeZ4IcFV5/HsLiJR/CwP5n0p3i1uxiBDijondesiXK0e/2
IxhDXgi1f8/KQIwLAQLpCHnheQHgAhU1z2oIhbV4GroR2ZaJ8XeGPHsmEl2Jb3CP
Tk+bgIXmr3G/UfyOpaGfjRSzgn3y6r93kQ69qgMU4w5Eqka+RNeNMbK8P5OIQKW/
SWavi1J+sdXcizZBz5SdDZXpjAjs/mfdismEVJsfKmGDb/AG8YEa9B7FF7lRC4Za
649qUQPQC3HEmTekcGucsbGMlr9ZUn/bUZXFZ99kyl4TWlr6QwiPKR7Z9sNrPifp
FQdZulvl+ZSXzSUuHdjFvxFvvbYwgNhas642KsEkWYoMo9B8NWhdky/bySz7GUr3
zDXQ7zIxbSxASLdg4sTMU+p0MbE1FdYH8IJQl51WtS+wYiXWmfkgEqsvX8QMMcGO
j77eJkaUluTegEdsuVLfmdPDCNkAobytF7sqY/4CHC/F3nxu6Bkpa/YBjK4Us+nP
gHNRudpfc7iXoP1vAsynUcB0KNEaVAh7UsDa6wN7NiIkqsGq7PJTV7/ooqsvIPPv
yoXVPRIqwCCfKyxhf8Q/5LqPLuxnv8uWyJnpb0GrsTtTQqky15U+QQaSSKi2Isnm
VThxw6TJuqzHNvPxV3L0X2h8lPZZ75vbZEzQGVSjIF0UtK1nLugYOkv6/RuOm0GO
Bv7cRgTFLCuU7i6NfA37fjjHVAIvkDNO/8DQ3WLuvat1MT16JFBUsBj2EAoL6Aoo
7G9Ls6Mwr3IWeCus35ipNlG0B9oyosHHsgZZa8fZ/dpkLRVlXotbNI1rK0ovBxLI
Ty4CkNbWQNyDftjBSpPrehzk8hK+4n+L7QTRP1YP/+w0VFL82uD0TVTHpjtr9k98
aDQaKW+/5M+WpusPjr9pDq3wej9xh01XivOg/Ro6/L85Gtr9r/IF9jXymeZV8PX+
vfjs9+bkBYenF8sPzO9Js8N+Ji8Ku95i7QEPyOdmo3cjYOHS++6Cr9ukG4SviWxx
V6lYIyJPX9JbnW59ByVqHi5eEiQsmukYPZwLLaLXJS1fPRum/KsfzB8heShujYBR
ja8R8bwDUfMgb/E8qgzQ9chmvrvkcf9nh39S/ocy01arZLhG6vdT/gSFSVmgwtFp
NJixaNHzH7/6Fd+2Aj43p9sjXH6nCQ4rkcETb0PFJjuOTWPgWentNTUsELnaczWr
ChRFKxdAKmaZrX/JtG1eips0v8bj9sJkeWLaIcsGSS3Wn4YAQcIH1lj7LADeik00
HupifvIVNWTyDca5DPPtWrnbXxAJJIAmub2Ff7dSybeVbc/TfeouZqZogOBrBvQb
nng03EzLxVp2lbzzqRUVNZ5PIhitvSk9bQKLPjNBmXRV+MAcjMcMz4ENDAVDjxsy
wvgHPGlgpbLNd3NndDOtV1W/WT5Q/hWcEZzGQU58fsJj9tt3mEBTgymClfkW0lVX
KqWpCW1Vt10jzYJbfPZ0RAtlw9/BCuFDe5qduHMISx4blzo9FCOIFsng2z+PGkHp
5ixKf1mqN/Lhd1iiOwk+Amtc7xAMP35MnZfk1Kmda25lb4qH0jNBD95G6g+yPuQM
Bxx/0yVdCXV4gKco6TyNF7RFzIOtOimkkuVkfKy0YOwBOqFA8ePDQnImmbqwzVzS
SI6FgaNZcNDiQ5LUvG1lwvh2B4zIR+qg/RVj1Zq/jj82is9GTbj75+ZPEee6kC5h
ZLgAXYazlM3oKFOyCa9DdSwES5b08q7E9lJ5sULBanc257Tw5iv9aqr6IkS4oljn
YAy6RrzLYzOH5Pw7aZEktUml9B44m70EHGqsUx7I/p82hOOzip6GGccXOTmBz/KC
o56TtVGc+kQM0UoWHmL3Z1cKxoythGtm28hia5wjelEy5LZEkeTUiC9BhjNMRaG7
t4ms2JDqFTj+2b5DHWKSiH9wf8CypamTLXioWZyfTWCoEoq/EZjTcDYPoK2IhOHr
MWcduGTiFCry96MKavaq1ZYMhGOKa7pXtBNeVir4579yZZNTqIfXSA5XM3Jv+kjW
epr39IYA4loG1vWYqeTDVjJREa5vFSn7v56zpblIbFpfj6tSIY//McUAMTpoWlJD
OPpbIxvZAHAX46WOIsJ5gZrh/Gc2ZSqVi4Fkto2Tt8F/UrwWnXC7BrT2QQizX2Uc
Wd7N2GPkeDdKill+CuMwIczsVxWr98gm23L3Jf2EHzhU0xSybWFbVBqG0L1LmEUx
BjsPLZDvuQBVac+mAfp5t4b1CqtNnBjNFqI3JXtxZ38CEsyq34wrQ2TRqyJFvS8q
qdrA7P+i+cfEWniqY9HsJNZeeT7AqyiHBP0gy7Q5soSA+DltmWchXfTPqeJnMZUQ
u16+VsBQUzCwZLNRReqkXpML54JgqlcJvMKRsGSwMKa//1MGxJA9p+hgG1oj4XTs
+z8j6bLqNwPIsywjGT+1jGBvlpO/pKYLexkueCvSbJUAbJc6rir5fI2R/rCTZGO8
WcVbIuUSDvLXr80sIZOZT/3+Zj9NVMpt9+DNvuaNck5YsaeJlEpIltHqH99RPtOv
irRxicIBaltHhdqaQuHZzGWCVldPrCKi7pQ0NbE6v3nwTignzBXYH0mw5hWFzkkM
3xnu7THIeRwRrEZkYK7JIX4Hz9fp/KZ8AVblSh4SkW36D6xAd4dZz9kLX72+902Z
fRSlybgc+0o5Qh5TH/F9ouGsGIiJuNlE+MnLU9ob2J4mRgMYN1F6+WoRTrAFZ6F2
gF/QUYkSd0gSYGexBacWppxWvmMcm3wM+zh830p7Rm2XrHu+iovdm/uu+rxu3uls
h/1vrIadsDHex5tBy1g5bpxwiBExhsb4xtiLeo3XqhT38WkXgWk+vEHcuaYZx6gb
lmWeY2SjeTXYR2pkmPLFgQsXMfChyJWkP3VhcrzTc9M0viThZ/aCPDp3gYz+v9es
knolpqyxCa/iEUjRSePJJ+SQwG9fdGInErO71B53gYGdmbYaa5PYtbWJrrETQwSo
85xtcdwFmf5779n9KMjNUZooejUzfGotiuj/MRURBv3HRFes9F14Hg5lckZJzFxk
zc5ncFKb4RrtjEL9tqXft/NKy7AK0vskiMAdk3ISO50bX4cOsErTg6oH08RgWXtK
1lFxCka7pH/3HaDWXqKYve1W6FZGV6y01t9inoOOs4VZcCvyWofJZRH86FCpMC9m
qoZWCvC0GG+sR0ockrZdQQAsDIfWZrvlNEGKDc/TbshjERrmsJApjlvs78SmfPId
jGVSkANGEvz3oZHApVAsYFBTaoGKphul/W2uMaWzY+BOa4Q0gcmmFDafJpBMs097
AxamPaoBWBPRuNbVTws8/cUGDyxx/ZpcqKkNRldRTUd8aMfGhO/dtoqOoVq8pZEg
XsrHTCvodkrzh+XNe+4luv1Wr5dKZVBOWnu4jemfY500rhnVccuKKAYBevV22eQW
UclPFgnjZscGk96mnqF1Su5ubOiL0LaCtKKW7BGwJS27/6P7s4i5RffR54Xw4nbT
6GbgqT/L/9+zGnzIMOHLMuXlhLPx5NdjKmexKeijpIjin4A+Gxa2TeGJ9n53RZMh
C/AlWZpXrXmkTCrFt5NSeTOQr/41/E7X7enzMYHt+QgcjJiho1hsbNdCjEqEOqxa
cYY8dypUNBSuRszsFrRg//m4UsrRSLEgBL9sW3bOzJpnfSzvfjTRFMVlwXXlW6N3
MK2cp2Zh1KQmiGdCdmBV0uy57xEZG2ccgmq8C5EXKtbDqYsh5xewtqT619J+QhEK
R6jLJ0ZXME/kWFm8+mMQVSCxCYjZA89RTBE87ED7oqUI7aMt1TX2dpR6lSLcEWtl
wlNnBPqq6WEChqDcswp0KF9d1P7nPzP8BH9pOhEOqMSr9hhqnaXuk7HWeom0bhYw
dzx1fSwhJtui8uW+BB7UNfQpviIMMGwxiQ49wRkpxNWynYqc7gsjbs01DIUcvxjl
DrofXwCT0IU4UDfN2kPzqI/vcxIuV/kOp9eKUXDo29Fri8xfdXt5SULkjt5yCfnJ
Z3YmEDYXaB/ETHdJs+DRQrzz7PZR1M1+oyuRbSLJRSaE+e4NZZoOPE48Yt6H3tiW
8uuxUMDQAid0nMpEV2Vvlnx9XK5vZnOxxD7DCh238MVHIwDSCaK4TdLDQKKOAL6L
FCcMo4EFNELWpbIsVf+cKnOIoo5fDyo4aIWPVS8tDB0dkfep11e+wzyl3Bv8H2o8
LYHw12c0OGH6mMbA3+mcZablalXPKRMblzxRnykJ9HolyNqxK/PhbchkUzsz8G1p
UY6XqnT2rq2ViI3HJmHQ5/Fx7YGx4y37+Yjx3BcYCx6B5FwoEHM6s8TkXKDVPPsW
FAmvUX39Fib6DjeMdISDUD8KQmDS2KtIQJ43bA2Ihuiq6YGp5EkdX/VZiPk4mEvB
xh4qA+gGc3aITVW0+r+KOsOIj+0UTLksR5DqmuHy+ioP+7+D3N3GEFcDWmgFRHi5
WHAp01MvCcSTb6Ecyj6/yH4Vv7aQ2r35HwsNaSTNtasI3USQeDz9w35W19bvf6QJ
6d/pB8jSgSk5rvGxo+vSgvZ67SSV46fpPyxP8jMNj/U5haIrnaCn84h2Q1Ou/XWJ
j/sqICIo3DePhbl5yVVVE2E/T9Kd1Rnl1gYmWjvYmwsWKQkcj3mXmg42K13JYeCT
L9mqDPY7LnBhmflgKCc5CQRJbVXyhAWziw9/BwzZ8OPHz7n6wh2aZyi/jPoomcMt
uSO6XcQ2N069b6iIdEPCY5nwA2eouEyuhszF6iJmkB1MVtB8YLyPyZZoaMbKdT8b
9q/ANYonLV3xZtCVbJTmgfb5QBGPx7Kuos+HyPyt2hBuKIyd8L9Ff8f6Snp6/jMY
nhVWGVYNKuSk3wBUOuo1/QBHzDpCk9PHFKO6TXtt0sSgoQMQDuJgMvZ3M3jB832G
vbK636RkltEKmYhCN2Owwoyni9LsUUHgLf7GmBKkc+dNpZre8T2PJIWuMlTG+uSt
Trmvn3IlIqRCgphnvJbf3v4eqkT3IJT2w2Uo2Gf4JIbtyDDZOuq9tqU11UWVkXsc
fvF2YmgEHuQwzjhOD5NRzvhrPXzAda4953FRY7bR0HeuGzZsyNdl7v989hy4vl7x
SXN8tJcqgl3z/oXuSCWKskZ7fs1UFlekcgM9ZWAZKF9ts8APsCjjmJ3hRfRUbQMU
u+HzFZ4EHkeCn5VWEpowlW1hPhVgLAiXcBmJFGSVqkE+1+7bNgLNxWUXcKQnmItL
HOx2FRKwNyjHXiIijMm7AYL1FwNhPCqXSdQhyNGsH/RZ4qjgjtb0IkpyNMuiiRhl
RtnBpGNQifRPJtNnQ6qEoEt3B76dDU5wGhjWPtK7dErILVnrAHw11EbgbpYNQGfs
5vaqPBuS+PgYKny18if3GzdI3d5G73BFgIJZSNLjqgCY5ZdjkWQY864eNteB+vKc
A+C7R718KM7ruWYEX7bOJun8BYFsN4C4IpmLg0k1lDLS0EOeyWtLmflOZaC5J7H3
YacG/e4+Inse8JtGJbN9iDQUoJnC/cHJiWofmlWE8mhe63MYgM4nNnCU7/O6NarW
+FrO6ywTLr1xu7KFm0r/rNQoInWS94C51H8rgIzRLMqtfcMNfjGV/GXsYy8uiqsx
AwJzgrUrWrS4XxuBO/hVPtLx5Rju6J7v1ulzhQRilRXq8isvAttVh0OvkxsbfQrY
xhcufatMwPx88PnmjS3WA3GR3J/u6C7MZWcN7sSebP3EfIy2WmG3q4htEfA/wc72
/JWx21kNnolLCO4O5ETXlMwFHMbBxFQ9SdxM5DZsAmubQdIeNIQIyLNbzc4RPg31
fqVFH/uYtNqMfmzUT+bVhKCUgJH6QAoCFPT2LzLkkmBrV9kk7spA6csv55vrrdBt
5SDluSFP0QdAOsbjE6FtGiFca2hNVPRpL24VkKb79WLQg+/2qnO/74gP00YCVrzN
BRql7xSRGNdNexx1bgL//QV/xAC6rvcRCwj+6b1G5xRV1g9yL3cb3ax6q74CjaPV
XNq67Xy8l/f4DopJPx39FwSx5VySPK6fhXYOFqeqOPqIG8aJmjFSiP8m3Cea4lBo
p9inL9UQctw/qFuNydCRjPEPUi9uxFKNoZMtSFfKElj2a9tiX+uvo5lN35OKVyEp
qJwYszgdcXLQVholqVa3OeutDN4k9NP26dk2KjIp8rGeVAEhWzWHBe4376RLhsvb
V/Jk2qpZGRWRDIUSPuahp31wYPdN9WADqG5FWwSf4qW+WqPnu3ZeN7Zw3UehvcgN
TFvlGTtsfZUFUjSF2ppMigMy0mvdqtPKNFqf/o2J3Bhj9vaS+aNj7ehq2caVX8tO
sP0S5ByLbFkNrb/K7d7fnJaCjAPezd3G7FH1PxQTAQpl2qYx46N2eXiBSbUfZpZy
e8ZTY63JNXA3cb4/czVvORE6xC8WJQhvOJ8UNvgyb6sqM9KPSz89F0cxaV36DjGI
a3sBObxcfxBrAwNwwybfu/zLBU7YDEdR3+dB7oXZAxP5ILOewlGrhhWKJHeITHIs
fvKZ90r4BGoXrQu7jz3FgaVkHMTsVqcJhD1IZxhFQcs6Mvr96jOTh0Yv7vuGkqkd
B6Lt3frUHTtYjhfv9Fj6N9F4L9D9a1PV6jkzw4jxXn+dS2fteJn3IoDcThniKrFJ
qjN0GH+lbDCTX74N9WmM8xW94ajlM3uS8Hr61KE/wlBKTksG65lBlG5M59aEzgC9
zlTjuTMN3ztVUQ2n5qPuD2HOdqK9REbhY5OHv5jREEYk6gh7GDMd5JwTBCbCpQmj
Sin6XIbxyIrQC+WPVRudt7c4mVyaKY7ZvkSGVj1pebd/jQx9wiA8wCotxSuS12+R
bb4/gUbznWWcqYEMLHORXyyM1l7yfkqzUxN9nZKTvEnHgTUk5aG+x+x6Ra2LDkMN
Pgz1t1vb6nPlHQxymSPXOTM3MIjJ7RjYlw4WC/YuCGjxPdeLfl3FjWPRKYZbkjMQ
7dQnHJRmB0aO25a94JyeamRfioJ96L7+EE6vDs62vJKQT/9nzJPhLrLH+PZOg8V8
L5WKCX4hDWyJRyps7Cs+oqjPRwTsyTg3LUnoBIr9euIX/6jb4M6k/cgrjbmWdPmg
wG+SleQhz63HPwEnhJmyDq1m6e9HtpeQNeZgLG1K4p+QT2bdK5A/WUA0hPQi3yd+
Yrgo8cLYj1nYBMfR+H9PRfIUZQRCu8WTZbSLI7N6VziS44xp/cTezNVzZibqP6L7
rMVmt7kQXu0M5F6FpUgub4xT+QA78QAcnImhxdu03ARaeBui/0PmqClwlqevukGX
Al8GJ1xKY0vLItgaC5uMPfzbrQjvZ59RX9MnalkzbPA/swZDyNVjQ4n7GMm+uh/V
FvD9mOldrwZ7PimZO9jRtTlHRmt//VPZc9CcKjRe3pCeXz7Xk/DRbEmf/bNdxtGs
sjKoUYxD6dCvUJyWWYaPXH14RHQTQUQ3XvW6mZXfe2gVjbVvvR72Z7bKvzb0pmmy
MQWW/QPtfECuKL8JgQZ1kNPh5JgICpxYGcZGcek51LlsNlzPVNlTlwgWDZ/weXEW
Hhup8RbhI5ax9ie6fxt4DM4zKeTZS81aCJXtdECgzW3H+nFihjsSTOAmEjN032FQ
Mkw/2Ie1nAzcwyMjnuRCkn4q2HiaSyiUbJQUze9xaeQN47N6ttef+yZdS7NUD5HJ
j/Os3LTo+T4Gd2Hm+AhuLypjZUfU+QRbHZ+Xl9YfXZBHA1Kt4dDDvqn2/D9rA5Dd
F9H5mLIfeey8g8YYrrX6feyiAZPlLM0SCgFNllCZuXND9BZ3Pt+OuMkcuiJCxxFg
thJ8u64FXwiRC49s4tEXEFo/j+eFx73LCK/LVzrzqSt6yQuY1NQ5EtsLo8x+1Dtt
dQ29hm9266PzEK+yQOT7RL/rkQM+ybZ2y7vDm7OwwYWeAnX62XkwRDxxtsbbigDk
0KF9eqA+a5qz+DxS0327fgliJsQiHIfUuHilR+kqIfHkaVQOvxkAkO9ZnDbHbRq8
11GoyP5iuHBuhe8HnumDzhr+anNHe3SqO0DLkbgdfxGtaLol9Yq0N2zh1WpJUy7G
WFH7Cz5lBI3oRzmtPT1JNB2CtYuCXB5KH/ah+hwnEGznjbzeSWfKgqL4khFzva0Z
tAmXwVrsAP7GZ0s3VWZSS3L9h1g30Jz3R5f9S92WSgYsVWxaeHkGHVYASLdpjxCg
T2RYI2YLIUt58hF9zrgwxGguIUXZK9Bkm5cgGPId269Y0S2lck1tzzNo+Pw+3eS4
BbWMuSF/SbddX6cLk9j7BT5HDI/VqktBbboJ+KmWvpSbVgQ5szcBV9vRkz5wk/YT
eZFuRHBdtXK21F/cGr3G0lgtAJj3m2xefjjVTBqs/noZPWvosyppVYbRB1BAofND
fRZBLs94RMbPtLPTBaDPzWXn0zeP/vg65WHO7wIvS7y3XIZj3RPh6XDXeYEoLxnO
EghWaDzMlbYHAGlZWO/cfujCqGqtyikyIwlsu4QQ+Dol4g941FLir5SGXSU+PtjY
g5LE2lJSPlxSdZshzQ4VWTbqhyFMHGuLsWQ30YEM0zdpsbJMy+EUcNPH7c+aQJf4
E7Kyji9L+mwsq3iPNa+lV8cUE/nOEU7sXz5V9akavgZO25lo//9HsoUv+4gLMeim
sKvZtqvENOHI/MvprLsZF4UDxKQdEyALTaChCamk1Kz5HWjqEuGlXt0nLi9+UeNf
SypJgtnjqPEBNNDy/1R8rFcWs/bVBkgkT+8STk6lTO9sB+qYTEe88z4iYVy/P0EE
DrxolVwZNx0HDwwqNwzMutc1tyhFjeMr1OeX1t9N5uMhyfgissrKSRPeT5uI4to8
8C+/6GQYp5XvZdTq6LZXF99MAYdOaOTl7fy8vVlXXQbJNhmafFJusoQdY9/9q/Qw
4l0k5E8IumZqd5fa4UaOnbKLogwqH6q6e0p7Ry6O9bTnae3O75t/vuADAnVRiAUg
imOkwYUo/5qQ8iM/QTfhu+YHuQpNbxVh0mCg/2gHrnf3GntGXOdzlN/jmQW2DtVo
8d22SQdQGSBjbgafmMgflKxoUKoDTpQnXTPGEEkMUsUDUe8RycJbm1vfVmXJ64pN
UKp4F36G5egUiTbtj4OFmiG+mTBpY4UpaXCkVx/NXgOf5V+OpndajIx2GeSyPvl7
DiCzF3I3+lfxjpAbmLh1ICFelbnNY7LiDLupQFlIoZzcbre6pnLMeFNNhlGtswP3
bzhyb4p0CMxkZmcy02K9CF4nbH61fA+uOr8UQeOD6ZF/o2Wi4J9v2UX5nrRIqJb4
MECRWP5nfOpRb67BtNrauTjMVNsGmN4WU7reopKLThy25nIxcCc6s9PkcVJLsbcv
yrnEW05JIrMBMFY3p45d2e09P1HJn1azKT3Pmx5TU5vWXRS1bSNZ9DBgafS7V9s/
8JaUc7ugxm8FMvt7h/gqZxiSv17xtNqGuCSNHYuJnpcYu8oeiouBvo3VvLmbqQE4
99gzE9l9k5JKxgE5nHW2GnqYST0KkpR8e84/8vcZfs3qNiqkH4t3sjXAspoqZ8iv
xp3KXtImXxnYVVh2hk6JFJY9ZOqwZLkrvmlvQfuHn8d7Gm4PGRnCgCr0YESb704e
/fGK07lMyUVEsup5x2jNKULFKMhx6TiEbXB6psLh2vCYj//4LARMaJ/4Yb2rK8tR
3l4h8EA3cmcZT37+vq+Hwi3J0/HS6uI6EIs+Hs2RCi9i1TUbnjekZvwRhjprYPex
DCvgDsxKXCDgzHDtb7kQOAIFcnOGJCX0hILWHh8adF8k7ND754sOJa16rYvRrk0j
bjKQgFwAnPielJLjiSlQZW3rCcvMQZe7Jv1pIfLn1VXORZLbLrH02nCtE8UWGlGZ
5nT9IXYyHIxVSW5xEvNrtcs6Rnxd6HN1IiXqOO7TVjLahr2mpnZqLz4OzufKdg/4
t6uE1+OY+eW3nvGkJf1SmMfylK+U3vUVCaQelV9yPIJCUVgaW6BPhifvb6Es++kQ
5OBfRdJ+IPmFC+lZR1XesjR7OD/kUVvlICuc/UOB+veyowbvlRxIyHJsBv63uYV5
ZV0l/l9jTgA5hF5nSfXLioxowhkJqREB/y2/Y5W/EWJ5Qux7SesUM+zDr01nV0rh
ON0Xz0J77/K/lns4uRz4keHF5nwiLgHygv5l7RnCciNI/r4PRkHkp4DQE/DFqxez
kdo3LsMgdxm+igThS/c/1AGqXNVG6RY38q6oNa01iSUUEbAWbUOlqDatCoFOhnKH
/u17C9B3wXPFYew8YJfDV2f6Y5llDn3oSjA0MIGyjyrlfZRPlqcKqK5+uv18ZQcD
KF/nJCMj0Sm7bf7dz+YLQxfE0zh5waXsoqsVd0FxuYenHpch0DpbSqLJWFUNU38n
dPb7G7BEkmX0quG2nO6ohMtiCKhuZvj79UuknONZfCajPZjtbN6XulLchPKTQew3
fu7xl29+oIas01aY1Dr4kLEfJFUzW6sXFldNejMWiuhTVdEOosbbj4QF50jDfGU4
mO0aM68ZEMUXVi4pcXiZIxTQWdhRUWEM8i/sJ82IWoZw4XbTtEemA/AV6eQJBK7z
56Tu0777Y8YVnJ/uRLNU6JD711S9c85MgHWfDHvvLsQCuAVO2yffUZMDLMlxm8pD
Gd0opR1WCXL+2GI4qJLN/qEGMeUCRRQAQMffwAlkEDOXyG2QVzw5tnq78GGvG4z9
MQeLS88Vuqt/XBLihqD9e13y5JOEfKvKdzH9PICfCGR5Poy0bYfsCUbvu3w9P3bp
Ltm/TWriwnw0DwCzNxwa97rhCHJB9O6zETim7z+tFyt6iwm//F9Z6rkNDkXPeKTF
Mu2tqKCvTjt/b4aW0r8mxSJDfj7JUgDBgEEhHqcB1PUwFAxz9BJ0vOyR3SmNNyhV
WurlQAbiLMkBybzK7CKqUgd7I4lSo8Zis78Q/U8nr+lgLy3imiqONxWDK6YV8ML8
d0x7env+txq2DypvkU/rpc28obAysNid8LWmEEZCbH6EOzK9ZfndMdatk3mSshwq
+pJhOZTuFd1MVXgRNM/0m5I83+d1VKowy1jaepNJ5a5NJ9XEhY5x1pZqeGpQyw49
oV9aq+xPfSy59Hhcii5I2ujfGHEbtxlkabyyfABAn03/Fg7B0BzYigSZQcN6A0mm
U2/sxV000b4A0OH/wCIf5Eq6HDFZPLkiNqc7tRBQktoeKmKe3kUOhElGb5UqDCJj
b9+RiGZ73cpOREpRC5UIeSBaJR/61PmfFN5RMYCIKBkDnomj6dbX2oqFHyhHp6JM
refbbVG450dLtizFmmhyZTsy/ggzgQwvNRGta4IAw5b9a6c2+2uqWEkfKgS0PONw
Xw/2n21xkhr+yl33JRB1RJcYexUNpYhbjMl4jwxFix7FNJzLxr2r5EHxut/Aia/H
aEqdi+3Am3UElYyiPkwVq3xS3X1m9r25SahNHvOccJLDO360mBjIZxkUZASE+e4a
JZtKd+AQLTKbNT40DKobfyh5h6GdxSCX2q/DTWjEK+0X9csOSAv5Qn7zCCBRzigG
QbWqr2vz1vr7QYMcrBmsno601RL4y1V5aeu8d5lm+gx2I34JbRJII3jyi+f8BayJ
HJeAYMF3qJhSGOsDKvuZ06udoTkpckxLI2NDnAFH6ZyFy1i3AV9bT16ass/6IGF0
whpyfjNcM/5g6PLvwVQVnhP9XcsKWb66uc8uuhSFOXU1tbdU09JrNQSj0WQMsVTM
cs3mZz7YFljDpE97Cfs4hoXsCH75uecMRiVYTT5H1uwZbW8ave+iHMZu5EQeNK2t
U699v74hmniNKh9ir0653AN/ReY7NIoG8XtHe43uDKP8WwkjItqEOXnAbm/A0hLn
RvGrZ2Fu5EoqGjTT1UqUjEsiCEJPWx+lNLYTAi+cdmQ9648z0h1A/9vjGc3CnuaV
3FGCuh9vEL3WFe54FgEbnIjgkfz3rF84uohC0fPYi6W2lYzPdxE9qK5j8eRSP2lK
5/KxOEUaheF0nyWlxN6RPWFHQkC6kXR95Ek3SRGYYt1AFv8knOc6BgWNK33VWZex
AmLX37pIEYZTvpm1q8t2kuxPMRVDnDVoUVZrmjyPPDj5dyLyKA9PX3zWhucUJRHq
ORkZDRKxK6EG3EA9b5JNhmUnWPl7fTxOGhwNvNxWkgZDzdoaJNfXVjW7pRIlmJKT
pWTA7KYXP8FQouliqC96uPCnQgqJbMH6LYMegZOnsLOHgz3rWFmcHeqlEHDIzJzY
z9L/wA1Yp2vSex2J4DJNy+dLUPoI7LyvkqcKTluYLG+3zQ7lfg3xIN4xY0+ouRID
1QGB3gC/a9fSHSc6IfTXyyYaquTegQH28EqwtpnbcWRoMCOECFvY0yaJPqiwiyJG
2qGz5noNZdw35/mGY9I2JSy0EJJMrV15O3q9cruFmupdocrJ2O4YvxzIWJYR/yAp
oqgRW5l3kAcStgpdF5CkcPM+wHg6rTE3ktDszyJAPOk5+MvvPpI5cl7l/uqgchVS
pZ83Xk+zGjNDsW6C7BXLu/2LC/H6XOwLT1Fz4hO6wxQyb4QoRRp8zy2IUXUp5JMg
y9NdNP6q5wszLVwqU+nDzwgXdW7VxXy+1ARcvO5bEElePnaDJcPo2LgGZI7lu9xg
Qw/pCVodl/gOf1mi9qwcNRoqUnGlc31Hr1XOM21sBJC48yYVdhTSjonHCktNs5C+
JhAi8+HVuzLEEBjYY5sL8MyPdnHu739i6E272P3LhfLptyKGqo6JnipdTD71pwoX
unwM8r1sXsa8IjDFJsJF/euiFAUSsRpN5HsMGoDgkQk/uB2cDgt7Jm6KC1OcXSUq
vV9CNt50/2Uljj0lhQFzULWQEY+pOeEIG2G++bEI7PK6GXif/TJOfkiTIQj/Gx9Y
NJCmBagjEKMNOEhCT1NbFK0TDgZ4Lo1qshfvaN8dieuLX6F8xa7DUmjKJ/bXeX4e
yEmtg3gF81UayAJf3MmLSoLKRG84SwEiKNnBAStZOlzk3lW3pA7xHfVB9ziIIoQj
GRGxXzHAp3/8FAJkFmf7ywTiFBIEAvjQ0cAqhBuYpnrPxYtVDoEXHzG9npBZZRYZ
b5fLFG6jHjHkpzA+SWO5vWjwiEdddM5q3rJ7/8HM30tpAcA2gY6KpZtuEZIIZIQm
+Vk8tF+XJucyHywoiAg2f85bdJiZLCKV6bs5tPVRfvD4l48cUzbtjfXimmYLoUSn
7F/vzRKpvOrvPulbaZl2SWtFODK6rVSznbJ3Jm7Q4sOhwYM/P3OQoeFx6CUs14/R
G2dFxhinU2UtEHVIdRJyDwmCZhdfhaVn/gGXcgLcuII5DvLbhBqpeB8Riahtc7PF
lvZXegVOifrtauKzGEfS/Rv846aez+tEX1ghhVMdEBmE8gn5sp+UNp1N8HvYR/0A
QjNd9grUxzN7nKCWQEYLwmiFu0FBEh6Cr0FTNrSY8IwayEWwX08O54ZDG7CYho8b
ILSbzcCLXgG/CI0/V8a0jU1yfJBc88ed4udrua0MsWdMyiAnlfu/eziYWLrmsJpG
gCbRopwqk6oqQq/pi+MRO6MlUY6GOHHRXeTQcEU3ibi1YDoxp9nqs4x/qYtTbLix
RmNUl4Ru1ps2d2u4z5hzR4GruX3my5mmsW6yVwwj8w3zzTTAP8HMLZDOdHFvBwBR
fLHfcldaDsDZpzj3235s3Bhe2rBW6ibTy69XVD3RolA3AT0AohTlgBYoa6dHwJ/l
1Sp6GW/cexabSc1jEMjNGTRpVniJC4R2y7iQXfxY63Co+KD8ForEUxV/JXLMfVUu
UjShzyX8aHto67e+geY0dFG1X/8Jg8th5z1SEzLGy+ppDJRgGhL0eSuDYHKpEvNz
UnhWxkO6KUwrnrm43TXX6Bu/BUUqxQJXC9V+hz1L8KeunT1gl4N58N7mDsgwJD63
XLON/7/82iZKhJ1RWB9B18Q2AsmVGSxqcTudtQNIhEyzcrWuu5I5kw7YWSQu2Pur
CGwlSsI1p3WaHJdajMTmR/6py3YRMxSwWKk+BBnotr4jWlKSUMp5XXZcPk9xkuwV
bnmgO5w2TwdSD/4bQeP72Kj0OHgwfX8UyzNIkMoMpkh5STntfAgtdOJTdPYVgCvo
/dzJtEMGy2u+/c3Z3iET7vcRjUzAQ4LebhylnzClvCjR0pCQFTVqEKLcR42EWgSj
gLgrSApRs/Cidx5VH5gp9FMvlATXXY8/oU7uotiko4nHnxaDhKFWJIOj2iR1P7Wo
IE3DrRotU86Y8IUYsoNKS79njTp2KzAG5TajLEOYfMlfZO/nGMEAAWQuNeF2OCDV
VHWcqh/vO+VeifqP/PM1kmpeNfLTaG0cBGq6Dz1GqwEw6cBTAPfiSQOLXc+6p5ix
tTGRWiXNNuG4rAGZWZa6YzP1WqPH+vw8p+3XcWx6/TZaSx8ZAQ0HJpTZ6jqQFkXl
m0NuVJguWzISh1mKpP2NU4XomT8y1rv6w5Wis+wLQiei01HyELjaqfYQrcdh9BgY
3wI/vk9BWvF2YWbHpCg6F/Sj9aWx8w9n0VyeZhUiCP3e593fAqNrbpLT+jDu0tdd
g1tLRCeD++ZtYZ+M7xKjaR+Rry138z1hCaizPXgg0YNMgLGlOVeBDRYcMac1Mdzp
ws2y8CQE9pCcEQ2iAd1wZWm2IbkG/wqX5DstH/gkqyZl/lqRDwFQgrmYwZLW2J3Z
t6OxHw2ETuelqK3Ly96wtS4+6gZj75BR3Eezc+hi8/afDowaVkn7lg6Ap0ovo4Ck
k8h+myB1KJP9AiZeNaGV+ZRKC4Odbwo5rfUypJiz7xzH/o/k0T+wtxydOElXLprv
fj51Tv62jrjKSus0uzZOI3DtjFIf4GsMXQbbzZeWvMPC1JAq/GJ9BBQZDc/pD4Nw
sAtxZJbeTGNjyWkwDvRYItF4QWVPTOjeBDVQ+S3+1AYMVD6c8K+g4RAhcAPKh+ig
xroYZ8NIbHUvuFq6Uq/7ipyAnmGs2OuienuEFKXOkirTaU51O4qm+grGIGrwGxtK
2MMGrYJPvhpNnPrcVc+0FDkxdbPtG+phf0zozBOH2xdfCd8VjYhksfxULTO+9UgV
ayEjhFRAc/Q9iFTj97/C/sE55IJeGszmhAAh6tmZvv1oAihvZg49ZtSdw0H1lhAk
g8FV2ZEfO4lRjw9vqLcVWTxKPy0fRRNY9bU0sQhKbR+V5+tD04k9Yh36/XgYVIcT
GpYA4NZWz5e7uHI9hA7sYSXuxyOJ+D3ID/5DVt//iDvbAcXfZTO4Fyqz/jQlgKn1
DBG18MV6B6Ze1xMTCutO5c0fk5e+qgRvzt0lEvR05GlJs1MAB8ljTs0Z6tDzdovW
b+RxyXVmD5eFASJFn9jNQ//0Z7ZshgpljkA4p0xpzr+qibW6F33C0guDU1k+sXKa
FpDxy+dRSETH7pHTCvaYmpnTLNCiM/S4qcevf4zHnqs/efV+0nPRMkNf90PD8rj3
iBwWAPgbtFFUr0i3hDFY9SIVkXmGkryB8wR4Dw/tkSnv8r7MocGNwswLRTooxprq
UlEbCbnYkcASvZ0GM1qfnh4f4qdq5IkAJLYbXiuK/muVIORF15f7vEdgnS0iGn9U
fj1tbECuPNnU3Rru1pdY75pE70NzqfvVIog52wYQpuxCWUM1HqJ0pTgMkmkJfSA3
uRyXFnVFOSighez/Y9L9VCsaFQYW71JNqGhpCBv+p1Kzkhp3ten9tI2Tv0oanrYm
p0+QVpsSmyByttPbgLN1fHtu7D1lXFJBd8jbB0ClBNHu2Cz+4lxtGZ2CCsX0i4s5
XEcuqVTg5s1OD0+5G8KHK9e0I6HE+BLzAoLNjHJXghr5Lk6LyE1hAAeZZTPB4Dz8
O44X4lBS71vQtmnT0Iz21t9Gar0Ute1cYG9V9gMWF5bOXzbfGHl3+2TjSWtToVxr
/BUJlnxBJdIX8P4Lp4BlEQhiWP+twr5EoTeHsn6/2WUbjcQqTnqYLMTYbEOxD1yO
/dYp3PgAWokD5oxBQfh+E6kGOqqeXjmGOOGtqw+L3Jtb7TPAJb25EOMuOnzeXtip
19Kn5CK1N7xEravLda2EHqlevZzPZm8ZW5eCbQ5FGbTsInsjgybtRnB2/xmLFkWX
d3uGWefKrTEEWniEM3SL4psozB4/Lm5V/ISLK8kxsAbbb3v9CdxNfHkTKv6/iMaR
DKrm6FkvITu0+z5/es+3qMVN/aiOoMn7CRXGFTHwvk7wuXmaX28ymDwU/vCbohe9
RzDkAQoBXFwgAGWrYG4ye44zIRGuBpLcc4m160Ef2z+NsUCWBrRj3oDZiFRSBbSA
JJDuobcRUsWQpsaSYgtIcFDf9i4doeRJa3FQumZ8d7q/IAI9KnOmnifnpgmBG36b
P5OkPEOZXuhIZmTPTqdsS0vSoSd/KkDdThz1pSIT7AA54+Ih7q0LZeAUmJ2CtoZy
eCjximhY3SXNH3fFFZ1IUhCguuKLXKx7Ze6t7U/1XtGc3nbnITZHCycj/02L9TT6
qPR+F1KoAMDwuC49D2OYBO56q5LYfURKEzP1v5K7rh6+Y+j8WTnhbB8o0GBsVLKO
QXvDLedlYm2diRfmQs4iEpT7m3wkCXxtOtBsoV+UBJEyffki0f3MlQQ9AEObvwIp
l2E4sKoMva/CY4qm7kjp87flChI0WR5C5RODKKERIwUe1Q9BxxsjIo5/bydWE2dr
1N6hNQdwghs4OMqgBORBcd439423XP/xYGZfxZhJ0M8ChcFslFI8vlNUYBI6zcxn
Vgc7CQZaVQ+m7LSZGrcVtRSsDTLyH0Uomq3CmrHiTa6LQlDyt3lLyKdum57XkNvO
0+SuzBbJer/7epZ1bJHYe2C8FR91c/5hOc/mTJvKXPJLslhbKgMgoxVuLgsgFyW1
GOIZoAuAtNecUlfoL9Mxh78FBhnuTLJtqcZR9DoOkTEJcToH+2o1agKiGJRB1qOo
1mO/BM6/QcGaGEUtge6ocSGnw/7hQex0vuIF6Z3bGqlaYDWoe5dSObF7b1uMOmTu
UOAbKxOQJiH1KU+UIi8PMYJck6nl/gNfoQcZAXoE4PbHtm6hPC5nGydsdAFoFk6W
r8Cc4tHrJAkNyi7gd0yyK5EGzqXNrA86qdo3v27F1mcHdVZpVk7y8ETVgIBgwiSg
kDZzffXvvwTh1+xwQo7pAY6wyFP7pHdx0SwRGgux/XbXds8jyNOHXe1Tkk/QaSi2
1d6Pmld0aKurifxciymLvAWwD9FYNdPeXzVfGxSkJ4KYn+sPPB4d6qvtdB7XKMVD
/MnFL7JOSkhmm/MYfqLFk/zQ+KoZ8dQK4WphraVn40Kg/if+hMn+m6sxOwRkD6r6
2hTLg7sW1hExhjh/Puix3AQX4qLxwkehdl7F029ez2ETsHAyPVxD3bdVQIlRPRbr
R2CcFemVV1G7PjCdT01aWq/gJS+mpAmzw59yHPJO3wqEEJbPJRM3OW6Nof4ZujqM
9iUL08ujJii5/lTtWz/+YTJLoG6foJTirup5NiYQttbraIDX8eYMEigVxlisIel3
dwYW/fcUWQIa3ndNRZN0rMPRrlwrm/2guLznw+hcsAuIvnhh9ffByE03Ae5HmXi6
Hq3KqgJefBgwKyw+M8XU8h2Al9q3L/S3+IyAHawvQ9Wd2b2g4ioKdcV/qxmJH7+E
JanVCL/o+ZU0MgG/WmHIXZMdZKG9yJ/fLPOHkIkKDvsuhcbwBvDQ496/d0RnZmcb
G8xDZxr3Y68fZW59BNMi1JOplBZces+oW0n3iw6Ao/TCPEE8ZUo9DSs1wiIxmleL
P00XvSAnAtOWJ6Hs8wbzYuKdPuhLZudLNAoM0j+7SXWsN8YEfnrjilwzcJ6nyEA8
8Ja8drB0IzjVPQtUK/Wyxvt9ji25AgXXCvStQdVmbdHqmFkblbi5xtS3Am4PSS0u
bLyvIyjo7U2SRb9U2IccS6zgAoCe03PVPENB/oJimEkmc2QPFhscwtobmtQnRt4E
ndO95nAlbZS5SMP6hOKlfTZn5agpDX4xwdYtkfc/X9Ym+QruFNjEDElfwSY7wAWN
XD8W9BdK9/AM2AEP6GW0j7LRNyKI9zuE9qImn8krphoLPFBTrPOUE+P2sRw6r6d1
XJ/tI40bn7QcNKiYDMtMTeYXj3VVFzjdidHFgw/NeYME/iYWePpqZo98DXdTqOSi
bkpfdLCP574r2yi11PlEmNJZ0Bu7Gzs3C8v4szxKEkG1exH5uXwF1Y9IRoTe9rlf
Ucv6XPELhiLmwRTd1ZnfJsOx6I8jzi+3JO9MV+V9fDpGB66/WFkv6e4zc6oHY1RT
2HndAvbA4Va1mVrGYumPWqiIW06q0VJHjUK7G1Oj1wWY7SjjZ/hS7E0yyDZ4TvdQ
iDtvruelYp9Pl8YN+5P5sKWcko7fzUsAZ6r6UaHXolUdVxfFkE2WPBIGCcUleoHX
fw6TKIXUdutNkfajeJ9+FX77Mu7QTvrx8IUwby2w7Sw06U8sExV3LjHnal860VfR
VK3a4k9Xv8BV9TiQB/c5jICdta1rO8O87bbFhUkxr9rIqTgRqywpd0ywiFuKbTt+
tZ5dgNdQjjoIgaKxiQqyVCLhQFjBHmRSOgNmhbzn69eQqPqxxCx57p3jFL5Off0e
YTXqaQbu6CUPt5lW1VE+RZt+fmOjx0xF2vwtfYckhBk80u1iSyHndtEMJXNS050N
AvoHg0wqNk7cR/sR67G/4QzJC/1few1GqyK8JysdkODHFCS7fePsZjjBhnUfI34V
eUG4ELxK2yO756ZMiIINoOic41LAZV8tM2FRPwDk6a57D3YF99s72mwDmWoE7JyY
rV+pl27WaVOaot6mLvgGWmNhE5I11+B8+96yWu0nHAu8OeQlNqDztA0OH0cHx/yE
dgKuLXOO2pbWgmUoQgUSi9saMslDyrBrSe0mQazcFw71pIG7De8Lm5o3gXdWC1sP
fR3uEU5L01kmFRMcayrHfm7hpST2wRpCjSPyX+4T1crEhKveyJ0hSfxQ7Ijt4Pzb
pBG7lrFg47mmxRV3fhUOOvUe685n3pf3A0jCzW3kjfDC4uOh7syt4nXWVTG6N//K
UFqXs3cGiP8WfZPkN3zBuRtDaldbyIsb1ZEkiKsybrNfcZgKgK6ofwRgFsTXztz1
TZQLE0+tudMAQkJqIrOig96T/RljFMfDpw+2me8Kn2VmEf7IwqE1UsR27eg7oSad
423awtL3ET2fnxwTWSCiUEvaqbwRh9We3oyYLZD911VXAGEHReTx+HQClQBKTew0
BYyci+0B+r/dSEX3ANk9bR6m3wmZ6SyHPQYNhNwij/ka3LVeoQpmUdVhAACdBOm1
adGF86xynCMOud05Qg5Mep4XstrbPqynUzf/MMo5OZ5WuVG840cV5+9Afr3Qv/si
0568Wttag0OMkXDnsv+4sLmATjRbyWd0ZsD/u8JN8SOjKctXwF8X7fcBVIEbimbp
Llox2/AdHEjiAuGBgWn0XEofrr31XEq5qxXw84szV8Jh5K/r5fAnms9KopG02b1N
Byypww007J07OwqvGjGmejeIxS8rNkrbMN0NmYL5xt2ofkDVV7WXudcGECIEmbJF
K+QNfQLh3AdggDDsjYs/uEE1C4EHnpbhwm7FDJ2eRgrcdHExr1OaV/fNbtxlddX7
WAvdiy0R9yc0CX+1CgL2sKgc/RPAHZ9uay4xwT7PxEHF88b4Uzqg3ApW1JYiVvgV
CcCKwQnCPi65ZFIrfbIeLYTYAO4tndRqNjPXgNQEfXtqMly4imUjVYdbnz5O9jX+
krlstnfwAYHmk2gyd3il4W9ziFn62U7SZXfnaoafluR/VwcUbsM7jbJeM5G/k518
fGUFp/c2ZGVp/L29ESXEjOE6BapHOqpVipwKpdYJZkGuXNZdGEsHHPAM0uLrVZx5
lpvx5s76I1JajHmM6WYC1gt2K7LomyGWEhUyFfNjiUQolcUW3BSVrfjJKwfLn0ZP
c0bn/8ctdb8GOPHcu6gZz2YWxGpLgXRY/EyBjzjYpdMFQfiQJhkYcYyflXS89rI3
ASqxvwi2OEoG/tRqwC07eZdaViE3q+r/g+H6URX38NcFTqw5Tnw9yvKcAQSQxvYr
aI/IVsOQyF4kyn/plDfLcj6r57XxwFJP9lYIK7ZEHzRlLqtHRy32o8+bPwbIdzmz
XpyXyYMKAydIGcLKQ10AXzLnhmVzYtNH6YHeIBuJfne8xRWfrIqj5ER0mx8vKA/Q
DJWkUXoZEN5Jt5DcY/26lbukN4CycVYJa+8HVH67NwdG0LxjvJLB74y1O4z9uL4w
brNf8oqZlh02hbB4Bg9uBDUxNsGZ5YUB9fL/TxaPrI6Dxi8qwbTNse7VG4IwU9fU
hmk3ULSjlaFdjBT8hc3sOz1HJ9w8IQ+ODyPrwXI8AYLKmBv1vjq8cd9kya7ezUm6
GjANBT/yad5nmJnMHAysM81laXxPEz+v7ytX8BagFGpcKCmT04pPmcq16MehdSfY
w/BG/YicPw/vskRNhb56m+pWvDqxrdLBH/NCYjbcrJXu1aGjpHx3ff6ocrBk3IOm
I4KYt73oronUaoTBNBGjK7NS0O0CbyHw8yaqV8ub+r3CPWLuxMxTD1Zz2eXFu39q
k6qxz5as3gK3CjTo/WcyyjxYqf8qaeSttXlnCzMqXrBzGFOayxWEAwWeBYpImAqz
9VTSzM3ex1H6bzzPqxK4j6x6/+4BalorMWB6oBclUdAzr+sF3g8SEjNEbYsF9OEL
LDov+KRu8nwdKkxp7ct3omOmrJ1tot0rxGZwxAw2GMJ/BJS2t7dWZ4e8Ers/UbaS
2z/dyZC1SBccKiBZ6jTV3ZioyEbMXmj6sBvQOn3jDYHu88CFyWFvfyMLj3PxdpLX
n06j0E8kWyJNyNAYb0G5P8d4PhFXVM6OSbgbPPHFxY1sk/XpZ1oeAOsMmsxAy/4t
uWzO4M1hhW9iFLZNQ32JnDrf4p3hONVhxu+n5yj2APOeYIX+EnesjJy3dl7HT1XF
aa7FLVrCh/DWSrqfwOxkSMBb8FfNQ7hGOnsdJmnV7uQUKoZURNsdyMVo36c2IZpD
w0c24XuEefySaNXGj5eNo9vII9xGHzjF2Ls4fwqepfE1mH6R5EnjRHrCHj5bNnYW
Z+PeNSYbmBE98h/mI7HFLp9kgnWtJ+R1OWCNIYhsWXWwMvl/mvQ5V9SKd3G7y7yl
GyfgGbNphxTGx9Vb9ZeuYAWLtvMhDqpCeaaHhSPhu+XnRljpb8kgxXRrrLLUwhxL
kygRs9rWJGGd8bwDoOcT4foz+gNZrSxd0dk7SiJXjtdl2I7bl6n+ymfoFGOCVIGs
mBRq1QCpqManD7+zSRg8Sbq+rdUrLU3ioo71RCVdz06Dtx4OC4WGkTJsAySDPfcl
vDvwSKtT5tldmEzgFCGwMaYX6y75dweBeGUbYzqjk8VsVFJnCi6a3y08P2fJAKmR
VYeZohbjLjU75VyqnsYyXJzbtMz54KYigRjy+NhSKLQPSYN4l3p0SYXe9g27HAHG
aSJTzqeDrwkUaomExwR7taRjR/381LRLE3GJq/tmT4jha/Mm0HCxiIs/4E0Ami1C
4bL1giC6dYDShkIHeYg7T8nZPOElWRs2SuT+V0/acOOdJvw6cFlDGrd/6EwiMbyU
PeZhnDgxu1APC3hwXQklqGHX0qh46dcR7kq+G7SIjRn1/O5XdVY7PM929/z6nrwu
btaEa5xe3z0pP5/mbLlV8kW70b5zjBVpkBm78oAzarxjuVUPxKt1wZuiowZFUvvr
GQ/OWHrYk8HhLznyZm8mVKzAtHQCvTruiIPIZHyMN3KnkJCSpkAgtvvx24/QKHgP
nngMxuzGxjuCCHCsYqrjdpEBJv0F4/BOo1wF1gaFJ58g1DYhP33TeEPwbaOgWrqL
ZiYPybrDZsPtkwB6Kt2aIvdMgV0/lqbD7IgpSxhDLhPi9BOReYcZT7JUMWDiy4kw
L3hMJV/PGxh8CqzhqUVnXvP+0DBzLr6I9eWANse3BxLoiwviy004a187mIrLrGFO
fiQMJeVexWhuYtZOHU6DQg+u3syu1iNU/BSZFDZZbFLyRhDa2EQqfj3F5L8OW5n3
qDwEzP27urekLHOx2FJ78o4T0eXiBi75zvCfUL4GIkxhKOJqOixDhFjvhGhG/Rbc
vjql9EDDspczWb6yOk5c3hL+HaJiSSOx+/p/kLBRkqyI1UU2jtL4PmpM1QxGqoTf
wOi7tiso/SJTN5X4+NLWWtlkjOHpG0YDNriZMY/m4qbtJe5aAt3ifgprweKIzo6C
BSg5zrzX9vw+JEqbMliSzZNJ23Mlm9dmrejDPXqKYh7i0V3wCa/az+J1fImuZliY
1YjbZmFcvmLVSfQMpYmB7E3OniWE8504ztQ7AX0BCriLnLzZboFHQbNNebBahhsp
lk6f7eD7+lgAD07UxZAgUfrR+S5lBaME9GCxPaSSu52hcCtrXsonYpIYgpDT2bmV
Nb3kJT7S8KgATa3AxTBPkdcqqxSEqt6ZpJPDqQ+loy9shoXfxXfcTkBj1CWpmMYU
qxEFUvgOD3R/wLRSeKA7FdnF+DeYHjijEpOynJpUUf5y90UfWL9Lfhse1BHKd6yH
vFy0/icjp3P2l5DweOz5QaLmrD3Q3YKnPfrCEk1QSZXw/hrZp+JVZiVdBizyUmVD
4vEzyYuWT53hggBFDLcij2ejdtZJM1k+5A2+GgPZ+W0XlJfLhhxSFIWTc+Eo1xI9
Qzy/eXm6Xrj75V7YsDRdBBXrBXd37dgsfNAVFVQXwjNVzFn6NXc3wewhrf73Ppgc
6ArczJj3CB+ZLeQjBhGuR4An3nr94IGPSdVdzE6yLa+6zUTQKodKvvRnHWMJl+hE
byWs4vGqZbE+ZR48h3IwomdLq9h3uApkOpYwUiJuvsMIMIIB6IV5PhU1ABfx0r80
Y0+yR3qSGS7vx9y5hrN1jVQmqg/hZIE123sj+3DA+huoKCO4yi1p+MrGTl/Kb0wY
rrW6y/nS6x6cL2ZpRbdYuX5efkuDDFnScAYmLXc/dE1EgSWJ8fDNAMdYyuUXodij
H2MUJsj2s+dP1WxSCscq5VI9lhVJXk968J1qvUQgrzUtJ9MZMQXC2eyYj21xr6tn
EMBD4Z/WFK9VFn6d2qyxXpG68GHCYzvG0BLHFgtSWH8hwseKi48F3gvzIk892Fr5
NKq6A0/3LB0EeYlNrISzqc/Bvimv1fKZZ9MIqcf7RafRwRvvt61GgccMbpQjLB8z
VtoVL/2/pxeosN8CJOb2mPEPq/QoWDDyln+/OesiXLTwYS9WJt8MdE3npctXFSb5
IPSri3ESp+Ko/jBWwfhA+VAh7exO2CByAP8KVBKuz19zLbiVa8arzjbvV8FvT5ub
uyVRGhoABFpCcA1ol/44iyvCKY8zJCOdVCCJwPs5jyVJRs/mmezpUQL1pAAjZleL
CwekMGq75IX5wSzg54g+C26UcsnEjzCAqsX59mWsZkcqB2KE1fvM7rdXbxNgDQp7
31iR1T4BzNNQvrSszLXCkYoa4RyPoE0YTMh6IYkPvy7Iv1dZWL0lrawnijeZaXhn
cL4UWc1A7oGIVrj5W3D9DLtqSt32Aaj+3MDCdeR+g9I+bp9Ek8+XzTnKaDANRD9k
XlSS9jRaPWdmXGDZJ+CwkFawwRh2DxUw6cGwKMw7s5aZnHtnBSHi8THb3pMq2NoJ
XwOBciYgWDgtQEWUhQHikHLBiMXxRL5UPB6caXGLAYhBTHrWmXrOdnEGLnbDW6Nc
v0PvbYq8XbiESBpHqqiP4edHRfytF10fjT3lIm+tuyerLeAijx3Zx3Qu1UMo/M2/
qsMV1Fa/oPzv7VacKkRiLrWyLIaZVYLPxK9SPRG2MqwiHUfX4CnZCgK3Leu2Sgvs
UPt0i1T/p5HaC3FZMJ2/8CYp+aScgi+5RRggmSQOnVUpr52ZxRSv7O3cemypi+0Z
sSoK0pPHM77j0qDrSrUr/w5CCA/cc8UaZkB794iD7y2DEpUmGHAWNo2vaXxzxDHr
zgIGSpUfQORzUEgy5NgqXSk7Uz12GsCNNQHw90ixAg9zmFBNs8Uyil3axXD1qvBi
O+qQuZPZqvWojEZK/RbJ4MPkhGU0W+lB6PH2OpJROjltY846foQjJO5Le0uPKLsa
mvILZv6Dc+TigzBGINDrBLLaH8DuChQBkPfzkdeFlyhM3iM6sO+Tj4zNH2IOpXQc
VFTPYfwKT9UOSnqhXix+CFDcwAEYkpgX3plZHNDX2oThlIaYY01eWm7mZAzcmDzZ
DL6xvaGubl1yWxPtX3QE8e1jcbuEHd9BunlpMcLHY9H9depcr0m1bSS3SQdfUJ8n
XdPxQkCY8Fxb00sVpsSzWYcAMyFC5tiXOPXGd4knFA8nKQ9YRTDkAAkwxKS5VxWO
lqaUc1aVsn2jGW0cb7tHjO2yG7wPkmExQja3oTezw0ka8lsLg7xw4ZkW0eeHfZOz
oDqEgNNCRnqXiHE5aXrItMHqYM+zqUSJNyEGOqEjfNEuv7GbAdFg7aOTrkppnXbm
ZLhyxrGSGFXxbqJB3X8Xz/zJTbVDQBQdOH+8lAg3vAXiXodwm/KBFQwVs8Tio0Qf
aPoPFt9vvDWi4kv4zHHxMA6/yPwC4TfTO6dQahII/mYZhwSiS2AHbV1xI+aARJV9
OH7Yvq9Cy1y05ZZj/TegIGXcDgRiVngguODM+Bkb9WkQwdz5cf5PK/ZILhami1ah
S+Oth/jFk+rsf9WSF6xr01W5z0/qhNztUzzVWqeO9JsZFIRzEro+Jdxg3kopfb7v
6tZ+UGJVBJn9A2OQ+8kC24/HnPpQnYOWs4IEjeVF+eyKnwsimClD/U2UDtLjMuWC
jlCQDZWcXVoexYdB9MYoVICotS2Z587XGBJlT1Q8N+MZZQ4KkNn/iTS1Ox5eS5w7
miF4AQfd30tdEeknq3STo+a62zdaqfEPHYaz+O8UbckfDTiYUQ0tnmlKj5awBv4u
fftzKMaQA440lKC49zGaLwhUCFgegNyQXL7DF4Q24W1cHxbJOyIw9D7qUUzpFHP6
vpJUOZri5C8IlT1GYceSOvvWjt25g7b21OEzJN6ZrrM876QYxFYysJPFIV0ZY7CR
4cLJ68flEctQzqBieoW445kGWGkgQi7aUY3D1F22yTziimh7lVsdO2UMBY1/LbNG
Yc2f5mV+CbyZMRMnnT9fq+2rbh9sdqO5rO6mW79O7o9TCx41u1kItzPMFIY/QkLa
8Oouvdn9DxSqAG9ei4+QBxV3sf1DnEcUp3mBqx/WYvl0ochXAL4fG12blXm+/2LD
FQgfCd2l0HoQMiYcpeuV8uepF4g+Z1iJLzQRdtYN9UpWzHxXA/jFcByMXrThxkl0
LydQAeKHw/Z8w2Zg4ocS03bU8bYBZa9UmOcjFRxJTvOdD+GMQkN2ean/CmJrtnBi
MbCIk8TBnBA0j2GCmcb6wChccWy/YScH2D1Pb880RP1IZnulD2jYQif1CrYsIwlQ
IoEzluGJIfFWxMbyrIRW8+xYSM/gTle36UhiBPEq+o8vuEbPwoTEexm7C0AFmVki
/AQswj5L1hRFF6e36Nd774VkF2lkECJwwtJwU7M8l9EKuhOqb6hLZBlBDBf1UL0w
1PArSpfdG6GJgyXxFUXNcRdfqE+05uG913GMuG6deil4ADc8CPWPa2CRTw6FYvnC
JwFSoA3igW6GbRGKpeXS1uAf9Cm2abMH2zmt8QMRncoNeq6PtdWagMePKTRXiWO5
i+6CBUC/bx5aWjQRCmJMRxqPCiq3GbAmC59iZ12tU5Nsuwgq3gX9B9wubGXEs8aJ
r+nNkL6r/4h6gFnhU0YBEbBvX1aC5pqsxuZcGNYqMN4lHRXfh4gEtocTulf44xmx
eKauNMBwPlVhg8+3xGfVMULhhsm7cPEXPzYvqNxxjjHX0m6FOHYUT4ealyxcJaxS
229EocBL0Pz0nyCxpWBnhqOdK0dtEynVJF0bEn5ttN5t5EeB/Qu8QpYjHxeBFNC4
i1pq3daQH8XytZ2UPiU5TsciZNt19i2C/GKPLdvkj3LTMl3ZmJZsfda1rszsu7/l
e2aiAqDXatOj7/59W7YdeAw2MPhGDeJHoE+EWfKH6dg2KzuuRrF7oLNcWWB7ire1
+qJrG6RYcZpVUlNOW0xxnnATK7LORp3lRIsb2ybG7CWUGlOPIiJGE1k02LRaxJox
2kYDmltPO/WfJ32U4zObWvL9lalOuPymVd5Xr0pgDz8kBEx4yKuvWDNqu4znEsEx
e+ac4iJCu+ALrGm7CcY6Y3AQS0+A6LQ3uFjVJqNEuc/XwWHv5KJLb9B753FynbCT
jsaat/rMb7RoLfnoz27DDAQqHl4d+Gmo0s4YQfuAvKgQvjK2dmNmI+/ofxbbJhaL
mSNYJGST50URpA4P8RfuEUv1UTK04SW4chTr4aktcBdhRDugRhSE2/GKMqvZad09
ALaWwHpGoFN540GZCGQTyWeiwmrbhQdkpfcNB7yPiymHu5I8daRCst8lxdzBlFPW
w7Y5HClSZ4h/b3/8V9ObbgLUDXIvkdR6oYsFcFPBdEh+P1/f7+DheEdHK+P3JJbu
4WEuffTcKfzwsXSGifUNOqrm+YNB7nDJqdJ990lO/fjLHjzZEZtNHONhvt4FDPqi
F/pr08IOMs5vijHhamF0GtYmTaO3Izc60sNxD6hnnVB9nJJW+4KD80bwEVZkts9B
uzcAqZRWCc06MHMqrF65hKOV+jMteWpCq0aoAyVd9WkKrC89Sj3XI4Q8aS08kmvP
SCl+b3ZmYoqMwzOkNmqmQ3/Xujdkyzt4hPFxQlD7k7yEvxHVJM3uO3jOme3RBx2w
6GJ9llh/7Miv5HJxnUu+UtJ8ISNZEESFEsBMZBVSe3a+oCrZbq+m33TnOGeFwVah
zVL09DW3rwqe4uim/ssZAUIo14K7dxcPyDoKOJ0MwMcGMsm5BGiTxPHvH1uUGSc9
h0nuvp4cfPyTpvzJSBTyPhBFnTWGXYxf330f/45jHDgBTU6IOcAG2qfGWtlYBWFw
mfCGaZ9IduAGB4BX9Z+T5Lc/sjZaKtHePvaWuZcPzKzafjpoPqcNCJFMybGdsUly
LhASkDQkNjC9TTych9mlPTGIm/xjMMWjxlxorWH6uCpooOLC0RxvI7dHWPxMoKNo
yGpkj2KmPNunHUOIHZun+5xbS/f7J5atupf6sXUsxc9pcmmNCzA8eN7OWB2iWqq4
qy3mL6+LnbIjYKsCUjp3kqNRXyKeY01OV8AbCD1+rEh5isx+Zifd8sd5KCpIpTG2
sDur80I+GVIraj3jE0XA1YcN0fJUPCeW7K2n6fR2OUJWJwXoHJf7ykdWNXTAIXPV
Zj/VOA+oeW6HytwphWiOuxgCOQw5WpzG/HRJjJ3spkz1qnZjJ+JM5fz3URD33PVR
FVOGd9nxu3ybsa97Hfdgnzl5z5zdwDcID/Nzr+nqNAwLFuULUdkx0I9Zw68EbSBD
qhi4A3TxhZtAtYHhYxAR19y/pGos7K+322k4KrtQYWw4OvBsxsOo4k4nB0gPALoX
oUr0zi7M531Hl1a+bTnf0pPLy+JXV41q2dSmu1XA7JJ8OcuGyYMNXJ1H5NgpjxO7
oem8HkTkliiJj/YFx6csCJKPfDcS2yPz88DFqjAF8NG/UdCKV6TIg3yIJHBUA+sj
JMIYBp4Lr0CzDh/UjykMqWDuFXeNa1YBFLNofd3+ZwLUsw5lV0NYlSJGp/fimCtp
3yBUEQCM6yZr0YcWdOnru+Zp5TVhz//nbEEzzlVbky+A84rZUueiCfvvmjbtQ6Xd
tBTUpizoOQy9avFIEWok5LQeNT2hXpcE0+Rw7BpoDlVHPAMV3nvosUhts37n1aVY
/jYZvLPs2SQz0AyIshiewChPjgCn3QQBszu8efW/TWBZ9aJR+oj9eg+RNEVxUAVD
MmwrgLJ52ER06847p093Kco+EM0hssVgAQtjtObXX7uCmTHtF1ILZt74Qj/aF1zM
JlTHK8vtJI6x/btLqRSDuYLEDamfqZMl7v7loFgXEgu1PzZfxw61wsPxsQ5bsB23
A1Mpf5dCw9eMI9yAMXScgH1sAF4tzzcG63CFFFtKRNT1Zqqvm/JpU+drXDgjJWM+
J3NFVpO+hfzt0mUHvXuJxrt9pGnrJOW+RF72GXw/lPdHrpd0tbZj8P4B7wPCQbXO
10qt7kNm3Sx7ecjSiG/hN0OlTTXwMUSNZaeaSU2kV/GNI4SVf3SsQ5SMdQtLgkra
8s+Ro5FHFfcSTed1LeA6AVV1NmO1UIXLL8yo2Nc5zid3hdl5WsAgQVtPkebY5AW9
l41AlUORLA1yutwaaIwnD6SE2oNdr9+eXcW1JHDsOJy8NqgiFxjtzbKvq5zVXWuE
fQDuNxGBad/xShijSzrt+p/b3L95yQDh0C0zD0jV3iTPd1qsdAjZspExEMOF1sEO
xFA/WblZyJqp0bfXUwUFyvuwvOVJfDOIfJKDAiTu3KHtui5wRX3QCxYlKzbDWkAB
mCHl/fp5T1UNoftoFqBbBdAN2zfJ4Io8u4W3bh+ERC0yxaye1hZ6du4fUMVZotka
i39GPJgVlLYHiRwmz92MF6U96FnSATx8eGcfccZXBAJAdSjym0L+cntZdDRpgQsN
SPNQDmyxB7w7HKlsqUGA7jSxg7YOzdKy/TtaYhSuSoc+nzwDPpnq6nQD2mLyB/rL
TECHMqOFsMAiEi2lHVUaOG9XqkQrHPxKAeGIM4mq2saAChzDh/Yj9KUhfMFdA3wu
ATtRTlork41EtYfN6qvogFVk7BIy0LVdlyw5Wb2muJnf0hmv2aj5KtfNrNtFXGGC
18Rm3mPAVmZM8Io2o3zTr/C2lvyRstriRCyhc8vQTFVhLNsSm+1q1kvcJ6x9jvQn
LZncbw7vT736VZIZNu5V/dtkQae8TxdNq1SFQZT2Qfsis9A9W1sB8W5EBe9oneAr
xinmkNvaqoprmrpFdLoYFdgIKEIoSVKMgunOwIpqXVDsjJ0jSUKDmmbalWuYQM08
QXz5C6KcDlVZThx0Xb3OGI6q9w0KfU4IJudYACL8UltX3byiXZmF3PqOMR6IKqIA
oPGXnRcRmlaDxdC+Iq+eYaGHEm3SM/lLO4COOtc/BEbkCT/qoBA/dPqwrPnZUv15
Ql+DF3F/RSdmKmxZDPsh6Hzb7xdN7ht5C0QgRrOZvqtuOcuygQPMwsqaNpt4750D
cjim6vBZiC8iLE4S7DowSvRLcvgLt1oQolxoAioebCqm9AeWhtxbbF7WQVHUux47
+DjZlRCMiHTuqgYSHri6FRUST8AeYydebV1AxA3aP0pKkjhpBcz3p/GPLOvvHtnJ
u0EUQyJx8f1aQia1tJn5b2J0UzEQ1nRUJjlbadjjBRD6cR+QZhpBTM4YwxzptKlY
zAajn2q6NC0rFCWJ8SFStWh6q6o1onPr+IxzBzI6l5dBcNFZvSin3LvzixCteQJT
El5yDndD/LKP9eP1ahb85xIoInWQ5Ie3nlrHEgC+g7AYM2ldIqiTLr5Md06YwTps
uCHkr2n3GJyE3qjptzMDZRXGQB+hrORZGtU3fakznsY0BZaG+xu2FSkX/wEYxsU1
etyNSch0KNkbLtYl6b/w6AgeVoxWQo0WYg0EZt5OHuZgR3GCceyrNO7kugEKirGL
fgmYZQ0mvGOb015rl8ic8bNCpn7FRvREUDbia8ixcUSG1mX6D/npQDr4/8Lc+D02
RxQEnWcCwZwxq/k4CS1Z8sJ/6BMeM1+MDq6mbb10MKT8anQfE87mOtcRh2zFYHAf
Ycy0Sa4t5DH4UMa3QxxY8fFMwUqflLwgXMbHdPLUGZxKKZuVSiwOl85F512Mdymj
pm24IL8tVLRfmfJ8+stoEUnjm7XCQoRXK7Q/7ISZx+ZpEnvF8czA19RfGQ5jFwZf
698PYKmDXXu2zO7NfEiowXaDlO01MxvtrFnIwajcXm00Zm41uu6yl+1BZ1JkJQeh
K1f4YTrUkkkxQITJXm4ANa0wud4oc+SPy99B7Sdchgu5QCht4bEIqMXcICI7FWbB
e2nglu3bSSOIpTZzbJbougjm8dLI+TaS/ll2V+DE7VU00pIjdjKc+bh1asrRenV1
2G2Z6s+Sa3xoVPkcu8XzAPSbmD6DlQjjQ4U7vnIMgWP3wib9IAQoz9II5NArACR8
CSFjrzy3Wta2O0MzrvObsIxylGMh+otfn+yZ16Q5sfCT4XUJiezpDAMnsMqBWXAn
sVdPmYLNxnPO3b/JD7CEwczWViX6YqXwDkyqe+ULzvhXZ+EZm+J4WZ+7IpGwo5f7
cS/ZI0MTRbomeQ3YbfPl7Ivdqlpxj1cmbLIi5FYmbVPQFOsNpbOm7dO3v0qeyHT8
30/xHgLcwSUQuXRiLijq4tHsmWoJDqT5eCnFx1e8Hf2BJe2WDOdBbBbg4v+hUomy
jmVHQLVnJ8SrlXvsz8Bphs9T1XvPqs1FMak4vyiIAEZBbvg4yhKqwQg35C+JCLoU
vIEr7pFjVRUxspTL+LXjf3ZRuW08A/xbeON5NDXkO7NaSvnBkLlhk91C4V8tVoeo
ibBQfZeFWmZe0k1Mk2DofCuvzOoHRJkimfSUQYSZk8JZg5P2IWw2qBBNhnAjiext
iGQ97bP6qGSp8S8p7SiXjR/An0ILLLwncpAEUsSWnvBPn2uNn+B+PCwLjA0g01xA
NZ4nGAl74pisCK6FkUFL15o0KkyoivrannesGvVApJ7wZ6lFQUUZfOxJ96ikaEvb
P7AyFlJxV5PK1RcmXWE+O0bhTbG9Fjn5q16xyqWBaf5uVTyMVt/9Q5fdUnmGzae5
iRU2GUFXR2O9n6swI0FYwpr90CzUt4iAbqyGFLXAmRcH5qvlWUzQ65cspAU2iQar
bjLacvgbkFMHA/s3cw+6FlBOZ9zLiFzjU4M987KOw7AQjeo8QDyB5Lp4nI8OmS5e
E4oER3ngjBZnNyWm5BBjakRuRN+Pl9VOe3H9sG7RNrQZ06W6jkZX3IuEY4ZFnLMP
++j9f9DhbR2u1682hMi5NTGWSIPVRSitKy1x7QSwzQSEiRtMVdpWyXXIjCF17kac
fkd66amSaKdUJ8JzYZDKzL/8TWit0/toX2V2cXUjPt9IJU+Ewol9psZxziR7H80g
LHc0IrjQdyadDsiGHvvwYxAdsEVOHzSnO55DBZHoSqDkYLgtKoyCzpw/g0E3xti0
Q9QOfdeT864nUrAljmhw68XU7IUebJAo1WMq9iIWP5TXhEgY84BJAPT1Wc5sj/jr
0dO6J0c7FpIaWgu/7xA0fbJyAKG71czrn26/4jvyS7UJB80Gfszxp5LyBIXL2CuD
HKyF2vQ6A0LdozLruiKFscF7ZLdK2GlScJ/3QdCwkaWqzHEm2LPfvrEOGXTAb4mf
0Y50HbF4+Jo4aiDXI+73jdqVnZZd+HQ8VPL+DdT2xgJ/Lr51ZTwGRiIU44DZg9VO
iBh+Gr5QQLc6PNISKtWL278UM5Io4ygmPfuDmlZoHpXpWhuEhvFycopDtWuST+mT
7ptqJIclVK2Gw18NodA98vjnekpfMjaHHxeaxmbSRj/GrwQqZ1n1EiMTdD+q0H47
gSxQ2FrVjQl0v1GDks5ci3TcuJAicGcz/8JXwDvZNmZ9pp9Q0YLD4yTjTb/HM0t5
cYb9F7HxX3S+51qiu5sYPuxlvp6COFipRWY3npjSmRGpZpo2uuDiO7027ef24XFn
N3B7hNEO/2PUyk57S8rJ+G7Ek3PmB16DLMDmErABy1+n7J0TqWFRvJf9TVqUaqOw
d0jbtapOGNr9D10rwNV8XrW/jLlZAAe0WqQGufk67LTpxAvaafNAuOwRgnktrI13
De1+wlrsZUVyFWCjJVVCKXYJyR5XO2Qlj3yYtm95WNkMYQrEOVFtB43r9wDkNDg7
OA/qX7gwyl3NYtsd177R1boNZE/Rwo/eOc7XY0RUeS0EwWwcmPsQ3RXb3rC1eNi+
a0dAIdD8+ZWLMAW0neK/aVsUUXlFTU0qP2eBMI/MHjLgTSCXkyaiI8UvSNnHxi4M
7k7uocLbyjcTniOE2xd5Np0nhIh5vhTxEk5MT8Y2c5pr2ZQO0QZ1UhgFng4OMdTv
F3cwKe8EzW4iF3Ntpe6+01JIbZg+qvCjDwkjBdn2xLfXykJ4lnekyhVqhniDPTgu
dDOhHgUnWb3sEn7nLQkApqoAT+yrTobwOqsdNxtQmqTuMOdMpCIcpHNSMjmDnydg
fHztaejY3V4tyv53Ql/E1/nQWtm0OuUEvhPh87p8bQ86LGIZzFw7P+bbJF7T8zhn
PKvPraqfuoMq/cx1Kp4WT7Rl8cbw5o9H0+OvvrmWMcRpaIvzh096K31FUNU8c1VM
gWxSzeqLKMxv1bE+aos59CmVOQ+m2UwW1eWrtR0we+oLbO5VHcxZlzs7nt3dj3o9
yqj8wrBZKeev5U37jVGMB/g660VtW+Z6g+N6l/FzawC9Ow0cBIBq+dsz3Tottm8n
uazGs5H4BkzHKrkbXIFHM67ccLvw4QvGhxfVGniYBmq6hGVygAKgXtPr8jCe5VFv
UcyZoAG3EO921kkzVFXMw6J/FV25DeKylsVfa1v1SM+Wz512qaO9L2Tg6HSEk2Ho
Yak8xidYYUGAtJo76oOddsg3oLKGBB9ONuOAB/SfsHwH9Y+2QXbyR2AF06Y7iv0j
L8Pw9Apn53gtKrPwuaoMnp+fW72JsUxgBA2KEoMfZNwt6jwHCuk2dNl2hASFwfrE
I4LBFtANBfNsVvqmEnkRsFHX+bd2DJf/5FHdVNi6+vBT5OOCNo1/V58N8pFEIPEQ
NxLdjaE8p56THq0rPyYSFqfhLvaKiJn7UwwAGzPjSDgrmvgPN/PC/+w2Qfg3+gWR
xGp/3PY2Koreh3syG828AgPllAbPGMu0cm/z20fD71KZazWMvfmlfhKao7V0neF5
gP/tE42qbovLWXM2vql8u56UWpMY8YIKuygmAeXBOY0cihMlFwHZKjP5zHarHyiE
cBwR7T9wr5KnOr3ZnZD9/aEmJDljELmFD8uTNNSvXVWdYSWWKG/t4RoM8KlMLR76
KkD28+EdJ+TGMkSYu6qTjNifqY4DMvBbFVNFzkCjQsk1OVDbIe98/VWXmNWXhJoG
BB49lbMdm4HjeUSk/+EOF2gpQN4j/NWLQI3XpPtT1zbJPYlvgJLSfzw9C66hnObY
nJqzxV0Y9yA+Ozgu53leLA7fjFhBN0XKkE3qGu0EYGJWAusNA7N8YzIzESe4pGL1
IOTY/cWdduEErGyy22vxE9c6LU5V9ECgH8VWI6ClCUAYjGuHrK72tulme9rbfP6C
emdRQJSVfY2tx0j8uJgf34Ay3CQr3OrJQE95b4dZq0bZfpem9uQ2e5tfL6mwjQOt
cENN9y/SUZAcCkNM58ILcaSUoa+r6aPQvlu1CUb0g3Z3f4I+9SHjqhflyoSYHabj
ESSCxZ3aJonGGBvkXRn4XdPiRYCO3Y1BagaNTyowrdrIQeOp8GMfMpPVwmV5m6Vy
7wN3/xUzhw5A5HIibt5kFg0HmJAK1Yu/HkEgKMEYrJNtyD/ePLjgVmdEQ65MlQgU
i/K4KByACyTQ6PqV2KL/tVjewGpoXACQzrsxmG0cr1RlcoQwLMlADKlnRX1NpQQX
zQs+Dgv2IHGvnuALlxzEPaFQF2f505WwATIXeY60N1x7JZGANi9C94ukLZDqBIYx
hkfp3SDMHVz9ibVJtUazws9YETv2+cdGm7S1F59S+UAndkin/n4hUpFPKay04RQt
HYZH8dkjyePzC0iUQUGcqy7qE+9P0xDvjYizCE5dHOvf4iDJJAzBKXbkPGBreL8G
W2Uk+wMRyRJ0y6ZsAF+AnA7vSzmou9P+BtPDEEWrYvJIvQRDPpK6TtsQBIBwm65j
Sk7b5FumAebN2xM6oCQRpWL5UDAuutYZO7/Gso+hKIOmXtgts5k+ujU8w0Ik1chl
wDNrRhfcOAfPZvRka6nVZhkHK9+5ZJZOn98DvvTwRtiSK3LX6ULPNiIdLhUzZXFl
lq3IOcBwqsLPkpz1EqRgpLSHw2mimNwA+v0uyhaJAVnDbhsn+AJUqW9kVbG4KSFi
t6hf53KkMARfwbls9hx4i52kzNgq3A0XIIA9M3IXnIJjphIiGa5thP9jyxUhPyJ2
OibKSXu17Z8O3cX20uavmpzWSCW/FY9P3edqK/W6XomIRBBc/DIRNH4Qay2IRP4a
cbYHqOiDKFvzVauZAHSLDqmvlwBnC7wR6zqWVLGo8MLvtPQDGKneNU67D9erEK0p
NvAvL9oMYRwY45Z7HBBSkBrxX1+w4/VOCmRetu7mpnhNSlVP/uzyyJ9DxsGWovfE
MNMIv+wpd6ZMqLTGYcP5VI70ewny+DIFjb+rQuknD8l+WbevSksaLvtsNObp7B5f
I2MYFuRhB0RdbjeFlyLO9ewOB+RB70V702BVOxQWISWTWrk2vnb3EZi6uhD3c5El
TinnHqwySKB6wrKJ1KIC44+BxjrrsIZc+SdReuuLnmq8DCVVHXQqXMd9Gh4XRkVk
1kDb5lih1oPAOmKQ+ILWStCMaQ7xlvSwAu0jLDDuM2w0km1yvNxMMHnlUxJlxOwC
pP0fiuhv8okkNeUly6IvxPWcGeipIEwnqECbPDCYXEiKGHcqC6pbL2LMFnY3wArY
jZrVmbJ82YooukAjWdXNMquUcbHi9rEFtgRl/NgNO1AEdsaFLDA80k+5CZuYh0mk
yURI7AjamCV46spAVNLIvXs6xfKsdIXmOG/SZtVbWnmixXwAV+BnrBXb+sZ2wl/u
yhY09KbghoFnmpoTb6Dhrv3nqRzkUKf/9cmqDV/sRzcEU5izd+YS+xfCdQupowpd
mWZPk0rBnfFVPmOW/AfDIjmPJmZVdxU0otcmmSy9lgmTF+U/PDFV5SL+fwPacDxV
W38BD4uEihY3nkmDdmM0+e+1WmE9n524ci+IZAo3UbkohsXybIm9v+0mxeIa8k/b
5+Y80D98H8Fn3TT/Yh8AXb9LOiHRkLmRoXQW2dgiUyrRyG++SK4yRntBO4bHNJGi
6VzeFsU1SEBFXLns5PAybQy7lv4E+e9Jz0XPcheGrBs4407fYTJhRIZ3aPyskdBb
YgJtX83zEIZPmj5oEVVVjgqvnUgfT1zaKFlyprfDYuCZoZla5IrcxWzkWpWEXSWl
fqiNCoFuKWIMu6hZ9LE7cEgOquEKecQi5TXFu/3+6NsByYKX5whmc7joPlw8lplG
E3GDgTe1LtVAocODYIfMP4nTmcgoUYSKyORXcCy3shg3txyOfXDuuireoq1RG+zZ
krRSdD5roI/1kj/6aCEBOvM+Fu8VxKvoa1F5+O48PvQC8f602/ZMOfT0KZb9MfUN
G45iNazK2OnBHxfQX7apcyFDiGj2eHcmp7TE0zi92ZE4IPWC36pzk8n57sZ9FaPo
mpYkxA+jeFN1QrGpz43C2ywx6GHdmiIJU3VAzrnqbP3VX4F6HmPIshfKzUe8EO3T
PV6t1p1Pg8hEo99dSmaVuSQWt7fNPS5GZH+45LqPf9nV1nOc/SKUSVDdnyWfEa0V
s3/9dS2FpCqdnKw+ZB4qnH7dWOzospERFHrJuCHHJZu5wckZvpMGUh1WIhfrLkCC
hzu0BnLagNIATYGSJSm9XuMWeQZI9N1OBU0hDAxU0+aHkyD5aD0mWKhTyTrhnHah
diviel3uWfp/tDJB7pEwZRoKStsIhTkA1HLBWINJ0Jsy9JLPEO6ZwVSubzfi6+LD
OXvBz59Lgucf7HZBh/His9xX8XVPGnsSlaUOdPAEt4fUwZlQOp4ncJFp7UrleIr0
sCW8gRfrapER1BApAGZG1jq/LACLxvdUgXd6/x2F65QFNTPkeL07GCjJeFREbaAL
7DJlZmFI5e8Fs9YfQNE13s3Fba8+ewP4DgJiT3OUvC/fZjAkSlQnuJuCe5T8E5aY
CVYI/p9dvLDslQ07NGGkf7xSZwEETv5uoMOBETjtTFidYU+9HKcqeUbbSs38SeZz
oDY4RnIRka5RulJ7Y289mM6VgNIfpkCTWCD5IZKSxYv0w2hhX8tv+Lub+tbOw5aT
Q0/RZYjP4EgBXIVLhN5izUzK0SuQCXWe0DEUOT5rFGG2zYZRlaCKzIEaDLQNdPRU
GJ8yKwdINRhjOaGDbcLHyH4X7up6nfSbQV44Qiz39AN80c8icwzzb8xsjwsb9w/t
FO6OslK3EiDmOI8r454uo9qt/EliZkAVgZc9q3tXIPQcafQlfOEPIEtG8y2Mbt7c
jZnxfTLV5JbXytwHOTEFa+PSZKL/18T8UPmfl4EmOmad/OSVKYESa7jPbFsLBrEL
otGvyBxcHE3i4VWyuN4Wbb4BiChzWw81PIGPLHB9/nn0OFAVV/oy/jn9T6afyavd
cnDeDaSMdZqhRGO3PodV6IM6ga/oigu4Zh4jin0XoJbjkdBw6apKhDdMKiPykjVq
VEyE6dXM4ZxSyq7HZ8fo15DAlCx5HTVjZkaJEC3vVpk7vDyW24Oq/668oDMZD26j
9GLkGbmE7P4VwSDpPSL1SNZZtjJeluBNeIJt3BWLk7BU/SYKbcTVHKhMAbvM8Oh6
ASbAepNWVGzBuRK1UAhDW9iobr1DFhduWrkP888PCgSh1/fVrRoN1OM0GKugxaqS
CFb5r2MwVbSmfCrxtJojqoAbdfeWSErkI09RwUib6dEk9y1nT1P6yl+OTKCmh4ss
QrTMPf0SKpbGiHlP2v+tGXwH/jboGuuJ0vlSXITChUuk8ZEq4zRlYc0kHCCpiVe2
AavvGqOkCtGEdhBTldOnmQWK+zVa+u+xwqjXQxw3zBCRYdemxnNZsLfwYfDC/Q4V
TTA0CDrFomF6VQJ2ct8RT3Ha4msSARnvqXF2TSnZZtDOpMFSUYNOW3dyN3Cj/h6n
1xOSGSF0G3uTyyxFwvFdXjxeTJwcqzRJHErMiYnSwGcd/PamBYOzDTP7BM8mjy6R
a8tDJCggDgoUzQ9MSzhmQNL4312sYWj//CpLQXs83f58AB9z7lZRtcXkd7DbVEWu
LTbfvV8ppkrmrTbpUxeXpC7jaClqlMqjpaHc9wgCzulqeEMCdjcpTcGm3zRh6zUW
NKkfmovzwuO876vI28rh8KMn34wWWM/REZJY0paEx46aVMwItS+y5RXHYR1b3LJt
nKMxACC13TWeDIWJ9gijXeQaSKPNP+Sx/Q0ZtyT59kV6os4cyr3kdjB3tszLn+Xi
/EiPySnk/ZZ1pXt3cxYbcFRl6acwfNotPAqO0FcS2wnTJkFYWigICvzsGVd/2VaN
JTlhkq2uqJxONdo3JMREg1WneCZp8mG4cyOftG5rTw/EQIWeh7MRrjJGT+9i9Wbc
umvgykMRG5tFjBdqkyFPo7BIXmarmsYj6f732T3HSvrnf8jd/S5xot5V+VNXpxmQ
lwXI44BD59NSZu4cWE0BnT2nLBQiaKBI6TPDKcuPUabLgWJyfEg5p1g+AykHe/3Z
AvGMtxbiMPrMRIEucYIR3T2MOO3731Cd1HFKeU+xHZJckCn2IoaGPUI0nT2Run93
JERoXA+UnoxpkQV0LVv9jkvx9X/qPWpCifYnTXC4XLO0Ok4PzCPKGQZnPcXw6s0/
pYw6Xpc7UMM5o9pXvuyNbdIsrreeawlpPveZ5UdOdazFN0Sg450r0DgEoj+8gB0G
XnD74gwp8mwr74SAzef0e8uRikkoAkR2iB0e542xEh6cjy0VfcH6jiz6Tz0Pcj8W
zh7aSMsHWRDuEyeTH6Q4DhORO1GGiv/Fbwy9bZuulfxjwoPYH35tg9Y+8yA3mwyM
DYQNf8Y4sKKXXOzsKpm68VUXLP25qmnrSzWqtSH1HaoLgAzW0gK5ApIOzcKlfAU1
TE31vWNZ1PC6MVXyFo3tS+yxDROasfz0lzIOxnLeq3mXZkXwwm13Ubrlzif4YYT1
1rIqF/RSb3kchE0mFbZpvR9BWp1S2vznloB6c38FlUL1nogjQkkpE7xc8OnUESFy
WisCd8hVFIfV993FOqa90zQm4JJLbBegcTQXrrU4IQjsWcZu9uFRvbseOubndSJQ
W1MvacIrM0+bUP4TIfCUVb30KOmzn4c1WRfvTg92igFlxW500BQxgpXdED+28vWo
f/iOKnXY+ER8anwWUteRV3lh+7ux+4AM25Xvb0aqtXXFrIZKYsmKIPZ1cilRpVgc
uRQXoen34X1ylZ62vkMnds0wqYzDWWaDnEvHbRR0W97mV2yayANNToNq1OuhYKxi
XaNpRsKdhcW/niAeoBQI3WS77OHdayJ0MlzIZizF/BHZKq9QznGxfT8c1pC3HRwF
hnnuTiTVIentroqwfvC70thxSPJgUVefbPtrLx171FE7wnFysHyJVtCkEI+NeXQ3
blXupnjnP4QgrlIm5qNLXjKdWXD79mCv+pJTxaGN81bCVUpEjwdoDUEekIV1lCLp
irHLMPxP9UjgzgMEWYJobqbyDwFzoJRB5AW/feAw1siZTctQ83Sp15xNEOWZzvmE
t0Ttapi8C7Gu6BXwLYVT7GjBKP0SKz0G5yI+H50YfJ4FJPeO3LaxljQmPYUu5tIF
j5vYceYUtIUz3z1Yf9FU1lXdCvUCYsNolyqBtBaRinzZ7UZ+pFUPyEnYAfeELptM
6yY8Nl8ZGfQDAYthL6vOb+6eBo2ZhiS6gU2wnogQo2GEHpWJjLhM4RShnfns6VD6
4f+086CA0R2+wYByWnlimn4L697daW0YC4xqUG8kyfbKJSGp/25RAX8rDX002k9I
038etnH7ShLVzvdnV9cFoIM6TmTZwrzYeN/DO0sNRjH9qM/0pSCkXlVdbbG8o3Sp
QZ1sx2JCgdpTrIaC/hVIHB5aGWmL7zmUdifhgy6XTWEWisF8ZoR0SHk4E0ZHFxdP
nh/VsR9TMriAQ4Pezw21AK79boWUX5xqpptKiyx/t/CqmBqkhTAi/hDvrBzUL1P7
ObnyfEy0Kn7Ry3tNaofLSRPv1lAUdD7Fxu7LSc0L6H3CbpQiQkddbN6zx9zCmuJr
VIeM7Yh82miHN1VneNKrxel+81k9GC5HaJMS4snF8PCak9h8RxLcS75LkkXVqZkE
NFMJ/WqgmdhnKmhbmBjDFw+LjL8B9JzRWevsp2IJ2/LbZ8qL8AhDigp5Wes0Hmwl
awO5MixzYaZtFMnhD5LvRupS+TzmbHc6s47w7lVimAd8miJME5vUsL7xtou9efnh
Ym2bG+yqloWyD2FkVdW+5KGMHZ3y6GvQtdwIGmvvz8ljIX8pToG/YjalvkEEIi+P
teJf68AVzpKelY8R3KI/4cAFj8KwViI8B7FTHfESlFreNTaJZ/DsRnaoCpvrdhGf
qVAxGBrUBeUwiSMNBBo/3eTt2a6a/7Kw35xaojIZClNsBUCZMOp/2x5uWGHsEI3D
0E1YCil39u9RWag3QGSchYpG/PtSRu8DRa9/KFOzrG4X620+RaAZcY12mCg6sizu
vG2M6TbQUonCbq3bjHhnQmubU+68xEIVnIw16YyclDCKihqD5qqVwGbxhu7Fvqx3
dIRDaZNY/ylWRa0wcz1Db2HCbA+Ikc/57JR3def6Lh00/guvKAeeI0FN0ADC8nsG
X4lwCoEJNMLg7RcULQn8pvs2nQlE4HMuZfsj+LRjaE18Ha8KAi8EnDbSBJ/ZxTaG
VgHEoh3E8j75zToI2s1ohSidGZ1Xgin+r4QD4WmBNfOpKok1OprMhJGs00gZI1lY
qj+bXKeP0e88xYOa5Rw7oK43OBbDRtFCiBtjdzZqdE7br16TuIwuNLsMF+kBqVNn
Mi3omrXwp5K8q09k64DXkjEBAKKELjU9ubXGIXvn2hBV9pxC4fCCGtQXA7KjKwKu
sm8rxTaMu2XEX2anrU4K2fzHPBbakT6NAHlGB+AygVh1Nfx8P3yLhJ4vHzyeZztE
OeciXIuGe+BMpBeL852QPhN3Bef3nfgizGZuK+ENO9Ue5o51LflzfAehb5rWWVA/
3lgdrI495b7K3YaYZOgZF/31fGM9FFf46y03wwv2MeDAqEojf5Dm3ul5RE9K2wtN
/ZoudWcf2+8/opxTgQQNkchGAo/jpRzWo+kI8TfcYRYyf8HNW0txno5NPJvnq3rx
3ifUXkYu/2eatE9M9Q1Lvo+xwnQnRqbtE40q/c0/yrQaJWJENADUrRoIlqiCtgPL
hTO34qkIKo3wvhxU4K/V62Rj3NE8p4abWzULe4aALI7WrLyGbRxlLuKY/IqAK2qg
GB/9vpjfjmYdYUqUz5LtzSWQALZIHfC46z24glFxA7pT+ic/Q+5ba+KSi59iHs5/
7LTxX3qm0NKbqi8fBDfvC/Y9fU7dsDkmQ2VXeElEjsOiVWC88LwTwVyDFMri29ht
p7pcN29aBNbyFdACQVDRDfTlqKsxwSVXJFQRuyDwLTMUJiOlIm1nKoFjODRcdLV2
kRBqvlMX11XQcOgwlnqyWE1Zr/8u/OsTN+NPOhv2IyGVu9HN/qgUSlUSzN6QA5q3
A4ENjenXlxYGbVwe80cXwvtv0LHFtkOco+UNdYcUA8WhzhaCjtD75vXMxj3h5xbA
WPK6d02v6G/ZBBpCoALxanOarCFVo1b+BTgfYJT+jlgXPXE0QeS8wtzOxyYTyNET
nn/b4dSU4GLcvbzXpRbEIOfoKLa+BWRpODrPZIowkpqX2r1KJoQNKUeqlCphu/Si
fKPNanEg+uNcri3cKlCEEuYnxfejEgkw/SHUv9u1PSIupC2FeCIF8mPEaVR/U2qf
y85SpmJYKV6jcgk8FAAFqxuJAvkPewEgvL6lkpamk5+deOb1ODi6W7Q0q50NgkpZ
JOcPi23d9GrNq1/VFVpJLgbRgHdUH7leo98hbQs8Yb6MZrxeYefVb7DCCZBRk9mi
UFZJhmkfQgbizdpF1qUHsPAR69xrFNWpijSIKVgVKcejWy/GnLbrtloiodtbENzK
0bemrKCSznWUAbkE5ZyJ/F/su0H0oIb+dhGcbHVYBC0Ldq9+RbHSNNenkh0CKM1g
aCVxf1N3eElEmcomiz3Db8mxFQlwB5cgnLMy1/zswtFdpIDQgjve7Kx5Yqi4IkjA
d0YPNbpL+Uh/hCEgktX09nzdmrvuJfpSS1bbpAhgIRZZzLt9hAoGQ7sOIE2LHQBK
VQFKUGwEiVyATCbM8gpTX/GFso/CTDWGKhyK6tD0LyOTFRy504ix5rF799tZqyCN
b7g677qNe0P01t5MG6gQmjtYO2Cw4tOLFOXg0nk6gnU5SlphLqBeV2mxaQb1b7RO
NnDSyR9pnaoIr0y77LpJEhk11lmtJgTeqLxpG908H4eRavKMmHcWN+vpty3FgXT7
ZOK/yjD4GLFpn9IUzTk0c/Fu8DQUyQZbOY/AwkoOsqFPymbNiB0aHPcnKn7kB3h5
s16BidwlAFrP57k/AsUOnH8rrMV9AYbRDlVluiG5ISwjP9InVgqzFXUCTpYXuhSV
zlvPM1zMu8EVB3DB9Axwg4fy8GFMY2jLqD6AvrODtJkknpDNqOLcxwNTv1WgUAFl
AnB9ypu2mU++54TnTakyFSfJswo7AxW2ik50aSvjwlWbg4GrrU/egiEj/RHEHT9U
QnlTIvc5u+Ga1rSxps10Oe6ShWMRz4Iv8HYqVn3N237v0xx6/AuC0do0N9GVXKhN
CnsEOcXmQmTpYdnTJafGS5zrB32t5eRwSO2GhUzcFeHLIwp+ZokSbBYq0aRa5F1P
om9+thz0TfpeZzrQ7tqWvQ99PaHcYCGoWe3jUgwrftpygYoZl53a8rlQJrhastD8
SK953up2TOZp+yYa4HOWxMZ2VBguQ0JY1pnFl1kr5Wakm9PvmGTSW0SvO56D8dIJ
tB42sAVg6M+wuozPWTrArcjSkgiErQ5KhiQ7g72/BbDwHg0/jMJtFXCqDmjCwYpE
JZai1GUni0WAiVbF6G8xRzYM7PKjxc/KgC3/ov8WuUWEiJiAlmJ+Uy06pyf1AJJg
otZz9MWTKNKJZatpcsk1Y74sC1YJ7YwZxLcHs7KRKjavtRLfXnYcoXoUE/zaQxfi
PMaqYUUuys4bxmsv03iYpslnv90zMkTrazk/qE7DbwaCrqYaVpZO73Il7opmF/1x
BSB1zCC1vWKQvKuLnnytvuVRgspW/N8Yr0CR/Hgf5zvcAH+M6XluPB+a09Y0M5zf
fLdTGrJNURdchiI1IdS623FLxJrh7RWEdaUAVUc8sK/awQYWpLPpSGZvy+Ooexen
ecdgKCWCs+ltUBb8giXXhmtLPfc8UMmImh4nDcpxwU/W+0z7iED9VonTlSKD+69J
mMcBMPDyHth0TbVbckotYGZngZSCmOS22g5QiBYO+S5f1R6GsZuRbb6QxrfSmFX/
M2cwIa+O6CWqZPnlY8j5DmToKPGFBk04izPsX/DjeePuktS5hrcIZKY6Sf1EKzbU
OD2FBSNXHCaKTZyC/E7l6C7v5xfH+29HUAhelvtYLkMOlxpr9n/M/c8AQ8iGWluD
i+ELZzH1RYJvX0sNCoy/emJL8PofwEJAql+HLNca9pg+EyXAvJY36IfBMOoQ+BeV
OQ6Q/om5FYVGs4PJMRmE8pkfTm5MWkogEtjkPbKDkQaWLQ3WYM/1Joiz08AXwZ+t
umMvIJmmgeDHmOa3Sl6nXUxOqXVpmFUMnMdkQg8sURqsrWuy/XJNRbucDvcDNSjZ
UjQzEBVUTe1bZeIoiNGk5RkjxdKSlwJTljuYebiPmuYmVCpTkXE7dL9kX1jWdHIw
aJD/qh8ol3esNXiESC9SlEaCizHvTG5rCe3+Pw1G20pa19GBQBIaq3EVb8cfi5eZ
y2D9OgsKEElyZTyhcl8ZGqDIQOunWFadqltSk3p+ChpF1LWOuymH2OW9ICEqHRc7
NGCPAe/3b8TEyAZWjjaZ5uGPPGTSENMQAY7tvVoc0SxtT7dkeywnSFT4uwaYl/xb
L2e5S9LeTCLpVauyGEYoFOTcl7E7BQcqVJAvwnrgCnHzKC8JfupuLLydF2ujycXF
DHPvozpeZzmNjm7yLluRHLDxd7zYqXPXUmyNd2EHcqTGKwMX3SgSJcxT16HJS4A2
cGc7W7LGmrhSi3IuaIChJlZeddM7tiLnm6aImqB8GNqqs1eCPwz1EscX4BV/TKzx
xsFOdPB4ZnM8+X1Q0OK7j3Q5EYtJw586ETPEc/TvJ/YhyZ+2yHCfKWOQ/xi/1/Lt
m08NXUCs5AMz9+va9fwTr5JpQz9YOgRb9LsDgfm5gYrkU7/E7ER3Y3R2G636PW/M
lPYykdRi1jlSug9+oKLAaVs1ymeIm468qePYoVw4cE94NblXWCgIJgeeOLerLwcx
vh4YDNT1jN+ML3sQb7gsJzfqvqJlcWR5maTBccv8aEbXCWkvxoerA748Zz8uXgRB
7h7asRdSW3Gemk/9nhZTo4/KMx2CPPecdF4mX7BLCmF4qbZMskwCKqWIxhWlUfZv
juqToDJoDojSxJf+oUv2uHlPLJb75EDBVeSiC0iZyqBGoZSjcfcRcHZW4fnwnjBc
Z876wuYJW/Cui0lWNGHv++wwWePqEYryGsd0Gktu0aJ/fxQM9h6criJTHwfjX5h6
YdmHIdJW+6n4i9kykoxt5V3HW2sLkCcM84N+/g9xE5bCz93omAcI/g7M22EeAlOY
c+5Amf/sKQC7KVWS7gILd/uItrSByrFwyL+gSbPo+uxIFya3fOKU7+0kQ9fRy9GW
vUIJ69L3psxXDN5oBto7O2PhTATeSaCyuDtMmZn4jrXgZgYNTPzHK+Rr5u3Iud6X
vVazLWDvHnF2V51sBVobBNZo9ARThll9zkqfafM4bvrKjvmu7xsqgOoAqQoM1OOo
Qpa4lNwmq1fJl3oKRrxq0es/0RA6xdkMcOC2c9iABrkHqmqJ7mDErE3Ooa/aqopv
EnH+vYcReE4O0HovBtwvj/Z0t37+N1oeNucjWxwPsj3nTpGyKIKBa0wmsDLPQpte
GzrsYLH6DqPEQQ80khe93xNqdvwxGhrqYYD0hdP7tOGT6RVmZJqL+vOlotJ0V72z
NOZsX5ieJaESXEPCn2cpYZdDUAZlB/9xXEKq9nQwWRuSBWzQoEra1Td9mOoMwA0I
pKX2AwffCoPy2X2HQpDnRdEUYNcgu/G9wDxeE/lk7F2C2RMRTz8N/DzGGs8/yrlO
Radxskv27HrpyOt+6FAOZyBDA6JjCC4kcr8COvtkUlSXTaFGFaw9u5KIcWtP+T3U
y66Kay/m787ugHbsKqUyMM+/sUEm6lcASKZltGDX0CJuOmgKJ19s5eEMCHTMhJE/
jQDVz9SuhLLQ8DdjcequV5m0rtr0uRG8H3bzjuDQaguMCl4nGlRj358NCwn5Ey5u
rE7PiuozQQx74YkLiTqoFPjDl/3LC87DARvicfjt7eV5KUgctnemqpGUsmy9KK/x
fhn+/63+noddrb4bz+xVetmyiGgM2QfNgGiEtCaN5ICtSf1u8j672h64jsBsU+VN
fDNo74S/jyjs2OdvTFwyWSCUywlPSj+/Ml0KV2vV3o9aWhPGYXbgsBS6hrl0YJtA
FoniZg3xIyFo/u7xdV1WjPG7anDBqwtH/9CBNLHNVsCzJDmv9SJQkMSn7d5RX1gK
OP4cBjK0UJ7IJXUn89i48fpWDLAlZpn3GfNUaUnT68EW326Pfo0SPppQIGvMyYRe
Q+1/f3rIFw4Nf6EBosklHa9hYLaO6Gi+F4T+p2R+nzxeS4tJKv7iJ5hogvs7Xra6
ikZedAa7nzrAdt3a0ftOhMU5NTA5xTHH/yiXTNMzMQ+AM+dP+99bIOAGqPuGvaRF
Qd+oQ+W0jcZthhKMhbtWE9jqOHX0wWG83iZzlzT1nWKpnJJd9GQAOqJ96F2Mne5n
oaJPvZvk45sKUL51cqAiIeXaL5CbzZAf6L0ekWDs/zJoYvQivroOxLaIKiSUEV2q
lwBBSl/mUeVivaKFiuwJ1YDZ9WOdSsHNYUgUBjndSpAmCYWuGGFZM2gQBH8GEYoi
7Hil2uzq+W/FKGgUAD2Z44mup4A1zXNMEjZB6w5a/0fJKTVHt/A0DxiVZDE4xvU3
BG7F9anx6qu9WfDCBQ/3tUpCd3i2bkcOEt7eHaStqTVrBZKSUDzE9yQoSIJEUvE9
LMpitVusm//zeLfVPRXoiFCYE1XD1qPxZ9N+qTJPtTBNcsoH0CzZvEEAI36b9BfN
VnpwaQ6bQmVxD0ktQDVUu49ahDnaRWT6QJiR4Hht1rkBENGBUJw1UGQnfTNDe2L/
1re2YmAzRcwQQDou3GNe7O25xJgZUezl4mRgHNBNMUFq0PXfRuTM5U05Syij+Qgu
BoF949VV/3mswNgz0LQiLlof5w0utKIieYEAkJtOfTjJzv04Yp7/mrb4A+UrImEm
mL3EvA6fsFTfxkb0fKc4PCqxdgvIIKSMTa2oBsApy5MLLmGZcPQQR7DdsrCC3yOV
jC9lulH3j4zT7a13h5qdTnyqUJmUJBGhbHytRRwQLpI0DOyYDXF7c5OT4l/dPu14
ODKOxnGAvdUJqroYnnW1YsiyB7XFPqdfpMi84QAbJQIKsS+dYMxt2YaiZTnj7vXr
ZTdeT6BECn93ghj2CR0wBBxW0aPLnwWY6Gb7WN3ukJaYyYAj627k+iTtxnaxwSuf
sZWXZ01NVMvvSC4cGNESy42sexjbx8pzqOAmh6E5u3D9J0p8usgTM4RqjRFdo1U1
HG5rjaR8x1mVD3F3iVXq+ZQ6ZuN4Bgq0EAlTlmQcKBkf56DnAWwPnniUIrUPHTCE
TVLpNkrYZKymkWEH0d8LSKP7nbN8j+FHoGtrB2sGjgIJNy2gNgTkydPSvDTmS0iB
BmX1h4gbaz1Fe15ArIRSVxRH406K+P7TZUnVm/R2itZNr25g7V2ibZTu8CE0uy23
B/xag2V1o97NLQ4oAixK2rMe7WOMQFc7qps2g5zGCcgcXCRTNbdTbhK70HcdkA8M
f7mOl+tcu32V4pLMblu8JGV4iSAFI4B4P9bkrA66TMO5C97rwZj++2a2L+3vt4cJ
UlNOp2r4gHF+CIjQ2DkRMTHG0fy7qie8uJe+q3iD27GXsFeI+utsGlSxzuspNCXk
JrmNHOMhYO9vnlaH7oXgeOs3/vEJhS499xgMgYBCXZ5VGzv1FxmvPnXGR1rzTLN7
aFRhb1O13MTK3+Vf62xq3w/C0QItKnmTwN7MY3MC/jqqGrV+Kw9V111nn8IPMMVZ
Jz2j2lcBJvfbaH0Ps4sf8EBDYNLgnNPiW4nbG75GBzbX17iaGuD0bKJsnn7ZBDrj
NUb9l3pUHYESdSMueabTJUcwIGrYxdtGfScJdhyq6D3m14WpIJP1nYgAdafZ7bEG
CQfvRl027u45p7ywMWty8MdaPZBcTyIUwZxPaUYC/REbBIhzVewxvPALgxs/FH0G
M94erfG3S9EZ0a5uVR3xoUevTrENWa6Zqyr9A3DxN25rcXdIXwXl1nf90BzCrq6x
QqrYuxOkB1/+5T8CWwabpH3BSokavsh3hXdnQ44BcNC1D7I+nNQCkUvjm/58/LOd
MAy6EgKHIN6yadRLFLBVPNQsnanfPKY9rjhPukVb4PQ9Pxro33nYWRPQQEyNPVdt
GzmLguWPa1oA9aqY0+qxslgF4IJ5N50qCiHNDVZ6gOlVyD2PUznjGBXfgxASHdIy
6UOxh/TzaGPOZmPprxsXq6gZeP9kOtqkGF21uP8ZqI01XILfApScBq5HjEXzUrS1
T/Kpz9XmpMeykS84ZpE5Qx6yPdRLJLAJ6vr3dpMpWcTbDdvanm9mm+xqzPiI6V6E
buQcG1w7BofKsV7P9wv0PA/hwp0xI0uUUnrmuiKvMMlWduGbPQpX8N7jxzyXYQMy
X93nD6/MyAF7KxmQi4TMipAJK8AuYlUQ+yIwYW5sszBgHd7lX/Rrnn4Tx4MT0/3M
TfzD2bq2lwgtqyIQliQTehLMoxASa5fqlTjto1WfbbNtX4S5HWYBBzrMY0esOfKl
5Fu4cBLX6MkcLU7/XA2QGGSY6A5SEv2zZ2Zp7gM9ouk3xzah8O2uCvHzpU6Qw5up
bwu7jIrLqiRqFHGdlB64OY16jVxG89RZ+YQlEvDdOFQ9u6Z+Y4ugv84bMr1q/DME
5ngW9cmxOSq6x/Z0wMTZQz6CTN7EhFCgZGnv1LMLAAdqpkMO0ju1LpP071EQqoog
NgRdY5XCk5s7yiLKEH3uwZeMVwc/UpxJJpYF0A57WgmvkHAYBtogiCOG0tDSlazl
A1vm3i47i9Xigoe+fgOd7NDVstvXw9qI7oo14ATK32F5KnRbPLNjsJSTwbgc7YvI
pI9p6Gu09dI5qM85OJ90gjLrlcjacEurEGcySipA/Q58W/9Ku9ZWQQX/4C+YiXyp
40njrWw1qdLNKZIuojx1X34Y1AvO0uZRuYAyF0z3yvyiE2JDoNdB4OJqka48KUFR
nfYEXJR40z5VjZCs6K4im3h7xzIYVjSxcbgLY42fz+GFanhy0zcYD6xo315740JT
pRVWCkxeIf4kLelT6sYoMhptn6b+W6334nijItOBC+9qPbjLXc4BA0bthAEJueac
W4TyieXmAKER8MR46zk7B3vbhIh1FynfZLimkyRSrUQ3f5Cb+1ZpzTLNTELXNnkE
ByVxIqKuB0bqu38CvKbCIOrvzrn5C7F/FaGPMLqyUxgTy85TrbTBkIcH9bjXp2gA
aNgEGdHnL9AGYJr7fJCEwk8zFfqMOexrNhDBgO8n//KsprLVdybLAgPMMqIsOhuE
Zlmn+ZvEzHqhdsJPAa0sFYzX8OF68o9hvhXnSoxxljl0EpV+b6G8us4MpoxXEn+T
NGFjhG6LCEwwmBaWOHArUjmlyVApCFo1kd2Bjtn9o13Xt7iV5shpMG0Ilz/jsUJT
X80QTBqGin7w+J9fS2/b5SsWNtvkEB+4zpq8FK0BrUxMohKN76V1iXsxJ052yjWl
WMQLgv5Wf6FLEgqyhu53Vs0KTgGBFu8vBIm6NWrypnfAipm6Bx8wPaC7K0F/ny0t
o9ZQJ/FNHTfLFOJh8g6rfqVeUydv/xKZUXS816jFrZLY2fRB7Pp/1Rr4yRXZ798W
f9KzMYR8SWkBFZkZ/QvZkKWxabkzEDvETbjK918N2bcbOLEyrK2AP46gwiFf4gQY
2MrfZWsnFvTMP6PYjeaKSPX2rhXXmx9z33mNzCeLcDfEQbWup/mhdNSBmAi3hiUG
0J88VAuG0DYCXt1qtvFJbp8QkUyLmGMRt5WspLydoThhNj164xGNyHNYeSVoWg2Q
ml6XHtxjoJXI/brxOlbOA8xvxjXSlUtxu7h0NfYV/4dwUMpeK71vZsoHwLP3qBJZ
dpKiIMeBpqq0HhmWkRMApjK+TGfVGrhm5UmGyOUu7PRzAph2gZHSQWzd4VvibOsy
5OOPZMCKFHbtSB6MVGEaFWTjZlqwmrtzFm9RlcTL00c9J6BAEc4S3PNcs70gkZu8
WjMdknP7STSyBTpAhoHNb0udep9ZaM+FOj3GllS+pXVU701Yd7gScm3vTNlYuWYZ
VDAACLEm/+bG1KR7p4wopdkySJBLB2WiJFfvKyb0Odu/8fGOznmJOagLV82eTOUx
cGzeOALKGXHcXXZ5JI9vt8twee+prPCqC/PAxe4g2yhwx1SOeojDRfaST5pEIPmE
IqaaA6rfIiv8D5Rd6W1WU445icqfauvzEYRG0qTVTExwg6n/VGISrDS2r8yK4eYP
sUniRV7d586AdRG6cCbMAbgzy6lPWM0Rcwg7IjtPjLhPVLtZ5TF2+zKQOolC3/6o
iRU1G4+Vw9Pbso/jnYKTHBaOClEo6C3XVixaNuOKtyxOTZ7VZQu++myJe/l1OSL3
ufO81lNipSrJdXEEnelRFrG6f/eLhqqV2C5pkFXuF6NLsvp0fCpHnsQoubbjqwUF
qargQbL1zCHeO04mO3xk6UOYLTnKvIvfZ6KP5bk6eP5PC8+KT+k46PlLFwEbYNS1
8YVEj7HwhMfAF80RsDhL/YG8GdgFJ0ollm5BERiBwGXNWJjuOXlxrdTgEawapuu9
BGvKXNK/JqVHs1LRsLT1fgMWa/Lc06qVT4Tsf+7aVQUeKWI9zDbC16mSzRebtPvX
IbBVSiFg76QhEb7+BGtuXL5tv47IXoOQkSVZdcyN4MrTTukrNCt1S0rgaat1Zz1t
Vgbjqh/F/kDG0k9GDVjBbtSb318IzclL9WQYRFA8cesMP46nlNiPhqQ2ypF/YlKt
2VgMlLd6LiYzZWH8LZRB6PzVQsWvVOYhyuNO3Qvuag+x0K2LYCoYda2A7q+7JlAT
ujIu3PyyHz9f2R85G7zaW7YDAQUS7/ey8OsfkfIbRKTUJ3KETZnYtPrqVAGS9zSW
3O7dqcneC2fMqR5QfWA7O45vOoEITSjrA/SMEwC3YpzJ9SoQmuXQkbcdgn3D/GOD
bsr96MIDzXn93/ncEXQcwQbGqRLNTJPFNSSeDFksqMReT9LkgP12UvL6wyIEnoeZ
tgNgWaq1n7eai72I/fhRA8OXjrE14fjgkmi60lMwtAlCCb4vFPvNB+/XaIoPDU4Q
YERdI/N7INsygRAe7/KmoWtYw6EBpQGfuCMkkC3ozQgpcsmew/zChLT9UKyGoG4N
6PhS9aub916QvXJa6DH58JgRFerLu/qDfjZMU4/zDZHrN5k/2HbiQOeN8ywJFHUK
POZ+bPRyiKUv9EHzecktUIXWv7j8qOokwosPzOHVmtRiqRa9LeAvhwcQPAQnZsFH
qcxPdfev8qagQw5GJXCDx6d85AqmVIwcCxmLm9r5kWsolTg97oE9aE1btsIYwoVW
ZTQWk03lvQP2sRvPvOk2PRPsj0vWrgn8ZYQsuQI8eHSvIsT+FDp5BZNISKZYKj6c
RK7GCIFbj4tmtpJguswPOJw08cMXe57rRnLfNUuU+o7ubheWyGxzEGAK0exQitZl
MgN7aWgUvcdXLmxKxkfCozo8b5/dYE9im05OGurqscxOE30ps17O1du4vXZTT6KA
WZx5db04EjKpVV0uloflFM1gCn/0i2SHzWQCS+dJZ+ujkpDCbeUV/UeDE4DnTWP7
hTtSxdQSMLSkEYH7Py7Wv//hCm8IVqtcQY3aa3OGIwAk9SC1iaVd23qtT9Ooyk3b
E7Z2grfT2fVH6zpAxjf0KkjJwyuvZlSPrKRe2RsMDg3vbcOAHhyjOBt+nqw04cHT
8MBYBRYseG2PrortgOpi6twron6bym31pGCjJJ+Ls9mpe1svofV2B+XJz+ygzBkQ
vxPHVGuG4HBnar5IN1GAyAQZRDgLekxLi9rENrH/3y748EyevSU75MzJLJYLfQoa
r6vEAmHTf7qZUXNLhEisYzLRPuc7TnrrM3JwSeljt+Sc0YhW/juoi6F1ay3nMMDy
vboIkgJ1IdLbBbxfJKfs+TPFYoEeZ+XoavXOmwfjJ/RIMBYKt6Eu5hB/akMpU8VT
ZAQcxzkWvDlzgfjQohy2ycu9NzdnjQ8Yuuhwpxk8yE+th4p1sGNhqknrLo2Omp9y
y7XdVn3ZXZ1o7/iTlYiVIGiMxcUi2OR7USRqtJKCqPjE35qhdjCDtIvuU/bb56HP
ARERnDTEo0PNBsJZ2zAtP34aQzzcDQ/5uSLeTNaZMn+LMMXWgWDeU3oDtZqrwI0S
zPxgD1A4Zg9HOZIzadv2TifdrUxHYqFgeJHsoutShJiPHeb9NGzhrWwngMx8uVAy
Bp+bmYXBsqLhZFy4XBl0kOqK5gzMlz37HW/ZRuCiLyNQlTtdxu8eB9IqfL6EqBmX
D/CaJ3/iRO9UVJVZW9PFdt/aROPfg3Q7ha8Y8ViCTNrBGD8uQbIDVFu4b/cFx+85
0zN+adUs2B3mOGoIAhIxM+VqrvaciA9bsYdWrG5GF0gEfv2aB8l0jgeTxXtQvpEe
ZlDgC0di/AffERQMj/3UCLufCUA2iAwlgGniSl0W4wHk6xL6gE2h8Y7SbvoFf18b
jX4Cc2p65yc6AMXN824K6WDjeJvI+yfBGFC88qZmcwfgdLA8Nm4csfKHm14BwAV8
w3tJe0fgckTexstXfNCbhvkR4GHmshPuqxpqV3ppcg2/vH2kUR7NyoxsY7K/scs9
m2NjU3gq4hSk64l9lz2IJpSBTG/Rjqw60guwQkpiijj5Zy+qg6J7/fj7u0T8N9Jt
uhuCJfJ76PlAQ08+nf6yP07f3SVAy3Aff1taWMebfQKYjehazyANB/FK+1DTq48F
XGyerZ17MzXK2+99+bz3Sdp9d82Y0XbUus8R1UVlODqEbjOewUaErIaNuQSWSXV8
Xa1D53cY/hfGGS9OedCwbmn6Q3m2DBQFvXtXkOITslHkqLvW/qP5gkX/IZBe+oG+
cUkOdWY6aOt7QRssVWX7C0lQB9Kp0tyBkx38UpNYqctFHcJyTCVm7H8eA/nPurnC
bcEiuCKK7addfJ3jXAlm3CRFg/++csvD4paN6RH39nhKt5QRxsdFByWkcl+WYlVp
/+S4p/9HTkTLfqr8ILm38Ks1OAnk9JeoDwpQPbrHUMBrzxKXN3tC1udNhVKW7B0J
HcXE1vFJBJmoqQFwmdqCek9u9pFK3DzroBgGVjucL7Ybb7WlOuZ1k9UCP3Swl8+g
ipr9kx47ABgAnZ3Gw6v7azHsaXhfYKBisUg8MAQ2lYH9J1y47prWkUr42Yg+ZhnD
Xs+Vk6jUbUmAHmX+snbjI9dVMHc7U3Ez6jVs4/zJh4VIL+uiUTa31PjGc+iW+CUp
pxaYbfzConzLrSNbeQHcFSlNMDh38Ouffa9/qZ3p+tFRZM0nN16YsinNRvQeVm2W
n3U5wh84aO3sY7QlgtyRe9EBqYCSAaAz1SAPNYtEyAAPnRSqLBTRIlVCPcViHDaL
ZlPugXtbI/8HWit6ba0CoRFFBn/0NSK//0TQTwJSlY/xQ1kRm0ecsDZEpqmx7cpN
6xLHotUzfLIwS7VTOc1afpXdwauyLjhRPvUP833mbW8DNgNWZDwMuAmM6mHMBLmX
TXMJq46dLhkP6zPvbXAn4iquBdLP137L5kY3cHmMaNeolISz/vgXuCKMZhidujKk
CiqGD4TAv75NSEYc2i0fM317YuuzH7O4BxFzmPAcvWQ1eZlikJfXllV1QT7WPONP
r8sSUmg5ICDW2OwdJeTJez9bIhpDQMd+4IVarUasfg/itw1CXQ2kZB0KU2KQ3T+M
BdFx+74CsA1XUpT/2rVPco5QzsCTVtt82PnWy5/h38xOR9hpqeTDaKoe6paWP1ug
dEySvauYWJQm3TaqDjxgVgDkA6AOQtf5xKLxShRCrY27VpNrngiDcT8O6EfIruWb
qmeKI7qzRXy6dN9/+A+umOgy84p1CXkq/DPAJwendMm1xOZWyta8indTcv7vmtwz
HdeOSE3YDOXmmN+PUIHBmI4ZMjPHuI//6jIlmSfn0wVMKa6hc+pobQQqNuP2SmPT
EjafGv8G2D7fn2XtUQIOZqODUagUiK2IoRvfCbQsVFuGDleZuH8VrCHNMaCqdMJg
HGeGdxrnGNVtNXUeK00R56SfXEZUNC8sUhdkJABNOxP3Teb6qu1zpjfOX9OHgiWx
xNxlDey9U1EtGakapuz9SDT2Hp1Rnf+o5108/nOz1/H2h84mwkrKTJng9XEgikjh
mUUgHTydYPCFtsKL9KupLFAII7Ux51/le+ycx78DVlIaM2uesjTye40N9k6uEyg6
xAgHV89CNqW8EAxC0XMXYajLlj9bjA5ggPXdRoR14pF3hfJC4ga6F8qpRSrFngzR
1Oalo6vWIq0Sq+Pz/DWtrjXBSS23OAAeeA0q0tExEMEsM0HUPLHj2aZUr+CQlWV6
rfGUWuV3feo4Er7dDTImvpMcGgqtdEYWYi1PadQsq/ANa1DDvuRr6FQ572JAAvOw
c2B7o6hZrvxFNPPnZyPD9iqD96aWRv5/GyW7l2S82tH92el0lNrPoL/DT1HZlwir
qi2CjG0oXeWffjsFMrG98OkE9UDPQYnenN9fOCoUtqT7iEX8cBQtI7wPPsJ6fzKC
aQVYsfFJpW56/NVyQ6lXnwkrNN9UrlFBYuIEwTio7+J9gLc0IlgcOSLwQBSU0IfB
vrwk8AHCaoR24iesTCgovijZi27O6XmEoflq0KdSs7j0bQVZtASK7DuUqsNKnk65
3mIe6/jCMn1H4fpkhmuS/cCj+m12Lz9dPDki6/6XZsiOJRIxuXBWWHP2WucbYa7b
ssDMxXvPPNw8UVp0pejCpHJySpaE6sNm/SUHnGFLzU9XcHAI24CiDTTaQuIRr/MN
pxZ8eHYISem0jcEyagtQVU7ras9uK1FQVkmL3octmwK367pe77KFf+ODO+a62lAL
iH1QK+0gtnSMQa/RKRJZSt+4y4OSebWDEmDIF6G8hHJk+jIJvBN8CY4K6np6Kr9j
/6juDlo22YnnzuKVJdAXlbjGWaomAOTdiLOqNFqlD58oAG6B1kpBkX64ZMhuF0xW
qJNhsAgp3a2YVoZZ0Xou0gvHj6SSTDd37TFNvDYRtG+JgYKWyAPzVpajdxXOzvUj
gWhOcjSmO9RhtCcVcem1AVecdlxeFfPcXZeLfnDvD8LhiNgfEsfkzC5Yhj07bpGq
6KuX9f4fnA+AZxTWRUQDQGAngje/r8rA+X07IhXV2kK2cWTIArvMhxkCeM2INiby
2mzMj/jKgzN61UQaBi6KETJJfsHH+qaEHq6XnZOEn0VE1Kis6jGyG89ZfkObyJp3
C7IBtdoqvrnQsXrsvPEJV+7BOdwtZSED84Fl1Oe9x4pjtm3PBqVWC8Gu+luBdC/M
gK0v2i0woEpLCKcuO6C9RHopYiEFF0GZE9HM9xT3VzIQ1Y60zqrHOQ3ODT6HDBWB
SXxPdxE+WFzhqQFZ5qaOeAEk9ktYlV3GZFMVYux0zLyQo8cdJntX8UWufFo2ZCqV
0GRP73WJPGqEomCA4nTfmJz7b+UgEQ/BkLIP1rJzfBInYK2FYB3Kede2Ev+sDlP9
C5iBY+1lOxwZCCfX/LeVmm/0WhMNC3aBaQ1lVkENM1v5+juTsamfbksWRI4qJy3g
ee1f134zWiJiF2Ax7GpAmrMw09gX2hnNQW6/bOEWFgiapiAoCXaN2HVQ7SAakZYk
BATbpn1t6zWe5/dpmUq5W4B9RvggRVtOnCRauJ7L9PPQ9Y+/HlFPr1H6KZV20ZJl
LiUxZT0b0txz+h7IxezLWsPKrq4M1gmrTkGj9fXk2pOro1vhpz29ZHWW/XnUbHqk
yJSlXEMTmw2KgXcgiVTVmnbtNO/jut6UjzLxjX1mkzVGkmxbspastOhNGRQPRcrP
p7g1iBmvioRmOjmBM8C4aKkujvwd6qrGAugsF6eARZqaVnhapS5iLgsVLaLpHV70
+k2PRN4RxHaJzhlNqk6UDuTgziGKtqbs7XItRI1JR+BooFSxl6ZxSPTPt7y29Mq6
UiYTOqgCZUtJmgBOwuV+CSWo/j8/5EWmg2vtFFbYso35ZWzHur1XijtfMppzxnzZ
A/SYIRIpvnaSNP6NP+aKQY5ZIGZUJa4w5+wdTZUD/U6Ps/sBm/SdTy19L5ySeLVS
uhw+sEilelF/aWQtcc6eNW7WNeczSK6Vhy5ECcO6zH0ly1ZPF5dd9D+8OykDcG/I
nF3NsafdEMAvKKCwdD5f6PPj7qEzQU782Ovv7dj8jhPPrhSgpGt/kM8ayQpguPsf
bGMM4o7GRRAoQtQeCEZpwCOqd6aLRr75iC8pt7GJhx/JOv0g54HZReN1qBIxvrst
XJQE5yfAMGiCFU43B817HwuMO0FDNfDoqZiq06+jQ+e5afWqrmbeT2D+iUxoirBu
TpgKaI3Qs3e0wJm8DVkGKCEpinZ2ox/qFw8v3QmrEKtdXvnup5iGgnsFamnc5l5j
KzgxqUOJnbsig/2/V/qS9pUH4a50oz42IHYuNDeSjJ+7+db1a/kwOyANLswTiKKn
PXZzVM+Uz3VXUT8tFgefJv2Uk2xcPzsqD555+2cnGS5NrSuEOEsCBVDTF3AnLOsE
Qpko6En7VMrTbSCTMGq3EnaCJi5+27UXWeLEaX06ZFmTFioL0W7pK2NXnxUERjge
8dqSR+SN4r/bvk+3u0Ox/7uHD2x51dzQaS2OrkBzsPFjy4UQV8LrMPCDlrDHnrgo
Y9hR1Hael0BYrPbqU8cG93tssSD8K0IjkGku08+vvC5fIM5o3a/8ZLL7kfExe46s
ZBYnGXHyAWDUf5lCsQmgnts2rakoC3w4aIbnGvGw4O6GrT0ZGtvoh+VD2xEyRMw/
f/Py4v9tQRwdyKvc4i19N0WXHzMcJRIhexjIRk78+xzkByh12apIGEic/djm5Kz4
TZ6UEORo8fm5cOEOo3Qo1FAJNMru4W/TjUmOqbQuofprlA7bcDTO045jPf+M7K1q
vR7F+Kq6KmSDqR9H6nVfwi0gX/YIoeQClDAgpZSEiMnPQQms3FU0sgA5c+AlDDlp
z/s2Yx7fomuvO/bAiMMmSxeFB4MR1YCR1e0fTVcSaL5l4sPDpA8paGWoxPeK9Pf9
W6YT7QmzlfGe+lJz7XvtGXsAFZPvO2azIkMYihtwaGSLjmdiQh4Oe+B79ef9/BND
Ob0hz3vEuBdrVCtQSA6kJaQuIwB7ucq5hl3cF4CzlOCTvc1AEG9YHOe4FiYPxYMa
0TsvV4x/D5mHq2pgqTVYo2PUifPFQUkioKcLK2jR0oNriEQrtnSpBrRX51JNV9er
eywhaMPjD3tZYosnTKxAgsyUM8gSZRsADFcydazg5p+bylkobgAGp19SKN7IfIEo
MKleDVhxwTsDjsqAwS2tDch9ZCNYuXd6j+wKxwVPa6sSFhDAtydrfVobGMlMDmqo
kYheqamHuEmRUuoXhMyj4UcFSHhgQKHYLyGkHssYmcM79FuVTRUHo6aqgHR5pZ2L
eXCETJvs38TdopuML90iSWJlQM7VmzawdjcC17xwPafrDFhD7cbX8vgsSQRy6eKP
+bKDx9Rk0N40c95ORW81+Q2c1B9tZbV08Va4lnCMplBGhIWMOJGpoSGyEFEHCR3F
iAiTs5VABazybceJ16MXAuThIbArRKeU3P82MRs0Lo9A/XOPDJpkSZSlL9ofl8Ig
jWVhkmCs/TH0frJxDYVhLQ3MvMCEKYwtGGpcpoltI3tA4b4/oCF769gvnAxd3gWc
pqEqn6C45nQ5JzBOzc1wI5wIaqkvd2tnDlqImIsdg4RbAlY3Th8aK+rvuo65LUrG
lK0NpdvoXLWGqKZEkxr8H28W+C7KwLqrdrqmjEWPv4DEp4E2aF7syXAW7J8MBhEs
Aj8cZd/vdG6dxHno2eQP8S2Ap+ZQ4k2Q4UhyVEvaGvdHyG4wYFeTrXTtQe+H1Vb1
NdRgZzsc1TNOlX3SDxKdhFcGFwj9CMOGfjoSynzuQqqVn5M014GIZKSPnetUYO/a
x2uKApoSiBpyN/tQ+Shm4nRhpK6jWGYD20Qcc6QDY5LJhuWfcSCYlPcsXbUG/fDs
yAhVwe5QOx5uS0pyqMhnlArNON4jUqmPeFxr1IdfJcVfAkfIq16qPUw/ZbCF77bY
NtH9V1AFAKmEW/M5cAEv5Dl7nQ+p3akrvC6naluR9rQ/o0pDmZdbomfy0llmoJdW
eFMvEDrBXg/M+CcoZhb05/JNFATC/SF8BJHslUy6J2b55Cn8c8qQyuwokWT3yGll
NlEOAOzBL9TDBTfijVwLfR5DJhLVdZNvbxvBbAaPreUxCUphfO2Nd5JxcBZNatBW
Sv8PNZ0ABQ4rJ8is/zik+/m6hN0x3r6YGTyDHRJgDUnshzCUWuaFWnmDmZfZTZsU
pMOMeAs23A7Fu57M+6tZ5g1TKZaODnRh7QN91P8kO0HZ41RI19gEliquJsZrPwRy
UN0lNiad8bXVdUvCCyQQsdrxOtBOACJJDeS2urq8Khh9SANrIFF0nzo1h0QmBIvL
kw8/s6OdPdRyGyk7YYK+LqolB25kyXNpRSpIQvqwPM8tOGlbJYk9xBNwQKmUWSCG
bIR8EhJfyMbmPdmHP7sPy17KGQIc4KPwE7j7JdMHhoP/CXmU+t9DgADo/F746pje
4CJCky9iAdaUSrP37fdWA/rbcZ9hQwo73tkfTHP9ahn21ff31vzdm5m2BN35Z5LI
4Fetfm6krA3QY3hr1vH4LzMReLZ4LeYMCCYWsH6woSCOX3dSarWqRR312oz7DW8z
+/3M+oz/Xp+er/SMmkejyBvT/HhNNg9mgGVI2rE3CeMLlTiac/EEv6q4B/lXtoKk
eMC1bqH5fNvoMNVHxjnoaZkIlLgpya0dZ4gYoGJohMwqIrJBt3+qfoViaMVeFhdr
noGZmNwPwICrumMEX7X69aU6fttagKubHf4wi9aU6BcHz2zq7OFc84Z9Uglmsdtj
D+5ORC+UCb7+t2a982B22AL5UheczwZrg7gIHsTkon0XksOLjuBU8dEUSNH8Js5R
WV30WKP7oaI/0FkaPbjmta4S4rNMbqUmmxnFPK0tlxpN8cp7UEw9PKHL0vUX79+f
CpwtgSf7y3ZGAz5Jxfi5TTAKLP8R7KOmzMm0u8d+dfmwgTS9T4SvDHOzgvr/wdsv
+fybjCxsFn/hzwlcjKGycxr9CfmjqaCz0/8fNrFDc3jSlKq4sUgvZQHwAGpq6sJk
WxVXIDslR8yq7kPbJtKcciH/2gIYLcqj4x0QVs4s31azV+2yatFI4UgjnUh83Mdh
OZW3K9WNFoO5EmYSV6TNAhxYtzQljjPtCDC997JLVe/1MCffFps02d6seJSK/1Ak
UEaQNaZ9UaHb9dT00/4Dh0K+QdYYcF7KtdjUWq96upl1/YUlzbCm/YRk2MdQXwgF
w63bRChGF9anjs9mWUkvS7Le97DqUh4S2F1BphelLG/FeN1ZO/5I5AbHxflXAaH4
4D7G2NaLSqNNP4xSBYMdjnLELoeiAEP6alKrPJUEtaVNYjdFNfTWLvTDut6r18s/
nX0G9Bcql5GuUE8i56W93wTUGMllsAViqoYJp9CH+QvsgoASxkHEoSPby+JZXiGL
9BZMOBZei6wdLpLh4yV/tXCpSm2GCxWBzNCUjnoSE2QDShzz3CGUbvQIRXSzFglT
r+byJUbwNcD7vkY6GJli/HlVTDCsTu5gHcTh1L++jGSwyTyoJUerYaT74BEJeLm2
C2rps5PwBBGMkFL5h7bliA5um3GQpDG1jiCzpEMf2IRSjRPQ6Kf1EyucOCaiMmPz
RPPWZ2j9gY71d3xiljndxHG3ZJKPv3B03+GXMA0GDTqqTbrmegCcE255jQflZodO
6yv55kNb3sWzh/NJrTMZmzVxOk24PvPhq43798cJSgJjyWNE+tdgan8uzDJkfExj
EQuaf4bwB3ep9jhnfTX1kmXmC8CUB3YSijeCJVHP3ukuP3a4ziuRuZZfPS4wV5h3
8MZW11Yu5vmQ9Yw+Jn5Fhwu8fgCD2eldHiEEAnXGkDgM8t6BKiwQYotQfeghz5pq
MPQM2x6J82kp8C7fCgKoT0qEPeFCDKlEezEOHKdzUDNscWvflUWkdo14BPJPxCYE
WEz3bleo4S5auLhDpixQeS/pTnawVow5JSRR2TVSdHOlQq5Y1GidHx2Wv2AsM9aQ
bdFN0MFtWK7pNn8P9xvjFYxmiFtWUnT76OMSqpqYqCmI/PEdXHuYCFkIJg+6Fvmb
KZWLBhq/dJtSmk4naU8wl4OI4c5cwTiCPWQvDd8ybC0N+K+qGsRmoxluc+oUedde
JCKv2qccU9R8OFC2i+TnyHs4HKbjGHW25d4k+660AG6BgVgHv2ltc9Eh3s2mLwei
qiOU36XllahefggDj3UWmvwUhqFgbbnA6urA68KCEFSLsN6eggwtp3PKAOes+hVT
s2hciJGe4XwmSyjFu2g0QmlAnfMuRTNkBfsD6g8sPtolvrDVRPsE+fKwEzQHO8DI
DEjdT/eYh0Yms5GB/K3n1eJG5M/ce+so+k3ZTCWZOfwoVtXZNkEg1vQincatdQ+3
sjE1wk0yFXijYa+E5d/uxJ4GlJy07eoke346BDaoLSIvlA8vC9qGesYET7l01qn8
Mj0+eeRVReqFgUmTpL0RTyC7nTOjmmILwD+rKWeDCzzsFdTRW/2hA/3jIRlWojX2
J8OZqNm32n4KAtNDaaALLcyYqJsM5Gw8btWxgAtws12MnLrU12wqo0O8keKzUAsd
8/enRvuxGiAYWUcilhhFFPFI8Kwgy4qU9A9bGcEPnVmeLvlUQrYTmQwAuwm4hLqq
4oevufDi4nXnosr6KJwwu0cvqAkSp/31/t1JTBJ+JvZ58ePLwFo9gMCa49nqS3Xk
7SHdlgEhDuORTx576zk5BxnWzayFBWY9PkFoC0aHVUV1pKu9olyOzpK6nBo5231t
UmlHN1VgJG4Tff4syZHQ1i8ccvSagwV6nhy5C7aqPiG2mWyWoYD4bo+XWDzjnwGF
e8cVfTp2JUVeXcDIo2GkpaHj5YmxcdFjzQsgt7lu2nVa75pjiDCktjSHm23soQKN
FOJLlv7OeY18H2w5hb59ER86og9Iu9h5P0oqwzSr8SFWkRm62aR8Gi/3TmfzNnF4
/32UlDY63Mt97hhAKHp2v6usYblLC1s3gubXNieAaAWIi/d/XoMfqnl5XxvxReqX
BXbo+j+3zcjygz+hUwVhIWFUypFQXsCLyE7mC1dJumNZn9q2U0TR2+8EkdaIcpC2
aPqwMUuZRq+QKiweUJRpNB8bTzy3dca9mjgbvXAolAPGrpFW0gtTvxUCimSOeKAY
01KlqSZAI8cKcHz/g+Hy0VlPYwxxofqnivtT0cN7uQyAEV5wpifeErKPO4zMBYQx
HxmP6i12IAGBVIv0SxKJeU003JvpWNbh70e1p3Mvr46GyRVK0MA/lDZlbx4Soq0v
pktrFrQDBBhPdITBbqG6u/VV1Q82YSOOs/XzEHWAF49WsYId9juJPeHieANJo6Us
3ZAyHBAFle72N+Vvee7PPn7AQHhQEi7v2w3376BPvEwsXNWV0wlGo5rsnwM4Hdvs
Pu9S4P9CjlmlkFoFNJ2m1fdC8vTmfLG6bWmYhcbv7pQ4J80WPxOfvFELs0D3l98k
5x9Tv6NwfVhzMFY62lwZ0dDAoy7TAoJ9h+ZweIgU2J3vqKrcKJ3mWOAtNhE9iYHA
kSIFeRNNyuaz/aotTWoHTDZfDpr7kKyBJVYMX7GrDBRvvaZ88LWXA0YD/YD78dex
zZ+B6qXKx0c1xYg0CC2Ip6VLhg2XBd2uG8xyBnrG7fZ7KjKA9TWWarrbNsFdTeYD
vdcGN2AYSGTIIr4mRrpSdKDUjpnVvJbF5/VNBHQNWdcE35D02WFxXZsYUb77uUSL
7xvDVDhSLHq+IJgW6Z86FjRfX2rDG1wmiim+h6VpCSYBdhivJfS5q6vzlts4fCaV
uNpYI/zVk3AeojRhfN7qCzQWH05wqPYazP/rKKRHXBeDs4FrgAZc3RllX1gcHzMo
PwfcJjDpcCIx/m5Zx60lvrlHyKIrEEelmJqJEGK9rzTnvI46JMopIK1qkQaN7NkS
ALA8tCPWZ1Hj8TwMnB1/yGCSS78ktSoph6ivLW8scDAGeV1qylfXia15HW69yNvg
FnqtwhaCZGvyKpSP/tTGwFyKxSeY/HJL1lFcKsbyuP32wor9TYuiddXmhXQhn+pr
dU6jyZjjzv3cjFAmv4mv4oHSov9ZkcQLtu+5x8v2SB6lJ4+NMei8TftSqmr7IRU3
aVe6b9lZesTtLzLyljrY7FwYW6tGBIlXWcV0wpxdOFHSaWZDLODjnUzJUmG7186g
G4gTws9iE9ZJsGnJJfgupD/I3FZ2ddRGs8m1nq5s6/s4TZzaGYUFDqDlqWCeZtOG
HXsEp4oFj1DfNsqz1D0jON8cJmRxYv6n278nlof70YbPZ/8IOF0xQsqbAm/gmNge
DPzAW4QOWP5bWzxheJUoFq5cODygRqtvtbDO4Vkozvw3nnOLfGy2S8Y9vXdgfFvk
wG/d6UI6F0OORPTenZi96+ITdpLAck/yCUu6R8k3v5jTaUSj8oDinOIB1IJFtkZB
eTvG0EzKonoAwzZmSWdmmYCDScyVIOJg6D0uw87hErqdS4SUQWSOsJPHWjIM0LwC
9d9Y60SsJn4XvJ4Gdj+FghXrwUdCcDOKRkSKvyjFDltLNOO7PRiqysN3d7gvTyoe
Hdp3CFB9BZeIbrU6b+w6hyTc6GHC3+jbIGpffvFKOe8fVx+0SUPjvwdQE52dLK8E
qvme9vum5UgTvmNHg5OKRBaPtLgC1UQEDiu77LClw4ZYN2kQMgFib+LKnpxdNRP4
dV45iOtrtbXPUAUjf/99wJTwSa6O9hT7oiVdvaxxnaaquXu3noK/Zv3NGbn/TuHZ
JPMY02P6tDUTMUOkRr6jzLQedDyAEHo0wQAcsbLL9FC0okTKqpPcAXLyqMPoA0EN
Szj066YBQ9r8Oy3HucS+JNjEoyRjrn3u6FqpyXf1pYnsbX/mr/h64SkT+T/lwYIU
9am5VvwiLNqw21eoIAdSIHkx/ijeuYIuQeY2dOWBsyaVtPossINI/CsZg794FqDX
Ajn6EfCjNt80GOk5Jnxl7ClsXUIOJ9071UFS+BkWagAadUmnDWyBLes7IPsM4huj
o0tohsfDQqXEucuhBzqlIlhKNTw6nNdzbfP/T0AAJn0yVjukxUyLSQe9T1hrMEe3
UwNjRAeY38Gnt2BsbLPCVnFcNGyoTYU4RjlJrAZQJ4fOnR9XRsx/VjBWLRbSi1Ex
1/Y1J7I6Hju9qViJc92Akq1bk+FFmzk2q8T2LicoDL9JjWYx0Zwd+OSw65PmkevE
l1Zs81n6YW+UcjYCz/mO5SGfm1GIN2Wb5n0/NR0HXhl3+PlNNVLkVM0PgMqZKjdb
qXzxsypNSRyMP6TeCFR9V+kcJVmZ6+i1y2bYm/ZW2O4WkQjsPX+HEXMZaQSfRJnj
gFNFDKjZnUpjp7y2l8mnlKN0VqE32e3kThbG85uHyF9dF7ctomoUD1rXKURr3nmZ
5/6UCXj+NyZxbhbz+Pv4hvIbAv//bjikzTeuOl57RQjnW/LF18Sgc7gsoNor/CEi
dHXnaiB3lR/8cYjGc8kCrPgb66NP3MOF+qx++o/wwjif7C5fyiKZpNH0P3zQAo8c
xwU177Ld/P+yEPNhHMWXlJoEuyLbKA/NWufYGkZ7EM+3SilwyRmmRHh4slfrHkqs
ilqfFnbRC0Tv6h1SlT/JgR5AQyhsw8/CE9zWWARzHwIlPxkZfeqodDDNehH2p3lX
9y3r36yVCKgX3gd//BgXL2SB/MUOBYq3ORiBBFqnGI93q5mnx20LT2CTW8Kwtzkr
1GmZFfPAdb/uA3fvTcEJupqV7O++XNGu7AxGUhnKvD2vjBPGHNzgOeGIa+XLH+Kp
WTsVWloRi8r305Non9UOECRvNqj2wAvlmb28YUssXM4fWucDP83Im41sSaVZHI8M
HMJSCno8AUOwiG33qGyRLBhyLGSR010H6kdBvSsftgXASeBD5Fe3oUaTKc/2sz0F
3cNCMtYalstecEGfRjZi+KFIh+Y4PmgJAlkuEnPjIOq1KIY7WJWTrold9A+W8LV9
q8YqYdfUWh00+8trxrwe2ifB0mxjnlawL38DVhc2GFf4JMoRxKRHeOL1DDhTn8+s
6vxHAjz4vMR0/inpELr/RoRVORaBkdi2sVTqIzR7kmjrvsHgdd4xD8RfMcNkvKrG
Yz5d4x2k8y61LpDy0N/FF4/09QEUfcg6fKIQNDhbSD2Gz9wN0w5q/XHp6EVjrzoi
k9oP0kYCjvbLPpzFf8B7A8STPYiBQqlnbOKzbxl2v3SjE9Iv+IputD8VJbGUwROE
bejgZ58mqqbyleHZgzfER5s9waCrB5jTMaIakvhOOKhur92+ER9M0bQCpFPz62aV
RiTUL26foLDDPiYqCJtSBSAlbNjcrpS/0OjrDJSxpaLUa9Qfp72XxwtTo07r+cQJ
unR8GlcSlUYVHkvMluwZ9su3i9uWE+ZLwB9TalzVJWp6EyYOyeSzuyDgoVeDvbqw
eNxeQCfLdz6zxW8sWvah45NI3iWwnoTxl6fnNQaFcPWEmzRuAATPyJt5zQyGc6DR
kKM3H39re2U5521IJGZI+RZYP3En4ZeBxPNEKDXN/fvOtnA/fay31AO6iNqJ/YF/
mQCfYolMJfntPY6sMO0HrK9u0xZE03Izjf8TpBtN2dhglWCjftwEoPlbnSb4I1dd
3CsW9dGaXOdia/UrTKtRqBvwBB2HK/INrypzUfuJA93rDKAb1q9FPvmmLGOdTq6x
+aQKpoWi4g+eoGBKX+LE+m9pwIRTtwt4fCHkICj5tQdp0NgNnbpAtLMYxjww7KbW
TjoEFVTz7CxHFcq9ZT6+zsBHn9lMBeFFQeaEzjXaxMFJFxePyCSc95aHm1fSiSbd
D1q3j2uducTzAwDk5jWeZx4ZniFgIpJgC/foqdjuPLM/UOFZTXsJGu8CgfWGqxq5
tx5/z7yVuF0a/SI2spXXEEkSLeYNEYVaXiN9O20DF4pEMMpMWpSoNYJO4CQ9M6jO
90adB7AipHH7/wvTP13yHXYVTfabnsYmOH2f45vxzQ49/OQf9pALRXU4mI/tp+fx
U3i5aDzBXtOpGWdfITMUSaL+o7TPha5KJ/y7Q14CRBRJSRVhau3WFh0YgD8F3cEj
s7rhLaihtvGZKJo+HvjU6NG5M0xR3Ri+g5k7cbF6mb3ie4Ym4KVAiToOiheJQX7d
E2/DOZ7PI/wCfdmNH+8PEGS+l++UOKGgTncRCh7lpkLIccfb/FtwTzgZ5Qupi+ML
h4Iw6ZEI14BMgHBw+aE7dxdpSDlEvanAPJwjDbNmRhGeSjKjy0cP90zs3VqEuy3d
ypykDgEJvnMDOkwjFDBLQaWpowepZF4r5UBtatYH4AGt+7QDxDAU9BMo4Q+Qk/gL
E0hIE+k3gAC8QSpf04riN73VtJfCF58+4uaZAbshW+LLCKE0591cruv5U4PnyB3G
0IzK/ZxGsGw7QQwRZwgp4oPBsEyxq0lsjQDJUkr6+QvqL7XY5UgyJr+uHPiXZwHv
uNYTo0+b+HFk5+Lyu4dGKqTM3IXH/+RDNKYppJT46sch57826DrylOUuxRVmspps
+tNi+L6Nux+FXt3u9C6TdfAgleSd9PeZpNSs2k2qrwimfXp9n63wkQTokca3ENdi
b1isDiRJlCi5K45ZstUOTu+sNcuyIwbsel98b5MojrYBSgYxkwNsQqL3+NA+yATj
2Cp+rnyOcR520JtxMLl7/kMc4ojKjVbH3Mu3czIl5PgsCMRyoLtHQfBk0BVfsjpq
1JDa1arLChjb7Q2BzNLZqMDvYI5yTBJkh8owZ3jvvgYh5vgPGsJbCHMzUyDHeAGK
6ihn+jBFFDfI5jQAU2IHWw3LnkfWaHPtef5rO8Gn+A4d0p0q4PQ/8VOVsq1J2Vf4
5ftU7mAf+zpHHcGQJahDXVbgJG8law0wINVkKX2DSErBv0zJ8X/pEEciLLWpmcik
uVUs35rSBYO/RXZfYPFy2lB6Q70t5ilgMvmPxlu35aljCq7Pa7TiTXhgXHvqJJWA
Y/URvliyy9ET9wxAGN18ntlt0jUrfBgg34KKSxUO0MMW76DlF+gBb2BZnH3tkHf2
nFKhmyILvo4zAwl4FrKECaZ4pjnntM2ii6o3aCNgDo1RMAIT282c3q+hUUql6P3D
S1ng0LJ0ulVYceJDP+1VG2rh6Y36JhuQ5tF8APGWSTW5Fpb+lZ++0RQb+dWoVb1G
eoEBvu+dSnOrApf6x3NAEAVm5h3bELQbQR6s1NQHol4OvrNkW4eKySwIIrkL1rZ0
lcDkn6VXCB4btCjM42LisFkPjn95pbv12vS2/BFPuOus3pZpKZrXoWpyA1tj7swJ
rc2j7GvHqD8T+bWBSCVh5olBN24Fov4KqjKQCfs36TPHrhRAuo5ehhhf8ka44n9q
M3ZDatkjCVwe4YGrZVzzmzcIvlcDvD6qs22+Kcgyi7+Us8Wp23I2X5OFd2eH/6TW
qDdah+JTtLJnCeF9JJVwWmuGP3LkxPO4zLGJcR68n/vXcXA0JUQbRrKIxXHovPIW
4phkz2KcWXAwEiCUWzUEAoJGr3F+Hd6P+4qjok5Bso4t6tTtjjE8f9zNJjPmQnJc
cLJ59wT+k3SHk9S2WZt2z+gftZoHq66zILbLv5hQbYKPxidi+vABZXus3a1BnmO3
fS2tcSeGO1rEq6G3C9MrbxQQjIeXMjK5ytFYLtKEfDvcdYZyLmAt1VB9BprgVHP4
YuTmacjT8LgZf2UauT74y3eiSdevH1niRPffxeyFeieQi8V8FVhhzMIZFmWA7O7Y
1ZuHk+cB5gPS4/dmM7AnUu1E5HYdg20Jrkiy2CTO8l1Qpyk+yqyWel71Zd4//J6x
bCQpknMwfU1+YPyU9jV6Q8B7fb3wykjaQC8KDe/l4ayaz42Zihf90w9CxDOjX0zr
zawl39PV75w5+wib+oPBBPCSvrnpHbEpGmXE/qdKarUHfMsRshHyqrgGvpZtTBI9
/AAIdQkQueugrVyhYO6i067x6SvcxYcDRi20EG6u83QTrb+qcOEoUEWTpMZewjDP
r9njAISNsbNoxOqi88zVrN6YWaEZHZsYKpQ1WJozTSiu7vRyzLO8gwslH4eKszo1
mRhPMVF9h8TqYJvgwknTaZzhQ7N8yyxFF4rZb44bcZpSPiQj8jQ1lnxEDZhMJeUn
G2wy8+lgsiDbRHyDlKHJJM+azxox98X3uV1oubyMWLu0ff4O0RkSQ35TT95EJX5q
6pFezUUNgLn1TCZlehQcS540t12q2D8y5RVMQ2Dj3NJiMcPX+YCF6S6CwDB9tI+Q
kZH2pGyCf4tFsLcuQUQmjykcklB1GkevinpNkKBZOLwBDvbQzT4zjDPxPejrQl7Y
8VgyJCqqNn3XuMIxc8pImbomdUHa92JaInPkMDpkRtT/Tjt1oXGIzfcC/ZWs9zGE
LfT9k1OJ4tLr5vxogU1XujrTsLvDHrKjiejh7Bvogd2ADNClBj/Fe2fy+ao6U2JQ
GGmatpWWxptQ5Dps9WYQVsNe369NqP0lgnc9YjXOWyJBHSlJxXQS16RJ/uZsrOw4
N98waslMu3wJ+gUAEQT4JwSH3g1WrV5IAWaaC8Jpfv+qpcQUYTW0irEEYbcmi7St
mky9Sq+VqBVQdhCnQgF1xkV09UAcJVgMOu8nxs5oX0TV1XGsdLTN4qjlhvukTm8L
VQtXwU4fikM2gb9a212KOLkNIGA3MCsXLGzHJfKTBwENQnJfdyV495Nky1VWQnkk
JrmkHZHanR2TucLWRRji4FkuThGCWG7xO+3yoAPPTGx8JmvAtBfTmvPtsLgcfpu9
jFmJY104b6SieQ8igUp3kzVAvQAsoCQlI3mN45vYDcFKNzRFcQjRzn6Nd3Adbznp
1/O6hTgdi9oSyWIIWu5VyP88TkHIn6Z9N+E2uycoO7BsuSgzuUmYQ5MxktzfQ6mZ
JKVHoxdz/J6qVQRca3WVY6lhiXxRaFmUOSAPkbslJydRh/W8CD5F6+w16GpjD7nu
p1Nzy+Nx36xE8zeL7kStYlmT2eUeIklx48bYJ2884M1ygue3vcVy4mf4TIWUtmtI
KZwmRQoYQwGyMR4gd7DOtt9/GEZKeQhs8Fz6JvZeFgPJQIyxLwts3Awuejd/gRQ9
nFjrc0ubkmntOVkuVg/2VSEyWdJDZ405UYGKQPBB0UTRn4jQc0IfWagotB6AHg9E
ZRfgVhMQ7/c0oNkbwqqa4XX+1jQ+6ZlLdKzUUhApMNolaBNbeof35ONmY8Bd3fDo
RlZpFQ4KCuVgzkbPNUnklI4cNbPzbily6h9FZAvGN4XPo/F5PJloNWhD9ZdAOi3j
eVbe6o2CYTCOczfYjx9Ae6BxAwjwe+22Shhm24ziVBcJxqIG6Go9EtTXX0c5SzKL
l8BIshTwHBRIfND8snKrDpSO0bT0ZFLR8caW07f+Wwc4nqMKAcRUDUZiRGgsL6wR
dnyNTyOgSjfRB1/r/h3HzfcJEvFzpZ8BBTh5V2bdhoWnUUSPJV11U8R+Agr6PjQa
qCWpPVVF+lFPQCfwOzx6hWDzWueJe/GZOFlD3TP7sFxRSfgblkMUdUB9H2/61D2M
b7ND82QbgGPyTx5j/WRcjog47wPuIZD7z6lD8+4K+DwWceFvdXkxA00icJV0tCKo
/gWz8kL2OPC6LMsog/dICFEz/uRs8LX+2j8sZOP/5SX1auFB0db/SsYwabjSQZ0e
ZjUCSvwzMsAN4UsWmA8f0et8cCXZLYI5ajOOznIpIrNFe+BEpmzUpgzFoqL1YjYB
0ow0DEW3ILxyQHsejZo2IraO3clNdLO3HxgRCryw3+d5xgM6ItpbsnAOFZ03RnZL
l9PfTBejmAvKhCB6z2MrBUwfgQVPtEO4g23/KO0kXNjGZtRd9SK3RbzAtddUU31f
XHLgA6EgcSX3ATr0f71URyRqJ7WRTYMrOWsTf0okT1YHkkuyWMptAwqzJGNxedKf
GIfYwOxMfWhFjZWSCd1q4PEw0pEB20n1X20Izt8xaWmRfeq0F0L9rqu7lBNhpO9N
vATon5k5TEcWZacGikZn0+KPX2tWZf0JZ0nWRc5RTUkxDm1W/8wD3EXZGCvYjmjs
4Qkqt+XkypQazQ4bF+vXZuQtms77Xx2plm1mMI4Kl0scjJfXJrCHP8N1fuXkrV8P
8/nG6y21Ky6cq6YKIJ5c86Fyk+anQLI9kFu4OTjOUOLwqhB1zR2VB1p4o0gv1moV
mzqqbuVmwlnlYdb/ULsyIKQEm6eKNR6dpRv980+E9ky4+TVQ2oL+oFQ8y5TE8/wb
naZMF8IbaafopRzPkT73zABzvsNaMVoQ7RrquCxc3FfJ24A/IxSxlcGySWE/lqix
v4Dbb0CcnN6SjxHU5K+nphF2iVIaTvtZOaLcLAh6e+POP4KlGVEX+mKGi2SMg3KB
RmW6iuak8MntLFFUtiDvM/lY1dD2mNK7panMaVTX6gEnWSh30obKCgyLZx5O61n+
+tHM6wzy6OxsxOTVWj5jw9sgilqPUK2NytnzHkiXLAMiEK2CrKgvaIsJgdei1J7r
pSjyQwaZ9LZaxEd0G+y9SJX7I/6ayVgKr8RnzABwQ42Dfv6fBpQfWUmirnOxvByN
W/Yt6g3ZqLhtZii/dtXiAcHFkTSDXCOo0PRi8kMCazJkcQ5DN63p/0FitdrRK3lE
9qkk3nQHvttqv8qYrtpRMM7kPmIlmNaF9hwmd6K8xQcEYlPYGbi2F1CwM5gpFF85
3HYDaJeqHCGjUg8eBqeV+2fz5fSWkgN9B6xnnt4SZR/Vfea+UaD7/wx9Bk5vPj97
bkiAFmHiJMMsPKfOBzoAYIh9Q99R0wBVS4eoKfIz8MLWF100qlTYnlwy9lfHyj6/
Qm9qrXDiPcFBLd6OjQW1Y/J4FAhBYdFtNU7c25HMPjnxLGvJiTjDTHLYw3L7Hp6y
vdJ7wMoYteSxP2us5Kg9ipOhkbFdoAGU0DfX1uGjt8xn8jXWMfs4gccIo6TUwJBe
hUIWTlQSBmrsAjGpl19RXbA+ykj/VRKYIqys5W4js51Fx5BbvfH6xQIOwRxRn/wV
5S2GOXQodSULpTZofYcIq/YRUwwa6M6DCA6eXELm/2W7nXoWh2P1e/mC0DWpHHDK
fMOhz2ER3QSV/tAOdgFsvOeMJIN7tMYwPhfIIVY5nRGCv1T4XAnY8SX6I/m39C+S
uUbahabYJmkXyH0oEt0PKnRaDKkZ+aTSeLP5uN1itTCSQfYHVGOsKkSYyRYRa5vz
JykKT2RFA+B1DbsVMMHstOTUWOC+R8dKRKBpn2wLSqyiXvhcnL6rM5v9esStkT6n
/BA0hNz/2qw1QavPeDMiorF0ghAbJugEvApCBzZ5HUrpq3fGJM/FbQ17Q5IhVYW6
0Dmoam0taN0hQUfT0ISmkJ0t3yO9hR0lwSLVeV9d63VLT8AlRqYZGkxl3mQgXZIp
4EdoFmNmMr7sdZsrDFVFwP091nRrCTh0P1u8nDEKh5QAL5Yf8+8py+N9mxBbYQVl
94FJcGMJ/sB7Vtx/24DPapZKLM3J0dqSXZYd295MqxS1TtI7g7c6QeKDxnp/7R9v
rFcvja01yu//UcQB2WzVHOLeNWXkz9pDsWwHZ/P2tp2XAY3lKP2yplRbPpPKyi5A
WMOmI85KKsgUvz+IcSkML39lOnQVKc8OPCOr2qIPoArzo7hO3X7Q9OrfWLX2+x3r
ffY1wgIARGA5krpDt6t2YzMECOJSFeJo4q6S3s09r/36qNBMqRqxP5OW64N4HDCh
IB+mqiq4YTw1kp6xI5cXwBLymGLX8mTC9Hhce2Be9VkCDzd0XaQe8rwgPcX/I97V
UkTeaGb6H6T7RIBw3+I6Qbfz1vIxXg1fU0rCDRS6JLHoMQ8dtre84Oy9Bf5clnLv
8EadNTNlm3gTxEZBgMa1vHkoWUygowFvf457QLJHYDFQ4dADJQveQMk9CsykFLUu
El27d3ym2G/YYFEFJDjwrjUO67wWCdX66zIbjuKukiDX1k8cLwAkONqXmaqRW4M4
JH4wJHRMWB0Y0BnJ35K+E8LBzZYBWH6ZxfiFkV9xdPIHCXe4Bkq0g2+VPiK2BIpS
3KUtu9Nkwi1X+lTkafUObeHA4d01MeI9hYv68JH3RSDw7iocCsTr0LSEQ+LI2akG
un3GbP1rprNJ7ntx8Mkay0pI7aE4b5DL7C8krl/A0GA454bsa7rD7MrcmgxSSgOj
K0r7cQii/yI6Hs0S/vYKy/Yhr9MSsL7BBBJt0dzsy+2f64OpEMsNOEkRJDF1JQk8
bogyTaY0dgztqnm7C53uxC8xLwhsvqo4Nax0uqMzEp4Hc3HanZA2wfg6t0uDAUp2
LYyspVU/hg8bYD3Kd8/QCz2QY2MuleSJyrX/beGdK1zvOZmYYv/j4O1/7ueeYX2v
DEywUKkSHqDZbYVxYmJ6SWuMzeUxizupkK4dy3JWlQakhzIY0//PCJVl31RkGs+o
D07PHUaOxd0JNcmnCMJJ8U8Z1sT49GdhROR3wYJ5RyfORy5MDCf2CoTAfXX2Ch/m
78fUEH/qENGopHcQarIeMiu785pOXWIvMnq1AjjRjuZQ7SdzbbKyNB8y3wRkKNX1
8xq6tjjAUrvSp/Tgb1ocmQeSiM6Cj7KhWSU3VnN+ysp1vmrl9oWuZHVHgiSOEKZv
8fPE+5DJbx6E0uDTGV1ixJE4TNHJqU1kQMC6Qu2j3xeJiHpaWA79T7MUsX2RB9Vk
CygUGjeG85jHvSBsMpW2O+j5VIzRtcOP3WfQzjPXTzHCuCjvEtu3K5c0MwtPvE/f
joZH8hWv0QXxUgn6J9ZGlPHipDiY8KpWvxg+fXlongemdRXt0Fwzvj+telYUhYs8
pfh2f9g13perCRYcX3jxOu4EUnO67OKLxRvDeqPD4HqhnMHWShtJOX31emnbDpiP
Gh7tw9OLmJCpXE1hCD92qMmXEAin/y5uoyaC6vLFp2HarvI6kP1WbHLxMwLb1i57
Sb95KuRFHWZv0v4h2+tHl16ag84+UoDN2WOrEFMlezWHOC7sm0sKsvqwfWUMeIoF
UJO/+oSe3T1uj+Rsomapde6tBx2WpGqHS60NPUQALx87l5zMWKqrUntLtNFxXPJD
1E5Dz6Y5e08Redta7t3EzDDOKcjbvVoCWFg26LUpoL5W6uuyA4wgr5CJNoEK8gEp
xYAodlVy76QQcNGA2jHiz2Yf+RCqBmp5LbfUj6pbZ7aFA61QPzm8h1Q8jJz5rAW8
i01ODVa4aM4Y63CxSzwvAPtZd4Jc06ND648bKxDoRwHgOaMQfT15m71zh3l5XEAd
gxJUyz4H1I0m5rnxtXbMDDseTgpV1gWEC8zpRfseV0Ki1kSS+/yQcNerXkp/2iwq
TnZbG+7T3Yv55R+gzHde3Ff9kEvAbxyAWqGb4YW//SID8mVZfidjU+2+4WP1J5+A
6EpD8dUmXTsAHvPxufXMnTlQdhgtZ3dWW7Ye2gK0bs0JbHLfHNdc6kXPLTlHvs7K
WxR067f2UfT9B1pEsL6Vvp/dd7pxeJMaqemmOKcV/H89LMrT73kgsY7tFA2u69LV
wRP0r4MJKOWY4l7W1F1+R9OgjEt1vmBVPKDq1OfOT+9xeZlwojyu2HQ5yBSKrLPk
/aeNm1X8nfCv+cs9hx9VX/qHdy2WsXpkRxfCFDby6ET3SvO8DJx9sBclhEERY+FC
0zSDBwj9ojv8LXmxlgbAUy2meZ8CSWSH36Pmxcp6KB06BKHDNXjkNItrq8gLkvoh
1FKfV7+GQpCKzSkQuvidTU/qBdTf382+DNDJJykxKn3+En9oGo4rZE2HJea9GBlc
4smFpyyAEo0eTjCai8BAkJsc+IT9LI/1jh31ZgDec/uJ/WyEd9+4uV2bhKErVs/f
lPLpXuQ79eldTI3djDYUX25WAfOZ7wXyKlPbf+0dv4T6Z2Hizi/iScd7jlBN6dq9
9nvJx7x+cHassXDjVrZKfsIWLJUChFVTM12KvrocvYLpeZM5l+kzc6LP2PHB6S3C
/cqIyPe9tYqRaLUXhkMXzRaES5OWav9Ov+U2msPnubBuBqBo/Dh3q68ScikxfHue
eZKiAT4LJChErPosKXrI2YVxfuTuvecAJMTU7i8iVpusd13GPcKwSj1qjBHafNZV
lY6Vfn0Qb2Xg0JRg2YCx62yqScIDqV/tONGHxtzWu7bU6YjqHaRE4xexo+q+SsMo
dnQFKxgVj1EoHZamHJ7nZ62IJBqFdxhACQ4bROkDvgc+SdRKPsig1i0c0guPa//O
1HuKiQPQ7eFm2j9sDroCck4CC4qlG8giJHh2axV5CcR3E5pIZqm54dHaAg2wQA3L
mRnHWs9FOMVRBgdQMoZLZPGd6qO+PwuZKDEOt2tSGrcd9hlhD8sGKqQrxFQLwPoB
ofccXCkZDS9/hXUS3JUZanCx2E7i/SHthII+ISRtcaTkyglNMJeZ3yYljkCVAXeQ
2tchrlv2mBIcF0nyWsORIddk1BkNbIHtFvDJzo664UJzkLpbHwuKAygdCW23BebT
yBtU+fki8/Xod9qD7P4xf7JdOFR8pK+85u/um/3nylIbfeW8c7wk83NwSNiMRZ9k
QlJngFGYAtQg+R27GcLdt5HUMbHTIgteLTOuNJvHjhOUWwM2wu3ca/vKXrjXKPHA
JZqSIFM3w6wBzOYuL47+FaKd3aqo+dG7ruGfVNgvGcgkoHO5MxYZXWsiYFucm5DI
Y6DBbcyK8EXNdqKE8iDNAOwJxItsGYMtCTIgLtuaZu66Pkd7GyKKLVYD+b5Y/BmW
Xs4a53Fr04xr9bToobqYO+TcJ9nVi5peFwWHGFwQ/c6C0OtiEoIzb/WcMnxWP3tR
zAl8TnszRC0C7Q1Wgan6L7tViXZc6nkIEXNKcE4F9PGyzWRQ+G0ixVvaLNCb2h2F
S+GKAQWZRPgU+HlcS9QcO+DejVdNwE39j8jLJL3UobJSl1MiYTCrjo4CVpYhlZLx
WEaQkBqe/HN+IPR9GcUM4OoHv8/WFB+5aj+QtdiXZVFEshqJ7Efy3cC9ohbBWxy+
UTyfK6ZAFS1H5WMbeIdoHOx+BfvEVVSxEt5Jxv+1NzCdQ69SsiZP0YthGVBmiTMW
3VdFMnYzAobJA2XzNGHq0zacUcHWymsFOLjOqeMOIl82xU4YpNVkOJk5A9SiXCtW
tmbC8Arw+wTeBOwoGEsjMtuZJu/mS60BCFmkKxuSN01vQYE4LZBUdyBlwbHMe3Xt
FUipZGar7vvpKIyeud908eoOZ4dvhPpFjW6Y0oe5vujyHPsRYivIQ746OkNOkMMi
xruf51cVo6voHsk80wUBssp0H5QlYxmNQ9k7HjHomo/wSqm19G5lFCTasoz/iOs0
I7yzlifig1eB59kq/7J14TZ2BxrBgxFLgLn7ipjV8/CK5Haa4Q+iV23EnjFxuLBf
2ap3N9bIH4C4y3Lwv0D+cBlJEr2O8mxrIU/01lZ/Wk99dEZkDGrK+J/7jfSgpXMH
jRRS/LBhEPvxXqTajdu6z45m6nSMy7MyKfXGHDpKgAudB2NnrldKbKypsIt8ORsD
qmIV0frACJ6QIaEusSqYkwyvB6LKZpa2io5aEFP2DK7ivmq5957oJ5v8EqlPhr0q
U7C+C1urg4djXguWUp8B18tKDNylJDBW0vJB5e2ULsQjygSW+NbSNQDxDyNP6PoX
YGG3FWM1kDQuHlc6PpkKfq23zGW2KsGeTOl3fzzJNwfIc7dzF6jQ9K3ik6L6D3bN
BequUgk7pzCcm7RDkl3PLWXawUyHIqxRiXW3rttKEYGk627roLKIs7Nc4yNuZF2c
CohXvlmjx6d3639ap5s94ornbied8lnBCXPRNssWeWM5j29l20B5BsCN8TLW8q/M
01BnNhNNtLlNhqYOq4uDCqE3wE46cdY5dlw5HzoE9Fm9dxyEnAvxKTHBSs3D69ww
RqSJmwaGXEcG0yuPA+A5oyhBv/QVk/+cGaelyQlNaKoGP4/aSOz4O7luqfV/r4NH
vY8TTaij5CO/x1M5QAvOtGKi8eGlH/5A3UvoSzuoCgf+uFistTFs6qWz7TEh9NzC
WKH0rZ6QVK3GWH6+dSWUmKnRaeF5KkEdZYoBRoF4P3MOgPMOxr+LErpa3Rkz2IML
wwO4FO4motLKcKXFAlUsPRgBMPsQ8OFn/P5n3AJ8Hjl8DHOGiCxgoyl65HyMIzwJ
ODjTAcWSP1qPlsJmMD05/gfnbQ2qwQQeeQyhYK3/l8YajvK4NNYh7aAXSzsHCI5h
WFI6IzBmuIgFfP4dRpl2IaU2uni62tQGP+m86soUSjBwEZlOdrWkkJr4xz69WYlN
LA+5nuXLS6zn6ckf6RLLfoOuUv/Psm37dffjLst5JjB350KrNhzL8Pgxzrcd1lkM
8DRFzyvA4WEwjzfmbPRAnfMOtmgfNmzsQqdKY/j5+r1OuqP3JQiHqs2nJxBY5yGh
CMIE+EPoN1JFTKBsliIYqDkq83O/AVNoVSLZrkxcrs/jiR7oHGgVMGLKEUataUZt
1eD0FH+m89IfEqBVnk8QzecbxTcx8I5BxkTzq414QkEaLF1HeA9Nc2vSRyeIhTNM
Vw6+LUo9kps1hyAbFH/zjW/VdwccthRtlyri7mfZf+R0mLEgnxCQic7NSAlI0ol5
YbO5ZdRWCTnS3t7S9Z3eQRmzBJyGq6sy+5fS0Boazaa+DqrNzqZ4LGbV+n5WaMSo
p2LnxNyliH/SiixTpgOCRu2aX8oppSzhw7KLzLdHmFlavdqZfBGJICjkdQROtCex
OMVF+w+uIA2RCAHzLdpjMU2pHZsqD39igvWr4TjrMUL59SRJKQSe675g9PAD9G8f
8MBigaZb6cmILqfEf6rwuRjfrUg7/xn4jkvH5M/tno8wDFzEooxP9OpWnUCCvYPC
t7f/SaWuGybUHvD4j2vXUW5UHcst+5uvGzJvvWOJxe/fdvHIZ2FWfBLYPCmn44Tr
zxmUwGY4Byw00TwIc8xKhzfhCCpcQsarvWfVC+jIMgrdZL8Wf+/l5e52wpQYsP24
zyOikfWyVo8hD2sc2A0zM4ZW+zDmygaw1Z1Vx8xB+6CPucMUwRhgV5b+lKb2Ym85
3Ss1ogD6G+NYOnFWXFZxKGNx5AdTkmeTV0FLnFXrPBelAdSNTqJiohdK9CIGRrcr
g9Dx/658WCGYLsKppubRSZge8vG6IGzMpGmRKQl4kNruXn6qjt0Tn1gqIpr9m0/y
mBEMBxsbpGaTowV1vULZ5SgNjYaNUF0XQS2HgWcUmgCyxDIz9R+2VyUf7O2kH97G
SkOGSY4JMNt2PpHyivLlsCM0DD0eGiSGe/6MYp1VMxj20kQriyQpqhDzol5FlMWI
dWd5DWy/s9An2KVxD/rco6QRsdZzNGi8nZyeoPfaS7fg5GgrUtEJBMWQFcNv1c5A
esmKpvEjJ4FdiUwM6/NeG27ka0IHciv7MTOgqwR/LM8HIoE6wjOgmxmayKIjxb8t
zQVzRQEhxhFgMNwyE6agk0sKLfxj0Hcyz48MVaVD72o9DgZU1VndVBzF73O7m/8z
OvZWXaH9nnbUHXXw79gmfVfKT7ZMp2QzbDnBQe0qZgjYKNhRbbpme9IWhs5+JDjc
xjLnU7B3V2S+HdLEOhmzTzEzSL9NwQq9W3rchrtDU/ZTLC5Pv2JKefAB4jBJxGcC
peXU6ChsMqFD3F5ixw9ozhLDD/VCWchzQBIjte8IwQcQcPhRrWAfRCSkYaa/N0dJ
r/tYVzqn19OT2dUuZ3ptpuqaREDMRoxrmO6cXd8CkLpLGhW1TRDopsL8N7pVVEz4
yKxETNqNsFh4WR+ahWcaJSnS68esukq0OVCIaQ0tjxaJZVjPg5e0OMgMwxTIHUHY
CosUAsq9LYZ+QRzIO4WChsvIxzWY6i1N2FE4WrzoFIUQaXf5nWMnNBxm5aqU1z58
EwOm3ClNOk+oAaowtI2G6J/BGFxloPe6FLwFO//+TuTNUZvotZ8mrWtAphefFHVR
wRABz3s+lIE76HRPM4DZEIWKMgjoKTn5gSR0NkLFmxOOuI32NBWRZkQVTz/iBwad
qABzH4P+0D1p89INZZKD8yEZZrvdGwCcZbVizBq2Zw04u/ApKGFpYQWThYzCzXLy
4B0/M13thlHJz5/f/0OVdDjtSQA82yJ4fa9u1UJFp1m1w9kqEUnciHQbE/xN2R4C
Vz9czrs4Ug2zv+yR2g6BHPC7FSOXry0gFY0qFF2J0LBweveNkZ2nOyHsP+UOAeBb
qgBz9buqhdg1ss1407dt7ztdXx5YNsldlF1CsTZz2Q2vKZ+D8bqxcuQePCH7d5Sb
yF1DUzDxqWRNR19PW+1PgHd7NnQJns6OVyxiR69Yvy+oA+vFcp58YERcps0gjtOC
fFC7gL3tZSLytR91f2n5enIbUh5k0upRzcyyJlJkw5Gb3OpY/QqRptsqOxADe1gE
DZNAqDL3oIa78JuPKqZ+KGFRMA3DgANzU3aqKf6HdZe46v87b6kug1S2Wpwr1DY3
grYAf7Ht9pk+EBXexlcv9h5CsK2n+xui+oz7e+qzAA6ZvfkjWHQhQyjPpZF35wlq
WfLtIebJjCSzQBNDHTH0jEH9Xtb/Ko6J2ApmmGr20xcsrqhD1rVhn/O0Rim8FdO6
o4F8oIgBtpWMT20tTRoo82DbL3ETzMOsg5hfxj+Ops9JrO9KotApeiUMQJpAaDpt
AGObSantD4mrc8+xsfJzOuDJz48EAFt7dtBMJhy/MPxmOzhEIRuWalOvKx33ybS9
zHl2Gei6LjinYoL/8phkFQ/NFaVFflr3UpLHAouCO0AOuIP9dwiM1m/AlNZq6tb5
0AvDWFwkDm2u/2XQ1rFOxWoTnznEkE0psGNfVv/JXRt8P14P+RZIq1yIXwi1/74p
TfneAQg7LBZ75gosGcYCcLla+y5IpIgkJw26b621WQ5YhjR/Ot59Af7V7MoInETq
QsEHit3sdgxsR1p38t+ioJQjliMObjbda9LkKv6eJG8D04oPiPdzgLEPrQrWdA9W
7a5GY60Y/qjZKh2q7yWBUDBVrOVh+2mkYYYmq4dr+ZBsloP+0bAeJnA0sa9/h+11
oEDu8e3ZV3GNNw2/2TwTNInI8R45kF8gVO2kAV2BSxUr8VTGSK9hnKOE7S+XcKXX
7I43+xwYUkvv8Kk+osbLoYH7JOeBKJdi+AwRCeXK4chie0NtkE1f/vsENcO2H4Ve
dAEbzWChEbfX9e9B6KozuE3z1GG+P/T0BcXupzoLmLcNL8KN9CI4XS7imdGT50vv
dy3hxjgiIVTPQpaDej+abUGurH852R23szidQhqrzV2IVtoZ7z8ex2YJX/3yW3Ud
Qg54WNAAVG2OJWTsnHKMFN8DPreWNvUOKexAhBTm9CbFElX6wi6Nu6jZLZ3YVi7H
fAa+W7WFAsBw/HYhUAFpMblLU3PLw3o7vHv0dE9Cfb46PI2/gpfVkaFJs6BgGC3E
RhT6Vu7wC+gh3MD2zTTmnaXuC7DNZjZFXLcBTYbm6Xu7gMtw4OjFWBL4znyb/+qZ
OLrrEGUtU/J73KoyKDKpZnaio+TcYw+96jx5Qp3mU+pDpIz0Kp9nS06H9yUHK5yA
d015KWUY/SfadrK45n6JsuJM87yHtFfKQmMfYqAZtHLtWjiAUYRtZCcNtY9a7xZo
tXMeBSN89VFNVr8sCr71sEVmrx8XERBFPkKptyTOUbslRzwGsOsJJGViwd4i4DKB
VODWSDS2GLi7pt8cCKdOwp8JYjYgbXPOMW8cKEOBk5TCh9+3U5p5GAYJhagG2hon
A1kOtpNa+YSeIXcG+4eyvwubLfZM/9n1M64Yf5m3jK9x7CvctE7Bvimnr5DiEwQe
pVIOtXQ0x84GOcYnoQtSeK9HjuRzgzNLy87eVjlCBr5wg9W95XR6FsaHZpHu2OoX
Di9Npv/nBe8ZrPf4jvT4SpDewQyiV3/N8xgTekwO0WO5CADaw7eRSOUKvQAfWYNz
NR9YroA+TPVTX/ZpLHZEaQIHcZ9LxQ3BIfKhR8W1Pl1jAYMDYQLKVy7xUIaIDJOk
UHo8TZuDU/fanKBJwCS+ZNGQCBuDMvVafU95jabKFXeKVe6jdy3IdG5z++gbswOb
nG3+4mOp2iBZ6slIkrJh7I02E1QNwnqqdzyGshgiLXyF67NcyIRvSfB1gAjB63yG
ALJ+Wnd/ZttFrtrcodpvB+jpFxmLdRPwq5Q2DNrbsl/eXb06Y0XhyqspL8UKnbKC
Gy8wg6FhBFBqUwcjfSIzQpF6vq16o7zJ6QzYVH/ZZ7vZZ7cL2Y0f38Ok+ehjCGmn
k+74pWBp8iWv37rccSo0j/1yF3x9ivzgEfi6A6yhjG31p/+w5/xtn5Kx/G8ekolb
FBGSDnZuKf7W/TiNFvpWrC1uPSUiI9gbH8DRfgUFSPF+xJe1weiuZuTE/FVmvHtX
b2KPbTnNn3ccuG2urzl8Qj8ByZiLH43Li+kcrzPi4dt/q86HT0dZHihSnIjawiDw
NbReGnv6KSvdkmL4npdRs4gUglHvvyW4SbV4jKMDnpKYUAMqBbJHAj/yST4PfP46
YV2mo9CxsinWDfqe068sreTfC7YA4oCkv7xf9PgyJcqlGwhYjY12mCQyPSHbAtDk
8/AuEzcTIzxmzOI1auUEiIgkQg2dSyHpLgq8F7XQtfGK/rWX08nKgZDsHWkwcRz1
VRqcquJ1jcpycfJSKZwFJYU259iZaoOZe3+zghdoMnTVzTbLHC2w+6YNCgfeMBM8
mV64x8QR4dGm8g92YoqmTqKXR4/oUCzuwx1j7HbHgKPluxtRtLLFe7qBkflt4d8m
fKzQTxVq+6upI5LogotQttWWX9TsYDC6j84rviDkz/1nuC/XEm7Cr3zpWVCGdzIS
CI7FbKW7Ukc6hwrjOzIds1XGMvvSYGfwgmf0257Zw66FcJZfC2jQbMvhkxIdjZBs
qQ9CgD+Lf/AwtChlhuD+Xu3I2CgQPlX6x3T8XUkjxczprEdDeaGp1UyPEbuVvITg
mr8GFOZdIOgCY6TlLLd99mhCnyjTs9KXFex3Sr8A6SnHyVouWEMgPhiFaEoKsAp1
nvcnKidBGSx2wNQvqmqUkZc3jkCdCvvHBipItlRFJj9DivvY0UGv6douyQG/xwV+
7DslW7cVNj+Ad9x97vQ+BluVTXGIeSDmzt71wfiWJA5rScL1TC8hTGgYo9fJUAo4
XRrPbQRlc9Kjq4kbfV1ojhoHBkFexBeGglWXhvetjvkeda32tkG8ypO6xD59229g
b+Qjk/tKqfBUVgXDu5jPq3hr/bBqXm4JqniNfCnyv8rmkLGYi5y/00sssuppj31t
IsvlMjS7qJD646dZnXDFLMc2PnTloW3JRHPMw56sqEHqAU+cuxHW98JWncrtJpys
hd9GdTNtUDRqW9xfIeLK1njwALSO+lDNs3WZsDs310CpGUxFJNDzPFe+4twZ//gA
fBRLTjS3/mQFUYMUMPPkeGrf9IxmIyfK5USDyMVjPD+64oAVBRaKQUtxeLQZ7+Co
tDzKLWWQung9oetTIx9z4Kr7JDjFUY2+vgljUjcjnQPNdptkzlc3/OTMIfiKfEy+
Wo5p1HDlphzDJomiNrGtl5w5YTfsbJVrSKAviijWn4SnlWkhTWHwzabhOnVky/7k
cVDLZ/6OgqeRIEqGPXzoOWlOK2eP9wtFlz02UviAj+ZxF+3nqRDYgwZ/lKGqdHEm
An5L8emO5p9Mtmz2k/His2YRwIGwoHPaSu1cZqnJXgb+kVUlFpoikW8Xq+ADpxdF
JgOEd9saATrr5WGeJp7NTA+F7TAre3CxrQYIXUlMzBL7fPFXqcZzdXB+FlOvRps7
cGz4Yi97vU28BSjD6AoyAiJgbO5S3mCaKOtBqrZwWDszedv42O37fzKuv8v7ExN4
GRDWdrLqEklf8Usbyo84tTNoKq/vGYFTR3qisY1/ktor0QgPZAzjLexpVaK8h99j
MfXodfasJ6NVD+6sDA1cSOkorlD3Mw6fJNx1svIYWn/rSlQKNSfifyxFxReEjTQ4
ON4l052Aqf0pVVMeTIrtEHlz+6xWsNUzgEFDqfpVMHehMopp/RoWjATJ3CImY7Yr
GlzwLq3L2eWhiiPQFTRSIkp+8KVP2E7Rx3SpJxSuIlK3vCTDmdSiCya80v8lcAgO
nsg7qqg1ejCZ3YASLwzeyyJWhqbgSI0wk7i9j7R6pbaw/aKtgCL7EdTrm3AJPe9k
NtcRU05Xl32l6HX9gFenEIloagipulYN1WvoMrpWNU2TmwqdiRmOYyDtmJoqs2Y8
pEd8dH5rtvifDAILYosQi44xMbs46x9o1Yb4XkwYXeewxnbzvFvnuu4GFZSqdAhS
fArzcFFmj+2WogBlZgh/lXr1Zot3kpz1yElx77b3bjl4cvxnl15Rgc7vouYL1wyb
WJrgUScmKp5WBfKZhRhqCCqe6+R+34Jpd7tFhek3Bty7sFoMnQHH6g6wMnUQrNDb
a/8bAqpvGuN6ITExNV/PUMrw0F1fw5eg46+WbB7ZCKN5OVmB4SjgNWZC50KvYM6B
5Jc4cSEDNx9J1MOyuYbvlvH5j4cnTnptFdXD2Mq8TeDpm0/CJlc53EJocwAo2SIP
wTQ71iCqw3t7tCkY3ZBS4SdWLsDOMcZZSyk4VCykTQj/HCDZDLWod2mTs1UjSF6t
naExWy+vntsYdZFwiojfFPONiZF4+l0m4u6TOMLxsktK4xPBo9UPOD9QwtpDHRKJ
UneNUinrJpyVXCxixh4Xt1uccG6SCJPmyalfvvaJNfs7iTtCzSqMhqpicCW66q2w
qCcYmoXtkHnnmk0aKixWvBTqpBKjgXi5UnE0ahF+nlVM7aiUnArPcrbJWC0FHYeb
U5j4tWefZmSj4sKLnAspiTV8rKraG4qjWefqNN/Mu/tAIuH/YxHu8KcGKdpH9Hgf
tEcPJ4MzxmEgTJPh2zoAjYsqUqaQOzFfOuaRBzyGvGgqje8R/IuijhkZ3HG6h6Ba
nXu0vRUPZuegF8AKPwO6anWlivDIH2wMfgZDZrA0hHD4LyUfX3NvPrZVI3VXR0t6
gC7QDBBqtKnljv7qEb9TLbBbNQduaCxDSAHxfshOUZ9A8gTbcwJP1lr5Jg6XDwfn
nURmvtnaWb+loB3I8nfLWvRelTEJRRswrxmAFSddqYKiVm1+zGTA82Zfy2Ls7yhT
EzeX7cj5FEGNMbzvbs/Fa1LDm6q384RgO6cniRC7y7PSI3H2uSQq0skoDSLV3FEN
MgVR0cO7hotQ/KmFf0p4R6Yqv8XYeKgi7gJxMzkh6naPF5OwDUZhvxSWtfXk2ZXv
KfaT+npVUlWO/BWDROPDvdtb3wSYMVjPptix6xgJknVZ03b+3fAzrcJk2nNRDDdg
Ww/2vo5wUcPXZag8aBKrOWqAh/xiUatJN1CtxDcnVKEJbiU83patWbZ6pqMF5XD0
drgMdYWEU2lgsrsXZa7lM2dHH4psNID/0uZjnLzlavThh9HNwQFBn/4iyZA2uKQD
o3C5I0lVts7UWhmwXB0Uiw4vzcd1fhtI5QYTskSKoQk6jIBGAClVOD74/rKlU4n1
zThcuir71Zf0sX2jL8QB60VcvKn88YuoBV+i/TmOONwpovu6Q13kTynVjRm/wUVB
nUdKDZWyICu8eHcX+ba856oZOTrxTmmwHpW1BJ1zJ/t2D9jDuIoz46qjvbuXtzRz
azdDQ/oGK3o0+uXdWVUaDwIX6Js5rOiRKR8o9LcDGyxRiTbMKze7W6ekBUCG45U8
TRM6Vd5dv/a1Rmxuw7v8EMyYf+EyhBpdCjCyERpXW+mMe3yI6ibAmyPluRdXY1N7
wnrjw47D2+gmOpclLpzLYFmGzvWf6TdOlTWit0mAb7BoKInT9PE9fzSuUyxwIq1L
vGWa5IZ79V5hNb7Al5/iOg5JExgGjgQeP7W5ynXmLvmuhQ69fMNaH/7nfPegwsaV
D661DbysgbmwpUBBEOH65H7V1ptNKsDAbWaYztwksVAOmI3XwvVxLFgf4Xs42jKq
+HqshSGhgRnw+LUsl4PFQROR3Fpgqkyxz7KfazO73ZVBE9l2HUcim7Vwo8lJfRIn
cyDQTi7oJUHlBOQ4ltguJgNT4ICsiu4zORLEaIEA0oxbQvTXXcuj04X86AbZKRf5
m4DALo/USszJAXp0wBcGSzhlmI9m9BEXZ+8cjjkOP0gpn/J4B4ZXYQo3DHFvMsud
BRww/TSusiM/9V0I6Oy0qKRgmu8wSuWIdViVuHXhW+PRu1yA40pDm8QRkFrC0+Ia
fjMDuBveyL0Gnh9D0EyCA01ThrFxkhOrM2GFNnIL1e/rhy9P9vljQ4vJoE4qEwQQ
J3P/bgSAHeulwQgl1T3NN+uEJHI2qNCkHgmudxGoPjNMjz29mk3sfovSggpBNcuV
tR7hB69MbhcF0xILbwVnJ1SRFoTvvDs+OH2V7KnJ8A0UNsGZGZC91PhSUuiS4gGx
qMS6wsNmThsrnFelVqEvHgTrs3ubCns5mROL4Pk4q63ulyKIk8yL7IimOp8wx5RW
gQxLknlme58fm8mbrhqb2ZZ2hk5rlYOCsztANxA8Q9kCbyDEOhZ/Nl4yqhOwKrHB
yNyo4fwXf5MKqacaz49jzqp37SOk0JdOMsYnha+zV1/c6uVJBwijn4l9+qk5zQKe
DJxfncnRKH8YEAeSFS8ZM1Zxnmw0KbH3uAU+ouHasrjiVINSgWJFg7Z2su92oSI1
zh/E5pSaBHXPbGaZa9+pBm/e/rNeO0lVPrSh7bEJxyaLmyofQBT0hSDsWX8QlMu4
jOqitbMoHLFS48Sk9fcPyXar8SJl6p/41EsV9iE0ifau7ZtcKrkAd/S13WcJsGpu
hrzD+V0M3lE7gkpDGBv27UV8pax6+ufpDdHQC1Wi7JIMzXIMH6Y/fkZsRaxA7jPK
oSISFIt6ZoY1lurG8Dk+J8ofjWC5ttS4QFhoZzcqO6wdV/xdYFLU0ruShlD69gsU
+mGUqVdL0QJh3gYeWn2BdvCkwp010CaJggG3XSw8dSn5Xdw1GuP5Fp4oNLmH695y
C8WWFETSSPlPZg5AmpOaJP7DND6eFqUO4Vfc72nPxKvbQIV8WsBvFWCTd2CRoiYz
YhXJkXuGC0BvKrl8AlVLIGjsAIlaKgsnyt509miL2eFM8n/i85k0AxFRxH/gdAS5
6nyHVE5+Ak49DJrqfI9DHf6RNvPBjeIzrueyaPFoK93DIHOvh+nLEwOMaQZTDSiR
aMAr623hrdtf7pTd30VNu8fA9mxgEQbWfu+BjpBgbTkE/mZJvq1QY3dK7M4aVq1H
4upmEFvQYOM9xXIv3wFN7CqYzOMZEvHsiAEMk8S44hZDIBmUBYZPqDmfASorWpCB
at20jLouLeRo/h1J5ajDsfjrqmAwTmYjKr/j9vSWZ8swXrGTzCKn71CCJy8r9/x/
sgkNJthhi2rbIdg0aQ/4TOArTHKKo2vK7pk3KvbBST2zJzEhLX8xjK6REsd9/07r
oNU5kyumE1cYlvAiXe868EbhSeK1Juy1bfzIiI9VSz7RD7/GCz/vINdY7jlmUMpo
K067IsbWKST37iUpN2pbdt6MCIKZ721XIWpwtmfxYiGjeYyVWAN2TIgN0G3plyVd
eRqpfgGH0kDueVIV180mNLA91CvWqrCmiFlT2xJ7NBPHTffztIHNkjeCJ8hQcVe0
cr5JV+0FwwxYfS/jDSe5Q21R3VMyh1lnjAFJTqEhECgG+d8WQ+k+lv+gFe+AzJIM
ijAw/eZO+fKyl83solK3mNLrxn+41XOXsumjiVUO0lTt5F2sdGtXfnxjb8uI0MiR
B+s5lS72zHiJYV4to6um1UEp1gg3ds/3tbVaroDm7VfqGa3+5VwHU5uvWyvrf/ga
WBa4O7e08hqi0OB9WnMzFZ8Mig858/wAZh7VqfFBrVuYQ6XY/86hTEFw0HkSpqnF
qayS4AlYU3ggYhHDNxC2yrXqwGTVNjpTmactzmad1JS6PQx0iUp+D9ytaMBAsM7q
gfKYYAXVrH0uDTj14cPLmhu+3vkiUrwWC2gvIkEeHK4hKHvjc9Y85RVuVM9zITAR
zNP8i2+TUkW6BUNfn2vrElfpKysdSMScc3WOnE0AdNxbnsxZhrcco1iRKqoSTlSK
/VjgZpZIJqyXu5/51NAkke06WS1EqpKAs9KeheGY8ENnR1lmwglwbfeDKOcyItuY
nn2ldYBQj1Vx9dbuEz1AmsgzsGvH18gZO9OG2lmUgEszaYACPLZwRYqORYVNLd30
odNSldXJqnmjSLeklORR2MhVQGFjaaj3ZZq40oGepbUoJDoRuyg2zMOqkr2pz5gw
R0p/I0QljJwLZYSEz+bGaRnzgEnQANhw16czMwz6/qOY6AIPT3gy7tcqLupyJ3UR
f0ZkP+wa3ozDv1gGbUlwc7Im56PBEv2c9gYdkhf87DD13RHTzy4sJJR7f2DN51pv
xlPIXzZ1EfFJVydy9Hi6uMmmOTm9trRGVlh4OHOt/kTmiClnH/uzVteWstRmaazL
Sn5fdBiZ3gFSF8bkCXX8xSrCcJEon7X6gvglpJ9tzzi+UINqrxcKl2/8zNn+j6AQ
yEpP/KaLQW3daDO8Iy6y41PJlk7oafM0uHpzo+j841YSfdfdienb+29S6lNZjMSI
aM5EEG+873DBDDCDQALMd4X7cUkUU2uzhSANjzZOkoUxTmNQDksGkgKxktLf1Izg
3WVp3XHad+OCrm4ZPYLPbNJFxfuHcqwNhn0T9DYlQ3yLWWLAENk5gjMP2OyfTR+u
a/7XzUTzq4h3W9sjlRuoO52sW+EjQyJJOk6deUhJ8npUMplktJeOqGZtJR2+uyDT
UmezxBfzDJIdS2EKJRAGFw+0qIOAFRbse54HKeJhaq4lre93obLHSoUgeR/Rvkz6
iSxcqzg84FKQElCzGLfb4n4wFZ1pyUi47fnWvI4tpO0TK6aq5XUWspjqa8w86ZHn
2gPCZYcy/diVyXydJws92jLrN/9nuE1ZiaoyouV67ZWooAz9wJCt6PMm1vR14E2M
jOw8O+51VQgarLD617OhPMBjGYz61+tI7SUW0W1yPHAkuq0H039Y5IK4y52ZoRBO
uvbET5t6VXrQ1+DCyeOwB3fXCS/PuGUVw6t783l2ynmxOUF9e4UgZ70CtXjNQj7s
bhhbsP4G2qXXJII5mdVykZYTBdBUeWQQ+y5shXHpoLrLQTa71EYQMSf2T7Kk1bx4
SqKtbF/y3ZP+9BTEukU1R5QfBfMgVzly5xnhBDetjp4fYEgit71ZPsZnKMcZ/7LL
1ju6qGfpoAfK+1q0QXGvgGa7ggQWF9H4FDDVnkFjisxybXw5ZQseknjUTclWIG+h
q9lQIcUIgKmm6+/rITRptdZrd9f6z9tBg1brTNn9VOCsD4IBbkgh4UPc7DCd7bqM
iZcfMjjz0rLfjN7+sIpo73r/OJB2hyEkPWwFa2y5S7ilWcKBfD/vx3WoJxWfjlc2
3++qE+A8omnh/ZgxLp5ItkkBhNuCXzPNuDYOpIlARu9TiFGZk7TrTEWIavo26+Jr
BXBSxjzya8HEhd7qi11kJ8Affxjv4Xw2LEKCeQ/lavnPX6FxkYXjrQK3vytJ6LYl
dYM4qdHJygKJc4weZnQNB/6jsSdouqmnQC+8T2VQCTw2NnDcFxC80DEDH+yDxz5u
Etdl70PFPQSGArIWOkPHjJoVRAa7376JQbMVH2zjXxv2d+TFo0HzztsvM7daIL1R
HufKq5Z183ZP+LJuCXiSHUlb/EeKjjDku1SjS6vfrvxfQi3ebLwwUeLS1X/aI9ig
Wf+ihuYSU6qZRSLuvkazVj0OnETD1OewIJDI56dwblkH3ENBZKLxd5+si468qTQY
Y6SHZhRyKbPyPvBESCyXJ0CllstjWGL2DsNUfquxKhiPwDTiade8e2ba7gpq8RMt
drpV6u98N9WXB7lV3WtW6uEgViW1A/dWFbtoXzwmXUybm4+nDPjfMYHcenOnP5Z4
wyLDWUw4Uw9r7e217kuaTN/ZrUdjnX2xqgrpG1V74PHwj74/TkgE978aBG2ptZSC
4beXCC22enFABxAwY9zQFHH9aYYkGtNyNmtoJHfzi4Oi7xKamTD90dGNzdyShDtM
Vq34+7SnWsoIpnWockOEW2ECv7PQVHfAJsVbTID1abzSOVjZ0434xNYUZOMVIvAV
mc6z/9NBHjaTRWINjGT54fE97aEGtbLw+x89vcDgelw0Jc7hUUYlNvuGO0HMaDG5
Xo/CNH0XzMcvsDpsy9iOGECaHmXIGoEyhNE4KUafyj41q2TL5/6gi6vlUbgSdLex
HMSSCSun0Bz8ebF84EpjrAzj9qkAxjU0n52+VwAglFCSy3+GSnRTcF036UM9H9CW
jv/wGktk1Yfa1NJtIgfNIWcMeMjGXtDhsTpgPCP0bYOSDJVI18c/H1+X3AMbUmh/
zNB30V/oLxjoEFG80JBmLfl9uR8A27Q81/XfJGp3MbfVQan/RlDVCRGH/mJXMF63
gCt1nOoRgknc4WbD66YQuhK5vq/g7XLMS2XYGZEgam6GhEIvnKrLoQuL6ueBfukg
EGFZ9M4A17BhmaE3OBe0fM5uhByOE5lg4xsa93w9jvWeiVNTaH4oeoFER9aIo7zl
d3+nV5SgeUfMbhZtlbRCL7fhqgiiduAT2MwH21uRXkMW1lpND9cTmCJwJcMfgJI6
ROC6/Tmgkrt1tGb+5/UJtPMZ6X3hvNr7COnzLe+Tu5ND3kKTL5mdCrVV/ccRoEEE
rvEWTdWJIu1dRVSRjUH/BP88NT8+OTaCfUy51VPe3w4Ef5O0BgKEeRFqRaoMXcaC
FO0g3cpW1sLmab7JjoNZXOwlEbe07f5cI+Ge7ehq1q/oE43/hhoezfjPOZNZITFi
Ww0bv32UbRQI5o4K2zCAzugTz0uFUCZAqNfnS+g4zaLC2cOhpKEv1gZnJAglAebs
NSe9l8nM4B15I9ry4Yi5lW0Hy2Ao/biqrqmkLlcoYufEGvkz7CBUxw4m88vn6QGu
o1zT8DAuzhzEwBJrypG5U76Dc84e5tS5ZQE+oF9YlStdvE6GaheoftFufEHwfA9e
JqyejZO9p5vN20M6dGIlp+N7juGmpayLmWTdhdrJ3k9C88iM7f5ApwTzWp6Q+rzl
tUnmZgjjFgTlQn/Ta+Rc9Muijl93UynNa9571LjxAh93deuW20+Itw/2rPOQp74L
NqDmCLHr1ldv2dMGbyu9BDiMlrOk+fFmC4wwftzoLQzQz83bnXky4g4H3xwc5Yvx
r6RWWX0sxDw0whSkCWJtPZS6gBS5XTMNQfT+7vFELXU8B6syVYm7s0IgDrqxe8WI
tFSbALu9x0NVt4ST7/g8kYVBuiKkctaBfn45mGnWWl9hb/Awyx1xNRAA4WRVTyd8
TkeeSXn2rMuwKx2dnEVVh14g0A4zoz4siMK7vHw7XziNPfAxQ/Pn1NzhoMldNTXU
kV2eCjQW1GU6xKdyVg6nF8+fYY5+vo8A4R4YvRpFdiUiEAMYeT5nM/VV7LXO4Gj4
KqUbcqJDlA6YuCzuK2f+rWmx2MUba83qNoD1jhuBzSHPR9LzjcglQzDlf1fgVVcR
7Q1mQ2nfP6mY8uCmId74cTDLvSA0iqbbvi+OScDRgYzKp+FAx+FYXDN5FMqfzu/C
HSr6XUjh/ZhutoI9ait0SNN6KXgvCiLiSscsCcQRL+jtJ0SZlo5XwghtSDEaaQpV
5Z3Jm3/X1WdvGBYA0bcTdhgqLph51KtXD2cstUHNBr4fZTT2N0XPjZMXfeUDraxr
ZBh1d6zv5PkQwT8V1Q4lNRQGkomBRXw3qKwvlq8KFcW7GnA2Emcz84SLPzLOs7dB
Lg4AQy+VGDVm6upXiQ4odZLHlcEmShUHN9HXIvTTbxYrbQd6zEcQfjZE8CTHOPW0
T1dvazcWC62T46A2W8yFnP65576LHyrI0bZTdve+RehlWJLipY+0aT4x/9GKYb69
bpafBWC5C5my8qa22QEta6QLeOB2fFGpmwaS7QoNhUOKiBZ4nPU/sb42p96cvUGR
4hbNZoivW2zlC2a6CHpd0NKMKnHQr21rSiewCfnpM4Ngx+uOU0ivMP3j0zfADsca
Cq9G2Dz2/hg5izhD08AGPM05jK5Bip9rQKcHTylKc9riZ2wGM49uQRfQWYFCiBio
BdR5t94cfDMTgS90E6Dmvwom812L7u2hqmTeBVj1u+1HR77msn/Qdw/UQisZUWfq
0/C2butFGSqRNI26AmVT/800QvacBIZoPuo6a5kLwYTNVCT4UJagRentNNKjL4Fk
/Q04SBb4TQduS5ygsyTHr176cfbtIP6kwwBECY/Y27hlCH1669G9ll7WOWXe/3ky
CWXPGCGa3f7h85znZvWpneR4/sMAGUBsWNf2mszy7QDikjGV565/VDxhXR6LDfxp
7SHnjFHn5u5L0PjnbC2uq1PDg7bqL6OrCQKjHEPKDOJp+w7XqB6qeFfjiUXPqqPE
OiXPpHVOV0LKbl3+znd20hteHlMvuE41cl9GqlgZSvRKwJpedhyjYnYZ16zRlsQg
Ph+7AY6FW8CWsp7kVysQ6xTtNjCXt7t/nVa1z+NmAkETUKnC3uHYK+HWRZVfOcRw
bKlSr1jsNZ4O91xSZK+REYsiBWgVL22ooex+qDbCDECDRpbhWqWMKqGpPMXOcSnc
iD/etB5EDbkNuwE6Mbnvgs0jTqhjjuprLh1ncjX7FficdeU7cQYvDKmv7PGao83W
H+JtlABRgiz84WPX3u810OSssJc0PjKEIODsSFD7C2kJFfTjuM+Iw6KQCIXdUqG0
qI8ykNJ4Db2wgfy3QzY4TW8VKTmTGVlGP1ObatfvgzPW8gQRKhY/VjFb0j5oM+Dr
7wufxz8gxU3l/qAbWnqsd2skJibu1qjOAL++ISljRa015ZoVwG0cWO1G4Nh9RLEv
QIVqMZ3UvpTeCeLJYhOGSsadRQyhzNLfSBRZG9TFlK5NHqxS+p7RHt+W8f9WbGsw
096J73KybJXFwzKe3lPY7sxoztRDeJF5DqRqJ5zUs6A/d81u1tAMfNOussZ0AGI+
mzUvVGXgKFeZSiHQilbcUIoPW/2I5tEhxuUrP8Em5bmoDAErfrWGGg5sqpHiXH+9
sRIQZwNDJGvw7zQQuXDfdNDLpFiV3H0rjCk5cjXPrRXhbR4TcmKK+gEXOBw3K+mX
YPa5T+drCuTqXHbxZlr+4zlhEDtfIlKhT2n0swqUItxKcenQkwdrgxXbWDMwo0S8
JUao4Su8OyKFCe6qkBbeMCzntZ46wQF7rHUwisdcNDK8LHsBx85r8PzMIF6w5vrt
CdH70BApZaCpy6MDa9T7dcN9qPcUXsgfK1fMY+t+mcrYa8ssAvt+wPiIN7pg2GDn
MVAilIXHvn9KAloLenTAIJKvbwD3GiKHCZLzZIuraODjJ9Jd8BLyUycEHRtvcTLA
0DBhIT9t/hPZviaH+erA5344+s/2mHAjgglenJVt8Dg58JpFPenu9T3ziUhI2363
fkqzzR9kJ5gQ+HQIu0j/bGUA3q6t+EAmv2iuQdgiJ00/47Lct6ZzVcS7Rs3avEod
xjkZXzLcDaATqEaAoVaWhIvmAk1OC/evjcEeTr2SH5QIZBcEmcn3Siq4y4Xmzhf2
Kz2JivdYV/kiplm4ddj2iOBmTI86cUjEqUI0PgbaNreYtRcmU6WhN9kPkX51o8d3
EXyWoIxX/K+eDsB8UbXAC9z+lBpUbvFiXBt8R0+UVHNRW4QSYD6FSbYG6789E+LS
k2v2EigCkimALYeCHLSQNJyOPeWpX4P3wHU8HSbWAnnJ2JgD+L0ZITWnh+pH67EM
LsSW8Vqa3ANBJxVO/UQ3hukZ2au4qMfNNpvEkD5f6qlW2JlwWE8RjFUVJLXqKVfo
QqdNuaOKVnxQLzSmRU4zmU/NvAG9qa8t5svddCzdhIfjw0E1H8+eq+RL/B3lMJLu
JG8uJ4A+TtTBySovyu0DJjcCrMcC3XQBvMZhef/xqK+32hSwHf8bMTab0YtAyP1i
qLwebY5wq33rQEq1nVM9SSfU+aZPpuUoUGc5//sOk7OO31/SRXLua+vpj2qEEnx3
wdR/+BdxfINe93O0nYwwneuwYDj6l+8ol/6OtBODl1uMnvsUxic3qfCH9bU+jal8
6Wot4eoKFMAOpkYYo28gCnW8lIaas6qQfFZD6vXh+DAjQ2rzFlVrWT1yUjWECaqT
P5OpEMkiBmr9Q646Jo/Qanpyqls7VF6icPfl+evNUhhrJUykDk7ru36ZqIe9jhHr
Q+yzFtvenv5/C0uBNuKTdEKqqX3No7M0OVVMYRpuJbpX4YnUAYCbYCyD+aby6ylP
0t6VjvICzJlxrUztQeNluUCnapEK5WrkSwqy3rzT3erf04TZzZNvGRN54lXGubuP
5dg4hTa6cRfL0n01XMMxM4hUPt13KTjmyJy4rXonMbkHjYLWNHOUGOZeqafnLjW0
L9bQtQjNK1fcQkrRZtEvpoB+wi/CVER3rLvnD8DCOlIqPct+ayhZ7CifQ0RiFxI5
FnQW2wbSErgBz2Ud4r8QHWAMhv9wt1swtYLBXupNk/iRmOo2aImibu7hLAS+QMgN
8vtGcUcMSN6HAS4IyY0nO51tWb+sXK+6PRoF1QNRoP0Nhh6PCBotAtSXzoANPpzv
oIeZQ9LCN2acayRrFWEMyY52/qXuSkjG+BxyT3rWktPUkhizkpCuFOgLYI6ggbqG
QFuAH3jLWo3RYBJvYD/8T/+RKj3M8dF+X78qH464KS3GaS/AaMaq5uU22K+o516w
U4Q+hvD5lEEEt5fFsPoDA511DE6sjbEg8n2MbQTT1YOE+Tx4ub2/oMmtB9okaZzU
XBiECMMyr+OorA8EmFUourZ+Cx9UhJbtMX7xLeUJOCvfDnDRcYhku+Yxt3MMg2G6
CbEy8D/z8g6yvodtU6z0i5CRu4/swEi4J7ubvkwa6a/re6LaVDAft/W6K2Eytk4R
rFVJ/3VsZmpTqaQVy+BXxvSvq+QNve2xDMcoq5YrkH1PcFkS/LKO10qJWrQLwByH
XmoD45l+HswT4XeK5jbD3++P3ONEjoDnPeFPhNij/4DbZIAxGPruHLMk0d2aNNXe
aJ8C0JHqFDJVxxHJyhN6segv86J7hGZ1lyN0GfWyGd3yn2nPMHV+n5tcMwGTMW2C
4JPt5wis1RMjin1R926DhpfeQ9zQWPWuHPGmDnueOH7agL1ARmeXanZe7mmV8V19
dYMNWfWJ6QE/iqFuPQiQy8EGYiQczLQAfCFxa+XOltnqU1vR+fSy/Ctoh2nw43oJ
Ttp0ynjDjOXItQjvP/GUz5+Vub6UlfrRlWcN6ZcdwWEP7Ii3HqrqC9nZB0G/lie0
c5AKY60Hzt6bYaJD2XaH+KkSsJCeX/Tg796Y9KcYqFt5Y1QvWJy18Ft/3CJPudum
uIwUBXJFy5CpmyxJ5M1Jl/jVReA8rRYcJctiwmkgWlSWYk3o7cjk1bwhI6e/j4je
d4RGXqP9SxqYsAsEfrkzAfS4gkSAlRylBdr55lpxGKZApbAHe45F1Uo0HvSUJPpT
Kb20aZI4CR3IJjCsIrDl6g/hXkq7BR9IRlmBOJO+Qpc2oApee7YTk0BE0BnwLQIV
xPAi14o7Rh4glw+JXyQN4pTAFVwOXugMnJ8hcl5P7q3VoUM02dj2RXVujdIqFOgu
GAcibjRSwjX7uOkjUYRWWUG5feFUtogSaLA8XFdXsQHZ4xyyoXQAaU0/zb6byxiR
qx8HQoUvaHFcDWkAWr+7ilnfYk2AhR1GgYXQx8beNGEU5zOwmYvHHZnjoJYDuH9f
FhIJtp26e0VCR7DRhDhiOtkkspGfdONwvqG4nUfmcuRk4me6giNQs9HiAvDzgxEU
C/9PC5qxMrg4/q0dbPjB9fP2TZlr0RauWE4Sugql6Yc3ozQu6X/bMtvNqE5oyFKK
cbwVZGKLkXcQMKj0jfRZaTACt9RLurD5sZn9t4hEvrcs/NaWY70gI6uPD/i/GI6I
4bTrt6lHjCGqb/uXluz6wysbcclpZWJ1NMDek52/zyyjXOQthti69LL1U05Vsx75
WyVtL/yWJEeuduNVg+dwVi2EXJH32WGoRXYbu1vRTkrwZPtY0ElN7hQgD5Ddwah1
sZ5zVg5TOi7MYTDpRA/y2bKeH8I7kXJz5uHL0k0ONiy1pbu+tTz2tjZvwr/SKTGf
VjucHjOuPR2oP1/f/b/CBdpwre6l192CwJ5Rkk0hPG7VGI8yoV3+XtVXwUGVDHU3
NPqPEvUsjDO071XHPfNqvxnwL/aJS9Ks5p06r71rIZ6Sjt7IWQHk0lLfsZchGI4P
Kdk699+wxO3GzboS3klAs0YN6cOpKWwo0L3qyLvuAEKrPH72cVbMLi686p+G6tF2
xbvYiXUQytc9oY32mRtmPYfPWTAW6JDjQwXRqNAv4Sb0MpPV3vQmWShU0Apvfqbx
bftWy/Q50fW9iw0kSYUEMh7l6c8x7Vzo1UJJjIL6XZVtaeOCWavKSwZBemIKGY4F
2v2jrhlECivSYs2TtYkeabB+DMoXsDqOa0ywwGqhkHtPBJ+CvWockiPI9Q2vcxVq
Sc3rVLGyMAHukSq2hYb0GXujPr5BZfS/y9rh0V8a5MGeEtiONFr8DVIJVOwwiA7J
OSp+gYBEtFW5hXxTce0fb90MDQP0js8DH2dsyzSNHt0tXeBeqjhfRJQQUZDmvlL1
SUmO3dfXqTpc8X6tljigT1OS/FxwInS+VlUTqKUowWcLvOQXqM7ntEtG3APll2aa
VhilPIylfjG8wg9b+gtwSUIW72jpeV7x7RN/3t6MVy4wOdvKZCtbQ/0ie6G8YfBa
6BiZ0+h2Tbll3Q8Pr7s+74vrk/CMiBEYjDICt1GpcnhmGCYs3fJZr9JCvhVUCWHI
QKHOlX0Pt23V1N3UKBkvb1LQwz/J9Ox1UGXICC5kieKJUb2pVIat7L6Jczrs1Idm
UmbURaTXgM1Y+mRnm+T0HdXosIWQq5p371ZkPwirZgHIyKZ5n2fVLedhyXPuW5Lh
6y2wxiiRU2Dm04OwDTX3IqdCPgP9nnD3V3v4c6zDmiWkiA9GS0/gc12wdkDmMSTs
kCdOjnXrQkop4C46ln2vnNB5jnnkUKJK0lMSS4vtHuw14O/NHeM7bJRpD4rG3d5M
uPIbvqMEOPWiFUxE4SXR0/Uc3U59xw814l52GCoKrkXSk6Hn7Ov8a8c2LA7EcwvB
YLnBhorX9E4VUopQpZ9fkKa9UpByTJDQe6pAEjygqWVpJBrATjI50BT2VhonorPp
aWDMZIRtsFl05+Xi5BgohbRO2y0WjmJqdt02TlYKEn09e+esGSHuke+fHaqHU8By
pPNGMwO6zDuBU+zLgWIdXBAMshuGl1srq9rVbevotxprfhM+2PRgcW9J8Fd+cozZ
NsvjM7VuMMcZ+QnLpJzh2F5KdBNXztfmanHkNcfA/Svt2oibnBDFNehIGcvXz36f
skIbj01jJwwpVvUPKlw3qGyU+uqPPty2CPLDTB5Z5IQVle8Aj4YNSY4kCUPhSYPS
QPndt5TIwQOCbHceSOnhTrjoaFjM1zRtNmQsAVuq7rHB0TlFyPYlnwm520dfnVoA
TWW5Y5qowvlS01KukQX4hys7lqFHLvHKnKkLG4tp7052vGaBg827RjmRnORsxXvZ
mdIlopBW0WtYzLuqffE9tlPfawR6CXAsQVJLW2fUc7Z2L1omkasnjI3vkVE9iNzI
JYtO9VzcuTjNj527pRjD3nhMWOF2er/mVkFvoV+LITsyj16CQ2wwTHugIsvhLKcS
oGKT9QEB9fQ38h6639fi3/+/RjzGf1NiTgJPRVZxl1oQwqjLEIg6l/Bg/RQzB1oo
DPC2NV11ojbrwID5udJT8oV6Bul0AwUgYK4Ult76RAvEI2VhCKE53xObXWGunNy9
iC1IRsR7MmjwnpgsVHhAN3cvfg2qNT1WSSxvFlM951HvYdELNfxDOfUjbOFdl2ma
oNnyZaJygf3XCypKnl9ZPCOiOCWiUwWgH9lHigajhSHXB2n1Jpz4hzGhSpzeQNom
3316Hphgipi8qwrofzqZfgrZVZ0p8mEXehpwCmj/VE5fCbavUp/zL/HOoKn8jaFd
bA2DjpDzYsnjLXGF9PCJEzOgPL6AiyWTrhUCDhgvvWNkpho/zviQ5YUnHZi8tiRc
2vpkM+haDcJo5OjMFlaq6YoaEImBTgXClGJkWJ4AP9VcSQt5Qyn49cmNhumRZFvO
z/meyD2Yh1aq+UHXJ3WzMA2TDukVnd7X1bDkJ8hHioSluFvMBQ1z/xE8RxEftTne
bxMvdbqZbDjulacDDjsFvtNebWvo/ExnBsjErIBjGzEaDmw1TGXCjOHpGtHq/RZw
F+JiBEHHZdVGWeFQzkAeFM3fGciQC/X9dGaf+0jBXDUpm81rzu3+D3pZnOe1TYhK
KoBN6BQPeWi/5Rw+hrGEEZG3xcZk5nLYGBFYCRX6VjLZ8V6K+J/hLzsd3sS+pc4I
23xgjssmxjOqsyCGToAbaf/MwJarbJbUlkiWCSNNqSAYzQJ3EhNSAdC1oKyMwrZx
q1hl2FJGXz2PV7KRLjlyK2IfOOVvKW/eT3hSplrncNzzX7Ey8cQKt+uAvHBCWz8e
FhdrE8QyJomGfKcnRYER9Yn3uoLRcUAhEunCh0fYBr9pO3R/70l4+cogbp3A7Su4
D9MSoFvyw0BmwCkPI3QzgpcoR1U3z2XBpkZQ75Sd0XF8rXeUrnqqo8WZbTLyaFu6
SxsUd8jns+xWKBq9xWNgA99Tx5O7yEcLP/SE2xKp0YPDk1kfPYpKkb61+2N0g69J
95uevVlnsf0PS5G29OFDHcOcPsn0M9UOvAs2KEvbF8eES6w5muH6LJpBqGlv1OPj
qAg4lsO4Ap5i2lQXO7QaEXLwR2ISXQ/Vf+2V81rnpftkOTYjOW71+W7SzJz6j2g8
MkAyAl/owdUEZT+wVL7NImqsChpd+w4gHTzx7aCDGuXB/KI7Bt0sWP4KCY8jOkSH
motI1ifTYh6CSE+8PD35xCMqOvtK4/8wdLHi2C/QYUaOX99RDr1hWBo77g350mpV
uJ+480ZlHs7eY2p0ezStkxOfkff5txQ6S3NgsUQk6CtE0Eiys7hdSJ3cv6jiKMUE
bYqzcOVTmRhCUm3jjHKo6STCeFjEVCt7htLCGRPm0zRJA0NYPRURR5rcXwOtMqgT
yg4zaTvyPkEaUv+OC1GHWispLZVOVMaaNdQ4YLVBz3Y9z0SQ0GyQu4ORov2rovti
Jcg+L8NSkWy2bXZMwLMPRQuRF1I2kGdhM0QxrBX+Enk2XAETZGez65yUpXxw17IV
zk1GIUDqy0bmGKLRxWWWh3SedOj4BY5mfxD3v1jxij1HlHFHbzLCW6wSW9s0Z0ec
eu23MvxuPAB/pDYNWD+jWKy/TF9ecps5SFoD7xOUozfkvHN2bf247Ga0vlktyj78
X/XkO193zyyeBWUu2UrKIod/1siee9gsecT5JcEy8jDfcPV8v6phfq162R2mGaOG
phJEk1D8yuxozFVmN8qpjkrOtzgTSGrkPdFvGFAT3bjAXdkG3K+2ip2m/IryFBR+
ogLVho71ez/mgnogQheGShUCbSGsn8YWUmxSRwTfb/ZNGqg9AGa2p6ym7B0Hvokh
QqUig+3z78KcIAb8+rd0PKr4eTCk3QKp1jQaAZq7q9jHcQYZQ/RS5vYot9yGnX4g
M6ZZuNk+eSmboORmxwQejZaMtnh9enBxLWY04AKANzbObtwnHROT1s7rvdom8SCh
dvn8vVBKKoMkUTLycvU/YRM4CBxkXSxmX7DQXxhcawUewFAw4GfA12rqRcd0bXce
ZkCNfuzCZwMHh/0t8ERzbycpMEchWOz2LCGQ0lsEUMm/KVVR0P1od+TUirkxVTMT
UF6NeBC9FaXLzoOwUS4NZnzweBGVGeSahMbL+sKhUlFWwFdV2FkiQz+fLl6tWBhQ
hLAXFmkJsM13xAL7sKR4pvI5xDCfWV67getiVrx0e+NyPvxT+CpgdqNoXIyAp68E
C9uayyF6inn9rODthgbXWr+uPAcGqRnh1HNE3oceumhDlcgpXbbEirBsMO5QCP1p
bE3HT46MLUefPe+M2tVFFhN4i5AzDc4AU8sPLE3Kb4xAw/qWihc+3Mu6/hijyBn2
rFHIzQxisQ/YdnajgyzvpeZeaPESnchvB+LbLXOwxNXgdjR+nNAN6+hC6B6EkWd9
Ct43oQ7r9OjuciqvkOlMjpwxDNe9wzshP1i/wzeeIuFWUDVy89GhR4NNYloXmmCt
sdpR2HZwDRq9aDnUx7x5jC89rrrSu9IWF9rkMPdr3Om4l89ub5U/SbQDe8yAP0B8
CtcZUj/b0wZYxK3cKXNWRhozffEc4xyCbj+2n/vacjb+S0pp+jrIlfXCmGY80kPt
Z5OaUWdAKVeQtyAu/RhNOfGi6v+nFugxB+4pNjIkxHtcZPQEIv3xZbVE3g4sFOr8
cCWz0EU2pyGIj/FgPcGbrPbVaWHxWOt5Fh+oRfKkTxqarmD0bYhLJti5m7BSMURc
aE982sg+27//zyupmEliQCZ7OnQn8qjiVm5GRuBlqbANt4cxaphNb8DTb9kADHr9
jKSkA8w2994itCl7ExYsjoPHgWWCbg3XRlYg9wKOlMac+qexjxQ07LHu4Kg/TebB
4cInS6tcwms6YbLnRff6MH6nMJ3guIYumIJX9g4DOImg44lE2w5oyUnjsdDH86Eg
mNZO7bJdxSexAWCOYdbLaY1uRtYcOiGPnDRwHQnEo7DaLCo+2xnMA9NxvrDB2xhF
lqcbaFzXTIO6HGvb1COU3AmaAdW680Gy3N8821bwTptNNrFdmQ6yoqSMuQPWJ1dH
R5QGqn5pXH7xYauwLc8979N6vdyUkj3KL+MMwZXQko+JIokeAJjB4xQsc3KjdDYN
35TuFkdTcV8HaQ7SAMn0YkopbXL5hV93+aEAP0lxEa7UiJfIfiSZH2WcYkn7f86C
N+rQTT7ajFteMp57KX0nQ0udylVDSOQMIBTGT5uJ/vMc1h1iJ3Gj+H48C47Nwf4t
f2Z4GhqYE35kG4Ll6KZJH9zgYMmmMS1hoRwLcIuoBlGHKwj6MrSZd8Oqx3Ekc/F8
iqxCnLimnb2DQ6WIgmJHCIkLiUfcrrCn7KRSuYtv51TfqPOWizM7LrCpJTKQK34N
5r1CSsYfwHKIPq/gGtwn+Qu/r/3k5aSIfZGki3oypF/6kL8FF8k1MD37Uk4q1RhZ
N9uNYBegIxxqqS1AuzjFcGR+QNhIoG2SA2v6leDRGtxof7+LqGDThYROT6TsCnQA
2dfKQshim0QyL0GC/XpyhLDZyzyQfsRsxiwqyloUPc4Pw06lE/ICyIkeI7arCFtE
wfaL85OFC1lGpczMq5XMxVBGwNPDlQ/RwfqCxDu/0eRzDJ2RVJCWhNhoVJy8PiWH
EU8qzf9JRoK49wA0VC27mezbVf194xx2o6mDz6S6RCu9JDvuBVmTmsEZXQyhTEtj
mP3ql4/KcwIEjN4SRzFLyuXOzJWgBGbnso3k1dXWnn8RbkAV8W3+uheVhBVEJopv
BZrLRb1CGL+L7aqnvnBNQSZRS2tJENQOFepGv7vZCsB3CrcvZElbeThrfctTPbI0
GhJmjMJ1cSlkHy2ewwLGKp70i+Zqy3csEt2SU6D8scIupquqDHs859bPsGqd43eu
eRYPpWlGFOrJl/m2othcDa/4J11aQi+9CYmkKtDSf9vX4r+Wb0DLa+kP0ZimFYCN
9W/gNlwZiEIX6Od2EzHsOfwv0FN40Ll5LVKH3Gg0h1Yk2a3cZl3dlU+An1NMDnlT
3Lnf+h0Yl+Min/+6CxpQpK5EtRwWX0H5Tp9gek8XSI3n7TLvczOaW9mTpR//1kzI
tJ/humIFN7t/i+VGWQPV1unH4QAXGkdBPYF+JXunocT9FUdumYXiEYZ7XB4jUkk+
VpOevYowe+wOrrt7flRp7uLS+78rErQ8DgfiTSj2WF4tKipj1pqZPAmcwkM9gK2l
4NW2zAFc+E9Jz333OX5QpebwrZFr0XZpC0ymTyW/KzXYQSI146pWlpPc8LGnMR6V
pIk5ACVY7aiGeIIH4iTVlevanFI5jUhx3/eA23muDyCJ0ciKYjnm0iIjrUXDMz+q
6dOo1BTxpOaubZAHK+TrHjBOGe7kk53EF2/htJM7o+PgAwuUbRtkVy9z276sOcyo
jc9xEPBMwfjoR++0cmzU38dOCGAX3W6uTAfe/i/N4tLeo79jSOmwNw4iS0HqtACB
hMR+AuO2bLZcA7V8M4dR8Vde5fQjd8yfPRwVXOHo6s19kwlPT13X+9Ts0rPFeJa/
BC/pvCDf/rJieb+oVIt+2e/KjyFUk4ZRViiFADH7IFa244KLJSbBj09kaP+cIJfI
qQqCGIJ4XHium7uZumRqPuvBFl+7d8Bb19TbHXcWWx+u76zhB6t7ZxBX7F2KTZtf
0kkrB6YaFph8DM0uStK/SWpo3H8QCc0+ykbzF960hiaOSBPknpoQJrplwHSZWtfZ
eWrEHen77OYusQli0U8AN8lFtRQR9+PaO+gKTUbhiHPFmSjwZj9y9ChvC8EFrfaV
paPgfiWFX71L3gkRYlil+GFNfSSKpRVQ9vHR8CLhBvpnGtH+FzQSBctzkltjUkHG
6Y9uyJfAydoDevu9PtJHdoX/ZATtaCDvAbv7tzED6StR5WtPmgn5HLMZg8cASnSz
er62JaBWPUeYHDIo+vEv0fIe0XW5LPshdJBBRCOih0BMuNZ/TzvrfslpM/SFmbzl
nOaKxQBJOQOua5G47BeKs1lUn3GFOxqRz6uzN4z9YFQKaUMMBDolHsQhY6AVtfsy
LQaXFQIPvnTXRG8U9O3hhcDdKq5kNY+meVfVxxgmxdYYbo8GUK453QQTWoWVG+6T
NPSF58hEYPho/OKOo+ooaVlgugDlKnCQo7oYY3fQ20mpXsVYeoW9RdOrystHEXHX
E0Huk9+IhvnBU/g4dhHfy7WdZTbOIaVFTI4IBnLzQKFn6Tm7ZHyjVluuiwIsCr6d
icSqM3bNBtp2FPPTs/1sVVzxbXJWsQCvNbhpU6VEalM2m3XY/GW3OLVEBNJ9XI8x
+IiobxCbHfthQyZbcVg+nWY3KbDfVaXMBArxOF0iSJT0v/eaqnAMAQ/fsfJ8UFK6
DSlzN16yiaO9irrAriSRkZ1O/C60CksK32I93at9KVsC9H4/I5JeyyTk/WHvE0A7
gUIkF7E6F3Tqf16Ur/KKEMLuijgdZchmfXGaPAvfjfCtg5ZY1fYZUB+L9Fxkf7XM
hCOsDtkLUhU2w/BrZChIsTWU1YfeM7QbsOYnVaJfs7qEXs1CCMzKfCO+idHaa+OI
gv4zxYAB6auH0AO6m+jl1ceJrEqqT0wN2tRAwf+jOu0uGc9wDq4UWbiM1xmT7GSo
3H3439smA9GjRTBnXVLBWd1kHyP/vKrbJiFU32JCrFXELMMjidOKHVbcnLTdSktF
xWYTg2RxNv8u5yR3K4N5E9abhOEMOyBGnNYFlreI54d0Jj9lHxS0ZLbngRxuiE1J
kHkL4Q7BIdBaqiR2GpuaoL8xjEcqRp+tKAtJ7lD1ZOnbNXhCQnvYOHBiPRja7/9O
vbkgQT4i0NH0rBTaxJcJf+A0nTRJjEiCox+GJhUc/Nx166Pa6dmq0XTtVbMlEVzr
yZPKsdH7j12oWm9MHp/lqfgdDqUP6pi0WvqbWDMSn0Oh25VfXWw+tI1y7R9UZyK1
pnYtOQT30IASlEeoGcdWE3jwAvKY2UGpxCv5YpcPQXLmi0VdvjDjayaX6tSNqiun
l0km7dLov99eOX1ckJrceLQ70wq8rsz64Fs2A+Ft2LY16zmeyj4q6vlG/WhaCoCz
yLc0yOq8dJ0nDs9xR6ozbJySiTKKgRE7d+h41ZbdLR72GXHFRcsm7LK3YI2dx5vZ
d0owpV/q4xP+j/LwxoFiIb67cjYJ3LPI8S8Mp/XNYKry1FO71rH3Ik+5vBnLyl44
KdjgcbnSsC/hR65zl7Dv5tqkhrn+l7wu28mVzvvcU3U5H6VIitJ3R+FIXmr+B0AQ
x7HZBZ+lBzcbWSQex5ky0plm5GXltXQjNggSIlNaxmvYalvuk3BpblXC+t3QXiGE
8ehNaw4PRKAhpinLkBGmx1i7pO9qh6bZ8zRj9TGnG1Uud3a/4JRLnbSNxpJI3qzs
VY7GDtcrTtLyPx1TmUhZ3/atxS+a2g9tI0MKigY/Z7JcaVjwcQXIfOVAmAEMckwP
Vm/uL8BEO7UCyT3osgNvLMxBWUbmq+ZqDbM0Flurj8vt83cLeEQ9gFMLM6/aZkA7
mu+NeU39bmBxqyjPpxORjwkRTRJotVp4HPVAAcaIFANLXGVBCxcfOZig98Ut8BpN
xCVCA8XlrE5r1DN+Fs/mstPwRCfNEetnTHuLOjU7rr/+ZEQQkOfC1rXifrb/t6aS
j1hz2xhxdqQUqZBVaKi+GbAtqXSxeBCW6yr0nOCZhSXMRzL3M/OrAk/kdO0xA2gR
nZ4VgFrJPVYej+Zg8MesbwrX9X448rEjO6t0TNC64oA+PS2HAk7sGuzMZ43ekjH8
zWkpkWGLZAkK1MK3UnBu1MqgldSRHlgYjysvGnQ/2hCPG5FNLuRx73zTUJgR5CRD
W07OjZKJ9kJyoNVdi2KP5JmLaCxpVQoKYXvjaWfRtvp3AwkT8dt/LeEtpr3sS+Q2
gVKgkaNCUA0hfpuV2Sv8kIw2Bt0HOuJjFUG30GdKbrNrGwT6lhp/q1P7S1nXsgv4
9H4LXRhN4+/gUuC9e7dxNRxb2Bwbj+8ymPXRacINnc1pgWj56CjSZwV38U4P1+f+
hVNiznfNGJKI0fjr0JFQbqrUNlBgwcfCM9vXL6sBawNQicjRX2IZpfIg5mSks3K2
nw3dMuUHVRAbSln3yEcBQZBraw+/VNjM9ZwkpV4+Lybxc0w9YikaqPYZ/5VdLeen
gcqSwZ2URFluyRdZiAwQVM/xfjiITjk8Rd8f52YZgPvC+I7T5EzzSx+LgMA5PSL1
7KgGPwA4KmB6hD+jK+hsl0F5U74pcCL5tBP1mOCIleP7JFvQMIDpjhAIqgw9WiCV
UyTdRJYn2q7JUsc0NrHiyoIdexyCZMzRGErdqWLHlfvpzMYs0WADgObIfewPGYOe
SesShOuCBarMoP9Yee/GC0AEDppFcm+X0u2TB/LuNM3yj5b4FRupBlGdTT5AYcyQ
wXSAYKyCCNVAhREvEDEzbpkCoSDVyVZzEiq9C+xCM3iOu3mk5fOVD3koLttuZmsG
nkLhnAw8cFTPtv+Kq2cdwG9SEHxrTkKozQw3TQ5SBO1xsoPiVCitMO/CEDH8GwN3
fnDWJJf10RHJ1b8PwLPjK3VjujPdihRKHChIoN++aqliLgaesDmOSWZ1/BA1Gtuk
sc05glJYpflInrufE6ntt5/+m7eQiaEPQcwAaGgjyBPRXEoSPhp0HR5yBRyDjGcp
XRPnE6ApkHPfMf8uxpQ2EO/xaXtuhTnpfVhrqpnzy7MIJI9xW8vPS31VaUiApWP2
Vclh+biiGXbJ7EfguCat9uqbB0/GsLKLZBwEt6icgDDKXuPCRYjDKTMVlkcmnbAD
Z1mXZQOryv1elco51stKuYd+oEws+2TrHipacf22Opxm5wQSYVfqSJ9JuqFiUjQ7
BjdKy1o6LgxxjJ/40HqEeMLGIc+oAyBrkxBruJxNAg4zAUt6WRl9OLph5YsDYZlC
aFwObEy52tHW0nfHrsU10KeSg3pxkYUwQ3+QUy1M9l/UaH+NQvKEVze6nrxU7ge6
812q3oKwtBGDOmzZ/lq7tN2sRU4zPN+UigQY8aaQhvPfQpXYthsWS7CnlqrQOamj
EsnnQJ4MPL6Yg9AcmzFyBHrjjfP8yABnsDv3Ju/yn02pAK9iVBYDbKGOaZEphI5x
MEiBgLBTkfTDSlgbvx+CZVel8H5Ly4JHoDEMvG3r3cwFfthQCvex0dpqqcXCbi8a
Tggq/GhMnI7vKrz2mKR8yaPC1qYb6rQQ9WgMvX8zn/8vnB68Izy5zr3wDsPPxQgd
S6nut1oHD4bDUa7Zztm4q3dHd6ijZHUmw9QM/+/zj0tJJxT7z0YjGWPJiwLdSrF2
HzLEkgscjKYB7YJIax2Ko952dfcX0Qmk8HQ5qTLK7nG0JGv333DME0dQj+re1idp
vMPw76wxB419eYl7icmTD+VpwbJYFH0e/iwWoSzK8uhmKIzKZW8QEggdGsG/P1gv
3yQfm+en+TBtRdy0GLgC+tMMqRcFUXiMEFRPiLPPe82M1BB1zjaRZGA4CeFCwIU2
kmrcZcSEAYfkoL+asvOScwC4RDiM/Zeek2YrRqnBbRfwYz2BH+D2GEIn8XzC/HAh
D8jvtLENiUD378aQNd9JuDdWnvLDRpld9MVrd6YwAXLeqmRhim4Kb99GiFJQDaL7
TdsBjpLkL9JXl/fV5T3QmBZ6TyyohWhq7s/hL/z1BfnKpcApcyZvpCq5PWW7Hakq
8H1we7WIy9gtTxOFyMzjMDrRiXRBqdUSbB55FODvZHzDeD20uzsf9s8x3cM5FNsT
VJnyLmN0nITiis8UVbHw6SxmSmcAzLG4EGxtk9LlGeeKrirYsp06BX3sbOErz26x
gYpLJSUmXk0H/laK63DxHLJh2eSIsgcfhKr+2N+e4WmWe4l3hipaLBN7N8aiHAXe
PoMqtajiJBAQy6gv+liDagZFV58OScEeYcpsO1zenP06Xvrc4yqx70R+NNuahBBg
YV1Olma2BFtGxkYS8nrLlvtcThg08nZQdh89KW73/TXTJhtLcssoHqYmKiuJgdGV
aE8kOfcLZu1CgKdhKI3K9woBoApzDPHDG2Hp0TbTHEwJIrEplCXyjNUYuBb7HEe8
Q0HLHtyA9TNff3jjL397Z3+YH5cwH2VOs3nU+IOubdHD/M+XR0IErrZMzqRT1tVX
DpLSPJbt+YBffrkAmfvVLe5gn8H7/fghjnbuFhCVAEFe94BMUbYq6yP/HcE6R1DF
F5WmtF08Wq9f7E2NODgxk2F7njc+0LEVH67ImP+o8KKe0kPTvl7d6/3vmCoditDi
QoQsPFUQUun1eTMQrwFhDyzPm1DWX3n5g2uZKY+wc/ILqTou7qGBbY+0sqDrNy55
x4YNg1niZm10h7cofhN6vazmZIFiB+g16fyXJMWHMJeNHG75vf3F3QfvKEwV4aTt
Z8bV5KCkymtdP08tPFwM7ne5beGWLooDyIEN0wqHSxjXHeISvKx7B1wwzy6+2B8k
wKAZqi8Nac2YM4ketufSpfnBSLkyClqHj2d9DqgB81iBEayNqZAUaen+jHyyVJjk
ZKfMs9XbD2IsSmBF4f2eXbMTQmWyAy1yLYIav7pet7lRc0WIswnmrehC+TgKcQbJ
Q9xdwkKLJ4FlNM/7nNO81K4giOJtu+3TKQogToJqv2M4XRBZY+rtJU0+LXZUOGji
C2Ulk3zwfmDwpep8/mMnTmhQ/sfA39F3btCW3tFB+4Zj1dQMDd176kkXiIM5v098
hYn75kHthtgeMW0VDd7LJjwucZPeEQZNAw5ldAMCvBckKMaEaqZgvKKxNJ+lV8yW
F4m9d16LKDqnfd2ajWWAubsv0kQjEFzsSPA7Wlwq4fTXzM8KBq5Fw5dk8FHcA0MU
5kBl8Yje3sLX5/6l/aLgBD5jdHaHeMv2uaRyn0bqMjhBGrwAh//G8WPw/DNH4aWR
X0+Uoq//UuPtAhrR5yM6NXy04tAsLUU8TZIkkZarie6udJoP/ijzyd0PYmS1lJ92
FLRNIqyS0sTqsTmdMGRH/C1fvhE4xPHx8jdX8fh/Zu/HUw+MxfvbP5Jpw9OhgFdn
0njsBGz1f84/NucZ9EZEnyLi1aMCdfRkoH5ww79nx3boqNWMewapmity+0OH6Ifr
qjTQQntXMtf36dIKK+UeryJyocR1UKFiO4ianKZucOO1VLOcaZWcduZi7BCt0Rfy
sX6vC52rigRFQsxVc1NX1k1oErFHhOAfSfscIQvU+QZ2BH9F7ADfWlV/kMfyXIXu
1IiuZYWPWTNG4pXEpAESFN1wreEDoxTfYqT8zAI8rJ368mlfFhO6RE6yuCCtwM2z
JCpwvd+/+YvJt/P4ekeL0aHkoh43Ms6u6p/XElQYiwndUShvg/xWf9Ghh5W1XBiC
JDh87ld5B3ghhUGLDwVT7fmbPFPpfk77g5MgOOvn6Gz9uW1l1RAyRQpKAoEeKduG
Np2LL1XgdtCXDJdpL4QgbtzboySnY1FEllLcIqNS1p/Si43BRdX2t34zQTTowXzJ
C+T0EwXnNWvUyy4jr27zoKnG3YSlG4XAP0tGQNz2tWfWeSxtMOxrxhq037BMm/Cx
XhKbBGCywrIRBN0aIk9ZBE40eQJ7MV3ZW+cLz3K2LqQzDt01jW6rm/YWiP5RlxLL
C2QLyv7NBvPzxgum0QHyOZ+kHjXaeqpoRMyZCyIavtaQi2yChzIN366DAXiFPiHG
+8NBlwYfyw9ccqiEJQhfN1pj0b1QJuvA90oVe8crB7gTsw3mVTyK82LBVkJy71af
Sok51C4ditgYfVxeZ2/TvdqsPjFxyISPt58CpSYvANGvfFguhPQrahQFJq8FEQ8q
mZu8UaykOwX8nbgnqJdCzogfPqDHwBAJZ53W0GgM+DspGPhDpo0y9Q1wEljD0dpM
Fe+TpPyDusiCOmnelM6HLp9SEHgajtsYMhhnOvD5XUQwgszn7Z3mmdXXeAr5jC1p
eGZOKoKQ4yVECVrgnjL8LqnE/c0BWvfUFCPz6a5JUY2liAQHDYqefVwAswkZrQWm
QZalNO5OBoZAKG6ItyjIPqwifOK7r8QMRVSkeivdwKYYN+v4jTl99NWcaPBakwX0
nhW6uPQK03C1TqnFKSVH9yCmuaUYZbu+QAQcXb53ciZSiBnknYTuVakp6u2LZ7tR
4WOf+WJcYoeUmSe9HkDDPJ05TUBFv6ivfHM3vhdL1wSnosqex0zZ3/HoIB8AHMJk
hjL5UQXoivXxmxHDR1aT1HxSlT3WWwFL+H8C3jDpgwwkcCCmR3Gfp64NPN9aSzSx
mXAL//z0F6zpew0lJDH6qGhhjEPSxX7mTFGssfwAkTgBgFfcIuflUjns5oNn/LnA
FtIlNnU8K5YMJ0phFJXvlEuNhgtN/MDTX3OfSk3xEgNE3GMqa1bDC+mkYspxKlr1
yDoVPD0fl/4+coq234NBcHTzadEqBKbqurKBjiDf41CmrROGctc2lbZ9E+OVw7Y+
6w9mH1nqe8YZzf0PspxgcBGhxo5UqYsHYjzXCUdrh9oPoKD1hF/OvPyaTU0wU0u5
xLiLBoTryV45/JkyU2cVXikljCHMPgQ6kmckyEmLeiUZ5BYDxYzLIFZgErhftoG2
gprOZmabyy2407XXYNh96ZWtMLiIIAvmhek9MZvTWoqVAI8uWvBUxDJBxn9n+cyY
1vQm9uFxdYs92lNzdibuCrn1wGvcbBam7ABryygJKW2RXyk1FW7KDJPIOZDhwnzg
xGDmhNZFjccWVT9AowM/hOsoo+vrSs+JIlJW0U37NHsx7hsfDd7ZUncA7SkQN9hd
2vGeuRQm0N/Vvj9AwOOsCILvWw93Bz9UEUdC9nDv4Np2itHCmCMTNBp2QUiXA+g2
XUGdkiB1xm0QwXzXStCCcqMPToRaidMxyok5Mj4EZfQwnCm/GKgPGFkYX/6Uff59
XzhUJ6mkXKTW+s8Zs0aNx91hdx0S6WOrGw57/+MVcCR4UybD3JcqIE4Ogf4rxoOL
SFA4bh2ZCR/ZRTXvfsZJTTHG4LN+Dt9NsaH52GPM6VPH5z9b9mFOgAP0k/5+LwHO
Bmp0Uja+9wL14xfSl6qf4k6GMpLdFZ9HwejnfNaJtm7oGOEBJ85UFPneHrUepOc9
JSvmjaPcHjj1p5V0hVyDYgF1qYuHVE6lEw3+5fshSD7vbIz+UPbjfYjW9I5s/Qnv
Fip5LbTRmjIbrn8kPLPk1igRjrp03MGTMXpzuirIFfcHa0loCvEXdgapUk+8edyD
i55gMTX5wsVJDYBpeKQUyjO1Clr3e4yQ0eoIJtbjxqvo4rFkS74BMKq+nc3d+iPS
4N6W5K9zwCwrrz+23qVYQ3b1ohbIIRSL0EAAc3XPzH1uzX7E7b9CpT5YcqjLldKp
c9ZhT73i0BkzijkCt/KQsEsGJ+KMClcNQU2Xog8a/K+gN1m3aftNXVY3f0bDhIoS
2rfiIp2W0XLh1WOk4cNMp6SyqwbeaKIgGG7bjcAb11uhUlGTTlihll+g2Wnz4hzg
jG/qeMlqY3H/4fIPpz+dM4oapXjTMkeuLd1LNAWhJmRs/eRg3Jcnqlra/8mCfTFS
4sg0Y0z3tMYqutQ9J7+Kc4oKoof9hjYe5pam2YW/Fo/Puf6+LBDNufWpULOXR4lQ
WnVb6Tr/N2ud+Suy04WtiM/Z2PZc5+W7LTIUhZj4AS454CeQKdIi+uPMxD8HweQc
4Ehc1nnqlwOSXkEH2p3BWWSnDVn/oHFzyxtAqds0Nd8460loO6SEr0AyjWNY5aOq
UGhraMuX6pfsZhgAGX2tN1XRXhgVEzaoKh9vE05pVrownTKVV/EMZwhXKK4BPWGo
W1gfeMXX049kZQ2VnfUuKF80mUrjWe3KS/kk7/kN0tbssGN5e4dNzWGrSxfPcVRE
Bv9JKcpiJJns8J6RZ01mRr5ff7fPdB+b4BRv6YDJyjxIqEX5UakSXynSDYZmLwuT
FfLiojTBNPYblbJNsL9RrqaJZgpfdwQfquuNI/C3aOmFzOwuDD23XM03fRvg1rwQ
rP/dDvnPxW4h4NsIlxv12hDBQrY3/nljVRh8Gzl/B1ZmfJNz9jHSd9fix9wfd/3l
P/oEZRH3vgxSwcXkszUdqMHf12wlVq7QhWhleM8mA19NpNHH50bFgN+DRkw/7X0j
rEKuJrVPTXcii95A7Hmx9zCR/1Y1cxh1HhjIEQ4iXnZNx7TeaNSkL6N49vhUM/xi
Jzkqv09GCEBUu5Z7q35hP6ZK0qhwlRk6fZvxWLHRd/d2PL+cKVM48LTwI+rusRyV
POvo6kPEaEdp5PV4T2GnE7iLFV2DoqukKjNv0ObtYeH6pJXu3luQYHANz/4t1zNt
tYMmGoxr8MTDNbzGmdSEtn2coGznSbZiCgLfCs/lsAXgiPRbtQPNdhcUZKtiPqRu
tlrVQK6Ac2vWw25zxskuFq/zO1OquWTCNascK4vk29GP94+5j2fE2ZmgvxKNcmiT
GVgRbTgCtYkGOekOLEJ7n1EJn2vE97aklExWV2FiISfhLFgKvFPxTsRWX2sUhGOH
fMkr7loZYQwTxFGIA7Ve5NwcPqM5O9Gv2GJhdruP5xjIXt/BuzykOJoxoq0gGNGu
3eW2iYTGiq1GNsg1+YkstBsvdY4HchpPNzB+JMyqtQ5tVGzt2csbJyl/+kI6y6bH
mAfHCjhiex6iJ5BAZY487CQ4xK59SupGhWRySc3rfrWpNMlJ0+tdB1JPtKbPIWyX
djnvv4QYZGhHW5UVk3gqHmUsI5M8i7Xhb4R82VcQ+/MPyJgDGmHXT3XiD91RbTNg
kwEwkGiFHmdgzmI8JOddVKLlpS+SyDK9jsV0MAs8RA+sDY91Py51N2f0l2k3cuqQ
LNXWH0KnzRTwoNvfQ5YfYDcVh2gRd1CTAYzb3K0rCCUuZD7Di1y9umhtS9pfpnh9
1kcAJkIEY7Zjt7InrMJuZDQq/u2IJNNM43ttfQAq6d4G59+3Is4KkCVNeKbxwJWX
ezdxbACDltEzuZQbUwpQ0SFz4FZKSzyhdB/d90qothSCcdHpFVnoXyr5XQxAILd0
CtMZEP++L6dEdGApR45ZzdQ2el15S7Zdl84mN6Vvuy4FUzH4tKS2WzQ0Nd/qtjN6
AKnWhuwZvLKSiUrAW46YSxC16DxUAavUrnTGPoUgI9RGqwKfCRgvT7RWbjbv9zqC
RHQ+xrMJ92azNbza9xXV4frDTslLHNkK46aftIMdXiR9hKqtLMutH10KV2ItLngk
ZmxlRwWRdKNiKT67I3RgQvArM1R5cNBnlZzlgcoEv6UUeQCljAUN8jwynUY1FnP7
iF/FewRq/+ivWWFfbwMG6BHy7llWeliThJQOXd8bI/1CYN9MZoEN+R7xdCtoLDv9
7JkY1jnFwXOt6VjgjcrFRpkw3gjtiR85n1UPV0gsF7pSvaZSYG40bQYqPEzqgqYk
tmUW0o601mv81TbVFrRY21ZAp4hwykYJr6FhCuTBMit+h7m7OeQUYgaVfzjFySxV
haMl4xKOmekXQneIx6IrFw69MAlCgtbZVxtk9XD9tqIibUohltEyNRgnP4nedzCL
O+dd6OvMOwm2J/ySId7qMTFZRBlBtdLXuru6F3dS6YKWgU8d3KpMCktRSHtKaqV2
UdF7spQJj/K3Rh6wld/jnmEUugDHsH9rwwnqHxjRHiPPHUzpvN7yaIliInaikhFs
cWihYUmc6Q+n3YwKjRPiHItluhp3GW+3WL0LOWNKGiWWS33pQz7l7vselYRmQ3/Y
NrPSvctFscCFNcZv4YEowfchz05Qlg8WZGVx5OiNn9Bc0V9sMyc8d9PHxPOZxN1R
U2ael40SeK0ckt3un5vPsnuOUexBtcCZJH+kB9cOJPeTjieNPxaZKjPXJksH/9DV
D3YPtduELJQq4Zq31o5X92dOE7BCWQCHrOfH0pWCPiBmODH6iVihhFBlXzM2r4PI
uuZpa3XAhsX/8Wns+RmQueWUahCMn7oujlL/asMdukmi4nl4xC4EJ8bq+ZJiOb/s
8bB8c1DxQaVWRu5gewT4oE6+vg0S4/3T5QMFyNdVzp3fVrB5zS/d9Rwa6pkGSReB
P3Sq0NHGuwrJIGSsllqNP0pvStJRq2w7wjp0VXzJmialEKcbfbsZsaQBI7N0IWuJ
zq7bg8oD7hchMzx70bKCg9VeHIcUqmb9wy7dEqmUqk/tfFNpVHNpPxwBBP6hwqlE
O9FpBUE7lh3yqLQaMROc+F0+HDMNsy9XnSkeIv3Mq7QBfzEdmUbIJLtvVpA2iGxB
DaeUZKDNntpJOMUGgTMqVMptZcyTBaXzMv0XOlaVb4XWzpydveQ/UEqMKyA4vRg3
sKu3to+D6i9h5szk9pwBzXfjI2F9jRlkLirKGPvCtOBDSuMlg6El5YOtZN+9yAjc
FgyDaCwvwEM3eZL/5ITdgmF+ehDT6VrkEXbt0YulSpKa7uyxnWFR5MnomXcq/fvB
dl4h+ql1fqbIgECNs8H/l7YWc33U2spRCN2uPV43ifHinPFTyQSUhOVASvcFnapd
FFS8zQegkvCZ0RLjSaT9eV6qCpcfBmErET4KAaKdKKO53c6/7xhp7HhV6fnB5cz7
qL7OlZjtwNkF1IsOyUKvokcn0MNJN7e4LwxFzlOt9y+UufcMr2/SjhMbBrgwX0J0
qXXMBmtdjtXATgyYdLSAn/vUY6dnyN3E4tjjHf1owkbB5nJhhJcWREDnbmXkJRZP
SxvtRXtzDmSk7mELVQTt0TDBsrcrnn702VcB5ykCxI9wD1KOQh+kc3nWTjk+4kkE
yhgeoO1gtZNvoZDcBKSUBWSIoSAPgJaSGJWcNhUVBSktroPKIZpTJ2a1vriLaAC+
zoUz52fnn9vlLsC6/IgQ6eiUQ+1zvV0fbsMwU1KO1QD9TdWkaiVDVnWbZmissOsx
TxiDsbffX1j9LRYm2Ldz3RVYxf5bjtwiJD4J0AZZw0gdUwtH++jkNJrOZ1o6qvPo
uzCLinDmL4OZ4VB3ObstHbrW2mYCBevsDJBiGvzDLqQasZQRDj1nUZSf6ZnJB6iX
jvDeb+dWsrzmBBO4YSbpoi/1Pag1gQS6CZWtg2zM43KDe/ChKCV5NuoMxOK/pXHb
xShE1EgArzuJ/qs7DagaWLxBkJHMymzI1UkjGO6Ii1T7/EOEZym59wiWrED96Yfe
9a/K8RUXrmrdO4i6h6nZA01XEl7r56pOfPQHbFJhObIL3ue0ZGdGMQjmSMrG2aAa
2dlHUDkM8B5UpwiFs6knc/DRP7gbUPWc8wzqj9Zt1QMwICu7lRzk/VmCSAgDvPeg
Q6vlZrSnqMpLi6ckt92WQuwCpB8nAKFAAdMkeJPoFyapKWQUQGDl6vX0IHOg1s2Y
JGEae8ph68XxyRHshlzZiLhr4VAJO2O8f7j0tE5ZyRbzcFXiVs8Qk52lCqjQBszO
dias4IRf6K7JAzfQDH5B0zbyxkIoKabHuwYXxe3WWKovJlBqqVWVCXk1qjZgTinP
vYvpuaP/WSDf8WBStrqXoIzsoJ5Y5UdieO7nALe7SumhHIB4lBakv0DRL8qWnIk2
aduP1vhz0akWbqKo0zYpfQpZU++zIUbd2grO4TJLqzzdcsLCxuZ4gBV8rT8ojc4x
4JYjG0b6dqz40VhpUDXDLQifGcn3Hjvts0/5sryqKVtgoh6uUfQnuv+xi7TDXroJ
M9jU1gz3U0myMX5cPGaraGi3FnchGNP0Om0knTr80XDsij6v80xEy5GxLdHHxSfH
s7ysHGSY86S4Yt3+sUQiz2JLDgAaWkwgc7iACEYOmoRA24nxcp7I4DwHhH4e2gTE
BTRW09t4i2Ukj8Ta5kEID+SnKin1In72iVNGE3YlSslS5VfEsqyqGILE3lp4pR/7
dQe+CeI2y6HqtdGteCCKpjS1H9ajKkVYnTkCV67B+b/i3L+9n/F85dIABeER4pEw
aAUhGSwaSIcIC1ogcqhIivBWgDKtmzcqfMADCmK2MTiJmjpwTiKV73sXA+chM2Fc
PB+V398BpLSi29NK0Y2ddNM/9PY8X1yMNBXcBPvsjTQl7TbDpTZ9ZT7tVP9I6qSK
9rjDGnONoxc0k4QtI/H5VlmMC/h4qFHVvaD0nV9NlFIER5SXGLX6v5db0slVjwfQ
CAxJJ82gFe0pLt/4QL/431iLc89VgrhB1CB9Kp7hU16guC0ef9AtN19zTP5tZMbj
oeglg2tCadfOl2IunLZnInhdHMv6jmcWfBYkp1ljJB2qhb/21XULZdK464FV0X8F
I4omfJzIiCkZHZQFp5Y1V1CkGu5Nmp8wLKVpqgvdRsmWf1dJ9ZyxhmuF67JKCasK
13uSzJUCQcK5nGhOAtHzCvo1KTnwxy+T8DohAykqLtZjOZSd45jMo4kW2sAGbrR0
Ri/Is78amq68Ar6wAbfjq61Sm/Kxg0KyLbfiUdl7LeAPMMhcqgHks3e1o7BK+7FH
KqMsmrp0GFgA7IDkJBKTG+OKmj103R8WraDYEIB9IkQRACFOMD9ogP6l9Y+a7UeU
PD5/IUBVOKYKU2QTMWDJsiRpFHTzSjrnBcwG6GXrX0CTurxHAVQQUnjcrzq17GDM
L6a0jwoN5TpJm9ZOZiiIHU25ag9ohiFA0tgGaxwWOh/clRuplrnWxNEWIQqOJY2R
2IgjZ/u+BGNvpx2D8aNv4JAYksHZzdiaspZ9nGVycT6cFyWPLho/H64DO62TLygn
i+Kli72+U2xx5GEa0ET0uyz2mmZRabMl619wf3l5gpg/jiUWWw+uL12+af2F2yzO
VWgYTK5Dyv7oTJQRtivFSS/CENHUWJJKg/CswwSX6ZrEaCZRwbkXHeC/+/aOoBIW
FQaFmWie4kCWdCNdN2KwYo8XljVT53qEHb6iJA68oVuZRZZaJ1ASzN4u1SsoZjFQ
hNIUSVli5nn7jqRdYW+SdT3oq0MGnaxU/4mPApaa9FV5nCUNYFB9I/iclNrJlZzB
gNS+NUnEelI/cdiPmsg3ZPOE7VaP2IIPb8oifSpdNCivlRZ5lEJaZt1qTcEkuAVf
ZxMo3NKYgD9+IYAeos+pIMlqyGbIKaH93mynbPz98SJm4G52ClOgtI8Md/KQich8
LN+C4emz/EyIFETMmorGJDG077oXFN2QL8H16tNueCY1shTkMsx+xn8AVjAcZIRJ
KM7Yj5Dnuv5jbmiPkNGQy2330hDrb/+nJ+aUuJqMNYa/pFvHgIWRavHNr5+UeY4+
iULvzvFLbH0e4A2i7nySgxJGWG8uHIycSvU056wJO1u0g1hHseJUJf67FeivDiPJ
dFjTkmIogaz/KZzzNk4we/b/ziL/repXUV6KrSI4bK2D7mTQJWPJukiPXErtN6gc
//jBP89+rCIdAj6RaTKWoh/UqaxLjX/hf+D5wnfID2GNUDGOEMlPOXxYBDCsNG9Q
2uBH31z+Rxtx0CZDw35DC6Gz3rlUkT42DGqkxYDSS1QLr+RfSpnx+QaoW2+ZUNDh
JdI7tNIxS4CWDA/1kZlYrVf1ohhTcMiWF67wW9/zv3q878R2PohR2jCCSoeHIWAF
X+BxM2DPyLVISiCJtAHLXNuTUzf59ew+wpNWNfirAOpjqlayALO+5H9CzWy+rlJG
5Pw+wzdSRbfWbAAKC5N1N2RdgkJ1CBLEhb5pXWWyrSy5W8tab+37L5sGT/jb4j9g
dJA47eZSqpoi++Q7cTrpOk8CWJy6wkhQbFR1pi6a9/MjO5Aju89ySER25GoIlcp5
AqnBNIODaz0yvUavt3ebh6awzXOM6gMXTsgAgri1ptXBZFl6kb2WGq0pnIiRPlSl
808O5gRFXOkZ4xMQdwz+76d/NcEd5Atr2hYgSRyptBVYbqBH3lgtZk8M9IVsPPBX
ZAxk6IJ17PUL2DRZ+FOLaNRFlrAPWFa7iesUMH1JLMZ/L+leTKntQYm4FPovP/Qu
z6cMG17+4OUsZHmgUNFmwCNZHqe1nXSQrMyMJKnyiGJNhImE/MCfBg9ScajkQM8/
gTjyUbrIIF7/hMwfU3UbPcpSFwd0Kem9iW32EzWvHAOjWm9G2Obq5RzFvHbJp3Uf
4F1JbLCDUyU342NBuNAwfnYeuYFhtRQpimgbZz0vse3K/Uuo+oO2DTj8fF8AeYn/
g9fZBjSLqusQgIUyCRIHnbZqmD3oNQ0aCCPMdtsZEXHKa/aJ/Yesjyz76xXlXvEP
YiBY83h4xWs/5DLoufHio/qID7jYpI8cMY2QklYqNWkrTf6HQvobMp02eBVV+DIQ
qpZUTf0vXdFjD5iceuF8Z+Lq32j0OElm6GiXhGcIlwzD//ZCBDVFexMEMEZgYIkK
eRuooEr+wJujoBvCq+3T3EQGOBCLiVmOxwCkj5ZZrOVzFe1arWb3tHkqn0ppIJYy
kRCi2tGo8lpmlXqByyVWHoGUudgWMymduKb6Aq2p/FDLBgW94JeGWpam8weNRM1A
2qnxONL9X8jQ/K4iLjzInbNGj1DUu1D+OBiHj8UtDR5FL8UYK4Wt3Rl7h0tvm7zh
kImP1F3UhDNYTcsqh1fpAgN/lsHnULvFa6vcTWZ2CEJdbnSSu0NfZS2i0dK+gPsF
N8oxwaiqDs/bI7Pqwd3sBKzJYvn4GWeu7ePUITsfiREaHgHkNokYI9VWp246p4Oy
xbLFGMl68nozzIFV/CGUX/mdJ/uZnsgbBHi6fQKFI4uC7bB0yoTvojDSXCcHVsD5
okjoSMJjIo3d3WePACTxmsOkcTSTI0nMpy0isY82yJawUMEs0sHbMHTYK4bLz9zn
iKxIEeuZiYiMmaZWuq6V7E/8LvXI5I4uxcLhUARLMQOkCSOPhuteNW9rVK65bJb/
ZeKEqUFzKS30N+mhdLKeUe0LVz8Dj2zMxWiM0ZV7Y5ZkYjCIWwzgja3WxBVHnOqW
BXmfAVFaNZ0blJs99ZxVJFFPliLubGXzaxGhwIoGBkPDOEQgnscVFngEqnhqoUv2
OU1XgWYMqj/Oby9TAR/gGxDsuvXVe9ymL9PQJ2V8PNeVO2Vn9cP5Ayt+H5sSxePp
T1gDS08Dwsoo8oPliRSnUSCkH1bl32JCH2kt+DaHvzjgTJrnbT8PCH15gwl3TiMv
8K/f/xktx0TLQuYpVAM4mn89Zq2yQBeh+h1oDbz9A1RaLob1S3z45SZFmVOEWxI7
IuWvg8c8fhfOZ1JAccahd3DDOTg0IYlCAi7nJENOzEZpnIHIsJeHocrNjHMrPekW
cwfb6BzQppdIGylEjRTonnzyJC4H+POhfngkrHOoJ5Lp1iL0xR6hY7ymuHhyHjv2
3cpY0kWAzNCFNtC2RVX/IAcD24wAWIsy6yEzbADLlshjY504CkXxuTSaxK1OLc1M
TbV/YnD6Qb3ljhyjW5Aqj8RHyRNM4BXyMOIgpAZV25vw36JIdfn4+kU7cQgaoDbt
xLpAKHmv/sYhnIS9XlohMAKjUKG+847ii28lmkMqRffKOzz80GFrfo6nI7u3P4sx
bRPn/cnEVAJ0hFLfk7HJgrhtuCXlKXyJYmtuMx7aKpylW5X3iDBekXRv/9AAOEWY
1fU3IWvFbTWjlOVKGNF9RiB6pK9Q7SMMzWPSTqUSgdF2rt+vWV5POp+oGNqp7jXZ
psddd22BkP2e2/3nWFlSp4l97UrTHCOrVYTuceZaoVt+iqlPaeqFR90+c2hwj3vp
IMg9umw9ioeEwbUaPNn7O8CDsD4VFFXjMmcVZf7bSq0BHpRtCg2s+pt/XSzzrqwr
dhSXX0iXKN0ep2SlBFBLGPFY0Qk2zTBIhcO5SCIoaJ8pib8KkN9/Yp4BqWWjaxD0
bwfI5KPESzk4dG21ICJxuV+G+R2BOU8DMNgTcpOR9vufNM7rO1n7AJVNuaV9oINF
w9vMJf9QMwZJK4H8GQI4EpkMcdQrIRbTk84q8uM5vbje4+MLmxjoLGt9slJhuZql
5kGSHJFPkqUUIfV527CMhiAy3+4T/wT1VuedCbl0JjlGrEHU6Pj/nHZpRla8xXMc
KBT6WmleqTaILP6JIb8vvwJ+EL435jAPkv1VXWiCu9uCOFYEGoQT88DgRt7u+hZ5
e6QcTLcl25mgwjFFxnAqQDHOjSGN0n5DqcrO0lVwK3Wyv9+sunep2BIhsVxEC57w
ylPALMUkPL9YlDk2DBy2IexcwHRn91jJhFa8orHR0uJZlqBtaXKlsuWwZQWWXWz3
mpwP30cMTfWcyZdlbRxarc6DkdZtigASxtktdB2j1wBZibo9VD58o2a22H+KgSpO
00+VfJdfr4yWrkUtXeROoMHfA0e1dCgFmyLFjeA4mc03nD5p7jgYZOmTjsNa8hW9
1NSPihTUgoFSQgT4e/KqzVQ29aUCg/fXA7tUUDEVrVYy2tBAy9/YSMHt0XaSRKve
TR7419hIcHY/YUJ80uLsvImueaC65K0Zp3yoYuZ00mgliRkDx7lvyuCSbC6gdtVB
IOp3aQtqyCqDsAymbK66ynWaQjcmO5xWx4rg09WDqI8C/+Z6oIK+U7QZgiDMw0qo
NNvwua38cCitLEOTy8oPRFUTHdU9amlfAWuXjnV/MXXVaMhlMlnZDTA1B7e9y/u0
doYqMvaPge1nz4rVLpqo6LsJDIxnXoom8dw7RwhAC/RhwFwljbOJvYQvbFacDG9e
VvOq2ont3MgmmxxHUornmlwo3laBVOT9DF63Kw27zm6NMGJfIFKH/bI7S2TnV0AG
pc/llFN3Oc6aCNrnK3kqHLQCyUbCHdsufbs7fAqnAEmn4ZGdsvbXUwofiJmEGhET
1pu/rGUlZuWqvBhfB3tZytOljd2xqPgC4UmHldI0VPn3gvzXE8WD/DzATsz4DWct
Qx3niFciW6xuRZ2URqL+S/rvGRzxLrWdxDL5YGQbdqNGuYxuYgHa1sHGkznrV+d8
GXvy3uqGDi+lgFGJPiPHuMGaIuDW06XScgu0vjK1gMGMCiAFFaIfvYDuxAl+3P2T
zrCVt2soLuWk8shscztCXnOrhjW5kPA/hrsa017c44Ah5Vl05dnUwOfZz9nPEYJm
Evz/eLcQm4VhIkhvtMzqDYm3eHGuyRy96LoDwGtX3mNjNNv7KpfshcHivI8zD8T3
LzUDDFvucKBIyaCk6VoybqHbIR+LiS7CmtZBJHnRRxQxv1FccRR6UL8Ae7BY5H45
vp8ZNSPD4wI8x3RuQYEthAi6RyM1rYvN190SrPsc/RZpOO+ZUrHJEvQgcB75BrjU
mdC4OM4yoeYPyOr0Q1bZ2/JoIHYv1k9vJv2u7jMd/t8IOa6aP3daRs5u1dmoi0BG
Y8VvqHDNhfSlvBXs9eL6JLw4GXz6QQ1QJWwrkOK55GRzQ7/McFBzhKlNY7g1D5Ja
8DqviL6FLM/94NzgMbHcZj8sYpsT1WX5kZtrhdIgMLjPhmuhWJRjh/cVpP70L7NN
XBmdyIb8tmqMjkXzL/8ybAKK+MXc223CuBib5sWr5OJ7GwuzGFwuSKMIIYYRPAlL
dlN9duArnUJxPGs7OO4ZRc7r1Wl0lP/sPr3A1nNsMJxnSVuj/lmlFIJCcKPLCvnG
XBNCzS3gPlRQyhD+fMCzEN4dtF1kusYn8oDYsM14d8lcOEHGXYeN3Q0s7WUm3Zxc
UmgGxKlJ9rnuy+eVDB1xwU56Sy9hziE4QLkJKJa5kG2E6SWupxxQd5IPt4qYg9JQ
oqjrHEUOWES+k2vuLmgEY6N35eHpXuOWyZD7h/bV6YprbGJv0GafrjiG4xXxOVaG
78n5NgI7y442wY7vLSbI+ZwOS6XdGbY9B05zrxYc/D8JCOeVcpe/OACt6w3qC/cp
+wmZcGcrx6EeQfnqw8NTk5pwUwR80m6oYt+D/QaC2MdoTUSMdR/9yucZhnkAPWjV
mwfiqh2vc0LwWpN9rwfZfQDwcuGCz+Nym+ftfyhh6IV6RPxoI0cRpsp5tIB26hdV
V8xfmSSxo32Y5pOAUgdMaU4VySziAOOCCiizBgPjHH3svAKp6MKJvP1p0fL2x0fw
wgVXUwprUtCstAQvPJlOgzfzsUxn+lych+oeffrK4vFqfr3UM4TJ1Uj14Lfd0THc
Jp76oxSNCDxZ0b/7FYIR0aIRTrbl8s+bdtch6vpG5IQqIM6GFkBU+fE2KaoiHL/1
GVkUGrB96xraLam5SE6F/Gr13VCD5PHPXPm+royT3w2Fr+fVnQ+7Xc6+ndWQlZDX
QIC+5ecbkFZfPpEP2k9bcJ2kV9OH+gh0uITWMwjHBLSW24MnQblJhbAx94Mq6Lmf
061WmvZR5zEf+hsnAUYesfb7HMG0Ylz4QEIWkI5UGQZQDMQUcqyi2fN7zWrjcMxv
RCgnWSnRTfu+VbZ84ZtQKcNkdlUOyhtLKm9qBVpZvwzljuwQduJl2glvVK6dENrE
++dpZYyoAhxtiNdNnQvyhd4MlPcWtZe/vseA40ZjlTGTLBccPwNmlR02l1V6qtkM
fQb+EMcvULeg58sxq97Doeeaur0Hs/G+pRUlpYVrNXl/36WIKtvoEp8xPammckfe
ELBERyYSNZEgCpkDxPngrxNTaR3wgHffuetzPtzWyZkrpZO4YYYkaGFE3HI5Omwi
BRq3xikSBq69CrDYNJj3JAesmjpn7IMVcd0bCxfzsxVSs2z2qypV7W0GC7aYiz2T
OkOBsQL74wHXD9qyuDlHGFQscsjJLrs5nN5uuu7QZGynvukpFkf+8eiSecpiXAbq
m1sUDgkdWsisz5t2LNUrkcwkPo52XSj/8giuHauJWCAUE2Tn2uA84PAHsGXDIxqH
Tu12NlQ9MGg+91ZlAHA+KtFSV5jmgt0wi93PP3Rbkbc4ks+0uI6opwAgWG+9Lza2
Hkbn9nHovEAcZS+tLk9IC0ac2SxeuMUSwxN+Kx/sGsFE8w7ScN4iU/T/Ni7roIm4
bB3uF8MhHPY8SAXJHeB5r7caL7E5Y8Kjz70kje5EpT4pIZG9WNsXbnKeQg2PRjWo
lJzLYzKzselG4wvmPU0SQbmbe51+1zd1pZKAqZfvU90Uc/bOJ+/p0mYrwPbosYWe
yoDCqefGORNj2/QDEkvr05HrP+9IBMUXFfzdtJjx51Y764bUiqECnEgHfGvDPdiE
DnccL2HDMZnK8O4MQzUj/cw9dhbBmk5qfUJD4yTF84TEYr5fRv53CpmC4JkpOkPS
3Ugmoh+9FVb1xqqSlsjOb4NZkKVEMIgRDY73FQ+fqpcmptZn3wAEwPnTPQj2S+QC
Pmx1dRxr4HI/LCRqOhZMGjAi8Ovejb8QTcmvmsiSrT0fcEDUqK5z3ZIMAB9QBHPc
uA4NOSR3mCtFLtrgvy8cmrUiqm8Cd2+TZVKwXM5hr4TTJQygTF44v4AU5Ptsgbvj
OStsRBPckvGKMKLZUpHNgsXZ6XcLvM+d7Q42ZYnhlAH/224+g4fvn5yRPo4pcI5a
IIHsYiTxpnHWINPxFvTNrMBBpVgE173blJrWs41CCiYGNyUxznynCuHWm0ZiUDZ/
i9KYmuMC6xQnZGYFeup5C/JOU37H5NcsuiE53tlrk4vYFJyiwSL1Lc++tef7955n
ixFY23BiK+OUSpXmER5SRWLFBg9jnMrg30mQJawBCP1i32DIvrL4fmzawxDIOiAx
8Y1pQgLx+9JbZGNs+8jKmylwXK19XqxcdKBUEDtbhHmRL6bR19GInKbrI8roAih+
Zm8VLubeitzeCLkD/2JkIe2kHzTyt9WrhkxiyQmr81QcUNw0tw+zWE9yXFjMoCfC
ENYzBDQ9sI1vuzAzfdL2/sgoFcebWvhdTXxNtunPj4FxbAlXOcxtK1/oxibhxL4U
Ae5ndAZHdpT1PL+OQKNYCnHswSsqcfmYkwULyetLs3L8u2lbi1ETtrhTwkjd3r29
s9iO+wm5HTgW66Dn9GE+iJG+ZEUntMQk/LMiodkNtL/gZp+Yo85ZV/T7roLlPIAU
ID+/uUGnxTcSy2HVZnn6UsKS9+j1hzSPUk3mUDA961gfxaaDHvVw3QEFPAGuum3v
O7RDPinzdBE9XCFD5LWS0zjweFoGCK7H7zYxVbUlMFCpy4HB58qkwPXbP0YZGizy
+s1AkN+6bm8yUXcJehswT4aDQBN7/gLtc2/L1rCUI/wpxBc7QZ7jTxeQuxDKAa3X
DxYwbHRMZvBv6HpSGD9pW4JcmzC+aXHMJiwBvqvK+g6QVcOungIwMqXwu46PS1KD
MFu5vgG+CaFMjIMUjQ1ULeb57fxYypZF+dznORXQt7ro/xYphW0SOrjuq4tN4v9F
dRfY/wVWzSVfEALnTSNV1+I/JOZHo8wk0oQi8c2NEUBWZ4T4he2Xd/rRjglbM/U6
wQ8eW0Uqmb+N6Ipg1/l7OvEAIuBqrYEPSl5SDm/fhFz9K05JlhB3L3+1i2E9DgvK
WsAmQn2CfWi33IFTF5uBogkKOA0l4a4MISyUCTae2rtPuVlBYjxboDvCH7Kd6tAH
Qn6eZdiSB5g6Rjhc1SJpMiraeWqogZMBFPmouE6/eaUxyE8mffPFqo1z4SCr3NEG
b/i3jvOdgXwqDrQwEvVO9IVZzswqpmf695D2t+hoz21LisPwZfHWBjCL1E0JKVcy
s8Hrc/pgWWHPhyWYFlGvKWv9qTG68X4cHAf19gHw7zZkAsSDXaZBKDAl3xzXrsFL
jzkGo2nUz4mvHguuPQ+yUUB0iwxTe7pSsJpnWyHWimQJA4aqLYtQz9uTEUN4GvDV
j5lpl+f1BCQ9ELwnDOPVSgoZiEnB8RMFrsjBv1ZZwvXSSDHdq+XfssjIU1yN0pm2
jLjmX+CTAWxTXunLANrEZL3kOcnpay54dPNatHYJB3pj/wedS7UwqO8Gvdwc3y51
QiChHzBhMYii1GltEzxiR1YJ8Fu0wALlJZAy2/3pekZTUySHH5vM0ac31AJzzGIS
PnN6iGa3tUFMpg28PJe/l3J4gWb0yCv0dvUmdMAe5y7kNcED3kAOi7fOCLpgjK8G
ktMwEEr250kq8FOj0GZxOYChZmbxWaCXZF+Ui7ebhA3+NsSmXsmAcApK6uIZyp0B
quYz3NMdHEcEJz9Nd0/BMgRF4hfEP861ln2emYhOB2DEMaXGiGA3rgycATawkGo/
+O3Q/BHv8JzV14mHFqSTj8eP2ZggU0SaDSedrD08WsbELPyLeJynIouEycuJJvLb
Ut3Apo2U2DcKBet/pecEaD0E4g/E/i7IV2uIX13e6WBOJjYbctUBq/KK++w43OWh
V/m4SGM9DEg/r9oS4jy+9FYzHYYY0K9Kz2XBpcz3uLYeJvsHeAEB0NE7tWdUKdee
iilOf/Ulzgi9SeJGleJbR5firUln676U9YI9D44kX8QfVhfYp/p3rcgVnz7cDo0W
TC705fAQ2/9MbC3iFAxtirxd6GcMnOR7cSCqswkTYG224Wfq+AlEZSxsuQc1Yc0O
Q98oVXsjE1zRsPbWWLRUgGCK3L+fGixp2ugsjA3UaWPA0ug/fMM6JqrDX4rmCCG7
fjtIN9tyD4Lb4Lt7f+ob15Hq6erux2F7gRZW32DJ/c53UMOsQsZBv5V9cWrQxbO1
qaRuHWpaKZ7og4VLjIajymKYlwnV8wtwd3vUV1Wpbn4p/gDtgKeXKuUYokzpcbiS
jvyJHYruQE8q0hwXjsZG7uCZpIOPCNOFuq+O/Oha8q0gbzIZ8Jzx4MCY/v6cIR7e
ThyxbSttwQmPZZJWMJ4h1IQVQofZKys5HfA0g+fGSQ9iZ2vxJRF+POV0v3Rmyfmr
4ChRRYQFy1lJoNL7J4Z5uVNM3KB+hS6HMPERRf77yhxnCmq3Ov5dA7r3rhZToY35
TkHTJTkraNzYUeVPHoGqZw68/hKSgE6Y3g5l0ObUGud5BMrlsNGE6wP0Z2s0T1wR
UiRc3REpTHk8SsJS4iecYtjuEloynmrRU2CRhuTd7irKHyvpJHGHeHBe4Lt7Qrpm
iFzZoJ/OCTQKiR39pRorsiN8NDvjXX1vR4/6DehNFqV8iJhQsrA2aCLSNpwDdmmL
/5lNreIG3hpTXDSLDx+On2JB3fVpDl/26aHl/On1oPHhziesBjTUy5aQ/fAM0yXO
h46cir30KrzKCmAeg52S+Jupbv9yo8nrKgr9iDKD74ymouz5jEqE9RcRJ9G+uTyp
ipJA8qSVOa282XDrb4D8h9Vs1SXjJA5XJyGyHhrROS/ZzAUQy8KXh3RfC+jdQAZk
lp/KyxG0uK0eJcPBjE1HXBKFqb9Ms83qV0IVKivRisGQHErYuIMf9SUyjPEsbH3J
r1rFi3lo9msjg6RgbV4N10bt3rxaS41NsxpfB4+1Hl4yq7cyIJDBiakaC1Nvo/h1
PzA5h7zA87wwpIALno1dlTVzY++/kjgEdbWa1SrMulgLVm2Jvo3k7WXxS9wQBj4Q
yxJXdV7B45eYQwARCiLi13XtEiIeMf8OikLSOUOP7KIVnKBNhQOOIpLrY/Wnsbms
7UKqJYf8wRbEBWtRoGbrYGbbesZylwlsOVe5k+T5FN1zHB+LL8AkYllMJDhhLI+8
6n9JnYQrIXNK4kzsQ0acKXAlTm94MlGzC/bf7IlN8HBKuJ8GGuuoccyr8tHfmNO4
l3Ms9N8Zj4jSQQ8AWuMndiATVrosWJAYN7t2C1C/vMMkRmQ4SvdMgnJHfCUUTvxu
8LohSQ2tSrDlsmNJ2olnoY12eeX39s5zKXB32VtcFftw5Ul28GcJDYWDPMD63Uvl
+L4pL2FqaimpPWmePB2XDuzgYNbbOhsRHGpop7R3iQx59FPg49o/2QMt2uKT70sz
spZg+3QNsqLx9+N5jZglKQWNngZNUSLpnIHrn3rNDJACVCMxOLBQ2GLb/j9+BcwB
pRw8cuXr5S+ftXO+xEAfZYcwtLLDMM6/Wm5uceJLV99PNvx9c9sA1ruQrGCjgLVO
nDKplXNInRIVdSpKdhchZjH4Pz9Xn1vGUK/I3O/tQ1cSJp38whudKOVzKBRtIKmC
QcNFLD80OFdzH5SQlyVHrlNRZwOfTBP0QRlQpCH4GtbHvSVZGnXgZpyHYaN88HoG
EFdzffgSipFvXq/dtEhHDiPbMRX9eTt0TsmllNgfZbVbOW6/nlAC8y0Hx6jl9Vxe
G8ufsUMLJnXirwKaz5KQ+QZiFlB91S/ZswXReHGPTzdh9g0L5SYICf0LWGkkQgf2
ftmB5qHHfPBD/GtO2Ihz6grBWYNugiWhZO4pN79drTr/6L/UhJ0TiSM+Idy77J/m
LjgSElG0/nz9EX4DQX/ZG741/dOTD3tnvkrOmC56XH2XjQvvWt0TB22wPpS4VuLz
aWB5klF+Ia7poQABbCrupbiNShaZpR6JfloxpMNoYsjyKhojSDCpLpPJWeiXHruk
03QXwoBVStT5suclSsXwDwbG83RN0EgKwa1QJl+KyiJDn0mp6Bo8lNG/NElNOEaV
jWofOwLRxPwu0651YfOR3J3twv0Ne5g4LTqXo9+Og0pQwdb+23F4gFzKy4L3cKyo
9a4VMzyaOkUshsRfI8uiCws9Eo8LTLxZc9w3SI0kUqRjiMZ5HHpYnJKZrANy1/+S
WJP+gd0veec/txgjs3owIPil1UyF7EAYeEh3QHIksAjcuKQT9uocCktO8A2Ry3Sv
dkzl+uibMMwO6vAnUIYrMujFelS1maVMOMK3BPXqfNJvmvdk1gLlGcEHJ1yPUS8S
KH1kjJCGlGAg+79Xxqe5oZnIBzAtTNID/mIKEX4blq73ukkFengm5Yuf4glAQLYX
GK9akWXKf+H793CfFiQWQGr8//pGJ+rb3NrMTa1agLtZB2yyroMOH9Z9lmk0ip6k
4OaF4uyhNrUHQghks1cBwn1K12EljQLPLCy5EAthry4WPmnVjyPxuDyFscXay5Mp
TPps959XWK245K3mBmiZm7nffEh1OmRHvqSjIdmSO/bVS5fUzxecSUy9U0AqbcmZ
53yjuSxn7fmry6P2m5df3cxlTw4DDyen5U4h1MkhCgL4Z5+yaHTExvfmeYeUHWaY
C8NOWuukZUJFgrdLGe+a0MnzyGP6m9ID80PvlOQtQx2/WCNA+oiPwGPcov4SgTuS
XL1dcwUga9Tea/D2vOLa6G0hip+nijv4hvaCPDV+ycdESImMK+6eBMar8aunKzw4
zTiLy8M3IoSFjhOmLfa1akMdpPk7Vb89Fc1f8QhGM4bl7h6npd2dd13Qk4156t61
FkTq725ZoiuXeJP5tMBrcA45i1cVi6CeKVgmjme46h0YB+a6e6WAbAlhWlLKNh9U
j1K1eR3qC8g4qIUVYfNnUfjvD41HQ48MrR3VucCz6/U84Q8uRFjFFDvqMArL1+sn
6tgVOAXfToNqMijud5mWSOCFTGfAoIf1D4B1Qfr2hJve1cHsJylgZsUXJ7+SEvrj
fF8KrECbKfKzzmiaiK+pxYAZhnEQPm29sQ69A1pogTRDaqHE0o7497jeyC3t2qGX
/GxL9lm1KRc3uk3cz0OXwOlcNRZp6L87StxmDow1bgkVSnxyFQRaflFNdnKW53aW
3cU7C+ZS+/JosyE88DW0RUJaBD6Xrd3JTa+cBEtEzXtxCr3CiUKwZc6vQwYFizaT
HE0AtQZ0Ob50gMOEam3fJCZbt303qYq1R9Y6LIQWxLtjTfBqvM3VCLs7HjuPepCV
aZuO48oNpbkDOKNsqg+rp5rU8nOusl+p1aX+kc03tqXJ1keAIF4S2WYOt2bU387N
tHsE0MWZpPjZhZlgcipB49UBs8XEuNLx9SgVbsCCZa5NW3sX+CXK0tuk2x8AWiMp
D1V+/YdFnUqfONfhvY5HnfgqrIiEH5fL34NDhSXeWy/AwFCYWTa/z8/J2oQNY2d3
YInfR1+MNcNg4bdpew7x8M+7cc9oW0/cq3/I3DBo15sl96aFYYvb55wln9aYiUCp
bzPeA5jdiwpUEaxIVA8XNJ9VPZ6iaHeEsjgCYHHfhD9hXdWSWvP1RGhkLItQi4a6
DAjY9+07eqvlg+DaHdfeBL9tOToIsv0B6zSuoiGgHaU+tnlUZT9LP4WTIqDO8wzx
tFsZKEyX+c0th9ozsAgrtGGTa61HOJXor2b3BG5jo0uiREoizcEktlMpl8mN/sai
gpzRHOlZtnnEK4HaVTA/TD97hIv81p0aRZvJIQFPEAqoiwxBc88ZEf+06c6vxjO4
LXx6EJAsDer5juZO5S1awh4cKKIlaVHkBk5ZTQW9p1aXjJWpmv7nHkfGngfWRcxK
1WfEeWecl0Zt+QIVKZEyqG5WsOkfxUEn68o0oBwGL8zwGGpDSQPknrljPzGG3D0d
Ev0pcHDhq/XmfNAzGXzutJsj1z1Sb57406BNKXFK7ao0w0LrILutOUMDJBAJtHfd
lRSYbqHdJCtBRuaUk+GNkWleD7J8B/C7zvDET5cg/EJ17l5hTYWPeKNQ3XyoDOi5
n8dTNvJSvXp+ftFBCHuWwN/nBduXjyjm4TiPMI7htfgdgrSoX7a0vfMz3I9B8nfA
uLhDsD8WlTDOFJeBznGmdVLLLGMxTUre1rHpietXHImS3MXUWspX4R9Ehh/jifuo
wQAxXP9HF+fipoZ8VMsjzRrmkfp7gDRVCt0mIImC9iWOq86jdUdsJCp8IzGhrFwO
r7z0Jp8uOlZJUrqQ/mROm73dD3RPJQFs2rwjXurdZZ+fsDjkeUmX9LjkSyYitkMh
7ch8V3xZOgXpZhpjQMOk+742y9PVjjUAmCcQPAZnjfgoc61HScRvKwV4UmNOLiIR
PWwa9HyZj3rRc7mMvkEYdxs0N9eegNDLMESCuIrNA84KQPqbM6CTvOz6HyYW9Ch6
UEuyPb0norOAtbCWvC6M/95e0mcrSfsoOGa3H65ZD/npFulcceFPevRpdE1H1EAJ
GaegI/H2/uF99kpA4rFq42ItHe3QPe+hj7IlJkILqniKvnlyTiAw8eE3fDbJO9M4
tRBzvEK5oZxB7qZATkuGeoATtPfhdgnqWfdck4W3CPC2rGoe9ZgLzUwtCxHZCKK9
C9J0+BWZM1tpSRL8mHn45s47ILuzTyLUr/+4g+xWpnpV5+AMBL7Qjrr58tORx0sM
otC55eaZzKB5G/iYVUAn6Kmah61Fybw2KhcvbCx6+lPYDpttJRBHM18Uf5WMTyVA
NAwyo81thM8Nc2i4g/eT99xWoF8AvZTqYZ2s4qMHYCE7iNRAd4U7ietzE0kg/CiO
vuYMYVOBcP9BdUgZ3gDRsvpjsDmz5HZRuFewjpmNwIGLwCc2OW8mlk8hCMMXuAYR
XcyuhmfAFXRBkMml7vQjP/V17vlc/G8QhF/rd48Sixfg9jEEUSiBtE/249Vgrek/
+TdvKvsfn5ZylcVqpZD0CkAkNfDT+274ko1EQ6NEUtRuUYyxHIrfJsrm2cmsSRNp
wfemWgz8nZZkW7NLL3j+oGAxG0ZqnoYn0EGT9Ad2MOkzzUEYD9HlOqQjs6Sav+JT
BBVPZN3cdum4maPVS8XfXl12slHPMxLXg0jKszlRa8mY96CWLG/sdIsXdyeFKLSq
qy3KkQbKVn4bNN6p6Qq8hkVW6086zTpNabeLeihNyqgIRD4eKNxAW+PJE5qjkWik
CkAZsGEey55X7iyaFveX0xbRQUADde5/qTE+YkrCbLeHQZ1raDcRwmtdDLnfa6cY
6EBQcGPjal2IrJrkMF7fdjCUpBJh4QDfTVWMisR5TD9fdC8MRmCO2KchOAa+iWCy
XYmUwyfy2E9y8cXXL+bQDt+DwmmTZ8lIAU+KqGkhUXjd0tgZ5dZ3BOBQvzxMD1x/
JlxWSkDUKXjJGlbU8C8+8T+3eliEFkO6kDN7WkbN3v5jJLMC+OXAtI+PIu8I3GEh
tgnuXz2MTILUQes5/7CeFMc9T5cqg4g/2Tnx6FSoYAmRjvb6yJ4MLpGmR7/b1RCo
YC4c8ehzp/Yri+lzDyscpnJuQpMBKZKDlHpUAw1FxOxLaOA2gydoHLv4etVJ4LNC
m2DEsY98/1ZDPKnE7JsiNMOPSklSkXwIgbm9vzZo3/43LGZHH07sVb8/TqkWEz2X
1/VfTGOVV246IkB9cdUd1KGN51syw/5m4NuvVLvEMBJbCmWYnSHJ6QV9lESlJq12
qJGjHGRdEaEoXTG2UalU87E/PZEoAh7inOsZt1bSE2KGDQZNVhwyzUoCnSEmgTuK
lA9k+tqd+6MDU5dc0BINiPLLFqt88D5VYVpjcqjAJQ8HzuCqcYxG6/jQ8QHEw1jP
fbMXXZ9mNfHQblUcpWP4kU1M+QwmkcTjC1vPNd/5UzD/FFeVJLcGBikUK3G28hBO
eei8oaj3VKDtX0j2+A+hnLgD5DbwmPz4DVC3Oy/S7/wyFKsY5Il8WAN+/8rFAh29
kKMTCurZ+GdhYNUs6IcOXphKvIlnlRNsngQszzXSZBNwDjfxz649eQBl7ajZF81W
8k7GYzValdHgsTYJmzSKhfqG0BNDcBBu6bcLnsXGw/1J5ybPz8nx5H+c8mPxS142
TMa5UTVj2/hJ+3fSd/8DcSfDtWgHnEXIRJdRD3UNAeqkrkigJrx5wVq1NPuEiNB0
XmNINEUN4bTyX2GBGg2WhDLj46g6gBgorXJMUkJ3Unw0/EnqnmEpplIA9G5KyFKS
QvKfXchzwsZc4lZNpRIs9eSQ681cvsv1l+oaPFV/+ASorNckEtQCWaBe7S0wdJWc
EK43VuoVQ7frcjnXRZzi1uE1qL1gu3B7EHLWIUxfZk23ALtPkzFw5xb+h7RPvILj
Oemj/MVYs1fSQNhj/jvMSr0LnB7G7n5jRfHOnOzSpH0rN9/gvH/KkLTxM7YL+dB9
KL7dUyTt4uYHqqtYHXRVHh4EJ2czOFWWSJUxZPpIDKJu4RQ/yKgKptaqzX5ho28M
So14s+v6e0IpGOpRqRiloVOJqvykEN0NBPz2Z6WSHSGOzKyQEkbotOFecelZ+j+E
zRRrJxlUYnzN6oBu5r3CkKUDyYK3li7O07+WL6AeayK7++jOR7Jz3AM0ps8cNKIh
XMbkIvF8ue+L/3PHMHKQdOoPE0lMygVwrqBb0uXHYSE7UUsKEU5fUatovcEjLJ6j
j7UX0jKvI8Hur2SXrZXQ7Y18+pveGgNH84BKbFiHS2IdpeCjiQe4RLfYJHmDPH+O
jPF6xj+mSRGkTSeutHvaLr6Qo/Q/uJrh1/UDzL95igSwocNZXAX/z9rkivdnqHMP
ajpe9/FTNbvRTmu+Rw8yNYufAdwB7V2nschqugvipMmlSOKinIlnMc1Zy5p3+PZc
uYKbXEa14Xh1bSSDAG5G0tOeLMkXdDkdBkTIOjPOq3Cmu6raxeSm+dkwa0Jq0sDf
X8iCPNqEyNABQu+sMDSsY2pn9+G/apbfdfAHNjgwfCtTTh6kHNUhmNNC+Ip5fVjC
fVB2UNms77fn2bjC2Ehllrfid214+Rjbki4dGzq2el0cGDetdDzmAwjk3HaVR/Gk
rnoFa/9MVFh6WvFd+Vy/7mgcV7JuBeNaItymbVu04UAKW8qi0ZIISAWTL0I8lNrk
hk+rncAHnkowUWdDMKRcMDhNYn4tx3FYl8HW6JH4aKDOBVPSm1ryOvnSxaMnW0Nj
HQpYKhqXV9mol4KzrF9RP0VwlkWZHVt5J4aoaji3Hx+I7B1LzEu8pBIVYG5Lwj2o
kFtYqB3aKbpf4SvHphDWr6mcBGFRtKounKJrFArhqklVET/KxSaUgeIijTZgr7mB
Eo2Tc+lD03GdS6KkCo1s7HsdA3P0H2tmw2IkUW2ea/ZdbQhwpgcTW/JhONZzSKET
2qnuSXua6STd5Mn/Voguap1CROFCA7+mqZt5h5HnIm4/kz1prmPnF/CYVOKxWDiD
7G9FU9rtHNA/Si997YwCLzbr8iqfosPo1qH5JXGKJ+Ch8mF1AzX3ug1vTIVKP7kl
I4O7LZr1GS3x+1ZyWYWkpUPflCNfNsMj3bBMEqa9mZNjk7wIZ/cVh0ajvZBtFOTY
7MUSqsTwgjPHCGmIb4gNKq7ijADTf8Qr8GtVJcOll7UhHD1HHOeG9pCFfbFUjG/1
9041vnRAQKPB69oG71HIGIPHxXakJLFvVBywJdiW4disLvNV3ITps7t+d/ce7gbT
5FkN6hsnhZ8VcBPBqwv+VoLPh54/GzmHM8D1QOgg5qfV7rxhSjd0av1PJY2u/skE
JkLMo0Y8Yf2b8p7nNIdVXyZhtMFHZ8SAQJSceSeYE5BIVL/+o0rvV5Gk4ePuA81z
H23DFljD8u8DpIVnjvr2JVUTyIH7SnH+wH4m7QnEBFVz/99EcodUqZkkX+B8z8lu
AAgdjDLDMHqmVrUaLsVCpcN/gLri1xBRV4Zca1BP7BT33zyQ7hLCfmc5bRfmPZuB
dY0ggFmed8zhYlpC2juDB1qExKkjrjEK8N7lifM9bIDyALEoIcQOyrWojggm1ziv
y2ITMzbDl6b8ZvF7Wdj5eADZXg/+7Wu/bavIhFijRFbkK/lJuTPAhDbFXmQ1iTuQ
aGN+kBrklA+iYMti96rY1OOsaLlV4zXxwbPEuZEeqS8bIPTYRIeINn2RVFTTcdV6
ntAFBZSlBmjHcnPuINAjXiGxPL+p0YyfM19+q6AUb1f2F0XKe7CTiKl1mL3yVRme
k8EvmZbM9bw8S+5WXH7PqbpqXsIfdl1bNz3hwWmM4nqNT3VBoh55oH8rjM2O74gK
DmrW27bAkFT0ykfPTKouH8+txokMd2RVZx7aDDbUYVauT0IH/CQicJYNKNLcvBTu
OrQ6GGuZT5khU1HwRTsdY0z70QbWbGytA9ULftTCocxz3Zv23ufdM/M0HG6cIQrE
H8OyJUYsgCd3GdkqznhzeN/yyHPe+nEdTPqWdU1LDcr8759G0DPH4vDBDZxgD3PG
KPRESQyuXUAak4lmDJl3zhTI1iHy2SZXPf3dAcOY4mLho81LDVuZFxuoVV2KFPfe
fhKY74X7oeds9/swYkuV4pUMwjaISD7N6ZD08M7nJGKiZ5iicpEWITS+nZGTbykg
2UDZM1DXCYivTsLpMi/7T110SBsDsxt7nMl8WM8k6fpXRi8Ux0//qreOJu5up3VS
lPDlrqNysmlh18tDFIYqCNSDvDFA2B3gU4+p7ABpi753PV/LRcT+96xLxtre37Q/
xgIC8thONJloXrGWQ0BEf5EH9VOw3I4Eu3Yman/a43jhK2eTR14KQtIb9S3XABDX
rHrIL61R93SGDrN6NepnytlDgm1t4tnDEYyTsWcxyLhS5Dk21G5vMvb4+jA8UOWk
lA9aaqvcY2vCUU/2IBe+QF3In+kjd9/DwdEkdBd0TT6xpbRZEB2WhHwalHVWMc4g
dj9xc1xT4ngSc8uM7IcHXFGHTU+A4NvJSdy1zqowhmtwfAF1ZIjJPa1hfo2WOuHL
uogdhfAl/6p2d7oa7BLtY53QzhCm3BbcPZb/8Dcs/EIozXM++iVdtoiTY4ZZ25iH
hYrx4zzXyjSjHCj+AiNYO9JkP+tj5qXIHTIyA5FFz5HOzJdJCRXOalF+CK4hAuaP
m3rq8eCvwK9xpPHptrDjNBp8vkFPwHP9k5p3jR0szlXHZjmgr/N1dNngDjTgmlpi
5gqju9li0gE+zxy1ryDHmRtCynuTD70DmpwQquG+bFKpDhHqjIZKHyFlv2e4EHd7
jifiombrluAt6eJhHt9euLZOLk6qIlPS8IvvE3CQqIn/+pMa0vpNgTgS66zsnfrY
SretbYDd1Cd7sUJs0+kjD+m14S1100HfUzi7FvtjFJQwyjN02NiZ/VUxcHCltuUG
dR08q8F1KJ8Vn8AIf0q7GsDJ2CLiTZ53IcTUyVo9Ba92gbvAr2OG6VJXTiH9iA0E
jcN3pyooe3N9ObPkSaC4+gn0IEkBFNiMUv81gR6XDm8NZJftkOiWzJFErM55sdVn
MobP7dWVoRynbIBlY+Di5GZcLV8erG9O1axWc3Bi1DgeiG25272JzT8H4NuZMC4T
lJ4PBo83VENqriTNwPIv+/6DV44JEBQfNq3JujU0vWji5vZxg/ehve3tlHmk2RGT
dHm8wnhkPMn29jAZwp9U5OYQG8Opq4MadkrPyL/C/W5ZQbL/3QzaWoGHsjjqkG1F
Yh9e4OCzKe+vbRAYG2A4IesesP+9R8k+IlP09S4ENlsGvLW3A5wpNwrTMwYyxbr6
lNV/QqAgBmdccwgBxkFh8FCLSna5ehztf6QI9jxq92y5HgtR659OyWCmMVpR/CmH
PiK9KVqKJTKEMEnObC8BUAhPEMQm0icc2wxZtmzKEJgCvmKGMLU1lyB5LDJKNymo
jA+luL5XhJVS1vqH02YYVJpm6K/N5JgtiNpl76jKaXBGWg7hWDQx5tynbRvKPUyZ
0VsW8Ox8DzVxdjlZxljUF98CTQFs+KZGvh8vRl6Ug/Q1p6cTvey8lcIw4TPSL2Zg
t+zAOw8jGH8i7H/sZDkVpIH7vT1zHylnsiXiajpf12xvspyK8WFZX6N1hc3lFYzD
nP0UyC6BN9xX8dasgdlpe0x9UmrSygyYr0lhMZ0iBYM3b1t40aCTgPciqMI1TwxY
Nk0OLypFq9mI8IfkOwsVIcP6dR09BSwcGRvs/OGRk4iXbEP/oVdGBxunkC8QuFF+
CmzYZZrXVztmgoKmTiCEN6eGUH0lKVD5M/1Z0plijpRhnF6TFbA1NN+3P7vBsNlM
iUguvFNAGnYfULOuUyrbwzdc8cJLe8hOCuwL4b4uGio31sJTpB2bBzb016b3sbSW
NokEl+VSNFH30lCwd0ahP41J7zkb5/oPt0O5z4moIdNikuDbvetJ5Kt3CkTr7pMN
/hyaGV90/ev/SNJUyoixJ0keROvIYEeX5mupP6LO1DCX7Usj1UMhk6H9bMPKrZqw
YbN1qt5cDsgPLQNwJN+sYG3IkEq8aEa6XPpVUHlw1rzW1D00BWGgAgqEc+u7o4Bt
4bC/17HIIeBhcKj9bt+KZVqvEbLNO5wV4cp69d4TSHg9OtKfJAfInvPbVhSU7tXE
ANT90maJwUNUSo2XJ3+iVxYcRUkmWrKwJvgjGVbryjRTBKP8DpQuRlDjd4lRNuvc
aTF2CieV0myJGm12vIY5c0GC3hxXUN6qgohu+brvxj1Tk76k2btlmHi7r0+ONI0u
Rwdy/soM72tmg8uyBN5gG9OQCOkzYwqn7PHIna93KRMxzN7H3ky6T21QNfRBJ6Nb
Me+M5MWoesvazlyAuevGwH8okD8OWxk1Mz7shoZzLcKSUJQer+D9HqBh+41bKElf
cSoRVw1eDe3ZM7tRo18//4gPo0XSx9KRU2haZ1PYrBA5xNbvtXdLxGRbgbjKadMw
OEjdQfDMEOaeSHxoBHIC7qDFrcT/pkggWXJSLDJK7im+7DBXhVHfT/1cfMwRjvzB
VvC60Til17qy8BOt+B2l3Dev/VdYLUUCbrl8aV4ICq/yeTJaUDXze4KtVdHGtgR5
KY95AD+5wrz1zjKDH2rPebVqLvOck19P2S4gEjNlFVViWC1zL+A3FK1hOryN71jH
AUlAL1wXFZmQVjWTMPcVJWijCzJ7ZRG7y8xUqm+TbsqFR89Uydjw4KY5R7zli3ZW
H78Qqe4kmt3JaesjDp/jSbwDvRrl3U4PSt/B33ksVOikAjQhd8ye2CGOrY6flBIY
03Nipzqvkqh6o52ckzNpiPPRL/Hv15uU72iGQT+ImWJSI7XvAd/AMJKeTUk3zQhK
KO4wQQE1/s+atQ6ZCpTjZxWivSJFLDDzHl7ljqoegVY8hdNQVvdCHnJC79TSvc/N
BUlGXh3IJls2LFKMYKsdOSLT+abCIqN7qqP9r59o8g6I1xT8YTKiwbw08+2FomjE
l60GZEVEEZuFkMTGhJaX+i4v/216LQBYb+1RZf0HjdKVzklYYxJfCy7xF1QmkqV6
br5QlYG9IdIRVa1j6ob/ZoGukGlOsQpk54eSlu5xhy5QAoayv28rzhlECWrRtffP
Ex1KM2nF26KP9HqAcNt96bB9znNoZsulMC8lYqCXxqiLOirMwRFdOychWEH+Z1ZX
TpCEXfrIVIqCtFvhB6KTkiywbydE2DWOltiRMaSgN89dsDeqjGrCjzOr/G09BAMm
gVBxW+BHrWCARIFnSZITfP4AjqBJGJjTBvAah6lR4c4lthnykB8BZ+uXu+UoepfL
0votmCu0g0dvevyTYcgEMX/o6QrX0VdzC/TxzMF55lJ4vxrkhRP83bNltJSJ6bfj
RLoAKwY2usX9UX4v4kFMYfaP4xBh2UgZkHzmVgOG4idkFdSqnMCDx6TrKoSCZEcF
bur5L5IFZpH4ZALP9ucuJlAKDTrI0Wt8DGFYnSXZEdgfyb7mfM73T4WdpxZyd3Sx
IUCIXK12/ieVNquuwOXFiojZFPbiDnmTkGScifYxKrvzzopmRAgbPLbbRmIuFi8o
iFn00VBRl68P/GWTW+faqY1+R69QR0oJsvqm04KZAXnYlaYqh/sxvf6spW9O47F7
SSzEVXtmfPpunVOFC5npaaOHGm3Y14sr/6ki/rMAVJq39iZbV2b3wBl/nXv3cmRK
n5KXHyxi6xQEUo0L/xTIeJzavY9jOAZgy03qDNlsIAdmC63DwDF/dUfBe1sDRTiA
gklAOSidfsYnYbWeoi/bsa86P5H7dpyZ/xdlx7kqdk6RyKiNdB1W9SFT75PSrdeB
r5wQTNkgOqgjtMxRhRtOR7xMwx/2BMvRVZPD5Ie3oFcLcPpm7KUrD5cTRAG8NBlu
DIzFlGxD3H+PMSF7ywQCbK+wGbDC1NSMtHEzIpx2ke4A3BJ3YtDQ6VMTSLG0Op9T
vdR69Qxh9wYbGtqtTv4ZkWYJ/WsZrR3TqWk3Engu52tf0gV9fPruFWjp0nOELFMA
kEbgEFTVjI1Q/6bTb3YBj+Q1k4WzEnMrCsQgoUIesu4+KaHVhxUL3fCo5+IuujMc
d4AVjiiHmoLl8XHD0jL2bIz42spwm7/3PxvvSK3TUTInv5jm2mOn6KCogR2gGT2S
NkS51RLlsHbJm3OmU2I4NokgS+rMaGX0U34agx8rmATH0wF5p38d8a8MGvSRh8RZ
qI438JVw2xIyVK+C1iDZRfOBmumzmPwKaESrEqcDiyqtC1XuFSdz8HcdLmn4Cnr/
Skfiaw198jI40sc0VQY2GGO3DiFQ3GaxuFg46nS0DaiyOikZYIvJw268zQghAlrd
CRl2QSeRHEFpkihg91V93V8riLbU0oEGgY7YcEM+ZYeaN4LArO5opn90GdPTPDcn
d2qlW8NF3N+rTbbmU4tiDFlc492g6KKgXVqPuXyLgrwQ5mIsnrxDHFucVVOZp3tt
lAxqLJY+Ji5UenTIq+DY+VF4/+TAQqDjNsu5XNqsVeehhxIFKh4LjObMr7kmEMH2
bMksvreC8Gr7+3IkoO+Mk+0cg1s021PIXhYkXzWzJudKlEfkCd1BNfoBc1K2wqcM
x/pDwrtVpf75q2RxlV2h6T4qGnp3u56r6uHls1kBI+ASQIfSIKca+5THeOVj7Z4s
OLhB1vTFXKNn3woKP/BELtmh99RsVjf/qE9GISk1ORV8Jj7cZOXTnI1D4gsoudCQ
uPHg0QhUJFHITXCq03F8muR+7vkxy1qPcKzdfBFJTcoW4Gt7G76EZcj6k2L1RooJ
nHLTss61/Mk1HE6ouylC4+Wg9z1zwQrPOolxGZ4fBEHWuVypWHjOOVdkxVROUg3p
SbA3oqrL2AjztMcEmhWx1tZ7E2mB6P9aX/eLBeZc7zKM23d++3fWbyuAU+dh6LSY
ZE/DMviR2TtQMhoCYy4s5lKO106wmqWHO5gLAHpLs4Gecwyomd4uAa2knzbd1d+/
N0ug0Fylts/hafFnVkUWFUVkM6BntGXFyzomVIy4+ICuivHSdWvY15JrfDZzVVBp
Rth42wYz2ketr8RdOZjVF8GBD//S0/YM4WPFdegckqoixTlInJWxEVm8Q0qU77tR
lcfKHwfOxGu0YG2GAVUn87KHPCZp38cX/zLxrJFrouCxcx0qxv/KBol0i37MJvAX
s6DVQlfoNm3r285BmBV6oG0HjDQOw9BfoKfsyRL+5k2Rk1J+M26amZZKCDJ24OPA
vpK2pXJHsZN7tMFNe0gIER5ELrk4IJMKkREBrMsw95r7vdkPo+BHZTYyKkh+yJBA
I9pP4sxauAwTvGO1O5/FNBeAC7NBgr/dPbxHaK8sNIOXBLlm16ucHc7zASQ4p2HW
L7GJXGtcEJNipiudSICcpOeeyG7wpl+zNucwQ1MSYWEwZ8QPq34rI/cK6x1hEqz8
fH3w/nzrZzn8m+MKCBRhkPyTcitVylFufTxuueAnXDQoYP7h8RtZFNTMXOgkbwJD
i3+NgBie5d0YxqEdZSVm29B3ga1PZSVqb5nnoQT7k/S5Tb8RemmO1J6Blp0Uf/9Z
HbjHQxPnREY15vDwKOEcDwFEcuBD+4juHB+4hnSUIFsyLXYCB6jp9TN2ouzZaUXl
Bn9j3tn54AVx6hX+8r3hU5cEg+H7rGd+D2ke0uY+kSQPGsLfOfEVziK6NnfQTm4Z
EKGvWrfFpnxGcG5pcpWLsbyVrVHaREyhG7XxNGuODPCieQ29L/lM4NyLSG/1mr5y
XtOY6DQc91p1tf7hJwRIc31UqDf/reps0yZluFiT/7yH5I/XI6hb6lzXK8NhT+iO
N3wdHSQU1MGakWvAlI+Y4d5DQaJfIQQ2NthCUNQhG6IiKRs3uHiVALC65n7UDhpc
S544MwC8ISVu1LBZJ097YZQ1b3a3koCFlzPoFtpuy1FNPVLN52ymtGzAYE6BwmhH
9GV+/Uv2ZlTON4a6iCQE6h+o0LLx3xbXvEb0krBIGCKarcrbP6swSTrVJgA2RKfW
4ijV/SlnCFkQPIyJQMipzpct2ThB9WdrrETtMNYakS97+FYDVauFyb9ShJg4EI8O
0/qorgiO9IHToya/rjcvFys4relOn/HDPE0X3GXebadxbpKSErsx+dXVjhvW6Q6x
u+2dsTRwaD1aUQ9x/eC6OuKQupQR8gJs9vOFApZ4genC3E3ZjGq6kU4NqgoUyQDK
6vhi84W8dgRB8kCiyl+ax/LVL4t9Cqqt1Fgf6gwJvO3Q43FCI1xO0AFUJR7BGLV0
LvQOL7RRFMdLS7TwOPV+c3lWKCGtQxHFiDmol5H+Eu2VVkVQYdC277NFE6KvNRPm
L6La8mTGxDIZSf7PK1EVtrzS45pHqr0jdqMszrsagP5G71Tev/80840ni6FbRiEX
derTKUKwiZvj3KzPc2Wtdxh3QanGlXqYZDxt/FNY6ca7j08D0j2X1TPkVIIBIG2E
vRIBXvqgm8B08FIJL+KGNi780fd96MCRQjtiDTe4m89JuzPlyCaw/m8B8IXjy3a8
92q8HtCJdmxoJiD+bJy/0EK7U2myU0VEevu/YbONoKfnZ1zwHtxhZlmzVN4SRmEF
nqkjuSjnK4vimBjDmZLEcoxq5d5mqJdEWgopkof6HwGz/0Cft0E1Wp7SiLpzynh3
FjYRQbK49GFi4gRBvx0AQnJEpPUdniTFww2ZHr2ss0OdHgkSE+rQlHUUa22V3Pu/
/DbCV25oLtuxShCfPVfgrxlSkCP9nbz6ku6MVG8tzEvSsHqIfZEcF+53lWUSQ6Es
LfMXh+VmMW7Er4hQfPVaRKRJ1vkZChxNH1X19tvEDhd/mLS+LbDaLpRWuknywLuF
aDrAzqeqwaE6rnobTzvdpHHn/nyflEJdM6mvJ0BzxKHEPC9Q9e+KA0db+WdhN4Mh
YDEBkdsMzV310Y03yEtFjN7LTDCqdPZ4JIA/7WittxhkLugsixvlOFKOiLVQlgLW
T6f+m7eXnSlfbNOQcJlTPNEA7Y2wT9ajaqhH9aCN2Ngiu8aqz+Pbgv6LYDfXTUUj
coIZw/LktiKqqBtKGOOrlRw9/utD/VHaxHQM8/kbu1HdO3h7iU3V5FoYDsh9kGCZ
Z3UftGoEuFHRxgdHY9S0a50hb/f9gu57VwZpng2YQH4NLCiC66bAlyH8HH2w8BMk
a+7KsQjtQzOfD5nW6XTn0bbvtZ8ohQLDdStpwOIQHSfnWLzs1YPl0jYNsXLyssGS
RC/+8SJfr8vT22FuRMk00DttWPXQ0O3J5M7/d8a43m15nocEV0WI4xhBYq3xqNo5
saAUgPp/UT9Eh6qg/WVxMwfk7jD+mHl3HtGc4Rm/fspMpnZsUBE/xq+HPE4+PC8D
xoNBZVOmBGxSVp5flZmj+1MBfmMX0M8YjWEr6phA58Q97QbJH2ou/E8AJZMVcnsh
cMrjT10NMdXlrb2WlubN1pTqaTS/7r/Rlf7AzNlK7xJAuN8BJZoe7oce5PpTvs9n
ayajuHVsQBfyKTleX2wykvmEAApvE9ZMSd2EcUi1XS1Ez6V0QpawO731RQpyFDO/
QN/giD4Le2S4+wenpMbzKi+KZIEvu28hDz9XAnhpxPwlOwS3uxdcJj6w7J67lH6q
YgjNN2tkDCL0MF2/SovcTBLiVJVrl5oGrMmmKZ4i3RwLEIHQ0BHiWOPPe5A6ki0M
expocmtn3wnRBPoHo5grkUyMi0uzQa37pShH20WY8t+Di60eaboY7ShtFwTkdmx+
4YZD8315VT0oPHzIEoiEsPBnuVfQh1O1hhrt3NyoIShxYFncnL66OLn/KYmZdXae
MOtUnOURPxFL7JLyTv3p047Go1JxrtHC19yMUCCTE8LA0/bnFjogoZeRTJ6mX6Cg
eOVz/FsY8PV9hv8fbeieiDISOw4QrUENbFKJJ1wMPL90XwTRCySSPw2cCYlQxVJK
3xXkj/2PmhdwD+Pslv5KyjLy1cN9oea+fcT1H2gKNpVdQFAur3czuF0ogODci5Zy
xjI3cfCUTf0M049vJl5TwoCLvEfwOREt7Ttv+9YCDqJWgkqGAEb4rtyvYGZqzjKM
n+mLUx8QVNSeqlEmo/qNIbUsP7PdPDBWc43nBOOUDOE6kzEAJlo/KzDWGLOJF0kj
sYK4bVPKRJ+cPSWKZ3zBDBagP05NkB5pFxRs1zluSnHmsE5f5lrZrcdXzX2MQdAi
pMxi6XCnoO4/L7Dz+ATTir9vrE6itaP1EqUrcTpQm9r0bDAmKGko305/lMxJG6S+
YdUgQ7fg2+QLy6ehRsCQSEenWISfVcpwplNaTymwGxAcs+guLScySb+lcAENcoY6
3gW7ATzfONMuFaaj43z0OMLdFj/AF447rgTDIyrRMFz/9M/yZagn6BNR4HuIwdeY
Zv+jSNRlonxipZV28TLPeg00QdJ5cP1bKqwxGtmuATAx6RIKKLBUjWRG45hzYbIf
c6IJalO+pQ9XzFd3PRyy+fpjM5ogE1IiapoEYoI2CT5JtA4Z19SIBPSFBuVvaoOM
eXY1OZQywzrAkzvSk1y5/DlAEBqKGrh3u3/GiFP9/DMoLERyNs+ryOZxm/BtAFm2
owdBCATNrX+cu502o7MPosQKnbg8hKZHKDrCce5JVVMFkKCqjAD5G5zu6DY+BOEC
fAS2LJHA8fFU6+HqfE1oqjqMJeDfy5FzofXKhFjGXcob8DVHpIyyKX9jLtNEQhq3
jxScFi0apFs7jAeAf7cHaKgkvakVIBg5sZYCu1R3BE3NDs0whsFDlR5U5TW8IXGN
E2cYXL7CI+8Hpb6TPSF+jSraCELDde44s01LiBB/v7Cc10bBmNdgWq8IrGaAx8y+
g1VHXPrMy75kLpK81DwgOFgjnZy03X4vYEnisgbMD2o+siOaAuFAygP+MSGUJMiP
FlRuBRJJQ0YNespFCVOcroxE7TEXz2iZEvn/M6zM4DFbHKweAExLwLb/o2WXpilK
ZDb4mGqyibrGKjOyqIOUmBxL2+kQIHIzKe7y6pmIOF5DuHf//3MEdxauqClDmi+1
Ra5y1FQZlPEy2a3lUfXCUR09XKo16JZGhmZedD92bO2qHdGWn5E46Elti+o8HvH7
H2nvggHc2KLOUOhlXC9LqXgK8E8lt9/vCLp+mVnGuYIG5EGLJ9gRceyneKqXeEuk
Mu9IQGr+OgueYAS6rIbedJL+fTXNp76yQzzO//4s9pj0B8w6dYCToO+bg3lHjI4a
Jq+GPWneC11++Yqv8WPh09JxL7JAB4hGln3rQwAEeY2S4OgMo/GNAHWP7gL62D6g
0POxqX91ugP+m3yFOhogIZNdO1dpz48My+VZgvpSuvy9swL2XjzO8HkhMkkRFtuD
UfhNEbEOILu6mB3HQ82TKR5iRaOqRwKPv+ch8FWjKGvvK8WwvPrJArgXelsyqSY4
LW251Z3f59Aq42yIRIolFodOgMay77RisUuNJsdCS92Ltyrx1WCZM1YDru6AGlNJ
0cjs5OoxvSHc3ugiArGhwiIdizqgcFjW7siLh41AXkH8ikjcJbJPnCwV8CU+zzkA
DU817JYJ99S0Vpdfsw8WqLxboEqedO9av2N5apGbe8cPYUFq4S2ofSub8Moj+HSr
TzShqbdqtCTq6eVYgmHikUReHNow5MrOyzxIZtTIJnMtSXNtsA4faFex/ay6wLHg
QQoKjyi4QFKmS+7loEeyclM7uiYoR0qEAfX/+FNzF7bApl7aTZfngRabU21vNjOD
yWlVcFBXGsSqt2K4QYDNHhInjJbqmAB9v54J0vcEM7o4J+HYtzQa6THTgiOD7N3L
lXxF1ZPsdP4L9eAv5FjUJLzoo+xH/0ToEfsGD10Nd6Ed9jR7rpG+8jMKSad1ACIr
jHtw8avHfhdw2LXaUuWgNGi3w1NOD/IkQwy80+1ja18iqap81yE9f4x1I34dG//R
CcCNfuJgVf4cFa+QlpcGSS5murst/zzgOCm/yCiJdXViIQnEn1nSZSNwEthTAZhY
Lh2+Lsh7E4NvAikIJmmHsZk4UNruBFb6u63KbMOKArDADv/6E7z4E2wyfxnf+EqA
Rv0ffW42W2BkeEGDNz23UeqhcCTq5HAOk4kIKrAieMb3TrE/Fb0vtt8JSqP2HbIs
U5xpZB80qSypji8ZOMGeUYe544pZKhyXfJmH9mrIiFOD1Ioui07Va15c2zagsf2A
7o9Bj3hnTEpLl3gKYoFCffyyXZOQAscs7g7H39v/eyL21f4IvngRYuFu7YAeM1kD
L8+ejaNsn6CKCkwitAtiV6A5OE64ninuXbszpgUdRxOx8Hud2b5UL9p9LtiZcUvW
zvthERNOAGNq20iUwMMP3w5cC/3noZP6NiB3txiXYGY0u40vTVPWJMLD7VNpZi8x
IutXKKqN36y73CXthBuVGTUiPmHEAYie5AEgGOYSel4IDXCr8VLwEyr3rTbnfkIH
6vDB4QfVx9eYKwcV1FOLlUo46sASKfCogu0dBJbMQMisN/Cm6K63SwYCeoJfyRZn
r6MJEHXZG0408pmpMTPmG+EqEEpYVtDvNA5jjsOz9Xw7PSlmx6PkEuRlaKElrail
9TZTI02THAxAgmXXpm/dz5v2fKmNEiVGxo7Ry4I4BSxga8dar9f/wXN5nZ+Irpul
jdCJjRY4qiLq5JJPYJALAMowlI3ozaIcdBrgyHVT/rbItS4tS8CYvP5En42FyTWl
FUQxsPLYkIyHcGjYBfR9DHgT9p5zcC+b7r1dx3vKIMEcSFj6F9xPBhqBUVnSc9oV
HYtwJ3AliEtP4DqLyoE0UOLwO/5iRborKBFCTB/3IfRaQiTJbzk6rmdpf33f909f
HeUlUlBgOKd32NwMj9YyATVnOCDziZNmTUC3NoLnsURCtE3LZCyOS6NE1uVxc+VB
TEyP6We06KVw3N6VODlriIXUdTl/9CuGGnVNaUU99nTjPX5MEAE1ZgS6dO/eXcbS
Kgh5xg49ONMLmOltG9BWz87FvcSiAtVymn5vWCo/GHiagmeuYR1uQkDPtXbVFFOd
q5wUJzcPsWuI/Du1dzYXLtEHSMIUGG/o5FVxMBjTUGG/QtkGAbm9ZCda5Exgp8zh
lxoNiecJt4phldNmYz5hHKWAF5Q9yMDd/SE/azerZlr7J1OfNm2iymJiS+qrxxzb
hC/l8JGfFbDIHMo2d1UqHZ/1vxtpq7iQrHNMwrOQKpbOIGBqzv39qAaJD32L8EQo
M5l98PlciYoTa29vzSlF51ekG4L7i+7/KYyquRER/5KXsVHTYVicosmVUwNr88LP
3JhShBB5DSueSMw4EsW4Rg8GQGrrIRS8mQmpqYdfPLRkzm4gN4u380VTLwPRAYGe
r8Fu22Qajc8vLdGF/vuENo1WMqQhSwC6AkNfs3CnrZpej2zAUEOp4AvaYQj/9Krl
B7mfJWykrci7mOo0VIoBJGodVVUyU6xon/ORvz4x6AQWOuWzaN89wVgoJZzzEzDa
RnvaUqAJjiTSK4THkqaeasqiHOuiFEocBMQ7gj1hCpSeZoreQoFlVsn6wTXu5mVL
plyN5AIe/aiZLUmSRAMf6NSOJsA3CgNCDC9hdwFLSha4g8x8l/ecKisSo18mm7Nh
/i6ZgEPFC1K4EPSkyPNQBSoRpvMMy+01IjuOFtzdRJ2RWwU+HgzBPty3/ajNkAju
jJxhiVq03iL6GxdN3XyDb/hYo6SNSpDuxVuckru2otBKjiVeu8pplAjZ1NILebAV
gLDRcDMuMNjFZT5IJR7x00Db6gIKbJs9px0oQi1rDQa1pQrQxJRu8cF3CAN/FFL8
g28/ch740MEdGmTUVzHtKBFDjeEsfLSf7sCUthstsnJI6QnB3ZXlvOYcn6MpgnLO
89ga/BiaMIY4gnwlYdJz3PEeg17vj3gQ1KDd/FApVr93EwrbD4ZgU6kfr5RUPOHp
yaerQZBLzS6A+i2rqZ4lsUbMMbh5NU7evvdQijsVgVAI3GjZJVLf7C1H7tUh3RZZ
XcCwJ+YdNa5348gHXdEaJ9fgBLFB+yOE9a5t44W8ePPRALDJW61IL2AtN40clfS1
JlRTbmWfNpJdqDiBs+qAnh7tYbgyrZLHnHpWRnLGLhDIoMgfhsdQ03E8u2zL28V3
TwnnWj7RtfODxZ1pgt64H7vLYSg89YBiB2RtyfoKAxGGnmN4juNiJtskho/WQ0f9
L7X1t8nBn2KQW9s1DOwkz5tUX05bmKb4gTB4ehVph9QFB8GXCPOW5nni3T/VElaP
Ob6yoVShUa49f0LCD3pb+AHPPQeqQVY/iuniABul1IF/+9aFACjlb1NVYnqu9k8d
9GXIzJWfsMBhx9YotX80dLi8Icu8mcEdpILX0hROuOi77iewOkJ5vjBJ7ZxtYFeE
7ir7euXwKjwj1H7xzeUFfWYAaOpD4C1Uyp0Q33aBgHim8J+c3R7L6b6DkURECY9V
uC+gT07Hm5LwgbUXqzmOvh6Cbmc+KVAoQL0M6CZfq2EbPtHNkn38yzERZ8abY3HJ
Bte0+f7PfKc73mOVlrSgFiLkKF2F+DPAg45xn/loaTy7ioNZRahkhhIBReMRe8EI
MsM+BTNhP0eEMDjgE0NgHyy8JB5hqr7knmzQ520bYFVsN11T2WlBdPVQS4IL0L0L
rWG1+OT53p00bkIgXeXTpsPtqz6gQK+t/rMzj0OkTFLP4o+DUfwM4M3LbTjIzTwh
pXbxEz9lKu5+eclLCgy4JVoDp9Bw0rJUSnthUEHrOUG9em567/P+9rdi4sUulzZq
BOmFuxwg7shEwJH+obMDBXDmEr4gyd54lv+qcCog6IY2ZPPX5TALGq5P7TaT0lUn
DKm2+aMHYr6WUijkBkTez6Ur8eDIGLUJMxOHc7nD1SU000jwfQeF+6IwBrxdm0sP
Qiyw9rsXQxPc+qk/40lQQIr5JF3LthluV+Xk01U5s4KPflu4vxCH4ew8Xn1wro17
3CAv7YEvRVnEwbxslEyZeTzbIXiBNOWVf6jiql0cCMBsV/2g/BboIruodPDJDDmB
twg6SOfW6kD5lFxArcUc6/5Hml+Ekd22JLz3EYQzBxjXz3tNrN653+991VRBdjUw
U8yYVfYnFS3/M8XrxtL4K7sbqhCku4rCtAYla8HmuGR7GOLRT/pEY4AEqSDnnVqB
XL2qa8tlGm61iT1vAMSr5jYVB830Hm5z9+8NmVnHBdmAkPS6p3lZyX0YitO6JzRW
t9R6prN34s/18nWsf9eRMw7P2Caxww5kMG+wrgGAdDQ273M4fhCA8J/SoZb3uHh6
kOhEMfmvQqQy6kgRDfWfupDNOo+l8kwkk61WffK/ALe1S/OIlLjahgHLtLQtAK0p
7nsayADPGZm5AbQu8KuCpeN4KYxKzerT0/mFH4OGHTS27ks1D3Rnx3U8ZTDOURlR
8hm/a07ZHBlSE9/8hfVjJnE57OAbLFHPlYREu7A+7/MlYjX7U17CgUw2D1tQMSjv
ypxsMHwVYq4uOiXlVvg8uDG3VNpVdltrGGEobsLYJty7HnX24OJ3WFo/wAGfEdXR
QPpuphp8UZLm5y+WGR3yztEBop+v9IPIxytyP+MGlgdwjAYLx+oWKDoZlEzKpgQm
v30UvLktWGGXc6xPQCsLA6BG9Hh9ezOieoKjopJwCI4qpUvE/8dBr1DtJ5M1pIBC
4D1nI+KCDcDtiOdLIJD9YGjRv/70vbNuTMfUK/7YBvlp1/yyJJMrkiEwR8vtK7QB
rnTFIngN8LvQbcjFjyLaVfOAaXyk22orZC0+p+FloK20OV+nyD3b+JBWRR99Xsbh
U7Ie9JFU+pSop6do0aHzVsZkAkzQ4bl4CYYoU4lUYqEGVRpyRkG5IXomU30j2zJF
N/6MP66uELUduI8LHNoYjJ7EtICdrtgDh5v0OUlnmIq31yt/dJFB/wOF+5rIyP3w
vODe4tVZ/H5I+9G84Iqjek32UoxXa0f/Nxfsogr6nOiyR55CkSp8HIZeUk9CfZ2E
ZqLXO/003HBBhR3vgz90Q6FddzFPyH6JXKoxQclTBIU1a8xlkuMk3vlPqxewSCyS
46aCgb4y7LMS1rMyuPaMM42wzU2VKnxEaIzTIK09ACfkxifkmp9uOzYKDcKhmTbI
hzds7QL45afoAbKSSskoH5LW7A11D0rNqLqs6NcOQZzByxhlSbwGGUKGZcLRJ9TF
L1lpmLBNAD2YQPGUyfY02VCLMk+e34Kgbl7pvrI1bDwgq3c9pBydgcqKcB0/7X1y
PQoWtVoHrMYPr/1pz1YfL7NBSYngn0+IeFXmfU/8isG9CM5T1ZPT6iO75LXxDEkp
zPDsgn+3C5Pqd2dVNDllyc0Fze8phN+dnz3ldr4XU5lONCLxiQtWXPVMfwk3oByD
ZtCzaDzJuJitzZMEVC+ERveHWHumtF4WLEvUEhEAVX5DRzfuWpFHPt6hYOH3jY7l
g2sz14+J9U/IfSTmMSXSlzZJ3HvzaZ09X2yK6NKR0Pc9O43yZKkvWHIgy5fefZbe
v+CRhrc3GxIZTeUghIJm2G+Yi/PIpTVplLGz9urU7SJdzWIuSvaI69zNXz9cJ9jW
tt6vnUVstt8xveNMQPFFRmR6SoDz9C/DBPNJRmbgI0JoepicdGStOVOQ7UlD/5+i
nQiZQxCBXnVyGJ1NZuB2z0w2fe34I3aCmzlfV6MVcDzW3DyGxCHpdAwkRW5F9hKT
UprXzA7H5gqWldVeEDNNb/3ydqYvCOerm4O/bn02SHzqyK32sYe2Qv1+GjtFuaQA
LefYekmxSEMef8eJ1wsBvlB74VwX4pTbEK2U8Y42wwWqUMru67b3m2NNGp6HUoGm
OpmN0LC88MC+KsVSRnMEsRDM+sChuBsxBiZeqRf15Mr9Z/RyMDxbaFg0Mdg6S61y
NpRQ6ajpCx3mbphYhQlUw+fraLUTYCrAbXBEMjEUTgglLG5tt6rNjl/3W2KGfzab
274115MoI+/jFN5wrEtdNYk/Yafek/7doAbHwno83zbqZQX+ykd84tjwpcIHa4fI
pQrVedlQU6Z6ARvnbMPi41kvktYXEdVs6ZW7mDyvndhgLlXtaz6oCkRdJ45Gz6hd
UNjFq9NXGbBq+EUjTDiXEOReRXbbPZZPPtgTR0gtDh/gLAeKCztrJnNAhVQwXABq
unudCRzJZrJzoe4u8LsMnzzB9+0u76wCGDhwqGpuqdbZ2UJzbvkmfhOkKT3yatfz
hClajLGU7qmGZIpfNbsbJ/CMgmlfepvrhAmcFkAVSYcICuERTHy7UF3+In0s7uie
caSQahga3K5K2fMqkzfvMGFlYKjzjRHH0SCSFGLllGOnlYo7vbmvW1m0dy6lkF11
vX4nvsxuye39YT4e/IzBq5FJ7Ugk7wD+o1mt17EIKAbe42nJrF2upt52g3VlZK1J
sE9tlqjuPZAWlqchVFlTKWcVonxencKLp7l/OpaJYncwUB3f0WT6/UP1ENhxtgN1
gig0IoOcwi8zESo8uVvyUItgM4JdR8O2oirkIg9wVTxtJeXIzD0B/+iQ6K0Cp1mR
5oy17/LPVGjhSb5K8q2Dh/TO8omH36ey5mtC12tA1VoL3DpYOjO8jjoVMeUXrZws
p16ZYsfa+Sp3Y5fMEHXxXDiwpFrpdwgKUYo1ZI0rWk9mxrpsP+tbWQT1K4+PTyVn
EODgj/F2if1pcbvkatHJILE0op/oCtW6Ju/TZFa2gku4FaZ0ytYjbOJKqUvTvjxG
Wb3AmdRsh2cwQU8AdLOiUhkoyydifxzwNz9D9RK0LgXOOFpVcWXPnvvv+wGkKaAu
6KPOx2Om5ohVhyony9FzyAywG6DRmixlIUQiT1k9MrpqUV23kBbUbiOZQIONV/Ej
e0B9HkckpSvkZYi4J77Uh3H0wSBhLBH9r1MvIWL0vG+Ueiy1s+4jyDJul6kJGKV0
WTPgNAM9QzwSoCJdmFV683K/eA6dRkdUomStoFa+Meq2YoX2mSOvyhjlhCb71vYY
2CPvvJ9tIoMu106gpZ++5hctzhKuOzTx1eBup9ApB2x/a0W8VXL/KQsXZryQXhmW
dpzahxqqsBmBUhIRjODRmMALsOUgsZQAsn5mg5iQ24jx9gbmynV5HsJbVTFlUcWV
mEd2hJ0ntDA/1prlAlguO3EymhbYSnFmspEIcvJ7P+CA1ZAOoXGSnWQtKqYIB43K
7ZkTuUM79tYld7pumbpdlIuvln9Mt3Jtgs+vaLc25nNFeG8MjKVkBny8Gf7yLmlU
kGoV7N/I+08U7/VmWH8VwqylbF4ijUE014tDU8pBuSlDxfrA+HYH8bcKMs9u90bO
xu2t22r3RDzJqBRVhfP50esH3qn8RkLnDeU3TYQVKojSWhAEc1GlTzAhjv15lXKG
9OwrrQzi9JxnOdZVCDGwHXc3POrhe0ceuHB2ywBCmpzyuC7IipqMkE0tFGoA5jbC
xgiWmtrx6VwuM7Eq9u3fssKcLQ61pjII1FPS6kukxP5+tUTEoPobyrL87mg/qvXN
xn3StyTZOacSe7+5XP3lKJviuz+Ay96ROl/JcGMVLTIcTxfHHhsYb0VAtKw3AtpN
j7DLt0K8LHEGjdC7nm5Dz7Xwl3JpXJYkFEeO9vFGzSrpS7/11gsAXm/T2SZaufRr
rre3WKZS8EJfEHejciGWmUxnxyKsfVEEKjJgZgS7dqknZ31FEhlJsknf9YB5N/Va
FOdTN4dk7TtB+Nto5H/OczicG/UrV0ZV66o9zDsXIpBZypEmNvDgLQ+LwQ1CnyJy
XvyZhCt5RfYlfHR9C1cP+DsYUPA/XF8qGTVAQeDRtVPvI7/gFPT0LH+g01ndaZdP
HYXmB7furWx5rZ+ZvQlJYyumTUfkd5lpL0rTpgW5Y9HLzMpr9BtfWg8FJWAe94d+
CtTU0zxh2oHKiHyCOm7wBGjflrVs1c6KEi5r02ncTtuRedlo0eCR2oT7uH6Oy5ea
3tWAVJVbEc6Y8OlKmME/LYFamlys8mKFzwz79XLcSBg2h4AO+L61pjZ3Ruv0dxvj
szhx/9ixitUD+jsTzvep67BinTi84p3Unzn/A1iuzrBQuYVyMeruG28j3jyh4UT1
TfjZuH34RQqSx5wNhGj3uymivJc/r0sUgQsz84GJGhKiE3KSI8+k2quzdPIRx1Cj
EkP99AuzQooUqeKngPI+wpHLMCsUwYC6QVgntWH/j9X8cW6/Olc96/OjVQbvOWgs
OCfMcobbVeqS/eBUsHbmHLIo2HkU484KA1PCCpi9NCADup2mbFJ9LM7d3TjHezpu
L54EXGKRlhb9k5Oa+CbzAN5t0115Ti7ZDK2FDQ/rzJpz/Pg6E6yL2WLallKfGsed
qvuc5EXeMwqV24/PmlLeWXzDkNxdkLKygk4YThxZqXAhGWdhnhveOIsRHz4ogQv0
gYCvnMI4P9V4rfQz1wDawIHSXwqV+91c7H9cyWJ827aHZsWGr1jOzyTRG2NM+pg+
BqCjoGBcMZRqPDUlJZyU8mKytqJ1zLG230+qVIvQiHeC5u7kEJts0ff2eHcwgxEh
c/DWIoXKT4Ri3DT6kyNesbyQDFcowqk9pISVgsFTCGZZ1G+8GIwvy9civ6Gkgvle
l6Lg1zOwUJNEzqUg22Zmw01HgDlYgmkZm8Agwu+Qb0Nuo2y8nVY4kv/RM2CQlvp2
dW4pDQ+Cm4U82SDiPqcm2p0v+NcJrcz++T64gu/mFS12WZo8wAID40nkYu/GM+Nb
/rCHHpSfkJEBeeluQ7Uu+UGQ/bOzYcz2vZD8mw48gu75G65jH9br5z9o9Nb+ltOd
ssNHSG/tq3u4SZRMh6JFjjVmHQ7gyxZYQPt77sd3jVyP5Aaz3oHc9R67iu861u6Q
x7PfZ67Q9m3q4pkulrJn8uN5koAJTPrPxG//StgpQGjm9ckvzHz7vlJEMiTHAg0w
RizLi/t3JbQ73G5STv3nm50Mp3cs/cfil9ttHhihbZ17T5ZBV3xfbV45g5rUbvAA
Ug8THW7vYPlbzolKeQe9dBtoXnZhUj45X+lxEWD0XZr4/3Ee3x1cJfrQ1NpXbINa
LEp2xoVzsrcBAWvi51cGSDCzxKb4EY/8rZV0pJQIChuTBhheU7bgJmyorrvWlX8v
k6JfwT30C3pmdu4DER6+z3Ow+S0pVxCEjuROxQhsulqeGBKEprbUqOjpQ4Tcw1io
TDTw0TxBTfsjUgSc8iJH6YYvrHXUIKKqvV9dT6ZlC5pyx28995q7NwhDI4fdgu7h
fxI2XNEwlSN4YNjKR8oBag/Udt9Y/vMObftGkxs771ybJmge0etnxuIMUH0uvabV
R4498DpQV6lLxSbXqRoZx+XBKjHh9t3w+9HOzTc7Riy8Hppx804toD9w57mZFDnY
gD2ZZpr9WcFdyYxTTrkJs3WxMVlciD+91VukXFTcQb8pI5WTyiLegQjMWOc3QFeq
+uA8uWBStq+Ud+Woc7aCe2eIgi4uP56fgIOCyY1ZmE55XqQFzNynOdU0at64SYBW
l7ukgdqGYVDEBBiJDZh7FaMTnQepwcDYA30LM1JUYGuGo7gZulPGmqD7A967r9HM
DH368IllLtj/DnAr33fsc9GlvBiXa3UmBGK1wlxVx7Cwqm3K/AdMZ7fXAum88w9K
PWMjB5N28wuYFMDoIdFHtF8rVtPJuHWKJmNC9f8DvDPC+czZdQStXImiBN579EEx
11jt498BSdFICBCRMNnwok3QPGJKLpdxGndQMBPaB9x2jRvXOasQqcw1Mcuc/cOh
9FaozkXFK728HRj7T/ljatLPBHkVCdZeTfbuWvHUqpqd0mdpUvuv+bfiWE2CzAeU
q4CnsNz07+ZdoHR/SV1pYmQoEoBls2hrumErOtPuhBciEZhw4F/G5ouXgv74hJeX
cCYPpBjTZ+Kiq2m/busTZS/iktnmeLCMQMfdTIuWHPuIqLFCOC4Vcoz4e3JAGNTD
zheCpa4UNZceIHUHadWwOVPKwDXl2nOUtC6x6YbccVw1ztALIFldfuBEAB0pWdnk
CnWC77UMR8Kg3qy1Li5XAtBWmip/L8QxsH65UTV6S1uV1mFuesDOeHNj+c/oghAI
JG8voTcv6k2CgQOEJ0ob03Op91SKrVXad2tT0AB4Lb/NtVG9dJsOvaIrbVwyoVLP
BM58Dp/yhEELdVMVSw36fhqgOaha1kLjxLqQxhAk3DLMQbt1m8L5ZlaFRy59MlEr
ZChcDZ4ckq2UXmFDVi2mGEsRbMoOmDDv5ReN8daDc6956smVJXG0msLAZTHRV5VE
VYxxY+WVdAzAnQoTWWx6z8LlG7qkeKAd+NekUWQLOPBxCaT2k6zQgT837dAY6u+2
eVZo6bW9qfQjao5Y8xO57Ho/Ij6asLXVPAEC9YNpn+T+ki5eG2RlKAsaiwg6MQAP
QIukJWrjEnjjJ9nga10DvlPCq7Nxd3FXrej2zNzgeWvFrD8xbv6zP/6mmHlBiIZK
5kYamWSVZWb7VjWGtWMq5Y95q/XmtYGEcBHs/ca1B9rLav0CztoCOZi+LHXtDBoO
F/fSYb7jNdTrR9WDlbHKOot+N70GvXsZHu6Yc3Lh+XEna8Wdq5CPNRtB/pgJzVX6
P6MZmlUP4hxCCO9uISTxSRwqZBHQri8EbVwYUD1BdeYLRrz08cuU1UYJpwTzwL40
NP2Dsp5JaCNu28Zibi5HvQNyxaBuLFbdl70Bjtfw0HBFRl/WXsxjpaTiYJCo55r/
0TQmbeDRe47IliY5cluoOZn/TKfrKCPbNDtfUm0VJUdlfbGWfdEcOQo+ks13S1IP
EdXCIgodgSKZF2DiC9dGeDJl7pj4o5mhDnjaB8S6OQD8IrIBQU2KzN+ae8Tup9TY
zvn5TAP14rMGq41jbWcuJYXgX2joLq93vrov8NtPor0sGO6/2pm+VYG5kARY55V7
unfAMP6bTBNzCxHMOhzBa8BablSx//z0IDLEB71vwa/TYZxbq191cyPmyN1Ek50f
vStu7F49obF9SM7Fz9cbXHGnUoe/kUyOTxDk1j1/xKEMPumxMYm/ljmRSa8gzoji
JF/JFtwNUVYm6B2XDg7qunhY9A2F0qABmuNilrCBDD+9DV197fBzHB3VgKPyML0r
Jrc5v5NLpBpJjMRMxLtCS6wTNpBgd7x1A74ahmFf2ANNsvDsT/QmN1jTE7qIHgIZ
6QwBgZFutRO/LsywQjpjRiIdSl1dCd5dWHU4CIi5ubdgq/NyQqxkB3Cn+EW66zwE
6KDdkJQmmjw8la4gjJ75jfaquzt6jLxo+FOQia9FMK0H5XBLifv+wq39xmlQgqQv
QwpUXHNQb957c409Cnk1FxbljtuxQWb26uJkxAea5kmYGJJ8hENPjOKO2jh8jtHu
lWpmFCJPvBnLmne+QeY2E/TDC7hx4H/0EOb75zyhMzTM+LXUl9dAGDqFZhKPX7Sx
uoPFomkCZzfnpSVzm0jw+CU9LyLhPuWO4WVRAvr9IX2EYLsiwWFKpeeZ2D7yIR0H
UW1nXdpafHq8Io6cOtPyBvvBI70jBgGoJMq1BCVMsHVaZs8PCbPHIDPwftp17IPL
/7+LhvR4hpbxn3k4LvZQa4jc+3iN4bn27wBYfAbh3I0WM96r9Ft0Xw0hvfbaqwN6
qMo1lONJsg7QcT9DWvN60Ljm7HKAtop+iDysNP2zZ1SUgPRR1c9Ce+/KPtQzMNHy
k1xyk+YsgfRN30OlQrqBBW9VY2JIRcBxzepbYgt6gVCmoZBY3FP8Zc27nwJ1rkGR
fvZE5vlSDs7tPuug1+WyFWmKgIqKRAvRUTeyIVlDNu43k4HstXFV536s4c3xeiHb
HEGniZnxT8kfBUQNEqbLfqOGEfZ1zZEVCHv7L5EXqX7lEKYNnHMxMQXyT02Jjy9P
YZzE1azMgpwsRpyD5cHhRt+BD4Urrl0v0dTcYojqKdOM1J8oqo7HYxNkioZLrrGs
+nFuIcgBL4jY3/WAtQCQOazmEdsu8mX0BL5i3nYd11t+/YnHtcG9j7G6jnYLCNWu
frcHpg2cEq/scQus/+2TLsFUuwNm5OMzmmQ8hSywvUIIydkX5Bvr/EFsGQ3cdoYK
aUfrLVvhOc7gyrmGtqLn4diYVmmveBsrxmke63ogrLcLMsJxdPFfeE33YMPIv1y8
JrnOGYWSbQJrb6loV0dsSOqS8Is6fQePZLbBZFRr5bnBXpbiUjM1hiCMsRJQ0wPQ
if8f+tMA4lm+0+jpSV9mDiKhNY6tQRfTOs4VDHVUv39+3ZxVk9ROm4YsQTh1XBix
hT3Ima8svbgj0zTsg3U1SUtzebOpX+owkbRpNiaoMZxbopCFxeQnC8XryXjDv1T/
ZJpR2bed7W1VAjnFLll5JbAEWIyAxWv8enPiGt11YfOZCKk9X8zoLUGIPQr3qTo/
iUSq2zHetnMzQ7f47Qs+/KjkwmHCStMm7hDLeVuTC8+ERQwGJNFiWgO4uLyMNVub
AcxaawJvlpY9GlhsSQlBpzN+FjFrlRN/N/75tYIxJMdSgpPsHAQ80h4Jh/KIE/+k
6rirpllgf39F2CCk3AEppplVudmValw1vfMugJZQBkHHwimoWN4nOnUsHZKX85NU
M0WJXjcuTkvS8hns52l0nsLpPj4iE2Q8h2OVo+uo6AufV2kxpO65PoUgRDESmcV9
ja2dnJENVGurx7wRrcGkVYmUeo5Y7hw5+UYDSJSbi8UFQZZYp0joLOt2izzDpLQT
bfxMVuq5zB8wQXsGJT2fpQAlG4cWgfXEp7tN1PEDLhqwcUuy8TOjfKu7EjRCL9CX
dlZtF+xvXpftZNGbMX4MiKdDfj1oLzhXhy/OVxTw4n44UmY4V1hHsI3rXTXpqwIb
ahAknNkW0uaNQZ/GLVeJ2ZCV0MU6hAwkmvprfWyltXzY68EXwwjfclA1l+kPHLtj
p52DN8oPHgBZiXoGYFAyn3LIjuHwTJlvsc6ZbfgXi7/w8enzJUXnOz+mFKIDpwN/
WePAhxfrRVirVmFfIxCIadobnBAQ1iC1fezvfX1r9Op7OTBnWYdUQy3XHIxtz35c
eHmcDD8aQ1ymd6Ihd4G6wtZXyC/8vAPsytv+d8T1aDuWctVcwEtt/vxyP+ZN+LXP
IAA9qn5VRovvz6d8QLYI++DsslnTljLfULmF97CzBjFYLgNEHV78SclLLg+nKz4/
vqWDlUtAPi1wiVsi72rXNE59YGtjcprOYYJUpX2KQFinBloqQcLgAE8JkzW0QBVQ
I85DzE/nSSsth7GNoyAiMr7FfM92VKlhjAvkHWKzwDEha/LiHovV0scmgNqC/ag8
nSxENZ5YRL6GFtKaovr0hMwIRp15KEmPnMpH3rWQi3I3xoNj7/pIPEe/4J4kP9AI
GDvmOCzSckjOpyH1K3XGfddJ9GdEoAfEOaRFMt0lKeJaLOfI55hkjTLOy5vhXajX
98fSGHArKCgjzCC6x3U6XcIz8a0alwQlxgbuZVEgJVaB0lGW9K8L+DNlvRGOt95d
DTQNQMiF7o/nyuvluL0qYCY4/IwQ9mTWju9/N0ApLVTLDqfVlqHNhUNkKnbaDfIY
4BW2VKj7Qm1wQpW7CdTAfujXHPuU3qGYHN+bvQmb4t+EVBr9pnLs1cbKsuEJJf2O
WvAQcC8xEw2DGrGms56OkpoJd4apSieAvyyjF0hXxONQMTa5dyRsfh31PgzVm+5N
0EJYJ1mvh5Q/o9MoJLK6aIOSyMZgmMBvJxMiG6DlfydzC13LLidOvZFbNs7zN0hH
D5FyyT/X9jIa+NUv+LUbXCOIDapnDBf37ZkUZwsBUBzNXkeyxBOYXXqRKQga6TqM
Yx81MiQbcI9WLNIOMRyf4YeglSCeDPZPSacKfyPPXJ5i3lVpBzPX3jdw6N29mr/7
VdShGoQi29iGEe3oD7f+1QTWocLA+rjivI6hWeDem3CMx1BD8D4cl1IE+fY7HRIh
n7YC86v1QXGTbssCvpnKzWPyyiDgAtWzuLLzn3m02+7AiRR/t8N/4QWI/5v6a2l8
/jcXVXbRvbrFwv7O6xjCqfYi68wclHLJJeyTW4XUxCsi0vtIBZ6Z8XoV2NqMaqIX
gNfIsXGd+AE8GXMvCUKhBPc2CYWoEY2s31ZX9RWg14AvBqG8oLa30hX7+U9UPeqX
0Y/52LwCbKE2dbwt6MId+228RWAmLWYDY4aARLMVpOlvriTT661I6xeQuSn3KunC
aqCGZkFf1B2Ea+mZS0am8LlVbu9VH1SJq9v6NSco3+MrRpTFpPe0Q+Wsx96iMgh7
ZrLlEAadK/hygQbu7QOAIMD2XgLvpZRseohKf1xSwtGhmWto6YlZn7pveyyEgSY2
N2/gjJxcPIf3oCKYrYXQMqWYOgBic1rXsam2wdX8BfYI1A9+XCPjV4dmp0aPULcc
g7u+GguKUr0vvLGTtoWgCh5qgtqCfnXZfS4m1PW/fJCM0zjmrxXUnY1+cOsd8EEv
7sxkl4kI7hDGVt2FZi2hgmyN5dox/GHh9Bs43VD8O6/7t1++++3PN3tvTBS+0ObI
1IddulsHRDB6nOwmqthshhVnMHK3cvsxQ1by+6Dbxh75Lx294ilS5Z1javaFmVxJ
Cv98RArySjbozbkkW8FzjY62NUHzCzZvjIWyePZHELVQPYdr6Z6bOUC6lP/nD4ks
iRBDw7zQ7hzjHz54zTbpBv24Uobp5NudUn+Lbe6A0Mg05k9r0wNbyCXHPJFejTe/
xVdkh2zZnMPiVAKAaGDPvSDbq3CS+WprEJNmIr8+BJCRwfNiVpdRjAfyoXTXgM6L
57OP8KSFfiRaJVESLKNrmYn6jbGzhkjxgzGO9YS+zAKobdHgt8BWL1ChA8M575Mh
prqlgQJQFRCGyULlC8g3V/5KhG20dYiWDAlXUj0iIx94nYwMa27EYu12X+Zv8uZK
yD+hkLmobyISFixPvK5y7jq8brftj0nM0VdpGCbH1OSh7IXzc5MP3s1uEhZD6Ub+
0JLJyyVjJXCC7qJKisfKzXhAgg+m+JYSnbJhB/9A4B9gzn8O6Cw5Asuzd8e8uNO3
ZGQwADj+WhkwtEfez5aCraEgIsaYBrIa9BTYpUZ6+PdbAHk9X7UHwRX9yFmBeQyo
ZgQcOUg487rsR4IshlHnt8Aw6CTqA/xVXxuF1A2W7qj0T5wZL1tCwt/ZoQ++QE3Y
Mq9sTqt6NKmVlcq2r3V0AOvZK5ZvaxQ0ALb7FaZO2hVVdMRATMqLYshx6ID4b706
lYBySKdxuyn1abt19IWpOby0NBOhss3zWYKmrhIxCkplSsEyvrkkzSZxyN0/J5Q6
BXKCz0oJlYrTYbhtLsB7yPR4gUETO1Jza5fsm3nyXnhGD8nWyjFp25P33WUhUp0p
g1GbgNZVhTE1rJR1kbpAwgvF+xmcL8bWmWJhy96AAxt7P+06pZEYc94cp0IwtHL6
q+rFHVDct/gfbxpZuhECw+g1ucu2TD81jC4GwkYTnrRr0ugtaabWRZzEy8hVL0Pn
kDwMP9R+nxjRUPmjEyMRZ6pXwxFQCeOePDxIrr3D1ZE4pBXmGJ2JhTwr533rOjTA
YnlNTsXAY2h2+0IRgSFuxrvmi+RRYt0IOuLAwP7W/QkUe/pBlQwOdnnYM9Sf5Q4N
e5XWOTHRJB4Z1f2S1+83aE6ZuEF9oDGeeBgiz5GuTumYqSPcVb7Dga1TAZfAEA/X
3fq4rdPwnJy+YRNKU1jM7+eKDNbnEv6HUndTfCvbVBHPZyJfM/DOHW3hOffXCF7O
YJJD9qtvnFhf9ykcwR4zlSvqdilzXiMagkoxPZH0kJY1duKtLpUVU8aLI9kQgq/+
9jRJARy78s4fu0CWkUZfdeCp3iV6B6BSz61K38962UOmfnSsZvC1T9TNrLr0YMgL
zgsn9IrzqebxnO9ElHiqW9ga3u8md+Fq/AMSCF944L3WK9jlSYnhpaukMn3oyRe0
q/OUbfxGZNMJzXsnXt0ji0bqorG40MqyuTJzAImyB9vI94VI4opMOhxH1xmolhCc
z0YD6pLEdbra/jYYZ3exCThF750T3n0TdpJVB5TNc+M/pu1HvmtDQRzg0LNPaAzU
qqOnG0VxOG5WHEo2Mjr+df1Re4p8qxjFLDzFRmNRX7Pc1xKkErU7f8mi8Vq7qgek
XlQLktz+q5KwUvkp4/iWD2R2ymiEcz32lUyfiW4BYbjyEe5KN/1bJQgBt2QLQ1xN
Usb/NlQzbHfGVSPZcs1qMmK/yrOfUh983yGl2cAS9poYGKECkHLaNdioQHRHu4xb
H//vZUbY5pBZUJFrb+vhig2fa02a9ptORABC9rWWBoVg48+QwZhYm3EgIBdsnB6U
MdH2cwfpZNL3ymJ3WDO0SGuTOaImXZwsYylIn6rD1gSbIS6O8byE1IDYtpj3nl/G
fjvDlQTCQku61hjywzikJE/wj03OUyel/ALc7SrB6pFzr7lrgxPP4WZbzaHiH/KC
vy6ATgqnM3lgBl6ltphy7tPPPfRb+VszlaxG51gotsbicoI/iKpxsbO3+aRTUwXk
4mpznaUL9kMdvnDrMyprzAyBxv27TqCm4EhZVBa7rwWOZEpGqmsjqN5LbNK//xLE
7BlGY4THUf/EpscRmQYJCqiv/clVTy2b/hJ2H9vJtNECgsl7kP8+xJnwJuBB5Hig
09Rit9JWqsziBxQbRspcm5DQn749hyeii38j3c3XdtMCwpAZtwbxRgaclowj7ECO
uZ3Y2r05tupKHAUKPxtdyQ+U836zktsjmhujbY4de/DYQi8P7qmKyUKWI/hpZ00K
qOyyMw1K6kBytvMDVxKq9wx7UywBh87AcIk0mNuwSyeaa+IkIBEtJKCrNQjCbr77
0ms4H+uIwCFwrOaUEGHYvP720cRN+K/CVq2tBaaZoSJYIRwC8w88DK7AGZmDd8j9
oEww76+QVHVpnJAIWmECHZOaUkDTeYEMqkieRiEbpU/ehr/2u9c0WsW5CW+bF+qU
42pNAcOiY5d/PzwgZsZPaY4EArOI/CTBOBxMYt3IgoTBaQDq9L014/DxxP3SQpC9
c5HDVqXCHJaEmhQtL1JoxQLH1pEj3MdaREgZGJbedam4sHaao4S09hv/T1l/8WLT
l8YCBgKnYZuvCIqVct4+5TOy8CF+5UeKuD9dLKeM+vFGzeNmcWzV81HVEsvKo5Lx
3idmebk7xBSpa0Meg4EDOCzV0wUjKlPi+kczMmVmE5wCY6punB2ng6lRafQnkg2Y
1d0YhGECmGQnV0hS7eU0FuRd/12Uqrluqt/9FMz9+RRDrZHh/W9FqLnBjctP9Mfa
Ehw/EQ9BpLaTU3fwA2dFTlveS4Edxo6DG6fNe3Yt7U8wEKGgN1UoLErfqAYDMcx3
Jug4Mvjg//4eP/BRjV3cgXFCf1uuqjguCa69Dnrz1gJnElhMdVjmKZRv2GY7cxEj
tugDAQwpY4gbOCAEgMaBiFSxwltrv335acrE8SrrVpHnyLgQN2k1CSeumNt5m2B3
q9r9ZzaEeO0HumtU4t2UnrlG9eSO8vPa3PuEDDSqOLduafY1XK5vRrj64dV3Zwbl
piJDxngtoyjA7mlj/DBqz0vKyyMBuIMvZ0553MzBke2x2xjcp8WEhnk/jVyqyq1s
OkRiEbdlO0qSqvBDwyo11ENNWQsGs0JR2W2C45IhaeavXJGES+s6Ao2WkYubQk+z
POnjnqlCILXo5K1Ky7la3dCAjtnq731pzzQxO/LOKBLuJGwjKELc/nOg9d+bOp2t
dl0OrnvJLGDg61f81TjcujVl3bQnrBQckhE6gsQ8gH3e1KmmUdquxFM8AFCgQceL
I/sk2ZFI4aydhhnBRtS3w3Swd4KDfjWb66Dwr7xmhAA1MLQapKDqcw/8UepVoPW+
wIahApiSAJ0UQOFFlUsf5C63+70xxhLJNFPLVLgj2Gm2ust0zHeOtDbq0LpbnSpl
vZsb62PiiMqydUlJRHU3/qETxvsMx/ezx2Cg8XlTwMDhNzGsv7BPpKMnzgH3Yei1
2eSbeB8DbEgO7joYP0D45cQx45VHRKofE9kou/MslMBeyvg2BKXtO17HRMKshu3u
qfps0IP9bosmxbpQ8C2onTY6XDjhqyvS/VeXaGiMwkp5oDTw6GdFZLuj3BzZymIv
s1tYZP3oQVAUdREWQSZ6fLEo2b9/+l6Ml1YjRqVRka96nvm0J2dgcZk2GQ5v7RUJ
03ZYm/UqdwazpCWbK+ci2Xrjk9bSI/bKghiEb3r+VIUJNTMWCxyVGneIALxgrrXA
b1uqBFTRi8P+m6pm0cp8X767+LhvxFVYNtMsyq5OugW/qQX98C1QLDjwj3cIh+iM
3NIsEWz74kpDS96sWqEcbhLEr4R2Myneiqsd7BmALH6mzWxfFLlBTFFWsWdNS8ZJ
V4LJkvCiZTtKk6q/EiEDgyPblAfugWM2wHHOBTTsZIzRAub4qbHXwmwE2e10JD0B
w3oBXh3o7UWl+Uzfu2d1UuRhl7k/2UBs3vAUtNfRVXrnFQLgY74siAfx2C0kt/eI
cr/jlTDBle9JQkVnb6+JhxgCtV4q0+Y4JXsP9h002+hVTaH/CIyTnjBoa34ImZi1
ekVA/Gsd8VWDdp5jHG6y/Xtaus0lkWZix6rdEbJ1U0f/Lk53T7gjOYgIO9zxVs7d
IR0JLf4/kozMu6fkxrGKdrpBr1bG4AIBlkJiSt1ZW187kEoA0tN4g+McevAehm84
tMEoItqMhRrnXkeEwSq+hxQ6rkP2aEwSeTiau/PysxMFC6XLwALLtFSGJWl8/6EE
nULz1kUAH9HQmF/rykBB4j44fTeFidmYggHGCpsxzpf3JtFil3UtID/KzVdrIbYQ
9YVhDBEHMdxc5fGFHqv6evA6S893XsQMe0kJqHdJy6GRJWnZWDPL7NwcqAGUM5eA
Q37MBa+tTF32trINib5mcqEsKWTeN7Q7WIlVKk9a9H+3j3ASLRHW9OqlqFf2lOlx
YLm+Kt+Md890rBYmWPhwcmXfHdEQyorrmUgEyPBok4s3vgXWUygPnEHmwneldh4A
cUmz7qT7uT6WMKFc2I0wqBBPlJrvRcV58vbVLLx6IqCslVmglqGagXbba0YEnaTA
5mk08zPKbMEOkSlEzPboV10BBIopYYYia8+Ln27kDHXxZL1Tpd7PCeeN8lbi3QIo
GzFXq6YB6dxmZgxQbMKk3GfK9QjTZL4ujts8juQODNDhvk9uOlo6qiN7VARVcMn1
0VjVbWLp+uS4C9CzHunae7d3Xyh+LlKaUjkNjUeLlgfQJHW0Qm2fjggybZkSf0DS
c95tqbRYXb3QjtR+I9JN6zrlXnzVUajo3FErweEJ+NwuJd+pxeRA+bF2Z5v4uYC2
28rTj5mwp/5lvnQ5tADeJGGF/3o45Y/irFB0cBiDO27WAePJ+k26l8Rd8Y2oWf6j
NzFFTORfzSnzyNbHworK7YDheoslWdEQEDXwh4HDFzJAm1tcAB49avME7DTxUSQL
4C+rwbEkSaN2CteH0fiaDsphnxr4pY8VXJG5kZqCUhNum45FGPYGkmQ/ufYdMq6f
4KW333CWrCvXAqNyogU2wSJwp3HP885kbKRbyjFnqrPRV7BZlVy3osL1AqzJDn6w
t5LSVHHM19tUCvvwvkSz6BGbNP/+GzZaSVd1Nc0kzyBE/oZrtpW3gdYSnSGBEKSP
MQLSSlwoc+gRTAmpruBVQoSr9Aho1N6A03S3FJ0bhgYNFhn/Lek4Y3dJkgdxFbuH
tUK+ZC8QVze903LJTbLuXYpW3SKAy2WWhAac+MT+JnC6io9/c/rU9gBy6PaEzNYN
HVQkPh5I69lzwS4zip7gBdcIO3JLmx5IYY2PHCK6jLCJ0qY9y8YKUGdFaUcT4t0R
AN9lQpBhUEUb//pqYLzzmpiwhAkABcPTxn+Kp8W52PD3bAh1yqRe/uVrxnMBxyvr
ETbcw9mgGO+/4L9XkYOB2AdRzZrEv3oN49fFm/OslEuS3zw8LMVBZluBJts6eMaN
/irlh9pfk438kvPCAuX+YjnoGu2lLN0jHjeD6bjBp/6ZCQN1aDaAY5d0yDkNgrJW
tMf/EwgWhjnlIIBGKIMJtumdIkR5XP2MMK2n5e1oYzx10rvwSIiOwLF9JOghTxyy
P0FjAQp07FQuFdVJGeRQ2aDdSVe/Hgr2A2JUPjdkUhmgM9N8BtVsqHSd3htGmry8
c6neNoi4N08wmHLkpLIGEXNaWyb1l8/NOKVKICO/iY3VSrqaTaFHZDC+z3BrRnTe
dXqwTjkX+sdWHy6lNbfpoNyHizuZoTRwQ81Ft39GVDYVyO76oMA9rMHX+18K/n+T
ukaJdyczbZQjMVCOztSURzaPZEM9Mmb1lh2+tsdNDBY1Qh3D/zUuRDb9RzLYkGG6
FjM1zauEKWMrp2Ms0S5AC4xf3If2LG8K8E9iIXdP0zc6tGC7UMKGC8jnquLsvxdC
MOT+FgzBNToquXUhkifZn0M64nuGj0yW2+MqFQgE1kOqkpcuC4o87cWhPxu2Igvk
Z43nSBtKhfCocL81o662ADBdNk2RnsaLhUEl9VGjgfhpq3FlIAhR+UZ46lF1GE8P
gZoEQbbQwyEvRV0Q4vNcORqUvZ7SnZ8uISF8bFcBwiLobO7BVM04FKphLSE3ZXD1
BaI/ex39jvZBogwu/LWcrM5g3P96jZ21VMY7A7nfh7ruJLYRfAOLv7x26btkY6MN
iBa9kFMz/kFjRboL3Aq6k/nOpgXWEYPF+4e8V+lzWR5O+thYeWobsScL9bonS1Q8
+VjNdNqAD6aWbmdIF4q8UOgeMhTjVf1y4zQSFQE/s0aF94b9Hny+86vq7RsGhZtY
ugUlPRF57q9G3/SNsgYq61jFF5kR+YSCg2xKb51WZzLseIkIR7Vam/DbP/22yTap
vA43Ruyoxe6uBqViSW/pvd5B8BvjQ+wHlnf/S+P1AFZDDvki+kYsYh/TbzZ8f/+I
vAn29KFk5LKj1wYiGcYZjIFOvBxC59ZmOioGjQUUNZb3KCfYwT9hf+wt8s465/FF
pmrsKrHH88r/H9AJS8GlsGGoKCwWeAYGEfcj3LK6oByMGDcDGpZ491JNEtfmoxhD
5G+6IKE1Yf+lW6lypxGolRBxWxOpwBtb2HDT0aAwPmragOMTIoia9cIx+VhJholW
ky+TT24osQbdFzEd3iqtq3JVuHhwpNj6Dn1klH8msIB5kPRrFiR/ou3LYn7gSl5w
mhINE1BfpplIPYcRjrI5cy9+LRZcgyxXFZUNgPkKB/ZNHG0IXhKBjo+1hyTppHnH
S2Z+GKAK4pndKlSI1POYpaeS3KMqJeLT0zjX8CgKeqZ/+YdaIh/ymgLdrREhamEm
gHbaoXKzXywQBkaBskUd1GVnJslNlx0Eity39LfzHS8pzXOMkbkKKH7uCrdGJKvN
KSkG0bxvNWjYwdzGyFgdLZApFy/GxKytQw1y7jHPIWtTg5RT0LDLfVx8t7EEublL
UJr2Z5brkYOgQ0Z9oKYHBeWHXTjsxbAwUcFpPWjK8Sl5JGVut4t2IHRjxcncqhaL
NKsCe6eEbo2Rmbz0PEGy6IA9wI3sC0NBzCU22OSsQWoXHV1r2Ay3Nd5/RkCfgwr9
tiG0q5J9eaQ5Tkt3JWYsHj2HeHQslDhZdQZ5AVOt9ZYXx13+/C5ImTGf+xK/GyHF
lV1C4zT+DyEdqfcqDjLVTrH8EWDHiUwbiBLEj8aDfdIFpUs6ia5tn6DtdztkzcK6
ktfYi4HIsVzZTSFqSH2hLpTAko4uvLjCNm57QfPXknovK3vSNwrn2R0KO0tRsiXc
ZRJVIseufCFPs+UujmEn2sDZWfkazhPomeTAivUbfUOSUIrmAXrkibenZe7Iwbt0
7z8PfotFaFgpHZfcGVEANKsHETZo6EeUSUPwsd+19KSjbDZiY6e59fqXylqN+u+t
sTpb3fSar3yC57fWgTHyw00F4jCR/bRV6EfIj4lFOEflpVBf0Q0zP845xEEYVqot
jU7yfF33FWEjtAP4+ho/04v2l6nU9A30wX43tWH2ChvC0eOhXLbx3NxlWNeMBuVv
kcEf7Knj6OIFt5oMMEzUv4YoEzyROXxxcUkksfNnn+ITY6FgBNc+V9GOSiyUYfzb
krmLH40koN23lLH4dEthLtAwsSN0kb7J2NFSLnwNO8x+/wBquaT21xWEQzEQRJnZ
a+U4fw6oJhJ+S2DfaD+lyAstAYkYNuiE4UFnV+IyOQmCiHUnnGWj1OxiOzblLY59
fsLDq3aalPXXCPF7BuXbhPCPY3a0Kq0ZF3Ruo2XS/a8zmenZoDE46pYZ9m8gTCdS
lEuYL/N1vwxfKcCIBDC9sZX8imlCHEVhuwkh8Na14ICKmm/iwnNzbBFaIs5GGX/D
RVavGVLXUC/HY9qeNlTzz1Mhpx4K58JixzSGlf9jRYdfqGahcvRpg0pt9dE0dQcF
yuO+tsdXGsQMoz8ddY8WEZNt99+wq/MeEGxY6vtewBSRrRHzg69pnIKQknmHxwWg
9PTPU8VKNDEnRT2uPZJhVkMV+peO/VPBEFXMHnonD2/rQZxwp0DZCNrlx/05qLOZ
47Ozivn02aRt3QMetVfRXoUuQ/Ao7Tze7GfzOTw5nw+evk7sE659rZMPRdkL/GRb
DmWFX7EB8f55kx9udr2UjzraesEMzQixX3FEMBoO4HJQ+jKOXasPDwAibgw5c/nB
M2MamDqXd91pN+sm5W3wF/r6ti8WE7YvhbK4ZAP36Ydq7WV0KZKgqqE54jJyvXhJ
sZb+o3dqmJi0YVsfRmss88stOAhC5uvomyfS/AEjsbq2opfXXuTkgegixTKCH1ca
aiGi1q8qkpZdTPpbKZo0IVFZywD8xRt+PZ3QipWOp/8HK7B4Ib8ke2FKOtCgpBMm
EReq/W4IWF5ZB/CFxWnFIpxJ+9Te2432rcaqVNQKp3moEYXKW0FLWbK//e3uRTY5
daaiO1zJa+VyxcfkdrX2a/5NOsd4iN/NDrub94+PCdWX5+WNTFsMktEmCYbtK54r
eAwz7zIJQKSA7BHcvxmYCoyjfpv8lgJLbtHqUsH6ux7MbVq01DML8rhgJgGsikQR
hjv89lfulp9xflJEx0QW9OlbhftzSyaMcMuI5syY3eXSrOdG8/4nNmfuDH7NlgeS
PzJyiJ4h3rKWY9zKYNuKzRDwuLSDazELNmIO1bUOIklfo/M6Ge5pn05wBYfpfDfe
cNHeH4drLu4DNFsJPQf+8kTCndqMKJSv9+c17TK8iH7HqV1cPEa+WgK3uhITTfPy
ookZtUHAaSCc47cYD6iAMxmAfg911Ua/POPhsvNZwpM5QuYuuFU7S8CIo09g1CDE
qtOa6GlsW+C9zC4XVaIw5sGk56blY1jMTpol3RE9oc8BZkwXiFln1mGP10tJmURF
UMCk1oXBd0C8i+0QtPyv+e/xTuV8OmhAq/U4fQ2NhwMk/Idt/ATurvVwH/U8Cqct
mZZPzJ0BCyL/vqEBT7k6tGBlD3D/7QL/3/0+iQ862ZY9zMMfWYp/xrgsSbhWpFys
pTf9r0pVeLRZyXYK92pAYqhRU3Oi5GaKQhGpJ2Qt7u4uqGuCBIxRwYffvArmKRxm
0QCpZEWCzic5CbG6TE+F1+9e2H8RBX1YcTKd9GZt4BeFozsr3si3E0qTonUBDD2/
q1RFP++u3JL49HT4rwgkwWx26sS66eJFdY861nlH53apOBecVbttWf/w9lyTH3aQ
QeYG/tHVB7upPdEAX27FlQxpfnGbZAgDaeL2YFG16T7AO0bnajYdgmDByz/Ahm6f
V3AgiKci00KzA7bm0WE0wClLl7NOcMLp03TwHt+o3wo0Eyyb+EMMxHgA4N/ZjcL3
AZC9peQVQS/GwuL/HlgYaZKeVk8TAiThG2/1KDm4Lf/WQpYDjTcTsWfcDs7v05jj
Zgze2Xh26xygb7jh5/2epjKYIwLQtCam//oBlJBuM9I4RKVypah+fE9u3Qrf50nU
cZRN39NQfcKHK9pbWOUGfzWyFvi9kM6GEdV0EDAypTinRhWTFoHCy6xvgcreNNtL
y+MY+PiHgVwzro2zEqPoh/HIAMFQb3tnkkTYdUUNGLx1XZMvfMLAjTJcVp1Aoaqy
FzSWobrCvJAdejveZpmTZH6NZmmhxhebuEH6pMaOB//CkeOw89hBFeyJ/ErpqG7M
whBdz65oxvkMmJaTUJDa5TOCAslP7cOGkCHOd4kfTRW9whKtiv3/S0yOGH+e1H8R
2cjTHbHpPooHm9ueuKXGhtHECQndbBaIs/qnKeIHXUtGV5XTuhpn7fXNhJiRfeGL
BzIuK4DWFDqh3DDUR+QlauZvLmZM41T1l8VkpPPEAXfFlpqyQNPV3amPFO4dtZHg
86MQ9T+7GpJu68dyLCD6hMAvA/CpiQ4w4pAdhvg42NeizMJ8P1zR4FlRK0rApJii
dH8n52qhJ1Qn63anwPYna5u5z8UPugQw6lhJ2FWbooGoM4zUsEnqtNnz56ATD8zF
p9V/LKSfVUcJowO/1XGd5rvxAGWNSoO06lMqfcAoXK8ynUK90f7g5xNuNCD/yJcv
ilQK2ObFQoZ0ShNRJrB9GDJnnlTffZtTmr8nUGdeSUwb9X2Bd6elAbXODzWKIXUD
mRuO/cVzQTOvScLIZPvV250jEYkgxw4pb44IbqaJzwPU1Rc2FcfY2lv6NS6DnmdK
ED7M/Mz3X7+jcyXKt9WIp0G9302ga7gtuvPn89BZf21VlpUcS1EYUFhb+eCIB5bc
z90t0IAGlYqk13RBxtERvad2aEpr3FX2dBaCDetk7TOHJd+XlaBmnWj9G6O8HYl+
mJlmYSo3Ni/1BcnTGVicxpC12x5KfiesToih9DTw3mQz505TrF3YGzOy1MQnbOwf
Wk4Tk1BaSBfGP1VJElvvE2VezyrLtHhjGBwW7PjR2nbHX5rUdPSYMuN/vL/FgxA7
6mh8+bIHmn9u52SbcVCw11HWcbQTdx2xah0fpjojQ1jnPTNKa/Q61ZxpOLuvPiZW
S34Y+caI7fP37OXw3zQoteceEBBPvMVRNLNfsZTovMaau01z2RWcgeoCTyf7sbz3
A6a8erdZ7OAP9NWujTwSGTfNr79dyonDn5lWt3ILljZ7L74le1p+pf3j2r6RNHzw
dDeAI7bLIGNARv1wFR/JN9Bvs5q7WV/rtHcELohnN626nt88U37zpz+mi9mDLgab
zrCaoVeNCpF1dxuJFYNT+xj13JduB3CDO00jVsYNKguM5n5RpU7joJnoDLDH4X7s
nUm/7sqj8Bic0sTZ+kGA9n2xkznRY8KCFSDNcw/VHmNZESJNb1PWCCM3n6dZE6Ij
Y9TnOnPs52GWe1JvRkmm1KwqnffSOxlessCs/rt13GVKSdhQMcwkwUEuysZSTX6a
ua/QMDJ/sC6ZeU3WxNhfJcRyRVztNjkJlPy0DUW/dS/mo5HOpYgou6FgI+b5Bl5X
1Z3palhDMTbSa2Pdx+2orB9ZA4OI5ObOOaW1TCS3Hl614v0e/KKd/F7h9dC9NnDK
aIAXZIkekYnQJBV/GTeHhF7upyz+AA7CWV+LjveCHu35X9QvdVkgGHfVWKBubROK
UPIQ6nbg6W+GHsRHe/zq81CjH77lChoniu+PWn64CNLQ/HGV+y3e9xqdrUN2KI7i
ZrYIVfyHLHXzzBk0NzECRFWL46visvusjIBI/tG4YkwErtqe+c+K2s8MlqlhFfth
AQpIOF/UmPYONH2+mZYk0OKS6MVPS2Motx4gcnMO+jEUeC6/Jym3xwjeh9lKbEcu
LRqvj7q4H1hPBjzuL9/rj/QBBX1bwmak9z3MItPjC5igvIhhVSFZwzMi0gZSnE7x
9E53M/hI93J4RNwRK57QYh/2NrR6YqFL5X6F/kDkOKiebGrwzSYB3dhbEY9y7smS
hhLcOlAp4RjVDv+6obaraSmQTVdUu1Lor4duE4RRAzVmXHOjXk0+w+6lkDUiMP9l
2TBuuWinLtu8AJzOyF55/Lx8eig2v9WHEAvsjB98fYED0zPW9fc1pSJGBWcn5EDq
CUadg+cxkU2aOg83FWsOh57KsZdg46EvMJQqLfyMOsA6mgaccXh+BBI5uksKRepf
7TECDmHNpfMvmIxYYBy45mGNBRe6XGys0HMBClMWjXQaQGF3usYs34v9ol43dCiq
FrmiQMiaXUEkhZ6ADp0Q5AHCtl8GwtMD01JcQ/mHi+lCz2FNDyFU/nsEWul1nLlm
1ZaA20IXSAvFFrQuvibxHTlo8txP/4vYwp66fhq9d59GxqtKY4+b+iVnj+LyaPaO
aeW0i5nUQ0rtghL/RvIIiWJqGgW/SmhlvgxljeazGd03xgnv3hzTg2e+mB/A9pd1
HMXL9Keh7DiV/7G/Hn3L9IUoExa2Trqt7bWUMhfli8zd82Yn3qeaEBggInEw3ERE
aTl05KZO1DmhodiMCIlbUIDppvSxoS3O/5IXD+4meVXoxuRKq8w40Eadym0oFKgB
n0JIAAn2jFQjvtMkh++XX0HQyWbS+laoEXWTZ51v0jLLdw258CeRwcZTW4CrEBtj
ZjtwralQEIEeLHi/uo6wx/ZwXodFt3Fy8sqmB/SZfwpbUoG1JZgFdIJUxQul7yvO
1I4Mr13SQbtFR+p3hAxNWa638tv14qPpnZE4LqicEaO12iQtT1w4Ej7olUPJ0bBO
MS+fM7xpFPX+Im1u29pUhb53XqTllTHfrVTubjPuBDi8MzSwhpinal9+RgniQM3X
Zxqa/v2/MegsoU3XM2o0RFmz0ZvL28Qf389OD7GqzhOEcitiI9BufV9d7npMXv6y
QRDS+USvcsSd038mJjPzI8XcRKX9VViyeEey18phQx30taC4fhjTZ9xUQeD/M48E
jeWn/7uUOuHE0AHXiK8U540HZ/LI7cWFpr2NbIzCtgCWlGhqrXinjE8ddPS6kcxF
gRqSr4BP7rmNEIumDPWo+8IOo0k2UFVbqXzewxrKcA3/zqjMkItfSKjvKYVlkal0
y9EcecjOZUVuSIv2E4wQO61t27+Kkem/1OPnkmi5PnPioLlzdB4zDqHnAvw2FP3J
dIHpL3QO7nxov/yeLN0S6jWL4vwAKbAB7zsmozCyLhjdvamvPD7EwNboUyp29dfp
aZPVBdwO8Vx6Ioag9AhamO76a+U1ynu8aWtTPV5XTuAp/CWAFNs1u93M9Yj1NRXR
fpNmIBj2nbq9i6n9Gpi70bVA1e8mgRkiI+1Uov8ImFtsvAnNjmlmrPDvwiv3/3J9
trNNIDtr7HnsLTXm+IvRgleHjrk5LP8Kbi7ICGY6JF4tYfQDYMb1YbaA3JTkOZ3D
s4iFtK9NLWL8SzdhYJt2ZDiT7w84rSL0a+x3uPoSFktOoPzA00nNWANlCF9+6CY+
oqPDC0uPd/J1LUbvzTmVQ+dp8ySQ9YljyxSdOW353TPpKqBBIrY5y4oVjxJje+Yy
nmgZR4zYfdT+HoT3fVJ7IKIUqxdttWU63nFW7zkzloY+qMB2QEN7um+WreER69h+
M1eVnF3oojGyTMOCUqIKAEgK1sYp1V0G/VYuY6VdT7MpWMXMzmhk7lHEN9WpiANa
FDB0vLzymIdDGMgzSBsnQ6mpe7oaJdCPkXC+T75NkagRfa4Y7LPVJ2UA+z1PBoDM
V2zcrpYLmf3HvyDJXarWGQpR1ETc5qFMEKl7UkvhMUFxpZ5T/Slu+slOI4afg2sr
UHvwlLs25+NQaucWmHzmkjG96TSa2N913lkYoItdJJzyfSr+LzeAEJnfsXo7GSkv
luN/dxYh1CLbC8Z3vhyNFFolgZlf8Zr2mADF+3blSYosHg5/r0l7KFex5rYYH+Uu
7Y5rNNQt5YtiQY4u6pcbNdgItlG/jDh7TuzVg3kQCTnDGw/EiRAe3GuZCZ+HwWRE
n1XUGZ2KSo4zGecBi1FgKfd+NaJBoq/OhfT+X8PMJ27BKt0ztwr8UEKpZx9Do1t2
WJ+6aWB8EFBNIL37fgA/z22gFchoI55DjTYwQOEKRXBNnnLLP4HLtJSQVD26LNdw
VzqMdgbkmvUplh1NnDY23yZQlrlzT7kIKG2aA7lwbjx6catVoX4qFwYsFzTREyCZ
gtLN0sTGOq2xRCRg1PEShrLQUeKhW2UTAW4l5ERxlhYuq/xldktVuCnDq61vgWaX
84Y2D+3yGFn0ockSA0Kgcj/+qEUqLBxC8K+AdJ6vMWbXHXFKUXG5LDzuJomr5x9Z
cmDiTTCdql+kuWWRJbEQ5ETAuY9EK8NqHIxByH5u2TUlMyUQmMPiCR40Wz48sYm8
7SyZhgH8Ez4fKS78NURYuo+bE4D0/Pn9/TaZCsi+MLD238yqhK2SUFzcV+1gqsfw
/XjZVTi3zahIyhoezAc+etl2k9R+Vh+D2X8ks0UrCmlnq4TW7R9ZMDa2cmhraMLF
SMlzm5wahCH3nwLdswpxS+actxJ1M5GxnPLQV7k5ydu3raKXN7QWcJfBlz/6aFh8
9eGcqZS7FkS4mV73yeL9wMe4p/iRURooH0aEHb58qq7viquWWSty/Egqmc5kNonF
QBA3o+74oi/BQJvFggTDhCshZABJik6cfqNyMaT0lSIlmLIqY07dAC1KLP7cIzBf
e+RkyBR0d6J8bVMiwhIB4+xJzl2kVPafqA92Tmgbalac7xPexMcuPmgaNNCmJ/Br
n4DWAwyybUXmz1AkbG7ukBEkWCOI84F606b9N9AiGiVG2eXqs65ssrX22IOZsjX7
fnBL+p2zjs9Vff5FiU9u3g4ihhjkRbbiE02IPNkNcrsceYjefa+YpJfez/B9xmar
lhiXN+HIgu6F5EqrQXuc8jxtKBYJZGGoa86mp0CbpkDjiYHTnHIiQoBHd6Smw75v
P1koUaLlrdsq5cri+44aasbRE1fyVkAu0ebexGWNmfejGTLzjNZLCJ50Bbs7v9n3
LFvUEhyiYe8mk0vCFl7CfnHS7+1PpsctC/bPlFIIyqCmvr5oAcyWIiOthAAkjboH
rkmN0W9V/FS2JYa11E4gZIG3rYVJW2Z5CmphSsy/HI0D9grGQkOyThgckikfzFXl
ZKpf5rzQiw4y+rm+jHLQEwsI6vdNlEQ7jpDf63Lr2s7CWy0/xZO0cN+NjzLicGxP
7r20qmar2ZNEm+0anCypFGGwSbcn2wDk3+uUZ+4oTPa7tgaGtwsIpnOf+uqqjgJG
k1sDM+/RrYZ4AT81/6qsf3TtgX5HObLUjTtV/EhfGB2wCRqjff4Bn0/W+78A5xJY
YLz7eU8S69FjvEmZnBgJjasFhBGUmZR415kLBdy3+OatUZnj3rYBBMgCC6/qDBU2
52VvJU54AEO2jFwj+Kj006MDffcTaK3yIpXHUvfwm5g8aCH21WidqDW81FKBNcN0
osZ0SNtLaGNWBq0zcnxZZYa4sWte1nmkoyo/pF7Sp4kQxbHwQNH9I6Eiwx1Z3+5T
V0IuDwyGk75p6aPIRNrly9Jh69b7jqs2cFZ+ety6t140ZwvAqIj2DAyqcryioMOd
7i32B5AymJfRE7n+FZi6ABuAc15NgF6VVFregyPBAOQk5kXLDU8dyExIHWdah5mm
9CbRgzjKGDJfX62RnEgvk95EeJRHQVNHDtX1Amlwlmevh7/gYPjgdmohGG3a/tPo
1F8pUtj9a8ZlIPNU3iFEXObZVfqhTwCtVW61wiNKVbTVcsLNHOV2iaYh8ZLPX5f4
z3LZ7XKEhe9oE0LLAS+3XBbDGgZoU9v2/EgExuVKoxTn/z0Wlja2nxJAGkU+BpCF
ohCpF5ukUnsnXfnwH/wECFTmd5tHx29gCvyaGSlp48ReGOVBMeqWpjHMEvqfgp0A
XKAFFq9eA6VgLaGfd450r3JmcpUjyFxgug1DsoGDDwTZnAFpUYDxC5QvflE1AqbH
VTCql+kAjkZR+Qmbz3YZdv7r+TftITUTXzRDsbiuny7mSNcIBUvF1EbOSGjz93XP
zKxmFaTbhBLk9OofB/0D0ZKuKLjC4Ylx16si/zBarp6VUui52fkD/4JiDCEkVbal
YUpJ+Athwmh9ANCMGh0Su9TuChE9ZJno/NezuoDT8luSOk8mlHObgPmGLx/h5D4z
rbCjbXw6oUHRtmfc8+Rov5TYJcw0Corglhqjc1TnjG8bqtzbIUtldWjgOhxNeXVh
FsEOacCuymLLB2SVpamx+3Znfau1UjznlBwVRtwhVdfUroFs2+AHZhtA8kRXdQhr
ioqfhxalIB+0gQwE5Ewo5pyzDyLCuigqSxTt3pAUJtQX9gH3C0sNONJcGkJyrSuo
YobRpp/JwxBS2J36o8qniCll2CWwL/gI4Ie0YbafC8ikM9Hs9jXfgW171TeNAW+U
cyykhcj4l6qZRKu4FgIBsx63Fg6QqnDxu8W/khu+0gk91b8sOv/oK3yJ8uWcbGjR
iLn7ahMaSf38tidJu4Lkr/pFwgcnQ+DplwbuY8tV5paUKjTRvsFkuskhk4JYbCQ/
CHrtfTm7DTsKx2j7VOemEH0SeDiNdoxUjcDApMxD/TRVn3eJgYa9OFqVO4AY9n1T
yqkW1PPFSBIXBtauYqSTSTK8GFyKbkH73s3ZduYzZ4bTI5TaE9rMC7raMspY97Lu
btacJiv4IU1e/XHmhgflVYlMk5zFq3MeZmhsMNZaL6fVHh6IIvKBBar/HP8lvJDM
IeE9wohAZxccAPZwi326cqEYChGvZN2B/8D+GooZlT2fbJvtVvsUfaFGByHF56/K
jISn4eBqmuI2iOp1HEf9cODWw//ndrhW0E3SM5arv2jRQGPiU/thRPgJbsDEfMH0
YguyN05UTPhLKal0cJv16dS7s4ANixtArF+l+LS8F3aQnHP/vLeCM7XlCCJ3A6G/
emqjwmIZEbRQ/0jqPydeOh8OVG8zdULf4ruEqciJGCYS0diHZs2yMU8Vm4hl/0oW
qg0eTNawk2vCiUeNXw4EbsIooBL3UFZAuQHppUcMw1ftvrNmyUoEYDpstu3zBIxK
Jsq9CnlBKtzy7+yM/0dcW0M1qQVE6h34zfMHnqqTHAc8IM+cXyCq9pv93hU2k6LZ
kcjx9ucim35kMkZ/gSbgrgiaFNNbqJ2W74BEmNWxYSOWPEe/1A8MMfIRX/BVtTxO
826opD6lHRjqJNazkBJgYVY9yau9BdNvPXl0nfS1ZnvMyb4101s3iEoK6QfGF/LM
xV0I+qEeW8PBCmpS1tTcYnllG1oyk5UxWefmKZgo6vg1cBip06Pe+VHLUwEsqBUr
vq8RzI1S/GAAS/hpaZ1glcsD2ckq1NGrkxGnXgRMmt4j0O0lcgdfJDULaeDb645V
yodpAsJ5Jp0NbK1+lTeaCDZ0+EzJFgJDQvYVC9Q2bK+A0KKeeksSyat+QfHgSk5t
arHkfAtMianlu05tP1Spun07LSXFd4WHa0evVEYA2ZjqtEh7aa7nnMsVm0lSOE6E
Y/1+0/cbud4gz8b4mLUdVOcc5tmsdfcIvimnm9o8oOxaargOHMXcz+lWnio8ZCxr
HO3QumZpkuSkj0tbaTbK6GuRdATfACnl3rokT36ApwoU8kORfHpAeYwehonyo+Vv
+o6Fv5QA1RJ7qXg9vFK7vtNAb991i1pNsRBai/cFVuNGJfS0h694Dvx5XhuZaTWX
SLeowpWLVwIEyUEY4UJgi9WXo9MdF0+M/6OaDPOKTdnND2Vd/nPNwbNryunmpc5+
wUevJdpk+aYpYSHOzPSoXfdLUpqi/5Ly7kx8vFLsMW2wAwOKavVatw3MF02JC+I6
vo0VQoqb6MLh3pZidfmiDY+uN4VawaRVaoaxBOkFXWOxCLvigh9CfT6mJJ9vdBdr
XiHtQh3AYJoDQy+a/ytM7awWSv7QtLUKvztQ1G6X3IChgn6zZTOm7x8owyw2ONi4
vZcYgzXou/ol7xTAWiIeMIvPf7+rKo5TLwZwdDZ6oEBn5aDpGKk8L6IO0QxjZcuj
o74JqY15Ip9fvHwdS7dP3MxVNv3VKf7ncpUT6nPNoeeL5NDRQSwNtAGIzzD8OkkD
dplkAdNWoMeALDWXVSkyzSVhp5e/bNXG5DU0YRmkWyz3fbx6HM6IhBbyE4+4aDl+
aFbrbdQYzyMf7q5dW/EUdcjUHMDMGKTLFHYubPL4XwocceJAZrBC7CJdzCvwLope
GB4oUGUjkBcLdX3utbrUJUDbLwRRe7j3R7C0ww106N3qFIFzjRZccwMaom7tfm+b
9yro+AxpUiMIDDXpn9+f9KSU08FmbsqchDx4sagRH14ZasTvZpQoqKuLZAqpEVzs
NiH4C/bcpu8T3P3kpL9mwMQDOyekJ4dGYf5coFkoQaIp7pYyq/+VggxzU9ZZL0VR
o9A5s5e8V61DFKBHYa494cdlHwumtSViVxuy+h1ApsC2PmHOEzVezjlgjg6djEpB
K/U+c+9Ur+HbHitBPpUgWmHk3XL1NUNwk0/+6lR3QZx7z63R5/E7bc4+AlrqPosZ
cgPzTZRpiLGPQARBgYW9yYCMtIrKwfQ4LYBZ9BcwA9bUMC3nR8Av9LAofnMb2UsB
Pgq7rgt7Cms5HdPS9HG1PR9khno7ys4W4ba2qdBM22raI5p+5EvFho4MRR5L+Mv8
p5ABuGxgru+tWJ6er6yw40wYl5waZyi34tLewS4+qzhEppEqw8NKE9jT9SkO6kp7
Ijsul1Lxbn2ZOiJz7HqZVMyXbyP2GLgmsXgyLOkLzT52VcCUqKpb1LAugJJfPjVg
WUfaYt/pClpGZdKRIWlAGn4UbjsIxVM8vNXOEtPY14wICRzUZ4j3LHwhnlmnjAVI
M1/5sQ7lgtF9bsRiXjnaGSOs6+A7cYLvUeJCwUpOahkWYxZr3rnpn3ojxPiBshfv
1xlwb+UJl9AJhMHvg4hQ8noE7gnnjP90FolusqnONLaKxu0xYYx6SAO3sNho9VQA
rJukLW0EDjQozkM9ihgJRpthe41EIyVlaEhLQo8hQQbPA+3GJ/TYC8hEEd0GdQFd
EzBTdHOpmkkDByVGcBvLhGmyfSfDMTgTpqZ81N/9ZUUkyUIA7a6vdSfhqZT7+wiA
VJVKv26HY2XJhu30wqOqMxlc8TQzAd0A7CY4q1ABdEjmqERDXnRWlDUH//Jt3wo2
yoXZ/E6GT/du11Wc2o1qfaYv3yOUgWf9WUy3th4Ja9pnwG7OlsmlacN4eOk8bw8o
eomb8yzGYcDUtMEpvSU073GhVlN8jnTMocCVU9r++/HL2/q1jMsttolkIU+M3CLH
cfusSbTP1ofsdlRgZTuZ9Ja0euOEy5FOx3vxlarDmqRZlRi9hclanATf7DegZKMT
Vw/0xf+PwxhrdI5iHaed28Vnjo3YndmDarajvrmVaFbQLWql3BfyFgQJ7z+UVdds
iFzJbgNiI1FbgHRViC82jUwYL0GIOqeQSAVgYu9c7Nlo5WlWoxET/M2gEklTzV50
twNA7PQ+N8XYb6hW3IZlyI3vhjFe7s8Q576dr6D+DrU/BIYH4unYOvimOy0GI5Mj
C8XqWWEUnNkizb5eJBsWydokC279OzfP1yib2t5DNdJZfFSc5pIzD9vP6AsgQdJL
ji/rAUHy6r2Z/yRNxHayNKPI+VptSX3uRvPWtyK6vp6RPud0iZQNlvK7jFWHlWFj
GOEX3QJxlKS0y4f0Y/z/tx0DRNyuPiPJDpLC3e4+B8YZowH4K+bxZcFx//kj7MnF
3Kv7npwpZlWaS0lOBrM4lySvEcQNkWO5uMBn+/9pRSolllpjyZ0GgqA2YckiZ7F6
1BS5ZtGJBhVfQNan49BWDgKmtn8ZYaseQk0tlNrPXN+otNqKq39lX144PTAOLiR2
fsCQ60Qs64mlMjEeEYdAmJ9xe3lzPkGw2KrftlzwHu4orzx2RKY6CWxsAvQTytlU
0waYRGxHbN88s/dgQfW3PekIGxDqeHD1d/Gh3lbd/PmpV2prZN0zIFckISBnPHLj
Gp/BtyQESeyE/qqdbzIgMGxqMHahxEerTQkp9zILW9PiT4VtDqxnMD88oZlcuIks
aO3+1oowZqd/AIoQFOmCvcwkKMkULVOUkuACA4HwT1mY4smcZjM/4lAdh5jgRbXq
KZLyMcdK6sKm4PZPkp1p/4/cFt2xVbweB1aJWT6Rj7Ia+aGG+K9FnC/UXlPtwaTC
9RuAI8xYJkpg5FzkYvjoghU37s2QAbfqw0EexwzFChIzuORtfWHWPLM9KF3QWh9l
J84ax/fkNQJw0crDCV6apChvdtXjT6whpHuvWPZTq3ySBSMaPHBHd7dOnAzkJGoP
EVY1MNiBwcJSHRdOwzLNZnrcRkUjk/HEnjE98/cbu2p0aLqynDpAWsIfjk710sK8
UMJzGZUDheC3OXs6tl00YlFua7pMhX/bOop2eMofBfVZFl15oqRtELvj4w1GUlTs
hy8xhcT+jLo07ZacXTIXjj9BIdHsRACcyxbuUZKiLhUWIhoV59ps2J89owPJU3DD
00EQt7CZvJD8ndZjnPQ6hHekaas61bU2eOZUl0x+8CDsrA0qCr/027oEWwitmDtM
m3L0IP953/RhaOv0Jnip+pFZFxac7mGt8lMstcHmO/Kl13bJZkLm+U6hcMnt6sM5
sqmjtokqsPcbRrSYHvXCIR8dFsc0c+T52Rsk8jP/F6fPYtHe7eLVyxCJmAS0sa86
d5BUsGbMHTuDmLAni3XKISpkL9obqHUndlYEIqwQXYNTHKPHf50Y6rHfN4+cAwcC
E9nicYD9rtJe2NwTLEhBLgFhCC1fRuraSzzriIPogZQZOU+js3pS3Yjt84E8NGew
Hi0MTRNt0OunHwLTtz0aiujI31yEer0xDLmaD7E0xA0WZHnvUttiBBz7TqxAGxMq
MUvHynsCzJrZLXZuXlESbIRpkNIlAyRxOY/UR/FZbzQE/B3yMQiDGHSmaSzeRhIf
KeKqmheaCRUb92qtrGDHQ9/FjB6LGbYFzpwEskSemr9XEOcQYqs/9Xxq5LYLJgpz
2Mzvg2RVzKcXaLc9OO3LM7jottFPCvopHdc+qZwFU33P9zuJql4ZhiDPu2m8qvx8
3qaWjUABzSCAT4uF82nvIcG0P2zjfgs5FTLBuRlZqubK5ifxdHCUI8yUvM3bjcv1
NIG2rN2jAKKW5BindDT2g/cX8pgaUYG6zq/nLZBKJmzIrMRjIVlha6LdB5ucGFtw
k2nP+6t3FXX1rqFRUjpFt0EY6EsRzEi008FgWUyJbhq6cmm4f0/0jddMyMqEfDi2
ZxhaWXUx/QvHMr2NKd9KkzNi63fJWsdVBuroH3v2ni4hneHv7xNGLa5KDsRGdtxZ
nngUGn9eDinQrvbhylgc6dGtD/I91TCqBovIN+pv0L4Oxa6ExQOVKiJTL2xlUTU0
oSk140ic0FCacafXKGHt/RKTaFqIKAceQptLAHj4ZAKmYT/r5a6LCddep2/WDj5k
HPB+ziZXSgXlEBoNgvFTYoTwwexZJKRDLmy+5bvjSU41Ty6x36qTDavpWF2lvY0/
c9ki3q8bf/14i0QdJKTiKExL7Cbx83GVa0WpTG5heO2zNH4hOwhvWOvyp+6lEBek
dwClhlylkVrd7FdheTj3BOuXUxe8h4Mw1+nZjLu7r2s/8cLwdwesHdtSME5ATU8y
zg+aFxQYg/UZEoXEjOmPOmaFHtjWoySZxQZX+uCD6l2IuJPyEXtfoY12TsXJ27lV
cU1mVuQwwVDwxwl6Y2ZCwZoQxUoQMoBfQt95bF3bB9ZtyG5weWrXLJV2HT+4UBjE
7RglaLbVz0/A2LoWvhE7RstpM3XJ2MIc6EcFaQ278nYPRvi81Q5GS0UHdMkhumEq
Ny/n/wSycmcSvxFgiUCDLuLJpgxzFdvDXnE1Xr2hZUfzSUKoDMfqN3EiL7VVMZ05
B5TNyCeIdhw5a7FQ3wg1+xtgs4Hhqa5/lPZxH2INvBu7e37+5SwqPUiquOu0uRuK
a8dlYm1+jMP/+jvfYo3gTvoLNEBls8MzaXxiAuGnh9JKVjp7K1sL+Xy/nQEQB94F
A8uKh6GSAejqWpQ90ECSPnKeRz4lilO5yvQ3cYcvk7wfH6eL1ydNEw8jgKpTDOhQ
3jM5kpSNORfLrFckThcHoAGGEVrYrgxL2Kzv6XYQNIGTVrZgsMK3yBrBR48oVV19
nT8HeQh0dBQc+zIjCSMBJhkuVSjLzTXt1C/klVmsWkXTBVDqqCLFCTetZIfg8mHu
m1xIVQdZdfFRIFikFengfUQt4m3d1ftg0sXtbo0I6ijWfH+Q0PvkZu5oj2yZgW3u
3/WbXhyP6cFpOb5ETSYO9T6nRpgMugDRNGhMtnhHr5XQAMHvHGjauNdhq0qpSypz
r6gjpXp7eYiX9wSQ1FaIKM69L0JRlS14d99XByJolcOE7w91jncEK0jIE/9mabaG
heZAaUk2L6S84lf7ONboaVqfRqOKjyHrA2xxL+oH5mCqjRNc886XtHmVO44TGKOA
qsldkibZXp2M1BQ8vL54b31lARmvMQZxOgcWZknLY2eC6knuuTFRQ4R4QWxAUIhu
UIS/1C5lsq9t4lMBXQ+qXEEdcE84alEUMVtcVif8vEWSIL8w1EUOdRWrSxuN2tst
uIrzl2W3PZsxcuauoNfp7aGbWOWoYuaCVdLah+RzzA0UerctZZBArGRUNrkZAVZn
mVU08eBy4+LLhMooUCd/gYLGYtnFqSsujDrITc+jAhOs1bQ1qlcd+mhWboHl1IGe
0w43k1IOcLvfyV+CpcNq96EGDcrROJ6yKVjbJtuHZGeskrsODP24gubw7ERx/PkM
QhL7rIZWHwZ2iu+5Ads6ZKZFKa2gr5vfp74bgK86M04/td52BqRZGQXFiAKI4nu4
vWWTUeeWKDiNjDseDCDxAYQAdzgnN/QQf3S45ao8NrRI54bgRCeTQ6lhBjSeqGRQ
06UoTcidd/mB3cEK+gt51vSk1sYjGu8B/K4cHd3zMEhsEJVuFYseIvpzbbB4tmN9
afq8OXXagaj4dm39KNC/5Ru/vfk3X5JIcJ0EHFlOsEsP2Dlg3i4TESXP6N4N5k0L
cwD5aoiaSDvb9x08qczW/DZwBjyYpoj/nGoLfqY58zNgr7yXigq4s+fF07xpqEfO
K1b7Jk8F8n6U1tIhlMhS700tRy9JXO2YWIuhgLJp6TRkuptMn73uj0yw1bdc4zt5
Qmituz2IQhjQj2EgIk9l+I9ceK1Jq9a+RGYDgb9sSMe+CPiD++vUjKFEugbN2EpX
WxBpjvSHHYrAvsijuqd0b0rNBuPt5BD6tOesLKoDQy2hHI6QcbXISPk3k9wf9a7g
s7p+dGRXlltFrAfN08XC1b1VZc5ZGcowrpHoWnpqV9EG165h67OyCdj485y20F57
A7WFUuBJIC9M9yJRNZPOjhw96DPOSjkK7gPN2ePTgPyqsXuEt8rNjjE1oL+pc7Td
StEHdK4yBpRZJgskylYsmFp4zB6d/mAX8vnZ54M9eWRr+43/FNQrnafBs99nidN5
0SLcrPLg/b0JWPto8Mm26zRH4xoJ3lpEdT+Nu+HmkLFzfKhpqORdzgZg9hvVJ0yH
PwcjYMNzJPaxoE6HpRnImcZ0/51c5bqdJT4rj9RA14dEiXv6XFdjY3l3pb2THgWL
hWKzMpZ0Tj6ZOnj3N0CobplXYx+KCk72t2tlOyT1giG2ucbPkZgmZAargHwqZlI6
4Gqs36kJYohQD95FdAISY51PyzdtdZXFDsPGtX8yXqM8ZN2U0LV1M+rjPtMjD90t
+5KOWSi0yEKqsjKZs3HYT7Xj60VCZ20wsjOWyotiDpAI66y+Lf9sFXcWFDYkt04Q
3BT9c/E9x52ecuCuM0ApHhVh796aAoRCwv8MRxRSAuDv88mRneHsAXsjoXv3yKJJ
7DhmxjNj/imttroQ2rnYA18m1A1cz/9QXB8iQ3zAfdVKxSsNGQJ5FFU6GXVQ0lfd
NIxNRFcNZK+yK/i1DMtFKuOdbLM2w5qnV5C6jAExs5glAwtAb6XgslMtGCWX0l8q
MjIIQah+sEAIrkVlDuPxPU/wpNcN1p2P6ZF4rZ9RKS0q3WpBg+rv9hZrec2gt8uD
BPGokOhn/67fr79Bgrm8vuyZEhhPh59/oaPWrD6q8pPyecfNdchPFm4vb7KKbFAC
oS0ZWT5OLhAZPXZCIo9kBnJqjdMZUvLrEVQqe+xS/LAwJaipacubpfWS1Ex0tzu3
BDCuOhyDDF1oAvyIeagwDEF+yp/+lFJUcGMroMiX1VejnwIgHFCw5hE2Hh6nLMim
3JL0dNY86HZzH+n1f5wITAjHzvTlb3vCLOwApxqQW0EpnjVFaVAzz1VTRO3K671q
5t1YGgnIC1X+4NpTa9QZ6NrAZpfh6EE+ti61SNx6kL/r5xdJL6xQsuPhm+led5Sl
DyKX03+bCiI5vN4JmDNXmszGuCz/3/BuWHko+ixEq22AI0DmxKpsWW30kFPWYKHL
r3O+JUNfZv3cT0E2rND1mpdCePkjZWxRXd+XrT44OmPTZZs0qXUfsZspoH29C2p3
BoToksXsYWzHCH3lA+2Iij5vQIRBNkLsbR67xKxBVOl5y2jkb/MnFavX5vAwF6jN
Cr48HO9pg1k8xDPczA0qQPiOAZzgo5zwtY6/A8if1p1Vpe7R0qtLAAMsGvO7MImk
AC5KZElDbSHG3gOt7pJc2d7jj/Rm8OHcs5PEO7rNOr44ptZRBPafGrn2kP8Ns+VC
6BPkshuot8qIvOHUcEktjuUMfjxGSQ19PNCzRXqeIAEwH/LIo2Nfoq9uljkBRDgo
aWZ/hxTGSw9JIdNABRc0VNw00PqZP8tj+mfu4BdxtYMyA2W1U+JvFaZXZdxfvrJ9
Bx/Fz99pNzvLKn9UM/hSih2psndJq6kzZkkJpCoc32W2IQ8M4WDg795MEj2ejUv1
hVtJXHdJUjKfQzbud0zDg3jH4S/4E7/Y54JNWQsdZh3tTtmIujO0kheHw41C6J1D
jOgO1yQope1d2m1TAa//ITIRcuFxLmaW8c5eyRel9Fl+YPp8e1/fjpipUGbguD5l
kAoMo9efnAsSqT8AQFSNaoW/gJw7Thad30qRa9TXkJfRZnq+wpm9uFY1Bwy5GwDO
mCLHn6+GqDS5EyPzOgQDjsy29dwf4RzE3nnoNt5ggUbPjRSSexg99MRPD3cBWGFt
MZnGpCSmsmzNhBXue9YW1vmzyxm7sQmr1edh4q+RTa57j5fCIL/F6Tfq/LWkLypy
iw0D3aqaibVq8pyRCmGXBljZTghRCJlIE9WsUHrfYVkwt2Gx/tEJ6OGibS+hW5xd
6uECvNkJqllvSUCfcQP8a0QS2tBDgTfdV4k/h3JUm3KNSaYVV/WDoLM37nGCkegf
dw1Oe52nBULImSlHhHR5K2iNwzLvJfoqZGuvb7evntBoeGU4BNzWJcaOs+xWHsop
LPl7FaFuInB8yIAgUD2vkRIYDeCw+/aDxvl3qkJnlzaa1p2JRf2cw6loGu+V4RpD
GBurT6C4GwjUdlgOYo/cC//naoexJjSqqOym5vdQUtsffhCOK4Is10HhGE68F/XM
9uLN0Ekm/3xoacEsDQMuY3nX+ie1dz/rZnTbzIypTTRBYGw7sEz4Ayegqf/znMHQ
33lx8wZKBfn1nAV69jroncWUh/XxQwpp1MhZZoRULVQD3HQnyqB0B/3INbv/tTR/
zKSDoX4jK4ihhFO2sSSnyzhKoUNIAkn30yGnTdP2Sq3FinD5HeZEDzFrnjUC2au0
MUrWA8qG22C5IHmcTaImrOjHRjdeuN0paQWd7tdJ9VZ05LJx1O8hNXaj1VpNdXt6
outmd8iRtO7yXwJ1WhGTJjOwyx0dQkDLuLQuazIn69g1ePv1Bf1mbKSVRoh0BY5v
WSioKlcDQGqmR96NerRicm1lpaMviOyerM7SnWqU9jRr4+2DEN5dEOha5et0n06b
6SrSUDwbVYKhCT0DwIlgfPwhVZwE90aIYFf8zunB6Qou68PBD0TL7HCGeQvpEzea
INUhCcEUtvru8rIfZqGKNCxCHuvf1GByquJbTTlD5uWXgdt7HbuEuAtVrCS55Tsn
tDwrPtaFR97Ut4HNyx8xEmtQ92Akf0Xnpj4iMpSzdpa3zinLzT0Zijb2Vq+wrkyf
/r9+QkGGcqdnghK52PUnxMIwKiiQjjf7nu1y4fZMgaaAMkeQtM6p7MLj2IVDkL9B
6yzBbLL0YsIaZ1x010KW9pY1geAILeY+M1iSPti4XRa0b6NjbtQxvzn2+MFhTdAN
xqFCPHf8uChZch70pJpyehCzVeYYip/LV2J9UQ2olkrC5MEyJfBPZWqGy68UiYdS
06l4oeka+4CP4jJzb5ngQcwxHmgvrGYf1on4zfHdYXHSXiRfiKGJK/hNifa2XSkq
avFhs23UYslm7ok0nQP/CaDoRfiNWapyPaEd87Dt/oT0WlJdQTrW1TIBdM4NR0Wk
nCJCeJ9l0CLHjpSIRTqP4Yq525URQPvDLH8YuH7+eAtKsZdrAWTVNKSaxwcbR8+9
kWVjXGJdz9xgx/NXqgyK534V1kL9iHz5P6jpav299ADsCOzB2vzgqFbIS5eSaWNw
dPJDeOHUpGPzbfWysWyjy4jzkVL5h5ia3ZSMoQajHQsH7/WDjLGOyWhL7xR3r+Oj
UvBiJBlcsVdsv/FCntUG7hCR2svvQ2RVWl3dG2vjlH576If0m2gNSaDrcqi8kDRU
ubujbnc+E8MJQk29ZN18UfX25TlrTdCaG5lF+MRoKzLt71+KEpuraU2pfc7OzDZl
pbp9iFopeA5UtdO5E8qxwOG+xTPjSArhnzj0VzmY5qYrrfKCEChBgM2LNbg9eyXp
Fw5hZSMBR/nF70gxr0AuEwvPyj80M5WwFKE9yJ/SaGLTsFVlt5NIBEZR9KdNtuT6
F3erZuqBkWgZqNr/65u7cOqWutbgLgLei+PxSypPcCn6PKYr2/uhJcAWKFLKfjNg
UC2f3Kl54bzIE6Xl9EbTu+FKj92zqGaCVNqMJbfkNUJtvMWOeWyAxlPR+UQq6o7o
UZJV4twEGM+jbEmBKDXHXvViI6BBTBDFZicvpfiGnd9BLhbkHgAu8f3DwtRSuE0G
/wdQ+IZJ5piFyuaBAAYEYRDIriXVRB1j4PhndOE1kwKRlDTOfZZWcLxKXUzGZ0WO
wncIR2Bfr/TV1NPkRBezvET98AE9JIEGLCzUHOEUeSjanhJkBqJxZ36b72udQW/U
Xt8+/4bTZlpaGKdmZ1CW4NYxHJjDno/3t1gFeofkmhI2ZxMSyLKzVE6wknyMnuzG
YDG/1TM7aoh0HECsXD7wT4JRd2lbN1m7Y1ppHUI93lhJIXlJtTJZvarDUsEEfFPA
ZbaNpAFJ2aVGcGgSIg7C9MJiFG4s+VfwDRNHxt/EM6CJKF7RZxOeCv+w9OEbcIk2
llwc4W39OK2nkiKrN6qpyURBlHSmRwBY9KhW1wRXh9Zag270TTBHmph+Yg6ZSKLx
aTj+KId4hjUZqWoX8LWAxpkZwtDaLPUZmWxUD3h2Cp3HBY8dINfNdFkQVApSOXW1
0gXtqamcJlAoizXR+gAjqSDXB358BMryw7c+LYBl+hxRThqWjjKOQ2hJa9mDIgZh
V4AHslXs6N2pvrNuDlYYxQVQ4JldRFlgCYlATppYKRxsynOhiPoCvgrkM1BlzXo9
2EoFs3IUmw/Dn1aOZp8hE8kJ0J5KyY7H2jcqhBASd0dksexOkEUIYyBpMWVr/LK3
pl1UDz2zbxUSgFhDn2pJGKzGP5dtKF+U3/Mpwv/VUmC9V3TsqwJPv7VsnpAPB1ne
/MIGh3Pvz/al0RiFx1vhjWV1VhO/9K/c8kUOy1EmDG2y1apDmT6++mCKdirvpHQ4
pWAeEj/nwIznWVtLPiJ8+41F7Lh7eOM0+Lt9PFrpvWdv+1PPlrsssf6J1+cap/CZ
jidKa0jAyMH+0w6PNvOLciZmQlo3rbv373YeJGF3lz/o6USFaqqJN6UHmGZtv8Ky
O/PYLn3QyYPz7mCRqheP97Z62GKfXzrVO023xGhaj9g8fms6Okq/BPjNQJiYyVd5
LsRNEjL/ToLYjQ5+dv58Qut/bJKI0zpnLfGhEp7+z8QUChmnufxa1tDN1nZ52/TQ
9BiO/TVDE4OKMEELXaHERnPrZIih7GCM76jPjbu/R8LtOZItMQ2It5vkVNXnsjBQ
YMfEadLwy2Uj3G4JA6o0BS4Az8K9OSYsa6kmlvdvcLl1pcfVMip4tvXhaahXCi+l
CWd/VrFG0r58JsQP1uGmvy+Xk/iQkQpuPvSLqZRzasUTGuclAm/sSFnUvTmbDZij
14/8Pl8j3NpCVuJzYkSyEINIxM5pLdGymIVqt0wDu3yoU1422mzytc0CIefv8z6S
LSGvwtg1rq/YUhioUY1bTs7gMSFo0EzZfOokjC078CR0Z1KqjVvZhuzwvxpJCz2e
EaF2LWVbTiRgXpQMkVaX/zI2NZySaPBLLz+5ybsJRCan05qINPkqjc571gZO1G/R
CtuLzQ2EmRlcR8emnKSbc9AZDbHSq9XTFooqqqPFOZk3nFc0vN4sBOZTBNiPf8lZ
OtUivoIjXNVg9zsvcQvHalwI3b6Q1QdACL1AYnxV/AHKI09UR0oXMNuP2Vzo896E
wjPgnLWdGLEytvbUMvroj1/IyQhbWGVcQBDqHML26WqJNDiWtQF7zGPAwGK5wQkp
u+qB5XOJf1fCDXQ4hz5+FXBPLC3SDU16MyQlfa+CTa5NGUxVhwngexOYoURaDcbP
Z3aq8Rxq5xJ6/8Gopi9+5cOX/g6/ddIxMceeZyeVu4bC9x9B/KcTMg15nFHFKbVs
uqWShzXQWSvvL3+3ibDezo+qfsau08YUx5qIbxhXH4hNZQqcYrNVdAJ8dJZ2Dq8F
IOWbRO8nIsHHMLpWe+zfR+9ZUYUru9G+kO6PDc2NkF9bWiUrfgBNVuniouwzEiPT
KGyA3pMOlBOttRGutnLjSLFjc6jjcw01sF5oL0vZgpNVWTqiWKbQ1ODrag07+1/y
E1+qmQqoSMja48gSeSnzXeb/Dcv0Qlct93KW2e4yHv8DJmPIurPuJtv8GVAgH7MY
swDNiBo1C96En4U90znxQSjm/z5ljdopuyJwnlvUwfPIXuYohYbQxCLpLH28QOKM
U8DByOmvd0BG+BqeR4Ul6GDiZHCzIaDSICBR2Wfqj1NQYRqk/dFsNhOEDDkxOAaQ
/euGciCXnHiKYHFDhbITZUeEEM7sjcwVWb4CKFr8gAXlDCjy+R3y3f8VjljOCbui
sqlyU4LnMQTNd+xSEYuQfxEMigqC3tuYtCMdUJm2lshvVJkkdhOjNLGd2PMYsTE8
caQQJnZy3N0Rt5RDipVUhxY4NeIPfToPi2Lh/g7seyxmBmE5ztqw7gMm8PxBSEGm
T/yNFJrhRQJJBu8J09Iohi68pN/JXywtDT5T0v4TO4It9zR5Eth7Su5lGPTFYfT7
fFzBlR3XM0OldQOJom/Lh/tK8xwa2Hwk0C5V7EBc0pvUsbRR1kfeRWXondm1Oe7f
mvFLGsYsjPozZyhy2S+zPcYbY8aGNDzPRCWYbtp6umJWeZwTLtiyF8Tw1NhGjyhz
SbaoUxAeKsWq8+e7HsxnKVt9B2Fm2XH1hs9wVl+Lj5T8Xv3Zf44thI6ER8goN8zi
IJTLOq2QAQDQrTDX5b3xzuCg16go5oO1ZP78lQ6eNdR8Tyg3NMJhWL13HYTmx8kb
7BibVqx0NgNrYJtnQ/PBISmpDAc6jQEp8UKoiDUGDMDL1COh4gbFwWZCxMSA8NBx
iz5uI1PorUhKBByI9TnhxAsUW7dSgsetNzuyGb8plAEJZqQN4cbg3ruvql6qNYye
a6vzf5tsGxtO2jqreQ69COsABs6ia6gt1w9H+BYB6z0+IEsWV7cLB3iLfZHfuSG/
olQsFVMVdWfNLT2MapBRfjPDZrjeUWglJV9iXMRfJg5vHlhruI9EA8rZjqWaZoRM
ClXTV2ZB9YkV0FtDS12tLgHi94Xqki1q7qbfXRV2AArLNZFwipm8jn8OUbkEPF03
0raXvzevWdHbsBd8Fe7qRSzbMNAg/BN/d/TZefTC7ns8OHXr2lZ61+26svQKtzt9
AtWYIY2dQ3mLvsurgMbxViKB4qvg6MKYEtycCnIdtdiFqJeAt9l+KNcMFM5nzhaq
Hn5MTfY35kUeSLBMcf8DL5dU/riDFW5G8bV2adkuNQfakmjbzfg3JWs9u7FmXQG9
FXAYmAVEj5QpVv8jCRngiWycu+dZttg3GXbVhnHoRXYSoeVdG9IO2tc2lHp2L4lQ
ZCkZZa5wahbIxD95ddzRYqDLAuUZFEY9sjDZVraBZVnz4BsmU/R3ndt7ipD/Qqla
OIdfWOhxsj75LZvKG5BpkGUmsth49z/STJ9ZpDAaIYP0Eq1P4sJe9IMS59vtbHqX
p7xUGD6VfhQ0yjL8VFLb9xZW66IGvonEBG3FzGHCMr6DYxlcfSwIgtyGTQq2uKLE
ucht0RoHtdi5bEXcrxX6lv5mPNTe5r3RGlFqUuhuhC+kZxjoSPsBvp9WvNoprdKQ
WfFEXIsUEMD2p1Hq2naIPiWbsQyF9j487u8v9DqwXFv9rOTobTarxgS2Svg9/lnj
SbxcUdqgQorkiHWoePh+MkSeBY02II5Y3+DzT+6ZmyHNznVxi1vg/HjUHkGTKuiP
mNQPPKhUIwahHJWNG7UMTjnYErLFR3vzlwvWKyOWeTwyxYV5tjveuRGhUL6hbo0/
xXrg/VOP82CCTMfUakZs6Z2bG1MQuUxeUun/6aTLHIt/2b7UGG4IURvRhqIQGxsJ
X8nMMRILxxmrwOOFnJe68+Nm4P/X/ScWFOCQan9Gi0iXxjJpI4BYWwZG7xHNnrDH
NbYeBLvVfQ5CadslLvzsTaMOFaF7G/6DXwVJP1XdxVTzQvmXtoaAzwTNyWxmRAS+
y3FZ9jFSHOsQAykYkPiGc+9ELVbWlfQBYirWP3ADXRYtDczpSuWbNFatYyZlTaw6
9Ieu5MFBqCwSXrzQmxsTRgz7+gYZGXCIjshzruAFZU3JQ59ZOCTxPtRGF23unDQB
4bA1lLMGcq6aD1HQhhal/5Knak6wlORLf5nSJzDZ/tQ1wX/xJgzGaL7cyq1++RXc
PcA6hJeGTcHr8alSrqNzEJSdjRDl9ZM6qdb+IJJeXLgEewMU9Ie0z6iaHOA4PoGX
rw7tEobjuAdgCnHgOGmfg9DAwLT1MczY8CgeEUFcfbD4f98qSGLBiYXPbZBrVR9a
B8VfKrDgc4JEzwRsa+Ut28m/7CQVSzFb1Yp3rQ9741DXA6NCksUJup4zPuVVarik
SdL+Mw+28s1WFUTaPjNXJSCXQwYUmqASSBx1j5vzzvkmFu3krCXqu6zS0GpUsIfp
rhJ+dhR8zhdBAF5ZX/DjdwPrxXST+knTPuy4efd4cTuRPl87eIAFa0ajfPEFFdvI
93ilc25a/mrcV9wGCD+wsPTxp89M5El9E83LujQPmN71POVQTwywDcXx7o583lTK
at8X1IQHFPx3SSguuf4N92SQUfKXkoslLcXWeHCABY1NfAEylsVzpoqUqsPaN9LX
OlIvdAQL4mxU35/HN/prBMbYpxvmF86F5gLDCkRNifdK89Ztmk3RxAMPwjy2KbpA
da+s1kHXB+GiijqlSSAHMHGc5UAXQK+GjAxF70gSj6qbQZVBsqY+5Id4IpaRP1LW
JN7BybDIe4f6+Uwe4CcZ73a4MQehNWiVny9CrwbZX0OUvka1UXsEUESqLT5uCSKT
rE4jAriQZiOCg4AGJKNjKmWLwN86ogS/Tr1/Ut1p9pgsOOHnpNv6iL0dHmNEJzFy
e6Ju2hANm2zXNQLZNVdHHAnMBG1yCCStSDgsHvM76UKtnxd4jjycha1u9QmsGpGE
M/LvERr6AjutIP9XcsTxDdt50iXLLxaL8K4vQXM3hSk1dqCl5LjRjeaBJO6UD/9L
n/9zq+7nIQ6OSbPvlG/gYdIjEBCCBRPhew8sZoK1fFEhpipWr/n2+1E5GwRCRmY1
17C3kcTTnO2MBAvGEfE1j+vbN+n2sR/rMygsRieKOKu1LpnOTPRKjVvzyxiC1u6D
qaeek4IKrZE6uK3WgS+FDqR4jxmqneaWtKLcX7ODcXjO5Wqt5+njWMp1wnt2NRfm
v08Lxn+It+JU/rTCKWBnf1CPNnPRzS4SU5dYjSiC58r4LhGGbVARRTTenJndI9cg
T//9x9l/0RK0ijDxk2flZTLWH3e1y6qNVVaab+D2+HsqckV+HwO4pAAoeqko2eI4
Eym+PG5EmsOID3uMR9am60a5vTKD7X684dZWweBprZQNHxzA8DDLVatOoIdk+TGI
zPSiBBk72m+Zsj3McDCyO1mLOy4hTT7z7+ypJu8WsJYG7cLdxnglLqN14oF+tzCT
NyAJBNrRO+rFlT0XywE1wRI7GytpGGikxN8OLei5r7zpiPC+448VX6ggZ64xna5m
0znmMyhglHxu2iuCh90adczcSX8eeUCSfcyVN+YrivX4xXXWXhOyTZmkVFs3X2xD
k7j/NMByTm9o+aSaQGlMrIsbZvg6DFAAkaNe9QFWsDpPv+VPT+TpZkFQv3t7irQT
FCdIyNd0IkXHVe06bjaLFlnT8y0TomS/vKk+8lqO6mqgOpRxIN6CLb4KpBGV/60Y
IOhz3XG1LTp3JQzEmQL1atL3+o+1UQ+BYy7E0UqL0EP3rZeJ0sI3yjIUb2/TKHY4
3t5hkUzi9aZVYW/nRuiz6bzXU5FBvjBj0OMk8ur8dbpMNYCpFibBbH/PWt6/ta6Y
z6jERzSOv5j/XFHz1h6dEOVUOMK3Vcin0SNKf6v8dZtB55h0YWjuKQZiYvXG55Q2
0AbiKiVMRCAptSAI7vgErwLXKL2EhABKzjBjXYFn/1uXmNjQrqkLT06HNzPjnE2/
dm9W+2q1ZMSoeHjod0b54vnG1CMnSjxzM7WVdYofRNZU1CeCXKG0/n32poX+Zykk
0dY2eZunAN4gp8r4zfJjHGATTUVdeJI19Ag1a4fltxbTmz9V3NqLvKXHQH+kCv6W
LKesd8sj/G5zeG0Xbo+Bd5Ce3CHC5lZe6g4TUblT8ctKnDhfZt1f3VOrnE3rttrm
JNuL5dIBDkI4HYmVJ6mOWQ7u4s3ojTTl9ERJqfu/l68+GQH+QBObgUFSnvAKSSMg
i+Fpda00IcvPr9OdbeYyq0pkq/Y2txHxtPRYGwlXX/umiVCJKu6xbcMiflDzG8yK
rcJsPpLxNV9vCOZdVEv39GqfK4FiTH6oeuM8Wwg9KrmEwY35pcL3399J8x14FuB3
Oxr1vbw73F5Ik9pTK/4aAMI8tbcgnj4MTGdQ8k0qFVSbDVyPwMZ66ehLOYkp9Fyv
o9DNf7FwzBnxa1S+KWiJA3YdOhIU/fT5esODfNCzLiLMj2B+yVbYwtBKGKfnLNAK
I5srFt+3Bzh4TcLuN+8FjGL002pzGzGKorqQ/ImTN5/VNJArdg06lN3hOsVrivaS
CInguAbNFPI0v9fIEFPowl7Mha+SxzarHdoYHSSqnDOw8QgbFeGBIR1Rbrt1/tDN
TVDX030eeqtrqspmpuSrktnrk/T4OryHtiaV0rzSnzkXzLoh1fTl7sUX4MDrlXq2
6Rd4BAAAwqCXgmQ0p9TCFom78qq/DBjW6j35wQMcZa2+hrhJLg/OZ1YHk6xpRl+R
9CwLfUuKQZNlgr1NCa+tFdRxAq7yco+59e2RcR3K/zLfnx6yDKTjaML0YsUXfx9u
QvKJ6j0G6Q4H9m8TeJ3AqdKmGBBla/j4NfQnC6h2q1IKJUDytNY/g1sNSBZ2RPl8
rgzBvHMS/66b1Ld+JNOWNNv3glzsikIXRc3rCMsn8QHtuB1fvIp0eg12zS87FC4p
+/jdOzGCVzyA/k++kqQslF0LDX8v80rbfgmpgHoVVcFqBRZ60O8Nczn5fz6sRP39
J0EJ4Gqik8HEuL0kk+adDdPNiWEqiGMvj9Qpt6o1V7VqsTfZ3fJY5vXaWKqO3KH7
f6v0DjOKzIfDKGJiYlqWjxYY3JfIhyRGwN9g4+fFxVxpr6FbmM3xM0VNRwWJRxk8
lky1Ne+35UoKCnSrzFF+nc1j0ttXa68ICwlsbqP9Aaayqx8W5FU7eMAAJIOKLgcX
aEEPqQisn8A1cB2V98DtMVcY2PvX0Ey6VXyxbQJX3pHnEXiWFzkyHgXjjfdRAbYx
uPF44D9SJ9TjXjTEvKAM7PpPNkA5n3axolVv7T9RdnE8oDD6bm8/9Y5nnPhGGRG/
on/GvQ8L4KkVM8bSs1xuzYngfKuGmwgcLjqsw/e7ZEmvZ76FoSlojrgHzN4+K1sb
gP7nMeC1weqx5tMBgkoDSI2mUK1n5xOG8lLHa0VGJgwM6hTF7FHsWIO9efro8oOY
vHtSsjzdnHUYGAcNLaxCtFMS3o5adNUzkbvGLKH2UuNZTUGOKUbU64M/6sEzFo+p
vjzWhYUrylOkzArY048TlWmAxL2FBZWJPbf7cH8gJwnpUXwr9gs426tpn51Alkbo
4CdzaR89Hecjobi3PEVw/YDSXkspp73ZOLh/AZdN+KGrcFr/koePHXJEwT2i1D9A
zLeTqDimxZfvlFHX6a4SWbvYRBhbN8cpRelQkfi5CZRyILJ0x9JxPVMmZY5z7dnu
AhOSYeXUebYjwP0MAaB3UCpSCcqfF84fcGNTT0mnHAqCFHP18/LE6Z7H+n5rPEf7
7lniSYz+i53ZqPT70MSeIl8C4/b4tNZz/mf3+rQE8Wf8XQ1CTZaf1YUiNvP3/go9
HyBFPBi8qqUuhav2pBX6NJ069GIr9bktPBZ5EF5MeeMr9jIOBEo3YHWurfT+zgsk
v74JqMdQ1dO1p24oL39h6cwKkoNAfY6wgCNQrOgx4RBZjJVE1/cK6dELJrW1in7d
fxb446ztAUgYkDH1mfeuwa6blcjUOyux3Ma1c6vvtPa3i7cCQ5jWGbx2BA9I+qd7
MDguIScIsXOyuCrRiSLISNQexme1tP+dn/RRTl9dxU44NmAIbxq8hhYX7X7drHnw
LPo9iU0XVUCSqRD4spTZhnsXnhUSK0LqKX2MaSVO688aiiBHkOk9YmBJN/iUwXBY
XIOR4iB2Q6Z0KCzzq2434/NNWn9W6pqla+cUEneGZfLExpjYIT3iIow/nBKnZK9F
xPjYzAiIQg+Ea3t7JAMVaN5XNecvjvEoAtk/m3xhEnIeBUcWQ6Mk5qH+tXccFkzI
nGcmAzqLyZb4+W6SwaQi/xTzjSPOgh5uBlNJm/203No3u6a7lI1+a3H1ZFgtQnA8
inCAn8CcEMHgK9VkVYfdFBZGFDaLjr6O7KTmr9RHBKHGd9QIx3xjw6HmZxpCc7HU
w10MhczZUKghM7CL/Ch1OIiiSYg1OrZSddJFVykvHk4ln/vlWUty0TugREGMvY0H
V2nTjrhmhan8P+i6JSvLSeN046a5n7fSSYl77/EPcAkHUgKL3DSAOn/gt2bqF74z
klCX2xAae4hUpshPffAYhOxiEU1b0YbqJYlNALL9ZQO0WusrxKCbkS6x8F14pp+c
7TmnNxhu5l8lUWtu+pCLwqIE8GET9aGO6iqHFNvG6EiZnCHqCsxK5QWe/46953h6
8NBvJMIEas2yCianlguvpYI094tCuE/A73xS5JqPMcfxWWVExV30mT0Wmai2wBJv
RStNtNxiIi5WHBCAr/CbzIxC4P5DC9Erdpismwwe3XjZ2MReXTNO36RH66gl1JVY
UOBJL6Womr9N/49xfnMfyQZs1l14BQR/DjR3rGRnaQjjqQdzmO8G279IH6MPjTdr
U+5RCDdbs5f2esWclQnV1qh+s/ICtlaBMSeN+izJu6WazgiwDHmsFQHRCvvluitS
FvrvAhUNMYnCOUHEHvahe/gtEHM/XxJc9e9IdsL7C2Fzzb3/hL1/kVz9rgAVaJfv
O+YGjnKVYNx9jtMFIwjBaKvn7XFwvniVQk8/NEddlvCbkZ7i/z/ndOpMoQUGR0pG
mg+gkBf4IZ7rEBR6sVcxO9d6NrkgP7s+uXGEoXVFbSMxNFFLtboHKMsUH97VKb3c
N5SUCfOTceuCZpy4046YiDvy13Xt6t0W0ivUxqd9V+WJSxEGiBcAktNgqJ2pKhdf
ubvapjuprIL5+rWzbIJe95jTqcdHExyAiDToEKlZnq69JBGt5zlNPWl/SOfWU3fB
rb5fubTOU7oblum9+RZfFxgbcjG4WIZ2iVguisNcRhZYPAdS0KTN1Wa7pC2BK6kJ
GYIkTqFr+5dBIhdxewA3004cQ7s9JEBRExay7rKP3QAdYTe01zT4wag/xvfr9W/f
v/yfQF81l6TL3SnkgQfn5wV1XSHSICW83wam7wNBDKvzT/63nlYn2r5/6wSvQsWT
Sdt1WnZiqXZahVk/+QjyRW3wbmY1UlrU1xFfDrE/1nJjN1o0kDZ+qFW0ai+JSCyD
UarXCddvWir9XXxeFnPV4dSO8a6V4kFp1wcPk9DLonA4L/QAU8/nIxSmJh2lZAlM
7RRW3m/mY1frxa+iuSMEvM5I78+cdcmMj9UO/4y6zNdONF6XRTkmB8r5NVWEtar4
oo6rTjPMm2M/AKSFbpSyoyABoxg8FciGwMVOb4gwqUEp7PDfTIn/t5XTkzAkFgbf
4+p/2LmZXcaCJtpgSD2UrRYIniJXD8nYYnF5th9g0RrUevHwl1ceTZy5tJxrUooI
jQtJzIIHZjBSnJsAoKmu2DHU3cNRXetpOTavxttZxAf8M/B237lN0lxkft/0FtGd
YUWNmI71ACb68reruXJQnLb34jEbpON0tG1VDGQurHVOywtn2SRFWd0ita4lDwFL
pQSRPu6RrRjF3woJ6P0a2hqlUHltduQrZKiS8J0S7Z5C50Wzq+sJE3ShLjsJD+DL
/ac6qU1UWpYL0iqcciME9cEzHFd0fcHv4kFwB0yKi4QzJEAM986xladzZAjZ4ZXI
USJjMzakV8DYw7shLqMKZt8kIwQTwQ69mInyfGQg1i7cqlS63BBVYxXWaIuzrl2a
4UwbUKRXF2Rca8w27kMAqcbLXt0IuRekn99riG3e9JcKUY4CQO7eSkNxpDr+Ry84
o6YimZwsrCn6JOsT98Ici9m04/O3rWRrAMsT86iF0yqFkk5x7c9JWIGE/OpGZSJS
pduRSvOkUVAkizzVITJ8+kZVebI4W7IMKuFaDO775dl+xJzqorl/FSJMv76srnqF
wlG+mgRPqMM97nn8P8BarymjM4pAGvABcuzTANbj3EEq8HLKNlwz/v3q64NQaUx/
iX8MoiobTWiTgcxym8quat5EwlKpnMJm2Ep/gaMt/2TtRXhQ1bwY9kwEI92EoS39
cGmNq1ind7FO6N4qdP1KlA6p/fBQ2vTVzRVL0kqvelSOjURNCGq8EWc/T6taS8D8
svCSfVYpJqp37VLV5oNpQ5/5pN8XvTD+6IyPXoXH9FFrhTOj+201gaJeheMnAQV+
M0hpbCj7AVILuxE2o/bRiziBBen7GPohejMi8BXF3NCLaMKoZWgS8nQ6rkjJZ41V
aDTe9yL/L1Rv6WHeYXD6QmubbAQ5ajlF9Jfc4qV5MRjGxLNai6fYipAZF8auHdEm
ee+kilym++vlaLtOhf5Y9JFfpRGiMton9wh1KHys1huoRd6lYMhQvxDcsIelAGgs
s9kXl+bzkHgX+TOxzFOV1rguhisN2n6Z0TjiCO2V50y9j7cSNvSrnLLWn4GaILY0
4OzFUBu0cYYcEthnZytdjs9H5o9ehhFbzVnCDUFYd8KEvu+TN9VCgxhkJOc2Z/r+
69es5SboP0XOmHVl+B2i7KFDccexLwOZfN4NcL0Z+OeIsWOyOweJWNpHEV2lIcGn
x6TDuyK3iJo48TrVzGxkU2mZHxMOSH4v4dF2Se3KMB4AEFqRsA8cH60bN3pN1oxJ
DVa6V7wqnGvkKBb6b5izhfE/Mtb9fPcrL/oxCee8x4YROAJ1Ldeirq1GyZeAqz93
17//VqythpO8UOwVa/xObQhcvT9MwU3ZwHladbc//hgTyk4uRQrTOD6AgOO/uSis
w5WpO26yJL1SEy8rhukwI6fFvAjeL1KAcxKdlf2ASrPV5vyqjmN4O/f+p1pGQwcD
jCsOgm0l6RR7mD1kg1CoGZLAKOAcTnAlAatjzuN47JIY362pBH0UzXzB1bXDdWuN
KutfvdiQu5y0+1tZ71bhqVVaWJfoZbfScsjc2MN1TyKkVo9V+nr6dTzLcAj8L59w
7WJ2mUPiiSSso5zpijH5UpiyyQnR8jvR0AM9pYgo9tDvsPkSq2xPTTM3atOKfx4L
Uv64Kh622jQwey0dT9OJCktlnOEr82doI73KB3wW5hITWgwj+F78TRBKncmebgMV
q67RShUrEmC5O8/5k6WLuNS8YlmFM6D0W03KJABif47nBftJRHtivdFa28dbUrJo
KBbYJ56qUxOpKzRWSzDomTDx/21aT8T/oyfmLiVUvgpouqlRXfjQSUCZTEEAZvlo
qh2/zX954sTXtFizn1WaU4tyLd+PpBRKp7d5DjveVgaDR92O7rczFFhqEyCwap6J
d9NAzVnzibhgRqtQYxtMYIyuJixQQh8NIZV4ZK7e8/l1dJuNaDyt7H4xhL+6CX3P
KQzMt/OMCHM0cVgbTFZgZfoX1SmR77m3uqG/ip6J+7hhYrFH8YfYRGI39UiSEqAm
vBkr8QeiQxmH1zk6aWZWJGwx+IBD1I1Z9Rxoe2e/0oHUEXUIcvXEgQb6+OgYTVG/
rRv3/406x7KnjbdwZYgbaCaIneg1wSTzDHY3u/25RGOk9e/Re0N2EHf6+8csYwS6
zOrH/pJIS/QhCav4eGMmzFWs9OtjX4/oVe0DjnhtgGQw/4+D0q8GIUKL4MIqd2fM
EoW4LMhYybkUNnWR7pQGFq4keum28ywpu/IfYlkd0XmtItyC78iL8Za4wyIEky/u
6ghqz/3co0A+MKFUPP9zSPgSLmH9pidMllXdIfR0KGWQR/YYtuADife2EyWUpPfk
1adkJ/zlyBiBoxkSMBSyaU+0wVRZoU74oufvmFBdmqovq07OsSBDyl+u7ydQi8ir
+1mOS++TPZeCeKwgI/C5qLE79LOWnzUv+tE+mXbCz2Ur9z3C/NgrRvTGF0aYv9a6
S0y43cOfeNN886M+CDm5zmOOc/zNpK1C61RVwklQGuwH341VOj0YSXOufQ4ln7DE
Dbb7x5jeZxIL9kdSLT7hEGuCB/MZwOd1dQ05CF7pyxTZiUsc/XPPSYvtsZt73unW
1VLQLYsHPxY45NHQkcSnALpudLqT+Acieh0v6RTapWfNf4M1NSGr7Cm00iv4qyQD
sbz/j0NaOasJXtOuGWfLKFzv4OJnFXAJdNw4MtsGYuI3CwxXOTCmPkAKFvNvPdtt
Y415Uac6ldVcvpEGcE4XJjH8CTcYQTwrffUFHMbWL3QUGk0AnVHUlS6xoiqaAzjc
Ej4Zdsj9GnQMbtV6oGqi36Hso8UOKbEJT1a/Iv+vp+dDNJNnYTstoNezP4C7GU5i
4RESy4sRyxSWoPCq9gmrsv71evy09bLtpKa3ltJrmCU5bwYKIWHvb87MHoV6QqEP
qoxWAk+uwsHZVlMZZhGUKZzWDAo7G0ab8N9CItro5OKQYabja75tG0p3GhgMiYt4
MFtekckfsTk2aOsOBYJJaNpnXZLG899yqmNVyROfLSbeD3/UGXjJQBTxcr8aGRjA
LWoxZMJdfSnmRuOBAXnIxtv2v7sQ/qv79XuzMSqDGWZN6dHtDhTSeHupBSlrU3Ds
l+6MFdSmvAciG6eVLjwt2YAiOpimOF63cOJ3p4frTW41Vwh+En9DlATd+0ESwZPt
yk5F7vAbz3+E4tC2FmkCfpPOqf7hClMHI/cBOgRiSQbAtDuLcDWOxR+K3LDVaVib
yTXWCoZUbBRUDUKmDoBAqZqLnmNqPb/FD75UbHaHebya2wu3IA0q+DFNpLGZj7Cz
7X9HXvSUmNgtei/XaAzVdpj+IlE8QFV//JUU5fCfnI54cC7YLsxo/1mJoxi/Y1Of
ldTlzyyjRxhVNUCH3CHZ4JgAD0ib/09MqtXP0ZEm2zOIv2+vazU1MnOe9L54EOSB
SNDKea9XGP2si4lpJxeNruGGlWR66WYlfOOxJVcCbxtROBlQV+EZ5G7HAfY4r7HD
9qkjcjix0dbVx6w4xz3vCMiEnNKblAOL0G4Jy10RfgfanmakGpbLZ//cSHqxpm4L
MbawtAjhuwTb+VkMZ3AhitfXbl8rpmaCOVSalcGQojd1dmmROV1G8t1h3rkW5OJW
WSr6EueUtzNKfo3wGb7ZBeiVpuj70T9zPbkOqtMKTHxfXQORW7fKtfKiyuBbK4Dr
8Y2JiO5pTdmJCkH+C+Zb0d2YzQG392FkwIppSU8fxpq7hh12FMaZBGCdOi+1jIlX
qEYg0xT/oRsF+XjLJPXBOy5z5UhO6ojqWb242BTPgpW8CLiYy1cyHAiiTg6XC+N6
gt+diPLnEp4hXHTprVfJ+H85/0ah/w9cy01gUKWrjMVMpwxJM1mkKCxVPpoAwkRi
lOPHWJ2GbvCfgqu810hc0/7fQxQRCXmq2iv/RLV/fyASoGfkgzT6tDzefAuL44ht
AEBs//SLXNPQQKjcC6FzlXZkq7rga5gyzoByOSKpC+FISyJCLh9I0tmePwp+Is7k
/KGcsvrCBrlAuLgp40pJHXLp50gyRQQ9SAl9X4nLxVERtJQHa7O/VvCLn4HmEX8I
hJJVWq2OWK9RlJGawQayoFRxZA0gEf8LJzds9QuhHHqfF64ZrM/KLHrKovdu1fPA
kvQVGWpFjbtSqjWwk5ljV+MflN6WQ2a0sUkX33b2F/nOF48oQSWZWO5RpnZFIf91
oiSPK8lvj47/70GC1JOzfRjNCcslWq/xTSGx9BGRTnvnJBG23nYP2y6huMiS9pt7
Bdnb8JvdfpKM2CnyZw/trrcdwteoaRgxgCp3CHxsIx7rbzDi3dhTcxjGzMHY5oKj
X1gsCHJ7uS8q3E9Ady/JQz67Y6l1I0THTqXnPVephIjLrvbpXnm9tn/UgDPJztzQ
6pGWTcHG4NUVBo5WkqSwb3veCeEYF/exUIvZd76Nj3D4zr8HYmV01OqtmPo20Ji9
6S+Tz/82wnQwJrV/zfrKGt895QvH9tIBrIIHgH+4as9zFdbzbPcqNxz4O0W1PPZp
fO385Yijkaf/9pnn08lJmg7xFDv2vgyW2Tz0fl6ujYmuPykRIjqOfNsOXZUSLSYR
PrRCnnNkgD6L3XdC9z0dHc5+EQLjJ3spLQnVX1+ahohiXXx3h7wLxVH8uQaxvvYx
w6c4aLMvysqUgXv7355L9Ce1jsbn6F8lB5PfSWxKRL2R2lUCPSsC8ePQs0aWAzd2
SPze0EryNN7GEXJXdsy5dMyUfpw2QsaXPlEI8KGT+Z7Fvg13SsY92waQqadsGmay
h5LMLaY8zMC2TSyaA80aWuXZuJPxtxhtoam9WKckKbvxRsuZ3RHJncGbUlHva4PT
pIvOcITluHBYLlZPyQBktRWRjaHASrm45xrh4agLmrmNqKm9zASnxd2QQmLMv0nl
FRAY+xIDhXBWxu93JfLzGcILuAIS5dKhVj1790GxVP4Oq1I8VHAYC5vUjPC8Nquh
ZXYByga3n7HIEIfrGI9pWoVls8PMBdezXVxRLKhkC1bUL//Ypo3NM0dYzzeHjsJj
57fwe/gGhXUTTN150gjwxa5Hec2G0ORrYlQbP09xDgiqF+4L0hlr2DIW35C5w3Jd
u1ATWxJVc7ZkAJEfUzOnTtE+OrKG0+0QYjmKtaWblQn81K1Roh9ys0rtMZufv4mL
sbzyOx7+0LGZ8mMuTD+PUBAg/cha4FOs42N9Mgr8NEDJ+0gVUTpxjmK+KzaFrXGC
IYNjiPMay6XNn+TgVeAvbFwQe3cKZLb0Twm2fuhzw6lSj2fbBZ06NOs9Rt9dAZIQ
fEVZxta3tk7mL8fLRxIcs5U7l891Nca930g+dyECysY/KAHI2DLnAy2YOwubPK5k
VUBmBqS4Qx1FzAkVzP7IH7zDloViYBrT6hlYp1d6vBhPAoArZjBugQknVnvO5mYb
VjjNrWeOb8P0ORzzbR2W0hDjR2ai2/LjLGTmRUN0Bv3gbflsETqduqLa85NJBDky
qA8ChnIRSCtpionKf5CV41NQNafZroepNaH+btdYTEb5RhQJ7ThvflKtFvGtWEcn
l55HI5xRczbKb360IbbScGwg5cjhTPmZ2q3pFkH7fMIMfj1IOn0fRoqzf7UQEUCi
2hQIiws/CqjL1IEpgCmhqGDj7EXAODWgZaS1lbiZjSNwd2ajJl8bFedUbhN2SvPN
3T1Y2tv0kvzFgF1XzmY0W3laU5TZclimmChkJklMQzX1UGre7lqcgfc2x+IQFoSJ
ODCHwHdTj1ZjJVgfKpy7CPJ6+ys/zeHGuAVBQQCwnszb+dS35ekz8SiALwrOL+4f
RzW+8Wm28Rj4D+pJ87oESoeUQ2hIBSAHT1GB7z9XPqGL+/J0C4WGNKU5q65IkdtN
r4pq/w3ZMAYOPhKcOddUVIEuBhG8mfawmUUh0QOELYnKQ4CXC8skh4zKiZLPmduJ
nAXoanMn360xN8attUgh6SgvABZP2FGsd9+IlWihXT8+JXnxK3kIHVb9OIRJZdlr
6lW0K5DFuBYiKW/B1P0FIiHw5Vp+7g/i6wFOJO6zG81pa1KaoS0X80kigwoBWvPE
4eThsqFMDX1QPu4xkfpVsMJaKKIRlZ9awFdapY3scoOFY9GeWfx7r90Ww4aFWM2+
10RWelBdL/cSaPHO23HRLsRRQ433IR0AH8VWM412Z/IrFomwfOnXNWuOrdlStbuP
41H8on3a0i0Qkge3rDXt3zRZ2/SVr1VrsZOGJV6INnYl5NVTrkE/BJ7ovSSuAmI3
ulpXGun8V/SzZFGk+/831DtLr+AQS8vr9w51i69MTaDozGE+ML49ccl/uD74uvi2
DlVvf6GUdpQHJWAeuni8QHO7HFHC7ysU1zwSeltB/l7K/lqrHt2tWIkRwXt//VTf
XwY6Luk+mPJ5Ze05PwpT3TImrTy7g8+3Q+tU6uqX7qrs3lREib8LAPUzRuTIDj2m
GSugTw15dkRbGQ6YvVZkrhVTHbbOOTc17ztWWHCTGFIRDF7r5mSs1GHKO0Fjfs0Z
zFox028h34dP+J+6trCNxDlhsvxg3JWhkESmptr/CGvLC7KPAQ0obDFjkrlH18N+
ObJUov1R0A3x5CMSTdlOJ6t8L+/tT+me/chfS2P84zOZzEvxji7sTpkSdXNRCO5O
zEPX8H9O8EwQ+ZGjK/YS44kOBixz5yo3Asy1HY79FJ6M9OPjGPS53RsvVJII4oLs
f4EN1cPEqjMIacUKIOqMOWriovmB4ZrVICkFeCp1hvvOYip8GOGyPTvnYANgqvud
iLnV7uiIA5yiofC7fwLi1pLZBcVZcno9yN30cxzKxY9bpqDi/x4WDq37UC+no8Y1
86NY9ONW7FmG6cZq5hyHLFh4slcc5kuHythk1rvU5WA4FJX8cvZ6E13QIU4F9MMO
mjux07nfP7y4Db7g8v50waHBjBFy0P74xXEfx3bpC2crKF/puHCuwyB5kPdcHaOI
ZjOnQWFbtu4miXtjIZW77+pctZuHnNZvjLQYLr1okRkwCGkdJGLID0LyuGWEIlrr
8zbKVw+eXQ9cvF6xpeOpEhc30Lo3dEvs5FwJyNhZLJuCZI2fr9uA3WBMfEammh8K
zwhbJ932wGLGkOdLrKcK44QcNHaPBA2kr/0DOK062LE+vIxZpMf0NjYUaGBY5MRY
znpcwPr6HicuiLmROBx2flX5/mdKj1JFXwAkDyDlcRGiU1oGkahsp4cCcDxCxGE9
WsBsAx7JCxiO6zxQdGBw99viMazjid/Ji/UKhPToUDKMx5iJTGIse2v2ULeTI3c2
AYRh6CzQ6lIT72AxlIx67AKFzDDSFTwnbf8Cf9lnQJzrMGaXTejS6gfe84kmWCXV
zsXOXjYFRCDuUFEOWm2iBKJA9L4eKgSLVAKpZpdTuDAyBhA5MvT6GAFBU1XAshyD
h7ex+DSjHwLhGeYMZf4ZXIrTfMDdSoipekVMZ5mn33uzY6HAz/hzgsI4zttQfcTP
443AdYSkgJPFqIcA9r8tHMFiy5Iq409vq7qXZMn4xWp+L5S4gUmher31bKxPfE6z
FtI0K4ZdG2GYy7yJf29/TZHKqP803UMJX1lsdbgV5lo4FW9QQ0s8MpyUN+6VkdMs
rkepE8GfChDmSypXDjjCBhbI5+wriDR8558DS1s6IlZfyDAJJDGzmaGyzo20pQOG
UZ5CgFBlUi3gcUnEBdDf6QtEOfW1UvG3FR7FOKcwIDp3eeSUWSNJNmAcd2gdMndS
3cBpIhHWyri/V9r4oHbMQVPwCQ61VB/1IIMXtb45afAPx4d0sECEC7j/NW14HmSS
rqZX1pSeECxy7dwk4SFQK2Ijj9NhCNeLBHBrXAYvImTnj5weFRpl8FF5o2Gh6zW2
KEBa9Alhj5TBMKAMHjzheohBHcHt/+EbBmo/6lrRHD8bNVpMGZKtVTeufVMUb2S2
wBf/5f+giTvfw3w1w3Jx63QppHSc/aH2Zu9zL0WxfXK6tjZ3CzECakRIA45oL3DW
bnOuFu/gjK+qrl29lBx/rktU8GG+VueEFBT/ds02pRLAjBYrA4h8JHYdbJSobF9U
Dobn6FQjxE5mLYYKXEoOo9lRsqHK9OkSWj3TF5LzkGiorwMEUtM6s3ceXMjl5tyZ
ESIuFqqCxWr4Q8acUAIFLRalMreI9zsyWXVkdUmcDOJh2RM3JjLoJXHalg2zzkcZ
M3Gztezab50izbH2FvrcnQdXF/wfwD5IHwT3zUklGNfzfHAEb38+hOKDlcAPFVP1
UcmPh9o8T31Z4urM39lI9chZOSaBDXB2/1uj2+mdk8kuwUDDW4hrRkUCTFi8/Kjv
/WIWXs6TFShrW5WrnDC8AOYGwzO9jT1po8vHSLu267ehv3uBemDE0zA+P3oRr7+d
MSRvxMuQKW8KYmTbqAf1zvY9jqo+Lo30582Br8k9fgcpRSY5jymGm/jI56wGsDJk
Fu38dA+qpXxTz0NVoTtB1MbuzROY8BPw8TRg1wcZ+ldAZKR8Z0jR94cvRXY/pUVy
XOEDKaxB1kSA+1bcTQ1ErWu9dy/MQpXPvxwep2SM5LS1Byl240TETyvM2UZVRKW5
ZV9rdBxEi9l5KphfRHPhbrG9PyyH4azuNRlAdhno2Alk2ySxnfFJzHG1zJ9xL26L
vP+Ir/QzGYMh/lk1vvrHQOSTIuipVCK6QLnohfqEchyT+rMmsi+KDkUNXiirLZiu
+U+/yrGlNg47ulgXGGGs/cq4cnIelBjeR0YqZ6hn2LAnkGNhbIdWWOfgrOTMvJmI
rv82CY2TEskI5+YPQRheCJlj1QoZzjFpBJia+If77hvbeqo49pJTRYgu9FaOSgVv
R3+c76g+FhfJBvR4toqZiB1rZBdsTfc983FzETtefbV9NkbOquaEdBUQWYgsu+vd
Fby+5Tbc78gnUAtkRam91jmmi88JhETNbG1MfVv9oJJGEHB2pK1RTPlBGwJbG0mF
Vk1KsTN7RjE3ND+xk9ON+td+q+aCOkKIQ9BCZyztkNie0XHV5VTkArNVUeC4naAB
Tng/8wEQwziqLTMfvktStCtRchA3u8x5a95ASQ7cljpfgkcDwk4LYob8fC37z3qL
XHbhQP4RHEhNBDiuxGLUOAJmxaqoTwHpG3xcO8HLtpx2BE6nOXDJC8BdiLbFc958
9inPKjfP99JoOiyt1HtrPnAovdThTKJ5U8Teoi+rqzXKAAL7XSEXtEy+XeG4qXzY
Fc7uU4qoiWevfbH7wyVmYE1mBXaPQFx56cIpArE771A8hWAIscX4AUxIr4pYfIe3
Cd9UhTtdsu97JDVDziySX4YC6dZlDy3An5bDhSUFe7fJDAZi5QKCi6BEPfO7ODRm
3HZVbEafX2MCf6acOQbBi5bZgPgakB+cP1nqLURQ/ocYdqnrsTTFexFJV7DaZVq4
OiCSPmBqrjy/PXdJMtKx5TLReU2rrZ+m9N+RzDQoMAOR+5uofsyPTrpshm/btism
Yye42XGGOcTxdcrKnUUCFEBUt+E+4Uhle7h5DABhphUL2PkUajPFhfu8egnhs5iB
AwvYEmkc1w3kEVyrFXexol5idG5Xwi6yrrWdrwHULWy3jlBFESne+sXll7SNO//W
ffymFlGs7akrCIN/RWh/9OhMdQfWnuyZvAmZ34pKAzXUtDxbcx64+aYJbmT3UMsH
M1GPK/M5sb6d/4rOv2d+rV+GE98bzudZzZ2h2Mol8zebokOFH4w4QWLRDEcn592q
nqMWt7UvpXizUJ8sIRUX2tkyCX8P5Sne+IIaKtSfKg83nSF/nLjgIYVL6LsxdyWN
BxrH0dKoRbYsarTSxnm1v6717x6lpcVO3595554zT2RHHFxGRNTJwhe35ji0aAqg
MezgT0WhPKDbJWcUuTIUI83eIIaDTv5dSq4OuekZYTQahH9IkQS+Y4U6cmsdtbGv
hv8LRlmMWUEx1TB7be2Ig6gIPs4tGUyI0lW8C3xGLsDMqosRB6/yebxRsjxVWQqF
7SAj9c0aWebaEr2/xBtQ4MV9lKZAgrsnyfTmxvIDfWiDDqrHLlpTOcVsRJcBxCRW
kOn+q7j9ig3x1Dxy3TNsqG00S8Bs/t83M4GRnTADhXNc+YG3p0roegWQT6wM0Ta/
Uft/55U3lVhAf0jC+cFLeitwNhEwM9b64l7uNbKKUXNlsISUg979Yhf/M5f56ayv
aOnt2EGeW52syltZwmy3hVfxuiFukj6opaR5Pl47V2a19TH7hx2ldGfoZmFDpe8n
FH4RlY8ce5HMtgrz0eOwAHnAcTWTrQV7kL31h+3UKp4N6fy7G7QK5SkVoykiz/5Q
NVUIUOGQyYm2YAQmEugIzspP/Xgj19YvU2Vh13gEtKg55B/YrRhEh0hNHaxF2e8f
KKh6k2hVGl5iCCbAvpVjCVwaXO1eAXE2KR+W6Aajd9m61cy1PWVKdB/LgTDVF7O/
lGhrsnXDRJ03QujMW1Q6Zs8ZRg9ttqnswj3KQYb2aJOdKdFMzWR1QjMYR/FhJJoB
0za9Vva3vcfCDM8vYVSnQbXHSbwAtEDFFuS9b4nFTFsSlLi3JpeKBHC2H9WE2N4Z
ofuzQKq672YqJeExNRH0kjApQaBU8tvPu/4JEbBjeSzOi7v6bCIawKHb5T6+zSaq
86GUnkbdJ6Y+bFCnwAAefbacRPDUK/s6SwMJo8JlzSW8NF7koMx0CgIJcsdW2dUC
X2XZi8tngUpERsdiJ/pa8XTS4fkazh7gRs36fERIbnT1NrbLN05oMPtYUQofPCLv
BKi0Ks9B1rdnF2vbVleFe8lwYmd3SeddFic1C54eueuIjOXxPuRr5L1AW9KLI7MU
YHbBs0qqpasxBZ9Nk7jbkvMkzqpmmfW7QgkuGP9925GatxkgNtALtmXeGPjvWaqv
3XnYuSkmz2/5ATfAf7a8sh6B+rv4ZwUEtWbesI0MoC2u5sQ2Z09ykgMXZYKXIpUQ
6fhYTagH3FBFbRb2HWDvTNn2PBpUImlVosA9NMYG6CapzbxEALir/L0hOlUeSmOZ
RjkYuoJMpjbiTVZqZvCSMLX8THwyWkt4ea/C2Njak/3kclXrxpQpIU/lfsUjiv3j
f659/wTIAjYh6+m0H8dIXL2GBhsas2hKbiZ7UzWa2Z5gj0QnJoUaXhfB92jTPgqm
xYNsnFh80b0V4R1yfYnb6WBuDWbPP0SSkKLAXurVh1DPpodTmLBjFW2P+rGW2svf
FqMcFYrxOchYJqzhrcJkisTQufXin15iXvTUZoleFHAE42qqrvZAQstJM/Kf3/UG
0jGEnGm3UHD3W5ga159CwXXJY7n5ga/kFXNjaPaKxI/oD/ltQRNHA1VWCyNsdYJV
KSfn8Hqp14qRMZzrBxjoBqjM/8Fi7Fq9xHGD0Sa62wlttsApFhZ2kPRxQfJhEpNU
7c1UGOw26dK083E5Kb7116Y9ML6lDzzsT2Oux5DWF+d+EAWOMST424M/SUznWZIQ
cejCMGHFdSj9kQU448LqcLkhFanfOXwAFRDfSG4CvKIC+cEBz6736/IXz31qGs+P
P2rf3+Bnq7ih+mCPuJaZFp3wFAv0x0KiTuJt6j2hZQwjN51MTPdxyAbYhvIFqy/K
dkJkhOB3+TUZ/SWoBpS+6qq0AlHF7ynOBKZFMSUzOKSL/SU8gzWP15gWMaZw7x9d
1KqW6MSqsfj9qLJEuJzlQSZdSGoLr6uxT1K9njayIsynQWtNo7BAAgToOgqz7Z2k
F078nkvEWmCtzRSx1yZEqkYnOxvEUGppq+dfK0u/5o+RsQOCh4Il4etxpHc8hVk3
0EsmyaJDm9pJ8wylc79mgkU6KYpYuZht0O52faXK1qzZeLEpSmwK2kY27BdscEKA
AzDzSvK+Hla5BrpL/7//J6ESxnESuXE711akQyVAfEyoV8O+Kt76WuLaZpU1v5IL
P4nSTdbNKij/ViSoLDNQ26meWdnXwGl7ghkH2f+wt4fBlNTmJiDPUx8zFTb95KNq
QkQBArgRLre0u7pu51cG8M7Wu22l59i0FcpUtjI83RHiyn/Ynbx/mR5L635vnvZp
mSQe5AhJwyY7xKPtvACtrY2wKZ+R7c7hRboNXaGBaOTaMrBErJtW798Gy0PJ7piS
g9s2uVSLQkEjbeOhkdE0/YgiksIfekxIp4N9KdhQK6kWXUDh6DEC68UaHqVMatyx
u1Ow0yppD+a1aSB5eyYM33zs7W3S5PUFVLXhS5WGofyYbxr9jymjmZoOyEMeoYp9
cSP8XgJHvPbvqwC6MFh6SPoJpkBpg3AzxLAbDRjM1at13qlt/hE1mTHdJlBMdN/i
3Mv0nJYVELfsF6Qkq3ThjTZwvh5t7oI+GmvHDDusPQOhXQbiAQSQv77U9RiNOpcs
jCpYNwSppNDboTIFibamTZcpyU6hg3PDWv0aso22qxs8k7+FOX0ZiTnn34omHAxt
cQ9Jwhy3wBWuqc7nYsObBhYXFLFM7f9tsUsuRztn1zQwJ1XMcqdb7hRrdENKj09g
COGYpR+4zNjtQ5H+WHlgRnkOn5pJMkdz9tiCMvLwnn6LJ9wsNE8qn/vaW6YOaw4x
LbNxk3TKgHmOAweTgvdIe4kamNA+dxCEOXESwvjlfk4Po+bmEZNM4vSDBMj87vyq
Jli5hCyWYGjNk/m+3fFpdeYmE8dl6KTSJmTexBRYuppXE7SHS5wpufC4WeChB7xV
k0cXqxcfOHwMHQPWoClxHsrHxkho+eXBb6rO2pk8gs1n/cUwbJaLXxIC9f43aXph
khfMr0irVg39ezy8PYaj0dOjyUnjp0LJIDCR2pNZ7GCZAufNpJ9spFGeLdDDRfNE
nR7TlFq+vSNHeV3z9LZYdcYiCwGfvbjy2kdnRMW67pPMQ5CV6c8BA1fwZ0C8ReN4
c/OA/9E+DliwUlN7tGGA0+xXTryCeCvZGGPzUSmVmZmIMQy5KX8GQTFiHbYC+u03
qUQRTnh17PM6MulCQ5bpPrGcvKceB3r9KJxfx9RiVpnlxDlVW+42ly/dhjtQqlUW
6S8HmW4RwSRMow4uLRPCzfxJyR3CFsOq1XOk7TTWiBjDTHL9B9Cdy7bVCR9Xw+1q
i13N9BlMy99ipgN5DvVEI1c70FlewHjgqanjlxieagZutG1z0SNoRn9uM+TFN0ou
EgfkjZH4WHfGKE1aNmQ7NY+wYldPkxPcq9yWa3sKizAnIWU84xab/wyLTMe4kZcW
sD9BSt7OFyojlgygZuCWOwF/miOIQjDhkeBGNbVgSybwsBx3xhHAQABIfPwg27Rb
Wc/NlTFf4y+325XzBYPYOqWbDaf2vUJIure9W0pYngCLc2oOY27wnvV3BFWKiJJ1
q7e850vBpZj/gMBJjnKu3CJj5cAGV4FvXxlTtZGY0uojluZjfsuTLruX+mWhWl2/
TJooskXUomiBLOatc+bQ+vLs0pNKq4JvGkPLBJ3/kNUOQvUeiqF16mupFrtT9KQx
ynN+PJbJoNV/IJHzcy24yqfWwH0OA/wEGgtM2F4bXdYvz3tX5QKDbv18I9Ft4IGz
qID4E+4ovIuQ1DhURztGPeHevFuN6udE+vlaw+Z9iMVLBkCcHjEgtZI1L/sG378e
ndNMx9k/OOlU70KZ0mEsyhop6VPVViMQz6VIzJdxnWEGVOCeL96XHxLTn+8EZa8x
cIuUoFcPd/sdhXeV7MafulTwU4XIXTCez1OxZyMRVXC6lsCt0bQHxPGt4N3AtMeE
bxcD1Mb0tutdj/Lqadv58zqaWzCvc1MhGltzurkALlqYdF+mzCW2MsIGlO5uq+by
hIm//JKTPKaJbS4ySjmbyYfuj49T5QxYEIi8a6q1I5cTOBIzwuh82zYkjWUXCV6w
cDNfoeA6GC3jnrGG+3yCOhoNkmmZWY1ZT2yZS0Wzmrk125fM7clasJU48vWL0Qdx
5l4SBR8fnwOcGyWTi4rAA20hOhfFHHryHiP994gNGWRskgOHvtYLcSC4VWsxNgB/
z8EiZBBFNelZ3JEQgLuah7USwIGOEmIiPstFJmEAKp1svIvFNR8m57O3IW3aDCtz
Zd+lMFbTMlYKF8F2Jr503jyQmDfd/UiDRnQabYOAbNnWjp62JT5Krwr21S6otL39
6whArz1gtNlFz77/C1n86749fOpc0afP5V4cxeGienyhOBx05KHZPvIgrVydnOCn
vCpdE8myJft2Xq2ANFeFNryoN75jkfJDC+xCnN0g9k6WEmpNobRh5T41nRgMM3je
wjSIKpjRm7jfxIxG0EXtZMr5I9v2Ign9aK52lwPakndFHsU528s96LGFA0NfQxqh
c2IsaMnd14N0YlM0ieAqkLWfsjOmMMGFumaPj5AlzVwGAz35wUVqeFPe8rW/YSTH
tqIFhxtIizl8NtaGNNq6JwTapxK03WDVzsMmYvO3ZbM2D4NI/Nk3YgnPfK15fipJ
HzscFrQoU5e5M8FqIb3AzBUdwizTNxSUql4yrMTddCtrsgqeswaX+c2Q7bIPzKAc
Y97yLgOo5fZhN0WUn9R0DXFFHuHwVzmY1q4QeUIErzeiu1giZc2VJ20FpGUgS+dm
zh9zISvycAZKZlWPc8+nTLqvI6gPPLCfWF9vsxKTl/yFZJy2WyKfsdPHCu4bTB+j
zAefpIQ0aZ4RhatT0RjBmIy8nFvjE+ZjO5BMINcflLM5bZi5z4a66WkrdTI4XkiY
gnCgOk5oZN2YAfmpvPr4n0SCUb3qm6+EMt5jaYfPylQ26NYrJb2eGbt3WwVcPSR3
yffqyD90USpIvAodKHIaGI0wCEvAIIcAEAgBYhYgWGdRHwQKXa5Nm4WzBs+NLhrD
J2QtmHi/fcG7GNuGhs/kYldpJjbyH6LensOy/ykSPCau1ABQj5tzi+rD72E1o54Z
uRSvZzgQvxotl3/VjQ1TqLIoR2s8XlliTnNQBGCd+XQlDhkzh27RDCcyJgkVH0cf
iJMP3gs+M2QUJffBUUbpXajiCBOYA6pTihKNvwqlz/aRh5DcoyH8M9e3zlB+SiS9
1f3T2RhuqbWxhBOunkaKIB9//GkaNslQy6cDO7aRObKAEkTe8ojcvy5WQ/9cyfRV
+WplVLK8y5/8ZmlDuhuALc3ByaSJPyt1iQZbiTfqMvNqvMSoDqagT8DBtOOsiGaN
XLTlMJQJmDd0+BgRGm433mHCYwLjeZtGEWBMRk88YKmw9/gYjcszGfpNynW3naL3
cHXTYmhd/JclXyhZDswJantg7NPN7s9mCkbOrm8+VvGwpo/awM1yofUfFzQy1wYS
keyh/r/jYRJz2mcOHuZOmi58i6NKfrlO8gIuamoGARMYWE71Bg4J+yGdmvbv62XJ
NL79pcAUIBL5NGAgHp2nS4DilnCCwVsUxIWb0MQKhtcfoNd/hApL9BOI4eSb9DWy
sHoEmHsrLW5oN4ggYKF7QsLwbcKj8wL4T8tCD3sq1flEagJ1zGudqzhw6dmVeucv
XaLNf2RZtt6o8Sa3j+EqSBc9j7Rkj4JLtaGRg+ectbyrxfnr/+fpnVjopa6MXn7a
UkG7V0rlyCQxy0xNtOooVQH/ZADb1LXONoPqYIxeh7bleH5DzOQ3r9NmSlPkVW7N
L6iLEAc2TV/q4EJqnK4mjdioarHe30K+x4TptiVjq0WktVUjFuP6aMk3B4p0nyGQ
SEt1tYRvmzjUwu9cZVMGrlv7lUMo2mCk6zDef7UJtIBP8DoQrh+6Ohon/u2B1xg/
gP5I0c1swBKuT0lxPw+iGMky8rTkaSM8sXqlh8di18vlfSt439m6uiREPwKUbhVi
lU/uplmNeau4I3luu2WLa2FQfCChugfetJao+aYtdIUsnIzvju1sqcmQ7l/MbuMi
bj7HFxqwKNN7fRcw3ASOvL6lNi3rdV/kxryzxy/YSq/ubC1FoEtalE/51JrPTNoF
8qwhJ8ea2IxoaGk9EHIhMKQJdqnJe4ZN5kUX5L2g1jV6zz9799F/sQyy138relLx
x48osPm1NdjzAYxViBLdFNp1YOMBW8/TumFkX2VlLTxD/Sw4bwlU0Wg8IEidQ8Nh
LDyXD3+TsFQhue4i/k2GfPM05HFTvtFhwF1TR/eUpiiC5JCRthhYvkmBIW5HIJ50
dIWFSVl0/NFdjkbtZqun6RNC/aw4ZCKWcmT37VuKm0Nm+m45++t106UF3iThluM6
Wwn5FyD6Xc8EdTJwUQZO+yPsApJYyNxMEQrX6Qcoado8EGCoG/s+M+hjX68sKjHa
L5ty8C/ytqKZdtYPlty4tujF2S0OPaDTweRloRiqaSnUn2vsKZAFnuuYo/TIjwKj
knpXVxoTqpsgWIU98H+fW1kwl2XepqREVGzn0lsA3WuDEvXOT56mTVmdvZhThE5K
RLVi3LrYmLOS/3OZoIhcIu26u6qg7ZnGVYHf6wF3UlfBOU7zmThKg4n15AUWa7yz
SDV11dMO3jFFdnnDCpqba76305FHWo8s+wf0xe/uwfKYxZy17F5rfNlPKkAGOhU1
J3azLy+sEAqZgGLq+MtGir5ohpBlhm1jn2AQDL1kwglcbwYkFwB8rf9B6YDYvZGW
2VFp40Pl2pWWFqhKIsPwIuUJoLvKTu+qJpoHt8xnD77GDFjvDfVc15b0s+lzhQac
abXQVmNgibD/FAADXX8rPTQF1WIMVm58qOkpq34PPBQfZwKWUPvnF5JehZEFx0pu
tVhZ+stUGGBdXTqJ2BAoHi6in13nHJF01k1liUw45kOG7+7v+ineQk4wmikOqqw0
pSjd1dS5CvPRgqM2eh72py7Jo9ShwTz0RYqFGHloZ144hl8bC64i6n2U4jZuhM1R
RAIkx+UsrHObGkpox/txl/EAxk/5RoMaPzEALfc4dGa8wlCKZITICXaVXya2Q3Dk
84QCZRfBWP027hp0N1llB5SJE54Edn7fI/q5rQ8NlfQn53O2PG4YQctwpdMvsIaE
bkyVvaqK+QxzTonM2QthLDx5jL+4NgTBFJHfbCI5fKQzni6ZwK84SwnrIQm/H429
3CI/XaP+GvRw+f9Erbh6dGc2uZ/AU3CPUpzbJEDjB77jmAXugmiruIRbEWkYiGHg
AMPaeAREPRKHk5O08qt6/otg45CJRKtj/FBrIOgGjzewglJ2vREr4orGmgKIe0Lt
/iUvqXQghtU09jilCE7iEUDB4/xsykPw6QHCT+ojMNROjNQUvdshlkfqbZEYh0vP
lfWs+mW9GiXsadQzk1Xodfg1rwvZ01lpR9+GhCRFfpdldKyJ9ph0TH4Yvpae7QDg
21KraRhKj25xHSZF1U59SqEoYdb/10dCKMllPGl1ScZElp0LWPjjJrhrEoH7QZu0
9tNHVZ908LrDBu6PNKa+K4hwhxYluK2S5PqoqGDYrKqmE2K+/Ekccpw4ek/lHs2X
Q4Zun6sSOuDNiOaBF+hYXy1FHHf6b47hd9ZbO2I1YnOdhiaTO4lBQFUSqKiYl6Gc
1wmBoGfYBUFC80a2s0bBds5I7ErCEMQnuxbVRfiKB8vmY5S9Qi9tb02aJjuGcLOd
jsxQCoRk5a0tw2jECFUVt+qS/hOB2zYJRc7l2/0mQ1L2SUgd2TUperF8TeaIIFZa
GhNCC0q+496+DZc6CyIbAGryPwPcL85o9RIr5hM8uiRb6uaFIlvwmsrULpSh3tgx
T+E366jFdo01WZhM+gShbV5vv5PRnhXdAoRa1Z97h+G4238vEIF7dnFo8g+8NCr4
Vzbq4cBZTBlCB8vHqLZBBsiNZq5l6Gc+x2NMbykL4na6ZcLcI0+I6eVxdAgeOCHM
T97dCIWcrv0xnxTDOcJPlZRX7ZvtjMneuvlBHbFL/trmOH00q+ND3WACvWBT6Xj9
G/Qz7DW3rvUGYBlxoyaXtfXiYqemo+fUEvmiplldZ0pKYhE40FLTHHf7dJsX9AxF
t4iiLHR2XyhMwaArJeRFwoRDUvJzU11JdIQ4gzZroMPdrdfK5EDgTX/J8kCgoHVj
OFp4nnP2ZjO02u72NfVWlcUZaNV1+psRusBB5IECd6ieBMlpR58e4jmmUYJOphcp
sxJEkf/bJx5O20sLqeo6MUS8t4K4O59X9CF9n7BhA9M/UNvU2NIB3q0cvx+df6nl
//9KSTLr2J97PAnP/LdYE6O+AA59fRpfGfQMfnhNGsiLrAv7D0pYl75FfuFyqNPG
6tu3jVwEHjZG1aE+3btAkV6GufeKAHrckkL5fdI5FECjsc3uEa8IXOBxoq61fdRI
oqOI8kYNKBw6BWfKDMmAQFUyvtg9nxvSKem5C1qLWayncTztD4zzQqyi2Mhh0H5q
OpXp+YwGoq9KtzM+Aupzk8JW/MHx3dkoTOErt2Cr3bbJhykNQXTQgmZ53kXZ9nDg
oo+ABabBrczioW1dgUF4Q4VTO6L6GhKj9vAUcCTKlIQBXEtQ4qZEwKVO40GM/VJ9
Unja/DZ7fmoYVV8NPkcRP4YqngOjrnXLXc8dkBOUhJAyq+nsrs8Fsch/Ukjk85Sf
s68krq7gE/P/HjjL+wTlKkCzKhCi4jKRlDFX8AaZlKlnOfkE43VmuKtWTqVgN/Zg
oihsf31N6F66JttnahjAmTOvUF9QXlflSsLzrIASH3M4LBUiowOa8iAwoTkPxTIH
aIuzE7HOtvx/o6jH63OALn9sQZE3R2SCkPUoMseaJS2BPBiB+TySJyIpyJa7Pckj
2+rFwIdMFUWQhfIgcoypQmgTZPHbofz9ifc0zsVB0aL5Bmi4Zw1lVWd6WuNH9Eoh
uGLXcQ2oIkwHByoKk47qNQqR+zr+1FfyhpV+RdXISO91TIJRi4TxITjtjgczokAJ
8M/x8KCb79H71nPdxenLHoiYxrPxNEsuBn7NzYFrFFYNsNjxnsi5jbLVBFBWCFPG
oJfAElXASOqBFVjbe05Eso1hb31gh1QBTWwAjqlJbBVd6C6dRcbyhjAPmfXshTc1
WKhy3vhZtzeeZ5YIo55AH0ZjF/2y03gHpfmaYP3N0rRRaQ8ZhiOUhmgfYSd1T0MI
L2yZ7SI4/VI+dOxVAdMhFpow5Htc/ytrDoQRdZFpv7sBvXQRU4pknUVcBUoFYclm
cpGHM6bstyXpAOW+2IZYEccceF9Dl6LFHX/hL9FpzeCQ1dtFqnZPV7TjZQ+SoGQy
77+Mm8ImUhLU9/kw/HX0ljJaPGhwCtwPVX8W2YyZWRsNKmevHRw6IpVp24du3/FE
fAHarohByJmpa+9HCfrhXDhg1OfCV6UpoQqoRen8JQtoRfY9oMPQtzrbTteJ+CRk
iQITkuytXpMMm7Gu6wdTh9Mlz2GjetNxckCGC3rnYVZ/leENGx3tFIchXIhyoKsu
glt4ZxPSnspYPmsd+KmAT5nwBG8Jr6O6djW41MqwA6eekpWRRw+J8ZXhQR8xX69V
Y6yIyhdrNNTRCu/2ZiOdL391ghfOinLqsptnBvGmZO2GRuu8Ekz4lUnetRimuhQq
QFFpKmgFfid2sm7VyhhldycZbiCN+y8CfGF2HnudTxNwE5smTEMe93AbOLDBNmXY
ra7920MUTB3gb28O7m2a9qNcCKqMisjLhqNGNae+CfpG7gAK4f6E+/d9NPLI1+o8
Dig8txRD8jOOk1cXxqTYcUHFkJS+XRk9hRnRSbX5EHQFXUvcd3DZf7y9syWeBXcA
JrYhqhqzNLfUQQP6PSxfQg3eNF//RfSmVazy3Ip1YPmUeAxCYYEM4wacEVco8VgG
jfP0WPNXdfRnZbJJ19V4Q0OBrWwFQxSC2j4ru9S641IZNpyvnF/vDEvQGz1h2hsy
D0C1KkdMuxssrCFhfMQcqdANc9h5qwh0wdG0iIbCAA23FTp4v9yNCkmxV9bQXe5G
R0NmyipMnwcI7ZEYJD17aRiDBXcNpkYcXQJ1BlRIYPnzIK8PNbmyvLFLwSrkKbeE
zAa6+nYOdxOr4g1GLduQ0jq/T5BybOvWV/IBVeqxFfW4CsYEqfYmS4t4TxWnsY+f
lO94MzTEzQ0SyR1/Vihy6DBJRfPLi5CMe8blEmQVe0XRxtVmGaGBclqQfMnPV/Ua
t40CQlsAoanR3+yq8c49bnVymy5vHXqh3UCmhtskQix5xI6HiTYENR18Fd/Fq5Cq
WHznf/isy3w29XU/+I3mxj4kCb3c8p/l3Kldu06KuPneM83sdJO8r7ZUfQLb2yYk
K2ILsPoIJWSB7wmpj5jzQYIOKrO+Ku4+JCP9J6HQ7ZwMNJb7Oh/wlqC3JKb8Lsj6
3jABMO6gGzbmFZX6jab7yqD15Qr/fldHKS3sPf71IckpeIuCAp5q9x6U03pOgZiZ
tHAODURRa3FEKW/SPQHPaXu3giR07c0V4iO5cRY0jFB763JvHMLnFMYtxgOoLhHV
zVYZYcAxJPCakV9wFpJdVG8jRyW8QylSOwJJ/brs9+2nJm7+1Kq5Q1NccyqTX9Ku
mhc+/UyfbDEEKLuPbCWwhYS499gWasoSbBIRWCSbbfmMBme6EM8qh+6lnLLCfZ2x
g7bPlYIIyb2tqJYYz701NE3q2ZJ3YbbF2Y7pd6uTnn3KUBYlp9EqtCa1cSR6wsmm
7MEz85mSAYJQ1IYeL/WhtiL4qxEcFMPBQfBSNKocjQb9myuBVrUKn+NHJkkGnCDl
RGbyBKkYqYcGDij/FtoM+f7dPf/McQ9b8DadIo1FvbbTnBsA+QzSRIkdDWuouFUM
cHPv0egoVpK84apAii80I2uNbsaRkNEXUSDrij1S2koq87uRKGr7reLtWcfZ8Bte
fLFZTlkumSflcU23JzDiMuisONmmE5HTe7J4dkcWB9ymKsRLKWZ+Y4VujTJkiP2a
1YUpv90oLFH5maXcnJpiKePvvsrM6fWXdOwpAA5TthkwXGWwsifIq56u1d6ExPbB
5CVGUX0JbuNHWDJyREGAIRQwUNg8LmytOtfz6ud9r0ZXNDiM+gdIbmuRpxt2/h+R
U1NJIRc3MOv4FsP+EbGE8g93Vq9qK+VbZGIA281PhVZkc/M6mvowBolbcXBM7IKN
GkFTrqPJlW2VexvPMj61u0WaQ3qVR4+9WWK8+XzinlAzbfrjErtGgJOBCDQq3R/A
mBwG2Xg+OAT2wpuD46J4IpjYam4P1nZwXttwUN3c6C8jfjArn2Quw2ogLmgeYGXS
d90AmObXW+XE9FDcPDS9W49bpUSng38A8/x3lSAm3JjtCWCmjELoieGxHUR7C0vH
vFeiDpE4dkx1kkZH9ViTBWzT9W9e4tZipuYvFPiBtaph8eRcQI16z3VdF4v8/oCe
VgWgzekdrIOXKT7OzhTcx1ci45Je11iBUZeI+NpaE8QN3BVFYN/Ff/CU4Y1QzwpH
rXkBTKsYg6+vo1g1LXq7r9Xim9sLOW2v5GdAsvW3vfyy+5BIgoaPeIpb+Jdjlniq
qWuP3YwHsO/gb71npPrekcbzuaQZx3zn13qFr3DxPh6ysTVJ2sdsaizMymUm8/ZE
pDEcvprU3IRR2HgpwCpyQQ/ElDNw8QFLxUqWCkGL4GBHFwqdojUiC5RyFeprr6Jp
ELIGy7hzjcl5RbBNdQi577JFlOiItfyNa1S4G+wuzbKMw08Ao6yTva/C6XLdHUFN
7iKu3Emv7KeN4bH1avE9nL8kB+sx9EnQRxLhNbJ8J8z8h8tHOmmkFLGSz+rwsIiX
frDT1UA4ufc8TDs5lYUpYL0y+Ev2m+zkwaD27viDUePbr5Fgr8tBHH3NejrwFb3L
MAqclQraKz5AlR1VbrzIFxMFBw7FT+b9yaidcOIKaDJqfNYuwYeyzGECWjkPddYU
J8vTQh2DXMV8PpLJrg1KJRlCL76mSpvpJpeMO0J3yj4PUhW5HkmG8SD0OnaiWV8p
16A2LlAekUZjCksroxBPJvzf7D28p2iHdhKRA7Fn3Kud77wvnUDbedq1oTZ4RAZB
bTH0h4e4KmmSQzE3rZYMnNSOxUxZsHhl6q7i19hBvt7wHnOBByj9RpjajGKBKGOb
G2iRPjYZeAKFXXNCirZQzWa+F8bWCY+6l8kWKqBYdldgJ2USzMPKvoK6VN8W2Yox
FzYAFHVvdDGUt4XrRcjIUPTvTdPnE2yxZ2xTNoUy60mfo8iKv75SIKNSsj04va0/
yfY7Sf3nvrPy62iwuhsnw4YFG+eYeQPYlc41yL7TehZwCGuJThvANrRic2YzuSq6
ouBed+UiYVgQgXw5ntN5Lk4eeCl8in70PBGxVqYwE0v+gOYp+qnOcKky8VHtwNhp
4xqLhmzMY9tyOQqRaMuImmM+di2vGLJjeKqV8dyNjSPwCWjZi3Qdpy9st8SJK47J
8DL+krKyigoXnZ78FcW8ag1U09too+jQGbOSt6rW+RoQZBhrm8iuFFbp7MZb0jHs
7IaHAkEI2C/LDfS5Q6Q+MjXTis5LneA0Pe47x2zLITUM+mO74NhZP6vZU6cADBJz
YncjS8nTgf+iCwBYYJTHuwR1JqhUnPV4mGVtyiqHj7YUw6uJ2h+W94psrrJF/i9w
uL4RIrCyd4rZfsRVbtYctCPBcGPxOW6SJjuNQ+eq4viCpD/+lWbegnRIF8Dl7WtJ
84eCMVaXOESkZGYpXepHnJ68DWZ92zGLaCHhBc8DT9cQr957NlKCSnVdPqkEGDLk
F+VOGxtq6UU7nnbDHfq9sxRiKutgAf88dlno0lv3dXF7NssLPhCE67IToDvFv5O3
ajmrEwoPRTkX624B8HKAglx772M0TSsaxDLTuzcRqm86sAsaQJOqJ5t2YPdrVda/
Uj/M9jAmL6dBbb4/d/h811IAzbcRzhBusC4GByVzRCUaLjwogB1A00nykb7OewBQ
t2jh/OsqzPOwPdM+Vilj01yNCnx5m3d0xr+jj0r7SsdCDe2Es6yRRMQ5TEP6R0U2
zEOazUY0KMG1I5qUpDu5eaV1+phqFV7Cw1C4URTKWxpW07Yw5w6NHZOqeDn3J1G4
qucYTHvhHdMGsZ17GPWJKp+Xgbqg1XxtN/XOIdKrdjEBd0MwT0GJQStqzu+Q3isG
0TXFgVhNlPltbh87FEp3eopLugqtaQFIvB6qHQ9BJi9AWc9pVWbfPBkwaTaLvfsj
2OVW/htmOBx3VZbfXVO0ztjUZtqnXWwcipWg2zpmLAeHE/j+2thNzFd1rdWUTO5C
0LJJgGA5CVJJhdiy936b2Kg3q3PGbe3D8aQuriKJW2+ZFxpbdKF5aFnZOkk2FA3V
P9N1JhNHGR0FE0CQnHB02DmTxB8dFkBaTmuDDZtbzC0STclmMOiHP94bcVRfXn2E
6DNQ8WthpjijDm9+6zpr9Jt3933P1Lwtg2m5XcJFlK1vXh2GfQvwztag8aTcQRWX
hxg9s9UGKd3ce8nQZIvS4sfwwfvIqtaAh+49h/2u5kqcRIxJpKQ3HH87d/tfRp5/
Pg2PLQ5CioEDtK/QDrDKIUhVjVXn16RJ9eY+hyz+oyPFDSUWi2BkV6+xYADVjOKz
irJleRugXi/0Cdy8o7/sKpc5Ma3IoLQnENghwyvWKFsPFth1An8qratDevVJaTmC
9F0rrCpEO+ghEmNumdndYaAszOy4tCZb7FRJKG82+daOHhkc69p4X7ls5UBVAi71
f2U2Aj2cQ+CjPCRn/NqOiTi7EHKo9K4ttDMSKdx+xniMPTKdn7m3LmA+4SLhIrRb
7wSJT7MYrOnR9+IhuNIgSKDRV6F7xnJFM962tsNlNKhN4W6OphN+uIknLQjMmMC+
fQCC7hoZrRnw++NDFnBgrx0m1EeyA2Izqu9VBjGfWGSBJX4klvkv7nbS6wfUTnMN
iCX61bEd9rBq1TYWpuct5jeD0AXs+xQGKio6g0P68cubh9KThgtCQh6rzh3z/iaD
zhb0acZwiwk4nvBk3DG7HrUaSSXy6XqrsX2gFCHz3MenkOiftvleUFtMt2iD74YJ
EdBX4Ma+q2fv6ZsTb+nfjbdlni8M8tHVoaJA3Caexzcsf5ct5UoCs3Cx3b5tFXTw
WcRzqGYBqUp4hVHR6ofD8oFzd4KZTQjsZoV7doA0fdRKzBQtrXDophC/u5JEmMmB
RkAO/0C4/6XCNhJHj8YZXun4glWjZmOIRRSQhUy9aGj2CDY7oHKyhJYP9bGgYH25
W4xcv2svRjQVuxKDAogm72dbN1zn7yy1uSBXEjLYGagtuJlZG6T+tmrMo6EXESwn
le5qXxX2wUEqbmbkL2cJ2ezFhCTNOb4ON08vywpjgVJo1RLDAmmA9pGWrl6bbaPk
qm2fjZFQ9K+Lwkgq8YocJqhtuYdBrMxYyL/b3upsUQ6E0juuu9HMB2Fcz9K23Jvk
I9tYvtErS+hAixeOgZi0LYMbtAIUIC2/0Mztr7TYEHFFIHtD9SbR8HGLYl9CL7mn
/pIavMnl18gyBh87JEbhBJEUSgFAJrBRz2S6K4FrB25sUUt66yZekp7a/aaEgFGB
21psv4RuYXPYTsP9FOP/C34nqJBrkrP4+LF3HJH6e63AzUwrWP9WJIhgkDMlLsEk
KDaTjOtGxMp8M9PWasu3HKRNNcXfLL4CN23C7rhUxiSRIVfNo6oY4dVCAbG+BJf1
I377mkkVxPHDVxcULuxQUiUd7kADUt5iJDJSaTZDaje9DKODUnoGUCHqYhur6S2H
D7UmQMtIRA2jD+W6UKYw4/Cb+mpAYMOeRxoZjxcDGWN2XHyezzIY7Xf0Bk7kXrfs
cEHyIOR3CXmUEItQt+Oe4AA7+qyMlbCQazBDdT0397J549pgunGAB/Wdg2ICTmHZ
qHRqIeELMic1fay3Zr9CUzCGMDyaVYPiSJoL2yW5LZnj5+83RKz0m99sBQReRfQi
H5CrXEmnqwgXLUKE4BotCojt2WRQtVPzAM7WKshMY5PFXq4DCHfdQbT6+PIy/jkC
TqKO1f/CdYhCh+mba6KYTAd08NNyCcMhbUslyKKKOMSe5ZECIYqr6f6wEB07afdL
V/CaxusNlyjtrXF51OY+mlWuCsO88P3srpezcYpjWlVFlljm3Ez2l88FC9QNRqpb
/Ga+mjJBT6fwdzvlTV81xcjW4hAhzeBiDB0CXNT5snBzUopw8LkSU+y5Wh+N7QHi
4NJYwuUE1ycuv6C/iNVkE7rreBXw/aEKhA4XHG1kJS0Iq+MgLzLoDc0I+4Bpg+QA
YF5pheWZWn+5vD4zaqADn1x1u+2AObEpqv8tYGb+4gUSaQORd40GV5NQ9Z8IDaDK
fHRmUezVhBMk3iSygWikSokpF/8mTqd7fdWg1j9NCC975BQB2wnxA2Yh4WyU/ZeH
3JU37s7QoMoAHyIMBtjhviMI5TUwBi1+WJEtg9QcxlN9nhp9jJ1Aw6p+amGlbmDh
CpsXb3rnkQ2kJopEzgtYXVGCFFqAuWoUhbLAIWKBKE9kQgC0+oqOavqMZu6kSdfB
53Y3uQzczL8Fgoru+mafZXnW9G5TQMBqmpc5mZXal/sGoRcP4tWagJKYkWnJ/Sk7
oZMT35+8ogOeWTW6tc5UdmeDnHBkOi51/avSf2SieTrdXxNQTc1bj1eAly1dwyMw
K5m0qH/jw6POjVP7mdIRhh05b9Z5cb+KIt5ujHURawfqmtbP8qzk1hr+wmNBWlce
saSQhWEqPlwazTd+NkvyMXTyje52aCB4XkVYqkndbq2F8CmtvLKf40bnRgupnKJr
zRIVXFrblo+cdQo42H0prfNbNBTod806OywiBGDlTiXdAl6M0ucni/uZ5jnAfAe6
n0pWkXXtqApgXIzpGxYpD3jnJoee0a41YExbe6fazBraG5FojUmI7NCEL3eGFMLj
uI2TvZRa+XPLGtV/K/+9l0Huo94iw7JNQ3wblBDrN33rnzc+neLAniF/RFCLPGjU
Y6n4uQGhqXuRkaIWv7vukRBis7wdJVoi7aIFM2hntnOIFumlocmfCR0Jg8vsGjds
T4a7+Kn3knA3Rv4hVx+Aqo0O3dmeAktdczEcfi17V3MIP7olegEH/RKS0uMzZgH7
vqlsik/najhAh9GVZDdaA3y6KEeqJGdG4xeY4P/DWGA6CmIXzqxshZ00kMgJVG1V
tp7kH+Q9UFFJ8XOlr1unXnKp0FqSiOckunfM2H9REhbQbIIDgYdXEM9s7fCgCP7O
PSTGIWOOuOzU5Qx7v2Tbwd+W95CBtWT/BH7j4vkmAM04Ug7Ps2VB81CpqBntO/qi
Tn0vWenQH1Zy4nIZspvZZMuDDoAHPT1v8W7yxRue3d0+5m5NMgfEHZlY3OMtP10B
gQ+SU+vkftizjhJrS0NjkGQ6X78Qrf80TxW6CDgQFk9cRr9/XMzqfdwNpl1+DtBr
AkM2M+CbpHyHjkg9gte6/59RoyXV9vRPq70pR0te1WvB1r3C8uJb81NF9g5xW5zr
dBmkQqCZVs73By7MfD4ycXaE3dhzxKpJXBSzXNoI5xs4CCzSQMry61VxxhhBIjO9
PB5MIQ1rhnB7HJadvCaYScAW7Te+LGfkZ1kO44xpH3hOmHocDSg0OHCNPt7xlDEN
+WH3OiOIae4OnCdvG9MQEOUtlqidKVDUeDQoFl2x/IBjN1b1PQAaJrshD6y6pL2v
WFJxn406tUOhzicu0eh3hPvDoBTM7Fde/pkvk86VXEz2CMQMG/JE1ZI0LyAmLUrM
1kVj7oGHOUfuwT0yfKTxGX7WxuvvMKoGiR4bVxH8Ls9axHW/mEVLxul+TWbWijUl
oiisvbxU1rzrR/kbufHIdQlWIol9anJwO5wHl8stpgKboC4xeBfjl625QIyumT0K
WiwmAR+qUtegYVAKbu5ZNHrpXvXyi8ufnWXhLDTTmvyN7vPmhP/jHaq0vIaGJs76
0JH5bTGdfTHirKzGwl/BJRrnvERQ7C/P56UFSliAd7uEPKnOc11PHyRI0ftKkGTp
2qJdhMkUhyYCKnxPBC6zBZUQmGeVSr+wgB3RdJE0rscuMLl5zsTitViM79sw86AR
NsxAtf/HEcUaspoeHaD3g1UgeXNti63aJgtb1AY/v8w78yygiNL5MkyO09//R96M
wFof38xrIwiCgG7aKBD079DTjLcI2RFoiJGVf8zq98X3En9cBRoNXFVv9i2EINJB
xXlZdG4hrnDZbLPgZxD5LuXzTR8w8tbkkAn9J6VUuOLv8/i0faiRByHbPE236c0E
Wt/omJmAPkdxyDlu3X9eM7tK3kCLX2aqwUY1unwMLjd6zm7naD6S1clhRCMbifVR
SeWIoBwCY9MtvXxYx8yMvo1RwSg4XrPBVh5Lzes1A19Cy+BPs2msAUf5dtdpNy3u
gJno3HU0/F0ud4J9lSVYIFFD2P3BiOmcU9M8rNk3cH9SRrCJnLudqqxnQ8jLSKP1
2ONPloPCxaQFHypVvRyaj2eXABOux2G4WqDlwopsDMUEgmqx9Rs9bC93DnpAQboy
Gt4ewnoKTkxocjrKuAvpvnkUgOecCRqY1ueJNosU8kkxBNFN6Yn2QyuBaEAZU4mz
1lqGvuHOy6uzhXu6r22TVHyMbtrlZii9KxTg7G2moTn8Jg2pIOaA+QUKwgeqQd6I
jdsCAYXCPQGKH0PKmvEdPats/1mj+4zYas4eoUdhTAWASMJRsWT/ohy78c34APta
uZkW8KACr1vyM3p1dUm6DdiUBKQWPf8OasHawExYH3A0pg6pEY/Ti7OfJUJlQYlc
uCw6hlXZ29RSCQjGWaSbiHbKwXJVsYCVW72n7Yton2DEp7y4pMI1oTodcWbkdekx
aUF3jJ5Jiuf+yFOEvd2OjOJ1N1q1Bd95/lYIfUxnnj8/iJoHLCIpSyWnSbMxbuLw
5SalAYy8xSoalAiLupeKdf5zNSROgJxWAiaZqH7NpC60C54EkA3a7OU3R0wiqTiv
4a1BmRkiFz8WH8huLW4EEqjP4QVw/3i0+jYjSkxXtSFmLQtOnIvfEbmn1DOjXNVQ
FJRrMKumFTc3kclnqr/SsNxKhcKM0DkyWPGI0R+sy1W0JrCQ68UKR1SNe4J0sOTM
hbr5ND26UwPgKisx3Dfxys0u4LPEZtxLPuR3SuUHxK/WsDvw11HbgDp1lzbdWn+l
9XEWhfaLNR62vDVUioi0+07oSTb6q02yw4UmAAyVUyPc2E9rSh1zc8+Kfe8BObAU
FYF7lFFjddpZ4N/pXSaOS9/qC9+vGCBezswbKq2ogtV0YPq5jrO4fAYmhhPCv25L
bx7SHcw2qnc9nuMEyRCpqEt0ihuIhifx7pzXA32/xjdjQoOUR8at8Z93z96mUBZJ
Gk7pEG9XTTG1tSnBjrCP0lHGq97FhEVW3xeKISUga83gcTXM8uDWNzDBudj5XxL3
D61xEw8vEu2UB8AwgtDxqiDinfQ6H8P80Hcg2/wKx7nmOQDLJbSmqwDgZuujbVJ7
zY0yEAQ1YR0Bv+UtJZLUIxWejh+yTY33hR4OUF8kCQE6h4lp9PH4Gfklmd6T8Uud
ka05fdYSIpC0kib7TezZ5IaM8Apvv9me4kTZXzULxbQsgfVh05kG2ZZTuNYHMwhG
Aq9Hd6gQWfl5TSznLaeDgJGDic8QR35vLfyCZ0dGg2mjteHcFMlJAqwRyg4PseTS
GlCWwKdUgoVo6Rp37FUNLrBQW9OAhdv0UvfaZBz2+Tra6g9JCG7UUrYNOqy5XMNX
NOXxxKkmam5kP5aO9P3sfFcB9m49kaQDS73wxjMxipSYJKgN2yCgefcNKb1lZkIS
C4tNffhf0yjhkz5Ax9Y5I5abUhWJ5glejwRuEw2c5BE+bhUD0Gwk4+jrbNGBjc3S
FWptI9c+lfpfMsh9yH9sR1FTmJKwFogAp+wkHJNs3vm96mW1bE233o+OAOQoKG+2
rNdr6F8mymY+3BcfBGBtavnfIY3yBiniMcN1G8/kMIzzLzoc2XYuepmHa2FO8sXg
MvVIHo4nK2Bg7jeaYnsN5tvQprKyghPYtYqmYLiATKmDAHbKnbKZzvbRfm8C+Joh
v+iTeXkVe6RBw7+8EfogBdcRs9rsm/ix/TOt2GXFNvt8r2o0cWF+Hp1+k7WukJ39
Nc0rZwzMZhUYWyMtS6Vbkmtbl5h7f1ud/MMwRSOEnMu9+8X7D6E8K7OszCtOMgeu
MqkecneISeuUthvEAglJepraQltPSi/ufob+DgrSPz3LRDsD8YxpibXossM+mUdj
IuceIpo8qI2B/vuG6MD4xoe+YntIexDlBaX2BLYqOlOtdxBh0Di+5AXDiHyRtzry
8KRKbz4hRWJ6cftLJNlo9Ns3tkrEu7ggfQ85aonkzVZG7Wa+ZVCBj2Uq07i+fC/6
0l41yVnbgQckN7moJ7hIWMsvvft6HBaBujzYoqHu15oiiQhmhZHIzKhbD0TJh2PO
CqjpF13GJuy0f0IsrDLdGTzlaXuWKNWdYEf/6kPZPDvsqsxkxLUlXZCcaTuIAk4e
g5wlPf1pQ0wt0MWEiHBYpBmW4e2EIXGNQGGxh/5Ajb0ZabLtiwe1ne1yKKwYBOme
rMudXkbC3uy+FBhw5epeDwHVe6PMuGiBg5x8uuQj9OeBfpUXZi8Di02FrdstRBCw
4PgP3FCGnVwgqB1KL78jVjD2+nI81zGth0+WVMl1c3FcCeocU+8g8Nd3ad20dloI
KFsqAHV2ZAPAE/UFn6tFd4Tc+3FNCOZCFk3nVxj4hdSf81gg7a5+9jstFEkkkBu3
926yXPCqrRd4XOQEtp+asO2uu1+0VakPJUrCw/rMRLBlmPW/8nNBUVE36eSEwpq9
8vIpAz6DYs6pNtGOdKwpXz31/8YDTiPHpg6yA1mQYoQetkuX3vISN24I2DOWwvL1
rlY5ZWLjeNovN109VmC9Pwt0qxuQyXY1LZZ07fxAKd9T/k9zi5koR3Wym0t21ckQ
zpXhPS7Leqzljka+gSmDlxlqpFdBlKWnnMMhE2CSGOo4XZ05T0uW63Lkdws+ugT0
gXHzLKpZ0LeS0a7Qz6IEyr55o/va1mzF+CQ1CI6WPvm7Xi/XxDVcriCopDVmFDOU
6DfEf2CY1whlGJr8L3FBrpYxLunnplUB9OjctQekaGf41GKdgYwRPYPMly4A/M22
yPULT7EDb+91W0pEXmdmq2biVKoHyOqal7XvgdUs4/vatrSBSciZ4meQdpxCfNM3
IIPXKGK2ZZdvQQjLZMVO4r5G3+SjsXsNGTu/evNYPd4Nj4PjRebnpvf6kdy4vy2o
qWZI/i5+SShcoiYP2EbK8WWAWxHmjyQuFG2ZiFQ0ZGCI0esAlLJkCD+UrywfAHiO
/d0aUYBAhqgpqiX4MBxVEDmIWDPguqL1H55dMvOHk6AXwHURX91wVl/DKt0/4DhL
sIbuQNWDwJwIVhdTmj809JisPMoLISUHLiGB8okSF5+3RiT474fH1j6yrbJGt5T1
5g3riKJ8qwJl1dY7+HsVZt6wHdjcELaNDNMh89y5yykUIRw9UZ4f8zjaNe196c8U
Zb2HVZ1X3Q+Hrkxqq8OR9zlUSwZSGb0qOiBXWfFIXyXYzO0qyNCu5wx4rXeBv1Ic
A1cGnqBUCEPC9C/MkHkiwq3hwneT9OvoPr6KRLqk/UdM1jaGo5PmSNCUpYfQ5kCT
keKjM1Iv51NqxTd9T4G5odphaWb+qJprUWTm4clMN5OrWeMF7f5SDDBcuX3MfH2x
STVTQsVTI65uNMDBCtr/5yiGW+CvUfmCZmx/zgauM0N5MBB9WsONYmJ74WEqpcYo
AIR/vIcTwL5D9TiW4sN/DK3je/zkUCzifarvpvk+34G/VbO1YUonWThvUA1zJgPg
5TCaZApLIbjMQ73LfDvPZpa8dcumcc1DZgIvZ1/LZ2I29Uvb4kdcrAlCbLgy6VrV
/h2oqr5w5VeQgMzrplWHNrpyltPFTWDLXeFQ6e+On+xZrtj8NA8LywPwEn0CToNz
tAPURmt+il48Z4ftmipdgYk06Xr30r9kWV9UNHEiStStdCH1cB+UkGT9GNvxyoTr
2Gk6lmD1pKd2eV7snen6S1ZyDZEyG8OQMPB/NQu9XmjLDcBi2fXALS5ovQx8MO8T
l8W5jCOgEnP/HXgp5ampbDODdGpdAZqWy1VOLNqfo7tdAtVOjzYq/U2PB/47YY0Y
TBMpYMCRmKAiIgZEhKPtGKBTRjdG9ef3vuwtdXuRrVkhWq0nLruRqUDPYSOfc8Aq
CGmqqGgCCwVXu0GtLG80oE3a74/y2WtEBcYXthB6L7phqXq+OnAxPVzp9DwpNfET
d6jfTb003sZ7dUaxhNPNWSO3o4hJuBcUAgQxyzLlA8e5ck5mlCTm+N6xCzC3lQJT
G4EiosDW9PPoIwB5LeaaGeY2z/regGuPoLSFnQ+WM/H7QNElfMgBLpvHlkPDyqOv
V3kbVPUjc8zxVTvjtrhIofN1VnWfsnyT8+PGsQtj6ogakW5NLF11vB4t5o/R3KY8
zigichwlxrnlnvwBXbXDjDXKiTc/nPfOQl2xyhefhwLCDOyb+m7TFCRxKWSJSi87
mxpYsWdrSWePD0DO1ccF0lcW51eocjLUZTnHp0b9jXXR7tYu1KTNaGXtKEHG9OC8
2k08CsUAEU/juhO3DJKtswCubj7/W5M4vmMiHoBZ1mJoihv3Nq+RbVpwSzkhPSLO
qVegeX0/OQv785VetVhJ57ioQA4QME3loBW7iSpRJXXjAp8II8wiV+REvRKDGHXt
GEyIbjACY9YX682p9gQ6/HnTb5a0cnB5uTctC6/VMVhnw87Wp3CmCeSL5lbejiyZ
JRvLL4wnOzKgjWet+GTE+nfKGeX8vGrdDpGuZp8r0sTDCDzP1kv/izTcCZuh6kMG
lPgWfs2eNyaOUQUMTncp66Tehdqa9Tl8rROS98/VVKSXztXrV0E9CWaWF6yPb+T+
4rVoBwNocEz29l9iDJu+fN9MeDwccbg1AoQEs9JpWX0FaZGLiTl11E5mRkUf6TGx
BYgA2WBXwFZbLGA9Y1CXisbrvmRfvohNBQrq/sKMKVE=
`pragma protect end_protected
