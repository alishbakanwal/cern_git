// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:05:43 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
gmUARTLNaJDHJS7L8NYMQ0+9S7CEEjmKuNB2I23kGk4LVD4cMMfVoirscBfJY2jX
xjsMxYnKTXchLqkQfM6eQIdOGX0gNl9baDM779Zg+9EgBIU89HOWadCu6BsYHwHp
OIO/HfbBAoLRycIv3s/WXYlihYOj0M+cv+htXSDH14o=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8320)
vZ9vfrfluVDP6Kpcp5ftOvgJ4pfdsdzf7VdHaEqRtgmNl1YC1/1GqT7K74SGIrHA
KLeuu4CTUxT/07gtEeBv5RlbwCs/JdyWLh/VqVCnRfSsWpF5whNJpTzonI2/VYsF
tEiW1BKLkoWfYUsSQENzknbxYhkHBlRbbjR2ULhAV8ccp+HL4jO46UfZMrZCYkV8
NVjqPupdGjiJEjioqH8ZTyjmYp2LPBXTj6aLnqElBq/xTNwmOHzQFvq9sVMHa7Pw
VhBKZi3f5mYq9Z3RVc6V1K5zqe5Lf4bEjYz7Bf8q3Rk9nvSEpoDY04ZxHWWlGux0
oPMbHvYYYQLhk0G23aIiLxYFKXiMfqDlMolOrVrb1tRMEAIsCXX2276vWp++l+C2
pu8pESG9I4eDK1AfEb8IvOt5Hq+dwwpznS93WZ5UBD+SNGiG/86gB1MT/du4aI1a
J/3QZTTTr3KTN242XLfCKZYaybQnpSK/lS2jgdirBMMgJQjVa3yK9kXWel1ipZrP
BJ43azr+8nohszR14zbsmBNU2redv9Mj9BVPLQdyAInpRvwaXhvJrFkAN+GqKfb7
Z+YeXHQrkGDpf2g8IiwWG5EvIXP+vj9woNwn4otZUgT5XDK4bx4Fpl/BFL/X8k0k
yCFeK5f1IJa9OSLhUuEPOUxfqjg56bfx8kb6lmhRFpRzFGmGlz0h1N5VBLoBSnRC
xbec8Ce5F+pmJZvr02iCmXgIhz2fINBv6KT38o0t246wt1RimlF8IT+8FhQeGkRv
jpNRDXZyH/8LpabYOVAAH8z/X3d6oGsb8WO8szmIZZ6B3SeWFI1i+8pBcT+0ewW6
D4bPJJ3xoJy2RJxv/626T2K8HKviod/7EdFtjAu5VjCiXpUYlT84QBsziyKwmx6i
Ncf22CPZQflGeO/58jyufg363tENrGEDYzjr8dqBP1QggDnpBDZfhfl1XM4BaFz9
x70YU6dM0HZ1F9+pJDrHq7fksYCIbm28gAMAG5GNLt0znUqexFEQNEmn61mw8zZi
n+f1GdGEr6HQxvINx4VIieYfdA82qZpcoLua7ktk8LPoLIvNYjj3NQWaLXTXJDSa
KFLrPt7x9mg8+SFD1RkIaX9j7kmxgYHg3rj0HWAmTGUx7b58gS9C0PtCtJqLiYb/
ZPgikChtRCumLtOZc4BdzjizA6ZiIElvo3wxuEV3WdOiGVjSJ0EWCeTzt0iBJorx
xu+3EtB1tEzGO8gkIDiKZpEE1BYxngj+e0nrntkRdMHLw0KqjtYCsNmLv9RSMyGQ
2+ANWD9x7EXJZa2nZc/o8iuRpRv6ak8UZnYmsF2DPbUU22r7gDmc0jUv4Y5zaJ39
KGDo/MRAY5o7MEUa3Qiz/CmvFqtamTrcC9tMNtetnyg7HMgSJIEKFgAFuVQcxb3n
9lSZyDurrTtPvqwMquga07z+U0SDmiPvSwq6gKjvQCY8+5KEPLPRCjOrInVyIAip
PyH41PPx+QqMtITeGmVbA0QI1JT4R03P3bYvElKoO9OXygI6dJPeBFm0GeRagSax
qtTQwC9mCT2CM7GMno3LxdGzg4XQIA2wdZvLN2peCldjFMBUincEVnPPCCB4FHSX
KPx/ulw1XnpJOUtomPaBYzW6Sof2gwfVNMrqtj7Ak+QaICBR+hpyOQFtEXiaxHmV
bY+y1P2xBkxfjxaaDNN4UzmP7mLs3Pzm4PiEY3D5SnN5ZC5ncYhmic16nImgB3U0
WGl9wHbJUFnMrqa0NvaUH+gvyEuUW1glGrUAAg8oYY2qU9BdWQfv8nODbvU8T9jq
JslcWtbQRdP21P5F+BB6QTY4Lz9I9LHtPdAkLLqz2TYsHtjkb3jJCf1IPOZNZVz8
2g48rM4gfX8lWdtZqRHLF+VVBh/SqPlleXXrI8wjDtmM9F2Ky7/ehk8MAQAeXrVi
QY7tGPr9TZYZlMBS/RIEcsj2BM/gYkPPONXz2/GUuF4Wi03Spce5VgyemfXLKYOt
y+gVzBwQYHxEdql38fgCapnL9QLzPks3EBNBb0F7MF8cDypmbucQkhZ0RO6skxPu
VsW+ZPeWGgtCfP2aCcD0vxOJa+m/Xr5PQI+P1FW0+9U8R0fM7FUfHIntOvpX1YQs
DdkRsEvxg3TRTITEiHD3gpJJV+ZOhpk51p+jqVJPqoLJ74jktiicTBdyjVz0bBgD
QTdb2Pm8VpBtgn7uDEgl79SDpwg1Ra/kEGapqzfVQTDnKa4yZfOahlt/D0y9wk0J
Ra0K2+a7Ky4PZpwb+LuLdUt+cfTtlGlwTGw8pQpDWdaY5xPsacmJ1b/biQBKvatr
ZCU15jcaDA7diOUbIj9di6Tf5kDPtnlM7UYY8NMfA0cBItUD6TzJkE7UxyAFRB7F
G6zbIch4oT2k36RFd3FvV7xU1Ejejw7f10VrI8BIX5/jULaBPJbYzgK9BjHUsH76
mtSMBvCokBV90LJjNoKOZ9HGOMzMoEYIm3KPtcQwjI/zaS3KbS4z0W52hp3X0LEj
i6s1i/0g/KqxmUmOhY+uePmBTDI88SsrxXhnQ7FNyCKNKZYARn+/KrKiXXFy6dCW
2e+dBWLwo9I4NLsWeEM0f5bDCFnAayOsZ4g/69hioiS4CRq4+MfXbaA3TYOwIIAn
ZoZ1wLDcBlbYl1kcxKV9XUL53WOuqsf/RiHHuCtX5fBXsnnRFxw1Yd7SNdF4PKBT
7anIfGMpAUBRO9ZRzvi2KkADdDEXxlaN5wkzgIGyXx9pdWZsW7AsQh/gwQWr/U0P
ZMdlVi4O6djM4bk0XMWR81e91+n56+LXZ9eHlzDjWOJ1Qqmn0Djcq0JjyH5QCbOR
j+O1+pCtbSqr4IKVzrYpEKWUL1sGDRG4ded/HJ7+8VZLR6aK0jxTTERH5K4+s6MN
9Sm/YgqRzCiG9+E5IHbwHm8uOSJ7irrf9gvpa6NfAFs48wm15X+BdDhvtvx/9BGK
BpXxUqqhRFJcAS0QqvCkipk70rtN8CuTpkwy+GRbKB51jBAUPxCjySlbTovZ+GCx
tKFqQboCLugKl8963eOn8GewxRI11ortpSvreL71Ydp74oIRX5UQ2XoxP3ihmHPK
uFNIGO+e0oAr/arlv+elCqtMHI9nANNPeOjfTXNsVmzl7OOGm0B5IcTI/wIxUIku
jE6bIXO5W1RlNFxeeeP6intdGtH0iwSpaGkhvzofh6gT80u0wxDlGfiSdK4b6cI5
7nk9dKJrPjc025DetY2aAUm22vqJSXXT7iWOcQIs75/tAggdiZt9cLAq9KppLOYb
KODN7RX/cFezvu0MzsUMeBq3D9pbf4zVorHqzox/pD6/PwZRngBIvN8uQ0sGE9mP
tpLTI0UHl0SOJraoVMjxtorNHonXmSi1wEDMLfl0jIaP8yIH0pIC7IXr9yW5JIp/
WnOKHAV2oXz08Rio9aP97PSIXDTkPttbmDYogvM66HzzraGAOzs30dDyPsGeXIOG
SCiL5xscic47IiLQZtTyxpRK4yDjzh6xv0SFUdlLM+SX4KDvvFxNGKTuvzI9oxCg
63bmr7F47+opZUxubuC37QxKIAEIuxn+TXkvUUjNpsIFMRJchQ7/9Zr2aFIJ9op5
Bno3a8vVtHadM2cmwNuU55xP3dXZ/u4/XavIeHlNQl/lNoiY9ePzKIkV8WzZ4sgU
+OfaHdHav6i5jdc4JvT4TsU6r12iDnraGdU8oj97EzQKyuzstJqil0rJe5OEX4UA
EkgTbmE2WhRk3zuB0QxExEeEJq8H4d2UdsSpMLPYVWwprjGIVZ1x7iEzXJal+jIN
8wTMVl0fEXVXmlkhmSc9pLunpMQfXXVVMT04ljRB7NOEtdDmWp410v0mA1yxoSYm
SZJP9SjEtu/aecQxy3JYbkkw+kvVAg4nKdGwQgMBFxeVJnK33MuNMpSfFxzsxNA/
hELGGU84XiDY0ff63H54qqgpVfxIvBJbRlgtnKZ2sP7k9GBI1dBllNDn5PMkIKlZ
K0l/THMb4dfdb788nQ3EL/d3ZA6qnw6C2Hour/RO8fbA7oTbwNVyrl7QhkF04IZM
HJ2cZStajzD1ay7fU0kVnABcMObKWCThFn2G15LNcjOSN+oiLjlsSgztluo8RcFN
jQ+HNqF6YDKJDN+oLcqt5FsBpR53ms+vUh2pQqGbcmLpVCOWhztwliVZww6e1gwo
okoUtn6sP9HJTZn0fO//lPTVz+jsY4R/VouKWvzo2qtM7irQEU+uBHfmu7z/d7kN
5/zShm6wIlePlOMika3EalRZuMAgis72ySkAP3JqB6mucLymbgcSzLrXi/aFejQP
gDC39jxyEb1chbt24ULUWijAKBd5UmqexaNiECJLDnPlHdjAwFwLKGxf46RuWTmT
QERsOMjPUXaL1f3I7NBkonYfJnksB6KYKrNT/B5VHHISqztpqwnHWLupd70cq44u
X1SdnMZ/8QosCNsbuBc42500cdeaqLFW8N7GxBjKZBjemGguEWmNE0QlTxM2vuYs
q9ZHBwlcXkkZyOG5gEPZHHL6hpSzcu0Iej/9AgcEuAvzFyKNI9EFGkt7h4U9gTGI
7gvRCeLoVBVXGZFzYRJdZocFLIIwcNWTdW7JKJFzEknHZDASpaj6fLzijPUXihY/
9GmyUX2/le/6GG7tL+TOIHRpHAiPlrhPa1NHs/knHldLV/hNnDV94U4Z6baRPe2n
5t7HxAloJlWeTSa1mUfzJJuihNIUkLAVsbJvMGCZVIv2XKK4pMYnOjcLGFd2Ka7i
dN3IZykTCJCFqdn7neSizALLfak6TORFhyhdjz5j7Dfpxe/tKSjsvAODHUi6xu0a
sGhYehd74lYeqAj5d9Qbk0eyevDHpoK9UFqlzw1cj8xoilWIXwJvpOImluXfbUkP
c4GP2foWJdbxuBAUIk+PR20OLUlz2Qn+b5/IrBF+ssny4hdg29MhjtDTuVkVS6VI
sFxQ/xBBM1Ip7chrqJEzuJ3lLvuTmTzVs1x20fr+z+6olCYdSSUdLneIRlgtjoiF
j1YTJ0vGdfbeU+yf8hnpLl55wotQ17Q339MO4TLzA1EvRHVBoTtlxZ1DHfrIHZAJ
nk7yKmrpWE12mbWrp6ib8zo+AIl5trmrULyjV3A+0M/r5Y1CB/JolrVAYX4rgFI9
JJsdhfcNXQU7wn2Qi+M/o9Y7rEdCjiPrZ+oyNH8gxpMrlJaZymyrY+TLb/8OtiRD
0+76rIdGUCJNB93nv81ujV4R9LIz1h2xlYGI09E57QVL53Ccx6pUlKZyC1+RFje3
pfbjkkUvVZNOyom5ACVkdc52TQ5HHESVVUpJ+vFK0JmRint0j8Zl72u01N4/g25B
xITx9rtYDs2Sg8uD+nl/hX18QKnMvS0ZyPRAgF96PmQ4FFUssAXt1ja8NV8hgduY
detRfYOoEtXexVs26mFthGK98hGslh/nqVQ926+ugJp/H5U3mB/y+PTwZHkYHw4Q
tuAvwwqCw7EJ9lJ0rdgkJduwU/xdEstfpWiyF9WqK/fx7h5BEIeAN5tmry55hHV8
gbwRTfpKIj4CoWKGgkYy7qTxF1qOTBJsF47muRhkBMp9H29NRYyAEIrXoPLicxkc
TZ+HcWeuF25kiciWXWFq3u87IbXivgo6YeceJrGoSt6U3yhOWHeROfJTLYjmpg48
yr0og4KU/3AZOqHXLTHi1s5beKgFCWLDxDrtU0SWz/kguK0sU8PhHOHphWdWNYqk
e/wyg5CPwp6lEqxbqwZ9JDzDdCkXlFuN696XqeW9OTPW/HNbprMR2iYSs1Kfpksa
7V1TbReHFD6Jto73cv9Kp/9pP8k4dbCul8CADaHnfgA041IovTmZEvBu+0UHF84E
KeDBCmnJH51OqmFIl59EnLYefLRjU3WGlXU2z2LXr5i/pjUwK1nwoCU+IJ4YRUbu
YVFg0PsYP9aZyFmKRNUMdfbLjQQCJDxpLHGHSv9oiQk3a9qymOhMld5gMgOd33lL
canELOSq5ssHJOPlnM3kLVhO/Wd+NNvqIxqQUNEZ8+hjg8LtCHQTgtDHoa16fx0q
zbzJitEbXL1bOQ8tpW0MbPwKMg5JlOdu8bLKsyD1eOxw3rsiyn0ScTzL+i7NBK+/
unV/3j04/oTD6Y0SF4JB4BSGNtwyJDU1fzCtZg7Vg0DrMrhZ9TZNSsUFwyDODnf6
xDxjvgZQqUogfdVi3xGEUWKoHD6uhTxFzgfbfkvhkRE2ZgUh1HzkFvIhRoRBBXXz
Gtkg0ynKJ85AewH1cPSrMnY3qubJRIoJ0rYn7eaNP3rwLVsH6OAeZKzjkcLO9REE
VBZakgNZFLwCU8RqIDbPWXfTT0cVoNCcUnYZb1V66KAzLhvTykPI1U/01LrLGYQP
p241PnQoUyJHwPYlgvgxxh6CZzR0sUaCZ5m2eHYifU7LdxqDe7hxIS8iOBzgFvss
M6Dta2AL1thZfmcmt1NH9hqcz2HgPAU2lMMEy+qAFbmVymV54rJMWu9ARK3Ftcbi
DpIuv4Ry8kf5qLlPlg64drCuirxkYu1JG0NXtgjWkhTb7h0WelQvm22tagMMNYy1
ucJjJRGGoc5V9G+wtxH2664ffMDhDAj0kiLoDWuUoeazBjjGKnMfpHZQlkQpXbRU
ER9TSLa1BBxtYEOEXzkPIBNlQZSRPirmd5v1+TKABVuIA4TMdw8ULqX0Fv9MKpxX
SF9IOCWmADs96Vqm1kLptXmXKpe0l9aKyd9lLv8ueWZOpmEHdSVlgjNgmDJOdOdK
+jy+SQ+Tw89y06SU4cvYeSM+UK+iXMp1pleaLB6Wk47y/l/pEUj3/MwDv+GCivzA
cJWI270TA/t2M+quPq2DUguecCtl6T5Ce/n6HOdacAJnVpUsrkp6ndD/MWiHY5kd
Bc7gyPrmGBmEIscQci86r/PFU+GUZacek0ymfy5TFD4cXFEsb3luScdOlyor94iA
FzQhiTGnQpT3o1VYnzwCIq/9Q//9y+yQMFMiuG/gSpzxEjyileRFXSm4tSv+6K+5
hXcValU1R89v6DP3159sZApk0GOcP+7uAuFQFrjtqgwN0S+7YGjoxMnrR5r2SnGt
6ntfY/QN2qM4cwtV4flBAomfreH1RsPezEdAc2WhyWTcwZO/j7tDJAHzVmq4JqVf
lzvI8rKIRivJMu1G+FSbLgUFdZ+1waBt3DHuLsMHN6Kf4Tvh7Qy/Iq4eVcW0wtAO
4waAyZAN2wV6uE2RGij5zTa/Co9SSh8JMYc4dKuBAfjh12uViftGA6BbsVUSYb+A
uihTkXyUOaZ6vXDyX8aiwuSAFutgMC/Y4cNT0h39oKhnoFXmqQ3FTx8ADX3lMXNl
JH80FPyLA9/eegDhNK7KhRoOlJ4Kg59ILcwcVaqu+F1CQfgNrOoq2wNkKt5sEe2d
o1LQYxKw0ZYdA76msqeQ97cWcNWGQTBezJ6fTkDiTOzroqDxN5Ok6CvUxhgoCC5l
AjxOokeNTwFQK+Jv9KoIPIDgmWj5IjifE6JcJUaMJxUFfOSTGfeZu4B3D6qvJ/gk
xFTpQPCfiitkPnXiSuxiGWPQfJGgo4a4nDA8fzLcP+lfDLhIGWte2FQH0umN+wOx
W/Pq8MzDeBBG2J3Jldqd87VFZQEQKnSfjY4DfA1TmPcp0hkqKm5PHdm3nGNqltOG
jFlQAAtasaaKLqHhyROjiboS0QPMnl/xAMK9VsW6flugRdIVwEUuijzbHGMESmhA
YAbmSueqMJ90re2mh3jStCmKOGIJf5HgN3lTmHRMOtV23yMTOj0WWRyMaSJGOEvJ
HYPgOdHLgoA9tuY7YNE7ulmPuk0vAjKKA6HOuu8QJpi+l8pk/hd0DVVzSmkOhS02
mTUjk0VfNo9+oBLf+7hpNA1qUevyr/S7muskjHEDhUl5DyTwTAItnLQfMd5bOWsN
lSiD5ZpZ20gI1OS8G4f4EgCh1lt5CzmsJdw5HiZWsU80jN84u65wgL4dxbyg+gDf
GegfCatp6cv090uwYfiiXoLEx2TLeKvYZ7y8az5rM60DTvwa6Hy/c6OyxjjMFYZU
sdrgMWB0rLD9x6lK6H9X2Y4bLTGZ480amaIr9Y96pPA+2ftmoDyHDZVN6t6LTRKt
kEhew39FYaKxPABFJj86LHiyFqdx16CuKlQ7LCI01A6xan1wgRQxHaZbPSJ1G3YH
0p3r0pRbeUJs8YRPjaHcMfcpvK9zXpvsAcacFdv4YJCtoISwgGlx4zZ5/JjPTnxJ
3jZqiXuAxXqOFhfXDd0KbE5I/uU78UHbbWVvLYiL1Nx1BHvuKaX48LUf8UXFj7V5
+2WcDOa6QjVAqfM6nIfv9/vDRJaYjZboYQl1Ir+u41vgj4m+1VRb8TCQZ9AZD2qK
MEofGnNfxZbF9jGrRZWbrkDuIgMyWspUl9pF3pEY0PyvXVMip/sja3jiy1USSqp3
yML+WeOkdP6vDHEo4PzaY+GcHUsd3XEJ8ntuNLu+tX8ic2r0R1t8FzfIEeH+HTtg
qU5e83PrFWe9wrvWrM+VOk3XMcGdAchih8BRKMc+2Rqzx1EVJl6fqc8W6e2RJJiX
We2MYBZHtAgWJ5QNCHncaEDsJJ+qezkoGeI0Ew5AQ8TGE/MKgqDm/j+FKknNkxAM
Rcn7T8S9NAQnIYRYy3eeSa7t0KuOTSue6sZygksyQZcqcVewRfQsZSxq60ZmhSVM
7uGnIeF5ggKEs2lwxef1CVJHRYdOjGHf4MZ2Z0/0VwmroeunbRAlByxKAz7qIpoC
CeSOUV7apYeUXD1v1lv49aGdFkL9PrkWBJLKRBsIubCgXn51X+6qSRxXZj/f7pBc
H8PfzYLOoJ1/3UXSj+i1kOYHpuC+u/AZ1cpZS1PPtKtFu0+i63xN4iwKItdlny/P
J5jVeGV6fO+OdcDix8ggOrhEtqklK/sTok8yw2OdV2XzsOH8dl5ySIPrWJZFanXh
CHgEohYBDSpahda6oYt/LgwVEWJh/N5c4En/zr6mL+rAiqPC/0OxSxv/tN0w/KEu
vN/E0uZNY7I9fX8jLhShFKMXD4qqy8Fjl5smRappiisVH92GM25y52/MQ1TihNLd
M967DM5U85FOiNj1Faf1jdcUxwlPg/XY8/LfhtJlnXGwnQ6RUcdQ0ar72CLtYufI
rwdPoJxjPM4poxFwzYSDTUOIMJAf4ddlCUMxD4OBvzHHeZQpFgehUXX6ZFSalbMI
RcbmxLDnPprYVXhX66NmKxzQ3TUX9EpkgZl/T9RmLa3CWbCQh7YH3gXcSpFf2azk
X3HC7YRGoH7q+Dcz/L5bWJf9xF4dyCGVvuTxMkJZudN0qeDyQDV41ioNlKa4Zkn7
KmfvMw7jSiAT/Jup2meWo6TIWGiwC7/cNsrUk/SobThVDLzdeeYVWgoQXUqSbVQB
qNWANRnsvWXwNPbW5wpeeAhqKv8y8ujVd21SUzIHRWgFvwEyVhbIFSayywaSRVyw
rzq9DQTtyyb8GrTY7A/sIO20KKpepqa7/DuN0I/NjYZpuX5kOAlqMJPGU9VEEdke
ZB+mqmBIULjRrg6IPDU2Msa67oWKAC/izlHLcG6YCDd1faV55ag/EwkAqoYE/Bw4
+dbeIejbh8Lw2htQQGs5ug0z6EfhXnHiga4oONvNb9TjMsveE5FEhxaqwltabhng
jeu2yjt5c7Ve2HXqU65ZBwOeczQ6euHJnq3y2PY+EcdxO0MeqmfKFroOY7zfAGCL
4tJm/ISv9+bjAsGbvLYn814PjXgdNX0sZh0jGnxXL54GrQxIF+Yj7aWRto4EVN4J
YUuf03kydb8VFJhePm6oNhwBTGbkgjDA7egIe1RF7/QoRMOA2ee5uoRt1Os/69yD
tt6YBObaRrRFB0CQdYlL+EvhcjDRmDK5k+oK6uKJeLC096uYgX3SZgDhnxl4NAC+
JWuqhtUloNA6/VIuOR/g6abDg+8UgZdv9aet5OrPbg9gHs/tZs62rjfdtN9FgPXj
bhrm1Lsc7GM4aMX9UbL7s7hdnFL6YgOF6dsiiwG1UV2V+ZY688xQEGlgk0O6wJbr
tVyMOjCoTDo4n76JFXDasRrUrVv/fjRFN0iJC3WrIfx6h0lyQ+bpIXHKow6WgQW1
oeViu0pIO4/ClZwvW2VvCtEOeR+n24zJUioMnQPIbzhFgiCY+n3keDLCRMPM3ONv
WTbmFD+YPbKMol5Mq2Drkj9Lc4pOCS0O47HB5WswmHMGQeNCMLIXsylKtvc3onhV
e7TFsTMNGF7BAX6aiUr9RwimmvpqQae7LM6rHjcN4YygVqt5Uv18kDJvYsHLRHeV
xJniw+HPmB4k6T3V1Q4MLvjuUqIyyRfwDlT+/XDEI6U4Zh/AYz7q6vSkpz96idLD
jfBTtr+he33c1rmCtY90DYtl4ArG/XfHcKT8OhhEVvVRzK1YmBh6TNcHCOE3btX2
nrETOXeMWGZnl40NNdeamBRschHs7SGVMSvuk//ucg1YTdJnUI/JeOpv+x+sedcz
LhglyYSMshK8KdQs9CySOGyynQc2RpAjWwh5VLX7ZyEPF+xpFRh7hfCvejUPpOD7
D2t9P7Q76EgOcSb1G1iiCcIugoNZtm0TXdo2mxpL4xQRDZWRee1OVeBpLL/14pHo
EwOiij8H9qlhxXgSDMFzYbTrhki9uDlW/EZtNzdofro9ftfYUAHtlIs4As8H3SWC
31skzN6M/uXU8pmmUe9/Si5FFV09cE6XXVhfq5DxrcJyk6E+Gj0oy6fLbStQXJTC
Vh6/iyaasMNlXhBx75YBDIph3MnUrDuqwNkI66lfMlJhwoEiOqebvU3ShCpsDwbA
FmDTGeXhf6VInzt7ZWY7iZsMnOlbzk/6m4XCHJ9T5o7LSgKHt0r//LgXmsZd+q+q
FsalPMn95zB7fjijBR9Ckcy/XRGi6KbMR/3w+ydoNQ+qD0+EwC7jXTC9xzmr8Oy5
5snrXG+Y2RIv93tNr13K/r+fpRRvnFbYrmZf3hjvCPS+I/d3nLGRMNtBtEEJUEiy
/q3/NQmZ4vdigct0Xjtkv3qYiQFlnFWS3uIKjZ2pVddGOZRjQKZ4shtun3FfHP/x
XKgiuIsoaZ5J8i0E/jOKRBiNxT1adphp+dp8lSyllPPcXZpy93fbakdNdQhg08lq
eCxPJpuA+QyURfWIrsznFw==
`pragma protect end_protected
