// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:02:09 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
EHIm961KcWNyIP9BKUUkJGK+XE6E3+jrG8uoMrj4eqeJaF2p+SJ0vb0dmbcCIR79
/a2elbK4nDRAHsWcqsbRyqc4P2Gpgq1Kj6VHI79KVYKm+nhgnCvIL2yNi2mbaIVB
OlRujyTraPiBBiZ+T4S4EWKU7pBG5DJqhI/1/7gxM2Y=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 33712)
p07jDUja8Rsrj3dC603mrpk1p7IrRTQQlij5fsOYC8QKOSgc9Xnfzl4tbnmXd5dD
yteKxWTTFbZP25LcJVMYZg4rPmMqvPZo21869Z/mYgbRZkYbrVQ946knJfvV9+lT
1WsmWzyoXxQ5cAxhe8WUolnqnQr4E+p0gdesPp8BdFHbev6LttrrcFnqQsArtr1C
v9rLiUf1QpuKs2J9tQPNBVtpeE7IXQ9KXh6FABON9aQ7rSjvH6NlkXr2OZOPoGJu
mx18TgMIvjhh9RADCewrlR0CT31gNciivQ/Hpm6Q4ZuBMfLW//yABccOUQkos1TY
xYSI5jAu6vPUMw5LZ/8O6m92iKXc80EeNWqpSyNyhK0NKvzCX3/syYdIuhHpG9B6
iTHOiYyutSq2PJIULG4Q2b9OQgBHZBnUoAPjZpE2L/RkBEF/UyV8JphRJuXlCbU9
aYeeCgQ+W4JKMXTaMaxZ4oqu4hIt8z38WZ8W57WjGfF83x6IcQStbJeg2AnVBZGQ
LZunHmwETIkQiUaG+uGXaKKgzEosBcU4OCa0xviU1VNXZ6iZfnnmyTYRC5ULMA0I
AIs2dottRRKhg37tlCtO6HaedMtmGDmPTzpgJjAgx/XIC5t1Zx20Ex9eJCpIkKCR
7ROP3odJunmOumDmaF4fl2FowVsLH9twzK20yIt6KvODhnJa2/1whexkMjoiJeeY
7kNH15wnb+B2PHHUkFUAjFNTUNGlaWFwzdp2UM/XkblbboMOLsbs/qaAbYdTEfkT
0xnKJzef/SCbUy+N+T9wwd0XR1nAZS1O1M8p9aDvXMo56gMo8NIG9BzRv0n6o/Up
y8QbTiWErCZ7ea4lc7CzkfHFq5kF+gWjTmOPNX3X2ii05gHX4vXD/5NsdEysmHrf
LVKof88ks8WAw5EhSgeo4HyPLM48UU+EvTkfTYAKfCnGxa2wqsnB4a+P8bM+VKLj
sys33y/lvUTXfvCaFFcN+CYG090ucriM8dcviIaLl/ILyqRaUhuwDTKl3ZCX856l
RmF7dLhBLXho2xqxxUQcM0YfmfAX7ACkGVKBKL9bR/QU6pymlPeySofPcp+FJ0ly
QFEAt86tDAWX6VbMtwhVpL8MtJ2Qvj7Hat/TvYszMoKHT0hL2bAVVCpRGdUKTw0M
7xZM0XGNPPDdQ2JDAaKmr1rQunTYcgP1QIDw/dnP0IGlCC1AAJFibM2tS384w54B
CiRAmwpqnQ3ZfUFWxMGKMGSpMzIyUE8y/M21NLXrpfRyT1oHCsxyaUjEih0kpin6
LXG168YhDCNGSqPDdHB/oYmo+hA4lkiV5YMPMoszkL2qpnithzbzO45XXcnO5eKF
XZSNpBiIgV4wgoh1KpWKlaDjfUgxaFr6nhamEv2VNp83DM1nNwjvIVDXQVZu/dKY
RAd2rBAwRHQrrOBb+IcBCGErPprdE5Gn0qRH6GvC2jeTt7+2y7SKp5jUdERX+Ve2
At6JbPR63ZmYOedhGSeYUZhAVzMFC5E9C9dF96OdExO8jtcJ302DE5ucineb0lSB
hXkuRh+oEyJzoxzdmZw86EdNFJAiRY6yf0Rr0zarEKbCbzXpJzglUHtbXgNhoXv7
WwrPAglbO2it97/rY+ZH8ZnxuEri3Cj3cZ8n5mmQK4e4nNkvZdKbYhiFJL+G2zyW
Q+SXDLo53GpjjUD+kzFgMOKA3J9tieyp2+lotz9Nh9JQgVUZyP2RIY7UxN5SL5e8
ok6CFenFHKCdVDwJI+rEZIDtbqpUX3tpFquElubMnViMNpKa8E523WVf6VVfIc2t
r+PQuX4wyLVFjOeuXzOUklsavNOqARWVaho7WkMoyoG2W37YzyT4d3SII6HIPUTW
6+FIYGohpEsvaCpvMBWywku5HiHxmvhvfl4/zEGpMYzGE6vG2g/yk+WBqMl7mE/m
DrzB7PY40jm35rinLCNH3B4cML5JgfFfl3fqK+OlzSFuhqoNhuJle2utqAtJp7lD
E7LDTtOy5htF58A1VzLFmynOaNRCRKJH4cjh+ExpgRN+jY+hqJGmfl4nMf7aBAI5
Eip7GEWYhQrHf6hdEtP+L7m2Tu6jEXm6T9iGrd1gWb0BXClVHiDPCHOTbUcLSqqp
4QskG3R4pHLCf4rcN/ZgmacVDJUJF2xJAn9ekTqoTp5mXweeOkQ6vQamncbrYHvg
GeNNZZPhFa+0k1kHyAZJ43rO1RVsmkLHkaHU2PdYC0QLzjSIPeAeHpPe55SKqPae
mr4FD9cuHxQSC7+twmNGpZmG2i+UMHcJJOTgXg9GxlnG9jVNGBRhK8PRfa7m18t9
iV3g5fro9O0ZTIhHdVACnPX8TFuZxpp3l+kfHPCSHEyUDrSORFUFkI10ZqFK82Kh
qZXND5prNAB0NjJSvNqCUa94vF4qfZm58vHT583PL7F3q5rw6XmqVxGXQeOgU/u8
t8qW4sXe2KFAQSafS8HuJv/QTqy01jocXQkhtuBbtWi6MCPqV6Mhk1t3puq2imEi
3slWF0fyNmmxJ9AQtVyvQxmBUdRugkh3mE+ksqv1SBmUO3AEvzEGTRRZHcsHzZix
hWJiLB/WS68DWluZMQrDoZQhoSyMuC8eG5CVGoCyfyU3SyfQ33UKi0hIPAjB7DU4
yc7zv7bmrsoWWj97VydDsKVHtY0dHoHPas8FeA97ylvqjZIn7+wlb3VSfyPdkdvN
ETHTbKUMDA5THd03lBJtcoGcDD8wX6sUfUfxnojANwE10IWMwYqKn28+u79VtwET
tUb4qs2P8QK6LQHSIMrctO5/LV1JI4B5UOEhtu+7LwYgP1irhzZvb4bTNVj3ZfyJ
JvSz40mr60p6iPaHTYRTGhEVfc56U0OciFatsAmUBcvOvLYh+YFNitsOr/moNnLt
Qg6lN6Ncwt10d5/K145IRW6ZEfc0UzeyuBcZy29epymhgibYrgOq1amZAN6zBxsG
qbHLpUytZKiWc+3uIjkw5rScVVRpDEkhUhaASQ6CkobAAWONOLYQg0Go8uAplivl
4FpbrarihQN9+p3Bm1+KtDzkwo4pS4WmiGKnFo8sSOzp6UM8odq4fclVb6cDovaL
UAKXEnRYEWHPPbKCKacq2Hk/GTASf5zrAdLUrO114Zjk4xqpPxXH8/YIdYF8jqGU
xhuF6p95uRfY5ORZPpK2iri/U68J5QzLd+R/1dT2788CNfnpcbEqYCvlBN6i5MjN
8OcZClCKpwls599bnAJLvmEEQCAYvmirvp7ZUoZ/7FTJF30dhB/8XSjlMiykTR9z
nVoXQV9o1VjjR7YAlQt/MG1vdYBY5VoG/QEm3bDW2WkX3Z4kxkyhgnvXx/BXUM8Z
Vs4Ay8al9oekRw+WT6PlZqGG52jLuWN1vhPJkJ3DaYt1tWNdeK7JgWfu7e6sjhWa
swVaSrr5xnTqxPkHePUZGrPXtu55m5gMpnhT9Cj/rYYeoq4YvdBuosTLx8vous4W
sKXlzcSE9vgiNSE9fAqcNMPXNRh3fpvR/8tIoYBhQ6MgpkGprnmtxbloW6EU+aC5
82xuioxF49MxMKZLZ+SbyyL/Sn+/UVYx8pOera3A0Dxy28qExHoXi7D4FgqpovG+
c2vkw6TlSJY0Kgdq7AJYhM1rY44uAD0W2p5BufwpeZ3o6yhTSgdq57YXGg9hj5r7
r0ha5dBJnHpyvSPHrisB6CmZW7FxZ0T1cWInWcjSbap2w8pF2We23cUENxUt0Pg2
d81IEC7X7Asfc3qQJ12y/r4BJAWLasGaZT1fOdUVIOTDJNrqWHBZ3Oy0INlxzw+e
rV88djsVa13Z259ieKXGfUfO1CRzEcKe4xs8rdCqtG73mVu1lLwZILq/h1mdt9pq
R/z1hq/fWdMvOWHi8O7q/oKOz15MKykYLw86GN+ec3XLqQNfsajibEI5tBTrvT3/
z42pTYrcShGQyiQ0uyfp+kyLpSEdCrXMll4bc9aHs9dMit4aUgDbtKYpmRnYoa82
rqN0Iz/mGTM+0N/u7VfzJEkUfKx+zhUvCTYWglGXHL8CPeXWjNqfxso9T8gtf/Rn
gV0E6uMbb2KxyRSUGuHIfewQhYzGwhp2EViY08a/p74U6PwVJj8acqctsYveo9dF
47p9EA6skV14UYgfjGQaNvwl5j6JO3xlsWu5GjDoGh/DRaV+Yfcx+awBKwIxQQJu
EtaWKLbSPLShclawZikkupuZNFjQ+oTMJk/O0jJ1W7X/yP04X5sSR+K8+2by0lnt
aooViokXkrrivSbO8sCJeSC6xFT22Si1/d/hvRljCX9etAeBtWj2G2tay6pyQuBN
qTEb3Sjk8do6VhbLWvMFMhXgqoKDU0rXn4A/xB3PFlbk49Zn7cPj3zJGUMVgu/Rl
FuPOOiXUCFo7KRBpdzwniUomic4Y1J+0+5lYMMgJ6Gex+P75CcNldHFFNT5d0Iyc
svzMBgs0WhLe7PK6lACNMROCidXKfl+br4gEsRLcBJo+faxOaYzfp29Mjg+IiO2s
udMo4w8MwruOrW32ZU/2vJeKV7ZhGLd/sVIrHH7ZWWceUzjSSazTABqyq76MwHWE
fLsbc57isYalGh4WrLmUcZLz4E21mIa2Q2hHS1WFHENzOM5QHZeDhUo7PDtRacKe
OevIDYHADlAQoyefz2Icy4r7SdQVQY1xTyduh/4QrP0Ze2+cmU9M0Ck0p1iowVgN
B+9e1vV4YHmjCuKocTsp29lWXyN0IBQ8LVV/1t4hZskNFcV+dz0ArzYNEnljIG0a
kzn09pK2e/yCrM1rFf+7WdsPL7+EWpRPyEYOAs+KIzj8paHm/9ycu2wS+qx6fosV
Dp9ESySlFxRDYnBYQ9paWVi+s8X4WZ8fRiVZa31suhAYOhGDEGnz3AZSw+/CPYc5
iJnMsBFHmL/c+ZVzbneQZjHoiWGI6chm9d/cn4Zeib+Vyl0+d7oTleQ3YcvJH1yi
Iva1hJvu+igkKbPgTP1Gcxw4i5fPdnEnPpxAyiXInGE3PFsX8ZkEfMdCHUC5q3PQ
bn7ZWegUrKjI/aFCCikTTF0ypEXXbmvmw4K4TDyEAlD6h0Mj8F20q9rwkbvUPzAs
ReM0NCNxzSXl3i84FAFTC1BAFQbLnj8Q6D5ddljO/ExXy8I9UBF9xPAGa1EQhG0R
/ikE26GvL6VZBO2rBGSP76nYyUUNCwy0BLvVuBmLTN3ISP4Ca5B5tX0d1hpZoHjL
pob04H4OE1iGDU0VxaPzZDILVcY5ERpzw89TX/vq/9KSQGy4qdazgiAP7A2Vr11d
20C5kqNeOoztBrXRmAgDI45W/dbfql5YcQXzvm2q9UsBwoNPvfUI+/d/dONr3x1H
q45C12S6Zrua/pSO+Sr57RpJ+n78F8eov7xm6+OlDaJkBPSxIPwfCaIYiSaaDbi/
xcb49/TYuRhO7Myh+7yV0AbO4JgedgHM35it+4lowWWmKKOHJB1N4xprmm3WRgQg
/E5nLAOdBYO9nGL5inY30Dn8JiG+CN0fAa0QbQ1d4QKXnP3Wef9y4i2/k5gP+89O
TqRh6JsrPQXfP1E+wC0oTDSF178wHJxZM+amMMoWsDYC0IjonsGuTvYT7VjSlwI8
6Kz3WrO0uc95c+PLr3K4Qc1/uldCGR+B2/4Rz7OF9fHVAUhORVDqhHfB+HyrRrlC
XQMkaqwH1761WV4DJ5SMTGz4RU1oJGuXNvUlLkfim0wOLVoR8DWyrlQRw+mR/qsS
w3YQxDekPY+ojlYmJ1noAY6Z5a46AN7tb53irgovGjfmB8bYpqqv+MEkGtrIsx4r
5g91pukX0OQj2E1sJdWGlybWTe/dL3thqcOMHLgD/3rDyqPgCOGFZwUMdrCFlgrM
nS3eK+jv8Cj+i9ntJZCX1Lf03tstFOZBCI2lS/PitW0D2wpn/vm+2mFZkFQlSzJ7
s4y4edwzH0+3NCBZcH7iBikrEMIwf/fI3Toi1bDEIKglYh/4ibe9eXpza4YaLNH2
jqA9rsBv/7snFz3Fza9fy1okrLQ8Mj6xbSvP0hddb4r/rpqR5oMtZ2D7jN4/sK/x
3SHiBCPPPymOPU1ceDCOm6Z3S3AvYkYKzq0KU6I0of+oTNHympI5CiNGhKMCDkVf
eVJx8Fq5h9jGOMoaUQnx9Iu6lPowV8sVuYAxkofcPLMd/x3fZylN0HWBp739jbkn
NFr+8KJXcux6DgTFXOjlAvHYDI/RvPnERnvDqfpTkDIZvghnAglau2eDSBgKsJg/
wIo1vUuFSF5DAATnAf00gcDxs3ctzZhT4T0PUXt6cgA7RKPYBvQhERVsP3YlSZ0r
unjAn4JsdQzji8W5dEOzleBBnS/VBeDcFnBCvqzbeh249KyRH7ti+bXUShffqPxt
lmsQahSFJzMJUu8PEe2S6boq9nN58hR3ZzSVctxLuSk6bqtL18LAYJojJ4lmub9X
CuGouzQzEQsNF4vQh3oL6nJ2e7bYsb4vXPSYkObaLB5HRAryafbYvj8fMyIZKwq7
yjfHNL6sKDKFxiDYed/TovqsyOa2p/qtYwX26mM4PCE7T+IC0HX12iz0a4UiuNs+
hZHGOcIB6h+6LjdIff/pCiVO31HwDI6kUwQs0+yAUkksajsGdjdN/Ia6RgoQxG30
KgHXdF4dPEevYD8oIbB8eE6gT+05THz1sCsEihqtw/l2ZdY62BFzc6hdWZ/Glkv3
nels6HTteJ0j0OqnX2CvBxAQV8C90iO8B88YsRJaRI7SOk2t91yG9Y67onxROWnL
6GWMK9BF45DY5gUSJBrLE48JAM1or9qwCdT/K3v83u0FSQAqRxh/Kr5g5j0T9Nzg
l6+VJ+UhxzaJ5r1kK/g/d99RdrppUWkBg7T29IAnxloXV8hSC/1G9/gDhYIaUZkj
U+RGvcEuN9jsG7rT6cEUPMizxgNTZz2rK7LkU+TTjBMp0wy6UEEOwRoNjqtDcef8
44N/vOMeHXWql4CQGdiwOe+H9MSQcFZZLjqma/+M4KaY9yANSReekcXjr0rrnBGq
rz4cztMYP5aHHGBqKIzuuFDjUjE9ZQ9wfRiCEDgG8wFTSdfEUUaVCRLzFURe5eud
TkDHgG9iKZSuuMfaU2+SpoGcXxCfDoU2LL9krU6fusK20h7o6IjcYMnSMnCxaILu
0ZVMSXFrXD14//lTSrzmE34GP10gbaJKLq0IVp78lb7zids8MtoH6o5fWThZ0KAe
N0qeOQZf7hZypJ0csTVUVX5CO+QJxrqZhqF3ylrBaXrarWWIPiWFbMjYfz6QJs4N
lc1nh8oasQqZ9aTpClvSe1UN8Hke/e75ntltUR766VdkNQawQ6/7S8VPz4KOOqDO
ymBtiezGk3DVmNqu3FVdxBhDbF/omWmoBuKatOTw441Js6iIUt+CpqrQqebc6BKz
rWtvRlcB9pVIjIvU7hj5AjYoiFouj/Boik64keAj2PVxI8tpsrTS9b69DwHzgJNp
Ja4Oja78b5omFonuQMYZeDPLX/5EE6GZK2yew4Zf0Jq4KI/aaKgJmbRC46twM8Pl
tWIkz48zrWbjp9PEbO3lWOr79Ax2E6fspJYd/0ox+F1StJWVikrHaKcVWTTsCtni
e//XZAaAOQFrIcid7W0BjFJTCZRLnHT2JDrhkeRhDuu8BHy7Lc8kmSQpHqKOqVPi
WUD9z8W6YT2HyNM7DH1YfULakCLlqXiDvmMfa88EeRuHqZiJd8Gok/+6Q+zaYdtM
l7f4t48F7lrYq6WGwtN8Yyu3StSIbV7JsKWQVcspGpGy9J3YwrynGS5y8Kefe1Jn
xHl0coG/vQrKGhOp4jK15NXK9IfYRYmIB/awwCe0AjHWsQpYgArrhVIXxKpZbl9y
eSQDSteh5v78h1oT5Om2p0SBmjR7CBDzW9gox73wLYxJI2a6ItY/2byDzOniav6Y
JpadspWyDVvazinM24b9qqIkvQo0mnrCibXTZsYiRuY5DnFnLi/MeuAx6mtV6s0q
pchJramLnVbvDjRGevTlqt1NeQwyxpkQWjBNkutl1bASAk7kGA0T5wlCFFObKETw
6RGM10PINSvv5ET0784lvClrpzbTDVRi25W0VlWxXz/QlixJKPoI5xTbtiWI4Tm+
AIneap6d/KgdCZMqWqxDRlS/KiB/eLJ48LVB0rUUqKUWJLX0cjLADUd/ugkgnblQ
cnBLzbHMcIabHYUMKxxvvVm9cjfxUTNeZppokJKl76FQm8BUnoVFEoV/4D0TbTY2
mqAjBaXai8pVJ/RTutKV9qJaKhHk949xPXS+u70Jvi21fcq56Cqwy/tZMFQrIUDL
8EZcx2DsLHpNGRfUCDrQAIxaC/AisWXSwLeUQksTRiAEIWL6mOj8tLJyHI0XOiEB
QCpUH/KqhSDVpEF7yar1jbLq+kjbe2bjkr3sL2KtG6LVp+du0TDsGM9f40CVVtRF
AhS6xxDh3+GjXioVOaeQVHLl/Pylv3vIw8LOEoFGP29a1dBi5bvN5DvmkKLl6Nmj
xfgAILIpAuu6ESnbqkFl9fWbGJ9KTf7L3TLjplQKWaxb8fva1FI7NvlWUohmrNev
4LvvZ2Vg3nobWNgdgKbT1emV+inqXCqjFDf02x3G8G4Dp3UD0TeOjkZ0E3rh1iBK
6bXGOLspkVNREe8PTjV0DUdDN41iLsLYV75Jbg5ZUXdX5GBv1LEEg8l27fadHtNz
jQtEWyXf+5gq0bPFZDYGnZCIfyITZifHnYvHfsknXsH1H6V5S9T2N2tPdQKEFaH7
Hs2PfRKykCQ2Kwi4YBXSH0Q9vSICvu734jLzs14bNwy2uSIUDff/bwkGYin5kPMV
PGBAniaMEvFbe2TjYfQHhQxhFGLKnSWeJz2KZpzw0zwzPPuwza+/N2YexoiXMc/9
JJRzawVG1KLn7uLmW+aZlmwvuRAwUnP3S3n5CuFWU9+9unOYhCUZa/X/7LxRwr9q
r1O4pO0mcn+AyWN+eYHvG3tL6iy3D+ECQeeTXX6LZsQeRFsHcPgoyizLwkOe70ve
9nTO3mgmDqJNLyknKXNmPpmOV5AGseSP7Ko6EvfbSd1nFOBtwglihc1hqsjHr0Y/
9eOgTu10Gw9rh2aklMExyfacMhaR047VIRmfWKACUwEfus+EG8bflPSJyz9HrlA+
TYwbzBKHPotpgwZ1fFqum5O7WxWPn1wI1FJP8aaX+OUbCIDhRLb66xcFGKYASGC7
Atfw6Xp4SvIns03ztiM0rve9hXs5PI1jhJtCBLlmdvwic20u4R7Qf06LJ4eAEkxg
2u+ApCrS67W4B0Sb0D3GiEvhgD1Ol4I0AVFJJJii+fezmhkzviAC4lsdzpZvCgwP
0EADvRAjL46AX+OfV4h9cYf5YMEj1ZCmLZw6veAzhSc0q/6G+ODPlELn75lLCmzO
vl+dIEPTYIE9mN5bXi2qdSpXrcjNOFHo3A5JUXHTHhRQR9mbsm+yPMzkjwV6Xh1a
uvE3aTqYd/+u4PKNTu+0th9KQ4VaVPIyrqb6BqEVOR73TpoL9G7tLZ9lLmQtwTAJ
d2tRMHrCvxZK6p9Ogbgpgz38x/k7zwi5FPw1nT8AJLgSkQaUzwncILCHKIHIQZKp
mL6aPHRIFOGEHWgGFmquOCBLQGCb6qjNjUEde8CxPpLR/zcb6g8Ckx/0aI9YTro/
ZGEMMqXsIjtr73rBJof41+2URM/6xTlbD3FjLGWkfzklg8K4UhCvQo85Y5vGXeOp
1jH75LE6+XTEW+Z55xX2IwWmJ5tix2zkSY4G0Tnl+1oGThHGDUPV3balwQTrevhO
rFeOuGUeUNY6tGbY3kcbkr60Ew5gPt/RIsVSZ0yxb6mux87Jgi3c+EtlSCcQ8S6c
pl5O9kbLctKA5OcPVuxJEwVQYUrn3YtHSamcUVflL8xSNCbuptmCCa0W8Ji0fXDG
hTTjAf8My8jN5uFJH2A14T6aPnRPN5CkeS79Z2GXy5D327pOk4dbwWOLMBemjzBE
UbLhIMVXe0Mi2FYSN9qbkbIp7slHV/Rt0+f1sAEC1gyHxEiE1zw5P87gOD5hICNA
B2Zyk/82hX1l7qp26hxjA326d38i97hTT3JOrcbm+/oi5NauwbUV6Up2lE5F8S7h
w+vvLwzAfnzd3E6yCntww5IWVSr3vOe/wqlq0fc4DHJ2aOE2yHYhEkdt1eN7lljT
nrCCCalPyOpILMJbpfByyZee6BToVux9Hu7XlpQurXgzJF4Xj1KFocpeGogf4FVh
uv8DtNOa/aD40TD4YhORJjOjL1alWqat5GbxIBnXE8U0iCaNG212IFjl8bxr7qxM
GvQLOYpQsXJqX4MQWC/Sksf7+meLhoLcTexdIx+B5VvZMMfraXN5+ISq09t8xfwS
TtRh6a4sz7PD/EOqD/8ubQVZnJBg5ARe4RHkndckO2DW0/NEbsA9i4+9gzbZfZZB
21YNpsaKnDV0eJH6kfPe+/Vg345MWNpWJxoo5LhKV+XflnVl45CZy69wTuDITD16
t/11UvvI/JHdDu+MqmU09cbvSmyc6TkSXaIrSNOfAwT2bXJunZFCXgXi6bJKS+0u
vd83x6fjPViDUkxSpvHzd0+AKIRs/LJ9sQzgPCU5im63fmVF5r4zL/5Uu8abTpSD
D4vCKf3MJ9fEf2P59nTOMitTPfSjCZsfS74MfBttqFmfy5x5YU9vBR0N4vP/Rdgk
drQ61FBlxWFU1/ne7o3oAJwtzMnIzawfQ08aVonqJBkh2nVRXSlwcyfm0CiDGaz0
2QK/TbWVkbFwKmIBCxpABPBxpsUgd2li9V2t6CFO4+3583O95294j+MPrBXRc6GF
NyInUG6YkwI7TvMJv2bTpCXVDZB/S3Ixk/GSIRylhGWH73QPvtVZmLRrEDfw973K
l7NzMD/7cm8SysAX7IMI5WwvvQVqaDOd4cLG9cT85eQWAuut1EvNR+8nOzwE6VxR
0x1ZEcvmvDEq6bAYMBf6C/MEDJumlnc6ufmlWasrxt1YembQYli8QFK/ykwq2rdd
CKv3hFV0sqKudP9XuoU0uef4Ig7pnWN1onVbKRb1SUhbXFq+GSiQOUcTYHsGxWLc
5NtMMaXYUbkFnx1KqbfOQx830WEkueS5CLzn1RRuXrNj4qXEdweTNgufx+yum4q3
rzhA2EFHu76zAzpcm/e3lkBN6kJtEAvY8F1QPzWxbir5tXfn+uM2kBqiGjF9STjg
KVb5Kt8r0PCdxPWxXfW+y2208ZhMWKN4QesCW/Kip2j973B/v1WYi2l5qBtwmJTP
L7wuuJxEaSoGcb6hBSK3o4GqabNojd+w+go1jlVJTLxFswDSjWc6meuzvbPbn7T9
53Jy8NU+vwmrW4lGVpF2G+4SDw5X2mFaFKxl8AITMXqKKjvxInVz67dnVDZbWfXw
GT2Wrjc6ovTx3YjdZuHwr7ayCotBpZoxxMbuBdOwq50IjS5l2+DHypfMxAsyxOb4
e0kYKGvb0qVcHDKNvstheIqsPXotDGdiewMFNq5G7b7DiiTPCXHgjQ/hcST1n5KO
CSiHVZAMzoIINCh1sap7YRhoHKOw9Os5PRZIH1wH5UImkIj9VFAj8+7tSEozgki2
NbAbR9+ehjIVTQCeRopxKX8tQCua3bucaqeTM+rn3s8I91ZCIptdKmd7eaBOV3Um
bSnvBx/QoJLQ80jsvvapnnPwwxSqgwZhfOfmr+xnnjepnk9qlbrjQ149nMQy4/SV
253pLRatGtAdEW98GU5PMeuARNxOU6Y9NW/uG+KtYbw5mCZIfkONz+hRuM4nMfst
AT0of79zKSffmCTBUwHJfV6CPn+DLvDQb/IVyour1MKCX3B0Kz9hY8MbCe4UgRTu
SFEyXW1W3iCrysbSVgi3qbJKZw1K4LYJEL6KIXGYeZb1cq+U6InxXG+ITqIEP3kY
Nc1Z4UOquCsJ7FtyAr68e1pL2Yykhs/XlQvI+LocQYPKJNrucvtwKQJrmZliR5Vs
Exc7ZYWdrX3XlXW1f6UA0eqy7GvxiTa48dJ7iRdD377G9MH9oMtLwQOhhmMhlHxq
kvuNzlfN7IPQPYgRNrs4X5TbYSHcNovDkJ5Nur3dUZa8xlMUjbDS5Nq9OlvpLQiY
ZzZ3CHXNYlCQbho0dE+mhyBhaNuWjeMR68R1l1QuC+qz8EaE7SY/H1RGyi+KWuEK
jRzmcq0eHbWIz0wwA4QamGQtiTigtPHK7UXrASi97m6IblrgbnJddcVkNgIFjAnD
XPrl6VFUb+pJTHnTIeXlpNXVYUF7AqNGmw8JBzvPOOxYAjMlJgO7zHFksl/an/go
VZ/1zGO9dQXU026uojWM3SYLJbIZevHoHidt3eqhT80l9S9U8P5CPfGFRrAdtPkb
+3YsgVw2etQgo0vh5JEiCyz4NOTaUzf/3p0KRAvXOl5c0VHl2TEdwYVTmj/JWILL
44xVaJzQnoztUaIcMmNVfxpFtCydhmj+jKVqBfUNYojFeEaJPm6ZJvGYQe/1JYeb
v7piEcrOBvBKlrQ/VUKUTvGXrzh24LytuT3PzUTuCHIk2s2S55tt0qguV0jrCBTz
Kke+0c12OkFuAt1mGl579mMavFfUNRM1nC9BN1HNBjqOB+Nvtyn3dXrqLMYJtG7b
/JTEBXu+JmB4JaznD31WMm+OoSIi7caFLoTjGYJkZ43dlFODenmJBjqt9U7AmdrB
NhrWrRzHVJ7I5r3y0bbexRdPYoG2ySI2tcePDkegCOoVbwrHOg4uXjEQVhdVgo04
j6lcVbgP2UwBAzyJcqh315/hIVagcKx44dDcvby2H4wRFuuE1yb0Jn//dYHBq183
xmWdtEQYvaFKe9I5Tvc291IlEr1dadsT4dP7Qfn9ERUtU0v/6xEuBHxq1KWoZ15f
vRMROgcNYpY8wcp5vzrZ+Oyr31oTcYuLeWI8MIjY5g9zNPBkqvimVIZJh7dlm2Cg
ZrRPZkJix0jZHESFQdkiu+feZoin8dh62I51T7uX3ACETR04zenxoNeRFAWvOJmv
4yJgX10Ezua2FtoT+igWXjkVu3iWJOf0YShYGBO6Cmn6/TXjCTFf6JVYDlSi9LcU
5kClqgr8zbuU2zJu9g+bKGXtvNxRvbH4ukt8ZqWIOziFKOjwM+xGUO4X1HPq/+zN
newXAMNeUWrAhoum34s/4BGmmvKTrPqixCCqIFJw9SeCXAjPR4VHiCEd5o+M2QlS
HHQvM582iw5zMR5bPKfO+YgLooAX+nJzq0O8jGRfFBDJR24m7No6BbjpB2ZGPSzz
nWYVzGNm3J+fnyCTG7n0bWKJsHP0tVRwTju+2DzLpb+G7IuSa2ggBZuW/WagWbNi
C/8aO24quJxdlIvOGHkSZVSD/PQpY6UBBVamLuw8G6XSOSfD7M6SyEiuyfYORJuN
WAKsZoD2wrVXc/BAldGF5ztq6S0qale+VaXKqFmkH+s6nJJE7+vlsCJAWseL4Eac
Nir/Dr2GhpYUgdgYhIhUaJcaOcwVZFFtXDhJWvvp+tjVDBIydjfK0ad20h4OX8lp
rDM7L9rbwFpREde2z0gn0LxsfQqECpey4r8JljK6mRaZvI336BkmgFsTDCDYgmio
GDx2NackfyoIlkFuJp5HQvFfyjM+wd4ZC1yWs1HcMjlARoI803x/jusV5mJwCBFM
4Leva2ZWtAtg8I8+jE+gqzkigoPYM+VY1EXt0PV6ZbHd6hXgv0V6yMz7WhC41wXc
NvaU1kNkSOfKWWp6QnVMBVnC5KcbZNJ/+cNDYtcIdTLSL5IwmcZdDK6EDs3sEjR/
vqVroaH6dnUEBPn5oSm92agSkEXwxmd0mT7h0KCkyBu35yzkaFXzDelnuWz5IjSs
ho/RJMWjZ07pJ/VZjKIGwL1urAeo2364Llj9c4F6uPARL6DJeO1+g16rJ0q/OPAU
WWiF9VOdBq6oYQKLwgYJpjNnUfXl2M7rijIE5/eyaDfbWYI0xdR43TQJYXnSJZjv
ErNiN3uz0YLur06aUUrQuJOSoGwrdLvzZOBT3LJrjeIcI04COMyzbT1Yt0uy53yl
lLgWHGPhHKtrH8d0EuzBl6A+MmP4GHz9v4xVB/l/Xsd399eaxHGRTKbuKSimrZNU
1+H6RO7/vi1yq2BjCDKWk7asWrUS4EH7tJzs+QtJMUFTChWvOEqBTGJrp2MpOp7b
lBtV+ZI5jV21m7gQfk9wG0R51Hfq1wBXYfWj/z6NCkSlOs6oWOrZ2oPzgZ/n1xnk
CbIZCYJPveIbkndF9m9e9Hi7F6mswSjgxWA868szLvja0gxSJyQmTKpvm/N+9Aq0
47c6lJu9YnBDP5wi5mlprTtJBsyAm+vF1GyarsJd9szgiX6s/eZ+9OIvFiJ1C6bK
gEV+OLv7aiPmZQnmvTi8CEeZAuEYRibN4PTYnd8Yj1VNjH7Y7A7jt8oSPKVYTSF0
YL+3MdOeYyTE6XN8idlJ6HBEY67Hub/zX5NIbRihk9miudGrkokDYlhuof8X0bKm
iuJ6ihlkahQywJ+v8jaSFpsXkRzzPnCWgyhMgKSTv39fI8J4tZn4n1NdNDCsy9yI
ysaDf1oD+VuT7Kbx0YEJylU6z8VVsTI2dc6jys0IQzX7CkRunxrQqMVg8Ug8WA2s
tFDhdbx6iLWcSir5iomb9LXWdQTHBuWUuSbITI/f/3z3UxzaobnUaVlu9Y9nbwzx
vsTuswbfGpuYnRy2RiUrYyg6eLq/NKHCm1xyJI9EedwBN9Ymnc5DmbSzLUFpVvMp
TCjAnMassBPnoeVKrymCCNaRO2hlNCXj5tOPIQXNu1b1MKjhbbsPyg5g0hbOEmot
aswuhzaN03R614Q/PY4rDLD+7x5MQZlhqWg9nVjMO0QyabYOWj05BbJYM+SWZbhn
TWbncY71Wex3AH2fsdYT0APf0opWQXbeQY/tYsZDoy+zyrmYh/YB9T/DS4vnJp+4
wl6xKXUBdaPQE0Ssme9WQOd1nzDCoE/fTzswrKpOwOS/6nU0uIWrSKYQeS88D7ma
FWK/xO4d4Q3U4OlUO6Fc4sVupSvfSAvKvHrmQ5l6Cc0Ywi4ZS1jUPCfhc1Cr/6UZ
zB+lMh0fva2yFBT3wgnFnsTzLnuqfD6Yp8UvtkyXXAjn6I9c0FWYKeLt2mq6wbOz
+/fxY1AvtfyqiTubTpzMIfA8yGJp8fd/qyemqVAkJkkNR9XeZFcIiJ5G63SBpSWo
cDJhJPhxgGBZYN4imJiiP84GniMizecsewW/xgSNhJFEfKFrqUKQNErjSSulAjDg
AHNcvXB6tM7WV/fYJjlif5XWBrtfrl+9DQ4RpHbK0oEQCsb2zc2G5Lkdb9LnuQCa
fmKAmjeDd+sUA4uF0YWfmLxXJ7tuogj92kyPiJ7q6g9aJdLxbtUBJD2MHKHN2HGQ
pGPvn+IY4JYBIBlKecCS0LSNEIHmh1HP7i7KrwoqVI9X33Z9/x7Tr3JkpBbNLGCF
qsEe1PRkEqBnZPPWtvb+EFyQfPp7zP9rwtcqqX+Q1UlRFSLWEc4lBjlEHQ9vnF1A
KgpO5NSVSx+1vaScx2+SfBNNvcmg+nJ6UtHw6SzduRmcB5bmb2OvziBcoJwDd4dT
X5NdTA3DVqy94cmmhy2xJ6uXZJuYJadd8Py4QDJ9d8vrniBuKZWf5/pEA4S3IJen
cqWqEK3DWym8memgPuLjU1Sdgh+49sl9VypEvTaCw+B7VIaNHtouap5ZB9Q9f2kz
xFbfLso1dsjyTgbDDuSr4ojE1be6gU9cnTK+rMpEuRODbWKDGaesPYiHY3+E7FGg
y7yExtwU/wRyyDbvMDirp+hJuUiQLmJPp6Gr3wWDPetbLMyKOHt++K0EFFAC2eXC
anzhg2JwTyGfczk/pZS/UK1IfuyKCP2vflUun71op7y45yj1t6+67sbBu4MMcnae
JlLpgXOSfoDCuzFYELZHo5D6E1WSzlg/9Pryq+gOjD0uOvoj37R0ZcCRVflfZ4wR
wl2AUo0vhqKiypafHrPAdqK7WabCfozNsy898dnoFFKc/VYJIeNy3tCmUWmHZIap
VF7DjDbyIRVQMs5/Yl1rxlX3IVYf+GkDzo6kvoBgbXmDLHv2mpxZUg8e2l4vF9Sr
oKhM5fTxyWwS/1DiQrbwbZgMG+yg4opBoOEXMBCutOwl73J2fSVQ9kP84pYgCi+S
g7wk/FLKcXcOXmAGVydJx37lcZVz5P9GRsFiLQWHn/6g7ocnoaHndDDHnndy+gQ5
qJjj5OfkicuJo+07B2SoqN2ASUqsxFB984zFfQPoGcJMiNGEibAulSQurTX6aeVO
fEZ4+3zkhafxstB/OgTaYzHragxvfMCjSC88/VcvE/iurgSAwH3gmVnXdmvaLPyq
pTjn0az7TRuq9wIP8GHqE8l1iD9zCsEYqjSckp59qsKMzgTo+jelfQrbnT+ZTKzG
4Gs26Z9yCchiVIqe3eIeebbVVz3hibHa3i+800qskNQ6t3uS82WLaREAdkx1rooM
biO5c/+ONcDwlVCqncKhy6213Do7m3SP4SGgnL5cp5vqpUS1BjDRUea9ctT5Tz5x
rnyPpvTGE4X1d0kvVgV7PQZnlihoz8G6jS7Ds1RHqOEAlVQvge4WOHFTVoRCHrGT
1j8910BjwmmP2rE+f4EYGlGZWryIEX2SYTS4cFHvfzrWKKEAHvPr/OpM7+AP5nNX
Li//F3ohrKoNOAxQ4vtf28CYkswVQnY/mnukScTFXGM1oqxP5wOiv9j47ttx7c1S
Ajq3gKLpHt7iPRyhSoq5hCRx1c51ONcej4UKV5RCccJhMeWfMCK/PZA9oTUSuUbl
YzcN1FuP1qB4jiDm1+k56AEDzQ9vFxcAAOtxoRq/pBmnEkI/Lg0cMZLj1t3PVq03
zexsIT5h/k99mlnJFawQcMrFoNuz9dV4VuLIbDulwz4XhhGKdkUw6b9DO1pzfxW6
0+Sc2ZX/f2fCV9bTGefl2taHqvIIhKsHe7EwA0RHO3rMjuQ4/OnZ8ARrFjnQ79gU
JTSFm9IrKCz15udxM8tlxie4bQXwTj7a0gbKoIWKZKxyTIFKI0etOckxy+JgKBck
SZnhDIEPzX0DRsxWKwVQ+w6XFVZOSeYFBylvWkP8IZC4XIxpoUIOXuprKi2V4eEh
Pdif2eo52Lp99Fv6CC5wJwAO4sjJlx2ZyoP6bkbcI3nWLEwoYeG7CLuiHHSb283C
PAG+b2mF9dk89RYVjnC3BsR+xUkpT5ycqntGDaaZ6PDPgs8SOUYcWP5pSC4TNDtK
bdJgOxQiGjegvD9CNpzBOb5h+7ESQHUZHOaynYBUf5yLC96Dpc89jcbQrpeKDA/w
6d7BMVT9k5OHHkOmEVJpEL6h9uE0Bqfq/H7mXv/IxbRODhIR6aI2txYJ7qNCExAc
RFZQmSw0Xb3cpS+vcdEcZXW8CKU3aMj0mK/PK/4g/QjHVJGHIQoqvklo3yMxq5Nd
dxPtmEtf7OSCivkSPjwnvt6jUofSTQzQ/mK638v/aw1kQ36ZrSYkh12v868bxy9F
13Wnr6fRxVndg3WbGexdINNfHiyYWpDClyV7LlUEnmgcBBI2mbXPxYmNDmCh2IWA
/8Fa+d3Yvj6+DjKxdSd7mxrlBEjTlJnEovq1T45ePF/enhN+opHYubyqDEsC4aza
GABu69t/70+QDbJUBMtn5W0t3sgBJscOvAtQ5MXRnKf0aHM9Sw+UcYsBkjhH29D9
nz0PdyWfi6NPZo9AdTgfgRpC7b84QlP6fz9V+JrcfAfIfNqhxlPDRfrED5nbQZZ6
Oqcx3VyW+XDrApJoj41R4BG28AqSPiOpkb/UAnOfCzPt1gNjDmdwTSK1dstXT1YD
DyyLfcVWPpoFGn7WKfV05aaqt2EWYu7cTc8hZW3SuGlVVqPll7h4VbYO3F7vvy03
Ono/jkUcBRNwRlxijyAKS4Q3BDE9ZWRdyuxD/O/5MWU4PPoDqE70K63egz4uJKzY
dOhKjrtbxy9nOyeotDgrc3qaYWbva2wp9l4ths3NxSyHdmbEjcpRCAU/npd+z5X8
3frb+HXTITXKOZpAbQPufkHaUX4HvL5FiDz4kCB2pBu2yCdhZ3e5yp1ERsDx7cLL
V0niBxQnR0qPulMcmwXtLNtVuuJ7cnKAFDp3wMUxLESG0ZoIMEpSsKzNAZlRWWT7
zRYci1IYrkRMPC7jusq4nPfsLUBPZ6oUhGdZC5U/yCIIgF0FTy4yDdHbwMJke6Sk
8oivZch4YpNEeH/oRl/N+Hgvfp0Mwt4gQFKgeRLzTFlslG+kykD5oTryc18Zi0Or
djel8UAxHNLD81mL557JgpHjv5lmPz+TuCdozB5Q9JbZwjNgq3roFs3XrX6nbLZx
om3B/0YwYmThbDV5Dx5adz0KVI6AywEgtc1/uVW0RdO07aUqtkeKYBU92ZMAiO01
irnjz5ULjTzDgnkDVJGeTJNHldhH+U1rtfGMWAcVYR42hg1OuYvFnfLWywxIA9lz
N/KHZjUhiXFi/7UvcPQeBkXLwQeh8rp2k77EMaB1HjfTk7N8gT3GlQQrf412U8wv
6vWN/txNQJBRKGjys3YeYAuha8GlAY5Q9O13g8UBw2tefwoVNl2sYAOugnBVKKAb
6jAoy+Umjqs8fSLSvI9Wtom0GjgfJcsAPzCn4DFsKJdRA5n8q5LHLyKGpHU0NXWd
tGEvvQB16pEEIpYXB4kE2XxHb9gUY3a9PNNzynRVM2cpwaUQsx6noe46hrX352Wu
zpVU2R6JhbpFDTvVAAvLWvup8D2KXM2KRo85LK/h5WeSy6GQHp1boX3cSnwxaYzL
XtEtlrsmcSQ5hrBL1aqE7kT3d1THlJbaLXoEjnXyQuMoOZlKU5xwspFgwrmpgACI
JFprTs1XT+p4pJDSrAPsNzC5bO+/FDbmg1ZIpakYX0lglkJUwfWpn3tZ1HjUWzUb
LCtDNYLvcP3AOhs1CKWT5MeWvGGnnsOyCn3aOzU5Qayx3K+aHECRKotiTawgwt1V
vMDaBazS0VdKT3+YBeAhLzB0xA/MfKTKStAKEPLb2jdkxEb8NxbdZRSqWDUKWH6e
hyKRizX3Oz6LfAwWstODT6gpa8CENRRf0PWgNepjfJjdPtsQgWEJUVRp47xI3lzh
dYYqeVHOUKG4ciDmc8Vp2KXGCgO0yoDh5YCqMexiTphnQt6vQFPnTmvrmhBAm99f
Ho+dP8W08P4bq+6BaAjFc++6vjVdtRhrRvWKXSVs9J1ItJ3iSw30QhSzsLCzUGt0
sue2Qb5w1IOlfpmh+goYGoK1cKsW56yxx7TOcHLD3uxwCooT8sGjjTwPkFuKSspa
HXLf0hQGbR3nVcb0QjGjsFqCBfcV2OmvY6oxctZ/KLL2eXyLsah4cdcj6JuvxFto
YeoPUY4IYLN3JDYceAtnjIt9VVZOCjHwQPX7fg8BgLvTMVlPZs0dd0/dEinbTEsx
MJAxChTIawebcJjS8Oc6WpaWtQen7xjs3AmfLDqG4ccv8UbEdGcTDqB29Z+MLWPi
yMA4SN2mmVXtMNfw3cB7rao+nDXvhP5ozhDFpsU1popzVrw0X5txxgVrbQBZASTl
czL6XzMyUNjsJaMkY51nHpm2dfWhszWAQW0IQJioQfVdxZ4og+fQGcVJwpDCAoZF
vvWn3Ffm9a2mXDnlgt6ySk8CnsnLdS8Mr3Xl66NpXvh55vOw65aby4oO9QR5nWMI
1F2PzQ3BghkDyfWVwXewAIKplgOj1wUEA/IvQEnlCBeX1gGCxTN4WVijcO97N1yA
KxrcxBe/qDuO+xQVML65eBlr3yQrrNpLZ5o2lmFbnP5vEvu+rTniMWiwWEK0rD0v
Qc8gTkMcZ3L0UzLd2HSCcjBDGcM+HObz5ed3V4fuxksZt1zMkJAa3I3hEwKQQJVJ
2p7BCDRgJqb6uIy6zc5ily5RnMzl+BwnGTWJImouXEl+b3OeK9swPmf0GHzsuF+D
SO6eur0XTSprTRQ3gxTp+8F4NkQKICcIlzd4gzGk86U21ouUDdN1x43xFK5a1Rug
PBuQySAC0pH7nbBNPm1KBoRZFdL/P+dtUYGKWiQB9EirTFDLeIbUQPyzYX5rLmR0
GbkTs3t69BQcuRC/1QrjQRgCwuQHPfIjcTNS71z8ZGGbRi+XxLSYQyxaSQ4W60Ey
8P9naCpJAmYWroOg+V5uHrZ3hs7RK6kSOzNaRAb640CmMixIdEezz7Gc6RTuXnvG
bvltv6c6iJjw6ehkbRB/lqWLXhSHIOzU72BnQaIoNtAoQmEkPL8o0DSl7ih5cf4z
QWW5eEfVwnhAQgp6lJEpDJeXaIluoZhbQUdgebbk2GTm4n2P3tq7HHkAPdQBvhOg
SPT/X3d4hM/GL5Rpa3nSy89vSj+KAZnsY7XonZYN+dIKzRRw72t95Rn+osd7CKn3
B0wtAnTfO+ra5/khSBuo79qM9+vT617iUBwHzQ3gdU5Pho1AdN5ByWwEHN8EV5Cj
hlcHGDPwWL21DUZI0L3BXypHVQQrlmrsoQ+NNZUB+I4uyeTqCxyEfc/uzgRg5uPz
RZke9NYY//oK4H+xoe/Lx4fS5wQ0Ki+MXBihRZKb2R4z0hbHFzfhtVq22lVZZgRJ
1x41q6/511V3f/yDN+r5c1yyq5yiqhGm8sWu3UOVKwGoHH4GWyOJyVFkCn1WQp8e
szpfvZyymuS6XYefsT/G1GCb/ZxX7JNkwOSVtcVQ46DmWC2cDInBIlBl1whETYf2
e0aIATLEmlvGNH1R+0VS6h/WRh6fTezDhYTM9mK9xiyHOX6zi1dG7NOiYrC/8GUE
VUIuc1EhCeHuQYcMc9tA63vJEAZ8HflLgLQBkTZ9lFLJpRds1NHEbV+InI1DF95H
Q97NMJlZFd9HYNH3H7vr8yMp7zU3Ar9UaeVrqzhPMLP9bgAXSTdjsG7q+K40rAAI
m3nrNj6t0LUAC+O/vSIEq7xqjXOvq6iNp4MpJvauyR8i+cgLwKVuHiZ83wHefaOm
BFRISSsf2oZD0C83LFldoHVEBfs0RU8pDYSuoi02YdzbA9HOEv7ayqwrBZnskr+G
e/sRBn/5DnJMsb6MOF9wQZ0ztIYyici5tzdyjD9uSu6gSouq+XJpWnacQvskYR61
6SBR5CJDqMNu/MjIP367zl1/pYzIyy/6C9r43cLagOnw9NsluWGeMBWGspwHakYT
CAB25lgTVk5xUAcKzacHphW+gPLuvzVgpavUE1oAyg3J9Wep//BM4YvSvXDiwoWF
TCW4UV2JuRoFVT7+M3p/0Z/cDbvLi+lA19m+LJT27hxland2iaoDiblN/Eohz+Fx
Am3ts3NL++S4QFG+KqOP/9pk/oCMciN/iFYBSzpYa+6kGYBCwh7Th9XXQ6zSvkgw
pAmVRRbGD3Uz30RbmbFzAA03U2tO3KpP4foXeZSAVlvQHBYEUy1x487xSdqVCMU4
HhD+pc63CVdGbsLdzTgGRToXYGeJJOlqTRao/EnX7/uqKxtzto9IulL+Iamt74pw
+GCwlPiPUw3+3tKGkjoVbGN5mgzPhf+L1SlCm6puLT371RCFZ4jPnQ2Z5GBnHbHi
uHYU755LyAaYPrbs9l/D8G+EsF2O3YOtzUxmVpCF1cUIrX9aA9jaU5cD9g2mnYqW
Kym+0jvm0AwGuU9yOTkYAS1pF+K6f+T0m80lDVOOzCLQNrFAJGQs++kwxxtXxgnZ
k7CzQ+ckaeWkX6+YdtidifCZyX2IHjdjLEGtAqe8VJC5/UYuJw3muAKV+tXBt7fF
BH8ZiReNu1UBVyLdlZSHPBSvO49xRUwY8arxfGrEi7WsW3XaWjt67snUs9GuMGUY
JBNNVt9K5hoTgRV3+kff9F34Hn43HoNPg9T86mF/tUVregluT7nIF643KZPAgpov
+pTHZAtQXzuHu5oDDVkPdODobggMBrV13mEeq9Ku3Gddi1Z6Aaur84Hbl6C4DVCe
MXOQTxea5ZA2zqDZumtwQmP37tGPLpJ8XTbG5UpRFFNKFb9W5mz8jKXpSPxY7y+Y
C/cA/SGkXbGqBX4yj9v6E/4NN1k2YWn0kGj6Bb74FfZCw7mvsUUQkHKR21X/eG8Z
bwDTRxkkYvXg/fwV+v5bbYUjCQf5Di9C95zU3BFqNaUTyzjpwyKxUq9uhUTOK489
5bL710+2hNt++MRESEr8GdPIbHnqCFb6BL9MrB6F3S9+0lY/S1YDMSK2hrRqwvLG
sOX21j1EXR0FEYPV1AlEezdruXcjWrcYM1Aa0RPavL+lC6YCWidXA/JSPrDM8Qbg
RUfwou78JMJkBJxykSj4aeoAMI3TjG6iDqN7/C09Ax2a8Npc5CMb0fIX5J2sYlFk
CVR8fv9mBAs0iXbo8FWyjdpAA3txjJtNVly4YaS/0tb6u+rP5ngQebC8WHjBKAg5
mAbrRAw+lXcyg+KybSDISbwSF6sgyMDq2aDA+JV17o4AhJqavwMyiS/jAsGDcAoc
LOjJUG9Znh9SDsW4koRTA5iZGym8P+13/7Up0/u1dSyHUE/wHVms/m023FVeJKLX
n9xXu5/bh3PKZpVXXqGtrX4VDBeLuf+ZliaHi+m0Bq1BwwBOv7yYKHH1atQkPouk
7KSmGlp/GaMAxLn/NvlYRifeUHspluP8bdG3/tyBqKg+vIq54k5u4/Nl0NORqv0T
JCL4h1SVPzGhgjJ5qckfdQshv/4nEf59NwunV9xMia8h+wlCFrpGO2qe/MWR3f4e
EiyMkWSGj9jplZSIsAJUuhEkapotuj0aKv8dwIZkGi1SydapRt6LGr7PkTbtLqPb
d9Z5bUeX8fKFryhbPBN/NAHz7nmxuSfD8dKQTZHwph9E848HyJsjTCn/iaKEmmSA
Ry5ltLx/LbNteFf+kmU+9e09UTmdk9pdGo8QUmNJKlWx5bMJWbPJpqDHlZmj76rt
9q3O9SlrwdKrpZEbZlIhSZw3UBfeeu2rpfUf8mdNkBf5clceNm1UlXSM4bmvjXEJ
+Ktie9Qn6hg6QCj/ym90L+mFEfpFTHTOxVasZ5Q7NOiOYH0I8RJpvHhiFN6hsS23
WajMz1kQ65X4OrvZbgu3Bq06wqrqfXpHLVoEcwWqlUJtLiMnsxAuweHGYhcAU/+W
Y7qEbUlGNKhqs7AcZA2JEjGXPK/z2orr4a8NlBB90EJsZcb5PvienqRLMjErpa53
BaU9s0SSAB9kXYoELMq7P2+LUnjdFixuLzWljf7kdyjM6ZG/LYkMIUSeFdACf7E6
qDgCu+3eFnduQCadqopeECVnoyuyecgZmzFLCSSO/8ryNThCkqVELh/C2/2QCDDe
mVYkVTQjbxj/LEI42qIoXl7nL8GpveD43pOeLpazpB+v6ocBtEWmhycg9cnWzhpX
KjIiekJ5sgO6AYhreHiotvHUUB/IFiX5RBlO9BOhv0exBeWI8qbBdwz9wA9wnqag
Y/1u5CmcpJjkaJBSnOyYi0U48orwNfJ5qjTFodP89aCRIY59YconTAQAv0+casxL
lv3g1FgMOp/bUgEV2Qj2jDgxlIJDpk/b9aUqEq+l6eTM9TgRFXQw2HHpDpgUL9rL
BGVFHp9ITJ3qVv9RwGsNf1iClwkwaKQDqRQR21lrmiTA4Fp4DdNvx9BbbucsAHvj
bIaOd2wqZq0C2sJNsotwWmYckDHwjfuLdkWGVu4TG+3WyNz1tCOJRoeDnEYCsfO4
SYZ7Ha2j/en29bJ07ZQ7ZuEZuTvQfNXFyt+PWUb0t/zYuGK9J/4w+ipbFXc/OijK
q7JOwknIFoeHlfRCMDabx/s0Az78GHkbQsYV7cLNCNHksgruPgZmUGa8DhHJJH+f
lMDCXa2WB8dT8JKL9SXkdlgmUo+BoxzOJXsxA1V/75/OBpjVHfunxzrEIo4fz/V7
VYbCVQvZHsPvziybtO4RkHRSQPRoON14huPrV2lyTcVIqvoxit3kvnSAIWChKUAA
vrMYacgdt6FZp28xaLcRErg+BsW8kSvc9sLdWQcayO3yhOR8KqoR30UZOWsFwgSC
xqsEpGYLXPoix/6zGNpZDz2yUe7iTY978eQXUa5XPQrwi4emXbTfYH2kS+Zk+GKD
4Daus9D2R+mIZgl1f41AoGZwXzxhWl9elSx2iYftE793S9mFWfH86AZdYj+e6vle
jEgQEpANaR6jkpUae3M79Swc3hje4zO7+rFsuQfuyezem0rkqA5Os1+M9NsyWah2
LozWTpBc/NKOIS9QsW8v/CGqAY/ow5vBII0P5SjUamL7QoAA3U+hRZBb8iVoz4Pk
7wc5h6w0RUjUPZ5H12vaWJ63O9j8KeC3R0Dd231Xt3/eWrmm04qpzXWo9yS4eUNL
zUgsF7wmAiYX+w1kOxvgwNM6sID0gOic8eT4kwIvSlHcv4WzxeAOuQTYkvK7g48P
MixkEnCvxHhf0BLueidM1yxcgVPhGpo9PcyVO9zc1RM210tU2/K5NUI+D7dBkVDx
yiV7KDhg1fxMYldNDOmh4jamrmEr4IqTfYvn6E+rDtB2GF0vT8Zu4TQcvh2n3s1Y
bnVngo9RZyVO6DRFr1BsdSMKAg8/J0+rVqPQfPvCllbTLNBY9OUCZ6mjTGfGX1td
PNtS94Jy1mbl+KW14vHx8jGwEqzg9b6gLYGfSYGd3Lt71396HN+26fOVl/9AAW4q
WlpUSCvwgvcObEv7LJLe9FRl6AwGNn+irnJlg498OtdNq8jdYdwKnt1W2ku/2hWr
UNoLpo5yGD1TuT4rEsvcR5+IjcteZ7ekboC3ef5g3UWMDDpIUFIKlI+4JS1GqHiA
/0acgo5EPnKfxytJOaSVGivgWPyM0ZbszteTOQrIkq4pFyhoXdIUzUonUqShNSKz
4Ed7v/3NJc4Wbz8T5bci+fmKFyM4vTCNd0d5IyM1rlSZR2196bDJL8kHpXVDET50
vi8IErCIQW3kBzlQ4oBIm13bUQ9jbxJvkbVwIIN9DMAabeOPsAP1wvH4NFbO8yjt
GZUtYE69g02vaMa4mfrOSWKd0GEJzocioiFBXNwiDSE4pnUVF7UglV4u/Dso7zjg
aOXuSwJOuo+mxGsJndByvkkBEmc6WgblCzKyfK2F/kV4/5G/7kFvE7EqZ6Cy3icC
WId1Wj5ib63OWWgvsSwDMDhBhYiOqdm60aU3KbIzTV30pQdyRRkRc8TiOG9+CCIV
aL0DZkEhMdNCmSbFYbYd0WejIlpnk0DvvpeBoIPBuk7fkB7kOsmikVKa35ffAxkQ
rGMKhm/M5a+/+SWkljQN6ylKHE2y+y+OT6YJ2sQMYS2QmQmthIrCZ/7gHDG6anck
k1gpMz9F5dSk06sVAaAcoaMGzQtS5w0G6PB9/11iq7mVZKEHxwPKiHLvFjj8dQWa
il9ykuvAS+k4mLMfD4HaLEqeW5XV7T0T1Hhp3fXUs793cVs9MP2wOxcQC8MYm/aR
S21ji2J85TZ/y38+XDqVtj6zQLeX6NebGWLe04qQRPzM1pRXclJIbKXWR4HXPkfa
9l314GlguQz+2PbUzLMT96VQAcp9lNsR+j4ogu/0yibDDlvH331n96BYrZU/7sAm
XeN1exWE9Jo+bAMXxwEP8pJbV7GI69I4jwoOXyl2O8A8uD27hxGNr2gzu9I7T3AP
W6N6UpQFKGlhVtSUEvQl21/AN3Sd5vdeqSIu0ibm+ovc7sm4fii+n+FxdmOoltrr
z+X1oqVHHw072eHvVawKju7MPPvsJoTHNWmsMBRGzhEHiPWI7N4JRrPsOucLzXjo
C/8yk4IM+DlfJ45DXCIlUyln9hpmcGM2Aq0O39+MPgpvwH4beakt4SX/L3ZQmfnb
+8Fn4d9X1NiPrZubkwW6Z/R4pajHicp7myEaOChv/Nrv47tv2vA1/zDJRa768Xtw
6HrYf5K64OXILPwV5WPOkq7UemcORQkCDoHh/3L3ei2WpGxn59Oao3fupVsvg/4D
tmVrel1zUooCFO7T2Zq3svPl7bW8IONLaYM/bUKLZRghRoZJbyVfTZ36CIy9vjTz
j3gtyzbLMOSvOgyKJWG1QfQXQ7twnLod5VYqmYwHxwq47JlUPU5yLITUvhtL8s4x
h4NpJWMGRIqVmvH9Nhl3g8amSMbD47zCRRmNQ58mHsD63eT/s3RWpiMG695ZrEIk
m+SCozi+Nj7mO0EppGNQAXsuklHOV/UMoY6KrWUSMcv+J/d3DjcJScZJEsm+hcoI
sZfj9UmkLzyVb856qOVMh2Z8UzCZzPtVEdoOaQ5+RfxyCrlp6Z1oxJCXh1wxbnD1
jJV2de5xV5AywtzfhJfmd364tKMeLzJIGLO36bxW+7Zmx3s+oYHWXFSV5VoNJQbw
alX/W7w99e3BW1LNYB1m2nmb0B+No8+g3YVM9Mt+OK829jc14Xy9fhFWmvfxO8IJ
Ivd/hFre1Dza16egzt6MA0fcUOhUSHr2c4JohENgZd/Kb7snPmW/FAPwIy/h9ubA
80HkuQMv8zk5sfxPW21ItImsJEHALPFXtK+6jXLh6mA7rPc/wZdZZrcxBq7R8ZUL
q5R0FBnjDC6xzpWnjvIY5alVtR4jMacOFOiskxRw6yjjm5jYtJxXRc8ocj8RmFB5
fA5EnpTTaa+YF4hDHa8HY+L2rP1GL6dLKsybl9+QwlS7TOvY72mN6/9bB7uYonfz
E0ah1bez3XkRzk4hymC07HuLmtY4q9EcFozIuOMb7z/I19QBAE6ETfieH2yHwevm
Y/+I2FP+ylccwr63jJcybdFyXnVGI/hecYjP/9kz0f7UpTINXsvlnmSvrOX8Iqen
WWes5odFCnztJ09f5bcOB1V3EqSfYEZ0+SiFdyvUZqGPBzURYyuLO/g9IDv2xWyE
1aR4EdTnk3kozmjdrABXfh4rLnMI4kE7uuxF2noD8O1MSD9QdGpdsQiLU9b/aAKZ
7pSHvZ58IJhcZFabpHXUBLrgOPSYhmciHuthn3/WAsdQjwvxmkFSZgVscVZe27C2
CUT7fHS6nHBYdV/l51fiTDluJYPRcXFvTKdb685KPdW/+1mkobv7zcnpotUuc6Fe
mAwXJCAluZfEePhJh9G+MsYclHXhBFeHZX6rimEZ8a8Tet3EP/QIvAMeSo8LqRXf
bKwq1suNIc8bXX+HqSXmIjqt2dsOfSWuwMD22WS6/VkckAW5Ma7C2uGYnaUGsgIf
LGu/DZtwwqotKxLc74YmrobQpUNoI28byCeOP22XX2dVRizzkCKEC2iEgyOLCeO+
3++4GAI3dS9wsEbnmjgxAM/qrrrKB1D6Gdt1VLE7shkq5rULkpsNxopZXnv284u2
BICz6uR56ll0C7oDQGjONUgu1qcJpcXS126UQ2I8XKTDDlnf4p+13oYvE03asbBc
Nh+oyzXRTYOzOMBP0CEts88VEfq2QzBulRHYT4YIk8ItsN27HJg8Y+fRxis6P401
lWDdXlQP9+I9DgnQ4Fr2Mn7o3UfVw+vURbLdrDhpKAO/4gfE0gNc60QfDKxeM0MF
QcJZc83p0K8NfzmMHSiHLVbasG3eFcD/4eF2CmKkfoApPVesY7Gw2pWxwBJCncVf
rgfOT800G0n2ChPDSX1bZbigjrYCWso2e6o9/S4iIap/4oWlq8MbPYBgQKX3/XPJ
mGroxXd1+l6kYq+J5+zoHeSH42wRgy+9zd7OzKcz4gR00hVALB+6AoRAL8xgUahl
Ya7odIl/iBDwNSfOYABG+R4ZBsnxZoHPH2UeHCv31WO8eMsYiOZCr7OXRsvqyHkZ
2q2age/RwhzgjomESZAKEBvTK28zsJdg6f4LOB1oeYSrWSEHEtghGDwJiV2+PxQg
CbTruVOn3Zm01uiFh46ehaY+lchCVwbDTxtIUFVBYt+9xyq/Pq8pd8pbZ/0rJxFt
+Vu69nf0fCnLTKaGtRw6bjx5RT5Hy62EnKmcTG+nR23dW9FpUxwbfVW8eWp3c9tK
FoapwTKkBys4Hy5+7CH7LuwkaHEA9esjHdPvmFYlOVyQhgrkywqDZgh95LeGZHST
oAxC6G222541/+5nPmFQaAPD3lCVKOMzSsEz7tF27bsIdYYxcIXorjyvSUo9jek7
Zkcj+4xVknt18iE4WQS+Yx+rMb+OglOZVm4TBQNF6i/5lYO3Z8soPGXhfkYD6YAf
jOIl74rkTOXGfw7824qMNH+leutylfedU2sz+J4OJF098MHHNPGc3koIozNuFP7J
3fvc9b1luP0sTRgXWbLJOjkAljUB4gTrPt75Gcwv87930wPzYmRn0sXCfYDhxJl2
CANtRl6DMgoDzL608LtVe2cmiv7m/3mPBiOdQvlNHz4kqjzlN9kQmKyjcu9OHGUe
XKGrnqxwK/HeO6VwXWD1DOW0la15OEgNk1PIlCeMfMrWURI4inQCYMLUdWxXJHcR
DXvXU+vwxOZn93l3B4MZ3lYnn4+2q9qE6mk1bZDg3y0P2zD7AmWB9zn3gmRlvbMJ
ysrPnm8++MPjzJK8W2CUS/WFddfXDOfZILqOWPfBUYIWNdfkBkYqb/MWMUVuoY0F
WHI+P36DvoqQe6qQGrPCdpJBz32u2oIKaUgeHFneOkrjdxPJo+pCG5sdn0K+sYMD
3il5Pa/1zyKFcDOPp330GMICncV3DxQi4B1o3pJaIzOp7OfK7wd9qj9R+3DpeoYA
gKIJw/Xlp8PK8olBNhJ7j4I2C4CyWWTSzeTfasgbrJM55ByRSFwnKYds6kpSemZS
yWWdFN+pufonLPDStFUKzdl5F96Om9smQyWoPzRm11JGQgtXAYodHus2bU9lmfHZ
m7inQqwwZKCahospKSd8hOu9OyXt2rqOyWiM6C+G9wBTuj+3K/3dWJxU0mRjtC+D
NCik5efZU3eaZ8nAiIOfOEmtCcP3rEJsPB58s/VwSlruG0KrfklB+os6eIbVYaI2
R4ubRQ0NHS7YX8dKy79hEKTT34akqlVg1Miz08oIAJlXEjFmYQttun6gPX0hYzBH
s3oHhhfArno4RF/qk4b+f8Kt9CRRfbXsgILXpyUPvQwScoaCEgfA/WLYAQJVmE0I
EZN65X6cxVLnxsG0h5GXiFwU4L0bHAm43sI3RnxbcBrh4CAYBfwC+vYNhc82rlM7
PCqNAWxOoVN6IItjtR8Hl9RPLg4EetPecpJ7tMi4JeRK8GoOJCEPTZcAwOP148B8
gaw0gL3M3VmmLlTv7ZVIhPfgwfaBSnRUfXWhfpk6M21/dlLA5k/w/8plAzIoFD6C
UTlDT8WR+fIkbGe2k2347MtU9gr6/N+uo4bHGVTnzyx4/6bUS/JLmKytBE+ZbkDq
dJsTfmIbimuRrupnfHvjiGX9NMcm54diWHjGCV/mUljC1czKYshL85RnSY/jTDQm
o5fhLI3aALIDanpguZ4zBIQ+SIhCaNfoPr5FJJgxgr4kEP9ARN2huZR4RXIJjX6z
x7hMTQpYCr4GU0yRbPTOKS3HS8DcoBoE2TyYoOpZ40L/pWlAm6iaxbn/qY01Z9Ju
e/ucYHzy7y17gfHn75sdCU2SD3VwkDkLl5g6ZusySSNsNKbHZnzZ2C2PRmNXpwZX
PwpE4Ydltw0HI1ZTkFBRwad76zB3MJOIi6Sxehc0lWm4O90jvIpO8prJte5vB1xa
QjFqLzPnd9vawbgfxS1b2yUzcTXtNOruhpXSg/gQMIGPU1XktgrRiz0ncrdohFeK
utcZuWJbDQjXfA6o72zNwiFiXmpYgp2/4uVMSnHFQJ2ZGnQqLnlmRfMVL3f/067r
7nirF3Fj4F/MMFnUc94ls6ia/5yuJggrkVmMu4ma2BBaQ/TSQaeWSM3PNpVCKaQs
Eqn7Qa4MiQ44q3p/YkKv+N3be4+FGDLvx7ygvMGXiLcgrFVVw3bZzj822jC0S9fM
c6XnwU+JNOgZDx5nkHxo/gnAITXXa3qHvbCG5WpwNadRXx2FDAXhRajEl4jLCosV
KMeFnpH/wCJ/G0E7RrA01zS352xc7xFGtehnmyIS+8+nWhd8BjXdxIyKkjamaMAg
kUteTGM6zsoIWMjFz0C472mhqW4LKB6aSMPjjAsx5sT2GWJUBC5m9L/JqZDGAlMl
40nnw9PMW9igtFCEVk0UqbFJUFwJuNhzarvErPdhOql5S+GriY4sDaMbqNv5VI2v
Ji0xS5aLUU7p4ROiQxyS1q1R9g+El/hdbuJI+CCIw6hM98L5XK9g12QwYLDNkZ3K
+aqkJzgkU0d8bmyNur6McSgl/B++QCE7xpOxfnK1zYxUy8Yoj0eos1Y2EfuNyVtO
RdYksGOyklvywdKbQnwl/I+iSS45ehZ6+HdjP5OhmqCuStiP51DDD5Qq9pDZqQy2
xtZ8tmdCjSZJDcYiJeFxMk8rIbwtWa8qsNC7wF8yXaIfNGF1nOE2cJyZK+S7tX6o
IJ+4URyn3KIQn6RO1LCmRetfh1is6OiwaA1oD/9MmYdyalsZqgTbKByPCb44PPhC
nTCIG4yHjxTGLJxFNB51/HP7GwncURjqbYE5CHbVZWnjNmr/tUGzvDh3fxbhUlpY
H8xNVXTBYKCiYVZU4bUHwRA5NAs/A6wNUgtPc/OBQpBZulUz1WDVfDVLBfMpOOdA
sm/uznvlGT75mDWCNttOek5kMViFXzxIrwKYuDF/17TIyrnfky7KQYSqh4eKHi5S
aArL98gMOBEc8dCu8RnoG2rDL+es4xNeVuWj1i9wQIAXhwoguufwd5PJboyDNyBJ
QJ8LIEaiglZ4O6RUEc0UOyS1w50QWxotZ7xcLAqAhUSFj4aHCl9VRGGItNvq77pq
mhqB9vP2ak51Dl3/re6I5aNIMqkV0/FHrOALT1XFmfxdv+YZyTpLpK8vUZxZj0L7
osVKzV3AKuCNGAxDtTbLWv4XiB9va9XZHBrSKinmidmfJNIrPVRyUdaqQlV0Ll+G
qTFFwzAaBp9kqy7gyxgN8+8GSPfXTm+PZCBMJ3NOoZge0oGLvjF1ovEX3lK7biQl
Gt+U+EgIDIQYaWTiL4oo3cEdcvyU69HdB1703jPEBbnoH/t8eU89SpclY3MDjTEv
JxDAqJeg0CWc/sXf64a06dwhm2PDPtbDUbjZ1Rz1MMm+0vjLTGViFWrcI2nslIPO
6jFQT9c/sJa1Jn8NQCfRU2PaFWlYhzs7XUkimATQsheeilrV1E9VI1XaNdlPaLNN
uB49/vAjQmDcSiVhoMn858YUnlAMui7wvFzMe1dxs+r/WLXSzuvrYPmVix0494yC
EjCdFlrdrO9mRyVxkX26I7AwWCuAULBcqL4n6SAKs93lbyTH8QprhXURomIJF+5s
DfiULqABzRET8OOAGb/zHMUAF+9cdDBIptRWs4dCVD4ZOdLU65nneEoYCuzGcVV/
fKn7zJ77vI00StITc6AZOYIUAio7vEWpIPUG1k0UUHsvDWj8ApV5BHFoR7+EBMlf
f3+tlT4Vs7kcaXP2Dy3hpeXFuGbzOC7LP3zZk/1xsf+e3UKBa+XMC5QSULTrnq6Z
9NVGImgutGvPcbK6SLTAWUborLF/rJHXOdOL85iheHLWfASr771jQ15qlDMLpH7S
rp6MdmFQ9kBm15VPXrv9Ec1WmCVjRxdIOl2N5oGMKfI0+6cFS7yLwT2QQusBH9fy
ygwoly/lfr8gWBAhfiFMl3BEX1Zxspp64lrR6Q6NLlZYAZOxnbB8QcHTMRLAWgTk
VeDPN/rgHnUwWm1NopNeMjdxkPhHHfH2TI6wFlbBnnEjOHetfiKsY3BJcx++itgQ
OSPfngUL8j7PHf3d+liFqoOvS4N4VK9CCpzgUroiB50Coj0AY3IuPjllzMi+DdN3
H1UpfGzm6fcGQ4MLYVMg37i404uSh9s40GnQOTMLO3DJx2DAurMOevQWMfDH9fOe
FgW9xzneRMNkOlnuislIKx8JEaugixnLLWbEGQ4iUT3ZB+podEwYEhLOSJfHMbpA
tw1bTdr0vaVeTMSiBDAJ2/2kfAkO42Oj6oGjqS7Cr65aF8WjnxgZkGaeRGUwkWc8
j39yxG37nlcBhBDEnRRSqORuuKXZolt/j4rbg+/ILVGoyZVMoa1hh9jJSpKLyG+r
5EdZ2XVyvJNSAfiZsA25nTyp2c3983EwW7BEb89qRaaVNp2DQiAq9cDfqBgmh3qe
wHFUzp+4Vficl2znzaOSPmUMnc7oKVgzxLfQAJ/cBkDJD59NDqd84YERMzq1uqwH
Y0qTd7cltxNFkQtMVgxrzVR1VijO02iys+XjvWFcBB4n3AdUonJgzP3lmVC07N4q
1qFrzeYIj+V3BVojxYVDviWjIdLwLAdqc7EXJ7g7E0c0z0NA/SnmeAvTgFsQSjHT
3FyV1oghVPI7F7Hku/bl+IgsdqZSmmPnzlF9uhKTvoCmJq5FqQMdDpQqgMkI1j5R
zoKvlxTMPzN12idCS23cq2CrIfrQsGYgHN5STL3VIkstUua91emobRw8D85jl7l9
Ibqwg+QlYfu7k0oArKreJ+HkbwMPnO+4OWXuvuM6x6t6W1GQCXTlZi2ycbu8WZOH
qZtXXMILkU47U2QlA4JTBzoniI6b4fvPct+3JTFUO/TCZSTrPcpxLwGUVt/5k5b7
/6HyytyhQVBEOYkD6epmubDzv0q8AtRN9ntkTiH3Xl0A5IU15WZ2kJtGu1ZmcpYD
60KKOmTw8tD9as3lnwaiIAehhoY9aLrgClF0Rvtbig+uOgPzsd5g7XS71kNEZFVS
GNZXtuXcnRfaQuNaphqNcpM4S6aLk2PIwTAX7PN9sztDMRz424z7j7L/u4XC1tWV
6x2R6kwhO3NBOT4GDSSlDP+z35n94lNhzi9lwBdnfx0kn4DnrVsw5lo1MvvM4RT9
2ZRVoRXeb0NxWARX2UxB0Oa28BoB/UxwygekQ86pMH5lzEBPjnJsnmxETxrbx+eS
wyrjPINBoxN3KQROjm7zr+EZCbteNsg5g/JCoqipask2osuOqwymLylZrFXIlWR/
oqBJUnCzTwQxDervgqeJFzrSTudjWUyCvObLkkGX9iIZgu8I0ywoWL/Wv35mx5+i
pTFJ9fqWEuO+tF62huAUur1P9FYOn+v4N+PaBJqNin2J3i8FcV6HH/wCRi2dX/gT
Fl6U3oayH2ErJ3vfimmDXrM5PuBpbnsZAPD1NjJYx2ThcdjcPaokmg9AnrAA3pin
Qo1GfV/qIHCWZoAxdFI1i9+q4zwCRO66UKS8lu3WJSqurg6DphQzITB4fwHHBGvo
qXHJ1kyzuxo8A/myIfVXCZjHwrXhw3BFGxkSDL32Y+3B8BIj/tTIDmTxlsUQlp3g
LdrjinSLm9PHAJVD0nd2Z0sUKSXlus9jCowuxwtphDkIGfmLV4X0W3RgrRdeF5hn
Y9uFC8s9tnl5on5S2ypt+N0NDm90IRhayOROnV3IrZjDxk9hxl1AE/TUEih8V9B8
oLv/ZEcansRL7m8oHb3iHnFrgFGuXh53M55k6pFsJj4w7bXRH+OlvI4TTNnZOgrX
4vMmKAx8+AGV9tclQEHg/toVFzeTSJth5p+DTAPugtSN1UDf1rmNjycU1c3XxsXl
ktHEufWnPc79EKI5jkz5fETmU2DH1pEm5eAnLiZ0LvOGS9ypNXGRsrrgYcbtvRSS
DI1U9OweYINtQ1s4NulZw86J0gjmMXAP0/ZJhr7fvYdIzTZS3usitoi76bQ6XFrQ
sRhLKrREvxKr/YmnuF5T7yR824CFemNpb4iURfOnXQrrv0evtNoA901CqriTB9Hk
/JXxT+vG/xJ/02grA2if3qM7o+2HyALY+B9DWswuef5D1IYZXNY91GGo2IZmdcjp
zgojsAoki0nBQ6hT8+WSV7IDtviswlL9VefznzpxnyRFND6FzEXFI+sZbHjvcLoW
AgR4SlnGIE1JkEWrwH59ZgD1Yo9cKmEI8SQBvZdIB2jjRmEwABSZ/8P/32ZKkAF5
DGe21Co7jwIknXjoo9h8FopZ5DoL5kXgLwuvptARk0pCv3HWvIM7BB+pUrV0oIGY
GCVhxVpfhr11RiViASI18uaztOvZB99rTonRhAv2etnX93H2kA8POZhlXBMJTP2P
CPUanHuXa6B5L86Sgx4G0mIzYnToF+fjsrEZCF+6sZzCLiOIpSV42GEnXa0Tpqbi
MPY//Z+19X+j1bYPniUG8j1sv0jPU1lQPwP/aSe2ZcdM8dP9A3Nyut8PymV23ItS
xFrVTWB4UgJjaNRNOCsXG5ciuZ1Rv2egUrjCc2R+NAHBQIXBBWA+/6Rcu73OvQqE
l5/YI3aezxL3xT1XucICcy/s9ioGjcO6hsu07711dDqKkNVt+U0Sq9Inctr76vNx
HIf7jyzsTtNQFmANsfrmRNewnvfs6tYg34hFNk9vrzSnzUvN9rNrEg35QKgUHLub
TlK35CB+QOKtq02gcqe/yJL83tg10gKjFWb/f6kJuvGr6+h8A2pnedfPRE2uUhkA
6g9lKXeM6VwTQiU+HUQSWyGXE9lBUqwUzn0ysdEBkqRlRhTDxIZDZIDDFmS/UqXh
c8mUMxPz1+hR/yERz7/x6UwYGd602i4Dhguw+WfDt6ves6GBmHl5BwuqviZFnL/2
2jvaEqIuEvGyCbaYGhkqWyUjdqKAS5qVPNq+BRT5nMj1Y7p1zTDg1jSOPNSC5AlF
q+9gFR6P5qtRzN1Hy1DHdki+EdyUbD+8w1u0qX73OcsKP15OsaruegiYvnTZ73ki
Av4HD6uLTpjTbwCT3FC9QpTCM4jbu0fiwrKSQfaBol5FFp/0abTXS2E9j5Ast57A
Emwkg6GLkhnqaHWT5+5wC1SVa3g/J21sBWiVA9WCA3HSFukmDq7tV98OYWlR3++n
qxxvyHOim9Jb1V5ar3mZ/aGBW0DcYHro5cfTL1+k3o1OUFvIBmnMdlqPTiRkG68W
fNrj2sREa3e2pz37vdKwsQLF2HnuPg1jUoqomA5Yj3KegKwQ9i1wpDSz2Ky/k+qC
EcJdg+iA/EIQC3FfCOklzlXorrWUgVptpnyJy6ffDxNeq/RAAfverR4nB8YBEyyo
cfOsJJ0AvI/xzKSd2knHsCEKHj1l8TRwKCDhPj0yQx+yKSSXp3i6zXV6SXBVH32g
gEHFVgVtNVZoUOUEXQgftjXWNB5LEKos9MJnWX88eXviTnuHQnCHRXITaLRbmPHu
mSGUH51M56c410ELDws/jCkyyORU/V+IDqVoxBQ/6/4+sZ7SRH6E+f5bO7qPWMDj
cw6d/YB9e1FlYdHrpjr8kQohcTGGHprDDvudyrbVnrZehkq0zHwehFz0eh0U3m1l
aaG/PCzsjTn/BS4adBHLMkNoDsQOYf2OlHfKsJ+NoEuG9eA/+JDDgyXaWSj2VWwL
m3oE768nNSlEYxj2Z3eCCaSSOtL98kFfkQYiP4hQ/MwXMi2LUk83Qmbo12SPqcBh
z+NEXsKU0Fbapd5zZoaq1kpCtuIIkF41AVGquZNPOr349MrXJeyVqAKUdHEEH/ZT
mfe+b7lTyzCEpGKYjacQVOxIJbKBIdTxILiAmbIAVtVf91GFtC7RiUW/UslTEtH1
ea2Zb9F5SPKpJsz3moy889O84NHVspNdxmK+jTbq9Duz5dVkEhGHLZrtwuptOwqi
9iUpS7SZYTnQQ9nxOLBQFWt+3Gpu5e1on72KUimssN4XyPZ5iTcVzMLCpBY+Zcsf
OFYwn57ujgdLfYq9ZdE0gqfVOvPKbX7zREjRdVbDcjAbkHbmljT/cgNI1rNayeGs
u4pSbs1Os7s76twnrnt0m9Uuy37tf8uJAHBF4WfxHmt69fcPKa3KNzQU52XJ35uV
M+fyaw6xxFaTHdtgf0y0vdHQInHvOdrtBRDl19DEsjPKUbvqUBUo1f8cxe/wCMgH
mOqCOIXSGm2hvBKSQuJP6fFIMuI+InbhLbu4h0VYxHwWeVwX1mGJwdWPhdwmleCc
yNAMD/gomQo/KNHdLtukL2LauFMfhRq5fzPMJl2gxv79y3JI/Q3U4mM6vJPLKR1j
zw8QP842wZLkHgTzVQdNiV1f7QLhs9jPAL92LnYeRnTOG6i/XA2wm7Cptsbof0uJ
r6mTgd81o+8QMNKU5PQKp5Kk195JZLGGHdlsy3h0DcPHH7RYRkonGnkvwxoiNyt3
03l/GlDtN8ixZBG5ApZADhe4rmOh3Jnb8j3Uc+eG2kBDTnXK8C0s4YIFGqooZj1w
4wMkYIB6hhjIZcbmUUQTeYEHUjuUIalkKz70VNMnEIqyVd563uE5qFKkn8M4kWBM
g/KLnt2bKudACMlW2Z3XS7vpZcuR6e+iuDWgaM4ETvPlVO2dthcmpChrom7faDM0
rMtTA71zA7cDjUIUetks1GNgjB0n+k9GZoyog/MqjagsalyBy2JYaCFrz+l8kRXc
OeLlzKT+fJFiM88VWHEoWIIMnIvopcfARZnDCUjVrIn8Ofjno3Mq9YsFOFCvsNUk
j3sqR54Bgl32xkaJ2+mvDByWywqwO53QDZCnxMispbysdZXJgAPYLviVAa+ehtII
N2l1pxzt0Wez95stUah+UQFMDS8p6unbc6Wed8/TJ12NQQl6WBltmRwaDh7dIA0b
ILhYOeNK5NQWsmt0Eit5MZc6clmuOtYr9fHe8tMfWpHqZXJiHrfvnFm1S3pHu6MM
VhHqd9c8sk38qLUJFfUjwOnhyjVZ3DXiaF+hyJ1n8vNEi/MCLNANqAUZNf4RXJhs
i2DNYMLDsvshE2xFN5zW9EyFCbMYjmcTkavfLIBfJDKGb4CoctTpUhTUcvGEm+I1
5dTzUwbZbMkFd/Q2ZU96wcY/XdtAV0smQklyGFK1YzENZTaXrEIL2rgXdBKz1aKA
0ny5n+onGKdkjG77E0swIdzdWejA5oqxLQzAUJiVSTj0kGqJ9yWPAcme9cnfUtd5
OHaWhriZMHg7GfGxAjIjpY+3FVMM3BPMxf45MRklTOm37CmSkcGG/iiy7S0z+TYA
J+2p0zHemfL4oZ0Yhq/wrdDd8aBVgwvrRmLp0COXFmsTCkUaYQbmrW0vO2DdcQrD
uqXir0/EG4UAp16wAu80XqE1Nzhvy4GMpZGaXe6JKyv4JxeJQVEUPbhjZnbFx5Wh
223YF10XNUSOT5ZRLcYQfuRzEFmtcsGtZVt574pEmd1q2Er0Ksq9wttGA7gXn5Hx
faYpLrl7EEZ2Ys7Pozzu8OjQI/LsAOwZ1uM8fEoQeGn8vMeBMe7IU3GB9D8d1BIf
0LmG810yWcto+MNowqGdf64z8nLJMz7Y3n0XCsSBftXHbSnD+9o6t9binnggFwe5
YyVxnPpEOg8T6eGYV5Ia/hs/IbSItsyX3zY/Zh/khG1Bri1ZwNYWm3CFogXcH2t9
lNPJZAO1ikv6pOsG361ALzuxkr098jUa+05+8f2kBrv+/2XHxW7sej3aChjelxsP
QySiYkXCvkleULZeZgk1QU76uIz4d2jwXKtoig179FEkVHmo5Wf8qi4B7JD3L4nk
LLqb4G1dLpv6itpB84StzBcJjy1235q/bYrm8fu5ApuIW6lI6zxhfjRdUYeEvUyq
qowIZJZIHEqRV3mPzHjgGQrKXGr9AbuKk8F3cMShlQMovVkF544yyS2hBYRAtnQS
GU1qK/IEB6PlBhQkz5xhHBfzzfz7FWQaD+lCE0DL5+mjd28eHCXGAN58/cdhlPxd
J9+d4I5EdXoFmZs1wXQKSJecROOidtWIGmS9/2gZ7+eMK1x2PvHSdaNiN50E4uD4
GEwjfewy5jyJNcLNKULHJgARLscyAmz8cU+eESZFKUbI6x0A7+g8AzpjVJFoCgoY
/Nc+KwTqpssBVO9lMMGxpU7ngzh1sKFw0uR8bzVCbtBF/Qsn5KXwgdxzvGBXubT5
JQqCeN3RK/XkPj1q+tqB1hGaStRYopyyWkq/cadCSBOd9ZXE8A/kXwTnKAMWC8bV
xHrDuGgIXw4KNhgYhd6hOxGBazTkXQpMlRqvYXtrY/L41mg9TMzF1oX9mT0FSTca
LwPOwFnvKHWAN9AKFdWLmdnOE/gRbKsZKhcPP3WBQmyFTt1z3JRJXIanYpbNOBq4
LI+s9DxT+hunkKS1BAMWphf2tAcHGBKd5Mn4pJ6zYsDfImE/nWFuermhejtCj/li
tJa033gAja77CHMKFaXJS6bGvZjVWnkYjvFxvNWVEVTChSTcXvq/+WhgOAMTvfMO
RFrK0acCPSWNpQrr2P44VjYDvEal6y1Gx1ZzSWrIcbkJV84+mqSNYg/oieT6+9JH
0Fes66mYVHRSgq/utWnNezBlMq+139untcdrfhkRwez8Xl/ZIoEkvLJRiMgnrwwk
KQ7UqgrEND6XfQ12eHWbJt8jAUNqBAo2ky9JHJ4urA/4B4yVjpBkOPc/B5YcypxC
eov7l6hXCjMLAa/JwZe+7k0QoNj3upn//o2Z64mHg1O+srt3rzyih22EY0GB7Z2O
93fUZZlG7EpiQ5vw4AtLariXSnut0JRidhNOHNBuH6WTnX7vUjjUsaLtck8sSitK
PcknWwEoi3E9XzR7vVlVHyeIuC3PAdEoPZnafLbp00c8l5HtqWTLHjopszr+tWGv
/8ongOutcVfYXyw1JNYBdhQKu2gcuhmznfx88QPTyUoWraYVFyG+R8UvsKdxbw+u
e+MZKyIVyL8qJAq7SshNf8m18BoZTyYPnQ099fHJgHHQk5NsHQ4p/BO22FsxYSpq
5/v7Tjoz9sMvF22pu5bW/B8gErJID413CXSSP6bDXFgIRGaSqVM/vpJyXDXCg8da
yaGGef1/E7pO54iudiy5TisiO+mY/P2fL/WhOVSF1yP6BljMBF7zcIeWAHrQBBha
YP+6jBtmFfYJjZ3B467QI+KAQJ06Kk1R1YfXhhHayxXce35eThas9XPc8S9x5K5K
hN6NLDZVJt/W6eO0P7w3acFQCI3wYgfIQwz5aQ+ZIkbIMlKtZ4UhzuoCkN9AGRs/
YPF4zCjYolQKjkpDDi3uayYE0TdeaOfAur8a9gPMoWGBJSg5CaYgXWWr6sUwS0zT
osIDrJK6j7TFRXyDXESNcq+YWgnfMbh7ACOSZ6iuH9VIsO1s/YHxpkKukx5JHad+
vpQhngfOhEphk+iEmiLdTEbuPjoIfrn3ab8Bf24wIJU7ZfuGLLVETWDt/VFDB9CV
NhopyQQI4o8Dt3NNja0+PfyFHhLmQfO76lZgyWLdv6vGx2wgqZW+tOZnk/rUXFH1
4Si3OwIbENPD+GYTH4cU2sfk1OUNVtl+FlKhmu502eJgITvhJWlq6OrcP1MPniYD
ddFKNJaZ+rMHawP2mgTILL8g1UdBplzHb6uL2wGqQH8o3FaQJ4y7rF7mowkeSAKV
3VRC2Owheqr3TOioCuChHwlp4e44hjCvLrX7v1g6JjEoEuXTojw00rJ0pOIeHgK1
Y1DBWPrihjrlt83j3T4VYn6GFIXFVN4sTSGymIQLGGSkt4SehcPuS34ccSfwb5AN
9ocUYV8SD6+nkiPqSWhaZbyMczGkY5blfasOjAOzTJe32rM/tO/4Ok6pPSYg6p+1
PmKRaZHnwI2LprBtBE3NTFATtzqZPayw/YPul2fosnQd49zJcGL5mTX3rkhSnMQL
kO0GZLWiEh8Aqfxj522SpskDUyaq6QhrIMlibKuLw7RhYtpLE/kAN/igiuBWDfdj
R1nj94m1agphN4HxbpR/yqd1ii4cCtq7ZC683M3CjUAS2R6odoCJFyJ0ehqsAH1o
kLmCZDefTYeLPpls0Kcw2benikCFLTA89z24uG4rG/xfqYM5hlAeZRzVFaBF/z6W
i7VtuvmsWzB9SXXlI/Oo28LZ6mtcLfmNlAG1pdWqmMTWp79P8t3mtrp3nOGqECH9
hygsQ82UtY6+MnpeY8gc1WIKdjsRwfTjpHI91zaZDO9hc5GufjVkVLHjMX7Am+RX
hJPU5QJTrZ4rSnwic3XcN5hXv9rw+i0tzTIRFWegq4ugJcbKpKkTkRugyFuP5TlG
6tF/M8wPhGC1aXGbpuCcdC7bOjfgBv8SbglDoumlSGmQyyFZUS2f5YbJ7Dfvw40o
b6ltE0ioXToyT8K12Ft6jqpZo565HUTOtR8htNXg/6a06HAsa/JW4HJ4fPODXdGD
3TXcP8kxXsMV7MQRO6vR2qBw9hEHWxEZ8wgBkv0oUvQ1GnTbYJY8259nDfiaygLP
RJLBLYR10BHzowvKEGQES2aAPfwVwurpfeZ9qHOcMXHOrEmdBIWAmwlDJeTXaIsl
MmCCx2+ws1DuDkiWbTYRLOLZHOw6TB7NqOGBqrDNh0SgRmg7jqdjr8ybEvs0Z3r8
0urZ5NCt4UVT6LuoK/eWhAvuxjVwgoPQYUq6BZc3pDRGnFGMgbL0WgCvLqNwYn57
6QetAFNi9QdbdYGr0VAsuM4ZMfP2EiCXpOR48U4m7bhOBA8gRMS7FmUWXe5KDsUk
1c2XNUoi4JWeYwixfWn3jpIuImyWyzwxJgcloz8hP23Arw0ZZ/Gei6OCqKxAU4Ef
IZnGecd0vMvJp0/upgbcVheBPOJExfqLUmGGbYRYiXgmHJYsa8E7EqYtgqn/hcYz
kVtyp4tzos/OJyWlfCMSs7k3ZyyV0UTmTKe3gSd6S7kIoNf+10ghLYgYJHNxr/30
GKssJxGWqTBvI6dRX20lwlNtHg/+IsIsFAmbk483XLxaJmxfzZDsDe3Ib4DzOSBz
Zo81zM0vfjecV5JNdS57H0OIgqNdiMz9zkZL/sI60KnmV+78xizZap4zN3zPcFix
2VwFg6+QH+91PhNCwibIf+SKxmOrvswjUiXZOkpsPJPX0b5eVIW4X3m1krPMrgA8
86D9iiMJwvU/Ux9Umy5NZKjeabJv+pTE8h+fPgkMqvqfHdZVLrr0Rkn5/t6I+/1F
M9v08aSHa9l3hZW7lTylyyLGOtaa8FuBvtYCpiezR1rkjNyS1QqmhPjMt0lmpJlg
z3Y4mm3fkhQhI+2sQh+wo9MKRtH1q3xnuH0ywJpeZkN7nEYvZNxjskbtA5nLeeuy
Ev3wf5WrJUraErlXE4KHyP1BLeoF5tNkp/rqsK1U3HYM34Mm1DiJrZgjCDo4pEGr
9nmBheLH2aaShl9F49ZbL8Mey1ydkirT80iNfPNaONY7smaYlKyZrN/ll3weOGIT
oxIa8XlgyofriFfs9y8HXH8xb+3tenDf4DLCZqmT8Exb3Hhskf9pIrwYGUA998/R
nNxB+hOuQSIUgb0KXgu8REHtS2cC3Po/o5CARHNbqfVWJXyFekTm09hN/C93Y43N
SNvbQFq6roE8XWTs/0L8XnpAfzljLVZeUqvb+PWUiPBNKnpL7QAakz6A7jZFp2Tp
fDty1/TTnSYxabGVbZpODQTT2Stuk3JTPHwOxWRQJGoSsezdDJoGKtpngFwy25ow
LFLM9yGZRSlHlYsgZ/TIF4XI/7Lrq7i5dcloDQoEBS7xNIMKW7D0azt4JttVTktp
EicR+XxMufa0R5jn5jkexAtrH+xMYFCYllkYin0PCw3b6xm4DxghA0sTZq8BFahF
ECgBKFDuC5L5aVa6L654pCp5AkmnWjh29UxxQIQcWxb9Z0p7xw8yHxNZoezP0zMh
x5L8DNHyXLBrtORTljjrxjl5xiuAeh0yhfTYqqFi27aUrDOqKToI1VOzfNn2F+zD
CcqUzZo+1O/Cr/ygeuDuJtjMlc1vEdQ+f+zIO0D+D35eu7vtCnwLAya0zlPvY+42
LKYtwoSKI3GTegFw3/69udxFzYhiAoE+rTj/2Kpuh2EmXUZdY+WhYW/BOSKJ+1Nu
tCmVFpI3XjY8QTSLb42vso4v5E7Z6Q+gUfBqnsc9Zg0mHsn5gfeyCg7eSFF0SZGf
x6WdsAOE2dpCjXXkdKbgivbjRxokYkPI4yXPTDkdW+E/YavfXuRKV52kXyJ8XG5N
TJcT3Q8+ymikI2Yp93dPfoQEFdp8oXL8IHUTjCeqAd36Ue4m77zW3wF20VqRnC7A
KNLo8Ek00WNblblSCtRtpnXXx3qdJes4ygCudAnWJWkWmleWRvNB/mtZiM9hoJs+
TbFdgkfB6DDIPEvHVzCUe5421e8ecuafNdoLehzCfFHPj1be/EDGDgrb0ejy9tTL
WIh8Agiuz/kNXfe7oSbmdECUVy8EoxY3E0+cjvzRCwd1R5aHp57jmXFbOd5k/5So
25dpBMtYm6Fj+2Q7K5aT33IdbzxxQXrCRMDEqwbDNRvvwL+W+GUFAkTntraQgxyu
c3vvMFVeOynNJgfVKurSRhrv/OD//+k+qX1xFVHkHXd/g0cPwZQEj89X+qrBJ+Bs
hYyhMRKk/n15hVtZs4zFcNYfs73ql5TRPRdf1qdRbP/HXYEfgzzjoAWw+1Sv+OL5
0dtqjbB7RR8EKFz72AryvyC+RMaFa9zjNqTmt9UOrJHjOmX+YbPs4LcydQjX69z/
EsO0DRS+K6qMsM8mCdwTNkZwUbiKXf/kZk+DsrV6/lzfBQxyaMz08ybgjHt3uEs7
eVf8oD6490ckAeVrklPy4yukEVgEwrtswTYlN6gc9baLsqqwLd2ALQM6vacYJ56s
b7XplQa/TugcLb/vvHWk8lEmfqph5Y4PnjDR9zW7F3I5urp6ItGK5QuwQPGCr9gT
nSGlVNJYgfcbEvlgyrEJcx3wvB/pdfkzs04KvECh0eDlJtOXY6UETbRgeXeRQhl4
8x/8+XbC9ug9vlS4DjVZ15nZFqaLAEs8uwSQFW+TsCZK14+2wvlQ7CixNB6/oy98
Zq43Jld0GmgcWGRvzbtX5j9DaRF+zN8jL9P6ohyPFHXBo/ZUnYnSN9xeNtv+FXJl
leTng1EN1y82xLX+fWnd/g2+7Wredlvl9Iqr+F0hhT/TquWVoxPpK3xhBCB0pdt5
qOJaZ7RCUGbeQTRHJH9ZFCIWdyeEQfeDMx35HdK/85hAwn1DCVFjtT7tcgHjVtU5
01JCtnOxSYeLtzDIITPhs70Vq5YmWxXJYUGxHdYJiH+dcgDwR7f6Kq5j0XsKH+Sg
WxGCdXHItKAeHQSxqrKA26yOuxHjL461cOIT5S0tVdeZYLwDrtcbrstqQ+qGXb5H
gnghi1ex/cMIGBtgvhbHzB3SIWggalB1FLlEbfxvocME9ndXUUvSqSWPuL1QTcV7
LXEEDQUuDHgOQW3SSXJKpteajfGRQsUnKfNJUdeJVVufyBKy5KzSGCq/4T2bMJdG
ZGaxRc8WMjbdbiCaaJscnz4mboGistudMmsPQy3+YK5kd8gUohWZ0j4+KiN7z1g3
vt9XOJqatsCtWOuUiQgSSHqqVDPr6940DVfzVlmXp2wuMNaycqsGDWceeRTNNBY5
2NFuqCmE8NLLRc8qd2MsYodRoZilIdgIoBp48otKn7XgpXpWn78CcgUz0br0Q1M6
jOErGlx9gKNM7S1CV9DHtL2kwptbghbaOKv91Ln5dEuubQsNiEUbuWQzk96nheWI
hwZyNxzbWskCqOXXm+go69t9qyTU6IoE3anO5Peap0Y24ya5tCrYJIf7uEx0h7iq
5YWhVMMiRcR06Pfd1sxjwttvnagNCvuR6DJMD65k7+8mV+FOEVPi4FcNaeuSkit3
5yThk2v8Pgk9FD4S3m8GNN88RUODQyVgmklQFTsrAWncwi4vjnciNeAStegi9auA
ew2Sff3raAujFwjCN11ir0kdsnuW22KNDTFdtFlujcs7kbyFT2KZdKBgzIfdfIIk
p9Sohpmts+aCBoxu4Ki/oZurd0u/Tt/zLXnc/jY214t1tajSVF0jdG9pBFXiKXJs
BkvN2XTaLb7wDPQEklYB/ozyXVJ1dRPT09XFMgRxOaadhwccw+vcr1xU/ukLakTn
UTTb/rMogGzUUVzNO9P+04+pppDPJaKRHVhHtfqQQvZ5viisTCpWcpvUzHE3uPid
8tOfy8UY8B/Z6oQQP2EqjsiiPGaN8LFUe0SJKctqf6FIJbXPWB7VAA/BKJHeTQg9
xxTOop2A6Q8iK33jwZGZ2XGO88cFBIaX1H+o3HTG9FTAPPUKL4tynx2PjCGqJm9W
6h4gftEkWsuxGnXQdo5JWuCJ5UHNYVcuCk0R3z8aSrWy09/V+LqIy2C4Ae1b9BGT
lP2QZBT1e9UFqBhMwvM8Ouq5MAX58XP0fCeZ5LCayNTVNBk2dsZLaMTT49NWr9w+
E+prr+kSDzgSJdx2Hnw5U1kaaMfalQVT9sBx7LIs6L8UcFCu8m9+7kqpUhN+Va7p
Z750uHYKZXjrdEhYb+UG2aob++1CLGXp2akWb8E880inWp+UmqtTK9jlPluEegwG
nu+GKMnpFSkfWDCEJQXgci5IbOTG5TVH3qUmspZ+xc+3gxtd3w4rFzLxYGSM/FPx
eWPIIb6uDKx5WZoEv8QPTYI+/lSmPl2JgKTuh0pe4tDeKwY6sst3m7oVHEoTsaTN
8GO6ri/HeMqWs9yotgGaLIftChK9LbvBMgpK3QgvFSED3RghW1g8ah1yv5dfjBD5
FSzwTr9pSA9RxsV0guSazV4ROXp5Z/KHChBbz2Bfpo/IyMBccjOz758sWvvQuMYn
yH1DIkGzgnz7t8TJQdmgAn2TkFThYskISfy6+hQd4CeLZ1ycYyj6Ixjq1dXQtWTB
LMbhK9BAsNLjgdcTRz3T1oEx+wLylgNxhunCBmcJ/Pq9woT/nsmug+QLVsZ6g0Fb
wP91CoSk8iutuOebjPm5pvK9TYXRbHlehdSkTkgcBIW7WcBTi8PNrMsDYfuclXyU
QbTwNzxtY3y4NMU/dh3jp3LSu7kvyNxzh9Bf9aXE6D1GvXS1QsEnNV/GbXFsh9a3
RiSEflGvIbgV6k4vK3iza7/VauuMC0Xvs+H/zPK4217RFfUh8YmRSoQgGZ8aIlRC
N4888SXvPWTUar3FdOIPGYsfL+zP3Y8IQPGvqCEtHsuYcB06ehj5wdduSyZVLU4C
GHqfQE9HHJCiHu0SUr9eUIa8IJBB7sie4bFo25adOrktgCBBxxFpdDMARlegmDag
6pdubTk+wZynTx61W8kPiyYYcStmU04O+Lv6H9TujxIGkkVv6nd+9F7UQcq7++wx
3Y5nHWd30hvi9mCX+6AW8WHWwpXGZ+kn4IyGaLnpiQjgyyxWKO1ohrZ7WNNgMscP
lE3Yksjg0ouhYCpRx9R8MRIMVaC6O/32nad9WMH4NzyU9qZjkHhsG/YtVBn73qPG
8+QuQOpP2k83zHknMdLg3Q==
`pragma protect end_protected
