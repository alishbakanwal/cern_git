-- gx_std_x4.vhd

-- Generated using ACDS version 16.0 211

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity gx_std_x4 is
	port (
		pll_powerdown           : in  std_logic_vector(0 downto 0)  := (others => '0'); --           pll_powerdown.pll_powerdown
		tx_analogreset          : in  std_logic_vector(0 downto 0)  := (others => '0'); --          tx_analogreset.tx_analogreset
		tx_digitalreset         : in  std_logic_vector(0 downto 0)  := (others => '0'); --         tx_digitalreset.tx_digitalreset
		tx_serial_data          : out std_logic_vector(0 downto 0);                     --          tx_serial_data.tx_serial_data
		ext_pll_clk             : in  std_logic_vector(0 downto 0)  := (others => '0'); --             ext_pll_clk.ext_pll_clk
		rx_analogreset          : in  std_logic_vector(0 downto 0)  := (others => '0'); --          rx_analogreset.rx_analogreset
		rx_digitalreset         : in  std_logic_vector(0 downto 0)  := (others => '0'); --         rx_digitalreset.rx_digitalreset
		rx_cdr_refclk           : in  std_logic_vector(0 downto 0)  := (others => '0'); --           rx_cdr_refclk.rx_cdr_refclk
		rx_serial_data          : in  std_logic_vector(0 downto 0)  := (others => '0'); --          rx_serial_data.rx_serial_data
		rx_is_lockedtoref       : out std_logic_vector(0 downto 0);                     --       rx_is_lockedtoref.rx_is_lockedtoref
		rx_is_lockedtodata      : out std_logic_vector(0 downto 0);                     --      rx_is_lockedtodata.rx_is_lockedtodata
		rx_seriallpbken         : in  std_logic_vector(0 downto 0)  := (others => '0'); --         rx_seriallpbken.rx_seriallpbken
		tx_std_coreclkin        : in  std_logic_vector(0 downto 0)  := (others => '0'); --        tx_std_coreclkin.tx_std_coreclkin
		rx_std_coreclkin        : in  std_logic_vector(0 downto 0)  := (others => '0'); --        rx_std_coreclkin.rx_std_coreclkin
		tx_std_clkout           : out std_logic_vector(0 downto 0);                     --           tx_std_clkout.tx_std_clkout
		rx_std_clkout           : out std_logic_vector(0 downto 0);                     --           rx_std_clkout.rx_std_clkout
		tx_std_polinv           : in  std_logic_vector(0 downto 0)  := (others => '0'); --           tx_std_polinv.tx_std_polinv
		rx_std_polinv           : in  std_logic_vector(0 downto 0)  := (others => '0'); --           rx_std_polinv.rx_std_polinv
		tx_cal_busy             : out std_logic_vector(0 downto 0);                     --             tx_cal_busy.tx_cal_busy
		rx_cal_busy             : out std_logic_vector(0 downto 0);                     --             rx_cal_busy.rx_cal_busy
		reconfig_to_xcvr        : in  std_logic_vector(69 downto 0) := (others => '0'); --        reconfig_to_xcvr.reconfig_to_xcvr
		reconfig_from_xcvr      : out std_logic_vector(45 downto 0);                    --      reconfig_from_xcvr.reconfig_from_xcvr
		tx_parallel_data        : in  std_logic_vector(39 downto 0) := (others => '0'); --        tx_parallel_data.tx_parallel_data
		unused_tx_parallel_data : in  std_logic_vector(23 downto 0) := (others => '0'); -- unused_tx_parallel_data.unused_tx_parallel_data
		rx_parallel_data        : out std_logic_vector(39 downto 0);                    --        rx_parallel_data.rx_parallel_data
		unused_rx_parallel_data : out std_logic_vector(23 downto 0)                     -- unused_rx_parallel_data.unused_rx_parallel_data
	);
end entity gx_std_x4;

architecture rtl of gx_std_x4 is
	component altera_xcvr_native_sv is
		generic (
			tx_enable                       : integer := 1;
			rx_enable                       : integer := 1;
			enable_std                      : integer := 0;
			enable_teng                     : integer := 0;
			data_path_select                : string  := "pma_direct";
			channels                        : integer := 1;
			bonded_mode                     : string  := "non_bonded";
			data_rate                       : string  := "";
			pma_width                       : integer := 80;
			tx_pma_clk_div                  : integer := 1;
			tx_pma_txdetectrx_ctrl          : integer := 0;
			pll_reconfig_enable             : integer := 0;
			pll_external_enable             : integer := 0;
			pll_data_rate                   : string  := "0 Mbps";
			pll_type                        : string  := "CMU";
			pll_network_select              : string  := "x1";
			plls                            : integer := 1;
			pll_select                      : integer := 0;
			pll_refclk_cnt                  : integer := 1;
			pll_refclk_select               : string  := "0";
			pll_refclk_freq                 : string  := "125.0 MHz";
			pll_feedback_path               : string  := "internal";
			cdr_reconfig_enable             : integer := 0;
			cdr_refclk_cnt                  : integer := 1;
			cdr_refclk_select               : integer := 0;
			cdr_refclk_freq                 : string  := "";
			rx_ppm_detect_threshold         : string  := "1000";
			rx_clkslip_enable               : integer := 0;
			std_protocol_hint               : string  := "basic";
			std_pcs_pma_width               : integer := 10;
			std_low_latency_bypass_enable   : integer := 0;
			std_tx_pcfifo_mode              : string  := "low_latency";
			std_rx_pcfifo_mode              : string  := "low_latency";
			std_rx_byte_order_enable        : integer := 0;
			std_rx_byte_order_mode          : string  := "manual";
			std_rx_byte_order_width         : integer := 10;
			std_rx_byte_order_symbol_count  : integer := 1;
			std_rx_byte_order_pattern       : string  := "0";
			std_rx_byte_order_pad           : string  := "0";
			std_tx_byte_ser_enable          : integer := 0;
			std_rx_byte_deser_enable        : integer := 0;
			std_tx_8b10b_enable             : integer := 0;
			std_tx_8b10b_disp_ctrl_enable   : integer := 0;
			std_rx_8b10b_enable             : integer := 0;
			std_rx_rmfifo_enable            : integer := 0;
			std_rx_rmfifo_pattern_p         : string  := "00000";
			std_rx_rmfifo_pattern_n         : string  := "00000";
			std_tx_bitslip_enable           : integer := 0;
			std_rx_word_aligner_mode        : string  := "bit_slip";
			std_rx_word_aligner_pattern_len : integer := 7;
			std_rx_word_aligner_pattern     : string  := "0000000000";
			std_rx_word_aligner_rknumber    : integer := 3;
			std_rx_word_aligner_renumber    : integer := 3;
			std_rx_word_aligner_rgnumber    : integer := 3;
			std_rx_run_length_val           : integer := 31;
			std_tx_bitrev_enable            : integer := 0;
			std_rx_bitrev_enable            : integer := 0;
			std_tx_byterev_enable           : integer := 0;
			std_rx_byterev_enable           : integer := 0;
			std_tx_polinv_enable            : integer := 0;
			std_rx_polinv_enable            : integer := 0;
			teng_protocol_hint              : string  := "basic";
			teng_pcs_pma_width              : integer := 40;
			teng_pld_pcs_width              : integer := 40;
			teng_txfifo_mode                : string  := "phase_comp";
			teng_txfifo_full                : integer := 31;
			teng_txfifo_empty               : integer := 0;
			teng_txfifo_pfull               : integer := 23;
			teng_txfifo_pempty              : integer := 2;
			teng_rxfifo_mode                : string  := "phase_comp";
			teng_rxfifo_full                : integer := 31;
			teng_rxfifo_empty               : integer := 0;
			teng_rxfifo_pfull               : integer := 23;
			teng_rxfifo_pempty              : integer := 2;
			teng_rxfifo_align_del           : integer := 0;
			teng_rxfifo_control_del         : integer := 0;
			teng_tx_frmgen_enable           : integer := 0;
			teng_tx_frmgen_user_length      : integer := 2048;
			teng_tx_frmgen_burst_enable     : integer := 0;
			teng_rx_frmsync_enable          : integer := 0;
			teng_rx_frmsync_user_length     : integer := 2048;
			teng_frmgensync_diag_word       : string  := "6400000000000000";
			teng_frmgensync_scrm_word       : string  := "2800000000000000";
			teng_frmgensync_skip_word       : string  := "1e1e1e1e1e1e1e1e";
			teng_frmgensync_sync_word       : string  := "78f678f678f678f6";
			teng_tx_sh_err                  : integer := 0;
			teng_tx_crcgen_enable           : integer := 0;
			teng_rx_crcchk_enable           : integer := 0;
			teng_tx_64b66b_enable           : integer := 0;
			teng_rx_64b66b_enable           : integer := 0;
			teng_tx_scram_enable            : integer := 0;
			teng_tx_scram_user_seed         : string  := "000000000000000";
			teng_rx_descram_enable          : integer := 0;
			teng_tx_dispgen_enable          : integer := 0;
			teng_rx_dispchk_enable          : integer := 0;
			teng_rx_blksync_enable          : integer := 0;
			teng_tx_polinv_enable           : integer := 0;
			teng_tx_bitslip_enable          : integer := 0;
			teng_rx_polinv_enable           : integer := 0;
			teng_rx_bitslip_enable          : integer := 0
		);
		port (
			pll_powerdown             : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- pll_powerdown
			tx_analogreset            : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- tx_analogreset
			tx_digitalreset           : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- tx_digitalreset
			tx_serial_data            : out std_logic_vector(0 downto 0);                     -- tx_serial_data
			ext_pll_clk               : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- ext_pll_clk
			rx_analogreset            : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- rx_analogreset
			rx_digitalreset           : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- rx_digitalreset
			rx_cdr_refclk             : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- rx_cdr_refclk
			rx_serial_data            : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- rx_serial_data
			rx_is_lockedtoref         : out std_logic_vector(0 downto 0);                     -- rx_is_lockedtoref
			rx_is_lockedtodata        : out std_logic_vector(0 downto 0);                     -- rx_is_lockedtodata
			rx_seriallpbken           : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- rx_seriallpbken
			tx_std_coreclkin          : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- tx_std_coreclkin
			rx_std_coreclkin          : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- rx_std_coreclkin
			tx_std_clkout             : out std_logic_vector(0 downto 0);                     -- tx_std_clkout
			rx_std_clkout             : out std_logic_vector(0 downto 0);                     -- rx_std_clkout
			tx_std_polinv             : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- tx_std_polinv
			rx_std_polinv             : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- rx_std_polinv
			tx_cal_busy               : out std_logic_vector(0 downto 0);                     -- tx_cal_busy
			rx_cal_busy               : out std_logic_vector(0 downto 0);                     -- rx_cal_busy
			reconfig_to_xcvr          : in  std_logic_vector(69 downto 0) := (others => 'X'); -- reconfig_to_xcvr
			reconfig_from_xcvr        : out std_logic_vector(45 downto 0);                    -- reconfig_from_xcvr
			tx_parallel_data          : in  std_logic_vector(63 downto 0) := (others => 'X'); -- unused_tx_parallel_data
			rx_parallel_data          : out std_logic_vector(63 downto 0);                    -- unused_rx_parallel_data
			tx_pll_refclk             : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- tx_pll_refclk
			tx_pma_clkout             : out std_logic_vector(0 downto 0);                     -- tx_pma_clkout
			tx_pma_pclk               : out std_logic_vector(0 downto 0);                     -- tx_pma_pclk
			tx_pma_parallel_data      : in  std_logic_vector(79 downto 0) := (others => 'X'); -- tx_pma_parallel_data
			pll_locked                : out std_logic_vector(0 downto 0);                     -- pll_locked
			rx_pma_clkout             : out std_logic_vector(0 downto 0);                     -- rx_pma_clkout
			rx_pma_pclk               : out std_logic_vector(0 downto 0);                     -- rx_pma_pclk
			rx_pma_parallel_data      : out std_logic_vector(79 downto 0);                    -- rx_pma_parallel_data
			rx_clkslip                : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- rx_clkslip
			rx_clklow                 : out std_logic_vector(0 downto 0);                     -- rx_clklow
			rx_fref                   : out std_logic_vector(0 downto 0);                     -- rx_fref
			rx_set_locktodata         : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- rx_set_locktodata
			rx_set_locktoref          : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- rx_set_locktoref
			rx_signaldetect           : out std_logic_vector(0 downto 0);                     -- rx_signaldetect
			rx_pma_qpipulldn          : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- rx_pma_qpipulldn
			tx_pma_qpipullup          : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- tx_pma_qpipullup
			tx_pma_qpipulldn          : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- tx_pma_qpipulldn
			tx_pma_txdetectrx         : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- tx_pma_txdetectrx
			tx_pma_rxfound            : out std_logic_vector(0 downto 0);                     -- tx_pma_rxfound
			rx_std_prbs_done          : out std_logic_vector(0 downto 0);                     -- rx_std_prbs_done
			rx_std_prbs_err           : out std_logic_vector(0 downto 0);                     -- rx_std_prbs_err
			tx_std_pcfifo_full        : out std_logic_vector(0 downto 0);                     -- tx_std_pcfifo_full
			tx_std_pcfifo_empty       : out std_logic_vector(0 downto 0);                     -- tx_std_pcfifo_empty
			rx_std_pcfifo_full        : out std_logic_vector(0 downto 0);                     -- rx_std_pcfifo_full
			rx_std_pcfifo_empty       : out std_logic_vector(0 downto 0);                     -- rx_std_pcfifo_empty
			rx_std_byteorder_ena      : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- rx_std_byteorder_ena
			rx_std_byteorder_flag     : out std_logic_vector(0 downto 0);                     -- rx_std_byteorder_flag
			rx_std_rmfifo_full        : out std_logic_vector(0 downto 0);                     -- rx_std_rmfifo_full
			rx_std_rmfifo_empty       : out std_logic_vector(0 downto 0);                     -- rx_std_rmfifo_empty
			rx_std_wa_patternalign    : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- rx_std_wa_patternalign
			rx_std_wa_a1a2size        : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- rx_std_wa_a1a2size
			tx_std_bitslipboundarysel : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- tx_std_bitslipboundarysel
			rx_std_bitslipboundarysel : out std_logic_vector(4 downto 0);                     -- rx_std_bitslipboundarysel
			rx_std_bitslip            : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- rx_std_bitslip
			rx_std_runlength_err      : out std_logic_vector(0 downto 0);                     -- rx_std_runlength_err
			rx_std_bitrev_ena         : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- rx_std_bitrev_ena
			rx_std_byterev_ena        : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- rx_std_byterev_ena
			tx_std_elecidle           : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- tx_std_elecidle
			rx_std_signaldetect       : out std_logic_vector(0 downto 0);                     -- rx_std_signaldetect
			tx_10g_coreclkin          : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- tx_10g_coreclkin
			rx_10g_coreclkin          : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- rx_10g_coreclkin
			tx_10g_clkout             : out std_logic_vector(0 downto 0);                     -- tx_10g_clkout
			rx_10g_clkout             : out std_logic_vector(0 downto 0);                     -- rx_10g_clkout
			rx_10g_clk33out           : out std_logic_vector(0 downto 0);                     -- rx_10g_clk33out
			rx_10g_prbs_err_clr       : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- rx_10g_prbs_err_clr
			rx_10g_prbs_done          : out std_logic_vector(0 downto 0);                     -- rx_10g_prbs_done
			rx_10g_prbs_err           : out std_logic_vector(0 downto 0);                     -- rx_10g_prbs_err
			tx_10g_control            : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- tx_10g_control
			rx_10g_control            : out std_logic_vector(9 downto 0);                     -- rx_10g_control
			tx_10g_data_valid         : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- tx_10g_data_valid
			tx_10g_fifo_full          : out std_logic_vector(0 downto 0);                     -- tx_10g_fifo_full
			tx_10g_fifo_pfull         : out std_logic_vector(0 downto 0);                     -- tx_10g_fifo_pfull
			tx_10g_fifo_empty         : out std_logic_vector(0 downto 0);                     -- tx_10g_fifo_empty
			tx_10g_fifo_pempty        : out std_logic_vector(0 downto 0);                     -- tx_10g_fifo_pempty
			tx_10g_fifo_del           : out std_logic_vector(0 downto 0);                     -- tx_10g_fifo_del
			tx_10g_fifo_insert        : out std_logic_vector(0 downto 0);                     -- tx_10g_fifo_insert
			rx_10g_fifo_rd_en         : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- rx_10g_fifo_rd_en
			rx_10g_data_valid         : out std_logic_vector(0 downto 0);                     -- rx_10g_data_valid
			rx_10g_fifo_full          : out std_logic_vector(0 downto 0);                     -- rx_10g_fifo_full
			rx_10g_fifo_pfull         : out std_logic_vector(0 downto 0);                     -- rx_10g_fifo_pfull
			rx_10g_fifo_empty         : out std_logic_vector(0 downto 0);                     -- rx_10g_fifo_empty
			rx_10g_fifo_pempty        : out std_logic_vector(0 downto 0);                     -- rx_10g_fifo_pempty
			rx_10g_fifo_del           : out std_logic_vector(0 downto 0);                     -- rx_10g_fifo_del
			rx_10g_fifo_insert        : out std_logic_vector(0 downto 0);                     -- rx_10g_fifo_insert
			rx_10g_fifo_align_val     : out std_logic_vector(0 downto 0);                     -- rx_10g_fifo_align_val
			rx_10g_fifo_align_clr     : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- rx_10g_fifo_align_clr
			rx_10g_fifo_align_en      : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- rx_10g_fifo_align_en
			tx_10g_frame              : out std_logic_vector(0 downto 0);                     -- tx_10g_frame
			tx_10g_frame_diag_status  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- tx_10g_frame_diag_status
			tx_10g_frame_burst_en     : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- tx_10g_frame_burst_en
			rx_10g_frame              : out std_logic_vector(0 downto 0);                     -- rx_10g_frame
			rx_10g_frame_lock         : out std_logic_vector(0 downto 0);                     -- rx_10g_frame_lock
			rx_10g_frame_mfrm_err     : out std_logic_vector(0 downto 0);                     -- rx_10g_frame_mfrm_err
			rx_10g_frame_sync_err     : out std_logic_vector(0 downto 0);                     -- rx_10g_frame_sync_err
			rx_10g_frame_skip_ins     : out std_logic_vector(0 downto 0);                     -- rx_10g_frame_skip_ins
			rx_10g_frame_pyld_ins     : out std_logic_vector(0 downto 0);                     -- rx_10g_frame_pyld_ins
			rx_10g_frame_skip_err     : out std_logic_vector(0 downto 0);                     -- rx_10g_frame_skip_err
			rx_10g_frame_diag_err     : out std_logic_vector(0 downto 0);                     -- rx_10g_frame_diag_err
			rx_10g_frame_diag_status  : out std_logic_vector(1 downto 0);                     -- rx_10g_frame_diag_status
			rx_10g_crc32_err          : out std_logic_vector(0 downto 0);                     -- rx_10g_crc32err
			rx_10g_descram_err        : out std_logic_vector(0 downto 0);                     -- rx_10g_descram_err
			rx_10g_blk_lock           : out std_logic_vector(0 downto 0);                     -- rx_10g_blk_lock
			rx_10g_blk_sh_err         : out std_logic_vector(0 downto 0);                     -- rx_10g_blk_sh_err
			tx_10g_bitslip            : in  std_logic_vector(6 downto 0)  := (others => 'X'); -- tx_10g_bitslip
			rx_10g_bitslip            : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- rx_10g_bitslip
			rx_10g_highber            : out std_logic_vector(0 downto 0);                     -- rx_10g_highber
			rx_10g_highber_clr_cnt    : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- rx_10g_highber_clr_cnt
			rx_10g_clr_errblk_count   : in  std_logic_vector(0 downto 0)  := (others => 'X')  -- rx_10g_clr_errblk_count
		);
	end component altera_xcvr_native_sv;

	signal gx_std_x4_inst_rx_parallel_data : std_logic_vector(63 downto 0); -- port fragment

begin

	gx_std_x4_inst : component altera_xcvr_native_sv
		generic map (
			tx_enable                       => 1,
			rx_enable                       => 1,
			enable_std                      => 1,
			enable_teng                     => 0,
			data_path_select                => "standard",
			channels                        => 1,
			bonded_mode                     => "xN",
			data_rate                       => "4800 Mbps",
			pma_width                       => 20,
			tx_pma_clk_div                  => 1,
			tx_pma_txdetectrx_ctrl          => 0,
			pll_reconfig_enable             => 0,
			pll_external_enable             => 1,
			pll_data_rate                   => "4800 Mbps",
			pll_type                        => "CMU",
			pll_network_select              => "x1",
			plls                            => 1,
			pll_select                      => 0,
			pll_refclk_cnt                  => 1,
			pll_refclk_select               => "0",
			pll_refclk_freq                 => "125.0 MHz",
			pll_feedback_path               => "internal",
			cdr_reconfig_enable             => 0,
			cdr_refclk_cnt                  => 1,
			cdr_refclk_select               => 0,
			cdr_refclk_freq                 => "120.0 MHz",
			rx_ppm_detect_threshold         => "1000",
			rx_clkslip_enable               => 0,
			std_protocol_hint               => "basic",
			std_pcs_pma_width               => 20,
			std_low_latency_bypass_enable   => 0,
			std_tx_pcfifo_mode              => "low_latency",
			std_rx_pcfifo_mode              => "low_latency",
			std_rx_byte_order_enable        => 0,
			std_rx_byte_order_mode          => "manual",
			std_rx_byte_order_width         => 10,
			std_rx_byte_order_symbol_count  => 1,
			std_rx_byte_order_pattern       => "0",
			std_rx_byte_order_pad           => "0",
			std_tx_byte_ser_enable          => 1,
			std_rx_byte_deser_enable        => 1,
			std_tx_8b10b_enable             => 0,
			std_tx_8b10b_disp_ctrl_enable   => 0,
			std_rx_8b10b_enable             => 0,
			std_rx_rmfifo_enable            => 0,
			std_rx_rmfifo_pattern_p         => "00000",
			std_rx_rmfifo_pattern_n         => "00000",
			std_tx_bitslip_enable           => 0,
			std_rx_word_aligner_mode        => "bit_slip",
			std_rx_word_aligner_pattern_len => 7,
			std_rx_word_aligner_pattern     => "0000000000",
			std_rx_word_aligner_rknumber    => 3,
			std_rx_word_aligner_renumber    => 3,
			std_rx_word_aligner_rgnumber    => 3,
			std_rx_run_length_val           => 31,
			std_tx_bitrev_enable            => 0,
			std_rx_bitrev_enable            => 0,
			std_tx_byterev_enable           => 0,
			std_rx_byterev_enable           => 0,
			std_tx_polinv_enable            => 1,
			std_rx_polinv_enable            => 1,
			teng_protocol_hint              => "basic",
			teng_pcs_pma_width              => 40,
			teng_pld_pcs_width              => 40,
			teng_txfifo_mode                => "phase_comp",
			teng_txfifo_full                => 31,
			teng_txfifo_empty               => 0,
			teng_txfifo_pfull               => 23,
			teng_txfifo_pempty              => 2,
			teng_rxfifo_mode                => "phase_comp",
			teng_rxfifo_full                => 31,
			teng_rxfifo_empty               => 0,
			teng_rxfifo_pfull               => 23,
			teng_rxfifo_pempty              => 2,
			teng_rxfifo_align_del           => 0,
			teng_rxfifo_control_del         => 0,
			teng_tx_frmgen_enable           => 0,
			teng_tx_frmgen_user_length      => 2048,
			teng_tx_frmgen_burst_enable     => 0,
			teng_rx_frmsync_enable          => 0,
			teng_rx_frmsync_user_length     => 2048,
			teng_frmgensync_diag_word       => "6400000000000000",
			teng_frmgensync_scrm_word       => "2800000000000000",
			teng_frmgensync_skip_word       => "1e1e1e1e1e1e1e1e",
			teng_frmgensync_sync_word       => "78f678f678f678f6",
			teng_tx_sh_err                  => 0,
			teng_tx_crcgen_enable           => 0,
			teng_rx_crcchk_enable           => 0,
			teng_tx_64b66b_enable           => 0,
			teng_rx_64b66b_enable           => 0,
			teng_tx_scram_enable            => 0,
			teng_tx_scram_user_seed         => "000000000000000",
			teng_rx_descram_enable          => 0,
			teng_tx_dispgen_enable          => 0,
			teng_rx_dispchk_enable          => 0,
			teng_rx_blksync_enable          => 0,
			teng_tx_polinv_enable           => 0,
			teng_tx_bitslip_enable          => 0,
			teng_rx_polinv_enable           => 0,
			teng_rx_bitslip_enable          => 0
		)
		port map (
			pll_powerdown             => pll_powerdown,                                                                      --      pll_powerdown.pll_powerdown
			tx_analogreset            => tx_analogreset,                                                                     --     tx_analogreset.tx_analogreset
			tx_digitalreset           => tx_digitalreset,                                                                    --    tx_digitalreset.tx_digitalreset
			tx_serial_data            => tx_serial_data,                                                                     --     tx_serial_data.tx_serial_data
			ext_pll_clk               => ext_pll_clk,                                                                        --        ext_pll_clk.ext_pll_clk
			rx_analogreset            => rx_analogreset,                                                                     --     rx_analogreset.rx_analogreset
			rx_digitalreset           => rx_digitalreset,                                                                    --    rx_digitalreset.rx_digitalreset
			rx_cdr_refclk             => rx_cdr_refclk,                                                                      --      rx_cdr_refclk.rx_cdr_refclk
			rx_serial_data            => rx_serial_data,                                                                     --     rx_serial_data.rx_serial_data
			rx_is_lockedtoref         => rx_is_lockedtoref,                                                                  --  rx_is_lockedtoref.rx_is_lockedtoref
			rx_is_lockedtodata        => rx_is_lockedtodata,                                                                 -- rx_is_lockedtodata.rx_is_lockedtodata
			rx_seriallpbken           => rx_seriallpbken,                                                                    --    rx_seriallpbken.rx_seriallpbken
			tx_std_coreclkin          => tx_std_coreclkin,                                                                   --   tx_std_coreclkin.tx_std_coreclkin
			rx_std_coreclkin          => rx_std_coreclkin,                                                                   --   rx_std_coreclkin.rx_std_coreclkin
			tx_std_clkout             => tx_std_clkout,                                                                      --      tx_std_clkout.tx_std_clkout
			rx_std_clkout             => rx_std_clkout,                                                                      --      rx_std_clkout.rx_std_clkout
			tx_std_polinv             => tx_std_polinv,                                                                      --      tx_std_polinv.tx_std_polinv
			rx_std_polinv             => rx_std_polinv,                                                                      --      rx_std_polinv.rx_std_polinv
			tx_cal_busy               => tx_cal_busy,                                                                        --        tx_cal_busy.tx_cal_busy
			rx_cal_busy               => rx_cal_busy,                                                                        --        rx_cal_busy.rx_cal_busy
			reconfig_to_xcvr          => reconfig_to_xcvr,                                                                   --   reconfig_to_xcvr.reconfig_to_xcvr
			reconfig_from_xcvr        => reconfig_from_xcvr,                                                                 -- reconfig_from_xcvr.reconfig_from_xcvr
			tx_parallel_data(0)       => tx_parallel_data(0),                                                                --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(1)       => tx_parallel_data(1),                                                                --                   .tx_parallel_data
			tx_parallel_data(2)       => tx_parallel_data(2),                                                                --                   .tx_parallel_data
			tx_parallel_data(3)       => tx_parallel_data(3),                                                                --                   .tx_parallel_data
			tx_parallel_data(4)       => tx_parallel_data(4),                                                                --                   .tx_parallel_data
			tx_parallel_data(5)       => tx_parallel_data(5),                                                                --                   .tx_parallel_data
			tx_parallel_data(6)       => tx_parallel_data(6),                                                                --                   .tx_parallel_data
			tx_parallel_data(7)       => tx_parallel_data(7),                                                                --                   .tx_parallel_data
			tx_parallel_data(8)       => tx_parallel_data(8),                                                                --                   .tx_parallel_data
			tx_parallel_data(9)       => tx_parallel_data(9),                                                                --                   .tx_parallel_data
			tx_parallel_data(10)      => unused_tx_parallel_data(0),                                                         --                   .tx_parallel_data
			tx_parallel_data(11)      => tx_parallel_data(10),                                                               --                   .tx_parallel_data
			tx_parallel_data(12)      => tx_parallel_data(11),                                                               --                   .tx_parallel_data
			tx_parallel_data(13)      => tx_parallel_data(12),                                                               --                   .tx_parallel_data
			tx_parallel_data(14)      => tx_parallel_data(13),                                                               --                   .tx_parallel_data
			tx_parallel_data(15)      => tx_parallel_data(14),                                                               --                   .tx_parallel_data
			tx_parallel_data(16)      => tx_parallel_data(15),                                                               --                   .tx_parallel_data
			tx_parallel_data(17)      => tx_parallel_data(16),                                                               --                   .tx_parallel_data
			tx_parallel_data(18)      => tx_parallel_data(17),                                                               --                   .tx_parallel_data
			tx_parallel_data(19)      => tx_parallel_data(18),                                                               --                   .tx_parallel_data
			tx_parallel_data(20)      => tx_parallel_data(19),                                                               --                   .tx_parallel_data
			tx_parallel_data(21)      => unused_tx_parallel_data(1),                                                         --                   .tx_parallel_data
			tx_parallel_data(22)      => tx_parallel_data(20),                                                               --                   .tx_parallel_data
			tx_parallel_data(23)      => tx_parallel_data(21),                                                               --                   .tx_parallel_data
			tx_parallel_data(24)      => tx_parallel_data(22),                                                               --                   .tx_parallel_data
			tx_parallel_data(25)      => tx_parallel_data(23),                                                               --                   .tx_parallel_data
			tx_parallel_data(26)      => tx_parallel_data(24),                                                               --                   .tx_parallel_data
			tx_parallel_data(27)      => tx_parallel_data(25),                                                               --                   .tx_parallel_data
			tx_parallel_data(28)      => tx_parallel_data(26),                                                               --                   .tx_parallel_data
			tx_parallel_data(29)      => tx_parallel_data(27),                                                               --                   .tx_parallel_data
			tx_parallel_data(30)      => tx_parallel_data(28),                                                               --                   .tx_parallel_data
			tx_parallel_data(31)      => tx_parallel_data(29),                                                               --                   .tx_parallel_data
			tx_parallel_data(32)      => unused_tx_parallel_data(2),                                                         --                   .tx_parallel_data
			tx_parallel_data(33)      => tx_parallel_data(30),                                                               --                   .tx_parallel_data
			tx_parallel_data(34)      => tx_parallel_data(31),                                                               --                   .tx_parallel_data
			tx_parallel_data(35)      => tx_parallel_data(32),                                                               --                   .tx_parallel_data
			tx_parallel_data(36)      => tx_parallel_data(33),                                                               --                   .tx_parallel_data
			tx_parallel_data(37)      => tx_parallel_data(34),                                                               --                   .tx_parallel_data
			tx_parallel_data(38)      => tx_parallel_data(35),                                                               --                   .tx_parallel_data
			tx_parallel_data(39)      => tx_parallel_data(36),                                                               --                   .tx_parallel_data
			tx_parallel_data(40)      => tx_parallel_data(37),                                                               --                   .tx_parallel_data
			tx_parallel_data(41)      => tx_parallel_data(38),                                                               --                   .tx_parallel_data
			tx_parallel_data(42)      => tx_parallel_data(39),                                                               --                   .tx_parallel_data
			tx_parallel_data(43)      => unused_tx_parallel_data(3),                                                         --                   .tx_parallel_data
			tx_parallel_data(44)      => unused_tx_parallel_data(4),                                                         --                   .tx_parallel_data
			tx_parallel_data(45)      => unused_tx_parallel_data(5),                                                         --                   .tx_parallel_data
			tx_parallel_data(46)      => unused_tx_parallel_data(6),                                                         --                   .tx_parallel_data
			tx_parallel_data(47)      => unused_tx_parallel_data(7),                                                         --                   .tx_parallel_data
			tx_parallel_data(48)      => unused_tx_parallel_data(8),                                                         --                   .tx_parallel_data
			tx_parallel_data(49)      => unused_tx_parallel_data(9),                                                         --                   .tx_parallel_data
			tx_parallel_data(50)      => unused_tx_parallel_data(10),                                                        --                   .tx_parallel_data
			tx_parallel_data(51)      => unused_tx_parallel_data(11),                                                        --                   .tx_parallel_data
			tx_parallel_data(52)      => unused_tx_parallel_data(12),                                                        --                   .tx_parallel_data
			tx_parallel_data(53)      => unused_tx_parallel_data(13),                                                        --                   .tx_parallel_data
			tx_parallel_data(54)      => unused_tx_parallel_data(14),                                                        --                   .tx_parallel_data
			tx_parallel_data(55)      => unused_tx_parallel_data(15),                                                        --                   .tx_parallel_data
			tx_parallel_data(56)      => unused_tx_parallel_data(16),                                                        --                   .tx_parallel_data
			tx_parallel_data(57)      => unused_tx_parallel_data(17),                                                        --                   .tx_parallel_data
			tx_parallel_data(58)      => unused_tx_parallel_data(18),                                                        --                   .tx_parallel_data
			tx_parallel_data(59)      => unused_tx_parallel_data(19),                                                        --                   .tx_parallel_data
			tx_parallel_data(60)      => unused_tx_parallel_data(20),                                                        --                   .tx_parallel_data
			tx_parallel_data(61)      => unused_tx_parallel_data(21),                                                        --                   .tx_parallel_data
			tx_parallel_data(62)      => unused_tx_parallel_data(22),                                                        --                   .tx_parallel_data
			tx_parallel_data(63)      => unused_tx_parallel_data(23),                                                        --                   .tx_parallel_data
			rx_parallel_data(0)       => gx_std_x4_inst_rx_parallel_data(0),                                                 --   rx_parallel_data.rx_parallel_data
			rx_parallel_data(1)       => gx_std_x4_inst_rx_parallel_data(1),                                                 --                   .rx_parallel_data
			rx_parallel_data(2)       => gx_std_x4_inst_rx_parallel_data(2),                                                 --                   .rx_parallel_data
			rx_parallel_data(3)       => gx_std_x4_inst_rx_parallel_data(3),                                                 --                   .rx_parallel_data
			rx_parallel_data(4)       => gx_std_x4_inst_rx_parallel_data(4),                                                 --                   .rx_parallel_data
			rx_parallel_data(5)       => gx_std_x4_inst_rx_parallel_data(5),                                                 --                   .rx_parallel_data
			rx_parallel_data(6)       => gx_std_x4_inst_rx_parallel_data(6),                                                 --                   .rx_parallel_data
			rx_parallel_data(7)       => gx_std_x4_inst_rx_parallel_data(7),                                                 --                   .rx_parallel_data
			rx_parallel_data(8)       => gx_std_x4_inst_rx_parallel_data(8),                                                 --                   .rx_parallel_data
			rx_parallel_data(9)       => gx_std_x4_inst_rx_parallel_data(9),                                                 --                   .rx_parallel_data
			rx_parallel_data(10)      => gx_std_x4_inst_rx_parallel_data(10),                                                --                   .rx_parallel_data
			rx_parallel_data(11)      => gx_std_x4_inst_rx_parallel_data(11),                                                --                   .rx_parallel_data
			rx_parallel_data(12)      => gx_std_x4_inst_rx_parallel_data(12),                                                --                   .rx_parallel_data
			rx_parallel_data(13)      => gx_std_x4_inst_rx_parallel_data(13),                                                --                   .rx_parallel_data
			rx_parallel_data(14)      => gx_std_x4_inst_rx_parallel_data(14),                                                --                   .rx_parallel_data
			rx_parallel_data(15)      => gx_std_x4_inst_rx_parallel_data(15),                                                --                   .rx_parallel_data
			rx_parallel_data(16)      => gx_std_x4_inst_rx_parallel_data(16),                                                --                   .rx_parallel_data
			rx_parallel_data(17)      => gx_std_x4_inst_rx_parallel_data(17),                                                --                   .rx_parallel_data
			rx_parallel_data(18)      => gx_std_x4_inst_rx_parallel_data(18),                                                --                   .rx_parallel_data
			rx_parallel_data(19)      => gx_std_x4_inst_rx_parallel_data(19),                                                --                   .rx_parallel_data
			rx_parallel_data(20)      => gx_std_x4_inst_rx_parallel_data(20),                                                --                   .rx_parallel_data
			rx_parallel_data(21)      => gx_std_x4_inst_rx_parallel_data(21),                                                --                   .rx_parallel_data
			rx_parallel_data(22)      => gx_std_x4_inst_rx_parallel_data(22),                                                --                   .rx_parallel_data
			rx_parallel_data(23)      => gx_std_x4_inst_rx_parallel_data(23),                                                --                   .rx_parallel_data
			rx_parallel_data(24)      => gx_std_x4_inst_rx_parallel_data(24),                                                --                   .rx_parallel_data
			rx_parallel_data(25)      => gx_std_x4_inst_rx_parallel_data(25),                                                --                   .rx_parallel_data
			rx_parallel_data(26)      => gx_std_x4_inst_rx_parallel_data(26),                                                --                   .rx_parallel_data
			rx_parallel_data(27)      => gx_std_x4_inst_rx_parallel_data(27),                                                --                   .rx_parallel_data
			rx_parallel_data(28)      => gx_std_x4_inst_rx_parallel_data(28),                                                --                   .rx_parallel_data
			rx_parallel_data(29)      => gx_std_x4_inst_rx_parallel_data(29),                                                --                   .rx_parallel_data
			rx_parallel_data(30)      => gx_std_x4_inst_rx_parallel_data(30),                                                --                   .rx_parallel_data
			rx_parallel_data(31)      => gx_std_x4_inst_rx_parallel_data(31),                                                --                   .rx_parallel_data
			rx_parallel_data(32)      => gx_std_x4_inst_rx_parallel_data(32),                                                --                   .rx_parallel_data
			rx_parallel_data(33)      => gx_std_x4_inst_rx_parallel_data(33),                                                --                   .rx_parallel_data
			rx_parallel_data(34)      => gx_std_x4_inst_rx_parallel_data(34),                                                --                   .rx_parallel_data
			rx_parallel_data(35)      => gx_std_x4_inst_rx_parallel_data(35),                                                --                   .rx_parallel_data
			rx_parallel_data(36)      => gx_std_x4_inst_rx_parallel_data(36),                                                --                   .rx_parallel_data
			rx_parallel_data(37)      => gx_std_x4_inst_rx_parallel_data(37),                                                --                   .rx_parallel_data
			rx_parallel_data(38)      => gx_std_x4_inst_rx_parallel_data(38),                                                --                   .rx_parallel_data
			rx_parallel_data(39)      => gx_std_x4_inst_rx_parallel_data(39),                                                --                   .rx_parallel_data
			rx_parallel_data(40)      => gx_std_x4_inst_rx_parallel_data(40),                                                --                   .rx_parallel_data
			rx_parallel_data(41)      => gx_std_x4_inst_rx_parallel_data(41),                                                --                   .rx_parallel_data
			rx_parallel_data(42)      => gx_std_x4_inst_rx_parallel_data(42),                                                --                   .rx_parallel_data
			rx_parallel_data(43)      => gx_std_x4_inst_rx_parallel_data(43),                                                --                   .rx_parallel_data
			rx_parallel_data(44)      => gx_std_x4_inst_rx_parallel_data(44),                                                --                   .rx_parallel_data
			rx_parallel_data(45)      => gx_std_x4_inst_rx_parallel_data(45),                                                --                   .rx_parallel_data
			rx_parallel_data(46)      => gx_std_x4_inst_rx_parallel_data(46),                                                --                   .rx_parallel_data
			rx_parallel_data(47)      => gx_std_x4_inst_rx_parallel_data(47),                                                --                   .rx_parallel_data
			rx_parallel_data(48)      => gx_std_x4_inst_rx_parallel_data(48),                                                --                   .rx_parallel_data
			rx_parallel_data(49)      => gx_std_x4_inst_rx_parallel_data(49),                                                --                   .rx_parallel_data
			rx_parallel_data(50)      => gx_std_x4_inst_rx_parallel_data(50),                                                --                   .rx_parallel_data
			rx_parallel_data(51)      => gx_std_x4_inst_rx_parallel_data(51),                                                --                   .rx_parallel_data
			rx_parallel_data(52)      => gx_std_x4_inst_rx_parallel_data(52),                                                --                   .rx_parallel_data
			rx_parallel_data(53)      => gx_std_x4_inst_rx_parallel_data(53),                                                --                   .rx_parallel_data
			rx_parallel_data(54)      => gx_std_x4_inst_rx_parallel_data(54),                                                --                   .rx_parallel_data
			rx_parallel_data(55)      => gx_std_x4_inst_rx_parallel_data(55),                                                --                   .rx_parallel_data
			rx_parallel_data(56)      => gx_std_x4_inst_rx_parallel_data(56),                                                --                   .rx_parallel_data
			rx_parallel_data(57)      => gx_std_x4_inst_rx_parallel_data(57),                                                --                   .rx_parallel_data
			rx_parallel_data(58)      => gx_std_x4_inst_rx_parallel_data(58),                                                --                   .rx_parallel_data
			rx_parallel_data(59)      => gx_std_x4_inst_rx_parallel_data(59),                                                --                   .rx_parallel_data
			rx_parallel_data(60)      => gx_std_x4_inst_rx_parallel_data(60),                                                --                   .rx_parallel_data
			rx_parallel_data(61)      => gx_std_x4_inst_rx_parallel_data(61),                                                --                   .rx_parallel_data
			rx_parallel_data(62)      => gx_std_x4_inst_rx_parallel_data(62),                                                --                   .rx_parallel_data
			rx_parallel_data(63)      => gx_std_x4_inst_rx_parallel_data(63),                                                --                   .rx_parallel_data
			tx_pll_refclk             => "0",                                                                                --        (terminated)
			tx_pma_clkout             => open,                                                                               --        (terminated)
			tx_pma_pclk               => open,                                                                               --        (terminated)
			tx_pma_parallel_data      => "00000000000000000000000000000000000000000000000000000000000000000000000000000000", --        (terminated)
			pll_locked                => open,                                                                               --        (terminated)
			rx_pma_clkout             => open,                                                                               --        (terminated)
			rx_pma_pclk               => open,                                                                               --        (terminated)
			rx_pma_parallel_data      => open,                                                                               --        (terminated)
			rx_clkslip                => "0",                                                                                --        (terminated)
			rx_clklow                 => open,                                                                               --        (terminated)
			rx_fref                   => open,                                                                               --        (terminated)
			rx_set_locktodata         => "0",                                                                                --        (terminated)
			rx_set_locktoref          => "0",                                                                                --        (terminated)
			rx_signaldetect           => open,                                                                               --        (terminated)
			rx_pma_qpipulldn          => "0",                                                                                --        (terminated)
			tx_pma_qpipullup          => "0",                                                                                --        (terminated)
			tx_pma_qpipulldn          => "0",                                                                                --        (terminated)
			tx_pma_txdetectrx         => "0",                                                                                --        (terminated)
			tx_pma_rxfound            => open,                                                                               --        (terminated)
			rx_std_prbs_done          => open,                                                                               --        (terminated)
			rx_std_prbs_err           => open,                                                                               --        (terminated)
			tx_std_pcfifo_full        => open,                                                                               --        (terminated)
			tx_std_pcfifo_empty       => open,                                                                               --        (terminated)
			rx_std_pcfifo_full        => open,                                                                               --        (terminated)
			rx_std_pcfifo_empty       => open,                                                                               --        (terminated)
			rx_std_byteorder_ena      => "0",                                                                                --        (terminated)
			rx_std_byteorder_flag     => open,                                                                               --        (terminated)
			rx_std_rmfifo_full        => open,                                                                               --        (terminated)
			rx_std_rmfifo_empty       => open,                                                                               --        (terminated)
			rx_std_wa_patternalign    => "0",                                                                                --        (terminated)
			rx_std_wa_a1a2size        => "0",                                                                                --        (terminated)
			tx_std_bitslipboundarysel => "00000",                                                                            --        (terminated)
			rx_std_bitslipboundarysel => open,                                                                               --        (terminated)
			rx_std_bitslip            => "0",                                                                                --        (terminated)
			rx_std_runlength_err      => open,                                                                               --        (terminated)
			rx_std_bitrev_ena         => "0",                                                                                --        (terminated)
			rx_std_byterev_ena        => "0",                                                                                --        (terminated)
			tx_std_elecidle           => "0",                                                                                --        (terminated)
			rx_std_signaldetect       => open,                                                                               --        (terminated)
			tx_10g_coreclkin          => "0",                                                                                --        (terminated)
			rx_10g_coreclkin          => "0",                                                                                --        (terminated)
			tx_10g_clkout             => open,                                                                               --        (terminated)
			rx_10g_clkout             => open,                                                                               --        (terminated)
			rx_10g_clk33out           => open,                                                                               --        (terminated)
			rx_10g_prbs_err_clr       => "0",                                                                                --        (terminated)
			rx_10g_prbs_done          => open,                                                                               --        (terminated)
			rx_10g_prbs_err           => open,                                                                               --        (terminated)
			tx_10g_control            => "000000000",                                                                        --        (terminated)
			rx_10g_control            => open,                                                                               --        (terminated)
			tx_10g_data_valid         => "0",                                                                                --        (terminated)
			tx_10g_fifo_full          => open,                                                                               --        (terminated)
			tx_10g_fifo_pfull         => open,                                                                               --        (terminated)
			tx_10g_fifo_empty         => open,                                                                               --        (terminated)
			tx_10g_fifo_pempty        => open,                                                                               --        (terminated)
			tx_10g_fifo_del           => open,                                                                               --        (terminated)
			tx_10g_fifo_insert        => open,                                                                               --        (terminated)
			rx_10g_fifo_rd_en         => "0",                                                                                --        (terminated)
			rx_10g_data_valid         => open,                                                                               --        (terminated)
			rx_10g_fifo_full          => open,                                                                               --        (terminated)
			rx_10g_fifo_pfull         => open,                                                                               --        (terminated)
			rx_10g_fifo_empty         => open,                                                                               --        (terminated)
			rx_10g_fifo_pempty        => open,                                                                               --        (terminated)
			rx_10g_fifo_del           => open,                                                                               --        (terminated)
			rx_10g_fifo_insert        => open,                                                                               --        (terminated)
			rx_10g_fifo_align_val     => open,                                                                               --        (terminated)
			rx_10g_fifo_align_clr     => "0",                                                                                --        (terminated)
			rx_10g_fifo_align_en      => "0",                                                                                --        (terminated)
			tx_10g_frame              => open,                                                                               --        (terminated)
			tx_10g_frame_diag_status  => "00",                                                                               --        (terminated)
			tx_10g_frame_burst_en     => "0",                                                                                --        (terminated)
			rx_10g_frame              => open,                                                                               --        (terminated)
			rx_10g_frame_lock         => open,                                                                               --        (terminated)
			rx_10g_frame_mfrm_err     => open,                                                                               --        (terminated)
			rx_10g_frame_sync_err     => open,                                                                               --        (terminated)
			rx_10g_frame_skip_ins     => open,                                                                               --        (terminated)
			rx_10g_frame_pyld_ins     => open,                                                                               --        (terminated)
			rx_10g_frame_skip_err     => open,                                                                               --        (terminated)
			rx_10g_frame_diag_err     => open,                                                                               --        (terminated)
			rx_10g_frame_diag_status  => open,                                                                               --        (terminated)
			rx_10g_crc32_err          => open,                                                                               --        (terminated)
			rx_10g_descram_err        => open,                                                                               --        (terminated)
			rx_10g_blk_lock           => open,                                                                               --        (terminated)
			rx_10g_blk_sh_err         => open,                                                                               --        (terminated)
			tx_10g_bitslip            => "0000000",                                                                          --        (terminated)
			rx_10g_bitslip            => "0",                                                                                --        (terminated)
			rx_10g_highber            => open,                                                                               --        (terminated)
			rx_10g_highber_clr_cnt    => "0",                                                                                --        (terminated)
			rx_10g_clr_errblk_count   => "0"                                                                                 --        (terminated)
		);

	unused_rx_parallel_data <= gx_std_x4_inst_rx_parallel_data(63) & gx_std_x4_inst_rx_parallel_data(62) & gx_std_x4_inst_rx_parallel_data(61) & gx_std_x4_inst_rx_parallel_data(60) & gx_std_x4_inst_rx_parallel_data(59) & gx_std_x4_inst_rx_parallel_data(58) & gx_std_x4_inst_rx_parallel_data(47) & gx_std_x4_inst_rx_parallel_data(46) & gx_std_x4_inst_rx_parallel_data(45) & gx_std_x4_inst_rx_parallel_data(44) & gx_std_x4_inst_rx_parallel_data(43) & gx_std_x4_inst_rx_parallel_data(42) & gx_std_x4_inst_rx_parallel_data(31) & gx_std_x4_inst_rx_parallel_data(30) & gx_std_x4_inst_rx_parallel_data(29) & gx_std_x4_inst_rx_parallel_data(28) & gx_std_x4_inst_rx_parallel_data(27) & gx_std_x4_inst_rx_parallel_data(26) & gx_std_x4_inst_rx_parallel_data(15) & gx_std_x4_inst_rx_parallel_data(14) & gx_std_x4_inst_rx_parallel_data(13) & gx_std_x4_inst_rx_parallel_data(12) & gx_std_x4_inst_rx_parallel_data(11) & gx_std_x4_inst_rx_parallel_data(10);

	rx_parallel_data <= gx_std_x4_inst_rx_parallel_data(57) & gx_std_x4_inst_rx_parallel_data(56) & gx_std_x4_inst_rx_parallel_data(55) & gx_std_x4_inst_rx_parallel_data(54) & gx_std_x4_inst_rx_parallel_data(53) & gx_std_x4_inst_rx_parallel_data(52) & gx_std_x4_inst_rx_parallel_data(51) & gx_std_x4_inst_rx_parallel_data(50) & gx_std_x4_inst_rx_parallel_data(49) & gx_std_x4_inst_rx_parallel_data(48) & gx_std_x4_inst_rx_parallel_data(41) & gx_std_x4_inst_rx_parallel_data(40) & gx_std_x4_inst_rx_parallel_data(39) & gx_std_x4_inst_rx_parallel_data(38) & gx_std_x4_inst_rx_parallel_data(37) & gx_std_x4_inst_rx_parallel_data(36) & gx_std_x4_inst_rx_parallel_data(35) & gx_std_x4_inst_rx_parallel_data(34) & gx_std_x4_inst_rx_parallel_data(33) & gx_std_x4_inst_rx_parallel_data(32) & gx_std_x4_inst_rx_parallel_data(25) & gx_std_x4_inst_rx_parallel_data(24) & gx_std_x4_inst_rx_parallel_data(23) & gx_std_x4_inst_rx_parallel_data(22) & gx_std_x4_inst_rx_parallel_data(21) & gx_std_x4_inst_rx_parallel_data(20) & gx_std_x4_inst_rx_parallel_data(19) & gx_std_x4_inst_rx_parallel_data(18) & gx_std_x4_inst_rx_parallel_data(17) & gx_std_x4_inst_rx_parallel_data(16) & gx_std_x4_inst_rx_parallel_data(9) & gx_std_x4_inst_rx_parallel_data(8) & gx_std_x4_inst_rx_parallel_data(7) & gx_std_x4_inst_rx_parallel_data(6) & gx_std_x4_inst_rx_parallel_data(5) & gx_std_x4_inst_rx_parallel_data(4) & gx_std_x4_inst_rx_parallel_data(3) & gx_std_x4_inst_rx_parallel_data(2) & gx_std_x4_inst_rx_parallel_data(1) & gx_std_x4_inst_rx_parallel_data(0);

end architecture rtl; -- of gx_std_x4
