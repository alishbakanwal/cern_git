-- mgt_pll.vhd

-- Generated using ACDS version 15.1 185

library IEEE;
library mgt_pll_altera_xcvr_fpll_a10_151;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity mgt_pll is
	port (
		mcgb_rst          : in  std_logic                    := '0'; --          mcgb_rst.mcgb_rst
		pll_cal_busy      : out std_logic;                           --      pll_cal_busy.pll_cal_busy
		pll_locked        : out std_logic;                           --        pll_locked.pll_locked
		pll_powerdown     : in  std_logic                    := '0'; --     pll_powerdown.pll_powerdown
		pll_refclk0       : in  std_logic                    := '0'; --       pll_refclk0.clk
		tx_bonding_clocks : out std_logic_vector(5 downto 0);        -- tx_bonding_clocks.clk
		tx_serial_clk     : out std_logic                            --     tx_serial_clk.clk
	);
end entity mgt_pll;

architecture rtl of mgt_pll is
	component altera_xcvr_fpll_a10 is
		generic (
			enable_pll_reconfig                                                          : integer := 0;
			rcfg_jtag_enable                                                             : integer := 0;
			rcfg_separate_avmm_busy                                                      : integer := 0;
			dbg_embedded_debug_enable                                                    : integer := 0;
			dbg_capability_reg_enable                                                    : integer := 0;
			dbg_user_identifier                                                          : integer := 0;
			dbg_stat_soft_logic_enable                                                   : integer := 0;
			dbg_ctrl_soft_logic_enable                                                   : integer := 0;
			cmu_fpll_silicon_rev                                                         : string  := "20nm5es";
			cmu_fpll_f_max_vco                                                           : string  := "1";
			cmu_fpll_f_min_vco                                                           : string  := "1";
			cmu_fpll_feedback                                                            : string  := "normal";
			cmu_fpll_fpll_cas_out_enable                                                 : string  := "fpll_cas_out_disable";
			cmu_fpll_fpll_hclk_out_enable                                                : string  := "fpll_hclk_out_disable";
			cmu_fpll_fpll_iqtxrxclk_out_enable                                           : string  := "fpll_iqtxrxclk_out_disable";
			cmu_fpll_l_counter                                                           : integer := 1;
			cmu_fpll_m_counter                                                           : integer := 1;
			cmu_fpll_n_counter                                                           : integer := 1;
			cmu_fpll_out_freq_hz                                                         : string  := "0 hz";
			cmu_fpll_out_freq                                                            : string  := "1";
			cmu_fpll_pll_vco_freq_band_0                                                 : string  := "pll_freq_band0";
			cmu_fpll_pll_vco_freq_band_1                                                 : string  := "pll_freq_band0_1";
			cmu_fpll_primary_use                                                         : string  := "tx";
			cmu_fpll_prot_mode                                                           : string  := "basic_tx";
			cmu_fpll_reference_clock_frequency_scratch                                   : string  := "0 hz";
			cmu_fpll_vco_freq_hz                                                         : string  := "0 hz";
			cmu_fpll_vco_freq                                                            : string  := "1";
			cmu_fpll_pll_bw_mode                                                         : string  := "high";
			cmu_fpll_datarate                                                            : string  := "0 bps";
			cmu_fpll_pll_cmu_rstn_value                                                  : string  := "true";
			cmu_fpll_pll_lpf_rstn_value                                                  : string  := "lpf_normal";
			cmu_fpll_pll_ppm_clk0_src                                                    : string  := "ppm_clk0_vss";
			cmu_fpll_pll_ppm_clk1_src                                                    : string  := "ppm_clk1_vss";
			cmu_fpll_pll_rstn_override                                                   : string  := "false";
			cmu_fpll_pll_op_mode                                                         : string  := "false";
			cmu_fpll_pll_optimal                                                         : string  := "true";
			cmu_fpll_is_pa_core                                                          : string  := "false";
			cmu_fpll_pll_powerdown_mode                                                  : string  := "false";
			cmu_fpll_pll_sup_mode                                                        : string  := "user_mode";
			cmu_fpll_pll_c0_pllcout_enable                                               : string  := "false";
			cmu_fpll_pll_c_counter_0                                                     : integer := 1;
			cmu_fpll_pll_c_counter_0_min_tco_enable                                      : string  := "true";
			cmu_fpll_pll_c_counter_0_in_src                                              : string  := "m_cnt_in_src_test_clk";
			cmu_fpll_pll_c_counter_0_ph_mux_prst                                         : integer := 0;
			cmu_fpll_pll_c_counter_0_prst                                                : integer := 1;
			cmu_fpll_pll_c_counter_0_coarse_dly                                          : string  := "0 ps";
			cmu_fpll_pll_c_counter_0_fine_dly                                            : string  := "0 ps";
			cmu_fpll_pll_c1_pllcout_enable                                               : string  := "false";
			cmu_fpll_pll_c_counter_1                                                     : integer := 1;
			cmu_fpll_pll_c_counter_1_min_tco_enable                                      : string  := "true";
			cmu_fpll_pll_c_counter_1_in_src                                              : string  := "m_cnt_in_src_test_clk";
			cmu_fpll_pll_c_counter_1_ph_mux_prst                                         : integer := 0;
			cmu_fpll_pll_c_counter_1_prst                                                : integer := 1;
			cmu_fpll_pll_c_counter_1_coarse_dly                                          : string  := "0 ps";
			cmu_fpll_pll_c_counter_1_fine_dly                                            : string  := "0 ps";
			cmu_fpll_pll_c2_pllcout_enable                                               : string  := "false";
			cmu_fpll_pll_c_counter_2                                                     : integer := 1;
			cmu_fpll_pll_c_counter_2_min_tco_enable                                      : string  := "true";
			cmu_fpll_pll_c_counter_2_in_src                                              : string  := "m_cnt_in_src_test_clk";
			cmu_fpll_pll_c_counter_2_ph_mux_prst                                         : integer := 0;
			cmu_fpll_pll_c_counter_2_prst                                                : integer := 1;
			cmu_fpll_pll_c_counter_2_coarse_dly                                          : string  := "0 ps";
			cmu_fpll_pll_c_counter_2_fine_dly                                            : string  := "0 ps";
			cmu_fpll_pll_c3_pllcout_enable                                               : string  := "false";
			cmu_fpll_pll_c_counter_3                                                     : integer := 1;
			cmu_fpll_pll_c_counter_3_min_tco_enable                                      : string  := "true";
			cmu_fpll_pll_c_counter_3_in_src                                              : string  := "m_cnt_in_src_test_clk";
			cmu_fpll_pll_c_counter_3_ph_mux_prst                                         : integer := 0;
			cmu_fpll_pll_c_counter_3_prst                                                : integer := 1;
			cmu_fpll_pll_c_counter_3_coarse_dly                                          : string  := "0 ps";
			cmu_fpll_pll_c_counter_3_fine_dly                                            : string  := "0 ps";
			cmu_fpll_pll_atb                                                             : string  := "atb_selectdisable";
			cmu_fpll_pll_fbclk_mux_1                                                     : string  := "pll_fbclk_mux_1_glb";
			cmu_fpll_pll_fbclk_mux_2                                                     : string  := "pll_fbclk_mux_2_fb_1";
			cmu_fpll_pll_iqclk_mux_sel                                                   : string  := "power_down";
			cmu_fpll_pll_cp_compensation                                                 : string  := "true";
			cmu_fpll_pll_cp_current_setting                                              : string  := "cp_current_setting0";
			cmu_fpll_pll_cp_testmode                                                     : string  := "cp_normal";
			cmu_fpll_pll_cp_lf_3rd_pole_freq                                             : string  := "lf_3rd_pole_setting0";
			cmu_fpll_pll_lf_cbig                                                         : string  := "lf_cbig_setting0";
			cmu_fpll_pll_cp_lf_order                                                     : string  := "lf_2nd_order";
			cmu_fpll_pll_lf_resistance                                                   : string  := "lf_res_setting0";
			cmu_fpll_pll_lf_ripplecap                                                    : string  := "lf_ripple_enabled_0";
			cmu_fpll_pll_vco_ph0_en                                                      : string  := "false";
			cmu_fpll_pll_vco_ph0_value                                                   : string  := "pll_vco_ph0_vss";
			cmu_fpll_pll_vco_ph1_en                                                      : string  := "false";
			cmu_fpll_pll_vco_ph1_value                                                   : string  := "pll_vco_ph1_vss";
			cmu_fpll_pll_vco_ph2_en                                                      : string  := "false";
			cmu_fpll_pll_vco_ph2_value                                                   : string  := "pll_vco_ph2_vss";
			cmu_fpll_pll_vco_ph3_en                                                      : string  := "false";
			cmu_fpll_pll_vco_ph3_value                                                   : string  := "pll_vco_ph3_vss";
			cmu_fpll_pll_dsm_mode                                                        : string  := "dsm_mode_integer";
			cmu_fpll_pll_dsm_out_sel                                                     : string  := "pll_dsm_disable";
			cmu_fpll_pll_dsm_ecn_bypass                                                  : string  := "false";
			cmu_fpll_pll_dsm_ecn_test_en                                                 : string  := "false";
			cmu_fpll_pll_dsm_fractional_division                                         : string  := "0";
			cmu_fpll_pll_dsm_fractional_value_ready                                      : string  := "pll_k_ready";
			cmu_fpll_pll_l_counter_bypass                                                : string  := "false";
			cmu_fpll_pll_l_counter                                                       : integer := 1;
			cmu_fpll_pll_l_counter_enable                                                : string  := "true";
			cmu_fpll_pll_lock_fltr_cfg                                                   : integer := 1;
			cmu_fpll_pll_lock_fltr_test                                                  : string  := "pll_lock_fltr_nrm";
			cmu_fpll_pll_unlock_fltr_cfg                                                 : integer := 0;
			cmu_fpll_pll_m_counter                                                       : integer := 1;
			cmu_fpll_pll_m_counter_min_tco_enable                                        : string  := "true";
			cmu_fpll_pll_m_counter_in_src                                                : string  := "m_cnt_in_src_test_clk";
			cmu_fpll_pll_n_counter                                                       : integer := 1;
			cmu_fpll_pll_tclk_mux_en                                                     : string  := "false";
			cmu_fpll_pll_tclk_sel                                                        : string  := "pll_tclk_m_src";
			cmu_fpll_pll_dprio_base_addr                                                 : integer := 256;
			cmu_fpll_pll_dprio_broadcast_en                                              : string  := "false";
			cmu_fpll_pll_dprio_cvp_inter_sel                                             : string  := "true";
			cmu_fpll_pll_dprio_force_inter_sel                                           : string  := "false";
			cmu_fpll_pll_dprio_power_iso_en                                              : string  := "true";
			cmu_fpll_pll_dprio_status_select                                             : string  := "dprio_normal_status";
			cmu_fpll_pll_extra_csr                                                       : integer := 0;
			cmu_fpll_pll_nreset_invert                                                   : string  := "false";
			cmu_fpll_pll_ctrl_override_setting                                           : string  := "true";
			cmu_fpll_pll_enable                                                          : string  := "false";
			cmu_fpll_pll_test_enable                                                     : string  := "false";
			cmu_fpll_pll_ctrl_plniotri_override                                          : string  := "false";
			cmu_fpll_pll_vccr_pd_en                                                      : string  := "false";
			cmu_fpll_bw_sel                                                              : string  := "auto";
			cmu_fpll_compensation_mode                                                   : string  := "direct";
			cmu_fpll_duty_cycle_0                                                        : integer := 50;
			cmu_fpll_duty_cycle_1                                                        : integer := 50;
			cmu_fpll_duty_cycle_2                                                        : integer := 50;
			cmu_fpll_duty_cycle_3                                                        : integer := 50;
			cmu_fpll_hssi_output_clock_frequency                                         : string  := "0 ps";
			cmu_fpll_is_cascaded_pll                                                     : string  := "false";
			cmu_fpll_output_clock_frequency_0                                            : string  := "0 ps";
			cmu_fpll_output_clock_frequency_1                                            : string  := "0 ps";
			cmu_fpll_output_clock_frequency_2                                            : string  := "0 ps";
			cmu_fpll_output_clock_frequency_3                                            : string  := "0 ps";
			cmu_fpll_phase_shift_0                                                       : string  := "0 ps";
			cmu_fpll_phase_shift_1                                                       : string  := "0 ps";
			cmu_fpll_phase_shift_2                                                       : string  := "0 ps";
			cmu_fpll_phase_shift_3                                                       : string  := "0 ps";
			cmu_fpll_reference_clock_frequency                                           : string  := "0 ps";
			cmu_fpll_vco_frequency                                                       : string  := "0 ps";
			cmu_fpll_cgb_div                                                             : integer := 1;
			cmu_fpll_pma_width                                                           : integer := 8;
			cmu_fpll_f_out_c3_hz                                                         : string  := "0 hz";
			cmu_fpll_f_out_c1_hz                                                         : string  := "0 hz";
			cmu_fpll_f_out_c0_hz                                                         : string  := "0 hz";
			cmu_fpll_f_out_c2_hz                                                         : string  := "0 hz";
			cmu_fpll_f_out_c3                                                            : string  := "1";
			cmu_fpll_f_out_c1                                                            : string  := "1";
			cmu_fpll_f_out_c0                                                            : string  := "1";
			cmu_fpll_f_out_c2                                                            : string  := "1";
			cmu_fpll_initial_settings                                                    : string  := "true";
			cmu_fpll_m_counter_c2                                                        : integer := 0;
			cmu_fpll_m_counter_c3                                                        : integer := 0;
			cmu_fpll_m_counter_c0                                                        : integer := 0;
			cmu_fpll_m_counter_c1                                                        : integer := 0;
			cmu_fpll_pfd_freq                                                            : string  := "1";
			cmu_fpll_pll_vco_freq_band_0_fix_high                                        : string  := "pll_vco_freq_band_0_fix_high_0";
			cmu_fpll_pll_vco_freq_band_1_fix_high                                        : string  := "pll_vco_freq_band_1_fix_high_0";
			cmu_fpll_xpm_cmu_fpll_core_cal_vco_count_length                              : string  := "sel_8b_count";
			cmu_fpll_xpm_cmu_fpll_core_pfd_pulse_width                                   : string  := "pulse_width_setting0";
			cmu_fpll_pll_vco_freq_band_1_dyn_high_bits                                   : integer := 0;
			cmu_fpll_set_fpll_input_freq_range                                           : integer := 0;
			cmu_fpll_pll_vco_freq_band_0_fix                                             : integer := 1;
			cmu_fpll_pll_vco_freq_band_0_dyn_high_bits                                   : integer := 0;
			cmu_fpll_pll_vco_freq_band_1_fix                                             : integer := 1;
			cmu_fpll_xpm_cmu_fpll_core_xpm_cpvco_fpll_xpm_chgpmplf_fpll_cp_current_boost : string  := "normal_setting";
			cmu_fpll_xpm_cmu_fpll_core_fpll_refclk_source                                : string  := "normal_refclk";
			cmu_fpll_pll_vco_freq_band_0_dyn_low_bits                                    : integer := 0;
			cmu_fpll_pll_vco_freq_band_1_dyn_low_bits                                    : integer := 0;
			cmu_fpll_refclk_select_mux_pll_clk_sel_override                              : string  := "normal";
			cmu_fpll_refclk_select_mux_pll_clk_sel_override_value                        : string  := "select_clk0";
			cmu_fpll_refclk_select_mux_pll_auto_clk_sw_en                                : string  := "false";
			cmu_fpll_refclk_select_mux_pll_clk_loss_edge                                 : string  := "pll_clk_loss_both_edges";
			cmu_fpll_refclk_select_mux_pll_clk_loss_sw_en                                : string  := "false";
			cmu_fpll_refclk_select_mux_pll_clk_sw_dly                                    : integer := 0;
			cmu_fpll_refclk_select_mux_pll_manu_clk_sw_en                                : string  := "false";
			cmu_fpll_refclk_select_mux_pll_sw_refclk_src                                 : string  := "pll_sw_refclk_src_clk_0";
			cmu_fpll_refclk_select_mux_silicon_rev                                       : string  := "20nm5es";
			cmu_fpll_refclk_select_mux_refclk_select0                                    : string  := "ref_iqclk0";
			cmu_fpll_refclk_select_mux_refclk_select1                                    : string  := "ref_iqclk0";
			cmu_fpll_refclk_select_mux_mux0_inclk0_logical_to_physical_mapping           : string  := "ref_iqclk0";
			cmu_fpll_refclk_select_mux_mux0_inclk1_logical_to_physical_mapping           : string  := "ref_iqclk0";
			cmu_fpll_refclk_select_mux_mux0_inclk2_logical_to_physical_mapping           : string  := "ref_iqclk0";
			cmu_fpll_refclk_select_mux_mux0_inclk3_logical_to_physical_mapping           : string  := "ref_iqclk0";
			cmu_fpll_refclk_select_mux_mux0_inclk4_logical_to_physical_mapping           : string  := "ref_iqclk0";
			cmu_fpll_refclk_select_mux_mux1_inclk0_logical_to_physical_mapping           : string  := "ref_iqclk0";
			cmu_fpll_refclk_select_mux_mux1_inclk1_logical_to_physical_mapping           : string  := "ref_iqclk0";
			cmu_fpll_refclk_select_mux_mux1_inclk2_logical_to_physical_mapping           : string  := "ref_iqclk0";
			cmu_fpll_refclk_select_mux_mux1_inclk3_logical_to_physical_mapping           : string  := "ref_iqclk0";
			cmu_fpll_refclk_select_mux_mux1_inclk4_logical_to_physical_mapping           : string  := "ref_iqclk0";
			enable_analog_resets                                                         : integer := 0;
			hip_cal_en                                                                   : string  := "disable";
			cmu_fpll_reconfig_en                                                         : string  := "";
			cmu_fpll_dps_en                                                              : string  := "";
			cmu_fpll_calibration_en                                                      : string  := "";
			cmu_fpll_refclk_freq                                                         : string  := "";
			enable_mcgb                                                                  : integer := 0;
			enable_mcgb_debug_ports_parameters                                           : integer := 0;
			hssi_pma_cgb_master_prot_mode                                                : string  := "";
			hssi_pma_cgb_master_silicon_rev                                              : string  := "";
			hssi_pma_cgb_master_x1_div_m_sel                                             : string  := "";
			hssi_pma_cgb_master_cgb_enable_iqtxrxclk                                     : string  := "";
			hssi_pma_cgb_master_ser_mode                                                 : string  := "";
			hssi_pma_cgb_master_datarate                                                 : string  := "";
			hssi_pma_cgb_master_cgb_power_down                                           : string  := "normal_cgb";
			hssi_pma_cgb_master_observe_cgb_clocks                                       : string  := "observe_nothing";
			hssi_pma_cgb_master_op_mode                                                  : string  := "enabled";
			hssi_pma_cgb_master_tx_ucontrol_reset_pcie                                   : string  := "pcscorehip_controls_mcgb";
			hssi_pma_cgb_master_vccdreg_output                                           : string  := "vccdreg_nominal";
			hssi_pma_cgb_master_input_select                                             : string  := "lcpll_top";
			hssi_pma_cgb_master_input_select_gen3                                        : string  := "unused"
		);
		port (
			pll_refclk0              : in  std_logic                     := 'X';             -- clk
			pll_powerdown            : in  std_logic                     := 'X';             -- pll_powerdown
			pll_locked               : out std_logic;                                        -- pll_locked
			tx_serial_clk            : out std_logic;                                        -- clk
			pll_cal_busy             : out std_logic;                                        -- pll_cal_busy
			mcgb_rst                 : in  std_logic                     := 'X';             -- mcgb_rst
			tx_bonding_clocks        : out std_logic_vector(5 downto 0);                     -- clk
			pll_refclk1              : in  std_logic                     := 'X';             -- clk
			pll_refclk2              : in  std_logic                     := 'X';             -- clk
			pll_refclk3              : in  std_logic                     := 'X';             -- clk
			pll_refclk4              : in  std_logic                     := 'X';             -- clk
			outclk0                  : out std_logic;                                        -- clk
			outclk1                  : out std_logic;                                        -- clk
			outclk2                  : out std_logic;                                        -- clk
			outclk3                  : out std_logic;                                        -- clk
			pll_pcie_clk             : out std_logic;                                        -- pll_pcie_clk
			fpll_to_fpll_cascade_clk : out std_logic;                                        -- clk
			hssi_pll_cascade_clk     : out std_logic;                                        -- clk
			atx_to_fpll_cascade_clk  : in  std_logic                     := 'X';             -- clk
			reconfig_clk0            : in  std_logic                     := 'X';             -- clk
			reconfig_reset0          : in  std_logic                     := 'X';             -- reset
			reconfig_write0          : in  std_logic                     := 'X';             -- write
			reconfig_read0           : in  std_logic                     := 'X';             -- read
			reconfig_address0        : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- address
			reconfig_writedata0      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			reconfig_readdata0       : out std_logic_vector(31 downto 0);                    -- readdata
			reconfig_waitrequest0    : out std_logic;                                        -- waitrequest
			avmm_busy0               : out std_logic;                                        -- avmm_busy0
			hip_cal_done             : out std_logic;                                        -- hip_cal_done
			phase_reset              : in  std_logic                     := 'X';             -- phase_reset
			phase_en                 : in  std_logic                     := 'X';             -- phase_en
			updn                     : in  std_logic                     := 'X';             -- updn
			cntsel                   : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- cntsel
			phase_done               : out std_logic;                                        -- phase_done
			extswitch                : in  std_logic                     := 'X';             -- extswitch
			activeclk                : out std_logic;                                        -- activeclk
			clkbad                   : out std_logic_vector(1 downto 0);                     -- clkbad
			mcgb_aux_clk0            : in  std_logic                     := 'X';             -- tx_serial_clk
			mcgb_aux_clk1            : in  std_logic                     := 'X';             -- tx_serial_clk
			mcgb_aux_clk2            : in  std_logic                     := 'X';             -- tx_serial_clk
			mcgb_serial_clk          : out std_logic;                                        -- clk
			pcie_sw                  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- pcie_sw
			pcie_sw_done             : out std_logic_vector(1 downto 0);                     -- pcie_sw_done
			reconfig_clk1            : in  std_logic                     := 'X';             -- clk
			reconfig_reset1          : in  std_logic                     := 'X';             -- reset
			reconfig_write1          : in  std_logic                     := 'X';             -- write
			reconfig_read1           : in  std_logic                     := 'X';             -- read
			reconfig_address1        : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- address
			reconfig_writedata1      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			reconfig_readdata1       : out std_logic_vector(31 downto 0);                    -- readdata
			reconfig_waitrequest1    : out std_logic;                                        -- waitrequest
			mcgb_cal_busy            : out std_logic;                                        -- mcgb_cal_busy
			mcgb_hip_cal_done        : out std_logic                                         -- hip_cal_done
		);
	end component altera_xcvr_fpll_a10;

	for xcvr_fpll_a10_0 : altera_xcvr_fpll_a10
		use entity mgt_pll_altera_xcvr_fpll_a10_151.altera_xcvr_fpll_a10;
begin

	xcvr_fpll_a10_0 : component altera_xcvr_fpll_a10
		generic map (
			enable_pll_reconfig                                                          => 0,
			rcfg_jtag_enable                                                             => 0,
			rcfg_separate_avmm_busy                                                      => 0,
			dbg_embedded_debug_enable                                                    => 0,
			dbg_capability_reg_enable                                                    => 0,
			dbg_user_identifier                                                          => 0,
			dbg_stat_soft_logic_enable                                                   => 0,
			dbg_ctrl_soft_logic_enable                                                   => 0,
			cmu_fpll_silicon_rev                                                         => "20nm5",
			cmu_fpll_f_max_vco                                                           => "12500000000",
			cmu_fpll_f_min_vco                                                           => "6000000000",
			cmu_fpll_feedback                                                            => "iqtxrxclk",
			cmu_fpll_fpll_cas_out_enable                                                 => "fpll_cas_out_disable",
			cmu_fpll_fpll_hclk_out_enable                                                => "fpll_hclk_out_disable",
			cmu_fpll_fpll_iqtxrxclk_out_enable                                           => "fpll_iqtxrxclk_out_disable",
			cmu_fpll_l_counter                                                           => 2,
			cmu_fpll_m_counter                                                           => 20,
			cmu_fpll_n_counter                                                           => 1,
			cmu_fpll_out_freq_hz                                                         => "0 hz",
			cmu_fpll_out_freq                                                            => "000010001111000011010001100000000000",
			cmu_fpll_pll_vco_freq_band_0                                                 => "pll_freq_band0",
			cmu_fpll_pll_vco_freq_band_1                                                 => "pll_freq_band0_1",
			cmu_fpll_primary_use                                                         => "tx",
			cmu_fpll_prot_mode                                                           => "basic_tx",
			cmu_fpll_reference_clock_frequency_scratch                                   => "0 hz",
			cmu_fpll_vco_freq_hz                                                         => "9600000000",
			cmu_fpll_vco_freq                                                            => "001000111100001101000110000000000000",
			cmu_fpll_pll_bw_mode                                                         => "hi_bw",
			cmu_fpll_datarate                                                            => "4800000000 bps",
			cmu_fpll_pll_cmu_rstn_value                                                  => "true",
			cmu_fpll_pll_lpf_rstn_value                                                  => "lpf_normal",
			cmu_fpll_pll_ppm_clk0_src                                                    => "ppm_clk0_vss",
			cmu_fpll_pll_ppm_clk1_src                                                    => "ppm_clk1_vss",
			cmu_fpll_pll_rstn_override                                                   => "false",
			cmu_fpll_pll_op_mode                                                         => "false",
			cmu_fpll_pll_optimal                                                         => "true",
			cmu_fpll_is_pa_core                                                          => "false",
			cmu_fpll_pll_powerdown_mode                                                  => "false",
			cmu_fpll_pll_sup_mode                                                        => "user_mode",
			cmu_fpll_pll_c0_pllcout_enable                                               => "false",
			cmu_fpll_pll_c_counter_0                                                     => 1,
			cmu_fpll_pll_c_counter_0_min_tco_enable                                      => "false",
			cmu_fpll_pll_c_counter_0_in_src                                              => "m_cnt_in_src_test_clk",
			cmu_fpll_pll_c_counter_0_ph_mux_prst                                         => 0,
			cmu_fpll_pll_c_counter_0_prst                                                => 1,
			cmu_fpll_pll_c_counter_0_coarse_dly                                          => "0 ps",
			cmu_fpll_pll_c_counter_0_fine_dly                                            => "0 ps",
			cmu_fpll_pll_c1_pllcout_enable                                               => "false",
			cmu_fpll_pll_c_counter_1                                                     => 1,
			cmu_fpll_pll_c_counter_1_min_tco_enable                                      => "false",
			cmu_fpll_pll_c_counter_1_in_src                                              => "m_cnt_in_src_test_clk",
			cmu_fpll_pll_c_counter_1_ph_mux_prst                                         => 0,
			cmu_fpll_pll_c_counter_1_prst                                                => 1,
			cmu_fpll_pll_c_counter_1_coarse_dly                                          => "0 ps",
			cmu_fpll_pll_c_counter_1_fine_dly                                            => "0 ps",
			cmu_fpll_pll_c2_pllcout_enable                                               => "false",
			cmu_fpll_pll_c_counter_2                                                     => 1,
			cmu_fpll_pll_c_counter_2_min_tco_enable                                      => "false",
			cmu_fpll_pll_c_counter_2_in_src                                              => "m_cnt_in_src_test_clk",
			cmu_fpll_pll_c_counter_2_ph_mux_prst                                         => 0,
			cmu_fpll_pll_c_counter_2_prst                                                => 1,
			cmu_fpll_pll_c_counter_2_coarse_dly                                          => "0 ps",
			cmu_fpll_pll_c_counter_2_fine_dly                                            => "0 ps",
			cmu_fpll_pll_c3_pllcout_enable                                               => "false",
			cmu_fpll_pll_c_counter_3                                                     => 1,
			cmu_fpll_pll_c_counter_3_min_tco_enable                                      => "false",
			cmu_fpll_pll_c_counter_3_in_src                                              => "m_cnt_in_src_test_clk",
			cmu_fpll_pll_c_counter_3_ph_mux_prst                                         => 0,
			cmu_fpll_pll_c_counter_3_prst                                                => 1,
			cmu_fpll_pll_c_counter_3_coarse_dly                                          => "0 ps",
			cmu_fpll_pll_c_counter_3_fine_dly                                            => "0 ps",
			cmu_fpll_pll_atb                                                             => "atb_selectdisable",
			cmu_fpll_pll_fbclk_mux_1                                                     => "pll_fbclk_mux_1_fbclk_pll",
			cmu_fpll_pll_fbclk_mux_2                                                     => "pll_fbclk_mux_2_fb_1",
			cmu_fpll_pll_iqclk_mux_sel                                                   => "iqtxrxclk0",
			cmu_fpll_pll_cp_compensation                                                 => "true",
			cmu_fpll_pll_cp_current_setting                                              => "cp_current_setting26",
			cmu_fpll_pll_cp_testmode                                                     => "cp_normal",
			cmu_fpll_pll_cp_lf_3rd_pole_freq                                             => "lf_3rd_pole_setting0",
			cmu_fpll_pll_lf_cbig                                                         => "lf_cbig_setting4",
			cmu_fpll_pll_cp_lf_order                                                     => "lf_2nd_order",
			cmu_fpll_pll_lf_resistance                                                   => "lf_res_setting0",
			cmu_fpll_pll_lf_ripplecap                                                    => "lf_no_ripple",
			cmu_fpll_pll_vco_ph0_en                                                      => "true",
			cmu_fpll_pll_vco_ph0_value                                                   => "pll_vco_ph0_vss",
			cmu_fpll_pll_vco_ph1_en                                                      => "false",
			cmu_fpll_pll_vco_ph1_value                                                   => "pll_vco_ph1_vss",
			cmu_fpll_pll_vco_ph2_en                                                      => "false",
			cmu_fpll_pll_vco_ph2_value                                                   => "pll_vco_ph2_vss",
			cmu_fpll_pll_vco_ph3_en                                                      => "false",
			cmu_fpll_pll_vco_ph3_value                                                   => "pll_vco_ph3_vss",
			cmu_fpll_pll_dsm_mode                                                        => "dsm_mode_integer",
			cmu_fpll_pll_dsm_out_sel                                                     => "pll_dsm_disable",
			cmu_fpll_pll_dsm_ecn_bypass                                                  => "false",
			cmu_fpll_pll_dsm_ecn_test_en                                                 => "false",
			cmu_fpll_pll_dsm_fractional_division                                         => "1",
			cmu_fpll_pll_dsm_fractional_value_ready                                      => "pll_k_ready",
			cmu_fpll_pll_l_counter_bypass                                                => "false",
			cmu_fpll_pll_l_counter                                                       => 2,
			cmu_fpll_pll_l_counter_enable                                                => "true",
			cmu_fpll_pll_lock_fltr_cfg                                                   => 25,
			cmu_fpll_pll_lock_fltr_test                                                  => "pll_lock_fltr_nrm",
			cmu_fpll_pll_unlock_fltr_cfg                                                 => 2,
			cmu_fpll_pll_m_counter                                                       => 20,
			cmu_fpll_pll_m_counter_min_tco_enable                                        => "false",
			cmu_fpll_pll_m_counter_in_src                                                => "m_cnt_in_src_ph_mux_clk",
			cmu_fpll_pll_n_counter                                                       => 1,
			cmu_fpll_pll_tclk_mux_en                                                     => "false",
			cmu_fpll_pll_tclk_sel                                                        => "pll_tclk_m_src",
			cmu_fpll_pll_dprio_base_addr                                                 => 256,
			cmu_fpll_pll_dprio_broadcast_en                                              => "false",
			cmu_fpll_pll_dprio_cvp_inter_sel                                             => "false",
			cmu_fpll_pll_dprio_force_inter_sel                                           => "false",
			cmu_fpll_pll_dprio_power_iso_en                                              => "false",
			cmu_fpll_pll_dprio_status_select                                             => "dprio_normal_status",
			cmu_fpll_pll_extra_csr                                                       => 0,
			cmu_fpll_pll_nreset_invert                                                   => "false",
			cmu_fpll_pll_ctrl_override_setting                                           => "true",
			cmu_fpll_pll_enable                                                          => "true",
			cmu_fpll_pll_test_enable                                                     => "false",
			cmu_fpll_pll_ctrl_plniotri_override                                          => "false",
			cmu_fpll_pll_vccr_pd_en                                                      => "true",
			cmu_fpll_bw_sel                                                              => "high",
			cmu_fpll_compensation_mode                                                   => "fpll_bonding",
			cmu_fpll_duty_cycle_0                                                        => 50,
			cmu_fpll_duty_cycle_1                                                        => 50,
			cmu_fpll_duty_cycle_2                                                        => 50,
			cmu_fpll_duty_cycle_3                                                        => 50,
			cmu_fpll_hssi_output_clock_frequency                                         => "2400.0 MHz",
			cmu_fpll_is_cascaded_pll                                                     => "false",
			cmu_fpll_output_clock_frequency_0                                            => "0 ps",
			cmu_fpll_output_clock_frequency_1                                            => "0 ps",
			cmu_fpll_output_clock_frequency_2                                            => "0 ps",
			cmu_fpll_output_clock_frequency_3                                            => "0 ps",
			cmu_fpll_phase_shift_0                                                       => "0 ps",
			cmu_fpll_phase_shift_1                                                       => "0 ps",
			cmu_fpll_phase_shift_2                                                       => "0 ps",
			cmu_fpll_phase_shift_3                                                       => "0 ps",
			cmu_fpll_reference_clock_frequency                                           => "240.0 MHz",
			cmu_fpll_vco_frequency                                                       => "9600.0 MHz",
			cmu_fpll_cgb_div                                                             => 1,
			cmu_fpll_pma_width                                                           => 20,
			cmu_fpll_f_out_c3_hz                                                         => "0 hz",
			cmu_fpll_f_out_c1_hz                                                         => "0 hz",
			cmu_fpll_f_out_c0_hz                                                         => "0 hz",
			cmu_fpll_f_out_c2_hz                                                         => "0 hz",
			cmu_fpll_f_out_c3                                                            => "000000000000000000000000000000000000",
			cmu_fpll_f_out_c1                                                            => "000000000000000000000000000000000000",
			cmu_fpll_f_out_c0                                                            => "000000000000000000000000000000000000",
			cmu_fpll_f_out_c2                                                            => "000000000000000000000000000000000000",
			cmu_fpll_initial_settings                                                    => "true",
			cmu_fpll_m_counter_c2                                                        => 1,
			cmu_fpll_m_counter_c3                                                        => 1,
			cmu_fpll_m_counter_c0                                                        => 1,
			cmu_fpll_m_counter_c1                                                        => 1,
			cmu_fpll_pfd_freq                                                            => "000000001110010011100001110000000000",
			cmu_fpll_pll_vco_freq_band_0_fix_high                                        => "pll_vco_freq_band_0_fix_high_0",
			cmu_fpll_pll_vco_freq_band_1_fix_high                                        => "pll_vco_freq_band_1_fix_high_0",
			cmu_fpll_xpm_cmu_fpll_core_cal_vco_count_length                              => "sel_8b_count",
			cmu_fpll_xpm_cmu_fpll_core_pfd_pulse_width                                   => "pulse_width_setting0",
			cmu_fpll_pll_vco_freq_band_1_dyn_high_bits                                   => 0,
			cmu_fpll_set_fpll_input_freq_range                                           => 0,
			cmu_fpll_pll_vco_freq_band_0_fix                                             => 1,
			cmu_fpll_pll_vco_freq_band_0_dyn_high_bits                                   => 0,
			cmu_fpll_pll_vco_freq_band_1_fix                                             => 1,
			cmu_fpll_xpm_cmu_fpll_core_xpm_cpvco_fpll_xpm_chgpmplf_fpll_cp_current_boost => "normal_setting",
			cmu_fpll_xpm_cmu_fpll_core_fpll_refclk_source                                => "normal_refclk",
			cmu_fpll_pll_vco_freq_band_0_dyn_low_bits                                    => 0,
			cmu_fpll_pll_vco_freq_band_1_dyn_low_bits                                    => 0,
			cmu_fpll_refclk_select_mux_pll_clk_sel_override                              => "normal",
			cmu_fpll_refclk_select_mux_pll_clk_sel_override_value                        => "select_clk0",
			cmu_fpll_refclk_select_mux_pll_auto_clk_sw_en                                => "false",
			cmu_fpll_refclk_select_mux_pll_clk_loss_edge                                 => "pll_clk_loss_both_edges",
			cmu_fpll_refclk_select_mux_pll_clk_loss_sw_en                                => "false",
			cmu_fpll_refclk_select_mux_pll_clk_sw_dly                                    => 0,
			cmu_fpll_refclk_select_mux_pll_manu_clk_sw_en                                => "false",
			cmu_fpll_refclk_select_mux_pll_sw_refclk_src                                 => "pll_sw_refclk_src_clk_0",
			cmu_fpll_refclk_select_mux_silicon_rev                                       => "20nm5es",
			cmu_fpll_refclk_select_mux_refclk_select0                                    => "lvpecl",
			cmu_fpll_refclk_select_mux_refclk_select1                                    => "ref_iqclk0",
			cmu_fpll_refclk_select_mux_mux0_inclk0_logical_to_physical_mapping           => "lvpecl",
			cmu_fpll_refclk_select_mux_mux0_inclk1_logical_to_physical_mapping           => "power_down",
			cmu_fpll_refclk_select_mux_mux0_inclk2_logical_to_physical_mapping           => "power_down",
			cmu_fpll_refclk_select_mux_mux0_inclk3_logical_to_physical_mapping           => "power_down",
			cmu_fpll_refclk_select_mux_mux0_inclk4_logical_to_physical_mapping           => "power_down",
			cmu_fpll_refclk_select_mux_mux1_inclk0_logical_to_physical_mapping           => "lvpecl",
			cmu_fpll_refclk_select_mux_mux1_inclk1_logical_to_physical_mapping           => "power_down",
			cmu_fpll_refclk_select_mux_mux1_inclk2_logical_to_physical_mapping           => "power_down",
			cmu_fpll_refclk_select_mux_mux1_inclk3_logical_to_physical_mapping           => "power_down",
			cmu_fpll_refclk_select_mux_mux1_inclk4_logical_to_physical_mapping           => "power_down",
			enable_analog_resets                                                         => 0,
			hip_cal_en                                                                   => "disable",
			cmu_fpll_reconfig_en                                                         => "0",
			cmu_fpll_dps_en                                                              => "false",
			cmu_fpll_calibration_en                                                      => "enable",
			cmu_fpll_refclk_freq                                                         => "000000001110010011100001110000000000",
			enable_mcgb                                                                  => 1,
			enable_mcgb_debug_ports_parameters                                           => 0,
			hssi_pma_cgb_master_prot_mode                                                => "basic_tx",
			hssi_pma_cgb_master_silicon_rev                                              => "20nm5",
			hssi_pma_cgb_master_x1_div_m_sel                                             => "divbypass",
			hssi_pma_cgb_master_cgb_enable_iqtxrxclk                                     => "enable_iqtxrxclk",
			hssi_pma_cgb_master_ser_mode                                                 => "twenty_bit",
			hssi_pma_cgb_master_datarate                                                 => "4800000000 bps",
			hssi_pma_cgb_master_cgb_power_down                                           => "normal_cgb",
			hssi_pma_cgb_master_observe_cgb_clocks                                       => "observe_nothing",
			hssi_pma_cgb_master_op_mode                                                  => "enabled",
			hssi_pma_cgb_master_tx_ucontrol_reset_pcie                                   => "pcscorehip_controls_mcgb",
			hssi_pma_cgb_master_vccdreg_output                                           => "vccdreg_nominal",
			hssi_pma_cgb_master_input_select                                             => "lcpll_top",
			hssi_pma_cgb_master_input_select_gen3                                        => "unused"
		)
		port map (
			pll_refclk0              => pll_refclk0,                        --       pll_refclk0.clk
			pll_powerdown            => pll_powerdown,                      --     pll_powerdown.pll_powerdown
			pll_locked               => pll_locked,                         --        pll_locked.pll_locked
			tx_serial_clk            => tx_serial_clk,                      --     tx_serial_clk.clk
			pll_cal_busy             => pll_cal_busy,                       --      pll_cal_busy.pll_cal_busy
			mcgb_rst                 => mcgb_rst,                           --          mcgb_rst.mcgb_rst
			tx_bonding_clocks        => tx_bonding_clocks,                  -- tx_bonding_clocks.clk
			pll_refclk1              => '0',                                --       (terminated)
			pll_refclk2              => '0',                                --       (terminated)
			pll_refclk3              => '0',                                --       (terminated)
			pll_refclk4              => '0',                                --       (terminated)
			outclk0                  => open,                               --       (terminated)
			outclk1                  => open,                               --       (terminated)
			outclk2                  => open,                               --       (terminated)
			outclk3                  => open,                               --       (terminated)
			pll_pcie_clk             => open,                               --       (terminated)
			fpll_to_fpll_cascade_clk => open,                               --       (terminated)
			hssi_pll_cascade_clk     => open,                               --       (terminated)
			atx_to_fpll_cascade_clk  => '0',                                --       (terminated)
			reconfig_clk0            => '0',                                --       (terminated)
			reconfig_reset0          => '0',                                --       (terminated)
			reconfig_write0          => '0',                                --       (terminated)
			reconfig_read0           => '0',                                --       (terminated)
			reconfig_address0        => "0000000000",                       --       (terminated)
			reconfig_writedata0      => "00000000000000000000000000000000", --       (terminated)
			reconfig_readdata0       => open,                               --       (terminated)
			reconfig_waitrequest0    => open,                               --       (terminated)
			avmm_busy0               => open,                               --       (terminated)
			hip_cal_done             => open,                               --       (terminated)
			phase_reset              => '0',                                --       (terminated)
			phase_en                 => '0',                                --       (terminated)
			updn                     => '0',                                --       (terminated)
			cntsel                   => "0000",                             --       (terminated)
			phase_done               => open,                               --       (terminated)
			extswitch                => '0',                                --       (terminated)
			activeclk                => open,                               --       (terminated)
			clkbad                   => open,                               --       (terminated)
			mcgb_aux_clk0            => '0',                                --       (terminated)
			mcgb_aux_clk1            => '0',                                --       (terminated)
			mcgb_aux_clk2            => '0',                                --       (terminated)
			mcgb_serial_clk          => open,                               --       (terminated)
			pcie_sw                  => "00",                               --       (terminated)
			pcie_sw_done             => open,                               --       (terminated)
			reconfig_clk1            => '0',                                --       (terminated)
			reconfig_reset1          => '0',                                --       (terminated)
			reconfig_write1          => '0',                                --       (terminated)
			reconfig_read1           => '0',                                --       (terminated)
			reconfig_address1        => "0000000000",                       --       (terminated)
			reconfig_writedata1      => "00000000000000000000000000000000", --       (terminated)
			reconfig_readdata1       => open,                               --       (terminated)
			reconfig_waitrequest1    => open,                               --       (terminated)
			mcgb_cal_busy            => open,                               --       (terminated)
			mcgb_hip_cal_done        => open                                --       (terminated)
		);

end architecture rtl; -- of mgt_pll
