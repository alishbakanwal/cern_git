// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:02:17 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
MFjRGzoeB0GLC/xmGpY81eYqKxL0bbddZyuZId9zU0O71Oxa/q3uxqznecoOxSop
AIxXxFEoPSSNr6wC0KhnTTS3c/KWjsGeUt3lVvn8uKPRQrKLx7+07lgmxFeg9+rQ
ccb8r9xsHWJNZ1WN7G+jJawLMGsWSbgKCA6Jbm7vsZg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 31024)
TnUJM695Hvob9uCV7Ok4/EuH9sC69oCaWiFaWNo1VXo565OSLilttq/vkd/OFhhe
KH4TYJkiKiN0OC5WpMj58CYqowz1ohOGPtMn5L8Be4gVAmCU0hP0tvZzpvKAf9Ge
1wS9/cBqkDRX20EntoSnYGz4FGrJuEnQgiENaQrK8y/4KXcN22N6ULxWpDCWzAQx
VvxuTYMySDNYHqKA7AjTO78nasKO1lTOKGsZypXnCSYc7U+LO2gfPBr2iAF/Wh3u
0mOzc6AtxYec0pV/Vyeaw4mAzkv0hNvh3iJhJP4i/nhrdSWtogyl7DqSlkRZK0D8
xTahE/d9Z4jSsLqg2TbwATGuIzJBwfAvheQk+qZaJzwEF4rwwXlk4TjHqQC4X7jQ
5Ya9ZCvxbpnhOTUXk1V/Et2qRJ+7pvwJWfCN2+LS3Ptvmw/2T1nXWpyvdOgD+tN2
zmoOlHH+oXvqwNpVr6ik+8gRmLZFwGr2s42Q/tmVgxxxHxTbskBM/VMGPxxgX8AZ
9SCyMJl18vaSL913B+fOmL86emYjr40mJ+pllsyBKVg1QFOswQSTwIjQUCO50gtn
k7fOl1JmRZ4GL0aacJt7En1VIV8wpjkfBb3w/DapWcKsA0IOElaK+Dn/lX7JAJsi
gmAZ7yKJnCqI7xv0mvjcUylcddDKcR0BeM7a4UuFDSvsAWta8xJE9V6rLcUK6XAz
Ovd11lqdzFqOwn3VeyZ01Nguj80sw4xM+5AjONizfc1MaqVwCkbpV3fRmJM0ZuCD
iteeLNfEiW/ERQ0L+44tVGkZg5o8lKp+HYcwQGs0M+GLvq3qlu8sQc1VmeGGSnhU
QqdgGXqr+TV8csG4bwvWuDxuCfVwPER7Np0gtlLk2KpfW/LaPTPGlhZ5IhQIwics
rcbLthU8iNzwkQ5f8QEoY7gw/gDUwsJyBBa+mZj6rkUaiWDKbwmTehGJOyICpz56
+0jwxLPhScMd1UDjk1fC8IBYOuv2Dk2Uk3ixT5SFpCXxBxrNosESK5/hQ2Bog4Rm
ZRCaQAj/6iOVKONGc81hkIJxc9NQovkYjnbFqz/H7uPx1Qg8JSGHHQ3Om+rzw2w8
P26HPrWstZbQ+6ChgNo2mf02YisEo6vwZYA5hmscRRSDYfXkEBcQwYPSkcZprVER
sGOrGxrKHB8whf4ZRn848unYaPZabZHp9Gwi3E12AfcaqQhs8rEN2/B0f0ykQyfF
z39timpI8UIs++TgibxhB8MHxaY6dc8uBUfRoUN/w5uFGoXksJvKIFv/igDI2BBH
zyluQZlnh0aSi3KBwLLZjGg1q0CV9KnqCd3pTw7x2z09agJ1MNAsKWqdA9Wc9KIB
VCk0jfy1JFo5fHr8bJzs1sxnKZ7z16xZ9JGHAU6RkBhyhTEhbmhqQzgkfaydU/f1
MYvZPDXZSXClCqQnLfqEJGgh13V8vZVJ74PorKxNrNWroOTtuaQmFdybH5ykKAqH
+uFgM5cQh1JtBJXE8rd1CGisG5BRdXcm9RhPIO9rfrSGyknZFFmYCAi2+kqbay4A
CqElmPB0uhZ+80moaANX4eZGEoYdpt23r2xHW4Y3OTdD8/zEC2wSqZMlJOH4ZSfH
cNDShaEQ7xCWHwU3lo/Hxpgc0VFRnZhwzIYQjoeTlUMrliQXICqBagoCjMX9KEV5
9Z93LxB7tcr4mkX82urBmpIcVkofr1fVrNFYWA7FtQUcY4E6UH2J8WfeiFXnSxe8
sT5JeHFOcDu2+rgGPEzfQUHLUducdU5+6KtIg0piKUbgR53yodqDDfjHXCbvd3re
tgjEZjY35CxnQT2dHWJNdNv62SrHagdO3l+mqhifrq8LqWbJZ/02rq0f5c7QPkeW
wW311FHsKu+6d9xNTGGs+M+H/2aj/c7hjOBu2oRrpqiycTGnstft2sjHAy5PUHqt
IdQnxol81iFmUKtJtuCdrBfzV98Wi3aFOHNC6GJ6gV2umXY/TZqWqnqaDNzMJmTl
2AHpiTNBpyUXYWebuFiYRG3RLcSm2kGLfcR7jnp9XYay2RXCGILk7EZ8mhlOZeH/
ssFh1wWOoDGGO35FPjDFARnvUxW7SJU5+RNy4NHz0ICRzNagvry3/+45xIkpiVFa
nNuxMip+6dH3FvFbZWMTZ1VsowJc08wzvJdTc2o5o0VuKRuvLrpRS7krmgEXKhll
OsXnVZmrqUDpA0Lt0qhI1mWfXeavvdi7QiQKDgArbSs5/rU5oPX8r1JYAMLGiHfp
YaeaMZtb1qGACbtKolMwfmS94tWnfEsd91NbP8RcA2IKJkk0ZMGvDQmF/GsgSKrG
1INbWslKUQKsq5+qd8izkjBnE4iizc9YzWNxSneH4MkFb+46anaEh1CDaTVsEHyO
jnP7PGMuPnryGFCL9XX3MAK1hksiRt8lmb7dkKyaRcUE0ddvQb6nj8mWNtJDHt7c
u7ZnsgJ6hUagg5GBtyL6J236x7TAofbrCyzA83A7blzaJB0Uv/fFc1GIStbwW6ck
WNExTr9xSVhz9x5n/L8mhnAhYmZNcbQUP5UpYgY4guuEZhWCdoKg/VI4SHpMB9BE
t1PC5gWsbtjg810xDV0dFXH5/ypSYsRucukfRNALW2KF8ttniYmiPvcIPdQBw1Lh
f5WnZhicHBDEjH6y5Y2c5pZ1hS4WMRnAofPRiRLs61dt2WCtIRaMkjayAu+4uqR0
ohify0j6G8QkhFR+wM0cCUyZkQcRcG3czY8+yNgZxGy6zQaYHKfEU2bCUgGL0fXL
rSe8ziGGHwk+UU6A8P022DsDyfooXx7WWyy9y5undovb8NX1mlRzL1nt83jIFnah
fOZZ3lSKxVpnXSxYdaqpKo3IfYUcpZEB7qCDsT6niWwQyiiudiCj8Je8Os3zxMQj
0keGmrMIo8Jwz7OV7/dV0xpBN9YgNhfEclJ19teX4lGXPNfDB83PelZ6+3TKo4II
n8RDrfelmJzBAq3cY4HqMNQm3UDp9to4wzAJtlqdo3LG5DdsaAJIF9yIMtD45wnj
nmIj42Zi4z5/SCPPdoLVTm0tCUREJl3xV1JVuoLLkUezEaNs7qTY045nXeDZWn5f
sK4Uwmx1IUxd7VNww0nLLHGt4Kl7eHqYTGo2dJLgjR5zWLDvC3HlOrLSav3n+TeD
KhYi6TxkPi50FseALD0cwrogbxtXCZVwgso8SPjFG0R4g5CJPKuI2VzpZ533zGN+
FPay/NDI79//apaBasMJLr2NEfwoWVMMqEr9hM8yqHzHHhIYgWh1SR28zzh+2Bwi
zJERHY2znTcxzLPCJmd+sEb7FKlEdPtm7pHGuZHX/l/l1IonR4oaksS+ewkQXrG1
1cTET8bHcBIFIZlD+6Oa7RG/8gHODkOpv+xBXkAhD9/L3X1HTAtFEWXYvrADIRFY
dae78P0KG8/ZtDF7g05hGt71z8a8Akhtgwjbq2B3RMv2BY7LuD4Nq2le2W+/JTMU
7lE3+RrKjjNiO7fJdjovX7PMVPBuY5HWeDBRFwWw6tyquzv5MO3nLv8LCWNcunII
EHsyFpcUoMzxeR5hUvu9h4OZK3aV17No6xISxHGinIvkkqAFp2mxc2Ih42VgEMbh
ro+H5/uKwLCSV3qGcaxh43i3b0HNW5BDbdUckw43nTlz8WzV3MEMTPcvIdZyxwNX
REygNcM4gy+ydTcvV2R+7wUUGsqdzyKfp5VPaVdHhuiIGLRsY7P6PJPEQvDvBD3F
aljyHaeIUBW/tnu5SL5v8RLSc+G1AiXZ6d9JUAh6adOnUd0GxyrfpIiHRHWs/6yV
DHBJ2q8luUJrpRmoTsUjaTeyMbgK4JZC0HkdVAdtBmVL+UqKfvaqZ85IqLNoDA1z
PDoABLy6VgZo1pQZKE+JOeMwtKCfktii3k1sBDNteHJchaXYnGoYWCeWOHZYztpK
5tUAMxeQycuozbMoTDZaf/nkl6z31HkB3mIwQu6vje+E8yj/NuoELwXBiLao292t
tx1ykvGQ0bKV24gdNDIyNJs1KQayeHIbXDlg1M7XeYnVRdLDIfcyZuHAlBFYVlgo
KdXuuqvGhRaYL0bkX9vDSgvI/jXZir/C/DtezQck233oW1XqvW4lbiwi7lB+rm3Z
F8lgdhdm2f3EwD9AoKXU8XVrHKfC5zHCtDVZCvBC92VPorqUIDn2B+iFHwB+hujI
MN/fBLWHMy7wMeClc3p9FXCO3BzTW6igk/WSKCh2ABkPDuA8OA/yggz8r5gMErl3
FMNH8fFj6npmQdEq9Y+3vcFjbWPxTVJMdC0xo18/QquQj6HPu4YmdEVK/LiH6v2U
X73N7lB9JU3FmWZVMsSmrDb+ZzNlONSy35Jy7s8DjgVc9gml1Mc1xcutdRE7Mv5P
Y0kHJZA5AbI3xmyWqADNzIDPmym+phAkgoa+AEZJ8KS4HcOCaBxK3tj0a/AzEv6m
BQdNRrvwoa+JNhkHS5SQv91wCtBcR8PtFA5hbBsSLBbskrMnzbILqJX6u9ECTVWg
TFa0Zk69kcm7I34mGegL+e8YvD/EdG1/OrRdYW+rjIWV+FHx6MFziUHG9f/sbuUw
HNE4FkjQqq6XKF9OBbCGNlLnWJWE7sbbsZ+ZqrasjmgQMPBy16Bz9GrpQ0wU4UR8
7BqjRAgc+4e1tUwnil+WAGS4n/nU9AxOea4mXQcXriPEafvlsf69PrGhsJHqgcSb
qH69JULx1OR5pDXG2OtuWhuTU6yrL+cfox4EyE1EFSfI8FJNgBqmivoVgc1IJEtf
SipncFan6dUQAqaVbY7X15DI4GtNOcbVU3zneX33MmblxqoctmIWiHw129JUIlrY
22MBq9fpNjM2zsLKQNfdry8OOnkgjSZ5KBN53fiscJPdlPhp37JQHB6nKz4yOAfg
QLMqxKfJYVy/fIHV2WxOAVC0x6t/owugf3RnOfAtdDj6Wd7l4g/XDV7zMUvZH9kj
uDlqhZL4bVr2YKtnzJWH2+K3hjaYCH9NLpTkDounINCHnTKne9NO9JtGoyVSWxFB
wNqYI8WFPFM6t7uL3odnxy05xcv0PJrxFj5UtD6BgolC02ZF+4eT1dV3FjuDj9FR
0RCnplq4HB+2wGwJrnbwvVXMnWaHW8uBnWtcDIdw+FWlH36+Vi13v4hQNKeIBmH7
k2O7IGDQP8UVNVD944DIEQxsVuliUvXA8xIIxeRsONVuLlOT3FXEZ6Ibl9y5d1Q3
+Jp0dKXdVmgYpVNUcw+Wp4MY99fFFMary42JzjPZKF++aokobhfEEnPd2jNH4m5J
Tjuj/qZrvq6rtKxJJOFp+iOA+ROs4llIQMV4/IUuIrxuLUb7Cz/fxhM0YJJ1c1rN
v/WTBZpIuQoFydzdsK8dAc7d6L29BtxwNaY3YWy3mtk4AmoqoS80Y2yqldvubDZv
WPcz0cpYcIH8x0zFQhtsBBIPDVUqpNc5WEzaWsO9/seLdN/hKAj7Q9vFsBYzRNRs
CJ+DrIGuLCu8KOSLl5EBlDLYn8JFO9XABmVFR7fDvFF4radqHyYG+CNtoSeI3OGa
Qp/glojqVM+Y3j6/5Ex05Ec6nxcvSOR2i7Bxt3jF2FkdvzhHpoflODLjeOqw8WWX
b7awHI2Gtg1qMMgfnIEO27Kz4fVd6NAOgJ6HmxgXwWt5Xv8yTOwpLfp3XwpZXMbs
pApFz68+0Q4spv7JX9NRxaDPZ0uImY2EJZ3MOTAw7Xb7MrjffV8vlwWuJ28+MCxv
3xGEkcqAP12dnesiV2YCu5EifWWPzs/RpXEtVYmedgGCq9+QDXf3vu7+nPrAyUtC
NzyF++C2x002a40V8yS8SlUHG4Zhv8WZj/JuowlsxNGDnnD58wd/AIPVu4gYv++q
trzaZWoXE5Aunb4PmrxREq3/V7M9fC7zXEK43FSeDhJR8cw5t3qOwHAGfAe4/DL1
9POmmKVdOUvOVgJrleZ1VNOtJok3n47qcp2DgRU6NJAJoDlvUyuJmpGyGHmZ8j9Y
5qy4KfEnH+fpTifKJ0KT2e9cfytksO8e2u4PPKDOxnnSYRJLFkBr4HoUPg3WwwNa
srxhfB0au1k92qivvuOG5JkgW7tVpG09bFaFkY3MjB6BPFGp5I7LHEhiDgvClZAn
w6EAaMQXbuV3lpFGZqhIp66szklEFnBegW8GprUex/L4aSXi3It539LT6SCIcOx3
yNrdDZhvh2UeY+ZivyBZobeRjkMA+tjKtiQ8qWed8Jdd0DOvIuu0b+21ISxBQiJJ
SajK9tsZh/oANwn5YHKvooIqIDoNV6txXuR7wuAqAnJN/ZfEUSWWXZ3O54j8sSgd
ePHXSZY3UoWpSrey8uptM08a67OKCjg8rJf76vX63rnO0ZMKDLFiVjuKzoFLB6Cj
BvVPRdaAXNpgfXu4apM2b7lI7dOfwEoi9PglyUVsatOUmrZst5EFSmR5t4+qXfyD
AvEemzu/pczC2uRSIOtHR/Wqxfrlpq7YeF9OQ6F95y9GvrCl4TspGQYgfrySuX7N
XqwPSTo8zcIjWR9At7cWaBbQny5Xx9ONxW/Ccd6my8FCZGHqrSuHgNU6VeNrMNd/
9jUmDpQcRQAH1l65Xu0vJAAHcZOCGe2ORJh275J7tuA1lNJSV6suJqC1ASGTxwE9
F2hsCDbhXOXiV6Tnno4UTB2O4LzwOqOce/I7Kct6mzkBkKJmSe6wGvTWjMPg6Q+R
EJmDIrRckD70o7c6mcY4pbcyHASUqU7h7Jojr2jygW+Gn2YZinRcmCPlGj9Ive5Y
3h7897h3yHYQ0LHuuK48+PtaGLWkn2U4Ogxt0/0fvqtklFSD0MDiVbPPPGTUBRqd
+SCCLVQPB8H6xKmw3+FxnX70S7alWl24KKjM+0G/hcOdMdGXZ7dKDRFuilWFTb1F
lkFmFJUL96zy06N1FHZAi/0HxS8PVNxX8yZTDRWSoYLJY2gzzQx+fhwHrmA95k7o
JQJ5H8mwH6aDnVbCzVvuQdsAP1HYdeF8tnaX5kwI7qFCikSbJk2fGLlGfurfr2hp
ONK0KwdztzEZ6yeO1Y5w81ULiaX0Fi11gbWtVK7PovzMF4rJ842ilbbwe0oequob
NY5ofykXg50hengcST3v0Kt8DgCAntGV8ak5oXoeS11TZD5cbFwRFmf6clxGZ5bx
0e9IHLeRe1DCZCl8II8j/Z7NDcGdsuJLn4Pj7eGv3oDhd89JW2Nf7oBkaEaP2k6c
osW7wDyGWqVAX0GA1CS1NTF5qMtcHXA9IUGzS1vsJ0jPJZ9XtO5CUnyPTXF2qOxw
AWrNyXKBm3gxlm1fwWzTr9EOhLBpZyBL4maObztv9ZVUHYmVLaD296lDn3C7N/pD
vj9WiUFccZ3wL1J3d54syUO3ZSi0OLvviyi2sYU0fIcMBqFhsZrjmMorcubFv3Rc
DhJv0WySuw3q+ajXguWPBx1PCX9KCn9ZPawKzhxcUWGSioeC2Q4f/nqZVbozaJ0I
d53ANADJhg6SrgJm5rifWbeDmnF+ZqW0tMdBTRcyblq+FdCIug+sTCz7hfVCdIUJ
HLCbYxuGXHl/oew7VtFd3GFnkxaYnoddwatj+Brx+sv45W5SQKTbWOIIL1+Bd2U5
1yuQDAYL/Egnyk6zIMgqLCm5YKy2Nf4XaV8WphHAU50y0NXJAytWj+fjotRkUwk3
3FL4/Nog0MFopjuZ1F2mgV9EY1JO6IBjbf4haQsSuleNyrVYXELtCqSxjFSZvR5/
NSUdCh1N8DltmDHtt7g48srQ41tmZV0JXByXj+hviPnvefA/XdDxNrhQB40rYIfc
H2elsG/gN+CRXhnp7al6pHXl/p7a5IacT9lkAJZrR2H+Bt3Q1/uB0ThSE/6cDkBx
6fLC+WDFtHWy7nQZoBi28J1xsgnyTFXJMUpNs3nBNcHbK0obvAOdlDMKYCD7gw5M
CHjSIWjnjevy2CSv60yeUYbiuOpgJ+vWuy1sxLnJiuwHYezez21/ee99hSabIxOv
ZiNl66k1Sjj1B+y4QLrD7gAPKj6L+9+J79fD0UvJ637Xwe3nrlXqXBf9AS3nqYWt
+N9+JnAID3C8xZYB/RIIzAKhiENkK8NWCqj5YkvX+kABOPk04+mIvFPzKMQnwq4o
yCxbtOrYBj4s1g/i3hjME/HZzB9j1czDMGSjSUgQ534vwPs0p7AiyeldI9YGiEX/
z1byovN5dFzdQpRgAmPB81mwQvIeI8zRjJXL6WKel9pCyHYREXv6xi6IL9MJrwua
z0iWNwDCAST7/lis9uHrjpvntpYB8oHGxe8HHnQ3c7LNZc3D8mGsicRZAZiQI1Ly
z88EpF+KjeXUpPNrfli5yHC8FmskDhjUWjcyv4SjQmukC33coyFQmEhTO5x9jCAG
tF1cnc+/VBBslcyu2M/XhAcKmITP42EAA/ZCzjMv6mpg9uPA0nHrzEnLvfEgLXcS
koRg3Jk4g93X1H8iLQG5+7DGuGXqQUa1aGgmAm6507lKJ9Z+LKZJUt2lCZ0NNJZJ
CcyaZ4+lvtxfEiFZS9Zc+XotHydcu1WqUK4gm/f98HhyJFd5iaxnoQtopUjLLqXn
RkTnogUAYSuc5sFGzVRyJt9q5ovclhgPAJa6JfOtvGsSxNqv/DAn/sBo0qr3hN4G
ZgpkKCRv+seSgQlrUbUgxgDGZ7oSgLACsQfT+VGBP694s0u90WPxEsZZzR4BACV7
p1o1/ZPEGcZ+rur9ESVClUWyoXQHlYDTwi4kwx/xEfuPVnxfiIX9YlMHejqrDlgM
AhsP+bHCjysV1ThaF4bpGKuapy92sO1Br4TiNSsMdwsQj706jqP0jhc6+CIo53tb
tbkxY9WYSYgf3ufJUnfFSiZv8Nb01PyWhrL1O5UZKxMpRuy4e4rPm/uqnKEEjK7G
Q1wl/KeVWSJMB2rDROfMUg3nYFU5+2YTYRoQz43Tml5pQS6gWAhXZN8e8RpDMsZs
dBHXee338JRDJq1i4wJQxG30yKpZVUHO7lx9llUibBZpVyYb0+TPxeGXv93jikU1
+oPoFAN5t9x9ODgmj8fqe2tmQP+x6XvyNSpYbcsP/24eDRtMGGemdH8HcxxM+JAz
W8vFZSppN5CJiOh4kCwkGiiysZtWmDijckKj59SD2IpDi84ShSKZol5XjBg0WGNE
UZ6GTBdZr4E11gOZJcLQrjGYSAdqMRP73IgwBzpdWhg8mmIRJhwOU6v+MZ2fhexv
iZbewiKAT9BWkFsvfBYiNuom2uL+wjkctL6WlQr51pcdJc/lyrFqBL7ThnmSfUSC
rsrLMw+WkwFgZwxhmfXLnIo77Lnw1gbgWVBzRCVCYLGME+gVvtD6a1MlTMD5HoSp
pDAPyNJhjsfbWw9A0ihKrsCinMD95XJ7esQzIShNe5VtlT9H1JT/j1RddtmsQ9B+
p8jx+a8hn6hpOVgUuJ+GfSNdc9y8AnSP28rYFhq1YXmHc6hJWUqnD9NBN+e7x9fe
2bWwB64cFLckPtKnFNn46nP0+G1xpavt4lcn83gJm/ekru/6H84BXZEpdf5+RM+2
QY03Xayqcu9cLLXAaixO6yfaFIzptoWb6MtQGo47xi6FvNLFlWRdpqc8M9Wowcg6
BYAG3O4QGqtvwBILZDA89tEO8kF2Qoof+WRqdRmirFHy/X/zIwIy8qaxUhsAuYco
Kpzvd/BWtstyVpVve+68WaT2yXh903lyCzH7avU/DF2XVsjiMbM69+KW1L+TfpLn
57qepnbPuCYbNFbQwjRERwWfhCMXW9e7Gj7mw8ylglqArWOrLXznlG1aakm5XQIT
cgHr/2In4IFiTb+HIqTrUXCPn5Z9jXYmnaypRtOvByhdI5qph8237sZZYZfheXYQ
Xh1kTaJJXDS1IQzgBdeWh5798jFsby1/AH2FhxuAcZdzvGThQFwMHNNvm5Dn48CK
VXmyZMyBnDb4F7OMUnW/VlY9MK4jfJTgHWeWxOgbOy7/u4nq5bvhNXi98lrtlbxJ
AADOk4dX/rDAFW4VbLnkFUXI28BpGE69cET7jTIAawXfqsBttBlQrMRjambwVNjn
xxhnJKQyg/w+Gl14DCzZDdGcKfnao2q7Y5j/xKRRFakBFAiYQniUw7kKDSmfR9LY
87H2u37XEkbas0xV60VNcUjBFtwHOc5KH1Rsq8HlL8/QL7oECiXBG7iwT7dDqf5S
FRT2KXO9gFiSMAOLFFiPjaq1qqW3vhQTDx7xnhZQqpoegoaor7jq6d/zEcZoWYF1
rKuQBCudVKTG7N2ztqbsFd8U31KcCFdjZj1oBcuJLDSEp021w1FWebW45gtyIcq0
LAqwSsSzz0J91h8Vx4motiZC8OjzDItbQCNg/38LxZ+Urh2S5kw3EoyOoV+OmsQP
MQ97HhmaFlOpU6LjihL0Ozca4Dwx1IfCmfrlLUj+p7jfe1EtZeBFPbuBlK4fL67j
3XPU/bFYgiI8x1cSVLlo9TC85MMMFb86TbAv1UfyKTt92E3LFiGHsfqQcE44lYbM
pm25N0UoQlLpl0O3fSDXGNyV865DHbQpcjRFK2Iuu7GpFtESRsw6ZdjPaZXSiOtS
iu465jVzoM9UfIFRE37SqQsvP2FtK7sNppCY7trP87pdRY9CVNN87kHZ9+EwBACU
naHa8s6UM9NJyUQbDv3b8CGAPqfF5g9+e5UgZlZFzIdYh7qiqK/C52eKjyLrRDfg
0C/OkrPibm95fBcLzm8ElgWeYnDlGF2Aw710H9/7Tg/makabHPxEknXRCO8mO/2k
mA8AMPcZmw5q2+iNq7uprGNMMD46SpS1ClN6cFrIzgCm5rpEer6iXIY3t+w48Od+
BR3FzIhAGIk+MLMpeoOyEss7S+ODHun8SxYsVUNB7W9Fel0GSUs9bfwn9p9qnbS9
uXF30ZJAjeXBuDfyVWdqc6Vl7kemcvufTdOxZ3gUgAN3TlzD43mOcy1aOKP/ZAMF
7rd8/mHohT3GQJAppvrSXxck6VjZrVIsPHmV0DmajzLJjPrPqV5iWZ9ngfuOgDik
EwCqpf1tuVJYlIZRcPj8IlB0aWYNmoxcQ/F31UOdxTaBfS1lLHAlLVpxv/81/ORC
b+fIb2QmD5wEJ0uhgozadHZXXehRKe5KMFD2eyodpW/xFh7tgRhJYh0OIckPL14n
QEOtp6Ju77hgGH1n7GIMNeZvDEv1G9E5SzK9c36+mpwpTrvKAMQfYj1muQsbkB2A
D8c+HFqj/tdVMmQKwZXLO7R1lCmxN0Adqq1CsIRTLQbdLPcLAFeyB5lQ2naY7ykf
rPT96G/QY0bxWJ4PnrzMHxFZ9Hdb5KbW3fn1YWi23HdwfC7tCHQ87goOSB08yxh4
+QbxHSBveVADZHSfCAfChcLmCQg1X1QSFA7qNDT+G/Xm2v8lHtKjz8uq4rmZ7O80
ZUJIC/MjQgt3dzzbXdLgcCGDnel9hFzwiAQbVeTYPfOH9kkVC5Sk0gVKR8uxlgtL
9XqwScvQdyh/qMwHMe9hEGXxQuSkI+a4NX7bcr9hprzUlaHFXVIOZao3SP1kOGeY
X1Fu80QXLEV36xcC/PTopFviCgZ1S1y+u3hZQlubIGs96wLRmnvNGN+K7z7+ioZg
TSqRxTdAQK28Hy0Mw7mSHsEgGaytIKkVMPQx6kIkxXlY5VP1tS6odCReFq3RMiY9
QTwoy7F4PfPh6lKwf6uin5K1OJ0TNOQpNQ8sZf7bs676GKUsQGEsHqq/rtDnPxld
EcjihGknz3PF9Y4EQovF/dINzL+vCO+cvrk83c0xohycM1QKdGG8qJ7wqAeK3iFO
HVw/38pgIx2helesLfMtCQ5oGH5rde0cZlUTxJmyuH63OJ/S1rOOQfNm3ek6IRoC
uT2ZCmamTf97Z0AcD1ppToqN7QQTyBHBRb8avftE3mOZhR32+AFXgsuWoLfcZFVl
7D5T/ap0mH6lUmwc/lKn4y49reT10i476WeSM6Qt0Dja3TvJQVSZnTa9oq8TA/rH
MxlTrRmm11F192vCeWjnMKUR8k1FuE/TUKEPfXxAn2amm3hRLKqL/Ty/Dqkqp4Zz
kLWf65lkoAbPpWAxUm7qvCOiZCMjQAzbU8C3PUX5zMq77sK+BBKiwCd7D+EI/Bho
0vcV2liboAaGMAE19QVe6B5xhlPFXaB/qnRKdNqy2z6D9iSaDToYhH72CxKggq+m
agncp0gmp3bMgN9nlIu9pB9pLSRNP02DI+H1XEzvPkECgsKlVmeM5Ah2BRJMAZQX
8Jtq8FNPNkSaSHKd1W7D97RHbx5gfymiMcaYWhFfye+h2jWF5jY/kG1Njnl49Wab
+QixjND+t/eCxWj66cIAJAhC9sd7C2NHBULZHhoOOokYLFZ83raZrMHCJvEN8H+6
e7wl80wKnabVs8ZXKPDGFxPQTLYI7tjctNMjX5W95Rxt+TOLfzjnPun4nP2Q2BxC
kA9xWV2+aLDOboOTySQnXXFw58KRINKPS1nnjIuBhNCfyQ8AzPDP6UmTlBQqkZm5
coIfRSvg4uPnrN9/SSdzU4EgBnsjNwjwAWNw5kYRT84Lgse0gf4Ezwvzl+vOcDvB
k5FSAtQDBefz8OQTYu9gkQZek/aOD0F3SaDwrY9xoZgdwDUO6zuUC/HyJfAg/xGA
yBW6xj7XRxuwArfWAFL790cku9OB7/8py0gVvu+nReEXpsjrhHH75VXSQdJnswVY
tkwn/sG5EUOKOMNZnYeBiIdbj6UTKcSB5z32ec7GINxOUlprWivuLadSReMtD+KY
m/9uCa2lU0KaZhEY0z0sbUm4x4RX4nyCTWXE4yThzSO0yLMakxFEAk8N2U1gSwbY
HX0op0RDxZFca+62eTNfWOfiNhZbkKcqq+b9AltDxrepeHCyXbBl4E6Lt/qFM1FH
PXIWu48EKTgb+JdgZsApxgzfVtHcFSPk9wRFLKVACqeVWfbITwbKtJYRXPvlXtj9
cmA7c8ppvujda03/Bzh42wy3TSzIJ0T3e9Vh41T2kOsnxgpSqKxCTGRKZPT3hzNZ
y0gO7dpyZ8uM1fMU0dpdjCzJeNK0EbLfz/oN4b5D3zino20WXscuG54DuxyPO6d/
OZWHaIYebAcPlbctK7D5oxJMv945/shaCjQNvWk3QEyB/C3i5ob3AOYzYnqti9LM
0UWjHoQVXg2ypJtCqqCNB/sTL2VXvic3EEaLjRO/sr1HU/oAbYw7QjPySzLkSNWw
FQ3teAn01FwBrnMsWKsGk9uSal6b5H7sGo2lXcEtgiBDCxXHzLxf2cGHqLgTDpBd
ZDqQ16d6x3nZU3vRPnSy9mPZ0qfFIzcyEUT5yLJvaovd286DKcJraxk9MRJS5Opp
iJZpqsjNK5cbzBFft+Kw7tJ0V6ZFCqGmKB1OmfF/MEcM/dVvc6f4SOXROXjqARA+
3p72JAOUNxYTTLASJTmGd4FOzS73QK7QQKwF/jTrUL1bvV5Ge+NZIM8RvdZnF01+
0kIIf6/v7uYHdWIDGgM5hn4MNhXmbTeumOui0c/GMyv6CBZT9YJlaGta5G2rbEOi
mf9NpRszSur4kYcrmC6EHIiQEam0khou/xZd0yRYSVvs1mGwevpxQMMSt6HuWE9Y
kfWMYxCg9f3qZ/vx3GWkx1wlwVvZsQQth5oV2CuarO6Da3dsdnyxdJCwYETYsW8o
+yiryCmvYmnUM+yVRPVbQafQZNB7u6+tzJWs65N6RXctNW+lSXEOaRpsxA7QBfAS
ciRo46Yc/kXsFLWNOn1gc63ZqfTVksoF6csnXfvn4khE5jAmkCaK1RX9yzqVa0DI
CveK9EOkOljea1HBEfLCQWhCGRU7WL+SZaKsLQPNM/KcGyeMye9JEih+FdQ8seuX
KkP7NMEPxPkbzP1XpwF2WpW+yT8qm+W0QNMsNOjpTopF+a5dqZo4wWkQ6sd84LWY
FzmVKJSZZw4+VDxP7oFLw4rSkLYkKRPeRtY9i+8lxx4lvrpZcTGQNw4wwhXm61SI
Yhc5fiehg8D2rLiTMCq3kFS5AuX8hqGJGbiINdkTs6Z0xwT4NDaB2Xgdj32skjLL
8sUlzrTAPNNo4cRoQ5awmJuBY7YL8tTwgV1Xbh4R+GP7v3d7eAoRsoX6mrHsLK1V
goYUfKQyEFAJSJ2SoDopIpqdzicR6hjASa8FU47jy9I9dUTPPSvXu3IbVKU4lHhO
eT5F9cAnzxzbQwdGDwr/heWkPvwZTHVO7lmcraHRJmqc9s/jzOBmANJg/3RrxXEZ
ZJE8h5c211/RcawLRYYdw+O6bi4X7Olg4u+4DFbk5X5DTlW+uVil4i+8a1bIzweP
NC2gCyfsXe4ykJ/gBG0JGCVzjmYHP6Aj8o/uJJaAXd8hGjz8PP0VDKkK3L+H5I4Z
voiX53oh11saUhSucKwp3gQfZikK21cY/VPq/Fu+rnmnr3u1fc3oFcwLv2SnhjQx
EmB+2Rc8uYvfHXtU572+YN8WY6qIRNqJeadGvOcw6yDXbGUYC5E729y0KJewy6+D
GdCdeYefYQ3I51b6N7r3+I78GMEREuQYDaFw8BDjjV1+Q0LFtqRwVpMjfQ8bDu27
Cwm4nGn1hPCKifHDF3YhBgJ6d5Amh0PLX+ZsxflSCTA1egXaR6ZMYrJ+JggfveDb
tKiW/PG+mCsW9KsissHSW3dmBbztt7R9U+M9B/cm8UwJVDslngMKI2dcViP1KplH
w7EqEO2w7sYcdn9viUSYyc3TJ1dTjLavz7DaDMO1A08rhZ8gsUJ+JkAtVO7qvpq5
RsFmIt1ITtHnd87MHzRe4dlQSbdZelxKu/hq222qOB0rE4mKtPuOaLD+iThy8muN
N49BhygbFlpL2uDzrChzrnpBRI0sjMW30i9deiqOPTldE/hvW5CkKjVijTP2rlxX
mPMrrkDhvTCUTSoBUXCWMTJ0VmW6HGYQrlYqmAGktH5wwut9D9QTbmNtNlyWSbVw
3CsbljIAucQic6u18llUohybr8TpIyQ2YypcsHlz649Y3dkA3q9bIJCd+hEBeVFY
D1EijkZdEP2NRXtVZaaRBeMspq/sqCAD0bRm5qjVy9977gnAnxyDXuSd36NQZZlu
Qe3jIz/VnZa7aAb+H3NFjKpuKyAjBqlKqsDMssnW/SRZrMkDNQEScPZM1Yl+ukHE
qR9zcRUc4LZHhqBhYWQr234zm1i+aXKede66owmr59NpuHQtNuJ2rb2bhtN2rZ2o
O1WLF31HLSUPPNp7wXREfcGH/qn/j5/6mO+0zcmB/DhRg6qwMWgDxEc4OvWID8HX
VDDktCPuazFmltfWmtoVDrqTNj5G1uSTrLlr+FQrU9WGrMVqm/GJ6xSnhZ3dLMI4
afGSjoeaV7dRngaxMfO4pVDCNg6pAD72Zhc2cSAUcG9CG6KhPIqkdIiSv/uFQR/E
tiEeD0jFKw8mDfzyFj4Gf7c3BOEPT7h/P9fKYxHOA4RIbkkgtqjAwQPEjs1U1K55
alQUQU1KrWi3HTgWuM63Whhg7Lyk4JAP8FEk52LrRAVDs1l3YU1X80AC04j4HEKC
VXJLcDFe8vatG2jj36YqsxPa84DxIU8Xh3XIQGkmAzdN+GquzuyZEhuVtJhNFa/L
nlOYBAiPh4IvuIt065NQHuDPeLWJJsYjHqH1VrPFQ9G47NX3wkp4WzTDJ0mrMhvM
0ox4sAhO1JIHL9XivK0Rf5Y6jzp2mixntZJ17LPG6H7OF9/ZWVaiHBQojYCfSw3v
5StYA92PuGmcz3rAF/jpYE9t6hy7UnwOI+0iD7KqMc8XCCDZKTOC8a/MWGGv+2FK
WrgCGvJ0xvw+UGOg1kJvO8g3NFyEnXOs9WqPDpDqEyJXzB18LRCWQ2Ia48NHwuD7
TgYxAaHZ8jXpQLoYJbg12Yt9mczobo5792sIHhvLeh7wTMtVNF7XMEiOVSWC4C3m
O8lMYmX1pvtPLDJ0fFvJ7P+PPp/qr2gVe27VR8+gxg66BZzwmKwNN4fLEq+dZXKm
MNcmNZ8OT3JDpwFh5kW/SsqD49YH0uRenoev8nPmbw5ureti0qY4R6k9AiIHh31P
rjZ6ySc3+B+Qy0jtBBYKO6/7iGcUZ5uDYQX0Ix2yQybSPjsmE6MQBGKPMVeyOBmk
V4Ivt0jtf6Fa98BVbxkSCeJhny8uQskbbA+ZuswFeKHkRrwZhFAiQkoIhbig1W1O
ABGepbSGWDVlBqLom8KSHevFe7rQW//jbV1EeErMeDMovHiHTe6oTjBrGi+DPzfw
a+I3W9U++YvBa8cX4R0ctWzZZuiVgPUjCQ4BzbTQiEqAbFjvE+MNH3kigiwFXjn2
acl/hJHdJI2aZ+ss6n4H2tjFiJbDyKhPFnJUCb6hiXwu0PFimtVHb+ssIrCT4TnF
OBN42OBn5sOd1c2NE3kr653TrPUB8loa6ld6uclBOYfnfrPOKZdMYNwlVSQvCG7w
h2vP2p19PYKHwQ8px9O5SQVU/VBdDXAuKPSU7PCmAu8+l+LyOMeFlXQnJagT/j2x
VqdmKzNGo8LNIquTkjqy7bxmEypisiwrhi1ffa67Yybn6cRIVLKNX5BeN7FUjOMB
MxWude21bRJGrccgQGkzixXEjnZKLM+NQrx5eVf+R7LX1z+lQONxJz3nbx0W7BD3
qRv0ayq5Q4nTntPAKe3ozmunZlp3j0H+bYK2ctea6+IcUTy6mVVsO7jGgBJzMfMJ
9eEGVGsb69MN/rQA1I1RKdLzbGZIu+S4l6zWnJNPGwY66IzkYxWN14XX4m6U/aTX
sOHsAW7kOYkm7JMQcfF5p30waR+bRU0mz8fFFJqJZXEXTcpwDHdxZvtLBG1q2BEe
CBFi/V2z2an6MCQt3fVlptaJMrDSv0poy6IGyRg1+VUVAlbYHbTOq+O79woER0hj
kLj+5LUuyLgQLVCl8m0PxjQeFm3z/COJ2fsgAAeGgtKhIjDFY178TtWC/JQbC7X3
8x2dy219Keun3tcKPO8lkscYzIRJtA4NU30FUy0zggLiDnfoW6K2Phm1ILgQTQbR
1WGG/AFnsHztdhsPBF3QCySOVm6oAMWvF0FfWBiU/X61S7aP0Z3yJEVp7qdUmAF4
da2pRh5vRUZp5aFbWcgmYFvggeBEv5rUnsyKQMdwaa8ATwK3R0+mIVU4zXvDTdXB
GvJjVG7Odfofw3X73c43RK5QIs0NSa6KJauxJ/8ZbJoTBUeKS8tIP+Qzl0NKNesY
bSfdwKf7+i1X7W4Z0mSURxtQV9QSYQpdiR4W1kLEmgL6sWJvRevD/AWtCglXEPh1
XnF0YVuNGDI1hTTXBKprscuvMEvsNlQs8EQ40TWit8WaBhutCjN5Sybzf2Gp+1jB
njiv2tK95PYHVwyYeSUIRFtIjcuq+iJMDolkp4npVpth50qi6HJ0OXrKbK5weGE5
WZAcUdLvHsf/VZWi/sIfbCX30q04++lvSkXZq8C1vhOUMlSQ4GF2ZVeglTDh195i
oS8S7SkXU8xNFMJyXR0MBAqGIaAUH6MatOGqYGBUlrHJieBhO1qImCiG/AVqjRkB
SkxyhRenPgR7Nzhqc1dNg2qoBrVhPMTv6MfrhPDbKMMxmjITSLdD3vqeWRDLtL4D
WlFDxBjG1asBfnURxD0nQhSaZh1SKgQPDTbOzd23dQXg+GNNM+3O++Tu2FevcNHy
IwS0nqrmY2or4mRHf/ypT7rqsCl/7Wv4CAYHMYY/kdc/NtbN3AE1/nzNbcn25Pbq
dr8dpTdYXJNBhPJzr3Pp6UsV9GmLO/KVKn8NeAr6NIZKRnj9bCOI5nXNUVPQi/Wr
3q3iuHaYeab/3epNbVkOJEMhBeG+wvAVKPLaA8j6A86XBq/dlbS7WtdQS2r4pj7e
OPjgXlEtnqsQKss1uaqCPOLQfxbqJzFzUEL23B6EvAI6G7II6IXNsPiVCfJe/FuH
c1KOqfzqR6nNrWgVzW5FVYaCCypvMlI6/PqXC4FMOZpVCNIEc2jf6J2Zd+dO4xd0
RPvl3rV7EhLO7kcTp9QG2FWW9El15B60I17qskOrZmd1ugtwb4h2/aeHRJodAdg9
4hf2U8gDT+WupLp89waUDmLsYAtEEq0Gjd3Nt3KhoHobat0M3IvqKt9YUbwB6bfG
QW0tU/ffR30RgwX55hk0PdMUV9fAVdC3RNr6NSUAVoA8qdcZr1laeSUU3/pNy6mK
P1WhysJFes88E8TciW1VhzdrMvPFTVqLvqAkSlYb8ljvqNuaMNiy+RxYm6XcOc+T
jOYnngtmbSGRC2Vnv7h60EigBEn3J0FaXWi9TocYeuHvQIUwR7QFcy47AATkrX4S
/QYeZVawHRUzgY18cH0sNYCgFkJhU8evXZeGhePphAt1di9kexj2qdwix2tYRyq6
+0F8XQub/Z2s3TKdtJdPyZs6uLBWkvnvil1wBmz7Q+vbzn3aw2vLqWYXFI7mwXVF
uBlBw6gk4d84ZmIyX826Ul7I+Dskw6NPq1c/OQpo/3j8wgXwrWfNtj0dDOx+zWXB
sOLpwpd2wQ8cYTNaZc5GB/RJACo6Y4jI5djRzNqkkwGdS+hinHrwkyTwVWM+9mXG
6Ou++g4B0ge14vVejGxf313LmWTxyDS9tQdjsvTmLu84XB6lfbr/Fc8tbfCDW1Aw
Dk1Y86VeY5AAYFOnJkDW97+C8N4VAuALJ7Xgv+nF4s0COlKC9512sPywIr8HBkJ4
zeKrTZLnpFVz4lUcT8rp2fg5oxbkfjexeLn+4n9FSKJMwr3+U+o6/7Km3qt3IdRR
lxko9FGx9WCXtl3Fw/MJ4gKk0z8vXGHzEDFfin6L7RFVtIE/UIYT0sr/33msyGZI
nlBcmVHOq2PznsETjDQeeQ44XT5WEFjzzuDkwM9uNWX/z5/wuffmkfMmaaZlohNE
71YrNWT74U3gbSxjR11GpGNhriWLEw+zaefBvpOz/sX/nYy0CfdAi3BcNiFmZrUw
RSjcifpBq1dVJv/cVe15IW8tYPxdpLpPzK2wJgqglJvljvF+/iyFKgDDY70Aj/zS
bteoLbzT8wkEo6sI18VyO+jrk4xrMdCL4Rt3qfJxd/WvByjFGpEn1N/2nEE7QiKt
yl/vAOB633LP10enQ7GXOEnM7KWOmS/lDX0+gAqrbD/gt6uMO31Fy9G4UUbjp0Rb
x259y1+5fXjo44fOfyuBCNUU2MqPeicq6WoWQn2QLEIG3CGcRKoozRMnPdqpNFuB
GqHaepUUjGd9BXbatPfI2vu8MIlt5El6X9nE0amAs3QmpC8ceQxCZPtlHeNkyoCi
uWAi6jjLgSO6elCiYA6a4CS07EQGr0ItnYQ0bfvONjR9QIhS/pJlGSS2Jra98F0/
+4nwM3pfSKZZ/K8kNHkKRFUJbBYNPXDXr/bntDXXbm6Go44YxnZHWwPRr8Ow8eq+
LM+g9xbKgonOfwsRfBLPs5eL0BgSfYrtdJP0cEx+Vf4hmvCBi89U7Zz1caJAzIbn
16jkmKOi7aFvIamvb+GA26st0usQ6jig/w45PH3Ki+qfEJVP/R/wKX4AAZqvTGjy
6jS1gvowzWmIe2DKba8reGn8b6HPT+ikx33KsiVM+YXzfY8hG8LI5hIZ4Aq1PXiu
nCO88ph1ouiK6Uez/A1JZlJVjXqOC5Mc/G7TnTBQs13T0UX2rYK/m6SZ9Dq1lwo7
xkjXaXU2aipM5p++W1GmO+pk9hfD4O37klUngjrfpnqW/iUw88ktfx4mvPRU4Umf
BJzcAnO8ZJLV773Vkp140ucY7vtfzAddjFtdJ/mZXFQrzJwt7z4Y5YudG3R14xSP
FIYo7/P56+gTM408HqoQT8ggsVUENlKE7N9Uir8GzUqxnpA4XBFUVh3hO6YX2PoV
+6ILEEALEXy03vgEg0siflWLv60XNEAoLEq79+Hc0Zoy7xSvkvmp5j63qaGb0sAp
78pQSmLiw88wg9lyBn1ZMhSME9NOwhGE/NzbL5yuOf0hgESBfcmE92LKRglVnxu+
6FeS3NCLvOWcQiD5GszRTy6Rx2588AdvYJQZnTzI7m1OISXuRJeAhODdVr2QQUzL
cC87JQM2t8fqWrZP5nKZU9XaELjBQMaeNjjwTEaK9MgCvpDLUD+yxI9BkOba2HTv
LnLfs8NIlgZS7udAV2QEsjmasjdszeshDfV+wM64Q/WfBF73yl8R9f3oChcZpY/C
g8nQtzDfnShG3UyxGzi+2N2FVln63FwhflR1eA9RamDkfbjVXyxJkuUqf0Cc0g51
9iCV5Rb9l3OizI2OkrHMZGLJ7olcfCsY8ZpxtVOGYDg8HFq2kCXHcpwpXQs3lVsU
+l0ibesif9yP0kQFg8iHDcyrLdKrMmn/Rm8RXT6uVp987BbzQaKlGjMfUP8uEqO9
TjrUxdD9Ao1LAO+dRMIk0OUYmYGeVVBr2gYddJIky6KGN+D53JXkzeZybon+leKK
uGP49wSpZWmJW5CnuUqXRGlC1JaApn1OJPj0ML8XVyTZBA0MRNA5qJzQ529c4bc6
/sTbje9ahAVy7Z4hDJXFTQ4nWcQFAb/YRvIKQ6fQCVQEyY8Ec43AY5m6DNRNlXjV
7/HAFwm/L1ASRl4GYwD9Y1wD6p7ubkVPcp1w2PXzWbaHjvWqGfEAa57RgNQLyAg8
Umi6ABYZ9KnKE3PrcucaEWgkO8rPPdiXj4yQ62V535gOATcxXccxeb7Kbu6hu9MT
sQO7RQbMF8Oh9qp53Bu12ljEoa+AvmyXd4hkbsVWDCB2BPKwLrsEPubZiWA7Y+r3
XlnJK/ll7kwF/4tvnCTGfPrKszVcbAPwX3wCMUavzTDgSi1xCndCpPmKt2heGuST
QfkuLdCSFA55v3AQeG5Wy1fNEWdE1ltY1PROBLqZUq6Xa9m8nORGMdIPZQLZ59ro
3+jz7gu1pBEVQOJIwyFGmObmZVsF0Vx8o4gzkczbEyeFJbo6jtpMFdUaXsYN9Kv2
/RVJWuHDf1s2qFeOsv7qbHJwiLy3nXrmBSdT2Z+2wdor1E0BqoaipIq3PYcjRXLp
8DG0/3whfUGJHvlvucyYAZ6ACeVUFkDQ07v3dWdMlTE4v9lpkgJ8iIrl2OUP734J
LZ4FG5ZWx2nKZ5t0qDrPF83guFy2tJIWASQ3Ipkp3fI8OMXBUW3H+taMOTgt06nR
g8dOfml6MtmUr5308Dv3mYrsKoTuUqyVwAGafIUWNmcVUF6LVj4Q67JKNrlXEeO9
ChrZwe9hJBo/eKdC0sYsRHaZDq4HHLhk2viRWK35zyJhK5+rYXV8pGynBkmL2CAx
MU0X2lTK/QX9KmnolLPEWjFileAdfn4HaMwMJ2Cr/BwqVUqxYIvwuoRfHKsvboGD
pdccA51K1nKuG2m5IKHprUOWCGp059g9AIwJlJEZR6MOTErUbQY10i4b5KNTq/UL
wXFezF8/fgFGyKnTp51IorHTlTbBQx2kSn/w/Akd5bCwElg5vBXLn+TcAIVV3Ilu
FeN9GJBULLOZtRcVP+43eqzhI+GvZrSgmvga4cBAEc2X+ZuWLlUXgPnZnovkXxCk
1sWyby1yhhE6oQW9ETY3H0SxrqOFmh4y2SB2MmywLh29FNmLVD+CL5RVBPqLYJZ/
JRm7lgX7NT8seAm1OERPy30e7vMpWcTwXFjIM4THu75HA6jbrhdWOa8l+Cm+k1p/
pzGySkfEHI08gyCCCWF9Y1SAkHBZnPb6Udx/9+hEBFNWZ9rL7QGstRkIM0VkQGRK
3yrx5i6JMs7dIV0wsR11YtJJcG2Doxd2qgtKt48oeaDM93OfKx4j5Q/hDqGPDzis
zeXD21taHSZ3OlNX+2A7qAzpSkifbTRyH6ubxf+zvPukB0ov4f8pDS2NXqBRQNIv
8iWANjrojBx3out5leAeN3LusFgf3ZP/JDgq/yiBNK3QiDpCO0BUWYLVzef8kLBH
IQqzDFb+JjdHOXQDvd2UQFa8OhYO1z3DPlP7MZhO5Cw3e7BSpTO1+Q5jVP3wfzkM
bksab6jdqN4GC/txNo2B786nFfXP8dDe8ud21weYT3WRrBl67JCKN4xUvIfxRrzo
uYOhvpQ4MlKAMi2ZAclsF7NJhrrDkv/fUJnAHWYLozPpeXWAlve9ZZiTzvdIkecR
wL6mHrYFqms2yUK0+I4gxKC6NzjBVZ1eZEh5grj6Ct04pUJ0jOhBXQis+3qfrB1n
czXcJuNVnYKgbJpGI5paJK8O180Hx3E9cBegSP2oJH6BXF6T7zISjfFLalQORD8m
bbfe+FBtpgCy7d6UnVzXVMBZykZ0i/ePBa3oS43QfxxifKrfYQUv4SQfkzClkrn/
YtmMeA5pBn7aLQTn5+3ujMhxpoM8fH7DSDgIBap4LltFZ5upbZEXIRncl/FKmh5y
XN+m2qjsRIeriSAiu6kjcZRFHt4Ybc/w43FSMVzkhQbwpGYZOX2//uHrZp+kCj5C
jceLlSF/7yW8eowjtGpyf/2LCOhVa0bcm1J/H90spXbufRJfXP54kw699RfMLdSa
N60YMrB4nTCdKmJXOtdR/dzc3qhaSaClrpocsUSFpQeWV/0BBSe1/ewr43432l6p
mx5jF35efCTPxrI1k8a0kQ5ZJaiPzBCFS694mPESIcyGYPuYcsL25E/WuZ7q0mVu
CrGct5f3KDm7CxCK7E1cP7o1tCv/si28vtNlJyx35I4+xG7ekoJJx29TjOZHKewq
44VobGB5aRF/ckjp8zIvq+Kxz/udQMWT5+8hB8Bj99Z7wSJ5GiLCVquh2Pohgx0Y
mjzAWtQ6b5cwamchHIdE9Y93LRXOmw7vardx2kj5hnRaZGMeLAhsO/jWqlXRrkCI
4p+q6BflPLX8x9X+A6+DO+Bii8WQ2ZTj9kG5EaWrhSvQ44PC0XBhbTlXCLWNpebM
B3XdNdjrXSG372cgI2dcpi5Kz776etnbd/peyTxG3ZoyMOjigUdQWCxQumvjx2j9
76qv2tuG7SvUEbZQ+eDijMVvRi9I1RfaBPnfi/MD7cMPKanvDTa0Sp+Dqx/fkQbg
SXKrvX8kzzCXZeeJWpSylxG/8vA04YxFMyAzff+gLcsP4THrJSYAKBiwA3TLXsCe
6XOFN6yQftXe9EkD2S4CxPwSzqZO2JkhOh45wDOzI55k5v4pNTsc2MJC55/L5qDw
AA0pRSnBpuE4G8G7KIC5H7rzjk33Z+B0PgSrq18zPwP1ktZGOi1AyhgRq8Q9z/9S
f61SW7EzrHIlXoiniz1caqr3pel1JmF+ytpROWVo4R6rwvH0iYJ1xn7A1YlJxsqg
s5sOuWfurlDjhLBNhsxggXpfzECJ8LrFKxtof7OqFN61MMlZAhvX3M00DLydx+xF
qALRYLoqw0XXBzC7MpoGsS5pi7VUGkiTc0Z+JyEynY89PgnZoe/yXGndEcF88Iiw
cehpooZHARzzRpkcTCvdaDZ3Q9N3Pe1VswnkjHx7J4U5D/lL4PUJC7h7kvxESkkf
aLv8E/GU5i0yC/tvR1bVs3YhoQ6PoDIYa4p+zyBBhHH/aOiAz4JXZ3mBVOn40Px2
hyJxjp9ccPy01DBjhm24/SAwWWMtRVB8qBZhHAXjrHZuKilzL+9ZoWC8RTQUtJKw
vr9fha7qXmOoC8Mhmixdz2OT6L//5JyILs3Q3LzjxGfv1NvtVtnqVwUuLMNpQN94
69+iMaeJN/4HDga+FZbO9U+zcaeGdDft39hXEFlsB+va48jH9HEEl5O0xE9af1qw
oLFopQXlAUDCyTNU5XUiiEuOftHXb09cJBrc52vQTs20W2xEX0+MDWYOCgoXQy18
KLPzAvd3n6z0K2CpIL5JJC4ICmH1cnrNQmMI6YqvxZCXJkmqzi+qL3p1vdj6Cptc
gRiSSwzK/a8MguGykU48VU4zQlZyHs+Jbq0tsf/cRLcx2WqkJ6v6TlLsw2kxys63
oZVExGHqKdIdDf3ioudlAOT177Gr8jAcmlmqjxyQw14kVymAaHonQmxpF26G1+sX
U085X7q6179rShefOWqiWB3hkmJ1U7KjTlcPxNetRyxX40JxuVOKUq5xex8LsfF2
kmDdAiE4+pYfs/+azJL8f3FaSY4ds25cZXZFeiS80nMBdgfITPG4mGO3hGtBTorc
ehIO0kCvRg213A71wx9lA3jHbJvmbZOEyhtpo7dcUBM4rSHFEnfZEfj/mJ8R+v1C
GP27GGusbpuecaMp24OdrftJrmMJ6FIxXZUUUxdFPP4yl7ZmMhaNQrfva3jiCv0E
RkYOC3uwxR7M7v/e6CXuk6m3DOJOkKDkVAwSxC1GEiEyPiXMz6WSWVZaNzJIoc6X
EwnI5AE7RLM9v4ZPTFiwlkC3NAjo0p+VfnPEc37BYzDtybu+42st+vrHMeHZJ3Uw
JM9SruBO6wW+BHL+WJ0gVxpWFpEHbHWLKZ1/451yHg4kV/dYGVyaHRdJHQ3B/t6d
2XZq7SDZPxtTTWz3Lw9hZ5QPW1bVPPQzjCYfSQraDELee6r7xGqvpSZvMDMB8Z/B
JWySs6Uq9mGSmfyYP8YSyJG/CwIq7Uqiz3Nvwmq9C2YVCIIuU10edp9G+gfu2ovF
55mRurPPdBMjtMBknQuR1yPpqQ+OXPsxfA4UXd9i6TqU4mwaywiG7/4G0gk47nmH
7XL7ZISLYLgy2ac4jWIjm00cdyhaHrIAutkK7AXhPTiA2F3HvMSEUcZMwsQ4bByd
kVVG3c4lHkVpcZxe5OdyHqEmpt4e0XSQBTH26SId284QZdrFz76x7GyU331ok1FF
Lw3nXNl4EPWdbnFxJVgBVmIMKN+xPg+FKO45Ro2my8KDbq+J+R0gNg+GcduD5lm1
4Qk4y4CBo8mWDpS36JCRRPUVwHLHSEhiOlOZYOyWlO/eLzKZz66Ze8+nbXKYZDo4
xfddnhppJ9NEanbKy+PEAS60WIcOVmvmtOTYmM8zsqsUenwzyohqLv3VG8edMc04
2/Xf+T8rjMWiRP3EiU6KCHGarBEYucAbbQChMShQg1lQ6fCqSE46uMT3MnaD44LY
MAT34MmBDSrcLSo9730UsuV1wE5BtS2CcLS1CwkSUo/onqGJMr5cmdYIq4AoS9Uy
IHmo2VrRG9kdAjVZvRPt6K//we1k74m9AaoR+STjXG8/7/KfY7EGskzVt1TMlWyT
NQCITcTYkcuKNCGhxFI3oVbG3sSKkpiYpmztUj+Q56usRuRUKzmdWt9a8iSvEe+v
Ck6tYzezCWwFGSJ5rnedZH+umzQf/HjsW6jR54s1ihNaXJgzaFtJYRogQlnkuzc+
vT0qNveVovPApAomgjhJgWgbU9HOpGs1v9PelgeSYmwu/uG8bGzYrTZdqq/Lq0UB
Z5lCt67qL5Q6L7XHnesvyRnSy/5eKwOWIHHuJ6R3IRBBYhuOMju+HXpCzvNG9tge
QkSx9zYM2hPWoZ4rTWE4euFn7UvNVzL52yvy9M3x3wevyemMorweafc8ixjwcgry
fKX/quoCrxMiwOD+f/rRcSMGOOttqPMOkeMVFwIvslB/ITzuoBjrk6hwKpVdLCgC
+2//h3pB/ZR6VweYDzQgoyynWzMpdtBe2k01oUJdVFf2mksQ5jTD07509qJOlGK3
lhwxKhUD6RW56n45ybiWCWULWapiydgkIKT6TjfQHUrN76uuuzxYrC000NGLXwIb
N/jfvsqfEVhhR5h1Fp13BWVB2ZI3hCNbFlW44ZI2Fwo50pchOa7xbsGfc169wsAU
m2uRqwLTiCYs1d9x9oq+PeQ3YDGSO16Rnn7PiELow4bJmczzNRbRRNQLJZjQ3tYI
wo75yqsBStYT2pCDxc4XuzV+7rCWj2SR9GmdOzET1ewzkHpeQY7dpNUo4cG7yPac
jLI4KHmkh/YqIiyFnO2nHKr8MMevn1jxfrAHpNqDFcR5D/i8seJ0NJUQy+cxo+6W
95gwtVkg+9EWl5tgf/hU0W6BgGS0ofCg5F74xpPX1InaGLs0x9OyaWvO2G8ZgPmo
gWAlWcq/CAh19/T0CZN8zmSYFrOz2/Xa6u2RFLcSZ9WWQTvUfQv7N7kOJVy9gLuV
aDHUMIvPHQPaDH+N3If/msnn0MIzCQC3T6pvSVsbQpdxk89JR4ba0fYq0o8vAPw8
iKLIEf5UQKa/67OWp9ndr4ycNp8WrdXicVoo3laPEI+6Ad2J0aT06AzgDvJjHp24
ssC9tNft4aXeS26ZoBykSTrAI343BZioQRuTGSF6jAVQPAwuBp3k3T+3H82vxJga
LfAyT1ht69sV55pxoJXDbHCpvHp/wK2OhkKM0KWeZtb/fkLi041LifLqjPBei0b0
VjdFBq2YrKRuOu1s8aAp1vB8yYVs6Y7eFYx1fIFLZ1dkY8wYcr0Rr0oSK69aD03F
Ne6tdeUOM1/k5tHfqlOPCM2OciwC0JBWbncyAfThNGuqUWnJS4N9XPKa74VHjrjJ
tYuueTLovvPtlSqenk3pHEsBHQcNNFJ1y6yIF5lk2c3uRVTlooFyqxtUfy961y+T
ftRHgVBw9QEn1q9qdcCPbV1/IpZZX/Q6ihoa4jtODJfELu5XvJmgd8FYRZKvcFbR
GaDD0MA2FxDkCYh+PUKhKAQR0nAdvQGRX25SBlXCa9VqLkANgEP7wtHZVVdJBlmW
123VEuT5KbKdX1UP/WhVBfyEKFC93rP86XTuzih4nQ2kMAmtqnvESetQjU10Aya7
VR205aAIwN4QF6Ig5r/0cQk5MdHCckTM2bk/19znFMhqREuDi3qJGXCtwwzPGLwN
m19VsN3lnF7XNitKjeE1RkDzO7BOw+jLWePymyFwSggFqz0ZSkb0GnX/QSPhwFdL
95/G6B93D4tkgO68sSFKXK/r8lZhD+BDKVZ9GIbM2te3Bp//Nb31XS+hImwriPbM
QWd8CsObwhrL7/W74h6q8UTj2v1dNPa0U2zT+c3fIoNN5xKC0vXO36YWifcZ5Hom
d3DlBLFLjayF34BdAklwtOX+ZngAu1YmGnVDlTkVPDjrsNGykiBCRi7p4lCTCC4E
csuZ/lbrKLBH9dawGuL6F+a2/U6RviV2bDxEqCBDIGpr/qASTAMV2K8fEIfWd6GB
udJM0AM5yCRV9RwqT2DqAP/5A+qn7NkT62TJJUsoC3aVDMAXw2Aiap3ThsZkNJhM
lzrx/tPj2+1NiSc8GhYiK7kW92HkX9eAXZMXkmy//d/p/rkztni9/QnqTR77dVgg
UOalymPB5k/7uIEHSFQpHHEnuP5l4ph7kyWL725xT6GNFT9bUwKhQO+ZD/2tz+vu
PA50j3wrg82rIul08vO86ydhQpR0Lke2VkgSoxBfVfN//28PDUyCGFv58QppcAhH
1BDChF9d4wRP1cZlT1s3tSurly66k3fXXLByfNbZz0NCxqeIqZYER8aVaGSKtjJz
il/sYKUUQqfBnCMLl7Cb8+6iLb4l3GAbu+NRXklj7u/8fz2sYf29s/OIN6tqj0ig
F0RKyclD6w8IOv1Wem6/fYfkwTcgAO173ithRMlpCYeI34FhSWXgHuKqp3VcDVu2
trGts09VEl5NSi5mmroN8uPgXosr2pH/XUta0r2zwrOIOQzChRgi0q3m41wnQ8Ql
U/KzzC3BCTqlX7f+/c7Xk/ukG5lgAYVjNDMZXQAgF9hqEQCIS5Ms3LGdkqpLtMdv
VDojgPPWOG4ksdlL+UqJZ1dtIxItAa8qBB9QtfjGDu78jzKzT9BaSI12DH/J7km8
En6cQ4bY5KXkU7F8pXkE99fZN4kzbGvBcOrbWipfLPDWoR2UnXLEpFZjsPhvpIKM
tZ7gsHVWI8LuTkd7H7h3TiwMFWJ9TL/OBg8hn2HoBXbsc7Z0jd4/vyp+52YSu0xm
FJAwmKx1X2S4/e6DmTvUZnLus2l0V+SVcB+H2U/ehqGCZXoJA2DXyeIvm7tN9xcs
iqXwwqkCI/SCS6XXbJjefj6dU3t/13xjdmebSGr7NZXG+wv5n9IAV7lAPaPoAbIJ
fhUZG6u5YYdhqaFTHMZR3TESTXMzrS0/t50sBgu98vl2LHMkqq+aW/vC/iVgdMNL
BGiBx2tJeM0MImIwO8BMWo8CsKqwJt5/EXjAT/HtkWffeBOhd2GkBNJj0Q4HyKiQ
M5z62SdGUq9Z+8xW7zZsZoW785++MtGhcyVai6UBrcjpfl/Lqz/XELLn6yUTMx8x
xQPHUGpiiD7OqmKOKW3M1yCWaqpyeIq5hl3xdG/Vm+kSFFO4r3k6p8Vy2lQdtEOU
wHY4Rh7Om4Y1fyoSo+dZAilaDEm5wYkbpqvgkMqANpyqPyKeUnFXfreEOFVCE/YL
fb28LYUkRKcnbeGfTJwiBHqh5LJpBExVgDUpMoCnQf0ikWKQ7QcajeGSalkkzQEg
+Ko3R0RZVcVzxHUG2ZTznQmAqWNyUzY85oS7lJ8fGp8HA3oYFBE4BTQtQ+R4qGz+
u24etFyG3XmOU8Xngpk3mcr7Md+aeAYae1/1IAmYpgFTwJW+uipC6FVKXaMwM38p
92vcHl1EHUAsrK742Qk9NnHs+mczmJaxveax2icx0312FxRFCXuWBY7zJPYfvzC7
yL6gCho8SxL8+1V+y1y9dAHpoSCaNh0jU46C3R6pyKi6vF8BWBIwpvJOaUcpQmcs
gyuyaFXRegIVUX/9fs5rb5bqRiBIVgM0h+r/13Pr560U+Jztb+1U6pfS2uGROxcI
JGeaT78KTuhhYhZ4De+hiG1bRdb/CDBpgCl3CbPhJM40MriywM+ha+cf11GhDT5O
STN2HuHoTr8I5ZxDueMPjIJo3wzQeZv3XRenWlC1K8kldl/sdfwFMTSaZrwhKjwb
yOch+mkHzlLVoSa8IBRW5Zx699DYM4NcG8+oqyCdnao5F6Qv7fYPTN/xuaf8O6KQ
9Vnigl/CGn6itbRj9cvy24vrpx0T2z6QFA8o1GaNlLJodVhQmD4f/C5g22AOm6W1
BgkbTnYE1Jb2X4a0qNG6QJPfRFdfYZUWdg51qCSAor1z97Ug2MCwDka5lZn39Thg
aZlqvbmnI6ypKoVCLLd2SefNjlWoSYNe9Ip+16X7/bc8jzyHZ9HGoSpldieqImdK
lWHJ2IrKu1SwlVRoMXLV4QeE3ehe3CwMSeOFUhHJ3BIDAD+zJ1CcNb0PJPCagh8G
N4CB18NE9BW0s6pXG0Fe/oMt/NSIGok6cVIwWLelgK9RJJ+iy0yaCb5cYaIf9Bb9
VJfGBM/EFauDf4+zoVFdoMJR0sSlmsI2tc5/LLchWHJiEvlqgrOaMJyzdTNd4J+G
DkAgtunU4prMPuAIQ7w9KmyHOQwsFuOWG6jLBIFVUOV5FkceBDk1pK64XfwJLbt6
+zELe2LHYWiffB5mqAqt9xBjj+obr4Bn5/Y7Qf3Znbe4q9cQy7WX/Sq7PU0K0Tz8
TBp0LOdR9MKfrCS7MBY+PPJW43Xl5Xsbtk+lNoBiJOLRP56ikD6P+t0j3W8urEFf
pyWA6rhLqeajO8q9BweqfrgyIF6Sss1qCbHSlPoAVum6O2IiUcD8K1HOOs+oxJXQ
qnDUB4Sh3ndtYSok6dTYMwYsYQt/3w6L2DARAG4HZl/V8S6vzZYFPCl/ChZ3CBjV
fx+iUlJcpJsYuBkyBQRKiZ/iqZNLjHi4gjtqNpg94yk1qz+2hZf1eWIzGR8zy3d2
MHZQfI+5DB8Fmj7oCIkHK6o7LWLhsI5V6u93mt7N5xZ+e34ME4gzZYSXijDzs2NI
0IlgNs7jghhnToxsatMqHIbzL210i554zjjIZgyaCNgE2Ao8Ma8dIijVGO415/0j
rI94QmKuiayasTfoyjsYaAig8z7NduSjr5BLg6igCvjVdtp/7KlBP0uxQ9qiucNt
aLfDL5ZozMLL8muboYZdjEHT8FBqAJPUOCDwiL9XqwKklu0EKgrt1A4jn9JCSU8F
paFyxMcHCjIOoaVNtDBin20RNrL+3OKrlS9Z5kz4aeNewlFH/vVxQJlqZO5W6emd
trO9Rts+rPyLQ20YXIQhs5rpKdKk5YoM/OPB2Ka2TTth3agf1+3DDsc4r9alb/PU
1dWMTld88fqOt2bGeegQtEDYlIdml/WTQuhSz/SOLTNMzQLGaRoY0HMm9PMKtY5U
6GbVRogZjXIuQoRCZsdbf6myvl97bIRDJwF6J9epgi7FnY7bpliVAslY8SZbaUK2
jpBKqra5S/O/5wIaS3i69D/yU3jLHkC9PFjXulWc3wYMSqGkrP/KdZCSRbZxKYsn
Hgi4EimDlkCQGby7+BXL0sHqZkdKbh5tCAQE5igEAWlh12lhDLNxRUMOu3m8JGxR
+Z/d6EVAUz/+++Vz4avw95UsBqxeRN5hKd16HpRA52fCe4JW4/XlEFr59llWmM5b
v0jE52DU7hLR9oHwznVT+UR1byes8qWJoQQCUKHLcJsLOiHIcCfppR9cUUs+6BYw
/ONcvIaCGALygpKMSEmc5t0XHjm+7pDTpRdpsEIODHOBEdoX6MSFUfrjrPJT0sg8
QNxEqV5dmB+Hl2YyWg4hoAWzNzwMH7pFspzonlkHQAyy7ycYsVJ/bbkz/AewvorW
iRr0CvntJLYV82TtHMgeg1AYXNW5DWMSi9CX1+S/31cozfoKvJUDBUQiNaLN8Ilj
eJkUt/Xs51ri2cPP/W11bujfkTXoxmnxApK/+fJ9oSeOW2U9R9ge1lcmXDVNnLsb
FH9DuCrpq/+vejNsI1h2vsY4TP+T8c47QS3qSJILrobIKC3ss6r70WnjSk671fZA
DfS5n7Sc5XiOmb9YZsAtr/W2jLHrW/G2PhAaqA16xUQlVZ4+L3ROK1CSG8LWDJXJ
+6TCSmRHzy75EBeiUIbwJdCt/2Fsc8hM+RgVlLMquDtE91X8C9+vK5HPhZ0TBSPK
NIVGe70oP2//mN1HkMlefzEDv1n4Maj2qGN9I7oWd5Pprv/S5wCm4UqSYz3iLwB2
02Fw5lEJFCo8+qxLidL6gV9KFf1az1jHWMdYOG/SxiMjFH8lcEdEF2S2MQQSNRyH
fL8BW0CvlNWI+acXNdcVw0cROJg0SeHR+oNEkOVVg0aW7YeNxG19JX8qYtKY4oHY
l6YauBhNOex07keu4S6ARgUU+UozqFr0G2vhCh6CfiWcmLLAAuDgSK2rtvXCGcow
3+IqUxNZJvF8FV/ifmkN85Is1Fmkz+mnyFYj+7gbgDPLoCxT+xcIdKvn4okct9ph
HH4gCfWLeWODF/vPvt2NffdKQ8fYrxkJldunpAiLUMbkWDwDZr85wC1+nWhnGBF6
vpHiYqKoWq0JqtWM+Xau1R8/5/lnEtmyuPAiKOS5kvBjR4ui8XHDwE/ixcDHntTM
WnzkxiNuRDYgh9r22KTg8WofQeECTEbRjgDQHrq8Nk+KgA1TyQhyhPEPckkZ26qv
zgRfUxrqawuvYkMOOKu84DNUmiz4wAHVaqM5hZP/YevSYg6mJA/2bbXM0j6xL4VS
0oO3UloiX+bHuzK56Qwmz9EN14XHsimHRGnKSrr1j4Fs8wfnM7jhAAzdhUryW0Kc
yrgJWEOnh4UF0P7KW9s0VlkVjV3eCxBw3WtfgU3Onrf/XO2T+r01jnNIMPrj3zpZ
uPc96hqZCkErOaUPMHhEpRL56vNAVu6BYGDL8JKvjRSi3SSu6PDvO7L4S7IpvtHW
kV8/pk3PyN/vVnTB51DxY6d3uwES/sQtYfe+a6M1j9tKN6YPXJZEnv9b0BPErnMr
6qeQ2FOUlmo0gQJQjUfQFqNCN179s8Qfljm/fpihQaX+pqno0qKd0Mn7eU5IXHHF
XS+SmTabjgG5DmPPjPmU8lhvggLDcVefJ3l9daojmqXy7flfWHAdkQyUeiZ/SLRG
fnonKRDfIsjDI4K7EkKcyzhTN2iqd7b2CK8KG4uZ6VF8cHsxdvRpPBAuGsVdK2Db
PtCJZSVoTkUG2t4AJuY305/z2Emdpjpfg/kneubjj0B5cAaJVz5OMo2bNwgGKtgK
RZGMqnQ28aumE/liKfZfBpWUqsD1K2Ayd3+FGqzZyrxxflIzt/fLtn3btBZnw+Gr
3oebdGVyT1hiwj6wnwy0lo5Rtfpkj82lpvdlGz81j6+Xc1VyLra5jy3sg+VCfq1e
wBZ0xlaoG9VpNidItoUXPEusSV2cFOUK1bxsQuFWruQHmAS41xVwcDUEhgKpOWqe
jmw9uUC9V4gbmSW8UXxZ1Z5fWfdTKnjuHEn8Y4irlk/eH/dkujaleZfRgm6RDZTE
xyWtGQfGeHdxpIbNSkTIIo/FQk3c5CSieWQP18k1HvUvxBCiL7kKAHIl0hScHF8Q
LqCXRzdm/8uYwPBlkil5vsB0vStpekR3+L13c9wTfsq6QfG4GoBlorjnu29L4I5H
G/Gyvd3vg6T3MWu4LaQrvAHMgKt3b2wfYFyAjD+npZUbeLfAKeFwvD2b77cYaNxJ
sQq+/9tEZkBZMGJuXmBl9BTodze7dMrlrLZNafWr8gDjnRUBq32IBvn2eKBVoOYL
9GDnHiG/8l/Kd9M/cwomtR5rTc/md/dEu+Qc5+hyc6jFbt9NHFBTlC92aDVZNqDt
aHYCPmqnllpmAYNp8B6YZSGSbEZt9Dk7UgVtnDrcGJyvC7RY8r9ljaxBCef1Juaz
VNIECRb8PFeGRG532Xn59u/sXkuOPIpm5Pbpj5vJkiqbmBjpBrOgUYEGcyelhTBa
5/QiOi5TO3PcZ4zTEKsNF6aPxbNEetEBqzn0dybwlFgbj349PyZfrmF28O2l04Pk
YFnmY88WSQY0ZBxlGlJk2iQgSKUzo6TXa4inQpTDUvlcZUoS3lhbJo/9q7HeE3IQ
YPEf4pijThp2hwmsdd3X3hAHqDTbXN0+XQ/5ep618pKNwkL6HRC729NnvL4z3n0v
emnYiPHwOHlMwAPPfL7aMrAqv2p4PZrK9UXzmNvNC5PbKB0wWX82SLNiq24xtzp/
QCHoQxOG/fHAwqYYxmQ7crDJAhp8VMOzuC0jcmENcyM2eN8cQWiGIA4ruDKzqCni
ZtAWNAPCVuBtFqu+Ucfu4cTV3GlmOzpCUjDfalfKB08wmS+gb05atszdJfx+OFMZ
d5TW5hrDiF109rOT+Stkno63nFaoySR5nvhSyQTPAaPgMmfl3k0YhP9RUn3qv6Pd
aOY9XDczs0Ogirc79JlE1xq4Gj50Y4PAVVqS76uFG5y9Y+VfCh8/V3suMuvhQQHb
gl0IaH4Gngwq2oVBHZf81j+Cobkg22BFWfbnd7DjnZNUIvjymVjgQilLOxHh1oEA
FjmAOpyEgMmuHTuigwyYtWhZBWRKpy0z6XO/vz0vABOD8Bn5AurIXnMNT/aPgYHE
0NDousmiSATxjXmAoTtgWKk0Cweg1LyeGm36NNYVjCrzIHgybQnazaZ2+3aCNk3J
QL37J5rEhWO+ZI44ZXl8tTwV1GTUA8mMYPLFlTL4jjUZ41QKzst+oR1NJtJCBrw9
3oxsFx1b1OwdUhGQ6iiuq+K52UhfPVBH1ihNogxpxGjoxKxjh5fZ+XyE2RaKTjFV
VOBhxWtrF7NGh3pHn2Zka3EdNW2bV51Vif/9FY6ZSCXc4o9DpUWOVv0smP0rQ7+T
yUwznSYBahYzfK8RuXt1MPBsU8zJUNL/pK26V9bRDcPXD1zy6cyIcPNVRyu1RNZ9
U3NYdk6PeiJMXo81qR5wUKZbg7jtZjgsi1FEgiSw9qeftd1vXvaWp3Z8Zuwd+xz0
/Hmx7g0JUlD5m1LevE/Y/pEx8RiikaBuP/9FomgukX7iV521z7WasvLUIQnCqVeZ
j/+uWHiIUNzmKrsSkn17NUgpHk4u6pvVisj3y7c1TWQNJ3ucCmco5eehCwwfFkdA
mFr8uV3JXHFHIx0zC8Xw2Ydb1LYrFLOon9wM08QqJWjl28HC3bDfN768OwEPxQQR
ukdXmD1KOqLv7tIrDDUhk3SSEzElfL/egNtCkrR4rFos+60meYCIwBvTFQRBWV0f
2BU9pipuEKfPa2+uIG6CThRn3M70dQ9g3yZeQVFa74LJkBOT75P0Gg/YM4d8P10R
niudQ2xP+BCV3IajY7DmKU/VvJFI5ASWLxstNJ6CDVTD0s4opp33LtMg92twLMce
ExnLwtI2AVq0iEOEHtfPgUrszMsrcso4Cwz1QkRseRJarH6lpFLIcXoUojQH8CZv
p/mNRA/+NrsDyEWf46IPcgXjJ8m0RZT7zx3a+sPMqLRNv5OC2/SNBRM6yNTq+Wq9
3VYjWhy/O06A5PTp+AAEnN22Pu4u2BtNjq7p6mF08v0fIQjC+EwRyrg4+Pk6ZXA4
fD2/hoVRmqlvkjOUwVIDZdzFgVDlA+c+vtw49ZdjW5hXFyxXuSy8fPm5PmENRPhx
qnLQImgavrQYfMOtWjj51KpQe58wO0WC01/SfOdzW39yrLfe9R/qZaChmUBi7oak
8CKm3i9//zFL8efPS4tBNGBatuNacR8RU9d/kfLG2Lci416IqBQtCOkBFX8zFZrR
lXp6OKh+GiTc54zZDRMwiC8kCq3/ZSvmUqSaWTCUU4KTVpSqLmLiRT24PaGC/9pu
JnJqROCwLki2ZeUaYAUqu/e+QQUhDCA2dKkUwFpJO5VUdRKX4noV0gSRk9KL7iGZ
/rq1A1wCteCNJ3amRAUAqAFMBgVq4LGGJREoANTGOjzHhK38GnCTWrRUStS9rVDh
ecJVrkW6a+mHpnzyxrMVzW2vE0HGbGGeOC6C1feZYxiwODONwfbk7P6UrdfDlUYg
/nUfG6klzpC9h6q9O3Gi8oMQpNg/0Dx4DyPr6nbxGCvMXoBBWr5NKmzDBAW5JUfF
xMisFYKT+VvFSmLw9JLI+cZnmW8gA17YZiJsIhUnym+wRlN5unM/3eo7wQo2XhlA
Dy59WzF3n5avCJPlgZBPPklzJ8j0iSqMc2VK2CCIWgITvyEmsasXSW5ajZwOvST2
5eZHW2SV8B4zjPyLdRwBn3K3K3todNa3qOGOVARPsPJ3ioeJsOBvo/0Vt+TmZfsK
ZBwSpbaBFBHes1JJ4ea7weRo/39B5TRLpd3wwzGSSlmC5gVthcJ45ePeIkrlHOGz
Ffbo1S/c8w/xkNTg3vi/s2d5GJ77Z0KOHK7JWWPjD68Fv8ADhPBP0sC080lONMvm
zMwzJQsLLdDAUNiUURpFCxtPoMXnOG3fozgfBDc8xGfrO+taTcY3SkZi0Dxa5VU2
MO3SjbmE1bnND2RMlyO+ob9dcYbFHeosrVTQI8jpxJHL/tneFcTjVYz2uSGhnRzx
01HNWwJYBSNXUmi09/RFzDtN9iMrevDuFgXQa9WfpPXqGeB8UmMokkoEFhCatRk2
vBSoLBgiDLUqI1LO8WTZYb1u73H8yc3A8VI/Ke3808BC1+uRCtloLbH1nZ1Bn7KA
W6l5J+eaUmEirXnJwVtKkxICmiwDy6fw636DvjTLt8Bmr/YLSD6IXLDCZqoK64KZ
H6bemL36khIp5jDl6rLrM5+1ot4XCUgw+Y1jXHGDasXdoRHn6CZyLVyvW4PjP89f
thKPGCcXEXQzp27SOOXwVVV0G12MiEBcJBPh+dOgNvuEcn82HbTRa+h++3exABzP
k5HsVhQVNJAjBYMCF3I9CC3MZum4J+yM4J9hhN2rYU+HyKkGGdAIl4BaUQVlOCMu
ECiQL2u98HI+70F8q0G1HmxpwWJPpinSUQD4zaAhOlJazCNDBYTAEWehMxjlRfyl
3ss4UPjmRr/bNG4hy+8DIjRQpGiSwo5onxkz/oT0oeHQLliCvJi6QByJKztD6H3l
USE2VDjpW+OuG+5B7Nq6JNlQP85NLpuIXD+rSfci+DiwQoiadtYT9hog62wHaWCC
+c3wsvWNz0YuF2JJL/DGa90MX+WCCpcEAzN3MRHrhcWptH0mb7IZOQZwfSOnkGIV
V7nojS38gO6NLKyjcTErg+ky/aXNJf0BjQBJfJETQASLkbZ/0vengEhgDfXxQnpN
yXv2zCJDQRbUaV9SHiae8xWjbIxA6z+D1vWfDmknwhYQC/0ag3Y5SsrqyZssz6pq
Xgul77xuguM4H/bP0oLiXI0zZmCav2Y1ghloqPeeElPq8F+4SLLTUCX9N4Q/VQF6
yiZ586i6hiI5J4g54lV3fP1MQhQ7uFHUPo2z/HRfxUaaFDLwIZieCDXpWonmrhsd
K1i6iIQaMJQFfi8c9xWpKOU6QVY/tcxcgK00qajJnJW2626JargbP3JnEZuTflDg
i7aQImavkqstcYWfTL6lviFI81yQbNhyy73XKtA4N68jIj24lPv17PsnNuNmWLME
xZaTtyXma24iKlZpsFc5UCeYN/dfsM8XL5+ewrgEIGlM8rm0kjQTHchV4gDGbCae
dn2B2vIacb33UsApiKPQITMKJwbg0jfNzx5ZaTm8fM387RFGuHqvZ0bJ8z4I/567
pqxZXYXrY09aRi1tkmN71NcVRS/juNLTB49XfBUYYUiOvuDXRMziqGdyDRVW0zUq
lV32TRULgJaIK6ILkF0Ksjd3fDh9IMprr1gJ48cQq8taRLbEiqEKhNVCYOVbYFhV
qdtIG6LLjIo+OKJN836nP+zQbNhj6cODgtfaqepdrk/Ff244Q2PbMYP2Fm/7YB/9
Rug6WtqzN+E0ynRYHiqfWJrJyVdcGGAq6vb+CjQvrSiHUqXgky8M0jtJ9e8uppVu
Yi1j1ay0wiXUQZruBYnQjikDssxLFWW51v7tXoi8/I3pk6hCrloJHI2bOb4JhPS+
LLDxKxN0hlsaJBG4zXuUBpXPljJg0/Mnyo+HfIWVdV6jpMN3qjiXGT+1xFfvvKpA
7QXzFV/lY1XmaIJne7sNxS7rtzu6pUtqQEdcGI7HzmQ2j9GQUTIwLEq0ct8rqT5M
jETFW8LX+VaaWcP9noLaQSkczeCYVAw0ZnP7bOY6BFq0aF20E3ftDS6O9vhKTQkV
rXTB993k9UnZJ0xLISiJNEA1PxMI571Szpa3fsg87Kj3Qot7GfxoH97nlZccj9Ke
fSSJjBTed+geyAb95EWT2oGQK8BTMR0OXJi2Nb0nI3L6V78HAxcS3d229ZWvMfEm
+aCDArGnPaMcsJGhoH8Umxcs6nHz+h5axvrxdU6awaE3MOjZtYqwbjB23YL46LUl
QdmmntIfiFhvLo7lnWCdBLhPU3tiZ8iTABeomnS7AzSh/ipR9whvDKzxikfEwVvp
LUyldiHjzkp9FN+Yt8esBionjTtUj+Kng/wwLUVHnumshNtMQcDhLdEZ/gL1A236
KDE+jOM0dmHainQ4qt+kP2qJLCDTLv1pP/w/oU1Y4ww9B5HO+dRmeI6xsOgdeP7n
FLz7AXTCUX/I7+gtxDcod7lkYQKNFX2DUTokFXkNcChU+TbQT31nY/8P7TQ8BlvT
dQZLUlu/EBEEGcssvhGinDptyznfaarAXiYYbotbtvZ2LmWwS64t98Y64XBcwOA6
nBZn04uTbO524VuQ8xjON9l7P1vALU3H3vDCFWdxt7vMWnG0nKVApoif4/nhnMe8
6FCoWDwrAbHUqUSbtVNwgtR/JAoD0JrCFymIrncIRK5E9ePe9yDodhmIA7UaW6f/
M6gzbxOoWtg79JN7oUzn9i3NTrcXEMCkymDILd5xUe/g+mEkQQPMQHgUZLQ20Clg
5OrViOyDww1NmAhvH1wHKsraBi69CuOq931x7ixm5GMflcB/b0S5xquFIxEZlGG/
QzIBVtfbhE8MuTFB9zhffy3s28sWyeUvc4wjtgiNtWwU9dkh+dnRjVDYOPZRvEMO
ZeRdwfG23eXJ+N+iDPyEniaSV2+nBb+ndsGHgpA9TGmpdu7ThICi23wQwwwVQTt7
c5krTqRMpnSMhXGQj1vrRtpRVPN5tFGUxemAsCU7f0UwMuQpXocas/6CmZ2Y/X2F
SyDSRWTDRNNFK68MTAoWArPeas5V5Wmz3/SuwDrhFy2bpD48ySduf3vqYLKFdlLY
MSDXpm8jC9zSM36wG9+UUu8jEFoBFsHAbnNobmcG6MmFiNkyISC7paN9Gy2mpl0x
nEKVOUOsRigj29XqmMlxG1Ag2jOjPq0QW/PBwpzI17b3xIMzbilaKZ1DcG4IxoLa
jDd+lZsFW7au0u+HiHtj43yyooiWpEjzW2pjxtJghYDbS0fAaIThyg9aiYtdx1uT
xriEe6rEWgg8mSt9G39o2/hy9JA7jgGQjFqcXiLNZHPhXqNUJj/dQpDNY7q0FoUv
Q76BuLZydxp9zRocbDOJCpqoXGjKSRKnNXAnMdzkUC8hb8hJH+9pdrf+QDssKzXv
0QwgqQZ3UbWCQ6jFXWha2SCLp5FfEeqaS7eYZha/gs3H8CHfBWeXH22kDmQHLy+4
+PPVPRw03+GzIjyyyZBEtkiGWPRtGQac+HZQzrRR4Zm0vLpUd4lYiOpsEzDYETNU
qmwzzIkd+NkefBzrqbcTVz3A5C2TqE830H/Njj9siwtoYuuYmmVOh79reYSvOpi8
mWGzHuptQpchlJmdPosT074Tc4TdviQDnQFJQMrM1VwYWAZKc7e5JnKgNKd6y8dy
jx3CZvouSwCJ+oLlsbW5jOMTq1RtFKPqrKxda0rS1qzEDKe6zWehysoNE4+nuwDx
ZWDB4qMcFg08lj/5XaZPRKHSbZwcq081emFZ++1d+ssG+axiivPQRBokPinPm69m
Pe0pnSRixT9OG/FQKC78E3YLhrC8ZwujCsPQt5EiEwdEuDYHfT+LIwZVEmvvorUR
2wUD55wUBqu4NgQmd8HGrk1iMy/4QKNmn+6pDZGMMHX7M25wFKTNN6cx7z5Lb+QV
JhmbMwHdyDKKOEirrgONIPwhtV2zIxDQLdYaBNY1ELoomY6UCeYKYRxXi9Swx72V
1qb3hCoDSNs0gzKQCOSw06Um7tLgKvGTKKmZ9pPNjtGmxeojRHxfxzpPfmVSEgr+
2VWrFDn4uOenIWXIEQdL0LHrPW+I4y14rg3KmNcjJNlw3HFItbxj/qjY7SIQH7CX
8nVfHcWb17WtXzCBjwGTLYgx4VaZA8WRaruX2T4lAbbfwpmHRQ/k1ztfyOfO2tBm
lkc+eyfNGXuYGQTRS3QiQ+SxiUntWC1bu6InFhOhNgVdLQt0/5cNu+UOiXMf0ye7
RvAP0N/AAfgDvXCwaO/7Ln83ur/GgT/5i8eZGCqNcsKmdgK3snPCafW1Pw7ATTJ7
N1z8C15iiCUJ94eqBr1HETIcMbEJ1/OBh4wicEkTxnqKpneTr7NAZSy4P23m6YtP
HH4rRkAdyshhaiBre4lBMhpHLdn/4w78cDlK9RG6rv4xHr2891LY8mWPd3zgYDkx
0xgJEnzbFU/ckumyDiFNl0th9g5FpefEKUn+aq9p0zXXy+O/SxGOyby0qFYXQm+F
L5A6xjsv8cP1yYtZufN6SOFweIJtrQIui6UXRy811NQs61ilVD7/IvAlZW6As2jj
Qrhc1gV1GuL55GYzpUfleQ0jNn8NaRG2Se/9j69dBdpHRoQ0Eo9/H7bugdZ2ukSA
Q9p/Okf0rzk7EBFv6280S+jV/9YnhF8zp4G9jujbz+rx31xKEJQnsiVHPse4/ZTr
5kp7TEJNX2MHJi6qUS1rOB6wkh1rPqCUJVhsM6mqC+Jh3ChT1K36QR5RFETIpdzd
F4tSSJoooO4xzf46VsYjZtzYlMRdF+kEz0pspyGq+y8wSsrJuWsOd7aHWEzBAxE+
x0TyfA19yqT5SrAJdJUty5sD9OWNwVGUiA48MIJEnmGuKLiJoviqeJwr7cKN4EB4
87zQZrkzs1bl7s7yt7PsTyt0VVjX12wjdpZFcIvDz1K6vbvlfa4TGP7A2+pLDWJO
+Slzuz+f57R5nRglmtFIlUu370BjLPj5aon7CUtP9e0dvYmhYFLcfRnFuRZzlXpA
Z+3QWca+Znh6P9tAsJZY9vwyh5hb7rwYOvKo7U4yZsUD4NZZ7A/FCBvRqtpGlqMq
dbHYXk+2ABJvcCg+/zKpgpi3Hz5cNhjI9neaRoQw/AYq76PKHL2V6lH8caHyvr+x
PfZPrkcjDhOAs7kKC+lZWXNxrTzNj0RNVBWWkPdR72Q0SMjBIylmzdSrEDcLZ1n8
o+Da/xqzZdxhPvOTbMWNsyrRVpsJjxa8WSPb8avq2l9VtsveVtSpPLcftqTYDoFx
u9yOlozzPogPKJRkhjRbEsqpLw2pKeh4keUTT5oEQZ4AnzRgvoTY6W7CbIiWfaXQ
4xvPPDrMp9XvEeC66/9po9mEqOKzI6wg6Wwe9LFegK7TRL/p5y7OJrOPOLi5jrEv
WRpQ2nNRGmJsyFmmitNutxcS4l9B1J2IChcztVKn1ClYvad69543S0z3hI515Q4s
766a2WyUhVlf1JKndhurzCWsvNQQL38FtI/8FOl4OHqeOW6lCflcSwjF+41CmCMM
03NZT/4QwmL29+Y3NMtOioyIG9SHHHEppYv0frYHWSBHRW2bAcUQApfXB+3iwiJG
PHniUUa2KolpA1XdEL2rHabraVHbGoeKW+GxE4s6f8QmRydcbKQtDcjw165YQBl5
GjLQo63b9jeTxGgA0M2bEz6pTaZ2AI7lY4mGs/ynod51mxiAqMYwECGv4E3l/wWd
OVG6YqGYP0jI58W1rnVb7hbjL2mJH2kteBly29hBm/yC+hEvlMfLTLpfBZ2miJhW
sHmSWzhmiAcgQ1BKN+MNyWNZnS4Qr79x6IIFaxKIH0WxZlcjkMvjPbHsqr4lxdr1
Rr5d3PUB3CGZdXJMLtF32eap/v8oFYYqBc6UeTZfxHeqoAawij4a6S0K6b0jYN/k
rg+RXZ7GdU+pi/AgEpOx/etI/7fjGYaNjnliA++4v3jtgvHGi4osf/ctTQQZBYB3
byx+c65Wlcohh7+dXti7A0v0FpHfYoJL3aIeLTJ33aXpb46GLor9cjGhnSkowib2
0u7hUcEn6pnmz+UX+prUiPPqtYDJOl/gwpE0coDrvTp9v3zW2260TP8JZsByyuCK
wi6XSzg8vBqEmKlMjEw3OO+HtwKOA6WBbMhaf6LCFciduFrx2Is2rd6wOv2usfJJ
0NLjko/1QMJoCm/RslORF+wP3gDHKuT2oHhaEoG61g4FNlAU3p36Rl20UZeQ8iUU
rffqfJIFChd9hv5q/PNPDWGGflSHsJILyVULSFMqv8f1vWFtq1Eiu1AoPdc1ukwd
Q1/2Ro/rmKH0sg8kJr05dRtU0rl2uOnz3KImqbUPsTM8Ib5oWZeupuN+fu4Fc6Sf
njENn6WmGpkOGsW1c/LP4JciMO3GsRnf0HoyZreb7Y8VneuBlsUrSrbGR/iG2CNW
j5Ya/JjkTXKbjUo50NYKbyxfJ7rJw0YROwkS3wDUdZDILqREzxtLZ+6V7Zzlv3pk
V4DLUzy61Ra8OQqWxidFGwQI8S7YT/hrYESNO5H2zmLnfmoUCcaFXG2Gw4Me9zyB
JiUqxS/ec3R3DP+gNG58FxcYK2HpJwuDRhhW8sYVr/UdCgV2mvbIUyWoYFGL6K9C
PLZpfYT1UQm4+4e+aj6DpoUO8hubVZb/hKk5vhBUOHpKl4db6ilYTJ+07kOeALHz
V0CC7CgskIM31MBH3SiTGzKq3Y3FLthcKxtdeh0HQn6hOo39h3xrrB8ll33mbDyt
u6tYYJTMLaZpB9ZP3toBcw==
`pragma protect end_protected
