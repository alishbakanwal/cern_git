// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 13:57:47 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
nHmXp2GJgxd41yjgFNK+3JYmkGiASEQUrdleT4CRpIzayNJg4TGBqMl1J6YOY3yh
LT49KbpElUV5S6u7VMMBBWe60Re3tvrQsEKZVoTIIcU51gHPLnDSKC+GmwmjGHVf
krPbYhnAZzY/H3d5Cicqu5qIX5U16oOfpsyfdeS+gmk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 104704)
PT2PpMd3Mr6HRdJs5YpFFjdO/jJGivv24UdSRORk7Vc36m89brJ88aVaeH5GXg6H
0YeF+QrvNCU4LEqjHO6KoaOj7AL4Ej6rhYZizUp7xtSF+PBwYLlKI7xpu3ro24x+
ZmxT/TTF++FtL5kKFt2tAi0Gsekg3DH6hjkLVR6fCM03Fnr8KBOBSdzgg5rWxDM8
kErAzBTTyxRprTgWYBkLMoCBwbf0Gm7ZEnVEP7mRbhWMmLLm+K3toJ29X/ecvvFd
ZZrbXmXgUaouTpW8xYBHxKKzXgWoKcvUBqRx2ekk5EBo+0JZub6XYYbyOg2q6X1Y
bHBNKzSmx5IvlwsW/lpuyE05+2DJLMnZaojaabKifON7iDfN0I9qBeBZnbeRE4Eq
ERCev3RWOwxdPRAxQI1y/XdOO55K7/MPlzIS5ZGW5Q3k9N39DHlezfYEMhjL1kIT
IBta+D4PH4PVSM5W8bFaomCuoCFuccCttRHYWV8cYcD6vTwGj+IkgDthNlMIgtLO
ad0D6BV7lBwtQrJxQlvpuC68b/9zLG+8kDhgjwFJU5EGDx9HJqn9xs5ZbdWg364D
Ag8pI446eF3EJPkr/1bB1ucHltmnOMzPtFxxahaSl3ffdQgaejAcfBxj5GuAR/hm
sRnTPmJhtcfiVwL0HJSDRfO9vnyXj2+66KmESSOsWf7SIuHttrhFjei0bZfcZPeG
c1QLQNgP7D9lpBxZ1sFER40Q31b4NqfiapICzFDqnBAZVEcdZwRD3OnhCiN2zS8R
Ny9+9XCgmVmkdXEjXIBg7Oxb6wo1r1+utRJUWAzJimQ7w0vO4NkPhQSpI/T40Bpa
o+js/bYxd2YgN48yAKHNs+9mJ0Y0dUFUEIlWo98/llI/nKifwAnL1Z63LRHhYhLV
zWE6TvrI4jnQvWq88GrpS9FL2yhl3XOCvlKyXCroQCYLgASJfb2pzWvx7WQG3H9i
Fin1aihvoBP5AbmgTHG9bV7XeaTRdOWat1WsknrWhkt8i1wZxvEqSSr0OjHQUHnf
1i98xvRg4zuWwytCNqGi/GZFH5eeaFQFQHCHDibQJoVSwrdYj1hea5cqdpoDw/Lz
oqO7Pz+UB9CPAR1WiM80sbIvWooyglXgEJx7OxgK5evNNO8W4yTquidU8TZWgUb6
WJ76lqIIYgsVz9QO+bTzpIEA2N7hgs9KqdKCUXOccH84fIFLKTBXV9zA6P7Zl6GG
ApdWsNW/YMM2wtPmqNd/6o1fqhv+TrRBkmsojM9TsupClNVFJTejTzyZ/LjAO9XG
wd6u83hoTEbTA1Ldrhfp+RTA6f1dwmFz29McwxOsT9HNatQ+Vku4d/Ss1JIBQP3m
LBer0HezUyAO9fZzI+I9T/fBXPJpd5WtpXa+sMlY2V04e8X2RPPYMr0bjDEevtbP
JT7an/NAMlQKVqE/IQoURTe5wqJgFrqS24xdhBhw9c/Ej4fYRlyg4AuOq0icKQxl
2NxEMNTw9XcEKYtuduJ3wwzuzOYK6ih8eJcsPKRN1n4sfB3lIvzLq5orkTp5sfwX
gkoDU8letqK+AAaBdHaRUCpaNE49SHCyiB2mqJYLsw+VmhT8DHMf/GuOH14+Yx/l
QFse7IcEG0sEsvO7xBbCyiuKruYc/acVKDnAgHjmRQCCELUV8aM6rXh1SEt0OS5D
Hqg4PiYms2WUiFupgjD+o13sk0/jA1cozbaxKy8P5OFY//uUxXm1O+sMmepyU3+i
7NrdVST9htFdHZymaPD56BLhAhK78d5cU8ABri7Rer2Z8I0xsHFv/aG+xXT1ngsX
0OgB9F3Hc0Qn4NGorAKg0N8YMAP5OtiMj9oSCGOSvnyseAMa0jXd8A+rQFA1nEVf
Q+YzuNYroxWSCbQywODidRVOA46TpFZPUmgTKGJYU3goEh+1xTkDzXYhzcIsmUDT
FsouNeWi0zqfhWwtmPYGu7r/i1t7O0YFf5R2xZA7BVVMZeGYL5FQU/hHqqlWbpmt
tO4UKOXBGxKmdW/8hVcn644Ql9cNAEM33tWdr75zfewxrzCWAu/hnfjeDcDcBENx
epZ9V1NM7DuVSVxQ3igp+lxsfODFPDoYrVwluGTIzz+u/T7SPxsMIhR7ERS+GMor
8RxcHwo8v+B+Tsewonu9/i0J3FMkxGzl+LP+AHgiDZqsL3w+yyxg64hvMTtUylhb
G2oYc8SHkHV4fg+ZPfR5h2O77gP5lcxHfmNUZaYq5FPeXecMlBQPDMTqtySdPmLA
irkn/XMOPa5bDnxVc5PMzjnO4ekSYemY4SVTCxll9C1sHz5i1My96LXxX1VkLEP+
KZSSMplTJJ41COPZbbWNXcrTUcAZ/o9TjFuzXQvdpfSEloGCLyexj5T4U4IgpAD5
OepgPYnD9DM/P9za1JEylSdHYrObbK+75aPhX9NN2Q0Qfk9iAD//jXb8haWgiPBH
pqC80cRagcl+6fj845q5nPn+zNF5oVw356PFNRJtDuEn3QD3txww/3CGSpMYgFSD
XemIdJpHEizo+4FyBblQXqRJJMxtC5S+F1mWj75ecuNmZm13xvfAttnfUcjFX3Gz
6ahJ81LnXZtrtppv598rTZ+nnHohLP43UXaLVwHSexNKf4FvV4l18Ujn7602T+AK
DR/BPkIDL9y5SSX4hD/1Y1pGtJFsTIiCFzGHqL5wVR4vOo55ELjOBG2LNApOLAwu
+zUrHdHej19WdqbAFJSQie3NeRdwNALTGWanuWlXln5Kx+GszpZZtD7LueLuMQ8a
87H9ei42OFmIPEVrf5lRPzVUfXM10MJAf5J5aAhvSYQgH0xYq7x2gy6kf55Xc5T/
FCuwXBL71h7slR1lzRGzMkMmcwsaCmDYvpiqmiJnOJmvjzeyUcV2SHOnsyI1X/rs
LqJntYxB4L0cUlNBDre8sszY5rZzHL+uSbRfVioK+eQj+ZD93QaLsKhrsjy6/FP7
3r2zPBI6uzZtWyoe0xRblVN1dQP0Mtmi7F8eDoY0fwSZw4eVHpsl818NW+BDE4Z/
VR6flZrJhc+vVe4zi1VHLYBCrt8mqWPmr3nF2QYE4ErAdeBp0KEq9SmGlTsIOplC
UoAd0w6oe5BERf9tU4Pr9yeCe+gu+SzdHjVjiLf2cnLyYHE0WE1ggSQ1Ob5/SZdT
8hNxY51TlGnlqZlvzxdbfvg2EBBv6L/6aJUuI/WyLWUfwJmN4aJHneJLFaCiopvC
0dLWXt6s96pSInqdoFeXn88kAzbJ/v3JuYx6u82DmDKXOKhP6V39//F43HksxpRP
tVhrIFnZdMMnWJJHOxSpF/htlUC2bVXz7rwuV3bOtzSffR/p2hAKuzAJgqf9i+IX
e7NQcOeGfg42rsGZtkq8itcwAkGZEN70V8Buc554AWRlw6pgn53MfWViP+jZg/a6
RVRlru3Szp5iqb3aAvRuJKMG3bc8qxw+GvUkGIblFpF0jlYrCHUwOOHBuVh4mUEj
cha061ToTgFbcripIxDUTXbekz0TLb9vCejnvq8fHZNN+vUAmNjWWveUUcbFovq1
KMPuagtgztxSL5VSb1e8e/akQuqzrg2mKOVOuorNABd3KVtnQjLgcIbxP8Gey8i/
QfgxisVUYL9PFlZ3fflivwQi4l4xjZ6Qz1kN/8MNm7TSzrKtdye9QAnq4xwY+ZWJ
5MRlwt0VcpXp6mWqQm3PJLNwJJYqkNa+TfKBVc58q/6pATwP/l3Y/qQRG7Bw2pEI
nMTLRP/7pJfhh0W32Co/osO2qbxQPWw+/WeP7Eq7kqhrkTRfqoWL6Uo1CU9C2kOm
NC2LDVWuE3sRjwRLQMiPwqYqeVfthxzlc+dDHVFX+BqbKC6hnDIHmap56jrb2ElN
BJdJ8ZdRQrwbzzXSsAp2elBvCgpsro5gPFlXe2awzoujwv8DoK6GpRBMZabVps3K
AvYZhWF5ktboEkB+m2R59RBfI+1gkXgW1yLSYnsJeRVAHkJb8MO0FqBqsy/F6C84
ISu4qOCTYjd8eqjVLDNI6ff4N6M3a8iCQTzuObuIm4nP6qLi/jLsaKieDNJH2Cr4
bljJCe9vrLdotdRODts380TZBvI+mGHEPP+6dkHbTPUId0k0GB0oJJsYm9IODjT1
qPVh+mn1fdJqY+pn5cssm1IT15NS8PTLVGkaKhQF0Cp5/R9NuRCMT91N1i36I3vt
swzxb4nurT/FNOzS8+SxIpua66aqT4JEv3x38hRD8MUMrBN9dD6gi83fizw52JwZ
zx5zD1IhKYYQUNvdnPdE79I3Rfrvi6kX9XhBG+pcYuE2Kk1wtacztoMvEMmPNu1t
OIKh0CMa/IHEOyYARsZNwuioA6IhhlEBfubWvcpc8OOh4aVGzP/MSc1PfkrCGttn
LLiKXlLgjo3SsokJyaJ5AdZMS4hMcOQVRqwclydki/dQZPaTyA01WjWHtQi7A9vt
AsAsJ3cbZnUcEd+m6+3vvbna9xUqSIO8HwcAL6xIc58GeZ1cWzH1vo1lXSez4fE7
mVSfGCWAl6kFZvgis6LPttCe+cD49RIjZ1auF/c2uz9Y3beU4YTteivS9dLybNOH
s4uA4lAlvYQDOgLluu5gRcfZ2ldlI1/54V7v5tFSohOczIDhMk8jBNz77YR7ohDY
XVDJG4gUCKliBJXg4E92qQEGhGw3rTvdzBbegJx14yoPlj2kqp+K39OdBzMHo+jz
he2grNyhcEyS9kyuP7lVoDzf2YcgpyaVE3imoRlAlyeF1xDqd7MtnevKRi5I6wt7
fVg1L4HEz+IoRJdnMWlFotuWH5L9UJCCGILDD2QbDwT32W2iWoSbmZvj0OoB8LA8
D/NA3wNlqC9O5yBG+X7ikn/YGbVwDBbrdBuq97EHr692ngWi/GIydKuM+Fxkpg9F
pc4a/KJEZjIoxJWSRuxPMetwJIzO7owPdtmIM7LrBGyYDhfCXFUVGxjWhypa1iFc
sZio5x7eVUQ0NKRqGqsKeKrw+3E0xOFVQfo9gNPnwgIgI/WkLq+FJltPmhFyTBRI
DfNOkWKZwahgo/eOigSjAjXm8BLbApzNYINJyS42MIuVneTWEVf/ikuNytLlr14x
GDmReXG3TkPPSyjCLIGHhi0GmjtllVNhxgbcqFUyR2jjHOuqMnCUBXp+0yw2zbBb
L5kYQjRvQXTcvL7/HygFKBobfN3O53sDAoMb6DPSnll605pEuITvBuEVvwAhqab1
fJg3uCdP+Yg0O+EQyKY2keg7R8Gi8cHT6jaMu2qkr/wqwZosUuZx4Ni5x8Pi7+Kt
pjwXI5MJojXp0XeGLGK3/pIZ7blnMD9hJaIF7EJGf7Vaulgwke4jG5dcvdR9dMbl
86+djSB+xFPACvf80TVY0Qu2vOx6UrSN4+8UZxzdXwPMIqvYOLPhKo5BteJ+5o6e
UkamxPGMBTFc4LMJt4aQq+3mGwT+LLEf6T8+w9Xc+kSmmBD8GXIhl/CljAOrJ3E4
0+nTKS0zhyTx1FkiLBpiyZPgZlOwJ3CsSPBanDGsyaZXd8BFwA53MdREcZRxMKwk
XJplRO8erZ5OoQ4ImV92Ljp+EhQF+KZfrq+U1mZf7Q2rLTL3JFYFxLk0+LJZ9Y4j
uOEfzs+Q6To2bMb0HivFEhcy/SOMsXHbMa8WldgSPA+URpmBK3eD/XOsbilE/VGK
nBWoOIxwHsCGsbC0/qw8eS+GWIiSh2KjuDMtvOkPTHWWrpHTqmcMjA52IZKcoYUc
revwdbe26ZhKnmdCyXZbSlRnK2Bk7NwSHdfMXJK6VtFzsscuGqxnuX5L2uGvyN/o
8Vr0RBE0tGf2JCOcnVZTJ8gl0gZ2LrHcqEFiQyW3WVBQ3Q8gRWF3OQYB9+L1QXSW
Bagf0oHawJdfZXKYwkxnqyaccj/GOPeLSxCtJ3beNAsUsRbz0D4MG1/7QnHEuIMo
FT9XdLbAFQbyrcVE/cg1MUBVp39xgVqrIH9vDicWVCJDuTNYjrlXcZRvazUOlTO4
//KT4gGQbyln/ZRYJwyeGLZTQuTOR0ydpUwMwe9v6LQOTWngp6T43LGe64W+Bthk
w00D8HzEFeVkz+aIHOxSJp5QqN3kG0ZxMZublh7MoPPKqb4riRhlWvXMiU9gBSAJ
rHqNozeXLxWaFj9XI3OxPRf/DrrYkZTuHArM2r5t3jSW1jiBzRAJt3qjp8CJ7+zp
kpsgseptvz6eEImenbLshtchbGbtQymuw8nQDJuBnyvEI7OZh4U+Qatip9GoOrLw
tEurj7etvPuwkAcBtL2mIjS5l2iS///qnU3CZrwHZPjcxvNSIapYueBJGPvLYYqj
fn90DnZpD4h1Ji5x6ueOyBLBa/E1LiXlTZzvVDXSHod1UAYO2Iq9uchHYvWX6v3f
XkWDWBbq8TxyKZkXaUYUEHTRYg7Ug0GRw5yinEmVeGaZHwgriyhWAjSDMNAaCYj3
ZLu/XHIvuaaP9IrkuO0afElwybT56zlqOlPKjg9MN/Cv6aEagucb5I+zNtc+3HR7
pU/CTurnSqIIs81Gtp/fFk5y26fjRtJYKcbxCj76MMsqj9/cCm2r0y7Pfbia3p+f
LFUbs/F0mF0yW8IPTRRjl8XWB/GUou/gDtKvCtEXnc4Z6s7/B6lVIjXCXDfxs/c4
2BsE5ur6zRW/GVt0PB06F4I5uu2ld0as1XEZKGr0N49bxrN+ursAZVIi2vy8YVoi
LRbqCzp7DRaIJps3MY/i3RqMHGK8zZb3CR9u0JhJqC22p3GgF6BqLU7B7K87KSQk
/Y/1trXlA7574HMY+c77wLWLATjNf8g6uXbQHl8ThCzjDjUIStmKtqGhQX1jsixT
2gkP5GfxbWpmVcyPjpcgw1z/5lRVzQGKfJWdJBeguh57P4PF/hK3P/HGDQZ33WwB
yC2wT+CDE0b4DtHjC74C1EVILUKEPHEVVPsDLI+jXHKB8HP5uQPgW2M4bkK12mCx
O9G0l8ssGFIxhkE+LDGPyVlPoE5y7qjBIp48hVZ8XEEu8UzRkRW9RIm+ZcTm3aeY
bbbJkrpxdcCImDVO72IISaTdCfghMMI7xNx7hzWxgLbwu58TuDXsIUFckyN0DqFX
CgmdnNF+5Rc2884sdIc0kRWRP2rzGIrq66VDi2CgE0R7N1aGdCsCJQDbu6eVLM6E
bDiOXA5mxJp9FOzelR9N59RWYKIIHwy9R2Giv5Bys7Fa4hkXgMTSgAQFdEFP+Yu3
movOXenbGWvFZD1TlEKvLp0BlIx2cQYVrjUrrjUQw/q4Hp4Y9LnUrOINmMSUHLw6
mDT9uOw7uxaENSSEuegEH22q4WsxTNMKUe3O/WrnUwRPbeM1HPyqZ8yJ2sj8l6eU
bcwygO/Hyw+mM5oWCYmD9kuo01dh2QIPj04AI036+c4/qP/OQAwdFksstD0xiGbn
TbkvmcUsnw00TKpimRck1v0t1JigUYe4k4juLMlmWm38dbadquOhhlhQE1+Oi8Eg
6Rtr5OFQDnIFgF/+E6OPe4mVljUTAR3JkSvQ2P8EZSmP0Ollbn08lzIrtcDSwEKL
VLpjF9k+afAwfGoF67xHkfCzKfcGpRsTPMMLGxN+FRkd5M2+xtkCo83QvJqJf3fc
kG5Ho7GE3CfeOnRUjerAiyUZiqDYyXfjQawfFu2NIhsQEjo9BqroUXT5Hmf19Ynb
Ib9ElwwqDYJYY0v1wbsG8s0f7JaAb9ww1GGxIoYTZG8PhLShJluhHtA7yA8d8iji
JyGW1aK/Sa/SbwLZHAx78c3Qhj7w2k1FyseNRlH2oZ0KuXoHBkdpNHXT/Ti+dh7S
rX3CyXTH3sIQa8bcW3frMcauClDdWAkh7/IJPlRMLTxoKHPNdmCeQDEUlo8PbMZG
WztJuCNZsDaKnbospOsRARqlSfrqqyZIS/UBxSfzi0y405pt0nupI+ZJ8ytUdE+N
juFQ49loyqlkB3nik0JnUi4WfJXHpz3LiF+mXgVrmMV4Ck63qIrIIItjRMCHtMX5
EAsL4uT3Pm42E/9KCZOW3GSD58SV34fTpTCIr7VkW+t45y8skyyQgJYgwk+yVDKn
iikKG6hc8IBwt+aIk0kyLoL0X1cTgKy+/+RKfzIC4fxgFuYnk/9o10PAhdX1NGVh
O2DJ/c0trjk3OYfw45i/0p0Ruwk8ju97ShkO1rLkxMyf1/scbAUzZiQvaGeDpH90
hC/Gy1qQet2kzmS/jl1QVz7dNvLRLg0go78VRo+aP1t9QOYRBYa/xWr6IS5iUnEq
YzNIemknFTMf3rdTVf8e8uW+xGJoaeEtmkIVNyNNxdIfud4eyAt/zGjG+0N/QY6N
Td4EMBx8VVSV+41Rl+DDhPbkL1VxyOzN0U1+CmNE23yKDqvPdG4k0AfY9JKvtvBH
BP/vzX5tT0xMUvbfEpMZA/m1QXcl0xBxEc/37kzEW6cISLIfL0VLyeKBkPmSRv3N
k8sEqlHeQ3i8ThnVkv+3LuwYU485HN/uo8l3hWdl1CrFyl4pX/6HfYLw8Il6KHE4
ixVmFRO2hwyfKtIi4ofhFCBfsvSOCilu0pMHuINM2Vp2ozrRKMwB259PKiHBwNf+
qfbPvZLGvxV1ohrXCoEDDRmN7vZz/mxn/hlXTHWTNxlnRM9gscD3FMF4XA1jcDRW
6e/e/mpl7T2fnGKsT9Z8CV2Wsero1fxLe+xTRw4H7UWYFu6agNi0gdxFUx/p0Wnd
mexeLKsgzOQSqEbaggpJXQ7UGqNLLpx9oVOe9hFKiieHMaK25qEU9dNOK77jgLKI
XWuOw8451OEnYUNArmplLGb2wprJnlaexHqjyQHjPBvAItfAnwJcUZ5RRpF9NRY5
hHHOqpNy8nEwg8uwv3Hg4jVn4T4Ir2Cbjjoea98eCs+khTIziDq+j8oL83RsR+aX
dD3ZXGYkjmtVrj+VhHLxq41IJeqprNxrAm9WxNWOJJ82VR8T53zo8afMmU1BhuNW
Tv/8G4TjZeMDhey5D1VN6ZsDwjPJRh2DtrJ2UI3PmiKv24Zd4OLg8T2Ie+0GsUUO
p2VktDt6Z4HL225hNJDwnTOXJdj90dEEXw65LULusHjpRpC+0kyGhfEwmVc1ZpPb
9mIHncQ93HciEelNeRdtinvlAHdg8QCMgtoB5deZpyCy4l7oLVZ8mOT0TUg9hOe1
3IXvCapUAQL4BmWtvxBhrZ6aiwHgZ+9JIpOKYPwgvmpQb7VzKBJu+mABNeyBgT65
lauNFwCa92P5EhidFxrT9sWcagk9RTQlGis895/W2XBvjV3bM4mbT6yN4RmDNza1
8RAM/6YSV1nR+nzDDw7BJ+DO1rB2br7U82gt9LXrz16cWdYAi3lLPkuDX4iOn4pr
k4N0QRbsGswFVYB9X3HSWfjwN/4ky+EED2M26DCu953fU/xu2zkbSIq8zdTGthmL
SppUB2YRH/NkcL5AeJp0kVYc6kNmQXAhN0xCV31kefGtRaM2zleU4pPe/pPhmlDw
9vaaLgclG8EVzNazCn3GQYyer2xRNL53IGi794BJxIgr+grPWST6GvatgLtX5++9
5Lf9e418FBCXPA2CUJxMQos6004Q9pVWLT3FyFNy96VgAm6tBT0NohXcmNjsu8in
5u/xi8//d0kOw+lAuFrLuMy+Fo8jZVONJ8EGQDz9hspcH1SqypHlSGyVvVKT9uHX
OPg12WYP/7hbiqUMMGgzwVSIx31owrG747g/8KsMSRi7U7uKDdZyse7EaCWkf0N5
jb6fpsAaHdCb3klKTSyN8yGEEJ6U6kLoxTuJCvgFcOj6dPQ0zVEk4ZdS75CK6gzb
ca4WzJLFKvLCWIBaK4i/DUcHgV8ntJyXkpapNnnw3VeYfST3Sii+eK7UMpYo5L72
suZY9MJlUfRGUztWnfy/8OlUjCFpb7uUHWm36AEdIQiQ4Uh6h1ybHCjNUDzf3jfD
SL8O9DONRy2cSbBJKqQlqY/2bhQKj8u4u2t7YNM3L0PBIY2ABObSj8M0XPOJHxCe
635cBlpU/a9OdB8JIA+2OoMDLV33hkP92KD4rSGCazi4vlZlKdMtRFgQ/eLKqGz9
Xo0Ta3fnlISZn32FuUjktoMuv2kC7hf0qHBOFWmKrT7lApvTPGhRbXJQ952FmSDw
IuNikmh6cckXCwa3bmgyf1BfiKEHd6JBd/+j1Ekwsj2WKfJih43aFfy02ZAgKvBW
20rXIb+TQPcWsWlJBZ27pBuPM+udbR29t1qttpntd7pHOYWtfjU+tYWu4bcLyzyg
3NX6HKonavZeGPXJ5nAoAByV9T6yCbiSslboqpCB+OhsfwzHnUh8HKBCMWSlBGtH
d3XGjmHgTH2xn/4dw15A4h1mgSL2WiLkeF/bUdqXrl8HYFegNP2pFXv+uYfLHVyZ
o73f4NFW6M73llUi79LsinKLVA5XdQ6Eb7NlaLzbxy96siKB0I/nipRwEGIprOec
b6emNXhj9tGj4ZWCWgWVaUQDLl9yEcQ+7FPpazGvN3KXd0la+agL84iwyWDIs/15
PD8SiXSmONIuumMI3dqsfRgwNc8HGZOQixe2vevs2FRUOgLfhshy6k3uSgivJnd0
JPIfI6PzGkRR4AElu8V6ZSoJ3ORh2g1hT5W9f2kCBjmOkm1Ckfvkfv9K4q0+AF2I
C3z8nK4qq/rgaycbeCWZ+Jeyu0ym37prm7DBIq0EKQKmbgoUKQLmChOT62bwC7pa
3APGt2/Z9u4LpwVaPhq5wYZwc4UqsYRCm2RpghoPBAqqYrGAPkG3L7lsnYcafK6x
Kr8vqRHmCmcTBNizuT/bw4IPSA9CJMVgmWhgz/QscHuLWEHs+OzCPKCY+ft4gBzm
nNL+gARkEWcQqT/Sa2rev0CvpFMaovl9WSYY/P+ahwEt0ytcl3kDXkxTiL1VVzWw
xC6HXTaDpjYa9Jqsim8LqhYP81+ROvaMjE6HmpWLyLCKcvEj0BYBxQm1Wqrz0Rkw
+9NY+/5RWkB3KzoqG7ApP+oa4aueQPA0GB2pLI1gOJxh7plFuovSMJd4yy5hBqJs
taPjKmd+Dqpkj8sCYduI78kSZfV0/DvqC5t2KaeiEWIG96hlcGNNbYfhWunmaeOL
kVPmnXjZamNKOPEhuSJQaEd4HaW3/6Be0dPKsFCW8I+0hamGHtSl1qv30eSmrCZE
R0V9w3pKV81S2cdjTYdmH7IjeAZl6oewCJkAEENuz+Nfrv6GSnuFbovv8CjmXJ0n
zmsZ5M/75nLHE3Ntn+jN9CEsum2gdF3cMqWLCpKvg+YIOe0E4Z1bFTWIAs1zxMhp
KAdQRKREAAgE5M5C8OOlQ+SNqPrLf/sSsF4wULikbYwqA3BEZGMt+kXBNxCjHVOz
MNWp0u0oL2MdvGX7kHtJMXHp4ypidyCm35EKgbeUyDFTfTdD9ADHu67Biku9O9e8
8iX+332ZNSQPIOexYevHCo6HmyZQZkwC8yEhmMEYDLoOiLq660tbkTZHsuH/7Ob4
V4ijo4ofKVrMKrC1q+Ch7fPDafse1+M3ESMXKXYus7YToeLo5WImBc+GYlNVMPCz
uE05vUt5FpcnP7Gb0e4fwDw0/d6PW/P5ejVyv7b9za4BVElYTlbfSFS90vZ0keDR
u3ZxvVe2MHGrGhy1Rrs+MSF7nIpqIiUDlVetlcNs49+0bX3xayn6sl/66MMz9MxV
cHoYkZ3913EL3TWdYiw9Tu2C/eL0M/FJetbxR0fa7PcFKrST9/X+bR5MnT09Ng/n
OEt9k891IkbvNMm0X9l9lCmsVa/DT8cE4t6WbOWXKUqLfvJyHOoE5x+3uSGItCcZ
dUhd4h2Gh9u0FhS5vO5KWv2/Fom0H5hTyrgSmEb+9lJ3Gh/YdtZ55xx2dalAanDt
nIQQ7WtuClOSxZR/HyjpBl6MD1t8UWMaparkwWM5bX7jomOv7U+CyiAk2OcHeLsM
Gp6OnL2QMQcjp68+hMB67LlpMxbNVKq8HFg6FBsrK/HRY6DeKJbXde880IOkIuVo
lu408qDnPcsXl85jnZBW7OCFovs40P0GvYgIeecqJy8dKt593aH2hMU8ZMhg+9hR
a9sZW4+o5M4i3Ugn7kfyHXupHSOMPQuNm6yr84TBWV94YkT5fU+P0bulViz60ZzV
EtegX4b8zkyyxw3TYSy7tQCXiUTLL8MmQat4/kuaW2fGLLm2O3y3LEIy/yj//VSF
RDppR3uhnPPQ+PbAE1Gammu8EoEjamy5Q4j1X6upYslpQE9Az9FPStBU4y5mRNer
8ds9j2FB/o99QuqFiwvRZGoBxyDYgIq9FrFti3vur3ys9jmFe9Vk8s8DVk/Wru/x
NW/HEvxdZMQ/URlFEuDC+d6cpnJz4z9TpTiDJcnsVTpeC8ohylsvrhgPFciufw2H
c1xrkqzB8+S3y0QsOVWsffx05GV3dlSu5lhTAg1XwXD5wbR9q3FvwcWN5dUHP0KG
fUr/0KNEIufHbCqFL57q06FGZUPwR4C12HOP9rkr+qAg7Moh8L4E46e0O71Wv29y
wSHjp6EMGASc7mAn/1EasZd9Foq2g0gfM2SXZl4Zt8YdHyuv/mXQDa5Ag592aHEa
FGqmbJz1WAWjOI2kbhMFvocqScSYFaMa7a31c9DjSpREz6q7lNNSAITkLv8vVxTE
GdubcN+iq9Z7Lx2jA9TEW+3SHxbXvtP3hEoySmEyTz2MhZaxzxclWuyUltGKPfXO
wE3xnpKbcRmuPlUGDhhXEJHn3ldlpsy1dAiVJck0zHgBuzLqorHlC5G7xythAXja
VHGZm3/WxSzEBgM+lplooYLr8ManHGKAczdqAjJ6pQuj8KXl4LSsyKgCZZlUN1Yx
l45fkwKiUFYnlcspP3rlFwWrDQVnJf7N3LvRJ+LOeqpk3PiSkUWZdjpSXVf+Jsvu
QCLohj64I+28z1fWyOF7oLSqJ6zfGf1MXVxkV4VIhx9swexd8r5EvUgKKwbJlzku
X8yK9/LwOCsOE9XPWTM+tiUsAx3T3Lchattcbu6QvSaMdwddYGMXC/vyxa39faCc
5+Tgv8bZwKmg03lS1H3A27hw2jxhvvXfC8BrUww4YY+kpbVN+TRiPiUCVhfYtVzs
Ss6DFjsIpidPBMIA7OSZWGDuBzLKXUlpgYPGyRiSp2LfrNjO3aLXfVkU4mKNWUrV
Gk3bx25DWXuixfUAsagJ8AUcUSCicQ86RgqnoGplXB+L7BVueJXZzTkxccw0et1z
ovh9G7QvMOCTlW29KASDlAxaQgPJz4fDIgK0RX7qLZJBRtpwQPLVGglRpB8rteGY
/uLVzkLXYIH7XNCOEXDYtOkpYc0Bn1nE4gdCzdiZ8AVe8/McPd8YmRmxs4Wj8NIn
TEMoSlNhvnD14QNxmHYi34dLOyIWvl3bhYgBrFGG628BWmdx03a9TZrejot/i4ih
NO1Z9gVvWaGMu/FVaSDnMYROmsLj7JSTbh2EKw0NMUgv8P0MutNLfsBvcxc6iNAm
UNDfmKWnPsNevmxGht2alQXyVAgfb5kcBDYqXzzvmrwtzkYODUpxFdzLbSTBZ8qE
2JW94pBHn1HLJId4R80UAHlDyqjHm0LAatqiW3LGHes2JvRxtCmoknte3B435IhE
zBeemJnPpVYcxsqGcxGAWGmNlNthSGOyS43k9VrO+xGdoPjs3alPALjBU0kkZYmJ
HE83kO10Es6ud3cHt6ilih1a0og2mauMUDGObLYH3RmhCIR8k9G6EDylpDSwOg2c
bRjZDZrUPV+yXFOt+vLUubOfIVUS/lLiFqB9n9ClrHjHdyyr+Q0yiiPLaFbx/OEU
/Ju39HUT7J1iYqjavSvfa+OYE4jQyUEt0DKJzpWI8t3eI6ouXnCkgd4QeQ687/IL
wCAjVR4B2gWuvyJz8Iot7GZneWpLXCSJvt8inTjBmO2U3Cnt55upzhuD4ngAKzfH
vYnP/YYcSEX6Qd3RJCjGUTtE0Xfsv21bBGvW7zRVXablWNeQbafzhSqCp3CPeNlz
QYYmp29BAxeqvP5sepwr+d8SxhkTW2hfYutypLeIQN2KXqGN4qQCtOf7W2ugTfYV
zarJzI1yh9Q5MD33mK/wr9/wanaL739GERu/a9lKCR2TGtfrLEd5pMymdblWpUq7
evRao2RRzmdWDYATuBShhaaTDCn4se+IcC4h+jY4ALuLenLAGJ2VB+aDdTDaTYAg
JsQIC/z3lYu4VYc5z2qewdnWN5/mJt98i43d3l9QL3eoZUpOWTpILMwq4Ao8MO14
NJllvJYc9rXuCATVArVm9n6oxewez43nwVnrUWNmPA+3aOHLMm+Vij+vBis2i/LH
gl2Lumr9tVcmiT1zLQfxHpdrahwB88eMwjFyca88kp4PVT7mYMDK+VpE+VmvdxEM
mKbxR1BjC5LNDyGVFUfxJyChwVTZVBFhclcU7rqZypgSzNFwJKN3v1UIgEtVrX+5
kuOMucMHBSp7aAf2u24x8tVvte1Ui31ma9ObT5oFh6PLxpU5wGbkGXIyU0/KsxoG
8KjyaQZqMD0jsJuUnDo3JVyj3UPlmJ0izJCq8oiJhMQwN2vNeP8oq1+M0PynIvV+
qbbIc46ZFy6uxHboAvu8SJuWCzdJ30qbFEWFKrYOggNYgT1GP+M5scJeQn3XiKPM
uUbKNeX0pxVkS5CxGQ97ku+qwZemPLAlEVt4eUw2Zlq+DfJHI5RXcepSe4ql6yCF
O4kQaGAnbmKMlCov70M7hNxUFGjRPHOuAUyxt+c50nsHv6SD1im+8oN+lsbVtPtv
XqdPb/XD6uZFuLxuHFnYB2GWYSxVYVxUfs1g+4zOF3YfZSSB5YLf60Br1/gX1+7z
rI9qv2mc1vqfblz1F++84Hfop4gnCd+qYwjNrS+FYIMVpW2VyASIPEuZW303tr+K
2ST7QSeI7hYScfWIpHD3T2UgrCsOq3fjc/gpZS/KOrpJhI1dR5ENKm1In38WdYH4
jya2Zu9LV9BNCkiR2ibdu7tvmq0uXtRZvhaLepk2NWYkjopS1Qh0rV1K9OpCkb6f
kQav9fPy8RsQwYfBp86cpMcX05iZ3caSCEY0KLQN+flmn+HQrE3uOvzKLDf2QDXG
wHDhSKHZF8zx5U4E0WI/N32K1LnQPx+fCgGG9nwo5rja7KiRe7jFpp6IBx+jKvQI
vxZTEwoYAfW13bI+jC395knALw5NvhgZc0u5LjNCoqhJtQoKGTpG/+BwaaRAnXGv
0zDXJjNbNoW/m6lcR39dgTftz1rzV5PtobOEXX4s/XzDUxCcEloZhktAJsaR7AXL
Dcb/pgEh/7CkcyXryv5ULNStPMx26NVpNrMO0gPysrDEA8zwMl9/NWH2auPJdZvj
xQ77+e8GM0bRSufOt8bu09yZJpNMDVusmqJwgSi0tpNimQuc7yf+2wpApaVRDlw6
U38y07aMePIJSMLKlvF6phSOoTeD4h1hbccM4IJiyWAUsBwAzvW/XwvQFb6so4cM
WcguoxE6Fa/eCcjNKSDSsZa7EuuIbR6XtOYTxk4qWgKw0Ux2HaqU/kkk8MAlkVqa
y6YmKXM0focakq+8N7PCfZ0L5zT15jg3KfUyCA29pKFkWepPph1OrnJRfWNq2iLk
iWTB0Up4MhMv3COAPRrRgfOi+okisNiXzwxuVpqhKUNk7B7UEgBifdljPtTNrgnq
PC/RjnIwJdY65QvxlW8gwXzQOLDrNn7qcYNUQ0ntXoDxt6+8L6d1N3nb4lOvXN4b
SmqzptqqzOTAfcHAzviw6QvRCC2p314maedSWOSEsm62RAaWYxPuMpp9x8MiV5o+
7wUko41BtCDU7ZG5MAHhmxHbNbKTanqLudhEo5Gnh5RkJzXRhshDAUAbezfO9cxK
yd+IGS90C8KrXDVVQAW4AvrVTGrl17dagCkC9QQ8/xfFVPm76l6L3kLqiqQr0vk1
1XhdBcws7cCawjAGY5N2jReNANouPOSqi4+BCHGDBS6JUaQiL6K4nJBx9+RbbQ+Y
PDwgPfaQn9obWW873youSkqRyhuDQh93NeR9m6lGSl0TQlPyki2W4YHYv6nG7GJM
eaR/MSxvC2SFZsUIWuRBWCo0cwhQGtwaVJGQA/V1Q6Yr4HTnhi+aZBcw31vyW4i8
U+GvLGG27fU3aSZU8hTvTarbw86mUp7KRmKUFVXzwmfId/abDx2yorxw3sQg9mP1
moSyMSRujIjXWesbckL3avOZ+2u3Vk1DyK0wzM9DkQp15odwHKnR0eTykTr0xYE+
ADrw99+kLB3uqTNsYIVg8lIjJre+LooOUV1Y3sV23e2BgDcRUOGitXkdspmjMLIG
2sC4rkGpMKxT+95Nxy7qFc5alRG/hybdJU8u9QP2CMVZQrKA8d01bl12f/uen66h
EGZ1kwdjr+jlaArLkqJLbVFC1awFAgReb6W4C3rutDiIU1Mfu3UKewMMfNaZo7l6
y0vOzDrFCt1zBDbFhcZGidYldPbNMR8FytYOVE6Xd/hbxOyyi+9n4eao0DzwAhVH
CEvERxcr207C7wg7YmdAXKFzicD6IMknKUF03G55oucUub3K5oqhwq68vegSwrnp
QJjMvDMIGivE17zSfLAPnOItYC1rkktulrf6Jalbfyb/67GbEL7/EhvqaSSp5HX1
ZYVnupVqd9Xx3nmfaYrjCJQ4q9brMraeuOl//l3sy5ChpV1biJH8MyVhsnpf54CP
duFT17+Y9LlKm84V7EzX5z9b9fkrkz/pR7dds4kzDSGkM5CFICEB+1kYQNPQikJl
+z0UZJiCQEVQ0VxzhPU7Dy725L0d2Cpn5OiLzJfzQtxWDOH0UXw3gCMyyP/tsUfx
vhe4OJMHyec+bO2KcO9ZTckeEj1LSxQ3QpiiZKpIPlK4/JVw0O2AcO/3sFQDwzoQ
pw+uLVnfM7klzaSFEWFY0lr/YMvL45PIB48d2ztFHF1FqRVQxGfRugu3KfCw72Tl
NCtw9FHQG6mKy9bP7eYVY8ogr1Do8/F8QKAZ93xc1vKcMOh/uN5UQMeFUqizn+4G
or9/Od6/TGZiaxbE8O2nDbO4QeKzYZhXdknE7tfSnW4lYJ2ihKBKPGQDFyX7X/63
mh34ppIO38+USCEuTlUaxoV10e2zL2IGz5t7wi6v8IDFO6TPdtgj4pYg9e32ZRnT
mxw6AjrxN6V1WkalLmQEo9ybI9VlOkXs3RICQddrcuoi82mAyE3071j/BVbWi25l
pG5hweh67CkkSgiWE28gwXNhhEOuwcml1cpK07owVK+Jd+W0SLKB5H+xnXeWhT9G
crlOX/5fuHuPtBaiTknB336W+xTksqWZnVt5ZeH8UuE4gPFspUsgoOCZnysNFKmc
zZ5tK77BhWXy1GnPgcv3EGGSq0q8hK7hp7b8QfMjW3jhIirrfFoyykSQfEOVLp9q
vDxwMpKjbq8ACszvMINQDt9V9g/MbmJbP0BJldrUo93gqv4Bickbnzs0W2t6oaQ4
T6b49HEc4cev4JHFcSEu5JftUes5Rh/GN4kpOGeQPcR3RoGXSmw/L2PSMkZ7e2In
SJ8L8ojjFF1sINyRLfSUtl0i2u+Y4EwyMqbSKnLsANaOnU1nZD6jyMqwkqHfBUTA
9o/Nowqmarkl/W623ED6B0DAduyGX2bQaALbY4uwP9JiNy+lwZBdnPfzQWRuPSMl
seOmxwRSeQG5ndyVmfkGMio+pqysTJ8L1bZtoV9i7QQ03DUaNgyCsdJToAwsF+Yy
i6+ogoS+RdLdhUWznTheLUrWYs/w0oWaKMOIYzvK4Y6oLNbaE93RUMc2acNEWemo
f27AjGyIzaosA2xfgzRBPYsyilWXbdM57hIzQQttRnpnGbgTUMpKNhaoyLdvn2Lf
Z2398lfaiFZOMt07qPh1vlRO5kJiMuEWo99wiyD/gtl2TVV8IEo8gzww+SZDVEDU
lQjC7nM0TgObjbqWFA95SG7s8y6De7oiFI4Ii9JfIhI6W4/OagiM4BOD1JEM0Dmi
ym3+4rteChf0w49SfhIZEFZRmBn0DRx4fcu9ghmhIgcChpZnxT1SKEY4dd3pVh6t
yIRlhow3FUDSUG6jp7/qvCEaoz+rsZG3FP2Pjc9TqcAVyx4iRcteg8eVXjQsQQ5D
jSCBnU5iV0M9KK1DDzOOivCGlM8WcernoHcZ0k0r7albjlSX90GWPsgXxyYtDuHg
UxW5IauvtRf4mdZgZ/HxdXfY/rryaAMTHYeJNjTSsQsTOSjws1qD3lxt4iBuTVpw
q3NezGYZi7C1YCqV/2LJLGQHcIwrb90BvwvaLL2DwIQUJx1Hgyg/TCE679fJ48Xh
H8QzjyIVp5AVXKhvSOT7q5TLHMSoZOLldpLMjUKL/geG7VALhVFXIHmQPm9EC3J6
wVTGGrtJ1+QZpJ6b6Fx9eceXxJcdtwiP5WVT7s5WMRTu5xh5QKpvNLCWCf+g/v2a
nSHpL+sIRm4CfWdeEe0K3+My/W7JPxlzub+EpBjBcJAzg0wu1k1uKMSJSjG59TJM
g7U1db/OjHry670Czafxd3So6HjBWmn6XZP3nfsf6+dtKEqvtGgH+NYGUSScE9v/
TWhIRekYhKNa/82+RCS9MXPtbF5kNSDb7LmFDAgYNeKeuXoDeHEv/iES5Y1YjkKT
NfMjgo5uEQegnJApzfDJfbas3iWODBMfsprANOKa5VX7pSoCc+2/VFSH4/YXSUPs
kMMm2uLCeGEb1AOeXz8zQPhBMwb/5e2ps9IOS5fgXZNxZFdBulol8rDw7BFaudPB
eYVlLH8esz4CpcT9cUA72dXf0fXDuiD6NeAWxmkTqJMdCEgNx5VTKzqncgkzK3qV
UEJHgC/cvlpHvyGUBMZxqRy0PlmVWz8kUAabRT6BSjAXucEy41hTtV22nUW9JGAJ
ULyc0F1YXaWYuOwBJE3ejIemMLrEo4si0oPy1AtRWOGLhLSSS1rZfmPy1AGT0IB6
aTpDL1PcUSBh7Z+AxIvOjnzvil1ZI+2xKOmiUdkdRGAjlQ4sdHMj39stdVYnGIcu
l1Rv6bOKy8NRAGIYCOGihUYAkFl0RY6p3ldhub1dE/Weer4lreIcQQV2Ev05nLvv
K+9ydpdfhlplkId4rx0rYEfZJpcOOW1UrUFFzV7TOvnQUvWszc68IrNTFU3/xr10
6V8n56a4MxcFpRTTt0pYR1ad4y+oVu/AeoaQLHzdK/FjgXrkC+Ibq7ISV/o4HAtV
T/25panhtheQj3eJaUI+BWv+POxQtdPAp5jVRnkU7NJM2df4ZjTj44AzNP1Hcdm/
yVVcPBeYcF/qm/rLofUoPY5whFtkIpAw6Ay1dt8ealVRA1YKzagGOspfp4Jqq+hx
mcG1ZsStdiAyumOpEXVZ0fcOMKzFRc23MghVuB7tq4jNnukM9oEu79+t0d3p+qVE
ZhGyvU7z8eBmI9BUid0Kv90RvMsypnL8uF2mAxSQdBrzmAgq3IMTvheHBoeJ6SDp
kEh6Ol8ohPX+PDQjkVjDX+fnesq5RpU5JeqE8eX5piYgfViE7CFrB91eu++vbngg
eH5hh1VQoKJO3UljZ3Q+ZVPs4tl/aGKJjnduuwEMbP+okky3PzfOYmrk+8kYFqIF
VAmgtOuDfD9c9b/lsTooVav8QWiNwnDuglLOWoYsIlvKbJhj07tLvL1OeuIyvAp1
aVN2E+GOGeZKwbMvL/vTLVKmG2S7nmIe5GvoqGXAU79B9pBf4KbNdsntX8V66S6I
n8L+2RWqrZ82P/HeNF0n52lQmwBfPHG4osgiIms1vpyuAx+LS3n8L1VED/LJBPOy
dMaoYz0+03cBv3yqSgmgp4WxxncyTsXt4RnW9BAQcTxd/grKzQFgPYhUAIWvfvnl
e6o+XUyACl0A7PH5UQ0paT5cuUvsIxqyxJQZeP4E8KCvP1JoBzv0HnU/5UIrdU9G
1i640LjRYuM++U8u6xg8yf1QM0NefiK9hKSXWWJAp0lVVkTOPzWZN5NBUeUnwS+q
xXrX6vTlwVBU48gsvkvEGeU9qFqAcJCVpXisZVoDiLC3YZwpa5b8/jRlhTMAt33m
W+tV+l9fPEpegKpwhtQLHS7nXfFKQuuvb0XMpxEsnDm5DRJqEu7Yjp/N2lVs+DPr
XQ5GIMluNdPaa21ax6cEdXEpCXfs8Nq0ffNqbSCL+3VGsOTtxPP48uNV2SFSsLlR
FWYMKc7fI8b6q3lFSJcHxZmFrsdQV2o2ZXV0NSFoDMDlSApkIImukGpKrdyRjp8p
jMv2s4JOjVU5lNzmN3kZha8W9J2i3Md+d/jStTvg6etz26+xuwPczYXy246plhi4
/bGt0jAGRaFKgpmncQQKTg9yJ6MO596pNRlzbKVFNb3b3jZ1Oxvg4v3AcK1FmArj
p5d0VkOBIIyYgINzCEGtaInOXcWFgfsP2Pv2/cezy9C8GniNTGGxgVRjAd2mYDoW
GxVbkI+nIjmsDhW9Ila9KQ80wfGbuiM7m+mEf6O8jDEBj03lKTy33mV2kLUlyg9y
DVRJku7O36GImcLdlqsIzHJiQz9UVhG2JVxKXS2m9TyanEZ2Gl8DmTm53mSKpFIj
dsm2uKPCkM17v2iv6X6WHPlBmWQkkj+Hx7dQxPkBRYNwmaJJsXXolQZ0c707lnyD
H3mLOe41dVy94hfqj61nLrZPyV6mnWxCLckyE27xYo5ZuImY1k6/7gAhOI6KgqWr
jKZ16b98dJhNnYVN1fhQLC/ZL0u1VmxRB4BSzERaOjSrOYFtNz7xMnBpCE1qxt5H
3yV3ICQYWRXiveONqfZN5xzKnrFKD+3BR0mHWVQeNIT2Tiq/OpiKHRj3pDJcHX/T
HefOs3zqM/WYzaEqeAX/bUhwqYyTl6jVs4CZNF8KDvf2WqmQBkrF7UhWdxQcIXCD
4enGUGTAR8/CoOeIvFSIOPcHhRuxkAnvt3bXOhPDYNMajl+lKUWbkZGoGpyXssXi
z3OXzBHCrYcw8+oG2OaGyCIJEkKzzq1abge+702Hqc8sMJqjfYO4rG+K+KwgxQie
NcO8ldJ9xPg23t9db0rbpa4W5n/Y4kOBlX3Ju9jOr13Ean+sAYtkUTQvAIPSt3AQ
FB6MzMzS/8WSAkZzeCptoA/GfzEbBp07fkVG/strRA/3vxgknrKsiJjLyxd58aqD
fL/x+NYSleAGNvNOxhj3i0MgPkkNsMrPYCZ9MZ5P5Catlpl254BXC7+fUWmKrlA9
vmhYr06re+C3m/M144gcVmevSA3/ckspAp70mAWheeEUhuYIIVpw5qCActPMvlpU
Zr0XQ8sbt0qT9R5lHbn5d1k26XoXXjOXB3flkQWxv7B8vMXhL02LEb8KKJGS3Vt5
++8cv9k5GMQWJjUY9yW+vD8TxJYyge75Own4pNeG3D/sfPZtnW94KlaixjaZPihx
vLMDbaze8CqWiqNZLzmNom56opeZq9Crg2kWkX7mtalktsZ/zrRgNLWcDtrCeMZn
7qEEGvFnASa3KJtsnDqtjD+tqiZlMGtzffW+ADwiU+W4aElPzl+qOD25PouEZLBD
QxiST8rwC5AXLcdqk7qPsLk70xEvETYTHavmqoGa8/vci0efJNvCPg/Uqb2Nka9p
616My7efDYXg5tz8xuehb2wV6HnQbeWJTXmba8agQjtnMAuc3d+L2F81TWgVpGHC
wOc/ECU/IpL/5/6l9hssn8yBtz2D2YzPh0g5VoU3mGUjNyp9Pne++1sgz18B78qS
GvAhlOHKlhOTupaMsbNGE9UbVuhtXJS754IlgX41LDRlqEwwvAWORJGuxs0Rtrj7
FFlcjIr2DDm5aNOBLlWHNTm7ckH0fTWliUn8MucunJuTh1NRwZ8eMZYs/4j8TLld
ZiKfc9R6zESioQuIgSPnRqEzuVGj82QBXr6alk2M2+0eZCemQO75jsERut08a0kE
sPTkxmezTjY0s/2FEILlXVsaIDcJQ9Q5EruJBlKnoY7OIHl/8aZV+Bhk6XUXAoT9
vTP4p5LktWWCZEruN0AT+tTeKYDTE+nuUzB7RVYuWplGOxM2VyG/6lUBA/mZQ2HX
NWrrq+LouNyMpBTqOUZ3lL8bBi08Wz0xHof3Kl937sNmZd0VF+31NFkbFtpLtPBg
eSNETaaU9615QuOSROeSc2HirMnoWUQhct+QJsGj9svDM+OgRR2lsPRXkaSWIzZZ
k934q2foN2wDX+p9NE0W9C1a8Spl+qDgMiMCorIFBj9DgGKqXgEoKwSIVIpyXpGd
LDUqiIR6wlBJ6SqpgoKWCXkKurd7oE1P4l5dVFmmkXpMgqKsdJPRHiTkixwPsBa9
5otUHQw8cV2YPd5vSXTFyJXQeJhIxgkGXwN4fMFRC34pyW+8bPgRbpoSHHUpn0Co
o4fxH0hcYbRoGLsPySNx1oXBw7idb4uPCUd8vEV8jUGwlglXRJ544rLK200fcDDs
RL34w5DQ1HJYjDHa/AWME8yUH501Vtgo9BYUXyhDuH3wkSSLkw2tAPVymFVY+5vh
mzCSEVumQOrDNd+1dEjnG4Vc67mcblAyp7nLUzUNHwDIL8fakAMlmpVNwNOwd5PZ
4aRdXdWiaLh58lJeyA33zlu9qKq/hWqoSi9qLhJCOgs/5VxKaS/ibW0Sb8LZJMXa
ajO2SwKJbny71dtDE7x1EliugmF5Px8gUuMRO8UHLNiW/6asmTEHciR/GZ4PZjp1
mFSw2fz0GNejiYi4QvZtVGIPHkYZhJ5dRFOVz+nAlCpB/ji5u1dGEfmAPIqKNap+
02hMkhxCKWNbPJLYCWGEMZOAF5D9IuNQy/czk3BEE3eRXxx4sjTmGEXUwD1uY/Bd
pOGQEpnraB9+gM3i4SJWaNCLLRFt0iTgpr3TxZSQqfvthBKUDhHqIvNnCcAuiZke
XU2UArOOjtCWtU18Qc3xHUlXkuVVJrj556PjSfzmiJIXqF7WcQe2ShrLmz+fOBG7
h2uq835sq7YSgpyKtm0fmMJnnZ2Tiw02SRyB2qcFjDL1fj5X2VISgcqgEq+m9hVB
OfYwA15awmn+zi+dobIBdJRk53PO/6ahEqx4cvYx95YD6APn0jp9FHuyJ8+2DeeB
vDlNklcUl24M81FWUSlqYSgCv1mqMXVzlCrYUrMtlvH3sfvW7FaZpyp+Q3ye1XvY
R4Ye/HLWjqnjVJSVR6QBJXrNZWhckwqdRFzoHf6gKJy7yaQWyKfDxWk5tql0e4jE
eg9w63ZKR4MQoOl6/NvHwAxK1CdtRPvHtvbt8voeo7jrZWg4aJ/+1KHRIoMyXlVn
OX7dn7798q6rYdOn5hTu01CQgzRJeILNoj+tyFjFOqlo2OmcQkGV2/lfkUfolElG
xfFnXpTN0CaMBg0twfj3MAxp0dowrjcLrXxIzJMzI2Lpn4iQ82Bm3Ukw2EYTFIp5
Pr0ki49XEkHVzpW2SWEMuGC8YkrNa6obj0jMsC5P7uNgwHHBRjMg28mDDyaH94Tz
xbuTFpPO4zCpyY8GD62uT0s6ySrsRMvCxKPdiqK1MZ71dWDBi69XEk7ZZEghoAfX
6qr26hKegBQHnR3Kfwg2yOciVwAQjOUm7Ax40vTDgTue+FaXn+mP0p0HNXJQoLYP
u7UNBslhV+E03MAAfhYEk37ZYjW/+yGPmP+U1r/hUkSfRF+00ImBpfRHF9Kt0EqY
8LwvqBLB1QAiPml6I0jWQ7x3sNJv+B8NhpipnjjWyS7FFKtuVdvt7yaejoON54zy
MHUfZDfJJ2QtnE9WBJRKPzKD/OfvuW8QqbaUR7QDnv2HzfHcEISwe1EhhTOwFuHj
1+Wx6fXQc72siLA2NWIbAcsMUBxUnjeazm16TyDYaKxv+6cIDpYEgAXQkBKz+Kps
zir+1t7luGbP44GGxTcTTLXN+LIhP8SMjaNwTt2AbNvzimIcUTE0yhuZ1+9V+9aM
V+gj59c+ojc9+xrIiMZs6GRVWJ5w52He4dzUzHPQq9t95MkGlkpwz+rdG0OB3tHY
XS24Ux3no8DO2umirs+5lkmjLluF6OIhbJwFDYUPxjZuMXnUJfnejTF6NJkGo/0v
cRMDAU1PqQrzFPFv92lBv9D+DlRevtcibo+HFuWBUduWVzhsAvGSxl00iMB9+RoH
EPqZAATJh1WGrZCPxoWsjSlA9U+PKosLuyYNL1VMrWLnanWRQrsdb2s6lqNIoFm+
Cn5ljFzeHICP+FOLrqdvnGFW7TXwMUVp8dE6HFUS/7CYMqQCEtTgR5jhRmoFvTsa
huquhxZOBiyaxdJfBHYPbV/CavQZyExzeca9tmOpi1yqxVDPgGQMU8vmqS4Rb3/N
lzZOUkTA1g3s1gpCgVSsDGwSecE7WYJ0GzajeL0+9IzGjVOd5atZJlGuKeaGOl8U
Qs7GFieT68/9jElebDqPnOLt96iq18m4/Z7NHf7nlFTFJoSpD7g36t1+dHnEzTFS
IsIu4jqDeSXpPwGSScMpku39StODWASNL+TpcauHAK4R+c7rmj1EPIUmJm2hz/PP
0xPUcuBJtCO4MT3hKOvV3goB3rxghsWWJQEa6s/8S4u2bnUtpTc9bnrQOuKjzvzC
5BcnGtrYqR9dz8tlRJxCKiwSSK8y1KdFg8N5p8zbGLLYURW+QluMbJOMKBFURwky
VgZaBSPmtFRZ+CztAAc8Ai6lj3sAgqjdTtLZ6dYcP/3uoj1V5NVX6VHkh5QQCvR2
TXBUMkFiMjzCUZaPA8KyLwjahQBCPIIInkS7OqyZaOUW76JTXJ/ropRggEb6vIYC
IFtpHnuTjvxhB7IPvd98k0QY6XS7BEtTdy/QnmUNiIzssTAAA91xbidgpBjgDER2
Ztu0MA6Dg+2cPLoddxF2JdZJ21dbbQoysVnbxXTus1Ofz4XVDAaRyAPwMgNoaUE7
TyIz7FlIT0iKUTIJDeoGVSMTv3/ls2xjGlnK0PBUkjqgapTtmCZSvnck5lFm2fwS
rCpIbG3XxeieBlXdGt1UodfhW/IWqzBI4UmfmWLmWUWXg6M49M4HuagZ0E3PQ8ro
PlleHptInyJzxqTWu5HplemodU1kLnBw4YXjRmoJCddUnUQNUlaxduHggeV/+b4O
HCCx6XebUbJ+qMCa83rL5816uQOaAKQMPhaXTyL22nsBrKdzVg3OtisiVyKiYNNz
UcnW7FhDdzWhE0iXQwtDfSRTN0c7PNjV4rBY75hrej/LM/yxOq7jSMuDRcmKZ5Zb
Xeclsb0xy7BIa12LKu1Z/+eebTJ/PPx6rzIvfBWlk7k+5vw/nfNwdTHCpw0HXe7R
8GiC+OVdNVeR58kixqhXCkKxAZUg+QvjlEr9N/psNNbPink44+UVjcuomoSEPh/X
naTFq8Wa4O3U7ewZs6YNhv2Uys6UMmm6zCjFeYoxgSWv78gpaK2OftYvC3Pbrlf1
xqDPG+NbOILAqTgAArxEGqHXDwuAbUE5USPHB9nH9NhEiellJvWEHRcgVlqPopnL
LzBZZAG4VcXG/fzV5lkaBNQobupxlmgmi8gvm08/ZLuLtPP/FcV/Z7lG4aRcwTZ5
tv1Bpufctsi2OPcKEfqF5le9NT2H/Kq1u5MiTfDn4o+oRfBAIab4dPcVUqIdwgRn
qyExlxrIXKb428m0EMBX7285X4YYjiCaQg7shke5ZCQQ+N0t3NypX8YnhU91hDq4
PCjkqN9QBDk+KF6iqQQqu+UuG514/tcOr9BgWvk2GtCKFDC6+W0aRtlI5YzKxHCg
bUNaRqlvpYJ0zRu3KesKmpL2wQQV8vEjP27LWGpXW5M2cGoL383Em5AFmOX+mbh+
6fnzrMQxxknpz1f1rlUF4sGbR2mDR83yXUANuhq00os5wP1vAxkBzYFNOHCfcLAJ
ifXwhFiQWBWQJ2pJ19yiacWabSsqgbK97EBsCZ6sUaCws0sNVfskqareqR64y+5u
LmS95eg9KJW1+fQB04liqMWTPVcyrs1wk1LQPq8BA3EOTVV1JrkEO/PcDZnu0r8X
a05JVXlJ1ir0THLARDGIoGVuXn+GMRqCQiNcE9PD4uVEMg2WTQ3Lq/K7Kk3fvFHD
qfZGbkhNC0V7jHpU6AubGZwoduzgW3WGqe53q5PUayyCCyTLYUFef95Z4NcgTKTL
tP30+d1y/2EXaZrsekcMAEiYcI4GuiYhZhxK/GxLZDvzuETc1U8bChq1yUgJZ2CQ
SxmyAJLfz9Ui4gaRAFuH8GOKLxQ2I5LVkkFLyBXznm1zo0bo1x49fnSo5hnbFSQH
SzTCdpeKHyRZY82JOy35sgfYiz3f4wuqcvq7ee++vKfz71dJDVZ/8JpV3S2yeOKJ
yKfT+es6Ev0KSmwESxJGn50sfYS4jmHh6eYSQJc+/VydBgK08+/Q4jH939b/K7DV
oenbDQFLWvM5qu23BHspyRveZOyYLV3uBCRG4A00E07jhC4JUD3K5JWh2n+EUubH
w2RCyxbrZanj6OVKSwTJ6Yw6nj2s9Weaa/fY5FI4Wokx5cdeLk93+bICblX5rdMT
C2usl6GLwqpsKyyPIafqKRITSFT8ViKkLFpN6lYUKgB6GB52Xauc3mONNmCbqn1R
jCVZpm0XcooxH2kazcXGNk0MKcl0zF+F8AWCGH4Jc6tQU1VKKi4+1R+D4SdzzJXV
pMri4JkITJdyzrKadA3MfLL8QulNjNt+h1zD1KHYA24lWVVrwVrXpKbIBgVOBB1M
ujagaL6pfeKCJiMrDUblxmPsnos+FbBeUutQTlP5461cW4MP9Mej+pCtgiLe6PPy
2ew80rilYsvGbMvcqZ/sIkFzCt/cQxvsJOjNWvygfmY6Wr/Gs2kB4oU9W3SRBr40
O/vIoKVzRfH9Puf0EfZcoBt6HUXigikrQ451iXZxuBFfyL+dYu4eOdp7tzec+1K+
Cw51Tty+WKMMlzq8VmeatUHr9A6iTI+MwI1qI7HF0GXD8XQtDIDlLHmFIEhKWScQ
dC/tVmzX3Ib8wiIgC6CT+NNin093FJlB+mOkWCNGt89q/ezbbQOnemHoNN8QLAHr
Bbz8e94Q/Mi9+3p2WfbAlZgPOy04coZr09le6SyENqtYNalvbcxhfIhHXjTGZdkZ
sCbC92AXsIKOZy2H9ZKOW3r81pWvtaxcPPLpYwe+H1hkNwjW+c0WzrWA1/F4A4Xh
qTHX0hXA8zRbJ703A3apR1YR2tZ6+mPY16NWMNfIK+DIEHN0zFUP52Bl7o8GBicB
I7z5HO5C+dTGMnSZSUW82CpZNckBalyofNE3kpe7ugBnvD5XdIM6DPktqIl8MHmN
9j5MLIP6DgCJ199lUazeCjHtdcvrimBQ5jB1sbvvDr890mHAEwC1XDDJ5ZSNGwvQ
VcN8RPZHuCi+7msgL+c2p7pE91MDcc6zS0lFP/zh0uNEN5vlEjVw+wWdlxWcEBVX
9G/xZmrXY+O0ZYxpa/ktR6yXijiLz13Ehkqqx2XtGwReE2eoR794gtLaoIp2oT1P
qMwr9LjpH3yLN5TnTvnFrVsQueJCqTC4CiGdbPuVYDbFLqqnxC31V0N4Z4VjXhZc
c9xWGopana4KGCZWtv4KjJiaNJEqPQHT1nMs0ghfQCoKDwDFnFb/mp4QJG20kJnZ
AMp7yd5XwzoASA5jYQS1fBgbpTpyY+XaFmZCRKPIzKRgmZhCdo6dXhIHZZw7LtSs
b8dghdAME+pKkndDFcS4ZDj5pkejXInm81k37YJbjMFfU5/gumfGmFPdH9MVMNuM
8Cr70KKBUlQUKlar/wq7hCZ+H7AWgh37O/ffVWGavMtzG1iXngw9whgaZLLDXZwE
JAijI5b9wi5iIPY5dhF9MgdQfG25JpJd0FRcVd3cpVfPIM3UxGPhiiNTqbTDyc5r
iAj/x07ss/7YatQ68scEnN8f+oFulqmtcOd6jbtRegDtoulFD4tZ7RPq7i2P4Fh4
zLPVDG7fOXyZwVBZxmYCovFHNeYPqjahSzJpgVajsRkvGTZvbICO7u1FG3QNR499
wr0MoLQprGLOftmnjWpelKngUqQys/RczIchdZA0qfYquab51nqQOZv2DOYGu5Zn
T6sAhGVsYxfHGvWon0Xh4bJNorRLYQMxlqhZ/965JaJohkziF9j8qyRVWqzbV3Ht
2Fv3vr0Fj88+dCgK0Se/Ui/1k1BeYjNGSLFh7QRlyksJWez47OOmGTjDEXVd+LNv
u2XGnyR52ApnZd9uS4zRmEm11RMNJhr0dsJxjTSF7QOzqhvTEugc1WdFzCj8uoU4
9BlM1q5wsGtYmbLbi+l9PJHGnvqeRsX1jfmWDJSP1ZejJTwDhKBNKnVo4WzzMQ4j
mgxuQI7h31qS2zVYFAqBvoivhiVWVBv8xFLpaDfP+sh0kD0ddIBAfGSqwCNJggQ+
R4VvpQzO6SbXehLhQNkzUDs/SqLJKHtcDChuJmUIL3xs3EkiyorHMaZrnEAjx9OE
mhqqE5yjuluqQS/tdl5cvb7rHc9Xf3WXQkYe0sIaY9u9cCv0/Re4Gq4ln028NCAF
TwNZ5cu3CGQ7+RVEblDCrovDPQzg4ir1os6nYtnX2TsmNT+ov7vVM414JDY3vBFt
7Lz3H4E0UAVY4/XM1sgQq0u5CeLl7Yglfj52c86rp10if/65o5WQjQIGosqtndXb
6ayNPl0To5dq/R7yOQ4DcnJyAFDi8OHeR/YbYPH3EXn4eqElCgwvljHSlUi7J6fK
XoAQnjeWhUly/dltZxXiAvFWRSR1iOUyS4L79xpJ62wzqlbxhSvhrgcUS1ZWOx9z
X8mwC6siaZpx9ZQcVY5SblHvJ0/Vjv/HtC3/TsD6fG2LXYeegBUx60cOPfYMSBFQ
KP+MIlp3XU82L6PKGX0GP1wl9hMjFyx/L++XozEDQmgjD6xcfEY4VI1l1zW1pUSP
1cRSXNsTACXOaWWXYRBASsaSbhdFTnwGeut/uUiTDC5tMKbsBYc9fZrDiNPOOwfe
rWSS/V9KB+4EBPCess0oCExxPhWBwnVOY5IUarR2ZZRXLcQdH8hZ3TTkLSECDKQ+
uQqZaIkcJx5Nv1ELg7uWVr5hAgiqMQ1LqmYV85X+mk0eB208vR+abvFWfNsRLN58
XReN/a8E50CHQ1OIYdeRHsk3aV11vOc4CniXtb6U9BXMH6uU8o3EM3FX771n7wxV
8/R6EqoZNnJk+G5XglK8nd3427S+RnsjCqPPYE1RIKxdXld/smiyXXtGOUkQq6wi
pFM2/4Ytrj9bZhdwWzIc3vxtmUP4yeejnIVs9RmhE49p70MIgScHuwV4Oib9Mtaa
/dcR6WRya8nGMoCvZPYOVjHlqf97vAY/QDGWQhPqYosjXzXM9OpAlZ3h5iumB1y/
cTJ9LJd9cBqR85Ig9C44nmI7acBqe067klzAVG4HO0A9LYooli5h2yBSsjzzChiV
82vvF1d6p+KQcCnigzu9WMakQXO76QkZi2HDJWXnrVMWKa2qrZbBqg3XN5R7nUyF
6a5I4j4N7DGE0CP1PEvePN/toBspr7GKhuC/3+uXiPskMMJSs9BfdvHLpEDOprx9
lAp6Fkqx+n/HkF8/awVZ26R58ObLDghsmeQuvMxqLz8Z0Abo+A4xGU1S1ct94SKc
xx3vI6voKn+IMkI3CI+fVem1H4xKWKxEPbFfiSZW+eTUAX0gCDgACR61Fd891Vzb
gAlSq235HmeEj4wxL9G8n+RYrqpufeNDnuJBD9lNLlbEAVER68khpDk0gPZLrftP
6qRPFE5kkzvqGB3ae5m3oSaOCYxehGgfqijqLDpfr7IX3NjOpDtnioHZJVtl7ykV
R2FItVQEHSWjZJBuCbdtbVLVCybUoCLnf5fUHgKTe8eJE6Q0BAnSh0oVRdxS4p+c
EJoETp1LY9f27EI1WbFHVIeBzRaGzUosvxAI4B1GApi7ljjVOilM7hgePg+RirpP
xhyuUW7JA6Ky9u7yAgeG31yXBASqobOMe/MDQv7Wp0zXc26h9AeQFU3VGSzHME1n
Ucp1NOKnesfX7FFw2+jF7+mbB1P1xE12t6CLXNrTYIl/870nEquTfSI6iG0bjoXz
hXXAktn0Lgckhl+TObjeRlJRLY4bPo1pAgVQv0nRGmpvEOhEGqq1faFvbLDwemF8
hdcoefKD/WdtNxrKtqsLP9ZX3hN1/mXLdKBckyjC71fRiWB7QdtTSXoS00mY6go4
p4yX+7a40P0QQbs0dBc3wCHif6x58HedODInEo1JzSGu7vRvvlr0NZ78ukTH+y3H
EyIqHOCcoroVuG4ImdOE4ZdFljDBJdBGeoXwzMG6uMBnlCbDsvOZdx5m7QEqhlZj
Pb7iiw53ZDXIoeWfoWwW4bY5cnwGRFdOf34yRAusxjMMHpey1NmCGNF4UZimnkIE
4JWu6+3i3UtD6mXGFCBUctws+y8FFbBL4dUkGWGPLgOu5PIeu7sqxelHGxghe7iL
7O9IKUs1YTwGa5WtI3U/aW/VzQJvo6kvHpxdevtL06WZzMne9yFc6HPMoOelhPZb
sUwhoYoamSDuVs6jjJKq0dO6fF4h/IamZARTn6TiWayZK0sSCFFSLt7QQb7TcvRo
dtMGG4JqttbcW9e5sQHcEC/5TFKUdUDAJrauXSZRF7l9K8IhVZGDOMPjBXSNFq5x
4fuV+7oAP3QCIlsoXU9IqnsadXIKneO82/TtqOf516xX1cYJjebIj+2o334fPBim
e0X4w1raG0/xXKujIuRbi9FGPWJkfq/j4uH0G60WXIQUWOGWljFzQlVVnwybPPRw
+oVYcsM0O2+7gzXtC8a2Z89c1ySMvVL5QmW/kjuYnKqc7/2Chwdr+uNH4HqJOBJb
abuwg436WfDegjt36DRgUu8e70ZqIFNQ1uf0VC9ltc8TbBu5NZ73Y++1dKQ1eSB7
QQVGDGucW/Ko8J12qw0wuqHrdcAHdu83Bj9XL0UhpZePqP1xSXQpp2Gah7wcj8xW
LwKnp9bYvtfil7M4fNSWZvdjmGfbR9DcTwhfkqTha0GnL9Kw++srPVruJXNcGt+C
xUr2X1ajIgTtpC0IX8iEMTRiWTNBE5hgH5SuMt6iyzkPJ9Kws+pNlu9m3ap+5EJ+
7gLF3k95ZdkCBrKi8DdGNVKNWKqBQ2IdRsyV7zAAy4/oQ1Osz4BMwl7wniqDOFBH
VRx3x6YDa89JnciCORLSd/pVXvYUu/FB+If9gmQLc71AaIZqlW24WGYvTf7KjfFd
Hx2cHJTu5y6CySyU2QAF/tpxGADLB5AFgKG34GiKmO3uQZe/cYymIFYIdhcGajYY
MDVGamEyZJ7rKvVsmU9UoqDKUPjXoS3WNXWv+BrLc7rQcvDGOJWmH7Oaetauh5ft
Mc0TwQDAvtZNwDoTZU4wAQihEB0qIfoI1NEtuy0WWbyJ1T71R/oQ2nk7g8FPKU/+
u+UmsIWK7Cv72tukH8Dkzzmv18W8UQPxDbn3ejjWBcZg5MQCv0qUWjcdXpcLlR+b
ULW8o1CdifPSaVKhieBuOH/Pr7u1mOmwxPtoQy3FDxTVm+KmCmwgAi7M47GuF7kX
5rPj/V8kGfkSX19xX0++Wg2qri2+x6GG0NUKXA9eCKbh+jYfFFEfy1c/SNH9hwal
+NkVZImsZOkLIi/1iNqqAYabT7stVoGcXjQWbbWZuQbjOJTmdrfKymXyBy22GRzS
9zY8YcDw3L2ksiLh6FSGPjDQzGn+TGLLMUShYLDvTbEb7NUWDR7SJruYm/8P14fv
4y15hqn7ebDuCNAndvBvC9NF+eN42L1eOa69sP0naOaiYJvWdY61C338PfLStnox
snndqQQskQYqyCIvKK2pht1v+dT5lgfFEjP6/kzNwUAVR6p45xLfGNHfDTXlIQap
iaO5+CTtL8Bs3OBhVTAz3VOgpw1q2/NU6mUVMrO3oZZHnaKwlkSq9UnlEvLUNefT
zYCZZ62jp8QPqX2vKn0SsvTgeLl1XWT2hHor064Ljq7Xm33/WTr72/a5ZK9LRClV
XilYm6PXBchGZ/rvm+5/SK3/WBTUgNF6SYNd6oJMjqOcK8wxN2VgxksT01Gg9jUI
cfYZEeheBiSxFiJG6IOnhc+5EwR3ZiI5dXWvqCd4jUR3vA6cU4K22Sc9mmfjtEaE
XD0kybJd62WRHZfSYxV+SEMG9KQ2KPtBvLVv95oAFuCZW+Kw6cdYJtT3RnMnRdNE
bpLg91lDUzCJNI9r8X/9CX0Tcr2ploikSOk3WUSBoGz1mkEbGfZjU/aYPZ8KXGA6
ZsSofKtT95Ms831+rR1XkZ7tZOdu0lbPnH9tfjtzL+OjOk/sdSrcoHqNQsisp9GY
oGQ1zqaxHT7KjxAE3P/t7XyiVskSLtsNC6NSdx11Vk96vFYa56IrsZoXTE8g6XPB
p+OfTy01VQEQveJv3mlteT4cYKJuYxsmt/+yOJ7KVnFPLAVYsJVHdjhp9VvS/gVS
t/lJE5HPvMpJ/ydAo3UMZrrWZlbK/W6VwETR6MfGgL/05EaOZxWCo4BA7PLrKEP8
0LSDC5Lq96t0TQ5utTg0eUSq31RPSKt0JVlh8DtFkXswWucgIiWQC3KRSsJ1cJa7
fifW0Xe6zZJrGFeR988IhUqxGFExUkGny03FgPAFlsQCw7BjF0JN8dvNUxRRyUwA
sZNNhbG5C/4Au8/JoyvgnsUdny5MMccHKw3y1n6f1mPr7P/4dFf52wZRLzJUY79q
6zagBGiInEIJnn9o2rpirm58lEzfpLcV7ETJedrAPzlcfytTbt3DPGWlHXF6i+22
HXufVU64Ln7+3C2GWbM+reRCQAG/npiLSu7k8Xuzv9gIl/X0Dm7D+8gfL2FzRLCP
EmDP++NPytAhYjQ1ArTR1Kf2PDLjzwdIgP/oS78wFrQEgJ+YkxpbMIQ11ZUfRKa+
LAtRhF3FJ/fa3cqC5oWWkmqV+ssQ7kYoVCKjNY0xkd/+l/vOkQxsFBEEWx1DP9jz
Yf/zhyG9df02kikcAz4dZEmJii6iE+LMPEkJ1da+z8/NXQ2CyInAjdYXZfCjSB52
V1PxVhhroTXFy/DjDVumoHmwqLe3reQvZnhDzarR+KxtGFfpxm1xwoISGVbo2Lly
kt9q4mvZFXYPWK0NGrrwX9J6074Ze4WD57e0ybT8OSQD6aMxQTSfPel2c37q6+Lk
CeMuz0BV7YhL6bGQ0ISHWWQUGT+HlGvAUOX3Y2bTnxmebcm/2wOCPd/cSORWBu2O
MBwnTiWMIKaChUp5rgoE9pqhzlKImxlLSXaTDJpoM5EgNOMAolajP6UUJQWMXASY
9zasCUJYDfSH8iALWqlgrYupMAMk7B5anFOvFKXQlijBJCnd/cY94FjdMmvp+9h0
hzpRz3BQcJ1QPEYze0LTvhwF+M9NbEf0NYBL6OAKU0zESZD0iJNPq0QIp4BwNg6a
7KXAuCkw+qXV8tV9fCFWdFXqpiJ7BUnZGcviBkhjoG66ObEoVTmnQ12+XQpVN1EA
iiCFV9A/u+TWHBPDAD8t2Ig9m3qzDp9aMVyMxG8Cmbis5INgXeiVsEpDADtLW9PI
ha5alBXOff1fL09bKmLvI2/TgowBhuCvqg/qhWgIzYdECXdV9GP/cX5aJgSUu5jY
mg0X7feTM9TM3QubzfTK0m6YJ9KK1OVHjNdOoTxwT1MIQ65lyf3PeI4fTUR/hI3f
Re2CjvuOlcU+zu45QSO0rosFNab4sI2s1ABlvKprMvgQJsQOgsC9xRSys6mEsz5W
/AH+mMTAu5C8h/mOXOOuyfH3rYjMvc14ecZorkkP0Vl8rO+eKKvsTKik12Zj3Ylo
fifawridpj/ydMbWuvPpRsSyqfuOc69K1SdEeYhQAcutc8uzIfO9C/zF2KwFo4Ow
mZZ8sdPgA2pmoqJxmrh57qMl//jVMRQslDs/n7zCEOOxnr/8mob8MgSJsByP+1+i
Qy2hjZ81ByD+iu+eus7q7ycqtPsZwX5XMDqfCk0bXqunESNrBhPeilLXg3i9Cfm8
tfeUr/MhQUOdv68Y6KFGBhWqv/bsKaPg2UZaHvUh3fesDr7TQpel6+oS70o4D1Nn
YpyqVNOX+fvadjJ6SbzPHCf8RthGJPWp84jB8Cf28WIOJUR5qhdHsXyo7O2w12sg
HeRrUVyekNkFpye6Yxqxdd9Jl2T1FuNpkJWHXBgo1/lofxwrTgmR//ZIAnO+eGpm
BAt7/nzEbV0S0oGD6YZjnJjAKIPACgXlKvWjf1cXUJcblsuTTG+mbLJ+7J+vz6D8
ayxWGX2zt28V6ccG1uRHKr1k/h4BhhJAOp7AYxl6pkwn4bBqzW6Q8J6C9nH7PUgO
atdxviIOAErJSP9gSwpOLBWdb77OIpzSy1vks5qHcPwZyERc6HS1zjHMqZsXbqdJ
pNPevk4q+hQddrslSbx6R670Z5vyYTvxeecYaH85CYz0mL5xhF424aBYm61ZGGfM
3D6jgGsFewLyTC7eRPHmHkeuaZ8z+qHxPK9wK0vpOmI5uOv0sLN8+YzrHwXn30Ap
8dX3aRAPSqRSXszQO3ZiRvpnmibc0QvmiVr+TDbMLe59z1p8gpy6Y493hlHeWNSH
RnRroS+rE9ajAEIQeJlDNaIhdy4Un6/XaJGB2ozEDXdlhJpb0pC5ZDWvWaSG2TQH
mVv2f8lxpBLpzsOQF0B8/X312/TnCTc1eoZmjH8h6bkvyFXmTL/9N2v3mLznABHG
uxtSksMK2Gh5KMR+IoQ9PjbERb0eWpzfox5WjA5Ntbo8jCFbWvin5/F+u61i9RZq
FGIOXqkcz24Fxie+5Vmqx58Td93aj69DZMzrYadNJ/3717on6MwZB+tgdJ/iE7kc
FlTML17eqYnV9vEw3+7XkclUgwR2BVkoa9Qfj3rufbxgZtfujBsG6u8tgh1P7Zmz
2kCTRsoaKwczjNzG7qWwXrrb34aYCGaHugdhMy17m57bSGiQzxscRBjkxUWl3IiY
dD7GlBwH8pEcN7DB+B8JPLPkMTIsuWgM8yTUZQe6WZNZ0mt+ZaefBn5Uh9Hm9MT5
YAr8069TwxHKRC2pcj3wq4KiZ3EVSuwk4zANNDupLe3WT3K3sUcGjztsr7v4fVEk
ADDJTi9FGATXNMNtBICk7NRxVe/T4dla67fGxdJQNU9ber0qNXC7vCFOQ8aSouHy
x0W4KBVz1wZMIVMJAzzRz8zDEAB5smZ6tUQ9QhPvLkvgOn4oca4iiQ86qrTgBdZa
tm5acHRTAein1iMDs9UbdqWIOX5EunVCO/PU1seFGIknjeNFzT2fQwb60LlrHZh5
qFn+kCDE6N7iFXiN4ML1Y8zhB55LUesHpHGhrPBJW0HqVIkGbNLxNfyfAp4B7M8Y
ICHJZR9CZ47Ql8nzgOGa8E/qnwngWHymogPwkOPq9yOaagNMFsbcKUwSODTelyDV
bABD1BSSHCIoyCx/igGnnc9jsoMN+vvBQVVSDBIxAPAgiqr+qZZKOxyLjmJhUlMJ
m1i1+lH0IBHeb4cMGlHY3NYXpMkHldGaTxpj1lAl1dTuRFHu1Tqu3ZvvwvEevG7Y
2EuapRPwyHauyu16qA4tGrRj64nke3s/Z7btv3gSwacmHJPdH6UnKTDdR3OO9lu8
Z0EseIbBnt00cDjoX0RY8pgRI9YOgpmi4hQRQtVutz/B9p2adBTX4zqOt84vmnCp
pmF1qIR/1tDOEOUBs+I0XxaqDwxenXihWnb5zqQtAxaOtGldu2/oxb7CN289eTBh
cPFMSy3L6HmO1V2Y/CaCqSS1i7uoMFjsHQbam6UdHCneZjCtjoyiyQ+YCFoGiJcv
tErzkUAW4VCPTSxnK4IrcQkdZfQZpURLghDJMa2buZFt/Xn1Lzf9uNeoEpj9Nbgu
6a+ZZspOJ2UGPXkws6NoZ09ZQ7wICLDZLU5X1IDHFwtXe+dd/UCaQawls2y//42r
wxJyeCmBo2ZnGEizJwnIbpttWRJ9MddP503LeCVkJJONfbAUCP0nbWgXj28zTJWN
bC8+qjeijkVLcq+inioCFeSLl0qOQbzUf/ut2hbjK3aXvsrUfmepK1J8I2m1c85A
uByrBx74j++XJ5IZpik7Vf5oTMzHMqoOZ4aJgvB70bEesCAmSy5S+cwT/2nSiGTQ
SQPLrgysbi3IERGCo3mXYqtkv4XoWIKwQy1T/3poX0/k1nzfSygqiou0C28I+abQ
+zW5vVB0ksf5p4Lvjk+KhNCRf9bj2sDm4BxluDj6dMbFlZBPnbfrTit0r/JngakB
k88gjAlDv/qCQ3pc29QhvkmcBs7XaghlWZh7aMTCPdPPWZj4UDFxmVN0bv3BDUNw
e3XKVP8qzYuwvZzlyy8nwAc8f5l00ang2ALEMzlHEmCPcBxphEnqj0Ja5f9Qc6o9
0TvRZq09c6eyDZebIFUGx7dno47HZstUBZtBUal67DBX1vdbVrfHnskiRZ1BespL
6TvPx+cLjxUvw+TKve7amjYDog4n6fi9Ky9g7r55qaK+GraNJjUhBOZjt/IjRdEn
r+gOLc/F2g/q8IK33MHfz83HL9cru5znWkqxjDqkZBtRl9WZHM5wUp6G3AWn1Rgv
G74vKDz2ZT46LZRKaqiQ0S2WaHzgyOrvTiRH2W0smGSDy774gSn+i4hiKJypVCIJ
fj0VyUBjPv0XxCgccUEZDJKptqUx5ZCePbkcvuDd5KT7AGsxvawxVnSSubvSoXEo
FSYcbUEEnyOOVmufwXm26pEwIunGR8gAImPwa47vTc68GftIp1TRZftWCcUq2598
3tIjwG+PlG1/HkjFlARH7XPr7ccA3ODBN5ThsCrTTbed5zEJvdcl2rOAT1WNaB0z
MAkszjNCSQ2xnUxBn7lU+T84agEufAP9O/LMSaAndhcCYDGXA4MJu49RTJMtuVcG
N3Ct7iVecIZyHpvPR0GIGf0yKISsNhSaLeXnq/iyRH8pp9efqhDWkM2FzWVHSvmj
JGFyFa2uNOAXax6xecvhEeiVoW/yeDUhghIY2WGg2z/9alTjIgymI3FKuOMAPKij
HaTm5MLU0SUL8PtipLvWnrC7hXnl3NSJuy5VhTVCbGBGZe7cTXvhQJi51GOC7au/
FEY8rSk48AQ8HzIrTdPTPfr/f1xeOCNdNyQgmwtS0J6MJFkg8BQsxyzIGxtGBCMu
yLOC0Lyukrc1X+sjAz/oO54kskER3bg6RWcF2h899CVxapA6qn/pSMh/PLDVUFvn
DYeJfIPWV1qALaUiKC+O+59dZDPkhMzyIrGONH+Tks7kSGBhe4V8W0bOCNmXQwRu
9Pap7cRVJ5jik8EUe3LN4WRwGBLzqGILflHLtB/7pk5oOiOcdXKfvgg0qm33oVPi
JXoufUV43rILd3ZgAdfcnbBAXYGMvw/aRKUWrJo+/xRbPQJf+2Y8M9vaPYEfzDjN
hkYhpLCTe7kqqVpKpOJXXe382A+gp1bkgPTWbSpnQ7XvR3nxVahm0VITdmsNPHhF
bCLNVjQpqAlUy5o+gg3hfQ2czInvF4Fj5C1DymCoHnaIDXnI1IZ8CYhONDrbMOz2
atay0f2YZdoTcg7+mEwZmeyAEKTuXrbmqS1/qunMOnpR3UIOwPCoDhMkjLqUfo3Q
//W41bW7V+LFc7xBPsI25AFrA8vSUonZAu0bVWLWJ0d2j2xpgoghMWZIfMz3Cudr
u+7wtKUvBOc0AO/qjUGCHQFMaQ2V6ePu0shj7BGConOoV/UXQshhREOPijVSARtw
lQKX1bNy2NynhB8xLGDIgGN6S0aC4ZvLpR0uCBqiaNCgX26R10Eo15LUKfriW2M9
sh6sBdQShBBG4Erukauod8+3VKx1YI+i+Qg5Lu/UxT88z8FpC6q7Cbl3Mozc0mil
CkoAclNWS28Zxjz07l8SjA76dwuKvF5xIfjvZT5x7FcBvadTaiJx31rEsh3o8i3D
WbUeLcyvsf3uwtZYbaT7p7WUAgp9Lf7f5s7jZBlQtMLH/XGryeawka3CksUJC/4f
PL5xyL+zfBThf5xZHr+Ku5ig332HjzoC+LqjVbCHNUZR+xPONLJtLjdRcXZ+S6UY
vGzv+NzN7rx0ioC30ZamAoOkj6Jz7Lm0/GxfmLFKzktS8UM6/jBZ0uDAI01JYEag
Wa5/0UBLJmIUTyBbFrSikFIoqdB2aBoA0lbv23aCjtHijL6qQgjokKGpOkGc9iFN
8h31hz/ixCLInCvRMSOGfNZL0gE7t8g3Xo2z/JaMhe5VSbT6qgE2QlOAyw9wrYYo
4AdRYJJCUyfo48x1c6zv3G5omsrGy3z6X6D5jLgOxL6h/xQ4k8LnkV+a2EUrUE1e
nyoQVxpu6hiG0YOCWPrG+z/5ez2+OysPS/d9tpW+l5CvR7PYJeNyYyrQ6S8qiFnY
gZ7ozRlHA86T5eGJV2jjuz4Z6L0xSFEa6MtIhd7jhfRdGu75RaTTON4V3rAmD2yW
7BVFgY6P1FhKMLNM0iEOYw1ykcWXkebN34xe2ynEHPbFi54rly/ABoZIJAjH0Vur
tX5Qn9hFoMl48aFRwsWXzIb/pOVJ9VZaLxXBko9n8UVBNQyPYnOZT0RkKYFI9TDU
f9jgoIE9hy57lYkAyAJNTGmD0EXy36al+at3YH+R0oAz33+tMXb5Bfo81KLtwWOc
f4mRYn0DVdzzKdhQuJgwKQCvUvZyR1uVumkzOLETcbU3rA4SUXz4ZwH9LwK29xkV
E6fOB1+7l4p0K9t++K1//0giu+V32tsEm8iaPox4OnCeNI4xr3ES96XNDbfz8f+/
BXarBdSzqzQLYcYRDDcW6T2Z4/5GGTM+3M9/p5xp+9RNeFZpt6HJ1e7vfhBazsf3
qGtvWLTNjMBDC2pk+BF/F0sHu8DPUW/bTJYFD+hGxWJwOY+ZpMn0VzNkAHwdQIsx
+mBVfFioprpTk/aVKoRzoqtiXqJ/Xea/mLZeoIxCXTN7P/2U+yVY/ZzEmWUXVZWy
dy8uZB/sEBgydlm5dmrem2HtTz28JLtlgdV/PftCDzlQDwf9/Imn+0y8Q1OGl5R6
h8umIOq1mslsJbt3sojjVPf6i02Ns43pqVFmdruY+G9k0xRorzarSX37vjbf1bcN
Ae5CS8a0q+W3gsryN+Q12vtIpyQtNe4bU/8R4za1ZGE1HLXx9qR2n5+Q5+y/ZPIM
XZ3HI78QDREjCmtWOMxDDc3urIknahGqbA+iAy1BHLdrAa58lbfLZGIJnbEhNwVw
PJndBWGfPIz74k0xJcITJlIEKaLLT4lQqRmNG0MVExY6MhR4Iw/0YRWLeapdhLcc
fehmRDBrEjtk6c7biLZ6Yo0FDWvws9IxBSpuF96X4BuPT8eWB3RJB/F6FAEu8Pgj
OSv6xPx8YCZpdfAIiGZ8ey2rKTWmEzNY/PdIo7SIHSEnoTYhlE0PBdf6uSWQpJIl
A+t8+GC4AKelcxmZUZU5Dm28U8BtVD/BYfeDY1RiZNZ2P7BBnFTNzfazFsDcxkfw
Kg7LwZT0iFMYHF7uvx5oYehhTFsMBD/pBvQip/VBPVUOJk1/yNIJmbOFYtmjwOA3
Y8l/Ul27npagM4hnENn+2s9y3JLUNgRiIL+ZQCwP9mWJKFiVUxVMk+BvwQykO8Zf
aHckCT2APptLaFMpcs9dYjtc4clO3VN+muUQtvHK+wkmEXjSpiDssg/a5YtdwpfD
/2dVhLI8sY61Ixdvy7wVSA1Y4w6wVp+lHHNsrA0FnynbqjCZdMCcSi8DLuosUco+
SmWrETvYiU6rReyjed2BsuM29/hvMhhiz9RgiIXHjGVFf+tT6ngP7Dg7KtqtFG/W
9W/UWhGMzHH6/wyl0NPSIe1k5MRjSFkxTVrjpILjZ3vnCNQV6+xVLODwM0BfdWpj
C5R/me97jsGozutnXQWBXFED6z+QVjHrtWlLl8wmDxLHkacaRnkw/SC4hr+SbPq4
p22/greaHntao6pBEMsRhgKx5Y7VzdV5q6RAUdcrfsXsIjYI/RPkMArmIox6a0PE
oDoNcQtxt9eWwRCLDZ4MrVCENhoP2+vGoY+F9JYG8FUMe+0LsKJvyozCHaiqZweJ
R4Ajl9ZKSS8AvPp8tZLzEPywv8A5qXtpb7Iddssb8l1UhEZPxWqDGrsnsIPVYZuW
+7zQnf/3wY1IdGjHY1gzvz0+e0UwHDf9UnweicQlL+XDXoZpEK0NwkzCBDJr81sY
JB4jPPo+2dhlbM8PxuDcjpKsU1k/8WWKp6VhirFJUGZyozDvYDeQnFcrnTVPREvF
JNVUwPrVLFhcmUqUfmnRGkbwTC85L25u5wVSevLX7YOLz2oygKeGsnMNkJLerehD
IALNv/lpOt5/Vd0EtY0hZDh6rC0pyO+bi1qUpmhnwOXr5stpgBMSbUn5t1GHoxiC
lqNHbKLGBj87xta7MC7a3JdyDNityzAQeohqzfg1h8MKexnzpuEu3o10p4Dafw6x
EBTryAq0oZH7J5P3+u9+3AOftzngUnuhdAN0SWIkdYQQhBWQD/MAOHds9MrAHIZj
9n/aea4lJtQiWxGAjpVgAS1YEwNI6/vVtwpE7EMqG/OpcwAxhTt6DL+bmuxQSbCi
jUJgAhVjGmQuvqjLvB9RR1+eVjekH3vy2lL03rzJuBaoB9WhWff4vscRqyNaeDjv
4BPL2dArSQiOBeMaKa7eFkNDmzRNbN1P/az0EYlw0OgR56ONGevHUKimENbsNiPe
Em36oVYoVVs0nwC+42FxuX8KKigkf6KIM4ifJ0/Xucvt/F0gczVnc/onUhhds6M6
SGVnMZgYnebD6zmrm9fK5IOetkFpe9jFJ6ap/y9rJaceWvZd/8+ha8TxtGY/6cqe
1KAVZzWAtLG10a/nzUOJP45cqxxXEAm8O+/SGVA6i6+BAX9ztNMOqmlguXStAq0i
b+CbZWpD1UXsuS9DsuCCv2OIJMNoUxXkU9hCoN11I+Rw2doUNefGati6TZuk4CJB
dN6ta2e6Jt7ggDuFq+vBNsZNz0czUj9X1s0/MPeEyhBOhDUxUayk097rXbhd+O9T
pKmQj6+HyUMj1RGbBcryqKCl6tMyAOOGDUOWT6a8EjO835VlAqNp3G1/10/POOIE
OzmHZFcaYexB6nPha5ESDcLnKG7AOy6CCDtm17yklrXYanKmtKtGafNtmChucIkM
uScWrg7pcR5pSZfBQ6IuY5pBVAIzUlxktkb/Pbvr+ULtMlK2QtBpz7mKiMhwndMa
3tQtYf8uw5ijYmXU8c55j3QyCFSUNt0NurwyfLNHm5HHBHv4EjsaSpoHbHI0p+z4
65znz2rzSYx89T7JgW+tt4r32cZxhytmtIb/jDrHnQ/qZ5of7uUxvterqnfBxSQG
cngxKGpqgV6C4NCSXt3yzUKQ50JG4M1f4ULdnaHxZtYFZdP2A+LUaXg51o+8uIU5
ZiqisLkcaRKDlMXz0DWRp5+GUhdyGsLp4MKyQB3LMCcAVK4yAOo5/rCgrHe3hVlT
A1/OuYBDiYU8x2w7IQU2K+WFNIaYez+stjV8eLa6Scphlq8wIbfGt3miRi+W1aOU
CdtbVfEiQuQMYxjo/psVbFHHjEBdR+A+Kj2MiQ6VEtA4nJg1ctR/f6JOcSKqiAME
tlm/H6GmmUXwEOa0A2X+go6UJQgm6R3EyoEH28GruSY45IrkV6HcZfx9Ar59nTOx
AqQ7QRCjG8N7i4tWcCXty+XrNv5PIIuCCUKoa2T68JUjPUygHg3H+ymMgZtqNcT9
exgFAk4n+lbxSVDzf2QFKwfWKeyJBcslGodt59EimD/5205vybcmjDqgN46IpkQ9
yHKpmFKWb64E+PUImRFFtCPJjWrnXbsIL7pmX5DCPgSj6iWi0MIeplkMTrq9J4Wz
ywOgX+42IZub/OWNfyCNyWhjKLVhsyeoBLGGTirRLX6IDJDatnAQXZ56T3369EJT
ZkOcoj4OLZusx0+SuoPp9JhnkFu7Z2teOMVL9l2SH5HOLDdWgS8HZnAXatiE1I+r
1rBOr0NF3ont29zpJ54Bv4GEp9P+AAKrHN5KlQphHQ4CwwSoPh8RhPUiSzV6/DmX
C4g1xQjF0ShBdgryNxZrDzZz5ZSyXFwVuuY8WMaBhSA5lqizL6jzGD5Rlp1V2tHZ
PZ77sJM6oAQNEvUJ3L0JXIkDUfjyal2UiotxsLN0w9Ml7/eYMF3S446MIMdpBCOx
wUvKtPkq/fqIxL0L4scSyvCCQJlhu5gLo2WaTvAvElUJg6thKSgaLTerjPm3iRpc
FXJRs5KqzAR8k0OFHn0x/1nn7NOjXzqvctTx8C1AY5csbtRCwKxtPr/6ku8TEfLt
/zsQ8r3hq8XdATRB9VT/mSoUCWNZhoHPpAZaiSL/DmxCl5XzLpslH+Z/PajM6t6t
Hp/Ryt9x2bb3KP1HRwU3pcpCnligMI4882RrmliOvmZJ15z1fkcxtP+tzo9e2yWo
oPBbrtoPdQwkyPxvkGOMSZQJ/7nEsm/PtkZvhzcCdTXxsLsRcWqdn9F9ZG57jrfB
OXJBaFQdkgFk+s8FRm+TsX6byKXcIVu9cZt3a3B70K/P4vBfX5TYL+RsBSmE/2ID
TIdpJIWpKOFMpsbb2ugzdcpzjuN2OvvvMLNcSns0CP9oxdJNSJPo7KRj6FKVMlus
H0nPtUGMWvzkToXT9FFYdbgmGrXdY82pHsv+bQv0RVn6cM+61vCnF3lJf7KG6K83
eSwBgah1N299mniGA5dTkog94Ue9D3vhVzXEeHu7ZJcUo8UJO1zbScPI/lZeomXD
LDjFmY9kPFfdwadkPRzGarrT9tyOey8sDnR0m31M9+WIRdc/ozimUTd6vWKoOEOr
DVErogj2Zd8cjJ5qDyeeBdACbqfa7fgTT0GcEA0csdm0tFpFrYOalHqlc+Emm+2r
Ozvi7oIubyD4kD4kxEK5/eZ166dv58VspSUZdUA4nb05Cs/v97ZbusMeKhPyk1j7
0PvQf+fvr7JktEF/B+EHBaj7bcOgQ5Y15BO9vhn4XjiphLEOIckSb4t/o6Bfbw3e
eOvqTEYe5hyZ4+IoHSFVTaDoR+jfRGh6pCYlfMsWfltfhFmlHKy9qpgF5F+voaOl
W19rGRNeDxLv9Iov/KHWNbULYT8zBIzekhiAcVighGQ8ThBeNR+tF5Nu+R6AjKUc
cyXJTDVI6FKKh+fURvOgvb+OL3OcLlkFzQGoNXyd0sJfAsjhrac3mGRQYLCBkd1v
fP76nlr09nMOkQMcSuhL1vLyS8tHxaGf9gtxqq7oYbK0u6WekFYRud8h0hZLPJBX
w5ERnfrEJDyVWYcuDr3b5l38PWWME3/lQjeu4YpiHY8PVbm/Njbw3FXxIfPOzA9e
UttmU0xuIKZ25ZOHni087W41TT7lvs56Bw29JG3Xv/dQi0G21aCZBcccihyj4v7P
OEZkdlILKp2STWLF4te5Rxfdrn0PKr4dPuRzW8GqdGrCBV7KvijWU5QFDAhtJraE
MiCTICUgqjenj5retvkKtVkFcgnrkV96x5iGnYZSZYHbx6BBb7/M2JkbqZ08Nkee
K7csebc3iTfNO5P2WINDuLfEYGMqhbjX8vKpoxifz+s7bK8txnnh+3k121nDdqQK
jSbFZeGqAPvAWp6LmpgFVpTmOKqVuy4gLtHbKAhZ1ey3sY5Se4IQlTdZOMKff5XT
jrYbd2BGbpKUujnLEUoTF4Yl1roH25MsarC6mb3igdFSDw2eoTHjv2pxVhy6amch
J0ywFODIQTZf367LOmsiF7xuYuOpyzF7FdNYiLeUmUC9mfEScT2v+bIlmHhp2Q3Q
Fh5oHF8RgnqThMGkm+Ysp4lOX9ymuHMbCs8vdCr6TXNAB4nRrp+2oDL9PuHN7wCm
ckGz1qGATOcXRV3pe1ycvxRGITYdyN2aQf5h3JJhjJqZy41511sOm8IdjeWP9jaT
v+nEE91Sux/+wVKuNY9Ex86hM0afGo20QlIfDrk0Mv5mtBj1cDh7373bTLSM6RnR
doMsWJvk6Ag4o0/GWQ7kcqNvTwe7zrO1YB/7y8vHjzvM6UsvR0206CUnZRs0dxQU
0uyQlJT6PhbKwvMUOsLl0P8kZFMjE62ti379pjS/TfHCAezjsW+6xFF5TDQUxZ1c
/miAaKMoJgloSBpfe/xs0+L1x00kdnFycKeZfTGKRmrA4UEHuxidPKW9JD+bKTdx
BTGjyw7aNbRMcIdU8I4azrv+TEYNgTVItIHqb0t4PzguTldtGdW+i/gV7Esp7zwq
fz7jiMrdGsYiNICPeF/YkCj1juPNNqhFcugA+Jx8Fswmi/LG3njveWJFQZy1yq3M
hjMxk4NH9X4g3d7rvFGn1I0S9dU+wdd6+0G4Ygv3vl13LvhYrrPwu03uwGK5fBvp
Log9H74uRbyWJ0oYDotnmrhbIsyW8A5FyBfDVUsNalr49v0otPqtyTWTRIUJcbg1
O/MxfPU33QUa5z5tkrSVtYoA0ASNDTODxRyAOBtcGSBFUqSEU/aeRajMJ1XiF/0g
/ZaUmHsEXcGZma8RSqT+JvbRYpCF2r490SxhMw/OKaduchQsVPrkfSRRp1VKRUUU
m0F/QQQKQKY8oKUAa9yZ7Qzkev4qtKGPu0Rgs7Ao7r4z/AvtpJuUty19tDms+zDu
0V035mtKitvcLBeXpaTopkF1p8dX2dXc9qDNW1Mvh7SaaGAUEZXhBoC923sl6ZNA
LRfYcEpBFQAM7G7vY/ZSs9oaAdvsWyMKhRBZEv0itX/X4bO7ynI17CSUIZKHMrWG
yxJZk8Ia/4wo2PSFAEACF8Uu0TnFVFXvtxu2AlGjy87o+y206gglz/pg9TJEN4Vi
ZXexvVRvrX4I6Ar+vXC7brCNis8I6EUdCzOAD8rR2YPdh3B1ii9ZBqic763m9SjN
5ziqLahSPAxOmkrq5vMQhg7dSC8DDIS3IKGk4oR3BahAQ2IUlCeQK5TwDPiktvIZ
hbv+5aSB5H6YHCwqvZe3+zQzuIyACAjrLKKh4Y5laZ0hWFWUAVFMlFS/91bbNSgL
VsnwsW8MzYKDGGOMtF6sdOc3ZlxPvkrMCpQwebf5r6evspgxnEszhcFWVxhFpVjS
nXMuRHtZG7gmG2ShrmMXXAYdO5hhluHoeqlcjoMCPXQv8Gs178bHstGTsix8da0z
5lEYA8oCC9+ps5RxyJXf+zFgtqpiEIJfBT2xOb0AonaBD1FljwUzTJyRLnmn1PWo
Xtfm2kuZciEjEY2RBFoHTlJyBvjLZqpLV7cPhc8/72Qfn/sfE+aSBx0r5SXFl6ON
vhD/VF68h6cMnjtGfatayt/TlfURpHFg1oLfURqTIveVM/x4yM/KK7muuIwYVu+g
Ge8A/VPoR8dU6/TowQlpqAgJdmHd0/8qYwlApjdtm2q/MutWKUUP0ZeU9ew7FR44
AkshdHpfc+Mpw8d7X5in64TmDubklb42BCHUHRI9eg4uHnnCHzYEwE/gfhC168NV
hRjh/rhW9GK44zrmQpzkVkBRY1v0XCMB4nQ/ADlvOaeAb/FF2mBZpwodU6tz6y/S
aHSiwm0gpgseq5ZSOYWYowmHBF2qzYDZAK4SjsSWgsD15VeTOHVWBpBg/+McKUjO
xJ5fkKNfYlDKA6ZgCHslCP/CjAnTTdOblIoiz37n6QXZxNB/yuPjkEvpimoRl5vD
vbmTPm6PtlQFmBulV1Fb/frNWEdkeh7M82ImIjbBd8kCWOCUUuM0V/i/fXx6GPoh
bFMsjee43K4AXFI7yPyB1tF5oJUkPdjtgfeSFh8U44xBeZsFQ5IYmAz6uq08ek7x
JnxA7vkAuc3py+Taree6wHUuyVQxRCW880d7ocSi/+w9uBprK0q7Casi2gv7NGsU
urZpuSzVb+apdYadWJiqmefKtYsiBO+EEkv1TySbfFwxV3IjVhvOrAhFVskgu3eR
bj14vicKxQMj589eWSd2XeXa3tsssaL+d7d7wJvNWYUtPOOnQZ/8yNxk/xMp9sC0
bvZzik1hix7CPPe4cmzAuTIFSt1Z4G68lfXv71jAtFRGfo0XrMRCAxncbtO0Vkpo
O9xGcFK+dzVQ0qAvn3Ztd2MGv2TLfVFdA7CUiNkPP6c6m2ql9xBDXM9KipE3Lf2T
N2rDc1JMw3kiOqj5Al1Q/pVDBhShZc7HxwBzl+aUmVmQAQRBp2N7FNv1pp0oackG
Bk922QY+R5Dy/YJty2NyOI54q7Qrdo9HvJsz0QYiZwwhnY41/bT2w443KqN6LsUw
tWDRE2G8bWq83pXrhBU47YjxQ8BGDs7rD67CQ2rWvsuX4byGBL0BlhyxFsNra8+6
kfhfaEpmQyZPT+EekNo2Ak9KMQnRfTSJlNSHGab+TopUthS2h7jW3GHRJ1A/BYrO
ECLRFxTbV0bDhkfe7/7284hqyOStjPRyW2ANp/0YAkT3lGS2IFvvbztSs1tj6idX
yN/8L0KKIbaK1D/RooB6/eEoFXiZ1AZ28ALZdSbWxwSpxTRPoR90cxehdPhxbjtm
oxSLYlvyknFJZNSl/3SagPe/V80P+AUlunWpgaP3be0dXRWEx4wFqRJ3FpeMSygJ
uHjKy3DSMsIq93NjTLlbuilSFAVdINiVpzAGeKdpJ0EIWKOxxQd2TpOb1c6lZ7Bi
GvXFAzW3cDRqLTVh3u9fHyhcL7Hy/h/OA3OPkr16iRUdjY/xSalNu2kMNwF69y4X
9D/P0fs8hXlGUw38Okzr6EtgfCj36MYVjKBg3D/JHxI0zcd5doIA1IiRvnDgrG5j
t6o80nXO+y6pOr/vyygLwhOn1KGpZB4qJP+WyzkOLnrvMxjQB35RbCbsKJv8Lq9a
tp70znAgS7Hcl/QxW2tGoUSOjlJggKh6y1C2vvQvYa6zZfdlL2tlcsPI22Dcq5dW
INQPX35XsXKtis9sTDJ8v82Gvpv4rwhQXp5VqFJwAFHW/hE+/3UuAX2G6f+m22K9
9l3P7inBwL/1LwY3ANPDSkKwbEO39WOOHyqIxe62lsrdV2Ue/q5CcvpEDdSEWdBV
KGchfk/LKoPfIx1Y1LjwsCaysbyX69y6TLvt/CRiMOgPZtDaWv5MrJ6rdSRzRqu4
bYc40Ra3F21uYH1DgcZblUv5enDCWclyxjlJwNsK9jndXLt171g9/btTjpoSgZ8E
sl438xwLLDY4SzlPgRBW3dQmwuR5PNNf8eV6X94XzwxWlaUD4FGQdZ05vBWTcBRJ
HPnOyPcvwMq7+mE8vzs/7wUcNCr9qOvscHslyqqtn6vYavCBYgo43JVqeX8pbou/
WXX755bsM4fpcvLZwU3OCF0MaTvlnf3MxlunDfyl4TfeXocJ2W2wH76F2Tb9NIsY
OXRHcCW1frmQ3PqtWRMDfhnvYhcJCqcQw7yMFNlpVhdAbiGKGsrR1mwHc3BfihpO
G6GnoJaO9d+sIPnvPhA8FHF8p6IvvHJGMvnY8gYJfwrSNloUDCMqONXgi8GimBmm
gJjkOvpNEt2USVs3h+2LSjoe3c91zGyWs4fSnEQguwM7UcF26Kep4YUeegFKqWXU
gpvj3txoiIknw+vcdnCKKy5sLGafnGNQIkksFhRac+xjy6Nkx83Bx2fPPQXO9iYL
jKpFXzrpSZW+bnZJXvpayThRzJppHalvh1jYQB5C6ShMc6gkvhpJhlvQpXhLzuZs
YStxDLt4LC3kuZRLrHdt1dh4+gCKAWuJNLfo8ORlk2TsBYEc7GyP9WBwfCpY22Vi
jes18dKLHZnYXUH25v+ouq1Cy0dKshWP1MwmAhotw7RuBXjksq2SmJ4nSa+YQxP9
9bEaWrPo/kKakig4CvvLSkWey4ucFyR8Sy2IyliW0l+VUI7tYrucWgVUeF6MvBw7
hfFM9mOSBiQ/IV2a1xXBKIRCXdmXfM/B5jGno6jk3pgQ/YxXwdR2hEVOmQhequcR
M16JC96lpkcPGiBrbXwQ/KW1xbzEQ5/hIwEvMcmWppro9T1rvX31Od8opn4UV/8X
h2CYFj2dDe5M7PKPs6e5FN19ZzXUBzvRxeqc0SZ5eSqaCtLvbnTpMn+z8mPxRmtt
V71dAEuD1CycE9LQFJqQhJD4Bnew4wPBxw7hNOsAo4p1f9KCt77YbwOnSWhJ2+op
4vbmf7h93zGAWgMoOkFYl4OM7VJRU+HUsi6o5BkRR1wZ4gbmr5d6o99i8QjFCXsD
Ihy9I4/t+6umnM/bLeEHCWUxvinLXB31H0i1y3SnSYSpb5Zm5kxHzpdYvfmEco7K
TyOjS4Vx74limqMcIGc5dNx5kkkaly5xWwlxg86Ae6NmB/5YzyhjeP0NadeLa2r0
2pK43Vq3RKJH3qt1aGIndAIvm0Cc9m+2FAV+YJ6xxj8lBkSCnF1VMv+1jIHyxrrg
1sytozIPkqT2/leuOWiYngRa/jH1v1qT4gPWwxqLgzla5FsRv6NBfVcP+1atYln5
UpUGt5kiejIAlb2eboM3MNS2d9PFNqpi9s+YKQDPzQOvRqKki37P/2a2UfpNxeAv
UHGMesr6Z3R4C72Hswz0GVziHOwr5c0+455u6isSAiDh4Cjl6jGZAvJ4mm5E2zBg
zwRhmxKTuVDyqXFeVND9CkQNhISG/GJuSgxdTWyn92Ww9YG5HagarGk56AbpBZXF
jK0W8OmDB0ybG9SfXj7LmkeO08eFx/6bb56FhSvUNNErTTORMLVKLlq4EhiJWGgX
iE7dWDYk5jzMCKEpkTGhsVUJRDeOp2lngMNfKuC8yvVCt1mtLTymkN1Cykr07T7Q
Okyn/mJiGRud6qoIs7ZJndSI9GcqxGqIHXlNqAvicWCnThmAvOhjpzjyyneoOVxD
trTaSbctmGc896kFuSz++S1wQMH0SG9x8eBGPA6x/IlMzeFDoX9k0vd9zhJN1W8C
P/fi6Muf0WWv/IJaresBI3905x9I4aVMth2f6I2k2XdpXAEMDinjZXaIbDzuzH3k
slNZepr5XjVsmkPD8Lrlkn34Ygo5zevTGom6xzYNQNokZR92uUyu7VTf5Zc6lhW/
UI6bP4H1ZHp6d7X/du4Tuav5iGYIcWsGj2/IF3v1OdgU+T+rhpZUcqbl32EMzY17
h0MqKnva6huYZBnHPF5lUQokf/aV5NIcCWgVRCkp6jL7v+aif/8rg4mPEC79bEl+
QnX9q9387J2RV7oTg+7oPJsz9sMn22PAILBAxpi4VBzN97o/dKHrNn5INFY/WEAf
0ZFniglS04XJIdwWsL9s88lHgZimu2Edpi80X8q/csqGJ5WtxOUNOA9i3si7kal1
HpvorUxhmCvfuC7lNQpyL9E+1C7dAw8z2IHYdxpNNrqn1wtMQAPjEglwH7S4tlbN
aOoqBv4M/PDA7psRovKMPN7I+5IY42dUXIs9f3M+Rb26LfORhqZAEBIlVG0kTrfl
JeQ9/lZKXFk6Y8/VXy/I17BRFzNXIhrrfSHv9pftW4EGLIIpORQwJjqBJ7Wxox4b
QuE7IxC932nyuWPc78PM5yMVE7X9i5+s2RKeqTPGkTYUmHQx0ABsxJO1tHO20Wb2
HxjTNqEDvCiCx0dj38MLOHto+2/jMoN3MdzQE2yU6VcdgoKvqdQLWZX+jYobcV5Q
pBo5NU1VLOkQQJmLZbIvl9Zp/cOPLv4LKie9fcP0z0afhEwpSp2rA/W2vnw7w0uJ
fKlJxmm5z++mI7E4xjDowG/eFcH6cJDzXa4ydwChvrrpaywTCKMwFbvCcXB7b3+S
NJpj4D7/YUEhzL5Jb1krCLyJXxwc5OeXxcGxZ8jNZ3VnMe6QXtQYTlSPu3ZGOvee
t9BOnwcDOiHb2HicHsfnmT0SL7zUBJ7eKbo+KyIdxyzDB50gAnUZZyNNlzpDmyfe
MlTJPtHzxl9uTXvCJiKWajVe8079iq35HIAoYtXqpDp1kowSr+6cBvCmHxyMWCf+
RkCuZFdT4YxcDa167V3vY+91esZoak6MGRQe1TwOFpyyUyhmaqVPTTJ1i3KYAluK
3LBhiMNS23C1S+SrZBIy3uyBJSM65W+EII9pz0ossQptRAXLuEpHN8NdvsQqGTld
HYk2eb7uIlpStfJMzzUQK7xt27u1ktlhJLroBrdVqYbDhCKVMOJYlE8VLyUzGnjW
cgTbWCTWLRsTj/asc7oOCMtc1McJymYEl8+r9+nEsrwQLgW4EtrheVPt6GbXbPQJ
CFF9tRVcYpjFNjqzP1SU2ztzBVs02vLGsipVrz2LZcsp/YcXMNA/Z8y9XJRlMP3B
q+UGu81BOCqIpM07pQ8vmuQMlEe2Ug9hBNBNtbpk+OHB04xxGI/EoZP7lrRWUb9x
6OdOvUTP5vPgFAkieM8VI8emm8ve51pbPpPuRNnrmOdJ2yfoJ/sNY6Ki5gMvPZp1
ns/nsM49vHNM8QIFXJim905UwSYRzDcrZadTQXVmO+qdrCvhvQ7yQKUZKTk0yDYp
Pcq+MJrrjtvg8/Ne978Xe7L5tbNAzbq9/XlOh/PXeEhHjOl+HQX3sdmcRRF7jP9w
lUmmwe9vARAfLF5oVuzEgrZ7/KC8MLNwLhbDPFIKHmFNulz0K9ksQQgWtoAXFZpO
aLvUuxyY0kxNJsR+5oBtm3ZpTQ0k9AddT45ZJLBQoD8sh4pleM61bF+xRQz27YkA
iWiVEVABLk8TZeGqiRoDtWOEkyB9Z3/W3oO2GDQ2ApZ0Mef+TH5ORzYirJkCgAgC
rXxcNq4PRsPu8bn4Lk1wDSXSxZYnlq4U7OO5nIbKvbQ0eA0eBP5z4gOBBTIUevLI
j8iDtFvRAroZkY7HSWC7z8ymeJnVsiKRBmyp3i/GtoaBdZFDF2fW7wEsBWs0ekiw
knCOo3Vn19BU4153VKmGy2Yrv5VQlfBIzt6jkqor7LADIPeyOLwpvH+0WCYtTCOu
UUsmNvFyPkfPp61pijrmk0JrPMoUk4EMsa5AH6JfrnOIhb2VMGyD8Ps0ZU/GtnOU
FGyzEeIl2wdQ0PycwL0qo8ujym//l1a7xoUH9vyqaLTimqJLc/ha1hS2kqT71VwN
3TSY0ryOhZ1psXRPW2rISFZWwer8gCB4ODTyOtTgyMK4oA55T/Z2jmGvUCqBU9cE
o/l1eYrzSM9dFl4q5CI5UKC7g1pQOkCUexCuPUBS0CBxgI92eO1Lry6VNBiXMi7e
cxSinNV/8158Hs2DAE87bbB+6PQzj4GHZh19+KxE4DoVdg2xKGkrHxh2WFfc+0gJ
dXRtygLqiwTAqPwupXq+wUn7TB2XPDZ5pDjVNBZeDeKmmr1DBYfiwassZnCoOX5Y
93ZzqTSj9iWjbDkGVAX80Tn99bkEX7eLrVCD7c04ouKAaZhQgEFt1+idawGnGRE/
PLu1XsWxL/jOCw+kNhIGG+w7GyYhC03h4TotZzTt4kHXMYydYmhCp6lyaSqh+XxV
pEJceaPJ13GxqB4LjIbUeGZDTxpSBbFlR+8kpY5gBhV16lesmRdhudMIZcGja654
OmgN4/8SDyOTMS09GQ5d7UDvJ+BEseeXpDS/06mVNR1Dvr3hH2Lxo260PaiXw1qj
vBykzxa4+C5Nh334w24LtxB3AZuPDXzdp8XYzglxjGi0ZxCZKjXGTwQF0m69/dmW
6uky9FG4i2hYBtllwydpaR7t4JBUL/kvTO6vD6QB/pIMV5VuN4ReIQ0mBvulvOMQ
4eL6xU2SBBku/n4HKR2h/18icS0Bc0XSIHnovWnd9WR8Qowrg8Dv0rl5uAns0E/x
20ckylXsbK2BGGO9BLGZxyUivI/jaFtJLIywIRl0Bqs43BY0DPC6tZqauikYek1z
E/WoJfLojXVOP5KWhoKeNcgqO5UJXQUkAbtzmRUtMffcJEOzO0kYkr/dexUUoyIe
C6AleEDWR6JI09tU0HlBuO1Gu7A+tI3khca80sE7da/VFgHx+I1AdbHYO3j0wHN3
aDuGMghC4Z29AfBeiLP2iwuj2ll/X7YkJ843kiNTqcFandtX42YKEAdu9uj1/dkj
RGmCesivpc5s9Zt/HzvbqaBFyvaP+KcoVJB9Og61jSFGzmAr04xn798Mthm9QP9b
XJHWaC8FhHBLDGCgc+T5lusTAJl61evWyuEcrFN52O2Ey2FezQBGbsaDXT3uSXFX
A6oGlYuhWc2mGK73TTNpgK6B2+Xh6B++TqGqPJZnaSZWi4z4pTk6e8H5g9y6ehhH
rRImBq2jXwpdH7Nlh/UurFmnSvgXzKyAtRB925U6EnMCAti2bAnA6OdBqt3vGniP
Clown2pkODa6La4EhDWsdMDPg7CxztNP8BUleGOLcQr/nzEFD3N3JTaTE0+8z7k0
O5Pq0JRYV3d+rW71Cy2ldJ3n1WHGlRbsn/r80LCLrkQGtUxvgNMP8fmNm194M4cK
xic7kpruYmk5JqhS+zYRXs0uoBqat96Hp6U5QkQBaLI9ZCM0PSHYuufs6fXPEmPv
5D0m5jIDg5JUQNIhrMPrrDOen9r2J/yOMccJvpByWIyxTpz8+WhmlWqEm+6W2afu
xzx5cXqHXaJ9kQbhWb6jq18uRvWPgWIaxqsW1LL6bIRt66+GGWws3orJk1AKF8ey
0/MoFepy1s7SfX5+k3Jff/U1hsd5APCnkX+7vKKtT1ngCu3SrOAEuVeWMo7WME2S
zHWMwtLr6T9JwM+tzSNm+VxluXDLFrNImQQAgXLV2/f1BPd7GoTumkF4nzMgdhO/
oeLB6Xg+WHIf/vJSxcjM+z/viZmnBSMJDJ8cr9IHk7S8dI123MV7eJnuEtxtAG5i
JPnuu6U1iXaEWFoFGkYCTE1AD/BSqlGIJxFlW1ceiC8sL6FdIARFwxghlrmUgGTL
fwiS2VBcB8utkeAcg2rYiGLG7qh4jELn8Mn/Kk0h5RJCaq7L5XOw/1EMsdm+v0pJ
WlmFGC9pqUSagt2C45mkJ+PQnFZZaYsOWNZGjDKV20rq0IyKuq2qr+2MGdWGONFL
Vk8UM7Vbcc5UxuMsq/Ogg+yz/vHpikthvETh1oN1EwhSxnMdvwdij9WEsA5smHze
c+I9B48bIIkr68/XJrhiVXIemg2jiSKREddhHbQTjjDG3V1mqWcu1Ful1sYUQ1k0
i7SqcX5Ea70Ey9aHW/WmtbTIZzaK1GQjQ+YCj9Pnk8MvDW6h4rNRRnQSocUFEvDH
QBx8dlkXH9K7xaPiB60ebc8pQ/0nNR2/GBkR4yAbV8j5wbL+PZ69ELhsj5acPTXK
uLgAhw9a3q2kw6Dyas8cCEUynEMYVwRp/7kpCcxQ+PJtDF8JLFaoN53vLaWWf+Mm
pZWbEHZGT193xPJ9CvP8xo+ybH8n6GxDSv0qTZ5JJZdPgqJdTWMQDORUvlkjooEL
sy5DAMPLRsZHe5I/pV3qo8NtzLGsl6eTwhJpoxAI//X6ZJFBiFOiUxeuKrGZemf+
tT/onjOafqfZUJxlSEnCJEO1DwuN0GwFEI0kW65LGU+hZDgGh5i4OCrTZplhMrEw
Luqj6E64tx4w4iwW+CwdU1MlZmXURWUqtJ8+BwJwuEg4wql3EO5/rTrRi/dLxGpj
cJHeRvejjZGNUgGNUHwdyggl2WhggTKYmBSHWdSjs4GXMJkko9wtEEeRKuwx/nGQ
CI2/HkGZVA+xEvsrfEd9+ArowWZc+NQggChcbSsu3cBXr8WRd0H4bYRClwGnjwyC
5HmoZdloUKQdIOhTUdZoyJoxSOERCfQwNT+28kocnDSrgoPIbuf3FI5Osd2NtZ08
i2GnkmhRbzfZJLZHe9w0t8Z8PZrpWTbthOxJ5L8tf4ipwzVZK3VmQ04ca0x3d0pq
p2pBqM1YInIgxuSfc4weZ8pn4jOOc5apA8cLj+hRvfCpOEeOGfhF1chdsBmPwTAi
5gL6s+Wx1tbxcElwRpHqN1QmbLTdyPdZc+55+aF0/MUL9/Cudu+hUBS40wfTuTeF
VR1Vy22tXKgRgb7RlgzteRJYis/vLbQOdCigAFUrZZu0T4ZLXcDSEcYktLXbMFVJ
vl5hzZzlkQOHpZRpcG7vreWy3dElVnuPNKArMwW2stM7Fr4sQfMzVxEmogNjS9rM
NrxRcjj9TPfNAKtPoGa3k6rZ0IvdzPKhhyavAyJCAlRWaPPS7mV1XrrKzQ1e60oi
Skk4nw1Ck/w8aTjsB28hf1H9Wxcd6CvhqreiXQchiGlJVH4NY+bVE+wzBUJKiHzk
OZW3k9h7RxTXLZYhLMmirax5TO0G/klyD/2q69aso4gCI/v2Z/Vy9dIYNx/d7jbb
cpZEaqPxWmhIQzHtbI01L2UiVJy9ABVPsTwdnBXtjbSu/R/uWCD6ACxg2BvH9bxV
kAwZeHYcQ94LvDG4Pol/iUd76vy5fEl0CeKHrquPIyIGVFZ4zUI4aPrYITIGF79c
HC6UO36jHtgZpXzzZUGCCdVHixAQf0TXsf+5Si0A3DBn6cs96ImznxkdLXRdFsMh
vK6dg0IeKmYPj7Sb+z/TxK3BcRMeldguy9qvNQjxd0RmqySRpkAiD56ReaG0VWy5
KvMzR8NdfGhUNWLtQcDnGMGBFU8i67A6VIdpHys0Vv5yU9h/XdDIqYUMFV/2Tq1c
91osV8jaGZ6ZdS4o73riQPHZLRacOLPMCNmG5p8JXJUDZ/SDkes1CX7rYHlU7Iv7
j1aMXMA+Fy7lXCfiJl/67fN9f5XVGxQSgM71Y0LKSuJqvmzhiX+t01oUdoxoHxT6
BoHiiCTI1lRoGnpbokvR+WzO3X+1XFtqo8cd4WAgk4X3lsu1w5/8UgeY7cq9wxxO
gVvXsY/p/o8IAX7I72bL5yP56JFdzE1i0S+eV6NMgRHFE6nZs2XeeHE17QOFpHn0
YRPGtvjCmf5TzFjuJLiKcpvWKdpdwh1PBgbpnIZtqkr3sy56jjPR+EvFBe3cnM2Z
O8u06axRfGruDkxSnS9bHd7Ewd9OxheWRq2SvtrI/ASJvgW63fDmMV4t8wEZfu40
8n3dM1iWYj6jFz0w9FOu2xCP0QOEZsRvGIa0EVngYQLXZjvx9ZW+ldeyh2jZ6LRk
8llxkQoDVEiaBvydASY/zhDgXEdqN1B6EPV3fYfY8IgPxoKGrwl7y69I3p+FunHZ
ONLmjWFEnW2ACvqKXJE+Ux/HwWtFMGlrHrrkym54QA/ln17zj3v+HZybbtvXDY0P
FJbyFsktAM7PBENmqAnl5md/RMhFswfxtdW6WP3yQjA82qP8hOkhSR5AY1xgkX1v
GbrVznIws7QPh8t/kfg3NvEDcSAMI7F9Rno+qs4Y+aSmeJuRFvFcFgmLx+sd9vbz
MErbRaLQA7BwsFbmasUewkRXE+0RvyXgBnGWpbSDsF65QDjmtkmC4Mw3NawOvEiM
V63BgEsuJzyDu1wqQMAwmMMpq8w6allNoRlFqNneeVK5pIQKY/dbDgVgFIj4gcw/
r53p8QCRQRWOTzAeB/Ji866qFZl/DTItMwSo1sCFF1Nsa9fuFlbJQGHm+G0WcCfV
5+HRFDPK/brHqr6vf7xle8rwJlE4IZPY9vx8qIOT8Vo425PoZDiJj3LbEEhBUXPV
qcnKmige44v0iZnGDmTtxHOvErs3WvqRcdPu4KrI22xv4Q7A4WGxnXrZ4yWCPJZ+
xH/NPEbXP4+2Fwfbg0KI3LwJ8uhWKJnXwxOyJ6pRG3Jm6alxmlxSP53SpyZFYGvd
K7eT/aPtu97lvhf04UQfNJWFRassL19sNDFjMYVUHewb2wX77std9XjQKwMXvdkE
bkd2tF5Lry5zsXBUWqYTmh05U6zy+Cnq6yLPvx1yBBp2GzSk0t58DLxk/wSDpvEn
mxAWjTKoJGtDknbsM0/MZb9SEL8fqOV6+AGtL/u7iH9VZ4JlBg7kahLJ7eCII/NI
x+PU00v0d/hBbUqIATmx9aq2JoBCEOvK5QmBZeLNtRn+Hrna3ysGaMmoWhl/jbO3
O0m1s2ew97k3LtgkWUD3O1bOL1Mto4zz0sch5eDlfPRMdlpR5m+VoCIQj/dd7280
9NVNbQeKXdJ8WIVFqP11ra9lm+G7As9Jtg+7SkI2joAJuZOE+HTKhPSPPXvMsTBG
lLeJuUG8L28l/XiLaBneaPRvMFkIlpRZz6rrhImqV26wtecjA1ae/KFKLAyPLAn9
d3Z8CY3cTsZmx2XNHwriwTIEJC4Gm7iHM9PefbNJEGwqxnT5XnZE+oXnxeFK3tEU
M8a0PY24W5lsHs5lwrD2WVlD03bEVMdPnJWaFb7ek4C0zLz+rb+vUTM3c8TSPkcO
46v+Ly4AV+HM+0W/2dasytWNo0KpZpJDtlMcKwoecRhhMbw0yDwg7IrdjjOfgQfU
tNai2sCTVbIF8rbGxNhCrstBeE9dHaceE3aildncc/UmfESZ7QPjmaMhzwbS1eib
FDDhsSJFq7pSJcerNXnvGvK60lsuSPIseaUWU4lNRcMVvB71kgB5IuJcHSVNTOV+
OQ9fjLvErQhO8iRkG+p7V4O2irnSuaRWGow+GjuNNglepalSU3v1b/38jXIbFPBC
35TXkkcaJjfGEbHGKCaf42TuYO5j9xqIh13avdCj9hLaA6UYft88O/D2bcPu5K+v
FC8B6Tob4KNX42gmySn4X2NfqsyfpqG1sJdv+OprIv3oC4x+pkeCwxv8itH+RsHN
fJDeE5bVeqWiEHTNgjUqt7bDpdptjeq0WX4HeuN5NYYgzCF0Nttdbhb24E9zC/zH
zIcprBYpamYa0vo4f7DWtiy43354pwvlHRKkzrxrEJ9IbT5/TRD0Bje6pNR14gVF
3R74ouFHnfBcGw82YARXCBNxsRJhqbZ8ubTz5/AmuXBPNfgYH9zSX7LUrrnXnzgU
Z6yZ7KNQBbXCaO90QV72RQG7xG4HsBRlP/RRhqGbMENvU1u79JEuX73xDGBv8nOc
qNFI+51d+ewgKK7q0sGlXvjmd3TjsdMl+SmfDVH/Pqof79JOils3frlJOIGjCTuY
gJXezE7cslz+twBCordSOBP+/KgoUaB76Ar8zQxf1lNBDctDXqvEqhwj0YiGnLHD
2YUWeFFulrowcVRYXEASsmbvZUpDnWP8IEt50s2ITHu+c4Sce9IWRs31vwWQ6HFj
draYvqn5cNdwxa7v1z+ip13UBE+/BwuRrrhAmhyr45rIcc6O096o5CnWU6P6ApqI
fD+DZ+udxh9isJwJN0HZ+hvEXJEX0gVqgoXQx1uSc7rxwXDzSSFp2isCYV84UYc4
2/zN7ROQ3n3MtQtMikknrbnfzeuI5euv8S9+tKpjfhYV2j6tJVQEZuW0CZ38xpql
yRop6UU4QBOwMsofYnYvQli+blCs/d3X+7ggazh1miE/o3bRALV0JzAcraVnNLF/
86MvJhTLKkN7xYv25q0s7QdRz9EC/54NaNEFWer3K9TLNpN3xDPimd80rc37yqQY
uqsb7xTfjhh6vTvBaH5jVOJaFu4Dq0FUsoyqk3a2e139tguR1gW7KawjBBm+bSLc
vCEWeV5LQdl1zq1CzuWx71kMwGOPKNSM4iBhAuc/3TLhO/MqufmEy+0FkK06UcEP
K+vuYeRw/kewy8xod2ZtY4SNtLbSI+ExdyOCgVdokEFovCieE8R45sM27+POa//B
pGT8FdNtfQlp8Hmhxezfmx0Z7OWDNOPJRc0mydfEEGYReMZojEho28jKUDS9IOJY
2hLlVgU1+Gjwd7Fqime8Mxudtm5eAGqJHIB0VMQczdL0+LVn9TbFCGSb/e9h4Rwa
pHEJ1KKpz6CWJsM9Bdm1rWDHI2UC+ncBYUWJh/0vA8R+Y6ONvkFeIHYzllpPvHr5
s8ay+jUKW0H9iJTs5woyNmm+d0LzLJb8DMAh+HIvc7rBWxgFn72yW1pS780a/d2k
7DU+jTw/FsqVKLW1emRj29RaGAUoYXx+ZTtHrQVzJT7wpo0YWgGVp8kWoAQOY4CH
J8LSa/dHhoiuWdxaArXG/i6tFGdUkfN5X4Rk5fYfvtGAh1reQsyugnFtouq6hPXQ
3/gtik/2OMw378n5Ds4kSNFz/24JqdnGuUhZlVFlev89x+sUa98fhpT/01HntnFk
pWU5qN3mWOBiqPvJ361CHS+RunleAyNSqUm0ioyxC/qQFUBucQQdA8m+aaZDhpKn
4cA6gPB1YkQbkuTulXLMqmGkL83sZ5HDy8Oc+4KZ/IjL7eXZRAbqVbO1SonOOA6H
m7zRBrGIiBPPnJ/f2g6HoRtr5ewslOe3TQ3iXy4wOooPvOhK4KUyClyOg5Dhu7WZ
I90EVOaEYLzxu/GTJHRT91CIUOmSRcwWK/a0vZpf37ATshF0VgnaXMIYzVG5yOcg
iSxyI2Vb9uievBhqZzcGMtJSRW7og2FKrXyNjkZFqAXWtWyG2aFN+d30hPpQeQwG
uV1PwsfK5fRR7Q0vMuWVwktfD5NZ67bCsGxKNmpAFLeRofuMrVI6nTUjuzWpOaD4
4FNZFFVFGJaAtzMmh2tFo2t1i4DWItq3upGVn3Cb5hVtvd+RJ8XDJoiDyfxJ2A6a
kO/Yz4wS5oGt3eoFcR0dxwYG18Jiiv9F8PTJIQB8n+spoeq2riNeaPkG/Tn5IZpm
mPh2fy760XdXyyOn8/wuUJN7MJKEnz1X09WIPAse5MXZQQOp02+4wmV6cldQiUAu
W8rGfsOQH0Y7p3IeY7lJFvxozeY44kYFWoMzEkhcr4n7pHTfPaZ9xUrHqFQLdWtC
1DwrqM//zPxnPYJl+inbBk7ixpeWbwSFlVN0+SFdp54FfYjN18m6qAPAKmCA7awy
MH/j3pXpB+4ZTUWUOfTDpuuWH3s9YCPDUiLX6p9Ie/yczBV1O8TLu5lkeF1+ZP5t
Qt42LulszPbG4Lw1UoLS2fowvYW9vm4YLWv9UhU2oMfkns92NC/r4Vk+ngCVUIoj
fSX4ckM5sovZZwV0Pxrrnyax23YUrA6JJfTLzBOoyGpT/Qs0Lk1sd2cxGfWbCk42
9mrVG1QdYG5GfDrrU6TBMFUDBUbZBPlduDHeCf+w/LRfLU2wGoUlj27EA73tAB4j
Sn6CqnY1sX0mKeL9MMcIMccKY7nqUAKg7unwNdEAozoRL0W2lBu0V94pvhXL0wY1
XbFAxcendzRvrx16Qd8Jk1TMTvW/vc7k7DPds74dATz3H6XfO2+jN0i2oalfd/bU
vBBCS65i+TjBQIuUL3WPuZO9kuwCdqN5+er7PtFpa8m7zKHE9je/R0dl/Huwq+SQ
XGEg9e0tPMmJvXxAmFHRsrWNaMDsur/008pfMVd4NYWnaLbO0GiIsTGB3orBSw0D
ZFr/fI4LQSM0ObhW/1P1IddRwSqkSdYKBQc8ISNHKXEcNWeAS9ntxY38MYsruy1B
2ISyuo7/AT9Bn3QCCRDv0E1oI8G59x3CIvMDTAqbkXD4nN1uZE+gPtGA6CG5zfyU
logVNbSCQpMieoAJMbhdDBtii4tx530jM7qA6pdSL6Hv7Kjwn2G6bVufFDpLCBBp
gYOUx5Yfa0kYJ1nAfawWJzjxYgSrMlHe/oaejPBpRxnpUw/CpbSNAGtgEb81DQQ2
pPTcE3sv3dGkhqMqP1Otor568mhE/DxFMGFI4mkOxPF1sXirI5OpFpbD/IHsx5kM
JgDtjp6FDP4D3ZBaCqI7K370UHCXdbiHZ7xe2IgQ/YYf0w1YZXOLt0KwqoncMrH1
SV0P3UZPiLcxnvtl3LxgJdNGpwCkN6NBeIyElXQPBOFJrwBF/ER0uHaXMm+TpL+v
llTuWYnEl3oDlsCOvWjUSRMwRanNe1X+CgmztwF1CKubdOnLuFlk1f7DSHDpuBE1
5qQBWBT4KKBXzT/1LIinxTVuVXu6QuTQPaz3anEMxbIJ+SfedgQ/AxCO4V9GhxLb
cmvRinC4mwTrna9YPCa81siGeMvTCV3tk3ToXfP5tghQ7pxNaOtFi+XbCog0NTFP
Jdkt5coWpIsJiOs76Xp6WhK7uzZRD11CSxujQmUeVKWCoSzTkfFlfH4h7OGKOd7D
thQuHz47QLVAlF0dbSyuA9ic5N1DiRl5gp8xN3oGjWfJ8ywqYskA6NwIjlg1o6ec
5+zCw3E2APOX9VjPfPAFGabHhmffTTCsmT6AcZv5+4Xscf5aI1jirgueaygXLBMP
Ha7FUkoWVVmW7CSYp/Fu2YDSctg41rq5SXbx2Gu9htK+cVa1h+7Km5bJ+WVCSt1k
wcGKV8TC/I45T64YEHThOEHulZBw9zxQoFi6OrpHClEddLPQ61oG9gRMMYNKLldF
mOCfU6IDdPTrBpaCRvs0VV9pP0ifKm7cf+FVNBFQqhsSsD86wRSW25xug6rlxpEM
MNhXHFBJqHYEShbmy2Lseqb10WQUut2TnMpQnDdpEBZMFLauh7pFIlJZKH2H6W88
4Ki80AIVrzzBH0K3MTd5+pRSOSJhmd4vBwDneEYdMje+tPNJL+1wBJ6uRz+D8s8A
cv/EZIglAjcVmsDx/k4NJTrNaofVYrP9wyra2fjtEDP8DyfjS4TwjdtNB5LN26EO
ZzuyftsJfCpF9i6ZAhV156i3DNr8Q98Bt67lXhuHVb1jR6ebmNpTnoWfmHEx6mJ6
Gvsl4usIqycw387CBFrGwV+6OnD2z6bFzxiRXMPSp566J39TvcBficlxB0LYrtCx
Wp/lrJd8eUJoli/eTXNVu5xHhbF4r23aVIK/t1qO0KMsHP4mNuL3unsn1bNO/yso
rksCyqiBFXam2tpG/NUts6YHd9UeHkKU6fEKh09/auq4F+WM0+QYeZWFF+WcgIiR
98kIA/uELEoHm06IOM2Nn1//T+VgA8AbHJRjamQNsVtQwtgckxWliTG50oI3Nj/m
RwdmtUtTt6CxVi3v8PDXNPWuZXF4GqtsrkRkoGJZDCF6bkhNFvuZKB+NALBaSPZZ
y+1ATqdRdncKHo+hCJ/2E+ikD8slM6UZxuiIpWwxKcQ0pQhKFY4hLebZxw1OfKGU
lqOQ9viARFJiPMRyp0h2QKxzddK22kmMXpKj/L+Eh4/LrWb4yBa2F+AlJ/TGDCZJ
NWpkTD0W/6VpAl0vP9hNuvgXEeO/L1TjylsgICZVEsNWvJVGN+UvRR2eqGVnr0NQ
K3KJOogn8g8rtudCN5dlvARVS3mcHifhVSM6kvGvysG6EYo9bo4fy6Y6Q+j1miSy
oO1zfSLoza1y8+sX6HlLYQl5hBWqML8Rmmq6Hh3ZqsXk0ri87ZjtVCdF8EHZl4p/
TXLDQOSqOoXXCGRu18gcYH9hTgkDvUMs2/UOK1EaEfShvhjNKrZZHc6VGReriuYW
iaA/HoP5bxpx0yOqwlwZHEqKuhUuRM3w4qJJZ8AQzqhJbYJb105szki2fcSzdx4+
/ydr1y34N/oUEAIsQpRiKnfDuLoFf+88FQpVM5EH5fkc8VwYWmBLfm+hi1kDPxO7
GZrE0W+SkxojrusfiJ/du235UVzFHwx16v3adrGWBstOm4+buz8JSrBcQlkl3vqB
2rALzHsKWkDWXw94NPZPhsyrGyktiNoHnwOvqg7cSRLJ0QoS5LqPuZUKZ5CRbVBA
q/q5jFRspl3v4woWH+6G0swU8RoxfhJhytfCeOuFV2it7j1XUaJ+4cLceAE5sJIg
tQT695kPk3KKSpD5okmArzg2mAb+8rdzweqIM1ayR81BZiRsBMrzb1cTd7rX62b1
AxcDx++2ie8co0ia2Bkk+B7nuVMWI2eo0t7J/jZJ2vti7ecevVFP1diPiYX7Ix24
XSzcwkgzGCZ3PnvUcMV6cHqgnnrea0Tkvehc0pIJOnqziWk5zL7ZgLPyXrSil8Wn
a/7diZ0vxwO1j3hKEu8UVc4tmQSpbCe9YFNk3BojfBL20UWRgA+RT9Caodfo9ksn
2oda6a5NrDDcMEiE/tIo2fRKx+A3YsK118CVBfkFoPn2Rj6DvjgtJdMnvZ1S+tyx
T4nloFMoFgkDeESVAmhMkxlTh5DipAS3V0+d2yc2QPKZYnJLXpjby/IwA0XD1NbE
QNqqBNQab1jGdDXP0sukB/g8hQjTl02DVF9f+77RQuFGu4EMZFZtAMw22zaSwoPt
o1PVt0AE9OTG1tgNhuY+4VN84JXmZkIzr5EQb+6P5HfRFm3iRFMnK9DdnPYk/5HK
yUamSw37r34imcsOH25kxa3ni91Dvys1IuZCJ7CwamLI4OlW8m6/ufCNM+i4CfLB
P0DTK/06+sUTDtzeL3moix6JMBq6NKAjOy/xWoa12rmVVirERstIqUgaqiB6cyf8
osILJ2y0NO0IKeODUGNgL4MjrxNtSBgYQYQpewCvSnba74lxwfaoVdEK8KDOYtsL
qBgOyai2vJ/wSM1uWKD/9B5MVR/CWqXOWegSDZW4Pl78GksZoNnAibyTXS5u/Kbe
FAIOUtC6nffvfXvQ9Qb/8P9RfYH+yzIa76VEUyxfuC0n6WVZAvR0jAoBApOaS53z
wzPy44Z15l6Br6faIHyyPnMkFUyAysIi/4u+1TgbahFQA/HC3IQxrU36UW/FTx6L
lSp+Yp06kdX51A1WgfERGe/ZXGPak/uPLGDUSBNWLoLPB1ZsQ47pAM5PAux7r24o
Ij56c56wO7WkCh+PFWxdTONeO8UvQ5bNIjP9wKZ1Po3ui+8ZKrXoW6OV35oN88PC
bFC61xTfAFpBcZbxMHvBQit5DmqoJiUwPYri+H12vEEev8vcMVqZcX9bpQSlbstq
xCTE90nZrnaSMCk3qToUiJNj0Rt1EQIOkuxLTC5uT1Pc2QUqfGwFadOnuXloOTbG
ize4A4DIS35+C0x94+kWw0taHyC4szwyzI8h0vodpgcg5XuxxvYHqJq+mCUxQnuX
a1Z0NNy+LeA+n2q7/bWy0ZNA/HJnolqRimHt2E5tG3teyf0weAQ2BhpWIMLkpF4K
MEjjxg/4Gju7M4hBXJzChjoiTlEazJanwCXqgT5CNDbKfU3oCOY1TJ0j8kyQrUW1
M/hJxC5CzGQc8ih+gw4UfUtPIMGv3EBVjfx/KSWJbibefT6Mq8IGYNIg7T3aeWhh
1xJ8APovP0kA1Q0Qa1A6uPKInZUlI7XyacVYlT/4a/EtR06rZIZwlPX6Xs5uc6Wj
ayt+c1hppcF2ai5ncbd9WQMPxf9gqsCSDU33n0RJ6xNZrCbSBtOu7+kgmjLiUF9K
+0TVyi3yh6jB3747F9B+hgNsRpjSp3m9Vpo2cTf32z/2BH+fN/B2gXQcuIeTqX+7
RdXEc6XttQEvDyApOnJ9eaKmlFQhM/wRSAZkMfFKFlaCy4JyPYUOrb+czEI9BGCl
hfn2GMuS7Fi1wEQevjbeLgIl6T5HvI7yPufPQGzBVGvpMeZ0N+QpISpRmgln4hu5
JBsPwtTkBWV1zY9WQghH0DtIr0j8VGoa86basVBC/iJza7YoqqA4Ux1JpY74/G0+
5Lyj2gDJOPTYRFK0XHp/eEVuvH525MDMt525oDt1Gdhm9TrqQDKejMz+vhsjGmZF
TC4PDBAHn/23LxVEWZKGskruUcNybF8dikj12xwUuGMJIAhkZr/H/yT7GNJQls9z
lJGkPd5SeA8Yz8G4qwk3AGftnq+sXhaulhdnjjhKvOHB9vvRfYJ5WMLwsRCHxrGb
rxYAy4qSdQT0ycRIcjppxTYnWqorsP7rqAr96nGPgi31PfqDhO2dXwA8Pgy7OeKJ
KNxyNQHTjEdFIFSSkiIm+rUA1HBSS/v8P9LZiS0rCdOoEVqdBZCjrXPTx9NJ2f4e
iPgx86Vw6iIhNZuznW4ECjkj7kiYwYBgtB1fUjQUzq1mop/iCqYuaDM6JpHCJipy
Eje0/zmFY9v7fzPfKAyQdV/5DR2YT+Dgxu9GCTaNjXNjYcD6MbxcjhnBiZBkRT6L
f6ZCHYXBRRwF8b9qKyyYEUgAhOjPs53QHazdlAeKjsbr+RrkERdqerA6nvg0o/r2
gT/DD0k9FmR6LnJ9nd7SavRR7ePnmsQH9M5CiGzb7tJQtjPKgcEbimFhsWSd0MNh
ewuKlFUAXPW7NvHySCLVbpUkIAEdW7+cd0T/nyxWcIllmJKvEN9g1HMTYTD589MQ
fyR2Np/yKb9faiJGxgFidbW4sh6nOYRmVH6xK7srG6n5OIx9sEE7mreMrGSyeNWU
bJdZygWWB6GWlGPIhghUrNAhAeJnJiFSzPyOXtir+W3f4Z3Ohyrn8jRZKi9Vh01C
6+BHWpVc5REThoJmJnIapsxWB+YGyjO2VpMyUGkYaaj0UQW+/QPguTg5a1uvc1W7
LET7LzSesMYcvaDoPpURaSJGjjzIhjfUmPNzSUDCWEytlN5OclVJeoCrDK+CY2ck
MbJY5PjFyYEDp8h+AKxavkZDvqSBgWA7yzf5L+A0+YBbU/ZF6bg/tC+9809+I2t9
SPikp5drpWRGJ2W3oiuy7hF/hqG9J8wkjfcb/aNWt2nl2R6GNMmRFeseHaVad5Rr
P51rZdIUlE2l6Gn7+oT1M37twnauTCQwRsjCP9JkaijL8XMGtrgasZ24QThbMHqL
Od8SQaRlS+qyqsGnQ05cT5E+Kaszbem8F3J1KAeMNlIVNacoiQOEgNz7v3aWpGWm
Nnzcfs9dMDllCfME8/U/ADkjYwM17LuSNLLw2ZgScwbB17Dnw/sJROzDH/SxTLdt
R/YOemT+T96hu19hVitOaUdGJrYIoZ03LJNqJJYHlotXtcM9JqjesjKSZtRltOR1
M1i7IBoWbhiKLmivMQ+igcZ/QLD0Oo/etGrLlspBCr+qizkRj6J3K/F1VrH9Bi7e
Dbdj8sp92w0r9kN8AFYUVJPBQD42EeCFXvDvDdJ7VMD/kioVaKJZDKoS9kjVa+em
j8wiv8HTsMpqqUb1tlBM0s4xVC2vS4Lpht2DvU58T7i/IjCW6U2LnyUKc6pqUgch
vxiASxB819z5bRd09iQ+HfttENlHXrzruU794YkK/+1yUqo8c2UQ59J+uCQ6V0KA
Yz8IV0VNGDcS49eehoUoPlWlGpBATTFz610we2gSEKfTTg2Mtiab4tqfHH7pRZl9
mctywEv3NAn9ziN6WROwqpgS6uG/E8GXs7V4vAEFFEXuqCpfYbM1GXpCN1ynjyn+
ORKTRvTb1Ne1b1ZuGJYeTy+pTIyGleOSOp2euUzV/hGQkttiLFkrlh9YqkbdJpEP
RlLrp1GPm2oqLya+qCcqnr0FCJ+od6UGEH0KSqIVvhBlKpYr5gD33kywqV7PmWxZ
A2BR/JB20CjufMDIg1b52meCWLtzofuafKusBi3eFkNFT3s731exO0rKO2mMAoUb
etlnL8vlgPbK7XGsaXCF+2VnRwRe0LlELvm8AC4pLdIOF1TxhedH5N+SWRbBILuB
bWE2wzPniXwbW5lI5wb+DST1obB7TRNWYG37l0ubfxbQ+pa/sgjGXNFIUjE8V9e0
0ey7bKJXxWmRHaVlhlAhcvWA+fzacawweDBhG/ZPFjwj5YKuBYN4BdN4UcJI0Wa3
Z7FWUsWBONRMNDFJiGoIYWc9dDgbsnO/iHWwGdc3GpH+otQ0WHCYkBC8ltcj4Qz2
RFRHD2HVbVzixeK8G7+toGmEaC40YUyCTgwYD1JZKElDnnDXT4g/UH8fl2wDfZIG
wCFiaZEKZXo+wrMNbKz2SXKttCHgwKxVv156TedB2/oI5V69hWQBMoKpSFV3Zw+Z
hhdVBOK60QKij6cxrx05zxJYmIyM7CGMlDbmRpksOap5IVR27EmHJ/jqgquQWAwd
fpGMjvkSf3AKX0j+5OPw6OYpqY3x1/SdJaM9X1xwjx0BIA4B8tPcvUXwmq+ePz0W
NwxHQhMPmjCi9riRhjLstFtiZyg3WsLkBvg/Duw3OQVXInTv3gQBpfZHMnWtjGqE
ZXBCZkvaUrOU334wibjCZ1QdlHKVVOk7HU/857CrVgqDdDEuIMFrizLwSoPGRqrX
ZgWUcQRhkjpuSdrn4/L/90GvE2k6LskdPlQFPnxyKx0Jly5lv2ZuCOPJwel0xRyn
pHP5GA3yA7y+9xl8Uf8zXyI8yrJzCrPjGoeFcN/H7vXKzo41jtXl/irYA33U/Cqn
1LK6J2PYhHHR+lfbUJgmljO7Wt5AI1o4BuiAp/zFbSnkBzfTMlALkSZ35T5F1+/6
WXadkum55uvLWxzIcLrendUJ3LLrOKhKObT2Paasm235gjLaZBEphFb/WAD7u/+c
ihWcAbuu/jkeUKO21hOT/m0XeonI2NmT/CqLHqSAM2wzGZ3mPRaEZjLR+el3eYBP
c/5RiTAaJWvXiUYkT4BE5Ox5LFgfyHRtxO0hceu9gENKaZA59ksGw3NqkePI2bY/
zn7LFLl4LDCIRbttvLF9EIZgycDmWsArqNkvAxSp8/XRuxBon6vwRv9+8wtyMsuQ
sst4T0f0d1E4fdp0V/k+7eN65Xd1CChOggvLAwBdTgx5a2SYL6clTazesFbakLC6
8SnNZOBbI8XWTTCPJrG8lGAqGB6EH9b3Pt04nNbrFVq9DJIR391KxDmfKGhAbKqj
BGznJnifgPqltvhei0PiVz/yK9XkVIAOaavbn6HHOxlaTV6twRsDtD6Mpm0AXtuN
L/xzOd0d8nmzKLzk4wPEFLBS/Iq2bKZucTf+HN6wCnwJZKSTzF33S2lW6uWEs88b
P6LRmmzStX6u6FyFQtX5eKiYw9+rqhnzK7ARb5g5E+45WA+BFvw10r17jDoUbOSw
HvMUFXBYWiDDK81XwiLR8qsOxpdnr1+ICeTceKcc5Lt/2G6LHmz0kOx2nf+JDM3a
pMvHeDHBjNhYpJgNl/T0pB84RNRYiWmmvcEBGftAgGgOD3qtXt49/LBHPKGljM8T
16CqDdzbGU0neoifru8V+Uz3LZ8tUsjd22vIV1SSMtq37ok4pGjntdSsHZ2zJ8M0
ePA9hbYfQmGvBMYzoLicTdguUJ7QglEz6bSTwmD6N62OzCDHLMxba2zfgz5Fzc5X
OQgo2LQRgYvL43j0aywvaPVboABFM03qDQ5NFcdywjQRg3Uoe7JrKt9vUJOV2Zny
N2h0YvY9Oj9zE0wE9qrGnzQan36AXtl+fdJh2y7uE8yF72CjCSa7Fm4fzBYEPu92
HjeSNjgdGQR7J2vJPUO//PKbMcC3O0fBQwhrErXuvSMLVnV3trIgCGRNtAWVtl8k
DL22UO2jgnAeANduYpCPD9UUZefdd4mkc6T1KzQsTMyVNsh87mPJSm5+a5/TvNuS
5JrivlhxujIlSjCanWJvO7mZvODhvjXZkydOMGovsd9PnFDi4q9nyAulUs7erO5F
nRAbuyZ1tDeuwPy9wJpWVhjAqLyZT4OcVTcRpDGfy00NX9oj+n1snve9mClSgwJi
NDE6lilJoXC2B5RaSdTviKRpEaqQRjuhBJcHusaszcVLikoYb8cndb80NcCO7AOr
tCNdIB3QEvr/bI9J5FlcYRZdQENY33eIiUEjP0ZGlRMWBVoWPL6Ha9EsolSBv5YE
/YGow8PRmQvxPI9dDmSxuh435QG2tvx62V19A8xZ5R3KnkBmFiY+PdtW6NZet/Ol
GcZEUDuEdjhuq2MMkuvhlJGxvPbsL0AK853uoA7jeL2unU37ZwdlvukzznRpxU7q
cxb9iWYxfVpJ8/drH00LbP3N+qQHj5m137cedqydoTISPs4PXiWMj85+7/SH1HuD
sYiOhtSh9qRFLGaFEXzy+83B8OZtYKgOP9J381e7cZy1XvNdQiph6RQH+faWoT0v
MGUqtaX7GW7KpSbUge9qby7U1S/v44U5qZsNFx4riSSu9hDZJ19G5zYRMYFat7R9
zXyv1jOD9kuGnd2t4PQIEhWS02LiKJcUG+FkA9wy0sr0piOsi4CY4XL8rrhttYtl
6ZP4LYFXEGSqGGByomCHr7x1d9qHWUBE1giLHq3fUiWKViSG7y9DkpMr8fAOP0FY
KiAFYr5vh4HvEMnk7d6TcKQSbih0NVbsOQWxhClkHHvWX61o++OJPeWhXhX4fBDB
NJGnqy065eIPLAa7AIsunMcqRIMJsAYp1Ypd7pJ0JTpR51ZLdW0wMdadjcFcc6mY
mghK3qMm8XiOv9+VLZbVQ721qjdJtM3ZAnX6W3j2K/QVInddsZaUc0vFcutp+eka
NsbmGnU+d9sjNfzXN8PCmMefzGxpUljA5Oi9mNK7gW+hCyJ5490leMhtEevKT9rk
QrrnbyisvfLNyFtgb2lUDxy2JFV1th2GGKcym5LzWI5E5l4mn3qOw151cYfpsMS1
CLV+1byM/DC1By/VTiFRWKtzq+tXHq/356BHhE3otGtXtwxmRPnLr2oi6rA4p9sZ
GoMyl9lFxom/0pN5jZS5RRcezy9+XUneXbGjQ/FoZTQYyHRr13durJc9a59zHdQf
bKD+YQswvy4pT9QLFSoTHAP2lFfYqEgpVJFN2piV/vdqUzXrGx9KakQEp8HbGMhh
JO21VpYhZN1M7DTQkgSYbDjXBD90HC48SDRvex5DcMDVdkScejohBdhsaRbGLB0o
rYpC4LTjTAWA3dcY5dIO8txxfp/MA4GDOrXNWbNBhXL/vk5g0kUgVHbkgB5AvE+S
p1W/fLtc+5ttKjEMCAGN5/hRAFq0JZgW1GVXv1paM8OmcUPQnU25Yx2VJgvDj7x7
nVJA1rPd6iw7yRuhQzYACSxyJRKLOsmNbx1f9QKi8DqzJFkDRUzHcNpWsi8Vzdmb
VYQpduaUv6BksK/hJyKVEu5wiOcv9padtK7RAj9Txg9lu3hcmkHei7OoUac5EqkQ
hL+N7sTNrFWjvF+mRdgbCl5nDXy9zhkFBy0xzc49ixlWMM6vqTRPUfE6rd98q4xg
tfKSe3GQYQNrIO1cVKbh0Cn+4E6zForl+vSrkrwH5xh9rhsBHrlDz9bdT7tBCDSj
HxLsl/6YYRY8igUiuEcrK1tPgIFcOSM88xZH4ePqwwg1AZYZFMaCvejgejez4zYV
6ofrkD02nI5CUmSLrORMUiW2Eq6qZgNPHhJ6ryTzxlc8uuQSJSWUk2kmkN+WKevM
fhY4kra/fKiZWZ0YAVj/9jh5dcfFqDmV1uFNWU18c/ONJXoupcDaUZT7VB+FLhl5
T8voM6VB7dnROv7VRACuO3/U5jJnyE8UovYiflKKZcNon4BrGKGq7sPBy8x0p+VK
GeSU2twwqbJIk/uHAAuN/1YT4DrqMYzOlYrP7gCS0+CCB3//Hte7zv5HBDk3RzaR
mLFS9O3MDhvlBlDqhAvmlgWpsrnD0MbcGa1KJ0VZsSqKNdjF7YvV3te5jRFXQyil
5XRdnsK6fE9imjpgWVgZqUhRDRZGyyaaiBCKd8W73Ab1ncpBCPvrJDHFRkJJH89e
fBTVr9SoSvsd/VRocV13d0WcnVEWr8FHR2F9LHNgvYMNbVShaWVScFH4j/zJltUt
0+Y4bV4Ju1iiGHEmqkQF6yqO4KeCWjf40YvQC40gyjhVMEXWaS84e0NpW7PIEGb9
saTRtC6DdUwvxm9RzuHZjGrRDhf9tPYBUnenq+QLPJ1ZZijBp3jscl4S9w+8VskK
ennsE5hkdJcKsk7ToOf7/d95hUFsyWqFjaTVLH9K4z5ITT91BOoUpoYrcSH3cek2
AGXsHsIeU+Oa52j5aGlhSTkFIKGqNc0BbzFunqmhCnqSrr0mXcFNB8quZyo0wAWh
M3QxmJkmZn6qlvnbYb2y/WwAAZwnX0fsAEh9u6dw7Ug7GsU8n89MOwU56M3ul0rr
pUH7HtJFUlI9JF0GAIrMXAdkum4o4Wsd+CITzrZjTu9YbgvGrQmLSZbAMCX//xrV
A6EXJVCxZ+EDZ/jgwPPUg4/b9Tz5321DVSPcXkUhM3K70cgOY8EqmBlJ6guldKPj
X/cnLOJ3+28x/HiPFOmQPtlYhMZuJUKEvtI/WjCityWqGnRczzomG7RCO7xNel1W
vOjdeGOgeU3G9MXA5/QGLYFzLy97l5OAe4uU8QyEtNUmHC0Cw4XanbWjpkV5j9x+
OjY1SpGy1JGG3uZQtOr4uLLs76iyPo2tgTOrEdijrCOHCkvYgZLMlygwSHfpUNKB
odi2kI143Ge8KKR/VgTrUsgvIPm6QUpoSkuZjmpD6nOzBbLZYgCS+gk8so3YBzt0
JQyKIuaSIxniQvtSCfya2tqeMhvOzD3tbOERT1pqh1bWTdOSw3afechCGPdC7AOe
aqgqkxxkG78CM9WvDG+EFsIZUnGVlfHc9AhLQjxiS6RGsajiHTkFP7a1UdCeH+6N
9e5S/gO0yoSc3zTNr377ITjqshYifhsJoauaHW1nRX7kRl1pybR4XPqv21Q0GQfU
Oel5XG+OecG67E/PzuChZt1h4UQajBqYx0Z7/Uz16xmyeU2jWRSYDBcv0eMq+eP+
57i4FlVhBZXCFF3Q0a9KCpNVoiSjqNnxPsvILVGtq/w3URhUpGPucL52ZmcuS+nM
E1lz0O6Gt6N4ibBBOhcdAB6a0nbhhs7cBlmcY6VUpsDvD54VNvjH6hrLm2sFD8w5
NAjq4Jk6XMfkhbprodyw0Cp4AxmNm0CsUjWo/EgsAsqQPzm6YAHziAI/rXjC2KwQ
hL5528UzZkXfJSj8hyNqli430HWE8ua68uhf0c2Uch4nCeZoWe554zkuVtkESSrR
p9deXwPd9VND+d0QHi2mjilJE9jif6Fbjpz9U3iy3NXz42GHczSvqf9GLHgMHEIV
EVsFI3nfQwO/an71K3VR6jt7UdhPq7c71XgD/wwtVszZn0+5y/jA7IMRznJL2VtN
/wjpyMOndmnoHm0N84wWPlWrU4ZPG+5EI8rgWDfrFkTpQ57LStSdND6N/dzjGuqq
3EenFO6auZdkwBdlm5nendj8Mj07jA6vJC1PQ68EDwwWJGKZWTpD+s1ZdZz+RbCw
rxDTmd5vStCzwArwoWQmFHz+/qMxU7uo0cKTsYkrrIr7IBAqGQFMDso67T8OPqN5
mdaWlrXx9btegV5td1HeqmwP++AMSTGPvIRFoaxOBuWkqsIRrtLUYbsqitkZXVax
9nUt1HG8y7E4MlyzLcF7Xy8ytkuGfqHgFCQvW+buPxc6kO81fhGEZFxjikzuR5gs
veGdDG44Nt/1vgKEVP3Ne7VEMZXj31Qb8W6UFceIBv3A+veS69K9WzxjaD1+QJIJ
2WOkrtKWoAilZdJGqnzZUqP1tigRJH/rUZSFSJueCZzc3HTTcLi2rmHVspZVzodE
Kb1ABF9tE9goPid0+hlONXeCukH/GUDZtGnjd0W0EiUjRceJaLbNpbegDHWsUwPD
QzWNWmqPhWjFo0xmN0XCHhS4ekYJyO2AFtQwdmYx6HNO4we62VTz2ZChosoKsvgn
X8tCHAjYrWOtbAHljERwoi+FtiqQA/decpSH2x4qhAO1l3+L/qfjxgJvoqAZsVsK
V1+L3kUmj46trlB5/v+GMFtrluf6qRsNE5t3qCKLuhCGxQ/B1+bT6bKXJsiQKxd7
vETgt/ULpOw5MR2yeegrwIByy1ehxBVsdRi/9pgfZ1O7yaHQL+2FKMntRjnuemG6
HWyauKq3im6Ic/4DG/DylbNG4FtFtjGe76zWYSRxH2oKUvm39KY2ZwKcD7RqchDc
5iAdW45SlFIE5ZDJ1EOvXBbRAllmV1r6fCe9mL58sfOeJDlMFi6tM89igGwWLye9
4N83pN2i3y43CFZ2jrw+8D0669ttF9exfPVWHk6og0CS5qBw8EmFIZ2RHgKDrtMt
1BkvDZmE64emB49/t1UcWe8GN1yDDKpbhgy1AUCE7NfBJi+H78jTD7wXklS9x87R
uOEjqbEfDFTStPPm5lhKWdpO7cjGHXwIX8bUq1PC+022BwEcj8tvKF38O3pIVnwk
Xr2xqxMq1UNTHgLVgZ91/8vp7HIhHYCIXIQkequ52W+hnA79dzQJb90UbWk0rYvJ
83gO/wOThU43QzFRhszONENRD+Va33jUANKeaWnyYewpSr/a6zjky1fdf/ICBOYL
zkpT5x53Jpq7Ax3pj0x45QyADpecfcxlToNSonjSx1smpT1p3YAfJ2uPXWqOjmGo
rXamDd9tTWYazfu78JIUVS1dWgJXEdBbtTV5LPPxLBkSvzq1vTTf+VKQ6Iahl8Qb
3Rcmsi5naJKxke9ZsbB5wUcsUuyF3fexEpRWA7eut9ZFmyDwDPq8X/8qRY/ifYoL
ASVKh2VLPOin4kBC9+tScsZOVYsxEIJStfyfVwCWl1WaRTO/lU1bHMYjKBGnRQ8H
lsKg7xR1GMmr5+tKpeIpS49nYA7mKDey2XK6Opd8ACTQT5qylQF4QoJtlCnJ7aG0
KGYg9KQOHWXuLpYhqM+tGhZp1CnX0CuOKcARqRI+yhd1THfF12PCC/9Zty9hKtAy
233Iabt8i62/iRc0mvm5EP1cW9QJx377d5yImjZMGw+ieMawWx/HoY6F/gEsVsdS
Fa1zHJUZZ22qpRYPrQkTzNn/NkzmU3TWFKk8pJgaxTKJcSusrq8oRADdVJ7rsvH1
mf2l0fs6j/ctS5wHhKD9H3ScqSgyehucZTUcnum4B3D0M0AGN/wOQA8lnU8tR7iZ
49tdKdRqCYqAy3sZlrEuMPr4rGEGXNCjQVJiRp5MPLXvBreSBX/nB2CyUCsJbtpm
SkvfRkD805fHIMgHOufSjHiwkG3tRoFDrKx+fNu1tKm2qoe2HIk1wkw0O0FVXVn/
aDAzbfIwUwFB9TEr9a+rR6H73erH76ZjEGFofzpDXMb7z2vw6TK++s/tNFhfAJ+H
UoE5fYzJjn+CFwOhvW75YDMxxTJQC6rhQSX9pJcBfN/W2nIbkiZp2pwnKZrVIP78
TcBLylqc+l+bv87AOR/RAs/f47O13SiEdN95pu8DwSW+DntOpgv/oVWhvuVds8mF
COMMPyPN9JdkLxVG0Ize0VaEIhHtNg8p9rlIfeYMsVZm1EqhuaTvwppRour87SGQ
L0zckZjyqZiV5XPavNFOIq4mmgYGt6+OsfL1JsbtiRinKBRWrLJYrlC4XqrMAYeX
xdowYa16lEoosdZha9esANb4DWvdFrRFr0eb5BTYw9w408xtHRukUjApAy5L0Isp
81V/tADv0B8MJMshHx5UR4zmSreON7Z8sCXNdaNvOyML1Uzo+1wYYFyik7v9slUL
UtTg2OW04/fkTYdA9KPJSk4nxbkckzVLUOqbPc+NUbMRHsAcwk9y/YpIIR63z26B
l7+SRacweYV+2W0jGq01tii7XF6d1U7j9Sh5c9TfjTvJM5UdrYkNO6u3RD/GFvjA
ZYdcRkjq9KTNFAbh1qXQQlerlh+dxtQYihUulKslRf9KG7jDOKLLP/DkWRDdkOW3
0k/aekCC5pwQl/7Loz3MT2mmGcxpaQPsxuWjMKLHyHKGxdsh8a/2Y/ZLCS4W/FL0
AyKZ3OfUYyU7VGLfPAFUPddIA5O72l2ih0ngPVGHuGWm76LZ8DQVFXmp6Qt25w36
wTGN/6yf/Z68hEtD3PpCMg3BWKSqXwTbXvi6wQXxie9R+a+dwkbYLJskpt79v/U/
5NcpBOBIMXhA+4efAGxbZqav33dOWXvbHa8AYTkxc6xwo4TdrOnjjKfrCuz5/1Hp
P+shuUK6v4rTv8sfmpuqzaq/uNTkr9zrHbRURrFUErYcjhM8pMsGWEfcYwd8BmUo
1YZv6VxxCENYNQRLCZ9tX3fTQDutFz2mvUBn8Wwje+cshkj1c3JU4LZr/1IhGI1/
gZZR89Hv7vRb26EzRZvcf4JdqP5BIpFeKGNraBUS6TSYwAqomkHEasvrMUvXqkso
bwnh8GVuuOXpaVWDeNl+kM99qcLRut7Vn+cqPVir3mruUk61Z4XQwOnM2Nnp19vF
rAr9y8eaFPqcldVg+6fM8ERAlhrrXMvl70iotp5Dru24KgJO7HOsz5o+sr8tpnBU
w5F1tuMBBmaW6C41IAZRHmarDDP5eeegkkSKy6LEW/7ve40cACplC4X38T7AWp3j
Tds3N6tCn18wdKiFzmmeG0zqYm5wGatrdhBQGv/cWKOQig1gfyVKW/itZkBKIm0d
H776hkcrVcnMNV2aCk3xhdUYo5J2ifOvEhZfnohRwTRzsfCx4aAfxJOw+suZfVUU
tX8GyzuDspZdYtrz2/xlXeR+DZn3B8G8GuOFF+DTFaqsMO5mtCDGlLzCQfz0mx0d
si63MyV+XcK5KOz70PmsTNIbEEEf4OG4KzwTTPTs0FsecsBSeKWOg1bSuedklbxj
38PUpiJd4R/MEZLbYeovNlgqtiY3a/YGHHvuHnN5qHah15m9MRAeHIEAtToX6AcD
LUPhTu8QLTXuF1IQBYAJ69spoL41h3MG4oTVU5wyh/mOObiYJ2uEfawp/LAprhfk
BLn9/Mb8G7nDUiruTj+L8FH0uHsjg8pNLMtfPgT5Odri08iebIB1GxMJfSd00jYx
2kgFGd1ewy3n+l70klN1rIGoIj4C31ghMWhdic7HYUFml6vGXOZjYtHkE/z8KwAm
R9cTOLl8X0x0dRFq1B2edU7u5ur7EKXQY+gsXLTW56L/OYq4IWuBi8091Pb3rHm3
/nUuKSw7e+hyV1ZyZZ7alJ2VqJ8VlBsQ06UDhbJDGhhE2ducg73pYJAD+LRrHWdz
LpUInjbtWQuOLuC3BLezi072JpjoxGJZxYd0Bw8em7SR9ce1wtODST9evd8ClzGf
0LVDdFr2ZSYw3Itgj20mhhg3wwhfGrGzasZVr6BNH3z/dWQQ+aKFtLU5hwwp1nkQ
qmoRofJE87LZhmrJVQgbNbD4TaHC+hKrj8JUVMjKyxjCA+veJdb9T1jHdx3XnXHU
9Rcl1X2V+nviC1VbeD9/SUZ+1F9u3apLzKlyxK8UJBB+s0dqivfZ2qKGo3DteHZ4
oFbmF6nMW9oLFekairMT4SpNr5KoiKd0IPy/a4Sxrp4mX2GTz/jeL8F8rLu/Hoxo
j8E5RNi/q3A91WTAjpMyD5oBxMT69/Q1TVClDBRhEndwIpRGEVIhPwGiTvoBz38s
mrkuowMoR0f9TQf1qZQqom33WQyyUa1JUAmV/o8DKZLc9zH4NbA9A+LenBh5PWQQ
qq+ic0E44JJ/w/29n5PI9Q5JCnht2B5H6VqmQbsvuGYfmAicFa6KgV/7EzO8gWrJ
DoXFB7YaLdkV2DaV5KbhqLEx1/K5EpN1j6krsw4RX/G8ESEVHdN/wq9K/Ky/jf2F
OBDV2gx581+SD0RaTM2FhRy53Yg9cGl903dSLX4GWQOJuMqw5aaCEDz9S9RqTbSS
EHrsOAcpsezpN7d9Zl5uZ5qoAH2l/eOv44LrY8T2wEQdRvHgXtf6bunGVaG/vs4P
PmNU5asYso88p5y4mi32Tr7ycOjrqDFw2NrCqgGwj0tUfSYyy4DVmX4pqcl2OiXm
TTubTqwbOGWPXFlM/xSbUW5Cw1fFaRotDwHsqRPXvxEEzF3u1Ln0ER090hbwIw5e
6LdgRA2+URxyjVwMBgzvskqdMjPc8Tb3KWhcwTdf30RFmr8X4AggNgxmib5zgIzw
PjeKR67uoGlSBh1WjNAx9rI+6xcMkpOXdCV2MIH1Czzy/83wOX74qWerAZL1YGtj
e7VwY2JcC/l1yJAas3pYOpfNp4sZddRp6L56cz2lGoqq/2LqPRd7s72iq7c9iI5/
9owXMSuxVIw2q5BmaiTEUgY+8xxyth9kV7m66toU8E11ucB4vkuajy7poG9ASY/o
+BE+SbPSAbrWUQg9Qai+b/57FouMy+kitk/KFVSsAg5yj+qcO80hao8IKX5s5JSo
8pWnAdR04K1qCwjiAH4JjZeTg7or5jSqEyLXQ542uME8Vu85hbcO++h4XId7smwR
EeygxZV9ANGFfmx9UT4uTX+XOHsJIMgY4d0B2jrVvtyUILxb+E5YXSzhUHfsj/be
x/lvoqR7345NhnGCpi8SDYuHdjwziirUczs9avDSuUB3d+t+unkZBIA1jtU7AMbR
iy+RVlPLCgP/FQ+JnNnTD0rui2mpx9CDNXvqOsajf29TuledrcL7FViavsCps6uP
7JNHwH30iy5IYaCkm1VN6X+A2isGw7xEGREKS1xNhwAUlz4xazP0JP27hrbvSy3y
Cp9nQkvDdxW5T/+Ke3X75Rn9ZSnXLPynzD4IWg94ZVhT2lHiATmh2/U85IXdRDws
D/u6g4K1pPs0cm23xM86GJQ7r669JDEKBrEtQ53WnHjqIc0fxt7n7jHD9PKAGoR7
nHuUG2LUm1dp32v54ftOgHcpFj/7TekTsYvi+Xceb7vmL8XYQYNXQbkUIzJijfH0
O8/h9yo8L4Chwm4SAEmcNlVxPN/GU9bhVqMcW3yCO74bwApvqTP0pBq313C864m4
DNC0ITvJKCbsPMmlNkyOYUxeolHWDE6CMde7vZWF9XExivRPU/Cs05yUZ3FhVQEW
tVGrqEgYWcTlbZUmEBX5Y72/bBFXGNWnUu/4VYf2UuRgyGiweOGUYvFdQrVKFH6i
ddCW2ulBdvjAFgxSP5mvziVzlQvGWG59TZLI/D61ZuxWXvB+iuVn9tF1Yz/UkkCa
VqWEX9JamaHmTt8XpZHlnPg8ZTXjzVIC8aSICxQ5a/+LxjouPP1bAkvSi3orlu8x
znxMXeDRb2EtJvEzleiMNJcYw4qbZU7cRKomSMrBJo56LPZ/SqnHfZ8iCWiSl1ho
gFmCaILkwviFH1uK7Bb7tq2/Mg1VUK7P9TLXs8rzuqpYgdffmqJb5jp4cFrAGTBj
mf3r0HeqgjSZuyfh62kqnU9uYDeE5CdIUxUau59cbnsr9LMcWoV8S7Uj0/S/Icrg
6EyuvtiPs1AV+CQQQc9CWzmumXf8Ic62fPrM6ImzJNxQ1Vwuo0rbWdK/cVUmqczW
Tmn6vg5TgHH3LUnWot6QfGq6mkjy0KSYvn5Ab9W/Dih69FrmJ+ygr+bLN5o3Y6BZ
mAreQmF5tntGu9wtD1jNdVumIdYw8l1qQE7E6J9f202yoal7LjXUVvTJulRuj9Ji
+1krQ8Z0iV7R4C3VpkxyF5U5Q3xmtbKyvECbjpHHJZLoV9rzvuc20V55NO9dYut0
qryZwJ3+brOuJBDnIYf0DzyuDMeULQVHDLWtJxINHnlvbI/GTr4sRQtsFopXoOgA
nJy83JxtK+KxmbreBAd/TURnaSff/OQO7y7J8mtGCWpI4KATQvwTyyROkaZh4RNW
WRBgDIeDiTsDT/SjWO4FDonybmyqe5qtScwYJQsWEI/1/cuBcudwFIqSZQOn/Aas
3qBX/xCOBPUyGFPDFg2rENarsNnMhMdhTIrR1Al/3a6MKDX9MpViZTEYWwr4duh/
4vjP8RdsTQ60436OEvBu7EjtCv16PU1A/PU100ZTJL2xSY6sqAl+ZyfcdJT13wSX
TniPbS+76l9dyeBxvrF88UQHm0g4LHl/nN+SUhGf0fo5z9E5KI7Ih6hYn1wHXj7l
BrGf4DRkwU1birNjvSYYeMl/bkFbLiiGP1HxceDst8kcrd+Bdtj/T/K3f9EFiudw
yLN5iWBHn1ZyyfVxODa4W69aRPUflNFES1T3Pmmj9qauv2L/nRFoNiWa/B4b3kVJ
sFQSUel2B0asPvTyXk4wIbmNHEQ2MMK6D+6TMgBWyfQUoM9WewVEu3Re8FrQEXrp
exmF++OUdNA11eK+ix4nxttBJD4vLmoXI8ezM+xQwT4oTXEvLza3VvHX2Svjz9V3
acrxNY+6Cq4aeBSNHTgj7RGHY2yd8hZ5tLiGRRQBbSt1BTM6w5PFYES98Y5WOg95
ELDNNVwVK5RhaIX2BOUeMCFvFyrtHZ9h/DX4UAruWlCVi8a/xNTtOuk1grRIp4Jq
cBthYasJ1D511ObHaE7mM2sYjqIN2LdEOjKNCVXAscaLVVOtCLppxZS54UB61CBQ
MTqXcNps82unRa4enSaOe6khAcZHCHAnT3ZXKLHrMOm0IwKIz3GeJTfOK0y3BMyR
A9jTmspoivAXByjcDwel9b1JebN39uxtpuiXWoXvgRUGOBjnFz/upPUlLZgZSM3/
TKbTc0SL0t8Fw+c8H+bvG8+CuLuwgXVi1L13b7F/JTWhhWqKicpRI5eL0hRwBvaB
9Omj2s8n/H9vnFEIJrCsivpddRvwWHqomwB9HSnC/gC4L27gO1vStsFSNe/yQVDA
9ugq0oAa1vYUAGHJWayuLgHpc72QXDHS1AXiwo3VbVzy1P906KSPE/icQAKsGOzA
Sy/fW8EP/xC6wOYMwZBlaXa5O67o8VRi46+DC89g3T5/SGz+r3yQnD9CkVTXMfm7
zt8Sf2s3uXQfv3K0SXSSzB08oxD1jXztHlbTci0DbS0dT4qhzYLfLPKzX26fh7Cu
CW1YPaKOiWSsALbsEyVs6VEW8p/LLoxv7kZrx8adNJOAsd/yGKfwwQAB9Zh9BzRr
B9UXplCmqbGgOaRJfWePRPAgqtACzbFJgx+hi/Bel7B+O01te66x+PsYOunTIefH
hShKghpmMci86oWW0PE2Ye4hGwVCMwwo4f/G4ain3I3EWBwMExOUcjmlBGGKrzb4
uU4Uwvsxi5oobfiHJEiFcO3mw5W8Eje7wGnlkgQ8XStU+sg79fOfZ/G3wht93dJF
6lX0mhn0WOFu0QMuwB7pJFc6AyWloH9QHGND5IYgSgzmJ5ngAtei6AbsfJ/b1Czn
R/V+UdzOcUCWGYzLa1Hg2TrK4Uv3WKwRTGj3yPQYL6VPt8GtjzmSQ3Cr5tWIpJML
OCXMGJ8g1Vciw3Hj9HPa0O2xGn3hYaFn0PFC+2FaY+IoCrjPduVdYy3ajzCyvRWP
NhFlnVPha6N0jG2r/szkra/ezZdru+dzOGSvHwtTXroXQFYci0ZH1ZpxR9Zxo9Ra
qr1DA7h0PXHZ6SdUQWPZNX9H1lnPeGSMcG6gjPfwjrnRx+B9ZZfykBjJlbPtZhjN
4dBSESE95tYaK6uI8m08QbDZPWJ1tnA/FA5lcF26wW4Utb6UxnbEowQhU61ZSn5i
y4Of3mzmjGlj+TBDpTodUVl0bik8jGyhwo3WZr58d3OQN3NrEwEAi87lNnfOEJJU
z4lvkaFb4eVZk8T4sYPH6phxqHOE33xKMjuQzsuP0tyj1xSj/FaA0E0r3GlE1XI/
CrdaUeLk8y43+asgXlUY07/RpYl6z5ejE9Vyl1vqb3jiVQphD27dmZl9BcduLjzY
e3lcajM7gsffPGqQLL6LbJrRQRQzVYFcCW5I8scCtc02YIxoefBU6FV4ZwIgd7hE
IAjf+I8mYZRHBZ2BZG2o7RP3xvSsQz3dd9XiffuKYTMVyWGkT/ASelbf7n1A7SbB
0q6jDLN2+v3qTtzl1NjXLmJNOQRM+rcs9RN65+RShrz5RMxCOAYnWETkvgxVN8mm
MS5UNqBlbjRBy/cnoEH1dL69elCxjyrNyIGUnJLOFGg71hgOIVw3Q36JABCCww2E
CyMhlP0lNYDgLf30hVx20UrEVwb2gEZuvAzV9Nk3gJ3AcJcMTLDoXABaQ1dZ6c+p
fZRBCNzTaK/uFfxenyPBhTS1Sm8WS4u0e9Tnu8D/b3WcB+HG3tXUxxxORWdLkQjz
FLeflDekDN4Ewp8qcKqpomdg9e+PgJkPP+J7NghCPcTuBztSXWnyrh1kkkeKkHKW
FiWu/klGVrLPj4xom2l5R7mfxbwI0/BdUaerNqYyw4hvU4zJmcwOHBQu/m8EiDMa
lEA8jLeazTorqLUwsgkeVcwbnceUOxSQ91NkyB2eTsNv/i4cVTDjJTMBu/LLi+oW
4UGuXrE8ZmWoktImSRVF3gSe7FPL8PeMKsONRUTGUomU7nefcuzOWmX0TiG2bqZN
iPMII86g/QSazw/eWaFowxJkDqsIeqTjjocUORrHfg22gAz+j5PvqAsEienxlRM3
Fu27i6iMcpfQV9UwVFuhrqlRK9Y6MeN00+T9+GlsZUuDIOlo7ypoDNbqJW+W8vMj
qUAbzAaFj+v8xn/Ly7a69jYqurgnVbH90DR7dctSimC5ejDyevgiRi14pRxOraq5
fpA6rY21z1mfK7tWxBsRq89h/57p2yxYIdS4w5yWFHTdZp+FFyyKwHKatH4rTS9C
3G3bKnNxeOYay3RNBTyyE5U63ki4zMxowxDuZ0me8NHfB4081Qqb3yiknUJQLC3x
xjxxC0xNBrx5UJ7mj/7TdGGjJvxu55QOAfVNQQb71/XV1AmO3+Lp8/T4Fc/7HZn7
lqPfm9BkdXN+xFB+PE3QmZeVbs4uE0ZQJLedu7aI8XEXpjryFaf9KICLrXNeT9lD
t71hhWuDIqKnQCY9H0xwWpzp+NxD16yJR4SbgQyI0w4ZNjrjnY1zixnA5fYdrhde
saDcr/p4i9nGLMv/ZCnUF0kParr/D5k2jZ85d+wjiA6T1WSWlwJ1b+tUo/f/pR+g
kgH5obaOxc55K/RoMd2bOM9T0p8AJ2W0r5X9HRGGaeVumn2cVIQpBhRulHIf2fqu
5Ub7yfJBqCM/B8aquO5GgApHsYZ8CHgjv2X4lLvB4K5hPAsGNL95AoQAK9WtPpOL
vQ1kSNVdvjpOCHaor6RL3KxTab/SPA3ElGvjVXsF18rdZ3wf7XLieQ7B/xzE2A8J
kkpj7MDyd5cl3MxUsq338TO8sUZYdppasA/p1bY/aB+p9o+x+NWqDkAqPS8aXic1
bYl0sCHGO5kbV+X3gCO/QSFYS4CuXqgVpABVn86Rf8s4jafuvEO7JBijwWoaqp7w
cII6ZHcFU6SKDNhVtDNobvrfnxRJHtOkyKfGliT1qooJXQe7bCG3+SwpQYowbXxt
iPaoXx2awBMq6K7e+eWHdmlmG188EZJQkA0IP3CLhWv91jjHiF5l2r7GN8QgzxiB
Sf7A4zxGfPikqjdMJ/vx3NDt3gjJ1LQ8uO79i8nYe2tKTIXBCyrXDf70AYv1LwT1
0vBGc4KfbQcr8+KHG+aAfxYNyhrKd345PbFMeDVaIplJ6S89rHZNbOLAT/nZ7rnK
hSJ3Ym4hMlzRSKAevzR82z/5qpSO3dhKhZen/H8Kasg0PXwk5+03Jnneid49sP44
WxvIBVkBcofxoVzrAZ8j3TmAeR98wBqwmy7y8KSMFbsdEfOM0n4nuEegalawJ0te
Fuf/fRVpfhxABSr7fJX6m9ogso10xb87/nzsWKv/KZswkDasB7vgvx5LQ4+o4oJk
rgm1MrbeFh5tOtzcN+ToQFW+DPZHKhp1fAUItnKHHXT0m8TJ+W1TYyt7JAd/t8LT
dJzFRVVRLHv9Y/7fGdSt9ThFld9T/wUgLXT/fkiBBUpTv2uoXs92zpv8XSWtWew+
PtcvEWwCxP/5jSagL/MMyFfV3QrnmrreFyeVRkd6VkD1zIYrZ5jmQg4VeFirB3ib
MJyO/ROyOa8MM4KQawKhlRPvMikhMqdKY3k5cN5LU8uv6CiQXfSv3ygtdJMZ3UQU
Oa/ZoJqOXJEwDLa2Eav7JVuIhzivJgw3pqRCUjlzeINbFCxtfQsOTmPBtfIZ3zNi
TnZ8l9mNtFnOuaJ+X0Ugp4upVtM5vO1lEMDpmWXO+0b6X1UsFCz4h8o5s/Rc31rx
1vAgBHanYOw8NBgbaXkp/Fy41XluMZhTP+T1NCd17DydLsW+s9LykeBg41bX30Rg
1cwqjx1zfLd+cmEAa4CXgdPbydypC8qxOACNNgGBjZ6o+PGGkh9dG6pmGzXbuQgn
XcAnOkYrbT4CG+FOAT9XhVPtIpqRQLXA1rYR6CHmEoODnv+bGEO7h/FOOHp27dD2
BF4JAuTIRpWRlKie/FfTpUzAWp4dpCj/VsYksMI0C3hScdMzw2J180KeVo+E3q+E
PCIFSgBMftjsTBLyanupSF6jTuNX2jsADzfRsDHZR7k3NoBJYnIXZSRfg0Lb1yzX
mApn7nM9NXT8hOJ6HePSGp0Ar/ERxoGalLRfTOE+hlO2S8CblBytb/m+gIOwD49z
WmvELR71L41SuZlbDxwPh/z5pPbiOehzzAa4r0qin5JfskAtVKiwPt64Qu1Mj6WW
qLQbwFIH+exxdnBuIqAhhw1YgqWU2bXyFT+QcMDhV8CTdTIt5hkH06Xig/KQVWsm
chpCEX9T5i2PfTS0vLfdCKEM26bDmbhls0vDt/+CoWgfZywfQJbdW2gSF1S4sbd7
4xKxY4ZkFq9Xl1F+XMKPlgfokaLZpP91OXaJSQsz7dvByD4Ke6ZFvJyKv+i6uOZH
55mT+XT5PkDTgSmDcQ2c5jSNTE2RztnfZ9QXQXmHFAydtePDTf0nEMcOcn751HWQ
Yn/hTVoHqdODKW/SU7JgyKVow2Sevs+vm8VEo1XJfoT14mfhGXeBtCfu25XYI3LQ
/LZZ9B53NZtyXOWulLYkgwgFdNLnCbjspE9IOqO/KJsTq3Id323rQdZiSL9EPQ5M
ZBq53iSzKyCL5suK0g/YE9tt32Zoc8uCtjG4UgziYex+WxOCA5SMgyWifVB7yFVz
4P8RBDWkZrVyCgY0kCrD7aKuGu3JFbxRoLzUN1DmWl+y0r1pr1MS9yCg5QDbMwR6
VZgGlL/aD5oqtrvafaXTETXsEBIBepV18Y+hhIa09WKfjGir1Kv0R8mdshYdjFE6
FBrXJ4qDyssk68dJBDl8999IqzaiWMVqsjzLIRSiDLikNFHVYLAlnq7lEO6w3dVp
K8Q4E1rSJtzLqBmHxffF54FLfjWAWZU+mcBperCOFiqVIfiMtMFqof3tfBB5gHjU
OLHXrVKfEJy6mrKBzCzsYQWaX6m4Cq5bBgttKs5TeWXrpH2lIEaN8ehiNcMwz6xW
kwXEv+L0PGONjNeDVCQu+ll6YLDQYy86ExSO00TfVQ3GQCe5geoOw5Q/KjClCAaG
QiXK2Du3nQjDkCf95XcnE11hGpuLsU7SRr3JbVp27el05Kza06/3R4OSLwIDrgf3
pSt8hXgTU6EmnuGsyLE0nRAoYt9/rg0VSCxM4w9Zd2Q2DPbE51nzO7rjMWVnD4CD
MFL5k3XP/zBNO4ScvkFjtyB29YjQp/7Gw/RbY6moomLGcyGBUcvK0T7rjiWo+lia
k8zLg5ifCt2sHuTo/GgIvIhKEAVixBPv6+7staOGeC4dEjRkgkuqH3cXvEO4CAa8
ENfvmHBpzrCyAynoNahlnxP0jw6I7fT99LnkvIIrnVsv5bjlNJbU3z1PTL7uVNWs
n+BlmFpK+HxciPLcWgl67Dv7IYDJEk3oD6m1jYdGwHZhacb++CXrOm5m3CHtd3bN
CtZSBSN036H2HVk7fx/FcXiNXFUDVwbimEhzLoIxkhLeRu3dA1WbWCvIDJ27/q3Z
8ctIGR4ieBrmn61/JyS4digpkNFM9ju1VOaC1OG/i3zQrKY6gBnvJGp1+VxkL08y
G3xTb6hiA2bQGw9olJ9wqLtHih9iiTefYoVO0MkEFZ7qLmJnNbZHAdTU25oZlgr1
q1bD1cuWtE6vTQa6geGmkXwAylDLLOz0P+ZafhLJqWGvNxfHmi8G/W0gFRvvk/PM
14/Slc1yR3MgUcqgFwLagOnpd4PV4RERJwDF5U1gopJXr9UU+y/xgmYK4Lb50/sW
Py9aom3VCZ0FhxC3/VyV+tLggfm6kcGh7byTGSs/VYdAcePyYKIrQU9lB5M/fNqk
7mYQU5M+7+J8vWyJLayq4sqUstbxsziHs+ZhpIwQfItws4lGfyY5A47jMkmkINuT
CuLyBed5SdRZ74QHqzuZud+5VXLuNbrUBq7lII2eaJuBDwuWk9NJTCwjNhK/jjim
S00atf5lL2iKTXCEi9wrSyc8H3Z4/qWUgxjeKTcX9bQ3RNnSit2zYb9Pa65GIN7Q
lLNt4on25sxBuN7EupSFMWs66QYLGnYd4HMNXtknwuiXkTKS9YOVpvXTA1VR18L/
auC5PvN1wOoQDkZipcRJuYeAkVqvAX68Fb0PWXaD+bDAJhjpySC/WzMkYtnmAGHh
YDg+87XfmCIvokKgyeuxpewSpntba947qMscgE54IxLN2Q4KRm+TTaiQTE8aR5wg
0eQkQa4sR/Dr2vIFF7yXUAyx35StOAwnMRu52IM8VlgX1SA98g50GCdzoKkoKuZ+
shr8j7eO8Wra+yHRFVwbagZkOG3u3UyS6KwtU2QM7j9t6/DmaUR2ev83qeYamqay
4XVqMewGZ0F65WRZbRsWJpfgFET0wCEXoPggDnqAfa6E3G8Fj8GoNmitKaOH6zKg
erN7FoBxYA+SIgFARQbNnBI0S8znWdffnpJRJySBDMFKakcO0luR7gmIKLBmXlCN
VHJaCghJXIamQ1NMTYCrSr3sFopTGCrcuciQ0UFOlCg+Jt2+NtAIbgMkLSjiwoAQ
96NlxTHcZx3eCSv865oqvwYfQxUlN3KooXOQDyYVew76ZlvOSjxwY6/BpSJjM1Ae
Ccb+EJcynNxAn5haRx8QklSolzzj3xBTbw4fJvpSXWKQG6sBo/qhXe+YxJXx/XqA
GFkxbaNan0CxS56QQC3YqF12YFTWH5KyuT0vduiogtkhfTuqWMEPKEF0anpFlTOo
6QHXG4ZRMvqErCyRjM+nljXEiGwlfGKpLkiE5PNFmbTGRWzgkqC43gFNpWbYp4RK
OkPszvNZSZJrMOLb1k0pph9GYf+5swiiM3YFsPucJsxsh+f9noZ9vYjxekV0Rx9g
0xxBOAC/lyv42hLeM0MolZtl2+r73zf75g15qy1I8JKMiJVnoE+ft4KPQwEzICsd
gsD2R4tzpXyTp8ph8OSrYIy7Y86QVsnl/8kG+5cdIjjDnTaWTPFxNR+L6L+/4oE7
zoikqKCqqQIVnMtGpEGejxk404TVefSI9eLQFCU4zYM4SZpr0z2e05JXr8uQY7BE
1KZ7/4m4xJ/5s1r//s8ynpYb+gUuBdPXfv4Rh90AzNCxj55zE982U/tXf3wPGEtb
z8pmnSHFWLZcBDOizydthHof2r4x4qs8DSSOF1gYWmDBDnfaDceOdceP47n6d79X
IxHgD/jsUBpd76hJh8/0sbfW2PBJOxuj4jxXVZsT2XTvEYUrrzwJRWCt1iqGcWUn
rbr3EE5KxX/Y65WtwDU5w+HU1HVbOyJfXUrbI2KWwY9s35MpoiGwdVMMuDa3K+dC
qYOQebm0KycR8tX+aZMQQNllrhQTX34PaLRd/fZOYIiFRTeVFvYLIweHOhzolGPH
mgaxENgvtlcX1A2yJMLuzhWelYHhN/4H5Z6LC9V7414G99QoJ9lgDo46PcR5gMFZ
Py4H8+YsCJ9G+SxISidRPBw3jRkctMeztRFRI78DiT0MudbiWBkK7U8GJo+WX4w+
l5je/0mw4XOKFILKPdNK/hEATZhTgmpwb+MVte3Rx4PZCCotR/lWuyUJKIkW224d
QAwtlx9Xc7O8B8bbjqEO5FyV/qz0w3h0yCTWRreiKuNO8VEm5T3MFltrKPhUWSpB
ZG0aFMDpfA6/T4PSSlp58tiE7YCGtGP5xVrLI5A2+qJsj1JeDKKHV8aGSg3t5aG0
N+TbPgxWjeHJQigj26wWx4ydaqZinFM4ndaYMw1LC+Sg1FmAucD7zoPXd/wUitNP
BEncu5osh/Mdgm4q/fl8IQpjRfAtcXe6/b3blls+Dqx/TnN9aHtobi5esTM7Byn5
hnVAyFGszaY1bcHGg/IYG8RZv0NU7crMtpxyt7P8wnhBFlRvTPTVdKj6kyoMpiBm
b3/xM4zurIgN09kaGz9zERYxvplg2CIgH8ko3QD9wAsp6/LflpOR/BHRZXtR0UZD
ox793kEFw0NKa/rTnDxtz9aXiCQpWO1DxLLt8eqnJ+w3GDtdhaMi+P6Hn/Bef1Eg
NW91CJSu+tSmjQ2bgIQFfu1j2POETtZyhi9NUJeTkrURi/KMRybde4BkC0zBhuR2
yHYsIkoT/46TwLq+iUSNa5YTB64iDFQWp9ODktNZZTyfVeiUZQDtBctRLL3cgkTE
7f8TTiCzhNV+NDRAbprdZ0a14HakJRqT6Gk68CsC1AOBsXnqOfyuUVtKVYUQG3kc
RC4EtAo7ODBqe3Ch46Xe3Dj28FR2FWVCKFso+7ZelBYy3aYIo274wD4xKL6U0gbg
eqMzUTcWs71510TyqYG4n9YXvP6wvk7Zsu53IbyNSpYYWBDEjSsUPS6S3X+gUFS1
h2+CdbMVsrB+rFxScqZOzn/7+8js0fnq7r6gyE53Dizatq2IFpAJcFiSNANrXSe2
K4yJzihA9RTTN6AAFwmK49EQs/bqmkHrcAC4cRCCoPajdsXWdjev46DBe49AmwKS
F7kHAErRSW+njYRyfjKTZrHQWGgnNMCHGpuOL9O2NQ1TrWs5mOhQpEmetSQ/VSD9
CPrJB5oLBIewwmGRVdbvTNeqEO/bCrRPFODFHPSVq2m+P14osRuskxLgnugOdn5D
5wdIjfu7HuPlujITjDO0IxuUPhUtXbKKRm0/2p93KUv5zdusI3pngpyoeI0UpFYb
JzNMbvgyBS2jVECeqFrveWM7h8HLhMmaJNUQKT78eueS8EzZLgpVYnn4MR6BDtnc
i9TrrR2ZPVpMDzzPGylEYT/ZF8MMMOnKCizw2gnrmHgpqElCCDxXE35hAGQGtJpz
mAf+aDzTZR0l3+JlySWSzasZjOAKKlFRnOD3ViKhLFfY+VNFeiIHixGL1XS6V9Po
uYEi0KEUfgQM7FnPg0zmfLESTQQ5IwzFlz244DIcH5G4CIvRAvdDxHCrbUTanB3u
nSNt+PndXtFmKn/OmY9S5jnO6l8cKnJQ78Z7T3+ywMEa/dge7Y0V/W3yJd6Mo78X
Sm/uvhMdhC4tQu/lP08FES8rEFVhfeUubRYCJzmkp+PAtF5np/KHuRkUfiQjbFVH
M+Pd+82qrObHJ8OKHENHGLuAtzvr8yTrYl9W11mfgNeJReWSZIVIv+vV6Nl65UAV
QhNziAG7pKYeMQ6zqTHSge48Y9cyR6u0jSdr5IsleCoN0FjT1nZKV3gtKAGauuM6
kYc6MrMLPHKrm5q0q66aoWaRNW4uq24BmxV2uuLImmOEn7QG0eJ0dj4VLXAgpAQ2
trzjNLN3nsspcDx8IVk4soLUCiARSMaXdTXTc0tPE57dPe7fr7dTz/Q5OPfeA0kA
/JLnRCIKwv/Wyoe3JdCNaZmUoyJ8GOgvePAIg1uqTGxM+mSct9SZs0CqTyNFnBfO
MZA6SmWuGFToFMuDeE6VCvn5tXDschPPmCD6XgfSyAavKxpUMyIi6Ne7Fogf5cgm
/rokM0evssLynR352SJn/u7+2tfwFnCeGNtIHARP0aSOpqminT2hU3iH9x+e3fke
qvmzs8nSbkCuZ0nf5UOqe2shSj61rT4Rd7oXZUkLwrjsLbMItprTKgAuUwy6wtlv
9elS/7fpa3IY19GP+Yi4WqWcw0ddfklEGq57yQN+y38E0d04CghqYprFI7DEHT8o
Xu+qu4qOjoPjHkT4J4/RWyFgzxitmuUFIRpi0Z2AKzS7bJVkMNL96XhxQVZlyVpG
iGq0DjAdlSsQeKtnOJErSR9JLa7uPSd1fH5w4VReBSg633QbCc1NMSzjJdjleMZA
0m1UEwAKg7sbplafgkNWfXHPCGuQIWZ7p176cRkqjD6GNZrtX+hpfdDRGHQL5Jt9
o4kzeOjNXERfsTKoGa9D8Q1Ygj1iZNyZST7LnO9DOLZLwLVFFWobAhFTLH1qsnGt
AV1bbSeT1Hi3GXmzHqiS1G7iUalvbCeORmDijqT0E7ko9UZssMyDcv3ZjoOcddPc
yC/FM9fIJp6DmBy209o2l58gNnXnnnjhxltm8K4uTZdth+ayIt0RXqPip22k9m8H
Roubo7gfQP+N6DEcSm6qIcez51JzEVqWJbc84GrbwReim+ZcwdkHbKOiGw4666GC
LOhTaCW5/WV48MJyZotCYUglpxW+WNCB31knX0XkcyOMJgOWCSal9M+QqdSmdYsx
VD1lZ8vUyMByk3y0ewgFLGAoAI16CLbI1tLxUcAsvlcI4OjNiOy+SC9rMw22heyz
AfREUuFk+AVPWF4SguGF8iqRQh3ZFNziM+weu5rYWlsDcWj4zwVsr74s5QJ1xr3J
BmrzmWq7quS9gWwo/jSmc2EFQNr+b5/za2KlV2l1UZYozGi7lkbE7ptlUfpqImKM
MgG7QtSo7wgCCeK9LjbhTKHL/GXxKMyxHQ+tQ3OKvPxZj98zIN0YE9yvpGHz5z0t
uKs676u8s2Afb+g8vY9ths39avK8+vpiQ5qlHiFa/A/L9WB+9NPZbGrmfFghljIP
9PoAn77NoI6jJxvhyEWevHta0D8awEXXB9/TPZrRAS9xeHqraH3zZ5i6u/kauvTT
NKTsjNHHbd64X9hfJgNKjqEj43qIBllPSw6SE7ndeEWZumAT9DfbFWr0nX4OCkRs
kKnRcEax3xmvPT/HyF3eOc/2D21k35I0TD8TFldjEt6kwjES4dQybkoL9j36tbxf
yO8+LCHNCcxPvhvaYaWELsZNxiiTMKDykUVEPeIMYzjshuYR0Lgu6V6JpY5tymA5
Bn4Grm/Lq/LUPf4tcfH5clhKAkHO1SkM3FKY9qtH4L3lSbSmrd/oGK17KJ+PlLXR
cmWo2ToUARCoB3g8kPknAem2R4HgzOXdNcK7RVl3+X1jD4iHTHMqQR90KmbNU0Ob
KxQnezgQnK07j/cuD+YVlPam/urYK/HZs1d0Uai64/Ny2c3bzUZ6rfGrMmbmnKqI
cNQFpRne14naxCSyYi2oiK/Ib4TiTy62Ktj8WmtKETuAIhhMOadJY2/JbFmNN4M0
7/uuOsQUYM06gZot9VJ1HjzKCgcqsbUEF/JaWQi+DaMJwAK5DjKhZq7MArg4b+oG
4tOI+yTMifoX6pD4gLOJXVhpTHvF2vHSSeMZpt9jXXGm0VdQJ59EY+Kdy1aLpuvI
In1Qix4rVuoHS0UpX3/sXTSDjy1D8kG0rZ8xAAQxP3Z3q6h5WMXqMSU47raZUarh
XkKK5GHeEM63eqrVtQ+ZuDC/6zKVVjgazc7PEVfsAB3vY7X+oXAQxpBpxAgBG0Wj
dLYA6vZGBHSNgHfqLxLv2aJ1Pb8uly4sEVDA4NbEPa96fKS9mUHkwQdLtRpPc6jh
JqiyTRjAM87/9IGnMLkrvLr7HioXxmLUifMXi+IT8i/eJ5oLHdJBlfupXGg20dyx
kx2YXnufHN/6dG05WgfTtM3UF1WuGTF0lZTqL1DAj0aEphUV1A0thA0HxQbdmQHO
ODyuEqtrmtwm1dC8MHxIn7vuj5itsdFgOudixUuKzq1y91t/7cbt+M6tkWMDzviy
Bb2mHD3nzeughW1vXgkX6r0yiRL02kDSRL76l0gGuYOQKjeaar4rvCvH+5WBKEIN
CGJpEeRYe2MZ8QWKhmLnnaaEqISZ1AXtVY+uFzPh6xKiqW8MLusd3sKoXtT+JS4y
eazLq4BbxtKnswlE/mNN+hTCFY3Zl7dFgAeywn0gBKTVB8nq3nw4HvvbbtoVFAqp
RDLwBxbqZ6uiMF8My1lLhRoc9WgFi5FKuLKD5k8PB+muEmPyxBFQkrzcOLcJBL0J
Doq9CJbL/tp7dDjjypYkYx+NvnPkX6zPO8H9zQ4hfhh33mtzqiMwEcfwxXTXc2Aw
ofHNw6RyDZOd0QZEwiwAkW+LbWtR/iMQcQNvZaSmEFD72HtWZxt08hesQWCDcoz3
LixzImHv4/coL1byHTP3gvz0t7zDuLIT18h9GH6/DFnIbb04zaDa8ZQce8U4kOCs
y+uM6L+0gvTcC4Phw5ZBuS8JN/FW7aFksdMcYWJPbJ3s1zIacprGBdDwaVa+oMOF
6RPTtrQOVGTHFL37WpJN9o5OmAL71RCwI0XrzgydwtZ6Mts1Y8wC8zkVshJgfCrM
8rjAKeO2mpvTNpyP3t62AW6uJMUv58zuCv98SNlFrLmhkcWDOlZI5Ra4n3EGuLqF
Aaa2H+NsOryDU1mGhSOXY2V/PUE8Vlc43fdc6GiTPauc5M2T46B6M2Cm1UAk5gy0
R96dvw3q5cEs5XLb0TABAHQd93MH9i3bD5biga/69tBR5feXuqJd8weOYqmX0wUJ
Zy522Mm/afSQdavLbFS8q1/r6YzZthxBzcCcJVB6Joevbvxyx2omLyObhSeKA+5H
2hrcIhzVcBRPlNGTYJHtgoUAP9638BOC1ZfNyyUvncYi+7VTBpkJsVs02zeBicCH
CAv0AyY1w/dfRSuPrsXQXw8lZpU2p7ZsHXJ3GkTmKmSKbpcS3mhAuZJzGFN7Uz8t
tZAR/oiTFlufDb9+dz54yDfHzLOQL5NsM6cltJLjOS7LjanpclLMm6ei3Ia7Akfr
QIlN5TU0qPh6C2sXAK+l6Y+xUzNbDBM2GCDzmulJLxjecEY4MJjDCOg9YFdFBZ64
sOkKY6jhJx8uiU30hfyB/tT4mwORCijsxoJ/F0+KfY3dG2P6Q6dXz/zdXe1BMeoy
s21e1s4ciCMGho23XVsCrhuqXIQ+ayOSARKG9n2WMXTvJKLZ1rflmeH09Xhl5v7v
fWobCfkPlTPdz2x58WVFqWSXC7RKSzFsiUM7gWSNUNRnDE01CQF3ogLoiYFITe2l
+i14RBGsq+jGNxvUSnIXXFAH9bNBu70wKgif79ONc3QkRRxplx+VMoHRT9Y37q0I
M+GWM92YaUB0QBCfwpcFknTyfP4BZYrrOnYfune3PZg68JWgMmRqxyvzgSUqQ38O
FdvR0C5qfQORsd0T3wTY8z9nSC3rPbWJ+L/nVZPtgf5PZGlVYwWjv59GoU+/DvWO
z7/7ZtlByQJQlOr4PVasZXrRolIdxeOrtrNO9WdCRKm7jk5v3X2Ia9meCaFXdQoQ
VpT1t+8gKy1X4FDT5okuNsc3ze/wVuI25jZYeb4WWz6czA+VB7Y/19nD29bPIX5o
ra2FxMmv84X7vy+yjQ977GGVf8X0cwbPkcivVVFlrtymt4dFP/dp8A6dXgWRHS7b
/mAkawCBF4BlNb+zevQuBlrfMybSFb9xcG/T4J7jO5BIRdMKdFSqbx8yXNVjFC0m
WI16f7LvqgvI4rjC5HJpPCeAgvo1Mp5My7RxZa/UnC3eC1HBAPDqdUpwKlDdmqPz
0Xh7LCBeFbM4sfJkSldEStP6yhD+gaLLGOA6dw/SD2VUcuq9F4iYv6OIm3I9Cu9z
+vuqETgi3AKvKSBmStzYf3ul5HoBeAzEqEqun+3WiUsDV8ybjk3IqHz9lvXhAQuQ
qnDImPc8937r6nISNbgJk8QzeMtKtbGlzfR2SvieWbOs2cW6LPe2Se2Q2kRFZoQR
TIB8IXf7092JosYx2iSs/6WWH7hwd/6eEU6jXGGQhCHACARnC/o/H/Jk3f7DX28I
XD1IpCigpim6eEyb2uNv5EiXj9tRvOSSp8juz4yppSAjhKYN0anEZ/+teyzOefYk
o5oFN8dGlRCttTNRkNRN+o0EPl6rXfKB3Ba74KSVwUR0A8JbxY+Obknj4wjBCNml
KyJO3/K1b8DIXEdSaMMU6e1xr71OZNmC7rUQRf2q1F70HEP1OuEnurbPzqwTAdf2
czIvfIKju9FXcsPjmNeziFQebJgkql19r+Bq9qaxSkPKUYRZYoScFiqZKO092LPS
Me0uGSCJobxEur+H3O2oRYvuDp5e+8EqadKJOtpwDlBhs8KwGur6xWcKLzunQA7V
kFWLeNUJNMmQlK2xumYwSjq+WUPz0TjKPFjPM3CkSCQMD20IjRadZX4xbjt72mfn
hwr3ybBl6VmNxB3DPzc4xGOie8AsZOiZr6r0NOnu71UHIATT3iuB5wnmjccP8lI5
SwAWJaUW7tkdOOGGsN1T0iHGMgYAiQTkgeCzoYj7ABBafMGJhUSvoMHCpd1ykHMK
A8qYOo16YfIViS83TRbAWQn6Gq0IvGubm2dqYeoUu2Ahv8w04xMAN+QbxLVinJKK
wS9hAeai1FWqyTJ9wkkd1kzkg7wOWh2dUSJssMd4kHMWdZ7R9yjUrEj9MlkjsjEI
4hiJb96xgCjk7ISUxiAlWk3cLCpiWSejlos3ML5hnAMj9vFz2IrQYgZonPgf/TaZ
Fg+kMjecWsjhSDrvUb2boXkf69LOd21vZvzzzvNC85H9SLPdf/8Utf7nApho2nwq
Xlp1DkgSMolauJbputfzpGYTsh1YdlJP+wV8VjXPQLVvLocTBHblcyaXM7hYxr0q
MhdU5r6h2lf3mNxZ00NY7QrGh34kGs9Fws0ifGeKnwnpy77gcpgdq7qXFwr5XNIs
ej73SGFNxPEn28NmoJuiclnchwNiMnC+nMg1iaY9WfgVapFZEP3k7I61HaB053p+
FjJ7r1XesR7BVdqmqq9CAQ8ZCqrIvXseyhkJuF3FvohwHKMLYXgDYV8zZJgo3oFW
fzRDPvikXiVSyqLzRICsIy2c3AEo1uf8GqoqVNwLdDbB7o1I46HPv6qzzbZp1QOQ
F7aYXT3dpg4d6MSIgeyYacSKBZ0EUm6DMAo7oVXeuEHMHEOA3zckFXYU9/M23B7Q
SEzPbHcPUIXWwV+e+5e+mbdwjcYlZOrm9BxXpTlbyMl9ARXsRLpbo9whjJjqJZjz
tRRsJ/YomS8RPcwstMcFDMScP/bBD+5XJ1PSoKmTjD5j+cmjUfmH83noD1dWo6ZQ
Rlp4azwL97avoX6uSEBqUzFcG+lvaRV/29lFlr1VdxMN9wImOJ+EYws5eo/ZntRr
lSRwdA1Wuw8xDOD5/BLfwkDxbq2N7/whQZSx+tLN8/hGOeVwwuz9Z1Ts3w0yt47z
VFatkj0wHbONJ5sp5GO3f46KuWX1yL7HpJ/Nw84BbKsmtDdFCA63UU/EbxQDXJ7i
T521mhPIcYSy6vaH9cST+tm4mN7MQwZd5o4mGbYn4ZW7u0+oO3VAMX3Zoz/j6Mt2
WKTidFJice9pR5DcL+giRPOrY6Vt57lgZn/bKoQilWXoQNuiHENAPlL4OF4lWaOo
4ma5M54vrKOW18hjp6FiMh3fg7391IVCWV3OhWMHHpI6EBoOw2nV8ZSwylkrgPI/
fbZdkNUg7nZQHoMKrrXy07H7/BmZXCl3lU/N0qdFnzeXzZ6kzngLxuLqcS6EOQkv
3sDL5ez6dIq8TxXMoP94R+vwEGiGr/R4/xduVCNnvCoFgdJc4plaw7HEzQ1oFTtm
IbVHJzmSDl/Aa4rJh4CvBp/npLWZgAPygRVUVXPipTx/xhpZ1KyAKHsNnDp063+9
rS21jz3ZRFmkaf1Sf9SU/OgW7DP9O1GFtRegTqQr7dA+Qjmu5LfUxBIyPtYxl52/
ECdCa0QrEv0YGNzB/jzSCPKhMzMiTwQwgysX1SU+ELC0UJE1bg9XB292gYPCoX5K
W2fuoo429ypHQa9rrnflPtpZsUEe5vqRxriZ2w3Mt7Hb4kjfN7aySS4GYBiGoa10
qt5erzLpReQQjqqQ8nIqeemGpRhQTcBizTXi+JnGfhDeQ8/bi1/di9VLuMXO1rKt
cP44/0uCyCz9jGVlh5tx+KwBJ6gD9RQkop1CFW0EH9ZrCWpFGyqhFAceL++sb8Ky
T4uPyH0Flwv8nse3D/71RFqFrfZDt6Y0jVqcCyFYo5lZ5EoC7z62+QEUeegdjN3u
yo1SGBF60YKcPD2ZQ3lXY1ye9OvWq8ROZlaoeOVfUECVX4MEaRWnEvPAe25l2E4e
uR5EIyfVDqBXIO3k78vBB1UpdywI7A2cKuUcUExXb1/ihjjdR57aVq7lQUnUtt9x
x/PQVhRTSgn4Vmbbj3OzSV2K5/TzVZD7EgEOumRDGsJ8+kG2kPfbMsYwKzf4RW5V
Om99A4HvxB9hldnX2lVl296LCwDZZqi6HG84yXJma3fPDgCoOsHqII/cAZfQ0JFy
sLqUtPFXs5gUh/p3JNunuYknw5eF4lhnEzQ/UDRCe0bO691or2+XbmfOY1ollKqK
XvH+1qvu8uegt86xoFEwoF3sX+K1KH+du22SPlfo+dINyEg++Evh3h0krcoOuBwT
IAAXURWxmqYo3FHMXlOu474pSn73AcaHc86Z7nRFBqMZniY8hCG3Kkof47lsioSO
i3ncxR8+1K5YCb/K3k4/0GaKpaXc5Nvpy85HtOORkEvzdzzFOyx3uPrxhtvklbjg
jWj/Q5ehgBR3Zn87aB6yGhQMv7xfkH1pNIuDMJH1al/1hRjoA2cYzeS+hTcqEKl7
c+2YEXf4aO1CA8Zy2JnyBxBWN0UQE1OHccRDFUOwalav6vo0pdGPMaOmzxfqBonm
w5sIDZ8kfv4LMruLaVsV/wyRaIzQAC5E+FDIVgXDxdawZg1bvAPST9ciHGh2hE6K
/aP2f0pHO0eAVCc7PudwJdZ4FuDXHDeh40RttD5KMlJnx9IHwLVSV+qFuvK744SH
TQmxo/rpCk0AsstMBx+iSPY09mApwe29kgMmZgYKh1iM5k+rp59Aq/0cnpUaXGZ9
vU7I3z3cicBls1wBcnh1Ju4DzQRpi23U1y2jBHGyXC1pC2gkZrpDDH4CPcn2RUWV
Zau8Hl2ZcwlQKmyUzNiWKL9U5fRryYCsatQkix3YIVioIW33Zol25cCsFO9gK0GM
EnE8eFYdAmUYCSuqQ/gNg6UrBxvCzhwVBLoQN0qmsU8Av0U34mtkCCP9Y4EeB/Td
/cKSU5tgI7fB2y3Vrmkz+TXTOkTWhVoIWlZ/W+jq/soaB35JIjGxdDZAzim1XCxp
yWZ4bpVqyaNaRgHt74QNC72LFgwF/hMGjKmT+LUX9QHrH3KDz4aHUlN1/yAU6Tcb
IY1D89eKFFtI6GRZKkuMnZDW1aAp2dc0Kkch3fVPG71lLmyTg4dT+uFRk1T54xD6
t2+2ZiGGfZpq1HoQ8HjR3zYtO3RHX+OeCflQDMowAqKgTIiO1rBt00pLWR0X+Z9e
Qj08cy0N0PdWaTKkeh0ctWK0/sJB5kqaTuoZX0smWxHu4IQ2K2KspEZBuv2QGi3i
u90ODiJRfoUpWAudmu1wd96mp3LlB1wU/9c6Q4hYXpY0MrRQO1PgrYSEDWE8VrdT
862U7PzE9wFUR8OP9FFRyl18axQTz/Az/t3veYZAraNKEhupTttzNvXjwQChGirq
tmcYJObRsZB++8hn7NKL9+a78UmIFWY0wWmaWJmbM0sc8E/59msq12NpTwMkSbLc
3hc3cD3yzlLLa87lspjsGp/M5hcEx9oAD0wfAZYUE+D2xjfXuj9Q+CPTNsKwDgDN
TqEsUKmScWjIY4zTf3/USJLckhJHrbcbom9V2YzCxsuMjZkroqpipko+CQofq0Of
DWbOqS1DpVXa4LtuWuqzj3N88yQfO9VhruC4fJAj/Up682Kw+yFVLUUJWVHm76Ig
vs6wlasXeycSrOI1Xz8YbQHcdTLBkLuy4WOIEp6FTyPTOTLUzngmL/Z1tpmV9ZsT
qD0cS1VsUuXT7vJbkGEWOQdL6Y+CbtIMSRKlVycfLOofv4acXBr3/1mFic9jT6nJ
Ngwx0cNGu/Q99tl20O6NMv3q1dl+0THLsnWkrnzTYDNB5ej9NMv+pJjEl/8nrGfS
B9xHGyyBcE36xucX8XsGbLaSHKyTG+wz5Fmx2ZfQHNLur0oAAhFthMhhBCqN6kCM
XE14CmBwyONG6rIfdodj9+XOPMDjMJGNJy/Vnp51YKdFREqm8HuKB4ZDQbRQZWPZ
xaHN8N5WA4T0KRkLfvo6Ogdl9mAMpWdJCzSLFuSdWmapkU5kOb1za9eZPLji8UJS
2MXCKqG04/hEaq7DeuAJSuo8Pi0JT2uGVRnH6ea4gOEr+wmkBoj6ytoMpzdO3XLF
6RFren4BnHknDrDePbTANcf9lhYd9gqIXzN8uxK5rix+PcIZlhniHB0105HqEdPA
UDFKTJt2+8fs5i7GI17sHOabkndC8/4aRMYTb6OgebOFXD5b41TJgjTYSEYzEQty
LmNu0HoKStkNrt1gO4a+B8dM8QKrs/X17nIfHpQbzuNalChGikjDItqiN0m7HBl0
Z73gj7mpfMxIlRfHDcKGfslM4NBPSCol68OkBAmiS3keECxev8hWQy1incc6MSZj
Q36RhlVPx71ls+El64joGAalO9N0ANIujxMvebIqiuiNfka7HiGAvL3ZoPtzcop6
DG7U29URRKKcdUKiKFWf1Z4NHh5zq+t+meQBB4ZHgs47rB5mBfIq0x5slHH8nPVs
P+xmqWiJZ9IlDWWuanFdLQ6imAIvmHt2KBtK/rJlS7y2BCAjQhIDdqhJXk2NjuRj
xBFsC8p14yLYvoYAICCebnXcJlEeD7Sfr/qlWwTRqt71iKSU364PvrZLbDKKuQec
VUfekAlVpBKIjy8ZBpEOKtOyikhUrEON0++pOgTCyKZTQTmG15ok+bWQl1IMnkPZ
aDs9nXQyPdcrUkTJ9ZLOq7aZHPAtkPhU3ioz0UutIIc+C8N9B0LFMfPewpxjvK9K
aKQRrOxv1qi9vGLrjVGP2c0HdKKboOUaj7vbOQkvJ3hqQvPalBdgBTkx6hwxSAM7
vl4LzAdB/PA9xi2CaLO+KhXkMgBKPDPIuLa861EAwCSAGJFSHp/fuJEWl80w5/6h
2mU3JHn7uhPVyDWxtU+LcxFEZn8hrxUNKZqJ+glbWT/jbZQJwYDTbpXuLW8X3fUK
ky60V1QICkfc4UQFbG5cY5atuN05jaSLGSzcedrryLQmHAw68KlDuzaeO5S4zmQB
USk/Ir82QkuBlsuXlT4GkSc3HozXp8oKFabukZRdyRmvM7z2oLgt4aAKV+LaWX0N
am2+QxoPyD0DnqA3BvlP3zcBsAUZk4TAcv2ctQcqZTK0Swms2BqIMbgC841sZ5Dn
tHhptrJBHMpVlj8gmht71Z4ZeQlWH0GXtC99zSO9mmPXGKW+L9i7vqrBskYkF3bM
BJbFxKQUypDGJxJ9wh7unRXTXklJs93AAxOmE92kuNQ2kh3AI1pDKcSbEuple41p
PitwuHvEl5vbjFueJG6Dl/Tuz9tHfQbEBcLSfxXphPvpcK8SnF3tllMDo9SkUqRN
8h0/qmEaEHzQRYw1gxRpW0MrSsB7vMuHDN/A4nH+kOj61S1mXrgBC2vrE4cGV/tT
+6z7my6SL3u29B3RSMeEg+s+RsYGe5EWOlocW0NCC+cP2kDJiPfuzMVi3qoPSuoW
5wK/YdVETDqHfaguZAlDOr8TcdzIUFR/wJgJFoPFHu51oQJNaf3Mx/MoBvBMlBPl
oDhar8/Yg4qbiND5bO15sZS9mkBsbQQCfbU4wu58ohXlubHeetWIVbyF0B+5x78f
gjiJ7FRDHKwGakB/BQop/0qncKPP73uLKJc54d6czO113TgzpjTR2xQ/TJZx7MeC
vTD1tp8qL1QyeZNt53fAtGAQgtmF2Nx40bHoI5g40Pa3xA7SQMe+5RwbE7rOWcKN
u3SzcfZZsf+TfMZoKHb6kt9YQvkAdX9xZCdcvuMTLJoI2HMVgKamyhdyaBqiSeM6
BjJ5BoGB2ule70x7QZRaqP8MsUipR0WOfYB+m/OAzFsRRagsiGidd+Go1OiKe1j5
d6nhcil7i3SSEtkfGP1QgT3xesFBIfo0bwl/yPKioEeoCviBl7DXytOpDwe5zxaY
yLFOjakUMIJxdPZ1Xy2fPoIkVGXErDi5A+zWKwvLQifvKcw3DlVzGeuVTnFRNkmx
V01ulsdm9E4O6XsrmA/BspHwg2s89q6ilBDSRqYccEfE8fO+9I4qK9W8c2NElj6z
VImcQk/V5JLVPCBUX55f/DTqnHozUS8T7DB3hXlApMj06U9iPQCJLfVEXj50n9bB
qzRt5hqKjxxk38YvedETwYxhQ8D5smULayfpbQCsSUFMcM7cpbqD4vP6tZF5KE5K
nCgCQuzsyCAJvvvrpFWh7mMZ63iMJQ5hyDAlVbgj08kTk54nIfptWSE5oNQzbi7g
E6h7xt4hdft01f038tLyIXXZ/jE8cBXv9R5EOGUc/ju6mT91c0FF2XSrtAYmKFEn
arxH8zmtc72RxmYfw4jUTtCnUwQASMPrzcn8nB6jB3+0aKhlWqwy92URBqBNaxDD
2QLvEl2MCruE+Odv53rfucjePv+ALgU186plOJUm5irl5F80Z7YXo2SOvH6P5fFn
AZRPpqArwcM3Tyx2o74rUoJxeiVLXPGpMGkLjc7RX/OrNhXaGONJq5tCanHUtHbG
Ynt3Gv/aeZPsrxxzWvFZk9/fsnSz23rt44SmXUSTdc//y4tFZhznLGOrdx+8305Y
j/KfWNJaNtYNYdvvMnYnL7Jy5fbQkWQjusMRoVVEArCHDkxr/s7G7Bp/dymB7UjS
pEHSnukf3uhsO7XJuTAdC/WXWvUloSnLj0YD8szzxXJyC2JluneOLx6Us+F1A8S3
fpQYFK/19O9FhVKVS45EZ3tnWNWxyCu0FNe+Pt5mhDmLzUIfpQokldCB6liBwW5C
P0XhoqnhZenjMRSwJO1N+zA4W9XNQKI7az0z+M6qW+6OwMnGCXTkXfPSlvX3AN55
XXsnWCtUQ/+UwHTh0qWV7rl10jcrxx0JvR0vcLvEqhtJooYoA+0V51OxJr540ow+
GDazvlsngoNWKOsW5n8D3EaKodtVHSbhgRrPGyF5JEMIyo55jYN6bwk6XJI4Kwhg
Fq9Di3oGw02+c5RTgeW0DuWSUORso/g7w0aRSfSnW7HE7JL2LMVYUuctvY+wgUbD
tm7DfcdkiyclokoG4BT24dsoIPVytpMe5OQhHCY2i4LHZrBzUzBSx9I2IGi3G6+F
D3amRPH7XiZQJ3njPSuXn7ddcrB8tNQsMjPLUBYAF4NJ/vb41tJm6PkZmcK1xkZl
47xwm0hfp462y5OVyOPGbgMWOhIqLICdewoa7s8HRJuFYaJKQOFp+i0MkTrgRwfX
VVD04e+26bMvAGy5f29fFrfQiKKSqMXA8qviywGguhmR56n+X4YHahQVXSEGC83i
AUnZI4KLJ8x6Hq0Vp7unfQF7d0gIcwcAQ/ixlNo0ZSDr3xFH8eRpAIoezr68M8hB
08IWI8LARy9eut3KCyTp+mXR5ynPKijj8Kdq4+3TVTG/PxZWv9kCKSaELDb7BvRh
JmdQet7wIBuFw6sq34Ssle4CbShQQSp0NVLmMYaLi00/ECdr3TRUaDmgNHcEzLD3
5V2ylFEj5zVTSSXLgewa8pXIskgWqpnEOMDcSnDKInPieCo7Gqeog0nb9WDxUhec
RS6BbfEa1ow7+cQg6NzATe+TgAvwcSdhbjKm5sTV6tsvyazbpGiB4HBZqBaNtJE6
yH0j9ziIkYrKYHsLOm9UN0HmdRivnW0rC4yn8zIuWryyyQGdPniKey8DXPjroukj
6NtXsqmUlRdsCFRdkMxvbR/xFeMLwaCtQy/bHsmxMkjJftjJ/jrvvgmYkAw+0x/E
5TPV+m3gUQ3FF90IJSwndTOZnIh9+oSMRxVzlaii5hyetahD8Ld1KbJWfB4Hvvdg
oi8hbewDb5MzelMRViEJIlCXDmx2Fy84upwBLHXO5A37Tk7tO4qiyL9CaXFx+jt7
pxvznx9aDNzmsWPtq+AfVWbHk6Crupgw8bOTzM4omtJ+b7bjKCyHcKX8XrJdRlKQ
GRm+kKqoxqkzn72I1IzcQAvQZzfN2+9xBmsEggaqADabD3/+7I/JfvV0ATnlenCn
/l+qrFvORx1qpTokeiI9p8hvNWBgMfhsabWf1kpGd1rioLrEYZJTkcnBRw98RHbl
dlf7tew4t8c+LvdRJXwgPsV1nm2guDqCKrnzAfC8KMCy7DyFcV3vzXn/fmUei2yE
mcW/H/vPhzKsVYNzTVLp/WFpcyBI1aziVBBZEflpN1JGhnhIYPnCQCfe4A5jMEO6
hYQ4EXs31pxaASVO32QJd+PE7+E68l9cynlQ4fJo6p69qLSA2gATH5XRnOwFUYiO
HUC92EFd2T2l+HG15NjyepUV0k1Yuv2+GMXPHp4iWJWuRnJNEOMP1n+y3gZliykL
dW5Ae26yzuMeetqE1871AyD0mpqHlSmFa6ZCuXrf23YeS0LOKUoGlY6WUrEjSMfA
uLXqo2S2sNnas87kravOJTerG6+4qpO7VXnp0RPy9KVGpWiD+ikCh2oTtbZkAUI4
2PXXkFA1L4VLjbld7joCzJlh/XRp6SMopZAicb1Qr+kFirDt+/9jnXXW+1mLxdUw
nqWw+wVLZw0LUw9ULz+hdksQkgAem0tBz2agXEaMMY+EWuGlf57C5PKABfNrWh0j
pGeN3e5PhAHrwxe4SbYasGkggKOa1I57rjNCX+S/yxZwTpxi0jer8cyrnMXr+3ey
uVYZO3nXjDxLBz01onDFNojBl1Rd0nA6n2X8b4KhIIr2/ijuvEpETd+VKfenKRtU
801rkoAWcWzh1pdg2Zovzm4QrGGYRU3aXKC8mJtlRsFAoZjx2C6Qy+VWyuoYuGx2
WW6Xd8EUGgo3Ngh+gRrAk5fXEfxyo1/2t6LjC7ZKGQ9d8U4aP5AjMi1n8hd9qsT/
FeHRxisJL8G8b0IUUkGpR9pC3D6qLuzBlZK5JGD5Wp5iVct3iMTbIliMFi+dwBq3
EfICTFa4BUNzW/tnSI7XueK1hPrGAseXUU0g7JyYroXovt7YbXfP+pRSXj1gcU1m
h/k+XHdoENIuQ/ZU8QriErdzZqmV0ic9JgEeK+kdtoMKZfszS59+k3gamgxzBF3G
F5fX/Vqv+ju1DoxEJCXowEKqu+DQ5X+ulS++MjocyIrrqmTKTP5tWPLumEdIRh9x
6JNbdzuD8e0KVHNXfZzIeOYyAE49fdzP3tU0rRxKJOD6Sx8nDJ8MnC2k30ChXXaj
9X8WZxaMvp1SGx3C2c+j1rz5VtRVfY59O6PJRqkve1SkILPTOmNsjPOxuK5tOBV2
RouiDogElNcZz97aiYsYVBNuupXfX9lopxNRVYsQR4L5VrfB+8yjQX8029AhwMYx
j4r8w2Yvp4Ea4TcBuxllODA30oBXIkDh3yhTviNw013MeAnTX18DGi+9V3IJUfRH
OuV1jyYstsFocFbZe7kz8Rqf4BrblukGcvZSIt5Sf1Z2uRI05xLYRhikjH8QKwZv
A0Zey44K+NPJ+PFbqf8UPZPzU/gP1i3G1vewGfRJZybpICWqw6+f76Ete+dA2Kpr
ryb0+gYfcFMA+CLC8kkbvLwh7ReDUCLZM4WPRzBZiuE65CEG/w5QbQDU/SJH945P
n/4UMnp08mq4Ru9zKIqIM4bp/N+QAwOsF87c747KZG8mtKhNbaM9az3pGinV+ONy
tJcizR+5cqmbZ8dLlHwNpF6JyOw9xkHUYfZB7Niw1/uS3Nsuco3NIclUU3kzLIOW
425C/C/R6nN9joDdBBlAn8Ib8+jTJMncBtHIhTMfnqVdrafgsXhv/lXrqNvEwvJI
wIRwRtCzP7gSHYgGfsy7l9JaEt156bDzmIrAHwYEepXh8n6KInQ+nXoUoRqgdgDB
VtRiNUTHLjqYjt9I3PMwYwukrjyvWDOQnMNosSzihtEMv6+sRA1vstHcUCMnUFd2
0QstjCUl6v+yH0xfitNnWriWmnFH9vXwYlXmdTJB7d+N2+BFJajrN1LfceQd8cc1
hAyGnCOK8su/yh2kQvNgV23FuIvUDqL8dcacY1hlLv1kKJ8ygD6lXv2LHXxTVIe4
rOd+YgcKkQW2i5OA6bda6NVmvyS3VEUXVKzIvb8c17xW1CHAdbpglrrcvucfcd/+
yQAXVAfEeL721vB1/dM7DwaUC6P9s4pYpy822x9ZascaID5KbsPJ+cC1ew7jNRYZ
/QbqDPgcLTlvXc+mY5meW/wc62ImXuHlZ9HOmAzZKq1w27X+dw2fJWUM5lehgxeB
Nbv5kBYLurgWRiKvuLeksHYKg/dtIfFK+wr4Zql5/fcJadQdd3NcDzFUBQNbuxgd
bkxJdXEzdQABPIuQSodwqbVbyrxSNRNsXdvFldj2KQ62xYZdCnCX/TxkN2xnoXao
C7mYKfCNqw9UsgMvD+yOn/StpP1eizon/PhjigaaTTcjxvkGKqy6y6g/AW77/vSD
VmJ8hi6PEDfEuz7i8HlwqPPs6/S7xTaORxkwF5b10rERpwGlcDH3BFpke783qhSi
m88KwR/zYKSP+yg9WXwolXtw1oBz+uGhK4g+eK4L9FURnymHHcgukWzLT4mSBYcP
mbGkNk2ZbDdrPMzXG6Es6blKL9M60cxutNfHmB1XamDLcPRi8MllgGeP3Gvuqy1E
RlybMqt4XN1uur6CieKIZXbwEJIUkS89g2/aRKXCdZ2D0hmXjwu/GFWjjKH+Rkdn
BVb+OQjSOeExn3VYKlFDsCBsLIqBrME3ALq8yxdbZDiWWFRFeC76jCpNfUV4oLTs
82LFoMP1H4aVl3skHkBUaOIXuTjipIVzn0o7NL++HlpBHr+tOaPZmYguFTbRJM1Z
PjAb3vpcsYDWttzu68JH0yNrEtkZ7ryFVPkSN+N32hsh/ltCFi2T2GB82eZScvzG
WcDwCZ/Xjk7kFhZalYJv1i6NRA44mUz4GMOo/EE5KFdWMkgsAhMbhN0ouKgtW9SJ
HjlRZb9eaRftmRUjQUxh2l1gC+RBhWTKg1Q8hRtH1rPDCFca4xKEsF8n7OHMUptB
WRHsYKnim8QXf6umPTn2bPuGH4Zd/GIiR0+dLZu+9dBA24m5HvDCHygVmRrG9oNq
9KYdOEjN3lTDp5KX+ToFtzlflWIermijuCbMB5eXFcgoB8NW+ZcXfZjHCKRRcsir
9K34xynZOD6PFMqIj695FiNTaKiw5+b0xVRTfPnBdqtoIaq/aQcEnsCTp1IeB6Ib
0Aj99tAB+Ii/eZSBdORNTAB4Swj+5fFsSiovpAT58m/o3DvALATxpmraGOYnGPHA
MFmRmV0OJjIb5YpxqLuxMriguwEPskoYKytPWxJZA43DCfjPvia1pY3MLG+KPTEk
jO4cmBN3VvYcEEeCbqmt0V3K7e8miuaTYm8WlGlh5+shjIEisw+LtFvTHwyMkzUS
Pl15ccWnsfhZia15jUbEM0hH0NxedV3QMbCD+SjILWcd43k2vgr2/Mhib9OuAZiE
4fWIQEu+WmYPA5D8GezP7o0DhlA2deywZFO6+Z0Cc3UuQ+ZKLbs6KQiFmmKTuBcK
4KntrpYXuIlHA0SJLRGmFz4AC7Gh5dFhhuTu4CikLweBadNJM+7U6GA/VmidDSBe
zcg7856n50TctLLIr7e9WtWPXSNv9OeiHQFqzC5zyR2shaCFuevoKO1Mkf9U9V6h
I+UlrFZh/1Yq41scG0JioJ3BcBuY8VyCvpxmG0hCgxu5KIJeJ7G4lQC5HKvrEpk6
Xiw7PuBuOpP9bZpCl/wIDah7baK+l4e0s9/6jtCKWju0CIfyS1+B7+2hq1CP11Qu
dIIF28Mb4L8gsAkrYEAH7wDLhGf/PFai9tHswvygJI77qzcFftwbQQn/QpCkCIkV
wMaLxHBzXC9JOBO/frI8a9frk3m3XMUZbprs2gxduTZB8p8b8qYUScgR/vblokn3
lRaxaUqqkt4WzaAE6UaBeFGFj+VQXESUxiK4IA9yg3gemI5pWRtZsauSHhSoyecG
LX/qOlqAZQnCiNuLbLG460Doiaolowg+LTAQZTBJIiEEsLX4iWCIWF7kavYMpHz0
rwiSxNTX+FJhqtkKfw6WJ0jWtwdfkZPg3h7aAyp0rEAdIgTmeX9se6kmzY+a0ad2
R9vuYsjDgTiRaPpt0nuG1575JHVRct/3Jxqs9/xiSA6ei5PsWeyporFuNkSnphrR
r2FGInwgPCnp/kiyLa66MAs/xyuNldLA4KV7r6XOEkltWxKcz8P51KR/hVWmRxWW
0xm4GJAAaVIXwmN0xl8RHuLhacw2/1yoJs95LLzRUvoxa6/zIIF+s7iEHTs5/MQu
ts+6iteZ+z9/RkIkgcGIfEI6Gm8GcUiBbbWDorhVmF1O1RFtbHsmh1f00XVPHoyY
ilKtPvrEBDPrJkpaRJl7nNXvnoRsuJKEI1OGHOh1vPhbRlD+P8lFe2oHFaqrCx+T
idKdbx8LmNo/gGU7s1Rsb4nMe3GSk7C26UOiG3qqOyGiAGghWeWlXBDtnb/fS0mt
t94chMiVXVM899VVTXXFxLbaUrBIRlzpasCK3g0gFtDlNxaAUcvs2Yj6mcPnRe9E
IOW3Z0/dSkWeIuZ3w7HgOt4cS4Z0GwOcdIEurw1eyNP+hogwvlpw9HmzsGF4PgNV
2hJ+UQTJQfEtvOE002EiGtEUjwko8FWS+L1uMiJU+ks/tC85btbaQdh7p+8OyyY5
uGn2cOyPvGFcUN4q/TmrDyL2uPHJTmQfnmw1auoezvKLzLREMEYA3Qk8VU6itXyV
hPfIfRB93zamZWFgIyAkN9GmQtmEGXpgTWZ69C6c7Xi8rOk7X1jhwh+ocFYkD49e
4KKBKY8McuemI01Fb8CCZqKEJeIlwCN63Bynd3ysx+XmS15CT5d/crfmv5hgI09Q
6cx4tAdZEGpDh+dkSIdswRsQk94EBFeiKCbGhTH77gcraVywolgGVdiZcTGxAdmM
TsuriWaVycF8p8eTtFoMD0b1MJucDJEDLN5Eu3diV6MNzLl0P9IZrXVjIR+YOgtS
ML1l/ZMB4jJG4/LugU0Sp52GBMStyyhYv+3wxIKVGo35p99SI2nAsGjAQz6CFWCF
VHxwfqDhFOH7rzBnnhbvuwgG0R7dnXcmZeONqcCkpWjcqzX8jnWlMwBDX1DBIVjH
xZouWOGY+ffm5GVArUkFWbszzFT6FPml9h8WOhUffI+rNAUzbjMBRqP7ZBmEkWFy
ZEdGlCwbeCwaC3ZVV1U1HYHCOZajYfttOZLCySUGcew9fSno/bpMUSrJz4xisA+2
ZXqyAoQMQQLaHtvIjAPVBmbPMo/JcDmqbd6G7BX2RxICmMZ/FFUD1EdiFPeID2J7
l5ThLhpzZ0/37mJ5RnLYeVc8O0gEMWWds36gIfU6h7iiQSr+PQSSuhrnowtdLRmm
or0oPKhz1vEMtQEBUrBXLbWU5NGCJDqWb5l7cQTPwmuOkUA6RaHhlM2iunHoLoA6
2VISc0fQRqvd6j6Uyh8czBTkS30KYOo0MfdWWBzou2kEHkD8aagCdTLyTbtGkhfL
GLAnGcxyWNj7BD4WVeoTJOjnu/d8DH8uCRLB3/GEs8pAl0SsJb+vIo8UjURG/Lf8
7Zh6/bT3uUrzb4z/sXCGgT1g0q7gjErjtBXn8EYwU1E44An1m/h7dyQzIgUJqDmi
yVnzzpJwVfdmGE8flC9xtvti8YPnLCAnxSoCEAUEFuqR6/XMtHM6vrAu/MZNUX9G
wxXnaq/4VSQ8IWrqJZQLqssTZudkXU9dUrlNjRLhBgMfbYRaIyFuTD/JedM3xPBx
QMBmbv9GgbLYaHwxPcAiTJl6srqA6xbE+iD0k87kiTdeN/BXrAcN5KvDwl2FKG06
fvkzOsXvqkYGe+61xA1h37To/rpnWxMnagH/zeBS4QR/U9ZOwW5c2ZysBGmqpTV1
3ViXpAbY0/2i/czXrDsnpH2pd5lENZmlqZ7GzUDy8w+rwXL2QfYwT+GUKdnjbspy
PE8LN034R4yDX2qCggZHACRKEHQvOkbU+ef7A5d5y+fYRzlts66SZWXu9phRaim7
DRRvEKFH1pLWW4T0c7Rz8d70TaHSZ3xAr212GCRv0o6EWkcNY/44CoJmfnOhGnBh
NjfT6RKdCW/uanrSN2mzjmoMkskNudeDrWdZAkG/l/HS+GLx0a4+7XvAY/s0rjiU
NvF5J4uwSiIiSAQFSHzv9XXSumwEw+8lkzbU459/kKUMsrqNtUyPf7K4qZ0LDEdr
4ds95JRJlS2B66e6tn0r3Qw05aeuloE4HYwutR4fgN4WSkkaE5/+wpp4IpdjSaUr
d2y69Smmm+1ptaHzE1mJPVWDBL21mAdquZ6LHPnfWND9WUR98pnFWP6Zhitlh8uq
+3VH+/ymzooczKvhD4Q6gJj0iK7XjgWp6etLRGM7N2gJSf6/TZ4CgyOtmu1pHcLc
NVkPFBEzg7AOcXGiZqAfrIII0uqAbvaVV+NXCuvdQCE25WLKWoB57M4jG+xVZ7t2
lpxqnf0CyHGWDAdItoYF6B5OBhbbi5hwGT7gkgRppntiQgrgvqyeB8hvhIGS9XbK
TT2o0H2RTYoWIrQPUCB2dHxiPNixUOdBlezjQALEDW0y4wmlbaodZCNuQKXqMrD4
NZ0MbvkQuRX30lN1jkqPuOY+cj5z/CUm9G5QuwtJntAwSk4EuzbxzTbMyS5CVf2h
QEEWDo7b2pjnDfO0UFEwO23Yb+u2idHPZ4gddZOb2VtGv/rI410yvDjmbv1XyYS9
CUsDC0N7XvuUdOMIO8BGoSZ4fud5yEPmKgTY0b/HcXQbxnEbupPXrIJ7VH2BKlBF
nDnQ3RzOLSiinGVYHr2ryYBAV8P5oMRc8f1Nej92GCVBOqEumhY7JdYxj2cZxphd
6gb0n1NNz65yqeWgSy/IwkhA6EXJ4luQJFFx3EFcW+y3QC0Vij2gp2Pge2YNXN3S
4kZAQndmnOszeV3NmVM5KoSv2fRC57TpX1VoJV7f0sar+XZOv8GD6vmFxxdA/dvh
PjXrWZkUeM6IVrjp6NklBuzqvrvw/BiUuFcspR8Qdb5/N2jTm4AAP0sjN6Gu8nkZ
8N5Zpczv3NAA/KGP4LtoQ0m9xkoh7EDL6zgI3ftC4pKIrGQUGsDxZtw/7ygpUMjS
JGW2H80wFe8tQU2BYPrTSRp3mem4ww5MZl5iY7kWL/YFX2pu1gBw115g8GkR/+3x
pElU7qQKwQN2VoL8AL+RJ/QUzZcKr3o+U6h7ZyaZlWJpU22ehhVaLotPzZ8RpYBh
QHFUqoVZnOJlr+s5iZ4NHRoF3Ap1bfZdAU40hz52GBwrjpNvFEzgmi1H1/GQ0YWy
7IUZprSCdw8s8zwlOkYtMj0vDSrZ65fi6mk8qxG3NjrKNJsiDnoYSc7T2lazGYd+
SiI2nFm7qV0qPfBRYDJ/VIjPJ+e8+07JWDJcTeWFASJn4cUhkkonJtCsl1Yr+VCL
FUh0oq9oCD1qSX/CkTpEuAvO4PrTCN/igHTyOiW5DZ6gkgC2kZuLc1aAjXNdnz0G
4vTfscFzoYP5+qnPjY+Bq+CZtE21jMpQybp9xu34J6or2TXyNJqe6+1DM5kC+7k8
5Hs7cSnSj0jswdw8ipyJVkmqydw/YwDA9jwHPEWu5BTutgNIftb5VqgUzf3PniIQ
juLkbaYQYik4aksu5sKycoeXNA2616mkvXyRllnagFW11OUNVeNrfUHuQ1ciA2HT
rPkMIa4zywySK039sMSZz/BRARs8q+s7vRRnGZ9ylObbg90QZwq1czxeBW4s7Rsx
VquzJSDRTY4NYjFpUTMtQQVdzTWiz8PjcpIcMMR+FFIwAgbOXtrVB062r6DfZ2L2
wqJRma5cGkvcoKygY8POpbEaYECYSZokUaeZiRvr/4Dg5yvwWpI4ZyCkK/NSrilx
5NDW6k5cxj7vQnUxVSl0xuhzTRZpw3MjutaE3+cfVZJTv7rHPJGfwxXczz/IRByl
xBXBH7qAAab8/I2wCzS6MKBfBKCiXTHiXzijM6Ij9LYHbYKgcaHQt2vq9kY96h5D
Ed1ENSMFcOX0ZXTTaQroFG1THe+b85msZASLFgq9cqSuqZLa6XcPTlabEjC+39XK
K82qJPrHami6tdrMJp1rXWfiV78Ay5xHVoEAwe0g4biZh2XNSapNw6p4AnBKy+oR
+KJiG8ZoGHNY8aJvs2S9Ye4lPf3p+uamX/vuaybi+lMYeB+5ablUoeT4t6+ySrUB
KB1fTbqzPIfVdWL9fXSt19OzJo7RVSzMWBpJnWlxRQvhT7pNd0CtIkmVyL31HPx0
gOu3BAZ4bcEc27XgFVGlyAfjXV3ca9rxV2hvrV1mfRLXLU0dv1ZDnd6PolK6rVWJ
gy/HEpcUckbkIxw03KHOr7qo5d//FHBM6Mf+ZaQelaWYLwwxVZzNYrWkV02GaOi5
gqUjPglg3Ll7R9E4CgVKOEo/cvBV3lmcw1nwOpa0w1lPkCg+71d6JfZEyCabxQpO
UyHvGm3D/Rg3snFwC4dByKJXw5rK1kSfKfm4df+KkQo7CjOChn+Ar6CnhE2lO2cI
zT8UUVgkxBBnqLk62KnSSb3FxeltsUuFrxQbKvv7sRMfnvTpcBVca8TO/p7xhc5O
O+0lhGP0V55q9d2a4Izhci9MCWZBj7QI/HZGjDbhhPKjUF+jwm31SDstYHZCo1Jr
XGIRURaw1Or2pFDHIyCkiD9vLjr74gYzqPBWi3v2ol3neTjt7A3An0YRLDoYgqhC
lRl+YQz6+7H8MzmdhCOzCZr6RUSqJK/wVbowHhvjyZDEi0bk0I72ba0nHlZfWOJ5
/zLs/iNJSi6WnCBIzSLrEOhJXjnV1tcdca3EktP/DV1BH1WrwVWzqD+ue6ChRyOb
M8CsCO7Tr0VqA+aMGQ/fBzJN00m8J+luKVP+JRdEz4LRzrF0b8VE77AKQ9K2tzsJ
hujF1l9/9aAjV/pCy/rpsVe0IGHxLiheuWrzvFaDrznc7pbnL2Onu9nJ1qG1Uip1
WmK4mkA7WXDDgkinfXiznygx50jTJbfIDWm4zj/qZUcr5wiVfG9somz4HBzfHnL3
keJ8fgwJJxU/hrgZelLDr8rkJQSxjA2t38D9OdmblI2sKK7jXcRE2l3kwp2AKL9n
mLJ7+Rl4Njk7ghgeszrKa7YofVcQWwyiXj42rfRj68hj37wOApXW6ZYoq60XhqBQ
cP2EWxNyQxWd0ThF0XZ/z5UUi0Ymii9ZS4KdmWYog2pCEYIj79jFxqj/JNLOtO0B
GXsuU52CCjRZ8NK1QchFKdOvi7Qr97emzsB9kTf1SZ8HobbTnBEhp+PkO1Mxv6OB
ZZLAHca0xCu29mJVVN91Wv4JTAsISAcrh1RBPdyayOnHD3+zflscuvUOplpdHECB
AAHxKvVmk/avLYu2Zs92w3vYG1FpnNLhSur8YauasUyAmNun/vfLHyQH/6e58mis
R429v7TiZuHOH8A2BsUwKJGJGMSlaal9Uo6vIVw140ojP+LKpeI3sVGeq3dDmX+H
L9um/PoXB2l6NPThjmnStQzwkJuEAgRlTU7oD7NVIhhA0vFtX+xzb4nIgkwhHN3o
2BGOe2/XsPNQ1ILoCRPYcdQbyPokQgGJrjK5NXy0B8Sk7RVQFwxlMniqF9CB6JRx
eFQ8sZncUhXBQAjyburW4P6lGtpO67B8xEy6hjThaznMoTQRPBwwAFKBdlN50obO
4HSNZuLKOJknrFh+e1SLvTUZyeoz/osTfeJ3baUC4xs5MI6XICUj9jzckPQuPvnO
G/084PZouRtk3VZhyfUEqRh9Ru3or8kmaQjdsaBN0ENeXWUSTxRT7mosSsB8pREt
W9SNPCsCMNSHNRE1AfhNEb2q2ssjT/LWVuIwoBY347yUiQPQw/pTFJknd1qQcvoN
CqSO/LUpQLa6kjHD82+THU5LoR82W2OWIADuKI7ew7yYnhQCDbnFx3YXpntezKMp
XZbVePvnxUr9J0x0oXPQ+Xqqwe2tzfkR6jurDwrFehu0CPWL7mvHeDgg88NPdC94
nWPBIZUQaAuqMj1SVGC6dL7yE9a7pHdVWVy2IsNdhaM7V9jYA3Q6rgFC18+QZYL8
+5ClSNHilfOcFlLfcJ4f8fUSsAZrbtvMAHsyz7eNlHJUVRQHNLoeChlloUzp5DUl
qvXOJdeRnTKHhms5sWwjZJBt+PUUSdIkGf3Ws80OeQ/VrRYiCvcOcLsuHwtjSc7T
T/cIqQOZLVl2bCGk2W6OxGCgdtzirKZ+uoaHwpRGYU0NUtq8nvg6PeFudK4evGkH
ZJfjwOLLyeNK+ynyTjlJZ/5zwe+mV58KPUk2RXorB6b9UvsubVbfulooJU2KBNl4
ldTHVi3aCaacXEZ9fw4l92Q4JlDgc/sLihohaAvMXf6zoO2isPhMWh8OOHgIC9y7
vigXandGNboz0B4Ymm0F7WA9+QhrnonJfyMHxU9NpGnrebiJ68m0kIgZO0zeZOuB
ln8hlY+i3kRnzq+cJIzZJ9oJEtyJHqe8dANbSpOjlRBITJHB8WRIcEJCXvbMMD9g
fH8Gj6lzdb2vAaib3FbObpqLNKqZASjHpGAVqA5lv6e/9GYueyVDC6JXjiU6OTKF
dp5izsczbmgmAJJUaXml3sCqRmI3LxWaXSN9tNzw6j4uw2Xx63/GQLy12h2RYUIO
7OzjB7ff0SRDcQhYT1fFr73j6jzb+7LhpTSmMlH2Z5CjoKu1+Vjz68NNB65a+O0K
a1Td7nVJzsMVkMNzbtKTfOBHgZ6TIbiA+B5mUCOZvPf62odaC5aIK93y9Qbn23LJ
EugktTkseLMHVPg1nI0IHYdJWJI3p+F1PIJmN4Sxko2StIUwWLEWSs72l9w/1I9D
ufxQCAPEfwMcDb9Nr7XcLYG2n97gmPNbNL26RodzZ/j7PSoE/FT5X0Knw4hKXxHa
GKDIQOHLpRSohvhra1Lj51FTKAXdIpTobDJpJWw0GmeT/EFu1le4CY1TSl1WiksA
BZeprNkvqbs/GRBMr8DNXvehS3uF/8HJMb0z1pPf2UhJWuDTgEO0/OYTFmQSm6B0
uUwEQvxqPx7rmuBnxup6OijZ4VZEFyfSThMhmEX4Zpo11dBOGU8GuHTI6Vi+j6CC
umH23W+kPnGI0DhQbowxXpGLcibfyJsV7/uddxRE5alr6H2hmU3L4YBRE9WnHby+
Pp9fcoTTq5Inq96Ur36pU60+t+YJGLiV1I1cYYJwQc4T639AmjkC0jeYPMkNB/eI
E1IBTX7WplP2+ekzzXxYqi92UwrJchRRPF8AnHgT6w8pwuWT1BLatbxpekt2sLBY
PW0vIYuGauK5sNheDP+vNa1HLrj+5KDdIsGVhMEUZQzP4KqKQ+yNrWerP0mCaTXo
gZru4k07B0fZk8Eepnn97RG7Cne/zIS/WoYizqzK1V0dcZS0Ksw770sBSVI9k/gL
2+GedC4E6vW1456+Ytal1dheQdiZ+MasujF6XCsGywunvq+R8iWkNtCD2jNeXvQd
KdiElaD7ItwgI0eBPBLJ/ttnQS6dCMaXATjPFlF9uXRbnnYPNHxn38ZijBB6Jf0y
A3eOeQ5zvVWtFdjGoIzgC5kwjReJjcZJL2WO4xSX+LM0ZhO6/sCV3vBd14omBpjt
tHoarPuJZM+z0IHiyieb8tmVtJSU2rkrEyY+u6dyYyRAZs5CuZ3XGAHbyPerEqdl
a83+y3pZcbzOYYUp1akNiCkY8+NRO4DPQ4up6ci/UUfxAb4zYvSX+xojSjOdTzfg
uugGp8zply39nwte9mpR7107VkphBoL8ae3eDnCaZ6gK1f/SdfcbpA0ogAH3M5Qg
PuvcrHfBcprnOM7VlTr/1lE7HSaUUDl9XZu3pWpKRDwdYIPBAjDxnuAFZdbWi+Wc
kavTNyXoxAYSPKBFqH+FE2QLK+yPwo1POUsF94G7QGzDhYcRQ1oHyFehQ4RJPbQN
wJcMJptgiUfKzKfKA6kJcF2hM9im4v+9CQjLGNfFAJrhRCy6ixjQlGfl8GrWLend
g2ipLce6+aoFwa7RJPf4G9iEO/0wrzGY1ZmyRWMsiqoy5G2GRs7DXr4EZEiZ4W+/
/OdV4b9jB3/Tl2v3oZGuyeDHOKTVijIoMGSpAk/ZXNnrGDABg3Z0pQw1DLk8ROEI
BPfq9LBRmoobZ+W7n3ZPVbOewCRh6xtm2eem+0z9UzURXzLxTQxBpE6uAYIiwmvO
GD5Lv/s4L8l87A4oGSjFVAunWzP73/ZaB+EAJkodCLrss/ooVNNpuFM8ohkmvNWz
M+EEcbmDa7qHPEKJAcVrjoaGwpjW8ZWkOrWEJ+4fbJbv205IDBlGj8brD2SbJK8M
+MSktVrWR/+uZRtT+CLzHOJi1q7uRU+ESnDj2KiCcE+mI81mYB98lkyBK78XPY7n
XiLXj+Zu+OOJd9kxwcnixx9SanQMh1Xw4UooOzB7aE7r4x98d1WLRU0M+MBJVRwY
wKMiubjIlKbjUyfh2m8bAR49HxeMQg3MiNuAtTAygcdLR0tWylRXHMTiPeUnxhgS
RA6qmVv/DF3sM2f0GpTpcXBozgVZSMrOePKbfrt/VX+AMSmJUy41/l532L/bKoql
ftrULF+f5g2EqNtidwE0enJtvlhUZqFb2BSF0juLETtVDCkXEGzNLA7NmpDfBhlf
fihUU22SCt1VKuQldY5D0TJreju535EeWe0JCQGTDwtL//4O5f631H/yQqjaFbXx
/gaOCQ2y0+uLM1y29m9HgDvX+aaUegkLhS7zmdzH7HejxDwgdA+QQW1ONQcEFwmn
oFTdNRghBWWZCRjxYcbxcQmKKQYOcgAJ6QByGIKNMwBp1kgWesyu1B+b2HFbAcEM
m8emQDtk+3eLOjR0EUu6iYpC0eVn/kd52h0s/z3lxMYN4n+OaEOqJWyRXgPp48f6
l/7ivtHDXizBnSQvuvbjE2yQWsRWQOgLCmEHGz0rfyvIXnVIJyFkVJnfhTd9rwj0
Qn3Wezj5ihUiBI1bHocRq3yLxUkNvT8NHAcwnNeQinFoN9g03d29KcszfZDXn/PC
SZPeNUczoOtwLtEZ6dVEclhr9c0qERtUIWpaeyN4w+yHoAvC+ZHSBYC0ct0HUaPK
yXvnRer4bgUSWWW2PdaPlS7fj6icBK4B7YhetTegeXx8jXj5UCarag351+nzDLyY
MBib3uRJMA2seSn5ty2gONdArjFVeXoyqRMhqY1P+n2wBZhG2pXRrKDfxCImsGA7
2eSFAswlxgc8FJabsPQXLbPSnKjUF8ROwVvrO4B4jbNP0oDaeq1qM99/AXt7b3WE
K4cKWD5iwOmab2m4iXvjqzL6+AQz7AjtjrejmEtPoJmzwN4+nBjqXvQMWVTVRown
IklYD2rpDYXz7jTeW7u0Xger3JaX2Jhzhx1iI7ZHdei3vPzCh65/KvHltPBpjSP9
z06hh3ffAN1xwKgQ2CEFAD79lX2tNTT/zrhczubJj68XLoOeRPWdHAJbbFhRaP35
uYccu9ENZiG5wKgDZ4Vx6oFjnc4wqMPF5E7E7DvfUvdg3M5iGgoYqrfh9Qap1T4v
UzrkNPV84yJYWluV7LfmMQvqT/7u6MaUApHYOvTeczIiHeLKJG/99QFEV+Cn8MrA
hHPWJ2kSxbJ9i8sYxJqUY0DHLJbGTTi7+xcFxm2Peo3/tBGKUs58PQP+aJ1Vr6cr
u/oYI4Xm6+Lqtx6a7f6EblA3n8XNmgSlY4l3IGuTNRCAdO+YNv0dGeAQ4K7yLTOc
/yx2FBVit734EgaxYKB+WyNsnPnZeVxaVwUXjgUIy+kiVp2mGAjesBtfQwh3W/z3
aSI5HCRF/j3WSSkZeucQGfzgcN7fhXA3iSIyzZ9SiW8PJNkCsk6XtpB15uYUJ2mH
7+Hf9SxtdSNH+PEXjIR7BuGpHwJ+0c8aLnNtqeDQJb+9XzRSeCOKwqQT8JIrQ9/S
DRZGecq/G1Ed/qnX8T2Tt54ZDa5Ld7KQkNcCgSf9i6HHwekIAvAllrBC9wXSd2Eo
rpUfpZKYxOkc6saMq3eH9kxV4LPSy+RGFQhrWQoUawKnO61abFxKqrQ6oRKFh9xO
tsXZki+r9eQHRtD/z98uVTs1zDG9W4tnovVd/SVDHSlP3502fUQ6EO2BoEVDCSi9
LhdjjQk3KZ1aPKZDInNnDAkDOgROxNuG+pSziOlIeH7ZHz2HTJO6vzHn0lDF3GxZ
EE9ekKaumFT3Jaf9et8+6ZlT641hWPCIEe8qQb7Vi4f+pp7FvqbVtCKh9AhP0tYe
FA/jeMI+x8osjTvyp/pNJAbMQHkMbL3YL0FusBO485EYJdCj2z5VRJnSRIc2ZkZD
sI2jkdYAj2KA9R6TSkJTdYbUcNx9hLZkSjCp+uxq0jwsxGIFy/llBmNjSvmfCTe9
d7wCGs1eWvae965JT4mmcDnNELe2Yyl+IXA+k6HNWoCmAiNOCzNWEI20WzyNIuuZ
AWnJdSxKnpN/d8CtQl46qgR1FlUwJB1dtsvMp0Ro63Y0mEy6Kk7leqesrMujAKaW
cG+NDAwQNPqZ2OIZACfkuizTeP8YoeEV74rbWxG4otgMgofdfDBHLkUno+buFB0e
F5RpBe+pJP7k/LXJ54wv6u+4cPf0cj8Ubo7zkRp71bzjX082HIOoPWBLlToX35oM
iqxh5SUvE1L/HP8YUlyVpgOgEDsjadlX7Sus8b22m4XPdDuMvaCWtGg95fwh4uIS
EaFmEGFguadCKyPJZLeek1EMztqh/lyerJsoyKVyEHn/neiSLDRJ42iVOxLa1Yzz
ACOqORe8H9RN0E+U0lzltOmTdvOwkeL1Hdv4w0s/Hz2DFIR9rIXN7CFkSZCXR2gC
lkrgLcMrQCXAhK9n26khNYP5tKMe+xtiCIJwzyS+78apAUI6/D2GuMryuFJORo+D
VWayd3XMC7+UmUDZ4HtiFp7Qwgm/h+dbO2TYAvfF98SlsKn3lWgfw98C7EfjfqDt
2V96+GdcE0wTHNGubwqZ1/WmQupuIzSczyEvNcjzBWKFxR8PfS7rWNoNyiBUYLPm
8mTsE3ogMSPSAY3470HgwneV+S/9VQsus6lZRrkDtdq6PPOAH5xFqU2UMHqri/Fn
I9GaVvwVkJIWYtiDG/OIlNeqhHpZ5OJz1l8jj3au+bYtMttUhzzysUFQCjeKjtCC
rIHfgGxZpbheSPSJAu5RWie/xdOpRtoxg8GKdM2Wk1vMcJAm8h6LcYpw5GAsZyzs
iWQ2gaUlXCVTg+u+lh3APwT76bWzKySP9J34d+FlKoNK2LXO1uQ1cWUqkIaWss4Z
7hSGI8CcaKys9rmXfxa2/1rUvZqWWDLcxJ6NlEFhDRP1YRPRm43FAfQ7g+tBxSTX
fzPShKOe+jxUuDTtix9tN2Y7klmuCRzrT+sDLLc3E8uTgDqiT7t8EXVb/obDhjRV
9VFryl1aM5/tGGEZhUCSca3HHthdsP2lpe8uEA+VBfM8d9e4J9jHnSrj4nZFIoVh
l5n8fOyRlMYRLfnFTfPO70vUwfGB31ICQjBgIW04QlAMPBGunaDUbgCIAtiew/8R
c50EsGwper7kpdih+bPH29Pjqm11HmT+9+wn7GsvzuY5nXfq9Kh9vSPCdz/Se3yx
WHss7m8WBoxLk/mDo2WHY1e2o+Epx81c4QK8AikmlyujHFEXfPG5XK7OKURdkyKA
h7XQEfWaM7wqQ7yAZcZmoMwWgBlZNZh6TuxjMZtgZStr6ioLGXzouQ0z8a8n69Hb
KJ3cLW74JjsHctDYpCoSuiAVi/HMQHL/dbPvMWAJlNL6O3JR5vuyddVPt1TqN5ZN
H/i1hd1Q8GUZJ1gZqiCwHwWi2VVZx8D7jQUG8C3xsKm/ualttwwWuii5ejsmBS31
ji1/Ms/iJTC3EPl4Z2CoVn4mOidvQ/UiIBV2MdL6ML+cN140MiAaP459elEEWt4b
a0rjLHgDjworJBIsrotutOyTdb0IAGBrMIodFMx7o0OGWdsZ/EVEXWxVYIdM8f2j
nQ3SqQd9iRRROMeKdddneIDVx0mGHgrDAIRE/IZ5EEHPeuiDlTo+3K8h4aUDk0bF
M/06vH4tqvNEULZ4Q42YmdtAqS0ZlzEpRYyeRjvGUnOZZ68HHiU8fWl0kQf0vxVb
hOw2pZmJr4123nfPqSAhHE922krPnSXuaLRP3ZFiDfLqlcB9pWvAlz7q8LdyLw/0
oNw/T8SSt3f+PHp/2+ffCkSxSURRCAkf8fwBP0tbz7DvJYY8JZxyWjsFvm6zAStW
9BFaxgVXW88shUnqI7QrbZyjfOlLoynpdKNHceQVtapVjHjenA3sfI3IGCY7smOY
sfLJ/TeVgaOfIA40M+nto+vjqrPHraZjDrFIF7gJg3CbJumnaUppHr5OCdD+m4gf
LUwpyi7w7j1BOHMv7g0O8YGU9sSbtykFJ0WdbxfDtVB+fpnwQt45LS1VvA9eAOSA
3POT5Fbv+RMJQOcdANgmXtkj4MCrRsMVGRS2qflSZC0VbWIPU4nYy+CGez+nO0J0
nzzi83aVFTOUMnvhuxLET3ssoebrdqXDo9zGUK06zIs09EjeeECBLHR9XAsJIldC
KaQCLfyjIKcaZTTxxz4YFfun4MX6klUMBXHsn8uEMq1SCq8zD9owLzRqUCHxqGIh
Ll/txajC1FJkG8NlGAKLiRLNXALF1dTt+5upmoss0bWx16YtP99ULvx3LNPQFQxv
oiio1FCcY5wa4W6nBYtxX6Ja9BeTyRbpOrtlKO6k+vvnvZidK1ZVoAAJ9B51EfWM
Zgu8X3y5S6Fa89kgptKPJHZ+ID5Xux9/powCji78fw4CprOqVd59v8DEwU29pPS+
1Kk2gCMHPWLPQt0oPcvBlt6yWJZDbKlE9d7LsJjTq6UNVGDyF3YXAhhYFFN2o1W9
BzRdBD1KdZ6aCbI237alO3R4aKlrSKFTut13unGXREDi+GXhEGXixE0PPx1fIOVz
dlonB5tgtetMfs50goMw/3pnHgyGGy/oTbTZskAQyYayOmknM5qzlh4aN4S9SMJ6
9zp4HoOrgOvd0Cp0T1BhEOPJLbPmGWBwSUo4Oxmqa2G3pkTSe6J/G/B+biI9vjAF
EWjfgRFGeNdlBZ6PmOzktSrRIbBD58075WR+NXOfrcbLYiE74X7Ky0bPwwZvDtEq
l/hDeLbzBEpajaSNlzqQ4qgOHNCF62UmS7nwyDYuD6z3/9NFATnJALszUv4YFyiO
DZyfafr563EV5julJ+/YnPn0PujzAyP207j8pwxuOiDrNTYlCs54ehu7boJV3ehr
9IMN+udUJA0tlyuoUGKq7zHV0K5ndDiz0L6Y33NZA1rynaVzwlucpYarnjSfIacP
tfC8+BcK+xcWfGh4hMRVUHDLRZ2jQfrkqhrqCQHVDsgwpmHPai4ja67DXxaZ5vTH
QPnE0l1FEsf3R9u6XfmRqorpNtIevoP+/iibrIY1oXQNrz5J0+9kopTeYFNmozgF
zRfzdc4ZPBsb0SUfBbYGZ3f7i8OSQI/beNLl1UZE6cd49g9Vk8UKdoO2tKvRraTY
0SdvXI2Enk/JT+w1mU6wpUvlOT9J0V6oWTeOW8gf1CwMn0uYj51aGj4kZXknPor1
g5tLFMj3e/zzbCq+j14jASBbmM4p5cgYhYIXJWZiCmdPzGim0XwSfOX75igJysqN
M8t8nFT4z63TMub9VO3UCzfor3I+PkeuXJ0fMuJ+u08/n4O5BmMarQpKbZ2QCy3a
cR8TzdsmVrFy0XspTm2jjQD4nUn+TiU1xL7HzEUcWQRKqKYvDbsJ4cI7f/bPiJzI
c6IyuHd221oYp8FEaUjTriS4btMaTxn3VS1qyVPXqzie9EuJVo/olR1gvNMEHZGL
EE8EBk+aLF5N3htKh+Ew87gaktVtwLl6AVsZTTaeYMG9vghnGDkMZlPiBkungK1F
KkhmGM7Gl8xr+EhaVcCy70IyldBLH0OBrLvK2CpWzkp0zeNKZO4XfWK88xrIws2v
kdOFtPDqkb6H0AL1ggXdcxpIBjDYBidEQvcC2DbkTgniQped4frJfvNMpzRvUkKy
2aBCCvoiehTbmjYZQlBGMMhMR9p6+kmtBYmV6KL0gmWyO4xhPiatudMua/1LGDoK
zRmwAyh2lY/WzfWpMW0fTmiJGD7hd6281jt/zjWNfNDi+2KZBPGqmEBo8W5ecdjw
+1WCf3lRBMA0KvjV3Gyu39k0IY6X3EGPSTOHqvQE1sDwuMOf1txBv0hR0nz3ppyl
O1kbCIp3MVUoAQTCAj+5QgiRdha9BTMHqte23esZ6Ev5LlgLRzAwKi8qtw9lRW3K
PQ7MDJThF3bBiyfKtUOq+EF84WKx5vty/ulRmniIs4hSxi7/vbeYzpV8ndFV7eUW
vIDF6TbBdI+P4oRqMs46irSQDJJpKPEhH3l3PncPxIhHPXrd+CmJSW7e46wu/avZ
ImN5bspLa8JcxpLmMWekwS8ET8bs98C+2QknjoY1YaxPj6zCbDR4Ajd8kasVBntm
O04LFre96+M2qy3Jt3ghOFhf6awJpUyU7o4Ug1aAGXBzZaDJPNLVRppTFk33+GI0
PSylZkpKChfia0Z+DcoBwNdS5jKdeatPQPct02FGBITJQrViJ2hIlJ4wmNKbWRtb
xXQLQv8Z931EhrKolzom/iKdi+S9C89TjsnlQQVpok89PDA/hWZJ2cdV81BlNgl7
LFrxdR02S0nf/fpNH8MN7QnO31MV2nhLTBm8rZY5DgQi1QKMJFEBdVw0Q4At/s8R
piDpHy/7hzVnOnA3VyYAYwBJiunVJD9NqWGV89mXUg4Gom3bomuzztrnyyh8XS8s
Uom/rd859eh7TmsAPb6dOvBgutI8wcCAXofSSdxW2LUXFeFgcDgpAMVUOhnS2OKI
xI7GVhL2j27ZAOx7N88Vrrwu3ASr9CMmNw4CK73zWwKsMkilGi0cR6hJ89PzS1gq
3qaR15E6wM6ldpY5tycjItB6p7RD20X2eLRYcENODBgOHh88jw3WNLaCnpEch2FF
QehrGwJqlB+Cr/uW3SLD9Sl5/fNT1KZ4W9F51AW1xcNcqQYZrXbuFv17RziE229U
VdI7x6TLNPQyoFtPNX9UInI0AdJ02eHwHI8k1imhO8xoTcuZUSopKB90qYvDvP34
GSSHUgcUQ33FGXCM4Wsa+QOX70lMhq2Oawu4AzheQhUUuElQk0LSbUyhKhFey5Z9
uZg5kPpYDdMa28sQpPkXf8EhsRB4MzhF2o1gBU9sL4tFC4n32gzZLH6ut0HsjO77
gRZsmgwDcPMjvdc33GTE6COhk9Xrf5Du0sCXL4L0v0tBJlaVCaZs0IF43ECt+nRE
FsFqabQbrzwoSKDRsKI8B77GNanCo8rLOi6oNem7h97eDNkLzxBzUcMEOxa1QCcX
Wo5qy3FOTAvkAYXHSstvV8TcPQS9oVoS+XmZRGgb6s29PzsVg2vOo74yBu6uynac
afPz+AACZU1kziDNSxI/SnDgdtW7CmPRN61gcqwWomXRcVsFcJEc0KKHDW9N8km0
2FrdbvUy7slfVWi5ATI9M/0X/lvUrQAnqmoay7FXwWrjnAGN3MN/Q9F2anW20eSY
9ezD/JU4LRuAQPtlDP6lxMpl19X//3UKM0+xv4SoHB8Qm6xzDKaYo3m/oh7N7dFC
FDAWI4nuG4Hjlc8PZiZB41zbN56U1Vo7hl27Sqwh5o+jpOpMyBjnia6PDnNE9w5i
M1IP9dp7xSGi1gXPdG1YEw6+fCxNYLaV6cleEb1fdS3eLO6lFm7MYhryMF+6MN9i
wSIFpgWZVE8I6Kx70fBQCZtqWqPUieOB4TEWzgW4DjZD/Rr/gB925yxE0pD1nsN7
GN74bQaRAMncmWTGW04b/NiCNQwOaY89dthBY1QH0vx/vhE2g3DJwH4eIkuxmh2z
Q6+2kfOE1svmtD4qpDwHGTqwmI7usWJKHP9QTO0ue215Y0b/EKVWfLXW/5L3r4lb
u+IABA5tUHT1904Ef+9IrERh7mt2DH+ms6AtYx7sys8Zu+L1e72KrsVI0WGnmrsa
mEmLZzAidQqqYLc0NYUw+3kHxdmNpTw0cMy/dNfgMEV946WMXiSBPu7kKhzmUz3K
GVzun2yw93j8J0lY08qaeX6ssaV5sqc08BYoiolVc2icpDsCRcVT1pq+KILIqX+n
M86O072f5/CWH6bsaonMk54Ei1VXCKoj0REM5rb2uoxt2Bd4l3xFUeEN+cIRryfj
uCkac9iIkNM3XhhWTEgO6tq9c3MOX/zpubNJUrTG5GPA9JgSN6NUtmh5iWDed6qr
ErT1hndaLe82wtS3a8Ppkob3MNQhAJIaiQe/aTwrb66r1vbhG7WeNZ1y4XSMPE+P
XdvnEYhZTmt7VFCRPzSpRl827/8rCit3kL0Xk9aWZaJmeo83Tzk8WFJ1dcSSvplP
p6nmI8V4PwIfMwtJVto3ibbRblK1OzK7ZVuyFcj1ZHHVl+UADQ2Nh1rHdwCsz6n0
hIHlByZGlhy2P7yJtRg7EdoHIi6Mtpl8Dm0VnuzoOsmSMDAfyeUKYNfotcC+Fxwa
w56MLndmYrnjUAdbWle8Pl9yWK0WUjuZbKVmgKz+pVCPnQVPUq7Yy2lCBwRlIZUF
W6ldIDZcaLM0vbKTXU6D+YJrjrFc4M2UamEo9Ddti2b5ezATkhh9amJarN3d3vr3
TL3zyPYaDL2uBNKpPj3w0ihLbf65mIV4O4TqGd/P2ddq+ij+33BlBgO4mq8roPPL
BNiIUiKFWCymuW4ZVVC1NjWJiCGtnp8V6sK4K9WD/V3x3uF+UA8ILvEpzfjWgX6h
pqkUY7jEx4dxmzZuim7uwm89WxnO7ShdnihIMQ2NKquZNkbIRlahQjn2d3OOhfKK
bv3ugaVhFUfgPY95bVd0HR+74Q2ZkegnFMKs2zPTiHhm+3W98xF7VRmFPolwvkow
xIqUlev0hVDfdVwkB4vL+Ke6EME1UCQirsjcHXx1O70AAm38E+yDoxNlauQ02k1r
VCiKUyQfgWXb215vwdRG3NDGB8IV5K/JNisLnXWB4mUEgam6rq7QPfh7Dbns8MRh
ThzA/nCI04K6V4pVIzr1u9sIN9+Dn4wd5JvXOY79SIl4bClwPwFDlSEYvo5HsTA8
g9cnSguve39wHe3KJPb0ecSVTkHprneQNL9m3lHFuFcQSj0dziQ0XlGpw3R662jy
REdbDeCF31dfoWkLJps8Ssy3+10q5QbJSg1ja29LiCoYgvkkWrMeAnLkcZIUMGyv
vZ7LesDs+EIqkWgfyKJmz/qgLWHGxmKhgjzi3HofNoscxu/iHeRVI2EwxLrb6kj6
NYMOQVF0DJK6m8dqcdcF5Vsc89wkv7LJLIWvtZyWrm8XkOAbPtTn0J1ECQjtA5aW
SUTu5zVbbdx0EBKc0esCIvyiLnEASNBjk8xoXuIq8TPwcn2HtCBSN88v2nkC6ovB
S8PXUDA9rxBwUoqIHb83O21l5WEaMGp7b/JcAd0eS30B4hb2LnH1kjDePZm+7YD3
UxPBIy+J0xmTRSx0BwWyK3yUbhMUxaxO60yBcpUfJv7LuEyFnqIVK/k6RoQvNaNE
d4oU+HURt5wjn+km70qYUEDTffCtQNn6BrrHJQQc1hwFWKumA/LjO71CjHzIMiKq
WoYy4XGdWwOdRScRw/0EJ/F4LuPF3s283ZVHv8eYIpF2Lq0OgRyhATOhDoezp2bS
jTbmTJzZNfGAoF6byc57vkTu78mqXSmmrjH23j/Yz7it/DSPoEnweu+7UTn6vmHQ
yRrtn17ar3uBMPcFsOpGdAep0PAe1S+vkJZ2rZFqpOTZgTNJIPj30CZOerbgQ/Cr
thEpppHCrWX61SlQ2jVmYbKHM3AlGaCgK8NHvQF4EFQme0NQ6PcgmwmgOwQOk9Er
HlsxeazCiK6u0CcVhtSyrDlPOnJ/0MDOZy5dXvtWp/vbdHR9wiZAl+X1tJi724kp
/Dc8vLmjo6HXlESpHn2Y7sFuRPuKVH1sxaungjhm9LnfT2uq7efPwoG38nnfgJ49
8UvWYSI3l+08Bm/YztlAT6EC1Pr6h1h9Ztbx+AbtnMsnnNzpmW/MwCD/7dTRR8kV
ecgDIp28K3coKN/3sPs7sZ4n7iCfhBHYel0dfDZ38o/Ccw+aEWmIvOXga+rLjJ3i
xRX0SVQfSx4izbgnKoXuabiS2/FdgAiWvmmpLObviCUaRS7TLqIJj4Zjr1eIXc62
dP3SsU6IGAPxQ2aAi+8kjXfKyVmPGcKapIAD/gSDrM07wixJKTsm0XVQZtUo2N24
6VYF4R0wbpHaja6ps0iSHLW0rAsk5i2Cet1stnChO2Oe04Ab85AfWBn1elklCp3G
IaETEYfmlbp9kmVTzj9aLzJMYJahb5zUMd49HHh/vM/d1Jm3ihUu3WnLDzaG5jBz
uxqgEDGYQeIOj9pPzbgob6K8YBSyyqb5EnLKnpmFZ/S5zhzSGJTO2SQk0DzB3HtU
fH5GKESCr15tX2U2L00QNHWsyEZ6p6vJ5CB05cBYuRDkBb/xk3GI2M2V+ONsnOuO
7VVGR04NdG8v39N2gl8b7sL57+WKTpkFU1hStgfzgFPAphnTlea5uGn4A3qgJg2t
TbVp87HQc/rvfZwmFEuFBN4Dry49T6B8ryzPStAd6wONsXpX/JbEJ0AoHd+JNGln
59ienFauvVLkRp8TvHP4oHf0g+Ve7sSo/yfwYCZ0tYMvsN4VJkAlabwbrLDFaAkn
U+ZuaWAbh4skvtlgSTZyvpTV13Rm6CqkquSeMYW8iN7JLx8EzRMNcKziKt0+Qs4r
3VPdzn0SNwOYK9c4VDBya1oVBWf8UaLB7TSmqcOLlIzJh38PRgzFbLckhS9qs475
ZKV34gEjCcIHcMgS6AXnNRISfJlwDnJk53s8VlJnvfltsxvPylCZjCxCB/GP+mt0
7/RI2PI7YIi9YeuXR74jW71RQdM8HwpkIQR5fp6y7SCTY9McfMDjiXwDH8+M8SKZ
AxguUS8UOWuZKPgvd8f2bnJpHvnXeGCikUI+WLTi4rr4P9U1pJYVm2fjPGYUAbyC
7zcF0zFBsqORHdBcDRvMZrh/rFegPNT0Mj3dWmgjdKP09CehW/Q3RI3uSZ2oHzl/
jOiqm6H1lqJ+/shTbFPoR2jPkfPsrQINphOhRM8xxEjhQlk34wi2AUu7VtpGuoWK
YyhFD94z+gC1ChIeVoUfCmwmGOg2EF651FW+eM3rh+YMUOiyxX9EPauadxnJL+9R
UX041Q47rcZKhNdUf7NiNohXWBc5d/wQ6kGkgarzyJvLPadkLCZ0l/JC8EbkYoRe
2kHe8dWfBTCvB0r660gSCjEBnvrs4CQxHEWqPnrlg4f8eEXDI6E7P6IoyFm8xHvw
Q3ax5ORz5YR5iGdYY2kxOlWS0cWjhixVuPijtzVNWWU/W6pV8WLELcFHj56/fCvx
9/kbn59M3w459hIJrDGeCMlNEiWqaIr6rgvLZHLMfXupFTSHE1SJ04Ii098mwvKC
HZVm2vvibAMnjElEtvrhfSZ6Zy+BNuOzX/EVwkXVzv9+H/kGKeNONtgZCISD9i98
XtX0M6zBeRZ16sNWoT4pf5ISigPKY4HZlRDbVKivhwneUObt66S6ejPpLmwL05hE
6ncxVH2HzZXOQQGTrpohWUNIwVqR8LyytFo5DWPo9bHylE6dgJDmT6pY6nJ0l4+v
13D+LDxXAxfIIsD33hDzeZCEsDjT3r/s742EIni/4cT5neYbgHvBH5ZmRsICvSNc
/lWJuBLo+hxDrwnyZaLtC1FJD6r/o/aFk1wKMEROCp7OEPEX9fLRLJys/CAGlO8n
TnWpub+gmApViyFyB3h55S7HRj5icjWmwNz11fMDpmIUX2QXglrNwCMuR3w6vdD8
zRxRxmUlhYgPBy4NhWuR9glejAtWqOmvdIMqpBmIYjuLGDXc/gV5wT4IQrs2xBxP
WHMNs+04HBt1FjkDMi1VX/GDEfStU7CZoUP7VuDaQfOkgBxnfIPZcpvIdRVFi6Tv
wXuiGvNg88pbi3geWiOY/c9LIXH2nJj+q+OwsJs+elsC+kwIPYl5NQ6ZYdvk/0SR
4iQgoweDqxCJoGpNH8GtsUP6vaXXv82nE7l7bTPtID7OIJPS9I58g4Lqe9hSdxLu
useQ5z4mHGe0nGKmXpknoMrMknPsQ0SYmpvR6e//9UK8y3dD/K1tBWDUCd57QA76
cbwNEO7C4A0eQJFvkGTTpxBwk5YEgbJ/RfI+q4Gahy2G7E7rE+WHFTT9tIoeoZpg
VD/I0mjEHKsSSTZkCzD/ceGtdZhjFeU0/18IwjpvZJ8UiarcdJ1XiOmaig1d5FFW
xLMauXd3BhN4CEDLcOf0dk8FJ1V9vpmRSoC3yZNGqnZa2Cjr1PZr5vAzNujWYaVO
weyGh+QDaiAjTc0bY0449iJqSV+ofIdBJ8NJXQSTVr5PLYgSjmEIR2ZuyH4Jfv6w
DqZnIl3JYXcucb1HQDgPeouJYf0NMjNpnQqXtvj53G17lkQDx8rnN9SSDu0Rwxm7
1PNRZ93tE5fzqUuNU3qpg8Yk9WKDfFytzh/icX6aRZJo+wDCYr4XTBsW4IoSB1Eh
ZLKOFxR/73W+HVKcE0/htm7Q1wAyIxpWkUxFjZTCpj9omLwRXmq2CMJjXOarE6oe
QfCcrFsk9eT6fO7WmLdWuIjY13RtDjxbhRo8xiuuoRxfUd0OpTp23JarrVeEkcqc
i1ci78ozr/KedHeVh0SHtGz/MTdgTf615k57yVNV7qEhWBCSPI9y8kkSVmFlAJ51
6PR5iRNBZu+aO53l1J1g7VJ8sHpt+jvj1devJ66tMbMBWGEf6B2RDR2OZzrnopVM
k1UqKHfPhUOeLVWoiGyjV4mASHLJtV1YnV3yTd8EuMLQBktDHL+Y/g+3noFViir5
M+lfo2RrEEvXE/5mpbfi++4fyqohi1Xw2TSdG7MvU5NGEJQlIJJuVC0wBzGfDivq
bfKhVT+jdS9xJl9QvJ/f0X+ayw5N16m6WEmlJHQ2+3NaYO2vVooT1uXPaNz5a0vT
3wbV0tH5PsUXmZychTi0MMFWbQp/inPGDLO52fLV1t3F/Wqp6T2eex6SE3fKvLol
A3+xmnxUKBJms8NaGRWLpvy+4zJdy+adebpX3Ok1LMZXYT/4tUBgbSXxdwaCvjwb
yKpg08/CHEcarFdY3xVT7aQzD3a0JFhYOk6YMLMMyMNEgiOIsihXXENMMnr3XlQC
ZqiRfjiN8PC/LvZOcAjmL23PwPfxWevuhtyQBSblWccPUy+DMBkKzLvuDfk0a+uB
QbRKZ0UtEte0fvFpxVmcrFbJIxo4aZw6WEZPyttn0s0r3dbSU59VhAueJi9EirZe
+squ+ksAoA8cbXMDgNH3c4Ag6JUMJ9F2XZxW6iBgbN9OzZIhZdVCdKSxxvSV9hIQ
36lAbbYBFMsZkJpe7m+1G8HfWSRM+OyD5Sdb28ZUO2RWGGCM4/q3ha00pwElJs6Z
IHv30HFPwgjY+gcEQO5KCIWYL0u9+uAUH4dBAVIK8Ofjp+okJaCxAl0uy/cyp/Un
Ql7lv6Xf0AhMhAqJPOkiT7ogaYFEX/HozmEKyKNb1k7I4WRGXMQclgAo5XKCEHSO
a9JuR+2I4Vvp5+wfBMkuP8s9Qo68y0M7lU5PEF86yhtFUa73MoJpHiuFLMC/pK+f
K3fwX+kTEmm4At3ugsuN9acrPQPSIxmIsVgs+d+vFLyQJVoEJsxmplsqPdHSIhMb
zpkVF9O04pZe4UY2XDbq7xUMHS+otwAGl73FIq3NFu3E+Ioq9tj6uyCnhXRYCRhV
/ochSpf2oTLH5e45mD0SpMESgQyA6VVVhZmVRqlQIoBsfdXPhX8DfwrQKwVViFQ1
Rwd7RttjDwVrX7iCLPYc4ojUBxgE0Gk5VCq7CEjKWTw+LCqSetsDGK0UNDja+3wz
nilj2j6cK2+3BbceQEb5ZEYZzMnZpycTvktong0lUS9We2hjNJ13KAQ7Ikksmag0
tDIJE0zo1fw6JvAqNIU172DZ6qOOrCOHAjhvMAHTJPzjswn0kumoqX+xWFliDR/m
znjcUE4VrXFGc7JcGP3Ob/Whi3akdEP/+C2IP2cud7Aj2TPu2HTOZWGvwyLp3WwV
D/AIuaU/4xSvqo2Djq3x4FuS9AaeC+1RQ/4bnu2pe6YgOtWz1sdZjuc/S5NgkhBj
OOKoykCNMCu0tbR6w/Zpjysd57GBUG0G2Sh3AoZWusFX6D+UZUa1DsPVS1bmWxOS
5oH+BbA63i2H0U/ah0iJrYJAtxlj4KEpLlvTRZTj4NSEDxk5bqPaqo/LtbOCp6ln
kvqBF9eg9LNVfS7lx6gqJ6Ly7YgeOitAgHQfBumj38GfA76RG0Luqs+ODAs/WTwP
o3xe9WgjCfpaFflL6ExGWNsUTABKpsGAbbN5PiTYJyDWly8hTtuan/3EHAlce0mI
V9meTj7cOIOLBCXhoyhWcpNwTEG843l/G2RZBZIOLesRp+JtYvbOoltxXPCPBeOd
xjQjXhab0OBJxMtxboI9aepRBUEGf8bHpSjuX4QSKK2i38qnzJRb9N6dSqSEhrx9
ZrkK+NZkW5OZ3hGX2osTD8E2IDGXt8KQXKsR2khYeMj5+BKahjZlbq915IIixvn6
NvL13BJZVS1utnPKDPpCoetCHCivBiySRs75izWAZKMeOtpR6hL3BxKk7biBc6Ji
WaNJuIDyNHaljOVqYjOllBVy3/0kNuE7PYqc5DOaVQPKj3Rx5NGkL9Gy6405j/ix
qFlz8qYcphyFTu50kO6D6FhQC5EZKNlpsZr2YNZogcE/6Y/g+YKrYRRq+LLAPQoN
AVBv5TaRDEAov73Lfc9R9eUQ3PGyD2HVCM9fAo891VBBCdE6E8nZqQkZDF65mX+t
ZTAF5ZXc/A8iIxUjOvglHnffMWIKWtPwQrm+S83jrUf6SOMmlSaBIIvEDmsFsoIy
UYl4e/81qOuHuXF6ftSJGNQYuft9Ps7bu0i2z1vYOPc1zqlcIrxsvxy29DLb/ZUK
4iHZdaMaeZ1GmjX/BYCSJgkU4QHKP0GbkTsh+9XPX44eTfyo71dZutZEn2Q7nsZ+
fVy7IS2m7t3ErLsimMHy6DJCLZGT2SwVsxKh9EsgniBExrPCSVmThSyr9gf9lZSi
I0XzBLXxDz2fr8vHS0I/8mY13hp7bd+uZsNcZOxLb8Fot7kYyy3hGKB2pNqWtoq0
U6nBH5trNa4goxWvWUetQfYtPCceexC1tJkzgY8r153e0jJAXdrjvShLe3wskG+N
x6DM+tW+uw8jbJzfqzzlopSsOxNqKFD5pGd1x2VSiiuXyCd/gIeM3gaadrrtGYWM
LrWA63zSl82noEUcpuMjRLy8Z6v4es49Gqhmpug7NwXrFaA9c8WFjx9okvm/JI8e
fJDS/w0fyLhG9vsJXQO9LARM7+Z0G+MAXlYcVl6n4EeAuLJ3XHcIGuZuL5HeKB5J
MPCIIxQL30EVe8eZVkZxBhufKprw8Z9JL2ErSigPWXJa13CyZ9D6ZU6RNVRTIrdg
xiQ5CVe8IusRA8oQ8QGc5PhvgcmeQVivKtRwu01wbCUoHg2Ha/oeou1gQFfbe8p6
2SHVaGgN5nDSKvpTMRuDYSzBWS1fPhu6TJa+EswLlMsNXxNwlXShnWdQ4b+51JBV
dNIK6Igoh88lea1bVG9irq971yu/7InYiT97MGaajjeEfGOLPiPkgTOqSizIAJEt
nNAq/ZPuZytLmMvJGEKk1rlrpy4tkZZfMFhoTW/VG0zoQnc01NBmKULE/iMP3ks7
dgSglp31335qfggBkmp/uvEQIXLzitURp88pdNPKAvh9c7bgiDy5G6Otdweoaj4D
cmyVlhYnJsNQeELgHpysUUG7Rykju0N8XbNiVKz+9SLViMbe+3RpQmiX82ADEHGs
TETf5U2yPL/9umVO3/+mKZO0ouhjb/5aom0Lo0F0UpaCD71ZZCez3GtMtD995T3v
yQcqAZn9bMw0Osx7BgE+o1Jc2f37VmRxrKAzdu0KrzJbSlfd9O7ypAKr7wiWzlcO
FpiuVVDV8ZR4wb7Z+3M4r6tR7bssmTEEsuxH95zxVbTUrd3I9RSJ91AMWruwYWQW
4YOIC3KT8GsdGjRqboUuZz9Dza96i017T3ob95WRG67BuBxSnHyDAuEI64pbXvX6
LOe3lT9qVwaPYmhc5lA86yZAUzikEZOw+bGYCB6EjUi3AOTifXJns2B+le/AHgR2
zy3TdEVL8LQcQcfLP4jRkM9N75YN8yjg0wohIbjRtkgm9z1Q6f/AhY8kEdLen/J3
oERsJ/yiCqjRK2jsQN8n95LGovJ7peQdwgY+VdBZA2MZztP/jUbyP2JdyDVJAigw
vTEdZj4pEyX80B9DG7dsiYCjHh2BOzfTFBhnXxuGr1RBxMxMPff1tLMMeBgwOUtW
bIRPz8b81XDcMWEddV59ZLFsckmzLXoACBN4gCyrM5k8tozLcq0A9G5DCxMKnCaP
WZp69mMHnYZdMesXRZMbJqMBdVr+6pVkZodShiYqU0PoW6nVwH4jEXJgIVoqCuGD
7bjQhrNLmmAc7cQTUXp00SePUFhEXw5VGWy//WTbPtSZFVG3yLvLyhtpVLvezRcs
rKgmXwQgL/ar/R17d84cG9uH4u+muquKoBEs/OBg87xfbNraAsxb02oAxB4aFnU6
NN8B4WsBBR4YJAIBvmxISzQHkeLYBGHxNcwH6nTHOIGr024if07aByM8BfKDP2fC
5QaqtU1x6bxjrgc0v+2AuKhH+EwD2XwJYa6zi+Op4ZjXnY3Q8CfhaQ68zCYK4C8K
1NMQr5pYFiEaZqC13W/d0gwlGV7SfVPN+8MxIAGwbvSlXK6UhHTi/JBBIocGb3+6
opXNBwFglaPmMBtDoAQDyblJQ0RAj0sjR37U9kS58ky8afhZDKSrhFdQECi5lkvU
IDyXX+k9Qfh09aDPerJw8QH03sckwRHewfX0MmRKB6Nev+TiqrI2QlqUedRa6P0y
qz5s+julKtb2b9kIq+kXcheQIrVFCTUDgcHXFqYbSiUPXhg2YJ7QXcAno1VanCz2
yoqM2hQHOtehXpHKrSLVDu4m2TMkxD4V9FDqHSwMp+hFml8BGneqfQUo5I38ERld
T/9gHEU1SZTtvDkRt3xoppS1GbwN5pnFAhp3whUrOi3j5IhN0OdPY9uFrbkpPVG6
xPEHPf1e97xRIh+AklWIbnK2kiud7iz/9b1rQFC7FAIHzIAJKvRPqKMiZFq4DqXd
iSzzcXjCmrnjuHS1436hotiQ4wCL6JeoscakhWXflEnQeLvoI3QA3iCNOwiVjLcP
HVahmdqhZPx0hYNRvyyyyPTG+ey5iWHjtasq9lwmkAE2eTn1E+FrqSmoPyIeq2ow
Gn6EY199BZReLkLsjedBic38AELvS1E2LZCLMJtWBHy4rUOq1yDdk9sDEJaMWbVf
dKkPMLWAglz+8oqKIK+tW/wcZZLo2i7JvCfoRMWdnSlVeyG7VrjUjFA8PIbgAsw7
FcDDiaMWTM+cExADRBvlTGpFlSGhEs7nQszxKCLHmxHs6vnhArowfRU00G/Mpaoq
3LkSFenYBpIrA/icZWJrW2OHS+B+MZSaqGdQIdwwvwsMQ41+RP8BCdhHRhEuSStq
WlwdWxcFCc5Fma+OzV9v40s4Nl+5in5n3KlXn0PLBgoxP5prymPKgxGuio/Q1awN
7j5XP7RfaNg0xHiw8iVTMc0vpBCrYshe20lqjHEuicJidF+8RDIgkQ7r23cq/HPH
UjXlRSiqALCJt6iekJd1eUZKBegYrXoDXI97/Y1mBpiW6DXQyfwOoXWkdcI2O1jQ
MPqVhQlBF1qh4nT+KzE1Oe4JH5I2qJVpM++M6zqwZyxiRM40HxajigPaCMHXOWVr
7m9/eeSws/vfS9r6po+kO6n7hCKvhywp07jn5Dl/KDW45YYYSgOcW3n/0UrFbGBh
l3sM0rjqYBYBCA7ikUGUdOUdWNjuoGdDHeBden9ff+bozjWmZOonBuoW2BQzgMiU
N9RS9eBqJOIPcfGfgUm0ULygfVJ0Dq0uBf70d8C/3vugsq9Dj7tZdKhgw5sLycpq
VMp48h0AoAO3xhulkr3cmSyaA4qZnJYsZ8wKdxUgCOAMVJFMkqZv2bdj7I4p6Oqr
jKT9TLWcGFPI52y5FGPjo31/BXoXx6VG5H+oev1FngZjenaPkMIkk7wYFf6PkO03
zp3DM4brSzOpHxF+50/lMOwaV2ImV5WU5OL2RJVC0GPVdpWqUvrJPDh6uaUmJLuK
umJEA4hps4W4G5ugDQl7I5lxNysxl0+vqLc5uMMSGnnqWCeDXNH5CldF41XzKE99
NXBDcDMFvNpr3qaKXqkgkD4K7FKjb7RDROUpTuymnzNUljSdllzqWIYueIPOPYkW
aDP2gdfXVDmAbycmubMHJWv21GOPbhY2kBswQP2wQrEvKxhcLsZNaZLJA8c2c2iR
T7l7bBfjlDD1bHkPkVo9wXk8OGFEWu+inLKP4mkQTmCPb70lCQRXgyC0gVFqMvv4
N9r9zmsZ41RT6wdGL9PL+fYbSqzlzyOSdeSxzYq3A2Wwm4UpHuN11cG6FK2MjTl1
Esv7ztQOEEO2Lm0aLx6AEKf4BOyWgcYfe2aQ84V04JAEe755RuMbPgCa3PGHeQbt
LkB/wT+ba6hPPHzMLcmZ443NQha1Th5XKPmGFMpFyfBnggZfLT/0Ac7qkdo08v2e
y8HkYXsWdd7D7hJcMTRq7qBhOeL+5fNZfO2HgjNKD+jkBwrUKs/T3MtqLnKB6Wre
DqzqM+nUoouELmFiUBAjvwYJGrkEoE5QpOrkKBymOLHPmdMyxSn3f1Akh8LXSPew
BGIBXCaeIc+r+eres2QKq4SbB8JnwuJ0m6NkKdVwQ/Dt7K9m+m7p+RJf7X8Zffa4
Go1HPrYVQ68Zki0s1CBOMhMT6tHDM8beGnjomGHJx3g6esiIhFoUGBEPgpJRCtaW
Ww6jEeuYr5GGUaXdq5ub42fNM6RJysZYjJgjktDv4y1VLqwtI01WFYKZtm232BG0
G7sD9NZdJ4APdBJ6vTxh5qpZ2anU8+7D/LgLWShUv62FFF1QvJiB0YLYLCu7SSQW
4N848ZdZt7BLfEv13SA/CRvqITrJet9RoHH03SdXe/Zghly7XPCPoN0ZFC2dz6A+
Soo8SJ2fmj34Ab7z5cPPu31NSCkh0LjNl7V8j0cYgTDgBg4QmYu7Co2IHUvgoxKY
n/J9UpkPvqbCWiE6GR9hUzr+uf14kSKLiPRvDjRtnnijlREZT7wKIqJ2P64W9U+r
fcZ07EPfC5BtQ1yo0ARyuuKEg1YvX/YDd+caG4Fp4+fZqvIVNonXUUyREdaGrPYP
Hy2SePKjEXaCPe9RY/OHf9d784cnrd2WbzcDq5K28ax90r8ubjnyLzNpCbet6x5n
lC1OKQRuWNpBFEXvgppd2FstEt+vGSwQ2d8mn5K+9FJQ2Vj3hf29TNNCurqsMBsP
xImXrCy5xLhV1fV8sOHvFFIJswwMgNaxjrxdMFxCjL0PpOO1kil/m8wxIa9YaZIq
3f3sVEGm9FD3ZgnV67uU/BhfE6yauFyuB/kjRYmKlqLZq4aS3epYIk8un0FnrHQl
vtNVd7Gtt0GNJMv38AjzB+YrY70Ks++51Iga5pcdGSOPfrQWMJpz04vYZSManEQD
TTQ9tWl21gKgkPP3VBhQs7YLBMmpmth03CTaWMRpzQ8WmwEdNJ0CwVVE8D3J0CG0
h2FssvGDu2wep3tzzJ9C0bubT/3DOKKIzN55jfKt2hty47zdPjFKdDwV5+W4axBI
Hoe/37osgqJ2KKv73DvegckYEmvMJxKw48D/0FwTviZP4b/lTBIq+8KXD4a04lMH
8LbkGBdLUfbVkEHq8NdP2+PmQm6MGVfTwY108axQbzmsdfKmDZoVHgAEY6M+mnS9
VZPI3J4jED82plmfAhvJGEGJFdklDY+ZLNgxUTtjOY/qOQxDNcx+UgA1RqAW35f2
hGNX5A1OEjdmRmP5I2FuizJubB3Z42i4AJo23IQ6z0aKmvDbhC3yoedWUPSkpRYt
AwazMnK5gSYW0cS8GFqatgjkE1Y3aPqRN5uWKToWG+KyuXItvVt1PQ8vf1ewTAH4
ZxwSZt/WxQsfpA5hMacUTzj9/quUoNXSG4i2LCuCR7yH0LCzrgd0SJg7eEE0ZNqE
v7pF6xYq9UZiKu46V52xBFsiukVoyhKCSqAen41OcIDwchAQy+2OysM7zdspJJCN
x4EEMbaNlNBw/cCPZVpu1D3sQ+cZJW8R7nFk69tMX4rbfpEaaWxmOlmMxRA7Q4hb
Ay56f2jltWxDpmB5e+9W+YscshBiiGTLYtBcDUIxiFoWOUKSXSPQBFQU2LbKDFnB
rnWLer/BoOkU5OUQygUn8qgoJULFEpagypx4dYL7ni93Mka6Z9r8oZfC9jCQOyZx
TtIsYUoNH2klwuqKCX3ZPp4bmP5VscE/+UgAjr48aiAlCafe1diecPZsGU/ywouj
pRQ/ixl66eBMkEbLpN8dA26v6vJLlHmSsC7y8irhjEOPpoSdNMNG/yq5G0/TJVgy
1nOi6n5CgmeKzx6lI3Rx0F4mCX91pOokr+Eny8JtGV8n0a88NOuMooObg2N7s6Jf
cNhqtEPKFMLe9LiYIE7vZKMTnO3Un0w55vVdakz8M+gbWW4LazZk7/VxWEJA9/wB
aISq0TlLCBTpxLc9uLfDl5Ro2ff15n0oSYk5gjHWLw9N7+vtHaVlk+4glf/iaHbe
nIhA6tEo6LSHSJ14abBcqO8m82F99MttsKf6wrtS1Fu5pczk0+OZNQqgxYXwmoc0
GIVRxV5Qb11PMS6zkiOG9RIkdAdEVpQh6jytpNpxHH2l7EtjFxBUNsIRVhT/iPqD
3mjn3QETgscrFc7nkmqlx5lhCPb+z4LZNzsFTjrD5sCKMKJI7tqxVu7JNmvRGiID
3NY8FXG7PJiaqrfxpzVu83B80oBhvn6JUH9LE2F8G6+IGI2mInjzkTZ22xClehWc
x0lId78dXNQLeUZ7fDkBWoWC4UUXlM+Gj0kyxwAQCFjeTwx5nrt9oN67m1cqvlCx
PbgD0GxgZ8RBdk0GkVdpV74QIDOON7O7GElmPo/UHVIZe5aCGSy4z3fCv6yKGJQs
tUty0W5ywcsaoIZbKUT8T9O8fkzNdEbyg790VHNK75jomimiLIE4hA+os6hhOK5l
F01Ll7z89ydOSrjMNaojqBMuz9yNYsYxWPm2XoJHH4ByngyBtwWwP3EdCFmH/Opn
ntjxhkUTSiQcoqRfWFjPehV7Erf2Hp/eGY2IbKqGS1WXPhstCqgjM72o6JU8+cEO
SLJvf/Uiwln4MvgAvZ8tXprRuvm0yPNuPLHmH1toAzo/NB38nIMqt6LVgQlmdAOC
SzwAH+pjEZmyhd0X4RubK5uERROEjsZe4gP2izgM6WkJquaaTM/BIxOq8BEtpLZv
7Si+mZDDyWlZbn8q/jeOEkyDuZZUVnJY2VR5V8FFl0nYFjWI9fWqYQgf0QW6ikvh
qQYLU9y6IsfFDf+FLAiR0Z6pjvfutOPOTvF2yGyr+U3/ftYYlD4tWQsKknY+cnWR
uhUAxw41yZT7oeqDB/nRxPYzvMfEZHgv/KSDPpbAV/fxI9JGWxnc9ZgamAVLvsQ8
Fl2ENf+NCB23ukRoNVND+7SZHM7QKxaHV6clclnZHHIswk9fTJ1B29ysF3p1mnK6
SgjDZCerBLgddVfH9yderiG5O3vS7Ae4dv9mxcVUsXWeqUpiY6pcxVDNXh530Yi6
I5cMjesXAebxtxg4bcjYDz0NAv/6GcVsrDOnakHZnpg4AQHzc72F+lZmOtp55Cza
M5q1oiCxBwau1+oiuagdAqj2scrLgOwhirkX6x1sT72MqKf/drGUpDJfBrUKLL84
S1KNMzkSGpIBoBg3i0oLyAFKo+SMGHEPebz+RNlQD4awHyeC1AyQWnVG43ngBZCy
v5/1oc/foTIHod7ZbKAJeA0wwCdHFCJQP5EeDSHCXowot/ql33pZFRBF+QppQ+Wl
qfcy48SUY3uYhk6+/w6h7s2vfnq2LAfoBT1w3gJZ/ziQzBbqFHqzractmboHOhrC
lAOUdrypEkCj+IuDtVz70nhuWrtiu6dxFzwfOkU8b5vwQWan083f+hOfxSQEjhO8
xJLY6QTTgPVi37hImzJ3jne8g1XPKFrGmbyA2dWHMf6XClXtHPH6KvF9AQUI3MVh
KeKjjlHlctBJx7SADlclXyO0AwOpzRLd4XWuTuIFlOqXw4NNl3wxPbRadkb7e2Vh
WSEPCDBHDhWrp8AldR8uXch7pX8CXGHgujdbjjXjGSJ8scMUVJmUI78FVPQjImYo
kOlnJIhgS369zm7iWEdr9B9fSLTCFHxueRYda0BxPt9KRQgmWvyve38PzSrYXJKF
j0502mml4N3/5u6bYoHiiPz79v/8+TuD9D/kKlSU38pAbGx521zqkjXy7f0ngtG1
Nsbs8GR4bRtYtyi0jhaSJ6bX1Ax2yFtvQMpMLID36wT1ND1IdSZd7lFCgJn8FQ/4
sCo7ttLejatwHcJ2gdX9DDw/iJsYdjrSTBGD2Igd9JiaY2D17QSkBnV8vwH+1ijG
DanwYcydpwqXU4dc3X9CV0Rzs4Bo5zFIN6UezjKn7sutyD/hH2CQp87+8OnRQMVE
1EdVqezKbbYcs5648U15RTjBF/IzGcrHAVR+A0wm5U3Oj2nE8ZIJ1scBGI8VUNWa
6IYGWgPkEh3fmKPQp6FloT9F3KwIQ9grEWIhWXxJZkTX+C0JwkSI1G/ebv69LcmP
RTVR5mWz+nuKrfKmjeblZhM6WILKxNtfSiMTfC7V/XtBLVjfeNFWgRkUVFPxrEzU
Lll++Azj/yOJyxDkBdCkluJuA4sJgzQd7QdT9AiRqbOuGZdj7l8bCZRBG+zodIew
9Z1F8QjHCzSTaDYXRNMteA4l/A0AjBzN59dmF1/MhOYT8US3YP/ct+Y1V89U+vBH
FfiyIRJwN9875+jgk1Lasl6OpoF/jwN2rFKnPpWcjsfodtcaZLuRqINcH58NH9hU
rhp4/0XjdbABFRuhIjCZVGXcUYg6mI/Zkbtf5kPMDLzI1PxHmfDlLQdlHKXbcESl
yIlF8s63IchHBJUkcu9/O+YItQvtNh+xj8WvlCh8k6nMsTwBfeb7v9FsofDbOEr4
DYRXZhR4ta5R8RJAIW/Tm7M1JyG+x5MyzwaBczTVwVnY38YmB1MyD5bo4nzlN+xg
5kMKy3cIMn9YSDNvJG2ge7g/cI2NW/qL1I0mUN6BLhzfB3yQPHyHuEctNUwGo2ie
7lbXFcsQkzWx6TtJ7CvJgRQnkZi8kFcdv+ex69lvu8x3QAi78jGcqChHme3mS4iz
Q3dE8bzg998nG/9uxqQYS05DG4dqV0tlLCGPNw4SjUp5kQUnIFqZQxoJax7YK3O8
x54crj+p1AjrnSLSqr/5Fh/Rh1fnfojJgANc96Hc13zRG/F/vhlWt3K10c+xdJyU
p5ZzayoS9Acw4HBnoxe+dfx4rtyl7end4H20/bHVxhc0IdT3GnRycq8vtqRdOuU9
ZS2vSsnQQBHAZuyH3YlljMJApzq+kROLMBmU0yfgbYES67uCCq7fkNLIZA4nl6c+
H247TRHeYe/AnTQTQPruF3kra1g0jjS6H5DtGsvn8r0W9rUqmSD9KK4hq1yMnsVZ
0IhN9+H3pvwJwWMDwbzY5JYg4yrqP3dZjbhDldOdkWYwxfth9u+VYvjEfWQX0vhK
rrQypNTq52Myk9cRpncUcQ13n0XY6kUy8bgYA+DWQCgANzLOK3pkCLfV0S0a3Ouh
YnWOxTh2vT/7y30yPueuJ1kzE2HnYMJO+xgnw3Z1YLiFZlL00sEWL4xuryNyiyiW
oogEplOnMSBw6HNVWDwUQsBAIX/EgOTn+HDLuyWIKh5O6c4enEYrTYe9UhmvO/9R
fXZitJOTyTKvK7zviwCpxfyEopwDMzZNCrCuBRvt8FOOFvtRoS4kqB2fJfwYjg1n
heZL8hEdD9LiXPtLR0YsOljUHR64Dez9QW1gsfyVfi37zANncRoBa5Z0xbr1Uf3T
OgRTzh9PrvWCkGshgRRPovcp+slynLK0vUxQ6ircAX7LOmwwz2qDIWDpwVVvwCbj
x/gwEeFhranbhx/DnMgP/q9jCSmEWASif1CW3sr8fXTtOdGJuRLaQlNexMtQixO2
yr0dFbHN0pAT6QEsERqIxkygtvICtfdPx3t9iPJwSP6x0qAk5S14OHHxcgrUAKxO
sRVcLemSKiUTIUd4ii7ld05eOrkDdatC///j4Z6ONhudOWaDNmXp+Y4PYUIE84m1
9Rf2jsSHVkkuzOVkGCrOMWtQNKJbsOJVZSd2YllVVHHAt/MKUXzLFdOF/l/MflcS
ORgkRZaYgqHT9lyU5lYE8hR8hzng3UnfruLXZkB6xP8eRaXv2Pcr40sbyecyh4Si
igrr7W76ib/lh8XDV069xfr+niXt2YTT5r6ABS75eqWIWlZXfCvy38ejVuNd/lPA
YQzPb/eQR+WMKtnGO0NJHPUEoW+7gxFOoty+2A2vAyxJ/j3cfyFRqtYTtNWO9G77
w1qTw91RukldIRfpQ3WaP3XDIc/1O6oWVQDmEcgO5ImuAxEi0l7T0+EKt7kQFVle
SN8tDVhAtcIm1EmWnsXy4LQQSLC2tNRcFCwl3U8Bf4S/lfq9Tl3fBWjadrniIg77
BlfjOJYXrMQEONS/Z/TX2Xrb/8InBUBTbx4EyyYLbBpjWDZ4g/EYdG5REKTCEyVO
HV4hWtJNm827VR2wCdaTVNzgsnCuCvzMlmk3qiEUb07P/qEV+MmtaHxCAfzAZskV
efszDvm6aiujAC5viPeN2QI/EUHz6klJUuhHe7mqQdKl8zBzLt40tY+dQjM7DNP4
qUAyY9BdV6vXpj0z4EuJpvQeMR7wMBBQRdXHs7cYVQyO28ZloNga18Kns8CdM6ch
ePIicyCmy7w0i2lERKcJcQ6NCQ0RXNleBen4/eeto/XoYKALbxrzPhD8ANSojj6u
lSK1X9nOrPET2wv6wmV8Rzvzhgc+z6gHCkiubt3nX5Y43Un8QYJLROX3Ct9xLn65
IF0roS8w35a2DjOYvvoFFmyUSp+xs1l8VtkI8XS4KgFOUr/CMz/vFk/AzHTdxJFy
FaN+uKcYyZMrPsiSvfcCzc89V7wM3U8w/J1CMUsCCDl8wL+I+1HX0A3ZYLiVLePr
n1pacqpnfdgZd+vnrfq7ghRtil+LioexVnEQ4BVAK3BQXjkM5frrtKoCH+nMeKQa
8NYqZykQPbnv7YCIhDcTApOitXHEzTNuPOChJHvXtmFaiKbao+s8RkQxvjPN5kx4
5VHBUBOABojUQXhB+83eM3ZFzsO3F3+Hxhr1B4EKpgWvhSe3LJG7gCc7x1KYFVzO
8Hcz0YyGz/MIirSTtU5V6KXDede0ms87AX/hP9BiOE9Cyi+5bvGy+0e8pcqPEkld
/uzkmoYDZiBitGcFFzgFu8ffSLkgJB7uxHq1Kre5p7eXv5wwV7a/hKMLPjMmosd9
sGRcN4OC3Kl58BqgmiSjs784LTRZiAzTOiZbqZYxdwVZ4fn2PKOKqLfYFYhcNVRz
dWrRewzGjSIAEup4/tBs3PuYKNnEksZqBb5W6wQEEFF52XIKv6LijeoIV42gQ7H1
fx3qXhnu9Zk2r7DZsapNTP7UItUc31NCKl33szyab3bk+kzbuHhvRo5EkDYjrAMV
yTgVJplIMftGYYBKt1vZ/fdjf133ttM2EFeXJjRQ66jrwBDEby7R+2WR/y9qkntr
36Jx34D0GXtg1V4Y1dQomB6ud/HEey/vL4Re8PAtl5YwYoFyRSFESAk4e16Kd+U0
K8dbQYRfVEbv/tt4PMJBI8JFkC5DHmVty0xSKX6rXAi9k3lY3igWdhPMv3pxKdYW
4WXzzOXLl6D7Sv4hr3d8jpjjJFR3ZNLnPBMNPVAZiG2mLsYezs3MoEub1tZ4PDGe
ZhauE+rBt3iDpfLuJiIp3M6QIHiossnDUz63Y0PpcNyyah70bILv90QKOp7yC/As
OrYNwyBQ2rAHLX8ZtclEmYeK0tv+B0PdcxJcziQvO4nIq4QqggXafTf2fSnQuF2G
rsCvjtlMUcgxFZiA7AEaShVXvn2s0ZWqtK/o/lLm2nXBGfyS8elsSfBT/jjGjmo2
rFd3K3sZK8JVULq2CTEs6M/OwAJZGv+64t3QCGaZrTG47s5h3gGZM5AfFXBB7U4v
QDWno1uXXQESqiyLgKWnpA6EZec8buFMWHlBAmLexpoQcn6lj96Ntt7gg8Hpu7pN
MK2y0cSu+t2F0x3QzOsrJCmAugAWzSr/tvZ9Srdlh9K0bTEZWSEKpO+SVQii8lwE
QposZJ/Qkf1OzgoIFY/PigEvb2Rxcfz4tc3BRqwbeYWh/bKASQRQ7yLEQEdkOnLE
+a+oK6Zt6TSKspkxmr7Hl+49CDG2WTP/xkN5tyMoA4BjNKReCUXqqgmpfwODhQrp
I0JKXm2ZFx08TNCFGTwi5jrdYjt/0MRGoOGKNINemXLtK/q68GE8IAB4K+s+1/Hw
0UumuNmUI1me0f7svtxNF/RYnLTBoXlJRA+KgVQssiHB3BbYR5wRo/BI1peUv8Zu
mP1xoxfqeLM3h0xbI1W+f8ygs1h/CNFkfrJLObu9eCLu3xIZedQCP2Z3vwCMUilh
0Y8ieGPWLR7gqp6aUfU4W0qcmrVwcYN5IVGSBDiN3GOeCJHhXTxz9kQfFIFb2ZVY
DEhVjuWZ3NhZFVJp9++5fqD6FIlgGLCk++xMjm1ISZ0P2P29kMJ1ki/Jjr29osnK
gfvoj+F24NAr++wO+82nQ+8qo0Ifbo3E1l1CMqjl5RfFWo00XqOX3ZbRd9ZwuLcq
00vftFAlRZYeGbgPjohqX0NivZRLzUOMw0AknfrILKTgbdhM9RXvN26KRnvHxZLG
65EsyLDC3fXGP7islSCp/LWWemGumarBa6BbzmONwJP6L/FUb39bBAf6/DvAtj1H
x0jcqTn8CSLTs54/czuWnPemVu2zHtJc5zMtip2iKvMJNy3auNpP1xK6qsQit55Q
gRYxU0FfTLa40A0TqaUufQ72kJxJ6fBPsbOjfY9V1XY7zb9nKXo5GT/KVAXUc7kU
EiuNiyqeRHAbYj8F70wVWTaDVQM4j5afze5sgfRf2yKsNB/YdERbMFRbXLwrwsix
PPHJQhGIqPh9PksPMxCozmTrD4YdaKKyfAMR66D8kQhtaPkeKeTHzyVk5xPxxk42
1VTP0CPBYJLihiFaQsPJPUyjgqfdVSKw1XAksRQ0CM6c68VcNreFp99kjW0Ro21X
8AAqbSoE85KtkWohtC41+CKhfsvnu9oNEwCw1UY87qRYqldptI9gDpFs2x/O3CRB
ZS7kJQBrcu8toEOmr2cmPJ4AZgiycTei3FgjUfp2+sCpehMZ5POmb3FxXBC8M6ew
3z4yYkJP59BnKH47nx8zVl001INv2J4dmSFHywRIyJBcoB1MB2lf8RD+Y4HNNwKW
zL6AQuUow8RK1MAVQ4XSwkrTpTHS7MvhsKRYIcbz/kqjaPeC1kSQk77H7La1ZJzy
DwRcOfOZxr9pAXMn5Pf6SAaIyNKn4PUVhOQxA3P7ivzpRhPBgEXD1dyQOGd+a24n
xaUmcmqbGCbdSfqc/V5R00JLj4EQQ1/dbPc5ZIJ2O5B1VJmtgFD/rWF2RV4HqS/b
FHEeoagDw9+EJqoRbhZBen4Wp3OWKi01lL719ndkRJKg/mPHNypqLjgi0BRRpRsB
M+wZmvC8QJqFZJQr3XbE2ZSGCPNdkg4gjbE51hk9tPXDgf4WffHZ7I7/j6sKPeOh
db8z1sGlwrhm0VP/MNjGJfU45rzdx245EFTkIS32rgyms2whs4c2uxz+D84Nry6a
QlVnijWFypV7zKXOgsLzHluzh/IBnJVjaNwvjkvckQhCj1BfxkwpxO9r77EhWnvo
h0GE1cHECxUJbAb0epGmi51Vbc7o2NsqMFqJy3Ditlx8MFDzYbwK77/CbO8RIkYO
KGZcYAiZiGieWyU5VqB4HlhubzZyjWYkB2c0Nl+k+XhnWc5wkzvcZyikicXL1a+y
epM3I54fpmlacqooxYnYkZCwUxImlUhEGrYNpmWbolmQxnzDvDD7LNVO6NiIfvZy
gAfMZy8CadRrO2xuLLiokrbs8w2bHPfumAhU2fnyPkUEuAqlNZU1KcZpBzg/X0y0
qF5PosRL3ur/Se81oGbY81+V+00TJzRDgKkQ5AzdY/bHRmG4lEcF8PZHM1racHeC
A5FGdRetfDBC3l3ZyO1Qx5R9IbFpiKHeq5v51t/yiQNnJU1P5vV9vomDd6Pm4wz8
PweEw33NTJF+FE6tubXjw6umVAmESu7qt6eJ8bcXiTFXFM77XRuegtHJMeu4m4k1
S5fwNg9NXyAYNZ4sUbmvNLF9ITf+UtNByVdQmhrAlu6fXENTNtWAR/Hrli1q/14q
7VceFHs+56PAVgcCPprbbrIawatcuwZYsuzWH+qkkuEYKk91t94XqGfwhakfrvQW
IWiA+67AVqS3/3F30C+mFr31DBjhzT6VzH0wAZ6NUD1fRgvyT25aVyeJ2FV3VRKo
F43q8FqP8oEcfnLsWOjW7YY5/NaXJIsWx6r8WX8TG9hFRDiiG77im14niGXSP1n+
HQ6RAVC3ZsUzTyznDvq/vIv916PvV1LnqjYei73kjlY4uyGCMkVMeIVfu6ec3RyR
4Q37zaRH5CoCOFyLLRl9Hw==
`pragma protect end_protected
