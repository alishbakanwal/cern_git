// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:05:39 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
RNoGH8rh2/3uwEqMldaI+rwRHC88i9CT3c1ArSyKz2DytMf3LmMupuSUwKBXIhHH
Y508ve4btCu6c1yTuDeKPNxLTB5aNwqDo/5HmoRH0xRA59pK/y/fQGojcOQyulaZ
0VlA/+TQEVWZE6rnf0fBfaVMLeVdxRcHW1Hs4fOFqkU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 20176)
3sY8hxG6ObkAJbdN8cj+egnrg63/03TyI5v0Qr43mIB5auM0yRDel2cLUgGkmqao
NhvqPjsG2xpuXpxXzTbSXAeggQ2I54QxgZAYkTXPNQAcSHWQ7y+JMaPykhkMH8ze
nzvc+vBOYVh2YCPvqCnzgyPu6BYdZZtSvQHfy1pPJTXkB8UnWG+TZ3pFqTIFV59Y
qjZ5buMZC/JbM6PvyRiLZL8oscXHdVIHm1CGSy0W4EWca15WNx9ZapbWFCGqTSXC
L1EGUnmDPVnpbxtOrqpyo8OZQwR60kisF6ZZdvxb3over3oItZM7VtgXh6OfhMBa
Ym44aNFWqI2ZL0OiIYK+4l3AAP+gR8y5J9DvmpMWo0EOpqgOSGYQLIm9LvuYZMH7
aKXyykUhOE/QUxnhxygsSnu9zxfFd0FuQhOjqUuo/yirwuOMyuLvHRQBQ+144HE+
AGQC/xufLj14T4NTsbLEcNu2YfqqJQUKG44IKPGQU3jDqTMgOI8kpiWd29bvpI8y
zQRO/kwtdmhtl0cRkADDfviDftqA2UBHAKMKWjkJsSoj7oR/HDJmmUy/t7X38P+a
Dhghz0RoQWAO5DVMN9uAdHiG4sax4hw1XzQtdOwar70+61dn4s38IDi9xBOUgTgP
fY8HD7V66sOyPmlxESeLHcwjCSK+noMAw+IvQHpv8XQBKalRUyepKRgdXFTO+ecQ
n2vd+LHy9iq80MP8+Xw3FVP8NfeoSamhxZ2fwV3RF0BA9Ee/9CfHERcrnoa0NB9M
ik1FjyrJvO8eXwzgg3c/5PMXtjXMtZyJZOFuFfZ0uy5VzLPAz2Fv96KbXW5bzIPv
GlIXySS1tk6q9fO/R+d9YCV41kw4OOP7vAfxSOvVVXTVVlnGWl5lsg+sCwgzmCpt
kxd0nuOClGZ45wKN9noE5aYchYuWt8qP3dS84YfYXnYBU2jfX098pDh3PUcmdFLZ
DalsMqLB/TClN++6B6iaDyT9svxczBJukrfZXw3xEPMoxTL38jn+9ER39rX6mlUz
mdNk+YHXfzGkSzPF2bLBx1fXykmDKq0ya5bxKDkSNszHvps3kqCo8Ss49556llRH
/EwHrtLp0/nD9LS894kbFJicDlTsKEb+NLslU8iYFNa3zQio/h9KgnvkmZ6QOvnR
TfJEOu0F2iGFr0Ax+rie+T3sUEGz6OAgsJxHazuRDmTje3m+FMBYsuqbO4Lsm2XP
azHdcDv2967/DMX71+HwosjiUgvmqKDXCjemZTxrowQjnwEPgBsWDliKPD02yrEZ
CFQO7l5xMdTR9O2bq189A9g1sZJjxxXUg0GckYpG+x7z+h2C3gqWOVplvMnW0LhO
LFKUh8/WHjWrd7BszgemRzCrnH2g2RxWKjin+hJw718PMS9Od3QYMO8/FEAOotcB
K+r7gHXrqByHZDgytr+50WsotvfwrgX7OJIU0eRvH08/gLf92WCyqPemObg1LY2M
oL9IcYv6GFBnlfjOg0jSLp+fHis01ltJULanDQ8wGJ58LkbGI4aJoXSqTS8m4FMZ
rhlxRapJZqZ5h++tX9cCza0U3fHXJBLAWObY64LttBa8xUAEiXiSRB9VHNdBVpS2
/Jt3j1I8pzCi1/0f+lfSDvP4x3XHZpipnb3JyCjcnMi75HBVSFP7VJFrEM66YhZX
At+AK5NIzeT5NbL+vlnG+Etvpu+gMfelFC1RGvXpUJBxisCbiEzeZnu0wDy+Ls8H
Ymj0yuBwxnS6q/Hy/X7XZO2GKdN6c9sXmhvFKmKaYaw6jujoP+0QjSbkyiH8xlBK
WWmHMeE2WRoI6hOxGWqcxjU7h8RsyN54vNmrdQUhTcGP/wEzbNiC6manFVqcippn
ltTPdwZ8ZOl8/JE2QkUYWIhPrP6bsCvrPt09FN9RzsdHFvx4hv2/8b3J1L9Kh3pR
Yrw1h25U6Pse1xnsBr6SKpFB/wBaC29y0mtg7swK33lUk5qD31wu/0F9aNzGSkOl
tvod2t5e35WWJdXkOUo40MNAinEIpPzkiFfPcW171cE0Mlg591mIlmhBKQeRA9EJ
ofws886NOOdhx/o7l6v2VQLAm4rO9/H9v0FKVkk2slbzhAKlwdDT8jzi/eXy7QJe
LoLIbyCsmOY/vds6O4PtplGn8SpDRpNq72DZH7lh7IPmkyRm7pwylAD5Gj8V7+P4
S7TwWNv/V+16a/U6MC+TEXmHzDV5lnnneZYaUDtUFOfc5t3Ucev8zzugV4pLUgPM
Go/PR1L+aM2Rr2ovjkE9AvEAVyuypFvH9WYZHzHlSsXAGXvyYkwsG4Ka0HVLhQp0
lJWppSzkOLGby/XQ7Li+wlHFoAtRJdzsIfdwJ9csyYGsXKI9Vp+3AQzFNu2aNSCg
1kevhI+hDk41VKCcTE9Q8aj3c8TgvpbsVIb6ztzjULWrShvuE9OR9BSRIBlBW4Ul
mKMPVDugYkONE0PtE/pWf5UQQUM31nMJZG1EWM/GJnbaE87l464TRH3x/QOG8Ww5
j9UATRV04ljIhQ6k+knZpJ6uv+6MBVy2G5p6kQRNvNHJK2fxgRtXY4Ac7Q1Mq0y1
Hh011d58hgYr99B15jAZwstVOVh6PThN7QWHQsNuKFQvkzyS2jFNnF4kiMgKvM+Q
TVOwRMw1KpaV6Zy0lYrkjFZUenFGOh1TJ0RJm3fD/c7+P5Rv8+KPdi4uRKvvMwj6
IDksjY3TbkiJdg05zZqq6yl2zOXfpjhLQFGuHZhJV5nMH8M1d8vH0h0gZ14sB7kt
G2GPHyFF37Io0bZnoJ3LlwxU2RSM+GCMIPy2hIQQ8bGjVUFdxAQhlgluP0trte5e
QupoILn0ngBjnXdpIdtXaOTT2b+XCSDgVloARuVKFppwMh9eF0jzR0qj88X9UcE3
WLQ5ObDz0pqQffqDM0ACIvHCSp2Ty4nSZ5Ui3HRbgrkXYIpVKIGBGdVZRhjfQYcD
m6DyN+v8pQnb6ydkIWhBuK2TCNeOg4O61Rg1WLcUMzpARN8IJ+PMPB3IVM/h5HAs
n60WeI4P+/Rlag60TT1oEEkrV6lHcNmV8KZFofVhXOC5cQycE1loPveaqrgJ3dHf
RdMcYXa3kGaoCni04RcupOBsksnWYHdScBDrlUnker4A5riRALn4LfzR8cgvlmfN
P/5dtm/y5kDPf3kWtotc+p+NgaVEH2Z7/28EUhBvxoydDdvhf/2RuExo2hDyRmB6
yYZFhsDb3apS0NQz4Og7mLtfu9Ub4LslwGp6UFBrthH5woCC7iMjvwK/EiwVoM06
m8NmZrq9gzbmglhCZvmxjsHj5TzSghgPT+ZAQ6DpHc+UpuCjuxg/v6M9AukCIpfE
Ruiz25HzVLRuklzjeulgL0ZLFzcvO0CPGFXtduNPh8LD/M/8WPACrudVX2lDh4LT
rvreZRlxVbSbcpbqD4IME7EbJ3n3iI6xxNJFNVouX45+/71nyQrGUEStwp0xVpCD
uoUbpAPcHy7vAlM0so8lrw+9RUXnMQHDfJPNTZ9H1uHAw4ny/3KCL9fEpNUiOPq3
M8ZIIeUPS7RCcoh98P2tqIzber+nzi4mpjVTBWQCsqCv9re9/qAQ2+NOYtqV3YOS
sc2bPqb0Juysyull3kS4ElYKwDSqrH0WpPK/yhOji30UD4k/oM1r1hdyzyR9nATh
P9cRNciSNcDo9yiMYKpReufs34W2YBpFdoaHs8UPcZDAY7ylN74DUkap+OVPZdQX
7vrjDlO7ypf7/LAdump5jAmwMbLbsjTwLAMgCGLzX8FlR3+1EoEIgzmxQ+AMVgBg
Et6YuiHZ8VrHoTnxvj9BKobmrEVEU5R/sX/CSR5XWl2sypYHS39mScyDrQcAciQI
3ifGPMkmG594MAAZYVyJhP4xlhOHmdbjiTzf7yUAls9EwA8i9L1hAeda2/WFSxmX
ESn1q156pTqlIIafQPM/TNXbBQ5xdSwBAqYYNxkDRkmMGuRGkRgm9eIH/tQVkyv2
zDsdRqe/qUeaI8BuovkUFpAV1EteTPTrMd5lHu5pOkUoL+frCJFde7kq1uJqkSeH
1HHku8aR/ojFy6f0zRB67sXQM69eJb6rZKNfqvyMf/JHNPAbjySboAnx1Jef8Q3A
gUq18ZEaNC/vHAjLBDIOG53SyUdKfHF99ctdnNBftbQidE4pC6UOYMK9R+t9UNmc
77lKMF0TfmP6i6Ng/ABMkKA2fAU94aCyyj24/VBaBRM8z8M60i+39BoJROftAhPG
lOUkYpPfeYwSpmRrCzYuXx2dw163lpY4PjC2LU2UixPRS3pWe8M+9LSaecvF+QsS
XvKjF1ZK3rSE+rs+8/twhR/MU/LLWgB1widdsBbPdQFoxcrveZ9EKvOl9jUa1A9L
yKV/HEJqbtE7WRnRN+6erR5FsG8BaIcxspDAtfzChosk+tks6z1+KhdAKO8+zNnE
wrpjW1qD5zVqrlrRnOasWgkoCqYtPqVGGxrheXdYjUGK1wWfrP6IJLGkTtGZKkuV
2hbbhcyEfAhT2QOp3/QAx3ln5SeEqbHtXBDefsalzq57RaIoauZt+xnyruB3F6/p
wZV8yXAQUKC3Rl+6VB0wBu0ANfmSiDq51VBbxxYipyH1kmWOVIRCdgaZXy6TK8ug
y3FeZuld7cR3+lKHe9V/lhONl+i+1jKjoK1QzpajeXe+Rjc8xKUwSCkELuy3XRye
bUeElEJxcj36GPcsLtlG4VCWXNcgm0MJO3ZjbN/M7s4Hc/pm9XUyRnjg4xSokdZW
JERXEQImIY+1q8OnrZ+mkY7Qy83xMV7RFZ3894UugLJv6E/e2+/om4BpUuQxHmxY
TSZww9V9HVs/HELAy8INBW5XhNTB+x6a9VEmM0GA9PrhywquuhGdGrfSSD8xvOZw
QEE1bL9d0AZxb9NueW3NIl2u/DqYS5g2+BsaMyyrmI3ce1JGlFAOV8YqL+baDHWS
J57cSU5y87ZuPuoPbo8SeIH+VHVMPOfx755qBiRD8EFD6xYToD8VJUTF02tGgJMV
5ZmgLPcoWXmm+9ECw6UoRxESqnQEcjtKNPphrOG0zIBvvwBl/J8Kkk7lbcCAaiAK
TPg2HNVs8C48vNTC/2aGtAb9iQOv6fAML/TeUwQkR3eZZXHP5fqtg3Qnc5V1P4+y
EmoEJu83yRD7fIcrSdj1TSNsmLLJWjjfrYO+nK8yxYLdTOLXLCqXQT0dKAH7P8MF
bakwZmeDDpDALQB9L011Aq2bCLVMJ6KCkK8+XcuTrGfzzJfqW8nk69qeaM2SrvWc
Y3XkEn9rIN/rkXzcZKVIDA1ohDrVhEzHNudthJHzrRoKxoCa+BbSU0QRgcZDU7Yr
IGmG1BYqHNIndVs01teavHFVqDxSz8VDEYuQIJ3hhprxSRNbdAh8WXu+assHN1bM
1G3x4tSQmGlksQHtm3r1HLO7RdV/VdMRz/4ODMKUN+mvJ8irt9rEU9adwutcqeiK
onl8xNJQSV/P7y4kNzjRDgZzNp12HGdOCwNIPvFwMAbKUeugvNzSnXfIDEQwlrkf
A1CIxjm7HNL4865h++B6xQY6n07ep7oDxfAKl785I4RIAkNdbrC5HZPIBjNd+hWJ
RIp1o0g1kv8eowoAcU0QxXMvZ0b/5A8J55RwtjvuNEjrCltIuMbWivJPS31LCR+w
QAupd1gD8PAsQ5aslZ1PTKaNm2oCNCd4kiImM0T6kFxUnWdpYumLfKkeEa+UWVKv
erAyoymEcJkyADcYjzI+89VqrulgOVcEoYroFvogVjdU5cNpBbVnSY7ejxgjgGpZ
v2KOewy0+jiKXtHUG3T58fIXaNFX9nAtlP8YYSLH5VENYxt0onrHzI66bdw5ScfW
SRF9zO14UdgP8fQSAN7p0eKB1cfBYCHxaP7kl9Mmyog3WrCJobTpvLAGonHDPyHa
kBDYULDgFlLxTIYyAwHjMj/77x8s8wm04d/W5ki6YZZmxKlIJ6982fvtwm4+dkhD
4lrJ3Odhexi/xYMLCENOczvjJnAqUKFe3Qc5fwZPcndSqWj+cbAPUwXFMLpLOPpo
mqkSLmYsZxlscU0Maaw4Ux9Tp77RtkKgItLOyeLQyCj/gQ7dS3GCAcFq4gZkbyEr
D/7xsLLwbj8zNVSYjEcXugnc4fNm3YzLGPKAlQOayZNRtoeWWnetob67JXv7u7Zv
lvtSpmEUuODzJ/mqP58sqZyNxPWm8YNDF1LIi1xPbAwx/hJabahljzq9dMa8ogQE
aIaULpGPeVMyBa30Y+FjsvwEgFZgqTAn+E6UtisC20/3eH+tI3KTECRDBFhEXR8g
Tt2S3dFg6mr6Ip2k1XYAH4yoe4LgR3Y133CvpywswMdPDmJvhYKY1GbNhy+CE4fL
iZaJbgErhO/w40tfBfhXB4zCYeBr6U3bpdt85tqDrabbH67zCdPNDpnGK5MTphRc
dTdGwUrDglHqCsVg8fnNNzVIkZkJoZy2mJTlWvEYe2xCy53Rmh7YsruJUoz+obFc
gqgjXdoRDfEkEND4By0OGrby6Xyvct0x510i4EWOfaFsdgFgIUgAOZa/ptY5omJD
Xmte048v7mEG9j4S9/5fD4IkD8kR925eH/gM1VFloRqYEQBgHPtRnmyC5O1Y7ajh
nf+tvR+9ky6A/l5sGwVvOtyD5T3oDNVNDb4b9RHPwiQ4C4l2nembN5KdiTvV5R/e
IYJtc5n+Ir/kp1bTtRHjbwEEoKOQ5KgClq6je6l6IR7TxoielLXP10fsHqG6Vj1Z
ygUHWgHBug9B30by55sRzrZd0tFDxMwcZ02q18deny250crh3YgpOZclwYsh3rGO
7/npXitvPQlfe9o4HUtqo3zkCmBDsge8t3UaJwwz8/M4Jyo5fTJegy0NHhaAtLOj
rIg8lyL6U0mtaD97iZYK3aOknCGpFsd0sQG3nefHxSeA3Zbtqje0iOWN9WwTfPA3
zNwvt1GfOFtu1S0DUxvsvi49elvjJwtNRz1HDXdFW3LwXEGaxNf6vASHQJOvgWyu
S+kDdfRTJvb39Cve4CZ3XfIgRi3DFd5uB0UgsM7aYGl7hTiDrIOFpRiG0g5BcdbH
58Yvia/QTVG9lQDpxxv2o3P4A1zATcbxmtnhA7QEqX2yWACfROlJ1H0YXJ9GdCRc
lBI8KS3NB7RYht+mv6mMdgk3QOqOfBIZeJ/D2ehY8N8bsxk4JXJmvKjJhvfrvLGw
jFsAHEpqSz+EnvxZYNGcwicNRQIjQPQjWfoEUbFgnxcnmF3WqKNW/twWyQEGed4o
dvTQdbkxJwA9X6ec1SWsj+IqKxgFnHrbqP4uR7zBEJpW/rOakUYszHieycUAabAV
l9coC9CZc7rscGSxXP8bIhJVcnFnLrU7Kr5+Ux/w/EHL9B0HNzlQnjF6Cq2RUeT6
jjhTvleInEmXqcG2es7hJPHxnzpTOjg9PviYWdghNaixvArs47SSZkpD5+d21mpe
MvPx1+9ckJU0pfgCwYJPlUQbHbKkz/LmW1xo4EQ15YsS5H/QkoIgaZ1BLIc0D3Jy
W8OgCPnDMtAZ4BGiJrVqF+j4+VBlKrnouAUgWD04ziIQybZuCwf9ytS2nWBhkxvi
7oV3GiYgdGADeGzZKnN49Wo1N93n3/Z+i5Hs5EW04BGBsPWKGFQWwdF7HCz5ksBM
vuKY0baTo9Y3eENJy8anPi+8h4OWzrti6RWq/5gyLFIdllIPZAWRH31HicoXW7o3
YZ9jwgZgPlDQpmorVC53JPZaXd78Zuq4T3cp210AYsfkTO6ZRq3U8Dgylh6OdUtf
0x73AzIeBhOYGBeonz8TlawcnuyQabvDuBLpsKRsASe0saFy7XkVOSVosW4Z7dHr
Zg1lWKIBBWSVGFEYVGx1TgtW6A0S7FfOuqJhqigCAPDE6eMgBFHu5zsKOdgD3wXl
IgabgpZG1vSWL3yaTSrkV/ziEKYtmNkk5Uk/ohSt1g8VGNvNS5ICQPBqZOXxvaFp
1LppBxCU8JuriBqtEGin+/L7F9F7rhO8FU+XcPzTfpfdYCy6nCLLuX2SbjYMUfLq
PLVcMdZdye097uCXbf8Y+HKY5AxJQJxq9LB1eFm8CZA6LZpi5CoFzlJ5YzOAlmob
wboJZEDwTchrNSH5e3yb4he7hnR86PSZGR9WxEW/caF1YY8q+ldT05FZ0KkT//Jf
5EL31/ODru9q5nuAqfbZD2sfSbw1M1kYDsgnb0Obl6kMJC+zxYZ8UcYm7M700oxT
F8soojYyjalsAMNOVmo21p1njaAg/VWs2sXDQEFA6/WoNjpxQzImQy8IV7vuy+4t
c9CrIWCsFpuja91CA7ko+qY+2yAvxwsvmapKSAMRikvv7YzDTm8J8jC/TZ6rPBNg
L88JAp7QFZxTblgIHlyQAbigp6RzT4tOUIof+O0tNd3tGRRiaZmjvZQQYNNSx1hT
HRHuZeLPN1kutq9ZinFtcfF9UA/lfQEwnVNRb+q03EZ1N3tZ0hT7TC3MA9qA0wAI
Wp/cEVavNZpTphch3piAuCCG+yQyY77s1rGX0a92xCWSZvYPfB+rW60ZMI2KgGxC
UNDidNbdashiDKyugH9r8wYvOHl6TCGOPMP9U0H3TLqc45kq26+925sX07gfpc3C
8xe/cJ/BC+0Qez3bayHidsbkfSXgXS2Qa0HE+KDRJprCB5o5hViWI11xOYa3LSBT
zes72kmEUIhmysht8vk7Hyu/09THdZNUbWvIvqmI2wI03xS/3rGdhxNSq6v+1y5n
niSoAdmaRK9xFXXA2NWIw6MiZWwsK7RNIQDWNo/8y38jqn6AQi1oy5ugqycIsw73
XIBp4RuDIMnLuligFYGmcCGvZvDOEn9y61BTzKQl4jbs/RhgHPgstd01UDDarYSv
Ia1JeqW1MsGhXuhvRxpb8/s222Tm6PljNyIDN0/CFbNXnfSochOEr9OYwUm+rChN
C5kELy+Ij4quBaxG3Fauxupyidny4sUVe2KuKDekTi4OBysA+YlutXdLNOu8/K1s
n7T4+nlv2MoUARKXCZMftEF47TlIDHevq/D/p6O2TxSWjyGxPkiW1TTIHL6ur3V8
c6rro/RtAqcVXS2ovj42GUkT30b9k/qQrbUIWpgWleVgfBkMuImHmQ2AHIr6lxqR
ugd2PHN8pukGtWtw59Oe29K6rfLZqSJiUR/TnpwyHdxBGiRCdqP72mewbHuUelaW
K/ZnAGENqtPRN2gMamhnPxQC+buszF85ocMTm0j0iox/BZueoXm4ZIR73WoIvHmM
ryXGFBrPtX71kpuxjHHasSWbnGmvlfzs/8/WGy5TtgHBG7b361l5wVvGDlU2+KSa
1JiT8STB0xmw4vAqWUdqAvkLYjJ93lZXjqdWexH/zDraXqPhvkXQg4RoUEI4b5Nt
zOUX9Mqfru1yHRApq0k6P8fsCXbt/Anebn8bFDo0psaO2v1QMRUViJ6x6TprZuQg
YshiqjnEr/lpdTEbQwd8k8Hid+i45ISGV0rfAsy44YmE/YF18aLSMl2fQ8xoArHH
kwJ/00gvNrSjlDR6Fbqvc80dGcESz++5Y+guS40xjvjrBmj2pxWJXEf3mgy2TDCt
UyLkSMAHrf8LyO95f3PeASxaZIUFduYr3y+tgjKbBQIH5KYnxGMIQvGAP7JHQios
U7UoH4kU+yylPCabCT47oaYozghB1e8OCJ+bwTYJwW+I8ks5xByesqtLOYiRgYfu
YAYKR8HYTtRzuGrDqv45eubSF5dPqJd2xG3EL8sCvNK0h5oKOkROJRaQhKQnBRAT
JOzE8R0Chnx6oiAEHayJcuYMBVYEoAV/T8G63vQJSg/sXSqwRUvzf2X9w5ri6fdM
/UXDY2XMbmlzOGU1KwqQ9oLmfi+FN9vyRsercGSNWjRqorn0t2a7oRijPxrx2pae
5EZ6EoGWW0sdU5vuFLqjMrap5xiTWhTHnwaEvJJBm31Bq2CHZIdlSoXf4b22uR//
wLUqlzJEKMKbrCfeHQaPy41mmZ4THUE/H/7UR15ugf/gCseRte507vIdF+NCxhZN
NKXd16xh3jEI47ZHdmD2Y8vbccWxvwk0AFnV8nusZ5QJCbDBB7uXVblHGMGvkqrx
m/rnf2WRZjwDY2iIst3FE65y1c8tAdYk4eS0Mh6xz5l2kCNM6JKcJgsF7OkUcRZ/
DE5qzafYm5MRiQF7aQu63iCJeBmX07eMdIGul6aU3qn8szo13/cpNVXzNWzmRyJf
zzpKdiIEswxFWoQNE/cXJ2OdBa84Lh4GQWPgxYdjz0Dr+mVsvuiRMe4DhcewDNet
fNhl4gc7Il0BZ4k1CX0EthPqWvu2F5GvoFscNKAcDBy9y8pjwwlXga9jq9tujgMb
ixTWlna8pgkQa4gjVMJqXMnuYMItAiFNnhJ9E8sa0Ijp+AtosfNtzxo8PWqkGe8E
I+k4zS0OOkqcHDkICOTAfcw9tfuB6u2nbDhedbCcyNxNG1EjEkVMhRxwy31TJBTP
JRqWf0wBRFFGMPGkWL32HV6doId3YuUEIFCdZ8DYuEE+JtefZWN8qHqzOHsbtWwG
nkBAosr6Di7/Wkd2fG2Hrw2wK5DoHLU6St3eOtF5CpDm0390irnlQk4vJhfxDBo1
sCk+4TTfsINa6Kxt3+giajk8yDPxy9EGFS92VvFuwoh3E+0uMCj/chW6K+DEr3Vc
2mCX6ajy8Kg2Y9RJr8lDajBwU35zqE3/KFjTvFi93iiEUCudoSkZkHABs8SXWqOE
uQnij6U8cZcnPbbpgEitEFJydEMM6VKUJmR//QLxhiKOid4TMKS5Dv5cGsNm0kiz
9TY/gsZxSE/wcRLCzVO3GAExjrraQH9SNQ03zRa+tUWhXgAsUvcrG7Mg8KoEUaOE
z5I8YjfiRadrd5Z8yM6J7EMIOY7pl+ahX0IrHV+GWFZmRIV89ZW3PI5GbemgDfYS
po95DokrH8747JU2D+MZaiS/d6kfVzO+vJE6Zz0JyqhgEQfgyB8sUju2QcrzQF9H
8qU3k1XDsRJo1oXtgi6h/zGPF/S7PtBFqGEd8MUERXzHYraJJM9bWuLpy8FRNYhY
SBoCNQ3MeaYsY0ABoXeNM2xOtw3ct0vm0FPopcw/LcOhLxM8nArtbIUjVZS9cFVq
BWgS5xxdd2GBGsDwnQspKdDDw5Fs8Vw0n950MLQvJelPcMVTGTTLplxbJt6/w3Jl
N5kIkieZhQuEEyCLOpbPkoO973856g4gmIwx55H+YRTbRa+gDSVPqArsW2QG9CWU
8L7T/h3b8sO9pbTLkuR2YXc+KkqsAEoLr0RowbvD2t60q8dyrCqy7tdgQg78OjZ5
BsZBuy7PcUBX71ITOWc3VK/ShTLeO174/sfVgOparGFpvsAcTNP9TXS5Uh2+rmyM
223jI8iGOx0DaRVZ38oggzj+svV0EKv7fBKhMwS9ryXeFWTnfRRMGzMeQ5EaHS7+
g2JJGt3dHqAsAlxGU/WyBRSKnjHoYvRIe+YrGIzrzb1C8W3JFebSq6sQHRiQlsoa
7sHsZ7gHhTaJewDtXo1arw6XHOG+AxsRKZBaXmPUNiSVy0fRgA6CvI28otRSYjmI
+eZuIgNgeJbIp6p9DkRRjI0/XNm9lR220vR7uyvoNAsTEv86YDEnn+nrPa88jlvB
QAC9xIDMULYe77/8eBcBXXN6JmNYvC2ruLgarTitbhuI9J5ZoFdpKwFR3zZIKK6y
/xWt2byD5OSKf0UR8Btz4kY5VNw/swN4Bl/g8eNDoYti1OAr4N/5rX+9t5XG+oMl
9dJg7h2Kph4qyVhX8NdjseA4oMsD/t5z/OlG/tPsymznxO3XmazagbR/E1i2bf9S
LIvNb7k2Ixcg56Pp6YOfHzqPGdoCeLuj2rvLeW5KvmSAdAodoYTlL0DQdC2N+yuw
RIVdTYg5J3afzNwKg2lo0qU6rlUylZZY0vJY/71mCjiWwSJhqqu7q5xvXMeqrvtE
WkD9j3G3qM0tPP7d6lduhjKUsUkcEFgqgNQE8jfSyEwpSbtQYCD8gK5WaYN+hy0W
191QfyylCKTGezQlNtATv03no6icQlfqdbwGFjfaBvIhnNSW0BXmepxImRUf4hk9
GWjhgxsRjTabMPxwvbpHpXwSW/ubgKfXyVamDeKtNKbm1ZEKQkT6eroHeCR+zrN/
MdoocvajMqd/BSLVfe6n5ci938tEKJjvZUJxTlp6iYWnz5btwdr0V7JtqtqsuZMp
HeLMyvMm457z8AS9vk4o8McpxHPzPCvG6UsiHGVqijmV/8IC7Ok4X06HygtDsmTh
XXzy/Rnls6gVEHLvqdBbBA08EoM7pUj7Fnva1sd2netIBzUyfxMBLVkRNCLsgY89
NIuQTPjTlXZRImnMVX3w08OgBxOeZMsme9ZiG5UxDaopbZkFA2zUc0Q/a+8Fp04d
0pwS47sZK3QV9totqMtN1mGR9OsjGZsGJCkSy2ScbZqxTZO5SMuVkEfpuJtCPX0f
HsZrSH7ZKQNzhh2KvLcuhG0Yyc3000MlsDEKcrE0+Xarpp0RzPwxW4peo85Nl+Yk
IinxCki58J/khV5lcplZ7o7UFD+8o6KkebUFAhmRAsAamQWapbuSarKQdgqkeTto
R6RbmWkzubR/VjB9eWomQIN+4NZ7t9gZfY2NEKPypdGz5fhrCjBDXV/FJSarOXSn
uxbDQsieuPCGyP1Saz66IlNA0R0RTEc5uitPF5NbwqAL8ddg19vaaYToXcVY/rFT
U3aqnt7nnsZUeNXoC4XU3Bhk40SQmRim+DugEOHjE3V/ulmoC15BaMdtdmMcDhtX
5DupYRg+rzwILvJpBc71dshlfg6R/00dlrgy40M4yoBSvdWECmPC+VjvOSlnuLtZ
smWSTjrXUoraAC/ozv1R0mnnj6nyrNMubyBIAqqm1H4pBSDfaczzkVzq1v+eDzdF
/algnrP2kcXitYE64UMPJIJLsPBw79SoF48fhkUENfziQv56i0bWOwEirXNTA/58
Ijdoe7UrJHLyOamJn5KxPxZ/1gk4ANNkuZTUrT5L0pQByq7xQxVxRlk4BCAHXqWV
r6NouYmz06swfBkMi8SaNgxfW1wPuhdY/7pH38xzmJHIj7uq267RUhLkh2EQUgwp
XeZyeP6iylx9Vv+cFlv4dzElTSjvlD9E+SeAa+zs6+0teN4I9VTyy4XF2w2tQlot
DBcbbHBCX392lxIxiwor9gHpdjSh5k5N79oU9XOZstiqCeLIBCjFR3bggA22q8nX
RCAZs/zudD3VgLRiIbmudOHH5jmTfzMuAjg9hKtIhwumnlIs+/5aklF8fsy1JZiC
YyqO1XC0lV0VpFa2XCh6GJ7r4Vex3VFh0afBMfVvm6a8Zd/7/JqH4yBcQHjf/+oN
6t8ymlv5+9cuq/BG4Ep9AZgCwcoThmxYzIUNWvhnSp+LU00tPW1mpL/dQkBhHrtm
FwsYxdbF0dWrBZVQuhAdP7TDBuwpDvHQrfoDN2y0gOLQB5QJiy0soareXlNmWwcH
B3e14nBM3bZ6wR2Lnq9mwuv8zrpZEpMuKoDbir/RJUf1ZXbWR8WJq00JP9W7NJdY
2url/WWTjLwG6kGlH/v8fe9j4L5Vm8N0ylRYcPb3f+obOLDmLxP0hI/RvL5nrIz4
Dw1+XwaFMQ6zX+zJHID9W+T92GoO4reqSKV9VOIIIdbkvmXDJ9yW2msZLYptoOlA
pMpIQ5sabfa80PXZcSDoi6leaFwX+IlVlu55i8SAzbCMgkrybX7W5MBsIXgnFFZh
zzOtis+xxuuWo/vU8bdc+NOMdRPM56ef+FsZEWbudpPe9CEOW7MKRGH4PMtZ8Pkx
oR8oLzZtdXoWLNwAtZ4coIivK66z5NQSXNKefB014j/cU5PQqPEpKSnpM0xm91NB
uAvzJ6C1acUFnivSTI5mVb8756gDTYzqLh9jp85CXLfI9Ke1FB4sNHO0oWFjwqHI
hepCPQZspn7gRnX+TWUDo1AMw5+lrUDvE0GOb/5hTzauQNH/UofYLwT6TqbDhEmS
qCsKV/iYxCspYtey7619GOMdHjeHZ00G8zwzOyz+qj9zcn9lersjFvI06xMflPIH
cNHL4k2tEDWiToXt0iCXfR+x4TEg6djqjf3TKxPyX/0+zhNvmVmyccG5oAFlcuAT
MrO793PNCQnDNChYw8smo1aD5ED4f5z5gGl2Hxcb2A5izAgrjavTzfK799LqJ11T
GjEmXm/U4a+qXjNxTQNE/niCt5f1QiaVP4vDwGA8aoI+xE/GD4UxHk/Y8WAK5mJR
/lBK70cJqjqi+U46IY8CmTU6iyczie3dprkZl1xu0q/2UrQX+vXy2Ksuec6JOXmj
FuZgnS8mBV4nGbJRS7Nzs+vVyccJfr7WlOYxBoGikKsj1jnwAz6nEHcup2jbHmsL
ODiYEtITcRkrjqDeFnhkHPCVOWXcaVP52hDEU7GzdvAJez/zO7hzNIzxRt1wSYqv
7eFCaur8xN8YMEzh3zVyqLklZf4twC82lZt3LvfwAUsGoEG7rSMdFzE8TmK7G30i
U4NgiEfMGfEqjrfM2vggVkTUydLX1HGNLMxl6oaQqWeWnQpxXicxrzgvGZdxZOr3
w408LNI2KeXPPEf+KHfkBuznd5XxcFxNlBcfJHdXNZAJm8WFcYzyF/aqmHb4xiAP
tbsuPML2xirvkTWQcPEc5DHjVkBsu2cp20nLxRqGlpCcN3TTEXp/2IT7q/CRc6mJ
gIE4K7tm69vurVrrIuRLFZqocrVMHsw5uFRou3EYKO/PpReIT1UzWAyGZ1iZx2Fq
DgSkL+FQ5qn5Bk4b9CHpT/VVMGFbJtACSSHAERg8U+kPqMkiDeHo4aI8XkyAOGSf
mJgC+TrzkcSW2vVH8zXUFh8lXvdvEHRwVNP01pLhgjzwbuO9Ul3C1Xq1+nSa4o60
QKpfp4i2R8FI6zI/QKM4c1qyH37br269sj3/6cjsJX0+5/2cKpkfWZQ2o8G6G+mI
VoeyXElMQTHfL4wRVEoLCtDbaEmHv/TeAYpNZ8HQs9XMCSO05DAkNW1n70uXsCtP
WoH00f3i9svSL5r+297629XLHAMg101uQTnhVsxk2Au0p80/XKFgBa5BSfzrwKN4
SVcEApqFkSn07lwVDjZjR/OJZqGxT+btdkgMs1DTSamR/Ex31KlREhvqylQ5Dlak
VL1H97+ma+MIGQo0fUAhdftg7bOSl0G3OK/Op4oGGmyFptfVER/dwMneUFYA9kuh
GrosoiwbaFKcEafa5P+ykOvK5HC6BLUmDDmAoTMQiLnmjx/hVjwfrzmS+M7Xi+gp
g0qwcnkCfeswthgdBcQo1nMzyym09xhf9O7/ZiLcUPN1B80rAdkkSvqLyLP5E+9f
gLCYSx/sdWLeYOl6nOh7TAvUQlCkLbS6lJ3HHX3WFQTM1zJRpMUyjMHxQtY7oQoX
/3AlFY+WyOSR6cBJ3YbBdkwk6QemGN0s0oxRI2MuzTma0lvHUemlBshbe0dD/cfb
d54GkKNMGoAYjOMKXlRTDtCUCNVDruI/48DacO6+NwtYbzKYa8RkBnU2ARSW7mBs
io9MvKoZwYEfsEMvTRsu1YSMv9UDHINSSfJ9jJ8l27sH0DnOo95GpIEcXVs14jJu
NPWDtW5hImEhDukCV7c26o4rQQUiwN1x6p0ECHl8eK87ZGt6FWWzBFOWdy4ZwWX3
0rTJCleZwvr3uf1qQfNfqA2UXzS0DLxrbaTrJqUb8BPitkeE24c2rjPbeBHtRvX+
oe5GfQYxksii7osmo85nkjhzcWfux/RUWLP7TNitT7mN37JJ7zLGc/smbL9tXdVH
hZExOu9jW3mYw0KF37HAllxAfZavMtDZVovAKZp9VZztIFUznzFcxATuqf5ZCliT
fvTohQ04w2Lj/QR4MGu6hPBZtKAZDq88AeeAiyAZZj086jVn8Dfid1MzbDP/dmOg
AfYNfBFzscLe7fCmuTzzUazBkApx1xLmajP4COpu28zKNC2+kVjfXuIJ3Mg/EHlZ
GLLBeqPeyLF27YNCM42Ooh5nmnWbp64R45Nr1LPdnk0D2qoWI2oe0zzBK26vR4hG
J6khNdJIbZcwjqntJqnsRIX/LGXWIInWbpCmF2urOvxLA3T7NK7PPWqDng7fyqIH
S4DIVeIxfRYz61HC9VgKfPBdM1oE2Su/+4duNzG0rGphrKSrJlCwoCAAWOHJyZPb
nM3FYlZVTG641yDuE0000zLoymfxuim13qbGijMY8hkrQ9/0wLJJ32zx9uW58o7U
LDhoJLz37b7ReM9mwD42Vy9YI23PqptDvHuf5gn5IM1TWhBXO5G+Thdi2jkBvX2N
bRhsgfVRrANhMYm/qitY6KqkH9dkooftelGcAk/uAo/yGRaJKtQS/vOHL2FZLt7X
89AKDEy3bnd3m9Pw0v1KG5SdrYGGWF1vazuzlPTG5whhF59mP8fq5KNGcb3nbHSZ
iF8G/Uh+ohhv7zjSkXsqGsESETde94nC1W/j4U+Ukq2vS9hwu38NyG6yk/o04QX+
Kv+uMPXeIuNgnpTI+5iLra1XKXLVQ/G/alSkk/rVjPNd61LqxBOX/1ofDMLTYUwT
/QX83pt/yz/ALyuCw/BuwRinvURKLYiWBbSI1tWaQcKlK/tWx0wGy2fsCby/WxD0
8ei3jhLJbyn4VUh3U1oHFsXJ9SME1FPdqbMwwY8V1zDd5xHBhGrF7DyoRnrw2Ptb
t/ynNrblR3RB95vCWW+ImEOmMLdfsU8d1fVKw6Y2/+v3E/kEeIQTXYGdJbEPlqDw
9BVd+QUR778bZCeWN8EHL7hDcMjWgKpBMF8PYObg5vsU1GSkjdxmyXLJyeMQjqw3
s0O4+MrQDxKu2iWzSuPpSrKkAwxGb3MWg9fwkQ0CmUn1AnvRgWLZ9+AHvYWv2iwD
ihWworJm1Jx1qWI++Uq36aAusqo7EGXjlaz3Fkp2GOwcSPGcmkWTrKyaK+OjS4h3
iZ1TWuKzGxRTpRyYSI2UrAXzr+BYu2kpQz84WyE80Y65a2OwE4yeo/J8w2CpJyGk
uLfqF7Mf8pW93crO89l3Ys9h3h5sNuroBlaM+/TzE13uAC3p0LByzvZLs5Uuad7R
1zIsmWsWheUz4dnFj2gEnN/8yQFQDaGyECr06W213I8Omb8W7G4R//xPkn2pKKrw
N9DmitveZ8jlnIHNXkNJtm6935sP1W5ej017EI60rdLUqI9PWStIkYdMnvqwlS3u
2BHSGoO4xWsfSM+CGzEf9YB2kUS8QyXhM7Q+cxcE4V1JRivUcu0dM4I65tWN7oRm
E9n+QLjDzn5UFu3IytqAZwhZsZINBasTYJIkNKMTg/HYF1O+b0UMSCV6S4SxrWvN
DxJvmZjGohzBdzSphaN9oMvHgQt2VWrwanIZvnWTicacl5hDRWOiov90XPKQFIc3
U8Ahdl5q4rNzwkfCCfO63SXIdx7mkQKGJ5t0qL6jkwo7amoMeE9hXZyw2gVanqiV
/FG25P+zpxWGFFPDpb7Lyq4pIf9i+4zndki53iDrQpkC9BKd1uFki6UrjytpB3Vr
AWcgDqBUOfBRSWugsoB68o6Y/acybhVGhBV7m55BW4D6i7UIyNjj2hialLqST7Rm
PMol7+Q8SjpyIi0PDWdo1W2khroUzI/KsizmEOC6v2bxGJvLSAL0k7+h3bAikTmn
QSIavhecurMpreZE/9z0PfqAE7LUbAfRl/OjdFDS7YxDz+u0RMlBptde2cZVCQrV
ooZfI8zJXwJ6K5Z5hNG10gcXHUi94e3nPfYvEDmC4HWq6N9KTbVJmt8HU0zoEvZ2
TTfuNwEK96CVjUbR6PMsm5oqJjYJmZtAzZvUvIWo7XBzX6gFp796D9YYYpnSeW5b
evefDRPdNNuKG76mwqLA0F6kdwUL1sziwUbHIY5Fck+LF3MwvAUfLeWgm7SwWGJP
8Co6bQCdQlmniZMO51wb4OXNkbYDnCOforX5R5sBHCO6+kkibn8ymOqoLO3I13K1
wa0K9G8nyWp9CQFVk4brGOnb1RI/EfxP6TglzETXtdBYzZns08/LM5lCnnNMZgYK
PUgHJccT15FKlVz/9ELZdP4HEYU5HFWVYHCvF3msHa/RI6MoJPfPDNAymeedpt43
cslsYTrvEI7BpIgB5dhXDXRBl5LOPcPq/r8sYWjf70h9O6uKByTVnw4a9iKNPEVS
HoSN4G5vQg0cKBfoJxq2zDMgRDqN5lpQfYFAXfY1w32i0+0nIMXrA3rDD0dGDqsO
oHXa19x9apUEvf4KEhidCnUlnCQcCMZ3BWOvV+1qpjdws0JVC85hJqdSB74lIO57
TTT0Bs+prtd3hOFT+SUX+ujH2DK9i4i07YiBT2WmCiLeNAeKSDhaRfcrmYkvhmhm
QJN/0BAwSU7Kqq95ZgrN02LEEJJ2tQaAY/bcU3UTYHqJj/dY1HV0hSwMExM7lK+8
QC3PrBuuYWqNddeNCMYe0niiICe3F/VIDKovBboL6qkvfdSZG3kwyLC7Y/hRRqJ+
j+4j9abCEMS/W6iq2fJumGO9p5XEeDdKPYhb/WCGzNmAxphzidG8qyvVvaKI4ixE
AGW5ToZ6mCRPOc4m830QRE+x4w4ifNDo2Sqvb54NracK6dXeCdb0PoGYu1WZ6mKH
e7/m/eT1pD1JW2/c59UGOG/R5aRa+DsUkuXEkijtX/5yODJBBHtCvpXQVdtQ6eVh
ryieju5DmaSwpyxiQIU1fmAm7vhNnco5QIQUW4IM/fBbMxcUMCYLseeaupzKqRnl
laQr1xh4n+JXO+uRcJzhsdXXeu25fJrg01HKOFqxxQdY+ZrlguWUFJrxUZOXj5qs
kyxV8VyRJdA2bUP+CepnIZ6dnC9n5niTxRfXZ/YDLoq+Z7TCK+DtxrlrGPfM+LVI
A/u3T8O0o7wRvJEjq5ysZgWiQZqmbxHAeT4+/tD1d8cwp084NH5z8DKAxO6JkqXz
AMloDLzUFUHejXwevpgmr1tZTe4wITtE8ZFwXgY105ynfc/oUiNlC85PhSGA7+g9
Vm62EWKtpj2Slf+XXLy+cCq/IaNn6QicACq+sI3U4sXmgtoEo1v6F5cBvia98i+x
LW79PV9tdQoxrTd6dtHMe+qYEF30Uso/bonb2dn4esELMDd60Dwh+kh83p03UZRQ
5XoPmI521CUbxXsMwdjVMwx5Q26GclCH3zcp6QufavnO3hC7xezT0s0U4BWMH/Uz
+OUXLbbEQ/ExWId+UraufbBb1R+oz28hCsBKtdLbZhLaXiVIMsqZLhN3s/Hi1e21
zXSKrGQdtQ8edJYZGPNxASJ2fgmiSkulT+ro+4EMzq63JDp5FLvjYT2eRX0/ejfO
sWIkUQSkEZCxVor4qBk+V7/pKIpSBvTP4UHkCcX++/VTQpcEaomFyWIMvSEGNYsW
woZrYSHAbXzfr/VC3CmtkoOglNFBFSxoO7la9uazvMH06iuovrin7SVIghpj1wRd
hi+fWIsOqvg3+Cvjchzx1SARcN+y/SAraFPS2hbOMoSm4xYgUyO4S4xEK2COgiPt
s2LspS1ZllD1Npwa//LYJrozCgerZS877VywRox7khsOtpU30VCcMjLgVKzlQ5PG
YNw6Jw4vN1uQooImFqdgqZVLsai/XpqY/JVcnA9gF7avu7XDIeR/NN/3FG4i2Qjs
5/eNGglG1xW5vP3NLvZaHBneW2vyH4u/Yshcb1XynreHFYgcYZM6MD/N1r0MI1sv
/kRu2Gspg2oD5Z3iHKQRcO1lajnfmjCgvJQpgWnajAJuyje3gmG77yQecuDY/wcW
oZXHKsAe49ayq3z1YvH+pvxoTykdfkF9z5wb2U6DzRz2t2pr2QNlqLrmWGGHArSH
amGrQQiaaWV1NqJHVw1G1dc8IsVrvvSKjvI1qo0/Qj2PgIJOuwbi8jTUh5xoGl/o
kKEhxxn6QXYOb22wQwCh1QQoOcrxw1WQzQ4A1Jkqj7gobNRzg18JZLZ9fi3Hmfpt
5UIJ+OgFObc008sRujEvKrTB8tc5D3Y1GZhl/ACg1meP76zm/3NVDtbkwk3mVPdh
PIv2Dx//JgXABK2UtrdA/BSm5SxGkUXpSmWDdzI6pCxEuEpv/QmdIA5S+RA3rejd
mtzWVzlAHl3w5Wuz7HTdDNlBFWK6nU5LIcdzOc3oNHfDi7qVQ1nck+YJxWzpO9mY
JZ7BD/RND+cjlKDQBOPWuKLO1hS+JkxWRSN8lsxYjkjfBOdANjg5H2f0fvxDRm/l
yMqJVHMx8fIccfaPlUA6b7FqzHWl6nblyoT6uvnclIWMmty/7FBdTqxiiUaNAAGO
Q0EGFLBcUsxzH73zckHFDCUKGsTi51vwHvlESGBk01viD9dmzt53P4owZfd+I7lm
xb4ItBAsZ9tbUB2D+MNvsJ+dttSIDqYvg5QU3Un/ThOnDK9kLiZKhrLi5BjwW9n1
BCxtLeKYc0kOFcsD71McWImFzHhEQP9dTTZ6Yy++OcMf4eFpJ3RUJNXK8zhqmAN8
tYWwL2VslbJqrFrk2VmsXK9aghhuGsflo+2kfkNnOrbT86YV5OXDqx5xfs234NH1
zuJOs682VdtqIKrQ2C/ED5oZaUF1+B40fb1rA28DzSeRFma/sKTxudKIbJLq2LP2
3W41Fq4653Pi6HzM6MDEoozohK8HClf2yMoLOJ1tX1OTVva/I1p7uH6A+ZUFh9X2
HFhn0+Ijl5NNr6CVTbVxrn8qPdR5SjrhpDfUqJ/f0v7FixPVjo2hz0OZiXl0yK/u
9hnCnBQq/JmMTZe3ODF0znMIMnl8uX0kpyXIqu+8yr1heI3L+80met6qeEwkdGJv
ZBlRK8x7jpXpxL6l+7xrGzGAKdd5kyYiCBdeharPAfiG2ndd2KSWak3j+r/YiyhW
swHKus0qNhHeqEf3u6HqeQPnWw31GI9ZCgVNdTiPy0eGx1vv9DAykOp9L3y9RXBi
glDPcigN+PW/qFTuCFSeyyE/tQargNe4Vppi3rcIThOrCZjEHXqeCX9ddeRG4pxO
fTRPRdBtQXItL5449qm6dFDwk0D+ga+o9ugsby+nj9PkcYro8iWSQJCCgwGeo4NZ
saFCFJCpj7TjSmoouMZtwbI549RXZmWF7aWUyrY2sd2phej9S7sDC+TsR2KpbNeK
efqaXJhQ6JcXDIw1ftE8rpGBDIg2ZQWhwuKuCilXcGWX3udD59HLI4vAfVh89G95
9CyK27xAxZQtHvhJIEY9hU/OnuoMhhM2w10F9uB58F08SMfq87xqMwHZFx8G72UZ
nN7IYf7qW3m2ixZk3DBvKWxOAd8y4WzmutBgLjug5/i6CL7bDG/ghARHAmn9+0xV
vsCXmbS3H2qh06QMGSfW8SerF/Pp0S9MT4gNE/FQBRA8NxpKGIOFAzBzFu4iOAgj
WcTdZC7Vc95Y3u+/R4IxQpsnBEIcBhNEKA1jYKj0MDk1ZL4tk+L8kJR+CfIWXPZD
gGLVaET+ohUm3FERn6AnHWDFk5j5FmtiiXREqTrZz7mV5kjE4TNikPz2/rU5z9JQ
c0zUQYL4CXxwVfV+PYTiTNy0ht6weGFcm6oV2rzBmVNIDyn6N1mkztMA7SfF2+vX
sXRuDrle3exGYdQ5ZpeZXoBBSwlbyZJL1k6gzY7QyXKSLLO6pJDiRndjXzFqeX70
vNoHyVy8NtskvWTMMX2tmihoUyDVbeh0HRdTtWZbntXCPFMtFXY1rFjIl/Y7C1TG
iH89Zlz5PowaYOIUopBr6yWub/XwR1DZ7jSt8ElOmP3QaEkfpci1FBxGsbO9XBXj
84ISHzkqF9snHUbJxD8u0Sp1lor6FptZeqGwzk76Xp+ixf5QB7AWXW3lTx5Xa7S0
KcZOFt71u65QiseP6jYGeNHg8aGh4mtH3ncUf1p4Rf5jpkaAwzG0EbIeqSvFCs2E
gVWVFEfBpY4jt3fzG/Knck3qGSso9b61GKyT37pS1c/tsQttGNPMZxj32unF1xIu
69k28OeXQD/rsa3xRtQBf3NeXr3NjODwDiG/GwnZulsqxJiUtBRB7BlCpx4jKRxf
x9aCv9gmGfEgbRZogv4zcE1rj+LKQRmFvRxDoV/4SQ2gj/sv6ATjFYNucYYpdMfR
Q33lNJOlI3I8uskSNo5k+wX9D2P3mHav+4e0z70qQGVH9yYvie38Eh9hzgf/EvVB
hkBkn6fb6ICP0K13RENHHY00924QmFH3d1NcHm//GKAU/QPwsGqURgFnDMK96Lye
JLef3xMqTgQ5AHWOgu3fGWh4qbMLdx4qb5a/wHk4tNfTPS0yrxpH29PXw2vV1Zom
boQdeKmF99DfWYo/Eo6Ku8jYMTebh5fEVQbkr5V2EiX5fDL29+W/G6LMabMNfpjI
xBI32AzVNImf4Wk6ksYXBKyyz28RQDckWMGRrq2Z7abAczoz9d1gHqWZiBa6jTfU
373mD4bVu+evrwF8kOxyNVahIgOI0VKNsVZLbUm8kZRHeBOlQna3tn04K+6khr+E
eMMkyn4NdeYCNrcGQ3rQLWMcnBXlOAt7LJVwHJ7Tholx2xhBIG7hpToXGLGQgpjC
LTIilbopDS+jlS6e4t2dhlm5WeS49KPBQK8DOhDUk2obO+TsbZINnh2hGt3hTYAN
sFwdDtaC+WuGCbf/SWfZhtwxQtoaXwqtyMb0F5gkIiIgvCjFSOycnIWv/YwFKFAc
8a05Ko25Xv//8FN6QUHhop8rNCRMtttQfWvavbM15mTopfCMcPBd4lCRcOdHMfIw
syByK95rxZUk5QPbDXiQFlQAi/HwQYP8aCdyE/PofOXG0GZGbh6rMQSjqCy3deC4
hCE7Fqwb9tbI4fZfFBw90+zFWhKYwC7vLJdRCLNAf52SebD/6yhKXTx1uzP1pVWN
qF0ziDOaYywTYHMVOXznR32afgbuEUUn8Uy45MSIEdTWZlAvFH/M19fW5XZ16bsN
n+cUq3H9FHbH38d6ZCQmmV2QKBE6hx2uLMD3DBmdDX6ReecjGP9OiPQydpl1oPx5
pMzpLYvduvBfPHX+9PZqgZDvmKGGpfS0AU/nD5VV7yRF1JtqZVIzNWdgGzHMmSuE
LQUpVTgRsJItlqA+RrwUxkpvi1PIeeM7xVXLYIuq0WZUjaM5zJBPK0oTO0E1fCcg
mnaKtJrVANJavw2tQbnwtvLOwcqEejhhyA9NFTtlxy6DFLdmvvs6AyXnJWF3OqVo
PBmhHlGV8ecE07k/qZDsi3nExxiVkQRFYFRf7gedhJdBiqQicvMOxfEuGwgzhTzZ
vpbr4wCFlUf4ItZnxCyvdVywlf0VTE1iE1p4q+NsfZeMlPwUBMQfXO5U7duMFJvt
Tbr3ZYnxdXSK/CoOdSWkyrcB9fg7YIIhnQ4hRU24/xy6YhQaHq/cfX9bwQB2RRsu
qqnOpONAtS4FXo/ZHDDe541nN69vJHmdcV6ab3FK2ITBiakki5CkQ0IGzAS8X3dF
H48BsZCoYS229eWtCR0o7nDOKY2H5awyisvtaeVCliZMhd96TJHUVDJMqt5oFAVT
93ZJULwVGu3BOEEhcF26kYNmpZcWBABRUx12mQS7rHbWvROgZJRvDVzWU66FIfQz
By89ExDxY9sGBCk6JV5k3gAVZ4T+MDk4wIcb1n/BFMUERSfsBpw8hSrb97/8K09b
aVPJMoEh4jHfjDsXjUoBRF91yCQoUAPoa+3KtgUZdyDvJ5ANLzGCPAxnLHFYf4ci
MeO3ABKRaQFX59jxKg6G/ZVdKdL7XgfS3cdZnDd2DYBkQA/jhQY6GLr5HUApdBpN
E9Srfimr/wpCjXmSJo3QMdDRMwfQMyDrJOKo2gLzTA7Sv9gXRIC5ppS8mRpWsFQ3
tqNTXafnC4RHFb25642LmUSCTsNnV0CDfADexKAQ7fbHPL544dohzYITtvMABKZF
Q55nUAV/brwJEtLoSEWL5ILZcS2Bg0eejb69W3w8a8nYTdTw1SRDQldQGh/wQWmz
Q+hntNFEtCa8OowWf6PiJ5XJFLnpJwPz3ni5ujTggP48451es0mw5HA0H8orM8hr
UK/gI4kIicOseB85iR8+nLlLFvLOKpoppl2Ad8knwTSzIhbcChuI4Dg+5qnRllfK
kPXjIiwPMSHyE87jfpsG6JVQapaNuH+ulpFrPB/N6Hx6HDjGxSij7IPRs5BXEsFj
49tZU1vDwUUsQeetTwMLPU7t1jWELeZryKJ/qBklmAAVkh/WBiK/rBws4z5umgfB
wyUJLd78w73cJV4o8lsk6hdqC/k+ZRsq+5MDNfe9XiU6IoMBnIOxOqTcBf0AMVgk
lT8AbXqj9E8prEFA0vWtPsO39VKzeK7w1Kv4QbDdpysFqwm9PUDLy1fcDKr+EzDS
EYe4rtrhPwVBGvCbOmwWX6aIN90lFM3aPnS84SBiyFWMaAiuPiQx6eI5BZYyEJeC
afjlVINq7wv8qo8zrPt3e5U6pM07C3vOZJdhz+lfmeS3vWWnxYKfiM22RbnzNLI8
t9bcgPFXZCFLdUzfSvZVSwchp1G/Ejf62K0ktzYPYFZHY62ZRuYhpPtUP4EpeWYk
Gv22e/g5M3odD+Ltd7uiqd0wemZJSDg8K+BkOIcQgnGYebHvc8DweSnthM/oguUD
pY9rCbSp0zUexVA1EJkOEmPuBHLV93zt3Pl4VTcPtlhErYVfOBa/KtW8TYqllB9D
kBnN3hmpSgYtE2DnEjhxJ+FGq8HSAbW8hqSLdIHPkGGTl4JwJG2NP/kRNufmtqWn
5sRwGyRFuMbtyjB5RMTvM0JkyXa5htRPRng8udpDokj3qvCdR2rX1M8aeLRALgDO
P5bBaXIyFUnH/gxTg6hmAcaF3URgU8U/tDZ5++wxT8bLlurJjORtL3sl22pKV0QH
A2cShvycrX+/rqOKJxhDlynZT94FxQC3WBly+LCdk2Da+dFFSWzIjC2Xf9Lg7NUI
VLMEUfXp2+wniKqivuqxklsDAPf21ABcJcUEUF5B9rhTNyKKbW6AjN9245paUoyE
aMoakSrw0G/rCCrSsCeXhynedI4o6lLL7cc0cDJL3vsox+xlakPhkOci6vKcm50q
14b7E9113IujKA5bf9l3ePC/Ig0EL0JV0RmLU540gcOtj337xO7X6khnlxbVkIMp
aJzknNq7ppLQK0PEpsWVVAO1KFw9ynflB1JR21qompPbEg6S4/dno0VqDqpnR5iI
LVUieMgHrtr3XbdpBm9aCABfX4p6GrqOvjaDwOwXVrjsaIwlEKfAtyYtJzUhM1Nu
hTIvqxjgS23xUMfmP9QXpwZ5a53+BsJrnLWDJ0FVEtJnZycYLC2wZb1udukx6s7s
NOaatgEAv4sw2knPooVZvXjS4fVmROhXTIGdSCKaeffDz4C2I+ea4vIYjxtXguJI
FZSts9dEMMtWeookhj4OmqZkCoNtb4hAqG9SRZOwTXXm16Uf4gK0Lp7s+vGeL7c9
LGKhbZwtp7OaDKTmPoOlNmKFTj3GzrSX9NfLMuRfRMxzOV6m3APzW3pLn4bZUodG
1Cti4VJHSUR2qV0Xq+7jBIuSruq7thVfAwAK/aZ3znBYPODp9B8VsIqM55H5ysFK
Q7GZmQBuMQjk8cUMYm8qnlL+VPNcgQbZnPiaGlhmmkw9Dj+FXj4Q3ioiL+KoUWGg
oO5SkVzbvd/C5ccbSQfavsKJVV77qyyd9XenfCCOWpagYJhPcVyClBAJrOw+5ZEj
4P4qf63l3l7V5jUM3EcmiPPTyrG1bho/SwVkMeIonZGUeErntjYq/4DJgbwFjgn6
eKQvq5IX3/sPf6SX5jogpZEdqab1aO2Jt52DvUG7HzTzFPwY6QbJK/sAbS/shLGh
0qL6YR2BOZ2+Ab1Y1DS6qhR43vNCbDT3L1Z1t4EtbNPVS3dvm5atM4ziVoUvKO+X
1y5krOBkLBlNE0imHkUew1nSIGQfme31dXrDMs9HmasZwZwYnlTFxs2TZtvon8DZ
+fFACJ2hjO+vAH29VdHyCIrVGXUWS6U+bRtW3sGbaVQudEgUFVBhrG9qU+p7xSTQ
3V0BxcU3ngixRZI3V3Fs04LIMvXLVHU9Cw8E3kBgtDo8M8NYxAn7CHzUZ4LOVPDe
YnujZmzurEvbl+PsPrL8i3J/IO1Z+d5lL7myagx2y7qM1JJbaQWWZ5RHEmI+0xyy
8C+SmPozjnyDa90boFh0LmHWRq16QYe/mA8EIW22q+wVDWv4wmMdhH0hhLqrZvsC
nDCB1hukDSHi4s1Phpb7NHDP3EZuAAbdEnJ8uUXmJSea4q4aRo1S7gchsM+6TsV7
6hsnpupfZDOrCzqRRHG543D7lZNJvaYeMAYhRMZYDc8wrggAU2AGWZ2AYgOWxxfA
/fm080xG2ySCLH8BYoUTl0U27vokWsogxfFv43UzsgpAkgID1TuOySgNon3ZM4Iu
UFjHuJs871sezgsYKLgmvOW8NuANDjVDiZyojiz58EYCyyqfCjSlo8l++D582qCy
akCZZ6aHnd/y+DoONHir103HL0p8GbGzAv/wdC1UEJgbzp1nnzGFNCCRRo2tk3wm
cteQp2ftlKjUVBTvUA3Hsos7ICiBkItAO2d4reodgtUBodHbapoP9AfMQTpa4GIo
nJFaOsEak1MWsuAG4gM/l6uxbFpqSLAs7zXUm9RsqPUgeNMjndDcxa7I2vPlEYhb
HCAu05orMe2QNw6C3+ayn/epoa8uW+imJ/Lna+5ji1gRXn5dulChx4v0ZswtN077
Xj1L5stJjTzlISbDbXEJ4FNZjuOfcKrbk8js6/yvzRN1m9nA9B/V3tRXApidgsZf
LZ7IqMpoQlQW5TTkuWtBN4qlyx4waRdo9QWDe86MIR1c/smgR2+zMQiaqG/Z1qFz
3b68CXvd1Nb4NRifjYLnXWmZ/RpIA/ZUl1c/Q/3l2LsKN+xJcC55o9MnBKrsuolk
5JP6Nv7IqkDly8bT0n2mOBZFVG70tfIukf9UNnLB3mCHgrDzNQIeSnob5GOJyQ9g
vLUUHI4cvABIhf4eZcIgWg==
`pragma protect end_protected
