// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:05:43 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
UdhzChg4+qj6+5sX2uxQoi84sFSwbNV48CoXQrAzIoMNilloy9MlncgSprNaf5qg
a5zDN2NDuvV9b6jcmqkwoqrP7H6yXJBkmktojz9zs+BqlFanWvXodT0DJ4XuOzwm
BgIpx++DMlLfJK/NuIjNzoOgNIowe5rR7LEc9ycnGaE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 30144)
RUIAOfPxZhvE6qZ6WqvILU6svipSANc6YhNC2C+FS+rxt7G1WL4jOz7DJsCyZIYF
0AQ5H/LDuevERYBH2uFKBwewXsq+bNUeGUCL+Iw1iS7krsy4LJ8sfiFnqroaeCM1
j8LTWqwNZCi3uNlP45EESu4sJWPCNT7aPjMmCniq/iM+ZazENABKiRjOh46PZ/7h
hndiFOnwngdFQv12vkSKYSEKgKHU8U3w4z2TZ4X0NNdNGmOSnSOnbzFRXyf4RcVt
MLlTWKeSYwpkqqJc19Xp/oIiNqahYi0yklcPpsEG7y03OCsCkJj7g7fBtY1CY1NU
JjPdfSUU8NOaySEWi950IaRmUo/91bbu8eN9weSKtcOL4L5TyCUSIYYjsAUNTUY1
G8Ky3CWHlLZ6eS7VRQItk2tbMclajmQBEhgzTOt43gSjeYYsu4lYom9zLVn3WIgr
txc9ip+WkbjymhCdxnS6IOG+UKcX82DclwYlan2CjLPw2cj0QtEbdC2XuP4NRmz/
+71c7z0/9NSrHBzur9CNaoLYxw/43y9aQctTEOFcSMPl7qDdrOPnFQIdxLKcVQay
lhG3xWAVBq+f2T6C1bWRKYfeh3vscRGF71SEIwlAFoFVwV26NV7K/QBtmXYtGJqB
npYRRcv0BACaDPkJM43BIvT+x7BSGLmiGD53SBcaa5PPNy3lv0OGD97fmksPHEJK
mjySRDOqKjFirUdmJutTa44W0cSZDfazsCMGTrSuDXhmNjhjZk+oVypTwsQxqDlt
WMUkj5h9rAmOyuomiaM9fHnoAlTK/fijXUkDymrcDSdZEIxuw9Qo3iDu5cco58RM
D+SY7ZgrdSlGhbcoUWK2jGd6N2ks/c2bWOLBGKHZtKNBfhEDnuc4pcLRSAQEqX2b
x7ZxzCbAQm2Kh2b4VZN2UhKJVoopbduH/R3kbIDAdZZCQrwwKajGztvvmfa9VnNT
0ut7Ewlwdg9h7j3xYWLI3pw8PGAkSzcz1HO/2uCgO+apoIL2J4jYJcXF0jaoheDK
w4ON/gxrqs/ernaZALGbgdzMjCyJobUPLaph0bBTQMAyhI+3JokMSW5HAsmwuUGP
NG0TxqI7zmnKzYJofSM2Mf2uHrAfQXsS6xiErntLUJTgzbyFTAifBGAvGpuUniDm
rbvVsb3V9IYOLv4CMAmXJkhsAy0TgQkPrA6ug1jvRxsL653l1kt4qBOJREmfbKR2
zGBMbE0FFtliLMv3slZc6Adc89cQ9oiaXNHI8y3MKGnfS6dUdGZrlthlXCP2qLMF
tdPzWDBaCiGD3SyXFULvFMmBYNrDhbcD0XmPtS0jykkMuUKes6tBHtQQJVJXks5V
amT1X8/FZD2EZyWnhzo715xRNwfURH8vcjL/fs3Sr1RDtinJwsK5VZ9ARQTExx+W
PDjGmuVhR6k9bSBtDJDIqjjjW72nQz6ptBu39NLCFgwRZkGhjQb8pvKyaXLRxl2d
tWSAJ/hiNo+s9lnmhs+RcCwQNKVRIZzxBXLaPFPSkLeTJ/8No4uXd11a77rMddcT
sAmxeAflyEFpQ9n3QuvRavkDzyPFXf3eJWjTIGLk9vlmq6JxMIfpdE3oMvkN/hr4
NQRf+uDaF6982VNQLs9ngIhPGhJuHga4lUwRSwJpVixWkZXFVtCfMdRyIYOdeA/w
L0pg6NwXTXsVtsBDytUIQMu9i4MXwQVHoLndJ98QlLk8leKG6edz/4MjwMlot4Yo
49YiqRaAYEgCxTEyaXG/h8erGdVDMyaXyqo4fWr5QFPaJDFKOmZtZ/R2mm5X8RFV
tLEtR+DqfGIOwbwonulrD9YyRlTjslcIhJzuIdw0jd6LBuEWVK5xITXhqFwd75cB
jS28/f6m5WrXqA5SuT1azganCPwCdtUavTiK7hQ8GaSmLo0j25TKdrPXCe0xQMbs
4K/eWPkg4aAeHjuH2ndDUfF8tZtEkXyWNWFt6piSTjR1KZ43mZOH30ImR76gzybm
tvtmBRWAqe817m5p88j2r5ybWVdB0z/275QcrefBZo/sZIpKSd8trBWobe5JujwC
XHTFqO/o3rqEgUNSR9m0B8bU5RWXa5irmIUruJl0HHqJOv4cQ5TaxtYBZJTuewvt
5dSwoVBOuS4coxNiiRgN/9MhwMYPu9s2IhkjRmJy3AJrNT8WY3LBreHUm5VAzWCj
+9P3x61+n2pGoio5+rFdAcsVToc+2n4g8SWT0KGMpslvk/kpU2qhKl/t0eLBQE6S
Pma4a6H9LUQkIcbInLWupdmcKAPi3VpYxrpH4e+1bAmXaT9sY2Kb0raOzU622Lm7
n7La2pWk7p/2Ha6MpL9yEiFYSoEY+F4PsMztcr49P2oLBpfT1T3GVCCPHZ3bhzDE
gnb8yXCHwB9PZM/c2ZWGZtHgYKwRnWVg2JKSpXRMbzZCL9CvCql6lpVrgoXEAwej
uRlBslnkjo/+ff8sH6yhKNnjaHXU/glFBLKWwARpsnQ/h7ECv3Tpxgq91qBrfrxU
GgPWC3Zh1usBl0+Jp8VeHFAcjT+FYSx6Rk0uN1hkzow9GDA4+DerdSOFYvmlkdDm
tp6DzSqZm95CTirpw9KyJ/+IgYATkwhz066Uh+r5Om5W80JPerkouAgKa6eOdQ8n
cs6iyrtrd9GFI2UE8q5iSuwlAAAxM/GygfA82zhV1IKSZIiWMpUHsRcENk5kXo2O
3nPDrL0pPpOQFN8dJZ4bcTEVyU61KGermrIEN/HXR1hSF8NWIc7vgr2X3T3uFBSI
ARqpwRhstfamkGJU/xXArdkML7QRsmz5DjUVXCn8rn0S/aEH7il4DSl5nr8cqyIK
1m6qcrBSGuh8/AB3HiilLoRvMPYFK36Z5cbZtzxu2ioSmBhJzIDG1Ql0+1L0wKfS
oR0ifs86l82J+j921XRXCddF265+ATBoByiH6Q2NNJkOyookxhVb6N99T35wuLuD
jIR3hfbPOy8G0OS3dTzfjibrtpuLSHyRdz3W7vA5PEAlNfrxEfQijeRCSrCh2n/r
d0eYV4sAhe5EUs/+zm+OAZd62caeYF1RGjwSD7tbKIyqnLk6jQo+KxZ1GMyFcR18
sjDg/U4nEjo4eqWwzVMoD4ql4VF7OSd0yv8FC3aPkFJAdh7hjpYkU2vvExM8hvo1
Qh8NdL7KQQjdkpIrvL9MeM63I+8DVKtKf4EflIVJvA7xJ1deG4SqTEXFFCi6ssHW
83SyGzjo/sJuehxY8XD3A3ogViqqWhS2ynChjLQll8JRoA2mB25pRB7UIILde+O4
UdTkhogMiE+ekkE62hmIqbH+l7i8VrOFoa3cAPxEIl1svH6/u9Yr18yOw34J4mXl
IuAdTpiKFfFp4Jc7wyqgu40yYb8zid4zc56z9h5vn+6nm0D0yOA+wd1orxPygbu9
zd0Jrq59YhAbslnhDqstGFSTPJv8ZSxAhhK4cpoFn0eDcT7SrMQcC0Kz+T1Uhk6g
JtZ/423yCfGEw1cDll/UOAzABm/fhSr7porRCJd0LBWm2eLaaFed7LjonoX1wYLR
3isPxP8eRW1saRLPLAoaArMgbvk4rgiEMNvB7ir8CU84OYZb6tMZ58d0nFhj07V5
oIMgZjWdDnPdDEH99qOhcoAxOtncROv6oqKc2Fs/lgV5vkKhSwLBzgw+MN+ncZxV
seKCxwvJwrmBXwi0SvVRbVaLbHa6HD691374Gz4ozbw4Le7x3d7oK1MJLPlv4T4X
mFd3vdczSnIcSClgOqhjomf8VTkrY4d0HLd/cCeI+hRKIY1j5lQsZyR5Wpz23e/M
XCbkJveQY/QcBU68UTGSkVy9uyA4JymJgVGU4P1EuJHygVfvOIv+AT9UZlY70nt7
1ymiAJIVfnow1l8M4SIRiy67eXdKf7zHwiKiskDFVBTOh0RDN+8OPVfGwB1lfTrr
Y3XBQ9D7LZbLXutqu3fBfennwRKerRVp4OInCMze7bRmdvEdQ3cYypY5xLmu/tXT
l0p2IIez3sZ+x+1jbU0oy/mE30KW5qL+/Su3y66KUHVCn8CfxSgcS1R0VRiC88F5
72ksf1FRvih0+4RJ2bsKhCnEu3Y0RLRbPLct7R3XhY/mPKn36XStCLLUTLQ1p8lI
RzP5+mt2z58KE5z3pRPWGjVFpxNxrDLhiSzQxsAkCNdHPqb4GNXreB1CMN1Yh/RT
idJ9oxwBPCWy5Tcd5bg/lHAq9R3TOBoBGcwJPHZaWxm5esvwm1f6HzIAgzRCt0jw
py1SLZ/DUSoZr7SNlFkE8yQokq8NEHopurPCOggN003iV7IvMQh9vHBhgB1YqGTb
C1m8qfeMkoMewn8Nty1b4Ssi8izBh70YzkgVd8OUjjRu6w+VKUJaaJvhd7Bu4VWc
pT8JsZ/CqztKiak+ixZjRefU5rZ77wkU20mT6bnQuar3VDjzS5QjkWlWgYrqd2d5
6KwU/1s3yhKdWkrCyn8oWbQbGnmOQF6wdhvqYfEt2sknqj66/bLfs8fTQqwOj8IS
occxMAnP0gnRHRrTVDLh8yCPBtL3k6DCbfT5qI2eD8v96gZpK1Jl8GklzG0m+nUl
1G7kOC0MjCUw7vSnIdrr6JqR+Cvp6Uf2dDBROWd8nHAouV2RbqPLaqedsJ8Bo+Y4
4S6geQmUgKsKi9d+SH9W9RVZI6S89NEifQo5TnsDQ+jVyN0qLfe3f8/Y2CLl39Hj
3lvoCN7YNn+PVyu/eDWbACcthc8IdS/7L2TSFEQw+w7EudWP0jYU/lLsNb/U48i3
bh5S3yzjmdpVjfREWMzCQ3dt5Jy1xvNZA4aUjcrBvMQGrDKonQ1BPhPvqFbx8l4U
rfjNW7bcG8nA0F+cU9AoOTKv46kE6Uzy4o1L3WKpiYKp76pkpgETjKfemeCBhTbO
6+MgoFt6IGJ7UUwZekgJbTrhMRnwdkZCVroqDs2nI38zji8+Fv+wBKgpKs9+qi/U
jG6NDdx1sj9l4sbR3iXq2sp8EHRti21qDajhWhAeI2314Qj68pD5n7TppNf2sH49
hZX5SnzmLMAm5Ak4ExTbbDxIlu72nsuJ/wKvnmtMApulNPX4UzYOkQoAyt2K8RTa
zWXHrizMb5YQEHuwZ2lirzeWgyKp5w83FKmC/il0HvJpPXotjfzPuDlhmrbe2OKc
wo9tKjOnI4GA8uYwUbSWDsQaBWQ3yBjoFevAZ7zySlt5g0qty82RQsha3YsZ9a6P
ls9I7jWAzLXqHTtQhtZIA7iXs8wUZ9QTXneus4433Ae5HRMqAVGqo2rrW+etv9gK
7hAYDrlFP5y0CxwCkrDZQe0etYyVgUUxMw4s6Sq95HR45yxKZaeytfs0nIdjXxN6
Vwp/Z0V/JxNThc7wRPkK3KImA6bDRd5kjxHOUNVA0bIXaHLHgChztsCHmJigZ8gC
xDbuLmJi++6RvkiqAc95vJF0KPHCf6+jslpSYGIFNxdX8TWp0N1PbmrTwzfq5YoC
N72D6b2TvU5JvDDcD140iEgPzcO3OWx7V/FuQc2vKY+tCHaswDtfONzjAu6rVIqR
ofYUFEGyllgBIuLSIrFGyttBOAaCX2GSf6E2AhKKprljxgSTifhFVaDa6EhN08ls
/qWQ2DQFjx/yMvDlHOBqixTbdiDQCK6O7oWNyYpGPfst4uT8DoC1zPDSYRTmbe9N
qjGrmXyHhz7E9x9hGLsTJ/hGFzbpYFAur1xjfxoiwnx9+v5SHaIz/l3MV5RpUyOM
tZfdqf/Gej82L+ib9+Gq+6yXj/3JQYX/2aPKYrPDNymsF4LyjWOKhddLlN1TxYG5
1Tp0n1d4PnQo5ILMFLVhUsQe0sugTuW6HCXhy60tUVaeBppdYBfz3BSFRVSA0+VW
zjIOkbaRiq4vZyjGOGHz62hVOt2zLR6+4jSI2f7imZRPvYwE9uQK3rJQ/GnBTCli
WuYN67m7xYQ0IVngsanxPRrFyAtNQ6/LLM4zEgxCOM62KNTGDRlTD0zLUgT5NwpP
Trv2OHtY9T1d3+azMOX3n4SgvXSbroge7uWvr1TJ18Ll9pDNSYW0CbWU3wO3dkUN
8DHuFOfQeVqhAtdUGyV6x6oW55EYUducpsp440RRoGQCfwQqO9sd17wo3svGeUod
fFvEG04zezGSiWZbsxrU+ofoBm1wYMfBhgbYJcf5JodZgcDb/FOmELhsjawPIOVK
WaV2ll1TpIPrt8PD/8Nxjg8nJnAhCzql9sVC4w+hFJLjtyfLD10N9QGxlOq8x6f/
1h1+s0+J4izkAVtvVXFs/jymcKMtIvh9S6/bhJYBWzwnMl10ZPqeZuDwfzceKuXX
NuLDr4Pe2kHm+XbrHGukNZNfrcExx1cC5lCsw5cT91wil6QuugXJxyUuqNCGiDTj
JhOH5i1AOT5iPiYxBKAxHQypIY0YWsNmHB2qACbBJJA7B2kb997C8nWNqa2mMmXt
Vv2Qka3a2gxF+qtWLmMKR4D4447SQ7vbg62aFviakChOyc2OHnMgl+wgC21wJ5ax
2Em5Xy+0hyIEigjhTZrWoBMq+mRUemn+Y40PsyI4sKPbHQpOO6tQoi5jeJDcK467
Zq37d393HCDITTLhLMUPZKJfivlDJEmhlq2c9R2wwXXCKgGT5tNMoYjrtFf/mPqX
SPokrd8DIIBZia+OT2inSHz5Xk1vDH8BMEPjOQjdaymikJu7Mol7Vm6rMyZmV2xI
2j7GR/5eFHYCVYxlbAuTJ7pdfCccqWBdf1p8dKVoBhNR1zysqVma5wwiUX1YYMwN
0WeKzDtzcGjDqTAWeIOh++qSR72NUErzVB4c3T1RW3y96ADZp+5pT6uDZ/RoGuK+
tFB0/oYembFykJmNnqcWUeVwh4pxY49JZU9BGeuA7S8PMbwdKt6Ri+wSsYlsrFKz
SaH5dbvWT6THQFvo75duCAgpeqv45RvtDmMwEFe1scgfot+CfSQS1PzfRSlvJg3x
a91Q906ssitPZrt3miB+vBbZ9CKpprPr0AdYVch3BdoPy1xYJvAO4/thHrgoF76n
jZ72so+uKzZyPKnmIgal6QmqLI53YmSC3Zr7tBG2bfw1a/u6mTI7GMUmMQ0ABukN
7l9J3m1zJW1QVBa8v2UIshrnYIp0WwtOxwyQHNd2qhXEngbAgZfUFYWhPFkteTu6
ucLc3r2TLBTBIkCYf6eWSlRFD1FKTbJVLC3Ek3CbK79EH2/+KLcH3slQ3SdgnFUS
tRgZ8Vz6j/iNk/Nq7d5nw51M+RNWX7Dy3Jt1cV3QQfExoasO424e9as9i3wY89uC
fu88804dcTFqgYckh7Vw0wzudtVJBdO/ZtxQxiD/fyWBlRSYTW0LuPT6GMWo01EM
VO5vww598H5JfQhFGBW/tPmlcl47IW395OftCxKenhZbOjMVnT9P4QM+WDMzLHIU
vmbS/rurUhRkpxb8+MSFxZeJO+jvUxkosoZE3J6+etCdCB5XPx7BVJ7ER9ml5VmQ
sD2Q0QuvYWhiQupkp9OIRQsiKxJxqGrgAP++zNmnNC1aGsgZ9cgTn+15ycXDpyBX
u1oXU+1cTr5oTOUPOnKo453GTdBUBrm0Zan3HuoARiFwwrc0zW/Fn+xGR1Ii55YW
IL16Uuh6c1ZEILB3/dc44ZG0/BPtGYFWDafDveYlEOzNQHNYB771x8+SU0ybpIjV
mXl/Vfc1omemVSsMd8Wfa/V/lOmG4SOADJ8xvWffEVJ61rmDW41lvv0uSr+8zUms
ZOnt3DFvbJreVADlhxEmvCNtTlFqZQlySh/eJQgNR137pz+6vt85tTwYB3B/RhOn
rORXX6VHWX/upz3uPcp+Ak7M+h09jAyo8afNYlpQ/Ns9aTmtSuoiJx1IckFEqCJp
yxLi48VBTh5NFFDjhW5g3fZ8FefZGTr7Q6OA3N/RdJU+/Zx7QQAsc0tFeMhcu3oI
LVXU7AzmSUEbfRgxnTmpPeEylypJhsxtg8vYcdyLrycqH717ZQyd5bk3L/U0crLr
iQY1Z0i2P63TwUdw1fbFBJPLXbVlEB2K6SDBdTQtRSYHV1xtHOXtHzdePE3Yh2hv
SocddAuIZt+whBM+DTdLcoA/TUFa6wYa9q0KK8n9y29DeurpSKRLAgmmsqzfxPjq
9WYZiqecKAfG9y3SLI0+gfWqaksa2Q9Rl55SXmr2LOvALpq/FNGihY3KF3ow07kg
QsPX5nhBB13sLifnpanUw9tYi0gGE8ePL7l2QkBNfW5bJ4aG7DEruIIRreGhBTsi
esYJ90tzUE54749swb49TCBTDKqQ8/T709m8k4BPlfIa2j5KFFDnDZU40XopDWHe
xhP0Tw079PxO1B+QyJdN+bsob+hjIylMm/WUIeD3fSmmN2AGYNpmg7KMlE7GmNcK
hdtZ6MdYqHdzGwcyajXHW+dId3CO7XR9gwDnDtayMunrz0Sodrm1KdPpr7RHkCzb
cSI8+tC2t+J+gUoaAHVsJUCOeyHoOcn5qWdtLnp8zEQaXzQyJJOPfDR59j/QRwPT
LA32LoheOdLBtzaeJ58C4DmzM4QNn2JVIB6yZbY3A8uAKtxrjCFtKvrI366N1Vp4
CNgc45XpjJ3q5+J8bowfIe9v6l3rQK/tdQal1cJPtlLxiOlBJr9XG4UO16HdJS8L
Rz6VKlSBvT+F0ufutg/p1xZfdzQ3U+TmbzQOX7dE8dU14fnnQxWGOTHPUS/+Evpy
C7xrRMvqfzlQfPHt2P8/G20/URxMDxqI7lywqRbW1UKISza4jrAbVWffjva7bYOj
5Xx9ADzGYqEjL9pi9v4w3yL0JrUehhDxrsZIPobj3UymTg3UB7fkgwwrGC+zhKAt
hsAx6Wveok+mjTTE0IX7IL7y6X3LNNMDHuKtlnf4OWAsducrV/s0gwlGoSFrg6Cr
mlTaJvR41i23x3kej0sNXQqqryKlhD5iZyME9PCZncDano0faAcjGyeHCiy+CwEA
kbV+Ofp8OaCxJnUytHadnnaJbMRdQ5rgG1KVa7Fn+QhR5ufOn6TbCFEJuDSd1LXc
6JVnDXIpK7+bD+RaobqrJWShfqP/seKQDOTevPiW1nWvfOpcZdBYm//SMlK8PQHM
oeDQfIKZ/FeoD5KxhDBdyy5rmxxP3AEU5wW0JqA5tFoQVHk9N6PClEZhnnXr4Hvg
CSLhkmQ4G3gD+sSsjpUEcQIqEezAeXWGTEiyMuw6DHSp/meD43xvyhcwkwEtV2uf
8J3sdHY2B1DIz23De/RD9gDSKHVYViLaHfgzage0XDYhY/xmlt5HpF/BuYA1F1D/
3hYEOkq0V5rW4Db2fSRbquSEU2xpkvOfFoLzaBhjZe72Auy89WHK/LqRQsyeqlyd
28yfKC5O717nCo0fGgEskKYtQ+///sIXkSTCsa2iUwszAP4ROw3XtUCgqheRKBaA
P6v0aEfuIwvhBJJWFTXFSaWnof/Oi/nrG3jyd8lr4rKJFoOfNcX9Gxulw0I6Sn6n
yLESXCHmXSWflQS9iVOprZQ5ML56YferoAXHZIkBSpoH7+B3FmmFL7ApDg5cirg9
yH4wkmn885ZEFSpcYYqxCMHHyZcdOvMJ57vrWRWFopcIQWsX3IVJlYTWTVkmEwrG
YvKwJxiO73+4iSswsjVhBDf70haey2ruUn0idxi5krgpMv0+q3Oo26DRgK0CiVGT
bnzYCNPrAUvjHc5uQysvkgeXbwax8cnrnarfxZu21JcnzHvxd9zTvXzusAiE67Ya
n5mSOBjitmY2kKxo8ABPKFLr8EvyI9Ld95b3Zy8EVuvHb+H725MoAjDnafCrIKSV
BJ/6evmLBsVXf6EJ+nHNHVIXJDSsgnxQd53QHBCjcFCmauYoRiydzq2cfiZgKb44
ONyw2G8K1n7PNMRhTVa8GqTUwKM+mcW6/Idpa0H+FMyg8P/DQiufqTmCLEdpYSto
USRR/oa7+jaHsw06TLD7cjc4JCbiJGUKoC8iD7wN3LC0An3OpZGzY7IUZ8qTUZss
NR/HTyB2qev8a/3bn45ATfpiqTqDBEvf05gtw5olR2zEpXtjOPXdVI4509r6bMba
gAgVibb0e/Mr4MTAi9pvtC+nuCQIib23bEbs25jQzZk2IRN94U9B4ol8A3rrWPw+
nqlrdtZKnUNYFPPr+onCEmrbHhCZ3A7KRDsXvdRUNilAHVnq5Kpblp39dOFDGiR6
hZkwox7iIYThvZSsXG9SHEi87u7eY3IxIe75Q5h0ewwoe2FIj5ajjRP10LkYXSLO
vIxSZl0cKbVEgMuEww3iV9E6ao7tCksrbFRZ7j4arwYCwedkTGlT6YEUifInYj18
TSA94R5uAeFcEui8sz0YWROJCGcKAxDwIJ2hacSVcgv6IFHZjxBj/KUGA/OF+rhf
grcDwKzLrZMn0Jf+9C6tvDe+p6S9YnI2YLsyBj2u3CdfwdKeuJiO+4fbRI1ZtYcs
8mBbkGJ+exBvZPQOI+rDYdf7hn+kxXR+NqTB378Nw3YLhCOpIvlKM79kCQ7BD0VE
bynE00Iv//vHMjB4Gzk/XydvWLKms5/5wQKNtEJBAoEu0mNUE7XXfi9forBzv6MG
HKlpWbkvPqpus2LxeAuCareRG0XYMpMJ0oghBtb1Gb0LrGZhJCgsKGlezQ4C8fYq
dtjvIyLgs1Fbo4GIBlwgMAz90vDfDinNx0azghnZfrMHg/WOkwXCXuwgKNr+tYU/
50jgnVfV7vd2o/CIGxsPbpyxXE+capDooo0fGoYhDFpDpNXtTyGuM8dLdQzwaRSK
kNG6xhXM0Jhbq/QFpF3X7jRq+Htkbk10D8zKyvsZxfEkkFWb+X9QLFQaLsvQQotN
faCnlUnggZQlwM+XiAl62YJQfwHFs4KuTiIZDTRVE/UBi4ZfLos37101PaEQzcr+
4Z4Hw1HdTToCO6Ylua7e2V7G4FQYzyAlEu9A/w8xOx1cwkLWR+uazu0jfIqp3IE2
9LJ59IvJqq286f/ky6GNdal+e11F+T2G8zxZSpQ4kClJ6REvvhUl0QyHMEr23gNU
MGJ7+45jukMwSdfl964ZXS/JOUtBhXj+ovbMsqyz4zjeofdDzLyXT+vCpaKwQfkG
PaZ9eD7gELIJYgEX2EsRB9dXLBNvZbGH8C8CAsOSXHWNdOmUKdna4odveleBe0CW
dD4SZ0vXrhy5iNAaqzRQ9+0eC8tXf+af/Iewc1eKEQ3wMTmTX635N1G8mMbnCNlD
4qLvuj9+YDyvvyCHjRpvMGoNXVm4sOv99B7kIebecsuxbT7waIBvZqfsbYXLgwbV
QHO0vve740EA6QFvWrsr1jLd+Mc/MXe20dFJraAJDtcjvLg7Nl8h/F7Q00eQEeth
qLO59oQakPEU58b4xKb5rJnBw3TvoynZvuG/XpjG/Upy/93SnIrdww5X1/X+InqA
f/sr2c0Q1jZLonSBd5A1svr0ECwxWzfYU3hsLasHbcYsEoT2+Hnt8HwnrKzSM3oS
pQJXL0fsu00po5buleL+IdUYCvPcmGELxQcCvcrZqwMnm+ANIRC2F4H1yqPL54e6
+9pORz/oCwEhEpYc5ckaUkr5Gnw6BXLZsCbuiQgwclxt820SMQHUvIv6wOoOCLj6
MOuoGu6RxhI7YmSLFX4hvx4ixHI8vlqWu/5+2Q6Qqk5i0Mw5HTTSAvGZ1lmKvrwL
6Zw24Hb7tTmQnI7fiYEY1rkZsCNYrNgV/8ojZCGcgGUaYZCLgi3t6gb9h4bd5EP2
AK6jFOAUhkOziRparmsSq6DR/9+l/ZlvByliNf3VQzJfO9ZxtxxZpgiFoXYJO0kj
xWgoipRmW4P2QL8MIZI/ZyCeK3T6t4/+s+7c9FyjJHN9QzAlHa6vdJd5+qDb4JrI
p6GqpRZxxUHhlEc4a87cg9GN0Gcu6d4Uj0/FK10gqhRcuwHd4HYBPHcrmb9EP3DC
pwWIBfUMLtQWZehOyzOcA4NBMDejs18q6q4dXO3Yjti7zC4/1DBnqERQv7SrqihQ
abvr6wQuo0O6BdFTQpaSJQOZJ6wJvk/bEOBLWwHZLYVCqT+z28YbyAxIhIJPh2MZ
P7k6WqlCuW8G6S665/jc+qdguPnsvCljv3PuOK0fi3BFht3+U4a2QgLatQ0GWUM9
fC93Jdz13QiDl/E02AZ0SgYDYQyMMCoM90Fh64dZSwn+az56qx2kLaP4FvtUah9T
ceuDltVc1vOuUOLY059mxPH9YsRT6dvGPBEF0eOtycr9T+YXgQWIYeCTZojLPKmf
0XNdWnC100wgZtmBIc/j90gHwixcV502RpfHNNlciFdkcBVMx5zb6+Eg4ls0pkkD
NYPq2HUJq4AEcJChGOXN04Sx8l//U4MdLSeTcq9ba4bNHaOmWiI5VNJ5INsPa5+a
bzA6hIb4LdSMPpyKlk9grSSToLwrWk49NSFXD8qDSv3rI/10cRS5ARSINGDXxXie
u/9ioqR9lxeFkLzfhS1aV87weCZe6OTjgPVuF3hgzdTJTzpmpTiFjB6NmMrGunZl
ITPAkXYnE1HKtjxtjxTM4ZvKRQHxZNgR1L5VFcffWMORASq7QTfm/tG2t/Z93H8q
USAyOWv//YIl07VztQGT3joInIkoApuRqHuTo5gOLuuWV2C8AyqkGtvASRP4doOn
FicdFIpsqYcLdc66gu/D8P4pgOtGaLWho5NKqtA9J2+kf+RGyfHnxerAiPp7T6s7
6R0etsAowcdHDOn5UEZ0PAjD+KmXi7uhsEgOTodmUPOeeN6fpHfA04a6rzY8SJaz
OCnPKtQpXRS5PC+EQu6CBQPgmyJcjbCKZ5YYcmsf8M2dA/tsgB1N+CKlojMXNmq2
WU3P8AAFyShkrugP1vfZfJfWPlFR7eFPXaOeIysmJQa59TsRD7U8Vuqzm9T41Qxh
svRiy1CdJqGZHLk3WHKIqIV7DzUr9ML89v06ihPjhs171WBO4waWcGCqdD1/c1uc
sYvyBfHwdentlmWuwJhwVwE5+XqVl41czBTRvDwy3K3ERKGdOgJ/3CCUC1Fic51k
eDnak250/P5MzpYfnjPbzj6V0vkKIOhiWFsdAl+Z7cVG+v+IONg4RwDFhy6eeEOE
idA2tJ2A+CoGSQhBq760NOGeWW8oNObfOeRVvyc5PEhvXw9bPoCy0P/U3bciVIxz
GbbOMZSuslZXE2b4svoXq+cF8QAFp61o+lRtT9Ct9OJ/KV2oqdRPMSXF6BxkdJuN
i/v7j5UsWbW5+M48mZla+glPAD7GLsdlCz8C1RRTWrPq0YpQdjeEJAFbpB8TiowL
mTQxwg/w/jUAIiI9MY4o0l6/Sx1L3a5thiVopr7RCA9ilgYMAG7FPnLhh1TZUXZx
8VlQQ2d4G+l/NtX4xikKnDVAtDZZvCYh5mwrXaqhxqZbAaCYmuw1Pmm7iy+tEQUF
I/WiWkblF7UvzEFSr/M9fw/2+/fRFe+FJC7FvOhrQ2T7Ouw+cQVrqIhue9eJFQvv
pS/ywDJTLrSkWvSy9rCn/rwN+pF+MRji1rB/Fyqi7xMo6wKWrb+E8uyRF7IcMeVI
juMaqf9NEZ9/duTsZ1fQB1GxGaGOL7t2gBMBlLtx3MeGZsRKexHJY/t2mNRqWdqi
RBdQN0w0b371yj8ejHOkmiZDTc9znnbzb2D7+ad+GbhlAXMPNfwj3GBg+Z7MTcQR
WovjDv+f8J6GlrrJm4CaXUjnltrwfXx3Fy5wAVfTzk344ByDIl1GcLQdQBsSMnpH
6/Pc6kIitjSusZDCVydgIMRjONVOQNkQ/F3igiFMzwzkVghCcnwg3fSocogprdtO
4fJaXn1YfVrWGwNB56nXeoEg4zyOwYhHQzo5v4TvT0BwKHcJANQt/k7iRAAs/im9
+0+JQsWSp2a6c/LZr+fG+7kK20SQl8WEtbKhsj6opOFAwzzE2+8wTJQQCOqMSsva
uNmLm1xzsG/irbfjLgj/Qj8u5SVgy8OZcM1+10eZshxn4wLSCddCosavoS785S9W
c20jmsapcqfIt8RuaWDW7spdaB+MsgyIQUX2Df4hiyBSG+yUgSZDUp/z8ya3YarE
P2dFbUYjGPziqPRj03nJ82YuzFqM6KTYa6Grz00FlzZ8lfDd3lRjOCtrHXBtL2Xa
ugtp/DIYH8GKHerfSQ50+04h3N3qI2whnFzr3I5QQHNJ2OnbZqP4ny0baUzuCv3m
Zbe9p9o2gn8NU3FBtGBaiT5CcaLa/6qoVNyfrczUIsrBoU3g8yKtta+g1aJBm8mE
I1hCq+7Chth/JB4mn5YYEGYDxturyO8siUw0lXwaAzaaHqDXc5ODFFtIs7hrD7Pu
3VG9JUpr+Mk/H3/6pGEWekPcE2QUKtnzGyszBBOL/Pwti9P8j0IqgUA7BPRHwxGY
6AOv1ZE2p0EQVJziRyR0yp8dYdS4BEWuoWY90LPfAYBtwHmIJljSFe4A52uOUpPx
YskkvSz30JdSLzikPyHU7CMR3UEzn697fHiTZeHvFHmUlG31SqKsksu9gj/NblEU
O5fQGrEt3xn3ZvUXwhrwwDG6es+SKWRgL0SABjZUusfTKjTEE75ipmZzteh++7Ss
4o2daqV9POleNz1OMI52fnVaHm97oRkTPplkrU7iYqs4p8uofLq8Q6mT0ztgP42J
ilQyosE/yMOm3oU39N6jiP6G7u3bunheAvlWyed0tGcsVeEVfdge1gXyin7+J1gq
/33zrtTdIufhWc0qlKAqLLlVJA2XtbRdyS31qTkHlbynH6n3+2/H3+Y00fmiiOZi
pyGI/NEDeD7jO25BxlQn+Rr+gan0C+11z9Kr+Y90QYAlj6QR6qsJZbfWps5AqBFN
W8GAseFJMMvbEMs8ewCVzXKYiSWaRJu/4MS/vIsOd0LKaQ+scWq4nKoY8SP2l9xz
hVh3tJ9C0CFwJygScXXAkQN7pZ7B8vi63zznM5q3yI6yhcOSUPhY7qqQILpssRs7
UY7dykyDp4EkNlod6VxZ73jm0VsliZ29lFQv4Ahf6blaOrOltFonfDz1/ec/xHCn
oBvX8M2rjkAwuMa67W4a1KJtUmBEKd1ru7qCKCQGV/korM9GXfhhg33kcA8WHppD
J30jcMWMomjXIuyDxkDd++XxhBTC/1r5jlIb7oiQY4Kz7IiI5M3TDPU2pNB4jPZR
EfOq0OkXJBT8XVRC5nMcCDTvpbyzJd4689YfSnxnh7XEETHZ7LgVZk7R1EpE3F/n
z3+GeB3rUz5Y38LKa9BFaEc+tTh6sbFjqNJyZ643M6m8vdAp1yg782h9EtSIFh5E
HJ6bx59RgQ1yGjf2hrvtAkWbolpPS8TDwb27jsMuptiSLIMoxCQ2AiJt03V/naJT
iaOC3kkngR08dVt2wk56Rv6rTbL+225TwYmkknpfq3jpuGxy2555Bx8SW6u/ntID
4LJX0LRgBlEYKedojKabW0qTa1K+hdpVji0it3b9vw3xVHTn2D6EhPBxMd6dNl4z
8fXgaENULMjVBxWmyQNs5XfDla5fYqfhWkzuww+byGMGjI9+zcQTIOFC76X7ZP+R
GJ/5CbfJxInoOcOncZ7FFMUJhXonDTlCXl1bIMPN/qF3sSRZANAy/CWrGZHgTu8w
Hng6/nRfAzJykwu8dskLmTp6gM6fwUA+PVf1qXIhnMVgcY3pjdgJsZX1z7DAuGUc
ZvEsrmoHYp0VmPP9welBjxOVlvOk6rh6KsPNQNjXm521esW2VKGzca9BAZ8xGCeO
tcG/bXXtkp6lnAFWjtrLj6VDvxqedJnLK/TCb59NhYb9VkGiPhT1/Clss32Qe6jJ
ZmjFhAfFZHBdVoqJsenMncJNl6IAos9kynFif2ZN19eCq6lWEFqVcb6vaQmvYeP6
6OjCP/oynbYzHKxCJSxNh5r/UQ9U3VjO/gOGBdo3CjNPbWoSt0eczoP02dssairq
T1HrTbbGJOy83lli8c+sRPPa/BLtKxOtxlG8U6cbzqMBnEbo/aC7u7XNTaQlJ34P
Nd7jUdToF9fe/7MjSClNnTAHIz1bkuykA4gTDLoauRFB9J+X3OoINMjVnbxkCumT
/FlEiAwezWTUQI0NZ/Wgueaq+pAt27Kht+W6fI/FU04sLxxv98JMDWyK1oksCRGz
cMZLMhsKDHOxPNRmsHFXQdNAc34avXs86GlbawDTmHAlBKjoeqLkQjYY0s2ONyvU
GbNlKbRf5UMcben/KE8DgTCx8I5PHNqmiO6dudHQfMVrzI5wcabtR9zVCwVXaaW7
Xp5xp3I/BszPV5mFyHjltoQSF4poklpO2wbLCrXeSwHi6jn1uZNNPyuzkO1+pqO1
k8gZ0fy3TCnPc3sXgDwaBMmx8aF+c9LUM97cTLYsPoqqKZE76r8Vi+IlcuGPu5w/
/ph4JSKcDyyMRBb1TBwJ8nVQgCNZlu+8/wlB7jnXkzr3zvPegZPgzjYDa+ttmMKg
O6KkBEV9pU8Qi1kjIjNuruH/kltX9gSkOEdbco9yRTZG8dLLuQIIGsLbzhnXXxax
EeapLOyDIvt6/vTcQK/2mQ1liM5DBsekKpA9xDCh7n8yovD9ggBr47Sl0bDk23H5
4qnIdHTaKOREb2dwPU2g/pooivpo67vY9ZS6f/+ZUH4sxKESFATS7oP8JRK7QlPX
GzCKwJokvMbZGu+aC+dPOwNdqFS8+vs379yj/v9ZmOzTRA+jL3MKPHe3gAWnh5Df
ReFuAPXeqdx2pKeAibIGo8efwUWrG0Elp7qSau6cvIlt0KbeI5QP8zsaOYjmZI1y
0PPm5EQN0QsXbU7n2jf3d3+B0nHIqEZYlDGWlRB0KYTawmgPmubDphhamLcoj+eq
6CG2EQk7pYdcB6xdaJ9u/+w6J9f2vB16fxW/OjyeQ4VRaYYBWd9AEP5emiqawcoO
+EkrK9x2FBpDSvFjTJp5Y/1oEJ5yr6oDLjiTH6spyyoGcflC4SwT6vg5wR3WSa8Y
b4kjEJNYCOLgxtqNdNVu0750wdfweVAS6T2HoezCIbLGqUZDFfDMa+Oo39s9h198
Ht9nMXy4Wip2Fv6uC+Xm6DwKEajYdSYdXeKGFzGc77CNkHVukYcvW1VJZm2gJBl1
HVfKrqud5bGXziskjvnsOniga8FDxqEL/MkeReh/YGs74t+SPUUZLIXVfHFJZTvo
X8fXEqQbe3cjZqYlCaCdHDHOvg3DzkP9NcnC+gjrcUyRLUzDzgERTYjUhaevizfn
Xd7bBCHSLOdo1YpMASulKy1c+UggQaGZOq/mdYefCN7ZzfiIUUNBLPdTMFk/BLKv
QCQC7XjxunzK4oyJX4gu4pUMDO2sPLZ+wux+p8LN25W426h6BIZgQUgpbBxIaRf3
0BhRu472/lNIz9+PgJwCjT+ykb7n8HLJYBnTv1LF1dVpL89gkH/kPPQJ9G0prBhn
oUhEUe2Oklp5sSYikh4jsKqm5xRX1QyA5CyzIGcsbdJEALbk1bO01tbZFBcxRvSv
WEiCrXLIVQ29x6YrOzth7NErCBEZedB4ZjdWZB+9hgVZTY0LmO/TXOHDHJqGDuyK
0K6HXl5SwUYpDSMQL5NZ8jrLfMUL33ZO+C/JUstDXKithwgHR56pJ7dxIpa04pGA
imoYb3wQjsVUft3v9MiqboKwZiYrFng8zASkkTydONHdnxJKF9EYidd8+dZKOEUA
3SDVu84YGdN8nPK+t+zbvqfhJQYkkTHoHhjYbBMQ0kTkUiUDH9K4wTo7tmAxWF2n
O4VRx6oNic8TJ/Ps0SoCcgMkLjFuBKBPk/e+49nZh8bRRYQGcKRgU+ewoxDaplze
5QanLtIbybYi/FVTjRCzLhtaZBliorVz1P1XEUBLhuD9jV2qxW+YV+UGiLFkY8R4
2ROQfIYYq+5f7DHyjUNDLh3u6Cywd8qlNIGsohprz8Kbgl2cX3UoEkHM+rim+/jF
7KBiortO7E15ogIbSBYLroW5RyyClyiY+/Xu9QzZ0qRz3GXVncN+jCsI+mKeuXd4
GJ4sRWRpW/tk5EBoXSeFcWTUceidNwBIkiZn7/DvH5anDnjR88YZbikmY6K/ua66
3svD1lJpeTruGFyeUtLsSyLh10CIuvTXSm+fZNYxxSZhVtpV8BwbQ0xHfvzpALBE
RVDL5MU2/nSQnSwhtAURjERxo+L0Tr4VY2/CIw12VwvVUMJIO+M+1otKFjJt3lGr
eKxalpWfJKwAVF2SQMs9xzo0X7tCZSzt5GKJNUvRsf3FJno1uuGo0h+I0JhAhGZC
/2qGj2l+KdYsXOxkX8gYdjlPRdMkZovJxhUSKeAZ8VJ6UluHtI+9OwqMY15EnlT/
xpJu7k/h72xUEiPHFbUAqmkyCzoupM5HHoBtdJel0hbTUsyZlGjznDW8HrqM6E5s
9iYnmrPxmcLT0TDjT+NfGByDFL0e9ljvods/tw2Sx8oMFqY0e/Lf0+sZalNXDeSD
NCU5N/xEvyHhg9AuhowTXwI5Tnf/woqTCGJO52MU2hoMkoc1B/BlLPyCHyStyDYs
FZXNyZkYP1vWSdu/dNiQpKCf3IVMIgx+XSIub+L/W+2/pgAHl0c0pdEa6OToGCZg
K6iYnwGLt7yIoXe7BCoKU/PubSU7pkUnqfkrK+UqsLyefiC/pDjh/T4wkcYxpFnR
jFg7kAYFfvHSVQ5ehtk2I7jB7fNgqBxcu6OT9N5BN9gEGXUIHVke5dDmw1t4u2jx
ArD0EUqFoMbecclK0E2IHzPvWOHRAWXfUcQ4TUsb96TZk6e03DufQAQ3jqBQdkOj
WtLbBW0JHK7xFc4A+r2LcTWwNIhyISi7USK7Eu8Q9jr5FUVK2EoVup0zNDsPjHYh
YYhpWm9fvlz93Y+gxP7l2S8xQoGGZPsEgBuLz+PEPtAFrQdAFz1mAEYhd0PbGY6U
TRS35EVQsZiPwphqtT6OIYXlMipu62HRUDzuOnPwZHiOd42BybfgT1nqD3XkTEGz
HVWKk1bCOdhR96UuKMace81ALGOeEW94OoNHKvmFt7hW1Nm7JPFpC46kFxHNKdsd
YrckQn5riXhkP7ihVVJeFSxOZZThf7jIvAI/jU00jWNl3ApMVQL5dW4ftho6HfNZ
O38K5PLA9sCHg6Ap3C92I8WmK+CTR0TGeGWZyI/HJ4Ljnxul5fjbQzGgWX7LQ7Dc
LXkVbcCZmFQTrHfy0A/U21sLCyWOs/CdxIl0uLKee32Osa7PSGquzBQ2CXlgLeD+
KZGjS1yi7q3Jhngo+t+O/qH61Gpznrvi9E5jQ7JTelU0i18xw+dYsu/HxwfV/Be5
YPMQKX1gbQQ5GTl1IH6D3+zHgk6n/CpqnDFePMqmgSG9YG70EWQTMFXGC15mI+jP
JnF4dyjg+quRo+GnF3INWdhAnkCpRzTRBXi4F49pIde3t4UngzY8JpLxpBi25U4t
IgZR/500CkbM3l+DazK+Y93Bup1s6E/yGNOtP0rk9+3mKC80E62X4GhxZCq2x+bW
q18ZSwbNt3LkbTNvEVVzGRPhSC7o+DLFz8MT6FVTkdJXTE8QRiyvMD6xWfcEXX7n
tO3McluURTiReq7tj0aGC9caDUZGAdhg7V9FNKYfl4L2U9mri05Xk0pCi6pU6ByI
CSiAVogGYKeKpHo+Xoc7ovUVLBUyFq+MeT8hQ7DEWvxqqfOjvfJbvVdX1bc9Uu7P
ZdEETbGhLwYgGe4TH6gXVAaADsAIRQwcISvK3Qq6Ykq1OzzqgEzSo3wABYyLRrQn
AK3bK3mZT4Wbv8uVc5doDqFnV/QzLB1M33+oPoo/1cedGq/u/tKtoYgMtm/7/xYS
WgvQd3doOC5sIQGeyHhFEfAEfkOiw2AFxksYec32+fKSLDdlnSstZCiLMFW7JpY/
/7Sgb+pm0DEeH6KfUlxVSM9mJILaEE8SuH1SVU0xCmO+JFwWou2HO5ILCu89Y/nV
Hr6WHJYtWRONCEBObuP3CpguzaQ89850bWOrc/eEl31jt5YGnWMKy7pSGFc2AQqy
Str/eCjxo2YF2kwVd8oESEa3GIJylnzWKOMF85RU7qpjQRdNbPfpTmE8VeYrLMrx
awQnXfOcmS7C6XlYJTmVijlVVLVuyHxt6dNVJaO7VW49dsBvtR+JSNU8Kc4ux0O/
5VOIE/vXUjABYsRoEVbqEqGzkH5WlEq4nG89ZN5mMCLI/8MJnHj+STnal3XGrUJV
tm8IKZlPORQOWcMPMPXslQfty+SiF3iUFHusIo4Clo0qPRIM8KQFm5iJ0IHUBHhF
pseYF5kbFUNkkabenYXvs+gDWEyxGoE8OmFSJxxo5XKMCA2carbWGcQs2yZ6Z67k
0coiEH1P/EUMlnBBFpFz3nyRnqYkgdVsBPUEXl3yd8p/bTBoWAnJj1bCfCUpYxwq
0Uug/X41Zf4HMaj/BcpssR0XhM6dRaj5sf7IMntuU0blazKX9d/Q/A8lQCZWQ4XY
5VGABHS1hMdDpV3eH4zcIVRlS5sWslauQZZkS/Qz6uNwYpHINGgCpAbIW4pbhAmx
nb/o49iymzwVd+ATXBPzulJ1Z9aSiE8LMOVD7P9zpCmVXxSXSKYo8O4Db53e0O4C
hYeEYnVSd5XXY8QrrYuuAMBCjbqW1iQhRkuPgOUGb+RLDY5aF6Yd5uY/d3wlzD4E
tNZlyfi6qk1YkX+O3xbzjhuvY3MhgmgI101mZNAVo/U+tn3XQ9t2Sx7jLEoKqkm9
AFf0HESe2Fez1XKPj8hOAVAfODu5uvJRzUodoA+Mxe0UfslXFy8wRMiB8v5nGnLD
ydhm6m2MSRFfMkKlprc+sqSvUdrdLPvzPRaxu9W+y5/QxjaHIu+Yl6/NtOI11p1h
oqRlWu2jqpRoxs7d4zi/QmrG0BqlNDJwqkAMvrMUnm72mqdBtRxsIZqF/qohN93g
9Tx0dK+Vd26JOVYVRsatCUCwCcK5dPQEUy5JOvngG5f4rNVDxhkc2QLYCK1DDSzV
HTxyv2Eu9jQ/FkjzM5WfstawiPlTaacSBcrk0t4SB2wU5a0phdEqh/xFgap4MJOO
n4cMu8On/9IhKRZKyczn92FO/TVY8SKXWvOJsZp9BZRzr7wceM4ahZDHmMgaQJ2u
QYggPZXCksTuD5R87zrrH7Q2jCHbeFQKgz/lqsoHVmH+JdlTryLYvK/DYj+cx6Qh
pSxfFGM0NkGdIMIGJ14oYoKWod7Oyq3/uA4d4iy0valXdkHhz1YHdkgoq+EUovT8
9mL5gSHlD8+wBiVOuJ8zXHRwxdeliVLLx+DydHi+uMrwa0/4/A7rd63B4kK3/PXs
cDtWAu0hRvy3U3nlllFQ/TDfExQ9n9tDjuunCzrGIJgRPj28aqksfORAT8ASJcsX
VJIkCHnN7rdMJX3Tsyg0EW3WhNezuZG4we6s+MdajreKeRibAgfcFy6B/Mpckfh+
YXZbQBaARlLF8qjr8B3PVfixGRfzB8ebm86S9mQ9eeFWdXmMWSoNBnQx9deGjbCW
Rlr/GaBSknNOQbooOnKbOmuLCj1m5Xure26TL2ExHE5BBc0nyUaP0QsZv/qYlLlF
U3zR38axarqcorFzdriUs2EtW4vD/4rtRvyFCRBh3qnzU7PcHjf4wHkpyiKivQf5
ymFrc+uojh7BTBjvaJ1OvGrftXdklLIa7ddWTmP6Qvy5X3K5Q0kk4GAYoNL3Tlf4
wk7Ya8SCKwSpO29n/Ex67HRuI/lyMwdMi5oIOaw/dEVo3ZoJMAxdHmjack0DtpJr
WY87CZaRPB+taXThOvAYjc/ymYUO+sqRO7rfyIG/6CqInN2FOWn5Wj872zRRGkYM
m6vmYd4g+5s8zzBgaY5In1zDDfNZo1rcTDqHYuZaY7ZBbNGJTJv+6HknkoxiL9Lp
7NUiuKHdqRNtySmrPN7tJKYgvYmjAM8Q4SvGqPRa89otL957WIbyH2343l1VOTfu
6VzYduRCTsMF86daBVJMCpowGWgubA7rJGWzK2BZ+tuEm8wnzAInme+65IhfANQj
5QJIRlYO6AFR/FkK6NCqEjgOhr+d/ruK83bwaAqW37P51kbyD1Sw32MPwmfC6g6H
2wKNjl5imWTIWcg3JuQa6yFOgOd8Lu4C7C7G0CMVbywTXd68PpM6UJ0p5YFeCw6c
/YFiVslnXkY6I3QNYw441xsuKmpaOnAzrjul4RonZHsor1E+r8rsJ9Nf0ZNWx+Mm
Vk10gRyJoSz5tExGXIfTQs+od1PDhqjhD7id4bCyCD2elYkArYyEsu93e37OMaDH
NiXYgUCUaEQ6PSxuj6dnFhDY1sU5ZVz2TS7Se4zhW/v5q0KjPR+RA9Y0iTbTNodJ
8d8zcUPpd6owFPy1FGIe+lUe6J+mZ4Hiw9Y2M/zpvaqa3g6KWrX0rCPV/OfZgP2h
M4FV8F59O37dKPX6pleBvSFafFhzhgmRynk5kCFtQMaIr2v34DdNQXE8FFcXbmfz
/PPPNSyOPo7lzbYcj06sFeq8/bef3rOhbIUstuqbVFIh+PBEkspt3qz/TXD3Wxk7
DZNswAi8RgRU/4qYfGzSnhA72iyOQwDvTNiz9V/qt4L5N/YaR+y8iolFke3mE18g
WnCpHp+g6BExk8o6lKJ1oJvqRnMzjYwQDuut7VhndlIY80gAAM06mLzuUyyG3SwN
X96kzI6KMwjr71fWHWXQQ/YjM4Fr2d8AeE2njT54U22zx87DHEKPVaLkQkOnNBWe
JCvz0mnb4dwllet4nRlToOtyeg01J6qyruc9sQyy2q3pfyYgXx1Jx3jZI9KQaXwj
J2j6a/N+oCn5F4pCrXmCwpecpypVDojAxS03UwZ3FX6Xpax4Giyh9kQZyiVEM3mN
7Qt2oAjaG8XcFoqOcUfjouDXU8SuCIBwxvR3+zG47ZdXF99cKXI5pO4TpOLQiO8E
mztDPrbRAqzqLaUQqI5qf9XkK60HRhxNhgAeGHY5vQ5dlWmqS3F9tQE68LmvuvbF
DEibj/YtvRIfSKhwVChM5KINhuAMosYuQDHF2ZGuwpGlg7cF5RcR85sT9EkzALcu
Yxm870bj/5Oq+GWW/TGqahe5IqYq6yRo1FxCb5D8HJzynqNNZD/w3QVaWUgrF3uV
m4DjLZ5XwxWyltyd+HZmenW4pfGFUusoGREJ3dDw784vKM0xf9Ww7CV6ma1YrT0Q
MygmPnzZOLqgv3m+XmjCwNLlzMSpl8gekGsDtnqHH9qM7P/0OHEDv/FTU9gdpbPL
Y3ynz2PGOYFik+xZLMkKZORVd8RfyTieamJAe6uS84ECPw6luxdF5uAfrJ82J9ba
t08W4uJfuPmY1mcigQUDCEvZ/WTClLrmq72SO+RJGhL4bT9w6Vvc8YcvVqxiP8hh
avFsym5LoE5/TpvK7LxhkBXLCyIs46UVIuaCstM+C8oYgrbpVjMFH17HyFyl977n
UyDbj5ipy10LUVViHz3H+qSgzKMTQftJIGLYni+ur9EC0rQCmAsiEjj3rcJTikuw
IPiOmbh0/ZjvXrqalz+pAkqXlYgdj1JcHpkaa9bFlHb6OUVdkU5SHdoNHGlOFx8C
8qTRyXlH4PcXawdcWH1TJuEnlVfbMkl9KB0QT6QgPsAU5e9m8C6UbiEVQLtiS+xb
Pv4BapBQozdcqgT8kdTWBXsGLojbAloYRJABPA70rwu9KXwcL9A+IROtoC4Z7U7D
gSqj0yq7NG/EymHCjrehuejXAWLuEm4De+G6VF/lj33lmZr5tIhI9YuHFFDXwrNm
a8Oiz5ODvd8gVb/7aprylet7SCG6ZZA3tQMFiubH79QEHjpQUCRLmfg3rAhzyi4Q
y/orrS2jTrSiH+mb+SjG14KU50ld6jjmeBTlsm4o2n0GfPMPgc1uN9Q2TVvoXonz
yMqxW0FPG93zi5ExO2czzhNVkvFVG3fX0/TR73TUhhpw7529SwF7qjKoSGV22Ytj
clWWiQq94jbvGxlAlYZyFPcCiP7lFX7YuO0MeHHZNC2QXk9ZNriXaxvJW0lwlxeF
/01uMXdsvNarVqrj3KHQbrb8p7qgDHHO+ihhn/LO6+Be2KXBwl/M2vHk14tN/yXH
A+QjxMeOa+j9Js/b5ZliDSh5vx1ojE4fo9jtsqIuORzwyLbYrju5Yj1tbyo+r8HB
r6BQ+Q7YBz8iBHFvgd7LBG+rY+R2IvRb0mq/ikphvoGIdEpvJeEyawhCNtI3K0YH
35A70GyPleotsbA6jvwG7hEI+D0Cnh3rsOo90pYFPagxwBN3m2Dl++orHZXm6h8X
lSOAkKlLHSxHvv4Xtd2rd0SfXJGKNNjlw9uTAVAjC6IZ5kSARou0ZrGOUClS0fs8
Jhjh0GXYuswIqbQ878SzVhIVUubctMGYj4QQDBEL+sheFBOxIowvkPeD0jx8kqWw
i1lRMz8enwipVxBopnEqGgrP/8B/P81hgeLxPKVzsxbLAXqZjIhrUFB9Nm8ULQRk
VCkXTAILKzbtxqY5Zv1dk76BzJxDLLpQo0zbXsOz7Pc/IFAqXdDLXgNUfA193027
Ih/aP8T3Yl67ZUdiaCojGSwUHYSyStBxjgXd3Jmt7iN0MgLvS1499VUZ4FuhC/0V
nKmizLVjcInRo2w//4mxYd6/mc5TMKwUCia8k8VyRntneysF0UIN5FXNhWfpR96t
5xTJi7CMI+GZRVJMKtxf4WCecTMRx3UBakMyrD5kxSThXGPrlXLlHZ4BqDauGy1Q
Acjukj0+OCDAE3DKFZgF+e1dRVGPL/32aspcAzu4mK4pFU1QUTk/8vR3lSO2Z9Tr
BtdWwVWlKqksnbLNjHsTJ9Pp28YRg8DsyhrcFk71dBv6so7kE8sHpD9cOIyJR7wm
Xo0xUPjUAQTJcKQbQs9G8X1dS7wDA56OT4WgafkpzZvFNO0ypU/Wu3Wu4J/CsnmM
IuGehvdFrZypCjKUo20JGYoc1b155h8syOuOgNNbGw/S+i6h0T+wWAdn9nKzU31z
5wIpqYCbeOWQkRnKWV6OaKnYge40rn4Sw2SdBxnsWH/S+t9wfHo2fgaGNvuIHIhF
4f7J3mM6KZYMjAM2Mf7AhIWeugoO9dXh/El4puquUwZPp60KF175clMt6hZgHYA6
j360LRYzjCyKsrixKMsoH3vEmHJ0NgxwW5yxNEWOwrK49TAOjoqtRoss4xct1gzN
XEdMwNBsdVsSO1cSJsKF7Sy3CUKq02ikSuI8fXxWHFnRQiDvsEk8NZzVzkh9vPre
/h1qPZZRGOOgm7aogx2EOXPs2ac4Xd+v5GjhbAmQIt6m2uRG9UfExt4bTHFPvBYT
Ta95mhufrlqRIz9tj/H42GMcB9SRwDVWqAo0Jk3iifFQrWVCxNjlRJPAiDhgpD/i
u5UQTDpGKeFiErKp7PEO8s59pOGEn/iIbpD4TirzQzU0/Nv07FTucwrFEIV6aHwd
ghZSmNFyVGp7rU/NbT/RFa2F1cDzCLrtTreQtu+qil9+33pDcA+3sswx97lz2VZm
Ki0ZzQphJpcMc03zFEhu/NP5zr0l20SvOx0oGcXCXTI5kcD3W0E15/EdWsubvP2O
oxQ1AZY7lk1bO0a5n6l7s8i7baVrGdjD17HaOJj6uwqYz/haoSyVy6MMWbAWCGUc
1oWHVQIytw9TS7kcwzNP2YiHfJabEZ4xoIbhhXdgNDtFJNeWJe9UwoXSaQJSq9Yz
RAXRpFrc/XeRKQ8J/zIQcIY0cnNU4RwAEJZwGw+9vNtr+W5JS3VlTa85idX51yRm
oPLcxX35QIY7Os+uR8jfdwcxyWrZaoN9h/Oncs3c6Ah/1yC6SdXB0sOmPqFoXJCJ
8ipNhJfqgbQZsxDqV9lKVCh0gP33AeGTiwYi4UWDyafc/2Q33rrTzXnFLPzOKPSu
NPdmXTIHX0N6/vlPTK1oDXmkCq5ji5g0nUx14tJGIjICSm74SgMI++yoIWL14pU5
n0wCMkCMgzA7IcxHqVNtwP1MrbSb2kGPiAmEZKxQa4hN4YRvwjmSdqk2/OSJp+x0
RRMgRYd2tUS+NZ/n92Av9qggq3gjcw4P/YScuTXV2oj8+PTeES2PeER0LUG09d2/
s4sfwhZq14bt+hqG9T/bN2gldi2BWFKoMn6khdIWUfigxHXgwdio53xB8b2CwgAI
Y7PKWlr5C8p1fS6qGFrUcM1viUDal1u/7CbH6f+DNTcJV0mdgg7TPGv62vacyJLH
1hxcZBM2LOCVfvJ1A3hwKeUR5DMijVP0HesrHw6oc/o6HA+L9KaQAwMqMXn6pl0V
6mxQd5pKJIVQdbfnLgzw84o/SzJy1/AcaJT3+InC26PaIhSzifb1YZluvkr9Nrmy
73l+BWow5OBE0trIeLJ2DIAB3Nx6xbpO5SJQYminNq90MLG9gz1ZiF2yNZkXmaBn
NM2FNMuWAfr95KTMmOYQ61hm9ELzsbCXI5U0ayO3I2XeHvtNZz6Z7G3DBGLKj6gV
eQZsVvLYBNj02Iz6lSki/fGb+zRNl4ZgI2+g/2Gp3xjWBdGiDq9e6Out3v7E2w7b
BJccLCB26iBlYFB+Y+A13FZpH4tA+b0TfmHlk+kz4RBc9862hdIavAPmSpcyMLVo
EEBlL4vsOKkn5f94V+VDojQY4wzG0AR5GPwnnnOSMaG3uyUdzAKqnUvKsiMGuUqo
99VPznxlxb1cJqtrH2z6RUrTisxiI8L5CZtX1xt3eEnDTy/1CXDrBVxDad45S56Q
NknNXv0NDtWKfO1h5WLNlk3J5Q2Hch4hoclLa/Npx71dWhXFIrJ+Bon8t93+yyDB
IKwVj6yyp+gyaaNiIyH8LPqPHjcJklx+771yLwLuVpDNmjJ1kUu/CVv5F8RftJhU
+kUdsKuV3kNhenUkmSYYYiO5zLHTsVqwFPLQIKskSluVdvWTpn+uy+XmxsSBKwWE
R6gphF4od11mqTSg8Pe7Emnrd3guLgD8367aUHhBEwK2UUXMP9HFQL9FzywjJa2i
fT0xzR1Yr4PuQ216hy/cVKQvs3Z/CRHo0D8y4+kVnkbGK7UPJQRiP+M+/HnU88Am
z7iACmyY2zKViEVuKZd3mhVhtz+lbRl6qYr0k1tH1OSq/zn1xZreZXqoKQZBl1+t
mmhrtvpmT/DkmU675WajeM/28bWE8GLIbyhFn2+5aG0n1V/js6jtNVZuBe4yY3rT
5ISybt1dcbCw7jYKajsRKUgA/oXuw3X26DEfsHl/goMvik1IfZ+aJRU7Vq8ppBeh
H/phnnkw6bOWFyq/0260Fid9i1tlHpaoEqai9e83DHu9QpZ+hHKDPf/jkFgwHI3L
vRWGTEPO41wzykFDAyYjDjDkCWPK1Gk57n/eh/fgMq0j9yI7TkxG1oCfcqqGOUeH
WYEwrrS5L98HlWT+oRtH+W1ci9wAeHmzgLckolorVFvPgi3drTZ12FZgMKlusbQY
5OWyW1BTfdBiSBAHi8dhhPuyR8k2r5CLaP6JT8sJfMygHQ98qS3ELXN4W3wyCpe7
riF+byb/I3bf8oP05XL+rp9n7iNcZInc3y+uSze2GOZOd423huymWu6idDgLv5Mz
kMjNlXNOA6duoOm7Zir77ZPwqv1zm5ukypEU1r9QRuTgRJwEx74YuCJ4rbmTt0sw
6R24BlAPJJvihuYg/YMnzsg9baH1X4GnNg1zDerPXAZ7ZSqlRCt9/5iVVvWsFxBA
sed2kSvh6eu4t1SfbKr4jA95pGRXoZRVkdGnssCKyk5PLhj4EB1h7TP49J1y3fP7
OgCZ+fv67MQjowoyS1KQ2puAvCE6SChNIysOqNEVbo59/9mY18H857seplEbf7gr
Yz/qCUAV9hP19cNysnbHsdS1/d7giDKacKFD0S8xi4rerGYn3UMk1PcZ8sPc8z25
LTyfgIWg9Gr6VnCMpI/AQC6ezpxq6TjCYP5zJkTHRbFuinxs9Zg3erzPKaFaILec
e/pYBt7kHaJ/bBgRkhNEHuZ/h1FjXgGpYLU3MSvePp3yJN4xW2x++q9wWxw55uT2
G7UTEW46Du//IsP9MTGiBqlMgvAJ9BHa0uaGMAHj+dSO1160FqBhtum7KjD0/lx3
prj9qAwGeA+rphcPaB/tQwoQOW6l/dBDrDtWNFS87cEY4kyjC5/KlnBu1g6+iJo5
BGgqP8YbHdieft4PcT/lR+J1b1L/P/KL7TSCeNAwBlX+ckD3fDxGmOSYg9kcXeJa
E5NlInDhlsDUlP33NBxmDPBjlPsRkZYDiTVgdRzV6AkIR4XfF3qX3nmiXgO4Hb/2
cXYUBWD7vSabd2bSvrG7+j4kmTNpHYQhv4ifEpnY7dDrWVc1VkkeCLEnlWcKPX7d
zMyEImpF6n4/UlJYLGWaHJcYge40qc4/bE/oJIX9QGeXi1XQiqsWY74WQZvnhIZX
Ojgc/22pyPW2fbFD6wmRWO+ctw3kvVL5fhghZPUjx/w0P16WT+Aj0aipFl6FTI9e
c48eM6L/f5aUzHWOwLYZ8APJXSHOuhwhUCrzDiuxKzBLLLViTrpAYTMbVsgrhG8N
oke3HtL0neJTr5k4GoFaj+7BDwG/u/za5PIRicBQrMnESyQMvXs/n9EwwZMeyQV2
LeNWU8+robbMpwQpIUL0ZAke8lpEKJnN10s/SD3w+1IJzYFCSE5opG++IkrRvSdV
2TKK3hgC5NhBSi8ofIgrTGLoHtn8ytUH0tPCaTMZhqB2bB64xrw4fLltkwSB6gUw
fVjJ6sCpPh6Z6xiXPwoFtJwzhDOKe8dlHxEvjzAydtMpGmwt2rYk804RV6gzTzF4
jPN9GSXmGFlMkhdTOQGJdiwYweZMT+vYYBbPaGrro2b7eQF5vEIlOPTiR1W/wejU
ACnHn4F560KVv4d3v8aM5ZZKN0PsHdjen1rI0EDhYE/qI4q27oyThQ4XShayWw5Y
SmoFniv4ct+hLINKzI/XakNgylXm94AHbIQnhmo7rRxLQywtzVlZW1F8Eed4Fjol
di7A8ni8GJEvUAgbH6iqVMkaC4JkHJSwRBckqG8FOYHrEuORUBvVIOEQ2mKAQk9L
US/+aFY8QxM5QGOUJE1mMbzlglxfCERWNhNWD3iPGmc8TiCDP3/FcignRcXgkMCo
SWo7CC/D3cwF9nN1oa68OlM7EC/qK1nzZqGTU6PoPQR28AZ6AB54YGdNnrmaX6S9
JE2nfP3IGSHoWaqZq7zGc/q2Uptbb17hQctSedQ3WHxVMWmgTIWN4G9kmOxStPJR
GWWtCsA5ArMGbcFN6/fwutFonENL6K8lUb0aKjEIhJWdSa0HriIJxyR8F3FuWNme
OpzvMnRAXHZ0MlmQzm/TpEEEWN7GHyhIxZwLuAoL2l1YuW4EiUXiejhBaYzAhnQy
AKxHdM8R+NwK5TZWZ3eECp7vkZexW3Eus79FrWF97OiZuUDQ4MOk4NaVLoKVtG7j
82MrxdUpyeGrQL4Hg1IopijCQdwl1JnHbj0Pj0Exvl+V1386AjWi93A6lk/4qUmD
T/ztro1VO1PWLtmwyYvWd1DVdIhgkF8aBlt7HI+aG7POEDKRrJb4zWgluGdyiDw7
O3wErCmKDcgld1f+kRRI9D54wRTYDZ5Drxxqqn7GGoJ4bseuzROKwdzN6U11CUfa
1mey/OvvbAE6rxiQklUWCop59KGW7Y23bIddT8sGTZllnOM9+Q1xDEKO867ihdWf
sfhK71DJgH7s7DNSkv/ZZ+zECWnVYP3wJbJCm8GAaFzPthU9C6v0J4+xQlV3zPlT
g0xKpZo7yxKDJ54ReUxY/7jBIyxR4eXH4hSTsWc8ZHoi2fww8YyQ+f9515YTjFkA
gOBk55Jj1IdKWFpiXhX9UaWdgN4Hk6sRgSCjMRCcUnDBAV39jWVyb0LYSu7eIDC6
E7QX6xZNKFg/0p2+r3cpSJZfw5ixKTlaNCyz4eN0g47Liqbv4pWj77ehJ4ZynqiN
abeSGuKRVk71R2ua8D1xz4ddWf+x8kzo50ffvZHKClody4jO68ned6ALQMwjKT7+
DVv2VqIVotkRhJU3oiLqs14BMLwNCyyh28TyfKZ9zW3C5f9J1ofW1+hs+gTSug+l
QuCtArHCURX+B0I73IYSZ+lmIA0GSQcj0jlgIoV8wC+zyyrtqJCM8YIjppuy/e54
2HP7Dd+YEb+70TlNmK6OFM2ReoWN1qlXwhRyLzb4FXHfu9bzCFQFF9UfIYX6wTNz
C+4CFNyRdrF02tgNA+exP3Xj9etypErwYbUdWT9mSCyo3SZWjznOdhCbyAU5ceLA
hMyXqizLkimztSjNT/NVmKWaN7WufOfyYUzmPKab9uqlvrlEV1cZPUx+REuGMV+d
SIraSrCk8iJX5uvwub9CAsJOeNXoa93CuhSQ0g4mZBeAnkSXSnTPzIXby9Ijuhle
U+5BsXLzbThg0n4H+P/j2ljjFOiUAjdUKJWQJV1cNwXPTr0P1BHTLw5+ERePLFdB
1jaCF5ymScdvh7A96pWRhnltPcbjjomBfOJ7HduldD0dASvPAMxOTDLy/PwLSfXK
13qCqOGsQ82cvs7RVUs1jQ17A6m/CtN1Ked2cHTtxb+Tw7mlNjm8UH2Tpnl2Xbip
kD2cUzoL/4H/1qSjHKgTCXFDxpFlTButvIYZFpxw/jckIQwAXhL8iBLo+cZRKC2h
6MgJnfrzogjU+gT307jwb/3qouuSVtpW5MKDTNQ9ucymvGu9b7szHcikL4qS0d7I
R9IemrNpaJj3uusriDLCpzPaliGhSsN0M4VRLEYzFFDB+Wpmo9+NUb/CUQ5uTOUd
6xy/MDelEE7771FPAo8JofN0ZfRWwlIlsCqGd7HDStpZ/J3n+zn4mkPCRxSdkxD5
kVTNVjAMg/9DZR0x4YQL+tSQl06+n0sLLdohkvdMsMrSGpv0bTWyqKkd8TPDXj25
TdBzSxYQkwjNfn7/YDSUQlPz+3E0n3BlF+Ajxpn1YVTXceGCmdTWrjZNkaa0x13s
NzhzNFs0CPsA71ScwuWS+Cg96MUeqZZUnGHjKtVbdomU6LHpLjXfUD80ewK8rkct
BLCBt8sGTz9hpVjK7vmHw8ndZC1BUj4TmT67PWLE0iSM+QeF7LkiompHA0c9Cq7s
oCQWTDP6JDQwL3E6+wvRgUBkb0DUoKzqKOsS5/o1yhJ7k3z6DLMzYgn6aNuWcfL3
l+uAvT+SBPWruLV2TQXxax8RoUE+PGdXfqznOEojCY2xa9TrRRDTdDDIc8frW9gu
K9aDZsgM4BD9nsPhAHWpKSpld+imnIPVdEGt+Hip0UWFhSVpLtAT7LoLj6sHIbrg
ETQJOEGVmPFQCp6k6F40c/XcNAKPn32Rs1FeYY5EFJSaLgqhBVbf5zfhxZ0kkGzG
ghNXD6JpEqtplPcayiJOS8WStEG+fd/+1DOXJb9yGlaoBdTZhjBy3cEDwcp3T5jk
IYe9D5uEEe45MAhDZ5kIUiH0n4rXW53aKkZjywvy7XvSJqJX0IodrKx+SnMslKtM
GvEPMchZ4hr/4Piwwt8xX8szQATXrqEAbYwMoD/K495JWhWcxVNFyjpCn/0xqTza
932UYVnAyQNM1IgQ0P4C9/E5dO/6l4vGgSucfTf7D8NWBoaJWnp/6hE6zNS7rwkH
3BqYZNiySv40L677ovlZmygUWm8cefYFqQXNW2d+UWv/UhRYC2DN8RnVtZ7GG/5v
ikt3ppWWIgMVltl7ttZAcKM0bUNvWUVcmGoSr5id6Wze1bFl3hxLteCmSvShb9pz
WcHt7JC7fsxAJId7arpKtrHof4WOvo7KQButQ7fK+3mrTNf+99BAt32cXi4NzQy7
/X8Sf9Jsi5k8eHsfd+4cD5AdV/8sZ+GhWUznHZD79Ni2ABoVH7uS0BL2bUCI9rzr
GeD4sunHidgiKUAtFDeqiFho/0AwmqS1rlCEEL8583vgVQ2DZSHGhrkbETWl/TgZ
+jcQ89+uV27Vx1eeiOGQByHsrJbgWG9SVNbvgk3RYLdwP+Fq5FluFvP0Dc72m6wp
vtz7EtfbQYStogmTUmCUvimdfspj0eLnkMnMs+5ion8dTUOieSP9n6qwH9IoQ5CA
6KhJWlG2Zymqzgk1raXVK0oI0shjPwbkU3uNxg3aSxcfgc6NxR3j3rYq/9KwgbYq
p7kExPXOIgHgQz9t6UUtAOxNL1TctrXmjxkiU+K68ekxayTdSc0mjXYjUF1hMxW3
/U7AII5qH43SVgmWAi3bYu8PT7nlbFJqphrZNzvBnvwb2vTUjO13vVWhP2KiTcRA
R1ifx8ScjgFSZrBj8vBt35yO0GPyTo9HNwMuUGWEo36JIMPU7wScqN0em++tWwM1
OXEB/h1mIEJG9AoHyAfZ6AWFXR2hGnStCc+cmw14MMTQfp2GG/KIJohyb0fxHa5Q
QQDHOM7H4RkhqStxGRak5NJTPw0ra0oazPrRQnVKhsFIV5+Q49k0NWfza8FI3vv6
ofvC3ujcC9pWVa3qrw8D7S9hC1HXopQJy9hrdgBb2kVgGpcRuBXnbweVjDAqNSeS
G+sNLUrYkdXRaXJhsIGiNmI2jIRC+TAIJ10QUUr20tafX1KhYbdM3jf4wEsSK1sq
ryhnADu9ldS7M0Lf48DRhGt5GFEziPL74iYJ+/rcAvz8S7mxnmlS//KFZR7jrhE9
IPJ1R5W+Yol/1AKXrPWHU6eeNz9dvrNlssnDrIvIw/dG7+5vZNQAzqBKeOMSmTbD
hHqdPR47RwJUHv+hDzUxQgYtRAd1jJtRTW+w7lLsONTcPW4R7l+7RIL0m9k9C2ft
p4kpucL3e6a7T/0c4fMG5fZwGylcDSL5TPhV2ssYdqJe8ts055DKBq/XDqNUSt+x
tR+pAu/+lOhB+w0aYZDm9gfhmBkhDss70lV7FXbShb1OjQvMOYOPxRqUqEV8wuJC
ErAmzM5Kx2rYHLAW16ekahIvB5v0+E1XO02jxcRYJWTLpbjdMmR2Sriexg81d2rL
64GTaBAjJjSRKRrX4z8Qc+4qiHC70ERkpdGrCdM4LoPO7fc9rvGB+P4EJGizb+wT
y99S+DQGPs+LvCaLQ2dmDF4wdJu8OfE52VKeAoHPj37Ih2XIA+1GfAtgCwTciuCD
4FG8OVFyH7GX1JwlspVtB/61vqnMdriQ2Azho0XEESbDNA1B7bIk9WstakbSOTRT
pSyM+fQiPn1pBQOQ6VN4qu5jiQurzbR6OH+b7QVmN6xQ4BCzXHFhXz0ycoqtv8Xv
uuwy9zeoAB1mYHNt1e+yToQNZMr8eerkhZGQxufYuOWS/DQCNFgKtOwjQYGx597A
x5Z4n+GxvFCtqptroo6Sr4sqVubKTxMtBQAxBrGOkaOan61TLVkYIVDGJHgiPWEE
kVYgPbvnYbG8OI2iSv4gibth+Vc4nk5+tOTUT7MbOr/IZU6El23efMoz5i+6by0d
BhEKq7IGkmMVSpUEECeTaPocxtRYPqsZZB35v8OLBjHi0t0BF6BsPzbklxpVonbJ
mxCzeMuI4GGj1SX3WRm90BMMGR4ewN1NyaCUVc09kaaxywpImmZDhbgjO7mvOADq
4RKFKre1QanTet7wWmwmrCyZylgblvnhKGMZikx+pLIFQPz6m6tYWE3+G0FZmLI/
Q7oWu7AVXgeSHuTU97OcJHHYHnbXG6bQmyoRyj8ZZmg08WLBnJagULSCL1SFLmLI
78RtUYIqsBaNUwxzwKbmQnNG41sWh42dinW3yYinSgyLMX17Lx8vuwlzPVwWQi/Z
sIq606z+g9vz4OEPT/PcvBys7ymvwY/rGeJj6iLdPqSH8WxB7ENdrzdgkPbb7S5i
ZjkkvskHrCHPEHjCIbHAb4FaXW8VMI0yVuaLs9XqSspCquWhFwwdxWdsNrJ7XDuV
4kEUK2y06Sx9CJDORjMGkSKlxkd6g0HsmoCr9HsHG+wB25GzlKhGTUNXVxMDAe2l
NobxHkYLQBndHmYYKrwuloh9mphwEikMn2wr08mEe4J9WVq16XuyjjPOj3gkQAxS
VQV/6LIlw2KGp+Avo+IxLcm9TSAt3wmFXA4BkDyKAwV93Qq14E2mIrT3jmOkG/Zp
7nr1GyRHhUxtnVtbXlOv0yH55l3lt8evd6oPluHUGIuEnLlKRqKA48JD9bq71Np/
LRnOtks6JEdTlrAk32zahApQ1SiR/PaYaKOhFex4DRj5LBJMAQD570BM0g5yMIir
4humIgBE8zMZxv4iUf6+DO9JJPXuGQgACw3zpZQJpSkjX6OxK//2gE5FuvHCosMr
ivBtWJkTgq/dPGzDaCmdXAROsaWtaPnwkXbao5OKAnKSRm6He8hDMCM9RxYGsUa2
MVcW2KU1VLzkk1QfgOqzybAZMANpmjQBZ8vqjZH2hCpdKv+T5zXUVCSSiWuyAq4S
9Uuuzma9Y7TYWwFir9gxv3pLjRfOeT6nyLU58klEVR5hIARCAK0NDzdOHaVrCKuY
BqlrvbF1Ct5Nbp94eI6yQs61L/p/SU2yorxnEuszFmNeyAH/jbhxjuRhRlPj72XL
6FgM+30CUtOWSOK69zrSbOVbIvw2Nhwfnm5gUdX1iNITmVbNBLpkzaKLCgTaEvN8
NAq4MWXWmg8UNELlyj0DkLAGcqyIU/ZPLjYMtZcpLHOd48Hhk7/DACi1B++iNn7F
j08w1DxkDXkpkWa0O4JfpopagAliVu8yG6fysY46dYsnnhZOPK0vfXH7TkcEvZL/
Msr4wZ+dkCQ89/rX8QFT+rW+tmey+Ir6+pH3ka86HGUHOcq/fu1UJ2rqRF995nUi
YfMHYmuP7ipArVFAHe5eQFAoQGm1J8rHDJIQypwwyuspoJ8boMhykl9Bmr5Mk+Mu
IoAymmtnK7VHzsO4OBZBRMTnHkcFbJ8iC0/+mXSf46SR9sKdXEA6gr/+V8FxJyUj
l+vPuCZZrrE4SpVzYZTI0CCcmUvHZm4vkApM14/jBbjt9rtawwwjMMq+Lrmfiwe4
FNx9BwYO51ob9x60cSY1iGoRqqw0b8Mob5FoMa8Kg9b90NgJMRqhHr+yDW1wm3gq
mT30CgDr2a61SDmZEju6rVpUPyD6okFnsUjQL3Z+rTd1PWLzwAMSZTxVvF2Bftfl
ut/gfikZ0WSlOLEsnP0VAEaC3A3jzXgOWvGt2O6UWqNuTw88/0HPYFfMzInqua8v
381b2b/MCUcn4jsx/cCDM16XlbIcOJVBrPCi0sqUC6kVk7FJ1hMJeaSf4cJ7OJ9T
3YgKUuErWDSxssNzep997fnrJYaZ6vASdFt0LyONgbo9EKqgUInnbyxitEf8Ks/f
O4BhnG1IWNN1b7tQ/j5Ct4sIQBnASCZEPiYzMXszS7Ew8gNG6T7EcUCy5PBFEdlf
hDRSz4UJxTaQMsTPP2H7dvN3Ubi9VZByinCeyu97mWYeiQN8HQSaqMHEMODS7lGk
EUt/QQ30sV56x8o4/DF/+VOotOmXtOtdCQr6MKmJ75meFiP/5BobAEokcIFECFyM
e6KkntUWLcJu07SEYP+r4QxcePu6Ds2xStHklIKC2B+eRBRaWcLB3QJpl4pPjpOq
UaMJu4yapeFjwitea2iCkCTrEBoUP6FFhY5ozcvR5b7B8ixHEwGirZtXIwzyHgXv
GCbuPB23aJtO+1HwK+wInAeN9EKwmJi83jU9C5+Z4maYD4soHRdfvgXujtkjUtnX
WUfs7YbsfqW79j3RFW/cmcXDO5isPVli5IwXLJaQHBsiXswYOjQpbSZIAlyWaM0U
SiBGcUp5brINcQH3ZIVAQtvxYEuJO8KcI3Qo+4+WbFT6XWNZafVdXC7r4pb4JbG2
C8g8xxPunRVBfjjOe1qVcYTg+lxj5uZv669cP8nIbBc2tL1+KJM7VYw9yaTp9kfI
uVLgmDfRafRI5cwox790yb9siVdID3p+5zobsjSgFK5mtjyWNYxBTPtNRYbO2n95
776CEGAN6S30dDWCZjrZfPUC0a/+VyF3LceIyOvPcYnbozNVweVRB44A8VPoh69s
ECPl6EzY6Z9n1KAwrgePeoMAp756WcIwH0v//it8zOpezCWQBxKtp+rjlVQgGERn
TEufwHBt2DjP4AziA9BanqLnLiaMGYEzbP1N24MZqs/cyDf6aK02oMXFU4pHEg05
SGWwbIAOlal2Fj0X915ZnzdzAUt1FIARG48yQJXzCE1ZimkHQ02upEqkAo8qk8c1
laM8+zepGHMq+sWcXlXIsjqHJAFWkG45NPNq6i1nCTGXmJqaIdcNtht5vh8Ln9ft
7edoiySa7NENwkzrCd8DcaRQUfRWmD1pjVAH26UYg74f+hJFTjaBY2T0K4CeNY28
FWVAZsyb2vm51oF/eEWE9e++GVN7B32HJxLbKyCCeuuHsxRlF82KQxQkMLwLt6dM
YL2rf5dMgA9/n4EInqgxmP1fVphxIMcdpG4oaD8sy1i4BEDfVwFx+fbCNDZns9GP
h6Y4W/GHxW7w5eKc4Sc9r7p0KHCTX3KCrY5DXq41/zqp/L3W6jdscDrpX/ZdFqao
5JC0reitDlA+7wa0uTKo/CjCR9i6ziFeCuHhS3f038hQ5KYQdp6Y6ETY1MubH5vG
xeH9gjo/oR7qlBjQYi3Xq/wjBlN/ip0s5z7id0XuOvTVERgqEnqy/XnC/D5izthW
akWvfAtsDcmNteuvBrHSBTBAbSOBzlJsnab9Jkmrqzh+3BH/EVE8HnMWhtIXP6RB
HXTzXuvQTC65UvDeftdRIf+CK+DdfttTduWNYkyk3M7Yqx+V0/ricS2hIfHvmsd4
x1VgpSG7CK6w6b0KG2/0bAi5mSpu+25N8RYyAtJ1NfnpZtxNi7288zsn/CCavXWI
Oa7151vh09UlvKawFT5FORbX4ZOtCla5dcTwbhDrMeizITY4dLsvH6HneE+MA0Pl
yzFoD8pfvWku27hC0zszZAwPJzEbnn6o0PM0obWcBWyHGGWYPRfsRtSaD9KpcmeM
LnyFCs35a2KiQb63Etx8hew9APAb3ZUpguNMO4iGpXAKXGcJlmCr3dz1c7VtNkI6
G8rJP5LsDnd1PESTtMNT/cyOukBPmddT09EfHliDNXSLORXeWRDQVeoHlliOAL4u
a5DwWJmjG5cLXrphpy0XDkSSQlV3mfEsj0ZlM/T5GHVvCYVkgOtaYP4eC9ZYof/9
Pg8vtcDkFKhr4la0+8NGDML4/iJ8m/tD+b7gCFcCc+VaGDIH7nZatTLJSq8SIjUp
FwWd/jBy5xt28b4uIVhX+ycs+IVibGBoevhUC/5EtXpHfyfm0QIrTcP6t5M+z3H2
C2y/buEOL1kgEQ74dVaA14cv0kYrt8M69vM+EXagOEzS4GmszxMmyLGJttd+bV0l
AIyhoFaajoUIHE1Dz3rPzqqEI4k9uTV6FRZOKwqd/4HGZRqxlYq7o8UxreTT3r8U
m7jZT96aaafGdLyfVNIDxwhWp2GsTaKVtKeoej/QdRG9XhTcmoreYxfTrE4EHB3x
RNXPxYVYn8Bon+0rYd2UxjdbHCE3ejIK2Fl5ZtT0j8FZM8f9TjoYQnxWZkNbBg5e
Aj1Ke/q49/US+ivaAPwZbZYAqj90Y3xafioV+EurRby8ipPoOGN+ouvMw1VXBrat
mqW+/rVOed4B0FfB4jy21E8x6/+09BLzn21LetcHLgqXA7mRz4tOVlbSlM+mKHEZ
I6/sCDuMhKhX5zJdWCV0ESDGKoNFWRzSIGDkkKVFQRq1rptX8JX9oi2b93hu46Up
CrZamzmO2H6fpSxGvvjeTjC+BmUfTqXaMCX+IDigBUP0q+8jFOzo9Qw2c31PENbX
fP57OvV70ygOyJyO0rCVdPni6dX6N6KhUjvWOe/LuxqI1dW1347B6cgqg6itueUr
qJACvvpzi4sFb6vGfUB2WGNu1trYOpxeVaDpnBmkTKMQ/QI+1P47jlM86QBIUJ2X
xSEeypHSeDuVk+u7YqBd3l0SkH2ZsVjNuKcRvnToGz7+Kw+DL/e4IrIHbxhkjy4g
134nQ0OW6tvigbwaiITtTUMTJLetKl+hL6XiE0tHHz+ALHi1xedXUcUv5Zc1tFAJ
jXSCmPG06lSc8pIiU68lVLZy+8RRPOUnGUF/B8IFduu/9iIGIgsKQNJ6lRtih1lu
AMmXq62tJBMDJ/CLldXUbe6thK3vDz0ecS81XqN1poScVH8/P1TTW0W4SRSCkKOW
nuosO4mUjF5H2y731PSN2Om0RByQdoD/mr5UqC/RPx6gngaCEYsJs38fqV0V6T9I
3fXm/a9vRIIxuYXNpwTGbA0ozCvHgbqhZCrqN4s7NAoPjekH5gPp/2yqXxs9y2NZ
FAY26TRBJbowvn7y8WTSAywV9laJCP/Pqby5dHXTvPQzfLh9/EFmhLx3CAsXjlEY
eg4yv9a5JsLybd7d1L+zSaxcwM6qV1V+t8DJneWG8cytqRSsurBpB+ErC6vp9bPW
cMeAfti0iAqa0ENNQYhpfqqN45N/y8u8kM3ydPjug6Pg9UnP/8wc/Rp3IJf9DzjL
zHSoycav0Ip3Ky9v3jHVqn/2Kz1j1aNVj0dMr0xhB90JkJFYwFijP1AmsLnvNql6
skH2wCYMU8hKxP4gdhdsj8dkN6vvLGVaMDXyEvoH68dwvjuEauNBDpEK66MyojMk
59UUNEMdj2B7M6zLtmqF3119R0KJ+kUCusS5VZyZje5/1T2x0vR2uRnRuvbSMH9/
foVdcYC2HZJy8iFTOszl/SEVrqPw/rNy0/pS3T4wHDkrX/N6b0VSzJGIfayI98Fu
5aI37GoQz7AXxKOlZQTBfpDSF2LWPlvzbzEI/rOFwqlQbDGDWYPZ3Wy2m+UwyAvg
5OTukRqoZCuHlm2YvjefpkfTUqBzBpBjYy6hQs9uQbogYi5XENlhdYmxl/doOSYA
c9ZSjxp6RJgVFZlNl4XNrztmwzIl0tn3ldSr1ZxGIJiX5eFLw76L1oTTqmpVCGCt
SORbkUoc97M2QorqUZfSfzT1JHfr4gfxyfUqhut8z2xjcTFs2Wjrt5MBpjHsemDA
xQVYXbncNOOFhXVC+h0Hks2VgZdUlubQnXzLC2zSM+x5Ft2TiJpNFCPOl2U2jzhY
yDJm0/Bkdf5jTGzPAyvXOkCRM4eP2su6ddQvEyLnn4LDQk7INUJiItlGQT8fAogD
75aJC0VbM+yVDh3dA3dES/XPeCDHhPogXIUyBtDhH9/iGg3EE9TKDDp6HG+kd+1K
wXynOlpnkNzMixPGqtgFfRt0GzHUTIBmfiaFobYyVJU0e/ecgV+kjNQ3eHGl0n3y
HTNSPseGDB9loYq5RkhRFHm5nhVUDCRVC5yNRBYuDYV5xE51W0m3bFUexGoAb3z2
CWPOKUjwSrS00rE5d2Rjrq2ZrQGDB5ZMlb5tdJtn1VzzYT/14aouyfyVdQvv+zva
TC9Zt5+TLPy0B0O/o1dcPfvqr0Y+EjjbYgxqDZrs0lQIzOaNGxBjWZMuaHx4o/EA
UyKDVElKBK00FJ+LqH58ylhghNbAacQLpn6EHPr9XBwP8nKvSmxGbv+LMwLbRtC5
nM9GGaCnvzXNUXB5kT/uM3KMkzkqM/002N05hrCcruB6okahuQ81HjU4lMR7LkB1
FyT9Od5bH3AEhcPopAKeJ2zWmLnj0k57LQpAPN+SoY6B7hneTnd0hvGR7yWtNg3i
8ZBRatEJ3q6R5525WyTqmaQ9oDXW2O2cj1y5xb6bkWM6OgRaSFuHdHZiP+tLT8at
clX5QS38KsIuavtB/LXIyNhGBgVbZgFw50sAVFBA76dgCtGsH5Zfe8f1vCw7OqUo
u5+lvI5CFVF7HophbpfVzkr5tJt9/NQKTtszHQ2L5sH4XUqqTTe0LOQm9FAlu5C7
tQQqhKLNEHMKbDdOL7rQd5S8HO7NcDSAqsuhLoBpgnGv0LTtNVXxzR0N4aZToBOE
2mIUP94M8MZV/RN3YM6/yi8FaiCGg5yI+OChG+S6PBdoRFRYjqKjJ3uQ0UrFMkfJ
NYuh03csFcR/X8GXYSxzHZGMQZ3jhEhu6ErFcp24zrtqVNgLgnjHoHqLtqXG1Ldo
eNOEE6EyLtVvguDB8n+Y3X/E65fKBcinv2UV20Kef6EC0cgi/qxdL3g74PUErTlT
9nGkRZKlPLz5/l+1GMsXOGT6oKnsbOJOfrizVHWJX/SvGnAVPuSZ4DZsz7D5faRQ
71T+rUTvBXsYp6TbDLocK/kzgT1bRWTsfw6vvL0jFgrf3HtfSyg9r0UC0FchpY4h
9eKb2JupMXYFmeOhL2FvsxXDS34ID8Uc5HX4sBXhstbuXOHOxOre51q+IgNcjpqA
ZHj3zK77RZMoxCXWMIFUhhd3IINHAwKIw4ehW8SleCEbGs8363+XGcndB6V3Vcsm
nggc1FA6tYSqENKigFJYA8nupDLARNf7/eiKYgKzdgT/KSa2EvIf8STgBn+8DtF+
L7QQBhh6/HwjlUE2dXuXhzDLNbErmX4/6E0RSYsd+IGAIWifvUpwLiPsavFa2REZ
`pragma protect end_protected
