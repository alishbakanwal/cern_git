// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:05:39 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Ta9kFiU76on60fiL3K1XeE46NqrwqB1q/Ov81yHauRYsT/P/xrNSTrHQ26VuX347
wE9CDRn/dMb0vt4ZDSRHUshjtP0IXI+aYA2mpJ/OvJ6y3UsJK9n4sQILk3g4F6AP
8cgYb77fBRk6yJq5ouD99AzMLgrtHSeSLr360mqcZds=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11552)
6LsaLdTpZqw4C+o4KVq9tGf8BBq3JN5KIv/hakTl0tPIEN38Mm4Hhy5IzAYOPrMe
nR2UMsbWwe6ByAL+Sqte3PRRUZSr/uGpbIcf2Nz9FGGqzXuEFEwWI247tw0BvqDf
E4ZJHFt4gjSkbZZfInapH5gSrIG97/8CoHBNsj45FzMRpO8X+WpSDVl4pc2OBie7
r2KfIi6xYaHHrnr/nnKk46wtCmgCwJTuU+JXkzv13LEkfqE9oqBkePylnbTfTZ1b
e41ZJLJbQg5RfRQbAc35ocGJT2cbUSHPe8RnJjK9eBrQxbXXsGglFYx4sVi+yfWV
9iBTCSkoLN0kbYEGet/hCnozw5kY9h+67iuGWzV4oOhR/SU51oDNdO0JPMo8Yydv
ffSezpGwnRdJkBfqDMAs0H0QnJdx27531qQzM0GGospPwMpOVq80hKvbT6QaZdVh
buiHpsvb6BF+rmtGI468Bq64fBk8rNpEbRUtZxbrsTrd+gdgueSS6SuNSn9smR/3
qVHllIM0AWztaK6BZb7ZE2gfGQg6fv9Zkpina1wsj7h/CRziycwMqPUELH+Em/d2
2JkR9gQ44BF1sspPF+VHHOl9fWXtJalxPvSGU88X8p1YK+vVgtAUBkNpPW9rTAJx
IRmuBZM5I2WMC67fcYUYibDg1uvg/NvxN1ciesPJSxoRzxNPfhuqu97SHXZF6K8D
q47dYSFoSDiZHxOHYaCSGgzV/Akw9PgugzfcMS7Rz1/7pNbmo0IuVB3+i5oh2+xZ
BGacwDlObX3cYjpcOPpXMVeat/M+7zshVC8bi/NUqExPsupLVRgUiGRNDNfri0+N
uHe1/bv17+vnXmKN8v35alWXZ1yAYYcBTJ8VpqmnAA779Ex8YyFHM7slnvtr9FFL
S9AxOtZFNHZyTLvIq3Zwsh0WoLc8Ut3mXptaE15oG//3Vjk3WyU05Ljq7PWIBEMU
KMY0iO5TbGNgNPH/h3yC+eIO7P1i6V0u6FmaTdUnNCxojjzuTFBDjFy112nYRUQF
uW5ANwlM2kfNPzsl9Jsg3Ud6rMIEhI/oc2rbr15ZeoLzaDSn7iDn91rRkX/kCyN5
+sW5OKOC1aPwvC/TAQwP+RkT1zUWaeOn1lDt+OQjwK5KVyiGiJ0M+mZotIm3zHHH
bO/5gNxtyI55wQeGKE4qIiM8BtlHenveQ+qW4vvd2zY5AQHqF2zcKP/UVti/HimC
03gfhD1bMOlF3JFg5eTTsJZR7JHLWv1Fsc3IkiY1650bkiYFKi4FWDJL27B7PyUY
l7tYGI8PsWg2VhOze9e95b4xxjzZApIrm0mTkU9knsEbFvuAuh9y0gd9EhTqYdRR
med4WXQ+P/U0BeVP3b3wNoqIZf6j8nFw4NFRAD1rAJcRGlhHmwE1ZcmDogk0TViv
j9zUz7WJ+epEy/V3zIXOVjAVwXK5Yd71g6f/MYGsA6x/5Zt6rMlrc6YwKwLzvuWf
9Atw+AKM0Zzr850DHFxgQxBZ8HbOBmvcN6t/jzw3QbEKrNks287dcmift7XgW9pv
TZe4PAgwShtm/CySv54fVsviZsoOgRLiojwWR5Sb4AOah7aNVXZDEp4J05OtRPc5
Nu15bVwLOBl56EkBo/nQyx0UVk2oXtup+zQ3O57J66JQoJPpAvibMQmdZ8Ku98pN
N7BwpMEa8CtHHmPm/II50Iq9SbNboETh4BpAOsXwB/LuKMxDumgqxa8s7po5Y6n+
2S34XkJzoY08ntGDWoWM+Wm3Ao/Cx2kEbjOW4Ml4d7IuT1CEQseOoTw/bWX8bRcf
pkazxfWctmuvN4Z0dtZnDgJoYN/sN9RfLJ5tmM6gC8Q+cQV+mOye70/tb3dMvk2J
svGwe+hXq+otHZVs8VoASU662NpZ9CkFMJJbHBFBJxBRI4yi5UBG6sRqOQ1qA1lw
CMRSbRTfz0cWr+vKaUBIVN8+qNLMvbg0VZoM5rawRJZY5v2f5LMMfj/0HPCqCnLA
yvYMWi/dlK4Rh7WpddR+Og+4F0ROz9QCmPU7Nmb2lFrm7pELYsnm6lpHORTJANPA
SskcqTPGnMybYjCaIg53oDyfFzWOi2lmjkpMY5BJQnmX/ds6isjK7QBOxqv6DTfz
uBJe18YlHirXd3dATMk+T4wcqBNcFlufTmM1YFnBxPOx91lTGWJClrtZikgyfykd
S/IFQpzKsdOk1jTk3Krf2syfCFeRPOBD2ElGoB8CK2hd0qXRXu+E5OOSsS5TT8Cd
Zha0u3mWqE3VClcx9N+pAEjm/wybPjNLQrpav7h70ay/XZGxHDVYnjbmLnxfg4wX
rVRxPPTEgK1zPgsB+7ipXtC8HwogPNatb/ajXzTvWVsqpxdwKZPCj88s14C21TqQ
LcllPMFoA2ZhQhGIomx0261dzCiOlWgOB7SM3/H7rnGtlrzgcr9Rge2Do4M+3Hu/
iA0OGYzFybhUybRqjgvQ5msWOtZsB9Vj9a9Kv9+9WC17w+fyvYwdmzNYxs5Hb8T+
O6ydf2atUrrNDB8O7Sf0jvmbx2gdInX3mp/p1ewDHYf7gRDPO8hDdL8/1SjEKfW5
d3G8RsLFv+Bx3gYsCUT3h0f7r8FUjSe8e/6vPvRoR+zLe1XZm+kvmroIPkayX+63
/y7lD4s3NiVspHqTEqRVmofDrM4Kz+D7TlH6zec5GIfS77zZvpSsca2fWA2LlskU
sZuVMjWGimSTuozPefFRQ8R2F0gsml88AuYdB+c24jwF6IXbETYpbnzvhlIvxnXg
3Mp/pqxbErnWKESXVZZKqDPs4Zqaajqypn2/lxvzieTB6qLIosrhToVmXA2u54mR
+2KKd/npF14y/sWJd14o72UYgHiJZtvFqEDtrC7ogemo7vYfMjt7ASZ/57iIe4CF
HjV97IFPmncXrAjruN2rir0ejXbPeZur0QM5OrlK0UOZxmKOTvU0ABHHpkvi0/te
ekzM6/AAWmInBgdcPNEEUE6pF/vF5U7N+5q84ijQcVYzzgZ8ae3ygxLYmVxXJIVl
OxtoMc4YCuc2qc3Ckko2IxwSc3UcxcupoxFId0V4+qncbvJzFBZJh1945Y1Dhwcb
4AXecz8JODeab8L7lsdw0hNURUEFgOjmpEVHTmXmUH/RaoiDocCtUfkXmzFcVSE9
HGLQCRDaQfmc7XIhw14EA2c8cxzV8Hz1h04tGWEaaFPmaDYYxZqUQDXlQivPNcLa
k8bzbtMIw9a7Xm+8MRqyaMAIo1ayt0/LEoAUOiA28isL1uTxMSk6FucCVDLjleAD
nLyy/bMjnbD44NgV7fMIWz1/hlSyVpCUrbMt4TfbDNmKuqOCYoPRGy1sj0y2lJJ/
aTby7VZ9m4TfgVvbHrMgkJfgw1Ucae58/N5MxJBd/Eggy94lH9iXUmdhhzLSorC+
KiG6/BtP5KWckslTwc3u0Iv4zzCMm2VGK0sVOzwxttWxc53+RTEB7K24EOGawUAI
8nfcVfqbvcZgYOXSx1pk2dXq/EY2kp1IkWmjdlLXNoYNkmqLSSpfPFElSYJLdOrA
tuea3aoxY5gWJw7UmHsJJvJ81ML9UrkBfI5X6uNWdX15k9mfV0olhkQSnlbFoM5Z
lUsyeayIeWkOv/ha+vaFZ/nqZLljbr8bLAbAq30+vBfqd6AEjemUTqPimXkPMrgv
napS0hvTrRlmsW6PpAUFZg5uZxSbi2/HgHVyqiKQpiNnc4gXOpH2Ald1jCAIzHI1
Tnb3HvV93GD04J1ShEYHeZox+VnskJetfYWakcrJhpTORO5zzaOJ+jerMmPpe04s
tTIuIfxy8ldRsRSTZpM08k6ifEvDsKPp5VlSojrJkbMJ4cY8C9cJ75OYW1KXtGyg
fONMiS81wTunOmEr9Qee9GZvac0w7DcMgubWcTqGJ4VjUpUJqYHsnaqBYbhjSwq6
rnuTWEn9mlulR1yfhBj/9hIiO+a/sv5OYwuEo7cAixPt6Q9lWWXJA1Mlv/y8NrMt
ZL6TJZwRccUtQM7YisCSOjrkVmkanNhfY0EpfPFnN9Glzn+qeRqmNaG9Pa7zR+Xc
nbWr34A7UmNpy9ORxIA7YPQCadJ8ze5QqwkG6XVv8HhQDMIsrRHbWGwhBXoCGwdV
qFRm0qmK2hk8jhvYk8MxMo35If3/E92NoTyIpzewps5+6h6cy31bMERwMalKO8Co
ib3PtAAjxNAIh9eYfe5EPaz3pwi+BjSZsAaucxCPqjRf3fvvZOihZX8YIVskp847
Wvo+uJ/2Q6ySxTcDZqLgWsxekP5qsybsUUBgNw++Yyb5RLnQYXkMzJhUTfwZ83OL
VDc4qJV+Q7KC/5aulJgTBQFKY/Np4qNbjhIwtJN61+dcfWfGZY7XksLU05IQ86vM
7NY2qym5pNA54+3DWmg63h5W+WV+a+yCW/5jdSXk1unGejN03aDFhAThPEWOCAWm
8elHNJDbXnQ7XsVGy1HNzeDyDOQBHvY2ngKn3zIJsMkSs2vWXMS4xRfHV/lxaRTs
vh+B1rSmsT+U7Zth+YmAdxeahN+txg3hi76Kb4Ni8DLm1wIiaomOx2mgr5lWO++L
V/vSIaqhUWfTqMGdBS4rfZ4+HbEDK1eING8XTfLbUSdKNZKV4fecZpudmfaFQyvm
EwKeEqlR76aci01YNYs8zIthYqvSz9qQ1XZE6tXgw9qw/jSUiu+84DTpMFtppfRn
fm9N+gqUKv2tcudD9Qr9mtMtc0lUO/3sSDYChEeILaIr/p6z+SE5ux2POe5A5ALu
R9bp0BYwXcKDFTzoJw0dYH/QHOuW+71qzVcBHC3o9HpqMUbsOOr841vLSc2gPPjb
yufICcMaHk93On5dMOqiBgrThEOTpmlizZm13CRCkO3bPBBeE+J/FweN17/bwhH8
39AhGkmUkH/yPVftTzxdN0eWxvMUYZSpbcPHVAVSlfxWS0mho7mO64BIMxiUN1lq
FFBWD767vpcmntnycjA9wdIdAxV8kZPz8x6iKt/rhz8UHntbjVGhocjZtCNuP+K5
kG0sj0+0VbCORIZcoio0b/BZBz7+TTeyh4dZ5hT1ZlpFOcutMTSPIC1+SJ7iKttE
EQKbWPy6EyC3t0nzJYDH3zWcE3LjZz8ml278coLtpYgMsyBOaghh+e5r4ZobUtRQ
EI1s52d5SEvKBsXBVD23mCAlKrgXN3aE6cq7yOCCouyohGeUtp73wKkSKGqN+nKg
Uisgu/udYRE5AhtZypdqlBuIxgzGQT68TpVM8vGaDrhbJL6WIVyIFzkl+dthigKl
3spsTmWi1PTDKMlFEwBj5YPryngu4wnJDmMoGORsu5gvFIYXXi20i5X328QFQHTD
6Porcipjd9bielHjIvqzlSdU71kYXXmZUBXWvEp2uby+ulGNEx7qZA0FqQSPdHbM
9p03I5dVlPtgE6RQWpb/67Yb+ygSFTOfqDXgqRJTZ8vr/BB9L+YLcILkvrZWrGTZ
NdjTQsh/ml5CdrU96HXvoT7CVBsyiFLGYrEbWdNdnXT6iDe9gXIL7rsZF40Rprst
OG+Mdl/q9TRT2/xMnUHZ72Qhm/61tpqg5Cp/eofqBZqiyM416fhnG2obhxhKnV8g
05okoUabn7sQCtK4C+ZEWXQ3MTQlcVsAsD0vH/zMKDSncJFAwm9rYqTnR8L7gfxV
DjMwIE60FBNFGQVr1fbLUwd7wAyYypP6RLtX7UIPP/uDkjLlUbDuK7qx+QP/6Odc
Bfm9qAJMacY1ViyxgNVFMaDrYBp+Nwcg2mjSDZL0/Z+mInDIXaE9ZsSzvllba8c0
/tOrkVGXwds57REg+j4JfLAs+9DAIF82oNHZ9TaDjOaE2AKj4zzruwASigmDO85q
ldDZDowE0WKVFNoNRA6rFeUfUy0nZK8UdGEfrFAn3MGbVtsN3pFTptO1rPHZOADD
AEJoxn7p7mTW/npNWPAHzZcSsVnZeVihYVwurGVAQycKD3G2nappRiaWNlo6yhgY
U6S6friJjkl7t+Vw3/pLJP7wONfEe71rOuNqf5NqiZlkLAfvsssEZTfLayr+Qddr
OX/ik5TsvXVDwskHjnpZ69De2wzNpsK+0vdx81dtDk+6WJgjB5MqK9iVjLe4XQud
VV0WUzYJKGv3KOsh8MD1+AVvP7vDQISX/W+Qj2csgF7KVKYFAR5cy4nDXfP4V1G9
DeNA0d9eA/MNwBMCyHDqvBY2/ZLOh+u8CWQOCSncrtAKqKbA24C+7rYhm8kagl+4
ibzjd30yIKZ3Puz0ygWgqy1HETPOnLREs0wvdLDjuC4J2TkUoNB+YbrrIMvGu7Nl
+O8cm8ZrrUBIolvx1Ruvy9zfdvjm50qEGdufZW5tgy4qu7sVYxyDqJk7QNBMrxyx
UO6hFBDSCI98H3VDS5BkGboiCNHXQbAhJBkzX7VsW8MlnFTTFrctx5jkUr1vo10F
WeqXMqlO4a1hwhth1qckceFZvHEMyLl3laq5wGuGDPFS/wuKFA1TRzAr7p+Wb5f/
e0FZ5VUf0qoJ/NYXQ+VjEc3wV9xlm85MN+1GsNtvBcVGZduVPJe4cykvKdIK0Xdd
NOCRQOWKJAb/iWP6cS+ZLMKEBJHrjEeKYTG8lxUrxDGAnn2H/nmbqkuu/9fzbU9H
fmU3drhGbSmQKTCzPmC6TZMus9DfLc6i1D/kAwq9ZRuXxXzj9Ht+xDIq91zxY1IR
HDjJLBsPwIk6ZfVgN8+D93oCKi9Nsnjan3525FMAy90VbMZPpQbmEA1qVXzadPJN
wXiVPfQal183u8xlstD2DSC1S3bcqNmO1dFRxDPWlY11u6tsHOQNJXgLAM0NGzQE
29zvQqeDtQUOKlear+Ay1mhg+pYvKeF6nJXemFhtI37xMdyHMK5lPLYD+cufvgw+
RUmzxr8neKfWrJFwbAgmDdJXG5g5pl16qC3vd4MdS4WWXVV1Z6LblVLqbWmC/wP2
Ofdylx8jhph0UCZzfxLZ0ahhAtZiUe+lF04WbPOSIhRo3vT7FEUun/8NN4stgl0L
dQcXZRA9jvHQSJQNjjCLf2CnsZKF9rH1/vapZ04uHEQ9Crmr//C7sk/zSXGbon0n
M+eDUx90XzMrrEhRSsbCUiOqF1q0/ZTeT/QncToF8svPssP9LAEBmedqS1LXme8J
+PpSqW0RJb4JJEg5m+0bN9rNRdg3AAio7U7s6uO70+cMFXdPhCkjkdZKNn8TQzSr
tG3ltThZHMObHcPb0uOH+CL7JJkcorSLWTRTm3OW2OCNogsFs4D70RJwhWyZTbwk
SP6HvAzo3ON3LnNV/n6hcDLm4tiHFnYu4bWNIcGAPqGfytP37xbIPtPPQXfaDGHB
uHxMEYZlCNagr+Eq3b3j12Rykq604Q6M1RDzmHMyO3nyIrso4KKeAAu6miTwCX6K
1otklzKFonztYUPvtAho9xUw1nrTDaRBU+c86KgUTSYKfyMDOVpekWySnIrtTNLE
qIzpbnDKb6OItjHLFIafPA0vUFYWLTdFNDYqDqPEz8rK5UmjjnM16vV7/8oOvTwy
vRskvplfufFXPxnQWstignjjMcS+yT3bS5sgRIf2IeU0D4hMiFh8ezkVUYRkird7
m2j+coXorKs1jCm6BIUxlFRoidJe6tJgb492cWqXZgEO3qPcovmZQVvIEePyv+0v
2vXjf1kdD1PsUDviTcO/tAegs6TBrA/rq7GKo65pS7aliu1BQwoH9xnKxQtcUUdh
I/8HNkdy7pdewLmzOdeRbF+zzQ7rDnOOAoBRlqQ/95C7ADPVzpYAKgJlYGgoKFNM
7zU4BKwghWv6ASBoG6ZvZNNe7l8T1qjWi1CNrF4yio1t5gtEzwp678tOIbzoMlu7
2qvDiL2ED2K+EUsIDtxkog4u6AICNDNeTn3qGFhnhEXX0OGnhsQJEZyOC1mmN7Ya
4VKvsCZXL3yEuPQrDk6bjyRLgnc8EiOepaMYPkjLwUJjTXG55xWma4x9eCr0VaFF
88PXIL/9B8bwLn1/F9ypcuUD1mqB0K36v4uvXd9Jhb3QVyRtxp9IAMlBhy73ydSo
SKkM+M2UOfFD3Au5ike1Wu/hg3gt4gwe6VABp9nurTQLLrnfe4w61DP+mTYPIft6
auKHF7U5gQ3jpaA5kvbt0erFcULYsBFcsWugSkm/gN5Ib1EtAt4lz6ovxN43O3/r
WHSry25OIK/VqyIvlqEtW0TZQ0RVklHN9NVU2A/iLYg+3t5w0s24oTEC+612UTdy
oE41UrwBsVSbUYiF9yMWkdr98Fz+xbUUMvbuZp0AAM0HRvGzdjSJ9lirjBr8FxNh
mTRwx2kmTUqFcE/bZ90MRCo008EKUnnxXq8LyTCFiQ+f4ErDPVsiACPT1I5+DCSv
nwl1iMeppLC04v4Nd28aroN0R7a5UosdRJbcG88KoZvulfa5JLRsBvt2mfFSWomw
5+xRHKn5j7pVTxt+RseWaWGDf9/AmATHZGkQfb1Hs/IfShvYQ+DR+IDyMJt2kLbw
G5OtWGfLymkvbQ9PRXugvFFG96QEFWvC0GX0Rc8r70PhakQBfZt2ZijveIBRVVCf
hqqHDvHu8XmkmocsTZvv0IkffZQWPmI/GDu/MmikkS0ITpccmlTysf714Ju55lH2
OofX2USLbTen13vu1KJ/yTeGklc1sFpjdGxCewM1XWZzS+did0Se+9gdjoCf0mja
PfiMGdPh37C0mEaPEh58rS270ufotjFdU14Bvx4R/n04Bfckw4+u49L74F6kgblA
+YEt1mRoOf2n2QhL85Q5rX45B+sZhV6uZREf3ykbWXXOKv8G1DQhsSkfa8SyPcWt
BxxfZDhueGtOGKFNyG7gzViBwKrnDgs/Ev8onwZJ2YvbFlJWWLAEF2iin6psbd0U
RKH2/aNJEhnu8xpZgsZZC2VZwrvmZH+1iDZXhnpoG2/oSp4hvIxB/iu1FPcAB3E2
btjon4njUUfKvPyoHKwmLN63RK4vmKCAE3fPo3jiqiQe40BdyqYGpFgSNZQBeZpH
pJHAaucxRZKhKhhf2Y3M2Z2i3ekKGXsl2qm1Gyn01YBOpMeZC0EkKZ+w5HT9jPAB
vy1WlA3ky6JS9LDrzp2WYZziZZA+z4n0fKPxxZFULPhK19yAAi8KWCcNEISppc4K
n4fZZ/aNXoaVvyocfssMWO2iIW8U1RvT+L1kDDjVoY8136PHXKKLbGvuTcR9WV3H
s/5NLwXHuacpnZytUcMviQJsTF44LrHKcgKhbB1CnPh4kSNR20SLFHvuvRxKUM0A
Q+6WVEZaFCJxb/eUp/RSbEXok001q921/md267iXQcQbS2Ajjs40sUYPZgIfDSdg
jlS5p/LfKe47o+mvJgKi0cqrv50Zd5OkQn2QSnciq6p+29xp2jTs2TwgNL7W6G+M
tHDBNwSnb/xXHtMrtxWNXLba8gr69N4yxy6ZQdx5u8CEHtyxr+B91QN9NxJ9AR9R
5MRu+zCP+YoWyXz+Uvz9yZ6Ft/Y9p/9vMwzwKOmrLOs725a+Aw+cAUodEr9p+5+9
SZowlpCcRk9J0qkIQZrbRepTn5s58HrNncjN0+MCnu/22MxjsgVOkFw6YldGs1mD
duBH7tBsU4+gXBk+gqeuQ+fU9cN/RiBPSqChQOLNylev+Mm8z0iFoF0dCrz2ZFgq
mpqu2XyS5KE+Wx38BuNODAHDjQNwFLWRpfQgUVnxlPeJShTXTFPngCt0+hsW+Dny
J+bRYRlx6WkvWLv/xR/XseEd0tVH8/L2WsluvgBVcYVyDSA3KKIt5CWrpSNcvIGL
80FWe9vufxewGN43uARMvxNvx4RJTVF8DYjLdTHxgbSXLEscFeAuNgJiNddmRlCv
6UJefhrYTJmLH0NRvhP4uWncyR3ZcvN0wwJEhB6l6y3GTsGzthsbQ+kDTjTwmNvx
Ul4ltKULwDMD3jMm5IHcMBNAXD6q9Cc0V6NY/h8jv11nPKv2LHokYCjcCflYwZvT
SzHf9TlxnKe+lH1cVwqtjUWNn2BnkiPnOChVz5/ajdTW11axkz3lv07SMM4y7O1L
DB3wB2FxMJ4qa+MbBhi5J9eg4LCqqReJvUKt3IADrlzO3tm5WcSUSI2HLfFOn/99
XT1ozxGE/2MAPbN/c+AE1JLld4zC9DGcYsBd5VYz+Nay34FOv7cbn82VM56SQSOB
4qR+T+g2/NZ4pBvY8VDPmApDxxqw2JiGRlgJ120JAhrZakV3ciHgirQIDvHTMZWE
fM15B4dgfxYSX7q+jzz6mlilk50RS9WYzfPplTMDyW2nvFGOqcYbOwtz6zjvpY+q
AEL3KeS3QKFE6LXs0ipHmCmApQTsLOCApx/zLe2oh0c/nOM2q/EMqXaJlYAtOk7t
4Wde/sCvuzonjOhMC1w6gS8grh4nvXbve+EpRjCCD7xG0W3gg+vz+RwQMdhSThFM
zHjwWhtNhl7EG4+z4NGwlzs64COzLXJ0SY16Yn7j031EZDGZaQ4zIAqyKUWjM6I4
opJwImJwBQyiaVkvDBeYzy1put7mP+iQ76HcXMMXwf/V90Zq4dlXm564/y5MJxQE
83BhVBxvXm7yTS+B1O1I05Pt0ECrsOr9NgD2BAmawf1bEIK2yhnkTR/RKo8Pjh8o
N2I26w3LGCjlDPUc7j9cj6mXZAShgTX2qf1d0KeUg1ZQ50gokK7iGo8fGCH0m8hW
f2RFPGYZfKMGwmi/9BPLubOxJR4GVOwKg31AHWhRcyi95uRkl77cg5+8EUaLa76k
JkXRY2MDyL8Ed7vWvO2UQVvfXvBhg/D0SXoeHN29HAGC1ERAg+i1GEvdbz1TFXZc
mjOFB5Bubiw54fLKrCp8t4aq/pim3ymZfD4+GzToQCHo9mj8pMjoQc1WnhKA1bbU
K5bAW3V712Ttdgqxhd4Vi60hyVlkADgIv6m3lMAEyZ6ojQRnK8tHlcBajY+U9SeR
59xOfVkRWRqfEJCXiDqOqqMLVlsmireYK2Ox8gp9JtVB6qzmAQPPxaugotKG5/Fu
ZkVo2YHDmucBxTBrJUX1I0Jh+cRXWCP96v43wR0uIYX731TwSrM/326WNEEA3niz
UxnehsAdu3OvlRR6vyIxw+a0OQsVJF1ynAH3nrbr2GlNvW78okFpXEFcZKjfFUZo
Niw4lHy6GDVfVN7pWyaxpru0UAhPExNgDLfVtIKR/ZKjmv1BJCGO6kClriHm9Abn
qmNf/GMDU2y5CLN6TlmCYGuT3kUcuKMsjSl2EuM6a8H2kVRD8paWjzOR2gVJUytF
unIc6e5rHxHKF0trMTMmhhT8w5ccTd9XRwbde/zNZZ7Ia31vdbhoejBky8pCd3Oc
NJWk3ExeLxE/JVipUCiJ+4UfPhCIwU7VvC2oLfD5Vb0tDMvveDiur1umqBU8Lxwb
P8LLpd1EMC7RqMEzIvap4dvtqnp4og2Yf8sid5wB4SUhjVhxzbUto6wa58KL4phR
+BqaVHJ869fXNeFQF8BnA5kyDsyhauwAfyIun3V9M4FgzLzJvwLnM4YK0OK2yRc/
uejcRsbJzMEyHmivs8rikmeGnfuEFU/k2LTJi2CrLBlfyw5ag+y4ILNzdThCkpBl
/rU/WR+DqZjZYTqx7SlRgauOcxrDpPdZzSICV3PCZJaELnQU07xhkze2CkbMqOV3
Rmr+dvtk0bmayuH3pTcfFJW3/q6eidhlhpmKLNm2B/C/ZO18ouFTyFci+VBrTt3d
TAdg94meodnP8Z/pz51b3VQJ2iOZ/3KjUSkZkergk/EsKbsWImMXdrExhfswKdbg
J8SBjd09VoBfCcryrZxym7MkP20kqvnG0qkasjF5Wn+ocrJ9aPsdKsOijB8zWFX+
6CLFZvB8D1Rp9IkVnNVa7J6nQqkqLsKkIFIQfndOCvUs2mFpGXaYszOfyGAF0pyE
Qa4brT1Q2ds7SXwlMD5nlBJ7qO3zfQbVL1NQgWVn2YeDBl+jWQvOcK+N4ax4n8JG
nt/vQLe1Ju9TnigkWIL6EGvH/c/uwSbBBl1RQ0QjWsd2RHOcbu4E93gFNo32JpnO
CTw18dItctMzxXtzhnPGVqDyrFC1puOuxs97BXFHNj82hRNLvvuxzk/PvwEGle0D
jEyXJv0QTpZulG+sUtaYyiYX4MRpsjcyOwv9ZMlCXYd8dw+PQob2kqw+XsjhgOpy
6DWEMQG5jxZbKziDw4Ti5TV6BP9uLIausG7rpClnvQqBeMqJ85q0CESVpIjYREF3
82xAd2P2L1wcVjdfFUk/4QMOcA1h2/lTcgYd1ViD7+mXWDzpSdXOcuwh323tJ6K4
JLM+A6kC0F8N9d3nVkQ9sddrgNuctzhw+kGricAUOiifwF7x5RJCbThAtYxWHp/J
rEyGY1zF201z7g/bIDml7LHUaxR5CFMy3Hdu2saVXUEgbyhwiIFei0AhKdRp9KD+
awnzslmFgnucGjmvenrrxsAFv/PeAQrZUMFrcSXWdikGCA+732bQghfiT3IwCpoy
j5kGiE+b5qn/fzmRFL3s2KS5iZiNSl4hUveQGOOPrPtsVtwXJgi2uL+HTjufrtWO
srpH9+TJKMLW6oHntbFwwUU7E/KkakZbmCMlVl+mP2r6+BaAOON042+r8OEXjsTj
qF/Q+O4mo3zdY7hhvC97NBG2Qvu0P3J/I9qNTaalx0x3VCHQepThtLd6qUV8TGdU
eSraeV+Ayh2+wrAIm7+/xZ1XQWmimSVUBvF9Mac2dnQdFR2tIdY44PsNGCTjDu0d
OpC6lLVqikvP4qcdyFLOXCRS/cv+bi9Z9nTQpDjeQ+yFclZ7qXIXZYUSHc6p2dL/
GbZ7M4ZP/FAMWuJG4/rkQjp2ce0OYO5yUTFCG8EoufaT1RDpQBU1Pt7sfnL2BvQb
C4568i96ri+95OCUqklKqO1qhw1kB99gmkcXkMrfYqsKvwhOufPTYQDkKVCTRdBK
/FyhYQi0Bt6WsxXgU7zTN6rBABY6ISgPvGKZs0kkwIOUW0tRi0hO0y/u7Tad53PY
jeQFN4ODKT6Z7WT+4TjOkMYg0bkaPN5rZEmjf2+0eA72btVYf0tpVtSb1WGuLgRg
fTcrX4Z1DsCKj66O/VEFyXtHW3tl2qKoa5Yj/Av6dEf+1u8mCG/3OJGMBf6SU25K
05JABKjPOOAu2CZXkBJwqJKuq/EZJGVoHj/F0XEbEIqz8ZPRMHQDxhmIw36I8gBh
fpFZ4DI+RWcHzex8EQqwA260kzDZbbX/IKi8azPa1fVOebHGVxZOPKe9WXaSyvsC
mpf0cd9lEQxNJsnT49uMmbrSFwJXoVLmLn3nXLjc3eRq+C8YfCAPX65xJVhcHSX3
N1d80+A6xyqF5EFVW+kRV0PrdEHFA62nUGBgJCurwZxBn70rHklw7V33sSQHw8Ms
Iip9+yWr4ttcBvNC4QczX68vvPctC/IJvLvc9uceqUMOHzlYPiP1bXf60YNFZUEX
iiNJoKol7Yi17IBqiSyIfkNjERb1xMDkhYMQftE8ekzKK5uPK1vle2gL+9XTqvVp
X4YPDP/pAYo32eyZJ/6PObP4PeXDsmII+W9i0p7jBLH6WE756Bdz287hIFyizy++
/+W771oxHME3CAhuWXTZaSbTtB1Ya1n22NsfIx8tdREka3hQWqn+AhE5TP3bxH6d
tyv/9BgOKXfdckCl+O8LKxbZe12MDTOk3BBkgzBCOsbJa2WBFewk04Elh884ropo
kcHvzK/kS8ypbiKyssDjPyjLtoQil3koOR15kJTiYkFYlZDECcjQENSryFff0Fa/
Gh52GaQu7I5VYW7j+prxtt4ZJQ5vyLIWJ7nIptf4nvkEH6b55P2boVm2o5KzpIBA
gUXjeXMC+orw4mAn4Y1jTGpsEHwViGANJiTuao4yJSjJVGG5+y0YDZ+ILEGhn+IF
UfDBiRIbipjcVSXZd20uuXqgt9iiHEf3RCW9pvaFr68dXKMHeCVJzigYALh5eVrO
NbYq/Q2U0ocMV+NtBBfWqZUZFQV9LN93qlvdYiPsE1kX0YeAHQLTVyaQhgCIGk6d
/vbf3cjwg1M8Ga7Nf61sbkT6y5a0Ybj4irF85QcMhNnNK36ycjOboyLHM1cx/AJX
LqJkeFa6wEifSZJhsfurht/ub/BiHRD5uSa3xO7FGufm+/XuDEXx/iQtJ7p7gdtx
eZ85fBt/+Zs08nsu/jXojgWT0k9MapT3svRGyFS58xuj787slVwgDLus7O+rmeyV
+q5c31tW9Y0DZfkhOXGUBuVVRrzehE+byQkl1JnDqI4xryratVTqMEmwuBAG8N5F
v6ZedLkcqruCc74iUBnCXOyHTxwo8b0yezlKJTZjxghhty9rzgOYpognjS9RoJDu
7Lalhl/sFIQORPePO5Hc9Q+ItWDFAhypX8fvAbM49vHl+eHDI8vjpKppjqCcgPvd
GQvwr+4gNQXfuo5VreP/TWoxHmZao7XLwLtD9XpueLPvr40CrYwuWs3ze4jpMKTa
4i3kAurzWmObL9ga8qo41+GrjQNYrqDrgD16MmzWjA6G+ijHpXp5cvxlfI+1cWoS
8HI2uylLOggNDeGDG57T/1ry5a8vAKY2HcbOP7UOFQF40G07cC59XtCtqs2eWlOa
4VkhC0+tE5x9efbD7UTCDjrO+L7xASV3LgJI9Oy2gpCB3veYcogqiM7o0P/eQHqp
/lXL3ycZmERlEUzWLzoQl78qmnGnzEve68JSBhxjIq/yxFS7D8D4cLEejkzaST3b
yYxhCXcUtrL7ddZecoAjqrJyRO5lqs4SzQffubSA6zoFrQ6kibFq+sgaSvgdhR7l
OO4ldtl4kBCUsu9s4Z/bd6z9EtNwDICuahUUzEzN0fQOJio76J6fzjNths05fZ29
h+jy3q94W/2DFfDuWkReCNQmf9B6hVHmbNb9TWDDGklZp9hC20w9f8bE5r1IJKsS
mRkFwO2rYdd9JeS8PLamxpEP03/rjGrKQN2g+ulcSE904PI+abfDzjeY7hQPt8yl
tntlvMkr8AS4hJXhWlEpT91yDYE8bOMX1gBv67Y+VpYoHZrgsrqA5sPZ4PjYX139
ot+wALtda8I2DJ/BhTVx1Mk5rrIMRU7KkRGYz5MtO7B5emMhLHGs6pDITHslBtu7
mDU4VOQhg19VLBXVKCQTX5nNXu6O3VFOTe8fQV6RQG3a0hCutBkplCOxayBwMdwT
grGDgxBnydagMpvtWuiNRLayTPDRyCWRRh4GD4LVfEliM2t4QGTdTBi0OU6B95BL
JAZAy7qh2QsvODJeqczbMRo11anYpyIm/4MW8EKEsvsMueH0EQppPl/CfWgtKpC+
9GucCi9ZW95R01Vx+zVEgdL5svv2nSKl+vu1EdDrwfGyn/Y9hneizCk6gCGeO7XF
izSm1QcretkzPzFcUrdGeJjDYlHs/pIPPdbZi+jfB1Tssz26eu2iYHq9Qf3KkdMZ
iJ60QhsfFvT9fA93xQyYxjC6OcgxRRduIW/sF4qcNSs=
`pragma protect end_protected
