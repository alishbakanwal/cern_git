// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:02:08 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
NtL0X8NNEsml+vqShtzV2hv7BhiTKgpbptpi32dgSiE+TI/LomlTUu9eg7MTVMzR
t19SUbEMDfddSCAnZcaizVk5omtXSOHSrtfxlSv64BHrrAWIBPWF1ofF3l8cKxwb
qn7/0+CPOgYZpl3lb59+pC6QbDUg8sv/TFB72ir70LM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 22384)
5hBm5x3vlzr7JSbN2glMnVKUyX/kvZXFla2BtCAhTMcZwCIJMMyNj+UixZnSwy1m
mp+AxHJqdpXRkCTtV2812+Lqc7/EGG069p3amTEb+dTPJK88FvN+woXaJj2muStr
RyER68r38iK/L6O167W23/xNpRFek9wUL7N9WfnRy8us9wULzBgzKEX3752WhSQ6
YpH0aLi9g8VBpD3dzEByS8TZ8ydLYgytXydnuyF3nQV9spTDYhsR90fezlyIDlQg
vFrJM09HBR0ZJziMZuUGUD+LrBdiDLffOOwfoSztZQtygofPcFX2FIj4cO2ruvfY
4J8if3WU8V6TBjPhdX4o/ody4Vc2IcPxWB0aGtXNmNjOdOE2uVVJj/KMBb0QaGAL
6FiHA1El2uQK55hSNTvvhx19FkXEij7Bpmsph4uFaxVatqtaZiIkXsoGx0kIrOlP
3U70mfoUNdQ2VjTB7gGWmVzZ88tBFHI56o8J12bqepVdUgB19w3QF1P997YUbhSH
c/EXvssn+sLrh4KRk/4e4rVheANe/n2W5qPSKns5WqpnwyT/A/4TFN/sj+j2/fn8
GKWLgKTwqS/EATNNI/YKK7IelL3I5NqKPzIGjNBEKX5FTRwylnGH976mAwj8cKlQ
k+EXLSXgQEbQnzOJXMJPO2bZffhgWSZLtmFQLG0WUOkVAmafFvmghgDah8vt/L7d
4teS2XYpPa+X5pgO9gGkW+SrSBPR351RdXTT3St64dysiUdFOV8Zo7XL0NcTk3kX
1Qfwp322Uu5bJPMoEb0vYNVbobkj/Vqn7aYOYPgAiE0en4Nj+U5VqRd6uu1Ao6Dc
2iDMRfydxNsGAMP4RnB28iEuY+owIq7TciELAxQKsVJkrN028rdOo9yacRZnb0gy
8sB6N5fD/x9mzJURru2XevrFQHtvC3J/vGWJzzB+NQuaUsVBiHAwPsvvyAU6IoFq
bKm5ghOww88RO01545vkjSB4p3x1wL1xamvbpviUGKBumTEYbKasevGCRRSGjGr2
1tmTFHcNDP4HJFHQKuMprEHRv3/l39MPAtptKzsJAu1qBCHq6bXVGRmrEIxsyLVz
y8RKSm0EbHw4K+VUGlVjJX3ZprcbTOix+WQ+r9UNg7Q5YRoCo99BScLnwA44JymU
Q1C6IbjJxJ55nvY0eCbAbOIRFsh6i//Dzq3eQ1JKhupfvkjmPkizkDLxAoAl3o8z
ChpltgVv1NdDU9bBqhOL/esS7memKZZ692srDzkX3FhULdkgofo27LPfFoLffhQT
yPgumI/RKxAE7mcOP4bkkwzczo+BdpxVjcnLJfWAn86YB8PF0d1uHmFofmZP/rI3
TG2MtQgkKTBrtbqFEt/Cxbc8UotopTdK2ubOlL8UEbraqXxtuiPSIBoB5Nc3ACtW
GUShNiCNjkyKloSh3BapaXeckBWjPgrT2OsgcZaSnS7r8YsrZvgXG9ykfrupYPIS
RBwbyKe5axVOnByENXjSTE75bqihNTs+OYP2oOvLt2aTcgBBDkJTMlrjJN+vvp8F
3429qkI4fuTcv9iA/0yIdZPQRUHKk+D/mJR7GOQwdG1ojcX+GBu8oVCnWanpVuwe
e22YA+UEbGiH625XtQ1WaBvFTyvViVJ8UCk6BZb/lG4d+27umRUZp9Amhu68kIIs
qBxu9Th8xdlfJyl1efIc7+W+6FUHq6nxGDEyc5bwk709oeqr3s2tnhowjYj3dbSt
y2EX4jDak2OeA510+2nuDCD0sm+gIZblF/Zew+A9dJWSm6xbu1Rchn05XWrSpv06
3EYxK5DwNdxaeMqYObjHyiyu5bb4jKvuwueZI3C61iNpcvHZ7FO9I2hoW3SxJBTA
E0++f/v7uY/Y92rFVY6qwrHzbryqn4GZ8906lu88V6taJzyqQQ2+h+gIt7zPyRiY
PzpWbOxLPDYSacwyykKxbNKF7LcsPG3LG4ssiFNiHRBwag0mTfilOLIUsOhXWtk8
DpJLLH52hreWzh76PK4Rha/No6qptXVjAdWVBxuJ7ncw+0MZoEzeGIfTOEtLrKEd
ukyrrYjZ5gFUFUS/bKsTO3aridzhhzwYs3t1CvdxgVpvGw1MY4TgoklHaePs9hw3
bmHPL18kwvVPxJSuGU+YQvwFKcYiJtM9Umy1NfAITTKmTKIOYvuxRrOg8V5QPQa8
6Q09/Cp81GhzG3sGN8UUughv4RMSdA+nGIyT1T2eT8DxqmJr09+dYGnMW3qZc5Ri
SheopeEc6hUVRLcKE4FqZp8dszM1deVLPgDNTeOFrpRHCyFTyNLCv4V1LSQW7296
9yDSF9jyu4M8jo7CcRz9EuVFu60YFatIUkk1xWu4IGgpONx+oEtgb/esaU3i+1u9
oUNQH3nnF4GxzEB84kyCkrKT9jhaayQJTNduWpsrdzgTULnsOqCUhrLtx1EGQ7J8
/GyYuTEG6pQrKMk1nThIdbgQkioNY8iX/ee3MqPYfU5NPWF+E7QZ1lW9Ta7JtwYo
Xq67+ZWU+jh373yqfdVsYMAxBRvPDKudgPvYS6rUxLkmgiHCXPsoXHPw2cpbCoCc
jIZvirhoQRtcjNZ6potG+kEGOokOA6myjlGbuVOkHosuVYTfler+WqZiVO3I5Eyr
Y1crcMQ5Gkzm7kRaARzq+QcX4nIDdes8yLRUoJxVSREMXf9zeUjJIb+AdOlalF6v
XnkbxWiIUgzi0SuBgB5feQV2jSzJZli9jIullDGj2o5F73tni2OLEMJlj8dbyfDr
ephLV8cilR8AomlRZzj9s2pTAOSwCiMi8JEzue8Bh7vP6dsz80J4jjajYgcT7ziV
eKU+h6/1cvWk4Ab9qCua7wzlzZIaKbYOcQhskRL3OOvs92nTSvsT1i94qSsIXqJQ
ql2vzSvp+VfuPhxCpGFH/EG1W0s43l8tgvcsLZ/bU/sa8yALxA+R8v3nA7sq+/mF
Sg4EaANSCYfps9Qimtn7B9vxDOR04xOIXIdwkVKrCyxc9ycHgkOBai0v0317DfLe
9YMhzzaTLHLS57Ubs8iVLScqDTqJ++7d0tpcPQXwsEHtJ8IUuO7V1t4undSB6SUS
jMoecJ4cTJvAumCAH1qjwI9nfCStNR+uE3WihtMxRKxXenKlHA1evbG9uEpHDjaq
EYgZZBnnQOckqcAapZGKZlPIPUZnWj45pu7Ly692XaaHt1Wj3T5QmmEZdhJTpcSB
dKmDQOSXA0oUvbnw5iuK1KKnMbSSh5HaXEPTU+LjJ1gqxdoTcab7khfbQmVsGeZd
+84QHHWEKq2JW0CRcTM/V+N8L+jiRo9xynFiv99qo1jRJ3mhYu9sif0ddcPGHI1V
BceftFSOIssuI7C5KoZ+ReHTk0DQlk8eKt8zYct5xBJBVYeSYwM0aQQ/MYkyFtUQ
GkezmkrNNG1ri7hvOZGXA2xyMcDG2IQekAzUTqd9YPv41I6SCFdEWaljX8TMD2AW
UmfXvM1R7l2kk5TfvajzRMObCDMaWpycocCsBHgxiPBlXsd0YBmQ8QY//EBogRns
dS+0cpi+KcaRU760j5kOsVqvz3RAtLKvxO4fd14sL2LRnMRVf2zIFuLVpBTlMOAi
1Zc9G+h9vwxhQGpJIDsQ9LIYjahC4TMQLysTIvAfPB5p2W2DiI1mTYvVneqWUlUc
b7MQ4SyTO3u2NGGa22Id/EeoLKQKQEya2w22IkeynnKBcMcsO252W7cIrNtBiI0o
Mvj6FUXkFqIicnxmvfSiyd/QoptD3KGAqZMSQ1HRNH0aMGpwTzt5WOif1cdeiXie
MZ5MPw81eeiwrOpTK+UCb6iD03AJEuGrYdJ+wJ5rVvv2VFxKUuargNtl35LTaywS
ms6NPWV6a+D8XdisH9BylqPplTnzd7UN0LHpbeCONxz5E7eULedzsAmCEA7YSDzz
0GyfZ8x2G+gfeWAFFIzlYWsBzgB0BaHbdbD8CszHXwWWq84s55hXaplGuViWmkHx
lKEU6qOP4+t9mehci4ta2qnjKpFFMHCvWv3Xd9uy4WQkq2YkOyfQIQZ2k9pOIB3r
5km1PGLqJGYdJpg1fySJJ+EtOzzxRmrZIcrJ/PHtUXsiBqfw6JNOlgDdo+VSY4Ns
dCZ8TDwKyCqV3AM2yx3FYTPYw4VGOo2vPa4goAKSGC/3ees+0bWEn1R9zfupJmk3
GNdEEkZLmGrlsUkRika814uAenu15V1wZ90y0PoQG215EfgunwdpXvKZK2ZGph5c
qfC8zKdinrZw7idz2hkYdoutKR8DCXGZY3IN1yrlU4urg0ZJkD5jK0Eb+1fE9WER
WaEiFhjjbPGXo5aNrOeo0Feo2TPo/fxDEgTSqoNumNArxCDTCGfbjzb5rI1usp3y
ydljjUDLoavAAlVS4LFeydNKJcK4Ug4mD3TMHMZoyxzDySxyueaZG6JX7Go4GA+m
vWMsJGY2DEGHLgpMG4ReAgLKGEXfcfjzipVISCPYfGIbbN7cXug4OP37YWuuEAB+
DGi5sXEU0sXkyW9BucO20qkq8nBXuiU7yMM+oCvhc1OkuRo6UKLI7/FvAaGRjYSM
ZuAtO5az3M0+7VtL3hEJGi6qxACUHhQZy2lqv0CsHH3yUKlIAwXrOxcV92xDkYFr
A0jFYyyfNSq4cZmBReoWuww/oXAYAs3Zb5WmNu7LB7XhbFLXmChkYY4awEz2hw4+
M6GSWrJi9JsfLlK6fTJemGG5qxPIDEhvkmFyAraMyAIulIroaUE3abmXaOTAZGEK
5D9kD7c1W8yMrOvo1YopuJ8ycESt31xav059Cei1W4lD/oHFW3bKvA/iBEuqj/0L
nw7o4WGYOIPfbiJVoayWbflHDbBkmsylILjwHFy6KN3kWXAy1mVDX12EQ6kChRQw
0Lh3PFLGcC7uKpEMebY/+9BdtO18BQNQo8c2GRp83lTzhQ4TM5OpVQTXtfXNZaAO
oyZVUOOkrK/WnEoX8PpKQ00PZelwKvfF8iHVcYMhE5tPYjxT4D55+RISgy2Xwa4C
DSgYhzdlZr7vXgFaKkgZEOJGXvVb4apZ+eatrovNSDMpUtI6T1zc82qyYAwDbKbc
NqZ2PM7/MovzJb/jpQiZqTkFUtpKZJ+t7ODFIR9FhQ62S5VeYz50Q0GktuWf2o9Z
uqXEqto3Vi2F3X4W6dC8rc1ZH2LuDoYucYPJA7My0TmTf11RK2o914/WuXb4JSRG
5aaeGzhjrRIOSuBuTJpjSAWg3UaTHuReCLAljekOpMfWbTWegkplhQLhsKNSvMQY
ob8WKox9+NgDK70y73Do96sWbZsiWolSPrgkFl0GWhOV4MEQrfbDU4BBDiS1P1Bx
5Qmnk1X39+aIqmgpwwLd0sSx2evwaYb0esCwUZcL1E398X49JBRtFFvJEfl2RvRc
Tch1rNZqyzGbohI4Z1Nc6ZMthuNKSYo+97tf48OG4yIO4Et+fmexd0WPdLE8Lhqf
wohZMZ9TTYXXU8ax+v3kAJMPFivz56PT7SrLjlUGs9BPp1s7lcputIJxO8YW0SCf
Xeb2qvjUGi6TPf1AdTqfsT7wdLXO3WfmfZn51RIu4k3WsaYnnqLPfbxtIYlK8IEU
RcKQNVxIPPRnS2vqKS4eV5iLKRlqdg8K+Ot+/SxcUFKK3E1uFpa4kKEWuSzOdfo9
1yKdijqG5bjn4lDe/IVQ6cnOprQvJRJp3FZPVkR6JWI0R1SNDml3TxAmH2hqX0wy
1SwbxuyMT75ttXLZziWBJSjFQeGe4OFC7cCJoErkGaMePOnOFOi2F/krq+HcVols
5j9ikdUS5/LAg2eZEAvq4azTxBjkQslvkBHplMEnJeDd31bhaOBaUVFPnssM7D6P
RqoXd/diURYKsVaD20f0JwaP2nXFyoV7P6dDjhGCZdClhF/ixLl5Mpl1I2909Bg4
h7FK7jh2MTVhYTv3J7ShROp3pxbOLBJmTjUii7ZmFVYxNCSvFz8Unq8robNaerKq
iCIy+7zdlC4eToH6DyF7/Qv0Oatd3qc80Q6ADVks66nfSvmqHd6IzrfQT8oYtnSz
YeVhbufKOYhHbEV0NWa14G1fmlef+aeNYwwJSE6hGCeH1xztzQHZ02qJDFT/LebA
jjQvL5Qp+23t8xflki0Vmc+iPhG6PBbxxjBlNRdU/vssd69pqzgjs8MoZ42Bffgg
Pf9bB8SjSOcUjzo/gFv5/YZZSqknejul2czWJ2TA3sFLh2ivoGJ3n2pw1ftNwjLJ
Z/HCJyOjkCXZXCPKMDFuWgJ162h8+AY19Lgr9eWmHgarzMP2BQWTgFh8uWIqUeoL
wECw118/vYDeu2lqsxPqGNmbpBucfQ25qEoCQyN1AGpDu6/WOSQtARmCVcD1lf08
TA1mBioXLkLuL30vghOUeTTXN2z8BCMAMuCCjXsAsn8qi6w26Toqr6E0WJa7kCVc
OsW/83Rfff4KMDc9gjAF9Zj+UHBigFlG3HXqo5whw3PXizWG4WbZzh9Uotjy7vgG
i+NGWP9SBGjeAGnue6lXIhmL7v0K4oeUqN5ZwphIZrWnRG2bajPgMHXCJRSQnUlJ
JtoTKNp/kZtyA4tv7pySUXeKtQnYOirBVxfVtntI60Krmh2yEbChGFkrD2pnQLAE
008GTx35bWnLLD8DHSNUagIbWNY7LJ+9pdUN44jFZ7E1P8VPdBtoKDOPrpUkDRt/
Dn2ugc0x1aUbCUry6HTx+/NnTnQ9GJWyOvFLZhoGAxV9n2DhYz30DcVnhzHsjXgt
t2IGZFBAtWVrO0tGNOhYFDpKN386yOGuGt+ej90RcO35m95SLkWJus7zFRa+5vok
iscI7odsxVqQdY+Zf1xzVBEk0K2G0YQLL/Zc+ewIUMGC814LJcHSBHflJh+xCzQ2
dzxyT68dlLWrlCGcgCBNIi1ZVhnOkv2N76zFcme78Cso2Y1CCLMEeaN3GIXzkRtH
qTfkwybbdSErPrNXVSJYqXTJ1oSbXZYnbS3mV+jh/2u8t8Zh4AE3gsJUb83j1Plm
TUSswHhTjELPennHxL1Kw8BwquKTdMzEpnPm7nwcxkLnt5wxRlDZYurELzpYwUsO
8466U9/y/7+Db0G5rDB3Xn19XHUGELVR0D8IkaTtfBaVG0kKzC3IMKx2LGMkcgr5
LdLYryp2CsEbbFQZue7aU4S7fu1MZjsQ4Duo4SqfgBOMiaaaZI0UazFeScTtrei8
O5H39LUaYxi6VVEH+cyohJr/ypK0DFRgclBo2gp3zr1EyKkdUfKlUJhnNH/bgbE7
YWAJS4YD5H0CwtnQiYIdWEQYkl08P5QpFiNtu28d/p4E5pqOP/phYcYgg+OrO7oY
Eeo3/tskNPMDmTcApZT6xdBp0ull81VKFF9mOzFRPR0eTpmU9gf9CZC16+MR2N4h
5mafx3UvImnCVvwOl4/KwAkliqQGoN7jOBfgGGNaCV+reh2JfhF1c/FUwTPT9oqe
S7ra8BS1v+DBST3uP+CyiaEFiuXgyJ0f+fPzqRquElP2hKImYfNFRe5nHDPW30JK
Y8trWfkN/IASFlbgXb2W6al7ZmiqGQGAKVOWODsrCNfHU1oNLW0LkUWBn5BURtTR
1bIJsuaQ4Kkejoi/zYl857iFZwGUITMBqFBsuVnvxEt1nHH5N49LmgNN7ovrJYVk
bhIIoa7bel9AJE6S8q3A5JPjfip4OYBf8/SNaMjzuWzned3r0Da3YcYubKTgXtjf
WEEPRnHt7oYXpXOMHPb811Tm/BrcrLSZsooTTvg9JgEneAU6g73A0xVsNGe45FSi
9/k8pqUI2/ul3akuUb5BYQ0fGXO/QJY33WxnVp3CrqadVuzpYXq/S6CLwKAaUiF9
J2Rx/nJkjAXpS7iHRzqcMfF0Hq7Ac3trBMvsVqJTrQEyKkA4Z7d7EmuAyiR3g4Hi
DQbHoOnPsAcXHBtFsiditmSCTERdgkhGikfTbNjA94MjbJJ0pSSZf6emfquCdqfg
4D7Jqb7G+3SfckoJw3qN/xcXnvJ9TucNe8pDQoZMFPV4PFg9aI4qR/fBil34I1Zm
2FGBL6grBDpcEvoZbiF3rL7a+qP+eGcPfkl3emhBenzBsUAjziVFQziVGvvyiN7C
CVrt2hnOYmzaTox5DP5t75mjF5JRxFo3gkhx/SzDgqk8HvGSk3/P9DGhaagiCLEc
t9zw4/8vGefkRvuyu3uyS5nPQ7LhEyvPWso0w13IM49C+tSGizCQpBXg5qVWNEaZ
MTMT5g2RPfJJHG/GeU7Hkv2ZkdBY/CGbi2zgjx5Gqo5MJYCDRzj3Z0liwvsFoMPS
yJCZMWc7QkG5Rg6JAZILT5Tnl/F8ahWQInFaZkx+Se7aB8JA1Imcw9+0QVHuDEPH
QAripUMPrNQcFsYyiUHF4Elbpw7Y66vXFVPW87Ho/OeT0RNVB29jYpSFyw+fe/9w
AyqKUB8TzHCokD9OGGik80y59Spe7DAFJb4aQtXJ0JEWJnovEP9lapH8JjiwHCEP
ghFxHQ4uAJmk+0iwMGG4rHwc3OuaAXLgwgIDFnzwfQrsI1I1ubsFINgq3UVxKHmV
Cowyk1CVOVNvMwmnu4Vo5Kol6agA5/ikF9Kc60d5Y9Lp+nvGk1p0pbOZIrEtZ3vQ
BsuQEWOJ9G9DaKPn476ty+sydXiX4Ltt7RS+yo3c0zRJ5fA3Bjjqjn47R75NrLYG
7X0lKnFqW2vMWG53QVCGpEiJ9SUv9q/MkHlP7VwmHACUmhYOG5Ep/WdZ9hXwmX6H
ioDkQis3OvrmkZ7y3jD5tF0qbxL6WdVI+kmdzVfad4cTn5hos4u52vTezb92QM+Q
KhgB4MHbuZCpIJNTV14xSpqHVGvmsudnaOalQapbLfcqcc5YJYT7Ypb4EfDfjsSE
FDr4439wDsU4BdqKTBudSw4h/aNAtWDb0hQTFBcRPUXD+VZt7MEk58CMEW/gU32n
4F6Dr9jsnlw9sZEezC8PeFDDP/HiW6vm4X6GJy3jSfcNodSqHiU6OCelOtVft15s
2BUuBaBE1v4arOVQA2AMWzwwnl+GD1nkcatpxPvMX1PteB4Lo8NN8K5KH2qp9ZiL
CX2JBtsYZ8Zn4IkSBhTbPYcjF3/fd4lQprjBvfKKzujrJhaGo5xVsky+stZ3dyyN
wdOZphm8d88WRaMLDr69LQWjI/cHfoyneUiff0QkI9nXOEJ+GNW5D2D0UlYNVoFd
n6JDC+1fY8FLISY0sBA80fB/cwwrkYfv2YvaMHY45FQrjFNbjdIc0zJvziHhspo0
82S/e/SjlowpiB6CP5aMwB1y9wgc7xQNFX1iH6mzz3JcZGdCBX4RayKycGQutoEK
b3FF28yxw8Tu0I04EbtTloBNhVNmPnUTCHBj6y3yGWN2s39kWdn00sag3iRHBTDa
8VZ26HZMEPYs2swrGRZNW5djGh4dd9rpCiu73gXW6l8VRktH/mIU4SiHbv7ncVD0
xed4jzeK9r3KVuxOqJqFdTW+rin2sSRx/PUmVMdFM3ykWwDEoTVNnzEPma8XMbpq
ETE0UagwTfrb5/OOLyOpTCVM33tYPuAGwR61ti+Sq9Z/2dU79toUcqudoPt1P1ZP
8SIX2P6jmNeTes6x0ZhhOMDHN+z9JNpLalvbY94EeKNAUb/NOqjCzP6A7YjotHFs
H3WBLGWJ//vph0Jg95MkyMHI84Oeeu1ke/+tbVn5dfBlk+E37u23xHLxMJ8YR4kQ
tIruh3vIkR2m8rVLvGC7hZUqzefhsWy4ARtGCJby4wjQigkRZUoc+uCg9KzvoiCa
fB543iIJoo/ihF7wohUNg+gZ9srDrxp8OQGrupnqAf0yjQ5mL8RImn0M8OSgHB/E
4gZmCDOqni+pcdLykm8ut1THDx4UZfr60u83VwWbTiZgkSMhF6UtcIsaGDGUSito
BUI70+Zk7O+lYkqGxlBgbMplVndfmVV52/+1eKNKzJLWQGJHBnDRXESGFPd9m21F
BHUE9DcwyhtCa54DR6PK3jvmimrp4TPTsqJgZPA9T87xRzSwDgAbxWOdUpbosSHy
TgiP+913R4l5e0GsjWWRSujH+/w4tVeYZ7s2b54+6l0x7W1WNVcjzuP+Gz1sK7k+
bNa+grJe0eSTZVuUNj3pAgpJUtdztLCDzCC5I0bJSbllwKl6vOM34qBiWFoiOvbZ
YlBZripjmBbRPsKjjp2qltAOheEd8ZtXZZHiJXR1WO/RnJ2EmnRgqBnl8GYE8ks3
rbo6AMtewMp4x8ZVLSLqqOyTvsTZNGU6uNk3jU/D/6lFcTtWPraYNA9yqXn2DgKn
uizfnR73YkQqJCRpjc4qdmAyDpqNrFUclE8Sv7ZlF7KnCqeD9hJWfMOsetBSRFWR
faqqIAxLfNZRuf5wMtdU3V4aY6sqVXgPXn43CsFXQ9hK3ZIKZNwvi1nyKwob8Ukc
OEddBBbioFHEUDX64wZNb8CotQrug/YhJbN4i+J8D1V83rtDmmatMJgLqudhcBzx
4e/7149HcSfrjtys5vCIdxxK1nSYAKT9+3nHc/J5bonkFwND8CUzURwBk5od9Eg0
ZATHIg++CYb/4timR2ys8avyPgPFNdcST05gxpocp0oZcBe/7ckc9jMp4cMwnmos
k0S0ZYAVTlectO4aSI6TY6XQWeCYp++WollxJ1KHiH2od7yYfrDcQPBSqagIv5M9
HLmWbTS3yttzCAMgwY5T452Fl6KIpC2ynfdVX6GSEhqZ1QdLsYgpHzsPy28xGa5Y
bVAGUOr4dq1rdaEZXhafKVfXn8bpp67dSWPNi1Ah24kBmVUXyqCrf8AXgT+c58Ho
2A3u/bdcEGUvUEXn+NIkjnXTkVnvtLRwq3tXASJ/F3540HMOW4J1DgM7LIRr6TOf
wLc6/3k7YVoemy6bcotAc66tDxVk+IyRjuLgDKwsX7RhwvMtbjfBI8yjd298LzjV
mhLQ6BW62T1Cq7eEGOV1Q3PweoYMFiupmlZk24TWTCyC0bdIZjAr0KfFy60nomc0
g/z+okjhZTCF5qoev5HA2PIopDfjW9WwE9ptH9AAztUpmwysJJ6vIKt2FRTWp+tg
Tm+EDvJrj9d0deStyZsa6a0g2frPIEJiSBnx4u9me9Yr3li5qB4quZ4Hgy2MxhNS
jhCJoR/P6IAHBeHEjqRbl/e0hovLwEV8jDEJYM1FL0u1v0irPHao56PS2cXtD2kl
zn+D8N3srrgwFo4U0UgGA5IsEhbZ4wcdnwvRaRzZvnfHdVYLDGcwpJdcYfQ4nSlR
7wfM17SZUi3GmgfC3J1UGfiqFXpTIw9lZ9/+s/xl7A88iUkMWVAXoiFqpu0i4ugR
tV7z9fpvs3qLGSJ+cviAONK9Gf5KMuz6kel7YGxXcTcqKyG3qiB6mjdF8kWxRpkF
em5kaXJM53fHDuYSIlDX1nVvgzJbyQGdIoEPupL5hHYvM4vOOe1frDgkTqMyF8n7
0YIwtm6WHwbhJ/Fyb4/Mh1Ks1MkpCducZU6Hzu9DfYaRZ7z50u/AT4QsNbHzIkvq
4h//ZunvKz3QbwtXJK2WOuWhTLkjDL3fH48kgQrT5SdjrMatP3vlrhOoqcrjoEzT
R6m5vPpkJLacqB1TXX9WjKKh7qJg79nY+yu9yvUqUC5/bdtslEzsqcekvn0IJcF2
RqNEeXD/QvboeOkQas/HzXU9Taps9qLPk0Brc8tEi48ZUXTg3o/7HWKL9X4Z9X2a
6NQi3gGDywp9QjiPrviQh33ErMFtfMMvRX3aST7bOn8XUAcBkFmPPXRYHcNpmK9u
taTtcermsb8U8YimcPqQgpUctyC0KeMGKEvFkF5hCicZNkUCmMn2wvYiZKvmgpW2
6IyD1zUxwdjOwYdUzmi1eJKHRNtDptVKCOP5Jt8fGMQrQY1dn1kv1OlTqEM9HgYJ
uiouZacWTCFN2xdJybog5XpFfbNha3mpXIcyvoB0qI19ipV5rVZCqiAxoIwHACPK
WUKFJ5jhO2KiB3rMXz7MetatMZ43QzMXCyg1fHWVM/rpuFwQ1VeWGe380j8QOC4E
K00vwkRo7l2ft0HmI6FxQ6acIi0LdyfUB403L5BDUy+suIuYGT5o/9yzSEEJyVhY
Z0nuFZvwBtkS2x9swvj6Y9JlA+oowIfPwxjecfJjsIz3L5fxpLZNaKiSpICWudap
PLtEMzzeFhtuc1LakNaNoknUVRWbj1/wix/h90w2yPqZVLwGE5TUpe50GygviLGP
Me3wSFl9Bzm/s8rjEGj7BvtR7Z9y8G5ZPWne4vkhph3pdqoM/vRFkOrC3goji3qS
IeXKd2ue5l0jkNCa1KmKOJgh4uxHDeqM/Rxtfu0/IJhDIxuz0+FMaMd6h8GQcabu
w2QD7NwiLP/1ZWzCnHHCZLUXf6efKpm1tTwLRnCFzuLGsKn/xP35CtVtpGU10w7v
GKKMsXhnF30cGR9K8QorSdHa3dmyxOGh5ajvQhhz4YZ7DcKZbBUJhDO/SjwY7zab
JS+ncs5CIjXIAe7hCq7mCSFlYfRHceQD8ZLOswGLHX+cj5w4dwDn6kGK0N4aaXl+
sJBcJ34YK24xHHOiBoKpE5dn2WyPLUC89uRQjfFSG7zQSSjYkhNba8hrX4slAvfx
z86Ho0MgaZOHGeYoLn/oLN5eiu9Nmyfdqd3gu9b/k5DxhXGa2abOgciExvmCS2KK
R8xNvGo+yirAp5BHg5YRjnwGWdU/ccxh7tvSCu5zSJR+7Mq2QviQwykgo6zr8zHs
qnBG23dY6Zs24/GWyMmGkvcyGv45ygYAkhE2f3RNl/dG75u7r7lwmh6bpCU4dzCm
vbPdKduarypBq6Ejnx7HigMRQoLqCGWZfIQXNoD+7IyD5A631XB+Z3aS6yWgbbmG
4NUflrprpFXV1yLMuFdrU/nsr8a8+JSnxokecvOu5ujHFJg5/1x4gY/e28IOiHjP
CzjR/5w7Lr2YgJLjE52HtAmV8P7pbehlv5zHJU3Y/Av+nK12YhwqG2ivFlZTlCJB
5a93qWEqf6YXEGP/WnkjnRcJjw9fa/zATGlRBXfHBNSmpKYN2AvgIC+YPIv70g2K
xJbYWD7kcTOHw/NwW6FVeu1toSKzYomP/liMVTkgJJrO8zKA50wPw+dseCjBKKpm
OnNKemcgKVwa1vhOcPbPLl6ZSGLpEgzYrB23Tv9aYTLZBsJGn2Y9jeeh65o0DpGW
r3Y1kKwYFNejpOZnAUM49zRtuEFI7AKwgbBCyFa2dgEFmOakfAMSW6db2errV6M5
JESBgV0Rs7OyW3pH5yMRP3RZRw8lF542jo4NcW1cjPwzMbnNjd09TM3jAATbmMkQ
2c6fOC/OrPyqehLYs8Z6Un3zhLD9ke+24uvo3wYBqbD5vzpn+1bWQi2u8FsGviID
UpbHbkPbdv62yE3SII4z/+FwQmv0maaL90JMuK75DY0oui2szgHokksnr7IpvlwT
AuZuOZVEzL2efdJVtCqhIYl6WqCfG7tAPYpNk5k+WT8ReI613LDdNOG5fkJbHbzZ
Uzt+++hVttudWBwhdt6azCIY7v1O64Es2e95liWl6ceigokq14yOZ0nMUsjvLDMj
lFvl+euv0yUxMczBigpFxX0ESuCn+4uO1101NW7QwgRpDc6jkQuGixKeLrrrJ8oX
T2ltn3WrvJuLHKI0QydYRTm3+1Tu+IwezqfkxQfmN7cHY7Zvt3/X3SvIdsiRt/8R
Tgbp/WVAYe2oSLevWK1xbF/Pvp03lHgIWi/sQkUdp3w33PF713Ax76UXe8E8L+L/
Uz3U2MnigIiHcb9W17ZFQj9cWroHtkoFZJXq3A5haruCf1EkmYTe2jMMjy+AhKZt
grrSgf7pblzBScwzYsDbIXIcFYG9oJeHewUWMUyB6k+7yFDuxDXsQrsaByOyrV8e
BI8oRUCb7w0fbbq7l0MfXHNa0TmQKT2hI6Nd3KnbOMhe/MpHVMKhNIDNpeolMwtz
GpcZB6N27hBUSf+Uo8VF4hmbIzooU8/fCqMhsdF+snY4n87E7CrgPZFrvyedTytr
ECD7+AirsMB9LCZqS3AGYvGjb6AydDu9M4IuTge8IOQnijt/FtFeozVAHPwr7PFv
TzpRW0GgHqhqW0AMIa5W3mmRAZDcQ/ojHfcIlAoKefFrWaaaRa7Q8tC+Rq9B3wZU
Iey01IeMT2moI24bTLURQquuGbUFDZbk8r7KIg+rWHe5T6scgFTWcMnDUzctcSjJ
tBi9KPtDtEKLPeTekprv0Vvk+LDvw88IQsT6zBNMJgZGMX1kVQxKrhebY91UWyB1
gZMtxMg7dwPY7BNySMpxsHjVvikLACI1Mkro2XbrittwqGuLmQUX1a+Py5EX/Vg/
SqjOwc0Qm0Onh9wyVWjtwg0jLOh/UhyuzAfjVTM7u6Ajl86uw6v7lMMYcZwKuBje
ZN/GJSaJJk2hEJAMvYya4NgSNJZydVM1cRILgfhvJSyqg+NK34SiVqMMWnhpMecc
2qovfhvYMJU08Z5+HbvGdu2ejBogXZqaX7hON+XYnxO1Mwt1A2imzT1dgasXyrhC
fj+WpIIPDfBOZudfSv3a8+XkBmNB0mZXqVWPQfgSfWVGxrdxNpFV0YWFb41NwT92
hRHF6l4gqTynK5lWd/NimRb/ogpFXAOC1Zf+npalNYWu4M3lEfJ2d9lTNoFKNcnO
/dPwIxak4cK1/52B1xKWb6CxOJM2bDLLyhUgMJwYQGi+DXWrlsQHBX+hagMi5y6d
xM0yITSf36YdTs0n/HIGPi9iMAlRNyyMu4yY7biLV5LeGfQM9r5fyR5w7ARgWOQm
IR4kNhdCWsnL24i2KBmmMzVemP5VZQcD+W0yoJUGR4mvDuxum42V4ZiicWir/gLd
YpH3WoM5PV8fqECaGxuHvaIPKJVFFAGyMQlYZus4cLDyP0RFeK3TO2jHBaQHfIqw
b64dF1a8l4AdHMfd2gxa1Of7u8B8YhlfFymauehTn4UbPXXhboYA8P7uQ4Tg+nHE
TnuKHVg2+US6n6MUaUifqZlLm7lPmXQk9k3GEguISTloFZisGW9gQwsinbRfFTmO
b1iPmus5TB59yRc2Dr5ReoGZDhpF0MTKQPDf3JcjPga79kLDDFGYs5gJSp5L+9o2
gm+/+ZrhhbTmBXIqSGO7UPKn2rkMzo2OJULY9M6Aevzt9uGEGo8O3KK1ICBu/otX
uRiNPvtCrOJj9EmAavGxMh9446wDy18XpNsKsv2UP8pKUDOMxJlP67d0Ua80VxPr
hW1qeigjjNjyAz8j96206faDmjbxY4b/qVSqpqa1QX+oM7nRfiRSPkMYvqJ24mma
QXdVdeKKKyVO2IrcysrsyVocecUWAGF1QNlTYvVIKdjg9qHST4yp63VIBFrSu1ax
bAyz3dWCGKn7ocxk6hF2J0sJa1NbNTumRAQKGvP0BHOHWBpVxgQLtmobEM/eXJNk
ogG8gqsJjw6yD6kDskCeQYiKwSXCRTxw0G78OZDMRITPlvaY2tcrIfRpynKxLM1X
a0lk2QFsqP8uf3WsR8Ssm/w7tOn78KvvZuLFHnmtHOHIokKMGPmqIH7yLncWsGU4
tTGJvGijbXHCfZwMKkajL17ZuDxXDLR47CMQThDzUL+DpLiI2QXmnh+InQm3MuUM
Gk5YlaaMZi1aE57H5bsclC7SskGgmygt5VAbxlu23HAPpx1y+BTOz1y06U2guC7v
fgcfGeqU1Ye0fVmKNOaMysCGSA2Av/6Q6GGg+P695SqAzUYn8QrN34gTjtl1gNw0
JpBS2eg9OgNv6syGFLELqfxLY9yKDGtHdFW3QYxf9XEX1B/KBzrku1/I7FYSPqoP
v2ED+UERloSz0vQooNk4rd/aKX0ArN4c9DeRIKLizRdPOVoICH2WI9HqQjEOmtN/
AMove3zUu4gcLT4T3tjaBbo5mx2AXFEwF0MrzWDwxeMq1nI6L+tX6gzS62QHVBgg
ylzEAABVJiG0W7Mv2bBjn7nByF+cnwLT75WAkYy+REbDyXBmwKgSdiWhUD+ElJCj
sHiCIokk1OmRaD0CgWNegHz5pQX12LR/CIe/lC3mfZRpjc9RevbIp0Aaj2cn9yGs
tl3OgWpvev/RNFOc1MdZ+Gxg/4Ni5wcqvyxYCT8GPCQbUkLDsHlMbpv92oyQFqH6
gUpheJbPHlvk5Z5lmh4ldsbeTAuqmUVk0UMHq7SZtRLw+wYvNZddXnvfBBLfFE/r
tpY9ccmeEGudUtPT79u8vNl6SVtTIwnMNaaQkt9yzOoAudI58lfyo+Jw/+VTE0UT
NU0h9ZFFW188gvzC/CF/V2Cqo5r52WJRMZGrldh9bw0qdBQ7r+Os/yog/pT3O/Ma
2AbB3uPQmUnhYvGfozN5a51VxHS0NfuI5E6rFzlObDrlimjlz7K5vChXM+pn/Dch
gPPf3wf8qeq5nkrirWS6ccP705TNdsfm4EtWZO9MU6GPDdudEnnbXeR2zyTeekR9
K9MjrAdxw8eHPcjHwRgaaZaH7abc3EHXTL3ACnIo1bXgIRfDgBM/wNPAHa53E3VR
Nq0+2ONwWLI1aLHDFJ0eczK7lpcpqiP+NuTK5UnD7cEEzkDonZaPLOigjNkmNZo1
irOc4pr3ZBLsPIrlxNvJQ5iNYpFFFPgvPwVcDnH3SMWThogIAbPxo4YHLchrnQpg
hOAFODiO7HtYMK+fzadJ7LcMbt0BrqDJv6erQ85GAlNWM4xVYK9LnCBxE2yqNa5W
QjqDNXQte41sHkXsH3s5Fix7MHnYlfXuQHghCDbfeyXnKb/OPdyJgpIJvMpODdWe
zF7Gzkff723W6M5KOWFeERC4qIvYij+mHDzOVr3SDGHlVhFvIQFvGdU4Y5TrFlpn
3kchrLU+j/EMdt5LyKa7MZ/2RcFJlXLTAHh9azMel8nC6+Y6mkKLbo31HRI1Gc1f
7kYbh/7S1QhAbcgK6rzWf1XUmMa2jupG5f9jA2njbE4XR13TeExXbMw6c6eIs3vQ
/h1iICQMWdeQPR8tBjkMg6i2Qgy9OZbuvn7Gz2eIvhLEu6Gcf6ByBThcTfTo27Rw
TmPbLFfOTCudVcHNjI+JRujMeCGsE2uCxFzCL7/hIl+1p5sWZvJGeS0ey7vF2Uqc
2TvTHwXKFt0COtK4GMHoVf7P7pHUsD2r62jIEwBBQDcK0YlWAi5psxIh/8eCSFrS
hOfYbH1U5oG7PIvdYXaovkErt+/uII7HweBeuw+AfB2qF38WJ4tx4dKiNEYBqF+0
5mJL4NkO6otYbdmTEtk16sjo+gVoaPCyxucg0ihV1xYmu12jiLlqWSvm6pMj2y9r
c4UTlxXkBptmmWel87gqQNgIEhCiNg73tuatDTz4n8AY2tedgLgYMMrgvc1hGsFG
qPpty7gN3tCEJtLC6zcrQ6sRd6HXhcq+2ck2Oy3x3SXs5ujydkPEqm2QIzEfpuo5
ta+DWp3tHqhMgv0QESN/eky7nLo1+HvC78zB4sbBR1iNLU7zN2EBiC9dB87iHcWd
pEpkaX1lXLYZttm3otKF4TGKYyFH4Xeh36TJo9eUj0F0Q1x/ulgmRIPI+LDwhiMm
WQs+4SzqK1HufVa3vEwvxJzhyErzcUq5RqeP5xHlGwJoRkvW1KELfFnIWwB7/kws
qwrNw4HC4kgf1OfGHkThcFNLpCO0L4cnzV/fz0KiZvsFdxfEF4mS6JiFccdwdDPB
lxvoFIaMjisS+lRV4jTEOl6RBzjId69nxwil3la+hJCLFLmfb6Gc8sC0Y0AxRGwB
dJ5q+8dtWqJMSyG8kDfBAnQuYpzSm5fnFGovZyyIdrqAvXyW8iSuuLFneZsUWAbB
kOKJno/15EPmc82D5r1h995YrOVyPbdNv8guf7X2a100tQltXFP4hFsr2oLMXum5
Rtd7eSsH9+z6CWkPUiNQm2Au5RDnmBeW1lmM8VuNzZCS9tU/DP623Iv/n9xJk4ip
i5O92XfqbqKh4aga8Rx3ZcaAiKIOPyB7cui6MW8Op6L7Mj0N4fkHKWhVXALl6xiQ
maM6kyKSTSJhtjcAj8Suqw67zIvj6ffrDrgo03JNsWPYru53w6JOI4/EGYVoVHab
oXc/tr0O7HTy69Dsqm1mHuSxqqPXqE957+kWZpAoGzqlM5sfcrS2Tnh9ctMglmtB
pO8pVdVWFfbTMbUwLDEskkeJ5EgzkGOri59EGlMzIrrg56rYbhLPmp5ploajgLY1
QsdYGRpgZMe3RTa9z8Ex+45GmX9qEyRrIRJXo2yi22NHmO1Fdl7ibjRvmyBCa2kJ
c8IOLY58wiqmiBaym5agTquAaRglpCe9XlElJGqqrEnfNPulQU8yh9TyaC2AsjNU
uxQ78PCZphCesNOAM5oHO++B9PNj5tnzTOo+lF4HABGS4VIsQsz6B4NPqEAGxOHE
w5x0NWN6srGcWAROyXv0bDpgsFrQSi+LcH6MT9TlCKtg5GYiTLYis7eUM9Xb/tQC
1XjeOXzQAFApssDRpr8xZX99wyoyHjD+J+ZDPtraheGm5Zu5ALHxZ7YG1D4lBg2f
2z2pHFzJAEkceJjHiybkw4BpjjdgqeJPROlmSuHwCtugRDzpJapMJqpW6M6Wz9dV
ZMJUTqpzfTs54Ovft5QPltfhcOemLWTW/iTrMblHa+A5fwdm81AUobhtvqmkov/e
NLAd4fa7HWSN5VSKxSNxHKTB8J71w9H7b3rJAaD+v5OiryYmHimUp7gQfPhC6+O+
lH0hrsIACC35AlPHeZLYvwX9LfeCWVF0fwtMHuqfX6kqN+eZ6TS/Tfk3cKjQVGsX
7nBkPAOn5U5F57rRLCrwaVA/F66BCl8xyzZt8GxYO/eNRnn1wWTV5yLABdMTcUQQ
b6FamkmDQu5tEXt5SS08RqAyOgShIL7kwb7u8ntbrwMckhp6Y9UV83crUOKf4U+/
OCvs4EO48+zVYnXcmjryDwC7F/qq2TlWc0txEMZVR7c3Johc2QwvfEW8eG/BxXzH
m0cuJ0XFBMWWD0gF6sXYaltKCUwbkWHjvE3gNs8+zujePrA2em2AOT2zlo24faRZ
4w9soDW6p4pe8N6nxnNYl1/RzMt0kyqpHV1SrFbSoTm3vDG+p0GK8V0Yr6If/QsZ
6+mt3OnMw7DBmXPqqioKisF0SUVUbyvxmYZrjPhjSCZeZZqzBf3lIJSLet/3a9yS
TO3L7AYPNUETQPch2yeAvzMp4HC3eKMatCrmONRpU+WjbIzcmLhloVWpByuBGjed
L9y/W2HP3BW6LmgGcgSrAkh2oenTrfgHETT+lshEHxeVEw58USL6w3uqhce4OJVL
V7Z9zEd5P6ZAn/ZwNIRG71x0fKTSeJrT9Z96W/meyDnLY0BT94A8JfvCCqx0gTOv
cWJfDsF00vyIfZCG4S0opAXd6NPbXFAr2SFkXwiGoyPyR49QNO9EyCDSQevN+cvp
iMnRWuWNSvV8oyR3xxydrIMfUNo6+xBle1Gop/8awKjKuW14ho3VrLrQ1lyHz9Tv
rYS2tO+eu5dDC68hN2uEh27wirDoe4FEmrQviMPHaQeXAA4NFJ7aVuQn4TjAzJCy
kIXHJ44AS/1+KK7cFrrhKn8RKA0Ll8Dh3XZGIISYQ0URay3EQBENTOBu1UKX5jHP
L9MKnQ8eccwkPxqRi1avlVK1ZNphkMSe0FyfNqZfGYLwV5M31ztr94KDGoiKVVdX
rC5Qoo0yzeDD3F8o89UAJbtUKrrASouTR1iv5CBtPG28kDmQXVr059xRC4slg8kb
IbpOvCV1BeLQchq+ubgOABHb6gSJPCz/l8cXqnyfoT6Ls7Xdt6uOtWiOj5ZXBuLM
JaBn4ZIrqJI00FRjW0y1K5PIFkqEVFKNYcwRGyXt0ioX6zriGM5uV/PNpRyxXfze
LuYgxRfjPdssJjoHwpyY9GImZlCiJKEnNiY+fTLnZRYM0NXEKRggXJq00e8h8VnY
xwYKuJU8MfIsh2kB4JgOioEPzWj43ASVZQinU7lXMbqu5a63/yo+zYCyjZGTrAo1
93DPbwOwAPo/OOqagagSaFZ9gTSL+zSoW2v682VuFOTJCX7V2wYL/u3PAG2rwxK0
9X+ar2vXIG5nZsZ1ERy73cHwYKPpTBrH68qFQ2von2epTetZ98Yo5Qtpg7Zz6clb
Cej/GrXcyVrzVkU2vWsEyHB4BtSc7giArwjemXOeBwoeCD+im+OZn2zb0MNiVA1T
zpcPjvB2v8otn1k+UnE6PN1SiPqfaofiQfIn8WqbWk0haYOrUKBFfi9DUEtmRijp
qf7WXvVm694JvIW5TbZVlDzaZ828vxluHWW8KCXC4210Puj142dRwSkIhtYeWLbP
t8IU+hoy5aDr3UZAHQ1HaujeTrGpDd5cKr6EQG/4HdxEuzH0n5+XYF58RtRRUU0w
GYRuz2f2AvIniUKYdWwx/A4HF/lOcCHQeb/xUS9e+Uy+gsYvF5nacBBU8vvvn9oD
q8bqQQZpSYVCahQvUerOaT+ZSmZtEpRcHwb0xus/DW/lCJhfA3/FMfeNKU9r/pJB
u9TDeph+wpMMqZ1YYn+wk+tcJA4dvduF3/N+rdgobOzSos/VBCiBfEbEcANSfRK3
ykQODKjqdVqrHTH+MMqvIwRx8r9mEx0w87L16m5U49brYRmvf0HQ4h2zRlHNZHvd
jdhz8HK9CW6DMc7Yy+6A6KTP2qh8MhxMdMEmnajVjauF2tEnMVOdYHWOy0uRyDbJ
wQ0/crQcTVHJJLKGWZWs/MMBIYFDUgHY3DN6XdyGkGlBfx0WYhY6rW77zPPGUG6h
1DhYoerhHiMe17t5+d0vgjWoEOfU9rkcsHTgCEjFrHoQEshLPqn7Pa5G7qiWhJyJ
NrXugHQaeRpElrDYz7i8OH9jWjX/VKs0c6laW4ynrPiyBrsjNySj3Q1Ag5bW7Q/9
TTOWdI1cCuq3EC0B3RFxiTGyQB8UzwUdVsCDFhoNovhaHLSLh48LiJHQaMPOveSt
FD6seETpIk7TPxt9hQYsofuID+3LG1cTu/uQijyT2KmQaTF5XE+GrXyQJ65BptcY
3qq5a4PMQsEqUy2a8IWqASUI3lU1y/QWWGJWDIskRApOal/nOlxNtVfOwf15BmX+
Ha9CZxl3c98o0qHnh20hOY/S32TmhtNpUIf4ybpBT+fTL8PKY5n3dMpk/+u/vOU9
tEbFg4N2X6r/HhuhJFjT4ntUhDwaz1dvcxuBNO8TqkGZnR/N2WzLY8MrVpUcD0kF
xRAbK+psIUazKsr0rc+IPWcSezOqHtv5QYiOC+N0q3mINgjVhnmVOpuOPVxOlF30
lka4QPSwW6RA2Gg2+BDRmbeCEjre1hhC0/gyy1uyMyxv4lCjbIAC+feQTxIcyTOs
A3JIx+MCcEWR9I/LDST5Em6P/nvpYOXJTDBw73OHH/AVWcUFmvI2uQM2bRG82Vnj
9RfI+Qi850tGXYjSa1Yr8dlesZB4cqdrrhcSSddXOABEgDViiQfNxcrdooynlx7x
kWARt/Sdhrjof4h+EkSdIYgarlPDiS4UtN5/f002zZFCVHB3GYKObMukTB2eJzVK
5R7ZaH3I6KUmHUQzRwXg671oqhUYgSRc3yoNdKaK4OV1NZxKDWHzVYjjpdlks33K
5vMRv8z8VzatuIqHRrc+kjdr9bV1+kvrqTTstJYHZXaW01qZ+ZGWz1MNcokkJx+E
3MM846iVkd8fHLWpxc44DPqQrlc6elDAyPWraBnH9ETegbVPXT2DAACz0leBM5Ls
G9VNJjVNulyntx5ung7MMY0KtlLw+78UOjfsjpQXo++kNSzh4ZvlY0WVofKMuA7p
58HR3k72kiRV72dkVBI6GIIABo9Mafg+PyS3uG0zdIT0sBPoikjYfCF0eqA3v9dm
b7VZwmpOLkjXq1F8Q15iRFmN/ET7FswTd8kp7DOiyrbMe2qhxzYwfeJUj1JGx+60
+a6WVSrDWdZLbQmLdYs5QZH36Anz5gFLdJ4lgMIJ1iLLNRbpgATdUj6Qar96F/ba
0zeTKvh7y7aCVGCkjz3UTXT4tcHgyD033+3Az+KAhgQbafgruvKbZ1Ncm9MH8GEP
Ob6NGHvSKOfzcFt/a0q/wbR0tnzlFUr0q/JKjoLJXIxPI7L6ShgzoLPW9hgzhXmY
usdGJpJIsxRUwLY3lD7nPq46wHtZf12BL8B9V4kP6CYrLWtnppg4gkTrirrm2/Su
h7Sttl+awbPLs+2dDijGnXAMDViJx8dS6Waf/R+wd5pd7E770EsknWxPyHjhyuCg
pTr/gxHYwesvOhvZuWbW03NqB431QWTjzlzAHKMQ42mhAkfHy9OWE5PvBOl6ZLej
6f2oG+kVppLXlkts652T7FDk114zXMIlnJ/6mSRs/LKvZ2XBZiAccqn2Pph937M9
lmTmbDiTQwOomLxknmkJnfF2IlKjuJmDHrTO9rx1GjhV5/MH6J9l5OshmJ9PO9Ub
hdcoRyhW9cA5c5flf3coCF4e8NOwG9rWSyuTwsPP0VaAr0MTR6C4tERfg+pWSlGt
9i57uYfab4hU0P5MybWekOzTpVTq/xNwc3ybhfdw9amKGRnVFFO9OCcOvKrJ4who
n4XBZHDH62oESL1BRSSsMh0vjZ9SiN8ku17OxSRM+cDke/Ae1wj36h4VLqcpTO5J
sPjTgI/UiXFgWcU3sg+apjBqqh3zC2BTtByiHfPN0Spoqz0Kv+UAMTsxU2PujX14
ujVYsWMJaEh1C75ida8FeWyZqnl92G+9J0Gu4nkEn0oxEOJY7BwUol/w8jhK1w63
wOfTe0JTsuIiYwNKC/s7V1sWekH6l0s/xjJCv1Wf6OxLfyJz1qXUnzw2bw2gxe+4
fsjaOrcojGDzzeJfbQ5v09EqMSWyBmbrfnS7LiwWXzM6TQQNG8z2BdrWwni+3Cwo
c5UmRYSriLl7+dYOR5bvJOvPvpyNZR/UJkCGcN/vjw1a7WiGnrcnMO8DlzeD6mkv
WEKprH94sSIFFO/7zOc/OMFtZojl9AeCTjyqbvkSlT9ZCFd7UdYQ8YcnyNfMlSus
HfqDNwoGLvP0g3DYSb9iumK8/ZIny97Be0lYikocTEMrTUxUyMcIu7UJ4wsJrJn+
/kANdKHSq4il6ZOOucfnskhluMTw4fS0MfolzMRCPHhIqe/HoK2ZpzWzHkAG02Zk
AZ2IwCeSkmjIFCCuTZnXjqH6nJsfVY+MW5XS8oR9KyxMw3ez0kyZjKy6L4nYcxPC
5ynDSeVyC952VzqjXw2aWz0Ns0QnD9YzyYQCbMdg/L6+m8CfLEBJFAK+lGD7Tvqz
8obv/OqrQN0pPMeQobyhd36v7/LcvIc1wZwk1M5lG0Klteea4Rfy09xpU1Dz9B8J
d06+hiG+8PcqH3yiUD0AU+zOd5ohNJEQ/gC4Cn9VgwNLmXlMfTbltF8f0f1QiuJ1
L0GI+PtCldHWJb/IdgAQubnzacNTmcCnttrhCq9WkWCd8NFv0rpfPnH3lgYIhNp/
Yw+U2n1nCeWT/v48XItzyvnZZW2pjBAnsgUWHPn412K+Uny7meVLGMM2sRk5QhDA
YiGi5B0yYhuC3loGx10Zqrpz3uD8h4pOX2Kjt+kAVCcasJ8/ny4QbQU9wX124mL4
wPmzBw9w1JjgBJBtDyWEtCPdfiyb0Ju6kmJ+teyzZbAaLJJiYXvT5IoBaVqfyADx
SC0N/DjIC51CDxco1hlTluCcIif04MmmKntsIIv/AbM4fh4pOgMQo/Qq8th7EdO/
VbHWpv4DOXDt7XsyKBMp200x9mdDiSPmVRZVBoJcvTrg1nZEzomUwWs5s5A7krue
HA+4RYhsHGE71YWov8DlZIfkNYfa9XTEgIwp5ighNQ3YpA3HSMKBLA8yw3EyOBNp
2ecYn4cSr83a7fWiTt1aBfEJq6a2FujUKm76I6G8Svh3sInllTHjOFuOwL3tWmLM
DqiYLFHE+hf5H908z4bWoh6vSbtfNbkJtrRuc/mVBBKAqhz5wgoLxTVOS0V8FHaU
bdpI8Ex3KCoekkdq4SJO4QQhUTPjQK1YlREQs2/wWnbj/GbxyZz/4Fwdfz1ScOqf
QpNKh/HXXOSoJtdHCYUliyK4B7eZ64p6pgHgXuaMSd+8ULhFG4VSqax5mBF0t2MJ
STO4TrrVlr7xJ6DDX+2SQOBLWE2Al+YsTk2yt0/kL7BX2yxy0At8qHSX5BHEHCis
+h0begbs4T/BXHwa2nhVHBMfP8FWx7jz8Le6hJ2uO7T8WurNY810+ukkQkxVo8gx
sg+o35XJDhZYrssLH/7xEGWjwph04sXBvEcnV1WYyLDbTL2Pd8sCwRhuQz0dHkZI
KbUZvRw254wPdzZhufYkA6E1nb/tV6tumbrhhprM3MpajYs5fSCCWAZD0oHv9D9l
TckddqBpSXk3DFMyg37LSwU8cGo1Opa93JVjdC7ktN9A0A5npQiYbiSwFBhOpmbl
m6oTrVYmQgF8849O1k3iLhXwkwSXl5KvikkD13ayboOv+yD6uXraRZy1DyAKlwgw
Ooi6d5XYQFeJIYiNxqeig3EWlZS6OQfR/ntLHFatfCga8DOMADn1AJrifeCVXVWK
S5DKNApwcRJnEp1XDB/UkHdBTlty5xE7i30G9+0zsLIKG6E6XeuY/Nn1ofhyy6Wm
7WWMTOf3uIFdTRywmnSNPdvdlcIC6cToqOYwx0o77isXZf4ZJLsBt/gSf9CujbcT
8yUNi3gsd+jqyZ/enGUnoJCdmiKMyBk6oOdAfjSfRsJrFVdl5U6Z25ERt8t7CEac
7iXilKSJxWcd542+3h0WxBz1iOutr3gCqrxcf5g+QeLBV/QRvPbK5GponqfP3Z4i
rnJWYGx09mUvWCq0SCTzrHuFecV3MEavRLORtLNIuecdaX9q6ezT8q8/tN1CeN+I
k2Ow+iDWUuevajb4ALHn6AFP5/l4cb8vV/un0dHgJdb/yZ/iMva4pqRmaukeJMO3
lygYBa6UsfuiQYSBQOVVVXDdtOKfCzywnGyvaJr2tOCRrlCX2JT6NYZtu78Tc8VP
olSEcA2w4KKv79NW4hjyktbO1Cshki2IM7rMvzmKQDpSWpInXTBS8QO823wxQ7SM
1ABAHWKyAqoxH+phHzV0jMkjYv2RTkiDyWLrNnZcIbBJR/2XLL4ArDb76TvZoe5/
/6BHhn1/URTO317KV7g6M0vpfS0LodR0uAHfGfv/zb/myL6WgNYyJWbUMF1Zyu3Z
ycP5N2BZgQ7eU3nsO+rCD2VHIIwJPtLvJe7u+Yvdd8yE5UGR1H61H84tL0KLUB+G
m1ezk6q4XDNreJNRB0uzQhioyIhj/7qLo5XQe0J+S/cO77XgzhnlG5mSIFDuandH
MqQoo3VAJzyk1M6MxHAkLEuQZ9eBXj9rUMM4rwhGXV/njv+mjzyTWsIbbByBtGyQ
nBWuLmE5nCFYHXakqYouIzvstVHeGeWxn+m0lpd7g/m/v0jimHBBsQuTGYIqHj4Y
d2j+O6R8RtJo4HqLC5D8dVHyumRjlk6A07CBV+oTejz75IsBQFCvALya8LHXBZQ4
SF9Eu95MfIPAOKfTYfV+cea68oO3uKGrTmFJCk8X4tWBh2PKYT1oqhTpv3uFdK2u
wTUlFztrjPgt/u7K/uXzKqnBKtienWvralD7G4UGJYfYHwP/6qNKHSc3s8ugoKjn
+RQBIJqXLBj94p7zt6f+6JT2sbPnuAJb6pDNth8rxsmdvGZsWV3E4K8gPWg/K3TO
p78isz+hdVrasBeqvPoTUBCf1D0DLDNKZj7BZuGWRGugZmooUIDN+vM2fqbMOuL3
Uup40DffdRu267005kW0S9YK04TwqRlCDMGk4Ha8IerTA8UmVeJGTgRkGun9GfnT
r7B9dJYDBeW+QYPxoASauTDcvbQySpy7s8+wC4lFhmQtqWP/Hk7kbuXDIShV4LUV
S3KK6H8ZoecIcGtWAR4MNp4qbkwYEwumaADQ7ZJQ2j7wh2rZ4BhBEJwIyuzqVdG/
nY2n0xfXpyLJ9/Tw3yqhqoQd2s7UPRzObh9bfmOBicC6Gs6wTm4gWI5arwIUdJ60
zK9W68SY2Me5wUoLQHZpFkPSC2fwtFJerXJAhEwx58swBtjn1wkhIKtzHa8QIze5
YkceUtQMoMhYo8tW3aigXa90MxQAvcoH79N3QfNFYAJXxruzvnhkYB9ENAOXKKf0
32g6ospxmChQEOmXuvF4nJ2vnL1wEeFyovEPKhPIaM4WvjDJ8Frpgb36B4qSYpCv
9UBwPRbb/hAX8ZnZvTLGINto0LmZi2KGYFHqEckVIGTOq47T7E8QmRSI+Mib1RrO
hWoEyNr2DOWSizMC9bs4ZKANyl/y96fqnCJ6sbjt9QPEEiwabaeGOoqgPIgnat49
x+KqqaFgN4UAgqjl6KHwH9XiyvRMp3exAyc6xcXpH0CoWKMEHYp77guy/BHOKbj3
QUoh+uml5u45v+ALubHPKlIPhTVPR1L1FGylwNc/yFYumnzf6gEbNOfbqELu1NJs
pdsxwjAeCepwHgUQ9nlOt6s7uy3HjeOyWxlrEXQzJyoG8z1sljURjqFWD/Cuh5BW
DooBsTqvka4j9cS9nL/ubwrkGT4a5kPxMRphsYrTfjnqyynAyTrSxShKBk4uenkJ
strlP7C5pwA5gyI0s73+gRs4BtSf4hsouMn4nwzGbKKdyyTaZB65XWm2BXseECvI
jfp8vMqScZpq9nrwsEDDGg9y3SWPsBDHEM7Tz39zMmeA5gk5d5nB1Rhfl+b8FttB
wN080kjz8erhVianUyQLFZLOliYZq7BTmsechBwtM/B9HdGww7RoOS/m2mN2ubE3
V44mzAyJhmA3sSlYykFxqOApMoIjDCjNDkPgvDi3mRyHCfDZa6yc+qzpFMm8/nBY
ZMJtMdp0soVkGOgFzoHko72ZieaD4/UNftFxGToc4Nkd3+ibzca+wwxI/hQ7C/Cl
+bx6Ar4N7IRkqsJOoTv7F4rJBAwmXFf15EhW87+sp+jukGPKI0syOASX9Tlj2iRY
NVhiG0up+maOGDZ1k5RGT9jwwIBPgOcjAJN73YzCqzrWpqnPZkv8tOBO7juFU0Hx
Hnz+mJ/Ul4Q2gCapmUjf7X/mA0c33oZMVS+O+lBCQE0Ult8otAMzI4WnTlWaMEZp
o5ESA4O2YZ+xgkNY640SQorc1dSDq4qEeGu82X2GGJQIJ7Wj+8oNox/4unLOEPIV
JzsiREPm1IzUOwZCw+kKdl/2YQ+Q/NPH2IRe2thb/l56neKM5ZhG5vNmEVTgamOX
g9WtqoBzKsZQUJ8inEgWbQilMaUYKm065Hh2VUVQGT6k4GSR91iYpts2tGGRgHDD
JqpUEXDxLKqlOQfG/xfDpHFsYYJfrN7k1KS5V3mBDVkjrnO+Et/fTjU/urxJ1SyL
NOXOEMmjDEHvoeCUgyZlk6sMmogLdUJsY3lJgaxDnQz8Ddao8LHOhHR/oXcy7L9s
hJnpC51lCup6hlJMM1HRmylqDd947LPijjEeUhWnpDohaDzqVGcb3QjHzCMK+5Kr
oY1cQIgJPtL+yxDZHNDNjHvrlTRcMFQKYNaOEz3WFq2MMSAveQf0jMEecCURlTtZ
pyEUvkNFjnUTQnf1rWG/Qtf8upv1BcgT4zamzQTIpkC/jQo7kCJmEtavUericMK2
tv1GeIUkTfqiN4aIzmzXoEEsijNAdpmH0tDN/wN7PkKe00evil+NBoXsQz708pG3
FtZuZhNNBL2nuzjZ8Vk0l3QMmnz6OgeGMPLg0IXwePJkoVecyGdq3Q6K0epW0iV0
azFXzjCzoK6VxJeTY+OU6gjKr3ui4iX4gdAYbPUDycmvloepSVr+WibRBg5vgDqj
yQpC37Y6DKw6F/l1kl3DLlUQu0tCI5iofzmb60Tx8cbv3QQxPeoH3fgQq6zSrPCl
qpzzQmz1nIcL8badFFQ1Au8Ux4sreuGhPs2TNKN47AjEG5gQzIJqwDVnGUR3uVAe
xVzGN9bjgOQ2Gc3rx9y3Wcr23u7NCvUeq47b1SVrhENFx0OBHjE7uRutXsgpJhni
lqH+x2LcXH7lUj4eLFdAIrDAVGk+VUgNoWuoCgnDY5GXttCIjWGeU3wf+a+wAFSO
PcFel8PffPvYvjerBzD37QGUQ4HBCIC3I9Xb1hn/DUnUJtk4H5AGcELJO/HJg2s1
jbVP+yvonmVR05UM5vHcpy4GvuIsqY46w8VAlln5fzEskhYTlqBkvF7olJlGl/dF
BEEonMTLLSL4G7vsUovdvFzShjlo6tDcGr1SLUdmXanKnYetnRqdIqUr5p/0ke+C
fx3Khk7ocArzmIsYC5jYi2gPugYrm4kyE0FQH0vamoq9kONpa9aZcv3zoVVO4Fzx
gqY6Gh+K+2Nz9HyD5oPmiK4Zd8eVKaajUlqgEaeiJECvqZM0ZyZqcmU++mqrtcvz
y3JseVLmJkwciuRzQEa49ns4yUA9vSP50SAt2PbTRqS9HcXXbyoq/fvRAH8pYpYK
mRvsTMJ/I0V5SotcL3bntJS+0nlPyvUokYio9LaEglugxcykBnWDdWzxReSDiAz0
JmoDaYCnEhoZlYnXurx/4d6Rqx4ltl5rWCDW9AoXo67mIwdQ8pcSO8IXZZvFmgVa
tfpPoZduXYlzyNbizpdv5dq64Z3dARDYG4+qkA41dYnAbAMWusAUwNxWaMnGuGce
kX7+6r1vI2v/yv0+6U4pNww5Z2wfEy7Ik4tXvO2QshyaiASpPZeC9ofA8LmbTEIk
UVpD9+67/P53EvCvsslA2GzoMOB9Zu9AJ/skGvWd7x8xtn3x6PgW9XZ4/6Yyvc+m
8ceY+leWmkE1+ZdyWgdbjUyqTtZ5xdrVtwpq6Myrs5Ciea/zQ9zMFwsia8snz0kv
r0l7Be7ExfI84N26IAnHgHxRl+F/kFVRUjutc/5ygAK6jlHc5zbAOHuopMfYa3/B
9S0P0Ljmq2wQkRPy0jw1xhTtF2khugAEx5VWTp9guIdx7cofs0peB61IqQRJr8BX
riC6DP/43aJxpNqtLh5S8RaKF/e6Ea8aHASBvdL187aNFg/YyNCICN6pEXZZLBSW
IpLIUJQasxuI1YYcBYMn8lXNAM0oHbo+XPnofBkRRrUgBhs6kGDot0Z82CiuzkCF
LBQyuG5RIsNtj6AHi7jmweTCpV14xvh0tjVeSpgh2ATIb6jbYcjO6Ipc7e/q9dF5
XF/NYt3zQpX3yH9cJ/sU3VyrjFcXY2gKWhCEtGPl6QINu5GQNREGcOF+N0CNN7wN
a+W2kN/U3V44QbDthcVNDqFhBIITrFfB97K4RqclBoGfbja3x2Zs0OuLOUfEAOk8
nNx+5f3kdPmo99kiesmcDG141J/2sxTK9ijkHM5dw3joGhlGg78q1ly6T5GdBuIc
JvSLjALPSaET4HZWkVfUK+mnCbFNru42Cczd4rnA38TW+StgvwVfgb7c+vWHfSNg
KTzkWHOu13LUv17at5EMZGorLIPoRyM8JpM2wQyKvsPa2m+Tr/bPalSK3Og/fykQ
VPsKyOToVIdsQ0mUbx2NdDjfOhFkmzKABYIQPnHWvB0sUCsejf6YYM/1/HiSClL8
gPbtBM759e4KvU9VEd5qfJiZx0fiBaoBtJVu1p6J5EESnjWZVhob8xMdq94aj//4
htzKMyXfbHwPktacem4A/6/PBLBx434LEmvj0Pe6UcjElh4qE2LxxhHrlslhGlkn
gzMgF4/qaMWAk47BfH+xj7ReDGMZbZb4qe63KsQWPOAvdCMNY6hqHufHWIPm9rKv
4RV4F1p2ybqEC/zui5heoAUdzwFffF4/Pu51SX9PaHrUi9c3PA8c25j412lZOfeJ
0RO1S5rGUq6ZhD46XhGocGD6+5Ac88gqwtDdzPGGu4X1ieQExntd2EylLs9zctD0
aP3ABUSj1t1f6CJPlZnxJZuamO0ZuzeQbOB8lnEL1ptOc9Z6pcfkgymkVdpg9vDW
v5X09peUBjpn0LaQ9fOxag==
`pragma protect end_protected
