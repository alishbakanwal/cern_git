-- megafunction wizard: %Stratix V Transceiver Native PHY v16.0%
-- GENERATION: XML
-- alt_sv_gx_latopt_x3.vhd

-- Generated using ACDS version 16.0 211

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity alt_sv_gx_latopt_x3 is
	port (
		pll_powerdown           : in  std_logic_vector(0 downto 0)   := (others => '0'); --           pll_powerdown.pll_powerdown
		tx_analogreset          : in  std_logic_vector(2 downto 0)   := (others => '0'); --          tx_analogreset.tx_analogreset
		tx_digitalreset         : in  std_logic_vector(2 downto 0)   := (others => '0'); --         tx_digitalreset.tx_digitalreset
		tx_serial_data          : out std_logic_vector(2 downto 0);                      --          tx_serial_data.tx_serial_data
		ext_pll_clk             : in  std_logic_vector(2 downto 0)   := (others => '0'); --             ext_pll_clk.ext_pll_clk
		rx_analogreset          : in  std_logic_vector(2 downto 0)   := (others => '0'); --          rx_analogreset.rx_analogreset
		rx_digitalreset         : in  std_logic_vector(2 downto 0)   := (others => '0'); --         rx_digitalreset.rx_digitalreset
		rx_cdr_refclk           : in  std_logic_vector(0 downto 0)   := (others => '0'); --           rx_cdr_refclk.rx_cdr_refclk
		rx_serial_data          : in  std_logic_vector(2 downto 0)   := (others => '0'); --          rx_serial_data.rx_serial_data
		rx_clkslip              : in  std_logic_vector(2 downto 0)   := (others => '0'); --              rx_clkslip.rx_clkslip
		rx_is_lockedtoref       : out std_logic_vector(2 downto 0);                      --       rx_is_lockedtoref.rx_is_lockedtoref
		rx_is_lockedtodata      : out std_logic_vector(2 downto 0);                      --      rx_is_lockedtodata.rx_is_lockedtodata
		rx_seriallpbken         : in  std_logic_vector(2 downto 0)   := (others => '0'); --         rx_seriallpbken.rx_seriallpbken
		tx_std_coreclkin        : in  std_logic_vector(2 downto 0)   := (others => '0'); --        tx_std_coreclkin.tx_std_coreclkin
		rx_std_coreclkin        : in  std_logic_vector(2 downto 0)   := (others => '0'); --        rx_std_coreclkin.rx_std_coreclkin
		tx_std_clkout           : out std_logic_vector(2 downto 0);                      --           tx_std_clkout.tx_std_clkout
		rx_std_clkout           : out std_logic_vector(2 downto 0);                      --           rx_std_clkout.rx_std_clkout
		tx_std_polinv           : in  std_logic_vector(2 downto 0)   := (others => '0'); --           tx_std_polinv.tx_std_polinv
		rx_std_polinv           : in  std_logic_vector(2 downto 0)   := (others => '0'); --           rx_std_polinv.rx_std_polinv
		tx_cal_busy             : out std_logic_vector(2 downto 0);                      --             tx_cal_busy.tx_cal_busy
		rx_cal_busy             : out std_logic_vector(2 downto 0);                      --             rx_cal_busy.rx_cal_busy
		reconfig_to_xcvr        : in  std_logic_vector(209 downto 0) := (others => '0'); --        reconfig_to_xcvr.reconfig_to_xcvr
		reconfig_from_xcvr      : out std_logic_vector(137 downto 0);                    --      reconfig_from_xcvr.reconfig_from_xcvr
		tx_parallel_data        : in  std_logic_vector(119 downto 0) := (others => '0'); --        tx_parallel_data.tx_parallel_data
		unused_tx_parallel_data : in  std_logic_vector(71 downto 0)  := (others => '0'); -- unused_tx_parallel_data.unused_tx_parallel_data
		rx_parallel_data        : out std_logic_vector(119 downto 0);                    --        rx_parallel_data.rx_parallel_data
		unused_rx_parallel_data : out std_logic_vector(71 downto 0)                      -- unused_rx_parallel_data.unused_rx_parallel_data
	);
end entity alt_sv_gx_latopt_x3;

architecture rtl of alt_sv_gx_latopt_x3 is
	component altera_xcvr_native_sv is
		generic (
			tx_enable                       : integer := 1;
			rx_enable                       : integer := 1;
			enable_std                      : integer := 0;
			enable_teng                     : integer := 0;
			data_path_select                : string  := "pma_direct";
			channels                        : integer := 1;
			bonded_mode                     : string  := "non_bonded";
			data_rate                       : string  := "";
			pma_width                       : integer := 80;
			tx_pma_clk_div                  : integer := 1;
			tx_pma_txdetectrx_ctrl          : integer := 0;
			pll_reconfig_enable             : integer := 0;
			pll_external_enable             : integer := 0;
			pll_data_rate                   : string  := "0 Mbps";
			pll_type                        : string  := "CMU";
			pll_network_select              : string  := "x1";
			plls                            : integer := 1;
			pll_select                      : integer := 0;
			pll_refclk_cnt                  : integer := 1;
			pll_refclk_select               : string  := "0";
			pll_refclk_freq                 : string  := "125.0 MHz";
			pll_feedback_path               : string  := "internal";
			cdr_reconfig_enable             : integer := 0;
			cdr_refclk_cnt                  : integer := 1;
			cdr_refclk_select               : integer := 0;
			cdr_refclk_freq                 : string  := "";
			rx_ppm_detect_threshold         : string  := "1000";
			rx_clkslip_enable               : integer := 0;
			std_protocol_hint               : string  := "basic";
			std_pcs_pma_width               : integer := 10;
			std_low_latency_bypass_enable   : integer := 0;
			std_tx_pcfifo_mode              : string  := "low_latency";
			std_rx_pcfifo_mode              : string  := "low_latency";
			std_rx_byte_order_enable        : integer := 0;
			std_rx_byte_order_mode          : string  := "manual";
			std_rx_byte_order_width         : integer := 10;
			std_rx_byte_order_symbol_count  : integer := 1;
			std_rx_byte_order_pattern       : string  := "0";
			std_rx_byte_order_pad           : string  := "0";
			std_tx_byte_ser_enable          : integer := 0;
			std_rx_byte_deser_enable        : integer := 0;
			std_tx_8b10b_enable             : integer := 0;
			std_tx_8b10b_disp_ctrl_enable   : integer := 0;
			std_rx_8b10b_enable             : integer := 0;
			std_rx_rmfifo_enable            : integer := 0;
			std_rx_rmfifo_pattern_p         : string  := "00000";
			std_rx_rmfifo_pattern_n         : string  := "00000";
			std_tx_bitslip_enable           : integer := 0;
			std_rx_word_aligner_mode        : string  := "bit_slip";
			std_rx_word_aligner_pattern_len : integer := 7;
			std_rx_word_aligner_pattern     : string  := "0000000000";
			std_rx_word_aligner_rknumber    : integer := 3;
			std_rx_word_aligner_renumber    : integer := 3;
			std_rx_word_aligner_rgnumber    : integer := 3;
			std_rx_run_length_val           : integer := 31;
			std_tx_bitrev_enable            : integer := 0;
			std_rx_bitrev_enable            : integer := 0;
			std_tx_byterev_enable           : integer := 0;
			std_rx_byterev_enable           : integer := 0;
			std_tx_polinv_enable            : integer := 0;
			std_rx_polinv_enable            : integer := 0;
			teng_protocol_hint              : string  := "basic";
			teng_pcs_pma_width              : integer := 40;
			teng_pld_pcs_width              : integer := 40;
			teng_txfifo_mode                : string  := "phase_comp";
			teng_txfifo_full                : integer := 31;
			teng_txfifo_empty               : integer := 0;
			teng_txfifo_pfull               : integer := 23;
			teng_txfifo_pempty              : integer := 2;
			teng_rxfifo_mode                : string  := "phase_comp";
			teng_rxfifo_full                : integer := 31;
			teng_rxfifo_empty               : integer := 0;
			teng_rxfifo_pfull               : integer := 23;
			teng_rxfifo_pempty              : integer := 2;
			teng_rxfifo_align_del           : integer := 0;
			teng_rxfifo_control_del         : integer := 0;
			teng_tx_frmgen_enable           : integer := 0;
			teng_tx_frmgen_user_length      : integer := 2048;
			teng_tx_frmgen_burst_enable     : integer := 0;
			teng_rx_frmsync_enable          : integer := 0;
			teng_rx_frmsync_user_length     : integer := 2048;
			teng_frmgensync_diag_word       : string  := "6400000000000000";
			teng_frmgensync_scrm_word       : string  := "2800000000000000";
			teng_frmgensync_skip_word       : string  := "1e1e1e1e1e1e1e1e";
			teng_frmgensync_sync_word       : string  := "78f678f678f678f6";
			teng_tx_sh_err                  : integer := 0;
			teng_tx_crcgen_enable           : integer := 0;
			teng_rx_crcchk_enable           : integer := 0;
			teng_tx_64b66b_enable           : integer := 0;
			teng_rx_64b66b_enable           : integer := 0;
			teng_tx_scram_enable            : integer := 0;
			teng_tx_scram_user_seed         : string  := "000000000000000";
			teng_rx_descram_enable          : integer := 0;
			teng_tx_dispgen_enable          : integer := 0;
			teng_rx_dispchk_enable          : integer := 0;
			teng_rx_blksync_enable          : integer := 0;
			teng_tx_polinv_enable           : integer := 0;
			teng_tx_bitslip_enable          : integer := 0;
			teng_rx_polinv_enable           : integer := 0;
			teng_rx_bitslip_enable          : integer := 0
		);
		port (
			pll_powerdown             : in  std_logic_vector(0 downto 0)   := (others => 'X'); -- pll_powerdown
			tx_analogreset            : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- tx_analogreset
			tx_digitalreset           : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- tx_digitalreset
			tx_serial_data            : out std_logic_vector(2 downto 0);                      -- tx_serial_data
			ext_pll_clk               : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- ext_pll_clk
			rx_analogreset            : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- rx_analogreset
			rx_digitalreset           : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- rx_digitalreset
			rx_cdr_refclk             : in  std_logic_vector(0 downto 0)   := (others => 'X'); -- rx_cdr_refclk
			rx_serial_data            : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- rx_serial_data
			rx_clkslip                : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- rx_clkslip
			rx_is_lockedtoref         : out std_logic_vector(2 downto 0);                      -- rx_is_lockedtoref
			rx_is_lockedtodata        : out std_logic_vector(2 downto 0);                      -- rx_is_lockedtodata
			rx_seriallpbken           : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- rx_seriallpbken
			tx_std_coreclkin          : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- tx_std_coreclkin
			rx_std_coreclkin          : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- rx_std_coreclkin
			tx_std_clkout             : out std_logic_vector(2 downto 0);                      -- tx_std_clkout
			rx_std_clkout             : out std_logic_vector(2 downto 0);                      -- rx_std_clkout
			tx_std_polinv             : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- tx_std_polinv
			rx_std_polinv             : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- rx_std_polinv
			tx_cal_busy               : out std_logic_vector(2 downto 0);                      -- tx_cal_busy
			rx_cal_busy               : out std_logic_vector(2 downto 0);                      -- rx_cal_busy
			reconfig_to_xcvr          : in  std_logic_vector(209 downto 0) := (others => 'X'); -- reconfig_to_xcvr
			reconfig_from_xcvr        : out std_logic_vector(137 downto 0);                    -- reconfig_from_xcvr
			tx_parallel_data          : in  std_logic_vector(191 downto 0) := (others => 'X'); -- unused_tx_parallel_data
			rx_parallel_data          : out std_logic_vector(191 downto 0);                    -- unused_rx_parallel_data
			tx_pll_refclk             : in  std_logic_vector(0 downto 0)   := (others => 'X'); -- tx_pll_refclk
			tx_pma_clkout             : out std_logic_vector(2 downto 0);                      -- tx_pma_clkout
			tx_pma_pclk               : out std_logic_vector(2 downto 0);                      -- tx_pma_pclk
			tx_pma_parallel_data      : in  std_logic_vector(239 downto 0) := (others => 'X'); -- tx_pma_parallel_data
			pll_locked                : out std_logic_vector(0 downto 0);                      -- pll_locked
			rx_pma_clkout             : out std_logic_vector(2 downto 0);                      -- rx_pma_clkout
			rx_pma_pclk               : out std_logic_vector(2 downto 0);                      -- rx_pma_pclk
			rx_pma_parallel_data      : out std_logic_vector(239 downto 0);                    -- rx_pma_parallel_data
			rx_clklow                 : out std_logic_vector(2 downto 0);                      -- rx_clklow
			rx_fref                   : out std_logic_vector(2 downto 0);                      -- rx_fref
			rx_set_locktodata         : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- rx_set_locktodata
			rx_set_locktoref          : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- rx_set_locktoref
			rx_signaldetect           : out std_logic_vector(2 downto 0);                      -- rx_signaldetect
			rx_pma_qpipulldn          : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- rx_pma_qpipulldn
			tx_pma_qpipullup          : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- tx_pma_qpipullup
			tx_pma_qpipulldn          : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- tx_pma_qpipulldn
			tx_pma_txdetectrx         : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- tx_pma_txdetectrx
			tx_pma_rxfound            : out std_logic_vector(2 downto 0);                      -- tx_pma_rxfound
			rx_std_prbs_done          : out std_logic_vector(2 downto 0);                      -- rx_std_prbs_done
			rx_std_prbs_err           : out std_logic_vector(2 downto 0);                      -- rx_std_prbs_err
			tx_std_pcfifo_full        : out std_logic_vector(2 downto 0);                      -- tx_std_pcfifo_full
			tx_std_pcfifo_empty       : out std_logic_vector(2 downto 0);                      -- tx_std_pcfifo_empty
			rx_std_pcfifo_full        : out std_logic_vector(2 downto 0);                      -- rx_std_pcfifo_full
			rx_std_pcfifo_empty       : out std_logic_vector(2 downto 0);                      -- rx_std_pcfifo_empty
			rx_std_byteorder_ena      : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- rx_std_byteorder_ena
			rx_std_byteorder_flag     : out std_logic_vector(2 downto 0);                      -- rx_std_byteorder_flag
			rx_std_rmfifo_full        : out std_logic_vector(2 downto 0);                      -- rx_std_rmfifo_full
			rx_std_rmfifo_empty       : out std_logic_vector(2 downto 0);                      -- rx_std_rmfifo_empty
			rx_std_wa_patternalign    : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- rx_std_wa_patternalign
			rx_std_wa_a1a2size        : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- rx_std_wa_a1a2size
			tx_std_bitslipboundarysel : in  std_logic_vector(14 downto 0)  := (others => 'X'); -- tx_std_bitslipboundarysel
			rx_std_bitslipboundarysel : out std_logic_vector(14 downto 0);                     -- rx_std_bitslipboundarysel
			rx_std_bitslip            : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- rx_std_bitslip
			rx_std_runlength_err      : out std_logic_vector(2 downto 0);                      -- rx_std_runlength_err
			rx_std_bitrev_ena         : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- rx_std_bitrev_ena
			rx_std_byterev_ena        : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- rx_std_byterev_ena
			tx_std_elecidle           : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- tx_std_elecidle
			rx_std_signaldetect       : out std_logic_vector(2 downto 0);                      -- rx_std_signaldetect
			tx_10g_coreclkin          : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- tx_10g_coreclkin
			rx_10g_coreclkin          : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- rx_10g_coreclkin
			tx_10g_clkout             : out std_logic_vector(2 downto 0);                      -- tx_10g_clkout
			rx_10g_clkout             : out std_logic_vector(2 downto 0);                      -- rx_10g_clkout
			rx_10g_clk33out           : out std_logic_vector(2 downto 0);                      -- rx_10g_clk33out
			rx_10g_prbs_err_clr       : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- rx_10g_prbs_err_clr
			rx_10g_prbs_done          : out std_logic_vector(2 downto 0);                      -- rx_10g_prbs_done
			rx_10g_prbs_err           : out std_logic_vector(2 downto 0);                      -- rx_10g_prbs_err
			tx_10g_control            : in  std_logic_vector(26 downto 0)  := (others => 'X'); -- tx_10g_control
			rx_10g_control            : out std_logic_vector(29 downto 0);                     -- rx_10g_control
			tx_10g_data_valid         : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- tx_10g_data_valid
			tx_10g_fifo_full          : out std_logic_vector(2 downto 0);                      -- tx_10g_fifo_full
			tx_10g_fifo_pfull         : out std_logic_vector(2 downto 0);                      -- tx_10g_fifo_pfull
			tx_10g_fifo_empty         : out std_logic_vector(2 downto 0);                      -- tx_10g_fifo_empty
			tx_10g_fifo_pempty        : out std_logic_vector(2 downto 0);                      -- tx_10g_fifo_pempty
			tx_10g_fifo_del           : out std_logic_vector(2 downto 0);                      -- tx_10g_fifo_del
			tx_10g_fifo_insert        : out std_logic_vector(2 downto 0);                      -- tx_10g_fifo_insert
			rx_10g_fifo_rd_en         : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- rx_10g_fifo_rd_en
			rx_10g_data_valid         : out std_logic_vector(2 downto 0);                      -- rx_10g_data_valid
			rx_10g_fifo_full          : out std_logic_vector(2 downto 0);                      -- rx_10g_fifo_full
			rx_10g_fifo_pfull         : out std_logic_vector(2 downto 0);                      -- rx_10g_fifo_pfull
			rx_10g_fifo_empty         : out std_logic_vector(2 downto 0);                      -- rx_10g_fifo_empty
			rx_10g_fifo_pempty        : out std_logic_vector(2 downto 0);                      -- rx_10g_fifo_pempty
			rx_10g_fifo_del           : out std_logic_vector(2 downto 0);                      -- rx_10g_fifo_del
			rx_10g_fifo_insert        : out std_logic_vector(2 downto 0);                      -- rx_10g_fifo_insert
			rx_10g_fifo_align_val     : out std_logic_vector(2 downto 0);                      -- rx_10g_fifo_align_val
			rx_10g_fifo_align_clr     : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- rx_10g_fifo_align_clr
			rx_10g_fifo_align_en      : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- rx_10g_fifo_align_en
			tx_10g_frame              : out std_logic_vector(2 downto 0);                      -- tx_10g_frame
			tx_10g_frame_diag_status  : in  std_logic_vector(5 downto 0)   := (others => 'X'); -- tx_10g_frame_diag_status
			tx_10g_frame_burst_en     : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- tx_10g_frame_burst_en
			rx_10g_frame              : out std_logic_vector(2 downto 0);                      -- rx_10g_frame
			rx_10g_frame_lock         : out std_logic_vector(2 downto 0);                      -- rx_10g_frame_lock
			rx_10g_frame_mfrm_err     : out std_logic_vector(2 downto 0);                      -- rx_10g_frame_mfrm_err
			rx_10g_frame_sync_err     : out std_logic_vector(2 downto 0);                      -- rx_10g_frame_sync_err
			rx_10g_frame_skip_ins     : out std_logic_vector(2 downto 0);                      -- rx_10g_frame_skip_ins
			rx_10g_frame_pyld_ins     : out std_logic_vector(2 downto 0);                      -- rx_10g_frame_pyld_ins
			rx_10g_frame_skip_err     : out std_logic_vector(2 downto 0);                      -- rx_10g_frame_skip_err
			rx_10g_frame_diag_err     : out std_logic_vector(2 downto 0);                      -- rx_10g_frame_diag_err
			rx_10g_frame_diag_status  : out std_logic_vector(5 downto 0);                      -- rx_10g_frame_diag_status
			rx_10g_crc32_err          : out std_logic_vector(2 downto 0);                      -- rx_10g_crc32err
			rx_10g_descram_err        : out std_logic_vector(2 downto 0);                      -- rx_10g_descram_err
			rx_10g_blk_lock           : out std_logic_vector(2 downto 0);                      -- rx_10g_blk_lock
			rx_10g_blk_sh_err         : out std_logic_vector(2 downto 0);                      -- rx_10g_blk_sh_err
			tx_10g_bitslip            : in  std_logic_vector(20 downto 0)  := (others => 'X'); -- tx_10g_bitslip
			rx_10g_bitslip            : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- rx_10g_bitslip
			rx_10g_highber            : out std_logic_vector(2 downto 0);                      -- rx_10g_highber
			rx_10g_highber_clr_cnt    : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- rx_10g_highber_clr_cnt
			rx_10g_clr_errblk_count   : in  std_logic_vector(2 downto 0)   := (others => 'X')  -- rx_10g_clr_errblk_count
		);
	end component altera_xcvr_native_sv;

	signal alt_sv_gx_latopt_x3_inst_rx_parallel_data : std_logic_vector(191 downto 0); -- port fragment

begin

	alt_sv_gx_latopt_x3_inst : component altera_xcvr_native_sv
		generic map (
			tx_enable                       => 1,
			rx_enable                       => 1,
			enable_std                      => 1,
			enable_teng                     => 0,
			data_path_select                => "standard",
			channels                        => 3,
			bonded_mode                     => "xN",
			data_rate                       => "4800 Mbps",
			pma_width                       => 20,
			tx_pma_clk_div                  => 1,
			tx_pma_txdetectrx_ctrl          => 0,
			pll_reconfig_enable             => 0,
			pll_external_enable             => 1,
			pll_data_rate                   => "4800 Mbps",
			pll_type                        => "CMU",
			pll_network_select              => "x1",
			plls                            => 1,
			pll_select                      => 0,
			pll_refclk_cnt                  => 1,
			pll_refclk_select               => "0",
			pll_refclk_freq                 => "240.0 MHz",
			pll_feedback_path               => "internal",
			cdr_reconfig_enable             => 0,
			cdr_refclk_cnt                  => 1,
			cdr_refclk_select               => 0,
			cdr_refclk_freq                 => "120.0 MHz",
			rx_ppm_detect_threshold         => "1000",
			rx_clkslip_enable               => 1,
			std_protocol_hint               => "basic",
			std_pcs_pma_width               => 20,
			std_low_latency_bypass_enable   => 1,
			std_tx_pcfifo_mode              => "register_fifo",
			std_rx_pcfifo_mode              => "register_fifo",
			std_rx_byte_order_enable        => 0,
			std_rx_byte_order_mode          => "manual",
			std_rx_byte_order_width         => 10,
			std_rx_byte_order_symbol_count  => 1,
			std_rx_byte_order_pattern       => "0",
			std_rx_byte_order_pad           => "0",
			std_tx_byte_ser_enable          => 1,
			std_rx_byte_deser_enable        => 1,
			std_tx_8b10b_enable             => 0,
			std_tx_8b10b_disp_ctrl_enable   => 0,
			std_rx_8b10b_enable             => 0,
			std_rx_rmfifo_enable            => 0,
			std_rx_rmfifo_pattern_p         => "00000",
			std_rx_rmfifo_pattern_n         => "00000",
			std_tx_bitslip_enable           => 0,
			std_rx_word_aligner_mode        => "bit_slip",
			std_rx_word_aligner_pattern_len => 7,
			std_rx_word_aligner_pattern     => "0000000000",
			std_rx_word_aligner_rknumber    => 3,
			std_rx_word_aligner_renumber    => 3,
			std_rx_word_aligner_rgnumber    => 3,
			std_rx_run_length_val           => 31,
			std_tx_bitrev_enable            => 0,
			std_rx_bitrev_enable            => 0,
			std_tx_byterev_enable           => 0,
			std_rx_byterev_enable           => 0,
			std_tx_polinv_enable            => 1,
			std_rx_polinv_enable            => 1,
			teng_protocol_hint              => "basic",
			teng_pcs_pma_width              => 40,
			teng_pld_pcs_width              => 40,
			teng_txfifo_mode                => "phase_comp",
			teng_txfifo_full                => 31,
			teng_txfifo_empty               => 0,
			teng_txfifo_pfull               => 23,
			teng_txfifo_pempty              => 2,
			teng_rxfifo_mode                => "phase_comp",
			teng_rxfifo_full                => 31,
			teng_rxfifo_empty               => 0,
			teng_rxfifo_pfull               => 23,
			teng_rxfifo_pempty              => 2,
			teng_rxfifo_align_del           => 0,
			teng_rxfifo_control_del         => 0,
			teng_tx_frmgen_enable           => 0,
			teng_tx_frmgen_user_length      => 2048,
			teng_tx_frmgen_burst_enable     => 0,
			teng_rx_frmsync_enable          => 0,
			teng_rx_frmsync_user_length     => 2048,
			teng_frmgensync_diag_word       => "6400000000000000",
			teng_frmgensync_scrm_word       => "2800000000000000",
			teng_frmgensync_skip_word       => "1e1e1e1e1e1e1e1e",
			teng_frmgensync_sync_word       => "78f678f678f678f6",
			teng_tx_sh_err                  => 0,
			teng_tx_crcgen_enable           => 0,
			teng_rx_crcchk_enable           => 0,
			teng_tx_64b66b_enable           => 0,
			teng_rx_64b66b_enable           => 0,
			teng_tx_scram_enable            => 0,
			teng_tx_scram_user_seed         => "000000000000000",
			teng_rx_descram_enable          => 0,
			teng_tx_dispgen_enable          => 0,
			teng_rx_dispchk_enable          => 0,
			teng_rx_blksync_enable          => 0,
			teng_tx_polinv_enable           => 0,
			teng_tx_bitslip_enable          => 0,
			teng_rx_polinv_enable           => 0,
			teng_rx_bitslip_enable          => 0
		)
		port map (
			pll_powerdown             => pll_powerdown,                                                                                                                                                                                                                                      --      pll_powerdown.pll_powerdown
			tx_analogreset            => tx_analogreset,                                                                                                                                                                                                                                     --     tx_analogreset.tx_analogreset
			tx_digitalreset           => tx_digitalreset,                                                                                                                                                                                                                                    --    tx_digitalreset.tx_digitalreset
			tx_serial_data            => tx_serial_data,                                                                                                                                                                                                                                     --     tx_serial_data.tx_serial_data
			ext_pll_clk               => ext_pll_clk,                                                                                                                                                                                                                                        --        ext_pll_clk.ext_pll_clk
			rx_analogreset            => rx_analogreset,                                                                                                                                                                                                                                     --     rx_analogreset.rx_analogreset
			rx_digitalreset           => rx_digitalreset,                                                                                                                                                                                                                                    --    rx_digitalreset.rx_digitalreset
			rx_cdr_refclk             => rx_cdr_refclk,                                                                                                                                                                                                                                      --      rx_cdr_refclk.rx_cdr_refclk
			rx_serial_data            => rx_serial_data,                                                                                                                                                                                                                                     --     rx_serial_data.rx_serial_data
			rx_clkslip                => rx_clkslip,                                                                                                                                                                                                                                         --         rx_clkslip.rx_clkslip
			rx_is_lockedtoref         => rx_is_lockedtoref,                                                                                                                                                                                                                                  --  rx_is_lockedtoref.rx_is_lockedtoref
			rx_is_lockedtodata        => rx_is_lockedtodata,                                                                                                                                                                                                                                 -- rx_is_lockedtodata.rx_is_lockedtodata
			rx_seriallpbken           => rx_seriallpbken,                                                                                                                                                                                                                                    --    rx_seriallpbken.rx_seriallpbken
			tx_std_coreclkin          => tx_std_coreclkin,                                                                                                                                                                                                                                   --   tx_std_coreclkin.tx_std_coreclkin
			rx_std_coreclkin          => rx_std_coreclkin,                                                                                                                                                                                                                                   --   rx_std_coreclkin.rx_std_coreclkin
			tx_std_clkout             => tx_std_clkout,                                                                                                                                                                                                                                      --      tx_std_clkout.tx_std_clkout
			rx_std_clkout             => rx_std_clkout,                                                                                                                                                                                                                                      --      rx_std_clkout.rx_std_clkout
			tx_std_polinv             => tx_std_polinv,                                                                                                                                                                                                                                      --      tx_std_polinv.tx_std_polinv
			rx_std_polinv             => rx_std_polinv,                                                                                                                                                                                                                                      --      rx_std_polinv.rx_std_polinv
			tx_cal_busy               => tx_cal_busy,                                                                                                                                                                                                                                        --        tx_cal_busy.tx_cal_busy
			rx_cal_busy               => rx_cal_busy,                                                                                                                                                                                                                                        --        rx_cal_busy.rx_cal_busy
			reconfig_to_xcvr          => reconfig_to_xcvr,                                                                                                                                                                                                                                   --   reconfig_to_xcvr.reconfig_to_xcvr
			reconfig_from_xcvr        => reconfig_from_xcvr,                                                                                                                                                                                                                                 -- reconfig_from_xcvr.reconfig_from_xcvr
			tx_parallel_data(0)       => tx_parallel_data(0),                                                                                                                                                                                                                                --   tx_parallel_data.tx_parallel_data
			tx_parallel_data(1)       => tx_parallel_data(1),                                                                                                                                                                                                                                --                   .tx_parallel_data
			tx_parallel_data(2)       => tx_parallel_data(2),                                                                                                                                                                                                                                --                   .tx_parallel_data
			tx_parallel_data(3)       => tx_parallel_data(3),                                                                                                                                                                                                                                --                   .tx_parallel_data
			tx_parallel_data(4)       => tx_parallel_data(4),                                                                                                                                                                                                                                --                   .tx_parallel_data
			tx_parallel_data(5)       => tx_parallel_data(5),                                                                                                                                                                                                                                --                   .tx_parallel_data
			tx_parallel_data(6)       => tx_parallel_data(6),                                                                                                                                                                                                                                --                   .tx_parallel_data
			tx_parallel_data(7)       => tx_parallel_data(7),                                                                                                                                                                                                                                --                   .tx_parallel_data
			tx_parallel_data(8)       => tx_parallel_data(8),                                                                                                                                                                                                                                --                   .tx_parallel_data
			tx_parallel_data(9)       => tx_parallel_data(9),                                                                                                                                                                                                                                --                   .tx_parallel_data
			tx_parallel_data(10)      => unused_tx_parallel_data(0),                                                                                                                                                                                                                         --                   .tx_parallel_data
			tx_parallel_data(11)      => tx_parallel_data(10),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(12)      => tx_parallel_data(11),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(13)      => tx_parallel_data(12),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(14)      => tx_parallel_data(13),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(15)      => tx_parallel_data(14),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(16)      => tx_parallel_data(15),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(17)      => tx_parallel_data(16),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(18)      => tx_parallel_data(17),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(19)      => tx_parallel_data(18),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(20)      => tx_parallel_data(19),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(21)      => unused_tx_parallel_data(1),                                                                                                                                                                                                                         --                   .tx_parallel_data
			tx_parallel_data(22)      => tx_parallel_data(20),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(23)      => tx_parallel_data(21),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(24)      => tx_parallel_data(22),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(25)      => tx_parallel_data(23),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(26)      => tx_parallel_data(24),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(27)      => tx_parallel_data(25),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(28)      => tx_parallel_data(26),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(29)      => tx_parallel_data(27),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(30)      => tx_parallel_data(28),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(31)      => tx_parallel_data(29),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(32)      => unused_tx_parallel_data(2),                                                                                                                                                                                                                         --                   .tx_parallel_data
			tx_parallel_data(33)      => tx_parallel_data(30),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(34)      => tx_parallel_data(31),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(35)      => tx_parallel_data(32),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(36)      => tx_parallel_data(33),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(37)      => tx_parallel_data(34),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(38)      => tx_parallel_data(35),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(39)      => tx_parallel_data(36),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(40)      => tx_parallel_data(37),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(41)      => tx_parallel_data(38),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(42)      => tx_parallel_data(39),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(43)      => unused_tx_parallel_data(3),                                                                                                                                                                                                                         --                   .tx_parallel_data
			tx_parallel_data(44)      => unused_tx_parallel_data(4),                                                                                                                                                                                                                         --                   .tx_parallel_data
			tx_parallel_data(45)      => unused_tx_parallel_data(5),                                                                                                                                                                                                                         --                   .tx_parallel_data
			tx_parallel_data(46)      => unused_tx_parallel_data(6),                                                                                                                                                                                                                         --                   .tx_parallel_data
			tx_parallel_data(47)      => unused_tx_parallel_data(7),                                                                                                                                                                                                                         --                   .tx_parallel_data
			tx_parallel_data(48)      => unused_tx_parallel_data(8),                                                                                                                                                                                                                         --                   .tx_parallel_data
			tx_parallel_data(49)      => unused_tx_parallel_data(9),                                                                                                                                                                                                                         --                   .tx_parallel_data
			tx_parallel_data(50)      => unused_tx_parallel_data(10),                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(51)      => unused_tx_parallel_data(11),                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(52)      => unused_tx_parallel_data(12),                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(53)      => unused_tx_parallel_data(13),                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(54)      => unused_tx_parallel_data(14),                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(55)      => unused_tx_parallel_data(15),                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(56)      => unused_tx_parallel_data(16),                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(57)      => unused_tx_parallel_data(17),                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(58)      => unused_tx_parallel_data(18),                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(59)      => unused_tx_parallel_data(19),                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(60)      => unused_tx_parallel_data(20),                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(61)      => unused_tx_parallel_data(21),                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(62)      => unused_tx_parallel_data(22),                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(63)      => unused_tx_parallel_data(23),                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(64)      => tx_parallel_data(40),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(65)      => tx_parallel_data(41),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(66)      => tx_parallel_data(42),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(67)      => tx_parallel_data(43),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(68)      => tx_parallel_data(44),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(69)      => tx_parallel_data(45),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(70)      => tx_parallel_data(46),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(71)      => tx_parallel_data(47),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(72)      => tx_parallel_data(48),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(73)      => tx_parallel_data(49),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(74)      => unused_tx_parallel_data(24),                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(75)      => tx_parallel_data(50),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(76)      => tx_parallel_data(51),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(77)      => tx_parallel_data(52),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(78)      => tx_parallel_data(53),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(79)      => tx_parallel_data(54),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(80)      => tx_parallel_data(55),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(81)      => tx_parallel_data(56),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(82)      => tx_parallel_data(57),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(83)      => tx_parallel_data(58),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(84)      => tx_parallel_data(59),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(85)      => unused_tx_parallel_data(25),                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(86)      => tx_parallel_data(60),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(87)      => tx_parallel_data(61),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(88)      => tx_parallel_data(62),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(89)      => tx_parallel_data(63),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(90)      => tx_parallel_data(64),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(91)      => tx_parallel_data(65),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(92)      => tx_parallel_data(66),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(93)      => tx_parallel_data(67),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(94)      => tx_parallel_data(68),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(95)      => tx_parallel_data(69),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(96)      => unused_tx_parallel_data(26),                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(97)      => tx_parallel_data(70),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(98)      => tx_parallel_data(71),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(99)      => tx_parallel_data(72),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(100)     => tx_parallel_data(73),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(101)     => tx_parallel_data(74),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(102)     => tx_parallel_data(75),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(103)     => tx_parallel_data(76),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(104)     => tx_parallel_data(77),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(105)     => tx_parallel_data(78),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(106)     => tx_parallel_data(79),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(107)     => unused_tx_parallel_data(27),                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(108)     => unused_tx_parallel_data(28),                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(109)     => unused_tx_parallel_data(29),                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(110)     => unused_tx_parallel_data(30),                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(111)     => unused_tx_parallel_data(31),                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(112)     => unused_tx_parallel_data(32),                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(113)     => unused_tx_parallel_data(33),                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(114)     => unused_tx_parallel_data(34),                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(115)     => unused_tx_parallel_data(35),                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(116)     => unused_tx_parallel_data(36),                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(117)     => unused_tx_parallel_data(37),                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(118)     => unused_tx_parallel_data(38),                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(119)     => unused_tx_parallel_data(39),                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(120)     => unused_tx_parallel_data(40),                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(121)     => unused_tx_parallel_data(41),                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(122)     => unused_tx_parallel_data(42),                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(123)     => unused_tx_parallel_data(43),                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(124)     => unused_tx_parallel_data(44),                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(125)     => unused_tx_parallel_data(45),                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(126)     => unused_tx_parallel_data(46),                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(127)     => unused_tx_parallel_data(47),                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(128)     => tx_parallel_data(80),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(129)     => tx_parallel_data(81),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(130)     => tx_parallel_data(82),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(131)     => tx_parallel_data(83),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(132)     => tx_parallel_data(84),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(133)     => tx_parallel_data(85),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(134)     => tx_parallel_data(86),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(135)     => tx_parallel_data(87),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(136)     => tx_parallel_data(88),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(137)     => tx_parallel_data(89),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(138)     => unused_tx_parallel_data(48),                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(139)     => tx_parallel_data(90),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(140)     => tx_parallel_data(91),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(141)     => tx_parallel_data(92),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(142)     => tx_parallel_data(93),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(143)     => tx_parallel_data(94),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(144)     => tx_parallel_data(95),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(145)     => tx_parallel_data(96),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(146)     => tx_parallel_data(97),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(147)     => tx_parallel_data(98),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(148)     => tx_parallel_data(99),                                                                                                                                                                                                                               --                   .tx_parallel_data
			tx_parallel_data(149)     => unused_tx_parallel_data(49),                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(150)     => tx_parallel_data(100),                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(151)     => tx_parallel_data(101),                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(152)     => tx_parallel_data(102),                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(153)     => tx_parallel_data(103),                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(154)     => tx_parallel_data(104),                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(155)     => tx_parallel_data(105),                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(156)     => tx_parallel_data(106),                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(157)     => tx_parallel_data(107),                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(158)     => tx_parallel_data(108),                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(159)     => tx_parallel_data(109),                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(160)     => unused_tx_parallel_data(50),                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(161)     => tx_parallel_data(110),                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(162)     => tx_parallel_data(111),                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(163)     => tx_parallel_data(112),                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(164)     => tx_parallel_data(113),                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(165)     => tx_parallel_data(114),                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(166)     => tx_parallel_data(115),                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(167)     => tx_parallel_data(116),                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(168)     => tx_parallel_data(117),                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(169)     => tx_parallel_data(118),                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(170)     => tx_parallel_data(119),                                                                                                                                                                                                                              --                   .tx_parallel_data
			tx_parallel_data(171)     => unused_tx_parallel_data(51),                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(172)     => unused_tx_parallel_data(52),                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(173)     => unused_tx_parallel_data(53),                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(174)     => unused_tx_parallel_data(54),                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(175)     => unused_tx_parallel_data(55),                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(176)     => unused_tx_parallel_data(56),                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(177)     => unused_tx_parallel_data(57),                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(178)     => unused_tx_parallel_data(58),                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(179)     => unused_tx_parallel_data(59),                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(180)     => unused_tx_parallel_data(60),                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(181)     => unused_tx_parallel_data(61),                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(182)     => unused_tx_parallel_data(62),                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(183)     => unused_tx_parallel_data(63),                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(184)     => unused_tx_parallel_data(64),                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(185)     => unused_tx_parallel_data(65),                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(186)     => unused_tx_parallel_data(66),                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(187)     => unused_tx_parallel_data(67),                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(188)     => unused_tx_parallel_data(68),                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(189)     => unused_tx_parallel_data(69),                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(190)     => unused_tx_parallel_data(70),                                                                                                                                                                                                                        --                   .tx_parallel_data
			tx_parallel_data(191)     => unused_tx_parallel_data(71),                                                                                                                                                                                                                        --                   .tx_parallel_data
			rx_parallel_data(0)       => alt_sv_gx_latopt_x3_inst_rx_parallel_data(0),                                                                                                                                                                                                       --   rx_parallel_data.rx_parallel_data
			rx_parallel_data(1)       => alt_sv_gx_latopt_x3_inst_rx_parallel_data(1),                                                                                                                                                                                                       --                   .rx_parallel_data
			rx_parallel_data(2)       => alt_sv_gx_latopt_x3_inst_rx_parallel_data(2),                                                                                                                                                                                                       --                   .rx_parallel_data
			rx_parallel_data(3)       => alt_sv_gx_latopt_x3_inst_rx_parallel_data(3),                                                                                                                                                                                                       --                   .rx_parallel_data
			rx_parallel_data(4)       => alt_sv_gx_latopt_x3_inst_rx_parallel_data(4),                                                                                                                                                                                                       --                   .rx_parallel_data
			rx_parallel_data(5)       => alt_sv_gx_latopt_x3_inst_rx_parallel_data(5),                                                                                                                                                                                                       --                   .rx_parallel_data
			rx_parallel_data(6)       => alt_sv_gx_latopt_x3_inst_rx_parallel_data(6),                                                                                                                                                                                                       --                   .rx_parallel_data
			rx_parallel_data(7)       => alt_sv_gx_latopt_x3_inst_rx_parallel_data(7),                                                                                                                                                                                                       --                   .rx_parallel_data
			rx_parallel_data(8)       => alt_sv_gx_latopt_x3_inst_rx_parallel_data(8),                                                                                                                                                                                                       --                   .rx_parallel_data
			rx_parallel_data(9)       => alt_sv_gx_latopt_x3_inst_rx_parallel_data(9),                                                                                                                                                                                                       --                   .rx_parallel_data
			rx_parallel_data(10)      => alt_sv_gx_latopt_x3_inst_rx_parallel_data(10),                                                                                                                                                                                                      --                   .rx_parallel_data
			rx_parallel_data(11)      => alt_sv_gx_latopt_x3_inst_rx_parallel_data(11),                                                                                                                                                                                                      --                   .rx_parallel_data
			rx_parallel_data(12)      => alt_sv_gx_latopt_x3_inst_rx_parallel_data(12),                                                                                                                                                                                                      --                   .rx_parallel_data
			rx_parallel_data(13)      => alt_sv_gx_latopt_x3_inst_rx_parallel_data(13),                                                                                                                                                                                                      --                   .rx_parallel_data
			rx_parallel_data(14)      => alt_sv_gx_latopt_x3_inst_rx_parallel_data(14),                                                                                                                                                                                                      --                   .rx_parallel_data
			rx_parallel_data(15)      => alt_sv_gx_latopt_x3_inst_rx_parallel_data(15),                                                                                                                                                                                                      --                   .rx_parallel_data
			rx_parallel_data(16)      => alt_sv_gx_latopt_x3_inst_rx_parallel_data(16),                                                                                                                                                                                                      --                   .rx_parallel_data
			rx_parallel_data(17)      => alt_sv_gx_latopt_x3_inst_rx_parallel_data(17),                                                                                                                                                                                                      --                   .rx_parallel_data
			rx_parallel_data(18)      => alt_sv_gx_latopt_x3_inst_rx_parallel_data(18),                                                                                                                                                                                                      --                   .rx_parallel_data
			rx_parallel_data(19)      => alt_sv_gx_latopt_x3_inst_rx_parallel_data(19),                                                                                                                                                                                                      --                   .rx_parallel_data
			rx_parallel_data(20)      => alt_sv_gx_latopt_x3_inst_rx_parallel_data(20),                                                                                                                                                                                                      --                   .rx_parallel_data
			rx_parallel_data(21)      => alt_sv_gx_latopt_x3_inst_rx_parallel_data(21),                                                                                                                                                                                                      --                   .rx_parallel_data
			rx_parallel_data(22)      => alt_sv_gx_latopt_x3_inst_rx_parallel_data(22),                                                                                                                                                                                                      --                   .rx_parallel_data
			rx_parallel_data(23)      => alt_sv_gx_latopt_x3_inst_rx_parallel_data(23),                                                                                                                                                                                                      --                   .rx_parallel_data
			rx_parallel_data(24)      => alt_sv_gx_latopt_x3_inst_rx_parallel_data(24),                                                                                                                                                                                                      --                   .rx_parallel_data
			rx_parallel_data(25)      => alt_sv_gx_latopt_x3_inst_rx_parallel_data(25),                                                                                                                                                                                                      --                   .rx_parallel_data
			rx_parallel_data(26)      => alt_sv_gx_latopt_x3_inst_rx_parallel_data(26),                                                                                                                                                                                                      --                   .rx_parallel_data
			rx_parallel_data(27)      => alt_sv_gx_latopt_x3_inst_rx_parallel_data(27),                                                                                                                                                                                                      --                   .rx_parallel_data
			rx_parallel_data(28)      => alt_sv_gx_latopt_x3_inst_rx_parallel_data(28),                                                                                                                                                                                                      --                   .rx_parallel_data
			rx_parallel_data(29)      => alt_sv_gx_latopt_x3_inst_rx_parallel_data(29),                                                                                                                                                                                                      --                   .rx_parallel_data
			rx_parallel_data(30)      => alt_sv_gx_latopt_x3_inst_rx_parallel_data(30),                                                                                                                                                                                                      --                   .rx_parallel_data
			rx_parallel_data(31)      => alt_sv_gx_latopt_x3_inst_rx_parallel_data(31),                                                                                                                                                                                                      --                   .rx_parallel_data
			rx_parallel_data(32)      => alt_sv_gx_latopt_x3_inst_rx_parallel_data(32),                                                                                                                                                                                                      --                   .rx_parallel_data
			rx_parallel_data(33)      => alt_sv_gx_latopt_x3_inst_rx_parallel_data(33),                                                                                                                                                                                                      --                   .rx_parallel_data
			rx_parallel_data(34)      => alt_sv_gx_latopt_x3_inst_rx_parallel_data(34),                                                                                                                                                                                                      --                   .rx_parallel_data
			rx_parallel_data(35)      => alt_sv_gx_latopt_x3_inst_rx_parallel_data(35),                                                                                                                                                                                                      --                   .rx_parallel_data
			rx_parallel_data(36)      => alt_sv_gx_latopt_x3_inst_rx_parallel_data(36),                                                                                                                                                                                                      --                   .rx_parallel_data
			rx_parallel_data(37)      => alt_sv_gx_latopt_x3_inst_rx_parallel_data(37),                                                                                                                                                                                                      --                   .rx_parallel_data
			rx_parallel_data(38)      => alt_sv_gx_latopt_x3_inst_rx_parallel_data(38),                                                                                                                                                                                                      --                   .rx_parallel_data
			rx_parallel_data(39)      => alt_sv_gx_latopt_x3_inst_rx_parallel_data(39),                                                                                                                                                                                                      --                   .rx_parallel_data
			rx_parallel_data(40)      => alt_sv_gx_latopt_x3_inst_rx_parallel_data(40),                                                                                                                                                                                                      --                   .rx_parallel_data
			rx_parallel_data(41)      => alt_sv_gx_latopt_x3_inst_rx_parallel_data(41),                                                                                                                                                                                                      --                   .rx_parallel_data
			rx_parallel_data(42)      => alt_sv_gx_latopt_x3_inst_rx_parallel_data(42),                                                                                                                                                                                                      --                   .rx_parallel_data
			rx_parallel_data(43)      => alt_sv_gx_latopt_x3_inst_rx_parallel_data(43),                                                                                                                                                                                                      --                   .rx_parallel_data
			rx_parallel_data(44)      => alt_sv_gx_latopt_x3_inst_rx_parallel_data(44),                                                                                                                                                                                                      --                   .rx_parallel_data
			rx_parallel_data(45)      => alt_sv_gx_latopt_x3_inst_rx_parallel_data(45),                                                                                                                                                                                                      --                   .rx_parallel_data
			rx_parallel_data(46)      => alt_sv_gx_latopt_x3_inst_rx_parallel_data(46),                                                                                                                                                                                                      --                   .rx_parallel_data
			rx_parallel_data(47)      => alt_sv_gx_latopt_x3_inst_rx_parallel_data(47),                                                                                                                                                                                                      --                   .rx_parallel_data
			rx_parallel_data(48)      => alt_sv_gx_latopt_x3_inst_rx_parallel_data(48),                                                                                                                                                                                                      --                   .rx_parallel_data
			rx_parallel_data(49)      => alt_sv_gx_latopt_x3_inst_rx_parallel_data(49),                                                                                                                                                                                                      --                   .rx_parallel_data
			rx_parallel_data(50)      => alt_sv_gx_latopt_x3_inst_rx_parallel_data(50),                                                                                                                                                                                                      --                   .rx_parallel_data
			rx_parallel_data(51)      => alt_sv_gx_latopt_x3_inst_rx_parallel_data(51),                                                                                                                                                                                                      --                   .rx_parallel_data
			rx_parallel_data(52)      => alt_sv_gx_latopt_x3_inst_rx_parallel_data(52),                                                                                                                                                                                                      --                   .rx_parallel_data
			rx_parallel_data(53)      => alt_sv_gx_latopt_x3_inst_rx_parallel_data(53),                                                                                                                                                                                                      --                   .rx_parallel_data
			rx_parallel_data(54)      => alt_sv_gx_latopt_x3_inst_rx_parallel_data(54),                                                                                                                                                                                                      --                   .rx_parallel_data
			rx_parallel_data(55)      => alt_sv_gx_latopt_x3_inst_rx_parallel_data(55),                                                                                                                                                                                                      --                   .rx_parallel_data
			rx_parallel_data(56)      => alt_sv_gx_latopt_x3_inst_rx_parallel_data(56),                                                                                                                                                                                                      --                   .rx_parallel_data
			rx_parallel_data(57)      => alt_sv_gx_latopt_x3_inst_rx_parallel_data(57),                                                                                                                                                                                                      --                   .rx_parallel_data
			rx_parallel_data(58)      => alt_sv_gx_latopt_x3_inst_rx_parallel_data(58),                                                                                                                                                                                                      --                   .rx_parallel_data
			rx_parallel_data(59)      => alt_sv_gx_latopt_x3_inst_rx_parallel_data(59),                                                                                                                                                                                                      --                   .rx_parallel_data
			rx_parallel_data(60)      => alt_sv_gx_latopt_x3_inst_rx_parallel_data(60),                                                                                                                                                                                                      --                   .rx_parallel_data
			rx_parallel_data(61)      => alt_sv_gx_latopt_x3_inst_rx_parallel_data(61),                                                                                                                                                                                                      --                   .rx_parallel_data
			rx_parallel_data(62)      => alt_sv_gx_latopt_x3_inst_rx_parallel_data(62),                                                                                                                                                                                                      --                   .rx_parallel_data
			rx_parallel_data(63)      => alt_sv_gx_latopt_x3_inst_rx_parallel_data(63),                                                                                                                                                                                                      --                   .rx_parallel_data
			rx_parallel_data(64)      => alt_sv_gx_latopt_x3_inst_rx_parallel_data(64),                                                                                                                                                                                                      --                   .rx_parallel_data
			rx_parallel_data(65)      => alt_sv_gx_latopt_x3_inst_rx_parallel_data(65),                                                                                                                                                                                                      --                   .rx_parallel_data
			rx_parallel_data(66)      => alt_sv_gx_latopt_x3_inst_rx_parallel_data(66),                                                                                                                                                                                                      --                   .rx_parallel_data
			rx_parallel_data(67)      => alt_sv_gx_latopt_x3_inst_rx_parallel_data(67),                                                                                                                                                                                                      --                   .rx_parallel_data
			rx_parallel_data(68)      => alt_sv_gx_latopt_x3_inst_rx_parallel_data(68),                                                                                                                                                                                                      --                   .rx_parallel_data
			rx_parallel_data(69)      => alt_sv_gx_latopt_x3_inst_rx_parallel_data(69),                                                                                                                                                                                                      --                   .rx_parallel_data
			rx_parallel_data(70)      => alt_sv_gx_latopt_x3_inst_rx_parallel_data(70),                                                                                                                                                                                                      --                   .rx_parallel_data
			rx_parallel_data(71)      => alt_sv_gx_latopt_x3_inst_rx_parallel_data(71),                                                                                                                                                                                                      --                   .rx_parallel_data
			rx_parallel_data(72)      => alt_sv_gx_latopt_x3_inst_rx_parallel_data(72),                                                                                                                                                                                                      --                   .rx_parallel_data
			rx_parallel_data(73)      => alt_sv_gx_latopt_x3_inst_rx_parallel_data(73),                                                                                                                                                                                                      --                   .rx_parallel_data
			rx_parallel_data(74)      => alt_sv_gx_latopt_x3_inst_rx_parallel_data(74),                                                                                                                                                                                                      --                   .rx_parallel_data
			rx_parallel_data(75)      => alt_sv_gx_latopt_x3_inst_rx_parallel_data(75),                                                                                                                                                                                                      --                   .rx_parallel_data
			rx_parallel_data(76)      => alt_sv_gx_latopt_x3_inst_rx_parallel_data(76),                                                                                                                                                                                                      --                   .rx_parallel_data
			rx_parallel_data(77)      => alt_sv_gx_latopt_x3_inst_rx_parallel_data(77),                                                                                                                                                                                                      --                   .rx_parallel_data
			rx_parallel_data(78)      => alt_sv_gx_latopt_x3_inst_rx_parallel_data(78),                                                                                                                                                                                                      --                   .rx_parallel_data
			rx_parallel_data(79)      => alt_sv_gx_latopt_x3_inst_rx_parallel_data(79),                                                                                                                                                                                                      --                   .rx_parallel_data
			rx_parallel_data(80)      => alt_sv_gx_latopt_x3_inst_rx_parallel_data(80),                                                                                                                                                                                                      --                   .rx_parallel_data
			rx_parallel_data(81)      => alt_sv_gx_latopt_x3_inst_rx_parallel_data(81),                                                                                                                                                                                                      --                   .rx_parallel_data
			rx_parallel_data(82)      => alt_sv_gx_latopt_x3_inst_rx_parallel_data(82),                                                                                                                                                                                                      --                   .rx_parallel_data
			rx_parallel_data(83)      => alt_sv_gx_latopt_x3_inst_rx_parallel_data(83),                                                                                                                                                                                                      --                   .rx_parallel_data
			rx_parallel_data(84)      => alt_sv_gx_latopt_x3_inst_rx_parallel_data(84),                                                                                                                                                                                                      --                   .rx_parallel_data
			rx_parallel_data(85)      => alt_sv_gx_latopt_x3_inst_rx_parallel_data(85),                                                                                                                                                                                                      --                   .rx_parallel_data
			rx_parallel_data(86)      => alt_sv_gx_latopt_x3_inst_rx_parallel_data(86),                                                                                                                                                                                                      --                   .rx_parallel_data
			rx_parallel_data(87)      => alt_sv_gx_latopt_x3_inst_rx_parallel_data(87),                                                                                                                                                                                                      --                   .rx_parallel_data
			rx_parallel_data(88)      => alt_sv_gx_latopt_x3_inst_rx_parallel_data(88),                                                                                                                                                                                                      --                   .rx_parallel_data
			rx_parallel_data(89)      => alt_sv_gx_latopt_x3_inst_rx_parallel_data(89),                                                                                                                                                                                                      --                   .rx_parallel_data
			rx_parallel_data(90)      => alt_sv_gx_latopt_x3_inst_rx_parallel_data(90),                                                                                                                                                                                                      --                   .rx_parallel_data
			rx_parallel_data(91)      => alt_sv_gx_latopt_x3_inst_rx_parallel_data(91),                                                                                                                                                                                                      --                   .rx_parallel_data
			rx_parallel_data(92)      => alt_sv_gx_latopt_x3_inst_rx_parallel_data(92),                                                                                                                                                                                                      --                   .rx_parallel_data
			rx_parallel_data(93)      => alt_sv_gx_latopt_x3_inst_rx_parallel_data(93),                                                                                                                                                                                                      --                   .rx_parallel_data
			rx_parallel_data(94)      => alt_sv_gx_latopt_x3_inst_rx_parallel_data(94),                                                                                                                                                                                                      --                   .rx_parallel_data
			rx_parallel_data(95)      => alt_sv_gx_latopt_x3_inst_rx_parallel_data(95),                                                                                                                                                                                                      --                   .rx_parallel_data
			rx_parallel_data(96)      => alt_sv_gx_latopt_x3_inst_rx_parallel_data(96),                                                                                                                                                                                                      --                   .rx_parallel_data
			rx_parallel_data(97)      => alt_sv_gx_latopt_x3_inst_rx_parallel_data(97),                                                                                                                                                                                                      --                   .rx_parallel_data
			rx_parallel_data(98)      => alt_sv_gx_latopt_x3_inst_rx_parallel_data(98),                                                                                                                                                                                                      --                   .rx_parallel_data
			rx_parallel_data(99)      => alt_sv_gx_latopt_x3_inst_rx_parallel_data(99),                                                                                                                                                                                                      --                   .rx_parallel_data
			rx_parallel_data(100)     => alt_sv_gx_latopt_x3_inst_rx_parallel_data(100),                                                                                                                                                                                                     --                   .rx_parallel_data
			rx_parallel_data(101)     => alt_sv_gx_latopt_x3_inst_rx_parallel_data(101),                                                                                                                                                                                                     --                   .rx_parallel_data
			rx_parallel_data(102)     => alt_sv_gx_latopt_x3_inst_rx_parallel_data(102),                                                                                                                                                                                                     --                   .rx_parallel_data
			rx_parallel_data(103)     => alt_sv_gx_latopt_x3_inst_rx_parallel_data(103),                                                                                                                                                                                                     --                   .rx_parallel_data
			rx_parallel_data(104)     => alt_sv_gx_latopt_x3_inst_rx_parallel_data(104),                                                                                                                                                                                                     --                   .rx_parallel_data
			rx_parallel_data(105)     => alt_sv_gx_latopt_x3_inst_rx_parallel_data(105),                                                                                                                                                                                                     --                   .rx_parallel_data
			rx_parallel_data(106)     => alt_sv_gx_latopt_x3_inst_rx_parallel_data(106),                                                                                                                                                                                                     --                   .rx_parallel_data
			rx_parallel_data(107)     => alt_sv_gx_latopt_x3_inst_rx_parallel_data(107),                                                                                                                                                                                                     --                   .rx_parallel_data
			rx_parallel_data(108)     => alt_sv_gx_latopt_x3_inst_rx_parallel_data(108),                                                                                                                                                                                                     --                   .rx_parallel_data
			rx_parallel_data(109)     => alt_sv_gx_latopt_x3_inst_rx_parallel_data(109),                                                                                                                                                                                                     --                   .rx_parallel_data
			rx_parallel_data(110)     => alt_sv_gx_latopt_x3_inst_rx_parallel_data(110),                                                                                                                                                                                                     --                   .rx_parallel_data
			rx_parallel_data(111)     => alt_sv_gx_latopt_x3_inst_rx_parallel_data(111),                                                                                                                                                                                                     --                   .rx_parallel_data
			rx_parallel_data(112)     => alt_sv_gx_latopt_x3_inst_rx_parallel_data(112),                                                                                                                                                                                                     --                   .rx_parallel_data
			rx_parallel_data(113)     => alt_sv_gx_latopt_x3_inst_rx_parallel_data(113),                                                                                                                                                                                                     --                   .rx_parallel_data
			rx_parallel_data(114)     => alt_sv_gx_latopt_x3_inst_rx_parallel_data(114),                                                                                                                                                                                                     --                   .rx_parallel_data
			rx_parallel_data(115)     => alt_sv_gx_latopt_x3_inst_rx_parallel_data(115),                                                                                                                                                                                                     --                   .rx_parallel_data
			rx_parallel_data(116)     => alt_sv_gx_latopt_x3_inst_rx_parallel_data(116),                                                                                                                                                                                                     --                   .rx_parallel_data
			rx_parallel_data(117)     => alt_sv_gx_latopt_x3_inst_rx_parallel_data(117),                                                                                                                                                                                                     --                   .rx_parallel_data
			rx_parallel_data(118)     => alt_sv_gx_latopt_x3_inst_rx_parallel_data(118),                                                                                                                                                                                                     --                   .rx_parallel_data
			rx_parallel_data(119)     => alt_sv_gx_latopt_x3_inst_rx_parallel_data(119),                                                                                                                                                                                                     --                   .rx_parallel_data
			rx_parallel_data(120)     => alt_sv_gx_latopt_x3_inst_rx_parallel_data(120),                                                                                                                                                                                                     --                   .rx_parallel_data
			rx_parallel_data(121)     => alt_sv_gx_latopt_x3_inst_rx_parallel_data(121),                                                                                                                                                                                                     --                   .rx_parallel_data
			rx_parallel_data(122)     => alt_sv_gx_latopt_x3_inst_rx_parallel_data(122),                                                                                                                                                                                                     --                   .rx_parallel_data
			rx_parallel_data(123)     => alt_sv_gx_latopt_x3_inst_rx_parallel_data(123),                                                                                                                                                                                                     --                   .rx_parallel_data
			rx_parallel_data(124)     => alt_sv_gx_latopt_x3_inst_rx_parallel_data(124),                                                                                                                                                                                                     --                   .rx_parallel_data
			rx_parallel_data(125)     => alt_sv_gx_latopt_x3_inst_rx_parallel_data(125),                                                                                                                                                                                                     --                   .rx_parallel_data
			rx_parallel_data(126)     => alt_sv_gx_latopt_x3_inst_rx_parallel_data(126),                                                                                                                                                                                                     --                   .rx_parallel_data
			rx_parallel_data(127)     => alt_sv_gx_latopt_x3_inst_rx_parallel_data(127),                                                                                                                                                                                                     --                   .rx_parallel_data
			rx_parallel_data(128)     => alt_sv_gx_latopt_x3_inst_rx_parallel_data(128),                                                                                                                                                                                                     --                   .rx_parallel_data
			rx_parallel_data(129)     => alt_sv_gx_latopt_x3_inst_rx_parallel_data(129),                                                                                                                                                                                                     --                   .rx_parallel_data
			rx_parallel_data(130)     => alt_sv_gx_latopt_x3_inst_rx_parallel_data(130),                                                                                                                                                                                                     --                   .rx_parallel_data
			rx_parallel_data(131)     => alt_sv_gx_latopt_x3_inst_rx_parallel_data(131),                                                                                                                                                                                                     --                   .rx_parallel_data
			rx_parallel_data(132)     => alt_sv_gx_latopt_x3_inst_rx_parallel_data(132),                                                                                                                                                                                                     --                   .rx_parallel_data
			rx_parallel_data(133)     => alt_sv_gx_latopt_x3_inst_rx_parallel_data(133),                                                                                                                                                                                                     --                   .rx_parallel_data
			rx_parallel_data(134)     => alt_sv_gx_latopt_x3_inst_rx_parallel_data(134),                                                                                                                                                                                                     --                   .rx_parallel_data
			rx_parallel_data(135)     => alt_sv_gx_latopt_x3_inst_rx_parallel_data(135),                                                                                                                                                                                                     --                   .rx_parallel_data
			rx_parallel_data(136)     => alt_sv_gx_latopt_x3_inst_rx_parallel_data(136),                                                                                                                                                                                                     --                   .rx_parallel_data
			rx_parallel_data(137)     => alt_sv_gx_latopt_x3_inst_rx_parallel_data(137),                                                                                                                                                                                                     --                   .rx_parallel_data
			rx_parallel_data(138)     => alt_sv_gx_latopt_x3_inst_rx_parallel_data(138),                                                                                                                                                                                                     --                   .rx_parallel_data
			rx_parallel_data(139)     => alt_sv_gx_latopt_x3_inst_rx_parallel_data(139),                                                                                                                                                                                                     --                   .rx_parallel_data
			rx_parallel_data(140)     => alt_sv_gx_latopt_x3_inst_rx_parallel_data(140),                                                                                                                                                                                                     --                   .rx_parallel_data
			rx_parallel_data(141)     => alt_sv_gx_latopt_x3_inst_rx_parallel_data(141),                                                                                                                                                                                                     --                   .rx_parallel_data
			rx_parallel_data(142)     => alt_sv_gx_latopt_x3_inst_rx_parallel_data(142),                                                                                                                                                                                                     --                   .rx_parallel_data
			rx_parallel_data(143)     => alt_sv_gx_latopt_x3_inst_rx_parallel_data(143),                                                                                                                                                                                                     --                   .rx_parallel_data
			rx_parallel_data(144)     => alt_sv_gx_latopt_x3_inst_rx_parallel_data(144),                                                                                                                                                                                                     --                   .rx_parallel_data
			rx_parallel_data(145)     => alt_sv_gx_latopt_x3_inst_rx_parallel_data(145),                                                                                                                                                                                                     --                   .rx_parallel_data
			rx_parallel_data(146)     => alt_sv_gx_latopt_x3_inst_rx_parallel_data(146),                                                                                                                                                                                                     --                   .rx_parallel_data
			rx_parallel_data(147)     => alt_sv_gx_latopt_x3_inst_rx_parallel_data(147),                                                                                                                                                                                                     --                   .rx_parallel_data
			rx_parallel_data(148)     => alt_sv_gx_latopt_x3_inst_rx_parallel_data(148),                                                                                                                                                                                                     --                   .rx_parallel_data
			rx_parallel_data(149)     => alt_sv_gx_latopt_x3_inst_rx_parallel_data(149),                                                                                                                                                                                                     --                   .rx_parallel_data
			rx_parallel_data(150)     => alt_sv_gx_latopt_x3_inst_rx_parallel_data(150),                                                                                                                                                                                                     --                   .rx_parallel_data
			rx_parallel_data(151)     => alt_sv_gx_latopt_x3_inst_rx_parallel_data(151),                                                                                                                                                                                                     --                   .rx_parallel_data
			rx_parallel_data(152)     => alt_sv_gx_latopt_x3_inst_rx_parallel_data(152),                                                                                                                                                                                                     --                   .rx_parallel_data
			rx_parallel_data(153)     => alt_sv_gx_latopt_x3_inst_rx_parallel_data(153),                                                                                                                                                                                                     --                   .rx_parallel_data
			rx_parallel_data(154)     => alt_sv_gx_latopt_x3_inst_rx_parallel_data(154),                                                                                                                                                                                                     --                   .rx_parallel_data
			rx_parallel_data(155)     => alt_sv_gx_latopt_x3_inst_rx_parallel_data(155),                                                                                                                                                                                                     --                   .rx_parallel_data
			rx_parallel_data(156)     => alt_sv_gx_latopt_x3_inst_rx_parallel_data(156),                                                                                                                                                                                                     --                   .rx_parallel_data
			rx_parallel_data(157)     => alt_sv_gx_latopt_x3_inst_rx_parallel_data(157),                                                                                                                                                                                                     --                   .rx_parallel_data
			rx_parallel_data(158)     => alt_sv_gx_latopt_x3_inst_rx_parallel_data(158),                                                                                                                                                                                                     --                   .rx_parallel_data
			rx_parallel_data(159)     => alt_sv_gx_latopt_x3_inst_rx_parallel_data(159),                                                                                                                                                                                                     --                   .rx_parallel_data
			rx_parallel_data(160)     => alt_sv_gx_latopt_x3_inst_rx_parallel_data(160),                                                                                                                                                                                                     --                   .rx_parallel_data
			rx_parallel_data(161)     => alt_sv_gx_latopt_x3_inst_rx_parallel_data(161),                                                                                                                                                                                                     --                   .rx_parallel_data
			rx_parallel_data(162)     => alt_sv_gx_latopt_x3_inst_rx_parallel_data(162),                                                                                                                                                                                                     --                   .rx_parallel_data
			rx_parallel_data(163)     => alt_sv_gx_latopt_x3_inst_rx_parallel_data(163),                                                                                                                                                                                                     --                   .rx_parallel_data
			rx_parallel_data(164)     => alt_sv_gx_latopt_x3_inst_rx_parallel_data(164),                                                                                                                                                                                                     --                   .rx_parallel_data
			rx_parallel_data(165)     => alt_sv_gx_latopt_x3_inst_rx_parallel_data(165),                                                                                                                                                                                                     --                   .rx_parallel_data
			rx_parallel_data(166)     => alt_sv_gx_latopt_x3_inst_rx_parallel_data(166),                                                                                                                                                                                                     --                   .rx_parallel_data
			rx_parallel_data(167)     => alt_sv_gx_latopt_x3_inst_rx_parallel_data(167),                                                                                                                                                                                                     --                   .rx_parallel_data
			rx_parallel_data(168)     => alt_sv_gx_latopt_x3_inst_rx_parallel_data(168),                                                                                                                                                                                                     --                   .rx_parallel_data
			rx_parallel_data(169)     => alt_sv_gx_latopt_x3_inst_rx_parallel_data(169),                                                                                                                                                                                                     --                   .rx_parallel_data
			rx_parallel_data(170)     => alt_sv_gx_latopt_x3_inst_rx_parallel_data(170),                                                                                                                                                                                                     --                   .rx_parallel_data
			rx_parallel_data(171)     => alt_sv_gx_latopt_x3_inst_rx_parallel_data(171),                                                                                                                                                                                                     --                   .rx_parallel_data
			rx_parallel_data(172)     => alt_sv_gx_latopt_x3_inst_rx_parallel_data(172),                                                                                                                                                                                                     --                   .rx_parallel_data
			rx_parallel_data(173)     => alt_sv_gx_latopt_x3_inst_rx_parallel_data(173),                                                                                                                                                                                                     --                   .rx_parallel_data
			rx_parallel_data(174)     => alt_sv_gx_latopt_x3_inst_rx_parallel_data(174),                                                                                                                                                                                                     --                   .rx_parallel_data
			rx_parallel_data(175)     => alt_sv_gx_latopt_x3_inst_rx_parallel_data(175),                                                                                                                                                                                                     --                   .rx_parallel_data
			rx_parallel_data(176)     => alt_sv_gx_latopt_x3_inst_rx_parallel_data(176),                                                                                                                                                                                                     --                   .rx_parallel_data
			rx_parallel_data(177)     => alt_sv_gx_latopt_x3_inst_rx_parallel_data(177),                                                                                                                                                                                                     --                   .rx_parallel_data
			rx_parallel_data(178)     => alt_sv_gx_latopt_x3_inst_rx_parallel_data(178),                                                                                                                                                                                                     --                   .rx_parallel_data
			rx_parallel_data(179)     => alt_sv_gx_latopt_x3_inst_rx_parallel_data(179),                                                                                                                                                                                                     --                   .rx_parallel_data
			rx_parallel_data(180)     => alt_sv_gx_latopt_x3_inst_rx_parallel_data(180),                                                                                                                                                                                                     --                   .rx_parallel_data
			rx_parallel_data(181)     => alt_sv_gx_latopt_x3_inst_rx_parallel_data(181),                                                                                                                                                                                                     --                   .rx_parallel_data
			rx_parallel_data(182)     => alt_sv_gx_latopt_x3_inst_rx_parallel_data(182),                                                                                                                                                                                                     --                   .rx_parallel_data
			rx_parallel_data(183)     => alt_sv_gx_latopt_x3_inst_rx_parallel_data(183),                                                                                                                                                                                                     --                   .rx_parallel_data
			rx_parallel_data(184)     => alt_sv_gx_latopt_x3_inst_rx_parallel_data(184),                                                                                                                                                                                                     --                   .rx_parallel_data
			rx_parallel_data(185)     => alt_sv_gx_latopt_x3_inst_rx_parallel_data(185),                                                                                                                                                                                                     --                   .rx_parallel_data
			rx_parallel_data(186)     => alt_sv_gx_latopt_x3_inst_rx_parallel_data(186),                                                                                                                                                                                                     --                   .rx_parallel_data
			rx_parallel_data(187)     => alt_sv_gx_latopt_x3_inst_rx_parallel_data(187),                                                                                                                                                                                                     --                   .rx_parallel_data
			rx_parallel_data(188)     => alt_sv_gx_latopt_x3_inst_rx_parallel_data(188),                                                                                                                                                                                                     --                   .rx_parallel_data
			rx_parallel_data(189)     => alt_sv_gx_latopt_x3_inst_rx_parallel_data(189),                                                                                                                                                                                                     --                   .rx_parallel_data
			rx_parallel_data(190)     => alt_sv_gx_latopt_x3_inst_rx_parallel_data(190),                                                                                                                                                                                                     --                   .rx_parallel_data
			rx_parallel_data(191)     => alt_sv_gx_latopt_x3_inst_rx_parallel_data(191),                                                                                                                                                                                                     --                   .rx_parallel_data
			tx_pll_refclk             => "0",                                                                                                                                                                                                                                                --        (terminated)
			tx_pma_clkout             => open,                                                                                                                                                                                                                                               --        (terminated)
			tx_pma_pclk               => open,                                                                                                                                                                                                                                               --        (terminated)
			tx_pma_parallel_data      => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", --        (terminated)
			pll_locked                => open,                                                                                                                                                                                                                                               --        (terminated)
			rx_pma_clkout             => open,                                                                                                                                                                                                                                               --        (terminated)
			rx_pma_pclk               => open,                                                                                                                                                                                                                                               --        (terminated)
			rx_pma_parallel_data      => open,                                                                                                                                                                                                                                               --        (terminated)
			rx_clklow                 => open,                                                                                                                                                                                                                                               --        (terminated)
			rx_fref                   => open,                                                                                                                                                                                                                                               --        (terminated)
			rx_set_locktodata         => "000",                                                                                                                                                                                                                                              --        (terminated)
			rx_set_locktoref          => "000",                                                                                                                                                                                                                                              --        (terminated)
			rx_signaldetect           => open,                                                                                                                                                                                                                                               --        (terminated)
			rx_pma_qpipulldn          => "000",                                                                                                                                                                                                                                              --        (terminated)
			tx_pma_qpipullup          => "000",                                                                                                                                                                                                                                              --        (terminated)
			tx_pma_qpipulldn          => "000",                                                                                                                                                                                                                                              --        (terminated)
			tx_pma_txdetectrx         => "000",                                                                                                                                                                                                                                              --        (terminated)
			tx_pma_rxfound            => open,                                                                                                                                                                                                                                               --        (terminated)
			rx_std_prbs_done          => open,                                                                                                                                                                                                                                               --        (terminated)
			rx_std_prbs_err           => open,                                                                                                                                                                                                                                               --        (terminated)
			tx_std_pcfifo_full        => open,                                                                                                                                                                                                                                               --        (terminated)
			tx_std_pcfifo_empty       => open,                                                                                                                                                                                                                                               --        (terminated)
			rx_std_pcfifo_full        => open,                                                                                                                                                                                                                                               --        (terminated)
			rx_std_pcfifo_empty       => open,                                                                                                                                                                                                                                               --        (terminated)
			rx_std_byteorder_ena      => "000",                                                                                                                                                                                                                                              --        (terminated)
			rx_std_byteorder_flag     => open,                                                                                                                                                                                                                                               --        (terminated)
			rx_std_rmfifo_full        => open,                                                                                                                                                                                                                                               --        (terminated)
			rx_std_rmfifo_empty       => open,                                                                                                                                                                                                                                               --        (terminated)
			rx_std_wa_patternalign    => "000",                                                                                                                                                                                                                                              --        (terminated)
			rx_std_wa_a1a2size        => "000",                                                                                                                                                                                                                                              --        (terminated)
			tx_std_bitslipboundarysel => "000000000000000",                                                                                                                                                                                                                                  --        (terminated)
			rx_std_bitslipboundarysel => open,                                                                                                                                                                                                                                               --        (terminated)
			rx_std_bitslip            => "000",                                                                                                                                                                                                                                              --        (terminated)
			rx_std_runlength_err      => open,                                                                                                                                                                                                                                               --        (terminated)
			rx_std_bitrev_ena         => "000",                                                                                                                                                                                                                                              --        (terminated)
			rx_std_byterev_ena        => "000",                                                                                                                                                                                                                                              --        (terminated)
			tx_std_elecidle           => "000",                                                                                                                                                                                                                                              --        (terminated)
			rx_std_signaldetect       => open,                                                                                                                                                                                                                                               --        (terminated)
			tx_10g_coreclkin          => "000",                                                                                                                                                                                                                                              --        (terminated)
			rx_10g_coreclkin          => "000",                                                                                                                                                                                                                                              --        (terminated)
			tx_10g_clkout             => open,                                                                                                                                                                                                                                               --        (terminated)
			rx_10g_clkout             => open,                                                                                                                                                                                                                                               --        (terminated)
			rx_10g_clk33out           => open,                                                                                                                                                                                                                                               --        (terminated)
			rx_10g_prbs_err_clr       => "000",                                                                                                                                                                                                                                              --        (terminated)
			rx_10g_prbs_done          => open,                                                                                                                                                                                                                                               --        (terminated)
			rx_10g_prbs_err           => open,                                                                                                                                                                                                                                               --        (terminated)
			tx_10g_control            => "000000000000000000000000000",                                                                                                                                                                                                                      --        (terminated)
			rx_10g_control            => open,                                                                                                                                                                                                                                               --        (terminated)
			tx_10g_data_valid         => "000",                                                                                                                                                                                                                                              --        (terminated)
			tx_10g_fifo_full          => open,                                                                                                                                                                                                                                               --        (terminated)
			tx_10g_fifo_pfull         => open,                                                                                                                                                                                                                                               --        (terminated)
			tx_10g_fifo_empty         => open,                                                                                                                                                                                                                                               --        (terminated)
			tx_10g_fifo_pempty        => open,                                                                                                                                                                                                                                               --        (terminated)
			tx_10g_fifo_del           => open,                                                                                                                                                                                                                                               --        (terminated)
			tx_10g_fifo_insert        => open,                                                                                                                                                                                                                                               --        (terminated)
			rx_10g_fifo_rd_en         => "000",                                                                                                                                                                                                                                              --        (terminated)
			rx_10g_data_valid         => open,                                                                                                                                                                                                                                               --        (terminated)
			rx_10g_fifo_full          => open,                                                                                                                                                                                                                                               --        (terminated)
			rx_10g_fifo_pfull         => open,                                                                                                                                                                                                                                               --        (terminated)
			rx_10g_fifo_empty         => open,                                                                                                                                                                                                                                               --        (terminated)
			rx_10g_fifo_pempty        => open,                                                                                                                                                                                                                                               --        (terminated)
			rx_10g_fifo_del           => open,                                                                                                                                                                                                                                               --        (terminated)
			rx_10g_fifo_insert        => open,                                                                                                                                                                                                                                               --        (terminated)
			rx_10g_fifo_align_val     => open,                                                                                                                                                                                                                                               --        (terminated)
			rx_10g_fifo_align_clr     => "000",                                                                                                                                                                                                                                              --        (terminated)
			rx_10g_fifo_align_en      => "000",                                                                                                                                                                                                                                              --        (terminated)
			tx_10g_frame              => open,                                                                                                                                                                                                                                               --        (terminated)
			tx_10g_frame_diag_status  => "000000",                                                                                                                                                                                                                                           --        (terminated)
			tx_10g_frame_burst_en     => "000",                                                                                                                                                                                                                                              --        (terminated)
			rx_10g_frame              => open,                                                                                                                                                                                                                                               --        (terminated)
			rx_10g_frame_lock         => open,                                                                                                                                                                                                                                               --        (terminated)
			rx_10g_frame_mfrm_err     => open,                                                                                                                                                                                                                                               --        (terminated)
			rx_10g_frame_sync_err     => open,                                                                                                                                                                                                                                               --        (terminated)
			rx_10g_frame_skip_ins     => open,                                                                                                                                                                                                                                               --        (terminated)
			rx_10g_frame_pyld_ins     => open,                                                                                                                                                                                                                                               --        (terminated)
			rx_10g_frame_skip_err     => open,                                                                                                                                                                                                                                               --        (terminated)
			rx_10g_frame_diag_err     => open,                                                                                                                                                                                                                                               --        (terminated)
			rx_10g_frame_diag_status  => open,                                                                                                                                                                                                                                               --        (terminated)
			rx_10g_crc32_err          => open,                                                                                                                                                                                                                                               --        (terminated)
			rx_10g_descram_err        => open,                                                                                                                                                                                                                                               --        (terminated)
			rx_10g_blk_lock           => open,                                                                                                                                                                                                                                               --        (terminated)
			rx_10g_blk_sh_err         => open,                                                                                                                                                                                                                                               --        (terminated)
			tx_10g_bitslip            => "000000000000000000000",                                                                                                                                                                                                                            --        (terminated)
			rx_10g_bitslip            => "000",                                                                                                                                                                                                                                              --        (terminated)
			rx_10g_highber            => open,                                                                                                                                                                                                                                               --        (terminated)
			rx_10g_highber_clr_cnt    => "000",                                                                                                                                                                                                                                              --        (terminated)
			rx_10g_clr_errblk_count   => "000"                                                                                                                                                                                                                                               --        (terminated)
		);

	rx_parallel_data <= alt_sv_gx_latopt_x3_inst_rx_parallel_data(185) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(184) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(183) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(182) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(181) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(180) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(179) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(178) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(177) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(176) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(169) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(168) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(167) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(166) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(165) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(164) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(163) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(162) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(161) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(160) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(153) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(152) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(151) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(150) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(149) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(148) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(147) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(146) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(145) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(144) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(137) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(136) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(135) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(134) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(133) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(132) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(131) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(130) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(129) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(128) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(121) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(120) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(119) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(118) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(117) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(116) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(115) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(114) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(113) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(112) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(105) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(104) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(103) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(102) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(101) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(100) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(99) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(98) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(97) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(96) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(89) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(88) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(87) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(86) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(85) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(84) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(83) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(82) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(81) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(80) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(73) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(72) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(71) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(70) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(69) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(68) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(67) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(66) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(65) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(64) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(57) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(56) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(55) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(54) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(53) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(52) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(51) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(50) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(49) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(48) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(41) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(40) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(39) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(38) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(37) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(36) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(35) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(34) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(33) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(32) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(25) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(24) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(23) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(22) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(21) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(20) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(19) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(18) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(17) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(16) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(9) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(8) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(7) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(6) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(5) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(4) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(3) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(2) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(1) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(0);

	unused_rx_parallel_data <= alt_sv_gx_latopt_x3_inst_rx_parallel_data(191) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(190) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(189) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(188) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(187) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(186) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(175) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(174) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(173) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(172) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(171) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(170) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(159) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(158) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(157) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(156) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(155) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(154) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(143) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(142) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(141) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(140) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(139) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(138) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(127) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(126) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(125) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(124) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(123) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(122) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(111) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(110) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(109) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(108) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(107) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(106) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(95) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(94) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(93) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(92) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(91) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(90) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(79) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(78) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(77) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(76) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(75) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(74) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(63) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(62) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(61) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(60) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(59) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(58) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(47) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(46) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(45) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(44) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(43) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(42) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(31) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(30) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(29) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(28) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(27) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(26) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(15) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(14) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(13) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(12) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(11) & alt_sv_gx_latopt_x3_inst_rx_parallel_data(10);

end architecture rtl; -- of alt_sv_gx_latopt_x3
-- Retrieval info: <?xml version="1.0"?>
--<!--
--	Generated by Altera MegaWizard Launcher Utility version 1.0
--	************************************************************
--	THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--	************************************************************
--	Copyright (C) 1991-2016 Altera Corporation
--	Any megafunction design, and related net list (encrypted or decrypted),
--	support information, device programming or simulation file, and any other
--	associated documentation or information provided by Altera or a partner
--	under Altera's Megafunction Partnership Program may be used only to
--	program PLD devices (but not masked PLD devices) from Altera.  Any other
--	use of such megafunction design, net list, support information, device
--	programming or simulation file, or any other related documentation or
--	information is prohibited for any other purpose, including, but not
--	limited to modification, reverse engineering, de-compiling, or use with
--	any other silicon devices, unless such use is explicitly licensed under
--	a separate agreement with Altera or a megafunction partner.  Title to
--	the intellectual property, including patents, copyrights, trademarks,
--	trade secrets, or maskworks, embodied in any such megafunction design,
--	net list, support information, device programming or simulation file, or
--	any other related documentation or information provided by Altera or a
--	megafunction partner, remains with Altera, the megafunction partner, or
--	their respective licensors.  No other licenses, including any licenses
--	needed under any third party's intellectual property, are provided herein.
---->
-- Retrieval info: <instance entity-name="altera_xcvr_native_sv" version="16.0" >
-- Retrieval info: 	<generic name="device_family" value="Stratix V" />
-- Retrieval info: 	<generic name="show_advanced_features" value="0" />
-- Retrieval info: 	<generic name="device_speedgrade" value="fastest" />
-- Retrieval info: 	<generic name="message_level" value="error" />
-- Retrieval info: 	<generic name="tx_enable" value="1" />
-- Retrieval info: 	<generic name="rx_enable" value="1" />
-- Retrieval info: 	<generic name="enable_std" value="1" />
-- Retrieval info: 	<generic name="enable_teng" value="0" />
-- Retrieval info: 	<generic name="set_data_path_select" value="standard" />
-- Retrieval info: 	<generic name="channels" value="3" />
-- Retrieval info: 	<generic name="bonded_mode" value="xN" />
-- Retrieval info: 	<generic name="enable_simple_interface" value="1" />
-- Retrieval info: 	<generic name="set_data_rate" value="4800" />
-- Retrieval info: 	<generic name="pma_direct_width" value="80" />
-- Retrieval info: 	<generic name="tx_pma_clk_div" value="1" />
-- Retrieval info: 	<generic name="pll_reconfig_enable" value="0" />
-- Retrieval info: 	<generic name="pll_external_enable" value="1" />
-- Retrieval info: 	<generic name="plls" value="1" />
-- Retrieval info: 	<generic name="pll_select" value="0" />
-- Retrieval info: 	<generic name="pll_refclk_cnt" value="1" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll0_pll_type" value="CMU" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll1_pll_type" value="CMU" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll2_pll_type" value="CMU" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll3_pll_type" value="CMU" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll0_data_rate" value="1250 Mbps" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll1_data_rate" value="1250 Mbps" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll2_data_rate" value="1250 Mbps" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll3_data_rate" value="1250 Mbps" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll0_refclk_freq" value="240.0 MHz" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll1_refclk_freq" value="125.0 MHz" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll2_refclk_freq" value="125.0 MHz" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll3_refclk_freq" value="125.0 MHz" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll0_refclk_sel" value="0" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll1_refclk_sel" value="0" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll2_refclk_sel" value="0" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll3_refclk_sel" value="0" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll0_clk_network" value="x1" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll1_clk_network" value="x1" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll2_clk_network" value="x1" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll3_clk_network" value="x1" />
-- Retrieval info: 	<generic name="cdr_reconfig_enable" value="0" />
-- Retrieval info: 	<generic name="cdr_refclk_cnt" value="1" />
-- Retrieval info: 	<generic name="cdr_refclk_select" value="0" />
-- Retrieval info: 	<generic name="set_cdr_refclk_freq" value="120.0 MHz" />
-- Retrieval info: 	<generic name="rx_ppm_detect_threshold" value="1000" />
-- Retrieval info: 	<generic name="enable_port_tx_pma_qpipullup" value="0" />
-- Retrieval info: 	<generic name="enable_port_tx_pma_qpipulldn" value="0" />
-- Retrieval info: 	<generic name="enable_port_tx_pma_txdetectrx" value="0" />
-- Retrieval info: 	<generic name="enable_port_tx_pma_rxfound" value="0" />
-- Retrieval info: 	<generic name="enable_port_tx_pma_pclk" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_pma_qpipulldn" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_pma_clkout" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_pma_pclk" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_is_lockedtodata" value="1" />
-- Retrieval info: 	<generic name="enable_port_rx_is_lockedtoref" value="1" />
-- Retrieval info: 	<generic name="enable_ports_rx_manual_cdr_mode" value="0" />
-- Retrieval info: 	<generic name="rx_clkslip_enable" value="1" />
-- Retrieval info: 	<generic name="enable_port_rx_signaldetect" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_seriallpbken" value="1" />
-- Retrieval info: 	<generic name="std_protocol_hint" value="basic" />
-- Retrieval info: 	<generic name="std_pcs_pma_width" value="20" />
-- Retrieval info: 	<generic name="std_low_latency_bypass_enable" value="1" />
-- Retrieval info: 	<generic name="std_tx_pcfifo_mode" value="register_fifo" />
-- Retrieval info: 	<generic name="std_rx_pcfifo_mode" value="register_fifo" />
-- Retrieval info: 	<generic name="enable_port_tx_std_pcfifo_full" value="0" />
-- Retrieval info: 	<generic name="enable_port_tx_std_pcfifo_empty" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_std_pcfifo_full" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_std_pcfifo_empty" value="0" />
-- Retrieval info: 	<generic name="std_rx_byte_order_enable" value="0" />
-- Retrieval info: 	<generic name="std_rx_byte_order_mode" value="manual" />
-- Retrieval info: 	<generic name="std_rx_byte_order_symbol_count" value="1" />
-- Retrieval info: 	<generic name="std_rx_byte_order_pattern" value="0" />
-- Retrieval info: 	<generic name="std_rx_byte_order_pad" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_std_byteorder_ena" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_std_byteorder_flag" value="0" />
-- Retrieval info: 	<generic name="std_tx_byte_ser_enable" value="1" />
-- Retrieval info: 	<generic name="std_rx_byte_deser_enable" value="1" />
-- Retrieval info: 	<generic name="std_tx_8b10b_enable" value="0" />
-- Retrieval info: 	<generic name="std_tx_8b10b_disp_ctrl_enable" value="0" />
-- Retrieval info: 	<generic name="std_rx_8b10b_enable" value="0" />
-- Retrieval info: 	<generic name="std_rx_rmfifo_enable" value="0" />
-- Retrieval info: 	<generic name="std_rx_rmfifo_pattern_p" value="00000" />
-- Retrieval info: 	<generic name="std_rx_rmfifo_pattern_n" value="00000" />
-- Retrieval info: 	<generic name="enable_port_rx_std_rmfifo_full" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_std_rmfifo_empty" value="0" />
-- Retrieval info: 	<generic name="std_tx_bitslip_enable" value="0" />
-- Retrieval info: 	<generic name="enable_port_tx_std_bitslipboundarysel" value="0" />
-- Retrieval info: 	<generic name="std_rx_word_aligner_mode" value="bit_slip" />
-- Retrieval info: 	<generic name="std_rx_word_aligner_pattern_len" value="7" />
-- Retrieval info: 	<generic name="std_rx_word_aligner_pattern" value="0000000000" />
-- Retrieval info: 	<generic name="std_rx_word_aligner_rknumber" value="3" />
-- Retrieval info: 	<generic name="std_rx_word_aligner_renumber" value="3" />
-- Retrieval info: 	<generic name="std_rx_word_aligner_rgnumber" value="3" />
-- Retrieval info: 	<generic name="std_rx_run_length_val" value="31" />
-- Retrieval info: 	<generic name="enable_port_rx_std_wa_patternalign" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_std_wa_a1a2size" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_std_bitslipboundarysel" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_std_bitslip" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_std_runlength_err" value="0" />
-- Retrieval info: 	<generic name="std_tx_bitrev_enable" value="0" />
-- Retrieval info: 	<generic name="std_rx_bitrev_enable" value="0" />
-- Retrieval info: 	<generic name="std_tx_byterev_enable" value="0" />
-- Retrieval info: 	<generic name="std_rx_byterev_enable" value="0" />
-- Retrieval info: 	<generic name="std_tx_polinv_enable" value="1" />
-- Retrieval info: 	<generic name="std_rx_polinv_enable" value="1" />
-- Retrieval info: 	<generic name="enable_port_rx_std_bitrev_ena" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_std_byterev_ena" value="0" />
-- Retrieval info: 	<generic name="enable_port_tx_std_polinv" value="1" />
-- Retrieval info: 	<generic name="enable_port_rx_std_polinv" value="1" />
-- Retrieval info: 	<generic name="enable_port_tx_std_elecidle" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_std_signaldetect" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_std_prbs_status" value="0" />
-- Retrieval info: 	<generic name="teng_protocol_hint" value="basic" />
-- Retrieval info: 	<generic name="teng_pcs_pma_width" value="40" />
-- Retrieval info: 	<generic name="teng_pld_pcs_width" value="40" />
-- Retrieval info: 	<generic name="teng_txfifo_mode" value="phase_comp" />
-- Retrieval info: 	<generic name="teng_txfifo_full" value="31" />
-- Retrieval info: 	<generic name="teng_txfifo_empty" value="0" />
-- Retrieval info: 	<generic name="teng_txfifo_pfull" value="23" />
-- Retrieval info: 	<generic name="teng_txfifo_pempty" value="2" />
-- Retrieval info: 	<generic name="enable_port_tx_10g_fifo_full" value="0" />
-- Retrieval info: 	<generic name="enable_port_tx_10g_fifo_pfull" value="0" />
-- Retrieval info: 	<generic name="enable_port_tx_10g_fifo_empty" value="0" />
-- Retrieval info: 	<generic name="enable_port_tx_10g_fifo_pempty" value="0" />
-- Retrieval info: 	<generic name="enable_port_tx_10g_fifo_del" value="0" />
-- Retrieval info: 	<generic name="enable_port_tx_10g_fifo_insert" value="0" />
-- Retrieval info: 	<generic name="teng_rxfifo_mode" value="phase_comp" />
-- Retrieval info: 	<generic name="teng_rxfifo_full" value="31" />
-- Retrieval info: 	<generic name="teng_rxfifo_empty" value="0" />
-- Retrieval info: 	<generic name="teng_rxfifo_pfull" value="23" />
-- Retrieval info: 	<generic name="teng_rxfifo_pempty" value="2" />
-- Retrieval info: 	<generic name="teng_rxfifo_align_del" value="0" />
-- Retrieval info: 	<generic name="teng_rxfifo_control_del" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_10g_data_valid" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_10g_fifo_full" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_10g_fifo_pfull" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_10g_fifo_empty" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_10g_fifo_pempty" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_10g_fifo_del" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_10g_fifo_insert" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_10g_fifo_rd_en" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_10g_fifo_align_val" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_10g_fifo_align_clr" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_10g_fifo_align_en" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_10g_clk33out" value="0" />
-- Retrieval info: 	<generic name="teng_tx_frmgen_user_length" value="2048" />
-- Retrieval info: 	<generic name="teng_tx_frmgen_burst_enable" value="0" />
-- Retrieval info: 	<generic name="enable_port_tx_10g_frame" value="0" />
-- Retrieval info: 	<generic name="enable_port_tx_10g_frame_diag_status" value="0" />
-- Retrieval info: 	<generic name="enable_port_tx_10g_frame_burst_en" value="0" />
-- Retrieval info: 	<generic name="teng_rx_frmsync_user_length" value="2048" />
-- Retrieval info: 	<generic name="enable_port_rx_10g_frame" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_10g_frame_lock" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_10g_frame_mfrm_err" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_10g_frame_sync_err" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_10g_frame_pyld_ins" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_10g_frame_skip_ins" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_10g_frame_skip_err" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_10g_frame_diag_err" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_10g_frame_diag_status" value="0" />
-- Retrieval info: 	<generic name="teng_tx_sh_err" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_10g_crc32_err" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_10g_highber" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_10g_highber_clr_cnt" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_10g_clr_errblk_count" value="0" />
-- Retrieval info: 	<generic name="teng_tx_scram_user_seed" value="000000000000000" />
-- Retrieval info: 	<generic name="enable_port_rx_10g_descram_err" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_10g_blk_lock" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_10g_blk_sh_err" value="0" />
-- Retrieval info: 	<generic name="teng_tx_polinv_enable" value="0" />
-- Retrieval info: 	<generic name="teng_tx_bitslip_enable" value="0" />
-- Retrieval info: 	<generic name="teng_rx_polinv_enable" value="0" />
-- Retrieval info: 	<generic name="teng_rx_bitslip_enable" value="0" />
-- Retrieval info: 	<generic name="enable_port_tx_10g_bitslip" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_10g_bitslip" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_teng_prbs_status" value="0" />
-- Retrieval info: </instance>
-- IPFS_FILES : alt_sv_gx_latopt_x3.vho
-- RELATED_FILES: alt_sv_gx_latopt_x3.vhd, altera_xcvr_functions.sv, sv_pcs.sv, sv_pcs_ch.sv, sv_pma.sv, sv_reconfig_bundle_to_xcvr.sv, sv_reconfig_bundle_to_ip.sv, sv_reconfig_bundle_merger.sv, sv_rx_pma.sv, sv_tx_pma.sv, sv_tx_pma_ch.sv, sv_xcvr_h.sv, sv_xcvr_avmm_csr.sv, sv_xcvr_avmm_dcd.sv, sv_xcvr_avmm.sv, sv_xcvr_data_adapter.sv, sv_xcvr_native.sv, sv_xcvr_plls.sv, alt_xcvr_resync.sv, sv_hssi_10g_rx_pcs_rbc.sv, sv_hssi_10g_tx_pcs_rbc.sv, sv_hssi_8g_rx_pcs_rbc.sv, sv_hssi_8g_tx_pcs_rbc.sv, sv_hssi_8g_pcs_aggregate_rbc.sv, sv_hssi_common_pcs_pma_interface_rbc.sv, sv_hssi_common_pld_pcs_interface_rbc.sv, sv_hssi_pipe_gen1_2_rbc.sv, sv_hssi_pipe_gen3_rbc.sv, sv_hssi_rx_pcs_pma_interface_rbc.sv, sv_hssi_rx_pld_pcs_interface_rbc.sv, sv_hssi_tx_pcs_pma_interface_rbc.sv, sv_hssi_tx_pld_pcs_interface_rbc.sv, altera_xcvr_native_sv_functions_h.sv, altera_xcvr_native_sv.sv
