// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 14:01:27 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
jrpXJkQulR7naEsXxHpqe3wrPuvhDWFJZLYSSLrDAqh5zQ3IMbgyCMiyqZWhFzOb
0UOctaUz1iyHj0GqYn2Nt9nDZSz1bt36EHn1xhUG42UwJ4k1sBRw6WLUzymGF8Bn
aMBJ0CEUuxiDZL2zG8Wt6BqaATiB4luO0l9vAGXogyk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5664)
DJRMR0xp9CgfcIGSW+zBALOvVhWEzEj3u6o85f+hiKb9EEijaY1WJRaOIznk9yrf
AKC+JP2pqlVYWN7bM/5KwEsqG3cLAKt+zpslY3W/lvl004Me+NoG+LxVjKM/J6ms
pQWXr/nKnpQpKblphhlzG9L0tKr/TPHU/Gg2n9oaRHrs6aEqKpVFfELVEUmnvCK3
FAUc2KTZOVsWBtNCGItS3Al9okjwKrrAOjEcMa4irQDM5NEPkyg45r4mI2HfR0+a
vX2RKs5HEXxwcPnw2VXkfRMkXT6jS+/naErKwMaZ57recLwo+Y8YS4s/Xv9KyFYE
VsVd88TVg+olqlA0/cuFuE6iIcf5fmz4Mi75+IWjE68MaAhX4bIe8/97bA8ThGAX
Xb0jbHTHkqKa35Rzfw8UYBk7bfnt/wOourMIf6nMWU7+9RYf70y2TX929xo3rUJk
/egMXOGPp7OhlzDuc6znZ1xeQ1l6/DJ4VHS3chRYt2vlalF5nTuRp6FFcyIM7TK9
ujPzsDmEZOyImdEb9pd131GgBLlg95bsaFuQxbRl4GLbN9VQiR0uEvlOsFakkUip
OMqIWpuMHTOM0jg7QTKQeuPO+3ohUAq+DMZRAlbDpa8jX36iJeJXvBbjM/Vv2D0B
LeYBl+L11fi5qtPuEXxId0BeZWMPPNehmxUF3Mu780LGaUCHPm3THLltMHBKGpVZ
tT5K1T8Dhwls8mRUdo1Ye+iUqk9H029ZuYCR/xKwwEPb03+NypVm9KDZiydqkZSe
RdErYdz1YFDxtXHb06FhyX6nkISgMlGDmRRW6ifZg+TBkOZ3V8E8BeXLD2w+7H8o
ejLXqYLPYmUifJHc6vd855fT07QTRTODONH9W/FLvJUs09MJRz8Mzju7DbwpQR5M
wUHPlvRcokcQjlbms5m6lam+LAnijX9ufuDDIud16KVOfZCUJmyKU2cwCI37ZXyb
sl9kapc680aYmO4w2EdU01FtOZt7qyekoEn1pHl69OTCWFxCD7UOoYwuQy8AbFC9
DqzsBVqkAX0VWgHCStYSyB+7OTNL8OjJ/z4m63ngljo8fDI5fcsQEBz/fw4w6xvE
V2SZ8EFv7hXIpogQJYIhyoPgz3aEFBtaDLnEIpg7zr4AGySHZv2JYDXQU0cq9zEC
mWUlYh565CmcX41tJWS1z9Zn3DpU1sFQ0a4UVrsgeiEj3qJ1Uc6BPuUZjEaGeSEW
76XbsuZbrDD443Vx8d4/+qlNxC/HRmsD7kXzoLd4zoJW79WafALktx9AtqWnzOwn
KY8/Or2znGmkEhE+eOy/aoQ4LKnYV8tVA3ocvF/uHxKNdJ4c7FowXu1LBmczr4N1
CkUWVYCXZxt92Te3lVSDKPZhEM19dxHgEG4UGTRKpPhy9XYmRXit/pQpOjqL1W19
UnMIzWDraE93cDzPNrRvTtHa2BIFFKU2ziVgFvF96ZRiZCwRV3yTaScpJbNPu+2N
qrTKWkenzSmoulpjgpHac9KbEShTHCFICuds74+7KFglfuMkBtmt1vYDYMH13ZCX
1CzGY55Ip47pFhiEntXfWHQ4II1tIk6Vj1OonooyifSfXHWrOYB1R5wCJvwxKPgn
udaycN3H+n70eu4ExBqtc10RgNlhTllPey3yWa/VoetqIpmRNwXM3RKFqy4lsgm9
6Ha6H1iYqo4rIitKXhc6Uzf/bVEqjJQqx9VTOsgBOIcBfXtCnUDmSuC8KZ3okuSP
TyBa0PiAo7fIkRVGNMwXXqmAAH8Y8+SWNCtihTC3XkWAFYLJ989yk7nOm+fPghIv
gYt9p1/5D5RwqyKrcODlAACQd3RyAsiLhH+5tcHjvYCWtF6r/ddK8/goi2ENJVF0
1wcJ2xCfTdbfF3e6GkfGeSFG0CMR2ltgF1ByCLjwH8a8cqSDrvtTh+lzvlmL42c4
Qg3dhhNzgvt8DBXk6AncgLVKyqLPF18jXpTiQSfAGTPFvNT9LuvNpPl0N6bKemEh
oj/eLv/ECywS4X3XEi5qxSCaxl96Vzoly/F/nZAZDjtNDEadeh6qqGjBr0J2nUpk
ZFtj9236GCxOsZZrX6fdxWeX2Tbb5wCpDLKhjUsA4GkbvOG0mtVWQYRp7wEmVXUy
WR1/18uKPNmNjLWSqj0ZDiLz8r9yWqt9RvGUOttS07fXgBn4r4jFk/pWZt+ZKqXo
xb53heGXG4NmDWIkIYBKmGE8Wh4McuH/UHne+I4eA4fe+ELpidaS9LjakbE9nhTD
9CP9DPGKmCmBg9EAfkWUp0E4DsYCo6kxE1HGx2VgOhqJFWCPhEh94bmsRCgBIvCo
VBSmb/86qiOkgp0evqWzGT/5q5AJ5hjdqKGxXnDUKH1oRsj/lY8+sgUTqf4JBRk2
/t9XoSk3ugEKJdoQklbWluq1YexcRONKH2TXwU54iajdi3D+nFToVJqNLrcwWai/
nZgRZxYhqnl8CZJRX6bDdbJUeCjxrNkFqQNls6K9LXoTQKgpi+aQazBCbJmx304W
VfwpKrb4HYiIKk3/a27HL+fU4xPeFSmzMXvQwnUQJOJsJN7v9UHtnzuUpONHGBi/
YxUCo4i+oSxY5bu8ZlorzpEq1CgWF/o2DmBh2TrCFDPkdnrxu55f1sMJY1+JiX8Q
mLE8Czy5zVy09oOfbzMFxl5o4DbVGDSBVRaKAEp1w6YUveoDLRBFKhIRxjkdIIhc
M7BTn62Z71NwB7H2p0GEv2LuMgfCzndfc8Lt+eW5nO7FGm6l5LY/+vXeZv92mutT
T7aVFXr5LWbuY+CUW6reXX/Pi9Vk9o/hKMsFXDMjLRj1m9MbrYqX832EznSuaGxh
UpgYifhbSzj367OIbtU7WtLUXm+pf6w2nAI5wplMQc8lmGjVdYIMjiAvk5/+Of0L
/K0rMMf0GOLROVrsk7vxA5jXQ+H7+s2XYfVmvBV1xm4Gw+wew3Tt2Pt5KDgFhkSp
wyf0lsS+HYzM3bdt5anUMUB/8mKUjhfeByFkHgOKvVQrkiAcOrxG6qLTemgcbYaY
QXeh6+9hdl5eCqSuXv5nsHMwzXs0T/qSmxvOc+9KF7D+TfN6+ek9533HsoTMUUqh
hey3Ns1b5I4jU6d1nEKPxiNBncAklh/BLSNhh8+AXqAAS+hYeq7wdaoMHMBKjOE3
bOxxDQevO8RTchviG7jCjItGcclW64aYzT1AyKPNP5E+qixRQvDINpwIqxlPsuaT
r2NU+WoTKZR64zlSqDW6+2NUS3p5RBJGukKmfsIsrAC9JmbIKRnrz0vo/Ye+abN8
n8rFSAjCiN+Zlartc9LvXuEqey5LMAZnsp0HSqptK6xqGNcGl5BWu3hDoD2HMsl+
KkXXWJs63GUTU8joC0RG0czvEhSAkEvBELgoU35OOeodTnfw20RAwhFNHl3E9Rtf
pGvqe8KTVpNdgDZzB8j4c6aKyUm//Fg6EUmwbeo1hIy/N9XIaK5FEDP96+k2zIwz
MjnDdA/o0bOKSO8Paw0iDqrWkfr/KHgxKhNkKYaGpmM5NTdWBJ2ch6gucyhdUkXa
ueEEM8e4ZNXp/D/q6iCryGFMahHhIjDX6cqua/uFivXKTUvuWZTTgszm4YsJKdyp
tMi3Fo81V9eboRnUfF6pnsCywsYDYdVhrJPYBbGtm+ABmDMskDi2fWx4AQkN9Z91
nxlPNj8BFWymWAi1GxS5/1is6ouBtpN+XnOIAGq2plFmOVYtrZeD72NTzZvu6PEb
+l+Wb/+b2YH4ClieS6gt3IOLPztuhwyduHb4DzVDXm35erYCEhmyEhCRy4UDhzr+
LwSduUf7QAAv+WnMj+lunTx/gTDBERy6mSYKgGCmLsLGpjJfhtvBquWN9do4MetL
TU67m9q4vqOklgTyejhWRqtGmC9OwQ0k/HP8vKxuU/FFYC2a3DQYgLxdr8PrTbKK
bwcP7yBIs/pJ5fehzzfIgBJjSokXYy4GGRfVAM6FkU+3auZGJsHQ7G4/A4tGSfBC
QdCQqQgM7io4o2NprO5AUBLrbWkzQTUAHn0lPKtVsIe/29p39uSE/4eeJys1y2Ka
RDjHEMAVyZp42l0InhzxFUdl9d0A4AsQIzqZTltP0fNT0GX9cACsqk28MqRpIABd
Ibl0YlUGCFI1+uS/QpV8QAK9DuxnmTVuZ3i5qu0CmAAVAsiPKz2PBFqOAQDg6hhE
BEYMii2BdhdNx2tXxtpH4bww5N3pX7HJIl/YStrXvh40kvOGZBxNzcJFefR2SqLX
38x/9qG6/I3UOXp+txzKBRnABVBvQrNVlGqPU8NXocVVdRkhgcX9t9o0Sf/yMfOt
S2swMk5kd57iTVHW4dNzTzzSgbdQnBFWoLF3dqT5iVMF2WPOVjFYyXgff1uAURZb
jJJY5vFt1pi8pinLKN3WNxQiwZKyF6D+Knke0UQk4SJn1izhW2Pi2RWwPkUezxyb
iHZToVWRbIAV4mJIr/Cq2HLPl/M3tOfimCIK/Q0bicPDekYf+3NdHPJXRDoAPWtk
GZb2i4siX/OZwFSAd4Zwwr6WViTN5AkcGqibOAI1Gnohx+/3eDCxrmam/MFomhZs
Z7Ldthj3hktzQ25Gd9L1VgsV4KOOBjz7MngY5EZ9FVpoyKDyEQtzk/w7+FSX+c+C
f0dsZjEy6WEY2EXOkTawhFOxY4jA9LCOj/1GhlkVzadCVHRFxFAz/6mWyFzErWja
aMCMDuV012M8JHlJzxvEd04qKUUoiLPJsvbeGHAfYN82texG2jKMGruWMnCIq+Qq
W0onRCUJXzFjHu6MK35ed6CPMJ4kVaA7Bn1UdkyWq89gssheSrL3axBI2sn1FTgg
85YlpVsrJNr8HUtYgjjrDtVouReWdxKR3kuN8s38rjObfnyJU9750e+Uklxolbgg
6rLH1ScTgJf3EKHbq/YC3UHBFzppWHwZu6B794UZg2VpqbTKwqEWJqSaSCBuSA2J
a9XT75DDo+X79hdBr5kKWn+LU1r7trtbyuE5f178kWqAeE87Y7RWP0wlEs19QCE0
nhvWb7VNR1UZefQiHZxh2rVwF2QCtzkB3h1xf2jbhtfdirGDKaKBJAFVQ4xXfoS1
cqvZ9fjA0DUEa8cKj61jqxFIvbXVtAdeuK4CHMqzxTdv5BMRjo9UeaOgiGRxSCaS
EkJC4x1/h2FsvFbKr084PqnbmQX20r2//RHYgib8fr3Qsei6KCkI0GRvsE7VXXzL
0IV90s8RlQH7ZxiWrihGhGgZ9aROKQZjsntmVux2uplMfvboye8wXfkGXlJ4zaEs
vVsw2sMJbNoJD/Yq/et/ffyzknXtrBfTukVqlHxeJysiuzsnfSubsswiN28+H3bx
rAB4H+K9QbVTtE67CxcwJ7sIO5c5HJa9nVZolAUOdHG8TllHzI/WPCW6dj1S++Y2
xT13PzgMzcbGb0zrZ7GQFlG6sQ8kTzOmU7mEENreWO7q153Z38GBMnTSHQ+qQYnc
hzgv1PYupaJrACTjDOK0kwtJRbplCLMqf53kFfphEgvEiinhcytVcKSfISQB4gla
2JNuXNOo/3GOi+cheXZ87vH127sdEIwFM5JzyhabuUEAYprdtbUUkKL8IXd7Z8se
MOhaZw6RaBJJJNXWQpmQMCPpRg0zQZqBTYyT9PD2IvdRnZ6TF3hv6mj+pxlMx9E8
UoQJ8KJMyuJRe25RhUA9D8yHoXLq4JPAnz+r+IPoRpjSPRpV3k1G1TN4hxSp29q+
RXEVj1IYDis0wJRDVkDPXdlRo/uRn0oMaTH+/GHhShZ1yt7YQDDn6UjG57Pvw+Et
9hPdYP5kGgsGEGGNP5Zo9zvU4G1xBp8cY8FoUyY7TS7MMx56PGcPKTecthC0dp9I
wBthz5ikwPlYeAzaQm+EVDpk0Ai3BUjd6Ts6g+bCgyesDSsDl1iuDMpLT21Aunyu
X2AOXMqfxCNhSJm7COpqUSlnw/jd2XnnwXncBD+LUcwYrVqT86+Iv0wfCO/VGNbj
qvAmEBMCbfSva2i2z/zSrpMYU8dQqYSpxu8Xa3Ynobo6qdekE1h0cLCOS2T+RMh0
cUecC6gdGXHbneyAje3ITEkUWTRNbc0nJycklAYXHgi/qMZcW8rjRlV7iZ9xfUAy
ameX0dGNBSw3Nnih7E2goL5aff/IkaFXx1iboQOd2eZGoeyDww8RZG4ExuK8L3HP
bA410V+QA8GoscGheb+DzFoc7GG3WLtFWIndt9v4yR3ZU43TzVgC1MQ/WhlwrG6F
e+sgRvFu22CPJk06ZAuy/vaJ4NcqBLAw/JobuNRfcCPrX+w+bMfDh1NvR5JjH9Io
iSHHQMzHPo/M4qNeu9r66cO4yK1xCGt0ciCDrOY6YmXwWzi9e0IrhlHEGI2CW573
kfcWkQ6SFec2bwYcnFf48Ix81K6dpgNDxAtPMFEnm4RGjcjNT9DLgfrk/YJPmF/+
U1HVgD/WxeRFCcQ8Z6MllpgHUxRg1npDYSfdWJF/jod+/Hkuv9bb7X5lyvbA2eNK
y2awbavz3L260tuxdGZ1qmPMJEwY+QZq6yEvPWKXXGo35xOpOocY3HFPOgmr+Z00
rsOuKXiVjW/w/wdD3csCj5Amo6CUEBoQbAJORv/Sydryp1OCDmC/0KHj1BMFMxV+
79Vzf56A9ovbxb7ZrngqKCVnRHM2SGLDYSgCxCQvhDt0uLHAxmuC3th7KPhMs6rX
pLCCBpf+qVfI15lJaV83xZQmdMBivUIDZR1JoFRq4WyGFFHQkInmxpoR16vVsMYy
ZDzJEXYY+g6sjgy+AzUID+zvDzltNt1DYaBRcU3flBEHu76wqwzEozYrXaaQLxai
MF3oFy8I95SKpCpYaKh3Z2q5znqneRNqcSge1IxwrGow8/26/CFJpEVcw9Kb1Lhb
FcZJDgmjd5MTwvhRPGHK0N3KVwpdz3Wbq49i+3OdadO0GzrmwcNeczEryQC5OPZ/
xLR8lXxzdrN1UpobQGz5SMZKn6b/Lj5L/nx9MVD8eO0QpksKUNQI/JLDSu/Zd/Rc
f7UjIOvfAGw7Y64ieggOairC769N7afYduhLthh14zrYXIc+y2abdzRX/MFQJ2Rh
tiEgi4w+ilvCJVxTLSv8SoQhQOub6hRB+17QAl+cefpxE3Xl5cfrb2Iv0Vctuoob
U5JN6ITNs1yXOdbkv9Gn1f/r/0cdjHG/ZRKGLLQKZE3rPe8TqEvEePX1gx4oJZIp
zfml7igjaXxVNs/iICx+Z2vGUTHnQwfZzg/E5Zrlj7dOlG45AQCe6hyX0j1WpXkF
gtg8Q8k0pFMb6W4VMcTaFqMQPuPEjSQavzJvVU5xfa3yXhMj28oE2sZfKEL7Vuku
CFczzOyrtlQhd2V3CP+3v7zPp52+aSzoKXBVIMohSMaoZDwg9FMiDvNdNM0+aiNn
uQ5trEjrm+/jEBkwz+L4Ne6h4BtiO34W8TNkkYscbgm5o1QJAqzxF34CPlDFhrzE
BUcBgSy1YDHTlmgsvyGLR7DJunoXKCIRT+k0WZq4Lfxj0fWUbIToJ9Vb3/tBegbX
2IRjkjfhRsT4FhXoWUnYkZwo7MIorcMo+KvRLizKL0F6s7MFV4kAQXJYeXcZUIYA
`pragma protect end_protected
