// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:02:16 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
O/KSqC2QdUy17j2OC+oFOh+ipkPCgvAtPtKrVIkcFkR1nv8kBXIThfHTRVg9b5IR
5kTQjmotTLrb1uI04hYeKAcS0BjhhV+PFiaM0ztEuwuU3AWgd5ZBVPmNIoeOO/lg
tOX+fpt3gi6D646Lc+rn+mL3wcRsZ5NjQYArJHTHuQI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 183296)
56YbENbh2iALOBQedwCpfHBwIR3lHBV1SogsE+yOYXDB8ji9YJj73srqZJ0zGk1c
Q8FP9Br1MBW7iOTS2GiLDruAUnXVwDbc/6jYoFmjYH7Gmyhuhl3ISIhtsO2k8lBA
Ib4TPsm9lzaEy3t8j6zUun1YuqLHryh639wTh9LwbrSrwN24OLvnIWGUNspY5hoq
ctwWk2oquoPcjPVEL7gXCUw/wmxaSYP3cgIEs7PYvCziOIC/STtrO89YpqRqVSx2
ZdfueDEJJbPDYwgfH4YNw3lKcX6TYy/yhg+JwzSm32+1HgNQ1PjtFayVRdmQcBo/
UIif7xTP9zDmNK7lX7mrkb4ek5jhh0E83tKuSbpwzKywOaHFwEUyN/3trbqtd8GH
YsfgWrcPDzRyaw7OlSIbT/ApLA4gBRIT8xoTF1EcuzkET4lDdXe90KoK9tDJ0Gf0
Q5WZQGwtlR2l2GGi72EbdTUEskNUB26sUt7A5YEVSONWO1HHU+s5XIofBy8JdTrt
Z2odJES861shHJOXBoP02HlQG/gqFDbLTNT140mnQlh06k549ULce8qk7oZMHzTt
PpssfOgVg+c/PQBw3v5okBxKLxMYRURMqYeUwRz8d6+Q95Wf3rH8ZRxQEy6dlPIe
6e4w6p1xPudzELZoVkJIF0K1dayzmovAAtE3T1r2gvdKC7Gc6Wk+CG99yXk9j30h
8IGKHbTiRi7B8amzKbdZHoTDXdqqmZwTZVIQQln5ZfRqN62X6FyBwvj4LsYznw6E
hWoDSRxM1WPN9s0MHsDpDkU2LVa445aJC5n+fTwqnhPks3oISeg86JsdSmdvAIYV
RUw5f4peJ2ORiNT8jI7RZvNmsdBfMyYmXE5fDDIjSLepDI3UMQJcjG9LQw6D8z8x
NsOmCgU8cARENSDBdKGIu8W1ENqpV7xI0cY33FJdICXqytWAXn20j/XRJ5LH3sIV
pIkkJXoOzfIvTdVK0QdPVWAO7Ck4VRpNL2OijKTteFIhLJB7dOWQu3Lmh6+7ivrf
G8u1KePi6d0YpNw2DA3+1QespxURz/53kA0iDp9VqJWmsX+fu22ukg2IlIBUsz3P
TbPl/MKsTsPmSiolu4EcbcW77ZEMbC0CYyqjzWuq17I11J43ntUMrSEtvGI+fXPy
MMtGtTS4+AViHAdPJl4ANCkX1PBvTJmJPsbbggUlpcFbBldi9OpD6Mv8qC2jH5Qq
TonqjoOXd3oPbN8021GNHtHEQRpk4nQ4WlsD1bc5oUB2VXEF+/c9cNMwBiCUBmeX
ZY5pE1DGzDI/WOLx/w5UMqqjGGXT09Anfyoz+RWVwbi3zPs21oOGWuna0cJstU1c
+Wg65QQ+SjIFsovHFb2+Dhs1Mx+XorTbiC3PrYqB2DCExySMufjpE+u+M5j51TuX
Ge8Csf4JIxBoXMt+lGaiBJrUJzUwmNFi177WbM8R8CvjJZYT8LhbJ4bAnlfB1N8P
cZcE/ZwHmcw8Mf3bTH/uUIjHm1jEfh5ovRQPHk6Jn/URqDZEchxe3CMiL1sJ8Cs8
Fijjw1U/mj54I8o/c0LcXDsU64MwzECPrmIUHlzxdvtJgrnqaZyen1tCKiNaxkQF
2DzhfWAncKGF7jRzOPNlnkfYhQokGTABRYeJmz8uSFGSjRrNiDaQd9vyIAdvzFki
2i93NAXhDN6XFWd8It37hry+DycqKsrcHBjIY4WPD0A6SMgAJi+V0MX+pplEELaB
6UemDDQt7jlxXKd1E0cWFoA71+31eCNe95q2rf+xiHiIdKdALzVkJuL3u3NEVNq6
geWApokMRSs18xo4qv9pu8cZ9MjKpYNSEFHUp8ZbgtD7LxZ5VWi4TZhBqvWnlA9K
qPlfoDcPMQM/uspDYJ6+pO1NutDL3JdrbapnCFaGvlOhcCE7fU5C4Nx8ZzIGlBeG
d4fBI3WV+drcTtTFaq5BGjzQ3Rl+eFRCkzyvyVgdtnCkVCdOQCag1W+MVBYqU5vc
4GF0ka5a+ZLZIWVMBMfl2Bjg9VXMY6nxJyiNL5fmTj4lEZHwDdSbcR6INOb2FpTF
qh/2Zr3S7C2r5oa1JmTd2iu4Umvs3K+oQz972IWFouPsmMy8tzQNN+60NR58ni7Z
nfnS6IsNISzKAF4w+no3YVIfxJWLVGTBpo7a0OuUFNpM1AmdPaWpivblMGkIXG2n
aizp/RnWmycqh9iiRgURXZloe7CzAat7AO2om4k1gnI9wWqaUIOhYz7jqBTvKYw4
+z+LYye9WKqREzbF8QV5T1HBZcngFVYHV5Q1M6lKlWQys0ingLOgOm1/br7KWqJu
FrQCQCiAT4xYkt9mn5r2Py+EDlQ2VFhw0yS9rn7NsN1smY+hxZIzLteLGGStcGhC
WKLhSsv1Jy1NtSPThW6boT5jFaYvpRe/qPLvUOkm8sGxbsfdFhkT4nhsfkqreQPB
Ed2F2fRD+NgE09kTEgsUG483zeiXpQ4lgfobPrkovRPCEnoLfQDWr8lhjbjodsMy
VhvLgZQkaU/AJm6XL18Bk0dZjNKtiR5In2J9kihtDtZgitJyUv/QgAL9J/4bCKcC
F6EAw7BEwHz2vnIAZvL/LQn++KFHFtBAQ9B2RHO5JLOhwUh+bsV8GaW81piGXr79
VdEbqS0dDajGqMLGa0y1rsxILN7QVAXIMVc3RHlzyAehBdJXENR0Z1WbnlSIxBHc
Pj02KW2HNuhFKUkoWzBFJ577zMuZ1QWMAoacC2X3uxCVNpK84g73plLLc2iezwqC
AjxTQDimAtuXcSl24ow6lC6SZciInXxdXi6tnON3wk/Ryt4VxHw2bmjLzeOVIrC4
SA0O1NhzxKeTJ4pY4oNYY85CkinXgjfaQzTGMQdn28zKkuljXaSq+BwejC47Nm6e
28Q8jME4G2gz0D3H07cpSzeJcgn4i/KNQi+PTigSK4uMW6lg/0YxIUiZFFQdRI9B
GGKsPs4TuGVJcbB6TdUk1QEsCQilXU/P8xoYm7JF+gW2K1QGrl1kJMJju4OiquG1
BMbh7mSQUHccHFUVRuiXXrlI4NkrwUXpl+FtqwpYlBlmV5UiEgkkuRUeWmf6clYK
QDKgBxncZl+WjU8qGgggVweXZ8f3Ec3dwJ6XOWkPVGDuqFUqBBolBDj0vqo5/kxI
XGnPR0lbvP1bjLAcopLKdr0u2G8cc0rc3QTeoLdQMUx2WXVTNzON3xOSPqKZQID5
GIvjW0ku8myXAxG6L9Zp3M7UGKcBPvrCMZbRo6KR71KDEGJlfl96QXiYE7hXAHB4
u8uSWoZR9ipgQEPHGlT8MUP/oJ6Qtstj15M7PmDysb/MDMH+NC5NnXPJi24HhIw9
+B78Esea1jVyHd8uKLMjKGHutePGAgRzCWNr1wycZd/hlZX5rRuNEaOOp0jiNyFv
X13GCpE8KqWD6Yp69imK7MIgSzsc009NNvY90NkpXfAoJAhWp9UiY3DddxY7H/Vx
8x9YOWPiAfRPW17FhHx8MCxtrZBZYxrcIOJeyydGbk2jGPOUYO150FtROZdpJ//5
hfHQgNLq1r2ujWytm3JzpoDEV7Rzf8WfaL+4dNwV0oTIvGH4xikF0bwSeQINT6cK
hQsWaEoSQ6RMyBkcM7wk9Pn8VtBlSjSTcaUJ9akEu5KbJeDieMf4u5l5QYeRwoOz
SvXgI6Nv9Ta+/6nFeyN27XZBnLCK+BeEqsT2AegiN75YrHzTmR5zOl3+ZO7A2Smh
WWAzkk8q+COEo84mhdl7EqG6BC0xMnXBp52/UIkW/OyMYqN5QG6dOlpm8ybhLcbe
I81RKJ+s67illZNrRKGxlyN0pnabaAFuU++UKSGFj5qSP0V7rFRCcJy9BrmFV4ux
ge20UGrDkEgBKg3wyzyGuLFmgefocXv1glJ4uKTyehi/ey17rhmx34ABkFmiTj2l
Mi7/QskLqphEuTSk4malNFvWqlUN2tXnQvcYgNPNiRiKLKUHOb3MiPWtnUguibnz
IAiD/K1qsDGWkG0NlvJFJLS9z+w955ZqvdBcqHhs0JLOs8Y8blLe6y3QFmddfrKE
QHi3YoOCU0vc8bIQpH1Vx2fEv/aHiSGuGtQh3NeYnymS/FY4qwJDj4znfx14n0Vh
YxP/kay1VaKvt+cQ1t8SKXIXrd/nMTee/ZHAM32qBiZIBimUvpIj0/tSgXadCPcw
RsUGoJamHGSNB9ILkb4/lWucwc6X9jxR62DmIog56ELMBjrDFAakVCQyoPr7Dnd5
sxOX3yT38KdQMEZtcz54O0roXKP9dfsvOp8NbiROG7kfv5S5gNjWsA4+AhKr0rYo
dtq4ghnB467pIEkdm6VzVYJE3rFxmvkhlUBQTW6tPZOxKhySFaV9Y+QgyFdjE3Yi
Att964ZYrsCQ33PqaKx5WuymafVjDuAAjrot+78wAv3JnvKBMgcCHdv8nPuRi+Xk
GJ5DdmaWonO87XlYM3xuHz7JjF/qtkC+ce74i7OETE1HBSclnMup2aG1LfngvYVI
dm12QbGwgxDvUUSCGNOveXUIF/V0/vTTOrNShg6jWZx11e4mOAySqsG0cArjJBSs
InRrndDYO8r56rfxCjjv9hfeKzeR716kI3SA5JLSDCShz/1QRJCILoEU74mofpMK
+7oXvf3tjNUtZFoOUy3f5/cQARIhhTJl4Z2M5tPLZutVU8hPKdQjJ/XjUwi09Mc9
appODJ4XXX0XNGecv4Yak+lgTsA/WjsckMD5mpT25NqEIm96ZleHayueSZP33pWb
vDp4vx0xGtyXJj4TBRVA/AuhWYE5zuAasRRujJDvzCcYL+FUliVp6z2Mn1bf8tFf
KovSnTOmf6RC7PVIy6DiH0lFztFL3u3foT5k/rAns7MhraqRsDIMDSsC8BJ3YRpB
WUwiHCRFvn7jxhnTuVHN8hWegk+5J9K4st9qOl6pHlRTb3Eeb+Mvkvno7+1RfbQc
HtWrmSyRl7+j5IPIQjqczU77v6YH/6vGP37KT3tdkGo0pQ/TJw1NZHqCgtNGaE3g
dcPbV0vwEeq+YVwbQHq5HG+oj8iAW5lv4fggj4nDviApCdMg1OK8lNNzTesSb8wy
L22VXkgFFu26aZ7Ix1mJDz/ozuaKq1n8dKsLhnGe/XlzYyH+p9BOku3CXYY/olHp
73IO7412Vpt8foiwVdCP3BeF7Uq8zDIX1Jy5vEJoG+CvwB8J40OPTsjcBnpVou95
9zcWK5ijPbBiRIs+UOIKjkHtRvo068Jgwoo83eQiqGzO8jhb1is0BnZyRVIiLwVb
jv6/DXuacVw4ifyeB+oQYTsqec9+msKA+V0NuMg/MVqB4sywAY7o9Vdip/6NtcNl
ODgXimmQlSVc3sIgm9d8TBK9qZQcI0nXyaCATO60F0glvWLUqvU2T98Bzf89KJ1v
uewA39Kmq5RHiNDanKuaqWBrjuuLPGFLYn8Fr/4fVOvQIXdKNP2dOW5jsV9u/4Qn
/eb1/CRwshgMMU53IW3gqry9Yg2KWjSS+Rc4WzgJiGRzYTs6outppl7omWSHtZDK
eSHiogUTet2pnW+sAakburl+Bu4w9Szr9cRgsBgI0Vei2jklRov1B20gG3i3KTnD
IuUKGjCR1uo2D0fA6PDSgT6Ojqrd1T6iRXvan5qNsIDYbaZyG9xS7EPiHg0Eg+qG
7l3zedy7M1p2dBOaCY0k/QcHdxSaf3i9Wl7AlEMMBO4cQZeakxSJ1NK7KTl/IaLk
hijHHFgMNM7h5eIukBQuz7iTe4GIKzvGBEe6nqOS1wNJG/KRhO2bjpp1AW+qe0ny
aL3prFJOGKYgnizZ4BeB+rXlgdAC5l5qCXjkW7FCCjnXeD2gzi1rdx8mFeEcZvkY
63zA6uIFKhvHm4lMDVHT837ALotXKHaq0GaF5ebMg0MxrcARF+Vo+AZ5RltmpuwO
mUrCWddnnv1fomd/rVUNqSjDHuJJS+RldnwpT2Xeta3Wbq9ZU6O5yBlpVwBj52mB
SwHuOniuHnznhOQHgb+4X/0hW5+Cn/vk8DtEio4m8b5CNaf60pK4CFrseGpciRjN
t1EuXsoQbVR63S2VsOkemt4Ql3bbNdYdHd+8sfz0eOmt3FbSJJ6iymunmgtb1LG5
jk71u5iFQBlyE9UmjZERT0zx8L1SK/7z6vAvX8+27+COSi/0KOqgfMMvQv5w6tV5
4pb/wT/SBscoYLmBsqm+VZ/8xdlRI8TkEytphs5B/0LA/CWYKO7wtxDYiOJmGLFI
XHpr6uTvFRTOmXiv6Z1ekJwz9i1wD59kTQPuo8QmTOPIsgVXYWjoddt2Xc0/B/l+
7Bx9NLVyi2SJWxoljFaU2iKgoRX/lRrGJmdSD+RaLeL616CJT0v9dapQUzWd/kPr
EcZo2ZvKpJnxnTrdpwXPrmdvwCnOlv5hsOLaPcyK4I95PlOKXz/Ev0jgoquZCjKF
YlEl1wnHhE6n8x8k2oLu25Cyd/nqkFWOJa8iVrY7hKTgV+kLGeS/jIFC9F/v5XVF
z8Y74iHg09xMQ/1wUmE29QrD9dApOdeibPQK9PidcClydOpvGqM8Ttz+R64DWbxX
m2cYBw73/kHSDNK+BMHvYo4G6c7xvgp6Z4Sia18imLY+mmsINnNANNNoATyBSBrx
vxjRGGx4rexy4bCvV6PATC/l0J25mIoomSJRhF4+c8SLV+awolfDglJZ6VsuHWXQ
CXHWOvKSeT2dViVmUi5NaEtEjr9oXLwwKU7fRalvleGy0Syly9fef4F47YQxuIKi
GJLUfzdMLqGkylB+6FTx0lGKAS6qcfOLoBQRi6yAlK3jOg8f1awY+cmmXN2JS3DE
Sbypifvf+25vdeqcha51A4LNe1Bg/nDTJ9XTzdFomA/EiAGpb/aSXJBlrs8S06WH
EAx5xiiCIqlQr+FiHJA4ki9qLp3yNrj1ZFXz1PppziMkS8dUJUaeBvfJsRCHYddz
N2aB3MMg+DjuYsDlTvr07IXyLfljNsCyKgCxQn02ILYHAvTqsDGLBwVZWq2GHmzk
+/bKQYUOiUayZz2pqwn4BNJZNyWVN6NHd0JV+QICVcQ1XNVDVPsU0C1543NmjHR5
wyO7Y4XjI7nNqnOHLk8vPcEIyyU6l6AvXp2njr0kI/6BKRlJWN126/bGOSPC4exB
Fc53KleTd33T4PNTsKyWMfiCu8Mv3LPFTkV4nF8O1lrwxyFFgfx2glOfM77ciz5q
lE3EoDnurpXIHq+z/y72baB4VufdgLI61E3/yCeMGQ1pomlqeuCQOWyrF/ffBITL
1D2rUkSd4P5cjAIqhDgW7prp2VfvnVbzkqtCVZtGaQdUj0WkEKUouxsrm4CabBTV
O00c41n6mz9E+SpacH6waMl4QlP/SOGs6yqLjYft3jCZ3SWz9pH8jIZsvn0A8Ixd
J1VBCbR2yAmPzrBoHg+cHgJ9p0htVO5qb5qTOsEyOZKP05Oel4yeTrLoDn+UeCAc
2lhZ6uiICy+dR+GJMhg35TqVdbvmEKxiXnNOfeWfwXVAssYqGEphrvSgVm/FPeVE
OvhsfvwKtqVzDkJaSb9nhMS8W/rGdVd2+5jrnKn5XQsQN4PxpYqwJQYN4dJEmLRj
XTgClvqrzkUD+iVsKFgz64nwMCm+NXPJNZkQamuk3hVRWHcb9Fg4Xxu31KcxA0aj
96AdA1TL/zMA5kt5jWw/yzHmWd/8+OfbgWn3EPOpuzTsPcw9RdfoH/ePmLASRaxn
APg+9JrioXCBFrYdxk/6TviLH3sXjNX7sptWbxLC0NXWL5hx5QPcMOeSmnZFkGt4
GdY/X4UFBTU20D6+3+hv3PEB7wZFtMWzYUywwwJYdpz/9GUSSm8GgNZ0XThmPdRk
h991O3Ld8yzl2g1xhx2Ft1hYPJqCpwRsXHC3WjQz971TBNFpbCFNkHDwGxD5foUq
qtqUYHFnBcrl8HcvdLyMKmrSVp5xBK69Z4Mu/BMWri10UfnS+44Sljtfrp9XSvjr
AOfhF4YYZJJ0ISKPR5zomxFZc8P+repEVYwhrxoFvZbGL2/LwEG5K1FzozBL5/40
poXhPbBvz3RswD918ZbR9uTTC5BnI7oxSTcZCaX3tcmDCn+w2spfZHzsz0fBT0ld
PPZAsRd7mmL1o0JryZOThR09doLybHbxztan64WIs3cR2AeF+N8vLGodZFaKjjzv
/expOFiV4GAtCKrEqZLJBtr/qecvj81i2RpOF4r8KD3r+PvRE7+F4o/N/U0QAGQ/
+wgVip7C0zH8uukFGRIzvvKDdbCfeh03a0igNJP8OFfp77cUXPauVroFhwWeA8MR
scMSANSU3JJ97rHB6nf1vqxMA/12SsZFWiR8Nv/Coobqm1vteMX0nMA565lYD4d/
P6W4B4LADATI7XKGZN/sM25u0hd+Ao5zOfHzrXW9FJXN6k+4uUUtUWVWM2XpuGGr
M2tkehSyPN+YtKsrPpZGxbjGcazqYXMp7nMxPEtBo8cACrl++gR11SBx6bammt6a
h1BNTLiWuCuNf67UiFKNJ/I5/uBq8IRHsxcr6bGWglQ/tz3pCAqa149yWCjf8QyN
/jvhLTlSv796mMY1wSk2+/aJ4D+a8kAOhwmd9QQwLCJYVcPnDaWsCouCE2gmkPhO
B07Btvh6bYDbTDFfSIzjdOvAZuk1KQ/gQAuOi2LYbr09whrWmW1MZ08rC8rAD6R3
tIjlt8bDC3mPRE/ltvmxVHkGQsz/sjYjQeg48fPGWAacAnWLxCoSo49TgH2SO6t6
q8EX1hZwKya26zabSqT0B0scitPR1X0Rz8p8kcmfAla9D+sC2+HMXZwprg2CbWKZ
jrfsPJ7eiBUZEyFHAL1X0n775t5i0Uxgovz6uA3/iLy2cUQAZFqlmcoWxyON1yOv
c1nOK1c1BxT04K/vEFPxkMoshdoYa5iO8bUcOWSeT1cbQNn3gv+8To5JPHtQvUiz
mzy7AdwVOWNzZmBNkbvJRVP34cMHq7mrf6vDsO4uvj5LzPf6kOtDyFHIRH3f5QPa
qHvr/p+kO0vl34IFl7Fi0Im2r1iF5U7k+V6eKNFBBo2Szkub3u5B7t8YMLSaRrlK
45B0jhoaxpIewGcaHru2LTZK7KFBckz+NnI10p2eCQgARVrmfnZojS1gGKmljzze
JnT+I12uqiV5rUpQJ2MOR3BHiXu0LKhoOwajb4s3580qMl8fKPuVOwARCANZ2ZyX
2dQ+vl7dGcxWkdvNt1lC4ORBgVjh1cAEvtbUmjH1x/Dd/oa63LT0CViE/nbpP0Ew
taBPcJsPNxRpe60SxgUbCe/L/iZp/6n2bhYbH9Gyg2xPmh+2qOm/dOrV6cEDEDoF
+AsPGCoHRqJFXw97NnVFN6A5wwfXyH0G6Nh3qgjywy58Cacu6fnnr6wD7Qi170yd
LYP9l1jyLtCoxqwrGOy6Eu1TXQ2zqh30FxeUHpNsGQQxqDVLmQU2VJ0YVxyUN74O
ADFsM1s2duyujX9W5L5p1/nELLca91b7c8LGO/h9LN9+goyJT81bMbl2Xv1nKFUN
Is5xSFQl4hd+hIBEwBiRrG8PuciVNm/6LlLQM/bhizPEi/KpRDlWgdDBSWbhMiZ1
F8c/x11WHBr5HpSuKWmL6fGlJf/DWuoL2JFwdowzoaGBWz9oc2TrXjxlOGrMfGNq
Yhux80Uo9J+Q5jJmNqzd/gXXS9mvLJ3jZF5KccUBHur6v0B6jDi7uOQOqHNlm1jX
JiwGH1O2XJqoj/8L23KsIkFOGOUwbTPaMADNR8ujKNd4ZdF5d7b4iaDK9tIdcxW+
7LaJSSyJ4u/nPrQEPE/QgeOvGDkJQwh1Lr9DHK5QYhahR6w30GpO/rhhn1E3Cx9m
AUn4Iy7GJNbbn9yGE56ZsyQG/DDUmCKfujT39C5jrLOMuPTktngamRyoUpmW87qz
Z7OCWrTSiKCvaWooOY4p0VfaLO+W278tvtrS2Hpbl7Q4OFU3eElrYaSJZ2UygY8w
LItwQ1/xo/Odys159BbAA9umHCZDl8v6s+gtbVsxsU8WdJRxYQPmcdNQANbB6q82
dXq8bKjktqeKIFEYb6U33+Wm4SXLSVMyQsRaAHPprraJPk8QNEqGXDfPNe5CoH5D
ViTtlNYmfed8EPlC/+AiXQYNzwiR5k1Z9hsqO5TwgE0Scga6TkCkQa3z9TYWSwkd
fsvu6L4ncL50UdpH39AwccZUN4uq2OQRv9wSoZch1ooq4ObWep4vqtUzV62xFY9h
+BcEtZUHBOOLSgj+Aqy4F2NKFam//au/Ku+8lOROLg4O7xNqbt/vQBgVwL+KZ1Do
Q69hSN6JsvgbxLmlkLi2xPHbKXuJ/cERA/YoqwxOa/cK00ocEIGHigclIkaFUYm4
yuih28bmJNv3Xq9hpCg4yj9Q/L5tmncIh2U/ud80aKxGGDxDNttPbssG8fKRNab0
wuM3YhS+akI23rGn4E7ViTGiFzvdJwDo1NrFnM2KQh5g73WNvCnGkWVWl9+GMxnK
AF7kPGgfvjloEka80HJNDhiDnyGXXlAF8fNTYD1kUwC7e2r6kRtDq+EM4Y93mUnm
XuaNkQUGqm/qyDbneMUdBwBBtZNlF3+c9HiKjgpQESELN5EsS+OcXOP7lOzHJO5j
tywdfTfcwZuebjMoK5VwFisSRJVZDfasXBbEF4tJflIE1dhKC2kgpWO4FUcFtW0P
3KoCHy7h8M/0+I0MVu7/75+lriEpVtQRKYhWFOG74JnAuuwQfm/gMmWf4WU5GOpn
zvuBCqSJYpEcbaB3O6bHFXccKKPgvUG+Nx4NZ9MinNi6UrvdpZH+SEHZUlLFawDL
k0o1WM+x5ehha3XvGCoc+KsTLJotr1CoVL1J4UhSFJggj+dkU/xVlDY8xk4i49WS
uq+BCPAF6FH2gvvtS5Z+JVFAyUfnBORpGBca/DqXFC23w2wVKUvcsRc472ykrC2/
Iy/O29yotqOcE5cGU2k7tYZexRokbX0my1Wv2W15IhlUjMWJwUFslyBTWShh5Yyb
z1r9WM7YfC3Wm7VcaIHRDyZ4+UsWvYg3aMDkEUrBYoAQXVqQeQESIF+3KHsCbTDA
aCT0V1v0Xc9DANF4JaBqgEf1SshEJPf+JqKDWaHosCB78DtJEoqQUiKIJsrKmMX/
0OlOvCYY3c/7iWYBntbvXhgcL5l+CWVsaidEeOFqNyktsFQYNCt557bQv6LWntJQ
iHFUEDLwFLRqtkBIaxl91dKwUXlL20BsTzBMJJn18tgBEQMZrH6NAKaNEMOjyPdv
ol8RhpMQt0aYFzOq+KR1W0SVCC25IBLRLwQATGfzqfM7BErT3RRf9oWgLfKTbox3
SRi69tbxpHlGIUDcJvOunZV6xHDN9Yu8LldayMd9KbnuKOtmi6r3CWAxSWvfPeAf
IduFeCT+hEKaTYy6rMI9ElaRA8fU+9+13Z7yZrS2HADFUAw1vJMwdFCIOtP3JBhF
YlCLL1CvtcFcCjtTqCK4RrfyKH/a7NOh25ylHrisBBp4G3oHpVcLGvJhGl24NRne
1R7QFp4b0mNxxFctfCo5K7iTFTcxA86gse64WIL+mVY5TgYCEs87pkxyQh43Pgxf
AAJD33KxEbV09qAMeZ1GTCZU925AiQHF7eR+J9XddzDrxtzbrAdaiJarJJ0hLhOv
LrjvAXlyYT3gtfFkbESDPcGHfLRyZPu0ggg/QBujO1KMJS+wzDYvKEjSk0QkYlUi
bRm/CbGJzIs743d+LBJfKTHHaJ2pR5lV+HV4zB/JXS3X7s7hxiEhgYW3D04M4z6Z
gJss1xjsSwpNBmFcZjaeQO1DzN5UwaPjWNxijzIvbwLuiH5E/dHYDNrtVBK9sOc7
jVXDJhkTx6vgJk0s0XKNyd9U6jsXUnq6O2yW6eJGIQ7lJo1+m+2rt7izNDSby4NL
n4iIa8bsIT+2Q8DMJkhsobC396zZH5MfOefTkvOqftUgrmVK9/n/b6xh2q+So0B9
eelcd6+CIp/9Rumg5BPt78L5jLnNJyGaa3dbVzOxTNb8XnqmPpKtx72e9AgmjhTX
991u5P/MToDWeS5NFw/Rs1ZU7QlaOCfDVHry+t1mDgC9hXMDUi4R/Jl3UxlQ5oHx
E+QCgD6Qf3SXR4v16kusBiD2k3YQVJ7lVV4aijIIovcFRv90xEAToXIU3qnyW0S4
i2zQOC00CWAal4M/TiNkDp+8Q11VMymzQzkyHa58ST0oaLBT2Ver86GOLpsfqR0t
E3eJMfU/idN8MzOP2VyeSAhb4JHSVkb9i1uypOeNMxPPNi5tmiIwnJ7bODD9m7gC
0tquA6oLfi2t5V+Pd2fzXHRaqXAS1GC7/N6ZvGFcrsRKkCH1DEjRnaumel6HxG/8
7Bf1A5falYLtmvnxpM32tOFjRJQ9xRx1YMVHrEdsO5AQf0uhGpfXeOCBL5JbDVaN
gNZPk4z1abZ3bVNZX7kaXJ8xTZEvfYJ/BsfSXxMm6WqXH7jDuLI6MB2LgAPzSrKo
XOqFbUw5S2h5IEz8JGZymhqfQsrQg2iNEYcnH3PkKCpJSaz4h0ZkDHrLoy+Y+SH9
oe83khCzKZXQ0PmHOqhOYKo63emBqYfTGjdDJ2EtZOMTFt+EMvq9lNWdcBxX0sr1
XJX/o9r9bqrNhtcnZWkd+JB1NyR+/y1cSmhvZcjh8VDwof8eanwoov7uCcbTH8A4
oi35J/8Tg1yW/2v1DiUEeD04HCOGANhBHc2OBSrRuTIod56AD2PWf0zdIg7oyQTt
yoSEnORtmtFiWPMAGWZTaZDQLo1icWzS+jwdxB0DaUnd51a5QsSzNL0q1h0x6+wf
WTfJl1WXwFXvgr735bKXiZw9Pzpp5cNpltHYoW9BjFBwRSmpfUnfMvLh8UH4E6QX
hB3HYYvn5sK0qN1zPTVi6KJbxRGJ+W/8DtDLRWlYR64qz9/LApGI43jpMZEhIBbl
CRJq4w+WkiDbLu76MjyFCKH4jBAvgkTcgKBOcgRLvEoRR5GqXZfgWsFVMoEaV15s
kHS2DaXVo5rThl6ZNZCKnQe/627mrBcnlnvlvMSY5CR9vAchvsCNsAeiJMvXBW8O
Xjx+wNSGjo0EWVNsi/ovGoYpozOPYn60Cly3G2FkK3IGPFk9SI/N0xjCRr1vreGB
Qn59GYFPRQF4i0sGDfBVfe0HEPfxtxIc2PvspGLVeL/gkEgvLb8S9d/W5cdSRQ7X
Cw35jI5vrLIxKKR01LzbdmCBZfhoe+9+Zb4zCOpFjkuae/3j/sd6/saweV1Qzee5
VPRMIvrZjshI3b93/+5g+1pWMMh2Xmly7sWhLjx2dj7pAMHNR2tYyUpthg4EoVsD
tHVHk/IRWQSrYYYrVP+xMruL/1CwULsw0KpykyuOSRbSo5wrGQ7im5yj1nAK81pz
xCQASlp3dxQCQC0H9qajqsr1NdZksTPMWcTKRp1xGIBNB8jWVE8WnKgd0gIdQ4M2
/PoYCwmzlhBSksFKgQCnCSVkOOrqj9uGX5osr3QZitDmD7vddCefqz19OsA1yNES
XcIm+Q9rLvgm0yMAxeFt34GSGKHxJSZB1okCQxE4yeDsvo0o98XyddiBBO4Srx/D
H8KxkGi3X+s/jXj8hnU/YzC8TRqSoqtiljuoWxGwMuyyJBX4J9liyROMvplGCAJ5
OMkQGpfsyVmBqTi0bDioQ1hOSlAHl6f7VRIU6jFG05PtDRO9kM0Yprkik7n16iGZ
rZEHzcUMkU6JLd9YlQffsojyWLLDrGyd0DG3MidxdyEmx2k7OgglKXKyUSzflQ62
6oN5v/WxJQVnNQOhcLKhhYbse3Kdn6tT+bSFuFryUuc/4oTCSKbGDCqFZQP3+duh
PRO9h9dn0sRHPPbxzoY0GM6hNCeLaWEIzTci0xGeEHJvRpiZaTj0HuvwJ/IhualQ
tVQvLz3Kd887V+F7xdoNG5EsrclnLQFEiN6KL0IjncLADXFbdR86c7JzpK6fKutB
dYFV63+iy3lcN11wpvgdXzDCSbocw2dSErgE2MzfB+S3+gh5i0vavcfof96bh9E6
gQhmxpLZmn2wMxCYRcVWG6D3lENXnryRPSXkm8AmDjnwHQ1M7uIwV69ZrebP0evt
UepKQjPqXGe2KndzcmUSNJKgNBrx6OXoOoIf6VwvVJV0Vu9xQj0oifDgb/tkFDS9
i5iutMTM5UaUihRtc2AcIY9vH0myoSbHp2UnCJ/lOH9C1hJw9NX89No1xrVEXguu
7UH6QeptUGhyt/gnnUptKth0FbeDMMbQ7+1YHHLq+sT+AOOOUVX0jfEbrbvmLqnE
t6D/qJ5VfIXSrcB/v4bc8y0DL4qIIQmddHVgiV9CW+gPfG2IiaDDMY9PgTXJ/w0t
7Hy8qa/Ej7CtnWfJQk8Mt/3JTa/Rw+PWg9pGyvTEXrIU5ZaB4fgIABlwcBnMBwNf
A93U20TcNYvpmEQhWW/IMveZRACkcVpdluxmwF/h5cI7kZXSmUL/G+JT/h3a8Ijt
/SHHmSCUzzj8us9BibbxpxU3XpHn+clpXnm5gp7Co7AXkyjjqOm1IM16mVUKMENZ
UqNRNgoekC0sB6sdhBmf3eJVGbFBN6y3gzBeREAYSvyztbQCCg1V5Th/6zoZ3wfr
bZIORQZ8Hq+HaAddDJ61C+nthG8GZ9CFZXDz55OfoUTArnQNtbOpDHiHanEGALkS
fvBL02DfOKpDQc9O1qs71daq/a0N+ya71j20ycfVTp2VoXWJcPWKQbDLieqgxLaT
lTWEqw72lbkVWc/3JRqMAM7+lJXeb++z8jLbRAsSPwDBhWTcaKRHbaTRncyGCRWW
Q7n1hTlqqUw4faSqQi79B7YcsdJWLHW3K6hK2B61cikzlvC9qc+R2F+GqAwlnB2d
g9Q9N0OclTpFZ2XxACq7FEk9JpOO0AA9P7xgEnednmAW1ApFaUbJHMuBoKZEJ9G8
qV+VGLFlokp8A0lq7iZrijWE7RFka06Jp6mWwXn/32PMkEfUWBVfBoK1t9CiK+wx
XhY8WUBGlj3zOpPok/uYTrtxpB6SeKllZEA3tbhiJsCft/8OhBcjpHsRsDg0yTF9
AvPnVAQi/5DmQxZv5dEHNkQy36ERJGvIUF0xj76vUo3n2d38FpY6/+1z5bHvTGE1
1Sgod5rsUfnSCkWrzFs4hi+BjDat9lMaCKmeC1VQlODlYr/3hcT8lTxgmmxU+rWx
jOkRTAJOUD/vKbrsIpVxiNzvlWra4jYZjWTZz96snV2soxAcYkcGkDA+HqVpHeDf
FZ8xfIl23WT/xvPfuscRkO1QhhiiM4XkHeROsnBbhrPgqzAkgWTAd4f6r7+7eGNs
HkyazhZyUl3Y150wHviDcHgrjwIy9S++HpoNrNppqnDpi/fTgC/U8xgmKL/w8NFy
KVilzSmpDmwzUpphfI6sKerWs3BGJTapSfxJRVe5M+zmPgkFw/SEqT6DTdT+y2+F
GqoMXoQRzPAo8tzY/gmdWNviV9j8krwm/oGUltLLdEi2A6TTQHqKZrPjY5A38bDd
qO/QbyPWLG2FVlwzA7IZBuLE3kvqgLJ/046axBQ+nYEnSEycYU/WEIyxaXfHpt1K
9Yx2F4/fWYmCIdBp8RiB++9Go9Rgk5QHDAO4fdLAUL69s2DnL+hkLMu/UTdcE4sD
LC0XvUIsFOIZ5buV7+2l7LplH660VgZQ2JLiwpKHP0B29PG1sOfTEF6SK6xHC9A6
2UE4HABdVHpt97ztWMURKvnvH/3q5qMBz5xOytyRFViOISTsMm1I7zdWHN1aACAX
FVtxj1OD3PZ34fGw4HQktUfwIrNRgQAWqYUFF5jTrTsvOrgUjbWz578TXq2+pVzs
Tw4zxo4jjpO+RFN2QhTcgdJkfXi1vkdstw3zOkTUpmzhJKxU/y7rFzCrEEkNkWlG
uqoHWfDldEF90wvzjdHmy0LYBNGDPCcq4gVQv1RC6Q6m5YNgI8knOpnlNmHM+XaH
LTvTomYxZsoETTVzXWzUYxfyIl3PRzHbioeEuLr2/sCbOCbC1Xvxxx+KayTiwwMr
rRr1LCNYIiZMNiIpNRKfPadzCzETr8SsuEawWhG0YMx4qxEc39dyPW5TwSaTmqwr
KQuGHnQbFNW142yX+xukDIEQz2IYATWmbRJ5WYf1Wzc8lwK8vbHWl5KXmRbeXXz8
X9wTohipQ/B3i6NmH6Aa1i2K+jrbu9zWL95+1Yd4dDsATeLqf0c1A8XpTSzR92TO
u/OqhTYnfpTkfa5DrgUAIqrdsZaIWNoFsPpr9AfzdnxfSKe0weXHNGq4UTIU45M8
ewEvtpFUplMYwugkI2lZSOmla2RgAx7F+hKEvrk171Ni49cCVii+ZeYYJQU+DRhH
eNKmGlpKPZ4evC4OmgHTKwCUbfPNkyIr0fLZjaUHIqC28CgCrgeb61lCU3EBJ67s
iHxqClmiinHNHV2a49yDFPZ0/fvP/K9bthpvMgiTZPfxLyRkaWsxQb7MiSfVOo4w
lxqJ8IOfBZj3WiB/Y2Mcfaa4r1BPP0EWg3hQQYtjazR2YBd02i3o45ireb38+kdO
HKT2UJN4v/sVpWeISYfTYl02hYK+E1nFj5YtdCjluKSOiMIo39ATY4mKD2+aqykL
8kuOwUfzXbWAFj3ffYgd8/yneZ2UtC2H8GX6Otq8SHMHkHosoyrrIjsdM9Dys0gD
wb4uZtRhiRVbE8RfbmSpUQGz8WCCW870XeS6x5e34PiGKknifkM6OSUePnGXNePR
TrEOmCwb8MUMOsfPDMQ66Te9D7rtkYzAiYQTtwgNG1RwKMBxLfcw/UG64hK/y58l
Waf8q/SKaY6GyV26URMIBABZjnaZd2TdVRVWthRDobNOH3h3ZTgLpaJfFsUSXNQR
ycUSxQw5INQWjk0dYHWs/Fg5UERvfRqIUgvuBFQ/rozkGpF38j4m1XqwwAyqd1A/
GlIktbmpREbeMrTb3uFUzCkl7rdrOVcXHlmunQZhzJdpC0B/ct4IxU6Yo2yEvk70
Jf9CX9c6KBZWTKX9mlA0rtAb8iVxhxyx9ccP0RB3U3X5d/kV1i01AP/jRylmG/UL
Pl5/qe1dRcjceRkugW17tm3eOgu7ywePWPfdK72KiXMZIxcQ3R5Cr4OtAB1a7T0B
cXGv3flKZgBBHcKYwKc9gMEhNCByzJQMAa0z67UGtMsCvevmhkEpSqhmxhEp686D
+P1N4H4Po7Jr/czRO5B0luTioQitT+xf3t8Z2nqXhJ2qRzq9DKF5P4ADdyEeMgsC
yxlMndba6yOOYnlnJ/sBTjQkAOvmaC1fv0uVRxdZKiL20OPlPs6iUDvA8rOyJbZH
3HOynYOacmtz19B+L3AnYiKwgVVVRMSNJksfntzPNc/qLGqPpj+LveSKq9rDatSa
k96IC05SVfRKYhtLKtoYBOSu4M3POr6s9jtWBTGTMMe5k9gLpNxPO9SCc8X2+l9l
ekAbiF/Pl0KwvOo5dLt2g00/6MtMVaDmBR+qYiTxiZj4ob1QJZXVwMn6zx6kXhv0
f4h9boHcNi4iEGFoYzaJ6DkrNQZTwAuW4ulRhNOUlg2hWs7gJzgQE1lVUj7I7rS9
IELULUOHSTJh7tdgt4fAtvHn6pFMe0+y189a6aiwvqXJ1BEfvdC3H6tW78NhUFbG
MxcOhGMK7B8enyubFKSUorEtdcXU53RV+UWDNxACovyVQtPxQNzQTNWajXdC1HRy
FkWDhWorNHWGHvUlMGbls4QI5yWtnTpyWjZuBnsfQ6qcjSLgIFtvvwPSmfybFQZE
MK+WE8p8EtB96Q1LxNCJZgM6pzL+WQhlnO1Ht3rhruyCb0c1Bo/L+vJPQgCcBeMz
FO12bmYFRBpFJG/Jgc6VJioUhyKLfXOj93sUHbH38AtFAPSFDNB1mqxc13TrOCTk
OY4/itk/BSNvPpLERhnOagJb9qREln6alf/0wPbM+HE1c72otSvsLJ0F74MAbs3h
E9yth275WLmJpi8+XofhDMWM/ktRooXVXmGxRYVQP99cY24Iefh8osON6rnNUi6n
c/UHnEekq8yKY0Chzgbxuf6ONRvDy2JakKPGyuxQpQSlYS7txS3TDaozt7Cboh3q
tvxxbVxvYJkiotR5cpRVrBXBz9FVmoJe8PBiGWz1OWPvMMMC2qv7T2Y1RUdX7VwF
RUX+qkpAmTtKP2js3Y0tYEe9QkyvHEvteV5guaqdvO07D2hO1+rYoLCKjI4oWuTO
E1A+Qb6R3pyc6sgz2j8FD4l2tP7DjRBvuLlHY24qvoPh8iOBHYN8FweoYKUb0fMb
6YBioH6iQ5SSte/fNBkxbnoClJ13jKkmbOmbYTBHHcZ2xTjMaXi6ze0sY9HVBC8j
e4cjbRfVFcYhmsUsu6k5NcPinaWUzqUs8jowXE8otggQTWcEv4LoUGQXZJlALZJu
Q5y1xQrlf5ijh2kH82nKzeW8XIIxztjZy61xLdbtb/a52KtwHQm7zQUtcg2mFWPh
XkQvjYVyaiEt7mVpBUaYh8DqRhmWIBgYZ3Mb9OpIMyQ+WTPTs1txm3cBWZz8aple
x7XkdAEh3uyW7saT83mhu0aFYLEyDXsT48oAY1uHpTfzRW8c+7bqNFID8uGneTRt
nRGtufv9I2nVgQw20+GiYG3c5MW5DAfLv0OLTVmx+T/HfxvOdaW2lbtajHHBRZdV
gx7rPXsczmfzjTv/Tl1uNEvUrDs+6xmSe2Q3jJ6u82ilw4n9nq9kccJpBD/navIb
RDZiXiq2oCZO+m+0KQPD+cLuver/nsGrG4GlhbqRJsyFdliSsAlb+eZ8WN7XxvTC
5g3x++VMX3QEDkh36hentOF04uOLs4ebxS+mL01O44JMBuSmSE5/c2WCkVZMIpkZ
MBP/0WOws9VsjnZ3aefDQVe8i8Pa25H2akwh9NpXEfAo2lR7owiXaAlPs3OyU8P4
0dk1+hJuQ18CS7Ftx434EWfNVVx7SxZ7zFsx8w5wwJCwcIIrPSV4hOkIw+uGYivy
1X8yeFFd+bZlsMBOoUlUNJ/lmhPDuDtBvKGYYVSSZCz1lP2jH1+nk22A8WX2Zuuu
C++T65DDZUp/3iWOr1E2pZ3j76oPCYVw4ZGVoVgHFcHhn+KUoL4L4lcedTNbrt9W
XCzHdzCl5lo6+Vp5w5/SSlyyuxdb5LGdWXNqy0Y+ftmlsEVHEW47wlzq/UvnoKxd
m+Zta3Ut3FVfRmxyq7jZ3AYJE22/2zWssEbBLrKaNDJOq9N2u221GZ2LKpaHg0YZ
5lQqFC+WkQ7rcDQIFmpohGVfoQDeKW1MfvlfE7qyQCgTXDFnXn0Y0pJ6HYvUMThf
kWY541ba9z1vwV2ZEzh+2oHgNpA+6ttcejW8fgt0LQsZntF6Ha71DGh2X7ddqKY4
w0U9SfeDIYZYdvFcfa9/GbGMJmbITiKtH08WUWYp5elieev0k2c1V8xEy3J6wQaB
EUpacZ6VDgDi+K3db6t9Zlx71cxLF9xMPLa7QWTx6mj1Stf/8ED2ajsu00Ds2ayD
0Y0859qiGOD/pJ84GLPkIEYDYNQBVCMR2jZty8i71GEkfRPm/rje3qH6OROzFCkK
4cYPYRNVHAI1a6hV14fhMpO8kk9GGCkcCtZGSKxxRbQrMNp2cLA4RLvamDjiYrYg
OXJNWeTw5G8DKvVw9wWxbg4HB1+KazZRMfJLlc84vMLTVjepheXXqNfKNgLEXaIs
otS2J6/OoNJTd/ue82UIyuaMGM5A3TLCkxOFd9WKM5uu0jFQDGmMrCvkPi0ib5kM
hVcU1HxwU5AGNTLFkm31rXradDNrXeCaRM8wfJE1vgEWUrNhIEW6Ybk4vPxhoVGM
EwT6XkXZgs1nVl+ZMh5h9+59fa+K+0VbASgDyYCF/LbMQKksQB9wHuwaylJl8HNM
rQogV3aB9x+HVycF1G1/+LuQzknOlE+1r3UXWkcIldb0Y7fXz42bEjw8uRpaAOEZ
difTc2miOaaR2XYvdQ46P77bzxSjhMPn1jQ3DNslDzG+peGyWO/lgRUEvu5HjKKm
QQj3lixHAfoYN7r3iR7iwLbfkWl+hjCsQTV91TAplxWzlpei8EmhwX4MBosRJcFW
kLL16KIVK7q1bBZ6nAwZWFBgJ4MTK4annWo7guTVXjO3knibfqMv+rdBAzy8SGKu
BB3M1E8lczLnJRS04rwzwxsLzA2xRHNbLfE2MNOIFrX1U854ZzJTi/k3mgI/08ro
Lhs98tpdDf81nAcgRAOzLLhPSNJWoYh+nb3JjhVNxw1Lf8noNazV3iHuD11kkWET
uIFB0i4NqHHOw6W+gVzyQyg8EPLeSI2B3xB2IpnXyvnB9TLPsCdYtgL4VIKba8Ye
GChynaOhFoCF97z1hOkI9KiGwt3DCubbz6xcxInonP4Y6/FqursrYJM4XcIpxXOA
KWXX72gJ2Z4Uol03jXAggT0VR3CUbQX3J0NzkJoFqrJQgehQrU8YCDJ/ZG5Mkki0
LOZmp3aal8BEM2+OD9NUmIB1JBX0E0qgCkQmZ8rp890XeJivBRzWvasGdDwRF0p3
oQQcR5x51tr8lkqhOn9gprm/qbcy4YT7f26tbHvgH3R8d7z9YGpzedATfCwPZ7/Z
vjiPshUdfmj46CSo0zFtAcIKkH/IYH3DpYEKDb93sl4nblCWp0gZB3RM2w47JD27
aCUXoXYKWBJGA+ljRYRdiCRC2+6a2n4cPJ0FVqC0b7kYw8whGh+jyHpnPJRk3D6K
CL1YuhSBUdptmsRGXaZpszGTnoayzT9wL2PsqNsSPWZCF5a0mxMy2y0Sf7ZpkK3z
iLe/7wu5VoFzqJyAWomdn2WJ/hH1ByxW2pirVGF2WqeIsW/5T+odguVyvSUL8cBw
QLvW1Og6AqaB/RYcbEhVlqxddj+0wW965KgWuL4QRSrzWpMthxTXohg0mr8qKhaO
B6AKVAsaW48EsMonDDRkgZ1lOg92gU3pY/YfM8eTU8uJpVgbneVhpBHMiQWXw4O8
B732+YSwjiDJBaIYNeATfOrCFuXAo671Pxp1DjAkWoysiabwj0JyM38NFaB2PLcC
t+HfRbMc3EhdMXUsOIlq/jTkJGKEwh/Oy2RTsuip6R0Krd9d+5+77q/a3c5RJJIz
+gD0GqonzNvyiWkuz2wBW539PHQRayczXHquChg5qI9hqVQnZDbDBkaVmFnAKg+g
XoV4blAyGo5GEoprqFloyNNqtV+YfoTs/7cUCyDX0AkEACXTojE2QLnlf9Qu5EwA
Do31eXxxdeiKGDXmltfVA1IhWVFuESSJ6qkoz5pm51MJMK65haoD+lEsAv8MjBW3
ZHE2STf3JsiMOD0Aj8AlbWa7hvXAG/tbHqZWkMYUtV+zavV1TJJ+0CVH1xl39iDo
UGgnNBYBthdEAvhrdBe+qnnuiGw6cbJkJBrjuGLz2NpppXVroPeM5xXhtzGKi+T+
vCsoraStG0qUYrOrCWwQYXeKf6IwpkaGWsS2D7vMYuXARH1c8RpAqN2L9B5K1f6h
gVjl+bOyji5u3FIPhjOCBVrgdgcKgW+ScnhbfwBIOzZ5UEk/Lh7XLcFRXEqllfrH
ZvFSsd4FPt1fh5L3kno6Jvm44sMl6S7GxrHa5AGa4GbstEdELU/P9RjuhSihSYGN
SCSkKwbKO5lpXEN1HmG2ejEAEplXS0uKDu2QNti6FbEA7naQDBBxYNzX9qsUIUt6
KjroAVPu7m7pEe6pW0ETNvYidyLsLX9PJd9wQxCzSUm+Qahp+aLzo+2B5qOSY0PI
4Zuu5m45Yi8ADRjWqJvqJy9U4yV96fiM2lqJyD3Pr0HwHDEk1Y6HlD44OFUgRSIy
y3zAkraOFHxH5PVQ7950FVTn2mbvW5Y384bB+oS/bdBisz/VeLhUJhzbbeFU45JM
J+mLpUEoWz33GRSiLOGtIO8vAI0X6PBARB5FM8CzRK2b1/LOsuBrSzzJ/BCVbQ6W
JHLhmy2a+oKAo/IWRcyKZScnDub1c6eVN4xuLHAdkLXbZ55x3fdQtyPy8sDOK7Gx
ME0RlF5ZBt1rlu9k84Ow7fz6niT4OUhhFsxZgaZPucK/Lzye1MSzoBDc7aDb3HUJ
PZKRaKqMoBXQmlYAY0XGJ/TGSlOSgfM3JMFiV6Y2DGFROqz3CbSiEebdVIPNdAEk
V9EeQv0mc1NeivcPLcvibFPrZB1Mq5TaXnS5R/I5BziKsWvDTQO3bPEl/axYB+cb
8er3uuh+56dNVGd+rSNQNR4n9EUzszwEiHm15EgfM736RqYuQAlXsk1qo2fOmQtu
dYiD22Szimm5KY5GXNv4YVSeaV1jwtojf/5S2E4zWJDIXNYMbHKBEZd+KTt4RGCr
gZVQ57y95Zn0KuzYhDRddDXU/v5Gbvz/CpV8BEy8l+JuRbFe9WWhbnfLBynTXqoE
M/zM37CX7s07aqVf6NFfq5FjyKqmDVMO4Jvx64lFc75eYoQMD+Akul7TUXCQh0Ls
803IpVbNcipHZetU47B88+36Qxvyh4AklbjP9RaDSNOhZysgtmc8iPJagPJJ1xvC
k7c+xIk5MvZ3lGPJPDdUyTnexmyL71JQDH9lv0qBKuz5LIMm3Bkl4alrAoL8clbP
Q/PqyAAPISLhQt7evXiI03UdTjMIxiuRnfryMkRm8+42gztxtnX5AnPUYCAKFQiM
k15VQZIwUqgpeHVXSqkNxI2HC6rx3bOKJYwvSg7Ox6TN5DeiBtcaYj39CumyTt1U
2bo0QlXzs7E21NGAc3wu31dT7eGwapQseBTamQjFO8yxGxiGBZfGAwxlJvszipIV
Av6+3+zHMbBF1R/E5a2IZmvB5ytKp2c2nNf7XUvbUM1Omp2Phdf6FirQt0N5jiOQ
dRkM3HI5lFsTNeW2aPvwnFSj6/cIkn5trRe0/9D8Rsug/OYVOd26d+H9OaS+EaTU
4p7Fwug6UHDn5IspZ31VnoxeYbHjXH16t5ghpVVNLIQzmhLqInXYNCJFasZgnnqm
di4b1yWLLR5um1PKmYB6iN+76vRB90jIJiHAIOWDRpBBAE6bwjVpr4bfEx1m1KHP
7txCHxUzJvbJ3EJ11oSQNJAieE5z5e/BeZYd62sw9cBbn2uTxoDjDwu99NNnOXB4
K3dX0v/J8Hk9AtnWAZxQcBgYma+uGCX7SB/HXLerNi7m0U1eqVXWJ3g5Kxk3BIvm
ZoCTBLeQr/aM5DT6hPkSxs9HUp6RITy1CYSu/imsQixy4aQwsPi9Kr8tGoLR/ruU
2iM10WQwi9QLaLb600BI0tyomMrACMOBe++EMUC10fsWOD8cQ4IDK0+v2UMZ9OaM
d2wF28vqMKZ4AruQs+pbva8LyoVIRJoCvezrp7Cr0PsI3Dn0TKUyDvNPwh9/2fdx
8OCWVV/fpgCoNxI5OktJd+Y51DyxW435TnMNhx6Q5C+tBSmIEMxQcsJo3Yloqmh5
WrZEAeei4JdVjMw59dpZcP30lW94+Mm/uBs+PlOzthGmXR9d9GAZGyT3MuIPNrzo
ZNtnjdGDdDU8m85Z2qM0Gg5LVkPd5qtk5w1BzuERYD/qeog7IrPOuFZRy/gl2lhe
qW3tLdQuDXm1q/uuE9RvXOmn30iz2D8cc0mRkpC3IoCis/kRkk1y/4IF9d+g9lAV
iteZAJQ+ECUwtwRzNTKxYaBZhdQuq4euo5Es3mNNqCNbgmWeOXlTaIPrTmxU4DJz
rprH9h2P9Pu02pZLP3ySgBqLTSdpSL4iDGxT6FKI81g2dpBGyUhexEkMylAwDNX/
6sOeQo0cPjWgIZsj1dkz+xq42439vgA8OHya2LHDgE1r8GqYvappDxEUC5NhGD5C
lXWww0N9vJz0PBJqQ0H2bZK87rukr+eoV1XJis1xf530Y6tnl8CaZTwTG6JJQk9h
S1B12YfOwGS5xo7PSAECBQGHlyI6MOzaICPx0P+1WgrhNVtmwNjhOsByeE0rScfP
oYKzroun8wa1Wz8BFQyvRHnMGEpfderPchXnXwjOjTBMpKMCGMgvLvLRqE1z/5Kn
n2+TvzcM9F29H/9JiAqDjvOd0bJRW6pIRpCS+GsBH1DmWwggycgmL7FLNiK6Z81n
08iE6Rig7ov0F7kGfHtjUEeQTB9vOrtjbYsbmBuWsPpsaxhVbmyrqIbJYJaDDuRW
F8+Iak3dLW/xiGOPR1+nhmyFCEEThWkgMOHn3u0zJNh1lxzKXZnezdTBvfgJfkly
Q38XfnUu+GP6Cwytl1SumsmkQp3qVSiIsNOu1CXhMctPbE46H/ue+VilrqPhsVW4
BGSHgB9yftcjM2V4DhXvw5m7Eh8cJM3CqR3AHskRJZ1bfj2dwDwB18zCgZsF2SW+
Lmq/8M78BorYkvXPjJvP3ETp5SKRYZBos209oZqQGFBM1dgCXplGTP4IX3tj+sY+
WTXrH8W0LD6RoCAjPYaKzxJ+ewokXfd8A1bzVbWp1McOIpsOUZBNivaCQCBKvtHw
tMaHpBf7mV6znbfgDz5hemwh2XFFr7ah2gDpXUv3V6LotfIvERVz0Fg4cgSQYOIw
djhJduGZFz8hVd9lDxExoaHR/11Q07AJhyzX8zXP8qn8hV94nN6ZtlyYIapaxF3J
24jQaz1pZv53dST/a4Icclh6ShpG+Ai6nw2TbbIXb7hBSYaWItKeJbfXJfCmfwGC
7MM1UlovyR+3K8W7oRzmqTUaMtdKfWlmPZiH5/553cMeDahF4MJpgB7IpIifq7JZ
37VQZi5bDS/Q4fLzVVezgHmcaVv5fzJQ1hiqkr/n1dTkcCNEhnybphFDTAnZkPLH
0E7rt+XHXwLlVcKKU2wTMOIiSxJRyDeHHKb15QgRpn6rj1IlDLgaS+iskEFqIUwR
qjqpOGOi6ugop4Y1JJx9n1HNZbjob0iaKww3Vq3RtzCNKjAcc0aIGFG0zKg0SHHI
g2geLwqpIGrfXR4GAgEeSNPGmdClvJZ0wRbqzjmYtyb8haww1nZrZC6JEwdavhGS
MceM3HPKMkLmfqDyH1S11DAuI3IEnX+6InqEr5C+fptcVCLdn3dD7SI21KN3rW+a
zE3iG3F/heMoC1HuWBAfi2R8kgckyifvm0lz9wlMihbrMTm0RhtRtoVIy7k4blxP
4Z6YWRunDOYWpE9eenDG7Lxhay/WFcZpL0XxVPXBeT6PF0wQFqkAOztjL54Fx++q
Rs84bpYbwTND1gCVwzhVUZb3tpGib+kHY6ju/Ygh8seEXOOd7FA8KD8fqKylOnU4
JbqGJ16Bug946en59tqVBy791m6IVENkTYN121vDNb1J20k50u8PvxUgu4zxzgNb
w5++9fQz+vTE0/J5JGvtexOiRA9Z+UmRUiBPV3kfFI0xCVvr7K7MusuH3PPZbNd6
DygNZwzGGr8O9W+Uvqe+R2YRRBhR+RPtzonwl6goBX926Ia7+26rW9nXv9dymlk4
/dKBQRnxPqwLxel/5JqYWy5r62DPjIZeibloNKUSn+sx7v8oHEdTuYEuvdNUMUgV
DjgP+LetoMJb42/Ckf5YpkE+uTL77cukGk/uTdBQxLZoW0JHnQ7+0kILiFrLDWrk
Vf4tDaMgVP2TEfMEex3pbvhEfosHiVMQyU+ABxyt5QXfjcDXtmVOF/cnhetVoqNf
Yow+VbuWVpmy6fjEqC5vh7a860Ez9JxdgiY4jWVbib/3aJtdXV5xRLMDLNJkDEFf
/hyc8DFKYW5IsYe1wzLAbFmHPEtUe/pEhmhrdNoSCDt3LFGFIYCNDLsR9zGIDppt
seIABbtBW2WnJCPjQHRRyAn6/kA6IQPquQ4FZ+M5yyA7Q4MEV6nC0GpdeGgbEWPo
+sBpJ+Ai40WbSB+Po/WntXlIgLf/kq05+ir2rhrQCQvHIVEuMRmj43p0g4da6m0O
z8R4l2VHiTUJUzoKI+a0L1/ZjX53tTGpIxLr9vVIJKi9RXViLe6FHdsBPD4bNIts
geT+goSBASuwy7lDuyuQQ/rIBKNXXhHSvRLFI7BLzHMT1Mi4eTXfE5wih3xR07GS
061ZM1dB0jUkcuGfR9Fgp0IP/VevBdBgxlMuM29dthpZN2jwcWcbjFueYkLlHgXG
le7eFTaQwJEOTtFqQAClaxgLSMag59ljw8xgUKEkFwBwAnNlPEIIfbWxLE7+haRb
jvu1fFNtTaF3x8t5Zlh4LQoAxWU73NVBi3VtKU5kB8XtbcwzKsJoeXD98d8846Sp
Gj27ARqa/PPZkMaZmLhSgxZrb4qnDesVwGgpPOsEjs8nsLhE9eS1nSDnp/nOBlq8
b+mAYm+47AILtXgzNBdLyJUHlgkhnsRxvcsWTcuX8SxfUS5dR1ncR9Lb1EiL+sH2
7K+/OMn2rOEbFxGpeO2eVpAfvyLioOCZguBPr4PxBPlRFDts2g07rjGmS5ef2Bhi
baAwxak5SS713V4xp6HXkRSwP5ASRkjmPEgmpHcgaREG6NJPdOmqq7Ma42AdCng/
dniHb1OXof3GaPv0uun4vrJAoBVaKcg6I5T8qf5MIIB6CV6jRQNrlXb2N3/c8Cl8
lzNRR1UrqtPdtPETIRLjjEUZwEZLB6+6SBWtS2TLf1dRW+eSSpBsbgVht1Pi90XG
dzRTkyOllX2VKuaa72NUkIOSPOq1CMSqaJwUYR5kRts3Pt0mH9ZemuEyXFY4IABO
KvXhAOVxwBdAPocmJlXvnmOq0qqIUihSULu040bITe7TBpPst86sKOlsNhPXJARz
bfoFobh+ew+9YdGXU59gJkB1NYVzEChkgHSqQtkH75XDilzSWi+19uOnJUAMGHKn
nVvQx9UCUYTAvIuc/DurfWNodwbC2hPxmHRdU2IxSnw9jxA1cWSAAXhFRcGz+23z
2ExqyaHIJieR4hbm4NY6DEoX8MJePhJX9jLHN0H0OZIRCvzts84dVpvgIF0iAZiC
8dXQCpPUpGd0srCCTlY1mSANL4MNTI+qqdWMN4qtisiLEW365KfxG+Al0WmYh4lu
aIi0ysGPrdiriW0viBu0P4gNt3Bc6HqY8wX+EKJZj7Il3ooMwWamzx4NSu8fxLCg
Y+smkgIPVKEiYNXIzk99qAnAG3AIEiyMvC+/GJb4SXw6FKxeNCz6kTKc8/6yH0dP
CxsuXGC/CDrF0c3H93Pt42rXiJhhX/jA6ZD6RpCfgTJuEGl5Q5dI0TeseOumV6Wp
Ju8+bm5eKBL+F8620cBUmAPufwlZAaqzvRhjGPTy6wprtP9ZEF9cwGv46/tHvB8U
ASzFWD0TYBuW2/UVfPHF9cqeQEuo1uiww7K8t9diy4guP2+wkrn9C4ylvMPKo/ok
3tUD7z71cmlF0P3lRjU00JPZ3U3gS1wck/lMPl5LQupo2oaLUc72jnDFsfKN2rsr
z3tV68+x5t4PqnQvdpp5tkNavbo3IK6qDrJabLKR9arEI8EENmYrn+4450C/Uy0e
Js+n//9oQv08hXl47Z4lCdA8R7TxXJnjYP3j9YUw4XNUfySgQJUrb7j8PWwBCp6L
qt2zl9HgvryTGWkxVHxD8RmqfDD4eUapJiEfdKKwPm2TIyrhX7v4UMtdPIcvlu+f
j55kKokypEnSP44arj8zRJArmEe4+x7oDflJI3j3hbxK9LgtnwiEDPXulpehAwso
ELnrT7NJVBOYOeoXuKKt1OBt7ywdVOyQ8nrPzmMoviXvjbp6h99zLbd+9YC+aC7P
7be67a7oCmHRqFwpV829UZ8jECVUFyWRD9GckU3UxT+qPhBMgWbGlV2shL6dbwkQ
8niQUw6OGaz8Un1Fdjs85PXVe63xCR9u4q+tvMOuFU6CBFaZfdpAPxEeLx2kA7CP
0bU0Y6xWkFQFciAypqQznoNsGBgVVhf/l2k1zJWVvJp7dRtI8fVOb3qCP+mNLEgi
hrpqSEuh3NuSRyQ5nL4d901bHjkCmrQuoM49KwQ7tNFWRVZYoQSaN4YjjeKaCLiS
tr3vH9jJ39Ovvc+mZvZsYDV/NWuFR2xbXFVmMClimUqAj6HFjs2bgHjA9nqb67iu
Bu3S+15hblZoTZwVlpk8+DL8yrSNJGwp7BD0e33A/0khLaiB56JDSqJ3OOI9QyQ8
KpdpofaRkWM3vH0eCdgvB3OEx3Hl6NupiUePViZjqVHbXm4jPSpbDz3F1/ygxwd3
Amd67R0Vb9HOwXWwmu6YbrZLrRhnvbHGKdMoCPCz0e7qGK1Iii88MzgLFvDqQWmz
pHiziE8n8dgrkn9qENCqZbbn65sZ3ZA0GfoQO2vNhbTWwG8RoG4bzXZwN0MFcBn9
ICfNAafJM275oWzoDVfVLQ1YEeL4005UlnkTSFbpoN9zzTJNH6xW8nN8rAY+eFc0
5ClFlCSIsy/r4uQ3dhRGmW+txqn79xWUPqydsoKfIdZrT5ajuUOscHuhnXJG1xBv
I2sSvpi8u23mFrhpva9AdQl2QOYqNE0WcW/nfxo/P/0aAsDNAYPAJ5ZQ3bTZnEB+
esM3zy0k3h6Y/8GWvAajaWGNCR2GqCLEqU2gk7yzg7jYlPfR+d+DQo81GwQ+bogm
VsOfU6jea/WJnwjzLvC/iVy7UXQd1HPnHea/WMgHwY2gloosylDFemIGcvrV98za
yWSuG0qdnsouakcS4v0xjQTBGu0amAOSq8JifpNlfeXBD0EBAYJrK+rayjl46Z+s
dmq/ovjpbmyLErJEu5TQO3X8SBNzOlfQBsaJAT2Fuw5VIOB0iq+80htCqVddpugH
Az6Ko0Tn1x4BgABBWqnnrsbK8JMpwpnos/3gBXkRWWwhN3Ibe8KT37RnM4KYjKPH
mM4URmyTwm7aYwXCmveX3Lmi9fbkv9oblqLSabg6x6z+3IGj0rS5QNANYhpkrqM3
oHuy4cVC3Oqc1EExVx8J+FcO30+HygeoRWhX9c+4IFrjdmUierAxX4yExz7qPN8o
b1S1sbFpvqVIe4xf7J47TqPFTd8dg9ufxdu9+GBLR6ZtD6MdDpMbEOyob92pNTM3
DolNnKW3Uuje+klp5mc+k5DVEwBCqLTcPcp6MSN32toNBF+8FpeI69rB+EjX1W3L
xedHG5Fte0LXYCloRoRHMvVoZcLAgy0GqHy77JRH3koDVzkNt4pqJg9VwHwqAPLk
tD/se8BXoXDcQLPutPAgaUxKMh4ul63HCpYNHAkA+Bmg1pTw8cx629PUL21y82FB
vnXzfcb7pC47A+udFYjdTwjEfrrwfkYg9hRVtvnuCIMEu0sDVhG4M1ZwcxH6H6p9
JUfkTbb2bIzildmxLXD1nsi4fL0Kag8G5ypq4DDEg8fJV9CPhuNFF7GwIp3BAQFV
ymZp785DrFojvCCCCldiVoOcR3H7UIS6KmQ7DhZg8iZF74xkGaieHPLtKjacRrBz
qcpqzY3gbwNCOGTFE7d40DYbpPHfCm18wxzI7s+RggaPcuS9/3SATDQE5uXo2mLG
fTcsQwcdWSzn/RtCOjm6omA1TjeRuUzdgs7WSSyWkM2VSLqFkiu4n5j4ZQjbPONc
IvP3ypHKvni5hX43TfkL554o7AjFnUpSLWR4fx2XUpB5mjgWmaRT2PXl+iYK4u0F
rtAFg5Mzu/rK/qhEoQBWXYMHg7ld90fWFIF9ySBKswZ11Fys8PvW11H+2AKERHyY
T/9EbAxXHZid/rV2GFjM1fL6U0F0j6AAqBn2R2wB9rIyG8tYU4v+rKe3fLE+iBAR
/CQu4z8YgVKitpk47b0DnMOSYLutSeep3tTyi/9MuEFFSl0gFD+QCZN8Jin6k6RX
PLWriErxyb9EhYFgn6nItb+PweA7g2F9FoZ+0g2wk/PhLs+2xuyDMotaWRaITabG
QzVttS+nGkpFlfj3pxz7cq79y34WJagHS18AXbWjDRsLi1KLDG8UH97st+SsOEIn
QkUS7x/S6jtm00Dfpedl7cP5v1uAezfX0GrI+/JTRrlxnkuQRXU0kUk/fuKzq+4E
ECSczu7s/MZN1Dp/eFRjXNnRmql1ghk8FraMhaS2q7G0AlPanYE/KiperWCR5zoW
PiKwwv5/vP0roZRNpsxMgnbcsB0TmBX89M9BiTmgYVA6OIM8u9amN+/7rusnAysu
0zHEa4GqSwg1M7MJLpVxMrv78r8fNWY6gAtmFJw+7g2Xw8Qp1QHLqUDYOkgL7uRn
BGEBXV+HkpuJYxZxDDZYCrYnJhvxXMHuVn/J3nysBDRdX+NZ/+PnE08CpuUFg8zK
Kro3cuJdi4fKdnKlX68pv5nul5cSmP1Uf2hd2J50TacrIHjnYk5XU3/sYK21g0tr
3I9F19GSJG5Mtm1tf6W2TpfMFDy9p92Amk7iWQyOuH3UWzlUsy8dmYFgUfthB7GN
9CURAU6s0Em6tNGag7Zn613J826IXBVt3KqPtPuXmSr7fjAorkOFq0q7bh/hzKUy
h96l6C4FGjOGjcJYcR7T8qzmjoo5dsw4v4GML0zDg1zKFXUI6QIOqROMPTgnZnLh
HwNvZfFp6o+PiEoE7qOciOWD+KObcqYWuGabs4aGg4h9Dp7XPtHgEBmisK/K3KMk
4uN4AyXlbwjfWf3vVKsNbjcMEkBVsz7AQD/3gBTenv7hagIogcLFFIIAXxEtp6B/
fOiDGWJIXchxPjRPw/attq8Zk8XppFgGSNO+E8dD4/X8ERFHLNlBzJZT5l4pXDr0
TtcsJRqyCUL7HXD52RMnE22RouQbQIONscO/Rhzxb/aB0f9piE3Mz5uQHxvXjkM7
3/PbBAW5E2lzupIVxIrmGRW6mVedy2Zw94p/tlFzJTAOioHwN+xpUob+dkZEdikO
2CU5iL+MJ5fIYh+21xyEoa/edFHf8ymseYrLPR2cuGPwWyA7UzwM2LHzN/t50iJx
HSI+S99YISbpZJfISIjNam5qVpx+8iUMshyUfRb0jq/qPPAo/HzJxd5H+qLPWDDO
Q7mnbhUjyX6d8Atp2iqN3YbhSmRUqUlYUjT1IRskqwTpTav8ZaT9LJanwc3MEzUy
5wdVoabL7ouY7SvSBAy5yjeQe7AK0exo6cQVbkJi9zMzySQf+CR3tbIBO5sirAiD
J0Qnf4jalxuPDqtVANOp0fxoxyWlSTJxUrn5NbQ5LkXEEF22plC2e/xR0rpwJgdh
7e+Pt/pWvq3ccq1QrUw0KyAwkrB/+dv/mSPqCgDrWTV/6LmBT/IWZvwJ/KdSkxnL
9nA1GvZdre/nQlZWADNSeY4xN2WXi4nRlSzbt/G4MbdOKUFAWU3KGCM9NpExkYbO
j74Rp+ElAe9X+V8KLQ6Fy9SJzhRHN3b4HFNh9AfsW7u8fymCasmacYEpO0zYLDbn
fYmlhmv8JMidDtULKkpu+9SwT8vgM+h1z35X0b8/oREuF7CKeKlIgpgSnVWK2YVl
9F5AH6YqgZVbRFGgXqm84xd2EF/DZ3ygiB5/VAVYiFudSwn1QyV3WvAiwabyoZEy
kXfSTjR6fZysa8VZqKsYaKGgjVqVldjLNVhqnOf/ORUwKZmULDyk8Giv3334fR4V
89BqAWd7Gcl95E4IWPLMafGMe++2i5CCyXVQXmLsh076hGA0EObkxLhRyCeeucvF
L8Rs6bXcuiHNZxaRnT3l4diS+HLP5bztbxfLSzYBiHbNwj9njQfAiPYq+LwlIAxg
FW+oJVJ4sKFlsp/YyLGZsSvP0nxAb+amNAcAjiFfv103Kr39dFRUSgGCU/e7rV6P
clpFhqfC6Vaqt3qbtm7QqUfPtH16GfpjEJOdxGxs0mJiPrT8l77xHu5kzBgZp1KF
/73K44YewUYKcio7CWheDccZGheeDOWSBOQXW63YGiVSK80wanVJh0FuobaeQQ7F
d7Xqrmv5R013+61do+rN4j0XPRevB70hAnt4q9snp6RO+SWofce2kfItbkWWBKtk
kYvHti4srix00a5oRnKjm6TUcuEzXNFjY0t4x7o1lotQHFLbqVqQQVE4QyFrPTSS
pZDLRTZGdxsx5mmtdoQ/dc9YO8SnYzUOl0rVrhxT2FVfJnCzGDUs8hdn5OVstUXw
3C2Aje90vwfa2VYUzWiBL5gYoVnzER2LfSFaK5kNi0zgyXn0r64oJNOrKGhMtknJ
dhw30XFLvdBzNmYjZ5GtoCPR6n0kOfSZCbEVmKvlDmjmZcAldtzKNm+ZezSA/AgF
CiIlHQ3MixTLnprJjaHK0TZqMEhChLIHwpW6Ii7x3CMbCtA1SpUjTA2HPBCBhFSo
YOYCajb5md89vJlSBFEfMFM8hsp1xgxZJ/LlPUkfFlnR88zdUWgfhsoGXTtC3xkQ
QFUTbv8fljoAsArrcWi8CpBLKvWe9s9+YUPA2RhMKAUI06mnqCl2xwhxXuXVZJks
lSzfu22+kjf4KIQbXMj0YRymcLvZN/1kmNnsWp4bhpQReBBaQtbkYDaAKXHn+WmV
hvfqlQrXGol/45UcBnd97Hpq8ix/iGpWCFK8bGC3nZrr+6AH2D1U2CYn3cHljP9b
4aGu2GingEQoauMASsGpXGv2CqpMq8Dw7rFj1P2359J7iYIkBIIjKMiWxiEcwaQA
mLwoUcLPg+WYDK6SBYBpl32pFGWCFA48w7ysasF47VBCr1lKgkhhQmqyulaWUmCL
/muRoBqOH6psCCvRUmIZvmrTJ7KctIGUX2KJUUpgyaea3OGL/Av5NkrwFExlInO9
NJY/8a156JENKAzC6jRAoi70Fw8byFer104fIR5Kmc2NJT4e3uOwoWyrBaEPI60o
jVj5jw/pUPLSD6kskRcRLUqsgJbC2Q00a2fpttZLoCVaz0mlnbfby9BtKO1B0KfV
oRFhz3Vz3oagByHEUW6DQ1Sc9eynKB25llhN/d0Nd1ymK2L5W3Pe+bD23QtXg4Et
GSakYaoYsxQqrQqSxHoqkg++qIxVjCqTT+ylsGWahQmhwbk28Sub/SAMSaFXrt9t
t/Ei6J9ghGWqLns5xvs1cRNdGFTxydnpSgQG7x6UfU1Kv5yp3a/sF+ewCIyIHigl
Ses7b2NH5Kpjofp2PRFyrgx4USM9R/idecVUa9LY/1mj9ykyXlexSS0fyvHV85cX
u+37b8woj1xM8lXJc8arGqNbU5Pr1CRPEqltveDpXlBqVbv3qUIvSa382sg65Lfo
iyckt9zdMyf0XS2K00Yu2I6S2aLp+TsPKNrilqwy49bpsJPSS0GT2K6HITFEDvJ+
1rEQRuhwpiXSO8YXWjKcIV6HpLblJycH9Hb8o/0F916NEYlhxS5fRNvXWz7VZiGN
rmsymLlXTK9sZTYTS3Pg9oVIbXimRJoqqnn/0AvkIaOwahoOgCdS6rotm7M62f+4
0ltLTF+koa4dMtabw51ZDOHUFNJ0SdwR6MmwzcIeIoUcr8ODdm4fU0QOtwWXF06S
pxbxgfuhThL8diXkWQkBmHpFdTDAS24TWe/zF2jKQPFs8/ZaP/L1fu3dQSCXVaNP
c7S8Yq4788Eem0ZNx6VrjwsHrsMqtl/EaSBAFM48TNZYIH1Ryl4+/2TX7iy8ZjrU
OrtmypYBXtRtKhDkYkiGEm2yLxIZnGVsROiIWg/cJNPmD9x4FHIXvqIl785EzX3B
WrRSxP19PgPheM3C/W0hycWlm9VsyAp5ejLwfzQF8oLRm2x17WESZ+HrM2eb1dIm
gLGHuSWp0Xu8MKdC4BpLFwXDdwnojRys66XuFrjlOwolk/2cNbN6V90fZuE2P1yJ
2qDYkJwmtKqmWiK41cDgzqR2/obBfmDS90JJHAFY0fU17EfthIqvH1z3NeiQDXKz
PhU6Em6TMRDz0QsoKJOT281gfjMAfMSgdLuzu6xzwU9BAbS08RM1NA2H0MEXJ4il
OTFclp5TbQQ63p0jObGa1QtsiAQkRPjq4UT2CbJFjacDq+f8rEdb2wQJZH/ENvUw
Ds09f/IPjO4HJhO+MK+HGkvFE9omTZUcp6irLtC4JOfSoRFuFySYstPSJ64yjkYB
fjgu+7zkk4RS+Sj84D4OS8Fdib4ox2ucLC65Xu7E+tVihGP0SaIlqYRSi8kv2Q83
1prsqaRW380pf4t4vd1aQKFAFjT9SR6NTzx48FXv6BZMNvqJ/p+NEvzCRa4PnAwL
8a/UZoEhNRwRgPJqU9kLS526ck+H/9Ypes7rai1GtBA6TXvvSy11sfaXA0FgZJdE
H4WUXxH6FfmIH8hr5wGGzcor/l1DMRGh6ejzweh1+G02yo0LPfDnDc2o9Eaut65X
+hInVfwpNC+BPQgTSyFGAspG5umX/wAkMRNLeYww/bOv8FR5ISMmbWFYrRrrj41l
jOn/11z609b+7gzL8H57YoFeTabaCPh+dPvoUag6weorPrCeskWqYr4kemb4DGQ4
rcJDFeZrNqOrAMlIzYqN21L6EiTVjxqqXZdzNYZB1vh6Y/YS/aMdSHQt5E/Af3sF
WMoKnFCQkKCzBKnMtJn5aaaXwEHQUTW9RG4N7mDRE6HO3Xz0I9jq/pP+EF4+LSXg
vEuQlmS/YT9pWwRNU57pQWyHkfQIWrsZ5xoLGCPCwnGo44emQc1radM4gjdJ0dfM
CFHNZfS+KC0B+D2o4tSnLRhBXw7KTFBWdCbfF5R+uvS9q9lWaxq3+SM9SczxUz1+
rr8mTI/2+jtc0m3S+BJh45WR+Z00O6iRcNUqEhFkqQgNBALrKBX5cTxKChnQmvZg
To4Dx/30tenGBmQ46I299sx8LAaJXFa1zGkaMYqa5tG0nFbteDeGTnzNTe8WF2kq
EvmipwQQdXyCdtZ2ui4BdtIYR4Y4Ynokatm/2zj2gNBCgYJC+yGjPeCSNlH7fPBh
PPoNGa7vFOAs3FdEaubkg7W5mzzuTkKyyZq65edVjhMAeHRNWibO5eFkkCMJI6vp
bkMT/4jLlJuduVdDtR2gpE5Hv6nf6voXt06RA5uvM0facpRm1AVnDg6RJUkLb6DG
OH/VU33rb5iv0rl/W7kzuE6X3K+2P7LbPVaQTn4kMSx096Ztx964ndlc0Agiji+o
z6sVAivVNxx+TkR7MQ4xgwdsKOlNu2danJFY3CBiTYI54paxve95hpe7hI7G5cYD
SY8be0kfX9e46ersQikoxDYJ2NN1cr/gSC6pLctKcERcyl5IIAeumFuEJDsZajPC
4tyBTT4cQMvsTI9Oqe2uYYndAtYHSASPLlvoqWvGgjT/AsdZU0Iij8ll8iWCZGCv
zSKtI9jnvzszTMZfSHBkHqrAdwWZuXGhaEabZLwvmeeoiNL8MWYYwYj40KIgt3b6
octeRpZdgTMhU7reB/PEqiGUBUGTFfjGI3oUc4NMB7psnO5kqqlySt+Nvqj5beFV
67BTe5vvsf6wxQ5yK716nDu5NPRPR9RJppIir/3iuq/Uuqd4dLQPwxLIZjIEbc1T
w+CzjO2p9uqLcHTvrBaDfnvuj39TJsw/fKYGOAeRd2J+CY8v3LIplsOJkG3YU7Jo
hNMr0pPyPNM9xO3z9m25KNrGN0Etdh3/WFLfw3iXtvnEEGUmrcp7dnTm0YTa5gZm
Q8PUojLlhVmdPl0MC6e8mwLxZrHgdKQ5Ss6apPoVP1M5VZyuEDmgiVxaSHNR27CM
sV9BXVkVyx2+fRbfRAQqQDQ5ppF8XfLxS6+KpMLNeyQsWN0DFu1wsIz8ldSpC5YS
aD3NCYtHddC6jgkGkjCtANQlrD9sBXvQqGEldskU6KtXNQW1H7bjtZ6OZqghzA5l
0c0cC208Wd/vv3OD8EawbAovPm/ioNKRNpPmlL0XDD5gAJhsuR5KuLM5WMPsNVSz
6PXvS8R18QByNLENJO4ogjY0iZBml73SuT925AhexLU2iCPeDLL41nkMZIYLZnPV
fMgJg39594dBlKsN9iTwuBQ+7v5QNr2sCnT/FO1CpyYiRH40lzrXDgAXPp899MvC
aYj1gmkHtyKBDThSt0/4yOVQuvbdIaeRAX4sP/G4mpjeGupM5dMlx3Ich6Gs5NOS
enEepUbaKI90H1k9Nu+iWO7nqEFTT5ZAuAUBh84mmN+D14uU0AV1vvStRSCw0pHr
AS93YvorAXmJJMZ8zG/KwddrxqtI/EcLxwDuEByFZ7ifO4r9xAJRTd1GrYWA8ISC
mvEzT6s20c53pWCyQVkKWciX1nELCTdwMML8kILuJCGgHqiQDbhnY6ySSDiqXq3o
uVoH+hs8/xSTe1yk9T8UKc8dY3IVRflcbJGdVMyti13c2F0JXHLDkQvZTUWOvsYk
DFg7Am+Dor7MOLF1jVSUEbcogpBLe09Qd1pTe0+og13TajjUpI+FGo2DdBpaS/zh
S77MWk8tJh2QGP4jebUb09hdHfxY9um7BUfWuVME96iz3kOUaRgooN8GJumeDgCS
MQ4hNe9Hg4wPDE7UafBXr+UJ5BCPgQTQIOvw2B9p24S3pR1ltJL/MhB7Z/muum28
/oPxpLeBD91lOXNzQuY6mmL3m8dgjOe9o4jUPFBgYGXEkIQyD6zo6enG9IKf/3Ua
BRPfgFr/SihxYzBZJ9KsR/78o1TxvRFu05ALkf9kkUR28k1eT2apcOAYrJrrlUCv
J64YbgxHZlKF7zVMhvOHGmrT0c5j+QoAFxlVDCT8MYsWbAdndyJNO2VYY0qML6uJ
a9VDtADkRSv5nlK/qhXJgRtSGNd4Fud+18nxsKnqPMHakcrYzgjBOQ2+4LVBrWs0
alvRxfdfSuh79FPiaQuE6hfuxDaP4huVhgyxd6Oipo740LNesHgadTGB72z4Vl0T
o8621FKteVYV4qg+s/Ao+TKbQkAt8rV3kifLP/cgTh5Jf/1iM8x453uX00hn0hr6
dwpuN8scPWQAO/GJ7wi0W5GiaVfAgCSYW373axnPM3MxkFKdeafGCktzUvyfdz7S
Kx2NMUx0jfghbBQAgNlXWdIaEATKFRdOhVyaETsc1rCFthfjqKnZF9YlHUGFvJlF
fn0Qsy0ps65fFqTFI30C2AMrk4mvaNNDq+mtjAkouGPM95C81LIhVJCrpKEfdasi
fV1626gunsvuPhelEidK7xOrJ0T4DZgJa+23ccx6KXNTbmLwpvKJOTj4uVTnoqAo
gUpnEb2k1AxcQKNrygeifiJF7TbMIT/gTYLC2EUN1GqGVEZSQiV1zjlndFSG5dY8
bpX8nLgTl+LrgVd5C2pZXSnlBdFNIwmgz3JejlfTO2coWRFYzO6B1hH64TxW1i/0
hLTWd2M5VwWE5YV98oUfGr4N1DsVFqUsol2HMlh3bv9TZL2fUnbT8/Jd6mt/fL+h
vbzDGRjWTwrmfQ6uJWSQjg7wsCPzSF4/Fna7dKnsqmmJWjR88R9ABzEV7QUmYG7h
1b6YsjqrPdBPtgqOpxI0CNSDnXeBfiL/urQaZpT6kKZrC12eiNdaK3hWQeimUv6V
emoL5bNROIO9TNUH8/YtWbiPy/8YpH5WYgXzgN0Tp6OOJXl3VvveuDFt1R8M+QR7
DSShvYs3bhDmj0Gxz6qX5Kj0BjnllKVG4wjs6tdLy8ayakGBqB63mmH7ScjQJa8x
iAxk0vYPV+vbIJGNUeW0+1Y2au7c9LnvHaWhwX7wzECWboDi0/QRJ0MPisbGY5SL
L1sQAjsfyZUCKutZS4QMZaaR8CKY8VtgxWnuswqNBr93T3mie92cqWMiejpxReZW
NbAbkj7PEIaxOraZQ/M8xVzgT5pFuqagOhogbUuF4eRH2jN0uv/w+AtfIoqgiS05
eMmtQxbycGZ7h8/n0vKcr1J8Kyuz1reztPy+OA3oaaNfRw6E73jNERKm9CUmbCDC
TsOVrntbfGKs1i6E/LMcEd5Vnl2srQ9A/emTT/g9Q0oYxCLNpp1yUYRgVXARA9hY
sUfXc7+E0z5pmWVASH8MkNDqkQQWYtKipuuBU5WyBgIYjjLxKejTDFWJZjKKtbeg
WT0fxarzdtdR5KDAau/AGV53d8cBFPu5E4hHK2xsFF+0hH3xirciDWmoVv88Nvjq
81R8rJkpWA5K0EH2xw9dyxggSdY5zkiFPEiUyUN7lxbQCdw/U8v6klYtgWLAK+MT
00hrRHrjB22kNDftVy/tqYo65eYYvKnHoN0MX2A91WW6tA2teBpBMqMLtcaity6n
jdc4Z+v4ouHDWJzOEh47LwzTrM/PKi8CaUKUwKvcDLS4+v2pwMrQUhvklomMXgy7
eUpB39zE0oc/jFBJXDhAKKz8wghoMBk+pN1H6+VmUwYtnv9mOqdEdVvuEKXt3CfU
wHA2rr8NM6DpGp90qXqBpsOBG9PH4po+QnF7Ewi9OTeUnG+ritf9u0tH9m0DdPKk
/sx6ltLNIoZS/nIcIIN9FnEXR3Z8zNjq1KLs/cKBR446Kxu0HMkbrrQDQbtyAAY1
2R52DmnFFgA8Uk+y5RWb95F1mkagV0BTgG2c77EqMTXJs/UKuevXndHDDngqLo8o
8C60dyghGe66wZN17Zz6AP8qCXxl96QkEP6FmDf5rk4I7FIGj/G2FCqtq7J12MPE
SvCFye3GjlLxSiY1zlQQ6aoiy7Hri8oDb+NkzJoMLATNq4DZ0Q61PzUxmgDiBzCF
gBjp3+aZ0IELykHQY9VsQbeY/xDwJ8Im+I4wgQ6Epa3mE2hWzNaqhwW63xiRic/C
75GwT8M4pLhVNC2a5lmHfVRTc9ia8YmbnYzABKRU+ovKZEp1wqcS/vVdxW0qYafr
l1zVyuQRH7ckK6OQj33nsnrHuB559IA7b69XhVcAjlb3x/Vuys58O0TY/lByKWbw
dF1WUFRZniwqQ2yY/GyiNEuQIbm6AZzhpm+r26Xey+dvvoRaLQeDnc/sE3OLzdud
7mbbXvYEgpvphTd45CeI8S05oTRa90fy/BmTbsEFVyGLysXoyofCwzOIOEv1KE0a
r21kAUG1pAb27SL2GSOvYVxjDzynWWo6TwaS/4f9+F9xfjC+s7rVTIKPuWkiuf2x
cvTHnMC1LC4t0yCruJLC8swj0NZzdnxbi8kPfJEXpHdDgcmMNKOCoM/mYAQjKknm
Zd18rzyLf8ku015wKXIg+h8GD9tP5KxUfQEqS0PKkTUk5O4Qih8+o7zoC4tI3uSG
0Or+1zao1snQ03IFfGgFA0Wucwc14iHd5aEXvlfKTW+3Rn+diqlX93qzZniI5+yN
5Z0iDfW2QIv45D5BUWDAZhz+RhghjY/mOBspdWLQf4hpWV4bkS3Uu2olrUhDcTuo
aTPabXEZHQ4VVb968ckYJeS/RLhXqgcZNtZNaeWdh9rVmT2ae7vwLW3fMllz07Wm
ix8FHHgSQp9LyK/e/tcCBmL/YKnA0jFc76ANGjQNhE8QVnDbpB7qWE5WWsDAKjYb
nFtB/lkx2PMXvBud6+i7In3gvcMl375FU6bUdmmIwMRH25bjyTrd1RbN6l5MIWZb
nRSssk+OOl3J4z+LIAd5eWBSN3z6xqKgqEB5yOZYo0H8g3rDyuvJYykcNm2ivkbv
vz93qQcDvhB5DRxxlJ0uZtmCzuUKc7+s0191ohx/GSkk0AmSW1mqHiuYQHDCTmPT
NiZM1UcVLljWx7nbmm8bXMnVWwMGlE9hwHvY7VTBv+M8XEnoSsUjrgpGIjllB4Kr
iZxdS737Ml/r4fZxwEgCB1pUP3z0l9yFlr0HtVfTFU3rSRTmk4pGxrFsw2bNl8Zo
lHfrjHRAKzL2ptt5R0uzWn4ga9qslVRxvf40xdtfS7vEed1JoGKJD2kx2Zf8QX2J
UEC1RBSFPI9lkYNAnyhzsJICspBii4p3LuQLiV6w72v0qckn68WHFZDRNvkV7ULn
pXvI/gmsIfTsUb9EawlH2WS1x30D0xgXll2m0uxp2nOewLo/92Vx/aA2ekJcUWrc
GCkb5/mb3DLAO8432j9hALb56H1uVGl3dvujYoJ1GWk3d5XG+lD2Np2jGPXP25tJ
qscQjmWNHBZ7qhtWjGZx234Kkti+RQXOcZtG/RjUagZVzhmKEE3IqDdGg2bKSqd5
rdJsLwHeRbw5iaXRlAZKgdZ8UQZDYb5PUGjSj3AnvaHs9eK9Jj4KrbvRKwunTjFn
7ecrs8oq7qNM+lB2knnKZ1pkc3ecoytz8zz47wxTgJn2rDqmwhRLtJ+42WkdFrXp
rFHj4njmbDBUzvgdyRPVIZ2SoAJVOFuNDNOY1ir/4+jDI6ElVgLaZyMoTijHpcQk
HMP3wYFapAdwaQThuCOJLrljuGLpqNDpca/RD6Er78/+SBinS/+tbfjtIm2EjQWT
p/y5Lx0KL1/Myovz91+vYMTw3DU+WUPDVOSyakx1QinpQRUy0pUZR3nXewY/HKpO
G2cleGcsDxyLUd+8QDAp6hW46xGAsY8QvIdbFdCX3PW3lUcjaLJBLHbxP5ZCOo1p
KuujfwTuEFx6pm0LXGsrJhAbaJalTVcBsKjhPjM5xxfVj80Dr2T1sK6b/oflqgo3
81ddrkd9pO2XgndkwLUmR/BZne5FapNGoMzuqMzaDEvLp747WmI3iIeXy8cRMm7O
6qgJVzCW1rQLqp/JGdIuOPnHfRiKrCEcWAm39KUR0vhV3n4zGY79bDrYM7HZqqUA
AtU0CIohJf0+bbiVj1T9UXeRJNw6OPO2/qMF0LsONtDfo4fSYbrMrUOAvyntuqr/
wDw7Z/nztEdAoLRvnRqEEAHx6OUG3/lE7aqkrckulnixj82OozD3dipFM0S9syls
ADmpNpAMaQCkYmxIGTrBWPxaZJUYSq4TMljWAy0C0jWOMmiuRVX3HQbkE44ImSxG
SAKIMCRHATXQSQZAo0DRzsTWFSSVtdRD1z/4Zj4U72togIgSnN35Iks4AQGQBKaF
PA2c/lJnLN1apTWmRPXL12gSq1yAoBP8iobnjMRRLkOshslUcateBIAwKKx/vhCr
93uie9YdVbyGjJ2QHmYPF7LtRZFOaxXMQFshPCB+7pzekAX7oAiedYTDnnxnrsqX
Yz3DUnuUwrNFgyzz1dgObnGIMr29wYMyuaZf44smhSAMH9z7fbFrFo2Bufl8ezpx
/bK0VM/5lPeucSigYTd35vQp8Ldw6qg9Un2bCCyZV6+/d/z8cBKAA3yyiM8PAGpJ
G1+5LWoPMUTW4zGzRLww+4tszqy9Isj0xZPjqWarHIBrmZ4fZbLMDadSNfvo6ZcZ
aUaCLMheX3w4MdBq04Fpuv7aHAxTX66awJ6TqHbGeOSM5R308eWMGGbNhqtRZjcV
2AV5s36Dq4quW5XmMluuiJkhFz3MNOzGwhebNh3WI3OlU13fzWyZ8WW0fn6KgaRT
b7M5wJE/sFIuI8C/5Sr1oLZ5WDgc8a82Cee6iFPFww/IHOZw93yWy+slWvVLdN39
zrH2ZMbmQvdjt7u66biQ9UCUKOlyYHYTGQ5mo46xCTsrKHsEyQlVi/xFAb03EtZW
YgkIZOy+mNv/0kMk+oz79uZKo4ZfR1hQpZz+9HOvn3fQtrt6L5rNzdRaNn0LoIa/
Uxa3FNga6nI6XOt2R5wOQyJu6NKnPsP6dn9YRXEWocZhBlOb3SK0i0N+LEn9o7tw
bpkB6MVew93iAenZQnVVWaSsKbRJGuDf1EReTlWPBC2G0eudTwFzhTUt7HglGskK
qY44xtbBrksigv6fNi85+7UPJIX588qhrHQgvm1HYEIAvSFbqv6u7G5kajyJK1qQ
k2ECTpMsBya74Db1vMPy6GqlMPwQG9C1496rE1rqShPZtXl3B8weHqyXWqDeb4cV
AHLq9j6gkYD7C2fIR3jLlxfa2Bo5qJDAsFENzzrPf7FLnq0LPOu4Ndl+5yHPVBtE
lZzK5EWdGEWu5F69DIpT3yanB5qYD6RMu6uEFCZsobVA1txk12Ku+lu6PvCBRl/J
Vti+FJyma3Z3sEpGX6qJWaNXeVFlJ0s53grtVkIKu/TdRIhODXe6A/cNB0wSkp7/
nMNIY9kFg+QR3qnzoDkjCa9TqYhDIf4MAcnXLqYVH3kBGXrc4rRHHmlWe7BGBDnJ
HRWPJw61ndY2zHq4yVTg1t1EEUcmi+sgplnMZjrbgZSCpBYfSzxKLoengQecsZk9
7O44qIvt/CPZV5O8XQhP3/holc6U68Voib2Clakse8eLQvCbWVQkvhCXnDVZskf3
AXGGXQ1h7PMij4VzV0ElHrNnSE/D1qcfniKTPZxqxBkUQMm9OokIxvbdlvG6enkJ
8eSJ3l5uYZac9xgp/SdkAlMkYX0PVWwh+4aWN8KfIPqQ7zebRvZ51VJwOvnl2tey
qd9izlwiwFio7QJZkObFodsQ9TPDDF7gDUv/3jcUSiHSlbaBoobGKLGQcAh/JztG
+6TND0c2XLTxecyrA3K+w+Nvkro3M5pfqIyiBwKQ7XqAyj9r+jxCGql01+hb5vw6
Xb597+8GVN13+5xYRYVzduVie2B6JCg6BpLQ2ryK5+qy5bBcw4dlW4qgbLnZST2k
uEFqYlwhZlQz6hTVGBF3oNpeme+gQg4+13Ccsk0Ef50gZ73XSq/dMfEcqd3pzQJ+
9Iz7JrMW/i6ivQ2GoqSoLsH0XIus0/1E9q9oAgqejt6JPRn6Yc16ecudrSlqK27I
rloa1HrzhXEc5tNwKG9qcIchWj0SLq8yZ+CSIDMGf26fpsfbLY3vlJJ5FxgRawrh
iD2pGbv4KLYn8zU5REHR7AW/x7d9uEuDCR+YLCikOrFIPZMi0SijzAQ75bk+2xBG
IZ8PtPDghmrPIo6RKdNdcA1IlLmPjWv75OSAyKsJWRFKC+EzXE1zU6DRg+/zUEQa
8iwrKzVIlbglrzLvsk45EABMHnbnxJu2yQ8LEgRON/LIYiIlEM0hFu+3glF7pI4J
9E7AhGSA2+xPFGzueUXMLrBGU7/w0Wfba1cAdDzvMsKJe9P1X006Rn8hDwxD451v
5VolX401ZhgVh+QJDC04U2lYUjYSNwMWE4ChLk0vfxSa3z/Xt6IQsFVyVzq+V50M
2Q9k5S0S7GrNzis0Qab9OnYHHpK8d/HY/G1D4hgpEXkYqxOTeATL79Pe00u2QyBY
YxkQQH6ih/TtLO9UHgQ3uuKAKEw5+fb5wKCxLFqH7iSoL9WnYxiOF2i6TpRCoizA
0OnxfRUc9ykgT4xUfn+yfZauTWNOJ/N478Mn9NLuwQ9gefmswgqXFc4HcpT/u7vQ
4iENffjHuvzDHrRn9v8I4aqFGlSOLosuOvOgu7MGy+/j3vf3Ke7sQ7bo7+a4zTd3
y/X8v5SFgD6neQr6GDzTx0rypAPLJD+u074mCX9v5y8kp7Du+Gbx48zQ/nld9T+K
sFQPKXtq+p9Y7ouG059crk6DiHyfJTTnpQLDa8IITNPlVEvwNdQnY8MmAYegPrzP
ERgkdXtOIGaMiivEb8pPdfsokFida6rz74hh9tf/CD1wCdsoKSjl8nUGzuBp8Iai
XfcCtaBRkEr/MWOckjXFlHylYfN44GvUHB+QQHqta12BS87NNA5rpX5i+lD7HQVd
DWXZXRxR6QAZB1Qxu9uNm8tP1KfMluvo/f1dIRqVD3UmYt5Oofmvm+ipzBJY4WHq
kDY/xhpPfvqYWhSyWSAY2KKfy2jXdO7J7vGckinOxNdnebFb4Adz76ZTdSc+GTpX
Mhq0wINqMkXWIKS8NCIeYcTGqmLs8492e3GeFknPo3GtEFkULxXXEgx+sMCtvdYA
WP3M+OY7uR1d2l7BTcfJSm84tv8nKOzTzaLBlUZY4Gj1P+qFFG4gtf/UJpN981yF
6upvU721TohkBF4c8Px7RxT3xHixn2G/zCKFNbt5/RDagkCKEDPMO/knJf4Bt5aE
PSbwH6XOq/yqHbePUIzYvzViVom3s2B8aizo/66DuHUrhm/V2SvFwqwhHXxyN0xB
NnXYWrV9o+vcHgRMhII1DidzuWIhgsCc3KJ0WxatQ9TmA/kFSIO4fFsV5udiI1LM
kZNJrNwMorOGN1UFEEeiQos3Tuhd25HeOppl5tuX28tMAtEkG51Xnd4JEJwixWl5
z7OlPqHLV6XOopvHFxJ3qoVE8JsU8ff2006RL6paF9Kw0XJjYXM2bw+67OoUzw3h
dYOGbQc6pkb5g5/5hnC81AStDZ/SKaAJ72XSwr/QwXz400SqLT+JE6Y7pVSm0jTI
H8hhVlolk662kftk8a+LixIqLLtScFr/RXtGjrKmAJTprpPBPmpyhLlGEQ/o09bQ
cONTKbukaFWcM9HRVzYekQ9Sgu1DsAJD4Wu7nwGLNDk3QXqsqW5nXy0+6b3Dj/VF
lK7WXVC5IOPfa58/k2xPdWLlFbPdNhJFG9G1Yltxe/X2gKOFYL8kHY1P7pvlrdFb
8J+q1A+y3dxeDh7SH+QGHBbo0gA3Ky9pDB4cjJ2s3xV9LzKYN0tdKZCUrwUuXEvp
drKG5ySDNn2lcCdosySDA2LVafpIVf/Og/TO8u4gJewELDVpN0AerUgFK4jw9h8G
2gwbpfq8bMqNJMtTTeDfcgYrqlMkAfou2lKb876oNNW9lkT36ZR/q728HDnXi4cb
ukIHQadChmKa/97dHzZCgsaPN/+6zrPufyyR29Dpc4TGDbDwjTgGtcUnKuX+3cIN
p7m29EqXM/zS0nHrpiTRY0WKIQ1D730pJk4lvBtW8ACpBkVNfnd8zDgQCU5xo1th
48nrHCsM/pQG3Lg//2vh8dKmnCa1DUqlm3xgjbS//hq6MldbuLzvzhDzKyNwrgvw
nlZ0lbeY/7+RpTrSbN6djH/PSAR0xVOqo42jo6vOIGZchkrvP76SlIp84drZM7yj
fDWVDZ9sXqw9dnl4jmZOror+Mg3JbH9qtrYnIyEP7tw5Y9n4+7VQ5ztiTrxkWuyz
tMORqxMhT+RnyNZa8GdJ503FEfBSDFpce+lIYlbw+bakt7G9NKLb6bChrvwsbLPQ
gOVfGx9+e24e64Ov37mODzAbdQzxrqv7CiGh6ic3bAlWU1KVGl1r/aDHhE0iHN8D
yHV6+u1JL4WQYmoLChhfI58Njd7ltwKwCXeRIvKqMqRSASNyTRZrsscNOToUXMBy
xWg3a71tB+dQzCYapbxTxCTo86R1Y9515rXf0MWlTPvdYPrsQNPm7S9pce2TxqvD
lJPisEun+OPQAUxAEXmzYqIc54jQac9wSBhTuBJ7W+FrfY9JtlPTc+RIh4kffN+i
nobs0cQ6K7Jh9dFv7E6c6cDM2wcDKSOvL9YpvJHyrdrXFIwPOg9qkyPfhWvMi9A3
AcTiN5Su3ZWHFwMKCJAIRKq9RStkSzGZcRqAVLKZxhwpnhUNYzi6FTcUlMDR9WQx
HUSPnXYWkAITWu9Wv4DkzzdHCqnzuCYv4qXqO4bYZwnovrfl371GUM8cryz5T4dk
F5BS3+MZTdqVte07q5ze2l9H9Z9jOLqe0qu55gOYw7LndCHWZIlXlghrIifnsbL5
WPtzsq+MnZMkFUNg67yFbn8ZgpTC/Es5QGO5/hC6g5doL7Kchs5k2zmRobf4fM6P
NLUonqXU5RaO6xgHJEOOyU2+Wkc3DlztaPNVRbZKRGss0fnfxOMjnv0BtW4Yd4O7
ctCJWiNgOHv00/SmdTCTdOTQnhPS6RG0YqgjRZ5H5JuSjILI9GRlrrylPt9jNvHO
vfSnIwZ+VwEblNVQyiJb5TtMI+ekpxt6VEpvXZqHYB2dmFAjPoAObaJ1i0P4yJ1O
jabZiOBUq/IEGrQZNp8hDx9lF5SgsY2LVA+d4KPReuekv+wuByx6KZBz22MF8VE+
1xs6tQWxLCl/HdG0JDAOI2QrzkQZ5FhkoOYnr8uKGMus/39ShGDEPUedzYe5fXWr
6r9YuoJCIF2cefy36UB5vQsqiVp+DDlKrAIWqexANuHIdT3mUSCnc05rC2bLHB1I
NF/9rzJfU0CfuVhsiY3FXUFE1xYF6RebiHEIBjZgz2/YdpHRDpau4Pfvo5HFUbOl
tEWSwSaAVV2FllfqvPnvJQsmuoaFsUi9uDqlU8vcHlHDzZ78i9eMmA2wzl+BhilB
DD3gfUspkfg4auwcYfcEV0Zq2fRylxadW91JkxS1TiwlHDdrke0TquRfP52nMl3R
+u6EIdboZTBfp6qxXjPL29MeArqZSxlafhyUuxnloFa0LjOQjlm0MNoCDzcaSYJ4
/xSTGtLQEnMD3yk9qgzWxTnxlL6/cMq69zVdI4e1ot2ZJ9JW2N0MtShTfq2KFqms
vyxHH2X8HiT+HjOjQH4ByP0+jCkQL8PQ2dGDpSbfjeCWvB5UUtHOR7QdUpov5LZD
NeNdkoFbuxIshJzR7+bRNCxyuHBApE8qNsX1vGQa3c0ZIsxqLpUId6XMJN+PKV75
XtnZj/1hWPAlHAv2Z57GwUR/a6GK7S73Uj2geUKKoB/evvBgmc/Nx4UTJxQ0vhMh
FL9+piknmrBGTNLTKU7t1RiCwNgOof1F8aSt+A+jrJnMLustPo+/bxr+VotIayRL
5XvhogsvZ3gvLTL/3r/lyyckstPSQjnYKyCyfiVSo7waj/EgST8uplXg5MJA3x0o
keuZYIatmv+MWN2hyn0Y8O1OxkE0TnFxTnU0MnlrvGhhi0BjOWjHzrJ4dz/vkewo
vlOY2UU6ql3iO6GGiKKyurRj8L6LnWKjQfOqAlUta/tscBfLRqRa3jRl25tkXhbw
k/HEO3v0wvPFngF6mT0YD6x2eTHGvC4yjsu+8gB7vHmvl7V3C67r/q3dJhKXF7f3
twaHGpL7o+r4ecpP0T1ighw0C+zD01SexcPx4Tu2YGeaGTAWafMkmNERtlukAO8C
929z21MqWRoMqrZCIoOiAlD1VBM9Yj1loZ2DEO8iqzAybMaA1wsGkfObq3WD0zdB
YwdBKQaqozG2w0mS7bz280TMwB4Xl4GQWgWflSQUuzQlxAJ8KmLEkCH4Wm9Ue0Gz
jt7FLnm5NkUHEcnd4nLPD04m345bqiBi1BnlCIQ8qs1b4pCnPGRyACXQOSLHM+dF
XCJVflVErXT/UOcKuOfqIK0uk2ZFAoOcyqbnRS7y1UFrroJ/sL+oF412UI3gKrR9
BW8XZJKcjpV4+CrM2GZ3nZaepWdo8g0DQnELbH2o3XFwsZ/3GBJhTDHJTTSiyTMU
SHKBWC7WExsGU167NoIxg3qfsNwLBvj98RLK/Krw+3SI9bx2bMUUPCoR78Zjtvla
2nWQZq2QbqMlseKzlINFHQIQYFuhsXjZJ0m7gz7I9ZBS5ZCmw0v7Bl9MVmaQjCZE
k9OPbLvoq2Q0P+DQPlNNPSPAI+x+Sg+OgN/z+HCyoU1p+iP2RRET8h/g1wU2KnFU
G/pvcrR9pjqZZ9jyFdxC/IDELdwhM4UeD3Uw9R7zhkp3gk+4kibGwQ2v2NnZNwJr
pksqb4L7ul8CrdFY1/Vw8lzc/PlczaoyPBO785PZnfOK1BsB6rKMl6tE3I10Kyfg
kgDTsjEUSvcjuV+tYuuZpSGSgxGs4tlozjbtiSf0E9DfK1eulsybM8B4sJTvhR9K
EcDUqYsbf2qw9M/e+PQ3Jw5dpGZwXioO9pmE/20aVNYRH+nDIghuYJnLFfmRaU7Z
SQT1keG0VeGYjIKvv5+i4MiaxVlAK+rAMxzq5hDYEgZxYh6fuIlAS5p9Gd16hTmP
3Xh1UcDMFZWPyE+1XJOn517aTdBJm2aG95b+CBmckI2wH5vVaV+WHcf+y06bsN6D
KMXG8/k8yCuX/IeEi+x4ZJowtmDWAIlmKnQdESlw9Chp3qCI+4N+9Picn1i72R4Q
oG5RHi9BNAgTDX2pegDIKgWTLth5t5z7T/3LXu491p5jhYYdRtkk33hohVSJ2bfd
M7uIZsTJTvLN2sFD9JmMBNOE/NdMrbTqwlXoMltt2Ze8ECxZYG0vn5vXaq8QIxqb
fHgtPIPZFPaoGJ4KUcFPF3CaUblYUoa0I31j85OiNXbhs4mIzG9NAuP6uV+9mMSU
ABLkYgSGKR9mFANf10tEWmoHjCf2PP9rM2S1cQ2Tf+kOp5P/+IaBdt/o1Trv+NJh
5GsnnFHzs19RLmQD2l9azbhHX0UNQTkQwa4HhSqoUOIx6qr+7vKu8s4hh8vxVq/E
EP7olCYWKwMtUyncTT0mAR76W3MBcTOnHElRZlnYHcRI6YjcVSgt1Q8UVlB6J9Eu
BhLksg3ubNA1/6nt9iQ4tQTlC54pzV+QBxHU7tSDyZN+YWAs4nw5fhKlwbHnYWsM
4R7VRS42ht7+g5v7FM9PXpm1R6nFDK347GBh2IUAcGpIB1zByXEAjW8vNSvx0/x1
4bpK8My+Bg1xdfbq0srhCgZjdTwro29izSJgXOJXOS129ydagrotasYw21j/LYop
3aLPoKShkuyPIln+nUJnNBY8IjclQygNEURqrCYAlIw7ZkVj+NUhJvN20Q3GtIxW
ql66o2jez27Y5j2esv7O0aKKaSY7rlqGwHQ0nQRtq5NAXA4D6u4HYjfMzkpsFcTf
MYqrA6ytAOo1v9R59TwqFp/VUdW6xumnr+UxwOuSWmfXbJYv5FA6cVKaFglR2eAP
rAveow9vI36pYlwH/UtQK8eTIkTMQP2l3MwjMWpEgFzBSoEO9hW3UgH1kTUf83t8
SOW6OgfcziwvwC7JOwQDGBco2vNuOhuPEkiXGCva1Wu5VxB56dCjYGCobLAwRBz0
mXxpaWI7jyu+kwJpS21PpgXqmA4lWQqX/Ft+Mi2rr+iN717hKy+JzoYvQjk1Iefi
nM9bb1LWAHLq0R2KMsS8XtmjVoyeV4v+J1fgaw2XwjoGCTw7gwyD0c7Q7abB5j4c
RYDZI4qhkhswn9mjtFeX/W9EFwZtlIxpZ59PoqKlj4V06UjRZSONLMiDYc5LX1+b
CqEwIqhhhCGdw4Fg9En/qLL16weUOLFr2uoVwfPl791WwKEF6Pa42Zpps+iL/o4a
qXcwg1+mnD7EotEK7JotuYzVFcKuJtQ//TFc7JIaXr2Ov54sW9vBDQZ3vlZddo65
MUuZ5Ul7aAUIW4+vgWkUy4zpzws/qgINDWro2rAUGI9JtT6iPjA+CA+oh6inLeGR
YMEp6aEPpkxjC1VHY8bpbJONV9we+z7PRJ9mN7rYcp3BUOuCrXNTKy1UtXnFKHOK
Pb6Sqoid4l/CDWYyjKp8aXK2+lNqjpEHThJ5XOkNotQkGV2aEiQeFhGqkCEtlw1H
TMwg9a2oWJ4V6WcjdE6X+A6jnnCNukehHt26GhrVFczr79bW26bpB64KllOLAA4s
L07sCxw+3t2lenUqT4/y3oPTbWMan6VdZyedlspzNfZr9IUWI/oez4gTJ35/2EJY
Gk/XMemQrL67xJKHQ67R6NTwseAkHiiospzaIvtJkiYOf9WqrJ9yi8xkQKOrnhgK
wDgp+XnPLP6Ne75VNWrvvKSi7YGHuS/hsDRJ1BE5rN0f1z7RBNxS2FStjU/rv6Sl
uDm1qkgUDHeKNCLK37v3lElt2Qy2j/xf/5LGB2GLVVjR1PFu5h8a8Ju4wEo5/dv9
mmeLXM5D5emZUyLluGHNd8dbW0XvdsP9WUWVB/s2jANP33XFYRz73Sxeit76ed19
LSTuzsouQn4fNlCvBplW+WJyPJ1+2BM25WOxK8PFlzRb8cXldf3A4PWcY5S/SGY8
rytqmyjwlb5TipPmHbvFHKJoYM9empsjClXWIzIpbj2y3qGb4xZfp8YOG2Mw/a9t
CaHaSdl+49lh+wpjln8xkAMic5gk3E4Kigiwh1zIoL14k8H290r8OgCGoPvTa1Ju
1NWj2NySer2xDf3FKsVOmqc6blO0QwIMNUdQ2a7NgRhlIGBbEYOsaOqVveizn27Y
Gj+waNuVJQI6ybAdyyho7/na7ZVE7Ldebz/0qaNHUtMTb8kPqgCsiOpv4ukFuFlA
fHU4nukRqUe1pBXl7C5dphjgamoEhyZe9cDqBPaJ6Srbk59uQ2S5zZN5+0nkwPM5
dJfWlhUWV9it4RLFnq41pYVr8CVVmURowdTvyFoC+8yJL1RaR20Chppto6jP/XbU
5iEzPM6ByRKqj8tSKQah2r2NCFGiMyxJqY5AVgWYa7iHsVgfr52GZvcNRb9V2V7C
xJphS1qKreVD7LTJXcx4n7NeAQPyF1JP+7JcXfYBga5LAw2zINMRDHZ0EayhiZuF
TBVj44zGyN+PWo42sxozS+kkVmttaOpMqaFI23g4/ouZkRl6HIamXTwWOq51PDYv
mvql1A+iYYhVSVthNDnVc5fOJ7FC4T2jx7+Q6p7j94QGTwwtYTagsID07urqqhAA
0PhM2MniAMbfZZukicmJxcT8wJ0vWGDFjzuyRmjK5Fj+hHcITr4Y4x7XPbSJm/vV
DfzbQ0ZQlzn4ybbI1oyTE7VmRoi8O3JQ3ZwIntLOAvpVRl7G1+mtij0NluYrGIYB
RezzTcxk/SObO5Em0pJzcx2UUIJcEc4LYn8/fZzlwGSKpgoJsBxCkhgEi4iwRkKg
OLhkNrwlSoqPM8uVpYcXcg3tQN1hdx6j3HaXN37PeSMlqD/u9UkTlhww3h/DIIUP
iUJDvQOwTywQHZTd/8xMChS8nHgYlYAgv9L7RYDHy8JmsWgLiLO7JwxineQ7dENY
1/DVetAbd47U2mtBzGG9i+0XDPJmXpIp9ZWTcWFafqzzLcjzKKijsYOlQbLnK1ui
CCN8ts7KhjJRiKCX0dJ5c5zCcL1q0TMQqAz8fjXCDmA4qvx/BBjjemG4g1epIH/p
E0i/9Mp4Z7kAxSVDZ7dnuEW4yjvqjQkkl5qLnYmoSAY+rusRaJC0Uuw9UsbrFIvp
OIEX4cxZBWa+iXTJyN8/wSwJuOsx15eFoTRyUMOBeekbA0nte1wiJfmQhJTmFxL3
mvrPgrr+ibj4BOMtXbhfI+ARyz7i3Az0Dsa0hjbRdpcQCDo1fLPszFZQ7JAAsJgB
LKa49z5wd3yfjtV+tOWjjDJsVZ/MpQM3M0l1xg3is2+Q9zcxSgSK6nwTf3/iVBPP
Oh1aa7BEEDpUVELpuUzT6/mZZQg6+R+Yvx6JGFBqgw2gDoXUvanZaDMla3t51rNe
Dpul2sH2F0C/dZnthaN/8y2JZWbLeM/6poyMhRGdX3YQZSzIBKKnatPWoQ4a2c3u
xtyPfQOKqYneaFWJZ8TiPzxA/1qH6QDUi0kdGSJcB41W02s6SZS02snAb+TquZa1
TpjJzUoN3XQnziES/PH+j3YIFo5LHEHhm291kHITOjCJh6bGoxtKLmd46g0IJjLI
Sr+pqofSinPUO2hTBeapqw7CJxs3ZrJaCVLTSQTUEnzQYJ9xTQqy3/OZ1Pw8q/bQ
iXhh1ZU0gBnUmiQ4+ZQgrDFBM2zK/38GMYUllQcUtmtKHA1vor2rk9YuZ7wwPiwS
10X3RoFl3seOg8VA9ygXqvUci7N1XylkXmtHQ+cMiUvRnC9ENqjon9dXl/tch3EB
UgPbqrlfD2KPXFHPVz+1GLa4Vi2bhrvQnaN6lCAkmK4vl04cNycWFSikyqja28Co
NB7dIw8WRy3JnGdTbgAJgdxXjMn44Non8AiVblTu7Aok1M+9U7K7g6w2Do0a/Ji1
N7KL7kgweAwsbveUjj9q+u0GFsDNTOhylv6wH9l4EouuIwnJUzCBHG48JyXAo9OG
3rROfl3wO5HaBzIkNrxprwX01Fctj9Hb0+yXl5eBqQFaTSBPdzxxKJ/BfyRftom/
hDM4HK50c60eTjdsjmd1G9z7zPLOQ2nUwkaqVxtPfBmuAapcvgHkcl7+rbZzpE0H
OqN+ecnnrXQMtDSw39gNWVcZXHv7pVuk85pwRE/csvF1tZvJpFu5b4VaP5MB4jMA
GkGzteGLjhML8g5d59/B0rBWPqkZDJVF7IN7JmMJj7B/WwCy2mQ0AKkc1PEcobUp
EDt1MCcOJpMpr2Y6uvrWVqtkauPe+9RXP6ELG1txfECfydQPKhyuZPrYUOCNZe+R
nsdGi9SGOsAO2t5a3I67YOciDb8veAyMiPCVh4JYMuUabfcd3TLQ/a+0gENs86dE
UJj2sm4mDDoscx5NEIifOskklwrAEABV2aX/a/X9n6xqDtx85toynx1K8+B9amMh
9RlS2Nd2r61w9uwpXPjPvTxcxc68gdAKOTjRlBS6U87q5hOalnXv8Va+r6y6M/Zi
t8vmqgSY55SnBwoAXJsltgUR9AxnmnB7E/c9Pign57Xgj9gufc3hEXqCUEsq07sR
0Td3urcpLnpBis8jI6lP1eCBRXiC/jm+gdwPpZxR76PAQ8FL1bI48DNGU6Ey2re+
JdHaC9cq13PVojQ2XMLmjtbaKBzz9fg20bPn4DC0n3n14x6MVcV5QY4Q7eWsxrdz
Qp81lOAfeNPy+Ope3gm5xoYYow+DXgbslZB8eXPcT5LfJ9FJT5gipF1lS+95QxTq
ey0KtMyuk43nZiU5OyKP3WqC0GFQrYaXm8h3uPJPr99ol1IWlegIOluubjWijIey
9b1vg3YL4mjsph6q6AkmSk0VLs5xbu46dS1earT0C0bwFRTew7ocSHSExejnQZ6F
ZTErY9umtZMu+wZnRmdDOAFmTUZ/e6f6ErPiDEvT7e0RNtU59+tr8Uu8FZF3bgLp
9b0FiS5lk8Tu2JIzE+KeyMJrAWeGCMx6vvwHVEhwHInR08d5gdYNnBYvEPcm8Y49
qy5OUAp6HPfKPzZR+UEk22xh1KdAZygBNRZEv057EFG5Gl3PE6XLp42849ZmMhfh
qAFDmXOsLe9fPHF3nkwtwRjr7KcIRuqd47nxy6BrqyO1gFpopQKWBcL/24PqimTl
DyA8XTGRsMhAAsgQDDMgTm0NDZJCyEVQubk5J8y40eTYByXOi7pqvJZDTxSj8l0i
hfb7PYtGMh7r0okmRY5taxWXGlbrxaFdpJnfcFfb9GsA0TXgf/zcb5YXATj4gvLC
IzPUvqYp/trOp8TFQyimZ3EvDOjWLVUfX3sMQNwMIq99b1Sii07B4oYldma7SA0O
va+CEEpketfq3pxXNarh5yWox0Y94Gs5q+a0RKXyR6jVYKueYpC6O+wxqMaM1FlV
goNjWt2UbkuI27dhCMCcPs1mV57G/LZnsj2sGXKBx1oUeNtWDMoMmlhSwFBvOy4G
jnMGVG4Z2ru5dluG/ztEg7+dhaG6T4yD1bhWS+EQtSk/LuPZtVgi5hD/mdn8Er4y
N3n9zZxK9AxLKu24uKRGmooGHDm06XoTIBO/1JyijktHgxge30Ng9+RXKQbSkcTJ
4dwIWLWjPELax4qSLTyvVR96SLmtlLWUGDJdMH2lgD6ypw/nJdKdIO+DVtX5sy7e
tnPqfv74ho4NwAniplIwQkPELafY6wOx4FRAax7Miws75NM7q14mmX/f1S7lgdAf
svPW+FhQpNRmHUsOEd61povAbXYB5lQLcBlMhfBhjjjNCPoKHFlKfrysmOtbWnD0
JO3VtBOgZCp99ujv/E8fH74IUe96MDDWPLw9PKRJGH6ffGEuyhO4Ju2GIatVwYom
IQ3AblDbjQIf4z9aAW4PWPuP8d1hUyGOp50/sQujS3uX6977i7z3hbcmNQV1MzEz
qG3DgX0JuUM+PvhZEMwStJnXGyzS4OeZx4Mb1wABi0lJDJeH6Q+mCqtk0B1Tvv5I
mF8oGRvGya/yumYPv50W9tXiY22wLmCOX2ztW5xnRnTuc9p17ZWB5nOcPAMhEejj
7UTLIkKmCbFtO2dDeHLAT9ZPRL9imK/2nCHpTXRAzMb4YR/cvcbsBUOM1KjetgSL
MQCstHoeZptq8N8hoNPDEEcQ1wZppxnsHE6CPRDvVCzbyyCrTQzy/WiCDJhUVgGd
8kxxqoNoV5lzRfACY+aabJJoY0ut5hYTOILyORe7IWl+6qTMDyHHM1ZYoxtWR0bY
2fZBc2wL/qZmqGsqY5l+fjsbLXq/Qd8Ygt5Kc7tC4KNte9Mkx9PmEuvckoz/sRGp
Vz25qiRQBf3OgZ9iFuC3QgYijQcAzxG9oeBuTu1IcBFLWfvCfWeaa45SSAOhQhEM
1Zo3FqRf67PmO6rt272b8aIjp7zWuFFALevZk/yLsvEm3LO+QZ3wsjr8SCam98ES
Aij+VN5Wg6LLqZSPZTtA9BoOf18SOYYMUc4u3PlZB13aCYTTwdqBbbUx0NnXFS/A
W7qR4stvSSa6V2wYGzB6jiesZPtC9C4Ry1KWMJHuwcx5de0vHWamk6lwgYb2XFBo
jQd3d/G/OTsKMap4ezyIouiomeN2fwU3DFHxbUqCgtRwif81P+UQ+Pej4FRL0LB5
yVSNC12kNDTTAar4PfFZwwj8JxNerZNurTbSBQkHFbmkKnmZs0HOxxsJZIN66g0b
SrzAoNbIWNgc1PLWGl6RiIE5oi0HnjuGcg5YC2qVox8qB3rTw8efP5eqa8e9s6tF
OqAoozhxLwhpCAizDk6EUBfgicKYMd+dyG2lt2IkgpjRkw0YJi0ecl6Vgj/Gs3t/
4DQFaK2WQIDTc6ydxVyHclvhL3QHRLyTfHUbzAAwTVN32e2xmTlZa/J16p2ROsjv
yuzlhabqnospOnweMFOtcZ0GBG/+7euZyikL2xDoRRLyzCET/KinFFtZ5WiTTN+P
TCEEeOJdyhEbhaglHOBbhif+NyNVdsCRVARI/P6yljX5SMFXkG++rU7rHDyj88dp
zh2/z+ltFT5w/V8aNU3FafRpcu6ukFb6v43hWbILB4ebRT4pWuV2wTYSrPbMz99K
89XwkVDQbApk+yqJ+QwVtcG7Wml+lO4cewh868hRL9jaO0nzuZJR3MpSx02zUbpJ
whXBW9pJCNN6g5/bs9ptOgxPfunST9PURNKQmRYbDxt49bjhLECxdK/O427dibhl
0EVKOBX2sPGYesf3Evb0mh33x+zNYUuOQI8AWYzC6Qz1uwrq81AsV/TdxAsYhev4
mePURCfLuHQ/6eTgJi0OHXAmhE/RU9Eb9nM0K6clHO/BSpoINEmPy+o2ENC/9SUE
igXV2PRs3SO1g1I/nO8SLLWCs9/+G2T1OJpASjrKURdWWfxkLRVK8AgNrj8kbfCB
Cf1ia+dIbanzpldh8YrtrViImYnR6h79exAIa/3ABaF7XYFagwsRVZXV4Qzys9q+
54e7srwkCcqtRMKhT7SZ+i5NifFOEwQxs0l52qR90RPlH/YNUv5omGib4H2Xij3Q
KZ7wrmaTGvMpHc8OfzmquCrIqb7Wp3RB7ZsmjUVH4vk+fkD5KUDtiVDaO6brr9yG
AyBwPixdkj76ZsnMmhmvQ8X/kfYyuwLJuWA3Q+FMgqZdyDL8202IZm/AP6/Zl/rg
84B2i3dZvxRFrbWsmXojKzEhErdrzTP0NouKF44Oaz5PnoPZotn+Y/7ti8xfb/m9
o4hwao1N9A2nOo/f8eJpGpeYpcZqu2QyAgx++OyKxWCQfJUtfVsGYkPeoQIX+0ED
Q878RCKF7bBbFeyeJMdLhjocZ4WeeCY3JKB44BozgJ8zlrsIZLmuMfK3YSmUR+8/
UdhmDdyV8w3zPT66lqsYjWYu7m3AVY/jex970BLo63BEcT80KGBDIpwzEZeXvk5E
7Xct6svstQydjx9MUgLNN/20736bAfIDSQqf4jRgKfoHf+VuavJUi+d5zs3OLBLf
pmOX1Swsor5xO8+5iaRHmMuUIvyb/oMeK6Uhpsn188X81IyRReIGDN3RmoXgIm+b
3rQYNJ79vlWOMq8rKJGKOs3JlkuPWK6ASUNZKiLEfdU27lVE7n+JhwSUJ45LaM0F
1a1m2EgMIeAjnCAzsKGv5Njx4z2DUZAZExd4wGxEfZHfXzpdx9R7Bb7Xb4rq7SqZ
atVTx6R8lWe5ec5PymfDx/BV80g6YapZHl0cU5kqCpnohJ0fABsNA+2fg19eWvL9
W2PBgywL58YCWinhZlYf3rqXRXK78Ki37hX4YmX/bjxKdkbi9bPLkA/b7ThdUE2b
Jf05/2/yhdbZg/9B5WByGHkGB69BosR7IryzNNSxkaHBXgtuOlikgwN0rqkHef5G
gN7+SIesrUUGk52Y7uIGZqDfLqz9dK2oEYBxnrndKmGuE5l1j15vFA1tK3FjwIW0
6wJplBJH79xCp09QbE7oUFjaGAMo+tlqTg3MXJPCLK2TvSv/ETBRSToBscdjdQvh
u+hfJfGj8jLOBGnN//vdy4fjjErCGdE5LpikDKXwizEtQ8Ad+8lrmI4OtYiXa1Wx
V2EmPS/QgXASLDXqi2lvR+SIAAc1dDEiWHUqrn3/jkbVlmqIH7EVnY9H/tqaQrpG
ePCreeSzNitmjVdB+ZcugzGVvbgFloAS/7Si+r9+yRH1IZXm3ynaiKzB3vjZdteP
cdBoE1nn8X1Dph4n8pdKiY2iMNXKF7lZw3mAdLjeQ9K/5ujjiTyNPU0FKQCajDPc
9ui6mtk80vcHtCSkyldXszw5XPVFve2bRuuuGtmhLy8Y6sFMBHOu14qNceBo1lb5
CRR4J63MBk7jLNX8FRmJJnuA3AlxcDd0I8Bl44ldHERtiFhVK7taWQ+SLk+xKeVz
OKxQ94LQy3g1/aXzmzQy8HqARGCSjUbU54yNEpluZrM+fQ/LPFlYuBsh+EuROQ8g
WebX1f7BGggod3RBybBwjNOKzkohO/KpSwUHXvTfbOSIgikAyfi3YcGkVXKoNiQe
dpuXbGW3NN9PfxpdFPFgv3EblCOy048JwVILL9k++DbwCeSrn+K/HqXgP9j/Nm6Z
/+eV4odhMHrSrsugn1rFQWK2dGK/0L4yd1So90+vWkFD4N+lHaeXLgtNjX3jYvqr
1fBtt/N+pc5LHPRHvJXCVkfq+H8yRYnlo7tXC4ICjN9rsfluPbl1cpVkNjSgL2Tg
tJOBoZzevfZ+9X6PHdOsm46Po+io5+lm0HdNao8DEiwWfe0EYcvKD9Yt8NzZ/sr4
xIHne97xWir9dRkxdS3b/GSRAa31hvuMo1vhJCgRE5guWfytCFZ258doNm4HQ/vO
Crj6ACCU0hB34+aLmwD5PyGdi33otc0zIl2VovYDyUNdRga57NEdvQ1MMDkHdqys
OKm22pGWISQU9jCqpgUS3MGc0AwKNUa0p7KFeG65X8ac2oKRPnpHsEEH/8zpKWPK
Vc7TokcitExYgOVM/O13/Sl3Q9yVdLzHGSrk7rNl2mc0hpf11NnT82aq+BGqQdqZ
41Gik0uDGrQQvhMrEmrO4knn1TQbos5O2uc7Xae5Zwt7wDE3vl6G4IsmnVYwtulA
hXaPy5TLUQsqNAXsnmXj8aqsq7j3d49p85lwDMGOdMT0BRmtN647fzZGswHX/VaF
Xn0u7S2VfcJUOmk1/FjJQmK2OQGGv8Pm27c1BAGP8RzUQtGR7jweZAkuRkE5dHV2
EJmn/yH13oqH+Ui00w0lkZd8xMfiNMWq6W+/ITjjQwiVHejzbKFPzHKEdbMGr2s7
d3e0MCYYSDApPg7TNhynZzz//Ekfaw2eMOyorrg6oER6EnOOB76le5JPbbrWk7rN
hgP6N4DVHHVtdhiQ9fkOE3uWglSjXWO9GQxEYr1somSp058PLD0Sg11gzyQC/qST
P8rKAwx0mrTMfdLLBq8kQxeLRLeOPD+tmhSof9YTWFxEJYnOr+r3yuGnXIi9NYMu
cjItm1K/PFzp6RhhqH2aS7T5+gkcTKjxyRmMHALzMzjcc0NOTUGmQ7Q1ltHMiacT
hbCxZhYCOQlYiDbtMbFs8llZFuvhkQJmr82DyXyJVAgQLud8douilArhf0rEK6HL
fUH8CiipEmx6UIfwWxvrmUxdOtigXSZ1HdFnEA36E7AqozUb9C2GGwfGbp6MQkFv
MQBk/fcVrVcrt1rAFiFToDFb/2sNC8x99xYIo5eF/B67rqmQwB6PbckK9V8SW8LZ
tVcPPyazEBGwf/q/ANNRW4w3tDlbiy7zp2pIJJe0IZA1cFJv+mAoEkXVGjpMrHQk
OxFmcNdzTI69GfLzMsPHWFbzYZnYKO72PlRwK9c3CkOT09MqorQ9yRhpLWqSi5dE
1J8e2m23wMabKmT2YEu97xfQ81vcZIxdE5200Zba64DByr75A4Jg7nADVdGbLcz7
VDItcpVpEbjGv0NKn8jqVrvOz9ZWbl/e9BE5Cg+ICK549+JDx14PafihnaN9D10I
OMM+gD5Kn9vRMsstfwps2uH05yXQ7me0YKb1nB2F3NlybDzwzkA2KaUH6bJj8BjJ
/+nCwMsntLsvhXjI48WOQ6WGw+Xn7HtcdZaSdm5/WCw+Y24dMlygg69POfFdR8oV
pZ6V1tci8ntQ41yEo9Vt1rj7/+AbqeIq8iwQDCNGmUwx9IC7VeE+11iUftJ5g/be
3BhpmTqOUeHiFxM2BawvqSORCHjcp2dHCpH0T+nyCnCOvC9a1L5ETM8UIf3X8dJG
iK4SYuFe0qXufKlmP2UJwqoRTEQ2akrc7XhYR6Ur6h8Y/tdFuk+54cZvrZR5Ss57
LRnTgmmGDJC6fCvb/rV9XyHuf8FmH/YMLbnO2JmMKPsyAXkB1oVDUMrYXU6DDSwV
3hD2g9OFSCN75g+aVaAzifP7ciCdutMz9AFz/uFjoNglhhiI6ocOVszvV2dYOggL
BZgiv6FnEBmXWfRYZfMI7ujFmlLcnMghZzcqskL9Or2zODWHNstZaIiQZ+mp/GUK
p74/OVdE13N4fcCVrDUfcuBDBrLQlzJsyhMxVckZ3VjFxgRW5FHlcuzF3GeN77Qs
V7ZGhoGLwVyBjev9bIpFSJxMpgoXZP9xDkLUhkvb8cC5+qSUSgkaAzXezusGteFp
ajV2wj6etuYRqf/j7Vh31tcrpsAEPNq11Oq82m4BQ1jzZIlF/Fj/iWPXrjoxuTW7
DOdmR8NLqHTG9Vv/1/QA4F37QEgGPcBf4En1cfR8KkXkywEKUHC5mFVlrRsYDGxr
q/INFfdVr7pPWz2p8+s217Jr1+ENJYYqvwXPjPMhg0Zm+n95DYk2Y5UJ9EOJqUmd
vPq3U9yiceQfsuxK+yZCgIiiem11fodUCh506baY0OMSV9vN8GgyhE7DL9r3iKvR
2+ncxJzAzLixB5m0uSXaI9efXRcQguQtyEo6Js71YAtswyJjfArXuyEt2/u0XPjT
7Ybsc9dYyWTWQyYqlE3QKnKXiEC2pmwutF5+zv9cV8tSRv0ad5Pb4H7NDwT6p0c6
Bp2oBmkyfoAwvLPKsENoA3AGEKVOpioUYGDLJL0GQr3ODfH/V6UHio9V2NflgPWy
6olRMPhiAIpMiDjVKwY6f/Wd+VGWFzNnMBkYV2eetSpU4GHXK4GerQBPrdWxkcLV
NTZarmYQ6KLMLoC8f2ZE/gI+fUQMnOrp/UEtEZhOATWYpksgNsT9EYve0iCwa3R5
ZMrBzbSxiZYi5RrBIESGyE2/E7u17DVFYzGOq6LkofDz5wwYXjcCOy5Kt39sdUYV
DS/USgdHw57ehfBmwqvxUiAmfHI1RDEJYN5G6kXdxeduHgu9lO9Bo42iSHJvphwb
aZGNQ0k3dtriXpEoszVG/n19Ciq0I2uU5OqI5ZSyevCvRWffPtjgLMWpgZDk7Z1x
EyHtyanmhrT/wZmhkUK0rpnu4Bc4dJn2t8O4ELXFRQxlLcggA0YuIn4/yjaqHZST
RZY1ayTrXElDYiCBry/h2/c9W1OUz752aIIgVfgqULNfmTJAhXx21PCt6j2jgzqV
q4zPtGvBNSzlMdpBaTWeWWpr9FysNts1qwcvMI6yB98Y6PAH0V85kwlyPfKqwn0y
ykY0QcDwOSlBpO99yDM/r27BC/8I7Q3Q/MjHh0/2BPd+C33mO315TWIu2/OR/8bi
Ids92W0bMWjZYw08O/zlbIh1Za2X4hQFPz+B1zqKAWnPD3i0zOxbFYRWCP6iNF9B
4MH802haaMt6vrE2fWga7rM+7L0mPDo/Q9Sc22vn7t3fJKIpvt7zEUIRC+LJu11P
zJFhkWdnTm3tQrW4wk/90AsaI7oEA8hIxcaG+DQfriUNl1UsgP3c3e5N4ObovUaP
21Dnx8mugbv/Fn/hXyQ5xHBpdTjFkqZLjHpZRTVkIo/nF+lXE77gfIv46jtv2mnw
+v1KYMzZeOV2cMC1VPcLUfqXwcER7JjLpPk2lkTrP1ztcZGBuif6Yz/lB2kCSKfA
V3kEY7mZbVJ/4nTIPgATzY/9TyfKMieO20mEvHCN4Aejv/9DbGDh7Dh7DR6FfBwN
hPLJAWKb9x74CZqJ5y3Y753hTZFB4RePTj9BxvC4P+OIlyRIi5N17f8U7l47xjRh
Q1tuEPEmhj4X50yyKIc8XUkuEsaQBD0YmjS4Cv3SL7xYZaYUxm5EjXN+Lc+uSUMg
gMPCl2Ej0LqAypLIjLsTIvTCgyqkz3uAah24WqS/iHCqw8ZMViJ2AKS0NR1aQV/0
sUpxZpl+rhKsP8+1mmpAWQMW6qa7pQ3c4+oDDT6AERNW/OtmRsZ2shWOC9Ox+4Xh
TONoLvV/dE21RfxrrpCX+x0ITPUMajU6ntLXXkpp+Jl3DF+NKSM+EIJsCC4CJblE
XsF3cIiIYHMMZXFGAx5kL4Dc7Q/oh/gY2yIkJhkz4UAe7EROWXjjaSNbEPCS+/JL
xhcTo0JUBWKn06032CAcDhh/FEsVj2aWAUZE/TejPdJxDpK5ZzEqWSTpZOB8SUAm
dJlMUG/PayzEt1WUc8ub+o/fHJ6oTNoa7+2tyawwtzETUGMHWN0PQIAw8rK3PXbi
44D8ODr0xVwedparoDkpfG1IhKMYMzQK1u1aeXaZbz/h5xyBL1xJC8yJNceayFqj
E9amkvUp8P4qTxr+49nbqRs92aIyLxmhh7XurCgBMDka493JoQNeTFpVu6m0kFwd
4/vKPCceCeWxw6Ii14lCmUu9NQNVcEKUwEh62o71KiJhYKXN4DmtSIewzalO/g2a
+TCNvbhLefYLsATcCGQhoEk7FJLn+oifh05mOwiAAt4gi1R9gW37CY9KzeD7IquP
6uaf/+Q3ZHvs0w2CKMz05KFQLKt93UwxjIstJLyOdw72IxCxcvzMoHaecLB+afhX
5DhbBaWQIIlWarrhuhJTjcsM/7vOu8aVvJ0a+MRHrgwSlGg9hDHbb3ElVQOCpNRf
IhHs/rAgh8b6QgulNeF5Pqrsxkw0O0LWcddK9Q81jqqYTnIDVOCCF6OA9nv3uibH
TS6c+uPoQT2Mu8ZJpyAJvSDkgrHdkcv04PnBpGLbIn9nn9mnbkShvZc2qsRjNG0J
L9IkS7+OppdsVOuilBY4NXTYAsaTBAi6vsZfpowNd/IGIh3NxHEGtUaPiQgVQS6V
uMAzHAKk7wTyT1zyjhVoKpD6Xfe8SYWUsS56d5yoFCN4oleQc3SKA210qrYuoU1I
/mVFLqKpKbAbpDkilKgoDncSQ6HNydv2aTxsiQpI3+gPQKs6P2wlDWUTjKOHwIGS
k3ZmEH5e5tnW6OZxo85IS7twGTMLfZ3pYne7Y/0uCjOoXJVuhj+TRyRuGJELp0KZ
+MTfBQyu+FDJ6K5vzC0RWq5SJjrfdsO+guOyhfwkZoX+gkKGwRsJzqIl6kb3v2ln
S+6QWuCtvyfuvurem/VD2Y+GMapQB9RYtKF4nHKQ1hntKL6xx349Awu455NyBaNP
TaGj1271mF8UL7CVZAxi6scaqrVOFEzik1B2+ZTLOcbT2hMdv9edMA7ar7OkMFnZ
ERToih0NWZxY6Hn4cB5ngvCGYbe8sSEJJxYlkYoiP/sN/LzlcDiQtnVLsFaT2I6R
+28nE0Myxd5elQqFwjeICA9V5nyYP7NOaC5g6mcV7g8Dau9FVl/FUZ5UPJWHNTTe
fNFdfwDH/zG44W60gQqVS0Pu3ftT2e6U/4W8RXgw9iInh7tlpjQvAYDbANc+qE9R
RuHyhm8eQi3jZbbJWOKQjboYJizlyflSJfFCn3bU6rdbuUYNqMXxNmKKPPhElde7
TVyMXB+wmjcPggwQo+M40zgeZ8CT1525H/XMxxJERvwftSdLgqM7B8RrIrZmLf7S
Oli/Hm3akYolQa6Omp4LqryeACSHgEIkIkYrSNC5FQegvo/O3AzG4a6AABxDpW5b
0RX1mqALqyJK+NLuWYkbZbMLRLhxAQpdnTJqXJglqo4Z3nd2/oJpt4hI19VQF00K
ZU+XuKLIRUa4+3VksU3HO/aw3iZpAmgvUnB/LeN21Ytr4advaPIeAJayEo/wNB2G
phBtYrch7nw7ouBpPTHWUqzcS/OTSBFQ8GpXSMLx1OB3Xa34OJDoFgVa2dc6dstu
sT6gvutuvOKG33d0yTeu9fSKgi0uRFmsokGFLe1aLvpBuoP1UnlAQuxxYaV2kXjA
KJL8XVw9QZTX9L3bHPwgbqttR9xRWSq2l5V0XkepuDDSq9Oz3F1Pl47zk5xsqgkB
QvF3+4K2QwElxIU05Wz6C/3E7ZhSax1bH5uChcoC42g63/kFXQEK6+HhnTHekU8q
GMmSsPSdDrrC0YGQZB1HhXNs2iyaeSCquj+CzlZvU79Lugca+EvBa5AW7/mLKV8a
bpteY2awQyERqcDCkybgTvpXPuvm3jxKlqkD4VChAuivoys81CXPKtUm03m0d8Ev
lflCTDyZ9nytFS0tQ9falCZ83izqEXzeh973a2R/OQh82E7KsADscplymxAaXz7q
1Wvfwa2K/a14nq6BpvG5SawCTab1Nv/DVw4FbEghXBsz7ZosYE9fKCKXnjOGdGHn
PI4QjEx0iG35/HmFnlNHwLmJVbxqGNA0uUTgMLZE0aTVVFqvtSoN3yv33cMNEwrf
ePuo3Q+8tSh1LtHN60p+36PH5c5n28V6ghj/z1OsHeNBi/Y9jK+BxwB5WNCv2bTA
tH8a1eFtG3ExX4/QPcswqTHYbuOgW4yunAfupaxfjmuMoNJ/z8lNkNAn0MQSaMjj
xjtwDgFc2IOW76a4Ddoiobz3RNNkEiDdVY7BUrVj8UZ1CthJWULmJz0JylyWB0pW
+E190QvoyhwHGo7zK/kEBku8DXSUnt+zYPIwKIGeTY1Y2HRGUCPiyXLInbUM9p8w
A39ZB6D3QtbSXADE9j3wnvNxltOi07bN07DmtWeh4FEdaoDJU6kUMLMUUtxPQM01
+n7LCHyALUvObTo8u83KaLjzg4uPd6JH1R2aQfzSoUFSSozqPmP3SpoRxDBepexj
4MiuQwvuN7uNcYOS2rBCdX4ht8l6K95nchMd5KM54atdEH8FZzIHsvTnUfzWY+ml
joqLoiwIpZHEt9DjZaOWFmkzMOnt3PXyZP81auZjCDyk3TDwD4pvcTUsMYc/Mf9i
Zjf8Qa9Jv1w/EUa03NEYFuGoOMRG7qJW+xR4MnQQKSpsimJ5xDQJ7KxtqO7swWDm
w0ppP+i4GyuNuC1FR2mKiymLcSkJPlUkRon6+B/cCXOAmg0zQZ7XiPOPiTq32pAl
6qyvxj+7tTj1vkDfmXipVX1OQGVHcJWJ92dUylFmlVZfN1PXRGR0z573VsTGatYI
UyxS3O/hlLURIPsO0wLvTZGxeW3WRbAKPa65W42Q1xPaknKtbYu1kf90DIUFNlT/
Oz135rEKthkXqr5lZdeIgSxBlrhV9VxHVSASxpuk7lE7+nZF8siXQhNlw2Y7N4SZ
P0dZR5IC0QRArcMST8Fk9RxwitM0Hr5v2QsXO1x3/NYUS3fT0WUAcHolJA16j7JE
VtycajyeNBLAnVGsrOaYqtzv+gFxiCQGrzHZKUMdwZkYB1hUXMbABqq8XlYeA++e
ISBraE2Y+9WhEuNKl7GNdlr9uqkxjpLjWeJRWA+kWWnYHt361JnSj0HzJm23cvVc
tMFSMwxlIdlql7fWQWBrBQVgeVeZYPfCKs12x8X4AwNf/wNyr05/UwttCHBrej6I
5ImV7kkZWBBQeUyU6rzt5U3HFoanCGOf+Lc9wwKCd0ju+ng2wKgzJbMf4NIf+r6v
AUFQgEbg90fNNk4UW4fDBNJIVR4HNsd063m4pMGReR0WaE40OWjFmBuiZTQQU73E
f8VfqYswbmuYykV3QJNgnXUNjgCG4vSJf5JRjcIcWz8/uWDPbmnZf0mAZrxE9jbe
sCDOb0ejch3KTAheMrp0ldZXPIASFcb4wpaQU8OQ1O+X5TycUvch4ghGivFx8NL2
J3hmIjxT7GxaJTNkx2aAAiKuRNt4jGTDUlKU/DVRdOUgOCd+a7HNG8PeIMN+2QcD
Q+/Sex9BpOUsWTt4oaDqatbuToQhYOIc8fKDmaoXi6MVyEsLfRiGvOQjvtsAkVT1
MBXeKL/G6WiHaZxMhjOmd3wUFRiZB7Z2O6G9yOE0AogOnCaUUaz3Cmad6lLWhkj8
eK5123iyk84Dqdv18RQGEJs7q5shyOssZBl58KFudzJNvqpv2f2XD8kfAeHO4zn3
7/u38yFq25fv35vddSzpQvIitoAgdEZxjjmorynMAqn0eTq6mYMb9JewEX45KXrO
lP8tFXB3rLMjpxbhqKyngZuOXahfM4vx0LJFd4M43X4xlKu8E23XGUATvthgnZIP
QN5L7fRPqAoy8bIStuRwM1fwEpYQY2nOAxgHl/XWiRHAoQEb6eDf1m/BzO16o4Jl
u6OkAnEqb4cHcnYT40hHkZ2vY5uGkmrTvx6LXq378LEYzkhKEBTXofCCa0t1Qgnp
Or1pDjZN4lH2Oaj2O2hOVN+bfb/RwRMh+n6jdRKY93vmRwhCGVn9EgUj6J5mCfXO
bonQtT81xA8rcyMGHv6McgyPYMoYZwCJwToOLc6pMBvEYUn3B2HVC32e8Z59df1b
kYemoz3YMtq16fPkVxCcFKovG+pTvFe0fE2C9NukZ4ARc5RXiNruptL9ll85BF0Y
0V37WxI5tR88jtbe6GPtRJzMX1huyIBOXNU55wFcrp2WoPIlnR/4bHJRJvXTu1BF
WGiNlJ3lSOi+vPLgzBzcKrqfyL1fFaNvCo8/E5EXfs5AzqzO0p1Z1gj7nglQtiGu
azEaNE4ApCVV8Z8kTH8cQgCO2R41fv8/97ElKMKlFimsEa3D3Ua7t1VFZ1nGE914
2gZM1CO2h3Ahbryq07ooWI9wq5uMxZwwTfSkSH+rmpBqzICQHPQotrjxclKp+2uY
iM1dZwMsgDgZGhE37wZLWo9DjLzgbLIS2AFWvvRpyS/UNj9aeOOWBkDsQgJyWr7F
jFm5OPxkn2n+19JU5ZHsLGgBflb7MLmr2D3Y7w47CCeyjXr7kUN+uiv061C48ctX
nXY22kA9EK0veWy3VVJht8WZ6EhwOAP24uYi/gXDdKgGPbHGm4jHUCzewoK2fCat
EVOQIDFKEbzswEs8mp8rgtEMdP0W3/WCPGrNtdQBIrLrmhBnlpBStOU1dzdgy+fC
KpINdnsZG3ttRxKof6SskRVhaTqTRwpbSEcFzRBA8xXM6FPjfP0q+zGtVHB3yFbT
R4ZljKwy2tB4QpVSBDJS+p9bWi9m+AgQsSfYQNUl1HcNQUrMQ4h+MCj9GPE/ngVM
UOLoTL7q+tlpQ6NPBe3AKInbha7iR0plt+9buwhqkJuBTN0XDgWH6cWBfQ8up5N4
lhbU83NGmMWiED0vok+SLEBAsNednL8OjfrX8GqCtvXkgd/K1D8lWbqH3dudPmmv
I2Zl2C5ViuHUxTAUufHWLRpmHJhIdjviGFTZpYch/GLcFNmLle/Bj2AYYv8Bi/Py
+lLI7mCuiSaELswUe7RDh688vcsenoZFclll2v8vKtFclm42i+IjXhMWphRieXL7
Zb/GhIJs5elqpo6MjtQBD+UKXvU1aZ4txexR8akT3B0bUxR+oQJDJ5eLCs4UaU2M
avXDT9jG4TQnlAHLCkQ/Bi/ScSu9LtsB+FBLSsx4HegZMIzabMNmrsqe8E6h5qUz
9c4JyM8s16KzmE4/ZOf7EkIw1xwD8ADOxmOr/EntUEMXGGed4Z8r+Spy2upIFrL5
R8Las5ufOO7B3Z4UuaDIEgX8/DKs36x0f6fWNuvkUsyrdskNwcL5N1IVtWimPZz+
rsyGwzY6/wrgtwINLzkTCMAKGWwFccCNm3LAjidF/GtW+e4WGuUjMGJoX7CIOetq
3iv+I4RKsvIermPLbU9uC0uCPRaf+o7AxMRB9Jtle9IO2UnGuLz1/cFzbnBhROH6
J+2vQWvO/63TUm7MfhwEjKW87P1W6JQCHHFzb03ckpDhL/ttWyo1hM/yZvpj8OOr
i+zxznFOihwpjzEv7YfGV4GSmrvFHSFxDIupfZeS5XSRXJNcefzdJF0LYeZ7+wQA
EK+F7zajV69MjcxbcCeQM4M5UkJyfipcAxz/rabb9584rAQVeUcxQxqAqtvaaHq8
LG2teOpKy93A+qgJad70TV6N/PjUtBL1Z1LTmIBiv4Dd5qE1T9c2Hf/N/okxw3Gr
7sNUtnJuxhlPQkWTBQVrryQ6jWKmwGts+ajuSF3rASy5iHL776gbvJS+R51BXLWD
uN8FqXshJeckaVsdURQox3NZpgn9+jqx58engcX7yGtvkWvwvR+k5i3gPf+Sldxh
XSotosV7gAwH8UVg7qvixTUNPpQMsAm6ymbYg4nBVbOWQtX6p3kzsQzWXOk3ocdU
C5BbvP3VZnKmuJeKCeyMkKCBbfpfq9dBP5G7SythHz5fLvHOcnKrNaUkNSKXvHo8
9y/MJSkYyUvq7rONQpgBPTZ52bNfHIl5vdNnU4FCPmQS2ssckIIbjYOtd95c8VUy
ysZdNv+MPa0AhgeCqOenZYDRDJySVOD5uH3xO+gkL3tkB5yqHMTyDiL8uIoydMb5
Iogs9EgQePNUVF0qseZcnbsaPs01BEHxP9aVbDXhbtxCSEJIRU30SiA5ctDmFg9W
Z7kqBo6n7p6xaIPb4KY8tgq07BylhZNwwxzPZrwa7kYtob5y6rwCSb+HVspIQp0k
uMBtRcXfSe6aDl2mWtAku+xz/66HwD1gFUlET5Jd7OmI3AnsswWhDMmNsQyd03TB
bAt5w9N3ydy7iZ04/oZt9+o7a23WXl552UgjTYYJJvuTCt9o0Vx4PU544E85e2Vb
8c+IUXH5WeYv5Ww/dRWTYKDCMgkjqU8MHfUJGIx1vKd/dX0ADs3A0cnEGVPZglsa
OxE1/VTKDNrO3VJw6d9RrApXunxlPrdaG1UINYN8CskNIBi0WD9YIvQj5CvsGZhQ
rYywCv+CcxN4L+Kai61kkfW1K/Pf3Y4eGxk3IHseSnz5oR3JCTCT+tgqW6TYvBj3
PIzPOTq7HCPYNhVShHY8/VhjjxiGjXvbHQ+9GH8YZQvqsk/2Wecc4twB0wE8Zdqs
dFSV6GfBWO2LbloVu3TUuyfeQbSsg3GM2/odct6fnQhfIikt/q+poUJ95ACjbM58
aC/t1A9aX0yz20WQOTznYyrImCkui05hfDcWlvU8PfKK1UKBHZYRHAdRrIkV0lvb
X+p9YxeUSVUMqW9EIeYPCaua5fG5naGiOLnkDtR0Qt2A8vHr5o4W5jmDE0+ph6pd
PKJv1UPYSps7Sy7uHrYfoaxyV6kd9Zhvn+JQOcx7iWUyDIE9C2LbTn4JWghiDOaM
ZyH7TtMDcAByX4SyxY1fgRKMI8YlgViejNpaAKg3PBp4s9MJo+yKZyr5h50uvhG5
AhKJuexreMWcmdTd57ZeAMKA1SidI5AlsZPIiRjwocpbO/rIyZMatPmOrP+ZuToT
HxDh73b281qKkkwQa07wt3NlCu1Id7f1Tb2XcmDN+j0sgacnZJhSJkerhZ/1rth2
lxe6m4NH1kAYOBRF0ObZjz/G6hcp+7t+L/6wtbUoJ7u/xz3lHqsuIWOn/oYQKMlI
QuaSHBWGz+UOJTznSCq7q/xtdokFybfu8euIaiX5x4CHXD8YZ/U/Y8A02jjN4NBq
3ok4WTyP2oD+PtEaULU3U9Hgcd6udfVwIi+L06racoqFurzfnRcuYmyd70FEgbPu
kQdnkdX59Z8HYDTo+2HlTKPFHue9ZbpPSiyNQZ58VL2Zf9svEVQ955EzveeFDq3s
Y3WqjOgnnv9t+ovP330bJ/8jlPvmw3voll/cpSy9SVhSeSu823g5WOqVi8KacdB4
5KWvKX0KjhlbN6FbkzWa/oVNayrBMgBxh2m6B6f3Bsbxs7RFA7WNAIaDYSlQPha6
hSwVdLAXvdQHVdId1sfBvoRRw1Wg4iZamgusENZwFyBakKJT+Vx4vaxNJBb9oQVt
L1LYOzR2Br1Mye3Vs4DP2G5fFfMo1cWWksRUETzIDWhf63FpWjgtP/fIzuNWxFxQ
1FL5l3B1Bcllc7O5u4rRpNrsvXerVEPfz+fVgMto9aXVwd0kq8xIfPu1PUNcjsR+
iAnXpVoYEwa/FmUPpuQcOFMSTNcOU337k7DNj+P0Hf00jDBgBMwvji7gtXbh2sFq
HbUO+zeYRxYEGEj7F0UQ/8cGisjEh8zXHaKVAoau6W42SGws+t+pHzhL5iKN3ZZ8
mGmBbAOaS/YUPNE5usAdLiAPqU43MlabiCyqQiQ9XNwuQZ62XeWKZZtvIHf5O+Vh
h1yFvflpYOyeSfuhaV2r/Zow4WiJuXsJSrTuONT9y1h78ZintDgZBtM5IedwjG+U
QctH5a/PyhL0aQ6NYtkEM8ol6GrJ1qgROf/5f8Vc1Y2pA2L65dHPSEF39xFJKeuH
4qEHnDE4OSE/XANaGRke6O58xpQhyiU7NYVBODJIbkMUfKakeniu+h7fE9bTdi5Y
9YYmedkDw9EQcQLe1r95IGF2G2ZQdafdh0C1s74CJPZaAHNTFDc5lnPsEs3MBGSy
/iuYi99TLa+KmzDLWejUdD2MeybXKgvJptmgDl2lBySGxsEKbhzHWXnxf9Z9J0W2
nNy8Z6RbnWP+20koVxGjjBq0f8LIpfEmHUvDng9N3+gbBrY5BIPu2HJy4GT7A2mI
zTR6bE1eyVjNmpE35EiJfJZghyoY2q6NmRAEq8o6+YSarii5ohF/OFfrZePtUGMk
gY7UHTrCY9Jh5YAIkCOhScrbvqf6LWQWUVfvucX1sIvEDfyHHstaakrdIucfDYme
r4Hh5GC7CCkDyKnnJTJUUQ4rstSMl3/Zi1kpqD9Z9+nWWm1rTb///ymW7Ca+0r6F
YFeH6cQlEHoWG19Oh6lQEeFR8edaIxpxb3ihxp0H8PSBpd1mYzgsNFH+XmxSLccf
PGzQftocN3cYWP3IHuwTmEkvSRB1L0H4LELq6IbXDlY5iKdC/UFfzYIwHAiG3KwC
mG5i7oS9vh/5A8plAFYFz0dNi44iyeuYh0M5hZ8u5XvsoB7HhWlbevE/z1+EN5t0
S4G6GgtbmwGYu8rz5hg2u2BL3BSc574w+kp9RwoWlf59jzt3iGo5WNXACJ3bljp7
8Y7rQqg7z+t8iC+YtE52VqCvw98G2o9DLr2f+Y7vCbaDBXW8bYaZc+DdFpdKhi+d
LutualrCMFSVBKDGrwNiYu/qe9ykELZUwUYDLmj0Iegm0ighIepvNLoDwYH89qQP
T7oUL4lKVuIkjWv81hUssZGFbtE2K4QHJ7/lVYy4Zrt4KBzOV1360Um0mC8K0TgW
tltNmYmOP6PKUNvXYqcD3IIecpwFevbSpKRi+1UhV6SXKkDdo4iNYn1rZnDY87TA
t/SHi4oF1OWXRtCUDuC2zYK0E58GOhrs7y8INERiSjZ7BcF1lNiXWm++7F8N95PL
Ah2yuenJpKYQL0v3pNXyXcJBVuuvAROWzLlM343z6Uh684U5oeGmJTzhp4c2O0Bb
P97k/FGf6EzRx5mzmRhGH/dtGr+Sbh0KnylfCf7+O+GXz3JXutZALqkYefZjIOhl
nqx34p7gYArKN94WWAvr3a65RmEEpwSuwS8BxrdjEpSxzKNvVx0bDSiqtv6V6Yxv
lfMufntC5sa3wIFGRqjOHdXw90HUlXuBmPAkWje6s3HoAOh8n8jHEkyUas9PKD4Y
aykA2X1+v4/CAHTpVqX3QdX/DgW7jAiAtSuFxqqV3krr83VEPL9gFISND4LoGMtm
xBnrE7nXs8Iv8RqptRRZ/dFfUrO86bvuDSp3wm3fRCqmOno5Wtv8D1y4ol9/2Kmw
jYA+wz7acofvnHe8VRcHHEVxDcRAa9CFYcSytCLBrMEay8YdPqSBhtyJiFUDYi8M
2s4FUdraUk/BYU7dJ1rrQoZgR7OlhFVxbL/9Bc2U719Grw6WZc0wh9bDGne0iumI
Wi0IR8uKXaLhgGqwptIJLcF3TU9Qwgry5SdYI7BgW+agrkZwF69SxW5ChxN4G3dI
MUbunGEbQM9WkQuh/7ghDfCtWRvsNJFdJjsa/nD4WGqBHPiYo21I/5R/hrJPbqjc
P+/wFnLa7lA3AHom2BCZ/x6i4f+8VKkwHlubrgPC0JpbZg8CerNbVGbi++XNJ3jA
B8pBUBJcwKWTHUbNNXgilCnVTMhip3KKrPCZUYP2ms/IAmAJzCaG19DxSiti0EiA
HUyIAL3Bx/eacH7BPcsjQqFchJChqcGLSpJ3iPgqD2JcCk1+qFcWJXy9Gt8L3diL
ylAhrg9AqduE2D5kCDyeJQr7PQtheB83Qt0PEpbo2yjP+q+vOGBbrq7rRKyaRaNv
+i6A/iCISdbxc4SNrcPIi1SBSIuXihTEvrojncHL/byILGwXaGyTdFXcF9SgiQCo
FKeTLCxb6W4OnaQ5Im9nf/EylvEifRcGNi1WCTJgAEQCd1XTorUJB2j2dIkrErMP
1BX7zOC3rE7r3mLg3D+oOjjmhPJUfbBy0iA0Dk/vZ6q4YGGJ1gwjfTE8PTpNGyot
sUxu/25sMw9XZ+eWjdWE5SbxLDIYX0MlUoNPPRfFGvaJv3ogOiKtJOgzaMnd23Wx
gW9nlqPZvcMJ18GamGlft+QS4Ks6+Wb6eHKVfRgNo/2MiUGm4Yg2Uci7wCm+eUiv
WFZBQ5c01nUlf3mHWCu/TRcSySB8c+hBahU6EQvhlr/rTo0Nfzz9cPQJ9eJsfE+U
p5kP6uiysYRfzvVk8zxjZ4fWFvixTd+4YcjXeVkdu3kZRix04VTJVs7+jRj/xIij
Y8/9krmRQdIbO8azIw12agTsHCXDBWjWWO1FSUAAb515UgrfAqI7MH9PeRKs1jfd
RsujGW+x+I/Fz+FSQChBb59h0LFTlRMV7eQCVLtNw+b4FImRQ0FJhw/0/O+6N1A3
nM0eCkkBEVUSJD15Sq+y27S3/AQ/rBK7M03FZn/TgHaPfJQLAhnHBB8TvHaTHE9R
7QUPR/4FWKTY3PYAfWGCCju3Rp4AG+9u1upozgobJ371QA/8IOovS85S9ZGaC2ia
704+iHpcOKsLOmK61OvhCWe7VFdkSRDOpz58BF/u2zeyLfaclC6loPjgjZJuD6zP
FRfIhqueg+6cIRdA6l2i2FKHXe6NOpbDmU712ktcYfx3nSMxj5iKN+zOgKQFCoY8
UMhiA8FS1z8wJOqTjDupbSWBlMry/fEwo2NkEJcCMasQRT1jg4Ydq6fJVEdU7d+4
PqQUV+pITu5tPKh0qsEe4gCcMEDWih3ctLQh67QlHpC27jrdWaEPv60bQRfvciY0
LvLQG7l5SlvnFdQtPQtRNCZqNBSLX87jtp0+GtJhWUBZGd1PXjdsjyUZwDQRYEbq
fhLsbdITVJUskiqdq2qtAlWgvxYaZSNZ22EOiB1w7GJKavpDiUSuoB7r4u2lRfCw
sxLJbyh9D7hJ66Bo7cbP2ypgMYvpo+7sbWbPtpgFi39tg1M3GqPAzO0uOzs3xt0C
VnHo4g4K9cQ6GdY39txsC8eH7ANNShHu/e2v0uz2mVv1RYU0iMcyMY/M2je3i/FK
MVC+OVsiqeNeqQgM7GTgzaXEcGuuYx9PH9/z+gxEwpxUBsEqmcS8xSI7a393WNHe
Wu9Xz6aJfvzxEzRjOmspKNMF+PVu5clwwNBgen4vZKE8EO8RmzLd89YlWb39dXuS
f5ZInen3fv9uMjEl+2SzL3GZihJtKjY0xaYgfiWBN2JxikTGOMJmmokyLWfx9TXl
hUNirScGbTN78bRl8co/4BQWYfXX+PAs4IG5BG9RH65+VVaD+DJ5iGaEbv6z7xd0
CPjrTr439dDcDe20T9aIzGP6H9gCwQBwZ2Hj1Hpyuan9NImBXUYCTI5F6GCCs0MR
s4CUfwGYlsu4eYpRaiR5NROJjMU51VefR90lOWo3IT4K2n8qb73d0J/0CcXzAsiw
O9GTkZFDFmSwD8ev2dBj62t2DDTZQ4azIZzSzaDXWJHGK0XAA7TwaFmZ4+GFNWBT
ZwaeHVHexZg1pmVDYdGbNctdPMh/OxLG/fhKJtPKSrgP62+CQlGuus8fzlFX0gKA
+IVaTWK9DI0YLN3Ecui3l7MnbmIlSuaAgwvhj9zcjVb3GkSxrURnAbpVW1nLatK0
QGwTkLNPRK4bJKnjvVn8k9ensz2z6PoIVyZFxBuPIZWwRMyUvudaD+v9eKWKPj2G
b3XM6JD5PshqF1mcsEL5Zm6Qt5Ffkz3qs/k/JLD+eRIJCc+BKYD+DgNbMK93sUl0
ox+6Uqq15QBvnALEVk4X9xUnzmNHa33oAy8wgpLDAGi+qrtBuFTnK227tj8CDYPe
GZklIdH3MfyXui1w1yph49BAddniLkPKMYgM3Nf5AXqpgE+khz1Qgie1nTkdYbAD
OjMXizPdMOJB1RJAt2wWbzReCCKcDG3mLQHLarnuEtOMjGxExQbNNBcd0wce+c6k
GsDKtu092aO6yZQpW7wWIjp1HGvLwSXjkHBwoZYrrfKew9LafMZuiciO5qK5yxHF
LBmHXI59D7JDfZDPBUNOptjc4zYiVplSozKHRvtdV7C6LMU+ZQLBHR6GuysRwJiw
boBd6EjoALfoDP24uOgZsAlIzE4jvxaCcqL6iE2gCjQmAp0FAxKTV1nRoNn2Mc88
kaREfGDI3mm/VX5o+j8QVvmvoRGRKZO8OVQsJ+469Gqg6Q1xEcbP9FJwc+3STezI
Tihtny7SS0xkc49A5dkqp7Rsg3y2DRpc/ortaYTXJnhIT5j57zWvWybFQPy8Ne5h
Uk/Kt1gHT+w22iL5weOfeWtJVxTGPJFnehioYPpvc7MiqCrBwnUulLLk70ed9mrM
G9cVgYYnhcnELGynhuEnYSDLG+32pN4XUGt2RAbppsWhLr43gaURp1F5N876+cwW
leI975OTllEEmPrvOKJcxZdmlRp0Js2d05DqKqvYpw44N1R0bAH6NF+61VP607Ju
MNsif4KiRyVdxirtIddxWlLS54+ydATRdR64iT2iCzonlvJyVFeeCR8O/IuboFTo
OKx2Lscq1O2fIAFbUFFxIHpsyOHolEqmVDSPja0QnCTqy5lgTl0kSNnZFqkS8BBZ
WTuex9jv1Yvc6l1kfsviEs6SmOv4iXg2ODTDCfw+DA3Xmidkj16+pbEPWqU9uYJ6
K4VnhpxJLy4PAmaW8mHQ4FqsRympqj0cruwhrwVFT9nZ51t6s/W/w2r5+VXP/W/r
fo86X9nKbIRGq1LSm9uL/uYLXAFu8EPPIpTU7xtPXNjDhwqH3MK0w7rFOWq26yZM
w2IdWXrrhYU/PTsnNNikRIWdT06sn8Y1gAsx39bVtjlIy2qABxQaknluP5KHm9FB
trUJk0RdFnqxfJqb2Jm3rKsWY5AM7A37l/GuLUx69LQXmn+fPtPirkbJ/6VdifzI
lgLV9v610nNyxMAflD+F+MDrvB//cSgkrHHncLieBJUkCJR9u4Y8KUY/4RhW29I9
J7EdXcWb0U2Ck/uLppjHWEoRhe+59T9YA+gM+HAPMuNqdiaLCIIag2okLw41OdA1
eOshX2J3EdkHHeS95sFPRqEA2SDiF3TWBpREX6O4upLBwS35nOOa32ShtWVoEYAN
GF1VxlXQCodWcWr1U2NHDhQzGjD+KFFhyAAoxtIF8lrBBVqWyNuP1i+P9+uaCLNT
wlYLdEJ7jL0Ex4Y+tZqYUG4xoeyyF9vta1Mq7yU1WnGz18cPWnd39rz7+sb9QqgB
nEBDwsJHo00+TVXQJxuqUa3g2jqFLS8Ce9NJ9OHVL1KfmD2PhygcCr4uvsOp1XSU
Y6Uj+ZWMUgVqyUC0uaGaSWhYurxkW+a8R9IJzfuYdTHfix7uFXxMPD4PrrEuW2hl
UGunHsOl88anJyj/LX20kURaZN3uRCXa9ejv9EmDn6+t+AOvPVMxXidSgX9af0TB
bu8xD6+daLNjvU5lM1EpPufQU3bk9oif5CtHXM+aakXfDnkYexeTQhrs/HmlF7/W
znRoyJqkgpV3DCIAyDJV5fhRTrlFqrVwwpJzqHOGWTCOJSEueBRk8tRBToR+V8hp
SVWaWQrBuaF41fUHWnvT9XzPz/CdmvvuOEGwTQuIQABBwuBtjXphU9jCtvF9Os0c
L3v0n3REm0yrKglDLYDTqFSYRMEuSHvSJaLnZRo/pv34jN1XbzSCzPC/5/EnVTlB
HG2zFEL4oSGG4AefhxmB84jMX5PNIL4Ki1s7NBGIrSVD8Vn3jdBmj47z8Ii9HYHu
e0Zpc2tQ3moDjt+wwq8QbUdoLS10S4z4OYdPOz+uwKWEaHqKEWUdf1FggtGftx0v
Arry8qdQroNMju+8WJ1TWzbyB4fasVg0pKLaumZ3jWP5wWeZl0Pz/QAHTIfesdK9
uS7riTTWq+yKPhno3ZAeLna+WAvzV9sye3CyrDMmCZzMheoy3ZltOZAd5DVu30ZX
9OL0e+8VxMF9gYdPCfHoni3anKfiTwd6WA/CLH8gMvddo1a6rKi7ExMDlZIaJdW8
EECowAF5JFTgl3RDkiXuWdWY0/01XxkRDRpTs3aEcDlfT7rIA1eN1na0tXdzl8LW
ymEPzEQbgUFiWyX5j+dvN3plETIO5ZDMUo9CxMGOBQ63sceV5XdavUGzHx+QoP8X
ej5o9eHtaq0OKnsJARecgHDuLKFOmJCOJBFhqSA1w392HkTlw6mIJ1IAIeqjVEdX
4A6FM3w2wbCDzLOjWBB2EWP8j6vkJuOHMEckQzVjiqwUl3Bgva+dDva9AdLJZZTh
2V3PrUtYqx/1SR7m/I1Bx3L/36yJPprGsHqrgRdRspTvD/1J63o2U7WhOWOgbRMb
6tCKrH53xbIfzcTE31IQ8J/e9olYsHb67rLv5ChrV41zwm/vKVZS8w1C3CRrM8lJ
qEmoWZ1eeUUty5oskWJmpvgknGDyHEkw3K4w4lA+Lp20ij0+LcZnVtUtvMUtuNhy
iN6UWNzAi19vADDjPvoxFNYx1eNqH6jzYBnYnfYc19mENOYkFCDL9frOzfRR9xOl
kCeCwap5eOn1yrGcS3rcCizJHcyepVGCqqP9rJOp+Jel7f6+1JetgPfZqZ5WW1zw
X37zNlgWeubBdWK1sY6QYlHIuhYDl2lxixxJaNBh3IK7tbognhyMX1g1iPkni2Kx
TiZL0rcYXXG91vTuvvwu6AwFOubK2lfdYECInZK1T5ZN4WJdgfYlq4MtJWREsbJh
gtJturYNkmjlZXNd7UGpFypK26DzzLs7SzaXObCRvGrtrd+DmxiUP0V5TqHyP0HY
BhRbp2aam4GdEP0ttk3f5l95P1MpMB3vZCVTaNh9OkJlgyxH0tSA28upJMnUGyns
4aGuvbKd/VUn3A6C/gzmBmz18Vb3V6Lbndeu4WLQJWcAiis+dLFpcX/fveKMV1wW
vJUIaooB8LhXc4jTho1gUJ0D+Zu4HURsJ+isks96HajTtyFEC0F/ozQ86yH6r6pA
XBBuBz4req98+zke/3EoGr1/mQ4+3W62DT2hjIYc6dGn7CSPWulr9mbxqLWsO/D2
K4NLZ6GuvRh03vRRpmL/ltJn1+5nRooILdDsfr/+RozNoVAm8omhCt7gUUx2wE8f
PrTdQEYB34BqjhiIt1HVOiW5bB3xHUdxLnBUg8JXMfa33HTKEod7ymy+EnsMb6iz
K6W7Ke78ZIJMIzr7wBNG/qBu4Yc6B8cjl0FEup+cDyvBiuXC1skBPiRiT/jx2tBd
OLeLP6bRCSoYJX8abCWI1SjhF8WkM4c6hjjuAmey/SlCNjVl16CMlgUfFWsNiCij
NEB+AZ4gXqxVKfn2qua1K71WXWxEhhNNlMEs6oUgovwSTDZwikXmA/qOnUal6Er+
KupSDaICehr1YGIYAORdCDvOHaidA+H4ZDdz+CcPcZ1U4r3/Uu1hSo+Ur3JAKZXE
zMEHbfOBVoMXuNlX9u5i+KDZOPcF33/WPy1r/lMHvWD2TtAtGmrJxYjfctaRCoBR
R7SUjlTxmJcRmwBFvciLY8Vo29T324j7jbQT+TfGNWLs4mpzPvp3fscgQpP1D0yx
P0k0IhfxbLoSFoTgdEAoWw14f+fO4AyFjr4j1ACrc7rJHgcVXPTNI1pHQNHEhNRg
0NRGLOoBOwFsha6TtPuBpwN/9hhTkVq7od04ZLdJ2inZ6P2Yq2fz5jlCK5UIvnDS
ephzg9yfLOpIy2qFgkK103j6pPW9sreeeWGlqtmmyf2t5tfQIhhFc0687VrtTO3L
V9i9+bcDLFqp6ycYLzuvPZQJ3R0UJg2BiMrBb+Y+WMzk9/FPo5pRR6GHQKabR005
jeZNZcHvr+V+yjRmGuRLlFYx7TnytE6s6GY7JrSJaWElpBuy0ck2gx/ocA9+7bCa
vl+5GLvLdSU0rRtSz1oiUAj5IfFUgrrLxe6HQPYcy7ymOmj7dUACUTMmg81qUgS4
11rKIsslUwdev8SVWwmNS4SezrfZmeBzbDJIbzxYAyGMPcca/9vw79efar2321Wf
lr96sFtgHvUDhM4YDJaE+luC7webKxwnFX65cPINn5wPpYE77zbAFlXRahADor1l
J+8Aych423LSQdHP54BuU8Zs+JfwD4+hvkrrKdfROgF9wuq3Vk93Sn2gALSmZVXb
PJDbwhu3lQRl03SsBym3XgfzKTfrV+RJ0HpYF1Veig+pWiXjQoMgM/l6+SaLXlZt
jkSNJ3Il7FNV1jfWT195Yszcs6f98bd2yUbQhKqo4csYP26SEUzoSqpSr8U+7OZ/
HjAVINqFQk4avDbOJBogrnv5ASbdOLBvvXCREfUNNFygSQRZgc5wnYsjA+a4xmCo
APnpwMwlpAOUiJsdmQcsf0GKJHQf0/Z4ojYD0BUevWeWD0wbjCS2xnC3aK0xxJmw
Ag9yIPvbgFJJj+sRK/aOhQ2baJLM9cRpbG+vXB4uEw3YYca1nXDBsCG/ibyM0rLW
DMTUABptJAtBw8FxLcgQmqxyW3hBVT7RLlULPAye9adf/dGV4SlIHjacysLcesrR
1Vsoo+Ap/HZTEaFAozWPZsfoWWM2jcj++POaJRHdUnGXEjZ4QnUm7Dam2lAd7L1R
Kv8NSeoPpVOBgxVF+bPZxP5bTro5KGgYg9lsRlDJRFMIKpoeUu+lkUB+A04M0NeI
FZAb157jKDhvrQmnRh8TJuZ1WGJfCv1NgUDkGgwLilYs5dBoWgWctwbfQJikqmej
LspZXp/ORyxM4hSwDAHdPd/Yhtp1kHlfXeMbbk/3gymRdNnEQ9xZiiyxn/TAHoYR
VseDA9yktm9nqMUOxwz8XUUfcuVZXaNO2u3eY8ompEUmS9CDntaTO7E47u1c4Msx
6nFsPdy3eLvegw6N+H2wh8ll+hxqhUtS3VRiLcsn1O5ZCY9/iBoY97AQENoKZ0gz
13rmT1MMOfZFVvW/eVbbcYlSm58M0MlqaJVK4Ah3CDrkS3d9yLw63EJ91uU2KFDb
lQ0kQKEcBxCw6l3iqUPgnQH4wtf/VzdHpkGsLg16fIjXr6PZx2UbDJTcTuQwh4ac
Cm9UL2hFc4JyIR1Qmn1N78UNGV5ih1djB9JoZBeOixiii1Fezydzho/+FNK7WzU8
viGyuz4R93BwfRxGW6iux0UD1HukST3VF9nWEn9c3QRmzI8NXt1Z4rNUR/rxwLUH
SEZWRmm7jFHOtkZ2DwwZ1Yj97ix2yzScjzoxBESCy6lD3azzlqCzDIk+zsXzkUxq
I82/lSnAE2rZdumldsIrn+NqGPq/cWwES4FfIJ7gYRvt1iIQMw1Al+OIkVln2Kjh
jLxCEPOkkv1quzeNOSKQhStyZgoUUUhklaSbnABRRfzp3r6W7q5bey4F4VIbqbyM
xrPOay345NJqbSj9LoG/DDAq9wrPigZd6T/E4EmejfpGkvan8RWv86IQPGJFdNSk
uoEbOWpyncaF8KEkmpyKd5xRDnc+9ztDGv7kdfcAsq9M21Qfr1C8JYAjWgXisP7x
AN3BC3lrOR1zFp836vnFg+vKiPZiNBiunn1TOKzMOCkDb6mB/o8WCRKOIWRRoU1X
t5Id6IKZgmX9EhzD4IMoV2bAzbemARGwkBpZl2ooMbMi2CpCQlYO37c9zvkh+2c1
ux1UIc6e7hesoaS8X+sYnBWqmWR8S0QVnw30CA4hx4tPhFAIjENbrQ/eQQJVkJUj
qS3OPeGPE6O9DW2AeWWeD8A0yVOzffNIwCjZvgxMj8v5jZWY5oT/+XBuNyHxd+rm
QHbIROfPxXVMRb83GWdgSwzNVLandzgANB+rNBDruoUAD76qoZankT/4uoIy9rvM
pTdYPu2kvpdyZ1KKI6hLsDfdVyf8r6QlXcRz5yHCuwrKnRriNsRgGvdXj7Zdsoi/
8Vgx+5iege+uUcfxR8/lyGPeGVKyFT6toSvLrCexchEawBnDQdNBysx2xwvL8gjW
uSVfyZfAPM088Kh7xLjEUkHjQbVaBRq/eD3JuLBI10R9RxzF3L17T5sBQTVH6C0f
USeQ5mVZB6w2hIIhDgMzxlJkXK9KROBdPW1x+32FzFATmHUAfqxzPkRWWuD0bAGo
MikTOdyCCIWk7Kd202xHicwQQgx8AXtU/hSQZ8kIkmhBZylBAg7HrEH8BPqwpfIv
DsLLLkEofbKUwYdyJILgj+e9CCpvc5jefQUeRW+5g8gm89/zEOontMNXRghTXKHx
GsYf2FKUFW02gYIq5oEr7Sr7rZQKjUBPUOM6Xd/7OA/Hv6N2ZyN4tOBPBfu+RKlk
VRArYuEH51vYmorh638Iz9vw9SYgiVrqAAW5bNzCWZAIOxSrp5CMRCbC4vdEDkvB
uCGMiDmH3g7ogS9lYont5PeD2V3NwtZ4/FdDv/N4v61c0imzcybb42RbdN4HsBUL
NrxmDZbf0S+TsgwRBudiaZNvhO3mmQIdEDrg0n40AQp68ERzGH1PxFMvaurms4KJ
Y9z33tYcXTzMo/gUPug3JajRuS4DlFvlYBI4v33N4aaJCb9oaNlNiNnlTVwi3lRG
1lLInn0xc4vSjULlO7IaEQWWpm+nOGebSOeJYV7GRXhmNkEyi352nL0MX11c/Pdb
NEC/JZ2WzWpcSPRPTh/SbSJmrpt2XMMY/DjzqEp1CiNQGQxYVd100Ms7IDlwdael
lX+rv2jNn2S2TjEHDwRcmVFYJgfOppWR4/5HB1oxLLd7ozbCjIf1sdkQuFYxS1Jk
Qwf5+4F/H9kjVO1WzO+AMoCaX8eD+adBWFFgm5CSmhFlxcNvo2y6OKjwAYi8lAfb
X0BqX63uM9/m8wOLRk9eF/enWj2Kj+LQSWW0/Yk9QEEnI+o7usRou9/Z1sL6XJFj
urgRB1Dr0+NTtT4WrXBFLlpxO3qLHJnWrNRejstU6WjaWHUbYyNFvJGiNQH8oV2o
pvwghwnogaeX18azRBD+krAGO36AZ1FKxgcmPW+7VL3uOBOCriIBfKNZ7A2+CX1R
83GoJk0iODN9jIXAVt8qhK/PpOovkl+hCY+7lhAujCjoWXOLAe2ZDzOOkxs77ZwT
YNqv49LQt46Ws8SZO36xfehQJLpCVei21KKAUusu6cekln7K/0p/+5JVuyiOve+G
1mOHFpShLGyhv5rguTt2h/l7ZD3Kk/Mj82QdI/ff6rqe47GTKQM+oG/qR+GlCmtT
7kzotwefGPyBr1crpz3QwY+cZLOBSfIy1ICT1EAKFx/qHYY/x03msEjHb4rNiFhK
Zp6YXlzqKSn2iyAggGqwTn0oUhxeF3tCpoieReklhed4cHYHCCk8WFxd3UINjjgc
xRzesaTfF6woPIRCcQShAwa4cwb3lxIRMxX+T5QkL587TX/6IZUk0COlY5jviMvM
KXq7DoXlKxMkgzeSUYLATok5qSHBx5XYjXynn2UgXUH1ZVcYKtvVPUQN4GAWY2+/
+0X+6oosEUSyRb5zjHZfklVQpr9JkNotql4/jmEy0pOVzmgxI2+bjd3VyMe6QHpg
qyVzKPMLc+R1XFw06zQk9eChwXjenEfRECz0IFCu72Bj6RnsfjD+sO39m6U8pp/a
h32EQrxQC6Ow/mji1wxBsgfehg/KaWomndH/4KUbCRIU7zEAXikd40vsIioARjOR
Ftafqlry08bAxEYFRQRgFUSic5auO0bmndo6q9AH2idpRenn2VxiUMUb4Qwdrd6W
1S94B3WSFWrNdS/DszPivrDkw0Vh7CcceqKT/Hk6wyenJ8GHlSQ51LQZJocjHEHf
/X9YHPc+iDPeMCfG2Fv09udgXC/kTrdARWWeAcNbFgqi+MgM1723S798sWCp/Vy8
od2mDaB83NQVAOOo+RCqq4DwGEwQwHOlkzgWGoa/QBVFdLXY7o5Cwy6O+wQSX9ML
bXed7W11unVeBsvaL+lxIIou6rX9x5dcTJGy1lIEKVFKeuYOSSMHVAesDoJEsygn
QWrQqtorSDQRYRJdkpf2ZC5VoVUMPbLF9aHhgQrFLQKUeqvXXkgNRWztbfoxVXqz
x367ahhWGdOPWBeTszavQaPsgppktxdaFynfAd2oIf85vbolwyHzOaKJ0mD/ImNC
bjJBZqJ7U0tGaLT2yGZczlGvSyv8dyCo/zH+IZQQb8jbCjjrSgz5KgbsSCHo/kti
gdKb77C/RND9l6rUhYWguxLOWs5EtpFJlhBGyDeG2eTnqIzVzH1vIHCqMtYn4dmY
toyXOG+pW/+WNlJl8q2Z2/ZXI4blbrWM04Vgr92C8ypy4s3gIv9nWb9o6Dko6S1q
ixcMyOAli3JKS8p7ecvlC16ci/Yx4rXJtGBxBQ3t3HG3gt7UfQLNPWLwNYFrZ6Ho
zbo5aOUW9UMRlUsYsHzeTzPzFPM9fmCzZThNLHji/vnQqlVo3Ckxz+m6Vn6BxTpM
Zx+qUY8ddRG1uYNVSDfdPCd4QVQjeiRrmh0lVnZiJQaYhrb5bIMac+E/UaQJsJsX
G0dLhkuzmdFRnrUknNPUzut0GMJSjj1uMFWrEa5TSWUENzVqnylykdOBufmYbr0O
CWsZXQnp/sO7AW/EQVeaw1hsk3SkLPy5276M6W5+ax1DZHvcxSJJr+XLcbe6Vf9Q
6jFiZUtHQR//jKT717S4boi1XMwlcXe9MR7GP6fSBKRhHrDG0EVjRir4sI8wEfIn
+AJ8zn+qau+JRsI+SDeM8w4boPR30HeabbeaRCMrW7C7Tu2YIVX3p4cX2cv+zbrF
FIp8PnEdFY8bTZ11BHdYwz8LRMsAFxhLmXG5IyXW8mr7Ifd5ZCouGK79lRfu0qlC
+ltsU30sWzdovBwjTP2vIrOWVk/Jk20GBjd0VCZWDOTH0BOC5/EuWj0+o8/wbo/a
FUpaSeCpQBdnzqPBfR6wzAQfucwd/vR+b9KW7rufAQhXr3xU32UaOEPQEMCrwxmk
AVZ5XA1JRqMwnenkxR2v7I5UzIPZkh/7How8YPeysQjVWrq+BehSF3rmHxv/FpnR
enrYpUXZZJUkzCqxx2TUBuxBJQgjGpg+ZRNeuYODpGtX3TrBebtLwhrlw/bLSuDw
4G7s2Sv6Pm53Mb+K7ZUhgvIYRGBxV+mLZQEqUuYYsCPGVPqsgGop0uLlupeW8fG1
mD3hRnS1N3FglFwIEhuycq/kcaeA8KwG5/hyXxhW6u0xHaFHdkQFfRiJuC9juRoT
PbpAFTkm6w6COi3S5y2b8Tz6gmur9TKH0gX1mcY5OfLiuxgAqxBJWl0s26DRfa9V
L48+BU/rBGc2AC15g7XHrSLLWjRgYf18RrV9y25MCxbU+SdQntL2RMb5Z4iRzpbq
eE3Br3xcV0NbluAUmyLgJAyIk1Bo0gW89dzX2YfAaeXC5/yPQ/swLqTJNyMxbxps
t/EmdPhsaGsJ34jQA40A5K9bLwESEtadRZQ8YlXSMxyrm9r7cUJsc5cHT/axIpcU
jt0L46hjnCLthHhSUWTBakZRRnqi1pwiEvutUydCjcxon7upU14OHEUMQc9nDEYI
yuGy6fzR6JaHudAj/WbSVvh7M6WAOz2898M/QWYKyHB84XvFukAw0W6filV76Hwp
PP/8dNXA0AwLn1oKZUwtS7POsXPsXF8/SujsWVrtNMWLyv6Vp+0lsVaDlbfJLzDz
+EGeFoj8CHAuhKKVpY8/m8bqhpPjehL4jL9BCM42rAekh+ZJIxF3ZnXH4Q6tWQmw
ts+CavHsv20/I1vY/tkVjwDTM2jbw8tKBFclBFHv/A6L6WAEvrB07WSovmjRD8Aa
0nVtmodTRoQ7rnmhqOSQ0A4FlPH9QT0Uvebt24gxh1/kBVfWu/6SF3IWVmyX4tGW
fFVUcospT7UoLNedktNu2bWgKOkqPm/ALPmZoCj8/fADPSs8SOxqj1K/rKOpaznO
kr/oZ+1cl4q6j51jf7NRnEcJbbaB4fcy9z0MvcHv4VnNZHtD86JAAk4FE+XjffQO
i07pyiaz5r4sXRpxGfNjEe0ItzybL6a9pM6ivgvPowYVpbsJ7X+w+xqnnI+UdolY
QI0qIjfxi0vlInRB9ZW8YF3DpseK0oLwYuRTVB6TU6Q+OkGhkt2p2qIhLlmeW6C+
uNI4uk5y4hORbzznjHsN3aET+qf5iSxM3/c+acyur77yjnwSKWaMZd3+bhgsUWIh
heo/wXQCBjE27C1CLvtQeG97QeKqiyPeV98h3BL8HZZA82rHq2uZk1eDmQe7TUsZ
7bVLMh6J9qKlmmnaDvRamcz3iyNpdMNiabQa1Nq0YB2KypljFtFLJHpqtAkRpdd2
iIvZjbb4f8x4p51YwXkVzZUfnZfdofwGNGe7IwQh8bFxarm+nfJIax3vspQeYTFu
yszt1793LiODjp2bV/4y/Vlfp3n+Pf/cYfDyiPHBCmi4dbw4fLit2L47TajheWxy
70tnLtltuOErwTOoVZJ2bDR/rEr0rWrfYxQwFmSrU/48lj5NL6N4jKiVdv6Y1d7H
/Q8N5Z6dGFS4ybl1PrBjr70ugEgUHwxy/5j+TxBfLszVP6ttNNYhIzgEYLNZPPIu
OWkzRBhQxC118oiP5f3m6n9H8JHyAfbNnlGEcyzFkZBWrF2/MXGBV5O5kqIR1Afh
ceF1mz2BdzrYyy0q6+TuZ2psv1ji8vqrGw/s1QhumXK8+wJXo4SidnqWdVP2KbdJ
ZoBnmHLt/339a3Vte06FgCMjWEPTDugr/2oL2hAl2/5ZhZoXYaYyGL0JHM1ZDSR4
MwRRcK3UblpBX0HdTnaEg0w6vm/PGpctxZdYxmxfTcnah9W5CGorvxDN7ayc1Ngc
V6Z5uhuNZOXQer4pbsvVYq+zKb7GI16SLhdTxBXGVPQrD3YkAaJs3fq4Suqcwtuv
uKeCfuXrEX9xa4dDIPIZ2/CFKc56h+yQK+lDgjGkRR8JMtFJbnqokPHQGdZwOxic
ZWYn/TWMj/8nhj4n+Z2PrZZXTLTr1BlFVv01WewUx9hsZUIBlFUDGIZXQmaRDIlr
md4v6dk8cG1r3sGoa7ESU+WzOTyNVS0SyEx8J9BfvrX0UaeNWvyD1l3JzhMcnlKD
YWYRUCl5Feqw6iY4y/erwBKS20nxtIkV+oEluQr8jUuL+lbOdnG4K14QV76uBPYX
ZIKNSbHZnzCOOrqZ72KOiaD7lc8iK0qM6WVySrBxl2Wn359c/IygregbYHzclVKP
bhWyTTmeIgAj+AqUD3iUtQ0VtmreCVn+qlBdLfcjVO+mMjG4gbHqzVlxMPMz/PTA
ZcJa+9LayCDeqOJ99VINMHKglp7gxDQ5ZPUQSkqFaSmNeptkF/VFgKz05L9H+KWy
qXUro1Re0hEimp+SP7Gs4FK4oAR9h1UXBIMOhkLLs6E0SNdxRICJ151eTaY0OgQS
KIbNaOZncg/RTlZJa1+0hEniHbtK5FMmbRITbCwyqxuOlMzXNUl0x4w/oPNYFieC
k9m8sPqwU2+LbyzmmMBPF4TZMimNik+Fp56lhGH+E5VPkPU1SpOZJ+UTwSvRnTs+
nc5kRqfMVK+vEbuPMK9J+GD/nZREP67PCcPFerEvPoi9zeI+vDgHSJPvsbivDcaw
qZ8P8sjVdyIDV2XW7fxc2naEnIZy74nwSxP7+OzDGK8XraetAmcKmh6bVf2Q1gF+
YTIW9ask663y5QyyuMNvhr/Obeg1/TobsuAuPMlBDlGdLt0/mvEqSsJr7VPQYY67
cwWIwX9spRO2eekubPt7328nbceq29jy7LGLoaaDAf7Vsu83DcDbC+cCDRUviSxG
EEOyM+ULWalirG2xRtg6S4HZ+SRrbM1rYRKr/FzNheJA5SSFZHBqDkN6yBHdILXa
OxfL/I0rZhhModJd0ZYf1ix6XNGCGrqbSJr9ASsR72cdYPDZO/9wkSkp1TMHtsXK
Z4/QsSh8QgFKzbHDmjWIv/smmFTMNlY7sr17f+Q8Wd2TMAj6IUayO2jqKzzexyHL
8bzzG4D+kSYYYZuurikjHMIXzAV76YLaW6rk7H2pHJQTip7Vh1oQ0IrzTotXaVyw
l7E51YdoclHC0eUo1RCsaJtCVwj4qO+FkCu04uTqWOKF5JYO/xLZyiM+yfsOIuA/
prRSHy/pVL96UVj0CtjLgKz5zhf5MkyG9DHlazJqDmFIAVfvHf+xadvDHx1ZNcl9
uwAjqYz0FYwJsGq/2rpJuGEPxvPtzc/498pjwiWhg1AsCzTdSDS2qsL0lI7mrizH
qHq0FbkuHvAAvZ8WzcHXgKNfNQEVIQEmYvza3qm5vIj987+Tbn+l1lIS+XbHfG/N
z2XoD0FWPT5ROYhSOy1pPAuU2oUvdoETxMGtynA94C32Viuuyr+WtKmabuNRgZlF
aJjQ2tXy5GM9ACprZ9S5iMcKUDK8ATGW1kXM7hep8X6ApCW7cuu/Fu/EALSvtswk
tAoY9oMKiMNWQsZabhnD1dO29QsvfhLmgNWm4pSVDhBFlLeJPSTDiwN2He1xFtqi
J9JUvHLJTQYTlDySAhNR4VrGR0DHPw2I6qN/p3mmPSM2cXmY+/Ywm1YPeYazZkrT
xgQNyixM2xju3rGsE9JJ783U5ea6T0iIVhWDmN7th80TjvGnJJZWFg+kdhisYtj6
C66W9mNdNF23usLoutEaUHBsaf0sSCKh9WXIuDEicE96Ax0WwMCkYo+y+yi1EhSL
F2XESCjqLYscV9myPxnS8TPB/2Pj93TQUfN54dhLfw6uxoGfHUPn5qSyO++24mEO
Wc8IsjacpJQVPQhYLk5Z8Z16/NTX/WJ7cg1MPLOsI3BfAl4Z1ml1ddLPeX/ooWDK
1URg//ZKQpmJojTTCfJQvCmW2pMcq21X5CQRXV+Eo4pLjECMgi3Y4e+MB8c3VxhL
fdyG6uATD9pVD6RrullHTCLMjTMa3aqjhF6zLZhUK0voMvNK3oNwkO6DWjFiBo7F
/WVsiCoky2JpkRdWw9xypiciPTg64PBRw+Oi+qIMm+yD/d3qlvAjaFQ/KwKRGELI
bJds+tavVoJKbH+kUGrdA7sEmwTfh12LeZvjGdHA0Z8Ip/Gq6KjxOhBxrwsYxSc9
2yNjV4dMRwac57jCl4Z06nz7c3XPoSeOFHpSHWHCUkXGdeJ5tqhLfNf1Bp3DlwFM
Xe6KwuVBLDcGXyqMu7t7MmQOFZGqJUhbJtUNwM8ZgYS5cmYPejiuSarbAPUF78ov
/omzA2FNg2qh61+VTVHktSbNpClUS9FlM5IezGFvZLzk6Vtti07ge5caiaQJe9z5
GKd1Xbjz6N0YW6UKz5ARL+uatBwuXbWjXnHKvlv8glo2B9U5Bz5RrNhk9OFyq3tG
f18XZ6nODQRL4EQaA3aGd4mxHsUU6JV/vtMYCKsqmkHazwJQplD6zffSqfeEnc5T
Jq4HCI/uQ+7Uya9u6PXA02uU5dBehG+4W1mIi4vKWV+LZ1KJBDF4eDk/ssx+g6Rl
pEMjh9TI8zemx0pNYSDIqoobsQKKtbAujDJolLyA2+HUIssMdOi109+64fCxojMr
PKfBSrkLig8kXRjg/ZGCK52GEAmuPpUl7fYAmWlPOuIq3rg4AUbcP144K1mCLBCE
0VaGoSj9jzXPSoZCnMBbHUZj4U5nKNnDzdOjuT0t1Lwal49aOHZ+ZjFd+AQE6zM9
gN7epcuQ0IhAhRZBCKZBfwzIzWIA35UyQHm6J0fYkaayMvlcstKIRAbAcS0ItJ/+
1NI7pjHcCPUEwNtZAmG7hbmq7kP3LlFGaji7bEPGxb2gn+1yVuPl+1dqYqFpeRhg
tQpZT5/hXck8X4Yy7AQAQVZmrvlC/ddBdAgHlfi9I/jSQQcWbHt+3jPxSj2rNxFI
TNjDHharWrGRRtRbY1vPPzsviFLIwfDgZzm0tiRqcF8jJxWqgDXFdZzfFJoZ7acn
J05BtWhnL2D66bvjEm/chRz1+lKzd3d2wEUVNSx1YFqO7LEtCb5pkjHzzZ7sRkKX
aOQCE0ENDnaCWi0enpqoFPEAqjT8tx6VI/ttcFy+Pon7IxfrMmZqkqeUXFqjD/2h
tg2iybbf7qnvPGyEtHEVra06OF58OVA2jIV5dFyVRfi+TvpIpB5+KZ4EqEaRYTi+
c8l4km8dP23f1oZnHORITwOUMMp626/vTTwTfrA7Wj1/MbdpYRqQrAYyZu77/CbO
EO45x66a9OCGclIL+cIAX2I+yeGbEmBIA7FBKxfVFv/XsuaoJ5oQ9kCtCIbmsrYA
UA6zbpaSdZJlRVlx8LxzWnmYCsqtKc3Cjo9xkhFitjcGC+imXVB+NhvSKTCJrvJr
KRNpTvWdRjp8EQTDCJtInNyG7hTeS0u97oNW1+4UiTUQZ6+EOrsVgwC4IDlSFS43
llCiEABBNeIHMHTjmyDqnE0vpdnUtnJlWQdLc+lwFG/5c6kQcV4rrfpw63/rS6ui
zjPRpr5tUFnxpHHP95jVx/fY1RP4irLL32BkmlNkugz+Bv9PCgloB0HA810Kht2s
shFFzHgWpg9hcuzlDITAsi15ERf7tlL3ccWfUWM9ppXOj0fKgS9NeTGfbpKkNOQ7
SM9ux5SS/Tp+vniWEezNKGWfXEQFoT2drxzGm01qGAgLO/gOMfaUHDe6BAvQXA0A
aSl/YPBcK4b15ko6Y4uIaqC7dz+uIj+8jW6IMb4WXXtsdFx10Mecg9IsDOJWsS7/
X+lnMzm57N2AIWhAs+9FnaSAz7bg3Qmi1TxGQp4t/qaVC2a3WLfn3b1i1SHsH5NX
QlpU4hmSAvh6ngJLakXn8BqLdLYFZt1+z2gwIYc7zBIY7zBl979XwBpq1UM/oQfH
QF3BnIuzdxSRajAfPyjLHORNGi/U0Xl/Xf37P3jI4yEo+T9HlAraQk6ctNS+Rm96
v5l5GHksCu2AT/bgvcM1KH9lrRG9S1RE0J2kKW0MrW28Q1z6zZLjfDvDS9y3F3R0
dInGT0R43nFRBFwLZdU1j2ujz2kZEEuovyHnsqs7K0vlVVUYnjxZcIYgClcR2a8p
dc2xUMo56RULUVuyeWidQeAdLDMbiCS6Kz8g9unT32CnHA8SSgZXFJF9U53GhWiY
64iFZClFB/DuT3gL7ciP1pwi0ZOThxmwfiY4m3giBkK3GYBOXdz2QdFdbBQDvC/b
9O2ySGsmdGmJf++G5KdbqAynHQZBUABFCx2pLDHcK+hq3dS2u5Wvg4o7czacZBUs
ECeotlXSqGK613pQX2TRIpD4+a1ekYyjWlNH0UF3zUrgIy3rVt882G/n0pswJVs4
YqsF94AcjQ41E3ClSN9ukwWDVAdcf90nRZvDm/P+Z9vsAQkiDUUP064r71qU2N8R
f04VsqUEvJKzqV8kxZArk9lrgwAaaMe910Z6mnNLHTfYsvko49nDXbKtapgCwKlD
fBbni2IzocMAPznY5OSbckZeWrHJKtve9wWe74wnTejAfW2AUGkC+Vh69ETSJ+7W
wZ0E/mJ1OuBWVL2qya36KtvxXRrrplXzJLileH8ViXTokigA3PSDqrrCrQQ04TiG
hwH8E/XF9cQ9ssxbqB1oeOj4Rl0QGHDX8dTJTYP7cNHXsroTTCs4HDpqt4WGrtbw
1dplitVzFIO+GHQSu0coG3/xYCv3GlEsCYhCYAr4ZJ4l7t6LPwlQC5ZnEwP6cpRK
9TbEaT2lJ6UoR62sc/rTuEzhllj6JmgitsvnmnroYf3GR4bO74G4m9LNug8aWLyt
xhcPBeqHhhFl5aKjihbDGXAprPWJK6wUGurN79sZPNddZ+bkkKAmdlaleLE4323d
a1aYkq7xc3yEfDShOjGuwA6tcSMakt7idScJVbMX0dXmdvn+g4Ji3YPLACWGfkhX
39IULYhSXssXv1UK+LFMVYhNbJBH9Jk+sCBzfG5+qh8BbdPiq3i+Ol52h5TlEJkc
rDznFQDoJJWNmwDTol8Y5PjwqdFbGXPEmYoiKyxipgkIag36uzozrymsn63h5hm0
vvzwWXW7LnYKqNqXwVcslkAkOTKgMso+K34C5X0TxkQSSOw98b1l4PFzO8srebY3
vhsFC4JPxVy6xhNVtJtgWGHjT2r9H+HDtYExiZ51G1CkS9MTiv2ZY4wYKnvx2dTh
YNRo+k9T4lbifO7C/9TJZM2otM26W2WYD9NIhITUix+SknX7o3kClBzrxMbOnUJd
qTM3hI+VUL3W6G6Gxy0nQ/GxPSCHRI5g3ZqnkOT8i5oER6FbO1cen7GuPoPA2Q/5
YQ3JL8BZigkxMxhoFBX/2gPZuCV8JqWm9Md22RLB1e8UeQpIthMp0QGzOyYtLLQU
GCp4w37rqxe2QxWrSabGVqHzoMBrh9i9xr+MyQJH4JfFoc1ySHXssk0yRE47sKa1
2skGjo+WHq0slYdHKkQpruMGPx6pmUD5bg7sKlLwgtU+t/O8YtnBvw7u8FGAfvPd
vJVSBwqtgIiveWr6ItJHfEYP+I9ioVgmZCdKFo9ndR1N/fDvkNM8YFKGMvyUiUss
XgwNfKgyNn8lq06GE9uQtKH6Djc3nspr8TumAt8n2E13aNy8ELTm1uxB+tLtYeUq
B8JJdDDZ1NX5jkgqVHfLf3fiSFF83eKw3cqt20NOq7eh967CQnY0NdaQU1m+LAc0
B5DTwiNZazG9UM4fh06Ve+cxTPC2C/o75yJw8j27/b5+egyLniSqZxgwKEoZf9Fn
31G9KJg059udMmC94OltaPAHhrcO/LE9t1vUoQI327LUOAawXo+nMFbwXKo48szX
BJj5JI+VScVQfx/7z+9RW9aPULt6IgbaqpeF3M22PcuHLri7T8pwrT81AWr6shPQ
AXvjDD0Clx4CHSoTAFwkAusqPbGtrHkWbXk1fdYRysQGs1n5nH1b+xmSRAbAonmH
psKbFKazBN4CP8xK1FGcHeGjCClhTTtSq6Jh/dPkU4lFmFQ9xne6Y9Df9dXCa5+7
Y3rCPHMCw+8E8xaXpbJR2BHbwqTWxkw/zZ0lMncsFfpIBltp/+xF7aeAZEfDpJKz
GmpCix9RVYjXKrRbjf8LCOyvliJquxlqBkCSvRfzthd1pyuA0FhEPouZfjgUc9rU
Pdh3Gh/Dc+CN1b7SYamtVqS2DZ+0I/lK8B1EXcEcGu9YDIsmEuDgnOxT8ZmI1IcR
g5IPqOlq3uFAYVIZHdNx8XZO4Xgy36uhN5EGYEd2KWCtm17dkWkw+6ql9UwKm7F/
ZdYWPmNtdoSbNo+j5MRQLuwbdrKz8hPiVcSRq4HX9EtCsdi1Nh7WfToNNGzwcFR/
dbfoGjlTg3LU95YXJrCkkZbQDO6GJyVQfeU8AU2yw/t6dVFMYCCD+Re0Ff8c7yrI
sKf1LJfdu/9bqsm0wwMg1hO6avWywjdDPN3fGBx9LamH9g4hHlP1pdTCCoj4JFK3
S2s8eaEmcvcf4cs8otngUMlJQaURuC98JqkIqJPsFEgvh7/GNHTd6X+VYNQgPKYQ
Hvkr4CeceKmoOHx684dWcP5UMGTSsWOpy+ofE2NhvjfgHg+ovRSlnbgQXpHjg1Rl
SffTGc/+B3ziEj0DZqIadiejdM+g1F2BAe3c9X2ngeXMaL5cMSZjnyTXKaSB1tmd
r53BKtvInyXyWG0BL5WFS4LmM2FIxkJghEk9Ibn6+yhGQs6GSZ2OSd5SPKlrv4Cd
ZzEIm7gmZMB6LpQ7c3ayQchHQgVaMnl2Ykx8FfNAOslbVyC55WlGicWwFnbzeR2Q
XfJwXRYUS0D+fRKUKCwpnVfiEMScFfCppiKSPHvF43G+Fjbf2rRVTgIsMcN1YyQE
IXqtvWPhY46XDu/4svFBcovuASRHULnB5bu0VFtq6Y9TUNCR0StPSDAmGIhvHHUh
QvrNQqiojtr+C4b08h6HWQkZ3Ferg+Tm8gpC/YQl40DnvyR7bPHFvd/hklLlJuI4
APJ034uKly8gJgFvMj9jKd+knjPP2w9LcBBuouiiO1sCYu8CNc/Q4PkIX/h/LUrl
jPueylITe276JKme5SJFpLaNvtfB5DCOy++Rbwp+jvNd6CNcrV5NjDOljEtPa/q/
IMyBjKFIhK+xTD4TvPbgmup/L7y+ftbUKgXYUJB77wo7jEzn+lajWcr7fNjjBQP6
AOoFz+eP5mB1+wSHeo+vpewqdxif9w3BlWQmur+nGinNfVBAWSKyycXhTUiIbAd5
zazSKeIjt9tBFu9+3m+e9GCYLHEbrx4VqA30sEjRBObDNFKqJHUk8EubPWwRaXEm
wrXpXrP5s4oQud5h7EzuHaY2s9Xf60Gzh7rFfWegRI0ARscbSye1reD1kdZR0SIQ
jPwoxOIjRpIzbgrKUKPZ/IfCyMfuXUYoJ9xnh3seM5noD5WTu9KQrHa0LR6r5Stf
qU72ZdF1xbBgTEWZg5BcSmdTwkgSBnbLjxUYM9Ry8l9CjyqaGpK+2YzhV0x+GhZ5
KTmZwbz0kCfkPqqU2oUC2S81Yy26wFXtCvPnIKZ+0n/HBRF83bo7IV91zQAGIUMR
lQSikXaAQ/M9OJbtYS5CBVv9XsoGxEycsPh224VLH7z2g1ZxOi6E4J+iEorR2bjL
RFiBlKHln3nGRzB28A+kqVAZdRmXf69qg7i2MgSQvANRmMI+pLk26AdAQhnViyxa
+Yh/siPqh+ybf5ftQ7LYffUI2NMUTeAQHplG0Duff8CFl7USLx6jnkYN/l7pkzko
pmkOoMbC93BovR72cqOJ/9p1Slw2a52wOHFqKoIwwmyT9k20irB2X+zLVIpNl/OU
qZt4ynXNgdpM+SXCoH7mjjty+8juv1lwBkDfuPcLv2BL3N606Dx3Zomvs4l35hQe
6y7UEcDfQM2vuuzm/108CsIYpJMlyaGuhjvwu6nF01CajTTyGc4FTZWIjxuRGxtO
tsi6ac6fJRFch8dX3YWUzOc1WdubfAO9HhIiWKIQvCFmvdyHXQdgBbF7pOj++gZf
XXAlRzsn4Gexqz3aFw6KH6x43XMdG9WNIQg2S0zG2fJ0IJEJ2E4uT2/7EaSjwi+P
wtIMSIeI3a1EVnCXwmTGNHPrtWZMKaVuE9xxoDUITMqP7s4h1LwhS8G4m2FuU8MH
AsQRd8hbBi7FxOimDEyFUoWUQvVUFbTfSqhM2ie+43eTMYtQaeHT222LkYHupZjx
dF9u6LrZN58NLfXOo24vyhkZOQWSX/C3qLPrf8oi1UvmEQHXsyurUMklubgcrkFw
pn3bdkGnpatD8a1F/iPHJdAL9rckzXT4M/8sD8QgFG4T+iuBQGzs9x1BhiQgeCdX
bIfBlNJRoJpQA5W1P023a8CemVtpMg+/+Bf0uVRr1XtqWbYCb0SoW6SpbzzD64FW
Tlbq8aqV2Y/lo+JASc3lyNn2bo3fpVSnEYpk00VRlljcp2X7MULqUuBi5hn7RJdq
F646n2YI9UG9Z+aoUvxHci/YZB7nX5KCiF+3mG6cNJ3voSsmLO2L7SOZPsAgjg5N
74GS28inoSqb3/LysZrAEesDS2c/06OI9PLneDysRWJFNueJXSwUNIUA8cGl5ed/
p3OTHapaY79E+DZ2N7JD6LpeAE2cNwRhjzItjjhP/DTL7Et9ooSZKFxkwETDgbVj
or5QBFWLsID+TMWtaTTgSah38g+/PIYwQstXHfETzXIGd0uDeeWqU2fcg69MYdRC
YAAWm//tvoGAs/8LZ7tKDnorW7X9gAsxpvjLvlHP3YFUQBDSb9903xtGBVnGCQ8l
hRTOcOzCeV+IicTWrugwp+toFsT3ugWtZ7Ut0m29o8BS8SOvlBKzM0lngVxO8qR7
L9YD9LYMsnVSB/M0botw+0OhI6By5s0ch4jdgkdAZIfrqHeVo7mncBawT1MQj28A
eQcnVDy8oM3n2SytYfWJ5kL7mBMOBuYGLKp1SmwTjcZNxF+3zStLM1dbI5WHWPHJ
adNJpr8yuxTnDvp/byevqYr9KUjOlV0u68sg9XjhWQ4Z2zhW69Y/K9fJtJlB8jIU
NAQvxyiSEC/7qq9/lB6MH4lwX0sL3HwjMXOo+2+xAPlswH3WLemkeka8AUsj3erR
95wBKTkQzhVxGERV584ap6XasOcBUvyVOotFtrqAq8/yJq1HJBlY6QCMM1P3oAgJ
qxHLt73vML5lZba1LweR6cYhv0gCNSs89o2TUdUEkK6tcoQt1NFEe1cYtR/eaPW5
rDIMcj3vtvMOfbaBwt6JL4ZyGY0wk7WPUMMd1OCX41uoEtYg532GOx1VT/d0WpJa
jYnw47HFSc0NWu95H0y72aJ2+CXDEVVOTKeU2jss1Ps19BHXLudJ3X05wwOC9tJ+
k+FdZDkzJgL/KouN5KWF/hPLWFc9kcCnRnS7p+W+gJdxMIxXP3TpjbkmJ3wrIdOr
nVAUIBZRF4oX52booYJTMvllquDuUvq8XUmBhrkfa19vhGPBnaEXh5MTfrN2I/P0
bf4592szAf5mWXZGMvnQZfesjJGsgdl5GRsudVCXQb83zOugr7woy0JCdnaLMMYM
nQi3YPD4P5seCXch4ZRvv2as8qUdt4RPjuoYCEPL99JLwmfhO/jHxC0nZHMx0EOz
TX3e++wOrtL8rgjitCrQubZjehT6AJ8iCK/usSePsTxgvtu8kGd91q0xawuXR3J6
OuXBEel3NGYRIwC0lR166zpoMr53bxQCtWKLDu5tL8eG++/n4+lgURdjoClfAqh8
c6foY7kAdPbmd4W4S2jUdyQzB46iYWvOL3HHYE475dCuBcleAcd1C0iJ0eLN1hcE
sGwHH49v8HPmAdzaTmaf2g2pgfjWBvdnTD0Dr2CIKongGhT88pROMp79cAt5nl/d
LaZdya65jNqfgzpi3qnj4QoLIC5ALR4+JUcHh2I4VBkyB225GMhJyHSIlrAr69Rj
NThoxX0XwYxHwB5nvsHgieY6UVwYtYvEjw14c6DE6+Ly1LsgcF2Z3AKxF3xdIA6g
xSCFfgPgkhrQ/ZcVX3ha5Owb5jJBjEQvf6PRozPN0jL7DYserX5JaXDe3HOABSVX
qeOe9CcZbjlL9er9ZtDgVLBxjDXisATJZ2vzVc1FsOjN7djj3NBVO76RSrURDGPY
eT+PfQVoS2mCSi3lPm823+VdegY/A0awPKPcxbSWnN4zk0Ln7j9ml1jGiDMj82zk
MR+aXzwtoJAHp/RYDLOwB0pzn436vbGXoh1YoxuZsSVtbKrUXGVvcBOhhVWTJs4+
29XK49pMo8cYGGiLgG3dCVtNfeOzFkGFY2pPLE9BE+RR7TT/fZIQCnOHHw4zCyOi
gbetUXV7bBNl3ci9wsTOplDWMIeUcOO1nS7RDQ5vBv+aHMT8n0g60nkyQvHpkVJ9
DWIrcLb7FdqaNErgOOGTQXkR+As+YBBplaQjQ9ocV4gPGqIJFYaS3qidjOfqo7U8
mq9OE7GsGWqPDggfB6kxfeguodSpqBjsIJdvdT/VCa0s6eMf8qUKuxDvYx8zvyOM
m4Agbw/BPr0mtHQsAD/hbxEkjuy8yaSFjxFQbyoaeR6hrpi7/n9LNoa5niTxlIh6
VHTa0EaopCfU0J+cz+kQSEF2JgW+ZsOlesHP1LXAwmYEntDkjdFtFKaE9ZRlfDpc
TL1vBljbnPVE4u66HMTixAqNzoRDQI1L4omumRFo/eHa1zz5ByP09yr3et6mqQLr
YOWylvqew0fEcZno96jxXNiav7uWr2xGK+fhS2mV/dwLcs17U4Q1onMbcwnXtpOO
yrq1gMZQNFyb1dufQH7ujxU3GYeEqfJ8vEMnBUKPEOaUHOs4elfuYIZ7wDPuyNGn
0zo8GAhSLkuC6yiIAd6XZBN/5g1WjzF4G8454cEbraYWeA2BKQLi7hhU8vaK6ScL
dUO4AC9QasJoiRq4lNWgs82JPvLm6E51yHN6XMVnDnmbQGS+2TQKh4gO3lVwUoBh
JbanNxgj8qLco4oO/YJyOxbp04QMKhBR8fAJjQSucgpYtjmm9krT91jt8rh/cglX
oXhah77tYBZsDtj+4XKgC3eJ8pV3r/jE6N6HMOws/qLHs4BZU8WsMC4ShSzTOUR9
CQUB2bwm8kQqaWBP/ofdZxboe2ubDgaSiAKuaFj8KnBcOhKqZ5RVaR1eWqT2lnjf
IOS+7QhIil+iMnLs+uu0vhJbQtONFVMPVMjpHftW3NZteD1k4L/npoWGlBBxY3Dk
FyMyFc8oG0GULoC+CQGQfD4PB9YRZFcegRU3NkWtIrnImy9AT5B16ctSGWvbH+t3
YCjwHT0Ui+ecH6kC4ZSlSjPUw8cCz+GhEYuxaiDW67W1DXGwhipEu4GRxPXL6unB
4UX7pcfj6Nw0sfcYU1pPyeAFqzDl69bd4O/D8Rl6wMcZEK0vUS8TjLVdwfnn6fo8
LjhPd1Cpsug31bp/vivo1dI7lF85JMexiZmiHRlbU6IJIu7anSOxbklUSn7JgIaf
CKjKCkjMaD1xCN3/zLA4oyeYQdSahr7mV4HvHxEb6eCkFsR96s0Ii15e3HqrifR0
fadNKIr5/pDcVvZ/RLU8IRtaqUW2WcTsZ0rpc39pvxraTU84/HxzO8gPbkOOP8o0
fb1VIrZaHtnWcXIsmNGC1hU4vOy30wa+nre5OIBR19Jt1RhDFu6TSpuMMV9fGCb3
OzVhxPxcnYszNr/g0LEdnXuKL1She/56/L2g3Bayq9o9j45GkpEPX6rTjwOyQiTZ
ZRLPTPYWd8Y69k+nAeGf8oUmRL7Yg2BwipFN0KtoZ/SvNK1rzqAPVwYdpVON3gCX
c25s6VTb33hoQ5mn09fz/PT2D3ubWrtE+da8pJrv1ArZ1GjxkgHYZb7ejMf8m7L6
u3hl15HOIIJeSMY3fkbv3C2tElcWSKbI+vJusL42RMRZmtnwbNZAYCgcuxnnARFx
SDORh4Gd8qu0RfoMKSzXctzaN+jDH9EkpqXgQBdW/lP3EfZpLxioQKsArkMh2V+J
H+6DCOFAWMJWZOQLMFh2JWW49YFiIx+qMQWVfwA7xXRJD0tjgY/4by7z2nuMmmYZ
IfPKXV/wCl+Ovi1tOsXGsVYsKT8jzSGATiZOGe5UH3hMvV1z8FbMi6WJZW7zxucV
SSa65ddo5s96CMxy5EJBz+dDjc5hA0G95sCZ3sfwY++r6cy0F+HaepzgeSm+QO4d
eUYblimb3AB+sc6I6agGuDS/jSGMMOOAgYMA3UtOWTO8nMegFwodtiOk7GIgsM0O
QcAMsfiDCo7zwpzO9fUF7hUu+a1Cp8wKH7Zryc0e2bA2C7VqLzV3QupxAvdqwdP2
s4GtyAyqMsGU/80AJ7EXjgg7fWvd5/miT1OwXQyBRG1ZIWrHmIUS47TelZGb5/0G
rupXfEWenF2DsXfi4tRioOO2K93E7QL9r/4cTTukyoPN9Rhl7LVe5gga4LQv1Ouj
Yt2uoqdxEJ5DTYXmrakx9ItKa3i1fzL8AEOSiRMWXTpanv+292RWC2DyHtKkfDeL
n1+mJQJPNdYD+uUAqOT3SkrSf+FRkwUsmh5Q/KJ9M5l3Bs1BEYbp4gjdXLVLbeF/
Rp3lHu/ISpVhE83/fOPr9TM3CbxFloPsRCWv5E6rQAzoPWXHRtt9etK0VfNQwWHb
4hYp59ha8DReW6Y7+EcWmmjn+6wa8T/BlW/2utPp4so20U4DK85uioZn76PbHkM/
fZStZeCDvNncN8cl5328NaO+/3vx+HrMffdtIAUcsRnJNSeVQBuZ9UwL5C8rIRM/
rduvys9lNa74d0q+eucBIYU++FJ1werAa2hlBtvtwEkMDnSduI4R6279ki5mltjw
OzPkH62NdkeZpZLyMFeSNzL4iSZ4O3VHPoD8Wz9b5FsCCBD9rGFWH+PWXxnvjouD
oSyB8btFB/BebK7avq3UnunAysR3x5sqvPYZl6NQXow/cHur75Ayn+WC4AP13aQl
d91WANetkuXEmYlnLi44jm1igbho23zP3MNgZB5v49NZ1mPkBkYTtTrns7MsVPLD
bm4ONB1GKA+2bkLGmZh6zTrDQe2U9oLqByMgm8abve/H3U3LmcnUG9M1pULWqiLi
G/z8PLWJAIyp+v/4t4RDW6UUCofH4fFwfhEo5grF6boMyn9bcWEWlIPhMvg4Kcqs
/IgjiKejaHgWXNrlQs9fYcZFQOqs1a4QIEcSzr6fYxVWEX4wTiF5A2cWbeeCewgm
51Wa+z6Jz8qE/Xv9LijGEd7C6iljpabtKSJbu/CM1n4PYUfwYSiuxcK5O1iOFJrw
Nhr78yC/fLJwRAjuXrHST23ADV1BK8yJmptgTb/oNbmwgcsrhSKGvgQVhx0usPs3
z2j0cQng+nWBgoMn3murX6VVdmScgcsiQO4F+DGuMYaRxGDo7goxVy2EMsawD4CA
nRPsB/3ubZ87gOnuLaBnNFRIYsCNQ/lx5+IFN+gO8kqUTd8FIaO/St4M8YObvoHu
5OxP2jSLiSBEvRf39rc41xKpwma11XQ9CeCqAyQrI7Q9wISVcHpCUQoVtPba0wov
1rB6vUfW1t0q8B496TpJOx2qsjbAaq11oXBTWpW8Fi3hrNmPMrlwcHmRK812EEGB
EA0dwsTrNEg4BDuaj6eP93vkHX+823hui+4ZF1bAC/HgnWt0ZoJOa29CmpWPQSSx
XZ5SYSJnOuCvmVBW1J0hQ+Iwh3lTiAdM2l14WpdDTMYMnhiNmaoj0/sTY3zX8BZs
DrNqPhVnzUTjDAGauY9fLyKmKTvBffqyq0C+ls7s5cQT3BBrL+U/aLGcah7+2rlZ
lKKceHvIZEVlut3fYEwwJZ+OURdQvvUg5cLNqmZco90al3zMuSiPQa9kcfVC/ZUx
5vNemGzTAo8XjgSmQ3dGsCsnz+lO3ZAirp2JKOcqrt2T7gSUFtqZ3Uj4Tvp3PXv2
57gNSfF7VE2sqLsBLEFQd83yxtKdYCYavqFzK+dcSJRLVO6LIKNTttfqibBwr8su
ZKqq6NJo52wW5zlMUnncSqpNIdtY57VnwV2VI8cuALphQOoIpkdLmKz2i37NIywq
zZWDxZl/hhhk7WmF0b3stVRsv3BNNMOcit5AtwhDZ4nNrrzP7mq1RyJNc+i8reng
BSz6bizfUTjo8P7F2LyZ9DklPcFYjMZ43YADizmyhhBgMHdCmRdYBq2tM0b8vF6X
YnkBAAFNi794BlKlGhzrCJPK8cZja+Bo/wmqraJ0yz2/Hks3jF93Hxv6kj3d2fQd
1c7f763YzMJVoW9ua+UzGIWkzN/Nga4PKcqvziTrTte7fkRa3uvzfY4VV1kyA9KT
YqWouDE9dUHW1L48zYWMfSxylESxIQlnGpZsyqf6SWlmcfMbcVBrVpYRT797CJYK
jGYgutCNxMI5IEreInnHLM9GMvY25gJp4OXuehvSO84U13ziY39d/sIcl3VtatBB
mbYVkdxeD1mnCmxIVY8llPaETeMCzJbQx2TannFyQN9W4Io4/GIFe3vOkmYRQp+J
S6uOSX685tnKTGrVoxXWuEt5BcRF804/EaHMfyXDq5xY7xW/Gx4fBXPzC5iMSnZV
RYuIaJLGWady1yPHV3EsOotvw32VDYZ5Lp9jk1/CkXDmoqb997pcsXFCAt99WRQ9
r02/JzK41AB0fOGO0YGNv/ybGRdzyNhxNreZfxw+YYEyv5zLpq7wzCEfprjeAzuo
OCq4cSJI95b3CBOmCQS/sdtr+jwn/qlIlgShP5E+cTQ31wzl1cAp9+/kD2fufWvH
1Ak70SeRTXUKjhcaJ1TrY3UyZbxunBfUIFo+VXRQVA+/LJahqpIGYhuC51gq3PdI
EOL048q4EE1nfcV4Epio3Ui62VEO5u4L1rX7uvMvV5SF11Awq2hHW0VdqpgplyqN
NUjC4PsKqUX9zyurh319epzL+TFKJdURZdFWzyfhjKNqucTrJwOX0n9vc92VCpaR
mAldHmPC0Lef/zrAZirpYrzelh7RX0LaBkcv1iLWW1G2er0GKyRyKz3SGdnKA1mc
Z+esiL0p4SOPlTC9Zp/v51I6ljUeS/Lt6aOJ7nNQ8AT1e+EWX5MftDbre29Q+3ZB
kTSVOd8rZbDzk5gLHHXeucxXW8LhGd+1IYncTDU4ztNVBsQjjFM0zEVnC6GLq/Xn
5gbrCua8boUdLRcV6sR03q35RkSiaruUXuUSz4L0DTQ0HlPFOdNxHKZt5YNxbCni
53b/A1zseB6J0b5yhXEN89SgFcpYyfHJ2dc+7M/eYnawnJe1GoY5+OtZt6tgRb/T
rXeGQsukOqFu2bmHqlSHW4k1moFH1IYHHAkbhFG+Ce1B+KlQWY0/Y7klbF8DGAcD
DGN+V/0dRFnxkLtOK1TGMgJeLaEcCd6S6+9a3azgI9ZyioPeDpc1GNxm5huvtP+7
dCBrcBq0Qb17N8cTVn9+cG0LfreWhwxYObLRTTshpJeFe9HICqbQqJB+fPfSaPVv
ADw8yOXo9VLiqWVghsvymAr7oKFTw/e/X2V1lFm8emlVwO2KgMPW4zi9/wiZaHcO
eQf8F4nZL0P7QCiyjeHYNQifaqdZ28gK9iL7ZyDnKQScyMLCkPsnzZq1t1ps2SGP
8ndtBDAXoh38KQCZAmW5nak76QqMZi0t6bvuLz9yHV6Tk+gvjEbHwNFYv8YcYL7N
43orugLPZhLFdM6RR7U3mA8o1VGfhygcWnbmt8ClPgN27imXuY2HEFZyGQzSOsTP
lMMYiy5d4DepJm38/GkxqgKCdKPH/B9cQRjCigSTYIz7MYWPda1XZhpS6oTyMet4
bTzxHpX3aezx4G8dP8dKiO+28wxkrVIy93nZ+MxqhuNTTqZXGZoCYPd1sbltRxfh
mv2kgoBE/1fU3NSVbSF+h7CF8cvzBYgRFK8uobqMRb6A3XohyJwIlmHa25mb8RGT
RCl1zL7VYQ/fRTDCwXY3R+WcZSCAWR1e59VN5rv9IxgSyWv+K85VjqKmZAfrBvDC
IMJyT2Sb6grtdOdzKxu3+6CzblqpKMU9aw/jR5b3pkezHxvUUNXbiCvj6ZxisXgO
jxSXQKOdEl7obPdY3Z4iadnG5N1G8Y5BR7j+coSzxs9p9PYQ2m6S8vHpXvyCiT+M
yFo9GgCj0Ujr6fiYI5RnYgeU4G926Dn27h8KGqvDU4KdrmxgqEiW6dg80AHzyJ4k
Xi6N75bUdMyJGxKlVRQFc2Zd9OLLehb4uGR8ZeZ213zMTzP9HZiugMcT+zONfkvv
BzwzYDVEeQaUL2T2gVc5dSbxD+Prxhmp873+GC7Jm7+rlQxO29qVSM764iMs1bow
XoOVQp8Z8TfsvbOEyRqI3423h4Y1s6TxqGfK7qRSzoq31f5FCAzO2bXbIfkG622N
4+LraFsRh+frMtVtuTbEnXTMmjYLu0sewYfW/6g3r8O273hF8W7xEHEv26qh8seG
wd46tsDahf5huFG2QzwL4l3Bb1PL0fjV4IplNdSLIDISSFnL7SJH/JC3ZdUHJfvU
hoOjwC48Xxk/E7Cl9vthrSaHB8lkAKYttY2TltCEjz2x5jhjcTGO8ien+SXYCFxt
iWshY/PmkOaZpBhEL/M2zxaWgN49sF70BqRVEU56tb01bN1+6VWuHNZls1knFA9F
2K4bgmdjWeY1f5HOxWxVgMEmcCvw7R8vXPJMtxoASIp269Nr6Pjdmi3at66apG4N
+pImwNdjX4NHMAByY8z6679r/36Lq8slXFHfk0WFSqfoeASRsrIWKOiK0OmAYWFM
qfWYSaH/p8SCyvx+YZB4u2Y4jJ+YmOpNEjDk1w1pyomWbMveoBD+LMGqEN1wHS5k
gCXE+UsL6tqV0xLuCLm5ZW6TYS4c7BvVndfVLweSX1dNry0x6tjip5VL21A4qmqj
HKbUsdV3JxsbQokooUDiHUU0pk6YwkJsBH+P3IkR7d1FvEQDxIhdxKENwQHoAzRR
J0Xmy1YouWXuVcT5gFkGH+EhTR7JeT6U0NeF3UQ+9lMHJbJfm+PDVEjMMjXjslaX
qsL7+2HwIejfl+v2NrhC2kGckmQGyzd4u671fwJT1xkZSqJiTOsHCMpg21xgfQ5t
GGzwkO8VOSsi/IDfyFZYX8T4S9od4JDz9RiHQbfrjrmWDA3aYuwViazUi9HJ4RzQ
ZglLX0KfngAFkMAwDuK2n4joJk0v3nnJimLqf4w27wplITnAHF/Xu4JiGJ3dKo1C
xkwe2PpUE3IFy++eJWW8Tzp87+1s8GDEZWrHqtaxbCHlfIyg0uj2sT2mA5V4DUFk
JK7g3SZaCNN9OGvVIu4r9LWwovLiP+5D54lBoR+cLi4emwokZ38sToreWm3Tilt1
r9vYkd6xrcV/sPk9TB6oskQjVw/UOFhp8g48nX2as7j39IZpgvFY0TrB5onMTsko
YcssD7orUk1RbTXXHxC674tVQYt0fy2sJfT5k7wCtqRYNgrEa2zy70m0QCv3gqCs
i/KNTvWGadHhlTX6+GznK3X1rSc2As6ldBnuNsDBn+TmIFRyET/djEk/UP8Pwi20
6juXtzM/bPxcHERQXwEDQjnitiD6Qq8aPOS/BKY2M+4fRf/gZuQDtBl0jT6MyII8
175aT4yFvOp2NgTBDeK0u+KPHoPMxmv7lJ/N8Vgq2fVsNVLOq8RWpKCS/cv4hkW2
5bHiXD6/ytEs40XqQb0753QQB4CNhU/ihyucIAY4Lhtc1J+5t/Fm1ZfWMLhX9kLt
CmotVNufJroWzdqZojZ1cHKOtCOyns6OjPnFSAOWMes+8BOqB6pN6HMfAcsyTu7y
vuPUGEkz2tQEpeNeco5po3+ugVfwGRXbVf+wzONysFOGBY05cSzzniWu3ka9f6aY
0pVgFgCbnikoAh4cn06bkyLsU0zBtoh/1yhNv4oNq2Uvcj3E2GTOOB9VlJBb6MUU
6sZdSG+4I9eo6sc6irHgiUUo66BwRbwMxn8wFUzs8F7c7o0j9mq95Z9niSgfWsPF
hyuKqLeAjzmMH7XsoW3KcxsN8+76I5tIhnEq1Rjmavibm/6tNWqsGF0gO+CP1cUw
PsxBx27wmAnbYreuCMLOgbyIaEidF2DJoYkKhLTDPo1Asjae4+zs/UkRQ5PzgXZS
aZVKrixae23FJBHAWpAEBWe9vVB8Eyk57yetWGAtJOD3yeqSTzN995IjTrrX6voT
wNmcspUsTerAoxBThoX+sRzMQB9j2WY7BRgbTa125VX5FwBiCEM8WeS5zD85BlAS
4/qR+nhfwPjzaZK/s3iE4xwdZtjNN7Gma485QbiSp05v1GOcYHGo7rxIedD7d5Fg
9H3jzFKc9tdM8ocCLt7CkLnimmboCBJIdD5vxCSEbLAdLR8nJ8arv/pfN1UzfWHc
AZm23YZNxtvkmsQcXR1TFhJnaXGSJc5kw2hZMp+Cj4iuV/+KJoUmqn3grwKBqBva
U7OHuo0lIy3Eh1Ih9oj8C+JSWjv01PIfmzAqS/Nu4jPV19hylosMX1rz5CxgR1Nr
LXHysJwb2NQl9jnW4KnKcEzKWtWiqxlLgDaoNRRe13ZFesmpVrKmNp5DQC5+mFO9
YDzr30ndh+uhNpdkis9ZkTvpBHZp4SAbMV1jMnSorKypw/wZH7lysk73QjEjonnl
xbZQn8g8R9kGlFyko7DUXylI9IJOOlwnn3kG77cyo0G8V713BbqYqgyk24hj0i6C
wfpbTcejwa0levNy7usIwN4y87ltBC2GHgyC2tuWb2j723MVSJxOw8aew9VLREi2
kIca/rk4LhMzEcl4Hb9zatqtBwoGuDhe/tFjn5X/2KaB7sReN99x2+zIyMMExBEy
btyrzEZp5rQCez+3KFd6eQKbq16GE3Zk7pI1hDCBBm3oarggyFGhHeHDWQ0kqIgk
mma2WSh16dVtX+YiWJ2ftvCgFkosyuQcdbqmi/xtSLPDZhKYOurmGMwNtwaH/Hen
pmxPFSHo7CLUduBZMg8TBeNz5lNzMYiESH5VTAun+Fd1uFVrvWBIRyw97laimLyQ
+AIWoebcUNUttBc2JcclBjvswt3rylvABwf966x1oX7Mtjp4eZPmn8AIz/+omrkW
nM0LU3oDEub0eXZSTcXyLvRT72sVda+PkIvbepavCajQCmHNFjfPewCws4CFa2hY
KI1tfmbflX8xwK7qd2+YqpspedJxbjVs291lRiGtVKW5lODNcIqdxzi7EhUIW4Wj
eZ0FkUVrstwgpNFbhoylaevGg1e9rOJZ4qwP+sBYZuDS9atpKAHxSGs9y3TkNPWj
pUuErkyPwpcWwwBUqzOsnjI4CSXktSMim5SiM31/o4N7t8Mg5ibdUnU+6om6wpQG
0YOIV3OMuqWLkTnR5U1EMlaVYz0xZ2QoQ6P6h5et+BuJyEgSwZn306VdNljvAWif
hznBAcSOWY77QEv07R6ohlEMLNuDMY3Yv82rufyFSYKh8wvsLWVTtc3wivmYy4YX
2ZRoFopBpMst7DywFgXNVAlOq+mNvBmLR20afLlPSyYVucjr+HinnZsWEQbn9KiL
64NzwDlISXQgpNoJtm3y5QF8GknUqDcslTp/mRls6jf71LZRxbOqnh4aV4JrlZnc
mUK1crRfEaK6hWRVOvXI9aRgWQ6y0gcqafO+Oc59zBfJpIUMfuRjjK4T4cRm5rbF
gWK8uNr7q/ZxLcsiyTCod0OyZlnbdyCpHoXP9lMvw3XFn7rhj0TyJ+qrAYQiUMer
FqVg/zlSWPYxtjv94QKqaNceLzsmZkDFTR9dL551FKsLPzKVJc0ADXTWl4dC0Mwd
BNvuAuBzxrVFGuJO+2yp8fgeXv/zFUCItdONu8z5s0MDihRyrcSXWO2mGgGVOfwr
mdr67ZE0aWy4UKUTzLACUCNkd1JBJEKCf92YSiKG7btJkt5DO+jr/RFXvkJIoMjq
TOS8Bsa0zGuK8CJ3L2kZECm3a/WMlwPwyPkUZgRr0OCwvz9k/8aq0ScEfhYHeUsB
lVJO17/i3zOGXKNqJWOrFx/T8IrQMiFWOx6s9awXzZPjmtq306cuUC26dBrVRjEO
5/5i7niCDB3VELvTcPcAXRHaqllBHnQBcQBoxCdwDsrMU/yTk9VXp4g9IYp5orH/
6lervKL68ZBAX9viMwnoSvaG3dsGKPDkwJebJ1i5/to24A7ODEaxingaKng9Twqi
9AlBnssx7bUyDGRQXvtGdkibN5G9DN69T0hj4FXwKToQAJaX19flZIa1kOxEY0Xe
m47FS/H//+RRghsdt3IBLlBEi0VolLZF95rVOj1PK79xIDapSlWzJM1LEGRGdnqd
tRMv6O+30Gi5+yKwLzxZS3lDTkHGX7V2h0RyrmyEPoVLAv2eRLOyYAoLbpmDleTU
8ah0V3czKu0y83InTKf+O55nb4eDUbEFtiz0wQ2Tcq2hvbL50N2m7I8Yxcg2l1MW
NrVHO0ZDMGFuEphA7500A9exDZpQfmKsV5B2lGaKX3Z0ZFGL4aaXmquGNy3fmHPG
gDqolYR58gh5PFaha1R/9mvCT3oet146MrMKsIDL1ECCt+21u5naYv2Bw80YOem+
Ebo/PO6ItLqmYOnzn7aAbXnSJN/XDH85YaFL0QomBjriCynoqhOEZ//2HZZNMoUD
BE3JaLRJ5/3/AJR/zOSC8OxFp10ZBX7Ni9w0K+dQIzp9tK7XWMbDmMV3lsvLofvr
9c/HuStR2KyBDiPyBJ0mn5jRHOsAh1S+8qDiqvs9LokR1dCbfM9RzhddxG89ohXu
XY5qssoyqWe5t6xm/GEhYXPsorx+v5TSkUWFIKNIwIVE79ACglK1ly5LjcKkONL1
4n5Orw0M873BbNOGu/c44lQhLpSdpRXiYFaVaLDMr7tOpfPNSaCceMMR+bjGb/Lj
HRqsnR7YR1QNPUSShYa4z+6XFxAZhB4wyXBIpXLIzVMTSKSxMVucTcOWxVPT1suT
/BaoXGjB4qT+C0PEh1PasPrwWeBaENu/dQipm8nkn4Mlin00gIhQtq5JjpVZGgyN
J6TL/DIHN/HbPlJX/1mBOBM+4QN+VTTQzxZISA27AUT8oAoxz7Zg2uVMyHP/fOFv
5lvxC4VzJPG2uip69EPR7KBigBy3S5IRCTnsIlfJN/+tpbkxZQ0FVSnerxMfIdZm
FnwY3gNZRkiuIIlcKmpXMwKUfUM/n4JJTaVB1Ba/L5d8f8EVLmEg5vFnn8hA4Mnm
5DjEMzqMmPUor3dY+2UKkvOtklts6+AVRLU5cFnFhWLf83j4q1TnqdoeVklHUomU
Qoq1Nbmz8SY2pR5HAWTmY01miZikwYGttoSwLeslomILYqKBQN/SFzbd1Vmr3+wt
xP/s3eUENiG0LXqDGLhmbgl5KbmzME2LUy17hXwNpBWblBDTF8WNo1KrptsqG9pa
OfttAHmLwpBeQIYwcDQrKfzPOWNnHBHvniBzjpnxjfUjgG3dRdtMtXqSdWxYRPzQ
04AIBkQcyXEXBrn8BSqiZUiY06GcKlctwwrSd2MPVoepxkSeVBFHmeqS0yFnkWFs
RICSvsIunY9GmkMdSpGBQ9JbzakMi9Rv6EWhgE2G3UTfxrRoTi6Bc44XYMcj9n9D
otW20pVABc7F7dZYh8xKZ8DsHimxRkARQZkY3FY+n3W1GJREstnHEl3xDWSQUU/7
IyVa/w08h5Aw9bwUVYongkM6QSpd0Sz6GVtj4MHuUqfbfOGuUy4+2ms15hpOLEOb
oWmlLPmy983aUUZiJfutWCDxMuuu8V1s9mLZ/JKepSClqV5LIGmw44V+CcBot45p
jbk2GsOGyQE8A6dhpzbWEVXhVQdEYdIxOh38wYx6mAJEA5pJUGmp4QIjjl7YDKZM
r7fZ6bUyoL9NFfCj0lNAFKcwTShhWb5ZNar/ktxEiZMV5mhXR6PyN5UI36ZHsUSl
Rf1oUdFWbNPhYLRSg+bODqx9S4SiRZ5KhyPAx51nWsHUih1ULRH+BlhRIh4pCoCV
PBCH0q+9IXY/uaIOJ9zlS222yeejBWoYSPbVIJHQTE7HzAIwSsgJopnWpXsqus6Z
WyqE4OGEZ+AcyiWDBZZ2BYYBC+zEhmQBCZeCTx4twlTd/9C1QUtKY8jTSJ9Jdezh
VdoofOUSEUpkgeqoAQ5jN6HSrzdiJPo3JMndHXIohU9vE/YoFeHXRyjyMxLWpATN
gSp3jKOZv9UamNKWLDU1buEr1WXNejUlEmzonvkAQ5UgG8A+6tjbpeedKbro7OxB
VG+3ALpfema0ay8Aus22KbbMZU82wo/HBUyGTd5sKmamzOvQUvog5ojLz62+oo5X
zJFYRI/5L3+f2ZzOrehTlEy8e3/0JUIhUT67y4qUniVJCgGg9vqMzk2N5NHGnBSE
NsDX1k4E3A0WTbWMKIKSpO20wy1ZkHT9+CugLBKxePVvjXxwl/Vx40ebTk+jrh9z
Ww6ZScKuNpde+8BVySzNFSX7S0pxrY5LP4En2eKBQyrqdFXErr22UKoPIn3fhH0p
mpRc7KgCZ5DUqnwe+83i//jAstrUjtZBfaW+jyzzYiowVA+fa1J6cgoJa0jD68LD
WaszzRfWagLWMOYp53EAuqzvRpTaNkkca1TrnwtQ8EZTf7z+qND8s1vxWNjqT6xG
+VqIQJv3LmuJ5n2J/bbad+DuwbFeKO/RHeQ91nT5sZxxhQ4S4dNf2GQqQH/gKwPh
ZMSjNfwPYX29x7Gmes1Tiwb2KAp79DCuacOK2rl8Ye0rCCmjXOUxYJhEtO/2PVMI
GLcgHahRRsx4B0U5/fek6XfbK3oSBTT7eVn52Ny20SpYYbienZoYd+hCmdvFyxk9
5g8NE5hRvLg4JSGnR6VXO8ZiJqbsvyj0RmSds6CclZY7QGP99HGLngUVD11yNy+r
GnjXR6oF7JQ/Cu+DGZAFX52LGXIj5Zd+SjofBtE6rrkTftdEcN2peL9WdIUWEWuG
xnzc9hI3k5ke2PXAjL01S3pCdWV09mX++Vy+q9QRRc5AjNs4tq0LfJMY1IDiPH3Z
0ZwNiBhF8OgQV1sxaYDO921Cq5cg0KcokJ7BVPAjOq71SErcINWcOwteogJJ41ga
aUZq6BrbIdvLxLpH+zc1N6yzxSEp5JNHaRmwwWNfQveu4GLYTZKStZhAGYy85kWf
nNJOwsd7p9+QM7nne55KaAA6avCYzHhS/NMrGT9Y1Ix9vKJQom4fP3L+hE4fPR+U
jC6Sre6rlO3Misp/cN9BfkWyOVImDvnMKtYwAPq9Rb1DRLAYhPJgFU99R8OuZHG8
HpJ9eWtvNx0cohc6f83sBEKPtFOGdvvrQymylMSwDbBsHGA883RN8e+1AAxtAI0V
sVKLxcxF8HRD0MZqyVvsn4biqWFqrfovz86n93k53hYFU/xCg5nMXy7BpGDI+wT+
QgLcfV94hOTAkHjnbBdKhKG8tQtazykPdcuFHGZwbguy1gxRv3qDq/ZGwxCVWXQu
Fm0rJqONaxNRfBGlxAbtL6CKUWiGzhuelZKhPSxCGGEeuUMGBugCWREQaQ/bD8Lu
Z3F+MWuWgj1jOUxCeB0B8/MUaUmNK0uUeQaJcnKvn7SP4qceIV43qwBH1lUgDZYT
8B3oikUYipzTvRT8o7JSXdLzX/LxGUGtyZBBnBFHrqud0SHzNSXpY1/nPzuLjmVC
N1cySnSBF9oXWmdNLoj54+hs2AFKEmtyFbitb4sztWiAOdVaYN0AfKPYt9AuO426
0AMsF2AtgT87QuaW2tcM4/taY3CRPhLMaNGLVsNdHBGMYvmUWbwI/u6N5kWUThbw
GM5a7yoI9cOtnsY9P2ND6Yo7J1+Iy+t7X6A4LiC7DOlD7l5R4jV1uBbLgsE+Pzyh
X28qZ5q8jb0YR9rq2AzOCaX4JxapF9+b2SSEXS1J3b3qRN49pKWmgfqcsw6AYQT1
qvjFsodawGb3PDqFSGSBE2pZrK//GjFJvjoKqHm9tvqe3vPSvc9mDiNFuiNCJoDm
IcuuDma9Mc6tyq0pEHi/K33X4wN5Gkb/5+I6RJzQwH0JUiOfCmWw/XhmAslCe4q7
E0frfDas//iYkPOsk2EPd3+e3E52UuO5X1UZ8woRwSYiDf5naAMy1Xsmb6zTfBIv
5GQpNtANkiVqPOzLVQ0TZ/icBwJB6tIOOxtTAEk7TggPzkGW3VDwLxCBIDsZQ60k
j7OmVyq66F6fXmqaCyRcSgi7w/wmY2cbIUJCdbfTikJobgj+bO3+d0LDMpBbgl6B
G7LLiFA+Mq2eVS6dh7D4QTd3oavteGpW6uW1swQKD2Ba0NcPSoRGLAFiMnGuG1Pv
tDDOYzSlaiVIsM7wT3aDA18AY1xoIyz25iWO67tGLPwMFc8VtXvPQ7h0U34n0ELp
kI3W6jyGXvt94bnuDKwhmrvHem9TWr7trigy8s52jS6kILWLtw2V+/78PMM6R4D0
PugXTI7O0t/ZW4iYGxT8pYnda1if3rSgJJpOjSyqdbyo59teiQHtz3wPNg/qfRch
fZkiYDx7CbAnXa2FPI7cOolIb93wK150AGlSRSPnd9cv/K1nlEkZ/0yhV80u4zP/
WMJyc9XoQaAXBm+UnmnqJ7Kk0kL6H7wfcMSHV4eTedrAJjvVuX4hoOkWGHvRALpc
cHVMJ0QutyS6MEZOU4jIr9tsCiqzDGGp3nWMbsGX7W0oOHO/zeStzJ1a8LHwLqjR
0ppIo5NFgKB/SqXCkWB8r68vS4LmncBRTMH0S4LSZjC+jDYakykFHTf750oId3he
1PGNbLN70sJrbb3hSdLhyIXgMk3Wvv5SnIY2SSgBbZKcKPkffRREmRvAgTa1xqZr
SK31gdVh52bY47je0QnVXyIxuDtaike9BFcR/uQuwr6NlX8pIhQq35/QwIFjTM9F
a5zSq/vUBZ46fC/J5FXpi1AFpVSJtvO5xODhKa7sgOUUjbVOb8N5Hy1yBeTp5STH
JbRNswMVNZmSDMK2OeBRLW+/pjWoCfeNgbTcvm6zsmRY7cQtnXBwDsqq/Fwpllob
IqVSAfSVUiGtBDL4Lyv15XP1IB+z9mrSU9mjcvUR48uIBFpMSHNXVPaCXthvD4SY
REaZDZcFkFQu4yMBP3hwSDcV3s48wIGxbmQ6KotvHGcl8hZQHrnQB81Obw2QxM7t
EPtgXsR6YfiimiLnrIz3vuV0GfPYg5WXAPdJ8ckAP94mInGGfnezo9kiTyTVY/Ao
WKdsmEzvej0roj3IZ8U3ltY6yG35FDoKvyRQncUTmyIN2U/2HbY40XRzaSkrnr+u
sQSgPjvytJmgkCucDLwaXk4rzwXNd3hhtLUrh02D435s0ERXyP9CHBOiSATE1CvM
efdMSnZjGmABDAoJ1GShYkspCqSNOo15IKKZ3dt26olRnbQE1QN3TroBSH4NY6Is
zpvlUvkR8ZcYMcaUrOx3PMRjRIITClOGiI0eKtOy3hlCRaEenvT9TEnevfOpkPmi
oEwGYfNR4ASen1JZ7k0ZyCE/g4SR+gm+szOdS76Rcu1SNOeyDgt88dFXmf/fsnhe
qCttfhIW7YEbfRCOuBnGUAqpABQJWQaOplnvPYsKTom4/oE4M/gBbpvbY97Q62Yn
o4qL1qqsI4WIaZvaha+3rC23RXFiFAmW1u70v5Q/tAvLmJEMfaXJqkjx8lKGwPqx
2NyEEH2T0C1Pq5OUsHJ7P5gPv0uoG/hqe9kFrYvr05O+LauEoOm1oMgot4G8slgg
EeHDqi7KMBA3NypWemeNk8dZJYoguiCx+RUHUlctMiXGXGX9nGvKap/fhONgJfAU
bKmZUCjGAIMQORSUGa6PRTSnkxESBFTsLvw9/0tZNbcXMNnbjBds5PJJRLah35D6
yKNWNLyEL9/9ygymwc+t2crJ7n+2qBhufzxH1MZDUW6PnFgfEKcZjjZr9aBBILwL
354C9Tiw4P+NPSnjQBTcXkr1Y+V0qyL3ic4FU4cTktUazXonMQ9fIX2LfYxgDpFo
ASTj2O0DKZ/D20RoKn1znlA9R7GGaQ7ILM8SiXInMlK8PVVERbwNGh0d4+Djz1o9
5c2baeRotICGP1SaEJxDQWvlr+bJoHflzknm5iODmiP1iu6ao8C+9uawXwLSEGIQ
7GlgxhI1OJVLZCXFSO6J3SleZeA5deb2ArUTEaV279x5E7WWKvNlhlqbuV6WIZVJ
xdSz6ULroi2O1zZMsQze5DgDPj0gIYnjU1gPkykcLF3VR2LFR9yR7nGY94mDqCFl
WvDxvY/wzqsjhSEaITwSWcL0o9610O5b33NxE+FzZx1DwWJGrUxyBUPoLMxT/va7
Zu7mBCUI74DG9AFiXgfuYCPSj/YCLvml0BWOWfOIvwEif7DOEa3ISBmi1k7e492a
aahTADdK3m1hwBvR11mK/0SRyaH2KISLhrYlB4TsLihpn9GDsrx2V3wvwRwf6blm
za2o7JNcRif6W16MZJqzEZCZrqqzlOXxK41FYvnKHzh7D2mJBbU6OMmY+zVhS76G
OpSLiOdXkgOpqnlVZHjdFVLt7LfFsny7syRsiWMrhgrp94xrWU+THPrGDO9JISDS
75gu8p1j7OViDfjh8PJ+W+aQ4tSD0XgL713lRwUiRmp1PTHcjVqXd/eBDBSC7zhI
aC28rBTfF4Sns1Xaf681Vs6vjHYKrBZj4AZNcpySyPj8gI1rBqMQAFW97nEWfwSF
PgVgC4DH8cFXvhwUwz8FlU66LJBoW64Ux6JKN7SIn+4hgI2dCuyfxyjwZUDTVZxZ
MB4pmyGoIh2UrnmdwKhALkC2AZFRbXFJYzdNue9XulO1zXQKAyrQtcu3kM9rJ43p
i1DTZg8JL3U4GxT18RUMYdnWDiPBMAeAQ2NIC7CjGr5o5bQdQZaFEw3gLMEBsPOJ
rA0wz51mGzJzTSXTM6fizdrrdP6hrIiNzPNAd4S6LuBEWohkVrav6+zWjfogyKuG
6EZYGP3XyEFSnYC88FN1yr0l3546IKOcXUVQDfjaTlHObCRZVR4bicPqajcINDv8
bAM48rO+PMA9yuW7uCwgiHMLyFqPabKwHapd5qGqlRuAj2PYsxIbqgQEOwSJTXxg
Iw5IBJlI1WhIxtmIAeKkJebei2KQuFpmmTpctKHrhI70ydrCYqtj3Qda83Eg9Hrx
UDEucGq1LR4EiJHdqpf5LkRSjIHhCLBDX8dV6tFnnr42uRSKGvxkolNBbirunL/D
7omi/7qQ1OBAGHwUjn094/umUiymwHBxCZuYk2nyOjpINFqxhDW9A2zuTyS0mqP3
BsKFn8RjKE1UQ7pQHx6iTiW7anSGmlmu8Ipfh/uUk5XboOlF2+RgRIjfh6x4eGC9
PHHshOoN7h8N5uiu09AJt8eBt3QlfcvmL9Zp8bjATHnCcoSZYsO8MpQlQC7Z+HZH
8TYwiCs9kKZbwobpfD63tzecFyQ1hFJPKqss4Q5fuNAb51Bo4B9gx/wXwDfaPqz2
XHosvQfJFo+x4BTfEieI/Ii/VQoZBH/UqBhBDsYyZO1Kn/GdczeD1k3unBIIY4nu
VtWZ05cSiRYvT1m6zDvF5cLNaRxjs5p2MGlrOcQtkQbiJ4bk9YRUUVazSuGkZkDA
LEXqgaHCY/xLUIxT4+L5s/3WGRP8rdwn4HeLsjlaGU02a6pyoFauHiogMTR043m0
+lxLE9UnUWccj5jbp1xLX/RcBufhK+5lHu9x8VTt6KWjBsKBG5BvnefrgKM/KJIZ
DRDm3ViYHcQouYOAhv+LmU2X5lNo01qIvllMV9ae+h+Dn5mQGVgy7XoDxOSDLPfz
E3yPLILNS1FHFeT/nDrQ/ETczlqhCvjvzvdzOQ0KYuz41rIY6i+Df8q+OR2H2Hr+
UsfLxxbb/25FecuR8oIEGhRNP20Yn9iZsfE3XTybwCH9p0ZaYGc9VaumEgu9cj5L
LNfYD20wnGota1r2PAf0k73g5584CD5LfQiXM5KxJxVdfyrxZy/GOYjaVGoEz3F/
XPubxjkl3U2PxOx7rI3wTZ+Vfh2DPSwCdYJii7tCa3B8cvEr/AdqPBIjrXyhq3Y4
Si8itkpGqJyup/if3sw7AqfUgmSXixxFPvSEorN7Z4W0B0V3M0+p5vgQHcf+ECGR
fQTxyV7vF4UN2wRNL3x9wC2HcJtTy9CDlIyKezy1DvEKz2uo5xC7gcQcMjJ+X6BP
UpqPIzKmtGXXyg4jFsyGeWmuBiK5UacYfFWG0aS5k6IRnelwRoeQIE02zRwz5YFm
Aqd/6sA04sgyC2E9m7HxBf1596lFP6C+9PUgbQne7rdCZmOf8EQ4rCwAs+EQxhC5
SnzQ05+I4wCvyigUjSZGrBysySlOqaBBtolx6xm1Qr/ODKxJtEJxnqCpfhEAGEp7
KvXmFoKuyG5djoW+7O11g/nd1kWuPGOTIfXWzbi09hhKO7m6e+fMegoepStvd0vC
LD3WQQf+K0GNgkf1lpUMc8Y7V4RAruZ9vUldTXBYVPGKhVRMrosfj++HzBxTLXBf
Q8WRsTgayDoGvnAoUxFlvR7irRcmu8pi+ACzp7C6WmiJHwZlRQLkwhzK1hjsHd9L
SfmUbbDOmzHsXSHXveIa+RTohgzKZX9fX/ubVpKpJ2vCRP+7QIRG962cJg4LhpcU
/U+tRyDeBeTEmogrgYYi59D+51YzUjUmUTKmzEEsdD8A8bw+E4fuKiAGDQHHGzVN
GSb8FAK4AaBzZWP4c5BLLEAtn9ljgNvkxVrh7oI7qpxXMtJGy+LTFzhnZ2BfVY4M
Ijosl4DU77Da12cTfOF7ion3hO9Kg6bomyO3pxHBsceSHasCJnzjrKqMOjwlm7Nx
e+YAj+uAeaix1rpxJHn5INeAFar4iMYK5Ey8rxiE7OtH723I1bGS+Ak2+GoI6Rdr
UYjyMehyHJpTchL2ZAb51+eEzUVC0XacHccl+KBk9o3toen/GIOJcQowGius85Zp
Syp3xQ+n+dDsyTAE9tmit+wmkaRY8xLETAmD/5ibFp5SeFs5DRDNieRTaM7lpSM4
NxoQGuYAGegMCaC1W7qQUygA/1aIjTbrpIUyUgBnL5fQz6UwAHqRoth9om1kwGQE
XsSbG9wyS9YQYhp4rInaVyvVpW+ik1vpHppVlP4+02yr/fRYtAvIsTD7gqRlkf8o
SeNoodi3ziTKP/aEyfIJ2gQRVDC1xjWmlRDlaiW1twfItKJOc9wDUSHACP6xt+6K
4qcHHsjUIXBufaXb4ak4QC8Qn568j5xL8xWLjJIM3FYeh+hEL6buJBxjxGKJISYh
3NmdogGHybt0MIOatnm13pUZfvjK0TNPgz3xClNdNKvNKdhc51iuLx3d2pzJJoHU
yvmr1h2BzJL19kyjgvKqQ3NWcpVzsBWV1Fgki6qF6FKiW6W0Lxjr9tjkwObuqTGB
zErMPCCzmnQxTCDhX/4opA0l50l7aTWtZKQMSEbmz+OlNBMFbkw36AnR15oB+eEw
t3TP7/0es6S8Sr5u33xdD1Kw4WoYZsdCdy+OP+cblDlFbrXpPfPBqlkPBYVQ921H
LcEoWJNAHu1o0GyCBUYwm76G/7QznLTly3G9Se/4OkvQ0nzDWBcJTlgGUp8nwN+A
r5GqmG84pku6Z25mtDDoa9eEfKJdFuRVR/O6vrbAzpwRXbvkGfwYvcpaypTqCCP5
JLUmiNJvPunRaYJaM4KpZPeupCW9wJLnM2Uxx7795r4P8YCUYsm0ozl3kpPcnEiT
ZIhgvOXeNr3Ro/qdFzx/8sfCXeKRsWi1OrmGqbI4OkxGlvxllhYk2QSmMags9KmP
7J6ggL29ZEa+wHRiemAE1tOLVIsREtyXS5NOyZhf+4rH5rifXbgDMZeucoqAd7+5
znqZ55WHkDrkrjhqfz7iGhv/odSFAklh/aGtlZVorkeDabPF1p67/JLmSQT/6Nyd
d6xi4A7R9/hABh+sgknEV/5B6GnMmAODwTvsh2gzDow/MBQM7wnGiE2BDyM/m33T
SzWm9hkiW3UAr6Mn7nccWrbD7VIWqjvPSLyS06nqCWdsvpdgUFG7k5rKADWhxYpK
Hah8ubN3hdJzX3dp/dGIuhPQDlWj4V1sCAMN3eGsBwBHP94hdrh9NxWE/TPYIRpw
60WaX/ghxayS08JOj4qsbVv/wiFYiu1pq/pFrSl9G62lj6usNP0xfCgk0fjLbnHn
PyTLB6R2X8FRe9JBs+I/UjZuj8cIwbLvn+H8LxsB6h/msw2PWqQUzOMf00846oBw
95AZTOmznJSAr+XaXW7cin2SEBHdPLBDUq5mGBRy2jSemGEjXIa+kj4+vZ34N0+N
1fDhfsCuKJv/u4qfiArVOdplzz8pDkiEg7yn32mWy8DFOjotM+Qj4CImemk89uwO
g1SeIz38iH8B2kCUs+zLlYVoJBWO/ov2qgUYqDDx67Qxp5MqdQSEc5kjOEjm6+NF
0LrYwO3+YrqpRSCvrCvV/T6XNJgBnzz5b+rbmoA4aANG+OwtgJXTasR2J4DvWfPZ
DLP1MSpyeu4pV5J7njV4MqmqcNwGbXWiRoXW6yjNINTlBgpryC1dVbgFDX3aijHk
KxkHz8boE2j/VOv4bzQplvT4WeY1/O93waYxeWLW4oG4wnTyHmgnt90Q/5XMMaa6
uYZswlWzTkv1Fc1jI/Ko0v8p2rQ3O4WWO6Ryf1ir0hGkizPTY54mqvsTk3Iq/8Xe
UJoo0CBI1jKQ4BXw2p4OsjOHyQ4E35FBscavqw5GUtfwn1MFAXcca7I0RfZ8VNF/
WcInlmo+OGx9oXHGB+FuWoPlrDtV4SH80A8J8p97JNc0q4HcEAirsiitz9LL/W0x
IBL88F9MEH9udjjxa17HTxBid307l42TRc0VEGOJq95yLjInHX7VVNau1X4cKPjC
4P0dvWe52yqk3jVTqpA7jH70bD6NhxOeEYweDrAJVq2tQbubzTMzusof96wK2uzv
uhSE4QA6Ot4TYMu2kIx3PI1Zqs7xK3OPeEIz/xZumsE1SccG+v5FnNeO76zHnqBj
DjJitezcMGuf6FUUzvI3S5m4W6FAt30pNKj6d9yfJQLd3Cy2AGoHC3Fh9bFu2qtq
pezF5/uXDSljDCfTkTq5VJLXfbFU/uU50tI1r/+kRP2J3iOXp2iV3a5lbKwhfwab
xjEJpEgXltG7/FBnQ0XkSQcqZtjlfasqpHKL80MBF+8u1d/ZydvZe8924RD6CX3W
krtNPQQnWi8GFTj3+iHyiIF6aPN10T7gl7gXq0qXQZXprQpU2KFvNUJ4Fn0Y5iNM
WIgGQhuYlFIlxr4osj+EgeKg37Bg1lIoIr8WL5d31LGIY11EGe1LlxlNA/g1bgeI
BPAsvYQc7asit1Nj/sPtXu2pi3LuR5DYUGpdJ7W3huonWp8b5Vji0SIfoZ/LRVK+
IgxBF4l+GFy5BKQ6+0Z7x28ApWHLvj5ZFS1UQ4XSKjEQH+L4kZYVQcchhav4lu/F
DdqvVm4m2Lzr+hneZvcm0ZpAd6YalhxCjUjz8R9VwGiQsyRwpGMAA+kC/dtrFgOW
j5FrqioVj+/v9x32Limi6tvb/BocNPhUgy4/ILmqZ3+xYvltODN4YeIShrETmyG4
l5Q1A/GW7dRFgxmMsCTrO6bgv0riN884GIsImjSgZpeJFlpQkU5GWSaLPr3z410J
YT0Oa7gqBKCHPBtKRVxCzGPSHdKZ5LPYoicSnMeDPMsALj2ZoGkQv2zl0rVnjXgC
I/dakQN4TnEV1D2diMa0P0uHwG9fqGA0C7S/+GeWFrTrFqQ8QANoPWCi7y1ZBT+R
beFAzGKrpA22twPPQdnrQso85036Tp79DnCnZ3j6SO0bsIAg9FOUY1uSd3PlJvUz
NBfo1QqgNIGj32/FY/M5n2S3sHZ+WQGWiEFLY4/htEqHChn5g0mDlm/htLzjTr0d
e9ggBinlrc0HnKEVHQx1tqQklUzVVMSLKI9ZvgykKPBD7bmv8iCiUyqNGlhvpN0j
UPfYKbqkq0WfIyybvxLKXxM/kAyWSKsILHnT2J5Pfeps31LAIAUImowZ9XixssJA
NNDX0H6vy8muxSiBrVV/22imnaId6UFNXeSjqpDbVuhWbf7Yo7yUQlyvAios5mXA
a8j3kxjWIRGzW+bjsrrF9rWnv4/8v+E3fe8tuIasXxcI6q5lq6HwQPQMZpkjD8Bf
ZUEjFZ6j2sZy95D0iBcV8617MfambYngQGrOXmGOYP6iCPEpVIh94IGu2VYHGlKP
mEiO9oiyCTH7xYIgrq+N28qHjQkTGKkq05t3qQexMdbg7Ge/kIsflqyjtpPBXM1z
nGfVAL/kdHmd6LSERqGnCZMAQFYODlfYfy9Tkwyfu51dynaanVhe7quzZWdL4B27
oSsp6nrTT1nVc/eSywmKMZlQ64VHkKeGwsR55Go8Koo2msCnH+JptAMIrhXGeLP5
ru9wEyz/j9f2Qcygdd5ILbwVywZUMwSTVrYHz75O7pOwaeKFm+LhOYkmQcuopdoM
O3n4rgYjeWKZCPoDQQcR8GXhzWmdeUkGuQ59Y4MrtqlUVktH62J/8HahnBOL6BBs
RZqADd714yBRZD8ChlecEPI20nB2M9Z0V1Bv0Ar1cBEQ1XhD63toUKtpG9P+RG2z
H+fROIJPIQZaqNngGkajDl9whjIcHBm04iFzOePKv117EnpX2o4Qzpx4SlI9RxVg
UKJzYr0GT9ziY8HLBQRKE2qgT1wwLTOql24W50QYYnHUFqWN+eabEcJh1w6Ieuoj
4jLwJLg37vQ274mJ/4PaMyeyrYsuel2vhV3BStVVuqYgW504BUc/YwxB2tGtODN/
WxzCI9GIeRLzc0GDSXvqEWwtHkrxR8YkNcHUISWcx7J3xsNRF0V3ekOOSKjrdkrh
VB3ucfFAIORIk2B4fSNrvElJA0Bmo+xH8lGdAck4r5yW5NUdZXz3h7S2MlbqzysD
/SDlL/qoAED9QL6iUZxNNNjuvdEy0Wfc8pre64uNOLTSwTWW0/MjdKaoeDFTgICT
YC9j9v8dUS6GwBrg6X5y1NVFICZDCMUf3ADp+LIpyXHsodE8Hzsc1ofJQ3QhDLoE
5FZnTsTwrB/+61zsB4cix3uEGpjWTTxWEW93UgV7kdYSh77dEUtgWNVnRXHQ8WrC
X3itFFOCLKFsnHtyuanDXfoOoZo+FQFM05BWSWaq8SDmYivifhwR1F37Yz5BQx1K
Z/uNLN4t4rWLhiBxiGDrhCuMdq8iOvfxLLhefW2LN8Y14L852nhaF9A5YTBsr2s2
UhCFWz6hZ7u1phgiA76QJWdabBONyrwV9W9CgncKNcD3O36o2rkyZoldyigpetI0
kptmvH7nUaTU1fv/EXiqBiZTDOK7G69QxKWIwKsqAwvUol9RgSFKAuDsNGinkmLZ
WQhdNd1A8hLLJ7JLw2vmLrZKpzz6YTKs3OmsKrzeIj1AHY95LuhwDp3btwYzHvUe
jtvmvmglBZCQOLkrJuFJ7BUr2QRQawwMwH/+Q72WrUmXwBWgoE7jGt4yr0oEh1GH
dm58SLiuOMgaqvEepc1cS48LFYP1spZXzOAQJMC1/TqcSVRc4SIxWR4d7Up4eX7d
RdsU4iJLkPpsvbnjDVXn4+epAKIMUWIjYkedTgrMpcT+Vs6GgdinUcy4oqcUIUqe
982tEQ9jxyXH4uWH4oOuA6osw4Za20io+ucC0R2+DsxI652hUbCrgoetV7xvAuXR
WjeNzX0VWztkaHlCfT77UM744zR2UmPVKR7Vxf9U4gdIH8/uCbgnKiHIcXHvRtvW
ptrfBJLp355Ky6FYxVf8HdKFaxDgThMIjqs6DBHwold/bKXYDiCKVUuEvDKFsZXk
lsmxHdMnPqVWvbnyqMg6ag9YnCP/1husgJp7ufDYdJQY3edcNAHFLFybyntR1jk9
HTFnEwTPOL8G/DNHXQol3RYd6PRB4X14Vny4Gm1XlEieugzkIBy++fyECW2viKUd
SKwwt6pZEcGxVMz68mSzVWIQWJCS7Xphph1XVEBzWvJPwNzspPteGDnLPQP3FkMr
k/mlGCHVkrrHrLk47VaXvppTm2v7PBywkGWdQIIl61erBBE5mOVAtFufT37w9ZVA
g9Zrb/PIOeZ7XRmTbzi5bZzez/U0kDstFxtZnkwCT8625gBNNjpp/rJ6ADhZT2Gv
zQBz6Paaf1Rd4O2eN/3npnECxiRCehRflpg895D5Fs/gmaWufIddE/A19mRS5HX4
6nTotBphE9gaSHomdRTI0xohDezrlW6UiBoip7Gp1YX7gN+1KI1mdGhINbLlbCr+
IbenfzpnHHVF6kp9qBtej6yg9ckcw1EP+18A7s7OTcDwfo9ui18fPDPntCfjQlPB
QPjG0bY2ul2kM4pj0hVr2VZU+Sb4K0/Lv/HajanjA/COh9mLwA8kh38mKPy9juSM
/iLjDhLfxzFd0zKJUravq0x313kclo32ACnWCmTFBZkrCY9y4wum9Thndg5Y1KOI
lfL9TCOPLFw2e5uyPAOzdR1n916ZKYpZqgANVFAkx9n+crXQQyvbP/AcwbS0Wrzi
T35JArEH/QU10BGqINmpGYAttS+wHdDxCryM0ilZxH8zrcHz2jsEOLfDTOpCYxhq
SuAB6tJr2Tpu+knWpDUUXNJivql2njzunZagLMz7DrsLSdjhuJurow51/Qkh8tVH
Rt/Yn5devhOVjx/uCTLjsz+WiCYoEf8nB9SVtWkWinfypVdbxZ9pjxdGcnj3Zn9m
yLKOYQa11TH7D+pnRRX60fTe8mqjwhYfiawlKgWohtv7gEqwiL3zqc1S6T1o/fa/
13tD63+mbIQnSG6fwrISdUng2w3Tamqyri/mE3DSJvMFqHnSb4YEc7J8Le8Enxc2
LCMgp7fr3AB9Rb9BcKQ7zMnQnqSqllm5nzH3bboL4Rgiu12BOJjiT4ehb/xSaB0d
DhHCwlcLHz/5ahIJqJEnDaPB05JKxx6tPHcdhH08QkyPaf1QshVXqz0OG54PqbC0
1VHqkEXirX086m7HBnOu+3KXyKFhs+FPIHm5Nn5RSI0ILfSmCuQcZeBeu7Lqz6ET
RNw/+NnLDu99vHkg8ZRpX44wlQhAgDg19HEvM7OA1qdBl8IMCtqUCB1C/sPnMtdC
TT9NMw/XHTpi0e1nmQTuATfEkfOdHeLlFaFLbRPtoVNkNdO9WNrkDLPS4mEfXieU
Wna7KurzvHZgwu+E7lP1n9J1kz/9ylbGuSXl1KL/tvIM+H1guUrQ1wD/jy4CSUL6
QVz8fVnYZao805DBBCS9alMfHFG6lOxLDKwvpS/3XO+wmM716vdufg/fzrk7naTx
1mSBeMHAd8IYsjdWvmY4L6zfwzsRrT9zzB7Gdc+0wjXnfouGTwjmiMdIHg/MbOdI
KUtadtfxqrBzWSbk8IoiSOGg9izhfnvN7bOUlrFD03D6d8TbpsUcvLjy21YJDOpG
c031Fs38MZt0DRtxVHaot4/3hIV9IjHNTsfysXofLjCcLXCevf2bmxQpMJ+en0JD
XL5uQz3D7DmfDNUV9YYX6ueZQJ8p116tztT4LaLHLjKz6NG9BLfoD9uKwensqvdh
LXpU7s/rjBSxWQVuRdoAmAqIX5nfHDB/9fBVPutsYv3SfkMdBx9dJ9U7Q1fTBusH
8cA/CR/dJXlEtNZkXZ22PW+oSsTlDBUkGh8w+MG3vffmmA0Q/048EPIhT6g3fn6w
arKKud49370b1VakFlrFW5o3VOK8NccjacVU9OxF5fq4WyJUq8PnVaZDDJv8mm9t
nUlS1jBp6trBFsjK+5dfOIA1+nQEIYM6bzwC+m7g8W46KEVD13ifeXW0TuZvIB+h
GNRm81Ef63SL9DHLWY6GWSINsYyZKDYE+3TuJG22jzTyxklj+ebkNMsHj+GkrYFY
YjUIipPWxyBScIO3gCxQatIl/8Em1prQwYxflyhDCRU+Tvmzlk5cqe1i8wK2DqjX
Yy3iAknYFiZ/fKRjF+VITT68aqEPYt17Ii5M/0Hnpxj3Z3UoRRu1LXQfBk+ymJCk
ucUIYNi8pBP121gDFlyYVT4GMqIL30JBg/ryRI3Y7QQLCb6FPtS+RYnB3UJNKEhY
1Y/xmxvGDHfczmhs6Ha4kPczwfMPRfSvETvv6IkHqgCM4ihnUpeLljcb4q6YEjR0
gbKq+JUigMveBHGbN/Ock1JsqD1r4pSg8n0U73/pKPoEKP6fA18ch5OgK6B/rnyv
KwUYywINwCnKM/BrlGJRD9ws8sF8UzWp+MApkuyZ4dxV+baeNYL4QWHmxop7fnBx
ESt3NoUqxiclIkwVYTJ9G8aWnrXlI0X8YSPkqj63W83QCPZte4ZpeYJeP90UhLSt
5KIn1kTjUGg3BERjUF8HEMcXJp212xR00wLJRuLvURnBc/f5RX2PrVaf+PK8dvId
sh9Ho1uC+DkqNRdYGdedAnJVXXEvnWXIcJ/33ekgXoaAABFWqJjLvEnYT/O9xP02
d+GgDozbBptU76qZC42mXqGb7ghkrYZeiB0NI8hk7gJFxpux/ZkbxJS6Rm/nGwup
9IS62tOW2dOO++JIHlPyh+/exyapmLzKd10i7cgTtIjSztWup3MOaRUYEfRlruld
aBRrhH18q4J9YeXKUJEcz0jzTIfStxA+NVwjFHImLOMLY3NPEy37HbTUo8p9w3n1
DGNRDzDF49teb1sadxyU0g8KvIv8/DxRnfvuVxCXB1kcMuyIoZ9fZT/IYtNCu2h+
abQ0FPK0y39OwcTv7h2UoF0EhMfTQu9JmL+/nhZJfsxq6NBKOT4WJ7T+Dd9VfCxw
5FuMRNtQbvbq6Xnr/DjU1sAG8RBBqQKcoCM7FZ/UDtoXIOb06xjwhWvrMUnRV72S
n5LQmn87zypE7FIfITmunRA5Dt8Bs0kZGtFEboynubI/064OvCvjpGFaJGNUhmlb
tXOo44nIKiTAG1SxV+icRxvxRyS8P4gomS+SNSTjZ3GJW8GqvvIUSmJYqHV4lw1r
3hxwt/L80BsaBqLR2Y0itBkWEZiZ8hGknwHV4py2lF/F6fntSOPZPXrFvC9Nro/E
VPr4ubPO7Z0E+hPFXnRe1LD6dli6LQLAqLk6pnAOHy/BXlYLluwznRJT+mQzwuiC
3Jb+Vcv+RV3h48vqxBcT5TX10tiryUtQO3hbIs2jww10gJM/2NYzUwzSjtba4VDK
Sl+lyBHO4gn+abhoMEp9OkBLy4uASkLojYZNRTjtaQGlDHWPslGdWljG+EdE5P3F
PqAQU2+A5eJMBxB/eaFiuQykMExrTJzeIfulqzR7V4Dv1PWZ7YghC8swd8Jb4gUI
W/HH+wiIVV4XukgjOFcWHmF6BmNHgRuA8n9a9rJj2JqBVr5o20cKuPhvSfTkfjWw
eVhZeBpqGBpGpFuYzYspFNRCsIXVH1FgKZswYLHq0J2mpeLN5kiACL0PD0MyTYLw
kbYjU6bWzUWlI3JD1M1RIlHDDkQWBUXjI4EB/PR6umTBgX/I8hd508VhS4neecQn
V1rvmX8huKfwHhAFTcyarTAAUy5/HoZhWadooTKRklFoKriesbvmmG5D1GQQrp58
YhF056ibUomD1ygS0HIrwyIWXVBTAfNBMlYIGh0g3ghbJI84xiy1M5Yn0RRp91hT
y50ekv7bJICufZbDLkjRBzNBV3+OdKUqw3FigiJv0h/CClH4THdSm0c7FRMwmlim
tr2LEvAV1uC0GQ5mR2CtSZh3vL3H6BXRoIF78dFSYcEkbDgMfpQk8NgsPR9ahcz/
ZvLXfDxPP1Crk+ICU2aKFbGbUkdiMfHZQID5vZyd4drdcLUOxc6Sc9+9B17BWsr5
TGVJAxAOYk0oVUsVyWJVFLUSOQ9LO/fWsuIaL+vljaGhz5Abh1xKl+u1+2GPrFTZ
5JZpG+aItLkhaYD1dq5GDMPqFecnJOFItJr2YU3M3lqLakOTWrwqaOmykBU7chZm
9wrIPmvyRlfziP6iZEabMLs9qLLDRw7ZvdiYo06hPVOkFMyNVDOS49duP0anI8Yi
UTc4naW8LjbstLHxFHpyvG0cOXUPP7IFl6Zyypgtl/jyw4MC/rhSrRSyBfcU5xFE
M9TvG3OepuvbejzC4fwbcCnBU607LYpFv7KNFx7fPGVp94KGWmzYJNSDVJmvYYRq
y8HMyC5eXRiSZfpeAt1566UTGY7iOiIOCgIHQED11K/Cw9cSs0Bq9bKjopubQC19
aNmKlM8P+LGBBfJOtCpvI9wg38OJQS+ANovChThNkWsBvq80jwyMnMnozCVF332A
bHu6iJyjz4jdfePh/NBa5K328wq1ULhFEK1UyK1f52vohpNArrtezEJxDuMi9yTV
8qlxZlDvF6bWjQcyJJdJOGqxtHkwlDC1EDxA1r9vjI/bupbFwoTuPovc1d+4HWMA
QhDyY47Lf7Ni1URT5VQa5tmCRIaJFxEQw06Vnp9EXlep58nzVFkQFFa4rlWmeJo3
flrfz6meqoJ/8Bm73M5ySc4XnI9tO1nwHuzD5sqeuizJ7C/IgNGOS8cAuiNSU2Nw
JUKwQWjcEgE+EZmqAZllDgB7FrHwZ0DN5YiNTc/UtWn73oG+jW0DsU7Gs8wNF0wn
QswMQlgVAtVfAyubhRZyM2FFUA+JxKC+Fx/ishYQwWb7ykpV+AnjjVG9DcCtrE/5
SLrqPXGAKIZk6rDceWArgPJ4IQVD1Qnh2HsJmZwkgj79KrbFYICUXSOnKZfbUoIp
H4S3HkapAkac/Im6jm68HpIo/dGUCE25XZp2FGBXtRI/aJDEuweqUkmCEOK9F7ZL
+z/pXByMBaBkfIY0Wm8o8ujwIUtqpnOr/8qiQ9M/YlQGhyDDJezsaABwuxATH89t
AFlKm6rQTGAKDVo7XKsgkYVHdN3zJm/A4atFbM3Nu6diKG5Owkm2zqyV34P4xrDh
n1cro0G+rUO/bLMSGEn9IEKS1Qk5Pl+MBmfXD2owgu/qV4Nr37TKp7jlb07sSNtq
qptjaIac7TOYSCT2L+w2apBBNpbJJaNGYgEqaSZtQAj0LkoyotRLJ7E/llAuyNF6
bcuY6cBQ1MQy+DNgI3F8Jwakgiig+QMuhehu7NqSi2lb7WPHKr8cwMavZAEVpbpt
vN88Ix7FaV32lSHv/7e+cq5rfngA/JeBXTHHYJMCpBy/BIKSsWbppRPk2kB04Hk6
Bpw5VehMfnWFq0BxxxZiGrQsDasBeRD7lOiRa3JGnLliLvhPyGjt1NQwF5rvIpET
VxICHksQHjNH7J9wTHHPlbkr899oGHalpr2gedzl23afPEAzQ9cgDlc/0db5BPei
oh1O9cUa6jWeZH8oBTanjNFtiF6zoakhyQDFgL653uXVAZ6W/iXZKRoCiMFTRLQ5
H5hzRriG96pNQzEL66Fyc6dgzoDXZO4/WEDpQbPg1z14cSY48OGBNNmd7GvSTq7v
5xvwSVXiuVY4IBZkpfR2KIHukWAw6IG1ivIg0o8v4HSGpgVFa79S8gtERKtUB2Mh
xP5teOkks6y2Z9/dCq3fYjftmIp99c0TYwg2wq7qFTuJc6p5/fJVIu9j4L7s1jFC
1kyrhtbDE8i8u2ygbHyCgze++Sjza+Ieff583+vYqeP0y/EGkx2/4kjJ5zY3JcKF
jwzzySqS78qk+WHpN/XDa1/5gkAHvXce0Rk5hZNdWVZ022aQ5oaK3mkIB7cGUifl
uY18SH2e6MwXppGju6HrRJSC4YGFDGZoVorbSkFCS6l73ZehrHiqXWlLN8sGwRZf
5h4t366OPC9gmNAQ1HE4OfRDX95QgpK76Mx/lF51SRbcyx7QIxQUq28edL75yjIt
VgbBioXPOJnz9SAFbYKf7eFSwo04WELBdalyr68acsF+bd85hU66HHUnsKmnZydT
vva6qT+QQy0gK6uICGJfih5HifrzUAGDsHB8qznq7usxu6UxDbrb1cJGIcG8IdSR
Hpt5cbZJFfqh7KmjMltVypn+vEAhHKnsPLdlisVDGqenhjD9tIXoqy4u2nGO3cgu
jP1T7xoyOROFRaE4PzXFhwxzT0BHfSX6AM4beepGq6WlPAiGCNBeEQkg06kdybsc
18MGwUjRwtE03Hz3oF8ScZ9aWVDPQcOX81FX4OZY0JdiIO04WvLv0iU8lalU7kPg
ujnII8CFvdh+jMXmo2FGnw5cYQK7PJYhw99gaFWz9DCpNHZXPwZeC3bzYjHzo3zt
iSrWA1/q2YF8OXKzstkL684iWN8RDhHOmOa+QYWzWD7hc9PZ2gc4uuxHOpugPztE
WDEPIyWnQFsH+g5mfu20kdVXiJyTaUSgg1cxzPJ+BSRD3Z9dRlrKL4MO+AayaTT9
MCm4ClUhL+7vnUBKyipNQ2n3rwJwcot/uX6mCzDhLO7gXIDziiO/jvWi8WgTHRZ+
O7inrs2xveZ5D54UxeJ1nyvnpgMjjzB/dZ9OO3vWMglENTdNInjmJra63BznkkTW
atXsgh1qcEZ4UyXW6rKsbsLZqExn0xHwvqUqlGf3tA8P4IRs7feSrNhshilmASzW
RKOrT/zmC760QvUi9fvUlyoZv+90nNVC32CnLEqG7/4BUC4iNnQE1SDp07tMbUoc
YQACac4Gus+K78xc0C2p63SFWbA6w07IccpjF3spDD94sWbRyFW8+Osfl8bILkV+
XXp6nYoqRf7SVAwg9UxZeJ3JUgnHt+P4fBT+DKAgLNDD1ssfdFdV+1I0z1MWBIAV
JP5flODO62jPXd1iEOpJd9bBCVP82SMaGDbvopR0a0Kv7CmaL/kBiIVt1UrcYUHA
tLqYuegiS74uv0qN/+hCtdRkzL6/IkDj1l9SqY3qOFCwmt0VLsGk37iRddg8LetR
kTzyaFOzawQQbHS+Kks6Igv5OCjhpaUQlaYs2lKiXF/Ke0R1rB9ulS95wcN/iDsd
FZrMSNAlXPuwlFYdO/g3IsgRf+GyDxmtu8cwOuB8Ndz1bxX/86prV9hNu+4Jg81H
TP4zWpP4vsajyd16kUnu3CuVBWL9W+Do8HWDGyDY9vSHZgkwoIVe3OIUxpsBdLg0
3wMoPbSdDK7xBCKjpXBe1ifdFzyBJl99ZAFoLFa45gSaUxNmZgfonOHSYhFy3L4R
+R9BKC1dEyVVMH4bwXmQk8QzGS8/0Na6k8J09HWNtHC/igX4w8Ajb9NWzwOaNldW
LQHZWMihbQJB1hfSI0glNv2EOzwZrQXCtTwaWPVniGVgzb8PhKW1t32jl6Zn3V9J
pEhGpbLdAomZA1d1EFebqUjuvC9XXrAFCK1Z/WgCXACyTZr0bRRv2yoZtYcp5CED
TpYfXHYUNeByv9UzFr5pooq8ZhZ2RS3bRg6oZcAgzBYeFKTl9VcnG+Quua9tQk41
owglfnvHdc8K4B6SYK+SdjAYmRkJy5ab8gdL5bM4LaTrcc5VS5tjhJHPnOlU5wmo
WDJSuGcYNmoQpApq4UW07G5O/0Sp5HIqWp9WfSEyEc2dTUAizWv3Oh4yW9EATSRp
XOIlPmmZVc+aFdPq8JolUJypoMmiVJgMMWLGi2PL2P3QO1lY27COUbivlPh2hbCp
wZMByu693SgOJwQ+MQ2g7QXRB34aN8djbqglnSBgxGGcem5bH15n/jE5xgxM7wps
hiE5Psos+t4bVaIKH8xz83VnIYPJfsaPqhsf3sL4sAgVBr6xulLAbUk3/FT09sET
Mj37uy+9zVlIKgrKDHS2KVIVFlz7/1mAUycX2R8L91zH1ORNuOix+RGQHiwA+Q3m
Sj50pMBCttAKxq+QtpWejoWjOX+2/cUD64ZVm4zz09YMrDpr3TDYdoCEgUxXyWTY
SjE5PtJ8JSxD2e6Sr728to45DRk4Ga0Th1Zn4w//kk2TytM9zjPiaBQsk/R+zOJG
LIPaSsxjhNl2UHqEVGkpkwZPmM88o/gG/dDYh9UTWmmJM5W2Y6N3Vfn+2u6TpvYS
4H3o19P9xzWvo5YaEsooX/fEVhF3Wy1eXw/tdukV/oLOR+sBU10iN2MpGxsNtjp8
M0zBClDW58Krr36NwYiKVK6BbjuQc7kPTO8AgLY20jcNlM6xogn9wUnfKBvU6ywO
k2sMOhemK3SF033gOcqfoZ4fx8ZH+QgdAbEffssblUJZgcyUPmJ9i+xfbupbBsQl
FmPTQbBURvtPlTmvtHAxMrbKtmfk9U/K7lLzBUFuMje0VaduGgzIQ4v6ImrnNNSn
FurNZKv1yFeXSNQ1sblQnoyjLwxqJCNAmrssz31TQUnKIXk90fEg+HwSe0jI2eiN
8GzBWw5fpicdztLIqczGOJtvyzVavjkvPgdqYiWwkdKZw8c740mVwOtrTamIPyMC
noDNMunSqgDrDxnngCClbCMzPp5XVWFR7NImPmr7bCoXCKA8vfdcsMeiXCXSEJWd
k2VjEWvELSeQpGQ8026yxfeWG/w2C46j1gb7V3ruZUy6UACwkVdVTRC6qPoV7Yid
e5GlBlmVKua1C8BYwWKBq5hEOP8VcITefXyAubWQlBFjUxNcQ4NNlFrzxH46xi8d
0wdjJlKRMjCcaEgis5IKAafxH54wmc0vH+p9Y3AXu//7LBNdbviV10sxHgoowRr6
rbsGn9iicP9ysXOp9vWpyfxSKu2wlmL6ffTLe2lN1Jh/LoBIjRMd0ITtdofAGR53
UCrsxg1RVRHYiTaanmo4tKpkghAf1/gCcPucrACkm0Ca7puXHT+HIkrXJ466dRlF
njMZAj+5LSfkH1KlC+10L4euPuZ65Z0Hp6z6wDck9b2sHyCRGXVfqAqQnGUHdn+h
c9LQBThlrSfe7XOZF5CwV8b31Zr68MoGuMOe3gMjEUoZMIbuOKupbxOSLZ+uwH9P
3+qozNGlcgGJUXtE26pLNNYhEfc2eGn/5Vumoa3Z7NPATty3eyJcbDLRoK+zaoSY
aPtkmdH40jXm3yn1O2syueGO+rtMKeOhj3BvYPaOdQIyJ9senAdnxyar/u+7CjVn
vEiiHmGf2BQ0UITOhyT0WdXsuZb5M9ao6IrOIMPjOzyJAFARHxb35Tu7P7HeZ4qK
d0XgDef8aoPuK5Lg15gAGad6QxmZ/8aETiAkqTbutcT1UPab7H9TzZSOpII/h/DN
BsaQFzJIEcz3gEv4psG6ioNuL5cLXqlbaF3jkmJhxsHwticJ538yXCqFPPZHmwCJ
Hq138rdQkLl2lfMVJJ6RlqhoV0uKQTnEABSyD7C8E2pSdK24/HoQJRKqmsIK23A/
2CXveZV02idrck99t5nGRXMEz5xS1cHZMMsCcYnQ0/u9uGyRTidUS8xAT5rjJCcW
UefM0OvbF80PdQ19zV86Pj+k8O5XEZv/UjlcHdzAsSlxncw8/TWnqdoI0YvGZVWV
MVEr0RQiIze0SJKzXDarmbgtHnUbTLK7AIG2c5NGS8MhddJB4dYwH/Y6zzhynDKj
YofMbYbHjgdxU87oxxqbwysAQP+GzneHuAfGBuMDDPzmZzZfx9ItRVTwJdj9Zk1N
39jAOTBxnAHFQ81yx3ieXJ7UvZ8LGRgdKOlG5ZWtSZ+g682gI/8FWYkBhj1jkDvq
Y7Bv2x5Jvse/W9nSn2VmBuoNFQqzcGdj/Ux8EepivqqVM+lNP3T4I+48DXRiS0IH
t4VC80VUQek0QVAe+PTc5+GdWuH/fLUaqkNEQ/gtXLk0w6I5iCwJc254xEnLMJIe
AaJgfl/rIaL7QujtGuXaYLCVnuvuBJ4vPF+YYY30iZlTv+8jv+72CHCDBw+Hw2B5
Kx8Kf6U70JEkIxDST3FK7raZLWHXlhPRQfHZXAfjw6KwGbDGR1Q8gJdmawIZLDS2
Zzjt6pnFe4MbVuEi02CrQhDV7hxxjiPibTJj5SIoXbRkcWRHYe7foFNlWaGXxsZO
230X4yeSj4WzJJuZ9zkduikYJg1ZBTSUaizRjgJh9ol7gBqlxd9TaviijmNktNOS
PC4pQBW9Cesyvp1Kny4OAXTQiII5pFLMRIdaKgIj76EFMgp8neWnSu3DdZlvkLZG
0st5JczR5Xqw6Wi7vHAT+08rPFnUU4IqFdZ1KJvgqG7AlYpQg9kEHeIXPRXcrB/G
I1IJkrYJcuzLB4NJuEcj2VX+m0o21qqcvhfvUjf2PT4sGxstDUnm/tXwpj9lLzDF
XEgRhWJ+msOubEsjA0zqkh6HQMS+8vgGaaPbMNkQS2DsU9sgGulfPbGlT5pU93kL
ggBlqeINHo7SIDPUn9jnDbPWB7X9Jezb5dF0YKAYNV5nrwDyZ2K8oLk4jX/LKgSE
WDPKS4aOQA1j+nK56abYgcpfCESugkbraHg5gLacTOZglo9yFQOGTjGxzsPV0wjo
OuEJrcIyC/UtZ6B4jXbZWKg9HycaxRswwtPi5r9PVrf5/RTCI654bgSnnGY4DT2W
MAxKjVetiNTk7P8uKee/ea99LuzlpsDYvJNWnAIXiR3tYBrG3qPZTJh/cpqC4HOo
YZ9DY2C72nMIxQom74XYgW7s9kWt9AfCV72BcOmNyTVg+eQQSPegiDRWiXQt9jrN
Vuqt5W45dlDemdKw0iz3WFGYS6wgzjLEHZEprl2xQsa5zPvc1tg1qEW09kQkws9i
mgCw2r8ufUkhnQkXblfYNO9pRodq9R1/dsmDb4eP9kkdAiyDt8Gs8JAAkVaUXrq0
Rn7Z5StiaXxI5Aa6EWMB4KDZOST2vPoLSLCwj1zHdmy5sToX78aBsGKo8xb2lDrl
spZjFV/bOGRTt0x8teDh6DgbWGWNczEZAM5VhjG+GCUTPdiH5GTA3UUPLa44SReP
scjGBWfHkAQXkxcLwzcldpHU6j0M/EKeipPEgcBD1joKezauCNaSdergE9Vbmrmc
iFUtwwS7Q6I7C3hGo2y4c8ayQzXGIW9BEX8qlRzRb6n0/6clBQhFL5DHS8wbIBRY
uUJ2EFoBfnvR3/Td2D3DozfxAngRrzLHOe4MNgOFVhBeCg1Xe44HMD69mqQoXqXI
UPn+8E020bGvgT3gIrFSTZJ2JwX/Fa73+tcHPFPJCFL1HCHhxDr8XyCF7Wyc8PlH
K9YqAfPEgL2xpS0025ULqf+XZT+POzyMm2Lpj/zDCB/UZnLzZYM3XLRiDCuP0p/f
bJnUH1NXY+SB3sCG/Ut1RAwY+GCEhoZrNdgJ6i5z7XHJ/aJnOI4rZGuaofDZBUWh
ByUbsmlnMFyF9+NgLhmGbxzy8jHpynhSyaH5hQ1BCtWaX6rZ9z5LcZwcfrxux4FG
D02pX6wyXxnMVOuJRMZtNWKflS24KpznPvl86AdmuVYRB/9EpahDR4m50Uq+0NMG
gh3m+mdlOqoHXAn3mntBtcVjFh2V8pqaMyLtZ9LsYApxKYf2v18VAZ5LcZPHxiuZ
HBcyimp1Q9TZ3N6jh1mWxmbvvnp+7+EpYoHqV2OlknhnFlXG0P4gOJSSg7sXXr+E
3PWahdcoqWFd5sDCBtneFON8NSlQeljAwxbtCCbRMt/CRrO90X3+v1JFRQ/4N/Ty
1hltakkXwmItbYgRkQUb0SuCxOrmFBbm+tsa7Zsy9noXWGiw1T36lOJUJ0RceXEq
nE/AXC2FO07miJ2XGA1gPlQwN8WuM/UHPB5yc5sU5tYlguFJusmk+oCzTosedzVO
j1YJFDTTdaTDVggrphgCtWbZaKg9PwFy6cij6xKLcVpJDkG/4Mf6ugUQVZtMQBaf
kqCsot7vDq4n5PKnPIulGA7AmbHMkk4UorGFkPTB/wn2oGGbvIVcFhLt3tF97AZa
G6ZFvKnwYO4mIxnOtGFDAL3qV+ug58vH9WbKQCK4c6l9A2hx83PBfZIidcOodHJD
YsXHpfphHLq+EOljcz14d6ly8lUvAwW9EgMI2FLnnDDKyGnBWaldz57BcEeR+XGW
gPHw/xzKeulhvX/ooH4xqqtwmM0QWRM3N5BYAvFattxmgg0NIAD7CFKz8ewXE4hr
WbtgIRmFqbtCVDLmWIBAk2MESEq6WT0dvh+ZNUwV1oCt6cvuLBQn4Mp7PNmbT6Pi
nV6lwhuzLtd5ThYf2Hm1IfZiPdgYBshsmoMzGUYNYiJWx39AI4ZsjropmnJZJXQB
A/xEab5TEVM4c9KCRJEa2Nc7usvAEePB70ktwBi4cmIi2Sf1dRlH8d7psSBcqlzx
CbakkvE+bHmwgCOv/R1n17sRmwYscvvpNS0Uc1Bu9Duxqkip2g7LuhVIZ14C/9aE
YWvlt6Hi2KJZQ7kSOQObUgxW3mwZO2Z5tewGtEK4rS7xAc4HKD56LI6WaC7PNQQI
Z0ce3zct+iLumQy9lRyYrZCt9pf3wtyVGralA200WFL1Nr4l4qrVL52t1t5eSEKN
MICHvqI8Q1vrkoLuiXgMcjZ6ij2jjUhRn11EWluzERSOYQw3ifwTfzuWZBVp5Qid
K4EoH+50lyJLzDYo70Ww0fp733iNomXzRZXdBgRF7x0dvfoxhIRLj/ImUGniLhtJ
1AyTGlxGYRZOXmRZRr5tWYXvXVM75QDUKIcqRdY6zZ8gZR2UzHFBZtETJ7ym45Da
ULAOBDSl2mXvZTXVhjGsfrNXqlm3xSNceIkB9Gs3+Ij48rdpS26bwVwt0nam4iow
tua8YuLGnEpwvKeK3ucekKFXq1NUXgKVuX5V0k4fL0Lj6n8mO6Oq9Iyip7HKk1Ur
ZcR6DcD7ZzU/2DeABz6JMZVtudo7BQUjadgfQoivCfIBNW1ZNwaCam5MPNSfiajR
uuXSB0GzEwjy/xKc9yeHXzAlrJNAYN9FygD0VB6oSjKtRB54IZo1Kba6ETX+13tN
GaVIBvM6XdkhildSe6C+BjHEJylLzrKyoG3GodxaD7sQotOFq+I4/BQpd0Gvv17I
73PHZPsDCz6d4BWjdabRJFHR1IvQq/KR+Gh/9taoWUEnp4xy9pnGUvuTl9H/S3PE
DluLvcouxd/ZiWaHkhyBtcFoh7f+xLcKdJXNg9L1WDchnO8Qzl+SawtzawZxAbmD
l7SrPQLnI+Sl3UtFoQI8VAWSkNJ7B+WmFev3p/cuLzyrZ2bfVgy3QZT84LAh4imC
fVBraqz5UZ72vd6uV0lV3TaOdDjjwO+a75HgEj38go4oqUmj6Pm/HmXnTuno0oXi
F/lg0GW4+XA3So2wRViVtkk2S94CO3YSSNUvyOts3pllWvuHF+7HHA7E1syUWcR6
SEaH+945gSH3HUSScZZqGdm/Y1nIC5jtF8rtaIIdHbFNxVnRFCLIRwD51dHXRvlW
PykytVgeUiukV/Yex+QCvYd4BN61MbAoqdoHEy2ySMIKNcsRTLsMzBtmshZIbDRX
vJW3DSXqItn56LKPLwOmvwoc6vnB2Dqtlb+kr58iFjxtAnhYaida39TmaPRgCRW8
VT+qpLNGxLyFq7NLYLVgppWRkW8g/WeYNP6MDNcKkvlkGxV5K36ujYnmKAposmu7
peCgyNGo4wya/sF3XOzSXKg3swTc2GJFFi0/eHfFuXTHpOHUrdXPp1FPfzHNpoox
J6bIDjy2V7rmVkgAaFHJOdD3RBLxikFAgGLd1pMQDXTrGzTSik3bKzOttnAn1RO4
uUzAGjcUG0LW/iGDySrFxFS6KSNyGixPDN4+66nMX5gcMne1Bp/mgmjeZ58USYqK
86KMVO6nBpsYMTqEGW6szHszHnAC+NT5LB+WDrHFM+KKdk5oMEAA8pgtILrRwAYs
l2p5c4iqevR0kCrKSX5wbDk8BNf+UI+3cYNRtaThVv9TOBCSOJxSOZ5Wk/0J0Gmx
rVc24zvSLQ/H5a48pSpaW3/c26jPhj+snmVP3bmSfW8BLFSVA9y9GLvfPi52QpVC
3yxKYhTRl4vw1DAkE3pTb43LZu5XZ4AusZ9RV6m2mFMDdPm3ZePAt2B09+TQpSpi
mxVQAbnVKTiFKXVyPYg9k6rXuYTXnzZhE2xUVLKkdXcpsSLrdYZlvlQAxjm/4XJ2
Oh+2+5GL3APvUGL9fubWSW358uYAAptrPsbpb1qTHaHU5US5pi8HD50jsDeVNc2g
OLSP/HtecyTNSNlWjD1ig1K4LpQ68V/+tFAMAn6HebiNUTsgRXVJocR4B/wIvkOy
LEYLYGG6t4SFACuEeIDy/jKWVWCLqgL/rRXouQCMsl9shMHFbt53l9MHYFynNg2X
LB1B8UVdxiEqGq7jfRq2kdmxDLRUsbClVOin1ejK/4hXSDVs1RSrQOIGL0dT3aXL
bZKkNro3+3Wc+c+vFugM71rJSVKDZGpmhxXgBbNGOVXhFsPKCZP1oY+R8/892Cqd
87/aj88hsGTnbXc5HHusQxUrRk9FEi6cs4nLaLKc+M29ohapvjRvNpKYtCCdd6Rj
NLdKY6lg0K9iBJukMPhBbV3Mt+ZtVnTReevhoqj+pyVvaAMJanYuXO/thyV5FgTU
mtbXs9vKjpvT0JSIdD7JRFWhPd1z8pMunMgLdMgAAxPWLVearkuJ2lYgpfygP7na
wvMIbycnQlnnmlNgiuhfq8a126DyCbyLg6Ui+ULyqvlmqmAAvMcehoOVrUtSNqIZ
jsWhoCqIHMQgIJOaAssNUdwQPmOi+FCyFvOK5hOafyDV6cdbV6C1hAnqWKxoFBxH
DoP7YhVmjgmmTGTi+7yCB/zZ1dVmAF3I0lDJgxJarP5AgEhauGLHygp4RpJkdOqD
fWG4semLtx+DZPF4o6H992NcCMs76PlqEc2lpexFvlv7hm7SJpYvZ8PX5W9zP+l2
NPaJRrL5t2R2ywE/AHgJQI7PA4PxnxLzlnH7zLS8BIJvZdJRVYoJ1Rq1hK3b3+aZ
8/OeCwbn5EBtZcvTQeP0JjsFCGrDh5s3a6YzqaitHM9YpvRGoXHFU7V6yzg9Q/Wj
HFAgdBNU2CCR9u9GidHEOXOYY2JXYwz/T79Xi0tT7PtljRpoOBLCSqLfX73mhwmc
iBAcgmWVfxv9ZcbsUooOye0flYZ/2PHdw1vtEuYy42kkWP8TPn5BMGxhyhYPcvNk
h+8dxh5nV2wAOHPIzoUsYMHjAOjCm+dLAhI3aE7DbfDsu1zwlHOqfDUIGMtk/5ta
4RpOVceS6Ano8irM8alVYwNdJwUimXFEveVom2rTTpm8nY9d0WyKVILCbBj9cOT9
sg6zYZ7a/g6zXOngB7j/97JbnZeE0F3igmF1FacLEvJKfNGguq/M6SkKmsYdXTVQ
WOYEPv3A7LbdFmuTd4SmL/fL90HBY3QOj5+wg+DmQmPxoQNto0dDb80aGDljBOR6
PSkdtol0P0/Surj9SzDHskEOATl5WImRD3u3zLKe+VrwYUEWqkqdmmGeuk+rHFsa
RvRRwvwMo6k+NM9cSib6tBygvryCwcnKZB1m6YR8yRUad/pFVPHrbjKrKdn4F8zy
uUAB/MHVPpOCuj46cd+PmzzXqa+QOA24RYQdWBa7vaqBcHzmLumo70k6EE32jAiu
wdtEPvje+n7QxA8rOTd3ZM4Q9SKvnLHZ9yl9et7ZmfHWMZNr5zTvOdUMB5sf4nO/
LNgOG4/1KjURg/hhRvJ3yVUV/ckOyvhXqn6BNVxOkFJBxxfdPM1XGe6O2+M1+Byu
J03xtgiVkLQWTecxrT3s7Miu5EfPXG8nTtqs3ZVf0kzhbFBocS1HunR0F2qJX1Wt
Uo8CUnCURg1z77BK5A/2+Fl2wOTyvZHjL9/ILrOUKdT4Gk5atoKC+PPpl+KbZp0l
f562L/oLLk5yJ7CF03ltrV9O5DqADA6Rk9Bcp1I4ztITBAdW/qcs03WcvSqlYoSO
UH4GBa3qvu29z5xgpvQCDBLx6HFCNiSXS77oOb216/BVNyexHlXNrHEdthWHlIMR
zk0zv42rTfI0VESADQlC9/08oVnESkfqc953uthhzlh4yi9N5p7M3lcUi1D0IFO0
MtCaKY+sLkTfonSFQZf/pU+K8IpDa14nqXQpwPZY+lasFpSb5dJj89XMce8qsQeg
AHqgV9+8QPFm9lzOouFBD1aH2R2+RBT1nXN0JKwf3Ku2s7gVpPXBKVQfU2qb0La5
FAv40juhm1O7UvAyk2+OS3gLFVXCDavHdAmgoF8IJ7hxxcJd+Y8wAGa92sZahP4u
xawgC9YTew/sXKaSt+gIqcN+ONIQ8mgD9F0MN6yBdAdGadXwy/xaNB2SLcSisV8M
patn2bDr4c25ISi3F+FGO4QsmWfp6IJVf0VVYZrLPzTSVidt1yIpY3oBRM2DQ2NS
N9PI8reaAd8xgCn1pIXzTxPMfRQSlMd9EtszsQ8tLUKlnR8CdXhS4+PzK9/xzFtr
G9iOQ0U2E1Mh8dSpP7aj2dvDb6M70O1f8sNtlFdT8ezUx3himEwNPdpftDw6aFAu
XLG99pSInilQrXzsqvuEY4CHRs09FiClMMbpvK2Jf8HtkLRBllx9ZGwSyq5oLBXF
rA9KWmzRzL0+nErEXpPov1DEp+ZSfpWSgAFzHvui+0x1ExSXQmEfy8+vcrSsHray
7yna3h74oo22q46YWwYwLWnoro0utf72ekqSPdwZmtfhgAnEvwDzy9NWJlY9Nj2s
j86lR9Yu/K9g40ny49+GNnwhvZDTB1N+I1vW5jveHP3byagFIu0MRnfdOYsQ3uHq
WjSrckSUdXCtOS0yH81YW4biLmbypgGa7f1TrvBQW3M0+fU8G6MgksHrCUGDh8Rl
KnllJY3tofwX9HIYsTMf330wv1q/YJdkhce/HVQXm7cLLhj7WF5ersoibfmWfcKJ
G7rIOWpaEDft7hKdMKtiryLcieh4Nb/Pmm8XwXtEI/aF7GnCNTrQYu8faGh9w67S
69k8gjuIpEEZwgheUSn45moBcBcIqTvfaE2iyxjIgjQifLsNKIdkpZJB2aoqbYDz
8RMfPvy3q/5iv7KuoDEPLre4JrmugOK5JTlGx0DBzuGLpU9yaX4wx/WmrXzBJe6G
xizbw1vWLTsYq1rRAvRwEKIrktb765p9zppVmokN/QGz+niAnzhFbaJ+ujqxOF0z
DRFygkq4cwCC1smzmKCvYl+63epafreJes4G7Msuxx34S/y5p38D+8+VXHbMjZza
TetQtC5nqwpYVFoDFnQkC3oX51o5F3Bp6QiQ9ePr2Q08fNEMKWBKP+tSqnfYxLF0
ylsbZCyfTQW71NP7JL1dSUuCRm96UGQcLBdOkm2Ad9p8beN8UUINar0o8nY3NS+O
by3wQiuTvdItvfWTswIk1uZNz9r6CDgion9c8vnguaGsE1GeRuSBRvJkVfRyaOLK
PMZyTCDoNEckgmiRO+R7Eg2A6syIrolWLnD7xl7s1mF/xNigWmH2DqgqWxLeLDwH
UTX23pjvbXRYHRISqM+BjIYY33Rqpe/0Psy09XAjTxbRjcJdKsPRLci2n5qNYlHw
LsFPrMD0ukAcnQ3sQPdxn0uJpen6NdHObF6wxrmYo339a1hLwCBNeFXzsUFX/EY8
iAaVYs6kkn7A3J/BAUA4bto7poXtdarvKTrMHPaXdY4oB0jdRxzAK6mtVK+niaEw
OcHj4kd6nFvAspwhDJ2cYBVMFmAkTZ7oMnE+RfR1w1yBvs/9xiqdkZznogAjnYmq
I7hGmXNdMavRukjmCW1dMsOyPmj+ec2V1jlSc9pHyMf/rDwSDsdckLwRoAvIjZLy
gavvsOrZsL/NW2qVkhfsLAGUikOiE5lDj5MTN9TrnR1hfq2uPUZV0MW5OAx4RfcP
XetuVnnR0HbQQYXD3eKUAJthO7oTjO1+I2GYr69OAy7BLA5yc+8hhBNJb5Um9R9C
fI0LI1Jmj8GtyRJ/Vhzx29XRC0ffgXLKQvvmc12M6XmMIf4ccZjppnWIxlMTYjiL
DXPeUZTRqcCkyLoxidZZyOtBCDoxpWtfs5Kq77LPGPtUatAeMWAAl6b7ZDPpflas
00n3Q3zJlqXxFcCcJVRpUkU0uCbsHU5Cko6/DtJnPj6oYxp0yOcnkH7HZu2jjF38
DM+5a7mSkUmprU8z77bPFhVpjTJDW9HJoOSVFIoKHojrWpy6ZYXNptivAWxzwvRZ
iDBZ/VXeR8r0Ep/wk69oSQHola2BCgZOMtM0fYp8Jp63etib6XbDocHkoqn20K+G
USSNWsjq0B1L0vpM6tJqYsnnxdjlX/c7fUssgwH2U6GrV2yW0cBbCxxX5Vh13Wqv
onJnc/zIi3rvgr+/RvJnKZEo9TJ5YzW3AKsmDHI/HbaHpKLOdb8tdQtXgPJbM0G4
Hh+dBrpXNxC38i4xbveL15wd0hrygWEZGfAc0oCm4OcZ+JPK9NnMTBwIil3heDbi
tzUBQHJ3Tkb8lOU/6NxuxXW8hdIFTUaqApArpnhdczPlHP60WjvSUVxErQhjGY12
zpSHl48GbXKFswZCOALD49xwVqaZZJjGbI41kU1jmeZct4SZYKHjBOzc8h31F0Dx
uNJ2mOEoHMK9yZHC2jGKGvlzKlnxXJI0LeoFGkJFvhLHa98LndWkevuww/9VmsDM
Wo3TffnubnQGHk0uGY8x3AoewLIyM6RaQtTlKa1HOmvIK6dr5XjwDCi7ftBkkC0P
mHl056ZPQrU2uYlmH2ttgtsUgVMLf467Nns0SghG789M8eX3uC9vyoLDGIvFlJE9
8FhIH6Vxjb9VyRVY7Z8Llx64p3aePJKKok2Vu7tNZGvQh2Hmv/shQHsMOnv5/5sw
tEWW+vWJSvHge4sV13tgdZ1nCo/Y15x4Q2RtQnF6z0M6nTSIiX26SALRWKZEnZoy
BwiKR0lAMW2V0V+xtWBOkXRmMGFAOIEhH0i0orqQn+hd9gjp4/sYwle9KVOuDFOs
34USrDkO0NcaVw8Du8NZsoEmqj5Q8Zm7Mx5EoMNPtwWxhWIiWZfTLr7kJ9FzE4OQ
eHTYTm2BRya5Pi+NfabOmMgEtrIcGCHueiNNinWiEjnYyC73clIpL1LRWKAqrjn0
jNAzkkflNrm/ou42PTGSziWLwmG12R47mE/AytrbtZJOI6Td7p8FwiNqFvl0pV5M
byuoOUoFW60J9Fpi/lASxHJVEQr8aHGsV9O86t9sJD+r2IVZf93IqZVr3zzcTNT1
07SnxlBhn4aGv3wD40FTytIZSW0ctlMgX+rVEcqPGFR/SRielmyQ3XTCUgEG6shJ
iVrFDqMg8BUUWp/365YyMIxhfDlwFeMIO7L6neqJJ2+O0Fqpdv6Bsc6IBoXHDEyy
RC8sGhAQcdqraNGAhx5V2H6fl+HfVTI+PalWXE73YQUle+xMWPlpjLykXT1a7yx4
uPfs+ZauhmCcJ9qN9G9BhtcblUrYbHOU4aXeyG/06jGeFW3DE2MgK9/PUorhy5xe
GUbWjsAvOl8/dEHaGYMogSG2hNG8xIwwrI3tNXH6OSvPryf8ORHpxO00o2IP/ntq
H5DxUfD/f8OQG8VM/1HY7FgVUy7ljRL4jkYjR3E+pS+vAEqAjAX9JI7WitjYX7eL
bhRqHlm42v06lHw5j8NM4KRuA+ILGQvXy/202zca9TThc2ZgJ1lfdaOGZiV2YR1g
ud/IHqGnpElaBKpTiyie/jyO+LADsW3K5dqeY6kjVx+W/NGmqX4FAnUcQuwL8gEA
M67+czvexWNaFUgLERYVDOFQw+tTZYCrX4wCVZ43DuaxRFm1ty98zmpaTRfviMPt
Rs15bNQH8UCp7V9r1ngh0Uq+XdTMDO+IFp/W1YD+q7qlT+qYPWx12crn3ooXC13a
6LBHW8YDa1X05C6OpP3p5p8lQuc8SgxTHlZ3mZSn7yxNPryOOY49Q0cBRv3uhtrc
xspIc8IFdjq6PGpcjgAKwtpkRNhEYneTlkJhUbAUobWZz9j9Sim3zdG75FIwyNkQ
rzfd0DZdmq6PDVj+3XdfdsOwyPf0Y6IHsrW0KpvMnG5fHbcEf4ChHBy8FBaz1kqD
D2MfBLYPI5o0FZGyiWMPmkbz1mLkKMbSnop0I2CWdQY/ORqRsaDOIM49q/xZEuEV
SKL4SXb1Ye091CULvHvYL+YHccPhibcLLCd0dPKfAqKGQYxJQpFYEV3Q+Mq7n24R
rJgZiejBH65D2+VIji4gzLN2n+eql16stZximcZQXdWA0JvxbKCpYs5g8rJi9q/T
QDLGiOh6xfWQ5uwVcVeeneiGxamTqDwL9+94TJzi5tERPfcsdhAozmaP9xlPekY0
co0A1q0tJSE9IkOh7HwyKzG56kju4AoWB33CNLbIu0qslIu1n2wu6UGATirscHYb
wmAKmv+gKvUTvXnBlUOIzaPMjotqzhvLAYGMbRoCUokfrFFK9T+fK0QaO1JpBKls
2uYCyHdk7l7p9JLEwIL0qpzVtM7jRakqhlW7YKhg76J/tCfx27uTDy8P3qyDobhR
abxDfnXRPVNI7en6Jb7ZPUYCIWeuFPtIzTEX16RLJM2ScEL3MxjlYqOaX3pBZ1Co
z2qtkT73bBGELTixi6j9vjxykMqBwDVo06fZu9jsToDpkHd/kBeCYbDHIQw7wcsP
AUinL7g/yR+vErnngkqN1E4tkFmwKH+oTPsMBAOtXJM+W0DyoMVwnikEAcUsUOcG
9/BRNCajBJ1/HW/+w9shL9RdTvSIc8gvPXa+sbveVFVvMBIBwpUyFF0JDZn6Md+H
FceU5p6HtpEPYLzTxry3DIIwrGkjpM4P7G4MdcvsA9Pr1wc30zf504VDbGFVNWrE
EeDQANM5c1jdtGnowKWnK0j898bc72CmRtPOjpQyP36GA6cbOUy5OlzoXODjhL9P
znZsdR4PwmdVxh5dBfcLzcN2zxWLGUGUNaFlIXDvCDIKT8KK5YoHEQIyU6MmGwx3
PTVJaQdGyRatJv3Q+J2OxvZtLuWfxo3JW1w2QHtZkQGkq7IYJKF6mxD/7zrkx+P5
27bhWIW7dV3lNzrefAmeL7+ol0Vt729yc4O0GmC3dBlyu52RNQ4UdUoK+GW5S4MI
tcUD0umSPK3rOARQCLeRUBgHKGqCARiQ6euc2dsvxv64u33H2bzAkwXxg97oGn9v
p+vo3X1tpNIVg333zIJkjiWUAP3MXypb2ji8/gkr75lKN65ahKFBAbZWK6JAOp+U
a1TLUtqjA+E7IkDwFoYpLkBT8mUhnOFN8dnkpgfcBQhK0E7OO7FBM6KuOP/hafy3
HmirmE85q+9DTpOH5QB8WMcd46rZfMkSsGjE0qJAfvu3fpwgxMJEd8NYFNFJmnHr
D8ZLa75g0vvHO30Pt6jHl2YaS3nTCdKOzcuOqhX3lMMXzh0cybZ3c05jKOFU56AQ
vs9jkjTspjuPOfzXzO8I2iWZkNOqKesneYZC4eLWhIlP8Unkx/EYHZS9A2aq+e2r
pESQ4jk/30SYIEMiAD6+VOpVlYjEEtvIRgjSqTm27UACUfuARnsnsNPY1p1B0455
8UZw/kmSMsPQ7YyuN03qrbY+L9VSw3Ka4QnbBJ3/dRnJVSZfgIV8kqLh//b8Q9LI
8W2xmvbPR7y3q63xsIoqnmbZQjVG4biUKKQGu60XJ7KNHpXjuVBguGuOW02ys/oa
E2FpXm1qyislGiDsAUTOi0W4wuZhKJpBO8ZFonixmREwPQa9fQCFIAZn7I2hav2+
vEDjmH2MAAKETOjh9sdNQmowHiJnCqxaxNoBYvcpZ27apte61OlirOyALDLxbuVN
mka7sK2coJmL2GKioBfQiQGEeWTq8zC4HOEoJbIX/7J/xV7uOF0VW1cJ4hWTnW4u
xeEr8XN7jg/cWXS1lmW/WKMn02AOQRfao3VLBK4sU2I+7nretpXNQX+/zVGemde8
IOAsuc7ZUmNN5ASLO2rjpb0dR3FxLo4MIffw5f6xpvS+FnSEo5sa0B2UPV8Peq1h
AlBWoxjh/W6JjrsWAbmnsCkdIXtFeLLhsL4YiQB/PLOiK97OmFa/Lcc0V2/w+KZm
JuDwLfFyIYg1hgfNGRmc+D5Vb/zSbaBLdUKG8Hv306LFmMwT8eP9HxhYoVnTwV6l
CA48iqc4TniOBw2T/nKB/JmLgYJ4KFy0CYEqVfUnSWMbigkjyJoT9o67fmjv3L6P
VI1Xy7EvXNP/OSS6FjrrvaUqvYuslRxRDyQ6WqTwmbgrkoVT++5TSS77llEPEpe8
DB5abYrVLvGMlWrbOy5YbiM8sYESjcJuifZVnieSORYQFgUsZc1z5U+hLqFAHvRQ
kGqSheKYPulfzYiAdnlyIBtAZd/lezx6lCTKYLdiwWYSO+fZ55izpa5syUOkyRAn
+7KRu6xTa2G2ErIA/rWkOdLzujl1HVLCHJoyGXueiD+1Cp58itnmADWzUXu1ZS/K
HFSPOUTTmW1VY1P/m1cyCEtJGT2yd9s7f6x/c/ouVgyjkNHtBRBBJiVCcdCjGyeJ
M+nVX3j0RrNNtYBI3LqZERQ0Nool+/KBJI3L3GH8sY84J5zzzQXzSrKCIEHgpmH4
mn3Rpo4fFsIEpdzTbO3IHzcGp2eOe/hF0V2pbmbspVPYP4+KbFknEUhwgFbyO8+d
y++89eXarAB1V3VcfzWcdMclLvJfINbvEJ/E0U3frEkxftGvbKSGIPRMdNyeM8Hn
IpT+4bsaOuYw9dS35dSPKQWtkYiL6XLTJwGZ/LQnAeaCstRI41kkE5fBWacAveKA
yKfhAqM/R/h/BdG51qrcRrjnXIHvjdy5h1ugMf44U23MdIhYvaMc8Wun9pA9KmI8
wCz0CdEsBVEQsKLd9wbhclo3F4d8zNxl4jU+9gFjnelI8zNj2Q9bkhG1w2/vI6dx
fFcqgrWSDVEEVE0/O+ex0WhJjJlTs8uiFQXuwFBWLja1iEQD8vU2zNtHf2u7IDlc
mCDNt7GpEP9PUGBfzgK6ihlTje5EKThPcmu6PUjB+ZRxkXUODO+fxc0XVFGN7sFF
We1S4wWyX0DQ3lzHn9M56aJtg5wjI1NB8HeGPvEZNToNkIRELevesJVAJRE+kukv
8N1w8J8auuL+IXMlpAvr8cTXvi17q6BjJ7DYlUsEhiF90l6emasaN66QiBLIkIwi
mocCKFVIdIzVQZoaeKDG4NORfYnAUaPlqfsKWssGWTzN+1NW4c0pMwq0Vi8Tuk6R
q5OqCAxMhNfGiyM3i7doo2Q6l+/4bJLMVvVTzf2XFOqggrENa9b8qQifzEG+TITS
KR+0u4aPJhSFNdh3qBp7nTt6O0g18t/QCjKt/ZgC6es44MMxlZQTULW1/pKRfwQb
CJUZ1iL3phs5gbGrJ38lQsGcW6PhfGKFsxEZqs4qyXZhSR74qzR5QVX8AZHm8oZ1
hKeLOX0EkvTkdRQpYPnaKR8hVF/uXK6apCqoqIxQJVE0hOJEz4tGXEIr6qrs42wq
QGW9WmvMc3cAnG6WtMTnamMCGuXorbp1gh4uMpumm9s7i7poiC6A+PbysXbAp7PO
1G2DwaYbDzrhMdqHW/7OgSdGo1MT+YcH5tngHe0lQdzX1uqbcfr9YhoCIwJtCrcs
ArVQU8Mw5H1tQxsocvTNIFoxsNsf9YGN77S4JXlsloKbMOFMNN+N7hEsj8t6fy6p
NQSixQVKVfZOW6CSihJ6dOoorJLXXkF68fcIfS+9Ge+npSBp0XtCj3I14pDnpjhn
yikvWtx1v8uHQieq62/4ebQr/iua7z+TPdxOcV2lTuu/rUOvM6jQT+tjjQwxPoJP
NDS5pWboEClvJBWm06EkNpc0qIHK3lNMdWHbdgctlz0erAa50CA3M3R6Y687LrF+
PfUynQ31CYkwCRbkxQKsk/JV6h9CDFGnPqgTG4HKBVx2V223UCZ+Jtae6haaP6T5
RHBcOYbDQR26wum1bglcdhB6xl6iBKR7mM3lhDeZX7VaaOHNwpHkzKrpnc4TlfNu
PmhdZvzy83jhQ85rQT3ODI7DRdvZK/8oLm6goVjffb9/PQEe9Wz8/k8UhLoop/zy
tiJNKB3es/IMnMpd2DPM4iOt29sHos/TxxXGmLj0WKdcl3An9IrW0tPpuhNXmnho
9Aakz7xY6hYe9whCzBx4ZIITUwZash+vktzxuGbzPFEkOPFfxq5hJs2eUjoi77+U
lotWZ02bOblYXALWN/p2kGC0zwg/Y5yUygRWfdXVWufug0YC7YBNmpnnfb2lUEWJ
R7SX0HiFvG7gm6xMihEmuUQvbsvO1ji6qMmp9z2Ub2C4emdMXUzh3jWU0D1P5SDO
kzcDqvIwjSzzyRuPTl4cPJ2UnGVgXy5e/zZRMewdyXcbdFyQb7rrHjUYz5oCrkPS
Ik0uIcqqX+2mWR2Ekzl8Y23tdaiQ3miF5AKuNvv2zNE6mZgB/XFRnCC6xyIjKA8a
jDRblPJHuDczQXRgZcrKP24SrX/bjK4YSbKPWXhfwzXyzuMEGLk8i6yl9tfG9ldH
7XG8F5G5qWHH9F5R/btcTCfqW2SRRAkARKrxCyfv219Hej+wFjuvfht0lP3LnYa0
UydZVvl4pN/SKoLAziweHaEDpm8EUuPECNl6xiRGsESSsexdrbIXwFTyKrdy6D2V
pIYBTKC7Zt0BnB0kfOZPQ4MwSnrnNJAXo+ZV8iVaAJ1jvo0BCq9jkcQPhFtftKNL
/L+mOUFd8xzpX6NtsgdOpy0kV1xMQgd9t58nfeGBU5yZjTQgPqP7wmCTsn+j93gH
GkwULCszUt7VEuG2Ar2kAmHNMFUXt9i0cfuqFZ7J8sZGWDksxuKNPk1ToQblBk65
ggysIraK+5o91WPrwqTZEtzzpONILIF8wbR40X/voaEnnpM0SZio4YWsuKT4cQl2
aiq1pSeyxTa3dLCKqDBjQTPZh09b/JVMXaiQEFxcs0o+9U9zkMEZyLmV/0NDNQ2u
M5EHJX+W0DkfJ3Lw2MkamV5MtXFZZhp3i4Yskiy/1sQ+gyxTIHOpJqDnTMKMgjI7
OHeyeqmwR4LFoSiMXYMkL0wRBD/JY0l+CpW1DTXBJtS50qgkwJwZCpJScgC/XYgD
gTZtsYu3zUJOR7D4z4v7LYgYfkxi7B/vjZPyNKkYt9Ty3niJuybkrqNeBL+CDTam
P1pKjajrOOElWo526tcmDxijkJDb36G7EeL3SY5+AnA787Nfe3oP3hLc0Ac/HcHj
M5HyPWbI0birsvRY4RPo+cLURDirOa55smUuUlbM6A+6tlE1XiARnpm8aapbZ8OR
NrzsTMrHy3q1RzhFMnA+RTNPpGVZj0iJB29BcTN3/SA00GjYTNmzQVeIjFghczfA
sbkyuSXUvR3HU0XaS4L1TrtBeG+is8bh9zlN8/m2klYXpUZXJB+q+iGxJ7kCYAPF
89ECFH7kAtQf3X3mBOg4DGOjGKEvH4XH/oxOvTusPUzCYDgQ/JKU7w+ss6RMcLhy
mZ3z+IyhgF1eB9kVy7JuNtkbX5OCHP1DcGeE1lWPHHUMSqKIzE3X1K8Uu4rVQoCX
5yVg7GBW2X+xNp3KE/pcz1HTOKnWzQKVNgyv9UDgc2MOzoQAEkeG7WDGKXoC/GDT
he8B1eVhQuPgrNVRKmAeoZ0KSYBk2DdAbJ93YbvQBpbP2rNpPm87eKjqzVZC8uWu
lao/zXG6tXdZejIrjK2oo1tjGLahhxC6T3zWYTCm/pC2gYo+MvYIjlFvNYQz9RFb
j73e6c3r0oGaryx5WCDDmrwl7v/LrLUN5ERR2aLASdg5UJMPdC/CRTOzQwE7qFe/
D0F31qX+IQYoMufC8ncs3tbXroxRqs+ZdskH9EDMN6QGQfRUMr89+/HPNkqlUBLL
eCM3b3TXKT9FZW2+vXtdR6kxxGc8FDvPWKVlTEJUzvBb1+LEs2qXUYOcwNraZZec
HPkhwHY4QPBSrl4Lg0zP8otAvK37ThvIbft5ByQc6G2nlRc8lM+zgFEkQ77tFlX4
oVX7Jusw5oWUbcRE1UZjDq60MQfZTXb9yHXNZ205Mkauywk9spIiEXitlHE5LU0p
1kGtrWg1iRQC8hkqAOMgJhRxEGquP/Mg2jMQRTEYgAHHtnntMLKI5w4FwvbjsnwP
OI7J/MpAM8ceMFsZXPcAVNSZrLynwZrtN0+ZFs1xSKdGLKIjGRXESaJhl2FAouEJ
Wkjc/Gp1+O0lxW9r7PL+oTANsp3mdeVJllal+a4WjZjEAXOyoJrMnzRIh7qGf5zZ
iPvikPavtbsyKTIYFNWEFdsvAZjbEn0N+TYaaYtHrG3DqSS/wc61TMZhQrcCQboO
cxSqfokJIvHn4DwyrXHfQABsHpLRErp787yWiB1oxLgmaA2bYaC0pao3RGlhFPy9
nebyLwwlM1gBDT19WkfFBE7jWQRHM3+/d99N/oH7yAnBO7i34CeGZrH9iRbSgfx/
s186suxWVL/Uz0fRyM4l7YwmbvM8Dq8Xs57nYXAKrh6g/4P2hjqiDGB+A8zZzhT0
EH97rUZtvpwJ/JrXkXmjJWfOX4nGIDAm5wHuJqquD8S5h3CsKNuHeT2RF39xL++e
SG9wElNbxTfeQw6ceK584Nr7VzpIlOuGzhVVzry5bZ2KfKwcz+kzOswZD+ILrdIs
dGjwJy0YFX+jnobPfa0lb0h/8cFk8ai1VuATsnxZEyidNr1Ig1InM7zID+KLWh2p
CzCiofkyNC06ujpY4X5if590679lsYtZrqDdZRUXRBlU8QRoVloGceSByE80Y5bM
tlAbCzJ1rAlsNVhDBU9ii9mWbWPGYpJzdXLGM/bAK+WJyZkVGPDiFmGFD8h/GQJt
pEKZ1qIb1D8mRrec4kUrbCGPQgLFfl0Ow2bKZyf/4iZTYBABxMz5j+53LKx3zw5A
oAaoM1BfHLv5DUsQTm80td82PZR7NWbaf1k3opq0jIUKDsZOm/owwAI9ZeLUQto2
M19c9wXB0J79qlMhOVgwglf1ItKOx8y0N9cwazQFbb1DqewwNnsMxp/UY1qRhBLZ
8AtiaBHFRN7BjDnbpr5MGU6hvlTc09AAtN2hZ3rs1xawNPy/KuL5nONc6haF+WAS
mvHjaZvNf0OyocTXZwxe8hoMIrWcNHDj54FT2AtBPpZvhpeAU7SH6hkdcHLoBZNY
z2Uja/beD74A081C6VngliQRbVoQnHLz6YiJ1h5mc+JcElIW9bd2pqefVfe/qvHa
CgNnIyODLzXVZ2LqNLajCtE9YimFOxcqqbh8D61LtRzgFbSKHvodyxa81pT467oc
v20aP8BQb/YzlwweBJsbAcDyE9u2p4Y0k0810bvbHR+DcuSW60Z8n4oRmTjmiAp+
yxXjKpuZNc8BaWXzGf3qGMcAmpgi+O+x8xsP38OchXbVb4b/aKmAEzVNrUCC5t+m
fCDeG+RTbyZNkWMIru2zkLi2+I7gTYeCXwWGv9ed5YIi3m4bY7OJHFXedhtM685i
eLWxyYYWRyyqnba3L1aR4yJGWJn62ncRqvZsHGF8EirF65Cq3HNbxGX9u4BMYp5c
/EBC9MtWcsvaL6pS+5k/W6uuHaa98gSy086fWN0xsxRR1w4DURNkiZp6QCvp+tSA
v+Uk83DHo2+g/ne3qXmIjkr/Dkz1/raxEaMAu+RrRV6MEiser0aFATN3gzpLD6Pp
H5ipbrFpjlXR+geGzJMd2UVvH1rMzfh68PzuwFm/5gCzPCrr5Z4zMVQzIDQtCRho
1XuyuxLm9cuN09yItwalPmvlHxJTRM0Ja+9ZLSEMdJ4McQPoMQKjJ5i4j+KO+/Yp
yTEzG+VVU3mwmjZqnFyKHlcjaVcjA2YUPnLGGTB2WfF9l/LdQtInttHCjaNjOenw
mRgUMl/iX8A+neYI1pQNUuLlVt9Cmqka8mzaeXSs0FGQnv2++WLn/HA4xl+ugIi2
8kpgeezb5tsY+R7vYTjG7sAtSU1w43K9LTqHox/EgujAHXB1yGVmAuyW1AXQucV9
9Fjc1TQ4f++K3eb+CE+CXV+pCvqHkhpmJva8PzrpsIhCigj8q729uLKYJLjP+8gy
LjBVXPlL6sehVb6yzPQtgRkTTyRHn/cyuFEwyb0w54YTzAoAjmi+h+JZnrfYFlTg
NzublW+EYQYp4CVsF4dkHmapRsKXBd400g2j0RWgMkKt0dmzSKwf+UMkQ6ifl5R0
CobcWcp8uvYyhxK6JSNW7dmGkBnjeh4zXv6FOZj1A3vH+GS8j+yV1hRvHp8rZ39v
WKVv1XNEYlNCKvS8F+IPA6bHHwPUKqI5qIrG7WSXxPTiRVWg4qOXpp/UPbf8SsOX
+psjF1iNfSjqCYrJE6BK2bHGkhXoCI4gk8C4O948o9SzX2RRUNib4NPDT/a+ch4d
Lh6YEXtylUfy8zlHVOKgs0wjoU3mQZ+KvCvNVuufdziNgjYDEGegibAXQdb/J8w4
KyrsJ8+pErJka5/9AKolovf8Wao48bmfQurgmViGKSX11Sp2+lwpcdBk7ap1yHqo
fz7S/XVcuxDwdlGNJdAi2g0JRH65DOMmXT1yJ7l2FShpZV7oP6QsuOgmnk1rdmpp
49csKyXEn44oeLQmq1jcfh66QuITZBx1f8aw00cghF1rZOg86SXqD5STyMi7701G
tncv4oWrSoVXa9U99TiJHt8kbv5MKMGJ7Ire0WRjVpsDGKTfAMW21r2Ebkf+kkCU
q5QcSQHH9BLWajKQE79hK5EXSUBABWzUdOO5aKpV2+u1A/8DAFhkQHNODDOquhai
3yqmJKCgnu/ZoWKsGdCWlM8s80SOrGgcGOXXzYhR2bcREkvFTExspxBXH4ycUqgo
4LjBBYlh55f3s3lniuqWbJ2IQXSCi1Cd9mnUUh1/TySsJI1xscFzfAdO021OArrO
H3buzPIIUiH30acm3lNLJG1uZlyyIPaqJIGQD+BY6G0ORGOBmqiZukJ26/VNNWxk
sXhGfSw4rfwAjj86j0VFSiEJDt+3zPCLAGMh2n/g+H3X+KxD2fhgNeYhkYYi3xH0
Lf9Ae6nIy9EC9HayxH18y9q7OMoDE0kfiZkdG4tn/1xYVn4yv6Cw8dwmHpHPKGyr
PCTOy14rGrXp53FmC672VVhxNI1hrR5S50y93xU2fx0OIkPi720oU1xyhTI2GIii
+Tzp2xklmgGaWIveqUDacTg1EZUwIVURmaAH6AQ9GnOYpjuJcL5NGyDjtQeylpPl
06zdVnV0xVfuqFXsVjHLGp7UXziZUJip0wyWuW27ol8kB0n7r8O2YzgI5BbONyL3
vZehIoOKvd7CtY6p/OVoZj63y+cTBQvRJVjYzL8TuRjIKWU5S9Yge/sPMNDkLiE3
iuhP97+TacjrRAF5HigijZHyKyBeNeOel7nN082gyA3CF2ME8ToWY/tkG0FOQn+3
Noih2ycGFRBezPiopCdpHiiAOsmMVCjztV+jq2wD27kEjk+9kMzUeFcisrBrGnrL
Wo3TF7ug0yJpibxlIx4nGkd3m1eBbFIIgKsvXWrT6++DNFDq33pWWxgPYk3Qq+0P
DFDI4oQB3CrC8G6GTdCkD+ccnx0AvS4/+5hPLzdGeBy339AfyiIR/whctjN7otS0
l89tMU/397XyZuvj7FB2ArtUZr/7lbBhAN1g1bdEKXRuwa2KfbTGih84SLm+gzNr
sGK0QkxpTgdlmy+h800/Uz4+Lv4pYTrF9Q6Usl55tZEL8305qoHp52TruebUBtck
j5zaCmlx2oB6CIONuaJ4KEZ7GofJhtWDoB78rCt2LqEjlZAM25na57xsTwNvdD3p
hYvjttzaIAAh5/i4m2DFcWApOLRAdzgmp/zJGAzO00d4FlQsfAhOv0HS2nCAl30u
62UNYXV6INfvnrF4LKUcB/shklMnetb2Qap7BVUo08MiMQ2x7c3ZpJeui0W9AG2e
gVs5XxwZhmeuztdwZbhqMb39x5xYQEYu0boZRlTSm0tx0BcIyW+bDbkYF23B5/vY
xiNh7JdUhJCku5kKRQCIK25ewLAEV7HIQj5nmsfgVDo4mMSlaQ8g4rT/4qV9l6hY
jdL+P4R3Vdm8fxQv+wNuEKLxStuMH4CRj7Y/RRYp4Bb2i9rHfQB4BJAYSfD8VVbL
FUVM1X9nwiUePQY86mw8DeDG7DtUuZJc54zXzkBimedk3LIGZxBfOKjbDMDvRvnB
zFwdmHhzH18y7KTJxhwHAwmRCAWX3o/2DX6prSRghTD4JwUdfwjc3hBEuIjEXs9R
0rEdaej0Ioc8vKy65BSDdtTYP3yxsyQcXD0xNsZzBOA38SAwCvDVOcFHF69/08LW
VmuaHjT3K8qLfKrkDKFDTcfGSNsBKGoPafEF1SNzr3dnyf7WdNVHGzgeIS1t0Tfu
B9mIs0WDsLcKeQATCV9g3SUgdC+K/B43BeNzV2gg5sWm0uYYTNKwoFgqeV0uTUft
k6m1SjcZnnihsxPwZzbpf6njqxr7v9fxToBKQAVBOxZVCGJ9gTbwzdbyKZRsc81G
4wn0HjDMW6qoW3T9UusqaEYUOrCJLD1Wmu0zdwDRwZmDPVS+VfrWT2AD1i+cS6op
ZPglRj+iGXu66YaAXMylBG+nGDhhRD0/G6PMcp6jaKq25VaWtXFxhLpvs7N9lLan
r9RSixKmFc7YT6/Ggy5GIFAxVUtYvfvol18ckxSJcZKFSlCTk/NlBAFRdIB8yFOI
iXsjRFhCn+Zbqq+6N9MVYJGVYoTTmBaIuh/8CSdwuByQVoqZags5h2U8g18TTpoO
J16rBhoMQmPNPamnHP164tLrCh05M8SEOHHEoWhE1nwkr8OvE9K8J7kAu9cvP6co
LIMkZ5wO9XrhHyZqDUhAGDOBisZnZi9b5XEJ03cuzrrQbRLSkALEit2D3O5mpSWW
OwlSMbwfOMzi9gGIDmq78nCF7nhtmn98SkR0purdrbD1FdJQL9Yctck40U4bGbL8
5HxQVXmCmTyV5WzR94AdrGn/Hoi8t5Zd88PK/0vs3AI1CMsdigI2dMU8hb1h0UvW
RLJZX71Xt7wfozKwsZi1rDXYZHhdH4yttGkNhjcCwHWrZ98JObqH+MzLcJTtU5fi
gOQQNA2DyimSzmmZyXEMMAOOkatwyqU/3uOsnf8Efrx7qVSg8sIm09nNwMw+4bdx
0Ww52vMG6myiNXkmlr/F67pFmY7/lj1vJfPvclWONWnxLG+be1WLxO6D4CTfDApg
i4rzEvqQlK/aq0nMQDVZfhdmbcVatzDw9o5YAIniPBzwP7nl8Th/oOO0XmAqomEh
1HjWg7vO18YTQ30JL1hmDYOHBuhqdS2rXWGnfL40K0P9NTJUczAO4D/772d7P4ON
yuIOUVi6KL7XNe4DmSXAeQNgJ+Ujx8ji8sngkZWXPUkWdXXJUJp07BvLDjvNmwqS
iGwWHq71tIr8Buy3JnvolN2b0p/ka/zQsWsarwB4rfj+R4ETupbr/KxYurG+epHC
rJYKDW8a3mRmbEGnqFHDdO/i1eOXGfoqxpgUcFi4XzN6YF60/cbRvD52jDy4eR6s
onvDtbdaV2UbyEuzx0zfkdl6qQkrdLE4TtnVNtCgEJrHv0odZ9pF1zoO4HRCIQEk
L34MIeFm9da3DxiEOq04MW0JYpRFQW5o6IqHuEWoRuSPmsMPAw10/HnMhA3b6E+J
OWfC1Aqwf78+4cCYOEnIRy3IpgyX7Xvusk9+sMO6AFOqyW0R8iuLkg9z+MCGaNSZ
I8WWaNxiDc+Epqu7uw/78CYDDOL6AbCgPEduCOWiUna2gWYy7lX0j4G3sqfte5Zv
6pTJtmih4xPF6wZi917O/Cl/lp7/u5ssyQgdvg3lAlELQK1FKSaSkCqvA8hGWF3I
XwdgjkoNU5n1TrWDF3WjpizWqHZZZojsTnyMTnIfuD6Y47GV9J0mf756ZZp0AInr
LHsWckdROFsHGz6UjDaW70Krv6nMuGX9Q9N3TUdR0AIv/6VNTFj18U6DnmJpBWru
qvuRMPiDX5n2kti+IJnYwZKEctlkmZxY9vphZw8ntHmdmxd0eIZnApBeCl2J4zpz
XF8nxB88FF9SmUFoJcUiMm2OGwwTkwWwJ8+ZOjI7HwVL9vEzoBCdOHTjSxZ6soDG
MwE2+HLgA4my/3k0NKH4lgKtTJ3qEl39mqa8F+6RPBnVz1u9eyVcZHEu1SIYg4G5
6SdM0jkTjBhm9EV7CZWIN2v7f+b1rxZvtASnIG4YdUqDQZXKntqfN27sz4NXqZUC
erl5XNx/PFoQHj2UhubU8mXxruPTdaCJwWqk4QxKhkQRAeKATz6nR2z7sfoHaIJ7
mJMwIkoUscG3nIH8FLqtjGzktaovMxTozT5sxaMyZ+3HgJOJnfLx2hYSKxQLFBjR
Yheef7L1kA27FKW3FqJrQl8QE9Q8Ky7MyNVo1aFzBrTJr6g+dvNYkudwcvHC2rlV
hnBybljCiGq5pxPKX5+7xk7W3T+0j2a9RiXiREnQ1k9ORu/jO0cegPSp5IUOyuEB
56UcQiL+XmYtbbD9TFhg5dukNjcNW9mxawBgHDOkSAY7juzqM5LNP9Gsp1giurCa
Y7NqwJmYD6UIz5AHEJWTBndINRsrPrjNvEpJGPAMlkDov4fDyitpM70SOpI3T5xb
sEM0HVxRiemrIzgau3umw0VNN5xb4KHxW6/w785eBBd9GazPSm+Uiia22nLz02YH
zMK2njEiJL7jgT3GTlg8mG06DB5VEDw+t/E7v7bQhq4iMMbSdUOumwyxtiWhqPry
6Stq7vMyN/fC1x6MrKbiZDjmOcnI1cfuAlZ+baZ7yfImd+vFddL0KfYxv/CRblNb
WBN62oIGcFSkD73cofdavb3kzmgVv4yCOopMbLq3OgEh/n5Wsc1eKWg7NSqZEwuV
vay3bn+3q+wLpeQorWdwJEndmCeL8QlcYeO2YwJo0i59lQGr7mfc7vkrXrCOpYjN
9rvpJKpJEsjFpbFsmlbl8+SjMVmcItW9AL0Bti6J9aHwOf3p2f/aZhWiuwQrVmvY
sI6Z8c65AfbRJ4R1SVNHIfQV8/H98LBtGlacfuJmpZh2R2w17dbKUEnQ4UER0gq3
xh+lZVMva9th3IxEJCYO1tP0ECG3P9Rvi+DG5uHcBhd77AsI+wi+cdDjz7xdur4d
RS0arxWg7ZRp6ZaIYWHwozV7MEojXSY3OCNQlPOz6aeDDg57sZiBEiXsDIPtq/b9
2P6AvSM9x2VQr6pXxL93GTZQLcP7WK484JLQ5O9ovBKtoXni0wQahYRfL7hoIu+s
f9/koTQJuiFDcX7EldbCQHtDyrs2Vej9YsMjh+6/hGBzIFTT3rEekMgh0ZPmAZ24
Lrv5K5GM4pbavX/Ipim0lLiUX4Lkt4Zvpb5IR0Whq4SfOo4b6ybpHH++10Xhtktc
pydROYSdZHoxXJ5gPN/ZH2Ih7xGKGThFUjtml801K2ND6Vmjp+HloAkQNTrYdtYY
KHMNAYhGkWNujgWwYeX91Q9D0Ax8oonaagYadxotPkKyGbyym6LQo6bwcNDpnWJv
BGC5G0bwPZ40klw3qtpi0ztRTLF3pUJlZGR+UblJHDKBUO4exAkME0jZhdXYUGhg
biGcyIhSGjdSvdKL9DtmMiObgjAy0Eb/4FTtWrv/NlRS/WkwlrULs2a24R3aYKqc
ZZCNRRlUzRObayLU1lO2U03dSuEDflGItz5hhzBvTWPaQtEAOdCgFXatIJQMVT8c
uRTRORHgKB+n9nCoqBvf7Z3CT62ZQ1QsCp4coXe6fklrrRwZgEm/6IsKASaysE9T
BPBZre9Ft2Q804Yc6sd6v6e/l79tenjruGnzfVFdpGiAFW1Z+7W6LV/dJ7/BXCSY
nhS4KSAGEB9baA+HJLtnuMwutialCOzKGd+hmSbsXZvjAAc4mMs6dTwnFqU8ZVr4
Fi2hWtX3L2zBznAz7UAjcUC8KSTFk3f/7YOqCtgcSZ1iuqrh3QlF7ueBG4duR+t2
aQ0bqx+ah+RDsJBGgcaj8imYvjBmyfEl0qXUxlvJld9QTuLDFRZWz/dNodCwMvt4
mzH13jh9YOd2GeRx/JEqteMyV6PD2wcxfUa8hPSQTIhPJD3uH4kHaRft7Ue//zt8
JSlPylsWIQC7fjnlGN2fpkINCJ29Xkp87vMhQd/CWI0p19zCruMT8y9oA5qegah1
yKkofjTYtx7Hcw1kBoycx/ySxvJk97A9MT04tseY/2Eg5VHLSImQOz+n/cvWGcIn
ZpBJS/JHv7K323PloOoM0OLWZD7llXn5nZvP3ZBJbklx+2YqOh/JdBc4n9l1mCJ/
F9hpfE7bW9jTwMGOzFWPtCg4fOHE9015Bk6jxNnxFzbf5wEpaiboxxixWQinqybK
XIL2O5znRYmMbWWZIEAgnOHcNKtA89IvOv/gQcVLm3WCVu/d8wM5sIam1f2qrwcL
FdZfFNO6lkHFcwH/y39Er+ZIEHxG2NJW1d2jUxUo/KZYeDpwMMFtNhfiNIhmsaq4
OQUd0t/xl4DtirDEcYgJgpm2fjseZGAqwzEDDHNq20HUhN56c7lN7aS8kX2+/Pme
f96dTzFJriIAfMU5slLDTuPONN+qcS7CVtd/h6TVPh6U+sZYTU40uKNdqddajxuq
uQ9E54cNOWZUboyl+zvqUdYGw4K25KoRCazy2ppyLW3DpoCceGLAsX1gd2yBgRt1
QAIie1IcF4WLE6nOAnFqlrmA2rCxWCDrP0TI89MYHBjiPVljZEzYgPKVe6IXoo3p
gztc1KIxf0c9w8SYAJuQPooIDCsbGt/if1c2xvxfTsvWhTVIsVTIrEZm2pyuNH1x
45M6+RMC0nbGiWSE5U/9igLpwWkHdIzjrQfoHlPMA+Sg2fwvvXudIu4VVEOoA+j/
yRUx0TRZ5P471TNQHOs5JlG73G5PK4v7BQZsQTcJJubnNLvFnCFHuaaQhL+mSETl
8dd7It1PSjFUqYYilt25L6u6r9NYd1n8vTX8Ront+bzbGygJxG9CJZP9F6F4YHGj
pfpeUW/PFhG0j3MSKbBB4OxkIbiH6Zkpld0fuAffGl5ZAIS3mDoMy5sx5mo1MPpc
yxTtRU/vUhgBO6xT/EyBPdDIswYatcwKRdC0jX9ZthNjHJ0vaKoopoQBJSPqAcHI
m24xYlKEZ+tZBCoH0/uScSSYzn7MQISthkmRd1p81ku6TyuwqzkRpmOZ/z5VOWom
cVFTQU1OiCGLn/GKn9wsBl/EyorDynyfRiF2AC3Wps6/bSTXHB3qBQ21God0VDUy
CWfW9h1+G8mxuJA0bayuEcb8pCaeVNEJQgo1h6UBA5bY5tbf+CLpvttPLRW9Lbsp
z2moYn4ACB7BOxcn3lnhPhCE6cxQMdCKXf+apCwDV144U08k4F+yAbEtGoUyhoFg
iWCkdy6h0xnYfinnOPLN26fWeqrzS7A3toXGtdlLclDSicxK80WeXypHvJGdwzo9
ycwWUPJmDD8idQkuIlF5u1XBNBZfw9VtjivqdxGFkLvcl3x8BnrpV9jwZpHi6d5z
P86vVdfUw74kMlX+m+iT9dEHGa2kWnfBt+L2Y32v+e6zkFY9IoLJCpU7d4qNYtl4
dfrmgo4UGv6TFLMbejahiXPwYubxOLQZLCN4dcH0eip8M/9DDeKAA9FXo9tr/jeB
ObXNTx4C7iyjn+208Qn5uCRa8cypFbqEMrWQNtsSrCOdr7vbeL/vKaIT/2IR4dhd
oda/qwEAjvoKPx4lQdHKsDITtj3CIVHD6It4RXfJRAwb1W3FctjdWAZZhkYdCElH
vTDKjiRAtrkr5X1eaHPueN8PgrpwYjEfs0EHtMjg4PeGiqmjRvDkfBdxj7iZ2Ejl
I85F6yAvNBU/dqQNMqC7LVI89QTY35wpQrLuckolhPoZ4j4vBW0l1kYTHrbcS1Rq
8I3bZ0MigBDoLw9YGmAE7ry91tl0lsZApyy4c4+KyVxCByQLMnZulfqzEpN+8maU
7VGnv/HOyM29mN7YYlhFl7g0AdnT0VH03JfIeMe8/UpOgmGRtKLty9BCq2yyTHad
ZQ/2JWOHVM6YJ2mKk7cWRJV38Elai69v0i8SDiulRCxjkFd71wE2lSDxCQxGZ8Tb
/q452h+OzYrhD2CUJNgo0eEhN6jJD414zi8smqQMrNtwVyqKTLvkEXNl+vfRFQ62
laiQPAQmY2xS/ivgBJ56VWocqsLhYxvSjRHf5fSfJWjK24tgGLM6dUvp7ItVAiRA
GPTZ8Vjk0z0iQQZL+QZ6E8emd+mHbdU4Tiz8vfBLkrtAXnu36zZpR8g+VFgRoYYD
DOf9qnaxetLTU4I4KCdtHFyVjX1hU9zVG1x/sdyMXVTW/6sCNb1bX4piq/h4K8PB
Vk/+FGP4N40TYx6N7GqGcTIbOIRH2MFRzshsaL5d79tcDPwscDK3AI8GAzx4/zhh
rQXavoBKPOgOuBOgbumDJVJAcfiW8hs6mAb5d9pnnjxFP2gYQOC5FfiqTebLyV+M
ZGacmejZDJF9c4PRK+03Q83YF++6iPo0rPuJjhC58X75sFnTtY0dC9fLv0R4/oXA
wKHKBrX3whIF5RicOKi7sexC8gn8KA65S6Yb0jf6wqoPfDhUUM2vRkhtYKGsJbN7
OXHhTJZjhfWf3ukAA+jLFKrBNdi9LAouXng1iZ0F6ca/Jd/50nPFn945oyT4zpdb
xdRo0WLeXZLeoNHBDe+blbkUlsizGOObM1Gk4kSOFjGX7v370ce1b/N8BReRcx7g
32Wfl4Jfh/gQSVBCSxMIVxyozid5ndcMod86aMBNZZD8Gz5hSyvjMEL4PWAxCDfz
H9KFipTy+8/+WvBXH4S1UnG9AKhJhwpuJR9uF+JQQdk5zLeGQ2rj/uVwjxKpXgva
WKbagwA5W2wnQiJwRYA2FgLhuvysWjJU4uWNEr7aOM9aRJYfh/xnCD3o1M62Y+Hk
0gpDZ6PnQBt74gXbbeOL64oNqKcDSSFFcAHopmzZjj3uysFPc2nEfDTmJplManRH
pbqTwQizk9sJ4q8X/VPtFbPRLUHMYhptBcIBo/KsFayZ2p7o4RwqfJ1PHoPt9OOB
vcxaYC35pQKISRZhRktAB+JLKDloVPJiLJ4SV8JOjI3VN2kOSgIJ/FhaXr1RmNQk
oATIj6894s6QYODYRTVilE1qnJI59DlJQn+V/nShfyYZ0GK6S6yhaB/Pj5MhiDpO
zSrty4HInkCq4YI8MeZI+yLp20dJao+FkNQPavl46iCCtjRmht52ZqnmNpf5XHh6
CWBZQX86wNFr4vPZY0tum4nhPFO2zjSWGO2kEShqzwB9hUO/F8kdUOPLEkhr3dG0
AtkgoaVtNfWq754p0b1LrVIR5xMRKNMi4i3u41fCMCnotdsFSPHexQ+1vT6rUcTu
8Z0Yj40A1n9ROwMaddHuvET2huw1LZ/PrV0WZESSzePjSgSYmh2nHQtsYqzf8Dkf
Xla/BVpdUJx0l6DyVcMnFvPpv+GKvLmGIzU+KXZkZhjtQsBxoKrRxJ+VCmNcXj3n
W9HoX/SWGj/R0dZiOSfpcx7+6mLAPIGi4JrO9ky7x+zC1ZlGMwmvirpgzOrYbrbr
yWJxFEWnjz7h3xTdi2k3YxIPs+v/YStd4XQ//Nn+yNdqHrWHSlM/MJfpl4aIFRQl
6qwbo9airJPbpAO68G5PmaCCnkbGz4mIi3moI9iA7SXFdMv3aE+yyG0J6BCEHeNt
EQBUTqebUNZB5g/7FknYRKdkxeFv7zkf+LLZW/K6MbXWCkqu6oRhZihYNLOXC+27
e5aTCdpySW6Zq5xu0JxbGwxucEeUykf5QOVDbRrA97zL8ap8EJl0qzUdPYpqw7U7
gQXRB2qfHKN6j5USHt//EuqCmkru6oD4LQnEztwNFTtpAcsuOzda+YwgJR20HTQ+
EFYIS4TlKImIq2hqIy4sq98TqGOhxFwa1/Ygk6i1TQQo1pbU7cdj427yyKMWnQJ4
eCWaqKnLpiFQ2emBsSDrKI4bSarVYPdNkLBHiCTlmGG3o9CLjAp7U2umS5jimFwT
N6DFLOjF3U5c2NmKvpXie0VKXpaJ4XB58frtUIU6Rlva++mgqeZwYTDrSyemvKae
g1JX8cxFg6hFOokwei9ulNxxTOFPrejNtX6m1bIBfo9xJ53boQN7xAdmBjDGUiG4
oYMUwkrF5Sl5wHHCDyvk3g28AXxpO8+ONM8iNmgm35JoPk0iyMwIFtkKbSFOaVzN
ZlmHBzaVevqzZ2OKS0dLiGedMjN7E91MAELgrPeAkKHDN0YXUfz0A0N+YzGFxQB+
Aarv3ECITJosZLD/g3T6ZPJSivi2tUSPHgMba25PS1W2yeNiv0/71jYter4/AXw4
AeDwB3M+Qp90BJi5RGLNLO4DvZxPm53plUIP33qw8quoLdgUg024TAbzF1PD1jWe
ejYSjZ1nsI+9qFiDhJOx2Ci8bDODi620Rb1XJl3/L6MrGZKxyiRFVzwxkiABuDce
EWp5S54HTOOd/iIgvxj1Kw+Zm55XktEysE0PR1GgiLNt/F9MC7EQcJ3jLF9a9oWw
wFHROjm3mPzVH2XBis7ay5HqKj9ZWYHbLwvu2wmw4PZljhfPUEQffKr4ScZvwZXe
DqRneHaqgIut715hziDTufQSJeG71H6BlS4kWGuVDEx5mgs+F9A9DBgY0pYXvE5y
Bdg3EFBCuQPGn+7utTXfYQBe3UykEKFJE2IdI0/ndqO2T2JArrzpvlQBFH63qawH
KZMxQ1FOEIY3rUgOcNFo2x/YmiB3Ag6xI+ieG0SUW1wDMt5Qbx+cfKQGLwbOfx7H
O+pPgF/ZNi2DMxKgjsVsq3ZYqHNvArqjVw0UgXzZcHUhbgIJPaZRLOit58eQhvZH
rMDC7RftCDtJJFgOKFUeT6lPNRroVfL1/W5sxjgT5KQjXcPrFocRajk9hNzlqm4H
53peYLDJQylyUAKKPl5DdzpyxqAp5Gd56yaVPrIfqWRzGlhJbC+RFtBpGPrJUsQj
pJloD1ril/WQrq/XMXCnpQqqNEgeJAk8QVhCIlycsIuDM1/j9I+vcmhvV5UqHXJS
5EKAcx5vGuzKdge1ozfbDnU35LnY1I7/GLedHejjmAckasCYY1E5YXO7iOFKklPX
HeUvTDoHtevJlIklr5jzryY3r8yFl+30c5TUm1QkuBMVUc8bbTqQXeEoOxT0045a
nEkJwIep0dXuiu7ELMZMYaHDheDdwJIY/BLE29QbIW9y62CkGncyAWHUsJsJu8wr
QN/jwVuqBHjehHAKIoTB8rHxt+tCnPapLbpL/TJ0kQcTFuewNChbqll28ZkIfMBW
3UNKvfHrzBo5vJjMtozLSEt+wkKJNy4ooHLI6UqtqL01ywns6WqBKwnlIxrEU73J
yZ7W4qop0j+AXfH8B01+2rxxmqllzqpmHx+BLSwO6iaAaZ8Bk9oO3fo9XftK9DHr
Sjh2AeCDszg1pbpV/awK/jbU3lmyvBqJ+31V1e4FpfKtEPiSmT2kQKXWeI98n79C
wPyTSPDUDDgFUh/IkB0erYXuhstu4JIVQdY/snhyPWE0kqeWOmvAc0IOdGn7IIOH
DGOnrFaF6Up+MfV+fgrogFhEm8VLeO9EIiEPv1RE6SreHPajVaFJJ1wrVwasMygp
5h0mmazXdtCrwg/2oZht595LJY5L8DbwOxq4f+mSkUuYcYIu3Jv39TYeOxqId5s+
rYZvfg2gCsZpxGGE69T1mjZKPo3zMCU63sxvChdxmeA4mBRdG31VC9AlQtTdZyrS
I2uXnBTH33c+Y/bvAdxdf8qjAohyu4Xrs84nKfXZwmIncnA6pPozanYqfj1g/nlc
o+7XEsVd1ORPcGmW5jzGqR+eQkTBJy3SRZ6ZK458pdfzF1z2qrGZjHP+zYcRM7L9
RHam7+a+GKgIxGzUQ3TAOzyr/bF6qoqkrZp2/SKEA65FvG6xvlkPXTnAaXIQJzyr
htOoQUxwHJXbCCRKi8TLf6cUW2G356yY7rprGwbm6vusM2UU+JsI6banszAzBRHD
YbhXql3/6cnD3cOk3e5CY5rvK0nQ1tllT9xxveMRnJeDRfSPffj3oL4Dro0SYQ4g
JIqcqlJBXk0mOjugHI9GjhvTAz48pIt3WoVosg6Q+RgTCZRRYGFuCyiWaSi5xWTv
ZGWbONLnWFREllySpqEYa73IgjOVaZa+Lwe0ix2PcDpluZSpCcHJrdi36oJg+yzk
9UmZTmOBGI56M4VtFyl/W5LdbWJNS9+f0cAfTRLCEqkdyRESjfQ1j9QvCMgaJKer
DB8qbb5itzDQPM/gHO1vO85ijG2bERaO5ccNUe7F9HSarxFrVvUiicHTC/0dH8Vd
hT1dBHWWcX9w2FCoAehXWl1T3SrXOw5bo5Sn2qUF11ryYO8+jRki8sr1r7Ps9pyx
HSszVXOgfquvnatonaDzqBzRgUgITVs5x1TjXUYOQQyjvx+Im0c3Y63swHM1LfC9
D/55fb+VSTkKAKqhF3s5M7PpjHyLAUWsGRZfymLjK3jB+7tQ+2o7RRs4Pgfu0YmO
fsdg2U/+cS/7HzZQRmNjCSbWnC3s5fuXxrdgLhg6jXtscT/x9TobrlYk57EHv9WH
oSrUBwM4a62ox9SYOI/iT0or5E8Tic549mNpZjJEQRGWxnzwshOq2jeMD7J1M2bO
L4ZhlTyKC4YEEFyE9C+xtsEIDogOT3meKmgo7rIM26i2mh9/2BXApoAF+EjxjyAC
NFdTV5tq0vD4Vfq/9lJXYYwcz5tl3b1gEspaFT2v0ZzkzujpCsEOXWcFe6ZtZI9p
41PJTbKclFPeR3cGMKWUIJYailuoJiQswg7f339PQ06IjhzwNgTbjp16EivFB82b
zjVn7cna5xeJqLt7GFmPqmOJIIF9K22191BidbJdDV4avWoS8P/be8tsQxljfLZL
4oPu6q+qSM1QU9/8HbL7fqDihhOKQn6R4lqbA6RD5xl17iScuiNS27/cDUjkW6xo
FmzzJVhhea1TcNGxNM1/rNJy+B5a1BsITle5yWW7hHmKtwSzI+iONLg5+SEv2kJQ
YnzP5pSLjXrVG81afACMLFSrjnO+KSK3+CXFA7+2u82DP+mp29bCxxwFmcbzfpo0
WqMzMpDo+UlHpUp2QrbNCgjkQOIh8yWuRYbzc/4jiwoIHhPPry/M66SGgfzdxwED
gTaB809TpIXF5y9dXUSqqF3dJZcGJ7miB+RvBqJvldCmsxH3oTpXHOGu7ZEuowok
6UwFex8Bfc1ZTwS9LZWqtTworgWC5EGkn73k/Vd+NaQl0o2U2pV0BKd1PzdUcI+c
28ORlFXmjxYErIX4APRg2uYlBDakrzBeEfPzcS/ToPrwzW0mkmSdpnDE+E+NenIB
4sk9VKLfy9R0jVVLmmD1WxBRfwYdeR2agUuZHXyp7WyuWkfsspHrkDLqtWJTunEH
qskNvW18wnfL+PtoXowLHs3v0DqJJRrPJQJ2nq3DHET1oWM3NN7t1uh3BTR4t3Ai
Eyteg764NU8OlfBigq8iKctQGe3VpxT5bY2A0+eqX+d3OWOAC2u2yPZCRJdRc+Qy
Tnmmgp4JSCU9RDdXHDj6XYapSBkPE0kQ1zH7UXfc/sWJwePybJ7cj/OywJIdEdXd
r8rl9YX53Ng5elPq9wqy21+r58pZSctmAtsx1JMsK5qM77AlbrKqih+rAevjhkzX
7+SpDuy/8OcVDgCbnKInpP07cz0WP0VP6y9oCXXe6g0eyf24BE62g3gTJyUCDu7A
Dgck9ZBlyJcpBrXMbuf6jGP3e8XJ7DZDAN0LFSLvXXqwYJyPoVoHes4P013K42I7
qjIPUKF4kaXJ9YMElQk2wIOT6rHMluw++9rx1wcGKALo7Q426dwR9vCxeguT1tKA
U/bfdkAkRVPQsY8mwdaITju5XBFZgwfSmo84k4lGNdr68z8UxdlmaZG8C3S7TgUk
pqvLh43MF0+VCZ7rD9Zbv5+/rxKqW7EoC53heAU2fu7Pll8l99CdKKB14jBKuEaZ
1yIcuHj0ksdenIB+muPc2C97ZTka45u/04rNOVRR45zXuE88mbXhQv2wczZgg+VW
ZT8DV/2sRfcxsV+oBwi9SnMLhEixuLZPb5OmprrvJq1TcmKYriKKcx+uNWvVr3HP
CLa1xbDJZlkFwSeK5gK6h2Na+7h73QaF8dRzC8SFLvQVVEKzM7/4lEA/gWfk6BPm
v4M9Dze5gx225TQSVdyFggyLeqgC+5YO85cRW9mfLI6hOnRzUMZP9DxcJ5gTBEHU
/URZJcR9cFSLvKE9xj146CCsIFdVV5MZk3ALJNTRlt/BBdwD2EVujtCh7Hu7DGSM
X+mCiw0adPjghVToYA8jcmjPyzuIZHF/fsh5hc1KITO4oEjleM40eVSkPnSsj+g+
N53qMpYSyg2BzFK7o8uQQIEUbPFQbe8TCOZhzPhWdvVVjLNGBrbfaGVhWNTQG/St
C0OZ+3c9MQColU1d/TUl78Q+EBbgLVEocbFDl91e2kMwNaDSMObjBwcCNC2AUHBS
k2Fsbyvyf1zYEjJHH2LDQ/C3VxhWj7zLnanlVLxQUCRRtZLhS5k7GfuGOz7E4fuX
zxPlwpPlMOzI4zYChoG7QEBTW2FCGv4nja3CyWBkiaNJg62/YqhmbgoJuNficnNc
GBpAH68rT3m/MhTrqU+wc85klFcAgJn7nGoWrfXTtYasaf2tfD4RhNChNcxgOxWw
3g87UlRz789PO8XLZTFhkx3OEHx3NWvOfDN4FKFnoqtroI+pR2JJZBhNk8PESHWm
2N5uvPoJTCD72C20Sv3busn2yxbQJt1ljsFSe93Mx54LAlDjzfilVOJXKDQQwIfX
eGHUggVTgWq/QkJMmdDmD12xkWPUWE+uKF+f4dJ/03PryV7MwHy2M03cMt9DrkHg
9runQKUlFWgxRkGlGOfWb0huTj8Lrm2LYzZ5fGjoPNosWeGqg648o7uDrPDF+P3g
JbN48vA4Iq5DbiGbtnU9rMOj4UxDAiuXXpI5EB76/OLWqv1u+Lf41s7zNisHD3D6
e0aTom1m+1F+OGuJKoRAjwupqWZa5UGXq+ayxjHWNRCZ3MW8yKlggBYOv/pHJGpL
5GX/DNIW+Epd9CeXAQOKQgvGXFSUY1XEWTUfRiIYploQCkXvnzrSlXiJu7QbK8Jv
LpvHP+KsQFSkvdHxtCkoRjkiuFiAQgHg3Lv0Yvx8FPGRr695m59LTuYZcOuhbK6v
mPfV4yVSizmuHOlsUJepQwTUr5tmdswjC7imN98SJ/zin14lIxswCgJsaIQiQPma
hWqpIts7sCEBQyifstyvcV80J7acNa/VfuwMonSz4AJKBkqudU6G24qUYbSHindU
cS0k3aUjxOYMuqzs68qi07mtEjggs4joQ3sobe2VKT74ryz8ejzWYlUTPF1JD+sH
ovVqg1xVAlXcSYkW40Ue04Gbh3XJHY7q1Ht7UwiIZrOcIJkxbrfhBo5FZ2+J26g/
UHrg6aNaKruOF3Q90VbUTAHH9Erjf/XTjlwea0vPb5/mcubpd2mH4mvQGxiYkBQl
3EzVEbaKb7pd2uMoI8oH/nCfuD5F6UAT4lYRtFeuvcsq6pJhDJHUBeVDU22KPoLI
ndSf9lC//Cs5B0a/iBtRByXW3dcU/XRtjFHUY9S2MHXZMjnfLe+xeLhhpe8aNtzg
/SSD4bW+7UvjWxquR1jN4Z+/RBosPGen4ZSWUQ9hE0vUf616rXZWTjoReTpLWHa8
Cq/Li0fZT0cunXFiKGsHjYlSan3I0+X0/7oZHJf3Oy30e2+baoWd3wagcmPkDC96
6JOudr4isejgR3ihNWMML76ygXX8Zl8Y+F6qagYLLbXQwJJup3uloHgO6NxuX5rR
Cj6LANms1Gi3l4Vp7uByVaBt9k9+zG7UNtLsbqW99VuVUVkIr4aMTqkK445kfhO8
mNiaX8PhlOSjyDg+Wyh1UiB24+whZFcMjTTwduVItTADKY4ysZB36P3OedpTBoJR
SG1amhPJzB6hJQudlkKw9yAkbKLoXE1FDFCszNtx07Z/Xb0chF/VQI2a6cK23hf4
CxQ46sCkpQDbiN+ezu996cMYhYr+A0l+jBwSnU0mDEo5kTQEx8pezKFRLehFv9Ih
MOm0/owKUk+p61UEitcjZPsNeIx8HvqSQ6SsCF9k4C2yKVXa4Fr+3I0tlhQxUB9O
1Jk/lHcUnV4ww3p8yDu3fk+UNzB58pEshn9CFPNziY6JsyW8anvmxk6di+d6iWwm
4meLZ0TzYJWxB3Oahl1GffNNCGXpplfIgQ/DvJtZUEPQDTam6zG7hTeU3Ytt38tx
iCeuUR+FB0YHqsCwpe+eSBPL7A/uy7UxkUGQ3AomkZQ1Sqe+0zCNWQe7EnSb0h4x
dy6qpG9aZ3vqZ1Oi1/Ih6wDBxjiNHVj/x28WMBj54zQqGCV61D0PvFRFuBRHEySd
ba/j0wSH7up5R5CMUh7M79zglvqki9w76ltlU9lBu8Gk2f54ToSVKlQYMiyD6VyK
+9neLgO4BtghCP2P9zPJC/Qd9TAefm5eiZI4Pn89/GiHYnfpT7NwPKELt5Xi5lfQ
iwbqe42UUiigbpgaNq619wbCOEOrxGKwHh9g/qxW7K7iMQ6m/xkYfH784RpcsP6u
M6ithe72Q9hdRqVxMyCFj2fTRU+V2VlnV3dF86jgAEE72zfzF4jj5w10mDWyNwdU
xxZcrFN+ALoLU0CW9kpBLkZqYDqV8qQVZYc9LSQJpnvPmoeTxGJYabmgYGH4r8c1
MsSbjB+JmuWR/GepDsXTLRWpvyFl+Mb7Klya4QliC3PxqIDub93A0CKP1A0TlqKU
G1vEO6YF4YdBVsEfW3dwuwJPpA7CQ/e912mlPILMX+Pba74XSzW6HY335w0Aknft
8U0Qcfbips13ch/7cSAANVWKy4CbRId4gv+pd5/3zsCXuTpJjQ/AA4/0jj5535/q
+HEv5yRt5EGQYnLYce+FWiFPa8o2jfj/JABij0/rheJWx4kUrPecTaqPEvsMZVjr
+p1P3QwCFBhwhLvuwRbQiLatb7Mki0XsBFWke7oM5ANKd4vyjDqrHkzXic3RA7ho
1krT36PtkfEtmNsZ2FgCny/BaShcLHHTjQLcD+jhYF5NozHHfti5WrixCgHNtvyO
SSUzBdDupM3Hc6vK4ZZOHRS+qiuJkAcq8/E8UzADXI+0QE+EygHV77JCPPtdUl1S
akHghmKOcaaYSNtCuSxGMAhTDNrz0woNwj6IXjtNDa17s8k5fnfkiJQAHI1IGVx/
v8zrICNZk11BtEyusbAAP/9JWlXyvfFyhNVwdlLc+1GONdtCBmyVB5ow++P/Q1CG
2S/EoShwCKeCngTFzwHEFThqGTkRpsP9QRovGz0xq4EImknO05P5lalH28StZKhS
jM/IKkhH7IgPbi3uLZQQIwb2I1fuTxndkLdbQMG6hP4D+MH41JlhfGTqi8ogt/45
aaBvQQqmx5OrBACEIOhdkuwMpqJXGgKHiyhp/X9c7xGl+L/NvJafvcAh1IleFUNY
fiAp81XQsaIq78kmV/pLCn5yRdXUvUkFsajecK5DOuFxj8Emtmf0rQx4FGbSctTd
6XdPTI1gTuKPZNKzVLypz1iXyvKr701FecZtVlGBgI/zoznvbQYVR/PPg+DgPcJY
bh72CK9r835fUzhKeW0bQlEsyMbfjUfGOOFow+Cb9p3RNYB05Z/YmBBsRPwuXX6r
3rbU4Jd7epOd9u9LgzHW7G8M6c4tpjFczwGRSmp+4DXPDmFBwM+Dg+Z7lr1fh+1c
NJJZyjE2wBkR1Z5C9c/NCMoKCPCRz0K/NMkob/bbKtWQDIBApeLd+0vold20vzRe
EZlfbkXchuZdIA8EXtzFO5/TIagCHOAAFFYzFaNiWtm4Y4cPkT5UKQ07wFakBDvn
flRi0MN4eGWGXWCNgt7pHvgU6fITtKGlKpMt5h5uqtfVnOsdBYFJPQi+zzuDqKBj
u4OUC/PWg8zXERIY3iJChrLZBOfAklMHvwmrcnqVsNp/66OqxNkNIh4ZuvVaRiyl
Y4AP7iKjz9JZ1Vo7Ki7IZRFHW+7QLR67j80Iei6kO3OYkUN7iBccp5IxMDmN2o3L
FpfRZ65qfq4KFjT3UZtud7AQsoNQ62rL/CxzjOkYy370sa+mFrzbDOCQPMJyU9wI
ZS4FMgfwGyeMSDeXg8LFq6KrUIZxRe+rJ9jJnbYIiqDOlKPPIxPUgk2qKTwGusPQ
4Wri6lZKuepLw0TppKk+3R43J0DBePCamBvH05+olxGCMa7pvCffksSbOjGV6eNU
We0yzqzqyr7WLh5Gviyck+N3QO+O3CJttgyzpjLeE9PtqocBgTkpajZaMxTyQgSM
jR2LIFmOf0GEDf02qlJD8qDlp/DtFJi3R9doEj9gQmaoLIbmkp51EQqaO9Ypop3p
gzK4loBdXTSE/jWDzvem0xs8kCLBc8EDh+oqFK44Pxzrrq/ta4E/ebyJLqqoqBpv
gIuQpFdK8Jxko8XzkUuQCJ9wVgBRQO9k9JJ63Cncew4J6yQq89dweJXfhxGgvgqZ
DWWVIMAi67h91k8IqbcUL65SgCwvnSPfyGiSGG5NE67lo3gMsHaUmUPlBhNz5Lft
odZAX4K/RbEM5yrZhtesxT/gtbY/HwiX+UoSQ7OJ2Ip2sDlzB90c5AjmSaRiUJnN
8rr+5DB32c9kuMUhKyT4B0OJEVXfvdvXPis2y9iad69tchfMbAGoeeoZ8UBMOKlI
e+c29vjRfYI3VqV5BIyWgpJqVtOL16z0jf3BrwPi1OHelHEU+Sa4R+T+AkEIhNX/
eOhyslxUMsqxnuE0kMj4g2yPJ1VSu6ww2aFaYsOsz2RWEG5cgMSDA0qEVEkc9k2I
H4OtcgXxqQnqMTPuM0I7AJruhN9Kw1FKhC4OknjGFtbTFM3pmp4IGcaqc+s0pk/5
AW/V4KqL5MK8hBfoIvVzFaTUTWgtVkUP8asczWI1Zwu0QLUjRFnGPYcrmrxy0ii/
Tesk73857A52NrAxw0QQtqDHDJ5m3dXPSau0FShzjkmTLVjJl7P0P0Dx0Rvn8tl7
fzjaGF76OCIVMT/mcLlzeb45GO/yTgihuqVOmFWCa1Kn83wbDrjNTkR8DKblBOKG
A4YU3EUDlD9xmT1mEccGV7J/WbJPa4WamIXffrUpXxs93Ss4vA/mViJZmCaoqyyt
1QIl0osbqNgYaE06l2S/FfNyN8vpyh+DShnbmNUsB9qLkUYat9QZp6QJwBoMepgD
H8HmZwm7XuWT9RBfJIsLw6Odpwow3r6VVNe2lJJg8NBt625FaswiS6y/jX5qfkNb
bYjxSOfCExplaPLM6ksJnJxt4OCGFUacZlpFo2aYIDEFGzzFfwBBjtOX69ptQb2v
2EfT5y1rQwBvKsa06zXXtJky1KUuqhordfGrm1yVpKb/nnTqoY5VshaM30l/lBY9
LNTc9uzQRwAKBpmby6pQWPns95KeBaGpONbGE/9aRs8KBRKADlgKEsxvN562/3+s
AS2RSPN4WagdAE9VbQ0Ku2QuOSDFtfsymneHCpRReUc65bx1dTgkiaahfeZYzb1Z
Dk4PQP1rM82bSASfrNSjsxj4t0e4PfpCs43WqMs3/iGmVjHBl/l9diBfBi5+3m5s
IusUKvlwKtxXU9Rl6ZiaLCtWXcxnaPyifIehOC8l3H0TQfGhmKZmEN8IPZGD69XJ
YeJFb+35PN7MxlAIXWd8cR7txqJ7gGK826qOWu9X86QsOrckt1kSMUQcrdLleuvG
A/kT5fXddktZZJZVrjiNlBtacPe5YnKTg7f+XN8+ie5ZBZ7kCvVjg2gKR5hVDEiw
CMjM0wneNNd/CpzUImvVFm2DhF4KCjHSjhzsN1p4iKHAPH3DWG4AbWr5eS4MfKWI
qBFkWXVjqoxCU8IfMTiYVh+1NzTcHEHF03IdcnDRPQ0J5ATyHsfW7s56mXq29Eim
p2mGC2Q2r4ApMDCcqwFTE6sXOpd5DUVjwrQ8MIpRdR736+wtcsJXnzuFcnMv2qrF
mTh7ZKW/tzSKXcrzW79WvXksI2kc3/ekd4Dc367keAvB6DZ4rjeGVQeqk5DPjYET
J7oMj8C5fqdycXPKvh9lW1AC1YIAeuAjFmNuWVB04FFTjhX+rP2zfaC8kNXJce/o
/ZtbcJYHuo91sIMpR/9O35oB09YUfk7wvxEl7ScK1WFhGpPEPJa7SQf8UV+Dphb/
/mtHOkqqtEGBlptjLwdbqApdc76f9Wdq0+bewdejd+3q+yhWBDxn+i9EtijUWs4Z
oI7L3N+lJOAhW+0HkEo6MDKNBUtOAKTq0VlmoSmho1oFmQVDtByJH00q0WlugxuW
CZKpQ8SmrQI7q7QTykI4mV+OOuaszXMsYKAYzuK/E2SGF+ossD+kUVkGnlis7hIz
gRYjv2NlPJFV3qNZjze9942nsMHGSj+dRJIJh10fTP/Y28qq1w04AyWhnvi3QM6G
7/jYTXIw8rvvue8lGSU7OYU+zl61KzojsFW1w6q1RFwOx9hT0gcPY6LHxJTSFZMo
a9bZqGLKJBwRJI0cRyOVchcT4iqWVFxwaMDNdYzdh4PIci1GQkvNykTeAx5O64jF
7Rj0gnqdTK646xmsNY63SkGjBdS/z8EW+afrx6XK5jMxFcdkXFua+2OvvwM8Y8hT
aeNpNL6i1Gr1+8/AVR0Lrip4rz/MWlVIa4pfehU5Ahmj8Aun3NKOf4HvQRT7hgVp
UuDYUbVFDk+j/IVOb5hwu/Df+58jadrENF2hGvB/6xN3qAAb/9s7JWalFIYDnwRq
c86ger3NO+Qx+VkrXCThd36oOp+v38rXvWcyhrbf6Ou93NUjC1+VW/R6XSUCU87q
0u7KU/yJSaIWp5XqQHTKWcjQvbqqdNUeNM3j0kmzsTEMmBKJVpEnbShJpPKOzrmK
gG55qi0vZIzNV/86d1YiM7RlniM9Vg6WF0z82WiXHPo6mEuhLPISv+JxMjhrcLQK
O3MBYKy9350m9a3z3Nr/VcXD0pdbuQOxgtzjogPqEtHg32IxKYhA+TU8erVYkHhn
UOByaiQzpfmtU4Z2pjyI0Xeoh6nWkdQ52RhtKbVxzka+4hasna309us+FkQZ7stl
guMHcrwzCkIjt3ENWWetK9QMHZDhcE/SyGpGv//bru4ic8ltq5G7tHhHQ5ddCZ+R
go+Nq3A3sJdCa6J9l4LlUh8XtCyr3yz8VsSTvhw5RVcS2qhBYHB7WyaY73fD9dVW
M2aJlosxDvWzasJNC8TUhvRKPAvbfPoz944gS+y+6jdi+/2quaP8aih6n3fkNCBz
TrliND4ahxoeNaCrrL1qf7+zL3oj+4Sa6JzIjhq26PARY4o5ByFvcrCCYQ2TVhhP
6T3nWgQqYBEqF2cayaSAAIVFH2ytISmeXMSyYYGNcS0BJ5jqiNbc94wO1lBShwzH
t0Tb5ZJ4gPZMJ3YwqvIAfzF34BShHSFRIvAxL7d8x4B2DJwNz5Asa80GGFDsw/bw
XZCvik+XHrUJtpK9YGsQ736LGTiUM11zbYB5DwKMjMXRyUip3Bbmou30cHj6dN2+
F1tViU+/c+4/jGKmWp7HDNy4P9ESNY8nj4cV72bytOOXf1LGwjux0aTLZHaP16kz
7g50RzDW29lEKjs6n8kP+5aPa4dlLmxjMLsYFNggT1NLHx/PS3l+u2lbUxYYTjXG
qIoUjKjKLWMvdRgZPWTrozsF6izsUOydzadiB65ots/iZqTnZbMOdTVYlPQyrWq5
rEUjQ5NPTvvLlLMwRrXhyr4v+kpjCzrh6LkgXA6jz3sc4yBTW8shRSEYMzIkjwVs
wRmHPhK6tBB3IS0eMKAK/pP/ZUIR8ahQsciQfX7rxEGHqrNiWb04OOz5CJAFg3Ch
6HJdtKScH9rmInTDFzRzA1RhGgJPy+3+yQYoczBhS05Km3u61DOlsOV8GbkSSEUU
7deQ8FpG6AwY3MbQQtZAn38991FmGbZVw4cKG8uc21h7MqaUihyFWMtNrG6WPjKV
QAIO09cgDZjx3zPceoPszMfoAcqs45P4JsTzNVdR+Xk3BE6w2rZGJyEip2Wyzhou
kSDPbCYvnovvsvSYlhGfoUCvtXqul8L5oLpoDFwo1KUhM3jsrftX/Mz/vvtNVzJ1
IlVLBjZ+CJCOj0XINC54igJzrr3JDyZXYXZKGHjzECoqLCyd/p4IWT08uiCmr2Tj
DNbPV/avJ8GmPVocqI0veJ5df3PuYmZ709Gax44flx8uYpILLidpJu5h+TgUOg+P
Bpdnk5/YEwxqUdlH4hgr+LfgW6PHiuQv+sBsI5VhNeOqkMR0EV/TDRW8ltpjt92S
2cMAXptmcrofhqdApewuoLUdr688cIK8o2PbyP1sOvYtC/tOnkhU+BA8gzrPvOg/
EpQdNgooH1TIxEz98oZ4Hyu9cn7jiI3HvXaPv97j78WrhxdkeRoVfaDVTDTXperR
HstvobC/rubi/B9IW0ITT4f1x2UHKUzI2yVasmMSI/8T5x1o149uMZDG8ERFqAnS
SBKHn9gXzrlZQNkZC3F8u1B0winbB+4W89M/PA+G3HmtqUqNOqFA/6/j5Ww7/lOD
g6sdH+tCzPY5Oluuwl8vLcvuYricmbLUdYPkHpKlmn9mOn+7gG0Z+Dkf2ELl7Zpn
W65+s4zbmntMXch5DgTcU6a4qZdPCUMG74j6xRheKhUTZCF8XiSCNvohNFBUIeaA
uHLcD4SGAyEzKjeElKfgvJSDfsUSw2QtbJUfX3yIGg81q3lmYOdtYUX1YxfCtAiy
18Qhbb5YP1tIUpNihxrNR3ZrRLvN+ZsRd+Ks4dWyfB8X6euzJ4VkpHz3aTQVs79/
reldiHnmTYKnMEuylNCoqQUEIqBNvnJv5Wa83DKv4R8YE0Mkz5GPJiOU+a9SvR32
+QhbwAPd/sOlhRfoeglSOS+quqi3yO0h7HXvFpRkOIWTYDsSKvgZyyOk/uuEJV1g
/HW6GykwC62HK6ThzOc4D93ZPwNplKtL3SmSuauQ41Bts4gMCEr7hNMcGcEyjJ2n
eqVAW6A8HifRw+jCSloXZ1cw4wjNnpNbM3UyPau+oC/23lX5JXef6gWSouJ1Sdx/
rLps6eR6kcU22X5wdcQkrH7CMogCoFDd4Es2i/hSlKuVIBUsu3bkV/nAhJMsto5u
aBOGtNkcUz9c9Eqe16fSa3Sf/8NSdKlUe/deh21js3fPvrdZigYfcsbCtSzxXOnu
qUfnX0NrghWmo/senuGeklgl0YSlWBXp/4p8VtqCWHxUFZcAmv8vmeK2EhzFVvPM
iSLYbokV6KIN845vbTFYCftRogBbUtXvWuZpRXm9amfQFTF2RUSAAXoYc/ptbadg
LAoeiMKGBKfKT2QiKp7t2py5k/b3ffobAiHLO1sRawisIE1DZ4WP8d3F4i/MxXN1
Ubifg/HXzTMZoIx2v7jL5Ql296+WrrFBwzvr/ib9dyDhMFAFPjRCsH60WNHLc/bs
H3v2NsZSBY3ix8mvJz2VMvh2/jyxcn0P/6vjkjdDH4aGNZtYtZzzYiiYHI6Saj1G
RgvfwBnbog1kwESYqzln5T2uxH7pyOW04domg2Sn28mJ/sXTdHv4JYda5b7Nq/7b
6NjYw87G9mH6uE7i8RogrMrhfNhLdApHDqPoPodGAYoY1CyrXd85ATCSzs+5P15z
DYF7NAos7Q338F44qxEdoOIBFQn/t3DzApPrsQJvegg/pH8oVPXuAKtA/8H+9IkQ
4XiI65V6htwVNYNpSDJVQlVojE1fQJrX/0lLHSIMznm36KUNgnK5gAedySIcmE/k
H5Kim60NfF1YQKABfS6mB4kje08GWf1XPWmyz4ok+k7kTAyrtHx6rsHl3uU09uvJ
yaku/N4YAkzCD9PFXKUga6aVdb5UZm5nHhGq+5Q+gt5ikeorO5Q/zGzLPCQgApqY
2vOtkCbNlcj5eFnDsdSfYUHJM0yx/TGMbnNQZvP0mmnyJ2+lN9nLnFmIJNJvuvWT
2ZybsNT+6YVZDjNix37qsNrqftT9GxrV0piHAkTXN/A0wia2ffqQaZuHIMBVusVl
tbeWyYriM2zuXfVs1AbIRg3aN7GVS0YexlS+FceSNiprZMmRBgTafd62bx3aGPU1
C5iG6WTFbFBfgewdendfJ1DJmioLTIe0m57gyaG/kwTVF6kbpzN7uEM6w0VhMW6q
y8wXmGJsJ5cAJD/s0rwos/ZihIZxwhyj4MBbmg6Mv+kzQuFbN4FqnLT2PJer0Nei
8HMGYQXiX7DZzEP3K0kyR6i6PNsPcSU13u7uM9c0v7vn3/eDF70f2M4tMhxhAnVd
F2KwZ2YspCR6o76Mryn7bKU3P1qnUut9BlLlkGvBfY9VDga/YocOZbrnpZMBAl4M
8y532lobWZxRmjZqlwB0cr4wxUGsWnEVDUFlwvq5TBmYhoh/LwNBdoOhqJ/yTB8R
mzy1NASOZ+w1PP3LdRWxp7ezbexuapMbCCfHwUsY8G7nENtcUKUILqtm9UVgIexN
aMO8nKl0RXBA+0VMRUdpQE/3/TUd2J6ZedfgWbx9w+Y9sO43fa9umoTpOqPWTa29
L1URmcw5c09wrImWMZjKuQagWyIe3NOBKaoieB6TZ05NazXuPUf8oG7odsAiGgSQ
pDjH0lcSmLvs82saR2b5bTHLjBKGqJk9IiiJ+fLxh57YJHTF5hKUsiEC3Xvq+D2/
NzVl+IKs9jeFjYmHxh0U4JejPyAq2+w1R82Wacaqzl3STo3xGnpT2pXi0v1+0+Pm
sXFuGX6EAdR1VQ+NOKlrpdFctW8pqFkU3fxAjzGb9QstPIZ08d+J5py2tg1MJZtb
VZIU56BmrBX+BqRaRzGmRnmbKOyX2TLy3D7cABg5mz3NeglN8L9v/3sEQWmnbjEc
AZt/zFrQxCOwOxxtQT2VMPAjTG8rquvLSx0I/dH+tbgP5wb4BRe6cQtqwttXFJXr
yq6+ptrF47cbV/93DzgG6Ea0gyM5ApOgs0ZRyWIoGGmE7W6g3Asspkuz5okqpA9P
Rib2XdmvZaU3jGwMCSAII8ro1tWNC26tTQkbTxp5TVH676VfwVhj0FcXinzcBBlt
3eVG/9Vd7ymrY+VjjF7DJwIZ3dAlet4sQ0L/aUS2gIWij2pIj3mYY0jH/9rzvM0a
hLRBPNmC3Gy0A5Jv1xDQBJcd1Uz7GtCUFTUxS/HgvUq4tvUZQWTn0ZaCfNYMhYfx
+XvJgiNabH4svddEKEhXyNIgI1KJmKJYfIBau95ppYcBe1igrRWJLZ7Mz8JvBvfQ
OidiK2OXW1vqt2vH3h/YUhDb8fvSow7q60UJAyI7MTkjLnGEv9NitubLcOhDhiYQ
wx/bdecoIE8fqjAqlZsVWZxQGdusRQY6V8hBfPEH9Avkmx956UoEbKS9wwoC9KG7
ZM+Ny35iOpzw3SH1dC0h1PnA9gNzhgdPe45nTworQ/qaFDwz4UfrGNWblSOzrrf+
3JSvy5x7Q+K9ZRIOR+yGeGeMmOzeRsFBNS2YhcuTWfPxa3TBEZyJiY+rQ0J5EfDc
yEfQfSFRLUt4GehpJ63rCE/yNch4T/Lz/x5wMEOVAEHetRv1BKg2UNazxK2hyQKq
xcRZ6NjfKY5phtligliFGHORPRUzN7XDUYmTDIdtesDE0bPYahNu+xMUwshY//S3
EltHtcREXVIlehYDZy82lTdR6mnUJwFDZYyRz2g3FXWfkzL6YBvBVrBX4cBtIK9l
NVBAeXFhlDkiIHLoG6zzA2LFme51z5cEVz9bN4lPzCBGmW8D/mF9W3AfpkyfcawH
FWrG+alrrNSNovuNYMbIR5UHquqWu1gsib3bqxtwg4zWX8LmJ2Nvm1i/kHMjmRH/
3WLaYxY03/THh0OwA891ZIHcZROoF88AdzksNzmsppKE6Dqwzi+A/6FZ50AIO55h
XVrovG6MAmgLMIrXN928aTlCTcuC+SnJA/mx4WJawreiPwowBEP4SRgmEjS89/sW
CPvfgZe03tFvE02NYVwByo9+R7hT91CJxxT3MLZe2mfNa5jetUdFMOg4rGt1gQeY
gyMvJpEMdUFXHbxxfZuaLnvgPLMn23s8qsf8Txat92skYvsrfe1ry0T82Ta5ZamW
xwRUrT60gLlwJz/qpD1gYsR+7ywnqi2dsF3CbTEcmN07ro4H8UkvDV4hK2QtgkhX
C3WSyI/cWlP1wmDZuez/a060eAVvDbJcB+JhmbX1z+Cw8teHVYewor0oY0JZmlZM
gw3NxtdTNo/0UxoIiyIoVPOWd6u/t1mou/gc1JXd0S1CkYS30Q3GAVIvARhcAu8q
i28Hfy+ez3ejFMj1f0lEWGVvsyzvE/nj0YoIPJMDUDWs6J74yQNc4Fq+2WFMrPJW
Y0PEQ10GsDLVUAhQQ9QORDsnu7kLY52d4dYSGGH+yUz9XVLu+AWugQ//3K2wqous
xQiOSbWlS02wnhhIXMWhiTpEFWpTzJyDNsHhJwf6gQLe45u0nJwsFvqf30IUu26Z
qjRB2TB9ApRHnY0A+Z02e+ox3WNbx3lI6GQ8F8PQKMiG3jCbZkueVZlwNW0qs7L3
Bw0Fts2V8edg8EyycwvX7E6oxksYdh+I+uK341xB4V+YWyWwDEvW3fSXoiRXT54t
rXjvaAACR3lLfo+J248hM54vHCq+sZUp5IIAb34hwzW9kkzjbGRXDt3ic9GcnOUW
8lSVacFcckiIhb7Vh/Bk3TNYNydIDkUGLi5u7ScXtLgzy8/EsRrvltDx9rWwf4u4
v+MZxaw08mHnknMjXBHCw7auKkAsFVSGEy8BBkeVZRf+YPFA9V2jZZNMCXuhrUIe
mm0bh4fZrX22p2NYXyKNBdhfZSv8/q2YHeD151y7olCHJffmP94ijat6VCSNURZ3
RWq3lezwKaIaqXFvRG7AppXxIly2Qd4+SeMdPxemEu8QGlcLYu/37ShaOAj0AT01
BRIzfoT/eafCDZkLXqFURdwv+ceXj/ChhPYPZDaPhohfzKb84xJcYTUt13iMDH3R
xQ+05hDQaszNoeAOy6BmtMrHR5k6RObP6rqoFVZ9Yuy2oSgRcW1J7sWm1ltn+WJx
5BWjmZISzsXptk8FwipXlW9WydTYFF3l3F4/L118u8TS4pPnBkKQctWVJQFAxBgW
JbLCCY0Ohuf7uPPdzweKLHdMUKAc7VmIQ8+IXOC913p0x2mJm91Ub7GuAADPlKFQ
R0HYVYwZrN0pHZPGZMdsTrOBRLciTzzCi0qOVAY1x8scoNijXIuvkKoHUr6sr7G7
mel1D/MaOHZf1xzwdFpb9xdE8ZNVutxcMRBpwGE2ez7Ux84wdJ4PCuQxCHQda5+Z
BUZKIXiTpR/bRSmcl3h26UfPYA+ii3b6ReN2nCJEn49Ujq1/cM6VC3E759uOmHqm
gS/SpV5jW3APv0H9ICPiFpJbq23LD7W49MFfiLSpOolbmIO2GspFa8HUGDsaOHnK
nB4cTwLHu+N4Q/Zc14pcpKOw86p5YEY3qz4QKjx2kcexGyB5CUc4qSJVZyWXOgvC
ix6Nrq4iZdLjj89AqWMBKtGO5pwXQGN3+HyoS/xlTxEP34NSde2j5h7uExm450lV
xfUMXoyTnEdQANuvwuPHNKFNdZP6HJIdBl5NwDWqUrElgPXakoBE6SyH7SclNLDj
tqW9hfzAqTqN+96rtXpdzs7hyac7Uy2xD+/0nF1zn3At020EQ3+bhfgC9ztHkHR8
wYDmHR7W2x4HwuP8ThvWpRKk1YaQ/YDSb5U9aL8YB9D8cPQSjLSt+ublzCIW6omA
eVWoMkrVts0tQpmoCDAkgnkor4rFVEuV1WqFZH5+HjnTLa9t8brd9ZBGkTFcy7e0
9SoYPpNJroXdSNSJPZAyPz7uN6E2WZGP/AKTUTKMqStuacf+hyZBvL6i0z6bCYYY
tRP78zXCqlUean0DgrwmAuEg6u9+VsqHgV1XZjtRUTwQtDL7yRU/rIJF0oopAe6J
bpURmLbdikDlkfWYd91r18HQhDKzsxU/EKlqJUrZhR9R7yLVBpYh2/j4ZkcipKoD
VrwUosKuG9mzKQzC+l22g/SK+5cTHrBdEK3FRFM+71hktwj5lAZkSnnuzkUMwB2k
1fDRtZFB7A83sSuTRVvJfPAw2GZ++CKaGJsFQOQar+AaLQ5aqM4LSi+W1zxk43U4
vhP2lNk5nH48vJHPs+ex5q6kGvf1fAJO1yqtJV36FWsRNIWKgHM5tlWKeWaxcwZg
4X6wDk69ByPJ3HgMBE0lJ/TNbOYkPFUIEaTDiDCHRsaU7JpJ+cDhNqpIHnjr0hL9
dXE9niKHi36vzt7dsx5EINL2cWmgnl70LdFUtTpqAintbuKtGzUAeH4yV6+mz3YK
TqGbqhENv5hKwN3so1HAnKiVI3UChtEBR60gMjissjSvSfLVRSmQBZM1S9LPaEVH
LJnUuE5rIUEu8jTRnGD5twwKIuVxo53WBRixCl8QiKetxU+z7uMm7BIHoGLHyfNI
cT6p0ygSqkj1Aw6A93PYbnRFBupj2I1XJoMR3Jms4pdhaehGX3aGgBKs3lSfyvCg
CD9d0ALF5h2G+RumfNzMLVIDz5WpljbgNvRo30c2ahrYVrDvrqJLYiHPDLZDRnc1
bZn1+XZjMgrC+leMTJxGxpTfqQMM0I2xMzJQi/DzqS9YZNj0Dtb0rt3pwgnb3WVz
ixzAlxvbHIyKPd2UqTW1I6K629PxTsZLMU00nYKnPsYpsLLT+zFKoqyEjBaZN6pC
762SFFFXDEQ6i6FoVlZZ9s1y1OyucjvhSx7MRYGpEkYvpEtCkhPK5x4teVIGvCiD
tnHcSyXfen4mBDCYL6zwIKkMwuT3Z6HyXu28b7cJk93LVhXNQ5MNI3rRlRNNJbpX
9t6H/ki5oGKdhnDd8C3AWsB0HgcUwZY6FGcuni57TwlYer9p4LlhrJgyu4Z4o4Jn
ThEPEny9+17rH4eewZwSntzuJO+HG0kyqf7CS2eO8jl8JXqH6g0Dl5IUWa7R1XJw
Kh0LolNQ/iCv5TQdEYjYvt9oR4Wou3Dj/YRK7oa4hArH5oloWR6Tw4tF+oMa1jvv
oDigjcvnzpvAQ9lsJh+wSksV7G3YSfrapm14ohE37Nv5j1TUvguyFb/gt6/AreE2
1fZqIIQxCktL3w68KRyU9lvDoTyz83ayqBAuYbbS+KkVhBrcIYboZEcUuLIPSRY7
Rv+urpmEaeisaVwyS4RCOZay+xvqgj9FEkAmOpwJRbwfmGwZ7/84vY6jcGCXSIjo
NkX5xl1QVkOq6/HIZ7gV+iYQYBG4fvDgVliANs/pe34vYUwoy3Hovp8H7kHoL3k1
QTQ7kjfb4NNt4vba87nhSHK7TuTaHRfUh7WLjf+vCq009JwzZ2tznnYofH3qCTF+
XnAOb1zoD3E64747HAlp7ZXYOHMxHsySgS2YXD3OKUno7s0ogfyjoWyXg1aRS0qU
ys2eCDvCQGpO4KzhgwUoqiTLHxfN+tCnAmPNwZvXYm44AGt9O40kyOyJ6VNwnfwj
8V/acRAeG9MvAB9Mca2FAiMxK7OyGDkYTca0+6LAuqe+K7JVuHiggqgJa52OZmhg
fEZWlQMV9IzEZZKqCOjXUH7D1JnUB8MGxE03rGSWXGqXwLtQjHVMU36Jr95RjMoj
jsEnJfvZIwsqxqneiqyMNKJTqNhltMamGUOwJ/EYjoCpxhvFXI17/6JsG1dgM5Vu
PjCq2ZvYRWLnIvaEt1W61ZtD+wDfqgIbF0JVR7Q+A3L5r64n8OzGeZUArBl8aU7/
rRXPrnT+txZsRCprXlGzg1s5npWi70gR8sXrROfHJ/kga9sUD7uSJdL7SE6f2qfP
IQU4ScPm0Pv26PFgYsmRY5alS3o/1p25kCXu5H3KdjZ2It9AMzWmwhsCiGAV35ma
sneM0HCIXBq2DoP1OPKEppi7m4cUVEelg95QkZkdNBxdZr+Tlf7po9LXzHeySnxA
CjKql7J1fttu+mYsdb1ODfr2mm+SIgDaJ1SP0hOGBCvbtiVw6Kyoyz/lFYZxy9H/
4Yrq9ywyLZST5qkYFjgkfkXbKid5/wae3RTBJ1P4F0EBbx1VPjzCf/9jVGBZ5IqS
TIUgDegAua8gw8l+NqUkp6BH+4cFFlKZW2sHALb4nJY7SJIhLSNZSKcqWMfwLqqZ
y7Lebv6QXrCJWEapPe++GleYyAk5U+Wpn9I/Un7hJnNusuve6UQX1bmycBotEggj
23LTTqbpgFY3IDrGJPsYxtG8fg/WV/+dvomxbcmB63JY2MkKMpD0pOG8bdsFCg54
HruHhCiMhEdSFaWVbSSHmALukbRbi16wLKgZJ6aL4X3nEOW/QE3X6nclOM+/8YlO
+1KXkunfjZR8Eu5Qusqc3IK34fuHpdEkf6hd1f/OnyTYS7fXoKWtn7Kk57Y8OM6j
fJnr9wPmVrYQHnItrqGl5HHeAEkbk2Mqj5T+5CGTqDXJ3LGAv8z/Kmgb3EbKT/kS
gK4nqIbacHZ744A5Zo7ZZFtJqli2KQMol1fEo4PgXrevSMhjmhM35iHHDlqd0Ges
IAZlBh6g2YHEYKJaUyQ7UOiOrrZtdgyYZBIyJkh+vMF/vpN7IEVETgT61V/BO+1T
101rkMpH5bn7v9QiUqrNHP7qWS+qPf5+e3Uf3AX33tpcXpbAzpriPtFmf28Hs09y
EhUQ5mLLyiKHXqRi4uecoQb7V8BeNbeEJWgXfr9t4b15kdZOzn5Eb8ENQWIVMdhQ
c9bV/UzsJtUWGNRYin942RX6X6fzlOCwGdd4eayO05Tx6+f1N2I/jERgaZkNyKes
WCLORd7KbFqzQnaIAEnIzx04jws0NLzH7pTOAZlIk9YIg+kB/gsyj52EeVvmRXgX
1fqvUVNXRV3rN4CdcMvM1BjfnV71DLo2wlrskzm48kj6pE9Gaf9xy16sPP51amDt
EbCrD0GnAHSyhf6mseG+X/HNVnS5LPrARrh45NbfC3/8yPZ0+/fSscSJFM8OVcIj
K74lrfXB85zS/uS41ZyPYewFBO80yMxEwh1CXircw5mZPrsmhpJhpAfkNNBFl+fx
63x/QVRDgX0lJFiV5H49wbGumICmHmsSDZZTpjLzY/40zNz24UZyUWl2Iuk7gJNO
GaS1DtAy3YkeIufzuQFVUB+HPiTBgJfni36snTCbG4LuSVwCQ9NubV+Dsamf0xX9
sPv/ep/fdILoGqIL4DOs4hDQOKVxTBEBLDWng/z/t9BO7ODhtej58FiHKkrq+j1Z
tfxddd8xl6Gu+WPXLdqezqQvPJbZegw1shclOT6LpOloYhJkGhdSPHJfvQ6oNCF0
Dp4VCYtliFjTWj0l0DezFi6UZajzl930ExRJ6t5azMbL0iAxKiWjng6k5rI+1TZh
qd2s3uARsF9627NT7nBUrOy3bCnDq/SD/lU4WjTr6D0mgVM4qrbUUQgomtm/71B2
qrdqNRFhplnQEc1bT8bXZTTFx6uKYD9BTZHXX4c06AGrS4jMKVgGhBP+aZs5/TZ3
LUeMdXUmFbom1ZzALuU8keaAK8VuxPgGZ+p/0ehT3stAg0obbvaN1Featc8XUfaU
5FLlLWt5GvMHylRar4vsjZ4vnVsgftieKXfnbHCKiqdtAppOpsvfcmwDjWxVh8Eq
OO6mWfUMwbQTXTrXDv6woKDBxpIgarJ5t/eObb9pyOHcHju94FBgZFhyNMFeNbjc
Aii7LX5BYGORN442nq70NLc5jWZ/nAVf6xK1EZLeC1SX0m4PIlMaoErynbL7qzDD
owLbgFNcry2EKiurDMgNjP0rzsN3NsKErYVojUcC3B/M7pSCE/g+7tL3MjZsSRbx
lztTs1Z5GBzeoR9Pqy5gON+OqBkkuPN/oSsTHhaUksmFr+qc3SmXbEAQwVd5tpHF
gIhTRuXmaztaQu405+6Bh2+xJhOKHEOuRRvRtxIPcW+Bxp9ToiuI5+Sa4TjLsjnQ
izQ4gG5cjSHIbVSv56R9pWQ+6aT174YvpyiaSdwm7mrWsRDMrOOaGDl6YfNAGBfd
sspJ7WFbyfffw5H8kWsAdZ9Crzfx7vmr4z8jZBuz/+E0TQOnBkwuE35kQa/oawCp
Z1S1X/bb/yEfff3UQLv2yWlRf9ONx2PRRsNxq9DVLinuqG5PN9v60A2P5ryMDhyW
LI7X0TjtjBcd1QWOfZIof2jeWwDYFlqoGl+qd68hwy0EdLuWQcuPB2QMCvnEttF6
9GciN7+wGe4OZZ3qgqpDRD83KzaknoGHWTqxOadqhEQJDRrPaKlWpFoB8SU+IHSe
9IksYLjGQjjAIrc34a9T8UEvGGQzWCuRXHOqXD8jH4UAwr3X2JfyY39WoRq+GecG
0jKXGaFS1hQ+ZTtWG2T0EtqTenhv8sRZHtl246kSlzmDNY0BVUKdy/Ko86LHdxZJ
0mMsg4VtPlGlqnVgQdyB/7Ysdj87t2Z6Ldm0EWIOzPcFLzDs2fFSldCS7c3bYFaC
X1t9afez0JtskbhzrYbPwyOkK0+/KuvnyYMv5sNN/fe9Lyux2ZVcCrBrhpFnR/a3
6frUZjG6h2Cpq+sZBaHUlpim9LJrFhiSCKDHDxk86cUm48Yp+5maxuXteoSLpGWC
G/0rffDPkLnQ5BLYKzXcCrOjkxVUOrk+F21ZRkckPdeArl3HCHDW/vSk8d7cOKZO
7+qltqHaF0MudedGZH9iO+2LPnIEzzJNW2413jKFYr8Sb8u+q3qCF/8eWcURLRSh
VwSBxgcFkaecSAjwATmnpVVmP5IbOPQM9/joPFyK3k0sjqujTeyYrsACLOKCQNbE
gsyTn+TV4B5i6jJG/I7YmY7Fa6J129LSY7LtJlewf56j7xxVC5KuONekgFB+G1nu
7E5Wm/hRQwMoGvVsaUyn2WFbwjTThkJlUo/HY11bA/ynq/yd8mBduYh/aL1EEz61
EIyhafiMTDle7E/iu+GTSsyY+FbNK5rzvxaXWeQDgFuiIP/4CzULx6TbwkaxI/VH
7sBREdfGVS2j7nPCGlvkNvzs1hCNVwmz4FYkh6C9GJ4LSz50yYu7RB+3MUJltyMG
IrQHabTy4L7qVsrw+pxiFk6PjjLRENPToVJum9pepn7foUT8+uqzrAnQqYwS9aCk
iBLQzePRNLkS0xx42b3H3dkWcWTdWSaPOHaUFCkxrDxgwHvIMK1gwr2fK5j0tO9d
MEtvmGQVuG8i6W3c8p+l0HqqFgH6QwBlLYxfyyzh6v6aJJ7V5D0Dx8y8gPTFPgPu
IMb32Xc5VUjmXG+fJ2QiCcOfK8gVwTskwjkKU45HQ1UtaK50WfYP8VCtVAvSO9v0
AdGZlB9CvOb0XLKL5NiHZfo4q0akAk4stx7Hbe4Mm/d4vPip6hvDMYYLfCPixRs4
i/TWOcoeLGbxeXgQrGbsgQ7JBl1PDX+7mQU9xgT+4rf0a0zOsaTsl3tQ72gwB3vF
jfhzXGWM752PIRNrI3dhmMuCu9jowTPqRnzuZVWyWLqnIjv0Y7xCsTF9LtZQlZip
W0zvca83SoMiJklNaSrDpRMMwMBT3jm5gS3UPF4MeDhIHgUWY3YLgG1H2rbF73Cm
roXCBOGzMOdGW8+ibzOY17sXBBjpcUPCAmab2xz+8G9UHYeDRcbbSdVlpyMtKYuB
S/gXJ961bIZHl3QAD1c1aDwCLXSz0Rvf4gNvL/zdRRcKrG3VrF6LJPTZZXAkSfzO
tD3gFpI04TwDRYdginDuG4b/oboxVN+Buu8skz34Qw04NJa/Rzu17Jwdsf41FP5U
B0Cxd65wDwBz/z0TRsAyCAXC5t6uxqSS2xldwKBLJCecJYpzrPlSoGkhPAVBaXq0
Qwx384MsxXeugfucqqs8dTE1WztEDVX2etIuCi9adVujmq/5ofuqs8/t21foV1Tx
ANqduP7y+OQvVeQP15zYTVZEniRYZOHQAInD3Q7Nk0QF7I0MbpZqZzR0We1a8tcD
z3idWEPYiwgq5TyaM5dRE2NM575N55+7iIUZa3GbsGJjT34pLHxI4PVebv465qJI
Xga0z2MC9zNtfo9pC3mY++lsVrNmH44XkS96AWtqUtrTfyF0kakdCNkoXAOGHDZq
maQDnvBpZDFeNcABn/kHE1tP+3+5jNg3HqkttNHlL823AMfOWVbFjzZmwJNlS5He
AwXgdfqfolwFpNAp/crIsy2qG0e/E/9fYngAr11FFRvZRixWT52lRzQE7AnkSRvU
Tbnvt3Hx4FTbqsz3ZdwleIJ89ntWtPvOHOm2Y+oodjr1aGwn3Ea+Uu5L8VAnfwOX
iKOswDUmsQiq0wPS4NPDwRdAZrPBNvH57Lf3jFEpP/EiBElb2CdyZDkSszfuNdI+
95b7GTS5rIZ9gwF/5b61aPtAVAqoccjlQMV1JRXaTG8istJB0ggXYI6FOCBSWYjF
wxXHcwVCvMJO/R4zQiODfnK2lLgeFa/ieWtwknIJUQ5r2RQMSBpvXBS0fVaCgU1x
G9je9inIJolDiA2ja335sanOqg/n7LqsA6utNxpFI0tv43KOZGxXArO6is1PV4sC
o0kAAfOs05RRrM33CidyHEy+SyTy9spEtiuFafqNl6bDUgPHT/f6oTfQuZq3JKXC
hWa+CFjbErx9t8PBIxkIEYk9g9KMnQlDejn1OIQfo1csuodsEscBIMDn3pjFkG3q
WvUXG8u3pEbCW30RxNIP4wtvnMFMD83a4ChYyOU8WHWDGcLRDNr+JHQd6pLV9s1P
xalyuO+wXXuyuX/AQWlRafsmRQEV5ZWc9x2L62Yoh9sVlqkk0A/noC/QkX3azqiC
kNvRa9g5bREH7Mo0rer295pPkqM4CdsxZ7pG/elHhqAbh8G6TB9nIiLMATidQQNl
uo+MPMmcPx0hGX6gZ54O1Wbdfd3gIN7fyj6+vvjbnIGRCylUHaeEGraCZv36sZgO
D9CxzuuXVwn6nnXIJfwTgiyP7wa+XH26JGKpOB6kZu+lKm9mvuRJbmVItO51gw90
lzCUU6aTW/lLF5abV4npFaP1WXR6l3xbWN7/+y4NeOoeepBHG3kuc+WCmu31mddf
BDbWAdtpuDWiCq8RxujjDm1xF1mxEbVgZgxyPV1t8G6mE52daG0BJuYkox71kioW
+/ql6VM5QhMl9GsqEDy5HJsvd28h5DAynixo/R/jKh8zSj8KsZGbAHbgxsZV7b4Y
RCBMexsqTJhRsJpgnCTHmRS4bMTw7DyPaq41N1zSO6Zqwp0N1zg4C/MG4mRbWCMa
nHG69sfU2mpeVwBmj43bnDnmM8pyfcDRub/w2U1Xvs/uvRaefQ5vYIHiHF+lRuq8
Pv/3/z1XYUlnYkXAhPrBlWx8n1xnVjmxtb0GPPmjWdb9islrYLNo28t9dBoFKx0S
cLM3JOhGwdhRrQVZWZIe4VP8ZsB5KHvQQyaNuxl211K8Gg4gz6I/O09HYyjp9TCO
C5mhnIRMtJ1VhRgZeP7oGcZofwmS6gWjKfts9Ft0Aq1c07Iu4NMtCc3FXLG4AUp8
ZthGU5RbdF0+OV85lBrEtWTOrZokGSzOqQC20d+zi1J1SW8UX3AalgNw9xRjzPqs
BRkEqQGcQFqLdJupfBxPIjeal+A0E2pblH/ZVYooe0Z29PjvDdhFvO6d2JfmFtGR
hWFoE/vgER2WfF68hiu2VjNGXC4VXpynaFNJecWeXAl2wRS2nL+573CM3/wioAvp
leaIMaESdsNtTfRHMcEqVa9qozd+KRSb/lIaLpHZu9jC27E+q+BV9ChzySBkkGly
jXFDT8GJ+ww3OFkHNyXzcDUdAk5CFgT+SNKjrk5hbvR/XnbQW28yNw5xoT6wPy6S
7EvbNoIlfrKC5IbxhjTF92c1lEQQjgld02MHv/9gShALckZq1enWmwV6VoNQnSxW
FalzBlhgIjkoK5Jh3+D3Dv9CtU9uJG0/iOaVfXrfGEQWuAMd/lUdICU+fyyLyT7U
O+suz68YRSk3ELL1qB+Kh3U8XlLKzkFGdxYYjLKUMs+WqQu5rbVcqTcOhie2Vi1B
vNhFCUep4dQgEUHr1ilkFHw6gJ9xHn16egXe6uMC2cSLr3+3h5ksG0Y3rdzVYeAX
SoLMQIeptNNdzG0bqscM4KOO/LQVujZpT0U85o1aPn+rCKW6/MRdjD2DsNh88XME
xn4kuey9zNxlJTT2sATwPInRQebqS6EwZxJKn/4O79qzQohc8fEN0QgkOHwsgruC
IFUqQpt++kA6wsTOnR0q6A7XfyOmKlFd+EL3hmXmva1sibnP65KPxINBIT/nsJMQ
UC7qqv4+/DZ6aGFC1JBmMT1ACW3MEGvRw06IKN+5f3DvgUWrjtiu7FGiob7MsqIy
NUs4EXPfO4D3CRfyNhIjP0nXPIaz7SRkxWdWqyAJ1XFnOS6V/6B+GBOumxBcxhzq
1OZXKSCrHJgcKl8PVd3VY8V6dGU9IZJ681slA+sfPg4PTnH8TsswB8LTIsKy0zNW
Fq7afJ+rDvbfSElyoN0fiaz6sOEeIiHf9ajulQQmWM/ylb0g1xFDIDKRd/1rCjXM
oAd06WwapkuTTs3FilceS8D0aozcOSSc7+4tL0Qq7FJGiuxLBelp131JLLuoCdCg
oiO6eap+Q4xUPgV1lp8J++7+MP1682UA2+UPtgvGHUJCf5WrVoKEAnxTN/yGbEMp
9q1CAQ9iVoAX8EqhmYUcHTBxTvREpt1jY4wqf5qrU6wRpw2UCCOy18MAEV/4/vse
8/twKwKMtMSnXLHS38WDBLOOIJtVsMUklNREdvXKcsIpIOZEQUxcfmMzDTtUSi5z
5o7LWFNutWWCB3hFfcHUTskOmcCPn8TKf4mVU99qqWYNyuxS/RHavSn7onyJUPVu
YyN9ABENi1JYWsSXFF8GumCoIdyBVQ+NsHhrLY/BD1EUo/rWtRC330OVdUpq8H0u
TlqrjAP2uwXpkHlqHfTCmbHIe9UyCkTUBVZg/DbAV9MVt4KJG4hQ6yfNoZP/sTx4
lRFKd8EgMiGyHDa0cfUGNd+y3jytC8D01bUqribh9OlJEguoC+6zTZk/KIJPs5D5
WCejrwM4+WKe1DXKGix9/JQsghwQt/Z3VKtXw/D9li6D3+18jFvLAB4jvT0mpFMo
wvjMi+GzVsr6WdI79Yl6o+PsX0NegAX9nqdxLKtT83XUOuPF3+09tF+CNIlPH7RX
PLNuCyATzK4pdQnLpHpktWFL8zv/DSnH7tZvQNewKmuXhupi+VcBFC90XKcJdp07
vuNd/ut8zjjdzKOwBsOAdv2bdU0MGaQP6Cx55/k11t90yCT84dHuhk4lHpKNKTiz
ZdMbdxZhnTJKMYru4QTuff2gm7C7xHU5qnAx5ppQzp4ksgHuvSWYSLxE7k2JCa6U
ZvoeEordPVVRul59NTgcgJkIcUIFLYvNS3C4ucR6+CGnGgDS4e7T2WhA3fqZmlde
zX3xolwRCbrqxT3Qx1Eg8KE7NoqdGHhaSTWYsENaDcHZWnbTTa7VvTZMOtjxj4SZ
EXiR2SkxnuvA6xLc1Pq+xdjT0OJwok38iwBgngSE016KAS+b6laoXiSpnAwI+jBc
c9j5yw8ZQuVEmqqXVlaORxGnJY3gGJtrTYFEyiiFyeGK1JOlTF+fCQ2haD+3Y2yS
g0gHSsSY0TmeqisuypsAxucaDz22F5vfwCnAJN+7uaFZhXxL4aC41xsU4deCYyrb
ZFkE4hlu9sHSKjDwn7htjdZDJxfMrf7P995d95gBPqwQQ6bFyvgGM3ZALGTvmmBw
1UHrUcn4WfR6hejz2eK6awLWGaDmRhuKdc8Bn1PuOj6Ie96TpdDuY7lECc/sWihE
Q4IKwOIwViuAAUTDJtHK+IKSvM1dQ3GeHDVKoS9OSyW+X3+qDcQjTxnktvKbZPRT
+5asI9ltJdV7dQRN4IjhekwjdrrASF5IfJ3CJdxAPxM55aVOZgbSjXmU5sL2m41F
dlsHOc46I07AP3ruaC6wOZZmoKxGhqpLrbJw+U00rxYI+lic4MjOlwuhyncM6hs8
cNg5UDs5gzjO+FLrYh2e1QMdEeI22Ocn9EWsspd4P0JWi0gIrOCUMvDBlK+uJPKg
3uClwiDFLqFeLGhlQIgg8Mj3kHg6mZLK0GNtWxR8YOdbFMkOJmJoUlwgTmWgA5fV
3sr7ujglXRpwRH0RqokwqIL6RdCiVZtKjWkmsnTVumXAJO+WBCGVnMXinftUP7dE
as75QN6eKHiR9bQaLYDTx+0+md1oFnSlNcrMxsjuOPUYZ6OyKfHJ95/1P9XKD1wZ
5s6HLpYR6mv5wxt5DAjpPNS9rBuvdNJWxEmj6M8pzP86rfii0fEzFmvA2DnBMx0t
ZGzGTn6bhRkrpyGy15rCnxFyD6OsQz6WSgKTOcgIqGhZdrTnBsjA704lnKVM2OHh
ssrCBELOxW6BLp6N2aYmSB/gT5r3LUd5hd/OAGTTz9tBkd8bTradvZr8mkcNrRV+
i7Cx8U36fGEJjhTYK8Qtc1asBsWi6BAILViUPCMpfaLP07kaI3HpqS8lqfXKE+Wn
+n4Gf+7bDi8nHGgvWX4k51XbXxSoUpsv5CdLYdhJm9ySDD2kSsSxsGaDrzKghmBa
5+eoMCqzhjKi8iPYS/ADUnVVRVour5ywpsAvhCZIgqb8vWQn/UXtco/MvKrzY+7Z
NHOoCC58r9HC7JYFiT4BOjYw4gsf4dZkoWDVZXcN1ESqmWkL1mHb++eaJigtdI5z
uFH+0UpwJMXocF1p38WP7VjCqfH1yxlUzWVjcgSmYpsIGgYrpO5jCcEno+WZ6N4K
U2A1tRVx4SIw7qdzpmQ7Gr7Ue5LnipGFd0Zg/MA79LUTsc2ZoL0Mh5KFMZjS6hd2
KSh6lISz4PeaMtSsd5sbYm74RT7Q0BWdugnpibw7NMd9O6YdjTKOTTSQTpgP0ZpQ
vhnQi/QSgnteKqYWLx51yM8f6hZ/erZaQ4VkLShTn0Of43Jjue2lF+w4kqh5my+i
T6STfLWqI/X/FFj9mTymehadmpV4xiBKjjClH4tv27ak1V5z9Ceh/qC3rZXzUwVw
V5ICAXUKpufD/j82vec+/fzZR70L8nlUxFkkeMYAX1B0enBCqT+r8KeuubZ3r7Oy
eviMgh0OFTXy6CLMCG6iwlqDO6FLFPmaRNnzl135IBSbmcY7IzJdAck+qRRRQaSy
W6MGD9+waMtHfMm1NVoEoHc+vgLRqoNYfxA3NHoUbJ4aTqtdOjSpz7YjQOdMV3Ep
CbCrPiwzLbYWKlFHpsuzJQK3CVbMlXHelNJwY52c4zxVV8IA66/eAj1dsxnTzvXz
MoczT6Ob3wYzeyn6IbKHlNNeLBCop6Q+dTrLGF0E0eleONxVSJv+9RpuNIUmlELx
cj/0gKty0TpWyB4Cw/i7R+UoVKGJwRGHcFrGMpyloY5kHKiFEYZIbrjgkiB3nm5a
Eni6RE2Dyi0Y8cSjosNykBqDZROPyTKMJkcwTaIPBGhqXIniCD2atLDpiQKBBmw9
ksM3UEszqxijdxf4+i5JJY8jN3MBknr/Sqx5PBprVqS6/I9e7is1ZQFW0WeVgZma
rC75++Wz5ufLzlhOQUgl75PVlZVCr6H8eRJ3DrDvEqG1obbH80aP3NFdxK/U4UxP
zHLwT928RBrUFFpuNZy7KezgniQ2tEoodxXp3M0bQR44WSHp44f04e4mu/nOtbn+
POU2aZctK0CdfNMvMp6boQ7c9eJOgxcO1Tc6bskPWdQNEPCGUb9M71hi2XXF9QDz
WnIc5esN5z8xlIA/5SVXtHWNwo+N/YvEgviXXNEwdCRhH1eFyrazbvPDg6ukWPbi
0vtEPlozlxvsieO9Y9DQybr2SmqWLOY7rrhqy5tXJoFb91yJPKNm9+0cGAjl/nTC
uPm84Ex+/vUEON0EzI2qz57tysFqpDwg9MILjmxxxW1E23eSGWnAtUuGGod3pxYO
1LnpMkZlvFxOumPhJea9TLiTpb6G8FBcKRpc3PaPzMe1+4ZJHi5YL+1dadTzIjCN
w2MyqBP3ZajCv5qtF8iDv0x41hgP/GSgpveL7cOrlF1Ag35x64ob0mgcgdRxtMVw
QxI6CCpIb7jxCKzhu5ufN27y2nN0W0KLNgWVnUtrgXsF32/fUSIsfcbImTCPfLkk
57NfWAvpzDwup0uZzbkVoLy18KUxzGriFk9VK3X7xDH/91SNxEVQkUoiak36s+iA
/vb4+6Y+YMQDyXYhLYT1ROqKWAZZmXrNO6sONCfA6n6yJZ1X/xnej+yEZGPWTHj6
8TQGRXmo65ClF6FxYzX5w6QZAt4/i1jiJTuk8YHFmlQ8HKwG8zLPd48VbCOSjkyF
k1I9ArsX1mdQ2+Sqf4VY9zwIHb2X9JzEN7tQP8CEyIYhs+zP78+JkTlccGMVY/br
2+Gm01Daczt4LLgEIyi6BNYVleCZiJysR0M8gvKEs3pmwxK8oTmf68M7dn69c5Li
Vzmki5CFAk8s/9NAwbb2WPOi3ugN8d92tviH0bxl9uiOJ/LccPy9w3HLwViswESK
UWWcNMXP8A13fhCFNhMNB83dEE4IhI+0iAGDFTvluUPCphViTHeI0Cqdo2t6mybO
T/1xXsE3Su/q6xLHTTm5J/ejV+/uwrNfuJ2qwBtQUZqJV12o9/WF+Zm3FtfP4Iqb
WBjjLS3ByQRRqEoozTmI+GLy2tGqxLoYJz0x4CcEAfABMolWntsK9A4t4Aw+bpi2
6087Lj4ltpxZPi7JwcOVXQP9WONW+hVuzsSs6KWu6+Qhe7v/7GLI6MFKKUsqiicv
uvWcuf3DWwEIQPU9yQYHKT6GwW/5CJLldgj7KZGCB8bPa7CE0csYuDnH0Iv+ARQE
UuiHPmc/O1fjiAVeCtJcYOQjt56IvchCRomlD73kQGLRuQ70VNR+21Sebikv9YUy
aUxjJqBhHEzwqsRcpMk4GKYMopDqDZf7QnJXr4qkHduMj5QS32pq9D7LHyj32vLC
FLAbMhNifOhBnmdIZdScgynAjsMdMKn8kbxU4pPL2oRenW5tNTnHQkxYUf2ViPIN
TeyOFbVSOXzlYkpCpewri2n9gVpmY43O4Kfc+C8VsiY/BqLF86EbkhDetHGPpqvm
mVODDQ6O7pLf3KwhS3ydykttNILUbn9U2USFOp7LwPzwd/5gcNIfgTPwk+qmh6l1
oqquSFYTTaFd4SgtQ16TWk4i2nAs9LX75wE3AUBuaHV/UbNIcRnvNdo+Zbr6kEBo
bPg7Y9uTg/e89LKDl0dr8tf/hdE2gTFdF6WZwtJti0bfzPDJO59qvebfNggSBSiM
YntZxQMQCQm/lngVQeNUiY1Hmgi7x6QVdcLYUSIRLbT5aOTxYPGiQswd0ORn9Xlz
+hVx+qe7/C02jjUiEOAkOfV2eF29gLG+B2s0PHv9ttbVIUoNuiV2xahwOOWiIK8F
6i9j6gp6AZu3Qj97qs0xrv0UQyQUhH7J5GBedQkyqag06y8d70e+UtqNRe664S4j
LzwOAjV//eVi+sLF5RbAagukWtfgutkX0EIT/oMfu7q6vLmQRjkDfthpxI3yws58
hCaH2Zd+0rpFKGez13Ms5mIufQwV/qd0HfzEMuVGXwNrwHteBYw7VrKvFtvnmKUu
7xEf8JIybGHQfh4W+6mKcTaEIaxk2ieZFTtbsiXUMWZQr+TrrvYDcLOem8uerSY3
sNpdpNJmhgkvNSVlU6VAvFlLSsw/zSYHV13bHXzcIg8cCF/i8C6vqAtuIZ/C/hou
3Ghpe0GPJG3fMAArAsxRU5LDNNW0Fkj+MtK/mIydwpb+tuYGjt9DkbP36LUa6XQe
zt+KogXjg+k3fXRmVysIe281fI+ftHLfU+C8KtNdK9y+HVOdrj3KYiTgRzO+ftIA
6uAMQQnUUJojhpukqGIaoocjBnscBVLX6WZO1Gdx0/eCUdGFyuF/REeUFCPSD7nO
vGfsOJiMHaFTBOgj9ofnNDskmjeMy+d9WS7blSkWgHsDYKnzEduZZC5zGwsxvqfq
BZSuvRUAWsDm7zj00wTG0NcyxtaxYk+vEywhzn3W9Y0DlYU+KVELlEQPIjDbcnyy
X+Zur9SdLEmPxZw1xW47jH9PCIys4q9dRzMg5tvT/wXvrBWPe/MUpIFBWGxfL6w4
jSG38Q154LHX0cxFu3ae6hojCF3EWTFBPBDdXjbIS6hFBxkGbfIDzGwEbr34QPJf
K5Jw6hylp6r3OaX+u6e7aa+4BVc/Nj0iv+07UGXjv6NiE6WnCK0St/BXZldmuPA1
++LSES0JSEJJGSL7w7wpPSluQmOkrkHYzsv8dBniFh787u5sNGZaLUdGfyizKGHr
8slQlE7Hdr5oP0tWahjCVbf15hBv1fmbPl3g35l4coEYrvRCvVVVZ1aGapcw8JFO
qjS94rE34ofBMc8qgXxeWq45QtHSpjHzD5dMYBWmf7BgDslSoAJSLw5YAVBYknn9
fGjOxFlw39D5zbNS0YnP+izptSjuWXlq9kFXVKktcD/TrU5pMriPJNqDdjz5io2i
x8c64pkiqWyP7Zdc5UrAxuVqCpDH3QYeLaHiWY7v3GmtfspU4Nnq4S4s87bJFcM5
N/qTmXfUV0l2/aKRyZEiDN09WuhTA8WsqeSwVK08YgsVjjZoMPjSb7zuqwOUUafJ
aF7wXKdIeEO3pvVH813hKMzlXT4Csxm848VmExum0NN0j5YNxFQCWZQKrPlsm4pP
jJ/KgZ1e0BKZ+J/S5ldZ3AjSuSjT+C6RFE5M038A/I+UMAPXy3Ji47ZEHz1ikBv/
ohP5eNLvFdANrjT73awkLgJuxidZyaXFxSRzd7yvH48R9im4cbmmEsxG//NzxsMX
BIDKXuPbwcwP+63IHVp2I7wf+zrjArZLMVoTeHRP9mVN54n07etTHhkrrT9eQlH7
92HCy3IQWf+CTvHL4iduwzhIICJJ9Gwy0JaAxlsxDxhmHd29YPVvdaREzGB/XFt/
B3xb9DCAl1KJKpuS+h04Rg7TRxPGoDLiAHIichY7dViRFTip8Efor6CNkydm7Qvg
JPtDxJ/IpNFQj/ToxOLRewLmI3a9KAvDfxKoPBB2yxbtruw6pWnQZ+guq/rJCfI5
fyJU4gaxIqim4VtMmUqfQol4GiHym61YOXwccIdT/BoO7idk4yhofgBXMrC8J6lU
jTTf8tio8C9q4NB7fCiCGacKy9a6l4KR9zx5uqndZSQeIpexOiqCUEiVQDmaqrB4
ko5tymwog06SrqWrXcxn1sQn9N1/JniVp45PuzxN5So1uIGCTW3bM6P31W1rFYBf
HhRy25MSRnPr2VWvrxNWy101tRn4QsdsRGgi/KPxOzY1oZ4jCdYO5sa+xX7PbOq5
mN5WtE2xjNmjz4KpFEr29txyPugLNdC2ChnzGiZJPw1oPHDOP/qVpwRgrH9rbGsI
sHwKweCfLR9Ay/CIUOwovxnvjQ7uhgdg1sE/R3RvHJYZTXZ3LbNyCvDSJpX26Ki0
xuWR8CoDaFwUqxT6EhyYTJQyWU22vJ/dnkG/iFx8D3Yr1gKj7Um1OTUaYwSWqcxy
BrryZdWH0lAiZ/8VOo6VkKtHa4RHL7hq+I+ouLxmDsYxymviiMVZFohGYkhCd3G1
8mpNV5uXdzMqhwa68jSsgkMpSDH2k7fNvoQZJ+KJPbKNKOL2R1wCXeTM2ZvuNFS1
dTLZjB18JlKTKih0htyIHRbVs+DbrtXaMOUBJij3m5k2Ab5OSxVCrOy/4JkfIk79
55ihNrQSVdgtIbgPEmekji8TSAU6dizJ/YdkAzWOjZK0v0Ndl9+7U+e7spr6nnsK
UI9yuhZo/h+u7uwypJSIdB/50kJZ8gX7gxi5XOxJ31nGzSsRa/HSqt9C79hlE+Xp
c5GRR19cLzF/z1j0p+HsKcmDhs0NLMWPWCYHnjVpUPrN2NO2fM1Kx0yuB6mzfgly
P3yXuG543PQSdMODFLlgcloHHu0ZuiwprREDMGTV58qs2abfEDxHqOD/i2/HZYNh
Bh8TUNH1abLdDcYJ/CvZmuZSLMj+NgMTqq21+vNQpTrDDV+zid/LzoCcJeYyz1cp
OTSd4Tu+tgb/yafrxZ8vXfmQTFNTSLHCnQjdY6ffsFQ1YeD0PnEhPKMHaPBjyY3n
yd9EJcxsNsYjy1Fxw+oRqurPwYzpcEdaFsGQUtiOdAAYVfMzdy1Z6jt6nxCELdyK
PI4l4S0pEBm5KF+jbKoOI6Ire7ul8qFnnS0OPHk3N/GI4UBCklZtc9kfJ4GbgmJE
vDn7wt36WuJMydoM/bVeRuEeNa8yp7fB+sSUM9UCur4siBQ7sF/lFnI5q5CfhLxe
qA3B+4bYQGJKa3jiaIdwQHFoeuLF5DJg4T4ddiFaQDKzFp29QmXgU6Yl/vApqGNX
xrzPnyvmwm13ll3UdCtDKe12dcBjdA6puFKYPeur8wMGY+hS6fSDX57X5neg5bjk
Yoc5XzoRmjezipygGCwNMcIbO/qpRn3wXU5cJUwZWbqGTCdep0EASa3AgtbLI5T6
ixoxBfMDEtE/BxIhxirT8P5hZ3ywbVyIU2gfrDYZoHzQOu3ScTYwPL9dKKL5ZCR9
bbsnZAPGfLJmJQG8UUWi9bET1hMIU+99mxZ9aqdawjDxvKM6Dkbps9B+m8AnXwHX
j29BG+mCuzKNbKCEi4TgUCtm4bKfhhvpNohTe4s5BcsjtSOwUDa8sPTc620hzRkE
SFs1IsgOnX0ftFAo8RdSahpy0PQMB/U974wffho8HxIJURuB4He8WeXtJuEBlTcm
QokaBHhJbBMSl76ktprPIUK69RjUsXJ68xbhT4sa7U0TAdNFu7I/XTuRLajHag3M
EmaUktTUgVd84Bv+UbeFvHWu901I4IYMzQihdZXYlC8f5ko5vXX9aJJ8kFWqNAey
pjSxYpqQW6XVQ28lV+JB9W76wgnKhYXvAqLT2BrznYhu0RjSmaULciCPFTtLB2dg
ArxWHPuXGTl95Ylq1fp+8Y1bvzveM2sgvXP/wP7CZ8Nc3FcUuDBORatiHNvHpCtq
uONNWVZPzt4JOy8oAvAxMTloxwtymHHr2L2D3R5RCzL2k+DjQqYSleyG5j5cDYIP
rcHhAmCo7MKeZmSpiIcdBWLrlSP/E8cdquy356f/P9cqp9WlhZx5fOHpUnsMmsCk
3aiakgvKNuAPtm0jvLjgs5Oo0NuuX1QBJnmInBbzidbUg0Kt7rcQ6vwv0Ti4Vcoa
9VZACSBkWaVgUVB1tXTe+LZTPNCzPr1N2c4FXW4SovgUseJiF2MzdbGE5U5W3/w+
eY9cHMRai0q7PTVDUN3jD2LjfTV/C9WriKgnvSFkkV1TxG7c/3gFSGMeNxSZOOAf
/YPVHQq22DA6oljLj4DHrPzr7aEIhfgIi8L1rn43/iiYu5IpTIUBvQruWCQTY0zI
Cr09JhplJLoaevhfvejbgY70A4nX7NDxu6a2GJPUZ2kTk1w5j3t4CnkAlXdh5wlM
Tg6YVNj2ask72RbBDT45amdy2JDXd5rMEGo0BQzOoUOVERHqThNsGPBrUTEBUzAL
dZxkNDSUR2TAJBH2PWa0FaHywj/EGZ+6JpcgYNG8RizcfzagIIoC9Aon9l7nvyTI
CsLL4XgUkOTU47Vn+Fh5WS46g6iD4UlbMsUEvrSkkh05FybHo25S43howc5IqYJB
PSPz67y59umGZl+KYi8WfGl+5mN7VbZujqgm53K/j4//j3kLCpZtR9N7qpciiqUC
vbyqtp7gnFD7cz5QJH1jhmXdRMtUNoHivE70HOM8EpfdbQB8Djy+5yDCH/9t6uR4
ITB1S6zaz5yQN3ngirQHRh/SZMmpllDyy2cIauiA8VYwSsVp9ay6iVZAPYyI8E4A
R9lQ5zzfj2U5UkQx1zvuswQYnqXp3UWluglKXb/4v9DO/WmPyAnb3F+fpxRk4uJ/
SUjPWxgxsIne+VIoBhgOMM1OafsH9J8pL0qEoG60DHqxpmcSrJGo/JrH3mue5CIR
EOPFE9kzceUOjdW4BMbtJGMvu+wctpb5w/lnkQLj8pkxxMWp7KSRHELBDLkyVtJW
Afqh6uFOwisu4MkDMkKAuVbVOTYxDhsNVSW1HAz4dqO4L7xBLCXLwtBuSTpGrEUT
DXJ8tAeyWOvKE5UdIqbmg+/LtL/MQKkVi1UF9fjzomm0rqUpPIiEjtFVHuILWIo2
eDBlYng5XjGzqW9qnRv9Us4r+nBD+dv3KIKLBF/lL8bTwBdGkK1HIV09jCOY+FQF
pxvmaGp/7mH9g1CmQgRx5zbP/v5/r1UIjn1cgXjv8DXWn/qUcMUXq5eCYjsNt9jP
8+0l+t55VxCUrwyFkJzi45Tg5Uo0cfpDuC5HKS5wNAA1ogPtoZpqjt4ZtORSaPGR
mFySKmqCsue1JJEjfVgKXln5YDcPNGISWg2i1RXHOMYKH9wjybY3UcP4aYL0IwSa
fPc23x7OONXj4Gc845ajIkC4x2BIpUOTlHA6LoEREv/EMfii93pMkyTyGszfNuPf
4Ab2yWdZNiuFKw4oHClm+WCX3CjDdwibnK+s9FKgm+ZnCiklPoCOwuKcsPwXAASt
iYDtMnT9mB3Si/5VkH0OfzuzsctAEx6VPnv3vjBlnUZ0aIYS+tH+PGKnGxGFpvQZ
3JyqOjt6pnb7b2mga/uGGKy4CX+z7wBMVsReJFb0R9x7nIQccKmRjxsUwG2nQtoX
XTu8AG2qZDkJKVyirE6MlHE621nvYrP3CGLsw522GA0UKxfS9I8zVgHdqB+0WuD0
/IS2wTczSO02K8Zk+ZdpSHnb6biXzSneiH6ORAY6qTdgeHvziHbelo/Fq8rvcuGF
g8y6oUIqfPuCEn2aAh52U7OGUo8+ps9uQDYSZBtcsomqjL5zV16xxp9QdRq5jWwE
x5l2/+OcBYmmhFgUdKeDuDN7FNwOtrFia+UXh1O28THqAAj1sNLJG6dSA4M6Dqd0
BRJQF5SK67IlaLF7sQxg51y+KeyFOrnOm6Rvnx2NIFCN4zqMC/cNbrG46MOJi31S
TdztufPL5Uw/6BEndIF5WRUQaEozvuDok+4SoXgKm9k3I2mGEFjKQDkNhsbhxV/N
xVZ+EcIp3VChEsp4dZ8A9hRTYkhYb5GE5ZBLktpSLQevDVP44x11c2lqR80Fg5Ig
Z1KCNXV45GG61Z9JLwmYvhFf/GCFNugaHka6DdGlcGWYBpDFZCnQxL9bJGTp6ZT/
XjIQbw1QqOXW5hl9Bfb46qd7RmNUTA4RIMkrzaxIrq5pH4jONmZ2xMb10UFKG4dm
QfGmb5Mr6vZJ1U2/en4DfeJWi1X552u8CXK7rv4c+lviIecjDRF+yl96Y4/4DffG
v//D56PTMAE6moAy/VBJT+RBwBB+ewmBX2eobNRbrMjng6vRCVybEWze3LeiUF0g
9IqGRhjshKYjTBmaT1KLbBJCeXle6scdbla9lmiNny9TsVZugLu/RcDgkjH+pgVq
ethoWp3+KfxO3VvqRQNKHpEAtQlqeInbc87AL4KJdFMaHN3ZtIwWhNFxXgDw7R/9
I1Mema1Hf+zcQnXf0a9JsCMphDTxAsKEhGaX7ac9sKN/nzNuRGRhRAN+N3yp2nxS
Q74iDSdyWf73KQJ6MbQGRXNKxzGJ0tbfFmZ19AKGjpRy4yS5E6UJIRrV+OnJLGGG
lJEoOffe8CMMgmtCEEf6zYDYtNgOhxGW/zUD1CScBpzAW/qWutMeN1d8bsMSG+HX
hM30w6HCy0DvIrS0ZnUTUuWS5ZYKpfCZ7VgKw0Uu5q/H2SpEAJhWSaCXgYTBkdj1
y7tF53BrStGkiobCE5wswHkPp215HfGkQTDjQiTrYT7DX7XZxOu7+yZsI727Cv1P
KarEE97IrPGfc8qPcx5IviSmu525swcME0GNBSHw/+UreH1akRXl5rGb/2OMHWIn
Hk77zgTjSJJe+RDQIqfgLZQKU7aQlZ08T3MCZ6qRnH2g5SIcwuSr/fIYQoa5gusb
3vZH2xnQFsqX1NbRoloQEcQcgqCewd09p8fYFjd3MDjFq3ULi8ND7t9QWpdRLi4C
8NFm0I588axF2ZMGQNzyjQ1pYZ96whi5H7BuufuNFJmbaof0mODPGXhH21YvyDXz
phhfJfF1kr/x74ut4M9Dfenet85wNvMrqYC0tzOyiJ9YhTVrGL1y+7Y46bbJdKQ4
MYfiEcopUYyVNu0PMMgyq4xOdPMRE4mZ5tuSReXOy9W8djw1Pp0ynFdKLJg4O9vZ
AQ+wPFzPXbhq/MJBhUEH3MEU/qPn6+DuMOG64MZ9fMsK14d0h+YlhD9GiVnPLloH
DfCzffW4JjkoRrtZcjS510n3D3hkBtSXm0+sqzLt+N5f5nhcb58pG4cywASehqWl
jiHtM/P38v58kPOD9TvDAQYIRvPzrUB8BFNZnCNjN3ZKn4zv8G29bwN7QvNuwvqd
A5BOwWAeodG2hdjrllOtTw0+mIqsgR7qmcRw1wq+An8rwTCo8CbA1UQiJyLAqVvd
HEWFAI8yvbvLCEOueMdgKK6wcE2TCYO5CJfQuJyxCc+a6tlKZomniS06x/RD4n//
lMKVAqUoJc3wMJMkOzHOeCsnZcKgwuWzIGLiesmBGSqeKFOTtTYLiR1vrWbM53co
DkNjIR2DBNbRHRa2oy6BEc7fDr/jg76jYmXLuQEEzCJhZ9UWVZ7QtklF2k5nuMNc
F6sYAz1KO+/pYObZ823uHppSVM8r07NVo9cR7oBJ5I31NuVS0EgIVeBG+ENpeKLr
MlQqKLZ/MqESEXw3QQ0t9gxToi1hpsCnRPQsEWopIPA25iGfCoifaC51xUJAQ5/P
+Yzefk7+J4vWhK8frR/BgWs7z6qk7MHGXtgb1gCoOc1On8ffyQzW51eVrMnkahf+
pBhTvjWOT6cp6HCT2lKuYf7YZy/la7t4pUiBoydcSKGo1f66LdovFyFZAM0csCHw
kOgFosTMsXzIm8BzN6o3v++yh6xgvRhy/gmNOw1WpUA/38Lnu85DmkjQeUylnzwS
TXFN3+If38HVVldIuSiGQBJH+XKWehKu/QEQ4Iq1kr3Iz3Vpbb2y9lwPsOyILvBo
84lz1WV2ILYCxMV/nPAF//FMUitTksmACYWDEBt00E1rAIWL83/TQLOMfTewgT7C
UCOjg2GXdKCi+is11bydcE43rXU2G5i0rmqWr3FyGw8q83vyjukbSyo/gVoIySNl
40NnpuVOOAmmPNxTsqT+yMCLk90GnkwVKUKCDG7mYeYAn9egnSp9mNpjWhMZyx8Z
jn5z94KA2V2iLQUf4QQKEilukzSF1FILzUIliNgT/75Ly0kaVJzYWURVugiPt0dP
bRXcNR+1FdN5iIg4FfM0bms/NIgwWePrcTUU9z7ApGcVxyY3UB/f2hSrovkPASGF
RiWbTUQaWG/uSmNTtCEXyGi9GzPaWYBm2StLZbP9aV+4pe1lWW0vPOal5SxRum8d
au1sd9kAN/vdcKK90nkkDolyFBK4pbjpaGv87N3SPK81B7FQARo9ieJ3Lq6QMM+R
nb8ae7nkKbU8k+r37UdKYIhOSIuNyW0UWRhIN5HtHS6qDT3h9nyfmBn+O6yuuGYK
piLN4hcRPL7HD42wnzr7bXBHxbao8rfQQiSr+88Fk2ATRpVD47NWlTmkTmK/5R03
SB+lS7tmHuH4Zhq4rITJBVtPTluQpGmXPgKcl0Zlz5dgAEo/+UChKVx6ZdAOowQM
8PO0RQ7EBXwq1hLYj5BG9XcNrTTXV5nZ3pcOvaYNOSX/Tj+2+aSTvi9fH8r8Bnus
Rtfjn93CJpR+K/7R19JM35WYA3rBXc1kaYwiJpm72Upy3HQN7v1u0ovV/a6crsBq
CFgwGuWBB5YPv2NLSjB4lqSAlBz+6Xiwlmb0aNtXN5shl7AiDLcOr5KdAay2BwPV
dlCZ8ZnoymUdTKgaxZy922kEMAj1E9rChPiAh5cbUiFkTGcybKHhwgn0/JYRUkN1
HQRUWwr2tlrnbumWi/AlBhq6t6hmDcpDvvI465aMn4hMuC+IlhCOPZB14eZCQuxI
kmajdrYaw7iPEr9pTdjzvbj+mA31HVtY8Nn5qfXKnqV6e4WB9L9p4A6Ek8uJnBUY
Cv37jpM0u8IdjhwHOUkqk7DYQ3BENtuyGHYkhsaDWEb8BIMiKIA4LgWkMk3RbQSp
EZlgSTF9rmCnpGwA+nCMP9Gn0c6NFXZvpQ7LasEQ3Ymkx9wAbN84Yk7yszRtb9jg
2O9WRTKPJMeZV9pI5ZPjek3/EbiAAmzonw9kOtKMcHC1GZgmHAxihO1eRxpCPm9r
72IMt+7kCT5ABEzPuQ4ax7BbYGYS2HDs/DHD7NcDB9HkErhY9hx5l8T/35WaeY4B
L0Ml/TOaZsPdoW6qimsjFmIUaSIbTg/5ZlXwdLMbweq2FW6+Ba8jI2rglp4UXNnF
chNSkghezu9xmZWBsvLVh3HU60/dJFPqNRvEY5/XBh4S8ndB8Ik8z+Y4Fa8en21L
lnYVMm81lhlYCZcEVvACSXY/A19mdMlVcHyTe7VtQGvRJ07xUcxaBe3wVRma8J0Q
bA4Z8WYcfvXKCP8F+4uIo5aBqo4Z9Ax2NcwUe5BS77h/IFJDF/h//YmXRs2TbMXi
PcfIezN1CBEBPVGN4mNg4hSxAhNVhdkjBLfOBgF7u5eXMO5V4GuHdTD0mxpHhaDt
cyk1gl5Bx1MWYdXXtQuagXaJrfe9DfcUmnkG9KPhd5kXamxL5kmYQSW+rMvhu0lo
oCyeRVdUDz5XZXQYxnHdDtckem9Siz1UiV/rrOHX8KGiJNNWp+YiogC4sg0ajuCy
QA3ru8DdxSFF5bPNn3qdwjFCtOuFsLqcRU1feHG+YbIlbEj/hY5DPZxjblyFKEhG
lC2UZsMsgPi3MuvwR00mEAItTNg+lHodw7UgTKU9t4Q0RRbYCOoYYvlede3PpIP1
Ck8eKFbO4utlTguKiObOozU7n7BFNTcFB2dPJBttbW0z2lu1HcRBNQ/9GOHdXCMJ
FVx/CmbrrNqrklvp0kA+NNLV93+ZnrNz/dKL59EHgmvyT2NSpZYU8Qx9WXCi6y2V
4UeAZ9BItTVxgevg/ZN5v6YXAanEHTEJJpAm77BWofZseOY8Br41hNaXQeU/amc3
zoWpjPFUOvX/9p9G8L30IoPbBORMUnSqrf1DnvH6ZOdkx/YRCLgtoeVscHMPwG+v
brycUvBT4jDTV9V4kNs3yQD0YE6a4tGPDrZ5cq4Z3Rv0kI4cVUTdr6i+KKrmmoKf
J2HIld2SpVnsOETeEk6vAOaWzHznLFeZrhmgn5T/ZYM53aCCOqkQ08buZXqYQnhi
bnfE3StKX2BZJhCFZSAAaKOoGFLp00nZ2q1dpbzhh/NevkBDml+tCXdfoS4mZeX0
dmXO7aSxX3lLNGzqdE5VUwlRpcs7tk5Rh/m2xWxDK8uQl57NfCculYayFlcq5eBX
ESEmH0n1e3c9HAgqq2vjYdWf73NLRFd1YPyGbRzNnSyKxywNdIw7KF+S1//hRVR4
PCG4JNSt9BUQXTfdyxaC3wzk1Pqh6i3SoGPMiadedYx5D8Pox0fnlAekP4ZdE2V2
sJn56z5FR4KsbBvB5ZDQ4r+XwbZL2Yu7t25zG7vvUKnzMar5LqpeKUeMZR/29Aj6
Qx48hFYjogYY8H09wwNPLacjWY8Hdx7f7paGFXZlht3uc2J/lLcz0ZGu6McguCap
dcrZyCoOxC330/sKuD2ojl/j48ixr05G3ZPpb+DqaVJqoGLJC6IlyMRKfVXmHvDt
uf8pYT7x13zvodBI/2GhR0elY3hp5xk7ix2jldeaX1CwngukC6zkf3U+WQb9t+4L
MlJIIv7pBkeiMChHVk9MRs6JCHdbATn1NHyXn5YR0Er2Xj1YeWq1bj1CurccCjzx
aOGAL66pmuwq5C7Je3EY/GRAMJzJxGCgz+yVMB/JFR8GnHJ013xzN9rJngUynjx2
x8E5QonmZixmChEPO2V8cj0TILunrPYKFlS6VqL2HKld/zc+ZNuQRRWP5WCJaNT+
VypcUIUIFbWfYvINH0VWezhPzGp3n2jVX5uQx1TAlAN8Xq3G/2Pd2gFsjJey+6Pn
FCSGskmF6Wu6xrHAYbYqVteD5iU82EjHmfQcdjrOS4pCDcqoD3kJexo7rZJBA81n
nTn+ZYu3Ti0o3nqJvyL1TB3HDLOjj3yWYnhXzkhLt+Shk6lBmhxGhzxvlGWo4Iwj
/wc9dskM7RvsNN8h7fGXy7qznOvSs+TqK9S9hjCl3xcqISZXfRBTL+GogNI1vVRl
SFZZ50K8WnMELq+5pbViaFofDqY3JRoko9ygy6W41RAKwFtXt8dPltokR+zhuz/7
nXo3wMQ5w/wHpLAeC+956xaAn/sN4BhY7pRU6kkeHo8qCsIomYcUIfb0y2kuukVJ
lVPbnoalFSDZ9GL9WGZHaN2hRAmhJXebv23K2BldoD3m2XYSd66xmHiSCIbYFeOO
HFlaJ90LlsrtasGn9rxMHYylT9uROLxlV0umaClAmo/qdaNpbA5vUH59jUOCKZ1I
ApOzPe1aLXJQUUBqhQO7wRlYfekWh4mJ//ymSuLF3MgFeCYDbJ0Re7DXXGZR8DV/
VCNoZRUEtktY0CfYzb4IOSOfWN/THb+W/5AHLtO64ml69ABK1xIo4gc6DowM+wjz
QMvvH9Z/Atko90HE6FYUeOp2LSCSmAeS0bdpzH+kfwAv/W3OnkfhVMlfaVJGTedh
zZT03pjJ0Jdb995xNX1i2uWq08Q5HkGe+tc1RojHHqHJFXooPCa1oOMLlLquHngA
b2FL0jHOeMZ4mgYWIcjHrSczdHd6xhpBEjubsvikyGtNs46WrBAG57tggkWxCWuD
Te7Ep9UBEDCp9kFoY7bp9Ww2d1THEVlunNGq04WX2Vhp3Fy81Br+x/va7VW22F8f
SkWv1WV1ghW2FAVQIt7G/iPh+CCbD2QMLnEl2+caYW6KXdrxqBtStRKPE9On32si
+c2wxC8CZj4jC19OZxzURyAsAJ1FAB4D2/4hHAdxTZa65gFNNA6BCCN2QCQZ0gCX
8Wim+NWdUiR5iD1pCSJE1vbga+PZ6bLqphu0VY3yTmskMVYAb2xl3oZB1X+KHIFy
ArePjdHKGBs/BBysByHo2ZWqeSysN30hJsD1BuZG/0oCS/fh3QMjhubWluNfmn/K
o1fFuHBYziNdeDexpVWJza/Xp/0e92RESiJ0GmkbkJR3Mzf/tmYXUm/Py6ovrtXW
4MYWRFdC5jMQqUdmJDUhcy0iWI//ueukKcCvqdXUt4UgXJVJK+d1Xfjn7XbvkjsK
Pe0VmuuJAFlByegM0GO5w7wr4X/Lab6SgP1ziSlr/lMWIAQHMm5mR1xVDsKX+CjE
pVPcJ35yuTRuSyk75+qieziFJGoOEn1feIgq98F5zVFiHld4HFLdeyxg/ZLp4qkQ
xNP2L5KJ3gpvGJlJJ88boynIhorCDW0Pk+oRlQvb/r6JR0bhZPYxxAF+YcIyPL1B
TOTojGODvvTKucS5Y+DdyW72cheAyf1OZdqXQ7RqYOemtzDdFhzksMGVWzWOv/Nm
xjTX7SfZOIOpqpg7Q8ZVLwZnheLXLVMZmTY8UJBkRe8mBLdJIshIjBlu0LCQwfyU
T4M8xtXtetdhKW/+QwF9DnTheV6owg4VB+4OdGN4OVB10hC2FTgZtmg6Xbg4Jfbd
T4MR6Z3rZdtoGtnia0YRaLtFX7aMw/FJWCM0A4rhmn/SA9Wn9COPbvBfkQhf/ZwL
mCKZzLoerSRzeMO+Yl1jltW9BjPLZxq7IAWfHGZz7QhVQ2hBs6tA4zV/7b4rrom8
yRNji/oWbhIrZ260uSvEiI8Z5B/G4+l4zMYlubGyMJGoJwnUb3fpNMdwfIgBwBEe
YLDfzb+lzg0Mh2tUEo4+L83EnFrQIV8WNFxLtNEF5GFGM7udaIvnppWmTTWhgxS4
DvtAstOuB3iU4Qt/++Jddp2hZop5TG7yCLClCOw/cIUIl/Z63501Vn6a5g6MseRg
w2oQ36QbymtYwxbhzF/EkuIWnnnzvwbt3DUnUU8JKpUB83pAEsXIXGe7b5HTdutS
hIgrxs4oc4Do3e49nW2Mpd1Dm814DtkFdOGrVBz+Ngxml77cWMzFQTKxLMZJ/GS4
ZxiGUh0z+3dbMmPyVOe02XB28wuCrdCq0ifAr7weYPnXkPmzoC5PowX2bLQeKMKL
k2TFF4BEhs1dRoENdRw1t/ANMU0/5tu+KViVODyZt0cZrfHZsVshpDpz/8E47/eg
epCWp0hrEfoQSH2rpxwwbUkounkb3fPWAT8ciZSMFEoxE0EoUME8b6BEI2U2T20j
ibaCdpkvaCl0LvK/GHi1/wTt87aoUVPpvT+bn1uU53gJemmU9IZ+29CLhgmzclKv
sWdjhjt0GXM5xK1HImsxSb0LLsUZHEX9VqYrOlnV42tS+lOANQ7Uhp6UkpbiEf7L
XLL7EK5Csbq5JoljqGcbDd6Fca4TneCuV46c2hugfCM6ab7YfT5QjK8+GqnBQTdN
SfEzFqoyWftsz8WWCUKc65ir7mZchC3p8wgvIFB/1z1smB34NA5PaQT3nRXkxeZp
p2qRJ/NritP2OsUu6iT5dmQ+6hv/V3zjhNs/5YvFCNLszpo9GH8CqJx0vLAiykWb
fgBNT9bfid3jMTbt079VNS6QvjjhlhopNWAY6B7hS26SOisw75lvKaRdv4k2m7dR
JkBvZX2hN+n1O5PAFTZm/VkHczkakosZsUxmorB9GGGBVfsGll+CRmTU/qCDDSZI
pVg1QRw6ArFmApx1omOV+uS+YKuyz1y7vy2Z0cRnx9UlBxOFkATPXmlKWauX1mLN
XfadMzidx20EK76w0kGkv0vY+i/gr8Xc805roJZCyEwvDriZNH4DijmyJpCRJtoV
mzcgsTfRKmV17o1DyK5z7MhEcudMhYhxqDcdMq3UNNeloXLY/ztJNZQgcX6tPewU
bM6J2kW2CmH0M9YArYgAE3BTYCT/CwSrR3euHr0+BkzxLPtHz1AwZ/TURUv//jhX
hIgkTEhrIYx9zpqAFNGmsRZ2vJZLQG8q04QAAWOrZZxSGdtbT4CEQS3cqbeadTaQ
N//usMfK3euzXMw4TPVusiR6bxK9CFxb1mkWrwx5NaiFISVwC0YFZ31lKdiCs+Zo
c3NyIrOW1CUnqHyTbY81vGUSQTm5Ysk+MIjRAkqcb+79hzATsi1JTCIzU2QvwMy9
HGwJY11ZoBmGG4Q88i9dR6HlCLWTdru/3tV65WeHs78vv6AeBruB2q+6YSdHlPCw
fUIkKtfdPfIc6wJ+N6zkVcDioUcZzryxSN/0QY912C6eYJjGIctfcLVGXLR5q692
kP7CNSIK/FhspHw5v+dZkJ3cu4R6hLbueWSAalpdbiTyFMuKzZueCUCGSnhcfSXs
W+2f7f/48SQoWd7qTUWgT5DevbLPIEHpWBvZUfRqomVTNA5y7akOMSlApXIfu1DF
D5C51qBmiKneO1uMbNBo4CTYGOiSLBMVueZ9vu5Gs+eHDrHssIFQvNJ12WS1lWSy
ohkvLiPqUievzJz09L4UHEtv1KaBpcaVgWJANYfixbi8WI6+PzGVyf6Cz6yGDp7j
zoslRwJG8BdR6EvePwMQvTaw0uyqz9lILpuNdvpy+TBbbQA/PD1DuJOFs9tqpg3v
5omvxkeL8kcr2GXPZlqisw3suDYk7tco26LmrEP7ph3eImuc2bP01HdljbpYWHha
96Hkuau4Xr5jWdcLFKCR/uK1NAF7aZcbPKt+p5seKxa+9zCKY4iNNL9z4I54x4Ax
iAJoMIYlW6+f381YJhzeGWX8DMzv127UxzgVqXXtHvZJkjklSjYgwqGJkSZpELm/
ukYKftd46eftzz0vuCXy3MLspQFsS+4HsJKWQlkvC+yN77SCc1ZYb7tU+NrI/Z6x
RxXGh6/VNgnCHv4ufFJK5A3HdckEW4We6z9nrmC+nanUEBlPtChmYMQcg1WqCxdH
Hgn/gASo18pjqHDW/k0GV1OmeyqEgGpsjkx/lEh9yUPltC6WyH8IGcNt3mCE7uUe
Ps6fizeR2girIZyhFwX8sCmy/WQ8TsZeRjE9N20NaUGXO1IRqO57JNwXB6gar6mV
88Y/H0kss6xsmQQ6BPHqB8uYLtHYxaOFw38PVYx5kDlPZK4Vyz0rCPkvNuzyEXHh
syYMYIef1OZlCxVg958+BDf8ZniXsHRYWvj8aej0aKFtZDxTi8k4AGB3oOqmW4Et
wCUKu2ZnOFOtg1Zp4Fb4Vh513ll1NR4XS0ELcYmPWUd0yMT5zTDP/THyL083dqd1
cDldcwCmjtmVvMMwL08i00ikCfs5fPmPny+Hi5MoezEptnEEgalUZCSwWTu6GRGK
do2lVey+RRA1Ec8vqIo6He3PxUvSzJZD6HwlvaxfDILbDViEzhR4c1CvM4QXv3II
klpjksCP1Idr5KybdVPavm8uPxD4jTM1Tge1uSaJaZfu/LNh2DvZiiDeI8xhFGXv
zdIG3Te6OyMaaZR3KFXgR7pIvKL75BX7IIljiPZMlGkoixKQE8Q+xWOzYhz2tHba
ZaawNprHOQ5wPh7HkQc6irClU2K2AbUfboIu6hOaQmIzhJyzz1dX3VkCeenYKwkm
K1sK/hEcxrCMWf0sOo34BRmd71N10jIUEw7XcJKuAyjGym2T6JnP1pEAp4wYrgOF
V251/E9yTpPahewCtWkVXoTmefn9jNxq0Hjql6VIFZThdv3ugA5y3v6315m5FBs8
+QSNRIrh8Y3PCoBOD+j0E61o8FRftfoZiZ9J+r6I1PUzX1KZLiB3Z8Vnka+ZF8od
N/4EGFgL4UN8Pn42QDTFpsj5LXf21F+u1ACo0EwucXOg20O0ynJ7re2l3Zn83f3x
M3qKjeQ+QVAt8iJ1/I4oUcSIYarj2PmjPIeBBISOcT1cgvkLRDlKF6dSSRt9bKAy
zwEETO76skh0hkdjHL2JhK/e8Ufo3zBB717kC0QQBZfKjnw9q0q074hq2M+Chglz
nGFZjK68AobbmaKTgfJKrP5Y7UHFv6H9b+gEFyvnbYs6zRrzNicg/PhaYIdYwkN2
j96oJ8CEVvEwEH8CNeJTq4WjXjPi+z4D8aYDzJZAPkG4eMkJL7e3yi6GdsdQD3OT
BjI2bzGyifxvn+oe6HnuEurJc2UdYxq+49gempTeABsgm5ZrKs62kWsWLkblvQV5
mdTrV8rSjZZkiaUo/uetmb+MKzYw9ibOKZRRkkcDlpkkt97Jrc1HTOVhgYHyVPcM
hyMLaAzpMeP1yewLDNJZvE2Zr6T7p9Yi/1U7yUeMpDiztGTnKqmAgLwQhfkLdnxo
5QE7FYfKEeQqvVcVCeSmtnEfqF+Z86GkHQEN9OpwyfQYnej9C1PP84wBoaNyCkZB
maf/EFwtQ5kMIqB8boCCMAAHd4XmXUH9ek6IPgk2XbqJ0EZ2YGeOb/MktYCCC1DH
57ZQ9JxyMEJ08MZ9liH1SaAXpNqJ6il2wWCsv96s3c92vz/niRrW4BVZxQORjRgr
ZFn30wKlNtaZfmew94hLggmzkTbB+Kd6u0FumN5VznOBiVlCcHzQci0Hwxun2fup
yPTGPt1afBGEJ00O3lGRGfOMshB0pnjsox9RseLSzh0lBmJzm3f0LPTWqM+kwjbt
Tr7pSmuO/uymV8mRGSAWwHqRfkCO2rA/jhp2xTOk/qomrqpbDFnEnUKppp1JQdLb
SQatYiSG5n2pizMm9ZsbJcsNh91jb4/fcf+cPsq6kD9bEQR/HliJTfRnp5F+JtQ8
2sgTmgK6dP6zfklBD15YLVhpHR0AtC3hz1m0argcyxtzGdBqKZc2RDBhkMSW3v0X
xnuD6ehEqnZTrlJYl+zlivoXkvXFfvVZ5/l3G5iw6WosMgaVPb60jLvQktHELFYw
nFC38BMqWO64tmLef63eSUSTZ2FPo8EA+Y6/AqKzL1vE7gF0e5Lcqch8TpIrwZYx
2wbnmU4g2PG5db+ya9/AMxyeIG3Z/nWp4yYRpuW06YbLemPZS3EGJDVYRl/Tl+z6
lpHPRBOki8bJ6CEf/MOpPRkU6VBMw9gxCNqElfPwp0BFJcN0+/6HRNvBTPJyE9k1
l9SNZA8fEp0tVYJJ244lAbsotfLRSH040ZZmAt8/ry3WfI3mfbdBs9CTEb1cZQlX
4fEnnclwhFgNe2yF1rMd6WyyKfN3AF8rNW1vJRxRVuSNPLcJUA1HLx4J8hWWnF83
Zrpi+2dkRewKS1prTA4GAgB2i1jVeAb15Z8SGgciKeFXrCijzUn14eWDhzAqYBC2
QpFgGkbJucNWAWC3Eg9IXQBXOzCurfIUsI3lnLPnI8hjTjwzuL6ADaE6b0jT27Ei
WAc728TYiRzw3Afs5144pPRxrqF34NkFCygMvQCaCZ45NKUxWWTaO2GuNtIFUaBK
g2/GZLf9WkhqM4ebjQdq/UM3bv57YzH1tKjEAjAe0AHia44vtwl6gIDa98SpIchl
RxOpiB2H8AQGhgltMVdHPYYIAaqKZxphhAzCCXi08zkrkqQ6CZ4ndB+7ymQX38tO
tV36ha8WTdNxADGTk8GcuSS58n7KpZjErMamn/byX+4jx88frTJI++qyEP7iUKIX
v/VV8qFK9mzX1H9QGjI36gqie6z3eTsyFNmhove63EfhDlZtkcR6P1Btsc/BYzPK
qx3whmOlH9rmOllZz9HGVBRjxrAqaLsMmvyeFcdAhsl1r1Zrk2YSzBI1kMfaWuet
gBE1KozKl6lTJZtzP4UtB8uo86O3zyn/vhjCaNZjJ4fjBZIjIzApD5nq+KO0b1gl
8i5dTuSpaHgjixMobfFswEKZi4FbvQrAelkUZ6W/L9gXj0d1CQmfnY5U9mBBQMx5
02QZSbfN+dmivd6P5qXF+BeLc4zhnZaSW6ooQdmJBC5V4LhmpS7+l/iCHlmzmcXq
ipbYYVIXgD3wB2CuiiaS5L1X5Llx+HoU2hVHhJM+lCkWM5Bw1g2YHJmTUGjNIy9J
hL/7Uax+UJLHwEnjmOZbX6osL3V0gE465qUz+o9zomd45fDQLjtX2yokKipS3dUG
ZjpLLsfIbUp0+0hlQ4+KGbTNDccreBYJVgB2yyammhVworcZg+TGbLsNOUsVnCZG
G7HjjMRjX9pzuLvCn5nDWiEPNPcOq4Jsm1iV06OpDbGScQzbIQyiUDyP5WjI+9tm
n8dQaCFnPOOYLM6nhWv/QVIF7O/6tvxbY1XMt6irmuQVuDR7FLWw/NIStb1FYj/v
eCZZ8G9wEwr6TmJ/YLw7RkSK9HpFoZkAT5hM+nCESHqRzi2SQVovWwC/jAPMYBct
qaHAmhkmWlxDEGUWlx1l9Gu4KxxcVBJefvAW2he2onziBIQiZrJhCURQdtKHeC/e
ArUBYkXvwr/3UEHb6Oe3KSzHL6biW6USPAoFWywwNlJV9O8Nz94AxRJnokAQ/aE1
Wu+qSKbYiwlxq2YyYW9F04jRZGp54j98w2Mhyw6wZC9KHUM2BDQ/PQv6M9F0RhPt
SH9oigv4qEHnEVyNr1ammkc5hIswOcDNAZVHZXhJnFc8ukIE67KBxdFZPYEBw+RZ
Fhmxu4GeIIZ69mth3VhsLZEfLGw9+07vSbmlN/vQEnCiE41i43nfEYY9LR4CuaMQ
372bKf5W9qFkVGLvWoVTC8CT7IsnzZ7i75sonCNqZmnCXt5lf5hm/hh8evmNGDu4
1aw6AaDztW+UqQ9nhXqAWK9rBbtuskzRQkDylOJHOhL9Iuy0VNhfBJNhS1OQd/e3
tby8XxdPFI9k2tOEoCJehR+JpXczqHvIBqGntZiKg6pgVIJpZSLFTNQIeDUghDzB
X6rYa4lckpCJsVjeC6GOExtWcz75a/SKT59CgABxrQ0qpm2n/K1/rUcRJOuKOlfr
CHSz3Z6Gf5d7RtKcFvX26FI8rEgvgzpmxQkyWdGfgnlitocrWLgLCeIbVA8K4MCD
H+gFz8sdpJsQ2WDTKnB8MgJnhARkvKpPZmmhOWG9ssoCgNOoJdDWyk5AkOod7nL0
84/lqJ6ky+RSUL5hNi3mC44HcQnsA6kgXeod4iRDbRS7qAYEppWzG9UM19zV+kMm
S+LAhKX8kyNwLQQQFWdBz0fWa19iWOXj2m2Oz5dQFSBpyU/jLMFOeXmmDXzoA/vP
FCplCpkbgXzUc0v0k8DchMyOzWCIs0qxtRFM+Xlzo9ka+1S05mdDOiKdCmWJDjZL
XIOCXNFBqAYig2WXjpEcqpVGBisCdac07M9i9EwLEYaOe72feBAD1QhoBY2hmnvt
EqvAYogr+9mPyYwuKlL1Ur4XBGfJ3HZcm6lS8qohEVwrS0oEfGen8eEZEAJ0FAev
ggbhD6+PrvAOov0PtMvB3xFQGt0fXTPKiqCqHkbsgvB23abi8LI/9oYYrkkU8ZCk
IxTMMllwtUVfWzZICTKmkSMGbUqJUZcnsMz2qHvO5gktQ8/b8qOY/VlX21b+Ry3p
iC5PRkUKqb9XDZ1Mnyu6jb+LI9RPk7F2o1r8FoucO/A6kmIZE/RMjOkhX0KDaUw5
AE5p+5DucPp39W1jhksAx8fS4UzQLxGN+iJFOcFd7wHVzWfmrT2f3FGv7YQfqyk7
9A11mESEXw980TrQ9hYWHSwvW2w7dBhXWkHieF26ix1yGzhWaeixrtMk2hbTUhW+
pFBz76NN2f2hTksu25V7gfdVyBcuFKjIKoq2RgO82cU5ooXuPgR1dRmnQxeomgBR
gHXbTAKMBtS4/2LJZ7960DVWp0XJYD20vdizDPk4VLnXgF56wG0Xi4gmrk357pK8
yfBWEveG9vzg0195Io0QC1RwxOvQu2GjjuAA3XIMdrnrA2ibXjL+5o+JLHCzV/zG
PQW8/O2MoTaotJvfoEeuMY53NYcyJ0y6YSwpNy02XxmMxde/RUn3ByxuwjRO+mfD
54la7afzXhY0Y3Sod/vUQ4+L7+1EscTulMSoNMlDkXp1ApiITApygL2rxqh70avJ
QomlqPT1EvXnezOV0etYgw7eCQk7CMeBMJCZ6GI1C17NAf8Lu6RZEpmi1phPMYun
YNv1AIUN4WRe7QT1am1atAjaVOxjmhoAGvQe6d2x79mGGnPWTLEb6tY5LGzGH2rP
U2Q384ONdk5t1D/fMZ4kzcC3JAT6SUMWVMQq2I70Dmydzd1pswV+jaBkuTf0j33e
N0intvwxNbdW016xgoIHyzO+m+Pe80YXc2SzCy+O+YVZRifNqkocbZb+G1HZvjy7
e7MgW5+zByO1Xps1lOGUHiZU7/xCCh0nsoyf0A9nMHDBEAeJGz9evC3vUAySmkxM
KinJdXnRFfmsneBdctvp5vSrLHLn72C8ZC1qL9AtYDpwOhstKpGwiKVmny/4VsJK
+cJBOWGNA01eaBFrIuLOPVqzRjWB1l9SpeUdWYA6CGFqlBh/yyQpvx4b+jpU1/QJ
Gw4rN/p2NkOQF0xzFH9iW7rv7687UiSOXibyz1Ab4qcIJN6iJrhjZVxIg1eB5lnI
sH9To+kLgDaq2IJO8aSYz19JpuuHc6qPcjycFSdyTp0JXZnBGgiEJMhtgDapD0z5
CajHC5pWw/45xcRYq3FQl/pEnc0SX2UOGX34221td3rVeYvXdcgzs/pXwlRcddrM
XIaPxXrMuwpaPn0IilVIT7zBAKyQYP/hEP/R+5073p62khQrSKm10GS0ggbAhaH2
XFXH9V0s8LKfHSLKI1irhztzXtbO/+Kg+WbBynia0gRCPBdlDpua2YuzGHm/whqH
b3WM7VJttUvmmZNOavFScI0UkHy4DERND0AoxHx+mq6eYyGosr2YPSd3vs9fw2aG
J4bZg1tMJh0VA8kw3hQwqLTYL5MRk3NWS2UzsOzytsqDW8ehC3PoDEWgZ0vWUvVg
z6RRObFIZpyULRQXhug3TUf7PxOFWl8yXCxgzr5tN1MoTPg3tLI4AXdZFxKRLF/8
WU2ATViWRKwhx+Jn5X93Pgp4N2RdV0Fehs3cOVPstkFBpVsePNPI+RanjeSToxCp
1DKO9tUEJw8ZtbhpyGvcUw4DHpB2K5PFVx/DQMCifyifIXzulSlUXPVNbCRjEQ85
lSP7Jylbej87B6HF5Hos6IScNwnkQ/VRiRjyhz4xRBRFqkfDaDBLeCrB6q89fr/Y
REGiNnaGRS5AHEB3E2kFBNFA0hCDP3SZN3+5kQqYA18Q8+Zbadx7B/gYWeJI+G5K
nXYAIkL3mGKthnyDMjPHrEs0imkaSMEvCsaerflKK2W9xYb8gUfYWhd+30eeq5DV
f+tKYx6XVKtCZRphN5LZ/gu2UkU3RipW1NGOkOx7l6GOoNTy2tOYMBqmZu3dfaSb
gTiciJM/hzvZh4TnRbceS7yuh47228Vsl8jrqVUMHWLGXrKCRm9JPplQQx6B7xdD
KAfMPlfIdnUNoZlVSooq7SRBXyEqlLvUhiqVoi7btXJ40DM/TYBpQXx2kjp2frUl
+5RHEk/sYfvBnEBcmDmQDH2d1UBYsCuiQCKnE9/5oRY+BkV36Z3MIZGBA3n+iPgY
0RFFkG5dBaWfYq/oGADg4e5AtPOyGE9QTmsaBF1afzpS5Xnm+iJWT8TfU6R7ALvY
R41+k3YbJkrucCY7aJcT5Orx4WPF8dOA87xdOw4wpoaKTdv+wbYt8Tnx2u9ZulBU
/NsRGfhzCMuNHfJe3ZBWDpx/oIqf1n5Y9kPMzATg/eW7kLLO/GJQlZsJ5WfkhAm2
BNwkUvXy8uv4tElocrgh40HEIiZh/n1WRk7Uamg+5sE52Rjk6N5DW5d6MkfkVNdu
LY/NGvs+p1IzwIrL5fAx4zT5MnpCj9PvVswrHtcD6HR8bpf38yP3i7Y3o07amCZx
udc3d0WG7j7cIznCVdx+0YG73+drIpJpFliHi2Qt4HLaSQbgrM3IwrpDpJEdNFW7
6xqCKtPcADryI60TSOMtPqDSbqMOOhcRdydRghBdUfW6qB6zSr8AR/mSJM5fMlZ7
GreN6Yc3p/hBnJhG7mM99YjafFnyptznhhs2R32iuVenb7+LYbdKv4EzZ/UlO6Lx
xE/nfJSnyT0AegSEPboD6oEyulFAIjFXUkC7e15VT3WzuKJAqRf+JcxPkvbdULir
CSCcAPAQagMtm376ZkoW6PMYaK1JumoRJjAx0/C+ZNJ58xzTKgT2pvDFECAtEMMm
Jb3G3fOHfk/qC9QgWYzUpGUyLY4Y1qMtqbA3GiJCXdwdneFLMtT5XGg56XlGdA+q
PB9b7f/Q2W/aPTToS05XuDYZYzp+UWEEK7kChXWO2bqoLbwgHzmPz1V6p43FVNIv
y6pOe/B3k9QiyendIn9VqBkwUfLuf/YGe3ZYs1g0kP+U1dbDqX18UMRvbRmGaNS9
/lJDJyvkQvwIZHpXVzcmMFMxdY6pEYgRO010BedeKxC2LkhPKCLribMVDQEC3Lfa
B442hnrCXGeEQF4QvRpPcUaR263Jkm//rg+49Rs0knfJsbq87W/aHvxvpmKPP7G2
EZ5AdIcRdqicHkKJWW8wgujkOyhi/4LxkhSbAw4seP25/2xTsdWvHiy1RyVtxyZt
ECz2e8Zy9MkKaao8oRDp/VTQwrhGdSQcoYLENGjJJxGELeESsUmB9XWmeIM6qacf
q3FCKQ8TSVnUsWJ9zBpl7cbx/AyiczwYaQyNoMS69j8fs8cywYLdKgy/EU4avnsS
kshzPVSeHixvuME+wDEcLrEE0P9ulCbJYhxNsFAMmCyQWVyeNsHi9QMWBHihiORD
3SYYYqIUta27q65gi81UR3iU48oV/tNpdR78yoaA/UCeZlXHQV6Sp8MddfCmxpiy
wWLKugQKhKcDlsNUDF65g8dW6jhy1sl0yGYYMcjPDwsNil+MOPlpzEztAwSZxFfA
YMBWd6BHMgkNnSXcptrsqv0HiPfKzHj0stgTFVZ5Nzkh04PXimOSIP/9ZosS09BN
cf5C4euitibED5vcOA7FJWVBuicp+sKZVAOv62xPSQ31zfocqKTac1yDPX5B/Fzl
uS+qsRnAxXJoUOFRY7lVnS76ydTY2FFJ6pkypXMmmXInUODf3kB9MVgz7mrUiqZC
gqNJBlAkXv52ME+n8ddmDNMY1F7JWhxfyohSPrbuFTBXnU8r6B8WtFGun4qlKcry
ke39oBPHkjRi0PKw87eCz6mSCDSkiUQapfnTHtl0Ub/V+onCPh+5qtG/Tv9XDokj
SNcospmyHHq1zlDVYgbSIo4ZKU5YB5mIq3oB+jbpgKz4H9M0yh4JRLshfRMnRQJX
xOahxyFzT9e0G7DKVRJF/wuHSnSSwoEYObE1oKLFMEawOIP6MYn25+TtsWCFTn5g
i6o/UkFNRCdh/zxHxgJ5Lo4tklUX+YC/5Eac8LZZYOa71QQWynGZJzrbqnAr/r/x
XRuNdlXBj9KOuis5qnczD4LVuD6UbNKJiUlhWZtwU87AE36byCdrLrSYiuEAtXH7
Zqnps/h5FAkcgVo7GUqt7XogzH/UMBgHp3RlWTXxd9PXr9LD3f48cDxvFgJBP5EA
KBRLs7snOMtKhOu2TRdL7t54BnftDHMRcqaiUtwSzVlwcM4p+gaFhV4WpH1A7sAK
p8wTN8BIVq+9G2aHT7KGsVruNFNCEkv7atNV6NIltidGX06pzGuGQX3u9ploFgOr
ck7RVrhKbt2QZxd4HaaKi0eMW4kHCZQkh2DaUHZi5/Ns5pvMnVJdOxUkWTAh6+VR
2vlq6NgX8aMpZleWp/Ga2ALeJWxriQiLGEBAOyW0GDanNnqbwB2lAu3TQR9fkrPP
aVCb4tfXQBapyis8neCjvlE2GejVb5xFyQtdX/97IL4aIE2tD1BbjcpZ6G6jjDTu
cZdYLQyOdebzJ4BdtkkjXq9FZCpSor3zMko3OT/U80TyP2UpEErogCzd2qKndEHe
hMQN56WJJ2lnTtTxeXPSjU6l+TVW4534RmxXqEZda+07ZvXM45f0dUhliguYCJlq
NOdYCCj8d4fOwJDyJ9tYWTcZP/fl7AUbuB4U+I6ILORkcx6bH132goyNuP0yRAig
YkeeAutW3AdkeANuXUR+iJsACL4eODkPUk6ukRurKXHYaVkLJixOkonDyvYbej7+
/RH8Owfh4IMQhTIWNm6AMrXBhBSvTp9yk47XBrB5DIRUtD4Wk1qaHAkD40XHJ4ie
kwSswl8aq9z4NICcIg96duD7tSDAwrlCem9en18G8DLQyc+TuLAy6rtO0qnqR5MC
Lq36QZgxFNxe+bMTriu4b/9JtBTPAvajRg/xw15a+Pay2a/Fzq7mMuT9VR5K4Hv/
2kf1/alMR7lVFY6c1FOZJ/qh2gQQY2CjXQznJbG7wmr61+I6wKnlnZ5X2WLVh0wR
PhQsFDVOgZnfJ04KHTk6iGB+EZ0IHBTwsjgkMPIn9MGDsYFfUP97aFyO86ChvqRF
FZcOpHy3fQm4YHjBpaldrIPPAXe4B0ME8EUp3oY00PheuP2ePfZDsS/voYdYJ7Hi
pitkyBvvQTq9ThAmdgdOl9RdW7VRu7zgyg1BAz7+CzDh7iIbJMpGX3c0fjmoST8c
WaOe9JY3IpKLw4Aaw61fMunB7Gi5W0T49e8QXMdJ3xAtB73jkXk1UILtMCvL3MIK
u89wqtvex+0utc0Iu8Vhl2e9cdGe4glYgQOCiTPz3o1KMjz1D8SnuyC3AdqllasA
bgkGa4r7EEESHITqDno/mExvG5AbqFlS/7uJIbdwqQPUloMnAb8NiOpKxc/RV4Dt
RqrVTaqr6cemZPbW0W2E2eOrGYFZt6Q1T3z5Vjt/x82/q6kpGcX+2d2jr87S+JL4
9MWD/uOzh+CtRfPivRo9dNQ1Mii/e9Ul2Td8fPDEz1YhUnC1CVatq41N/QcpJHBM
u+NPEiKvnoGILwlR+w49dkxEC2bEL+6nOPXfZX10pYG/qYgxTNRm4fxuwFx5rKf9
yc6a1ccFcOZR4+4owLwK4IIYneKOSWUwXcqpgFplTepHQkOsb/KHv825qKAd9MiC
LenNPR0l086Kc2ETqnrynYiXFsY+wdqap5d/n7i6s+e0MfBMbrEQUqfWAIXoE6mF
MTLu4vLdNfI0i4lrG0RkjXdR9a7CGftQMVFiQ2kZJGvB0Vr0LxF6LVOsznhX/o/V
BA98zEJKm+KdzMr6D6G/hU1Y5T/93WCHg+N4tne8x/HzlQ0KDHS7AZ33SGQ6lsAm
UXPYUXsz8pa5fzmnBwMDVKB9F7eg36Kw+4H8qz/01/pDuk3OQEAmcREXj3oAmsYT
BQjqfV/Liu6aVW0gzSWf8A9xFQoQEOYVwIQDgdqyL4EBFIAtx5jnH7sxq7R5kKkW
/ryam7/3NKVo3jGVacYIxCdokQ5ahfH9CiVqiMWqhjheBFvXooD6hOsayyJFG19x
ouoZLvXOBewzem9jpipnRcAbfVSdsqc+dyUP1RBkY7H49sv9YrbHdjtRXE31H0gX
AOx3plSqrVE3La3sOBmpoHMSPMNH3Tgudm8FklPtfMhyAVmkV49rsZ1Gonc4PSpB
kSxIOj8jhfIg15CsoecmKhoWs8qux5Y8EzT4TUQfcBrs5nIf6AO2egO1ZYlW/HJ0
4626aGMv7s5Mt8XQ0gSyhmDyObP47/+uE7kbaslI7I+ebWP3x8IIbB+G81nefryj
BKHSsLCt2o399RUqu0puqNoXagWuoLTndwD8eP1IZejCw5YO9rAnHOU2dima0e8R
HJUmz0msn4wKt8r2p8KgLXefkPAb9eLDyFDXE7vmcLYGZqOSpON9OMUBRcn67N5c
zskfnsRbxxzahN8/p7Jv6M3dMja7Jgije9kWO/CQt1uAagQsRwJ73wGfyaKBebUD
ZFkpR4OYG+QcXyQZ5Ctqhzy6fPYUfergUFAYz5CJ9MYBCY05MEV//X+j3woYSA4N
j1okLHtRDRq/G36u08B8Qo8yO9zGdFPrZ06+m+Px3/E9lJrVAW5KCXU8yUMB6hXh
knxWPpIO/mdfO8uu6eU5PBJWtI9/aN3EmdATC7l6sofYgNEbd/yN5QEp9zCwxNXk
erAI30tjA8KmZsMLNjamfuK0e4+DmO7meYL9SdHoPwiB2CFmk5Y9s8L2fZDmuRfj
4bRhrLVMrtG5spo4hm8nXwqTpfUvSUjb2t9d2ajXQF2kKAAcLgF3jY1V9UClDI3A
JWhBFRh86PK95S1PcdxiCx1GNOl8JqWvm7jogK43WIdJjpB7CgVczpcf2UtNCM9E
A4FL1w/9GNsnnEVsKJY+z9sjy+0vg3nQOo/01GomT8YlIkkGYM6GOE9M+Dps15te
eM5TPdU3hAVnIBr1EFJPpWKSd2W3Hjfd5P1Y9pPwE2eTopWbDUaeGfk1Gh274wnE
NxDz8Zx4utbFgIZ8cyKFGQeQufUTq8agmzQmrxvqKtRTrS4NFNiKEWAqC5PjIHNL
rf9DUU+pFWa1nBtA4lmHruwStwu5m4BuvA2SbV5Rq+fVMG4GiyJeq0Pkkvk6e4jo
2r+GskPcuKFf+wXclB1O7oaS2JyQQd+NJR1o/xcv9yj8rVhmSe16rzRlbJhBPkv8
3LQWwwkZJVAdA46nof31muhW+y63ABDukF+1RtG1+pIakug7QFCCtYKIWB6nZxWb
THJ7Fip+9u2Hza1zA+3bYb3fhn6pPk+/t1R0Ix6GBoPPYSXxYuE3r0iQ+7trmng/
X4xyKCMjHh6X0h3Uc4oa69C06RB60HqODgJ84bgFrX1Ski456T95u5HfVZx80cjo
o653SuA2fwIxPFelPMmhmZrv2r/ctMrbbFy8HIFABEK+F7+a2Q8IMBn13wqB7x8C
W5d1LlboUeRu5RswJOawFDi9TkyjcBDdZ7KeeQ1y6obBlftV2mhX32j8fJWSOqf1
UCDxuDts7iAwKb/0LdV53vBqP/2a51z57ZYVudaLvIF4FgLfrXUxhRnbAXLIuJDD
Tx74i/cwZfLjFK35T02k2GDbHxrIS22mi4EoY7U9QC3tdLYCq3ZsSvCQPW0bvBxb
vqpYXE66GHXyGu/46zibF4Xrmgypo/xoK39ZwJCzcZl+bYoUCxeOh6+BTq+8XYRG
NvahQKduO7P0okhQ3MHwfstTxBBeJb8nPlLcD05zf+v7XoTX9HmH1/Nk/2cpExsl
mVtxRR4g/yLmCzuEIFqULJC7+4YU/c35KRMPXl1MdcKRxChGQw4Z3FsSAhXkqRpH
G2sHJ/LqutA4nRUxLyNHzJ9mYSUQz4n0MVDhMPSg/dMBE30bpi9CsR/L3CH8tJpd
n8p47piQJScpUdCMGFD6nj5sTS5mPkTMi3eZh2kU9qCaj3GfO71z/Jhm7szDAQaG
wUQ7Azvz78esj+fUa+d+w9382mbrs1UdFVCLC9PAgOv97kL1AR690yjynTDm0ghU
xheP5Lho6+yY2eXdTGA/sCRARIw3aKBLqtbgrY8yApwBcF7BCNygUeen1n532HDQ
ZM+BUwlhqRWKwtducX8MCh4OVDlQ3xhiBVo3ijKYgwVYLAxMQnFk/seE7+BO8hjM
gqMmJazTc4F5uH6I1b/Hs6HD2CsFRmCU3OYsNTU4qGJuW8wxEtHgqx2ztPsI6aFo
I3uA99OhEUZcDvaEid5l/piuKw53iIdRrzxqIZwpMU4ta4XPfYEc3ohcx3FLGAem
pv8nm5MDwu9TQPrHO3vpORAlVSID2UVQpXX8Bmfe2GRbDohgWR/BLbqcuooRNv8+
0R3rD0SM//TzsDOl46TYaNa7GZ01VzxKyNEroYt1SLgDjrzBNKrLWjveJ95gpUKp
yhR4pe1+VSf39lwDH2jXYEfswEdB0GkfkEvrdoz2HzB15gEM7U9C7B8V7qcuUOaD
hx01/EpV3Hk0Cwg0g9ibIcv4z8+hlGUn8pDAx1ZncaXnVhb4neVd97dxQB909W81
UmyaAmbertMlFD4ww+dXu6S7nGQGhvI6BWzfeXeZKjLHmy+3czu8lIR3Yj47777g
xRQuW6sZXtE9CQN5e2mBubiaVBx7+GTlAbBWUspLI3bGWuM8Y946/bFLNPNdSGOW
wZfBIbtmnMPmxbusiNqa8qHqH6c0HwzG+kHbS2sx1jEPH3TsePs7mFtVbFW8gAzb
ir9KL1nFSTD4u4Y66e+/wpaY1v59IyMgwh0sLuKHJJXQH1V0C0wVXT9DKP+f3LRv
hQDuXpgpW2HBYR1Q1fWxr6yNjnLlfNIvYOpbTqlaYTy0/JRPfcPjt+P8wDJ9AtNk
FCtBXnHu5xTweXMz72b/qbafbS3dytzSCqi9q82a0njVkzd7wMH5Rnb3/f101PpL
LD6iAD1g7drkmGuv54kj/bwAYeyBEh4SmJAvrGQe7lhLcHvOAm6/P+zM8UdKupjx
FnYQo5fcospE4SqdQ2XKMm5eTUUrVgbnjiPBeIIiKv60SJme9ucwfEJ3b/uRCQRV
f5OdiIJhqcbdgCsNEbYR6nq9X5AqXDYF6IiBI3GkonQeF3cx5PRxmK4Np5ls02wN
6ObCI0lRuzXofGChXJTreSJwzEOHpjpGY0HUZsraqv2KZLOsmme6eSgaXL0LC1lS
ZeGctpFzGh+G7NQ1CafBkaQJG3PWLr/ev6nrhaK/i0e4+/T5TbmD5jqwX5/Jmx2S
A/kkSxAXPOvdYE/HqFD0p5w30aHuhIyS1FFIwJD0rJgvd17FvL4rEa9GjGSyVZkE
ZIEutPzAVNUX0iLUy0L0GvCn9RRl3iM9R2E6YFZ/Bm/3x0VuPgOloYhVVg1RXzH3
9qgZwPoygh+/rP5XGCbfTUQKw4TQe5Zux7IT47Zje+oTTZM/to42DlMVnxy55p3Y
ujuAxo+DBTv1KKwDOmCWq8jaSXb1RvtL4ufM/dsny1/MIMxokafR2cgAeqs0LDSp
kgmnR8LQ1IjeLBDV/f6LGX5aKzvpgG73lTq9gfYSTVJlK01RI7zu+LJOhWcXrYAL
M32Oq+r+3mdqrU8q/Uwr6Rs+LjpOX3fvtDX0qeglcSW3GmU0iY2hWXPsBZr6VZEb
oSyTmLiIiN3zILKtlhWVuUv/jlHjmDdVQq0DBpHpqPqOQ7Eiqg3Yd2GPjh6nM3dg
o6oX2O1vDQXZtM8/T5g5MNnufHvRzmLG7ZLuVdCaiGNBdOdlcs0sZpJfyN26++2G
foAlbPxi9Egq38l/kCy8cAJKLQV2wE/maoMLQj3tsNgxGWiaGhv65pGDoJYq+Kgs
5A5bq1dltngg+1FRG5fcOGbTF9ewTL3KlqivIHr0pwS90/pN4S7ziQIo4eNwskib
vjc9j8He0oYOoO3m8s12piH69TGO31h/5x6Kg/PzKySlzJSkYDasBXhDb4OX5jfa
qN3h4X2qP2mApJrMBIjaDIwyjQVSIhN8gG1t9Exo2qhIJmAdwiE5OX9Qg5irWTTg
YBGq/pw92pzsbILarfzJ61P+Xu/x0sVHyTez1SACJ5PSCw2C9QM/pWbI6g8h+vj0
0uBL3NilZp+QRXjLQljdbWMZYcs4NOSkF4fnFU2TWC4CXAL1lcckldLaOW1s6UQ9
oBBWIbW+wtD9X9DdjLtojkV6cqM/BQ/RK7F2rLOyyLUgshK4ZjbypvjScuYj+O2j
wR4fbHEgwb2GA14IKFPr3YX2BwawhrZ7GvUHVJdxD/T8y8hLE+l74HU79Gx+2G8z
IFXnV4pwa2vXnWUsdOgE6QP4Esgep9KsohJucRSwdpeXKmJTH7I5YtPb908SSb9c
qOtNIgzfYCuBLIOfxF8I9CjyIo4T3bZazB/UkyjZpqTLa4D2/Jli80NiJKjVYUL1
KynE3uDRdX6Q9eOwWYIacfs7s1vsQadIIwgV5GaAITP6dYMOfhAglKEZjHxZZuyx
qc0ya8yiOi5E1hZ7kDBLZx1kT5eZUnNmOi36H5eMs4u8U/l2Z9Bon56ygY15CDaN
psDKpekvkCRYI48qfq7cy9FCckzhv1wzhw6cO1+zGBuTVvjH5EqkJRKI1HanhWnw
2AVp914Un3lyMiRACBgaW92If2rMZlKq7lFMgLAfl1cgPkVxYcH+dh7DsSb5zudc
lbjD8+tXeRRcylzOKjP6bknv2zQk8F73whpL2rRIQNYH+lleJsvQL4OJwUI0Twnf
nNMUT+4XlhSXxMrpJ547v7WNP0eWxO1LsCXkVCPjf4GwgYQhhk6GLqXpS7rurOm8
v0NAy4GINpNv+CdXbxmu/vSLXsgYh6L4m8EKZ2NtUJ+a1BwgSL/7IwDdrS54e5fM
4TIKg/WU9f7j7CJssjB326/ueBv5CKT1DSEPkWfG9U2FSflQOiKG+jYXmpqbbMXY
tgNDqLst9wdpw0y2FjcckpO6HuumGkrvp7lVoRrYsMsVsRI1P5Y+EBJFba4e2vVs
duFDwlY+ijJymUNXIR6njpidVHSAO50RUdgtWDJAcTa99wRJ8Su1fA7ufKfUkfA4
Jjrcy3l6ZyzlBHBtu5shonAK6yChhtqacp+rXdrVSgujjvY3rVhy9FEo8MCFHidI
Nb2+0mpfJGbP+IHJmkUILv4YgYTtJp8NDuizgxRRdxGSXEvYm1NJuXQeCcFvlQeR
u857WdaNfRNcU6gzQ+PeQwVTTXB9Og5xfR3xsuZAASma94C91KQdPVPAJdElewpf
TwVrgtahUmLm8i6X1pKpJynW5IjDBrPijCcytZDOmKoCIbu9rbDCEBHsx0D7LLAx
7pXw7ufgs4eCyyXu1MJ8Q7tF21zsPZ6XSV41UU1zq28x6ficmjMDBR7kRBVSoZEc
udxkev7LuGsW56kEbn6fPBDuRozcHbwqpTlpMOB2r1Xo811EDRRuqjm6x5nb1MLf
C7S5E/ppByj5JRGJtzsdox5b7Aaw3tFj92/c5vtevK6w7wYYR25l2CxUh59RGsly
sjfFoRpTJw/FehYEF2OFAdgcLjShOvWGSqbqWAO+mSKWbSugbQTDYgX9uTrTLdS3
f0JhM9EoiODhSQk4AWQh87tOfwM8Vb35vIxZKY+KoiJxcNHCtvm7O9zhfk1fHLM/
CqxEPyT4rADi5jvIZx11T2OO25GTJwmGr5Hat+c9Ssp+hiLnw5bgo0nzHIzHZWuZ
8JKrS6nFRh9qSFlKMK16l1gZvmbroRWbJCxGGqmiib4HR+Mbi26rqIMvL8662/mO
C1OGQ04RZPGuyjX4dOth004Wr3C9mqiFGpKZFgM8E7+gDsdy69DWiT3K+1BV0fp+
83MRZKg6bjBBhXWIRA5+/WqgtKjOsOINR9vA2AsogZEjHcACt9UFdPBUJKMXPkAy
9BQ2JNja2r5SuqOa0aUSt4PB3M1spOYuywBMK+mNeCUQ0LewXxrMWGSHIbxoVyai
l1YUbTn5eyf4mzwucgh1dO2RNPybtFRl+wsfoaQvQM8A9IOJHKQ7xgeE2NpUmcE5
E+TLSZ/7kq0hFFMGK0M8odvZON0i6EwvUS03VWwlUl1V4DUIyjFLDGAZoNaBrtGi
AaalDyEQFmkuD7oUeCPad1GiGPnOEM4NZdm9A9wfUbUF+r937kNcjt8wEMDsVleE
a5fG0Oef9FByUsIBIw2mcTh3uFXBMM1Sx/t2NwtSfQtD954NGOS1bZHEZrQVLZTR
NtSSMSQuwcp5qw9grgyzz+jYzHy0BXuUTVhISp2K/3v2Uz/QLsuFcHqK/GcYN/rF
TAIRZrpqJ1BnPtABfQY7fPuVgOvS0nRi7/+mY9q33wK4MEy+TS3jW53gy0UOySIX
E+aaSitPiW3TkIllQMjq18wbtwydEWg6za4MAqX2prvTtuHDImBkccXKzrZ2qS8O
+aN4y4DDA5eVphYgh98h2vEhMlrqgVUZjegIcwkdD2RXPEhHna9/p0kxgPbSi0bD
aSlq1nxUEIEFIHHpTxG9m2nn0yKdJO+MjAXQi0jEDOAc2Se1aruyHtMEQCzDO5m2
B0QZ2+ZyQKUCdu8MhQ9gPfW6UBLXlq35XkbJPUwiHc1TbiWAlta06+7krbIacxWF
xhmbK2Iup+yQf0QIurPwEOXIoRr7wLsssy73AxjrZTC8FuOsJXvh+N/LtQEPyWLH
8Vs3E2p/gZu0Lul4X6YpwZyZQTtJkpGK1QgmTkcX0ucBU3nkV/IhwIdEQaArctr7
zQE2fIVNwvQuSdPq8Of2Gk9fN62JxQKDQILk4/dw20XaUWgSk4fDNhccfZu5S3Nd
lYSzlEy3p9Z5tNPndQAj+pFBJQK7HDo+Bi9w54UBBmzJnhgvtbA8iUHA0ykaDbif
9G/BNki5ZkYSQ2j1YKUoQLsZJcjgnTJidsET50OodIolh/reaFPlyr6mdBuX+07E
7d2vVransBIyCLfoxMgsOLvnJwvxKXZ70bOaahNi6D0pY2HK4IHoIyHxVyP2FL2R
Yl/AwZpG3Pw3O/XO8wwDwGgJLTL1KbTme2RZP44zQY1zayXHyZ/XS8qep+SMJB+R
8Ofb7+GeYJc6Kf2vmfhu7qVk0RMldBlWseEChwgathK9Tcmqp6BuUWhrZZjVGEfL
BoTBsZWeSv4ubRzLVK3ELQw68+mF31RgqpoakA8RXemmjmTPAPQhjKi2OX7tTB8L
Qy5BvKs4FmimhbGZKX/HuezfwU9ILVLXS9qIp14mWQlVHZa6DCqK3ghDaCMQfjk3
xXtWrDqwm4hfw6qLamAaNEAZcRv8n4flfGDmbP4k4xR+UV6vPqdYwKQPfq+Utxls
oZgsasqOrSd/ZbL81arZcQg4uIaR71mUttG26eW+l8RgR2hdTC3RFcdOzNoapVHu
6Uz6/7c6/EAyJRTMj1/Y4hxPW2cG8Z0eqzP69tJojwFyBVB+Qx2QTgVgsL1viPM1
YeLNFvNW0t39IObr3IiraMnFqMqPJkSXDE3rpuGi3X3dza4OShfSsQyl4eRMVHZB
3lnKaw6R7sbhOzHspb771rihbc+9BV2bg9lyHaonp9NNfSowmUWNMzTu8n41iUzp
2RNWQBb6cxRNrkezGmszgD4Yj2fSMDJeWjz8f1/4Kqnt2WDuakAWWH7hCx4uSen2
3ABkWtdhPBS7gBkn6IBVuFLzmoisY9hFag/lhcP1717yRldZGUXcftKI5d4i0Vci
Ug8VFnm1Jsreq0v/zO+wTAy2CbMkRvGbR4xyr3gNASDm4EIxmpzCRZFcCcdFtDsr
BCiTf27H3mliHb6yeCCzsN1IxgDVsPWuUpD6UZgSi4xYSWxmXieHMjCGaaNkqJlh
/ANzEuzXuUBSIzCh3oWtb4WNFrhaQvl2EJk/fgKX4N2mtguc3iz23jYVlQv6j5Oo
XiJP3UiIkVFynWpCOCUdCfMukHkvg77bpum93xxnHjvU6uUH+knZSrcEwm66n0dN
509m+HbwnV6zz4QCoJeA/pMn2cBOkm5cE+nV6aLAfEc3M3XyeB82z6PqYu3KSLrB
kDDoYvGgNJEmMDFXtYY0UCFvs+LpBbnX3hswKUHjH36Q4vlQOdoxqQvzJWyTefq9
zYwUR7NmGExi1cBTSJPaJqZC72k1GYqU7bpBdH6DzqamCjT0q62oiuOYDtJed/Vv
WBpsQfP8s0bK/C0QE4fHlQwJpz4dJ0bkg5Fwg/UENLeQB9V9W6RdUwoPiV/23ycX
mjClGMvkuPdOFqbeOmctd/GIgt1H8PgXnzY+LqFXo2Iu/hWVFxYo09MtitgKIqot
1pJUolpyCpWpinGXxdc8XjwK0K0MrGVKvVPb12nGsa3niruzpQK+hRA++VMUsxZp
SNK96MBQfd4uCym610IiMIaFNj3yH8bkgwLxMwrD3HRqMso0EpmJKMLcYhDzkn/O
Y3Vh5eSStIy/lguAJ/GNVmzD29UHhqfn3xcHUrc8N5JEsE8pfDDT32ybfl807EnB
pI4AAk5YM/n+xG1eKliso/cBA5uNc57F+twEyxObUBv+nNVeItnAMdkhQHFvh25X
07KhFkx2HlBBgIn8lNIrL6qIu2MHSFMs+LWh0wmzG+hes+l5u4AoprbX/j3sPLSJ
FzzRd1fW7Xr3/x6qkEEBj9RJHilBub8QDxdWiRgcND/Gw5Bd92Nd5wnRyj76YgbF
kmFvAyCwK+V9GCtNPHrjwXQAmP7YWynWHy34D3uVhgtgc8ZQk0+OKjY1GZKgL5Hm
m2NmCFmesTgEV99I2bRhphnZ5WRaXYPLx10SWXjJd5sXSw4AZy5pBZL9MFpSIB8G
t+jQX7nDfFquOv4sUz36gvYswMuLzkFLsONit/u7g4EGmqC73psNAUg/BDYwro9z
rx0p2zmxsPHgHkk5jdEOxAzCaoMUR8HfxNfry67XSYl+kMlgA2MSh6hMGW0bLY70
LH9/lrnCBEuJu1L1KZvoiYDZIGuDE234uxYcVwhLsPQLq6L4bSw+X8jnBqhVQBXx
F59kOZC2ZvfMT8UUeKyBKbO291HINzkNCjxKxtV1qbKJJULt1i2t2Z8fkmUlulii
45T7L3QKKLyAWKWRZiGZ4S4flpkrBbJSnAGOsQi7ykAMxATb1gBmsQ90XDVy0eto
cIgrni4TWHKP0zPFuu7PqZ65LsWuLJdV8RActn6M9wT1qbVV9TepWn6I4snkpZzD
JXgaFMlYn6STWQF5K8p7502xnSNEqsE9sE8apBspad5s7okOwaKX0yHgKoRBUIi8
braw/WqvmpM2TgHfo9TEXw1woirW1dVBvyCdNs4n9xk4gmxZxQiq0ev67iWOgnze
t3ZV3VJ2pSMfK5DupIyj+JxbxQl04wTDLRacYOHB7f13xz2FnsPKe4tlhyZ278Cx
dlZPd7s4JX0lFIxgH8K3KzYPvgCypbyYn4QZisy7df+KHOGW/lIWzT2kF+8yEeO7
n/v17fF19oH9UJwqRlzVaGH235ndc5LS8ArADPxZhy0Jy3DrNeNsOPq62+6cUCw0
4onQrBHk1MwW5eMdRKRhbYHwY3w8VTDlHEaIsj1WZD8qCC/WWHRONqxPqWYn0IBQ
wm/OfxbCcp4spZ8lRA63pXJc+FUYU8wYgfi7fVNPX+eSxH56VNrQwYYq0Y9QjIRA
doWNRHLqrJ6SpK7RsLesom971RIh19XEXrmig7Zae1z9oUQEjkcBSEq1Y8ACGyno
/mIBMCpI2K5+nd38viVJdP5ZMMPjz/FuzsXWbC6/g1/RLDbWDGT58XlHUQfWUa1s
FXEUe4rMyQzDb377IAe68Mm1FihTXx9I68QP+NHQxCrlMybTcj3XJgLLNwe+UYvO
T19s3Sd4R6tlxad1dhuiqfj7UALJ3fHwliS3GN6MgStzhSS9gJtpoWPZie/6SXd4
OnlUibnDkJ+apXG+s70UA/VoqlJeRZyDYQ2wpsfmyUC5ofI12IHsFFoWpSFH8SGi
pgcXQE4aAW4soIl9pXOfYswS1fC2J9vpH19cinZolGIkeKFdurkFlVsN61NY++bm
XyOmxQDUnMu4DL1w5jnooFq149UZ27sSStVxYA6hX33Sb2Rkioetr2UAviSvmxxj
RAzsE+vgKe0KWxCacBHbjjbPYw+rEv9ZZv+2d/60cpBqw8CVCHLCY4ooztLPfbtM
DcH59YcOXh7Vt4n6IgpiyHLGetjBNCIrQethonPER+Ekv3p3ozBHHcqhAnt/IkBz
z18c97ocoMBCkHQ9hp7zE0rAXl+amvtv9cHBNK+b2Xm3zsiJut/nutooE6gvCQXo
+bxinKz7WphggnuB3Hd9UUXmpR8ED3Sklz3GyFJWZp7KdIhuwnNnzDpzsT5tKTNo
T+HsHuFzGaL+P8qh/gieeLvj3EWNvSPaiYrmym6Qr0eYIEBcCJWZJKFJMYvWaPSp
iD4Y+W8LrPz5swXO/DqdR3q56UktT+1TIaFYC/Xmc2BjnlW+FFNAJ9KNZ+b6BasK
N5zQU1nQE6x4e5IsY58VcEZwtIwO8DLBcmsgBagLDmv+7i31zBgWEwE71LOvnNbI
w3ihkELfdM7kjwi3OE978Wf2kXTfxnfyAEgCqMbOCPA+6tzVMsCYaCIyprv1RNz4
+EWf5c6bVGXAuPpzmpCcdD/GrjxnQRNJmdgVNykdN9FfIKzG3qcJ9nPd5V2kHXWv
KVrkVFR936WecnYjZ8WufQFZIBS4A2Zm6INXjonn9MlG9WSLOoeCMMg3OlXv3SCO
1cRAimSh+wPyd6kyhlwnimDWoCYnImrdRbcLpaGIIB67H7/o1FrnPTicoGCxqPjJ
svBhT3e6M+Bov91PeEDt7UPyTZEoTkfTqk34EDqPgJBN877FY51pAZhhC0zBmLLX
xvzNo/uBXrV4+VB69YEHADpWi5WxZ1CrQL2lURiohaQOPiH4cP6tQvn7D03nCR+h
S6y4OJ5lbHaEPaF5lX/CAokml3/xwp9JusmADT1jgqSS3gr6k9dpXdTy1nBYJEE8
EycZSla60nA9l55Iig/ZEVNrj3/oPaJMOkIxl0X7kTO4HWIdN14Nd9ne/bTVT512
jJSawBQqS4/uAgr8Um9x21/S7SKRnPkFSsESdCiAfX/zvvhtoRxsZx5l08yARfNk
6AV7ZRf9XNJK9g9CKmQDIOozVza0cy0QqLWLCn1vhr7jkHavM2OEmQl43LzqxXlH
A+dK46BHHykuxOtBBtQy6p9TFKna8mjfgSVbAFpQJj8xR5WzJPJxU7J556GxE6Jv
jTEmb4q+h0/ys0C8N/rX8P7g4rU2ravM4uABLjY/CacTCoGeBLyx8Fr1d4jzsNOw
ZLpIk6Ia7aDEixnmZI+kXRtV9Nw8bMYtAcxW50Tv8i3UyP311jJJdfSWzAair+Y1
VyKSlvnWr/zsUviX2+n4LrH1WIMt917shogOLGdxFOEdi7CPiXnXnaD1qQGhBe2M
mSxwIka0p3ivTK916ru4SjiPKqUWrsSyfkwBIqmR/m/io0sQ7I3sPh0v1e1v04Go
xzlazH3uKfC/WQmVvTRNzDfmgpSc7wAV5ctn+FESGVQrDm0a17+FI8TCEw7lLAaS
1QQNFcnYiSNaMh/kL6Ku3kucv3rjCvzgGnEEsxSHtgAYbuoiPbodL6UYQAZxf8IN
I/PN3IytpqMWsY8Vj2NJdu+a+2PKccv2g2+LIkprw2rN5/kh+TVLhpCQZa7Ovih6
euZPpIFd/cuShSIks9VXOWUdspxSkQAmL1OKzPvHcS8A84khDgDKH6jkjPS3coWH
5cETvRFEVO9ARy7EQ36uubztexKXWvHU71v3EtP6WH2zaUQydSJkN+AQjidfImno
BlLGeZcJJCJMJOWhEzeaTJz+8vt3J+MlaVRLZLEfOV4bUSTcLOjoWypFR0dy5HMl
ghb7AxxEwjTbZGk9BIARsp4oZ4gsZHXp6aSx8jyMNVZP9RldFOi7yXyjQooSmshw
y1Slfo/PaCt3I6QjGQSe5jlMLCU4UQcZF4wWu5MLhWArbRLF8deZFCmwzqitZID1
lqwYu5ZZpliA6IJ6Qs+rKpA0TGbfjrPuNJtX80HwVJcpuQk/dogncaPyKi9a5Ix1
0wVg78qT7SgQrReMl6jvW90jdJjuMQclQm9XteCQZagxWCkvL4KNZw+nowIN6XG+
Rx6HrKHk21eBqV5+WO4Kcl+IS6Up8pO24Z+Xn7tl4FeIdwcnqJNVy0Js6rSQ4u7x
/B154Xx1Yr/WAGgKEudbUaEA09xaiO9CUCSh8PbIoBUY2vIvqMCNnR73AOndpZDa
fxn8fLVaFAtW9q/AM0pwVodUfSuItbktOEp1DMTm3WWfqPKdq247iRt0DhPVhByk
soCBAVEWmcYjhtghLyfz37WPq0V9Osh1syF2y+I0wpEOYNbbQ8a0YD9gI8Y6UCm+
8F5FLQmzyvL3AyxAXf4tSby3m+XeQMdyxM8cdbOpvd6CzuSgtiz5BZIG8kSxt5PW
vykrY5CbAmb3GdzLXV+smFBGjzAInskucpzOInFzWwpsHOjdrdA4u13wwyIyUHj+
K9mTf7MsdLk5f/+1G+r5i94nr201Jr1/lnSiKXmJ/TE3SXFHjOk2QHSWTC9joyMb
AfVRH1xOgmp25WRsOgrfmos2flcB+r+h0ezf8iw+gPuJoz4KYEEure4+Lne5C6VQ
4G6oeDC696vibDQuhFa6I5mzhyGXLk8TYZhCFk5MYqJIeIiGTuhCy/DspPIV4TZd
aw0GhZChdO5tqsizYGvqGWARwdxwn1++Rd/fqX3hBQVhQnLyM/eAuVrvFlGD1rT9
iF2Aau+qRUUKRN+MGsXOi+ZU1YNkHOl2F/2Y+RpuPJ1C/n4DbDLgF8d5G/GLwRxW
JkN0zc98kmdYfAySyVXghGoHfAeiDMCrq8lHS2ZfQbMJXrUOGA3uPoDJCeMKRHVs
BwvWqMBzXISnWHLLA9iBYkiAzXAxvT23B5bXaaOl5x0R6CGA4Fz2v0Z2SbEHVXix
wHLq9rvpmzAXzC8Ceo5zo/Rk5OBK7EfITDoLrZRI6rJOEUVXvE4h5gXJMO/vCele
NPUz50YxPH5IZAihmLavUbJCgE1pqq9eb/YElPtk5wzPT1dTIeQuudtEdnTLTwB7
ws6M7/758jfnXG2mZ2Atib08L2/14wAR+dxoX7XdghRIuQa68AxqDBo3YnAHzG1H
BuqTx7KqUZCHpbCvziyPdo4xWHglqTyTth6TSeijag70g9RESeHjR9NXjqLDaWpB
z+Cj4gQWVbK5gVZuyf6rvaMzgN9wusaODYtFIJDX7g2OAcfgVkUrTkxt4Pp6LbU7
mA6NRekFdh028D7zE3VpVrzFlFrMQO3c+L8QcD+bSX7XNkTSYy4LYccZp4n7dmla
Y7oR78WxJWAr66I7ZXo4ALy3ruDh8TOPgAayDcGu4cKxiC5sVBKXQjcOqukCvGFN
ObHRUJA4Umh/SibP8dCbxAPfYzzfxS8t+rzknAfJLSJvELgnajtdVPx8UwV/CrqX
wY0Laj8mUYQ3m5ynHesuAodX9/rxSBRc8WZmToKSn8qNd9//GIs3qIJffIrtT5qX
nz6GmXdSlOwpIlGu6FLEcKndYZhI7xmVojsyRO8EGi2apqW96CUtqoKN6ugbIsXD
urxyTJBvzZNAXpPzLnecQ5mUAUaLMxTRsyD2GSj+JpxCRhivk9O7cGEa+R4nV57U
RfuX7kaPwjwCTXwfSDswRP8nKNx6WaAYhhUm/o0epYXWm8QYqusCxKqVEqcxjxcT
QsHVjJd8cz/gv+eyepvYuqL9OqZe9JKSIWpanE4xVpolKSOw2K9xFK26h4G4qmp6
2eA7ghZY1qRKAT5V1RwtL5UPlsRmyIzTTD66Krum54IW4+5TLFmf3+I/qeoeLqgb
/JVIt0tDD2Nm3Ic83o4METM8QFgi0MjQ9fpcXNYmvKikQHrhusIBHuRt85syl6CN
DzT4l1kVNTKbpkF17q9fnmX6IaZyVLMApbeyhw5mQxSGvUKOoKEcTs3BEXWT9gKS
x/y70YS813V+Oi6pe9FvyAEB/aI3pGfTFtJfY9gKd6gWZAfHGPB4pPUQbo7dIXDE
FlT7r7DtXb3IG+ypxDvxmasbM1StcULauLVXo5ePsr7b1DbVk90yv9MQkpcodKGG
c+T6wEcM09VUdnYu3nYNonAuXrv2oW/J5Laz24GtOfea4fqeoUHHTfHsmeo+ig/5
qZYrtNHTd/tUAvbCpf5347uwuALRZAxx1u8IUGXHsVwDsSCHX2LqNNMJKY/4ps2Z
bvnFTHSCmF5kEr8dIs8z4Zhxr2KuJ1xHk/168bq0baNQiTPF8xM4m8bUOWHRU3RV
eZ+L7vFevsa/zI8N8vzLPhraxOpSR8ygcaDwnL+H0ky4qvO42G4Kpom8TEmu8GQH
/ZwcaijsiPg1nxvVaSa6ABoTWWg2PnVM4W+FkUUHlv80pkV9eFqo3lVjz8rWPkC7
xOunSQSp069kxJzw2BFfFxnwoSMABgK13d606cB6ve/DSQj3rXptShrawAz5uH8o
dqpf9QGVSu+C6ks9yhfKiKF63YEmSPQ8/niMB14ok4Cg8HkV4UQOsprLKROXcqes
SaYlGxHXV+0E5wb2FUhymj+h9WQtnQQXHlO9hJ6KyQBHf5IMkzpJwKB2V5gB4E/i
JVnMbBUPdkQVO097K6l8J7Xl6ffkM9tGKQFaurR6n7KGIA/5MU4ibsyd1GSGmEtC
gOXRQvBfU+0iDkJH+zysBcfQ5j4F4ybUIXYOYM1Tt7TGnfabPKfeAi0qw5km9O/T
Ybt7Is6IJSlSiULxY+3MauuLtQKkegDqTIZAsOfPfWr6yzd8sTqfvz8K/Xo9Vge3
m8ZPV4VRjXT6JqZPYG5Cnb+hO7uaDCE6qbaRv2qCE7pAhFlV7wuCxIyMO8oexVfC
FTIGD+iK61phGOOKv/Yt/sIkQQ8Ln2hgSfKaFjLWCx8nJwRbuYDs8SsqdavM1hXa
u+f1ApKHg4Ds4NcC1uKycUNm1VU4M+9W8JhqWclxOWv6V9gYZfmJXf5GdmPbqIB/
d77NemIqjcgLDeFvCE3vfREbaZCWQtboADnmT/7zQdeIFVqwlL+178671tKkAlpM
V7oJhq0++ewNmWFZH4q9ntbSWJMt7jaxLEijIHk5MFiuEYvjeiQEOr4fS8zKQC53
Xn2vmb+MD+KB7KHQCeBROL91J1Z3SjKnnEaj9kZo69lq/BQ4PsZrR0OiPs+B6n5x
r5ikKSb7c9JCld4Mqh22MqKLctupft69j/hXMJqeh47cu/0+F2G9g8NVOQMl+Ftw
iZ4tpzXQ5bw5vIAd5qJwfiBqRnR53VnVukfMVAU7lVRV01efdjC2nv9q/6fcTcb7
eW3nyqHkkXcyGBe69lZ2bzvh2TZLhSzU1N7bTN3jt/bozTjmv86CB0ueutyKKoUN
zaWeu/Y2DzMkap2uGsP8FrtzA9Zv8JvOhVocex3y6bPZ+DMFV+oouaQCLIHPZF9n
f578j6l7eF9oqbK+T1qY5p/KvcxHuFw/apKFGZUPuXy3lmEmfbstlwt1hc69yVMd
SOKFY1KYWJadMqQcGVuPcaWQmk1ZM53qmKcYY1MIp7B0y8Ekwugcrhu56mKBKCPJ
Ruy/oPj1pSQ6eMtHbjsPfijv8PNi78DeNu0QF2+Gf5AoNEw2MkyZNx4xRBv5Vuww
PvSAAtCtp8fGXE78kRT8RSOT23CCUvuI6lVpHe5JxxL11Ka64z5dX7GO2mRmqyBX
oPuM3zQw2Uyi5FYFWCx8MFNRV1Eqazrg1lXXphcAPKUNB0tlXoBv2FxtP7q+jST3
yTlcALLwCNIy299i3AwetitEW8HBWo3BjPL42XqRQBFzPPpHDQ/MSoba7I0BWVXf
qei/A4aFc+JEjV1bJ5N31MWsK6SAundZEG57sxk0YnF1KE8UMX5uZ02M12yDRy48
RGlbyaVkaxbGzsX44qDtZgdrQJRcSW83lr0HUcrjage0VJzCDrLVbK05jjjyatOI
Z2bfFtDSpJp5/T+54+5rFUbMLn940L6e465A5palRfoWoSFO8torxpRKs7XOdFl9
aPjdUIZcFG9PlHzXs9OfRmRA8MQYN6V1WhlzhS4gwLkSJa8rEsbbZJHm5JsGCmPW
TliaMRRgr7QJ7n2Zs8QoSsgw9lj+I/ohriEi28YTQbRDlQ1IWA1n0ATMseMoyQvj
znLQlrLNS14X5Lth2z/braoA/lDzkkBV1ia6WPv+LDjGyWpde332jDMz5IRfTJAC
8Fkb90KeUQmbS+tlk++LFHqgBrBBcnWSImzARpVLzUfK39dF22r4QeXQH0u3KB8Z
L/y261eOnuFRxYRjslGq1BF2vtubK0cVj2tRQquYclgiAJg+fvD8kw7/tDN5TbP9
XVjwJyaJNPMzOiPmbjd0ijS6Q2ccGQNaLHUVTAyqoQYl2z+fvkhEP3tCAlAUMvLB
3XJXzjDy9P8SVkBHvaS4xOCxNNJJXsIKuG5hOnDf14HU9Bs08lRPuZOB4msRRmS+
D48rYOMHAz3dHfPVXNFI+DPJchppJ/RDnNaRIKeJCeqkHeHw/aad5iRZpc63QT/I
sYYJ0R++VOWoSnck1oAwgAQEyGzdBTLq14eQy8+AT31BbFkxux8qlEUcXEyRh23A
JUopVvfdjNyqDiZAYKIyq50lnn6/ee248EkRDAQaWXZg9dTUtZSyBBBO9U9ZPwbP
f4JsW68mSmgYPhfZMV3JMeqow2JYl7dQfSJDw8ubAM5YLJXFM1aIXhNrDJyXlvQn
mH5YgsugMx3ok0sQ26QmKX6eCQM65IeXXx2YPqnPPhzeqL8+upPdCrVKEloKVL+y
Tzi+UMn1rYbT7Jbf3PHxj+LWVkMz3sX0EJxmaVfh8Rfx/C5gLWBuOedjm6XcKYMX
QSpMrKKT5TgVMWNobSXkRbEmq6TmjLSU74qAIaMcsm6VVc5z5mYh4aU0Sinuipg3
eanfMXWYafvaW+L3NoWqupWj4lfKiWyzM2KKjgduH694dRipNOyDpJZMtKcdHSnX
XIni9w52KfjzWDPbhZILo6+e7XiLaVMfeEltuNXkIG6VNWE7lHgQhZeGGxZNha/Z
s4lZk3E1Ypjl3FI0xpdKKIFS3iTmW1s0cDXzsB3aSPyex6CcB67AJPe/eb/VY2/N
51JN1j2/7ojKS2A/JHKaFMrNa/ar5Rx3AkSyyNd4ecmnkddEWvkuauvjTLLUXxk/
mDNygDYFoTgTt+qSLvAOFSd9nW1ka/On0AOu7i4Qeo87yKwPYD1ph4YpEuJoUFoi
dCYONkALHJ50Jiw9HmrUP/DPF06EbfohWdC355neIb0a3OuyXPbMx/+XvUfEdkzg
/9xN/I6EUfgPAZAM4V0KioyKzmrbXPuMkq15ZlSd+g2GgEpWMI5dk/aTKMtI/gx1
lsw4XPjoaANt83ljnpybnbO7KrX/yrzK1kNUhXHzO07S6OGXVgxZPt/Op3E8LDyN
f5MF+nzFxgCRhiU+K/L7xaYhA1emLYYkrJMRSik/aWqR3GOs1lwkP1rIXsHycTKZ
p3yfnXHqix7/D1RpSvOhldUohbikl8Wj2RvmhEZiRJBmbv0V2t9jUtyF2xFlG1hM
D+ad7lZW7a7nLRARow5pzJbkdVNW3bYBhVRwOnSZkkYI7xFxjAm3irb5pdzBYnzR
y//xA8PJGfeaBvuCnoR0KayN7sDjGn1EuKi2gzyYhMD+8t/fBdmQ+r/UdGuvQYDv
DHjXHYoxRuLTbjejnb3LVCmkjfFWovpWLCCB3Z2oJrV5RztDxAIvTyWd2MGx+DNk
MHq/y7nhEgPgzGq8LYTWJkCjKlG09MlsE2QTVoaYzRFGdHrgEHo/ZyYLqlEL22Sx
kP3SWe5r9PU6sZtv8NbRGBgUkbI5BUqj7J5eAbQTNBS93OWvuikSoADmyuap72/M
lTtyD2yf2seIZvAnX2cbtVOU/iF9us5QjgRuys7P8VAFI/MTM7NBRVOMprwlrZIx
cYh431mjtFlOh2ATc7Xo/cpr2vvf6MWMo+LvSkMVZyQprZKcaCHc0apj43cOHjD3
EZhKi+A0mx9wQskUXjoKjlD5VDwTFNunnu9JhzlJ/k6RygBMsbHE771YaUNK9TNn
JO/b29WscGOaFkY15/mnaJezNCEPYdpWftw+PyEZFLDd+bMhXcJ43rTdNU/qCkvI
EULutUTO433X2JFPVUWgl6fxq6UX8IZjQs0RQuvV1LwJ1zTcBdJ74gK42xWwDLeP
9xky+RpCzBchHtw+gIK2v78+kXO8Ik/xoKtI0G+aqVY5uCSxBET51o2gFlyVk89m
muAf7UYJ07LeQvcUEOASR+z+ZVhk5vwMTRXjaV+yhiGglx64FSG8m6RmN0xKMRUP
58hOR2um+NvVgXyn3yP4kPvXQMHrGDlgksgtch5Dk3GEJrwxYC8aRXjnnO7g4ScX
u0oOxRwVzg3aTL6c6OxFtdtp57r307rOR9rbmMzu9CnuUdvlD9df06f3njnlEzk7
hJ679uBmRXhkIobUWD/vtOROL3h52qyX4WBwQhoyngTHVk+cd/gwVZj64GJCfbpe
40OKj4iKEoP1zUitGCIY4wbLDiCe20DnTbBujXLlIOpooah32686dv+lYPsAcSMg
LLRSfRQDmFeGk+oVW1dVRLHb0zgfUKSnFSIHd0FXzA6Ee51Ow6kCHTjNbkv37v0F
Zi7A9Ko581dSTS7DQZ3o0x76TK8t36D+vz86NpLpu5NSdLhmJBo1HnIvVd3zgbFB
Hy7v2m6I3BtcqbUOAu/Pw3tgDwwFBKaguQmGqvllybHYRrMLEx6HlJiWFma/kWse
XOBX3g91029won8fevI56kEN3ScfVykxxAwxfAH0GXYPOse8XHpYZ1eDOhNs28LJ
Iu2vUGdBOOeoByXJ2wc5n5FovsIEPK/XwqSZLFr8BZR0Oqcddw9tCbQBX+jGCW7i
8OTYUegUPSvYOSO4UnziT/c3v4gXhyPc0/94hi7MjhBtVKx4o15rnGIKTN0HIA4+
k8bMkclXqFrg93rDAHmLnjXeCukXRaEVTXgSawPg2oHWiYsiHGziAvyHOxs9jbXo
SgM/Kk+KblDhgSAI7631E00a+SBnAsQdrCP8cPHGEbmGUC/ROFhl9ZmsQjUuJfLJ
Lyszj+0UOhH5jORZv+P7OBZFmR7qtwpvUbaiQd5K3M8JnAqZwViieFkO//1hU98S
EhnI3VI4N8g0lMVllWGIbQFoFRdnnX7pnuawj9nsdgn0PFwtzzs5w0eFNxm8nHlU
6YkH1/usoS2MiyFgK8l00PlDNz3Xd4FxeowavjiJXWXnrfEfi/2EKN03g6ykrbAM
GK+ExrWtA8e9nliEOfITlLKC25zF2wxRCES+3dJ5+8VsbKzWKF+etP/xrV1EXYFm
kHGEA/8cbmipn621yyHSe+Bf3e96Gtd3qJ3QHXvXeMCBHw8GCUyjII6DjfgPSU+Q
cn4Senhz4LkbcnO0JBDTfdIji+HgjbDRv0mNz5EfKJy1qHsqGIkh05fk+TTol5zE
EnYso9tjQg1IhCSdy7Nv7pZMyCUJBV6Jxa1T6Q8olrYoCWPSZQ5tdGaTcsq/9PQS
bvasVDyqV6epNqg8vghsSK3iFbnB16hUiHrqqquIS/8zS4pNHgB/JfttgGRZ1+jr
Wy6PKYZp2A25w3Y4RACBgc7gMX7MYDbokAQvBExT5xa0smBDui6rHKqc/dROaK8V
hs9xoV1jmewX5imXn+YPpdLX+TkNQu6hbCa9DgqlFK+DiTIbHsw4Zys9lLzRLByE
Sv/lGgyF2DJZ+2l/3JAfRYqcoCX8js/L6BOAIwRdmwzlzMJlfJPg2xyQH9Yn7YGz
egK+neFsY1Vek9BlnnnIg6MHH7YbbCd+g9yVA5B2VOwkB7FsIjwMzo3LvKLfosRu
WmHBLc/5e3KLHQjEUJxb9w8k1Awn7g2S66lDL0LuVf+OlQMoV+d8N6fhvLhGKQlN
vqstgPjS1K89Pbkwq0ORo1ZgxRmYHjPPBJj0JDY/6XIkF+INqJ6QFp6FItsdm4k5
GafagtKRCOzASQsS6qb8zVUYDjTzOjrPlyyfxF3WIJzWCtcvq1jeIG7AfPNiq3RT
wnEcTKXzw0WA+2ekzam1GqNU5+YkK7YSMj/PUq1yUv0Xe4o5F0Ak+S0CwxAPOgdr
3E4USryIEdNeC1btlWOTtPweXZGpJMi9kryBPhAab1gBu+Rh/AptnW+DuTynotIX
R4Ygy5o04UD3nKwWlWcKR3VfjYz8GAQ55Tsn4EPM/9PxTKRT40Iy1akeBKmYljiq
Qdr8Bm6S2F7qfw0RMDCP3yvy19vqI+czyrVSpDvZbeNVpVHNF43FP044cxW4QOSY
JEmPSjk3sLYccrRL5AgyXNHFaMLGXpgaBZMakvLnpfpd02xwf/P1WlApSDJMwohE
sKGOshdX2qmcU44XpFQlCE+LT6ZIx7HF0zLER+LU5bMAvr2cHMZHDmYZ6EpVg0WZ
gC0UQrEQCDG/Gif6QQeCY1aUcJVb2e0ugvhEBGxQfC+dla5lYGoyr2tYcobs++z1
kUdu6hbmw2KYOq7NzJsU0k9cpidxk1dfXrfwj8tULAwgYhP/xZqo1hbc2rppj7q+
HyEKata7+huHaRdoGhOZ8YekoQEZjRodpaAJYA+d9SIZMnsyq0XrGCFrLEmqzgDT
1/LYU0z4FtM5n2RKZyN1d/ugNUWjmj6pcqOtVIndGc6BlwhvjChxHPNZtN+iV1hu
KNBviPxd+H53/cOW5aUg2P5I/p0t+quYInmsKIF5TG3h2hQXm0iHDqc8DYk9KBPh
Uff5j+0S+/YlNjsbYE88jeNNsmjmEAAkBxn2Soe/pTaespVhT+vfSGl1olhnclNP
JhdZ5L2zFldt/f5LwdEuyDhwqHQ3zifJbiPKUtK5sUobweRPb1nShdCk9O2+Ob60
JTgYN4+AXZaUNZ6qh9GXNZwroBSOlr0KrGD92nY7x+tXvs0FXnElRUdHrpj1TSn6
rgARBf6dMX+e+hjxXi5rsU74b1n2Jz1KugWcGu5CdSDi6/uZqLHu/MO+jfswWWVa
5fHyYchTFaEUUQb14lfcZm3bv4kngE0W2JN4qIa63RRPPJ3dXdkxbVzCJ2hTCnV+
O8MqROvraLetKlaKgfP9mQ8HDaIxTriKI5Ss4LQkF1dXfUc5vosUuYSZ4wvLoMk9
8EDgUhk8n4FcBRdh45etqeuI3Jabb/yu3Qob4WA2Z17Wz1Y+Y9StJWiC5BBgC/Mn
1ZU0ZxQBtaHq4uytYr6HI4XRUjyX5MeBQUoPRWFmTsD3lF1CVj5S4U+rZ9CADu8f
xU7ul4d7zhyZ9A71e17F4ZXL7lv1SrnaPgqzW4FehbYw6K3A+23svWCsMh1mZUXy
LpLuir8u7RjNbzLQIYmKerJnfztab3uFeuS+/mGrhCdeTLwCnlltq3dwcRFhGqdG
hIYG5BRa5VsUeq/KcAvZSPt8oeVP0CWM0F4IrFrO6vj3Hnol3VbJwxEuVLsOhI4B
dXvfbXN+Tzgf4akCTi/EomN4oZhpPSQvnSrbfQopK7BqB8wc5rzPiu0SQlZeI/Gz
ShAu6pW8bExWCtRw52NAitZBg1w1lid+eWpViziF2wiUpwoR3UiNdyt+JSkmqs/r
LZNEMjy17q70klbE4CAuUJ2OnPnXyT4za/jtn/XdgPjS/et96Vzo6ij42AiKhOdJ
EmAnxBYHjqH6fj7b2elyxoySYUUVPz7mMTz34w028o3mL4bQluj+okna74D4+zR7
lma5mDF2r6th28pyjclKDzDCVbOPXrSM9nOtmsMoyPum9Iqk8l+L/FeI5rtZQLmK
Z4yILkg62vTLfb5UaCEjBuiI46abHdbPPry93YkqJipXEC2/kIGHEMnlGel/nTfh
njtxt9Yau09ttVpziMgV0fs53/G6CIPuROZp2/J9otmTwCRIGh+z+OqfJhjjM2RY
12PeyRrAe/f14O/wctcaQQHNYKmE6dgic2h4tqHocot+orfHQwQv/M/mni6dp2y+
B6n7Zrni06bA+RMnfjXC1We8EH/+73AyqkwhnELzTawKZclYBzvcf5RYlmczXt9Q
Mgv6/0dsZ20uD/Rplr/N4qDLEDlVlElG2j4kgm7NTzriD1Kt65IfDS2H2oekDB3n
MoWVBhMh6eBFaxZsMWIixywmS2n+UvBvLPlr0vd47jPuSkyOImIAT/elQo50keNP
O2FwdY69/93LWjtm29TvWigL9RfJfEkHnEQFT+xj5Ar4bmbKkORMGIF2mA/W4x5w
5Hlp1fRFtFvqTMnLK6Crsb6xPIyWIn70vm9AszAAZnZzJeUGwSFwZ5xo7KQfD3H+
IKMq+DdI3KIPXHcVWB1f/qjV8lwtY8oek50W7L3NKGPloxE/uHo0mIYH9bIfxmF1
zO9U+9moUjaLUeKPUaCQdlZqRnFQCknLjPUGSmlvX6ZnUkH6YJVqIRV8UqhxHM6+
ufLLFJQRT2xY9Mfb5tbqwpfZO6OJlOtqhkwY5veQ9mWYkWwjL10xDQejid/WdgJo
4rFvnc17QTGtDky4dXvUF962FdA5ZFblYj+Hs71EL7M3yoproSzfKYJN4iFGp3bH
oLniFgrhuTvpeswgICthelFo1BTdrSH3ARjs4hOTlHs/S1D+7WtAUAc2zj1vN0ma
xXjK10jMi3OHmV1qtY+reKqKjuV5kvS5Zl0gr/1yGt+tDlR6HwVMCSwj1PXcWvux
P166lhVojwLNWs+8WE/Yk/xDm/t85hHULjTlQYGTT3mB+ImsPgGnTqLBM7ofV7ON
aqtZKz01x7XRg6DTEBY5idI+5GDnnk+5kZrulVKmMCRfysNGCMWhlL0jz8lPKuLT
OW4XcxzRR/5Ug50dJotenj218HDQU0S6mTBBx8yNeeo9jG0yLCckh4mTNA1P6VSU
1QkRLwOqfphAjS3VuXGCevaY5D5TMRKW8x/cm7xhSyZUBBDD5wRueEVqerWoCs1o
n7IiMeiZ17GqeVN3gGm2g86ohiqsc0mRViSyqpIH1RccXjqi4gZ0J1ZKFtG8Lylx
1EN9kuU5H0TOEztNsfAkrKWdV3L98oRsxgZH1s8Amfsu8aHin6qfn2N5RiLkxWW0
bx76DLSyRN4My9+TMz3wkqII6iZrfTXzp47jbZrz3ThGb92rgjNYTCO0+MWhLKEy
7CEEMNNy1QBhgqZoo/gxGw2ywyyclMyKr9PXYcrobiYeym42/RrBwpE1+zyAhpSo
4D4PHB/zri45Fh6IRgxhmjSGdSV1XYy8n+OIGKiyhZH96OflFBuxTTdBIzvIch4e
/rPDXCI/EZ2X6W4N/+5nOySYQfoPM7b2mSxO8/5p6RzbV6BVm+i+o7BqjiB/tzBx
YsEO5oZVogPAix50F6hDLgRUGlD/VWQVPzTBQ98hnhXnveNwcb803L9EPIRS1Qp8
ZKYeghDVJpMKVHjjkw3pj8R8bEWhzpb+3+k0MFyfCtwtPqGpXcxen1ndQjNySfmJ
w12SCEmN1kktdfAYJccTAeSYQQY5BBqZDvfD4sdun0/0io/6njwM/Jc1oecZ+iIW
2LImONzaapDwMEDJ3VsPZpO1arf+R+uTTQ/u/h6vGVXNpCzAIyifZ0qASfhB3+Og
+ARLOp0zJX6Qiev3CjiLjwFfXWlZkJXmVNHAfDmVtyhg8VnzA6yiMBikMkis+J+9
fbdwiI82aONW6KxhYeTvjB8Bhbfg1qx60Zj0xgnulZz02dRVFBJauwLMNrBmTxm2
vtRF07MrJBvTZbunM8EAJgrvnOKYOA0ZHlNCodahBwy/iGgnagmbB52Kx5YQjiI3
V8m5E+N8/z0uQNAUiWzchgmcXjI4WCRpOFa7m0JhnunuyK7DWuSGwXDNzhA2oapo
6lst/vVO5vi2X2TFq6EW/elkRtR2wPfI09S7h0XQA9HdoqsA5i0Odd0dvNDA6Z4U
mBmHaDsOip+/r0Q2nH5U2JOfhP0zar0m89G9aR4sgs4xBFaIT/7vSGoIoJ1h72En
F45MHC7a/Z8RVh+muBlOGQ/1SiQFj/pWjqYpkCr519YsrjOXDa8MFSFbyIBAF8Qz
iyesmG4XXZn4oZzPrY3svSx/+a/ehcko2Wpk/J6HtBv9srYQzagHm/GtMAB5LbGK
OmYiQ6PMkA565LHi0tq8+j8mYKMhimx8zd6+sKZ3oZ1+Z10HCj13Un8R1YkzbeZh
8WY/EXgpE30MMPyxUGTlR6XCasETIWadN8hO89PVoU5XmJKyWhgcICCdmspexxfs
zZKxLXP074pPxdWSAsIFo8LL1R0jqefTQXLIrAgt+9BAcXaHIzAqtlxeAfBwfyne
aAcGkGpnjebDGPUGygvF4y7PP5LxSvWbhntaaupvjLRiCXbNiQlOWvTAMozqC6c4
YqXZj7IB59P47YO+pz1sHhxvbbTjyED1S4Mmu9gIml4SlxkP51BoKA44W+w8bPpq
OT3RQft5sgO9AzkmJhjVL0Wn/ve3UL4UqTaOqCiYE/eTV5IP4dOaFNc7Sfj0o/Gu
A0ndKHAzbjHEtwjK8O1HkIxAe0RGMEifJxulSjII9j1IkecJkCLJmsgZIpBLcaVI
zt1TD12f194U0BJyg4QBDdJaPstF8pNj48Rp9SneaQm4KKdAllISR7UKBRbuM5bG
D/ul6SlWbUhE5uHTiI9PpXTEVHxKYHLU8Y9rC5N1ubwmWteWriBxGlxA8QVTbKwW
icrtYDZkaKa5BjJ+egx3xwv60ezqYvYP9ZIqVeM4yDPdv/N7SOWA/GR3tsYwkLZy
hwNlFyCVrU4VJZvh4dfFEkiQN8IjSBpknpq3dantL/9c/xM3QQg/CQX9FpbOYn+U
rtn12Jez2E62icw0ld5UDbeKgg3eUWkRir5dDyQfqTWF2LTJ6uAyIj7vfmpnwoww
rNGa1XeFpgWS/EFHCuCASgfoX7lvK+akj8uc08vv2LjZPK4qLpu5e2atsy7oEzZ4
Yg4weSOt+NpHAE2zPoUF3gCkaiurAPYQXlW56Met/rwR1IA2W1sOAF6wtoP2wOjH
NJg6eiUxBOYtRqpl4rYeYiR3rOC5J8/EmOKdj+TlUGIzr0d9UTHKXQ0Pkx65+0RI
8wssRIs5D3E3tuq09PLhdGKb9fRWI4c6Kxwfs596xuqrwVcpDfmuRj3xxDDF8XIn
NKuz5a0aSGLFYlOZN9X0h3r91NBr9yRmzHA2a4O/zrs0PfrFp/6vKb1eS8fNsSGL
HLVKmKMqBOYkg9zyfR1rP8SklcFhQUYK2h7ouPs/sTRHStbk5mLrdQRy83s2NGpZ
77qdjRO/uqYyZLGs1O8JNzW9U4mkZ8cPEswDYrGxyMkuimJz2PLjfGwVYnv8GcX+
sFqk3QSFjo1Io3MkXsPovzFT8mTKVkFV1urNY/rTm3RyUnv5Tv6E1HWrfE57Krad
xPXH+d/FWrE/n1OHQv1lE/xQVHxtRLHs6AQlJEp5DLb6/r6c91uu4eCSZ9wmcqub
OkECTUOSmOtHzzFZn7YYSruPZXLUM6Cg6BQNgsxGAWABXIgP7n18/ACrysm0qLKR
vKQgmYGcayceWUOcMZiED8pnzA0xw+s/gLhKRn5D0mscf2gTGU6jQ/B+RIc63/fU
InLv3Re7xGR1Ejlgz3Cme71hqS4ZsSIe8PT0fEMUxyJJl+ZTfSss4EKjLpDtHA8D
XKsZN9HY/rWlFBY5Tg9+UtXJDxlPiUHowdEnkHXOYtkJmDuXVED0/OAWi2SW7e9z
o6k1IsRLc9sPgBoMl8GI2Hwp9w/c+8z37mS8cCY6Bcm4Ks2Eej2f71UF7295D1jf
tZo+y4gIJLB9wAQaxbYw1Z2+FObNsHewgSTwUYjSoHsXfc/dp15TDHaFNmJxpNek
Ve8I9ACA613xGVoZy8stsreQ9Lp2JT0FbL6+8taEdSKTUAE5+h3cUI59SbB3lkBy
H61CRggdwggMmnnwQXYNQWY4VIzXV0G8QR/WU1nlAch6jB8GcgQWzTP6Gbnf96x5
qQxwPCanuVuIx80l186keDHhUhsTcm4X3P/ePAFeti5/rRj6XL7crno08sil3CIz
AxosvEzKymdgoAbhL7hAUhd8uy1K8mfC1E0c7O7TKG0kqkeNrWDERu8bI7cK777U
mLcOvMUgq+aYVOUNixlonRRzOrNmZQcIWPMFi7IwHNagf3iZzybqfTE3aPIQKEW+
UOQUUspcYxHweFW6ddYkvG0vltcyF2aqb6cJjSUvImmLjFwQmv1zDs7uZgY9tXd0
FoiGnCSyjcLHNKrPWdIVJ2i6UGFFo8Nmmll4JpPwfnSYH9gkJhpAcKlZ16o2pCKP
plBV0MoRyknCw1v9TQR3tJ+dofaaWhllPmSkeMJ22y1jvbEns+W+FJXdRMdvcI+X
mNrYKvcwkVzhK76pML6UpBfyQJZxWTHiSbLjVLY5J+KzWRDV6CzeiwLQo2CQqF79
kJ5rW0YxzWQK707BGMiBRYOkfTALOISyj5qoZUXtdZCPnhYPGx2bu24TnnUkUPfI
BQxhzIsAbKqU01eJ7/C0cUZQBR0ROP8AWAepfrGcGS73mrcxsv3lalfFH7wUh+Ko
Z/eX4iYg906I/Rn8ZFKPfGuwgVfuYh8Lq9rfqIT3LWxAy8yGVdtHp9ch+9GXjLUo
l/lihGnyAljQ7Ou9VdZ3hT/Y2vpF00oZC0CP7NncJPqtZ2VMq1v9V/08MgLeZR9P
0DJon8d/o5F5cRujwuoryvGA4Iscd28sd+tyyPX7jItA8cVDF0Wb29ur/JJYJ5ce
cuMz+kiMcT6yYwLmT8MC7fRUP4Ph5Rzx043M1oQDyDT/6pUpY9e9k3rPWXL5+pGG
mUgatFE+D6spZbWz/OReg/9iu2Gmkr+BK716s1Wn0yN4ezPRglvbv79iaTf7uRuj
6RKmB5MPfNgyg4IUn9UAKuhDnPxZyihar0y2+LYUZDx+TLgNy57PA39QNSsZpvCg
QaPo4vuftqFvLgfWQejglBzpRksQN8YJHdSx8c4/O0A+gCjV+wFFQMu8Bh13XOAL
gtAQ/dzNvPwLaILiB4nGZYZczm9rvnUwq0NZbcCUUSd2ecelrmN6IR77l2I6pRr1
1ohItbgSNv3fDl71owvx6hufC5P6lIARG8jfj3zdrsJOMmacU/d9U72i7VXk6WRI
WontZzHTbZP3vZl+2nmrqD1IcYvqBUytgezJrdgQgD01/hO3IwHWDZfJKSa7ZhnK
RGGHzOpYEr+FIfHuygKjNYrx4fGnO90yf/cpvT+bjh/2R8qEMaLaDURVWDNcuWa2
8lQSrKfZdcWJeY1Pz2iIhaZmh8Ziw9NCoX4hK9lfb0+Colrbq7dAzEyAUY5FPYO2
ehzAr287QtrY20znNkcXOIiEzqXoG4WkevKqmEvw5q5Mkgxr00bT0KJa9W2aoftu
YK5hfK594i0v+tUoexuVOHyTo2QkpP9rA+XiP//mdEtrFM1KUTdcaaWc0vO9z8Gl
MUQvNRDRvPp8GWw/JjxVuc6ouWjYUzG3OLfCd7Lka0KDuRve19bqD6Tj2MPeE5JN
i7MMVQ+dbSyJuMUqiXajgN5dzhy/SLs1Z0HNC+LMU+NpgMRaRJnZam4ZYpPqKBnS
3f3bvZogch9G38N/TjVfEKOjLyor8iaE9rHza7QlA5ScrplZoFeCysBYQ3YZ5s1p
rR5/amp3jeCUFi21J3WeCHiJSz6AVaFbT/a9WO5rmDfzHH7hKv+XTXSaCfz1hvc/
Sns4g315730rVEZBIT3YLZ3MQUzKoSeQC3lrjr1zrJplAPHHmNvcXLSsya8YaTsn
N0UTLBRREteIkzhANTM9PvtXddwrwJCsjPO/hENSx4FYVAyl8pNfPHNJ0m4tYgF6
ilfzUAx/wPMX6EpGNTYr6+bj1aW+NMiejlv8tz5qXwxzHtsxbclFTXZtaeGdkkND
7omLjAkE5wQjdrJFElqcnIHwcnOXuIg/CPmzaY8e5KG0N7UyBLieBq//TvzrH8dW
WhpyWmm98oAbEO+eVz4zgxe5vNR0i8JSCMeqvjh74JVVT7CdChAz8CWXKwD7u/sB
bCJzUdaN+gXAVouZBhVjEq856g3nU9BLgM49NNF7aC5FOHQ9GRoRnjPRzDsFqE8B
+VctWNlyuzm6U/SmiSqbYXQFdV209f1GTDoizTM/ZXFSOymBt3T11Ltj9fykzxev
J3sqRWB7z76p/k7nemOtAgMByffpMua4EwxyA8wYqmW9oAddbUcGp6qb8R6WybW2
+sNU/d9uJ22tPJiWTQvxhSwLGnpcXm1yaJQS4e3I1eGgj1qj+U0nWDfWxHImu243
unfVjiz4/6YtLPBxaGkRPGnbLFDTICDVT5WlJ+VPCyPsxs86LVI0EqCYHAsGHG2Q
oWiWrCalWARlX4BHkE34FvGdE2y9IMMCMV+YJf+QY9PI5MvmRc8f32Ag88i1H6l0
PpUIJkYjhhXEfbqcy5pzdHed3ZDkEO72GQugEx3KS8wEcsZXGTD+0FSjxlGn4BA0
j2W1r5EHIzfX0lrLpByeM+/3RQaL45sebTGxKP2kxv7AfYjE/WC64r4mNgGsumnj
QaZ7byNcxMAi56xsanxROwCuNqWJWHbtslwP0G9GRN3Ss+mmA2dmkwZFF0Go2SjY
4AqZPADxqh9gJ9YKmiIHxWbHq5Fk9t5ZeGloMfERq11uxgYJsAGrUZ7+zLArKrcg
HkAgIKuUvWwx083kwfW4zmHvcmItY98OHilB7VuUbR2VdSVMds1H6UGeAF6dn7XI
N1wh6YpvWYmI0klyGKdqBe79bq16HxFBPwvRgVKWkzljQpNOv4CkZcisBuXRzuNC
MhBBQaNHfYwURQp4c8mbtEjk5pm6OdPaeOJNFVZUoqllr44Uypk8KPNs6I7AdV+8
hf7KwjeixCrTh+s2kyfATbIScwSw1vHrwHORtPiHS7MyFzsZkJlxJ+fLnkvIFTG4
l4dc3GV6826DfbxQo0KySn9KLLxtaEpxTQaB4JxtslGluKKJV+K4igplW2/Nt+Yf
nxubFSYHpRn+qovDy4dJY3qwLys59ledpqApv99UMmzbrvndkLgkAdUZZN8xGk3x
AR/a+7dRXqzgIPfLHXh45GmYD/wugJm2ZabNSg/Ouf24XNc1YU8AnV/s0/rkpIJM
Jj3WB3BXMdSHS2GSsBl93k76CioC5UH+keZndpTGC4JVQmHYxAKrwQg1xovn6Cje
F93omrjRJIuNROPYb/tRlnCiAk2mGOdT5y+llub/B4yocc6y0xS/BpJtN9mP49sW
MxGKPcJPiguNqzk/hok8AVUmjgqCVPijZz/JAryuCD+yrow/Pd+wnrLeNL5fCh19
8PMz9AqGJRP0Ox9YqW4SiLIhf0nDIm0/Jw2R4B2IG32U32GQghUfBOIW13GKR4UF
ZdbMNf8emtcsZ+aK0avhkgyAvK1/6/fHO1XCs+qHDn723YZn6PsTZJutLHHykuKx
jIEZem4I9pdPPF10uFDXEDmvi8vM0rWdkAez8VGAiafZzltN2IiruAlaEP1mGbdW
wF7rhUOSaxfc+YMaUEaMMt7RUinrNZyzQdu6TujEqY3fpBbQ7kc83icZyKiK84Ff
i1thzp82Uc3ASuiidciCBImQCO7Dh+qONaxplGL3KPE1JyCVPua3XXn77bmVRcv4
alBB+gwXMNkipCMA4tSeQYC0TJaTnX7PTdUJSpRnONToI9ldW+sTJSKXQZb2g6F/
okWhuALX2z3mRXUxT5UR4zggHgDgdLh0yQKD8j+Q+OuBdka+f7W14WHWsvlbZc79
bTddh1RQAA/Jg3+39R8cwwRLvtno6hvz2y/c2yEejZIMb8rT0D6kT4tOdx91xLwA
YKXeUo8E6agktwFp1PO8qOAdPtxvuW7EtTEH2U6lkly1RWBdiuivFIL6wJAsqOdY
58isONd2Lcs07Nu1WKAdZyu+jeKKeaVvVNtI3ZBp0KUe7E+rL/dTCGuc8jx2FsbI
bxjWawojTlC6O72WlkIay2C8QP/gv5guYnYS2GULUaJ8fMtsz7NhMFcM/zp5RHK2
DZgDU4YK7XaFTxbjsquiWCQrNSQI8CA6RrhVNN4XfDPaJ5uLJXhaTarRM2b47e6f
W+nMEVfZSXtQZF10NuA9EPYIV6JBQCFMZMkT5+0vbxkUw93qw7VEBRci3PmJ+/Gn
4h/Sxxq9Ago2WjlmiGb/Zc0mK4N/0b2LN3tK1Fbm5nqOganb/qtsfr172DLJPoeq
2qlZvJbtQ1cYLGiuTdviKxsDt8kzmn4lTomZ364l7QU8RwryktACBmSFF3d6qWjx
XrMJKZjGtFnGNzNXJp4vq2mGzQqHLV6jEoSk24A9s7drnzBhxL8BYqDWRhLRD16M
bXG6JXb6MwVLenjaLvvB3iu06xmGmJ1VnVQp5OIOgr3EVDr1YRLmDg8+wGKkQp4m
p9zR+xvJyL8ZPYlRquiHrxjmQl3vvCOXF6QYNtXXO8R2Hpplld1/CvWJ/khnxxaG
qHf19YcgGH6XgQFGIZFbmFp3AC+/yTloI5mC1lqPnYQj5yxGnEEmvD/teeDjEnAA
dm8ex+wXQEvIM268ShBWlrb6+x/tM6r21X7om+oC1Qqs4Y9BxVULrjXJN/BcIQmq
/PoFXUYeMn+BJ3oy0BTQ1frEoUg0eFNJ1Di7MT5oJBcYPL6ttlmmFCMJOtyEzU0d
fkVhQ6BRaXu67vfMx+rl3UBzonJNFydbs7iZvQjGnwy8Fs13YokxGQ+fDWi91YLg
WJz+ZM5sxIHHDHPn+XaMmmZMpxgRZNhMRbpf1lSzwPwU2DX3pX/EeN69Qx5QzQAw
hzK/Kyu4kgIlsqMd3Oe0qNm1Z8Cm9HBRqWYUlaKLzCsV7xQiMIot/d8kNh8WJ/GO
CmW7pYCesyJnVsCrrVxavUp0bXblzJv/je1GVk0aYuV02is5YuR4ZN9dxtkUjdXN
myKpEC43+wdy0+7CjUXYtG7rQM9bXiuie9R3Hqp9fRg7hsm79P1JLOOT5s80mNvR
/EeJNIFLKGa29RRwv0eLHKfBJNkx6a3WKtnnlH884grKWN7BCDGEjcMtLkePCebl
tZTHS279uRAoVuUyfeJaiXjRbHkU8DezUKe/0zJjfE6N4N/1NLeNubnN4VgvyjKa
Kz3zrnKqIklXZ7AeMKKO/5Ebdm2nIzk0yRTKIhm5mren0Ork8K9rxvVGxGPcu0+A
NaR4anjBBPoWmYZ9XUcRGgUQQesFzg7IrXUXw/74oZHJEDgIltVyGn9xnJNdxvKR
RiMu85P+tTXgNxZEPrQxyYueAw9kCI8O+0bgQjxGwJCoHVESrFLGGiYv4GivvlwE
2WZfsldMoerqkNfAS4ix89LCn3TRgOd03aZ/EdYfvJM77jj8BnnHGQxF35nDVnOq
RPhceTA92CWpW/sAfsGDcMW3Dp56X5UhzQdDUK9Dpaqq8SWydVG/eBS1P06jfVs+
6LCfMGq7np0XbuNECiffTQiM2eLpiCyxO0fzCmsqodqlHHyvd3Rgd4L0+3qqdQUj
WVodN9FGgnypKbcpKrFNJ6qeRQFujlv0airYT/IbJhzthm1amZH4Drif1SJCSBCE
KXa5bQpBFCjHaEqK6IK3UNLrfQXw6KnrQuRotNmny4f9Xip1IjTpVlDCZ5XetjO5
nydgWILhKIFRfm+f+rD+LFcN0VU6ABdrfAnIxTJmEY0zV5N4jtXdVIS0jQ276dUS
pYYvRIkwB+kPg14hwbSO6wO0iGoGVcaWPWkKHv3E6YmzFBY3arWRFQkHBCpN8LzN
4gHdHgNvN0I6tNgbznGi/FmsZVTvW6JuTudA/rfm+uuZVep3cR+l44+PznVVAZlU
TSQ3eZE80tm3LPR0cwFvWQ7ymzouwVCGpqLzGv/k2/YFwE7/7ZCQ6hhwn/Drlejg
5idokLpWU+EjAOhD1jlMMzHNGZ0vRC/yOwFVqZLABhxfWxU0lC1iQBBpmIN59veO
gZZyREw/tUeJzHU/oaCPNBlrYt8KQ/LfDHNSsz4cQQfbqTxbZnqFXuldOeUu1h2U
WpwzftlTqV9VR+yFrPjw6Q2oXxdBOTgNWNgWbFOOwMV0dYiTKJr8jt0gMDYawhKn
YYz0M+wGD5mi8naebB6RS4igqZlMFLoRdpR6uv34CspOaRQ6GV47Vd22KVqotEeP
JVGXqtZGxBfUI0rRgEUifGtP5FLoBvDGmvXuaSrm1012y9GAc0oSKOgQggiWD782
7UNMxfglZH/10vTT/poxBhv1OcYOoCMABYSqLLkUYnjYzphG9yNwmtgCVu/GmLca
w9ZV+7m/LSF/JUnA1xdc7O+gA31x8HypgPytDCE6XuxV7EpXIgCERMptafEFcpYh
zT9twnsO0QGAGKiqLB1D41kw1oFbLH2p3GlYtQYcvur5e8N0sRuDruX6t+PHV4mz
ZCGW77uhjZFmwsW+f0M9CnJwOPVa2SrgEcs43B2P2dh+0OkoV6YI16gJk6S73eSs
AyZXJ+tuzZNaGXmjdDKEWPkeSyy61SFLAtZcXEpj05iB2iS0+T88cM0uef38Ez+i
wwiBRxsl3p46ODKHTpeyqwnCILmEIzlsvs+pOQH5w79p1Fa8cUBF5sObIrJyQeHS
onOhnE9Ib0gWj36jYb7qcCGt6qTIVy+nOFjRMfPvYYlROXP2chzcNU67eLtf4gte
WEmcpqA1O3SKO+itRT3at2VlMUQjgmvES5a173yg23O83wUAKGT1IzLZ93ulgRN6
5h2RSMahbhJjoetC6/kUdF5CRAwxSE7Z9ZOVuoQ0DGCkz8RkKUcOYyKLt8kH4yUy
rk4b44dkQg9zK5M31tldjeMWwIi5Fs59/ysp6RVZXvCjWtP0ztIV72QNrfffhAUf
NxOZ6ZXOaPKVBCp32L3miYdrx6Go+tx8qCJ451laAdOd1mursU9MVIhzhSxW4S3S
6gz9YsDE3dF2IYVtfszXWLhnfjsMssxXhKPRa3Zm8SK8Jlc0bpKgtykr6PEqswi5
Sm9NHo+c3nCwUWLd6ABhfm/hXSzGxvKrDsn2oFhec8CKwW27UEPgBlFBhgSO6NeK
+EsgA7DM0WCNKtV2e7fKoCR9nRcy3GGvcARDlAJKfv3h/l/yt3zEaYzjDU2E1Oau
TzCEz5fzJ0c4HRRZzMHQ0m30jlAspCizUU6fxbxCWgQycmPksRsOWyNuEk+PlGYC
40iE1/2tjtSqheTb5T2Pr8udd2CrAiCombUgLAvIJNNNjSdwpZBig66VT/DEXiWE
zfNI+X/UM8YwitHpRIl1/0zYs+S/gIuRancfVQqYvTQuSE1IHbLRQ1P/zhXDvhHn
rVOtvOyDWYqXbiZYCRlNl6UAznfiFpdgQwZEbW+MFnBfrskEw3qVKlIUMosUskug
InCqoj57P2yB0WaJFXqLu6gG5HFQgJ7hgRukT4LpE3ph+8ePSy1jaqht+6FpcCsE
Ynw3u3NBRffqRTST4KCSfe1BFkc1iITwX72FZj62sHZP3E0kIek65ya+pNQam4rL
gaxKxyTAUQXUAJIVHQkp0QccY7Cm6UhPs4o1HodK4TNGPXmh9LYmDtBDFxw26xJk
9noQyMP7hzt+Yfy69Rej1R24rm/LbWnRy94t7hq0R2/ZO5H8xkCqHn5+60LCYPE7
NLoGjpxwXYQM6ze/6uB5+wSuS1KSyydw6e3j0owfcKnF7+btJHjsWzkZh1OSoSBW
is0Jk0US4jU84/fHKupWIa7F5/Od09o1BXpCJ0JUDdzbAW/zRhn2e94cvQnNzQ1N
KApK4QaSHDDpKWjH+fxUxkfVtRnOMfqQYX5JVdfCbQDmOv3QXP/RfN4+u56JXYBB
STFVLi3KiSxrhQalg0p/bcUTy/914QatMTTh7wwz89TO5tz+hkGXhvQVEv6SpZ+f
Z8T8eendpNNwjBTCTslp0rHE/Z11ThE0ogE61AoGODtFSa9Bw2Px2MOtSoeApPFN
rhPn+55N4HA2Ndlk5okNLo+Hv7N/R38TFouY/IycnTM=
`pragma protect end_protected
