// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 14:01:36 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
M6ScEWdDc5ZVqrV9l5xKt6sxln1PnznSsGlPRICppwlOuH//xp2BCeltA9bSYRZQ
huRUg9RnOI8mjPxLdJGbu+QSOe+WLRmsde0spcZctjqDSoB+8f2N/x5gYN61b6WQ
2fqX0DLze8F+YYgjzd0Wo30jhXiHhnyJOYbhANZURmM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5600)
02YTj71yJUrJYkzg00VsnG7CNk1Bz1T5VhovwP6t9RiztpLKnWJPWEmF2M9D8Rya
XeHSWgVI9CPftXS/LcKWDSGM9SqfhfDl6jAWNJgY9bFoUDKf8kzkKnQszzQL/7lZ
voBDOuaP06ZqhnGj5vebNrl2ujo8GzucNnwEwrtmhTaSJ8kaFIrO7DTXmBcIDQji
cjVUJ5hQut8X2NOI/NTaPFbfmc4pKvMquBLrwUNgUjb6jK8MaPpwKMN9jF9KddWs
yUreJZU8Q8pU3NJh+7phnnusEBd98YuGkVicn7PgKvcR99WY1k0SMiZJvYtVJF8L
L3SWTA8JgeB/NgyJgLl23f9054YgmqSQoJR0dniZw1PPD91om24aJQPAyNEqOtJE
u1xo1xUJus4l4aiJpkhh2hNfPqJcRFr5JNy3fEBhuUPunhsqBL4v0VcUUivw070T
tsa8OxcasORWrShWBssTGR5yVqGu8r//30YSjG80vo9nZOY0xpzRjAshhyeo3ATs
5rc7CjI26XQY8eHHvv3Yy0Sy2JqAqNs13XRZxyt45hWuU924xFV9gSNUE5v+Cmix
ArPhm40VAJrXyXLYDb8FBDozsVzn3HruOiu73okfb62fWruAYptE4XqsmRJ6pV11
krULYUcyMM/H6qZel1wdyt3CH0MbgHJ0AtrMGDu6of55KPJ1aIIBNcai7H1dsmcx
C7qU7R3wkiGLn0eFQgrotvCCPnWakbdaPDOMDnPJNan6CfwWHQkckbD/8/K1eJyM
CMTHiGGfxhYiSj7VgqdC4LYmKl5e1JUvdmHPdCuO3/rB2q44I929AHdWv727ur+0
eVCLYiCWZsaTs6bwkAdb6thdUYlx8lD+/gaob0qQ/2rZThfa1323Mdn/m7vI9F8j
swhWXl4qNCmd5uOG6UDpo/HoTx3kKdYP3PqG3/sa6WltPQkmDPAR6CxWLLNk2TNF
w1ASmgU8r0/dWmhZZHAGhdRieR/xWeOlhA3Enj/ynkxSO8bH9dbcYVIFduCKEOPC
9Cj1ccd4Wjicata9V+p+Lytc343rv1LmUAuZJgl1PsqLqBYP14wB9dpAslUJ8dA2
TuSfvR2SuLsR1WzR0eV0Go4qdxQ+JBQAuIRz6zItLC8ZZVq+wbXW3ApamDnj1ITO
v8atLXkxPn/8cZqSx+F9zuyxAYInrWqC7YimyDPheHVaVxwbxb4D2xQAELKsY+ZG
jJUwWTxM7pUkxM09ec8rIEq85UJNNw6y0kCOncUxtchXqgO8WALxt5CQtM/PrawG
AODg8KxxlGJJEyFrgSyI0sG6uib5datwpJ423DCR97S3gqbC/XO0WTbsInXNld7r
4h1LVwAlM8ifQiDucgihsbC6SMLmjYUI7tmIIERllzuJPfnGJnv5YfC88KxRLEPc
jqBqPVC+3gMd8htCHJh3ICwqcPA+8n084oNRLLjRD1cy2A4Kd1Fyq4VwfUYo2cd1
c/e+ydgv8h8wy/J3ESw7opelZuMOSZpWTSnZt3sFA6B4yLZ4gM/GplnpZhGfWggG
UajyUyoXgkNAGnl+dq6RlcURdSk+Si01+wui3/xgk5g8IzWKvXTrUqQ0xRPu+O55
+rXMfKMNaMyK+KnHN0fC4q1+hn6XtTqkGAPc1+WJIpgG3OMUIopnG+oBiQZxqXW0
BKoCdpRyzOHY+E7AHwfIe0kMoB4G95YbmJcLxwdE1V64nKTOKvQeSpw5/jr/XKPY
/CTlg5RE9W3O4gJD2RLADQ4vaUO+gbQTyprzIn8aiLQlsdGqrLeyiKDYmd0R2FXu
cyf0ZUohW4P0Xu+Fx5oPYmwx5inkX8GmnGgVmwDT5sDzAw2A0ZbZZ02OjH93WAN2
Ww11+pPIMb157sG02Lh3YxX3WXNToob0VG8VzDXDwQyIaDRqOc3O0dPuLuJZoSTl
nEvR6QhjNvPVx2+WOBFI+FDh00YGU3rW0hKi3XpelJaW2PlY24sQp3Wx3yF9fbtN
xGOC0C4PTs1D4L+vdKhXfPgwIKD9TT8Ztr9pVzERW34FCDKrMvDiISkUnDZafKsV
VzZ5xafsYqm6Su9dvzTOhGNan1RyghnM87E3M5tHCRrBo2m8Htak4WgINbEpnHf+
617VcwuSQDs6x4csgEzgr7JRudVxCy9nlbIL07YDkhjE0rROURtizdttVrK/wfkQ
ph8gXFOZmraA+GwUepASaimsqOauQeZ3CWmj/iQ/MgTiToJutNgFI6d3VDy3Mky7
aSqiH4b4gr6TOIBOf3tFkKUI5uLRyS7r37zhq+KC6rhYeAneoDRTqhUjHrjAuCeh
uT8XxPyJ58PPTMPQLGF5Fj6fRQ6d6tuhK4SZNx9njqbRu93p0WLlXNgEabsyAH8c
961yYE1mh27gjyjtvN1Zv1pBxeQVreyNUEbUp6BpekCzZDPsjQj9/s7lMUzDjiKj
vCxgOd2eTsjjJRzZ00wQAFIrN2Y1q+84RypkqcDjtRlaXvGcJf6ThbbvJdfoD2Vy
ynl9G7COoucGVc0cbJRkJMSv/tk/Wszs60kKmsTvVTDw8whMOWIcl28bt8UntcyR
wARpf/qla5ybJIfoHfZR9sDrjwqfoNLUOtUCBxKHTojAFcIPxNQR/9ttjcmax3W3
bqsFcTpgShi4VRsFhXnjshkirAJNAKsSEI2wTfICqfnVHjnA+q8WF/VKb2xPfnlP
rSP084lnln7H9dWcShPOlQERFsKG1biOA6DWNKr/UZF9wiH0M8w6TI0xjdIrSbDh
LeznjXuqmaMCI9oIyxkFBX47eAC7z9yTCtl1e5j8J+AIWihDZ93qBIFi+gfjIssp
H78LBk0H2RO5KKPKWABj8oOelXZzOJYFcXyhHWw83yIQjZi6/fwkOAsBo0OQPJdf
btYaMq6XeoY7CRqv2rndzrCIrfxkQZT5pmpDeYGpToVbfkYcYCJ6bnK9T6JlYqFU
oDU7UTrRHb0OQCCejJBIpuc2mFN/A//BNrv5Jbbk5B8T48MxALDc/XB+PKJfM2Td
cGqkdU9K0RJgra/hzPHnb4WDY9VE80c6jIRZnvBUvrfa0Z9F58zTQayV1AIxc82l
soeKd3bErPDNunpgxPGc5yRUIDWgE0yctXZU/zmYV4MbBM7ub5Qw2cteXflQDNpJ
w9R2TxXjGHQN6y2i7nYY1IFPGh9xCj3g51kXHdlYqCSK/r+O3gjMTy7eiptqlboc
b6ZHZNstjZX/wus9t+NKRGZSJswgZrXw+aivPBaXYF4W/ET00N+Mnn8tRoiReFDd
i1QDUynOOIIkABoMdx/7Dq+npdTis6Iy51bD6K8apUq034VuYuQhwzbfIghlJm7l
zhwt15tFJRHwjbnNMHiUYAmxgKpTk0JB1pyn1XG/4lyRj+f/N7ViQXJ7FbGvv7qi
ZvOVMgm0L/MAS3Pj2PWqhy1U81TmQFDZUq+RYCnsDRrkak/g3oD2suQ5teJZ/QuX
vJGe2tV/atsDFh6oSw2uY4FBxOoTsCu47RSRr0IXzob2idJ0aOdwMd6/cb2vH8jD
WNwRPUs1lUHMHZ37LLcS4PVYVjr1TEvHVZv3NeKfEb75VGu/HUjsTdsYw6poHMxP
gi4xy1+qB17kINngE5BNbiJ0fdjh0KlfbpE1rm+jUlmjg9LZ2B+6JfWKAffoJQmy
+akonWp8O2Cma+KqFv1aL5ZA/iocLOyxqJTmAMKi64AijR7c9Mg2medP4OYFxMsS
iP0Cb3AlpZA7sDQ0vGlyOWZ/j/hlXee97+mKAK0jdiT5WUoU0n8VKI9dsjxID+3m
eGu/3EyzYCwS4wvIE7SYLNScYLDNr38kXOvG0J+c+vjcdNQhiTtKUJUnhyht+xb0
kpfhMcfsCFoCxgBQqZMzFREdz93H5RCB8ZMWN4TxnHgmJPFQbMFm81ZKHANXW0GT
tz/mlX6blOrcqoA9q3PjJp7eWdellpuRWu3j/qnYC/Q8BiFiIBlPgU8sRVMMgnRF
3gMYPq58vJJ7bK4zWBOPVG2daxmYzFR4fVywkquPPOUhsNJIWNTwDpGbknIMTdhj
Nc5ANN5h8+x7vZHzuDnLGX+p9uonlINMDphak0RJNp2yYCZdWMdWiKTYgaM3DO6M
fKU4uiiFaNVhmidZeHkPTV7b4VrjZ0ViAn4pXczxyB4GvtTQkFQESgHhPRElTWhn
8MMVbJlCTtej45wUkcFYv+9IICk9INd+8viaoN7GpWTG2s1I3Zv2GME9oi0/lDmC
hLn8dppQfA9wfYfo7/lVNDmNryRSY4iq69wbCCBte0TFKCIzpwNCkc38miSkAfeZ
z3FGVH83B44CKMqUXeLl1iULv3EJ1ylK41tiVC806dmmgRuMHD4JQxbuFncoJCt/
wLJgewQ4lfuyq5F7AQZa4nevBVlrVyJgFr0KgmfSWLJKPwVKd/BVV1xkvCJY9Nlm
WVLZGWXTcDQFpO5sTXRuwqHdJcBEkrvAS1kzErBf5txawKBolvttSS0ZExCxipYM
lirZVT+x4wVlwZdjvmc+edG63Jt+r0NjTTx2x9tBmTVPkrmBoQm5ancs+qMhcOlg
XDwIx6IQh87uPrYrSncYsGZ/iAdGKp7S4QOmTPvwVv+Xy8io0TBRXvfFqRn0+pC5
QoNB7H5uECfu9yU1m9hYda6y0V3lqgkF7QTHV5mgbbXHCHa4mB5D4pf3uYap2oEg
4GZl7r9pBKfc7N2XKJHXR0QQCXn6yIKKfbnsL27hKZNw7aDK53inDO/F3HRkrpYY
fGbqQ+Bi/kXTl+jVE8JXgu5BiZbIo1syfnloq76ehk5m3fNpDUu6yAo4mm+/U/ot
NwOJQV3CMe+hPjr7oi7XioDzpQq7W2psCml8o12GFRKCT/1VGawW+bUV0qcp39zz
26MmzBeaTAk4DSlUwDW4AgRVGOvGMr0diPdXrXl7Ws4QawOGLs8q7L99vu+qnQZH
ajizq901B99jO4e0ycuxK5P1VhHn0Etu+fl44EFtfk0sBPGsSXGQHgKYHINdRISF
iiUF6d1WI97fTNosRW3KAwhlYlQWH5KJ5Ejr2itp1Ze6f5msttbUl0GdSW9R+vZE
unGP1+i667f7epHNZt1cr9pHDsRo9FWC7tELtGBY1lYmQrJvNM1ZMEgFu3nukcXe
QzTK0YrariarcY2j0KoLiO2NlF8mJkrJZCuZfwxg5bH4+28pkIkFv/usTJbjgMzK
HL2wfjFRs/uzt4+YkVxtyJXNWs7pPF2zH+PjnXkUXeTG/i1WEFf5Aj5XdGPLqK+F
ikc7eW3c15gfFNyU19/9C8uIzs2aboT71HU6dK7n4QhN5E9FycjwP92RGElAjrCX
KDiYxdJABTeZvStMTbjCWplVkf2iQo3Tkvy4ykz/jjQO/YxKcj7IqDnLtwEoJbUf
RXsyyF+BF/zR3Xsi2zAgGh/CAFDBdSSI7GxYNgQY+SlqQ72c05PuyQ/vexvVtcOV
tfLsPUTLVwtbN6OygYr1bhot5FcGgP6tukSCYVyjwF5+eVJ2GypXvuMsgZlsrIbv
rBOMi3LllzIl/dycJlNkg8mh1yGs+KV7e4Epdydkp1HckgAWvi3edeOJo0aC+XND
PtU1KvDsZb0YSofMTIZbSP+8vGyxtcvkNsW68mNA5DaSiCWogVk2iv8Eq/BHFnyp
LlNceGAz5QqCz1DgvUK9JVZEQNd9ynuQCO9SLzuGwdlp+Q1i/reCpo93lSi5QNt5
Q3s3UMQqd29f+rjgGeZ93XZYB4IZnWHYfo5LfEOXxlgcAddDjwDyB+rvSQ8lFCXx
M1DqYycIa6be8st0hM0GqADl3m8O0Ldr4/jcAumCLccyng1U4N+ugJEKcv2t53ek
Qq4hoB31KRpH82nUlEp3QSmdh2jz3gx9aNU/qD3vhotNZJyg+4hQgnOH3MtZRX5K
lXDr24ZMWEW4l3xbAQ+LYFJMX8mhvOnO6nracjFsmzNJLbGiBa3k3nRm3jOhwsIx
r39QSGL7K6iLN5BE+HHC1PWTKXg8bImcfivX3MlYqI/myNesCAkya6tMExs9ZPQO
bph5Yao9MQe+2ABB6lKWVC9E0asou1cWVwOg26wtxha5No2zvaxmu1OoCKk8sdWp
YTL+sT4KrvQDHUtidZ7uIpKbXJdDKEhWQQvw0y20RStiLWI0tM7Twems5dE+Z0gf
fV2gEk65/mqmjIjqVdr+X/ERk1VqsAX1f6g3ZDp22cTfSFd+n+/t80QckoJmpIeO
c2I13xOrB86b9UbKbs4C8k/WfvMAWCP6bCqsKmfcyvOj1V3Xg+7KmuzmHXsjqdgU
44dsnOeJnvBE9ofZa1EUEQX87Mtm78z+TFABfB+OUl5/FW2UW78ngeEJByZqiKcb
8T9godJuup+qHFEt5upnlzte0H1XEdsN34Vtv/0Ir8N4eVJXaJKWf6uyAx+Mhx+Z
iQ6qZAM5vj+KrokIgdkm1B9XJ5Orue/vSNkxlazOkM7UMjbtVKMvfGkFgJgbTWmW
Pt57EhbemrB+f8WbD3cMx8KOYYfnT+TmXsQ1z3g9w+jhYqbJ98S4Dpj+TLYTaqhF
8J1dNBDuAFi+XNyrgDNbyU+PePta0Bkk2QITGWQx1Q+cQXp5q4zENieNSh4Pw1GT
DtZyDx8Rs7bzSpmDB1oQ0dr7/zlc6l36gexomMiKOvBOICTVNwjn2JcDbiRA1cOR
J1B47qu1Np193tJ//MV+DZwLzjfMDv0+o69sb9eW99R1mLu/dODEcdef0avJXxK8
jcp6yFbA7SK223DRojxy4ooXdzaur3QGZpO0aEAXs+hwRI9LxtJkHPx3uFVlOXiJ
UGWdfB6vaA+3h/pFGfntPLN998tiR7OWTMIT6T4baFhXc4f0yt/zHYw0h7bL6c7v
gvC9f2HxcZsyJzv8jnqjxJ4Qy4clKyfUm3NSexoLvc4HGRaqZOojOsITUJZTS2C5
A4trxMv4/9nY/ISwEBkwwIUMC2i5lQoWXZwwnr0RnwkiSQuVJUIUEN3815AE1Df/
VqUxxcTkenapgG664fGQUOcF6a6xT66JQrzud0DK4TxlXM4dFYmZreYLuj9ceEA8
5KZZj81MGMjC3VGbeld0qNXw+TCe25RFayHEKH8QTB7QHZpflRvz5LvVeH7OhmHH
EcFsAHRAsjs6mcVgNhw3pn4Iqd/jpiR4frDayNPcIEMgc40LO0BHIrZkXoFNQrE1
6wOu2G6+dLlKVfaxYDm0BzMD8eBPBhcegKxwLW+kZQWfCLnt9BgTOiK6nql3U+Eu
VoHXnTMKiDMI8d4cpziTciiqCxK7sGtXcsGk2Zy0QjFYNm6gDC6n83gidB2kFCNP
5E3mpp9zm7lXAaV0qNo9d+HyfejoBsMnVd3N9Bm7sm70UhrH7p/Oox5+vlBiMe0/
RQnSA8cfK6Meuxn+JlQqn81ctDSQ8zUTGftm2Y7uEr88rkvA92HrWQ7WekX/A3Xt
rz+6t1j+QSeG6XA08yBTdGPpM+VR9CYaMSquwwxNyFQ=
`pragma protect end_protected
