// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:05:40 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
azQusnIBs8Kl4Iq8JxY1QqQ1rEHgYwCA5HJcTkW2QWqz3669RAmsUu2jHZr9KoQj
IhWNfYqKebqMGeMBHZq6SvxLjiMvUGMngRPsjMvIrW+chrLirC43ykgeKewGkQLv
1nmeLzEJ+xuJglMeK1y+LHLQTsigVkke1L+t3X7e1dU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7072)
LdnTqO2HltHAdH3mYZSQQoz+fT5bVO8qpeII1j6Aq8Z44Nh6vk0SdpBKsKZKxclr
sRi/9a9NSGF+TCuptdb+nZtjyzfbbty+SAL9/bNWGm00aveuAd+FBDqR/sAritlF
bB86AEAUGKkMkR2G49QXogevV7lSJCvh3wM1Ciwaylo1mEV8AROcHIrnmoc/Y+3l
AVv8iGyZIc41KLgB5GAzIzkRVizWJD88J4B2Ilx49I9HvLFfRaqJLWOM2vbnwAfY
8e8M2CJSvGgYxapzMUBr+QagQWOulGK54GM6w6rgi6LaJjK1OV4gT5i0EGJRV1bF
VCKaljZE7n9i+UpIYQnRV5XJLQB6tFYy5DWaM+W3pfKBUOzyE2LLdoCzbdSbc7pd
TzEpKfuKDjB5TephX6ZqPL4OatRjJwJxES42bbs87MtvgCp8DO3uKfmDQ6FB1//Z
/LCfgh/KJJJAHJw3QzXNe2izAMsEnuEFdq4mrnHJuamzQ/QU2q/H85q1Tns1Gd/Y
PtnPDJU8iXDE8CxRJob5QGkm32wOzmOM7wQXbl4EDhukcRpDyRgwj7iJRVYYTVc0
ojxz56t4X1su9zCWLpFQDeIid0o02qH1E/Jef3RjtJ22VB/6zQ+HI/ss7btuHoXs
HaEz9QdjCg7WAEgI1wA+X6n4w5tENryrgKaa/Y6HHiHEazW+aT7XTWEQpq+G4D0r
xBgYXP7icEUE4zFUiOW8ix3zP0pzUtGSDkj6DEbOhrloo0LevMCi4/2VsLy26yIX
sSmBTWsDZB7EqSaldwvGHXFkchuxLvrccR3yydh74Gv4VM1s8KLTLuPr0VkpNxp/
4h2wbPAOXYR8npsVFQ7JjaGZTgAfGHLA8/AC+Az/3t0So2SgA7oxKMvkaLyy+UFT
eX7YQOmVNqi5cgVvwUV8+RavYJpORFC2B7KUfonY7wcqrnsedPE82E2SczidnpUV
78kp10KWeLc/9VB2SyySmHtaiBfe1U19ilJdQkNtpab/fUc9poYJT7LOXuLYlSst
dAOXqZPBOwsYqdsSgDlzOCHIW11AqhjZu4UAQh+bEeIE7Fy1OP3ROAugpc2DckXs
TEYVBQob20YAmP+vujwlJuiqWSDkvkkfJIBlvJctvTjJuo6XZXhyFOm8dWxL8dzi
GG56mN9LmwqO1W02GCMOM93JSE/pSSR6nfBk6vXbO4RGRT/begdDUAE/w+i2apr5
ieCCZJ9cNG5dEMfts24EFQ9A5fuXNNap3N34/Ciy4wqBJD59RxTnZoDGvL89ACD6
PqcwU1oCiK5BuCMExOE86utvHscECGgrwsQecaTqSV496mx1VxlXkPV9QbpXZ/2A
wYQiinXMatBP/TA15lCn3ecVZX95OTaOP264yWp3C5YXaxoPqxF/eb4azR56zk8N
FunN989KsrWLVKT1nhlwoMuIDpSLH6qlQiCoSnNlsXshZ/7TxXhv6e+wuH8S/F8g
V8yNyZwhVb3aNESFjOPopwkfzoF9KoQ5271RFXHdG4Kdm5Lv9nS3gYW/i06cPHVo
g86u9FG+LagKkJXwrUja6xPz9Upkm+1K3mzRzT8ghrNDTnnpTkWkn81TlNp4wfu6
RF+5QBqXyGyImhlQQmJSAaxcid7SUMAVpDwd/s+wwVlMSn0YKFckZABGbk6d2OGi
5/KM8vtdy5sirukT6vgLv54DcAExlIUjqd+uBbQ6NFwBYvVej+6x/VdKLmLwUI5S
KnDXoEfpWfF/rsWdvVsLq/b3wi6jkF5f4JQsBVkINZ0gMBdCDzJhNPaJuHmy6d6N
keTmKFDRKF8VuxlPqMkFrzLjrisiQCeiEGycLUrYFAzgF1NpwZbY1sQ5Nzf5Mvi1
1+RIwIpHVZDjmQPvyVY/3/UEkc7f/75Xywh2Lfpeoy0W9ZqP/FLAmhqQ8ACsc8mQ
WiVLgBLG4qLyaVAFd4CMXDT11ayApti9s3BtePks335MqRvwwnREfn2Ww4sWshXn
ww7hpNRhbds1e8wKLxtOlxVZ0Om9BFiBM2ljiNIZyWGbNciiEHhr64X3wFv4tPzU
WnurXsKlJKozu5/LjaFbdwcLcg0F65ZVI7uQvaw2/vx1BSgmyBCx84fpIsmtDQnF
fchWRTZl7B9fj2401/vinR4bgmQsxvEwYTSWJcvO1AO5+plydAXGZXWWF9VwNHWI
x54IC0z5SSH//41pEtOJGHETZH5xSNdr6Zh0al7z+7tAthAeqm5ux1GEkKEk0m7L
rl5Obi+oTxycVZyWhZmBbcf99AQ6TtFmtHTvjmY6mvKLffGi1oPZRHd8lqlQRbYH
QbETR35nwl6YDO+0jy9mImzRjsn/2lWf0AyDsfmdqyY2qpkUq2RO+Xdtgc3si0VJ
HoEg4o2EbjqQeXy4cMLbSCyvZwFIz8BZ8SwaRBMX9UruaVYk2uqSm68F+xMDTKBw
hhkJYkiZVnAUKr2tA9GZzrwJ40vapAD7xLdtb+GavL5YtRKBxIGz5ymo/cz/nKft
VxM7fkvxVguJ+OfYuSZNijiHGtU1yntRcHtJmO834ZLUBoE0EFnkLRqMmCIrBFT8
yX/yIfnYL1Q42lv2G7uAdZPOsf+nKGde/bLaC1WM8+NoP2DpKrr1sPY6FbMfsSjh
Nd5phuHJY8SNWSurdE/t0ph/zWA0Tjae5MiHvcok7r+0B5AEDSqyCLtVHtlT7izr
qWf2cwzu0aJWcalLsGMv4MSIBwQTVWmZFTTUD7UnQAaEqtqtaeqjHeH+jK3C6V+Z
99r3dfBzS81YYJnOWpuS5KsvGX2SjsyxyD/0WYvvM91kEa5q+d7wHl6r8s4fQDEm
Z/wQh4/IeBecGlyBXaK2ig+NeH118zbU41YFUfiO5f4qlXxZO5qjfeZDv4JzWfsg
DNzOrh4jBZNtDhfS0vQ1hjqecf/Sd/2xfe+IVirWniUftEXDk4VqlrjIgvCjUmKx
pILblJmzB5pO9oEA84ppHTzgjU8/OKBDx3n+Elas3tJg88amA5GI/rt4d47VijSR
kgXE5Eiwhsu+KCs0C7OInH2irzOVwePXmUIUAvEe62aRV40LNHSWMXi3mx5c3KZT
ZchqlBX7nopd29wpXjlJ7/jtp5ltNxZ/nEaP3/AIywUAsm8BJDCGm9MqwQq44/Kk
ULCy1VxmkM8JLPTF/3PdDqO95DMsjf4jtUHqYibMa3uVTPg9tfBm2wu2Th7WAcm4
pwt1jrVr0dhC+2PpY/DDYWRnJZ1+vD3tqfAZ51cHvquyOKPNk3OLA2q8BcayYcpY
tLovRStf8RHxCjoNudgax5XyOXe2d+yn8ceHxleG+uLD7Ufu8TYu2brvD/WLawNu
58YghQDau3iKMfT5ObW8SNuLUNVkvBaHSNBxdSQB0gLIZ5LwUlSrYh76RuumkawZ
fv+tyRK923kLZH0ojSPChccg4gFJbekp+PUXAaNzl3U2JUOzrIn3gV699nKADUqT
+ro1Mf2/UZ2TtjKCHgtrX6+EDPIXnvZyepT5wU/gopsX+X0fuzAGesd+YTj7psnD
jZniIkidkte9n+HCIYMHOYtOswbpBtdZyYL/B7YodoXYP9Z0tHFEtuxv8Bx4YnP9
V4VYsFy3dLirwLhNdtjj3k9q2WC1h/F5RCJ1/MW9y4dL4jq2fAiz6Nz1wHndbTFf
eA9CUYqBg1JpGL24AKmkDgmSfsuS7AoGa6Sq8BjvjGPlh3Ixjt0tNDrEutdCN51d
COFrIsk3q3hh6sWHwtT73RKqL6pY2L0AmkZZByVq4HA5P4oy9vADORFQySxz12w+
glN9E8dYvfLccDINCxThPbpGWhLmDv6Udo6Sv/yKJmzIZqlY03Ifz6huKU2D388U
z0FX7usvWl/Wse+NH2RiyHqYFJqxSDahLg5mPYHa0zPJyAe+qTGNW53wKlfGaBlA
bTd8kX+dCGYcfvD5bTUb6QDdLR8Banrextv/HNOBgXi1lPd7IBQESHsv2T2Grpyz
eblCF/Bzi4Z+dmtpeHQ8VvKcooFNf+Bw7tCEYoSktKNuHlDKGbKvSGi9jkOymA2O
XRndaF2cGSbbboPEZ2HfAFLJK9J3Ombr6WoASQG7bqqPMaM43bi5/v4YQNCg02Oo
bulp09d00gDxH8QFFR2Kjbzzz5MRv0UG5SfXDVTOnjGUjJNobMjhTzTtb6Q6h/2M
T6HPdH/WFQmXVXZ45t0jGHRlhxCI1n4ArAiUTrEPbeh2PMzNJg2x9Z5OgODwmHfz
o6QZ7vqiMuXu+hXeZN7BejaPHx1ssbGNtDXbvzLSJuE/oihazAeV4xSfXOw/v1FH
EwUOGCmRH/Hoi+zSxVNx0tdNscliYYveRbVm9fkEVAr8lzjay8f3D+6LrugBOKvk
uB7ER/joTgS8yHDEvMgqkDZDYeK7tGF3Wchzr1cYIcj+866vwyCqqos221VpJp8d
JVeAE6LfQTHiVcmhW5X+ZrstwXsv9gcDMe2wj/N+Pf9XzkJQMFEBew87Bl4s2+q8
Qjvjsnu+0ggMLepdbzwXx0kSFoxa+arZzHj4BX5AIMk0gd4g/5nnlbyFKp/0N1b1
q4MfSM2xGH7ZVPVmP+J33RgQ4jQN9Fma7Jp3D9QXI1pfI0sPSAecGZJ2tUtNnTgb
Bl+VwOgpRKnI70y/jvjpdu6fhOp7OHE3EHgcafV37/bOpirnxnqiK+e0+p5hUFti
wIi85umJc4gRZe48n8SfD51p/oc3hLtlV5Ic3/ndnP3cPW5OMinlIoiefKsIRTtA
ITXtAJD7423+XkUVIDMhs0K/qIgjrMON43PFS0MrPB5I/8ToQfpUeBQMcB80Dadp
ZmRRpaOaRMoKPa3Mu7Ziv0I385LvkHQgDoTUGc/g6rVtvAURFamNZEZwhzZCc3O5
kN9K5SilhPC2GdTJrQI0hhPtyV7Rsua1hWKZ5Acddmh4hK7huGEG7PYVcXA27FI8
w7qU9NPpEKV4WJVOwFjH6Nd/o6yG7FNEhOjp3uYrtpNXZn/Yf9Py3L2TTMnVJG6E
+XxMeeXAhfwATInAQEurfqUQ66g3uDbsCfx6MfIt+5NDkeIZ8umV1I4zdnsEezFH
BAeWb3BVV9QPrInMn/lFmrLlGd2Jx2OPkArAIbtfYTbBdlXq2pvXyQo5eTIcAPlT
MD0RaDbn+Bp2ofsnr74D+pUZeATR5mmQPoErfMlw5IIKeUoyAEl2ajtcn9aufwaD
TwpfcxbrKtH5TMnVnfD2L1nmg3oreZZztyEEqNk6WGk3k1VwH1rPrI0ObBunP8+u
wmwuWBeZMorueM0qaOr3EdMPDq3dhUDcHmhGNPgutpjTPTbU/fRp4psAZ0NjdozD
EnkaplD1BkTWxq2bremVYhQswpspCQAz4ntiGnMRa29dWUxGWbqa4E9UZ+BKrNG2
EZYlt28ur573Gg3tmKQiQ3tCqFVUnUHsp3oWW3IUU+W+sp1UELziBXLVoPpiRsQN
lQEomNCLI9plOJhYBhEfjUOthAuVuVQxN3uUBePhF5GSExmaroo/2pw2hl+xpe6c
wUn8k30Q1Uyn/DRDaQufq5jaRO8K8bnrN+n5329pqDUv4GeZxdzwpw0OQq2tk6kq
nAspdDzIhVBDrDMZF4l7ozGY5vi1rIymyw1GimBL1Cdz7cIWPmCS7qkkmEcfitY+
9CgjWklUl4c764SbP0uagodOyd1oZrBdONgBfu/BryASeoPAn2y95chQQsWQlwMu
94fmJaJ2xrzkNeX/yx+tAnLfIobYnrjh0kP2w4OtPcKVDal0tS9AwUwp780qahK7
o0qLpVOaTSWPTQuhbunPYjBhl9V2BHr9WaCcY5Kw1p5jL6vJi8MnAcGgaupwP2qZ
l/vsp/cewSr7ttfzUkrdQeG2G7XQ4jb0stI9KxI+NUVYKtKl96UFZZOj4YgZBbZU
seo+KNnvVGOw994kCpq2u9O/bw6IMW4LtBADaBLf6jpqwCugiBhs7mxsn4tINN+R
Y6bccOgrp91GJ1N1rWphJf13lmfTbjgIbjmmqELljWnj3fhxEZBPaVcZFhSREwaa
gAwWGndMlSsUisO6wnKOXxb5zaf+0Q7RPa4aDF3jrNtSjSnWM48X5zqFhhpWscRq
T1nHKPFYcfV3X/HObGQ6TiLvCX4s8wJyJwiZPQ98V5j3arhEc0hnfG2Bf6F1Bxnh
J68bBj9hEWmnv2op6DHn1xJiA/uY1DrnrUteAdvv6ZZpYc8uCSaWkQK0wGfxAVfA
oVjKadUgbZHSJSMIzTBbwd/bQr3jzP6rSwXmw9ruYWD7XZiQ6DD/aJ124NlO88Vh
609Bi1StBLtmcKhamLUhaT/lUutsyhbIqPEzFfdJiDtY9LqUN0Uzs7Hob9JFi8jx
RUuY5b6cqmyzOQVU1AXajPolSDSNsj6KqgY8riWomr8CDGbc4P0PvXD0F9JD7mUR
p7LaXVNkV1X2sHG2nKsUScIpH95Y7so7AwnKfheXgl1jZzxx7jaKUANTPGECUpXV
xJPmsj+hcbyWms3L7WP3Cmq5XTAelaNt88wkwShBjQaFLPCnLQA/j3niq1PrnkdJ
CIQoDl1vVQpyON4dWlEyWxuXZEVfktMgRjrKoamOFuhJbLmQLuXVmLGIecJpWY+E
nfhcRSkyKzmjTOvvR08WO5+eFUvOCH+iGUqjyfuxr9dyDSazZmAh+UpDi+rv4NaK
xQnATwKVP3QN8su6O5qIuzVgYrasXbSGajXWPLF5udCDCiH231c/bhbbJhjHBDVq
oCUjt9U5OkgtuL+g2Gx7+9DGTXgo/VZf0y/7TFQDjp7c1Rw4qKu4x4YL5fxuy7ld
kLjoxvSpVsZmDGbgJ9S8n1e+rDLlPmuzXlxj9hZ2KQPzyxF3zYm7rHTbRhaMZomT
lELtp4JvegcyrwW0Ma7pOyNnyM63U8w9SoEWsTclY6Go7X0MzFuro3GLnfklTQx9
oKIKiJFGAmEk7RbFQ1lNfHf7oV2q2k6hUnnEX197HCE/00YZAbO0nXJ4DRU/zZrH
/ZvG/ZbOsWxR/TphlblMfbbXmN1+ln6kyfkXtR11dEgQDMzaV0Dm0lZcxHvowB7g
9+h2mOFpLqOj9tBofBg3Bzoa4FEXOItPFNsZymlTy3jHZdfCb0/BOcAMWnd+Tif+
aXiJZs/Q8NM03k+Zk8ss9HJZUSd9y7BpWYwyYDnDz/RWbzNgICjCeJ30wWNHzOZa
/KkFJYpXinm5V8CaGZo58B3N2gyXVZMAMcLpTk8QNuhJncCXVZ9DQVjs3xpkDAfI
+v0fT2SMWTEV40+izrIUJh5C5hbcyY9StNDRm99jJm40mwbcAMG+XEab0iU/2vg6
QhdV1dD6n3LqeAkufVNePVGFLhz4tCtwx90AElNo4VxXyRFr8MOuFDwJOyF+V+g0
3+bH+vE7DHKmPY7npF15x0cNbSLSaoQvJ5TKFR0nKnDwhV5mQ0VmeCBFQOYW5QVn
kmEOR0GFl7KsntKmLmLc+aDtWOu/M0S53Jeh4LtbuzBU6Wchd/XpJepH5EMd9O+Z
4HWjKETSek1NxVDCv80GpvuWAAXTcdlX2m8SinqgTfQLyqBtM/R3SHyOe2STWjIm
TgR9kFlP8Q9lual+byFuc5i+GQSQypBUbo6hkyqdBX6MTqZqAYRGb4XT2TAd270l
4CprCHHg4jFShQU1e4vnoERPWLU+7f5Exo0qYOp7DFnVGaxaOrjUXpYBLPdilBQv
0ZRXgOEfHz2UbTGFXaql2j7PxXaaE1TFzCjdwCOOjWRTARmGF/JIVVZkkSKHVouN
DsIlGxhoodotrbZIXC+n4BvIfobkRSXMos7HAbpZ7uORC+AnPE92dUoSuLZPho7o
vqag+J+ZgOE6jvqqLL1/b0qe/YvpOZgE4u/ydTmL78csUI3Rj4pRcnh9eFFRlw7s
FKOX5Vw90rFTRdLXHKp0N4jP7ZZEFgFFlsn0m+s7YjdDRKiaQBP9XcuDjd7lrocU
a4KVVDkCGytCkEzaXaoTZVFRsVoQsppOkqm1MxwId13OFAdRKxUo5KEGSjWTNnuu
QEe3cBzVF2OwlhS+o/0pXoRpvF1wjBZ6KX/1Myq4sMN0RPs9AhR9av94mnZz7gHt
wI0cYNhI3ufT6sGMpe6SdCie5fzxt3uqa1jbuJvn1LFAXmVBVQT+y8FiSmDTv44j
SKFnB1upu+Jkh8NWeryKJ9tR5s81B8XRuqg/kcMDC+dt1m81Gwsa9xX2rWUgcg+B
tnYOT6nlk+UbCsbm1Dy6PyTel+ZeoWdqiJH/R8jE2mOMIEiWJMEi2JKbNBUO2Q+E
g+8/mkZj1xcSDa0M8YpasLFmHJnlUMoul8v/UcoowOVsATyJSFow0JZw2rYX7FmV
djox7ue5CgtZJSwhugJnk8AeqsvBKoohUpe7UNb/iy1YWMUpIf7Nz1B9RrLWUQjG
nTQ+JSbAp4VDw9Oa4VV+iivIaeLzP3zyEtLQwTD0RqSkDL/4B5va88ftgiBdqdGa
+zHSVkqfiHj5a+wVmy1PmC4YeLpjqXAnnqdqvKBLNvsuOVQoujMvi/+enDLtoNkH
kTmFdiPfInxX0hRYZMQsYJJ+JAOw0Sp0hiZwWlAZjQlQEdSGIJLZZJQvb6vrTasc
fCk3i+x4wCt5kTKN83IeMXSAUmM7scPzCmahIzDTyIoyrvRMgiNfy5ggtO9PxXxu
EwaLdzGUOfIkXhAfkXTYPow7KL71lhihwJC9HXD0Ud2GdWzmfkTnG25GKp+pxutR
XvR3/iq3tUuVhjcnRC8Aw6gsI6wbMizQ+baMc9mrvkTWRNZ1e/K9beQ0lcFi1A2Q
I9m6ZNG+SsKjHvZBVpuIU7AWj6OBxRn8oy0UKApWG5xgooIm4exMgY0QOS3Y6+K0
XRXldTC2xXwwfo+hpI0iBNg97YQnR7yxLNIJz+FNfYRO5It9IYZDqpuzKgQwW+fk
rAl0bH4KZ97c9v30XHJudkH+ECs5r7LVvoKqZfJ99J9u2NeqfmQ4RXlF/8VBnCe0
G6X/vUAi6Pa48SzJFQ39L/UN/QmOozUsH/KSEoPBOvEXrPZdj5BF+h7k4OCMiWTg
D5/AFy3O7C7wphewRjElKjpFsnR0SWo0bXaAVW3eOicKdxfcnm/NDqMDOa/T11Rw
/g87Hennd2J7S3+Ye5hnTAR1NMo5cWXlGmqZb+05MeHudOVfnjqzEAkZkoXINK8v
KY93q0IVYYJ/ve39+mQjmg5Qz+c6oRbS35O3uswabmOKY+Gzm2Q1NfixwhnHzsMo
VMpM2hQLUEa3oP5eiuxf5KJo2R/bq6zrfTGc1ELvv46hXMm3SKBvCRj1HoTmjYog
bBGUvojVXze3yg9ffbLjvVqCSgky+4/atcJx7LGsoXyuJudC1h6BE4KNmo0OTV6F
9dI8H6ZS7RZadmtje6LScMNxrp6W24s9F78G3gFxoUCdaFbLo+530sI+mRFSwLZ5
D+WsIee+7teb9u6mYBO0tA==
`pragma protect end_protected
