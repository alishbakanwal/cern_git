// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 13:57:48 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ghqTPpAySkq675xiw84wkUth9hLNTdoFZqGknSjlr0EFfcYrRqWbB5I0lOPW6LpK
WR87kFCKPeZXEDw3ZdjKC1+PDgDLGwRnX6LEVyOV4xV4H2u4Ovkxxj4EwUNEScOu
CiPR2YBTrLuDio0sgwTa745HPbT0UfJC7HxUvzVfyYs=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 57760)
uH+SgQc8R6ZTcR4WmZU9PTgDSxZ+vphnXeAgwZGeMXwMdu+9uJXaeSrgWr5XF8nr
mRVCcNINzpEE7IoR95lUn5zvb33Um51WFZQnDHX8XaD4hClS/XBLZ6nDwtF1Tryn
v/XIMG9NHkGrjPJZ5aMmWHb428guLF3nhkQK0wGxXoRqxYFWIYcJ1g4hArGGbfhy
RGp/3j6LAhZz2cdCCxFX3DZqnLMzerfNo4ZVMzgOhpp+H98KI4RUAutFQP/ZPCec
sKb/ckHCunfs7pTsJYeoB1vefkk/0doa2A2CjRbNXIDz/WMDLmFkQ4xUs3lGIle7
vVBtrygLLOKL/jLeHsBUhtgREkpY/Gp5egynm6kS1xPOH8VXfJE1X4YmCM6u/lHI
h4mivoNOvGjEV74dVV2nyMPo9pxkkxk9RTer4A8HAFScIqVvbv4Taqzf8A7+Q2Ue
WleccCD+Ads0sjCjkLhKZ07aNgUAbzYYRG/GS/0Cri0c54+17sZnhhOhPI/gAVxf
aM48IR2I6P4TWq/0KZUf3IlK3DZBWKUm2DUOMw5qRF9omo2xYXGk88OFghje1h2g
PUSG5qVmyUHqzivBz/+5PVpLlZK4Vib9bN5UR3X9xkD0GL2HCjW8UG72NCQ7CBow
3FGMZ3VQbQz9MiXPtD77k7TGfPRgIufI7Rp1ilriGcBr+e56vgEwpgHcv9CeZrcE
hYwopk6UJVzWbTYtMzjsi5798NhGQsSPpz34o1hKmihnZ81i7ByhZ983iZjXKPts
h8AowZ2b2NzpI9jqciNFGnQ6ZE1xnkoWNIXSWSuOg8l6ktgjCcCPbUhOOgJ5NU6w
eGHKzQ71/TwV9re7gOoSf4OPNgz1ZrfNz2Z7IypzyXUyilq1FzSniRW/Id6SL3/h
3OTK0d4/13Mw8U2/u3LI/lQwcA04x1YYg9MAB2BlRBhyZ8dP0CTNCv4iMawQHxfR
Jq1r3g0Vhe0nthfQ86S3bqJY3KOFKzw4GSTjp8RWFZ0N8Pa/vdguPZYhDGGMknED
kKqeCkDrf1BYXKvrPgtjY3I/PL3suOn5Ak5ZVyUB+ZN0TfnlsQrpLvTtEfS/Nmp7
bOJyg7SSu4jNqLKhnS92HhlEJ/wi6haDC6Kmg8XokAaOU4oP3sLeOTmwv3gziLkB
NvKRy3bC2O9hcHuiXUhJRRSCvl7CcxdYl7N+QHklQyfPX04nF098gMSVwzZtVuQl
w2HGEsIRVO7V2eBOZ4LqlTDfrnseODpFFDc4VbNoCIiYRiOikl5dz39R9daETXhj
7vCDeReo84cg3+7LRwKZ2952TT5rpebYsf4Pw3da2Tz50uvtbwd2HsDjMcm4SVFO
JzS2LFp7VCzI6/LB3he6NiBZgGSoL5WEDFLsPdOAquUx/Gc3iCm9zAwoutadmwzv
AQYFC8SXyMeg83akGH88mWVrC65fCBUTsBjgnJ3eLR4O3u6jwxnkdBeICQdsX8pv
k33bWTCdthkKQ4pqIZlU6xT8/km2C9KAmyjfsIfptx1/WXmVXw1j8+trXr4XvRIs
O1AluwkxhWqMOr7KbwFnsA/MfYkti/WktmDZE+2quwxdPg255UUAqnbYUixpMqc7
tQoSfODwwSBIq+MAoWuy4TQZgZQKH4/ZmK9j/zMm0m5aEK6+aXjqGfLt2CiRDEXQ
iZj0kPasqMTac7Z8I26J/mnJxXF70DufVaFymhdGLccWUDKlLzM0Tp04Vcpd6e5K
tAIf2Ua9PosgYxRblGR9D02UBiARsS7KHLtvssWo0MQ2Br1ufDqs6HJgZ7NFXlNQ
MuaOcsKycWRXKqUds/AbmNrYTXNC+0WB09pjexElYy8b2EwuSW1zX5BkZPxwr767
1R8YH+hRm7GM2CVKOC7T9rB1yEj6oNfql7DdDyXRBzLKBN7XGkjhulbcxSSeNyzx
VyFwy2oppQjFDdlup2EdO301LXFPalbc6NzqstJ8NEMp9QdbnCi+k2AgAIhL/N8o
B11sMznP0H7Qblqn0SqhWL/VKU7XWTVUDiDy1UEv/tI9hyw7XHw3IcDv/AK0ljwf
PNBxocHWwwfsbdRpFU1CzWSiqJbERFCmjQcnc0jZPalPJ5zxInLXQWjN/MCYChCG
UoeCFPnvauP+pUQqU8qWWX91Srv1rD7LOqgGeSk7OjNbG8hDMmptg4uhKG/A5hYN
DOgFhJXHTN0YUCZEH3C7SKzarzS4jgwg9DGHzr1TO+QDrgcoCMrIeB5pgxI3fjbj
vFipvSp84GvRnqs4edaXlH7JGXb6A+F6z05pFOpTOQq2z4uANL0t1rpoTAHrS/mM
ZAbmaj7Yudawu/fS/12gwqgjSxbWJMzzRxBd+ljv0MtOt1q5FQfctO5FZpAEEU4t
NjYv1YLva+5sxZ3CO9ucUC8E9d9kXaFKoijicx6Dny6b9V0OVFFkpP/bRy14FphK
FtUZDD9fQE0F6u+9w+JAVJup5bATEtveIPwSqUER4N1WLP+SPpjicYMEoU8n6/ro
KUs2gUPUN5cDMN11bx8Ener+ga3c+Pz3gyhSXj6SlWtnfmkv6pqV2SSvqdup3avB
hHOxsQ1/mU2sAtePtmNQikieI+nGpyI7aSU/QT7BmOb8miDSVzGlFDffj3P2Vpe0
mG2F8ENctVJ56cjjQcdjBD8HiwXZaOVed4HOx0HmL7jg4pfxipQXCWIoVaBz78j1
277GWkwYQhCF/kLAH4aYX5j6dSqocxeD164hS51dH7Ozr8bcEVwhjb9Y+VgQ5Euv
XqolpHr18We2dhoip08Jb/A3UcFvve/AxtWfFrBWBlRD4Kc1HdwYjhomvUoggejk
n4Qj6w1OhIsfGylzuXMadzMLDPe9AUbFQ7e/xM5hvWUh+2RNuMeHVlLqlRu2PJNn
2uMllBMoYOedfSS/Om6888aR7O8sVBYHOhTHno5vdne1ZYITFYw4owtLTmhKNJkj
OQ78+dkX1n7DyzWBpjN4odfua5v6FkrXFLcHibmdVptMurJmm2OLdKHcl6Exozg6
B8UQ6i5Lz/FWtdkQYH0ODGiUn/2m+Tmy7dIEBxGb8N4D88z0eRlxEZ8QAUH2bXLg
V8wSaVAJZXT1IGII382dgGXCUTrPJmiSCYQr+gtNKZEFfTh8c4r+J5xINXBUHmi5
pfyL3UGn5riz7TJTjkKLw8265Kxdkp6r7xf4aBkjtrv6iqlbzWOCjSB4DmeNsfXQ
fIG2A/zP1YUqVBvw6l7aurr1iF4eqJ8wCT6rTrXXMkoRkHVF0PP0zbaRP1XgucNn
5OS5pHOeTO8kFv5JCzGqhC24RR1tar3YHl5B/l/KQfQhpVo0c4HH+V9CK62Bql0S
MAtzJvOz2OEepPZ3JTqEHREMVb4M/cMYTJl0fqNCO+qHYGqprcFp9nDca8QmGxuB
QVvCIbLN7eeoqk+Bm+65UupmKHD489zjVUh60mwMMKPVJPBGZQxKOFOwQnB8aJfL
+iSUoWrlZzGi5u1z2TMifSyb6BIDA3pRTjg9Tge27Xwe8EPvc6d41AGUwPpzSlbL
u+UL5EvlmN81ZB56nCng3n/0JOURq9BWzJDUUoe8AUpTZSCnvAA0NV/PWO0BaToC
8zNTAtq1XY3G4Cc9T7al/AWWKR/G5s6eQPF/Arn3cZONceCQ8i2nD6ArYRsqkGe3
i4Flml9jQq5CjTVEjQo9GKFn/xmKcu8rgNlgSCJ78SuZKZzUi4zkzVU0KTnUMgiw
fmleCm/j/XNOuLKNV4wBMA7g7YgAm+vcI5kzOYagf36QYRJtZqdhltED9zimlEAy
iUN0Pp5WHMy31jR5+8foaH/oLWIl1CzMH+8y0Z/E8L5eKyciW4lSL8W5k0CvmvoX
zKqRpiy3rI7kiClAQTOM+Nv3M/puKuEq3vZw3gsE6KbETdxcwkWNhAaBXMJTh7zq
fQsNazxxflQSF/dgrL26EqduYZUlsoPiTiH7PlNbb4AVo8ofQ8ms8RSCR1iw1dK5
KBnQ98GqpdX1YrB0pd4LI+f5Mr4y7Kqw2O8RjJ79kTyM3u85wLCbqce0Fctj9Cxf
7LFH3VwejKPxMqTUgrfKuJhqIFs4X9QPguJvWzCppQkDehC73ey/MX+V/IGNMoRv
1gcIYGT4kKFwE+SkYY0C5mLk3/auI8stm22uVH+mbqD2ibfEovU8i7GbZ3xijrme
p3gtRB86VfPZIewpRuaPi6epSLdCjkiH8OxZsx7dYr0bPf14AD7AaPJEgC7MothR
gkXINX3nSe8JXkCutY2zcXJ0DetIWd9B96Xr0RCz0LWHyZpQRTj7drOLmxSSAMZ3
nnXabSzVGJ0kxF2kH6BZJiXwAyg7NJRAFxxbIumfTRBuw8BkiUZsalK2WoFUJOJM
1/sG5rHkLKro2v0KVZGiRL3OD/It4dkHYu6rD3Qr/LkeR56pbQn/Ultmgrrei23D
7KGiVWuywfoiknw51MPHY01SLAWM6vRtA0h2e3qA+6x2hL+14KDGW5Ii0R57Pyrt
yGdSvFTVZVeBdRbp6Xn2oiwfOr7cxnwuL8scTNdyl+k6xd4IU+DBDsWdrIEsYePE
WU0NoFXksEkp/UxqFaCFfadQ324/oHkyq8timaPGFwDdgTcH7Hw+gyitKWO51RIW
JRMn7ot58MJyHi7HVfrYwFCQE8VQDq9G8C5dDj1FnTRsfn4hHUnBhTM4WnkeMHyG
spQKBisPiV8pVSKFBlktEHddwfgnPLoYiQv4XeCrz8BjEXrdM4r/DuB2O7U4yXar
H0olYqw0H58BwftqKlByuMNywk7OAUrAzPbRuLSF6iUrFvRkG3h+O3dcuLMZ2vvS
uyoowr6NMtncpNznftb2OqpXo38AwR3mlyXZP4umfqeO0Jx2b/AybL5b2TTNeXBA
q/6bHyYHieXloBd38JZMeKfSFlEHx6dKzm3i7Pvn2XoBl+DiIl7U/aja7e9jS5DQ
es1HbrS1K/vQMU/6zbEl1h3KmGB9KsHXHF3d0sFHcuAFgVxYxWT5/cejTqBAfAnO
pbI+5unlARx4gt4yW+5LC+1r5ZV8s8GaqOEiXkcX3VbUl39RSw/iUu93HOpuv2Kn
adKd7YnHs+cv8F3GCybCgrZ54/wFQDjXpF1T3kTdXDdm1YNjEfGLpsl05rMOv0Q8
QPqY1OPZoSjAqFOsAkvVInuSKEC8Q4Jw3R6dVJ7+gqGRjrP3x7DiDImms7Byxdz0
W4HLuPWwzUR9lUapG0kuRROk4X4eLqXY5n0KRpIksi4lYbowNsX91nQGJGxHv7qj
r3lUwro2anmc7g8an4qcU3MvqSfuQy0ZOIzukkZ83S1+YAT49dZ6ieuMqC99zCDZ
zs/1EUcUcKLZ02iINW78ul1bdeK6sRi+U1apaG7cIeMGoYdQTtR/cE6g8fK0WUQ5
17IBrltXccHU6QeiYXJNv0ZgngzgfKBqK61H2rX3av2G6Nj+leVhF9whxxNKvX8d
LDGeLXzBis1t10P67CPk17dZ4HMbBAJUhc+NiLXYNNQ9/OLvuDlwo3MmPSI8E3rC
6sOa8LMELGp0GsaRhUx5RVssLimVh2Ztni4XpTAziaJXqWWZb5ykpGaU4pGC10aR
2BAnTvm8wyo0Dkz4L7h5pwjVmN20Dadie8ApldBxCosRbG23tYoHNj9JcyaBU8AL
238W9xZDKlWhG4dR+r7zISumSmvXlXUzGTA25QQs7u6V3MZip3+HKoT3MP0k8oK+
2120YSOmINmgTipadm3uC2PnDuYqvHwZgNRXP6/LA5WGehoBKrJvoHXM6OeHiO4o
be4Pbeq+zEZOyV2P5Eykt3OMNGkOGqBxsq6xMZzjst0/cLcPLxvqN3EeU2EYT1EK
Hqe/3tOn4ExnZa9ZbtRPRvh89fh85gUQyuGKfD411lDiiiD2QSCfceV6niyxXTf8
NEoBwQCWbMy8g7jfwa1D1mgrtM2kHM71UwMhxq2/2qdIpoTem4CaEH4M8DUirKr5
Fa0Mub9Fag1Dii26piQV9WWQ5x4CvGp4av6o431VKl/JQySmhe9XI9p+IMgWWq1W
v2TYttpsIu0fX/JfCkbQw63bkIpLfAdOW5mOZhmUDqoAccb1zVekaoBvKkRkGSM5
XbZo932SJ0s0s2JJ+mb3X/l8LK5MLLK+dpb5LXgUqYvmzJ9FMtRiP79Wn+TRBLUg
rFSnSnVPzeQ1Am/J6KnwUP3bowEjXcyIWFTqJ2rvkASBm/ESPRM/PgIyNxmBMEr4
mGvjNBg2Gbm1ZHDTlw2ul2ZaCE3rkT2hEWQGRyKMbyb7AUq2LhgIvS+p0ZZc5+IY
2iZNEQLYUpL9NOtDwi3enNrqvojyMF9asg2r6VS0AMZDd/c6wM4Ks7G1V+exUzcp
lfcqK9UDn8awKHm1rmhUfTLgYPBJdXUes96fDJOQ+XMvKigqplf5PAGuL2rKluFd
pDSM44aNuu+1XoaZxHyzATNws35NF6hYMXbfS34aPfA0rOJIYDftv3yEtjdKrmLT
+v6G8vZRwsegW7Ojt8INxY1iJFbVTueXyAoh0X5a/gJsAMfRKSC0N3ngrlgBvmfh
skOS3/NFopol+HCuJgU15p0iEkI4LTifo2d9UE/y1Q9KoR+jhTfLNwfVxd298g7w
aQWzC6rqvCwR7PXBAM9HMqThSVTUCnvjxlenai9Jpr5kYCT5DKK/wirmLfNSc6O/
GvlZOtdGn7dZwXhsrJXg2/krtXHPG4fYQ5Udj587n+yXC8+6Xe6OpnX1vSFJO6Z8
eKnuVVBRU5YVPdanpkNiQIk/nr4ZXBKW7dkriIKn4nX9TS3UpddOq/B47yVa60+F
CykSR4iZBkS6onpP4ECbX4dpO5jIEPwKl/HF3w/+zDrH5ilNspWxLWBTlmrDHAx+
eNscolQ1qrsQYKf69HwWLwOoSXEMOLnhK3ZjvXw+uMQ5pDuglcv2v7/ErzuJ+5+R
8XLnCow/GYwipTAcjRKZzAKJ277Ob3ptrTZmF1Z30usg5PJQwVVvB8miUaHXzCTC
lV9rBjl0RN4xQGHjtmabqYWqFV9bM0Ssg6OKfkMZzvRKQpL+u9lbpIP90SQ7/hjT
KtqS0wt1CD3LtKScz5StXFCKMGrikHF368WH1Qbvo7tsOq2L5W9PyxrgxF6FpX5S
NxP0kQHYfxbDHENZqlhmugm3OZvQGQaWHfd3Nb798LFyS9GiRZbwPLQfQ1Abfe8d
2M9+5QLKxNgUzlA4ENMCayyLlLccxrqIx/lxUdov7ghVR/nYM9RpwXsimVcNTw7p
uXVMUPHeu4QOTwK5XdLUlRbI4sWxEshEgJm5qOfo43bNkRgjtqvIfODjElKFBp6I
sw3K+XfkiaJYWcwUewuVRU27RPuLpDbRmryVWFJeSQHo8u2JeMIk4g92kl+6z89D
rKKSgNhjPs4qzhPA6HrPcBe5WWAx0c22hh0e3nyRqP9TpBwG0ZGhD4fIw0lvEwj+
0gESabBGHNpMz8rJCkpPAwL4XUkg2WCdWJk1YFP5W9HWvf2q2weQo35jk+/NSCsG
z+La2Ue6aut265YY0KxdnARG6ehcywyVCwNHHJhSQpCOPEhM/ai44YrBA3SjEnWP
zT6WfvbnY2SzsRBEMtXlgCNQf8RRv0ouppLDtm01OrEFSZyrCB4iQpZ/hd3MMJ1x
pmm5A9j6cfCmGU/CxW5ZHUuIp9HEKfLUtvjMN8Tvk+eg5NZGR3xGfXfHku6v7Z1u
df2OhOiRQ1GtD+x0JRTritbwhQj0mop+BcvUQXDiQ1z1Hl92KxCtVcmCNAobNYTD
yv8j0avgzRybW8lq0C9ioCmYOb+ATNGMfztv89nvf3nGQtKjPYaHJkaPoVpwxFeJ
8TwMhQpHkeqyc+qy3pcuyB4p2ZAUgrKGQ4Y8pCvVeqMxJobk2cBrz9yBQsIGMcQ7
IaE3RGBLq+Kmx93KeoS4e+71z09q2R9V7sNWAMyhl6mUxMxPrDTkY7LOgvFaqiAe
1GMVueIwittGxWKvN9CyXEKBJdab+UMZCtg3Ga27YlcxlQGeZtsES4NETVOsz5Rp
FcoPtC8qv0oNMq1Cqhp8YJDXPj3HUmIc2U5Z2eKfGadRShR5tJNsu3UE1J8oe0u9
MN7oD/geFIA2ouLVX0KO26jzl5YXgdVfScP1gj2ftobl3JPDyP4SJOnNCze9av2i
HhI+7+vN3kxqCV/N6kD8meAcLCliL0vZH+/7cEL/wSdqmtpUiPxyfBacA8pk4aTT
Rk+h9/phEoC2pDXxzZemh8HUOF07Fz3qoQJnz8y9/nONOn3vuhwUoLxhGB+hyNmH
U0QtClXvH237Hro9bX7EDnCx9FL2VI1dFeDBnbxviZIj4LabLULPnTbRhLrG52Pp
JCRH86/iihCTeIAhe2mdkMvyrEp+8jU0fAZJjbdch+cyLz2AdAjr9oC2eHHYzmfa
ipdp5l5k9r6GsR0OgpCfAE28MiUjZDG3SoUqMBUY51PdsaS9jbwV/8pcSJTmqavu
2hwZNKrzhw9X90r4tMDQ857Jmn92VMHum65YaMAVwZ7ja+EkavIIrlWAgd+26fa/
lYIZQIRjvv+46u65e5At1uOL/OVu7OLMtMlcLSiqEG2S8Qv0mKkKqMbnttQKxDbE
wbLYEeGK2o3+Hq4Nqu1spFgUF++xyPgBvxGlmPp5Xw2RMC8slFtnJSyEkm3YkGdH
yg7jsrJen79th8RhLQyo2Loz5FAWFN1AEr+D3UrGTC6KS3ujSvexW3U2VTH2AacP
jnRCrlwEaK0na+DoXrdtPbGyeTmcKArnGpIUNeZzfweiTrmYJeHy0tB9cEvLbNZB
tnrPth6Xz05JSIpFAUKbG4KQKgDG6CQCRh1z6sTwUPCzS1bxdM6oc9Dwq69d/jmW
6RslX8Lus1VL9ZFOhJBhRUNSONcDThc1+VEh22r2E22NF88fHIgM8LeXvy6SDrtm
1PZdDdj1BCIpuIxPimjZmgv4BlURNK757TzerPL9fKFTlvg4C8lxV5RtF0DfZiHh
MwC+Jn/FYTvLPu9SJLDw7DRLq3YCcZBcqEsikCo753M+RzCSt7nS8FgxffCZzorV
zq6UeTUnKSleKxHMMb0dsmf2UEyxXX0tfmxqEJPfJthqY/Na3zyory5Bwkj7COUR
FhGG6EkGS1jIjyF1o9ihIEilBMi9kRts7gH6RojpIky3XVJjH1Gw5w1uEhk7lN52
OHtxEd0vYR8tWlAeL2TRDWxxzKeyb5q9qwfiWwUFgJIRqaDoshXqb7IGGbjTmyCM
lu3RO3XvOFwg9TLMDCl7H5oVwDwVAFbWO1ENWQqe4JxV0KZqJL79st5LVAT4H2FL
WqYZ723UI4cMT6VJHAUxjRDl4gTCwb7ADqxNA0RSSYkbXoIgU32Z354iGn72Id64
qBaINm44LEUuzbiDKrw+C/2tcPBxjNNTQd9lvCuYZwLKvMFjf/IFmGqGccGb6UEd
J9kJ6hAGj7D/L5MmRQrepIswWKrSNtKKa6AlERBSi4DQYE0nMNakOPLkN8BhNsxK
oVeSawjDJMfPondKkGvEWjdBLSUs9hqeq1rtVgLd6Jz33EMcwdn53+lzkvB1kClj
q7Q9ldSjX1GaC6wVEOyILqSP+JCU7klZu44pfbEoi9YLbxvCnmhxo7k5SS5vgGoG
t3gb0jYfB7wKaoEQAFm259WHLq8NyyGNPBZW48Ll5k5YZ60V4gVRENFJzs6ZjfjW
3jqS0L7B/YFY8NWJ9nEPnu1ixqsGkVLlF0KCxpzcNyWU2r3Dg4iSAewL0YPaSnoU
nSDHsQWzOG1SM29nQANghGz9Bl8us4tStD7wA79uePnr3SY2xz3E/1H+sjjpeT1F
VIgw4ZPrURCE9X+D86FcctvmNGmVnZicY0M8DY+vlJJ3AHZqRNOyXm4ZalVT+j86
UNzLaBeS1t00qFCsHnsGDhtsqb0MSGFi9gytjzD3yqX7Nf+ZsEavfAvbA/8OgFvL
6QHIxg+rkh6KbBNqQaZHj+ZZ675g02WixFUluObAXen4rfZ6xshqTAtFe3fkbvPC
FDe7dlFneLOi4cgOQn6OX0HPFUBsPZftGc4ysktFfJGqAM9pP2XWoC1Wsf3aD61A
cI/ZsJmdpN2sw+xXLpDYYBHRCK5nDmf2v+1DWXekI1nsDwjXbzPNaDXv2wO54A7u
mjOWDAYd6HwOQ9c8Fmgosuc+GqNeminGU92D7AkERyHa2KNZ8Z1HxRdf5Gerjzng
whNxz28L/M5HkDNu0NFgYaPtNKDZhqRyO+RJE1MW/e3Px6r5kNRmgZg5o3L0dGOK
adl4bds6dqQw63FaZFcrbstr9rPjNSWWiWbTwnxUwKjKgdSmmtB2i22ImEcgE2sa
n/wOMBCrqN1kiBhWad7+ww0LpUUf7H2Rw0SCdSw0sxIqVtm/CRkFQRpD/Iku3ras
jX0cFoI0M/A8VQVkxGdA9y3SvcJfq3ZJ1737IEqxHxXlNeQGoMoNaxzNg7vD8fLi
MHWLdJwl2T3ZhQW/eV6GqBUYGf7ktrW0IBAKq2DoYWeGKXONOWziv/nih/e0wOYH
nWZm6TomB9+x5YQCe88VInEOXjoUd04D3grID5IYbbK30bKaT5H/+9btajx47+K1
rqUZ822GwIUoRwwndFkaCVMWfTTLCwM2JvwI6rnRVjceBwFRVUgzn0DVkvClMZsX
eN4GpPMIYqt84FdR+lb7rCMp1zV9GBgzeEKfyy2tRla/JbikqXT6Z5Z1AKZKy8bL
WmJoVSkDyKwpRfFGhrYM3EQadd/uIxr9QqMUhiJQ93I/GMR0Qhbxrteuyt7hsDH5
mPacmPo5B4ayZgbW3Sv5RnTbVAcaZeD1esQHtyQ/QSQG3NNE4e/ZemN/AMRYmED9
g/jfrvtwOCi1m5qh9j/aowTpy/REApG+UO2E6YDqXmHndIA0QssLoSAcoxe3IjTw
FIPzjk0367BLtrabm26BdSMPsiik3VgE9MBnUVK8gh/XZK3hJdvGhHIC45v2N8Tw
QMlj+1kRy8N4mcTop/4Xbu+aJmAgLbvvLKGXvEWpSIW3BD7pACrOEnc1pV+LvbsD
jKoTkq3U8UHA3S7hT1SA33gZB5yKTaKZdk4GwbjBjSz5UCc3UAOaW2jq9QEJ6oyf
ZVMBu2ZOcBu+uUXV7IyPGA2G5Sg+YYuqN9GEJjEQRKAu7Dbb2F1nRIrzWOMpi4Qf
1PEWlME/1a2NqGnBcOhQs1l7rzWNd4AsKWAocW3sRstARzqfJ0PXij0KLL1rrVYo
Q/tyAPefPSy5MnXWKyxp4DLME+TBbAW4bdAYLcO+x6q6APhU26Chu3pGpxLlQ4Y6
tDrsujrmBxm5DafXmhtG899aoiTJN9pon7tsyLi5j+qEYS+l1oorMaghLsOziHBL
50/aiMfpXA/r+ZtG3CE5MCHYPojCLzCJGV6cRIKtqo7QBAUsub2bQf+/evm3jhan
VWJm4VlRqge5Tg8aqUwzl9TLDjBR1xIAOWzRK+F2GU2hx+nKmdNAz9n3Z3bsEMa4
s61FjX4Xv0w7JEAvBtxFWEl7zwSNFsyvhxqvS/jwT50Y7Vg46rbVrPnpyYZaYag1
UNHd3YcG2BrzAv89XFJhDbhmAoSFUfogq6iVDdFYRSjW14pIxyO4OpR2Mp+YdCkD
2Z4K+j5GQPGzqonKBlw72WXVxK0IoJuiH4BJpFBU0d3LNnAT2WP7wkpaEq/8/VdG
kHelgwvW+//htSWMMFIOSK5LD9QXB83pVSJQpwzzT5h0wasuTS63QocdUXs/AcnD
TcMAFBp3TVQAywMCoYxl3VlHPgMShW6rSixofwthKmvdHSoBoYKuHbQoFO0PyVr/
yZm2B1b17+WSPEhNaaQ/Cm2dngqi4PiVrfDpyn+PTdGAI6Cu/ygCn0UkTUXdYw9B
JuxrYvGFO9EkgvgLGv0DWcZRAmzM+tMkojNRUdAUBsCIDmg81nBrmbSP5b0JlFiA
/54mirRfIdlpGvsjdDCAO9LU9gTaw6MW9JfwgynJ22cUcgGsT69TCcJ3Bp/oTR3Q
gph7jehTaathoDIIrgMoJlqWgQAd/sP3Xxs3fDTwxyCnqH1BJMVbF2EBInEyA+jU
37ogINyEbt31htWDtGXW2T5CIkclTX6a3Mu+N/C3qZQDfynWXYvYVGvMH4Py4GP0
KPj+KTWxo/dxZKPvTu7MbwAwtouBJV3Gu7GpEzPoIHvvWeTNfZNUwe0ZCFZ9hoID
/OywWZXDiXxt8bnBW+Nrz7izV9TcCr8idoV8hNfHiYw9NhLCPwLvX/PMmA38TQD8
HwEhEaDvtCeuES/0gfJxFAUeOztdor6CIV5TNUf/y3LkDYLgL/ExX4qdojnAjHIP
z+FcSTfsQ+oEijyewZy2kSNX22VR9yvqOKdbpf4eQIbxuTB1e/YgienkhZNd9BeQ
rOuoM6G6IG+jnZ2VRxqqS8O+F6npwUQEChhZDKyJ1h0iuqCBR5X4RnBpJO8442VS
3VpnLbO8xzZm8RcwI0mjt/12bqi4VFTlP76RVjr7OvYEBwY17eOJqdzFFfKCntDT
De98YxapjWziDLZ2f8faySkmig4ruA+z9gFjT3BveYChmKe7wgkz0N9TFxJlnMEZ
3elvMoklNxBoSlcvR9dcrqrJE4KIl0vb6j66ynAm+XhHqcZr2OmIiTcseALEqt0s
Zg2SZQCUOhfM7XvexTsie8xnM5ibosENK6tUP+StD4LZR6PDAu5adnAN1aDS60BI
uUjlvkoRpSJAQ8dxbWFYoQk2CMSy8xD95mP7TEzOrMeTmq0CHbK4+luWs1hkJzLR
qL2wFIDOPJCIBRepFK24HxzGryStOuXa2f/JQi2MBv5XHg1vXLxo62WkVJS0QDX1
6jJN3EzqLo/uXnqAguGaGOB2aNJd0L05lh9dHADjSAf8vttXG4J7zF4xUaNe5N3k
makA4Tjq5m9Q1rgDAvfpJK2uwsbw6/+hqcP+3FTJkjzXXN6sl/QKhEvUOfYMLB1a
elD6orx7iVj/JxVCQD0+juo+b+Bq8a3Nxj3IiqYI/WVNTgc7n+nRuR3fo5gtluDZ
4RVMvbh3j6HiwYHDrSPaRKBguEjI7wWg2dVmp8gAINFxH2oKtHml7p4+G4SuZHhr
TB7Gzfwf+aMMnvyDhssOSth83ItpUoFPGX4Ri2iZSXItiFgU/nYR+gQDFGgLqQRs
IzO2E1wCzeOU9dngDSPtdXO55aKqyC0urjzOdagK01sTXhWFVbj9ZJO0eFPOUC17
rBaDnB9j1j7qtkBngaEZPPdtkB6CB2Ueok6+QA1SDPgqkW+HPAwz+lpItaBD82yM
RuCZW1m9NuGr4RawuA5qCODhVg56XJsvnCOx6e+DKTK5VkbV3dTFurVQPqxsR/bI
lVrMBQyCDjrEk7CDIVdh3gO0i3zAmC1irv1xrxuMEfM/ueF3qs3spKAXTvBAitKb
zBwkxUWLTP13nRlJQWHKJKO77JRzAtry612+PDauu8q/EYEJxO0GdCRPDk3VVuLj
0DmHvAbg7y9UuDysm5s8ixCDZpviFO2U1q6DCITcuw2na1opjVzhqDKfpksC3jMh
3nmrE8uJepZ6+Y6Cd2ex8QtigCQds51+SGSvZoSQtDD944E5sL7ubtCI/NFOUvYE
pXgeyg9LktBy/s826Jn6UKJ/iUCKRNqaoFsGB3YUO8qFPktgfkAR1zAVua1qNb4Y
u+yALGFBg9w97voSfOaK5dFprBgUdo08+hCLkMdWe2zfP/wToiE9TANQGN39Iebg
ka9q8E5xpzWGWbYPEpk6RiiZKmavRFKD/EwdIat1iZoJmojUAHjxuA+JCs6bho+/
cAAnxAw+y1j/H6WxTxIDRKz7/hSZoLhoxjXSOCpRDGfu1NjOj6gdgEb7gJiKFzog
FGIFmxsucWRt87kuHlZELgTf2/D2Nypp+jDm4LhpAON51rpndd64vc+Rq+xfGW+L
/ZiUaRrq3fQBbYx0bMT8pXXLgkuBo9XerYMfnhi0pwTYf/ArRMVFcjwdJQs/w3gr
ghUQEunhaW8dGnbCTvk0BJWjdceoN+n10EQrkbNrAuhN3n1HLrjQS4Nkmu5TBVhD
zeA0J7uGKwo95smi4bRo47w7MvtvayTnLuuhbtEgayWiqHwKyt3mHVySNoh5MP2+
REWnzEYzTcXyU83qU6ixY3aZr4xnOSjvlons4l3GqJaB/ow+woDGRDs1OKlWNJMx
QIscTe2JdwwV4aGXwlVaRYCrjT8M3cZVIA1dU8EicpuuRsE6w7pIIFqrFMOGWSIs
oOAd5ASdD4SQHG1FQoU1SDAJrWRz3IFzL0s1EHYmWiIC3/E94/Pl4dXGYiG//0hU
Bwubxokh3lRZDUjsnpEMQEl1RgHIbQPA9fqVXnCwc5q2+RPYLsK2GRl3I7IpYflA
uaw6bXMI06aRuSr0cr1Hhp2Q1TMODS6euoxXzfFSdErdfEmZsdFe1RWfvomE/6XZ
mQmDGwNzZRPUiteudL55ix9vT/UcU9OCGXlnBo+MvhgQXx5KMllLQESikJpUiMGq
jhUEVncMq+CoYtlKL0MdNT4Ok+/llteefYyBuHPWDspRatfMaQ4nJcTbyrvjjzzi
1+X4eFAYJca1Xgsa3kPICjefz9rJsZEdcW96Yo4Q6rraw/EIWJH1dNQkJKG/rwt+
vp/YTlvQZmVWxmxJJjAyMvNOe14pxBhccK8LIT7Y4DT4jf1JSVLK9C4xoJp0seiP
c1MmECF4fpKuA2CrdyyGVJv8ZgkAGYlFMy9FXuF38iccaSrXJP4QBWAOaQvkJ38j
p1UZXNRQ+t8bP2pLbRaBf7ygLeKO6HRKUBIrBUwxoBM+dQvh0H4/ehTiKez9kwQU
ESi9nwendUssL4jlkMpH0FqCNsKqYy0iEd8J5KigHjDUa3NOcI7dVQzLEIeoLuPz
y3LcazLdo6IlMm0tNudKMJ3gnERW22dTx381lXlPv2jS2gn85DgPljTb6l3YtpHV
vHxoof408VUpQEz/dvcrEj7P9BzXeVxEWfy5Pj+C2whaymsOnUEXeYpF0g6JpfUF
xGDRlVpnPfKYqsuW+/6xRCofDkjbZvSg5vPNcgQ9dx7DrLQ+QfJuB+rw+FUZhrfZ
XwQ52wU8GrDK9eAimecETLHs0E9BLp2Rj0ohuKTA1Eb430ss3pYj7YjtTS78E7NY
Z22J1DbCOyjNDJ8zUAtxUjNuWmP9CgUAfR6DQn2Fw/57XHo0efbrkWv84WqTonrc
sXXHulnkYF3EOEZQonaupNHrXYX6V2tBD4fcKhu/1hHuxa48Pj/RERBAOQiyJzOY
weTSXOOqTPxrocTYILptm2cIf6M9IwvWQW7xk9yLP9+CU0jrBrf17sIibG6isSSv
LrX7jK7uJ/5PBAGWODADwfhnD6igHW3h50+faN41Sykb5Sciyt1tnZK0vwKMtYKX
EtkK/FKy6SYHM4UasO/iHqWeJgJ90VYwFf9Iek45ZSFXYLpEjebyoMFYv9t6LWvk
9u9+Mc8f0lCmXCUgKghTyiZcIZ7qRtbkOtuExrHetNwHZMueOZJPkFgIi14EJQRo
pwVBdJaf4as9Eid2e0p7Bq4N70l73BQYSC2ijSEY8vEF6xd/hbz3wpWHMBF9yn2G
oTYfHIUTI9XNSPqAVAofa2rmfMCuabE0QjPLa6dKGg38zKaP0z66tb8YBeQOF1cc
3mDVMhZ5YENNEYwit2NE2bfp781tGKRIqnt2ajvwhmvmzVcjHzuJ23X+3d3Pp5M4
ldAIm24MtOVRbd9CrLQFPODvYdvJcQdE09nulST23uYF62iS2H47DqylL2fQic9A
OGQMutxOc91KG7GB2HRfzfCboEMRvhfO3VLCcYSG4RwQIBqglhp5gBhmNMmFzA9h
FWlNMwxeS2a6LMxIVKgsKzd8VUrWSFKeMzmtpgyEhzCYic10yU5jdjOdr9l7ikun
cMNSKkMw5nna7GzXDhlwCulXmzQ0bXc2OdGdB5n8hJbCaBCe6qnTDFospQq0o0yK
vn96TipyMhiA1lYKLBlPy9QZ1A+0eF2FJJCoSoiEp8GRlZtw6RX5yAFg3Tajz/ac
DEFykRd+eC+i8uYa5Hx6oHrf6ug1tG1Fx8Jul8Uz04/SfkEN1EtZeCGpqtXZtfcd
lwHv1Uvt82adG5UnOORLnDakjYENx1ZIFfvrD5hjSs/rC3sOpWCq5xQrNLeVx2f8
QnFeOA5H6RtDKR1lGtWVP5vKuTXe09EgxeV5Op2gsMX/fFwPkmvICXMsd8JsPOgC
3TMNSyQH+vpDFQnAQKaiHsLo44kuJlCwSa7smbI5O8DbGrmHsySz1+DloYV6P/1C
uXXAW9ZLTxN2NGrYxZ66IEP+lZuIkwDv50C/WMX2ogUb3QYNyFg1r4jBljBDT4rh
tNvjUBROpnJvXLl/HVtgbopQCIyMFtGkoMsB3m64QH2RH8uPhEfJBN90b/ZTnivz
uscObe0h/e4sqWVaWALdOEdlkBjfAXAdjBll8mTWDMgEsdeQPTwBeyJwk0obDw15
Pjjzz1BnE47iL155wIhv4Hq9d9Hp1ytggf/uiZA7IxG2WFnnpXFH8Hca+Kco09gC
np4UR/qQGLNbYEkgqjql6/l+lZovyM89KoLuVFsLCryDvzNTW0W/pO6PCSxaEpvy
aDXfCVMmSSylIGlKt8e0XpzWfW+1n+EFp3RReO/dvlzClR5EFSS86BJFdWldB9xV
59kbTZ9X5v682hXNJ+XNC5He7EpRXyM/md1W0X0Algkt3MtoCOwXnWyfUN6V8Zc9
CYnuV5V48BRkHhXVeqlwmRPZQ111ACb1Hyc4VgRaxZ3/AgGJjQxicsKzwgPhMjSJ
B7HFQ+wtN2c8W8O0QevgZD+mVeJszYA+cGSPbRBd3TLTOUzvWrBenLYNnNs5OrkN
ToI1K3KRiaKtcFXVQ+uJgcBdNQDI2M16L9LCX5/o8PBOP0rta3xpLnbKZHzZNSZC
3zPKhDpm8/sce/ndoWTLhysJ3fhsif7NdxcDDyWdcJp+cH3SvboCKxuUZJJ5YrST
SDZmCVi1H1BPANo/xV7WvYZypbxsqh0SFBZPO8rcwUDJkMJYaUKtMSNoLbtDHnoG
Ft3nv3KFQt3HEBqc+kQqC3J/kS5n/nf+KNy4v77dpyoUvWZJEglytjHg5Xi24Jvd
9bw949UGnogwQy0KfOYarwzJ97e1UwT1nVE1xOR9siJ7ATgOgj7/yOFrlkYnysFW
+Nj14+Te5Gs05yjUFoXhZ5FRVbIX9EgIeZn0E57MhuXoLJWz6rhQSvtlY5AN/yjq
biIVS3BbCy0d5kMCKCvJbIJdlI5oMvdAxkY6qoFigv88zUnD/Vntii0W4ZCO4f9P
kj6CJNsnI+BJOEla+gmIsAGOLww329hrT9PPVGngNPGdqe13RRe/OaKWtfj9+vuU
e+MEhA9CYYgdKkOr+f7taam29mesdUkLt+1I0wYlkHhIrvsTpxm6URBkNdGr2lPC
xOhJpOJXB3uisUb3eML6MQEtPLrGCbMyW7lNG/XKAFsQIVn3nnOE/Q8iIp3RttFU
+bODyVNrY8a0G1nwGKz68AB/A6iiA0Ha90KeQzWSiSfimya6+Ik6wky++svUJai4
aqO7FnlTbrIolvLf7YiZJd8EdyBFVSdMmgclUfeJdgt72vUnVv/SG82L3aj+oVqV
TBXh9kwoGxVB2HtRdA2QkCl72t5REeo1zdhGfIUyzde7nZI97Y0erMLMP5iA9LNc
AyOD2auT5xXPizgqybIH+G0Ex30mRno53Sm3RoZ0hZOz8vCDwqyuVCiFu4jI0HAP
XoXAhQvO3YZwSc6Ef1E/1Z4d5x2HIYL44N4shRTPwa2sr82YPya0EwR1RQo26hap
LGW1ujpqxffwjphl87fMmAsK4aTm/xqczooHoEuW7rqS38y0ilYFKL9Ulk1fPKc7
1mzxy5CGTOtMYnI8tM11VQ43xb8EGseJvnpuKDVf0igcdntMJ2vQsEb2aeSvJtDV
Jx8bzHeLkW+bb2Iy/1z9EPq36ihN/jUp7BTetqRyizpuTZMJujtlOS3NqAUIyk9S
2ISe999rpbiVnkrnt0h2O0+RItwJ9f5Gy+ajTACtzb09gqyhmw00GOn2u3k4rnFn
MlqeJs7B5LeqYjLnCeNjD2rVYZBWglajw6pkxBCHhNabtZReXvv27/NKb1c6MXxZ
lyUUIsJf12DdvYkNN5b/9qJHpEAB4Br5pQMEpKDx4YekQYqavNX36jDlhbQGc+GX
QKQ/HrPhYB71Uj7FBau6NqcaRcGPmoyWJ2WW0pcl4GKFyCMMbpeKXMh3KPwYhFYD
KRS+h4oWdOocEIGdAVON2zrmCx+1oVB0T/EldlzEhg/YSKVXTNpey0zfLVfqk83L
OPMc6bXaw5doGyTvEd75KiDhNw54ijkOmSBKvAXILFloCOXPQNjUNg4xOosfGguA
pvl5B9CczvzpgBVApfSsxrwmFKVX0oSF0U64Z+/GTBuEfjuV0rN6zwjfxU2hD1nD
r+V1R3lWQ7rrlXhKYDTDbeU7Vj18kbTDrzmSvfgf38MOo0BAoS3N80+c51ZJRIQY
3QWYvY63xUNaPbD858B5rbNLmRmbe8pIpZYOrggLk2wq1hDVL4Tf8nJH1IRA9oGW
mqLRxk3eDd393J8Hax/smdDtO/VQ0JWgDmNngCywyTaup7mGzeVtJbg4cC6T95Ya
ytZ7CY78RSSiUPdzXf7rtwCus/JWsFISs2ZUirDGyO31+guquDWrMCuqbV764O/B
fDBNewXonuCWME1COeuOpGqwk6zx+xXOeAyolk5LgSRcJB/cP/Hi/KLo16P5/u8U
a82SHuBuhlsiKwavsmCbyjhHIyQLbU1rTf/FnBIOTd2G5xz3mFLg7KzVLI+pLOc6
synMLwF0XrjoWfhYD1wDc9aBaO1b8ZuY2RxvpsCEYqtPPNhQy9yVAUGhbRLWEcpN
F2aALDMWSOti03ie0KNYzQfQRvBnBe1emU3upNgooTqc3opWI6Sg10LrmQXMg0ws
H/BLx5ucyok4Dkw/FEfLxASdd10JHlmdgylNN4WjBbr0oTJB+HJMyoytmE01+zVe
PxQ1OeOCRs9Fg3Y27NtXj+DfmFcnln5GkOR0dN+VkzhPZFE5osTmJx60nFU/h/4/
BPdqcaKowkn5fdDB85x5doFwNEKKvPv2vfQ4iQtBpZZyZ75HA2iuh9oqdlOFchnE
Mho/gI/6ZjH952e6Zr5HxJ7IJkyk7dzKi5D0+yf9v6tYXYcm9eZSHbVcn8wqFWDL
2sisEgmZzre4UyEkCX0wZ9+64/Zh4I5nLuCJ8HYppcf3FiD33Ic4eK/eIT6yZ7Rv
O4Ak3TArQxPn9PP8kz59KlrbCwfpJhhVu7L2RmO2oiLEO8GuvmJyfOhKn4O8Tb35
d/MVcBU7h5IZicxjwovpmqof9QVXjRGQMskyH4GaAmuSdPkNE4cyZPTZdcKSTGav
b4rRWHrgwn1ZnCD4VyyDKa3KtH+3jUItXhfbRyxJBdw+5DE2y/2NqCPKdrXNo4OL
HMJwtbRy+3DDJ/Gg25xx3ZQhsrCbc6owWJCRaqXj1FY6HCKQECoh5+OxaOJNeOvu
fQoaZokVohQggAI8W3GzzCgwkW8s01p5OxXuo3ISekXBojUO9u9WHXT312aM2Upl
zgAA/0Zo8Ra3aP2990rUJp7ZEyVMNz4iy/pXcLHlXwWfyb+oS4fY6LCzZV4c562V
PKhpDPL4i7scFZfQZAE1cdGGMy+DYY8X59wkne81C1p01PxT3yIkArI8k/Rmum34
d6vn31DIO6TfSAKaOE/WPrRkHeRdYkuXnqhA30kB3P+y6qIZ9TJsyvX0gtV5ajnA
zvgVUHS371ACeGXazZigQ4HGufsYgPeBXtiy0japEcjiSE8XTGmy4jzwtXMjaNf1
FwLQ+k5+gKG5Jrj573OLzyQF83U1O4GYKRlaZu6EGonvfe+YrfOMLdqUdLDP24Lf
mPzSFtStG1KgRthDbyK4mHriBMeRVbheKt+H30amGP8bNq4R+oFVJt/ELvHtC0bg
uB936eX1yIOM+0kcSkXUn0uBttrYVoSuwcnPZGeYQSknb8uz4bM6uGTN5WyKaMF0
kmJK8UbUlRYY0t/fSnPo1N9j1DjF5c1/zqySHwP5xEYBhUQL/DB3ntF1s+lBYury
8/ZQ7Sj0dQwJ/PF9LCgNd78bxuF9z9VgxMGMIOe8vjTz1MmEZkCu1F8r6zUGUnhz
c/w7t++pJhhtC+KhCjOwNa+1effF7Aww/lVeQV20WgVByjskD1hf81H68BrjEb7g
eF9u/aSApKI/BhgW85cF6wFgYytbT8QYBYVNOOvpFTbXRWzCckBBZKIbNVGbGbu7
Ymm+Y0ucwJV8jQGcgMr+aRbJJDFMo1YehkRCoVdBUHaBb9bkON4+zSX75vH+dUaH
+hh3iNOZu1yC3PgNCLl0ULpkP4ywwpCqn4XNTbCZHde0jfvEGMRv6Z1LqRuzQMf6
N6yHaGg38Z5CyJrrmuOPC7DDG6GN2vH9WtsVryeKoJzL+Onn4FYSubk/oiy5sKE2
/ZQG0B5c5kZCBto0XUdbM9ZHXGSQvf43PqPakrp0/9alzUddqbwVaZna4SThfBiY
iFjsI6zTbIJ4Dq7DCBvs92hWme1sXRXxD45Wx/HxgvZ4fWF+8fM467V++28g70BT
DVcf77idun1dwRzMdtoOjm6rMmEdR/ne77KfX+S7ktSJA4kwangq02Jzu26JXr2H
XVU1+yOP44Au/zyLXn7TlV1mPD/Lsvmi5ktjIAN1m13lBvCg++PgIFuQnpej3kVR
gjjh5r81hB02SAX37M6a/aJk5/Ub760jikZ+ygrSTCbbLcrVSxUzYuBWF0KSPYNq
cxJy/Sl6mT2zHzUzKuCh1nZip19q/lnMrvx306o4Nss8V5Lyumr3n2N8IMxWDWjA
K3SsgUFMfDdB284TLYQSRs0WWJMC5VSUFRs94igZtZs6nmMki/UI0tBp486cSQu7
CwMsr+fSHdfC58g/3+BgeQ2wPxNjXTc/xHEHXReJgk+hvvZXlIZXCdSp9f3t+zRK
rwU6YCdDYwy6cYyAWMGbL5WMR4Wvf86zdWb/r2lwvCsjjQ4YzfxHF7lISaCzfbYQ
j+MJ/QPs0PN48i42OVu5mrumGnt9PZ2aJt2wOgZHqVUIxSOObX6rSZn0aJj3oD7p
Zqk4440KjdZtNI+Uebx4g3eN+afasdjZWqOuQVuUBEQyxKwbN/sN9uFMHMJjVGYS
soYKpBOb2TX9k1yTcGtPhs33EVoLbneTMk3eFGDpyYMk1Jau5HORiPF0MzZskPEq
tTEkDElai+fx+sCo1Qptx/t2j3nq1ywPwe2/T/T6ZFdU+SoAvdhCXceDUv+SATM2
PhV9Gy9XUPzis1DQ9RiJGgSqq9nSPQ0rjxq4kPvZI0OXyjQXUdQNfGnbM/UFbb2Z
B9U2UPwnmGJnif44pP0z4bWQkz+6J/H2Yorcn8EBoE17B22KEhQynP8Hq18eVyk7
E9lQSmddY61EpRWYiklOSUUMQRi041iCBdT05XhJjF1EigET0a0FwMyAjVFodBOG
TNJTGV3sMxY4e4lMHDE/HePWBvsFeh0ipVjVWja/x8Qr2cpux8GdAWM7zuU/B3Hj
BT14hHAGRJtbAm4y5Tb4BK4sDVXCnEhvQMJssVuYettAyz2LBfAB/UIAXDP+D+lc
DE/r9vN5jXmI/t/W4E69GhZ/Qc6JoYn8YqYhv4nIyrIIP3r1nnSTpHloyZX2P25V
Ms+oq4GzBm7R7McoVeEiC/LplwS2s4NbJiyZzz0lZ4B6XAZTq+CPXMdfe63Tv6A5
JhQlgsJelyECd92bVvPAWtKhAfvyHyWDurwr3H/18shH0D1RlITVlWzuYV/D+c7Y
jHTjNh5DC8Isc7kMB7HThz9RSiqjSyTo1/rh3BRK6zBQKNWuD2FHCK1dIAtmQ2Hg
y9d7Cl/eSxtqtLI7rw/tysnyVtMi/elUzzt3cRV9WuLURLM50TDsL+aihVb39Xuy
ie9o/8q7QejVrblxb6nP1EO9hzUngtj4h+B35b3mABThXq46sMLorkyIcKhwYt9V
sueOmCBAEclWyI6j8kaUqRESmG9BS/fUyRK7i88BX+IE0nJVkuqoMSGeoBaiXjXo
lC7MjCg/tOI/0A3gC1AjBKjZeUnBGNVppRQbvUBEmgENaGjnrObofQpf6B6KPQoT
fnQNoG8z1cB/cQ4irwkSlW9i4ivkqqg0ZaXsyil/RmDY7URgrggdCkBxFooaK1ST
LZ92NK/wkBd8Qx2vNjzOZbFw1W9EdyaVggysM/Jzl8mXpgI/lmAiaoiVU4zbmds+
BxEnr1KgIZLDX1Bd7Y8GKfyBCKVsA1Gj8mZOqmuqiWsI0czuo6cr0kw0SQsLyHEw
cJunb3Ddnw74SCopv6/knaJReO0pxp0gSiTXzfo4mmbw8Bd3q1SWO4TJPBfxteLW
Ny4+POAv4HEscwCfM6Am9fPs8FeH1dgvc+oCz4bO0Y7KrTBaS6aZTtLPsF2J6hNl
LxWYC1Z/1r2hvsEIreDaZ89KHsz8SNTU8/XHPgssCcx/Q2fiSAgxOjqgCes9TSqM
dSmKUfhqjONpSnG5VxpmU++Dvrtpn/yP49Yyuel7q8w6dAScmSU4B7wC5dcMqtfi
NWSaoo82v8wK6ipJdZgy41AgjiGD1GUcWeUsbHYhDOVnFnukHiLMyfDMCfwu2+A/
ZRkeidfsQLFlugXDJI9gj2gmFMsZJAnfySFkgLPZkkocmvnmhX5kYZ2bRl746i3y
Bv2+piE6OWOGb7KvtqBkibk5zoat1ghd/DF1/QNfd9xnmIEstsFpembujwwGTjbo
nhVfEDxav7dpbXVK/GgHyZzt12SxX4x7MLtPurkAC+oKSJZydTuoyK2BmWGsDXaG
daKS1w2dBusUlOLZ6XtIIfAJx4my7F5CMtuBS5I+hG++yKAjW/Z9zfa3bZ7/Uzdo
CbwZMMsh/ZGqG54TXLEBe/MWeOsM/LfZUaeXldX7D6WGuA4bVw6D9sQax3qw6Pgg
UYpDUUbF56RmKMYOWWcTDTtWTTYMU6NdSMtDtIsrhK94j3FO7oRsPU1hRpQOSxW+
7P+51/51CXscR4r3zAGgv6MSbTdGtMgTamkgGRzanYvsL4sNJmBtwbtc7xNfPqRw
pnJcQlETnfIUTz1bCQBCKIrC7oT34xiYAO75grKCVA7ruekCtoNU24s6Uk9p/9O4
NCeTDxjiWdEMB6GqWDPK/UCLoCpplv5DnOexR52zVxCMCQyBQOv4UXanroc2uNeH
T8ha1tGLxjfU+qV1TGTcUwrj4fnLJkNrnkPHdAvlbABeEgWQCFQRhRLr4dHtyxzp
NtTmcksK6jrCuKPLnOuGoLy8w/w0ZzjpRdvitAg96vYJ0/fySvqlMhlQY3Ssrq2/
i3O2/4gJ9WFO47Yu14nT09raQzddE9vtabjFO5XY8RW61ebaDoabwexlXjbOHf7A
IVp6zsjMu3ly1FXYYycehN0z/2voeXT6ZnHJE8E1byamWBuWlpiIKKhdeQLd5fE+
fLXQnuc24X7IROPoxRxMv7pgZMdg6H3/5IeaHkR2bQMVuINRRvOwsTKHdcVPF7vw
vV01Fohxf0UiLCr6+C5wDYJMRc7cbqR2USxC56ur83EAXKwbKDqnz3YTzdBrP9ed
oVf9iIlWrgVs5Y0Vy+uEr8Xu4SgTyhjULcDNdM4+jLbSiNriUcmgcgTsnXZbHfbD
ajZzLUtPV8fDL9O+SOz0qa4DoL/VamnQKeBQmNi2XcaUwbcmn2VWb/72oSRlMUEp
E0H7WDgkVJRZAo+1SMiy0fAkljNmvIwvdc4LT621Nde5Qdqe70l9OPddLx9E5JW1
DjcMvFnqdbgDdqSE86yBFX1zTVRAq62b3rAa8FJTO5wHZ22wK9R3z4hNJrhVlt77
bubcDenFjUj4+82q33uM58yzZKo6F9quVeE3YFTnZ+Wuh071Ynzv4NBlJ3rQAHzQ
RfWsNlNpMWfcTmRiGza7eFxz3Id8AMknkqA+4Y0tOJ+GYcOJKuqhuel9W0HnAPtt
+l4fqQgyuK1rBOLSKSX1HA29mlA2zKGA/ZAnn+a0Bikuv1GKqw+/sbM5JgtLGwVr
LrQFv+2/Jtsgk74kW1TYIwMk4xB92mBaVSAfuqenVf17BGQ/jfZ+4oSW1E8czzlk
eQHmrz07tmwC3+BdelExhd0YYBLWCyq57gdlRqVLxkTu1pGCWHUvj8Mzb+bkJMzk
OgUn3kG38z3MnLdSSc/wsHTSIPn4Olevhk4QZggENwx/T1O7o98X4MHPlBoy+igL
xZhvfgJcaX5ljTfLC6QL6Wt1HeNuD8oFQvaFzzPe8slWJ9knEBAay+/IPrZpcXcE
LWCHgxEFinnuWOeKUHpGP3JZ2RcifvidepI6EhYBcYIyzfGXXlhf/uUqlH0uhYJA
XS1TdvDPDKqZwqxN/iDIKTtM/uip13NPXs2MPGNqx8qG5eO3u5d692UFfz3+ffSp
DJpdd8al9+1vh9amFpmpAtBfzxDNonIMl8zKmcUdmpzGlMfIbO2uylwI+ruXPOFK
1mECdD7kzs/nLIuw5Bn9TeW63CLWGam4PW017MgePnAt2GoScvKCwREkYxYyrvuY
XpU4VPMpgJlmrkS/meqBgj6chJUEGHGQCB9o2wT79SKbjww1sEk9xNgg+HkfRdL2
rGFxP4d76Rahz29cFRmktQ0m82eFm9rOeb/Ofoyh31HwUYnF+NQqxcOanGU4jal6
Ct5R2T4qMROFEhbYPRxxk9PVXoBh5/C6w8RyT92+GO65dypQCw1ndIUzfe1hptin
jihkgEC7hvbAlT2lccZ2wu5Dn5yY8O1dqFvB8tR7s2ny9HAmFL1qb9wWZTlm+yKX
XvQ8nA77tO8VM/B0ibbL1zfRXgi/43EXaprd+XTsKKOoWoikZCYSMOGGP4myF54w
aiLvsFR4nTHTzK+5JQB1v2Qfx9Uy3SDYVUx16qCjaAAwGLb0VZO5v38/JzO5FqAf
mDpXBrcWCwm8tDRhqfbW4pL0z34D/8c+iHHxXYfI19AP1oZGevughYJn+IUHski4
G7Iyc+ASh/SN7DsXYjf7mYvzfmLAZhzJaRbyHSCrO4foOnr/SVadNbmxwC9K5wwf
cT0noBinGcbf6Cv2CxgmUrAg5sEXDXDH5SvD5kJjRiMkWR0y4bPwM7YaQOoDhdtI
umAeJ2aAyWC/k+qYRLLlqlSQtZGridyoapaPI3MNamXfGSgX92rmkJEeLCcxBK/O
uOknj9P3idYvscWnrEjzAF578O8UdSaAmnON9t5KeB4y/uWnVWCXKa+YA5DRUxOY
DI4BpDF/yV21r29rviNT/akmmaYZNsnyHOh5Bt4oCxH6oeyijtX1zcT1tky/Vuql
esnEgauMQXsxy2vfvytM6ZFKuAEkeCp6OndOFOEaGn1v0TL8HhvhRNa/TA7cso6U
ifdDN4C2f7L6U6RfgZ2COGDpiGblaV3/FoaBrG70eciq8KhpnevycxKPLUeZ3uJN
gwmG9vd0yuKjZ/UJoAr6S3mFyW00EAg9D2/NaPoiqhku3wVUNFrOuf4/TDf8SXz/
UmhqauFZw+CbbeRUvZQ8LBxUESNTsrXR0GaHJ8HAzsIGguTWZjnnqzJKHUfjZush
vJzZ+AUtcLhFy3EvYWFcTsz4XZVIfR1Dkn29zahdOD/iEJZOipA9OnvANzhf5iJl
6rdYVrW0nlzFZHGhihB+PuLSbEFu5OjxLUTVaZ8aCyevzt2iiflFqh98VCPNKfYl
iNIMRlrrprOP74nr37OvmqnzWRoxr02XuQNazq27TWCSjrcVjIuUhnqOf5PDzq/4
SjsVsrQ1j2f3VKw9Krry6H4zKggG55hws27MA4+2pN2b6Zhe4OcRrxNGh6uuOHph
MdgG9B/241WCq4i4ftTfnv0a/r3KwxNzUO1+ZoDbNToM/wPSTQZQE+87K/i5K580
JQvB42w2UImR0sV2+bbuaKpEtHfxK3A5VFPU191e3AT/YkkvgZSmqx/mZtbuqeSj
lkLOFpujtC7vBPnUmLpfm3jv68NjZeeC50jHNk7E0e6fqWL9EsGuekxo/7+JvT9i
l6eIHxoZBLJztWaTLDkBv0HcSZOzxxfgAFryD5podFmrn8DAl1mmnTdy6oPCeeqv
c5YXmBuJ+96CS8gGdiPYfXmFfn7OE3+3MHvJxmndCgZCY0Rrzk5ZDtoGxok2rbZy
QWLMempq2n7V37To7+uJxMc3/+8pQhmACMM1k/h1hQtPIf936dBeBTxPaZ2SEvia
kVpkeeKqqRRt0goTp0kKUswFTNbt5KWL4EDhzOD5EB7gcvQbZYY/8nBs5syXBP/I
HhdiM+EwbUhY7AhsZpWmqRPx4NI99f0Q+tRUGHvsLjvBRImqsu0t98/YTFu/fixU
J3XegLXEirMLp81jFBsQTqrz98h/ASxjCyDmhVZSKq5HIH7HI5ATO91p6z3Mjz6R
aBaXkoCWx7XMjcxIK9M1NoFwD1bJuQGh79y8qixqa30g9sT7s2ldrK2JiR79t7ag
ORVvbaj4QsHL1P8eqJVk2RN/FlYmRTBy7S2psifox5zaBMPFVrGvpNGPczuPq+QC
GjwRHmhV/f1L2+LPRwX28tKtfkcb899A6lLeOogw9OH0qDzTN7tDAU21YSWKnXoF
n+c9kaHpy8wsHplU2KNMRFHad1RIJEfK2FxI/u4TS6naQ+SZ1QoYT1CeRddoKLSO
8KDM1ICO0GLe6Tw0ageFdpRXYAW67qWciTpCi6ks6kGK1fOAHGzLLVEQ6qID9z6Q
rWYKhcBzngXOpV0IfZcc2zKGYWJcBsFKHCpit/Tk9TR3DCssZzFF21SI6LCZEIBV
E0qoVS4RG0jAoF0wECgw1ZFfE0ilqrpoRDrbSxrubO3rO6EV+dP3uy8ylza33Oqc
X4Nu/u/Xe7aSN42aeMCW/Lib4d86QaJpOa3fCr/V+HW6rI3v31X/OiZW4LZOosE6
323oxmSurKQtpklOgRxu6j7aB7lRQIE9Sd+kgjkbrE5Da/p+yR6vN4A+S8PlcvHH
ngQhsh/4cAculzANjNc5WhPwFR3uBHIJzwpuzaJ1A7Zzk6h3ViqfUYt/ic9h6ZMg
TliDMYl6fHMDbGfLFj6GerdI6bcgkGGhFgl+ExSboCaRItENIdvHrDHdyZdO0uOW
sSgecbBG5xf3wFDLCrkl1ltEhohZEAHNFmXEluwUBP2gnOHab1MUtHT8S9fptyvL
tgbWuweTMOyKWxUyWxV2PJxh3QnR/kYZjzSg4IxGct4hsrfzNO96CA7tiT1einhZ
HwUV+en4O8DNvwSqi0V78hGac7OgchaTfDn/r7t6JDURWBkp3hAjXQhWVpurt89d
wtFTvQ2SSVE517HOku5HNOYm5NEXVRyr4zJnvsPgvhyLVPsBAoEeCmrlyrEJmDDF
dj452lGgFXrwxfimNYBVaVgjqlRqAvbHRAIE3nN4pR/bS10InLQAknAfzVvRN1FQ
TPXxoe+NUV6vZ0nlgS59RsepRYiDKQvQqJdNAjRFuTddWvHyfs0dKvyxpH2V4Nw1
1d2kYD0UnqvSFfHm1YWPL4JivoKV8LQITJTDpDeekSZZulBo/elupWRR81Bu7OE5
Yrh+b6gG3FHsLQYXbfOlBZQ1Gef6VTIC8Dsl91CbejWVCqiiXYTwckv2BaGm29Hh
jZphbL92HBqhY9YGuS7WBV0vwj+Nu6oOCHdvdrRnJMXJrneZF4LX9v9habHa+amR
RnVrw6N9e2nAh24ZXL1kGpp+uoAjV+TCwuFmDVbhCYos+BYc7AGcVgoCV18svjfx
HSyT6mw73JUfp7TiRbDBD7vo3GhiSxXSEVsj/u3c14PmCoKwo8gYpetSDTGwLllB
GEhulxnt9V+183gax6M7MI6vQCEQym1Fa6bzxOGxUylNoz48kYHJv2HfNXF+BdIf
x//LmYU4pGSDf1X1oFOovOScvEoW3ZN+IjgIuxihXobCGF7+Rn5DNZY1SNGEXcHe
ZEcyp/76YqjqNkmU6N087lTS0TkYQIQO01YP6u+RlQQdj0SajWUCRxJY3o8pZKKp
JmvkVQGBvEoOYMHTQtsgHEQsldtqFzfmIstbcRN7IHSYZGqeEfyEO6IP/jRtiUNp
Gmp6uwAN4VJsGR1kjq6uOdwEVPS0SeuVlMtKezGnDaww9Vms/wruypefLiCJHPlk
ydIh8qk0K1JYWmrqauT3TY+934KzeqzGckH7vgbrKO7GaxZwiIFh16Hq2G2J3hIQ
HFTe40m3xCpX5uO5hnFtvwi5BSXqOu9hl7y1lOMhn/Uuk9K5OlVa+E00NMSGWMgv
iWFRqSt/ZWJ7/1JDPG0+wr1dRTdW+tCRH6h5ng97VmtwJsX6N/0D6bFF6G0T/+lL
fbXaopOVIgpzzpzC8IvRb3uZC3hG2WTecY9GMBGZeomH/zwMQZ/iQUKrUwNHwNzP
JakS8or0F8JMt3MQQdY+UaEavCp5pshaLtg/a3FsTC54vk7eeP2IBQFFbrKeVunz
DNbl4y4hzr8qYlCwZm/TpxA42u5BluVwT1jKiR/IMH83KfPi2hj6wLmB6o401Dv4
oAA6FEXAbh5B4tVfrv+fyBKG6WJnm+9h5cckuhE6b71te27WPOVLyOKDu6YHIL+h
ZxhLozyVWDX1CiDi13l79htaLg2OtZIVweakXSZcFJDv6xCMzHoEwxn476v0M/SC
jUU3zxV2U8vJwQfeUPqNgitVztJF0SgetgLJha1chIq2smKBIxiYjQQZaXF14FLU
kWMQnRo3A8VkNNv59rExpmTCclm957GnUEaQs+GOkx70O3LiZnbsvIuY45kUH/nU
lylBVJB79QSSr+zSJ41TlgAgGL9Skp05VGDhyADzETD8j7h2IhXI46vHqTXGT1YB
JfHtBVq83jCAKBaUUqOgq8lnCAAwGYVh9bkz0yq6ytKBIhe93b/DJJYo0bp703+E
3FC+swyOXFNsMTH9VoIE2ysETF6KqmivlpxNSkuK7hM1bwgvAAz4M638JP7u5Muh
NX4MljALDALHvWX5WiA3sc9z47afLNDvd5k2IcdLJ/dIzw2Ig0MDpM9EJXDLvLxJ
wAifa7oMsw73mdvYbFxb7PoPFVWQ1gZXjQCEijbFqLcqC6UM8unAZB05ocjJfuqN
L4RDDmOaRu7NSW1nP4X7u3dObfp8gMHlHuRXrOdMy1Z4cges8CddeWFc+r+q2yg+
7AmEyhmKEVrLEDyQHc08Yyhhk21KUSi5dSLkeOVPGwpzk9JAZE2EBPaFH1mzKMff
OsdOR+EOxvIOL9mYXnTBd52tJ3HbtBsxvrHvs7eKMZrZ0pr678OZENNaCLqfl31V
+teMswZhMdjF95pA2tWdcG9AUdojoWorfDIu8PBBNUbh5jmYvj/Eliaqx6KF2RWo
zilo6iBSbgnXzzf8TdwNBaPcx12GGQeXlYGyMaTLgVkiLvr8WKHnnKzeJdjvkvuV
UF/bevw+XwkWPS2BinuwYS15bOb9cmsZoOOqghCx02NiyKitqPEWIViiDqw5pi7e
XVrARapPTu0m5W5cutkt06OCuPlKTlGCbeZy6N3IgQ8E4DdNy08cObqltNUZEkta
aSZ9gEZEhQSq5eH3D6H8Ryo/RSd+bss6CycmjU3nt5/q1wzCgsHfUL8IVy78NHOG
mrt8zbHtZ21KVgaQKQBhV+CkJPUJ5MTDqGZ0Pu/Mqm7rHiJLrcZVZERn0utiBRQ4
Z9agi8n04AE1GDb/MZhXrtrsTtHxgrHHeFGw6RQyUSKC8hbXspc48QPK7ELEytO6
3grsV1GGnTWkdV3Kz3AnHySy6ULfP7V59BdnbuGI63JF5iXbiJvB6wnVj4p2zYri
uh5XqmtRPKjBpsYX+a0yx0/Qsr7gxWsFlgv+4+cOmSQw8BF9s2gOQowaJMXnS4U6
8LPLZ6+uaKtKo++t6CZkpE7F+tREhthGYCB5PJWlFoKTFf5fVqlfjZLzYmb+wvNq
VQAqVx2QbAT7+LhXRjAYqno1mzlbPbhX1+ixgN9V4X09Yp5y9pzhzIL+MexdYDSS
ha3pD8/3kcfq2rOGih8FrEEGY/FkWU2Efl0gUk6jHZB8oeiYd6ruuAjtnpje5vqG
Iq27vQjqAs9uzHVaiyqTinAh/CN0OjCHFQCf0Ru5eTIyfFPXSrf6uzE5ztyDV/A/
KPqd0PL5ptqhqiL6Qj+bpkWki+++qqyEjLeKUxgabVwIIEfFSa17V9anEtP8xvSo
Hqgw+IEA9be2nNHtbdG57D+6HgZQwFIOVpb22gDzlDmDagfL8/uHOMmKrrzmbKS1
3ua6m0nF2EXE+XlYD5hOEKe8PrbFA/r6J1AOkrNjhwlMEgMsIl1+E3ivwhy49RPY
uIfptp8SwOMbNPl24u3wV4Kv9+K3RqeeEf/d78QQD49vcXDxuWhfWDrGckAhbjtU
eWpsfO5Ve2KsloJnv2JMqIzYTQ/WSnlCSZ8WEtIYR/Sd2c7mOqCXVRZZg8HmULZZ
yzpCzteOSR11GgXztnnF4f9VxNz22MdkMsXgMF6xTB8/cKZzDQVZKp7Qqp9wbvkA
9cmubcN8VbqPTpxmzKap/JKRt87/UAASvU+fVjvodfZL3ybDeFcuAQ43eBA7C7pG
WX7l975Uxm8+tWyQ2rPLHF9myjjlRDrSnqaFVyPbY1GVzGIFHK4r12/vm4dtSYCL
Mbvhdot4XjAZPam4j3bF5HNJCi42pQt6SYU07Druq9583Cz9U5LbL1z5pFewFpAL
3xYuW8WVb7QJb4ZN1tjYNwyjyq6C/G5ccj//9UUdUGriaxbC13hAA5GB+5uczfjo
tD6iGvzt2yRAzNllFvSBXXbIFgIn1E8SgCP7jcB6RIt3FibTnHHRYVfun/ZfQesK
JN2z8VA3YRJTDwkVZZT1qGLG1onxGGhJ06oAbWLP55sovCW4TgPepjw4h48cU6mO
hxilrQ1SJaVatLoa22z842ejmN1AqLW+463HJ79tu9tfN8IuP4FaLRP9Et6Ygpo3
s3a4ug9mC29hK9MXfiLRlZckJtz4U7LxNPccPKic/2gd6aeUQ9i0MLq9tHMWu3LN
v44O5lTVEeEJGDBzGMzE2hoXmElU3QAYvcam2H0sP23ftm3WmVy0OYAXD11GqpJo
921IyQkE3Vw7Ia2Mn/KWfef6ae8DlytViqjhJrVm4s3wShTa+8h6i0l5XvKiZU1Q
9eewOLw5YLnNBq/syr8QthH/iYiEisDNbA91VIAercdu9fRYJphJ31ioRgS9el5B
cVh3W7hSDZrr0a1zTo6RtLRURhTBKf4RI8M2FM0N8jJBMwGt1eetDu5CpzkntDTd
EGvJPiDn6b4LFlEXoBoM7r+zOVTK+F3UMFzBUGiOCi3YD7F1QV2TrvWYdY5M1X8o
fdWNf4sRuC2soROsqcP33w27taV3ePKPpOoGNZ7yyplzKmatIHtV1qNaXuRWNL8v
SC/6x+sNtuJxd31YkxgOcqh2/glRWx3+NFS49r3Skgov9gyKulSmbGQdk/LB47Hq
aI+9vrSMV6cA0p3xI6DypFhHMdNxHXBEIOH8VPUD+gFaGBSZDNJOXWYZoEYL17vb
xDDWzQyhcIRhB2mJbN0atMxFm8k+dOVKvBAFs6AZE1lTilXNZW76Dwb7Nxxl3AfK
58iOPgLaJHFN/U8rMBYLxI0NbKvLstUqtzAdk1q/CgSNoLUW8xrBffMaQ62rUc2W
USuL5g10EcPLnX8NzFs/mPvDq0qnUjz6qX0VyTnT9hcmQ7WrzYtrqkCDMARotPCB
pVesGFjMt3lXjvbuZ5U/66GkpgCE/pExcPmFdlrfEjA+pL7Km60UvEjJNFTIzfc/
FsPW3tVX1wgeH1bAANBitJpCf7B/au/GU31O0PrDxDyfFfAjKgrgM1tMNvZGCbkZ
lx0ayCGCtRSHKk6VOTP9d97nmzyCnMuetlqv492hLsLieKUOIIxLk7rusM6J+fOx
DiBnnezP9D1U2tQEwj3g90D/eQSR3owaNv1T6p/aLfy563J268NU7EEA81yjfywu
l2xXhg8eXinAAn9cPkKrOaNk3HIVAQEneG7uD7jkAJa2pRqwxKucSaprxGdb0mDJ
ONO28VAmvUTtofdYvBV46lOBWNDKDfnPvncm0PpaXfgynZ/2J3Xfa9sB95NdLMnb
dHmcwMebaytbRv6/34unZfP8R0WCu+8/xmlcHF4I8/B2sGFCMnLvowzkK7DnHi3s
5TxuL0hIurajS+uhdjvCA/NoJRZvY+EkFut1zqiZ5lZ7vB9v1qqGDejaTapkFQWD
B3WCrldzAdy2YUGYI3rDA33u2L+TrjZX6OR3yU+ROGwoaCGulF6mWP9qabMJWU3t
wWCQ4jhdhPAEjgIfU7mHbXrk/y01tVFYFIB9aHS3dyU3iKc7OipU2UwlIF6bP0In
/roxenQ6hVLgUchWTwx+WAZ9nqPOtStiQSD5YchCerOwJMykQgGTqsisTr/zqoFq
Gg5y5JlxZWRje2SGmdip/d0eGaxUYkuDl8U877Q6RUV05gxMSsY0HfxGlON1kLP/
JsPkI+HUfMKLvlHDJElkXoLcu2+qm3km+1XGcaWyqYGOUiaM+IzBgVbjkvxr7lGx
45SncMGcSGZDdlSiqOGNPvdCjLicsQlUKwrSVkBB7NMeO8EqIclBdnYjw/LREJeX
RpUUIbaks103usuXxbnaztIqDHEGXR5W98E36xYnw9cDISSX71FIOj+oBMD+H9bx
t1wCoXcjgDqSrc2jYB9HrHcrLeFWMa/H4ot5BDYUSFa7DXPxbGkt+mLai8zcsKa5
auid/KA9IIag0IqlXkGYcIaiSWEKhuBpMY0ed5JecQg0eg8IeJS00DdCZyvjhnSx
Fi6+KDS77PthvknjOkm7s7CFHm5j4y7v9JyUMaGJYOOclhVALjIZE/WX6Wg+IZ/x
Iq9pVSAGVrDr+Y/831bWTxhnHg0ZHViAdJ09p8OXip1cPTqC6IK6C6+8tyckcfWQ
rZ/fpTOAdjUX4jKUtEhq/9QiFAAiAqLCcmsUs5UqmKCjfI7T/VhvoTuYZmsfOhzO
1fSWF+d3y+ojxZDBhRPBfzFIWo+oWc86R6LuVG7EF9lPqC52Iwkleg0Ohe5ZWNC3
9RitSv9u+nxBDdnfvDn6hR0s9MgKCZzVRZsVmFk/1Qe70wSEylYZr2/wbn4Tgvoo
kQeBrPZs15G4IW5ifLJ9d4xIxPhXX2f2Mg7ZO2x6b43ds8vqtp7B/8m34lZLKyvW
B9DlL0K3cMnkNX/rSJ/Qhrf+fmcCPSGDYzXJT3/HXCCGZIA9MFE27z2OEh2WxxEi
l/5oqsgyLK5gUjDsKYw6/jGxRcUniJqfnhm1F4j1CW2UWiwQXTFspurJsqbSWQ3p
5/aD/pG3auUgASMmYM/Lx9COhCgIxh9WgFAHOh1HrjwI5nz0yoMA2tRq7BrMcggD
jTvMOsiwRbahT1AiywkyCj1e7QJBiDS2XeIX1ElNRRoIhSH3S94rPy630TtYoN4U
Z3L8SjlcGTV1WS7Ygez8uJPGV222FkeLlyNdwYb6xgckj+N6/wDZxityE/r5Qm3B
C8E0bprimeh7ieD8xHB6LPEfpaY5RhsM/Lx+HpkK4smZXUfJ0Bd5E1GqEBza53nB
YW27NsHrUkzxtbGZV3/cNfNhpcmgCy8OKhU+19uWacNwa5kuB+BH5mPmz5B0rp0I
J3eSqH2MgMb4vFzOL2glMHQhtkli6r4ORwBW1c4NN8Eb8LZlCRBn33AgjAmo8yUQ
tfkABaf1ghTLUbdnbwPc2mBmo0O+6a4UThl8xLscD4jiDYZBtr3azuC1WnWilSjy
3J6vaYLhmixOljCXOodQYJfViCvr2KRd59YWifLsMWtwWZmIAJIz/BivYTdXoBu/
guG6rBBEYbn4VDi8DxmIzp4YS1MrItf1ufFO556IzX5vFklbbY/JFAhILq/Hm6bo
V36q8OkOR90tPuOY2RJfLOcUDkYB6tXSkbV7N8oKvp3Pz5s0BIcCtp6jEO9gFzcz
3oNoG9jIprKU//mV39e4aTJHiSdGo6gk0q6MaAbdHtTO1f8s10bdq01AbZh1RguX
klr9ZjEar2b6LbrpdbnVissTaRJcg40xhKSwTL+Y+8pue3RbJ+o5wyp+vrfcjTQw
SlogJzMHdEQaKxZGxVaUvryV3/uGsINZRexGhlYLeH1xz7E1R18plUV06lJak1DM
8xNVHSob4SzZ45FMc53LUdlPrxH6pLHYJGbeaWaXCN6UhXVEdG7v0eXiYCcwcbOV
Z0a0ww5wNhjnZ/+76XbcFzr4Y3EHa6GwmOEhqRuGdHHeCmRrh6wkMSkRK1Zm/6rc
pKHk1eH1T8eyZrY+esGyyXoItCFgdBU9c5e4MpzFP9KnZzB8+ZVKey7CsnxGNTDR
rhu5iq3cPnsNW3Y7dwVviX+HDIiLx2jKz1oA4A0NOCuSqjZtGQc5pqHpxZVHGrC2
wAOIedPxwsUDJ0QhVyZRzNONkogfnru3yE3OBw9SC926sx4aAt3jBLMq3NBIeSOz
xlhPLaVkkVGWoLClMobNcgIH7hWBMgApbstmaraCbWdjvGoTLZDrxA0Zv5equyP3
DgKntoiPC2rDSHMLKgGn25OV8kNn/zzDHscNrtougqaiYJLvVFjwAAt62H708MdF
ORKp0kEt+BtVMvUh0l/Icj2OwMlEUWWROEQYyrPE1cgrLm9RW3n+nmw/CZfnlo2j
S6a4olmmaR+rT5PLWqyx9VPkTnVOqQfrGh8K3pspbKEP9iw1QmbkiLwTQfGhHX/H
BeHXsw6oHPxLXo0cGX7+mbWwZJefSHnobE0JsP+ZuVUfYm7CVxlY8wKDmfxFzdmB
tS5UikDkqnZiL8gCZpgZ8bwYT86M2hIcIId/dAmPbjgWW7UXu9NEGYdSf6S4cTwF
6yBLNbRsdWjXqOT9AsTFSm3YfIOtSEXtZqIbworGW5TaIMguEjIhiCYRFE4ABFSH
0PrVu+388ROew3NADl7+fWItrUtxat38oAAdCfNo4LjOfpkowFFPrhT0qQO7bDri
xdjPiDBJWVUVUdoY2lmGIhCVmV7Wnfp+7kr03LrslB1miWqD6fBKIkmhA9yC8sJQ
FPX+L+DmjKZvUkLJMB5xYoKIIlXtDvYLxiZjXxCEed5+T4WIvgkCyAMnO7ICdgaO
RW8jAmevJbgh3fbL1cMTpCVXcc2vrAQjjysJ6KVZB0eJJTLxLcsu1xOVrEHNQe/h
Q6S9HoMMY75qKZMzvgSvhpwdAqEwaObHC/+OssbVruAZGtIRHFyBtK3U+MzN6FDd
q17hYnyZAo76HRngWobkRFQFqmYuAVcZVsPh++cp/Me+XDgd7I6TjNXzScqXEmRJ
uzMcNFaRObO4c8fJJatoeYftGpp5voaADtOUacXIO3o9Vlkqt9ekBmKtxIUL+VxH
7bJEHJlHRcYovyTJrBi8u8aT8+3qBodfyKB0iNqMXVCGQK9e1TGtblSi1t6ckoPG
jag6k5PRN0bSlGmQoiXo63TrdkQm+8LUMOTcx1ml1wE6vvcbAnwoPLRpkM4wlAMS
mzVeUP2+FlDkeTEl9tD2WnBizBT6CgenMgQ+eDdjq9EDCM7SAGzlkkXpa8IGMcGO
xbXQyjfIWbPpc9S7EBh33hjT5vdmGTGc7FevYsaXdCX1zkfNPdF/VBqHbkYOlknw
5+7yHpP4f7l3TBRAx6adMZCUxDn6RsWzs9bd2ksun7kbwCPQAOhYKiOHpbjFSAmq
Y2ZyaJWV4QYAKBq98vLMSDbYD8ewdH+hsnXfrCzYC7zvA7/11LenCW/IpdK8jOw8
4xSHtCuJU8Scu4wdkwRGTD0W6dl6+ovtQzeNObc6WawuKhTQusgDl9NHWF2D8oYi
+eX13G+A798Sk0OQViTqBUHxLF/UWl4SX9Esj++EkYB390wzp2U/Zv1ItSgxidSI
UZ6wkwm5jsb7qpxKcNWQOE+gE3TPbVnDN/8vBetWDHIMnQbkcq5mojFBfxgZu7OK
YNtgs/xByVK58sJhsKst5xQFnNWNipkd1F42XO1rm4kb59I0XD4nuDZiWGbQgIyp
OMdc/UKtcLueUo4W9BmGLWGqWBBD3zz94HmxLN9AXXcH/yWsI/CPAm+EuIsLrfg0
jUjRoqPT734Wl4QSYoah47XjrhpdOqI5PExgC36Z0gCfzNZ3K+vSlx9AJu9rLZ5c
P6NPHDSamYViSTXbJ86L96XM5d+4BWXYrcmravdIxU1IVTxWMOTZooYukRu0ueGN
/XoHNuvz2Y46AzH3ifkkc2td1IXZ+hEbr8oBKQC5uYSr/OyKs6ED+DM8uEOBMa8/
p+pOV1xlz0NutVMLOhVk2hPBHPwDNAHEM0OyH/B8gbpmkoU6WlzpVEEQj2UAHywQ
bZa4yX0FIb5qD0HbZLw8PBgk0uFFuMLZrG7iQ8dyig4j2BpTbwdzkFZAYgMBXDAb
wBNpTnnSTCuQTOFOATSoFLjDAW1OtEYrfJak0hjmbvgnq3K+pXA8hSZkiMXzkEwl
QQLm2FOKTGTtHSkFgKfdHeaSdpNaiY4C9GJRJbsX/gic/3vwhnwzj1IscS6u1kuK
e8aLkGNuZiqeyUjOdRQhCr3wSWU75YaZ31G9tHpAofMzUWAYjJB0+/Kmft2wdGvj
5M6xX/9JlXBBUE2CPfxPh5rrSiRNx2mWyZQORwTJjz0A1kEX1LgVPQx5p0bVlz6r
5YdlX6IfTjs+gRR5t+2hJlVK9sgByjXQj7JbVrMyfOdJ+zNOJ4GnH3L2pWUUAtVP
AbOJ9mgSP41/sQxuKUoFK7nOFUflG2VyndvzJpZoP7UGD18S0a1v9HCSdnWOD+hc
vWiNy5hm3kZbDPpQaziWEekQjhTJ1v+Zw54cRVQu5x81kUatk8pOZTvr/Lisz+Ek
xcyllMo2pt3ki8vHB/RfzgB2BhueroSpcoD1nXaaGR9+YTYy3Ie9+SsAkRJMn2Fg
UDKzZPsyswJ1s24v46TLLCsj0LSOMWFBThA2yzjPhcseiziYeelCh4uyn/cLKVcp
2jZQ51li/wSv7BfBos1Nf9i+7+c92jgHUmc7wWM9Ibzw7TmRRTCsdEWz0PipWhfh
g/nDR6ZtSOV9Vwiu98Wo7yOzYwW9Oeh2xUqkrKQE6BNIzf/jNTn9+3e1G9wdHmm8
XM781L+7oNcvKT+/HtyZQEdzFpX1ZzYRG9qCpU9Yve7tBb1qJM3iZhMRInyPx3mZ
rXaRX0QVfDNXfCHuuqUN02pMDmfeMRK+RayZfsaZop1Vx8G9pboPsXKpy3wnYgmw
qXKjb1y8R5X4rsypyVekl2AlOtNRPe2xi5OEcMdpj8XXbo4RWM6a+zWRqIeqsF5X
Y2RNQkaZXxMoqMOPbFsBzswpPz0Pn3gFc1KZEtmJO6ZGaQifLjTVT9nqRTU8Xqnl
hEI3JDdmjRdQBDheonDwRVVgpVHS3ea6IpJ9TSqWnOeeA4jUdEpBfll1AvpJNAp0
BRlNSN/RWj/EpjyQKvQdfbnZGQS9xM+OFtYfQJz8Iy7Bgc+p+QY2HMBx2icYBMiH
IEFjyqahioU6kjt7rjJ4wFHgJUFBbvOoTlg+q5zAYff+0JFp21PuuFwsQlbSGQ4/
ROIez+PoKvHI3rs4GCqXikp88i/YZDvgeyQ/lnn4rALmbXEwTKYYRyn+PwxfBbnz
QndM/keHrNWAWe8V/Va3lp4lM36Xy2fnzSB91da8gS6W7yS8WvzO3b+vatShdDVd
zjEXEG2esOZ/4dz0dEJTQUypSXp79e23vT4qE+hc983SmYIXxUU27GIpZ+AsF7S/
MKe8ZZVCQWZZxlQuaCQaz6JxX3qcBFbQ7Gr/8dGuvKrnqQUaIod7+Pb3pT5qWjIP
sH4TbfYkXNPGqmSCSosVk8nwrmA53mkX5tzJ0AEGAmrRzAGGaNRezAFKhMzJRX1n
qeHmTh1GsD+lqSo1ExuZXliJHiZK8zodR3dLFrE+DfHIWOFkdkPXT9EuyA6aHdcc
0L+7HOeRDM6FcbTPaMPjFFEkEQ/200kcjBnWeSWm6NCoNrZomskZhWwj3+We67n0
78UIa10N1kYPwTHLDBQBUmhW/qUt6EJOLcnfTQNdGvixFGrNDSxXJ4M9q5JLgwzM
tFv8ThteLxaRtMWoWGx2LaIqYQw+rlW/N5/ISa4DCkYBNFdCSYWM+dDw5f6ObR/G
dRJQC/lK1Nt3KVr0hir31TQZyrOleOCENRht8ORTVYdvwZ8C1hCUAWcjfQM04U/I
1+8gVIUFzqd/OD2FISN5Db8j0lFP+5g4LH3UC3jVsn77xuVakIP4CDLiV85As/LD
/Av3bt3mJdJ5R/gptvP/21xd6d/2qZXMeOGIcPGdQF53RYaFF1UjOc20hLyQRZeq
NUZOFX0cO9FWDBzZ17Knp8x+bK0cHOKhFK88/7yI3aNE+stRpEbwRpkZUGcQ2Qt3
DOOwU+AUQvllxkMv3QBZxjKj+yAmCPmjp7doTe9JayZtTXMPEQPrx2RYUtuj9Xi3
Foks7+ck5DOnrgvCUr0hGfAiHx2Za7lewagP5mOOKgh27Y3csVIe7qryRXKIAh4p
s7j+ZkWTCJ+fYJS8Ul2HEq9DnIcFuT1ppVR4L4GpC1oC7j9TPbQ7bMw/fFVwgdbl
7lWFrCw3px0G3xrmOnnoIlDwexGS2xvqUFTQggagf64Szz6pS04poTImqsBvgi74
pyAO0D3YPHM9Wj2dLSrqTgKCcYQ1C7+e3B/Vo2SHaELnP0XGLuB61xCWyAoqRC4L
ehbkIcU9OQomBwHeGC3UUeuySI+B1K5ufQPVjcgjLPToAjERQ3g+fZNRCEtvf1g9
XfYwYu8Mitcj38WNpXkdcl2RYGRqIxYHBhOa6kj3JRw8+jDWtkd61bJ3g0L5xVHH
ZPG7i1SoL2lY5t7+sC2XJg/EVo4r0FyfExPr0orZf4d+TNCnU2ejld3mAl3rkoC7
W7hbO5BmGN+f7A5CU1BoyZ4PBF2IyRnVuBgrM+gwbUgZ9HIKkjKYWU+PeZynoTW1
ad/tR50o4/ekfnmmzkrDs3D1dCLNzp4VwhaTNKXnakZuQruxZrd2SpIdSkYSvDty
IoxxkT1Z9+rgmgjqMIXespRmdShSRUdZ0kb5rZUoeQ1kd9/Ni9pAAcKx8NNpAIlN
qopOCrizDJogxPT2RDVKvOxZ4VP+1tTLxQ+cJc9abtI+j/Pdl2cKegrf+XWDrv58
B6Mc/Bgz+ltojYwshDryWhmdRQaVtJMIOrcn11Jm5WC4LtmJP8/K24KI0CTc88JP
TrjecjgTZufy6vlTXUv6pW7wKfJFr05s4Tb5kq40+NFnZbHGugMxfVFX//wceKS9
N57JXy+9oYnqZUeKpPFFCfW1bdZp6Fiz5suOPiyPb+6UPH4/Rr1278EawWLe5pxH
YEGhiVUO3ymKwjfzGUL6T4878Ubh0J2SqdH4nuGtzL0+HEx9DIPLXMOWSUWxRIoK
vd2tmxZQBLWqJWd+zpPa9j6RBlxrfSEWrXYLHhM0gIsL2widKSPHO7OvVXS/EbT9
ls/iKmIjK0DQN8yRRWQMG6vw7Mbo8VgEt1XyWRhAPYahyHcAHqavAKp8TzT0iH2O
RAjtZYQGH4Reg+sJzyrsDR6M3fKgBIaQgTQvNWIp17hgs6CUKd5uvHy6dZbQGrR9
ccVQmDX7szrfa2kntmua3hJyOz3iR98OfnM4TAOOx933YKs9IeboACsU2OZmC0MB
Kcp4Z4tHH8nm67fLnvsv1DHVWQqJj7ehmN/F6dChFY3kq7AZbg0Dc7LGRa7ZB38d
Caig3o1VMgIm+qfUQ4M4tIr1sA5yYZU3n+rNiBuXvTXtwr7cFHOwEcSZD4slp5rD
QwwbfgFtMOV2dQqJC09Am0daE6+desjRbggA+OcsZuD+2jq6b1ds29kX/mJTvlSQ
OUsKn6bIv5xPLlto7FJe4j5PuTsaJHwNgwwU838orZbwBLu2tPQzZlsZWW2E8rHS
6GABEkKQD2nKx5w7yxpY8KZl93Qp8LPHDNFyabNUTo/k9XQcTe72BWOp2opkDgJ2
w9EQ30iA861RlGn4mRFYaxb+MNZdPbqDZAVgJycHUGbbAn53JZ35Bb9lzM4FhlvI
WPAxVoKKLgEbyWZBcSqoHWZcjn8mB6YaJQo/Kp4/jA6vIkxX57yA+t9UFEibRxDZ
gGWWY23/jRUa04q6/IwHxWKpd5uazeaeKovYFOtK0efN18tg/hlcsL4b89hxG/Dm
agMzfwh1kqFpQfjwBcD01JT9v+Ua4AbZ76ojP6BnSQEEP0TTnY3Pl8oLK29M3287
NxW+wJ3pgTP554vY9xZ62/z5ka6w6ZJ+Thq/5Wps/HpOY0wvCZWnLyypgFlOuJHT
ymhI9S1qBgeS4vymR5k3dhG0bnIjlJ6PGGnGqmOEyp+iA7a6HErSLhAfMtA8RzqG
ZSLlwS7ipfbfZytgDxdbkCl522CeUGpS73UrdRjoxkCpElqoGvka1xinYrn/vtkX
vHW9atEqn8A1PApxov8BQW1C0QvIVos48HCS9wQRw7mIqs7ROeYx1PgyGTQFvfec
Oi6KOuSWlP/Mv6eGT7X4kjOHy76jmivHMMd/vEzknE3xhKmaru1d63yaA8iJRv6P
P7hLWIgLjLrMITg4RJzyqRwIR39I3LVhnLRg5+cAat86JyHBAOBfquweagouKQ7x
vQ6uWRbeNHADjLNt0dIWXdLNEwOkZ+7jAAhIxYbs8eUKZV714GHog4wAF+1hAphq
sBDozxI3h8k3oiQ1EhtzQsxFvBfecHf2vkn1PE9BpGNn/UNop8cs5jPI4HjSVDhc
iT4OCxOANSDeJcVIwMN/EZBbH5YeL+MaN4HF6uGg4pskAWvsmic1/Mjv1qOoiy9l
SlfdmSoWPLNWmX3rYVfO/CIl2gn+cSpqVq3RVrLRrrIWGtdUmhrPIRj+ArcG9dBI
//1auWFc6BeZBG10OY0xAfnscMwE7te0S3sRo6crtg7oFryvwqTu4KzD/rVFp4d6
IDIJclEgU4xsUGUILnqsP7l4DyAS+n+fD8qIBFU1Jd8v9qZAiPgvq/YYoNdYjZ1y
DVqCMM+lOaQKRqBUxlV56p0ylDj0HJVsv3Otl73s76gmXGJ2hT4a+sQPP4br/rid
+SLcqi1e1cBGnkFKiq6Ig0EwNSZrnjqxyvMyXc8wQ3JRJXzPDLtC9cd3BYmU/P7S
VI16520+g1k/Vdi+OFDyt/C8aHfgedYV6b5U0Jf2gm3G5P/Gs8POVUx63PTPC3Q5
nxt3nVCUDMpjN2iEeOrttqALuuiLBK21HNk7vLbuzN46T1T7Qwfx8ix0GCpsvq8B
9nM09o9OTjnHN7v47t1fkvsfY6bmSpuop1i3wstjdBJOgrh4+2oI8NX3oQXPUSfG
eHiRY5MvYGiAWM6Ji/X/781t5GRe+3k25yhoTRCFTnRNXoodrIaA3cMzg685CVvX
ESKE3NiklvbX7B51uk2W+zkZKamyyB2zr6BxRZWuZR50DhNnRZyfwkcGK4rnp9Uo
DSvjQOAvbNEy44bvq9luiz59jXLTiG0I9vT5q5PWVzt2KmlzhZGeQxSidSV7/CtR
mASk+VgavscWkjboiRp8iZCgllkSGoy4mHXB5xWhRAV7DxJoXge26r1HXtQdEDkt
NIJFFb3v4v/TC5D5AsHQf/wbCH5SVmkAnDSs8qkYADSQtwvF/f2wdMfGpfmZE8uw
CtNAi5qTSawvFk0sujAijL3epppwGncZH8xXRTF4xMASg1fnnN6WcDwt5GbwX8vN
2gucEn2ngkmSD9grhm7c/blzl7r1MIHrMypG/tZddsdtsDEznCsD3A+m7usvgNla
4Xtx8wbjcrmuJR3L4GlPo+brlTxl3Rrx7DoltqEL3nrrXxTnpm8pOfXtW8WF30UN
+WWYNQV//5GEmf+Ix4MKE2GRWOUZZdzjTKIaalnyvFtMVV0QFOx2zOd6frMjI8WT
VqxsRWFeFbqCik2MioSIuH8mjYz6DWJ05mlBHSsbwd3SJViJXJ4Y+uQ1GGsDC/iv
EhKh1D6cQrpdi4s103znjWOLjg55uKBphvLNgZvLGFJpm5LI3T1Y99E9O5O1cY/K
De4gq4xPC2E7b1A3lwdvJjvbb+z2l6AaAr0ALvOeCIQpu04A7774pvbXtJw0DsNk
NB4FpqTKuiuQf0znNMzANyx48DX40Ym0Oq7FRtr6LQSJjAdMJ3m4tp+XCvgMHSB4
yzu9tYTaMJ8wVXc8fpyqW2baLbWurLHtr1o46wrgLLo40uFW1gd91CEU0/fadUoa
8mO+j/G8xiwi+em+UumEw6clmNh7WlhBW6N5KJt8/D0FWzzG/BqGYlxtVTUXjqPQ
E3RSpjNEiBpTTC3tPwWwlyGhqUbI4v3b+fz3F/DzFkv3eHvI56LYF1i6R3kfOl7Z
lQ5uQRkn8yKRXTZrp8zGZJjXWW/+jx7cyqX14DzuoJnlubuflIW4tB4nLYOLeCHN
mReexejag3o0xf05SjIXYXISx7Yp8GH6LAC04FF9us08KOwkJtYvsDpnsGzos+e1
YUv7OQIsFFBw8/zficJpiQkLAD/gialk9YAp5ee/MSfV3IHfWK2B0BV+VEG/Idzi
Fosh+y6YH4OnMgyXoktt1REOUC7EL93s10o1NkyZbpemBE9ifrNzMc8WdBe99lno
a1DT+JTANSeKdeC4kGvCU+IU8m1CLpBM26pYWSXLJNrgPMna3xZYNTD7W0d2C/XT
5rxdBNJ5B26/rghPRhdcZW6E+t2WV8oSOqlTveJ9yHf5SsGeAhhC9h4ViyqknJ+L
bPYXmBzdKV+U0cL6XggaLvxrIS3iWl/2U66TX1bWCBxLxVWv7ceEa6uk55MofVIh
8qc10N2sQ7TEtxFgwPzrq+X4oJzLb0pfenpyX8Sh05fnmKs6Xu/YhDuNNizgs3E3
6OrAP8VqgloHh1OVF43hhGm2Hwo2oC7wuqbhj5ODN8CHXP84G6sn5LpkvWrkRp0Y
B6MbahpsAUGp9l9MgJjyAMLDsK84ktTwW93snvH5H1rCvC1OI5/wo19A/FIli/Is
eZOKl7HRezRqrnVycNfPyhm9LegN8/hKBCZtcqLbnbbE16P2Mg8xjOPxGTTHBnMf
JLp88XbdVPoDKZfoOs4nPyeirHS3ZqGkpefJW4oSh8cDp+tCyR898PpQzrYIVQo1
liCq4WMZmM47iqnFRW1jr+4sr29cbEVe/J+T/pDMPpU2JlKaBnYLuLpZNLwq1MyK
ceeRP7O15WSOaYOQFJdThQNyjL0hkDXgyVIhLp/CkRpWtZFE1MhtGOtP4gN0jOct
5QKthQZGIaUntj2ZOioRjhreoyuonzdFJq/EoORnZEUHWnXMT6tRBd0ddpj2qY37
Q2BQkzm+spVIxxc7U0qr4/Ulita7De1KxIUH3fbOzim8KxrfhYVqgk9RdJgdJeWu
JKTLgEeobF8edCuKo9sqbvp8k+/yymFSfwnF0pFnqNHK4kXbKHb/4sfkLQLqFQQ0
hub6xHJeyFPl2DcgT5skjCULudeWXztp5yReaUmM/XtaMiSZkUwdnGh6qTYHiU1E
nw6xnS6FxtYHLifI4ZGL3EqIU6KKj4+hiIG365YpQftgAtKmSoRr0YFlRbtUC1I6
ygDqo92wwCb/H2atfHQdGqzT7z3D6zI6NfptraavtvYyMZFVr+lQNBy83MvtX0qu
HkrqHS5IU6GtPhEDHP2USaVRucvJgpa1K5dXSl6yv/Kc8uHWeMD7iarBGPQ66NBP
1mbLRtwa8qMSseW9QbKNNjdO6ICSvnS8cpV1P7aXL5CUaboqJI8nYtvMlEC0IehU
mW0E8P4xnFGABciMM321ce32wuhBAz0c+8A1s+iLg2jMuVnND5LygciWUVuC0K1M
UiYgxaxvY8eINDpskn4lTL/S3KR0Q+wX5Cv/gabDRsRzStTVFnOitEKYxI29wgoP
708IvuvKVL3nYYHRUFe/HvnJ6QevyOvc4eCyqZtu1YjaC2lCmWM36v9moXHCDEtk
e360bv38rC5uvXjfTzo51HyH7gnigMpU5VdQEggTCGNjHYPAJQWnMZLSMRtFnIne
CcRIqiOm2dTfnL1eZVL3WJJEvOdgjshO1lUo1B8zMVSbg8uJM5+RLRG+510c7HkG
LouqIyJ0yUIZQCCvhb0OKY/WGCBeaszjizHsw5mr/yXYwfW0GskxgALkPrdKwqdu
tJ9hRDT7aWiq4sFJHLnwF4q2t6irO5yVJw8JZx9NpVTEMcAxTOy47f6Uk2YksYbu
Zw5tQ+RTohTfJu/H364jv2g65WtPiX9UghjxueB3xsXmrS0Wz+UqfGICvDDri6Sh
6cT6EVBRQvltDkD1gAHAWDpeI0ZXm4HWnWzFfRp0kaY0O6S4AI6fJR1w4uTc598O
tORFP2M1wqIqvX0ZaqALThj11TUky/NXWa2tblEh45OEMddgAS8+t1wyIlJ3fTqt
ImbEW2VVLVFUkfYsmRbTepqQXJ1R0GTe+0OGmrp+bk9JdkSUUT4gwsIeUk1pK1J5
QOi+nmwGV4f14ZSIxqi6QVqFVP+ZUZQdBHj5YiV/mGL/IHz7OIbOnsXShUP6XzTm
PJ5YVZUG2H5zwqXyOls8DP0QkeBcjqfJIPIQ0bPhWTIlH6BkjqegLVaVjZynxuo3
s+mxJmYuiUG/79KZPVco3UOMXGmwh48uiYcUTXpqXJI8/dFUy3rR4vbvB+Niz/vE
IvqSRJRv9+q7EoCCgtjqkSRC6ov3vsp/R61ffWH2GakfNot/iAcr5763SesfJu08
E6CNJEnECkok1zmxUr5MDi24HqJXRnEOH4ikAv3MPwa+P2EB0vXk3xxtijU1Djvk
v1FODdq8POo6gINUjMb5+bKMuA4oYuyEYke2cru5xe82W0n+urcmD2B47c8uao2/
UBQ1L6MLamN1oUDWNS9bHsegbWewLJkrPRnDIDLih1XHH0fWWinyhiojKpCWNymZ
vqGZChugknIETAe5QxQwml1R/RqbWElEKeMWtW+dOJTFfnvE2Q391WivLtaVII7f
XAGvl/0EPGIkvVUKEyMtpAjZ1NyzxrkvRzvzq91QXqQBpTJHo6CcrJF5rfiSj95L
2Lbh08IV2atE33HZfHwHIIVxpuWkAiloJAmxYGV9jD0yDnYgrTR+Uv5GgE/12rc1
bSKF/twYCWTkQ5sZnq36wIH4dZFhEC5S0LXyl/bacU5czM79WM5Yh7aI2glIauqQ
i1sxnGu/pbI595RfpM0V0zPBQ5R7sJBTjppg7moBj+9Hkxt1KR+uKFbSMD02Tzqj
xc7Tm9GzybcVrA7b12ngI88sS1WuYsJz0vHGSkjMrK1jWshKA4Lr1yGqc6Rs2eav
gFJ8Mv/h/HUyB2JOTNVhE4SI+FVlNogAeCR+7ICgeNJfvk5/3kBKYgql0NxHLG5s
q01XoMQff1F9jC6MOU9vruXDSRCtUev8YePIhWvX7Cu/nIQMMek9z88QarWlTeH8
ui77d8SKuRJv+GdqYZ32V4VZ+RTnPWCDM6FBg6+hHXzoDuF7Ubzh2j1NN4LlPUg3
cWl9PxrHeclQ8+6aq1GLpkI6Tp2fXnMZgFgh09sjUBZwzUPiSo84ulQmv4VqyoIW
IKial/SR6kZ1ZqMVZWkUZxBGraGnyNfd19NsIFkADDga7HYOmBMR/SixNnJSpw0s
ZWR9pQ70U/eRw79jjNYnV/EYdQ9jhI7kyjaA4We8cOohH9KpkfWvID5WTzMd2tAq
bMJYYK06KznE216siVSYp6lz5QzwpDLiM3z6LPPa3OukUs2Np/yp/kUDwTPnsJKJ
Y2uq09i0viTfVH6HgDz6JDu6l4cLljM6YH884A9yhlQbLBl2xFP1Qq+UfrLUNJTS
BJhmvMn6VP42AttXpvZtvhPZIO4EOc2Mi6OSgy7ixwxVCtMv0edLnZuWWu7LTcww
JrsNzfLbKLltUByLdF14kD4arNjbigBBG2F8vWpyeDUrAL8SaZxG0gYjIv5oscY6
MrQPc2BDA7oyB9B52OZJDNK0eCq2sEno6Z8UMKZ2HICtqZxblyYnO7eqHRLLhadm
A8wQzQluvdCuAltafDBCEPcs0z2UDeBTMk56OzseLRSTnhfDmlRG0myaJ+Ke2bvA
YllXQEoO4WIw1/IdO+VvdlEuqZvQRq7K+AcO6HOcfijOE5uHrjVF4KPWVNptPcar
We7JUWW1W5kWMTERIKmeEDxrdchQCT3bgLNPZ3MhVpoeWxEFqhD+U43BKP2jd6gh
OZqIjXnFsYQoV40xO+nF943tHyvwWrft16R6RwH2+fOBfhZV+ouv31DUxOVBD6gi
CaBAtKrwl2q8dA2SCl/jbCazNBzbgG7ReI2fo0Ym3QReRjfvzKuobgEArqJRkqAu
HQLA1PsQfKjHRUWdYFxqeSlNupDfHruKhrFgdwgbCfQBFwFPxnWwUQAk2+dRUOLF
aWlbZ2rNcARTwsiJk8P53HH6YHDO7pOaCyeEzPAAiSUUt3ECm7/CrXBLM96/R5Tu
sP+iWVg/WWanUIww5XftryR2MrHrcrqoHokm36BbxPjMhvU+KuqBz2WmvvCru3dq
rMxhoW7/lMZVttmjAgJxiaKkaMgo5E3F6Dyof+pxpAMIWe7+mODBkErZqHab0HGQ
5BgON+vhRnpfZwUyPmWKzr5YT17oON1RP758B4oS0sJLPo99CbG0MKkPf9aRf/jy
JMkQW4FHAd3fSTKamBzJCvDnU6uDjoohgRod0WxuFcuSfd7HsLy2y8X3CH8lVe/U
UUVAOE5RebEAtIC1MPngIbA1nkLpQqKb2B2SOaQkWcPNHzblSrZpmLEjh2yd8Bp1
mKwJD/xTFPIl7PmaC7/iPIEtdqASwiBsG7/c/DBQcAtNhH1fDQppDnxlvf8EGCZt
u6rDNP/oGW7AK6o2pNrQItcKJ3yNc7FtSOf7DwpCaosvU6ZgxCKNSVvT/A+vN2US
YJNgmggoqZ17LJWO4oI+uYVLjdYo5eNliRmwVgkp+UX8MAJZZeRSuOgqILI485B5
m/9T4WE5iCTFy4VLkmKDNUYB55pCrQikqpdCxeKxrcpoFIIuO7HDFw6PVl0sUaM6
faSX3Y9vqri1mkhAMT3WjUHOJdV6W3lk7aPvzVDJk5E9z0+DcUTUrqo1Dt73iVr/
kYywzs3KP0xFfYUNFJoJczGqF1k1sAL2VMRVylQhVSz0KGrQ5YxeR+hDXgFdXKPw
ly5mC8j/p56MsLwtBsqrdtma1SwxnrBiyqTI6s2tMq3j+Hocj8kvin/tzkRHiOy2
yq3Du+NoJznqnhTvrKb+9rHWjOvGNRxYAJDwTYOeepXa9vHefAJ6Lk2lLjpjbVix
eDPPKO/gJo+KfzsbUWye4idFCna6ZO6rA7Q98EcgghWryGhpCD54peZrBxWSXNuA
wp9lQbvExGc2EoCPGqcuOmLgSnXr1qVuDHC46ySihzvsbzAwrT1mr6mlW8La06De
VG1OFiB6hx1cyQgBeQNcP/dQYZo05eHj+T3EWH974fryOkTM4Jez/cLB2PVp0V3g
qgi75FRCjRFDvWm/WEbh4A+Jb2J1abkfyTXG/YHbo48uJ3hvnEHfJbVqAx83BVAm
OLFJ5WhHrImalNfqh0iTxvL8vl6yJPf286rGlFfmdlbrSFUvLkXkYhuClgvIcbcv
zjOqNp4BrexuZ3PFP8qJzBNYvT1tEFF9FWj8wYfIFvhpRu2NbUDHpGulJ9/TD6sG
MbGikIarNDGxeBhpYfJjCOoRKcQtJb+fPymXRIq5/L/1D9Lgon5PklIHzUJXyMw3
WMQQGQ4AWa7XnP5Mm9P+gNq27g9erBsv2RNGWmK/0+cHFGiGorHUgQ2zAaxCtPec
m2mscBzXnyL/olSCwx/wirfTSQtvP+tQ6isQpL4B4KCl2N9bpfNybdEo4HtlL5q8
XOFQOCjWZfrTlttHwN68lKZ7rGOk2aHJskPKTM5WnI5lKSCheg4J4JBkHJhit58k
J3LljjywlLCZ1JkIrKuisZOHg84r53cdQqcfnUqGX8LutHdasppgx7Evp6SV1ed8
N2s9xPQkcJAL/6plNK0a5abbeTPyK7A+6/NnASatnRUxtBTuCOtWx07LBObhladM
zYjzw6G3ymOYw5QKaps9vuthIb8wl51bWCzVn33hKATpLlC1o05IWozIJJ5Vmk5L
omFaKeDC/WcW7d2fDw/5VA2U3BeJSNB4ntmiOVb1UKiFL8eAUPFDCZeQQfEZsOJf
M/ncGsTgGj7HIYGLEmQsnvAndDzQsV6c/pLWNnjVu1BHBOXXWtFS9Xg63uBihoc3
dgAmGpAy9yBHwV772rBOza7arBPlz86FUTxr75dOeVVb0NcorMa+VQI436s5uDIi
vYm6Bgz14kt1NYVZn0aK59WK4Y/88Ek3b3irGDUmd4iXXe2XFqr9jq6Q1drU1Qm/
0BZ1bEJHuK/3zy3p3uwJXnYch5K05tHWA8PgIXKfoV/U9uXgdthAgfJzvUM7L3ZC
XO6GUYF9VHn9QpsFzDumQIBS3heyhe1Jse4jETa08efLdMKLSz9CvrC3b3Ak+/kj
RQDFzJfKr5BFSH9HtHzLA5SbHOeUcGKkK387J6JSQoHG4SScQvfuTXlzyPuOgrUh
N5MUMTX5rMvo6xjpyAMVQsy5a+jRHxlzUGC/BYw24m5XlrrIbbHaw2derWB1gL/S
tsqbg7FYDlMvX6Tyh7eln0s6V6TAshAqvXWUfgZ01cX1EpJkaZ0KEwFq1pOFWs2n
wqFuoElBUepqqaGL/Iby5WMpFoqaB3xDWmGlB63bq7fgdrmKm6kruywPJq5hlfHT
zWjak2/SlJf3wFTHPRvUyWPbkT5xhoWcBFiVV18W7EYm4bvLBWSgi8muVck2EEES
kBVgEV0OAPpUjBtxucAB62BreI7ugcy/ksVJs7W6pM8i4eSAQx5unoSlcyNUKibt
4fYvJUnmRsJSTxg5k+LAzFDgOQ+L009yUCJ91K1386YM7+sPLz1hoAn3aBzSo5r0
c0xnWsxyG4R48qxwv/0EL751tI1KFQdfnWwSf+CZ1qQLf7012A7k6LcauxaMQ/3A
9q3ixPqgJyCb0shDQHq3s7Q1M1CV4J9Gr5QSJNSsg4st4yadtgoGbAOiM50str5o
Cen2IUqbi85gah7Xyt3CHZo/91n7248Nzc37qpHcIXgiatNbdvbV2jw/0Q6ELDz6
S6GNZXZtMtImvbVtuou9SkcLsqswNn1Pc2MB1woQuY4QKEc0ak8SbvOVh3kpY97E
0Gm9WuiW/okC/x1vreYs0EN9VviYjgW6cYzN7NEqESTzmA2aTM+/NcXwwZ7u4WDh
eNdNgHWO7P82A5HanLM6fdG5Bl90wVRymaSEbRrPNclljCEN4/2IDxAyh8LSeEyA
XLXvurMluudDNyQexP3d+zZP9w8NamtLtbOtdn6Crk0dqWPgl0mObBSbskgOGRWq
M8aJ2yO8Yt5MMNWwX/P9aFBPJ/ByaiZF9I7/KnNqwdf/UwmXDJGRBUKku0ha+UdM
/3VAU/XMUVRmR7+pK4EpHsO9WRc1BFFV+xaguMHqIyk9G2Fs8LIEqxebZVM0Y9ny
c7M1iHydQn/hH5LmFvbj1/oXinp4VuCpfWpmswXCfCxrkeosBemg6Gaiyjxl9x/R
kz7BSIRXd3L8kql6AU5sf6ibI3p4n3BFeOE7QmkHFddShH8a1SNuHzDpfJm/dtQp
uEUaNJaWQOQR2zWPjLZPFmo+oUy2AUpfW383iGfgBcJ5VmsngLLbn7kj2uQYvOf4
yeK4P98AtOoITUENvBN5Rj+r04H8i+ZjMGQquewiUX9UdIcQOd7YDm1ayF6SOeWz
qfmSAVaPB0d+7euw6TslKizdc+O2t4UbRMmaS+JGPXJpQHIbLrOc+2MHpr9K0/wW
fKk4V6AR2RUBH1fkvhmXv/NLzQbweHV6mGDVzsaZ6TkkhaPHzna6yLscZVL87FZr
LhEqzDbdogKDQx8NKQ24wb0dLgeeyvLFkGzWPEz3aH+9a/I7tzzXMVr9lv+gd0IK
VhhQedRMkwLQBQVHqLXAnijI3HfDf2Qm6zZbg6B7xsyOr0lg7AaGFA2A8SFPf7/o
tdQvaCCUCXnx6cdzgP9KD9SloArS68+Ac8/sgrsGFWUqx9e6CqdXX6OI2ckyVQEh
yEuVpxn/YSXJdhVN4IWcc3ky+9ImcNxxY0ny037b0hFtrxWwnOxJVP0yoMCaV60u
DucBFka0Iwc2rM39LSd6yCpUdpDN1OBJjDHgKrb1diH8kiok5pgtHWqHt3cufMi3
Qo4db5PaA4esBgxtoATsUSpbBh1pojaJ2hJB6+HU2m1syEW+nT7hbWXobZPv9DH8
2p3BMQqTs0O+TQxC2ZS6sloSwbe/7OLYKLWyHjATcxLXR45s1M921j0LcBCAWoXy
CisEsnQihSY0SbORaJRyRjNDE9mowrT83YGsvA8XdOdPxLkVybzZen7pA+M5tR4m
PbyENGLmaF0OaPgaHfogfw/KFNphJa/j8pn1hOSgfxc0WTIEoyxftccHn1VZ30Ye
x+qsq1KMCbdslkPrNREiQUqL0q+BaB7uk8jfrf2De57izvbZbqwqQ+skcK7Ibzey
et5l5PnUKy85pBr+JyFfTO8XdasthioytScKOTZ05EMJOVOE2mU6KeinvjyaRNbm
0JhDdQH0xWTOcj8p8eiKd0nPp34D5omy7lpK+TysQIBaWP0YEnp8kxZlXBxQb5Ls
/zFq829mKKg989rbQLC00ScbkH8GkSzYA2JP1CEvtPjrK8xKw2Im3BCj5ptgcsQM
nO8DmhaaVK9gvY8niqjR7ifgT07iziBCmTDT74IPHbkVJhQre0c4+GYVDci1H4Ju
G1qQ6YjZqgZL09RyQN7IinVdMTemSCMaU8W+0BKoHcICN+IRLaiQCZF6VGPdjRgi
EoTMGNUF8M68aDpQzg678p724Mm6GHrcT+Ma+5n0Z/R3rug5k+kfECKwqmnAONgG
avLhn4hR0RqXezO0Gk2rQ91shzuHY7UbFQwBfUEicVWnALb2IU41mOOWVGvUR4hW
wtJpTecgMEW4TyjRsPK1P7tkg6ZHfgwrI5z3RChD1eiUe9/q1JA3DpLY+ZxjUato
Y0ghStKPo4ie+x86ckHOkl8lXvPL81u4Ajikye9R5EDNF0sl8K/DNj/pD0rZcngk
qsrASW8R8MqHMkLFxmxrTMHVof8XqieGOLJJ9UYo44cpjKx8E91Ob7dh47kXIjZq
7ZEAiIuIfNQSzYtOn4CcGSooIVf+rySY4tJoxGZQVVOqqiWA4ORoeYWauDhLvu5+
jSlfqKbILruQsFJWErAvwnK8AwAc/HnuAhJyppHETo0q5YDf8C3ccSEDvXiPEja6
YOgP2McFpZTWePa+xVRTNxyGmFW2bciDI3o+rzbFuC/d9oPntBskmPm1WdBDbE8x
mzEyPhG9G6NctaXiAwLCxNfAxf/jY8M0x3+6HjuBRAW+tTSue5N023U+IA33qacj
NmF8LMSTjPm+rfHZFOLokv66BLuT3zc1itcAD0GSWpxT7N/fokDgBL4u9Xc42D2D
ktbfwKxe9Y6KLLqDfLOZ3vUr2hWV3EowuuopeIfL/MHpr2hcLgSB0rUgSoooL9ax
dZly+i94vpdXIVAi6BMtMoWmsWMfiWLoBU2YIVjh5qVcdIdnXWQDWk5K808a2+Ge
pMK114kEw5lOSfNQUKmRPS5oiBs3C84qtQYtiiOPrD3pHQIntRhRxcvcWGXwb8Et
IwBgdOEWEJy5E3JF11XT86BZWoigL8R+zzQiYZum6hR4rIXgd9OIQ6tj/eZlANtr
HDg4rTGGKw7ibMkP1CrghrX9yS/vuE7WSdddgccsB89WH8IidaKvm8z04nWJShsP
YTF8aWIDtT0IY4poXp9IhZ1Jv/3Vg0Yt1dobJAz7QBBBWj8KeHCemlm3NPHdSvKa
GAHIWPaToh6hbSj7nJbyQTHlDO38Nda8qIM6QQQbla2pMwLIz3sHc4SWH8xcYdjW
s3c3jqxlFzu3hrnfixtL61+D8nHP1B1VKassdMtdsMFg+Toi1av4jUKhOL55+aNE
H28EhSmQqg3oz0C3kS5oiIZCS9RXjxQ18ZaX/PkP/aKY7mAV8Vjhm8Z93VOvmsFU
da1TMlXOCZWklFWhfMQSU+zFeV8jiiogm0uA3inceLXX5Eg8uWowbeTRwlrgkSja
a17M+4RKLaRkhslHQm6dzMBq5NjmkbQ3STNRgSwc9w0TxRHXetjcZ1Q2H1NzV9M2
RXN7rjjfn1u8FRp0D/T5CQKyB1KitHnsraatz9uCuMTybPgM7gxo+cKzlxOuv5Yc
KNePW37MjQmFXhi4j3n/gb9CTZKne654dh1Xr1ABS38A3uWkcBhvFT1yCN2e26pS
4XKvbOZ8fnTMV7krhdpeM2OtCTnBjZAlcuyyLy2Vay/A7kP53OWGJ9l726CiUeiy
rWp9scgVH/viJWrjlR0vU3ghDJzBLpv9oMS6gNumaHImV6ilPtfiqrS4htXWnnDr
Jplyg2/zb4HvkxdxZ2KvxOAgGc/ri8QvQkRgE0pSUCfRDLrHT98l0r8rUbUxQB4j
i/fmOVaKHKFdqywBkQr6Vx8y3U+OFzWenVrcvuFUNf47ZW1jk11cueTzrDwEibqp
Ah3qd0PL7R10vofJjP3+4N7bmZ95QcOQrW3Jv1L++sd9CtlVqIjQuWOXgNW7HyKF
sK3xPu9i3s+oQT/V2+Nu5LT/YHVyMphniymIv9FduriYDwJSTY6iZXzwkaHXOk7v
XLw4u4TsEwTiumREw9prVdwBuKBCdIRsmX1NIVu/qm9l1rHTeWcezWIWir3Ms7O4
L2jSguNPq4wHWciFalaAIPXjCKcjMYv+EpnW8eyOkmPlhua/E6WQFWsoZOlKY0Vk
4CDsFPnS9FvDfHxl3Zll/cv+ZCqmI0vm50fPAYrCxZFJYjAj2b8982NSFlEFoM1Y
igCehA5WtP+/A0ZyczL1l9Qfy8Uc9IjGCf7BlMuV4oUpbxsL7lAMpwUm28mD0sih
V98bbWUW4v2BXTF4fiLH4tX/ZwKhwGGbS4iWZ28wFSdJk+ZGAD0U7QrJ+rgCRqWY
Uc+E4VrG8+/5fJeoRsxvrcBhBE613E997g5G6tn0sTX0In2ytEJefDzuaDrhIwvt
WxxbVnB3zA1tPOFzxVqqKmLrg27esUl8A7o/5ixAnCESW0q2ZGmOXA82JEfpunJJ
WVmcuWtmCMYseo2HJWCiZ0s3jdG8ut8lMy5x9nUfDUF4kDWJNNtpGyMLaKz095G9
AClXkd96OCVP+w/jiqxSt5xP+27AGyEaOjQtE4Yjg5eVqeZED9DcrwLkuYAuWxRy
pWZ8LBXedtO2gReQnGrMOesQ7nVqm3LeIFD0lQ9WmJ1Xv5uoI7/HIYmeFE0OVXVW
0eW1W0cfhJ+Z+pE5fXsxq6fEBuNu7oZOkrZMTY2CsQ+/1Pt4tyt6/3/DvMViGoXb
38wqbZikubFNenqb/qjNCk7r1mdmpSXV7p3SOdg3KE4kHmtoBXL7AA1qsvSoJJPm
mqe15TyN0MCQfFccA11bEfsvj0tklhA27+dUy8Qb0ZncZJ3KrpLRQpEMBjAaQGEh
VlA7fh1Y9cZxUCY8SNo1Uka1fchxCY/xFcK7sEbHhSK8TuW+JX7fYuZe1CBA5Gc5
PaR+7HuJlrUFEMw7QNkfkrNfMWUAvBWn8PKOvzVhIJv+hJv8dKOZollcqLjq4f0R
hqH29rBYg56bTbGnXclemReGFsH57k/I37tnIzif8bGyseGlBC6oC/iF7FTtjehc
E+hCMFD+nTb4E/aq6Ss0peErFMPFwG1w1n6xYCOicNpBXzWM/4loCKHAwCLxu8rW
X+kAtOWVtsZDbqp2Q5c9cTG4GwwNuwJVeq10+tcniXhImV28fX1VW51rktKvcq/M
zreTx+l43czrkk3h0rgrUkU/ypMl82GFm4udw5Z3437TqrVc0v9r0ffo7qRXPqVi
VjH92a6WKO4Jgs5csfrieg64r7iwzXFKU3dgNoiAp/9zNECQdNXAlOcOQuknOwjr
rJsBnvUfTKn+sDasDHhUJV3M0M4otgB8RR/E0vj4U7FpqxoVLNjATA0byKCHZ4T2
eJltBLZc0xbipByH6lHWgsPvjpvT0fIunRfQcfABG38PYkAzr2wPO1uu6NgBUJST
4Ou+NolphFxcWxqiKB3B7A7inu283vxaDqrx+61KaNUOVq66q2WALVRFqo6adtl8
4P3/TVLFeMOFyhXp5kLsoO9letRGrcQDQi9rrrivQtqJeoGWgGhYif708lAD24Uh
erTA2u2/SM7MwMbZ7StpcKfYVP4AMopyTrWz04bJ6IO2veegRZjJ4me805U4w8Ew
8yEW4AEWF10EzqA6kMwOJHplcsPKPavayMFvckaXG3TjDvpqZv665nYyU+0m4uRo
JG2jnPhMTygWBlL3vTjhH2VhHaq/nhj7KLD6x4L9ZHtZKC//DEO6F5yZ5pIFQxTe
ZqqHYu0g6ULh0LbOOTXooL/R6P0VXBZZ3BPCHGS/rWU3YvGDb0wpYzJJmr36Astz
lmbPTmfJ9NTJAicXuGwB6J/BQkgI5irox6Q3CQW+lDrh2e1XicZJU/KO5QAnF9/l
8kJ/b+Ox/ppiow4pIjGognsU6FDF4JORCCLdowfo9hoHzS90IO7U4UPD6YLzIqUy
kA0YKzgMRcInKIzG+WOjYwfYzKXXPKuI2GAsK3vAzqoACFFRAfGBfCUDk2y4xukB
Xj27QNtLfVKa+6EtTaS2hykL/Civr3IPPa8gYNvisqFRHiL9whWVeRynOo29So5U
tJkWMLiOYWiBoi19VQl8CdzeKbE7UQy3sONOP2DRdPUnXmO/jQJkYd4kOokdPjxX
ZaNTsf685e6Q5+3QxcplDSz5kFg2qM1oC2pT6Fdpi/ETR7KBITo+GA+zcSYTF0He
ehuLQH43yHG8Y5eBfyT7iK4i51TahHfY0GvmRMs1xbnJDzNfxuRPZHr/ap3TLqDg
z3zfXYMWiZVCZWDmJjlX57iAOIsCyj2Bjm1WREmk0pLSBA9RbiIcYB2dQZv/ve8A
UtZtE/XgfsSsx8t7u6BuCYWByf5YWt0GU+JaREVamA1DUjJeiTmtOFkHC7xohPUm
CnAXf2hBOCQVg9ItZHB4lhibgNi1tKHbWmeVLrIT3t/mgdCXheko+ICKYgGVummd
7yN+3ZFtJxjKwIA1m9Jk/Z5xm89Pkn8fvDfpbGWOZXYRful0jBXHAFZMBbZY9gDl
ZM9V9jO4Sgg/wz7Eu8jIN+iThSi5pZaSjWQXgwL9f4yXQxZFtJ6tuC/HCkocl7X8
1B8BeJQ17ELoLPbpLPniyIKUmGkOU9utQuc46gqv4iyUNeoW8QvlTE2a9TTdxemG
dfCnJx9N3QXxSmIJTjvvJFn3IaELAhDXntVPSBhXjxutNU1ah7ZYmZg8f6Ju8JAr
vh+rbszTVTWUioynttoPCvce7C+8IjUFAA9v2diewfAeJ2wZmPwXkSXLUEvPiqHh
jiPA4duZTEKKtAflqQtv874Jf7dAec0rlv/sTlu2bZ91asWxaWCZALW+Fg7ERP+N
tKSQRoTgfkgJJdT3u78gumpho3pru0dWD3gyTqtpU+Nt2dm2y0/8V6OQG1L9b4G6
QeZ4p7LK/ajn1POm4QSq1HuM8rzy09FZ8H8SHhDvpgq9s/HBRrUi4HXUSVqTxjip
me7zEfTqinm3PeSmhI+LfE4WPeFnu0ylas0tfrJzTgLglxBoOh4C6oEIPAxA0Z2C
5vwEXIfZTWgQOiFbrCZNGCbArPI1Huq8LfcWQRvvvEc5wHAHLpCtAl3yuTeFKzKn
PdsBgRMrjoDpdZeTuufZEO+TgcbpcK4ydktDLNwus1HG/HK4irUPY+NlqEemeU9w
/RgIEQeax6wrJrmpx9YJuFyJ9P+7roimm/cU//QbmMxSYyM2AbCthOG8TM6HKR4p
qujZ0zJmQhncGo0GXaUcPfF0QaFtNENnB0kj0sfIXRyVswSfeE7smtKlh3VylIyh
bN5xowmMsnm24pkM45Gm1D2QcJzA3S/mN0TBtp5BZ+1caBkkdJ3t+P8/e/Owh8el
hMpvorY8L6iKI3Kb8qDqHjrEqoMSP5nBdc/NuSS8p6yXtdCunCrYqmdnPxPuJIaV
8MlNKo3/IzsPZ41moxWMoZE28zL657HOyG95R1uHCDNeK0+pQv3SsQqckV9Q1PKM
S/BB5QYTXY3o3vsrC0g5EjFGvooyPS/AhkZpdpEcsftemofjvyuAdpnaA5brXAUG
8ma4Y2d2e/6bIS/N8aRpiYbPOouDEN+LiehubC23JWqps0R0OTlUMrAg52pN8Oev
gNf5FbZKqHafDBk9qIbuaQPBTTLWiBvioFDVvYjvw52YIwyuoj4l4oVemHK8JZwn
Ml26EDnSvbWJz6Nbej7HtZRSrCSAoJyjY+Fs9gTGdUGVqa53kLBJWPeqqXYKdT+r
1+lM1EqjLYNtbhyOTS2+2gK2oO8lMeTBq1tIhlmDJgIY1UlqCBcJE/83nA1Xlm6e
iDZ4rJy0onHTazaXtOfH2n0IVnVEc/bWsfpK72+AThdUvRG1DF8yDIOjOv3uyZNv
L3tKwXb5ffuyaItFz5tncOYB9jc71h0Akj0pexZgdeSMUduA9gn7gVIVNHNkSV29
DlDZWmsEfuMBjrzPSuBj8NMzYlg8XAzRkGAfm+dAaHGoqzbhRgvUNw1WWxH5cpst
J0ESw5u101pq9LLCZ5eID0l0vn4cQ2iIFbxV4awxv2b4h2aI2FayiT+S0M25eqQG
hJUx6sTu0/SpmlU4NQ5ENF2OFB9MK5INzHb+i8hndjoBr2DtuSZb0rxa+BCdsKZ0
y4BdhqFxP54ZPFW4ogXJ+y2/aAxc4FD8JRbuLJnLF32kzUavapXPUuQAttoiW0y+
KXtk76QDiQdTJcSEHEd2F7DXsKpXYcXlusDdBafm3pQffirl4w7/ereBdEUmeIaJ
1eBWnkxmL4N+fLt1ufgrwzPVFHF4UkfdzrzgJREpMxr9HjSTso7wtnt72MN4vRWd
FfRNydXy2MOEg2n41MH03jEIwyXKCkW7lOQCkYNsZP+GaQBkmJ0e+eeiexXPAP3C
8JqHVOdVZeOP29M150+/fQHpim47xXBRRxOGrT1InewjhoN1b2PCQO6KP02DXt/u
VZF9We7oCFZa4fSH9uasyGMUkRw4fTli6IC5ZLkwdmwgPqVUSeQWy4esIbAEVpdV
UJ3mv61eA6p/wm8Blk2isk8TK1wEfGH5C+4/RlBR1J09n95UBqfHFbHQCLieoDVV
ixxj5R4aSd8lT4hmoKIJSDum0e1tTCPYc77SjHWMU/qTx3lZO1vtmY7OALmQ9rgc
mmAPCrIuEGmGDlmRu2AI5Vxr/dE0eRjL8Kd83NbZUfC1JqFES2IqZ2tVhkzyWLxp
Ca3k6y23VA5SuiwI6bR1xLAN3u2PJYt23EXk83gCwFBKtYYq4pKu/abHZ4Sv6Qqj
1gLMJCr/0Xwr8iVPslsxxi8RJT8vT2Hlx7YzHr1TKtK0XSe3rOqFep9Ju8mkK/iH
b5AzGXc8UN5fyg0bbDgWB8tcaAZIxLfDt2uxQc0c8NfM1S4nW/qXe+WT4vYUCAKS
QO4Az9SWwVSgJwMupABsJqM017e+5UBP/I3l1mSe/K+Rnyy1c8YHUxkrWwZXSNOq
SNcEv6tRdY1kp7Bsa4gm71StCESh2DabrgBHoamCA/iLHBuA0YDTfK6B+JsPnD6D
u/RsHwls3VX6yP23SN6HNtxhWTT47XeZKB6nfj15on30o2YJVUluNIeKYpFSXFV8
Ol5Ob17EgqZisXcsceZAfMk4XUj5kQCtNJrDhEwAIehz98+6o0oo4xFBl4gBK2+F
70MYq+4IVgI4eNBUqeOtO7hK4wzdsW/4ZejGMop/3yysS4YGs1uvFMfwcvg3Vcoo
WMNiBGuUbBb3clKAwDzAfnGE4kYCoCOfnT6U0PfTstZD0YqRi66NlvqwzfQY2smG
Cax2aikW9otMou6UPEm3PCzJ51/ulAmInOIhKk7XTjzWaXx2pO9I/b9mfwy8gL49
jsrs8oCSX2YQYCgfEhEJtPIqiquc4VVndZ2DKlWsha8NSQY1WZ4B86UMb0L7tbp+
XuvbGR+nU6G8RODWFsk3r3024ZRoQU0qzpnIrYrGPmUwnmi6me/7sEjMfvB61vcc
rK8SN2nR5mofTBX85mf/5zYLtX1+trvGNQ7k+BCUWcqKHWS65TBv9b3TkSFGq/KW
QAYGBearYGHiXR5uXSpnSD4IEGO83QkLnex3YaFg/LO7jVTagQ/dQT2SsJ+pJKdn
0cm2GI+RDsZWM8TDaBcRuv//iSSIW1MBqCmQwUvYK3e4AqWvovXjb5l0JNrs9zzn
K0QhQgTB3GW3HxOf6yU+qt7TGMhZWb6j5lglf8Ufwwe0OcgsUcXjcWEEA+BxWOUe
knNRWnJRVctyOhhTImiR6BVdPuPBkFCADYnn5nRYDXkVAhf+SnwEwKFtkGbw03dc
Rm0sMFjOYv3UDpbmYEX5uxbBd2VLfj1+R+gD/V+xGjfLQ61zqgaKKtC4r9ZYxVqc
T5qfZvhCS0D7GIa8TPbPftSm8stqFBT5RAJ8OP8uUkaEfT02zx/7zi9SOmC5xbea
kGebmRLap9CZ3EtmGEC0DSVGoQpz//jkpjHChtBPdG4rkKjjmFi9ThIDO0emm+ne
JZeL6Yq0c/JaqjBg7b8GpjEKyL/LmsSTX8Qzkh/gVRUngifm+4MwGuKKQitImvKk
l4e0kfHxHTqmkQOgFI1RFZdKXOCIv0RLYXvApi48o901hZcjfymD2lf94f2DzQXh
4dopWecgLe2IitQ0Gp75GR886e3jIPlOXxuM4R7U9TEC/ZvBitynXHvaHsHlH23p
rMzEv/4L8q2TEKPllCKjo37wiKXk/1R82ojoZjUtVSIo2TiEONGgIDGppJR9tHRQ
F+CxanUEZwvYCY/eCF6SU2x1sjtIS3mAFMM7y3bsdcY8ksNpwDeWzaOZ+LZGQvQR
jesHxRwoz1Ee5A3R06yUObOBpkzAJeGhiThRTmh5P+3p8Ngzd8HQHg2ycAactZ+N
L8w3vmif3yQhUf/CPH1PsOFOgcQ3RpU3t5waNS0dljZKxAhYRdSFLY6ol4tF8TUg
2xD1f9mlfxps/cLYfS56txg8F/kCoRX5/Uhi+7OVy0BcEl90D7wVPpgx3cQtmjzt
LQP3Lo6JNe7z70Ano1i3QqZiPVyRmUTzJtk/RsgbqLH0rlVGr24cfTuFUrDFNrH6
s76Yr52OTq5yyL/IYZjmjuXVHdvgC2wg102Vv3hkYcmTDcnjbm0Zkuu+vQtgH62v
Q2WOrJrybTeERN0BDjs1jL9gSv2j1j0R3tDfw1uCbcUag3KQ8RxU0BuWmoBn0/3X
rvkbljSqzgDpXyNieF28n0pDoN0aF6il/XgaDdu9OHR6+3DlV3HcR4ta0W/Ci5B8
Lpkj1NatAv8SZTP4zW/iDXfM3NY00osQnkyU3pK1gN2N7RU3I2HFtTkPWKFqKFrv
m6BqVzvqX/emgBJDrsTbu9ENW8SnGBQ32jyBR1jeymi8NUPIkCBYagB6At17Au2l
m5Cn2kk5GivLyulhL2z3M4wqgQvjSa5VRqdh+aCq0dWLBA/Xgppg7/mofecof3Z3
HgwfZoGRf228/XJa/OOxsg+dMH/Xz18OHAujBMybkAdaVMbzPiOtus2F/AZfkSmK
EU3yE+YznZLG8L/O+tBxpIxNNYgbkVjyM69bWfMmqqhlQWhEpoo4QRtUvPP9MUfl
PNBmxDxZN/wduCVMAgQ1Z9f757xzaWUk0LPbpro14pC0QToCfnXMTWiomAVEPG2V
yHDSQvPVgBVUrfo7Kku+yiwsYgJU6k4pcNYuYxS4Q0eu+9gfECxqKi9Pzl+w4Okc
pU4ak/kqWzUp5mV+cbehgams5Z3n1sQFVKJ8Sjf9cRTG3tWYq6jBuIQ1dfJiqd0v
yKGhuTDAMOEZOmk29BWlMikM2kf7zLWcw6s5GSOnpbyJv6uGOkXNoXvqrBF2rUVi
UVsrwFd+AP/eelwb+9rmEnJhWvins0BssBIWVGLQ1fxyjyh0pR6BcWKcrsRvXPBV
wafZIjWXl03BsvyCsvPlP20HLWIYqdDX+Vv6VVEvtUGJ519peG9rQiHbAGHoA5JF
o3j5JZee548e2W+/qaJEme17PRpGKpBwELCZJNSOQs9uB9nfBYjHkNZY9B7UeBf4
Hr7mw+VNbhoAjw1d86NJ1b6y2EIfzwKxLI9aWf+ItiQJabCwvrIzGTrZPWQ0Afbe
mbxFD9JF3Tm3Zlap1lRBKN8RUkWjFBAteQcgGvAQfMxv/5jGsX8BVOk6KF6Li/Rm
k4FWfEm7TCd0ds1NJ71WY+I9xha2/idWVJNZy7dyvmGftD+YF9QX8Xdx9q2bW9zK
W/iRKfuS7p7cABTJWA+uBdyavtzliiaRlS72sXbrtmewkhLf+i1zo5w/73zHX4RQ
QWTbg2coVSaOF2xk79+jYJEDh1fh06d7bU1uaxLv1AWMjcEpV0qabxvfYPGj7an/
QV19e5oIIomty74QHOih15G1wO0drZka1OUDYsnrzcofCHLyFr21XY2MowhoTZU4
e/YXXVhlio/8nUOJ7l5pJO+oHKVM1zqtmoPUwC0IJ5SoMhNsMtx0RCmcTy/zJIzK
pBfiX+MaRNyeHyLG//PnAI8Aeo0uv1q5XJ2ELGjhn86X6HViVQF/yMGU+/KlDhuC
3NGhqyVmjZrmxVHBVAPuuhxH8ZZVoDtoUgk19l4u3lPY1dJl53XWw7+jEdFtDKYN
cm6jhRo4ehQ6S1GXumcWADLwmvsnNczYivCBfmw1uHYKZj3D+cJpdpIFVYmU8dFF
BpxLl35vEJENODtfGggWGB6wKjPjiRnKJyP/rUjNSaDloC49ZmjF8bRbaKBiPfuN
byL7mBWbUIbQtc9ndh3w3NbA3v6uWjDEwlDjKHqR8yjJ85RCGX3713/sTWeJRKCM
XXrHTVo460JHyDLQ3+QRMzLDUIJ7U2X3i574YRuKCMOtJOI34rXQpk9Id46wjQn+
RNe4Hgn9l/u3h7Vk5ce/759JY/GUmsdqG7LCMahYYiOy6o1C+/1CHZzuKsEgTdAA
roifAqpVXUZSicvp7B5ntGyat3p39K2Y1/kE85UMOPKatlC5ernHX+t70M01BAXn
XHX87xGV8ljkroy5atXRySfHIRbQC3WsCC/pkHmXcKrEqBhTxnrqeMdO5eDxaoi5
a5+BMvE4dmZOSyxZIpPAR3n0ee/zrjp6SiRjXsbuVh8SrzBAguALILuCV1ccVMa3
yAhJLvu46sxKq6JJ9qlFHAg+bptE8ZuDBW4W2v75lts5iR4Jb1ZTki8GBgbNq3P9
73zyHYNMVr9+fJ+lG12yGpzmfM2nMZ6C4WD2QsK5QaCx2arbzxIrWRjpGZA0QYeZ
7UmY/e7ndzhj32FyAuj4StWcuddF4AhDFYV9DkU0r3oCrjjYpkWATnQJCAuW6z82
nBmhUhWdAdFfAEVKripzyLbn+9vbjXt4BCsAohFmQoybeaOKO3CVvOy+9i4jx1Fm
G25MuqIM0V2DeQGNSEkz57IUuaQEm+8JjzbRdRyNScTn5ATYvI6A4scr8fk5N1KS
09zU6X/yoPEXA5BnUl186ePDMrGKRJf33jjWWa5H1GHbfjl0RTedCTS13euYmgX0
ShQ8Rtaznn3t/GnC28NZ5K4WhL51/TfQDM5KFLrTxzlX6YPpE6MhQohPz0a/JB1l
/6UHZeBNwmo8PBZvo8rsvEPCPzbESR49Oe6EDIy3xdL7w9SIA4/ncjkmbx2glyi1
qTFvu/27xT2BBapCq3Z35r3RHzVSCI1N6QFveMYtX5ELOhABblnZZ+vfy2FsKlvL
s5B/zOG8Vht8MGesb5/nNLz2wuIwIg8X+zop1uplGdkHe4rA6d5uOCH0mYk07C2s
JYkZbxlkVnFOlBnsfbwFCXyzjjeCTHOIq7/FC8osj/DkTDreftJYjnn9CLbIf6X6
RYidvNZxgeRv3m0uCL/mjUFs4tPayaojYCGu0lG2BSAQJIrAtjKLPb1TZ8Iz95Y+
TDAmzdEr54+24tVqdM9orODjV+awphgP8jbOn+4tfii1ZQUUy4wCYNjDOaQktkRw
P9kVz7b2swo4XfcRVyK5CgHJ0IaRWo0f3nxNU5z/zWyPvy31QhpdI7XOA9yEHFsI
n4ySgZGOY2q4d1RNUdxiyGW4hE8vRfSMBAOnMVVZSCxpeQAuWi9Ql91QX9c0eDgh
SqbFuQkfkI7zzo76nb4LPF6GhJVjcugleVsqkP1X+J6XvLn/4aJPkeSkZfUYX5EZ
eMVAQyZ2jmuVACuhWsFjR14ADLWBO1sbWPbD3tZVJweRUwZ4wPNTiuMW+tFr8vsQ
BRxtiSOYZCEhhAo+Xz2oJOPsBmuMTODSwjLGW+w3Gef9CTx805aXD29DEKhZP/Yw
+kLTdOp8y652Zey7SELNlesZUqac2JkmoBUUCVYL3jyY01VUi7y120aT16orpyzl
IueOBmCA027gFRpXFlTXfI73X5CQS8nvrm/9jvL1n4YG2MtWUk0PpOZRkq3YnS+0
LM1oI9INPxaHXGO7yXTu2arPhbaIQgH8yy2D172LKR4NmPCphB6FaASKQT6MztPr
nkprRIziLdB206JuS6NN6vhqXZIACD2uKOgn9VhmrPqIZird5aMG8IwsHWBCuSDa
80clSkAWyOIdYrrC65jLlkcQlj2lhc3F/w3cV9RdoFUrrjtqbkVeKoWuikPVu11k
2m2BiTfyPoLty1wUQf34mChJdndQDvevek6AuDfF5swB2qC18yGi7RP6IjHDMpyV
YyhRuvBTUQd9hDDQdXXjLWaNkIFUgA0364HZEkceVxwxrm34VYOYY2ld115vfFlA
VMb64I0qAw4SNbd0wkVTBMmlaaR3fVYk+QO/jzpB5FLS9C4RdO9g4aKgZgB1I47j
VTBLwZ7BCuHMTiOFsI2riD+ffsJmhRUZxOFqIvjB7eV9P5b6+dPwS6/EXpD4vuEt
rX3juNZ/zaKsA0PzD6CuRw+8PYyLGaZy/+no9AJ91s8LV0b7g7Twq74h/7/55O11
6V/xojPCDFmSrUVOjWQRm6bS4T7hCf1MNZaaHW+VHlIrGl+Sr+JSpGPCS1qqyYtc
AR+pmnZDT7h3IGZS7bJreVQiwNrcjTCok/FHzXzg4b3W+hbl4w2vf2IBl0zcCWYe
f0FcH/q8nhNrhbNz4y95nCgMnr7v+f+8hSjLQ0TVOX1zHCb7oYXdl6FUh4MAqhq7
sGfwcC2VANZ0rrQ1yYKcTobIloJHlC6EFSbBNBiTxlShu18loudosad4tRKtRXLT
nxQLatz0IM87/RgPT8xgx3GhVl8PUi06Gl3tFOknxt/CjGSdYtBekZ2V2w1O2t1x
vNkwB984D/yUGwncxsmCSYLDw+GgmKwBwmIVje1JP6n26ekzhA+nk0Z9YNSejBPF
uQ0q0HcojTf9VtLfEkgcEdM92fQuF1+1lpygOVBiun3ntRIXYw++DaGPAWYwYrI7
iPyES/+xRCnKXXTthjpEysEBssp2DV7bATAD1XIihWAcN2TwWd5d9liYjpKmoV18
xUtVZ292AY4F64MMb/bFVdEAeL11UyQoBIhByueLBS6ENB9BmXq7f9wdxtBm+M2s
OjIvG4j71QhKJDPfaW++HCvD7QMwrfYRVuooOdYTlynN/Z0+7pKQfVxEqL20acxF
TOLbR4Ygo6AONeR1iNidj7T75+8wuxrYVU85Oe/GQ1iSahUAjv6IwUKjvrVyCDnM
2mey3RZ1fSKlRWQ4SCt91Z8lpMQJ5Bumwd8QgK0YWnDq8uf74cBcusLsTukF5hXP
oyHzNfib6TKA257oqDkEpPsXR7W8LglrBBPk36blxo34P6PuSk4TBOLR3XUPjQps
OlfKQc3uFpWof8C0xZVlltx8P0TOPArMu9xNzeWk0anGfGAywu1Jzxxqa3UgOofv
7B74TMPAd7tEdVBHlyrpuKY87/Nt0tAwZZlxtlY/TQqCm17h3jyxVW0t6U4+tMeH
n/pLIOREN7NCfmq2H9e6N1Lt2VNjOWzI0Rufv5AmPaIMPI9p0RF36o/rSM7/A5Dq
7CJ8WxlwXgycX/DJ8H6/wkUmkvJvvlWhs+qMn2b0bNuRQ8Ju1n9BNeoni8j/jm9X
+aiBStJo/vUhN+kHZutkpevm0m9SZue3l71roVvFVQzA9ke6FB87O3Fqf9QkXK4b
gNoxQFA4IUPD5QgdLP8KHiDBQXO+JhPLwq7eRQ1VUm1C4J6FN3PdaxdjrMq1M15k
nyywX0VBqF3FyKAsKTlN1T4UA8XQpHibPNtIlaOPl9gvSBRxXoofEc4qh2eksVfQ
SW9PK2+n2OyMXlPtSt6fTe2Xmh5c9DWMLno401QVvnBvKbPmdwoDGEoOa7RHgVzj
3eBf14CbyWO6yMuz+tDm891xylygAiqw5rLe4GYyVwvx8kNY+GmVDUvnvC/Ic0Wn
mboRGIzmlrP1yhmNnvpocN/jY+a20GYWJnbIIE8ASIiuDiMKaIfnBTmE0lUp9t6U
bk7M9hTZBl8sJfOEM8Im6ZNZAJ02EFMglu0NHTYNHUwMSEloYf1GbyVfop7ANGYw
HfQRt44pN0XFu4TWhfpfA0Dg+lzMEfRhqAPwM1hb6TKJmw+Wg1kWMttdPumxa6PS
W1nF3PeWZZ70L+iNOEa5LUyodz+qsq+1+Y77iM/uGCoceqVJZcxs1r0qz4bNPMGT
UTPGYVt/3pXwD/IBU2001hJwyRZ1jV/hPZWkiWLdtqvqUGaprHARbHX8YZGsD4Kf
yzFN08b3ifRHbIfv4iIcymQdafz+tTXvQRrKuUqtvHb3wZQU8nPssqdp1z4IiaJd
xjnURXHrWKvk3edEvwuxXBBmzUC302QUMKZ4QWdpg1U5Cbo525ZGQlXJKwGexuJU
IFwH/eHh7uhiFOXc1PWpsCrUQUwJi+TipIM4t0Q16a/pW9qpfqNShLraKiHN94hT
Hh9E5ObWHGwKcPTQuX2IzpKy3cYp9dj0BWSQ1jtbXQB8sfXGwQJPe+jMtc1v4b2L
zOH6abCBgC6kBy3BAvl7DU81AMPO553TCjdev97J4huqCdBdktKA7O1tA53tabAx
byn+nJUiJrSNj+9PUqlq8alfhf+rkQUyWdmvHCEsw50Ab6u1CIYM65nhgUvg8ds7
XTjRfUu5t9huIek/r1uw5nMZagpRTqJuJc//haIWsACnfsvUgq1xmsS1J6nMP/kL
pg/JTr5pN9MoFLCKjIRC9uZp2L4PssvhjmcYPQ6Zx5smCPTvEagDzwTvHVTULBXl
2u7VrkVUFc23OwqfbGyccwm/d0KqiIt9E7U2Pkh8hSXITwM7px1MzqNOm/A+Nnoa
4hbVYjm83fJwwZ9xAgcMTOHnEIgqttuWBKjCsV5YJlJ3JOR/ky+prSEThBn/sM4h
n4A8XP4t2tA5Ohd73ygwnlGu61c4b2UNBdt6lI4U6Yz71jHtwDJwIMnPLifM1BfN
dgj3sYs9aL5lqhPrsiIHnTW+n8PvyTrH9HeHr/MtIjVWC/y0DjNQCfCnen2smvSA
Nb/4EPej/tK1zqhkRQdN0Jo/kZAyexI5eKIE7CbMARe10s7LsoMzyUn5YnFR2T4M
k0DK6ymEvWrCsmLbMYd9Dzap5+qvZ3PMNlo+TXik4xQSDLOfdPfIGxO7BhqCjrdY
pvRgYrOxL7oqHRK4SFWhdg2B+CJmJAhtg5PSSJBYXDU+JCzGbPeODvk06r32Kzmh
PaX8zMkK0ZbAbfoqAi8+cqo5DolkmmzqGmkxa1yRmHhCaJT2ewsWcxIcLNngQc+w
TUNri/IMt5F6WkI4p9A/hUJO7w5cPNZ/qnmjcemURNThoMhTYeXmpsV00M5ok4t/
fNyipHEdt/VsyiOP7UZmXFsJm7SkE/Kxx26hk8TGyuwuN3NwuEtsURz1CgHMYfDW
xeMzamIxeM3TMWIJS6Mz/u//kYE2INwoyxtB6GyvcJMC962cKXHP5uwvoNlO61CR
42CLflJVaSquv+LV7Okuv9BRz7PYEuvEppA+K+w/G+P4Lr9I2/PBnVOyGpqW6IPP
wErIhAdzm9ihrs0qMamv7HUnVzR6LspN6dUgDhiPCWwqfdPLO115FyqClGCV6Krd
b+J45s3EvQzwoLkgqPSPRwraSsjOiKZNU+K8OWmU+FY63HsnRHt8gwjyW5TA7xL+
wtL7i1z2ProUCkBSkz+E0OYJtuE4twtUJrD6GXEZmpSTPQ/jUBGkV6T59X3bU891
wAVuC9PnKR+5RkdvcdGdQcS+LMFhE8pSgo+ajJXxjM0TkM4Mxq8Iz75AI3tbyIwX
ycCcVqRvJYwmzQ9NCIiRBtxwtINVz/HUb6Grm6v/kAN7cLwpB+ZBPYjKZ2yvOIK3
f7q97AzBLAkJjcFTWW4+SoAvVN4uRBnqzZ/iOD6IhD+Q7xN8u4VjA68TguurH1Tg
/f8Jv3QfzxTYK9a9qzQcYVn5c+DeooPlbNzEPSJpz0U5b92YqcHAhU0sH12M4TJF
sj4lS0+WuMzCvSu/vI6PseUH/W30FYAzm7SG0lzwlC4jS7AGN6VykKhOFxJnNTls
018aPEbVaGlTCDNMvpVSesEkzG1vLBy1fRSFTy+0f68ghE+ismfCoUDGVGiMe8cX
cZcYs4rP10LSziKnk4if4gS1225SskqT1IqCWqMnTh4iQEEPU2xPbN7fJd9SjOa7
W5cLi49zH1liYGWBB6VwzQDMPmCYlaIaRFzUmOQl+DSoUYjCCTU4XjQjf/Tp41HI
+i5rZByBmazhXc8rbzRdfJ25+p9YOLMHu2YTS1ajZRA1WJkCMmTgr/feWMUn6APR
gxfOd7DVU/9sIt8zlHj+xoEhrm0prU+ANoyZySwnEWMpmHRV+k1znY51IRsxkKP2
lPws4z1PaeZwCnTmMaGnUfgpc+O48QTgYpuSE9/FF6c0ujG0jUnckZc82PkuMp8h
lGirpXGckhzRJP9FSrzEfiwlInlSJpyoYwuf8r8Bsm33R3eBns7T8UfzdIdzAk5x
eGmFhggLtcI+zObB/iGpQuOzOFhT1J1XPppWxSUbR7P2xrDOwgZKIkSMkDrMELIh
kTSmlg/wyLXqsB2gLBq1jAVdhq+PM/QRV6sgXzpmh5yhMgB6b8+XME9+vcQ+JKuP
cN06aZRyjqo0E5hYuQYTHjLsnntw8Xywb1e3UiTIhv3PzyRmtsweQE8IOHZJRURr
kEoXxPBFQbPC4xkc+EbC7XvRWiXZWUe+/6Dhq1wiFG1zIJ4k9fUr2EzqhqTJxXl2
WJZNGU9zjFzpMLBVcS+xErOfN0rwCILuFbieGiU1yvtTH8wV/Vc7B9cWOnfAVuwZ
CzTpWO4znNRL8j4CJVucwjCO7s5bJ41KIYN/21srZQvn8HPgU3igLMr+QyzAJy4O
O6tZ8iThmwEd0gv2xtGxVb9Lg5t8LwijAzYGcIMHkZRBqrcgT+E5m64+eUABSNwf
GhRxFY4p0mlJIRIVQQeqcFfnRp5zOpN5FpnB6HxGTgMzvsDcjkOCGIVPDQcxacnk
5RSUIBGwyMVWHrlSvfgtFJWqt992CbQWESEHWhqQDCQKpWVjVVJolZVDPSdg3H+a
FI3MGtNO6reo3X9RZbTrVfkAkLEr84Y9mWUiNKJrJLOenUPstCeVQiyNQwiDRr2+
WAtNCpmdn8ZebWfl1bAQdGriXbAVOBfGwcd1GKssyNI5ZxD2gF3u/l7y3wek+pez
d/6rpZ89kJvNN88Je6oxf/28b1YbeC4BAXCY0tkJqzE6PieuuDtVh4Fw/ag/3iKo
ENBlXuNINzdbMi8gdgBFnFaEmKiynnCDpkeQQunjnsc0E/Gw5jaYmhW3DtSPdyLy
5P/fGsSReikCEyxJebZiRJ+2cMNey5qpy7FGcPEA+be6JCDpS6Vmyg4sqTtJps2s
brDuHy4/uW74Ns1K7iX6w9f7SLS7RGa3Q2a70a1sk8FXL1Tn/3sHtxjU7PuKE2gS
eOz9WRvXXvsPsmC5rhXb54Q9bnpvdj7/pJ561sU8KkKRufYaHNYXwXhyG37lNJv4
UQguS9L6FgIa0/KSIg9EETjuDI+d0F1KMgVoPaycazIgfFOk7EpQjTcNSQHfN0YW
3aoA7fMv8FfqBPzc2r3GlZZvV5R6Z2RsQedMOmScLLnT4wpFUpLsg8NCkKOJ9iYE
erAobBp4+RaAjN6iWfzzrZAxN7//KFv1Xt42EbS3LQCaa0JK+Qi90RMclnI6XZ5m
xtzwlFF7xEmmhVMWBSb62p6jAzw++FtA0n9jAc+qj8RctjYGN3Fp4girdsC+sTtp
8/hRVbZRmqxz7dSQBeQr3X8sOBTr8kXsjxvIcnk8tCffLY7mmWS3PHQ2aDAkL4S+
UL8CoShz1ZEmH73RQTMUqwjoOZiw55JCX+NSvzTu3M+Gs+t/nJDWt2xHOVDdDd5l
iBFTyxEd+P33VZ6Lzl3XCuJ+xzZxKGCAqIImKEaX4ioajpz+sjdjSwG+lh4pDDao
FqUWgfJtysSeCg3WBI0ffrtLk02QkzxZ5iL4xgtGU2AYSlgIIVnmW0rOYlGApt8Q
AadXCcBn2JLlfw0FIkJIDA3OMW8H27/ZhULqYMXaqNdvgYNUKRSXYk0rZwPbP/vf
TtuFdZO4L0uYJMWU89JSk5HmPrmpnRsgpRJw+3FWl+0N+MMcFwORwQYfihN7VmIR
SIrsKHUK98BgdGL1kAi5JJiXPmmVtDRKzQcQtYrNyK04kWGTHotBqRPn78QkuMCk
PaOFsX7qcu926ZQEh2o8GCoy4v1kHZaJMWVH8Vc95yjIfKraOZ9GUvEVOjbLq43s
rOnTCPzBIks+tjmx1TP0cvNEPDZy3KYXwo9bjOq+RrNPSMFdpoUO5vc4cb8GMd0K
z64eu6PjdmYWDuTpgn50rGQnKt6SKLY0b09vQveX1gBgOdWzUS1vx32GXHPyTDps
3h9wWKeJtLTV4ZG7Zxcpil8j6lginiksrcs0Hq1bNVQ4cIn6LIok1y7xDWFdH1Ww
fo9yLHlE0DEFlv0FF0GIMFRGkTV0cQQsjh4bm7wg0/Viv3q1uJiaIS+sAbelgOKe
QrKMbaRCkrsY9F/PE3OWItuJ62ZBwYJ3oZTX4oQ7HKxijuvX5QPsB/v3wyYnZj7O
fMkLEY/MauE/hKnH8tVGlE8hvyrwOef5Jsrh6nMS8mN/c09PGqhHcQtX1C6rClu3
jCzufIWH3u+sR7wERm6lNmW/YEn+ngM6yglWfSVltesA0QDyiPQTy66wvDSZswLr
KX9vRt+Z3K4g/sGuj8Us2tW+ciiXLtCTQrTinRA+6MM2wS+xyASiY5writj+DgWp
1QQ7VWx6+XifmQm4L3aCbRa3HSAwfRgpw6WLdrEPVcNkjUlrtjD0jCJyU4wqEQxi
QEQ6YBndYoK2bGySrxGJib2crhMj2g1SOR3Y5Zp+kI/dQ5pBgqDTkbwawLwqg7sI
5EqvksbqG64IC2OQ8Ujk2UtJxAWt3a70xkA7lDMMSIiFbQs3d07j1LaWM+AzfGH9
H9Sv3hpOoFReEM9hFPCkrIqh+3q680MqhlFHuiTr2jAJ5Bc99FO7+PtrPiejnkdP
bf6ah0kPneP0BZ8wV86ZkJ7De/xnqoZJjwT4Ov38HQTGt0Kfy3G4UTCFJXVhUbKw
QZFBIs0ydVEdEHhV7hVsM9DIS27Zd0ei+YD2XCIIQQ9WrCzHdTzVP/gVEa7Ucx2T
Lxot4f88avtCEUUJKjv8MhHh2gI3gU8FxnJV64MuMI4NEGGpIGAvK4phR+Ozk0yr
cCxl1EA2bpgRPHqlGWU9Xs6aeiRijtEETARWcrzmEIROeKQn/DLe6c4vHAe2gL6q
zKjKi+2yy3LaCOxCBP21QUUGWLe+r33Xu+JAWjdFBt9IbkrvEy9w5olnE7GH3yaH
wm9etMWBNWkZaz44E2fKuXNcQJkR8SI2mZAvEiaFeueXOpJEvadp5ux4InQYdnrE
cdHXERkJn7jNBDIBt/36wD9uk36Zz5Yys1uaGdzjXCOC3G8KWYz8qvtL1E1+GUrj
sm7wrvs/8EBKHv0XUIe3ri5s82M5YB39wbwfm3t/WrenDgVMcimqU7hVZEog/sYN
NZ7KGTapiByA0CUlbCu4/IF9GbcTEsyNFgGQn5CJX2oZ5m4YeUJsyXb9/LgOgWhh
Qe+QNribmc+l7xM14YPi2Bf34Xq3A8JxK795CMiaz+CVO/GOoP5jo2nouR/aqNn8
hKTiz7bgkM9ByMEySze7PherxxXoTqhCe+wC4oLsIIU/RDQjCL8hqfjn9htoqZaM
mjAa8vH90l65l3/L3P0hk5poXhVkW+Nb8c9UMkSDRtnfVxaTghlIdpLxbwbrApZc
JQwQFuQdwsNQ1kZqk9QzgCcw4NWvtL82Nn0sFgRpQ8oVguzFvBqfjq53ACBBiA8u
yvxknxMG8MnbjzxA0SAraN3pizYPDdNDvkcP6rEpVZl61k7Qh+2cMhfyYepyoIC1
5hBfmIBpsBd3QpcA6fJiMu69wFQOy2wB71/uWjCF9+p2LRuwXKSK9L2AdE4p+LXI
SNP5kk+b+5fhOd4VJuI5a8vajWxrZRvNTLbdd4WgT3SXCDLw9qUjAjLsYSjdVHCA
GdgnsngdKyXJXnmJA4tT8wBGHy2qNzf7Mm6LEpv5eohFolcHQJDYAXOBmi6BjsMb
tyq3esVFHA3WwUqGZs+ZqtA23ggUGxSthK/hZJBpaZxYfyk6ajD2nPoOX7W9ExQG
oEk3SjKS2Ez8PlRpqvsdLCpy6ZuxUCzHImUipbyeWVbhFqjYR5guJEjMXYBmEaEx
yVGHY3/fsdCdisUn6ViiB8BxmXbr1sjchVRTxAXpQ2/1EyMll+tYf7wIDNls6TwJ
6o6oOg+PKT6f3O1NqBNeXqaxmk7vrw7Z1x+F8PEj1Dcgq6ZbVc+sJvjzBEdL4iHL
gaToHppbPyooOPwW925dSiR/gNr9vFjd/trneQ2NfQsf3sfeJcYnjYSX2vMNXPJE
zFV6PTGIbI/M0GNyoMGCwM7Wq6c86cC47E+O1liuwsUsG8/Wv8yvuk8vyJYoy9DM
kaANkn1B9pzq88+VAbHfnxvewOIiLsNzZeNYCETbosgYdwH5FAKxVjT9t3rEEUbu
YJ0ywcfcgSWuT6DbrPAJkKc29FcOqexqmm9ucWWCFQbQe9LOsLiiy1HxJseCvVOF
8n/wTaXfv9xwZz49/XtuahJLtJmVC4ZlUJNTQlzJmJ6ULaNaW2ybe1xP1F6VMWL/
gwh2h3wXStMTv+HLcnaVFFpX8g+UiTz4FlKM8haDWRdM+hL0cNVnpJzHYopQWq/W
l+mdLhclA7BDbdUzSwL2ovWfHuWIEkerAefCSVsANl/DeBzuosZk7BlY1qxH6139
xnNGX1dYEqKm69EURUnA8/aMbbKPbtrsJvgp5505MVwSCCB8uXIPX/LQXra427Vk
5tsX5ygR605IdHaQ+u1UZ0eTPPW5GelVKZ5pRbl+fJ1ErTy7Pn9nH1Rc3dGIcHMv
fHtGnQOulF8AmKfs2mmCW01f8K31YlEQgVPc3AOXzlrcIf/vYAj2pLVUB+WT93WC
MozGOqPVf8sPFiCrksFBXM/bpFtlDqhHd2PzheH7nwNMaZkGzN5mUuEN9zoCztS8
KpgNvWMOaHS4yTBh87MmHiKPfkdF9/rrdG80u6mYgBxXyIxInSG6V17JCvRfU4LI
oqqr63AmY19axMkpxqY89qcZUn+WG/onfHmk7Lc9QcYHYNF0Kxjzyv6n9165LGQD
/9WjpMjomNXz1lL85NeCdb6irQpqQKEogeaztklkIMcHuwloff8GjfMS1mvHbPOe
qOuxpqjHyRnzlgaAqm58boAUEqSId0G4+/2wbERdE/rumBsn8eiDGX6XNtyXCdLl
6zRtiMrJAL003eKwomGp/RHM8QPN43Qx8qNQqRdxuwp88egXKZCr4F4dlQ5sB9E0
X0RA4Jv8Se/jzXBVj4XyzG5+B6XobKFo8L97xoYU0XSuduPdRpJ83gvLJ7FPLnh7
otAtFBVVYLlCiWRXyqcLUsgPKUyGmH8lgAkxNMEYnETmLuCZU7crFv62z1RGY5Z3
DD5IobDIbdwvTSLUpstpKpQa59Ip4Fv/1o1iZdVfdnjAdT/9rsBXHnyWm9xn1DHD
YGYKTcsIktehR6aZPFkyLxq7MVZAOtt2/yAQch9uvShBwUxtRRpAAyPNhk500HmN
id/3HrTxtKwPu+bsTHjhdEv9yHY+Wc4nE8czaG7C9vXbobzkN3oO3dWQ50jXcZWN
CO/eujpMggQGbxH8UUgQKWc8U28jdTLRpO9Eh21PRhl20T81nFUbomMVZW5gLY7U
L9h6Zej9E3bM3QowHnU9ps9vdPHWHtXXNGPyE5Wt3P6e4qatYZPcdi85SZ6o8Ecf
7hs5wuQctLu9uvSnH/cUtPMfTFzEFTv20byt4ok4/BRpo0Zc20+FeM5HJdLJKjzt
9De25Xq6yVA+8YR890G51zUuLQmE2eYVTF3DdpmUPAhayuddy7tnyeuFNjbPWVe3
eOmAJyShMUSUqCeckwcQIe8JH/kKNYpUqHhr1UZXqE6T4izy9P4/0kKVfulc9M/+
qNAG1J9LFCECbJEwG0A1457Baj5ysZ7hXhJ+z3TWD0r7T3rf6DihgGqPwSnHUXPO
tZD3Tuplaqh0yjiLackuseoP9wm0Vmn/TBIPPrNWfsFZsDv1qm5+K2E9QwbxQmxg
BDqexl4s1C1kh3bGNtJveu0Scdw8vK8Q7+J0K91D9JKbr63Kandc+0mcu16cZ/H2
BLYqE7RuczGSDuxDG0Y9G3Ar2I6sEmzCqwNzkH9q8IHh2yrfMYn+eqZV6/La5u9s
5CfpA8QHqhtzxjuN5rT8wwr5BbO8NI3r1DzhDhGCdDjH2dkRirQ76QJt6SvdDJ7j
9R0rfVxKYU7cGm2feouLF4mDpdYMvBXvaY5jSxIMXZx+b5YOYK0hNAkET+ToWFhU
yIKe2FQzylIkyhVSUtI/31awWZDi9/yZ4Vt56/bQwuG0PwhIdc2xma/ge+Gb6IlB
XYN04/IAKZRkt8Jmmrw2nyGYzoIx5Xp14DE6cJK+zKHMZ89aDl/nepdyxp218aPo
CcvPp1y3cIZXFRTw3plLAkf2xnJRwuPPV27KBcbqE2eSMZTBu+L2u9izeCLh0zT5
880aqr0tFejJdzIyTI+/PCuCjh8iXWtXy9650C6U86uN/UhGrXc0EQesxwipZ9Ro
I9Fkn0oT7qKkb2KtW6tEJTvhYx6GWNf3JJpq8Avhp7apfVGMzyOR1YX5DAqDwcyY
Whc1G5aKcGZ8MS7FIi8pCHK7TYC8mjSl1oSAiLBXuf9/ix+qOoxYU99YmxeHTEyc
41fhW2D3hbtB2vNMuOlUW5iQvnwj+Nw8yPckqKOg8MmCogMd9OjfYL1Asybyg2qV
PpPlElsz890eURj8JPihNBwjsmq4+8JxEJDDI4LwiK7NuiI/P+c/PhfiRkl3cmeT
p53QS02TPbmrS7GP2bnRT4nQlN6vlRp6MRTSkE6gPm+qq2P5fGph/mYWgOoybcpc
Y69mktqKmvzQm0sEUGuJF6WZQPQeY39gGsQRbheAtTDd8G5skUeSnLegY4ObS0rY
e1C0/vCjhrfDEpMFDapqolxS0yCAL/ScMZfBgm7WZ5UUKeVsvFnpAmqEMJvtVpNd
tBapRklG1NxU9tLzz/M2B2S67Aajb6DVCnjvEVGOxNRBBDv4HSqZx+5TJGtqsV3P
8sDxoi3IxOlni/crdImB50nAoqUWdwmIE8S3xlpTg1pvF4VO056Ckk7ogfD10aZG
yvgF6mY5k42IfLZuSr7KlQPbG0cdWgGUo214dxGO6egMog3V/pKTd7VbezyDVM8B
z2zJ3QSGl2yABARAZagOO1/f/sU2uLMdslomFlEvf6b7QxZbkG0xIU/8eSZmYVU0
k29Tk7JM/GI97qLLGye9oQrehGZLzHpv6DFalcjIle/OK5fsMTb4VDg5jkx5kqxE
N8GQtzxuyloVA+7fURXrIywp+i9QDgkBLw5PSRt47e8fwbC9TWfnKZCJVHbJATvq
XHbGzMnbYAdpppQktqv4mvsCymF9+7SRwacPdzw/lK5SZfCWoz+fF18kNQRN60bP
jEAm4gD4RB2NWBYkNrpp7umQlJaItHAhJZLwwBksK9ZYHQrNHo79eCWG9YQzEXBx
IacMJh8uKhQ+O5xkpzg2gPNstKme4Uy8ZeIW7Mdj5L51goZ/zIJQDc+YMKoGCH2t
WXFLiwV9jyTBGuE1lpmqwMFyI+m+zPjOVWr13gnM2nfQG6Gxxe6+zMCg7cRyu/LE
e1rlYHUE05SF+L8y53yGO+t1gT6JhmUFM1fvWb/4silyCjB81GhWdF+g+3+DkLUW
UslHe7F/BrKyyLxIMt/hpL8o6uo2vqsAJu1l1YZbKW1cwmYlHbw0SA/yvTXdpU9P
e4vJkageJPdLbxClzPTjBKTXpbAKUuTyZk1hYe8wPS5n0edDi+tCYUPu9wDdS99F
b/ndWaAqk/Ez44DQvenbuvFrjlWYaJgld/nfdq4v+NfEHFCruvGXdZO6C+8Ys/23
4/QnOb1T1grNYGuKrNf7wy+pVqKSD8/wqRV6sLOQEly+qXJmuWAtZdz0C38YO1O3
jYTxvstkFCgXoX1mhYmTUxz41SIOrL8Zn7Z7vza0da8GZRlHvg4z0qM2I/bJE9mq
pfdfGD37sRQYeExWOCeQ2wFL+qmQk6Qd0uyXAZtCv3yCWPyO2+JvCJVi+vV9BK2T
BScsSwRY3/b0xkSlj8JDCQCecWB/ZyrHh3A+ExxiG1gvRojnUArB/7Lg8uOUHJLc
5uqwd+tsulQMtkPtY3aii1q50f95KTbgGuU1UgmUZBxlNtuMn6DY2HzAg09Uml2u
otRwoU+F23ZVr71OkiECrlmiOrnbHiLtCpoyiWhpYTK9mjrITWOG12NNpKoKX4Kw
Oj9tY9nKyUyildVIabW3/JxCHXsCf1orC9k07qtWYT4FT8bUnrwiRtRlwhhdtFLp
7wtw/Wp+LDHvRs2rnZYIB10UNW9ivOAE+5W07bxlINr4+4BI5JSnJQB24Cde0tjT
x20LY6Z0Nq0gEoOoKBk6I1EGuBUMAnKYcfd8SWoIEH9FFBg4E6vSgkyOa6K48fH/
QR7BWr7DXWh0X9RdwNbioCpyfeePal+f/0bYCZDeFz/AXjMUXaIhK4k7GnCR2BBd
Kc8Bx8MgA/SO8FL/ApDgGO5p+pZkBBvMdTW8saS52VYOy7ywSMxq3KCVH9gUfjqD
9lYK4Qxjor6q8Ghdmqj1u4q5dwkOxrw0B/xgawrCE+vzmgVxZ4290uOEz72c9Q5d
eoxCATGfpaUmATA6a2WphbebcAaYWbGac8CtYycQwrrYSVE2pe1rBrQT9KBPno+e
NZCI7Uf1IhCB6hP5zBDOV2mI62ej7o3yqahrcgBCemz66Gw4Asz2VHxeYrQ3J36p
uxUFBh0bQBDR1+NnisYsRUMatEiiLwFnSJ0lLXZwjO/nSBwNmeX3k84BSjoYKmME
uUObd31R+8BBgAHP1bi8V4AUkLIGr0e7aDX+FYiV60lhcx4KTXZcIclU3E540GXy
6+kTE3I2NlQpN0qUci6YEdFYRD4bs0ATSuPQg9dAE7vPUUK0mQvGzHqREr1vv2Xt
nQaAwEwxG0GI6uE8GEEYGryrjc30JmXgf1nPtDhse9GZwQL5d1AMQR0W7V3jzU96
EVBwfbfIbcUATzGPfu/F4djq3rYXKvBAtDxOSvTB9SJ+m1vWBNDWuhhtYNkFro4B
dQmM1Pcp9wayA5YSFmeGT2zSVIabioNKIL25HZLfnZ2f1Jp90zeG9NvDtcLhFO6e
rcwd0RfpgvyxLud2AnixEVCjXFwLYQ/GDxjffazKttZ21NWtuXJCAW3uRRIdYycj
jHFkNs8X67S8ojJwk6dE8sy146o1ZT+Te1gb24fJT0gUqO8gHfcQEOfaK8NJkuR5
41CLfdNegH/F7ykTqYoMyvQQFWYc/GyVVJ/LPDFIAaQPEtrZuyzESSLsgCwHptZk
g6vhqCoQ8ezEtInTpbNUYRxagur2fhvIQSR5fDh4xmn/ArHTxEV++TrEATYzlhA7
ynYjiQiBd08Cg8HJ+Q50pOyJc+efyIp8xw0IqeYM3JkNc0c0IK2grnI0rAP9DCDK
Os830512zU7WTAvQGMebYbPx7/Sm5SrKeKcBI6KxQ0hxRCK8N8iTWs8s1tl4ViIB
3dssy+lMcv5HlmSQqDhPu2cYp+XSacNOa+nrrzWc2bEIj2DblFgZ7Ihmi9Y1/oJq
ehCwOnpE70iDcOxwJsSiuRQqWehw9d1fZYHcUXp/cN520kNQ5kDGP/BkuLT69U4K
MKX84kLL1zGcRgIjWcxWYzLPZuE8nr3qu5v5trsMaaWD1N/JzjVuJmTmLtDtGZC7
xr5he+XMkKNAsUFyen8ZBfCpsDwzUV5pWpD7wdKtRF1bQH8IXZsSkwwg0cIjjtyW
NZB1KlDwq59e3CvalucAaCz+lWKrXIK2/uiozDNg0ZRUucG/qDsEFPFCvKI66QbI
koSnJO0/uqxkQs82gsPxYst/8rzCUzABAjNk8E4NmADnbtKgA8B1DLbLDwERx3m+
nDANkpzihC2h/URTNA6doKW+Bg4OEP3NxDb3a0N9PUjXoD4Sc1zWmSSfr3cv6O1P
9ladnTz4KOMHrmyj1d8mhF1++1lQ3gQtL/RKdO8A/OYP+Sgwanx56SGE+yLggB8n
raA7CPB4cuWjAybSH1gfpHenEds4/RD7L74FEOeNldkN89nvG54nVDvdX81Z6ddu
yIjQRPs5ucNjsVko8dJ6AHfkAZRaPRPDqabe6K3MK94EAO2npbutPulwD72UK1iJ
U2wsoaaw1ZOPs0ilCa36jT25AZ6YXS0yO78yM7K52m5avkig9GKlwhU8s6t1QF0H
ml2ibp+AmEEGRACZzaDMmQ==
`pragma protect end_protected
