// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 14:01:30 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
MqBuayxE2r8oJvd7FxShCQNJIoig9ZRQkkS3D+dNbGDk8AMan/RcCdfXpvZHRQy8
zLxysqQTOgCkvkPT2CZkX5mV1l38SLT0Nv69ny4h/O4IpbP5Wy1EPST7fgZSLLuj
5bv3iuxFhljkQDrAN1vDw3of4z6IjJwSaKuTYZSDLDM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3280)
C0MqkY6AHkHrmK9+n6DcUQb8zBlpsVYtMaz0ylAPvlRb5l5ydQDuig78UYqRbolM
jviNmvX2jAVzx0S9+4i+4jv4N6fn+4KLQry9bRVrfDXCRKHPVP6T8jjxueY/GLPW
lut4XWecddL0i5tyseuQEV7SdzpdND1h2ebzR2DS3rUMcaEM2v+hRQQ4P8MgQQE2
XNvDIfBYA+8uxYkeGhGpR/2OWnyp4sCwkqvwb7Dr/Orhk8p6uQ5+VbABm/u4Bas/
3k1UUiaVI12tlC6LQVq/b/RaVPGVvqTHvaW0/wvvBcaAFL+cumreNSX9k+kkE+xE
6ZUKPChbhIFGtIgjpnXYtvnB5XwClK0xVFswAcYrmg9ucOmE1CwOxca8kDoj+Jl1
SvAXMx8d/Q0QxDSHWdD99UymD9bwM7U3lIWy/hJaaJGRnhkweCkbijLGWxlaxsYx
qcVRUglwc6J5QVJRq+flTNafKkE2FIct133DzjRRnihXKI/UdAsPcz1H5mU4C6ep
iiWTdV1P76bBy3Xq/YE5Qg0BnTjdsGCIHCQ6HFOK2CNFjs/P5kwXtS9PLuWd7K5N
Q4hh49X1lA5Zpc2bPtl9XNrsaheCuah8U3qxlCuBi+mFfNzIfMiXgO4EOVOYbbvv
6NJI82fY6t4wxLi5LWCmtetfS/F7ZckvjOPKqW3D9DM2xP7GstmKX2VjZl7U0f83
jfwxkTlAZZUxS+XgJnmt243Hzl9Rjp5s/gnBrFlWIiZ373LqTsSf35S45c13mgyU
X7kEn89NgCVFzR+WTOdf8Up5XgXU/N64YyTuTESLzgzze4CljZ/i75KJRm4DXv/5
dll1S39onpYUqTy1l/BVw59jJw+9z4x4H512lpEMGZ3J+Cu/upnQ3xB1pXq2wJYE
bh0go3kqQwz3T0YeCEgsWtUG6WAPToNAEkI5Db6YHD7jb+GlnJc7vM6O36Abi5ST
DQxYtobyykYvSNN59Yfy8tTPbByuvAfT04sS2SA0FcAowU5GCpZv1dqZD1V04eGd
zp9HGgfdAuKfRE/7vtcZfZSXHBAasPjB3TYyDdQAiyo7BEwtF4rdpDJdAtPA+IH9
eO28n9TpqPOvCg7v2KDkRza8CGY/a6a+uW8EPqGvVbGp665me5A4cqC9amB3d+4e
wko7CQAER4s35fSAP1qoPR1rzCaa324wuXGyH65SGLKVE7m4rrXUr4+Ntz1LPF74
P3ySnhaN1HSErcSfZznYPz+HWu/S79d83mEPhjnOaDael2++UPbSy+I7JQPeOvRs
2b+/44Hxa7WJAluEdEo4Dsg5YZRAG9bSa7wm7DiQXcdGiEfNigrQy+GjNctC/LZI
5NPXaodDR/qh16WyRc/Mzv1C9bNvzf8LbB4RwL9vXNwPmau94eheLbLoRMDfu34h
S/8dPfC3tYUTEFDzOm1z7J5/imvoHxuEoKy6DrBBwAXfp9tSbpGjYm6EUtSbqg7r
3ocVPYhEGFefJbSp8Ze5tF9BaZagpS/cMhnObJxfhg8IYa6yIikwDCTpJqBCo7Lt
dCCBGezW0e61c0Hvoi9f+TJP+63GPDcI+tpHl+9Bdyo1yHvcJ2g+5KZZ4soYCsqf
a2oA0ksE7msC50SSfLPYrMh+z+ny8Fp06GYiU9bmO967KjNKihDvMWGY8MKrTLYW
ZrsEXiW2KHscU+JNX6pkS7r6/AnC4cB/oxS2ZkMVT6bFPSICgpjQ7c/GcHxPdZ9w
qqfnPjZ5YDQEl31HKC9Q3W2yY39U5N4B1vPR7EX9s4JzQbWrwKy+1dG5fLEGqXYQ
FuLWgrMR8jomJ/W+Mqnvgyei7bCDSiqSx3NfYozXn9Ih2FZw+Z6J5V1liJQWudUd
XXztZPIi9j061j3NAOncwMQoYV2Q5mIPkqW7IphHV2V01aZcSHJvgqXWd1XOJ/eh
mCXH5NcLVfz/IpFeyzMe6YAQsBff82Mj1gPXOfZ0gI6SH9M764kyVG8QPjJ35pi8
qrpwcmX1S10K1hXfw80OJZV9xnRhtikIf3QbSb6JUZj7OmQnVlhjiDQp8Gwisbzp
cf57yyqKlAMBxawjgMabYoCGjoDGoljCaiuY11wyb6Vj+bni+u4P7nuPc1xQBg30
t5pLj/Rug/dQFiYQfQxmUxx8ns0UiOqLYJyhrYXWDsCKbUai4W3wEFVlktPcw+qM
r7ICKQD00wFDy4N5DK0qLn8bqo55T1Fzf8PO25Mna5v+aDXgZxmsMBWXmjEOj+RY
Lp68RaUCdy1Mrn+Y+PGt1XpsB9msZg0/fA5w8nCcoxkwHQf1IhEQY1ldhX1hAYOE
QpU6GPntVqhbH6PTQ4ofSZgXawCf22SnHz9JdTEHXYvRb1uxxF09qk3KEnOr7clx
B/WWbwe2fvZX/ktyr4I3dJshUk2DWpJeEJGh8lfFxSUVcfOcjBaPfbC7p1/vZQeL
d1pK5GwrWWEqHpXltPAxpJ98RIiCz79BCU9ROS/p80q4+jTirPo8Yzm2vbyT5hqk
Wn35l2Uy1WsOOhiF77uIwo+GWGIuN1WKjH/WGkW6d5MFVIuWrlaUfQg8fv7LXnHq
eY9fmkMey/tZ24p8P2bSHdf+wMf2nVoAmIIiW4UkmQkCmGxodpQw+bETgZ2u+0Hu
oNgdVVj8rqk+sPHQHlHvEw2taEbSmAY7Ps1h2Ujn4cnFlyL/F7Ick4aMgEXpkVfp
R9BFpCM0or7nXgP+L57RCJxO1qzzc5MECtYK5ogWrpmMnrrjKOtVSKYXHCov2cr0
TTOXTv3WdQKow0Ny9+NS7Ks2/46JPEFKlY/9CLw//hOP1IlBRS/D4OK1U4gx7Uwl
VGZCFAFMPuWLGw93bb1wByDj2K34Ob1zgVQo1vCcyEZA22YKFb6u6Xq7Wx103Oe9
/XqZomUs/4JG1Vl6C6PaD22TtnnGZQhJgEaodkCYCu5bwJdWZMUBEjRp0s8aYlKC
ZEYG2vUi/PURd89Vars7Tv/EymRdMszP/oMNexgtoTXlwpnxbn0YpDir0/7sx88D
kRkW/0+O2IkIoHuuUyX0lvYi71SbKQTupe9fAteeg9MEBU+kngmH68wg9LO1Yi0U
dn2MwUaozr7MljffYofYn09Nqg6VZf9It1kROP14Xba2VeCLvU0iqkTK/lCbmJA2
61OECksHmoiWJGN5Vf/pfLAY2Rvdb35ezjJ5KIgWGsPdRk7JIAq1OP4R/mrtL54Z
+EVgVVTlt5/7XAyolN6fMYmdDK2D4uhaX/gnbEmkKQAbXol2y04/lxmQFFlxYfFL
ymNhrtJ43ieVB2acVe3V9L7XytIhcBq1litfzP5g4w+9cP/a1XdJy8TcTpn0ur5z
57heCjIrs2VpxXf0B9Sd0rAWuXvlqfaghkEudeeUKTSDTxVuCaQBK5Vdihs0wMGL
8Zx+9TsN5ClsBDXsXObokzO1s1Of0P+iYrd4Q3XhucedgRnyv47UjbTimTBT8cw2
6TTXo35v5awlDWSebnVcvwxuOANhoDIszmpLpyoJkP7S5hEmLBN++cAYHgX1MDw6
WZs7UUCIgenG99OmUcr60NY5AdvtvNF1PcknFH/3MMt/9wvgWJIFPMF3aB4JCRK6
0tv/XT6AmbEJ9PUkbJYmbDg/aXWqLuV9yN27qaGCHbhx7S/uyuogvNn1QDa30CbD
4D5ZfB78uXeSIWBCqsvOgYeZL9f7/76WQMkU7RrcLxc9lm4YycucXOYNS2G70BQW
yiWHHSeCw3fsly+4sMqU4ks20G5tsq7xrkSoTzIjWaY70dSZS1IFqcNPG52Od62n
bRyn7A2dOGzM0XGN4nJ/iNThJJDVk2e23R2f0PjevRhEhrHqyd3BOUDfGdwBH5jQ
QwEbfg4xjmgcKuQnkZ9v1dsBXn4oODYd1vULGKT2qF9d1ETsCiUyB+q2YPIbzcHw
cQCYBNBnDmrNeLW4V/EveJMDCMVrt27BEIZNvHSMW5CFSKApkUiVPUB6ikKwbBiM
Avp1wUMgkCZPdnVpwSWEizC0UYr0ChVgrmZz7KetnpxKfjeuIjmaVl3N4jgJQY/+
Wa5K5dcYNIQmeLCgY3IQejqV9eaYMIIf2Dpeq9OqAgqtymV/CtsKAs5a367aqtx2
tvsTBzUCJg10CF/zJ0KOsXrjESVYjBuE/U6s6UaePE4JdvDZ3cN/ZlDW1jfgb+2l
MXoajpIRfTZJxXm0lofGsf6L5kekFXFa6wKRF6LXy2oXjoz8yV6I+uTyDljwMYO7
0W44hTxDpn6YH8CzXT1Vz95v0KtCH4RNKhOKQotcsJOiRnEZCAjANaDY5qlpIg71
7mMMy9okteB2/hmzjjTyMRWpqM45QuY3C9MEqKYDoGwKyUD+gFpWO+YjJCKls41y
d7rQoL3Y7takqkUftKFNhw==
`pragma protect end_protected
