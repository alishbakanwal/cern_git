// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 14:01:23 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Eb19j1rQzEEnnGIi/VqgVlXzptYnRCW6yVLyfJSnymXcd5tPKqsFP+eAhDvMc2cA
MikC/V6WSvl6keiRNGbAXDMkzQByYm9i+2TlLb18gEO/V9RL37m5CFgKnErYugrN
aCH30CuGbLisXuGglW5nzWvZzocKrAZ9bp+gZyyf8OM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 47952)
GJiTrvCuzcH9f518TBs7VJeJZEkkJI2A70kjsWb4gDL3EeGrMoE+aDZ+b1yjFy7Z
OSxupHDBxiJvux8QugrzH9H89S4SpiII9fEkz58a+G01xOIFZc4aVD4ttfH3y1kX
FFEfbpX3ptsN5HYSJo7U6WjbgrxbVhVJly0Pxmwrl7k6QxlWHIEUxohis4Kh9ymB
DGzupkoqUtM6r/IAXimTiPiHInvUDo7P4tPkLxdBb/Cp/Ghm6rM+J5XyoqI9zdpn
FzQSWO+atx/bSUgGgFzhqTLhBYTEub3P3LxSNrp20gLHG+6c98/rN+oIL/k44HeQ
Iippm98eoC2jupO+uT6gCANSXXXZlg2jQXuqLGA6Hu5aLOPNAVIXgZgkT7L0CfVa
beGRtgDAwhMYbe/sXJ6nT4sjGlR2a1Aej37D8N6VTH2oHAw1Bcl+FwPfZUc7luFw
ru4CxQVrjiRFOr6TTb9bmbB8J4s45fd6wNYDYPY+zP6W5skTgXnfC1Nt/UJCkbKg
0JQeumFJQ0yqaRjh7ZRZdRWm3xv4nx/MMHCn9sdSR0XuMbk6Nys0ix0Hw14ZnHlG
mFNauAK3MOjwG4Sl/pHc+attLElxHZ9gwAr5QCRKxeD7hKQSToxHhI5N4tvuVVgS
Ba+oK3Fvgasbacuw3XjglmmShB7RkD/Zl1lTVSuWI1Ih/HY4aCGYumVVy7oqQ9IC
iM1BmJPGXXmXNFxDhG9YZZLPq0U3cx3Uj2mqpOJBH80Rn3Htyb4wuxDBFNPB2sNb
UVhqBPL+fORC/eR/cT+N6liKjIINTWyLPAnAQ2rqRjW5qlq17c4SHNC5j4MjQSDu
V/c2pmGNtzXHcvJ4HLw6zQ8eIfpbhqqmPDkRXw4BD/ZY1Q9f2PUPRDVt2rlMvbB+
GeMLNNK1jDS41D99aDs0JAtHWSMzIatt4nmHmiju7+yB0xH5ls23p+ATmfkFQqfF
Mwabj8zk8lGLxYdlJt7i1UUcR8uj4FkcFJYHq8kCoukEr8R2Ww2TRa7kC7uVQRtf
QT0K5lsPiNtM38goZ4srjmQGC4eQi8a4xa3Ukcf8fsRo+TAH0rbBZ5A5k9nPkLzX
K/CuSKhtweqlfIJ7TsdYy1oMjIJdMi5oi2VH7U0xucl4uptDyaxrcUrLk7noNaLE
4y3qVyM38W6WoVqo3RNzIJfXZf9TymlDyrKtMyB2hq+RUDlNf1Z5SZ+B/ypVvK+d
GpF9zGWoXmBTf001xUHsJ1ezn7rKtkxAlHX8X3edhH2WgA2vhSGr6jlz944F51xi
5DbSaLd09T3v3DwHBngRDK1MZ+U+0WSiWj+K5rESq6ApMG8lPXvd9gPKvAucUZZ1
XH7fFkhU3LMMryEXJGBpORrLlQlJ18/QV6IoPyCwEXekyMdrKTJxwDl5l51DmXuP
jrYh0VvPuGLGCiPk/IzVqxu8Aqm/k3YtDZQLYjiHQCNyazrF1dozFBcbjv0UTe3G
KPHDw/oJgMQ1WmxkVz3lBdr9edqqr1clVhzK3hmyjOmMpKVgpvpWi5bW9iMuCw7f
1cJbNQGJuVUVv268/gUi4I2GVX09RHsUa1sQDI3a3g9HQLO5kHJadXF74xdlI2GK
1e0+Ky3l7d9IR6ah4dlToe9cQAwDZaNwyL//v8jxgD13lJO7fZS/nUZoB0BRhTwV
kt0+BNuio9AA4NDtQCyvQPNuJJyOhKSmGpQdQuPP2eCRLv3kq7pnyykcfZ38nUk7
fXFPJmypj5I6YwruUpaAmF6Rz5l1IOXGYOJslZrjBynMJ5dCX/GGCijwMYekjfD6
7q2RZ7bkYuHFuDGNtWlkPTfO9k+zTAKwblSsLxKkfamREE5O0NRiJj1u/uRwydwJ
HRiOMJYZ6ST0SC5CUG+Su9hSkvJIh+E025BmcK56mFKZrDa4oktAM2xKGYaMUBKw
GI418XKODlY9xVjYPVuOwuqtOwoIvA/TKhL1IHoKojrrhQlhnI16OTJdlnGajrXD
gNfbIwuNmor9VEPAwVS4FG90D6fCIY2pJXVUgpLQfKUtd0ccncbwAB5VFnGyy8M0
ywc88rasNjxWjOQR/65y+QQxmkhqE0tkRSKGsYNdTZIsnyTUuz/PVvD72YZWalv+
XX5DgGH8hkpcBsalPeI7w/GTsLCzUXBrUp+fK9p/itpp1pJbaDuIoBmvzHC3cWtR
iLfjCNcEn6hC3D1zTJQ63FF5wrtyff7VCg9a8mVpLnP/5DNAbPJO1DjdwbgjMe/e
mcxftgKrz8HdscXXl6cyxwplCfg1S71GR0GTT88CTga7o0zPJIkP1LhgeZl6l1a9
iorDsUEDxIS3BEdTPWp8Ycfabv4tgnqwuL4Sen93EhejOu9ArwdTouBu65ypNawc
Ucjb7kjREiPs8v5Aw0BLRcqbfKyvA2hjpjkMhRHAFTNAXbjNO0/D16fXgSjWdgrp
Br+WYdBEpTWZKFds7IZo2tEBb1Zu7QxgPN9E9IPID2jP4dXFd16YYJrHRT9/rqEU
3PFoVpx2GAtDvQVRFa5J1Oal8v/gb/z9X9L++JBSrXKxMpeT5tx9gaWR4nrbUR1A
3ai2Wg+8zCfvntLJThlGnvFj1Oxs6z3785oixU6cHYkZrxD3pn+Dk1frNutH5Zpk
4/zObWjqsE4DuUGI3OwHgJ92qmb1TbnIF2dAo9+T6AFgwNZj6gWQVKN2mTqnlxqY
imqtJGomkrmflxpRL4I5oO90bGETBmoPGJMtObyoNojLMaXx+2sdQpa/ayPyoTw0
Cs90xPINt0FSrwVbVWPLT25lSIkBkv0CYKaBJv6AFyRo+kWHV1WRQdMcBoPOs2FV
CrSAWK1o+ISoh5SdjhCOG9GCIItx4JUC4Eg8hK6yythMieiCu80qHZWWrUNEYJEv
dgpvmGIQGF1MQnVtHXfiCYhd1MraMx8yEqFyw97YDcNbPIJb4YWVP8s+qgjg39ZJ
tNoiwoVQR92hVUH8UKE+LPEsS9QJJdUPRRyiZ7ykVLNY48uw5oG3LkQRtV0ZvBbj
3MhIItr7eW4SbWlif6vR8ocYbbAmYE6GMbrdHWEBo0P/swhh5fLP0GfNDVpgC2wn
kmaG1GXVKrB+Z3O839UOAJVf0/8mk5W6hjFVi0CxawJpZXZeIKAUQxtZJxSx8a+P
R/Ypy4FQoCGlo25XFB6RGikXkpKpcN1fbXt5Es30++edBKl79UVtoHt9U+1P4G4e
GSh/g6Hs3PkNtdCRRrhZrgXXlHigek5IF/qHIx0aeCdYwuwSoDr/H8yBxrnkXPAI
AbY7T9JJ1Qkh47W2V0ixvaOlsO3WnG1Ti9QFRFdrT69zuFhDxM0NPPjUuyOZs7a3
vGzKHNY2o2KeAn7YgsKGki/F2quZWA1oEc4ZzVIyeY4kmxWFi0fv/ANvb1uX4aiK
SO6EyoS1lnsRTEvzK5Q+lELqk65APkF7f/5mj2lXfEgmNzhKQoFOA1jRdCNYvgYF
BJSs327DljiP66uQa+P65ky3u2ehDTJ8DZ/jndOEKtMAPcnI/CM/7FZBUeJVQGar
qkY0HUohuF9aK0n19t5abh4q2NfzRlTvIPgw/m+r9I9ZrroXAA5MHceURJHC2X/V
4+aZIbTRvUfaGgJ7rojQTHZ0gzDZ8ywssO3X9R+ZTchychvEGVEAxUtb1QoEgAvK
Ouosm9OTk48QFst+RrH/bz+B1bgBA6BE0N/J401q58GZVjiH6izAnKu5jj8caH4P
nU+wiG6jsCFICvKFGXmdDsovsHthob1Zb9bDl03Tfs+IJFJfZlBXvb6Ps8FSlgaX
bgtplI9CVrg7mHWUIu+SGETGAktBPpsglm2LO89uZyRZMjL5BhgL/jqyuK2taZiD
GgjXN5HBNXZuQnQkJmGVHEAgkT5/IyB1nG130E7O1GsUMBPTAALm5haYQcboiSnd
6y6ugyMPsskh9RFz8547Is4rMo1ClDdyQMZTO7RTjNGSeUeAer5aEyuRPwfFHyOd
7sQpNF0TJX4tM/AkUz639QstmFFPqORY33ArUTsRmcovf7DW7ACumsLql0xtqU13
yJw3o6OjyGdr7pdvhzYYQbVUnJFeoVeBV0N8NQT5sEURTOgA6XAix8yHUbtEiu5U
UOFgcE0OOOH40+7D86iqaJr9ZhfoZcifxqZCRtECqqAEDFHX8Fn+wLBIguj/eDmg
PEWe6o3U59u5J9cst4Vl9QhL1NkEesdM/rBJXxYsQ5NXmjQjBzOnDLlHvHLIi5zM
K2PnCRKPNBs6nkEHFos1LWy40WxI738m13EjOToP9LFek3NNv6KgbhfM6A/w6Pgr
moFlZKvARiFPMh8UcztU9nNzyTserOtMUGRKy8vkh+hzjX/EAwwAkB/i1zhWs3oh
GGwESFrjAN/mBwdgMdByqo3coQY1xljHecb5Fc+XDxkMSYO9+glzCjwbjz20jfYU
juJw/sRV6VForydAUWndPnW8VhPOZKweXyj13NhWCuVuaCOuLaizeueaMWb7HrIy
YiWswhfJFwQslaIdJpMAyLZTrfdrMoFSm0+1Hkdo5B4BDGf21L+PyMLzHkFRRn18
PLRFKLcVunGFaFSsfXq/zZIf+KtAxz59cbRveO0HllG/RMNJBwLVLXddNqrNlDls
sYVzGmsYwML/Mi6uFAeVngTCwiTlJyxD4Yk/gA1qOjkDE1qcF4bOjp2C2y4p3hmu
p78l6sfFwq4w3mEJunN47xZ7a0QZXNYYIFZxYKkzcNTd2AgOIMiXpiFqopV6QUCZ
i8CxHBHx7tagHXgzD6WCs9m1k+nk0a902d/hzMsLsGRMvzOAwZiLMSUxOpv1F261
5kq6E/GIt1/YRUYysK4VT2T4cM08Zsp5S4yItStj4VHwaz3c3/UW/Qn0LflnoDu1
rv9IVmIdWWHFYs2/vDOsjJMmdbGT1hghRaIL/Whf+yD615iq6BSt6G3gNIIE75qv
O+wRhVVKA9KEc5rXP1yfaPm6pvbYaq8yIlbWfGqX2lXejVDvpaAQG6HXLU4GG4OJ
sdxpjveAjg4ET1ZsfJ6d6KqIpF+AUMPGuN3Vac483MqqDX2JVsxVbg7fwAjMJRh9
uQ9jhTYmNPN9TsW9HvvvKiPmoNWQ5jjA8tS20VL1hGKSMLUXD9J1grDD5FRv5uwT
ChhPL5hPiw0ToP5lV7qpwjeAThvYkCTMYcDIfSYvb6wFzu+N3QzAun0zb+rIIp+M
u5UL9qLRS4HXahSQmf836OMudDuvgb1O5UNMIjGnDOTLhzfjBgVx0w1sdHo71lz/
KMdPKT5NyhlhsD8MNc+y5b/mAUTiDVcAdu1WJRGSxpY5YGJJyTuuusT5adbrqeZn
NCtI02u/qJlryzR49q4U2oNNSuXzymt/4zcJIM637FlIEDXR5gUMrYw2SysEdauo
iwTtXT9Z7ZAP/5Mzcwce55amUFwg7tYo1lHRlRpM+CW8D085rt9ocQ8XiX88tb1W
KAsii4tjP+dfmtcFJpYz8korSp0wQ/8Oo2wwFQjYd8FxYl70cStAM3FyRpicuMf2
AbUp1v4sD186w/pgXZXT2sGTMOC/VWXV7TYQ5+i5ev5ftbXPBS99EhaT8vw5a8qP
Np/mgJFUTwMcyCOa+oG/bgOZrcqsPxifgOWsgVUrAqs53xlkG1PnPR6FnkDJCR1Q
mTm+xRCRLG6D7Fw50nuiCAia7Rd0II/n9UwkuoEzDUxDLK22oOhO8hIgF397TqSG
Dq8V5V8ioKqvf+U7g8gPWJyjTUeV+9LBCE687comAqiLmmM7gbNkEBC36RZUws0+
W8JrZTU0Pi8oQ28q83rFnBtZ+a21cNmZjxpAWTBpuV6q85K46M+si70y9U9ffWfa
iC+92TSN1n/1et5IlXnk7xx3Yr3UoNdiAQNm6u23dJtC8SYnPF1x93jc0Lfu815W
zkOskYA2DorMOemX29W/ilBhFmY1Nz9BqSyZupyE7tfewIpvwQ3v6tIhEo/3E0Dc
OsmF5ir7Ge2oQz9JNCsco3M2zWk9eSTX1GVj9ehjHD/CsHacsfJVTq7UdzmY5v3v
NSQc0q/iM0J3PjTUDa+Oka1KEHeVk54a0KjJxGmnEKLvSRO5FTJKXgmmPOORn7yT
Agms8eTHio+u/IKA6h/Vy4YgFtqkS69vre0vzlVucft4e4Dc5lfz55DlfjivEgqV
trj7j+NoY6GbpFor76QgUOgJhTuUpsx2+26HBhmJJHKugaeLU9Xk64xw1Z4Xmyaz
rD/Dj1q5YXujKjFTwT911E5TayLKD/VaOrx9MGV2nWm2ZVh8gzMBjIcwDZTQYpJg
BQaWzDzgDvYMzBtMDJQn0lwalyLj5y0FkRV2Ooi45+VqSVourx5I0GmnK3o/b3ND
ucWE7tPiwHQOkTU6QbLtl2kHjj9CNV2BNnqkWlEmHftDKF9fw/1UR4WVGGQ8JALn
ZACLeH2cfcGrSMTFufeY1rPbXk0GEldzU28q4hXuzzSawJJxLDloG+NZx7dy4FK1
dyRUOiIv/dNmSfwX56Sw7djr25ENRLd7jyE58Q4rHhIEuwSwjfEbCpDbSZfwef22
lMJ/BRB+bXYgtKtT7uQtIXFsKtkw8WVoVBS5M/rpT1TSa8ERVMzLfRQFxpAiBvY8
gJhVzdIaTdQCzWNnuqfJJXHY8iQZ1mJXU/AFhTHcZwmupWeZkOcAp59nLQSVjzO3
NMOHnN9qAuG4G2xAbefLen9FJ92wP/nPyLDfdsO5kbrChuqR7yNVfEKRhYrOCPns
qLnCbdeAs7wkoPmHDUWGG/XJZAFItjKBegq0Tp0clsbOud5sRp8C9HgSCZ6oSeRy
1ZYJ64h+JAu92vt30LDpfV4DMrgx0ze24Ui2Lsu5ydZRSmZmox/4LsmjtrpYhkLc
/rWHZaHzF9FDhZvH56j4n41Ji+ko2f6QfSzEs+GkvnkFnuPG/ATchOQa9ug/npo6
uxczEUYQ9GRALb9fNgUJX+GRf8+94uVtoOUe9oRIjUqWIb9ZASTrVVPbVLQXzED1
QDncbr5CMcv0pNaB5YuNsJzKRhJkgkZz7qTjvK7paAhB0kepc+4+R+/fj8ZBHOHz
KHHfe/CltWOJFJObIAbfJf7EYlDWWUNTjD+xQ6t8ydHGVkDBReky84FSQi84JpX8
n5msmnIZXWKviDHsmom/WrR9Oogoq/RttzBwuIi9Ya7rBWm4QvU6Ho7AQIi8o9cY
gUHa2LTVtsywo6gNJHrD5NGWFU7HsujLKK+ef4q+pkvGw+8lEPYO64qZZkuTHqmu
7ZKnz7k7jgYJvuQffTZ89vjX4+dTVaE98V7s9d7K36D7utIuucJB8Rztto6kC+uI
Jjs+HBp5yaC+jSM67xyeAPhb8S60L54Sjt2GjKku3vRtmeZYKJN50fLWy7Cgloqv
KAoXbCQVkUvzgxyMhdNvwtIy7IC/KnqZgw5EyBJFnazUfPho/+pp2hWbz5pki6nM
7fnW0xEt+HVboD9zawqDmz4dPZNjnS0bXrud8sm/utbCfTDzIEJ/+07QkjrNVdms
gKFFFaH3c/dNYgfrBSUqTy5g64oLG1FGOZEckBFPOShBRxA1YfGnB5xDpq2KdLZY
h9F6+t0jUQXnjqaRsorS3W0CKchQc95ebsA9HdUe4w3NtkvxnGqP2RSUH+5TUuSL
l7wIBdojytUYr4rOaloxXVjO1hkW74mE6Xrg7xSCxfGYH/wvL7g22dCcPbJNs+T0
EXvRUy71WPRvep6IJP4rUt7VnXK+5aiUpny4y2TBotXrxi0j2vSq4YtiCvTQHX8E
HvIV8dKT9lTAEDLnOMrFeuihlw39KDgcb6Ldh5axfF7HUN0fWoSgXTo6B1DyaKUC
XQDJnescNbQDmiKNZvb8hUUmoic+8VzfCki/b0dQqH3vzIGwlo4coaT6hUC/Q1E2
4xK18A4c5alNISeu0tA/gy8cnaCaUNDrZo4hpbgkXhcwW5ZVKc8GmK5/snWSSzJ6
zycFB9th4B3dj4csS8taBUclVVdUGziqCV2U2Y0eLRonrYdNh2HcsqHEifASNUJv
pV/Xkxrh+U6aFoAMuPBLijdZtffAYPCZRnwrKGptG7rz1CTvvEKtl7dCOgpSDmU0
ff4Nix5T83W1NXwtiJMpFWljE2c+KkjbSbKI7RkxhYR5QW8s5wj+HT9FhkIwPu4j
uD0/xaC5QwAPiOh7SG/nlAjMgI5cexQz/PXfHpt3sd0JFoqgr5J+93ugqqR00d1v
X7gHE3Dgsz1SkWKfdICNZ+wz7mNlCxMg/p607fYDBWlhpj3tBIZcAt1uZUvT6ICW
RnzFTv7mcJ9hDVlELqNc08MZcAPhqVoHFLRqKyWSP9sKBYWmOf2KVXiaFTB1MLnr
Bs4wWtw9d8Z0vHvhxA9Uhr/3rGM/O3Smg1IUovFXMzUfg+QBq4W76UB//exWLK/H
OkHAKqgLpR96XuL/zVDS/BJciwFaY9oLHhqJbUMFCYWjUb9a0RLTtF7Lv3tfRKfz
5EmFHxNDDaBs06KT/9EA0qxCWcAyvVCJQFaXeUnYvWBy1bFHsKaOsLl1c0Jg9tiy
+Cv3skWmvR3UP6tnO/LA4QZY39R+FdVm4MxrmTQRjaqP5mZdoLLVMEOXrFJk4c50
aV06D6kykLWef3abxA9/MoXw/GJv+hVC8nPCHERlGCatJyaN9mt6AH9LZm9R9a+O
fDyBzgILThxkh3o+6fEyMuvFiPT1VxwqS4ioIFWwP7H2MLBmjs6GbAmAS5lWEGtJ
8n0n2JhRSiQfgQEHs3z/45AdCCrfb39lPyCtygeEOaZdpD7vOvxAS7gxpPOoBloN
dulb1WCCZRPb+v4q9ZQcHTuiHfutCTWO4fAxnxbDcbBz/38sUqU7r5TrjkLawRfT
DBtH4rcofk208n4wrXwheKiEzJK9lEbzWWl/Ggzv0jlzQNu+ABTYQ0a56wbLs60G
kbWdCIQAV6eOJKZa/d+jxUdKx4Ur6m5sMv5c6CtcQiLo2FqfESKCEPKccGuGXkuH
LxPyXWMTCD7KccXkUZ4HJ4JdVFf0cTJwgWye/8bJoLfCLjdeXdNuhYy0L5b2ORE/
fbUhSNobz0yDVG9wEms4gbzNGKSr3ns51x1XJ5SeXCDY1kUK5SrBGO3oSFHC80MW
72ZdrJfdnmvLdtWVXo9DMVQ1ERX68dZcFIF3LnlSIKFkx21AnXDCMUtm/TppSHtq
+AG+F8LC4mFKYRr8DP8GQPR7RAQVQfQPJK/rhwYTaTJL5Z809lnBlOQYYkKI+FrV
+8EBeKat2TkX+snLocezsHvmzAME4Oor+qs9NxGrgaBZje9XDkjc9XaDEJYqpJ58
6VStkdC9iTvx37XS9Fh/19s28vZo3utOS4ZxRltL31Us/q+DAxlB4J1kAt1nS5no
0dSFraksIQKVI3FXQhYhP4KzWQ4Iwe25TX6uwe3e+u3HF72AhCF7Qx0nJz70lyBk
kAM5X6xLwVJeXpix0HA7JZ9A1qJWwzIwDjvr3oU/24qPtSKhJiyLtcRzLYA63idj
BbG9gutyU2paf5SgetnHyelLmtUcPueDYJi90AVBU765mDHngccVcbs6u3vbv+AC
hM//GpW3m51D5NAF0t//fcw/3XTnxdDK75qMFS+Lx4G+uyzFssuFdWbzchOZ4ALK
VdWDSw997hXgSWRAFcNyzHEtmB3cOLCBXpwbEPTUpyMWNv3GX7oLBamnnrAJhe9j
P2tkPLiL9QXf74rGxNL/bi07qC3jw/R/X/gLIxS3966IqFsvOyNlCoQrLLJMSJQt
ve/KyHyqEkLFI6nzzfRuW0myQjkNsRWSWE5xkWSjNAd9e5nvQXqY31mTtFq6ruEs
va4nOkwJyYSIAcE8BkiHJ3UyU3QQpCua3hQkCOzYsWe5snpsOpnRPFoydpLzQGZ8
72ViVVyEnsTLa5ZGr7C9IOA/OZQeoPBf64cHAeMaidnO1DJvwdk6DyIzqrKHFz9a
C9xVuhKh78bStijdMGwMaba/GDlU8TfonzFRJpxs63pI4gywbXYTPYYJ0Ek6bA1f
V4gW6fOkT7zOSKxGtGgAgnSpR1/E2z0UeF2HO0+KiEN6rVGFhATFJCadRxguc3y7
BRgFLzqhUiu2RtMKUZCOn/NcJTuK6UXmcbn3Jxhi9cJgTYXnhJqtdeqM3RPjk966
t5j3aRohJeqg/P0Z8QiUK3ELPibNqy2PbMdBKSUvViCl8YE/sf2IzAsIVr9F2TTr
4C2MXVYWxaz0E0zt28T+Cqw8tWvSt39CFEZmC8HigXIAIsyMWNHACIvhKg7ZO0cH
R93BP7kS4I37YeyRaGnIdATu0PWGs64NzdzxxpvWhzr00JMN5ZMCR2Wq9Hpi7pt0
heWcDQcbGA9tX4qT4NMs37amV1dYoKlq79mj9VTaoxoOiMPxI40yDcMx4seuhu0v
bbGVZ3ZS/Ll5Gpf7O4WCBcmK635G+3H9pkfxLXQ8krvVjbRK4PQFcLdl+RJCrNh2
mNLg8JCIJEZVS47ie5LeZJvSVXWs4z0cldeD76V3iNSJ67GlpKuzzITJZb4PuAtB
Zrc8XMCZKZmD+dejmFRrbBah2XIPjiMMrbIIs17QxeH2gLH7liTxIqjqIqzjQAj4
698SaQq+VnGR/1nVAk+e+BhlkAtqDeshQXAlmMuadOUBiVQlDtv4otiO3ErqhEZW
2Mi6g05VJu7FAmND8uCzONUaQrN+HvlnaHzW7dIbxkkBIv2EfeWlr3u+aZPOk+vX
T6ZbPeiNY0D5iPWRTF+U1ZkW2sAdkGYIgoO9Xrd9swFYFi0ieoc6L/pni0/Sog+3
IL/JRW8FDIt8PUDFQLYNJXWUk8J0qes/qlGi0kVhM3s9NGfEltr4GRjJZVXI7aSN
cc9WvNjhrgam9jSYjngCIY5qNdzbM4XGdeiknwfszX6aAaUsMIvk2dRNu45ErmDf
V2/00pKH/knW0Je2ABprOK/tgnyg+qV8y0hB3xUU426ulUUHwXPE462Dds2iLHBj
VWajCD9r0KSt4F4d+c+xZEzQiSsqK6GLjWMwUWxKTPN7RrekJZMzn86hj3NxmcX+
kNhaL7tEN/mGxhY03YfsOD6LbjXVlx0M33xMgU+z7e0Hax/LNSZjeCkwSGfvfDFS
gahSENZn02BpEn/s17Sg6qvKzxGnhKDchKMiplyER247kGUwZTNZsMuSxKt+izGL
a3KyKlz77QsjJHSrO6E+l/UG3zHYJ8KCcGcDIqv7nye8S6xZn3Z05O2ah7cTPKyM
difcLwE89wvlOiiTbyc8wD37aXR7CuOTc+qHk0t0gqsuccz34n/WYsvfdVUUsqx1
xLiscFRqPvcsC0JJde/XLfoAcL/wYOiMqFoN70tFOw7UdpGipRL1A/4wxjQwrAHl
oXeBgEv/fEHcRUMNiY99GO+Cnl5HUZffRXygEGHszhdNNlW20mwHJQ/vM/Mzh29O
rVb0XdJnfw0MuO/Vb2bVMj+W0M3f4QwSRUyGLD4XC1xrQeXyrReZZquwR26dtT8c
QOHwQ3asNiPWUSv7VFgbcBWFlC0KbFs4gBVwAOQxuZd2m0kiBm9hP0/w38VtJN+u
UKBilJLQ9/m0SvLUYq+Ht2CFvk4ho5N8GqECajOWnXOuXCxdzqfzAzUbCNKy/3bQ
Drkt55k9jcxgbgCgMLZTEJ4OYOE27KfHx5WPb2IJDhbr3396QhXK6mm0J4QakEk+
OsLYpgR0GYbtncWLd5wkKzaKGSxFPyTazD3V8xU6t3Klh1WGRBpQkrcYfr70t+M5
7JaAhKD14It5AQChppNqj1K4n4EHQPYQCHflRcJvdmzt3mPbywvebT2gNxUtNrba
TU7uYMpLAU4apaHx8k/X2cjfwDUyb8fsYayt5LzGW7JkmZS16gGogl9nIdbuIOFh
W4d51In5H1ZevXvS6JcPA4qUQpxaMFW/gYnnZ+Zqc+OdJ2TUb8RusPGZ/8i6KmGA
w/YdmBtwYTY1TIzdqNP202HkPh15QwISl2YWjDXs0I2r8ly4a97QozhFQsEgZ/JO
LSKMrNST8rKHTjYZQxx4BNoFujMAK7RN5lFzmlwkA7GGNwKUwf8zh/7gtTUIiTQi
DcMlmmLnTdhsbqwSuX40KdfWSnOk2T1rzyzi8u+pTMqSrd0ySXTC/rzBWC0Q+No3
PoHaYQl3J4LAYWn5WtaKgkw6m91YTANG88UfHhAOZV1Dug0acESZjD5ay+wM1/2T
mCdQAup6tTKXbfkNlbHFtpD1c9fB1dXSsATH+LlSrTZHSYgcgebpQWRS5BbWdMNU
g9YoGb5/sMxhxdhtZ6bQ+VMAlfJ5sUP9Nv2YQVifXbdqt1ag2es3mQCPvdIvuL6W
mUz4r3fMlKEqn00I4U0a2CWAWuM5S5KjvYDNA7kksEhV3wmcPKbpooP4DvpfrsVu
wqjguF9GWIxGeWta1z6yH+ywi18vccGC/z6fsjlZMVbFG5vgkNyPnbwhDCsvo1Go
oU7vBEnCH61TkIWl9OBUWTfPpnkB5ikiBRtcycTHMUnxc0KnkBXBt2rtjJ9GW+3Z
nZOyxeaUnCWkQiDrf/yOvycukyv7+IrxJxRfGieA9ixW74wik3+SI33r/j37EjrM
MBoR0HiegvbNtboOgg31ICJ8OKRuebbqOvzIOH0ymLfe6pxJz99LkdZYsCkCyFyG
Xn06upEE3LnjyNlheJAlbfnzv4RnD9qnIP3rslEjbB4K6vP7Enn8qrwm5CCt/Wic
5pJRd4OEYce0Hso3saTSLNCjoTwHm5D7UlNsld9XF8vQ2eo2kJ81WPDyRhnfQVSa
GG0b8SoZjhkIWKaScVdmcGLttFbSXnmcDlTDFGet1/ex3LjskRLInk35hmTqGpkB
zg4Q0n+cykfurez7ouJObrIin/y2aOvAxNMVbrgn0knOvbOCFuofs3SUcIHHv9Z1
GXzaRBB9S/PYtzOH+z23YG6xPF88KZ4hjb41vn7H116Bv7dhV5e2FXZ8o6Rx9pd/
Fqn6GBd/UhxoNCnCmD+/jI/63ZEaOmDSUd7GZw5dUYti+ooVRJsKcbmiYGP7PJPX
0mN/PPs/CeW921vxb0ADoferUa1hWdIFPa7xQAVztmiaA6ryN/CL++5V1bChbu2Z
fH33SIjra1z4O6AbHdu2LwzX7nap5l0V3tC2b0uYaVTD5ekXH6KcH4G09nF9yHVe
0F0bSiQlIR/sZcN1LKEx2yBrm93iuaMhANh3Gjx7gRCmO5YxwOTrWAdkP7NbnZYl
3nhxPzWIoaHrj7nvrf1FbLBI6EP05e467tQdg3fY/l5F2YMc1tcLEA1sAruUWncK
cXKsZW8qDgwVc02Mfhq216ZM880PEqSwSNpqpWq2BCmbL/bo4lxk7TpM7Bplu7Rs
PrUh+hi0R0+avs1zZMt1fynRKI+Jv87MA+jG7mLfZLQmsq1iLcfXXgn+LXyci4V0
hLYgrigg+09LzP0Epbe0intgxPGzcjnrB2c/w5TeMsA4UQ+1zlbamv6Twsq+4ucB
dhIdxTwxQIozBgzhXNYuyddWp4s6bkkhl2ame0JeR1jevQZOiQnPhK5n4xXo84Zj
dGYsY3KtMC/y0EeZuK714RXjlWxxwu6E701/nPIu8EvpPUWcVldI39OC1j6M3fpb
/L5lUdKTGEam7zT7vrVa3iVTY7sLtGGh2dYlWiA+lHTzpbMmtrdp3SBDWEaQB8vE
mX5ndWkiVI0uPKvFPoX2we9icm/Any9EKBWaa1Of7UpQPynnTcl+AknB25tm8qgq
7tguQGVr6TYdumYeRQoZXoJayAf+AdmSTMwB2G+SCG3HgwWcHZTaiA0yvJp6ycom
LNNvfojl9Z8N78WHQm5l7gUVSX8N/2MAQ2lBXqNKR39iR9BtyyUmVBb8ovQS+1QN
btGERmtpu5wk3saMqNyiskmGTOIeiZz5GwvVqxOWfEAGpQaLGMac3nDiSFjILIWM
qPzL3ImtR2NW+wfYIe9llqMF5gbWkFLP2d+/+EcFAD1G7yyy3zeyvkYN7m6d65IZ
09B45L/pQjfFgYXGmoLboYEiawPOUxzmYFWmwgQKnW++XN31lqGDGCspz6cBajU4
Sak3GVhqOFmfxUxDZdfmcSSkVG/iOo0jpG4aLYH+lP5H2La2NUERQJ5udcSlKkwl
FAOVcCDp/zd9LVx6MCYigItHLVldmzj8nt7joWR8ws10DOmc6tqXFqJGoyfeQ/49
qU+VdPvoWnS5PVUUYQliNWrgy5VHIBHGWIEG7VBGRxr/l9QsorRJoT6U5nRfvQic
GcLQUVS9OzgKKztWZSjWUbqyasQgulsV5VeenfXTKwX+fMjcEmrXfn4cW8qafzg7
YStG96jeVZaEVguHzt/PzLN7/D8N90ZzLWIHB53b9GEv7Cl1pNuAWF/WExFcCqtc
SaNqCCkuOriK2zqWHAQxuInRoMRBb3m+yDB45v3tdoYhNaRxU7Z7S9azWCO/5Q6j
vL4mQiRyoGFfg6FjpFqMUbL6aQ6mSQ56KYLtdfkNEHzXqiZq1/n8eIDZ9ypqjjFU
dERFo7My3hEzuLk/gmFnIx1NUZORi2O+zJrUvEl8Po534Xp55I8FzuqCpP69dG5i
EgHvmzN58NlNnp/q4kvkDf2gLliEheOmIxFdceGTgJyv5t7gpunDah8N4XwwBWH9
lSlnh79fYSCKsBTB4s8RdHhQGL3IkY3dxwKiIvllke6+3AdLo4fEAg9qzgbY/66E
AyPeCDcZt3gnJySPid5xyjmkuw0grlKPAFlU1mBz/LuCskOTT1shRBuFykxx+epB
T576BdaAEzRXGr9gAOLFXJfsJ1m0hEi7bHDY3XSFbptGhYCH/+FRuiOQfp7vZhDw
LfijP0b+vf/uicNtMJ2+nbH3m8x9NACwkyXU+HFC0K2qVFcIubjcLAaPf8ulv5/d
5rVqeJGBhb4XUbCTmQNUEqjfSPtQuTlChwzFws1Uc5SXWztcLxGAj5OBom2Cg+gI
emnuAmWrTUee2S03HxN3DkvHBrct6bXTNYsNxhI4kY7Ug+XZnyRPg/X4ghc/NYk+
Nd/Nz52Iy3ATM+d6JQR+uVO+bR8DlsoSJJVwa2Grkih37AJ7dBe/YssriMLSCDnc
OJvTTrhp9oIQLa3E1pbqpqs2+Z2e/5oK772tR30RTYVKhTHrQMpCdb5/FF9SrT2Q
SL0UuT0yfbvvTX/pTITkuLLdfO6DCBu5xRZOsO+peCIHoQmYcN75PQOshq/vvP/I
NhZutKDTTLtubQKiorzQCxJ/SgCr23j9kyf/nmeG7mSZNj4ts0DS9oDcfKqDAo6A
33MudJgtms1sBBccBoCpLa5d7SNGOLwr47rnKAvSiZuEpL+Hg8NJtccJ5d72xGpN
zWXSVXdGhsV7w0Ea2Cq/ZfBl6eUMkeGjANnEe5m2PKc13WFhscn55M5lnm3XHmrH
HHYPzSCz0IBex01g849kzqGa5Z2i5dGcsNA80AWVNMBDBOhCsmolM/ualOQ7wESs
2/sYExfwDOla3Bfw2A/oO+4hN73YcShlvz7PX++dP0WQOmt/ZhfrijEEoDdZ7c7Q
TFK1Ya8Q2WUQ+KP/ryI9ScysODVAewQ5IMUwUkG9wW8lgCv1wtuNtaONjyWXLOCA
SoYxmN4wOLju+EadQ5MWZ+yvowK5Aa0ty3nfQqikdB2KgDp+UnhVY3J1rU3lXKGk
tyaTkbV/vIOn1LEYY21Il4UcufnEhhZ0FIvggFD7x8oPrMuP8mfF8kaeuAUU/2XC
SeCZNSOZ9stLhdNc1oKyPaErUZylD+XbAIiwQYVEZm4PDziuYI6QtsgMgmt1KVSB
u/6qFbPdlxohfJIArHVt5gamN3iAXUmajPvr5tmarqMl5jcB5BSYnZ5ZDDFlGuwD
jLlxTGjygOzf4dG8MqpJPAhzko2oXHLm/8W+aA8f8JrQ0jQpoURr0KoMOJbTQgk+
2dbJdw2tanT1wUuUlDvkERIAVYkiO9pCPdKiv+co9DB53rIWAZ70+RZl8DlGCfiT
VnOn7cfmdQXtLJb8df2rOw7PoAdXfpRGB/9aKXW5MVIXbYr7xYgaUFcINy9xSeh5
GgtQTIN6UCubynVmaUYUcWJmBD7QByis53lD+NPoyLmJ86uCtG+eZ8jb79oVXd30
FVnewLuy5bw5vAiZ2BN4FpXPZxXowYptzHRnmvlyDd+R5RSN22ZnSG9XPpGHOHn/
mmJIp6xU4gVOftAWuuA/rVsJiKQWp61EZBR2vfUzVKwhX8+OimjrhHPMMWskdAqZ
Xu8KICkMYnLIxWkVcrLyOkx1uTiZXtnrwqpV/B0GH6ohZ57m+A8xYfuIwfZD5g0Q
hgCRaPh3zN1XXFH9bbK7ivlXa0O/5JbeSYQ3E0QIs+2Yvj0AHheh8smlzNE8Jtvx
qHfMwxog/az8Pc4nDr2yPlmd49wBnXSYxmamTkc7xnXp6dKBSVqkX8NDYLy4kRKF
yTlbjJ8QN4kjhmf3DoZvPxevtgO2DGKj3ofqksqidAt3EoTfw5hFFP29xj4VhHrq
9PyTg373FVETeB2okW+uaIWGh0MrAw44pzK1RStrQmlpX0oW+SsYYOdk/SPT2yW3
/4iB65x5yHZdz5XcKQKiwO04vpiyQubcEtmLdhE6goE0VcnGGEG++86I1nhcmHlv
DNnXvqAhiUfTAm59h96K94eDVNM6GcNW2VQ/wLB2rWjd7VY+zJ59gDhCboGKFOXL
GC7h5xny5eF0Kj1RGRekhprzcguBEDSzI/UZRef75mA5gnFW+URtz4epZVVifTdc
/NERS93VEs3vTXUACFajpcb5VjPAa+LPHIQTfmvQ4jpIHoBPFozCC+Ec4XF2eipX
8gZqMt9S1kAnKXicVJHbwUkMSb3qhtB/V/UdVQm1Kp6WCNP6f+OmjFoYJWg+Ud/Q
fENTCDvDme8rb8TGGg7JlUfc6lN12jjWXJvB+6I1xR07XwYHioeYQORCpKf4TLWe
MFDGaNKw1Qwd2cv//mjg5cvuWNKG22cQIctehGOTSy25oiUDkxc+f7DJACM0/cwB
VtSpUaloS5cykN7FJ1cexKmvfuDTEdoqZAvdTN3VwLFg1f8G9qZoMu2wr8ec7Zbb
MhdsEzQDBGxsmCn3sInwWeqey40XNIqwT3t2+dg4S/UifHca6ICIRAJIqb10JlJa
i9siQIXgiaYE9+V0AKBLs6jQ15lYNiBOGc6DYpDa4gheQaVTbf/pyf2/5bp3RqL0
+9MxJXw12OE1ZoNWqteLvxSVEX/CECtpV5FlD7GaKgjKDjW60Hzf8euveE8ZZmOd
SuXaJu81G0C/ZD/Wdxt16niHgoP2E2VLguNOInk5em6DPSrbq7VZVNLSCsO65eWw
YFgypxEuasjd2C3YBXvj/sam/NNfJbwVGtYeEnSt7wvJDV33QMmDFrSrN2k+flGd
hOlBtpZCLER5qyvsj+Pz0bnhQTInijhxhi0qeJfX51r19AyXNt0didEXpC9Bd02H
gjOOZN2q7RVz6Vh1ieuqzA/iI+WVzdORNykhwueRMmPVGcoKgzHOpWWW1UUrpNvI
xVULWXhN7EC7g8gkMAxG5kYbLK4FicCEpZEbtNVBi31i/cF3L6FWQ3Ff2VGAMtEe
vlcaOyi+Vd+NXzG7Pu5HzuYi5kuYx8ATASA1cGcpKhJM7kUfYyicXOuoCNvOJoha
E1i/sr4Z+it1zX2GJnDtBVF5AfZ85+as7nVgQXOKrtVPcudC4ceLT/y0OKDUk0yk
IEyJYJfY0BF+d4xGEjQWy6PZzCX8A7j4Eql7UfZpoKBuLsJbpdRs28bbfrPcljRS
+Zi6/hps/3bqsimndaFjoTDqbHDkaznwzWb0rWF/RQ0dtgAdRndM0VVuDiRaBglz
6cyDsiWSFXT+MPIrngE7bHP8Z+BW6Hekpo6zODzjb+u6rLuv43+6CWOihva4SE1W
L8yu/t5w2lVHgGq3YI69iTVJA4rJOHYJmCWjsCSRz8PQ37mKqIKE4B7hfq5OLYlE
nJBm/1uyV9vyjnSyAkpLcob9pJrglP5bj94KSWpaFt+lWj4NCKyIHE8Xd2ItTIKt
rdZaafsQlEKzYDp5ELGIPdrqTgw6mJUJpUBd8zEoHvYohHfiAfl6CIHgWdC7EmhD
1mq9ocj1AP/PlQdBVUg/OWbvhga1FdS0wstUFTMQjlWxVmJdqRGu0zc+JjpQncXB
6qKGspTkohOmqctDnKRgS2uHraxRjKQPXLdkz1jncaAPBiN2sIEJ4a5gP45RkuEF
TLnm9e6iSvNT9dfA9MRx04Uc1wvhgL6vhH+2zN1K1q+3rIDMVARq4oIoTaS+Y63b
eZ0BuQT0bHH92BZGTSLucjDBfJmqVxA8qpsgJv0YKNm8Sb2gSJrrkUCQl1QPGbCd
7MpkrMEq6yCBZ72C6+tGq2+xGckB6DL85ZcmEV6VFBYu49Cm4etS2fIRHWn3z3Pk
BCAbWpTJ7Ah2bXjM+0SWn+7dkzJRO+RZAksS6rC0BcS/2yJlQ/CBOP505RoFkCVh
YM2Bp2FZz/i1BThcqgy/oAkNoLVhI/v0iUH6UucH8WjCfCYnO2CQhpvBpX8c9Viq
mB/ZAoFTA1KuRLixe0x+twr4kx7gYWVpc/MxfvkhPhPYFVq5WuW0RDfLBozZPRu1
2jCtQ0I4l3OzBS4+aiCyfFs27/59bDUizjM2dimBpLy07A6iu7vRc5p1uegY3mFF
xmv5WoaRiMWk32t6w07kXv42lKTEj+LmVrpBj/4Ik2yevRMNy8ufyTN3muWJfhJ1
ZOcRnJk1U0sWfjxBlm+9o6RoCnr6WsTh8ybcz5WUCeoXOEwcgoFjFxBOATyw9M9f
DXVYlVQL68cqNINxsj1RY4k5kVxI+j/Tq04Mga029wZPT0t45WuYYEpIVEpegtZI
3VE9JCOqpVJJUhLW7WI6Qq9N7a0NV+TLGQ62JW8zN+HKK9i2dirFx9GkTL/+xPTy
beDjlMNIRA9N28Cx7dT/ccE93G4Xt8KMqxhlYkRGnSrZ9F/BeToq+Bcgov4f4ogl
VihhPMdOlse3keXOfa5gNhqcM0Yw7PRm9muya0mFe9DTiwArXLX03bXYouwHKmKa
2ObGzzFZb1eEI0lQX8PGEknwj1hwIxhYlErRzOepKt9wIRDB+SLlW+Vl9qulpK/n
Ai8h2Ni4YrJj4I37cs6nk4s5/lTy6wNTvtwVU4cqAyMf//hlCImF7LO2RfqXu0Fi
ieaI3yYymHdfQ9lCDXjaoe/vc34JyuHUWhh/cfHPL79L2Z9fbz5wAS9W3J60Ddqg
VA6Z0G08YuxGQCoQpwJc0nrAnb8An0aiphWaEfeVQETB8ZJZHSU4P3FaVTpew14f
CyKYQYgN8FvvQxvPw6irnFdum38S5/1ydxWY108P2FZVn0SDprvEuqZafh+rUJWL
hTi/VAR666gnr3R567kJb43ZjP8lugG2O2wVVEhn3dGPkA0t6L3aMyf0nA79cPOd
2dfudDZM+qjHLyZOzV73D6q/ndUDHwSXBX7G++03ahV2Y5Hq8OeA+Z+iPWB1O2be
KTv6qLGvV4GLLJprtWGm/ZgKE87u5OOoY1ik8uFBwrJIBlibUAH3lEhKi3Y1vAuM
mMoSBAU92a1dAoztmz5hRK91UkYpMzBLGTFhyI0TDd+jG8EKs20xcxE+517eJMTp
v6NsJML6qjoTlo7OdD7MovOJMlkBGeQAW0BGRI7etINCbLIh+vuEMUeW6nALfq7k
kTcHd3iab3oKY+FPmulErLCiSkC7QmyX+3LLn1m7XLB6HxzCbHZD+HD9Spmv5AEy
eij1/q9hnvQeRyXZnS9yzMqYwPO0mvHP4KN1wJy+X5wMafROwvFSn1AJHO+o/PGA
58XMdUONSZ49oJ8MLYt6boI+a5Vc9J16WRx6lXoQpsFrMp5wxGjtRdFZ5cEA+sKS
PzUUaMKhWtpLavNnZ9RKwWAc2+SXQ4NcsxyxH6udlbLYbWTUr+yMaAgdlJxvFsJA
KjDbcVTJOpulFI56Eq5OOa7rxiE6j67wZfZNFJt5smu7Ps5+khAbR/i+8gC6vBd1
QeIWkFQro+IH73M8Za8HEiTDKtQqdGJWsxOasSTIi5h0AlVHyWX1YorlfKx8C9YA
Ls/JusebWwUnWK+cdZSV3YLFS7BRhNo/gK6KyxfScW6MVtzETDTOv9BzxKNeHoeL
WpT/gpsfLovX5AUhOAUS7NJ+M0tdWvKgWYbzZvwyfLHd1Dnfn5eG2c25zkoRof7N
7Y78q4eSk4qCiCJfRmddkC6YVde2v31PP/DV2vvwgotoTSnsgYoKWW9wMmORoV8w
NHdqLzZovJ+LOskrK4LVbRWw918tuzlUw9kjBiqxgopoi1Y66U95QBHiQ3qu09LT
17q/CyKMvLMik6hoS7aIxObu4xW2pxj6oVbXfofHARNDNcSp51jZsfxrd0C6N/6Y
0dhBvJwhj4YKr7+vn6XsCEPTzgQywTsYabX35fIdHd02TRF262facBmGEbDaJlH/
9mpU5iTlar/Uvc/ClNSeHXgcGRR6kU02OOjD03mZaY5ieicE3Z9VTr+7LgylJvxH
NBT/lh0gSoQRyNKURfOq60o2UOnDPRkZ8iW2YkrSyFErHFBA5F7GRTUNf0R6e8Qs
6Ft39I7+HYrpwo02/9mQ3doudUDT7S0XibUeoGW3CJI/2p4/evXe35NgbEsoQjCe
IlRhwUkM1igpPIaZXmfMCTigMCL4Gr+SmB7Za7wclTfyD2TAjLTjI7SLjF8fe8Es
MQ8PMoyZC16btZ97S9bD7H3pI164reyZpZOFyUOxlBNjJPB0cWzSu9BR6RFHZQt6
IxK9P4QA/3voBBO5yOUrIeMxbEQ72N98eJBJ9x93AH8+UaR3LNlA00Xy46WYTrUu
36ZEEvuIeLZFY7MKlAnyxKGTJISCiBnwa8hHpAtPjYBgVHurMyN71hRB1NzfDJP/
XjbruVqEOfCmBhss8ZMilVU6IRzILvRTu9PWV83I0V295SZKC6R4/c+WxqtIpwn+
lggcBzfR73Tkm5EZHYMlkcvjd0URqi13HmptLMWwBTUGO6j2qTz5U055KeRIVZWe
NO85PcVlDCuGZn7jwzkl8F1MnupCAZWIrXOcY4XdJ+obITdArVHqaw0P1bKoer2b
jrlxNwkhn8wPK/dKzm0JaciRNtC28q7hTRzBKSkKfvMd3RLyXDGuhyKtnXEXyVjX
87yb97CuFw8iEWEcWPSByiEXT+AlOqtsc+bfYMhO3CCZR3CPmu/7L/fIZU/MIgGK
WkA5Kdlf+jsx2DLeBlG45iBRiLFFh2XbZ0et+OfK/gBRvGO49IuyE2QncSFP5D6H
dfHIuA8ZodriBzVzCAomxRy7LOiq/i7lR8FjTYPYLFBcRTP6DGztQWeRYxj5qFh8
tdQu+EiPPqqLYLk3Ixsmjo3AbOV4BNtsxUB1w2BSvvojhJA1BQdp6gPbMdKnXUir
y98v3CDY6IQNSPUq+cCdR71Ti5aAcSn9iqcWKQbAq3L08HEV9nlCykHCTm0uSqdx
VkC34pOItxjMoWc45VHq6xru7aGDkspyTMfc69xgCzsLEM5ATzESHMeSDQg8nc4t
UH4ygpbKQ9Y+lXLLzdzzWVDHKYeXVwZOCuf4eyDlmy78/vg0EW72ywBpPy3XxI6C
gTFQ2XlOBuGCv93wDk60FGlWbKLZFnVofoQtUbiAWRfJi2ik3Vta/Vi8RoeO85D5
LoalVgpHO/bWc4N/gm0/TJ9Bibs+gv5/cbhysIbz3tMXF5nhC5fk5p5WFOZeuJvr
0Gy0N7qsSwrbi/ZjcP1Ci2vVjfWSWwcDe1EjH1vq8xdgnKLP6jedMQ5AtiTaSD4U
YTwfD8zC0PohNLXNOjUVwZENOCrbxi09m/afbdGJpxE+d6LW4cOEFNqk69qv14RR
do4neqLDdK0BQeSGs/++AeH8F+RMF8D1WQz7jzLOEAS19Ui2Eug7SdrqaxtH53mL
DD1DXiyRJN7dbDiknkveSvYDOnlV8Uwpedtv86vTyBhY3wRas2/LnmDbh43F9gNU
Q3ojHV0Mozi8CzritrWdrlG6ITa2IbhH8FJZTje5ZlOG3NIMKdXevx2CdiacJCgt
eBhW0m1QUeCV/BKjkf4m7JHJ2V19qWuwrnNt96xZCUdM/+PDzIUwEflehWq3nuVl
B8JOVpm3D72hQ4uWqFdXFW45BqOJ4QFEqwafI+B73lrR2neZJLdPY7wRIvNMvnZt
fJX2SL9++hQuYzT+Pcp6jkev1Cmj/QEwFn38RFg8v5AMRju1PYrkqOjY1cn8h5UG
FMGSyjImqOxtxOmHb7COtKjY1dPLkK3jnHwaCLHuJ/ksxqLhkS8fpkyWL5OgD5IS
tPC8SLPaIQURcVeQppdUn1QiiVUCijMO+mgvrPMiTtx2OFvjjsTDDhwwTxKbUU+Y
msYowIYRWeeFBC8YHgTIQZ8iuL/BWffoGBxJkZ68xJKZtFUPQYycL6ersSTVpnab
lnBZCAS3bwyxcEwpf7RQn8deBiCnuyn0hvtBXo3O9/EYurVWj+uDlPUkhR2fqI4n
ZoT8qwPgToysQLENS1wEzqlQ16K7BLsYSj7NiKeZUegSwUwqXTIUs8G2LtXeZ8Gn
6zmGMaaGdvXv0x+drQTTwWGH+N7r1z2hF3kAs+D9A877hFwK1fBWuLYcGBjoeJ/s
HL+3a2kd5fRW7FStL7CRNLQ20j1VqKvkVKs0KGkb+C0ugkGWZIOcsCHw6PWFzo2Q
rd5p3+HeOTBZiu2M5XKSbK1gk9qL8IGjQso5tXBmcmlZEssyQU6+TADDhVIK8ZWF
b9LEgMnZ2tvMYwmi83rgxO+RBwhPxvruEi0XtPbVMmgY138FIydVR5l4MxO7SaJ3
xVPMD5gFlC6QFzc5ohcD5AKEA2Ct62llTUa+Cc69bdIRQyB8jd2RlS0M4tEH9aYz
JAd3sjq39j/awX8HpyziT51fo+PhogfeJUar1Bl2utHGP6r2oXpCfwJrTOy7iEvj
0kQcMdvmf9UtpjPShH+nF2LEuMD7bLJQbM97UKWUX4QEVVOURSaVRQZyCqWbNdsJ
gfA4QWMsdz2UzapuM7rRkWx9NqY/B8vrZCRLNzQ82IiDWCCer+ovcO48U8MYOPFy
6dQsrqEYky5bKmZjKEVt2cldr+bxy9cXj3lY1Ph7KYmZgB+O/KhGU3SGunMuRpNS
GW0u+W853moRLU3y63ug2r8sxNTMmrIpQY7MPV/ArVsnP5Qqbt/WDKrNVXts7K/v
ZEz93Sk7CuDTYKpdpBY7IQ4dfSPz8VsvnD5cTBOlj4aJ6K6MMuPqcGRoyUaiiRxA
JT4qYCMJISAXIgyNWEt9oH1k2hFnAidb8QqkELBQir6J/qY3UYuqQijIFd7Ce+Xr
AGmXANBUBWov7i9ikQbr7IEN6A6PF5f6TfH1yiQ4jU47EYzxhJN0LtXV9EwWLZJC
BQrbi3kGMp0SAFB28T9+84ApXy3pt1g3QxtM5jevTyYWShGRvWde6nzHi6PuvPJ0
74wFiTRcrEK0yfHAdhwLaXVguLXxd7881uzdQJNWEM47EJHONG50w+l8oT9ozeUt
H4EwHP1YaGkUGP39Pjo90HsZnyb4HcjACYyvEC/pEudeKRDT2Dvxh1hnVk9g5pxP
uupXuExOEql4RSOcmnzRjb6XEVVVRkK/4oy4pSEbFUcFMVfCcnQl3eIjjzdK1bfJ
RxO5Rvt4AAV9XDcAa0TTtlTUmzRggtmPvWg0BzFYqI7X95slfUX+9qoanmAlMVZp
SM7j7Avc26xxwk3i31GCT6OG8SR3yXcCAgqwe40Qv4tX7a78JfUjqQ07W+AWkXpc
zkNyw3x+MC/taYI4ydYwAEclld28MTVeA6ZTc/QmOSOMsrTp2EXzI5NEYFWE73xW
5/yHDCo2ts/0ZAA0dUXWfShP8kxuf9XTsnfBGXDQQDfLsXms9DOjwe9Ocx2vlgiH
NWpcDGBei6e9TZORTJ6abnmaa1du4KHi1S4eKKqVLphwABTFAilITc+uoOxvGLRE
LWiMZiFKZhORy924NPjmzETMCBPCjowfvoeulxJz8DSNeXsT6Jmh0byFBvH3jBmu
bOPkcwqz76+T8az7a4LvbvSDBO1b/u+vVRgTpSD/9vDhN+BBhgEKB3rq7aslHJNS
dWiz158bvgbbU50/PYiZ0+1fa3jLtlRU8MZtPs3DwntuzPMn3drBWlNYcKaWiSqV
DAfpROrO1AjXOC6YsDPiPmIS3dTXKbabK0IA4ybKNyeaMUMbhidcPcLcYmH6U3qp
aWb99+KTfEFLSmRa3VzFw6EoXjjSv7Gi8jhohkohPWQ6GivGi+Ulr2r2tG+XMqz+
LAf9/yiRQ3OFG/1GYIaDSYBiRXZvBYUCBcaLTVRYw64JL0Tr4iRZfirDQ8G9ZEBy
V0z92Ptt136pOnsZmpfLzA1bCiLRKOvj3+3j0NYT6nuMh3XFlC+jDb8mXLFWQBVE
d8iiJ1irfSCl4BNx150KsboijW+O/8xof96ZJZGUx4f5eZjIpsWb0pFCSyAQfdyf
mHemGkUOanruTcU0vYak0B6I+xBcFGXL2wpJO/CYGgyW0wOpnZknpb4blapbcCSG
iv4iI/BvBm71f7xw/Q00aypmS3zbBUxKZdQdwhg9OT/IuFcCYDdAhg53IDbncIgO
FzGfVzemqU0mQxbIUL02EnVWU8kYHcBKIYTJ48NetGm6GpT3Vvhq9RfE0+mIL/MK
fMmtwFHLh/uIwqbp4RRyBZ+A13wKwqQ9kebtgocb2mmJyvnqOVsNRmt4pURefUNU
VZEiRkQC0p5qK4EGRm3pd2GNP9A+0AzUkoIkhmoIDXvpvOCNmLhL7e6rABuWt+2X
dq4dNFg0SgUJdU0KjB1q7uoG+dB7TsokA6KCamNcA5h/DufICNBEJHBR2A/OJ/bX
miBDHWbWrTglvD144RRrKwWSS7hz3N4t2jHWTsR9QSfIdL9eu8h33rCLGDIGYYVw
/VT03CcZ1ISdl7HV3akEmNztpcDXCqMI/zWqF09772acqvmLnNAiPodShWrCqKRA
f6LGDqd0H7q34CvebQurBxSatKlZr0g+8CBX2vDKBGaoAwkzVHLd0vboYLVszJei
JUKC/KNAIttoBLNMGQxfdayCjQU1aukE73ZoI+fU4P6uYoGnKRYKoDopWOAQsy/v
z4K0NNHVIMFQhVsMoHqzRxEOyRgzMDDX3gsP/Bh6OejDRt+harCiRaL+NtojrNkH
RWnPe/oSHdY6bFdiYzP9dGbeiWPPf7IpXGkrRqMRJfYC8QX2esp83BleClYeij2R
8Z2MRMLbYKuUwS9m3GkL9BXKLXD8oNBt68vzb6neGarOGXripf+AVpoTOyWKFj/8
2mb25XhQdYNR211/hzVD29rr1EqEYNF7J1oOOuu0MGeeLe4aGcO3ImzSvMDz/b0E
Q2wwkBpzlxoJS96tiXnuoPdkW3rX10RI7Yu0LFkf7bL1NX5JmwG6kugJkHMeS0nD
Z+EzJcme84ZD6T/0AJu7eXCokpEhQv1DZ6go8RU5y3ib37x0L2oXBIyDIiZQ7ezI
STS63Z901Fw+ffxDzB20Q1j53NVBvgyNqRbuMsSX9xh6HuJayCRLoNMdtjCgagbV
VJv7fXA/mrCFKIQ45U3tmtP6zr205ObQ7xpAVfOCUyuditbZJeetArvmqOUvTZQz
60OAVx9qKIHU4DuZsQ4TtKuO/eVDAxie5vt6/LrdLuupoMJ03jifp0UG8n82SLra
8MoBM6Kj/+wblGxS5/bG7SRF4GEIojyFDtBXiItEEAyIGUqaxN1u6jPIyeXrVvGR
dabto22OEG68xYtGf6ZKcy0NmCrJ68oDLeLdCg5ef7jSNJMl127oHgFDWFU4R33h
OLoNk2dErsO0YgfCrbMLzy288WFOmeXUV3E2D0EpBjPnwkggtAEc+HjGf0QZnsBC
rdlNAwsZkq1JhsSM+x/1W5itDD453jNeXe57ai4SJtrLwZ8uWX8/+FGkpbfxdB6M
HFuy2HWJsCm93OGKVIeGr2eDnnryJ6AjQw0MsjRzRMDdFmMC4avjjfGbsYruyqeW
zQx9tmv2sWcSlk9uyjoqLC7J3XrNLIHeS2ru+g3/bMrV2M1SdXP3Yo88fx9zwayV
DPAXdvtKZOMzYbnCTPiDQ4mVckWTnYEtFgooJq85LdFSuXM/iHlhWmDK2pgP3FbR
Jy3oKTEGDOViQI7Pi7f5cofg2gxOxyCNPZVyrTvj70z2tYEJ6B6oLdaahsW0fdgf
Y9Pc7OxRj0D/yyf8x2G/CaFXrWLF/OTQCkjgrT1Y9ZldhlOSi7J0oE+mlP5nD7ns
d+y5Sy2RMx3IgvIuW7x5hvYHniPlLNdOG+WEW6AOBm/gxy4dUAV0e63W+7amiM9Y
urvPTuIFed3vpUDx/k5xpFO4QspcZzpH/eWuWs1i+ameJ8wIAGwGmeeOfF4Yd7Na
QOvhnBU5G1OoMtphLwLR6M8MnXgOX+1G0KKHmOrMvPwE/J88wjTKIF4isSUS7cjq
kDzH2q0ms1zXNEKRxiS7Usx/vXW/Eu0aTk/cMsMD22tDp3ZMIhTcx21S+LWuiu0k
OyUZlz1RVSaFMUOCfhYw7FpDgp7Rmr61+NQ41NwJhWb5hAoiDXMBzJ0MI+n1D6KO
A44zA/fmvvVtkw4n/+AoFrePI0YXTMGJUR7JZgSq4YWAmv+9T5gExyH8YeK7Pfrf
DJ7ayi20vd1jZNTNDbTbSEH3/esLDe6BYA74EfUK4+UUQpcGeeG/KcbXr6+OvA4K
4BhHJXNjlWAil/FTIUfhgmQ4bH207Ve0pCu+NI/iOt/4XgCNH98XIecprUcadm41
7Bhj0n03t/2Mxo4+rpJS1B1pEo8oP/Ug7j2uqlxsyh+KqrdmokTL9SDlFUzpBGeV
JOveSYM8B5HxNDnhVzUmcxaAxwUHoNZFaLa6vUy58pdLKy68vJClZ1CCT6h1FHKb
u1jSHVdzD6nDha2ufLia7G41C291Y+5gySvJjJukrvwDoMWnHkrq5/3tAbVQwHg/
XZLOm2VNWSrYvNFYBmg2xDx+F2K0GRjW6TcnZEDdzUkopVlzTSsc3Q/o+U+BGZAf
ebZWg7eTdD7oN/kDWSYyZPL3ipi0/lnLFs49K7dWHQ1pwWheYsOgYmyxnNiGIqxx
lV1fG+iaS8lho4T4sq4CAsYXwqUEfHzIrFQ78s7jeH/mfxgFIzjulKtIUdgSQdJh
hXpez8MpYI9ZiNdFh+HG4magXYG1vV7LbWErbWFTmhJJ4DK5/jIN799clFczTryb
HOQCwAG1cRHT3dBCI4TE0fcQjAQiR6skOP52B/vlFWDRDPHI/An4SPr8NPazKJEp
d4nJc6lQqE3t7yfFdlLInmCu3dPQ/k6G1Rek3Mc14DtuO86tzzyTYh2J6YYbhamV
oxvk0xuT9Tmk3lCIKXnSG8ZwevSZr3CUnFDhQJGa6GGLxy994UT5GvrF4bcy8j+M
hm9lyAZTsD9no+QL7Re6tr8/ENVlRb8koH5yRFZukWXYrzVcJQ115wfQj4Ty1FET
8AncsIwiYLF560khl5OmV0SF9mhS68Ixbx+fbnZeDLOdjmNc6vepDCgud5MflfjK
qmGhbU/bwgLVMw/NkbowCWSqIMtNm4UTCW592rHzfh7051F4NDu3TyHJxeUTnNn6
WZUJXws7TB/L6cvJavmBCAGkF9yz8IWaF+r/ZGdem6fk5hYwQ3ihu7ot0QebPJc/
U6iR0fo/zbsbRWN+vN/LA9RIfaFJ/gSUtYAjosgpiVZhcwSs1PEuObD05macw+Zj
ggzwBEPWj6QwRZxNBtMO931PHROZvsY3shWcQjUItp7ZhxmsnyO5W/Ft76ipl9ts
Q+MNLyyr2nyj9HEe5XzwUMtKrCTC+K/kx4jMArexmPhAGIZ+qZAIjR4JlRIoUcHf
hNQAnkEl7fSE9apvqpgAuX4aCXDw7XOrn5wRfiAT6hzlBLcy+8XNFaPG2Jx9WpnE
qusBbmBF8HsA8RYx37Bcl5YONkxtTVa6+GcB/p8WdaQdG8luH8j6WwU3DGbYJy4Q
MEMkHImkb6z6KEikGd2DxP6HpSKd95nyK1qanH3W182Me4Ne9HbILuePQ9/MK7vD
dhjk0CFryOtQ1//94VHQ6TZ1ufEwn/80uSc6/As1DwJtqky3SoNJcHc33HY0tGLS
fiF1WVY2CHMbarAJcB45tOwuing8KncBnz5yPYvAzRSU+Z6IRybARY378oY8FZHw
ac3+5jTjHIC/rHj7HtxB2vuNHJyx18LeTRajWurKD5Ktz+8kXPx6HAZ4FB4J8727
Nu0WtU5vR1pLuwsoUR5u6cmti4P5LE7ot2+mn5GHVK7VxjPOZ46O0txaF84LXkx2
aQp3Ek8bZDgAJX+/DSb7HiMOeU8ku++MLi1ecEXIMtcweS8ubUYbKTx9jz3Razvr
QyC3zJdyx4s3qk9O+DYoImMEitd5BE6o3TRAtUp+iSArkFnuLt5JlBP2rRi+8/+O
LCG10B+d9NQ0rxq1QV4gGjLUIng7ZTwyuuRi+TWZop/I4M+K7cdnBQEp8+xzHMHV
3T8Q0OZeg08kEpt5NGSk8sC+ojf84pHDyW+32pNpK6sYGxj4cfyKE1G6W4tNMFp4
duowK8/UYDn8phBvmlTC4MYN8rCvup5nd3imFm6ofVuXMCmq8bnYaq6C90P4V1q5
w1z1GQ7AWkeww9/Gg1uTKnWH+Z+z6PIL67KE7H01t3jIQOUahu/Uhs66dVbeIlfm
9YcLbX2/8mMAVDRjqDBP0Q48X0frAPSo7NV1LB8kYuxCXIxlmA1qJ5sK0IIz99i3
3SqTjiuneLfxUeXiZu63SNLriPP9fDLmQOvpvr/hHSGIf7Yl0Qet80FIKmqqRgVx
7F5fCnxKW3UzDwNhUF2U0YTmzhd4ybDUFq6QGcGxaU3GInkLz70qAuxeP2Ldtj+N
eJ4zkmK+4u5Z5vEFCZ9URZdt6OwrJXWMSlj+bdn5pRRiW/hqT6aQzjup6KoTBM+f
t4Pgw+giGMh13Pl2H2ErsofhyOyXa0+Mx9OONEkz44qCvxb8AmqCNujcKVuLxn/P
LiLi79I7F5ctpLrprJ7ZzrM7V6Vl33gEKLAZeh1Pc4kpyopqD3XdLFDBWVVUgXjy
W8LPttWCJof9yLqfzFjFy2g9i/4G1D3Y5B2EHsWhi4rJlHMKeP0YgJuBuW1zBliB
gOF2ZDa0dfjcVsS10diTfI/7JAd5SofktFxwvTD7bm/Wd3fl73lGna15Nh4yTTaq
fSdidgZtxfE7ZtnAPObEdnzTbfNlEdX+5eb2Z8JQTfUrbcXfGQ4WaO4zrLcbAS1x
z29p5tYB4pgOyohHszeI5JpmtTrpg8UN02EQJPq+OeQU4Z1PbCLLLi172f5sMOaV
s7eGDVHGrn2sN3TQ35SmbymoWN6MZ3rT+ae3SMWBvvJycZoysIqhgjt9qzUTp9L4
8+JzterwalVqodeA/MR2B2ekvAvrAR3LjG2g/YJpv7//PNPk2O/zBgyjuW4urzfA
twpD3SII4p7ye9p9AUWER1FBcEvKeQalX8RTga0xhVFTMPMhMXa6bGiT+9YM2ptR
i++ddE7LrkMN3LItOWa7u3o6NWP2vQrRj9XZjlTRIp/5ufQ5scywTcvYXp3pVfRj
FZbtj+veRzzmAqpr1kyjDA/QMNAOMwO5dtTQu1hexagD2WZWmgTuqEAv8mDZ3WrB
w69vcFsa//DmLNF44eM+BpXr29+Or6H1COaEKMYf6S/GRRj0mh2ynSNMvL6qqjci
jKN/zUHf2s9FYP5oRNOgiIwKsiSzS7A3zMPorThE75bHNJ/MObL+hVrdclVpLCES
98UAqWWrH8ZqE6K2pEN9EPM74iIgXcB40o0KUQYGyXtYsgllqCHudE86jsqsnxif
+kq1NN6vm0qmkjqzvJBmYVgbWU+7EIwvO6mFJ/EaUtNWijtyuC6WnMCMrunZ5crU
vZ+C3G9qTf/nbg4KT6038wnHHOpoCDMYLGd0OAuw2Oi1HAHLO9q6+oXmmguonjJg
umyD0/tvv495vLRLXGmXmGK75RTA9lB44wpOi67kThSfNklwMdEfRLs9hwR1Fhgu
6DQV8EmRSKq0wUcKtqzoICmLPbOB4TVgTmJQGZC9KyDxsSRj0IvUuEO5O+soam7t
PzOaBH7fUxy2QnllTswL8uGsbAkwKDbNVAL56jfmWGhHVmHjBaeYvUePLJPYQvC3
2+4PG+2eW+V0qINcZ7901iVbpF1anjLJZBy8gw6eoWIFtY0TZPT+2FcHzT1scSHh
WkGUp4++zS+h3UqvGo75BGyRtV/g32A8dVKJzsB1a+OcaoJ48c04DkPYWmYY+cTN
ZGiZVb8fA2uZjW3cBRsWlTauHBSMYL4qd6Uid06aKenKixBcYbPsnGTyNGhOcKsm
X1js+Yj3dGWNI/TPNzOu2EF9GEFcIUa9yqmwvzEQSJ+9rjBaaArgO5QXtlL97Bsy
PL/retvr8emSKdYYxDyrU0xZzOd2SoLSD4iy4DvSXFjsCcU15FTI0sOjZcW4onIK
LUxV5QJoQZwZmfROU4VoS2w0882p/UAg7lwVC7UOYFC55Ct7ZA39JCAcPXkmjlMO
LMimU/zTJJ3g7yPqJPV7nuYZl0pudxNfO7uiz/lsbkgIWYasj8GqXjV9QHT8yYAN
GWy8wyQuTpoQ4w2DlhsGKrS+4GXYpAA1tZTXplBWFPJ5B8Mz8R2wgyU5u9wZCN/+
qiOsDwQwCsTZ6JdGqLe1wL3dtp4RbeaIrEU9+eAKAybDnmwgQ9rncX5YBwW+VRQz
HGr7gmcdjw77YvvbXiCFMg69k5RwAW/IE2T9MzgCocR6gwsVwW90D5gk+jYpHhpT
6o2An7te5UzxvI+LctdEcFfAnbrJWe/jL4tOaDfBFmmftrB6hx/RT5WdWQvIZR14
u+V5y73aEKN7ormYhI5rL7j2GjGmLtuc5OgG+On9HaP7BtJm0+VgPBI1slUZ3rzM
+rYOo3OvvOnrRouXah2hx4sD4PgcOPRwVnKvl0dT19+cTnyXDS9bwaQh2ds4/8WY
xK5JfUhvpD73jsqjuyLJVsVQ0FeU89+9EnZ/i74MG1L6L56sjOTG/BOwQQYTGuYm
iQECWbkQ9dOZ0jT9Sjf0VbWDvkOYWQ4afqldtbf9YhOYCMCkgKK9JEfTY6QSA6Ql
D9xNI9Rs+Vrh0mNDtg9+PkyMmdx9flemR1s5ql0Sf1XtLWA7C/QbygU4EZ7jlkY2
05fCq6IA64Sah9UbBvmB94YcXcRf394GntUNirEqerMj+WZJv6gmWuH1NpShPbY5
/Z2rWB66n8SsoDEYAKcJvUyzLaJR1B+Z3zn7s3exf3D0lu1D9y3W6E5uO2pUUURy
iiLfBgzReF3h6yZ0zDhpkacV1s1Tq47H/Sm0tNjqy6GET1Eg5Q1vYT+5U3xzwSa0
1LDECLGnZoTnCHAoblLFdDh2E6q0L7JQXDwlkv8XSrA2zXwgmk/ZI7rV1IcNc3ma
nn42TC4IhqXmV7VIdjHjQ+9y3FFyhWsJV4QcP4s6T25ytSgYhtgSI2fuFx6Z4mUS
ep5YK5PxW4J36/eOScZiPqrWxFGrrOeKQGQrLirB9xbfsEpeCBkV3OueKeshae5h
L1SICo2zufrpWM7ZIgjXKz+rMk6/hbRlpKouWfOGC93IY0njLWxLeO8j4cMQ0pmN
xzHxR2jV8mZ03mPN1AB3CCdkbZLYcBD/Jq0kY/uIAaCrPJWnz9Q860aBGgytrVl3
1z9IskhED5dGBbq4E8aQDvDKm8rWxl6vh3K3lftTpjz7wvNOmByRkpzivToROeHo
d00xJK1YF1jEzyAuWpW91pQXclOPtFTZSlWjZaqUO1qFdgjbU0gMMZMHRGEq7QOw
VmIaQCqOyVrPxo+gNvWuD1gvQ/YeSCZmRMVDhsi72K56BvjuhZ1NQRP4hcqkZl2s
5S62WexdWiVwryPpm7JU1kf8v6BKvc9WC+aWJScNehR7Z7gt1sRnPs56e+HkF5R4
W4qktxF+miBjxY2rAVi0Od8k3F1XtdWCMImSTDbbo1TBPu/IHuFYHORk1uph/Lpj
3ebcUd9JNcph8TVEclyIa+L4Ad4Q6kR5X1JSMQ5jjKLEM1+iTJkzQw2cszGlFp9u
wyVKA01bP0UCDfe1y+VVzF8KLC3RrJUC947a9t+7W77JuQGIt4KZ4jrF4JTVJcC+
R/8OazFeso9nVtgNu3guJbr3VXg8WhepWmG/IHqeNGxipPSbWvbVYd0FNl/Pa8kn
vepfo1INHO/tcLQe6vOhQFM9Seloyx6j0DvLBCy2QWNLe49+ap609Mz69p+4gzfi
IH3qE8D+HbX8doiAe/XI3xWWqXrNAOhCCrn8A5A073FpAK9yarasg8W3Gl0axD4Q
f3oJgqyQwtBh9JBz7MPRhGuVzSbQPBOJMf3VFOTlDmZxpbZ7BBbNZzBBiX5WEXz+
fWm4Fs8GX7ZnsMNBnvAaCZu8CYfMsSzFE9VaVK1VpTXay0ftlxwWvdA1Rg+32kr8
H2d1KedEI5XAKAJvgIy8Q8sb5gSMYMWb0lIuWjLm0GZN8h0Ua0fWRzcwc1SCapHp
Z+LX6zA/shXW33k1OJYmlszUImMY2ilfljjMhblCE0UkHftdSG5wIJl8FX9/NMts
ZDkdeVMPbssiagTSnBIp0nz7xrHbuftPmz3u0njpq+/E1vjdbq6TAo6vffE9+LRS
xucBOI5DHvbPe2J8znVoyEXb2x3uCEV+DMuEgnuIsXH48xUEclaXtU9IX8aPsrOc
Ad4Q6rQP8Y5SsUCrzSX3E5CtTUDfOQi2gPshYPjLeK3F40rmBGa+f8hhNim/u0HM
ytf7oV/SXb/7wPqlpiAQtM+L/+C5apdK3Y0Aj2V5SqwJFV0JPErcWLID/uzNsYs9
cJPkMQi24GOtLYezeoxJV+OEyHN48jnds6AtilIQIqZcRdVSL5+nBQisFEBkss1t
JPa04NBZ/vG5aF62K4jLmJ1hPA3NxQ3Ie8nDZqkBfjWwrUHuiwPa1UIO5T0klwyh
V945NtvIVVKlIiV2w+LHHdRAhGOmWCDbqpEGOh+w/xd296FR51z9+XsXcGPmkYws
Mi/ntiC+0ZycCWmvyFfAYsxHAXZLFviCaDjs985c3QaOh+OpJ/nIaWH2bPCQOQeA
rtJgjRoAyNKHGSpocQIckRV1O7dgYzxj01Mh1V3rvr87Qna23mqwbNcKXpnRY0OR
vLbzhAwVyTtyngxIJj2Ss4uV4jCaCbnkpBRZDBmunOXCNUiwCgNvOwUqTGzf6HXl
eD2ZwEe4roq1aI1pHxyJlP2UHrDlC360Bs6fNSP8KxPB8h7+D7HUKvqygZx0Q5Qf
bgo+xiPDvuB14qTjjktRnoTfGFUIeTxvNA8pv2CGMlYRJyapE7pZFTEyrCEdEElb
+FlcvWcKQ/5p70gc4kbdUaoFX7kAnMgJxSOnSGU7X77j4UaWu3aWGWctf3r8qX1C
hW5Fl2wdCK5jgLC7TrQjfBGHus52OBg/12LXjiXE+YT08GG1AITieIBU5h6Mq9Fm
liANpFVbEReXNNWxlNZzfst8ud2D44I7qdqpTcgFesuPUV/GslDnOgaTPZkUBzkS
0m7LcVeuKNe1aM/TS7rnW8oqJkbvIBmDmKg9dmdRLjABYbkNFLEzxMqTspkSxyHs
aOeRh1P4Mjcae1jYHoiN4CkZLVkJiJX4FsJHZmrHyglAzBIQJK9kMiHwUYxyuZgI
IDqUc8S8QwL4yWJnNE4mFWulOuuhn4R/XFlwXzR2iekYi/2LaXnG6c9KPg2oW8vV
COQvE1wv3J9Y4RVqzAWjE9lYGGNU4IriYA4S2oYouMmnn0LKVit0i03ybSFsER3q
Dcg0XNew/DV9BocU52X5AJ/a+DTYzxSvc+7l83cg1FX5iHagNSFWSxXDWsUgf1WQ
02nvo3m+EcA24u48KzRtPQQ9MQeQWuZX1KK7fHoqFhcbvvxIiLgoStAo1nWEWDrs
QCPFer7fy/3SzerC6sASedDoSmMosbFmThG9GVxVu9g6pjIhJhkyCpzEkE3McALm
Jz/rCxq1evkaPGX/U27FEIYuNaIEJYxQ0O+j8laJnFiYgBkcoaUAUTWmgRR64hAh
bNo/fyrPtg5XEpVs0Oj7JrRkTGV6fJ340avKLgJWJZCbKbHUPQfoAH7jktCh5TKF
G5DimUaDmARmhgioThJl8vpuNxa1DVfQg5OM717VIci/S79QVaGbfAuM/pRaA1K9
E2Y3VoiQtTM8kOk4kFuf00oNJLcaoDhyw8KLamg7WN0CHqHlJPUPxHKn2vVt+cV/
h2Fsij98LWaDaBKaP28WdS6pMB45sTDz+9TU61Ikg7J4f8V/aoiqsezqaiUm6rI/
dnOSwtwrQpPhDs0jDSw/pJDwV7ruP1Tfy6v1SwetdlfPGJsRGUtpf22Wh5B6y9x2
nKrMTT+cwR5Z/S8X/ct0oFr0KvyCg6DxeIwc2X13/pD4HCpNwUYRRR1R/2a7TB2x
5JG+kuevJ/G6gFiK7tqIuybYNUpW59sD6111nQAMqdTtQnXsjMxJNUR5AoZ+YYKE
wO1PSDJHxqRc+Ceutfe6U6Rdpgfy1NR3OsXGqEpixUM+pkzKaBTeXJL19pHKm9du
FgtgTD9fsYKyUtC0c8tImLLEZYxtivfudHV3llnkKrjyWtjoE/malw38yjQL26ei
KQGjenICt2yJcmnU+p4FIl20tZVsAdfnuaQBd54Hna2bpSLpECejnA7yZfQKldWi
/iKgGJRX0M2J66/vH132lVWZgHl5ih1+D0Tu+F41s9oLDsIgyfIroD2fqEPl6p7b
59dinNi/Lpq750lCpfOYOPRgcTeFmC9b0czFj19jdleaizs9lNyzN81acAt+dQkm
+348N7RAF9GP81QT/yFsHm1/wjsKl3PQw1KicncPOItkUCwiNNj+RLksqmYksFWu
xFylTsgJfOe3AeAw4bsXzhTzx1Pq6WFedW+PHxYuEjbli50z+W0/NmdgbCXjqUch
nzlJQNla5CJiw6OwnA6Z7Sqb4kxsdA8BVH7gdMkTuMIhCJXpcvTpBMk/+Vr/r/qx
3p7kKPh1C2PjvFZDt77SWzQwUbuHVZ4u3dksEOE9hgZDa0FKcgteyaUAV0s14PIX
AQHiCJFvXaDsWcvx/dEfhpy+cTLAANr6XpTNYxLB4Dkq5MgAoXTzwWijvl/nodMU
i10JPZZxR2Xkna6bGOdHL3tuemSKtwaoHvV+jVqMq3QDUsELwcnd1i18cK2I+3Zr
0A9FR89a5E0jgt0J3y2oDMfrIjmHGJQWHnfW8x6+fTpxtBGvmFUta8SskTDGbJF/
sz10i8jLA/lh3FZhSgLu+fEZ8jAcGmxBXMByKs4QtI4TRfsyz+KzX+yiWkvOwvze
OR75fvcKha2xjxC9wUu5EZEcp5MmCACxGcF3xYaLDhmTvAb7SkjiyHshCJ/z/Zwx
4kz6GUnijo/RYyCm9W4KZidJ6QhxnsnIHD5LXECrpVtk1PMVqRMInidEy4220RJQ
rzSkxL4pe2BuWUVp+wTbu0eOwjXTk4cUIaLGSHKtjMR0OaETtN2Z7zSgzJTuYzXY
8diHUZC2cjfAx7ABYmsC6dttezweB3DkCR86ldepR3IKalBI7PKXEA3Lr/E1jRUm
vkIPJa54bsV+HLVTbf8YDNCsY4JB57yMKUvaXSGxJgBLn8TMpXJvJOoyKTvZQs7F
d1TXkXyTnKwPv5H6reQY5noskuDeBvJBLGlM81yZ05R+XiLyotj7aemiClsCQ2lg
U+E0+lu4u1etbUsMB8dc2VjNEaXqRdPcYoI8z7CODhTDfwPwFvAFaN0V2HpEBVYH
G9t6u8u7vSixBm4dRFcDTAfS2POZnTj9He9jMKnpBnaWQYbupXgb6wtbmqv2oR5i
IbA5b0/FDsUR+JvRr06wgXMX4h44TCgov4vEQobtomFD0CuYTIcDy52wXLtFZik3
qBczdKNFIlYKmYysEnPqY1O13ZmqOggWLwGNM6QFeTwb2Lk6WKJHZf6laNK59j1o
JUqdhHQc3atMepH6TUYBKaSzd1U51CiAwzrxcPlRf/MrnETdHk8xEcmFf8PJLpVt
9vnBlmvYUJXsW7MhGxs2v5ShnqA2yRKEL25vS9CrFlLMbO7raFL4etPRfA/nM8xl
3cE+SYJb7kkWr7C6Vv/Yp1S0gXiIpTA47j6gJvpT4U5M7kBwbkaUMzuU+jaJJFER
nmRwjfXBte+wAMs1eqlMSQzWf3BmxesW1fX5Tufvsgvdk1zBNsD2TtNpDp7hjdGO
hjZ4fB5SXvAmusIyVfB7/CGFj/X2eS8w/P37KYbvq7FaI3ch82GMU8cKOQQewodW
a938nPgE5KO+oBTglsH4nOFsEfG0FEy/LuhnADW5KzkiyJydVTSL9NOv0PrvkD0p
GMsqnZpMfMD72SA6vHsiic0CGDGPHwR+Ra5GzHDcXomgMYi1gc4y09tVvqBbY49F
QeEYMxBQuIpXyop1sVuz5/+XkWyv7b6UwWJB7iEKsXue6+22y2TJdXFmi1VyNzP9
4pu/L4dbzVRCpup//ru7cu0i1tNgiMK9JQZaHCwaa33ix/lrXyakXfo+/+af3fyb
oVqs/640kXriums+S6hc5+sCzDTcL7GlCDqAad8JimOxX0cr+KKp3qM2h7/WSHaU
opO3AW4j3lv58PsSgZcUiTsID9v+sVJuA+/HuyNozdknFTkx1Z+RsqYyuJo5lrsg
fmjWtkX3LOr+SEpZQqSA9iI/rTk4XBUEX1BLFK+ywkBrCWYDBBPN83ZzO6uuT5BC
HMbaF76W5hHNRmmuHOHecUAPKvCeFfwQXqN1ZpxKDcjdwWAtAcU1iCSx+PEuUnnI
9gsCSYvxrxEp3bGs7LEPnNs+OQU+wNhNJ62x/GmUZRr/0KlmFqENTwsNWAGnDWu1
GnmMv4SfGubuCxNbGjohJpZRatvsPLJc8KNKK142OtEMEnCmx1yjbLNnCOzJ1NNZ
TCGa3pO5qX6lBJJodW469oonXtno16MWcJqIZpgLF0bYhsboCsTazZFXjd1bvNgV
HFaqIhfbZKX0bDjN3m6xwXSovBQljA8MFMcmEZxaJ09YufDNbqC5/tB8WZ99ils6
ELojnDr85tIHQ8E3iMfw1pQcaSLBW8SX00tue+KLEH3GRr9QmteTPay6XLa8GcAD
xKWmsUvLrvXl1Xxx6DFI8Ns0e2igAdu4HjsRoWa1LDbuO0kv5wSko6YqX+ATJ5vq
qjg2FZqto4VtOnSA5CrN02kC5ZaVnqRBjGJ4cPSXCLGWNxl8lKGDvmitr2WPC0pl
6yQnvkL2vcHe1LfqtGJVO0ow0N3iOGWHznA80dDPvNBLnVj3a+Wa2yJkLR9IGOpI
P1wagdRo4ACKYVzgbYKHb/w2rXl8rrcUWVs9qZAlL+QY3Mk51oclHr2YqcjyhL1+
oWFAqiGmH/gML4c3mqXG3oKY9EDsSGNRBzDIgGfOZizu88hWoMeeaDyDwRdtvqiq
N8utPBmkUOeum7J4qVbI/QCNJH4cdmytT6mDckN4XFlKXoEXnKXGvErD/Rt5LKay
cL0Ov/8BlFIxM7nZ656MowvWACmBL09ECM0+gOuNWOD3qCvLm/v0kmWT4cPxwbVp
lX8XOQ8CRpN3EvEZuDidywmbvLiNxwGxEFu2j52lE+gXrWgdMi0a44rFEM+/Vvud
mtQmbRKTZ898ozVXKqN+RGNuVpVo//nQQCfu0DPxvbYsN733guVTrB27MvlHG9Ox
kv4Mb9Blj4d7nHCJXZZ+z3srT0vD0BZhm5krROanaSrkDUr489JDAjaOyfh+X17q
PHQXEztn53/uMrQRQbbEILqGA/KWAI3EZRoHjydm7sPyP22FIOmU/WHEumZacwxV
easPYYxX9smslAEaNYKlzjcVIUgzkFNRTpE7uZx+voN1PX105KhCaj8ws/8m6Uqz
IqoORu3YPzByV+OHiooY2fuxzRKIZ/HI4I13e0XCEpJSyx/UlXlnQT/J07WVSvmi
GQWPYASJ6lu07AAf9rySYNp961PBI2DR6fY67oQEpEna1E5EsB4ztKAdf4QPHwgM
VWnZWq2C1fmI26TqisJam2VQEQHmGFJwKappdyYcUnpp7OaB5ic9aVJ8s17UfSVV
baHm4gSSYwX4m2MS3Fw2tWz3wN8L97XPKwlBXVIts66PIzQVq4sKWe0vAzujjnQf
fSZmyfTKXhpXp0MMDR0dP/xVO0WqD5ccRN5zwvwP84zjyyoKCIQ+sh/Q8YISTlxd
Z+o3UP9/FhC4jrHk/2QTjUlf/MnvCUjbTZnlGPLzL1epm9JKP4aTswlDfH2naxDD
iD/0AOawYnEGSRDheyzTbk61FjmT0PZmxbI5+yVT2svWw4dlrZj2sjMp8d/GVE6F
+GIJkI2osiEoPKuJTx46+KxeScrS1VzfmhcTkJPz4PSn8LmtdeEwNomviS7TDftY
Y8dLk3nId2Pms1pnIV8OPOdLHFksX6WsRSTu0KhaEP/70QDEmVXLYvU1kYf/KkyW
zk3jrBtulMH8sjAnKlmxfeuMGJC+i1rJ2cy3KyY+9ZX/TMMr3sfcNAq74ammU1qe
LbUwuBT639tj3l8Gy6hE2u95O1/5V+bZXZZa3Ja+OmxZS9f4QsAmWDGpkPeI/5Cc
0SzH0iFt4d7eY0SCm57zH/qaNoZ7QM+HeptEkItfRetYuEgkeVAKL4Vi0LlRoWoB
pCilGXlIYHM7cR5WjBnW0sbyv9BDcz+PC3aSfmBrOghA3UZCRxdQhhQi3Zeq9qi5
ryOW5ifNmQkuXU26icvfY+T2Hqv+N9y4IXwCX5yIqM28sRuywQzNCD14asTJqI9C
VpDKbgb10G/brKZFUukNhPO9Q93HrUgJu0vmb8owsHbEk1JpxAa/GAtNQJY5yzpw
bE8tY5yrHXVU2D/wl/a4Q9UeNOds8gbKy/IKTAUD/LKmaQXc9drHgYrBpqriibl/
4ZSDMo6MLYDmp8GFXzDFp26o40WU+PqeeekkCL/a8Q3kcP8gQnDUkF+aoVakmzR3
z2mL2Cgl2LPBjzf64ulbTUnCCJ5gtQSl5pcmUIDJZBwub2c4r/zdL3aWy31FY8U1
OjOMrWlmB5LBaOENjbWlQYlWWDl/LASRlgZzZbuDKqHoo1h8Whg5uUOOKnuy/euQ
elF4bF+hQ/vood/JWCzFZGIViDZH40fOMHBArGM6QH+XoV0u/wJN+HngpkVDwI2c
csKbfQu4uIpKlNvkiVbdyxNSx4V4tNeCt9g+fslS24jUxpS66KtOBOA+Qr18vAiG
NpF8i6w35Tu5GNZz2O28/KHt8zCrq0tuKlFO68Q/3WGPSdAGl3eN6dsDAO7pPcK9
MLgeOdA0a1/clKMCl/0aA2DNFQaK0VbbByfLVQ8dQsWiP4yx6hlHLEW4fx+6iI6q
kf9jqSo8IWdMkIlD62wKdOfPtBZgCZlvkKyBH32/OJ07vxW6CRZdPlc5lvB3aIPS
1l9yU3w1BC7tL0kKQoYT8LptgWANMfUujxLjIOtUA2nhqsy91vcur9SDCa7akFoW
uK0aO3E26kMmkqAinOHmme7GYATdv30EfJsnHoFWDrez+dArZjiXdClKl5n7k/00
npzZbgPJiF89pYGR0Ru4MSa8wJFodB2dYiU1zD3kb0fW89K8z4ksAgAe0Ix1/knM
wB335eKShnyLf5SyoRNUh24vTwd7Sjap6Ni9fMtA5nfA3SimxZb3WOe8WDtyvoKq
KJt/gpMlzzJyNjLjV5vE1wnnVcVc/HsSp8JXhQsgmqtlV0icei3KvER2JEnbkRyw
c7nnq4mpVdTZxieq4359WaASA0PuZw1+I+Z0w5b0goc0wggdATJZqKuk4J9Bje0C
dC4Ob6dXDZR9WOfeCrdxPp1BlCIeEbp/6b6XjwlzNUVJ/M9XArgO9X8Cbz5swfLj
swpgdWvzemhNIKf8AzSH+oCqRijECdSrW9vWyYN3I9A8ojgFuhHr2sSdbw4bnvXB
Jjn7PyayQk6FDXtruaJPgg2DN+qHHR+T87U9acSlPSXZku+hK4Ivdmi1PdUvKiEl
hSe+0V6tyk4UFQ2EF1pHtrewrZghDDJw+rx0TmnFWfq6qmeMwI2TGO8ukEx5liw0
gG2NhEujzAoZQ6pFT0jOgj+Jh/blLzIjCvc7+s4C6cS3RXmtuaM9wAZjCYLN/WbO
21BFTlsXxkHwkNpuWHiaiTwdiEOJimK1z3ae3eLrb8hFGDLU485SPhjc5o1ZFhYe
CYeQEb0HtdnLrcIXv3j0d54F1CPt1vlyMDUW3PL/tl5w+02ZnxbdTmHVsQpcbrZe
Ai6dVXZJywjPoKeunq5ch/RbeaWBxcS2PHZIFvqulqgd92HsTVvn23EKSOpmBUmz
Nx9pXfw/yuWeBO3zx/tn4oNmoK9zph0MdciixnXQBSgjO5KMmV+m01n5ss65w1vw
aTHH7u0d0NjkepeQjr97F0Gt/kwk1eiIU8eGHJxWN7SQBAAcyUqhRq+qzFgaCrgw
OAKbC3TCcMzJoUFN//9TFnYrM0bSookrGryblzB8jBY/tHO79ElnzrXVweHcIFOp
gxzMlV2BxdBmEDaftPeAU8WXzWVoDSsd2dhmpuEWqCMa3b6yGtSxWmSKNZvJ5ecu
jjoCpRH/24L7LdDWLAq2PKBXPeTzj30QHUaV+cCQM8VIO+1IXGZ6wdF6HCpfQYmi
8FEHDyeDk0gqJnkWkHJKJoTXfWM5G3agt7N6cubtx0UlOxMFHHUenSjuyIXWa3KM
LpCxVrG8z4oQJibuQQLhFzwkqEwHhl9nbTcgzEpxRxfFEDxCAZL9yKNY6IWCSvqo
lh7Tyl+91hTCdd+o1lABV79bCxMghvD0VmCARy7Wz1TMxW3ZlJ9w9D0pyjPVUydl
Bi0IRdx21XQ3jYyFv0s7KFilEGB1KVyZ7DOW4mUANnnByMU95GvTJ09o4vgBCvdd
z5F2TSg0DSx+ZP4KdyQUcLWRXHls1naHlRvA8Yq7P3Uq1j0RIhZIMGUMVAQxswiz
sPGGgStIZuI8HTTsGBisLJogO751zaFew/J/9X2UewF6G8n2j11BuKU9OLU9Bjms
mZ4mw7MkJLnzFIO9nW3zdsZfOUTRm+wj2APmW08Q98NCV2qi4UUwDtEr9Z87AeeS
WG2QBCvkFK3KGYbmmKOdm50KQsReD2eNp3q388t1uuXjYfvUttoS/7w+w2+/1t4v
VGv9Z4FbZpFtzLBt2l/1vKWjpEG/xw3e2Cj2o9/xtb7S6DVq1xfy70mHOcnsahUU
RI6a58tjhbzg5Hy/5L5oNaN30hhJUMpdCg3X3L3rUdqbvzGZKBRmuwNmEGi2eci2
oUDA9Ck2s2S84IT/EKqea/RgjVDdkXqC3rBdDgvAxOwaoPFyLBEbcwoNWRcsPy3o
MCJPv/wLlkFbKwJ3Sg1JgBQKUUNUl+tsGEgN0QsHmg64MOKYaKWcizR1Ah1Dc3KH
xc9+dcqkvbirpGAOZ2PWj6WRELPXZ6kQFFt1jSK5yuvwstNV61h/lbzQ0n8M74I9
Oy+4LwxsumXm0RIwE1cuE1VpnbNRnxO9bKz4annfQWXwjiVm9hKIp7kuuvn+b6fS
QSgwc0ZPx8NB/bmD4Ym1SYWst0ZD3Rf/ceWbLAXVhtFxTa6x4aOHMnTGM12XrO2K
rMFcn69zkJetSIUXBAREoV5E7f0brx80+5jpNp2fmo4xzapsRys/Q8CwapbVmDNz
LWL71NfaldDQ0ghc46uec6Oe3T2lo4QZN4rNA79pUZ2OsBwY8Fx2AUchPzj3KdCN
3xBjuxpGYh1W15sHeCYYueUmiKUkUTQ71ZeA58V07jM9TzpB3kCDIwXn+BfiGjX0
QoOT1ZGjvtUrMCunPrhoMFnaLr1Mx953p3P/xXlFVNYC0wzqelafkRXO2Ys50iwl
iQ6ozLM1fTgkkd6bglsos8NhP8EugwtRD7mQmlrlkhBlMrRdJygg9DIvX7d2HxzD
Gq2mtq1bZDgHTBRaUB3vSySCb+yOyNM1ms94cyPaUMdLhrjB4zgnvm856N0zAYe6
hxKeZz9PWmgoMZ2fV0kXoLm24ElVXkCxUkIE3IOzVEhZEwO5Ncrw+doVht2LQWU8
GdS7H+g47jbT5mTmvqmwXegh7uIX/r2bWqdn4LSDsQjBVeWo2J1FXjXCYEZC8K4I
rmE7nao8m5KeyYHZR54sCgbrD39mNph8Ce7TrtV69+IvzxJg7beYrynYBcXvx52M
yfp8LyW45LyLZbl6QyImNAfw+4wyT2zmKY5I+V0/NB3Z6p7nahH8yeVAtVfYkXTo
XxZ14llUZQdZmT+xu+qqsVoFTLhzLnD1IpMl492qF22v1ae67aCsGTzBUQEeyBy6
I39I5iV1gZqgyUN21pRwoFaWVdmlfhfjxqXvV/ICw+hlcBMumHtB2QSloRPIOlKk
bIQbb9aP7yx7D+Zq6hAq/qTvs32c1i9n4ihLL7Fh13SA22IwWfcYS/qRkUPC65HR
NaWbboXmrheX/tTvnRms78noXAmj4w64lLRaVQCdD2MHCl5Jf9S9ZGo6xDK17ma0
sTlsbOhY9ofzKQPM2mI750TqaSBcsokIWghKpZ9VSKPp+xvhXCYDLNmX3rR5rr/v
Xlul/hCYMvqrpYhEOWuJ4ZN8ggKfpYxh0M1f7GeU8BRimsVmaLY+1cYvt/pwd9W5
0omqjYajlpbd4byOGV50ZmdjXv9Q8z4G/9HuG/W0+hv1sQOHtR6wEcvbgDi2sPst
aXn88t9v36twazxcWHBTK86YTd4DXADxw8ikNB3BPAlAYZdri88DrYbH9089Jdo4
HyMyczLnY/vFC6T7Ms3EvqcFpHdyR8jta/vqfoMIO4ex1ZMqUdPnEYVVDFDbg8CM
17Pgtyes+FmcfCQ/XukvWnE82eqwQGqmdHKVkYtq+QMYuI1+ZgCY2mhzyu/6VBuS
XuUD7dYsZDkiYUdGWNea7yeBWMjQJnm82ESqDoiW6DmIq6VicsKLViQY7fzt9jXH
IDnWymVAUyhxuG9kNAVXDFqK3y3FmyjEvPkpkPznV4D309vpfUAyUmB7YqawphjY
LDj4RuJ689YXfao2rBoR+PlV4Dnup+WYqU14ndyUsZJX52/a51zxMQ2G4D75Vuqn
RL5HwVBvzPiSDJBROcRt8uUOwX0spWrhgAzCA8tKICdGkwxJ/Z9Mz0YLnaDLvOqQ
yAiziAVdFIO8pRawVZanvWHAUuupEsHQbcMLTBkZcwt1ZOXuXyKLVcpmA0hOL3tN
+cJwE54d+sLyrEoG9QJC+Zk0bjfrpM4ITZrVO8wwnAUPYKia8QyfAqvf32vU8cDA
niSxIAMIUFDRwX9xoDyv4mPpfnZpat0duBoMR6gJdRjaNYwm6H7q/Gty1ANbf4mx
jDvZy9HlswcRbRvvIRE65XvfNhFcqPoUCFz6fAfqUxz6K6A44ZpqGF2HccpoBJbn
/Bo2GTpyNaMW6CNWr5d3kxGtsP0HYDkSFb4DgmveF+3lg8XFNE+yKZo276MIhk9Q
Qis+0Hw/F4SEncAACQvoVeq/qMHHjJ0aXg/RYqr9gHLFR/lE637BqvWgY64LEQVD
0asULyx8yyx58ikngo9w3Yl5oG6NJuXqt2zMiV0dOQIizZ8CWJ1LZcfzoYSE4+kL
XT6wDf1XWkhgnw7ULuQ2pQmNDBrIgSAE4sMnlRDf+pW8Zucy4VVRYcBCKKnF9LYz
pjuf/YTDj23FqZlHdqfGbMW9GJ/4NmHjdS4GarRwI1FioE2TL1GWi6gFN+J7+aWo
WyNEzwinZznOxNCf00ALLwhkRjWsZ3FmZ/bjLmyvuB5kktd0m8ZR+UyiifoqHEE3
SC2dMPjvTVLcVxrfN0fcMkYQcdH6bEHbs4R8gRhRZmE2lPR3cHou8TvGWH+qRJ1X
Mf3ukkellBLpoPfRoVGzGBpDHdZmduc0m/mr55FdEEbf+zSAXMVpPmgzQhpomtFC
gyBMM5HBH3qUnV5DOoMGkLYt6/puh0PSpWShpBCoa7I5Mapn59sXesGpYQiATfBY
vn5n3ExOh7BwOhL0Hd3/n5mvgVn+E7iNpcOCYpZvL6xRzUP/sbSegeAcwlbx/3Gu
BZ1tsBHShU8bmGSdsJcqqatBQkorpaSdOFPMiaXbaKr/WZAE5b8b3QlBA0OfHRgV
MA20ovA+NJ4akGM05n1w86f6wJwsJw5esvaYGI2lQ1/ls3LVXzly5bIGb6qiyZ/9
DXIoxbcGGlZwvFcQGPB7hn3XJUXGka1y2XXz4LuToyazDenHfntH0UzBCKDwo5ev
ZJ+HFtAiqFSeMId6AMJQNG7uHL+AvbtYxn7OT5k9bKp/VUwpLikKmuKuvktkmcLw
ll2YV2ruXL4hkKHhsnRi6kTHU55MctaO9ugYUKPpb55CChjCD6DgbK20BcmMZ1hw
kT7uzbf8TwKydr0YMdkrTzVvhqBIGOx11Zn+MgQ0VFOkA6x3zRLMTrukZN+SFgeg
hmomG02Rs2nGFfOXAYe14iV4R0Pv97hM7+PVQnR9gra6LZrP3Elu0p/2kqEQVzDq
+ke98dgs8TXhbnlpg9qYQ5S7AxsB7GjBAm27izRsaFAmjpQesdwrp3VTJ0Ne65az
87d1p+idUcZ+kgTxg4H8RWlblkUN+bp/eP6w58nWYOl/UsqqJDmoeYMS8VHflThR
9tni9YOJbISw224uGpaIiDRODGa49PIq0F//S4fSF75GrdcpqDGvrQpEQT96RXWl
7DPcpGfG72YsYw+uKq/F+PciKCeGDEAW1em5HdC1i2Qe/IJhFx/zoiW3LkHsDZIU
FgCOaX0b0sqbeZO2w84FdngpFuiRBgdJC+SLdZYm/h0IgJFWZsqsQGmfE1Zs073J
yfkOdVB8x+KiTQaoiGLguzaBZB0gEzXlHIILx5TdYKTHhsfT1wSDgYJqwGrC+AvK
y/F48k9/vNHYgWA4pvzfltmNnLrCXcW/FWmeJPCzngAgbQvhMvpUOcnCHBpRE76Y
iDjLIg77FTk1mKeJHJ/B28NGGTn8HvWZlvUG3751Du3UPrnTeMLpNzVf5FJ3FGDw
nJa9QL0DB9Qo36cljveApyfj5nXRbOh8sWB/CxU7mK/VKZ3irGHT6DiJeTmSgcj2
2TIM7Xmmf62j0A+atHMrcFztLa9cPHJL+zbMJnCTCi1SZ68/kD/hshRRygPwtDAi
PkGggMDYfJg2cGpTra7Zkr69haeE4Jp9YoNMmiFNqqGaQlHuGq/lqbVqoPW2trFX
SvSz6Dtq5NiUSe3AE8W/cLwR+pc6HD2uqjLt2olu4GtbVNIonVV7vIjF2FE41W2R
80aAIY5Rky9T+xlieksfF5KfKYDL4MsKrA0CpRvMiSJf2i0Lfft+MStpjUOuMN9T
d26q4qL/gG20Ic27OCQeg+inMNn+4EEirkzBhoRNXm+NHcW+PhaVdpcYET3aLFzc
UzbITukH9kO/+z1+qEABQZwtSFi5QdnB917FH+X/Y+uH3pUCCtoU+hhQy+mqnt7V
lFDVr4trpStRl3kX6RfFupvCXzGK2kvyPNDxbZO/clv5JbQ0L6kk8HVDNT4FrY/B
eczbO55w8ccilfdrwnHw8VcP8/e1qYP7BDKzubbD/dcO3YbFb+fdl6umTSVMn0J/
ptBhSNyXdk1lZsL7JEckkoqaQcX44BCxLdfNz9ILaEJnDGBlKTtUR9Jy3o7fffuV
Dp9gUg4AL0RB94GxbHnjc7VJJwxf4fdV/dvcjLXogTXh2XYqkT4uEfSAp9vrh73h
gLKmJETa+J7YZUPsnHg3UWyfnpI7N/JQ/0MdQHLbd/J5WCpxNb3Rk10zM0DcXaE2
yO2rzIcvhtvHnbtPWmzyaDc9RoC22AKwy14fR+g2v3BRE49Z5vzE7H54Ln5hPO/Y
bGIYFmf8CIanyO1uUoO5M4XvrYD62Yf2ixLNZvXLrd7IgYlqkEWprv/z7v4sDk4n
jHz79v1tcM1X3TIRbLeMdUEAGPC4d4p5dV4Z80UEvDX3zwGOjFoEmgK5V0J0cN6S
44Yf/NaFzOTD6gDEDk6xgZ9V1G4GzOA6jD1ZWytJxU10qE1z5oOw/7iKjY4VQJLg
+pE5UuIxSnvAFSknhXQxDFqIkLlT7JT1hbi5rOluBY3y4YI2pqmyL+Clj3mQ8piv
rMATMplPk7xyDiqfELEX0iSdzkr2I8lG0c6n7oPesL08/F9EBARBvv4lBETaqY2y
csxjBD64x9EHh8xwT7jSj4LvfI8ZqKrDZS0FuFQhXD02vW7zeOA9klcnop7tVnS5
/+dKALAhrAKCh9A8r1HXjJyChu1U3EXSgmkyec2zMkHzjj4N2HMdGLHyxSXYIncv
MydwkAdWzxw4g+IDasctAHdf7dVJim1g25+vAYbzMRqCOAYPuJ+vkuQfo120yJJQ
8Dnfm3jfyJ0MwGT8nNHl8iCkZPf/DPck3GXztfMBonY8wgw0bkbLt8QlQg/EUUu2
Cg8uXE/3Dpx81ONEiO095+2Jm+axSqHrvjFwzKDd+38H3xp7RkLmc/9rIMTTJVIk
adDNTx/yB004Avz9KA7L4BWmdpaVsCY+fdIZgIVJRqtXvpSrEEqzKIX4Wu1477IO
9xNqfZXUKw4pWbvIbB5E1H4WPSJ8zH9SJuT5ZvEdQ8uSBP72c1f5VATtoc28ovDn
RHGXamxUQ/JknWRLVCYWAQdVpvS8iaolZUloZ+5jLUaiEitp2W79CUCIqmmMNNEe
m8QHErhl5EHkencEnc5fO5o5udoG0G68lw851nLMNLR5k+qEzof4ww3y2A4f79q/
NNwlyTLqLbcFjLW21/sWQdD/eVrm90OGG/Hsep5M2SgQshTVllKiQEkrwpJu/C4Y
kDGKW+gM+RCUNnrQf4Jwik5I3vlmpA58EXrOJK5ddcTd6Ofl4Jww12urlKulNVX8
iKlogOjemFXRIlzWtI8EsUDFtyc51WE+P9jtlbd7z2JPN5vLiqlnJDbgSbgqX2dU
jbzRcvpYtRdSUGjLfcinTRa8hx5sSOBrgemnlvMo1O79OdqLtaNeqYKhDDRQ2S4e
FMSokq+dI5rdU4lzIyJj1N+dY0qK1CoaIIx+iTzh7jQsregp0a2vUXYjIIbHgWYR
iAx3TpOd72URslIHS4Sx8J7POs2MezSBKLQKpam4TTXpl7ptjxT5IYghmrLmKI+K
JACINiNfEp6qlgYpbdbtxJSOa59n1+Ljp7LQcp1ZCmTnU+OQXii6MlXj7BzitPJU
u5kM0y0NPMXDiISICmSK+vwicFC0iqHyxot4VD87B+u0bOT3Y527HkIGrVyqtQdP
k+oWoXUf2NiH6DR9fN2Nga+b3n3cifb7zW8slbVA321yLDGkQPIsQygd+0uJJDB+
D7yvTkMotgOuu4diyciqAUSUPc3pDABV7gpgll3Cnp1YCZt9tOarxuEy8sm2SpF6
EsKkDrFeBujYo99yGqRn4Wds9KaJJwxtURZeIO/ejti5UuiuHAkqnrYUK1LGYky3
5hA3GO4FTMd/0TcWovJ+AnaG9tXbAhwyzrpK6hg7HFr2LyYjuE0A2nrNsfKoJYQa
t80sgpu+z0retaZoy/wurefgcm4kshJh8ecZ9eE2W5eMC15mhzZHtrAs3USr/rKc
8is5WI24FlmMRHcaF/S0v707kpFiCHh0XoPyOgD5m855FU+YwQUO/vTSBYD70F4A
rSJEBTOC8/aWu3OcxTo+3aCPvkYATdAMwRXRV9RLr9YrXek/RKqjRpWyBxP8cNOR
gxVEgNsKFKbJJLKgtRIIu0nayAIejNYWxTiXb2Bwv6NPwYyjb/cRZeX36eTHnDXp
fcQxCOl7CI+/avDIZ5/HvKnUWyH9Way9rgTtcZxREaN4h63SIqB/Qu7ztUhcD/kC
ogCWni0la9JkTXTnU9GAFJlZqFoVR+PwYHIULLx4baTAxOdbBGpX3gVC2MrzMC2N
WeOl8jdKbePUduftJY72MxH1qMQzzdnnJKFNgb+BVozASvRgROGgclW9Qa2WZYEl
nxS2AIo0FbSgjEE7zCLMvbMJpBf8DgamP8ZPo3CMPd5B+KWgA/BICKHwz62KBwha
h88NIX84u56m4Dg1E/opaVDTmvJJ98D0sJbKE5AOYiOAhjcYi1ofGdXWs6jkuXZk
C2K5bgsRlPsf9ynHEAmbZsG4EWGPOJCYP5+rv64f601VNaxiUo8mf3P4D4w1Jxl0
VT/dQCmHpEKcyu5dIs8u9bYE8NthMyVOxIDDkzFBG94L7fAriZTehFbTc6OpzZME
UE5tJNck6mTkt2tS7EaZiU+mdw4e8SfqZrGUgGSABfl9wNDB9xVFxFRgFkANKReP
mpBYTBfdpnASfTObZaOTDGfPyNyH/AUvykmezID6MZAr0Hw+v50pnwosn4QcJkRG
8KXFQYdNjUoUatpU95OINCnDMIfvzu9mq5dEiVwOAHm90uKEX1i57D3QX4jR27vG
TiXi5SJpy5KLR84Dtv8r/PrqTXT4LMVAqz5SyKOuG1+yg4zbdWFlEoWvLrROh6MX
axDgKV6WP19CxIsByv2ZkfGLRgNNkHeQgYBsbn4O3l3J9k6ghn8yRPZ9HmDGDl7i
RW3/ZuOYQFuaU0153gfwR2+ratZsI4tMCFfXdv4AIkqoLNDMmJQdpNQt96hPB56s
6k86qPDFGBRapMTq5TzzfubHGo19G4CLr2euJj2f9enqb49wZBhdtnFfg7qd0KMm
8/vG533qbTNIDKB3bDhSV5VbIUGDqa06qdcaLTB5uabLyU9iXlOyALvPMdUjX9Up
Xr0HZl8FaSAtrx6Ejp9MlwgJPMSFsA7Ggi70joeCb9bXK/wHStHYfQoFt4mgHzuY
Vn2OnTS3j8BiLGaK+MFlNeaBpo4m4oZpjrSPd3UW53y38KhaJJB1NcOVtMFXuwEG
qRSKydpxVRpc1y14c5TEjiAkVdjLSJHHkI4i+o66UE/kGML/T7NGGpb6ZW9QTiQW
c0HTvIOAVunhmxjzoXwgndQkNsBurpT7n2WjFGeS97cNoVFqhkxoZTD5ddFhitw4
k8lUbQHk8EbGH6VohfqYv4TJbj6P6mcsinvKCOmgpwv3tpRqFHplu1v4Ru2XL+Xw
v8BZcg0UhUPVumE0uI37pLQ0exDJXBH24KoPHOAcSN3Xqc/XcJ946+KkNmiUHMXZ
WQb32hnHLctGFx3ZIHQtS86uOd6X+PkjsJQ9dgU5sBQDf44frQhC4CEqyq8RqXTP
QWKia09K7UIMyrKmiuAMyQyKj4aJEZWp1dYlAtlz7UA7NfW6eG/5XJ0vhp/C+Qtw
nOvTKT278jUFWHCDHu1k42YGVz0le6jdEg4a0EzeOcoYiZfDxwW+qnHkSieDDZGr
miaOFjqeaEhKkN8++1OIb3wE7oW22BSmnCuXXSuCWwJaWWUkHDZJLI/k26fPKOH5
NxCzBl0TaHVEmAMw5N8iOfgaSdqo5P7j52auxnzIx0Xq9B1RCgiDS+ECYvXGYNsa
ZQNApdBMwQ0pLOVSJ70Iye6aPxx5iEgsb94rh+UQ7p3aTdRzejIw5JqCtfi3Fj+w
u/ZhDdI6skpxa8O5+mr5SGZHodJz764RqUbdRJPSiwZzLeuxO/06NTZz4QyayDFB
+CZmRrYdJ1OcVDw6oO3YrVTjuj4XvwquafOLcJQjpRV+zgdqY/AR5F6VyU36Vrbu
t27GOefE8jov3CBveO2uERN1dtW/41LcUM/0C5wDENynnv0nxbSbWTci0x8mSDnh
OWVyWCoZ+F2ldiyTdRy5R16Rl4HkBKtnjHoAbSG9XteUqEb5i/6mrn90EDVpSKGb
oE02okveJHy8xZ8/nOXXuf6sBS71sy4uRz0HYr3KT0di4Cp4HkjTgCiubmEh1bs7
dkKEa+bSXSlL+YsOuMY8GnVvD7Xb42O9OQVtwMmoa2N8JNWrbFOQ4htWrG/NncQp
BjjpguWMyNPfjLHCnXyD/Q+O74O1avxSuvZ6EHmJrBvTs5AJ4zNzIrjVZfn0gD0g
71RCRkfc2KGgOs4Fl0Ss7vQVYJU4irWdHjaDxZlEV1e8/G+Z+qR9sRC97SyIFjMV
yRYJAMnk2h0KWdox3eRujOtpneycCwBlBNMLJFvMtG+ypqJrhE8WzC2VF/OXBYx+
hLbrNvey/R0GEHbuZ3CtKwbkcgRQ3In2ZrTCXBNBE7GZBdPqYt2ZE0cI/65HwnkD
KemRBNfrVoLwzsmQGaNxuVIo94UsEqII9ONYN66c2TksITrQBX5vqR/gUQhuyQuH
0f/u5kYlOYLf9dP9URFFLcrZi0IMvWHGkqMDljA98JZ9YpT2zPMfBKXg/m/VfKt4
A0Z1s+2TImipdHF6miavbBuJgkFHD4BMG4RADNJO7nrmRLI3JInsze2PtqPo9JuC
Kb4dZOCSpAlKeiNZmb94yuk+RiwgvlERx08znrs4tREdXklOM1gvR7Sq+PLmqiL8
bIBBaESnOtr/9bAP7fvhLiyelAtdZNsyDedfMwhcGJQ6pVHDXpZo7rO9t/44eS4D
WT1aIkCGJQpFM1W8StC9/Sc80uIQOhXqbT0dUfCns8v919cM+wsoAf3wupvCHan9
Xl9wDqJlFq5n1XYMltnvy4XOctTyMmw8owJfDPTBQXoyytRqmvaRUODsoHpXgyJX
m9YhM1xgaT8MPqN6ekTk3Q07csHvyfMLU+uKPETYiUOOm+DS+CPO4LvcCaa2tq+r
Jwr4NWuLPZbCB36VOvRLyJXb0ABdEGlzRPckqIlVn4t16lfeP4HcIxSVeUiYzvjo
fOXQUHcInSwtR1YWP5fUlIR5L7Zu0C1e1PImgHHLjka+/2Ds+nX5gcNHd1TqcNBq
7KkeT7I4FJRoPqQN23T8VknAZwLMNx6W0MeVCEbxdeFYjfjXgdmiqQTLCf33BkJp
NKozDVy9M/7rvhFvY0Zx0l+N6i+0yUyOoEkavfUqtoIkHgWrRcjbWM7nYHYV5a8G
EjYVJ23pfXBf+mJ1wkandu67E3rzR/jnpH3KWVp1SYyd5CEZnArkXzCrVLEO0jn7
zUPCvtnqWNs6udekDHnhPDR5UJ8yNu4nvAdlCrTkcicmomf/FSpWtMbLvphAh6Fq
RzflZzOPLFT9j9kzMhPxkDBPDOpToRgZsS1mZ0DlMuYC3a2iNbKWnXbA7vkVQs9e
MQTOopwtPFr+HDTdXSxMRd5oJfBtcH8Aa+7ZeApSRSpRO+OcibJP5+ijeu5CeAcq
gl0zl+QTv708/3Zw1IczUMakntwqU+7dT29Y07v4i1RbGNe3WJhq9MRqKUu/bh8m
L9AKL4KQ7Tk30RzK1bh2QgZ3pMnqknAtli5B3/vVvf+0p/nMKu+79fO+8A4RMYBE
hW01aISmjTyMFnkQ/Up166g1RNODM0ysepsMeMlPbmgmP2bt2XpGrRsPuD/AvFdT
fU5LKcPRggGmtb25fJgTp/l9oJ1NDr5D6//p6TnamwQ9J93oC2/82FC6JhfDCcnW
ejEAKLL28dvCBsaHgrpMeBA7FjFvNHidAcZMqkVgAE/9JeIesn0d/a+headKYFPI
7kDpH2gqTtB79JilVneflo3U7vb81Gwn9L3Qi4UNneiELfqIzXX3MY5gNMyAvRiT
oYuCc0U2vOWFbsFgMfQO/He0KbGCVpwQ832X73lFKDeOKu6ficFyhqKemZtPM6/r
wLe5p2NPwMM+9q3axf0vCz1yCsBSvuq3hSrbO2MFPLOdSyo2dHdWb8KSPa2fYVsg
GJrmONJcIpgDG0+SHOeazRdSE7BzsIf8bnj6r8G2sb3ejmYbsJiXTlSvJOYk9U5i
/JUaNqvogRdMasSYTf4K8KQ+AnXN6gcvXt4uKt/5fvREqO5f/5YwqLI7cxDo/xGP
B/fAlTacc77wvI8UKCg3ENZnZ3aeZyNTMr44KHBF/qXREk6aSkBnO88g393ILOJ1
35xDx/eb2mfG1PA2vPmHEg8e1dSSujpRnUP6XqR5hWiL+XcPzQGlTa0xAW4qbuUJ
1aTdICqH+qo1QDqSEGeSiXXRUjpGzEz6Gyh0sbkt8S1FIo4CV/MIa9lzX/igJmc5
GHWZ+fL/r3YkSL3grJ+dF3gKITtasw+IrArpTwJnNev7vXM5t4lIHAITqwzdZEy5
yFXW449NAcU7Mqm779w8qHNkHjc1vUNGuw9oUaUXKn2spmqi1K6k5SezNoXE9wLr
lm4b1Tjsyld89/5UwAVAZNe6HDBY5SHu914m5mWm+JS9Jnj+tr+v0tBgjOMpcgZv
pZKG93JPqqD6UGqDWMEbQ+Pn3bKU4T4CSDVmX9Y8UgMYzr7lbiLsyu7iAVU93Ofu
4W7pwOVnGZrz2fTYNxyNHba1+BKdmPENjYqo8GRZ6/nh4lwjGqp5W9uz9v8FrKr0
rHMnAlmvHiktOUXvMaKfrv8/uuK5BO1sGow4M3vj3k3YVMDJfPI+T7UO4mlzOgg4
UsC5grs4C6eYNkEia8lf5Ok9CECUWNl6bnjV2qo+o8okl1tWvmJ6YmY1XHD+7mNf
c0gY+2wCrwFklS5cm0SOmaTem9Ek7NJe5S6UhZg5b6yjFkSZfRedVnl1LnrMEok4
76CRhECxVtX2zAOld5OGwRRPpZD7lkF+hAwGePDC6MgvuRiYd146kAmh+8yDelPl
ZFk/T4bnmCnVv0U56MMjS1DsC/n/fdUs/kiEO+LPdE6cXLmSvFLFSBBiJIH3Fy8Q
ZlzgIvoJmVBla5wvpmGjzC2izyUVPULr/CSHuoMG+3bEXt+KJ3nTOTw1J9MXVVX8
ARKRS7dvndWEnUi4TFmedlhib+oGORUbVBcKW52ZADYibW7yIS/k8VU+xZXmL50x
lRinw2ACEfPjzBDNlko8AtNamDPZ5c5nb4lwcckrhCzfJnRxfcZ9gP0WxUejvlGv
K1B/7xxeu3rywCCkHnUrPAhg5BcWF1w0/6Sy5z/QiMOTNHfTsEDaW54XL9RnnnQ8
Ho0Q9nPP5UjFoTHpB/Y95wTlU3wqrysfa/MBHU6zve6nxJilagFjJZYNoYOnRiVX
ZBWp5jdwh1mV/nurg+Kh/wIne/w8cqM1VbKnJE25gD2+ukrp8N5oDI/ZR/0uF4zs
1dri5Xl9y22BHil/udsNFQ4MnEUUxMcaNeWrB0mLMCaodIbIXXuXPIsYXJkxLeCr
rMGaZB7rptPyMQ1elK5rvufrPUVp44WhmvzRbAhGRTgMRigDB0ZQGSVB4H2B0mQG
qM2OerB1MnO7rQV6J0luaiCcnCpxIPpg/B1FB//WEPKBh34WX+2HwvT0+43WQLg/
EX8e4oAjaueb0RnS7sxp4Wfo5Af0mnwRaCL+OLWUrivEKk7BoWdRW8rqj2PLTVTe
jMxRo5PhVeaG2bLgUr/Vo1apN7iqMBHMGLfvcM3XsQDCMonLI3GpvLGZ/UpGD7Jp
ITVoTVOx5cgGdFx9zmxwHT7bKf1PCpNu1amFrMA5ItUrxoheRbv1rDhJdu9FSBDX
pFr+PlyrmJj8uW7rOykY+qJCQ2DdaW5uY3tjE5tZF12JtPrIG6OmJbmvbTparmWS
6ANcinhljLUpOBJ5ZOGeFDsyrjzCURALyd8mpGF1KqM9WA3y43FqWEo42/YobetK
Z/uqRGYwT4jShFraAedJ6BwqFth6jW3jM051GdMLXjPfXK0C2qd7HE3BbMe8oz1C
Lo1bi2fdfsCTM+dQe0bova+ZaL0BK4TKj+JnkF7LsX8x9p533soENQrV65bSkykD
R/6TtYT6kcxOmznLqmyOZekPvHhe6xvwVf83uz18IfVyq2QeSUG+Jp5FpUAqat6S
MMLj8bvS3VUfZy3o0EjCxFRjQiql0GdIp2figofZ9Dx1GoRus9JJDvrF4MJV3iJ2
lCtJae2Y4TLvXlxIgHiYTvWyvPzxob0aAwzvoL9IfsUAxbCJcsOTBl9P3Wc7EKf7
EOjPQ3iYhkjtTnhW6gTQgBZjpmHIoq8g3Q8MG44UfXKEsm5g6qo8BXJaTt7Cw1ag
XRlW22npUi+n0zBWsD+hKM0nFeC8XV1acjarkBbTr7iPH2GRA9lyRX2ouK1z3Waz
Z757eDLg/vkCjJ24BX1Es4n3jyxejJSrZeujP63/RP6rE2KQI9fxQoeAeB8lLjwm
hE/eiZKtEyklgvtOty5pWejBVRrqHXj44Gxk+ub99C01vomUK6hsDtPJoFICKdlU
4HCESI0MidaBGHoMsVJBIENnPglVv6k47b4DjSBxBMJfNtYzUGDkaCXq1TeY4h7N
Anv4OvG0IGm6WrZH3zV/5mtEg/QGH0aKFjUrD0bzmBKOgZ+UkTsa21emEEUDwD0b
y+hadlDJiFy4GpyOUHHaa7GlBvGGKUde0F0Uf8mC94Fly0jSjuCMTvEZcfplngT4
T5Bw2WagWEpQcjzSoXsOV2HtoOzuft5spmia0IOSxnM1C7RXGgAqBdHkC/WSwDqR
UjO6giBeVt0VrWRKBBdbWKo7hr3m/Ufs+Vvkb8mS81uzyLadKtvn4uqbGMrfkum2
0XupLtzex8EiJd/EMt+CN+NBpZnKMOD8TAbvRqHYnQyK6Fda/Hs57nP+ukTVialP
+WnvlWMUEJthsfVfL/XtTdjnnN7YO+bKVZvXccpbqqOee4y56j7N01yA/lXHnmUn
Kko+rdEhkFnTx5y7PA7vwsQo5VCREMlVqMFelJMY8Oy3GfNmwHai3kia3UIMfa0S
bDHJYiEP7y/JXYsSVg8Kld4Ns3jFrWS7Q5QeM1z8gTCw0mp6OMQOFsjIWwUmfY0Z
WcK/9DlmbOa5KGwSBBCNTKWgGeHpCD/Ahr1Q+2rGu9pb5jSDXoujyOuDu0bs42Iu
N/IbzXQ213w60cbFXX5tYmpbRljaGfcLeDwdnzF5CtWbVG4bhLI9YIsmN87O7X1z
Gd6R9zYyexObbSliUrqxqrBRSRjrPJN3SSlo4er4ZmPIW3RWUBWTXjjOY7KavM2u
Ucjlm9nJPeDtDZXBaKiX5dnkgkse1op2IQgZJ9V6hNmCj46OOFBslqVOltwF5IAT
JIhGUJZNHWAirXpmMqCtu3lehIND6dw0NBISRn+G8tCO39VloHlEj/7fUaU5+XgD
mM/qNcV7bQDcWnxMugJVqwOrYiDz+S9Fw3437bVJ7lIC6f+a96uD0sxmdNt6vWt/
JePjQ+8sKKFwMEOqzlduR3CZpkA2zHw9JaZZgfvWKR0y2TJWSe/e7jx/LH9mflob
YPEEXUvQiDlkzw7MiyBQDyR7rWM2ed22hG9jgIlwb/T6sOdgurf/Hmo7C1zdl7Hd
RBVh86aABqy290Fgb6M3okNXt2WAxKw7snDgz6zkHy36FGm3UKqQ3Hf/yO5S7JQG
tacTByGvfkvM+MtwfMOof+tiLMHn2Z45rVlu0R9rQszK081iLyrIItMYu1CfSQZW
exA4QLrAo8D6VOjTbXEIfn9tOTrJC+YhM7bP6kI0ILa/vj+qjBcWniZd8jrUaODv
kj8QSuPzkKd/yzKj3uZlm5HGuxC7K7kPybV/UmXTM+ujPqy1MbXmi3z+c+lecSzX
EXUYEmNncIetK0yBZGCpqWaRuPRUOIxMludm5+Xxa3tIE0Gpdm4HLQzHkbU/bE4e
++nRIkAAaCqi0UH4YofQeHZyjvuG7dYr7tLhRZsVRrDspFQ+9AVS3ph4vGKaWkfL
mpjdt3Ba9T14dkvpQW2khho6064fVJJ2VOQZNPPtPAApUBbwodrDvNsDkLbiaCQi
ZGkv9P79EXKqfVBO5xZqBYjDM/fL+n/Mg1cT0OCPX9XbhmrnwRL+Pewswl056ehp
UKL9/4Mqr+QGHqTQExwKyBwbX6BDsoYt9akHdUhJY8HbPWs2a30LMq8RlPhyiCSw
rnoiKsFNhqhsnzuUxQ1I+jiy3l/fYvVx5AXNKVbx7Timst51gD4VgpOAFF8stkR0
tTD3U0O0JlfWSguO4dgmcl8R+RcDQS4DsNNQAULZ6gNwVf+XiRyJD71EBMwGpSRv
ut9bNEb7GERF+RSm9Los0NPvHkS0yfKxhcW1xuBUKsW9jJ/7KyHHKIQhGO8ux14L
DonlK+UaN1gv5sU9WfXO8IadvI2Zj3a04lZNGuutGPXPsA4oJsg55jgmi4WZAllt
PLThCBBKkBEUgZRLhCq/aOk2q1ntkX8mCv/ObH2+sF35tbznDOQFih4IgL/SXTpF
aCRB8fO+5teSEYSNtyfFnLUQLtvqvZb/nfqg5JynZ1BhYHJFtVWRXcB9U2P2/YTu
6AJcnwSEq0tW0hSKyIm9eno0eqydyOW8F78sDC1/AFiLCYU9XwdT6CgUa2buTEfO
VONfruhJ5pUpLQRTOTdlhu9S/SO8M8RgtJIx7JGEU0GQKq0xdxqSk/3STOt3BQxR
pgfmcuI2YxWhOHEIbs+t+qAHtXaEM+xWzNsjdfcAQ39qfSoddqdzviupYUqZOhJv
R5OlqYdFKmUEka8W0/ceOqacYMmZ7/ExMdrYrIBwJVFx6jUofAqRm0ssu750hlPs
Xyu9lILitQCZNB3B5vAEawmww7+bqXSn1w+xmHnCXUf/PhFx6CFt7laUUQpbxJTU
JH8rB+DFlmq2YLzarfuYF8BfXSk30Jg3MYbvK8cuxnU+7jcWB+MpyndqWmcPQ+6g
yvJasLcy+JlSCCRIoZP0XcKnDZFcXI4B4V9SCnMj0m6N8AaqHcY711p9QBVqtSEz
rSSdQXO8acOjXc2ML31/pNqHwfSusAuf5xM4B948zfopZrwKaDQ6MbYpehD8iQQN
nw8rrIUYNfvxhUChZE2D83VUI1NDDUT3lWhMa+FhSwKSNYaqoO3Dw03y/3ajfObF
Ho7EeE6oT3WjlyoA6JKwJTHRVzUDafzv6tRiL3Oa8n6aVHteE72Ju/4d5U+qZwT2
2dcHiVKQZTymCXz4yQP+62Vicsv3dIyKxY+Qg8xJUPbessm/1LBsYzXMgHHBDPf0
+WklkEE/AcU+zdMyvWLYWGMxDuE/FBXWA/T3XgyI/Ra+Stg7d8HPPeTRk3jX+J9M
2wPauOxsu8//BkRIslAEk6XmC91ErVkIxyM5GXbxlQsYrdC02NMkb9cxcgndV6Ht
tIp09rsx3qmMKos97n3wW7VJQkfy9rkaiaJF07ou9MDtThlsacnZddbNng3ewZ3D
LaWcT+Zl3dvVg8Az/0z2HUsEcQYtrBy59dZgUtheO+Au/oXHrDuw9Sv2XtAU5VZ/
srEZt6EqyKHk3v6DVuFO9xtXqIO8d3e9/9K5d547FjR8kiH80CmN7SNdMaPQBuMw
j5DoPjBBWR53QM0XLSPuzIyddlZ1Wt5WthqPSBuja+gO2QMerbokBmO11/cXV4GP
nRX34eSTXUjRETpdfyFbSGzvoN/zwUdXs0DjwUynbcqb1e0yguxnw5Tn8GYLI4X2
lhJ6Ne0TIChQpdYe6bVH3ZdMPtUHaspE6jMyHUltyhofhdFSnAAQE4Q2JbUIwkH1
oeq4UNVw6QOw5zkSVWu8STsBiW5MT2K8qsfafYbbB3p8WWHUH1l+a4Vn2Bnon4+z
Fgzh2wg/+Szo4Pg+utoBzptEJNPCZAxZ+90M04PU8v1zO/KEcm/hpL3k2gkL/QC+
D4wKJBFMCrjOv3o1eWDD1Tczq9SlHJPRQ5hp0LUZoEj3ZDm2nyLwf+tpqNPCjQes
dQ4WkzcIsoJbp+mcbLiPq+j031a6UMllPgOpv/sjNssTLTZcnj5L1Xmx9wB4p+Dz
vpscKw4Vrv1oID1iA78dqiuStHoPizfN2EOFQWXv0OUz3+btk9W7m4I9uOJCviKd
3yWEcl4gm0lnlG0c+HzLDnmYayyF4MS2Z7YZf9dgNLzCp0H162PlKskG14uryjLC
IU9glswUOcFsZdHuGMaPqFklPqcRr2KEOrhjJibMVUGCTQzpCgDElK5ncLukO1Zd
upxulIGYfNMD4+oBl3GQ4q7sDnMv4VT1BWP9CH6rioJgO7zKBPxhkLTIswIaNXoa
QjecWaj9SdD+BBYOLpbPotK6Uo3nwuH3HsT6xdINJA5CYFo2YYopaxdjkfz+oZSm
pQJR2AaYU2mjVINqv12r3ivWXxcJKqpZMhowKRhbpfopZ/i4Rs/ecbn0X/0HC7Fm
JyGOhytMrFSBFZ1z4OV7OWk3tZi6TyeYt2SHMGTojF+juDE1eA3wZk5L3vtyfRdf
0099HzUKp1UVG4DnTBEk06PmG8g9rcU8MyZIYfjcyDaI41Omxf7885gJJyufiY9v
r3Mcr2/JWeEKWcK92g0d5L4brehpTZmpz+H2BNAubdjrYhZzmPCeVudy54bHLpLW
iVJ+yhlgxTCj0ugCCCZIJMohw4NzPqg98fOGzTJAB0+XX2i1ECADacAbuErXfZE/
I9BRisn2OG+zpe+yHs0NJJar2uNVxmvQu6ZC0DgKg3JiiBNpb0/qbtMBf6k7m+kI
BzqrLwVxTlGXQdQ7uiqOwOZm4SLQ40wjGNg/zRefcerNRrd6upVn0Yr1aFDvVhHO
Jty8HKeCdL3Nm9B3fIi/F1/m8ADmoIMBW7fzGOLOXEW059Dzv7TP/vQatTV6OJWu
FK03pSHBWIAxgmz6qKVef6m7bVEKoZwcFOsz3brV3RWrxwRWc4eFYIRqTBtzN3O+
vAyHuTzvihHuYdFqSIYgJiv6Y6BqFZaUbnEXoaAW63OlMw7h7ovf309QVtO/BZZh
hWv4Dqd1hMklKqYJy6Byi4SXgBHUY+XtgjPRfZm1u3uHtbKMgA4UCRg7I4A0cowe
3i9fABohA3RlM/TdbV91iAt9pqF7tlSzg6qX0RjTBVtaT/OHztUlNSCKPMsVFIRu
DbzXueB/Uo29LvUFgMhk0UPOyhosH7NosjhrovCZ3teumpIHx6n2iZ4JIXsB24oT
BVOIVCIciY9EzE7rCk/Np5LwBJyeyhebfNVlvb+qGpLEppTArrjinmj+dH0N4Qy4
XpN47MwGWTI2+WTVcyQncC+R5cxsscpVcrQ2POAONsyWbJrixAhtrHpG2+FQApFM
xVwGrwvwrHiPD81RmSEu6/PqsEmgfTn16TNmzCDRTMv5QQ2UsnnV5wfdzThy1gXv
C86ThHW2hPtNYm9CxwTSIq8Eyu0fAQXu/hMCC2/+oo1vnB0GW2muQOKPk6tx7AC1
BVJwNz148DpLA8NPa91N0IoZ/BmuacZUie/TkIdaxDKAKEQ+Fenm/Tm3nBqIUY2C
NpTZJ9V1lON3PXZa5MMHe6BKecosZ+6L8d5Sl/q8b1lHWZ78L0RWqx2AO+YASvTg
KLMvOFYf284Q54329t1SYFh6NTzR739AcUofwbfsAR/j18abUrtnJR2UkU+xwkKh
t6EikFwVVLUNqIrJ3T4wJxwcGKEJiCnGCJlVZM9ac/IYBG6k06+UVhA6AJzrqKKO
7VoEm19Am5rsCgkAViY/8/SWbP+rwtVp2IobbGe1QxkHf/yVPO30NF8XX8fUXviZ
ZtVs9n4nPDZthq9PB0isP6t/4jmynRpZwAv6Ozv+R92Df6yfwd5HrHu3iG8lfzdv
oWxpOkP1yJMkz1+d0k4xQvvPybPO86keCYyfDBlSSC6kuHkjUCANrlZkMU797OJC
RZ3Rjm4dkme5gLzZZwHk+Rv4TdBNrEiNQ9l2TFlMiMO/QsShyHZnXAhj14+8aszn
PCcNYJskjqsUCHXHcM04RFiTNzedFJau1vmTlqD9EE5mUjBjoWzkJQytdHYGRkfy
03FMVzkx0soL5Sg3Z9K4xY9Cbl1hShRMNQE+QVGy/GEVQqIbjnh5FfnDDUMHpitS
w1xARR7uonQ3XKtg5DnaC4F8JlCMLh/8yxTuQ3LSie1mCKAHjwcaMTBqah+VIKwh
cMlCqrUmh79ETgT63omUB//hk+UrGtk/2400oXg6ar4oCCXK6OaGCs687fSaB72o
lBdo5gMj4mhVP0ZUfDnErDtrAm5bW4Ov0przVvC40+2U767FDzLRYaxR2StDxA/b
hFCjO8m9bUBueSq4fX2lfE0SR+hxvfH7h0pQfEJejN5pMhk/MvFHETTUIi1ooEg4
ehHCHolqNwcNhmsadRDE1tMv37xqzQSYBXlDa/T5eJbtp9ZzucVmmS68PInitSPM
0u9jVBVgKCas0BTcQ3Pt4rxuk0yZboLesolh+9PLjxFAlbo9eXCzbXEJAcnyIvZP
OjbDLT4BYAtDYJOABoT7lluvzQhSxXxt0dgPf1V4s3BetbnfUqkAS5BorbbOWWw+
Me6OiZ5PZ5lflP1AfOiBDwaurofjJlZ4HrOcUgNsxJF5HmCacyTA5yKezcqJZuxL
9gk+T8wxOdu9nIMDw6zqqGkC5NIa4DvLLvlwHtJKwmyR5Jlcpmctc8YdpllLQZzo
f1vTdwbDQnxhK6W8j129THGd64ktNF96+zWptCzYcub+9+H06O4b1894wWoItAvV
/6kpMskHwAYr3LKpoHDZUtCPqXIiSfzKrLcAscJKF+veSnfiaF73gyV4TjK7R8gh
S9eWJH+OXzCbZW0lXO3A5NbaiJixiU4H3TyleokkHFWgdsDbUM5rm1zL90TPx6kW
ikQvEHb/meHNCSFZ5DmBnVhTuyDcl93FrqtJxsuPlF69JtOmZH0BNUAUIR8D9HCK
OA7Mx8juOvw9Khxh2dRBFIhwIbReli7z8QZ0QdL8PLLsLs8cEoSLNP2wzh6X0ZYR
Zuv79RyI3vCHbDeRnyrTU5CnUBn+XsgSbECO9y+c7DLMf29ERJMJmOoD3pf2vA9h
vlpXZCDsDJ28lNOmTFU9fq80uffRQ5dtVxMnusmY04HsQ+NkNZknySbXTMy0YjnI
2aAGPlG9S2xiOMzhxCvSr4cKl6djEH2BwvHwyezYkhuGy7QqLr4+y6ueYc3rNAbG
wuHT1EEnSdA7NHqNE7TNPaGQlhISHVwLnF/Pb4s6UtL6Yg0i9+H5M30pWTrdsbD8
w5BxfEJdDM3e5/S1sqQrU2Oct+jt3VhfL5VwDPFDDXHoYtpTsS7EogDJHvNo3oLC
CCAQJW+BGxTwGAD8j2F+9DK4NuaWN/4tgU+F7iq0NIiRv/Dz17aGnjUOg65FRah6
my8GOaahaM/fwaeDDZAS1QWAy6e4fXpYgei2Han05QZeNqk2huMujgGQcqnCkg5E
aCc9R/1R+fC/QBz96DnIr4TkzNX6NLqqzTx5A+iuFblyVLw+uB6e36etmwbFnq0r
GeURlO+KLUDaLymy6MkniuEEchNZNZ6F0swPeoUJWDMZ8lHTudKFvfj6Ge6fhvSK
fDKgov7XpGrTf1zOYNn0CwwQI3hP6vNJ0OVBLgoF9n0hPCN/GRahR9d8jQIU+VUR
cNegpEBGCgAZe9NGCA5Os4tJ1UgHFEkQu3vgg7jsA5Bq2p3tZgQy0lcyAeJOdJ4u
U4FIUQJQ0mB/nJvCv1RbMfKJuRUPbdBtBEK1u4VBvZxtw0T7cdikEz+tXFjk6JaW
zKfIU6Yo1WecG2y6HsZNExkVZfzogdWdHymk6eRmYBWL20c3F8fslEUZfyodQ8gG
kBWdN66TObNddq0UIVTcrU5oY9SDGif28nFX9wwO5feYAQO1tk/2dmVolAp+vokB
WakraaLMPVkJGEQM0H3yfl8dzBUd0ghdDO+J0kHbuIWqynusU5iHEphV2Zv8Lu5s
B9QBRMCHsvvmT9bdErfVvTnMHp1p1CLf7ARMQ7Xd5iROtU+gSIkVo9/9H9oR468p
N4sXwnLvEcYYwi6CPsN/3SNA+FxsTKfgx/2w1NnYYBDfzdxWX8o+3gkJ3+kRj2Ve
GE5dRS4770d8FJ+Mzf7pmKiplQ2aPF6EqmXQd8DQpUCZQF2I67b/JxEWx7f4/7gG
VYf/NqOzWUqtksxKREwY+eaaPiuUhiJCMslaOGncB0xtLANP5LvC/mp3F+hFua6F
fpNOhCVrUB+WAhfVQR/nRffECT5LWWtLPpU+7/gVnOyNNZ1/UigsG5ZelcURtYVy
N5ZCU+DJYIIje8wyfEsOYHa+PUVrD9ddc5HozXfbKmuphrIXY0ZJA67BowAY32p1
TuC3Ik4d5MYNsHD46kTjraGzB+uowpja2bwaNospxhHdH1on2LImmH8VVpxaNgP4
R1KIRUXBQkikC2Znz9HsbGhsEGdwJSnD/VHmvof7a1UIkxrIN6OyQuDLZYNbiw6g
2Nm0prqTOklhmNnn2XNx9GN8sCpwJw/59Kk/qRq+Srn6oXAwhIXXx9/4nZxlGfAh
jUBArsQW6fN8meGV5NpEIqnSVIDj1mstX6X10A9BenRBS6g1oNNcEKnfvcUX+MW8
tJvSxAng7adQO4rg8fRq90X/UtSqocMUEI10Wo/rPTFW2jesPvKl0x4gxBje07TQ
X3BXbDUtdyQ3sFqOBaXKQNUVk18Q3wxhMyU+RNjhtw+kWWaW2CWd0J5gDVTXweDZ
GnPXgrJR4a6FOGU0I1CTnDPcMbxtxjJRJT4Az/8vgrkmpeEBHyqMdXhlHgSkInaM
0DuLCNiLdOdKRsxNqMuNpq9MSAetLoQyMRiw1XcjpoJZQJox9eATu4MRanhbg+9g
GOTkv7jZYOz6aM6wSRyrh5ARG/a9Y745m3YT9E4h2hHs4sjd61Im2rPQX1KEOZSz
eIRODqLK33ek2KlB8OhqGcETNmcqLu3fdmjm3hbICz+MombhU7WZ28HUXxSuUwDa
IpoRjNObLMfBvXfwcwoJ51IfRjC4hCm95lJfA4vdmnu9ZyqJpYaGv9bwKFJ29RSn
UfHNNlb0P8kD6LFvINlqBl9DoAJvT/oEIFNUTX6V/c41NPVSujm2aM6/R1Hb6jNu
UDfTQ+VhMo53RgKd6jdxRu8LDcz8HgKDAwwbGNLDJvbQ9m4ojuZ8yAu8RWrKXH5D
CFSzq8GDB2GFbJC7YIBRbODBTuAz/LufLfMCHpV+gWxlnZ2aZSYTjhT/X4SO+hMi
L8i5RZDZOUUY8is8POp8OWrqDqmPdkqx6aElzJdxfKKrG9m8zk7mXV1INrzeL+aX
3jL3eE9GIjx8uLlc135k6DOEWvSnkLDfExO7R83ksvrOJGLmEsA5TllKj1Lyotu1
66RV+f8x7udKkf1SO9JYGieeELsQSBQVhIAqmecbvTprTdwpO1TXqSa1u+foEiB4
uRBmO2qD6r8qgvy5P8g+6ZUdvkytd/wEs/k6EFmjrEHK7cfOBZrz3dtL4yly+Rkh
jSSe+sb2U5ovqdYO5eIG0dFCzV2dqPN/SthYMN8x+YrBhJvVb7XlXpGLP4Y/dm6j
ZDbGBddGrO/YLyPXCW72Yu1++RCQy16Ud/dgcf1dLdaLNQgSt1U1EPeT0j3W361S
pXhmsAR0ULkT5RiaOBGXQpajPp40et0jZEfDVsNCtKxSYH9WtEzibc4ouIs2fTN4
0roIl02JQB9SykpMRowyz4J4SaOKReqwu/HUkhXFFQhYbweRcJ3s66muecqZXijM
OZSJ718n49FSbESXNlvQD/aY6SdoqhzIDIFaavqbNWtj0mG5WOmvHmjD4tC1/MUa
RCZcEMx8c6Zk502ogATEaLBafP0tQRXpbQtGTNeMBgV/RWAU5nfZr+Svysd5ZK/h
i6fygaX0L0HSlLw8Y34Pm9bhEbdP/D23dl/CmxkUgxAS7duw+Fb5PGIcts0bLWnL
8KlA6zxtBpAu5UDTbi1FzUO1jmLQqAvLryfAVTPD8rSB8i7RBqGKo46uSXy9rAeN
ncZMHNia3d19w78d4aTgY6ILQNICVCGpH050Mh5EB9nZXp/rNNuG9Uf9J9CEW54I
BKFtiH/3h6taM4b6iUfWfCa+28JQb82QIS1WANMeh80oqhg8M/8C4e5b2FQKHnJQ
SugH/0QrKKcpH8TBaaq+9HutETD/w1ma5IQRTPZVbw4iVNl8qjHtPoc0/nyfCaj4
0jPGZcERMuPtGGFhB/fky2ZtCap1Vu7PQIQ8S1KBiqvp54URBY+srXJOZSVF/tbm
jGtcep1XkalSrPX+MrGmciKF9A3ZaXcggV8s19JJCBveriszL4FTQP9M6DEgvqB2
Z+2ARA51KMi6zquzq83RjdM802GGVHOYyLwz9GzJRtgkW7P1X8uY4x7bvTzvJLtf
`pragma protect end_protected
