// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:02:15 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
UxHbQAjUOrORvAoGP/GpbAF/oyC1AUx2yW4Io7gKFofiLGNaxB5paL8f8yYu4FcO
OWLw+Dc3v2rGIr0hVPQwRSi/QH8H1uR6dx1xnb9Rdqe7441TtKQguqafRpz9zwGV
6pn7gITMZK+7ZSKkpBhBe9TkTH+9FMOpbUI8mzplXj0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5296)
IjNaUZpBFr0NTbMDLnuDHVkdyNUe5Cw/Qmw0sh5p6ndhjIYgKO5tSEHSP6SN6wmE
IDBClMpQTIFtVlOEUMP4PhC9G7y+/eUDUO6nfef5I7qYE4PosVfg3Up7N8pGVXWA
1ySKPOvgnSLaDJYtYBbj6DyJbTr94vEu5amOQ7D7N3lXk96PHa9e3nrDihCh3P+i
wyxm6NFtyUreVcMuVosVUtuhTiz7Ooy4sis2m3gltD9b6xEYtnuBXHPmGpysruEc
l5cTTmfbulZNnfEZ7Lsf5I25mA7rsNOXh85KFyyVw4sd1C2PDkz8XI4n7jLUTGVO
Ho8Snk9+B7EhVvUgPok/HZEAbO4o3+wTWBfydZpFL7IFKj0+267Nrq2sAd8u/V8M
ehpi449fxFWa2scJpfc8fgKY6R82ftKaodxkFkAc/CGV+9IB1jYZmBqH3o/BDzU8
BwHLdZKMtuzftO/umimsh3bIPLXvcn5m3/h3p8gq73vWLh3Z196utxARzcrHf31G
AvRdZTiXH1gl1aTgLuzQIiLr5t3hqZws7VdVd7mbvesmxY0tue7V04atLac3PHHz
C/RXuabEKKfE0kJ4rX9ylEhJNixf0ZqDATyEiNVpaKlAjNLKBwjhQGniVf0C6WLD
aFqH4SwPexMZdNWPqRNuEcdHbYGCHuTovWMdgMlcGYVF1H5EhvDtswPaBrWihOZ4
O2TpVwfduH7PMDOnSlCIMqO+XBKuaZ/YVf8fObWU8TfJfIYZJktJqYPE+e1n8xUN
kX4BqohYBaqv0n6Xr+8zixUDZnin5PRE0zQgDxrfR94Y0SvR2YMCtTh8MgKPjh08
NXx6GGka8b2qZfLX8nN8Cqou0ZKwDIn3rrYaLAwK/99eFcPdqyEU6dSQcNxB36/Y
kllVcsjzvSy8od8ImMDJhkKGouQt6oJFoXaqCkOqMOMYUBkvxtNThQ/td4e/AIJm
rr7mhQxGgjA4XNNMgGjA3+pGKbR9Y25ZxE9vEDgD/0tTCxawLgjoAZ3YrhV66cgz
nL8G/PPcqV31qDR17rW489f1yAMxL3zrpSrJPGpoG7c/ceZZigZg9GnMsZ/wlTmX
TQ3chwlglVjHqfoEXS9ERCDf65DeIr3Qh2kp83xNBhLJ7SSm8yng+KT91/8COV0R
T67BA1EYB/zWq/DVz7ZcfP7dgQPrBk9itV2HuZhiOYXHw6b57LsNwsEOiTk5DlXc
SMegEIxDixhwtIhy5qRzgKN3O99SwG2LRySEjixipl+0c+yhMy5xWn9bfvX1EpEy
UNS+mE+bV7n2WLOT+6Nfh0gys9YBgr0tNLptXkXSWxCKdmFGaJmkeTXBQ4p2WmMV
avaNJtwLVnGhgHh3NJnY0XanXOa4yun/5DAHQnNUyFZ6pV6xL/303mis3GBOYOiK
vzXckia7dFSKmWiQRh79gv1zE64X63Rn8VBdHAPYixDJHte1ILbMZO9JW/yCxELa
yvBZGemzh/QHSxelm4mVm1OFN0uqaxQuHfrRa1DBFSFtkYinBgoOKPv/2t5SVNFZ
P/s53W2IyR9bRnEPgBEPYu4Br1Cz2a95KVzqE5CQ/c8apaCj2/UxZkQ+roO3OEx5
GbgOh17jYVMHo0QDtYi1/z8sNWBcbU0gTq5pBK3LApJ+k+SFbXSfBLqWGdSLdc/o
fvubWI8ORQZvrpnZ9w46DPecS51XxGJ+v7/Yk3C1nP0quMVm0mXxGpohptMMhN/E
kBL6ZGgpiWGFP/KIS2KXjZerp3JudilCsCNClcizkw+Nig92MHqG/l8u5DKi3RDL
VtzDzpy0IoZIXi43Qgfk+fbZeH4ZiBeXAqv+PNGxz/beHuz+aJvfUQOAuiFrry9R
tQut8EMRqaJtJfdDyU0kZi0b7tmzjVaM8D7gzoS9ONRJnjUwiM430FWiOc2lcO/E
B8kW/tchtvQ2Yrxp+jMiGgk+dCQIGfFiLHZTgvHTyHI0SrGvpg8mKaljEdgvUb/x
x3cALUdgvqJljCIHfIV2zKXLwGqrOa2ARmiYSFJ0LMHqPXPRyDh04D++tgyhVcEB
z4p6t0andtwL8v9/GLJtljDkHfq76MSmzSMCD3SLi+lG2JzdMF80rfehYIOesHbo
XkFJb9w5DtYEQjCD/h9QO5nR6KlqeH8rsjLRM4B9HC1cMkHrxEuIqr6PKR8CZI59
QWRXRCr53KTcIlX8Vi/Nz39ZpDCYegK5ve05jp8Q+jutbxN/JXJiCrszbKkJhgj6
TXAbrvimgU2TBwXyFHUK9lXGLS5GOAttREcI6gR+VAYpHbhuZIXQM8fYVxfQ95oN
cBRS6FkFucG8ezQgmw5zRUnZnuZrxUIiAL14PI6xW684JAFI7ospbqD3vo7/O0Nd
i62cdgMFfJHH/n8xnfwWxJ1feDOcW6slXX1ur7gbmwFaVz8BDRg8zQsTiGAnjQk0
x2zY2yScfcr4KcqYDW4uia0CODDYvNQfxadMQcy/aRLhX0vkwjnUv/UNSRwFF2TE
qVK3Z6hmVYBLhQr7ejymcDYp5WP6danDCi01eiZuzRVSZpr98NwmplT/QeYvhxCI
7O5dbo0x7KFJvQ7A9svk+JVHVqeip/fn6Dx7heLNTyPAKeaqT4ZC6NgflmkGWVXs
7osNfLJPnEbjGeKttQ808DPnkXPzSxXypwYScHLp96pILY2oKmaWMWRSmJNmznWf
OB3U49RR4Wkbthxg+cwT8nT2Bhv8ry1AkvAhcI47d6GoMC85hE6qkPCLjZ6Ypavn
WHguvZ5szHAX6TjTG82jxzjJ606O9awBxppUDTp0W4plGIjUkFjlx8QhTKLxrv6p
drEv1EVLtzjAseM1p4DTrd4CfG2r6lp7xd3Yjyu5VdSXjv81MI9JzsckIf62f+gL
SVhQARIaZ0F4FJ3Eerd3+p53sW3Wy6UUQusV2EtmZgBhL2+s99IwAF9K0Z0IApZa
mlGr7C9c4HSWGibgGhV9rln2SR7X/OxtSpgpyZBNPHSvksKP6/Um5UedVKiw970j
DT6nIEN+5tx78FM9qLy1j1OTaLwrmfYOAJHhIVRMkKQA8YdJ49tCl3/vxKJroWc/
+AyfuyDXfDK6ma0hjDM0QzkZe41tW3t1Qk/ATSY/FiTVXRb0INES9c2uxem5/hZc
6r+Egd2QbCA6MdvDvJMsgn/EJnDUnLGHA4Eu/RUhJ2LmcGOdK70Pb/hn1Kn6ni8J
L0n3HPwpIiolzjP4xlFxgZy9DmRpwM3teb/e3L2HHbYQfcwSp7VIUCdm4AZ/FGvV
0mpiVwdWI0KKzWwt/aAaZw1TtSxtyZ0ci386v7z0d7ny3EqNNrkMrnTINl/hXnT8
InNn2xcXrbkZbYUhedu3XXVlFrLK/oFw4FAPcPdjCRPXXiFlcf2TCbLMX0zIyM1d
aaKglQCEHyVtPW5H+V1Mr/17wd7mtX/lHxIhhkdRdPuTRnWJccioiy0+Be1jBMKR
xP1BCY54fIOIPsOh+j+FMtVhlU4itYUzqHpEIpPTwcOZogtvxHH4b8Pzi5jNUpsc
COAm8WsZp/1q6nerPhLD4UcC83JN7o4dYMq0egOjVzAt4jN/b0ErxtbLwolJKbHy
EebiM9bryis8IkZTvr8o4VeTy/+aA/WsaHNIPrwLhYoC66iuTQv5Fu9jAFQikx/J
Lz5F25lzgawcNmlhMnbPzsnF3SF1It4JKODO631mXWdrqfq/NniUEwKxIxQYrYF+
By1s40So6FQ1LxkiOIVP19804hLRcwvijSqGWwC3p2KgqdfKyOlw6/6Nw7WvurV4
2IdaZgjSRmX3Je+yGwEVzVInIL4GdRvpIU2uJ1G1/ea3idfiBNppuH1VChgd3Iz2
Stsjlw7dPCo65qs7IxW7yFkZlZP+IloKLHFvzDBN+pWZXeb/SHNSrminllab4GaJ
lw2XyOKWJmMvBq91Wd4MxYEAOH6I+QGWc9R3R5NDNgNP3mGwzXVdWBaqH/FdGsZI
8MCTf67OVrG19f+2Qy6XMbsL0wJMJJTsq3YeMU3MtKKfCV36XjkpzcxTlP+XI6Zi
kDoudVD4Fb3PEIlH2JhFEPLe4dHZPttIKTvuJ4aNMfxQEfMI1TgCZMco4gACTR3A
uE9lW6MB0o5nQZ1aeDBEB2SfEpVsWHjCaRDuh/uGvSCVn5r8Q2Yh8kQzYH2Nt3mF
au8+GA6NlgIijp3lFuRboH60785J/KbEfwQ9/a3pQoh50ZFn83fiASU1G9v3+jVv
Xi1ujGElKDTXTX0YnU2y7fYTP12LLoKcJ/YuDvJvREgBEmRnssd50KnGSyENDXEH
+x3VE8bLmuviNkawx7DLKZV/n/Mv0DH55oe7O7rvceYl4W+1IeFtKzuRKP0Dj9Ub
z1hLrJJPkWSS8hvyIAl4p8XgmUXt7QkhMUgVker+W3p/WjP/YTLw6pX7Z9SJ/MD6
kNdUbejgbH4+GNumnY0UanCZBn0sXvsfpSi6DBqTHX5GsCEcJO3UpvrQDlrdtlxT
vrMrXHwvsLUoTS5+bD+XQC+JIZczczSXzdpV3n/BQVtPrTeCcz/FYJN5vPy+Taq2
j/omH91BTTM2WYzEvfyHBeU3CSZ84s2OyD5TdTldX38SOQeZNocaHamFyJrAdFpJ
RNGzrJz+5nNmrGjYbsTArgJkEKUMJ48ZfdQZJ4aUBI0b5z/ojDbB7oioDDmuOVOE
aleBTsEw61aO+BoF8Xd/aKBJ/hN5pL9UMT5Ob2HVc3pB2YnXhHcbxF0Jiy2vvJhT
v5/ug0Irw3LzKlvqOxtDOJfw+naZu9vwER5rsjtKUVmJyw1FtYzTm3MTpz7xPgZc
18ZvenXN2i2yT/DMvHiuAnOQiQY0sUNtrVCnq+ZRxqUO3SbI3OcIZDfpgmgDQnVU
jheDHmo6/cbWTXehYK6ygwoUjY8ekzDJGalioXRWyXy6x0QSM2yygC0/4gjD73zQ
niIe0g9PpCgy81p4pMEb4qBXE4VP6l6nq0qHwX/E0+rR7un62+3Cgz9otEXsxHK8
wriiy6udx9QMF/fRhmRywwdVC0BSr9NuUFQ2R8GT0wd7XmeaMyXcdGq4X4iCWJ1w
9tBu9hRQD1tnIgRDZRvRLUYE8HcnxG3MOWk+4IRwcEFHCDthDDWXHLlyZoT/H0Ka
MuGDEFhd8H1p9p1zJZgh43pBNT9G1eGLut5uXgGM4qgpROZKvnoTcZvrPHHAKLpc
IXvM+jjP23VDW0+TlWnQ5isFJgdNrpukoyyyRJMmNxx9NcFlBJtNRFBwTvWR1TMN
IhI759UnTJY0ueqKBdnjBCOybskzt7vg4n7nEiCQ3zLJIV0+tHYhwzs2hA/YI8JY
U8NUusOmRqJKvFgYv9C+Qd8ET/i37i3GCCY8agU2zhOH5QjCwnunu6m2wP0kGdWb
e7jY0T6b7d1nrAbcEf/2WL2kWUCRaNIsnAL7mPzjqSMoBLIyvtmpuTIe+jvVuPGa
Pedjn46f1uoDArie9q/NCPKnJpiJb7Uf1KLovnqSe8SqE71tusWmXiy7GY/CsKrR
4Q252eUZXRAbER8t6atIc1FcphIdQDVqhKbhpjyngOvX2Eg1WGKCnbiH75HKBnhb
HKif07rXM20qGZyAntKDTiV4SYqIyxk2oMLRB2Kk1tJJZk4KfbDNlF8CS47ykBJT
OdX69J4mZHyS1eqGRHcb58wkaHvM6ooKQAsID/gIfGBm14E08IYaR54uAkw9b70w
iJKg47yI3U9Qe/2HxHRxl3dNj05FsmCf66Dejno5nH9KMvYUewp0twfM+Gv82ATl
LFIsDXtqH1bX9uv6bXqohiumlouxdStXU4RuGZoAnpLD4Pkjl6vxITEhb8Pobzcw
vGWd/xA+1hKoxQ+NGhKGKB3EOqYGQI+BmdYE/SByGHA3fhypjQ/ivbT1QGOi9Vgp
se33IeILWMNsV5KH0fTbFpNZC3+nObLVnekS9/hBHfzsW7mOBrma+fTWTiQ7MBdW
G7GSAZB8hpXpYrys9+Nn9ckxnKoYH6dk2SiTYul+587RfePnMuN3YBFVMRaL3h0J
AFd43NY6P8G9ABzY4s5Ife3f+ruBMTgRdLuDJ9FwnHVCNp/ovMV7wrojiWzasZ/1
mc0jE9K6IpF2fiv8uvZkD2mmOublWzQ9Nhy4uZ+3r4OuoUSvHagaUGJOz5+NCsW8
eHG0OPsRdcjD27Xzi92klTQmUoj5TITfLHg2xAy3uL7fPVaY/2GxAIht8Ml/AiTT
RW1yEPUKSII7han48k7CO8gXOJT130lD7obwEQXZqWCthe1Wa7GwBy1cXdc3JNnd
DRKUDoqmHgusVUim6Z7MR9gvjTCEOdoeZw7YureNSQjEnyKSG36CGDt2qFXe7iPj
bID/sodtwDIR9P62VrCKMtuhCyQw4kD6ck/yhgVExc4CHTMc4SasWUXuVU2I59xk
HS+g0NhEQTt3jSTANbB74PgjktFm0Mn9N7VbHn1Ufj7X8QlpusFxcjwUG2eWtOpp
RMJQYm0eGNeQt3z4ZwGR1NRcG7jN/wCYrUYXggYiS48ld00+jWa2ovUFo+o0J0RM
OlbDD6A6juxjATlj00LqiahZN4mS6MyEGu8PgoilNNWlS7zJVqm1Ku20RkgiVYiZ
//gKffDadaeXNNwxbw5nJQLbiD3nXPFXryt6C4WXlPbcI7xi7jPIFJcCdGLnODVe
GG4oYA0kpcRNDVZRz80pMm0z1oSvsux+MHACMYf/L8GOJgmyoxDi/53s5Ky61yyT
jF6GvL+1u/nTVLoJzdLo9QCdpi8/0A1SZtranUOZIhByj4jYpdVjcOEwO7q1PO9u
ZvssPozYlxsipkze3rlw1vcqPdET0bCVG68m20yw8ALzecRJ5a9LHgVKBbuvWA0k
la8Lkk0gT3wnxWwGFvl/aW3kuDR8fkBf1/lV05pfPnDxE/mHLITMMalbfBN6C5cN
DJVpc/lGg9JgaQmcihTQn/+YhHNi8bqEb+wNHxOxkEV5l9PfejnyI9flZVAMHvO0
YcPWsTA1BvqnylIjJ76rvSI4+1pzAKb9VT+uBauNqgYS8vwVEASRX0wcxWvWJ7MG
cBitrZzrVR2Qea/S9OLfZQ==
`pragma protect end_protected
