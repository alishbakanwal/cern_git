// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:05:28 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
RzNUZURPbh9lCHM1y6NWwhZHZnu4I+QqDaij3W461q1el5NuwDCOHLbTJ+/tk7Pu
khiQj1CGnJjgQHJCiX6kKlDvPz+qTCymdt85Z+2UQ4XQnUcH138ZRtrz4Cai0tAt
PI29QnLtuRvzI3yn3QVMCaVI3RdCoWQ8uHXyIZfco00=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 18752)
FZkyA55m4y583r1fxCQThB5x/wgPBRLytHfCpnClFYjK4dzRQC24nxQeDxdZsExp
Sd4C3jJf0AKX6FU5nogoH8gSeg7Rre09JvN318DqbSpcEjqZlWm3U9mgZLDDSf1T
DekQHLMx6tR6KRl1b57KnBTnoicyqeHoOupSiyOQK/j1conTPQ2QqNKR7rAlZogP
e374Jsykole/iN86J+OL44HM8fa2a/Y6Eb0IO5IVklUEZ0pqHy/LHgnaPjmcOI/g
KHfO63ALRFCL51WygwatMuXkCkT2w4h6XHWjswWS4itqztM63L7uLDyZE164g8Us
jR3wu/kqDVSyg2DdwI/1I90DgTUkrfmUpXMCe84MkNCMz+pEQadL1kHNiEcDx6Xb
3UMUfGGHrVnxa/zPAtKsO/QMH34I9y1njnRpAQJKGqxVw3jvR8fVKvP4zH1FVwQQ
YPFoV0ftogA5fDJOg2CqOwsZwxU8CaXkr2VgXW1Ac9TUzB05FY9oBSS2Bb5ii9LC
/1Xdh3Fs0Xgk5T8fDxYAcPVu7t8chAOKAcsa15Mh6e1m6w25ADZNdVn8IsV1SwXy
9AWXWJxiGyJwUCFVdIN9zNJSRMZJiNeDMK4E3kfMw468/xmIbUD0df3CZ6rWU+TU
sdaLG7f790+rIC9ESPoEEh+FX3SC8xUPaNSV8XMSg/Effwcdv+ZOshwA0An2QzT2
H0s2MzUa8K3Ouy4xIrKHKX56McbPKKTD2OkHvVxg6pCSTMJYwKSU78hY89Th3Yl9
FTAmi1wNm0VayfO1CUGZyCmwzhyHi36gAGIjNk08OmvqnjEplMSKM4nnU720dmyi
YJ3rsr/rMJXA1vAu0/5Z5jtHjOZB1ZzTgOBuCoL4yLLVjT1JSeY7rbOup4Pob2mJ
B3CVYPtvyMg4GlloueIiO5WaVicRy7ftwjVdCUpdf+G5irmM3HjQdBdP1DL7UXmr
HfSIJpWOp3Y2SGcinBmNQBUHM2+/d829SDRZQviE2uETj6eRpNp1DBJCr75eIFuK
kvg09rz0wrx5E6ViKUHBdY0H6MPLHd9ydoZIpWusLqp03oJndS3g92AO7+QDX+a4
2YbH6Pny5ovxLHyN5cNfA7UPmYMSNumC+GhrLV2bd0+zMaoYn9DBN43zJQUo+jwI
8Jo8ke1NUAgJiFAra1RS22/+Zgpx+AbcMPDwBP/j8cXCWY7Yf3+R7UeKsmPxOfer
onsphyFtsIuZeCguZqPLVYHGn/AM0Fw9Fa8NS0Cm3Thyrf5Ev4Fh6jy4hfYIFqGB
DI0fSReSRGDXL1nUTXfrdxYvU88JhsSVn5jsTFvnMvwF0vF6MWAR7B6/faTjzC6G
ReK3yo98sEUPzF0zbmkj+E5jF8xN753hbIFldaMW85YaAcbNvpjyNtk5W7igGpZb
248chpjslS2HF0VIEOPC3ghE1mxlsI5mQIG2/duVzguyKdo3WcgP9RlOpH/VX9YX
OYlnTbrClP43KMB98ygwL2J2i6GAPd3ASTW7xR07zfCCsDcLu4JBwfVJeTLuRh85
4ha7B05BmNuewHl1SZX3+HK7Uf0OUSgzlsG3NBKVyJ3zh3YYUqBGTcJ49XQVQyab
4lCVEJXa1sRKoQ3FYh2ZsxHnFmyQuBqJwhtfDTB5ypL3vyqSvyNUqp5I7IRYzQqU
CBLvr+z9u9ZiSzTJ0mUojOmephr7tyLAXo0Xr1xPBEkzWLBJaRR6TdevrMJGfMx8
Ir3TVU9reFE96BEE5ax1Yv02+uMFNKdslYtFdIUX/P0rV3jyH0pVd/tBosJYtNxK
4X1N85A4GaK9wKY3/CuMg7zCY6c68qhrHWgiXAS7Rn9+fVtFsrrwFhueAq4tuQW+
ZgW3S2F8wY/PZVaxFSsEF21ToGs6pfEjpZ9aTFc+h3E75a3XepGKHXG000UpXkyY
jDfvNCL3hklBIP+FSxHw728DYKmcUkTcbpCL+K6fzdF3m0hir78akXJfd4XauLt4
hThLWEZimKHhVXksHmvBSE/rvbQtkGAR6XfUDVYeX0JrVYPF8/lwbZtXQqKol82s
wfDqX2zduGvVPOCYEZBoquNC73Kf0PrqW5823Qk446sDkS3narESPvifQ1imu1Ne
J4gpq4co2as8jXmEf2W+uZCzyoAgSzUpA8JxIj6hRI+OvKJAzyWiQ6nDxE2whZBJ
bNFQ4e04El758DU1y1omEQzmGN/acDQdzhR0E3a4fuy18Qru2mq9rlvgcgCoi/le
z0B4m3CsPuJ+NGUuDPvMf+QnReUmX+aI8DQmKojq7aeyDu9Syxkal3XWt0KrUWQd
ju2BKfvX3N6FMDuD720BsaYxrRjUQi9FeTD1ppveOMgAFvvFqVd6tXQkXm+J18Mf
q9IXpgRETstOhGQpLXO+LjDw3b6nTVb9ge/Wp0RssPRGQZzg555HcdfgZab2/EuO
J4549ZUrn7/STFRvxC84CT67v0hQYGYvdOd3N3UkBroyGPLws2YoY644EDTNNwFi
NZeX6tjxvQeFEfcENqpP9NiHtsXbmcX4oXlSKNPnhywwmrcmTxsqpboJXe9ZYNn/
rI4GaPsa1S2hEDAOpb8kAcghtIjxQdYhzRG2ARzksIgnKjZuy0DAt8f48aTisTxh
NnE/iC1cMEHzEs1h7gd8tnEhawudpCZaaEdB+e1iJITDg8TEt+2KzIl5M3FQ0RCw
vZzX6b7dR8U/bZA8vSnGBbL1FpvE6xw0dP35nYkHM2UzgxXC5WjhsPATBcvjnGOh
4re+YUtMxgfB84RWz/pPSh4wBlDI8wMNSKkc2IszRCQiO4q07JTi0S3jLx2fJkj1
YfVP8ha1X7PR/AcX8XQqJcKH6cTwR0/Ur0jQJjasU7km9TAYV1hCbRVS5d4HQvdW
D62eFfYn4yToDgeJGD/4xDzn15FBHVPMa1D4Xlkd6bokpYJSTFrRA1hDYm28bLdQ
194KfgTws647VLm2PfkFm8YWOCQM9ILfYMJs7PVI96hL5fjpuqDrSgGMsvGpSlNN
DrD3I23PHMIb4jHy7N/7QFo4sm5aMxmLvP59gR5m67j4dw0QSLlFOIb7W/xeNjkm
DPxe9jEAE+hRz1gHUJI7UnW4UzZnlPggYGVMed+wtqDA1MIAa7E02G0sJ6piH9pt
RfJSxxVHckMhEy5sjmWmA0vWHkP0BkuQ8CEIjT2LgNuyEUloM7KCaH5S9n+4yNjK
eTHePhKq3Hh0HDhHnUx0QgcuuLV1SndUK1twSOzlFEWVCLc57GTK6oQp87sTS+qh
47af5vFcU6Gq0xe2gIRgXyU905UAK+ou1pKpVTfUmmFJ+7yWqa6BksllI3YQAt3v
7s9GUKdDMsidbhLA/cPaJV46003R+glOnz1Yht6Je2x0KcsaG1uxkietERVjXVjb
MEaYd6CRLIOiriPDL59yS+FyhhyD1MMKF6ZU/xCAg+kLDPi6VpVub1nk0UZ5UCo2
PCIJmUdxq/PdwkuyCbH/R0+zGLY+fWJxGyxCQGnADdi1AoaoDthdmswFhu/AhGeC
3eg0z4i/pj8EVlI3lxgTco+CS8GZauu9gAuIbWAr/S7c6B0NXRmQFzkRf/SfoWYU
oyxzF3dalBW9azGu+kLDTZat4L5TcWKJMkOknV6lY1sdyYyjX8RxhIgRI+bRTXZ4
+pSz25Po+XfndSXoH66EHLooWBfEvWPJ7mq9NlIxfy3gXvw746jM6K/Uwcyrprp/
WQwSa3cuRmpOROpmgkWbE0NLqngzZ8p2YSCR2ItS4glUm6cZ/DLQqnkJqvYNbdID
MFks7x1cAg1fzCVVHFi6S4SJlIyTSb7f4QuOP/AmByYKrbYW11sqjY2/3O+++iQ2
TViqmd0vUod2D61Z20WxI+J1f8yCqZid+UxQITuPb3MWZeZ36QW8nY+aBeUTTkpC
a1ikTB9ndmpXrjF2n7DhrGTahw2t53d0dGQ44bx1Z0uayv0kRDW9ZjFNlVsr/hPW
ibsSIX2Ce1ije2coI1sYEFrVGoPgwd8EvIoiN4L80gksvP3ajfz/AL3FWibmtHWy
XXFhPoXGtkDVzdC041SPstVi2vJ6abmPCMUTtdmG+8Sc+8Bou7+PzRT8V7hukvN1
aj41t9FJDoFJ0t5Y9nZd51EnpSU+2BTQY+/82L3urvr3Z7cMipQSObHTUQANIi2z
to+DBYVBKdX8dkEZTM8aWPjPbSNkDXhVcUhZ51ovoN93UDzcpeIsv0QfK+C8DDRE
5EuEZi8RqJ1ZV1uTvDqkwNW7lS3/KqW0M7YzR6fjm2CMTajKlnriprsoFwSC3+jC
petONfUXiIBEtA8LqlwO/EP8GuV+WZlVvRPoCe9hhZ5ei3Z/PDtf3u8M0HU1/OlT
SYgcZ7U6etHOehovpOgdFF5jfH6mE2qd04MtSCXxTsrPn4AtZFAoQ7qMGIzX4cAb
Re78yGsmbQe+8G7RQfO3ncxLWDcj0499VJsQ5XX89ZLBS5GvNAD54TnRw2ef9kw8
j/Ly1qGokyQGFFsGSxGwnpAHrYeW4j/GXEio/WdapW4wE3090J1k/cPhM1YeLXXt
UBZJy3Vt4MoOoYrC6z1RxjIJVxmf1N0JVWP7owdSFW05kw4h6bo12dPO2RiQo+TP
9qklYVZ6tw27fth7fWz8nqpuJ/HUrs+LnIPJVzqGo2LwRuDEvUTvCEglSX1sCS/5
uwUvCOh549XSkUW+i9s0b/QFq0XXN/rbP5DWr/Hp2g5b2QHD9oRoNBuKWzQq4H3B
k088wVXYnzakF7cb5jq/LPdg9N7gfeQYwtSMmygpz1fEEd65Iwjou8euYNQ/vFUA
uvvcwocXJcFrI7Y9O6uIgqqqzJXuoCsZkJGXtFU2URaX3KpPnFb9WFuJ7snDCD6w
VwdVzGigKvSuFCVVIJyDSlW1uO9TVVJVcCxWt3N5q8X37xpuKvnuswZOkwPjMcDZ
xhjiFCYnx6s6f1KBtOrWUgANOzEYB2lebYjjZc/IVpEkxCD07mAbjNe2jY1XLKKE
RX7Xv8KHGcPjRiCdEno74tQpkj16hH9ToaKSm6zB/AgRU9TQ9lIdNICFPUWGZier
SDNVZhrVFC6nbP+PM9OoQCCCwTjYlLJyaKp+OIBdHTq4NTGY63cIYS73gbQ860s3
M4Y4ns6EYcPFIZq/PLPdJNNIx1k/JzNPLQcOtZdh/Y03O4IV6TsxTZESJDXFNuop
9/dTrW21MaAYOWDTXUAse0HUhgL3/wKgs8/VPxI3LTt9o0Cgsioux7vJKpcdAesq
ug5Ce1S+lMq6jlts9CA/qEOAMzTJk5XbaGQ4snE9Tsfjr5YKYUxGRgx/MTYsS025
KgyQvVWQhdTQyDLE543DrkKOfvDvXi1gK5PuF69oZr53XT4xHzH2KTQ9HBiaI246
a5e4dATSCqwfOVit4JZYkOrGF2Qd0ihYutOe477MekAbmqOLkn0ctcr+IE3fhYiQ
d+ioHfS8zWfCZGu0xenD58KpHEWaGcnaWO9xH0p43yTAJrYAjOos3197q/8T+tEl
NrLtOJPlJW7nbYQ9VjaCJ59jwLAbkwLQRx3aVqashUVZoJvF7nUZmlxKg9ojp0zB
qSsyNxDlo9JZNi5pDvoBOa/cJpEeGp3liznCnznJG3qwtbo4wZG14E9M3cckDSmv
jKZdUf/To+uQoTnRs6u0BK5Y6t0LL6UYv/RB23+vnzjYFWovvsOmF41HcNgE7oss
tc9+tALkaxCIVf9cXr4eYiy/LMxk4KPL1V7Ba/X1Wzl9mP2ZrBtlkb+mk6rmdJJk
AyS9nYkd7kPvzkDBJB1rWRrJq+ltH77J2GNMm0lsvPiD+TxitDHhbhFQvq5ldvZ8
+XKG0yO8MAYSCTGsQUNyQ2vNJ0eEoLJohXA4JiOk897C52dnj2Ejvaav52XWBAan
OEPGpLR/+VqUkvdF+PnUu0esT9sh710Eoyn3r4zCoJqjxiY92pllsbFUzfNrvJm+
2cc5bqX0+fPCEP7Yn1wXtmsu2yU4vv/uiWeU3v+6hEyIzFjl3BURNm3loqvnmOL9
3aNucb5kUxkN7Z2XHkM3J6pB/AHreWmmcDth/5t1TfHsvMY7T+p4PjLlEg1gBVzB
7SxRDy6+F2kAs6UJOtXNa88YPe2Eh55egpRYNUuj7PJ2K3DzhMwqdVOH60bxRAcB
/bgw6P3T+CGN1PXl0iPJH5PBtQKIvbTDRs2pqU2c+o9si/yBsX7KOUlOR5aUfKfe
uGXIdY/A4FgoKgwfLMNfZd9F6ZslumK0RnWpzRMcASzgnmmK+RAhwnFSZc9haxET
7OTzMscWpHRutUe3M8xfIzqjMKkLX0AmddnsqyzcUsbokwVUNASpaTkIuKL9yM6Y
3TOEKILwLrI/pgvH1nrapz4aDd6AQsbq8ux+REQMVWDhGMoJvbqYaFigNL0VXD2m
BU272UuWqNjlKKBM3eyzKRSYcgSgHGNfn44zW4fahfZ756Q5cq9za552P0lt8FYe
DJEWW/skN1E76ZN0zOtmg87DLt3Rc75b7la77o+/bFYjjneYGbgEpIcDFPFcGZxa
74F2kIsDgryVlKYjO6N4/ZmIAVbp0p0Y8ZzDkwJKwOBeAAWXlrbvcMGeGPXppmBz
Nyo3r4y9fTT7gyeN9DSIIY3afmxgCs3uLugjyF8YizTzzpWParxw5gPvQGTQ0bQT
tAxuVRwgeQtwf6XGTO5G+GSRfYu1DA10Pmx/B6iof5ZsBgm4npT4Cp4yU1l1vVu7
b5hOzB4rWUZgXHVAW6pjwZzZzqOrZarsnm79zoQ6IWGqan/1VVdaupgD3Ssl3s7J
cRBXoy5uXTC1mjsunbRMj/AH3qcKDGfVlOR8Iuqjq/yJ3UVgCnK7C26ysmyhjtGG
VM9tPU1KNs4vKZmmvSJssxLUOOTAEI1zCVu8DgtIRH+hViCIMdwPb+iGbSIaCi6g
PZ7WWHx7uOPY8diHsxDVWkRl92f/FbHJmvTJ673thoY8wR2l6ldQS3wPNX6/2CHg
WHWN4LTDbmTU2j2xJobYKnK5YffI35RCd0ZJrH5/imdFDXJSKzfWJsefgORRCm3Y
ru33tseS0GZG9DPA6iGcIb6m0ONEFoytgAB3IYO00YwnU4h5WWNSOJ1YJwVKbY00
b0o5CMw5l5LKt7AoIPd7OOjxE9nPiNrOuvpp5cMmNMvmZO1kC5op4tpGgByK6d1C
ou5XHHB56wUw5ctf/FArSGC6uG+3qhJqq0Y0X0E/O3XPd4wIAarMmM6xnBryaznm
kMIIjUv3A/tyIQ2F3/YTt+zJ9OnVewX2SY8/BhwbfipDpc3DkgdoOE45Vpce8lWc
J6fCBBDCibFOjbmnv2pvoDyWPU67K8BCB/KZsNEn3mZDNg5na+jDIRKc4Gzfdqn1
DdG2q1xNSS+cXnvalNkl9QdBauB1hnT6s1Py8rV/ItkGcYg8qhYInwDpPMvY5hcx
BbE9EDEgmihLQMFwRDnG6wRdUfSa6552eo0gnECe5nI5lN4YXWGgspW2kulhx++d
fM2RXmBASMkMpnvD/wFmyI6NLFNqk2fdzLnRSN7u3uoVnNySr/A+haZnj/EDN9bB
Sq+/rVFgu7Kkd0zZ33cGycQl1mY+4UTa9WS83yRToeAl1q+PTheb8n6BSqGAnf0r
Dgax3pGBnZITSWLNj3ht+rjiu9odclKeiBR2NNLkH59hYKu4e7k5VEMPJ1+jOi4Q
Q8Doj0opdLmHRBQhssh+QvtjGkz6L78hAkMncv07XbkHTxuvN0scybWNMVwb0UiA
7KGVJ+KLqNYcvDuaPth+QNzA5IWFsQxwRTptNAbLXkbs+XoMaPfJTO3af32XI0Jz
NVr8c4nscd542yqr51nKaEhjxstYwEugfEMskzbu0sPRdX7gIIDbE5xRw8hYc8SQ
YUQLiO74UFqhSyrmI2wvELsnxJmsSRCCCEmzKtDD+soDYOOsnIrUIoJmTZzF1sRK
Hir/kta7751GzSiV1UAKuQuyqkdEcYTffR3NXyVV/8ViApArLV63pT1fAPEGpWzx
SheBQOclIy4XSn/lMWaNqiG4wkO72Qx9Lml5cMTwmvDQUBdR7CPwhwwFAP58YbzB
0HSfsr+RpRcme75GiyX/03Nn/4oO3Xavx+eyfJjVOEnXddkSwoG1Q256uTVhFf92
stRnOk+qIlOaRwuu/jNFcsAaT/W+wya2R8go9eD8f1G3g6ZKFtFjXdWr7HkaIZ8S
OT6rDuUOtx9+A18dnq9nlO6deHNsSHrVruawyQeuOSfkZVgndpIF1ZDn9+A2GQJq
G7S3CKld2proo9cWUmP2l7ArSGQR63YfENz8jb17GFrYZgwWoqmTP/brRs5LcA+U
rgI9WQyGHcvpP2ODhGxTpBIrPAt4whNSzNNVsuBDoDnV/2vj6JUT2HOeXJhg3Ilh
JnmB+vFoGd9ZUkWxiUeylrwn4u+Thffxol3PbW1WFPBcQo+9FuLkq5pFF5dv1X2g
ybh2u7OCIY8KZFOhdhmEsPz1uuA1qi3n0etT/r71fAcK9lcZd18vCEaOTywjVjBL
fxNWEPhspXV9gSdOIciMgrPQOmAFEUDP0rep+dYiOo7gSIR/A4w83iseRLQxS5B0
dZqshm6OGlUBskn39v+mdg7P9ziJR3NcWahBwoQ/jdWH+oFaFYm7bpJg+FhYW+Le
kyiwJvW7hKtc91dXZjNAgjJxWeMh/J+cHh8HQm+q6uv/x3lNJEV/xyj5cuce7zgM
cu7tP6egoufgCFuGk7udcwzvbHMLiwgSocqjlHaF1+qXXrW22URH0h9oxcB51Bgp
LwcGxXW91dxhW61ZQaDZWL1zkuvWGx1vd1syh60SEgWy93leRCQIT1obinfpdb04
1JM/3lkMfq3C5Gmf8rCApKuIDI1Km3pJPBlZ6LFC3cI8Wj+TrEj+XdAECgyOo28n
FeU1kdQJ+DPsNqm24Hpl8P7gsb5lQYzcylikJtESgjkLMghnN5anih+H3oGlgyW1
hmb7xl0MX68rIU4XTuz7iGaqFalkBOR8GzRFgkfGQrC+g2X2BrNjC2+LhQ6ctZv2
R5d6yOtNyOH/S1DYkuT0GyBGwlT49I/NdX5/DDXTJ8RmACrSpHHl4xldOBSPOhTE
2LG4XhP23Qr11DHcvmbNn9AANdnX3JDAvwBtfoZWQejlVECQx4Ux0u4eloulMkwx
MSbihp5783vg5tclqjvzrh1eHqHZPqD5WhpSmGcz90vVFifLktwhq1QPR6bdX8wM
Lmhmcxv1NbufwFaEQcW5gRUtKX3fBECjv8nywvAm5I1cm6NoSf+6KBJfMrlYeyW4
xLhWEhxx1QfJqvKqJzR/kJEH43rIiBiWetILRu46NqkLtKt73rZsBKPC9oWpCxrl
6pn+n50MWwJp0yhxSWZ/yWpgzcq2XXzdb6fyZU4cnJwn7gZezBTe1OgY8PTlWAER
/dpyevsPc0BMrSBbMvFYJ8PLj1l9TMmOGzHxj8QKeox7Bk80/OZ1xMnv89RMYZgl
QAy+2jPL+ALF7aG0BnJ1KsltX10TNHL+JtoS4aqJv89nLXowY28Sh0KesrE5NK8N
4mo0b9fZvfBL82QjkgnWsgl3Or0mzNYH4r28jHiLXXQUVtNqGU/pFiIRhy/ItFMA
ijdAw+5VEf33dTKgPUYx0w5+vWDlqLgqzAxx0r63EVfZ0gEv9LA9lxBOUYnhDJCa
NtVOVKeNls6RXfw2RcmtPmoRRPc2UE32TARp8j+Qtif4KV6Y0H/YiPOvtWHBHgRL
YbJm9WEOI/E5JmwipkDxXX0dWJ2RMVfdFd+cFWi2YmP/sNfNvlHoh3KANGcWm1Ko
FwxylEgDWivZ/JRgZvTRj2TjXVcMDXf7el4HcGDmFvUQ9o/UGTCuXgnwzbeNxBwT
q9MwF9RxDubzDoRKJleBwCcZhC00uuKYqfIxATK47uR8tNV+rMC8tv6WcCXs3tCW
skUc7JJvBLR7j3WDE5uhxRZeDtvDcC+UZ9GCB9lKnsl4iTmg24hT75jIGbxkB2ci
7y1KoS11BxNKXcX3qXPd8HyW9+QY7xyiZMur1DJmIbDu+FcC4pC+M6y2Rp9VV7Hu
sC55ScVMuN+QZOEaEgLneJwTHNWGHiAQlPE0d5qbAT2J+CYJiCm9s+NS6oe5kLmk
tBV4A5iu7zZsN9uwiGQsdPpFH+gCudEBuZ8Cdlz6QjzsuhJZu5F+daVDD6zavsYy
iI7Hq6sGzBUhZq5ZMSdGFbY9jNyaz2tMS1m+E/f5WUHAOjg3lpEYqbkwciLYCAns
OvccaGivolJmWO5MpVHlFKAkn/1uCdVN4XZMLbvhCBelL2uUeyCL4beZzURQ54b0
QS9RTMSWmCoKEcvNiuFPov7b4KAHe7c+5GNAtDuGqfCQhnAMqJiX0RzuexTqdKaR
2XS27FdU/vxC9dQimXeTknNhKrpPWh6fm7Fa1w6XkbXkQW1gS8mqlPmZ2L9M74yh
gxcqKomlFzAZey+kOtuj2jZHojNRlpNBLq+lFj/tFk4CahrruWGSj9CZk4Ce54fo
PHe6Qdg/91okYJr+CPkQZK9uZ81iQL9UgrEfz6iE0x/pbDqW6OKWyj0/sWhY1xfx
fLLlU68QihlE7qnVje0/6JQgv5ZvuarTgc6L6OWxJz0zaQMLzAt7o+HH8QZELUcT
az2rGoPUjOO8TNhegOG5002R6arVwn1WlLYftE7BIO4PjUald2SgfOgzN/vSHFyK
oc56MEoY1dwL7lAaPwOOm0+PPMkw6eGshdg/R1BsQa4A9VFvguoyvwEvl0SjHR5u
r/pqVQF4kTbSzhqxMEIZ/N0GmN4EIExeD/YF5gS92gozU8WUHyGlzcukclPemdsg
KZoZzQRBm5YEsgHdcFPp8Y6WpA8v64yfjLUtL8EElmS9X4Tqcg4ZnTOwe2pK3v1/
msqwKSOP5P6rqx3TiJHhsBSA4O4SjIRIt9WcNis3gTkQo1CaqSUJX7nWalwq56xu
ciTmqapyZG4Fez0GDjAX0C+6sVOgjDaPk3JdKJmpq4wtXcUJeZBp7bHYVWmwQXUd
fQb0mc8g/lENx/yfwnPPy02GTVNmn5uCaN5jzzksV7xda5b08142HFyy7scKA4+0
x9jUc5OAkkv5Qimcj7Vrt1UUlZ3VwpleAIvJl5ADzHOBI95edY29cVAxyGkfFXEm
Ps30zJdlxzLT5IR33HlxXThhcuQsnF6ZFVlyz/j9FR3nfSLESY0x7Gs8vHiNNp2H
3KC06KSy30Hjl/j1hlVJMB7NlDKGSv22uSCzLsflTMwtaYRipuiUSwKJ2HqmXVgi
/fI1tQ+9WIkr/fAvxniOY/p7IVZArSGNc57+d6eO+hs++66Xpp/T/8Dx5eLHJmwW
0/LGXexfUq+qLcSWTBYYx7bR5UwCeCCzxPHMyXPZkE3Qk7hRm7jlo8yRJnLI+sIg
MLluUab/twtXNpLVEYCuw7Ha5sUdUK/Iq43e6ElAR2ZBHuEnYvseMwRPaSqloqJy
nGTiGTAdPLMh+A4O5tuzXQN4MZL+Ep/cF/UVoYgJgREUWowMi/KdsTSk+cVxoxUu
OjezL0pH+IYmiWoPly4v8bGa5boA/yrkA0F48gbu5SbDnt476mv3wmNvoEBW3YCH
zjwxV1Zp/90Rvk+cmrchN++2dGhqzQfl800U21s/9bX1nAS9QGd3iABhcqQMBI7l
2af+3A8ztrTPfEPG7aNd3megeIuC1NB3xAovwUdmJM27F8+aWNlfbeyqtkRvEEPi
UFDkj1Ss1P1pFrin4pNOsQOidlYpNqJVAwo/BQtQOi48NZEcMx+Jl5EbD1HqgYEn
jHHLPO0q3U2JZN4U7lqFkt3ag83Gs2vYKzraA1Vge1HBudxX9i/HcC3TZgb6kCr5
+UVg5df1XIVHbRd/q2nIVZ4/KmVrG4zJWj9RfGa5pAx9mDXFlPJ/tH7dmD6xiRKF
T4j+G/JXcaYAxJIzvHEIFC6ADC9B4ew4S2AqfJebWl8ETUwzGiHM58CFIrwz6MBT
44RBUIBu4dLid8YwaJXgy9fEBY2u2LZsa4VVBzQoZoR5GGbmmrwwca5Dp03eGOyp
wumjr4ENykpmiWTTlIbcnd/A4E/LCiu14q7p7DDItcF6aZEuf879Av77v9tvqo5u
JU6gP4I8Qor3jCuvLrek/ELizpNELV4iRHVrZ+FhIIoiBL8aIBnWutUtnDDhk0oi
tnWfjXhDYrIiADoGZ5rr3Of1LnDT41nKUkmiE9tcvnJAQXthawl4SOr+oMdHs5Pa
m5Ovhz672w1KVD8rT7EWw7acF3fe0DH5JkdFQkeu3R/j6X+gx8ghWpYWwqwuuhYq
a1pSqgJuOAFDdy4bwmyhyZzLSiuwS4sMsLWOPe6tI0DhI+A8Ago9sp7p5gSIDiDJ
/wA2Xmv6VKFcNw2zhyx8fkAae44rZxvBNgCCpriC5jSKQdOYcXuwtNH+nJuIZvvi
R/0mGdqJww4Lv+IB7simL947zc9r1mk1to1tEuPGSVg5sM8VSHnabekxxKrBE+wE
RapF5ZeYuHzajBGLMmDGpdEhuVEsX8HF7XphnMKE6LH8eDPtYwvuSubdihUifvxc
zoMEtTvqJR47286BzhPWWRFSfeh42uE9rdJOkjcqfL7c52AQnngayzSQQNOSPVnf
UATqVSs+KPjFsHQMWXpDZel0z9e6Tbdrv5cJiTKtlINyDGv8CW8reLZveRWZ3fCm
JEWjA8TrMxiCNdyPoJJXySrAL7EaFpyvG+9n4Vp6b1SwU5WesIX65b5LUoWNQ5N9
hg8jSStPEDB0+1OQ3UqzaHyrU1XgXjA6pMjsXiXau+F/BP38iQVQv6PyXZ9gV2jJ
6UX5RrNCIauqXZgXn16UT1xlnEVojWT01qEzPhEUV1U8YpTpUkP73jJJ6Q7vvFPa
91kUiYZ4AEYrBz1PyoCsVjLeGIRUi891+4DptdhrQSjVXZPByzQKvJ1/CaiQ3oU6
oi+QBlbJB4faRrVE8/MTF4WdqBQ50qoggtKvUlvQ7HwIEJCO32Q/v7jLtQ/q6gMM
U0D40xkm5aNzM68RAEceTscC1jRJgsCDtYasWLqWUmsUdjY4+wOP7OhhsqloVwN1
FP1wfWCAcQDktAeLNtkgRCNcHYJuqQV+1mwSIiw/zvyAa+zoti2C4bWrBDx5u+fN
MRjbT4oXbAH2p9Oiv7I5AnNrR92vFDiTAcDfFwlf2bj5SYK/LQ0DLC9RF+C3TRZB
14aZ6hrwjw65UJZQaSOaWp2KTe5KwwHco5Zto+1OPXbOBH1He7iboVcgPigkjO48
KJPY7vpTTY4nm9c5q49n+uk1z/haNiIA+aoRE/7xmYeDioFxogWzSz0TO7PNhSwz
JK5XthN20Xtk9yaQ/W8EmXQTUAYEngpAksdbwojB6fQ3hyZdtjRPL5v3fUorO+8t
C5vFJ9KQa6YcL7LxI1IPhhPIowe5C3ZEhTIJjlWbaTr6Kb4vfeHX+fpjBfRGSMmE
0V+fAaE8Ef9kMmXBldkH0COHd93N33avBg6hHA6JH6sUalY89qmCDjiy/o6g/baR
mZZegS5uTehaZDb6bPSWyVZJ084quJqBsONVg+Pei1y9vIztAtvoTCd42UYa2XwQ
8uOBclz1HKD7B0DwsqdujsEi7bEMvOhNURVv0LdVn3HMyx965PMSzitSBc2dmDL2
1pfc76OW+LjdA9V5ZHbC38FsqVSvxH3P7Dg9r/sXthhMwME8W04KZg5YGqG3uLR/
+vRUDkVPy6RMavBq5FI/HTtkUXHkz6emE0hl8e2GIbgNGezSlCNM/RPMlZpOdsuf
XZGRq3BY+RSVSEc2KLkIzCTo5mhyH9TShUNRg26/GfUxOLsFNwBIZLCm30LxRTMc
8NdBrdoYqY/SgaViHEfVat3M/R2anNDV6ZQn2cy4WZdIU3m+sLYXl4svVfSoFOxr
xirrQxG6SoWR6J8sfdJLhQUz4bVJOZVCihKZ0VlyW0dO0pTJtqxBhLu2cEH+M4+n
0jepIk3Y0ae1wBnXQlKF3OafIjWu8aJffdWzxp7SRHza7YVjDT4WphtL97R//Pfx
bSh1TWlagx7F849D/J2My8gTrj5tlDKSE9Ssmj5qCH9kWb3rNHbCv0SYbkjTkV7G
IhWVrKSyK5kLAhf6IzpLnkKesWO/rlZXUTSo/ItcPlccdegp41ARnqAm/KYgBLzV
2ruWjZXTmUce7CIY2st4e0qq1RsvQy1q4kAih3LsgkMo/6jPXBK9FyW0seMnmyc2
oG5E2vt2HxozmPV4zwthqJu9luuko9RNUB42TDkEbSP/UaOezvPpOhGtgphrugSR
KuGj88WRLoxchXvMW8qzAXWcP/gZNYbSudHtbFtVogmO1ockuUlVHXFXZqTQIlSz
NKQo8C8UNG6t+IbVCUyzNXC3kMDrjQ+dF9x2NuXoI/8FVinuRrfNBIX1ys298eS4
QNr/dUpDq3yjSe3MdNWwZHFMLqZ8X/GYEumeRmZaw2bhpxrkpd0l0t+Omsl7iKzJ
KXBGG/r5eM4L4uiR6ZKdWt2egKkTc67lCMA5becuZP57VuG5QY5Ub+vMvsioycUM
l/bJwwWXG3uvmr0EVictOGbTZKaq3dtpKJVSH+QZfbWKDoIjqh83E4rEGTP6ZHyL
IINsYw/1OomG2nWbuqDq9dpUgbQ45U8Nx6mmoXF13HjC2kOg/FmjIs29V13EvA6R
5ti8PMtChxH5WeBzLVwn/Hc2ipfmRLUmzpV1prHA7sszZidDBeIhryoJ6bpvvwwn
rAJct1LyfEwA+JQqCKynlIouFh6X9rCNP5mlQsP5+zRUq/SCiq0xrVE9l5/9mnRj
eGsI7TUcCaUpIbcl4rBkNnPY95CNgQ39MAcy/RUlYrM9a6etDQZv9admkGrJ3oxs
49rgFilKsXWOxw7meqFb42hSgfHpzN+1Ijyuh/uxdHWxyal6If+xMvO3ra03a9Xo
8xqr1wZLwYrefVRNHOOMB44psvICjVOunMfMfEucVMaJGytLQg4iRdY0dsIBeVpQ
5dIPJoKiIZb185+Nvz1NkzovlJz9S6GfEntKclPVqZS17eDug7dDR3H1lGAx215J
slVMR54l5/Xi4Fs8P3AfmN6/B6/cAbkl6ZIeAZvgIvfTpy+EGtYKfsSyvvoVHpO+
w98uuGZLOJxBElYBc1aL3v4Cp7LxZRIv0Cy4kswFvm5zXWH51mHcdMJGGpXCgvBU
LdXMQakmSn+iptaEBEaBcivXg4whFkZIs2Vu9hFPyKzVkFtXuLLY5eQ6+yYXjB7l
+cEkAbKcVypDADf1ealqHna2WNyHD+/EaU4Cw9ssp4SLXCWLTLOeCu8G9sSVNwpF
wE9EINsB32G0eZGmKTrUnfCJmiYbuU5Yuez8px8DVZVL1ZJlu0OZoZ3rxLens849
Em02JgMCl/WleM+aC0bgFEZ/qlqN9CZk8IZbXXp+Rikprx6yNu3KyxKvkW9doEIT
FwtgJ5M9DBwjGazYHXedvKU4RYStXGig64+lX16vKn+fFbvMfXJPxPEF5YBDuNmm
f6YnC9BmTmSwokQDoBgUOvIX/WKucpBSRIa2xpn5g1Mw12D/fqaZNf78n8Q1avU6
W7zvI+FimDtkc8pF1C+jA6HfRGCSH+wynlCNjO9GHjhSoMyiUQcUFXcwvhs212MM
Z1pqF5C4bbbFVSlQkJfPaPuzjgtIbAVwUGscmPdVOq9igfMr3v0E7rAkLF1i1hMq
lCJcutqEoodUcIi1So7JZoefIwydIfb4iPNcK+FXk9iRd3V7mfGcZy63VBPqqQdu
Cvb1+iM19qvD9GgJ20xgZoaM59KK5aXt9LqTmLWTEzikTBx/KxRzSxCDt7re9QvP
wlKREUeG2FKk8hyuAqcYBDPWMIRyJmjhOe+2PHQ68CtI3bRgdZUPmDDDMLdr5Kfc
+P4Md3wkXsD7VJUSF9aHWNq9K9QEW7hirOLHTWGClWX8N8FBTdnTETtovp7o8V/Z
2lz44eEikvd0J48Ki2/1dpzLkBAEr+1b9TkcdlrsO7ctTD1miJBs1LinDVUolgvb
d9MHcrJjnA89edLFyFFBwbk3IWB6FdRXJypLcKvyv4SNs/bx4///fBttvbRuKEE/
44cxilEuPgtVovBY3ed+OmsnoSZuwrek+z3a/AW2sAaBnaWz83AG0Nt1VqeoYBOU
3G8TuC/OrqFSBJoEY+S9FTYiNLS/YUcZT0VKlcNvwlfub4e5nphIQoJEp3KO6nKc
RU2rE8HGcw4OUyBp6hb1YQxIxbLA0Pio9FujaySko2gb9hRfna8XpreWWX6HUlmr
bzuIP8TFIvm7MxNdMFZj24SPtSeIS8CP37QmvOs9zKy4++xsO134jd06BpqEaGoG
VnnnYrDSyFUWUK3LWeHUcOcWZOS0e4eU/cijtGctGsmTvMFYG+cb8+3Ie9/kFpUj
rMJQ1Dew868wRDvSKL+3B400JLqTDwYtw2xvPUTk3viFFpO26umtiidtdWe+JPHX
4zbtW5cjldQqAGMNXJBYbPojosjpxts0lkwwaCpV4VgxI9TVYXC/mNnz8VHCvium
yU8nq70sbIYvGe0oJxQw3hFpsqRHuF9SBoRxCSw4sEoF5In+2y1FfePqeJGoiO6E
VaJfcDrN5ICFTzp3UVOIvTjFejz5Tq7OpTlM/vwa4zA+BwiR+7HZexB+0u4Ia549
tC2IId1QE7ERuo5linAX+L+rSHGysh+kTlZGsAE/o0q7LFYillMIn1siz5Olj/yP
GONkY1PU6MMbFfhQ4G1eFMzzWrezZsfdqWbVJ2I3lc4zQPxP0muo71L10571rCLf
QLggafofqUEAneWMzdwUwQAUxLhVhCscTCw/mQzNd8dAK8rSRGWAUPJDtS8BeFfk
nTEa71kCpR1zpoGP6RgQqsqw18qbK8723nG4IS29mgFyDIZv1Qf4ytR6mro8EpbQ
mJOLwswaYbphCMIueh8oBejEtJW9lrRnGhOrIezbg39ZLc1nFCKPk57WpXxj9c8K
PwcRfyieSr5wtAZiuCZmytY0SNrv8wpQTjAAo9dCU778qgkZkGfob3dFnGFMbyvk
uplswlAmZ7eP+h9Y3H9AhD6XWclh48EGkwaThjHrV/xSuhc5Yr75YRIaDJYiNIIw
HTgEtdgCg1px9oXZsUcj/LZutYDiUB2yr4FzoRMVaTKDrbcXn+74M+NSFKY1tApH
RZ2gFUxXF0u49UdTa71PWSl4m6kyzAPnH0fPA1jtL2zey8FMSnm2/x15IA/G9aIh
KT0WJ6QF+wqE/d6XAzrLGQj3Kgyq3lNHHiAvIArzboESwJtQ37uMZG4XeMDwaBbN
eqKxEaAP1z48fcQRwolUsILUm3mV5jGGDmLfJEtjl+r3yBHxoJ6BeuJW1Xi3NkGI
TD5StrQjOQE7LEfZhU4f6oonwrylF3L8JmIU/l0HGCV2dxgJ1VxixCZ6v+bdjTrw
i4CNE9BBeEjPbNfUxdtQul0D6iHVqebewifiBG11ThZWGAXCMxWsyDPquM8l2gZx
CMp2sKcuwyghQ+CbtxxKZe7wLF9OCBv0R3xXnhv9f8Z18p6VpQcQB7UqmUJ2sUA3
xQyBTF/l5Q/+A6y0+mlnJNTzEl5sQj8FP7xjTcvHYVpkQ1GHkqydKLqJSGDD+ZIr
hXvpFk1w2msUwVgK0UGqJcRcOpCzdcGUxUvE6mXaVQ8xu2waWq4/9TDHumieAZC9
mASGF4AfWJO1fEg1hddN9C3P8eb09rsSVRNBs1ngDk1+BAmW0MJQIVqMCONhWhTC
/qgvBK1HYXQKdyGkWC+jIvhaTZvlMYXPnN5zRSl73q09cMfGcqX7189wMSW4uJcy
GKlwozmmgq0baX3OS6OCHIugpP/MO89jVKOse46BqSZXenR0+6RumM43GP31oziM
hRkSNomSyi1R/VFpI/wisUlhbQCp73rY0Rwu/JnKRxCkXYCU/MCWY8RWrBlUX6Zg
6CsY/Z8JU8aWUPJt7XOBcUHOOUGyUe6mSQ1iKrv+QDsTjowRZU8ESKl5soQuUMPu
FVTjORoL71RxsMdY0US0Pusx4/ZDs+7QcDPP1pQJKRuEuTpyLXVbVPQRqraNBviG
hBfNWoMnLnwOglAbrqnK4DcStpzJNhapAyWwt1K8lHi+Nazc/rE+oFnFlxcfXV2F
2jpgN6EF4ApX4BoRi+IcIjYAZ6sOW/JgFf1L6nDhK4YGZHtaH1Ke0gKWRVx35brs
dBVAtF6ADdNFexUY4uSbgZrK0S1eHdBw2b555DUQORKh9d/13pBobImZZhCiYIIi
P0LDLEhEaM9MYBxDBS7w3Q3qkaGNtmTQ/urJYmNJ3BY56KbB1sVv/mfXF5E8P9or
ulswFv38lP2G2yk2IppV3R2IsPjoeIKI8hRp2HZI5pzVae3v89vJrGE39Q3DxPCV
ayXD5HtISqs9heNMuK4IaLrcN970B5DoYvznU4DpBHhKBMInAZFEEl4Pd57LTgIX
uaU6QYrLU9qH2PdV8yw4w7tI+WQlZFa2T92TgPoik8RAMg6ifXc1OdNjvtXTc1q8
SVU856HYx1ZUjqQJ21reuEhvEyk+G4lc9wUUiv20hrxQE9xABzAJYt3ePTel9Hxz
MNWvLZI6vJkA41KzeWpSM2M7HY9k7zs8/rhLTAC4tlNkT73uGnPCN8HUF2kKQAh+
ks2ijvVLuWzK8TRxV9m7o/s0PP6nLWcw9wJAzreIdbNp2gScHJkIoSQ0tcvZRAIH
LE/6Nzb4RqMHo6qi5SSufC9tWgP/nh9LY5HlCu1A7x2QMNT2EgSP/g7h8Sb90oGz
Vh5XhweyPx96eCXvlmPbpUIyaoZU2my2l4ioKTbNzYBz8WhvGbifovJtiZI10hIj
YqSA/1vLVERDfONXYkevJ8h/ejcnI231sTjpQW1y1LbIqxvIZfgODwU/FsCuI9oj
6QCxR6bTPfIOFhfkJnKBQuMQN4PzKeCcCaWws/Ok5Fv9441Iz2NOgbx91QTZ0QAB
aNNzoiwm5ep/MQ92tf9FH9RGqKXmzBROJ1kZR8t4Xcn2fBY/utX1e5F+lnIhMXYh
VXGDsXhXxnSZAm558nttMgZ2kFx6EcY/CW6fB8uwtnSVblBWjzLpkqAfMd3iC+Px
iCRvvLFyLe6VeSf1tYIu16IXpCm9w6SxG8tK20Eqd2jXbe9X96tCrl+v3nKPRILq
XR0NIYCroopoiAqRhyN0c8k5g7cRAOliwtX1B2tj5AWILlejkE+0yVbTwuBq53bW
+Ky2Xy8WdB5EgLwtaUDb8ZANI6fIs4uwH0uTXwF4edBq8tsaCV0TmkIvHwBTxEMU
nEdf04wiNemIUWhaC3QRVCKa8nmkjKPtXCZHslCkcAEAyOjgTXQX4pr2QSd87PCv
8P2NY6NY8a/NiYAwV3OcmzSmpysMWftpAZudIwjR3odItEXMlbydVHiNRo1f7Ska
TDnLkZAuV1za/m8gh4BRZO3wvbdKZP/xYllicQT1ZuzCUb6MvgsgY+lltZDK2/ob
z1x0X4YLIpdCtdVnoYwpvDp5hq+RKTrzihWqVf/D2OmPTMNF9Scq8+AsHgyeiGAi
NMhvoKOKw4QI5e7QwGUNPy/TYLkKMZzxb22fPW4/bY6scodeKudfrg3zjteOH5O1
837V0bhNdq1FmyHTu61a2cb0TBklHjxO4upuEZawfaJPGWn1k2jptYxMHzlbe/ew
Fy1qx+QAhlQar6cpBqEFMN0NR7EJacpNuYVRO6d7WrJYkSJmwWiTMmWr6NN3EplG
jJ/Ocxk6QxmRK53M10dpiUroidsD3qL+KOkHMt7xBVX1sAXesTgkgMd57qaYDrYt
BRT8bXWhe2dcReW9nFCobwaLZrosndNG/hrX72q4SCqN02GoJJQAFZPRURYsSEY/
Up8rmFK2E8fEKG4Le51tKNv5opg6DtcahPnLW19hNtTSIIIKpolnAwEFGqpid8hK
ucWUrpEX1NOrch6YCIVd6JL6cqhhpnAIbSmZeObr2vga5ovELA41FSAPNG2nWwXa
sBn90W5tSmjyza4kDW174yKk6duaEFoeBuxrtrW90oPtodhT6wF7iaTXcUoGWS6i
rN4cCRjaFh0tCvSSHQgH7ab2DQj+1utbPxynTMZo9YZyBuG7rjgidFywb3alhuzL
o1Ilz+PNs+3jDBg32OIWW9xghfCmeoD5iYvm5mEDddXcgCWnWMvNjq5a3V1L2JIK
CkV8g3Qwfxw0whvwJZ/T0L8ZGotLx8FoeVh62FJqZHTyAKij6A9VScPHBgvX4ep5
DZVK/7nElVWICmTuvGSuUnRWTWq4zaB5rxLvkfqCgMSzNyRFg8Ng7/8tOLvIEUmb
8KEgsPgRGtXnCAoneYdY8UczVmIcl2Fy1hDBsKTTwgmS7hxEYkOUY5hGDh0uswIg
z2RD+CHaF6NILru1ZPcQvOIauRRRlTQpMKUCHvjbidh4WmVjiws7KQsfIrgydhMg
RnxKeLKZjO4lb5AQ+PFX2tdLvQqFDL6RZB7aZAxNeRhwbifh77Dst+s6rM7Xst4+
bIbycFEi4wo9UVAFbgs0K/f0llIw73GTbXNTrJiMI/CuqE7O3JXUKeQymAHaV6IG
Y5VifApDWaZE08cst0bdHlduC9XMN1lTRnPKtyfdBdlslZrn9AdYDTf+87VVCrtP
rLTpeIdhGnFRV3Qxv11NFPOG9mhPUA89R0C+aJmn4PrH/FmrdXKzma+JdxmwIilu
jGOi9thWqzd2RhFRA9uv/bw8BzBb9OOPx1gnpCTUcXeWCGl5F4wqa3X44YWfd6oK
LecrS6zJQ+26IxLhuY0QgJ6OPGkA9gQlPiJoRx8tRaCCB/3vpEFWzJ9jrwcgNOM4
Hh+w1nz1OhxIeryNgbMf+1BWvnzSHfdrAH5h+lnuiXZmYcyoPz/u2ZxxKxFq250n
udxXWamgH8u+gOsEaPWfg3PbOJIEp5bEnLCRgHEaWvNdNH5zSQ6151U5ePfKcnvh
nSgvlO3bPe47s+6HJjfDl0qGjn7C/uNZ4fUax3kwAt0NlXFDmXnMsLQVLafe1hkG
+9agWH4nnArnOTN6x2iwxDWQF1oyUWtNM8PUFp5+Gyn6N8BYDSz2Za0X0LGSUdvB
+3rc7PVm7swNAc+ZpFn42vGIJpO+zvpQRoRObmB/ljQnJzLqV5LoATPZzmyGXAwQ
NUawVb1XB0jP9V9KQa6gS+Hu6L9DtobRcalslAKcepMkeD7MXxl/dOt1q0yXqVoE
sQnkjpXtXpElxJXKjSKr+/20jrxIA5B9D5MUqGLXzSSyRtCtIuxxHH+UM0pyV3L2
bSLqzBqaP+pi51g8wRs/PJE0jcauAmW/S1H1yjcqsiboPYgoaRQJqWFhS9g+Xuct
KgBkaajTuXtK946AYjgwOVDklyCdq5QZ73k5TpKRlogBIsOO09OJVNSmpMJkoUad
9DgD45W5qGQ/nwlkaJW1nO2JiXuMUckY/Y6CUXqfY4mmW2HQNumQdyZvmT640xps
Cze00NL8Ku5/1y2JN/8A4P6eaE3gK21zl8C/6io+Yrddv0i9vIkmTg60H7ZcMdKE
SpP2VR2QorJDrnf6jRYvYPa3R3sz78G4+XiUqlz7l7DF2xLxYHjGe9B8CxEuEC+3
hjLycrMChTb6mi4Q2YztRd/l7s2MgpQOva3EcqG1fUtAs7hE2+mTE+yW9T3V709V
eqZGyF1A0l8sq1qpljj02DVtRbtGKfe+C2HzpNV4Vk5ABIOjdaVuj0dvf+Kk3ZEc
P2r5txDIkUEPNy5gkyOn3MHuEuEA4deRBCyrQZAjdfq38YMXoywwL/cKN6r8l2C+
fZem6+XkJg70R4/2N4wiVCzeKsWjxyl+FhC7FDbE6u831bmsks+B/dcKF0gdXRLt
2JNolfvlxnVHGdY/o5ZpoCRc2sNj8BHeBIo4vjRmB0lSIMvSlr4TelD6wp7qfFnJ
7uh0QnbSiC1LpSy+0TIVOs3qfMLERvJKzgGRuZtr1yyrA24MbB75xLLcRPNyG5sz
tL/Tqr/4oYvtQcMzsiJCPLo+uisKTFH+FCwjIg8nI/VBDNtqrqkTqdSCn2D0wZfp
O/Cl1euSSG/vCIdzkBYVS96oqAwHg32PLT+f7zQasdoNbEfpHO9mEEeO8KwJA0k7
TO42P+vzxSUO0qDY2v31aBW6orR0mdXoyTLMraA0+oWIZLmf4dCHum39pGLzbxmL
VU+6ZOCOXDnW3U1Nuzmu3RWWLWquiwiFFaWtNj30wUzvHU9GCt8XE+p3TWqy5idT
poTpFGj2mGCWuBDtMufN63iRO+KlLQlWJ9RSqV6o/NlvBfTcpL+x1PLrH5729HbO
/raAceNcqTuKJevzKlfsVe71Ee2Qj9EB3mI6pyr+5NIig/DRZs756CS2cdRtxRWD
61rYYjBPfQRSFiquk/UWCDOEgeWTQEYbgY417OSmVo4ftbYzEwYOrjeWpXxqF7+d
Om5gfNAAuCXTleubfyKn4/SUhj5gNCSI6HH60vYPbb+R/hfWQo5DBp5xX5oZc3QH
bXPZaxoMR8XMhwcJ3JXWotNA2f+IBYGI70zmLl52HA/kU1Mr1BOW5DLNpNsmDKmg
XHAsBpO6wdYxlx73KIHo21/JaPuEUcqX30EgPdQmvAooG8TSoZy+ZqTbp7io/v0u
fuSoTZuQEgR3YEVtst8bZEDgEIX2O2vJzxkASIWFlLF8rA/W98Lv9RCsosw47Kxj
7r559vVRI6QvH/C/apvID7Ddkqb24Y5ImC+VLl/WlL4ZM/ukKNW2hmlrxSYCedbS
HFWksyK1FofznZCLtc18aolMXgYsbGWLGuZ5cpEssnmOxGl0j5f0vdOmV+tZgQvf
p+0iiwX1MxuA6IvphcFeTA/JDp6Wnkx+q8wVYFEpsVtsg4sQ3EHA/Ul7Rz/LCW4V
FQNAD+4/1RfXlt2VtX8VSuA2Mg8PxM4jzd4IWFBmgsTWKC9CokgPKjREgQkeHXx7
xRudiJLvrpuxgeS554E92jztT4CCwOBvFUuC0s9JcSqWZr8uskwvolJhLvt5QQhq
BNCQORWNWjEGttXv3/ehtoZDGgb+83wRVlUat6PyP/26QbTUJJzPNU12QvNQn41J
0fl4Ab2yOKKSWNvwvtDv0CNBgu0//6uAKY+mmMx+Um6DNpa1cHWy94FTpa8Xgnlu
y3B3cDdAeIlGZBNk/WqZSDyFLz3lchcNOX6IE2AcQ7KX3+aWZaWCyjyJOF/VA+sD
thy5CC7ZXIZlZV5rY43UGE25FezdB36j6gVjy7/FAzmTVfmUyc6e3xVvD/kRvTA3
yw6M6fdEJB+6ttpZfMxuAefhulw0K+KCn2OEB99v+cqeuWb7m8uc1JM2IXCDtoFF
EsLNr46PdJOhtaQA5oSSanqXxVITMNw2sxcPd2SvKkQoz7gT5R/0dTyEXTcQq7ff
/6M8EZmKf6PwNFaMRsoqZLfQTUpcGpHE+/IWw+pfiRgyEhgsrhkLWZ3qgHIe+Dvn
yrdV/vHXtmK0Vhibgs9DGg0xfzOI5uCKiMCyrH3y04HplIToSCkc1wklRqdBe/xe
/EjpOLTVCXsW66Bp/3mYP1+lK+eLE1snt04iFCzo7dsu56QaUKVa7xVu2qCUUqVE
bDBdlfCzhNh9WuLaVIug7u4xXU4PHvycrMRyNh/Qj8ZdZVeDSwplaobCHP1a5klN
bsP2gNoAe6A3EDcvf+7l6a0f6w57MMa7RDMjl+OAOiczmhchrwI1O/IHmMWb7vjL
9Xf/0/JZvtKqUJGyfbCAuZw2YCkIXAI6rE3VGnL2exo/QRPCaf3nArUoiTuadRUm
dVyL5S+ogmgET76VLUFM4yzu+xJjurujLkBYiCYNEbuFGZWLcmoKsGj2oXW1Grmi
v7sD7Y05ooIcAXSeMafWd2wmdyVPnuOsdVH/0VrmWAzV0BJ5R7tsabSvUY8I0hLW
pFbqv15oOpLaFr6xAazl6XnctQ5AOqZtTG6tRNaBL7y4RgoT1xkRwSvKpksPjbP6
gAi5IK3f75lwN6hdoT3uF5VO25MS0vCXTNt/YW1NPHZ0xJG7c702BE62MJLKukiY
N+SS+J0JAMX2swIMKQjxZS/IB9lRsLtjjtJ8Ovbovdb6G4tPgiGeas82/tsBEWVA
036ptqSJ+C7kC/Ry2SXWUkT/J+hopsCet8bM0f10/SuXhh1MhF6egP2WbkuHFC43
7oGXEpZ/XgsO1cixhwSA5ujJzAAqrJjSmYTX/LHgoASI6Q77VUtlZZHCe8JOn6pa
dM5apjmZVcVmqqD3VF8GTKNTn97E5lEjEJSBhKtp/zWUe+ZC2kDyC3iNqZfANchb
YrUJsuekfldFsTwPoZ66dmzH6OJkS/XtTmYcSRaE/IylSXWzPPxdLZxlt+MUtmEx
3/r4v+rl0biZQatxsodsS5DxagLHGnKkzgDHug9WHfDGWLGhYubWsfXzOYY7FeX5
wb86hnTFk/ed5M2NzSiq3KGPjjZ1vI552xflwhlCjfAppS2G8bZjA39K3UgqhVUY
v01gDMWErSjuCy06Iq82u8hXVaGF/XBii/IsVM8UtoMQjw6e7TL0wheoWyLWTr1b
0CMvY/YYEMju15FShVa/0uJziyWy4TWdo14tNlAwt+/jT3ChY1mb9arz7RTXpmWl
mg6VvGK7O8xArD45hyVgysDVbeudnCR8iVSitmoEt6uYJdRD50Pwtz/0wv5vvdWx
4CQX3vV3yb3n5/CLSuPj1KTfFEdWU1K3ahVcy9BpedWIhmXk2US5KlUginAS5yqJ
aEE0kq6MHWiMHfYtUxQBNPuX1gnb59kJ7rnuGAxPgUz3yPlTNaCruG1hs1t5/RO5
HO7t5TqLNOxGoSKtOWUsd0LI3yi3FQq6ccuuuTw7rpy6Jn1bo2kRRp3NWeiFPmA7
yAoEQ7zD3/VmErU5rvkwsyCe6Ugho1NAqvMbOUmMFGHGNVtsAxItgcrcZsRD3byo
Az9+Dknwj6CMufbuyJcWTAYghmJMEZF6nX63xfnE8uLP7dR969hNePqbrhJBrXur
LPfToC29UWUvtIoHuITuPZNeQs71bs1V6gKrVMcbVbI=
`pragma protect end_protected
