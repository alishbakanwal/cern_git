// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 13:57:46 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
oa8PPd/G0A2+FGl9C8ZNXDUHPX4LAv70eQ0AXRaiFP/Sqi1RaYHKCNWIDME4nld8
R+MtQSx8b3lz4aq1vQ1Ki/ox5+sHfixD/JWTtCrXypeNKSxX+JfTgA2g/t2bWs0D
4HFi2Z0EKFF0KJcgtztrCuOMuGww9l1nFAAmqT6N1KE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 176784)
goXRcsnueHvvjH+/NAOocTfVxkiAr9PiuG/ug0R9ezrpt6WtlUS6tXkIfFZFfWy3
DrKBJNVeIGTiqExHn0RGZ475XmZF6aCYac2Mzv0L8shD+khSuwayrlxuK4jyJCWc
BonMbLUf9WvLJMWUARnrQOw3sDkR1tu5tzm70+YqMgVmZ6pxQPtrq46gtA6QhVAZ
FoMxkoxvhJeh8Xjw3pFzj0C2+77vbtQWpjKQ++YTItFbpTYFCeBKj8L6jWvU9TIE
Kyvppfvvc3BrcG77GElCNAg4pLt7LUIG0lnTnr7a+6dU1FXXBIZwjDey2KWvqltl
8VznaWs1xIWEFn8RAROkdCoI670pvMHrvQzT1YCIep0cjFvM8hz7ee8pS3XZe8u9
9DqhSei4A3Lui6MpmFp74g5JI5jxWg9fmLjd4RTURkh2xu1dYzYiueHZK3B792JE
cg5bkYJYI5oxKnVSPoG1A9+3S9J78Va19GmtzEwKoEmDsRx6vSs8+IwXTswV/3lo
+pK5VvFgxCOcNJwxHgkl4pqN5t7xD69lT2znFelsnp6xBSoB49frNufGHEZOAZJJ
AxzgN1u8xovwe3EyWqqOnZ7QSEd+F+vf+vIAPoFYBhHWO5J2SHCl9U5w0ePwH34L
ttZEZOgdhd74WExdDpkJn5sSaA6t2S/CTX1Apc6UqUruOM5C3zAj6+FfozQpb61E
hFOlmJiMV+rcpUNXv24ruPc1t1MJGrneZKc2w22pDNoweOY+89J7Ba1eOX5Fhcwq
qH//C8ABna/fklzHxm6c1lV8LiI9iv70iseQFXUL/F/m04YxziilvqR9hdnIyENx
U1yF+fKa3cx+J1RUqXscg/EOW+IUMCK6+1iGVQD+oGhy2Q6dUXF9fZ5G6hclly/U
xUXRS9A1y7+PYymlp3DGXtebMmCx9Ekybcgqgf1IG74SeeykQNzmeGjGuU4BlNp3
ePDN1dUw0mSI5Rdrg+DpOEtrVNa0kyr6WdTp8iY5oiRmXx/hUvA51peBWyE1Gp5D
7A0SjaBOwJRnPQJBm79EhvbufM0Kr8xnwv+pLEsE5LOa3DQC8zNz3knEsaWIAbCn
ZaaaCW2S7Ucm5mpmj3vSN+HGmSNZdf47wZJlLdiVpNte0oPy2DIiO3LSOjqG4iHZ
znRNsM9HQ2+PmlvXO/F/5OK0snOXeZv6Fbn97U0rNlChaZ3TmWM088OOCdMSlvZK
4GqtdciYb+YU9Y61y6CdiHyTsj4cPwwIhSrowGkdad20OqmxoQ8digctdmFEmc1m
PW1Bb/o0b5GDE4RBbc/hP0M7JrlixVXN0k8sxke0qKbTjhVq7+vR2yuu+zRQhhdx
UgxKpXck6Y+yVXhq/13J/cTR8wgdoWLQuo4ogHva1ed/o1V0GStruj6dJ70TeKn9
DvSDGK2acULhSc1hLeh9LIOXCpUf4Da4EZtqqihw9EkQoI+gY/AnGGZS/vaQYeTR
HfcS3eSTWXtRy0HfVd1TrU7OsAWXkK6Ep+89EJDMH4DGi3/Zu4xy+OL+RPK37b1c
+NGDCBDuTkCCAVgXfymNh01/0B4eCV002qaWnMkKZTerJRdcNLiKS9mJbAkoU7p6
OXxYFpqmLPeEHmmlGF6rOJ/xn+p6UuuqbPSCLfatXppErV5lji1XC69d8whf7NCm
IWe0zEB0vQLJApJtvZzntIHdmISubIlpZs5jMOY3ZMfkckczwW3c4385f8Y/nN8S
q8nhEyDJYrA4GbtpyYoValUk5xdbN5HxFb0BDF3+nYkbff1wUA1aVVwZzmfdE1x8
FWsRdKG02ewVcWDfZ/tbvQ6GiS5Eqnec+eqowhjHfU1ktbIf6JLhvO7wRecDS+Je
L2hMq7WwZmk94Cf4B096UU8WwHjshT9bMlW9Y+pw/vAFYx3/MH1AZZVP33SWZIvS
Wg4qG0CBfwDMNC0WKqAFZryunk2PEg4ouEVQpYMPZ/HhxLpNgnOpSi+e/+pwtVm6
SpDNFalin5C2VGA4hkjmKscO1fNrwiFP2+Ly638KnxhClgSFZxnqIx/gPld6UBMd
TaAALNdUcSQwGIEyl9De7y8Sf9LGMFTg/RkldaDxSbQefIchhRv1OdV93sZuPGf9
M6WnZYFXmzifsGDfJlvOi7nOKiQROZrfm9QFko8QbQhIAAtEVVpA/nRSrE9YY1Oe
O9xSbtn936XbgkBuw7zni3ArPYXfKTy8Xp+xQDj+sXn3U65H+ihCpVyoxJ2GJm4U
zIe8mRLmzVjfEacyLflLm/fjlPIXSrd/7K94TZtzHyICdMTwFxeB/1R3+8+zRxsm
RlMaUAqRlnxOkkZcZXpVB4KhixdyHhPXpRrGD5qXaLzsVoHfdOc1syl0lr8jExZ3
zc7RBK6OgjqN1v6AoakPBP0lAfRQ8t3WrWK96OUwCruEewGOS1srP6HkSUPfls9i
rFnx+8g/isxLQj0uIB0OargCWnq7LH3sbA53g1stk4hbkQS7uacpsVO8JHjaBWCH
oDKEvfFTjFL1uklZuEIN0Rs0i03CgjYvNx+1pFzDHXmS15rnnDTI3mt2qEZHs0Zn
iJWx3u7/tvBOJ55DhDgMg9qleKwoK8JXIKlcoyGqVvZ1COKEgIhqu+h96XguzkRE
42+8nut23t0YlGf+OvpwSC8aGBeBGb9pz7Bblz/13S9J31R08XCffg0knXWXV0y1
Dty1lLQrAcpoazaMJ+Fa/V825vQnEZxO4yGk/4/WRC8bvGhToiH2LS2/2owoChSR
NS5CHiHZE4QHnWm/fP8W+6NJTNRsmYuNc87ze0pjSG0isKCJX6qzsFn7AJ0rj9zv
pw5O5lDPUK+jP78oICKSVp9z2hf5LXazWSEz/IenzftIGlHZDP3Ror4Na4iMmGaz
9aM0EGeqc12W7lAh7Y7HyWVJywwPWWjwHoW5t8FzCFe3x/weXK9ynCxnerC7G0+o
uA/Y8e5CrtTIAo/KQu/wZj6/LyTvT4sBFQpC8/d4cxZbFpoDNRH3mQAkVBlmuWTO
7LAR/P6s9stJD6aJR5punHD0rZjEXpCs5UJc6DkyDr731KB4bWuB/huBV1Jqa2+s
rTMaCWCuvyL1uh7V92HQL4U5R37cTrNSOL6JmRk/qTd/b8YzKpMVRYnrMaXdimwN
S1lAVJ2Y3+4Ox1LAiLS+j3NjwMteDbyracDDNRK5AzfZNQkmCDbc12jLZ9rNx/n9
Wmxcv5QXRXZ0PEtygAlhn7ri/rZNXVD/AmtiSIoT86npn67lLb1I5NeYv9ChbePw
+08UURteGwia0Xjwn/7Mtmlm6Q9LBHu1rr8Jk9zA/wt8y/e5JH/agxiHOAklWWFe
bSVWXgwKntpkUs/iy7W6EJlhcdC0JF4sg6vWdtu1zzSVRQ8lzZGs7lBaa2L5MezT
cFaBI8ZBRRuvGll5fzKtHlKurgk0iuFmekVh1Zh2DtNcouU6Tl3voH9CB7TXsB9/
eKfu0ojyD/3YMzdI5QMn6alPsbUZ54hKJQhwZxulMIgwRNEnMogWJhIKNoP0fk47
EKX1aYwyDqk1PaM2MH8V2MRUXUD9OTn9GjaQTt61ywNGM/IzXGW0JpEVb1OO+H8g
1Ds2nz/RR9GUJv6Fz9cpOJzQjxBbbNKjUflpi56E0edoCkXvHmjYYuZFi4a0K3wG
MwBWXJOZSVghQSq8WCru7rZm8ghfHZdv53RZ9TI8P73PhRoEOWsbWhon9485Crnw
VVScFjOBt+9eDcie7XIuGGZzi4WRYkOdRZ7JSImsEfiHfPFLBUmJfuFseEHPrbE0
a+xof1ECShjlRW/oabfB6AyUdQhdy9KRwkWDYhDx/3Vvc1S++EYUQcjZK+JCbVbI
ELNOgqkvPMVFJt36qI2o44FASlc0Su9Z6sUbr3Men86Cx9FNvNXbTbqJMFpbdrhm
qNsW2NW/lNdgM4tvbjXjH0JWIBnaQLBsXnznlLFB/O3OSfc3AakvfWQhnUQTgNhK
1i/Ho9FxwIDiyRpHa+gTjMseYWlRbKk2R5mhrTJuUrbQXdLM/CQcfNxNJVrXMPmU
6aF6NYQQ1zJ4RYY5u9T03mrm1okGLLC/GNqntQJtqVok+APbdxEYryqaaeJe2pU9
kgqtVw0FxKQfnrILZlQ08iagHRrwZhz1YfzzAky3xsWmDT1gmJVqaK3x/nzbPIAg
PsEN/7rG+87CWf8NOxz47Mh0XYmF1dWowABn6ZUH5cuJPLI4FUP2Jw1uRimqpqYv
N6TJ4/kV5rivu6Os9SwELRCLddm2dKCZgNOeFyyyBdyR7lpLxfjS2C42ao2i2D5B
Cpqs+7YBKcT+yozs6qdeREuW3uwKvxUHvo0kMylP+ATduEy5MsDPeDg1FprCJ2z7
XRxmlg32VrnuavS7ik9ofpFyxOBjqX9NIvzxO8MkXevOd4fBdraSq77RzFponl6l
yERf92Zo3JJxQWll6gpX8DpTJorxGdrn7zTIfhzOdWwhX4BI9yE7JYpKa8Y+D0VV
jt/pa8Jru7+4P5pXiRdl3zpBkwZ8njYo/CmEWTztQ5koviEhe+uqj419Ljt1EOdZ
iMVyDYhzqG0ZuidbO6cTxAvTyh7XzGhM/H316Ayvzynq3WmyATO/+yv27RZRi14p
TNbU+tEP1j4jrogiwe3VWLd7buFjez7DeT4X38W0RMfbZ3SDAIlUjnYUyEzC7dR7
ojNcU97y/rtLCabuWpcYmDSGtcyYp3uGScXPnqaVoo9gaiYgjHg2mWEddlx5CfDO
Y9c9/2761KhWUv/PyU5iYDlRqMoqz25q4r3NSGWbZOIqz2yYTGwh+cLJseAPCf0U
//fw5UVSTE8D1GXb+meFKZtVlUB4Vli80lntJxwTT4Cx3QYQP2QykheOZJJ77UVX
tj+BLor8+GT266NCyH/1ewMX6NN/Rs0Su4zIPhbbD/gHtbHF3E2rYiZpm28UfjlO
R+Gh9NOZ+mHH/o3jyI5U3A5+JCRMV7hNZIDUtd0Q/cx3d7Nqi4J0tCoQ8QIXgs8K
G0SkMwFpp7+HBormmPoedJOHK0ulN01W7s1OinrKzcrlLiGtAE4QW8Y62dZPmoG/
S+DB5YlN0tzBl2haLkjcuxTzPybCLFwpXkvfKT9JT9DsU/mkGJaRVpt9NcmC2XFI
/urLyfw3WbU2NRVToBI6NKul7KNENY7IR+wJFLQ618NV4hurQaB/c0u8a3iusuzD
PHGyVJO4K+JYJOt6Gd5RWqiGJgdWERzQqY3HbQx/6CW0cMuZuX19duebICDitq4E
/liM+g6x1uN62bc2nS5BrCueiKx5mc5gJ+LjSDW2krOlCiWEA93xHwawMd5vPDiQ
zXjlTxxmePEeyXiIDKrS790/rPm+omiw1AZsMkH8VsAMzAWHvFKhoIZWAdgoaXZV
C7dmVywJhAjFpLqGQmtBxF+ljXxEYICUrbvsNke/htjmAJDPy9j3b8CqugmyMS6q
grXHKZP6wiLan/TC1A8Z7Dns23Sb9rO4lOSygCIA9CC7Vxwn8clNyx/q0VRwGwan
1nfnIxp1u+kKqif8XSV/MrC5G1Dneqg0qNdPNEvU+ScFEFb3YhALCykrUwdkz5q4
lt0c68x/ph+an+0sYvv8dJX7MZS+fvGm3QC74jRgNwqTGwIa0qa9PiAqQRzT2NlK
rfxOhtWRhcDAgJeuYKDMAzmBcJrkTzS0NNxKUYMbjrRxaxCwd+qS3T7P2cH0XBLS
FZQw+n1LZjSwxjRsb3oxfL8R2SPULURC+Yp09ehgq2rWMRxXUN0v7/lWW1UTPej9
wyURlowzVzKMEnE8o2zAvd8JqX+iC8ORF2mAcWF/kOBsmps0n8H+FACbE3tYeLq5
PG1napwNEmGg1x0hugJtJ+wf/6mLtl7RaJpoGIvddYoyKtAPoM5Oi2DNG0Yx0Zzg
cgwwH5q/BDRtggOHAYxClGdPEcKoaczk/7rWro/aFEGeDTtyI6Rik/PH/ZGQ/VTS
JrkhBsGQxrnHr5uQFpVOX+HhzDKMPqkSBn6TSTM0+UeewMjh4iemSUrI5ofclm2j
9gnp4w/4B+aNuxLi8QNDi8A6yjOtVHKtuWl6OlQIxoRNpQ+r2Aq7uHDQZ6mdlc38
sylueia0vHQcaaStwKAz8wUpuYKZ83DhP4ZZO1vZUIRBIjCwPRD9yvaf8zwmUjNR
kwUOAb1OCndSEKFeEEN0CSJ42REQ1TqU+MLavTrKOlnXr3KcAZNnf+u7rqNOlrf2
ZzdfTVuHiHK5XujTXGfTrNyHVgiEjsacEe3mgcpEf59/i0VSeMdUJw4GXwLvxAB/
DijrCE765nA9mXlHqmuaYBSxXdnMabnT5yo5F+C1kbTlkSdwxfCzd6AZq/m5AdOd
YIorSzwagMx3AogF54AzTUf3VxUuJxSp6zBY1wPcryOQALJUVzsnPPEWj1SHAerg
1Ij+VLNEaz3soQ/rwGpYesZ4BCHxOvdeTmuZKRgG9sKcmy1ftnnK5O1Ko6Nx0ehK
BNv0/vhX8gcemLYN2/hs7cDBg4cu4868nGkbOGmEq1FV21ZWDjLCpNJo/qGT5hu6
EiXfUOCGaJfD94gHlVsaMpvi7TpTSHHoWqmsQ3gldyrBMbban5KUmi+rtKAg2Vd/
Fgqfc8A3OKpaLqFyR7rIAZvrXvW1/5fL+6BlyOXZn+NCjq6FFM6dKmuljTEXyuQV
YvvMmVlGalsOqxMwp3vAyFOoSiXlcXs7MxgQzSnFQ1Lfwgf9xxspE88jl6MA59nI
6Nq2eeuF0J+OcyaJhldjMPzyJQWYYqgSdbaJwumuaduKBtkmW1G7i+/ZsrAEE5UN
9pL/Mtwu6Jd8KleTVkUgb+R10dIhAYmjuEy1FpFFHVMz01Qm/irCpfIRQTYKJjcE
YDzpmagw7OYhQawikpIOwnsN2wbZMVy8riI1SMhzKbT6kvVHr86LUfOS6PEbxm09
l9HGH4Th37J7JTrtLU+GQxoNNSkMS+v5fdJ32XFQBd+e4oYeOV6pzw5C0vrGP/76
D7Q/856Tu+uQrgcSjyR80F7gk1ktRj1smDmnM5VxRo5Dra83PFMM06EjiHpmWQWx
SK/da3PmO1UI8P4HcXzpeQ3ERZiqEi99L8z5i3wXbudy7fK+3xHze0hBCWF3L7n6
uZizR3IsEzQ/KuBzsA5KDVLrsEEaAWj/eP2N+h7I0bx54DXn3FtZlFgPRzGXMPnF
kPn1xLvkBi4SyKQnLdeuJfcgSFdcLWFXPcfDJ1NkulfnVDgztq8xiKfXXQzj7mnt
DlWLLKBFg75XzdSam+p+ZyPNwobBLaSIAtrjsoQoMURfqsIIbRwbz8IFrmDVEAxN
+olzmedPbC/FAAIqZFD7DldTfY5KgQtsi7Lxc2zX9CdF2bDzAaCeADOULxmiwNAs
BMqGbbW/lYlgE5twAdu3FnCkLxm8o8O5NTTgnjaACVPz0ySQ35hv36d1LSDeEOry
31iVvgva20oMmKiSxCKh2aMNKPugnBjBULbfrDBEJA3AozEhhGS4MNi3TE3DpYFt
YPgn+amlAAGtR54XpH+6RucFYVORfsdTkkFrHV7v5iCknPDOioqOAW0wbUo/ARpe
r5m+/YlIBPBKtC0UhkDYRRmxqnNA9n8LFE8/REyucq7Mnv7aDIVQVrFiRq2c01XP
OdyywJSu1Dv1cTxwDWix5R6tdl5kwpt95yzA5AaqSdNBnc8Xs79u94UeKVxDvYna
SThF8kP52UiLK1/bALtYa6V6lWn6J7tsGUYokFZLPbl7TAmeqLVW4qUY91XlbBI1
ikAEFRTKflI5+oXwsyKy8+/4ZfX5ks/z8WJXr7Po3Ry0pX64s5BtuDK6LARay6gs
pIKuwP+X5xD23O3VYFUrYSEq9T40M+iYZaE+7u2EOfkgweNroZNGcBRV4/22OISS
3fEXsAU284YbQsVp5/0NafUgPUeOwKkVm8aYYva2LUMKfZvVFwj/qR2HJ0L5Lpin
TigVe6Nvf8IL7CrWV94XGTjxOfNvPo/U+pYVAY/xvpB9ZnATalhQmaLVvCYBDgkr
xXNIuckOWTuv3uT6rGcgvT4GZ0D1dC7k2xC5zD4AfbhqCNXsYRUkrdOkwCNsNOWu
xa0t76uwrZfJx/h0mBdSuZLq4OT6sAogZIvzjhLqqYA85SA+riebPLage+WPmQb/
4PZWsOMls5Oc0rcN/kd0v14QPDRFvuL57k34ug69/gz+R8Pc9imdtG2wDv/GY29Y
dJaZL8/wqx6CINkc6swJK8IKrleE7q7i7sCXjNDUE31ulpPTOoPV7XQ8gEMmEOwZ
F8Wg4Dw2XZ3JC3Gn/ZNlGM5MaAO8RQeDiujiq1MyIB1AZhacTATOlkqfjBXhSd/8
plIFlNFrtvERIdVV73NgoI9GM5e+oo0seaLXm79mmBnoVlnILU4HaG+xDxvoCqO5
wdVaTXKA8Un4wGtQqO9UGvP7xOZ0x8OK0DBD8GuluIEsEt+lTX9p3H9FFVKIkqoD
6YlsDriTcI9BTWrhYBbYbmBGPU9wWEVHErWa93++BomduQZXA+6tLHkWo/G/ZK+2
1Y6W1frIiz9qTFWGSCUfH/SF+Z6HNtvVO8NvVOQnWYHM46dGCHsX8MJQ5i3QeuyO
PYecOfE/3kPONB5e9ThPnSPKuLIEwOxR7Cin2qoRmf3312EJMaw7Wr/drcnKtjqL
RNaHXmwdFnIwPxsheIcv0xcnl+j1fsrfb5zC0Fxu9aN3FBRDS7O8JGtfg4YRN0Ay
65ZW9J3UMRnIVZCgq3LdpZjkFwwhnNdbJIPZDYvBq3wXHx97DSgox9RGHtbXh8YW
tz7t4lAmvYlGJ8I+VM57cZxWnAcmF71G745mV6hOlMzeMEpkXOd69HdNVAWuUS4R
oJJMxh+2Oy/ZbC1DKKG7cPPVBQx47mNLuYJNmoer8VqWyTtZwVUdyC90Ncmsa5Ps
o+5C6p2C5+3E34ERnfXt900O0FVw4zwBv5rUyfbZ4VqemoqzS8yVY0xWuCR0BlMG
j831hfJ107H3lyQsFv3do/8HUEGguSBuKyMmvqPY67N2WNPvxKMazGJXdu7JDiwY
zjR+dlVlSrK7azpVELUPwVh+q2rhbYf47A88waLkmZUP4KrqZbvhA7osr/IfwH8Y
A+tidIKEsxCtmXwPkA+Wh9AN9Z5gb33zZWNQVeebTG0ktrh+QinqOlDxzYV2xi6M
KTLQEn/b1Vggl9WEgOSmbUEfAhRlpImDUcpL4FuK8b7NPqZlc+tuLlkXDfihqw31
If+s5z7RjwePBwdKFg8eWRNsRoADqOsAI2AZLLnMG6wPHi1sNAlOtuJ7DGfdcJh1
+BIfjj1agCrQWwqSgSUM9UKdobtAGoDqsea+TnOZKnShsqLPFLW7COBg6EjQ2We7
7aWTzhBYSclNWb97Q1ZjfoPLfSrm1b5PPf2LgAwQiGgOiFjQ/3ok4DdCt9U2SXIL
HHzFdcletzTh6j10MrhZKlPyxtxMAk7PJW9+/2yxrGHKMBNz1WW3f3hg0Ua4KVaZ
57cMX3PqD0yDV7/8ZJLIxg04+wVxHaYRf1WjMobJkBKEG1QVsykumcsbdpUyp32D
o4+EdCgsWcCE6KBczfRQ8aCPem1k2tZ8C5b2B8KDp5bb8HvUnjZ85fla4hlvTjQj
CCsj77sF1w/F3MqzkGeT/6G1w9U9AYrbSaH559eLu2EmhsGk6YvAMupzznfJmusm
v8eKjllxi09mxVhMx6x/2n2NrGOmioyxRK6agVqlH+svjBI3nXYuPHxWk+800Bfv
Bg8Lt1Fs6FsaKV8CJhoxh3t/USJs/G8zvRWqywyZgqlXOdu/Zr234wiX4fAd2SOE
456vbMdKVqmbhPeFyKv2dKMpzLpclKDEj0BkvatO87OILSwZ0h54t0gVmmyuE27c
9h8JtI4AwUte/Pb/OxqReDycYvCt3yaXAgkU35hJ0sppv0/QDz3qp+MItxhBFq4+
jvz1+9e0LSEim0l0DYAbMyfKRgVpwrJ+AZuTxx+FCD9icMAvnmmXBQuzl2kdl/F3
ohuWcZxRmVjhybrYdd3pAhi0JAsrsf60aZ6QO+Xw3W6iDFf18z8p16Gr8WWIoClX
OPWHOgzIa/CmMRoal8O05ubyuEX3+UIq07Lhczhx5/KcZydpnNpvUN7AQHbghO3j
0t8ZbRmjRqK8jA3LheyWcGHPnt+AYGgk6CiFqhgYsZdXnnBJi/8xNdLTQROCSr+2
K4Lk+HH9SZXN7IGhNUDPiLPEQO40Yy+zoWXsgEJP4Fc19heXw0k2yD+J7CHRIGvQ
UJ+KVd6p6Lw6ZIpbSVa6p0jLXLbumSF1xJ3Zg/XsN7veQJXMF/4oZUROpaYqqsDM
o37uI9q6V4qkEjEux0kq0gae3NJ5r2lvW7KkCX1AC2h55VFL9oYJEf1EMnzs/m8c
LDiwwcRKZw8n4/YoY1VHSnJz+scCucJYnK2oSfqvJsBKMpYRW4qfV4oDOmpYGh0y
U5wtfcU57tNPrwv760cFDDl6fZT6t/RIqOcdUpEdJezoO98xKMu6gSL8WJUprbLv
i31UQyR8ozrDK9PsHvgBMdHdwOYtCi43nEhmcaPQjqAVIa2yVeNQLIyJuKdcJ0NO
hLR8w2LDIq65Va50s+U1h2ePUffsLsPJfccdTmflcknoKRHcUugM3x0VaETH6FU0
ARucZ1iLi8iRHM5VbNhjdk0GQzGB9U9pgoK4Bbqcml+HgYVGIU7GzP7qd6EnwHdL
UuLNJHwqsF3K3fAxIGgQr/XtQwA++zKPJX0Nse4C+R8YhPlGulsKIpu5jVAKfX1t
D9P9aAV+CtnE/KPp9PxZMbqwKS92w1no7Dv+BK12Cph9fIqVCB0wqO/nHOTP95uJ
64Unj8L8z39mOXAygTMeBPFtqWJ6NVcCRo0N+5/19EqDn7rK2P//JHxoJAnkcr2h
A5fKNN2b+ONNZBRJvRrT+6e1OjWZoq/uC7+PW0dtqwZjbr7sm4BAqi+s9OlkhOuw
Dx7mSnsVgaOyOxQdgzt7KSpU1Ep+efBILm4wClyO+oA/1Wq79/OWYEWuGQJHSF4J
VCM91LydcRHX6xaE64dduBvTuUEY2hHSdvx1t064INnPCSpJdhNgj208HGpW5LdA
Ch+h5dP01RKAD9F9L1gBLPLti0c49i+jSjZSv5xfi2lpKN1ZWKwHhd/GOghpm5xX
DdH3Vqyzw+KMrybelHWWTR9oChX4XtabD/c9si6EdmDvAGlcK9cO/hrfqn4MQvui
8Ee9dfghm8uosqj02sSVbMFVzzzFXVE9UQpF9TYzHU/9/WxZ8UYsOGY14jUWl4S2
CUhaJZYtSThpcEE4UAjpMMyWcjuWvKy9nRc4+vX3P9JpzXHGigY/T5HbXrd1SuTM
hcZPw/sovgYNpkO2Uv6AVe3JBuca9ZTgBGkDtdCW5ILPWSwuAqp3KKnqNwdI1sB0
OnGF0c7O+JNNAptMH9gMDL69T0hZw3NOZn/tSpODF5FgYCbyRyKP5Cl0TPetbkBo
Ri3dnxnCAlVDZO0lprDxDX0vXCEBfvyV/EESzKiQgwkd41trVMxutW88k+gvBlUz
LkvgJUbY2t/eUJplZfrKTFlPMaw8CbYl93whG+RVIfY7dEFPAEWIw2mjJ3JtFDWJ
YOUqrS9Q6C58+mi7a0M2X2IwU4PqqOKkz3QNQViDycHNlHtRsN47E5evrzQ3czO8
rwOf94d/Pa1tyscm8gPhw9CMpcFvU62NVy4JIHH2UpI6Tw7NW6sJ02vhW07VcWlG
qjQiswn3xXC1N7R2L0pnK0GZyDJaXuPT2dpbQaz5/gjLfGBiPymz8ERnk7tGHEzs
Gmj2l4eKHfkFX0t5zsgJIxOG36irCvBWOT6WbxpQylsPhFZ0FiZ6sWVZ3FkFqTjs
5Fq6GKZhNfDXdlk16q/U/kbjBsJbXcX8EDiQw2QmA4X+P/o2heYzysF1CdSzjQjd
3PJakjwOKtZnfb1xesSUCaXt+28jhWY25gVFlZBAMB9EAxzKrMokQniu2m1teq3K
rwuxKmEDCPel08yyJUnCuIDbE6h4LonderaOJj8YCWRnloKNsSTPmZN9eOTzzs1x
92g13YogvQw2h2XaZbLEQcGhPVk3NgWvxg61vnVNPqGODp2CMn2T/saMydD9SMnP
KDWS9vH09ROYmyuvSyFmIXVRuv1x/s3IwwmMkcqhhmu8QmzQvCJpQtIzX7j2e11F
p66CTRRK2vExaOaxDsH9Joe4MYyUxoI/gsxSMgOcI4x7DOuvWN2fVXjj3JidMR9h
fb6aoEGdmqxaBUVjTUzIq3XDhnpPiwGUSZCUlG/gCbqUqhMQ6oRY1ylJbMgCeJW3
DKJYDEKbtd/UNrE++5x5bd7k6LtCvdUaqrHJB+LfPnug7kXlbGHNk0wcYeDUDYi8
J1PgImqKfk0nvshm71T7DcAxp+9DnqwnS7nfT4JvKWVL7ckgbbAN7/iShCpXMsFL
6y281tw+TyBcdVIxnCBsjVPGgGiwy5sqXN+7vdHTyqV5DxsQc3C3Uh1rrFQETAHd
RFDmczQ2EEiHhE4ckgRY4HW5L6EKcJACjPwDihrqRA1nbjw4VyWks4HFtMWMr3V+
oGLWQ7N/nSz1cNPS5x5JjB1T/g5p4BsD2gO3glO+3gOiMaLERm16NZRdJiI9J4Dc
aV5dGGRUwtK0VJ2PHCGhkNmpsiJ1e0lIZRmVnZ9QvvBdBsbT4j8uChkUzBwGejta
Jz7g5rAI4crkJ97s/+6iQzkL1ERMLSpD+YU/zv+twNE1S3wndii4Z6tqLx9+eagb
n5hei1VGE17z6xr8YW65Tag1AzZMNRZFCaaBZ8dfpGQvQE5VtvRjSRqEqsYDnNEV
N1UEP38yEI+xn/h76WZEQPd0pheJPAMwzbcAU+mveIsETtfgzylNcLyFsUEkA+Mg
+fIMLgEfyEg/C03TZfVzI5LSVBX/fym4tEUrRcgKcbE4xfiSLPl22k/yHqourvnk
nqRzv5amqtEaNHYAr6SnPrLduS47sbLsyiTZz6qWb3xMyBcu9B2wNtrP6+4zTJOB
z5/MNDbbwb4dMXSQKI9IJaUXZ5AKHZkciBs/FGAASipr40JIVkla15rOoFUjMXzd
hnQ4DIyybksc9SkmiHXyvJmQ2yJkwwRQlDs+dkQw61kTsMzo7402pR0ndMS4qAlQ
6LIrQQqyg4E/eHgnE6JGT5605KrXcf3R23i7+Xx/JTWqKZ1W4yCKN4J0T5xQQvOz
CFz+aYfzPvYrU4gpXz3flsaUyfeRsAuAgFYWebw7P73SXDDny49w+3KXJDRfNgcJ
MlDSiR7znUfn5dOLjqNAubBCmoHRGBJ0tYXd55r4EKEGv6xnL27/pKBsbzPDMLTk
2CmEWppgHFWjy/d5EDtXeCo0JKVKX54CZak98j2IJG4DpXJdX+OmooWWFiB3eOnV
GxqBQzuadktFtVE7Qbkmd/x3/Lg/DXR6XAxTnV2WKbIXwkE5YYrxF/tkhEfRj+cV
FNyMkHtYRePhDlQevWDVz3jDb9ynCnY2p+FKyEYb7Ik960ghKgA6TQNau9kKsvhv
jmdp7jG2VywLLdFHpmXx+fumfh/MxgVG+P9jQzd15I3pRgoRWavsQ/5TJ0jDr6Is
fbU5zm7HS2Hhh6oNgp6CrvPjyoD3OIrL0MuWAvl+oiSdvLpSxrf1STBrakJcit5K
T3Y/fdwzvlwg2npvC+OIPSMgPdbjyHyAx7+Q3X7zpkXCb4Wn+mn21vxGnqBgprz4
idTiqqmn6eA89tQP1B1h6FqKUya3V1H0bxyuDyC5iMZ+1xISVYCG62R14xE+8Jg7
FClHonOj50CluXHFsq3UHX4N6gYQHKi8E3adXGBeApCKuw3FjvcXonIje3htI7Tf
ENh1srYDFQwek572uc0hQdlw80hNqvuok2DXRMuGHGvDkDoL9oKzFXLYPwnKAcuT
YbSsaA83yLrFpngQczlC5rCuLV++rRPILmJB1yu+ZnYTzAmADtn6K+YiHGcyaXFq
GbWLoRDfg/jExpv/JBFInjCPv1n33/8r8WRc+hEvDIqMbUOJSdhqKmauTSrYh2v7
zPjGeAHxZA/xLCShx/0IclEuOg4bxx4XXK2dsBM88OLgS98fiwsx1WdXenJJAFOF
51Bs3KQyNwlQ/h6cWFeeV3Z6YZmpm3zw9vF5qv+uJomjYroBohrhAFVwMJu6VpwX
4xy7T32wnMAi3Adp6f5YCdGR/oZQXZgJnQ1/JLVf2sL82eo49rpOghsUIrVMrRUu
F/ksBimiWTXfBiaXF2hdz6+F8xiGY4jiLKM0GkAObXabtv8p5BPK8EZSwMNZs65L
tgb/+mY8k//KSxA4fU88R1cwwbPHMvnGrUXP1f5YPxfTeOUI1vp2+kNUJc4SypFA
KDE3hO25+gLr4UScFnNqPTDUaaEFlHJxzT8FglDFnlCdLMUBWH61w5myUa+NEr4p
lgFjLoMXmlujdXgHPfod1nQqARRimnOxPzLOt8AaJKwMvMbTtYnC/+E8AJGaq1yu
p6Sj1AYbYC3+QNxffr0MdenBTGET2DpMz4fshjiJ+dYonFl7sEXfdodOP7sIF4Jz
RzlNkjMBmz9lidMKhGzMpI6Q/Yv76Bf64oTUh1JOgmFvJLvedPVCP1UVQPPkYwDA
869OuErqoFEr6Y7ga4PViRvEJnm5d0LCGECU1tIvAtGBRA8qeH/scKLY1TVMWFRs
W6NiakzzcWCC4/esvc28HAHfILYIh04xQs07iQUTPJQ8J6NWYVNOZ3ULBJgSn5ru
sVsDvLbv5YgmIMWtyP9LpITANSXJgXvXwStBAa9sWFmi/zhfDrOjAIUmJT18SBBJ
BYPU0rHBbnx51bXzM4SL9UEhvMmZNjIDRWTmxZ6w1kexZ+8EaNv7ZOCX8lSK80pR
xxCn6Ke5KyKZxrtYApX+uJ2+RK2/JHbTcDDTRCzhI8vOykALgtoZi6ODMAj0IMSV
bbrj4fJ844+xjAv2bhl/1hFHv4hKOciw4ILcl/oo1BRggqJ7pjaI8zl/rSmS+34s
d881FqleV6qraebcrZg1dyA2XQ3PK3Oy1s3TYnEqWUC3LEscis5OaFHohEJsaa4k
t5nzv7RfZ4mtOg+67MnZ7opSepLIREQZaZBxVgDjgoh0i+5CaBMf9vP+xH9pG+JW
D1ITuXSgul29VZmXutBwU+dGZ1j0D9EWMY2DnK/NyfIlW8hYfol4m4ko638Tpfs4
MkqfOukkuSdfSubjBs/D799npMyiia66Ho8KA96FnuPweLDnEX4K9Mh5i5YWZBcc
4yyijPKi8evv21JWdS8G5J9HQv+LhRk1fmLZgQ/ywITTtn1OqrhNxmSSkPtw+p8z
/kRZMra8/6m3MthR+w76eWT6dGzL/CWOfneJLYWb+dD0nCodwMTVhtoS/j1hmPqn
mJlaGKfrm49AyWnouV5BN90PkTF2awrOEpZvgAoCN4AO6Z8BRlsAi8OgL4zr9S2Y
UB7AUkZuZP5+XCbpiijhVPRkc3iXEHi4kZ+ieBrfH4ODnPEObBt7i1WzM622L/OA
Hm/Op4kpgdvlHatfmR7/cL1EPh03f+3Lf+Tt3h5GAllqM4NJgonIcy+DhoeYjQ+g
ulyDq0JcNOooHEp0IP7sp2sk9md1gyC+KRL3i68IiZKD2DIdbiwJKR/s46YVNjOT
KpYNdwLATpyyFpbBW0M0SWmvVXswYl8yrv4niBCiVDFGBifPBz0HPaQZr0GP8+ds
XtM80Kv08wki1HSKpLyn6uAhls2C/aOJgof7Y8UIU4bVx2ST8ImkeCLOk094R+Sv
e4KrNuQGzjbgfUskUTpKDBD3atH2VPkmQqeJmr6ULxgFIvJeBpnU+Iw9mz3WKlpP
enq1X6o/3+rJjUaG3q9HGDmFOvBXA2yfuzQtu0qg2xtbunSky4QGx4B8C8WnzyOw
tPOVFspIvOHwSZIrZ9p6sFeerF5+MUUjHomaAsCSVKulfzd8fGeMdr71BJHffAAl
arLSUfeU0t/UKpmzVojE4HYIInSaugMt1zztlST6UpswEHqhfYxxO1X9ejjIIIMX
nzst7KhS+qxJiUYBTEEtpLkhH6819Xkzs1HL8hOnLMtcy7N7bybg99MWzEqcs2UJ
zAjJP4kYBQxwFJfXjpnw4oU8VC1JFwuWdill0M08s3Xk2am+oYRgirFo9zbAmjRD
3SBz0mMjeDeosis2JOiq0MoEdDafNydbUoAJ3CYYvstWhJeTnKoXO/YXN1Uecyql
KtmgtByXvhnbugLRatbiJzbxwFWBrq4/uMNBL9xmtYtmSh5FI8/Fnk/fxXB/Of1z
WoGj9DkinVI853u76JIOjtKosaM7XfewCLAEgP2UMZwpj/Ju96qNpaALYMy1iTEz
E8WHosPeplYh0vejYWW02AC/Qo5oT+9eRreE8N0Eqw0yfsPaua9LZS0VGAkQnkVA
h3C2gc9fWoVH5zWj0lKxzPWr8Sdy9Pm9PvIJ6ljoST6Af0yZ7TJm7UpGxsXdXcqG
18wl+AojBs+ZfqHKcc5kmcnGidzWPX9MYUtNHT3ko8klk/wrqriq+49bjNMgumrq
F92KncIqkvvqRXhQ41UPeA+wisGEfx6VBAT++EdW619myoryM2+2rSe2F554+pKs
cFnU561mNiufApNpExLwgPeoLDWMsLkolqcXTTgGO0kCMuHXcQywiwdagE1AXEpi
H7lbL0fRD1s4zRrh/YnYgy0EbhEG6au2t7FBA6IQH3QumLfs4EB6tE6UjM5IeXjk
2xCH02r2MrOPFaT3zyFoFLJZJRe2BrabXjPrescloP8IhPG5us2WA7x+DDc4kaUd
WUTAorRF5aIHjJNgCC6Jgzc3M7qKMi8dylT/yGjVBxDd50MOjZjOPQGSPfrRS4k3
84vQkySjefAo2OGsrXVoYXYg7yb9YCH8XZB7OSeSP7t8Pe6xwXp6W4jgp7CfMFYZ
cf37xRQsl8xnfJ89JrdMEscHjX8MFs+MGs6mbRbW6/dOiDARDNzuF5bfyiJzy9dR
2Cw7DtHBttoC8e1LJLD/i28EjpW8PWFdAYOsEPC5fvR9D+sVwX1+O9wei/+7g4P3
lVmwXIYVU27nCbgIhmHPlSBet9PNoKlLiK1O5IJnKtYA5mItcKP/UAGLQ5elZPrl
d8bezvl19iweSnvGfpq0Nb+TSz1DKbPoiQ7rbhlhGVb4HaBUxXCgxgXirn2oNrPs
fkJ5A2RYfUc+7zcAixvmrUZ52jaRPBXukJXXBReM6+c7idI+muA7xxiYzaY/UjXD
Uf2/LYKpVO2pQZP8eHN+QONxeZvYUVguvj3HBN9kcHx0qkFnKhulhYsP20GeHIAO
LwKHKNLpvXZz+QTu4c4ZPnFQDe0f1pZkZpFSWcPsarqFdlwPNRTZ17l80cCWq9cd
JVwafykWlIQ53On3+ZwghjdntJ6Rp7wHlpEYRXDwodCiDgaV3g7L8gbxOHEY4nWx
x2t/ER89n7W43CTOggv25R9Ord4d2e/F/r5DDqWu2jPh2O8nz6OeYobIWVp2mSr4
MP6JA3qj94IDjswdFp1c7ZPTuVqm0o+J6WnuOzdbnv8EnKIbxIWCXHM++ZNh3dYs
ex6YGRvyaM1U3ZHSIXR0mUV0pqTPyJOou1Rpp0smGOHM/AcNf7yVbc8cXbjV5d/5
KnhOWubCWeeCSe74N0MMQshDqfYLzXoaJsFz+1RbOtCv4j+l57pK2ThOp0U0gZKZ
ZaxexO68ZzW5StK/sAuOUBR6UyXI8lxHd5/6QOrgUre1/ZcSA2d/UWq7F7v1aOpQ
I++zVvv7R/3gsj9L5m0iNPEgR4YhbEbYCJ/LFEBVUNoADcOf82J9InL3ho7jgoD4
BFbuOFfju9EO6Uo2WdpowOnhw9oyNMWz50HcPJpSYd/yUuPNa3QR7NKyqH1Ppm8i
w7BOT5XrRAVHE1983MUdtXjBfzGocdfw3eacjc+9jitPOsyyyQ18k5smB5Vr4Eiv
uQ14JebGjDdrEhGm4moGEPAtDLOJ3XlDDE5kj4fnsJ8ob8XrNAyKDBQDsnjDRjnR
WwABOGmmGrU5wY8h/7YAfL6jpR4NS4nLUT8GyUhSEbdxaqjJ9y9166xtvUiNq1Zc
1bB0PGQEh4P5QdV4FGnymPlPPevJIWLAB6KWNB0xWOiZMFQaoiGMwT07fTNOXziL
LQ7bwsN0tLqwI2IjGoclbOKBLKIh3C0FC2zU92YdOY7bcyzdeHr/l3TwB4DefnN7
6N/qlDBWhw8or/xPeP08G4jb6WBuWOSfdSShfYOaNFcAh6S82W+8TDBjS8QNQgrG
iBC5b9zUHjSFfZAvsNv/xQrTQbDkGBGB/A04UcqaqFQydKqYADimNMYjnpHfyRkZ
wW6ObCp38tpL7T69jvsvMnP+wym9VjvbTY88j2x9/jO44FvyA0JwYWPl6HmL1z2M
U9EVR3NmaEPz0V+R/7tzj7XDF+1XBOCuYyq6E848Dg0WhTYxgsycCA/XsS4JZlrv
+VqnJ/bSSJqoZz/CAizHhbUoH6Ack7Hck3Uh3Q8bOOWd7wpGY29WekiO9aenCLbO
MLC70RTaS7pWocWaedsLYwn1Zh8YqRIxusYWCTk3TtoPq6cTNs4j/a6Bl6N8VtyD
J3x2pH3HgLvs61sJB3noneeYzCAYO3fyHcOYd0mWZQnyOB8TzyENbdIU/oPAhPq9
/OvB7pHtnzW8PvN6/LBOxA+Kv3asYbjoKu9+ZydvBNl16j63niI0JAbx02i160jB
QjcmJ0e3v5pWB+7niER9b8XpffKMXr/PHnlWQnHm4+P9W7/FksB7TT8v/j05s2DN
4eJDyvGGqUXylvuAOu/6Ur6tBjcnG/1q+ol/e7OX8V260xn28fAPxbKbMTqmokwt
TmJzTzNnBSvCUpPAapO62Uuf3Ha54sDe1/2TeClHzXNwhFlNg0QvAm88GZKb7kYW
fg5zvbfI7PLwXktxTTZd2xOYdBxrAa7Qor44Ck6me+HdUPx7uxBztZ3s87/frlAe
MEEV7UytvTaIMWXICco/2OYM3gX6ktmq02ojeJgaxvKIXmEML07y85FH51z7fdYo
MDnstE7V54e7tq30exkvhpRcd96q5yF2U7p4nzneespIGxAYPeCH770q2WPttegf
c3SZdXI0/iQAjHomki5yIp9hMSaMD6PbdLceSEk3FJBZkXBIkYnetXXWSK0jkWBD
AG1Cw5DDJs2mJ9R1pb1KyebN88vxKIM80bs0kPNsRI8alo+/OUKzEdRjWiM2WbTq
PX3xtREF8VcoeEMi78gh1FZFMmvVNXFntYWfGxvwPp/5jLcR3YUa0HU40BVx9BDU
xCNmC3ENzShjSvkRC1myn9P+2khInoRrd8vkRCeUXvaZCK2tVK9SBKAoFoqjBo+5
ZeGyzlIc58jtE8L9J6RQ7R398vdAVIEU2zxssCPNTU9s0NWLjKP6BsyHZMxMVNyv
6zUL0HhGhmLL68MU71F0WPjftKj6z/DAwQ2JPrggaeqUaMhVT52ce/Lsp3/181Zf
GUvdGszJeeHFyd2C2G0acKiSKPcaiT6qHA22SwEVVJgwgaVHnLOORPpkN5loNEKJ
ecE6wN9XcIQ22KuP7Zf55E8lvtOtb3ccq1EX29sEhDTe65akVnTOy1il0On5BHza
eZxnVRO7F0bqnl1vavi9OrEM+aASBGpMCDJiAm0iW63yFA1+MeFmPpcEiwGp6Ln4
vVkvHgm7ZtYlJ5h62sLx2wpfkdHi0JO4WZWARuXjIKIFmYvhcZhZC4BZOCTn9VaK
QQ3cj/pyxkuTMblitUAs+QATg4cHqd/d7rFLx3fX+vUcRWzKc8gjlLmYItsdFCA7
P9cefcaccD62Wuq5+1a1HeD//nmdvABuvWrcDiUHYoQBZhoPxywxR/4cfythq2zx
KcZiC7IL84yKXZTf+0HBF/WUym8dgc7bPyetfz/K3r6wttULe/H156skqQdfvsC/
/zPkQp1x6F//2kRrmg3roOnPwRPjT1VyPPc+4nkc/d+ExUTbMm3f/CQAdmPzES/7
hIIGMw7WWdiFyMgRWKmbRehle+tdwEFHF2qncZksDnMwUiF35lSZwM/V+FackFGK
cXuhg4FF9QavrHZ400gGo6OHtvhj0ioF0zM2EFf6Uga7pULLF/SllOMeWesSHAtq
cdYUO4LentWdNEZLkkVe8sWCiD+zYLl/cMnH6bTYSptW3nzrV9x9t6zwk43JeWl2
UUxG5SCMEQ9lcaNlOsZcWvseEFHPXocPn77Ekq8uEaDjRT7w7pHFmc+uMRdT72xf
1CNuAR1RG2CehVZOouvFa0s3+n5pkFuuXtLAWSGynvjyqi7pGB1/zEBDMQWxHaUH
hQ//3Hq19EJEHbHnYes7fWCeVeLn7XfDuTJiUmn2uuQwakFQjxZZwrFYmME3z9Pn
yD1UwHCFm0KBA0zGMiuPWMQE0B6KcPwmYinuamOAMwrAM9c7h7zKmYIMUtsQQ8Xi
JPSOoJgWty/MowS1iGpATm/J7Xqdw+nJMy7inHanpeXeeaTGX71ZR4/I9JbFvgCm
cornE/LWbdupweFaXdMYMzuKJtaTcHymrTTZ94cXgZ6Wfpd2Ijr0EBb92V3rZuPx
1rm0qmCHGSpSd420wAWN29fA+XhxBbkMadhgYNT8Vqj0ipa5V9L3AtCb/o+NWCfv
LXovDw+8eNoSoWe7CnIM27p/jlUtkduknoKuZFzN2/AnORtnTUH7rrglWhIRwJJ5
ySsOSHEawYTpv5mzoyWPnLjU9PgQfmOneuAooBF/DdigeWY6HETOsfT9D7TC6OTW
CoupUIt26AnXBZgMQwZtsrqkMjB2UIC9CaOQIkZB5Ai+uGQzsSlQHsqZCf4fuUeb
EvlO3QCvqAJXlGD2sdiO4/3aEfkcBns7JSl1IQbazLDLYBIwhGleTagOuQKLTRkU
6fTdSO7wEot7Z6By0nNfdA1k1omBbazAhnNmCt9cOAJP4NqVZ3Tx4CXy44dvbjyG
pPz6HCQ1fgkpfZzyGJ5LrxfFUh1an5UAYfDUTqHH1cIE4oUodia1hLFazURufEFH
UO7N0RGYIeZRWWvK/rz4FV2r5hXDh+DyDVO3jkZQ3eVwgYqEuIu+Hl04ZJFRBGfy
UE+u8iixwawUysX1IoF7/c3vVUF7chCtUHh5DXCRPB7B5zn24rEjy0nQWKJH9t1x
kSKZzSViv+wa5TzkpJs1vCfbir+aq3cAz8VLIbdotKsaQso+y7lo8eJhsiBfxC2+
0ihQyKYoUyjY7cPsxG3I/fbLIh9/9X0hXeG6wWxzHgRyixFaljMhQgqxIudeqFv2
6GkS14rlHbbjsT0zOd7C68I7QdENMmNka9hp+134eu9bSN9jPoCxwXk94rETXEc0
4hroxNpIXqpPedNegtGhPad799xmuw7laNT8aEuE+6txfJOskFK/WOsjmepTOe6q
W8xYe8bjVkjmwk/DZngZMCFsk+S4JE8X7IVkvUlck+6bJDLjaSNTKcO8umWZLA/x
xfFcOJ0rwVcJFI94zQFoSRNrGtxyTENskkzdvxFuqNm8ciWcSILlFqO+97fFJ67/
EWH6wcyYHj8Q0OD4KGtkEdUY+yEOcWxQY3nOSzIhvo5zgoldQsBiGG/3idbbFvu0
VX333dx0BIzaLnD5lNKuoqdDyPuyR3VmWAPncYdOtG8Ni4o2bIq5YjV9FRG8D9El
JCGeNEfbTs/nio5+shaaxPMbnjinfpGd+21ETZ82VxaHIBfLoGPnkiZLL9k9na8L
5V8cqTUD/3Rh+bXatsm4Vu92A0RZEjGy8g+9R23cInGS2wjCulK0tvv/2QF8uLXK
sqwUSl/rrbNFudq+Yx8R8W91Qo0MNVv6CkkA5HTRrVodnDAhHXGHIlVfG+4NKQZH
eHHfNHwas6KqO/pJx9FwOK9p4+/YkxKG0TCLvuAOrqwnN8q7/ZAShacP7VO4fpSz
IsiUzxHrCEG5rSjgHCErJV7wQF314StCXpASE7okf4cJMP19rMLRmLA4/Honybsf
hmSdBNPx4P4P5d8Vmz13Q/xYNh/7JiRym3xwe+tYN0D2UQZ1LNxxfAGMIaRfLwSZ
vmZWW1fjiK7XBM9vIX/MhFPC4d+hKkIRW80Q03TMMwDxU+6ZhseFeJlFLAyCmRvV
uc5OW9eHWe2cjgVQ7VM4N3rrD01JOsCrzdJc2UgCU0YxiOyg+sc0w7/nIo9r42G5
0KPMS5qTO68+ZAa0RmBl/qkuwHBw3I+E/+LpHklHks6q4d8TcH88P9zkGS91YWJS
Sqcs4qibeNpxvSUF/grF2d41cmr7vtmker+jNvC/xd+xQx9ofznb3fmAslA0V5Hp
0pgoezyyTWEoSzQbtUF3vEE+GXv2rd+5tqzNNLkhroIh9zuPNeCj2gjGkWQkIyuC
1IENkoEr7D997hmYZs6a6WZ3J8Py4f8lUG+c61OvsR1USF8ac0Jmt4WNtKvvWTcD
Vi50+76z0uHjNlqLDiRh/+X33UalOIkkk42VqJiRHXoqlNb2ULbIyHLwomvNbDlq
mOHX5LCvkr+73k7FjtgmjMyz7McNb/lYI0Ma46I/sZBfOXhTORpwKjLI1BPVPy/s
cKIXXWCpK0RE2fXikH5/p+XxnNGCPkqq9ZZB7sb6HxUB5ZR6L32J0ZUiN81OSQST
wyOrsop1V+ITJX4vmyXkiVF0njZ6KSJfxD43dyPgeNt888JoS82gY+i4gvlhs0GD
IJ3nFiP8Q0M9nLDovwRn8keoI1pHYI78sjHVOw+rMYXumpekxlXPd9xtWdorjNNI
ZVxI4xV8y+2EgdWSfrzwBzficphiSJA1fj+d/TWkgjDzHLlSJzxAqU3m2PRFX/+c
/2D2Gw+iAhzP7VC/Frw7aP6Sb/XYI3y0S7OVoKQyWItffmk2vfYvjg5DQnZ3OCwM
xr3zKOrzLgp3qD6yJXzIIlo5cnz1+4/XvT5ZfO+ua5CMmn9n3VQCCzqSOvgnDUQq
E5oMPpz9rxd42F7QDKFhleyAfaCvEwjNw/+LxqctU6sfBRLQQ09MPyNiSyZqNXHt
qYHQVq2+WMDFkDxRcFHP5BfY1ZITcyQkcnp3v1Gjg/+0woEBfaI+FoqBvHX/lcli
eujMHhYzX0Br6hCDL1ft6QiBkLDFgIcFKm8LN2cnV1LewI329sLzuk+FW4igDQPk
HPRTTKnBWYEs5yvk/t0k1BH7E+RSLNU3bTONEpbYrem0r6mna40iqtrP0FwZGULV
/1pM8xWE/Mdvznj/+zhU7ku2UJqdhzYoFdFVgLNHwrgTfNe/eEvuXVzOiDeVrTVS
gY/++Km7RGHQHiWWYQtBSQinml6xZ+pJnIhXpwzEjnEVDC8gelZpdwHqtXJa0AkC
27ckU4yQ2u+Tjg0r8KVWcig6XnJRDSn4bIWYmZmFwnxcLD0DhTx059YqwabLSYDl
RBzgYgMdBRYI9dcqlIp7VddkQyymEn6xn+KYngwfioFQgMY9Ql5TfO+0x+Hu7hBv
ocHkD15Kz8nkWHX251MFooSIJCvIeRrBroTxC9phXr7+my5jceUu+pbXViHZv4YM
c4erOCaiJiqdrHkK3mg+rpCNkqr6xzaXmgFGshET0p1Qtw2J7TqNPut7FjABe3U+
hpoQ3iZwsZhFNzz6bKycNbaoCNkpa55hIPi9xi4wgJUJr7Fzfi53tsQvhtjNc1mq
0v3cDcrVlltsjmb692VRwvfFhGcxFYMMb6ixXMXp/S6cLlzxvsxYNe63AT320dSF
hxJSenVAYvG7IvxfAbtuVNLIMAaxOWclz5ziWHaku50oxtbdvdl4O4qnt08n+/M2
NVKga55TL2SV9HXtjFGVQJnOglXipGBjSITgl3zpzGm+c+bivtPHVh8Z5A4rEUHa
oSzMa2Hw3e96c5jUizaeOAAKZfVsCv3nzdt+xz3lAbKDDrS1r4yDNRLw3YgVpB+e
Fy+8IKQ6oXg0pSwaMunGvx6oU/FhQRYbptNqEgJSLRPgzirK1Y+kr67YmBcdAI2T
UBn349wCC+E49MKzxDUH26rS7f2MpN34hF0Gng/rU1XAquP0cPmSu1KZRdbZAwA7
zyZPO4f7GeRGtBx991UK0gW7gHzidMzoU9VyPtVQRvXl0GWxQlDl0TzvMVtmYGo1
HrAhDNnSsaV4h8yrYnbouegaW10mmiBLwG0ifLFubAIFn0JuPetGl00fXP6RN2wM
KQMn14rh17S7zTjMCyQUVOkMPbT38r4hnN6c1hz4oXYDf+ZGPJFZXAT3y9kJVS98
rHvFdFZBdD52bThnk2wGdyzdZZp2gU68umyN2k/rwzSnJuVUFfDijyFioAOj0Spr
BOf8tO5N5uDoTozFTISBpO563GtVDKTAr9VuoVBKD0G++ggT7O1um5DAYJulGm93
XHHchqgUJuguZbfXhL4Yq+ba/VPYhuMkzOCD7Zx/SFNOdulOf0uIQ8s6O5K+wJUQ
9mSFzaHQMiemc9n9BKt9RxUiW8xowCK/uEQ/LGcRqkO/jiifyqgPTkWMK9yHuRHI
qDEZd3U0+T06sK82/24lk4tSSf49vfuLZ+tyLfaSWiMkPI27o5m/Btv4fbrCHbEe
DOzZ3xS7UvP26jknPZR2FbSqw3Bif6R01Yrpsh10Kre3/Nod7mWHVr+8JqJm08Xt
bz5kNsvesZZtThIgtfEj4CLgTpWHqxbBHmYYdY2QM4UlCLCl3ziy5DlJNFvp+Vjz
ykpQzYJ1Nsb+2FLwbukak1VXhBPiEglyXTLQW92Exd78unJBd+10N5uJx+P37rxj
z/B5wuTwYrMSBGQXtL65gqwrPRo2oR9ZBZfXtdExl40vRY9wPFjZqp55nNQXBVmi
1iR+L9i1dyX53j0v3acrbwDddF+/1Af/NQ+Sxvw0iV4cGwvI6smV5o29k8uT+h9g
1x4/oUi7RMfVFKUUnisE/1+OlucTvsRKF/VN6depevtwHSeDKqGTy2JCQQjS/Q3l
B/mc1pnrfRz8PIHO9RJxINGy73BI7RQvVGwBhenKFz4WLXg5PCXeG/FgvV+RBsZp
YnRvrwUCgsGF8musqQREF4DGURKO7pB3+5bXxBUS0/Rf5W1msy11IZn6hVsEEHgh
sU00aeGJ+hsDpNcQTnB/qtMvq2anfW0coEH1/GCS4JWCxi41a9azBK/0uYRDdJnR
xRGPUM0VA/uJuklljlj4mqmKhJIU25RbaV/FllCO38DxZPrHZ5Hn3voJlUIpJnUW
3JC9bQzsqdv6To4O8L6fJ60JZY8JPbnYNsOELll9yHlNoqaf5aZCvtOLaM56vvai
fmtGeBZq/YFKT8NailZ9F5ip967e3TnxYiJ7AOok9bUmtDY8C2CEQDdw2IFKM3J1
K8Q3PQ5q52EJZRH/YKJW6nDln+j7TE+iD7foWSSNPFBIdeqN1eqysOVRJDZNFWlj
1xFYGHuZaZ5xy5S5ToMbKl+07jAcmOJxf0+xV5AHZURlEE1g8gQYLuVDyyv3YWIE
V3dfsAPHz0w7IwwvsZxNO0If2EO1eUbkzINrhhn+zBP5tXtg/xj4cjx7piXw8Oxi
gy/bjpoVE03SoLC9BAAhwYp3/NpB7nGuqUxiwUjdE71dgfhwgKTGAuewutqEwQL/
L6M3PtQnEVDrILseUyawFzva9//wAnZQAKVC97MnHb9DRlF3qEHw77+ZjkA7Bs4D
U6eIXEt0GO6P6cz8RonkcMnn8m7Bz4zOHgqpapqw+u/6Iv9Uy3rJPZjeMdTGQ1R8
bX3IJ57SOikMXQH0UWPGS7zfjbE9htuHsxUc7iUsZZFLhzpI81PiI9ZrkSIuCNy3
ylhzQNruOoLFhyB+c3UePQ5TPt3na+GUx4iXk3eLCzwl8kMgMUz3caCE8uwWNnGE
nktIiOZldKof3KzzEJD+osRPkqciQs0dhbr1jdgs/ISLtnAa71a38/LDpTPUGfn7
kiscMKECOdbKRpY6dEivscjmdkk509Nq0A4nBzG9aHzf0OV5y4cfGLmD7vLimi9e
a9Zuik7VYqpwY5FsTmM56xFy6R72bcarjC1dZD1lUrkJaE2pud2vcsLxdcLLGpy8
kPI0ZDjmbFCnK1G8H+PiFFyKE460A5lsyYhRi7BdjQJIHVkvo2PbgXFuRdopRmE0
jG4t+XmKw180kHZR9PPDGsVgb2hMpErzNUiEEOKtwgqaACt6qbArzg9PnECWLc2D
4aDhYPrW6Po2YIp6oA00I5cghu7vJYV0Q/Z0eB1w5oPfJVRxzmKPYKHS0kHEnzd/
pfAHW/9WRa+0D0LyaBLEwFr5NGgV4Kr5sSiV+txeWDYjQTCaEtPFYi5q7qJVVNOM
XtUnNsioWmJKCD0mkDKavEp8gt6ilUpRiTXeqUE6HwlwhukyRoHgPi9fKyL30j3G
Pd+94RM7stq1o+ttd+No8eU20j32Jn0IyyY2FiD2r6oNZ3SEa8HtjV88opRDL9hp
fvcHKqXgGod/DWC7ljXuKhxEG7f5p7SGsB4TVNJY9lnWWRBiXmxQBfgmg7F5J6UU
BCKL9OH0IlF2c2FRPFclDuNaJuPcI1ue47cqb0RZR+vv2B2T+cYIc8mQ2mXyrnqy
DWl9EWlo5u3vMUDK04FJwne2fRnY+15JxQF/WhmhS2ldXFhrkdyZLFE7OXsvvfL8
GGXtxbCLUaLeRjI8VAAZyAMwVGrw05BrsbjD900SSNz16kCayhHXJ5N7YK21ee+O
pkzbS9cp4H0o7vnvgCyVhQgajA0s59TAsLntzu2pBAWBmF+0noLJHDJiCkDhjtsu
WhXxtPR2Cq+wl9EpRSx/d/vmSYXMAifyWVadpekg3h/04u/MIVIOdmUeNgAVRypS
5shN/uNawSC1neUa6Y0YQBvCDWQ6wKeZU/2Os4PDLfKjjNOtQ66MBX/KYg/38LLG
KCEN2ZDuV0YNcURyO22tZJOLvixOq4tRhumfEfax0Uxp6WgTIrmNLVbR2cQJAnZA
hsjDSazHUb+ORj4zILtpKGcBICCesTR4vFDS4fR64A0ZDZ08MWBk2YZNgS/KhsbI
sEzlj/Gu/8m0fmUQEMvx5ANwPah3rH4bwYUEabqGiiNw0EvV4YqC5n07JfgsaK6E
eXFKlArtZfCaRSTtVoMVqCLlAHMHXbzTg1/3Q7a6L+5eLzv4PqDAB9lEu/FP221j
aEVK59e3DZbV8MHXQ2Y49N4ZDPf9iBDuKg1GRJ3bDn/R8xzj/BvlBI0RjWOn53W+
6vrt43/Xt0DX5oM63uKGyyYPJb810Cc5oampSGif8Qyi3bNtBVf/DXCGuRzDsWvi
ahWkGTnEcB5qQqKyUB44+co7IQn0fBZu6d3JTEhkjMdmTiRuRnhpOUP6LNlm3DWu
7VIp+Ntwf9vDzIe0qQEQvZTUucf2Zg7PEDgnYV1JyzRSpQ8tqsy1rEJ75M5tgASd
VThPzVJrm0ONF5n2WXdqFqPUnIjqG63WIJRUh2hmmo8Attkx/E0kKecnsi3WYRa0
Y8YEcS03ZnihFSz0atjRRbK+uUYIt0tBD8gTJD1AY+3FCpleQLmIOkQsMiCBl+Tu
+VE/nHFzFNkFNxywhCKD5qZPjachEUDw0sponxjjNle8yprdqAxgeA3OIS1ljDl9
7/Z8IUYdWXZim1HtloEM97zETg9d0ENiy/ND1FfxNiZqohZbShIQ72UPS1KsPoYc
SR7pv5Q47+PHsZQMuBJv7DZdbOzEtuKiPf48SVghPPF3EBHJeMja08RJovsXFoKL
SxkcOxYJ2ssZ2PTjoB52r/kqkBzMJ/llpO0d2US1wzWs1ldRVm9zWIsb4u6yw4O1
cMEhMxQS6BeudhsmMBcdAdnFPp7f56mk50X62zzd+nyZjWJ++j7r7PnnUcgZ7LGe
0YCdtPLyZT3AZ/SvxfYOhbmqzBANM2AlwS+osfJNMxdUVUg8LZogGPuis9rHAzeo
JTcEmU+1nqtCXSstHsDs97nPhbimJwY0Mxqf7EhVUSaEedYO9UwrJeSzvldXeTrE
XuB3ChI3g2w502q0Q038aVKvv5J38xZHCgvt1sW1TAZZeZ3NG30rLaO+ey3I+gT6
TL6viR0/uZIkHMnhHJDwbVoopWrVKJQrm/Tlkqx2ZtsHF6Fl7K7ZF/BS/7X8kC63
EV/pKdGsS9sZFSg6V9ICmLoK7tqDZgfVv4XHiczC1ES2V5pxk7K9RQU/MhQ7e7s5
PkTrg4m3aRx6G9z1QuHD6+XbGGsNM9Zd5WHt9PCI8MBP/Vz9GToKVSKAemEzel9P
3yRoJJ/TPmv4k3fRHzxErS3AeQfhLdFwdo6FVqgHspVXpa46MJqmoEDQ7agO47Sj
uo67bHW6CB8khLuou2bfjKq8NSP6TE2aXtsTFcPhcRt+zorVx6MAn5jvqANxM0Om
L147FdZFuo47BKMOG6H/Tinc9xcs9UAKVUbCdRXc8Qfp6U7QqSBgXpeP9FZ+Uybw
cTDPRcnPkAvogNt7waNLa1mDUT+DKgRN+bZerQ3AktsQ2Q0tw3aOsqopRpBNxM42
izk/Wl1WSy1iYSAoFXVKrIgS5q6UFR89+iJl+8W2ajgib3xmWJTrogqjkXY+gNrJ
ZT/PgEzkjqnObFPG5hGv7J/MrqE0xOBorYIo3OqfxZQa1wOUTKD//Q8/r2ClkNaV
fZ+clpc4j47NMxXtmjV7yK+Yr86v6VvSLGCVY+JrazuzEt2lGruH8PCNs8FiXiqp
5Js+8C/PqYn/okoFq+eAJBowbEP3wIqoLXvLQ/+3QGkDXb9FoOdSpV9m+jJYtBWG
bieUbljA3F/zXpWd6sBwLoYjd9uJ0etr3afWb/DPv2O4SnOiuttm+T+XraHSpxK8
+9OOAoxBbxj/siBfXc98KtoT7hgbrZyq8LB/0QjLYm07UFtdncEHuQ2fadmknpY2
KOvMf4FOfYzezEsDza6YaFYtPWqh2u9rmi0uCR1YhdyEkG9N+IhuiaqgixMe0vyN
wt4DKmzoBb+EY9xWIZOVa3MIP6/sSnc9m3WhgBZqyRfbIhVMOA0UNTGVxoYKj2IF
b5t28NLt5WFcHmEbgq3BljCpSPxc4iOO1ymRSuKXZCrf7/t9h8sDM80spJ+IxcDP
HAvy8KnUXh+e2NkWqrp2BsMykGe/OjaLeBS0X2wCxLhpkpIaUVMvHqTkg3nCpiuE
S85Iq/6E8+tgwCN+og5fTN0/ZTWPVJVnrgaqVNFNB/Tg925SN3tdwetPy/qoCgih
Mmc0rSd0rdz+o2WCNQpY0ErZ+hNlBpHZkAXivDXIwqw7cfRgGCt9ZM9UdFVWb7Ch
o31Opn7OAboyeVB+RBlVAGEpv9jrZzguuUfx47UFHEiSggXjRr6FWqESs19NYv6U
rxUFTXj/Ujquaj1/mbTT5bjY0wv/l23jqCSlIYfN2mSeOrCF2bz+7HBz7ES3Evpt
S2puKytz1C9iHC3cBpXrI6P2uSpIf/Mq5N+LgkiB4eOxQGrusXwVzyhgxXUvjepw
YKklf70Oh5vHVgBqeY3sbyVTjqNIq3VYQR6hHW/8hCK/cT4qTHBGmsBjp0Ppzr8s
mWo6mvBKLmanZGdKbFtceRzFDJhjYcFA5ko2WMqfT30bkd4YRVwGiX7V6YYYT75c
JPqBbeD0bXAU2pEtsdewI6XEied0CiupYCZpsZzFQJVzx9VYeg8/XBx+Rbb7zJDG
bO4RDka1urEWxOmz6O+QlExGOOsLyKXBvkzU5BnxpbnFm5EQ81vcnmQq6Fqx/c6T
k6yM8bQmQwEMJW5TbpVCfXC+5VfcSUuRJdWsdUQAbNTutZBVSOimM0xbcT+DP4Vv
rCztNyT4ijOBhdybaYI6aC7Afhj9umn9EuEkvrNRe5EnxeNZT3ap7YW/4MOTpywS
AQ9V4LOghjzM4/6dOA+w0SlOiIrJ81vnrt5wQUEYzL14PHyDuVnN+aE6T99KmMVy
4zJmyzMbY4d66jxn5JBq/T3Fq5BxEaDzt2AizpOu0OMcU9uD5birWVb7ziyKAOeF
rhqq4p9SiyBTCj4LCpjg01/woZoTtSjyaFGHEonG091V0KIr9ZgDpxQEfnYPL41V
HWfJP5MxpspTR7tmsryfoSlaSx9irQ4AOM3KURk1hxk6Z3zrFtKYmPU6PZx5Gd2W
nq2Sr+zQgNt6HwR5IqguEyI9DiV/wt0ldhK4ydVAdoKQnTezaJpmIZc0QiqxdQ5j
F67Ut8HBqVHbX1MA8O4nY3CcvYuq5g38xTRDMgyq0iMQ7U512NYamVX2anOCycRy
KLj7OCjlOEVV7lfAU4JswQZxUxehnV5QKM63Z3B/A8DVLbcAtqgf4A0rwGNPug5T
OUOFxnlYOWNT2i57+V70Tgtlxb4v2j7DxA3POU0gO+KyY1wgIAvAhT99U1jgKnjv
ZqYjfwUZUJqVNmDJbZ5sEh4vni9AvjaV4U//kuXRvZnHFwXgu4FrZgWod+fN/wvX
Z2dODiV9dOBNUZ/5F3b5SJR/sjcjyBICaKj2dgWan6kLuGBQIcI+Yrzilj08WgUR
5Jawh4qTzHJE+61v11NcSwNfZK7UxeJCSHBLqyn6KjmRr/Wk3FgU+NGFa0W+YcJ2
43ZvSIMmQycCtzkchFli7BJhxzZUMabKpYDzhXczm/CiR3d8VRFLWROte6EfjvtL
sUM6R40SPjwx0U03GMrYjgAcjRinHVbHqSfhAjix1Ug9AsVcbQDrixlm7Ms1TPor
jVmlE4ykNdqTpwJah/OVtwJhn7yiQVqHbxpZlZOSk81N4WBTpdSTGFU4kTY9aKlh
8ZuzzFG2DauxscK3uajV09zkDL+hFQdqaVoXAkNGZ4Nabd+r/uUecOWoQFJS8lTw
B0fC4gclaDcRPK5gYhzDhseXtm2LWKM/AW1ivCU2hDBEYHr7Fa6D1b/dTsepippH
3FwWtVtUxrViLzzvNGEE+iaeypZop+bPwx4GlgKAOB8jzI7es8y9J9JyHzy4vqim
kXIBcBAnOnSY1RDGk3IiV2zP2vB1ihUjHhFS+qZ21Wfk+8/kofmRZ84PTpFCUhX6
iBPC0gHH89BMuvsmEcOv0MQQDVEUcBZw/m7mHQoVg5eipQTp6iDG+cT0GapKHNEw
70bSN+68y0YmMop3pW5QDyYp6BUpyBz6sA0Km/W6RTVXNsm7jrbwC5Vf5lT6nTW+
7jJp+BGxixENNZISETLxvYP2HQvCTseuOeMFyz/XamQVNMwF/Z5WUelB4F5BEjPS
ZbGmKrdP45ehPlupUbf1NmUfnIYAxQ0gBgYPKrmZ+QsVeD8mO7Bw+1wDUAP96BDy
CizARtZb500BKQ8w4c9iTAOcFVnyjq+sX4+xeklgs6UHHw4GE3bMJDP+MsAgMGAy
gEP95zG9AM5LmJJ3cfAl2DA7fIOGyO7qMtanhVrABawr+d3NeANslOiR+r/E5sRU
QQk6obXHVCirk/goNc5HutCqlwCJb5M3yKCJ+pZirnJwRQ6BdN6pw/Fn3wL+JUsn
qAh4NTeFg+t/tyzPtvUiwhwVMGdfmMDRA6P2pRsQ/BNDd0ZmJ8tEkze1MXZeelg8
OFfUrzYO/BLqYZHVAg1vfbBzztE1eUR4xXhbpZuA78uP2uh9lw5/tV6Jd8Gj4O51
aVWFlBP+ETT2JpMGk4cu8a5ZkOsYo2qUdRCk2sOTx+QqYsn/epowMk4jh8338AaF
Mj1lctWrGadh1hIa1L0eTri6RQrb7uKTvAQ2kXGSOgCBXCMAFLFgz6Ua3iUqsdMX
yaVhnizVYACVh40FudkXKJot/nwUUWSq8zEs5qTyM1g/Ry9rgeN38YdWf4gEERmI
Riu/uliw4qudLWoYMWFGmol8cUbLuNb5X4aqOeO7A8Ou7VXU/Yb7ZQPvUeOPVJEm
IplVT7DwHQDkR6e6+l7nuCi+WDFgKX3sqY9cbj40BmlJcVQB0kBnFlRxbWIonQnm
N2UwX/t+WidEVBNWR2eMyceuPO9KZHZHUGJ90NmiC+zhdK3keWajWiX6Lt215UAD
1e39YcWAOPwj8c3aj0MEsMRRu4SeFENpidCCmSddU70i4EOrG5hHV1pFnb2SJcgQ
35R21Q0kOYhDYM7o86lrn+ulF7v6FANpf3yfJPQCZneiuS+pfEGfnsvzEZQpiKwC
V2XPtx71HUPgDP/7w6NPDIHaw/0iIvS+MPy1HbZXA5gyC9xX2Melq6ayuEA8oR05
YfeP+yph4pv7FIpp53m1JrPNFmBbEQFvItgkgackoKEjvmHq1ehDSWlYup/d0gBX
dj/uRUDkrXvAou52HOgyl6jVITyjE2xJH3PpwntdHIHIlIo08/rWNmUs9GJKVV5d
G/J/05URt1PqgIkKzbmoNRWjRxbrtEiA4eKblqOKO2Q5X8B6kY6n8gXCJvXEQPrU
c2rJVUzGyl/F9H1Jgh0+3FroQRCn6go9KR5uXXi3b5fJPd9m8hiYrZ8C1Dk3m6lq
oDTIkIYDWaOm1hxXxb48fgjEaWoGqp0Q3qXH5R8QLnvV4/ttCTZ3qEmLzKLSpq3N
sviqMvhIUDtW00f01rqUnkxqf9i+gry+sAWjQp7aijiwFZN64aeyl6D5Op8s03H4
VP/3r5rub+Azwe6hWU+YN1rCIiPfQqTe7YBcHVDrdUOZaP7Mcq1uFyFVo29LFCgs
37FobgeRrHvdUlAM9JbSLiyVpXL6Hc13Xe4mTMdeNTb3RgqtVIwRhYd082b9NBQp
4XckXybUD/nLRPYgpoNzFpcvtU8xMh/kpLb+1c0bnGevAcgDZSXtxz9En3mA1O+g
Vk07aQ7YTbHJ0QW8JOv+NWRJqRzq7hEDjOW8XKvIXE/JyTgx/YtPri3v+wUNUU6S
LZAIBk5wZgJaqCPYXKlcvoQQBkSI22uY6D4X9MQzGn8diHylYu7Np/jGB4da2AG0
JZ82o4o38jLpIACRIvrRHbCYRB3bz3EnBkRJZL5NPafDJvc6uq7+p1kKTLdU9X3i
2tAnHcH/Q7WplOq/nQ0sbkHWQnOOmPiOfhzzR2acr5KGOc5RNO2lFtm9TVAP2QBn
fJobLhv+OILrDJuawkG+0nfSLQ/yEZXIF8xxXp8m92EFf5uFcLUfYltX+yJLtdQL
VQUBA0u1byPtr7Ym5YnqFJrPRYTjZqQeYJpYjSVw07pcwCPrFIhw2cd8Xu8ZeSHD
3YolZh9a9RHp02lUZfp9cYFRI5qGdFg9Mi7TBu/Asx3EjCKbZcanq4WftVrivBHz
by93xN90iSVefO6fg6CZ4Ox+rdrkxVSRdhtfIWoBEGT55QAProNLxdZ3oldwQVkm
GFo9Ihn3rxpC+8nqzjX3gRhzQ3jFceytNmmB3py9816Ss/WNdpnochLWjt2qDc7K
bvJFOM0ac0kFfoFqFtd73ipNjq+E9TywJkdJOsYOqkk4ICXgd5GxoLRa4TioxR93
bgEVmmK4vP/8TOYleE0omug1wWi3Copf87Yaj28ouuKYRykDDzoN1/sGz6jlSCVZ
2EoYE73t7c85gE6WYfTa29pvk7WUe9DaCMojGcEVIzqhkmIBSlWU4zGDU2fV5BNJ
hitY5xBiKeqmMvSX/UPQzf4A1/eJSD2B6acIYuTLb0gwdJowANA2ByWskB7usWBj
94dy3KHivSz615tRV85vRI7OhpZGtZFQgSce2lhV6Krk+oS/wDdX7pWnCazj696P
DidEr8o9N3yAaMlNjs5LEp0wr4aeqf/8JFxRGZzREOQ6snJZoeKd4jAxTQBx/ItL
J4/jhWCQn+zYqbbLo4mmQJ9M9loeNO+jckrloZnR8rlvZoOnk3LqSm/IhWbUR+Hg
z7phJHwE1QyPtS/LxygcZ1GvFqekNalmd1UJDuIoViyEd5QFkINjDH5IuwqFTHjg
fz97KHYJnWKKwi2UJJw5RABF+2j3i8UPp2iO44IQm5pJunIMGb5nt4F2EMGdY6Yp
N2lqRmnkE1X6FrqCLYGA618r1j9UUvrrk/TGkohnCGJIbRn/SrGBq2ekEfP78ihI
r9rY2R1iIlsm7My4Xkznu6s2dFV8EeDScUxRaB/UKcxktolVuWge705NvgaS5soJ
W00DOv6fR3RuCP3F6qi/VEKc+PyJ6QtWXyb7SUCFaxLrS7GjuyMrYFkQeJ2X1JQj
i1LqKt/sjFx1o7dyV1yIB35fc3bTjXGVRxhnplBvnDIHcaBkZdJdSrxspVhVp8hn
rBG7PcgJ73bq9M7aqnKCkGB87De5QP958h+BMb/t3BLpy1owZbQ8z1CVq0+f+3ko
PnmrPT/SWdz1TVFQEvi4/zDDC7RlGmD1emqVZtJf5Cb4BULaTLr9EpoQXIia+XHg
fWSfiUYdgIIbb9tF92na8OgSu7tuUeez/+pwTozIptoktGFJjXzq2vvBvx6XCFjX
06JkuLA3Imw5QlLknuIKLjRmOOqwbwxQJ6GuSBOQMFQkW0oDB+z7uPCAXpRH1761
hk7mvtrIsi7bcSbJ3ZbKsk+bv5+LCXDKz+lGxQ19MsiQEH9KBOL9pq4R8TkEmIA3
SMMUCLB8tyLIlPwl4Gi3D4IiHOuBK38Uxt4mInJZNahelicPjtR3+W8TKXcS77D1
+qrlp4gflrrrNv4a/4i1wTwfAr3vndhTyfJdQ9Va2R3RdsfZ9fhJnppb4J3XcoW8
3YYSthmcFZUiOpGwBQL0vKL9XoWn7kaH2ERyDkHK6eC/yzIQiNFAeGj1PqQk+7qq
mpRlAzQqQYeXQBPf+9IlpSQmc5MkUgPQiS0bgLDaqekPChIo928eEtqusqWDl0Nx
9d9FkalKQcqQ522kl08Rk6ol/RQr5a4n4CTiwwC7NSUoLD+FIpAHLiSWsq+tpMrL
dIpfvmbenWQwDVOAtJK9s+jEMXTgyNI0oAfpnNGbYEBnUSBi92RvwtcxLBl/U1Js
wcq9aVhf4z/+hsZP0DL2EuJ++/c+HmS08R+ZOm/r9yVW8rNrJN5rp0LGJSvsakKO
TDoDUZSGw2BaytliivIPpR9HlIx6uqxe3CXbnveTVMzvjbudpI1vaLac3IxhP4YM
UKE2wo0vz3naSm+QouF3gbLo8bBKoC7iOZfzes5M5hnLEJxbK8d9d9oZTJBHDBjk
4bmKdKXAcqd1m8r5Zbh6t0e1iG5Yky6d77wzKxSGfXRDJKzgXj6zlctmicBWsTzX
wpHb89+TCEHak8dJv05k6y0RETIYRIWNFRL19j8PMHA34ixcw1VU3iscHWBxHr0L
ewb0pH1JZReSILna1X3Jze1tiAz21Tv41G7DH1hiLuT04fPl3lzZ/PDcmeWAaq+o
TQJhMIKmHSfnByR6XDYaEqh6oUpcGNqDLuGy1OLcdNha5HvWIKOhlDyqu/ukb7Kc
jIMxn/xfFkc6xSKw4lxe16ekQKve38qQGOcKPbCFFls1NnEq8zE1RN8XA54wKxr4
zAl6UKEB1uz5typXgkBZKFSiT1HdTXUb1VggENxE6fRZwKBmrlbIfYm1EXr+wO9l
kOpwqpNPug1bnNz5JMvgajncqOoVzfxG8dBscOdl8u1Z1UpJDfj6+xAWyKC6i1Am
CKK+r0Q8aGBpkbNvdSqSVxpONlbcBbSxzvi5sPMpwPAu2YPeP1SbV/dSUnVYG+fN
8W59w1itqs2pZgoYPZBS6LFx9Nu5KhC9JmAW0UU24wgfqecMLoMlxKixX0flxT3H
PZZ2TEt10njutORP8hlHs39qmi36mE4RKgsop6e8aVMwEQPiOp2idJ4tl7FqpYKJ
4IOhTcBfrOSu8UyfN4M2By26YPfZmtJR1/Cf3HtaUaH7gEqAEBo2Xd2XSeKCd6/R
aV+TOCsdm6SKWrAfHe/2FB9/xqplW2kBBnVYtQup/v10eEGqSZNt85AyeJCX5zS+
E4YCnCvVjZxnS/ZMISKFo0GmPscmPkAd+JrdIv1V2E3KN9004Yd+YFIkY4gBjqXi
cO8eCW/rtuILr+orywi9Sc6Vp7VyJACz5653YvdGebIbpou54NZOMZKBiDpeUkOU
1PKPr7Ylt9fAR1qQsaG7xTu6fKOKMi4ofALSOu7K02/uDsdROWjLwFF1u2h0+qgs
stigI4kVUpqQqRvPmV0ClAC9CwugESgA/h/QTAii2dKtorOWsbYzLHmcCx7wwoqQ
OKcXxiLoEQNuYX5YyyUV0mFK0sDnjy7Qq4d6wGCV1Ebz0bLT13Tcgk0JH1Z8m4iO
1yiGmpUWiK4pkZaz0E36x+mdiLKwoEhYw4rRcbTnOBdOIE1nqkPZ6eMEWsKed7he
o8OTuGX2+pDHGE1c5DPf+H2lPztk7GUGSlrnsXUu6HeZOmYlHnFbp18sshn4w34F
lSHYKyLzTaMNIrRYmFm7cQ0eUqhptLs2WH2Bv78TvlWI88QTUAvg+DQFhZodR/C0
zXXvspgEAfjxqN8vJJFRSL+K2ULcNqCqcGLMvanjKL0P4jEyemAaHDlQZQIJpmq4
8jBe9Mp/lhVqqp71Hzw6IjPVZFvjqlzO1z7sqdPnVIaUrWqZPRZQoWErfr/763Xa
TKgHUHO3Tvqo8G6KBHnPyPSxqf16+RrRNt9PT0LIAvv24d9k0TGsGRmkpM+8tHCL
1GVYNL1liTv/YbJ0RxGr36o/mDUq304lF4I1CK2bW4P/WFYO+LtrH0pbHCgN3Y1D
niJBj8DSRtcn165sMNDPb0H616rEzHMJ8+ttJWG3GmGZDWjUNmCrvepVUHUIFH3e
+jQYkrZ3lZEAk1OP2GzRso0Zrj2ovipoziDYZht4FY2av+5Gl5Y3crRXthCGO66u
/TyyRaDh01sDMPWAGC9w0rfKvUPZE97YGRyxzOuRtPn7nHIS4P3VLO6Lavx6V3bp
S6SqJfs+cYoY5a9BjApcDARXzgZhenXoJZDgnhOB6QddIwD1PhYCPiZbpOzz/Qv+
mgOuNqOA97YapUGRYiCi8v62LkVQgcuUuTweaX8nKFqvXj06z0sd62eCxzJpNyeo
y811DTq9oa96DbLK/MrCw479122wxQKD/D6IUbiwoxmDdhDj+rstr9GeROsBuSxz
HcEgX7lTysk2ZQO3I38onJsCvnN7PcqKCiUeWwtra4hedWfWdLX6VHSaNTMb1UQh
+TJ8b8BhVrpOYFpSL3tf1HMnUZE1+RnabBPL5jwhTPPr8mdJqihE8HqK32zEVYd1
o41maNuO19Sd5t60m5/6eSVL/3G4uWovGOopX/Pc17b+s4mCt6TXi5qM7UAPiVpP
lfBn7NJ3SfjKAKScERg1OlMxPL/LF8zmRWYeQ1i1b2U4Qf9qSLARrrLN1FvBIK4B
d+Ejr6NvCtipd9DC5isQnO0buCU3qkvjochczcj6jN/lXtDec10na0+YiY2tHjOn
cnKK/+IMHMD3ezEpT+KZWz+I2L7LL7mCzXXOo+YWHpR5U/DRrdhAjigY8cC2xTVN
+fvrqAndMBm/0goi9pIjcAMudCbMEnRzbkotDiIOkj+7DJOx0y5maYTizqzfLcc8
KqEh/R/RYV1h++SUQC6xFmmSXHb1RGVZ8eduIjtQMF4M9ay6v5KVyiJ2ClShWyZC
yrLwyuuzaPWJzhSZNSKfmC7Wd6yG7JpkMfxoRL8oNN2YWUcOH3E/heNfPoTxILQE
VhSZwe9YqM0/nCjyBJJuNV5e9I9ybCBpwYpTsdTEyJ2okht8fNfP03ObMOK6dyl5
vypn0D93WbH71rjkZC1m8H5yM7m9hoBHySpICo8trboiwRrXo80Cu7o/t9y6lL0v
i+Acvmed8pX5vrBjPj6ielfYPAJogFliuCywnHKAddtiOsUcoq+m2kogH62Wx8iB
0jOtvM5GqF26pM9TSS3zpmG04GJhyb3ebHE/zLBlom8viyTB98m70vvHbgtRxeQ3
0pz8ueuyowBL3yDQjN/f33XIowDN0Zd66xpxfTDYZWMG2FXyI+fO0XpkWN/XJrW5
cdTpwYnA/toCIFjBXHpq9wjueMBNd61+eJfDNGxZr0CqioWEKBFWkkHBV/S7448U
fZ+3GIOpHWJxSgxNKIBVFrTUGDfmgSgi/ahsVH5UKftuzBmcDvx0LTBCmxmx9tOW
Oim02hyWeWMiiTEJdgsAwzq9KGF4eJEJPy4Lpeei8BDpsr1fOF3Dor6UW2A2dfb2
s58sV1qWZbvHxTqdES/KKDOdnV6mDc1+h34OsQxWBu9N8M/1gV/Z1E6fNfZ+F2K+
HlCFeHI0JkwaZ77GO+Iq5bhijVTB9KT0iWojymdaG8Y88WAHa2yqbBQqLkQkne86
TdGKxaGZs3PVlqRmJmTMZ3/BRDj7fkqXSbIYuovV4QftNYTfHY5ceE1Q5C5vWJ7H
sN9icweqU47TjV7hyrYESnf3uh3XIcMjJL4wkY4Lqd2VW/n6lllSVRjioIbtd0BR
qV5Oq54rqNrwPCQyQ/D2FNoey77z1Tql61NRRbOtvo3D+/3hytbjA6CPwjhDsicl
afQrKE0qvSbqXoQw1ZAw/aC2q+O3uxpvvF9OAr2SH8omEDeMou8KwiKUkw0Ro96z
JztgiUj2tJX7Pqjmp9aExFTY0mRLRL8CI0hjHxnuVowkENdxNC7Qj+XkWDz0vvAv
beIDkfrkJiYvzxWgpuVZsidHyXmFMThbSzJQKy4pG4daUTBtYRmcD4g5vLoalYug
H26gowNUCPVAC7XzXCzVFaaV/migN+h12j14/mvvPZSkCqJbLPQlXlVZmgGWKMMN
3kSbfDWDNNb1OQQiWtBjSd1cj9LCMLg2yvtVE/1irj5UnzD7IDn9T7WZen+te1ct
qUDZBu34wssaWlCVRyWOaHNwEd78n2xy7VW/V5AmdpizM0vKb05UQHYlnCRL37pF
qTWa05/FlwnxnG77Frh2/fgWQxngfwIHtAXVtQZtFlBxwB8wDplDDrx35QuI5Lr9
V1bLDgFhLAEY80t4e8MkUZIZXB4WSMfEGx5HYekHmVysUNKSlJ3ndyQzUyXVIFqk
wVXTauZhkYkgXg4I2BN6AUrFte3ArTOte87lo0Jifr+GdToNt3QfBvykCIc5ARD3
Wb3Obe8EeN2B/pOlNyRNowpFUB/Ik4DSwr57dwqO8MolpPO+N/yIbKLbMto7fqvU
iVvXJkfbMvGa21TOJcD7JL50UyBCSlnbE09gI3vcqpa4+a7GJePhWIhkyl0h8ipa
giyHoBue/3jFumny3aral1Uskk6EwF5OZJBBXsW/N4Q6PeYbiHiVijY4CCr/iREC
qiLDqGKCr/p9gAoLThJcP+IOwtSpobKc09jZo7Y3ETUkIxrniZ4j49RGvSxS1EZo
Ghcr//bXtjYhUtbLu+XAKB2sOHGm+6vLi4uKKk3p4a6jCgUjv1iLH9Qp+lo4gGOQ
qVHtXkBtQ8IcnPxMmFlBAmIUZRFo02uRPnESki9uj/dHOFfHjEWbnHBLYKGEE7om
MnFGUyWaCqwTrv/0EGNqrHw9GEmrhGzhIqxVye1oUy8iIYgWappByzzEoAYJGdC/
STajrIhn6IWtRoNH+FD+3WW2oh16a9p9Kintaw6yBG70/SItcNXFUYCinDvY2SAD
e+4I6D2FdMGqqQkFmYqdhI7V+ScI44ZVQGEGN3Vi9j4GENa1MmhozwhZL3Ri338X
/ck18m1gRlQGd++o+5t4Scq0fc7gF7nSWqXL3hckVWOREuS6WzorceAsebmLG4Ss
rhCywv3wAoNJw56T2nuZRQxkSFEIGxYebvXHCOrc8vDvmAb61PuBE5mv1qxfNypf
VVdx1o84rT14vDG+/N1Z+ApoCfXj+pDSrPtPjqK6BqIB6gE64RQKBaAmoUeFIzPq
oDpTGM2B6Pb45jTmVbHvObPCepBGRCjG7ZdKymxA3tBs4q7byDcP55NmNVQI4jNr
V8k8OfB2D8uNgaI83T62u5gGPj6STV9pslhWHazd4PDvc+nJ04+9nA4H9opoVwDt
nCcBIEBN7iq/3L48UekWB1w692lhYzMgXfGr399tIDJ3L9yi0xC8R575X48Dg7x8
P/5xuTPhFz8mtdVtdK9P58iyGCMnIVBJZJhUT5ECPU+Go8G96FZ+hTzU6m7kqrs2
PCK7TCF2CKD7X+SSqTKcnF2EwfFNTzTHAYpC+pPEWc8t9nc/XhdkBe2Hx6M5edos
ZU5kHn3C9FxUlViVHQKS/PJg/Xre8G9qa+T5mVhipBzbV0dBVmS53qYcKsoAjAqc
cr3rt1z2GF5wtAug7+2Ih2CZS7zUCo1Jh7q92cv/HFJdN2SQTzaC8ejDCpnMImWD
9XWPdVk3N3SN2WBIxVplhKGOY36GLyQgZdDq9T1gJ6lBuXrV/9LmTc1F39L71jTT
OY+Cwb83fCOIZgfH2tz1GXPKM9269KFiAgKG68ewR1Sap7j3iR9wmXnq9QIqQxff
3kuU85YjLefYTf2PiHTj7221yDY3BxUhkpEF0JPVTJMEPdz1llnMpRjIB2TNjXR2
6wlJkkIHO/yGM0B30XileHb8o3aaB0uauLpWhK6TpCQGtT9ozxoiumjRGdwUKz9X
dkLIoVZKA89PT90iHIZEUIz5xYfDmgy6sr+YYmYcOLK1mYfvCxw0q5PxPrsx8AI2
4qfgPO0sfkmLkjQRL0sFCDrQHEOxlOYbbYnwix3C3WDeRA8UoAUAzHu6Rl9F4JQ4
TAu0i26+Da4yYLYdO6fmOT39arZZlEj1Rg8EPxE8v8loqZLjdglpQimwoJfC86+Q
j2mDhjk665unuVWhGFP53oIzPCwK5tLrMD8x8EQ9GCdtqTVjCVXd3JCRJfFZGwSj
2Mpeg1D76yP78gqPdPbtJELeMgkRJtKyBs+UsIk4Rh7H/qbvgX2cZDflYlfw/Z98
r4owFpvaCGii8SPNRcckvQXvpfi24UPh6z8102XvPxHv4TWqcLuGDZc6mTtRD2cH
/lKbgKudcYGJGwye9ENvgRaGQLEmWwkEtdwj2icsrOZKUP5JcV8Sq5K+XFXGvmNN
1kPAv9WJ7HZhKZ6Q2mADL8bddOH4hf72EOYnix1mHn/35tIxCNFuwIpZTMookIhq
WmN9SZer+0jH2Fa8acrXmtnRAeXNAw3gVuAODcQek/+LpfRLRKF97omTANsCPxK+
Ilhz3AZuWBrGvwIMSg52TxdWRbjiml+J2kffq+obNiiHTpOByvd3GxcaNnEvyEAF
sBz2gOwvZKOQMWGUtJa90sPHxJQCvtCRVHVBtQeROOgUkBZURf5+QFsFm/AeTwje
uhB4eRI22Y+iIW+3a+GgpdNMMHbkZuCZcVi1wCZ6WcblOwcPZmN4OiM7TF1LqZCA
6apc3MjKG1MAJMXXuqOf1icsVNNhcWVmrCb2RhacdcM+CjVMLJpYD5zs9oIW8OZ9
nwM9SkhDO3WaSm5DppdAdWGO8ZgHNSvapMLB5mlOacrtLQN4nksZhyJaPQy33BN3
U4Dybxo+0kzJ6mu0dAEfROU/wWQ4xeXOMEXnUxIQqfSMs14Wjkv5FwUZgrthFyaz
TsYnEfgpNMmckDve1Jluk380k3g7rEt5j7xNjg3PDJX4fpP44AeE5kMIQ3pHvaZq
3cY494wWcHqey4ocTkxP09hys7imFmX1hY+L499thzw9TGBbP8xl2hh/F/cwXU55
2Kfkr9iVyN6QmOow3ZlVXWE30nvRlwGuyZBaA+MIaNHqnfoIqbodilVlvbJKVEm3
+sBv2ebmz+l1jvPxucZO3kSLaRgIIZhHkszFSsTPOSqHun9LRUy0mAvfg9S7/B2A
qEDux7D8r+Z1OAQr3US6OAquheTCHwSeYkZCf/f7z7GVs5BhN9NFkElxFO650gPD
YUWA/ZKcTo0gsV/NQvzWsSKgyepQBa21JJlCDU7y6+MyTrScDDhsdgNQuldEvi/+
2OnL/gC8sFH0H4ASxS8hpiijGOvLTw6pu18OmQqi1PCnXaE3xqp6jh5WDyb1nbRn
XTLwlRXaNMxF3U+uyp89jU9hJ9Tzl998bLMHq793MP70zRJMUvSJIUD+SLMFzS3Q
VLGrd2cCaQJ1dCaH84Q9yaIbk5V8WID2P92lelg8AeQaN1ly2pg6FZXW8xsJKp3H
xnTN53D+mOadjFIHtDjtkEY2sydkI4p8aiut5GSIF2tmetC3bY5qVUIaSdZpVh0j
tl6UHmL7Qm8EUyEH/N0ldF6NvFW+bLGfGMG7/ntapNuy03n2gevkvlNC10BLDphr
1vCm7BRPxa4wsjuJeWQmaGhDrOJUwWbwkU/4XfA6VDDspr55dUWdAuZU14T5bgxJ
wRhYDIbANkaJdYF/9hJereE41UwEaHIU26E105hdZf7MzzoUKXPdZK6FtyWG5otX
vOAB6dOVhMt29N0l98tNroaMpwV7m23y5ZcQ0XZIWP/a7C1PBDw3hLRtmdS9tNlp
gxM0joYPvNYVlRPsF8saGSVWjx7OfaSjiahZMla1wsZEnzvi6DbOqjdnBFYnb2fN
Sqet2yjtuAA86R2t5XSQrlVWax7dxJSsIniAkIFqulC6qTC9tMl2LZfPeM7zMus/
4LnkRRnPup23uxELtZkkCJc/9TBD2ROt84/4fckSLKZAxQncsl/eiEcFo0nhhcqC
T5kWdgnAmRjTxF9xcfbQGZqRFpHV5OWF8u79hL3wklmqu4LGt8stQJOHuIUh8ybB
zRO7vRGjZDLCa61NGl60Z0Re7lN5pN1ysW+pcn7rt1/HEdZSf13nGc0nws//oS/t
3RHWBBtJ+kuLuwhakTTdwSR7wOcvhTQrciECR08hXHVn/mxULz3TO2mIT4t0r6xf
0XG567SFsrg6mcwfUU+H+tT6StpBebgOS0IvOoTQ5ksdMeB/mmKKIzO2AG/eLPZQ
jmW0e6hnbysH92dV8XvHBTDwj01v0h6Q5XZ0YZL0+yu6zqrBE0jVe5e4x5AMqzqf
iNZORxcDubIqRBIygfsC+cPQQTBRKs4EqJDAxvSu5H1sJb6R9DlTmkDRorxWHcH3
egatycT6/exWaXV9ObzOjac0m/gpYoJtWs7nPaLk/kVWEYIlb4gvscC6KDAUdJnP
yInBJQ9watRFWU3vObIJCzSOwKkrnORqGV7tvg3TtGOG+6KsGHqgKaFXQrw778y1
6iU816vCuT81tjcdTIgJALh+0jQeYz+TLnKcCpnYh9wM2ffwuN+FmUftjTuvQidX
xImV5eHYAHt6nXHnI0ELaxAl4zAw8NoO7cKvIdyaA/TXv4O+jm+R12C8cHC5LM0K
nxllsEgnOFcAur3+ybwaDhZDHwi0DaiIRVs9YCicgF5CrGQc8SMUpbuM1hmLXXG+
yJGe0VA847z9pev8fHktpoIY1xbSjbkCP1J3MCK2VduwvcH439CIy/ri+36a4RLH
Jjz3TRxdYeEntKrLt6/tdpdjSvOyAC7jLL7WohtjGln9EcPKV4WvxZlCWef9Sf+A
fWrM2lcrnvh/yk7jKtqaXxXDVeaMs7dyJOIr2+oVpuHQHfZDcch2wXruJhk6F94o
LARGdPqz3xa0VU+J4YXtair/99V0FDXzZecKtrlHpwgYdEvMNJvNFtMPqLhng8WI
wPCpfuHwYLQlo80z3f0yOMeB3JBTvIG2YFauOs6k8u5Cu0CwfoTx5xnHsdOIBR+r
lX7TE5V8yLLHpagNLLnGVfh7Tq84UQ/YeU9hCF2Yd1A+HjZL5dWs8YfW7L1KRbX9
NswylyZblSO/GxlMvQqxcIQwdOr8vnsp+YU2uh5HN5NdjdnJIhfhsiMLR7Lg/doq
1LpExZTBEV41bfk5s+xu0VHVrGwvLQHntMIbOMwnSFUYq2QTjGhGuUIxhUdAFFQP
l0+DJSY4NrHcgfZ+G80CPC08F3kl0Ha9C9Khc/hNB+6UmjzOnmjsTlO6K4U4gUbv
icR5vH/JYD0SZFnnsPpyB2euKLxSyLoSsabJjO21SBDbDNFYadZeGvSZXyNTIZLx
eIgPUAwy/RHjRVbWg/rAXzSlgKTCkEeHblkXjZokZTrKFt5gN/LOh7Umbmo78Ira
Nn1eURUBL+3bjZGRqsooftx1MVXKRiZEE3xqansYJwikKAOMlSnpvnjYWTtUlsex
mcV96xkp3aI3crv7v5eDYeMA+hJ6fZzTk9lxVQ4cp+yi2MZxbMlCn6DJaRHGl3A3
9mnj5Z6vnmPuWRYI6V63Dvu/NxBvN6kZ/K/rTLGbGNu2xCzgQnW08Cyt5SnOZnLW
0OoKhHkrQCUc6iQa0t8xoC5vQQq0POltz4PizieK2f5v85apZiJezJESbWiuHTzB
gUr2IdheRW5arbwXqUZNvPlVrBBhLUdODP1iNivz+zUFMNa6D28yWJSHxRLWKaAF
DvFSGDVNknzfqg7rPb/FxkN6IWU+qghlgHDnHcUv2VFbFfmTmzJ58xtyHhyD8eP1
sMgid6gocnxRB3PnHFWesyo0yeLkPXA2J9cqTvnLVxGDORFXC1b7JweHnERRKsi3
z51M4Ydz70vu5mODn7S6E89afihPGEXFRdQNx8d/9BIyYINL5lzYdSNRsd8zNax+
JPw+FhoUdsz1f2Y/AErClhTYDFTO1vXaxVdgagGLcB0ICLSCy5ZOuHPfxogr2sim
mGgwC5HFMRoCi2efmbTG/2Z4RSBhoZ0bHCIBlwzvd2CBcyrS04vJArF14DOaUblB
llEfSEvRmzcIJO8Yfw7b2pfYv5LM+zJhwgje7YZyBb4fTBrIG0Wzt7Nepta3b0oX
cnyutYwaaAjyWmNmOi3cjnapN8RLqFszTG0tPL4E+aewZ2i0fvp79oMi+HjeODVQ
BRsnQze9rtvMoqfyhmOvzRpLFo+ZlBSCFgaLKevDXI/lHsn5uwVOrwgcYAQWFEEj
zILMl2VgWfs8cXiYQkDogz5poNF7druZa2HJNgYCcoCjHsmHk8q26q5K7+wvBSe+
5fq32hmvKdcit4a5pxdbc5a7NPxNF8NLMtcif63AL0xNDIwn6fTFZitmQ54rme2g
5Qwrhuuy9k4aApJCmyUVvrUUt+FQcukedIZs7ykg4kjpknTxsBe2acOcODnVUyma
Mqhv0jl0dKXA5ZpgFC+BrpcbJ5uynUPwT4de596MdHsdKYdvRNYs1rCqVLQzZd+e
xjzXFPH0sRFOoFcVanf7SY7+l5eOXT7m5btEPKah4y22b5wiywrOM5uGY1f8HDLE
++aH9JhoQH3JF3qAIfDq/2Y9Ow78Ybnqo6FV86JyFESyf9v8hVB0TGnal+0pFuo9
wPHOiFhLLOIqZDV8yv2ZcrH7GUciPfqpicS6lBFAkjFM16GNSG2PF4LYKArwScxN
V29WfuWdNEqnpiMEBPDHHW1gtoOrm5fE5KWcoO4QTCKBDHdnvXV6cQ4ce7xVS2s0
K+y68w01TEuAwpqzfj50zvSXfuSFQzmIUG4X7oj6foJ4DrSHjBPt85K+CYb12IQz
FeSh5duYITmX6dKfXCktH60n8wj7QA09GkMwAzixM0IaHvfJRoXwNpZ8Bcvqmcpw
XuzB4fU/EXSh9iEwzjCFqd/3MTSmWhoWjlGau7MRKD7T2rmGh+e0mQ76qL25UDAf
gf/q6tH8Bu3y8OaDNt8Avno8lnn4N4SiVB1fRWT5xKuGJ53CvUqKMfoXJqofQbH/
aAyV7/+3dhcsu4HUY8M/TE/J6S+HkUlUBgOM4IR6mEm25ZKqu/dTwrRv1/lhKsSd
GsGnzOT7hUxMa2I5F6dyPi+dYBZoTpIXIe03IUvUSOGjmp5XC1Bu3cX7eCy1RLE2
oe9AwgWGo8Xl9dmzwVbK9WaUjXJKS1T7VXYzFgbXzFBquahs046dRCf13hAvkZWC
ajJSbWBsIOJEeq6K+o8TxAaWzgsjwr6sdhuZrI3ml4h/WWIPo40dWltbV0/aP8/G
tqWkGb94gLER+EZKpfcUeEg0h+SQjy1A4EOigBCLyIH1tBFkiQuY4BZPugdIIrLA
YkoTQmYLMaCaDqGk7Q7Ksx+IbvgBNQm9ixd0K1VgMmtcNqVGJpAkfmRqR8upDsxE
gxW6VgInnm9IVFCeTpxJp5sNTB7VW4dDgOEhE/lqfXjN4sCokF6cZGso2hwf4emI
SkjHZB3oRkFmqvj+UluPifksD4/jCha2Jy0Q4fOostVZ1u7rdnCJaRJS49AoSoCA
T4KLhzzzQcSY+x5etpDX/CDhxLDAATm2FUqghqCap2+BDUu3ohnYBrjRdeyif0L9
2uQh5cRfgucAsJ3cdiGmEFv5eXPjwg85sH3m6nx4FRL/qGN8RDwdi141CqC/ylMs
CDArDI5IcSOnU3YxKQToO1FwRPkM0iwer2Z11r+/2+HoR/d6z4+jxOXhKgXiuZ5y
J8wmRctbqHo4VCYCbInFlBOX/i+RBoF/+4hzYRZ1XEMtPXXkOQxDo6TQ6Rv5T7zq
mpIwAKmAzxVP1Wg6YX7rVV1/GHBKhSMMZ8mtL+rRHRZzCsAVDmn31JN1PlO7uCJb
CHneD6EF/A+Ss61Hu/HK1tobkC/VyNBc79Vi43ghru2QPUtFW/sY2U4ZuSdvTYUf
zvm7Mfass23WuOpkv2JYt30XArpoxe4z3Zix7JAOEHqiZkry2w0yjwUmmQIDKZQ4
P6bWx+fcE4mHtVpsTbvuhiZNpA1OGEE9VJJqCoNiMLvUPDCDZEvS96KE8ZZg38q4
CWShA/UOcvXZbTiWxq0LMAFlA6otd6WE8rI0J1X7yIDvAJrtfQXaRLlFwbwfd2hs
Jj+qgYY04RNurwaBgfO7Mde8qMrVrGDjDSce0OJAlSTcopi8UeUH3jZWtQP5iWTb
qJAqTp6wE2SlM297R6/SQXfqp+LxBB2Fdsrt9Tq9MawErPe3lqeAf6FzbAmvcByp
ElJd4JsvDvEX68vsQnhSP7FqnB4HbJXKL6XrJWdq+OECCR9IkOFxv8YjwUWGyrgf
/R6i3dgnTSDsgCFzmxgy4DjCzbIPWtArACOqutnCocCIjRzjAHMc1lNgi7/9Y/Lj
we9INVY56r7mzTWtrWVvZUT9bke1wpgIVifnKoumoWQkXEDH9WU1E7au+VKqa6Pn
7872oT+5WJ9xwoVUedHDG71iBjcDI4rKiYCPdyz0crQGkHZttPu62ybxiWK6TnCK
Eo5QkM2qVU4vCt9N9K6VM5HjfaiqvWXJlq1vIjlFAWbusi1pDpDuY1pOABu4UPXi
YMcpKn/cDQFcJo2lLZ2CavWI5862XJSqCqh8JS5PqElnx+HaNF9t3OXUlgOYBrSI
gnHtvwR+3mQzcmfkP0uDEkZ5fBmotGVr46KsZ8fr2XW/B3cMswMzZfUffgFJeYBm
jqRdC1Rk6SzdGJdfOf30mI/awKbSKjTMqor9pdtR4/n3XQpluD2W2Vqjf0YsGxhB
s5UNnC0tPTHZIgcllfJ+MlsiWiwpJ5SpqkqnsMoXrH15++Joi/H+f+vM509vDU/u
jUi5JydQsus70PDLGHTCtARSuDePdfH/5loO3px7jBrqRj1imtRrx1g7NWVIlixp
CdCdzJbBlwbdcIo54VT77WtfgaSyWmGDSO6z+pYYM9AbLrfFlbQ6yktmk3F28ZD6
/momA4O0cHAlQFonwD5LS7/ow/CBrMDMqrlKaMldBQbBGhdTOOQOtgCkPszkywn5
CU4K2MS8GelZfGB/TrK2cUVxrOzbppifuMSSbWUXjzoZX4qDwYRMNSHE2j+shvp6
BW6vcaVFEo+THqxmbx7HBBU/62R4K2HsP770s1IPzEhMf+r3fazmssoxRkCTNv/b
hB3E5oDd4MNHzOIV+p8LE5RBAbxYN+hiNA1zyCopCID3kzWW1HEvNYdc5vMp8IUh
+K9trUUY20R34z4hAtnxM+Ef+aPhRkC+qGwFGbNfkFa0193SfTLG/Dlwvo/vJSth
2VgpjOS5+DiMVTAZJ/JXoaaenjaKh5298G72xNlhxciooS6CJD7zZs5H23NybvJb
dyTZo66Ca35S8W4R18c8edlIWrKZ1oGyHmxwxMSwEubfO5SYsAQIlMcm0K90PJpM
s4/147nYbEYdbifcRPvIL/IHOE+wuTKsn5vEfdcUJ9IGTEwowTvoRWyKzrjIKXI8
UdOs7ZQpaOEnXAIjRaqseehLfthAGsaV6FUQEG4Aj4DTEAPtUF12B+t25YLiy/VH
8pFSAbu4ZnCMVh+zDpUA6/JsPDVlafWnsA7EOPij82JilLgQxY+zztT1gl+3d7pW
ctaShrfHX/Opb12JiqKVg4qXEQPgR3uzGReOOPakjYtbKEe8iorYWW2AR6wMIZJ3
WXh+riaNXN3ARrKlLzBmljjN5IBPlHbHP4+MKJOiye2g6j1uVxoJW6I2IImWBWWP
rY9XYfu2WBkOlzDZgKtEEvvUlDtljfmB4Fogw8bxx6Pr2Zz5HgiCUyA5+aNSNo3E
xj7Hucoj8If7j1NIT+6glaV8SIF47loA2vBfItiLDtOUEFg42lsKv+HcQtGzPJM2
lj3u9Ntf63kcSGGHSbfBjadt5yTp/3KAu8S49BMo2mAjXiFTYHLz8VBh6sqneFZl
V1ACSuN+8F5b3LxwbvT0wHlJVCfJX8MKqqqPB01XR+zaYJJ10dqg7N2Pi6jerhap
HUuVbardxsAX11sTDYEEhUBWycwwojww8nDVaoM48ohL82DNNxA2l/VGnxuki8Ax
AyiyJl0PCaKaXZhoIJbPkqqi+MDiVddsa0LR3ggTVPK2x0jVvOQAG3i6sp3PeCZ4
n7UAhIS55Llv6+F88tTvEUNYcG6j0jYMGQYSWwMGo9iBYSlWWhOTA9TbYGtCCK7L
glpVF+iBL+zbC75IKzXXXJDpSoCeJOYvFjNs99nG9Njx0YrNcYD7Mauh9sk+erqf
szBRQyLWMrgUI0JokTrQvtLlKk0kcBAzPczkutrpA9u3XR3Mgx5ABBNQfuyEu1v+
BzjXKZnz2zruMG5NLuC4YqitsnCoPic+S8KbM6dNKsLMR9W+1T/g2fn5ghWEcwly
JMNEdU5pUerjc90xQFnVbR5x0QG4ZmqHVhjzgWU8Hhn/WcinY0+QX9yGUsJ0iMGl
FIQUFH8InHif5/lZvxW1CJfPNR45JYr+sXiIBpBxJHj7MTigkYh2/pzMarsfQ3Ig
QbiJLpaDGSMyLdWYf9U3/DpEwPjlUrVSVngeOZdSdJI7/L6ZCJrNFGD/HavyojDL
frxSQ88G/JYAjsxRvutnr84tM+WYUege0pD3TQ/85crX0RsSplnxj7KX2xlbeWSv
XvWjrrw84MHqcke4NOc8mw+/DnADHHAia1kIbKt9Ox8d87pRXesSpTiJN1VMMtcD
lcv5flKE7PGt3YJuejL4FO9ngwkiKEw7MI9u5DXQw+A+aPemZxQ2RI8ax0XN57K6
+DMqfmJ6X/gm/Wi5v5A8+680/kFg8s+AWlqn9qvvc4K1FFtG9R5JJUqjiTJvUPBP
+QWKlxU0orRwJwK4ZxrSJk8XKrVuxEEKx+Ba2oKdpJjBAboNE3KSh11zSoNt32Z5
8xDj08ZaPSDfN4JQEz1ypM9Y1m4ygxX3kdRwGqtl/h8tLCTFnxBOxjKXaSs3v6Ij
DqNFbX9Km0HhTc2ueNCDKDdzntLEX3OptpynUqZA0G5onhydiplldG3mMKZnzHiD
QO+MijhFWxwK3IneseIFq6OpwUUhepLjkl9FFqj4Do6bYyvFbCr6rQlvE5x+gX6X
wiX8RXgVcOlWtK+Q9KoETw3aR43EUFh++jJ5ZGO1k30DGGliAjukywVGrIFSI2/h
Fa/954pyhOp5OaZys6Yrc6NsSIU6qec/GmS1vPawB3QcSpkVHUeVs52qTDeEd+kK
/YH4NaJAoDQqE63UJi6ep5VMdxUDYZE7Bpn7TbB3xuYtRMqTnLc/pVo8Pf7lE43g
7rpRYHWIqlXQPSoKr+bcwE3bRJzSWs2E9NXUMi6DiJd6hBEUjNSi2PDAdFkFh9Ad
ZfhLz2ovH/hU2EUDSZxrpmKphN87Lwpcf0Gq/Xo7Y27VMbUta8O/nD8jKByZePTp
CHt17iHQpQaov0yPxL2OfEK4hDwVeJXYYPa0LoHOjDGaxBM5VsGtXcB9onCkwQNr
KqE5u8yS7mfZrAtbSm9iA9UgRV7dhgZMK5cKxTsWs2lXBbkd9yuCeSbG2sg8z01Q
O2vFXw9nGEVMrH9AVIMm2/XCszKgcAHeFrq+fDrBNB6oWD4PX4X8SzDD4gdeH2Ap
ShYFYMztURNMQLEb2f5GZVCiiqo0QebtPKIaJXgcBGxoVN3zdbajR/J1dFNlNLHf
BSDP/mcutieUhhBnL5YlJnIUTqukN8uYgza6QQfXOfhs9ljkgO0f2lME3CFl6xQY
GnGDx/Z45KIzvl5UqcxbD/k+PedhNM3iV0N6Lbxpb9IV9PirD8MDyAoY5f9g0NiW
gofjpgxF5Y8yi5qGMGdDu+7H09wS9wxNEtwq3h96qg907tWlxiuTZ8bB0iIws8Do
UPOiuGg1lLRyO3N8lLcmo0DUWBLv5DjVSSWMxFadySVZL7ZvBXdTimJYtebIxKW1
q6DaG2oLoxh2BZxaju3g9ePR3aDDUxkPnGnX4FhdyyiuWqHWdO1EXAicbqFfZ4wn
Yh8wQMhpNp+oOtnNpEgR+W1akaqepPuvM4PSjjMclJBLTcE3WgYk+ty91ivuKdU1
MEJd23tfdMEc0Z/rk4i+MfXMxTXUIdVdN9A2bwoh/gBuZLI77vlCStlZQ5Mjes3M
+uek7zXr/NGVPeHkMY0VhmNgYojJj2Ecg/zAZBU+xjakZ2l1Nd9fx/Pw5fHb1omo
Tssy2oN6xbV6UM41CcSuD7XmlAhgLn67ZRgqOboM1UpV/Es5nuPbwwQQY7QHr6Vm
QpajTgZscYOngNyN8PlLYZivJuO6zrh+CXkkd7w16Z10W0s1KlT5b4KWv8d8ESXa
EOgPoP90BBIGkAzmElNcKLyP93G7RjYS78w7xWxtZ9GoDgrT9l3q4FUDUJmANJnC
Ys6iw5dg+9dIdHiu7DS6Gn016quyr6Mz2s1HtrBqwTJ/yTykxScVcj/n86vkqlBq
4zbQvvb47CS3z4/wygOn9vg2tTo6uTwbxvsiYj2fLl2BVc1PrJ64H/+LUJS/tj7r
5/4tlGqZAW4b9xbx4/y6OavTUW8dQrggFjvMdW5/f48ICIELNHpu3BED5B0aZmSi
QVE4n4w+sgSOffmna+hs2vm++/3bLYdiRSCVA/k0ceUGzOGJgVNK9eXgmFjtqaHq
SHUjdnszIGE8jk7DbJO7uNPXF1e+wnnfgQS9agdRmFK+IQQ0rZ3GMcNL7HiAuLQb
klb1dFclfxIcECzMaZgNSkqLASlt3Mer2E5IEN3WMG038/adOJgehA1YHeTfKcy7
17tn3ZEpw7pvuJ+XkWxyd5mG4Dh5cDoUjOm9j0obqu89wg67oNOsvP592dF7LOxq
SFYdGFNCwSxtpj/a5GNAGITSy4N5iTBLe+ytlLzrUs5OzM9DkA6Xann6D7EobWv4
lCFPWrFeJqypUFHjDUKazmDc1Zkf9BkNVQDQ0JLL9fJRRo+8G8RupQyIQZsKXRL5
NHE/ZMAkX5fyWwCoq7RM36DulQpTBoSrQsV6jsilbr+AO7zYUaiDntB9MsP0tHfP
g+35llJplsBORK9mbLGuEkFWyqluloxC7gpREQ+rTpFFeJJZUYB+5245mDGr4JIm
JhRw8yVLzHHN570AWhmqtliwMXnq8flLH0Hy+3LUfQ6SxP9sNrLY5B7U2pFl9b6X
tInTTZKTvRSlyXhmjyTJpcgruPvXUA2TqosQHM+Yx+tLbP60Ozrz8X2M3hLH1ujo
RuOW/S/NmzvoGaXxx7eyvniI6++jj+t4cZhg7yoejnqIIKhTiLFKbh1WVGqC4hBR
s/KxTeT2SoaOmQQLp7KtuA0yOReOXz185e6cZNe4VrXEbvNS88AXnUhw7ZQck0uB
cVhsnIrgcuHAm6LXcdlx5Ar9qOHtcigPvhG94rsHftP2rlwx2AZ9NqN7jt922kWd
9EzV2y0oN+bBtc0iC0vdBO6cT41RSbkspu62msPsT5SZBVp0FZjBfL65TgLAWBT/
R7Tdjop1PIp8DTiXknBYDfQ63hl8SRY6Y7ynyz81ZO31x/q1y4t/+hGJOkRwJdWs
LQSzbJXaK+WgAO/pgVpZHtCEAZmtUTymBrlcyIJE3YO0Z9xQSL1eH0PoKBRsMZhP
7b4IgES1MgotK262pjXVQmTzlRjdkPOI3KaYl2asMKUcVfhzq+dkARkFM7U56Kjl
97kBjFwLyovKYQwMOAvoEeTq1xgTcrsGWvLLPUy1tLO6VnPEXRdi6dPE3eU17HDf
Nppg/fo0NOYIx8Chw7fnOROLzbZAqjBPPAQruWPmF1HPEs4aIuBhWg1bfcCQgLm9
WZFCdq8DeOGdaKu2Mquv/SYMA6l72OAANegiwR0abfphkhyR+mQSpLT5BnN24ttX
a6z0XGf6g0Z/y4k/q8bvMr1WAxMyYmcSwZT6mDbJNj859dQbzlLvqY+HNm4YdTOI
3VtPyBLDhVrQtpdPkdiegqkPjO7MxywK7bxcWlRvl1/RAyGDtJDlXrEy1DOd/vnI
BuB4GSUtetsy2qRGx12hp9TGFxsMkb7f0Z1ATZS3kucZrZJzJveb8nRP7Hc9uXok
ZAEzz7eKdWIMeV79LiWVQi984s9xKFYJTqZVd5bVCaofqh2N2w2NDMK2Cdojegyz
6x+VDL1bu5rGXivP9kTZc/ny/PRM8XACmyiS+heBgcUlFACpeDqw230bmYxT8Wal
0iLlGBYaeSe600L/Y08AizcMW9BilKuFL44cDzyyxVvBXKBno3iBTKRrVJ3bxbzt
7/Ac6+4oWZXm/NQU8npTIhnFMetsXuAq8iY1urrTDRcVzn8rJA0zVZMcLzfGzKWf
97scPTBYysvXNuEfaQSDpkfq7NlqH0z31sNOiqvgoY2ogDJjmWpdI0EN0w2gNWBE
KDh/YAakDjYFovssEzY73WTxwGazclUz6PctfCNBuTiOFMInztbjOZfUmCCuh7fG
QlfDh4qGFPAOZqojBeSwAQGIN9y2oahH+fKsgh9jgRl0aKLg67rB10ByLKCRq9cA
J6s5DwYrl5fg9JFMfNfwUmInGKQmaR6TOAx7QiAkf+8vgh6xNtOtZHSdm1bYNplQ
7HTs8xZXFx+rEE5vv4YMD1RsLkLPOg9UGiTXOkv7xEyLGmJfnanW8MsEmCQnjUp1
Q6AkLeG8KxxX9OXM8heppM5SO8HTz5eX4bHQNCjhSCu9dVxGXExPrZb450xDlNQj
BY3jl5abY8rnT1IPrlWFUbrsjbOlfBuvHNzsl9KJqr/Q+b903q40lccOppMipiX3
AMD6r5l9R5llne7ppqOL3Y8N5XI96HXtn4H2Ct33iXp7ZTRu1SG1BiEvLUvigWWD
PWFL/wl+QvwZEcpwoz83WbFRWQwhtCoDWb6JE4HSMzLE67KLyALjYs8KhcN3z31I
dFEv1pohl7tM3/LGh2QcJtuI/8wwXJHA6dgGxIce1bl03nlzt3nenXQcvBiWwS3y
iWUOrFJR1tDw60+TvVThzCL/DOVNFdQZfFfXtfz9Z05onL6EbaFvg4322U26XYLH
aiDU92WEX0QOIO7JlHABuNBfoRr80HWfcIZDgFvfrX66x1CWI3ZniEWXYvq6rVUG
+ZdizMMsOuUyl/PrYqWhcPg8dwFqLQ9Dtxnurl1Bk4q25qE8/8ef22FqnfPGPXsU
vpT+Ch5necgoeXhic+hHiFYa2pmlrbZrCrK3pbjS4p88vJwc/eVlT5IHyTeUWKkS
f6Xbu/iFuAKujvCI6o9gX8I3TGAyRFkOufaJXapvYfCewuLuBeLdpl4tphga2EUq
QWiycl6eo58nVMnxraRBsW5b0suJjQ6LPnY1UzHiQHZOIwz7r6DOk/f5W1wboVDi
HJmvfz/ZGlXtrzeJuCft1n663Sr4O2xYsKzyz7bvcWBUWqFuoBvEQ6LO2uG9nzeb
T4dG81UuE6nMZXJT9LDmsgwHG2DWvzm/zmujO7z/ORvqLLdHGpfeusGby7LdLVO9
QQ8powH8hqkU15KpIzA2DSR9KT4rEB4dj+uwRCUb+/RWIHALcw7Lktez53Qsxc/o
Gp+WuQs7IXqAW+/shqm4XjBCc3+4APCNgTGEiYGwhCmEpHTdU887i0ApvEErZn3e
y+SCL4Dp4fBeYdT4pudmC1VqNihknBk+WnDrJcVPX3QELli0X2+9skv4TV785e8j
JzDUPe6uKNZdbFQRWvFIc3YS82d9kEbjLSPzITMxqfWNgPWK4lDSMTHMXngiAJvp
KLEJif+XBZ6vNKERV/bj7hgVSnEleT9Ot44QAh+z3bQ/E+GuNuU5byv/h8rP/DBC
N+rvpqYI/Eu5HnHKlvs2FftFEmM557HflA7CaaiSxRWuFS9dgoEb8kZlZ+vW8QYS
FRrl1rWrLE87JCYLe0mZ2kAKg5dwwATizFp6wimRI6O807YGf4RYcYSmbtmy4wLA
Xb/wuNkwWYdEClAcTN9gNZYYIw5ev0fd3tLundTvVI2WMd1lt75hVxOZ1nA4MJyp
/nf9nE6TskiQ+RO1YtpR0Wzxq0RaQ3OOU8fHNsm/a7GZW/Uv6Z4wWfG/i44on2Zt
nUzRbbuEQYG6AXXCPzPJFL/wf2jVpKlODKG8L+gTtY0veK4/cAeHDHKkTsSSlkfb
iz0jXPE22t2IoaImOkDrOOcLjCf+O/ebhDLgxYSrN/1zKU5rBQYSTRvnN/ykq526
/jOQo5l6Ng/TEJdAaXeIy4sXdTZY2YFRmhCl/sHuzXG87tXSdwPPhPWUxNmpibin
+jFWOOCODlBvQc911lnwQqWIYVrGnrldckymrFJURvkhJoslWd1k+MYbi82eAxUF
vsTdv4TfnjuRtN9S+7UVtw3PjC47xo4/fvsHjFJD74xG/4612Fcm8omFgbYzhqS8
oRtX5jHX53jTO/bhTsAdTWcMBWKJi8WslGF6nHiZLh92Gspy2q68PHsVWQqkOgzr
rc/cH38vmNVs3g2DkZbK2Q4EsDluFL/mJDMhPdeMjIZGzbqf2Hv10azkRdLN/Tnx
4PQSP/C3zFu4A0IGALlStA04QUz9c33+RdzuxBAOuk4ie5cCYBW3Xim4ttpwxB5O
ss2IeZjblkJXRTbGk4rlsWBXup3V8MTjbV9kUC1+Jj6A9Rrbm5mIqNmCwCdMHNKw
O/pRNPhRJyssDOodYU0rZpX/YqIvK+cWV0cRmt0fdbcGMJtdBRjD8C+ddW7lwJBN
uGtsE5LZNjjSb2Jizz9OZIFxK5ZRjuwI7GgvO3L9aZ/NBU9XeryLJxSR8B9G2VTp
uTOcwyLehN/+lZ7ZN6zk9N0KwQ9ODJ2vCkF+VyGbhzt0i7YdhqyK3InvWeoEU84N
YTeFdL9Dt3B7TG9AOgGZVU6JEdJYwaqOI811Xo4z+8oFSRVF/jQbtztPXOGsPg8i
7FI3e93MrGox1ov13v1MfMH7bUP3UX+zKN/iHpm2MOmySwMxn5O5pUOXrfZFtcT+
lzEn3sBlZsK7DCjCCJL0nSjzxZz8D7eIKgWhTti9XKMfN76gYUx9lQZ9Q9etqlu8
mfCoMjaS9VX7x46C4HwtzZwk7ssgMj9T5SMjuwcvPa4nqDcvz7o1tfeCZfgyA70l
7KiYPXCtCKXS5KejmwvSkU/5cNif96bSB0UJHjNayA2Qfjy5nBPACMrlbhLfHOgM
nf60VH7OauOiFSC/iwUI6ZrqaWRoBOfzaYK+0xAedt+c5ewoiVJBDDysSqHVBrfK
oDj4vobHDdzMPU1EUQTfdNzgXBUEebe2N7JOCKGPKqWZFXO0iqpXqseyd7/M3dgj
8rjs0EhwYJG2YSzBvrb0UwPVx8cX7Dj+JZ2/EeCbCc4sApqz4b4tA8LOzS0Glz1N
WoXt1pu7HJQQJhREkcid6rSWjw1+c3IPK33uzHGLtAnFd3Qn6yJaD2l/J5xN/7kf
38f7wYWeQh4BaYQS6giALH1mkCKazje5XcUiBBCLUn4cpgSrRuY9WkgAbYZ2NkwU
PxVaVCELPUC2yRADnq1FrlHXeatfk7PvYN3ePcDJ5+Mus1IRZicm1J25KnFhTAOr
K9cVl69vcHWgOn7qDLEVuEJiX28RlCaxDBKGNMG6sPa5xMdQ7RiVx4lf8EQecQPR
oukrs2YH2S6d9026qaJt4YaAcTqmn6lAIgD7sHo/wFynOflX4EUFb3Y3lfj+iC5z
R8P6uiCBNZOaP+6+3wba7yo9mQQrf1Py9aIDSXKRqVIygRdliRCOgbL1QcqoYEdR
C0qH9QiH22kJS1u+nT/Os96pKNoIcJj9OLxoSMDk7UaqSRCk9IqBjdg4D5I8BHK0
YQnGro/zTiOJW8BF2ZW4Y3HoWEuLOn4s6v7ViYni23J5IeFp4JenFXsA6haJD7EK
D4sP1bZQKsWuLdbUIeCzysMZHx6F0CklbhHkGwHrbwy/AuahK77GEkAK4U7H9A7f
JwilYYDVoaPoqrHQiUWQvufcX54dqwbHYCRUOZqr1tWPARZlV93l8jLhV4P7nMvZ
lAHI64wYKLmUT0kUYzQI5QtaCQOQRlzznCDXRCom/95v58PC4JFLzmQ8e/n3nKcI
wDp8pTJcTDak+a+BbjFgOn5lrXMIPNpdPojXvPHBoKGlRDECx3j7vi4QQWS4zfzL
sUeuDe6Hi9WuJqg0RfT+xlbTP1wnR0wfeyIfYh3sH61Z9rPgkjE/xwz38HMUeTIP
65rBE1qcSuglaZSZOO4NRKphgk2RmB6h68NHIJX1RecgUnjY8icfQqHhvsLiDxQQ
SXV80cbrF2luwVwm8gppM4YWaj6lP3Dx4A4B7lCV3fjQKGCDEYvuXWrH8md6pqCv
edjDTgp4K8+0n7chrFZWqC0eCmJ+vXUvjDhC9EU3Yqi87ttiBtiVvFmQntk0mthA
pTHNAK1nealtE9+hP1XpJ5WvuoY0RZzQfGdTVZ3Nxf5VXSwLyn3N5hgVPUGGHk2J
aejArru6FvJts68+tOgpbGrMu6hVEf5zt5VPVerFHQxCHXD/QEXVDYcVavyA1KUR
RPnnWwSHQ/8L7/IrWGqhQBcMbZ422sQCOQKPIlOY1+EBOIA2GEtx3b7tkTibePbs
BqtOmz5zJwsY3UwO6RuMISH80xKc+sPOjGLrIN5NJjoS/M5rfZN9LpueEGKZHWGZ
Zo87y+iaEpeqMzqRgude3XLxTzcgByFQjnmZGrorWeRmui5XQQEjuDIc5w1qMQn1
46qK+YLtGqWmCy+1ojJo0XMR32WfcEgpYVBbBlrgqtFdmBpRRp3cPGBNV/OSFalU
t2hSpKeNwOw1zdWy09J55sg0IT3aBoslNzIvI4zLQETBc052YFLO2ONPFYHxc+k8
Up2CKi5ne6WUFAihCrcreZUmPR4uMDffufIj8PoHea6KpTs2jIo0m9Dg6gZ9IMrn
jtxsJCRImNz/4/8ADZ+HrvnFl1CoEc1XNw32zHOnEAGxjEvL6NAEnZOucT/Zn5G9
5SXdeYDmLwAvrPJ5ITawwrhE55jvR3LrhoW9o9xJ73oZU9BdKZXOMQo9FJ6rYIJc
C0eul4SVzoxmXy4+9CmZJhHHIVJxK4dqJTQbRquVW9NAYDSdKrVALp4i6+hrAy8c
MwfceFXHUabAnjs4qR9U19GnD6dtuj9g6Eq/Cu4ROkUl1iWDuIZwMFJ6spWxjP5A
JlghECjBDsBEckSnl1OnEskNNxPV7qCo/1TW1uFMiJ6onmcxOZxh1araGVR74Qnz
yzw1wB7Ke6vOmv0+Ws/yxrTxYk864SIxq5Z7eSBULtDu2vdgdQX4ux681JldqHlb
2RKDrKnySSKN2lBw0LOAW1OVd6YE9H/M+6YRNiRALk81S441ls51a6zCwY336rFH
akqJYP8dcUaWIuUopg2HDeKw8D0gGESibS+yz2G2d3hSyltQ5lrxT/hGUaX8n+mI
aKjbttKkUp2576vZY+ySCFaKACtd9O5/g2E3/geni7YDYjNp5wyPMYWz6xNo4bI0
kzYkMNQDGC1rTrxGEs8r8+x/LTK1rqq6Po1FnicdFVgT/iRAx+a6qm5oYqULRiH9
KVDy5jsQZvzCRJab2kkk94E6X9cGFZcyEBbcky5gHdIJhn+7EFaXy1c6O8TsZj3u
xYfBgCmKwdjvUaj/yxC2+DqUX+w64rC7beK+VDL0i6ox63VnkI9yxLDu1w0vYNYk
d+I2AkQV7dOQZ3zZ27oEP+Re25OZQv2PyDmmF78XrE4C4j8HXvI1tRVu68H9EGYn
G+yrftLk63TYh156MYoV07Sqg+dsvCw9PcM7FcCwNhOARsJBAY8NM1YSNffxODtN
zgEkfZhuoolUkHp8IOp81uwWv9sOmijNxw0TNkP5C7sy5Wi/j4NF3BrHjtc9u60w
ZBPOnbsiCbR3NQEB8B4Vy3DuygvYKJb8lbf7jb+CwDTQjlJvUZJP3EhoZYp9wgfz
7C0oma8aPpv0YJTcYdV/1NwVS21FssBxQNKZLZJplsy0hO2RQwqIAqXBBTzGLVGJ
PfehBzSF2GsziKTO161Eo/qwTBwMxB2IG0N+Qd1x+pLkh9ZR6PfRbIJ5635kIdin
sQXaNHAcmHKJNVGw+6q2rxZfkBmnd1y1GtaGR2EXDIuG1mL0QZHI5H/iqWiBMlgR
Ds6xEe6O12+eZxhD+hUUOBY86Mq9wN2kpNUzqG+LgOnqjg4ng8R1dtv3UQ61bmUM
tLoVaRBRwJq9mimS8z23oNcxvvZULKDeMG6vw4PijwZhASJ+Z/s+ZVgoCTM3W41T
f9ZCqw/efiQ0zMj3OoWiVnzQkEdg00aOK+rXRlQhWgjmpZQo9HEURBZNuhQ/R86N
q6Ll3wVjnW6cS6Gig/OU9AVlUvBvj8jqzmmSipVD4cBVSXfQ3AYYe4aQmoZ71N79
FdubSC6ojTKz+k9NR+ahhV4fI+lD5UfNf006nQecoNwtlMVZSEYBlQXBaK53tWps
oGstmyNvSbwWl//jn9MJcm2tKWOxagFx091UemRrUPZ3b4cuHTeQP52YVLFRa5pw
k3k75d6fy/AjKIDg+p1BMOguxLyy9OXUqhIIH1kToid34hRyBRbxoeacCC1lPyKi
IdLig/660WuwrZNbUP+zEO/cjyD2UP7zWXxVCaM21sYIpzttnF7fA94xYFpDoQbj
+GYoFj2PwevflrE65Q78Ef7qAnxfnApkmp0ZAdEM3TlqcLMm6iVl1mIdbxthypNq
yhts1KYIZzTArMXy4CxOiTMt+0L92WJPxoEzkrvPqvofg5rWXhrhyDFU1wcWHpTO
3KiulJrPdQDsirh1QyVMzy69+1Ok/2xnplr7fwVSha9wfRA08WxtTpgQD5GVv2Pb
r2OoNgaQ/XXmN2crR4z3WyY/8FT6jG6zq/WTY8YCnWkebQBu/JjBAJ8N675I/Xqb
/ZUYpWa/uNgdiMpLgC2RbcjakgJTZb8icd5Lxfe61KwVKCHmykEqL/7qJYDKrjtS
Te9+EVH2arWILd4bSSpGieoj1L1N9zGTSuHFd0fUnaj+1gOjtMtCHuCf+y3xqldn
U908YAIbbz+gNZ40knfImbTmIZXQGjpSxX5ghccAlU7idDigR6qa0Kq6kTlBjsoD
qoDys+MfNgHrn/M8Y7Gx+P87YMV5tD8Hvj7VmCUUpIHwmQifItlyHCgCYV79/j65
32BgcJRcTJSdp3LDgKi05jtnsVeSy8W+ulvsTVoaY+8yGcuPAiBlEol1lBrSr0bc
gPKybXwQjbJgkms15fnHdHZhJH4l64N8nPfhybUvvjAY2h+WGDQmEilbSid7lAo/
s7hJ4u/cbYKksxVn7WJbfwTQAC7X6XMhUidD8kFPNM5HZxPUjpBOhSLltgqmiT2s
rAmUwzehJHPj9+iQ1XbrCg43DzzAxmpsVlU0sBT3hNkgxqy0HMgRqCGhF040N0H9
OjK1qhl8YM7Zy88d49JPuGUQ6QbfrZdj4iMFwo2QQ5ozbnLMVChjTyBVAHXqkriB
HKXatqKUUyQ2tnrxPHNOiqT3IKBM+6bzGdRfKtSYzXXBZsB7G5QZXmI3F0fxwYNS
VrTSd+tn9X+VPWBIiPAIAetjd8NksBn8P6lg765oPQihsrosQZR/mqMa7U6eSxtK
7N5S7ashwOV4b+6El+BY4I2JG4hZEI8KUarV568pRaanYO8rSS0NxMlWzVAUicBC
5FmzQS+G1iZnYY9ez58sVw01HP+wMRp1ZO7QI92wBhTOgzaBsrBqqIwIzpuRTobY
+vpQPbEPMs1QAGIKAxZEoi2ozQgithJxhFH91NaqDxHTM5tcQ7gCeYWJa9bEwCk0
y6K2mK5m0AOFRMbHX4Eq+28JxaZs8z8sRrSsaKgDCB1Mhe/02dsbcypOi7s7EYA5
zuihahZaZX4U4w4F/IKkHO0bQkATipC7L89De3JQ4KYP5UpSRepamAOSgwEFP2eT
QmaXyLlaMgvMUTx2cOKGpm+85UGPJohVzUjJ/Wlqc7hP9qKG9+cn1taEAMmAKhD2
RMyMUcNWETwm2yEQNucOpCj4xZO1zqrW2ze4CPo67AJnUQ1ttUt+RrcIMUi3UI72
+QDYyPT6SaZSRNVpKIlp5Sio/4ewysRP9SN5k59DM03Y5vr/T564JV199L2wT+IJ
YuTHj4/2yWBU/oqanQGKxtaM8z8g7Q9RT6jV95+5Vml0FVSc6e47RUd+gZuousxq
cWXT89nJ/gOG0RPXzYpfB6MpUmMHkFkg7MWC1uecV1Fkdh2EbTT8tv0nv0UIrtBM
a47xacpxJNGWBUEhLkOIWoqw7M1lb2JDx6PTrYjV6hPQkbIketQdMpRCDcMezN2H
KL6TsahsFD9qbPyPgOKvbLmSIHTH5FHpjxUnn3+eUJ6n+MsFeFlbDJiw8kEgcojm
KlGI7zAQ1+I4kyEHcNmGtWwwtEV/QXEMd3rWd1MNdJRJAom7/5w7+qM0+SrhfcKH
vwwpwcZneSTIaMj6baGd20Yt4zhyQxxvWu7D7j1Rk4XN0BC6msGIOBVZRokFIWrs
GQEeNQKMMD4jLjihWIQC2U/rY2kYQFb7/sSgyE3jmwXct+EiIpC3blzvypBwkPWb
qguRC3R9VJxiuF0W4gb1w+Z/OtoLqRcqtjGF4raiii/ENE2917PKTpM0nOkTPBw9
aIP7e8ntw5ueHBointvd4iBXfvx4/6kq8hRxvZx7pRY/WFV+LsTyBj8G1aJa6qrr
PsizulqyfQFiVXM+UATU5gqiT4Rwx79c0RjeOxDaEm727b3PZEgWw73Gq5DrFTMK
xqKQcSGP1TbqtMjP/XasTa9ncK0YWvwd26xvhoKJhT6CKN60CeKrUCfXWLcie8Xi
9U3fq+ey1+Ng5C0vv3WzE+M9nvzpP2tOuVEQXIxYKe9RpZI0dWtiGnB0S8efuZvv
vKfagw8+4LraS0REILGk8ObiRgcktwMT9frzGV8Epp7JowFVUYtK38KExTArX+LN
1mIAnb3mbDoLQ7Le1tSnBkyPjsFndD2UPDAoMEDp4fzT1tgryhONaBXHx6SRqZIF
D5AUUcCw3V9/HRWoWhzcnuGZo77Nf9QFUo9E3IGvbNgnXAKAL/cf7LSgNUo+WDCS
2En8Ah4rCnwHUNzSQKHYJwylWlY0N/vrAnAUe8jDddfk05S14nj41wG/rJ4SXFId
7fSKIu7uyWDh6Fz9YPI4J+tkbW9TdsglnwtzS6/O22EQDdO5M3i3LRfOIMSnOUyO
4qb9nbOBV69cIeiH+hhDskCrEZ/PR2vAbuoh+Vi47KIDWBW31kkSkvGsDsAjP6XG
kW67nL3To3kf1UbP+gZtWoWEtvSQM2bBtSpYOnBY5DaPaBd5Boi8wDNXVcoCiLwj
tCJQKXWUNdefJeK5FyTSyGGgXsT1QAtb6w0SVeaEbuWxippGeqQKIdb9U1zHsHJZ
USQMip+1i7mMl6HCmqZVIwMhMFfWFcNDTrtP/ebjAqn00INpcgZN/vPj91LVYgWB
3Hkxw//gi/65nakgFaZLGbxQT/GnXQzaauHYwkyp3Np7Zk7FaeUTpXmet71gI9WS
qd0yRn3alskTRnK1D2F3U5g0GCPWgKUrSp93S6kh72ee/cqG41bt7w/NNf9RfuPV
rMErKQMbezJOFTKogYhUqqH881MTMwP4KriH2Rw/Fn7OZ6BifqXV8rOin5otbUwj
PZvWvGO8vVqgafSkYusui6D29UWfNiWgWLag1u4x+gFvlJC5ChpcSEttzvX3yxTt
AkSmYr8C6RqEQZbcQlJJiz5LIswV6bcg4Jab5As+qORvPRIhcSXgc21AtipLinXz
730Cw6kK+cW4XVfNIyrN6L9Ov/PbEFgAiwKk8n9Bg3Nk/5SWJr1ktj862pNT7io4
X3AIl1IDqqFVbWzkr0tc0EgoNqHJx37GjZTZ7KIueAxFd752zUubAozXm/o7nXAx
5iVA6L/mMeJ/ZTmgmt3MuKVUbZQIU0ku2hY83GFWSwET+8Tsw892iS1WSnMwpiND
RUUFpv5n12zIXWtgKCWWslyWiq7xBQKNz97gihlAzJ/8ICg6clty1ynH16HIFzjA
Mc5o2o90bgZmz6icB08X9PxxiUE7LBEJnPtGIi5/JeD/lXAOGC0ivartqHlW83Hl
3BXyu26yO3H8bqRnf6KGDMrNx51rcc5zPia0Mtz2N0usgiKHozFAqajmW3Ufrv2b
r/BTYnGNvjXYgI22SJzPcQ0GPJAWPFAkrUJlm/Ooaa5obLFZPPdTA35ppxhkO1Bc
0k+lQd8Y+Resjs3xj4Mrpb5TV66GjWqbFw/VRBSKaHRyAdjYm/wjkQBV3Vy7wIjV
Q6zC9Rn+I1OIxgJc88Vj6AtVQ6J2zYsiU0schXBOByavmJRR8imyaZ4PGWQIotog
7h2K+Id6daEwdTwhC4FB9iXZ0AOd02XraO7mhSDJ+y+o/bfIG09uLI4jfEvl+j1H
EEqbgbAonq+M34TvIFVANvcnhBerTvEkLdff4Tb/Kamfzh473WI3YX2eeFqEIgZ3
x0hLiEvu+c+mE220IrYbNXszSoshQCczW4pFAcmXkJNqQZaUkQ8QQQxD7UxbuJUj
svdOwuKbYRpyYExB/pI/5ARSK7aAweyQCw6BzSSgvZ/EJPhFPhZDZEnfbnvAFUJS
0tfy5zu4iLVgjFquPXguPR5XaLKiOFqHjuxCQwce4/MmycCIj8jbF/y4lWwaaW0s
6B50UBFLe6/kII3kBf0KARjL17wT0ABGAsWZPK3BmXNW2sK6Vw86tkRkR1Hlp8Uh
RQmeJIi8yaM2wrGUpIyxy8CKi81yeN8jiU2EC7DzDNt9NSHi4Hp5C9n5nKV3MNpL
69zjtS31yBvg3W6KZc1oRGk+qCPiubWroH7XM3Z1J8qRvfGtN0snf6PzmAcCH+cC
e3E3s7ypVJh/yVkyHsWFqDP9Vgt1rYK6uJuz0A5nocVwSYLdvLa4ZfU4EdI0ouQH
FW0nZ9yXL2SV2RUFGN8m+WezPw2Ge6XLfEGTgxEtAsrHo9+a4p64oEYkuCvBHzHn
Jf3YogOl9s2ws6dVzx8G1eamtlxjcGkj43P5K+PuJTVJVza4sQKjvByAaB8dbbB7
8nAiRN03GmBCp3HwCVMlZRqvqeKEgsY5/xJNZN4KUlAiTKIkBIv/5twspdnwN6lF
jd+r+TpCWNUsXwBH9+U/2QFml0kzz8xMPVJs1MUoGQ8GshawEB1lIacjGxkFPmkz
D7K4/zz3Q47ajoMF2HikhfJtNgTEv51dfNA6b6ak524WLiUoMa4hAgpFclE8FZb8
TDlgVy7eySbSIJmzC3i+8tMk01sUsUGr4r67GOFWVkqroOywmXnG3EG6lbyYF0ys
2Bw7jjE8nw/byhFmDy2xwMfAmhskdbmsb1RzryYsvND5H/HxAqaKUH39FV78a44q
L71UEVU5xqDM094Ju+dxZ6hQuq4Q0St8H5meRkvcNAKGxwHrGM4GniLJlOvlG3iZ
ZzJ6Np/n7Irzt6CGE0cfRsszbSpHGniRqcZn1kk0pfbEBk6Pi3kFcMbUhU33ipp+
4A5rR+OKXrxx1btw5fTM8PozPgyxzakygzHabq+bxNWFniY05e8SnpwfEimcDCAr
Oo6Pv5yaWX7hh32Cg6zMFeDtxINT872cty//IFGkua0c5BAZmZhmq85MNi99UORS
/mhNmO/PJLcocYYpZ89MYi7sSVFfp9FMKEp3AWr/6I0N3fxlLr0qsBHYIxENf73c
4eEWPEh/ksgi9m7ET0k/9Ezlx4N2he1/5MQThvVIctpopJGHtAfeKvG146PB4bhl
AxbUrTvy/pg3sIza+rBbd9JEih9ZFDzAM5hVvp+QlIXO5hK06k69Kd0SjVquqSB6
ZxHfPPnkBCKnR+FLyK6kOMHR5xrV6bOn0rtldfcbFxFgAZKVuEe2fG8YNPyYKk5Y
lIoQCH8GxiXYRtTgwOiQjWwOt7YpTNfmh1EIieqE72jeg/xrjnuWzy6K+aPnv8po
06ial/KCYSkjRzJca4Hp0TUogoKYxY9lnLc77YnNZ+3k7UBPUzLlcxnXro5Huet1
lioRVwT9Gx0uZ9abm4BZqkJ01FLRxu87CRi4x5rGKcRSCelt8ByGT4jsclauPieS
UtBsgV8hLKN20PWrQ8bg6UKZGnwPpbl8CQnD1AYP49NjZKDrsZgiRSoqi6Ig4yuY
77gfHCZKoVRHQBgvVCsEXVAtHX6BxNpfG1peDVjtEkbstclrUzcUjGSRS9R3yvvt
Hil7hzkuRL1wxeY1vOdRmDS02rvlV9cm9w7/qv8887TiyKLPwAcleGQiDA+TajnF
IKFsdjI2mgOcYMwmQRc0fe1OkjNiBn428SxBiZHJPv+UzwMQqdMxpbZC1pXI4OCl
pQiMGZ+ITvQGsKQsHiuCtvFTziCIOHDVlCTaUolDHKWcDObQJFSNhuIcvBzekvv4
FfxgsIFYISxlwyxiEJtILZeeyWWzTJegqr6qHjg0my1C9EMEm5hvIkwsFN4tvkXL
7IUK+PO0tBZ5VoYgJ1baO2T8hkQDh3F8FPV8JIuBC9zjyzCgXyC1C6kYPu1J70ME
gNc3l1e1F377Qm1oMY6IOtuumCV9ji1IEOordKAwGZr3u5iVZDjhvlD86kQJhj/L
hHzIf9tjpxM0zdfcyCz0+1XAWHUPAv/ahtk6GC9gKOm9NA7uzdFpBsEL9Ti2K1ik
WVJH2qJ+nWUNYHQQL4OWnLelbOgu/lnEOUInUrchm2tQ+dAt1VUbi6Y90afNSHol
OWdTnN41St3p9mJeMwAggxnzbS1esm7I0xOcsx9WeHMeiBI79gKBeJ3a7UlFsFWk
K/QyPP1VSI7K1QymTvSPnqlvr+xPH+z2mtLMs1xJJ90X1OVcnloYO1iMHUUvSk+y
rTp8Rq7LxRDhoGb5A7slnTN59jdv2PlHQkncKOt5R5Dwq9je5K2rRHbePH1ZFIKV
um1hfz6nkn5v1Vo37AbcawKrDMIO4KnVT8KXs9IVgqCZKhXgSP2Kt+Ej6c8E1Gok
qCAKiXlXNxpW2BMEuNdnkEQuOUVdApXWyhmx1Ot0vq9r6pTntSSrU8G7CDraRpj1
3eKO4ND11giSN3wQMGLF10RZ0YZXOR7GqLt5pGy4ezFfsDyme+eyXKvCv06mHRP1
CZx/6RGAEZ2MUywCb3c9A1XBXneyJCWIJyPIp0go1LqlwEiVlMqWy+4VAEXz8r6h
AWMmA3dAMI+XsJbGhxnie/5f3kh64fvkwJ4cJTFxkiNE3wHI6lT+yYe8cTjWOo7D
UkCaFJEyvoMoMEWm2+eS6ynZQoyzWZbqLroNQHYkDTiZOkeSeMwVo8uk1I/coWsQ
8BcAUu+hWI6aveZGvtsF8zDzso+xLQyuTN9mluYXeDZHCFxl+uz/lv1zCBV34tUR
m87twvhnzf+ESTf1DHV1eN15kLKpocxmwod4IQ4YmIiI3y4XlP3otqhYr91IdSvl
IWq9ODpRpGhLCtpLDHvhPfu+eqwo3poDZbdEeochvxMvUrg1ZKJxg6Kr7NXZVdjv
CE9oh+8YynSksdrpQ1cjEziftG4nF38XUUAFLUKf2UpHHfYEq+yo1XxPh0BTKt2M
sKvLHj+z5XKPWqEEnulRlOfWK3p9A38d+OZ9GqOwix252bQcV3ibRmShIsIMpIwU
nL5Wy6au/tI7T0I2ETIp2TCXZGo3TRpFNYw0RwMsg/NnT+T7W+MzfSibRsoDTb+G
QSPBHAC0i/qOlqyE3UxYyHRfvEiH25Ro2qOwbCd49xxRlOhAzaR7I9hyCNfv83oc
JFhBc6RpG6K0kpuUGU2oH0abK+5hES6L7Y6MBc7Q36LjQYRHBA4WKfzR0dSoI175
YEcT/Pde/24E+u5/NV5M3eEQLJxKCmsdLdlg8S8lh/QSbWGgbFZEBsVnBiYBkS8b
KMB3cqMTXVsuorFJwV7Jg+XDYnb8dWE5SbbIQ6ngoCjU6NVudqFGXgqEDBvnIJ2i
wsUU217Kq1OiR5SWhkHOCTVK8TWmtHJvE0x5QeuC4PPNUY/6guTpNKhUVQ+VxRD3
u4DUc8uTuzekUVM1xLt4QMT+cciRZlu4NjoaUCKfkb0V6KujolvgcGPe1cFxQI7j
DYBFEmYlMNSzHw0Rp1ZZ9LJlpxF3Wde8OGebASnrZYfcw+/ZjbLoKs3glVJpdQFQ
+6yeIgFwXtzeJbTMzbrlZkyEpwTJ4+biNNlxfh/NO4FyQrbdeFLIfOVd+bfCKJwT
Ty7WPmL+tvie44czCfaSCp8irxlsr0Wg18UAmoEKk9khqkgReuW2SyD7jGmnJ3/5
E1lkp4mzpffQ0jTGgLJEm1ajcAjSgfNTmtOXV+tSL8MAxd0ouLmt4GnK+WvB3lnP
QcXOEwZ3LQgpaBEGHEJKjma9pHKuTIbiBBhvi9sftO0szzcG6JkB7QeK+bstE980
Crl1nNkbKvBXODQwABe1l2gKvk7wO4286IqNfO12ugWNMDdrXcm6rb/nkVjUegss
Nr7j6iLaM0PtYyl8qS3ouH+qAPke+oZsHbUlWZZI8ZZxCk4b0fS2qstV2A0MnZa1
PouvDBb3EJE60YwOEQWh6yfid8OH/aLkcYSdLhSzevH9kKoCO2H3xb8F9kmaZyMM
r5Zye9eNmdETfyzDvIpiu+vrtldWWPo+dLMZVBSACPFb+WZnnm/LMa2N9Eai77NN
Nnop6WudGaWkMxEzUk1Jtiqzc+opnwKRJ/F6/rm76+r0CKWC/rohMlyITMwbTl5m
YfRAVykojbS5dflbUxFnGWRKpMns2R3ChyMkLr9uqTsr0hpvjyOANAJaUcQF77C1
TGHqWX1rel/GafPynnVaXIN3SGQOHU6m8BQ9hTmSkyDAH40YbPqd5EV2vyvT1zcO
4yb/Y/41wqRH9003Xs/1KZ+aaib5m3JPKFgiyJiIq8aqJSHBtVJ7z1BdkBy1WmZB
JDu50QKiDvvrbCFgoIG3DIYfg5GD3yZUf/NFYl7JFvilHesbKP3bQY3oZD+NnAz6
z6RjV483GgoVPIostt3PhWTMVUGRntHWc9OY/mcq7Eg5Fzrl/7Y7ckW0Hgp+XMxg
vhZhwP5kMWwRx4pjNaUsSCf/vVMla5X1So6kI/Mufwu5vth1aMN2/9KaRMx9C3L3
CLV900ejUxUlCCmcbafXCIFlPZxcVeYQyF3el2sT4rcRGEMJ9dvYW9E0CskDPk8E
igqWPXkg2n6Z1WvI/jX1yKVLEbmavSdZ3i6kQfqtKaOa9Qmt1r5XoecgnKhrKB45
SYadVLOc+NbrKnMm3I0H/Th/DEAjLvMhmDUHhkXeWmV4FYe9Q8ztNUDOt22CRbeo
upk9Ru9VwqifvAylXOTAd3VBMr2n0Uj/kmRa37vINhTJP1rLHNDSTrS4m69Tw9vg
uFso8iQ/ynOi+eS9Y1/vqtZhebV/QnAryLOcgNXVwMULHlENnZPM+BF7lmNBmcah
N4+HMMTgKi7BFGrW3/o5AttpeUWRby2II8smMDf77K2o3A3GtWh+Ad/3YfMtPu08
sNX6ohKIYps3EIWMvDG1tmDVPxHYS32S1Bko1fRgQfdpuXBPjk/hQHmTbWhS3BMW
BPrf9g826TTQ8iYjlWe1LAB6qCxdGVy89FeJUQ192dCrFeTuaUMbBxIuURLYtwtR
LsLsKCzX9R2zNgtkvsjvIy1L0WJrl/hnaN8WJ6C8G9dVx7HL0+yW05orQhNuHUAr
DQR4j3K6C+tODvgXi3RNoN7AXU+oEymDRqvnFFMNf7gRQflT7cOLLqg6Cof2x3Rx
Wp2PdNKK4iuO1Q1P1M2QZL3ifmZrkYBydlZKD9wIj+v0ssjqTPtk4lPdqpDLUjDx
ZI9+i8XH8vUZQLZdOvJ4yGOChD6yIVmMzptZgCJagCv5BbPvLrsULpNQpmJu8euu
BIWKPdSWQpwDMj7We4aNqjCj1njv+t0Ata39GjGxgp8cTz7xTS/p2qcmpxGh6Rev
SbeN/QIEs4bmLl1uhJ4ZN9Ov1cvAHLJZMAqVx1NzLlfsE2Pn7LsX6RRJc/N57aox
mVlxAH+Ol23asz9bmdL6Vl99lU10thwLRfSOzx2dUJvIQGZSAmqF692J5uOX8avn
CQOHuRXjn7zOhierr622MM2qYiLU5fswJM5JGX4N/xU7ZiRdEuqqBeRiOqClyCR+
NQHvgCiRRdNVPiwj3n/W1uMsZNmuhWPJA6KvwhaVvZCg9RADnnr2hHVBSfipu+Zm
tjlBl66PsMeaqWFvLla0t2sflY1xng7LnrUi/0cqKqrHbXfniTIKy9EEhbBcD6JD
fAtuj9JzRMrSsUo0eI+SZCa8Rl9QbkHIkvgdztm1JJKrZmPAPmeLUpmYGDOKVzog
wqC/wmmmgVLLwn8znUdZzq8Jw7hjxwLnIEgVR7hU7pnNl592r+tE1f4pR6P2AzE9
4O0lOSk6NiJoU5bOS35DDIbzXOR/fYbmkK91Mi0MbBDh5GHU5L0OywY0K8l0AFeE
9z3Bk6ToP1uQAiNWcv/o/AZX5v3p4KWFwB0+4vppb5UxPIBasn8kkmDoDQBJ/tCK
QPQxtKHnMLA0ENDjOCKyRt83A6w/Yk0Vil9vdKQEmGiXPpNqoJsAcsR6T9Fi4W8f
f0+cyIB/ZZymfo0gMhc6ZglgECFdDsPcDdZczckPt1+cKcyVSsBMo7Q0XOzJMwHw
yT+svhcpe5kGcPhu9i2MnUPbPPy6+mKJ2Sn1+znB8NcPkBpWskqGZAUU518lfyrr
yZ/3Xw0JSE7gYZvWxT6U7lAJ5d/tUExMehQnm/IH4cvfrPXqh9GiIiPUzAEYdDoX
J4FoDWSwboEPRa9LEspBMdddbfsahW8uApybLzgY3ZXtziauO5gfSsf04IKHACVb
qBvUMwGcUwNDj4IMcTg7tU4qA9RGoT6l3qV650rKEJbyYsUJCb1kUP/W4vKdwi41
RchYz+J8J3TCDY++yP43I2L1Pn1ut6joCa0WR8FBATOtbKi+NtsnqPihsTXnEipK
EZX60ES3cCLWeEyTUqL+fT66re50/5CCr8G003AgGrg4kBWJNtfO6aeNTZZvyXCm
3utXArpH7jotT8LTtRbr3rCGh7HeGFatq8wJvNbk5P39ZJhNK8d9TpJKTnQq3GNX
kS8OpXVleKACB2oSxCXimZ7b+FG1fwTVRGFS3x78qGXsKyjhgYYv8SAI6ombm1+b
DXhvuwh/RmA7EUcEj9PpAe4U3h9BAAz4p4YevtKzyz1AwdDKCqYLZsUQZitaM/oC
6hgfrKQdm2FhT8i744e8U8R+d7twD45+UEN9VX3q6+Rfp/MApsTc0HAUJhoW9et2
raV7HbiXqZNLkRNYcYmWaq56NuqJRn+PBgOy0ZDTzkbQ4idIu1g55eSmQR6OxBf/
yuSBUo+cW4BtT+x9T6EJLrwS+iLLqXyAwHMKbzgtGpe0BX9jxRy5Y9ZQscABmlsR
jzGmMenzQRUTWnmYVbmjsFiIRrTHCuiKyTHJ0GI954kGQwwxJlohkCzrwI56omf3
N/KehQf8AppNeBvp0qQX66SsO3ZY9uLJc75GuqjUUaRcg+WAwYlG4U7MobErE5sx
gvX+qOQ57Mvz5lYJSo3qXP74ZHOG+W0C6fXlPEj2pEHsulkTBqUpvsyoQlM1IQzF
Brg+wOYgepVvrONuRnNBypRauO7L/9z0OwvTHeLM0MKISqKQqksafm7U4lWcwMiV
hxU9Zx9yJYbqM84EN4aMmJvxFQMS/g1Kb6kDxFBbOq98iTJ9NI5PY6cAUbr3B3+e
L64IfNeJfG9X/IbYiqhbvq23OK+Fg6fJz2eYr1odK4KakoWtuU0LbCIsgy+KatAP
pd7gn+mLaK6I9VklAHcIhIa2Uf2PM0GvNTkMt6TAHh43fjx50Ut/Id6h/m0HbAL9
xCt8HQwSGHT1OJb9cZSq31cqsWyx0iN3ZCYlcx/6On+p3++8j5g8FGgJgT9zZOt1
xhAR7QGYq2+IbSnKN2NCf2E9i0C6P13hMl/KTiAyInYzukpgKWhgxPeFIY4xUF9n
NnB3ZQ6IhIspBxhbD1PB+r8eDmXnQ35NOftDkt4hHye3GkSbdzLOIMy0ZzyjucTR
pi3WDBWnJnVWr+5ScjsWqi+pNEREpNTQ7z1g8dOk6M9Jl7yKuFSdGy6W8XwJfWtl
MCm+qyerhKR/V6xFP2Wx4/i7/uA7VPJV7Ca3AOQ8P74QvuWMGknQH5pn3lj/lZWc
3blMk7OLPZa/wf2DEK447fD+crMhjF7I+1lMcYLNvqK6No/dzVCg4rl7Y8II8JUU
zSUg/pdHXA9CY0UD2JawZLMF5t83+KI3e39V5TIE2x0LPLqSW39Md7QwLbVbDGXY
QocO8OwZLOeC2eSFXxTVsyKYHkTX4Ers1UznIyBR5EqQYPDm8vlERpjvUPX4g8Ul
z1q+aWqQtCaWIZoV0wqpX9pd/Gc7dhEvOUo1+eIFc/RgcOKjOOVBmkeeMoLP6ygt
f9rZ33HeC4xgJjx59VsFXPhljBq+VNctTUUlQe0aN1uWpYBkainKoWL5iI+NYPSX
W0FL4nVb7a31RNjkJtU/3llHQUOa+r7+u1giOi4bm5SFEmZp3q31GLasjHeRWIFU
dsf+bSxJT65sD3KS0N4ezYlhIrKq2GNoJaY6S7GLKKg/wKDkJeDDppLqaLblw4ps
QbBqufjzPC7mxQOPo7GRwS4KDLsex4yeMjRzRrhVLSTusRp/loo5NIjrXVqOYzH7
FG6+u6fqT+4sPAaX/wf4dx+JGAMWDF5Gs66h18XYrTiVryA2tboQedPsW3J2O0jA
ZyuaRWb3VwGs3iHKWOViN31HxXWXDMWalTkSKbXOgcFVHbPUfI0W/wwxbDD6Nn/o
d+HFovsWLpa7OipziMlPvCh/ytyGhN9glIJFcGUE35qgJciAGWoN+RfDUhiw/74n
30BmX1zP4vYIlCse8T17xGjP5SzHgyFU91zKlqVgZQ+TgtptfGAfvbRbmlRPSd82
mElZqFJDuwt5hQBIK9S9YTfJkdSW/JzR1zc9/7BWXcv23gcCzxV9Lcu7eN4Wn33i
35bs53nh5VOR0Zv+qHX33RkNyRknVqbY49YBZ4j+39m9uOv0RjLdVIkihMvLvJv8
sIQjs0lzd7A6PQYizRHexOxwu15JJv7xx+6c4NTpb3LiLd+Q3jAFhB37EB19JZ0l
oEe/CSVi5ldi5rxOojoB/js5dA57ipRTJw230AIlLH+ZPXzlZxxrN4JewJHepfIv
ywt9lhZScLDs5gnQD2IdZnQ0ofyBoV2AntQWFNGklb/0Ya9TFtowvJqxf+a6AxKJ
mdltL2SIYwNpC3w1DeiUssF93+mrCB5I90fc3hnQbd4tYZ/05djMaS8Fd71U7fz4
Bc1Z0J7WehDyZEgKlrBcyaujHbHoNYW8hv1iTlA8WqwalPxpH1vmA8b9eU3RcUA/
WWd6KIqKg42JrFyK3HY4tfNPbzXV258e1EUqGCyEd0aWNZ32yfeMUdGJC5IeUPM/
EJrIl+Rv7p0B5D9b0UQj8biJ0c34ULzfJRZAX0DEGhi0W/fRMU0+wU60jPZmEBnf
TqR+9UUZaEdXkRDsrNfGmcvhW/INlU6Lxj0zdt+aJcqntJVTwU82X74FYwoaaxOH
EesvMQnqHEZt4OFh2Gqf6Bih2JKSoKKO0LzPDFJcA/41LiXFfex7BFXrujm89l3S
i373dbX7Jta0C8hEGrVBgAvl2u8n/rGc5a3NCCGUPSGEmia99qD6h/JzSikaqqOC
H1GGDW33CQwM9ouEbhGxFPhepC74ex+c97PVlkO7BSliUq6JjgGf/ArSySYD7sLc
WZjnK3DuQcu+pCA2a1a6LKCotD1QP9zg+Nopew8uB6RF9G00fBr9bg/QF4RWmybu
oynx+VuAkT+iAiLtmOi+CsIP65FXYplku4kotP91mRwuil6+6XqwvP6GCx3Ibtdr
jAxafXTgTSOX4PR21XU/aIokc7BrM9qT3vmvP7ZL7WFxvQlskD7PFHOpKlk3VC/T
hB69BCyU6LMByU45o8M2SnrRiWvprMfUpxWAv6B4FKXOeuJ65aeB7MhEyzaKPNQI
VVH3ThH0UsR8P5rwMkgXGPJ2equ/puKvgmaQ1fkiZsVg2sSWr5fU/D53d2xeQSsQ
gboMwkx9c4O9lf/C5shfo33uhAqYjaCOhfYpZOgtSFlivhWrn5Www/BdchSTTzVb
Dp+RKVFq+ZPxOXz1hY4CsNRnUWFWirmqcbQxMNhksGLxSx3FMzgOpDBZ2T5LRftO
Lno2Lgo3Ok6sI6hIVMh3l3+soGkeInTEXqOd0Yg2gwItICnODtomnThaJ2MDmG3X
ryFQurJzOnyCQu+bxSKg70Apsi6040JaoBS+jYlJfGjXXiasT2nIENxhMYhHBK1+
IV9K1SI35m3ZC7eFEKqvJw8eBDUq6wix20xnx8HW0NX3S046F49Oc+K6ckcANdFf
DnFmzs8W9p6MfS/XKdty/9Yri0Ow27fcPeUWytcZGL42Xh6DtwRUfvW3iWQrpB19
Fd+Cgt2q1gygzFoYr+4PoSAd7oxBG8OecgPsafB10ju+LV77SutSHde9jxKZyafZ
n9dlqWgQNI8VN5aQIvGVwaUwTVGZYaHvEe4g1b/TGQKCNt8DhK3rQ7Z3x7/+dpPA
vvtNGw7SH4agouBq2G6XTqQ36kqUU/F/Ed9nw4Z+85zIonSM3rN61WP1+GRYSg80
3ij0rfleuDh/BG+MCUJ76MYtGFuriNj3Of03r0qt+sRnUBt9h11XY7bef0VKKmei
6mRIKiwtRSPYvU3l/rO9HFE8CDHMQQ2OIlE1huCc77QN0jIkgHfvFyS4/YAdKrVn
9gmgmxm3COVJ5cgFm1/NXY9x6/8XyLsubdI/4qe4/JknZacI398lSN7VuvQXksW4
+ptC8ANxuM30ymVmmWZNObcqPUxGXjrjTVYQ2RgGWubp4RcPe28cWrY40odu7nYe
O/A++O2FoSMkQ+HnoLS2tLu2de+RsGiV4OLJR1JoVlUfctAMhAKJSS+X/y9V0nK4
PddfZSm4+zMfA+5AydiLDQpKrin2SRdSv8u20GN35UMiO4y0d+mLFCq8z8Qsz0OL
LaF2lvqqlX5161irZkcbnY96ZawDnBzficWqJSH81dwNGbRAx3xKqjmSXqBX039X
Mb0dlF2++IDkqFHP4aYDyL7rwGNZpjxDdpigMVKlYegSliP7FR2qS+d9mNs7rkYQ
2jiJ+3rh9caxIe1/VMpJANrh+QRfpRY0IgDz9f5hUkrD4J5kGsLl03EpC6rIRNaE
peBUcqFv8FH45jtoHNGLblmrXUu8wCpb5btaqEBtoXbN8C9DE5tVHkdSdKEs6qf7
kVv3fcldkOW0f1pC8LokFKYYe0dVQnS6hLJt2FPzO4shiD++sX5/HHUz63NQZec/
LFNtqPoKN932br6EG2jeBPZEeLScbO6oXzr1nj4+iqLX7Gq1ZHlofYWpBgO58hax
uALQZsFhY1AJ7k95gECG0HnNWFgs7UHBo5/6qtAjmBDk/2tv8ZQ4Y6A0utyc3TXe
P9H/AQIWps2X8tGmdnGJ6JWkgawRU/tkubDkAReV16G8iyvV9p0Jmz/qskbvzP0C
Y5h8onrlQ93ICqyqOz4jsDTuV8ep+UUXLP3dXJOcgQO7gfQlVFQPz5c7eWqEzOg3
NQf2ZvthI3w7yYxS5garYCZS4Sp5WNTA6D8LkiejeM/BG2qrf2tkgf6Xf18S0ljT
eQ2HRk5qyps+OFAiJx3KrXjnQSyiJaXEXXIGIPSLDgBkFUqaZGbfm4QsExZ1csKf
NV1fTzaHOOpmNbNMlsKCMWJavYSc8KRDgWqciGlXJ5ivrjy8ccFjq8HS0OrLM+rQ
3Fyvez6ez4dnuVtHVhrnyIgqH9BgY4J73R8bflov1wKuWEIVF2g/vMp1XQcZjy+R
5CyYcEjqSO8Hy/dKoHRA0yk3Z0vznxefkDu13Aszz8tXQou5m6/Iljj3QP8RzQRa
awTSygyo4HvKTduW10fDZ+EvuK24JJnrsWuhjzZsvb6Mpcj6errjwJm4HieKbYzV
hJN0N3IKk71hCvVYxfCK4JGYw0rTT8Q26HBM6HkfwD7S8iOCobnLH3G1SRW1qSzU
4rVAlPJXry6iPPTD1nLXLi5xyYg8OX1tTN0aMMPrW5RVSivP5rgCdl5woLCfuBDE
ThYZvBRnEQbl923jhXngvmHQHrJMWb0ZFpZ1ovbF89qYJRLNoL19QlcNjfxwOSzm
TIwENiEUvwGQ7Au4DpvZIoJG/1Y+LFVZD3HopMlhQKmz6xSUdNUJksZgZ0bFpaYn
2KgLinsLfe8VKJFVK0IYEw/GxFUZpOC0EEYPVeBe+iAJgLe+Lu3HfGrLcHCAYnOl
NgSA4SB/DCXurClOCOvwuzlxZEyYnQPisDLmRNrAg4/xHjlA3nVsjN3gsEJo914P
reFJz5VP+xGQrccAPpHiIvxMm5mR2PlCWgPtsPHxtSs8o3Ajc39Usva83E2wxhlW
Tg6OirytsTyR9iBYqmq7y2owUZK32hsFZuOlKUfQ39zGApMF0f5uRIYw/VfMnrnm
aSpCPUPisWJaFnlsA88XSY4hJw2CE+d7OotFLPPUpTXfWaIBSdqzSalmwXtogO9h
wUzHuBir+eTjmyIhvwjRB1BQqmHlfsVvkKlIX/rOEq3AuZcF1gp5Z/i1dcqs+d2i
ufWyjhpwHIAK6uW+SgtBZ8UQyR+4bJ53tcF8sCux+utlcFNbIGNoMIgpyg1BN2UO
b6Y8VmUrhBIjvETjU9IIs9yoW8/vI6/S+xYVoEwlKrAOcZ54RQI6LATUeRv+qDjM
4u2D+0OBH5paynd9z0tRwlpifeEy+AQE/gpspiwZubt09a9H7P1ZYZ0RLuoqelmD
kdXi0Vewuy+RiiuqtxmVQZNoAoCBk045/vHxpkbGchYmDygOrdS3i6g1jX4RX2F0
zecsqaFmJcqK7KyueYdQAHAx3jxpdq4hiJUpuuLcfMBTQIL3jot9CKQxSGGpVv3t
eSiiPHgqRSFEIO6UT+Q1wkYNS8zcNNIS20nFtRhTE1epaFqrKlXS9HaNBm5bISpA
1bdb2a0prP9e3P3JUyfq2unMH/hictHembRd7aRTHFJ+wfdTM06SYacgTNh95mUo
XQN44cYz6PU5vUg0asaVV6EfHhbRY0eEwpNHOS3MWF0j7NCHNMCtsldRqwvhRufV
bKgjT6SqWdya0HU5bPTakxZFQD4n4AOa7YEPBwrW1zrLF3lYPJnIgPR0yRNNiS1W
m4kVuxPwFrIXwx1IGiXsiN0oldoApDvZDRYQTJybR5MIjgMUnxx+glwA0iC7GTdZ
xwYQhIVypQp1SmQz3Pf0q2hxuTljM1GPmOIowcQkIAArTD/BK/7u1ggiYV10B9Bw
VrJ/XaSb9JB+Rr6O44rESFAC+f+tag+t6EWDodlvm4A4ke20X81bQO2RC1RW2rc+
mRcBkMa+3vJIkPkKhL/46DS3PCeZNXNiqhX6BzYgaa84xEPECMT5fsmsd83rARPZ
F3Ldw4R9cIs3nxoUAhDlq8yZzg8zuQ0sr7apQh12zBkYFhJt7X3ZhEKr3KRmuDZz
YshTLP9jpmn7lOq/GlpGZwAA54abwSEaAA1mV4L0NjzMTNKZq8GQVrsQCR68y883
qOr8OAQji2r/IPMO51jXJyTk9VqB3u2yc4QfR6f2BwD/kdG9IGZLEwAdu1jOiL9F
gMxTWhSXzOZeymelzDSKiUEaQD0ANWjzQUtvjnf/Uzg/A8uS9iazJjAIVjfOp7Bv
qL1kw1xI8JzPoctgrH8Os5sUI++tXgGePY5rJUehJ/AT8CHoep3ez9Vv85uK4+M1
h9iyi4P48cf2dcgPreamRJDphLZXA6ZIJeocRzB1fogIQMGZD6WkMJITPB62SSAm
Q2zkmuqsZHFv7RbrB9hNgGRuGZVrk3nkyLawvk7AI6LKmYEwJBNZZmgOhOs7712l
lthoJVJ5EdeVvUTcBw7VYSTQgkWvN77/10CbI7Nm77h6vbxTxTcB46mYXPKIrost
40oL1VumPoyqg1hn8COSksjJoQ1Z7IYvTIzwQ8nGWO/vrqMRhNiZo1jm/FqaYEeu
aqWctRAw9LRZ1apLoZ7LaZd8/DGvZ0fRN49KrGQ70iazdRdvm20wcZj6ZCUlbyBO
5KudhOgFGKSslgV04dJ9sSLIwdFuZedXP+tmcWUWRmQ15IAHDH/a9Y4mELsLAdEI
sotKp0SH+wYr7NCci9nQEvH4+0caUzS2tjOJ32C2UUy2LXeKHZXmAIrVqeMdHk+p
84tJflhg5dZ7YYAg3YKM6TpiLavUwqPpzPiHUMLnwHTjYeLQO2t6RlvxGJ+gI0ly
JfQBIPzKwwhDxWRpxNUeUAr4GTuJzGNn6jAbEEZd9FOOXYwuJrirqgdbeS2C5BMe
eLNmEpWEXEbO27EK2PNR4DzNF13L6/MbAx/INwf3kpulqAVuclrqCuj2aVWOS4I+
sp0UXTfBlvSoo5YI0924qI4x76gZOXyaCMxBQ4yz8fMMq8+3v6ly9alJM8p8WWUz
Y7w6gSCj6Abv2+BVRPVtsDckUjGIZRmrFS/bK0tOd42CMGwesI2TQxPYwPuqyrKp
f9b2XOTYj6IGs82UYm7a+B9cCzST4M1sLnnDjOz2LrKLjE5blkDDyzErymEctk/1
dY/Vwi2f+g7j92eSenlWcqWmzvXgfxg+FjQ71W087oOlQxXe/A+yMsitFZ3i7WSN
lWXa4NXq2GGWju3L6aEdaXtYPLeaOHVEwwL6LtPxfN/EtgAKOLGjvHdsvm1BYed7
2K8AV1tseeg/KYGjjM77LzyDGGRWbc97s658GjisWtKAWCK/MwH9r8OCv69kHKrB
6mj3zGWKDZ4gAf/4zglJE18m5Gcufp09J6g7/OcOH+oPh+7m9F9WhLHsqEHQOktu
78PzhuNraoRwk1N96vGhmJ85HdeP8lWTnsfycTLHP9j0RSF0sxmtZT9xxY4sEZdD
qzVAEuVPsSiZl6itDRRAngAnK5T+oWJXtEO9O0D3AYb+Q2OMHuWuxMUUWML83Pb2
3PZhKE208X+44NMTQ/IjFRglYTQTwQI8KIRP5asAACumEucmRzV4qrbI3rdZqVWD
dioTt4mzJaK+8lwzvllusbW3fksDVZmKy/UV5t2pbxJVCcGikmwB5WEc8Ztsn+HL
Tf33XxES5dwsb9D+bgnvNaS3AqVg/8txveYZS+pLIykWwlhtIqkr4qjMnRIvX59w
02T6wr7zeij8P+0YhW8MQX0wDBdJh4CaKl9MJaAjQ2GsEedJoT9TRsr3qqCFdn3x
I7GUabUh6Gtoa+FpIDav6+xgUJ8wav+Da/zVQeHyGOJzX6WfpnHWKh1RxLb2SBBX
QXnHBx3HGW6AXXjTa6ymgnD5ppLhYGgJmH9emgLiRDyMRdI5kUvpTrVhxOro0JAc
KAnqSqnC6y/4UDUACX1RI9dMbWmw3++HYxBcBYovsf790P3t+HHmuExGhG4VJw2K
ma3O/m7/SH8XLH0CQntzKVtpDy/oKgBdxXXIRmEFGNAyDKHbKxjmFiX3JpStC3Ld
A0nCuoLIQkidwxDb4J27mZ7wv8Uu0WcvJBUxuGEzVyO+Pb7yuR+czjDyMsu2YZk3
lpEmGc6fBuPuWpmeSArqNs1/1BJOgqzbSil9MrBu0bqQF/CDx/xjaBsgXi28Tp63
6hnAhphr9vLy9VkHh1QV/w+TaR9o2y2aclH5REdcATfSgGWea/arghRDu7TKeBkb
40mF8i69+GW/EMDTQvjCPtcQhg1FFd3MnIdid/5IDNY33PBJDosw5xYa3x683quf
cGiBhuMbhIw7G9ACEqwbvFRbyRV+2ZP7h175uFfubghzFSEUmC64JPk2x8YOhaUP
lBoMsXrKW5s2tzhjgPSkFhBSnUU6jx40XSVsg36ipaQbG5nbWT+v6NoY4HWSEJkr
UWgptfVKwZlKNOcTjkfzfVyCk3RZuRsMMhCeTiErLV4lAxRIXc44nnEk+LBdvscz
irpAZsIyCDc+rTC9xdQmdNMLtWIX5/PaOWsD3/kl5hE0EXp8BUqzA5pfeIM0Qdql
g5uqOt7LDpgziNDC9+rYkctjr+Vx0U04M6oZrHYInW8qyqbI2UyM/nQDqRb1+o0N
kL3edU6gAfKW6XzMVFwNALXS/CEEUXOUjy/DbT+HZN30YUu9sK+Zs9AoCHZSQYqm
5B/CSI1cVZRhPVRN2XGMuxPbSEJcKQ69olICDAdWm//yYudgfq0Cbl+fVZ0S1+Vr
PTCaXx9JoqZby4/LdhUN0TsFhxV8xYPncQANmV2EqFJcHA/dXQFVJlsPv4mEUMUc
9qcMYg6nmQXku6MYztGlPR9+DIHs56+fixsY0/Pci9En3S2Izj+HzQ1dM+tSKiFz
pUlZB2B5aLVgCAX5aQHy5UGCYJ0cyRS7lCH9DvgX/cM3pi+Mj6RHMnMJi6UfpI7d
4dS13udTOu9LusukzhQSviFUCfSEL3t0B3v6+6Eiqu36aX8DRrZF4pfjc4XyLEmt
f2vV0Oh2WA1unX5Bu8To0edELbUfCbDQLYE5wEvZQ3dk2JC7dqAHWmR5B2xkdBpE
loPbxVyGTLVCq01vzccCvxrUOucPO5GxIYHSdUs6/glWMzJccnouUHpcQSq/WSAR
POs77MM3d2qNsU0XGRA3ieUzrcrEel5oaHTCddJWFHMpXoAfO3INdOsbKtVXk79L
kJnnQ18QE3MqAD9Zxk0bCa+UJegxyvp+J8YQ8FtrWYC+BK65anbg2LxdrDN6e0lh
lYqWb7UwyBpkDjOO9zW95irJXZK1ygLK9BOdtnafG9EVoHRnSpAVx34gKC7cWv/I
63/f3hJm1U9V+KtfA9ktYhJLIT6L5fmcp45ozO/2neVLohKOJFw2c4Xdw08OBwh7
G6tO3Krn2kLrBttBvkrdT1Oi6KKy9+qlriGmCw70xJXcDLda0/7ObZ6wtafkD3c2
tLsD278otjfehdkXVqSWhWULr81QVq7z/KCPiJuog+vE3ZTm+8ZGpGKNiOUt7z3V
zB5456pSkdlINhFRhBZ/TDIxx7aqI/roFjdhoBKqk7GUtI6WGSnMQGbU0lFZira8
56dd4wDeeJlo+1jwT2q3TXtF+iq7Nlxjdl08afHomhGpqhDc3lDiZRbIkvQO4q4e
ORrBYyqw/i1UP+QDVdCMTFb1Ny1iUL6flgPEBeiRT9a2ExZaN9Pj1zVhdLlDa4zF
7miSnE2FAtTN1W2QvS90q6WIKZYb+/yciQ88ooGC9iHMX9m3dkbHPEnW7wfl9VTJ
UfClMrw6ZfviVi16gawmZlj1RLYCqKEOf8fZzOXvYgtxFD2cxdjhz5K42qWfC8/N
XN98BMb7kvRVuBluITvQJp1aYpnT0nzHfQj3vrddUdo5cCEdXGeeLnaTi/2vH16+
cb+cA4+qGk21i78/n+cuddQVmXGvXxOjvk4DhT3Xza2kqi8WN6sThKnHz9Kgyyfp
h60DEL/ubQNNSwdgiDl2bSGTko0qEjwW0EhcDB5LfqE9Fq7c3g+sCrtLZAe3HEby
bPI8m6dvuVgGspn0X+aKwKAqk7i6yrFXSX70zQa5zw2WVDswR2/9dcliTLrENmLf
EwyKg42iLN3GhM+WBClqjuNowQnMo/e+x01k2SpZQPyBR76/xCXCG3ZdAGud75kp
2AC+zvNQdMXXSaIOKofFIUIdhDRVgF650UsgvSbBwpdfttf7MRDvSWqJP0Le5+KQ
TzlmC7K6gNdxdTfsaUcajeLWHCc1i5doq4FlDb+DiYScE377+6sYUDCaFF4NH1Fx
tYJS6KHOaIYS9yYOl09/rDwVcDcc8gG6vJYuApTn5nUts68J0IhM+KgByZRU/hLr
OU0wRzPcn0wE2k6Jpo0a2KMtffBwXUQm7eeL6gcZPPC+YowH7YgWEfEqxsZVLVwq
wZscjOh1BHM6EHnAr5k6n8S74TBzZAj/mSoNJxw+QNUkO2E172nr9OsFOCBjjrYu
KZBwBiPcgwYcAXy1VT1aPtJytzvzqlP98lddIbOthnm5cCA86f72rHSbRAIBblJB
tZR8uTEUufZvvBUTMITzH/dNKTILF3dGo25c5bAKrq8lnER/Lb05MqsIHanYpYwo
FQbVBe8cX06RMG2M3dnXn2PPeehC46NbLss0f4NFYHEcNAapt841ctSz/1YVl0eo
+soSMET+vxydwP40eXVl54ZeUhrxPiWeSglvTQE04wFkDlV+c9EX9QYChBd++WxU
b1F0fNPXmkOyWmCnfYSsGV5tLpUf2T3aeJW6CHVWAgqxQa+sgBohh4DTV2NQXbmW
FL7BmAM4pcoojkwsQaPHePsHdwcoLi1IQkucZ1wX27CQ0lPpDKUWCRSp9mqXyMfA
3h2s1Ah5tdUpBbruYYJRUJ8kLDXfxrRMc3MM6qgcSt6Dg3/Xpc4+u7hDjkoMhQhw
4ugyoMuM3wXCP9/hVoCkO+LrRsFPuXqDrxrhvIzHI2UKce2PUdIRcyfYOdlehk3S
/1SZVe8Acn9EdRojSB54rMWr9gaIjfHhITHoZPAUOyhv/O6N9M6gEQvJnEwyf7P7
MGMw2NdBq0+ScrjD0k1lE4LrgcYo9f9WeGTUpWMYQIedjMlndI7iFqSd6DWr2CUi
Im7A/H1lOE2/bwRtXGOrIFaKvO3pMFBYz8qbWQ0d9WvsEcPj6JdlPe54GiUW4P8b
bkblCVZ6bMqk1l/bZGW1AeWsXYcpA5cmLHq62lORl20YgxVQo359LlYCBvNCIwp8
tZGMMFX4eWj/s9EeERMhygk5gvesTcI6swjEXyDsIpSrdbJnMLKYKnoVOqYg+FaV
ezqTzuFyTCRdyILFlSNiZqGs4CDDYDotuqQHD2fJ6J9f0LZRvd+nZA3Q8Dzns01o
ZOV5fKX1LpKqRHwbDvDkNq1UBtp3VRYXI0JJzr7Di1Vlzx+ApM6+viL99axEVzhJ
5JerxIN5mhgZCZhQeMDpT1J6Bm2r3k4mI2028Z/tvb8YRnQ04Ua7fbnho20MxDom
H1O56GOlZSkf7dbI77eaU+ZlG8Rr6uIhd0POCYJRqbQuV43LPc4bSkwtbHZ6KgG4
mJpYoy/6nrv/sE2QWmeVaAn/8o3ZyW3CxxVRveutRZqYiMu3K6wSDY0+WywyfR8c
/RVlPbRydj4XSaf/CGtBNP0cvEPo+Qh3sTTJ809pxY1g3dnhrZH1EP2u9oX+4K/0
PhWEWOnoTX8LSjDBXUjhIRsz9fgL12km4nam49634K2Iw9YcfPkGvtmO0q2qMGXH
vNg7J9bRWrUg84sCZKyY4OJN9keS6wYoBXd911qc5PXV4qXUobA3f9iVIhP+9ett
AA+EvxO1SblgPS72dfTmAu6fhdDNMLSHMwEghCDgnZJWO0d8Yw9xSj6cZGLopLNb
tVieOhwcThaGsW2MK5LYK4h+HT1FPiyZiR5rMhCrJeYSVlKqrQaQgBkfllL5EpL9
oi82qMkTrTCNBTtzKR1gVTIDpZfzRSItzBR2fRoHmEK+aDjO/7izs8oAPCwYjxna
+NLxdUZ+iXp5Pv4x+m6bfcgtPmdBnQx7ohI4scQecLX/k4fMUdq423P+QkKOZ2KP
PI+d7xMwIusXiWLQnfepJQIefHmHyLXwyk0i5F5ytWRHnAGUBdc6YhpR6NL24iC0
M/HwtnAmfgLSuehaNkamZ51H8D8V1gCs8HC3ajkbvmiyzrnUGqZtgAXPpqTEiOLA
P7Zr4rS5OYNg/XlHaefISVLtQcS1Y+XceQUFgFYORL9Q8Sajt3I5a+KvvcKgTS/P
kWNdXsd4fGuTuyOfPwCcrxOzug0DqtMjaeKj/a5bmhzZkZBDhRcZQ1Au7gDc7DSH
g5eST60Mu0gLb3BjLOJDzeUzW1rICs9sbBRQ4zDCFAy4LP6iiVD6HYQikEyPg8bn
Vd+7gCrftN3ox6yK/65v1JueTgFeixjX+/LUl4cpCs7vomgO9wwHR/P7cOkO6xIB
I10L5oGPsrnK1156pKDrryrWrV4jxQ+fBuUUuD106sbDUn9gm5t0L/cB449aA1O3
JLwr/MO4+qdyEzi71UuUFwdOscLOvOt/MnhL/TklRe1u5t9QZ/wbEuji2XklSRDy
Syd5UCN/OO1qXwOzJJ+CTPQwL+g6XO+A1N/NOi5yNOc1EnCIZcX3Lej9KXFn6OIr
xgPzGhGgwEfbmhPmDEAmAyZ5+d/yyAG2QwtHxOMz24LqteqEL8d3zI9TXZlLayTc
eD/2BwoozjwRQIp4xk83OQdYFy3JgieADBFrjwqcyv41q+Pg9NuLMHR7UW9tHmi4
xmeVsB+ldt2MyMzOnsuw0jjI30eOxropFaMlsVeT8NJs/mVhmwJKZpU3+//ZIt0V
KvEHTCBaWuRwkoBCWKrSo8/BcBEVY194PlgOKfBpHGz43zK3MAV4SEJOsGJj6TaF
Cwf9P7INcZMTut8395q2Xl3Zw5LXJg2QOj2EI/KexUaZ8ar1Qc0e5iZsH/pXX3JG
0342KsBKHGryFcL7OGrb66FgGCpv+6+9jmmSAJPYY1nUjX0/Xl3nLfi93DUzuXDb
j43aelFuBS1Cg1bzIv7jh2Tko7Zg/r8Ny5mYtjrOd4GoK+8xJVzUVxT7VptVIrZX
v9/8uPlikxjjto4pdghpglXYs5zPTjo58EfdJ9W0VxTMyv6p1uwLiGz/SvKRHqAu
1iPrWb8zwmqh2m9fmseGLms8ZtAH53ltVIktOrzE8utFykjtXdj3y2NhSaGFxhb0
rCEkGXoa0kbt/DHFv4WljkqoT6KhaglFI7lrCMF1FwvFwzai6EXUSflkUxZEafub
s+4lpsgO3XCQG+WOHphIK+EE/8RhbB8eNcE4jeqMWEsuFNDU0IKJC/eEgNXifV+V
ZhTEvKGywpxSUq5f1J0AxMxgprWmndyLzk4VKe09Z/4CE7NDvkq0xQD5Ru0oPvi+
akk8JBfJECH6ol5j+3uaYkGwPTJCyZlhpvFmTv6I183uziyl48YSuko6O+RcF8LA
+Kh62L2R1tmlMbhZZbsOnsaSiKDgFQGss7ByW9/JUfY4hlMztyQbikBNyMS+nodE
d5NBBgq0wlx+DZULSVBwqYwgbKCwXjt1NW5vBIRms+2tZKNJhFOlLfMHoIvA7luA
o6Ewyz/TR5TsS680sGWWxub+KA0YiVZ5m8+ZLig2n0+Yuiwi2Xo0Q8Q/M/xWlKAY
+oHyR6STRkmryIL9W8NtzJ6Dmz7xh8a+Pl3Xf0N55ZJLdNO5TQsrcGnAe/fSgDCD
WSiL6mVrHx+fYGF033LJN49EpbJsBBHWZf8tk6p05kskRU6xk8LyX0VL9+6DUQyh
7xLRsFz0Z3nNOxl/FkKmu7LRQkOFKRaDmtnhzjIQquQq6Wog+69NVXbOI4ILjp8B
7o6d1/FzDA0BYmjCJZ88KYLkF3+Q8EEjjCuPD7QRlcSmxVyvQ/gCzWwzjhlgEadA
GKAXZV+Mp8tCnc/tTiiIg5t8WYHh39Qum/DZZEBC+m7ckfN5LdamJyDDhsIHYzdT
SX1fgG3dHoRtZrFtLxojomR70V6Ug1nAcrbmmZniBOD9BcSyqtVefL6dblo9nXLV
mNrk3adRckAIWhFwVRneoP4e8Gn9q5LeJj6w2xVVtIlDaTSCurUfhzQvT3aTqxeh
K7utantIyHJr1pXpGlBvzkkXjUNF4MW+0fZ7g2HaL9X1BB0n5DrM/DxR9lksA/fm
O0wd0XCO59CaZ4NCIimQGwaknC80gfXbhf2B6PMxbJbPM3pVSGWbdyoHTj2U39oy
8OFEOC7AX/hBp4Kjr/GCrGQ324JJqcE7vT2qpQ1y5lUJZ/lzpYSE5iL4sB5hGfZc
yK1uffieX/mVlpAWE7RrhR4y+SZ8Botw52iV2xCQt9zhMeN0g0aXu2NifDquL04L
Jz00iD3csxHqjPLr6D6Ae8pQkyaSJPGlHvE0rW0yRxfcSyB6fESZ+xKIdFjv1QXt
3x1O6xJZrp5+Y4TMr/Ch4ICk8IaohLOjYOM35UqT86xCJLg7UlojjH/iRHVDRvnX
aZL/2/ouBmeRWT8yj9xjlf5qwyfVSfhxQe7vHaiB8r0IWvpRH7/pReNIN27vY+eJ
Z5U6ndXQ34Hw710u+vByfFQW+SP/svAGYO/r3oZXe+Lm5cMoWCxEJiNytK++ZqDC
9O0qsgotdg7G7Q3k02Bb2V8j8tiv0DAnbFmQlGgu+J4K1EDGsz2TPb9ZD+2eK1wF
M1CFYrBYiPjfmA8Bq5E/oN4LjOWxiLTF9SIDW99cZypfa0y8TVV31gTlNEeu1YIJ
iFr94Eje+r6vqcbVMiS6WKT2ZX+b1dTotB+I5SkczLZF67SbjAY45jUb8PuzvsqH
sS4VF459n0vfa+aPE1Km/b86yJfjxIG2zvqbQVlfWRcdLLuEYyyneQhLTt5HevVJ
qqu8KHEjVB2LThaVG8l+7LtQ0dTpZvd3gY3831i2OVOGsRPlMTvEZNTyDeNzvtRJ
r2mNVuKKQ1kdEp9gJM0jk4RzePtSqFKR9bkVDwbcSZ2f29SgIMEdR9i9LtlDb+zM
8NOD/9fbVmeX/qhtdoVmaHClaUxBSi4sgmME77QSfwC1KTbi/U4uNMKkiZayiPN8
YLPsLIX1GI/eXs+4kJ4DtGaTfhRfhVsXjbRc14u9EYhm9SDWCu/aVJTTHay9oSni
Txaw3bPAu10u7zs2dMIYyV0ggLrODjs6GgjeYnU9kV931hMn2n6HATuji7myHgsR
wK7MYHBWQeAwiSW3RuczezWIFryTi3TEJpazEo4TkukTD/0mPjh2wFYvxh6RJGzl
HoESeKNzm5hBFhCPBlxXLp9X8d5akzp6TkwzZ0AoSX5nXpqCKyS4wJmNbjoQfmkK
9QggSOrzTSwFLZo3pW8YmcF2o1KsPrMm7dzcd8t0+do/GgNm3NPY9yYDxFV+gzn6
R600f3b52KlLblEC/EwDB8N87cZJwHpnmeMzMeGJTHeCUlFY2uqPxIQAUskV/ugv
kr1KcrVtdgFWW6shPDIgZJOAJqB/zjvYWW4EzlzSQEpXUg/LqJ8ygDhREiLAqG2P
Be6AKJOS8pm+BzBnBSSw+GXjTyu57M2oTrlhmQkHY+CpONMRqYOSvn3D0qiGkmV4
TW6ru0XqvZhlkcMFtMLBeSInd5gZi0Okr91xnGwO8T9NEc/94e5j8tvNRgPFGyHY
/9LAFn9q9JS6zCX0DIe4v9SdnyPt+0p6/bPpZX9CGQS5nDruLZJMxcpFb2t7VenV
D18pG0+sdRKD8FBC4FpkRRT94x3VEndmgdoL6Vdef1wYObU7sFRsfoMolE9xXx31
RGJK6aetGA1tYnFxbwSh+KyyA0Y+2J8jwW/uiZynGSIvgzxsn4hwWsJiwI3Q153Z
O4pA2uQqzkVrv13hUbTlX1SlfD8U7UATRSHaWNbXIW6fIlQVU5lm9Bgsa8CCSlgW
W8s+mG9r0XcFupV0QJCPHfizvhgbsHKTPLV1Ba4s5l4kyLPJlzgO7z+Qtae9kti8
spTP14xVhhvslokLPVJP8KZs/gF+ykDzcWtKlBTe4Uo+AMpgGzx/n/eKlyXvrJEy
bQqcZ/pKYXAkoygWdI2CtwnyfG+XgLsg7g8WcAeBVkZOeTIuBEviL3j7ZNgOVuNO
Buhe0ml1unHKAvwRXbJ/XP9NjVuVWtybUDrqlf3OJ8gbdT/x9vO8JwvOjsqMpLL6
HinRusACUmKIFlSkPqxxVaHjT8XD0K60twQAnBSJBn0Nf2jV2Y6VtWzyeRpqKbO5
+P0wBgS1i2eiKx1D/EQJhkRLq4sklgKj9BKBRBWgWWhpQRdKRXbGgd6VZA1ix7LH
eOmto1KrXzOpW0rIlFqDcAVCQ4yxBi/zPgyjMcjSAcE4aks+aW0XyaQMUvlHCsMg
+carpY/JWbRq9vKXDhR3zCtcL4luO7nIEFfk8nPvEQMdrK/aGP5jWTZj0tdcHPJU
js1d/SNsq2IJVkXvr3uTLYQ4/PVALsEhgAr2w6Td6UVZ/a8lmjNpp0YgY7XryedD
aDI7L9vztkh6XbUVA2xHpV+MJHFN9jmU4ywVYLK662E7bOGlRNN/QX6P5r35GIYG
cZlnmziEiHVGZHBUBSKrvrMT3COXZ0vrZTWgUA8bMscjzlGO9TLMNp5CHueFW+6N
t/P6ig2m83F7/csTW9wz5pOB9e5vH150YZwLrrlkC7WYon+6re4pULZL9LYUr12S
beFn2aOEx7Uv7q2dOC2JrdMmDVpPj0UrsKTSR6Mg8DEMticULgJ/yNuLPraVUK3f
bYKsJe/C5giDLLfYI0OZGIrdZ8LWfWbWjxJBs99JQTfAoOBVQTWIcAxFaLoECRC8
+2HjQYozuznmH5CkAbgkg7CSmX3y9wh3IOTyAAiiAGT3HJpuh8VGj1S3SF0TYL49
t0KhzB+s8pf2MRoOgOA5ubJjQ7WCReXB3Wr6ure18pLUcLsmZ23FRj1kkzBw6yox
dY82paYD2OZZk4uIKzsWp3sCfgy5fM5ttdgarB0tqJ5vW75akeRomDKhQTK+a18j
bCsZPac+EgSGfV0hFtrwGc2YwOZNbOqxNntm1FTD+9OMY1Js9Lp3CUULAQXtn1VI
fh2rFfoZONfYFc2Oof6tI0Ik8EQ1WFxZynE+651/imy5p1x5sRFZjLn9ZnRroFGs
YLDCvNMMC/xg4xUEKcgnpr2GwH3nQW0y6s3TbmvE7HcG2uDzJMAPLqpMSGjUvPKb
IQQFd4zF3+MAh8DJuiTyVNqJxNOveDiqK1YQ8oWsW0Aq+HMlAijREVl1sJUhlP+K
af3tLsDGzLQnqadMpgE8OyNFgx5t/kXShaYZqE3BRU2jGm7RbXubc8i56BFGzcIj
qZDgJvxmbnU6Yc0c1rarCJPZBZU8jRZJKtJKg611STJXN0+qvVyyUiPq0DAocIW+
71KBXjdTL/jDCbynyVa89XVrOvAYqlu6SPa+NKVWlCNK/RP+xGb/+IIllzv47xGQ
0Jchizwec4SDGEbz1RUxVr+dQW0Q3HFg+0DZUowz1xKcakTdTkvfeXvtmKs2/ifG
RK+CvYF1gQVCSs3H9E4ShS4wYCjkHykQQoFh4XN6NsvJT8DF8ikgS8f86TXiwuUS
gbIvRcOC8jtukQKlU4rgNoF8s6H45iGyB2s7bHUgSdsFvb+VtHL8IMoT/UmA6ufk
9aLM51i/mBWSDlYAzKlXHTMMnIhHgO49YFm2Bxrc9Yb9yT4eyXTcku4K44Ou1dGZ
Ug8Q22wCFIzoDmGPd+Zs4GiE6921DtE3TyIYN2YZT7Y+KXXEaqJmaUPHkSvicXgk
cK9AArmYTFx8+TWLHoNgm4Y1OzQRQJsowlqySsRPDxRj23Li+45Ez9KkDTn5t+oj
YLj/n5kgQ/Wah7wj5E8saUCTPLuq+RbefwtmPhGqP4ZvSNA6jSG3Qk8LQOL6jCWm
0b6sLOngGTiQNaXYPY+FT/fiJeSLwUZxCAm8zJB9fWorqNd4O78Twh3LiTaBMD4V
fwNjQbHkJWupP4j1+BG/6kLjNPHCqE/02u4h+6daOcajLSROmRlaLhL18L6+Zd0P
l5kDm7XIqgBlAddiqqZ0jw20i347QgoA31me2bMOkv4Z1iJZf7bWOlftRDLAOtys
J/lsSIadXS6fehSMGukcH2tpvEcrKPNt+oBlKvbNi2NKiCaRBu84Uzvixy1pVZjc
rCfhGpBX1+LfyY6XjtqzHEqXhwwbiE1ySxNBQNLPljHDiljR90ijKL9xhyjkEX3N
CXvuyRtRRwvIOUFKh7S7wTZvnVgohAJzFGUCRnZ2ZF/j9zc3r/E0+4tzAhPYBrK7
AlhRd4m/gE4m7tkvjtkiwwYQb94YfGbx27pahjPEdd+mflWD/yxXQJ0vXYpRqgmZ
XrNlQ/36IahLKSFlsnj81VS1EWdReo/CEDtMFqjzpIbOMeVx96QfHi0KcN1lg77G
HHZXOueSju/g4Gs1f74PDHri1ooaPgnyw4Q763RCbXpZ3W/NfBfA5sOB7gDdJJo4
lB7bSwdY72lAm4dBCl6g3iHBCuA2Fw978KxdgiRq7MVzzVb0pYWpXEHNKCusXyVO
uqQjf+2KBMHVU8F8fK4XvroPWysEfbMlGWGjbw09rFyrD+yRaSmlezP/Dm5wJ32O
ZoLue/lb2yxgIXobb2csSqnOV062zvw+RNpDuXu0p5S8iFrAgeG4QF4sLnEVc9y/
Uud6ddZyTdQWUsTrrrGEtaQunyIhUB3dVKc4QyZfwcBI4NvyUJt7W4MiPdlxYVB/
MU3nWZEstwWOibNHQQzGeqe94vDThyiJEmvLQ3mZdymkODJriNgQOY0HFmhz7V6x
LplAyITyO3+NOG9g89fy104FuznYOV8NGu0U2DZpJ65yE0Ad1eLsE3cpGv5KushV
I63Mvqr9XX/hmyuQo2UH+7OuLNCBozpwf6iQZrsck5iaajixGYb3ywdduE1mFV0q
TDVTkWp9Doy5UqHqxbkmHaD66YxcOiGvjPCtXJLst90ghaGa3ki3G2eLfpcY852l
AgajJFE9+RvUAjiaVx3rrBMQ3BjF9J7rhdvVFp3sj13i88C2q9QyaLkl3cZMrAQq
Ir4ZuDluipE+wP/xTJJrPgGKStKNgTpo13ULV73oPaQ7NrkEDNe9hyX08MP/+aai
xJKjCp2m+nsGRIsy57hogrtDfHiCBbdM2sFsRFH1a+6oMOBfCdyoGyRbyu71BUKc
mSTIKIpSMoAJJG7MKFMqOHAVURQRaHn8igWAUIiMUGXrHWht7c7XKw0WlrV3REYT
d/h9exDNtuyncgpWCfMbzC1Z19+vKmc4ihYMtcez5xTKylLmN3Me6prfyZu/yb0x
2ETrt7CkqcpteT8/E71SZU+GLdxWo3+ZgE63/Y70OqD7W1fKZ+JlB905GnqXbFas
OrzMm+hGcDK1shKoy2pmEf1DO4lew83Xc+dxaaZNlwEDWYtgvlnhNVxv/SL38lAp
ramOrLmMJRF2Kt5S2pi5t3YYfldS0P5S/pM63avnJZwt4V7BYLMXXcC29SucJYoL
5ESdmxK2ytVVoRjpgG1EVYnfgUKgWU6lXNbWvptcIA/2tJE8qvh1bxZKupnakQK3
bJtNNkZl7nXwv39iSAaLzqVnoljerH5uXw0dPkOb7A6RsLEKYwdqX3b4UCsxmhpQ
P3VjC9boPpA6uaI4AKvfJvGVPWH1iyKFE9VttWVeoQEDzN3NWkPNXJMhZDew+cqd
aQ5+w2Yn6Kxa87zRZy+bHpddZlSDgTMMUQ2JXwsTUtxJlmI/ZR6NH0/U+OMQPohV
dAG2Zb1HdHUgzJA7IVxU4la7YInCG/dDznTjufmGQ/KyIjctS9P0H+F3Bu9NS6/X
AevuxlNIRHXJYn6fLZGIBw7BTHN32PrQYY4q6tJoKPXgNkQky7Hynj49U+1zGKoA
+VU47NRZyGdzt3hOtG6lDkqGwq+AIWMzR3PMk7RvWZhDd1UIWzWIdG9RoxBi8++L
Ve/hhCmRuQ/RKhGl3PYdLVvHJANga5It5/Ib6j5SHyLULYsnnWVx3VWVAZrj32M6
OSfg4S597YDAJXecFtMzYoFDsaaWi5f5pymKc9w3TubyxaFjyXdxcVzDfYPKoRUM
tLXJ831z1tPdFX0LVL0LP/qJNsYoUEvRvbFbxxefRUjzNkSGdi8sf+zbddFJ958p
LNxgZOb+wypJziMEIQYvR7cFGLeYE55qDDTYH5uIj3u3Zn/sCXm1/4cxViX6vNs1
Pbxj0Nxr1RaDwMyO1yDgQZfzUz74XAAGMjgNGvJ8g5DGJVOE2inF/HeKRaXxSBP+
f7+BF2Rs7ClH1AlIcwIVxTKfKc4SsW3ehJAkJ2gfEuudDsjvaxGq3ZQ6UjpLp6i4
9pRMJFLtmRzkCl2HkO/m2cznLeT7rf6g68/k+tnErTNWlRhyhsdGnf+w4IVrN2xi
KsN9HGZeduRwX55EsOcPDlDC1yWdrq52v/0tnPiqx79Y70E/Lp4IP+oAWdwR8/YU
JghWvF8pQYPApWkTYpt1mn190mPvmE+4pToNmKit+eE0eNBLGe0/6N5l9IQbwLXM
e8Dle0HCCLspCUhTU905L6shSaTKocsr/g3sxQIBgEj4ddfSBFcRI/PRRiH5SbII
d4ZQFtrLTozuoPTcFIKjQpvnqicXHWRlzWCvarODrWmW4hSQg/KpRuD6N4Qzljtk
gHB1GpSJv3jKg6Uc0EBmohH2ieGfGNY4DxUoBnPKmfsYXjUvK26MVh8ydvtXRnFB
46NJbb4xXLpPZjusyaSehrllZalTSBTsB74Tk9zwdcdFHVxjd2+R4RU+wEPPISp9
H+6rh3TShc3b9tCU+HsuONO01jJMmv3KX+yUcMKF/3FQtiDQwUOekJpltgY5uoyE
GaPJkAAEHyWPX+bK3g7+BZkOzkqyrK/If/1flDUpFMvoVu8U7c3dNvppN4Hk4/NN
hhcKPZo+PWsdX631DOLrJ4iyCvW4KyJdovHvBfLODBqUd/7MCm9Ypa9WjXUlrRp4
xhJc3r14GapRcqVyUcnB1y6dGrpGry6SA5Wiol/xBKM5z61WD3naLo0kCmk7sXQU
Pfv4FdClLKPN00gJWSDZF8HWCRIFq05RNUlE3Y49dhVvhjaWGVeFWOP1EF6vy42h
FlTHl5s/zZ8r1W7ujukB9DNSeFTQt8bOVgvJy99oexecgzcQER8MXv7zl5pzrNNE
1M0LCtGDimzmusOfLORN3DxI0nEGUn6+eQ+8Di3lV2YNs5G2EXXiZr8v5p+8xmCp
eDIs/bIKE8sqjftzRXimgwGyX5/V3o0SojsgehYNPoup/Ie6mBaKd88f7YANLxnl
rammx/stbniG+y01xvAZLqku4dWEaGag0noZWdYlpWIgnIouvoGWvh5YCqy+76WI
qe0kkibdIAltbtme2RVpiug4wWeNWoJQ1Y+5+/MQRDctr24Ion2polLs0bqvsTiw
d/uEjCaMcgTSXC0jAgzHX7rBaHw2xcOUk0ZOAkKb8DG0YAGQm5WR/5y7/7U9oCbz
CRC5XvjUbpdXlj4Mzx8jrlrW5EQoGXZRy/9xhSveDLMxFU0PhWFjvAGz5dx3UEA1
wW9XDw8+foDtpB6YptfvQM5qyGIuHqPjrt3VNMggNYQEJfTVC7WcGiI6aI5Zv7BK
KhfRAayPvoV65f/3W59Bjw6l7xtZJ71dedAFDYwRKEYBhEeU9jNkYiA3V5AlryfG
610DpsNJb4CaUUrcepzu+orODojfV/x+mXDMOV0YMJtLXL56Fah1Tq+mHXYidfMZ
dyXn3tHo2NWHkgmLjbE8sfpay9UmIFK5SmCAhMehaRpRMtxh2uC3UMX2ujc8/U3H
uOHE7NIGdLGsaoySoYrKHJ5UmJSXU3I/pFKLsJHj+iG9/vtiHK5ywuGLOUFNSrKA
71WwF/0s4f4XPedoCSvZxcYwF6OK+1MAcutDDQ3IVyJDkRGwnMXJpwf91RyiSR/I
1ILzPOQiyqqGDtpLtW2SNQYKdKOFE2p3ZdqyQuDxNk/Fq0xPoo/Zddh3uThaWZKo
WZc9zeP14qku75Lr70qchvWnyYmMWgBGM3LQYRytp3rl75s0mkDE3cOLI9fl3FG6
k3Hk3mYe+h+sRwiLfnO8k+sXQ10URkwCMmd6ThiyNQIz8Yw/wbl8lG3OKfAZ+DJl
SxQUigY80S4vEx1nd7FRaigQWloGyTbX9GtM2CsWypvL+zieFDatjCaafC95UHvR
f08ki/h40ZmPo2VckQVv1+Uj5Ok2DmGZX7NvfQ9n+63a3OvwJUgQSkjmpWMk8qyZ
mUsIxhhBnHw0rqZyY7vMjWK/suh7IyjDdruS5ZQa9NcFonRh+PLwRCHeLHquXoVz
UV4h4iKMjHn/uxU8o9ChpQKgKtmmCr97flATUYm5Ilyc6LYxW764jX/6ATx36eZ4
P7DV6VHwkSGhRVNccy1MzJK44ySji8sdy3LkZzUyWQR3l8cscCkrVga9uv4MW0J+
2pElz4fwUkZUHVh6xbtgpkHvAkOWdQuDWN6R+snS2vuhA0UAe2PuABULUdHx4AZ6
H3EqQE0IJvpYzuvENfjrgTnS5ixzDYlXCA4DjJMBa46jmrxs2bjNcsGo5pZmmWZi
t4FGV+2j79oxMzKm2lMTluly8jB9ldWrAUmb4q4/ZZjm1rPHjEXsrAj1vJ9ACziP
XtK+gvtPKTWaLXryUjjZzXBYBjHe6dBFB3x9oFQyISmdfKo1EIimawf7W7WtL0kc
vUzNxe3arC3kYkodWC5s3UNsnsMRiWYz28NTkbtOI5pcf0mXrTm5W/tnfm+HJG5V
5o3PGmjjWom3t8xgr8XzQtaS9XhTYK3kMsu5fg6AQfPSBQW92+2HftFsGtSIPhCJ
+V56nVkBEiLYvI8oY+4xHz5XPiJ7Q62g4UVytLMljK62cyeNPLxJZ0Dlz3t3m0TD
o+HbMhdJoKovUCelwDHnSFoKpch2PW2ncMoTKmXPxXsbTarloxHvgjg/hDQGt9a4
0Mw15HgtgXc3STjU4xeRnB7hAqt38FbiwJnANILR6tjzM4r6tegoGBW2FCrGC0xW
uP61+2mpPWaCxRXWsyg+rp/RZUJgP+tQZ4bWMVFx3MmrGCsyhsAKmADtarDhMIyW
d5euF/izNzTQF7BRmz8IUKtszqHx8cLDru68P97958tb7+adQThdQoRS/9sg5bYS
UuxZl2HeiKGgqt6qhFdg586SNnsX3+Hww8rhsiu/MrgFy8993Tv3Wz9KoEj/h342
BhrVGZt+dzJG45GjuJJSHoXju5hTdcUJgyBflAl8XdfyzoXLhxUvL3IVs7xWJIRY
W6ygm684RfrJ3iTCXaTMwRdXqRlcu9TifrSmH7nCj9njexnOLCWlpoQJ+0mDQ24w
cmog80bGYRLCdgKd2u/kDEVgPob/AjJ/tpHhBdDp86MbekrZg/vYVDwT2Ky0pVNd
qw2X5SIm/VXMf3ebLFZeqeXCIbTqE4mf/wIjxlFRqWAyuWFN4braQ+wt0jW3AkwJ
AtTBqQKIZWbbwaSS1+HztuTjqcW01N0HD6RjtUvWtL9K1kDFiQ371kWVmv7x9nqJ
IHizgjAIIO2uyFaAq/WBXxRysCvkRU1DQDSGCccGgH603d0dgnh9E2nNE/NNu3RW
VpHjBXZaXabK4GszdlDnUs041qIlQqYg+sTGyrCJneqWpcUY1/kTTcDDO2TPec0N
X+kwsISwPbCikxasVJZ0MPRBcP80v4ClrMAC4ULJJeCsQAPhtvmWSuIkSjrCujEg
9cIHlXE2b+8D0+pcndJkeTOUVj9Z3+TbOUZG5VuExGWVVqWJWN/t1/5cPJBI4Z7w
Y8uEQglqv2F/wBnVplqXn5LWm2N+ot4+vigspFvI8I18dbC8mvL12Urm82YP7neM
w68OhIqj9+G+I+GQ9ma0O+6CabcUlVt5j5SvEHusi4MF/5JTHuBAxMwT/i42KLjz
koLRbgoQLr5ubdCGbW/wtFrtrlroG1E9n3BCMDI4Wz3ZPppWxmvqYmZMkvNHizVM
XwKWzY2inG1R2Ft6Z6BlaBAJ4EYjKUEdPgppc9yH/hdOZ2FA8sSGAXR7P1f85Uro
bqk/C3P5VfKpMgEo3oM7Iul1+XeOrLiKJUHGSfxzJhqwHGDPMTOVljDWzFeZmzr6
yvLqBcoJlJKHBE6F7iZcDOJRSEVI3f630znsXFDw40+hSeJTNf1sHjuiC0IzWSy8
ImK8Ryp/bZPFjelvrAHVEqLPywJvSsiH1Q3IEjMFGRl53wmNks/J4I5qB9vKAwMb
jYyrO1cYP+TgTVhz+T/LtbnxlbzeaWbjqXCMjqnWP3PBEOiHleWXDMuxfLfY61m+
lNIdO4zbN7Uq0VkUw2tfaCNJFurDiJLZzdAdAKS3r/3fGvBOjX/XT7tPxmQ6Yg6Q
O7hQxvUZnGEP40zELs4QOD9CBfolGtWtAj/R3s5fpRmlgR69IKnShq047acDoc9n
Q71je9gPHkFMFt2g/bK7/a20ZkdqyOyArXG34aciUTKky8bQtu3SJWc6a4/aPeiM
jzq3vwjo4HsCKefC13dPIE0JbWlrE+E4mVuaEWEm8mBHEZuEzaQ/NNUaSPPyEdMb
D2fdW/0FhCQtAbZNAmhTv6JOwD3VV9BGlPYa42adkhqAPeocaEml0sXda3RKZoFQ
lxLcWuDYUXeh+icURrn9yabXaMOBPbq6Mhyb9Lc71nyWUCADYbJi57WdML513T3P
5sWvmfV//Yr/Wqt0JWs+qyFmJdFLZZi0lPZka4gKnYNrtqse+qkEt5nRgLdREG+k
P+1CR7rMrEGtAHHMwzKMWLCgSNQtOPgtfUQ4Wl8Bl0VSCSBuhsLi8yCntjQyrrrp
c27x3zYKxHltwutPQf+3FBKU6PHPf5LpOzVrCmDMG1fuP9L5OVZtu3nhiWTxfyhu
8Ubj2hS9Hgql432VtgQWnlENo+/sViMoMfi1b89UCFf1GYnhgVrJbbvpW4s123Ud
HuxXBL3DmYXYL/hPQLCvp9xvo5y/1H5A1l4LLaswqJKQAYRw8/RStUdB4YdhEEFG
KV43+oOZuex3bKSwd43ThmuLlNmVhIrdFubjXyR/5cWfeU7PO7bFZ6fBMr4Vchy3
Pv8/+NtEvUJBVVPo1NW1Q/d8sUJYUrcZcB4K3VjKklNdxbsTD4D//j4akZPT5jmW
ElzidMRmK2px1b1DskRlMx/7MJuNbmFgKJKGr/G6cO0ns+LMYjY79z0VSJnmGEli
QBWcv94ap0zEOQ3G1f674SbfuN8d4FWZwlAbmG7ntC4/emYZG5JZ+4eeMh5RjDG2
LPzXhk0Ce+N5VjmE6foKCJx49lsa0UidMhX/b6mnSiLdVm+jD5Rut78Z2xfjpMTE
TpxZCzkKNrTPexOMUu6Rr6xSPzMksUOZP/2cmaAVJfZtlV0P2bpZ0z7qn3ymzKfR
Ef5ibvNVz1sahPI9C8F/Y4EOQ+lo6C9MjNUGoqVcRzFr6x/NXtY00LBeG6vf0gU6
9YdT/PCsYas5KsuMGybzNCdSUqd9bmqed3u3sAhrrylgkGdUGAu5qzxGUQKxDoQK
VtLqUx/fP7U11K7V8SACbFXHpVrh5X1e2CK14OEMN8zMTlFMVYMJew5JTQjEyQUi
7+HSZ+3noeQJ5C6AC/SihFq6gFYFVP/NTRpg8x8CVVCzlih1lhGjw3D8SAfF7XOh
IJKlQNWzT/SSWzffhcSxaWOO6f5hSsKiAQ9nrPmLLkzJ5P9wQy8X844jdVJJtFZ0
yDJsXW8TW94DAQwD1130ULOnV0Q562JvKd5GTc8k2SIlPX0WRgBEK9VQ1W6/AeCM
jxe++7P+VF2hLnvLKsu26BxAj/z3q2Yz8x+tWX750R9DRQO+FW5SzGQ5GUzzt/ZC
WQsAfw7IIo0xMKmR4Kl42OrQvU5yQ+QkhOz0zEFmlSNbKYiGSM57xPBtSm2eX4JK
n1/FtOtxHUmWEKHvqBzc4FSVvCQHsTQ/wf0XnmzjF9xND8tEer+p5XqDnE0NCj3V
GPAr8/Sy70L9JWbOb9ILoVJgmzugSz8/kGMOs62Nt76u+VHgDUQLIYHibPga4Hck
HJs3EInORHCUKffozM3a0Df0mqJteMM+8vrxb2YwuD2DGhVCJzgaWutSVO0FEYTu
w3F4YP9N4yatw8xTbqq/q5dEVuE+FprHY1Zq1Igs3UYRO6SVrl3yMaLIdu3x1YpJ
NHp36trMzME826qZnKQApODJncC/h+9JSYmK4AvGoL6ML2jpvg0Gns3btm77kYmD
2OEko3YNWSbgalQgtpeJDrjM/8MaJfnSVbdS1Nu3GwC5lKnLmBPhcK45P0mTjy3P
0hGoqhTjQ0Hs2CbRIa5yin5VaxnEdVQ3XHmT13y6UNDd598YG7AlIs3ZL9gDiHH6
Kko/gbwpQm3E6OithAwkSGgEWJrCjNhFwtXeeZdvDfwi8ei/EgAvIZ6BNKIeS1WK
fGG5tytEwvRRDgWzIS8mF8V/psPzs8ztgeQG8RxvOHVdHOftRjl/YoTxkaf13lrw
IdN3Zz1lq1WhU+Vm/fTtN7FBK5CFrYjavILRL4bDQnrfILGtqtGL0Jcgse5cfPXM
48FsOoHU/wmA2UxD+4T+RZkcKVq/QulcSpmgw3pmQM00kY0wyBA7EuCHDR1D0Mex
b2S8Hnl6O7Cd2t0xtm+8az2x3QYy4z82b/q4kM91PzXFlMPElvQozDiQsSLRCv0r
Yxz6nDHM+FSXaJoX57I3IzcEsDbO0QSJ9/1Rw/NpX32P4Upz9qkGjzqNCekPjUKv
0tO1luUMO/pz9CU3UU3ZU0MP6pRbjKB+iPklc0fR1y3y8NPdLREwnJrIWs4B835r
Z3o376rh1tZkpC5gtsG4qentS2RsswhmKXYOKt/Q5XdvOIG/ABRpBjg8fvWmceJs
gRcoTocD6EHALn4MXoCmwA9jY7NckWsCweqXLlReEnXWndH7h9HKgA5eSR3aUy0D
OI/w2sbzAVm/2hY+BVDHAT39qVhvWli6HZTC2hfiaTTb+Z4Y2bT8OQ1j2+/JSn2h
eR1zs/YcRdoQCOuLU77lfJZ8F1ES+kjOAHjI2ETKfHh7vn2oqksDqgS7C//01G6n
ab1OWj13mEgAN5MdZq/AZpU8t6V7erKdsxoZH40p6drK3dlT2/D+0pOkQ3WZNok4
ZR0LMrKz9c07rGsn05x3XsRikdZBuM09Eq3lfe1n5tpqGSHdk2P3ceiJSQSOlZKT
B44stmX1hjCpr5SrQatukUnj8Osinc2YbZcu8FooKo9+Wgtf9+c9TiZUU5/3CMZK
2jTSFJV07EVMhXS6nKI1fhWj41xmcqwMdgRbvJzU2g6YHNKnDsAXVCNyG07M6WF+
0if2Hnjzg9jiL3o6+4ppFE+z4yFArXWhoWkdOkn93GfquUdGKAd9SvYQXvfBt1WL
cI7OoMP/UtiCbG+w9CBzlK2NWBbMH+xQKYdZUpXIDW6lxHyNG98LfFxyINX9E/M+
GBuXQugn2mTYk/FIxVqCnY38SyKR0m6MtN9Fht+c5g4TWGDe1mebGPOs5epZsBfy
eC4JhSt+a6e9sQmJ2LdAtMTq590Me9oHUPIA2fWmk35Cu2Isq/SF0M80ObErgUkU
a9kIzGPitsNrAjuU0OrpIiuAQJHwtjiHwLeRHWxmBtYiKTOY+AFMBgA+wx9U2Ioo
W367pkzLbNDJvXt2rhAL+fxtk7riQkt3fkVnbJRIXBabCxKZqblv6R6U22PCR+XJ
e1/IqndZuyl9JkSE6zd0rTOYS5D1zkrRwnfq+ky912LqBtQDAfe5uBsrju+9l8Bl
Y5fER8WpHEuszdptXSiRg5jI2VN2T8IvczuoLESNtCYQVenj2k/3UcDzjVD3Jb5U
bMIRTGjd8vBPDClL30K/jIWPf0ZbhwnmttEjFIEiBJLCgyKylkRgr1ZhtTBqtqdS
6qwMGt2LdFsthy8sQgUUuvi4Z+FKQOSWaVFFUcTkC5iOxypG96TR/ZbZ5Vnr01mo
GXlKzo0DbJ4msl0VSVBwat4XGaWG8+l26zWtBkIcy5JP56esHp+gi0Me716VKVih
zTUQ0dVP2PtlvN/8zYDSzcNSvTPe7S8yrZS3WMoBtRM+N7lGFYcyAYORjjMN8Z1o
46s1XCq/qEPGhwwHBLIQM9flj8PIJQgzl28GzwKVtBjA6AyZig1BVHL6NKJfUdcS
P5y1C5rOots1NBMZpAt0kLj8YEo8B9VMGcigx1cGikp7nnh5bM8hBtzk3xAsjQie
d4bzkXaAwdmKdYqmGsoU5EZEkEzCUtXvDrvr2u6GJxvHZ31TcO992LFnwa0R2qFZ
sinTCfN4c9pfRLtqtnT+2M8/LjNloCKUpq20iYku7/3D6zM/0nS4ug4zTUihEUkP
IZrr1ZRE6cwHZSr3n5FSakyoqVy8f7c2dLj2MJuPzxpETIjKKZHx7csMp/YLrctl
Ka22jb/BCRjUKOIdDdSAPz9xzyqQBjCOYaeP+xbe2Ybf9FkPSr/NcnDZVoR2/X6l
09Vu2O8rHnpvl0D/0mfXKGSbQA1CjamAAefJp4CQ8sajGFDeEKizW0g2Q9LZWmKf
FWiBtRqEjPigOuy79pkHYaCdmbXQCfQmi7Ns+e8j0BOnzjhm4qWnHKcFYN9YqCAL
EQYP/6dVcc14WbtYWkAB05YgsniKn4VMFuI2ZEBXffVr26yn+I+D1fe8udG0LJSq
x2Uf1sbah/pPfA8epi9dhhJLzPW37eUmqL0Ygzz4kpdtbEr5iXJO/nmLzIAgws6b
K5LCOmAC7mjn7Q74Sm9jnpKf9mdw18FS4Z7wPYCP2fwjlSXeEtqQ4MOTb6H8JOG8
+QYYHGt4kQBaHQExyi03o0m1dmzeD5a/qf8A1CkRZvRIbMMKAkqZJUEFZzvT6CTg
clnLuld6PZogVsdzruF/nEPO5ViIBK/VfNLMlovZm6q71cyBgIait2TlmpuIF6N8
tssaHqmjKS1S1Xo8iHOp0d80XHr864l2S0e8FdMTsxgF6vkQ4FwLA/W05CaNgrRU
19TzUYcdcHGlGR9PohHBCKeX7ZJCI5c8oqEDkCT0alJdDHy00OFfYhtBRmD/Ab1c
ha4JUIlNREaMQ8hbITSu6VUianB6JF5MAxx6+Jw6xz0x6wHPquTA047BH49R1Wpl
3TtjlZ1eB1zdoop60bwOayfTNYr5NYMKLk/gzEjI4WCDj0mM15FOv/vm9L1quhOo
VyQ+0gw6NT99diCg33eV+9FkzYmfWHYsGsb08uOdf/Sy7ADOUpCnw/V5t8s29NEE
NnmMgCIL4/jbTd2kujD6Yfwz1ha2LjDXIJeNzhj291DVwFsldZkDbEBX36qX0gwK
WwPAzst2KzvdSzQ+S1ZpnlSrv6pF3i43dNxaQQqx2LAnmDIc1x5U6Oy24EVcILsU
O1azfj5l+tbS4fdTILca6PZVg1YzXz03ctaxTeVO5ZL6iILAAWz/v+d6Gn92rXoh
eiTcyHN21HZ8DXcGSbfsE19ot8cGXK0NmFN753uDegu5TDV7j4xFDRFHPlZgRDod
VbS3tyjEPpK17HBn4HfsEkBox2oEIYAqiX9zuTcU3PGgXsqxPc+dIFt8o8FVBjzQ
jTMB34k2ng5p1TKejLVHntBfThiWOpd0PdXm9/80BpBD/t4Xb6REKwFCaUhVPV2e
TtHWJ6xbotsed3zV/LXLqMNg6XyVYziE5YG/cjdnPawecjjuemvNRnWaMw6w9TXZ
yYFoe5lH9lL64/WDAPNn2VWUOHB2xgZiXMWMSZ/kJw8l0R7zPZiigQq8CUgwajC1
EGGbYSouC3r90yUxnwKgDynGwt1SNrUzVHmi9f1xMSlvS3fC05FBEEcXCgpjdvqR
FSjk3nBJlLRi2+RwI6GYn1qC3c2rX7IcDDkyBem2n8darPzdRwSi9huBfQ//bk2Z
/boE+Vj/l4HdMxVfZUo/gXkcVT1ZBoCZqx0Hg8RXvsOLRcidkPRgkoUFFt64h6Tq
S0l8fYIMmjlRaG8Dmxs9pqLcgLzij/q9IzMyJcvIg5dza0AMQ/nAJAcGBoJwTRFq
Y23EcODLViC7KYZ7zf14QVSHNmz8++MxAF+EsOOBjyJD01LficgYqkVaJNDLCrqG
e8CBTaCHSi9/lILyk9/eoX9aHO6VAeRS89I4Vwwc+7z3G4+uXbKpwlqo6IQRCGnc
3ZWe6U06JqJpbE1lvwJrpcMK/dzFWm009pBAlFoUvKuyUyWWa6fKy0o0MpGn/dup
J8BHVMO4AbHfShwp2I1/eb9d/M7YBsCnbrk6GJryFLsT57QGT5EgmFVmiBrLJ53Y
gW9HN6R5lk4EQtsybFMmi0MljrBaAp7mxdLZwodkkwIm44vF8pXUWn0Mq0LemEvA
ct7Das9fq0jWAsUgNhuzUpq8fPgsuobKLtCpOx32b9DN6qP638E1ghF+mTWxBHMW
DtiLItVDOoJlWDHt63k9mAtaTvRooOtcVRcXvroxCFDeyBGWIw7x6tjm0hSVClK9
rKGruOBC/F8YIadHf9sZDQD/GwhRsDyoO8q4SVX2mYpKWwMTV1dnjxrVeK3S171M
h2z8DfNCSEnCsfKm9TceFDat/Pz9o6K/wbpT38QqJ8dAvPC0TzNMl6h7TuyVkPcN
p8Y1MLIIcuAp5B54o7UJ4s2SXyHV5dQBuLeKWMqQ3bvUCmLhIOqRWKTQmTB/G5A7
6Z8H2X2Ccfy5vV6MG963ty4WtpD1im9Z4LZeJrVeGvWiR9O49DJkJ1N2yQac43Gc
Jrpf0blzRe4UmYySDkEJLKKh/1nnwYxKGF5d7k02HD4B+mTBFNsn95z0UUqF7joS
uN12oyS80kK2q/gq8Z5Ptu3SLDHGYZ5TQC209e7+uoy3WnYPNYGW5XcK0Z6qCsLB
qoz3sAND+pBLWfJFMbkG1s9SjB5GlW7lKS/5FPCl0evrARP93Ua6JV+npTgG8Aq1
vLaT0f1qIGlo6PqTMjo6w5AesF5KYVKrTr0DLljSM6XWBgHZaAypaYVt8f1zVMnL
PHGrq0O/gQfqOE0cURmIk2E7sb8aXYvyiSb5nmKTgS9n/g9Oi6Al07Ig6nExu9eL
Df89uuJIVrjCLBwwBq+xh0Om9+X8PMEZdzScBND8ps+IQUa1O2wwOVS4DTXGTzf6
q5Kf3S/O6zVa9dalvE+516gQPTETCMqbs8JHXcZ+k8YeNpLTuVXodS7KIoZNRw4O
/5prnWW5DurVe8LfpHYC0Bgczz/oWGNR1WqE23KurhMDAxV46oUeow+BQLjJVCwy
ynwU+GRuVkwSwe5G5o4brpmhm3XJdrjjW9uMCjLhdpc2rd8wOk1cuzRTKBk698KM
NSJZNblovXmOd0hlXRLZacovpTvizR2pEAxy7w7CuPN+49eBG7VP3S2+dvuknKho
UwMX88nGy+pQur5KRifLHRg9e34PSfWER/DgsFk8R3Wu7GhAlRhZNbZyhG5Zpxhx
rg8mq68ZBdTn7euxq20c8GWOfBNazRektVEGfELfN/qIBOjnm8ppsimtIDNjfgYy
0V8PRcw3Kog4wQlJVS2nrfVRc53M+aK9fOJiKUR2qYQx80TdXqaQ0itwFsrOpvpY
wHQCErFjAt85rOalKk+nFwgH6ji0YVYqv307fDg0GrrEG2vy0XiUYcM2OmgaZw1c
7ScALkRVY4rpRj4qdtaQMqPwOY1R4SdoNr5gfaRZhlXKiLi1ntJD0u9LWuer1dXj
67hWFEQ46wmr0ykCwJwb0phpJ1OjKWbPONx32xCB/nTTBOg1gJwPaymOQ7B0vcB7
Vbur8gpVnAiLNLARzcftlcWlGxNYiXbjJw0CxNwfYT8UqQ5MI2SIf4uUD3lYjDp+
UMFpbGJDbo7IRQwtZqZ6rnZr6GaYF9qAd+9/gIkiQva16enn0zIEM6kfIEWm9k/2
MO73C103WC+aAqTo+DXViWM+J8IieFN7skg+9Yki2Ra+8qgTt0yf5GKIjpJ/oKXi
OsQxa0mPT7UIO5FmFsSgaPd964xWI6s+9LOcG+HzPbzBqioXW7/GlQ2yjT3zo6NM
+5GJTrFbKMR0C3rPU9pXzYFwiKvSn/eKLemrkN10kE9+n3+AkdFf9flo5Q685KC5
RJBe1rJYsuGzRUm7wyJK3Qdbx/NvVaid0xvwD3aDxIXpKFOCNZb5RFPGS5NuAilp
69zVJI6jJ8EwWxoUQikMZ7pafpGeVKfX0/YGXhUqhq7opbJxX29K1uo91OGZyKB3
3m9az5jqAfiQYlHhsUcI6aEAiovfL2ikMWj2ybcBG/z66FQfDIR3lBSfp8QikRfB
VnBfUFl5BCQ16xWp6YJ4/vOdbixNUwfmP2sfU56JKAAGrFllFvGipoH0A/alwD/9
mIDqeHkuWDe5Q47OkBmHm7o2sA6aR4HJSUW7gCZNwb04hXK9+D8hymPioQbUIzon
hsT61kZskIzimP7mICdkHzMK05aMiSLNtOAOGxhAP2rLQlTHPunzbe0FtLidSwuL
2+26lh9StHAB0nUcGBNdmdIEIc6R8AT+Iq9SUzv3j25jYgbDTkCERqaMkEAsTqaz
/9EPzPffQHSzWuS2dB0pLQxduw3JHr6VRbF//hOsW9P4fxu85Ngfv1yuqGyVJATH
9E9I2hbYXejsVXNO5mGCKT7RtMCRnBXsrnkEHhZwy8w3iqCo/hgVXcmZ9mVB68gH
2AZTKeVtqEc1GSuR9u0l9GpPwLp6IsBnHGke4rBoSPCgetW0oxoMhnOnFf5Dr48U
BtD0y7ntU8Aw77zWoGBjX4E1OtE8ATjOaBGMrEO7uPVMNXnyY/vOIma1w+GSsQk8
GDF74IwCDBT6UhTJC1Yz3aZ3iZPLTuB/MAktcPHr0fFZOy1ouQoh8brn1hP0rEWP
8sBnHkazN7cJD00PSyXDJOjENsp8Bi4V5J9ho1u+63fgOHu/L9cB4q/aNefR7PrN
WlnpYf+sqlQyMr3wtmYI6HCQmdkocoJOTCfwx/oOJ2j9WdemzsMcOnUg3GGztVck
dRZ8ZnYkLoYuxCdpJqWr4VUo11E40rirUsxwHGh99jh3RHmad5ztvjqfmzp8Nc8A
gWtX0rikq9W5Lfti2MDKWdMGJQ4ag8n8U0NzXftffQtaOAC4iRhxwFUtTB+bn4u1
jJuro9J+Ae209IBlzYJF41bCFTL+p8SqTDrHB/jJh8w0OkE/B8G/dSUhA8Ra6Zb4
3OGSw62lY0nSxl0gGXZGN7Gv5FPD8ySQMoYc00oggIPsTW+CLBKuMLmh3wB2eMVx
n1c2HlKanT1Qmq2sKNt4wxVgS5DYABtwKFzM6xlOvBHPHZjvAGffWP/wc5+nSiiF
//fvVlClEBdYdpddqUAiuinMTcnIJFeswZ2ZyV/AAMHeImFxyc//Kzw9vYt7TtFJ
GU9o1dRykYT3UAcAWF6efdTfWU775yGtxcPqeT6ARlnBl4LJ3iUAoUy/+seL9+WT
euo+GMckxdiym+X4JYiKANnjrAu7XOVnKehS5dpaz7NcvdPZvpcVSChG3Pb9sIIJ
/gc7vqEO066+U5yuqdHZWTy2VzHVAIt6Wp3i6prkhT4ISyYpaMkLliIyQTK8Johy
Fx8Pnjxk4z1AU98KakBnisW8NgFvuAlpKvG9MFBkPD4hBMSItw6u/uf/18XTMP+H
wHClDDG/yyyEjV32OUN/9rHabBcnm8T0Id0pu+3lPmVamVDZ2TJ/ppjsDpRa+By3
n+OSHimTd7u2wgcn1LWNECmgC5s1aJ/A04VUb6fkGokn/TLSabOxv2fCNQk3PgI5
mQcQG6Kpy4k+fOV2jPlDzY05ZsSNXqhXZwAQMkrw5vKZfcyvNE+yWhrxDcO28oKo
yVpWopt8hu91OZBSZWzjNimaX/6MlApRWJ4SZpzr4awafwlt4EBKLMOHkr0QeUKx
lPhVckj58ut1BRN42kBxvvavdBuKwnFABwDHVyTiE/qNVLxXG5PUvdal/hqSYJkJ
JJtxKp3XhDpVpaveD8fJxhp73kcTWW3guSfkhnUremzVlFqjxc913Ql3w0S9LHAR
ApFkAQ69DDNSWIdsREz/f3YQIj8RQu6QMDYC6m6vahTipF3rRbEiQF3/10QeEspp
0jOmhUp93k8t8EQR+GAi/GlCVtSeLgB45iFGBr7+1Rla79SzFXdFdH2T7dibyVbz
XjZxlzmBKlqDEgi39MDrOEFeFK6UbrZ9Lu46vxRVk7xyDv1tlDNIvdhWd2YRjvkJ
mCV0R92XRTMKafmxMeq4RHviKeLkMJxcefOEe2tSfRLLryWfqH+YIBFic8kvbyRs
Do2WV2iHV/NpbjgfujJ98LK+n6vzMvy7Sah/SudMBrtClz/VvYjL100/1utOfE2t
XYvyDOhMAETB2fE71vm4Vo5L2g4CwWtn+Iu22vSUjLhuUIym+Q7Odnae0A+lxCUU
NlDF3hwgnXRNzTrPEswQxwYBC8yQckLL/uAIwhNZZKp/xH5JbmT9WPggYZ1wJ6xY
sHGb89ZOAZIzOsIG9LY80zwJXJoPGjLB4DaBtzs1GsnkvBgh5QAgordkWcdsoSwe
lH7O7lEtf360XNfnF3YaYU2tS2E5olBsNx1N92xLDvkMLJ/gr+sZzC7FoSZtha0n
uFLobK7voSoZtglxqg6/HMtVHdma/H8vYzQcnlSfuk/M0IpDuNpitIpN/RhJxJuX
b0k7nDlogjB6SyYj3ToOQFUwfz1yCTNhFzR9SoEyc4u14CV9/lU29FrW4nGxJm0C
OAxqOuO+/COgQRYqBV4tGMY0a0ukiRxtydkqxoUuZfJnPM5gSLU2Eki1kTcijTbF
wKfzBw01kaHjiJPtPDzMBrQwovfaSCxq6/7fRmqKBLIKPFiZSZvK3uMzmV1pGrMF
65ZIMWsCKiokOeN9lZnHJ0v0RdWsTKEVP9UBAfpiMhuxGxYy3neibBleBo1uoI7j
QHl1ZaoZXX8Nyc/AyWZ2n9qea2h6rL41vpORCSd70YXEoLoSNY0U4ILBDZcnbNtl
M9xtTKTatwTtCxW1CyMEdkNoszvnPRnetU7dtS4af8RAyH0Hibb9G09Ssq0zjOlo
2bufd/K3g2lKT/IGuNQxU6DA6scdaaI1FA1+g+IU80l1SfqZPphX9pBY7zkPeu44
rbLEvF7KyB2bnou6wWCqQCsBbZqQosAcJnwmik1LWLrqunM6g/bAWgmYEWpudyL9
dHOxIi3fJ09CArZeL00Byd7LVV8o+QgoJ1EbuOHtEusd8OE56v0nR/Vm3kCBoKD3
D5UGWNEba463UeBaguhIbwZjwrROc/4dBvBeqQrp5bzKhKfQz/ma16axWE+CHCi7
PiRMj/Y9OtgbthV1cfzHjSyfHyhYbB23ljAu3jT+/ZFB9BjNaz94/l3VPEG4PrY+
pJZr6IKUoIF376VawVE030E5cOoQU3ye+x5QyIA45PbSFLTUY6uI+IqxNMX3zrxd
BEOTMr2o3aul+mW03W70XpzQCKIHg/6ijqmvm4b/etGP8U8irscpZ9LYbcVqq/2U
ZLReGinHh8joo4VvMPXquASxPZjvfhC7egu1cwf6LhuEPOHZm3c7nn9PIh6WDEsx
jT6bPnw+spPLaDSZGBCx0+c/BreTndcqVt88zx4nvAvhNeUT3xbDQ72b49pnFKwZ
ToGkkN8FcRgOlV/UPC4KflqwUzuyyL5R185TfQEqQArItNwccai551TcaX2Efh3o
mmLQNWrOr8CIOE/Jl0TNF16YYlvbl2B5E2Ng/hjzGchXTXLpvD0odbJnvsC2n593
agZw2/lCz4My3Mi0uz2Wqs+7erEzrJCuLjAfpA3EJQ2x01ZzdWu7vnyqlEX6bVgp
ZCiHYMt4ziSKdJRGqXI80+CutpClNprkyVH5WmpgvkwACwCmnfWA0ySaHyNq9P1W
OiD2z+VL5LU+Vj1t8rr2CJF0Ren9NPbWVEA+RLFF+jJk68qsa/xpP8B7xoA8Lr0u
648D1M/KBjXVn8d746w9ZWroSmLcHENo2VvgcRl5o+xO/XnHQ5QjLQ2TJDPNLj1y
IqhIH5VxaOxy5vjVUu++iAq7AbetMTSXQzKeCuldCTXndIrcWteo3akXw558lIkS
30ZN8G7Tes92SZ8sjM814LwYtA4N27vxjQJA4rd1p+VvqcMeg1XpcVzPQQML8ien
jjWv1L0vZYWRdGoT5P7e0wFF6AGymL0SSGVAhxgkx/Jy9xgRbGEzry9SGpoJ07u/
cgshwrS+FbeBywwKzIrr6G5A1ulOittux8E98FAAfuShMtqOgvi5BRYZWiA8fuF6
chESUpxriD2MYZn9QWNA6NZ9BD4yRBXRcK4fmtGanzQr7NmrKH6VLfXX6ZowJsRc
KK5T8dg+zIX2hLoxAUiW5z0fFRft7to8KPXnuRwPpz+83OM6bcgIkcKeYMl2rOur
800Di1LMmOySH2dQxEMCHWn4WTpBXoFezj7puMQDU0L60TBuKUhwlUPeGjbpIX8/
mPOOLan01/bZi1jSDWcRkpLsC8rRUHjEs2NJOHIK0IvwZtp88loGXVwLcz0pQ1iv
G/Q/71RUsi3CmMrWor6KAPhODU0/mx2tJum/aGDc+/Ai0dcJUI/fJdF/0dICwJbp
nU39lM7RwSGFtCWiAiHzjbE0RBy+SGAj1gfQPLuHbK6zzCIsT5a84/PfUJyEzS34
HoUsl1OvJA9d0nLDLOqnO2BS6Hspg88yonz3rm3WDh9Pup8bblS2nhPL4iMZ/Epj
ZkESPnTSt69Gv53P4yrTM+1K97DF4dtGbMDgHlJalTlU5RYgFPMR/3urCGhKcN3p
uiH31R28wALNSoyrIOqhaiwFsf/RbqyPyrFhpgXVZluV+MLFaBL3Ht6e6BuPJcEY
AdqG07OJL4hsHCFgwI5ZH7FwE5vd1AE5O5qQPaFuKh3gtlD4u8x4tbsyiSsFF2Xu
NXIXTBPnSYjpzgCUnMlAvMbJIJ+SuWDPKvGQcmYXoVOBiyIQNZoOq25wC9bnbSQI
FQEB3xnC1l7EJSbXzOikFtCfxxKsMMw59cKirSfXj3Dxvly2zjO3lVROheXo+9vv
+tzQVCr+Sn8Fc9gD5x1GPJc+BkSMW5V2x5i9ktymeEmwwvXe7r4ld93Abn4J9vxq
/Xjb2T4j0It4OMYyNcUBzj5jvceoYdGQ+gYXgki0/ZuxQHuueFW7NsLfQ4nv4Al3
WleGGSLP2RLKIRTvJxBUrsk6vYVwjwweT/NANjz6L4r5FkUDSG/ipOtjoMmNNOf7
9alpcDapYVhgrGPciLIAXQiMFIRtcyDiB7rmrekuLdXUlhW5hrfY+4bIeDNZOmyt
m3p22q8bA9EkvHT/dScTtsINH61puQ1CLH5sf3ROWVZdbxpE2S9H3RpUGivUKk3/
KTLA+eiVhRlTcIin5LTkjrdJRYOEWAO+qH0aFDhkbwnRt9+E8OCC5gwvYshgDvyH
frnAOSyRYxhMnIUfgSFHt1Xj/TZ2jKZ3omxRRKATs40WE+smUFM727Avx/5dhhTr
+D4v6vyOO4Z/7YlWOtIL8jIVb6MgGGk6uUIDvkNp9yDwF0+9wRXnptiaWZtRIRVe
upAH5IJ7QhROM+hg21Tz/HzpYZG+UWOX5mGJUb1d5QvU5jPLoudQ4fXDSzPO46qm
mTSTLjbnr+P5PeQM1zCfuMwGC3PMAyucBbcun9RkvBY+M/3Scf0g70ru0NJLbsfy
EMMDJIpTdON7TXpRT7t/4HQyrk3k57tTzF6uaBwn/dU24HDy2re9nPPB0wkvL8MX
Ydc2m0lPk+1zV877OfOw4hnE/Rnqe5ni+zvcB4lYQQ9YPsHg24q/LvqrWrLN3az/
pP5tMw5vdq9975ouO6CGLF1O/2S4g+n16P/rFAJCxZp5qM2aWhkRy1o6RTr0hVRq
nQPDr1ba7jzWNlA1iMxbhcZFXG0AwPZ2APcb/nVD8622qkChMQiory679Lu1Skgd
iFA0Kh0Jea+HVDf8vOVsBNywCqJOESN6yllGTtbMPNeky/Wf4rKzKvUjuiB8d3nA
/LxWMyofgP7xRqwdgbv/bH0NvxLs46ZHpoCB3Xv2X3Gu/PYE9QQmWe1jpWOkCAEf
h3DyWCkv/NXgcQYWSqkS4hKYnbLYSCRzdf3Yti6PPpkMPjkv4ld25ejB4Xhd3914
fycXyeoEOhPhJFvvg/pev7xso/QcWrPw+FslPUGGjpSiB9Eo8HyomIsRMArRmy35
yEfDHuj/46dj8hf4gOYimmJbKbRl+qx7CO3mm+eyZLRp6614t2GFaHnEiTojrila
chD36zVfHU9JE0AGPSU9lc4ompi7x8s48JAlubua34XOTW4en29zo58nH07yUoHJ
2zAQZmckq2F48Sgoq1NgwpzPdjfLrFgTCCb1FBmE2KGe/vVdhYRsJR+KwhZFi19t
CGQxvODsVYYu9PpWFehXo5zpmejFzJUJ/GJddyqikdO7BC96nLhW7/8azLfe3HLm
U6B2nhF8Wwiv8Mr8csAB6bJ8a8aK48u7QawREK0t0acoda0eep494WDk5OPBXbQw
i6TlqvwBsJvtpi7vRr5xiSXPFuTuYk0+9y5ZB80yRuh7Ly3HIh4d8N2KOTtRj1A6
bzsInEJ6C4q2NATHvSDis14pXO9KnyQclYRaEg6zvY2rO691Wp0xvCQg+Bgouh1v
H7Gip1RLFYz7j9isNgD7Tg7+hY/9v2DioQijrOvrzxVDKlroshzW5Eqo/0hy+dKf
wjKJJjdxjfnnxp903rdDNjX+oEaFYOkBdHb7QMJAeEa+ZdvTjEfBdua2tqnqX7f8
M3J7fMv8bppzsI0F7JJ8f2l+yEMGz2NtyLocAau/f39gXblUsapKbZyOTKMKfqKI
WSaBswpDvXo3p5tKggvaYBCzv5c3hBARs6vwhFVeOV9RVgZup0dgYxSnCzlvbx6g
RNymLF8us9d60s10PlbJEmK5uQvrT9lvhoevOpo//WozKYW6uP5ZBhukNCtdrGAN
FVpkPjja7J/rL5gVHZ/rOl/+TAzRl5CUQojJ8pE6Q3lxnd1aZFB1jpa3flzch1t/
gfUTIfkBqinZDTohXCchXIfamSHJcGNt7AuFj1A8p/GLaX9y84SXG4/x6XGAPT4v
r8YwoF7lxoI3Y0VOvU1imjyQvG9YsL8T0IhxPzbs5274liil1ZtrCUJttRsin9Rj
LxwYglhUrcE7go3W0dGMcOHbmRart9TR962q3ZC4WrxL0x8UFI+n3qTZnng9KgPN
86CIpAEEnMaqFBeXF13nW35HXFTqabfmJKYf48Vvl7tHoTc4FmbVvxVxmW0J0IFs
wQWVK/HpZs2eETTE4teTTKnz04SfeklnlxwsmKIo6TkrQdb7A21Esjk/SnWg+Qwg
1mat+oomaepmBQk23UhGLLsiuBnIdgfW8wiX4DIr7paXP0tzOtjqSNcBBs4li3hy
ojPxo9wjBnMqbVvv/ZGhXzRU4xGvjw3QImYXS5PMzhKd9EuW+2esg6rUzEodC74k
3u4U+CoJvL1q121WoMTZ+FsyDaMcpBtk6hWwVFmKZJzyirw7ZEESgEdPwvCJUsc8
FjQrPlOfWgL0D8xVLGscjhKNF3I78G4gxCqpe8bTo8XkeRlPU3aAgsCMWPJWW3W7
MgwEW1YrYyyJBYQq+hefqUm89e6JylK2FX6M4TARLjqa0XxzDmH6OIduviBrfh9z
H0vObbdgDsGXqCbrXFSZkKS4GfYVi3xLFXO2SUgk8e+qMsqfAV3TK97UYHVZSlgA
4vU4WBgYjyf4ERHjZ+Z9mX3YZosLh8fiM2CBGUgnDW7MmTZi3i/Ye53xBZ5RAfer
kxmiZQKDYtBqiw5x+OPcci/94FGOCHVnpx3EamSK0TIyrkd41vGX0m8nPCm+xAeR
5K+G8mWT3AeSluLgHpCRFDy6AhUtR4Hp3HoOSERKyR8DI9HwVF/kuysa2oXjXPeO
VX0JlvEdmwdlg8UnUe7zyjULejFdw/A5Z+GxBj30eqSdRPAHHHaPiURT6V/F42xM
okMu37dOsTeYT/wWK6v9v7PUiC5fDXWs1BNCIIcNBHQ2BG/bWRSdlwC6furd7mY4
SJcEjaDMPRHaYT2g8xXIbk2TfC3L/IDcQUW7D2guNjDIg4CHlF98x6ZGWA1EdZPJ
r2HUgWUtlfQygL+jFh+D4gO/wkDsd75VycXIMTA6/N+GO7/XoKdAUXySB0yhakIf
0hs8Av+V4D5zRL904ZBeCGbSBpW09ccT4NmWYMCfUeo7ImWj4dh9pMg0KpHcHNgP
AlzcCxEWhmhlTlMc8O8KdOdpwyFKHEDFXSs30UcU4qRCx7eZkef+iJ3IQyCqXVAd
wv5R36wZ6vYgUDwxF25u9yop77VceTXJhokadLW7gX7nTEIsS2/xavLb0zLmelxX
9lzYytQZy0JG/BZVuj3l0TGFJ9+d8AScX8C+4zMYynR71Yu287NblXtbiImN9gOB
biT0won1m8L25pMrDprXgv0pbsIgVa5tkikwA3nPeOlYkH04NCz3KC94emA+y6HM
/+MahLuorcafDezaKLhOxjiCGRCLtMwpg+fhVcZEfhK0CojRxggy9b6GEarBOw28
Xvxw8Tk9SiR9eGKtYhv3IqcE34JiXXnMU978Oq8bjxSBz2DL7ngkz1mZ9OA+onQt
2MwU/QgYQKA/kD2J34ax8Maszb3k/HAtdRyBsdZcDwBeTl9IPZcPMXl8XHQZHE6O
u9/9v6TWk9t15lo0TesJXP/k7+Jen4ZI2swhkQdfX5PWA2q+xMsTevvAx8Dal3VX
I8IGShGFcgmxsn9Zwc8tjNHkX48Sb1GGZfj3puctGgixDyW8m3ASGZ1Sn4ddwxD0
nXGT6G6sc8uc1c03tiG3g3u6IOuH8yVqfhKUbtBejDz1T91mjSv27wUCM4AB99Gs
bUovANZurqEcONblh+oFIg6FJk2J1Zej/XclWFlftQWkBYmKUdYCXFiz/uzqDwnw
QjmWYN+qRO3ZPMzPFRDkZ2NBN05Pt5mgZISyyIJXo8LI3jlurIk0DNPp6utI2b3e
MggNEtW0KUpbYRguBhIKomq+uE/J08nJx5pEESsQ76nCRMJzlp6YitZsOPLp0kw7
swRwbsDpoLcdBxP5O2SFoUsJvJn9/8cnGKTTtnL6w4yer0YYROO7LHdSVe920jO4
p6OsVF52c8f7AgbgAc7gVsWp8gUsMmcTIOlADUYWKmJ/Jo8++6pSNF07neJuJD/T
hum83H4Nu98z/IDGrkD0XO5+BOuIxOOb9Zik9ixq0now4tEL/g0qrMwO5l+L1m5k
JE+IRwMIXbN/6gpDlhc5RhcMOaTxj4OR3/aCqaLFNJhtj9jIiSoWbhFm4F6PuVpd
w5fP3WrBV8oGPxZtLw94Y9ZMk25fANEqZOkFFsN6IQUdG3w9r0jO7ff85tMST69J
pVZ1ZRzrZY5xCIRQGMsIwRvuH8FW0fCTnSczl/rT4YmVv7pxuhccwYdKDzoaFjOX
pKtKzKlUr7fLCD4ptcuUIYuqxDylkfA3Z+grX2IIRhUn5S65oZkfTxW2OTokXnzV
kTeGQr637sNI/RkkCT3YGpB2KjbZzipZEJqz4smq5eHTxslmPa7ZMuDNz9d+5cal
znY1RCgWc1ip0zlDa81ZOWADDxopZHgPRaaGaNsv+NWk53GgHaktYTtvcm+Wx7+1
U+nj2nLm5w0FtCBsuoiMMpp+Xz/256TeBYazwIyoo4eTsIXZUPmHW85uJSft5FaV
bXMFu6dBWpL6iVkJ8NgaLbprFQvm7I9aGWd2ipIkXVAp4HLTUBmki7WyzlIHnWe+
4qk25pbS7ortVUsb8YDrN/PeTNXIv1bGbyEYxiecbuR/ZAhxS2EzXK00AUnXNhSA
onyk/yAG1yW0ZgMcA63fNpgNXUgFGs29wN5yJ2wERAvoqpzDLXfNCb/QeLQ7Q3Of
k13ElRhiw1dFL1TOMMez9VOMDG2az2Otn/6IPqhLRR8OyXa4qpjrT+Z3U3zNXBsW
7gzu4BTzJwTadG+soFJjxTTSlOQlhIy+RqSnuwP+gvBkYiSlP0LzTAzMVga5ibgL
JyfITb949Q0/IOdqggQtehxUL/jaUBXTi+A42cKkJWSluUN16V3g0BkvIBqJuc0q
e0O8za/5RFmC09I797y/oi6qqM8llCX6HqjB2eU15X4KjVJQy1Lc3D+mkZmwkFZM
KngNo3lXp5w+3F7N0tUdtSBuCLru9IfhsPj44iI4UEJpeaiKtkS4haGKoYSjuIga
pnwNuSnlkceZEeDCpXYXa+K/635smJyH8FeTOufMQsy02VNwupbL2Ik/aZffIxt5
B0XbQ+rTSShSklXcBaYwYW735RiabSSioabQ5B6VoYyMYetydZ9L1dZqIEc8xNjS
uXiZ6GezXW6XdQSbLV/DNzLdod5w2KS846o+sdQAIXeBg+Zf8i7UjcogQuthTXOo
4aXTV0tVlITRp/ifLVT/m7M6kbNP0bJZf1asHGoT29uPTODNpq6RJlr4wBD+m/7v
Uqzv+5AFu+7880PBUKWckiL6cFBt2C5WGK1Duxloytg81pkpwct+TyUmIb7Onedr
BJp3RRZiwldnbBjwDa410GaBN030r+vYjI4LOyDxaOalXH7TZBLh3LSkd/T4JOky
D/cMAJiJuatUs2CkExejJbUn0K8nMl/R7xZB+YZiRxRtHEM37gZACF0dmDHBCT/b
o1RaEqY8n2e1GFoiUK0HwBB26iXTybFRM3texn5UH7yZyKCeJg/3bX2bFzSr9C7x
MKcOxty9/zevoPrgrtSC+t25S+4PzUuD8qSOAR28MAty2bi/mCXNim9INFeYtXg7
8M8PC9gkAg/n/m/wCkOZXoK9gy5c/mJBCvpqLgFrObFop0bb0DBzdOmRlMP/ouQM
nu4zhLG0tX/ZjwHpFa5dxvWmBTnmhtYZTvgPqoRnxaujA3BFnKRUdtD4E6XZsgMS
sXnQOQs/S6ZPyc9YL5LH6Q2/EvgfyNDlLY6UU+712ZAl0gah1he6Xcq3UdcQqCup
+YUJ5jEesULiNg2RVKC55modxp2KiIRwVT3uxNcdojnXnlUIc3jL02SwdAW5j2l+
KbIxpkCsT8eeUBQcuigVDktPioLV9NNuK/XAPicke+kHH5dkd1+HUFgX3I9FUap/
LwkTalOGH/ccKipfaNd/F6c6W+3RQGUG8VwyVuPRu0xsP2asDVkOYY482NtkXFjj
PhaW2liUECnGrjunYd9NRIRG1vj3spjO19sdT3Rk/sBJE0SBXOlWPmj/XoQVneJp
uxF5fv7uKvI+RyTEQfElHX+VYZu75pZXHgeQtwKVD53hv5a+jLwPOMRrdn0cYpuy
WoWAOOsIf5FzHBn0emqRuHl8RTnd6fNuzrQyv5b6NWNLM0/7xh3lNvhYYleAx6XD
4fH2/4d8xq51lbNkG0+tYFjFv1MDRp+9DGFhXFVWKRdiFjpfKQdl2h3fPVw+TERy
avn+vokrpugPFSPcx1so01a9ja3/AUxChagWmwrAE3ObNEifc4LnTjDanwoKYcZR
ZR4MaoEkUfNptbKvDz/mj7lp9/hegz/1obbvynbozCySawbK7FywxsQvlTLZr7kw
86oAtZAqANNKd2kV1Xjj5w+WgvrLhUT8rQKhtLvP8AgZcktX0NWHUYbgNbyZqfRh
YRBO/xqOFT3NoOs2fvutB+nhMpp824H2tEgwyZeYx+ZJR7cAcoSkqr9GBt2neBmp
U53bQ3kOqUX3mGFZEZAKPGfUFUqX2wDIs8pLYtvts/zRpxCHLu6V5AgnJyiuNCjK
ctbsQfwY9vkXr2DIm1bW2Tk96rfzBcnX1viGHnrVkgK5o7RkE6vIcTaDho0N0Ylw
WxFjMk/JlaQSYnmuhRBq9xs1+7BEYT6OknVcDZvGfVW3+xW9uxk8VK2xWPWDP0+M
EF5Cloc1W+dxDPhKoHXwuTd+HSiKCSC5V6tXqe+duGApOayxWvW0j50twf4ZVP6c
b/xepRHfvkYQ2S4w62Vk7oNEh0htg7wDRJAT6Kw8YgEOHTGEhfkSQWJsYq9iYL6G
lHGWnb/7TC0D8A15+pEOYXPqWMtD81PQEA6uVsy/l6tJCTnLnEdNQCKVPiQKuZea
wtb/F7twOf+7/QoccV33UStRvxQKV47apwyyqvBMHFm6vIoEGX7+dUwedGq6cUej
KuYgK+kndl/af4PE2kEGlZdJRv7G0q5C8hgQSPLpwlJHlwotnAhbXf+47OgMFskL
Cvud57p9g0WafTmlZivjRppIW1L31DniVKX/0l1VgDXk52yuugPRIhtelKf+7FTC
hDsQiJ9LWIY+FANgsemGzxmydA/oiD1R27zpGKmJhRJ8TYkIUW/xJMxADB77iFdg
mOR22qKE/oGgVm3JbdIOZdjfP8lZNiHmbEAwJGZZF3xcRBYpV+07DRQBqas1OqjT
z0vhrzJLCJw+Sxd3nFWs6sQKlELVs1eLh5KYYUj8ceU9VCPIJ+yxawOJAVRuHVen
Sequsmv4sB8l98XbHcrv5F7LK2SxAFSQLusCNIN/n4ufOkhhYRv1j4S0UBZAMoCJ
ecT3PxDUyu0OJsJxkZ3cIxUoNXnND7Jazu83H69OyqHIQam5OkWfFu6kX2eh63+h
aek1/qdOJy+t/LGvzhZ0P/PewVI8HcEeFcZ8l/y6pZe3eU5AaCqveK6G9DiE39WG
hfKACFBxMU1Is+sWO2ECfvLhRb0n9oT/HUikyX+QGNhUI/ckeEC1l/Aoy+UiKV2g
f3+7IT6cKmVRr3zaPC+3/zIlx1a3e7s4amJa+z0shibNsGO/Dmenyx9NjE1KnGu4
qMVi/cIGc61YWHyHxxzjRVv9NGQJ9dIRmJ3LpWzS71kzSeR3HWw92ByhE/gb2xJ5
nVL5L8Vkp8KaX3fjky5HaKL8OLMBdyiu8pB8KkWv3F3/QiYbEK2yKfqnN0RTPoct
pqPR6Bu/cCNqiNTZUSonvLRwT1jXxwhtcFC/zm07ueHNWvm2w3KFRy1nRQKNZW0a
ED0esOY2w6eKL8TqO6wDOulZft3Wdd2sXIj75Y38HN6EUsBbLe49xG9l9/LDijh8
HdUznvM9ZLSe34QJd0263yWlF1h7GcbBYu1OABgPaLAo2BQ0Y2Shug0sTyC1MI2G
6gSyELnZWh/Y2Jb95h9kZ4wBL9PQ4qRP7YTkT2fdPabe8XwFTCTfiK+B6Kfc3Gdb
BOztv5WgoVdfhkZSn4zcSg+eWDXNjmvvVa6e6hhYNB9mC1u5Bi2Kd+ceYu/7vN++
zs4/A3EEfDv95DlfFHUVPfPXdl8qIhypouQqaxVyS9zwySyNIL4DQTzyUhVmPGsP
qiDBxYUH1z1SGe3jw7BH8Xu3P3/+qVgvCPoJnJM257nXY6DRsmy5gIGVo5J+OB2J
2D/PpIyHBwwy2WzT24JgrQWONW8OVem0Xke9VP4cevERbV9IBEX4BjK+gf7X3Am6
OZ//o16ZU8LpOw/aXDuGVYsoX+C+u3A3BYJ9PFqncK3fL+sc33eQ8JcMPh4pk5Eg
rlEuJBXMXUt6B7HMsGPv564HHaZCgIoQakkcWipS1WcTWBDdJbbknT9d9xqrJP1q
miT/ppTCzewl/KYePF1SDbKfwmGZmFVNbsxr1ZK1DARTH9Je5dILhQuWdC8Rc7Rx
T4vehO7ThbYM5eXffKzPebqy5JlcjGPBuYFFKF0Qkr4iYX6/prNrclK8nCY/SAyb
Y+HJXNugA60hcmM4XF1oEdKFInze1CNAA2UwfeRSQsokgt/RPAVu7Gp3keQqmmva
C4WJNNG5e8Hg6Fcvsnf9T/rrVKazX4p8n4/7FsUwANuHg09YEAIT0Z7XH9NE1Uwc
8WXDGptnufmYRFLbuwK57AE9L6f3FD5l0EIU5u/yxWQi6K5ZD6/1xK/ta/Ll+Q8w
fdFFgmmYI/icXtcyqmFIs7nyIgh/DXrU3+7UwsZ0iK3P9id19Ud55oVom6B35wJa
p1HZMYnOotIpm5Yf2Lza5E4lp8XIfyut43qz2BnYDEHBuLD4v1N+Jds6yETGC796
gA2bALJWfbbjm333uizQoGDHkTq7DVyyL0VX2Ji8CvssJ9+7jWzIdftk69E1yutu
+VqlMxe66kT6OjR1OPRalGt3nPpX4THnsq/p8DmYozLTiq4xQA4qbG8DFGuo+v7H
mergJevsFi4Ad2VCMwAhD5XS3ZvYFt7ajsC1cOT4OxjJwswcEn00QuIcEpYnDloq
UPT7Lf5TY60U+TB45VLw73RFjfBdilQr7Ndpoe+jl7zSgc3AqcUJ9jV64hvLIVQ+
Fc4VLyRcDcniPAjzgzvNT+rzBlvDcoOFvgz7WCkzvojQjpEo+AYMGNzBEGeQwJep
0VQ+IaRF9z9fG9ZQuVJ+fwsmiLBTi7GXp6K0g2d8RK+p8OVmNsztW09z7WjcqdJn
z6q0TaWDO+PNfpjxNZ0B2dP2BAVjSgghDrceWcgwwjrha4PjOsR0pIXyvrxcFtz+
Jjppj4zHReNFLmbRaI8tdDzgElFZvkmyoLh8RmP8eQQSKKwJ6aOt5T30QrF1o+An
gEbua89PcnyHCAFlc/bLW90LcDCvqarDk80N8ZaCi/fLCU7i7XcDLyrZ5h1usvr3
nwXfTqhxwaLXtFeNpvnyCi7P280NFL+VqJIdTVx7PihwzC6UuINfECI1yxcN7a2m
zSGgqPdJGg49ukZQ7jrV1qG5Hnqr+s3v34PLLBd4M+tr5w7yzlOpKnX1uwUG/y+p
o/7ghLJq8bP17P7UkkH7cKsn5AcIwj6KJF/eEG2zadEF88QtLO+dUbGArw/yWFZG
6rfZE0uLAwhqUEKpS7hLrx0LX9b9vYIP4JM7fR57dNDTEKnTa/3ahoja6nb+odTl
cwsXxnsT3e6dA0RcW6p6+ZYJIYfxXSk+aFUU0iaNc0wpgE1qCxM7/WrMJmoO+aFi
WVAppJcv8gntfX7Q8eueXKMMyd2SwwW0DNQokqyiaos5Bm889YjwaEHG/uUKSUFo
RJxaV2HY8gnsp2YmEiqQ/uJqsniiGuTsOSBRt2XdSu9UPgMTd9QoYuaCZtBj4rQJ
UV+AJgeEPuAaZkXKBPxHVJ5UTZSCx/n7BXtVyAa/gc5MpLjQqY4vFkwig+eWoM46
wl1V9caPL6l6a12kCLG58mZqacc5dxrqzcsP+cFmbPX5AoAGdO7wtt3V15V+8559
tc7zqV8N3QzAXwbr0GZWtCODNEMJYwGsJq1CW5XzFwGEd8JEbvSo6eI7xYNiLPCM
idqxkTftBI6URLWB9doqjBGbOICuoObn1jY4ZtyEUCElY+7ExgsnDOb7vogu2//b
4SByOalsLLcET0yOYEQEK9ycjQ6+R+5jNAkdi4ujtQ3nFNRaklHoMSWFqqoXlXrJ
GdUKAQ0dpD0Ju6dpGGBtF93qtDVoAOtBevaPwjcytEUv2WJB2Uz0MwI0ovRxXOas
OBlUIg0vvL06YsWQrXpWqYaHY+hyVHojSX1KAoOP1gt5fVZwUR14IbfbNMNwyiI1
2QYgQkj7iUsqWhimt4K8fABmbgyhmwKOAJrpYd2eeOAcyGzEHvjpkUXqRT4O7As2
/zRNP2Drok21zPSmec8/eIu18nL/hwFsDpzXh398Dr/fyKLWb8Tsiop74634pibO
9yxiL7YBkAyAgBB1xW1SxyofTaWSrYC7wBTcUeeYFdrLuo47pqlZjmPQasjM6bae
ZzUDf2T9Qdbg9dASJrMvwIabGxDoRmf4r0IWQT0IsMah8orzqu+nPq4Mqzohw35p
daQfEW8OB7YZrAlpKC0JfjdSmCtD76EBTyHmKx60HVCs/v4Tki5XH61NfjUu2xUB
RkmaS0VdZIT1WK318QnWyHBCGMlp84a0TCPXADQZ2J+84pBhu3BkQPFVFheDAity
7SLBd5MbCyhog9ZefyJG44EnltZz6PbxhVxeTdbn1/ZLGU7jznlELlG7QFjWbcBz
fYSF15/jEIWO7J8W9yAqLXpzOaMPN0/1S3syNj5LsAW/bOi9MJsH4iq6ljlNo249
rJVQAE866Yk3CInK2WLdobnxApOahoBoZDgpPaWxc8j5YZsfoo8Y+0UnjpEf/Q9n
g8zu4DVoXuThVER2a8NHA8HQ97zx7OfrVZ4wGd+IQAg9bdSpLt1+Q0a8EnZHIBHe
KdHnYUR4SQmODpVfo0mxVNlnBsaQijuTvhGr98EaO/QLSNRTf/u78ejfwyuAT/4q
QH/NW+j9OZiaWXUE8e87LI3+RNPVBD8LCBnfJCVXGlpnGWyXfkqLn9lR8MH2/mP8
T9HtudyayCth2WHtzbzyGbXQoXxbQgfItPHYpt8cvvaG8fH76kVW5RKnrf9xjmdc
Ve4+AY4WVV7MuyEFvByGpXWOBXVpxTi53oukHOntMdI5z0sQ3dTgFz4o1rzfG0B1
gTpxESgu8I+wgP8n3M0jqU3WfyW8Q0fV/fiPSjTJWCksRusAFMK6k+LCS7je5thH
5R1yaamS6ibB4e7EUB23o14sdPSs6z3kItBMTx3ztT7UuV4NiwsnZ0HsjatPggmg
0Ha9WGR2+7e1a2kxTNtx7AA8xmq1Df+3kgjfCHhdyt8OtQulLbw2+RVwtU3nPhrN
ha2XZnPPdO9NgzhBVYQUrtnYqSQsyba4ly9ip+jXdbB+wA42j5807BR1rJrgKEA6
9OEWs4rljaxwpVs34JwZ0ZTwNw6qEKwomnx3UnwX6z1iVTKmtJlKjsePATRKC2Ze
bMjTB9kRTlMMnZAiiYYGinquWdbHHchl4vZT31ntg+Mm5+I0HuLRQHtfPARCVb1l
rpVOg0DTqeaoc4+0zZ1mwiOpe0SWMYLsmJ0va4d2ijmpuy/SVjB3utfhss7sj1xm
5ETC0g9ePsOL/nBGDN/io7hVpSWalTWuphL+kiQrFjaOgtqMxRATx4hvlpqp1PIR
u2yJcirlW5Ec1oSvZJXLdL/vX+Yac3TPWPs9lTPLVk6aIBs0jcY5KgrhNMQ+oeXT
nWn9FsLTMp0ehRXOngTEsdwb8OQ8s86zmIF3QBe5/HOOx8Di4RGW3cM7k7fOVlV3
8/BmLkgNEPyZ9kqQZPDFcc9CAWVNRPrpVZ2w4ZhY6IYj9Ma5zGN+gOQy/2j+9elR
YlQYldcM5mQ06XEK3BN24CSwGLWgTKmv39gK2NwAGVdFyJq3bXkMBZBzb7Gdgagw
jY3551+FGTa+B4g1ToIyss0aT8mWME9lgXwpvlpwslLG32RWH8ry5RE1VJZupSmo
j3asLgyfHrKEmBcKb3QmZ+Rq8ReeiUWAMRAbgohsbly+dHJrE4rOu7nYETsEKiu+
BmiMr249c5w5yNfwzvJOIojtyxA5YwiE+N8gMzYG4a9MmwFJUfLdGj5H5YyX1DFp
8JGpp5yTWUJY02jdLApLnUHyQ5mzsyaJTKk3Z69bt3dRA3iUCMnuNgV29Idt2uXC
mSr4BV7cQVuqQc7D2CoDr6RH8LFWL+r+BwUmi/uMEBrzCFSoGAVNBDLfszfTnQ3I
6b2uBHJWNKQYB9j11ByXfW+sV1vHfdIrkVRYKEGakv8N8572x2GRV+F1AJhrucWS
u6HSSlTW/ugZXY2rqFa2NFPlxGXw6EX7eTZBL4lx00lH7bSSGMtnehU1OXRZ/eKz
3yx6YT7ge3vmaIBXuE0MwSsl2ipynDYhURTZ0t1eZYprGFjBBDlZPa3VX46IcHeT
kwf+MmNjA+3cHbgTvNa8tUU6I2c2jSJp2a+jkb9lQwXQRIBWeUW+ybd+z3gLrI0j
iC88iVx9goyFt8OHAao1SCF8k/FPoJSIewKry+AxbrRSIqiQxqoCH/SzM5P2o2Mb
6/+SV6SPZHIfT/pyx7w5YMTsTPNd7vXlqNMqlZLXeLBjh6nYc4IQNRrl3VCJM1Yo
yu9WbPXwE7v3HdpG+r6EwKXcB7pQJEedLfsm/5NhtEg4rRQNQBSPrClfPuL+shUO
aWJLlW2cnC4fhWdRx1GvSndD2Yv2b2OG+3MOuMUVSCxZD1EjfLsKetdA/FWy0nz9
GNshMrgm46rX1mhgrrapsBZT7kk8jHwTIPeBFsmdKodzj+qew/xF2sutE46Z3NEz
k/1SO0T3qHwOoj8Hgp4GHS4VCpmQg0Gevj9JAG5SBLdb9BsaJOoedEwqQ4oudpkf
6qiEdDCHdV5wZe2Ho/D093d8r0aULkpP/OdH27w3CVyLxTUSnXkA6rY8ZAqeZqbU
rFtyzZ2hQUhcp1sP1uur4iTj4oqYNLt5pA64LwCygUEFBSyGwpRUb1IbfEm6yQxe
yyz0I/D874bekykfI0dvt296t5+ZE8AFmoyUhnQ+TOGdsmkuaPHhOg06syC4i7qc
4ThkfjlBR+LH9B63mje+J2Eq61eCalDjbjeauqLHPeAAlLnjP+HVxSKbJjea85V5
C1iZ3MU8IpjlBc99mxAoLdeitFYIb06mOGdawsEAvqfmH4vVRSZ6dF7CIOFTNV4c
+bg855DvmE03LsX+ffrPgQGLBsfZJg8eYSm8RK4fysj8MievOifYLONDyDwSU5RJ
Fx+QT7NdDWky8Z3A1sPxLgma/qc1M+AlLvwP9d/qyrQ/2q8Zv9s19jzv6y6eVaX5
dGp8hH2M0PTK1GMcE/nktCIt6/yHbndW3FdWccXMrvJC844xpxdgfyRQ9X2xDR3u
tNP3OjvLOFZnEFqj3aiVkn6wV7yK66n3IznsIRtOWOrBG3Ph/L0p3+erXamnQGCI
jqdc8vw4YeIJIgbhh2Ky11r1KfovQjvjEbkeVcGxtrwCE2MHjVhyCFIMlFSnC7IL
NgrlROa43bIWMNtmjlT7Oh9A2PvHTL/F0lFPAViSMlo0DNPI2DRPXJt3oD4Md8w1
j099Z9rYpJ/tmoDtJtjZ1tp96eJg7Z2sl2/ht/9qbbk9TFBQpyZJdZs50pOT0nWQ
6CnRccREpn7V1N/2oQskEiZvof+EMYNm+txk5z+tClUkoasazH2LeFfA60xF3Z0u
W3eqCksWgYlIY6tAu7Swq72JDlyi+E7pI6zk+sDB40aUYEgTsxJJbRo7Ag3QFGxM
K9ze9hgQbrZyiE9urwR0r3V1gcX40GwDNNHLiGeJXTE+NB4Ht2XeOUGvUQbHUlGc
bcLkuT0uNxDAlpXi0bD3vVZf9UilzmW1cC5FIsKzNpG+XqxoS6zcMrZBRSaIK5g8
WXfrH4tTggfcQTk0zjDTyM9uM9VJ2NWX0t0BNGKLUU1FxTV3+oh98Hrf1V7uCena
SelBBq+BoPzbBkNp5KR68x1o7bpmMaq34bT/AX4YMT9lrpQ5nnolrSfgDO3K1jAc
n9ll7r7sCQpxn/llbiwi95//jAJYlyLEG+UgJTDtZtnCvpOp7CrgOb9+2+qbv8Ve
NDABvNNY6leSbFBeM+eP2nYvCPqSSaMFtqG8XLBt9wJyLcjKFuTbmMJO4ZPNbK3O
GQ1/RISFyqaQKkgkr3dVCIxBK+LyUZjnMOHPfQ2PBU366hM3RiYBa4FcjtiWN3oF
Lzw78K/tGVNq7WOhhTyrwoACVo0IuHUp4gzlxy4AdGZ1hsoYGhMgfSXZC1XfFIs5
g4+IXr3NoLi/qFibM4qvi9Tcp+O4dcHTDnnQTLIBycQIw7dkNu6PkS6EVib7xwXZ
3nb7nTNDUTo1QpdUoViz81QDY/DRsKBI/0Osl5CLSYrgjbhlS+jpBJ9KnqfBDezF
GyPmF96C1tqYSIomAVCANtr6e/vcoNCFoy+vLYbj7f8e+BX6yeqtQreG1MoYwS1s
RoalpKA+RcVtrIWrPn66rVRQlFuklWg5e82VJwjqSadw6yxu3pk4GRMvz42XkQa+
Go4ipTmy5wE66HP90b1x2ubBcqY0+8yPxEgPuEpRbxFwgrrtb7X+t730rcigLzUE
0+5KQtTKeV5GnvpPl/zlX62U69OVwxXllkZUmbB0ShdI6W8cCa0GOnl0ykjZ8Vd3
tChTCmLW9wU1Z1WYiGI+DQRkrRevXh2ro94dLx9FHCSeFCzPRVpch+0d3hC2RAno
OBY13vXK+MY5OcFjuON0u4oh3dHq4sRotKtAF6qMDYDR7y4NfNC67vyzqlyjPFvr
msbAjOwCp+PHTcFisSSuqSRl4FccQgHdD/qD/k2MIknuBFJGpv+A6n1xxsr5FQEH
gZ/62DMxSPTL1PMGrmykx1Tqn3i6TVJ+gHD20sTZdHo6GgufLEh3c+VoS8FgMUz7
Gz9OYzzYgDs7nuhzkaR9LOxGG642Jjp1gjo4veZNWIP9HiZ4m1HYPOpcyDhI3w9b
40mcLO39xlbVfYcMubX3Cx4F1tHPD0R5aytxdgNyc6qXTFQGbBmleUK/Qf+COA9F
tXqSUF6lF3V6pH2OX+QrWLZ4fRhJnMosm5mccemRvnANvlAu1BNpQOLp+pHx7/1s
kkzo8eKyhzasOWIxOcoaCVR45gIYf2moemJC/1L0wG17gxq2Ci9UH/b1YYogVkUb
EhcTL2voVeVzCV5+9yZFuKgvjZj5s12fBBLIqtJeP0LxQu7C8AEUwx4zM6lgdQbN
WGFJqjbzEU3vVDvXNEAWt0fmSm2Z8xGNj2f/nPEJ6t2BIhb8e6cpAkpU1GZN9kHS
iy9sL1wy3V4wI9yXygACCgmUd7G7rommObZHUNMsRJsJGBvnUgH+8D/3viOHSTad
1KbQtRyVgovXU1pdZoYjrk5wEqY0cW+6W/x833tiw2KP7myapAx4OwfR/dxlmrtj
9DMCw0jZdS9ZnvEHIXenO1tBso1mUP9pXFp6axGeaFt5NZA+eJb+GByCymX1ag/z
A6yEl7ARGPCsyunN5ryEAcBuuwiI2lvoxSXHSMXnoEtIV5H5C8BpsWhksE4xnsMq
/DFRAnw7cGBPzmFqwb52dX105q/83c39fEz2Fi23UILaAM/oClNcy/xpe3QUX3MW
Xwincd6xgjCv5Ha7FFMpbdyDX1KIdDQVLgc3o/IkWGfATyECh5W9e85qdE8z/EDJ
cAFoxxYJjYym6NqQehSM9rUY7gsa0H3pXccXWOX+YjXM8j0MBHEEwSiONBwNu2hc
zOiyUeM9ZMG6QPSXyf+5fx5xDcpszabXiLPpywhRcB2U+dB+S4js9fqrPLN+3CKU
tuN3vEWJIY4JM+37FWAalJSCNwLElUog4bPqC4fMDuE4fFD+L2sKg04iMi12rIa+
PMa9BymcrgXj67Yg9mqOarRiaGjcaK/gUqXGxDCyEj7yEfKgGfL+m4CzYTOUcZmi
tfWSQVPzQCXbHTMRVGtaNPgD4gjIF7bGjttPB6Q7qcTTK7rAMHLmU1EWI+HFlJZj
v6gHs/6XFT8NxgzQ9QgSElEsqC8MfIrTZSupUonWWKw9Kj0711OQBvFZsxKnAFUQ
MMOi9RQ38H30lEA1V+FzxUl/vv7jaPTQrdWPZK+P5RgRNPx48+ge5hnzfCMswZYK
HZH6+UGaUKu5sAZzyqJ15QzsyhwbiiwknTqZT90cDWnEzLfY/xu9ufGHS66s2luZ
Bl8D9dtR2p8DghfzqWKB9JEt3KJLfSU4NRHKKML7CTsRkw5BeGYy0dS1QoIp+Yg1
fTAGtmFJ5K/lIJ3/Br01e7BD5mzP+uGqS8dpPObc8UAd+7CDpv4YohmxPiVgClP5
Dl3Q0kj9GnJPjkC6jy1bmnQRCuI3HoZzfoGV1+iqE0ALjVa8Vplgp01if9EQK7R5
ZgI09z9VvHT70GIxN8/ieWqfx0AQqXW0l+UlG844KAP2GwJRO9h7YEc9N3+egauo
n1ExjehnxOg+3USlIlJEBF5T1Q7fhqhWgCmVddmd2E2Rr71LdMxaePW0Pu4/FVya
Q6dq6OmwA0tfTTPWbxhEc7PkdQCrog7LQHuofiWKxJ/QDcO6Vromn8z7NX2LPNps
Du4YgIHxoJaLkfMCS7wytI46VGmfAjjkIS2R9p7UJMrdyTiI6LEP4uDjgSmm1Twp
hePCI7B9wAoOvP9rJBZabmFHOY+SgEbTl7OV5pcMwDCSM+G4aZaV/t3oYX9gdBhZ
/zPW0CiWU+c8FpIZxFmNnYfCeC1ETP5lKVKj5u4hL+F60ozGSKK1O1yluEHp1b3t
/sGKHF8u2lN4f9vyidWmcv8ebXObBRIPFP7BsgdPiEQ+Tb8UCtd/cJR+ZraczwH8
cIJoPMw3VnQVvN81T1wvQ+/h4Q4rcZrA9iAoSHiUOYGRuLVKwviZWUZ0I5MmAzsO
jVohPxDl5g1Uhvr/zPpGVqD6toPl6l4SvnXr3qMtDKVKS/17GxIEq66i44dbESeL
+3GAa/uSyLtyQlCHO6hqAfebMzmX3GWcvQAp9xi2nkzehK6Y9RO/UJM57OitWwiS
lpIgbagPRPDdOzbPW+ut1RL4i3UQwazYBFPJJKXXMo+6zUUuLwiOaJ5HubyXc6TU
cSBONDLSIxk4gCcRUncYh83nIx1ZTHZlK0t44JoL9Afvu5iJpUvYL8ISnrpMNfwO
ajzN8OyacBmThloN72Dv06h1Et9xOljQhyDh8P9eGZ2H8koLhxtYPJAqE7aBjydd
ghypNYk3KT+YQ0Ie3iUSG0+mzF3bupEPJjxoVXqLkaZ+NAVb//hz/Ug7gbLvS3d/
fim5JVVBXGYgyeR5+vPbg9YQswenNQw1wZwCAr3DAHAhonYCckz+1eZnJO97xH+A
et2hwJsMHUf/3dAkhMPgp8GWuJmPNj+W/6nPviQdz9KVYO/XtfwSIG5z+FB+Dc/r
tenFvkz0J0VQd4lGj/8HISs3iYsCFJ2iw44CN85g2cT1yeP/eFZK/C5hAEXY7btS
58IUW3IMtiY0ZyqyAMhbi2Y/Wu5OgnyRc4e95O0PmB+EuEUOcQHJ1qu30okgvu2/
O8OihpzZVPf5xuuecc7SEDP3g7heo+Eu8UEnnv1mPxbfWhMI6r4lG7ceVUCtfYic
K8re8a79FKgFkRzSP+vOipq+eG/LibEPwXC42kkFfrEJN0USjM1/gHkie5kQUUk0
PEKcjneTs6WVNHuwwaGmfdFiqVvhyJ7IEkAj1Luwa50X3o3qFe0HQ3uFA1X0TOay
rVYCSnY2CH1mtjBuWZCig+4AO6iHHxNI1UUk+m2I+P0GTuOgvZkIxDZqE4WxzjW+
iqGp7ofdLRvEtYgZiMq6ljotzSQQvUfuVz45Ji7QxFHTRhMhC1RduOsI0IbarDKT
wjNJ7TLeMBQ958Iz+XUCvrBYByF5OPP3joJUR6Y5Fy9FwdH1CVdMKaiPRNKMk/XG
MII/M7s0vXleCGRnI1EcaJAslfJxeeLtDb4aZDzVy3laPH+pIEG0wThX2Lu9oKLf
givlBzdbU+ld9j5mOSE1v9eV2WY4e1sNypTeV7Hk96qw5jGLkX5cQqf4gqA3GnEk
b3uhfRGjOxAmiE2uxqfBR9ncgVp3X5vBMZ1XpUOjZZC8w6EVuezyu3mh8m0yt5vl
LsRNh1bO3qUg6jLqR8cGIj3z/n+Jbnz/9xxA7pM3NNTuvZ55AdCCa6FE53I7I9u0
5BfjN6S5sz93syJtryRrHND7+3d20yFlTgZ5L4fZrW3brUmjJNfMO3u1gOrGhxmm
wxJ8uIpdg8yqMgMUCx4w9quu60+yNdzQnQdFW8c2xEo4SDXJ2mreHrd+iueH3dSw
1y7cda2btDIiKGiWb//uGPucEEqBxOrMWU1STXaHb4/k6djOovsgU8Ghl1czf+ss
DugFMWwzx5PdprOAN0iA3roIYbLtwOBJ9dsTMiYPJYNmvj0OTwgfDoFCx0BsaWYs
NY8Saku1YRoULjwygCy83hILr5/vHW15DmFidpchEx7WGvTooKJ5ebQia9BEe++I
CBoGvo3OomJ6FzcQ8EOOW6yLivW7c2XKJcxwWUXXmmfihB49BGh8GqwSQbFZWy2d
8LYd2fn3Tpt9Xmbi8YD+qky+zcIifO+JzAcVUUNiQnfuU4DCuUYtbR2ZbsdQSUAf
7GVfswD8e66dmVYThYh/PvLCjtIvoHt19hv/ducOQqMPZeIdn0DPOhNNuxHnXu1k
nV/rO3tKuaVsoD9d5xO8ehJsN+5fzm064FbluyYEXEo/e1zdbjhNSFC4Ch4JKsm6
v4nWqf9phov+zX+/4WmB3E8ikRec+iFAR0yX6EQK0lPCV8MW8nAaDnH1t9WX2hgB
NH5k5WcifZlnPsRMeb/W27hnLzkJEooMfESDKYzjO/QC1sUU7OXrZN0Z7a2MJb5m
hdNa3etwVLFiGL+JUm576fdq9KWdGjYnzq8CKyYcVpcKnjMmTZYuHyCUDwgOzkkL
NBWnD2at8uz4LZ38hzqBpczOg85YQ8QGh9fuN0eb3YqV+yIgZWR3DUlEhSFMBtuh
vLchynzYtEM1cZFTM8j4R/F2pvc4Yo0Ky1o13W7BS71XRL4aXkTC9XrmipGdKs7F
gGUX3lhpBLr84mSHKuWQeRrRuuHxtz8h5mOLOwoP8p+psEjJIBRpNwoE8BvjLb18
UxarwOMJtFM1c5xAAJ7I0F3N9ZiqPD42wuEcnZpCiy2E64YpQnx+ttKZ9SyxA2ZC
7dJl0fhB0QWr6b8g6Dp/d5PwCmurmI8m+gIizpP4jWorAAeqIyhH+To+RmgvtZga
AEb3Uoyq3zumMnSQc6SYFvaYx1bYjRVjAclT43OJ5iOp+NdLIXMWU0A41J+XanA9
7dG6VeDGfq4bNarQR59F/azIbWKtl+L/PmhgXqRQBXSRiTGAGH5EMKtWgPpTCAPH
vKPGPegPr30jEY8WUPbJqCUmdVtDpGdST2VnoTgswByulI/r6fN7WRzTYw/SXFE7
uRmtqoG3QCa6Lc7a/FnfP1LeMJH1Zf17Vf/fcgFk9jrG47Osh+f+NoWoWwcb8Oc+
by0rswce3U0MGfo19q+Gr6U37olEj3dGVzX/2duSluR0YIcZrJA29qzK2KHTYOz7
IGmXtmxgvKrkk3LCXvKZQKpE2hfFvRnDbwQwXYxodMmu6V16RFL7JLBA6ZqVf8iJ
QL7aJ0xNGSD1FJv6R/e9j7VnU6pkULOBF6kxOUR/kjerRvppoBL5I4dYckka0yyG
OtfnDV1F4tDPpsHZ0uFB2h2ULAhTl2JTJt3kvwkG7w7Er5wLDo+OMFJCs55WEqJM
I89ExpgTY1wAN4IXgpM6dGAJ4FCx939iu9Zr17C2cC5g9PH2hPCQglSVoTkUIu2b
3qrkkChSVfB3XZRSmrmLC3jyErfKiYwBf2vT9D182rCIulI7s0xem3GtDb1rnrwV
oYdjSiorn7r7bBhltRa7zQ37Av8r9r8oDVhF2TWUVeaKDcShMg2ZIIYaVJEFrWl7
jeDtvB9g7JoFgZXXf/FsfxMWnR9ShMJnmX5Djn6F+rrD6HGLbreZZdIPfigJZ42D
vJBGT155Qn6w/kHeIGZUyd0IeXKrACCnniY3Kyq+2N7eMrKhiBR+EzLQ+c9nogQq
uRLVGfzsvim6wlgMo+nEktPNS+lmhIQHkZkOEs3UZQM+XhiE5Aj1hcp90mpVe/6u
dvlOfpRAYCowVNVD7LYU0W6FDn3HS/cU2WvKuseRYahsSX81oj7OgPhJe1IlxvF2
c/IcH8cgRZVDsq7bchg1QgFETnco+IpluHiD1IqNKEwMXfRfpzK4tRlnrF+OJxjv
1V6utXgvzSvoTelPq4DQS/W1p/aCpxwPqlcaWDNjbaQlNEa91HVsIDsTLLg0wLuj
KIvQ5UtHQnJ5R/myx8ARNmpOrAD3SpcttcuAyXOPIgrtg55RrHQ1IkFrXaqJFOi5
QQ9i1b+xq6YbwCr7xR+vBi4H92rNcGfKRL9k8t48NM4/qMW7zlbRhNdh7NaePe0s
80JW9DhnIyWuKg6vpsjjE5YztxtK8wEeIeSFcy8y9GxUVDingoMnC+3qUQe40SJp
Byzou/mTlTcBsKW8btTbuTIfzD2KrlDdTAnu9bGmlqz0LanmD7s2Ke+jfo/bgR+x
VcjhABaHtbAQrlQwycHOjqNOHG+ui23ugMrLJnIf3/NdvggdijHmwx7jKMl1WvcZ
7itD+A6EwmL+Vh/NFeHcUBMS+DhPfnshhDoYsP9IuGmVVyM2DNgUcngNo72oXJ0G
cWojqL0RHGcvlROtpzmfMRqgAMK+EF1bFlj5hXKwgYVesEVu/gjXg8KQEXg4IeZb
mJc9ctefjtmq7OTzp66HgAnS4NauSR2Oif/1s5xjBJoHsWLleP72qjoljsgU2kiC
k84Ntf44PANUbVrXLZ26O38kJEe+qJMDF4P6A5a4iaoUmE+DZrQQRBowlOzOspjq
cskp9eg+7Vv8PCfqqtYHprfiT47R0YUofvzr0gWF6fUyB5hduFUrwxrYnF/W+Ymt
e+oByDekSaqEPLaczsxSHW0mUsVhFuWtJdOc6c2cdoStygPV6B9tFS8S2tAiwRJh
JnrJBfw3Qn+jhXfdGrv/jysFbRXiwlddxPkdnueXUe55oCAyrgU1Revzk+wqu9GB
BAwtpLU4WYUfX9Mq4I4uUaMjnsnmbKiZiNtKt6QzK79hXGmJoLoCneuQVIA/Jrl9
BVG+CgqPEAM9xPIRDBnKXk/vNRC9XvCMTQP0HOTDb189d4/cMMZm8cbcUOXKKrQk
Lh3usjC+eLNlKwEN9fA0vDaQrMmeXWAO8vfTXU5GZ+Q3QkQmQ6ES0bpCvf4gso7o
NTcWGzdviRi8rJLyB7WrWjWKi5akzdYWoApGfa9NOa0b0NK9oB7sCSnWAMfkZxbs
1MMI9y0L7z9bc19XWolHTEIn0kQQ0q3T7B09Q8Yh6A1tKAT/FFuOFKlvSEqGTgIP
KizbY0UYR/nqHaLt4KYkYlkMbqRjcqoPM58dAnVs7Wyrqy6ipDOjuqwQrdK3NFqQ
LhR8Ardkuf0PerbA5+CuftitNyoygm5QEqjgEwFE98dtMRBN+Yx25MfncIptAbyH
F1GQ/p4zPMGE54gXoJu0rXvxnnDmEzJdgeBEkM7Umv3bfmUtHzXtq4ZyORtWmCaq
KLULWT+HXSJLymyVPrXAIJmSUNN8nQGqoZSuAtFc3/lSBBdObN2aBTcmXlmx2FxW
G4A1KfF6XAXQAnmAgsanLjS+GNnjBtVDvzUMJf8xZjuDOXdx9Q7nled2yGrlB9Gw
1pFIYY85T276OAcjvakngDby7wGYBmm5hL7AA/b8eOgWN4WpCFqQzUQyO+g19Gzq
GHFuewERK97fUuxPz+dkx2NS2QRWItVm4AlYaCCeoKJ1ZdDHj1PfPXIqC/s5FXX5
56Fzk0Hs7L2zKARcT//HOh5AgBpzm9ba8SnseU1iixHssGv8AEJPB8M5JUCOm9Uc
VNIIBUR2yAI8yXSeouo1zvFDwChuwZcvnsE2h9TR+vOZOLlfgDROlwnFlHmJrJkv
IGTc5HgXpNB94cwUklxYGp5GwrIglkAt2sPI6VPSdBvCSJGN1ZZaCz8eGN+WsUKg
csTGHbjO4IiA0oIYyvV2WmhXJZPpkD5VSkrDh+mApejSnSxAQIDMB42fXl0BT2Wi
0UuYXU1GCoOuXroJoeWOmzaq3tzyzSXyEtoWMjB2UgLnAWUkxfuLpOH2wlb7nvpT
sKlcy5af7rdfbY3XgI4PKHcdh6+FEopK5TduHu1WQILwidROovBmOcv5Ih/TF4/L
eoRIHNjmD/z/snOEay7dZO3VPbK03oVjuGguxoToc1PtcyLNxTmj8LgVEj8oquUL
REJG+3mafsKU3maS9K3VPVS2zv3jkemYrbCMyFwwYwSpPTqeXey2i4pbReqRN7Ob
NqQv8Dv5j3GFOSpEtqiCyw+BBEbHq7bQIlJAvlXmVu+VwzIp+CARLd//qbfns1oq
7jUAEn8VJypCHncKIhqoiP1AbhjOBwmCSYJR3iOlUw3tPTaYEcAM6sNLAnyPUgzV
BFTvbtbQMBYI+ggkc+00g1CW3AX7zwXoQDjoERHicjX3vXe1lIuN6C/yzIXdKMux
Hk6F6ctGG+vS+ylhPOShaCa4pMbT8BMbbOOmJPZj/iKjO28+PcBjbtNi04N9m2og
ZfBlQ8GWiO8NRhCOqaaJ9MWTSLmLbTOnaw6A9pZppnWmILuSiWnGyAiBQJmQFeUi
0iIawFK6DQADXiKQ8rupML4OWBc47Xz1dY3HLw3RalOq2Gab+7bGS+lU2QanqrSt
yhFxn1YiQFEBPVeRqp5PwZ+IJAAo+hgvWt7gztE9hA+lJrHepHaMORSJXi32wRqg
Ud6kMuYkP+GW23Kd+/xFrDfsDRJ4nTN0XmSF0SNzwJ5AnXl0bEzkv7AGVGYi759y
hA52ZUR9OfKkVu3AcMtxKnR+B/gNKa5LuvGeykNLdQqeexfub1m3tOOzCqngvZfi
o8kIBBIbmbmpQnUitpboBzjfDVOvto8nm4GXBTxlBW/AHjuxfdD863117pTTluMV
Lc18JI2xRVRpItBNmHJehfk+bnUE6DQ8gAhzLMPvSIAcd7bbHoYqC6YT6dYgAvXL
a0zmYxIrjXayjKbpcxXB0ON7DBxpmQg9S6RXgATrsLOMWSyXMvSojI/YmybwZLsU
/XPXa66kooKXTURoiNSqgOGerFFO2P3MH7545aG///yK30GtD63tAY+Rq31TVgri
GgKEMDURNnY5RWGNSTmPIqmRt8BlTI9oP/i43WOgjKId9zHSPHizPZ2xEMzt9Qny
o9sg0Zi5PfZ+H/F1dNKPmiLv259OmYbW10MIXZy3OGJ1hY4/okn8UvAS/CDEtGh2
kfbXGBg0OJ/iuTza/Yf/EgCnTBnxpUOQSyTlqNqZSPZ3EmA9BoyT3WgeZRz+JwwC
5rw4m8/qjx9OZSlzP4hT+9bOpIiodplkvuTo7pEcWGd4MoOwnH/yYPfJPBEHAAyU
A3IgFG3PLREWwss57YdLZOWRvjZ2YG3YH94pTAG/i8WYl8xLE5B7eiF53QFc8R1t
K1Q/sQyXNXENGM6cL0W/QwYkH4m5PUsZqsPKW/2UNxRvBqUutQvM2paZTeaJXUQs
3wMnNZ0Dr2Go48N2Fx/Ru6kas69U4U88QoXo9gVBCKCi6hwQYdKlToMaEuOoaSqx
VJbD6Pqbu4p0tBmZkFx9tQsU7UmQAh7stffHIHGtuNR0XqZN+2ytVfogysikaA8w
2gE/20xZYL7lCq0Ijq5zrOi9Yn7ZnEsQE140qdrLMde5lvpoA2s2e0diOjL+XaND
hVY9m25PO+Qgd1YaIxKifXt+4rOTkYvSerMGUPdkh1gsVDp5KLuInWSFwKotO786
y/Y+dz4adr85C4aMA8xqTDbllEH+WjEjoN06GDhKw9nZnoOV8LrDWwmJB/WlPt1o
4/mL1WaMYlfl0vE7SUL4PapYzog1dG/OQzFut1Y0KUzbObHAcrUlYzDi0Bjh+msh
oZ5j9XslLtezs9WyohiZY9qAlPM9fJ85+lvTCjFv3II2oc1xQILjOV5THPERBN0s
3cTKZFkHZf4qkiL3QyDdY4oFkXKOWN/f//u1t3I1bOWaVCWc7PTC39twE4TLFg/M
jca9gTWYOHA+bu0Avkqg8amydZIn3Qsd8ECxzXYY6GHN8taq5YmDMgxgULVawUeZ
LBlB1a62mLhmV6z/uvbukkN7Yl8zAF82chbhjv60oagWKkS75uurw4ExpUJCNlbQ
ctDPhuW7BEL/b5xV9if2rKDh+5Ll74THSygaGb7qAmu/ZZ5npDfjKVrv/m0BGgyt
cqZNzgbwkAA4YdScaJhGv+SzWRyxYM7gtzrpAFpyuZj7AtrygJ7Jd5lq5aNiiOGG
klX7cXYuGRplP9wzpbzzRc9tV0+iAQevNGX3A90iW7RhoWSY5l8Hq3umTxWyY2gk
PkZ+b44ScRm6e4p8ENcYGjKageO81kOQhmXkCs85Msu9y3gOKVOeSk9NSjsuufGn
97jiDdPQj/PcAhRPT60IUloJ/LD4+My1GYb78HD1g72zATQypG9WcywX+GWiERkR
vup/Dqr2TV/rezlFySG2Y12C6fk0z9YO+oa0Ze3aApiy/5jOE/rxj38ETJ8ZKu/b
TvIZj3bvj0sq/5SwLVXvP4ZmFXpjasQU3fSwnGlXMLYXKduGXbsKMqVsmhYhy/Qg
+W299S59vwvSfEThkTzHGF6Zl4UXZYJZfnTdaAOjyuRz2AkwoKkiO1/x7psdihlI
+afX7UCFzBidnObtmnnUQluOlDG8+R/Ju5denC90hTlc3oGPUenVf8WkeefBiCZU
8UhMzTqKtdg/jYvELmkji0oM5+ho+ywCMq+jo3fJXIKdUOPprwiKPn7k20QnvhXj
eGZC9HrdQ5ez/JbUTnEcAeUlR3/FQPTbQ/Ij8dxvaO2Q52lvWM61uLAPngWAC8Wb
TWLojxMT2rDrcR+yzuCDjAvOJUHrkmpQ2V0AZwjDHmD4qPcq5vT/rMkoX82XdnVh
oyczO8btKuAAzh45xd4cpGSUEV6/j9jNQk9TTyc9IKBZT+COB9zg+v2vp9wX86nC
hybIBfzQFtvMx6STalV2dgmJHT94Lb1vsa0H0Z8IGAcR3qsESYZkmaxFMNjzaHDJ
CjQGmI06k13r2ecXFCuy1yD9uWkQ5sW5hd8h+2/pxuTAIzFS3iDTYoJmZm/CkRJ3
2qgv+VAeJh0eWBRNTSUhurqJJy0pUiweqGYJKFPWxAmD/f8lSQfGaX9hfA8WgWkL
Fom4udnHMwopnZ0u63EJo2IPKkxrbAgcRLfJLv6rpiAirtvu6SnqarSuTNupOBFC
00e8OX4vuQ61rGUOVcgQKrAuIBWDcOGiByr60pXp+QPJMXR7buMYQ0Yp1vZML15x
zELCoK7YtbCC92PUqnVgGExikbFitaY1eR5nxaVPYtipkPnpLpCYQdMI56fGVoa1
k08bYOqJAPqixbVx8XqSu7i3ly4xZrppZfJrSJq4WmYQB+goWDSskI7WUh8GTylg
zEMoUl43VgJBgzlWNuO37tLp8zLDfedIGh1NM0vex7O4Hbsl/bV1qgJBzNzdnFNK
PHisT+22xFetWZ81e4K8UPirC97+U7CsdwasbRN5gXe1E6+uMR6WtcSm756C7cF6
QIl5PTFskUT4Y9SG1IrPpXt50pqoUSTZ0YURb0/4PEsNEcobf5apm4oOWfQ8IT68
rV5IfSr/0g2u8Li2dVjsGZ96QvDDA3lYB357Ey/XktrMB4mii7u5THRP2CcByYJn
CSYfUzxqV0UhcDYUmNcDtFAzL3m73sC/FUePQiEIlXluZ4etZ2lPoRJcRtmORlSl
Vb1FWthbvLIl0XtA3cZB/tUjB7aOC/+l1wQZ19u6v118OsFtbirPfL4yQbi8g8yX
uVwbeEx7mnsbFG8towS5eJSz56h1zNscTzIy8l169X+8XsAsgmkd/PHC7UqUfT+M
73HRZn2/aQxMKWLO5JkJ/GQXh5qNo/1r2OiBfRl0Vh5oM+07Q9NVc4jJ2JGL7BG9
ipJLW1IAaqD88aKTlnlMtMMn+J7zjiFGov6zx1/AA/RtLsZ2m4JawKJEgiSmTVsS
LiwSC82AOAB299jSMe7SydlFwM95uTKfAoCVhC8cSn00ulLu0rR20jlyBFBJ7k+J
1v0Bf9wIekvJglvz0m7YAaNdt7IQRjjdDeFTiKX7g3v39cU93aWSHZXEby0n1KIS
4ZGriJvjQpR45VssoloRs6E86YLmgaKGfOYrRkSHE+70TAU3sYS7yQUGqmVBKgPL
P9CGt6PoUr6lgDVuhEQ0ghEl4qR9C5y3mpUXLmZOxrBa2SY/wvPUrbj0dw/IaKXr
UqIx8I1W/xPVe2ey6uvALMqfRKdzIRBQyEwunahBCLRCSqwqbJE6PvntKIsNjViw
KQ5U40cdOMqzOzhItpGWJz8A6mt7ph3XxG7dWnb34ESWzKwNPD6zfV7/VukU6YYk
mXXwj4cbMZo0MpKVfMUxDCpR4wtxCupZ27Du5QDdU/hzwRW1HfV2e2dPs7gBW+Qu
zS0Z3XYwTpFss//u/qgF2Uq/EYeH2pzpb96tAd5BQAjFToLAlUyQ4xLZ8VMXbU1G
xetdANRpInGXTpYEv0hQHq8jEN39/AkABSbflLevwQ3kMR8GOC4K8nJmvECZ9TUT
YmLWoFEixi7lkMvglWyDiXfZoJbzwzVMhiqs9zGYjohvoM3YOXT3enybpJCnH6wF
yrH7iZ3SUlJzpvwrjow6Zc4XHmiKBSi4bgAhSNpL5cDaF0C00HEsrHoEc12lOHaO
jEC+M5N68Vao3g1+OodVRA1H2UM4CcoKcJCkm623MAQPdU0uDxQgLLSo7+ajgXlJ
Z8453dQx1TePlngL3hiz3oRRyBigKFvroe3GAsmc5UI0yqgTCUggYWZuTpmdDVfE
uRbWZ4vpHaKnjSQsmulQen8BOVOzQ/gA+tRTK702hyzUIZSlYdP5oOCZBGB8VXX1
yeEwCg7ZgOyyrzUOxG5I5PTGs+95m5Li48OgBTu3H/sCG3XAihGwf5BOyKPrK97y
M1ylJhYKeM7dDPBYznJ+2YzvOfp86vU9ObWSvancui3Ykmsv/JsHulqgy6la4JqT
fpK48emSleAjCsI36vWz3qQM6hUCzK1ViFzX7O6nVoGu8iO/f9LhXrT7YY3OP7Is
BYjf8uXxfkJi3q+aoRZ09UKfWhlaomfu7mXT7GlIQsrfq/w2+LCc1zVd6lNK5gKb
pl/ulYApkyulTqe/dX8BKAaM36gdtVuzfUB663ASh9S962OeUqjZOR69F0ZIA0jG
Sel/1yAwY7ZaexXZyUspIA2yKw5MRPZZdveLub0+C9EHHWuleGDlsNREPq617oWx
54/X0OQt3m9fdhEc9Ri5Psajf72uZhAdWew2sYWrXHl+mPnbobIZC3JcV5455Pk2
gm9oaEWwROEmL1XtHdNIKa6nRBgzHx20QJh9F9awYw3JG7Kb9om058MAS5jDUIhZ
qXbNNyn79QwRzXArwiwiUwxLaVQjDxDexm7u0wEs2liR0lHOhvsfnOOZ2BAQrUz7
D7zPy+FgxBJWizj2gint2I37cAUzNygTYpBCn0ssRHxCr26ISmbx1o3ePkpahxi1
R05ZMQtbc+fvbKTGcLoXsPAUohyQVdxgKwwDBzpmjnIFZEnaOtaJXI7zs6cfQMyP
FUeVVS70ySjnt7x8m0NjRJPR5c+gegZjzNGMRBON4QKwePwO6ltueBHttbcafbyM
Xqn9zTuVccfRYqFzevnn6veGVcLWnTTiH/cs5OdbAeHcLs5WHDo/5ON/YtQ5BGwx
VbqEr+FZ7nJIyqPyJaYtuGOOeYUOqwFCzS2ES8YJm97MzbUfK05J1voc+rdrHRrL
x00wWsLbNeEbosFT0i5jRTg9P0f7Ef/l3GFEoIA4Y4my6mNQLTBBiaVJ/SmsZWxE
BK0+szhBvdMLBIfOrqYv0HksPcqypn1wg7GOuKtYWXPF+wfikrf2d6SDkwCCpFQr
DMDYtr93uFLSMC7652WZ/dEwWT6N/NgyAVyFr9/QQSx2fOuH8hudF06riCycBHkM
gMg6EvfZRULlRSECB9rQS/zhJlNuzZh+DyXWGKWX+mBLtWuQTeqpSxYAUNIsEki4
fTosutau4n5xBAP+fu4GXe9VJs705m7DBMN5sY/rwNZI/It+BOVTqvQJLsQqr4gm
VxDXvzlIA5DGvIFeQFjYbRbyDBKyPt+4bDRT6PtJ98nmvh5CdFV3114T4e8UB/zS
DbmUib2h3XAUzKq9MVvusZqdEUlUWJvItdaS4ep+llfzTaUmKkvaGh9ZX1q0Yz9h
dHO6JDuGdyN3LorL0ayXNQulJu+hzwcZr1plpVE3XQkSBUN1i/ft9o0pPqXt53go
jCe07NFbsJHbpsS89n6A/yunmFVIQAGZK0HHI3P+Ey2O4nsyxKL/tiRzYztE7kaN
FoQvzW4IgnLjtLSWMMNHs2R3u2pTcFnrEwE/pxqN4pTDpdWw03mtuZvyggPgg35J
KZWGgBhhvHJHLB01j3lc2c3YlyaLC/XSImqmprIuvZ07VhnhqoxbhtIxszxLYu3A
LSyAI4Llki9wSBFwvKynyG6qJqKKhY1vMFxsV6MKwnQlr9dSGAoQebjxEIYm5T9g
DmRiEtmFQbnD6I4tqcL1Do0P1mokpYSW2vIPo7xnKoq/FWbupF+myThYpL83KKJV
k1Hr5r7qg5sN+s8PHw5Oi4MADX9XQ5jNEHrEP0fJT8/l4ELIhzCBIZC84CsKLZ+j
z40NvLuL629Lb+fygXmEaftXP/AGd6tYpkrOEA70jkDUl0pG1ZCfhDRcCyOKJidL
qV3XptSrGfrK8LtbFkDnqfAZkrfG/TNtDBLIHHrz2Iy/SLiF3KmFoo49JAb+CDb8
dqSByWUgJd8y6VsprXk6sfB/KETWfAeqUO6BF8K3hVFcyfSV70yaaAdRENzJyTI5
BfQQPFVENOGG40o+i7Z3/N12ijadZSA3r1wuEA6D/weDId/N+lyt6hRi5JpX8kV9
nR37JoDv+C+ADRYS+lx8FxP2SpN0tOZVtyoQ6QRm1o2Wxxt8lNwYG+Ozmds20nVO
/UVFfdttI3nNdHq0VKiPDbB2FdkY3pN/OGT0OcxGuvBg+3KIdMkYfzluUksAcx+I
q2LVfckX+ku1jgsvF59Q84x5QZxUvyos35JIlmKXf7+aHucfKoUj0uPUmFMLopbK
SJLwAUTzgAAcYtNem/KP+vNgUYMFMrwZSQcVpqYZwlMnvWMLm2JSb0/n9rZPCOyQ
v18dawsztz4X86EIDYhkGbn1ARQqLsdpuKYuY12hUCkN+P0nLepCVh4ZgCvypMoa
GC/7liA0rM6Qgo8KM4jSC0/GA51tI80WVjzZ2DBUuIiidtYbb4gXNvsu6bkkL9QX
VxzeMAma0EgqYKxkdh4YnYscAhoPQPH9jeai7Df6Zjo5cipltbMbOmMkoUNmGgGE
/Mls0+AOCEiuIiZbOe7i894Q+OB93+zKh46VAOPWegx3dC70Np2MPnARbe9e2gpA
qUxNhGcF41X0GpNXkoOLWDmRes+UIOSChMQfyJUaa/U9N29vRzH2MmiIaYNmrmW4
Xd7M+ADkZw0Z10FPizZ1hQNPTRNgnJDYa5azD/qs87vkexaBl9Gy1wlJYWZJzhD8
tV2oNxNLF6LLIL9goX+dLMCKTPrn9IDeDfGgmGETYJhzOk/3/j23YRrk0M7B0PRI
0AEpJYsRD49qXsTBZYiQS1z9k9UY160NfNYkykO4OcNmXvhq+n7nHmUEfeRxmI1k
upo4BkrZnP9paugMTzyh3jt2gRkDByaq5hYm2VBAVSMGGvKTMZOQYthDqCZddLnf
Wg92n2scLQx4OXRvD24OAh2KbpE606iEi47CH9t1B3NjBKchYl4bkm/3W/Ee0ppM
qZpmodMOUeBsYI8d9Myb0OpCAc9XOEZAHy5vZvkCPI6KFSCYXKqo7dAJ/5PJEJ4+
Phyfbd6rRlFhXkUVdIJ9aBJ1gIauWG8gE1Cp+lfS60GEhVGdQM8L1+U+8yciqePi
FFRE6OaM7x24M4JmJuVf8fubVSKVx3mIuNQdUT4id7RhRB0ICOo4SR6dM3Eo28KN
YdtUpruVEEsDjVKj9TqxASUgzxUOu1wl+nvJRK+5hMasqsufAgn2uz9dVjCNHDFO
SEXl1n5kXMVyA04THoI82ic/kw685ngU9rfS6Ptfvc46725XWFuat7VyxbN6Inhg
739G5F5EIbr3oXNK1N9u0dRkm5sM7d6OAXywIe3Luoms4wdr08NgEV7xerAQq0Er
zY7SJj3YQMjf+c9rN+C3x3cMY2ioZkocIX32bKITZg8YRb5tbteJm2+Hkul4LKNg
Gi4iO90Goizs2Imtm2uPDrjUTCz3q5GXptr3xsMnpnp7zhdHlCz6NNIYfsB+jW7m
tRpTCdT9Cy/FVcF4TWQYCb5w7lrYYNidjtMuF8+FBb8XYhHzMqJmcT2FldL00Rtm
QyZ/FS/yiKXdu2ktL3fV0H2OCruuF00XhViunTMTGbSQ0nBlg/1v/fEPC8q53jP/
+TVYcuo+c0ZnGtMybKsHdLP3rNwt4cnATT+zjenGJ150co8tks6xcTPjA0me2A4S
ORhY4x/H72gVq/UAXTbv07lFBmTAX4GVR2iUKdPtXCZH4UGsTo/EicxEqsXhCRVO
85GZCMam8ASaqH4t36pJeFvDPF8c2O0rL8jcnS7xQDEb3Ow+QzioePKRD5IhqmbC
bsFiwTzSNKpTuy5zWtht/v5oTaFPJNra667X53PhY97GD/YDBZTfcoqty+EArKFc
frF3/8Hvpkb0fsZLgsFy4ZuN887nEKzTKVJTzshzek6TfPI6hGPIIDTe2FKrdH7/
paLU2DUd9FiU56tyXjGWswFgCWSGPMSQJHp9jSuZfRLDTrh4XjBnJzdr0uuL0axP
is9PvmEpFEky30kB8I85c5zQ7Y36cMrBAtCUbt2fzONqNmVmWMjWi+9ohRvKqH+H
4hg2+sXYKDKxd44HcfSI/MDDgHm6//XTwxN/x2O+ePtFkXxutk7ZmAfllsBc2et6
n2f8CEJRcnJk2updaQBPzpwN/Eomevj2nLF2TDIY+ATg8CPZOeDegG7kTHIw/HBU
31EEefX2q0PfQhUlCBLACqjdExbpALDIE30l2ZOywH4PoykF1cczIYueFNgD7gjk
5AFhggkC09DysZprZNVxCmVNZViNb8Dbow/MRZ80er7b6Me4Co8aQ/OBrcSIFw/5
w4uVtNpE4a7hDR6F3XKKEdcAPjVux1uZBNjEKQNJkhs7iOQODQI7m23roosXu6Lx
/nLupll4Jun6knq4CyRlk2Slp2RPHpCGIHdYFMywoOpZ8k3nNuOsI9Ht5oOGGJZE
bZAfXNwSGOx6T/4XB/PABDo5EZtvR3rPLLrGLrzYQo0G2+mhh4ZhRHVj0Kt8Euno
EOgxglhUEQ/eoXhCe3LAYYj3jD0v3R1ugJYIqrL4uSYkyvzIeGTdn1uKQJ8Kxn62
odcpwqrW/lb9xM47zbNINAAvZ5XfsGLsm/yR14R1TeB0GoqxewwjI39nw+Ur5VFW
Qb4wImsKc8e8WUPx4+JbUGqPv9ITjf3PAi7drH6II4z9lGBMmfFXzMQDUNsb4Kh/
rnljS6l6S8FI3aN0mwU6t3vqipMEGbAYfsBl8+JH6DUF6qUme4IWgPkW4Pmj+YOq
Cx7x5z7Epq2ViDBC7Ay5vR8PUw1avuOde3KkzQQI4RImf9+NqJf7MpdhbfM+MHb7
fvR5y068LOGiCU+hLOWTYEh4mywQW/ic+5f+S8jcfarFPLuiljCLNkGnIvrIoAqs
iI0Z3XQQu5BAPFMySRISWPYPZHYaRzRL4OMBFMfXqNqOj2MWC9+vyKcXaS5JGKn2
V0XRfU6j3+Q5aiWO5vn1DQEZESCuQWTbKZsdTk7rc72AJ9cuIPnAaA2gvgA9fApq
NkTDIc6qQhJJ+b4840DVehZIsb3NFzGJnR2Qo+tU/YBM/JZ8LvU0q2UwQ4tSEd/N
9J+QCvMSSMWKunexPWqcWG/2C/988as/CFraHbNVFiy4/sdY/5JbOk/EItJ9/bsN
JS5wfvuVRnLMYjueSZWtyaNSGRwymqEhyBPZ1oTOqkI97KHTExywI+Z3Ppmbhwrf
yXWNVYQvfN6xLs5itI2SmTWxynb/d+bmtrKdxk4a7K0NW7StF3VtRXak5vy6fvpE
5A8pLLHOCZDdTObvUvJs4TSk+y7iuX4oGRpdGfBTeuCcxjbM86ujr4ujx63AShiS
5CD25G7zcSdEBztyais1PV9cbqRiPNb9Nd89AkYEVtED3cdItqpl58eiuXsHn6rQ
93b41CUYISGVzJoJaBCXA6WaGKwxzcxttBqFnKPxqGy3+nmy5vKzhALdNiSMRwuV
/0BPzHzV7f9olebSolMmt3cnGL4cJPEtwZmJxrHt5n6jTaoCKqs/KokrqUtNhXgq
yS6iFs0AoA9NErjjdYk1jRPdEqFf070HQnaSxLIdBFNuT3BGtvp3wsywlaHiVawg
/mEQ6er4eTjAan4QlvvF0ytpMpV7ZfpKb1OojYAzia6yZ2dJZyzAEFe+kfkCRDdm
F6lpnPOwHyIDqdHPAPiGZWkZ+rVec3T13SjZV8MjT5BL0yzfwcFBhk+y3fzhwwbh
ZVDMVtsauvSA+PuRSGw3nwkK5aRQjkpqCQfAxjvrg1cbvCwt35r/ScS0PVhUQyhj
VqOQpq0+uVlUysiYDk6uGi/khgwYHgQ1MKDub0puCgXrdhWWcQC/H6ETxxdQhprQ
huBxm2N9IOf/kOT9bMgwlpeeomcoTK4R23ZxK+2IgZRUhSCn5J5GXX11jpnKv933
11Z+c84NI9UPxo2qr0AV7G6cVMI3gvxqsc4oiUxWKJvrSq0g8G2IGUu9g4yE0ix9
nfnAX2a3Fr5XNgiC6zYJY7ScBzoDGIlZPVz6T1ljkFoPm/haiOeQlBPLLwrbDs5I
fwzdYuKYQPHnSl6I0o6Jkl5kvTr86nfJD9YtSdpq/c4nYi0+myt3rs7Q7R+fxLRd
uTC/aKwTAH/GLgGYRy/stkHkQEvmyhPguxVGIpWX2jLeJmWIvrgFbemYikQEQYgn
CzEUZ1fM/VV1WwUlfToIbZS0C7qFwKM/KIsBhxRcm+WTWWHv+sjF+B/vHgeIuuVB
aOxa/ea0zOGo5qaEotPgkI7bCngLrw4txTlP0Z2rv640jGqJIwdDMISu1SE0tk8H
nhKmxnDvGDc7jhdmL0t12oLbUKcXSXpFakEwDgGdElyt9IkZN1YOcSMq8fUXx2Lu
cxw9p3PWpn82uiVFx/Edm781/GJKBew/KYVA+aEjb/TerVrni3mYcUm1xaNmj0Zu
GL5fvsFbvpdFRcKSbTkG60lTP5AntzT0kzGtZ0STOIsQn0ZSBCOy3mnjobl4pRMw
NI0fVM8PqPGyfwjMvH4vpZFwKq8UjPCAH/1IzX3bF5/aZ1sZX1K/gkxPPb57P5tC
F15zbJNqB4qpf+VYD4BhPGnppYEipFP2Mdcm7SVT/ZG5UXGPeJIF7v6QqKEUjJ2L
sqTl5RD8AYR4I+feODJwC2pzlv56l7ivurriQV5hH5q5FZNqJpIUAPJrhSzIxZXh
1VjcYzkUMVlMBzNRYUnJvKq6Y9RcWmUJPzZdwsPG3rg+havL10bxxI7xoiQZglsC
i7Qrw/fHPuP42dqAhEB7ljcJ2TIjv6z//apqUr+fn4zun4c6oCN5v/fWbTj63AnS
xP3zyJw/Mhh5n9w/sqa4J6yQseC+s6LNoMp2M7O9CH8EbfrMXn641uXRrPfZopHj
s1zrtHimHNbod5Kf4C/0RWaRHeKgkMxOMA1RdBLL7061FpdlwvkzwkZ/EmETmKTp
zQ2jZkEqYzdoQz5v0r/be8pJ8RQg4OUSr77gjV27g/mIpelWPsWpIQA6mXFTgqqv
CAZuZx/H+fN0Fhu1iM0yj+0+itPgNriSxgCnKTzi4TS1+J+D7zprsl+Ivfmk+lZv
0SgFFSdIJ7/jFyNQHxWhlq3AjGeacIMTngzPtU+Zuzu7z0NjN6PLeT7uzABkmi84
rMXFF69/wUW2pekkxqwS8t0wMGjsPGf80KwKl63Oix6PkOzwaVfVGsBFxmolIf0A
ne5k39YiuVY/P7USoh2hoyUFMinofZQ+C+yG/ybcNrMWWzEljHcPeQc8mYN1hsji
dY9KMFlBubPufAs94UwyKqFLxH1yoHESJNxGn7BBcyU6u/BNftLN2Q/OJ50Lu2vw
rUiQL+LZ/+ck2w3891PLwtIkeRQVwn6ntTyEmVXkNqU2OnLzhv9nslOUP8ylNAJd
W0nmgJsh6X/BCAj0ZOCMfz6WgxLLNBCQLLMhcCaBxKGh/OFQe8BLMmhHYdOTERsj
hGoQXofQLx10avUtlb0Cz3WClhm4nDVzlBscgEvp1hu+pYK5N7gIPwEkR7h4bUHy
2AMY/DzrY28fliHETrnpVS3JEzfWXeB6CcxzSW94GDEj33JWMH/MnQVUikenmRVm
HfILyWso0XyT8FusV/WGunO/SKwjZbFTyzG+JsWaoqyZUMEsAIjCMzMXCR3NrU4B
lOsygb3UIrJumR/CzDtjBitt3s45S0Lr0YJWIjl+mSd1LAL3zH986r37YoeAcekd
972Edmk5bJ3ZRGJlKiBdt72DXoHY47ddPXJDIk7mdiULWnzOI1mZBF0Glfc3jYpn
diNBUEzunEmOb77roI/gk1ny7Ju5MfthHzW66BGDjSCBv+CLgdz1Hppzntgdi7Sv
Cwkapx7nsno1y9czSgwFlOjcq9L9do2vUJBB1XY99Phe4UqUQp37StXzv5P/lp0d
o6mrl6nYYccP1AooiW5nnAZhcsmC1uuy8Jrmo0yPyHrlZsi6n4YH5u7DoasmqNzu
hQkBLbSZX+Nhp4Yq5pneGjVAKDFVbECjLx2ZDq46qqNQyp2jQYg7bYon5oDDaZH9
uF5pifkCWigdG1ScknjA7UwFf8bdP/ZTXI9dziP3PvpCiGehiVSLzk/kPPJ6oTzn
jJNEiMlZvzlmtmN4OkHxl2Q/uKgTKM9ZkrFT8/ZV+2wcMPsiKUKc5i1kXbiTGAxi
gQGQWu6feQyjadDJ7KSbMdgDqSJwk80yZEYqCEDGOpgxENw6wex5SA3w6iS4ImCj
ge8kdud4nmrfpd/dNI5PtcdXa90a0PBSUEq6d/nPx3+Hfj7xPPKRo6hoWprm9MOh
8L30B/+xX51lvdlPYNN8uRYyjQTmCmAATJBjy3ZtCX70RRSoHqQPXq9MS5jCha6+
D9GEQiFiRXvk1cj+0ZPZXSn55vtrr8/Zn+fXWVwKxUj1wfF4DnCxQgxj3ge6yCai
nkKTT3G8hxh08r+o2dqGkyBVvEM9pBLzHVpRLBHoEfwFLx/NbNOnVco9F7ENe3Y6
nLHlee+/3iQOXKixm3PmMwaELYM1OJxnU5mgcuV2oJoerW5vLjQQmeA6wFtwLnVD
cd43JYWHf81PTaTKTiqmVWqw781UK6QRK2Q6fSTU4MfmL4qgRujKBCydh8AaUlPY
84pWAeogw6cyM6LtTX1nAcf6NGmfzrPKjgEUWogKL3ExiE090S5f7WqQzjFKYOC+
VTKkZ5KcgM5WfIbYsLgnVpx/NXy45yuGKu84MS8+TnGxAq+NIGc/J3DE04yvLlnU
dhTwBFJoyf2YEy+YHLT9KIzmpnhJIzhIFfJ4voghQ7mN2Zwt2tIEGdmJ0Ux4MMYd
f0WJmGO2yySvV84D2ujV8uLyXinI2Tbl12r5DowXN6ffL/l40/Q8KD4xUEdsUsn0
k4vb/BxsM45meDreV/yhcjB3wy7vcy/J77fHB1wksmoHbNWKg+eSNJvy+BizTOkq
GVjI9dcFQf9fwdStVrVZBvXgvtjtawaZkQWiApnQaNyZBc3IK7OkpY2PnNvwIaPL
KHQge4DbBeRXmesdDIeEA46ztCFpPI9rL1OGumBLK/ynHtDwDJu/HGpW/DgzAwHF
l/MViOe9jvgS5RNK3TAUn2uT3Lo39HwPT5pten/9qyR/6zb4gNc+OSellMgiZha2
YMocKiLOXgJEu52lPkoXcpv4job8209ifxk2ST1OtNm8cMWMuxJKtB/2mVo3+AQi
X53tghJG3frGyV4H4p8N15IHUWQNX4BjfODQytczTA7jflahm2flM+1GaKM37uf8
aGJ5BuKrgU0HKuHlfuLBGI4qZ1ILqRA4RX+u8osJUWau+ZhQehlF7dvMvxW4yaAE
oge8JiFFOOsnAM5P8RJwet1dgtT1Aw8XHCIMB+Qb8qpAJJS6EIPm/gMa4JoRcuTf
pnLFmV/OlwDY0VqpbVYP9CWWUY/IIgL/qUT3xcT2yVS0eZZBPnSgpF6eRjaoktFp
55C3IK7UOlpAtTgEcsx7yqa5WZiMceLTIEaeNRwOsUjNBTLN1IBkEG1G2VXJOZXI
DmjwUcPVvZpGGgJOpjPpx5ucgqafJzeAaLryGio6KcifCbWfdyfz/YIkgmN1g7Ap
Q5+U/bJOcsnStMscYXz9ULAV37j0tYPDznyPo3CL3gcMN2mBxZQ7dcP/2nVgl6I2
ECxYUltFM4JUBybaWp5J9j0WLrK9kUONoyjqy8KP6u6JRpwPXA+CmuI9pGAphwnS
md9XpsrmL8t6jhjKidyYdcWf3+HnTdKaBm8YcTLDAmDVlCj7aziotR8JGXFf6Vbi
IFuUlN0bmSGUXeqCEEVey9g3IfpjwUM1v8BD5ictNz30wi/FSs5sRxekCcjvf6zR
ilSIz1i2W4Xj9xjVYi0OkkCeDGNuEQKfuXhnx3fP+ZxKA2xel+sgTilzMCMH1mhy
8EMxE8AXkpOfnQSwH/Lfx42LFfbeiPYZ3k7n/zHdzAjlLCwH3Cw2BjI8Ct3I1Ff/
n5IrZYzYEhL+hdh9kdczYRq5XrkX2ZkxTSGVxtTphVWN/BRSl4vgTLrkZZlT0oHB
xcscbzzuUGW3lkEbzzftMVov9gA9LEr/f2Q2BGr52/1bgEOvWoKE0uOyCe5SI25j
C9gtw6yrmnpdBxZqzbjCsfCGTG1wOz0TOeykzHWPOuE79GnqxK8YQe8+sPx/Bdll
QIBDiQobJWio4tbcXJp3Itz9cAmdE+aZXUP8i4Y8G7cNg9RvKjzaR6aVEy8xXVl2
udyx+Ef/dsSoZ7D1V6Hm0pcwYsyzyqCtMzyFmvFiR/Szd8rFZqhCwJN51ghZXi//
lJ98SgDag6op7YR4Lezs14WMAza1fO6gb+WGYK0r8KLqr7a9uITv86ga0pcpa6qn
aRSr9j6oW0h81qqrXAMYuq6Sv1LLoaV54EXDdH0fYHibYspCeXH8UIXMb4t0x/LA
U7SRkVjtoCfm8ouvWuPXPXS61UejSMJ+qiQsGdu/WQmE5Um5N9lFlotARnzRjGoA
FePNqBbjNEkjePibbRM5A1IBJfikp6Jg9Eb9obogbbcbYdMzYJOrOxRVJv1yCsBa
RBshyAraWEcVgM35Gjt3WnlUCK8VoNnCm8WctBLcMleBdYGkhYhG6jliHRBdmbun
DfM2KXPkmNpKA5MWkIn3anWHodiaCrzPinTnhuSUD5m0XNVg0yc3cOBpHi47lBF2
HO1A8K74am1Bz9M9pATdKyWXoiuT6okAUvVNocxmYez5hIG28aBcgL3DwZdIi5tb
5zn4Wvuj6SAH60UERiCh2Z3jAkKS56M9HzQYyj9ZhaQTBmaya9o+1Ba932fSPl7d
lPg7RzHZj5lPSGbGK/iRjHwK7OhaETIK0flIYrzlenc1dXeXZFo8wtI2Z9PUeUhc
wAudzGlHD4TXTd1BiBY6ChuBiAkE7n+jix+s8If1EAX+n3nGjH0RTcqb5bWn5eJC
2yMU2HzlYB+ZojH0DwNiIv1ycM9H68QmtPbrmx8xEjteP5UnTepStTx3nSMcMPGh
rnetIem1uUJEY+z8ol5FBIVzqUMgE21apWK71stEAvpUubhCSi1M6ho3r4j7/I16
romUKNJvkuCNtWefteY36C5yWU0CziwjBv5QQmbnKP+d0Ttbuybtq44hm9onKBQX
skwzaM/8IOXJvcGLuZOKDiEJwi9qaHpOJaegixDV5qUWicDtAWdVvtdxmPPbbEIq
Ptp9hsptvKXMv9hvuGosKqrbHyo8Y99llEzqmlZDvPWa5ZxyYfb36JpnOr66l0r2
usfT0+GIFLrHYE8F6d9U1M+3XYYQzwgdAjFlsADxhmSUar1oDMz8lt9l061KU2Y9
ec/pCiiht3RJ8hBUEaUT2iwgP1E3rTsY4yFOqPkjymE/OBxwoygTPl9WN3j4N3rx
vfPp0M4V0XTeo0GsHTcT/TbBilzm2u4Zivr05I2pqUvDVd8ggR81IyYHGI5i4zg5
32FkjPc3Z68HR4Kc1oLa8Rj+YuWHhjHQgp6C1wghTCdpQqsOD1qOonEYtzIoxX4I
2eUcpaDV/IihiLIUQrIo43TD41tgW1e+F0lQp7L76Q1VOsLlZWyzrIj4k2JGHg31
QC6/hu/2ug+DnfPz6RxUgJDg7Wm0koVyIaU3cHreF2yVUkmIsQ6QXaGMLIYR/bYe
+1QGtrR8OhO9gAvzmRLIaTrYnL3ifRvAJeDwS1W5T7ay4x5/V/XelKmfls8POLix
w4+9Ig9ewtSuGYwddP5sqfdoflEBzh0hGWNOtmjvkP3C8tU6TnUWF05CXNJbKLA1
XJJ3UUaYDjj1DVM+joQX9FXUBlTeG2IQLAWflcPOj8SEdloudTftATwWF+dzRC/q
cOXDi1MweYwSfqRQZbFheyzDWdAAWyyyoWRjoXBTAKjKuD+LViubxn+mOtDRremd
bVSJnMLTAZyoxSMVb9ZqumDc+yG58k3qQs6aeK/fJUr8Qp1O5qEnw/jdQQgOsz1M
adl4uY6iCOhiWPPRJWiSmN+21Z7rIuFy+DnQvmsu0p3Va8K1tbN2JxRTstVmd4Cx
desXNmihpZnlIDsR71US9U8Sh7djcrmKTfOPxCV+HPbLMArjst1/1PkRc66Eob7p
1ASO7wFWTJ3aAKjdCtjtLYdJSf624b+bF1pwqm1Deen/cd4GC91uUcJK4MVA3WoT
HHPPbDi35DtxjBH6W2aur9C1Fj8a6wnBh7ncPDp5VhqhJH3pYsUh2vOyoB2dflir
iKEAGnsmUle31Ws0g/Fy0/Ic3bBqZJr3HQoyVHzqQxAs4yqW9rL6e0pQr+t0LMoK
7G7Yt4tvXkOAWmfqHtxs5850kRWk8wXB2tyUvFYAKvYjejgcslGEsw7aMRAwDPnt
fdYR0RNMGTGkwtlUHTN6IgVipNs7hyopQ4xnUs3jVA5U0tyxi9w6J1ABivVgJ766
Nv9CxXq9IRRTfAbiJHVhY/WOMe8s/cImdvS+QWU3AhEm/pFNHmpY6HwsDUt13gbS
am4v4X/usTCMVUzcTDG4Dt5pgEZTaSCbSH5wE+UtCsnRtphIhn+lp6KgfO9XHasH
CDIOttjWY6dCrM5vR5o4gGUeM8NrHttyYvYmofV1RqqVu+/YFNUaWF/TJw+m+3zu
tOMt1zN0YlEukZnleyJ9of9VEZWSjcKFsYMzyDDs5GwIbZKm6HHBXvrcyNzut6PJ
3anot17FgxlhpNJ6YAQemvxBUMEYHVnt5z9pw0Wkg4wdMbM7wX3vDDlnYf+3CIm7
EOXjTbD33Omc6KvE1gEgrDLgmd5NfQ5Y1YXunzMlTszcLrIrzhEPFoKvasvgVNcZ
zrLoh8id4KwDHvjmPtiFtRo5pIe9/rk7MPSqEY0IyVqnV7ZS0rrz0BLcEVnoEtHB
burorydfbk0Ho/xXoN1e48GfSpXUEUSVglv9yT+ev83JDHpe7KkUysQS02uUhNbJ
+WpYbgfXnC8jjIOt+AccPgqq9AyoWo4WZA8QqsrC73qWd+tYU+RTOwCLt/Qmqjwe
4dFDZ/ql7CEPdVWj2GiiYqE4nOiRLdQ9of5+hnbUecVJQEFmBrF7vQUxrnVkxEEJ
dG04UpDBKtr45d4p7xk4gKqSr7Chk5niGcL74fjdLJfjFQyYbwglm/+YW/k4lIOi
/JOST5jUGY20txSwZ9aVr0MK90GjqoFRDbujBfceYpKV2eF0SZyBr3KCL/pX9ikB
ABKVFYfmSSuwreUFHRZjJdWzpb4STtcxEBz+6DOwmbrAgqGU2+BuSY4vyWJN5Kry
85QVhRPfgKBQmaEhu7Z3mMdLkvMwmUEbONh98EQomEoa/1Zb1q4IqdRR8FvSDpRl
+0lKrLNJ4RoP8IwPV8R2wVeLAYEA8cG+ZBb31hNR+AbROo5TMz0My42MZUbtXSAW
s8MVPVx/s15+wOloqVLuApWoKgz6xixfBCdpBUkzi5yxVwVcvQzp94lam33R9Rso
vH6gYiXA35jv0gNtQoOTwVbAIkjkyo+NCYam5SAyLlR10OF/yKHvTNYCH0eN9Yy2
2rGWPtGQDnX/OxRmSTOi16oolkgWLJbSBq8yFp315gTywWsJHDw6sJYv4IzWvCSq
SRjObxzjA+S3bWt8xpAEen4JoXTEW3l0XIHbKUOFef5IzyDq5wXossWeJKON1yfe
J4OYOptZO5Iib3RkUu2BJuU0qlS6WD4GoUo3r+xoP3dptLBiHr23ZDNeGL2iKw8E
zUjyix09iPzxGArSzAfB4RIwwITYyL55pLDnXV5buWuGwiIXt8d/Na3TXwWfFTTz
kVljisZ/PPtwXsvcus/himyz45BMsqQ/c0QZ0K8RFVZpcJJurPDLESoGS9UpMgWh
FBcqMt0nVYauqpcxxdXgtN7/aU4GvzHIK9alZaxsFzY8QbYquKTPdZf1mlbu/e/a
+VuFFazRlM6dOvqaB24zAm4Og960jKlzAxti05JshLlSRQ3atBBTnupwkLqvBhUa
hj+c7CEqNKd0hvubrWmsp3Cj//8JbbtMdOrNMqYzAJGkB/ZVqW49jNMbhHXCUn4E
4RTH4HN46YfTJfaTgt+CM12+mndB4WvIa0wYnFFNxZd8eIwjaQpqW8NfwGuolpCf
ZCBNl3M3+ww5OsuQ4jGoaeYnWOZGyGDO6X/7gLJmNFNVjlZ3/+5F1Dyg8rfwuGkY
uGsw1IGCs3upGlmIGll5ZOnOVs6+wJzEETGQAsNdT07siBXO7V0DY4vHkXkhYkRe
7VTvVXRGWUXZYOWy6OSoWW7e/Gt1jZzou+LhGX11NpuIK8/CxLcZXP08n7mlynvl
sjaQ/BVaCMN3r47RsEgcqZBFeFuHcMNL/9VFem6aGSc266/RcljiAPoW0AnDd8ch
ucG4JnV4EOHfZCW54QU+pSt/aPXcSbW5GJhUbU1pnZuWhTUEZDy16L4ugzkc7y6q
gWddlaQx+WifBp83lVTvNNr25EzwjZD8ftb4lnFMKsvbSqhFzpDtPqMjW0Zdr0K/
KQDwafqi4IaETUtj21Vtk61MWHWYB8GJa+nVvPJ3mgHPFr4Z5keMCyWhCdkF2Cil
NbGZE/MDff5rHCYyQg9sIUHfe0DZFGMlOx3GP8DpnZP5lcdYUklbl6wgMKxvefzT
af7l8c/8Agtbra7AsbHnREt4O6JlG0DhPLiIq+CwW79i5WsqH+hx5bq6vm8cW+LB
MRAaywfN8yghsLrLjaM/EvwqrSP7EwJIkb4i6wpUTYleZy26TZ5KqPfSlkF+Fgbd
FG5EMo7DZYWAZrpPStnhoj5r3YmpU6Fvizimyp5hq3qExqmHValODSfxD83T2p9+
zN4KOgvrRIgCqbceDrA+NEzHK2EA/6A/48sNqrnHTIxgfrXDUXjHRS8xxFEAabJq
+4dwAF6UlgjihruOveZVY0XFclZaafRZkjRtAomNWzjoli9WUhC+Zh4tJa5yI0W3
rDly+kcCqC7Ybdj/mgFqLy2lqtvQN69kZ9OASfIp8qrYkXQKrc5SLl0FAvDXihvD
9S/0uq5iHbCXIBAqvChzyogvX14NNRUGB9VjNTCmk99TKF2s7Yc7L5F4NJ9AdXep
dI9lLnpGncQE1UhgmC/tXl36vFidLoWaxtLkOzvWFO2kZhxaqkyCtDdAyxyMzQJ3
0j9f+S8fWFDcwDu5puZ+f9UqGX2puO7Fp5fN0IQLhmxzaWTYI8Eyq/FfLUB/vkr6
NLCNp8nk+5zvCokLdxuQULOsgqNvUHtTfh9eDZsb5RQ4L1nKOPRcs+LDl2xXItm7
6G9WCi8FakZi+CkVifKAgXhfM28/qIYPAf31vXWABgNSNX55kn07fKLYuIlT/fdF
JVxiL73WGqOvC0UvJuvo1Pacmb/7W4RMeeMKJFRvOgc86oVVYM1/jSaohqyeR40C
X0OSt3DPag1L97Gm0jl7IxLnUono9chB/yVQlz0xv5yRwhjFbH2vX7BkVNX1Y41D
LmL6L/r8nPWr+wCkXOgwoJtF7Z008DBHmvlPgxTMmaK5n9wMgdFx9jOSsEmhCqcv
laxrBt3Ed2HMqDDl7t9cYzlDQiT+74a+M1uIzPSJJxwcRoneLlg9arlxYa9WvKIe
UMoXNC6BQLGPDccKhaMNdPG83f68NqjqGk00u/ohpeNG8Z0lPA36sty0ve0Krt1x
qDMvpglr9fbL61F+zIP7apcl0bLvdkbK3zVKfnZBSkCuLBWNqP+XJKWCvvAKDqB/
fhy1FuVtkir9KKGq7Os4HBUaSBzjsFB5HLMbTjBsnnexuEqiqIsI2DbY7hTHtg4o
eHHGHcZeMGPeCkuMupHMcOL8DYgKPeBy60W9XCFeCX6KASJaGeXktJSa+X3b8lhv
GobfNcSoT3O7hu1aKOnCym1QbTBhooh3fFmN7Mn4jUqVWj3mahN9N6E1r+Rsh+s5
9UIrCVN/nY97D2m30gc8iBVwlfD1kn2p3WGqbNChTm7Z10PPJ0YRMEbCn/0dpZ7P
2N7NhuW5LuoHPUqIJ/9coIVAKL59dPWrWTo9SV5n8Z2I/CYN4D9pRN8yFqIlgnSM
kN9PSwzxcuiRrdc/9S0lDzR9sqUVeoQU875Beq0BCK+RDF7r9prYIp6N7YP5b6E5
SC7Af2NxDT8oYfsNzoPv2bkGbd47oEoFpkIvix0s36nlRKmbIlJs7HmRLiuidsv3
nRY+QZr8ylzWEmKzZwTWMJrdLXD3Dro+jV8j1/TPytJsyPkcv2WR5WKWYR+lzGsg
tL+tWeYnYJ1hZbcCdnpMVQC7Xz19PX5BHQulz2TLYHiinRTmDGe9WcYO7xoj5g/S
KRloUm+33OWmrPfBIV8pBCfeBCXgXg8p7ev+MyOQC58YLqccNUkTpbUr4DEK1hRh
VYrzZGFXPGD/lr4Z5qULPMu1lYRG2rXiSeFOM+ELLrqR7uDq5/jrtU7VPN6W0Gkl
H9QIGPqKcUCJj/e5cmA+rLueedUbzL5wmH4+Pi9YN7p35BumHJVR3u31EllN4+2g
CRtZq0enviH4BTIcpVlomtoxoz2cBDjMXU429zt9R+TIhhdugpuYKnbjtOZz8VhO
UazOxfgxdxfCdt4gfz2rYs+sq0CHdLQDMrmAQUML1S9KzMT/lv0W0pVNnB0egVnI
5Z20M76tOVe+YOb2VvbivfTYq6bQD3VsARg+yofquATmXMYWor/mIF4ixaqFPHkG
M8V5fKoT57hGY1tM7HrYYnl42ANlksrriClodl85skj41s8IPzx6SxEJft9DE5mH
K7QC1Buq0yCGjCXvWTwsYC0SkT7sco1764QQNUGoWyrdx+yFa7WXyab3MRT60zUR
FY75RghVct6P23bl49pR9ikWJuX1T9yAv3kCOip7V1mWMsvZH3G4vCX/SHofWtrB
X3Bkwrb5lM4gtdfz2XvzML0iTB9lVDXKRcA3UbfrHmaiY1vqAPTkNaAQrveK5FQg
RJf9Fdiltv5j3bFE1ihStLUqvkKYlJnt0CbTZuGRu7yuG4Ej003X6CgrgBt+eeyc
qJ/ylwXDqqp1OdFyt6aJvi/3Qu9wL1U2BVUul7lGAPoVyAd5xwH6zxs8BaEly9ow
9Uhts4jndmPI9b91zaLlqMAuec4efsULoS5P6jF1FUhz3/fAgCZ6JXytPqLbk+/w
3WRpZzdW1XnMmfF1miAjCuhwDFV1dBgGKC8owcSBMfhZyY7RyWF3Vy/dVusfOnG+
fm1h/RqzoY/IM53CVdyvPltgsAi4bVW+2C52hdfMuXvhUCWNBN+kDLPZRlUh//Pq
P+Z/sD1ibXkHDXLE+EAqasPbLxC8vOBK8vd/3m/dAFPXpDRyHZpaAE3Egjtj8Ksx
Dw4KdvTulndFIOk3VP+EAXueHRLDdWwCAuIgkw9UCbrRPMOvGR+v6pYrkWao2K75
DFh2KkFqb3dLFdJxyunxg4hAj6vhT29I1QG7XUuGcRW2zdKms3pTMUZx9yuTTHj0
rNOaOl52jrnCHt4iV11wM7eM3GQF3cRRjConU3IST3GAKXoDo21fHTYwLpSrDx2O
LAuiqNgTy2/i1WIK7iZQ3SKKKJY8G/R6u2uMvy6I/at1z+inzA2PXdgLsZ1H0hvV
wt8dL+VFu1Q8yv3oDCuUq/8OhA+xuh6JRYtqGXbedF/I/DjsDrfszgaknqo0IajF
WJUpvEz1zhgtUCBSy3aHfYw7B9cMiCFuqUGCBCXqqtwasrObuVmUOzgd11ArsLP3
EAaSmByvznRVAHHLdgMo5p/Pm3masQzNuZAjeVO5ykK6MvfLzUeQtQ32rxpsXqZt
8UuLI1GvDUntIozoBdK40IhBdKvLlDbHAwxcI4UiAoxnlJM+n5SkUmyMtibABC6e
klDIZnPSCYm77BMfTF5uSuwNk1jdDzEKRMffax0MXaBJmJxyXN1MjgKHUgsix8DD
QAUoJpU8UyilvHHvQ78kxIf4rsObtzq3cnaCEsDkccHVdNl38oE4z9kxF+7lUKm2
Oxq3bjPPsKiedyce5a1Yw6JjlzbMPYL9ImHCbHYTUsFdBnUSPUEWicxma513iBtc
vOAEUgMXy5WPQLPrmRH1HX75+zebobNIMlmNUw9VqVXiFAgNfWpPWP8Zy+r2j6vm
S3C8royxxZohLIMkVvMGMj+KsGDUqG7WlmpFsVlEkUbiji6xRzox8FDOR0z49EGV
D0/h0/TP9HBWHYuZezJ74X/SDpGFoxOBSfP1rHc1IAL49hSV4Ojl6MWv9AojYal7
ifLKulwgCD1jPm6tZLCnekqS8QjcpY+k0dIRpQK7eYRE0Ke911vbf+d6hM+XWojE
uVI58Uv2PdJEL3s8JTq/eeUEK9Op+Z2o51Sp66ABVDLcqYHPIBGznDj+uTpcz6F5
tHHkD9HAZCcUw0NHQthtR3ASG1DOeUJTyS3PT24GN58aZPtNhdt4TIwS1H45CG03
ABHq0SLAr349dI73V0qWzXLuJxbT5YZ9/glMrbhWVLevI/3CFb9yFjpqH02ehjwg
vLvqY/eha5r+ri2tGYYXWkkRNNGYgmcEPWwMm5pdIoorKLiigzBEk1AspF3KWiJm
rqTXDp30Gm/sIbPs34Z+894HsTD5dYMDT9g9aVC9Xri1Nhw/i6M0B2UaJ4qbXK/P
B7covEw+YHHMA972QhObn5j8/y5U61bBdh8fKkT92tp9FpYlie8MxN91LuJPuQKY
43/JN2EafkhmhKdE2730dZ628yJMklqMAaib9DAFhJ8DAX2Q9FGOtAFhfJA5+ehs
vXvhWwLh0n8H5Px49osplmLfVfbEXN2U+yTpYp6+rGFHi2hNdKMuW0MM1ClxOVwf
wHlLevHPl8jYELGLIV1A5OZWFYhuBfblI6d1pTMkYkStPjeMyRtPXUXMUCG4wiXc
v95n3Hdnv1mvmCmkksD0EJakwHD3aYKP/8kdWXNguSmynhV0/sV3zmpMA+fAP+HS
iyJpE744O2Qk4sl2GuxyWYo62nQ9cn+qqQ3IZmSOE5Wmnz5+RDq7ivxHqkPfW2TS
dd9MhZUZJM95Ron6h43eBQRhVYGZ603jGlb73utY9aN69FpqJNDXszkezf6gyrmO
nsMWbdSqQvl/S0FuqJ9F0ShbnVWwMS6IJ2NQXsDVSZivO23Jd3DKUEfDI6bp1DXI
f/qF6smsV0SQl2kH2a5B5tqjgI9a0PdxgSZGDqPxYPPBrstOH74ItdC12HvQ3S2G
7Ans4xxuET+9VDe1CPNWLlWOr3dC2Vm8bNyLNO/24+aaY1TLOo2/MvQ5g/mPkHxA
py6fJIglbBEwRoZTk/8u7vCS4k31/gjThpEtWlqSBdsQrg61NiCowL6WExMkAGKc
EmIg2RZGsg2Rz9sWCaDBOeoTCyRo1yoGX/x5w2XjDzUIKchzPZnrjuo0yt4W7qgz
+47w6YXkznLTXHHrobL6nBJ5XikSPkdxCduz4THJ+sh9PIg3E6kTGTxb0787g8pG
Qre5e1k5i5cPZMUYmlbdNanwOth711pwd2KOEV7XVvjT6+YeubouFMMOLmm8Ffi0
tbUGD5UYuKZ76c+jQnJVAORMIsVmmLsrcVG+E9Bbd539q2HxRdV8XOiJVHmdChxS
S/DxFaR/GUUZ/BoR2q1iRohzuHbnTDtWKbcILSbQW4tNpRlPM5uLsUv+LEGMxUtX
Jo/ZBl6XvoXOw7/epOprosDwXQEcsy5v6ARgi7WEFt3abAmnQfdE72lQgPYloceC
szvH2HuDhWNEy2s+XX+4sGukeSsYqUz79uZw24v7I8GrDwCvffaMGABgzerVAhNt
IHXm5z7zeyehQxOYAZBxPjNZ2bUQdNvt3/GsNBvYqdkNAh3pVcDsCJLsElec5KjY
gmEAq3LpvA/3ptj0aM3hrjyiby0FJ4xDICYos3spvOQ5k7jm58PgrLwiQpgHy9Ch
NzdaasFdtuDZWjetmFzzr67lI8i37vHcqGOq62sdYx1t152jbExcZfdXE4xeNgdT
HxfHgJHMRrggVYtPLlKZnHvJTuva9UThqVV8nL36/jhTRMZeEpfxVJS6yeZlDRcV
Bww3Wm6umLkBJIrGQ/grNgyJTDbaEzpXENxrdjsDoXEUEd5HGnXhiFA90aihbSyx
d+f7K4kma+l8u0xqx/n0dATfnvL/PTT1pAkieJPq6Jvu412ybzOlRe/WpII+hs3B
R5qfUtF0UVXdz2mE5Qpyagfc88JezIch3us+MkaG/Li7iidrpcOLM32IKXSlDf7Q
zWLGPDUGAW+tk1epkCj9LgkNqFvBHf2JSHhmB4pLSvK6wAwErVlo2tpmGGhHbm0e
AkFyFyqipLKsNE02cz6rZAWckESYrHS5TWKoqxOdq24tneTDuv5kKoVYsRQNWImr
mamp4gc5+BQcd1cWR5yZ6gbDbIsOIIhPyjOx6D/XcaGEWjRv5Sih9hbZvvLd+gji
+R+EdMgNqlJX7ldSBdegrxY5AcbSQByiNwqABB+CbUSAvxMt/pPBuzBB9oFaG7qr
2YSmg1qECTpLb0JBlHxiLksyU1AB7QM/2MzukxxU+J1uxqSTFUaYRUqqj+6p1vc+
ukyplZrVu7FwKWf8SZI2f5SLQ4eVBHNkrPmxeLTrRDorln+ZT4FbwmyXc2roMAQp
Fh9kmCaH5hi/9NhfVnaSAlvuzS26ztxjvSjqv36EHdkmSPO0htKFKyHm/LqtCDEF
n7Vcgm9iuJtxC9IAVCHziroOo70owjUSIaI8ADDOCwvA/7zwx3vrK7GtReBptAQ4
KqQ9puxOebfrMxlCUju2IfDuIGu7POgtOqjNCo4B+GTXkhh5r7DlzhQGduKsgUgj
KkcWaaAUk7NHGk1lBRvbLL80YLMD3BASsuQo6wHIBptdtUT8K2oiwn8Snq8EneV/
VJETCg5QoOXikKRDixVj2ZhKc7YLkAWE6ofOKW5g+g206Ku2iE5KM3k3MdgzoIX8
XaSyZ0S/MvD3qTTt+AC5MeNhbWziBbCCKWcFVIOjp8eEXx4cxu0MCWdJIiKPeTs7
nPlItPXF/7RrT4Y2Z5VLACyAuXCXehRT7YCJfzWG4zx4joUdQP3++xuwml7zfs3r
BXyMP0imGytUx2lNe5HE/mpBMy05AZw+qj0dbITUxt/sXg1dWAwJYzf/Omm/fbZU
wbW2eN7yXRcGhXlu0HDL0HlSC2XBLMGPiNGb+GWoIXKMzN5/OQK1Hjtria8UTAOj
tV6XAWIqlAftnWo2C6c9B8ShRmN0k4nxHETH8YJSWpL5Ft37/rEEMSCvKsfHZlpk
rrvPjhEV7qZ1ZiyU8MIlsPz0mkDH4OfAmCeyiNs93wpKnMO5EikzowK6p23Kh+fK
GAN0Q5koT7yCBRTBrBHKJgfaLrGDTZfOCXIUQDle+O1YDkJ2vLxYW4cZyp/urnBh
iblUPbV/YX5zYnmYDGBN04UA4JcHxfxdkjzfETrlNZJMVRoWECBUXXR2659IdNEj
4O6AXdiWNw0Kaqj9dqUxPCb5nGg1IXfPsa8pRTvsxozcx0H9k6BPwjLcX8BzROHJ
rmDrQpj0UVh2TAx2dd4m8mxxeazuJfI7vTSzQz1WvHc1fRBRe2JW9z7KPhiK2xRw
cvL7e10lgNHxBKcTIg6pgAolJIarpMNDcbUZioZfl087VllNOwHc6YGhapPsS4YI
rgBO/kWLsxzHL9k471nOpGYXvin1UuA87q8muglTIVUXKUcvBNg+v79mykT364vv
Acfii6oe5qVQB8JtJ9DGmninH+hU3W5FouXpfofivrze14UyHsIXfU9G2Phhiu1Q
TBasQmMdwZjpO0yi37KaMB1m0TlyGT4EdNgw2q70bVnX2ii9qGCikXC3NJZKt/io
sBbY4hUX1VQtRAgIUkfFVYJ7PPQ2qYktMy0NeQOrxk9GZeZclgeblZBhGnfujEYb
zZBC3zEcI9Vl5JlUU3rN7MqBhkILXtlSiwIig+O28Z24ysD8D/sILLrsRWnmfBxT
gxCgxBEb0MUVfmGNcIIsykHf6VPWbXknAuZh6Urji4cgIAgTSkqzM2bBjluziPv9
Wet1Vo/c7t1IAh9H9yuSewDU7EI4MdfQ8XGfFzFyiW1cuQBviD2nJ6rmDEsmbctK
U1pGaFrOER+iZ78ts8eARGS1EWAMK5FjJuw9SVh8t9+Yq3CgYVX5CtaxSZdssbPy
8S3zcFGjELP1yGiJMHUXknRdo55AHx/DmKzplMhPL+m6OMNv9QOEYB1TG9jsmopl
zKF6Qd6IbA7jVmQ646SK7PpE5Nsb8LmOoLBet75Xb19tUHWBgun5fFsj/gOYibaE
yvMcyYcGvFxK336qQtnx75UJCwgVr2cdkFiprxRzBekPtkT7XdfFcxO4f4KsJH9R
QvN1n7JL7b1B4eDNMTuplJumpq7qrkotsKpqJFA5aZERAOoIc+mtC+o08EAN8vZJ
galZZaMPX5gPPh0muLT33jIUp6x3YN6qmORlmxTgtrmzXpllUPX+MOkgT8L0zBSN
/0mYwGwOxmvz+d4IWyPJappkSK3PJISGEudwzJOIeEZ0WepyH/HBRS31+4k3Va2u
v3xj+O4L+M3el2vAvSPezWUM7l4xI6O1BIo/RU4rfvczOxx3+cHA0thajG1PSu+m
01MUSy5pR34ZOEY7g9dZsHccSBFyGEsTaJCsh7CQwdn5nn9Q8nQ3c6BkaEz57zCZ
AFqoMULWY9506PQnBbbsj2PIduSj+G9NtV0rR88ESdyqn8GARxabwnlJ4DK0c1PW
MZIHEh0sUpxIE1gINouuNTHLCpaDPaMxJonTVADdTPPRFSOGQ6BEuQWDbGrWyGid
pQv0VElBvHxY+5kgCQiNvBad2zo8oON/JFDHfy3EnAprItNhp2fip4+zipLHn5of
6kUP8O7FCDbt4+v9B0SY3Wn1P0a+QGKENe3t2WoT8IjIZ2aDMFphQTu1cVH00L6p
qya2875cGjHk7Cgohht8ZWbeHcOilhNA0VsCW0faslD6POpK2hKwnvsJwykZ9Hfj
IwF4U9hPj37OPo69xr3Eijvd9QnDkW0hElZ00ed0XxqSFrq2ecjSj2HMXhH9cUZ0
nGma/kpddK+Btg/vFKGuE6X5JCSw+IS5gKvvOdyjB8PWKse1xCI6gF50A7qgU9Au
dQ8zo+DFZbje2jwxmzFLrbnC/bbRPUq0T2l8/CULRrkeyv14Wz+uVXEEetdAWDoV
ood51Biy0+JAfO1s+8u6K0mOtSlP1xbIxsHKIYrRiYoGboVM71U2MmXUI/+no4kX
SYzn+xjK6VzGezTNhKWcGep4jjPctC7+0kaQ6rmCAShWtH70hEGFUjVy/PHHUcZC
QSYhAmH/V3lrmHCWSL/cFtZA38Yh9TtDH0LrLkcooygtZrc1OxS0AcPB3qzY9wrf
5YzgT0USt22PhYV04NUVfGevRY/eT0hmKWAm/DPKk3j4haFKJtLn9nrhTV1P/gzp
+ScmUBsLbv6u2OLD6lcEm4QWJA93ukrkpTFHlBl2Eu62V0DdF9ETtfE3+88pEF6t
7cLOGxGOTNmamNDWXRNpqLbP4qMzAKwzJ/wNGDaYsoOQfy5f5h6fcLTNCopd8R5b
wga/kk9da1HVlPn8ErYLfcqXS1f8c/B4G6AlVnwv2KxfLH8dYmsVTYqCnmeM2Yir
8/psVaJdXBcvrR6Yh1ZgxZv46f9LEoxUnBgVDaFxUM/3T8BSq8ETtOmK2OHzcBA6
vya8QDG/OTsxk2mp1KcIH4dmY6NKnGxkbOmBsO4AnW+Jmr8jJD1mT6ILjonHlnyl
C0dtldG5i5DjY743nH2grQ5xexJrO9FJXk00o0HxrYp2Kh2tgV3EWCQqeK+5zxAq
wAkl258EHDLA/ADJC1HaTfqmeeufiJPUutrOxSaI/B/1DMjXPyk2PAZIeyPnYQzR
nsdQFQJXBVfygjWXvTWgzl7e5Tsey6nc1K+vqc1G/p/Fb/KOrwVcl/UoALfjfYYk
FjN1co4kwyT34HR3xwx1Pi7FZSnc4dunEPPavOyfoSlc4fRJkMq7roMFVFZBbnPU
/v6HD9t0QUKb15Ryh5HFoGFA5AGpts6EDu+iJtRJFMWaEdCFbmSHj+N1wMP0FYaH
BK9Nm/Wl6AeSnICD8THT4dEQC5Zg9o765r5X12kB2yivbkhcLDE0KLKSkohEn15L
cRpDOE/WrRiIs/QyZSY93v3yx3sBnDlsKyhxyMfB4cQqPUUHee5rVhWP9P/JOJmn
ffVY3jGV6+u8cu4FSNwIrENqc0HsUQOL/dTaqOHBJMHxJ5rEdyMj3dA/r3TdLbpz
5z1Lje+nSsssODBOV9znrOmwNGF0Pj7WWs63kKadzQHdfu4jprNxfyrjceKabwWP
gdnAZSwjgUzuzAZ+aFzX4gABBa8q6wk67mhvqODVHyU6TCNkFI60PVNaRkg+jOWg
y1fhvhqE/fyRHNzEQ7W/nAoSZiK9Awk4YGCfkpj1gMcSSaubSrhDvh8zPQVAcmHA
jsaSeLiJjwPUs6kXwFtTOgVH/S8bDxPQ6uesk1sW1YBBQddVU4dgbP6DbKnoGUD0
dylEX4a1XtNCvDXBjq2lhHgm6uZyuGMFItGn2ayt7JyTiIyBeJg7Z6GRJf+id092
qnp4rx13fnhlY6GgZCb+oundPCLa5XmX/CfUkIcuXGDls4x3DM03ldcT/0Qnk1FU
ndU+VPbVfjHJs0A7FSqq3dCYSgR44XHnR9rKC9PDUVEyB2dyhYiSvvtt19keww8e
C5Ta4IEaHc3zSbKHaaN7FaEspyiPdhwrZVFq5t/TVHz3dsdgJXFemeAL+EzgN6LP
E5cYykdoRP6+VEXqMa0GMcjH8jdnBqIP5e2yDamP9SyLNT5BBL/La2H74nZdhRIi
xfF/Q9xEFLZprCZ5xh4WzIDGzKQSKniHDxBHaEPTfAmPdULqUefmLvVFNvmeI/lu
ohxpSFYfbMWhn4xAY+17BQLWARmjR1YZO/bqJZ7FFDe5ySkYsFsD4YbR6y9F3gmq
V32LUCtDzCwlNvQydecwkXQ3isvLznPG3E13Kb2Tc+AaH7jw9ZQWXTO57OFWm92o
k51NJS2Yk6X789ktSwL8LatkbCAQ78GhmlcOBfh7aI3UXCZcMoXwSn2SM5avyIx+
hHUsJkdhj77W3UkJ5BiLyz0kVV7KIkVtgRMVApAIo6modZt+VMlwYlTZW89zyGGv
/PW1anzbJgNnRB5JwhE3K1oDxH0r5A/cQ4IHOhEdbq4PdCAVcNBzRuAVaHwKcUfX
++jYXT8sRGHsF0Vs9B9P6D3/OeeChbKuoSNJfkUudm/oM2z++INq5B6wadOgdX+r
XKrNgOv4+YTvObIx30pH6QdWdi5IabAOg7JXS96D4J6NrXbcy2bF73IkXM2Esqb4
Ia4WlSeDCMXgGXBCpZJPaJ3i9o1WDDnz66FHCkrZiHWYg+wf7Tbe45Ec4Q5zYOud
pV312rJ++wUkEO572PDq3h6hfLINrPcG+hMbjj7cpXfEU/NdkMqlDj2/HfCFQb5b
uL6erz9IIX9uyL2Wa2uQBHkKWQJbJMK0EVuqGQVUvg9Ps2qeddw1kILYk/dmIh0H
bopnS4uyVmJJ4Et+6otmDfc0opcZ4iVsXjrfpVcUrt7awdN3HEVOSIGwmNzl+xSS
zyCD/vVA0r+qRp7ZA4EyFRJ+9sTzlaQ/uhyA3h1lVdIJi+sfPMfLwTvuDtnbyCnG
4ee1i9FvUhjfZFdXJc0fiOxdw6BJ7pVf+F3iTHB0BTuFQAnqcGNKx6OCVgtK5p+8
l0T1Qvbqbpk1BZJ06vK8UR+20pfFSAeH5j0wrNkEsz47HFqodUQ3bevFtEZFu7qt
pOjgyDn2wzF3V4SO61aifKdyCEdAWEQ1a1bwhR2x9c/FsVts+VKnvoHO5NC31YeJ
X7hXgk9lr3AT5ztzQKT0PaIzkeF4cJd8L7HadOY9SUVPOCeYbqyu/0ipOT9Mjufa
iTvX+/GMqC0iozJBEg5ByhH2FrRZqi6qEY7tLyY0krYk+OVnGg3i2mIh0eRYEJVB
ceheV9NccaJwvw4htwDZEvqe8Q7WY9QINAoQ5ogE2O/q/fHeSpFSH+ConEKgQt0B
qSROdHbRkesOYkMmZXRlhsusTDlvK5LLIEfVJHFQMrp3Ti5a6NTe7FRDTmulcWCe
fuY+kaxXe6rexG3t707lUay175CfjliAPq5Uw5U7M1xmyUnaeImCCTaF7fmj8eTb
9X/zvfWZ5nNd5C2YV/hQgHBqFybSREydpsoKd+ghBUx/EAJ06EIsjcT5lRqalc6Q
//YQULx2Gl74HR0QTEd3HFyL1osDRz2eDjDoaZMcyYYo3RXj3SAfwh4Hu1quxlOy
zRMwqKgxidQkOEU6LnNjhqnfTWukdVmnDA3gtIDQ92d163DiVWOKAsrwVFPBMds1
lKNJr7K0ez+oT5a+c8lJrQ+OGvYRt6o44SrV2DnUAkJY6HKIWUmKGstVB8hmS3Vk
d4AhwF2O/wO9nHQZ43xUY1flX0mSyoTIslTtQOKdqIO9Zz6U0n445IboGtmAiyfF
TxUiPQxRwZNw1HGdiHh0mpbP9glGpTSkDcTIiXKrR8GzNpaHU1AWbyOj+bYiJNo9
lnCceZIpsSgPd74U/XtMUy0t9YYoDV3qULsRqokh4gJtdfA4QEAr+xeB/uc8bAYm
fKYEeri6wTSlhcePUt21EKpmkV8zAnThc7pbQBDV2t8Ap7VU4w3T73JgXRwKFW9U
SbXIhAKhh2BNBOBzBe1Nx5U8PIU6pSOcOmD0yowpBsSzvcqEzBBkcpeK0fUCVzoQ
vg0RQ6wRXjKSia2t2w5PGIEjq01SKUNFdD30zJDFN9Sr+CaXsdNZjERacxR2f8lc
VqjvKJA0KnqTIFPuqEIjow0DJH6N0qYPpRttjLD85208nYRjj3q89q9ktsjhw8CK
D+/OWqfInx0QhmC/YmAoM2JR99bG5FF+jnPFsEq7g8qBhexw8tQQM3ym/6zzXBQG
EH+IyX5otKNrUEJxjjFGyMJITtcEG+7YV0V6cokAd308+7zdw0Kf8p7Qo+o7C7aJ
J/3VNsqdm2gOLGxIz+YG07ORgryXCLQWbNAhN2AZRxiyueFM2i3JZ3k7lv31PBZD
7htvHFdZ6OpKo19mqcBHNUarwAnP94Lj1+bkwfAuPQwUQO7EoklG3yAAh5CZ0G+N
Kh91b3RNgSXq7SYZoyQDYsb9E2+dZbiG+Sjl1FGMK5FYtzrDPtVR37WF91kdEEr9
RLZvK87Dr4yAV0/DcwWLdWz6vy9RX1PRtuk0my/jrn5a+pCXTLBUM7vUP6zFwdZT
rGoQ7xvOAHeiMnHmN+2aCqQOJH49qnBKDtizcSO/VYaV1aSx+2oMvV6tVHyJcLUp
enFtavTY5pP5PB7/ZKD3SFRbW/IhTZCQih5/sl64Iq0ZkIVwrGC1T17KmMKED756
Ah4RXHAjmfhnkgecUQd5jfTVIkYcpm5QhuOFgf8NI30CRn/lHSQnjvwSC3miac2G
K3B+af2mKLH2YTMvksmNdqbUjgwStoi034fJwtF0d0UgVcuT05pFkP9u8CXMvE6A
KMlJEIlKUMD6UYWeO/3t8rUOn7EP+EkDnoJwJpIu1IGHh/dmd88RGHvC/FrhzJP7
KEZMSirMI1NClor9/fm6vMOGIN95Fx4SDvInvMaZO0GpBa6Wzh9PnaxQShBG2kam
tyRxYTKwbJDmT9gaOkxqAlQ9ChQY06ieDrKSr/5UEymkbhXdBpPKF+z3J9ITVXGP
aYSv1u5r+Svv/8ZTS8A4rhVedi3x60763QNOqfUUPMFERfKeUXZNyVkJunuWvdco
7yU5D64VNni/S2uZ5JiMksTGTj87xwnwZxKlQ+VnqhAbhDa2K1G04p2efNUyo7EW
lN6DlrHwqFLoGQr/pBh0FOASckf2NTIGonUR4NpYFkrlBsmySjdR2TVncYo4gpt0
IxNy0mJ+l1OELJlK8KH2jp2MvTAIHmhN05cXrxdGFvx45JvgTxZzrfKS/bLRhTGe
nHg3ffgM7KvtItQtSlVgGgAaUsfMETPSHXW6EQztN6WGyKXQYckGcpUidcwKOUQv
LBk0oYeNuvVmloutbHJE5JbsoINR5P4XgrYQazT5MRY6/TjbWEwtNV/ryXh1AGgg
Or29ZxzwAFQNdcKGib50TKcXMmYZpN7ar46jgYzXNlGSxWxbzh5HI5X0ue6+gin8
GUL11fqHjIas2kO7OEU+kev1MH8u68o6VKlDwd7jHSf4L0YSAfbbacgXPEEHKPvh
r+H2CCH6hS4iA6uRwrBk88ymhT7qG5lTvBw2i4iJpTBiY9NOYfGMGgha6PE+GAKE
jy1mGE5svUl0TOViY6Q2reVI3jzntkZpYUrKkd+4uPAu98TOj2LeQEMcEexUtk8J
pw13ZT8uZ87hKaS0+8aoVMaetPPP9mtiemKu0Uqr+BW8Z12oCgShVCoCoJ5gWTx7
QHAogeqF5Hiyg/SQ8yF2Jpm6T5V3q5hlQx6xapCy1UM3iOvDNByv8/jFKbOwQoSe
4rLGHZ2vAdGKjbQTdtypD/Oa7hy+y32PPrYStTxolVOgZnZH0BQKAsWPx3FZ1NWp
DvqnIJZaKquqTlaeddEniSFbDmk247YwOt5E+GhP45XiyYXWC9aHhlhcypyE9pE9
rBQhPHGD8tDPKgzRP83KvZLi0DQK6//wXnH692aGjHWl+8XdeO0BS2gwL39b9BS2
620dbdlHwVVffca3doTBCsnKoYmW5hPXrgQ9aFEJxvY6JcDwBxZbwIr2H6xuvZFk
ZQ6LC8Tp4HDXPpwO7PlU1y3qOm5/RwzGGlJhz+mtO3L5N8VyOrCfKlQQHo2kQfya
JPiQsBC5cqcqr5eZKorAkK8jnDbtjegSrphLPCGdXo406QO3J6Zcm9QfsEe5/BYz
WMOOTmZMYN5RX3b9DGiBeEd4GP2IRl4YwG+mRo9Q9fEUlX1hMVWGJSDE+96C5+SN
zYfaxtBfBC5+WqAjYAOdd3rcosTFeoqYX3tLbhzWHZBfJMkJwKwtjIsBDhji75JO
L9RyAIkF9Oa45RMB7iDyg82dfWoZWsn/Xd5qNFrb/wr+qmpsgWaDq1faqMtk79Rn
iWk0C7R9Gx2oKw3sz9RvpckydmrthnpiB05uB3Knn6q6EWWIy5S3woizWoE7wTR+
cr8UTj8pxxcVUn3Kr3SNpug2n53QciJgf/TTk5/iuILfxvBnAebr5ivoUsGuQkxE
dJJtPO4UyH1v6wa3IwalfgR1lOtSDgdYY+76Tc6XD1VfwinFkzzfmvK8pyPBE9Jj
8ckyogEZ2E0A25SUlskl/lgfMXOjZr1Mbrhgn7eL8IwFowJoxfv1IptXdY2sqdsC
Kh2fgoNtz8H6/Ii8GTwC/FrFQxt6/3AZ28c/hrAeQnN79b3DrWu/qP2tBa7nz6TG
USr9yuACIiG/Oz00hz19c9d3U5W1VnGcLgmbQdwQriLZO+plXNQ0UyFtrmGWuLiL
V78mgReXgJjx0BD+5hEvVOED0mKpX0EDAwc0u4emIi4O1uJt/l5GVfp0KHKnNd9y
QyhypCV6HKuu2ADgYVZCLhswpSXYaydnYvCZk/M8XVLTyQQZ0T4NB8xZTkMlMi6x
2g3NLVyjkxBUNUCCD3TYMafpSq+KMG7dQEeNHQv1sa3gZeqzYcsP/hdqup9G1KjV
psmZY6XMXq/mtI4DJk3+VEmxUNvDVvNWPFFb73AnagBrpgBUDg58AaKK9H1Lh6Hz
M75LSwGEh83GKNdkvFveoDm7IUiVMM+XtnZwX/fAiSfrSCJEurjoG9jC+CT95Qz5
n4vup99ZmbIAMMA/d1KOCq9VKnCiY5LWK3d2crnXzpUGBCEXS4MWAKCbHdUC0B+8
ZGuYYJIuK/xZx/aNoXZaugGOdKZiMB6dx6VXOtX1zPYJgxDQ5FUmSzYbqnj94eVA
Dvn2RiwGmHOvEeyhVhmfkpFFED79fI3ehWz0FBllEbNKZcN9pZGpFYTPxRUtvO89
82wAYv/lwploldak3JO/6nI9D1ArZC5aJtMTwI2estBzbdhlxsDMudj+v7rS9JwS
vde5+vj8K9SNemTdA8HtCTKiRxWeLBdyf/dS7z0YW7ZORx7ZhPlTRQ4phETPuWPO
tgDuLTRRM6SPdL6VCjkKNKAOZcHj5mx5np3Rp5pjBPWDRhW0SxOL+XzZQT5BpNRC
UYclHARSRCtAsU8DNwTPH2D9X0HM8wqFrpMdwszKaK+E6jFMZ+kJ85ySNHs2wpIl
wnoVq5pSwAQIxHcSwKk+AvmGiWS1l5nvLwIafHuH4BGXo6X50BzDiodY1m3zF9xR
YJLDnTFNURfvuYOvaBNFCrWj2YSU4uDKRhKCdCR0YnOH164LLlAyQ9LdRH2jS6Zj
WD0Xbj4fjyflaQhBfQJ1bYP+qG0lwSFk8toRemSr99l7wOZSqR7aoBcLxHBZnunB
7TEHr37JGthfg5krB6G+p1YDv/iebtXkHzqhDpwPqLO+3VsTd3rTAeCFEmjLZlAE
y05L9Ct7iGjTsrQRn4urQcf7p/KiYuZ+bgV8ZH52CMwC8+paJDCkmKVGsx1ivByK
che1CxjOwLo1NQysexXj4YolyHEPEAg42SOYKNv+e3QG8HcNivH+lsYoFqvoOte9
zR+OlthOrFc19JokoU2c1h6yIHz+4jWg3LHrjBADl5HP+F4EleQfMTnszy0pWl10
rrMDEknWHNRR+TXmhulDHIfuYiAPvY9pUWf1ZqB3Q/9EJRqK62bFNDmt5BMur/zu
QDq2xuq2ldpocECyRYySM9h9KW8vwaYTQFmHg3MLhKNH2eitQ5xr0Sntt05qtd3v
9owv5BJjSQaE7i8KCpS6gNvdQNIS71o2/GCiG5KOsD5hbzPMd6BwnS9gDZ2M0YjH
MleKKipN25i97X5vexHzHE7ubFGRZ/Q9sskT6Yfl5bAocP2rfRdE6ZfMHXlR1yCJ
3meIm8/c3NivTiZnTdjf3++0eSIWMzSpphH76bm7Gu8T19kCTRHq7Hs+y4gj3S2p
gJ+c8i7TpfvYLtMB51TEvMNT5HUAVkY2u8mUvm+JkitL+DqXXNOG7h1ePYK64hjb
Kdnaali4NlrnjnwdsrdJYa3Ch7MjsA8msFqSX9oJHO1G/rh3Z/+AUU29JlB8g1ow
fiLdIixlu8GICjhGwCpMiN5r0rCLidjuyKly5hwg86IW55ySTSSRU052qPZ69nnV
gxZl75nE9ENFJh+J28qDDCAGXjuUHkdqpQdgb5vHQH77C45/9w55n+iW6kA+FQJG
ZtkopA+KpjxXRHuD8AR548YYAWYwtAzzIKZxukNzpHegMhLTl1LTX0CcYdDJCF7H
S8WnODZBLUEvSw9Rt1sDueTtT4AYtX3E/E/qRmyZsWTnAvUNwAilB1754qnsXho0
juxKcJyimGTOd1aHOe0ATvMAopez7zDKXXWuDIjJJGKAs0H93qyImUrGZLjNDMCT
/L/CGINziDUYJ7Aeb0A2rURfJxU1swvugn8jlNxhoeukZC0b6DsCmAnUO4MhvepQ
mu4IlST/Ft8ABXm2svQb4umNArBrqAd4HPqeB/IhVViDgDHqJiR60bMQgLSLA/Jq
RAAgVRVRxflrQ/60Bj62pIThgajs99CwwNH+BeGd6F2J1TofIBjeXi/rz9HUGWsk
KajjXDql/XkCR1ThsjdHrtqaTJ73flkBdNh34wn5YbW84b2WjqUIbSo4UOlqblUB
bEzOWAkty23rLFBEQeFcNzbc+eVbYgP4BnMYJqTdI9dxka2duzmXQd2pBn8nQPOv
vc0xq3fvuRK1fTMnrnT55t/k6rwVrMk6lKYduDOqPdEWSIkGgp8mF9HsTcaTCQ75
QBVhDVT6hI53Nk0t4zY1FoiWbhxfsHP8Wn/IGMC6e1qwcsacqpUKHUKnFTrjfcsp
GCQOsr3zovj1+/7r/cqeq7WqEu5WyPIJ3zS0Xd9Qye9/wUcsRtZ8Bt/tBWYmngJh
hW2enf2XiTQO8lh1s2YzNv1IZyY4wvUsGEJC1Z6Qa/4GP+ik+/+4+DF+vQlTf+Ab
HP0/ZqQO1A+F5iftQ+V/kEjr0CO80OdcJTHr/xj6LoEatElaWqTVq4ocWmo+FPlk
46fm6smVGCYDKz8C19uPLiXUkgeb48WqKilKSjRpw0dFbai1pIVWbIy9F+0Bg9og
ks1f2oezs0IQtu8hYDQ+jl1rwLNrxwnWIYlA1ja+m/elkcwkGKdjj3Kb3hPV+REi
GdTWoBVOHujuVkEY8VVDZAl4fUQ9Kko/HwVdHFFH23e3/dvXHegnWl26XvmwZuev
2ZkxGaFvbyevU6UgMt3V9AySydMBXEXlol0AmoDmpBBuWdJI9MU/MMSKjPPEg8vw
Oj58LZo9CAFB34xdaxMYA0I8cFxl50ZxHhclv6QpKG4XY/lge50w5sAfught106J
cUqt0lUgam0P13oBICeupaYULxLic8FxPyIb8yQXsWBhjffwCYFXa26bJ9J8KfC/
BxBpAdCOnohXzxtiXGjGa233ST7NjGzkYgHsZmwAGdzbH7dppL81PgnMkoTvv9B1
3nWY3Wus3zMgJrA0yJR2EpYKPgcKRfti3yy3FtTXyEb2t3UJ1ABx1jWShY02GhK0
qYngtg3ap2Kb948n+vJdJJSbDxLYItgWJ2GQbNEn8ONg8/+YMen9U8csPYav6gcD
qXg9ks46c/VNmIPvzKc59Q4Vkv7RdHcbzK19/p8HWacXHuEnHt2J5fV8kerXgAq3
3JMVwpqYdChSx39TsZ+NuHCbiD/8T1aPuox8pifXqzu230az+eG9cfWbhvUL4uaT
KttG4UELDvuZj8qWQGO9y5C0taIogykhkYw/v8oPLAWenK207GpBv9Af+4rQhlOd
Qw3EN2d0zfSx0eoRthSul+Jh4fDJmWFIauRg/8Sys47MneEdPJ0IbiGFeDDc5VD5
kWmhvzVfyl9WRsU8mu63TacTxv7n0ky/k/njsnZ1YXj3YkU4uihGrH73UMgnSQwp
MEUtQYZcIaI60ZgfHt5jcktUxAoBBQIMf3gRF9cxci1pV6lI3P7OCyrdyB6uYb9b
L8Mnfw3U8ARHdTufAhvgxAkNw/eG14bKnhSY6YiC8vQb6u8yhnhQzsLSAnUd8uCA
Trg1QVckIbPc8lFH+umKxtx/tcxj7rLWsAaijyqk6BTlZboT01unzOqFUZwGcktM
dZcIDYloYu/gp3cYqnKyjs8auQck045sMfCP3kveAhOuF1/LrMlbz6C/m/9RWrQ6
2vNdmF7SFSns4Um2Q/kl0xmA79kD4EXsMoLYrdj5WLtrEjlMFO/nR66zNN77HW5V
ty19sNxhzLKCNm6utWYP/QWx2DWw2c6s5piiBpE8brHp+Ey0k5Y07re95t1mGs1Z
Wni4IombJfBUH5m30yvi5JDv201lgQrQSJxXa1ctzzOj8rDCryx6NN2fQQIypGo4
cv76nUbvcBHp4U5lXF/JsT507EWMVYJ2eNFhzeIxg6BPN5gVmLXzifk+A9YD5dr8
huTtbWSwT4hd2sfsdKl3YBpuidZWoGTiBBZoWG/1B9N8XWC8wM63E3zJhVR+gNue
cGLQYDcI7LPaZqGDhU5hdUgmtW2yY9wC+bOicR/QttQK+lOhuxA9+EWXl3PJa2Re
3B4LMjZ/UbAlDfCUlBclW3PrxaGXkrHrbbX8C60UO175zVhlgFg7Ecn6Og0iBDUu
y0d5Kz88muUWoV9fNPD7iLvpBprcl1TfDqoXED4277xeK9TCiz2fpNrWlR1+L1Jx
wGY77Ssj3ZRyYyZB6WLJUFnDI8KcoD4+LF8llb6eWyMecwVoGsgg574r7CEb3RtF
aDlSg+gVS9ohzP/5NJGpAsPA3qp94Wi7TzDhlXP+0JlCmPE7QdTsFdYQ9LacIxDm
HEvnQAZ/MQ7WkOMII0hL1t3xRq3hPBYFakTCvta067oYO5zYZcfHuwDUoSuabqZy
G2T7YxoIYh8ehUfrDVymnOiWyo1gwi2W72G2B+0IbPMwypk5we9Ivz40kk36YFWq
CrfFTP6IRx9nc6Rs7ldd8FCvHZ1ierQwWWMD3Z56i+2ignoQRUW9DOrJIPtdwzL7
zlZqDs+DzS2cM/3S2fZOJC3lHXL9GHcBb10oiaMyj8OGjtI/j/rDwl8nVLtlqiFC
Cc2jgg4MLJM2dGhzGIKHawvHQ7MVixAs0NiqhQJ7vDlgGqddXqVgsoqeChU/uR2r
37M2FzSdHa5vLUAxV1vbH4JUrh9/MfkQQEO8fBtt9iNF+Pi7H/1MBMvgFma7Om+s
n86VAXnYXkDcxBUIg+c6cvp/Lc993RRCoGX/rt2O/JAkDZvdUbJ1vTVCYHYMjTDI
kirSHp374mloKeKQWvA9y+8k4Z9Sp4kjLFIW59S0CaQXiMHEbOlhFktUPfSqpw6N
Jd7vRmIkGqe8QsFa+rme5GMB7MpuQkgkjxthjHvX5HM3cC4hwu5g/nhvGzZQNqK7
Q4p6cOqBTkl6tsRk2Bldl5TDsk/Jhyl66frO6uTGgubiw/5UdSnaPhfDuRaJ2JOS
kvuJNKHJHrNhSpgAB0oc9SMMgo/pRX1ocgpNiwf2gnRVdvr3+fddkKCo7fXwcdhl
NvRV0HA85n469zFlsToDZe/zRk0mWIy34ot8olHZKKyRIbRCkoN3416GRkc710z0
seJaolB1/mlxzel9f+TlvFX4MK7lZtAjvugYlYwgUHmhCx8ie5JoWwLHL4+RUz94
TR7sTpuM7Q2VE5JGoxD4np2Aiyo/2IrloA1NJoLTKydFc6qOtPTKWRXl33eHHe7x
hLzDwwtYP19wY7gq8VrPfEHWBLgSI/ZQAU+Ok2iQif0Si8fHIj5Yi9GimPKtwlje
C1oYRrs+8jHNIBbFZOukFiBY6pqI9ZWT44vPJad5QYNhF2gnjKmtBJDL6I/+2mKJ
TJOtqWu+M6peBzNFbPo94Ph1PrbfSFGBBDZI8EIY9xovZI6fC0ixIt4SKKONEYoZ
1/dYHVDVQtpWWYpU30fArM1pDV7D6ukLd/Kc3alcDKlTVXJBHtFaAUHB00vMJjZH
Ax3hiK6EkvYEmXuLpAySQw2iKyduCf0v2hx1yDN10x7F7MdP491YVTNzqM4M2oSK
XQyFkQHzR0jKEFT8ClDr4HtimQj5LryNLyohindaln8ET3eyveYYJLK7zEQBioTI
OTzRX3mya+yWuxE1SsuI+S709Xh8DDnyH70RHVYxDJ1wEdjMp6RSZXfW1nmNU0QN
Ginxu2trgi+HljC93NK6mEkLZDxOQcq1TfNASCp16nKTNo3kROQamY0CkjkM3wF4
NxsarpV47QSLuq2dB0D5Luah4uk7yKUxqY0tKNYgAA46mUqSFuf+/0ZVdDi4S/41
YcS1RWlOpTkatLKZ41B+4JvADwEvia+7gy7HSSCanZJvPiYuzQm5ZeZZhxkCVOYF
GNBEdGnKSsLmnh3iCxfaNgBNGl0/7ILRMd5jaxMBog3yuE7KkGFFuzJz2LVOTvkK
1C3Uw9+GAaJTduJsOtQKAjtVy4B50FT/Z5LCoRUu7jp0drP25WHFSFyb9JqQC20Z
kBuPfnQLhA8uU/Cu3H+sOOwgpsZa+sXdZKb7RAPXrAO4tKN8dUzk2apJjaNuq7yf
cRtpnaU4r0CAG7Hni/cTz/ONSrtzaPWyi6H2bhfKpwI+FgrzibiwVE9phu2ofufa
YqXGysudtECaHbfcFF5nYTFlHqBsJ+Z1vVELukvw7OaOJaepW+RnXbIQL/4ro1u4
P89OJh8ZDod6vKzk9sKo30LWJwwiqKwq4iI6bfSfyX7q/RX5nMi+roigoDnFdNYw
C97JEeEc/dYqjVF+//nAQK/3TvoPY34hb1QEAl9n24M6Vv3QQzatfW5TDzASin/N
LxNPaqoWT6ed/eCATPdE0wBSXTHO9/+VH+5qh6lJAENWkFN82SJ6xWFSlNLGGLLd
n/hwVAW+sLJ/leeouyGdcW8fRSBuiAjCBR6xJR9ZK3qWpXw3+me8tIa7s+JXtkHP
tDc0icTpz1WGmrr4s1H8Wvdet2/Lk+ZBSv12zwyn6hihD/+zr/lizQIGSFIfKiOd
kURaULDm8I10jR4mhqRduguLp1X0ibA/I9Jt7Sb1r1zAzNAK7+i6ge5urJeJexyu
ZebGhqXcPktr4J4xtMw29sM6LjG1hQB1BqdaFMNuTzXAuTvGT1JmNcxs30D1tjXe
RzNx/Wo2ZrT5lWmoYKHjV08ApoHYakY1bRCXH6LikFtM6eYxgVCcORZuP7OlahZw
G9ABLprTdFw/gnG1YeWFf4M9VPaETwoVvXrpu2Cn9HLl0KDX1BWVhyl1WNfqrWt3
Td/M0s1aieZuG/3tDrWP1pwpzDhN2KX31KSG7v3jtp8Dimokwn8OelLmBfJC1vcH
UoNuIXtxfPjKRZX0KvwV8zrHKBJCeTkjZODfAJgftYhILXZhaGoJusxvrToCM68j
SGXzskpiFB0KRd4DHzLpRsGUDGZpY6WWQMiv1G2cR3FnhhQd0rPmqz8inNBproV4
e2jHqN8nN5/PSg3Zpe7iY8vZyPUFjB3Gh/3siWFUj0HzmNTDGcbL3oYD8jMYvW36
0vl/bWlFnqQyUmQPaBX3iGkmiBt4pSgeywRczXAvh9UNC1Rab+IQreBhvC8l/Cfu
/RzlBwVjeOuzcLttEGs1YeB+1BFaPPRlriBRTv84QTSGB9fuucm6jjs9bSdOoKKG
WJf0sT0RqFAhittQDJwJAMmfUXsk132irU7K63S8tNL+o+6xkrmeW50TwJNsAHNk
jCqASAu8cMz3C1zbJCmYqup8CTIRSAjIlhqxhG8ugDmi7kBL+fdMc9WmEEDE4vly
onKTNg3uy3pMCS/xblM2/PdprdKHHaxTvkEx/cIgdNixOQuiWM6imBV4XJYXVoSL
73B9RaZrx+iY6NcPqnZ+e19HC+60LhP2D5JP2N8F/s3zRmq667YAXnGusAPJePhN
t9N+9iXEXsLW2HQkG/K+Q2UDFMDOVy56qAC3PpPoRxi9BJLdRx7vFmZ3WA2jEagz
7ZmEKQWVRoy9lM0UBYMf5W8t7iKi9SWp4bqlM8WMleoLVgT4HVWryzAFFG1H5eqj
4PqOifgWQLHVYbE3Zn6T8OhWPtT5v5+G5Vo96NCgMBMPi1ixzlgL6EMO+oS8wUhp
oKrXDzauzp2ZcIQCCeJtaXh2v6a6BsMJNsdlaUpwmigdz9cIbXorFOez3dKHNUm4
/H7as/xcFHOeSO+aFydOGWqhYsKQmAUa0uAZ39a0a6V5SXv8xnEpKYcFpErqK3rl
M6g0NicGKVHH4SOAJ/MH/3UIG+NJ4kmWWD/+qiSmkGFVmgl1FdEDL9rCdEyBQVuv
HM58yKUe6L74jHrFPsMgDdRsEA87SAOR38glArOlelnYU94iAjATh8vBaUgfjVtQ
On3NRlhSrD3XUl5krVhoPIoJ5qsNlCK3aqni41YlKf9EjxXp4RvL63kCMjshEkdg
lQ31n2rj7uBBGW13+SFVEm5Q6Bf6CHFQAR8rRtVILkePfLaeEdfSz0CdFCvo15B6
NB2VvWhFeaTprvh7+peVGHJNgmnS4JITP4YL98m3rNZGpNOqBS4DnOWcCzJZlhIV
1At+gGE+DNvxqCb22loaMnr0oi0IfHkY2q4PDp5sHeYGEmn7/iFbPZhcGocnyU71
yNukIXdXprpdg/jR1AN6VSknI9lNY2liFywOYCXmZMbMg+pLuNuoMYwwPdrp51Hf
D/VTKKtpBAxzGPuHqDoRpOzZNha8O7tFhETSLacy7nM8IXmj0qHwKkHW+pWnSmD9
lkt6wfTWBEDYMsX1AHPlok3IMr4Cyz8tiw+qj1h7h1nMWUFfPEAOMsLCqRvU8VoS
XZDJd/1cCgyScYbx8cMWVtz46ld1Grnwr+vRPjHOONpPzMrS0AquvqZ+9TXCAXPl
GOYXYxhMWDniLxdnZBfFWKt/oE14+V3swaQT7aYhDVN9Ywhtv94JA2MbK3rViyi/
8TyxhhulqrFf2iHmatiDO5eO3SFtiElwrQTfzis6WJf8zRu5KaVMLyZAec9hEI3G
w6QWvFgZZJ6uRwoFhYVg3SBOB0FVRks1LXKra1pFfvqC1wnrANILNiNdUtaIzmGe
CdN+UpzFOY0I6n0yPUy8KE0fHKYnp2FZ0ONUdjPwbh3N1Mdp0tzWhDVUwj3jjyHN
GXwo3WFfeK5PW94GqkfaKtuPY/xFzRh+j6qMTWe1PSRAKGGTB1RnodjYEj6F9uSB
9V75vn9cZRwJyBZz/0RJyRNWM9LHntjIXrDsOb/Pbd0vmWAFeSxYf6GG2pWlLb1x
E3ixhbbfZ0CmbDpD55YJb9lQ3k1JiCHe8bKZu8xvT9FxyNMnsZOmdOCvEghVsc4/
gJtaHKaMrunGt5sZTjb2pCEq7DyfOi/2023n4WSHl1Kl1WSKfvvwnO7FrIjwd5Pm
O91txwuA/B5qDSDprVPDO/Na8ppLRYARfLIvJLoL8AdGOYcuMqmJcBTIyfcEtdsQ
shZ+vOMpXTUDMT3K4H9G803YOKnZRWh0AQeZZ6JRYxalv8zRIKG4AG5Fg09D3SO8
hmdHG6pdLhcclJHO253KFTx/86aeZBfXpuIeOileZ32d7H0nr6sJZeBNXw0jFjo8
dW1L8GoccSoW51QfTk8W9MIWkqfMq6lue7m/3xik3wkjtuJvZ5Bw7L5oyyLvzh0o
S98RiqNSc2jOHJlxw8QcuytxwL+QCmFsCaCsMQuUqkhv1tEYa90artJSLbIx/P7k
DZIYvM8tdeXo1lk/D+j29OXotTNsBD6vNgShAJ4rUn6U8hgkCLyf8Ic/6lx3RqwW
8BdM081XwJnv9a3DHrO9cUZ03YfwK6yltGHsbsi27Dni1Xq8jZPsqql3c/ezS8Mc
WCDeUKlU6LdcB6f3dWg83Eh46Zf9ERpCyb6pCGyfkJMdlO9+r0U3V3LSthXY6VS/
jFZFdBv0dTaQwj3/ljz45ANE/ZH8AVj0sOYo3yZ5/7fjvXRcCJyrkDDwbPz1/5Zn
oXNCJLVHFX4JCXa4zGAyB+FVEt6wT/EP0ZpFg98r3dldOYzSMSYAHhOrsS4wyz4W
NNZ5a/lRpAsVkqFnO7qYfyP/YvZr5yCGpij0+gG0tqBV/vyxH4sDO+4P6BfnuYg8
fYHufit2qbR4CO6Ph6KOCBTUspaS8djGjPU5dS9/wNdjU84m89lpf29Q7itUevFP
EL4IB3ro34lV2vXh9eB1Bd1Gtsg6sL6VN06BGBAk1WXtCo5UyU3GSzatITeaSMrD
uWp6JKmARxt4cOBd6JNmDd5fUlcs3J2U8sgN++Iitf2X8/7hhdie8SdQgY2HNiTa
8bgPqffl81+vwuRcXs5O2ylfh3zj1QiVMZCvXmBKnJUFzsZ0VtpF55dCPi+wmLhP
zxkle4FHiqdEHGWfPjrotP2cBMsEvJ21jiFWyw4mwK8cQg8k66rUPJKyvJMFHOcD
fq4LRaUyVo8DyncCGnW7VrRBXDKNCgOBjNxcHzwYAXQ/wzcQPameEbkT6rBAs/pb
3RLBXkWb+9tpukuqClNFgwxwWCZQbzNBoFzTOzmf051eTgvsPPAJn0sEd2oeOBJH
UeeT+hWDAYE2C3Xq2nu9NFeAaukUXM6HPe8AHtEgLEkvgOp2uah8nIm9VXYfVcSj
ynCAqInuxUk18b8xVqxrq0WmQOOiT7WeBkFklLIJc6cwj42e0WbzjuI8YhwcpdR9
Y5286E5lbFNbT93Kx/T0jQpIP5Q+xHAvLFSYIb84A0VKP1Ef77vmm/YUubWVs8e+
/1oA96sbM3Z2mZktu3ASC5jFvOSlLMSNTyTVQvoM9azvN+q55zhXtBXESf+DY2Lx
Y/ekeLjdO1HjDuVEFwfv63ilWzSHmLsj74yWC1hjBHqTX1SyNpoq5lKxMWHW/H9T
cGiqilMtO2TKzy9ROhc601nLBXnwdPOinA2OPdmyHjKDFBDThrDLbImfYafrXlq/
+Wa+pnSKn+FAoV5GdFpQWryv6zt5SWWQ7YvXWYu9unGHFwkOfiM/BL+4u0NVR0h9
4JNN2EE8AfmXkHjig+h6OmzUvG2Yl7VcnU4vbqPJCYZL8pl2nVDQ385fg2TL104v
RDdWVXpNo9thX6q1dKq0VVMl+Miosi9nMdzIMRl4/9KxCUl538o4xcg3LTtaWDYP
ACfMft+b4NQqndMdSnB21CuwpYkaA8Cbvxa4eN+s47nnZkC21CskBvHYYQVwEcd8
VAFE1YuP9xEnK1KLQW97mSi5rSUoaNJGOqIa02PAZde+nFx/awOxzvm7NatmRhup
5m4JOd7eo0YdiU+mJvD2sVV/GxgKLEHUoQC7Hu8ByVoLmPSApBr8WwZ7Ggg6Xocz
56cizz0cnNVACbWBTyDovzqWDThQceMImycj+bTJSwb0Q8LzORn5yOUKsOq+xqCV
Fn66LDih3IMlNpKFxc8xuSHYzje9wYwD2ykVLjlnqbfW5e+LZdyAr+2XbHsxIO6A
UaZEexV0pOe1BcdghZh0RYz+BJfT9Zio30hTA/fPgpcCS23i8VcVypP3NFro+2TH
lL0QmkxrJ0hAvxZ6OFoYoCYeK8Yf5GAnBydIEkZcF/b1hHqC1kz5Tfv1gIfI4Vp9
0KYan/HiDhsSd0yIcngrXdQQEvRi/dNqHhJZ5pyJihOxFAWyYKkLoIVLiLtLA1M9
D+qI4XjjezHf9L8SIxDnQpdIfaDuJ7h4mXHvpf8SB7iCi9NEtRKWmWX83GqJS3Xh
aUXvfwoUlDeYY/qJYv3+O2t+WwHCb+XGISf5kAFIBMfhJxUIF18Vup/cojJ2jiVn
jUQpANCanjX4hGkXx++jhMNuVcboWlllJudr7vZgncVgPKHSMxk/GOLqebCAdsAj
x51Zz77dmNtDCLuGvdmrnd/nt5vCOdlhGkPrwmYkrC0VN9tRWSefV1YYbbipFrYD
Z7hv3E09uRWcDtTZlJ7pBPr9ndlCzhwHwk7OrHorWjVc35F6M3KXsEKYuNi7m21l
XINv8pIcR25h64ocG2Krvv8qZx1ntcIAYodLtdfrbhdCYMKsj7YUC0Eop5DfRiYT
CdfQ+94y5TyXCeYe3B3WpTKfZi3+X8Ov9N5RH66tGpW7hFurdOjM/sjNVtuyjJ5y
MVxLwPJt//elO8JkVlkedacTDqjMB5Rm/WtQMbelTh5pV9OW/tg409D6InzlD098
JLi0Oj0CHBdb8VcTShSHl6Upx3ayEsoFLkydtNxoVDhxBba3aEZw5Kvc3MrzQjOF
rDUDDeQzW0fqvUHOG6iZ6YqY6SXxTRjqs7jB+9UvEJp+LJw7eeL37F2VZ7/AOVjX
56Omcl0VlZ8r93NszP3tMqcXcmeyV7WyED8xYC84M9+50KTztqdRhiKyURl1rSHQ
pqdV0p5HIOfKXhdVazq2ZLsm+LvKacDPZaP4qhsIcLeY7xZP3P++2Ff4Wxaz7U59
GmyLKr7NG97DN/LVs98QkRd4HxZi2xIlxrb0SyB9Bj2uzd/lNiepeAN8k4eHlB5k
v4PqzIyemicZvnF+IdTHtyBBW+NYduCCrASsWi1Abl/IklvyqE7jDgk6FXYC6ahO
MIrZZg+rEk79RtdDCGzzpOibyL9j/ml4xzMy3yUZEG96TC9Dhzz11E89T4L0E4WZ
+3r8MYhwAAlKYJn7fx5UO9AUtyDAgeDiMvc6T+ch6u3Se9CKJLGAPOIVdfNIeN2k
0QUICkhMY+zXJlvItJF4Wrp48A/UFNk45E+DMNFKwukwdaFE79dsaoNDkuHLIwt7
eRZYeDoWiBM4ea3uOoI/xyMND1zDWooZCgbquXrm2ArNAdqcrQlmSK9RarrvMMBY
dl0qgRgd9XHiaF2JK0u3JN7JIUXbOliILK6Gz3CygloXkqxdUQJBR7qe5ildgqm4
n50Hw4fVqIR5z1CkExIH6dFU7Ki90dWfR7rz5cwatOA3KQ3MW/YZLWLW96HiOU08
/iV1b/hTll8rxwMUZbsxpm/Z5cG+GBQDOzJrbHgQLVHnMj/RXet8Kl1lcYPZl4Zr
3IxnuPHhjgmlvxenm52RLz851GKHwECdDgg6oXIhFNOuCVeHPhnienM+/lrhmg+r
RG8DLWMq1yqyzEJZO4Hkbj/ip+Yk8T2UbJIPB3TPwJLDzrxDPWgso+BncokPpUuo
nWMWdg2QyiBLqWSfUph8z9+WeIiVwaNkiNqmcQuu/ZAHRfO9X1LYyP63O/bP5NXZ
XaNKjJq0ed1jaabfY1yqErey3UbYdh4xQpLDGsMqD4FnGhNm4t5jyvqpAVAfXSqs
b1Y09Z5z/kMVWgIUoTRlYHN6YlUmA9tSo3ewLckXoD8uI141f+0HOL+QogTR6Y9J
5ZqUfAXwrdBmMUT6BI7bv0JT9C8KN9MrkvEgbNRwg1c5oOJ97mmB3YklQSoeIwII
RtG9OKGM51urpfNpEnQ746E4eWVGXneiuRacEg5JdL1sR2Y4zsiUo7/cHKD5yeMO
G617LO2PUp9V7tcEsyMbCDnZo8vw6z7kdyyw1bFK2+ipP/05bwUnj4NBeZzKASWc
fGHO00phoyVSfdV8+7PAIYFi+kiJANRjKGC6Po/Axty+f1uM/eh3isRvWo1a1zZ5
9JXk3k+0bfuYxQ30CHYjDlA5cys6nb7S4c1aGkBxWNA2sBjTWt2qaF+W+EDdO2D6
0RWBkOFXupySkfcJM3H5OaWc4jwRRXZ9LdJ4RdgHx1IA9hbdrSfukgdNaFGYy76d
wvdOiABQ3o6JYPj9uD6jsMvIzKKrTMUgRGMeoViQ8JNwL/jwgVJio99u2yxMP1Ob
XD1lkTzgi6qtQhOw2+8i7DBJhRw2JJGMalXCovLnP2ae+SOdOY/kjCkA/INSFSdz
o3wqupLUWYzfKV6l00hWwJfeeGleswZACM4HL6VkUwrYxzN6z7GULu0rJwFQtwcm
hbmzdtA1ndkiMR12EAh95N0z1VBj1Y34+93er7bykv1eqtbhg3JSDCpn5APC4McF
/TkEjiTTR9+A/Yvb3uM0oKvQzdu4x8A73bfY+nGMqtfOJgU12typaQiFaeJ9JDHr
gVDpA6VimXVYjTsXwvkRwM8Pdr79jM143k9EZDpqyawhwAyGeWE+hK92KTceo161
Q0ZCaonyn3L8C07sJYmff5mrXiL3L7RePMT1vlLFdAV71lBMhVr33hanlOjvQH5B
bRnIawoLJVD43R7nE7o1auVA+q5FRzHX+ZCMutOilxdERG/p2fLSc6yINB5YDpWq
95GA2suYKAneFQhTIouh/u5WfrTJOyAkb35W2ssd7u11Pl06h8GsICciQaaZBuYp
uCbcRm8yj81ADLfFDgSvpRw3om37CPINIk4xWQP7OwHoXMd3yr4EaktSuxGvLrPS
FDEWudwG9FQTLIBM5aRPDwT2t0C1tb4sIn+rID5HuYliY+PFQ87xTXRJt7jplRUT
xZ42J9jSKr5mKhZpmvybt5YxR+z2xltvlOp7tGz0t0Kw4RMGcL5jC5oKVxo7q+Vv
oihngCuFnd/FqkobMozq9A81cGSEeHuDoOWvY8wo1umPl8COISUsA0cpQcAo6/wn
42bQf8s6qugTvGSJMPdm8L8pAf3RlQpJ5KfVvxM7n92W/kuxP1OOAl1ZdbvOsA6a
G2LjjF3JZgIdqTGFWW1P32OCrmQ9bojelCdq7+jkxvLD+Fcfco0gINXiCY8VUtXK
3buSt7EX54GeuGAx+iBPdUbJ6sRMGY7OL8qaSKEMHS04vT4tmmsMRXG6QbagjsXr
stRi+0m/Ab02r/IlpJpcI3+aTTOQtib5feEYxCEqwjwGyCB71H7Xa8eerhV7Aeki
4PWUy6BIxTEO7wt0mhtNEcLPxV6wrtCmaz5rkJWcZNQHbT+4+wHRc5gmUK/jZjmI
2j7Szs6TGq9frGxYFHYolxA/st4q01ixCyBBsiVzW0luQx9o5Sm3uRZ6QiQisLbx
Y3AiQQKOg+G2/nPxh1pfmlso15UiZIlbL/gcZnJD/JgaNEMRP8uSVyPpnM9h0BpY
x0sNO2HJOQTw3JuUZz5NA79ky0v7kja7PSEXHGR1bD18+HOIRoyGA0/KHlRbYwKe
7LI6To8CZIl7c5+9PIFqc4DyVkJf+PP+7Mn3/Fx5d3F5kdQT+EgDB38QZl5dBzSW
DTCIexqd480e94hXgkw1wkXYCUbs4AGHfJEeW57Ppvwm0YZKaVrAnl9uVoz2RBbS
fSZkF0C5cX10Yu0mgFrhLlljOYZkWB/8hBPIqcJxthT5VZuHUw/4S6kA1rmWi5xU
bio8uYTSXYfRxx+nIc3RgWT/zcfcfa/NcPct8KZEURwvPiGRQSultMWNXBCsXl7e
jrr8jP5Z2+xWb9+nsFLzmstH9YAe24/GM4cSsH5jrK/GJpBVftRlbaEDJdmx1gzw
cbd+bXp23WiAH7DUw0gvUlsjRFVnXqOJFS7pWBG4A8gl++NPgqS6wHLS2Z6fPxiu
K7HkBxlHGe+IN48tE1Efl3eGtE4gf7eER4l2MU35wEkh18zK603eaJ/SBR3klScp
JwvtDQWnsbNrwZpBkKyAdTgkeDL5fbYb8RwSARfdxTVJoq4uT0duRf9whZ/3KZYc
RMlpOf8OgpAJEjLBziJIQmROKsSycqG69PQIzwEPquY2cQ44Tp+IpBL+4GzwRX8K
qs42PfZexYSuTNcWnoO8eeIFDbovqPL0pK0leHXeQujfrfRs7pDrEpMXvlhJAKNq
Gabc19MB13OBcxmxIl7vfJNgKK7LRtywvV3aI6ZljT8F4/dbzO0VQpFIDyItC0LU
CErx5YAQVm+Y4k4p7NnDBxAK5M5Yuzr8spDF7kVFYTjjsPbN0LYrMUUMSGHOLGm8
oRwFpuyFLG79IBj5X9g6mddXljpXiQQGBRGn3ReXjYcv1/OvQU/ogqPaVXtILzmZ
Cq6h7LhtqyyrpVuvNdrS6tfJDaBjzssm+O1oCQMRF8lPYM0KZSasNGnFbf1/G8iI
zkQbJBQcm6aJFip4SqcMsxL67AcNkCicz/rEmwo1MnO0RFdwu+4Ic0PaGK+8yEop
jMRPC3OC1Vft4cK+gqHf8t2hr/HO3I2KNvjAZYwoAxLxf8Pevcxr3MwV8TJUf3GI
nzpy7OqxA5K7bmAXWlh47suwzsdTl16cqQDgF3n2NMwVqyJDQaW529X0o11fY0oE
SOpYfx6UddC8YHeimnx82i20KfiqoYu/dEyL0i3Wxjsyz4FLbAx1J7gL7N1SHB1d
kLanS9HxyOZTUNH8O11Vt0DmK9Vx9vW4sflXeg8OwCH4BZLksUjqWn/VTZcnxNPM
nJUOWUk373dNNiK17GK/kUnS/SWLx/TCRUyoOIbtbF5Pg9AdvifMTVktEdDDSK+f
VVtmcGjXcudXbVTIfPm0KjLIWBRntRgmz/l7ZZ3HVf3MjbIQchv3+MfoqYjY/Pua
DyaAeI8ti8ICSKRwZqRduO/zJCxOSqOoqe0F+CEm2RewwyuDV3HQzJm1QiarPa4E
EbshzmgS1IUCVhGm/jPkeIlBiJAX38UeuqjV/4nnLcRL4/ce/9ytCML1oUF8dN+l
3e1SEd74XtgbhKiL4oPfdjfZZHwI44OA3grLqtNGDt1AuvntlqNnMATxGARdgY2R
Q6zauAkGJrUsmekTz9QIw/EUiwuCBsG8uayg5rHey72kv5yNESBcP8Ib7UkZQFT3
dewNQC5+TPkGUYtcZ2FO7WM9j1+YSTzihGKKuJl2CLFDKhPEagACE29+R70h0sre
pLzGFx32uzysd+9q3/7W794wWnpXO/5Aqkr8IXrNNygL3nRHc5I1QTYWGETV3knm
fjfiP6PwtJ1+Yz2/ZKbpwSEEuZtUd1/mDGuV2l3dKljmwq3y3/P08ZZ2QpugfT2r
0lwWs+IaeS42QObJ/v4fWRQcBo5hYj+P7jsUPSzlMN+ijlrdkk61I/dXwohgoXaq
/hEAg+gGSL8PWxTrbQfyiRe8cRhHOw8yb8ZB4FVX1e2LuYDX00uiuRrGRkegXNzI
vigtsdJ4VdJD80qV4ONtrJeHM6dFbqc6NdCJJLFNv1Fc+JCx7jv9ZlDMvIUire5I
cZzOzwb6Uv903v2soQZh8ydtqihwrZGhEMvNBqjRZLM11b+XbADppHaqw58F7yp+
M5/iihZUtv8RiHqetQFx509/hDZ1r2DB2ZnezahpR+i5V6wLVKKaEwFO24eKS5SY
eBiDr2hVbnREAFdPLQguHzftj4t2l6KQmirdiEzYgBkJ+u7/d6304SGCUg64XeLU
4PyihzAAe2BL4LEuUnBBqRCywZiTaTBVZnB7X9js6T9jaTzZMTY+XRa2fPjRjI2j
79nvjvS+rsRrc/Du7fblu0LRXWmDLjW+DxCVhRAdBsqSrMFrElkcXUa2UFfcFCIx
GiBRONcbhuFd8niByqfON922YIvWtdGKImL3WQfHWi48jx21F1NAWzQEoLHCrfGH
gScL0+wyGi8B+p0PeFKwKDCuSsT7kePR44BQfhRXtUy+He5aImNI+dsNWaupBoQ1
FSyPQ1/+T3WQugdy87o8nVVTrzjdpZo7lJ2DKr30d6UFPK+DUGb+NGXaE6XlWGDT
B8RfCa9Y0aR7SwlkTNn+6iD2DqLx57KKc7JgNJBMeyQKPFCwZ4s7NcfGB2ATr7No
SKZ72QmPM2+HMj887WxvOhy82EiQ/Dog6x1/Ai0JpLEZM5UQu0dJElhjb1/9psAS
ZNoUHXWH4PVD6VA692J+LgtuIhF6wJNFV0xpN+DfZ9i31G2yvpG2vrvj0tNE8qc+
NBjgwKZtvB7E6QsUFcAW1BgSZ5if/HNGLaaDeM73Tjd4o++aLbTXywwOaJISyhym
aUQ5Hgd1Z8uydJYaVTKIpvLd9/ud30vaLhPOnXh9CcwvNu1bYR3sbA2Ws7ZA39Yz
ROlhCXcatHeI77bCpedu4j25NJIJzh9AdtgXAfZaQJurlBA3exfDjXklRuVptk8t
DNc0QJkf/QHe7xwmVHwsiKEd8SUYwF91D9uOtPfX3TpnsUayIBRP8skeKrSDQnhk
eZE5xMsQJmrrzw2hfE/AbiAzmPRDl+c6kKfCoZY3Nt94mDeQPa0GKeiQmlzPXXD2
qXTULmGdHt2Kt4oFyosE/tJ9s1MCNg6InD0EK1e9uU0g4EWmy8MJHRQz1JF0daiw
OaN/qeSFKSq2vDzCxZ7eUfz5UJl8f98M/ZZ1gudFvlWi1QEPPN0GxXOL4n70+7Zf
abrR/ukk0JL1FgCGa2tnA7crUmYLkv7t6HEgjCBN4qBqC7+ryGHT63R/58MANOwe
iubDqZ33H05hDrk/X0WE7FKHkTEZiRMXpogqovldbI9X1rldhTeF0ciItr6OpJcO
D09iARbnfBxjAE7NTTy/TuN/n7um4uBwrwPASFiUR92zUDMPYRdOCxk6lEhkZ9k2
ePAL0WzuwuHjqWCJyKVx8iPJGqNgsGQGsUJbEa+QaGtxFqWOuMmWMdmuGeDJ4RWB
TMLFFmI1iplezBUuhuDxVPz1de34spxBf3BjGBWfUD3+v32UE8fOnQbkfSXmWQm5
0M4hsI7fc4YXJWQd5U4SrWxKFxBdNNKooWzLkvH0BfzCYnuMMFAg8V3dXcP981Fx
m0QC8Dq1tkZs+NrSzBRLanDLqxQrPaDPWz1UmlnrnKuQyspmZE/KLggoNc7fMKwM
bMpAjHG9QT0dqhmsQn/Nbxw/47AFyxmyOhYxPqJawNE/JbeRpSbtnRP+81+gGDkk
Lyu7zE3X/uEa41Rpfr3jhJSsRHhaVDgQ1Dfu5GsIyxF5t3yD1gZAAvu/hkj+AGFV
z8JXcsq9dBzPengFR/4vipYOCqsWQaT2jBlldrmzVZPBC+yDDZpY+8GHLU09oB0U
hNWpOuCLBumzQ1kLzPzCBCS13sQiEykWO80nJhIEYiBuGir0h959IhJsJyPHS/aj
jV2wHQO3jBfharli8MOJ11Hl03GCXIpNYIJs0Gdw6mA+BPzYmn117WNwd4nLCG0C
AzMpjsyZ5WeqNH9w4pplyGk7I18DWvbra3f61o3LG76nlrJQqAtyCA8UfmSic/yc
0N5zb3Axka/RJpYtzL1Yffdv6Kvd6UEj9ZcJ/kdBa1lL3NJDOxevG2vfzGhEK/Q7
zOLrNNFclEVqHrUyAa9tomQR2VDvsXBbEEDo63wYuSO8GkmIIIy1OxHQPI5g2m/p
DaQbA64b2xDBaXx35ajm348D2pyyQy1G/ly3dPl2+V0pky238Z5AddmReekEfOJ1
G15411T+bs0yeaxWiBIL/OWYqtafnZhEQxXAftsTmZNtSCUumygxehLvvHu1BT/k
i8BOm/BRA2U3eVAN8PtSOUofgB1muSOQ4PWyE8X6aKIvX2tWUcGPQhkIzi36wJsN
9Eb6tp1pD+GbutSHcOgkjRCziXWX37mmp48ny3zTKBFA0Rq/d7HRGbJBKyu/HzuM
oDu68IuHU2dBsRn+Qpvp3ZzywLnyiikfuoUHZi+Hrc1KsyFSXgtHsBz8EzpJEpN5
G7l65vpepbccueD2jWMexd500IoU7asP0pFJmyo+OKYkNTT3iMEyXxMDccw2pWD0
4CePcgxGnxjoWoLBGGgjlF+q2A22u8bxlRTfH63aWIQK/NvqqKRbdpPBW1oWOyGX
nOxCE8mnf0KAdN2ohJQLOIt2RAAIa9lyatv+4hKGU7KML6ixepvzlG5S4h4nE7vF
ITp5gQUrqsqaLYE4Y6odRb+L5A1hyn++FzVs8EZuiXJb8jZqz/UhOYcw8gFtqZJc
EfU7Z3YvOvxTqbrwWRoYDH2Z2nsu/LjrYkHytA2/LVxZsIwMVqpdwqY95fdxxaVe
XqTIee9tPcchrON+6hQtwDNhkugC2MSasKuA2SOqo7I5ugJBxcwIZ84gVtDf+rEI
bP/5jnGuPoUbvSDNx84DBR3mDwIiU3C5MXN4aYbGYJfIhVI9dNdXVE06dgkgLjRw
rAIuZug1QjiouPFEKJ1btoplMjZHVZ5t5ap4E7YH5v9JCqsaj71SuzMksbZ04pjG
EsYeeV4Yq22EpN711uZtd+GpQSG+FVSE96CDk3rykhniXDhnRRHClaW0jD6gxBUu
VRqeSYIsW9xMoE5S/wCfY+v3jeVq+kMY4ajm60nquqJqR2YAphdTmmstdlt3zVxW
uxD+Z/aBsjNYLVUQzMFuOKLuVtVkySZdLJKA+Izh9G5ZgNX50+2vKL4/Dppxhdsu
wzDWMZtOJ2czzm5KsXKZdKEsomxxOccFpaStd2g36gXXUa1HZoXnbguwgTI1AhSQ
yFULbqlxw9kXsiC8BH2ACVuKvdGx6Xsiugz7ZaaLqNj1aNta/TBUf9fRBEFE2qiZ
WLqO1RQWpI28jUKPqsXOFjyNkBL7Nu2ApC+CCg0X3vb3wDsXCgUn32B5gJkqZlNP
kt0Ssq+b4QQM0l6vpakVOEuI5Pnp0WoJu04sZEkEYYaaDNycYocH+0GtpJzFcz8e
mHItbGpGJ/v2VymNR74cjC3AmpuUBN4504POL1U5c8qRHpC/h0ePr2nAraKJkZ4p
WlUK0hUfxjCo7v8EOle+Y7zHpo+1FL0Dy/R5pV6ne5H3RTTfQ4q1FXHdV7XF85yS
BKfeqwCON96XV6h78vav3bdBHA5kW2Zdygusr8ZoFz2QjEVamNdLDSI2DfaTRZ4v
Ki+D2yjy29UZ5lyNHfdY+5XYh57Rjy2oGEZkfjCrYufjk+NMsLh40+pjkrkXam7T
686cHiYJ2V9SG57Gv/rh55Z2DFlgdZGep24K06Y4Bq2j+9QRDpDFicz5qT8AdqyT
T/jwt0hqsubiXblfCCNmzSsVaBH9SmgxTiFtVsy/PHydjqYMjVMrJcmnY8GeUe34
98hJJpUitPQku6KnEFYHNOLUEbzX2o1dSUUzFo8uMsiOL7xXMQFWBPjsKuK9aFkg
9XMrDbtvFfuu5oJIX9bZ95PsM8DRAnOlA7wjpiwMqe90iT5xOSEroIBg36mrebqG
0FEYbh7DU37yP+Nz0JeJu93DHHOaCzJzxLQ0Lo2PcK70ecng1KWj4SJQ90S1LVC7
nOEQhYj8O4Y6HSPe7QBU11PJ7LWxrUf2nvFoZGnmtH6v0vK7Dpb2Sqsu3YgDcga1
rABxDRmDk00MPRCBKDqjzFAmKZiWVOYkuIK/+LfBR/Orv/LWGrrtyV0L2R8hzwvH
aUfaKyN96eiK9X+FTJCa0p2gu17G+ABIY3Ao4WiBYGngHRZumqZY8avVW9x/YVCs
M7ZV5MCeLZiYtAdQRoMT6lqAxiES/WQNmszQ/tIk6vtk+0O3sq0YYKdY5wWDmJTO
8o83tT5YdbW+wVho5Hgh8MZIT4KPtz146wStRF4Ri5WnJrpm5Zj0XZeMLWnYG4NJ
Biu3CxjLhG1JN0oG+ktvUx23GulskQVnWopIlJWCaxNGoh02pIHi7Hjc84R2TBNR
Qwqkr+NS4ZscJNWoI5Pk1PfHNB2rExn8EuDh1oq/OLai6AQNkF5e+pIk1e/LPvlp
Qe0cNetLqbh1gBGvkuJc8gOK+CveNEk6m9yjIRiaCZ8lYa3orYlHQHXAkXcWGkSn
psVE5h+todehseaHByeGNev445m15jVD/4kxQNyH8JB0tExEbR3u550UXff6wSUY
PINGYBusbuyoEbg/XDjdfuQHabCXcmbQCF78SWbsza/RMrZh6dDBk1DZpYuaSEok
LZek5p1++Qusz0Q84cYNFUhIeNmqA19cbJfta1uJqyk9FrNxl/kiC6SKJsU0DmKP
x6NFaGS1gueudf2REJCwTzZ7/ZTWBh5knqKlpgS4ZOgKao3c7q5KRObWtQPgAWik
c2rTWuGb/MFaTgP5dKj6t3l3j5mW0AKke/gTvSXAFJ+uAoVlhO2uunc2E9eqZ9tB
nqrRBVTTMsrqxRY7IE8JKtubeYAV8OH8eX8rCf/i0gPrrhd58C2VYNgdhJWfmHAE
FTOQWybSGkRG6iZpJ6qoSS2QP1r40LyisPLWQQG9msB0/mTCgiMTlz7yRKBVTbAO
unmDm4+gDTg2zkpl+y8nYSGjSK30IfuIGMWErScaKds1jwKyfX3j69XQYxvffPW5
ZMCNlILaPz1qx3pVYu4PNNCrnZXv47zcrmaLOCx1H2QvbTXsp0eGKpW58Vxk/PjI
mhorIC/9EvjUBWIq0yPyyARCA6cS+ROoOmxUBZkvGlAVMjQQXOjJbaIZnOGVwkbu
e7U1j3gK2Alc8TZUg7/xtU1U8kmMCAnlsx5XxJhvQwFyGsFacVq8LnlI129yUz2v
TmH/9ljgIdJklvb7NpfAZnYAbUTmV+OgD4BldbQezW4xCS0Y0jl6GhwMjxxYv7Y7
ORCRDG6Bya5I6EfghM0DuAv1Db8j8jxaGhdWZt3OLBF4DNs3B4nmlLRp4GopV+Ff
n5RxfNiTg7QgmpFZuHo3xDk28yuY2BilH49o6drNNbXqnoWeiNgTXLTKrp7HUIyf
30JI6OOqrzT8W5tXCLM/4sIgSqxI3HnCIdLExsnsXcGuxXlV6SMZww5JOhqFaJ24
Jrify5RVHhs+nIMvT8POjUL8mvT7UKU3JyoDM7sRlezb4sr7t5DE6RB+gCc750i4
21RU8MhsjiZ1MZ66nw5VIniAv4Aug9851Tj8lEigjLNW2y/byd598GZsTadQX2D9
WPfvIW34YYk6AmBNIljsL1rnvS+wNeeLJcbMs+xqcN3kgCDH+Udb8g4/IsXgvHsD
ilZtA2xIB4Nd+nwhJyu+KlS7+0QCt3CciiyKLJ7T0H7HI2u8cek2kk7EiMrqQ47t
jexoUV2K7fCQOou4u1rDbBbn4+uVmTs4V4Jlreka/g7t/wIWm5yz6ZSmNs4o983g
0RAn51CAvSYiivOWrlU1puIM60WsEHzdPrmg5Ha9dglYSP73MvuEfkQX694YrjKp
93j1tKg5dUizrE3ofwMGDaA1OLorwA6nba+0eNRzQiaiE1KlqVQeGXrpsoa2uxjD
sTjeWyME/yg5HcQ88hL/9Z5jHQPDoBWWC8UhxqZd7vPn61nADxWCi3Bve2koeAIk
+ctmECBpbMyh5oHlZsVSuePoStqd3rv8orJwIXzwXcdVokBzXzzVua21w77jFMmO
poGjsrSqRofyEMtSEhNzwBq8XWRlEe9LXmOJPQKghJhu0H1x3DKjNkcPla7tbCHS
+8SX9zKHKbG/g9J0a+bhSTMr+LM8kUcxeY/W9msY7Px20ZxTeXJlPM7vQrrkjyUE
4mPr2OtcUBHNjp2SilP5vPCN/967NaSm8CTO39v+YhgGWJIPkINluPmnVwlMhGlu
RIGe3EBJwkGSA/lKyc6WQtrcATfZipX9NTNNAOW4WJIGH07e1z5O3lURBrbXqlAg
Mk06QqVVybi8+nO5oSo3LDx+R6JophNntxIFO6RQdXnQGb3O77yCa543msh0oApj
SBl/XkCW5uIjQXnAVJV5+CQg9VV3PxW65+4kq0IJ5q3jrWI0y96yxHBvhC/BbrAc
P6xv8qZn1Nkh6L8uIPSNxLYsoRs+v+udkM+uX/jMnxB+KTT2PK+YaFiQPEf/Ummf
h9xJolyTXK7WHxZKNQ4I92Uiobra1F+0MKXpFugkUxhfy639VE3UFf90jehZQGeu
iv1+ueyknN2gdd2oNh/UNzauY59kBHPmMvDzZVLl6zQz/W/KZU1Y+u/D7ynYgSoY
zWFRONkAx//f6Xa10lUXZ1qUqizshTQPz32S2Voz+6ZfRVj+BPc3afQxyk4b1pXu
X5BTzH07iSamiS+QdjQe9Dtgy5vCw5NwQ8dlxvNhhJBksKeE/ZKBkVTHPcMe7BD/
4Msv9ikFt4IvzRywiyBaU4+AFElWDe3aKkLwGh3iMPdh+RKariG2TqTvNcKQxNjG
KglgaQzzd8cfPucIToARr8FlWNnMupIrl/CatpwF3gtyqM0JMHe3hbH6M9tvB0lG
NsYd4ifYjAOhGjM3j5SAQK9deovRDowJm0rfuauoN8djBLBp8NEr7/c2KTEfr+4l
LBeFPLCpJLeYLSw8AewEycCFXu/fttAW+w8IgMjpeJrZ9+VzyN8r237WOikGKB7m
6Gr8OSrEu4iERA4o+t6MYT2vOf4Cx6S47C/UEkuJpUg+G4xssM4PtDUsBiH1POo5
SLmSgTgO+8q0kkde4B3+stxwc2tueOGUIYB8nYMTZzm/i114tLvuAxKkvW5qRNx9
dOU9FwnBKDObOyHicwaNvUT319GCYwv9LAEWleypi3GLA9XiAzcXYS9Om0fsUwjG
A4qUZS8kYRGW/UpQz5FkmeczGC/SwpXWRWljaHxGLwR1GrznNFbolxxUx/DA6JYI
3UkReDeSsjz8lKtvhg/wtORUERZNB4dL+ZL0fS9wcqblw1N4LF415k8bM/cVbKx+
arhf1HsjnMSZKJibX6UMolxC8iLwQleykf0vxIMYzzkOTZgjphIsaHGm4jXTb+r/
dcJpRhAY1+o6Zgp9qIncK/Iei7+GAUOsvfBfHbmypGlGJeX3tATm+2dhzoOJxWE5
93yj4iV9xu9Z7+/laKVvmQYgfytkp9xJyMWkbDx58wnlTQFW+6/Pie7hECv2zXoB
f+dcbnWGtGXioINROgwTD2LsOHYhTVriq1LvaAFEpIvRh/OeW4wuPcEQmmtE60eh
JOneSdqxLJrIfq+ecG9LmKFU9lvPX6xB9e8ntGi7iQJp/g0q+n3xWExiN6PWnplf
mRSnep2/UmC2Ic7l6x10wC40FXzZ3uuflq0gq7c6YAFCroyolnvEG8zHbntp9YZ5
SZUtsvdDFNAmQ78i6qFleUc3lMUvUcO9Q3dImeoWqYCoQvOtAByqN0TVU769nU3k
1Go6o0Qq+55rxQBX5yAQP+dVA1LVMiC26zetW2i/v8Vz9IP6sETXiuXfZQ3MH6O2
5tMJMl9sHwJZxI+atqozY/76PB8u99rFJ6HO/OsYBdeqme1tNkIZv8UVQXFPjUUw
ZDibhP/zwjiW6397hg1rtyuV7umdaPMFtB22f49zV8e08AJ/ua9ophw9Iuf3GuAE
7Aq3xqF+3kwZBR15UHBhqWjbOp223C0wFZFHPgN4K1fe07Iy2RI9YIKAhn0A+KJV
0QbHI0860wqpjdDvI2sMAABjqHMOXl0RVGokDI2Ol5Q1b0IEfRdA5/8pTFz5QbLv
IV1Z+RSnuPPtLMgiJkyM5a/yUZzALG25VRL9I1KgbxZzRfwwve6HvWTleBIgBrou
ow5T7VHBGK26Az3aZesFBywr0/N/4IZ9wr9lRDetleOs1j5iY8fbE6G7wT4cBDi/
9hRgjcJcQ8/xhvKlydP0whEu45cx1l4eYdQA1vkNRvf8GziFAe5XX/p1DVpWKZQt
xto7vpUlG4Bqmyk1aOt6KSnvZjNKACR/116DOSNlyM2cRVTZb0T9WsXZjk3WHYyv
DGQuEbTr/K1WAqigKtxloFL4hK9a+J16wA9/kL+W49kRos5iLI1vGzIqAHcYTaUY
7sm0mhd7vKtVAcBQJwibmy15kbECcRHiikUO4Z9HN0d0NsIOINj3clBoB08/1AMB
2Qf7Q5P9VsGDYYPPXoAdIyo88RBgMRCH5iBEqf7lM+1ZH6bJSGxSiKlo4vYB0QNH
St/KRXx4sWXibSnZM9sfdjstW5JYN6H8wbzMX2Mi3ndEUZpJmgDwjtWme3HC4n2T
gQzxRBXRsu2mgfDkx6KWu8IAe+v1GYLNkSi+gS6BmH7u5JqnmK51m/Dwu3CVWBP3
4yCVYt+WoaZ8XEeZB9ARs7n2VyNGh8XedKNit0kK4MxrL1FuKqOU5+GoO/kw/QCe
c8hpA14iDzoLrByEeNEkxYhqj+9sddM+B4nDaPpR4T1es14k5Rwk/lMMphRtLcPu
He70oXvrfeVcDrdyfdd5Q0Kc8ixbmbXWtn9Yg5O0jyrVzuiG4b/herLMP2Fb07Fg
LOu+uRMmEECbSZaA0wd98m17+QgRF0WNmRqfWGqMlxXVkfieLH0YkCA4ohtT4SNX
8eubvARuC+ta6T/MFXuUk65y+5q4mM4HQ4wKRccrWmQ9KiBq0hQVP/cGpcC9ifD/
Q8AUWE+iB2PccWnw1Uc03d31XJpDQZTESASesrIy3WSvyX9qssirdiXOoQcXYxm9
ggNIG0hlImQEcBObLBHk5eSXDMzDUB4RrauxVkx6GAShwErCk9LYl6LokSYybfkh
fNLppI8092UwgCG1uPS4ACiKCP7hmn/Pq+sKpw7YkeDJBubnboSnPjDqV+V4Rq3X
fJh5lvqb6N9sn2qSOvxZ4X+cHua6Cn0UZEmAoSZb+9E30/ISdfBWpPhIwo34GKLs
AMH0mDGSzN3N5ZOK/cxn9FQ3NJz0dLGCpl6AAQbEe2XehKOOdkj1rFbpXr6nkEqe
qeFq0dyrXXW5tN8rRFkiVf/cIyDUD/xUHrFq6PiWRJbjZY1EqWhWHtjBkNEwxcLv
1zsUEjrDRFSpC3Ct2yru3uLLEPesY9HWTSQq/ukDDthOKIZUhzCQJzACm68AZR2F
Ut1qd/UTpShcXvBNLb4IZZlunUDeaHSzxqjcyyyFhWlkj9+q53u1DYMLut1zhOub
8QU2kDv4Hu5C9L9tbrAWH1obzdLsy6xcfXwlkr3WQGgp+/t4duJbPj4GGF3RYcjX
5G589zWnr8tP+Bge+jSIqGwWvirtLwO7500vY1AdDXeRXLF623Nu+A9CGm9Lu4GV
GBdvMWCyJFLjhhf5PYrql9fG9ycQeBaHDvw/g1C4X2QFqgtaXJ/HMBZEh6CyGYjR
ZSZp+Fi4uuMyVfGxu1quRZlk5UbuC4XKxKzBsc0qeQra7+j0vTQ3uVvNYN1rR0F/
nanQab5U2CU9CjBbtgLSR5p2G656sxQThM+U5Fk7r88MJXehubZ5pY9LkhU0ulk4
OCZvJTrv1q37AlhvJhYZ0Jt7zUv4ogtmlpTXNYNol6rPUCJqNQVjzgAiu57NHCAM
LPwCsGfo4DqRk3YE7kBx/4HKV4myVh8sLj1j2y88wA2cr/wpwz2YyLDKoUGnUgDI
coda5KeiysZwy1ovY4sxR5mUN6ZwqVEBhkUUSzOjtTZBYRKa/bTrpVzhT/GxpfJL
Wg/oDuhJ1k/WLkGoTbtavOyLMCQXg8YY+aGCThNOI92XyBFv48vzJ6jIOKE014As
mpPaM5ZLHve/rN/lvWGVs8cIl9LqM39w/LuCY+AJX7BkyLNWgfaKmfudBeIB2/yu
Ie6i1lPHR7P9jnRTxiAqTuDTgFCuvqR0JPUI1UPI61F3lHZybH/y8yDbw5xbofw0
cGmDS3s1kY8AeLpA/dNfjKMBnxML1b9Ol+3maVnK7w9+P2mxObEP/Zi6++96MaZt
8NGMGwJyEs91lRUY4m+KMAvlN1JapoyyN+yI7Epe5xu/CeZHMsHj/3DzTnT4ahhu
ZrHkqcLzplIEYnkr3vfcF2FWWIftoX07yCT6XabYKedZxIsSsf3Zw7hZrNE2RG9N
dGkZhiPTST5bYsi1dc3m4vKoh0+iOLcPEt/hGPMRygO38eYkigryTn/TFByvl5lt
+clut73upGTIO0kYFgbzqMBxQp+FejgKMMGhcOTO3DPCD7Re1zp4dijv3hOdux7J
5nRsKzp5kq+1hpzfGjduhDB5OKSVdUPDtWaf5H0L6T0DxYqEY/MbCIlWZT8NC7AI
7UWmdA0NkshDBTsqWHGrq4/sPo4iPOjmKUtOqqv0gVKfnegHI7N1s+BHX7gJtlvX
J2oHoYSberfm+a5GOTPpHJreZpleEME4a0wlWvzIw/ajIMZGS0CjTBaVw/yhmNym
pLyJCtt5cBsvk2IVC2KkW7qJgJN9c8YZHEzpSMa8AWEPkT2+PqscViUikbNSUFEK
5jLUWP5wXJAwI35t8riRjMqH+9QtT3M5c3WjuWUQ9rGp2haD+pf4/5eGWVVb+PGm
879u2iYVjETfMHL3LTU4M2DJrxZeZ95mPkeTervZVcaE4VZEgLxQKmxCNpNraEid
NysNu4AFZN1yzVJbEU0bmlQ/K58XL19jkXZo7vqc4keaL7QMhyJ09wYDA0b+i+lk
aU5CaCSmiBYYcwJLoIRo0+nt7N7VK+ae3i34XQsTZIVvB2W29BiO580Wjx9ANjhh
TyPJT9CnCmztXSLWecjGxpLdw0UKSVxbAyqbf62U1KYDyylTa8pO7SGu3xRINGlg
bWo53v/RsyXASzjPlza4Mfa1DlG1Ilad2VaM1If56SdXQnVIaefS7fZg+Z/Vgbhl
nGAQcMONiN3H0+ReEHskY2Uxj5aQ8h5WXtsY/RQqVJbuBZcqZ3+kofZCRcspPwp9
k5DV2Q4S2Ez8Au4rYWPpb23EqDLAmw3s+8e3uWvuwbFUWceKDQjpDj6z8Bb3IVg9
RlABX4Bg//sv7Ue/fpV9efoMPdL6dIE32fTtd0TtM5Iv7w/XJ0OOoipr68B60Sg5
9F5bafDwnOTyaNeeA7CcSKL2tPw/xX3KHEA0XJzIjfnDEQVb72X5m9Gad5a8AQJM
FDiIuVwYFmWG9kUowDJhZiCTQo9WYhJ9f5RiZ6QpPpVkU38GyL+9VkgRgAnEIL2Z
Srxb1uNXXZD7mK0sCfODM87WKPoZFArc+zB03n7v567c9TAF5DvF6QDGI9/3iUvB
WlInAbEVIi3deIo2HwvtDJCKhsJ1XipO5QWhUw2udcur4QxNDwHdXD3kxAgDAlBe
WGCBpn/Inpkhp+H0sYK7Eb9jn/St4dbXsXSrX/sLjKFHrzlE6pSnYIUTh5mi5nF9
rGONAwh3c98ryD40yq3M+Um7WRr00g+ocOJPXKht9TpaUdBBE83iMnonXJ3ZzmgA
rD7bdccb+qKPz86GR5xAUjnxzDkQ01XBjsgEqfEZqlnVwy4uMAXV7e/FjYqXznQb
DWP9SqoqLOt2ocSgEbx9dt/eTZfg1pIT+wt20wjBC9xAJzSZXaFOol4kt+nAYqzv
PcYbuJdFSyyVDHkLw91tz+GJseK2Rt1CbKWXrfRj98XafGyMSCMMIIm/tNNxQvwq
VY0HA2ToHY1Ww7LuupGFPMUHJhUF1WEA1+ku6vn1FFwXTFlQf9EP53fSaPZfXK7u
0JMJX+B0gtWgO9gOMZKuUDoFNiT+V95r8YLyu2pYTM3WsGKki4jtSiodL3oCbIrO
+NIrz51zPDqljv8YPUlLOaD1MbgrWWyUPySeWHq1BwoLuDVRKuuQSgjeCquxWv/O
lxZ7oFJSXGKnw7z7HKhOPGqgULsIu4TDSAJyc34WsgxrzE6VM3jH0gt3us8JB8YZ
bDOGbx+C4MnGp0qK1sZz0FDXwNaw/djdSrbBdiR/GwtMdJ54tCj8JZvYZ1/9VsJh
r8coek1Hio2sknAY82bpfC2o5zV1LIvt9VCEHRjJFUeGyYzFKMULWIie8m1Qb5eZ
c4h5SE/gbCWYfT8bJldueAxwko8kaRDlQ9RXPBoB6AbG8gh3Qce3mYJJBE8i8nM4
/w2k3UdyTfc/yIDuJjRB3XHR0xS12Ku8kvkoOAnm5V2sZsxc4p/1qnPxtnVyCVOT
+K1sQ4dQ83XpJAzMkIWLQxvQvcO1OiL5jKpUw65vlolYQxcnkLbvBKlBX2OzlJjB
bPIlceL82Spht8w3OoqYzuqrZ8O7M/mQ/0GioCQWwjTXEXcb4Y56mUkY2Gp0nZ/k
m/Go2ljeRv78eW9enMnVCJmdnfAnpW+/gWIkwlwvPFS5f5g7CX2dHAqKBKZZTlMS
zBMie3ArccLlyz4+vYZnW2xsxtYeInoBjDBC4Y236feqyVCdjYHZIUU1MEzNv/cp
OjiHAymr0PKOv1HGNJOEJgGw65HUhz4uN3tKpLo+7kcdAZX/fwvkmfzND0AJEDGQ
LQ/q3MFn2ArwBdJXxQCqOJnUQBfbTiXG/VREBAY5LInh6wqYyfqEjENGwmFgyyIx
lFc8DnzRptOHPCn+qSbdNvcxYdDO/9IWSBbF1WEFgMfOhJsrqIi8R2ry17BVfavS
VZ0ycpQKjnGYAx5hRZv8KO52mHlmlL31+lSrI9FIll4U1uIYA3Qy6pUegehGUFpC
0FtiAYzjVDH2x6kmUfmhTrUFUmRVEoOEztqb1YxufW+5pZXFrY6pELOZgB5kB1Uq
AhP7GaTetQBZqWOpPMchlqcBPrLp0YBjcsfGbBy1kIKbpjxAxn3/nKK5Xm+uGbsx
kwdWfDLD2DAysVq/tM9dp/kYIphgmJXFrtayOXo/JDm3qnr/mYWUVuFAzlBZ9Ive
gCkcpLmAPiyyF4/4bFf3/LrGtlF3SV9Zho4X4DGkcKJJa2p3K95ApPOL5GBSHzWB
zJdOxGb4cGDZHXtxiSynWNOwoL8fb3yxDAujINzGuW1O9qPWyJnjciStf40OMeoP
gTZJV0KWAjdAWJpbGz4iMNVfUAViWCipiIf1VSHBRuu3+SrBbs/LF9GYbosieZsY
i3rQBr+UuDsEK0p0pWVdTLCVBeNIEQ7CZyK7/js1eZr0XQFj47/Ykq82jCKY8Hq1
QF32nof8G/ppnLjI5XE4GV6jjB/+RwZBMhOQp2PjsriuERa8sN0oWn1hqYaoEn3n
j5//teKfhdyxajhTq6yzVXT9PvemqHQm8pk6KMEV5zFjg6R/ql2Eaecq9JmtjAvK
lZ46/sJyPlronpzht7VI3j4/fiDShx4LtrmKMgQCjUigfLt9/v6a+Mop8JAUZ+lw
qZEJeBginogW1yJeOHb1K1cAU258UuJGDWGnNGwcSeVvDceJzXq1VDO7ISJSKana
/nFbAZkq+klCacoTyUdpqpVf5tYsH20RUEZtArmyHoZlooAf9qu57JP1WvWJ0YIs
0/q4M25R3yqwVL8DoTrkb7o/yoKCIYoUGSUevAxOtkTb3tYbdrcQq4kLo9f1PeDd
9P5EvVD3yPbCmj4+EokpfcZ2wUW/d+/e0bq29HVWX3lYYh0YTikEMp9gNRx89l0z
qgu3BF3S/piVutdYieHGo9Peve5CYmmFqddjMtn7xdEiBilfwf9goMOILnnMH9h4
VgQ9xBk6rBb9q/sYociNR9gNmV5QKhKFz0mQCm7IdyeMVnYESKrxZJSPZ6I3+zrs
Jz+tEh527O5z3GxgEf1fBJzhX2KQIu2nj2uho0+C4eYSRZhXaJgBEYmflD/KKnho
jzndRvpjmkohlrZSDzCCz7Vhc+zVyzYidjh/nY4NOywg12kyZZHEDeBDO+7CFTJ4
MZumKoiKraSw417EBrro3V2aUponjD7bpxndj2UgR+Y+tYpTq2F+TN8Payjt0l6V
fGSt9xiapVFJDvso6naSMZyD8iQBvMOa1Ol5PXTgSMeTKjBLKU8hQujZzoob5Ifa
z70lXfBBrGyOlhPre3zTnpyU02urz+JtUThS1gleDjSabk+Q5Fk2bFdjOcJQuCSU
aHRAy1ClDCmgG9Rq35Ej4DFJ7voY57eIstz2mIdTdwgjHLUHBOdjaxWT/zqRvSPC
eiDwcfayzXKLUYTzdU5sfFfd9N5UDKGhtVZa2Rr5K2pLKDuZO10Z9mQL/dQyNzza
s2re1f6qsMzQTMtwDZSqgtwXGJ34vjnehxlDkTKZ3DyuVg74o2WVC2B4eKWq8ziA
gq6SSCjiVsjyy4QF+DlPiDhxJ3T6HgSLxbvhMN3zrMiFsL9H2zI4xaioBsadgYtR
cmnGlpIqbjgwkFy0L8z5B8AbAmva0j64H2avjvCNTs/qvdidQeRKxRQ3Q6hG0+ci
zsqeuLoLVyvULrDMblEQjRknuuRRVGKbIa6CeSE5ig9qgkkueZXgamM2HnjdoPfJ
ct005hpY+5GaFXle26lCc8ZbBA8FG97NU/q565I1k68VLva/kHstVUAtCGZxQnFh
ymxupy6ug/B3jVDflQUEahGJ0r1MgMnl5WWFb5JqSfDyLTDqWCNQlmP9YtKIjnoG
6B1Kfyd3PN0sBDOKwZIIc32+IBqclO28sw4lSJn1m9+XTb+GFVe1pJOOk9lACsOY
utlGkO4g7rbewBN4NlGUid1/0QfwRngHvcRIUz4wPnravhwQCZDp8HqmfIM5doEZ
dTQsUgzKJ/E+n8wbGKjuoApkoCgHzpKwHgAk1iLWLq/U96dgDf2Lp7oG00aME6Nu
NrGBlGLcIL0oeEdjvSLxi1joBjk0teA/qoHZQY+yfQ3St3hKsrCJVxyPmsoQrWTQ
9n2puTxu1g11ApWgkmwZcz+CdYgMgaX+15MuEb4YhZOnJc6iDASsZi3vwU5lLJTK
+Y82dRPsgfuEIzIBtG8kkgUbXSiVvxH9XmnhrtQSTmcy+L9y546olGPnPLElF+nQ
DLpQL8SV90rH9V3vXD6DDS64YVvue8lXr3hy34mBABY+Uzo8oMZemrej9ilm2R5R
YVYJFq+HfUQ4zspQz+dylP5FUwciJ5wt2bbRlPS0m7afac7Tnstgy72ajaJlq2Lm
cc55RoGjSCCgVdnD5hcbnlRPnI5JN/oWbivCudiDlC81P1+tLkMJt065N/IeOXMs
sP3ki0YfeL2FI77eER7No8AlpyetQ0suolALGepKM7+sgI+E1s4mLoTL489ftVmn
YdkeSeZ+dcrT+CkGDzHqFQse1FiYJ1E1gLM7U0U3k8uUT2zGUbKJArvN3gNmva8E
jRmw2thr0JGMmSEUhmIXTj/apmKnMOeuDjbubreOOHjmUJSxZeFTdkkNUC98zx1e
RxCNEyOyvwhwfPxkGKo0dC6m/gxbNrO2fZDACQKS2U0g9rnNUZ8v2c5KtSTgZ3bC
Ld0dE583OGCdNNnXkQJC7mb2kqtLGTH75rdqBjkXUqSPSMtkhKEG8Oeim7RU1Lfa
Sbgu17IDP/25tW8rW8SKMQJAmUwA/nhCreSGAFB+bJi/o9NKrYcWbNPLyKB8T/CV
21+QK4N9FTTSKs/Z84XUnHB19NxQ32XLLs5Zfx7490cDODvREweqG7jLPR3qzuZF
AasfnW4VfyxEt4PPhX+uwnphCfvwf6yjsK6/l34MZriGq0XUX42QQ52WHT5K23xV
NF8Ktuz3Rpxf72Q2g+072riaZvJrcoyH+/GTgeqd6gpaAxql0ZG0KxKdPkokyoOf
X+HcnnO6AHub07gMdmgRgCZjygrafdvOmQWd2NQpT798eUdnY3mGnrHjk9na32KR
5ubOEu9JzrUTWkiKhcNr5+Ku/M/XwyM7aH3JeS4TIQH2SPV9MaSrorONbKLXiM9O
LVpohDx2GgLccqsyxpZ5zsqsZTYFv1UAHRKYYb3yyAGTtTMucxOXjHZiFip6fKKL
K2cmm/gCxLUvH7nqct8n2q3bPa1JZMJ0wp14Xt3O2ZZM1NUvi2jl3kFjfnpzD9/c
klUcC2r4opnzoupg9XR051na5BSRKQSFEVl/FzepdPKTXnSP9suIO3ZBMy8n7thj
HBeHPAe0gDcN5osn5R5vSqiKXI6q1NhJ23zcnK5fJvTix/XHYK8PPqsr5JFXnWXI
gY8aIiCaAaiOOtJWrsi39zBqj4t9YWztyUCaFQ+q/t7R+evBxP70ppTGr6vylhQr
jMVnU/KTRO3pcBfk99uIblSTPU9slToN9ceKy9FatZnY9s8yufJfO+FD5YYYJ6hn
lZycLhoG4hbeOgJntPTG8Dzf1HQpKeLPg/y7pivM+mytmE/n8/o7BJk1go9Z19D6
PoOq8sjbd0vI8hplWszNOtUah2fnTWzBy2h4H35q3M/YeORvaSU5hnCkvT6kwxRV
4kzGmJ6b34g6PxlR5d3BiaVAs2iKLH49MW5uUiBKFitYfFNnOW1wJRSlqCmmj7d4
qmX9LCmyBz3NouJIXcf63xiXl/SCzXJD/YspKvlQzvPauBGYsWURXaGjMfb2w53C
lsZdkexFgp2byQnUXCbPh61pQuT8+60fdY1zUy6eLtlReWgJatVK4MH+PzPjr4P+
5vETjBj8Qfeen+ZOehF+VSn+085gpBNVaR2NFNQwbebxyB3HqM6V1kCe0mE+7eh5
F6hIYXDxKrFmHPTAernZd9VxfVV4lF5ceLxrKFKnZZqa9F2iJ3HRJnF7QWy1IYIB
bu8kccKSGiUkyayEh158ROHz61MPMYMd4afatG4wGCB1ynDRXOI60JsXpg9gMcW2
5XBoubTzkdW6tK3MLV3CRq0NWcGaVfw6HYSKB2Qgd8H5Sn9zgWRmV9yVPS3luCUF
tlyGGp5H+6UWg90mkWOQ3y3fweInvGkBtYLLIubvFjp+62droiSxctlZa6JLDn6V
BRFInWUHoKWGatq++3TYBksJ/hMZoVrVab/6JHys8zaIbpRAYW3xP73m169341O1
MIknejtIGChfjk+jjAq2pUF4S1O4akpJOXgRmZk1bB37Wu19PeDIh+5UZ9COjPbg
lk61rgU7lB3ZAjADCW1W2RmXDsCesSZAWvAS6i/Cw8Ii55Gen0qo33uFTFUgTalI
dLxJGmix1FJPAybARimW/miX5kG+jU40UC7XR2BWtaOs1vY77tdhc9dAUiLLddEo
PCsM4/dNlRIuDx1dgbfXvs8dKM7Of7rRRvMrI/9MA/JkxWcb1V/3teRccJNo+ESg
hya5uHy1/4W0ckuWNgcF8Ngd/AlhenHK2CY/IAK72yCDnkQb3qkAymlZeH4LY8y+
5vpgbpcA2CsEVJeV321PmuYROXcPgKtzWxcJZQsz41VEWssWvxgyfCTwmg6QnGaF
PC6kdnYCUfx/JixY1c3fkAn4USTYw/zBZsyf0N0pjYqXU/idx0pvx4mOAWNM+HVI
iSMZnrEYZ5FSd7wO1iaG51nlhig2IYk0NuZWNqFMwYP05/N3ptJgOXdXIP4lhKQk
9k8CzC+0XQtwKjTihco0FB49OjTGUd99poGN3FhoD9gs0Q5uctusf/mW1MfcUEsq
Js//9PzXTfPWvvXB3hmgTD+WGohgFcbmcyJkQtl2vd4Vr5TxjkZYjyuAIHNtMvX0
+JZUG+EyL7zPUG328ybmqPfv3hG8dvf+m7i4bspXRcPxYnHozUztk8cFYBW5bhR2
Z/qlxWJ7GInsj70L1PW74xHEJn6BG1QyZFmnX6/jjnXoCKnokq9mgq4mxhVeayZV
2wyjlerNSNdwrGlmJjXJACbFAU5zXa8s2yuF8dnvd8yFzB6tJe/wqC731sTiDlk0
fFDKC/6ja02O+4vIMCfyfdvyl8q1S3y3q/WCMfvI5dAxR5o3sT+1ReYkRiY6q0dQ
JtliuYduDRzpAHNYXpc2ts4M8X93o9KZm2SJryjCnHfJnIkrdCAUBlPe27Wzo/n0
pjc+AS4vD8CV3DmFY+628dXr/cJrzBTmVfGymlDntLi3As21KYlP4kioyZe/YCuz
sNLGjJWAnQ9ULWtstdxontYaWAnb3ahIJhEfXckAJb+1hXXqWc50XByV2CM99yx3
yuozPT5oScovnzA6+c4WVAsL4zPJF+Z/oWvM/s+Dw5ByxW3qSV1MuGzBRjKcn+KS
2auuO+7/Hx9HMCPOMRKaWsMCYPWvWp1ltVkEnLTMFl1/nZ661fKI8Il4BR/BPSBK
bZH+e0/eu9es3F+7tg/N5MVo3OUri1EZEHVlxF6oUg8f+RP/yLoGLmcRMVJSz1pY
W+gvc4hDIhy/W0cI1xsnwemcEtrKTiudJgjsTt1UzKE6+kAT9+lZTYDMDXEpfJlF
r+PV3/kjbiuSS6hzof8gRtWr/uf9/JKbyl2nGbvwMMOsUIKKJXC4a2WZ+2zq0bpJ
AFEshJcK9fGVz0evOpjAP6p6PjwIrrrW/VkRgCGcwB36j0Ao6HArtoXdWO+uQu0t
vmxkLNthoJ7BBYKsBGRMYL/Utky4RTsgweipVVbxgT1CQM/Ub7M/A75jjZyDm6P/
HRb5ZX9HxZh+MJaecZRUdRMIck+ell198ouNAPMrlHfclDis8ZhOEtivwYkZOmFh
+eO1/qbDUSUBpEZhHl+DIYL1HeHB+rYhMavTJMPORTBqA1Zro7giHtoYJK6BX19u
KDEUlnkmMe+3Acu2y0ShL8cV/ga8NHAVavq5QHqS6rqHy58NlbOMNHQWfKjMMFxz
G7BLV1fQsm+aDz9JO7Bs2TvAl0Cb1+8zi1tAhSlwY4+A/BMZ0+94ct6OjYwTMyyE
7ITBs4Fr2Hmr54YO8kvwkS8AYgre8rk5A5v3wtbksljE1YrYgtT0JSJMTFm96jkm
oDRsHOt1Mm8NxzAtbPWkEsptuVTpGAiw46dL2he/HR/4lTsoQjvgjiADwEnXO4lS
Fkvan8PY7e+lxdr2DCKz5K3L5GVEcDyWpbxZxbtYBdH2sqtUuzbHHty2oF3kqC4B
qBbDu82vvnMO0yDcTDIhf3LwXCYgRgvdN5J7jDX03Aq9KCS9IZpfaSVfh4hPLNT4
g+DLCP5nvyOlFWWZ6kalkuzCV9x61sMjCnYq4Y2Gk0qqMEO/tgt7bkkTgFPsEiJ8
4G2EYcSFNxsZjjLes+9MyoSndZqP5e6/GmH8Nnd2EJAjW74Me1yI49VZXxQKOWfL
u+qbw2+lg8/JaMZd5Zn4bODJ1i9rO9cxL5cMfV1c2mBqnA0B9uHeNEjR/Tnw7bci
IoQjMOIGiNO7khCi578tDCPdtqLYxhvYBZTHW2YIszi1xArJ86dO7wLhc5Rxv9BJ
99f2rtYTu0jbpNy/bHwVBMwBJUOCdrAh+FUPeaVllAKzeTWJP12aQTqpxUdQGQY7
csymfpYh5hbdIj6YMDQvgs1mLC4NQAMZDGdWbffIiD2v9A7rL1sdLrPSY81WyjL9
DF8Xvi47QnjKVDY2SeM0ADVtP2vKpjGy2TM3Wgd7hWmqeoWPpZ5kv3DeKIvWZGOX
fB4NU42syI9myK6BYIPt81zof1ZjvviozBOpw4VPXr9+j2Z10gXzBzq/Kt5twCOR
5WfLoUPDipwBKovFC3+i4Xy5Sa0POClv9HZ8PQqJHwKa1fns6oSQ+5Uf1bsZ+gtj
MzMHNQM+7AB39DJ7aE21qENvsomA07RSbFym42YX83mIn9FipFHrkRe0ihGlbzR3
JipThjA8/HcaGNbsRoiYcNVpyT9LCmyLwMJCeJw0jbEBiCBDmt7cEW/BEVr8eM4q
mIJNZdHqCrwFQ0HpapiPuuWzqpu/6+pe4g8YooqptCqHLCn4CPd8Co7o2zwgyWaN
6/hOXYWfakYszlZ2wALLmmm21rwFJOEnQsFd/+fjcPYYvYlOvwGKGQ07YVFpceBB
zAKjQWXxRycEvutssp7IRMVcrIMhgPpUfBf8FaQ0wIqhj2zgJkLPstGdsCO7rE1W
otTLMFZbTQYDZ+ALyEHZOk58JOQ7+7vGSPfzXy1XAD07e5/5nP7aTkbfW6UNJOtV
v0f7kS5azQVeEE3RsebqZrHnsZILIPs9+oMPnKx57yIIHXwGFXJJaw6phaMlQ7lJ
KN/t6rBDVqrL6WuRcZRsoagUQpD9vX/JV2vy/4UofBlBr7x6Wc1IlqGEIJRiLGf4
fhteirlm3N+Zw9BgQ329qeG63Mj4dRXsK2tkw1k0EA11BGIN8Trgg1Wk/0ot2aPW
xgB5IK3Pzm0oqcKqXCde9ojaItSucLOyirq0bR4PY8jdB/y94pnOJPnJDIDmxY25
riYvlxW0W+nK762FC1a0eYbaPL4QQiqwey+GvJ6ssZAVfstnZdw6iDDXeyxHQV07
fxCnseg7ZwMcCi87fTJ3sMRwqJ2lh7TM/RBzVJ1qlV4duJ1OtwjfUtVAZHvDlUum
DEO3mRxzfAy4I1M/Kjt7NglT3i4keCmWVv//OOT9jqczHqXkCu2jWweQs07QCgh+
Fn4mVHiB6AksCbRSrGDZ9UTsGBGDDRm0ds2yoeGeR3RJxlLWuC40VOv8PrVv6gu+
5FKf212yVodXKj/i7nsBHjOrJMtNCWu0vYOes3+bYrQMS/JPIBPZj9WzoGt670wf
kQzl4GW7RSi885Zs0Y5/QAJi3UVumG2AVcQ+q/5IxRUHxQCJepgGz8UCx32APoDD
XTavPG7366AUTdyV4o3JWAekUqVC37yM+33hN1a/xXmkuborwXMt1PM4xIPFl58u
O9iHCQmu6lYJc62jLGZppAOdBU6bIvi6nYU5WxycC5+UP83P4aja4yelrW86KOme
qt4h3EakiK+p1m9aUK2eqG+DBd4YWEZcjBE0BEQwiNNhoj6s12vFPgOh+sAwkIfS
lR7PG6dFlcSJq49pXIlKBzR2ip27BF3Q29m0JxRfcu0QVw6gklQ7+xVURvBiTXtB
vFD8YvEPNLJz60puFzgRxGDl2D6f55lTxmVL7hcM+dLEmAgmrqL86Kw6ydKjDTQb
CZRbaqQNgYMVy7oRFnwW8tu+JPVEDYdi4e2wQ/JEFuNQwupRKFLRRzrYp8B5CrKU
PmHCkjE7R8wdZde8LF2W0ZwXHWnEPtOB5rgD4crFTdjUpq4wLNex0u8mzgoPWTxP
QcpeNBlgIyIBnCj9bs4vUhon2kHUH4OEYAXihOCR7xeZuDBLpCODzU6fyrY6Q9ac
Ph38p9T1Je9TBLVMS8QvhQAowuD7IobhUfYghn2ePAVEmuuKrMtlY3xDVEofaYco
HU7O/4AOcHN0EhUz7B5EoNHyzCmsTLK98tc0XWZ+O284XRwry6yhqOLN74i42kHG
JZG22PBD5DRaK2r8eM1gycMwGMHH8M+De4ne8KUG5Mbo+kcnPnV8580noE8B7aHa
AGBk3MCeREcysYTELDt5KEmZNQ85oMqg1nJiEt1qNZplK2YDyn75yxX5KW5TYKnt
NllFijTWIulBE6OdUP/BZPS7tk424VAlpy6RCcpERrZljIfgUNA5ZwQKXv2MiW04
hzjgxThA+UkBoEc8wUNo0cZP8yQTPijFks/QAufLl+/2P2Tojwxh1GxISazh7rlO
woKojBNJMIB/fiLIPd834ChGuM7rJoZAseDyxoenTgxMKemEf/dl49QCkMQge9Ya
5mkW1Q9sydO+fQ+VdtO9+TIR6QZCR2sBaxfSgosaTTp1CpD3mXnBskq2S7AFzl7G
lrRZW+ezM7r7heunZDFh3lbMppyCyNlG62YUZRRllkOzZf7JxZ4wRsYX64r8F+6g
ksyZzuHcNCIZCAEcefbePvh+IZKpA8uuGASG7V2TVY8Cqylp8E2pQxd1wbJnooOC
wG9249vwOzVrsTY2GGHIRfLYmsxGCe4HP8JiZuJ6VQa56uId2lA8DksgsEuVbTuG
J/+Bg6dOhWrR2q28rAknAfmyjGdR5HO/q91/BfLtR8VhxeawuvbdNwvWqY4pAgtZ
hYGzOu1GNcPzrzhfUB+tuXlWmkd1KqJe9PCCsoF9a7voMTCTSOfTuMAWBBFk/FUx
Cg4DM7o1Ajh76Q0UlsrnSIEL/pKnAq9C75PPqvjOcUSm0GaJL3mpiCnZT6XdsDK7
YrQZkTU9DPutOmshu7RA9MfB2O1dn0nuiyC3V22x/cHtZKzCPbcqYr6n/Ta28o4T
HWyEsIkS5RVdfKw7Lee1xpHZgG7WHkCGKbXoR+7J+ScTvQlnxgRGHinYzsb3R89Q
MxLXUvFAsKoY46nMCmxvN18aaBU1O5d5yEEfTozGFr/En7FkWofIpPWnzLDNQ134
I8mgSjEUUz4a10U1QbH8M8M9cdLnN+eLX7CuZHLshpRu3UEQj+oGk3cig0HkSXQW
VF5hW1OJVNOOHKsLLMyrRXMWPv0V6RWsMjRiBegOGlP3kM6irYj0JuJ7VWPP185r
OxBZo/O9CQhIbENaKbFxtynE7LC2WDd/1UgavDxFwyhdThLK7KW3Ng9NsN73udwS
JRll4qKMlLV0XqhoS/lZhehJ+GbNsDJf1No1VnOtTo6haTCt5c97KB2Wd1ONgufN
zq1xIeLIjHBv5VWjIoTCg0vZSk3jATgqJaibnVZke2MdslQdBh0oKaiYyE1Wh5ge
hoLX2f6sggbk5lPaFgUaH1sGlYOeH/D1+txKzaC1jRu8vv5CMVPrVIjGaSYs/8Ai
VBO8ZT2BZ4pYYJCWiSIQPgB80/Qpm89VxPw38wRQE9FrlMDsUlz0fRmgoiLE3Mzu
mEqWyQlJ5W6+A1ib+4179lhB9BGTJkHIofwRsdS9u9jKrSursr2emJcrw61Xo+jc
AzQR5wl7JTfD3ZCMOvJIqOVjDjspLueWgto3DvjFsKnyl0BddBveiy8EwjOA4/wc
os8N3Zg+dWzqVSUnMwjFpXCHB12aoBKyb+NGNU70VdsltzGYbWV9Fwpnfsj33J7D
LBvdbe9zqHe1AEvsQTYTvCyC3rvL/cbx4QSTzK3rK5Xt8goFzggVtceWtOCxeiUu
E5/Xd95SB/PfbgEADRkVSQUvS+8IfSFmwtkLgXpYF0AxJ7WJIEj27JThmwkUtYl3
8umKodPsKjSam3SrP1K66CJYGmDnABwdmLFoIGrkcGLPC/92cWpoOIVOzd3mTHgK
jKk0SROFm6ugpxM5NUAAoCKRbF7Y0SJRio++5U5zrS//k4+Zr6OS/gi+z3xIxPar
zEiRb19pGGWrqCG4FQLu96QPtymkeP41pMA020CAGAHuTlcTkcvz9YEYE2RBGS+I
OZmrWWT4jXFRoBXgk0QaC5swbIEq2TiEJagr+Gl2t04qxXaqbGSj4VzT6yOdcmhj
zFZus62RgubwfYfxfyOMRihPkBgeHNXWlCCIS4JuW3KqF3uYGo/gbkcq5wch7CoZ
pwem5s93Fv98uykbdP8nHvw+qhoprh953vaos/KhCf65ucCDMVaJ71Wj3BuU/hXP
BdkBuJWiJTdnJ/ubA8OI/+oIVjhzIz9Ii0MmmWjLFVacXjdeO4/8NERZqXtv2EQL
mfCgvX5GcwNmW2b4LU5ssRI1Alocv8oyRwO8c702LD54lRKJqmx8L5Gwqo2mf/ox
lWTgrnlUwETM28JzyuaiZTNqDrAFN8NR9z3lMwbtU+eC+QSqOELuQwV5/VtybwVH
rQTGVt7ThABVkSvSNEQia19gtiAV+/ZHOvIpk4sAczMyG9gkxXOuuL+f6oMaPMi8
KsfHw4j1t7fD6gFb6aAPmVkpTmIpVX6AQwOjXKeZa6ifeGa69GMSe2h2cQn2Zq9o
GTTXoMiZLSiC6Ok/QKxM+qUpbZ6BnQ3QZKhgRwhVkIR39zuF8t0TvAQapROm4RfC
qv+Ok9wAN7jhXIGfZ4h8lmHusxx4lQP1fRz0wJSikx3ffNhmkjRHgD2sgap5l+yk
kVdIEj3bzFy6wSMVjrrIS7kJtxPD7wNGyPA7T5t3TRhouxNWyAKSgPPr80s7QuZW
ZBFcrTA6qpWaU0nvwjBisN7KTKNjWDLB9rfDR2YtvkWSAZqn0dcGHJHhQUzpKI+W
743g/rXeAbh7/XfmVq0loRdRQ8Za+VCN6rcffn8KHeW7NFCVfe8DKiE+Ekl+kV7E
Oq832Jkn+L8b2sAzLT/68UWrQ/JsanKCU8BDutg4JzvnFW3yZyl/JvRAnkL3uGWZ
2JVc1h/TwG/urH8PUursqLAC4vWYij2lIbbhavDOOk6pQg9B/lYNtpz8HnXhgK1P
n0BucSL7AV1Z4QksaGLT9hJOvXrtAxUjPQECqK2dLVSFQ5VMOE/vNStkzTJ6iDNQ
9c7qyrxkm8S+1hj335AM4+V4mmXe/LUXU8u/d7ws+kh978adWc2xNkYnQqnsURyU
KhZTQXBGI1tUJ/uu2ix7ff13vZ0/4DfXVPqtjI4f3GS8IcYsaf/7R8ZODDsNtkhu
y5WYt0OWSjTa52m9hclqqsVOX4uxJqbq+y4S15du5e6s7BRV1sDFO62UP6rF1FAE
H90yh0mMdc/O3miwwPS7CraUuBrbWjEkHGrElESFPC5JNalvLBGbSuYn+E1qO4bo
+sPeBkZIXYsbpJ51Lng+scAqmkeuNqdttQYfOKSUSJuotG793nNOUIdRP8ZQGvz/
ueal82//guMFLkMdPpVuMY2c/LN1aZP4E5Noom6MkuiAw9XCO4MjiH8VBK/Q05wl
6pQF/C3zswR/yEK4ppqCRV4h/J9Dl/13BTug0I4W2HM+R/mNBNQpD0AnUlKEUxpH
9S3nc45gzb3zZRXtPZdtlN8vrNMWkXXqsc4f8IoFdGTLYH+YMKN2iAPKTVq9idWd
ldmSHQT6zZFGwYDPK7jFAPaO/D4tMPU72pgCmRDnW6+0RmLOlisSFMxSpWuph48k
QVpbPEAbkxP4/heqExZEZCqZNT2db9AFSmhUIMw/iJnkKa9DVBZ13eIVnWaB2OJZ
seLPbbQyurR813+BT8U/IZUS5WSG1RWVydu8iEN3cLAOnyayTkWMOyYyYhhZJuM2
byFR/hhZ+tbDHuTDuU1cNIrNkV5B8bN7DtYDg64hwpJCB5aLgGhtiiIvL563EUTD
Ssmey+btgqKtysv980jOj/pk6KUAM9UGuSXP1rfoYelp3MxqGma/AE74P6KWW2fC
UQzsZrJUX8xgM+sl3+2oz/uLfpsAlQ1vGzznqpuP0pu81PLrfQ1keCOip1Upo0sH
U3d7ZTW7kMBDUlvovvjUR7RJk8Qz7mLuFfCN/6lMT9R+YFVLrs2mKWEWCt8Wsp02
LB2JPXMV1Vi3qwvk87nRWa6lxaArbz2mDhkiNdv59JX6UI3QEKg3KT8SgsODpAmE
FLXN6en09llfSURU2oXZjIwW5sUyoNldC+8Tok1Dk705TuPyBwFO9lpcspBEemXv
SCWtQ5kpT+3m7h/SQowqX7v17liSWgX4C2SVMPx1zRMczJwszLg46JgJ19hEik4j
OjWb144Yp+GBViaVgDS9bP1ASemSGEOnWFylThKidLxxK3WDWqKi/ZqooR2kNL9X
FQ9TUhz8XEzyi7zDpLu2cojqY3wZNtLRbAL8+SBO3vpQiJ/goiAIE6CTsDRC1S2a
euOKU00yQBC47yxeWtrN2QAxD6woqnnnlSls8Gw/y42QEqSFg73DQK1rpQ+e1Kdd
Kwc/J3xzdDYh/4msdBirpU+wtKMjBr+5jdqZUpKHskPYb+MKKGSglvK1oWXQwjvc
VED1rlJ44cwXtHn7zHl98nnccU3111HzwGK7SXg1iU5/y5Oz7mT+PtFzdS7Ni0ye
jAh2kEczZzkvsBV0bgltGL1Bj/VlyAmwV1uGRNvqi9a0fymbne0n8z2K0Vsia/RJ
a4CwsIFkGVHz21SVEoIynz4rZ0HUYtAZnpAsc6XQUQVGjEArRM0nsooD5n9Biv/p
dcMI41Nt6KolcuZl6pYQyKTTEEL+e/QD7L7KYIt9PArjyHOOhUay9v3YKBKbaGeU
52JofAN8gFu/wetuMTjNFJAuk+LZ9p1OuMFobO4lJ3XkbBKlBMfw90SqktVKlDfZ
lnbqgWg4FJIGx7TO9N4uy7OEObjDF/QQfCXJB54dOVe4fH70JyeFMHbY863jTYc8
45Jo+wDPicXfCgMsKE+xDgVdOsIEG++U6VMEw0COIBoe8ajrFWHXKs9ngCroeDOy
v96LWxosnaB9XWHFqOaxR4RMYFLHenIvSOB37nhZ6F6seAGE3StVX6LFzprg2L8x
7G3gp4jRYcLMeU1doCz/DPBHRotI9PLkT6zHBCY9L9o6GfsIU0yi8QOYi8fU33eR
w+3kXZia3bI+xXJn98ATPOrmJnHubn50lS8qy8hH2du5sZ1guZHPyHu07MAhnYQR
JIWFdJg+0ZIp+YcFf2BkHeE1o+PmmNWYXSt3lj7RNsCv73tReQ45In3+SfTzeCXd
v5SxeIs4CYPvBV+cdh3ft0ys+EBaFfUU+586MwwK6mxZXKNvaQcj8pCaDnagAkwG
v4HFWJhGKbOKBwBTJWqOvnEGPNB0EEB/YwB3gOyAhlJhCgHuC79DNhoCAVhjQJSE
Ksz6wHWSpzT9f2Lwquk+lJw/FzK+Cd030ctIHM/xpt7y7lBwtDxKethan6djlQ45
vxz3FRmR3qdUn/Nc5jhtcgczJoExXHmbTbWdb0heAjA4nyxf7Psqis0Zv0wQfqSb
BPTwAmrIthq28dgaMfW/aqRkBWFavfbfWGK5Bh7FXlEYg2FNA6J8ZxCJ/qtvjphM
DjpHLm1w6UN0DvWGpmwxemu7PTz29qnMzaMJillBCuxrNBzn5Oa8t47VEu1QYGIj
B/EhacAbtGNbVu0vTbUbeAhLlNLKPUaRV+9cJpAbmQ1m2JsOMyIWATynJ6oDAw4G
xq4ijWy/TtUqNp1ktQQ+8AsLi14M6hDT/2qp7AWOpfkcEkGpjuqbWD1lSdqe4kjJ
c7t6xGM96+uytEGyr8vaZIJbGkAYblYgJbt+lW44w6xB5v23GrH7nuOeQbXMElRs
44gq7JAZoNHRc+fP3z0C8ji83v01M5+RLkW9KFVR0GuskqAUsyMT7tBKT/SrP2b+
y7QGkcVUln9Uq2mGcWxZu5cu4ICrsv2rMmbyzvdaBbk90ZstsRsSjwVQ1waM1L70
5wtJ6IRcoWWxkVLS8NoSF1EyK2fstv91vsMvLqX+5J/Xe0bIgELLSHZRLqAL/wCQ
pFdEySphV1M+XKTB7mI+5vqPgLMcVltxuRGJM5jnIGR+NHsiZ7VxW2FR7jDGYXnV
qnm1H4e9wBht7JF4RRrgLyq8nHSyyybuVwsjzaexZUEP8tfeucr1IOTt0hEoX8J+
0xWITu+8/UXL0Mb9gFYekoVBExFVp7gjm2+hiEl3Pvs7hSswuADROolad8H0bRhv
Bqr0J1vKFBJlbdJpOBe7bhrtFosM4jHq5VFT+PBn1P61GGZmYiNKP7ZB6sUuCCSO
wyfRFjEummDuUSLaFcaTuLZ6BbyQO9r6OzaIaxWs+RFX/BBEO1qs3SoSXhAwU+s7
xuOq1nlCJXerRDW94KYqIgxi6WGcEHuPUpSkjkt0ai24qhUhSEQj54SE+ETQRF6R
9NTcSxV9q1o9XrPRIE2y0Te4nFlQnqCk9LrtEfk7w7mkt6YqQvTzvnDpDr3NPiRh
GMokprkpYjaHLTtx1T8xKR8Qg6jcpXtJXVBYQuXgnbyoSMcDWpH9TRBP2cnMMVYD
t9IA4gisrt0KXgVv+59NCRt3DBlQb1Gus/CipY/H4cM0zAmwUkraanZ5LVAd9p4g
TUxqU7XnogCzdIbyenik4KtmuPz2ZsGJz1CDN8DqxWcHMgSGkEdasruKvhF0nsnE
fpzZdlhSbSugrdnK3Qpk62/bI2NRT0xElOJKbwJdCM859GAkr7Um06fALW1F1WGW
V0YKj+eOmxFs37x2fyqSpJfgrxewULhCaWJ90GkdUGSBkDoenySgJkrIVduqJABL
yrYnW1jA4Xh4RcHKOlV1MZtUVS7imyM+dWd/YDn+J9mIF0W9+8x2jOfccuZGFlRm
tMkIpiMZwAnQ6/11wfne1ydGMCbWOJAv5ciqY6UKFZUts2F6G+lXJObjcHbrwdst
Cyhex+pxM15eln/vn3fMuodUOmWMM1pfM76bEYxskqRvxx4uFwyRaLZQfI4IjogG
lJeINK9nkVXU1Wax/+pbOZxsiMCwTdjaki591uBP4UlSqi4EqqL4YR6U3i1vtBNY
t4rQTO5o44VTByxJ7d3ZUInc5OTx4bqlAnvP4dM1uyc7JREqk6vMwt3CvgmJbUsB
hajyPOjJDumNBFonBUlpbCsG79mIAAn+lD12rNt0OcVwYvUNhYbimenzZiFPYh8T
fUKTLjw4qD/8On4rgkQI+2Y23EoH6hQ2qGAyekbFCJdC4H+4Cb6NT2ZwfESvMZ6J
9pL4IvNmfJ7zqM287+b/aB3x4ezfPmZ+I+REUh/2mUlHPwx6kLhdLPrxOQUnpcCz
XBYt+Cf4iQ36iE5lDr1tt+XcaMR7Z5LAnQi9ArmRqodDx47Q0eXsyNL9VkPtyLdc
sUUbVh5kSIuTdouBy3xVqy9Lvhx74tvsJjFmLknmDfWfTrz6s1pT9RgPUibVxSB1
Azlc5vL1Q4Pbtltd50dPA1xe5sc0xx8u9fuPKo9izobYZ5/jKf2lSvdswzLzTh4G
1azgZP1cD90ZqhI/dbryJ0MG9rWG8R+r+RcigBsI0ALhzty2HIXfJ7Y2p/X7ih/Z
97kt+JgNv6uL0dONMS+MrKW1EGZqnjQ/XzY6+NIQb50CYtYHrVgLKbVzMwlfXCZn
T82YCOE5YMNgGMocoW4wYk7kAqfO9dOqHB/C1BSI3b+9jNTQKn+k5AwihNBJwPpt
rLEAL0KWYYndMfz8Cz7Zprt1hDqZTRMEqIXEOA3A/W7fWNKlnxFtOCXPNu/RwJIo
67JLKx7hbn40Zp0GN1y1mhdSLCoTWSlj9nW65OLedDFIKKSBtafyo7CLbg+L8uJk
6LAmGAt9fLIYjHN1HVhXXJwKwhRkdwl3/Me26v2+RqXenciRqwbwPvtNxX0n9QIv
gA8TrR0GEUt8+6gqTPZ70fuyMkjTAGpA4hpITbnafgbZFY6osHP7OfB/n/lyuF+b
XkgtcXVNG0B0uvANMCdXckStUYp8qLI+wOhfvO1AifI943QzPgIr9v802qvmHjEN
hbZR4VXggS5PgE/yDGV4Q6uBM5ZDa2lNU7nL0huNhbGPL6uAK9YjnsgfMMHJfVFm
n3zmDKWjVxO6t5+sOAUtFf0BLemYvsDm6I5FCivDxOWz8ibsPUq3vMiBLMri2uY6
mQ67AZKDkdwN9YMKGN+oCx5yMockYVAbcQcskXvkBVLFtvHcBOQmgyT2kONtqacv
lecTG8RrQMoPkXdxEjClHRmz9KV5NnPdFScecCLSiijyHTAGBX1HNAzy9dG4WBrt
6Tk2HSF6yCO1eJM8qQ/gpFVvT6qIyA2Ju/I7M+LCTshpXwWTQCprsBtaq8nxx+DW
UbV+nkgsIHAf6lknPvc3w4qPgcFd40Px1z68/rKEC6zIZcvnkTmx7SbApCrTkTTn
KtIRcvEcReQQVXecTY+86nPoCwHNieTt9xRErf8H45KV3JhgUUPkuOxR6CezoIQp
oxmpm0cDFq+1B/QX24d+vQmTXTNx+fjl+uBlruCFMRL9PZEjK+4FrTU+kQLO6FA8
yLeq1B8P77lo+cEuR1EbPiIdt7hs2C8Ia52LxYkXgVuaXqX6kbqfv4SG7p9qBD/5
l8Cdc8zayV565bGQttnOlPpeAu0QLy3Ge0GXNrE6KP7ugdzPRSeFvnmU4BCDHZwJ
m6d3TI634ukg0UZPAO3GzZASuqfZGs8ovygQwBf92olDLY3COF46gqCT8AJ7DXzX
tmFF4V0YucYLIgay/LRPgujyUo8ZCQ9wvOpXQFjpega82M4NBUXeyXnOX2bp5hKE
WIB6a8+F7AkiuULTl5LmgJFLNSGx5nkeS/kNTNxjI+gfq4rN96e9xn0/D900FbGD
ysJ8O3CQkOgPnaMxSu4QrAkEw5b2IHom/IPQlPI9b1cwFA3qsqQI5Mkfv5ByY022
WSIKnig4QjQgGDvt7uv0xpZPnjuNi95je8OcXEZwVKI8qcKsenj3OxfPdX9ozjBa
nGOmCVkS+GAsZN7axjo/fndNvC8NES6mqyG4qLEsrs3Vzl9bqqBR5YSMZhfOqLLj
ZmvZspAsZhOv/VtkCswBRkMfwpPw+Rd3oHCmA2nEPwB4rluHOqxSOBdFDUi46dZg
E2LUg5wYUtqEtzwbH2vcDX0F96xJE+VMtoR3pefrHGbQBjJO7SXaGmIOaJdLsB/R
tJnBqEbGTcQGQkDcAZaqyMRJh4lAI1ZZmTrdDeYkKltTvkj66y/B+vJNvq2MCv/x
I/DWUeXqtUMfKsMQjjHiQmCdYzdIPGyxD4veUjSBfqBMKL54EDyua2INyk9wBOrG
EkRYoGvXau2Sx4aPe+8hKW3mr+p9eMR9ncLsd8B3aeryX9YiABS4QLGee2en64/c
pi6URc/+8rxT9cmPbd0tenBt0WYDVGvixTv4ZYFGKrWwaT7/JonfHjlfaIfFgynr
GJl9oIAw2ozSjyo4Gt+4HpgqqYVZ8kl5NUe0USBRVWfWvpWDQdm97Bj4e6L6Nsb4
zYDUyb20ykeGSUHvwL3nS4cqiZHTrjhg7Nv2cCCVxq5KiLNCzv+jUudYSUjkonfu
ekxnKMvfA8exE3rbi5rmhvnKzYIwMrbHLL2DP2Jq81zcswg7ivL2RsTmliXCoJ8n
CJRH3cOiHuQ0agW18DDwtq9a4F7wGfHM3O/IJpO+4ok3OXmdyqQxbzuMqj1o1BjT
ZoFYOSK2Kc5b/6cRi1xBH8MxQNQTlj/PMqsDT3f9OZ79WkuK00LNEhIOMpxiCD8Y
TglK7Z9BCRvlrwHEZWtuF0EdnhuTkez7CiDlMrjvzQ2WMWDDZ/gxZDuuguKrsFgy
iryNYwbrhR43Drtu/2KR+BCUAzZNKr2y81bxI1cLaYJShhHkLiB7ydzYUFpFs3L2
fAA5HG2Z3mi0jPIiqgIHs3qAJlQhI1goOgoIqN4xOkf5HNqRtGLWOdPVfE1riEO6
qkFWQQsNyxSS6z/v2UKUb6ZLG94sU4nBJ+RcSd9wrLS8BH6lnpS0QYjl5DM5xDWW
bgJEa8c4sXBImDZZoHf0wrfitxWwVKtHDn9CMnAHQ2gToWDTNssr8wD6ioBMR1wb
G8FbqMuLVI8WL2QKcMTxIRB2Rngr3lJKJu4sEY8yl9YQUy0NGnAcUzmD6M249fNh
x2+GhvIbyi6qrdtmnWlZswO+UMH1LZR3s9yYYvcdLyULCUFiXmGHz6qpQs+iMFj1
h9b9r9q2Tlo61KSxMDRuKalIs+yaAQhVE2nM8VSXToMI81uQnTOK3yDD8JZhpNiz
TxZsWr/q3dhkG/mjVMF8rXIwYbSFp1lH8bIvpHcSr2ZejDwE6aQ1ci8vG1iRi2xw
oXoU/qI13VVW49KsKj85IhMIli5fL0oFSkS10B8W6+NivKCQsneddangVWNCV73l
L4450UWJXaPaIonosqfaE89sjkMiE0EF3aL0dwwDPnD8q8951IccPZtcT7VncNwM
HxRRrmY7IsnVUE282yFp5hzH4T/uGeoDtfwuQ38PVoUyU+1cjc9hfPbsXVKWBl+1
uaqQGvPVBuE+jJLIYQuUCzHNv7CTkludOjMcgkhDB8cQT0ts3EWtLbGWzTYtqz0E
t69cm45OWY6O6+zdtqEkIKdRt+fpL5PMQNo3IK7C65vehCd+KMOjSSI/3i/ewj9k
5eeE0HoEpgkpEekLMmfNpxrJFGLa8Du2kCpBOVlzKk8B2CEmezGRSlLfzlS6tkaz
56JsfIyxzu5WaVMJpXdAiQoA5IrCZxCcUaHsMsCeS27z5q5NNd8W+EQPFhN4XfpK
KDpVRWi9iXHE7aUwS+/djBJ10/5VMna4a6m+lTpTU1o+oumc8vwRCtobylqBTD1U
dFXhwc4ECLPRjk1mqlJa4q6pzLuJCsFgLkhTuMixjcpsLA07Jqozj0gHtAc3Z6E7
5Z3dxz1R/MTDxuxT05zdFZREYolDECjTM58ltCaJuWgSjn70/898C4/NP3htVX4l
Wc6RVLrqlwZK4PQrfE4YcmKPvZJ87HB30j20tUSi5Rq4M7A2CTbtZLM8dTOrF8Wz
dGiHsLt3rr8fVMKDN6mnN+U+3bQH9xy5pLSO/FW57UEaFO4Oe8D4/HMFq5k2J+rJ
CLSK9ImpEom4V3Y2ldDIaE7LQRPRiBnSsc2Lv4bEIuO7gLmrlkHUnZdcj+3daURO
RBc8G1FbXmA1Wwyxu0k4lau/tb+3kh95cyNh72wNO8TQF3j4EFjX1UP6HI7/JPmH
8O4GTlyzHOL18+PzlHAHik9VnvxraazrxLznyptcG+ct8EwiElyxqrE5S1krNdg0
8i/XAvGPJMrGf9KKmXQIq5TqwbjtiFxGRmtwvoZrr0sNUv+jQXVrr2CrsKP+nQQY
olFWZnxvD6BM5esCloXYc11VtVODOvdjs5FPYozNCT8xA6/KqH2zsi6GbnPEFDq/
sUCvebLOHocL6LUil0gSJjqxqeXN/VsB81Fd1saKDbuoS20osUXArabACL1Hb2E2
v9d2Tc0CObBSc5BMI/jzar8L4MoohuV/jkGpZNYlFFJ7grwTUYZIDZt7y0iCNeFf
vKdiP0y+h77D+OFknsc9WTsGu1Z4RDKGVflfkY0vIjwsJBIcAvB2rydyNRsK0++G
34KEwQS/RWY+6cOB9C6mXjf7FlJ0uEUyMt0vzbwYxPQNa3oRraQhzYV4sSiO9ul3
ueELSr/RZnrYlKYBbKcGb6Kc0JPcqkQnP8kBFfuAaC10zWRqWll9K44iDaAfCAbp
0FDO/XuYCwojmbB3bDufkiecJhRGru9s+MZBVVSRglbkDqbeIDsdVY/KLDtYH9Qu
ynqrsXEavdDymUa63x4l2cWnWFJ4AV7b0qUXMLOICYtMF+OzU+zUNl0Gh22QJHEW
qspT3lLSI5nVm+WZ3Dfic+RVlap/LQ5Od6LXeNS8fAN14/GO3/lsAgJWpB1ZgCQT
R+gH/oLk4xOpZg94B9Ar+BtWXT9OVEqQSL+TVgNFljCZcJWbrYCW+OCQOW6FpXpd
Ht+nYRZoZ1ZSk5Xv7lo6WKB+Ig02BWcb59Ltu/ZL2bIZQYjLEGKrPBK8YoLOPx1d
SVcjhnZQc550FyQqiYpwc7Y9J3BJ79D9WOnAOzEXpkXh0M5sHxLZIxeN4gzWAxuH
2qTgt+pAeu5bVgcs4wHqBQ8wGqmomCiXJO4BAMQAf2QTMgryALUXPoxS4OgVAPbq
QTV+STSbOHdt+dfS9axbT1s9rJBNHR6SvELdhzSZ8h0I94aSC+1btv2oQ9oteAYJ
F0PYBZRw+kWwCMUyS6FDqoR4fDBxw3vfCevD6iHMIbw761ASikU6g3sUBsJjJ77i
8WGo8AaP8AxnaWfugY3pCVY/XIXl/mWliUFXaiR1YgFFidFfa+XPBiHrUUUajjXj
JNX2obQ/uFd0ltPdATVY5b+CSx9ELqtU9I5C9Bl1njDUQgQdqviishKnCkhYPz6o
eMrwregBCL91qNwlJBHKxBx1Up2+xE9vx9b+iYbbZcz60QpqOr9o4LWM19i/+y3q
wZV+PaguncI+fAzwX47UXffTeL7JHzVNSCCpEzDaI0crD3U7mhnk7WGfnol2z5o+
e1Dr4S0l23Qbmx9w0m1VRdz0BVlCdOtQN2Zyv08hHgkGzFYYG0R8hZ/kpUtERY4e
ywuoeZJH217xI8Rqa+bgD4AQJgRu+jpFZOdWiWObuyFw3+5qk4W5pTTrpE7E7lff
FQO08WEvO6Uxm1Y5+FfhBYzWYkIausIyB3lguHYa8adu8CegBw6mrqOUG8edAmy9
U281XJTF4Ybp/Nnn0EUYTD/Yk9qpMpwPlDUmjQkWIshFn/cKWiNLRwQBMOsly65t
BvGQPJoDm1qr0reTe/ZYM77dZ8TJAprHElF2Jt3rJYFYa9fSmz7uSIM26hDiTad7
DNCldRwVlw4N2fgTFFu9wWMOsuyvGE3lkz0zwMcWd1M2u8lwmblE+aKOt92G6uwq
cthGmqgxoEgGL4veaTuRp/djaforhmazVo2+77yxW/gQ9bONd/to9IdSrXDaIiaZ
Y7iBb7wVBc1MRaW8q0T+hwgMoQLRYigx8upJQUp9ZyyiOAMEb6RnG+WF696XuMZD
Hs48gFLC+TV41Sqj8QoQIYjVcCsz2hN4YCEXaLTHOv/KkDa8Fl71OUOIAGEegvo/
fZcnBAS0rNGyq/ZprpvoD3L7Kpi6f02fi3pQjN/kbLREmOHx+exVaz0y/xZvn44/
JJvxyeLYYCB0nCm7MzLyQn5098ZQfU5pUDHBHHS7Zw1plI7gHT9W45JBgbzd4QJg
zDbpvRTqb75OVu7ME1QaWJJItmZ5EEOesChaf99viUz78O7D08ZUiv0c6Qvelx0q
t9QpJgywus3eb8EX63P5QyQZJ5UxbPjg+EiguTUEKWMRIvvH5y6IV3Suq0QadTX5
CsxtD6uj5RzfaxhycV6OGEdcpIq7sI8gT3SERm9L8v2EAUCEGJ8uSmxmZPNA3YhQ
X6ASGkpo+TLUByKlgOBNxUsAowpXrg7wHmco4tmBJg1s5uMfizt/L2kkDcjaouOo
I3xe86Oen9ayd2/lrVVxcTwxB0exSe82YeuJYl4pIv87CJUVypH/BJ7dT1ANRYyo
7k+q8FXlhp5vy0iimOeSvVYZPwUWfaoRDuRwN/paid5gujpQjgGvlUkPPTpQShXH
APjJLNAZiXa7PVZ3Z71Wl7LjVSCbQ+kq1N0ydvwxJDbubdoy2UXctf1KM1i6xLPY
H9u8lW3l2N1FJbdl0aFUfRtjV+2iP5zVBCMHeM/A3bCIH+RozBXmdtj7sIJt4foV
XJNR2g+5+STUGu2UY2SAlNQCprcsSff0My3hjfnfeN+Is1FQT5eZi6MW8SMmXWXY
BunU1xYHryT3tfOVM2X7sLkWdyXor63uvRsFqhijlbhE0HgImy0BNVo9wkg0cl5/
VXgiHVfYbT+ZStm3oBSVcK5dQNko8q9AzYdJErJSZ62PtcFkcBIB3AW2G9lzwYMV
XYdCBwSweplwjn+m7OKirROJ4waw2+tv9CkXUmevAiGDdrxRfIAmTe06tF6pOsFk
VFdXLtV/tp6dUMdcd7Bw9vqA6pJN3eBF8vbn1KriFDoJlAt1SR/QXse34dfImVCO
8JjzGfRWDsAPI8QFw6frtOlMgJAEoYd96BFIvGg51g/X6VO4n5dZ13OrbZfkUvrj
eTPaQITqiC+7QDN88k0ld94XxH9kdFvcDHM9cEOglsYv2sF/sLkfrJTwVXaj6EKv
OKi4iZ1JdIDVEJ4WSGOS7Zy97DRwj7hbgEG/La8/nfigoZJo4s/64ULyxosXr/QH
FaNn4LslCDLdoxCPe+rvOywJ+GtZIU8SQDmPdHza0ojDDjET5RgOkYk/po1PAhDO
rLPaIGtDU7msGjFVPbDzmSkj7F7slv9BeWc7lpX3vZq8ls9wsUdWqckWUaseb1oZ
hE4JDFzToLSuGgsZWDjD4fH4FbxCG28ykSJ63ZPk3gxTUA0Xyh6dVXFVnulk3V6O
TaWMyK/6Cc6L9RZ2sglZK7xrJfJlRyVhdDLRu7WsniGuyLHto4h56X89tBeR7qjN
RCOuqYiNlWVvcghD7ibub6ro0iUYGYhIOBF+P8Cw61T2pHbsg4oY6WgEoxww8ycv
tIHCJAB8k5eX9mySeB6BNhCXI6zh4Qt4rV89ZGM4iY8xlJJ8AGFhO/ywgtzcKTDK
CWvj3MSb1NaQzdiPLkC6vcgZLOXBqeGq0Z0Bwf9/IW1c0VTBKLW9rti1+V4TRxDO
AabBnaUbqRBoSGzUUVZhMUuDHcxqZAlYBylTSt+YDNAUTCRlFX5iQ8Fb6ZBP9tQ0
8ZsMx6U1hNhv5G0+V5JoxxHmEH+3eW2PqX4lWvJSDGwXugB0PPMeN58DUCchj8re
fH1xb5FzTeri1/o963+9coK25RLGmsEXeK8p7VWWvT2DLGv4fsoxWGN4FNYNO0VI
oHLfCJi4AVe3KnRlYBuYpt7IdtFDHyi+GRZJuBK70MFYQqcIiGHfABiLN7erGlN7
S45g+clPle/qEY3AE/q3B/ExtdCprWJzA6IzAG4w0MKen0GDLBZOYUp2n3QJlrTd
4ERr/pQFjMEGXiWY9PAzC8YZYPqVzfzMdD/qg9WO/n+QrtvquBL3+eHwVxNFXJXB
Y0paQXEmGr/RyGpf/PE9zDnN0gDoHgrJ04TsN+rKVOvUR6eCoNsThZ74fAUDy4oE
YIiyENm7ALR7yuw8sW6G2r0ylf7CNI+jQSjX8HOTEVwkSiOYYOrzZesvzsgCvSi6
hJMg47kviL43wv1HDa/Vx2yKWbJ9JGm0X/JgIvjVo50rIiTf7mgYIPiZL/w0BQYF
FtATRlGYQZLuyU9SJEthdA3mKsTmFPVMmBcE/HHGyD/PRknNxAQhHTUJCEEeQVJ+
uLw5J0HoKwz4ZTO/wAqoFYceXZIBptiW2nEkdRxjxr38OJowcVAmTQ1ejnXc/3lO
uMkHnOv9lgnlQbOxLn4QqQboBFSuQIvjOqN6Grk6yokSNvStm533FQ2i6IOnWQaE
REOI3N1H4t62n5soJuv8twPUv3ZDnAXzyYTw0w0O5nTmTSLyd8awGpzPuMkjI5I3
T3dJfxkO5gdgK4UKAUH4CZfma9ypfKZxnTn45gOAlzPzH0wmN21a+JqbM2hcVMK8
Or/YWLOoI+lRXJS1L+BPate2n3lmWU+BXf2aIQIDZHm/udUzwZR2lSaG96Q8/COB
52pfTsxK48h4Qf+Q75PXBAgyKqCvyvXIOQfdmb6FJPzOn3L99lGReibI2P3M0hdo
jqtom9EfcjRLgsHjn9wNzn0bH6dru/RMe4tva8bfk7zBDyMm5vGAu5WYfQYjdNAA
GFSPARpB3mABN3e4kQYte+zS3HAcRckj1rUK+HOGimxjs33XPG57P76M4PhKa3Zq
XjdMDlm3hRHUpjeIpaR0Dec3XftGkSnzYI6hX92Ryml3RE3QkQ5VxKz2WeEwc29n
LGAQvai4bqY/58ojCqDjNIj3MEXoInidqtljOs2U7Ynap1P5vIyn4jMZfYX3bDXX
2R5ODhtz72O+BMohrDyOoAeYFtJgHpVEkCRvOoQEDQxeZUhSHjRXCt4hflcg5qMD
9XkSDL9lLg0WJ+9zarinYQMhBmLFxfPExRvzUux9DVpDNJXS2ZPAJhjVrXA1v1lw
xDL6Z6jrnueBaHOMzmbPwPmZNjlAPilOM8Uf8uxrxiG9k5J6dJFZ5EDmD+GJRNbG
5GJDJ7apYvzkXECG567dx6yOVYYccZLbafJM09hSaQWoMG4VUeq2R7CK94dKsQWS
kd8r6BEDQuC6MLfoLyDN4TExoDgpjDv0IXnmperlbf5ncjtInpkH42iI5QX49x5Q
6KmKAzRA54Qp9kzZbSGusmBnCgEgAzPRFALhCMyIkjK+TQo/gkcTObhEnNhiOsoo
BctdHYtaV23X0I6nS7EShB6u76OCmtqxvcO8o8zIyA3d88pNRp2d1/VS//EHLfzr
5O3CkIXMCOZ7vER+yMD2kCnKgs1kL5SgeIz29WjITEkaOG/jGsK8tamw+dwUALYR
54PE2mmA+MD9qOBnUvH70r409xqe/rgftkzHCh1uvGvKuFQI39mSe+4tHDosAHSN
9eh3DrBKzaU3vm9EQ0rHggWzPsi2CQyuCnDulyhu0xtJX8WH2ZGXeL/Y0mpVX1Mo
4fSTzsOGtHensMv+Yel8p3oTknMnXyItRHNUWcSQeITH+Niga1A/16XPBUfLc7Nw
hUD6Q46hdZ3j9bnl3CR4bUdw5GVPH+DOGEf0kJnJyj+FgzD1rQwAzZ7RN7c4Ewqp
ZAkM61vx8C/WBmGTXJeO/912G5zmX3yjbpO9IzoW7rqGSjcfnv3Ser8eslumeJJQ
DzeyEj3LptaRq/QR14SqUO0vR1fxgN0HwJP69Nlr/6VjOFWgKKixJfgpWnryfH8L
eOF8BvAYWZLLiF+GZo+hot+vH3HwbwXodD8VnGG+a+JIxHPH8GiVgmNP7AGDoXtv
ybtrVCiCSAJmXiacH2AfGYC2MaDBZN6ya5HPCFcmT0lPHkYhcZcnNMzK1MCTa3bv
dQ5wLFl3amqBuolY3FwT4meTKCH0S74GpGSi/iIAez1VIVtZkOJouoo8nLU4YOgd
/KURplL1rbPma8uMZZFtsqN5U5DFMKZQIRcPXTAMFoYw7XUloLI7Sg/WIQVOueXi
IAwtzqjDWV6WCuRFwnHXBNMRl7GOQghU/2UqndJRR03rx3iPp5pt+bwTnG+pADGt
eQIdHcaerVulYf2CMl3YOdzLTopWusN6+9ulbP8Vu15tlj9Yf28DjZsGMfQ5ylZG
Q0GM6t63KXbDqMkqo1TwxoTGgSEZ6+YElsuR86XHHMjuYxhUDvCAaemHj4ALLd65
YtM9J+61kpyGrPUxGqe2vZqDHYl2PESOwfzWXIuUIiMvg6f37+XzXNm3aZw6fMcX
xbWx9pSQtMLEbD0JHSRdXshCJ6pDafJ5CyzDZasWsCh2oY4mcOcAh7wzgAEW5gmD
CEF3xBXGmUzCMQV1yWvgoq5ALOxlLjP4GAQC75JCETE519a2HPAQKu/Hppe1pYha
LNcTewMXbwBGIvyB8wp5xkb+K+CkWhFuik7015iMb6Mu+BfKa18ItK5UoprgmkWK
ru/U9/ogrkTyIAonXW6Uf7iEhbWPHrP5d+5srb2/xmxIaZX7Zvjo7INTqrMrLNeu
60BmDBNaPMxXKcHd/enh+UQ0zrr5wfdsQyE45NWkiy069IB5Jy6yftw243q1IZof
BGvOpO2+Tvvr59VOvKt4XWwv/KPtydFLmoI0w2bAbeyG5eCvfBMIbvDMrMqz4EAc
juDqjzPJyOet7EN9PIT48PvPiYPmdMp7sLWugj1Hs6ODxllLYzvgFsAqY+C5oqA6
doZfln3QynakzHitDrwm94aB0kUek9JjPY6zQX+9+HVpsubnk5XpK3LOaqXO/CGw
2Wrfoql0sL1LG4R+wGFd2lRP1LG4/vTlKTT0Xms4G4Psgnr7yFFJQFQNoxeBKVOj
/W4RgiQQk7KC6uVSDzcVsjb/RHY2US8Kfwl00ar1bJdW+LNGLfnT83w52tVmfJI7
g3k5BSvf29xbOx0yYFGTxJY45M8jqqxLoPok3amU9+2cpuvrlm9j6NL/QgiHLqAl
cwpMCdFhQfGWUJc4zbZbQWXnwbklwxWGiN/vANeEQCvACttr++aQ3uUBJTzzscA1
WWrtRxrJteo3roQeXe+8rZwBiGZTbEz9chrqYk3tZE37d+DrqAm4cNizc3oQ081r
YE9PBFcCpp7/fYj/E95+0pmCqwDfXhVRZ0NqT4XfrT/JCtOAaZhueLEKkoWKmsbT
RJsad9a8GMesiqHzMu5H1N/0UvRh60sAxHRMXJoQL/M2XD6Ox/aUIDGFef2KOJQc
bqgCqRB4rc8lq73E0sdA16YPmH0crb/4e3FolByONfVFxiJ7jIc1GLRkkR9cv5ZY
xwnUE/caCbGKXWeerJT5toUr97YRdBT+r25JfB6oc/sVSRVLyo6KNB6AJ/kJSiUZ
i48LPS8a8pFm8QzzBaiJQWFTTkN1zfH/LmAwA1uk7jydS6ABv4kMMynxCHy8DTgx
+A4ElTKhwZsj5ynqmd3QkGzM89dMx/cOD11EpA3vDdK+2Iu8yDf9fm8T4X8kQnvT
+rzAGSYt0iCpHz8Ar6cGMu9uZXuFCFFozNWAh3oSRTKZhLzonXLk4NH7YIUf3O8j
eCNKVtePVPdrr5wpayeuNFQdeiXZk7490Wp5wsRBacpsvUf8FGAV83COWRpLIsUs
e+NBPASuLut+dgrLgkvj+nawJ1RRoaoejxyHFzFrvvUV7q0NmeVguNdTpAGmK+hU
UL3fYtDsemO6oTlfLvA0rpQLeaEieZ+ASGOtDV7NzncmnmJDT9gf9fKxfmmi/uK2
O2M4Fvcw3iSq4reRLSR88MtiVLp19b/Sdg6Iyhb3HFyORd8B2CvlF9zh5owRfkZR
x0qKtMx5GtdvdUC1kFvjmP/NyB6iaSM5qUtwqtt4w90dvWrB5JfDBNMEFVeoMJ37
KMorVm/h8iGVS8FJrOKAug/8INBhAfufKUC+Ps7rMFHqqCmYkQVMJhuZQHyEsyzd
Had54sWkKn9oVYXTa3DNJwXab9QsfT9jnOlgui3aWyzlBrW0VSF97xtUxtxp5wHY
0KICqk+Jk8sKsZZNNkkVjQkitt95zPd+iW7D6SB5DyPp5hzzraQGJAttzczfo9vM
Gyb4Z4vlh3bGVSSdikzGOgQ38sQxM9IA2U6CPdrayTFPI4TvBuVQMgTCYvbBO+4z
R9pjG5Qjn3ss+lWgwSN45/x57bfhV/uL8M42SRUz+VYUosZCh/ZE+u79Pk8o+p4R
IxMW6HEx5K1v3s15LwNcE9vAHPShTZvfoyQ1xSseRrb3gWcBB9yoCygHaFYCJ2vn
SUuFcQ698Ra+AtJSWIriZZaZZ9RBsL37CKhIggymB5SwMfHhJdCZIl660VbzGDdh
ahSQMlVfa54CSHuADXHuupCXV3D/5cLe32Jgxb5oBloiWl7b2Wy+/NCvVDvCuq5y
CqTZFjH7Q9/pb6OqB4W77gALUrcocjgIoJVSaftlt9mUtSbendWXLwWjX6c9GFsg
WIsjPdFvsJoiiwE7WqAm935T61PTUh2O4U5VCRdiErBTx2oHD6ztK/rCcHhtEl4H
CbZDNuye5mDkjELf2odtBzVFQFbyTstBOPobHSHfCF3U659l0US+SrBUOw7gACqL
G6qsv4eIC8a6fMidmImOfLk4BFdc5FTJgSNLls7Dc1phVPL/y+zX8ZbLJdaGl0go
MkjZaYqThaY43QIx8z7cAZpB6zlaHBYYuxIAVYOCjcGlqihn7Ug9WV29+B6M+3PR
vCjFNGYmTa4mMMpngkgOtkEqu306Y1Eo5zx4GWEAhy/wdTA9X7N2A5yp0NmTfj/P
0j7pG/+0st9ER4jlcczxx+RpDGXgtBYqIKwBbBoUIchDjUSAXl6NGXgsF2BEIOe4
DW7eB9BfLNpky7Rbp3jRiMcty2jteeI6HKPAq6yWI3+wlwxSF3rfwa2zQhoKcjE0
WTLJhGsyURjK1ldDi21J7GiAlnBkS0MXGH4QGpjXUjSE6Ew4x/KlL44FwOst2aPh
ZJgdGDdl2AwE9p3o1kNGoWHdfqu6VJmYyK5GnCSXr7okghjhM0YU88YLkTFMcw9J
ssRiilieBlpP4Eh3Y68s4wLOSYGhawfeDz2Z87oz5YLemd8NjCLKEQCf5hsNF1LF
/kJ2s4ot0DGUg0vjQwoYjs6Ahs8VxhKlB/6fP0SoYuahSksQFZ2afoVgBYuIwDlS
BiH+deCtJSkJhUYGVlkTeX3msMADV+Koaw68HEx1IzOLFuwyrpjIgS+jXG4Oh6YA
zimK1h1yy8nF6dFfg8RviohBJHxFF+rO8//GOaEfIUD+Kpi/TY3CWdMHxO7R85Ne
vYSBY4/UAeVsSGk2xOpIIa8d6pfbd5dhmtPRXLgJldR5/iRqf9xQ3ewxf4rBBXbr
Hm6YFU5H8XswsskR07vNiqmbuCff87KwIp/6UJS2nIR0D6uKLR752WGzmZ7XNiQM
ACoqg/l7UCcaOxY23tU2p2wInZL+kpFNGAy3gkRvS9Q5scWcaQBUnKcAT1zH3gNg
SojoIrgol/se2deh5qxVhM+dZCSKNn2S0Oem76q70u/7vvTSBD4nPtlD854GvBU2
MXgJGcj2ZeDN0cj7A5rJUiNFQDFZ4HUjRa7lHl+fm0bjhl3QdwrO2KAcuEeodjnY
crl2pP42VE7C83tAsKGvIsA6SxCv9IoPxazQZYQo/TklOxZ5LQzfWXl8hO03VW7C
HHCCSqDpZGRASSZzCB+xBtKeb+FGFzhyOEQKFu9aJZ7mTltXRDz8eervFKT9I5Yn
rSc6zmN/OZxDTl47dnJxRs0oWB0jEwLYdGw+uhyOZ19nGOnZiw2mXZ3jRG9x/QXN
O4B0oUWAfcEuxrCEONIKD/9K5YI3TySB24ccYmJ9xETQ1EDZeQMAC0OMC/bNSJi1
kVQajGZQy1lkrUo5hUREJbZWQvspDjat8+nvjJyIfHZNUPyOxvBXAo7HhzAap4HN
j1cCxzlXuPvXxpMM1qg0xnlv1FD9lDKvS9yihFnuffTt08isXGa9KzGN65Ytpo7e
nXZXWB7tluj5vEKM6rRTd9Ny2Yx9k38rz+pxrDYh+Q+SE1LEFebGoh7rTpMKhRVj
6pkI6Lrtm4yGhjwvb6SSp1pn3wMmdlWjfhi4nCwlhm6DvsrmW/RwOOE/OB9B8Kpm
WYQGV5OuV1FMizFSbplteArzuuEoSC/16uxne0ef4G9O/cn3YijNU8pNxPcEYB0d
UTnAdLAaUxkRZISWjzRG0bYNSg5pKYd69Ur/S44H/eXQRg+4sNx7SsNuWb3a0ifc
1sLuLyUkBo0SJXPdT/+NfPP/pSqkeTr6KpwCCEGrQdu/LaObejAbLQ1/+uZ0Rn09
gRAlxMusuYY9r4vREy0dyyj85qzZug0Yr08HppieSzd4UapyXEFRROhpS8RDP//m
QxtQhbGMmQNhsxvOVv7e+s9WduRJF5c/B7mvZDd2M7+Jmv4fRS+gVnhw8emlTXDW
tOrZKd4ROxpOgUxzRl51mkkdWc+DRF1O3aW3VzIZ7MuRtcQizwlkne07haUEMp4O
EwLMYnU7UgC/kD4heP1Qxz0XWlBGsOYbUoFpkgJalNpV4RY4YsbciN1+lWzysyEU
UHW97jpNnPGb0okW/qMl0uv7f35fkD9s+kueKdlhGbfWDODkDE0NpYEsFWFLzuNI
vYhPfeeVF93tv+eoCRLaY75QC1Gp01NN6czxPJisHRCr6zrJYweoaQEq+tO4eyKt
OQ5gUph0ulzgXkKCofwdIA2TOubARUGbGW5sYIVHtA20stp50vEDjd7rAsXZLgF5
EL0MewnM35hodqYBZyvWIL+XF0oZIdsiy7sSeagdPA7as9DSBxboWOB3g/78gsh9
9Kt3NhI799j/wCT1c/9cz6dC9BkovHrHcPSvJJOfnT2a4Q/sIHbMYq+TK8tg4nY6
SbLDnBRRxaQ6vNoUOUhszsDpdWI4qCtfkUK2rDdAw1HdlDKkPxXSuRPLoBpfRrRP
lYp0Yu8z2x4LcEvJ5oBd92yXytZ9IN9LlROKQhP/nr+jWNlUTqbov+CCKRzzSF0a
qZHX/jQfVDSbIFDoSFMxuSPaGJRS94qDy6/uQFKzDVOLP4t7RsuW/ZWWJBX5iaeq
KZ5h9Df8YwEdblZNg7F7FogdVmZlg81KiSoEosNF6M/F68VIY2MSXAd4glnV+3/0
64/r8QmksMjNp84D+i93UtU2RanRv8OBtgqRoIEiokApXFSSXmO3qUBzO6dbT0N2
gT8uiwS+lJr08yIVZyAwyXQGKEPvoyhSZjngqi2ZO8pXlDxWM2zBrz8jlvUcKG+D
4DWTs8Cw0UJ5/jUc3/rS7SyUp+SaTIw5MyDmCuReqz7wacWEYgaZzN9lMh05310w
02xsbvbo+XIEDNech9+O3Skc2WwFmn8GpWCLQIqBXObCyXfJwqIjIZpXxLGNsi+x
tWGuDlXbm4f9BU1eDcBiaQ9eCrOYmq6RNkC7ZvI8nrgrrgf1QKzRnnt2gZZyxO7l
VtwqQrb1hYc92fPnMqvtEFKQ4TlewTrhnwcSVJUZhMadWyckAyOn47beEmU7LXlq
DDeEoaXuRqkGXcp3fDwvrktnufTxx1TzWPxMV8NFJEwd1iS9hXF/WNV2lQLSddqe
sysDiRvIP24m2rDRgoIJOsYhePlo7eNFSlOMJ+pHJV2yJBM9aBjy1l97KbeJLEFT
M6eFir8qxhVBQ2gNM465K2PEMakWldQD+auT6wHc8L5Zs9lnh5ypCFQEIjLhHZnu
6gQPrEuGjax6YdMJT95zDiXekVpYnDoCEkirlMM6Qk0n3XMt9CFw86+/DsOWD94D
BK9F/x1KYZZxRVlut4FMhHNblNkJbVlqicd3ho4TXBV7aYOLKBwGmSO7delaNclC
p4QKCkRqZEVXwe5U9UeJgZLU92NqwcouTcoU0GUM27FG+v0iNYbxZ2ubHlqojCJ3
rYYH1kx4Xlrzpc7263zrVOpGPyXQdcVqP1PI0RLC1xgKSVZv0x0kxgYZSTvOtB38
Bf6wQ90uQL53QBZ8eQ07YGAK2ZE+cgSRT72JaNqoSiufs87nJDPd+nirplzE1EDV
2mOwzQYjkvrvqh9CYsvkDhA9xz0Ly76AT4r7e/pmuVSOru8f7+BiuIi+i2XDDnB3
hEQTjKFi0pYMibcDcgWWvidFRz0QxM5JsC9pzn57qan12j/Rdz9wWu/N9q44OhxA
wqGsqOPgxNA+9EbJjypGmjDUArfEXWxiJwGFVEA+BCnIH+ErGyVwEtSxqKTVauU7
JB63h+7u+gFmguiw9IGfEis7oyBSZ4sjnZGOWbE8xqTltQQDWNTELG5ZJFONKDBr
kZfF264FW0b4hsk14NgldzEObrl3rn96CxikhM/hJgaCxiKhd3jY0pfJbRdy5cP2
H+Cw9BLpysTdXgJ2OLj5bF4Jak4XClW6oILI95V6acTSzxnHGM8Ym4G2sYnXLOfl
YIhj4Gh0zgo1nSWPGfnJKEnhmIdIgJ6B92l9cNtJ2o+kK7BrpVAueCIQTk1oIlYH
uywRUz2FxVBaAgDuu2BH2Hj00oBw4nvB91rb+hFfTIMY7VHeKXvMoFDt/tBoCr9z
OLwAr5YPAfB+5FMr04GxzpPfbZjqsXdZBAQ4tu42TMBwxmrdVo/xEpMGwaNUl3lj
eaOqnso5DJbvZO0FZ87o1qiABheB3CXCO5jaarEZWA98wG576mVi+GnTA/mrxoHE
juCNsT2fWcvWJrZAPh2laQlXMu09zkTbIqyPNtwr3+Lez6oxr96PWKmqZFNd5Tvt
yKuTmlpkOenhcUDSJPtDsHOSUTUUYjmw0jQd8tR7+l1Lvedy3IrhBVoIZ1mOwp/d
uHwW3T3Krs+vjb9aqSF5xxrxiWg7D3DT/8efJpQ0n9ggpOUGWCQ6pXCS81jcg0cf
c1VeO9gzMCb+csAAqpgsos/NCu8xb+vyqE8miKdw/mZhoyxDgmLkN6vWSSYcNVs4
ZF4SlqBgT6f5zPlNG7FTzLDCP3A4YY/edsVP/AC42B0+GH0yn8xgBoVmNKaon6oB
4FW9JTiIXJXckm7Ftqh3F0YekmYWx68ewVr6KG+JxgxZxXbxEamlF3dE5B7pl6O5
HOB3aMmUVFTQ0raDYLNVrAi/PUq9fxbITNxDr9Ci2CvLuIzQ+qTmzlPht8Bf+rlQ
ZYWA5AdyMEdnEWTCL+sYeLT59RKIRk+3yTot0bJtqi9thQmi6aZWL2jHLAA/Fpwq
pAlsq25z2oxfPqpim53Az7z0vy2mTVgKz39jMHSB3QbKaMSK+YaHtUkYh1Rhmf69
Zl0Zup4pOvYn/HnjUSaZ75LnTPcZnyXW7qPZj/WrXt01FyFXAeal5pjpIt1Au5kR
j64uGaWl7HZiO7sQNedlL9+G4GURzC3ettnSkOc8wNb44fx3gWlr/0180E7SDD7X
89efbVmIXeOI09RViXchLsuDr1WEz8dPFOczbktdKBYT7FRotbeusI5JqLegZ/2a
uFpJf/JtechkUc5+ULCUnSWfOidS9z8Q+LihSReOeBOtfS7NImYHr/mRAEVNCj2k
cun4TlUZKh7vt+46QofB/9PaVVSaLoUtHMwc8QEM7WZDqbIzQpeHkX/h96+wX2sB
jERFWYW1gmt679z1VkYHA0NxGNUczrAaRICjAgNNRWpCFyv+wFFZ3Hyaz8LTYMrQ
k8jbHO9LHC6JFXKNcp6rzLfTbZJSirxPbc0ZclHcVN6HKwFWAh+28+aymyZ5Urrh
qVev29UPc1Dln0gmZMkazJxc4JvCBDWCscSurJ8XePAH2IDIihZELxOlkc/Y8bIy
pJN7Ayo9BTPV63rbOpKe6Qu9+cmZVqTHC6CXKhcaono0kwl0soH8eiRu3m0dg45g
vHDNidVQnu9oUh97HvUc0sKlOhZDOI0DHPG+juwjTE+jjALsso58dCu4n+BuuFou
NqZa/uQh7/srMVVQ1TaKsCjh4Td2ncT6pxioewh7u7VY6aoA6KOZzpkvLXkyVAs0
etSrh9H2IU7GsQxc/tKM7vkj/Rh8Em5ADw+77Vmd64tKa8xx8rcbNsmx7mYxLH1y
cBQEcpKxGaw9Mzbk5r7+1RUrybQTQM1GJtCXoikp5Vd/jtOTkOj4kM1ULu76wMR1
dYz2u1tmdowNNjtWe0sjCtA0RJciLTkWbjPQPAKbRveAjRlFkKTjWkgEZHEM9ZAz
/ihUjSwvbQq5+WtYu8+DEyaAbL9Hr4KieJWZmfJTKw88+blLxk4zjHEsqgS6xZqp
uB05Vg7kvlSPhUre0qfqPSOdyKKKIWL8/Otq2B228UGLZMHEb+8d9gHDDQlIRFYh
LtrDc/StXoAZ7nTLMyWrnFUp/vkgAjX/78wEgVuJvBQhSCDcuT18J65XnvmjjUtH
k9KdSrI8+gEaUYY3wd3CYwKOgV4vB0vUK2xAA+BgL3kZ4XBExAOIRD2ajSSh6xht
aT9OSw4AVSTDJu8avGKCVQ3n3bQ2DkavtnUsLCPu3ilc2zMs346pkrhhmwKnr2+B
//NEEX2mxl1K1zo6mA5Bn1jP9F7ioGbpzfVlCzLmmzRBzDFzEzNRP6xruJPKWc5a
lPT8XTackRQKp1/8OQWWX0HSyF1BUn5x+CSQsWbk6ET8Ris33Jd106Q9JOBfgPbs
L3Pw+MmX5jJ9cmOG5Vwl2uRWM2VHyrE5kKtarsPHSgBwtu1GpGoy8Z20a+shsoCh
ESqc3f87lYN0QDqtgL/sisAgxR3FY8qsJWbnsa04AvlmHpWEO2/MVLezd7DSjISA
TPeogAITG5uuQa7Nzwrfmk4jrdW6+rGMTLs50TxnY1CHZxspdFdRxzS0MWO5jgX9
IJAS9c8LbO96ZP8pxTTnHOviUCxrYUkta5wA+fnOfQbhONOW2oPcpd45AE7STSnb
xGSO9L1tYFclQ7KgK1tHSmjO/tyPp5de34wulJSgg75ZdUjsXgsxDqxrj8Qm9Duu
5CbUYoKk/urapBHmG8pRTZHztLlNlFCfGQ+BBJcWvmhITjAm57qC92IejXrX6kLV
F2zPzo+leQqtWN6FBRNNAvUIEoUxDc9aFBR2WRT1LEj2H10SnTPn6IKz0AamuO8m
5Dne/0g5oIBS+9DOm+LCXG/QcOPbPUm3WdgJxkLqP3QbGP2YVkby9wIMYh9ZKaGS
HrXcVYB82vMzifMYDUk/Vhih0dlaQg9Lba6qpQjlwjIgEpY23XduU89NDFG0yxV8
7Nq0dzLTN1fAZXazKAbVR7e3fqIdFJZ7f2YQh98UHBbOP+d+fCGpnvENJRcL1L8c
ttUSYv0uagqUyjKqzDWxZfsQBglaUstl4vEufupjnSm0e0W1/1V9EmwyciEW5B/T
7ZxfPEHCRQjnSm758uLo6DHdbt9cRLTQUpL5Vg+eXqc3qQJTVbDGkR3DZcweD1Iv
qu1VGaniMIDVBQnZvAeOxIx3CXZeMJJ6MIDDATWn1xROf6QhXTKO/6XEXdRd+cra
iKm4fE1rz8Qb8acn7G1T3i6/rKej833wK7oH7PH4VpeLkqxco8C/V3FSPaibrFlw
s9QUiIOwRW2GUGte/s38SujUx5SDd2xe54Q3pf1sbV9Xo7i0bUWr6Y51MDcnJ34h
E1zw3xxpIK/4/gj9Td/pQ44yPmmo3NWwodJZrKPKLUai6u4ufgVJHerB7B0pIv9u
FeiA7JeqI5lERLAacURAM/vY+mzJFKF2qYooJQSbdz2B0lfSbsg/AW239QgPbgUM
TdjrXENJsxPWrrnlUOpWvpBhJX1F5I12QivLHzW29SaiHQ2VD3cxE25cl1wik/yS
Ecu83XG0VmaN1T/R2CA2YzezO9Qoc5AvxfC0nqrFS4+AAjRUAhUmrWXTPF+cBVQD
iesSJYNGmIOfIEJtI3Osv9ZVKuxzs0Hb0c+YCbC0H9BmjL2fE60q9zihl5d5dc1s
NSTiQ+ycehyfOuPziCOH9HTMkLbdi04bwAQQ43rtL1GDb0SQP4p4poorrSbCvqM+
w6WrjTrkGURHNrrEQAwI1lJvNKd0lICF5JGFcI6Cs4HaZuwKQkrF4gRwgaRqP4+V
whVYZ9LppvRWR/4N7CcCoQs4lshJRlLh2wemXyYdy3pbi9V97f+SWhfFiMdG/GBX
0qaGqFQSpKxLfBf3vQPQeGj3EQTqn4X0aYwj4gbYhYA1VfWKirVTtykGwTPXR9to
DKp5n4E6Ur08xQ+K1bDYx5tLC5FXUGINwSEZJFZOA35aZwzybP7oH+Hv362asImV
coc1LJzpq5/a37tbYlb9EeO+MpT6Qt9ZngQWX8Qz3XYJ4weOl6FoNl6W6WulwAIF
6qite9VagpwxOm4L9Stf97tVNa6x8QhHLIsNns3sjm983+UHG5dgs2FrqfGlp1hg
6byZN9rUOx2dGGvjlzTUYeZtBWyPJkVe/wAf0OJo25g+h9vjLNa8sdguFIT1GB8M
5oOhhtjbxYOY95A7ZMHiIKy4XYqaGek3yA2X04RrGmoDnBfPWKDzd+0dkPdLShmT
zz8lcOAK2dB4c42d8zQBm3HtSHM1vXXqVvoak0EmrWsnVYPBnpAHxcMINbEGrdLV
utGIpdRZMfmlwTRS4o0PwHihy6Osswxly07ov1FPP6WAMHy2QNZ8urVOUqa6l+Q2
M0e7WG0iLbKZ41qCg3SdgOEqskt4fmBp/tVOWNjsso83SsUbto3kUpdquM686yDD
9rEu+eEfQc63Bv8Q/sNcGo2Ts8hFA9oSrwTU06kjNWkL2coOglVQrK0txMsFpQFY
O2KBIsus3culvSE9Yeu2Xiv/5fDB9Fq/qBS7eElyzAnJTVk/OD9tvMZWJ5FDYsXA
9cNt+iaJ0zrSYswgSJiG/CqptZElK6EZw3pGoNlDy4emfnksfKF/uxnyT6Q54u9A
zaMUWVpFj6F+krbFs+6LH0sLKWTUmKfi72qwigpxPGpz8FTjx1O7XCqy9a7PXiUZ
6Xb/AnXwedNWpUfhvqvZTN1oCYVyJC7BveOlvSHsM54rm9/3jY+2pzLtyb6YIeyC
V943F6aZjgU/5M3//DimiCYRF+zF0iZlIXsXPaIFkuG3HUpMncb2dam8tcrA6f9L
CyEdTPf1DZSZv8yfkbAhVBd/vyYNoGs/MXbk8wqj29m12w5LyU1c7xynW/tio6A9
BL0EjW/mBI3pChRJVrgVWPlhBUsgv019gcFAXB4tBqNX+z+Vd0kqi2+AdVhtET6J
oJVrN0USTDH23AdAU3MDGBAZXNJMU8JdjQIE0PKykSDeQf4DfTd9NKCu7P6N34li
gBYRpswXMdIJCraIjT3wqI5jIksFL/kdCvUdmI3cDxenNw7WAy8UoamMgsGdkvSL
iK9tQKGwyOITB+CII/x7xyJmgPY1wy+6UjqPwjJML/PBsmsAvObNA/UVOSMyd9tw
6Ycs8Q3ieTDbtReHWDg85XZ95vdAKuwjCpLcX8QLu66Dnv9EWQfBbCbJqBsgL2pK
GR7Ap2FvAK7qdfMm+Dwo3Oo0CevVNbB/T8ZTvKKP51KSTriIJShxfMEstpsmNpS+
G+o2akIBo6trKXSLbIEcsu2dDiAlHe0ts8S0dFy2dPiLuIdLao4WpzxmEdvJ9YAq
rrnHYxljmvxeIjC5IOqI1BlZQHC/ihnCF420qYReAiXT8M/XWp5XHPBPRafH42Lp
24ugYBcb2QdCDXo27IPxMK8oVHTYiiNFkwaZy+/Mk/VUVWrA9WtsJMPakXG7ihlQ
o4ovKZiGgHhzqc9DBumn3kgNSV/3o0BIWMT5gZokNXUrsQiXEvT7CrH5TljFdsT0
WvoO7SjOhFeBc67vBcPC9CZiWbytBExHHs3sLmunMd/IJpA+Df3vysHwYiKfPLHP
nYtjvT+nMQpXAmHlZWOv1V6D+Q73j80GpzZNxkIGWnY0GzLldYHA835ezK/xe2tc
ih+Xv/t5SkJp+HENDYBXUX1HcmFI0E7M4MxKxc2+mboRnwiqu89kUDz8bidhei02
+/Tw5i5ESJLr0mOTDabw7ZsSFe0AnUgOHWC8+pikzlaXeLsY8sT4k3/XphRXp+eL
2bcRjN6qs0SIR52kZ5Og8RdljG26aD6BgWG7T6KQVYehnD8U1+1tR9aQvzg3CN5I
ioIZRCkjL3dir9actDbkXrxCao/TXV7qy6XuvTCBMOBajFacF62KYtR5micdkafu
2oE1qF9ARcxaN4gAQDRjq60eDSc8ceACE6g7KNbpNW3IOuvaYu3qwVEmmNmV2UOS
GPUaJ8JIx+WpdByKeUAp1QYzmqNYqbVPx/cls//vbCffEC1pnYpuYnkvxZUdLNA+
ngEySWJUWsZQaR1Lop4DVIw0nCGFfalzn7j3AACrFZnDIcI5hKXE3lIc0XdOWym0
gWjpmCSR2z6NzklAetLBxFCtMsAKhV33tY81XkbXK3a01u3FgQiRw3QBqDavagmF
kh8hl/EEt0vyxLyZZlTXBa7haooAFQ2wbE0oIEiYxqcXiPKNPtcvz+e/c4Eya1Lg
RH16WHRhnE2NeK7d0UqmPvCFdd42fIFW22weu6GTgs5nLSuGGIGrejCBav6nNcrn
r0DF11sLj0cLYFjce4V/D8nHUpFtUEe737O1hEH3XEWhll54rQFEZKgGU+J/jntr
5w2Ng7yFGgim3u8sfryURO8G5La+uBIA0VhdkdgRyjXkIGYJKaUVP3LadvAtIEQu
b17IDJaHRY+fz5Iw4yh8zHHo5/4ZLqpC5CKSMef298fkU9aHMUN00Z4m0OHJDN2C
nrf9wI1HNs7u5d91Tfz2dGENtWo5IHw9CImlbsSZPfdCPFn1+g6OaE4zFyvcdxzj
6EjD7MyCw4FWaiCumYWq2s3r/857OrgiAG8kA7KMAkiHp9CKTrMO1Rz1jaROekIM
/3yGIRgdPzuHZsCJF+zgpkn8qTuKT+6/7Rxcz4Qbc9fQojNuGt57V8PiSSS6Jy1y
ihCgjuixKt06UPihZSG9sV+M2VFjVQ+PT3VOSG0ybvyIrXI2OZDsskNaMj8wJkVX
1rAxwpuBH/jfOwigAAMxQ8jsSd5cJGpbPO8K8MCaH4Etcan/qLTTHT1OU+9N6nni
b/vwfrOcx9toKCNwiZ/ZTYj50pWciczZLLFJ3+PZ7KlTlfrRFuNgf6SyHRu5CoDX
O7Z1U7AZ2XFkAqAabpBxpmdCKzPizlha7b/0kUfJ5hZJbs1Rsb3MQ/jRXVUwBCKq
X5KGgbn/yxitWuvzwrb0Tos3ERWwth29pu9S2o22TxYJ9cDJAuaacERbNbglg/V4
NamiOStjRgV36M3ePmdmPy4uWmjOrT/WYWZcSSJlo1dYGP/+8DRnGdq2/xcKrxye
Cqpirj0a6B2tmPBDt+9mBNGIjJ68Li7kNsqMX4gWvnHIu8f4n1QKDlcmXB0yzsAZ
RMM58Ek2z11PtJhtYyYiJelITsbiSSPL6sY9qlKjs+jWLkGTEi3gaax6CRZhmnZm
XR/P60spC1iRLeg9Ue55Drz7XxcM8UkTMQ5jnp08jizIE6vVCV7IJo4vjqUWYjcQ
L2vJOzVR8AwxOrGl6YpsgXVM1hE8QHYqnIRzR11s9tEi78Sl1n2688CfQ6U6mVnQ
4VxBrUokydoeXbQeRHBPJYriBT+ONnjwxCzzOLoPz3rgH4bY8utmndMKEgYXH9L6
a57EvBH5wSW9RIFI1x0MOEzkFsuClYEBioFL515hN1WmsrAEQ+vBchRHUImGUBGw
VPOjwY30osB73ZihsQqKeaA+LOPSBQ1XK922NDh3iW3wbbM4v7MtvDjX4R5wLp08
JT5W44IJRCu7lcHCt3s16j/gEqqIiw8jik4DKnXsNUV1wmmzbjItoZeVh/WgaYL6
aVX+Ohz04SMs8+x0MgGfTNVRLvTXSd9ifaoHs22VEQaor7UOD57Qari9VPIdqqRL
zmuS4VuSSSCBVkzDowMjYZJCCvppq1+XN57QqlOLdF4Ji4UhJuzwr0vEMVtGu1TF
o8Zw3SI3zMPggkk179+/BVAb6eEji6WrBtlpfizBcMD6SKKpUYScMAnTVvLi46cO
819/HtQdnf9ZQOgCfrHlTPQwwD7nBjcedXfZFPD4A4HGxufZ9OjRGt8YQeVEwem+
UmNcjAf2nKTj38Z8pGwJpTmVyBcqcI9yrbuzH8bPDXOzvapQ6Hq51hLOd4VV46qa
mhZqf7vr4sPYtzM1C/X/3LHE6ZrOQ3EHNewzNj+IxENJSX6f7+xY4hQdvgsHEDrg
e34B2cFQSbb4Me/0Dk0VSCA6y5z8CZ8uS+BqB24JXAkIZxQrDpV+s2olyg7wBQOr
bAkrU/OBi/4vNN6uniAgNbOJ5TpzxQZ08ws/Y8XbQui3B3eZbHZ4QhRF9Iyj9CZZ
psuHpIVD3/zdh79pXy5H/qbe5C6HbgpGmaDCR95lgp0Q8FP4P0hGqtsQg3lbwJhg
X9WLngO3reRvPxEUU/Tb0Wpm/flv/tGDkOA2VzLfjo+1PuaMW6iSJVi8Sqq5Oiy2
OF0yZDOCuLfH7xeiKnOQzjGZ330GUNmMNxbffvcz3wSHogcFp3dRoMdagL2eFnPL
FnZxziiblCCCrSSBJC1IRLpKeAFoNHsGh/oHcyQHWn4VDUzjuwBq77/ODpUBvIij
10Vk7o/CmX9jJaUKBr2owfLjZ95ulU/CtPYDMexiQphDQQxgknL+g77Z0OlA4lKn
f9+HA1r1EhZ0AF3/L/PhVU//vqtXJ9Kq7NdH97Wc+aaJcj4B7SpZKO5F3TgIpmth
EnJeiGA3YKvxvU3eTeqCyDP7gfbXii17uSfTEsvTbJiFnrovmtdBtpG5tNzn6VBN
on4+1O3Mt4drLuxF24uKwfUy+4PVLpxvn/zf6IMdTrgu6/oST0sxL5EtOucJIVgE
rAhvbpqo0IdSm6hSQlk+2PI5BIzmPla5PCJVA4cBJMrx2SrB6aJ0z3O9chMSAkwW
jnZMz/qsb0EMPpUPpu7JAkpYxz0tO6LTzXX8X9bgPETfkbK4ygL1VlBhQdFPArO1
r1YasP1sFhNSuP2TvDBWrG9yKmDiHST7N8so64jaS/LUUxp+tss4t7mGFfj0jD+E
ZAyrIQRFX1DuresWYeF22BU+jNdyJQ3yhLX4Reits1NUi0QoktECGJKjuhZYYzjn
yS6ScN+YYKG5thSBPjJGOZ+bLmwPqeKbijIJzk5FatoF/J98p7+5f/0tItdtHPG0
OrJ0zadv1bgv+P9sE/jv8lOINLzQV3JXd8wKdExmfj6M1Qbkw9CIpQ2+24biX8U6
WFHGIfSSCcheVg8kx93PKEV0QeQx4nGW1pbZp9Kc5bIDcfIMvuvda3PKFZZLqMa9
oDd679F4noWiWqmoUScpY8FxT4nCpWhzt5HWydxqRzXZX0DWF6zEPqkLe1p/JDtA
Yer39wPCulEafxlkflsrK3P44fLzKwpTAlMBVJGBdJ5s9+TyeTF33Txetg1bKS0C
6Fk+jECf84V57IZYHHeuEf2aCXu7aDpgQ0DwbsocpfntmjISVdnlbfL/ZnseXJGF
jbjEhdx4y55n9r6AXB/XwmKw6QvuW5suQydG5kv0y0+5RyGRhHKM9BKqr4BF4MY/
zn53sfw7cdF1SNld5+AWm9Rxb5p3wYVOex6/OXY8rYUmGtDlXE6FfPiORV7CNCEm
5BFGOeU7zIltESK0iT2MQzxpR7CnYvOZgegmsh6Z7eV9OnDplbmxbtbpbBBQl+Lq
r7Bckk+4UOgRG1IeLxafrQ2FzSoqYtcgJ6RET3Y4e5TJNCMLhLne9mMCpMOTkfEY
H8QyvdOoIQGilbbt5J5+B0H6n3fVbgLlG0OziNZKWQwFHuJ1wdehClC0ZZuOZug/
GBQTYQ7H1y5591rw6koff6SinEsXvdaksXjK2jXH+HeUqiKDTqB4o/tdkTpglM/O
NJJHZpHxRGxpSb1TVpReNq46Uqq9gOEqnwtR+nXiW2Q0gNO5pcn/ZvtWajHsN3zG
wo3iFfqF6N7t/4CWnD/s0Ypz9eGV0rpRMb1Z6YzLy+LzuNBYp5Qnlq/lhBoUrhMK
CewNqx/N+V4fhSKUnST9pgmhJX8gdOG+BSH0V9pdWymLexPMuEPwmGJgoKB1ycEs
JrQ4Z+p7L8A5Fq11GVSFg9Gt4HoI/YIMQhtN6Wden65E6RId2Oq9Ib9tBm/5wglv
0iA67Hpy4AIis2oYZGEUwR9opLGA6Vu+DJPRum9YAd2YEDnGHuwnQzUcykl+IhT3
QdEBu0VZJHb55sE2PoZKE54Fml78H7ihziQqA5SVjQnayg7SJXp2F1igHiocPr9X
oeX3kl5kOIjmKc78da7w8iFumkD0pu58ZvrALXnCjbXi033gLcelzonY8hs7zwpQ
5uvXcWa1aRUn9JP+im3IZEhaxwDz/WpIxp61bgyt3UnOqE5UMIXG/YFMwc3sQmKN
mGk5QttPAcGJh2FihUdFw4K8545vhHmKUN35+bwhhX8c3EnmVrI+CqSyBLZ1zDyK
gDyJlzmMox39GXg/sdrHgb2o258m7tv2wsbmf43PD2zVMuUTWuKC71I/elsrFLIN
KJ4ed5oaseZADucgA3a+bH3Q6s3MLn0mDWlTkTcos6IuivbP4caKSA9Dpq+BthM/
h3m12eplQY5dG5uONj9Il8mKZT4cTC5UxsIQIXOjKk42MXPd+JfsCvTI5T79X5vZ
2WXo5RqJe7jCsPlqStFDF+O0KyYVd2q6wMkKaQUrvuPMS2tGbN0wDQeWwBwMo4Ao
y77QAXYlEGYGc6FTrfrDN/ewPw7YG0iAJUpjCw9DuAwLP11mJqVOHshsN1Bt4xug
h4PXcy+tmHG4qV2oIQMtR9E/nrjXGfGugwWu6RQHyNouvVCpAcPzviSQPKp8ISM1
I/ZrFg2fB+TyeK1zr+hsHKIHMc5n6VFZlRJN4hp/miWeB6vbNhIisjJaQFXMMCM5
n0fBW8Yjd6RERBPM6SZcqNgXcHe/ME9XXUv5Cb4cuaFlRmTf8D6GFsEFz2VkFhjI
lSKItHDTqkm48swvg2Eh5Bk9hTRr4zrrEZ9w+Z+1C+telH5UfptqNBA4aBsI9n6w
BQfK5OmV4e7BGVczFFfnN7zwwOCir+YunwtZbvlQ1chzGsiFZFVIujMoAOzo3mvG
RXEFqxNREDBjic8Rja3f2BsQWjyv2Qy7I48w1ufRs4sWf7Eouz61Nu0DasArVQRD
5xw8TKTmxPYh4SsCPtVl7KaaU/qEF42VlREf6VWuMe1lH5C2IPMzq4TwLWe0Oobb
rzl79a9f/CyRAOehohLmyk1DtO40aIvxEpezj6/qh8IRhCbo3769Bnz27C6Tyvgs
LHgILK1GbhxgojAVl1IMHdEIVUIMehNr6m09cUq2H0H88By60PsQJgQr803RPEpm
2uoZ7HiP8oby62saIuttDveMG2HvD5OwRW052Gb4WDRK0EdBuDU3TYcfbOjATJcc
gOmfzDl/K4yVFyotKP42tjEBp+NT5LB1ozocFpnv1dCIOJlNuESgOrLcLzput86k
I98uT95WdE/imrL8wIBUI6J6U9NhhmzJ58HezKU3hl0Z6vQlX6aMY5QseZBQoyLe
WUS7bRcYQAGCiVoReam99j7wDF2WSpvDX5mW1QqYrvsjh4/D6HJA1T2z4CvrQPO8
`pragma protect end_protected
