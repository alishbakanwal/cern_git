-- rx_frameclk_pll.vhd

-- Generated using ACDS version 16.0 211

library IEEE;
library rx_frameclk_pll_altera_iopll_160;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity rx_frameclk_pll is
	port (
		cntsel           : in  std_logic_vector(4 downto 0) := (others => '0'); --           cntsel.cntsel
		locked           : out std_logic;                                       --           locked.export
		num_phase_shifts : in  std_logic_vector(2 downto 0) := (others => '0'); -- num_phase_shifts.num_phase_shifts
		outclk_0         : out std_logic;                                       --          outclk0.clk
		phase_done       : out std_logic;                                       --       phase_done.phase_done
		phase_en         : in  std_logic                    := '0';             --         phase_en.phase_en
		refclk           : in  std_logic                    := '0';             --           refclk.clk
		rst              : in  std_logic                    := '0';             --            reset.reset
		scanclk          : in  std_logic                    := '0';             --          scanclk.scanclk
		updn             : in  std_logic                    := '0'              --             updn.updn
	);
end entity rx_frameclk_pll;

architecture rtl of rx_frameclk_pll is
	component rx_frameclk_pll_altera_iopll_160_zwfcdta is
		port (
			rst              : in  std_logic                    := 'X';             -- reset
			refclk           : in  std_logic                    := 'X';             -- clk
			locked           : out std_logic;                                       -- export
			scanclk          : in  std_logic                    := 'X';             -- scanclk
			phase_en         : in  std_logic                    := 'X';             -- phase_en
			updn             : in  std_logic                    := 'X';             -- updn
			cntsel           : in  std_logic_vector(4 downto 0) := (others => 'X'); -- cntsel
			phase_done       : out std_logic;                                       -- phase_done
			num_phase_shifts : in  std_logic_vector(2 downto 0) := (others => 'X'); -- num_phase_shifts
			outclk_0         : out std_logic                                        -- clk
		);
	end component rx_frameclk_pll_altera_iopll_160_zwfcdta;

	for iopll_0 : rx_frameclk_pll_altera_iopll_160_zwfcdta
		use entity rx_frameclk_pll_altera_iopll_160.rx_frameclk_pll_altera_iopll_160_zwfcdta;
begin

	iopll_0 : component rx_frameclk_pll_altera_iopll_160_zwfcdta
		port map (
			rst              => rst,              --            reset.reset
			refclk           => refclk,           --           refclk.clk
			locked           => locked,           --           locked.export
			scanclk          => scanclk,          --          scanclk.scanclk
			phase_en         => phase_en,         --         phase_en.phase_en
			updn             => updn,             --             updn.updn
			cntsel           => cntsel,           --           cntsel.cntsel
			phase_done       => phase_done,       --       phase_done.phase_done
			num_phase_shifts => num_phase_shifts, -- num_phase_shifts.num_phase_shifts
			outclk_0         => outclk_0          --          outclk0.clk
		);

end architecture rtl; -- of rx_frameclk_pll
