// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:02:18 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
qcaIjLZ97SAZGmyGmrTJFGornaDu3j16xFQe9SGaxyT2QjX7CIABO3YjXc+T0lS/
bGyXxPAXVajI4PeErUnqM4sGxE7GKLhNQoe8tLQgbpd4RlTrPqc5+4R3WKACClRi
Da8h1zxVYgjGEjoN/HgBusymzfzKWQqwnW7+vtckCm0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5920)
ceFlDS/C+H5NvZdhLMyoXCn9itPqf/zg047gDM0z/+ZUL19Dda+jzYEJ3cel7j9Q
PzKWTyKV/BbZ9St1+VcCp9ZZOXoJPZybetJtYHiX/23F+fmbeuQbvxAR/2ha3wAa
DaK/nDiwgu9sNNTfyjKTZwd6BJaIC3kPeVdiwLWPd2CD8y8VKW2ItDkchXxYvDUm
sDSYAek8Rx7iHPRIhLFVsdUoSvZCa5RdVsBz6G6kNgxkSwP3rlCBY8q4+pedGojk
Tum25NP409XPR/BfIjEoP1K5h6RAMKjrtM4f4324uwgRjuojLuLNjyZRAO2PmDU1
3ms+tDCTxQImzJK5mz6U9M0ci2E/nXfHWxPdH0XgXKOZ2gXcxrvWyq39PGntIp6s
F1JZBxzGLrGgthqBwDWhDr+2JVVWVOfahccE9jeI28SMdNpgPflM4039mwa0L3Jx
QO1pfRaRZ8H3VQqvHiNacYJMiymqhFmXLmFdyOnEBPveOWlxeNAr4oRAc0MBtw3C
mLU3zCdxIakcgtXRPW4hD65beCTTjZSST2w3WhvEVfhNNCdWEJ6urtvDLjNWk1kM
LNDhRHvoX6GosVSwiK9y1hvD136Jq4ilXemAvWaYlvikvdTp/MpBCGvk9HWf247u
92FMyPB+IYPm3TLoj+xADqthuGJOqx0nH93aQ7FzZVPPyc187wMNhbMtr4xeSV6o
u684ma+r8GnmB91BfW6Y2u/sxomicaGPU8QvF0GvtbmZnyolNDjeyrBsNRUzjlnS
BaTstfWzgXRctcFTGHq4AYuBHliFKabMBYGIxbguEPAlwGZvXO6zsy6JisvsWmsV
JL7tlcVrW0IDqWeQRbw8v8KOF8rwaR5OfK6p7kKxssyV2dM+TvTG8Jav63m1tHy8
JP7ojLY/4wudOqSZkkZz9qo5TLHoMJfBiy9g8wytHj179bsOqX5jm1kwNuz7/cvv
niN9+m4vhTK5x9LMbmS+NXEW/SVuHGNGY1/GygNvTrtCC4nVsvYDOgDI0IdqAg/x
rIpL0v2NWm87mzrL5OpIVTK6HNTO7oidQsTRV1LSLrOlSkM9Re3MCuj5G+F7l66o
uIbke8SHx9E19ghDqU8lSLl5gDTG2wL0QxJcgw0VUlsg1JLhjUjVNKq0TYJg/moo
VY3SEbfW/nqrulHj5PDoeaRe1Ta0X6toQ/EWjIqK+iR0njLR9xUDW5Rni9q5U2ZM
hrm1qvYWrNE8/Z8eVo91YazbC71Nt89au0ElH6Rs+0CZ8JsJpyDxOU5yuXnGJzTs
/TeWxbEa9WXpBjAqh44uN0PszpcxfnEjlh2+pfEKUZPjHRa93a9aKVPaeVfEP+jt
sl1vmPhDpmSt3Ma1UKauzF15rvX8389f9piJ+jBrXXnfoVbqeYJz8F6IlzkWmABn
PGW0gRlmZRL6gaTRcXkyIYiU5J11gR6Zq9xGKP1uYHmLl+5Q7cKd0OJ4ySXWtn2r
3IWgwqrYpBVbK0XsYC8eaKKZns0b8/Iyp7Nj8A49csGS9NLZzey46JbJFznVyMyn
/Vt7V2ScaInaUPAM6BO/5oaK+9Rk8Ki/gTMJTrsaiVRGrlpxUwPNwxcYTHvi5cWv
Jor3yJB3a5Q4G1c2Unq2MGbb531m2cHPAs9O1Ol6LXsh2T2SDr2g9U9shFhUvDZG
8t9ol+6zrd6x2L3ylSMDKKYVgx9a9IlkXiRL2R1vke8qqQjasadEnDEabV2NazUy
omeRNjbM9du3gQkRSS/k3LOIqGfj9CKrn6AjziiXos1iZyyUn1YGmG/NPSv+vFtx
vbAEdw1ESt3OS9BKTnQ26dj1quWaopdrq5D/a+qGH6OaqDHXevKKE+G0IkUyNXKZ
QicXUr/CoaI3wK8ZBf4pfW3OpFDjUrncUwBaNTHixoDJL+f6xqBEs/M/1r5zVcfL
Uvd0yLSEfP2jD5/Z5eHkijUkU/GRwNH/RQe6sDWvHs4PJXAWXGXfczPixqgYmPKz
OWdBuGUSCS4naLUj4E4rmpCwPtHM4QM03CJp3536vcYwsv4yZv/5+O+2/ijxKHNm
RbKt3/6QKflVg0XA0j66gmytcsbGuSJhgjexFy8ZZBGPSJcCTyPIz24q1OMp19HT
s0BY4lnSbNsuivveTMBeSZBAtXt0QcbEfxj3Pq6ptWuNrYWPehVquSK93O9jqGWF
OUMgeJDrrb/lwmIiLYSpU01GabjLfqcAdKiTFIpHUiBab7s+cD9EXEfUE9FauH/+
0AB9P4mAMrbBzus1RPIZVTtnB7lX8p0pvGPWqYs+0IOXKw+7I0XhxfUq2dRS0rD0
Rcha4nNEyeVe3YBniqVKLeJ97ov90vgXltC2kfJz8xswYD70Wg6TkYnR3JHuZrNk
zP5MQPTgiKkGF6fOnWPjbt8tR4fRv5hBDtJOxe6njVQrsSprf303p4KGJz0sssUM
9SJaGe3yCGXNBVgvbpw9zjMR7XBacL/W7A5hksLiDSbg2v2mnjiDowAy1AMyz2J+
S7+8dd0RBo/gwuXGuHQFC6KMVZW5q6LkMGNjrO64dXLggX7C0UT08cc1DeRqAeRZ
wjcB3v6+7u+RhtrZaiUvVaZJWOiRxBCIpO2g3eLfAaNITLhgkwgFOaXMlXd0I7gh
j3LR1MmHQy7zKsGHLJxEAqOjFEwawuHMxBgTmFTbsue3vqD/B9zX3cPtXWPraNJ0
9BEEItP52Rjz0EfWilYq+tJTld+u+Jhscu+cD0ZOdEq8AyjWa8EjK/GZhS3xDzn5
kfv3MbfNkVuOuQ3TqLgzMFjYpiLPESk8mcpJXTtsdFKdK4w0OXXmN6yq+eF6LB+F
TmMxrsTGbi0MTMh0Ssw5kPU9e6srmJ3bsRkFxpDXUY/cbwJFQrY7LxOFjQZ5//vH
owxe+gcpLgAFGMQyqESMAT8br3IM8Rs4sxI6n8tZiYnuhUahfn74YqUCTRnwgeWk
JTN0PWEXj2a8FmiOX0b/FIVBK4602UqpBOXr8zUE9nvq9F3fTdLEm1V6sTI+Phts
Nr5zJPvW90qvQ7ujSzBQDtQmr76N3urMDJK8Am4fk6SR0Xce3maf2Mu8v1UJaVMC
p6+f0diZZa5Efra19nxl5KJz8SQx/0W7OVwcMSJ3T/oS6EJ3ESpiB/pXLZzwAlZ9
rmKgRGcG+DiE9Zs/Cq1GZjirMNqp0NBcvTzKtIWZaR4rphZbdRErlOa7NpGE90Py
oSuDtYZG9fWOJXMfMWoB5QHtA8JgsuOeCQK7pFxgMWr8T/EISjQ50narP6+CPzTr
0V37i9auApEgVhtG/uyAcGdH5Yl81Ovk3qBb/CiQ8VCp1N+q6k5kuvIpQOPBWbxT
IOvADd6L/G9bseNXgAenx2hxFTlP5HphoNWwynzvXGA1SvdPz9uyxOa1cXXeCGno
fQgrwBzkCb3JhLbV854N6HEm7t2vL7BH1glNX2Evds/KB8jepfFVJK9GVEEOi6ns
sml2yqd9C0Yqb+sMDWg1CetfetvqXdinE2MutwOYzz/scXNAG+KAOAZpBLsZDsE/
zWPz2wOj5NYrdrKsGdSbJqf5vtj2Zm7skVPnfcdCl3jYkFtO/2ahnRfsInEnC7P6
GZnJxTsu2EN8UdnzDQKAoGFAI99MmHCuAoDhShp5zo2V67+jaLrgBAbvx+9pY4rt
h/ZT0jTqc6YSJdhgn5gxyHOilMP/YzJAV09Pc06kzlRSHqpFtveQKfG+c9N3Pavf
2sfnXfx8a5LZsOHnbVYXLLl2KG6mBPC6F8XGnsdSG+XHg0PiGNYfj6vwJgHxpO3t
/Z89jId/pOazPq9ObLYrJF4AzstfxkXvGmo3qigyW+c/Bw7IEXsqa2au1gjtn0yz
16kRUHqYksTQOpBmZR3oAYuJQglv2sLSxaw678uGicHMQXaEZc3UfZSfUem9aPe8
5MK2TLa9u67BDyy/c9ZHJAEWKaRxzgOuySE7y1wyaVLBcj5981wWUS79ABCj+A45
qQdUN7zt0jzJgHtQo54jDjIw0riLGgmkyOuzLnGPP8d0QVMaWzedROThLLyWUUM4
ApSzM04K8Q5cVAiTna/jV7OZsQ4RwaK+nPUHY+uiTko8oC+AIp3kaNukWVtJt+0S
8J/KQLIYIdXu5V9dcREQ++Se7QVjjHS6wfre06/1XVCEKVybYxj4gjyqjklQSw6Y
qAuj9mVOP8w8U3aW023x6wvy5FOArJRfDtjQASAAQxC02SUXAvAC0Wlgd+tF5HOk
IIQeYgCIx0HnWcR+Ub/FrUAkh22Vf9t5ouwIm0Kh9AgVR7h5hshKgjbIcXPEhcs0
qEa10zeTJ0FZQ6znDwGPTYywmZnGsdm37sFiMaBGvzpb2tJEQvxX+qkWOdf5Q7yY
XnyXCbv7SV8N1toD0c+VZlpfm1M8jEl0syZ897qSOSkS0miSTsfcmIvNNaenM5Fw
Xw93vFFAet7hWuz667Nom4e/yyA+kNRFfeev9Cp7PjALjHb+cHX/AjGC2r8/V3i7
vTquV9OqC/RODG2NV3va1h6FLt0JZ7l7Wqst5OYLDItZWUrR7elY3HY31WFtQQAH
Mq8KSy/cf51k3gpKgBK25Ggpco1l9fEcc1sw1QOua1YBtvWWdZd3/NMBbf7cc4St
VBH6hAmo38dFgXN9l2vw8dhrHp0Xx4FNGYm/sfrWjimaAZlA7pzzINPfv9Uh2zfe
dXINVTlZOtm7ef7RsEnW4LaFBotluJd6Ct7nCJ0cS74BLYVC8wCmd2yeUtrZl+4F
M7sCCfeh4tl6/yvtjP7cUp5w2pmHFbQacd3Jko8lt/BMQsAqWMTCK5yCuiTL70sp
gWQ8KDjkPA8V+e+NoJ84SD85qaw+BgkAvbZpJtFnBOcx7EprhkMS77OEJcBapqGV
0yaMu4fXPSY3k9BXGioxPt4O8mrm9qt1qCuCqnXaUaVK9aXusMu7x2uq/7zTIudJ
rZ/JttTbIQe7z2uPar4i8UDurPwyJ2HYx8TwT1kWJmYRpxIuYr3d9kJB3nHvCyWv
fxodznpePQROR0/IQ15mop3rfQ7KSTIepuqKUAlwNEoUQhEfJvbcBcRcSlDABzkg
pBhmDQMkyPncroVqwQeoDzd8Uj1+tHSW3y9LZ3s5qDMwMKaIOnulWaVb8OEV33Iz
4sVUVRDQiBxzZF1Gak7ITd7fIgq7fExtAL9H9yuC0knD9T0dGjBYz4y4ATzdAM3s
7kkl7hV3AqwBo6WoHLo3A0kuzhV8UdiSU3SojXvHNuKvFbVp1HqwPw1u7Toj2r6F
bSiggVAu5bPsRYWs9csgj/YhKmuuANMTQ4gpGUIrPldO1nHYb/5haIiR4vuYUK6t
KlP8GABfmVsTCtXPAE/MI3sVDFFrJ1RuIrganJIUsFrRE04DzXSIQ8m7dCzQNIx5
gA+mCkoQQlEnQhygv4It5DO7vVQl5658J2T5gT71bs4zZJehZYNai0uif+DyyT7m
qdYtmexA8+u3m+snf6MC9ADCO2N5HbK7IHvuETn0r2SXffaNfg3h9qWJgBVSelZp
5NBzDNPG64h4/F2+q3zPkP24V2+5d6MBlOhW2Zahno3GTh0IGUybEXpYdnkByNWi
xial+YF5t9rpj0fiSzTDlndGofWtSVebgjO3jB7xsmcQ0/ad+I8b3x2dcsvl8Uim
tYqGJRJjhhIlN6ZDU/SGlIlTgxBXEFtBuL4T315DHhwuXH/aH7twlsrbtgIOCeRw
fQiNKp/mUgmNP2RN9Y3RgfqXxBQRTITZtt+GNVjre8E6mQpYGOMbQHEx6RwgWIK/
vx5dlvOtqmy8at7rPUfSGcJ6FclV1csa10ty2Mt+vkf7ZQsuX78zsr92JTlrRqjx
JtidsPY1KBaN2aA8TRv8LMBddheF8gd3zk3q2CFUsBNeEJ3mp3/lT5RzAEnf4mIT
c+tF4thLevAO99H2Y3xocfuBCVRY3MbfzIHWNtnGp7iV4Iztj/9U6u2XwJFYoiKs
YegFZrRKm93i3E/cGtzo2I7p4aFHLwqdD+1J0xl1QBFFhwDlNwabu5TpczMBVZ5H
8vzZZleWF7q9J1PiNmLMdtW4/lkjjDufdvl4BLnm0xfP45KkUCag/+/AqBGVrev1
cSNg5RXyqcZt2p20q4VIhwguMm0g8RA3dkHF5FujorqPkj/MBNgq2jfLjpglFynW
UrI00LaNrhtEQ6GNuAkOHrmVQhY52EPwpqsserV6yw4e1wQR0OSZ7x4O2+/j9QbC
FTAyLaPFdwRag1L4IqEpGxPNiBa1dQBAREbKppOEDVelHGCPROWeT27P7t2J08li
kbKw5u52s52ZG7S0CAASCYpfuE5ApfRkCdERe0AyYBolzB76mEyKIe4Ov81azMWn
r5R1U5wg2agOALn+ZHIBQGAn+t0pOZAUno2svkewSuFb6Oo//4XE28ZkeVNVbWY8
Gi9KyIjh0Okbwe2ZlxeBoZ8Oiy9XE9xQBIevQ1tJvaoJ439mTWkWYnJlUcI4Oiud
x/x3HI0xG4J8KHFjkK4TI0jc+ySq8W+hx/O3jScC+s9srBdGzOsmla58dIpxxsL2
FbKtUXAxVoGtITXTfv0YITXW5GxMTX5NlD9DEgBkzwGU3PRFj6+FPyDXFpQtNZ+m
aAP2lb7jnP+F062Pirhr9/C7zu+ne8Z3/LuTGtnUKfoKFxH2qioDGTMBNewWBRyi
qCSF/uq6/c9RdDN7hGaLnkGd/P5kOtNNLOEp1cJyanTBwj0JcZVXl3fIM0CPs16h
38pEGku7pVGl3Cjs2IX8W0nZa2pAk7snHYtmT5mc0G8KFm6epKPKE0bKqG4s54ME
AS1EF6TtpzhSOJEh5g3TonCPi4dp7MjBjNqCrgij+t2cAT38N4n8U3m7GIz2hO9q
HorgqrhGHgOt3EwMVEn8ER86d/XrqDg1Z8meOpKrglIN27fo8K07RuhWGR/gNyFX
t4MjuFz8nIiSsY7zUeA6StpXvVzRbyGR1e8m2dID+xcOnzqVbEoUoTn3jPwB/rTp
gfG9BjIk7huXdeBLrFD5O+zlCCsQOzKdm5maP+QFNc+dIdzJCxWJ978gc5+fFken
+GJqqN9Q2bme1/OFHiy3DirUk8wDgFrNOvxN/os4yasvDpLUyTVZwA9vTY/udTup
bGBYFERbQbS64dwXA2OeCYt0UaJn2lMpnq2g7jQyzrlbPdL56QYizwnJbR4lDdVA
8dA/ApsfwW6w8JZH9v8TBiAY7ZK/tSRk5b8Gp0XuGoApIatcetNRj9vyrogDVe3B
2r9nA/MeTNUgTESdul/Gl9dDyO8DQuK9C5mHTJiu1GO/0UDNce9nkp81MTypRx3z
NEXsWuwaCYANUJDLwdhIllsJSyDyvHIZfVLR/HG0igYrxZVDHM99egx9UUpZQNma
3t2qkWtjb0XW6IUEC3Yy4kK4XxtutMmf7KBncxOrwmjjqzER7DOcab5CH/Oq+krV
wkwyVk08/MNwkkgfsv5pIyAJYxKQUC5wLSWWFO0W5yHOTVZzcBtcdPBnWQjDiMB0
BNRFigLzvDYZ/mLE5YXmvHlAUDIn9AukBvCxUFKAzT804nJ44NJjy9JjNLial9Bg
CA5gx1Les2z25hkZCdgva/wf9b/7UNP/S2ZYmaWEcrm7PkycLHeqU1lcjxXj7e0G
1yeWeSoOmisLYJolSzZrpJy7ukSYhhXN/okIMujGQlQP0Ruk/cYVOk21WH3XHMrY
Nfp0t8AAIhaJj4WtYzsc5kvDVhrOoVQb6TscwFC+8MuB4b59lv0t/RPKa3kWZFc3
2/Z1P4OTknuSiWJ4EBiJM/oR0uk/UFyUkStJ/JYQFf2PXbaOAvPqjZaCJvQ+Zv8b
rGGjTsgp12jRF+B72Gi1WJJcDW9EFElib2CoRQg5nEV8qmlElmvZfZm/7Qeo7Ut7
320WldfyuuNLciJn0SuGAA==
`pragma protect end_protected
