// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:02:08 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
O72+96iSGHDm7cCONgZVZ4+URNwlkuHR2CxN3t/zvXsoTJvDA+5Zq9UMQ9e3h1yD
4E3JfhWlXaCcZPfNaNoWxELZ2qwL1Fkmy92O7EsU9dBAvukrCRkh71pW0VetiaHy
8KsD4fJMF/BFVi83fc0GP/5WEss5j5969Vxgbwpy0mY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 176784)
U304F0smbkrC40LBk94aHw78tHGKyhdXmy5cdwxwysNkzRzwV2TVpHh91I7hsWm0
B+NQaDeykJk7eoHPcRBjtfZUn0TE4/ceHQwQzVpCjuNhyu0ttSsv4IU69zaXF2Sl
Bxe3Si9ph74qesgX8+IFeUhoHK+AMmK2A3qH49hT8ud0XZJD4I32Q0I6SpYG8uRY
rOKt/Kobs9mE01fuuB4GLG/6n1TD6SGf2R3EGuKU70PnPT0mu7wbrh7s+IIOcJEi
E+1WJcHYqhwGVhgAsVAbZPFI251DMpNVDGOy7qU4phg36uMr0ZplYrOMU8tP6w6x
J2sbaB33M3WV5jiSqP6ZIalrdgNecR9caE3LyJaAGl/27pn2691hzyY2ui7mmimc
9gSrbITBOJJ+5tWmzHnVtMEAPhx/wB1TLc4AWKEFW/+QTPQR8r97lTnQN1+Fozha
BUoK7cCxP4LCmfdYSXIDTML6n+xl/V+myUVsW7ATjl1oFIvpkw/Mj7Gs6spvjteo
uHHjfODmDKAMkLAAiT2/ymhLmsmrW1NaFlESTdQsXJdaWfjKtgZ5TFWiAcKvjc5T
HbyG6KYqm7afJUCsiwRW/E4W3RnHCh+PKJAa18wm6u6AhEkfJXzhZSxTYU9DgTfP
kMT7vI3Zm8MF8Smhbc/qlcAUgloGkNKqtZQFWWtYnilv0SZtFVv2ImhuRvcxYA43
8fhC9xc+/SVtMQwfa+4Gvyll+QD1hkLs17u39t1+iN/Nk6UbcobJ+LUDaShRVRxd
0AmlAG7xGRYGH17pSu/gn5BMqI4tH2hc7zC9dNU7ZiuaKxflA7GQukDgFVUp4JEC
cB89PD2rP+8LFXWGNyR0oOuH7Y2ToXf9cBag2yevJO09ggWJomh1BFIrAhuxRVGQ
QOID4NB/Y3zhZ0N8//uHUh51kJ/woJ/gXxJPKFCZgE3IB7QsQ5VxFi7zkOpP6YB2
MvIwWszbZ1sReGAqeJJTUr7X/FeLSrsBCgCO7B5BiOdazpehGgjBKraZP5Tz3rbx
MclqO0Cad7KGjS1hwp17qPCz2xRnElvr4a0Xe/Mn1Nj+8EapiAeLqxmsSDB/yLur
j8Fp6BsIEM7liIs8FEvI6fI3ZrqjLt3fIVACOlUcYTuqRgaK2pMSATA33mSsJEF7
i0f6wihgoMsr3lq2uzP3OSgMIE1festmofnZRuAQ1Znt926C5Q3aOtLUQqIZcoQ3
JXGjZJdkSufsq66aciOo1FkE31q5QP/l9NfUJejBgJRfVC8BAY6IXW3BsujtZZ0Q
p8GMZ6wH66EURvcLaylDV7s5022KtEE76UNMM2nTY74R3pORAJAmOST+rKljAHBC
2RxWexPAsyzlKB+7hFzk/786Mo1O6+7kgOFppU+U4C6ob80qFrixeu42bGpOAQ/5
30l5uwPf6OjKZb9O9sYye7waWzoVSFhijAriHpaIPUwAZmvvcMk2v90sA40LMCii
ELHpWO6QFWzhy6qj3tFrwdYlLN1ok40p2NK3Y1DjxqJfuUhvH5panrf5HLVDog1p
n8s6DTlv9PsUnDQXawzrqHngjzEBIy12wHhCRRRtpCG5/oeDnIobLyAmhdHfF5Ut
aOyYWidWsWzgLLWlLxeZg4Uued6hKbnlIsQ4VtCJvh+HkzNF2pXgKH6aWVxXWqgl
+j4bkbm2tYjY9JJ5zTYwcs6dxz8eguW5A2U0fVR25hTn1sQt7DxR+juEIOSfiuiU
/fDug+dkmlcwiMkpfQ++d5uyhho0GqO3UNlxHTKKCUDWSVyXI+RGOl+2qESOG5Ld
6QgUDFgqUrorMF2M6ggQKcno+S2QLU2tA2ggYU3fhrlMdA5J0hC8myflIJl0fdJ5
Ari5OUV0EZZjgqO54neayaq3ieTZqLJQHqgkXZ8QiAPE959gUgTMFfjxOSh/hfvA
1NZo8PkoYWxwa6aQUMUROt/jAqc/hsEC9VLA8+GCtt6qaucydsmjmXbvVVjOPwYJ
nQ9Fa9JU1WMTFX1z4iZJrXCl4dbS1ApS4RfM1bEkJZ/Ik3hUM6/YnNEgCemiNTia
QCu92+E6e9AlZmnqCGKXeE8dTaBJ6rvkh27z09JNI6Et2isVMk4ChOn2HCzm5E+O
iORThsZhrBoQEk8d/XzA8WvM+NIEc8Zb0Vuat7uM/QBKQuvmEu6HA1/IHi24llwz
pAv3i0FT16DmtzPgc2FMlCj1uk7L7VJah34fawuOVf8rh3q5dqsjKrf8FMFbKv4A
QbIb673GMUdpayQwFfF9S/6BnpUzqB4/9qauFK7wI4Z+mamkSNiHmc4SJiDq+nQY
g0qvIwpj8w6/UV8SjXlQNke6XOcX+/58DP16PInhXzqgJ3klSqc9+fZ2Hi5CB2zB
V2h9ONghZuuACFXfJ07LIfO6KKKBTJTW2whPlYGgqIO2lnTFwpf7joJYee2YR1/E
4F/0wG4hhX5ts95v1P08g+3yqRl5Pj9ioJ2uRoYDIa/sHUJWjWrVqUl5eCAybTC6
xIkU6brk81SjyA18xu+CdFSka6mwBUlzJwdusPQyh8D4074mit9ASKL11zmwXJCX
w4P9g5zvh36UG7ARE5w9m+hyiEGt5E5Pk0PE6IdirAEBdsKb8/sY943AT5CV37qC
qUmUTQzma377WGeb2Wa6hLkJyo7EUtTb5zwnOyzQX1cXuj+3QvKdkpMtMNwpRvdj
5nZ6GY9+aevnWDJnPJ60drcDlu7Bb+YtYKMYLYeLh+yOlUaGCsoutq71xDPz8HVF
1js8aGUdC3eJONC97SVombRa+Whk5gcRRQ5f8NpaTkgb+G7i23zKsgleQFMPZXH3
Y5DoLDf4b0wknj5GyD13Aw5av8XV8uoU6/MRzr00d2hsjNtADpAviqo06NiZLBlK
+upr3VMQ1Pc8TFRk2YCTtGLPvt4mvyBH9eofKRFlh0IxJdiWoQQK8eZ8FhaYivXz
FlWv0PyLnKC38Y46ZX2t0u+kVKP6v38NE9p6mFdze2f9aTBXRAn4krnPB0zlAGja
RIxAxAvOLxwjBEoDMML7mSr9ZeioxAq/AfiMnFQJUFNFDL9G2dtZ6/zS/3ZlkhHd
IK0NRGQEM1uKqn2T2yqND8RnAEGOGscYcTXt/ieVL36POfHMZlkShxaJxuk8ksvP
3q7wN0IQaHpu8f6SJ+2jjbazGuBfTs2sd7QOXywXc4y3oummYfwsaf98VRSL7vwA
+0EdDRAOGkU+x7yypr//1VdaOXqXfHAGlJlJ+zuZSPwk4fHWV64S+Vr0Q7/bjZQY
C+SMD3m9fyQR7hktr2RuYDtR390k1OqtD17hjXe6JzaCQ67cEYhZ+GSqnUh+Inlr
yFmY+Ej2THk2glIRu5nI1nLh+7zveuli8warXJ2cMYeJ5ZiMMobNp53+Nw0KmDvi
wlJAST1cvixUWBQW1cmu1/sksS8f8tKKr2mcIiPRYIRYyQ0m3iagydtcBbgfdibZ
wv8BmiTUp/pTMjK8RuLGgRK2TidkEqQkHA3jFOq6ZTqgEqTHjRImRi/QTkGsZizd
zTqG9SETD04uZpSg7lG0OB9e4MXDRzBtnhq9HOEV3ySRpMyiq91QdhZnjDEuhH0o
7XR8tZcHN3jVQmo8Qbb2hPDjI3/Kfx8pTtl8wDikpQWpQsDhVPXAWArG2MVFiqdk
mAM1G5ecuXIGCuCNg3zgPtshhtVQr6Vq7qeLI11rL2knjPVqGRqOrcC01m9cntn8
+htXs+tjWVXBB/lyBUQQZuZwpwTFcilLXlWB39LbAvIhaaOFgHj9j9KRBgsHOScP
J22UdiYRjEGJcOibEriCKtpOUpma4Ao6TsCCbELW3/jCfvRZF/u8dznJ2Ih+ynHt
z10uel9rad4PJK/94EJKgp5IV9x+RpRkZhpD2gjX01KGFGytF9EPbmacxIKtX9Gg
SHWIZkzmR6YFE+BBnj+R9VkW6aWUDW5O24csQrPrKRHKY4eFmR7MgFZ8ptJWGtS0
/8KYgOREdMlkZiMthyhTGQcsnjntdDR8eIZy8A/1byk1qI+iow6yu53K5GsRJ7FB
xqe3l80ohui7sKm1wR2Zjtnv2H+vnnh289TPvpPraAHCr/CSv7RJ9evoyG9OneFs
Q6en0Ajp5GvbjsgPbApuUYBZTLTDWSe/M6ifbbf/n1AbjPlY2fV0orxeVrNDNayc
sxGsIMnMPoaXCfcCFTx4ZujO+0s6LMWp998buDnVh2G5vAAk9Tla20Ys63glxFXP
dqn6/HYk6Iu/XegzeZbeF61rrGC0a1p5UWcKkmZymgcM2hoaZ5ToCoO1gUQUC+2J
BPviZdRcEgp4YjNVLY4HrWdqrOM3DAIkxbreJqHPsj0LjHlHP4Ht2AeUmOhqB2YX
KmqyJ4picFl0cVRqW6JyVPZNJ64dDob3R0YmsESHriMmSifhOOOVsFjdyEpGCrBD
LgsC01QzOZl+8PWn6SrX1on1WTbcNqOnTtCGV40GmxiiDgeqOkGKCVY608n8jWJL
KJzjYqOfDXTdwUD513C/DDhVTIMVuc77bDUFiMy3ZrQLCrTkK+M9sk5j6f567wXi
ACc77wM00oR6cybiIv+mol6KaYj6wYeFZ4tSRBXJKS6nmjwibCADZ6e/WJKOkvGE
3YBLgw4LhDAtim+xpAdy2IpS8Ljkbms7evL3lm26LsdN2tCTxv00MiM0UBjkrHs+
diBc5LZ3Y2SgW0nktm9D3eY/OMucscz1+bsFp1PH+SJhFPuTP1leIgwmXvC04oq1
mYISYTCThr95dbKKQSw+DB0JTTIQ9dwsiQ+FTaKwBcDYlllOd5bue4ZVbjN2VxI7
41NJDT5954GUPE6vJx3P8/v/eaCuaEjrjw67BQnw7OMeFyS36oD1oBH7r/C01DHd
lPNspY/PGY7LQgn1b9p/jHtl8SCIsXbokZG+PNbf8aQMXWcurnkDPTUVCPuBu6+g
YF4yianqFMRkG8k0lpwfwNf7zqf3fUr3kdcDklofalqraixiUcXEu+XB3IYE/Rhd
ES2rjoGbstpwipFRaU8sGB7OvLI0ufkT99fnNWBeGkTkA+BRu7jBEapx+UKYY/Lr
y+2bUR3KcmN/qSZsVLom2JpaXYcARS/MjIVMZGaSsVMx/gLe88j3sIU899p+gKrU
uazSoimGn4zQlIpmhZxcuWL7h6YhDoXpLSNWve0H+V3adWJllZMaADnA2V2lUnpp
aUqVrTbmg+T+tyqRePR+Ceu+UwpuqLzAhS4Q4ES67Kg9eqGqocwUGRypD2TV7DXk
4OQcry1cryJEdSeFdrv3saE7ZgQM00QW9rhNhZ5FaS3Ioo4JCP0iY8O3SqG8KieX
mAwRX3xEoMw9w2oE3mEmuJPGD3rZp4Gp0Tv5EHRgIlFiXsK5YIaN1beX5/ZSB3vF
T3ORP7lcUGpBHdPGgITw38rACYIpWfoh87XvkeXjq2WgK4cKks5W9lsYbMv6vfax
+taWnFnxUNs71JwUheoSHQlwhOiMOIweAilSYiEcEv7+rlQ9R9z8O8KpSzNtGQ5f
5VuLMqp1XRs7FicrTcpXZZPd8v2wjdUZSetR0FTBjAWLVCU2x8CDzZVype5G1gGc
hsIaxabebG2P1aE/bHbxHlYr56mczbU+bfYUabo3Hc+Ug43VB9Q2R/MDMg5R7OBc
82Vr7xCbIcueo+xrB2rzfpKo5zBimECSPiYmmDlK6hBJ/azoYOvizGIKhmdFkoCE
QvEPRt47dn3lGuPMNqAoGrPUppJwJ8u15xWuef8CB1ve5hVlgl8jAMUL0St+cE6t
IW+GX3nfq3Tva2Hzr0PppLT2F0sD+VQ8gX3zqP4iGn4Oz5myHXHK3I0zDEQd80tK
1nnYfgGdLuaC+Vu5ByM9VzIVEWuzZsBVDSW/u3rUAyU7viUIqpewh6tyty6Wr9h0
qrLwHIZhA8yJx/lip3LY6CFxhrZVcNglo+X1hl2pHeDUMkveq2/gH/kZSRV+87I9
nAGA2tjqDwusN7R1XW49VMrIdmI5Li7DPmhnrgfSgNvgmaBvUwftGkP+sE5GQqsp
CaervApeGo+nBtNnBS12FNtLm/2NO6IYqB0o87FiqVe4z1qrSnKLoNmMLEcobCiG
Cq9aCsVw23w0UtsQ/Vc9mn6PUmDJD1G1EQfMbAqcFttCnTtYvW9F/KzzwSUn91N7
m8JjmtfY9PZNaisqREMEM3+8jeTlOClBnNrAKZ+XHPcQurryI4npP6e/n57IU9iV
6azQT5yW4/4+1FWkJb5g9V3usEkOiot5TOBeqqFx2ujiaQTLYcs2wnXuv5cTil4B
wjq1MZac1MuDZqEPGImjIB/aOcCL8chrdTgwumL46FQcRc6Q+GXUOqxW8yHNqYME
gIXnEFzGsh2/MQE8dHA6tcvnuxusS7pfXkxJIsFpQw2+bChNHI/gar/UUeodvIu7
wBQoYnNrzGsIb9Zz6g5XpDvVxxs8FGUxNaKZbshm877Lhdj1SjN/2ut5Bmzug1TA
fq1fChjCC23N5yI8nuVJbw7M+1Ne565Rhp5E04kYf4bL3O3B/eHmILc5bzcsfFlk
xS68LvvAHpEEZdF2naT0xiSvquSmGqtc60RLzEqIh8XLOfQlxqc8d1DbI6ubksS2
J+XDYVichZljsTT1qAsqG+QCta9zvHBM3vot7cOPZH0+BCmVcKO8Cl2q84+lXqlB
IAy4CwaOhJBGHyvz9H9/CL20WcyJI0+f/RHA1HgoAqZh09X2azEujUcGkEvsxRpu
3E1TRKF88/MPUlRG4FteebSEctEti35swpDZIEUJCOjHsbyh93p3T2Ixizet3Gvv
iIEk4ei9ax8mlXmFZdGf+dWXKAfR0jlA0LT5Hm3BctOVOO22CbaZRbgB8pHxJqVL
EzCzQkLua1fYmL/6q28951DyWYQ7TbVj0kgVxQ6qwRpl8JBM1jG6Js1GdaNhD2Eb
otpg1m/U8q8DZTFVDvC0QLEr2rdzwB8wHVhBLrlnnuwa0ZG4Svg6VcD9xhhTjAsU
kSe078eiz/TVkssFlBGZWfAc7NPC05zJuXjtYihnlq2HMMHzJ8hwxefep6HbMxU4
0cYTNOZMSaHcSQoXlNsECxSz4SS78LpozgItE/qWan3KJMGSj8qiTQJHJ73UqBZZ
QOT+w6NNGKYEVCaaI6eBU/Gdac7dWwu+tN2AQMvlsA7oEW3uue2ITtb4GY5P6m+7
tdamjc06J955OF607PuBKyA8TT+jy+g2VO5gGzmMoScqsLjEwV1tUuJxV7K6XGXf
yPC8DHiQ0C3h7j8l4vL6zYmm0miL/xct4kvp4OOCpuu2arqcN1CWy4nVRux79zIb
b0QK3kr4eA0Ft5UrkYnwe7sRVGv7Nf+enbNDDCv6oeymEAZfC/Xkr/Z1c7d0y4uN
KziZRcA9/WGwkgQaPW4n+oBnbCbG6Y5rmN4raALnEerou5wXmtzk9CxxjepL0Xy4
jzQyvTcwZ4Il4slr/hqoe29jXc3xHHUvAVZaSqgUqnJ1oFkFCHD9oU6WkvZHOlm2
FITvlosL5KaMjO+9y2VErBBNRJs2NdAKgeGbzDOfeqlWgm6J/ZwuK5nv1+6y9jGI
xUuutD8Db1KlMVH3x3+aSlQGiZnoLs5E2h9aitaoN7qRJ9RQ5nZTnUgk0+eUnZYb
rwQ4Wtu1Y8NGdvp3VYrXhjbW/SUrRXImtakMBqtBD6Lzt+R06g3T2kj5PTq/MAmU
k9T2MJoi71+q36OdeRs8F4xF5plUfo+mHGtEMdKUrpYmJBIcFY1OHK7ZYm/SqJjL
9sUx7bx2XQ+GFNtLZpfbOQDzh/KAM3976oPNw4gKUROXyVepSfanOQqpc2cqIxQp
BKSgqmQoy+XnbuPE9EZD4ko1l0kDNxw5M977MpcxkIKWDZAORxGLncht7F2FFiRJ
ltUgfUgXpdewqaI8bepllwh6ktEtvmwzHqxFvzBJbg5fa+8+TKc6G4G9qdlrR0la
VpL/V9o19DMRDus3+t8bmLqr1GyU+LrgP5SIcyGoGQ81/YzYoTTNdz7IP/Zr82TC
6Qi3X08GzQLcYu1PCVRGmxj+idt3YH1zkRp0g99GSw2Ohr2bm4xjWop2bYe5DpXU
5OO+op5Srod76j0BjwJK1A96qUd7tPm5ALS2W3TWWdbJ85ucq5MEMXODcEA3bwlv
01926r2GXLjjO9gBuMbGxQ0vcg578jkDuoyRsaQ6wkxi43Mpdmpj+eSKCrNo1br+
nLFDcZnnUXYbOdirftovQAHMUd8eD13GZWQ3tZsMV9mMqdE8mkOv5xqmvnofoljp
2+gKtiPm2ucbZdoToA4//5LKdGp9PqPn/B7dbkNPggh4tFPwxiEwMdaPmYrPkvl6
Vc6XSc0iSN5DLFAAxuKYd2nAJf2tL9kqHkGejxeVSdiIofZlTxbwQZFt5eXSDgl2
grT51B2zzSigHRw+xRt4KGECAPepHPZQljkG01o0PRGQfSK8ZgOwYn0A9N8Yvde7
0YR+7iOqtF+KvSKlBbj7DWz4v0ciL6JiSgf2dfTbzV7qOFXVw2gqWcX3xOsYGB5k
T5kT6UOEFIpZj6fLodlbOhEzC9VMVTx/h18qDh02WX7XU7tsszTHM38BgLbVekAJ
BHYz8lR0Ri80oUYcn82HDU8CczdUEQgVNDsZUzzePqgOzD2yN5eT1c8Kn8yyHJej
NRc/s0u1KFCJF4Buv8RrOtPkPaiMI0wLKyvM9Wop2BH1mjak4lWWPGlKha5N0YkM
ZX1xXmvFkLzTmHTwdY5ny+/O6XYpGF/MNjdRRozZw165/2m/XsHAVr6E14agt2GV
2SG7fkdTf8rldLOoG6QQUC2pxbZ3ftpURP2P8jk556WxR8ZSIST1fk79/ohY9tM8
lgRIcpcMy7chi8JK3KIgQhSAfTM1mldEF4gb2XkZBjah+yd9JCitlznxz1Tl7Xlv
Rk0mrTQmrdN1Ce/5E3LpYOSHxBAuASyItdNOX+rF/OYcoE8Zoh4dVEK2fp9F8g3f
cZcFmvgLLFsufTYeAZceACS/lu1ZJqq2ScwOGqBeqrS1vZVFgei9JPeWR+XyUrP4
e9YcHYGFXmhxWjwyN+lulHRMpjPdjaHtRO0pm9D2CyXh5mfAirNYN+0ZWVlfY0Tj
v2b6BsvWQHx/j8vEJr2JP4q8w11X1M4cPghyf0JgAyptC3Iqm48ZWTodTSqWXRvE
x16pCEWqD26Rx9KNAB7rhXo/21vygLLw868PBIm95r3B8NgKcOsZtSkuwwrfCR3/
UI001WOSFwDwxcuQVTCfit1mm+NHkHQnnEr1bYsJ3R2bGcLG7f0DqacEpQZiVzvw
i/3PGeEOyZcIGA6X6MdoCoje8XGVd9pYc8g6uVFfs6x65QuAljfa4/MhF3UycRwx
j5WQoScWG2qz8LeUtvDViPk4jZOBERWNRzMy7fmQCm+hrNd2FvSCzl7D1mIEA5l7
J5CduRt6RKv2ssWLtRa//Gw2hKUBWK6gi0IJFwTC5FrX8P68L/lGR6wiVtvh8M3p
Kb3QDkpxXqGFr8iVzcV7UZ90cuMNLOELqdC8UHbF4bi3zRm3qrRNq+lymOlbGEfP
cH1FDesCogc2BQYy1WwZDTXvlunquw/TDI37snOAigCSULC7xaoSfxXSwphYXmpp
n+gulutfQGmgWazLurLPYqQ5Eo1jvWDsYrXmyXkIgHNCs3at3JKv8ruu5EaLwaKP
jPa6lzB+Qmx1brbUaieQpW84oAs50thMc5adjxPxBwOvgLVIgPnIM6+Hjcnen7AU
/ulLpX15nS19nupytXNRKdVnHsDilWjdDnySp4qjAr32nVX/BexuddX5auYnAJ+Z
hTs5getUboHBSy+NWZgkR2KsPdGMMvxjGlz9y+gISSpEpJ71VQt+RM3cp40MwERF
zcEJhSXrPcqcUy0UJNd8amDtX2BH+Ez+5QpebGtyW3qfpty6btQBV8bkwAi5UChV
+fLOeo7hwh8f4CfnPlra6ldvBMPRa/bLnWuTtOcghQKtLZ/YRxRSmTU8aUxu0e8k
ZqTrC1ZyZRPrc8bc3VGqTo6+Y0qXUPTg0XdWeV40Tmd2KJsfRm8+dTgY/PQxQtQ1
3cMiRDwjloT0bn/4zVBklEqenFecriwlrnk8WX4LPfAFNIDXg6dlHBjcUI3CPW0A
cOz6Fk8H9lkFinnMg2r+QxnEpwenxfps+lM0EndUmzOz/6276dhsR4Og+/PGMUU5
2C0ahvnksh4+n54AesThOLgijhXVWxeWs50thdGxSVF32d3+z+WnxMCFD7Fpdner
SMj2HeL+POaJynxgR4LqcjET88/oyy8sNrcT10NkboMPnYpF3GA7iOzO1IvNJ6F0
PW98lz3xOOhG+EEbXs8YhBb2kEkCUiwBcQTm7oe54Cqbr923/cOLHhkyRWqeugVi
KYX96uYxuwmVbWGPsMEN/dq9sQkUc1K97AxGdb/x596WCvnoU90uNXNMp+qi2RaP
RUcGdb0yPvKmPc8o+WmGSH8DwnoIOHbZPV7GJ9QvN6X8tduFZOOmZd1PzaXerwzg
jaylbXaUUgfVBTEYTWbeY9BgACZGbPiTwhHOj3DTen06GEReQnKocudTotSLyW7S
2tHG8zmbmZBpQGqGxLmuBTikH/P0T3LcWsa5pyTpq9iWwxc6QXgfVO2yzrx6e1Hh
YcsGDO71ImR6aOp0dLB5FCeFmZzcGW+/1b2ayga4V+ugQmV48FpolmdC7R3xE8a7
40wO6koIaLOEPy6g5cB9H491+ExGd4FBVU/TCGdp4EUkZlHz1bOo91g8kAGcvwqe
eF6OOTJQx/8vmlYcgoAtRRplDVysxZRDoi1vTgzhBV4AgbKCwdGQTNA0sdFP2OgJ
TSgztC9M7BxmfbC9hBCIgsYafhoWR1WdnIh4rqcAuIJYQ+Iz5HoJJlZjUDKp9AMY
mFFVjw+ZfCAZQwmXvjoqa1Ba3T0s4z+D2jxNFLGk7kmsFcF/SLEgqUTVB9BRGum8
8jb0l7sZeTnflcz6VATAGmx/5citCnlirhzN9zHuy8OzM3FhCh+zYpytThF6xwwq
Jlo1JdPEgZx0usZApY56/18q4L2iRVzTZ1DbusvbG17Zy70FRY6P2wsXk/fr8HN0
inA1smU1jY493yh6YIbh07rAT4JHRpB9Y4qY1qmWyheo5SrRT45NYLU+uW4UeQPq
scCqbtpJzz6BhtyVbenkR1KPdhemWV8GXeM0bPCLj0ere1pnN7Z3SWF7pBCFNs/T
2QgP8I39wj4THe+kogrrggd5cPIhB3G2ev243ny8+zu8pIZ4b233y4TpkUNvi1JK
0S/8J+MPmkerhNWR15WZMVriE/Y1JC3F005OJfwRbfRiPyGqle9p+gjlXVTZ/mxC
ksM80iiHZd+50W0uBeU4uHLlkGAluwp1ZqtEJlNmKycFkyqIvGMhS+P0EUr4+uof
Yg42sg3mn6Q3QkQmQHbJQrjj9FbEGNiE/wl6+fdoBFd0oB16lkhMgHWR7ThCPVI/
C/2BJtkHofCPX3/yMwddhEidB6J7mYCoJpn+zNfoK+7DOOqZ2f9RFpq3yxxHkTdV
0LGmNAIjWwCi+NuIfww9TsRM3DQTTaY3lRJ5aypKuU+Xzs6p/dO7sGkSVUI2qw/w
nyl9pCWWl7MYDoAREZeCnE7qA4YkA090bxZFd1lxbaQQIvqDCuIFYa1kqgBkp2Wl
Lra81FT9wUfN1zmr18pcApi9n7WEeveWjUIunLdQYN3X8s0ZeRdrypkZ0aelXJjp
E5R0AFXu/Hd+f5gi8pMLJWm0Bzw9061gQEfRCAj2fR156C8o4gZz3gJ4iXJQn2Rh
tN4ZGt0lFnhrtHWAfLOTTDf8gmlU0hqP3H4L2AHEbdJ60YJQNoHXCMIvUhao5DML
ByjWBC2xhY7CkR+G+h3RaCW67BsVmv9+nfqhb7kcABqN+xF6EuGmJjWsXD/VXLga
pyhdVwLMgBWlEf652corliFr9v5WKx/7aoqkFVVT4LEFSUIRH4OTpNwHPIa8JMLs
Y+1hsCR2/exAI0ohgH/5OilhlkQcQrsR2WDhny02tTECsu7lZBTKEQWv2w3/Vubb
y7c10LPwq1Vcf7yxTgvTdV8CMVX3m61O5auPZ+JtKbchZQzBtxCOF/68LR2loXgN
FOao0OHGov71rBAhjrElDjCboH7YcfkvSLGuNDRf16MN9WGzFaYmgvM7ml1HXcdu
5tlnCDVJL8BZufqb42rZAIffjqxJJ7Qa/wNeVM8VEqGUx+/On5T6ISTcls8+b56m
997XHgJFd9UQqp+fN5zBHrWyyBfeA61iKqjbip1+UXgeGshCp4cvuFRecE0P3Nmu
7dgRIchlBMlITegxwTK3bJsl9HyvUqW6CMp9Ht9Pu1fhQbpRDMBvs6V+l9hSSHeP
rTAbLnBARzmkm2I5iGUHcApphn4PkO4aIaFSVv91O9kv0//hvaR8eR/T7lCEXZ+a
aL3ewaRN5pVR1Ru4ah4p6ST4UMcPSvkyDzDzca5hZhjjOxE71hzmAXxhD4qczEl0
CBpV8L0IqZE55y778ML1AXyHE1lci+QpWkWDoFUWDao5Nko2Zkiz3LcQA7qQxuxb
VSMiWC/9NGpqa3ZWF2fFATwgNrQpjdpkMtYkUNX9bgiNMTD+AgQJXHYRVFBREuN2
4buhbWseYTlKUV2iyoIPtKvn/DznCE3IuWf+1md+VgiQRHfZwarnYgIfqe/DEcsu
fhad/07U0/2Ug32AJT4l+eqs7twyAfd7G6cwCJE1klKKUu3rCYrlQMY1/MuL/Uy/
CExbCNfaQJphRQGZmHgPPTu+OSNN6bxV8MdyBqe0i9d4nGGIUUg/er3KuGxKzLO2
+GUxB4vyaoDEN4L/r1EYK5nkhj4mah/L4L8duvwoBi3x6kw+3t8C6U5E21NsVk8r
7k0lMbifF76++GHX/pyjPI0VEKhAR5svrZbjB/ybFArsD3HDtWnZp4vvZf2VvXyt
QntfluslFFPUiHfgC/MoBM11tkVsBZ0JX6AzGRxyCxSgX0hbYyY6gXaJ04yELVH9
r0/QFz/ZM1LUYpEy4TVCtpTtn1EPzOm9Tfa9sHmfe9qe8mErouf77nn1t9BqJzFN
aOOu8AhdaC23+5DPROYxoCOcBNQEYG9n5c0eVM3tb0/akD9aRIFTeGSzqdZ4jMld
3pXN34TKyIc8hgQ4MJ9rY4G+xGwxNtXyp7vkjVWS2FH1yPXH21mHWAUPiyCF5hbL
1miGL1gvsoRu9X9rQN97I6G4UnB1+oF0PMCtIfVrvpqXVhWpbDa17v/DTkSSualx
qid62IfwX/Ftzoahfi9OVRNT/+NmAq52hHwZKmDZ7Lt7A5D87G15FkPMkDtQ6N7E
ZMyNCssGevfih0B6HMIW4SsawI9Fx9hte4ya8t/w6gWYENoEreQi/Sa6IcvtLFSy
um77GztGpAJh36gLZAZX5PQO/mItFiaAs0bw3uAc4iGeNCQJahRx9qPcwNLdYdon
cu9oHMsRiXWNTtOor0duwIcxcwaMTdO0AoXiNuhOy4UGpworKYGI9SX6iVcRjeqW
6DJVP0ZyujZ/O6xsc51NQwXxHwKJq3s2C/oCxU/7S4m+V8GL1r3HiHkrHz7PqTuQ
mWFgjdqXQ6GKTss856rBRBedchhSyeMpxVBWhugwE9pxBilhEDwpL27fXcH2/Rxj
qNq6jPK3Cc/AZomCRsSQKw5EJBei83hwPc++Ot0+aW29XF2GYZe9oQXUzZ19QRW6
iuDDttWQQ0DS25wjunS4texoNhbz44gWnIeo4OCjkCB2r7CSTbBlxiL5xYSICX/B
Kzt49fujqvalXm49Hl0Jran5st/+FZ/3BkVMiv8u5GTn0INsQKL2uJrYjwC0+qbC
NSBCDot0g9UBgR6b06OVZi16+XK4n5H8UaD10yeivtOF3L8wJY8MUy8P0II4DwYy
lfJjWn9cnrNQuI57JRjxV9ffUWIm5On0z+tnuOSP4bQB50dSFENQp7IimZGGfcP1
jqczTi3VnARZ4Nsu1zl59oU6bQixJdIcZ8+Dc00KUCRjU1tDMyLbYfeK6T2KvTKH
R3fyMhenwsFtyLIvdHubO1I5Ha9JKI/Xpp9QvIxWOGEOkz1xoG3aLOBRfgF+91U7
QqlCCfsyyplMMSMQzjPmQQ6rA3jyAr0p1VX1PmBfR895pXDuZGaLfjObkn3MBbwU
phwMdM3p/uDeRP9/WNDvsfJufBR0UClxpPkH1zTskKq1HpsoJJYHBUhEB/3VP0wj
+ebXEk61WVhzLo9+F+CVG7C3XvAvU4t3IfnGLVTEHVH9ajFQ0XPRoC9jrKWNXJdq
YbpF9wIv5Uz9ijZ99Tn3PezUUyJScvgXHTx6Ot3ukYgPApfQH2c7cje1SuIJpvwU
nA7WTTQpbcmM2WudbdPLdFtu6G4iYO1p+7PYdG4v/RRldQhuW5xPiwMX4Pws3+Uh
Jea+ID0bHhR43xvD+u/p0/e7fHAWkU3PaYKE4plMIlaqL9Mooobk+FA4Ocsa9JOe
O65KEZ7nasyh9RufgpRmlzm+hI0t8S50rW8awfW0mD+qK2kmATdxpeXITls3uvIG
tBeZxU5NjGcs0dglVdM5rTEgyER2fy0FyAsV8oUEaIIwHjqVN+A0BpKS+15pjp6N
/Xl8J0PW8/bfhi7O9S3GAjUEh8rpN3zAPMNy55y963BA8WEJzMQZcc3FMSg7oG0O
nMWvKwk8GMwmEVNBtuCXUS9dcg3NkwoxRzT+aiJ/ziDjcOWlfy/DyB+vOwxVWLyh
G8QY3KqBECq5Sfk6ZAgU8TWlweUzjGF+qzSPda1lpOWlMaeroI3sGdHVmEyDG6gL
h93tm1WLt6QXl+3Dn8aQ12+B2mXHzqtaTJF9kb32e3B9XqLj0OadC1oPfTGI8E+2
OJ4UZEQxcoEOmE96LkmWQLKEm2cXmXFG3PCevpE1yQnPitWeq9ceVM2pMLNTgwlA
oejt5a7rfd7QaHxDlE280AT3mto4MPmx1+HI1inBdlYZVKXgmjmZywHkMqufeoGV
vsAWYAW/89VjVpaOHrWSkJuQPwlmjGNEiBi7C+ULC779aDUsV/mbGRFUiu10Gjm/
Whk4umyC0ALAiv0iDuTgtlrLH+RenGeawI6a/NtG34QJ5C/APtej5+OKBHcHvtBS
grUe0SytEIt68+wlXxAzytiG04Z0npQ5tcZlHuqa4BgDvJ+qgPbW8aHKuIdqCNZX
QrsctlcbbvFwP3Fz6JURITO4veiqbUgO+zthGL2NMSEFzIO6j7UywovvhitMCvgB
SKKYGU5KujjmQK5R0xYvDDBbVMexyZu4rCPUHlvnDAvueHs8EcG2tdpam6/gH95C
it0wmu92Nay9mRq0xTKMMPp9932u/z93MfsZDUrmRKinIi5f1xjVkFT2CTUuq3xm
eIX7oQo1jPu8k2uxGtqledkR4d1kY3S2mNp6Yrkhmz/k1BrcPbVJZidC2pz5SzBD
z/tWkQ46dWgrpMTG3N2M3EqIKFWy2oH7x7xh1QxTOTeO6c/sOS+iLKYl7nU17oxX
w1MZaKnqlJP0bj5SVGjkzqY4Uk3Hyhp7T15+4aUhYLkXa0yRa/LV2Plbv/X2C29Y
+L/9YXx1BF18ZNi6A5WLemZYG1SApDzQasiQejPwutl3eFYsPxx1+saGH6hdn+TL
fS6WIDpka8kqCoNHkndGvWu+bbTpn3D2xLoe18g0NqAWNeKLZxc69mmD1jPT/teW
UOcxyTM1EEOCQ9ggJZtefbmuhdDmLcOBaYbKDPMw210hQktMLtLq8Gt/huk+qMFS
gtRJkgta0f5TyGxgVSOtBF2gG/dzM4vBTABhgYgDv/NidDuEWXo/5KDE+bUM87Hs
B4k0uJGjd1JQrlZdnwgybZCv+eMISQ7WWra0melmop0M+0yc7owOZvXdW+pzCD+/
BlmwTut9CM3U+5bT0ihXReMINMBgHTGFH5ORN30PU8EMd4ngzOSiXFk5Cv0/T4MD
YED+J5xeziE0LFJHIdnedfquLMCONZHbxnXZkosvQEXmt7+izk14+g559jm2Kh82
BFMPuYEJKAhNuSNyyMurc5n9dIgnwomKGPJcc2T5MYv9ADL7QfUrDuRRdZnfU/PJ
sYe129dOq5DBuI17syjbqDPeZ0LLV3kAR0S7tItIH0/q48zv39d0R8DXPAbfOOLO
asDukkFjktSwmGoWLgANOSbv4VekYNTdeIi9a7AKh79vQgGLsqvBo6Nzg+w4Lo9G
Hrvze3foDqLR0+1LuLEsxSKn9Y55l0/XEFpuaMjyP42hfg1Ei3+432YNIGvMMw28
XYC2LH3kPSHbA0RPxT9fmlLHQNlMg1w9R7FXgAFBrQYDQVVviPOoq/vb3Mgvi9+h
P7C3esYpxQZtVZl0ZD28NHosWJcPsiW7SBrGxrM6h3SJkgSTDBl5EwLz+YbmCwCW
CFRaSWrhjy2fut0SQIvF2qIKXcZ+HcDQbkYgvd/hfhg3ckglrAVz31MQrkWrcUAi
k/IPd7rYxcZyPkhhgG93EEKg/0HaQfhvlr5Jd+/cLu3zfQlJbIcviBHTgP6/oc2w
4zSr5S1nRJF7dBzHTdudOnFAKkXxSdAZWLEP24/Ng/DLbO6PS+4StnWWPmyZXESU
yVFJm8zVSGZszenqcLWCjozBRTgW6RnptdabNUeYjQMSO97oilpPf36IMXBJOu5u
wkTAoh91SxCRClOdlC8ipdzP9D0JEuREwzKnVBoNTAJAFykqOtr1BDpeUYs0ZqcW
FxY7uQWLOc20U1NCOHuMxwjTxUu9b72LDxbIXgmIhvYUpMulbNHYmzKLwdkZ27Ps
uQpLoN/Uav4T0CzFbkSDWjZvMXvPokIS0zA70JHgg21Cc/+5UW6SzY6+zL6iF9YO
jvgpg9Br3vRDUP8oawt/kafAI0O3tNfmmWGN9M5yHGkd8QwJn1KCNrJaOqp8/b0m
aP2ET+J6QAa+ZdILVcV/5WNbpj9QPTrwYM86SPM6/1OVwa+shxvjhHPZztCBwBPx
P2YDoj6Q6hJyvROkOY5r7W3zKbN1K7TevihrH9AHfHl2UOmZi8+Rpq8qIzI1BO25
BzBBTVZjxCxxNMnQJXkImTOMPgrTUANHQstyNwX1ERkgIvn/c/nrZtL6egIVW59w
fCodhQLmA5PXl6yVyVVKtsT6jUssamf+SnSdIjC6QeiEhsARe7eSNgStj+hgRiNh
MZDeMzALs1Hm8o13pmcG7BIODsNjv2ZVJMeNDzolP40byp5kyzvFj01Ty4jD4mfU
zu63/Zu6q+fz5RUSmX0lHnmVjAYkZU/+AeNqH1TzlIe5YKqyDEOJzO1DoARVwjRC
tXqF4MJ4TYKBBpZA7WkvWlTK5r19Av9gm8nH56hwxlmsuYPfGSZVa+0ScR846VK8
VbYbweOs4MydKX2WXMMyY3JJNmeWrWDwAhrUkNZIdAKuBA8pYzCi6P8Z9GbcxnMD
DOEz2zQ20RujjZYv8+0KArsQyiWP9OcC4etyNVsm5jNXV0qkM4bYIr1h3v7AANzt
eyhf/IHB5/NrTxK1ceefLPncwvKypo02PqhwMlNHnCdPU8Upjt/xz0r2FRt+XlFO
8ZqcpI0kYBvgSUQc6IOvL/YmbjGEB7A5YFUTXMXBFf+xQVmMNG65EA8V7OVuWEMp
Do52Ce8IsaeXwEYYDYPpSZo+39UGPTgYWwbCrCIFDMy9Tcm/hAlEAYyYouWqjX66
o5/RGUDYRDq4bDCvB7uwr8d2j3wFSeRXckj0HzOUa6RdgPMMKE2RLg8JTLNtV6rs
Myv6CEuYpq3/9ZKq7yIfqB7CKtkSgJw26ZwObCm0eONYuAxuMiPeDPJT+mZHCGTI
pbH2FlF8poM4UxlhOFm3NtGMjjloLrSWDpsEuDjhvmqfR5WaiQ1zhsFXXJqKOCjd
2L4/H0IioN0/MpaTXCV6ANrVzp9imPmAgLP7CBfrcCd2y0nLQ68vvnaXS6svf2Ec
lSum+3ValQ2mN2VmjcjvRDOTbnjWNqs0PmJLKOwE4+F77q8mclRJjL6GZQoxEsxU
3sUjq07VBWeHKL3+PAjTjPsRLsrj+3qMNCyMgVp+S43b4L0XX4kbRsdyubEd4/zP
twD4rCiNnhH7qh4+grJshKK52K6lonY6mgit3A2CLemIro+YTmyFpmRbKpXTGRMM
ctCdL/RBEC9A7a7ysQnbO2KyzbE0zHEvtD7Ju+gZH1xPprQJ207hj31m8DghkBNr
rCCmbw2jFDe+WnIRTPe0ANphkLDgNBDTV8VotHXbP6DAoAn7Lzulb/2Iq+fakORb
7UHvXeTmuW81XLK5231d6EFGVkqIygnepdvJwf99MH/hfRTainsTT9ZNlaQ/T1Zk
wEqRJTlhoHx9vI0rt00W7RTxtbEZMYsnD62+Piyc0CXZcjdg2dPbUM/e/G7q+Aso
givVk4iar94vQeNnpfXkeCNCRFhqaLmCoo2mCJ8DmyjvpBiJh0ysjV0afRH/4EYA
I/BOKo+kquscn3mh7pFwQcOwZLY+tcPI+VCN3CjY0wNEH60ARYbLqA7kzz4JKNzO
LuRhgQFnTI0zT9+ppF+VHdcAnQknyGtQ6xb2Yh7gwDft3r/8TbqggkVsWqg32v0D
O3/968XhVzYrLYEphTvBA4Jjg4bYl4YUEoCSDrFB6j+paW+D2Ljm28v1H229KyDR
djvkHz2dgQdNP3VT7jwLr8fJZYDrBcMWb0/wml6BAp06BHk5iBkQ8Qw3eXUThlro
mhzTAGUURFQmsDFx+X/4zx18fY3a2013O7UE33wgZG8cbDSkBHktqBBVLAsND18n
Iz2YAa0Sid5K8Gq2kDMxwBCGuut1Vlwnkf7buxKpaVNBCPva19uISJhf9aMJ74rk
4KJJITfCUw8nlWOScCm4SkfAecJdV9XkV3BNvU8/exckpKWRkxSK7oDgHUy0NCJF
jRppItCrbtowsXoljK6YI8d1A0bwcPHgDhuCX5cGt1EqLrgAYtxo8tntuXwz06Cm
fNb1/WoRlOm1X7wdxXysuMtgjiFLNB755Mqejz+74rEgQ008SCc/wuddf3fth5s3
ZSRNHYiODvhM/nIfOU+Dyg3M6bmlj3TWMfKgkZ3EDkjKx+lpNN6Yvgeku8/ZEpLw
3qb172bSSXK8wnLk3rvfEd7/5V6WU6nTmOw/2BzvLtdq9ag+rPk5R5/kw8uE3+9c
R8k9LXYszLy5Cy/wEQ3Mn95MBkljiE2ZElK7pcn7inVmEWwW9gO5nglsei5+zLeQ
oJ6drUDLFCdJTAxur8ZEYJ1TBprr0JKqRal+sZOyOEZjravu+auXYnveLKop6oj7
laBFY/5iY0OWCf0VvwGKmvUxrZHg2v0pFUrkch89pOF1E/kEpVEf6k1HRmcrW5ZO
SrFJtitv0Wol8qFiQxyPmJkfsuETBJR4tNIhXXONOd9U8gHM8f9IQk71qIVzwEnS
1Jb+xtJtJg5Hya5IadDpTovlEXB6Q119ypn7Usg1GNCJfXwK01Efge0sQumi5rZf
WrSqUxlL9HwBHRI4qysk4iWmMu3bUn3uUFZ9N+/Nwx2Aw+puf2cO6Wipg1Dsqz0h
WcJ8QGgD8X5SAMkcwcTKoxPrS9Q+edu1aNlulNxyECLz+f7Adker6kE+7mVKZ4VI
qHDhccZNf18xl15opnQaOD1GJYnAzoWoseR3kzAPik6tUerWhlH9wAYsMrr2ARRs
BEW99DgI6iwwSzftaDkWItUQpR+jQMsxexcTYSRDmwoMcaQ93zrFndycUh2DoRXI
MZ6D4ygJWlplA01ulQ8UpW/YJ2LEHLGTB5oIr1J7g95S0F7Ml2bQDWnmRfsXb0Qn
KZqwa1yg2NzjHGPnwHQH8p3mEiYI9qr1w411pKt4qAhQx49mLaJLg7yunitXksnb
RefctPlKRFxXR3zxqGYNZeb5RhrGrV4pW0siFKWTss9CjTte6j+3M5vN5FKbNDIx
PqAlukK2OHQW9i4SPRC7Q98r8JYmGB9DyqxtF3rIF0NP7m6/cIIpnSmGs0AJdYE5
2bl8IDohT9kjCTa3UIQNw5qWInpzvtmPzaCGOUZXkijmK0bK96rTs9nktknGLcNr
0UMVKPGilwjcdElj9i8Vk+MFc4BdBgqYQ7Rzwm3W9ovWX/gN4Juu/oyOj6hpRKie
OoIXFjwPU+Enf87tM9CbjyQ6G97p5Mg/wuffmdEBQe2MRVvtjo1srQJ4Aedd43du
DhrgW3WSnp4LWrSKltkzhtRkSBXNjGvuXVTzPBPztf9HMUj1U7fr65szWbhzAvh2
VT7Yu0zrfNHPL/v+kLAlymwfYNaohJbJxXe2ZCXal62b+jBmCcpkfgoWbgVmfqbO
xwL6nN8Hx6e3ZBbOYZ+cztv9LG4byBGrxxq7RxnVtKvAs6AsmeNsjoJ22Xh13/VC
RtfcHZRYvpbBwjCA0BqtlqSnCSK0bsxUa3DQhjJC20r2W2BVAi6lmG1i0bDpIijc
R0yIOfBAEDVI60tHed3zSjbwlpkQ2oeHJH8PYqe//dI5HWaiwvDX64pSgKLnVRmU
MgeOomupfTPMrwfR8tCOfcoF9dx3tUOpa7vmqIE2EPDknJN4dzoELS0wctgaPWQc
K9T2bQVTDFWj+sYEFZPDj+bDExM1QpRGz00ynXkPcBpLLYmPrFS4ft7DbfDCHhMJ
yTpOluBgVGi5X49soaxAUEjkBK+aHCR64RH2Z326+mu8gCLRAntZ24ANCIRQgmXa
Z34Rauhl0EhaVub63/GKgMCzbknpiLLEna9P6knJ+jIbRh3H84AT3nDjbkFK6VZT
gPbbU0Mfwj2q3MzlaD0hICghLXIx1UTuJgxH0lQA/IbZVrik4WVZrDOt/RfMDo3r
AOFCNWPI8wIVMwGfz9sLoRWsvqwtlemkCpIQ/hAiek0EkzlVyjIdHLT/kOI6j8J4
CNgE3sFigKURznRGjQETU13rafzqVNoR8YONChs6cVYDOpMvYhe6n/MWq6PniAD2
g1l7/j/YEcmyXgiDil4gzYh6bkd9+ZU0AshSzXqIito9iON296o8UjRsUVRIjZsV
T9iDbHs9jiy8QqCdmH8dVfuaplikYbzGFyG37k2qudMLLkjvUyjUH2fKxWNkHFrZ
MmlEN5KYb/+ES4YCyfQN5UOqPrIFtCBkIuNoAqXy9v4D3f64LC0DhuMDle2Vr5Tr
HMwVoya8lMT8ohfEISm8+qKXExw2V6ZHR0kgnoN5qB0vt3NQvCbFOKlcMiHZXKkF
5/Alfw+hOB8ch6avudv6+3dL2aCiFNOd49BVEBit1wnpCzM3AokJ5XPU73gaHuqL
CYM2HD8lkSxFeqCOW8SJQ6SUFa5sRO8tvVZwEn/tRKFAkrR3l+GleZubIIjHVxZo
/ha/438BysQD7Q1zx9Segn8TXq7ftA9gc1+3+QCWRcY+xhYcZcUuE2w6Mh/EInHT
oi68uOKN5+wy0isIX5T/3Gh8vpVwpQfJ4EwCpoCmLJjEndsi64JWuSfwkguAhpDl
i3/4ZCN7G4mWerw3fM3pOIr9hM6C2ZlbmFgnWpIJscNXzRRH2ZelqtplBoNIAKlh
X74/T2g8w+UymvhTkAa1caT80XLnH8hKb2RtXKVfR07+riet4ljuNP5X4/pQMl+G
+o0n0N+KRrAcHr7fhWHUjDPs69UcGARkTI+lRoVC96/TvrqdpELAObsgsL/vySjH
4NgmB5KMqvXDPSCN3rvOOGGn4n1Af3Kr06z8NV3cdVp2Vzpmg6jsZp2JU1VhSxaM
IG84fUg0KCu7ItshWsZ2IorsvEoSz0PVLtwVwObp4nJGst9ChNL7E4FXSgj5g1+i
txBA4SjG8RBXjoxU1KEcJDsIxaqa+zjxwwb00uzdEm28VYWTqLf0w2UdH6ONrcJ9
KKHfT3oODdNC+yhfADJSbdCx4BPJYos8O+Xd28yQbJ35d1XPp2RHYejnFZA1CPuG
KvT5tBCZI45wKuCUwm5ah2bMgnEd1PIyrQCF0uKqZAkV4pnQ2YxU1KOrm3YV7jrJ
4pVJ2XJ+Ac4oz51TjTKvuCN8sF6ozUy9ZyuetkR0v3TRPgcwmKdqMeIJnxZ1bb8k
G3NBSyZRWwxiSrBWORyrm4ooUryQoLyjQ5793bNsO/8OZlAuoyCb59OSek03nxpz
BHwZfwGwhACceY4eq3AApazsPgbgXJgqJJKly1B/Sr+c0LvpLEXo+XIxHdZlXv5p
ajV4N/RPfouwWXzne4CVpsPZydd8xORCYw9QDQHHS4HUoTPmPZGb5I3JGGFfRtTQ
YuP2C1omNk5cgSOBW0dudGU8tK4kz75BU4/Wy36RSacfVp/ofz4b4dpwVbD4hW03
CjXxEDrM+WiRhzKvBhy4BFGy74A1QR5oYfVLhW2MQ1+d4v2wTfbLxV3BOAfUH8ts
cLThx8zW01qlaK8FGlwQPoW+c6r0rcHI7vDpalixvGsOrZTF1vCWxEKdkyCkCVal
RKfEWA4wnDC8yuTGEz/zVJJhukW6qFUKrpzUvr6r+TGHtoTpf+MthwzDDNT5dhC5
PE21fnWjuPDRWTwZLls8ZUyVOimT/OZg0Y+MlVVDZhefOdju1b6+41yPtwJtUAWA
vUBKBqzpjJqsTZ8WX6nLczZTLdM7bbTjU9Ek6RHI9rCslYPQLPOFTma1agFX8u1s
hKmLzz3MjufdeC2w4JpKpXLe85ZZYRLo09G/CjqUNncBlGbwvac/O/Aw7xWbtHlf
Izc0YvlRvAlClST6yefJJiYtHg9w4QXpDxfNyqeISv8HhHVffRTm/RfiD5F3Fk44
qMNWhTudIp9/Udv9kkMhDRIjaZots6yP8WVz7wYT7GPR0/40s2Z5nIzH3Me4lqEI
wgCoct3OsSCgGBSi5W4+fFEc9/YisOWfbfeIEW1tVQDAfPFsnboapIhWWkubWyi7
5NV32R7e+vBOPOxvhJdH9QbHZBTMAQNXFmYWvx5KIwwS7SJzVeOeFXbO5Uf0acPL
8iGHICW/f3hOlzlPL8rE0aDyYmzITKQQDNAin7M+qQsNBq4MOmIFrxkx1dY8sWQX
HAJd2oFR8ZcBVtFWOv1pBW5mghPiUhkOYLKmdRUrcaIUSa5rAdMcUO6lq97aJyXR
hUhwMdjRUHG7MIggeyAyOslV0VN4w1ZszOevJIHZXLyM0TelHnKVTtMc9D8uCck8
SJnA9FBzYI+JRGNQUG7vD224xGXp9L2zGHNkDXf+uBt4nug13GPwRnTvq3NVNOzR
N9a/fALlDOMudWqpFT40+EHsYImWGN9fsRpnB8pjPw2LzL/iZN8vAcBAg2CIxjqI
evvjgllYKrfMCcwa06GdEAotmZIb0g9WN4IHm9fT9gsIgiTd0HtU1JzmxbBsz9IX
mAshPGNpODlmTmjTqN8rD7bNJkTsuHnNELwG73xVh5xEU6xZmSnegrKdyeAkPzgM
/ygseoSgrgcQ/W8pTAkBaPA68W0uNeLoj/8/+lTixS7IHfqRrOu3iNiVCOmdy6mh
gZ0omIkn48ZZTtnJtgWNcgsocCZIFCC04n2As1SIxFoB5yoekAQ5WtvnF/WWk30e
KGhQ+wRk8FRW4fMYq0RUi2wYDkjc6kl/BXM35z8FgSkCbje0DtXc9ocYS45qL1WQ
teMvHR3yVMwcqwHNr0TD5bS09i39Qr+Zi4Ncbzb6q6rgynZ3SehvzOnzr4d93H6l
pgfjiXwKWA8XyJt5voAw2qKNzvZVKPm94H0bTXwi7jFNckMam3paDlsy0OM/ckOC
mMOyNbgE7yfnNH4dl/0TQdJmoj8tNffaDdsB4l4wrtlart/+q6e7bku8RG9eQRiu
4q3asMWdoaB2WjfzwenkpQg5EFvPxuTz1VNI4mIGNxI2HrdEGO/QJake06OVL92Y
3etlV1FZYj1tvQvqoEyT/Jebw/GbFS5h4GjAOgOGsnO6XxwKYOzMNrejgkG9oKw0
rCJ/fc35Z8kgrtr7Bbv+EWwIdXBgxbJ2NmhvLkcHCrf+p8yeYLSpMur4evyhh0EP
En+q1wU1RovWC/4u+CNpzDDPU/+Ssd0hIlqBXdVI51Gn84DrmJT/IPNzTxmkM992
9Iee2amnjps9tfGvNDlextZXBjO9SjsB+jjXV9uYITUpFPU4Yf5xt4eiIpmv3sUE
ORbyK+fQRcn8jPVKtpwtZDJDKD4VTVavvwGD6DOGX03Pq2mFc2+0Z2I6l3Q1XYJ8
N1xP0dpknMgiFj3TW5K9HZr6xkkqVZUinsLp7IJpJaJvqwu55h0Rev3tRdal0TgQ
Z5etPpRExujeQdZeDOTWjYmayaLOfuKHbacqnncfA28kGWHfQv1wnfk+zk032IZn
IU3WYCM5VRuSmJ5E6AMSNKwUgu9rRccrt9HlXnvPkQNke0f6UIeoOhI5NGhuP42e
Nj2iIYs178wWvZL3q1QqbgDJB4W3TozUAYFzfGd8me+RsO+xOzTm0H6GTimXcFFw
Wr0xgQTUWzNEgFTicUfzvl77dnRw5ufPuzA49WeKY4OGiMBGMwVO7q2uAmogeFZm
6iDoSkvooMGI0AogJYI3Z/K5blhmnupc/TpZwmg5vUwPh0rpjSkqrgT8qVmosWnc
/RGaYiIOhsvpE96tM7uBdTRVwd9s11wqA9xJnV+HOqcldR8e0ABUHYHPXf17c/fU
TmGmiQzgiRHWDba0aqNjxkBR/U3j+6Ivkc0ohLt1QjWk75DZfGexp5d8KXpHfoAk
TEvalyYCUqzz77pUjYvL1tV0HCD0rOFzfUqLXTsqxfnqUDGoO3W0O25MKDHJakxq
JzxrMmN668zHTdvXLMAkSg3KXcDKo2M2mCb4XUqiReeFwfFKc3D1KKNMlDH5R5If
DEjxwQA2tw0H4tPJDoruDMERvPoUDq1el4pRVkldgmTAso89T7GUr1Y+S6QuKNU4
46oDUDnKTvyMqQuE+mWEC9wHSoWfQ8brhhzjucIqqh9qA6bGT2OdaFc41BciHgys
dzR5gWLaKYmdxTMtRt/aL6e5vlV/Lp/z1N9d6gouAdjhjXwzFZIm14DfQkQPLzut
Q16oP8m9nY9WY+kXIeo2IhKXBcsiz6uqEHlNL7DNwuatgUCOJ5oTjDxCrzuke8Ka
kG5XkxnSzcZ6k2ofYanE7BL5ujQEBIL9PBj6sV9DqIexnYERKw8geKXeGTp1JAUM
hw9ZGEoECCHbUP80JXDOl0rQA48idXf1s5JXzda4STlgGxSIzvx8kW9op4i1GLfY
KHZNhDpbcsXcXrKhSejJNFJ+NbjnrQTluflc7emwLdaguaxfhYSWOzymr4iZrovu
Io/mix6S6OXSAiT1s/58306y+GMo4sdRCTyChoYmzyqbCkH+7JZWcepWnLHH3gjF
/+/bpsjJJrYtP7ZXy+u9PiD4TCJgDA/eq3Om6BzyUW4puiz4GWyJHBzGVbR9g5Cx
BjgbvJaIXecef23GdJilCfyRo4zOk0cS3Hh4RnAwCedCUVNop/cYBAYkBO1Q20YV
Wn1iCtYZDob3l2BYRGzTKQ3sQKyGjsS+zMgZ/1mH5j2Ir2443vbsnOBBUMue2ckL
GmumzqaRdK81MCKOg40gSJmIIMJr8Giq0FAPdh9j0kw2DCPVPqC1ezwih48p+zFP
CbJeM4WQ/yMJl3V2C01EJ22PME2MgaQpk6IJJ9htuKykAEl0yq5AFO26VtKWxEBK
GfjZOLMiZGGbFO/iGT/FlmHkW3Ycnn8ZLoqHj0VOBEjXxaHK57K+PqPJJiVDrdXh
le43eoBoaHi0vQN4dQeuOllMMkEd+WP4b0E4QwSPhlXf3isjspjlLb3VP8SbMUhV
SggzmaZwDTzqSs05IehEBoSIqqvRkOfU9ogADXesilWKu/fWTG8kx7aMe2OGKMCM
Ejggstxzngp4zO+Bvq1nPgq5ZQWsILrgSyB66NVl8AlaSSq1Lj5sS34bvYPVPWuR
wUOuFTDk/C8AmreLNu/iV1mg2c3/edSEy72Cv7g2TYND6hWZcG+JzdMu81Whl6nV
aCNqPKjkXsbd0wdcCDwDRAF3oeaUOINs7tqwVxcBQ2YaQ8s5vS0C94WC7FB07qTQ
rx6W7Q7L5imP2bukq20G886AnnZSdtooIgmmeMc+dYMEG4jnvIegoQeBz3bBoiCz
AiE0RgaxvUvCP9/Bav/0T5F3eR8aZiAMpOwL0RocT9Dm2fCoi0RhYDyleaTd6gy9
CCOfl61IR0186C0tZj8gRgcW+HVbwkKCmMX6JNKWlUAGTOaBXh3B7JUKR4Gs45hn
H76gGfdEF/G+evpGy/Uy+GoCGd6CSF4mUn8nomSiR6SuEo7BPKuYJDe4A2LrAJYg
6xFPKIqc/0JNp/FUMB0G/W1tNqW63bzXxQ93cqKjivGoPK2LDFareOSDUQcYRzq9
iPtq9oc13CaP67JtBXvPDgXwRTx4WVZbHi5t7MyDIH8PiAeO15oibdwZpwEsavMt
Ys5faJpyIp90C9Re0BtjpVU3zko4I+6M0QXm0Wrwi+19AwYg4GZwG+z7tDVxNyeZ
exnzG9ZdnejjF1+vDmhJmJHOI24WPgSv/2S/UojGK2qnc3qsJ8JqSO8+1SP5w2nb
RkQDHNoaaZlmh8Q5iH+nkzHHVxo+yzF6hXKKq94cpSytvFmEgJI7n6poCa7k7/uC
W0uYr6aKoKAIGIzrpuOnq5x2RPB4AWUm+zzoyxw4ZaNkH+0Wly3hvbmQcb4oWmHH
HyGo8TakXGtvutZAk6snqITQS8cdGyoIiSUorQp/xtE9RFVAqkgPMHm/Yh8EU6MX
VoGKK1ZKVymV8flf2aItycIIzVbHzDMy68bigMpIN26/vBGXdE1QIv1FvJMRORI4
4w9dr3now5pKh5scaEyOvCZbagM1G1lF5xlZXT/2kN3PDDA6/1RTiEac6Z+wPTJ9
KyDFDx6GZF29xw0roYCn3Hc6WLoI1NsgGhBnYQn4ENCk/mdT525MELHtUtOe38JK
KNJH5Zw6Vt/MGy9PEwKIcQSAPQVc2UfQO1emLhVdjEagcjICJytbeE0P7qxCYstv
Tt0jQ2ampRF+6LgpnYf6SnsIcuZBZ3C3YA6ryyj6mk7dP8oiKiOCD6WrI+sw04Jt
RvTg8geUyUzQYIHcDbxNnB0wq+EtH+66CRKVQl0/rDgPJxv8PMKPWALckCggZCg7
UaQOeStLmmBXF/ooRh/98UNTUUjgGwJIUIo2DDrABSFTD1Z3zhRwVQOzD2uwWGov
Hv+vX7JE22h0dpIiaUkNkJyWICastCfWZn5WvOACjzZQwMRO1C8IbL0fo4eXQIea
BQOUkafHcr3s9fxSBgBAsQtIjzjlltU/0e4sjw8mlWS7xxgKIKL/6uhgkcOKGL9H
yYUjP/O56fRLdaWpUDdxUhWEiW/4WXyt790oj+aeyGuTb0Q58jKfQFssHNqPhz6o
6LHAshJRE39tblGVS20biPqVmXnQZcqFd7v65sSE+9+DQw4p0f0wVLWn9101Dz0G
4z7beZw4ALAuigV4xUfvIwFPJAschg9bwkXonyxgeHA3+hl2elOJCpeXhzVgT+rW
GUusCnvTnpuAun9zXidZNEn3WALJUpyygUoMP/lRaP3l8okKjyfL3JE6rrK931g4
bSZSkqOL7PuquenLp/F3mtPqN78WNB2kNcfEYFqjU5j1XmKneZL5Shs9oCIpF40X
BHPqdvhK7xLajZO6QVWLrkfnwgf3/xv85l85DhQjkDUa9W0rIj1tq5zyZ3DNm2S3
p3rniIBZ5i0usPNIv5iwOv3KQ9d5NYd0KhNBwjqbtFd8oX/6hNmuXcy2fdwoYpZc
ARH+OF1l+VHatee3y934Ao15DTt7AtiNWBLuX63gmdwDi0xlDBnqhHkWxnGbvSoW
0l6Y6CEeocrS0oTJ32xYTY8pmpAkNLFZUmhmCBS1R7DyOFNcJEDtXYTwBnUsxxk2
//cESu5BDftfyIogQ572T9PTUQGYPu5ITOtA2ThFS1+uPmxsLtdkQmDhaloZM6C4
6VjpWROk+dfvMTlvwzti5X4bnFBKaQPu/BJr+tGkscs/OU1W38/l6SlZDkvqhHVd
gQogCTO2AK2avhUj5k/9rJQl0aOpr4ND/+7BVe9/yysGWQMB1vu0r3VwRR60N6hg
4mh8gbaqpI4lR4Ep65C2vb3NRCx1hUba792aGRJ/HsYI1OOLaJcPvLBtl5ew1e6P
ZtS+Q9+Ng4te4lUWNXFh2sQWxxBer+66jdFRGeLqUQDxNhJLsU/xABy7j2nx38MA
+a7Szyn4tfSnwHOqchsBZolccvfqUXexnbzAgD5hcLbRv5cuJMWx7RlCqVozS/+n
j5vAy2AV9jtd/Ruh26tljNz9WTm+XVCo4evXFP5INuEW6MJ6KwwM8ly7N42nnbmq
LzcMEuI7pJOG62wblpY38eEhBrK18Xgj+lzmb7iitW6ErEai+0pwUH2v9JgqrEQ0
5nM9rHNiKFz3ythE4u7haE/ajojGSpZUjYacxwCSzyPub2B1jg0g4/x9WOy26EsJ
ct/F0qONRdCyDdzAqj/ZUEI+143piF9+UIMSMk0WxMXJd6+HUrs9/vTTSmm/I+TW
bMJiXfRZ+lXdRHUDJQqrEvKOmxd3zep+eZHFTC/J3uvCmQ3/zcRhfYo1FOyFhMMJ
CmlSJ55Ccx9m2rLQ4eSBIg1JdvfPD72foqzA4o14NUK8eUztQoGkdZZhHQvGmPs0
aPvh0bizPEAwkrcGHFooodH/0L9BgSvZzxKayYRkEJUv8XyAeIPK+H2QMMUdbl3X
QVlO/rRJXOM+dXId1LXk7coVGgsV4Sib9f5CULe6B/q6cSc1aEWmXqWn+6Cqrx5R
gZXngmYImNSfqwCi2W9g37upQfDnnr/u6wzLEd5NVSUrFCjTo07FfZWhlSqSd3ZY
v0PioO57vLjzFDBWtH4WepPikktJ4J7izpVSpfWXEdJYrFzZWOIh8moHNyQHFU4w
NbfMmIo3kW3HGg+LM06CKQSzjCO55z0mrSFUYEIvzM/UaXTiyr2eHhePs7i6EqJi
Ywb4yybOaRPy+bhCv/AeWAzsPr+2TdPLFkr8PyFI9x99XHhUV+H7WBqQgeFIXswO
zc9OAXBkDVZQk/DzuWlHHgaxBWcCHfFA1U9Ah74BQrGcOtTDRyOLDsqstI4mhUDY
b1d/REmwKr2aqfi3hRDMPT8SnfzaDjLthLkmy0GTCqE3DBuZXAfpRlBqctB88ibb
S+PKZGin1dWfyKnMwTsQFqssi80grk+RDdRZkM0HFHPd8RDWO2mzljpkTAAj8Vh8
LSg0cebo4Hjir3Xh12x5ZvhHeY+ItL0PR5rpQQmupkgVmh7F0X4bo1U/R5gBpttu
lIuKnKmUB/K/c0jx0AqCKkywx1Rt7SF1Lrke9V5XOs8leAKVdZUAl+MM0yctxKZC
gvWolYiQe38eKmH1zo3ayYRtqeuSKx4kBvcPg2hSyENJvm5C5QmJswTIPzC+Ce/6
ptr6eSxAAD7xQbaAuhn42Kdim8DWVSpKrF1U17IKnFk0J16aDvWL8sZsv3XBoRxt
x/wr3LwKQkqm8WsspBidAxaW9O0eR/sXoNVe1DW5ZDBzwidi03t/R+iekVFMQ/zi
cjjZD7xEkk/LIDobx0NWvy7ICbLK0bPye9Y/BBAls8FbfnET2uEsuRJIqRxrfdp8
vCJBG1Ndb7GibV6Cy43Tptszyx/WVobWSC9IeSBODtsKhgAuEGaelthQyUO7S4DC
n27qPkOOIx2fiswJkgl6frMSOeKFU8+w1GOLnvzpq56trrfASu/nHbuYpiWkH8Yd
wfEHSUo2n4isTT6y/I8tj1V3QQTtsMS7qJEcLRK15hReebQq8++PfHZ2owHE5tQn
HGZk9ONEa7jSpyVOrwBYhbTEIHKpdGx+alvxlwdDsbqBQcqXhc6GvbJZICX6nGwT
OH36OkogauZW0cZgB7Fz5/xod/6X1slXf3G+JGoPPTjUwIq0SPj2RtdX/z9B+a9m
YCBMZ2zMk8VQ37YvX2ZpXGWwlTrTc8hyRNocE4USd3lzS5ZWZYkKkyq2/vdRK08F
zrl8cMGX02uOpSjw789M/p9r0WvLK3ARpny1IW9Fi/33cljKBiHGGY26TZMc5ECr
onAmP0Q8ZXw/dd1TsqNaDXiy1gblWc8eArPJrm+P3XrupgxwzkDuI/huw2Dw44Nr
WZu0V5ZwCLcqvxUyIoybPLJKwIahn6th1VNAffDTKDJbQCbpDS5/d7kHBbeNTx+K
0U6hIhkc9PqL4TQvsPmry0ML6XLAdoNnOyoJTzc+WDyrwEA5J9N2Us/+R1R5jUUR
af1LDfjI+FPfKxtHhRmiUpz6RBblsOOR8cLnDOrtuKFih5a8bYkso71XcAJS7gVI
ADKavHRZZ4F0F9kO61QyCJukFLsvpIHc4wSNMZVIuGkM4gaf8O7DNdfQ+GoLXSiS
xIp6Lb2KGBNuWMzSLER72wdr/SMkpaPezL0y7rLNQiAgyXqlPrv59G3RmHGI8T8a
apBNYT1OOoDjTnEPTDYec2ueFMcExJByzQTfTgdbTDNgWceRa3YWuSUdk4iseYAt
yGzuWhyz1TqPQdTENRTtvHyJcYcQU00HQ/pYrGqIkAGVu0iFZ6lz1GPGt4OX3PVf
3nk/Zgj9PM4V+3GbJQDdWgt38nZJrHgGaEJ0HV/BLMXFHF6Tl0yaC8oLMw34/7vp
y9jJHDggQYOipEqBtkV3Ivwp3OeMy0cbAUYPN0sBSGF8UXidkICBQLNu84LfaXbZ
hcyt4ecJaIImPVgyWCC3s/YBjlVOplYn5mahDDIRiuNoXdyxPbgrGMHTL1R8DxbT
VHwd/oEPpM70g15/9p2xH3eAGf8qKeqQW5wjnDV5Xw4bnkz3vlFdVjrcrWC1GNdI
fQdHHUNH37so8kaoKIg+3M9bQ05GRYGa69vRWBiyItlvPrzG16xapZAQmr/+mA86
elJTHIwrfFN56cEIvh9j/+zpKBEhReFyR187LMUTAwAJNfaW1nY0Pqz87SjJF4pL
CNXtJVqUlgaXjw8s9SNU+ph9fAfCyVDIhwwMEBtnQIzIRB+amZcATq1Z/L3/jacq
r1wm7ga6lpv25qEuTVTBEi4MMcgrBMd90Nfhu59IOjiPGQYLXyWsxDiJe4iUU0XL
HUDsyuGWtlCXfjjdQloGq5NCz0mJzVk1fN/Vvc8kWMB0jzF62E7qapUDhLR/DzE0
+xZRZfYGjeTXymcnRm3ZYu0bUqsQBqb9qyfg+cupfAi7JGPin+o6w2RxTX3CarBL
qZNvcwBh6YQitINgky+KjeV306cARbLwyRCFKLQikprjJlqugvD8PZ8zSR7EApRK
EqUkigX01M+U+2lGM7l8fK681Iyv18s+fh8rpmnz+Rj/Z0rHS8VYfXuRmY7rwTT3
5Yy7GGmlfbrvCgyLJKc16zIlFPfj9GohxI9caYzKHy+FIAekzDwnhatOexl7m7T+
073QKEUduqeBpHRLmgKuoD1QTqPKsvDsvb5TsD5A7tqoRe4tE8sFJetOJhWyVpeu
agtbuBqnAl2i9aewrLxMEg9dFklOrcXkT+xszhiIunnX3cKbI4y6FcRpFxzvlGde
8VXqaYVgs1JqwZgFF2Sjy9st4LkyHY5tFZSFRgqypUyBEH2dd/MKera18GUnsrIz
jZbgWVFcCVVK3Uw0XqYMTfGDs3x9o0r+EK3eSaCTBTsLYeRIb7JC9pbM/YZMcdOB
BCgbgz1mh41LRngf+iUUhyiqnUBU6iSBu5+wWaFkA59TWqp+NopvN5b3kM7lVlsc
n2s5HnXszJLQuTiyiZLXcZLW4GRxt9kqSkN6qVM8l7eBW5avA5ITRynEsdsq4D+8
f8R2bdhvltdxDeAQOiDWHkyYpuceGBekKbuJC4T4i8+zEjdoHOQvuiuyUmC5eTYR
crDxB4ljZng+RebsjPkmG5zGJMUuCtxoWpi8gA2dAcbbrCHKP07pz6ECOUy29vRk
dN3eyzfSfHhgIjPByP0EoA3bRi8UcZa4N4Jb+8QE5fM1uTUwQJTDbeMyxJ/lDnDH
9CNSUe2fioNPIoh9gE5Iy3BXJKpa5SFyhREokJ2kVKF/V6zi8CgPXykUq2aROP3y
P7rGay18oKF89R0IINxFodBTu8/GLkj6dEeT1BDtvacUZKmp5twTSQdI/uU4Kct2
HdTKGHyCIcjuTD7NXVeSTHJefDeOx+qbv99YH7hIZgttgf+qeJQYapVihJsCFHMO
7FNqtEhuOeQkYpRlZKmT5szVW49ydXjBLHLmWHkysBaScw1QvRCa07eLWxzNL1BN
CaWkR2SNSZ02zcNW1gOG0JK5RJSlJBQB1K0RyZ3SPXVWkxPy8TvQjnyMMSq6zsPJ
LX1m4lwf2KObP1fNYKFXd7OTwTwr05Cpi0aRYAwnT8N/NvpjfNMpc7arxPZZnPMP
8Rr5PCBmgaIoCMEPG6EteiIFjmAEjE2t+2YiOeqGRxenr8Itiz05JULQjoO2wzVt
TWWo0Vr9wai2Pk3ki/bjVjnOxQ3TlI6ODfZ69ClpPYm86UXHto8KFyAO6cazr4nK
c12wWfHhPRYgM9h3Cw1rGtdPxLtQnCT2XXmhkS6hDeyP+kq2UWLZIFl+uAxbAEwd
b1ov1kynzPwwFc1LRuXfg0bqNd9rvH81PLECbG54W/FM1IEzeVHj0WJxWOyJJJZQ
4BZjgjZYv1aKyq+nQWCGGA8h48oo6Yg802PAGebJAbe6cf4CGoSEs3mrQYezGBiu
z3LKpyj37SO+17gudu7foP1vVE4MKr+5j8qLwSBThVfYJCV5pW9WeLLOLUuKd+PY
3bx0Uz7BnIq9jWaKIWUHQ6T4i64VmyRCJUhu8a22w+gPOtbSRwL04u9pdJdRocVc
zHL4P3nDZPCs36/EQHdeP4upRkIQW/I3GGhhnysjG3OEAF3SH5ChCfvODJh1I2k0
4ZL0YJBRjw4ck83cEDxVdDEuHH4C7PVKRz6W2bd8x5gNXUlk+q+SEh7tEy+MsIgS
OGIKvOKLK5aUY2rM3u5heLB2G/KbdhbboCKT9HyplMoy5RiAJrXq7RR6WVZymj5T
FdiHAWW5o7iQEGl2uQSDzUqK0et+aa1wELU3MTpNT/+iIX/7xrzqJVC+IJ4tGVDM
dg8kG1rWxAcV/YLdWVXeil3irqH29KqurML6YsX9KPBtm0e4tsYHT1pv76FLHOuv
IFwj91FzIfwIWZTR2Elj8x2SI/5XtH0ve3mQWhMlP99Whn0BNtab85dMIQaPaRGA
k1TjPedZ82ua20d49tsbTpK4PXJ4NN6Eswl+ot0NTdQnLZpDfGSaS+QF2+CqFh7d
vCGZ5QEecq+wuaJ0fyEycpS+lrhz4Zt/2QHNc8bZRw2qKBE3yP+QaPwaeqI+LJBd
zCvQWGR18K/gTif+OiGT1jN8PrwgxsFtfAjyykRml9zTA83NDz5k7ocXn35YcW6o
N05pzuBeB+vsmKca4gasDrDNWrTbQIFsmIkd2+S1WXlwQQXxljVO2uR2f6woCphV
Yt7UEr/0GyoOGjxm1985GEUErhYPPPdp310KtIqVCsWtc71HTWtw0T9q6Z19C+Yu
TUzmGyXEddjkuVT05AfeHMADAoRYxb8ehPbfA1TqXnkXcOmTPPjVtM5isgewbo66
oM1dFUM+phz5r81auc0trJF7EAooJPKUWcOZ4qGjsC3vJSsbgEzhAdcbqjSGW1nN
Kq0oFaz1w1EBPiaWaf3VBDPIcQqCP7QUsdMcGgxJgEpJH849uomPmEtAR7eLSSY0
6bAj6zjgphRAmTrSMtTnSyAXFe5O9x0I5K1Ejl1Z80j3UknC/w5TBG25jor8NYfM
5nqkyJLdjGHv8dCwwOa0hrXyJzfVPxy+Xgh/8CRHZ/yzrzxr5S2x5dVxZf9CKDK4
ZQ5YtGSdXSV5MMLwRYx9hl1MiQsC2M0+Ym417/zSjjkOQlYfVSEpcVz1NKxUZHM2
nbs8OCvpBTMinTFMHcQPizXQhxA0/OZpD9eDINV2j1L8TwYA5naQvrBbn9QGAEn5
OEWpjKdvGtbbRaWBMCYGY8tqcuc2g3aTxUTxUIYi4RdivNNWXbO83/G6Pr9BZI4m
dxGTiikzxXQFe/pdUw8f1gqKhytVVlu9vlvho3WBfmtgwUAY+s5fG+JOt9UeuLUi
oNJnxHA7Wuar7w9pUMTdMVzwiHHnOGbAgUZyb0LAB4lNKub4POxlL1dLybSFvD61
o2nMPtgYGpCGDfy+h6Pi4ifH8Jd9FziuGKGP1vQLzmFC3EbxVJzpYsF7/rSV/9e3
OL1LdxcCsJ4CnmZ1++TtwtYDLSzDI/bqOBVxA6ojDReVKV6QkmaY4y/I44TLhLs2
OLdIH5QoWuHra6QIjs0AUD5o+FdJO/wH+g4CgRmeA3X2nZKLjFPggsFtf+Ic/6ik
XxVyQlM/Dd1f/5EonPJU/hpHB+wr2t/BhrAJgOcxPyq58WKDHjBG3HVJf5zZYgTj
omhMDPJ9If6gRGrFuUpVlpz09XjD3BQHbqaNsY/D/EKg5PuW9Sz1Er5zYVbvW2BR
1jriiDwDFqp2/Eo40qqC8BBm3u9YC1MNZNpJiVMjhu+MGfPMcmP747O8F9Tb2TMG
1E/hoU8iFWmXCLU0MABOe3603pz/rRwHoePrby3AOOduRlJt8LZm8lIjr8bmoQNk
DlyH94NTfFjr9+QOTSpMp0aTfVsTJcGSc6RBcb9TqoaX2zOqJkIUm5sWpWhO0Di9
UCO0+Wjcj/jl840XUYo2fljOJBYNxsqeXw+XeY6pMG7c4T4brV/9sVPuN+G+WM3X
QhwhaeqCVkNPg6uzSp0R+FIkaInyMkmD+TVyCovRNxZY3S3GYHHmWFCigJPcts5z
ARuq9Bf5CGCpc4hGkAL3OuhKTCTyBB4eQts4cqY3PaknOJE/cpGp66O+DWXwn4hp
w/IGzOo+iLYyAgweAqXzZM2626O4aQ6wuMYrBbaLzRUuXFIRt6RCwddFMaSAwXiN
9UGGj5pMT7VZK4c4tUcMqTIMJdpGO23Ys3UK5NJiVddl4bLgixUfhI7gkk8L10Pq
Z0Ayr7zPufqLSrA2ni6kjNuU/spKj+JCxaQmxFedGocPGsPprKxJGDFnExdeJKPr
De727wQiS5RTAFaz0luM91+OqlgI7UpBm/ALaWtNCsFKmk8Kovwx1P9bsPzVowhc
4T6PDdf3f5PgWqU0bjMfJumfBAY5xvksHhIZKVh5pAit8q9joWWWNasE9o4qsPfk
CnrOUOO+wXBd/+FRRy4NrYR63IgPJCY206+M0OdbbN4eYUl1HWGU/F6L4xq8mp8F
wVHbTuVfR4ItlS1CYMx+Y1bYcYCSQZmQWG1b+BbJ5/2rm3WpdLh9gVEeTwVMKn4v
lU7QFyjJXFlvT+ITMchXYrhmc8V1IfwT6DK7OFLsknID8G9EUEC+D8RpSHZ+zfnz
GOgdJvspqV1RoX2awx2XJN15l3kfEzy2sn31EYutcW3zvqWzrcGtES1uUoZOvrkW
RjR4eDH+RddcNF0gnCGI7a5y4iVi1mDpg2MTsiv4RtQ0ztuV7ogi+aC0BQIKwQ+m
XIZ/WEHHxYDHUjcSs5d/6kIKgyfGSu3ygk12P+WwayKMCobSms+fpjSxmV0/A338
2HVric46HVfXVQXIW/I3NMnM1UwjgMEIZAcCAFCQtXNg01Zw+yD9kczApmPj7fOD
yMVpDWmM+07HB1gHpfdvN2dzJ93P4B3N9zjvB7gfPc8QybKKDVWX+t3qckJLHdZ/
RfDy4wYL1I/3ZW0qrMg1mkYP0zslIuIk2KNnWJKRZBKjW3jUY8uEvsfGy2wEehIb
7dA08Qg1j0xiGqLqUtvIoy3+HAylewrFXzZXXG4ysnqv+fZ895aSzRShBOxXsreU
V9xpPB7HEIspSOP16iViglQ9CuqUt6V/IhNrTYn8fxwDu485/7ZbyXCIOE5q+DQv
ZpSMFX2YKFIwur1iT9sLDNyDv1jdDP8uAcfemq49SezBnVCVWxr9w1281eVPzefr
KBML2BvFKPrcrzDXAkfiOQiO3UAAOX78ExO5K4SOFr2Hftm0978GIjZrcFB9TcGG
jKqYAJmIJis5fbpvFl9Z4AWBp3JtfJOLAZANDwm+1TCPUwPuH94bDJQ5xgQrnJja
evTiNgYq/uTndEWKGbrSfFozcXA8hwCniyilTPmyJgijDRomUlvPzYB6AMC1Nv+F
IBE+0MIiPslwSm7n7w/ychrfih0uCFGy5nAe4ebNk4Z1DEEwFIPtl8wj3O/I/PmB
WXO1FnsWp77yNmKevsV66lhHILcK4fosF6JdJjlUwf5Aqym6mzuQJuWOKt2+76g3
fX5IYtxHpMD9/yjOfYMoiFJQH+LoSYnxvH3PWKKLFOY8cF+xH4V+z2E1LNfLAT/6
dG9pw0sOC1vViWDmrspjlcjLN6rd2PDRNoYeLptXoDID2kRF3Kp69SjryOUHru0/
qJp9wgSH4dHMdOEp2YYWjikTr1OltP17/zo1XghzfzTy0pfwsJcyNqiMEwyJl56P
8xbeD6ZzRBpK1D0ta056gOfnwQvRJvOtj1vzqQcQu2zH5OTferb8I5LIkIC0xbhP
cqS4d+WE5yfrl9L4RjWC0nZdf//SunWnRtKIehIZeeW1fI0Yo1vtDkAldBipcVp6
T5GflhCMGKBlfYLlSEfh1JHZv4zNU/UM2hPEwXVyzEBooWvaCKJM5roZShhA/JDH
iERKh1i9EhLvmKKp+ifVPZkr7rslBHe+BHvU4ODWjXpLlz3z8ZVdu/FnT1XiKmQU
50gSBzLh13E8vYcFSVgF1JKtB5jE6U+XiXIv5+TapDWjsMgG5spO7yO1XQ8V6Xd1
EMyo9tV3vQE+J8xE+KHqabQNi+KfNNVplg+akvtxadS5aCE2DeOgEz9frMtKF3w6
Mj6D5T76pQxTu1DgNETJ8N6FMmH+hJ/6mhjsyJnUcJYf76zt+NZtRDe/F+kyvLZ6
V9pkdXEfgeCd/hId4iKRYEzQ/DDZ93m6ECLBUCJMiECo5Hx1J/QChWkBgPATjRg/
4pS4pcgdagNS/t1xcy0G+EbptFwj3iG0vb13iN5zC6Wj/EiY/v6rs4ceijPU7qBh
R3XW0fJR4L7s5/69FZ6pMOcSMgnYQ1ndCLU0m5XjIwe0BUWBKkoorqBnOIyDEorY
/2BF0ALZUNwyHUnFIEzOsiqZVktugHAzoXOQ5HbySbPnQTRCQ0n0n++NJsDknfBH
auI8sdkIMNpSJWOSeP9mFV2nv55Uwe0FM51uj3sqNuNeFN9aUt48YUnieNoHlR4f
tD6B3TcW9v4ykR1q+JAqk2LXlwdL/WsJ+tX3pCc5yrPaTUzP3Twz5QOPtREjNx/5
x//iW8TveJ+KsK15Hn9Nr38bvLlvXXtTiY7dOQI9xq6bYlRH2VWL5mBuzQELD1ej
UNxKiXlT2qrcOP8C4f0hwSabeFXIn0DRL0M9dDQ6dUHYo9xmTWyqxkA+5hZUj5C0
NVWj0dFQmyfhryfQfV94TG3kGI1quIE6CGl7/MEAV+mVk6F4OqnQKEWripWzCSMz
Gt+2wvpmFcPqegFMEW05heoYqJf+tHFO/XLkSKfzC2AWIiRJw61zE5x7U1SvK/kX
TeKIuYUkwPGD1lv1q2s2AQT1avqR7pZu+dbItK3zoRg4jxuI3opIdNRUeOuhpiIW
dLNOAafc0gS1tQzlB58/Wrp0D/gCfn7DaFv7s/TDSjQR31yF+SC+DWHhk+nfF8Hc
V8l/Yn4Bq9RH2TqC0BXFFGWdIazvvcPXoapWR59SGH44w064RDUxx+8Ap76skjfm
rRQ8EIDUGPUQIILgOEkdqUGI1+0RjjrGmljsiv5Gwu3QME5GNAWculhBiXzR9v1v
TKMDmr3uzYfuJ/jh8MbWifkGU5LbNOIv36b/V0C3EIARzssZmbtfN7+qUyPBlTf6
FhEmbj4KLgss+3rK7klgWouE3iZ24IDmP/76H1lHsSUDfAabQIiXRVAk9slqDIO6
iA92hB6G9tuxj2uqjk8PlXNpzzwRKPHsBFWx/VanpMYK+UlZFEtOJvGKa5XIslmO
cmDE4pzJ4082hOpKuUA4m1eNz4GIp96knQLIm7y19RXOn1MjK79mhDbV+B3qFPZ9
aeG4P4cyoqWsFGk0MzGtfauBwlVSfEElLkDC693wEadEEarmTYD/OeQdHhyOfuDG
24I5r0Q6tzZsBBSqy8I9mUeK9YJ15QXKYNuODFJhK+iHybl91upIdFUVuSQ1ebvO
qTmFepn6dOjT7lr2OQLAoViqScfbx4ZaSgUcP+85PzHi3KBqNk5UfHthg77MFWRq
9vJe91ICi6x0g0mIsF2eAROFSNF1fF+MFzVuDp9OnoTPu5dIkWKP3nPxYFjD70KB
NsRi7G/i0AYLXYADskMh+vSg9D8r2SYyJzsyAz7f5wYbmSI2liYIzj7iVF1vQ1Yv
87EHAw9FpF6//dHGvKZOXBev4tpQEnZzWgJYU+JxszryVajhFCqKxfK9PW77e1jR
AcC2sFl0BipVRQAt5Rsi6hPSVmmduAjtyKie804KDcHaKxXjna0DG7oXicZOiYMl
tqdh7f0o+4yTUpNanQDr0S/mtvPbMLzVurruCLVz7YsOz8CuIy1ByYiJS4NJm7RY
1y7umDcNwHvrt23tK1uLMS5Ic/w/+OlbXQvjbBVpq5ospgowhx5VugnKA6EYzsul
M/gzg1faOPJZnbq0dLRgfA8eF3ejVZbRlTKpMmF90INOTY5U9JNoTBCvt/snj8JX
OWFiuEP0txvgFwrIE5CQx1ztvyN4J0/XKPR7cUZv5eS5z3CPHyvrhS5af/4LBGYV
QHAkS2mhuQrxWN8OFi4EqbwdCawEayCoX0eyF1g1B8xbxTZctX5MeJnXFtIfI0K3
Ly4Z/Gwohn+aF3Cws814RCY4RHPaqr6StKtW9+oP0UW7m0O0uzOG0apX1e6/Gh5i
kk9AjXmLFhMzcxJ3NMPQRRlmQOtgX+tbhmzKXyE2+f26W/kPBcNqZ+dt2qFJb345
BC8h9e/o69/E+BjiTw0v6/ZrDEA6/L0nii/0TS7M3HT2fuKCz9dkjsULgvKDHET9
9ZYlrL8DPDQ1/Axv+7AqmzO2gc+vD199ZLZ1FV1JeTqyVzQepOlVVWoE/P5bFtSg
BnOrKmdfOQGn9uamlxkcpPsWYsBpAYrev2gYYOejU5LbDJmeUdCmaouLr6cCSkAQ
IPhb8+mBqLz0A95jMfNBZCOpjZYVE8ZWy5Od8tH1C2b/b7ajEA1fBmcfNgA4NVJ7
g0czyIkyTs8cv45655YU1FnJ9rthltZGaPa2f/cE+qEykoZ2VhZLGoaNUo1wuaDr
TenazyHZfFAlDaruRacdlSx3ywOvxREyabfB+TdXxx5oI5QxVEk2WKwIBktnJU8d
bf4Wrnrs5ahDb1FxacJWgLlKlxqF6Yc/xakDZetRyqMAireG5TiYhBDqqV5wTUMZ
/ZQar9/6fLCOhl3ju32z+/0kzzY5DswKDSDGh9xc7VKA+zllW3NrIe0xU4mFtSv3
A690qY5HD4Wci0xVrMWLUuN5eJOcyJsfJmEd1X9BD2qwg/6nK//ylfp3hgqzLnp4
ns3JoEfAvkRNtRKRpUnxx7BtBStntDc/Mvr8H8YUrcBCIs+pC35GTxZMveoY3ni0
Ll90mDnZdL5GD1L5xmvWEAcQMx7yIQwL9czUeKxN/hfUUXZe8OFYSZFCDXFCj/tV
cKXhuV30x1kIz7bGfMj2/Z1fj3cid09kjpo40BrSX1GBEEt389ibtpix40VhJhQ8
51rJNFP+0satoqQ2tugyWdkYyiv//0M00Yyo1Ww/GChtEMRE6WubOY8aCdMBh6lE
TRZXFYr2CPIlalm9t3QE5bhLE8z8m2ozFJOMWht16curRuFGDl599TeJp5DlVrY4
1KDZdyavWiz3ogaZteqgXY8cr736UYCEhqB6Ti3XPwtYTxzI3u7osOF5nN1cSKi2
xpZffrpfy4+JyQrc0vAz+2cQ1R4O2jNPiZP4np7SrVw7czCMqkihj1IBs6UeCksJ
+Nx19KVc9p4JLpTJA1/TmRlnbDdpmIE7CppyF3naxOa19efqcG1vspapI7KZXrgk
+vTIMYsLVgH8EIqwLGxSXYllZV451ZFE+SfQCSV6VhKyqASW0f4ms/WNqC01FIOw
LFNJRSDZFO2pokPOsazOF/Lxlgk9vG6vDQ87NKJIaCMxnXraQ6RMy89HCYIxiLCk
CIulACE6LdBuSTpFC7Suy8hrAKYdDx4aR/0qwpFr8I3sv0n64eKhSg9JIsTyb9Ze
3gV58KqDpYR01QB8+1VYIWSTYT52KIJjAThUO4AnSnf5ol5EDrnyF3GEQJEF4Kwx
Y98Kn0HbiWWVLAwGkKHhA+xdup+TWoSCBVTzDIkswOQqjqQSKqRVOvn4VJAAwri/
H3v7sCv0ML9uL+DQUwq/HpCOWUT9N8H3iQwaAdmL2xV5XJBTPTgJj4nGKU1jtYO5
OeN1v6cyFNK41maHKIKGMICW5RKERFFvYPSjD/Kdihw1yCwMiz+1dr+rodEeDwV6
0vzAhwkYq4y1SbQGDeFZgv1JrYaZCNl2M9KEtjCXf76aIUbz3oE1LBkxv5TPdB5H
vyRio2KZyxh+geUkMbalX7s074J5G6wxD4wIcGGmrn3z9CkebPqFmOB3PUEhQ8zh
cT/BeuyZSmyjN5cFtcLluzM78UnZsMtmR5LIX88ordGfG7KDXlZV1d7Yh7Bocto7
u7zwiH9Ygi0BT0nHq/it5Td1Laqzl0xu7sf8I99ayiGLMeCnxvWibwtLQ2Lr6q0a
3tb4bw5QtGaOdIUvT5nka0+twTVaBdHfIFPTsvV/a+RwFN+D2GI7/Asnk5mqH+p4
R0DpBp7HQLvlE9Rl0RPwXS8yfkTPJ4F5QvkKaTp1UhmnE+jr+m3e0+JlbGGt3b1U
icV+VkyGmpgSvZ1k4PU9crUnakpmOlkL7dMOq86cNqMhDArxNs50SM0VNtrX3BkZ
vvW/QKGw6pi9RdXXOhjld2EcjldjXsPmb8U3t/UpGxA9HOglDrbs5pR6OtLYFa7D
TD5Y9LWe9pjVby+kTBvCHy+XuneO81pBL52R0zSY31/1E5PCUyuwXrR6smRHPbha
wyKEKSlX7HncFoYAgxtX235M0G+RgLtCARN5BTBpUSl5vX02jsRwurHvQlSPal/X
9RzqWCRGXEy8Tp6fRMg0IsHEE0d/peD/doGybabVrGGulTg2ZdIZkEes+ZD9vlGq
TqZdHchPxxlbFmCLjoSf4Iqx0auGcyPE47l+KMOwVw89NC7uWbd/H9YO/W/cXk8P
02r187WEwF9RSJwodrrgD5T0M8QCUndUHiq7bu07IqSOrnNk3eUdFQ2AkAffR6S/
nKpUbcEpLINQyry2DdCb6qiMGNSRadkoCRB6C0MxVn4/wnQvQwdF8eOSATJAxnt5
KoCG1BOlQv3sDJdq1017JaofpqJsq0rcYf9D3c//y8N8vYrzEzaleAo4H6Iz/7gq
nW7mk0wIT28Zd5BGQvvsfOeSDNtKQwDsBUJo+jy6arbY1RsGz3XYexD+Fxjhxki4
gF/DuCvn4p2KaUiCeQn+a4h8hGXHzQaebfDyWrvc+pWGeozKX1K/F3gp2QkOlpDX
GWm5j/szKXC1vqSYhKCLW4xwRc3blYh5uaVDzPEYIbN+CgHEB2kEmf0+0r1xDX66
2YFR0niDcK2Hivn+ih7bMCLV1W+Hrzk6wSSa3O4RKm2Gb6iP9F8Oy+OCBmnKRtZY
s0UUHwvL/LQ+rxj1w3mmgG2+YvOs6TnKZKpnwZONaqwOlbFltjTLa3eMzD3S3WRH
gCGfVy3G6H+DCPZJ8enWcawc3IY3oZUkNSFcw5Hom48qKLxF9zoFebnyKwFJ0xUS
QPE44LvsZUCmUFBAwHDLExYHxjvxm0OZC3AITx2BUYOOCGTtPGFcKXY8Sx/JOx7e
s9S3j1j80CJk9unq3S98tg3zegSykDFquwXVcWqCxICE4TrvQaaB1eRVq+iJbifl
7hlzA9WaXrysNBgGrrbG1j5Y8wArZNFDcfsQ7poMPd2zNub3N8+jcQTWSu+/7Xlc
DdJqHDAvX+2UY6LEdut6tgazC6ajGRoGV9yllkJkwPz7y9ygQgTor2p2LiCdTzeO
ZXACX3dl5hFQ8l858wdlPBhW3PbRuhSi4jNf6h0rwCLZFZp4SHZxVSIZU6I6MCOL
6vG57mANaTV2otvkhUryPi9N8DggZPqD/gxwIfbCppSZRfeO3I7rYzNcjaS0te4g
kWNCg7mby5McNtCO2dPE9edGVlOrL+lx1vCZvoSgqMrDGIhcG/tDd2ukB9s7xpMJ
cLbjuIjTvxeZgKxRViFSl86trhbwYv3zhXv6gNiBr/YwDUwQ+79GH8SgtT0ysNOh
56bMqOTV26IfVoW9RE2EnZmFfQigTcOheXm90m2zkqkaJypKbRxjiuVpJ+aV/PTF
ElMDSZU40Qfca08XcefYgA1uAVhCDTtZzl1L7q+IHWD672lwNCEFl/qP0WFCGYkd
zyTyaCUX5c8X/46iNL+H/7i/uEsw51UoH3d+a2jOyWcfD22IDt1+jIsBQz1U26E6
QBIAh64pPdQwYlFrXCo0ZhWz4d5ig8gojNrjreqIqR3NA8U7fQnNpUE05cyIUdMe
N5U0fgflX/KS84wIipcV6u27CLxznfehDZUZoaM6oEwz9QrI/TE87JY0+MXHqMGX
w5TrK64vIwejaSY4vm0f9pR49WDHfp1hQEWKI6OpYQD6xwde1oQDi+B68eTAdodf
loM1QhU4/VJKD+cDgdmV/bEJHwG2IuZrfUmUuQH4sZ+G4yahzNpuGpwlKfERifgB
yDUBbN+2wcD5JtJyENP0BXhw+avdjXwEVFlmOJQ3ndEJhfroNgsy1SteJ7XnMGws
5YHzt5Mcuu0OWaeq0O+OTZPHW7cfQPJ2aDJC2Jz0OybAEvyo65NVt9c+JNb4jzDe
Qj1QC8FnrXJlsjhdD9T0+10If2+4BLzl479gEoVfJo58sxoDRSIcu1rCGY4tSMrg
ykAW7RRotkEWlZa3G4+IXt+hPJ/ZQIcfWpZk+jjkOyBNjQ6AOsS/xOWBIT9VElqZ
ffZBGzS0sCFoBA/eLHe055br0rNHHG/l2riSJ1BXDBQ/Qx5p+EiiCJ7JeFtT3nhX
BzxnyiLfpSe+sM/0RLKmLHJ77VG1MkJNWQX+c8FcchB88mk2qNREWlb70HjqHOZW
mH+gemL7ooC8QNDKzQhZyWq8OdzAiXubThL8Ml45acqzp3/t3ajIvaZYwS7bcU+p
5YTieS6J2TqXPPYmrc5EgeeG6cyomRwl1oi7SiDNB4+Gn8JkNNCPuzYFFiUlFLqL
BNlGTKMDkb+ciOuv9cFFgKgmvyX3fOXVZ3TsXtxdKhwZWR5/naypMt/JUuy0NfWf
cSOJzwyikEnqhEg6eA1qkg3bFiJ2WTXUYo7LG3xuRfzOatWVem+stpCyF60P9koH
qsPyWTCNgMu4aQjKIwAVIrKcwjBpTb58ZPx6+T4AbrvG1ZVVCCNnjEeqXCeF1Isa
oNRY0Ru/1SONEvYyAeLNJFzFEBpwXVEX3uQzhCqyFCC72RfSn8Sm6dYd3tPKxdJE
pYQAx796zbYTBVcL+C/5gL1Vfo4LismC5oxx+HPT2kUnOqImadeAGryJNC4xhdme
D/irlTLMB8VcwDMPZIZiirxlUaV9kIvH7VzpzlDevxu9MIyKV2x2kzzY6UJg/1sB
9JG1+wv+C5V49GRargxwOSya1cxg30ufDGnz/ScD6nwlQcUGR1yG11EwshyxfGwK
/+iVl18V3LZgSoB3SaP6vvUvGjvo02rWldf5G/MBpcLSCwV6Zr6uxRsDPSZXO/3t
UErRXR3ZM6F8HRGQTsD8Ag/zgvxFI3NlZdresXwgE/X4ZXG0w9obX9KVWGgMBvgd
Vz7Q2iBNRMiNZ4rf7der3VPFoJidtWywIE2pCTaL87hXCzHGas5U8Nw0qM7jz7Md
l5m+n0FWSON4Iw2EALUdRGUuMKe+SLnj6bd6GYdmBMvMI0kn3WIzEvy5bBARBGjs
xSp5mX7QB6OT5dcdvgi+iht3oSy/bZZ29XFsSehb41sxoKW682AFje/QXHikUgW9
HnBWhsfDLyii21uh7UIpUY9p52M3skFjvNs/rXsVVkHYVqDPbuL1wP60U0yMTQf2
RmiT+Jdd5+c6UKcvFVsxfktRLmMpggW9gGVPbpK06z30RKNub29yQ870N8XQP3Tk
HTGzOzQ9oHbeIo+MdaZg0Jr3C5WS4Qu8Xx9dMDS65+yQIZGPYB0sbKQSVqXBXgND
BDGYQmyZumDP5CDAKyEoiAAy0LDfQfNbuocYWuzkeNTGqPggaeGegieZ1TINRf+n
6npe7dxZxGq8oR6XpYlHy9vV9wbsjqtAFXaqiyReCxoA27S7dNU6kCVdTlJeYX/d
md7JP6XQPv7rIdTuUDfVn1jX+bOYXDhxeYisV+vEy6/VHMohzNfEOlDuuNKs0INE
qcDXmO1tvwDDI4BoQskxfAvG1YaVli6FjUXQyu8d4ELPcz0MWIF8hsABS5+8i6M/
X96vU5CmjoexMsbhi7HOlyn+U5BQsWpFyNtf7uf4r6P2+peKRaDUX+DUER+2dICg
1i9RbzZjLSa/LnMfuyX1pCTlBw5UqDLKrfZmjQhRSK14ms08wYZ+wMz+Fl32kfvE
JRf7XOABBQcsqalmgm3sdVHlm9MZ3Kre0yWCaLk5jBoceGytNpWRGHHdTPWPd8Fn
BT8FA6UiiJVTg7OUtwH3buzuD6JPyzsJUX/JrB70/dTZ+VIJ5t+2PznWTl/AK6E5
ANBprd+TIHA7gl0utw2dv7iJRFQ9nGHEcf6k8+82S5lpdZCjcB4t0O5/g0omDQpc
oNB+Mfz2aqAp8SBtqy8r+1rs+ZyR8yfpfvf+ETeOI/kFDZV2Ii5Vka0dvHIqPTWo
czy/8/pkk8SyQvXzF7gcwlcCZa7IvQLDl9hmz2+juQH0+NGOPJfBz23L5gbOdIe1
J4uJio9Y2SWfUioMKAHTFcjDJmiZ1X9Ni0dUVwykCwYOePMcDrKQWdv6IOVhFFxD
JnGXnuvoTnoHJgb6UTqrSKZwpXQazYR4+gwqLR16i9xTo4ZzGQAIDXtw1We/EM4R
f+rRKRTU0g6I4wY2nZ3hB/r9hVGij23qU/wlZxQW9uooQg43ZaJu2vGIjpC5Auhk
RscAcc4EHrWdOwYm94g5JYxSeS7it1RES1ltdBNoouoirkxeUSQGs148/d/1zk4Z
pcZWfVto9uP1MmwZSVRkGna2bmNcObLN6tK1RRaoSOBPUiTLlYN8UtChQfYJOgVX
S6l0U2ftKBqkZgu7dhGp5hFkHG8PeKDFlZWb3KnVDa1lve1/XLpljnFCbTIBHXHQ
MFJ/FiYva5skgDyh80WXk4VGlROd3CyG0sge6ay7pQ4hVb6f3sTQA5wlEL8m2s4S
bD2LHjFpg7x/06ofwjhqX6nGtq4DwW3UWtWw7AQreHTDIPawwEWzZ+5nGV2DSj40
mNXAwQMae2nSi7DAZCtuJjMV2ne0xfW82cmaHl7qZSp4RFNxUURuIPgsB8v3MloW
lDOe0sRjD9nasteP49/E1f3K3ya+JIanb94dWSteJ2cxZFE4BPuOlEEkFO7DhnHy
o7sFwJQGZ7lGn5D7HdCHKV0YL9ILl7vsEV1rBF/oKjxhIWQw9T5xe3BDXu/fBaSy
PMkKb9KMe+1IN+crGD1SEtKgN3O21hBVc7PuiRmMZNyoiCNPc8SU26D1zIcP9Xmd
ZODocfeyzSWYtpACZ9gMZFVCktngSxjV5G4l663Y69JHJ914zpxYVKBe7SDvZ1Fx
5xSs1lJNN5i1yKLKLSflVhB1OvkXXyF7OjjNGkBDLFvl8LLSCsxPrEYNMTSTaxKx
yuTRIt01lQrVwg6LKqqm5lb7NzAwlaT2ry2QotgAflA5N9NlBrckby0E9t+6EmRI
SbUQBEwvsWlg0/pvSd4KZ9b/nW1QCdE47IZTT8/q8Dmhzuyi2h5lXZtY6l5ulMrQ
ClqtxbFIj3vw7PJDw6/4krrRBwXzjq1qNZHVSr4z1TZySCC7iEI5gXmQV2qRn41n
w43SIyKN7juwgWnaZYR33Jql1iZXZoreyu5eIvBzIpL+4ABm113pZk3H3KHbYcty
mifj9cfD1gbUEvOrv0YFI7ZptiU16cSCgU9HGQtO3xWmG5d6wbdDVsKatUCuCgjV
ONVFa8F1MgB1lsKolYq70mwW8vqwZ0SfJVZ1a/J36xfDtYyoUVCZ2cns39lhsqYf
5wEH52UvGKELmVRqzzd2tPjViiAkyWTDq8FtCF20ycdX1mqFRcYJywtMdlzPmE7x
3trHd5HMxJEJPHy+4wuGvaBNSR00kg7PqovYeLpHgOvI60TN8zH3jSctrepHJl3t
pAf3lNxTumti2ZlFlmN8awp1CcDyyeFYVcjNJUah4na+nTDTjJgTWitK8cosEFQF
C4W9v95BPLJ6gdAAIvvMNtAkyhaPiieMxaG7XZtpjrffWta7EO15pdP8m7uYvAK1
LLqwZb58xbORPQ36tVfDTFETccqF6RMtNX+1FXkR/YIlmN2fCMpo3HRdqgARJ2kt
GxeAo8nGepkOEPqJ2HNw3Pus4WwMc1Cw3dcAODUYok6vrYsOf2akL2G6zV9nowpI
D5nFd5kGwEl8rKjeuJV1Hfcjcr5ofFclMm4iRtiB1MlSobQ+n/nC2bCLVpy51Shm
HIf+39rjZ21i+Kg6AXfzZHnpEZvklI+dEhOajRnojOEJGAYW+pILTf2h3NAms5fR
MvtaoPz1bPaG/LcksXZQ606UC6tN3VzPE5HBFXTrBXHFVzCEAYjp76FNr18C5tGa
AE9votEVH2C/GwET1ltS3Y8Vv43/iWYYgnTanIhjDolnYYjTGMwUZZU8A12Cuv2X
V9BvvM0mqxt8W8PC8DLTqcxcP8IHkPB86DIgA3gVDloNy2oW3/g+yAlBcSJUJ0Ia
xfizZQic8TXsr6v/Bm/pKE4n884dVN+CmnQYY7E3yiPCgqTz1eJQlZ8tUrVSHAYS
/655yLvZmK4vBuA1gdbDRosP/harK/7GGroq+JMDQGTGROntAgu9NcwIkMGeCgTT
YCzqzR2XUar0OUV87EFO2p1Xgt4lCQPAwh9KlFwNcIZS1NLHmVUVtOxYgRN0Bzuc
cWVxEv8wvHPJoWx57aPs5gw8day13cr1MLy6Fd6BvktAX2RvsiRrPsTWkXszZ/tB
54WEW+BpIjwsnkk3kkJNyP79l10kok2ni/F2ZfT0zcKt7Lz0YWUFr9Ntv4hohuO4
06Ty6jpFXO4w1LzS7eCZsfrbuO/uaicjAoB2fZXUWp6AtjL7/apkOtIhDRVKnP3V
q1MBt4oNsRMWyKfll8gXM0k/XqdhuE/1Vt/WmBYp8RZt3JvHlOYBN49yaZBFPbBs
PMKQG9cnBWzSGAhN6QmNEdGAvn2AnlgSnnOqOW8zLvsshAfw1bOY0/np+RD6v6oB
zADLOxfaJdnHyn234gclNcFywTZFhMz709i68hc1KNeL8j+B3Hc5QP8VZf776Njj
UN/1mCS7QHbL3cKXXmgRmQIorGIu1z27433F1oB3P6dRhphndUcrBxzKO8Iff5Op
BkKPKNPnMzF6uF5tS9/CiGfECAD9I/4pin5jGWdOVxvkgt4tYl1TQnL/voARHBnj
mk+mFugOY/pjPULmbzyQ08CkCYn+LPumFntHWkHDdBydTHNTPvBqg3PKsPMeNMEg
f5iXTZgRGG3ZxQjKiO4u8ujE2uror/PIFeqlNKPUEjJeV8yTUWHvLQb7zseiukgA
GjEP3oHFF/uWj33Omf4ZBdEkSCWp4/amHSqT9lp2rtrp4jqS4DigodUhqQIzXhHh
LNpiojWGU978F6lItQ/hrsGmtfihpWvxCzqcnMXeI76BaKC5yR/zm1QMuCUrFtw2
jPnVCqlcdjwWgfXz3O0PBokQPbMAlO+LJ6nIRrQCuxFzl+5d3d9/8OnGfdG9wAq/
4BZHYTugHxZ/Sr44bRrvGBlAsATBssj602AVGqVEE8hgeh3/MIIPdwnxjjSzHgyf
DT6sFzqH3nudUe97Kum9R0zzJRVHU9auRNZlpqyMpKrSFov6azmm4Yo3plrWSvB1
BnfMMuUEqoeM1QgWqysNUg6EQnulgOA/rPdtvrrKMtJP5ACU9eitaxbIpPQoNjT4
0mH831lE+OxVL8SmTlZjhWXVp/pppvvziFqAvHxoFUrCQirVf10j80WrHUORlQWN
o0WjStynOh3xmhdXbX3JuGPAZ+NFzf2I23/ScuVs3l0DawhA0b71Ju5jWLvirzJn
w7zCG0D9L2MaU1ARQSLz+MwwDC3BiZ24Po++2lzIoci2d5JGMZbo8LJGDj9x5Lma
zkixoXtykOVxVQw7vO6x9r4Qjv5jS7qRDaAu2k5PCM6JyOLpjskUYCuNVMXb24Dq
WcjUPvt8yTjyJp2NhsjmtXsKi/karpe3sA6+RzzgS8go5NROCukPrmZPtuaHeQKT
ZUczYn+xtHHyn7k95GXn/4OmoA5GhvshWCl5bg7eiKSmrA5z3ao7fSs8UfAX7DY1
+PeZ4xQ8hrsiWEgzGqvw+TjMg51G/N0cc55daMYVfQN6gOIZXL7ZMEColzjEOuRQ
7D+fY+Zv4lmJzZbJXpnE4WZ5fMrMeBRHvf9JYitgD7HHOxvLe++xwuBr6OfsGSST
Sgj4dacLatS6ou0SPxRk9lHeJkPpe8cQjqNr/lZcw5L1Y1PgUO47buRbYpD+KCzw
NNq6h6MNmSwRs7/yPgLCl56kMyMBIMheCby846JA+moSJcLOKBpZgvlkFp/0eNsj
x4O0fWjtmIlKWbwv5Bb931Q+VihiT6SS3SXtrM3ptuIO0ETb2D0Nu4YwxGM/Zuz1
SlUqYWoTErre8MoIOHWp4ddef7qxzSLV/elzybgdtSROinV+D4Bl/s6UdrW/1Dku
x6JHSKI+2lesFs0X9ZEfpz/CvAYzdy3DJ0JKkC5WWNtoOf5uc+it3EA4ReYBJ51w
mKItSwhR9PpIqabZKLEGKAo6EPDQFkRb8anRaqTn2+ywjZaJieWAqp2LfKZub8cm
7VHuUYy1DJj3qUNWOEeig9BNUn/9UqMhHeQMedj9+ko5mUSU4rZKBSM3GVHkm3NN
gIQOjwyR00G7hy2T0sfhgtR6r7VrEKVH5DO3cbkXPQ0Lwj6jDctweMMJJfr+Kqg1
sHR7Ny00LO+SBKwyqMhhYYarljEOG1yRUqIJVAFHMD+CLEiO/IlqzLslhqNkAsXp
AwGQt334zNfYwgmjJy4Ydu44B8sp168yg77NO03Fv92MvI8XoYz7NeGbPY4AbNzS
0NM1RRUjTLF3E18Ll72fKJ535Y1fPeeUYRi9oUkLKwQJijgnSmf33Scig5UFX/fs
or02xYlmbdvfKZwoW6euQjRzqG+PJo4sbdMuIheOB9NUsOXtoKhMVguNxitT75MJ
NQWyqNfQyc8cnhBT3g56bSVLLckw1ROyrhrC1Y3jDdgeWeESA8M5UrLdMeJZzUCv
5Sv+l39UMbPT42mpKzn8ju7mmED6dnqgkt3R4oj/2X3g+9E+pS0fBqqAQYAMlwKU
GZGtIbWyLNCCE+kLN6tSIwSy5scIojwv5olXIxyfU6fro+adgG/J5L5+ynf8Gj4N
fl/WKdelCiGEKtm+0Vyrc85hrj7Jk3I1tDOBRq1bl2bEHrj2lWerkHBT/WgPHFaP
Sw/mFh9VSzb1DxPMh+YlZLZOV+yOS6DXtxBbB7YmLJboSMgnCmFuJ2kHg8t58eav
UPYgGH+G6SgPA9FmGyIk4RfbpKsu0Rghx+2lzvT1q28pGPagOVGRYVSu3YywcZZ5
+wRfUZHeAlJANVnnafCfY8i2WkVMjgsAQNRDYAxcYaLS74TiQHPaDqqE3YqpcUZ2
prJZMRtU3NbkKyNOZPbLnhIhD5fVbGNonbAsAZ7phhcH/kRXquyW20EvJytN55KJ
R1GgvGq8QvCyIiRoH9chI5twDnIXXiwP3ENFOKmvjNY0SY8qXO/nJddIIvpcz1NO
AuBAQkRjFx/vsbUskj+Uxr5uhGgM0E1izaNwTk/9BdrrsrVd1CruT/basl+Op0cp
EHNvT55LKFPEFKFSRR+sGfx5awdAOaMgqmHPmyDkVWfQmms1r/jm+zVpC2Q6JpQa
mrzYgHnlcKhM9K0e2INV0TVFu7MXiWzz+wlPsJqSY5PvbjM9Yb4J8uNpb/nXvQGo
RkrpOPcPuqDM2X93HwwCo2WyRvoYx+8Y2Qc0t9JA/ohHXFaH6bxoGEykjuQFE4V/
csVtN1X6OjmairsEm8wZYUED/uGv0sOSsTaGPe2k3h5NvbQ3dubD/jhMdU4dSe4O
q6hu3Zh7APOxqwqPqgv5QwMno/pIg18lkD7SH1/VxN5PrlIzYP7TXXx+q+NgY6YF
5gN8z4b4ZGanowX2fQQajsYDn1rn8BS4bB3wVpZ81DSjsBYchywG3iph+O7tHMIc
Gwf4dYE5zkoJvvpZNoKYpzBPxAcHltSVoQUV+xUr5N4afRjAtePgG149frXv3STq
tR0RYud7I+5/69FnVd3Hcp5ouZ09eC1MYthkU/3SrOWFQVz/EB/aTci/Xwg55Yqe
fS2N5wGjmxifVZyp8OoVu3RSdBvbxKp9obJk4DdjaS/umDDVK1ZgrttvS2TT2TpV
TSgvKo1RhED4lBDwiuXhAc/WPHfzMPbbrVBfTKe8KuIeESDi2s5YyPo+b99JcTWp
keikrDj7vA6EkSniuOfM7ETUUFoHr09hSLvoBbaqUObk+Vhsh2jPcgj5Bh/XPvRf
P1bAsE4JII1PcAvgN+RAK0LBgtUySV+XaqxCqp1SKzMQFioYcflq+yNW/a054rRf
X2mX7FHJVti5dWrY6r1AsE0HoQAymBiaYvQAsOrIqcPFksV+HyjxtIZzAEXsKI3O
DBaxq+qz6hDFd4Wr+3Rfc4N3Shl8Vgmudv+qpw5A+xQPcw+QOxD74kWRq0bT2KRB
cogjM95iQbOxJbEqkS+6Twprm4pbArby5I/s78/1aYkqvveEsIhqTzFrZYNhuGSn
G/QJE4colvJSKuUhsA2z8iF62WE5a6hCof2e62ipkWPvGk9wbvSL9btXQEfHzWVg
w8Ko3Y86JkY+kn5TYxl9srKB80AzHEoT3B9GV1pt7GHfU9NZkX4u7y3pFupKmU/G
kckiNXzTJigYjL3xACDQt46FdJdTUv47l5+MoOqOEu/J3DsEPCOciRLncZ0psgwE
6axfnZBLduCE6BNxF0Dwm/CXN2qQF66FNO2LQMnjm1T008l7fNNwOJSkBziB+oOk
zVI6/y603Ao/nvc7aVKK+xyM8/ugoU0jEuT8/zsGbfRVH4lXLzD2ihjvQH6+b0Cu
YW93aN5bM7m9UhfL98JGopZWWyDeFe8NhDS5HRHNTy71S50MlKY2hknftp15iac8
yTWGRjQELr+MZX+RgELwy7A4qGAVZzSMQjqyZjQOOTWiASvcEKN9HVO3Dz5DzW9q
ihnSZFukagn0N16Odi8LWslf0WZdG+2E0w1HbKhn03U9fSjKHppkIbCiSqibOnCT
G/qPLBZZ/qOR6luZ0qxQj8+im8beFRaaZW/ZD2ni7pHp9Omf+P6Nx4Ro1sCJ/Zir
Uml7N6WABdiXainvOTLucgAm/nCWIo0I1bdgucWZWh5LYw2Ckja4Suj0pjFrrWaU
G7vNPxthwW+MQPwU0a+KFkHgc10qduxQBrePCFb/2r2GDcqMxKIHk83dkLUMcd9s
3rOeFNY3gWq4+FDhiRWoAMHa3EWZ8b0zd7HBeTWi0MXl6HiryHOZXSpH1VM6ejuV
cxNNtUuZR0oB0bQtd8AbAE2mg2hjPYU3hARmNfdKGPWOQk3W26nJp4NJLoK+JKW9
hAAhqxEXfukmpvbOtHgvXezZ/sLImQEznMHuRP5wHwKtQFLmOP7uUBa0yz4+NhoW
H/5Dx0kFOBgQhGAOKnlNWHELEMQ5hQkL+M6tXzH+AKqzJl3CTqJCq/6KvXUXcfqc
wwJRwc8T3JC94uMsEa3Pm/HN1r2U1EYHbDznjsuFXZBN6qreVzVDsMMFGwLufEL9
ihHDuCAGfJj5AL+l+JOAZlWa4oQw8zrn1hvte3bZzvW5W0usYAmpJLcEOCKMidIj
EVF+HVnAo07MwD8WkZfwlNz1FXOO96j5dlxrqjK7tNJqJ8r11GghNZCDKWVuRNWa
kWDiM1R2SMzJLN43KcDlXqNdVGGRZQyticnoqJ/AwD+MNvzKZHZZc4wAIJ9GcFak
4z6WCRTl5ttyIWhz3if/YKsb5c0ElEch4er+WCwpo2LbfdYk0DhbW+8X5oV6IAIA
Bp5CzhH311uYLI7LZC9A+NSAtFOcLMnYnEszXjypnFhfACnW6Mzshcw7U8RJW27s
4Udr5lej4X7vT9nnoMiMuEOBT0a/1wE9NCDti0XbXnET9hZZhE5mc5maQm42EWU3
wWt5k/8ahTtjuFHfJ5TRperw3YYkCjmWT2lZC6OtRy36w3/VZjv5X397q+pYPRnr
6WK77zRGY/9bvzm1wCN3RtaqDPXpvhpS0X+sIPziCn9tMldSJjZm7KQRbrBsq+8O
O9VXIrt64RjCrNSg2vEpeqC9AcBstD1Py3CSBDIfd19age4RcsFfsG0U6pZkJ+/v
S2J5aVvChAmgptKikw+IryMqvH147RUsCf20sqSrCSg3YTly1k+WIk70KEIKNi+/
8U2CN3oOzrrMpKoXRdDKCr2RoX/dfp6t1kCviLbPImDFMLMajV01Na/8avuwcsOO
JWZrrC62FTa+pM5C6y1+4NI8DTol27ubr9XwaUF0kf096Q+ItQUcjOFa9lHtvToQ
1OnsUsqon6DFINi+I47QemziOf/YcR8zX5UpKINuOVvIbtidw1cTzpcK5oiZRinB
sa5As3w/VkreXykcQRhdpg2UhCGePUCuq/xp2HEbwsjKGxFD2pw+SyGHQ5M26hZP
y1Y9LB5zGYM3ysfBQwFB/foh4M98KTuANA7eRNm/CyZYw+u+afw1gJTiz6UZCysb
aRCMsnFp6m9qpb9g5DipvbEUZaHyXIzuJdN2+a48XvJe6dR4Gte5raVdkRMfNfoN
TTGfx2wbZHlrSbyk3MtoBWspI86k0niFmPRniC2LRf7jBpVnN2mB+rR1ePsR3Ltv
mnycMJnntJB2WNjK3lSZgWfBZo9yZYBtefbAybR6zP/uvqI4Ui9d/YhJf94ZUcXh
YAdjXeTl9ceUIjRzjT7yMT7dJO0dMwiwQJ++1ApKcyg39XcTnIfwFsMalvX+1fBO
vKxvVn9wdxaeUuGtRaq9FFnua8Uf74ihTGh+61MhKsEqfNsPUjVR246E7qJ5sDeo
ByTlK3oHgnw6ebqabul20P2OfGNgBhmHimDiWmTZlMdRJc1sbOQnYMYdvOsS5/Ae
BiWU+qrNw/UHB77NT+2/Ai20ss9ZOfZY9MWF63KbO06qEb/YJ85oZYTI4hppppM1
7I/qvKqKZgobDSkTQBuCN7DbnJAul79GklpkrcNopkNp4pHY/hlgE8j6UktoDi4L
bjOJumZua/WXqQZWfnXTY5Z2jg3uaZx5xcXz0NYAjBCNy2voXwX91GvNqZzYBtU+
CCbTosUw/81Nioc3R1DTz4qO8dguIrOQEiSMZ/SMvFDvSDUEVWBnMt/UQr+k8ThK
E5naOU6O5bf6OnXwL/bRwSoZcBNhfuU8I2hS3zr3kwZkk0b5zqbB/CtOj5jXarDg
KsF1VOf6ZDWOaMOTzQDIvtV/c/fl8TdnE674PDom9aRP3gEFQE9f9pCDSBDLRgD5
2OF8jIgfttzY0vQidkvBRa6w8BeytVRkxQb+DizjlBmeLlXCJQZ9N25jy+ItSvfv
PYuNAB8VJuuuVPVhmmHZFvuLHQzuJ77KwnW2AMIRb30bgJooFSCP6TMtOH7Mxzci
FewZliaGgeNRa9TewvPcKyT/dFwCXa183rVQaTs9SEVSnV1qX+MyXkxQOj7nBItD
pF4qjGjXBPTVgDZwB1tOKnMaPX0tCGlNB5G1yw/aBvZMSjHaBYQfNiUVqPImD/Cn
brGVyoevV8xRoo+dEhGPNrGd8Ljqm+W4niwpDyNs984Qv0P7/MsPkdEB+kCf3QFl
JFGChfpP/xPNR/4vBRQWnxsqbZenuUSWUDnhFtR+Sx863fDW9WERndmwigKvGjz9
dqTJz7VX9WRK38or8/v1/lgKjBdijgDWPN2uYKP4GIkYFLt8V1bZPrQJ6S0FiTSj
rxSHL6P6oNPxTDvcDu3eyCHuxXGa8ilJQkhIf4pA2U26V8XMfdkcQGUzUmOwENfm
tTLWAFcOEQxQrTXlpQvjFtH0gkzdhqh5EqInPOuFXQpBAP+AGMrcIold2S8sxMlj
SEbnfJThCzGn3o4j+KEzSt8j40LqouiRKDv8lkRcz7TCXtUQMWNR1s+H46dFU94V
WiTfSjNNlU2/nqjuAi0gQ5QRtJyZFbAyr/oWbmvEp5r0OLXcrNGDbRHDRURfNYRE
qNku8g7sPWgVFlVyAK8FomUITF/0Vl4emtLh3hxydKpPHidoOj0cvyl6Agl9OEJl
KrfCz/tHQRhpadBGaLmEM8w680FuZFX5EmfSlCIdxvK+O9qqOtwixnPDaseXmJke
u8/MDZK5ZY1urCXc99I4R+0dQXufx+Me5bRULuU6dtQcQOFFdCkUibHUI/Hmo3sY
PELYzzyXOe+KMVdH1z9DhFIUqtRKXyg+acuSDVVBe+oNBfw1XVUvmD0XNkno+kjx
qkciIptpd6+or6nZqFaQCVwr9sWLP18ixsnohZCgVV+SCiftbu/37GbGZbJpM1SJ
Da1kYpoycck31pfSopTylerMx+jK38Mf8GJC/kMKjBQq9INXxTE/BXeuAfgZhWZY
o4XzQwq5wDD9wOvwxx6azS0s56i2gp8YMwn1ui/PtElXtjDRBzGq74SRpEA8vtIz
GLacfJd94qD9GN3rRJODZwvSmNSCXSlrra7tSp+Ba4Dzog10T6qkBYOUL9ZeB45b
tWpo3uoLFk+xBo7mEMHqjMZbezqrPY2cmcM8x7oxfIFUYdGBUQxDr9dvzqbnTqxh
/L5/mNe0iRTM3SrGUdm3DaXjP85QASDVbQqmk1N819nPxTKeZ0xwa5hmEYKykR4F
I7WaO9ot5LhYTg+MhUKkHhfdKJJBsdeDz4e/Yj//LklUCtSgVpLfPG8BqcgrEJt2
4WnLbnwMTZoSlGR9u6ea5CMbqS7lX1LBLMzG7u/ucQNXCrB4CPd/peBIfEi3GgzO
Ymz8+mvtrH9bxzXl2mxD66ZA+5NhCzOofqAKWCyoq6jZMgVCDAYvtYDt2WDxH/MZ
2ObFs54wdvZl4dXI2czKCfsd5oxc2YmYz6pw6HvRESxCCVPASs65xgcFDTsNX0Fq
QJkX6VJaCFEaD1uRjxuxERw7lfTBoe5M7ZQRViz66Rqa9s8uSSk2KwOAG4AQO9ty
12tkdt0XkowEej8X0P4+l9ey0JasXv5mYhrpZKyfVWvK9+dhV4ca+7zzdA8LCnsC
JmEx2AQR5LB5VJw1hwXRUXLVH2GchzKIofoIuHqnJH78R2Qpw7b43J1VVEEghi2p
eVmbLpwQF/ehDYQQmQTKgHErogqqfUrOxJMBeeZ+aT5d4/zJDhE+G48AdAkkPVx8
r/HZUHYGoHJ1YSSAxPMAMYTbHP6Dp63+cFgvT6eKmoko1y/47f9qqqzUTViv3Itl
uSGFBzlrnk+/gnbA30VN8kULc2xHhiScsN8hdtbnuEBIGEmth9iza34Lg26phR5u
PYPGU5zpb3uNNdyNm1t3mDtxop6Hun9L97HyN2XCBGf7l0IQbahyD7RsRU45vrJG
zT4FAysYopYkHXOSGSSrGHqRCw7UOhgzL8VFMoGd4gngK+AzjVH6Ur4oj8ndOlZp
i4X5OlyDCIsmG5QuChM+1OaRkFuRU/PxpUND95CgX9cIZUnDeyxA2gqy7GJpYf/C
J9xUj33TUW2aS2lV9PrEL1BgRH4rHmAaeKCBPsMDdHH+S9im2c5MKNDck3v+sFmi
wdO5KQg+979Z81ZwSCjRFvz1U94uQadG+6VIWV7H+86yYa+sxQ7tnQCtLB8wMBVb
A4oOlt535c35HqMDUhL/g1YnKOqTesdjQvsstJ0z+8Cz1+72+ExnCAoVaiXOLUUX
jU4UUdAVCRehF+hgTGaSQbBuh8rcpm+QYXRQKBPHFvJ//bpsGAhZ3xcD8hT5cXzl
RPiuToRX4d2XylPe7jYEH8Xd5T+DLAw48J6rH40Hh/mv0NRmjf6Euv5FD3iT9AQt
DJDLSKtUAjC4ytc18hEeNC/5AlUrsxyyV7bgUFz+O7QJ9NOU8uwn0jye8ePTd2en
5pn2bMnMsDb271BfYgsMNiAuZ87+Xaccd02I5vIOKlW57HRSb6WufGTxsWk+u8hz
bY59fosFZH0YD1jI8P82zLYqWs4iKUe57UqX8q5+I9QATKn/+N7kK2l3ORbTh+qg
ZCTrGIsweX3HTYZvn61V5uJKBI/EoL2KB6Y28IQ71lwdocW5sJtmI7MNM/obVmmI
EF25MG/k0sSEBeMqiClNSVhdq8TF1WuYZgC1A3+6yDw+TjgrhD4JbO6vshh9fYxl
+yxZQvaTNDl4MVMQg5wPJbhgpCQyznv2Wlsfuz1Et5KQbbzzs8Kmcu3joF9t++Wd
2HAdqLNs8ahbDoG3vYdVKqr+mqgHFxm/PTJwleetyOdqTU7wmemb5Gzc8UsYAUMw
ZIFKXuShXYHZCNpXu2COaRk2ruP0Oqtm5zmEwaj3XgSd2vZv4XkSJG417H88x2hd
hSLHoToHOa1DjaX8bCzp2WarWQ9vz6IDGQa3uzuXpRmxWlVrAEB1Eb98JmgpOdJv
8DLul1IB16SxHZnw7b3Wqq0brfubTusTkgDn1l8HFMDpzybhRO6ixnC6UitDASlE
ebRG/GmG1s4zwKiuYM3sUWVmq1Yjvg2vL2/vOWDhMUgUQQIatrtlNKrpJDwWNTER
V2KsUjEGpL8r7hvoAeSVpq2KQCh6Bll/KTAkajBOrxN7sjsLmajiHfpTDjt+u4+k
fwNUEmwmoPLwkZcfnvBOcosGjjT8x+28cW6kJxvdWMqVRtBtIUWfNNSpQ6Bv9pUy
jJCAVdHpJNNF6pdZmxtYFZvCOpbgwspoFSbgO6P9m6bss9YObmlSEu7M21oCYndV
Qf1P1CdVKcDBo3woBjh6dzKh+xTe1D5n8Yiqve1/KvADKNHs5qwsx9w+jK4j6mbr
4Ean8vA0d9tT2btkYcrQqSnd6mrYYZXSsvrEA7XafAf6NWmin6/RroY6UMQKzjS+
kKC6OwAGmsOVImILxB1g74dfVdOE09UvZbo+VkW6LwSJODEZpYlRIdg2n+0zZAXv
lbI8ZU42VbYTLueykLe9ychifu69XUHiQK6V+Mm+RHYl5C2iJx06JJxwwTQGVAF1
npFl//1Y3cZsPD8qY/d4Rjmvn5g3S7kNWLuvXOnvN5lVPiXKj6iC1wGZIs810PIf
RL00HsbsLGcZrv8OvtkA/3lJMPKVaq61wYJ112S6G9VA8mSrZ3dLtie1RCTvu0r2
4qXQuInra7uWh8iTUDrs3OlaQmgyo0qLM6t2GhbKAzfYmKpEkkyqLXyd4uKr4oEs
a8LYWtgVPLm3ayRfDWIK3phvNTP5oXVTqkBVZ+HwbJdPUuOnoUCcbn+lofkpVTAQ
jvGVv7yLOfwbBUo0tpi0MohRwTwzzEgzi+a3yM6hGZtNybZ82BJvZ9E0D4sxiSAK
CD1zQdDzzcRSdybj8FwSA2pYqM4Yh/K3a3JphnUMIzKMObe9BdHOpdSCNbptlfkO
dJPzNDuwpnlMXmedfTLHTS4D1x33bbMpaoDTSerlkDgeYameDnYt3YZ1QsYhuwtF
5TUMYxZHeYwjUtYpurXxCbxIqoTWhmGuOkuMLflWFtIM4/0wpiXfihz2iaWlMPUl
5HalAUccrjnkm1+uJD2h8cEv5okKAZr2g9fduMrDHAo8kK31kmOKPxu9S21wHbP9
/XOK/EQ0y1UWzt3j7TSBbCPYjanOEi9MeTTXvu8tnO4OZEyr0Jhod7AVI7OHhaII
Yc6Fw1/dtmLnwbZ/fYi2oYBK/ETDNheMO1tOoo8ZUVgfLCHAE2XY/hbNp7GoXc26
wJR9te43b8OD77QdX7enR5/seCbis4QzLQkQzz3D/fbAVJ9lXhm8uw4TUj+9bI+Z
58Bz8vHOCoYcwWh9+tLYnUpd5KnkHdWBnPos/lHZn7E4llwyIV/a/9NvO6MPY4nJ
v4KQJkqfcNoXM9E0toxHArOI6Hx7RW37w5nnKoBKZD1Sog+ch25XHdPYHrdY9db1
RMHSxYh/AbAfMIDEEBNsU8DSRVH262fSlDwyD4C9m8u67cT+ow53v60WvURVP8kv
lUvGEptJlRL7xSvhSym64ivKttbhiF9TTAHvY7HIHeE9AI+M/Z2n/DPQ2IzIdnjM
pQ9kmT5T7esL3WNwB66qVZhe5QNQ4II7GZ7JibayyiLnIVxvuzJOL3v0VdTaoEHS
s1EIduh7viTg8MEKqniE8mLqHybXxx96Vpmi1VX2mTsqLdNkUPEGfW4Brw/DSBmQ
3+Ti7bibx6n5Dmn5PzqDw2xGbI3/PnkBtnGgdo/ocFuiN8W868F9BzR9YAMmUeO/
7t9cQCpU+TPDGHll5dYoedL4UShiOOQpENeiLENhVQyEDcysbYqkcqtwh/Afdhw2
6DJgna//4YBGr31hMoFSlRCrNNwfpIYLhRFr+D4RHpr8y7teZdBcCpVOF7Usrlok
dtDMgnQIPnMT9LT79cTn2JQeIFHGxcRYRS3wcSATVDFTa9sW1OdT3uAJh2d/GdWa
XTLqeQKDXHx07mWZuqshXxWXTpQlhSuyuQGY6Beyh0owAsYb77t45hKTg1l/HDAZ
4PKaLrEIQQERvAdvABCrQj2vCrhewPV7NvEUrjp18vIYMb/zm0C6/mzFh5YzUVGJ
vBD4pC+sVBycgDRijYYfCU6qdmHCzQJrKkuhi5lYZtdumOHSA21vCOLiUB255dyx
/rTbFK5VT/z7vYHTawyXb+F94VrrFUKMF59i4c+jz/VbOtFWmrdpsb57Bvv4QY3I
u9y7IzA9n+rCNY+RDmhIPB12XflaZG2ePNqkimw0NCVwsh3sYGeGHboduXrTvc8V
PLNebGb/6cmqNsUNEQ+u6TT7cFYkzO3SWIGnshZ8S4QNjx+avWgCYiKh7FbJyw49
PH8bKcXkeuj0p0Rs6H7jzJ+aLZq/6lnOYkR4HONuzWqbjBtatHm+F/LQ4mb8VapX
43Yc7TP6REtRtERR9JSInvoGtR1B74QuGoInRyeCWday19mi/NhOzymyp6W6t0QT
VXAHLYhVBXcy8qPmX6HbayYgEbPWU988jFyyTztHTNfD3lMi1OSQkI3BIj6nZKvT
aKmL2BRZTCW0vB5PvmGNATiZc4vQnEe2IMPfVPIv8/+f4xBhhMDENUsML4Lj8T6y
LtRWAom2j77r3D6gXTxHsYZAS78FpDQJzUSDn6VBg3u05eWvcmo4+sdQPBWwUtsA
AFz4GIiUrQR9NPL6KgOhxyaYiUTIwbcW/S25NxGUMEMMYLGOfvHjpZBhaoQ+aX36
ps8g+oJ1pF6aLiyVVBTNrpCA9/yNB87s5oAppcbxr6ijHIcNpWk0F+tOKBPYNcio
CRi7eTqcCG6O+jp05SjH8HprfjdN0iizPDCT7urcTXqx6wW3wtEuO8kf8NduGaGa
eufjOEy+UGnCq3TReFath8eGJ8lC7K2kzLRh3ptPo4u/qoZmAkeORvoS0Dyy2Gdk
C+I+oLY3qUajSHoArM58CSfO2xNbQnb+8Gg3lWZ9k8Ur/zfcisz3iGHqZLjpjD/w
qnnbln/ONEgBvrXf+mceP3RfpDcDRJacvPVFm12jhconu+W3QG96TqMwbGWRi8J2
U63iSdniOUcD8ehK5OBw+/wMdSq23BUiOf4d56O+JNl3C+T9ecc0FgZfQRvyZ6hP
czu5GK5xliJbuQ27As+dnpuIo78l4cUiLCdSz4Tg5cIC+m9tuQROZFbHoj+oK0bK
cBZ7M8fCeTV/g3EDN4c5VTbda0dLzu3VWrzEdK/4YFWozaHPkqZXsYoaYgGawTuc
nguxED6fsCrtUURfm/uu7v5XfX0iVJeyGPAEHaKS58p+J5Iu6VILu3FuQuMjacJi
gBWKfHY237WaCdzda0xOMMG7ymTQ2TzHhD6KH4nc+gtzanORUxxft0U7C3ApL+YU
+lRUOgUHWn7Q0HIKRBcQsvTzsI2IY2WkZX7uiTWrvilfQQk0xOPnrC/lTSphYaZO
LiU5awWaNIZdL0ONEweuEsRC6f9M9wvgVoBhQApgPs668ea5NdtjcsN+YKBVmuPC
+Dz+lGFqej7qdPN4Ut9vtpPq4JkU0lO0IOhzxUTBKkbDWzp4BTB1UJYfoyOP9i4Z
+kOwI1kKPBdVQWwZK6lr7ZBF2o4jBjxJwxvttTKj+HEQevqYv0PdOny1Ba/GBSX/
9yFgueXP/GnmxvqGjuwL5LigNqpOi88u9z4IO2JSHqMyyJv2gt2jpWCYcFhts2ju
k8nXNvt0j4topCxbEVUZVKObLEfIwtqDOI6g7vnyiq3zHGucBwWNNS02urFIvdT6
YZMgmS8Xw7zWLdJRh7I9W6A+qHgyHvVlEwArbtzmcotkkPypTpojHjLKuDCBx3Ih
c0FMn4PSUuBjrGLby0vEA1o6fn4EXu7Kg8ca21y+ozyt7FZjWB/rxGDikuR8uWMu
IfQMEFlGcr3CQSolf0U50IBG0xpyj7joFsRpXzukULuLC2LLR84OpeRwRhV+2bLC
4gkG1p6M5+kA+ejvLoB/OV8rMKAnzk9MMj8UjTajSmHo4ZIWnbqb+LZOhxFI6VQW
zKamt89JjTJnk6n47QH6tyiqJq55KrqUxNDlTrcp9F8dGI4IhlXpOVSPUBQorPz8
G5jMFuF4XkjTfdo96AtEr9WSVpR87RGquL2ZucGruyYpbQ7HJ9mmWPKquy3Qvy9X
jqKrEcI6gZRLW9NMGrOOglEgrm9dBBxUT30ANP0RL+AAhqaKpWQlbq59A0u2KDBw
pWdB5bWdIp3qYSSLhnUnsMcRzv7SzsvA0wObdd1s1xbVIMO5jJQpFmbtzOZaWJnI
hnpD01psbOXb9GWkA3NfqyKEgo+7WsyQ2jOgdQfuhnNJWOGkenFDD/lW+mWfGC+d
6xIvn4me784GYhBtzV6sohl4owxaZJhpysQPtt7ojAe6j1AfxV88f/RQDSATSQGT
C3BoXO2tPlh5UfuFLmTEKQHeAKUyJYLBy8N72x9EMdxUOzkVvL3LZKg0dQ387VRx
eYcsMpdqMzf26nXlyT2vcgpYTtgkvfRUak/7IVh+Lfo/YiEDygN+UIlwAW6ujyYI
X9O05KZgxrujzJUMHvdaQQM/eED6dNq0Qjwkrz5tDCfB8PZUUClja4wAhbxBK8Tx
eCl3Oc6qauOiCQIDsBibyt7+JWF26DLeUmxd2y52OX/P1iLCIwSaOJHT9/1ZdhFu
dNDXQPp+ddPxz8DBF7TqHJyawPWGAJeS2A+n8ggU3SzCmF8One7NcBHiFzn13Vmf
jE7lt01mGxIZ28A7ofaFPnQe5hMXXTYqmQIEjucP+5UW+FC3HDlhbN9hwKJL5Pmp
uPUWYcG4Jim2TQV7CVGBzmyN+M65SsQkob0/Ol1y9fOtBI8HLUy4wzzJIRiPuzQR
/6hAzmhL4obtotr4QPB0Vpc2X9vyk+MrzgYiTVUI8Yn0uFZGt5AzFeZ63keMk3B+
R05lmHVgxKYCnNX0Z7R38khhfUKswz+IPQhT1AFbuLUUK3aAY2v8uo6hcBYlVm/N
vpp0Dpoz9vW3HWV0quksnyrpwBa2OPpxlEWHSN+EP4fXqbkiAgTK8VL33DG7IyKC
U5nWOCVN5f1bgQDzKArAeSA4sU580cFfGvXTilRhgS3HsGHjZ3tY5TBYkF2SQNLE
mWoSvqLoyehk1bPEbpouIKuotE6XvWzypuL6A39BZHu5gvboHFMCq/CR1MTKm4ML
w2+OeiSLGUcqgudcmOh4oM57tZ5VqML5c8a6+V85sB1nqX4XEBHLIiqN6x0rtMh7
q3hjhgAymo0Gt9WfiPy5Iy4Z/NvCpG/qTr7WZ7VRJXdym/9+XjJvmZ8jDK5KLHxe
c5sizj6JfvqJO7AU1DE1IqsO+JN5bCMhem5B6CWdsmMSprlP5VEluP19Lu/VOjxm
64onRoCxGZ9KtJxU2fiQkRbo5fgzdUApEjnXpPWZOyKRVm5tbB3epwO92GHGVG9W
1uRv1st5AXc+YuY3ESl8Mp2xjn70UZ7qpvnrVMpYJ5CWJqovy0r9F0nZdEQ8j2D4
f+x7udu2umplDHcMn4YJNfffBOKaQCew6Ei0eEQczlQzY945t+znW8APZ5FJBpAC
y28IbSnNIPM/sNlue9+1kUBz3K50esL5VNNt1q2MGXVdqFE+V4POrjTCm5es8/Bz
VOOBD0REK/OAiDRyfdWTOHj/ECbUDkBxiSjNg8hMHwBGV/9wi6j//+RbCNVQwJ79
jPO1mKI0EXR1XZ+FR3wminieYE+JjWnCA//5Ykm7Xb8K3H3fN2G+IBDT6FbTih8z
wP9HB/343dofo8VOwWHd4SkncZCxFq1Ux+2mJs2gOdW8obY+sojKNe9J+lwBm0YW
JJF4jgBinsHl4BttxVFqJAQdNlrqyL4qCVrgj/cR4e5131w30pttHcmdK6zSrmHN
8g8iQErh2R9bRlIS0gJMQgtUpDMH8gYpU2cXEd+cj5sOStLl706iHQad+E958Btm
kpFzIPmhbBeeMCgXJcPmippYoMdkaQAnFt86WupWv0qhPCqpotr2/ZSscN0VfM8Y
OMUdo/9dMbTDFW46/XRsEOpbtwhlSORTusB/GQioNQYXVtT/11207v82+0kQS39n
QoS9oxHhdUUybbNeIuw7QmmOfUVYRYXTuCZrs8Bn+LOTgQsyfesA3Qr6NM5qiLyb
z7lTY5T6TYfnkMQQmea5YlNP71gCGtmIgWhWybhz/Z+JTNpEiploofR08ew7uvTf
x+MQgJi1I50IWd3uF7Ujaa1v6tfAgBv9hTs8Xo0+kQNfeIexW+muNtUbjSf8+GRP
y+CdvS/Z5fYY7rwyUCM3TgNQdbK3WSbB2Lgtob5eZ+tEXV/Xl4WZXNziYJlbYQiM
FTAb2+Rc38tKywql/vQWxNnRRT/iqJpZtQ1ynB6TTwAXi4qJ7Frr7JJEHqZt5A+p
2uYIlfeulPzw1XLyNa7eJgWDZ1Lnm+hp0bQFd2VHtOGMneD8A8ymzesPI28rsDII
Bh7BasdZwMZDM11aspHzX/QH2vwcdSXSltJMapK+vsAHq7rLUEhXz7pMlpK/ICNo
LFBpPkl4ZcUC22d+rakdOJZ2FCsVZ39t0b+CLawe7Ap8PQk8rhS5RU9UAxl4Juim
lb87JvKdxsJPPvOfDngRZA/Lii8F1pSvGEk28bXzbbI/ORgah52g7noQ06MtsQi9
XoKpB8eO4TAwUfVGQfyK1rxMbofN8KKY+WKEAo5dOMYp/Uz8cPcZtX1Q4LGCikSN
v0CyjIg0JdeWQa5t4+R8khPhlEF/52R0av5kKmiBDjwMly3lMxvLi3lxjsh5Nm/N
3k8k3l08hhbZZ6OcBOQfFoJCioZyBMz0rgPucZqqhiKIgsySdtx8JY8k4VSAnX2J
X5+NWm+mBRTGybW4Qnh/1yOKlaBDq764EqvLpZMmDQXc0YrqEc5wXA7mQblNZ57+
+6y7u2dFHMkU5FZITynyIvEtj+rpz7eCTCvir+eCUo7bveBgf+Zqn+bCEsLvuBDk
Z3W6lIBtXindY+cHiqeNnvwROM8qPH3UOt2cZhfToc1Bj1LEN4+NIP8XkaEJwVTC
+taVk36U5UW/Kw94isuj78eHUXZ8UiK1fjZgaMYBsORKoBsxua9B8Q8cJOeBh2Zb
IjqDbhQ5YiYgIToiwGy4UW5/2EXhc7HPUsOPjWTrpxdsQOLJwVUfr4bHYuO7BzHw
8uZniwO46Hf+o4uB3+plFzel5YFotYoBTBrwpUxxXs6MIKmby13weWM1I+d1z1hp
Q5whzKPYbGU3rFw0VWrppxp/7cLmRKV4JKmoDFKF2RHvRx82Hf/Yt4alMHyFfkwS
EgwiKDdgpAOf2Bd/fgQ8uPMfDs9rag4VCQGL71tyMwffhOsNn4bts2T2G20JzOA5
hxRl25VDBwf+vLU71eaG6/HaTvRbTpcd/pWzKtkxmAp1eqw9My6FBfi1mmSHbVL0
NXiOnb/4FxP/h9fjDs10UaNBN92+++V8Qt8A+XevnDQaJdsHK5hMLZKIqk3+aXru
NizT6o4WIjgWij4aWsEf81PgyKpQvMywvXRkRv+pZ3Ui1KDq2mlPZ+AOUshB3VxR
tuI10lXBKxj5Ql+6zoHms4s+uJAchJusJvoDMUdrFhTdPkXRb9eR6vkKofe0N3jV
8k8O/BMDa0WGSwJVf57YEg3kqgEVLr5XcISgb4stiWRn4rjf2xJUkc/MibrVxPDd
CKj7xf98A+8bY9WhegLEyVYvm+XGyazh1d9mmDYXag992Kv1Ja1qjRwq/RYbXFxW
8mrETkBTW3e8GIGbrtbrDbFCQ6F82rss7yPgUUEpdkVK8BLBImRjEngIOnLsJC8a
JToX53F85hLu3t5oH6gW/NjfC+J/plKq1XpxD627ItSGROc1okxLCIBbbuU6/ouZ
NWt/Jug3hK0c7M3hMlvKRsq+rx17Qm8GqLp/czrdGgn/bufZfwdcmzlJDq27BRVm
wz9XffWMpt967qiL1Z9oiEa9/KW91+SVYrTmOMbe2WY1FzxA62o86VQ10sA+A2SZ
p0bDsizserLD16ievnaQz7rAOyPuqesgF/x8ZVdihCA2NDGwAXx2DVuaJVa9atAE
JSlogg271g2kITQiwfQ7sU0dZ6X6y9wYXvqmNzRFep+8UGLinRZahSPTGWNNF6de
YDTA7rsXe+6aldWCI8So0VUSOxc8GOS0M6vO8qrQOH5xR74UZemjOa9dngmB5JdA
oS4FtqnCHwDLuxvgTU+q/a29Ue0N8Mum3TDUGIjAJGF76V+hBIOOdoxTlFG0/KBJ
xWLS8sfEWt5LV3oPg7qQikoSKYmSLjOrWIQvF5KAJY2HZyQjb+4dpaAK1QKto2wV
qRS1ctkpwauvPuLv/rt/7hw2Amo6nthxFVGDxHXkOKhixrv6lCf2/9RoNiK0NmNN
L9dn4eMuPxuO/E2/i8OBUBpdVx8Y1p7Kau8rAbOlIWErmhTT+F4JVNdBM1JA5eJe
OdojSWm8Y/25EcnOS4S9I3NgpJWw3FeAQRk3OhWxB5+m6EA69NvQvazpfDGIdmiL
MDvFapFG0hMB8zb3T7miT0hMCgj/xZ5A+q5b0miYHSOi1XlLXwTiUeS2DtOnV849
Y6Jfpzt2teceyc40yZavmRSvN8xQ3relP9UU1OqxmJYy7+ybaWEQ4pYXA2JmMGrb
IAsHaU7IvvY5J3nc/e8gFJ3uQ1PkFNj0aSuff9K/sFc/Jngx2T7XkUFThY9F4+Jg
g77l92hS7L5uHHMwi9fr+aF5EfBKQxlmi0gPHq/1NWMmJKteSIQXP3r3e6PssnA9
bEmFthh5mqPJLqLwxLJR2+UKGR66dTx/UQG0lx+YMbU/zFaML4yAX6EOZFukwNc1
Ly+0qNeXnIUOPfVVwxtcHs08QmfAoZaAuFq0Vc3Tt0rScu/o3EnW/gr/Si/FORSu
rOHJ92o0Xpjvp1F/R3CiCIJMLVxNpkplyk6rgkecZ+VCkZtGIsSzUBHTzhL8KUY3
pd6454BmDM+pbYH4avScrRuIDmAMxz1iFevDF3HA14MuFPdK9MmCdY7oV6MGXexd
1WkkIgW5Q/zqTKpFBlYkxAQyZ6D+nTvLDKk60oGNgQ2KPJhFLKK2g3jBQkwA9/1p
U0ucqkUTK1gcxRFsT2/Md6CxLE99G/iZS0TzR42VjQDMOdf6Nr2JdYG9Sg72ZVds
9XV357ON2zvRsih0dckUjNl7scZx1uc5UojemOFAqp523rovaYbsYn1i4f2IJJqW
A5Pf8UFfdqOx5qeFGur7QC/UwPv5KOAQMU8lI362UJPQKlxZBgPyNLipkvj5xal9
et9ZrCWB6Csfbv9YekeGoZHIgf4ZES2uKAe9+Ktgayj9cb8u1hp8y2b2fc2ZXXPK
xqoDekFd/+hK0gh4kv3jgO5ypgIrG+wUv6hct03pEgzgUHUwrQT+Rvz4WynNVOlC
s5KOCz/akytblUPwDa7pjeVo0TElJs3lodYD59joF7lDNMSSxz3FO0c9AGxZb5u/
yfinOk8foYBvpNQHtOwBi+1nNws7HgxcLlykNFmpb1UXiJtU6GS+aY+CjfxZoV8I
6imo77z5tEVFm3RB1o+B/9fzFPCjin82A2ILD46kkjOebJkXwiI39VjFyfRIsFVk
/vFOdFvCPWMkZiKK8K+F2V4eJnX6uh60Xop9ecCljErTjaEE0/hmIcr1wWABDr1p
f7O35eWFGdZV4F2rjRk6nsUwhm4A59Zh2ZTRI/9CjIay/P5CJnNaZebNoox5GRE3
XVeebmEormFagsr2FgE7048jcaN1o5dMzrkeG/HZl6wrtejVf9MLaPSZ4JivMJxO
1TLKB2iteuhHlEgTeWcYgKU2+5X0NxqmNAv6psIZVuJ4wvmu1U3RjtRGX7t4824O
c8Miz2Ok5KR/JUJWhHLjfEcDaYjpVS4lac7uyxrtSE/aC+Ep1KxboZ61MbsGDhfc
0TIJH+Ie5ZHFcl02A+nKTefmkyUDgv94Zv3N100HKRrb6gxKsfXBKVcxBksph9r4
oXcUaDNXpBXyK8WQVwCtwpcB5wwKBKuBkUPYhX/9cbyataxWfLZ0KDcMcfoXwoTB
/yz0RsJUHQi5yBdUirws0AED275j96yQy+RKtGxL4IJJGKcmArisF4YZwT6bnv2N
K9ioC8102NdlpzFYotF0VuuPvUmyCTdg5LkvkHExf7FyXjuGyeIM4jlVP1zIJOkt
koUrV4SYqyw9F4KeqMFSPJ8tyjWsfyBtxV1a6xQ7xhGi1L3YJeDLD0BgJXJutlys
9bPS/V8Hb5ifkLnRb4AAwSQgTm60PT1Ri2u/zZs9ejYnLpCDlCWyah3RCzRXLv7g
YkFk0iA0b7Myd97Uf9q2gHZYCPhcUihqpMRf5UKVerSekVHRhy5x0+ZqhY7AL1bV
rEBPSnZvbae7Qcaa8OiuHW4scJlMJdJrr+NAHbEhhViRBGbJnZv+YVus3OZCTSgM
YZRRAY1yBRZvuHv5HO+ds9S65i2Itfd8ixcJYKyo0w98cubPu/JLnASfIdZ+eKwU
EUYUUw/uRxmflPJGHwAYg6g5J0ktFEHtmwQTklvAYQ7KTuJtzbJThHkAOHsRDBs9
gBjQjc8PC/Tq2yLq9xWE1rANx3w9e5t1EUZXpZ02UMP6ClDu7wdUQmNAacnpvLdX
Jkx8LTMN3Q7LiedSCiraODedSy9U+u5X//YdrDZL+wU8c3SEyNLffpkuS7u98DiZ
00VdBpVwYo9JO8iSM5yg3FdmOn7XmFH97imYptznE6RVkEUMETWrwaZmhMUpMI9v
XiYJzUWsuMIlyUgJ5zgNepB7LgvdK18QwA6mTV1kfpo+naxtQsZnkT6KiFX5Z/Ha
JbWYDtnJSahRp0a70F1DQI3CvsRt0K899CRdANdEXwRCU67Y9sQ9Jh/2jufdvVmL
YQmBr98Y+xXgyZe72kE4SHZjqb6fYLta3kCr9mxyMWTrU2+fKeYPM84mWAdlfutk
x8DvB50LA779Aw8lEQLUTDkp5vPXkJME+R+pNVEh9+R4m7NoRc2LWGrF7AtNkd7w
XuE0+2a/wFh2xvHsSPFgJiax3aR2A5ZkYcwpmC4Hw+oMSs3E4PaB7LtDzQM5foDY
2oMyJEb4LFqPDl/w8YNHwvlmLMpax7e2sU0xgo82SrIYzE/quMKAcear6MeSZRTo
FQzaifbhjIcu7VINgYlvSrYS1QBBS7KwHVHaarkVKvz7uWyKpXblXQK5abfO2LN6
swUCUfCbpBejjeqA89uwp4VL/LB8siuvF0lB/1DUJ5vHe6ifLLChexURyjka/MZ0
aWAetgIFtvJa3BnWaQsw7f2IuGUlPa0yM4JrT1fzZXr4O6RKQZQBye7Jltl3n1Mj
wgVmQgt0fRAAosqV+dMafXn3kmtV9YVQIHlBAARMTEFm4ZeZ5Uv1ZlhBd2f0esou
VlCWlbWgJLCQLw8Ou5Hg2KmRKMUPbUU2fhTGR16Qh/abnANUwJEN2yUZEHLDr7LQ
UM38ZxdRdHFe8Y15IrTi5YGsr/ln3doVYKaWZXeN5U/iyrzCPGwk5Jv1QyTVOaWl
L1sbT2LG9K4MMGQWapiI/LA53My0rvu9eKKmcRjl4iT/ZtP/2URvyFLKfuAQXg0V
wlpkApfkRNYMwoPE3/iI4fqHHCSfUCgZJCVT1QDjxWjxvcM7WQGffaJVnJjDERGV
9xS7lsjXdaRyisC6kIp0d4RVNiiFep8YTlguVC5mdu0VAPTbJHneRX9lzJnPaPUJ
DU4RQhg4RzAxPH6JPIP+0UZ/WYnyB5SE1njV74F3EIa3JYfdK623a2mHMXbds4ic
yzg2i3x3Mz31tDz/onpWU7i3WNBs7KYKR44ky+HUC0aN2fmEkhiynaVvr6dKzYvO
2n2tsSa7bsYiIo6yslRQlImkCExtJDIJuTD6/e35XH2PQ0qiTwKLuxrK8Pww9uph
o2pJm/O6nI4NEM4EDlRBL0BTA7U9rFtMi/aS7PGzVwV/DA3GLeTKs6VoVBE/6/5Y
u2EKv6t08wYqss1Fz9C95/BgEwN3+Ne8yUe48J1PZWUYrybAVmtwS1AweWv3tSfn
xi8DXrLsLORmOFiJU3VU0Hy+AMP8+Rkjtlj9EPtEtCP7khIgyV5V1w8c2i67V/K8
bQQ/T1R04El9hRRKcWFF+SW+BvxrszJE1qR7zX6Po3YMG2e8ht1mPs6PYSopEWwm
dRQ6km7f/zC60ntdWYqGs/bw+zm4bjEXNbsiei3MVjQyuraYeVlv+z0idIbj6ryw
qEfutEU8P8QoR6qwz3LSPBtgnpyFOz78UbBFAyKfc261A8XAoeq3gsEwGQD1iKpG
HXJRXneeaOBiaHv+ZEhJ4gKJ60p5iH+3gx5s/cop/+bmEoH4+ZBe2P/Esay0IJ+C
FVqRGJpwi5/eUg2HAPrqnhn3aNYneXxfK05jst/v8Dqp55MNf5SDSlfaRZlRY9sA
75zGzGlhK2fnII7k3aZlStl2f77mv8Jez4vUzO9XODgT2jpG6VUPnATQpwGU6tlS
0LH8w9B2vTejV5Y92tJZrC7y3XzCMR5xi6cVf2ZNCkSsSHPWbvM00O88eC1/UI24
0eOQemz+ppEo1WgJ9VL2t9toauuqQe6SAHnGRa09ZwpqSNOkq6jgfLq0F0wSvnJ+
xSeVEF0LxdW+jp40lLf3IaldF86YpfJcJNjBNtBZCPVfHj18/0KJNBfkmj7dATxb
TCLVB+UKs94leBCJntq+yY/qn0vtSQPovHH1E0cn8jY2IuNFhA8Wcl7wOJYnvmnw
g49AoaQODtBD57uO4djAmDEV0HyQFo2H1vcN1T/QFotIYxC4bh+wBLvfzWgUzNlr
RK5TAQfxUX1VMHhFDoFGlG9sI97WOYmoc5dl5KRgOEtrqBPcAYEP816DcLo+0Ogm
wEZhRvL0u94c16+MtRPJCJd2fxDT61konifgQaEk7RD0V67fn5a8Culj0G5echex
X+d09Cd5RL0dNJC92Izpys2CEwQ6s42vQAPAwm0fOkJ98rFvlBnIxvfTPBE46VwN
iSwWN9crfayIBOKQOT3I35r4EMQv2UpALTVAsxix/Z5x2HDEPypfL9F3IMyUhdk1
BK8du8AVUS7Nu4Z12kCUUtXsWhhbxyBjj39oqgmrtken/AlXtLLVSTeYtREPlDoq
zE7NkRGkMpvXBXiP2q5HvQyahB2z3S4ho2KZ1hKVEj0+HYyCQhhW//Cvk0EqEDiC
fR8x0Sbaz42MrmL7CV/7kOzuOTmKlRILnoTkEx1fJV19B7emUpqv4vRi3BLTJBuo
y5+PyulJ8IH5+SEgjMJcxRbAwCAsTjisNNPDLKt8V/zZg2FBhaxLR/PWcUzH5UnQ
7skpHfBJJJ1RTSZhPErHFs4m+qzBpv1eQ2ZrNB0OascDSlfxMxpw6TmYZA9ai+7x
hR2wURKjzftp8z+QUqCyJtgnHfGeyixjx2lCpBNSIsPiLVdCE5AZNch7bJMCKVM/
7Fpb/XQA79hKttB/weEGMGDa0uTS9gLTjSXYTl4KBPXVDBdmdjOR1QS2eirLuFFY
6K8qjzYxjw+ENwq1pQQ+p6+o0jFcZbWb0o2Pxzbql+yaNwpEEuWNKg3pV/zGPqp7
uy0fktlIVIa+RKleOFaYrGRrEHn3OUdgE2dKxlCAoAg7w+rMGRNzPSvMBQwIabZq
bH2eZbrkSqhAYSYIqpO6IUlKUDnaggiFk+KAk6TOj/k/N2oQA/+iuPzBJxCW4RyD
7R3h4g+PP1MohUkOhaH5O2n44D7L0IfrN5hQ4Au0p53yED162/vWluvK0LCkEcNl
96argjUsFcVNmlHHtscZCEwt1ETXuR4bQoahZhTJA2RB3UKCM0WjYFgUech6zoq0
knZ2iIAHjoa3dMt/kGQAik0zb+ESK10M90l3eY/MSu8X5upcNuSBLrAXyaCZ9KPC
hY9jLxIRwSnoqqE9BslzvLEuo6EjRy3QOXhihlUn+5qa3xz6l4tLcO0CzY6MWIFq
WDwzj9jQWY5V4/8uAXGd2o7T0gvqYe+jvTNDjVD/X/1OdI6oOnB6hX9W2Ldk8TV/
k2CvA6qBYxHTUri2AVTL2a9hQfRdSnU+45wesKDnvw5c81t1ccRmGBFbamGnoZXV
qMsk1VCjjg1yi9wANRqcAEOyOKhTgrp36GX+iJQq+MD/bS/bd9lI2C/yvKmaaHnJ
Y2DEFzvbZMDE4n2TMX0RaYrq8oyOFY8TutTSMyQAYhKTkQsMLM73RnffLXztBdXi
Xc9oXMd7cm2osY8G1xC0bTfEUagev08Iof68DFbICtLVkihcBZPugorwcmWnRsN5
xRqAGVrj6JTIoBXAw1vELMBVbGpbABQOdwt0kThTa3AspH1FYTZ68pxquLwvL2sw
7E/pKD4GP/owGrg1FqoVt24YbJUi/MY/u9sxHBb8AHzZLtl4s31Qz4F8kKONttr4
j3b3DmIC8Aa3zZ8pLXVCk5aF2uQKio7zjdAeyT577KCUxMrG2KtZWIP5E3usEaD/
6PVi8ZZHCIFWmrZFT21vMSB+lCq4OlBYCb0eAqZ+oendzE7zoHxw9qN8bxFjuWAx
0vJSKRi8Pt2g/sVUFq+SZ2q4j5U9baPiMGzu1fgKDxAvnG1SPPD6mvk1RxOqElNX
XN4H/RE18Wrp83WufNY4ed2S9g0Rju08bHXgvje5LSG6qB2cQ7ORbBZv4cLDbye6
Gbl1mMAgy9/6XX7ZvEiOFLQ2oadi3BchB7u3j5m8tFeR2bPLs5EsDA1/cbmOoDt6
Fu0anVJPRiW4gPNlvsaebSf4vZh0QYvqXd1dshwOgo+GzxTyR34ZQZZ39IIyv4P1
1+Fx/S18WEyh3Aq3HDgpDPobwpMzYyNb+WTJfnEq2IPjLXeLitDSGBiBgyYUV5ZO
HU5si+Pwt7GUuAw/tC9PBR5kTukCOW4M7k9WPqO0GBdDsUrS9EMJ8AAhgw6mDhtF
f6YTAKCcgfCrAMAd1Um9SLA2Q6DMqrTcQ9LIEfJ+gdZVtP1jN3leieR7z+z36S12
OSd3MRBG2I4EYSAaQtJvuZDrOnkTrpWNyQ/4kSx2IpzXlR15uhyDhkXQdDmuSnZQ
Lv8GNL2GEtlVq/ENR4Bpyh/ZYuN/Pfl08FM4XaqjtcTQ+sYuae4Rrsf0rJqGIuQO
rtiLW7thHs8VXj8jUKy1SlMufTB0NK964pAwsIuKFTbkwlhRT/gS2O/CH6FVEx4M
+Wtu57m2svSSpu5Q5Wo3ieEQi5wJ5t+INYBc9oidLxKDZWh3rfXuR+pOh6S/5cHv
eiVqgFw3rT6ZT+hRg+wi4px7ccOdjH8YWCTGVETqaU0YZSrukhVUiaqb/j0NGYYP
wVfdQyyDo5ADfNAETNOx/n5A56+rIYp6+PU+e9A0GPsmj+BrsConNh0N2un69mnX
btAn7B0pIjwv/uaf3grx1e88+rJO9NybTGYIzqxAQ+lMVZOUqTFTlp+YTxWiVQL7
p9WOxHpqLHrhh3PEHi2k2OozPKjOrAym65DKTed0G9P99wAaHtv4VGtVVeD12Gpr
ziuTogrC64NHVdH23d3Z9Q52pR6IlBMYpVDku3/kxtqLp0Lp52QbAFX/1T686eSP
XByV0W3hz7b31qTKDCaeiaLvlaTaxx7559JgCLods3AZz+TIkzmWUtiq3/Dnrozf
zgYA9f4RH3QRG3BQahGeGgdAZkACBmIvZVWdmjuwAj2x5U+doJ7ineZ3VSMXrkg0
TNGO5wtfFyD/31/SYNP7H39v7PQgEV9cXwlq49qFdwVceeGOzrgXd5gabPuQPA6K
OBV9I4oAj/9bHVdFAsV9yOouroZvXuJT72po8cP9aVoI5pKvImJC1EUUKMYk5I+v
0H9YaMATO+Huv5onBXb7K2A68ssycNN0K1a1LMVeeYZtZOuNRwNeJwCb9Ya5GMNZ
gbnQGp/iXlbC3CCZ2JrSJA5Hma/hSdu/JRdb6BkFIYDTgCSOBNU0vE0g+PuSiVZu
Tt1VjIuRj7JE3RuthR99yVtlu6+ogfLbWF6PqswZbRtqVqbJea3DczcXUMb+4rNI
rRKM2VSQmdP0CsTcn1ET3I1nt82iLaC85hiadRhid4MoRdDfb2EyKKx0MUpAdbvU
M/WDrOw3woKmHCTN11dhw1hq+h7obsS2ruyHq8DpcSGfwQy3ANOUOPYrorIAQyhw
1vb1M6+IYSlOCUUnabb6XeQd34xkAihdPw4SRRijD2OZUtuSTDXoiKcssVCsWp2d
uuXhJq+OZIQQKLk56w9+ePiyWPJU0vohvPU85XE0XALeWCLj/+Br93aJte8z48xF
ZJPKg4a7xFgmjVdjoD+tb8UMQOtFPbrwsG9r7z3ytDV45Zzn+ffHYESBCH5kyDOj
w6XYSF5DEhEgaJRa2Z+EEnM6zqumbhuxzKUwtfuH1v/n9nM6d3gHZgsgqu4XH0Wd
LEaUUkragDwSZukEkpoGKyZqMmGtT+hGlACn4QITSA/qpl5DQbteLxaX6wUmMSw1
EIod9BOQA2vJOAdSgo9PvaRMwsgJLyf84lxVU1knCYgajCoJvnzFaF47sBeTx9GQ
5yxl3l6JNHOGcD/D9lMvcT1ZLRB8wFX+NmCAGygMOnUpIwqKAb4kS5ff4cImq8FS
Gftds7A8iQyl0c5vlrc/vDEEFSodia1oBWU16d83nV5hqDUdY4GgpbY/RDvmRvkV
W1pdbehpawHUtBJt6d877b7YouIUgGAwh4K01U1dzZf1AywbsDggjb+Z1XyIqtON
ObA4iZ3/GN498D4bc6uosAzvgPAYoYK++BcjVRwXZN5tcfZrQU/p29HNzDlDCefK
ZE4z3ispsdQDgUEWb/rtFtVnB78cuH3HxkyC06IBROUQnVX/kz+ZVmw+Y2hK1xdI
JGmEv9/LHHx09MaCq4MVEZrihts7gSxxrNZ1bl646Ikl5TpKY9efK9rbm32XK3R/
pifM6KeeXF6pGsPd422VWv0E7CKBszOrZccJpHgyTYOgunKkAwGvYDD11Gc7r1R+
u4wFl3IaFyRuxfp8T1+pFOwHPPrNesIH6KiCNV3iUEFnvnw+Bp7saPOkciuOXOxY
nTlX1RvO9etXEpueE73/67ThqyOZHcEO1d+EYU99JqKuMhwUiAtzihebJ57RpFq8
UI2f8Do5njy7Dc5ewxsAQBMTP4svJwdzT4Xihqmo6Gxyo31GRT31jrGor7g0w4y4
FnQY2xOrBoziIDnBTB18Jgxv9FqYfTBHAmT+rqibD+36umdONfhsDp0CGfSzX28u
ZoGu0AonCZpfGWtEn7qFu9MhY9t32FXocohcHPnnCpuWrW9NMxiW4gknMxlDeYEg
OgdYCpkwR5xsJjZA6ll57ilw2pnJiyM6V0lJASe1IpLX3elKG8hjzwY+AHL9IRh0
/GKgJvWq2Ce6pxthX2wUMr67G89L9x4K4tkPe7rQf5AFFG5XI2D9TOIY305bVPI/
PapFb802zbuFVFqGNwPAiy6HMbbZ1PiC036kCk6Ci9UbhGZnA96fZ6hZ5jd7Z/1b
hvokqF2oc9LZvGqvcVLAb1v5Xk8WwPO1GOegOgw87gCxl/Dkt/Ye8jJw/g/YlwEM
/KzE/SuwkjJUgPm7sMXw8+OMbiuCdxxTY1knbEjlm5edE6vK5U2t6i5ofCewCfTx
n4DhX/7PGs3JWPpDfH9m8NVtgnPPrH++wNbb1bdHKTOF80BHLbP0Szg3ad66+9N2
W09iiAdqgLce/P3MBgVrUHohJBGL4DSD49SMfhYGQCJcTiRirl5Cv8X2ZVcoodFz
UC2xKvC1dFfAmkGeQFyZGx5JoAGomDk15ezNXdsNP8lxdx6gAdTM3neH40jd8VGN
SIQ1afIlOKi1CpI1RhBexI6qISMGATB4h+VSeWg+rmf7Ju6TvMdk/UiKLOTaujlq
6vztkppT5b78wsWH3iPClnOoOUxbl2Dc4SLuP8ybuVtrqOFS9I0oq0GECUO8qIJN
hIhRstVNKO9EF+3ku1jh+gVWhhNPLlGejdLy2gX/o/qF4Zx+a5EzES4TTuqkSBdM
WyV0LzkZjMqNlz969oglweDy/YIfgcF2xSNHqntcaLZ/qBGmjvWreujjKFukappJ
Ja+wZkt0sOREr6ix2dbZ98DbuCMOHKl0UAREDXPTAj5EDuluWjgHSMRjLi4d4Y4+
VVWy5OdlLFJjAtW330a403KV56Iv01gyH/UCHNcaZuNDx9eQSMd4japlTLJToEYu
lidqcUURuWoLc6HWXBBGN0Nv0wCBzYDHaF139Fypi5aJMm/ZrGOr5E9agM8YFMJ4
HUWOePEiVQPUtiXIWDrEqQn4cntOSigY+LDzg5ImuaJqYYx1OwyuPgmM5OxFL/GL
iGbGU8rfZO/BtQ2piLjFZISQcnrk4/f73wPHlMg1YDK4urqIopc9kmr5PB94lyoj
S4DPIJ2NzzMGRRVrLcgjU1Au8AoG9a0BPZh7L9nc+mRzi0PBOBWUHFC63HgNdEcq
Mb/HYhbEtnhajXtPMFUwZAkZM0DALCfzYK8oVU9/Ide3ezQrMeCEh1eFyNH6uIVs
shXYJFQNqJI9tHJlluEPP5/l+b5fWsCjQUfXCYZ6VQ67Wuq9jN+pt10dZb/leQeO
D0esRhhhDk5sN0rpeURyKHIBEaBxmeYmZwB6GEB15zuH1aBCHwL+DL23/ubA4Dx/
VbkexY0eHFUIu3CGK1pcfayL1ein2ehnZqJu+b5CXLsoRpUkDhmw98Ry7bvelAoG
m6IElvmYcDns8tlTBrThF/HQAV0OTFIFvNJWTCgmqvjf/vIVk/bH8rzdYFkpPKEW
W1TwPUwrdUGYXyiGJ8WMUoAINrbfaC65F1xXDKs8ppv6bKq2HZxX8FtdZzLQ/lls
bRBjOvmVw20OKs/3API4lxUWD1mHFdiGDxWORz/ugwxlnx1wRBHK/9TtkC8CK9U7
o+7PZtCesmcqV/LAz2GGmknc4WYw2ka2oWktPY2OjRZjUXR93+0snsDwmauwPCXW
Ge0r6u0Ke6EZ2sch4Fmc7S7/U4XaTTrMtdzv9zZxZEpeyXUrct+ANzis0/YSBBaG
Q/bEnuc+G8tVNkfQMEyj+apn3zpCtZTEvjCiDNcc4+8pappCWuJW3LLbk815AApp
UYRWIyY3GycU00qGSWjhegDC8+6vG8YXPBQKtSU3XGGGIcaySna0VuX7K4vgiu3Q
mCacH7R/IT77Rilw2zBP+DVuvQU8Ou9UcV9pmeUkOMqm5N2qaqyv5yhH7tdtjE7o
2sdLBvswD9mSvgvL8hTh3n17ndsDKG91xxAc9ZwXSWM6t61NBRoiE3yMk/UV+/OJ
zmhC8Rs+tZcx9yxsDqikfLnX2VtYcMbSQuAKTNmGAZ6ZsNWBeBg/1o79AbfHJddE
prSbKAigmyiFP6bXAI3tMYc1FENT1CNXAu4zFLsPdOPGRz9ZsYwfbc1L1yb16i2K
p+6Nlr+cjNq478tVDmsBxv9AyForTzgPxBcl6bXjI1W+xFJnXrHXLJ5U2YrF0m7X
jolrEop4IuNVKNTZq9NrQS1LUW0+vCMj4BschpCgyvgjNOmBdXiB0s4SZZWu9Krv
ktoXhDqBxSdAFMy1TsPEsqobUmbhjrVYb1Cvf/fB0KXra3dlGIIhyfsbGKu/SQ20
ujzpRZLEzaxTzbfQXdQRuGQHNeWeYS9fBWHlYsB8mWUH67VDZo8njgcQsoDQ25hX
8kztpMe6+umaTJuX/D7iuO8QA0pHhPd6uijiJb8DnoYUtrA7rMQz27q5OBVNKXCR
PXhuSMTN9LIy03Wm1Iqb2FsUY39J4aJODInPy+9hphtbCjpDl1745Q82QrwbVVgw
AVtEyZYYxoF7kUsTtjCGiEk2iWYNcRx17auqSZOVhTV7pQFmYhZyRGaWfT9r9DQj
/dzRAuMPdzPNBMgzRTTkuGRvVr3WaoddJUlljKVnMX2qWlA296HDnY+p6PPrescF
T5o/lbvsLYjBFxdYZ+00tNPpw3bqnH3wcIMwLS21UBhCTK9NxpR0Rj2Rp0N4ZIse
C5BKnEoACwa8CgOXZcIj7As5KUl7+kBE6scvfBjTiV9zUK+2ikxUAnYbHDdrHKkK
M04jCGF9D2FQMI909k2LUTNVLl1ux2AlR6ggrAWepVrQd61DS3CJaaXBck8YgKt5
fIvWKPPEjuov8oD8ab1EUIXIztk6yfivW3ZpOAsc4+/5vMDWCi4Ijvjvlp1YsIZ+
vtPlVMAYkPc3BSuGbDe3jbNiCw/egOKvO7Nav/XiqV7NF481atj5C2WbRcFVsd37
VqElitC8kwV1CChG1f3qYiK33XHW4J0fgzyqnnyTvc7n4FzBAl0mRMA0xKt3CUKk
b9AAWqjBEfQB2KE5Sw0d+IX4IRyeYX6Gcv+pos99HWeyESyq8D5Cx35wZA0YVIao
ek8txT/maUie80BrbcX7WtFeMbzTqu+wpa6uJESA3hn5MaVmyCB58y8w/2sS1wLy
gxBTFOU07vbaeDV7l6+5K/wBfsJr+B9TiNE0itt6JNV6y/Gn9ZWmtMulx7KPwOIA
lt7FJ6R8S7HLbPLXGCCITshSBuWqborZX1LGm8a2m3QTBHY0xVs6UMF8+eefQDMx
4vducyNdXvygaQharpLjTXvWlsm28SegvND5mnn7p0Lft9cFf1WY3efdVb8xIi1T
8iar+++qoNq69u9dqi9MoaNeDzYrffDPfrulMkjt71mNrgoTZNgZV+IS7qMG/30u
rnB8eh2T/4r4OtTKBK0oa6tOfTMkExcD1sMQyhAAb/IRj+eLYqvjfg3ufatbaWzk
pKdgpqkIGrMN6FLdMJEv0oYwmoJq+DQQzaFCbFDyD7C7hlhz0Xcz2xQhC5Dqj2e8
CSfeKtvLxwgu7sdSX2VlLL2T9z1n0qcBO8ic2eR72rbJJ3n4zZT+6A+kRsMViVox
t1nqDLysZVEKSFhPtKsiwBe+eE0BIfQxnLLS8V8+DGdHwHUQD/yrFa6nZLjGUoNf
xYud5y9PwAnB+OdfcagTLjpgrNwO2Z6f+lKJJq98rFs2HBTbJFoiMfpdbFkMobXm
gs5HoGGMt+4IcsIZcriADpcSMj6p9E3m6uCWMbd8ir1CAKFUK5O3owj6Upe9IHbF
OUPwF64CbHu6W8687mvn/Opl9ZGtUTCHaRE+nqkPB5Ow8+sWFpzRYncS/LsbjbCO
xlLkAcOjyoqbx0O44rNF9Tmfbrgjvs8+Fsx6uAJQ+7ksb/+OBNOweeNqURear5ga
BIksfy4EZPc47NF4XQC1l6GkwpPzd0RmteeEl9MyH+1SzoPTlE/M5zf9z5XkOWft
OCsbXC4+8RJ0Wz099kgp4Bja96AnB7SkWCFjwBzGclowDykiyk07RzJtNVboHhVF
9oY5RQns7iv1Vpdj445Hi4PyUrbsolYWvM+1J6O18WVGbgxtRLSU4zlUQd9tZg9U
wN3pyLLKDNfVV8zLwGoR+WaqIWaOf8zfc4M/kkRz7HDuEIpCMBqW5u4guydBRzfh
Zq6ON7dqzaowlnFV/iqEnaoe6i5WbcF/PUk0NZhu+IsDjvH6D0iDPuwOLJVY+yfF
x46gt6PeVCcHGCNM995dQiGl0pMD5bKUs73fUHV/Mc/xPdY5uItKjiouXfhyu2em
XgkKc7pLaCh0xfQ1XKiIUTzCNAtg6u9H63GIelOx/k0rm32kXpi1xg55IK2ciE6I
D2+cyv7Ewf6dK0A7Mb4hV5O58WgvAgBjSfqa55JCNih1OlA9MkKcy8xMa8d2oFBC
Wy1xr3RKJpF0IMgxH7bsS0KoKe/e5LauJpJ03Hi/XtnGlcaXdN2iJmyYEQXKWbHj
VkHTWwGgZh16JR/EMrIVZOQQHpI9Cn0dNyX2aj96WdYRdRNKilzCSDbTEMCVQbeD
SrfkemNYvJzF0b6cAihQcJ6ro5w/wJ1XQBaSKkAehPmll7DzWcmyUoxn3i9gj/ti
5T/PxdmpwHOmmpp4SuEwPTrgZGNfm25Rn5ODdiVExv0NxS71nq2SkWzlwA8vFvSe
o8GzhpiTF8jB0R+4jzZdvVKDvvwEPrwnKe0MCjrrVwhs8L4P6sZlklrTCi4vjzuJ
vP7G0gjw6EkGbjcV7Jin7ByYS5wca7mATMv8QWvsif8Lw7L7QJIqxdeIYp/eTk1y
v+iaQHH5ZT/uuU0SoBwBfs5sNGIC45oGHU2fGeOwb8+6ItqJnCkFO4kspB70rzOp
5vbX6CYzaDBWz6FTL7DXGiGqM/xezWmFJHwk2baBmLQve7RkpIibVQaW3lflysCb
4j5x4Wn/vCwbScDduT4MfdbndRunkSocSdFIRIzMYOiBLFpLoAS1g+OehYgIQtxx
INWC5a1oMsAHqNTa2Xk+9ZBY9meH34XtvCvDSmwkrtfCZp/ZHAo92RlJnCLKypOd
LaRH13q1R/+sp+G/F2nPqCObGbTYNctnR+52oiSVd+7+V5zvqv9ajFQPbfeDGm4R
blgD0pQubBK7l9k3rVFwqDO8CRD+GWgjRH7TO9ngtdfQJfvuOOvHboO6Igevvvo8
fu/p80TxZyOJ0QFuQ1oZsrQBAed/PoaBMykbqJZlCZ9xc4PE5/y22r14BSz0YdGl
LyOK+vwxQqj65GPC0I1G2QmbM3pL6pch8m+hnWHygmck2phUdhIMebx42x93X5Fr
mX7QJrrW8a3fDVr/i6M4lJDNN6rHPElGFT7td4MN8fDx0nF9bf/SD0W39fkq14r+
5ymBSQTVU0Z5hmew5tPRZ1EB5Hhhm8Wl2RLnfA4gMWh7FsOVcEBc2eibsSEply5y
Uon+Bd9FEea5tkA5orfkHb1WS48oAo1g8G6EtVwFIdvf8BYPKMfDYuB+5RCYh6Id
yBM/74pwU/ItIF5GHizsODygKrN4WlOaDIkExIPwWmg3NhE0FuBojsTzMvLKBjOj
K/dpQ2sbPnY7x8YgNrYg4wyX+m7y37gjKq2/UDVu+vEUVCUvlTUcUVWKWmOt7Nf8
Lco1mD0FnZPWNFf+bzhi60sJq312HJYwcB+NAGI0VrgSuyyDda/3p/fAwrQaVSCS
t5MQF31PVh58XyqHxLk1Psx1gmGaK4WTG75AifYIq55hWp0+iawnPZ+7HNGeN7wW
XPz97cpbrjScp5+4ycbDSLr1BNLoywDSqsCX4z57INy/FhDktNqzl77VC011UZ1L
aNLWPUB/Xypli1b8IPfsvbJJxfg2BD1NGeM/4VDukuPDgSM/7CdIiKaQnUxV1D+N
3A3BLO44i+TZP1+lyXp0h4aLTdI1hM/xD51psinPndZ5f2gB5kx9gJCvuwTjNKga
clX9mbYB5z5ixx1wzaHxRYk8+SJDL/2FOmYV0KyJiSGekg3aLQ0IFkjfuOM68Nm/
HOfCO0aZnqk0M0Gw3z4Ll12HfO3VfEql7onwV2NxqB4m245cWn/NUFoCA4+BzHKX
y0qbuWE4GtvCSMq1enp5MUzStFKhfXJAJtKObWgARpeB9GOQsomfoVIhVlRlCbk8
RgN/VIOdunDvPJId6rp6mbnw1x6oXKSMqHbg9N8jJyGGmDV4mwxP0PiBMApjnY5g
OcBl4ebLsiva/8ArtQdccg/9OlibB8sfazptUaKzdbokgBSdScyFRivdkydCR0+f
qgsyyiqrZ+mJX1f4VFABqKV6jbKNY1f3xWA338AZzdys500mJsoFkLPs9wo1yFzz
Vsjer+47FhUBHFDDFzzo87qd9beUpQmeU3fsyQCgQpiF9pRKMoOK8I2+5G1MsmZj
y1ilq+taDkon04sm3zHu2vD1nnGLmNRulO3ARSjfPC8ihxrxYJnBQ3NnFH43yCo4
qS0LoOqC2TplI6IGIMQgumkICiTP+vODwpTKnRjFgeLuCwDPXG9MfxFaguNYKM0f
5+tJCKWpLfDa9LnvgANpf90zFRESJa4XWKEeswYW/q/uBxTPsC3fKt184bjU5pcb
8GNtcUbsQu/a2mnuNbiyHJQ4Aue35Io5liGnwUGnUY9Ng+EEzF/irFaxN0aR5u1e
LH3sJRzeElDu8C8/0j5q8Tkd7uTsjdSWMlC+bg0k0dqQDopRnfRQvVDwMhHbGFe7
uwlxtcsabMa6/67Xp/TvYAifm4U/9dH6rur0OA0glEfZf14GQsvQjb4T1gPEyuA5
SLNTd//zFboFdOtltxJHnxFl+rRXIl9KocPZxgHVKTajZISuPOBEXmOER7hWSEcC
v8m5ShinADqJMLd0v0Hj2T/pO4FzLHWSp/C2dv+XxAFoJMkprFo/yMFWp7j60Bcz
mbhFx8SEX+8hqf1IunFigkLILJ0550ndSGajbV076xnFpVs+AzlBahv3jGNKhkWh
30InpZA7HzHI3efjFugVlQEwKoocMrutes/CddIUjrcnp9uvQ0kS9mcSqcJpyDgT
1al+KOL8JJm1RymrpxYZnjcxfOY1dSZC7/BcdMKXW8rCcCWks0dNixw4ADctgqUC
b4mItdcsP+UPlyAyqOMZU7DwKN6PEEiAIBMafvQK/u3q1XtLuYXiRh+OXLvu2CTP
7hgXoWJ7m90dbK4Yd/SI6N8uAaZoY1Ob6+com4wOu1P3SZgPZwmHt8RBw3zWMvsy
k/Fgo2jXUj3MdnXAaFlR1mqkihG+U5g+arJalaMyXtAArkx9QSko8/7hGAAglI5O
t02Gs+lFFVdvZTEZSmUa/7dZ1NHGZBGh0pipUvyON01xUjsRjJr2UFDSwAM7/LGW
wDSZyuFh+XtMTLYlGHw5eGvHxsgSXAMoDV9GfvIl7dJTBGFdP/E4iCDXUp4mxUjm
//mw/cywDHQj7SSIpniZ0vFH/vAyBt+Spd167JT5C80XvQu2Rba1LsNKfjfatLMM
q6fEUjqaLj9vYF7ccO0Wgh2QWhkJZ2MpI+YxkMDprtgFNPEHpmNNDunCfb/lhFYj
KpZwCESOOuWyWQl+f9yXHrTMR1wFq3Z7ScmP+m1hC4Mw0AWM7pJzm/fxkYLdnFq6
xkmJDNqOuPlWRBJCT5OZwXdfa8fVbgMSLJBwNEdCY+nO8OUXtn6+gK1SUUS1pEWm
trK5hp29NwRuGzoyph4s/TWKkhUnc/uF2AuHCRemP/cq1VpUEsXxKFiyiYjU4Ifl
sLPFk7n4g9eRkbpBYEyvNhl8qA1n1yyiSzlj66FdHmxAZX1ejMoghE7EVQaa/0mL
TH9G30518a0TO5y3+Et9CEKUXtIgeBgTK+l0ZHP6TG9AYkmodCIixo88y6YkLkzK
PSy3/+4I6X8Sn7RAJRgh/d9yBPwWu0Dj+kH0oT5hvFMxwq3HvBi/CGI/DYRDWRUA
AL5z6RocZ3Q/Wrmqboj7FymKtARaRE70R41oEmUNlAlk6b24c/3NM7MU3kJ76Uaj
gqvEZwxqqqLIZZBmkftHx4L25X3SrKlXHMaG+woXjVN8woX5e89Yomj6KwsKruob
88k2yJKnrb/5JToKbK0X8H4BEeaRORsSnavbJxNmmKKU32qAHXFDTFlyOoUlos5u
SuBd+yzg7rLNTJV4XJcQLe/1mfsZlVH++xt+ijcqrPpJ1sOLmLsFT1XH2PykZamx
w3hGUo8pDvZI0V05h1bBpBOAhaGiCU6kVPuXGjtGr7b2DynYohkmUk+lCMW6rUf+
kic0ginW85KySqCGnwZQK9hRur6+33sc3M43ynCQZe+Az20U6vvPBT8JC2nO7hcK
ttKoxBb/pLqBlkJ9LOe/YxlMAN4Qdrd20/dnVsdAExFuFk9aDJVel8MEpVhh4lFC
ruvR/bJRyKkgCfj6h8bsID3aftdU+PYPjDfIVwpA9OMJ/VyDnGUj7mXyvxJqV2BG
dLxVjzG3J92m5wVC6ycfwJfGZoJjr1wrDHxZJ54U+VKgsAo3tkiM4Jd+J9bpScUm
8TESkeyWG5slmdJDu97rY5RiWX8pYzNW6VEqxEyXCCwoUF6LWlJXoMvEE1kAuUNu
TJmdjI7aWlv8/TY75AV8NzR3q1vBY8r/llDj9rDQ7ZUC9120BZ5gGKd2WpsO+xeS
VZU0mVufj1+9YCG6zlxI/n0lCXxSJbcJWOQne0A7MbYaEzbQ0OEugTYUvDbYCCI0
dZ8IlIEIA72DpHH0k1z6D8zn/tuhEUx4Ca4rsETxrYZ0g2PU7v0/kaxKElFLADSo
DkVF4AVCWpNAnRq8UzHDHdYzWzJakHITNOEyWjN/Q5MwMd0dIPfxoS0e0z0pxRkP
R1+7kBVALn539nD50D4yjNoyVmasN/Op+tPVM+Hzp90bri61jiB8wHF6OvnaTiUY
3hBUqdo4Y41zsM7TxoJTUL2eugfbz/nxrzTAYcyY7msc9LfHygF2Rw2EdNd9vJgk
b3vpvToxFsteOnsFhSaMPaO/g4RSrZqXrbUe3b41tbczQ3sqk0z0nhcTOzfugaO8
p5O2bTCqXxNLwZO/SQR7fYaz7TZhPGWJJNWCgeQxkwA8wafYAt5ecu0WOiy0RYAs
sKRB0/GHHepZ9xLnUcNQfC38kuMeY13mx1+UZaThjnw3VJZuYLuYPWKg9RdoIT0y
7NwvlSOihiAoyJl2gxAQdRT6OZ70ab9QTUOnBEmRpmBjM92/OiIv/6iVDzhUoAC0
zQ76YWo1gyPhTIj33uIqlRXHNtpKZOPPm/Nd15Yq6Wsg/C6EKswU2w3h2wEcw8vF
BHHwQif4/nD41BFZD3my5T6oZJ4vn5Kl8UIlGNbkZoX4jV7Ermbp+KJO/Fim+BlD
OWjGcNXZZc/gTHQKUPON69M22p9ML6m0sS92+tpLtVDgsiH475W9ZyA55+hx3COC
XSshQahZON/5meCo+Ft98MCY82wD0pwzBFgIcaTA9JE/2pb8mGlBM2VM1uDAEwYj
SfuKXqc3EY6r3Gt4uB0YQpuN7IWPyGP1k17ATKl1Uibs15/Tgxj8E+bNo+7hH4H7
3ifHI50Xu7MD/T7/fJEaJLdyYUTTfbdxmu1i7IbJdlI9Ue74yp/+T6l2o4TAPGgP
sM7svKAANa/pKdW1WHe7xCUAzL/1Pg5ndTuycaOdjyg9kiYT79b/1VE4e7JgruXO
LKx+wt7oSOUPQKJFGbgOerBGqiA9aaDxC5xqAm5gzs4+tZmJi5iRuUoqEtUZbRwx
DTJse2YZbIOgyqblIiVz7SJotoqPLb+Q+VmFbSQOF4oL1i7bS2iemGQ0WmfihQhU
vV8S3RqHHjj/dCmbCLGI+2ubxdWNOObz2W66gdjDpCpoEpY7sTiV+dyfWvV3cr48
8SmcwAv2XQNY5uZSMpco2hoE/VVz21s2PFNr17Q+GkrKfXGb9RLTJwBw1n4mR0AK
/vEr9qgY8j//CcCVQXCr952wTwGaZcr7sqUpe2V3p2U6VsxoLetomv5lxu8GJ/11
hdWzwQJguo3HO6j0VHlIcikFNfQsfi+5IsKHVst+J5Ro71JiBKiSXh1+Vzhlobs3
0LFLq3CAJBR99YT9fHpxvqAhtuBSMdTMueE/R69VfBdkjcCTO2Ve6NeLQtHX0GqM
FTcA8IScdt/VX7NjaSmluWBpZoXbIJZ2/T1LLFS80nyWE9pAdOEHzqXGp9b/0DMu
L2bvP8JemHgc2Vulcze1GaZbsmDap2Yq2LJBZ3Kqgcz6KtpU7fsAF/wjtyFooV6d
dLx94TaswmVcu2Z0kVxwpok9MSTUcJsx20BcZCpnLOYhmWOXOrhEt2WAKR56C/vD
AdjdsD4uUYSEHVNftZQGRCLbqbY+AE2fq8fvvqG/eJc05pe8VuzQV0Yik+hVizks
oPFvd4jkXuLsPuMFUqjxtLNIF0BFsJZ2QYcudzhRIJ+CzQ2FI+rhp+DNjc3IP3av
iQ7iXPAVgFTj54fxT6OhJwgXSxL1cjLzLqwSDRWtWd8kK5rHFa7I2aHUDsizClUu
59+pZiUfSmlLxYNkWDALwF1sNDF8HFrIfe7oIZMDolsueU+Xih3kABMnVY2+mCJ1
mABLH4Q/XQeFIKMOU3PSaxoueFsqfAMINhrl+83FZ5Wx2qQFhZ+8BqZ4xKIt3W36
jA3Ae+o0OLb9wYeC75JpXLYZhARNNMOZKsyJ4ebv+O+CGy9fQpTyXsHKAtvVpHfV
i1BETVlVp6/UCsjvBiEXi+9wxVef8fAdh+GkXY3ihg9H1UjBwZ++En5KSvuHNmZa
XLE8Kruvp3RmeGuM8VHv3Jj1/DSk3yFMDqsjIdrwPUNB95wFEd4yYI/rk6UlQLBy
CqgyHgt1AUut97jfjDRHPSjzJTKEPRf01/536Zxl6czeDmXnuy9+E/O9MSTI6uJL
UxNFJ1vXsYplCLurTYTnsKfoVCA8dcqgPtc0vIUqnUKSu3msxFrZguyS87CSYEJL
YAaICjKqC0ei7omxrJZvmOJYxMxTbaaprDM9RebTT6CaGC1Un6yLBkRSzZ+DT1HY
/zQV0ZRpxTn8uTYJfOYjoqVS+LcuKR4aH3RnEY2fG/sJeZlcX0wAmjpUFav/kI6G
a72L1QQV053MeeJg1nviv79xcf+7ILHZ4I2M15HLOiQdXlBcW2rLdy8ElLNc8uxn
3DZjdHS1lsXC3EYFpB94yqdNZx35oFT27anpneL/dcQBaNgThvswlBbiieGGoflA
G3KWQRaqbYBL5WnEl/gdpSNO6ULCQmJ54HhmZN69UoK7Zdr2fs2v8zUmG2ZY4NnE
N2Jr2oyQetgCT/1XXtXcACdLHsZ0hd1wScUExk6BTjJo2THj3UkE5xI5hapV9Xoz
HuE4ncqNhE10xT93b94s+kg6NsDfLwfp94UCDiOovKjwMrM66MYQOo5FKqsIIUKG
GTo9gwZLJOTqHGSBdhmREr5e10Giv0H4ktzS9TEiTSzaeqjbr6oUe6mrnPTE4FQM
CPNLKThFu24bdQ+NgjtzEWSvVFNzFrTg3JAxvZCG6QfyscIfEuxw06Q+eS0/qvgO
g3+ipRBctj84N+Vs5mvxYWyr5GSyn+NrP5i4iLx1LnIpv9/5136aN9Acqd0gFEiS
3vAWgwyDLRWyN2H/oCEYpLxSBqoL6uLNi3VLXMZGo19YT1dHRDZaLRgOdrVcMsav
3Tqa3qmSPjrH42LMQ9uUsEucdihBAef14Ux65+RXZBuas2GRT0ZH+0cAxDE8t6QE
+5wyMJZ5beJMdQgZjp3LWrnRpvrbAKtHtSfG7IdFCPHGu/V5/RiHUWiXNwWcQIoa
hhquP7PyBSi5tL/Jzui2eF3VWXrSVTs5w/NDVxxzbvL2+nii/C92+VAdn99hzMQr
qbMz+Lq0noRN+/9U6AbcoKsI1WgjeBU/5YMwWXHYXNG7w2kiKSX25qlABR/eW9tx
yuX+wm7zoTnkfIPQfL4fLR6XwqhlDOM+kifcQI9QquNLFpfXZASKcC8UPB+V/zE+
OLv5IPivo/o8avL71sd9NFvlMmifYWmraGWKJeRpWgRrTB8HwQc4e69pmAAmsGLE
yuykVK6yQRrlOlifbX5uJoYM5z/S1pupLHD/pIILy/RfPnlEhWrqYuC9pv625flR
QSwlrsZy0BCmmc/Bg/ArHQeV/wlSoJogUPRO7ozmcXN2eenAOrLUhFnh6kkzHoay
TJKAjqzKnKAMsqJ0Ya3AMMAkbkyQs9V1egaIPHDv6mJTYkO8sFwvJMXS1oAwuE+S
yyPJXnGOB2aoECzqCA6YftmwEJRUyxDaeBk3HJ3vz7t+U4kjvrIzjGxFtaDm9S2m
XCo02koDpjPCH8LsUdij4/zFaSW/8s8H/HyhlOCCrtYktzjVLrvyEX29QPkQLg7k
vZGOZ0A7dlvt99YuotT7of97xgn0nmIXkS3JyNBoGQIK0IbxjvIahgftJ64YNebv
qFlbtm5D5+14wRo3ifF3Id5529ruj6vysR44jLp+q9EoaBpbK4BETYOpfyCb4ytA
edW3CkCZlJhQLpNms5763GGl9+fhVD7oQk8nzQiVd/IHG5H143L9iFeuzmISBit0
Re8ppf3yUf/G0kZs1CROkCanNr7k16egzk7LpBkA+unfsBxT/sO0NygxH70itnW5
4nNRb9ZdIyqEPeikW0RCqMVqVEogqi4Yt3fHbQj3ts2XP10iqwJoBNdVcnxrYqwn
+FsSaaYRH/5/Ly3K2Smm5RDE8ZsqPpbHg6N+NtxPKAyrf72WDwyLA0k7zIn+Y3xU
+nMCqfGvAvKtINo9sIG5DukKRxhyrp+/wUMkLw2n0w1kpqUKoCxwGXRbO1+Qq7BV
9iDZ6RoLs0sqYzQqRln3vDgolU1nfDEkn9tkmzf3wylp97YqUBT9KIHOxELC2iqM
sAjLZiw/NPlZdcWQGgLSmEMtCT784+QKsdocLXWeUwaS64hFs9XV/FoYXa8vRKdB
wDSQbYqTYnsa1tucAxjyTorwsnWq0XheXKHjfG+8NPJ/3VHxQSqERmg0LH+Pmx8P
RGA7DIXeV7+vKQcp25HFlqqtkO87Ellf0pL8bvw95N/GUAs+KxoWNE2xtslu+SYs
hyHk+Phy58B/Y72MobsQgb/++BI/oSKpL315wtrzYVWgUyJmZlTM2ITXAqu3ZUks
uXUJfgCArFNwVlxvD1dOSsZDFDfFNvWGYMVSh1LSmpUqtt5WKZYrRjKl5auWIB6/
LskbqKlGZLApoPG9L96N9MSLag9UbFWcLljA2ZFMIwN31k1k1LWO7rH3evckM18/
np1qjrz1ftzYCBvQ8haNk+VwLndR39UzRyymxUBUAGOkfJgJdsXRns9HAlba6NwA
mI/mc3hwPixdDQivx+6T8tcZNMOBal5DFovkufHIz5GjLhJwSqsrdrpGV5Ydliur
JJzrjfPvYP82PjIkXq1etEr1WC5FoKWEalPi+vBJrRv9lFpu2H7IsjHX/70CuZJH
3IckaIZlj4Z3RRKTCqbAhDJew+1TZU9YleHpe9wYQAg8mjvJv2o+vn/K3B93w1W+
GP1ZGSQnSTXoArafZC6MCWFgWXNw73elhwVYSc1vYAHAr2zdAN8bQQXKMGk8T5J+
B9WGbMQ8vjOBnIXBYlxXyZWsd5hxArmT3vGokSsSnlvqQhGVNym0AKG51R1WciaV
3K0UGSUJfMXyxh5l4yv2u4lBUy4vyzNPhIQPmbxM15++eUabxAzietjawlihyfgo
XM9DM7l2QXUjszUI+aoXJqOw7Su4xzhG/eyIjkSuikywbERF2UQJJ5spLMFXX0Qi
9OcWQ7M11e5FG0KThe5hjreEvqHKrvtshLrEV3NoxaZVGKfGIzy/mdNwcE8MBCfg
IyrRT0wWyhaaqMmlGBmE3+TxkMMhAXx5yfhY4w2AQtmCUm7K7UGCvagFzzLF4op6
ckGcHWthkCnpnXBqF9zhOPHOXya1a7+c363NuET9cFOaEGO4u251/ZSqnOAuBAVh
7IB73rpFysIaEb/mKp5ODfscMMqrXDJhkyf3bDBno69w7fp4TLBswRyqLxZSQu4n
4y6yAwxO6OKq/M3DwHPogSau6eODWpXt3Uj6ZkrnLaGYJdjwMbJyA22GlItQ3Wji
fmKWxXks6ay0KhCBLkFttolLkL3Cnewy7SfEdzltq2iZHyC8LmYuhbAG1sDZrNbq
YwZaupuxhim7nS1R/vGS57jrR3tvYXWWLR1cZqmxhNnpzK3zOYQUazwZi9J6fDEw
J8ttOodOckCp512OYNW2itHtUJGemzeR4gqljUQtBQ71sAjL+r9TLJ1xp5WRlqq1
Dyojx1eCN6vVhWQERUXsG3Gw91nWb62a3G+D1gB8J7A4Nb84U/gVILMGlU/vzxAr
fljf54U15QO7g7vlotcYSiv4TKPKEA7v/qlsHAeGxwxE3UBYV303HuiLZrBaNyBj
JGtfXqPmRftWmBZJJ8/CnaBXMzlfY0APbThkdICoIf2lE2SG2F6tU8Wpd19Wa3Dg
1bnL0MR2C8kh53lqo9LINNZTydE8q+YmDhihbbgSpeegwOGcn2zwjLs/qK1xic4u
oJwqZNAoJFEx54prIFCsR3kgE+UkF38NBhR4Bdf5k45qN5/1ZHNn7/VwwTehtSkA
3GaGEMxcTgCM1sCCezRmzhNPUC8xRQ1JSZkk04HO2/nSxdKUCH1iKcVhcw3EBgAx
Oqss/iSiZsp8BKFYRov+OzEHuG3YCT5i7y0xNiLPZ8A5xaOA6iqjg2RtdUAOOIkn
z7+Qm/28+IobEuVzqciBv706aJm9Zq0NdzAMMiTujW3pzXKcR+CC4IgcTdWoy/nQ
J+kzH2EZkRHXlxJ0r5maDoiRK7WUsRaYfWH4nYsTxdpDBW7W9ePuvU5FcOpOWGnj
7ntLEfciSxxI+W0oYJYBmR3RAsVrcwFqD9qE1Pr5Kv8T41Sch/e+LSWz/GDIx1bk
NEAh3FN2A/v5Sv7LGiFkaNOe1dyHQ6AEaj6kRyLktTxWGjVGGoJkDXasuC76iHan
8dq68UNv0dx+4WIqj3Jgrd0scq5t7VB/3fo3SFIZn7LnTN85h+Nl8WvWXB//4KGs
ek2LQ/EMu56MytMxBw+2r7+RVrXtNDuCFZh8PTE7+8Kl10NhCXT2ZxJWa7RLfDvJ
tH5Wkfsr81Mz9iJjwQZHygqoiGUnJXh8wLH/7cjeaq035GxT1lIn6Zg0n6M3xd9t
2xvwI6hawVZItSq3pcMG93T8w2TfxIwGQF7p3ja4lIzUsTZlu7LE6pmcE5U4ytOf
uHV7xI3Cb3mQe84PMxH+Wph14Up6fINYPQrmSlwSqPFqVwb/20GKuoLiNNaD0w0I
2ITNE1fWLuGAH1y8I+Nfb/jKpbY0QMxOm5FA99Mz2faCsQjIgSzWnqQRKHa3d3T3
6Pf7c5LPpr/JXSTEI3MHU+O0/cMjlPDbGvPaI876SpGDgltR4AMmxK5wLSzSTn0Z
x7CiXpZ0Py/qt1d/GW1ysRU83OLYvmZGnQkDPDGl2xFfls37C/SRdVo6FT98kay2
RkhAWr/75lRfG5aowtNyVkzfrYVxFLGoq88SXsvvrfe2Vu6wdqoybwL8fJHkWvdI
QAh0MpwowYjSaM1IdgA42P8C725dDiv+seprAQ7sKjlhRXcE2ioHhG0LTDCLXWsN
g4nVcWqi/0tuoPk4tHoKoJ4/QdA99ArKcEGTUkR2xGfr5eq40hz6nQuKF1/H7DrN
SGPJcTIxYRSpzOnmWKVH9Th5LKQVS63buk3g4hpHJYCNfGAotm6+vFKEPVa0IuYP
81tyk+uAH51vCt0rSVafzaN0wDj7Rg2szwXIhCQDoG4rZnl+88iEIrB4ugCE7EAa
j4NC+ATGWLTIhBocMpCyDcAbylpyv9Go3GjVP5Z/VrfkdN7IWDeZEEjUMf9lmvEl
W0+9m3GYMye0MvReKYjYIECorrq5Bth+zSi10xy6klAXq6rr9Z3SBWlRaZY+7znK
DtQrk/EZnMV6lE7kCaQQHi3o7b9fC55+0VJABSXdaB5DgxJtefoHUf6lE1XQ975T
835E/rWhCZUmKFBpW8uo+VT/tH98hPJontOctx6dSJww9axlICOqkeFxpJfNoYPc
ZEbmgalRHNywMTfBcS3PDrdgpQAJ9C+CoOan5FZfBV8ONgRDpHTWq/CwIAdl2Lo6
JH1JnVifupGoZMvQrukW3VNhSR1SBbS3raUzApGwP7cctiAIG8oCw7cJnvpm7FfQ
wgK7nx9MMZNZP5FutJx57IrCDNTAontrPYIePUZclSLsv762ZaEOGQ2DyTfs/NZM
PBJw7T44iBdIJhZnpSX9w9wgCLobhGuGXOf5Yzf24ZnCQvOZe1a5DxuwzX/HAdKJ
jd5I09an31Nm4yIXEL83Sn2KgXGVgilGVGlPlEv7xBmvV2egFCaCETqT7e2XobHy
KLpRJbtX2SRRB7/kvnCG9tm9u2EmyvRRVqbWeKaVhi1SGNRSPlP5z+TkZuOwzLA2
L4gU3npf2WodDUrQjmzSnZ1RGqXYkeLo7xBABqqSLFWbTxOBzBXYu8kBZRWxJYUW
0nXbmWqmRqhYtcToL/HCD8zlaKr7z8b4stUCkZJdLYtRYoJTNNj1LfBFxu/7BmTI
oSa/zim1Xvyy0LEcHB0ZPo5Y0IGhdpftbRQF324yflf2XDnlTTJ/T5tdc4qGQx4N
w9PXMY6uC31TbmVK4dj2rZR6NO4OJbPVqHrIFY96v5zZ3lUxXsMOicAOZ0KjJmuJ
jQ6mku/iR1/43O0HeNaDCqHQ4uhFlX9srjTybp11dJbEYMapdGyVRXph8KKfC8dZ
5F/n8vd3Jfgi3jFQ1X1/GGOpCVnNXFopswcZmpKSVdIncg3K+T6i5Yhm3vIiHfRS
VgXfaawMWaFIcE9AHj6ZoSMConTlQupuMp4+v+jDiBB55FyUo8YJQMqhsGKODzTh
P2a1rf/rgYka/3JApOpwQTpmgX199frIEFHHjy8bweR7QBOFa/mHQzGDBsZZfdEp
T5AzHBZnIf1Hd659tJRU90HEcVw4LQEfmju8Mg/kePpqDHJiIHJWJkjPF29+Shqn
3E3qes1z3bv8iw/M6ExKSR3dAerMutvdvcG0Lf/HYzksxfPT1/wX5nSPbn4MSSN8
1JzLHV0XhxDtDEy/fZGg+LG0hzMmcPbx9sC+ijIfK1WBXUyaIkr7duDouYjBh1GB
QYag1uKmNJc0t6H2EPSINAA0PmwGbRfs9Y34O/oxYlPBoi067iasKzBxFwE+2snr
R2eBqsVmfK732LRaoiAfThkOPPQFTAO9En4OXIAV6id8tnShqIKaZox7kW9l41fN
TI5ZVD3coM7IdwttFyc+lRWdbyOxcg8ubZrNlu1TZAxk+5Fc3I7fdNr9TW4Y96oP
AHHIhT0VI+G8cifEuxq9bmIU3vIw4fQdav22ktXEJJk9HMU7RkWcy1Mi9DEMqSRR
h/N3fKmH9FFIjbCCbgV0DsnvYo6D4rBAUG2CMibu51Bl/kTguJybetXY0oxsWRgy
6DrVelE45dikbOqLb98MLIPPpmhRO85ZfKzvIF8X3A8eNH83bwKrUq7Mi18y8zo8
PARGGsPbn1u+AxsLfbDvEGBWks4xDUFuq2fd7e2uW+LZKQH8JlSvQ3CwXjM9E56+
MLljw5podfmMJ728Qvs0+4LG8yzFq0rrpGRZgcx5oFDc7Hf3brn4R9jam10nfoIO
5ahvv1/KzOD5aIVQfbKjH7FGDgkXddgq07YfnD8L3SD0zqkFhTi5gv9X63juYFGT
QJQJkN0DKBCAee44e2nfdA/yIJrM0ltTmx06KF8sf58XDcisJCZAxe4qG2+nZdZb
Q97sMBBy8x9+xs1/icS3LLbvecNpC43x6hV28EedbNBmO6rdIrUP0IxYEZBSKjrM
VbMx3Xs2ZkeDLtAFcxn1SDENUntha5opNnK2vQVSPD+Q6dwSID4b9XdYxPM0QpHG
xKNxIQaZoiTLK6vBSur2WL1hSakIJ9xX9SI+R/5V+ltcT1N+IeG9ozmvAvyzodko
nWveAv1Wufh2/x0bZHBKLOYzxuCb216URCJMtIRxouAQk+lEGDejvhNhvwm4JBm8
tVIBocBsBl16atk8iIljLuKckrSSNVRCWWBMy5araSEXP06ny9DIJW2K+hCpr8lY
m3HNs3FWA/+woY3tNoLbfhjyuyC+eYEY1w7wR90MzjwIQBEYVy3+2cYIwmt8UOld
ZFkoQNakjE7ixQDGasJ1OuG9uIgbjeSAWLpZSZO3/9qtP3Ttun9V3O7BcYQXezZS
Mj82/EaKDd6xj/W5xl/RIUgGp2Fd7O8Fz5ToPTTh/9RCi6jKAVwPSOR2SKziF1nG
hDsOqig93PtS5O6mef2FPCBSvw9P5X7lM99XckIPqNb2ZIeGKniAvbsnjYQ5IQHd
Aj2UzcdHBn2UiC4DkElyYHNrcbv1mrOzkgYbi3M+bZrtDDRktrkvwOIWWqTDHO8r
Y6oiLwosb8F03vlGd9yBSBh4hnTNy5LJr0fH4sWFL0D9c4DZuK/HjT127hosajZI
KLn9O3kxk1xUN4XjDi0+nSp6WzLaxVb3ABaxF04Y+SzBSnAS+ZxP8g0Op+rOazH+
aSE3UaVFtDHSsISzQNkP1hq97UuzEgDiGdSdWYhVPCInK7diovOTPjJTvdzV4H92
1k8bDgBAg6dg1aGOEA60S+y0eEChbzTHdHgWPfoTD9OiDAxa/hyMa0DrO1VMMMJJ
q82NTuWXWqlp1lML4FmQ2g4vbm6nsfUYdx4d9wiEaTl/vyWCKQNosoDvngnxbuF6
tkO5D3ggOZEfw8LbL/sPwxVi+he6oOFPbxQZ/tfQp736eLtsO8eoEe76nfcDQC/A
PWkt4AEr5OUGXqMeihWtsXJQMNlpZEo7EGT9GiUn6ay9MgSinpUxd/STd5rmqZkq
K+5zj4E5KDbqg2FsOJ6d1UrHgBo66bMbiYrCxY3AT6blxqRa5S+QvH0hHssSmbmy
L1FVE7squS2R+eiqklu7lJKvnwWTJrzPUGWmW4mecfmzEo6dSwpvqbOJw6GgvkXo
mHuH70Exi6K+OLKsiWOYrudsT3TQqHGJsFOnx1A48S/s9oTyIYUVurlhq0YLs2IW
EmotyFO6s+Q6Y7eu+wFjMGRgl/55ak/c4fj5oJGmeQsQIY8YEOrpu/0iqZ5uEs5J
G9qfqM2S8t9ksfFER/p/k7mfPWmxSRpx5eVA9wAGWFIaVJH5GRRS4Uhy3CdJCgw+
v8/TLIuxR4WZrIjkE2nHen4jC8Qam91bhsZGZagcGL7ZrUsJjNioLqQ1KyLzlOym
Al4kCb4z0nYwVSOIJ9SrvAM654t3ceQWVUHy5hYbhJFstJtL6nuKEz+2VXnxxYcf
XUUboU4DBAYupY4VERRTnH5eMJxf4BtdzCAYt3JnfJPbBM8IWhCWPHaX69/2+2kQ
cjlbc8ysSZOpCMZoIh5d3v0J2Lv2DURICpJmEyUXYxQKgJ5kn/CG1F49QcqA3/HM
VWwy0VIBTzd9a0kk1w0MvcE2DBR0/A0U7pjUYlpqyLtDie0dN4BChiuhRJlOK8K2
MtFFKRhAiw+5TlYzwuRdo1nnqAFEWgtfjOj/V5blq+8mBymbJTBiOGx+URHezuY3
8x1gOeyocAugCBWBFoE+Mr5RTPdT2fMNV9+xCNxh+S47NXq2KX7Hvl9rad1zZZJA
Lm7kknPVijPLyqywKUBwgNUl0keXob40LHhCMpKVfBAhc3JPz0tUIsnjPtQUYQm1
asKjVUwijbungpxfdNBRV60Q83sPE7xxOC98rYdZ0t6oiPxoskazd7AX+FaHzW2H
X1HbFRPEkRXtJ2mvxCuC11sSFIqSD+D2idJOKexqd3yYC4t/5WYmHiFnpqKpECcs
YRv0y76xvI+NUOTvkaPiNrAsmVsmRZvWLjIkme+fm3pfBYqYUICuazrXHSmXyAlu
eMGCrIVs2Wf20zrCw5HaLwWHEaQOag9Ra48V4AFzbSw26KwWpFyE+xLH8kmtgQBU
EWA4O7aHG45tbWTNPM6vhMn1bjqukGo4Z0Pq3FjWb9Ex7jerSS7vf4tiR6CYaCtl
haQqpam4m2sWXvpkC3LR0rZ/cHaOi+E1zExpo6Fzf3O/FGHyngZm+bYWE9TFO3at
Klu6iUvhg/260m8zEZJpT7xZqpaebXtf7QfTfrfKM6DX5UF3aOvoFbHkmOKYTe8N
Js3fIVkw9ly+7ric1mC0CDGgZ+ikifZ1taru+5+gUY2jc2VOxhogj5PEF2dgFwlo
7lvhu7l0ZZXP2mKd1xw6HmhBEOuGZIGu46oZOxE51LUn0ONCTrIH0n1hqJdMRz7R
quaiFVqyIH1FcxUSf/lPp5GKP+P88bNIZ2Ta4oaSfNDmaIdGGo28eFWmXpR7cbKq
Gb69Dn/dYXhjNTfef8jLRMR2vDuJyseTiXl4c1PsenzbpYJrGtOidPSLck1R51yi
Jcx5UnFoZUq5e7l+EEfoUssZOxpk+zMCslmJOZCd9YcPFOS7ZjdgzTiebqTTYiQx
DAU97bFPfHXB5mbqb2fLU5BMnNBGALyTS5pU6ebrqVWfDowegpvXUvYWk2y+zUuf
RDk2JyYdsAFG87TrE/PqMHvMltTiGC9FcGcWkY11f1GH2TZoQhUAPJRWbUmvgst1
vH6y88aCmPwIIuKriVSpJDsJHHKqwaTuYTTXk+wkNRAoupGnp5o5yWqig3S0THeY
4asbl4ITmrgr8KW4UaAjCQzg7ptm7ed2eLUUk3UxZUZu+nJI/Znnl8/kJ4C/eqxm
onCUXA+X0uIZoNMMEl52Xb8TLmC4pnQl7nTQLnG8Ooi6Tl4odiL1ZWeDShEPNuat
POEdKxCLr5Ju8aSz8p6hB1ig2q2cobHhsQ4Wv64Zhdfy9AzwmFt5jk3CkJIOHUiw
prAbowfeaMKy0XC68BoKRChLl8Onnd6Mpa+FU/4wQj1lEkjmgqzuqB1lFI5x7+VD
ri/PJmd+Kr/6gOr3ax1EIab+UmbZ/9JNtLyuKiNCuhal7uc+viatsK+2Fx6iiXw8
sMWvSEZU6mphEMtv4yiN7HzxIsvuRCvvplaqG4C73E63daOnf9HgiRMgrdC0TJKp
8J1dCqBz92qaGPFoEnHrgKswR8fO9lLLDtVQsm04cqnivjwyKAux5cHDpS48wpCY
u5SmWeygTg7An1UhKWN/uGJX1uLACbkTMh6uKZWPPpnC9Wd+TyggxSWmkeggsyga
tNLq780whwlHkw7T0pWvBCWJtx2FhGvstNRvnHOzVpLslFWC05TJafUr+DswrOAk
qqIzFwwD934BxtW6gqgnY87MCqb9N/RlEgQgFIdTNhlBB5bfOq5NIIKHMdy1wYNC
/e00XY5/iTXUtqmW24RqT+pvXUDshvYit8MHhsr3wqei50OiX/D3vNAmYfmIERZs
ytyx789hv0hw5UpDQb5IpTE1b6maRDV9aZRecLiRjXkbvcF04POYDz3B49jLhlZL
qsUox8wV8LFWBi2rc29sqtsFwt15PnimMBjnZFOc4q0ggJGoPUG6oA8W8ehwVCMw
MpklzZWzWTZGBm2Rg3UF5pnPnBaE6zSDPfIHEfUQtJYpTRIspdKhT9YOW5wQu/qH
o87GzQJ91NA9wVcMaostEmhVBqjE4y26gnoMBkMbZGkcuGdU5VLodBqWVwq2cjys
iyf/vjcVUkIXX+he1qgtAyfFevHEZBpQ8uPjQsZ8+B9LHTLq2vKwNbVH2wApQXpZ
O6CZWHIf+4jUDjw+S92qYwjhNK50XT1ibMzfb8QCtweM0pfYo8JhajR2VTPiJe2+
A76xnXy2tTFDpDwtxEFBdeo/zFu2GGuEYqzsK6QrJIukNPYXTDREjZI7yl/ozADO
cidmKn5Iy55XnL8SfKKr9UkC1LZcbIYfLwn61i5/HgEIrk2j2VHo/ELYZjb1TTQB
Sh+y7UjxKMH6xmf3fFRt1LLRykgALvxxdCHchNDVTJ6GEqUTCSwfEeeMnjRGNNuR
k/V0t+MTePcmEQDb7xKHw39z/PvAqL0A1jBMGPaOrPjaUcYEK6P5SYkCPkw57X/h
A94SSGxfWVhzU+IMaPLNsJj1I4/BP7ZZM7P3k2RwMo512wWeNbAoU9zF6D8Hd53j
n2sdyoeajxqDOxRE2XWVbsa8Ji6bvfIa1D6MvvEGNA28VtVFZQPMno1H8IE6zX9k
uezg/RuL/eu/b7qsS1yHuX8Y8a/38e7h1H6CTSikI0m7DDzdMLUjrGIbp/cAmS6w
X45jNjMI29/BbODB2UdbOcim72tN7wc7PQSfzGAzLb3sbqBCbDhbrgUUVz5QSPLr
XSkuchK1LMOPpCQogaCGFNjMgBU7qx56dPsk5KUvyQPN/CFsMGn0Im+Uf2Jjp64O
iLzLno5tqiqnBeiQ50WFuMuOsts8he3sE4lrMjMLi8S7JHpseq4YSvlW2+vF/rvp
DhEIkX4ycro8w2wwaAuqkdMzvrrK7c1F7reW81cq4BtOHfIx0X0K11V1jTNyLtOk
z3CZxFqX+UV4mfJXzgzQkXZ6Kaz3ToHHQQYQs9KdSj6w/WA+1PbwXitATB8y3mwa
TAgGOzXGj17BPtqBnstoYQUD55PamYVRtRhuEwOm4jriLsJbfInXKqVnQk1RDSRm
tNlWwg5H8iyWmxAQ6YvahI+dROmhA2V0My7UVtniwvkpcx7BkIEOYWDhYdipIRh0
3amO/m3z/NUXdkvve19E3y8J/h3hdcBIRqlf9BjvCXX6lbRs0souczKeFw1Kp74h
FrBBkZt4cga91AquLf40TU9Z0KFFoVV9h7htrcpV7y/s2Tyi1fGxmKPnF1rXrNVX
B3ttmKGWTNm4kOrlUm+3kPeHrJwIxSsHQEYwx4G1WZrbkCU4NhvbYXkwG+iTPpgR
WZeJbl66Qp7lfDwpDwvxWBu7s0osD6h8zQvrcutA5fylyfQMCSxqF1kprNQu+zkd
E4hmK1orXw0X66Lt70y2kkdbspVwigyl8vTi/RS4gUI6vT3PLtCt4uELRH4cBeYA
fokl+pKzWal1LXyd4U+jHvaVlXyifkD0j/ci9gAcFZnH8JMQebqcGBBfc8jrQZz7
GbNtzok+SdBOpOgMtxb+zQjdDTkuROB+TMakfWEljOUqvH66SiklMvlWnFzUMp4i
v/uzHxzdYxeJQuPVrRoU2yXRTaR/g0bf0N6w5Oh2Me2al332P4KN7Rx2WmUj6k2I
eva/elCFDjdzuTOaCFxegSDMdJcBnVKiSP1uc2pc++wqtK7nauCakhOeivJBLV0G
Dz6kbCAPKVgJQ7CL2UgDwvhxrYJvUZXgIRDDJ1b7lRaoV6VGQiO2rKpUQYq0wdkq
+96/t4ajW6txJyHaQNGBNH+4ml0DzjQliydTSpf066b0C5e5ofEbl4Roqv8+qFFG
WrBJNtZjqx4hsI8D9iBYGPpEXaQ+QK3Z0KS3uGGrEWUItGbUQXGJSlM77ZOke/0m
zKrYtN4kjwm9MCihQCRJ8vRHuI0Qo2rk4E033AWFCSPLoq/Jylxm2QkeDv29YYlf
wDGd3yg9MbWOmozdV3anh//cuA7opFzidfM9ssN9dHqjiZ3vXNS9YWI2izytmEke
cI7A8ryc+NAHrb0aO8u/4QVgMri2W9tyZHO4uVNYtjG3Tm41VV8UEveU+C5sRIGR
Uy03s0EXUBVAJvmAxpvJBLlLDVfRxGF4AcdNTD2C/fYbc/f73HiWoMOSwo+80gDy
Bb6Twt1AjI7Zp6hJIbr2e5mHMX+2ePLvMCO2GiWE/lei4N+cMuNVPiUAjnJZNa51
n/Nk4zq3pAKtesKaAd1GGmqfmRlPEpEr+01xFF0S4MEwVGOzQvolln82aLQAQHdB
h9NmgzdQYQzcM88+dgaRA6JBu7V4m0dZDd+ZkL+FQAe3l7xOoB9mK9IqOLp+n4vD
1dK+6WmjUO601IfOy1EjBmH1QOXo+qbMsCV8ufKczY/uL0K9xWdsPWoib93yZE00
TBNMGuyvYXMVMdEm9hAT5teB0nEXlZiGdRcC8tELpUtqqKkJM42F/n3hSR+YyAzg
sbcVRNNwYmPGGI6XMbkEsZYk8dBfUDrt3SoS4Yg2UzaLsOroqMnkDEXrQ1osbK6T
TsvT4Hn76s+J5SD8p3jOdvpNgZcwYncmVjhiPRoCDWCYBe1PubGEKOrnGVkul948
g8Pc5leMz+ziyrmhSH+7eEL1lcHwhajUTKHQ4DUgj3CdhkUp0QIRRFodqfXvs7/n
WVuTf5vbKSuPshXXyHT3JIt8xK5FiwIH2ti5B3MCG0G915t6PTabKQksdojJFudN
aNQq5wBEv8W8cqTVyVt0NrUU/jqFoRdzQAxjQ1jVwNBmWfyjCpYkAdoJQPU1b0Vv
kQdTMdYnQWieEC1b6ADUrC5LDx4gq3zlcacv84Hs2m/MUoBpDTsNrqzU2gDIgA7r
TE5Z3RGFdeQ7kyuQnOYyQfO6RfxDubxmRDAIIsUmwfA2rNnW4iBOKIzZEWK8EzId
9+pXKbnJ0pHvuPLKegcEU2PjJHTxzcV1gj33WF4LBArSrPm58mHCl1UyEjennl0L
klbA30HUixH2C6BZ8dDYPuPxAc1uPQ0rz7yJBuHI9QbPSFOcbZ9KrmXmzUSACAtJ
y4cSSgbW0gIJs4HXsDMT/5ma7MdAksQy5Pb91y62Cc0/QdXHlMjWxozTYnnK5Tqm
o1SWq3fEGnUgJ1KHJvPmVRMO2kEwAhclrdZlDPThGeHGbMvCPqWcq3JPGnOed+5s
bEYaoK8M2H6uZ+KkQgXiBXpG9IStnu5qnFTsQUCkqaoYh9kK2KmcDOTnGeRFDDpw
qtKkFurHtCjFZ/+n8ttZdGHRbfwqjrLTHwk8A+WChkSMtqfauj+UKuA01bL6E+yJ
Sb0ttbYKrzcKUdfuPiO03gmNC30N4+eqByJNvertET66JQ1n8ifMyvjLG031P9xG
dzBHfYecA746jSyhQ42aDFizMgSFVRMmrJ8tcPAtKTtjDSsY2mAuNLtDtC5lWu5S
6qa6WwK5up3fFfx8ZFEBMXh3nIJVFwXPLMkzcXs0CY4gdHx98bAd6b5AL/llqdYk
ggY7mnyUH1yyZVBK+SxzAlc56ZwGxlZUnYh2ICmHVkpy3AAX/ZhkaO5QJ8/968m8
QNtqChbmev99TIqXNL7tXXM56Zf+SoE+lsQpYNUO+AQUvwJHzYwU3+geWwr8IZB5
fF1bumcNc1fCbuu1/b8jNaoiLPZBSU1ElUF/EsPdYxgn9eAdWJZzPgWEZtEEhHaV
KHDRBbAJJLRqOgsSsOpVBR0y1T5bJ0XK4ZZaOsRenmsLvNWiZ5Y2LzdZFU4C7zoZ
TPysxnYgoqYDLTZuQu9M1TgCUb6kNU6Z+PpaS3H0K5D4rZRxwzW2I/guPJJOJcu4
zuAjESSaPYUoALxF8q8PYv61UOl/V1yW2uvC55vEDn/LwSIZQtD8rVZS6e00P6im
zE3q57D9y4+sIkevrKM7fOKOkAmFNA18etz9WmvXBQj+DCGw754G55SrpcUevzpq
Ks3vd0fb7E2HflC+NO9PJb3IWP/YOnoM2Srj3PUkNX5MiQtacVyHkjOdjZwNzOUx
xsYTbuOmut9quVFuwh55btiWK2g1J6pxg4UlnpAw4kfVcwsq18PSh8BD7IvGkMns
2X8ICcuH2rrJpzZXj9c7b8a3ryz8Bb0a1g8RlyuBCgkUljsSfQPupZ8Vauut/dbW
MpLuKzcYrcOXCx+70jCo1s3deDe+DL6LwwVGuaNiHir4sI0z67Pa2y7I1oiniWV3
YgE6FiAh7/MbdgVwrcn0iXcqoo3I6FQhDChjUnmKdq2WugTD+VHpdf57BxnLiq8R
7wrph7cKldkfY/bLZvmRSrXY7J+PNG7RsZV8ueUi5w7yQfbQ5epIJgX+vPRU2BRN
fgSAjXUCmGsTHY1+wRJhz7dUyR66F6Xywl+UxDf7IrTl9pLDrZPuoB0ebwsUrvV7
2Ft1Hmm2tlfRbXEqiuy0w9XanQ4O0tfi3+Z4ZxJZXz8zWwoSOaYhWRrVoN4v0Qz2
NCmeCw5mux8mXtPIED0Imq1udATbBVtI5yQaIdZYLCqjjbtDnwE0vxo8q048jA1o
9evL5mmdEavEYRbEsvq+K/1WkO0lmNMxtLaqL2UfxSN2qwgyCYHtgpb5rhLIRC9m
NuQIQiQaTo5ZQwRwU3th1E5pXvXk0THHfYhVXh6ey4hAWjhEio+xk1utDogSuKZp
O7YeXIly7tRreXQxI+nrnKmAl+69CMRWu3d33QA/xU9WinJDnpE1/mKUO6Aqg8fu
yTQyb5VQFkqkoTk/WshAavOwS2Te+QyBpfyUJrvZtMuxPTO0u+8rTmYVU8z7rZ0f
1CANbHVzFKqL70ECSiY3o6+CQM0+DZFg5bIr3W2Q/88st3nRc0DUUkqsWiY09bX8
wxT3D4/62LRTIQg4wPjxrNdLL9uV565fcJRu7O9BDkqwA5PRPti6Kde/fDdyBrcH
WGV7bmhCOV+n5NR9GcM4Z6Y8HNVorJfNKcmOoAwqrk9fb6heh8tZxarAEShUQMct
n9bUZpafx+6803TLEQXw/fPwWbCeYsPJku57mdAlAz2mwSlM4VTUjaK1cD8OCEPa
iZjs45P9fd57x+2ZeNSf5peHand7MTRyd0DkcevWE9jb4gMHXT7fahaCK8rU3+k2
i+nZ/RgonHhLxmuLpu41PIGyQWO+a6aNZTXjMCoGYfFGTug50nz9xj/oAwu//jrQ
dKRzs2wtTxFrHbxypfVo30d98upP19RGO8/13HYYwsnkjtGr7BQvqqO0PsFEEy7t
TBsI2zc/IeeWEDP6LQjLCG3V4L+a8mJb6KdFlAGNb0RH453lOZ+3VvUo0cI3tSWt
AUWNIpQqaO2p3JEAbMijpYs7Wx/k4vyQqC7J8kOcyNXMafSENRGLhVdOHkwwi+lp
pN16PKz55Eg1XBxGOWZYGHI2u8zDczVBGlEDUlkqRv/Tm6J5JQjoi8vfKq/IR7g/
l+0cY59363qGhnI9R8ohn5sVxpyjwJSJkOER1YKawJOxQV+5QR38Tm2EzB4TaZMq
YQNRojWkdOlpWjWpV+3SM42F6MhAavRBb5hISQjRtJCOf0YfGvXyQFfFkEGQFqOv
hnqmk83B6Ce2EZblQyHRILDByJnFNjU2TpKiLe2QhJm+GLohguoKmfpTlnBbjyTA
GsRUbzxTtzOvBoN1m98EhTZyHIW7pEcduobBzRTRE3mYx+Jw8Ny8e0/tMSwVl826
HDFEeHlTlACo1vMtQomR7iyXAeWKzpJ1vIVxnB9sdONURPzdoNq98d3aDmRAUU0U
Wuzk1rbuqyyQgovFpdvQWyLMPrNKwSXAWk+wuMUKlSStvgukFBgmiJVyYChpcypr
ukCR9zsTkuCYaWgOzsFYSYFoTM/OnNJsenkSlju5B341Gd3WWIO/6DymEtNF+81S
OnrSKj9conzgVCAdnGKkje9NpIGnlWaA3BgAP3DoCtKGzHeevxhh3fb/fPkldNV4
TWW/8PvQyNmURdT0mMoEQEFf8lFbfjSN1ijh34aGThsnuec4QJmQxJt/5tRNRscN
D0h5CJKDe9pb5VJgyRhyZYXTVE1fzK8CRPOUXT68D7CwdSGgKicjrj/9p4mPatZl
QuYD3eywu/ledv9bJ+OmuSZcYW2/ta/jwkcWaMQ0xoUX04xu7OV8ug10RBPKCM33
L3JlwNNSBFzkQweqjFF16f6kbuNs0OMHTx6Z5oNeel1lQuQM0Tb0B45tMLT1M7LP
HfGHyJwpS/NPwZ7dSyJybqiSoqsYOWrnDmIjarNS1U5+ouEHsE0+OJ+5xAMsIMN/
W7dCk/ODg6l6OCQc6QzDpArKeCcMoPWqDab/h9Z0SEQ+Ocxf9vs5E4hiYu4kdbzU
KD16/sJujFdnUgcohfgpt+adrw6qP1ujjHTGDIJ5v7q2c18U6AkrQe7vG4uSAd4T
ySotbBE53A/JbD90Gsph/+XBAOHcpYO2TnxCZamd7zpBxZP139D7Jd1k/Sy+hfcz
ajPIc8hNgLT+Z3rDS976DUGG9kxAaXQLQ+TudmrKVtIhZUl4uHfOEudvms3aaY7F
idka0D3mZ+dbuBmwlpaMDgw2WZW4a1tJxAo3JR1PhIKZi66ePQSJWmUmJNsRewO5
RR3Lv1EBXkt0YGyfUuigT1D2gidpmv+1VuxonR1f/PYd/tUhpiOR5qyzFJ3VQTG0
jGW3lbJrg4VYrD67WvMr/Lkl8uDZUEukurVTVZXPeX8GsRBki7HCgo4XVJn/ndX5
at/QVy64rPY+OiCCbV9Im/sK1v0ET9AOjRlqUIigzng2AGjY4m32t9hK49tU6IFb
3PoL8SjBhVF4/7aLEkcsgngVwqRvmz9E0Pn6GS/3Ezrxezr6L+8hho4kywydMUjv
u0Mi7mREaqpTAs3P3Dk3qrXC9fuNCq6vqB0FJ9WO5t7KwtcHjnMDx0B2OmFOIIUq
ovenBr4BPyGHcuVvYwZmpuEg43Xhbu1reeU93zJG+NqAuF8WTl1c/EvWXtyaKnTE
mmlQiF5KCn+qW4ff+kBkf7AOYAhNFMSXnZx2egTyAANvwO/WwwS7063FvMAIX3gp
j3N2hafGftg+jTvBEsl8mheN3Lb1g/OVMeu0fwWZFeI0SITuDUzFONiN0I3mfe3k
r9q2gheCXqtKX6MR1Y7rpC5hDoy+h93v4rf13mfCKYZras6DacZsOSgFfT7yFypr
g5NEn0c+U9BiSHr+27z/VP5LAptCXcYRhi9lCMGhuGDnnZdyxY4cmPvcbvnDoWil
YdS0k2MIwJ/Mup0MwT2OGL+XYCH6wQJinaxIwEnH5dCJ8TqLkxwgatpDkAGFFUtH
Hn6KNeRu+SVX+lCiPFm6d6+inDCF1Gpz6zZBAOU/bp6KR941VoOCm/FIT60vyueA
wuJUNjJzVsMjuvbbm/crpaAYkPAqDbRUCdF7CsOjz5gJMktcpXoSjI6C+Hw3HGjr
m7RSxLgmchXgS6MEhQhWqCG7QvmhTQ5wA6XvEFW4ibYIdCFT3Ersj0+U4WNqXFJd
2IyiemeBRTAnltrWgU89q1eaw2uRd7OUO5iWaY32v7GVM+i1d7u1GQjMdmVq26bw
ffj4MheBLfRi1mqac9nAMS+IEFo5tBzp6lLMeiBf748JAhDo1rYcEimcP97gClkk
gExeJvujb3VjJBEAhe1EMiF49ol3R1FnNZkfx9sMhdj/CCBGGkZwNVNDD+vznTvZ
pS7xZ5fX595Y9Ne//pHhW0g00I0FJIDsOMI/mJQGi31NdZXhrP5f5CIPzVWJZZsS
2JF6vK8SFkch9foUvyEZQ8MiVM4rVxAe4wFK1S+gFY4XoRm6IXaa+Z7sd5fc4mu1
uWMOu/JYfm1u1LrBOAR2GVCQZhesTuqT+GTpJoONDbWrNBtZfLFpfzmeYYIPbLKq
MoXmdflkkFPBJZlZ0MKb6WQU4NFgl3FJkfaWysc9ZDYk07U6UQtk/lnvj6QR6dtr
roPRmzzjXCN+tDpziJLRFrj9f0h9jHY58eB9FXjAjG9qAE+P0jKTfQvVkLgwPeed
pSF9Zyw6u9CeM255QtYUF/j/E72lXx7zTnmtA/oiOpqiPr8hW1MOn0DNx2qCNpP7
Eb8Lh1zMEvlZJ64q9k8a9J09Fm88ww7BCbiwTI/dzMnWxaTGdw/2CSv2fu1cuxQZ
NhTODz2ILQPu+3ypV+HHOCccS6adVIlcg4HbAXX0LWmqQYFtDXgFRe2CHjAGoKF5
zhBuufrg5mqtxqz1YcuLguLiTZY8b3UBInmEy+jfH/yKSpgsXdDXafWmmF4Z2p20
0hj1fhFmtB+6F6YK9U6mHhUu8yr4s13fRVWh4l9xjnaIYztF0QTLeEPuGzJmkFBw
SzS1KiEcyorQFl6ds6j1kTYFx70j6XcJctCvHOLID57bHASf7eFq8OkjJGd6X1dF
yyz19cLnEpd84YoVtPPZzLi7VNyRABo0tTjky3HYOtWJPyyjH6SO4opCz1dLBTCl
Htyg3uSJnfDl/pblq4Tt1DhNfueR11vxjcZ10xnGdHuqZG/MLzEoqmnQ0cuFDMFo
9uNiy/DOwZVw8HgfkbDUgvk4+hvrrf0u8VHY8V0AVE0gQGgoBlYG//X5RwtUcGfX
mMnQwB2uPZQSOBgVDwaMOsyMJG5aAyKLXsDwtCCugcFUqzwzuuMTlSeeTgERXtIZ
7h+bRKXMxIrpiMaC4G9dlntFHbrP59hvDDRHqbwAGG0I/SQhi68tBqtgkBzM7cpN
31fMsU5CVE9IADGhwgkmZbTFZXmCglj9H/BXKhdO2VwH1gOns3Wb13FTmroZcqVM
Un8DnQs0Qc9o3tRsrrbEzWQokzSygegVr8p7id+GktfVQjvamp0RTnn/2KfJ1kdR
UMYKypkJ/2cU3NpY+N/88tod7MXaNPUoY7lYivG0y0a3Ot09SH5zdPcKg/XLM08W
NpMod+gWTSIOsRbQioKEBhn5mCIhMuMETwDa/uHTkL3fxX/KxC1UIwdIl3VFU1Dx
5oD4YpC5nz8ytaYnLwIE043IhcpTjgTVa6jPezSVBK40R0bTgDIYDRWPsV3zTdBx
mxXoEKnrga3+3wLbixSiOSQ/rUesHwPj1mPk0U08uPZffpNJKCUxJmFm776MqlWG
1lTm4Vz1vFVFfflxcZuhDFrXlws5PuYixrjvsGvG2ZqrMBLHQOP5gxf07VP8hS/5
thZlsQSUjKlQtkqsX8VAqgG1om9uW/3HbCcPnI7U15naOiyqYg9cYodTVRplIxqG
MKEwEW7SpNg3x0kU3y4UrqkVxxEgewqGMekv4oABd2wucevmkuNqo34eMIbJ6uhs
n8yWtuXvYtwNRVG3FuDekRZwCLa/2GRLL0BdC3/9hTufwSWLTNJTnLzU5O89ZdUg
wj32AlgqEf27dWuxl8mAtdkmNla95iVVFGW/NKSq8Hde6u/KI4yDEqSKqAFm66l4
SP/nOC/TBPUISP7sckd4mPa6ozCCM+stR/13iSwFdD1iTLr582Z8+6yB1zi84aaq
8DXXSFJq3xUNbTchaaMSlLp4IsSmxs0ED2FnsOtxpfthEGEiw6sgSnNP7Q+YKqwC
8Iis9grmE4vFIAJzpBuSEQlTgm/bDWIxu0D6h/QNvukQE8oVIY54r6cdF56ykbHH
wwDbxnUkmeV9oaUHsmhg5qgECQ7flz9u8fO3prtR6kxBBM3L/N1coyZ7pbhrsJiJ
iR1V+xNcW/1SpqXhK2PQ/Vfm07Q6CQhT9w9J+VenFBL/bjzkdzs+kn/jgd9+fuY1
UKTn05Y1UYPwcqg0EWnUegyxGy1zRvgSN0kfyPSHuRFxdt2FtN/fLoYhX9Z+SJoh
QjGmlA1MjU+0qw+aU1OhIFkKNrAFWwoonFTPGRFN8kqq5sK7ls7NtDapyUWy/ChB
TbtIqksT/EI5gtVnqGuJ/GbG7FnxruOSTlX22jtlZ0wPUTFiPLy8TqJ4MTOyXbV7
RTSE89NldI/55qNCU6c7yhbO02tDLCb2yleoUXn/Wd0TNDCEkWtUFzC6Kdl5hs3J
cgMD15RXY224rixhFMShcuPp0Gj8CKkNEfO7u2ox5JCP/LPEbYsysCimqhWabxVB
imY6jXGuRdopKSeRyhnv3jJf5VDdUj3DEfr5xnIkz5Cif6pbrqmTV90isoGXIsxb
loqz6exjOZF7xxL6ZFC8xjS86Tko7SCyYhtBJV+UcarmiKknG+VWGd75TFHSbZai
UZNUj7KYqmespIO3SOKW9WiwqWBs1c5w7CXxvlviZGHeIDY3ZK5Rtm5GLfSpnVmG
+6PwK7U7yfJohvH3PlwwF4BI6EMBaDUyLbjoBq9REGIHwLxQV6a6HxlUS3TjcfEs
HGn1c+E9BYYexKfEI88f/2YqFa4LEBjsF0+2NxjqAqWxrBo0hIBLrPa6DNKEpesT
Ngsl80Cwh1cgN7Ib0EYMi6KHLarbFseeHm6VzXTO0Uk4gb2uVZrUfPbi44bHAbee
UUtXSTVgdnEE1PhADU0dSsw5NkgDntdN5y8RzDQ3bEzP1YOO+KVTfVBdyIRcSUcI
T5FniHu7fwhcu+zd+Ye2Ytyxe7SPjmditwX39gOz0SOsZhfLby8K3f7lA4Qtui2c
6WCnFzBZDszkgxqQDILPMre5fRwx/5xm20lm1Womt6HtGtJcgYDVEeB+eo1S2ytP
tJJrWdh37Jw+Rhy/J+apUCl6EQCv0HHEPnHASeCSqOhQQHA3Y7nF8rKkyjNOPkVZ
4UwaDxYlQIw0QT2HabgBComtquurEepUuc7B8b5NFMKzBrohZiG8WO7Y5xdtePlj
9YC9gBib8jkVnNKq/7MckEU4lasnaH/nBBrdBjurJfQ5kbNSnGzIhexNwLsIhRp7
vUE7bOj70Gf8W20wwJuiaNYf03noupjZanuzD6t3RRvuEbAPU30Z2LYea9NjwaH2
zADrdfl0UrXrwiIqWoHQMWf3PSTtWmqa1AgoPerYd3cY6GV6/5RqRNE/+W4U80aL
feH4KUuxyKrlrFMt5PQ1Fw+ebJY91tmav11Y1QHzDYWYw1cRuGghZb+TRd056JDE
hh+fpsekNGRI6ERePPBxHNDshzBIdNx81GPEQgP6NXv3AXFtabawU9WmABS2WSEj
qGIoQjcCWtI4P+U15CtXzM8mqqQK4oakV629MY6/bhnOtJXnBAgg/kqdyG+MxbUn
9uXW0MBN8T8Qerr7+zTTx9AffDmrIZtze3L3PvnmX64KaGi9DYfFCu9h1L/8BHTS
mBEpX+48jVZmVyMl3YUxlaT9Y1lSpKFzV/RrdjESQmH17uT4zl7Ohc6edTR7uBMP
ZPvbADmlV3JIR/hdesD0k1bHd2jsGgH3jTICNusg7PopnqzoCWw0tbWUyNTLAeGs
80PFvSeC39DwNLOgukHZa4PAnlRJFvuorYGNKYBl6ubRF8KdPbXCVxzyLrHEW+LW
kCdRtVobcvHyx+Ef4QQBGN5N5LDQUf5hUWx/31B3xY9bhwH7nEc9ihdStYDxMepg
9qODNukuydjINmJMD9VYCx756LOzZ1wX8RVnPngLO9sFAOrCAl4zixeDvci3gvuh
iyHbmYgqruzDEVwK7v4tWNbcCH37sbVyD2BIxfyhuYHSxJwgJ06r5RbLaRynCZ4G
3laDE7j5VmMOGMgCbdOjIVGqu4exMzkltOcEEZoJLDZwKEQqLn+RJ3oRo6fYoXot
O8frKx013l2HLYIfRtgNFPnPmTWCKykczCxobX6iLTyB8uTZQCu51MhkGkHin2GR
+VZPfTP/qAd/DU+NzcwjzmYm2iLseM1OvFBP44zlqxNCK2jkXD7disq8nYMzm7sf
tuByatBwmRQP5NjoHxHNRLE9bv5gN/1++Mz5CDQNJ8cZCjlt6IgjobhUhIg0DvL9
1psYILHFVMdxmegI2E3fXbxIbQsLyTd4FjQGxu2jKmp5DFiMremdYyNOJXs3PnMF
QAYc/AYMqEMTamUklqSThnJwMIrvJWRaNy/Io0fG9stHPHu6dI73+B1CY6rVYiTB
Fa0ZbboymR5HLPuCzIGXkgB3Sj5U2tw8SUkQ7fELSwqE2SvzRjEPZtSu3oX5tI8z
eO3wOAZdJySyqfKU/EOPU7kK+O15uX7QX4KxaNzHZLAcrZyo3XGd5zS4k0rgY9/4
Yq2q0DNh1PAO66+RHOCvNJHXtw1ToPH1G17s20C7z/NP0+T7nRRLIpTgOx9TVHTR
4sBV97khqiKZqg5qqKM7++4L775O5HXjHB/RioF5d3e8NliHCDeS9Vf5ITzjoywU
q3Pd7MfO5I1+38Mkn7HFWQLiRuLPRKuU7CKFu+CaK7D0lmnkXc7M5R72zlzzmFj/
7/1beu5HsFK4esh+8N5UWWLpUi0d0h+z3CMiCte0H5ffInzrDWA0tfJm8wfAJVI9
0ZnR2fUBYavBlcrF9nukTA0jrFaOg7wgaMkzeklDiVLcZfFqI3DVY3YFM7K8JVzb
5gDVvvj/teF4wbgcoVsHz8FEzmGos8d7wIkkxAZlTB57B5gbasyfoYLr3yDTkU/V
UHmNecm/0KdOVm1dbxubwmTGbh8DWprzjy9iY5yRmxalFpWxIQ0p6WodxrTZ90Ek
90MF4fG2Z+Id7J8V2DAZnAevS/fR/hWMsf+bQMq4EnuaanSwUN8c98adBlcapJF9
hOiEj6CRV+iqHu4Sb5o4XaMHa18h6aZ/6Ual1dQWM0E7UtXPjgfWgw+Pyp/6qF7y
A1+Lu9pVhu7o7xNW3JhsBfksJGrME33IusWIzH9Go8QqkPswkqmaC0Syg+Z9dAHV
R5DBogthELfx90Oyf8qTY5JhijySOznYWIwp8eg3FUHcKVvqhyW62GWE4N14M1hM
Se7ZjOfZeqIOirM/DTCuRGurPq6luOVfD+dEAhNx6Y9yDgmwbHXbw0aun8pSsZ58
dSrDC4gQFobCoSO7FREgiSwvO7r/YJgjYIWdaqNeXglWXIvH7RtIdl89Di/3d2cr
J6EJh1Rp/Aaarti8SwPKMQ8SBHB5hZoOkSnEPW7yZU53eV9tUw2DfWvnr1Nwbx5u
yvsLGr6LpovXs2FbP83hn5pb6XHBAD3Lmv3N7ioy/McjSmJ14b5lS9PNGu0Z/IV1
jqPS1EQu+nTH8qNwt+m+VttqIuKThOCAFkIlTAM6kZMEEPDn9O789MLPLfgJfAM5
OR3eOH1lvtUeYkpmhWL+D13vms+rurDydL0dbMgwAdTH8DgXt037BvOIpRvEM7Go
m6Yzxe+WFfuU05l07lYpus7yT9Zhv06RTnICvoTHwuliYZXoyi3weAxkSezUyYPe
FBEEekflZuuqPCE1nqjJ62XBdrgSLBH8j9eS6V4k+aSxlOKDdfMlzDLDPK2cvRVC
CkZl+9PoX95ERcXALdbfQneh9b0xk5XEp3BnxVL4fNFbbafvKRiCEf50EPJdreM4
/nkS2q5r4wNEq0E81jkpOlcivVjwbrTOSVux6Os/hUhYWFYOpNTYIJKBCvVzJKdC
Ep30AUWMJ6XhUURJkpXyGkqe98oilpsa1di/ZdS0YMPyAgDxL72KKW42BBYmsxty
C7OJlukusNLJs6FiPWSuWw5xOXBS1HTBr3Fvn93VMvsCRKSrDEwLCkrUIiezJ8U1
vjJP3+FbuZoEBtM9upuT+8b5m+jaHmZCwVHnEYiD+qhTpX0bACz6kxqYZu0IVp4h
6oeIFTiHlG4Ev3WBinhff4bKDbA5KbppwIJ2nodjdRVOMYlxj/VWmO4PnZTZGmGp
/DTJTMZd/vkgd6lbV3+7j1jh1oKDnsVCZ9ud1eKdjY9dD9fH5CVo9/+RAVXUTnov
iY0qrWbig2hxEgVAfeHoK8oUjqp8OXMUQJakazlIzydNr9J8QdFByGp7DxCiANtJ
udlpgnCjJqT5Jt/a0vaVu5OtHw9KbC0vl/W3CY3qwX3lQQJDyF7t2gj7aMTZfAfR
UnZZjzm9JekIpOlSzb7arfe642lP6InyTyRmNmbv2xxEG/uZ0Z8xBg8bXo5G4ghO
Iy6RUGuyP0wO1GnPtufb7lxhX81693qDRrjE67Rxtsbs2AP/Ucw+y9oTRidnuQSo
uyVQVUJtsPnl/xTG8FTGgP1Q3HUujjbDiEv1mhSLqecxZXkghQdnOMI5AQrPYrhE
7qM22ltWPm3DExez8F3ZTDO/MJbK1Q64EPHgoXVP/c+ihBwKtxaZvLiD03E34o5J
UvrCfPm8KTitA2XqWa1uDyplp86wgkGeClwUTBqJLdii+Mx3VVgayttPMkmSTiXP
j26QaBUcx5ZmC2X29ki3B9NUauuyQiJDO/O62EWfQZWK1AcGUpdU13riU7Hsswue
+TsbtkfngL/OplY4iANhqvZV830ry6evXRslutuO7VNoUbbDJw2bMOvt2XG2noxB
wd2Qo8z75xeKENfR0hrJodiGZwQ/TkSt6YR2TNIlpKot/dM0wNVPdrA7lTmxolu2
RmJ0Oneawf0Z7rH88uODbuPTZMF34zqGeDSv4OTuZFpd8Rel7tzttXEL8mROzATk
ML4QkyFRKOa2Ff9qr9XFoYM86c3h3EMAdQ1J+tp/8706j/QjlvvYPs5k3iLt1Cbb
gB/K2F6uvd6naZDTC0Daz5b+QEwMFn8tuoMgWnWfNR9QIJcjEhtRlfglYWhMnexy
huNBJdkQuHkherxu9cQWeqc6RiLoM85G83VeWPPjyAio7KSLOxPttYAKVS1x1TlY
0+VYv94QlqJnazMU803dcnukaHWpjL0K8ACdbi2CGTYM0SRNPGMD2lJl4iQ2iGTt
7jZXMRPzl5Y6CG613qyQ2BmV8CewbbjlVRVlsPq0Mo9XuRn49xOdLdUPdUpzhT/y
Vp/CJnyG2IRMwfu5xJiVKBZ7f7EPWXXmjyl2uMl8hITWXNh7PbeTUq/k3PFuv8cS
UUFajdvQXfwkwEgQwnymOypO6KxyUgKFedErJU4tEsosAwdV2c6ohVe04fm1oSnU
LIzcNgeeGtBQWJfqgnRGIA6m/ap3+0zZFi5rgYn2b5lDgz2C2Am0QlibsNk3+YUG
bl+CKYjotIt0rGumiUwCdCLVsi8ZAVDGJI94kiWhQc4FCQf+ltnLi9DnbClTd+Lk
PTiRS/7XZG9eGN5jwmzjabEuI864yxUGQUl/4G/BnbbArDV9dcbpLj3T0iHXjhD1
T/2m4LQY/wxcmkIdbbpQUDdcVAb+clSNifj/GknxLUir+S1bI2+EMYWXanW7C1YA
VSYoJIZKJuhubnMT9ipuvJ/SO3ElD5LghrGIYUi7kWIjivOLqxT+leobBH8+7X35
q8zTBzKYzI6CTccae0sUoPRI0I1xojFpvIBXxjF3O35H71P/wyOiuIpRip1ygbsX
IzLd1edVP7fU1bjx+7m0Tco2v8lc2D98E1U8vZ8Re3YiFuHb23IlF0pMtXSeB8ZB
Xv+V8nQU7TREm0vsijvH5eayXPIqdG4DOPKbvklT3ufSC+aQ79oIJL/6IegTDdyY
iBm/7JAl2vyrPjTbIUPEXksaos+iat/LUqo4V4sqO17XyEWaBNGCKj8LaAnCT3P0
UAVHtbA6G7w3RGvRZLTBFxSITd3VROWefcG1ZZ+w57kPXY5kZ7He3DVnXExZNQQz
iTfclDHfE5/u+qpAqzXwng4MfM9JPbjDl/7FHXeWEq8wR5RiCo4KaDnuzU7s9/MV
qL66kOwemkfitjFdOEq9PoJpApU36JLt4i9WglTQirQc7A1GHQZiwbcWEdK1H4FV
VX+mPgh46lchIuRpJH8SPa7TEYLMaDE/a4kPCJvqX/9vvPpQNkfc7qrZkRcs3YSF
WNjlGNTKzE/Wnh+OlRYVMJ4rEisbqZeYS3M2ktPD+mFmACq0rqCfZShuDYHrPVey
BAeWjAJPrU6jcCMu/ZlPL7dIh22a8JHNcozTs2qG1MEgO9hgZbkis65k4bAwZ0HH
yuJbPXdhJuxxiPP7lu5blVBhyOeNW/XknyLEC1o+jLZLoD1qW+lgdOceRTNJoSQx
Zy/2jFTXyuGWhLfaEj/acIud+yc0wrjOKI1Su40KoPal9s/2rufqLScQVHaHrSbw
U2tPsnqYgSKdfbIv065AiChSH6nGTUWS5qmAxpNbtvUC9LgmI7OJW5tn4eZbahdv
bPxP2ekC8WWn2NXmCCj5m4rtF8v3uoAiIFdIg8OnlI+qdiSGR5XuKafoW3ZAtCV3
RIJTPvBwZg5xXYu92pqfFBnSRLx7YjmTL/8stEef7sOqv4Wq5I1+KACnAIV6UFqS
FNnGrND3pXl/l8h9DMnZkPoAv55t7s5oubfQKZqrR2HJbpS4uNpzybGzrn0buvvR
jvRj3OPrkMcZDE8CM/k6ad4Evy+ER+YiJ8EToJbYAHGyWO78W5B8a30dyfZ2NGv2
ynH7ut829BlqiM7LPxnf1nRY59+ISVH/cpYYh0WBiFdqH+AAXAv0ksdM/rSaTIQM
DyhBETj//ZNiY054DQlZVdg+GJKAcCbiQZDxW7y/l4kZcrFgtWYkcWrLV9fVEtfN
MLGLa8EsMpE0ARGXnwraV89LEEaga/mXfrkh/WxR6o9jpMytk0lnPoFAXToh6c9i
LIK0kyBQL0/AYXbmGsUz+mDiDFP8PKJnKb+FE3jquLKEDdGUidfjGE22gDJJ+Cjp
N7SHuR+qiG+OMJnW5kZhxAXNPIcm7UYasTrQdO5UaTOFeAgStFyg9zi8epBUYgN1
697znTlnnmffx/y217k60pntFuNVY3I2S1NiOrY6z81jK2vwXJdPfqONxo+8XbC2
GjVAb4uD07e5ZGfsUIdRWdWPeqqheUcGG2rrN6DT6D6tsuOn0CM1EU2bdxf9LdC6
lY/it5JT6RSvdJCcnS/cZ1erRAJxKY6hN5hezyCvCaF5supf3sxaFpNuAYzOtRx3
ZLkvy4k5x82rsB/RclpUk+aUrtXppvnYeSiVOtRqKf1oDN3ki8BU09paSJG/Sthz
jzLgDBkMFXqZuUGqlU5bPBG+CGGfgXvuFbQkYU+0mqaPzMzK4O2pZX4WtW62Svzz
QeBog2XQnpnEOhNYjGRwCE+TIeQXQwx6JS5YLK0S1htGLJ3oVXpi9rI3T4Zveaoz
l9iRb1gZC4c5ogEhijdolLBwEW+jsqIx0Qrk+QY8LarRBP3jeh5QWyOpaErNtm6Q
sBe1QiNGNnQArTtUz2EsoWaG1xekOrAEmaJv1WvOCv4FAHxPgmyt2wclmwjYWALR
iJupHWJSMZEMI6Yps+unM1B4n8DoXjqIpjd1PX4rrEKMShVxTg8c1qNFumWYe0NX
p7zqpDvNF82jTs8vbmlpSgXidp1O1YIocf0RkhsdsDWaLaPfabc4Oq83rr+dpB3h
AkqcyhBe4yQr0t9hDE7GF6rFA0ExWwCV5PrVI3yWJuWBUOWnAk59K9p9aS2E063U
zXZoxSziHK3brGkJlesJV5ezJ1t6OJ2jBAzfOW29GnlKOOM7vIQVL1vlg0cEr6h8
rUCwuSna9Sq6MRSZGK8YOzabdpFKhSINsskuLWwJyyFzYbVy6c1xEY4ndlOaSZ4O
pSWCBInVAUorxmFw96ynI2xO4nAblcZlx4RKmH0glfrPDFfoMjn1DLaNH99x1BHw
FeLN9EmugPYTEdsxKSt3K82K52lkVKx+J1CWLjAFHyzgQFDI3NQHMYGVYtbD4gsp
GlDWRFN0ud3c8+ZSboweHo24mjGFTVv4T1lkddcohzH7e6I88VDdVdJ/4YRjAbGf
lGHKvuTSmLDsfJGqcmAUr6Nv4fMqkgiFmDixaHFxepcu26qdNSqUrPUp7iQ4bnKv
pohMcoWPHLG8qzm3SCTOKpPL5c5/Sjp6xYDxeKs6hfBRj02r8UDkB2WnGZLCB6Fp
hY4ONNL4CMcmDLTS14H3Ubr6PpmA2GtUeeh9l2LVLHfskF87Btg7QPFUPvGrdkUN
wjlaYgATOB9ZsBaNB9gkmZJWE6EeYnTW7xut6szIJEhbBWtUKpTES+EN9hHEZWYF
FFhzLbX7uVQ4/9INh18O32e6GiJywbxvg/ev8wecQVnhWEN5gHtfQ8SN1tLNBGtI
RId1b1ykDl9d3a/xSnJi/GcZ6VOZF2hoBzaPsfHIGw506I61BUuJ4MATg6ePw1se
YY1p17UNyXNeijxuCDIeXvcl+K0rMvY7VH2DaW8CVKGkaKZmqFurEzbg9AMIeK9Y
oTBcx2VVClbIbiMXW8BGG9RhjYpHGS8+gQj4dtUvQtCgnN+NcuUJeeX/PvLsd2YE
eieSc5eiDp67UJKfpprhexIRMF6+lmcJjg14p5yYcpEQhsXkO+SawQolVN/Gqat8
SVjbKMbOxG4Qrj8q9ycVrVe9RZLG+xqgYCMvLqbrqaG1T2wFDhsRpeYzfiIRKz3v
34eE8U2qfYbb07OTXjTVTov5aEHIr5A6mhp52Kh17BKhARBsByBn7CVmAnkmi7lo
Bdim78louVyAefLwEfE19ZXF5a7hDkvF4Kv6PlbKYJCwtrIxihi4xKTDB4Dk1Yp7
ZtEL0b5uCb8kDIYkIJhT2qfqEm90M1bgwedZ+uwCf+3AL5CTZX5m2hCsRoAypkRQ
EyHMrXA1qDfbsdbuMJmRznbTRX00JvrHTKftCwM154hpmlEc7whVob248GBCc+nu
6yEgqWllCc5qAHr2t4Go9QMge3i6xfhCeoxxugZBzNB7AeUVRYmPV7Fyaa6Y8Ujr
7DVApudmM38O9tU7zfzIUwAQXAALTXOEVDzWEJUZ1GQyS2XtUYvRJr3k3UG0L4R2
V9lZnjqB4n1TkW7nP3ePev943I4eYfTmZ+2sSsmRkvUriT41EfprrHz4i9KRBA30
6E2Dp814YK4j9UjJkP7ydoBDW/iUv/25WGf2zOtlCs16nbt6VtKKuWgJFN7Kk8jW
pum19vQLWOD17M4SzSzPzA9kraX0Uvgou2FFiqiZ1y955s1PrDV6m2E6eHKE/CDb
URM2N8dFE/KQdu9R4N4cWt89fGmEfG4BtxXZb0MS038CLgZ9yh7Kurcn/6tEVRsH
mex3GsJ/QfxWIz39ZHODGu5tJaWdHPBE20Ji/8hmYnRuPPEUh+i/hLtH9w2uu0bW
1LL37BY2S0KLUH4B9+G7J+M7TS0XJvNepAehDdQsEWqTAtuNUhgtO0WvvAQsdkyK
gsojDx34WcI/TBEf7sGUMPTFxBTwbM/LMrUF+OQ6KJdfaELEyXfEMMzF/Cr07Ggg
080ErhcW3+RpMEZePUdL637VKK60x/d/TPgo2A7tYmNyyib8ieZJxBYaO+ltvFOa
jbRl3DwM6KWpLJ4bP6dAdS7vC3QCmjAww1OfRDiUOQL+V1NO5bzig/KkO1yHpyio
Xnq+LaFwhkTeWeqUmVFIzO2uKrnsoEKGN9awr3WNYs4gbP6Sd5AO1yVsfVvEKNZK
+Btfu6s00JJNp44kZWJPC0lRSa31uLANUL06a2dzTHn4nqc5Vecca0fqdXTMTiUu
klbuhSmc5AzFBdj9M1l9AtZ+IH702k7MqTo1T68HbLVSbqVpCa8/aCSlkUl9F/U1
H3V9sEcDMIPePN6NwfbH4dwk0HNAjUKXsmq663rJyrrZ6JpUl0Sl4RWLhc9uDiSf
PqEZKJ9NC7cJbavk1I+OK3lWBCbph+KjpxaEepXioxnIaKL81sB7IIRBnWvM7tNC
Ao2I+JGuDISTgMVIuLFCZWH+JOcSaMlX/s2MjVh2CsUahqszhJasP6QXXNmg9LMp
BCHWhQzNignpA/ysa+Le+Bw7hZU02xr+5Pbck5RpnicZE0lhYNaIWTlka8nSmmaK
fgYM3tHGusw5hs9ORIMQc137IRzeejHbJOehq9b0JqhFme4C8yxb1+JMNXI/TM1p
GgJX8hY8iTwYyTeXkDWoWY5/ENbXWGd3767k24YskjxRxfBPEKtKiCyNg3E0Mc7d
kuW3wNfBBRX/ftu7ARsN26QY3MLD9KRZdcTzYp8BYm/kI2EmqHvIIs2dUrZuvyk0
YYzY30KWudHKHlcRrU2ZQhde0Y2hNI/VxDP20O5JHmD1WuSCht2PwG9C6IXneRok
NXcRCaf9DO8Zz/hTj+5jCWfvuP8+T9s5KFl1DXY0kNvROEdogIt1qk2awCY6/aZl
RVQqQUx5YKJU9Hx7dqespSTn5k71V9Re7KNoBNDVm6PgUhYjzMcOq5oaMW+6tX7M
opSm3JgVoVXb+dzArhxqwys91mxeYQcUhOksvKaxU7Ktj0dEX7NbNV068tnX7DFp
asGE4TpoYEPP9WZN2BRQKAem1S/bFZSnt0WmgweADeg0AOT5+a6ebsiCi7tPGyXz
vMrWoyQenOxjq2/vKoQMUPoTLNooxRchsUiI8iAHm7ZgjpWa6QReleQ82NyOBN6n
YETXKKmXV+85ulVDvkDF9oNE1sDroFwSQ/AdZeV9mnLuJ50Tj1pDO+Iu0GcC0iXO
/aiU3bBtwXJou0GV/Dm7UehwmKsIr7hJBCpk/9TI0k6pVKisDMDhbxiZDBiRLkUE
XOdexvgLlCieQEc/rpHww4XdfdMHV//Gw0ZoNR1Q7YfDvbgvdYWfbQCPKPiX1+SW
X4M8nZRCJ5s3WeNhFy2dGIBeGjZ5XRtQLBVM4oCxkr0rnmZ4cM0nSuZHDe2jgiPF
gXe/2zJtlEXYtoGuJ1fJsQFIWqY7p7P15mknua2H92C8Xsr7lFR66D6RP//QQibI
60t9094/JeOcI9QtuzYpVz3lz0SSvljKk+beYLPCY6AJo3BUyjaxMLCUvX2Yn1Aq
MjbtTUcCzxphatfZrBsgUG72gCeQkPEu3Gyp0HU84CYp0P2b1yG/NOoAm5IyWc4i
1KDBTaaIP9mpu4eAoJLnJC6i53Hu1bQNBWUtMxQ44/x4PBxqS4n3CcpAom1/HS0D
Z0m9/zjG4vuXZ3cgg0mbEPGsefCgYKf8Cm9E+QMlgzL5WYvt/dG3n0QVE78eWZPW
JLIoGZBpqxAW4X0flUyIUzS/wqM+aF0BklZJt9huMPPwmzXl3k/0Ne9k5ceAOeM1
Sb59O8ATLdSwbAkhlwe+lFXRSam9eZWODDB7NqF18HTdw+UIdYtbcQvTlpo24tI2
spXnGoc9hd6HHWL31MT8eDMRzUFNJl8yEgMoQx8GI47RgsXLBG5q16wJRE8KpCrM
Vsshd3hQFd/DMVWG59KRPhjBLqt8KnkEsoEnRUnlgccXnzebib42CE6gWAv5rNcc
XZ4slxDY6PIum+V2qQ4emuF1C6LNVB2baLYNK6twCyNwKC14NHqwTgrOX4IICY3/
eiRbtjzWo9chubEHAp92DHLWvF67dFmL6zsYB/WJjS4ldsQlPCZzAZ9EeOSPnL8E
9bUETrq69751VuNaMPM6LrHC2KTJOdB33gKUwRo/JvY8/XFLg1ecClzs/NwM8YIz
CcIJIr3UVvpzy/ZYilkV4j+JLJon6mD7wTRWb/9JRnGuwKZaxXk0WNzIXV232ZQh
h/5H79W8VlioDrOclGQA+pPBDyfjpLJPVWlSFtjtXXqVGwgyliy9zvmaQVOaUSC0
OizPd9AbPjTVaEbk73OJqA2AmgeDbpqt/NEv8y9vXauyAIQkGvZpC5OZmtd+gn0X
NM2k1/n9S01kRBzp1qgo7fCJ6iK3XfKBzWijEGchqq5FFlT4fBqv5IvuBEUhbGFb
uAg8Ir30DE4svfjw0AawOqGO5KqaK+35XrIM2H6UNp/wxinIug7Izd5t2GIGxnBP
3tf4bye7RYko6L65Eofh5mBm86WAeGTJB6/hgajQc5PxBi2hbhSDjWjvDi6/u/kJ
9hl0Xe+9shObqpaavj04+/bKY4CDEVHiTKu+7tTQpm8BvYZd2+ygsYsLm7sPuicK
AGN9piFMnbLD8gYSYwfvAa6oiM1NBMAk/k3U/BoL+Qy9dNoJEh+KtBpWGNgmw1DZ
Jx7EQo4vQ3dL9uX8R/+qfqB589Jeqy4UVI8ydkBelXW/RB9dZik6R+nT939aKYd+
hBEODdKTR5lduIp2ivDMQo9x/KGuG8XYJL5oZG4i+p2rJ3kHWeqD5IsrR/Aox5ja
kGCHn3jhO2jdelDnV+JR2lgW51vRnxUh24wZrb70BspqUrfE0OwgvlplVRfjihJf
/YUjGKESejrloah7BFqrpavozlyLeV+f6ZW2WmKf4/tL2q+GdlevMhlyfO7jBL/e
Jixapzg8OPN1puHZgI02e/zAFB+4LiYjUZSW6W/HaLs0pGOqIbFUoN/+nAYoMTHE
t6tlAIjOGsIVqfYOhJpxkDijyu+LAwju1hzNJt91oKAg32K9jScEE46bWG0XfRNR
lkJ12m7q9zRZW+twZW7SKGyuBXIMcfT1ONgueAd3GdjCaHfneIRmX0ntI5PdoO8f
V4lnvFrtB+gBdQIrs03f2M5vI0k82mu3nRqAOOJcnsBXzrnyRx6zJk2zoEbztApg
g1Ra1BFDA8Q/82U8MqQxmryNkGFCdpPaNzniNmHmUCQol1S5+n7pmb1vToxXj+Nx
hy9u5XgPCR0gK85X2pPwF31yJunoGCsC88TLMd/+O0pkl8Qzzb7AS41hL6AjM9g5
RQPsBm5O+dVVAnmV0yqLX2V2ZdUDYI38gjDv5CouD2+VSh5W3FBKLgQPQfRUP0Fe
B0BMK9ypYoPu2k9sxXV//P1OaUb/+JLI6ll5ojj9Elf27rhat8L2cT4FHedha6rQ
fsqxz/WI81fkrzK9Ax3CDInQ5MZoTHhOla95HnCONx1MWLJOTt6IEZTrkn5djdzd
l/F1CjV9HQ+7GxKPO38ivO2tAAowiZblf4ZsDVBPNLlMqBmrM5vwAiwBpKCfxoMr
7V94jzIugvL983QelciWcvc2X6bEVkHwkFVZEtOVYwRfsqPwwYMbAR/iGN0ya8Ux
UQjryx7ycFA6cudUg/E8xuEkdFqn8+77pvWvtYW0QCH5DF4eGhvfLSwN9D/pk8b1
OUpMRsehSuuFXBnESY4869I8urtP4igPfwKNwD92GPkOfLYXuC+HEAU4pgpR/Nut
nDUXAxdn8aoQcIROONI9/LE9ZQlhUZdwoQcKR0UpcoAgAxeUUZRnYHzttOaOFNlX
juZWHYQ/BXA6Ii8C6UmwWxvmLeq/DAkog+FsO9xJhgoi/ipI6CirB6ppMozBBNYb
+Ik9TZwNvTXa6TvxE6kVoOFGPPyqOZBbbRwaOLgLuIRGbDJNuhtg8TFbyUCSOXSd
1JVtIKz/+nzqziOE1sua0LbL00AUT9BB8W1aXEbZ9FwBkxmRz8ibDTk8nrpggWwk
3YEay7sdYN9s6l7cwpJEQ0Je7zNbcnrZy1tOLueQwijAty8sOFXlymG1RlMetZ0a
iSxxfyybuLQHgQyIBNpdjxF8k/YRsrg8Qrv/wnuQfvn81YlO6S2iOSZrqXvqE0c1
jVjtUntSlSIetYrkg9sPuaMHJ5Q3vh8ZyQwGQombofEivLz9lP2u4HOruxHLaH2R
lv5V1j4/+3jTGv7/kFMMPFJA3GR9/BInLROHBthZIjpkHOYIgmfl4w/GIjejS0X9
cwtHSUnUC3kNqVBPrDHAhmu4fYMVr6UIjBvG+edt46ag0X1xENF1ZkXOFxNoDF93
1EQtOchZ3vWC959Vs2sipruXpBS2iQ2v/RDxueAWJo/OjqUam7HElwFlqjzc7pTg
A1VuE/OYNe9KslgA7MweI/tXXsAUZRhl1Axk+g37PHwDH105s6YkIL6uHbm2ZlOg
BMLmda0izm2237rMZcP+duTElAwPC13PKgf98yb1rjLpvlZyRyef9JrXI77w8EBY
axGK7WEjX9CmMJIqJUZSXi32Qe5emTFf3ubEcm2omK6ueDfCGQyFNB3+YpIjpuaP
cKXWLRfSSk+U5s398X37jIt8zwYX2WfU1vDMlZyRlWnqlxEf22p3S0QR8D4H1gnt
uGBlV6uJos5EDny+3wO8oscisVaI6XkLSXbQNASMRt4+saNh4A2/tdX2i/n/Imli
Rho1s0pvoyqaBifcg1oyTG/4F/+uB988vKuON8JDU0bho7FjJLuzzVYbCPSWDusp
+giB4JSFBUcmxRDwGbY26s7AuWa+ECkKCF+V+3oZSpEPnr8OAunLkvjRkREUX/aQ
eN5t+14mZy2QDAK4HdFvnBfGe+V80JDS4GdJt+sbrKDYKNaqQzBeYre9n0+G8yQi
yX+E8Cr1xQ9nuPKzLkPTeG1K0uycp3LaoVAK6T9CyMFZcAFSeWYRBLgahQ33os63
mpAhUZtQ68eet+p7hbnI8XtLT3gTIlYVKAyplTk4GCVZwlq6fCFKR1YjL+2KIp43
z+y0SmgokKoHc1zqIG+Quciseseq6vJj9I7B01u4F2IAvh0/1FQqMrEqZA51iqlu
9LN4J3JZ2FfFTG8GHh4PvSjUGYZN+MPzXrvYqISv6ZjAeMb4DG5Llo+tQwPmESD2
iQJZefh9NIkfoJRgstt4GiL/tmo+zEtAJMWucOiegkDyVYZHZlvb/ebfSbeH94/r
Qjjwjzkx8qPCvWyP/2fISC+Fej9TrvCAZwbNN7Wb1TTZMfmANo6D2eHhFYxPmt+p
0sqHVlqdG5O+QttDn5CZ9ySwNH632E8+e2uYdHfJBYb0USH1XoV5MoC6h44B3A3h
kNIK5RNxmDt2p5F7pNG/p1/QC8QhuzcUGnPqbOoio2beLJc1uEffSwA1PszzSumv
nfx+jNL2CHwN5ghQ1t31ot+0BG48J1i7ny/WWW2/eIxMK6RDCCyI1VygPGFSzBmV
QPN+0Yt5XtwaG+pajgsGRIrnZMy18LYwFo1KWdmBMn/MERANg61RrPG94xXGaCe8
wqYpkkX2V4nydEtpkMRAAKo7rG9f4QT8b/ir64jFCF8Z7ZuLwQc0g9sFPpniF1wL
zy+SkJ1Km1+bQ0Mhok6GkFqvO/2kbEwKuASTjt3kbZGkXz711DMV25tgugXZcNs+
qwBF80doU/FoGO/+ABfEzftjR9wn8itNIg7oirnv85Qy8Ti7FHeFWNaY0ZC04/8b
UAWET2qrXi7F8bk59j+M/OkzuddeTZ3VRDvNv5kRScFdU5v1h7l5I2pMGPjG3CD0
GWruMXW1xHQcmiklPDKoGh74a+ddzZrDfe7obtN3aLsAHVqlP/O6m4mvCtzuJuSN
OLxHUnD1lGpcl7BWBM0HtecpiRy459ptShrlubACixLppmh2ZD+FgcoqzyQtSx4s
rHpo7LCsGQgU4yDa/c7kvAwg2jCg+ZtFTMXaIiEvhNy+xVHexB/yud8MUrFbc1y7
IXPknj3wmxXgVELhckfyx9Tc1xccVn/+XW0HcW//6tVuVS+psZA/HPVh+RutSjuK
bDAanXEwFpdqVAVvCzWjkiP96SoDeoPO6UOlt6cLXmowcX0a+wjraLngmUlDdpOF
+1AOaK3isBdZZp4/vSkE5rVN12qifJpfggJShT2yK5fxgl4sVhuG1GMiQhXyLFPY
Qz0wlhinHRpRVgPnrs2R3dDjV4Nrk4M1TcJOi3wxqyqETst+BEUn/jMxSAzfcKA1
ObjF3Gik4H5SLJHBZovVwqbshipYdzO4qu6eEChKieP13DZaK6il1R3C+o483qNy
5whZed9SJ6vA5ZiG7dbhKQAreBBgt3IYqg18N5GfTRpfZagaKNla5dMDFe7UTxQW
IiXM02NEEhwpwpCcnPVgINcRrJ4eh57RUuBtwyfTQGTU1b8RwIElHkehTgs2SajQ
+6tHW4515GhYFx5XLrzMsOs5XCs3csJNf0kiQeBnF9VeJT4BLVfDr63Z1oeCB1aF
0YWVQSfKXxKO56JWvZFgkUDhbnbBU7eUW4AFWoofa9IlYdFDIqUKkyKcpT1Z1BNk
zo/eiTy1MEPOIBHJfVxraiD/ypEUgAuKSiXdqSNIxvMNsZjRvTabpK2/AHERVS7o
dFcPhVtAPsMuS9ELPJwFhwq71UAPFh0hCU7/p1XoZJHR2twUIj70nDdG3TqaEWhv
NP5oeGMO1ixECzTWt6HSu2GZ+icPqTOCWyaXa6wU+b5r5Rn5muBGIAUW8xA3TE8t
Dzq737kT9DJZzvSyDj3I0/iyRPkWUjWXK1IT9mZ2libPITX08Hh3HGUgArSPKNqm
67zyklCRMNQlMZxnJCR0ta0xOSXST582g9F0EkJRolJ7E1ZFfscEvFrymJM/jJCW
pf8EwUqam5YtKJOefc4mcOSi487du/BJ+oMcFRGaxFeppTabhnG8sr16M61mrkX5
DXvilk72+9Xo2r1xaosvpp9W2ahEr+dwWrkyiU18IwwZh+QDDLLq+hxrlc/AIpMZ
9ZXrSbzC6MsEL6zfXP1fR84s0Q0BbBGXynnmTrpQkPdIawffaDuoneubC0ZfP9LZ
KQDHyCZJCWBoMOVvMQUjBESmqIN2Mc3BO8mjQWaKjMRgUQVKXWrOyOUrsf0OEaW2
H9bCbpgzM9xS1jDp1mqESbWLk0Yn70hsoTqa2gWM9vYoboB4Y+omGMU56sinokt+
P3mXWIRwPrqxUlnu4I1Ogpo1gQiY2Uq3d/T+Y9e7PnKkvP53sqUgbCbJo9oS463Q
UwvpbD+Fevq6Qqv8wXypsz4cnPLszq1WHoXvnfN11WU39Rnt64gAwYnm9um8V0+V
PlsJQrDkKh1dE731Vq2JrwNpKa2pLxFE8Z7ZZPuDbCVulCoWOYj6TD6/paTvuMZO
FGkYozEcthvwiO2qNHVyJ/lsF6pH6E7leYRCGCBC9huMOdBG/a8SKjvcBAERm47r
2zM6qTsagr61EWYZM2NmpkKoTKq4dFetYdKzYtszApXGDU2Zi4kEPiGNsU2nG+T/
gjE90hDGBiVq3w05ivKQk5Hgirez7WDRl5xSdUiVsbyfEHMdGpU2dddcf53zQlxF
IJmbYJCSO+BpGvdBou7fsETcU0SG825ZmJKxfhGI+ZyYgcorlIverovgWTCJkjrn
DYe2s5uF7+HMyVQKBFHublk8xMMHLyALNy027rH9tESqzEF9yWREd1o00eTFjqgW
4BGAxqvKGnc5FH/v+4k0WaAecuYlGxdXiZNjxTZmKPyeVX+d10k8UllBsdU/y17y
FIbipzuVU4QJOONcrBvHFdWhOQKvZ4XDR3/f07yvXpqCOnknYiy/+lJ0uwQdkAJ8
psJhEvEh/AiGZZZHJK7tsO71HH4ObSLGKAr+FMPavTyjqZ4EkcIagHL2fEo5ln9G
4sw/eqLrp3bg4renHoyvo1nJXq4qvdh+lWT0CW6X4QYI/+/0ZB9KKeyXGRkIWDyK
7OPf4XRw8/WoG0FkLxjJK/4JSFIVczQw77uoqjel+NNoqd9chxL1LeqJB2sazAWk
Ewm2IHZxa6gvfIMcDRw/bR/erKnW5LiDDxXRRRwKzuEZDwhcMmP2nuhQvuOyIieX
EiZxJGOQbSL5xd2wH2apBBq2poFHGaP+J8dPrsPhrppRCrNAdB76Rm5G4FbIodvo
BDwZLmvVc2guPI7PxIhgcE9xvlE+sU3v+JyXcLIUBkh2LvQ/XQPYUBxOz4aUYzHA
PF481stZISaovwlNcuOW5zf3Scv1cjGxiyIsGPdaR0jCtoxDri7yDxcSeFsI2hnt
uoMvqBUJFRAfboa/5HmNDjEpSRxdyPR0ohJ3/VRbcdWbVFSOEdlUZgxV60oFYgaN
TOwhpXIKTXYdteZczh+KWo21o3OGT896Z0EZe6tp3WpqEcM0uE0V9ut0jxQJeozb
IKu3hrTrNy31Ts65XQfiDZzNztHJU1ibSHl8jppCDcqyDCOasek3LgpRmXpxm5lF
rixVaLdApchBfEagfylLpr78UsT568jMrmd6Y9YGRe819IcgL8sXxDfG8gplWNnp
1Ft1ktOwCyW57ijez/UZmr7NeQHrWEyusp3mpzj3CKa2c38v4cyCm7cnc/Ph9aX6
0sumXCYD+W02VDpaPJ0W7ucCCczUgjvB4RMH2xKJ9/VTC2pk1d7xa9VYmyEpmm4j
WlKRoFiCuxHk1KhtKNGkf8yNNzysJXz6pyxp5+FKKPBa5ql2E0uSYmCwz7OV3Vie
emBzdUiRldnuNoR95boIVbDR22KSnurFBZ2JMQgjwwwgoYgAihsJAWmw6mQa3PPt
dT95lr4yfM/GXqUsQVucYPKZyvJZcv/RqVnfxKl/7mD6esr4BZHzuKgzoutO50rE
zlB5K71oIvokQtC7a1uxAUEVITwtUmPxOvvA7qf2+UKetCDrk2Vy2gd41dagte1W
v05vy3I8bthZJ/BV6Qi7myGD3MJoV6oeHT/2dT5CFTF1MClrU69Kp5O6Hi5oxuWG
dmzk7jcfHWkSW/ZMCUDj/URq08UhSGaLOIagfJq208sKZ7JW5s4ZUMMH+zYnn0YA
sg4wdR+vpwGtvARxqGeHWXhKzCrlCVE3uwvkEz508f2jid83MK1DabvBFapEnCrC
2v94Mv6TGQlw8MqblOOT0cz85i89FBs/LceQMVcz5IjUkjtORUjk3Ml2PeYNJnm5
FrS0O+vWSonvh6UFXFhvnschh2nIoiFxXGskRnhXVWLIwlXCyejTt43yTfkKhcHA
EFbG5Q0e1dQX+95BJMm2zLDheZANSE24srGGc/Id3hucbjNXj/IpwX/6Y9UeAJEV
xQ8pxsg2VzHbvdaBYHuW9Ot7sN6uVr4Xj3nNl+mTzdEaENvj4OMnjsa9Ql9EmQS5
yMPbR8ZX8kT237xWBKBO77Xin/UKrYCsE4yFkxK1+9+t95NDO7AhjtVTvUfxzKnr
PTkwTm486WE00z7DJHJ3+e6E8VMqjz7T6OfyG6gq3otbW0RTIhAOCfOhKFHd3Cjp
szwmh1DCHm4daDJnZyCRJsbYYkxjsVY6hqC9y4B4e3Tpy5pSfsig3p6lSW5YNgre
YxKKk0FL/EQ2/7OCS4LlCclPm1sLHG1RbbBpiTCUFIkz3WEWG9Jx/1bzU7zvF1ho
UcfpG8Paq7lkG5Bmq+ably9bu8tR1z4kA2RVuCtv9a2Ydl0RxSIKBxQIzDd+PGSL
UI6WfoCj2/ArE8g/W/93F8q0GID3VwEp0pXzGKamU4cLoSQa9k0Dns0TwCMto6bn
3uWJtgZuvc9G6Ae7b42LDW3lRD8ysC2J5gFh37GpwColhbi4o9AjJOw1KztY4aCR
YlRsjTnfM+LapT49IH0c72rGBHAEaQcgV4xjBmolr/+L3X2abSzeT5fugHw5IifX
HEcim6IsI/8K8sxYzBWtR11t93VQCMKalfN9H+ESCqRHKvO66P4ZSToqPMcmWOlz
pYYDrnlR6KpivucuEPPF+O7iIUaDWkWUvhocK0vRlwSGzJxqET8HRR+fAjr5H4Yi
XzOCxcs1aBgQar1tc9mWmyRNqtPSLQAGChuBRluD//EdCEuJoDmZRZCkS0M35fbP
8mx+HGsco2XyVgtz8YKnLDw8k7FWhFGPL0n2T2GKvbCsUcrXfhqUEWAC0YJP3Rqt
TeEUm7U4TWrQ+S5tnJfPwEFlkWl+KYtac2Qe4eYpacKNMNi3YGhq3j74J5eGebko
M28YRa3I6qWWj4qhUiL49ID2W1VHYNo3qVtDXh2E4pLzl4ip/3ILRWg3FIXGRsUb
6FYO7wAVtJJWWzA1aSas2fyDBWWO7MlVv495hyYG29Lu/Jvns908CwsyV13X3/XF
9U6g6lqiiSeNkSCk7lksEMLdxCHC8e7iNxY+mNDLQVLXPfxuEq43VTWqH1dCMVkr
5GYp1r+OQuFNueT1o6gMLjxNSkzXqHqjHy1etpR1x4sEjz1uH1HJrh20bxu5UpE7
nqqHe9DN/ojSe1SwJXc0xp+oBR97j0eSQDSQenm3kj3cbP252RCsvA6CI6kAVWwG
w4nydRUIjxozbkWuWfSSAHsIS6Zo0FfxJxwgEi5hFsQpNdwH53wXKdzzQXN7HUBo
KqSQXDG32nAzd7hjWTZ8Pgrlt7xEPmN9Xjl47+i5oOWAiM9hrfT1gZ9YCx2Sr+83
BK22QW4qVPOu44ORaFXjvM6T9AR6WvGpkrfR2ZQ7Lfy5exPIRUup0sNw7CgrHUac
i546GH49yx9pnX66NV0XOjH7MRBqa8EiKxB6n76UXCHhE+5uj5/iAcw38HwrwO2Z
/xQKYPUyH4+e1Y1P0MnEK0GUih8PxzAje/jwAE1aEOYFBzhRRANjauItCq/HUlXM
gIqjtwiFj/bqYSFm3oAdvgt8Hf5dveuINOCBv57eu1ON7ssFbkI69l/OaQ3x9po/
QTDxdRqNRoRH6tkwDkLGJdvFRAxmskJ//fANRYORXTTRUSTLLdYHH37Cu8BHRjOL
yzKXouHacPaERhOXCoFO/cNISfIR/rugtVwpPmBHPjbynqWCv3CBQgTsvQ8DpVK4
nFddwZXv3NrudliwjzzyuHiFs7ZgBcMC7R75RHncqxPEmsnKNJjS6hePo6Qs77QI
lvg0VNP6EdhhSGkBAjC6aCQsOizMtITD+VT7S5OqJSOTSeLwU53PoY+m4Q+ZeEPa
0k79YglUCNscoSGS0hSBr3PGp9GSu9J3hKRu3Uq/eH/7Kdro8m00ZZ4Srrqh4QSR
POvQgQNLhFf5p8uXSuPReVN5ykN39o7M77yitt9hZo4em2JZTe/HS0hXp9zNsl30
NXsrCwnVAecCM60MtnzupgBG3+7/DV8vQTG9xyoQfIrKjQHOqbz7Z/y78F2INRqo
gNYoJpkmHYvDo+Tr/rEcBAYEXe9jt+EkuvHRUVV7JV6Qo9pUJd+5XCnvwMmzH8NJ
Q18i0nvdH0H7rVsADSPqYyoozpttgXi/aIL0TPZLmlUPFupkgMWYVPIsoxkYcLrC
HIduKP/MFnGMq5ckiI9DSqXUuJ1Vt7mIuZfIu3GwrwwUDSiUNdmtltNBTtG0tl7U
b9XaoswWMo2dsoPvzg9UNJExEy0AJMv92ZP0gdS0nbMwl0lUm0FHHIe64thdcRKR
8RkjRgpZFY/j1YDwJd6/h2BJtgQVAL0XBn45dg+gMSYAcnlErP2oetY9Ry+xItcd
PRNS/CJP9qKAhi/qf8IAEgJhU13FifDxfmJ1lMOruogarwqyoxXNvzshyr3XowvD
49ZnTD3mXs1aSQPoeNb6wCEqhy5xBemGvV2CJOKiEodxf/pvZBBKoGIeCOzyNSr7
a2xQSdTOGi8P6j1r30Ia5fO0JloMk8Deztiq/GEJ7j+wHl5cuk02LPazWzPoA7zf
C9GWQtZxwq6NbRd1tHMpRkel6JljTp+HcEq1NY7iiVjB+iEywxvFCpRv+n4H7Yed
uEfoU20KMZ7m4hdgxhvtXe3MTGJFbOLzQMR8LbpnmxgY5Y1x/ssZ9ymcihy+vPJI
PBHdXIgnSwXtVXZDaK7joTdduwX4CJ8i3chx75jIARhnGI/pI9KywYoJsc3GWgLG
0O3WmhDp4t1gbnE6D2zg+H7WSVDhIEQM85qqnU2mKLixERVVzvbLHBaII0pHJzRU
leNP33XAu96W3JyCsMo2AFVMSTSO/I3+gd8pT2InCmsSGJmL5VhV0eO2A1G/ahRn
Ep5ab7MiwHu+ZeJV7a2ScpFM+2qfeCCGvre58vKuUfEI9Eb7wtAJMlWqfs14VZc+
FJkOx7qnvs8VgAIgv4V/kBpkH21xmpE8SvfhUaildajQR0x+KoOFbHRIoSXaxMDH
ZLnRLVs5enEe7SQpvwyC1JhNsNDSpCIZGbcvdYup7CJ/m6U5ik3Sfylhn+Adg9NF
tTbtAY1iiQ90HJQ5eVWpsq0Or21hEGijHrkyrzFRS8cZUxq1jlRkJoW/yJahAqyb
aIkFjWYSVlDONjTmKEw1Vc9+1duqJtZe8dEhXz9/lNhZyUqhuGuEOg1+RmRpbC8b
wMmnZTOVDiYdmAfgakqfiEGpl1smbQWmSPDrDQ0tX/lb4VzJD83NsRY9xe6Bx5oK
17xsYGBMRTbSUv6mXkdmxgAEMaOSmKymejRiOzodY0dkbbh6SGush3XwTcboR4Qh
6q4y+CsgsViT0wkDe9p9slxIcSi5v0CgZaJVSdmFp6Xvxbv3XvW6pTgaoEopDna3
LZny4RENphp/LUB01fxxY+gyVVCWr9LsQ2IZDZbcLqngGaUMfno4ORo1vqYo7Brq
EMBRNX2AUSB+FaieVC+BiINbU/8HuTRso1Yt+K14lx8rfYBMdziwmI0gAq8PvRBN
sfSDycReQJworIdsmC/mQUze/qeAb/OszHjacCHXxWIWuKpJdYlsedV/6W3B3o/3
RHQSP1x4xGCkXZgSv+ou75sxr1/12g7fuWqiyjPFBhFSxy6cHm+7SAyDzYBhGgGm
zzf/U8+mHqyj8tasnZUQqjyBKH3F+Mw+HOnumA1x+h2BVb2Ub0sMq5FtXjCUI4l+
TZjZSGnjtF06tHYjO8f1KWMss40j4f4eM+PH9MP6X8iG25eOdD28Sc47ZXW0kO4d
7OfrZURmdS2D2i0VGrjTN9Up+0zPWWFxZUK4fpIVw8B0ansACjsHU8S1EtPC6osE
63PcEnhDIQ12D96Tve6thLL4t+JKGTbwBCcDr/P7zjUddMzLPiCeFwf+jsknNaNz
IARKJbAjmG8zyd8RoGp9ZQFlrkqT63FFXWNsARhpQ/cnM9Q5NBDqGOturvjz3n0J
yYV94LApB7fI7ssjwhwYt9vmoilwHBif5HIXs9TXr6GrvTdQPAJXOL5fwynzKKjB
ntRHxIre1xmpA71VegBRPQjxPNiXkJWA0T2l0hzPIjdKx2olsvX938kzZz0W23+a
fLKttPWR59QZm4zzNvIOrvjd6MK5ijZHkPC25jgMxTiMuS6OqVjrdvie+B6FuN4P
MAGLU0uQ5mOrlCwMIB83ARAPdC/sK30dUv4X4ZN0hDXR1e2EoEfl6tD6Df0OUI7z
IOcbPQFkDmEzNAR9iqFZlZcE+vkbS6Df/sd8PdsXPjAfBzN+bhvK7AhgA8kzHK3f
ag/D796uVtQNUK2NCn1M3gaKXNedPH2OfRScpFnvAqW27JwN0DNenI0JfXoJbeRl
C6k56UjjwFngl1E07jTIdRPPMyJsvoMwZjjXaMQrjPP8GSDjslnwMWCA9IGQJg2q
Jp7DihBLuQ0hMMgoS7G+drCuwlrUOM2YljojtVkP2M49HZ8dZ1NDCauZOOIR7i3a
Ztg6B2DtPGH8t7cOa207nRF9pLk3cV8sF5gA6D4O1dr98ctEIGNz6GV0ljASiCKZ
FWIT4MoO4HL8QhheA+OfvcY7xx8Ys4sjaTykdNIXIiQ7SDstymSdMIHnpn3Dtjau
k2FH5BJbQCV+UxE6aRY7pbtdNF/1tUCsDI40SMNu6vFR9hEMJ40QViFTYDxNLaXe
+QyfMRvg419M/FDO9P2eJE2wEoHUXXKcxvgdD+JYv4iY0mPaI2wH0jNDqgqzx++A
qn5sLuK3PI+FegnXr8Ef9EGEnAnebYjLoyLxL95AnfZIWnWQlKXjwzRHhp7MRiLc
DsU/frNXQQInlKBujn8TpJO2o+VFlqNJEkxJiwij4Etd+Vzxdi9mAHd9TSmZtSw2
3wV42TAiVHiCBpPUFp56iDGZo01chhCxBt9WcXzuQT+D++40SxbIrMB+FKGr3GJf
gFFZuXQaGU9bAXnWFSgpE+9qFuC9JQsmBm0zublYcFm7Hc3Zu/vwvoAiToLiogIT
XpcFovHLRGqtN5/pTAInKD0HqGPPmNoybYlewnnqdqdNPONkChYdvczSuaFYz0X5
YhV5MrlCXwoC+i/h8ktv0SE3p1cIR9PejaT84d6cEDzvR+8dFnU2kiAajqlUIfJR
/bEtYCcfHMraEhQM35JBS/EiW0QL5c9G8opVYx5Fu4hS5EtpNrmmhwZL/P1JTylm
ACUWbgauIB3cw7frqh3yaeOq5dPFV5y6HFYhbQSo3K0AkKfspjugAMdmwfNSoT+k
PxoPYlxTEIvw3fx3/liTq7jQmvJs+O795aptnlv9deU7GL5o3C/ZYtRIrWMrenl0
T0qQ99Mo9X5UqUMwBAnfalgZ77TN5nZMS1AcMmvLDAhmX8eZlYHSi45rWZzqfqFa
5faCWmTKInHJlZ6hmQ5rPapmrjaSXh8j/UG4T0sR2FUV0jIa8pCZegvvyqRvCy88
9pgYeylsNS1imbFPnkciIKjifeU08w0LA8hKtsyLovkOulmIejhV21jp10lQRqGx
93NGSoqGiii1r9GvJGtNkfHOf0h0Wbt3k0LZfrSastIWzXWiGKvw4+yMTfvcJxs8
Ezx/q7RZIEc/t8fqMu/AMh3E+ARLCY/Zt8LMC4EPll1JfQTlwkEBMwu+QsP+eJfA
YBzevJYL6QHJ/1UJP2nMJUgG+sahWpErZZq2LPOwagoqylqv5c3RQWhiK7YwDX3v
1P78zvtEQEvsm+BHVweUJeloH4P+B50IwNmxC1Tg/keJ3z3pGfto7tahXbFRETS6
om1CwKpmLMkz0g32BoWAywNZj0J3NVuBvp98yepoXUDkpo5QSF3SsLlQ5bRIdOB9
YG3bvP1meou34zJpHVraAUzHjA7+w+KO8szOdaW5V/OT9RY+xZnNdKNX0VR0j2jj
wG3UsIYXydgmHAbOLPY3jwKMwy002GlHb+PQe/3QjpklNBw6opReIIyC2ylIHTno
O+WaTK7mNPTGN6tclcrZmyMEvrjbERB6rVOh1+1VqPMwb70nitbF27XRFVkhuVxI
AXbT/d/qANfcIBbc+IV2YZa+IwxuAti6mxn7SSTRxt2FyMi8t7Krf6LWe/f7k9/L
nxX7CbhE7enxx7ak524/IxfyeVfYzKMQv4cpCnKesAaTwFuIS0TQHyPdQZjcckRz
u6rYVlYREBwVxN5jkdqEK3CChHY2o2AnToKF8IH1I+XucrjIqQQjEBvZk4bFNXPM
l8tHjk9jynMugRFPrVNibw2OGwq0qQvcGDPRJGgWUmNB2TfK5WYAbgdnhwySIo3G
icVWBl6x+5H/rck/8xV+HeEn3Z9BcLTswFPdI28EOK97v9einlV8dFcT1hC3wKHN
nDMfIZytyunEVlqTB5FUAZ0JIrju9jpleK+i2/sjz3WgWzNQAGxGEABmR8v9QH+A
Jej6BbjAQAJfCEW13ChK8NmYv7OUAb3JjUNvMiDchEiJA8NE4d14kbjRQKVco1uB
FBoNA/3YfceYFm4YGvHJywTpQQdEre5nC2H3frpmJfHHpp99Dlnd3ENOGtO8DjjO
st1utcfy48612qF5fJjIYLUmgJ5enR5f5Bd8Bx3GKSvC8q54REXiSVxe+BkPcDim
JTi/6iQpEWj6NoN9T52zSrIW0m84CsxIbnaGdek7zmPXZkBAnJL8B5zwHA8aS/nl
mTdQsMfPsd4dt6wiXyGfHpyIwXT2eYWfh3P4yOIFtMVCE91RLoMd5MvYDHsmAr+y
X7Ry1SEFnbJuf0KRp4JTz3KMleTtJoBfg3ZynX4PSzQcBr/6//idaQiLtsTgPqYJ
dbSs5HWkdNg970EJ7z01xkfJYC7fncBkZiilxM3gPd3yGiBn08DHbeZyQZgXwyz8
GZXlHFqrNpu6nzbwWZH+7S+R8sYDr3S6hkpQtV2LqFVpN9IWrGP1wQqP5NR7FLs5
HrDg9lvdSJfEQgqsmxccodCyqTvVn6PQk9uCIjQTWwh5BDkKmbCLsrEFClHJiOD9
Ax7p7HFVKzBWnAOIMEKTZjRcN7aGVsSEDAJvQeWfSC0uchYkqx/etBZDJ4tDvYTY
toLO3FnMGG4/VNR7yxbGJMWoaksh4mlyMzxH3JDpglm5xzCqmhPlUxrdyyQW/20h
eAdj+3Q5VAdnDFZBJCNA5flExARa1zQr3uqdC2HuRihCsXzEk82KvwSI3V5UQlEQ
+bAHiwKt33FPjfU+00x3OuorAPoF2kjVxCy3V1piSZMY3UCTDOxIEM7xnCqAWmJO
g0CZ7KJWZH/8W7G2MeYKXqduK786Ashbh7E3gng0LeC6gTgJVKIfmFp+IAg8KXlP
J3tU3xFnQE5BzKVB1asfXvS5lkTkeL07SkPsRU2iq7PaBK1agETM/hSHtvArVWCC
fH52x6oy3mkdPeNj6V//0mLuYhMpGUr5M0/yZZ3G+lHnIiK9uTC5aC+Ca8Td815T
CQPPWVklBw55PMyOpE6V2zGQHuEuSw3aRtEuhwiD0NJtxbpk9PdEO4kQ5aloxf/X
E5rvDZHNm3jwnqLr7T8vYJ2eqOEzbHfg9ZejfwifJkXYupA8EaS5tgkAFewurUTY
ZOHUiGuPpu0GOWfXB3J8Aa6mNNziRqvg0w6LWDs5jX/4T1BGpcNzgBm7KhWRtzpO
bdmJ4mL9RgzCiCClA51AHlYUQUsS3+PbsBioiiFtHA0Pw69hE1Z9+6hsREyYF0j1
9asViSqtOaYBRNKmIZtU7ccuI/CEC1wdGKK2XN+Tcony6fRwS/jc5x0hv61rDV6s
1C7z20F1bDOtirsvDYLB70NPbeg3Ac+8W5l4FH3WZCVNI7rzy7XTTb3z200aZiNT
XUtreZbv1Hs5PglO/HEKvDXoHnSjF4du+pOXKxdzRELqILTqBPTgPCIYfNuM16cP
R3L87KFMP0GBC8SE3OXz/+s1BECOVT5sOOb3D3h1WB4tgGiur/uS/SUYH8xMT5ls
BK09yecypLm7DGosiiqKdjus40P2jfazEi/abdalg259R9KpXXmSGj6XlaqMRgqh
wNAPFmqOQalcDS9rXrkJZJI+mJ+EJk2rt9ptVtBU0s8Q+b1eH8aoDSuXTQtuiZhL
lc87NJYQCbzaYzih/3zJ2iGB+WfMFcSWiXRPpJn7eBplCI8CzcgmjfbWzTdFiFuQ
xmij7knNGsSjWumF2Uei0pBUp9ww2EHEjARLy7AgXDxKcbI0gNlTr+HQI0BjbQ5u
DyMaWzL4cyDwWuhVgcL/Rxzmmpc4ReGb7KPNIdWvzhlKgNzuBBSa6P8bSRHO7uqg
JZegG9fzwAPtyIjiTZcYc3wuIZo+bQizqW7RSPW3RBt3TNxWOJKOdux+pZiD13fV
RKyOpd+cB+1itC5FbAQCtIIHZqSr+aiNfov26vEoj+ZJXVeHm5kmFNTp7Mi/A6IB
yy06it9L1dYc1ICeWl//ju45OM5na8zIVPWJZqjFpGHdSgG/ttMHaFNwJpCzSXW6
AmQhI7Gp7CEmSPT21aOtUSSZD9u0dWO5NVhkxwEOGP/FSuXcyGOtbRXYdiiAPRxf
bLSXx6AqYMYhV/VBBHDdB3AcmCu0wPy2uCHAzJ3v6xE0d0cxNcxlZG+TkmDaHnE1
klolR8d+tHRlDHMoXJjgM9aOzDYKzNmdTC0jViTEB5ipCdS80oMvp5MdQCx3vKGu
djDJWdx2Aj/hDdK81FaFAYagoUWH7sU3ZupHTnzacYh25A2lnrPqs8MKQAZ1ATbV
tsC6AtCZLLX6Bv8811lavB38qsPkNQrk4vO+qPrk+PRjvYxUT6WgJGXQBF0q9vJf
EUCqPXRa/rGsts5KwHTKQm3u19IDOGqkOSVsjmKuJ+dUf2Q2DOqpbXX4yZhNgZ4N
TVXEx6QDhdoW41Dq1rl7eCnGvPKoRmZfGG8Bzg87XeVO4ZLgZ5p6xxf89IrKVvi8
DCaMGNLVrTTYIKubqQRtBpgW+EvVngr7QDANofD6CwOZqqdoPr6k6w+iExDnA8CV
SxlqL+IWlErLrxoi/hqZ27QjOU+iDFBoJz48mJlZyJOCxaImRlyNnSzVuUJ3O9c2
zLAki2mM7lrHBc+6CTV0YKjkOhFyVwy4Pq8MiK6oGlmzWblHBV6m/GLqQlI+BX6l
3oEE3ipmRq2UT9M29/jYlSxc62aDl02PQNMlJ32dF6DJMje1Ito1LAyTStGGV03C
GsiaEfuay2wgaNzmj/0MivgbxUe+MgLph3yVorUDo71BhGxqQVq42AJDfHLh1i0p
KIEv7hVrHj7LzJNLCMOS3z7MFhxMI8beyszSPikd4mWfIyOIjM0MUN+pITLVyRs1
z0s0Sm8jNENZpiW8QHy1bsEy7MWE9/K4hYqvXugPJNX1BozPJJ5LnWSfFfkNWmxK
t3i5u8b1eSHKdfmlOsJIjvHCiBARpaRo0hni1tJpzuukaUnzrbfMKTJum1bzQ8SK
FDuXZzGaeRJ+JWkfiS5qzjnKOERi+l3qF5zKcUc9FckU3Dgk9cDDVA4ZsuFWobaw
UTbUVcRWKlVjLGBUS7v1E3QqiInN4nU14tkb1m95e7aRQOahhwDfnJUMZfj9ql49
hE+DkIFejhygu7HvldyMaaZeeGzI5s7dkdSAhsSz9s5xwO3hqDtbF2qmfsicgjGE
iuiPCj52jahkJbHVofZpnbqw7XGeeseJseOcBhScey+mAY+s4PMlbXAUBM5D8osj
+9tEhUB1bYF5k0/aymEQsXHB9NGyl7pHwSbxNcKuU2K9rwqQF3lfrkmT7tFryeDq
4vsciNUSWOhzXdZspGZVOLHwQCJKcZpiphGWmX+r41gDBjzBRG6CtJIdfTGhn5I/
XagRBLVXVDd9DDd6C+efZoTjQmbbBppN6aG/yIj1X8FjdT/ocvw65Kyb+Mj8uQWJ
GqyxJlKx1HOl342hV0Sgf0KlyR0VfFld8mAljiDk05He+hKa41O7ZmNmECwO2fAX
bjShmCZkJ15LDOM1lhLvXvOk8xhUy3VOG8zRMZECcg3KFvOVWFx4/GutAL/LyO2a
Sivrk8z/VedRPbb4m1pJL379aFoMm0IoR0M9kgqyWO1Q3hPFHQk9NdsOPp+ZyZR/
Lf9SQVVkifNIpYBWkoCiKuMBagsOPXXhm0GpNrkBxsnAQoGFdBvMaDa8Gxx2UmtF
3e54SJb9X7wkAjFUJ/0uM8mffGbJ+ufG0D7hOpK3zfw9h33Tha7Hq4LaKQq1CHqz
nBl6xwJMr7DXMF9WWDHqhJ4oQob663vAVmXg4ivGHz6ms4TxZ8o6vX3D/DAtFXP1
Af//NWoKJeQFiThuWKjDbErT7WsGURBCTpKn7ovwwivLvbGD9wwAg2NZ5cJM6PjA
Ivw0AvcwrfdfkZo6MGtt9jZXG9vZbPo9kqXiOeFjheSsXsFog6oIL4VBGx8X5NpH
enu4jjTo7+/BRd9aANCg/OLqPktFYFDG5cONlPHT1PBpjGysWKq1slICsg21QYh2
SSo/n2rCT99iG42ALWJGcCDKenNmj1R32uLmtbOUfrGZzbiQUlzuk/56hUgJnuIZ
4VbrfMyXIH6DsyFEHHIDBZuwYkQMuPtdziZRrHbYmIZD8RX8aLSmAeSXkkh8MEA6
gvw6zSCCKQJ5JkVj9nwzb+eil6iLkaGYOBbj+8OmTH1XfynPy5Ls8Tqoclh6jyZQ
mhCQMzs/E2VlVdWlKajMhKl+N6RgTvDZxo4d+RO59GRcLdPpX1Fa1P+jPgiv9uXa
s4zk8tGhKIDn7jneCvM7BPTdlL8x9HMMfOjyskb6SBA+Afl/9j+t+tHaWWb+WEif
ns08NSRclZuupOmP5ZBhSiiXSgBujG1UHHALSGu+h5m0lIWVkrRWNS+Hv3e3XnIx
s2N4lFavft+avsQ3Zu/DLr0H0OCdHcg/EfPB5dRGEeQRG4gNUbOCvulIMdwbz714
+wKfhY2v8cUgeQub6RxADw/Twuiw7WL+6Cz6j+R5qIP3BG0bjo/NqE7vRlpneO4r
dzuynvDkViyfzDR6nHUHSUkapamczpkgKvl0mYw0rjY45xuXLbaSw+cV7WFaxE1b
tvXYeEIiwq/OGXU95IMfQLczbnWl0Nuw+9cdYaSZkaT6BVBPPOo3qZ+5lz8ewPw1
GNMaX8BzzuQas4dlnI7NEn3i8Xw0EVeWPLcNP2WJjiO3YvaGCoFrLRZ3CY7bsjF+
WNaQ7NjfZ1McomVvpL0e/cRdwv1z53Vnlg/Gq7/3O9ysOzpTqrhhUoPnBkMEHSkz
oTBclS+9izvng8gCT0QN8DyYhhrEHdSaRDvyYeACC3x4971Ud/hhkZP6Txy4uJIH
hFXWAcVtJsjp1OssHIlv/CDMaOqa/t6eXKfSUTItQKmIewKuORRkrEhEO+wK7RdN
QOKA7exT9dGaCMNG34GtmTTN4z0AVzh0jbmHPAFodMjSKpxbTaXkR3iSAx2mTTZo
IPaPkxwmHtcs1mz3RyxSIKCaxL5y2bLmqfYGwgcezGlOcp7GIyWmdtl1N4pE0ovl
+6cm8lsEjk0MUA8Rnb30rWxTpGqjuvGyiZ9+jnBriCpA3Uu7HP81YQrbrl4puQ39
tZjFfGa9is8ukjjUVGthAHQb5n//HIxwIme7EAzPO7tRisVGPn9JatOfbU/vV88J
WU7W9kqRqOG7qC1O4gZgPZ8YtE+FDoclI/375jRPedWzMvzUHdvH7EWkjyw28ux3
2tGtAn2d3XwTVZ4AiRwseMsBNwNcxrJQ3rwviVuWtZPSa7qHpX3ipw7czdS66Dd7
Zb88ZFktvzTePx6I8m8ZOXNR3KtLSLDp1z65Yr/I98iCr6SkUsYWy1mhJ9D9Jyya
ZaN6Tr1sqHxq6k3ii6NXy93jH5mtIB1fUAePqj/gTRQZhZSN6xyYgcP+gwa5TDQD
AAgX8emsVA780YUu7f4pIyjvSQEYMh0SaSYUoVcAuBKpfXGEcsPoyiIAqZTf9dgC
9kD1uFGP3BBlLgmsU0Z2n+rv+TPfiPC0k13+PVQvlCZx5TZALnu0DTEERpzP/2fk
Q20wk6cQQFyd0X3Lw0zCSBe4kkPog9yPenZe3+OCSY8fKBvy9inO90lSmOJYZXbR
+noV1BMwG1uFTQfyu/v3DSr1WqH+CiCma1I76W/vW4qiLiQkM02pnvCJcFefXIPM
qcYWMHQ8QMiXGZp9sjaZs98WxUywzkKZP5RrvjnmGtHCrPMur/iL6Smr5PWppbDM
nOw6CKV1knONF3uUjek8LXMb6FFMEYIGljrWL0NqxE/wK+Lvfq4muTihdJ7U8Qqu
TwRMOatfuHW8zQIyNSJdYqALcyr6zIdghW8eyVQCq7EZF345Ipb3G07edIT254iU
AZjqWsdFfhIf5dqYlpioJvi2y43ZeNvDXqjZR4ReEH0N7l3YfmJR1QOVGT4H0bJO
Bd2EjseqD3jiYMeb2hp+sH1LicagCMvU4kfWrDHRfqfXHI1t+GJdvAzsOHKcipx2
sCzNrQy/bZt9Np/eZh28R/MvPdpsOY5+R4bxv63/Ll+atNUnCka1GW1A5XHivhaj
OsXB0K1g/RpYzNRb75Ahj95HtFZtBEtq76OagJKPkLC3TJg86oWk7QmRIl2O/OZT
cLk9Coh4MJS00UEsis3Jw9jQXLiL7dUyzFqN+jgW9wy30F4TYvfczx2wXBbA9RPc
ywPjj/p0kSsBj3DJ2i5PQETf8fG4BSQxWKgan2wLvpTrR4+SnVhnD4gdKgHn9BXu
Nh9W/oNUYjOa5qtXquKU98KJCu6VEVYX5U4YdctSMH1bG8p8PJ8pFuEWtf3hxvsn
+CkQMMnfVQhfxviUKMPP5VREzcYpg3rRTZPGAgYr368qcvv0d1DTUOtGd2SFtEHd
J+zMRajYr8kYHdH8CCSYvABu2r9z0enYQL++jNRNtV0m4BjK6AKNXv+BL8q3+snl
0cveQ+1Z008G11GJniQttAF3ZdiJPi80L0/80e2JN3C+loCK35vxhNXguYor5vK/
Oq2Mi7LwaSuzMFlaXBtWTNdXHNcKqNWz52ILRKjrwILRgz0sxWEFtytDwabR8aFf
82PPwXMFjM9Rv3Q2d/fexu2GtZ3u0Rn6HDx4m3Q0A+kCiqnmoLkWo6aniGahQmMg
AK/rr4SFuq0lYq5PxUt1ELtTo5BNmCJhc7OaOVQMBkOrnLvMgDfqADbtiY0Ust2U
85PmQEZFLEqbcuzOAWscPITlJG/bJupbMZm5sI20ctVoeNFTos+RI4Lk6folWmRe
PdkL+7cFql1nT+YTqx1edN7BiBCbyOpDcqhFA1fKpRyczNk1CLF6rUM5oOdBd9Ch
UIHww7pqXNb+YIzhBuvKje9XKmhwnhzPnIIQnxcRm+vcWr+XJWljUaPoxAxsGy4a
4QgMqsDD0VJFt9oTTgFSTeY5a29diOXpSWBufyV2wnmPAWwVPPta+cuu4hTF9Qfk
7yjRox2cgufqALs6MdQle6J8EDgQ6ZG4tqKFwc5yyjEOvEqesD/ElVP3H4xoF8Dv
NNUk2P1NYtU8zh9ICpvYZJqiRe85w2mPtKx/Tg8E5w/r1lAMME/MWH+0sqw83hPW
qvHruLp6tP0NUyEOKbb+ukc9Cf3+zajl9Ehzzq5L7m2DzsejipjwCFG3wJ1UtDoE
RVvU/o1TbGYRShmH6UbK3vsPRqXRJzLzPrDFaAU7k/WzGjPoyTkrkJJwEMffD7/D
eP5Qv3QVh/567oHYDDPzkZbre6Zoc/vHuY7xebXqqcoOxuBzmf7d0rjRVbRx1X9S
09kbYyFHTuzWMZwCwggCFnTHxfR3bIRqzv11W2tHE3RVaP3WQ6h3CIeLYL8nnEsl
aJc3B6GUK23hDsvqX/2VdOfis/OAMMUNYy3QlDSUJmXjphJ4SIjqp5sebVRp3lFW
TjxxbOkA2Zm9sX0Vjc2sYrQaHr6BIjNWWPcxHTOBWj6Kv8Iez8QfcibHkoFpMt8a
Z9N68Auqe5Q/M1r5/cmBoRpHukQyfdgKm0aLCnzvh1KSzZbevO5YaBNxo630cWTR
nqH1FKCq+gUpy05NK9TNlUCRssH2LpgfS6k/2O8kVvvl1Nt4tcA/eq1yHbzLA1qU
YOKnOJf6gyp6WbHjYQz3yaTka5wU5Jk9fyPbHtChH7b5UqmbdKoBXEw1dDjLbZoC
sxmwUsTGZ3fKnyX+8Fv4MHYHniksPzyCrZxdG4218T/WG45H5wgy7z7SuVkTcYD2
fv2dLUbfOgC35lcFAe4/G1eYg80zhqJegFnNgd4QvCxufpVk1m3GfznPJ+NxYagu
Psy686yZNmjz1JMP6HyzxL8UFI2TMdXi3eSc9BsL8v9vLArZglXHh6Ep5H5YVslK
Nxlnt3Wj3gGZ6YZN4/jUFWMDsZcCpMng/G33bf0THUMf7g5f/nz/ucB8UH6Ha41n
BlSBxfDCoIf8LEQ2hhNlb/KmFS8koHC8Yz9owKyg4vRxCVBOUSxjTwjNxHbyB9ou
exEwm7xbgYKOhVEQGLH5KObWOOWV1YiW+JrXo4aUwVWo5m/vfMNpNW3CCpdWgYBD
zCI0itc93WtWgvzDHoDJgs58GHTkYIGE6DMzd+bLTJs88fJvcsHnUnKlkeojPXMk
4lq/mZASBj749Aijcye/67/KYhRHlV7rL/CaeE3zAm7tu5q5FjzbEcqC0siHm4I5
FaYohAy4SjAIGXj1Dh/YP7jfGH5V4zZqtvkYLLQTn+IzJ4B3pvmNpfa10IAstPtE
YOZoqU0WXHlm0BTKfJ/9lKcMjHntYToqgUzwHRmQuWx5P/rnHY6r51iHM1+oiiIi
+XmuWT2fQ5U5YjXLNxHf6tL3M7DvD3ci1sXspwN5aDGFPVrxtmAG2a4XZN03aLT9
eCJeybxxM82kXZuNkmvN8nRZtFVeVKOryx+muIk1AZg3HT6rNZ1oIj6wv5I74G5D
2jIK7F2Kbw1wiXSvV8rcb5L4yHNFnGBmyItz9CImQcszZ8jsMVMkERqPcjlloFrd
dLvzk8yIve4S6Rxpcw8GsrbMncQuu5HRTW6vESQz0okZjyuxUnGG6Rn5Y+Yoqcco
1fa5GdF4DNgeThc/nfJEGP0QAC5MGz0Xvitg9yifbwfpjErAkUapUm/sx4oPhF66
+TBRQ/5LlyPzljB/IxTZXXj99vMNWrIDg1LN843DJ/v4rl3dJTJpPabtnKn47cR3
To/m0xWi/n0gyaBZAdo71Q4Acoqc58rMmjwpD0zFEVzqCoJeUXVjzvISdQy+8jJM
CqM71BL9BHWKL+3bvOeRtD15BGVK3J/NEFFnWDMkajgMY7PHhkPQlCmVRDJssDBQ
6VTDu1bCEWEzoDS+BXWpdXrX5X2g7dNvfvyBjDiVQrDSHSNUOo09LkI7v6PMclLp
R6ULRAezkyNNKd2UNM0S9s3zexqbjCDNjrsEGJwaswd0TEnHv1Byr9OOBV4tQlHj
AkBGM4v8ISMwMrv1qUjoH6TRu2BiWB/Duy6M6vmemvQLRIOMylo/KUKmbYQdFez9
tYcXHoyeqXi3p182zKy3lslfR7MfAB7HBdFDeJ5Fp/vhdXbWcTiqPo9V28/QSbPW
tL3654DjSNO5VUpJHjUAfQrTryLWZTNIq40COvPtjsnwzKQArGI1EtT0bUbahijk
sWtUEm2Ap0Aa6sYCs4mht0BBy806CM9WmYTQJkfarPT9lqStYO319AlwUWqJkJWN
X9cOUdHp/T8x1jHy4sGGx/90RGeFn6v6hkXkp72KBvICfgwqlbSVxSpeGi5Lj3BJ
M0zViu32VFAQYsLpqhtprEwdcirSC3yr7lxbKZ0hNSb8nkSemhS7vkHJPiYc1LOG
oqdn24AiPuZrXwo3Q4FT64L6R7GpSVhSXyzMvk7MnhKADyVsoDPqQLl+iEITOorD
p5hBjpe9UrqjOf04iI/Z8++eSDeRK/syvpHlevz81qeu0jaT+P96/0srT7Mh7poX
+9OXGN9z260VZjlVgLSvYxoy4jkWQ3Qir8sYzLatoJ8jcBuD46U/TOMwsuhWEYmu
/ezibKztfgQbAe+HWhuWOJREfRKMQoAFk1Megw33EbRqDLU63JCM/hmkO8tNoXzM
FylwRJwls3/gKNbU0Lhw3KzdBHP5E17UD9P3EDXf5MWD817jKJh+S4eL//RQ2YQQ
zI5zfOUIj/aOd6FDvQ/E9UHWkbcs4R2j45MztQ75csaTKGZ7j56dKujx17HSNOAh
YqPyS2ytRzvMauqhH/biM0oRmsYty/DHWQMxRc/CeGq2fBWLGS0hZ+aevtElObOg
wToTNxXgVnP+XQOjZehzpywY/tZ5fqIHGEezip0gv3m93IouclXn1d1d1D6N0sBM
93roEjO1Kwl3/xvlkoiYQ+ssepvz6GmJrmjka1i9OFKPID2MNNzUqgkPjgqne/Wr
4pG3ceJs8AgHgTQqTQbmoxe+5+wATYrlutGPpedRLey/BIl2cUQZLfnjPUCuij/N
iZ5Y8m9J2xlT0STWa8hIaWDysrH7XqNEb8HEAdbfJK/Tn5B6NLvNOtFLKeNI9avC
mCBSwGbLfmkldWVDSYuD6AdwAOC6+IXM4CGViCK7O6kbqn7vyp0pgEl1/eAnvcFi
tEYa+8zx08TNbrX3GFjbSPEi3s9S4YllvX+PuL8khQhF31e3EFIClC1TdkLix3r2
nqMVlG42ee8KRgigd9HvRIYQqPuTra1/IgveqT7qiAoFOwrJQQwusAXKOzQ5pML+
Cz/yoTtMQGtQcZMQwgfK0LMZ35+NUFkuYIhamQ7l7kgHyHYFcuIiOnYmtm/OSHsi
HYiRmiDFoGUouPR2Tzc9h3PqV6q6TbPS6vtuOPiHge+kz++avbdBKB6QsEHDe1dZ
p5869Yc907cNx5SATj2sNDsMgDK1xJEXJYF5EsES9HnXAQi062vQ1Phe24eJhWEG
SeWxO8X9kqqGf4tP0PT8RJCjQm4/Lo+4xRtDAub+CqXmLXHqD+nTxTYhXZkHaYvw
+3xyh0ujO9tXjK3G6DBibFcfnKbGSQvutntgcTz6lJ4yKxO3AnRkrbdNdpJ0MnAw
KHTD51M6Cv0jqjwBmsC+THAMk2RERHRG2VPLRub7cZ9VbIkdqkxgeZFW8gHolqPN
h0qicaPJRk8goAOuQwxVyWtQvhi1EQwuDRE26DaIL2GYAvHxof9Uja+daGRifh/W
61TXtBIFqcZaM0rUGhQZgnZ4gBKoIxWMccEwh5u97GuNxNi/Pl8AvVZ3kGvgSy+r
WrZHprN96lQyTTq+4iQMl1TF5ROxkWgwdSS3K7s4UQXdclubLY6dP9Gn7V9+isgg
Us8J8PWx77X2qrokzc/6JSELZ1tEm2Nwtt8RGKxj0sUepfGjzNZtHyTIZa+2yHc0
v5q0Lrvn6l855b6lr1PRX7NvNMdUjjq03avxLMcNhKh7pDuUKJ9dVtpBZGT/lg9u
6TbVwaEznyG2Myga5Wf6Js0ZnPUOPb5PDq4RiK+PTrab4H+h7I3fDDwhdbGWo/gR
66JblLZnftnLlexWsbM14CNE/Q9YuqKztB35DQDh/y6+bCstm9p6KdSK2GsQm8/o
YgwWmGpatt0Xopb3sas0CBSvK8rIZOuOmpHrpmAmf6EtaJfvfeFHUjYb18IFtbOd
b8o16gPkX01tRjTCq86Wz+I6I2nlbgQ0e18VB/vHAVZL8WTooatRKHzM1oxAk4hv
vQ+uSAEa44bunOZO0dcCQVnZQ5tKqeASTMULSCkFBJpPy4Hf7U40nP+baE1WWAin
rD3+Cz0mCkKWR/KjzUIe6KDeKSRpiJX9alaulHvRI+zq00ZbaA6atQn69UVtvvdX
ejuxdJlL0K9Ys4EVt/8Wjay8PVmecNI9pJTzJRAIuBd+ELTyk4qvVo+zUZpXHW2f
zslWSeAQ9kRKuy8psCjq7JFG1DtC4AU5lv4vqkRMIy2gXPMvdzoNuzORPNdLiYvl
eDJMgPkEU/sA9dMdgo0qP0yKqaNmVA5qDCN+Ol2tiyQ+HSDo4EeDSjMk4AFYtMTP
uo+yumSuS04orQSLauaMwohLsbJZCcDXkNw8XnShsnEjNILCbyPIPHPzOIDOI8t0
xEPU6SSWbtGo6ATVa3Wo5V8BkwiDcBBwB85sZy+gn8aw0iJuCgkjYcIJtota+fOB
J2NUuG9r9VoHuNgKcSzb7j9YbiDxSP7Dyh7x8HXHr3+/HNU0Svm/wzB38rnO+Hns
AVC4bUxg9WNOwMrveJhSleUHM2hA/iVqxGweg6fI32g6nn3Z31+8mbs92b7/HqRo
w1GbH6TqgfpH0qDMonx55t7CZh8sBP2TcKjSY1hZQfn+kKPQGLMtvOhC4w/L65Fn
MyLFHHeCrCNaPGjnm55rdczTiVtisoVqBYMahoYpxyERTE+7UOjHabSwsiB71VEx
uv5Hu5uobDFRDpwNHDXM2vENxJohrbbLoTZ0I47/rHEmMmhIJl9XMaMSiJTjoEqi
Bncmv2ZtUqddglpqIhj/hwGEaHhYcvMFx2i1pputYsDkVYotEYzQWc6Nh0zzNLi+
r8SSm+w5yhcqYd425FyjtWi0wCVx6XC/OnQ5njQGiRdM41KkEoRmiRL+P4K5if3a
EYBqxcoigZ6wyKLwY/tC0a7Kr/o8cQP81YuPBLTF5wdpxVYqOicTxJ5aVeksKa42
LKrIKtn6tdjQmLFAOOzNMcWIjvF/QIs3nwlf/56VRkGLqePgP6xUt4osTkuyGoAx
S857m0zpxfL670ubyjoIHnhSzcEnOMJwHW7nCsSi/kqaKWLGSJvxxiPy4AugYQ2L
Y2tf42kWbzbMwYBXcJ8dwGlWmOesMLd0hIe9h/fr+lJrn+elo0RalIaM3Ezieacg
Xq4fph1RbcQsHP94J2mqgozaB8HN8JkixeKUCJSAM5gSeSQR7mwi17Nfj3qJLrUp
MoUFBwzYfKNQCsEjY5CWnTnRGAMsIdH8cccuiNlQTgGmUuTzaNPMAN92gSIJwM6e
jAkgIU+ssFqXHs9WDRJVQdgRWD5L0NHr8B0PSn74GEOS8GRnpPsLmdLrnZoB7ohk
qbIS9SR6oPajypFSDSHCM/BFVwkdFcPNw9N+dnaeX8XFCQOO/JRXcVpcxd5n+XRc
nWuMqOvfJIOd8t0Y99qS+nqyrDkrBgHzA8cdvbOjqNfOpcesOxOlOUmFrA753xFl
LU53NjLmI4P8bne0ICPUl8JlKUaY7TxdTWBtUSdb7vAfYeB4seTLpJc0nnCy/yVe
5dJraAyybAFQLRdD3jvdApDbNqczeg7DdHP/vKEufqw5JXBBxGxojtVm9tNjZpw7
I7X22ad7hJcOr3uBplDmlcRcP7OFdACzSacZtVuC1mJShnbNwTt1ZPF60fLYm/Kb
yyudCy1k01u0RpsciWQZqNsB26wH4gj9A5BOFvPLFHzV51+bTaSEBcXvmXO/BTA+
WXArdu8LkBa/0f3dq3LyozcPqy8FFeoyXrioSmOvl58bsczeB4/LMWuYFFEEfM+3
MZ6tSmlQ2tQF/XqiHpc8KvdgnDGmt/zy2qaLx77P1OMK9yJ0Rhk1KrF9LkhjCoqR
SmgulnxoTKGyNk3TIeHMf4NmmX9DF6yjERjnAW66UIrxwzSLYwgf0i8hvP2Z1MKv
1jmb9aix+eOL8uOFomqS4T00tvui6h4T9FSFSzNNYJNLYf/z7nEeogwOkc9sbOr1
re0FFcfb7WVQfMku7M/mzi+bo7WAkMLw7xCUSXBXizD/ce7EofpqK6DbtcC+tWyp
mKW4ISmUHikDJhc++56+jYUgKFh2VsYPrk3TeOiJYpnJg1qYDvTp8aY0WtKAUDEj
x+qyikGE3q6mZZU4FsjyH1Ex3A9mT2E5sUzyJspEW+NcHLPQ284d3uZZwqP/Q21U
6BIOKTPVIjWr2WuOfgaj926rEGpbrW5k/jfFQNoV5GEtxVNcfrv0AjVLscHYDhn+
AvMa/fuC+tNpcn8SuYIn5dLbIzTY59X2qrXHHOnm8EBbImiYc+T1BBEhKfiYyrhv
J5hkuFyo6Qv8QCEc2q12qyQeN2asL0o/89o3EI2dfKteRHZmCbeYmp+7od9451qC
NFTBC79KwbE8oWXrq9TlUKMtwgomBxen+8MnUOWWpS7hPlpgvKGp5Vfv18+D2vja
nZSNf2ERkYEx1/a4dLFBrdFMlg3quKpdnumEebrhKq1MdGIvOjbyEoVFaT49lWFL
EhBJUAfTeiil/KaHia0STjiWG4EGA3/MRj/neIyo115oyZHcQCDtlPEjnSDlsAnZ
ZG5hEzVx1O0YzYEET5/qTBkcvdEeZa3zCxOVkcwaEWwPeKGAo506P62CQWGyWLqS
SpqGBLfT562D5969fysU8gFBoaYjyJdGL0tAqmf1BZs9IfE4NZeXdlIGC3ncpM28
W2wCYLq+ggDIkFa8K6C4xMevxUtg4/mwXL7CdMFjAVbxQqCBZtWx0fYnTBbN5cnV
t9YxGz2pgcGua1hUzanLDdzqa6IFsnGoQOfd9+4LnDFvXU5lZ1KuDhnBWTQllX9i
sdvIU3TBxrD1aTomIBrIBYp4nE9mybw8OX6nqx2jJCQ+duZDdmL8ZW1mL1kvEX1a
0aHP3ElGwajIhnnk6P2O/eg8xZvQVJ5GPI1Nxc5ew3ICM5G24Y2yDq1k0US3zCaQ
aXZf9FMaCaCMbmfrszhRM0QjPfV6wV9fA4I7ZfyyJn9ve0wk58bXqSUMaotgkQo/
LwbUsKpMnHVc9qwBUsTa7Y3dGbj3c1I/5s0gCnGZu9kXDRfrrPpPoTRlnl0TAL0u
glntu/FYstJDuZmjL/jN9O9dLj3qqPPA1JYLbp63EVybqCKpppE6OOYUrlhd/op2
2K+/ka80QhulRD93iG3lKCBBA5Zci107PsIX3P5f6dI8GUt28mvv8cfzjzQjm61g
jYMzJRRZGgArMzn7KDkT+uBjXc8UHn5aHMx2j5Of3XnaxaL60cTQ+3Fr8KKfHAcW
iGfc/nvCiOPXxKkw3Y46LBZsATYFCiuR2WzcKpVRnRCBSC7jXr/+HAImliBcPxcc
HkFIyTQaODZP/jP7pQm5W+Cf3aCLRx86ZO60iiiojAKiSE4JA9x2CB+2iaxKLbd1
0vzwcXGcxiuWegIJJgu7DR5O3QkTYs8eRWtDqYXNojojSzg9vlCLzIY4d6BDm0fN
iNKQhbLm1rU1suJhBDNbIJUogPQlckYL5FjTAwmMVHAdFfkKSQAtYgpILXz4px48
L7e8sp3IVLShPBEGcS6S8kjIpK05fXknLWL7LUEYG/jbJfUeoNIkqEr5f7J6S8ra
SDyh2YJFUmiq9kogg9gd08KP1k97z151ZUYv2+DGD+tYv03c8iS9EYsrPpBs8vdk
F6MPKYi8ndUHwjUZ7kSBb0zgVmt6ZCTK9xiYT66QXcqj2njpQUqfb+GwG5CIbquc
HKvlQdp1oy7+EKAS+IeAdBrUoYLEWyYMdXX4pj5K9gcJj/PeFYOYAC4DriwIW/XL
hseSvdxSxH0PVymLH095QxMy1ba8uUFHqfsyoTpMdULlSmFXoXkjsRHwT9Pj28qU
pfYlIeWhZrZGS198uYQIMX80R2MCB5rIOUfyXTOhsvZsWJMkVdv4Negy0dSA2brj
iPmciA9KiYHWL45yeZlkK1ESh8o3F/nVNF4zvSD3trjinhEnBULc0EaljxOgZuCW
vXGUsmfEu7R2qANsSSN8TT1yjLa4mSCPijM/zOK+0CbAnJqoG45kRbsKxUgMlCTl
ikWs8IqdAOToEOoCGPmOAqZIq4q8B5mIVJRZZnbDTOusNWFDOAYVmTCaL+QR2kbx
c6AzL6SEh4jJ5eOyhfyQ8aKRmg9Wgzw9Bw4LtbDN2EDQQ+1pUy+SZ13HMOmtDrTU
RHFklQ6ym35Y9LcjOoyPIU6l7QyvUz12DXMndF/qGeXO0k/h6b+3g0UEL/6Y34eA
UBoqYehf5otIvjEo8linf7eQ0aG48FhLwoNk3oMazQCet4hH9AjUykv94sgBwjUu
LZjvKmt4uMCXBQ397jrI3+DMiBEAZuf5jFWqhdjwNW/lTBoVoIqFobPbTs4szYYL
KnXbiogo6u3q0l8leR0/T3s5McbeetluS5S1UKDPuhPAMYu7f8MR50tK1Wvwk7G9
xCK0Kkr9IqlnIf4pcg+E8k6x3OQtgPaLkIQw302WKClFaRFM3PIw3EjPTqNlO4kN
Hcrb4GiVKrIzKFNoXzOZiJJWemECmORiy4CbOGzkx2r4QKEnlpYbKz1LpyTXUdfQ
HeTnr4NTyhpo+PTN3kh7eyRn4yB33YdPQtp3M88ozEAZAGDZ52CVnCCAl5Ps2TKH
qNpNEG2+rIkxX+BvQJRBFEtoTwbQXwFalq2cryJNng9SQSQdiWkUJVxhbaifdcQX
S/hkUqTvV8N+kM6vi2dmyE6mgxgB43bx0J9T6frWqIrXUQzt9tKahW2KT/43AQhO
lo02XvJqVSQAb36Bu1Lt8AtDEMhnYDozoEysr2D7+9joDiApSEWIYwepLC6vgxPl
d0X7vhrK7dpHMpzHA/Z7TbFwMVFZjBwccvN5BVnlRDIfdZzWx7czoq1Rf0CfQIp1
gx6iSOhuRqWlXVg3D+Rl0+9x9LCjNCt9rYRnORNlhPUFOHQng+AW8gaE7HN+s06N
It0paaWws0ENty96YCztS7h0EbwgXxAnd2VYI+k+0kdwbrDWteh42Cy+Zrz40Dsc
Y1VDPTegr36+9Nl7y+QeSVbVosOfbQayBx/P6+8tTHkj5xYPPgGBp167tYfbZ+c0
p8UYq2gEbIv/J3/Cm2vGu1ySQQ+llDBEE+kq0DR4SenraLG7z+KpsYvOM12N1vCp
L8ge8RTaosU7UDZHducW8vHXaAfCi3Udgbh9g0DmOz5DOwFmugjybfGmGAbbkfNE
25OgGp0LelYmMrJ0HZaAIRdZchuy9dmT1ySmW54WLe3eO+yXzinNzkPRE7rwU+CI
EHa11wqjTD5d8sxMJOykvXR0BJnBNoYXOiOZdywGVikZ9XJm8/t1Ca04ugYUAN8g
JZD0mml6zRMJRdgaf+dzZY2gCKLHi7tnX+YQeTjVj2PDCwXznrc/RtiICrebg7aI
AkmZZG3z4bokomXaLAXxvqJxrSux2M1h+DV2cZrgeeeHuh8srY1eVKJqB9tUNOIx
SKRd/2PSgc5G+s44LIVxd0NlKTKLw71dn+HB68FLNRkFKy6Brre98wTZB3VBQIGn
Sv44WE1MAmY6qXfRTTjKvI0ZkeKQ/mPd8cZz4ifT8mYRW9UZIy0G+KOMDd3Y6q26
PP7qLB/9cFyuy9/wuiE7QeUa+VgPIK6qV6HCZyXOZyv4b2/aTrBcftzuhT/2Ljzw
ahnP1iIH/FlF7+pAhFmvhz5qFtSw23HjVrFDkoiEeWx4WetT8+TI8dTBOmC+Hv4d
btwDusYiUcO/W/mwoVyMkjShaBIZE8GraF39H2RT+0CoA07s8VE23E3VmTbaS/gj
EXuJaJV0I0CpNYrbNnQxBnrM3sNw6pc2/FgitB77tVMDjiZO1AF7mKuD0mqY+hZr
td6b1xhUs9DWXLB5pKhlaugt2NplEmbbary3gbG9Cqej5qI5rfnu4Kmmn3F0XpZM
rn/TUpXQdGiNjg2D0eWzKIWu9GQfO6MHsvfrSdx1i7fIgpz0IFrSP/iW4ULS556w
xtn+zQzi/DMShIX34HADF++DQiujc9efduQmZCV2e86oM7m7FDIoVYCTtYuLIDaf
q+5ec8noQ8//5ORj5LsTVpCjJtVwzcy4ssUNp1esO/qpDNVE1FSB9QefMnAG2xZY
X/VKUPl/W1EWda0ovpJZpFQFmPdLzLPFBHeYxE//w/KsZkEJgYwpfqBMlASMWJbT
UXKjX2kPhN3zM09OdVagCm1FlVll8NYNOxzMfDRYB8My7dx5NgB2BMEcpMmuj+SY
HBRtaEuF5Jcggx5BKEcCACa231MX+Y9sfNvh+IeRdiwXl3tYCYtzs3aF6r5c4OJ2
+O0A47drRnVwHFHzOAPTFMbBA6YUzuBd4VjtMFYrryKI6D8GZOM3axntapQf6FQ4
Nf7ZEgfHbB4gVcj5okKcixTNx7JtT7ssLqrtpVCnqOfj6Or3G2a5Z0x8JYor+l44
xc1vOFHSIhLS4eVq8+TdeEaZNWLFwDtvoI0vZPrq9hx2Cs+5oMJ7fXkUQiaN0YpC
7slfb4SWTOOzxnE0Q+5BmPMPOlH7vPMYeimbKVmAASD511fMk629dyp/bXJfL9D4
7ES8F24mh9GFmY19uvgI1otCChO1suJNNoeSvsThcU0MLk8CKwybyal7oYwiG2+l
nvslY1ybt8tx1PgfugwkcNmnvAdibU2jrzpz11zMRrLVS2tmNWyMvRuVzUSaTH9N
Wm8QbyN+mtd/NPwLC8nNPiPq23xYDuvMjkWFrgEiA2rwiHs0h7t17pK9CmJGkUy4
DM2y6e0Yg7UBKrUtNynbhZo/IpcTMMnHlpkzhRfqWopib5uRp6LO527z4c7VBwz5
PlzWZoXzdPgTultPen5he5ron67UxdB6d4ajZX9fDNuKaLJvyTiTK+3TuK/SUQ8K
cbPgCuxFWVCw2Pja7IIDGhlu03UVHzwpKCS9nH9sd3kRZ/WIhZvL4jtVPpR6ZrfS
0KP5TidIFacpUl5gENNcuUQdne/1u5KZ97eurQvLwYoM10ymi0L9r4KpWm4IxR7V
KDIGuOzR0W9uwoIH/neDz4ly40JJNkRv+F9eXLsaS42MB9KYDmAl3FUK02OLIe4b
vANESeFxFInZYPyKIe/fF9EOVI108urHSB2FVGVYcYzTyONvX8pg4NOwl2OO3Cfa
His32NyJt5hivu1ggggkSoiKAiKlS3drxTLZHvY8dw+JSYWfKVdcoQ06M4lr6XZh
jPxyDndHhx+W5fwH/BIU0KWt7DWmEvp0StweUyytMtAQqbt5AP8XiD9VbpEjrQi6
idahWpsNyu1yOI4IH2TArNiGrQsw6kZVkV21fj6XFJFlkROhXsW06/iuEBoo51yk
u5jtu6MOcJMhPUDfehmhXhid6xCU6A/+4EjHA9XjZo+b4TyWKXULSLsdbEtfydia
3HOrRtl1IjuXt68jsJufwgd0T60gpUgeCzxWrapJOu6IUNr9+dvMrEXPesuTj5wk
itOroO8aZ6viM1RmCPFvAcyE3db0asEZR5IuQErywsICGkSTf1K0ZI6azAp5PdqV
6c4nBGuBdeW0PDQa7ewECXz8qrw3Ecvz7N6EmTO3PwXV+mqh3QUNfqmxqmkQVEVQ
KB1HI58R2zpsueToRkWQTAsdHPWaPRKfzaTysbpJLeHefBzf8RrIRuefqLpXLkiT
HFODfj2wROfi6Kupj6mRco6xAwB25WiEQWo19ooMNAueVdfXvELu4s/61TiYb90/
7Y5PF+vAdg/mWs1atlxw9f4hUsDrJ04HLFcetp8vO4q9DF8EIa2vnBIgSa9h+I9x
/PHJFVPa4XmVK8XQscD/94OWTrjozmLa1Y3VilrgAR4A7a/vFwPtn1wgdqavsic/
MFWzedKJEuRqrwAIUAGOpSvTLnfcdgQ0gJJoIiOCJ+mZIwS+om9wQFaUQhlqT/mH
BYgYctm928FbHl0zJPaXIiXtY0NYT9GpqzC500OuA4yiWzlE1iTllE9kXSoSlFlL
nR4QGAWTTnhD4PbjhaZlU2Ry5YGLEO/ckUAlRbaNc96lmNpKQ1v86bX/eJGtVN47
wAoI4tSmn8oKRRXJOQsTutnL+ZAXJdQms+Cjtfg7kwdxX//+BFeTazwS43xirpCz
6SfftffRw6fNpgwV2N6e0mAOvMJO+s/6QzPoSFji+4sIXR6SgOKeEYJDco5DkBsc
U2gD4++I2mrF9awNYjfdq+0cf6IubVoHGTRqo69jVYK8N7QDUbPr8mIgZKW/5y2g
rwqzAHYpCEV086BJv8aFwsM8ExLTiCZEcMpnQTNyfZkEzX3p22/d44+k4AJtVzJM
LmC1WM7TStTQ8K0suZ0cKlgzgoSGHXAX0fpoU4J1J5ZJ08qhroJzPXj6K8dylurj
7pwy5fXR0RZSztA9QUravBAZHPFsuTV9/BsstARHksR4mmE+i4LxwmP1u0jHJug7
xIGAbm5ANv5wS0MUQ/592Ps4AwThnoirKCuQYz4aNrn9HPwKVNBjI/dHNTYwfzoE
wnxRe3eBUvSvoNb0s6R0CqlWbfK8JHkf7YGVm90f2q+G/Yx9FgzSHjSDK1e/rySV
WfAbiLnquSlP452uT9eNJbK/w6qI9uKi1WolWlXG887XxnZE+kjydUrSUJ5vYH/e
KCit+5t23rnJWQpXKGMntHF4iiIy81kl2PoSnvnX29BpTU/nbRFYw3EI4AaX0Hv6
emcBVgpErP3AkpjiGfbzMAj/MiT5Sp9w45M+uDCVWeZB0BK2rHpgbB+815R48lIX
QNfCFvz0anTZPXWtu5N6dDEcGf6gFePFb5SgB1accW25hjDenZ7T5MqFaH+WXcSV
LcgMWHxdSQa3cukXMb52BY9fFwW9E2Ff85QpHMzf+yCYpLdd8JGuHvn8aFIHSWs5
UG0iTTlNRyDvDF+AL80wLjMCFhqJlsfifVPDQpzYDwVdjuKf9nQFP3zlTiQKMBRf
6C+7YQDFPusDfNpPefp+uWJTdKVIKq1spr7EnOjfT0SMOvp/Up+r0U0kxOQ/kQkt
NEZflGqDG/tBdy2gaEUlnNh9Ta08oqaCg3RLFUtVDRQsFKtRwOs4DxKN5Fc3e+dT
GVjH+Gmbb6oh3Hvb8VrKlyY5ICJPgHyRl9Do2NM3PIC2qNIycS+fUCBOyp9gZayf
McFYGd1z9aYdOcSiMSwyV6XEdhyUh867XjpuNK6a+w29BBuq/LfpN/SG0R5NDitT
228p2NTWnx3DUuScn4IGsibaQiCmVUMXvN+rUrwBhbK99zeEmKj4Bq1RTbfwJO4h
dDEDYlMOhLgELCQHWEF0X87K3ZjCEA3r8L+CDEs7SLVPW392iwcjZ9PK/teCbNd0
rfMdODR5xXIP2ic7TWQmdoxSegToD5NIgBjHeKc+xC2o8tmmUUODmzbkViuau4f0
lydrXeuYb+M0YdFVCfe71Uu98+wMWQe/HM8vSDoz5QpFshPHmxiFXL9LRkr2G9ly
OxHy5ezmibesAErtq4w5uRtQFzywjjwWb4PsF7LFJpYKCls83wMBgnSUpfX7Lo0l
Yw5caqziSIU3CbHa+odDJ9o9TIQCISG0hgth4JpHuliiVEwniovv+vGNoL/Aui4w
M5wBtJUOdMdBrcIyZ8rAmtvvfsdecvZoMgW2+AOKbZHf0dBiUneFoFYzkdMcxtck
+i38pqCBd1avvNl5bM4QZh+lVjx1PO0x15i56PvYZPsqiU7FlwZwU8QYyrrBBoN1
ZmwSboZJ0XZdqai63B8sfdXfAqAT6e2i/Rw35IYuUNXrbgVrt4OeHdzn7bBk5ZZ2
FcTQZpw+uNkiKdMdzFGtlzMofc21IHyYN9PBSznfahKd5oJ+gY3JI6GAQxVTP+ar
KC/g1CwCVxrBulI4u4WPrcRO8RGKf3820Gm8NhLCyaNEaGAPYwq5TIGEM79icd/Q
9++mHHpTZUfdCSZGwgLB5nNb93jjXau2MuLwdZwGLJUIHOWIV3x9U2R2nQn9L87N
5ScS+G8HBGID0omBH1FrUATk07gKZu2NqoyfOusLIDcrU8sazenhwEu6yPU1VpmJ
tB5Y3bBCXRDS+WWId+o6LVxbE4OurUYnG4MCkuE2S0OerWpxVOjMfUYaiK9JF01/
61GHXeA6PXKKRvjdFyjleN9o+88t0LrOmAM8FttMyNRDZUEnzEHLDymtNIWhRbwj
Rs8sNDJQ3ZMFMu/Yti6v49LRselnd1Lcplgos1HUZW8QQYoFo/SlvYoW7JbrFJW1
74rGbttG+5os5pu2FuCUQPrL7vxJWEzVNOp/ikw2rkcxXSgn686hbXxSC+bBLqhE
vcu+sG6tWNf9hezpRFPhLBZ04ETplNdk124YffJMPXZjQ6Uhtv+16cGJ9+FRmM3t
yZ/ebot6a3kSfK6Tb9x6uWoubhMojegnKbACJ0mmdxnffqLjfmywFmv7jf1bEFB+
3f4mlUGnW/ydd8LYn5z14zAEfzpG+BU0zKpFNbuGM8RSgGf8wybT7E+7f30t7fZV
p0HdPhiPIn0M8EUZ2EJUV3GLc6WCpikfyew2fJTZFMTXFpCmfHWVQcAMkvke61G2
T45nYBpvXphSNkFP81fcnaQI3sj9Ppe47IEiKghBqty6NHVD/9YEN7e2pYD7ZHaT
lJFVFx5zjN7a2ZtIYXEjKNYLKMl88DEcXMj6CCkRugT2thtib+N/twdT35ICa6H7
pSD2DUBLXTyeeg8yryNM8++b73ISU9dgzn/N8m5gcfsgMAGYrSa/1LIQiJbdki40
bu2lXeegM0GoKYoCkGdtZ1nFl6Ej7lqeCyEtN3MDzUoVVY5Rygx0c87I0B2O+L58
Mge3NTBsjy2zZiqF7kGP4og5QhZePVy+1dKJHFyAiK+gxgThNS1FFosU3XY+LFzK
h4adJANEDfQsZ/IlG+VjTU0sAzQysx/12uPK/PUdidiUxBh11eL1Y09zrmSrKniR
PbJBtR20+aofUAwrT/W+AUHfP90+nDBKM9ai9X9yLvl44ONPHQ7wA7Wf+wUd3r3Y
1l7VurV/YUg6eIRKuG2WpI6pB8RZtfy9N63VMXEmvYGRX6PvqNU2GdwqogZqUAZi
Dw3QV980sSLmmB+M4eI17wIxXMLu3Q4/i1if2WIQppCaBqNE7+naLCdrU2VOwkM0
/tUEsO5kN/LaCc13982a3//5NGWvJfFKl8m2m/252Jue9/gAYcFzcsiM5LwPMXH3
jTw9ymQFPavhUoMmS2EYQDVpvjyCK5KCK58G4d0wj/PrzKZ8zLhh/3Tmew8XQaF2
Qtgy5PSYBxkEiJZj5PwjJWLT8zoLumH/XUFKPTQRbnJQXxjQQh7ZlwTPbNuzHllh
ItO6j/dltTY+7xq/U6nWflZNKBGXXbYuNYRk/r/3SpnP2ttbH4IcPnhEMIMTzcYd
Q1n1SCcQRYDtFcUkjCu123xkpnkbjs5kV5P28m8Qn1egp8syP7U73w26rV5ZGzqj
7vyLUDWp4A0K5TB5YT61GAZl2hwQnpSgGW/TPWo6rYLJ9goOHFfaS84aICpA4ALs
cOz1LuGIF2H06Suf0Z0TCXxMKYuhwEzpYzrLpmFAoayffdycgvcvdCBpOj+vGKvg
N4hIwCfM2kDPK4Mg4vT4rxFnC/RSYjirdo2Gh+Dvvg2JUF2YzaWRm3wE0Km3cMrw
tSmDUzizHMknWFgUxys+iZQI/qtH598p3IY2I+k4U+uEqUmz0Kj71V7TrXNCY4OV
DeWy1e3nC8k/DbwnaNPVtKlY2L2F8RCfvRpBcVzeKqsDPU/UhU7Jrt1w8gEHxN+H
w4QTIpK28weYbog9kIAGiCgVikLtRoxKAuB3JuJWq+mZWIIKZodqhlkVtW2sTEOl
WfFf2jZvVRNmGrSjgcZsN7eHjLgyA0JZuea9WhiE2AKCjtpA8d4zU/sUMy1uPhst
mCZrKEanOPmnLkW/2GHw9w08ogSoGv6fgm6R8fouwM2+Xz94oqq5lglq3wiH97GZ
X7yBxXbRPEBGgZjRYFe4ld/ny6LDutQowfRawARWp/g17oOj8fl5HJQGTSmEWuev
JzbGZH4vzez0FX1ZOm9r6/oP2hhA29oFjCruFFisfIpWlK8aAVN1owTwOilL7byC
7kCgSk9HLpEMrXDRWXH6T6l2suU9NdlQLoap/DV98iTac6EibGdiFX8hgyRSIV0A
Rumue/vzqo17hvkyawIDa/K28kwH7aBTKOErQcqi5941U0kv2a6TcGxUQF09GcEG
C5SL0mn0lBqIs/g7SPNidyjwkJZr9zeIJvZxj2SVZrSdfN8mKN+8TAETcgoQb6sv
i2eBrhC7ClqLoa55fO0GyUT92L79HMC5t2a/rAnnEsZg+tTBEh2D/QJOiNHQXv94
fxXziNv1om/awObGCOmhW5cyzAK+NO73pr0KdET6zpy3R0aVxF5I/Xe75eSTasCB
30cTsYOYNi+yg0CnYNbJrjBBa0vplz2WSpWw+ajDG9M4SV5xC0WHLJufUQBei89J
Mm+pGedCevBodykqDnPM9tfan+RfWnT67ipjRVy4f0q0VN1+mWAtgNXh5gHSZwUN
/O0k04AhgSBRM2B+egn3xRZVJ+SlEWdj5gnpKAwCRiwuTDwdddFPBXy0MoggEJc/
nnFalbsR3JZtVgXFvM5SapZ2uCnTUQ0zzi2w+EqKQwxYbbHLUqMXaGILDnLYTwKN
BjHOw2wJYjooAjRjd+WbG78496vy6yHFtHmLvWclRkcuvMJBhteZJsL6kJha+J6i
Zuzsy5/siZKUjIDnAM9L79dzQ6hXjFV1iGhqNhZ3LLPnfd1TF94g/e49jOiLuKOs
HYy16KWbI5glTCMTJbFcyvABjAsuSwzVbCPRQlL4Krpod1DqqP90W8ZXUaSvFbIR
PxhuXUbUUes1L9sdQzdg3srahvNUyb6cRIfwS+nmppwR9VVQbveEbX8tJxoQLzn+
eJ5d3LOAz1eDxf6bL1G+rPOnpiOOz+B51GXbaEYtNn3USTnuD9qgbAGc3XUZT2tv
rf9Y5OcVqEYrtcaJDBqQTXjiYnxWZf1o4aGqPQxUghvm1m1+Mq9+VC8zIxDsAj3A
ICOShwxPxmf7HZZbUTpW1BsGorfHC2guxQNPE6TaBdaq4yZf++ENn2k3y4wqTVme
u7GLPqD7yMmCYaSQSqZxUBGa4sKLA2yLjqe2cVA+rSc8z1jEJ3zWxNJTXOmTu8AC
mF3qL/7K7zl0LisFX0CVx1+qrESV59dTAYqyPuJ7c1J4gNbkj+Llm5GAI0u5cwR6
qtGK/9VvLyobLo6ZLGhQyd6YUwYrKPwJP+ITKbYRmaJjput7sr3gLWrNZBXVYdqu
CxmkXJA3c0N+UZBaTc+9eXlh98i0lb6DvK6IERlSM/ahIW4Pi54rwKYOQpV58607
AErgX9S1uRCLNG09064ssMp/3qxC72ESLQsVs1vOM131j23GTSs0kdxPdYuX1NsZ
kLWTvti/TiKDkCLzZ0+Dk2rYh4yc8Hwxrqr0rFYNjcrDfProYxl5zE2rGFDS4kH8
DDuBv3uRqAJMdm+9lphhUR3uUAeoZLnjnU+N3jYIQdTpB3fCSQzl0mXrnXlM7Lia
E7aypjdnwX5nCfUHApzIgV6oQjXFwBA0ps3abHVU+NCbso88MnF95SvFpHYEMCNB
gKv4dMUk46J+ub/UKVzMdPjqdETM7//wsbAExSizE3Izupy1Ps5bN2JNb9Sa4nO9
HTO8/300t4lDyyYIqNhX8hrDZ6JSOkuks5VPQ/1QtLQEpN2En4IMwntIDcVhslkk
DoKaf2Bpby3iG09gAqqn9Oa/2lYQXYic18gWlt3VEGK/YG3JqnWObRa0cnQNXGo9
PEo6eMlefp9f+BYJpIDMnNO5nSNoFgiS6avPHTwVshwUotlWcbmZgJ6kB7Dq7zOy
AhnBgeIpjr8b7sXsyKmkq3cWE0q3Pyq+v2ULpc+GBbdQput1t3DPk+afK44ZJUPf
AGDFrveUF/ppJ1qpKy1W83ZRTHlGtqWK5pUo+F/Axv0SDfGInwxzlr99KXYjFqtU
0IfRPDNF+BbuHN3+zaq2YpS/EcUrRwaKPhjUJSWKWkBD0WBqeECutiwETYbJ424Q
ir+WVGcvpV++YhNEACRmowsd2/8vf6ubT9CAL5rzEISmT/VnI/DUv3YoFG9XITJx
4Mss3JZRUAq2ReKfo0K0GuzpSBebW8B2d6zpziIkz3sekWV2cR1mms77CYeljYpr
MDW9eqsZkZJjwJeAV3jhFFQzIhnywciuGFH2Ek0+fDsd9knG9wKLJfwU+8akJhWE
8K7f548wSHY9rkm+Qyt+O/Tj1cMTPY28x64QVc+boOfFQTElWcULE5E8SV0w7U0K
s9nuXwB5R1ggN8gMHKxNQ8e8slZtkL28emBpv2NAGWBaB5ZOxsbEDhgR4qGKleDq
KHj9tyQckm5RIcy+9mJjF9IipJwqHcewYtquC4ue869b1LpXI5JBtpIDunFX8wbr
5udxcSgikqPSSRq7oUMJvBMXO8AgtOnHDW81pnHnJybgmOXCau4Pzz6r+MWQ8flb
Q2q1PINBQk3Kv3scs0inEfUvPI5BOUeEapxqRoMrlGWPRbZlI1xrbWJykCBkYQOs
Aa7N/yqjLxiXajueH+m5KfsIuea2xPajqdjyFqiOwx6Ofhh7UrUwY03dp0uVWNWk
HznYc7vR4Fj6OIDrJuQHP6t1kiBBrGNhXv3EQnEAXtHTcP5KB9Gg/bH5tmrfDPQ1
a5GPtJNPdJ5jUgZgxIO+cEtmzGS043fALwdOe3zSK199K3NOUhUb1qYMlrrLznAa
3gykotrNgeN+w0tioXXl4COuLyuVRatbmo4lwWrJRDldfepLAcN0NKaDKoshQQBM
PJUTkuRYCOKMU0XrsgiLaOxARQuw5ERWNQ7kpkYKHnFS34hZKbyvXaer9iMackHm
Zrsl4GwDmQZO2IpZRDYPhS8mt1vKYNhNeSlM+yBPh1tWrwkU9L19Y16577sOGEBU
a6okmHcS5RyEhcuUbMl/V8LXLCwgE/b65oyYpKYDZ/V6JQk/PWWM0GQvP5EndPkH
P8GLXq3QVOYL2L91LV9OyJt3ekc/YPwUeRqx9idQz1IEXuFxql+US+gnBxVkQAKQ
LtfAW49NyWs7S6A0yBYm8ZV6wH33iXUHsJygDh1BYH4GFRCcmqxhk3bzHBqvzCmH
Lict2gUbytzHyoNYk6q2SjvP3GOSg7b384d8bZWSl3RsOdBkZlTZyFvWm8nalymj
KE6pyMWEUn41BpjxlgVDRBCDgEx5AUoCxiVbU2QStoAJWCc1ge7AtQQssKsccsVX
P8Pzv6LMcRbV845eJ6NAfPP13JHP2uQyqoQK783Jt2X0xvhEpFcOdsa5BmbdWoOy
F338uURG/P2O2LZzXAw498yqhSxAKbM99fUiT/S3hWSxvbjGHy2v/qYNmUtCEpio
W1vOVJDZaNNbgkjcNHacnWRtFb0URiEc5M4/wCP2lOkQpYpmNlVCXQtOIuCqsh0q
vhoYYY9GFn4aBzpSr9Gq62BDBSjcKrfu3AcbuZgUdU9Pal76jiEGWBMpfTE7iAWK
hcmejxaqdnpO3+q2Y4pYaAlupqh4IGVM8hU2YIPKI0IDgs42rbj6NQcHp/7+/0lL
wDv+/sKuKBOZk/JEmzk86YH1q7V4AG9G+zlvqtwWE7uZz/pbonvcn4JOY4nYUJmN
VbUtUCzyjNQmmQNl8J4Ix3CqM1ImS3kdvUr1KLrjCfTgfAXp+7S0AuYS9XYVZ+Lg
eBja8uQz/alEPMNsD+IKubSWsr4pGBpbLi0c+kxea+AgGguz8Q0HyY9nM+7VYEJb
SwbShtMq7OJuPGnrBc7GZ2homTUqxVXCmMaT8ZKIEiHFEQjiFYIcuyPhyWgEPbnr
BFOMGVs/+QAk07kLsgwnKIkoj6Ub6PYB9LwM/VDrnpYwZzTGf+U7jtziPFYBHwDa
70OkdizOd9Dz4EGl6NYst4d6YS8vvY9VWr3nXP6NBWoWLFnlKfsdZtEBCicT1CJp
aNB4UUHTP46Q7VX2JkH/f0Su7+h4QqKt3LPTBUrupHA7Ke5duMtNOLjz7iWTc+MS
mxjCQsL1hwCmzh6LaOTqlV6tZsBOkVwUswoZ5/sI2IOqZ+uN4uHj9NO2sPckKhBm
+F7NVgapBTxvKzzUfDOyy+4nTlKDLHucR9dYubkOJV6wlDlTJCp+BtTuFJ6i0bG0
JnB4aAxUKBIKqHnTLt1jgHt6n+2iqJmApLpWpbbG72Axxp7W5e34iQ43IgH21s0K
okuVKchHcWDeUIUZJaiU908tQz5CSk0OClYyUPNGyeUqmUBjpWTZ6LkFY4678gQe
xC3zOGqMRatns1A5pHGF5WXj9nreKn1z1UO0cjjzbEwlE4+3ErHR7MI+u88asU5P
htYZePqhd9/ASzH/go7LKdU4451SdBGL/M7N5vEFhpV4HjLbyfS2hrrIjjJyuRPj
DP5nrsgQZAD8DQiYRQbpM6tT8UrHPOlBjudC63MOpVQQw/Nu7bhq/+x2s2eqzyZv
JVgZ812yjKm04wTFSTwM3KpvsoAe9seF4SD4eV6eLCnJXURlSQ+KaepRafL1RI1J
Jzqd/Vgj3EZ/IS6DmqNtByyWFGtaEPGjGtXa5VFeEQUBEkEe4qMb6evhn7zycznc
gldRE4yqDBvC1CG0l4iKl9yOabCRxnMbo8rW4rtuaSZRd4+HtUceCpcS8sKhee2F
Ww0c2wFXVtUvGWwTl9LbYaPF3UGjE5mqlyNxbe22A+q8hC5MKU1GBUlZ78Sy+4Ay
g9Fqt6Upxn644ItSdQOqZXmUoa/ktAxigl3lpJZ85IBQdMRgmSoqzYyUwq/om1We
TXquaVA2yfUTeu1hbRHvFdiRMGksm23/NruwxoKcOrOvkD606mupJyyVcrvBuCF4
M+aFqGVdSqOi0YSE3k3JlCrtdaD/NcmB16nKsxl0SWuwKx7tpgsYmL+7YILQHDLH
MQSnL788cc5Ea9HvFm1zXeTR8kCJYUXYKAvm/oNdYP/I75uHssad/UG5ftvSZgvp
MEdbEvkmxmVFJVf/8PJV6FZ7BGkNkPlVt7+b61sqUd55xX+1BttRUqgOodBDZ/8Z
HPej4PbPqUAzEZhhdh/PQbZZVrC1hJVl6n4F5Za5e9KDkYAnpDySLio3s0YnAvpn
+9+OroFhx9nFwtrw2rbxwSp3tLfZRTuYHjqJqitOUIj4BdGWf8CVUp5iDxnvgFDs
bX1Gz4yH/B3lyIoBSo37xst10qRXVRxBtZbPQjsCOpoc5Xdlr5ccoGtE2kR7yd3o
shT0EApNz6POJIuxfyk4p+tsnU1WLAwTebyzLRKUfyjbosuk+hiY3OvenIjRZJrv
jM607aPdmX4Tj3DEgh7sifF97hH5T8qr7EsU6JSWlZzjTI60JYxnuXH+w6gzoxr1
NABufkJqxu0nMhM0f4R9CA4wV/6jc7MEj7vi0nZUHW0SzZACQbGEsX1sH5DUI2Qc
aVJjL7spdu18i+D1XnK5gbpfCHPVjLTyn1RMvmD0Xi4hCpKZRmvefojhec5m+IuR
p4bxuEylr036hUUAHmcT/V+jueKNA4nC0K/9zD7RJlUzDd2I6y0D4xVOqZooo95J
I0kYYY+DFU+9o87WumReSV74lcnMtUVgcbyxANAUNP4TTCvhnfNUxZLEEck0bwio
I50uL1F7iG/tUiZgdhFF1nEMpZRUXK/pYHF0famSEEej6wBJOwN7tB9cCVB2ttuW
b7UhbMj8bahA7YuLfjvqBA/nTu2cpf1adw2eEB78SFV0mqrKv9FIC/yPJKFeV12U
bhek3AVGJb1NX/D9XJdjF2Lz+c/qyna42U0hHaZ44ncNv5cmqLegiqj38zCGsRcP
6J8I8O9/51Lumi3Z2VK964sogfBuN/YD1OHZgO+mhIFlLDn8vGr1KZgBOV1nKiG7
Ydsl4xWjIqIvDJsLfiAEkuTfjgUlj3mpQnvRk8aUFeWfZed1Zo6S5B82AY4abXBU
bf4f0udVbCupavQTbDgkuxkecDn0aoOsfIG/WyEE1q1PSKUQA7zcP+RS9DGDMqG5
irK8wqzOA6N0SHwJQZlLqaug/B5lznVEZpGF39aYajnnJYUHOT5q56/IsIJCEWK8
G1XkF0O/gmay2HxEJpDxbK7S1g8aVydl8qqNrvyDBNRV9Qe2SJNUnMiOGkX9PX+U
GyicaLx29PvjF5XV0mZOrowmhI9bE0+V5hPKF6oP4M9hzDhjXtXgt6ED64lKUs1K
eivMIfJxAl9yt87IkQJ4ga6sgHIUT4fC7qWbO4QLJRBH4ih0JbQrRnptndhwSLbv
aQYvYqxnvQeeiMzXXwl1o4wC3IjfSREIjRnUEp2pQ77D79nsxFk3ZdMCeBXf4VIS
z65rLJ4JeeJjm3BVuUa0XgNg+3iIsb2stsl4K8ZUpaS7guZX2K7aUoMXazU+OjJs
ZRqdvcu0654c3U/O2SJ8numv3ErFbJjBlElAU93VSVq/Ioqxbyqmt2rhIQ/YsbuA
2Znvx/vAYs78BrysA+Aj+wmjFx15D//9xsJhjbQlG/Xk2NhwhCqOoXbLxNv0ezPk
tzNR1AyLhM+5yIUZLHAQ9hFusra/sqv2y5dEgCJP3Ybk48oDeokRKIjvIuHsOKy8
B9e7ee6V1SJT1xum5JhdeeEb8KRW/yG6JRMkHNuN+EW4KCwgGTTZnUGEJfNX+IF/
FusGbyv1JMpkkzsNqH5MvXWEY1U0+M28Dex7LcJeTj423XYhf4A22gV1uEv7l1vZ
HkWjn5gSSbyu2ziVM7gAaotmFSN6pl85dz7XfLB51ThTcvR5x3QTd9EkKKMzrlfm
SSMhs9/mDNneFxesrh9KAN2X4MwOjFE+BPKP+we2T6/XS2SFmWOyZTn/5K9eeMCI
ZstomS4aVVkzlxq2zrXejp3INh2ojuAUOBPfo1KAK7THij3bWIFqOt67li44Fxv+
0suYGJKt9a07Y80KMIs8el+OiHLuAftnMXVhGw4ewMOAwuIEudSgkjXWofLmXZ5B
JbdsFuTBhcv0GVS1mSCNxQ6uRijGyWDD0+GFhhxxsRuolTCOtE/HyT3ofhxtTN7s
YZ47131d7OuQq7osJ2b+DY4rDJ0Pys+/4W6CyCFKj4/Q9pSgviaxBkM8BzvSK/WY
7VzZeG+/fTeK/mnXIkgrYCClpDiNKJ65BsuhZ9lmZeJWZRUz1tGqiXvIYt/sSUOb
tQqsGwWztFlo0qB2PNTX2pN2jdxYoTHH3SMesX9tNcUpzdLqgFyAzyy0u/ZUd+5Y
dg1IVETp62dM76gZwwDbePOBd6TuVNFZ/yq7H+xIUPY5ZwUdjt19/m6y/HoHmcei
4bi3Fg563NLMfJmauWc6417v4G5p1VudwR1lH4jQLhU3nMwy8wBWW+aulVVaRRr2
UDdMVsurnyIfByKDPDa3biHYY2wip2jmpLVdAW1NtG33s6FxJCqmqqQi5S13mZvN
M/KSvIryQwb9DBZzh6R2tG5fNqgfP5ZGBwbT06ltbDAL3v5VRqRBFKrXc0/UPTEw
wLkrbr8Vj/bpb+wetQ/pgK+Zj/YkoFSp6FIu6sx47r7yFOEY4izxEzIWaHU9eHOm
r6rHWquKysDiUm2/APd9xljKuWdV0Jc5jABy3MTzmMl8M3sLbzrNHFy0JUTRhQ6L
fs5inOvERdlU3WTMBNLftqSobcSQ/KX0tzdHoacRawzdesP7w8o/XEhn+4QfX8Jx
Vh95wIOPuC4qD75qg1cJ9qcX2ACOnzdY1KiLXu0zo314ervGuYqKgjHDHduDHw0V
G52WmY+DlUQjshOYR7vqUfCW7x0GkRvZ18gUEDJuoavGAeenxIgl7oQBAyL7d5Ea
bESRTo9EnSj528+gpi6bwjXSYtiZmpqB/h3A9T/EqRR4aaUA8KJolOA8dOmxN1Ge
jQH4rjgKywIqrNG5Xuh6BvV3p/aChWrl0jUvvyTJiFRZOlYcDFKbT6H6Xp83NU5f
85wo0tvNu+tw3JLOELKwFp5la4hvF+toTQOQB9fXk5Us7FOHFTttS9TKc5PNkeBe
JC+GtsepnXxSpdvRYexUglBlYOr1C2QWCgw+akCRTbdt6amtRJDTu/h9fpm/bU3O
m2ry+HrDh+W00uZpkaLU7+GpNCDK7X+94HQJcRvE/vNvJ6mNqJQZko+SGIwxdY2f
JPr8VBHcYM5yYPNqy6vCs1doEQivlznMA22nUJUsvTs6N+SzlAGEmeI/xEft7vYK
wWjVawXov+Li+nUCRWMONO9kpTXGavZ/oBOrQ2K9c3wrmyQMoFiVwa7F15FsXR6p
NME9pUzZaoBlX2JhEfPVHa6GwgP8ixodJR6Knh/IU03AaqRGE6ovdX+utYfPD522
SgLf0ZtrXDh/Ni49k8NXqIZJdznf28kwUA6yZfK0vBYGRbAJeAIKgcA54QGSqlp3
9ohwyLF1WDVW00cmIDH2GPf26ccMddEUI1hq6mssHlBXSGyPvtk3UDVrfuLjpccb
O/cM7muQY7ww2rdnm5X6GnutNKxLGHvM87S7hlWS/pr+Da29OvzbI72SZ3wKJA0u
8zYcy9orKpo8s7ry7RjRrxP55SfdsjFBR/OujDOixqYo2pR7DaieHGFrEFbboL+K
oeTbaVoG0JdCXgX8iU5JL3+0SrdUXH6nBa/QanBTv9zdOIzGv2xY7Yg/upbInqqY
sb1i1AR1KbzRdVIY34EPptSqhgauUyK4nq9ofMnyYS0/8qdkmPZqR0pCWeD9lk65
oL8sFepUDT8m4y/hOJQxj2so4PNHdoLYYHsFpYh61J8hvGjpnBV0cgec2L4kiNOO
/mdKJyIptDDNqqAO/NDgY6pZtgXM9mxGsYrP17SnZ+bW8ZKXmXReucrrfa0xQ6PZ
5wg2aVFvtac0VhBBVCMTvzkbCUlH9fSXVaytLGFyyztMLTB5DDLeA6PKb5gK5GDR
h/EKeIsC8OF3a9m0KiMxvB4uw9u/8KemHLzoS3e71tuJ5OUkNWOgyM0yZIvJDymv
woQE9evOaDD+HBhMvd8acJCIb6dNweXH0EvvZLLaKQfSf/CceWbMLbvWffZtO+Qq
ZmYcp5qbSa4bE7bCE+YiHi2BNZfLOTzLVf10eI05nOjo1SdxvkNomMBxaIQX6jAa
sUt31+eyL4rlpz34C1kBAd9VfNUg7dM++I8ui4znFBCS1BBsTjcK5Z9ync9OiALy
Rxmo0p7BtJPnvyjAmVHk+6Jtz26o9X15E5LnNY5VQpDRHMqNsPlgqKZRUMHjl3+K
fMaa3GPkyj8hCsl9oCtm5cc8WHUG7rxWsELTRJQt9q5Zc1muTSG4s/rJiuUFDwrR
6AVipdBNAWuCwj/EpJoYVOBfESiXWaY3yqZNXcRMCid4PUo8cbUR8oMip/EwE+WT
kdXWffgKMRsaa9m52Oik/mEc3Y1CDCLiy1MAooSLGolMwguLei4EBHK7LVGXC/Cl
wL2kkRUymTmBpM/zqezsKV/kxObqLP1lZRoVxhC2UJHpIEjRSE1lJ/foeOUvrSvm
GN5H30zMuNJ3pnlgFKOsCwtUXBbkwRJapGwiXRxeDxuIgzCWZg2f2FeE4004K7+n
EkAHAdLxDBq57zlrJAgSAYEisEuIDXmd2mv+RXnFWzyxfNPNWVUon08meDacptag
ze0UiKhwBc64lHegklr5dGoTn4V+PkYxqc73XtFIkAurkzOwVUTul6EbKCWYWHew
0JGM8X+qsuaOIkc9eBREcFlQdx/RsOep4PrcPHz8hWMzj75OTFctinLVlAW1PV8u
G7wep35GjBH3gEfp43jn+30nfYtDs3bOM31P7jR4LR8U7SD39auvFXP/4orqijhB
iDaNk8PiDqUpGE8emI7vOWLzgQ7CVhAcKTkMRj0tNeBWjwtCZ+4Rnefqg7hQboGj
vN5ZeiykrvtxlVB7E8B7j25JxQPCpW1qg7b+Ey76p02PWvhyQgJKxD87IoTBh3q2
wwco68zO1zEyWMAhKeas7POeBc3IbkS7+WsVMTHQ/vh4g359MWIsaCStWtuGgows
8oHqMi9hyJNkSyERnMbTRrTcFXLyuEY0+rK8s7+o8dAP0RxjDgfTimVYO7R7jiPm
KvCfxy6ZGnuEcbzt7H/zffc5n0lUZ8JZXXrmJLsbuYsTuEgH3z6ZG6l1v8rZHQbN
9fiCzK2IylzbF9HeT8bS5do+xjdlRAlZPVUBW5Xe1VfRuesC9G0dvMixbiuh4NLE
Xy/dd38sHJI3QWSS80AyAltjnYNYd/xtk94JLaSUNEeZj2T6si17o6DMGVzkQbn/
ggrA7DFpv61adFylJ+fbUvxfHzaRo2IC2VKihuYyPRKxTfgh583VHghqHw4YLTHj
EfNbvqzN/GkC+0H7nTPeCx1gHxZTn1t+dDhCJQTK6NyWDflth/K6Is+PphOLQB8f
vz43Vj0HkmlA7Rkq3ITSxvNEYeFw+8TyyMmItf5RfNwDppXNXR7faI6xf1Kc23h4
JoPB8Fn8lOVc1fWJ4q/htVN2d0jjxYV/3xoNrLztFWimoxWcRUCoN6RfilTzUprV
uF3mH7soFYv8Fo7AgsL9VK0ZNPOfBMxBHAu9y/Ci/bLuOHH3KfmeNyy7fW9ZGyWE
OSi4Y2KBS7WUWxXjJj+QnWkc4dFdPu9PeGB1mgxb0dCRNmwIHMubOTbhjqsqsueC
9Qr4BmiBqGHYH6vQ4CSVn7EeK8si6RJZ/4W0d/7IgNkLqUPx7YP3KNj3y1404cbi
/RSnbrNkwoqvpF6ODzswMxs24ust9kkZQQFAyOe+7lSs7B/Ik3ztsrRszT+nfbsl
M6E8tmUIKfiQEdQ5sLA9M1MFTiPtCQwPZAPirA80zFm0e0jlCptM+vOfzQLABjdE
nFwMP/ZqDoIWBNno7U1PL0hDqkeilX91WQ4RWklbVgzqQne5V6tlY3Y9mSO8NCeI
tgkTHEJKlpmVAQHNeMrfZYmjxVEAiFA7EUC8p/TpoY7SZwrRxlcEa95hSYtIsvz6
n56d0PkSEQnZnBMEtGY8zGBkXJVe5bOxIod+/wgLrF3fGBBqpzPNAgBPueFQXuMu
DHcuYY5J0b1dydRyzfiCQog/rUfPFuxUGZPhQzcbJ/3HTHFC7h9DLr8JS9eD0ZDM
soIk2RSVKQMB1kvwIZukGYKcaR7je8o/4sBM0FtdjbBIot9iP5Aw9nwf+oM9fs1x
ck8pqYP2LkQ1kRYStZZ3ctcms6w4TjLxnbmGqfyg8fqcI+MlJLde4/UcHoX4ap/Z
Ijq3Z4wFnN/ZA9V0DlvTeGg0ehPvUIo19nZraYQe29IATse+MML05R3PDR3fhQlX
NKc3YlAN+CvdunRCl838/3bRtg+4r9/3Z/l6UxPSlBpUhCptbEjUVNXmLhxnEWHP
mfty9sMYm/3VWdyPnLlgttw878k37EIPCtuQ3jmYUc/W7aACew9DsqrtumYNXjBY
xMUndkxC7KDdR2tEET1iLUQI5ppK29OPfFNhyEx011Au9Wd7AhKmKe0Bz9WjBcVo
ll56bNvMCuaaINCNfdHRIS5tzBepHOGjV4tJErJMMN1CxdJGRLkoCYveciDOUD3b
fmAdXGKriphQfRBpjRscmxgMGhIgLFvKEwshqfsPiuQoL7i55SNRTbwuwJM2SVWp
NIHC9Mt4239JMGek1u4NNy70kxlkfRSvh2AKy/iQRcZLZ0ozAvWqbfY1mZ/wFh19
OwPUfuN5yPM4zumsNPU6UUw0piVHKAKlDJzoHyebgt45zwlmrlWs20ZHhUwWtQkK
IVM2yExgPvwa/KE31sTZyMHASWaaE1NLZPlsmfRtOfXR8dHmAI5bVi6scQ/s1kTc
Wkd/N9oH03PYy06nEOZIitP7laJxlTOKYZ/kila1zwGFoRWkEoh5rsiPPW1E+mqB
zjd4hR2liOGDFVd6sUzq0jzfQhoKhidDNI2BKOURbbPXQJR2j35X6Dr3BBWQI+i6
tY714PMOR9fiY0jdMKx5ZxPJKasehEwHKPrTKoJWgDSik3LkaupKjZ58aSntZM+n
HVsI5UoNYRiXUmG9dpGoqiHi33eTv6sXKRhc7RFWhLJge0QM3NbWXOqTPKYKRr98
2Myc1nkWvvp1x+OL4GITs+S9ZGqd72WpigKqq7DlJw2/AkqeDYP1//Oy7eyOwoTM
44NCWezUOlo9cbLtTsUnsNNBPZ2rq4v5UH0qzG1W9XV68Z4K3qZ67msQy+N7UQM1
76RZk3jBw6c0tp4rjE7ATtI6WyxCgRKV0Bs6hwvqXf/lca/4ISQtbPKPUX8kQo26
1Anf1Ez9xmFvMH9fpayr9f49OEwwlrD+vTRS5ci830RgJeeHSzECGvCe4zqeCSzf
hW7g4zTFo18vjwSHeBX/QcnnDQ+caoVjpjfTSSAyCaO/f/a4MdN5VvLns5TuFxJW
cEeNH3fm1RluilHXlPfqZ1Pql0U13o1J6o7FPzsRTtIQ4QNt/JTefYP5lhViMzYB
3hQtVDhsooDJ5g3lb0J0Ny/lHwmBIcojz+zbtkwXJwllWaZbf5cBhrdvC/Fitrtd
jM4nyAhwkAfImSj5tHf2pxJ4cNCagmYyGXsLT923eQSO9po/GQkv/eGtEyVvy+dT
AvrvsVtUrfBOeRTkNayz4FGZBeJaX8NDFqnqz/jf/crUcQQuXiu/JBJKdRuAZSRK
ptW0INEPD6ZSJAUrVQ4r1gscIsBPwZ5Bp6zk584NK/9DPxqvrdIp843aqxtaq+T6
9w6j8REx/cvFbCRTlcFpUktNX0V0PCO+x3wHBI6FF0wyqIg5+f4d4naZ9bsukTjN
X9hHM8CM0qjNQ4gB8iNk/0TsZj9thERtRHWRYHo65Zuej6lnCNWFrDFbHjkMNtPK
JfaKNd/aayfRZ1TQg7B0ngw9bMJV2er38nDNmY63QmuzHoFxewu+IqBW2orCl1UC
HUR+UZjon4vY6pqHpTsKSZ/Z67yaN+3J/HjGBltpcrSnCICT0LCExdJb6Ea68Iqv
ZgvhmF7Mxr2fQFbv9Wty3fV00e99AePGenSbfUAQWHoGeDdZ3jU3S9hMSiCENGh0
s/kzBfg4aBreQRFfR1cUDCVgUnYM44wFn3WCGt80i3TkNzIjTuwf4EG5G0Prptkt
DsF9Fwj/MJR+2FnpoEt0hJDj9wGG41vdPnZrj+uovXbCT9fumtfRp3N6RKZgPTgo
N+Fb0QDwBga0Uw/23xwb4UNlseUGG81cnUxIF0qQI7tK5XFbqvV4/eeGrAKJb2NK
pFp9qUue1bFlheL5mdCRYPxMNTsEXUZJ8kXZylmDQh2fwXtJw5a93+KEhyaCGVky
kMvUdmL5bDG3kKbhnXu/1AkCNBCOaQfEPMMDHOCKY8F2ssyBcma0WWtX/oe2lufa
cEd6BCfoXqDjJoXNpDyaV0GJaRyzHCNZUBfWc2s6pC71bHDLOR5/NYZvpCJrM7m3
+agbRMxYQhBevkcyiLEJbZdh8f4RmOlTruR1oEXO0HKbhMS14qvsrYIveNal2hHJ
XomXk4NaqMc3NUGYrEw510HDaRNg0sEHAAupr70mJkz/CQxj+ADIlsyr9x8BDDS3
+ZESTkok3GcniMyxgqh0hrDsgekKkIn9P71gsZB76LApM81TTAKap02kLLc8LKBo
OqBMlDeyV2epufNAALZg5o0Vmk1dpxgAAbZzZ5p8e0/Jsdmnm3p3qFmSBz9t9O7X
e9692anrbdFAZpNhPm141FAEP5qeuypnF37nmVNv7PYeZ0a/yZrBNEfAgbcJqown
9l14uEjsxJWlXgOOKbHKCd3Gq0gGhkeaEAA3pVPvfIcY7vDmY07YMTpUuqFILUsX
k6aTVXnqRLQ4OM7ssGrmPxJ3/kr/HuOvVFH17YXvG6jfWcZQU4KD90vr+LxBU67+
R9qnxPGHH8i6qHCreMx3+2sjrtldlzegJhgTPfhc1pznXtBqufo9YSnIdrPkhyD3
8CpJQcXUgvvIQBkB/Em2zLYbU1T4aQE7KbYcmgc3G0fWbpny7G/OTgCm6L7J37cG
vvtg4vZHL+z5EX5d6LuMdq1jLdPXezGIZhR9FGJcm9x0nGR1FI9MFvz5R3jJXcQH
2SWI5JF98CddcDHQh/34jD4gJXSPta9TeGdQfxnVtXAcKovtmwxNbSQqyqwvSsXn
OeScGo4LocOe6AGgsIx2gnezBeSpwcVNKmc3m2KDmY+YqbILW6dSICBUg+Uc3sOM
I5Lrm6HKdrB+LpCkeDqBZamy1xA3+It/oWYiW3VZARgzPjqcAZoz5Hwd9Tqz/fJv
nsKJ+YI99i6OgQkNZIPBpPDFsbGcmL9IxEe+U5i4rgmLRVtrdQM5+jHE5BXtELC3
oq/N63svLgIcuv4eAzeBjXmUgoW1TS3XWp5Zfq+PFkfoY/4cfrfSbyGsvl2QjEIX
/iBaRI7mjswTJZD6PN37i8bASyienn44TNQOajbx8aVoCL2Y6KVNnfCwSZZmw2W+
djLBXhWhtv7TgkrGNruuDBkyHAN7r+MvCejT97bS2lISJiX0TM8am4NMrhb3CLGQ
puqHC82uPcAuHSkjDppfW63tZ4t1oWbgKZkxExC4rL5Og1qC8etFoodmzi9G/Sy1
5W9xLcx7lcaRgk7Ep7M92fKBln1VJN4QDHI1+RO+JgrdEpqC2gq4NeyyqfgQRLr5
psn1/+ZWRkIJ9NteJvg+YhoetMVNktNPdsicgW7sYWCoDewjV1YYQiNE8ZaDTwdH
YE04CNpRbA2rmbjLpxnkjZTxr8AXkaoAnx6gJ9INs7Vh7renv4iGTj316HH89wEU
kSDWXrAO1fzW5UDVobsNW4eYtQo0dIMyKa0cgIKQ6lBEHTe1notF+sM19d5QCMCR
NzNoeOT9CZ5Gq7DNvVIMbSqXIcwKvQFGuxQthqnjfVQOfkBoGbZhL7sbx/FrDssP
sucHLdBuULmoxCLohIB7SWZv6VDZdAS07FYtYgF8EBdz4mpFlyMre1GVuSW3DqMt
TvoudCjZ9ScHoGSHfOwp+ejkg4L34NAb+9Ay11SeDFV7AqAPtNjug3jo7uCTpq5B
3yw7mLHOFkqZGYOn/fsNUKsivk/8d3tvJvBvctlcR4l50CtlOUlM6j85crAYeOSy
+8W5sYU37ouX9YuLnh/8kZWF6m7szFCenV7/Jn7WJ3VGnb2BfALCScPpsQZByTbZ
UN87YgrzKzgClIFIdSv7NLVrvJ1VN0PlOyaQ4AP1eNXaZy7/ePThIeT1JbQdcXa6
HQtFbSxtcWKZ8dvhr4UjomT3eXTlJYJgsv8IqKyRF1g0ia/xsa9x7eIXZAfRHzp/
/UvcfwWmR6hILIVKEQZAhO8JgYJ2dJs/760hFefUVBpUrsY3x5sU74cheekS7j81
oab/LSPfaUH1AEFMbwMYBkwXwy1W+b5gtIIUJfIj6gqFqLYBDtV7Jy2SXVvuOsWv
zd9uNKL8bk1GrFKxEfqnIG1ECncJ0ROVKo49lVwNmb0OAdNPvYslb1Fuezsi/Wmj
HHPXNa3nKDhODpPH8BdAtgyByq1i/DjhHy3Nkr8ZYRpWe/7Ku9DzdjMFlmYuPiFh
zpRxyZH3JuVwcs/2LKWSNusK8u8bCYpiZeIf8lBs6V4p2O9bltstZOBNN3XGgRty
twO5FdsDlGhMz5m1fBu2T1wO/PlwfuSSyuF5Jdd6khYG+/uKpSboln4Zqzyt/aKg
c3PqZyBruJdBdcKtEOxQCq3Lh3WMuyJxui56EAkWg2MnfZoDkaouCDHSYZCsvU/X
UgUdi3w1RWr8a9TGtbgDy6KisbNrEdf5VrxCJk9DwoR5Jf+PqIrEnRipQEvsngPG
txUSKZHlpif9GmdyIWBWLa1lo1I22KzFtfMnYJNLzywXPCEp90I9jDvBDUKIZjX4
6xbPb5uamgtsCNt9fJdsIXJagNSYHiynECqrZYXTg351xFQ5nFvBq3KYH6V1PTEG
0MJXtpjIpu/fwUFZ35wtYyfOJAJIA+qGxpEd7NeKM0BsNOieUZ1hWharRP88wnpz
WASw3YXaCRD4NcATDf1wUp0KngvK0+DXKqYonSxK03cAUPhIkXQmjyJMfN7QCawR
3AgbsyXaldySPNjVDsUPg8/wsjq4tRY0yHbMqjcXjJHmzstNiJ0xCAIXA99AdBmI
OZVPXHD5l0m1xPiFeDkacD3kU9nRWIpyrTy3WdAmQy0Q3Q0fPMwIOl6QQ8b1LC9Y
L0TuRy5yft1goNnyEc4JPUQ2pzJStOO5p+qqqmIFkBR0d+vi8H/H2BCX7dLHgJed
WRtRz3c2xjvNQ0y3F2z4tnnOuBQbOIYB9Hu/JJqWsZryRphcdcMZxlYG72X3XKlw
3U18q4ePkEhUwVV1Rx0Ztjin5xPVfAVsvtPdgY7QXj5xHV1aT2V+LRZ/dTg6TeiN
Qn9YJwf9NLDRV3RQXtt2G94wXssT6WpDDMRj6qSJZXMkLXb3KX777DheP3TvpUyB
hCab6rU/Q+LOEcZp5maefMQqWb/TCo1iQi6jczTqXkYEWGff5BI5l9pHTAjaoXyp
LGjgevmuPrfHj4GUyAiUsNLJGFM7r0FcTm+f4iTON++0ITb99+FokKcEVgErAQhU
/DTwDgarHTHdPcGlEn2e9ZkiDnfkAuxcHHGtNVJuQw1RFMJ5QX7Mts15o3o16ruc
xuKgEAmQxFSWlhfoIsn+h38x8SSxaL0oZaTcpHp6UEujNxmy67B3oHLF3w191Qhd
Ec7dBMd6s65cYmJ5g2yDdjQv2rki7Vy5pH1HTkFlqazFwOHPCfXme6iGYs0ztVov
PEG/poNFKAL0366N7deTCD1g5WaMQqVjfPktVL4xHPWToJ0VG5tj/1dDaljiI8Iz
enZvI2VMwR7tLNB8GEN9MtemqbgKkHPzB8KpqwRy3bLSOUMrpR4za7yKKxU2sEkp
troAiSk2d4We50SHhh9RIFtbCkeiU5JhUKpHtHrLwfbxdf3FNQjgb+NODTM/8Wr7
e19uKZsrIM3xVYGZeIlPIlUC034mVjcO7WjXkhJw/vSUFSS80b4/ep9yiH4JFmZW
I7+XRH7uG7iN7gJSRsMgP+MomzZtQGfSqc2cWaW1JiB7etGnVFqlbqLEzopwKtca
qkMrW+y63bwFy8JvWNH2KhV9chewMoNFVdKCHx5y5kDFFAETZ+yBv7iqKg+o40SX
+xD7YTFYzMuGXJC5aAadT7FK6OCNvyngj/mjcYdT5FDRent4V7JNKJHEBO93Ddp7
3gPhjRj0z02XOXtIPIizNyJfW3QuA34meacnNHK7ewHrVs4fX8uSVRal1gGA+lAb
i4X8rxZzDol0lnQPspQwGIqH3qsPteKi1GEL71oxnKi0WPOgRyR75pKe7tvVhMIh
lKWC4qGeLk6lvcrJdON2wMV1wiKgFkQ807f8Dbak/EOb2Dhdz+x47nQWop3gIn2e
afbhKCbvSbeJpltORwURD5Kdtdjo4my2jF+tSPw5mF7QJm7Zn2ejp5yzbaJVFKZf
ECa1SlEFPZKxe3ievn5diAPZGs/kaMyUPiNtN+3AhNl8PYAmv77v8BynD2oMMqrA
JHUqq2TgoLW8gmkT5JvXhGgJEf6tsPylauS+bMeGHQcVVNusoYL4935L9Wce5Kz9
gYnw7FlVh91Wj2mEpklrTumxHOlUsvZEC0irj9Ry1IhsIwrjJCcrugpqfPpZ0dYN
/1qTNICPIEsYE8bP8KjGgiGn/S7LBrKbvt7UCgLPxTpkPYRTcfI09g70v+fhWbfj
xDxpEQEor2o3vy/EkZ0kf4iyN7GTVdW/6Zy63shnGyfYlqaOEHuJYZQEv95Arjnn
AFSp4JSnI9UFvfXkxQKhXhLpV7LAXaQxyxhan472HU9WAb7AJHYVSgCJT8MUfbUD
CKBkZWB7Ms7X3vbB9Y+cfD5MR02Tb5Syq8+NplNNTBgD11OIpiwn8EiZnEu8X67P
Sy5bEWwlKTJk54tlTJ/pHKjKjONAj0mk/woAJnmvkQJ93gOx0R5t8CvG89ycEkmJ
o39kWHvrqlRzUN45+rq0IU5Vr7myWrZIaYklb4PvZlRjUwWosu17bDAG5vK2joL7
h7RRx1v2A/cmImx2T/BFteA80NQZuU1xM7yxfa+8Nxk8cXekbSfEV8+bIjIF98Ki
+7U21zwMvULk65+CytRvdChHDcygJgcVkEa/s8mYWFneLILaELFMsAGNTK4RuVbQ
idn9BRqaNu2zmUiW1u034PBZkyc5MoxZoo5cIc2CzHdM9EW5zwhFXxnxIvToQuAW
pT7gFZ+JPqYyvoo15BWWJGdIwXNnyvQpaV120KQjwQkUMCYo/uZvXKcnoVL/qyV0
R/xfZEKGmFNsgd5K9umjTSGSCcE0vlcQvvZmTJ66WTfBcw312pd1b+eWn4zMTZ9T
0gDe+8fpUc7YL3TrkDQjfHXhX8oeYvRtUd+UnrvvTJ/0lljWJrGd3gTsaP469hJo
uuNCyirYg+P15OE0YOllyBM3xrmMd+kDco6QyjW/vU7gQkP7hwCjHTvXsby4uHe0
9NaHkn5LKFgT6qfrBFGLcgtVxSKn7p1u8k4YdKE4sYJqgeqzxJrvXDQ3qRnITATb
uc07/CfZAZq19kdLFzEhvz4rn4g/wKPh+bGb+U9A3UATikhtD3pM8r38tDwwUWTA
r7uUhp7ku9lrY4JFAYd4VP3F46pCVIUFVWoeQCoky0Sg4OZATjc1hUZfhb7xEEem
ZDQThrs1Yktc+1UOtSMpH0uFmoRoww1AG9nb+5/Mi6BoZTCbLo+lB9MOMBVvUoDZ
6ks3tSm7RO41+9KZLUGM3yN32m4qs5TPSHXTLEAg1SGXiPrXm3lPLK98Wj5pByHN
kksv4ZcPvlEFvkBzTzZ28rv9q2VCEzI3BvUX+8vmK0Aq8fApt8YIFdyjyJDOPKvn
0v4F4HUw3lFwgwh9n5mo3CGLFP/CrXRZCy3+X8JCqBIMObfrqapZ14ZoLyGZmJU8
jqYZXXY7p8jlA/59aUh+E/3sJsMbdxs6jVYvCThPC/C7UHIX7+zpzkQTOUc3BrJH
/JcqbOIlyyGpKK7Y8ujPNrXISBCuEDtyQJy9u6kFpOxEYyfHiLOeHV4ugNhfIhQ9
SaH2BUj6eJN+8Sg9Wnx3uB9qbE92ZfD68MbRgmN5r96+ttOOEGdP6Fw54c6QQsn9
EmOzDAP6Renl78XnovK/EAeQ2EfJZZSGJHh0fY594495vyj39ImWXgOk3HvJgMtW
uxYwXx3hiqKoQ2Yzss86rN04/khAUFKjgJJOpC6Eo8BKdYgmZLGk/To7GRflkNh5
yLkSUgNFdYGxy6Z8SZxVR05vTHKRY7Q23XkOg4IvKSSHf9UQTu4Yt9Idw+yiHwRa
N/hYUGW6aKi3e/DeZucpukzj5FDV4PSJO+hK/2FvZndX/N05efy8BRcWEhuFHg50
9lqalVKjkIxNbhEunHN57Qgjl7A0MHLlqJ24ldZzTKqI++5c+wzgfPI03sJhdL/0
ZwKwrmlQ+AKCC5EyVkmX5iCLnOcytXmjT44+sbfAY3i1MBVYKm399nRMbDeinQhJ
Z3iM+lLG4ZAn+mnmsQO0HmhWJ2aZG8beEjJA+uEo3CiRPyqU65+TdqjeADF3gPpH
HqBLd7MPjF4dxQMDbdk9ENU/XzP+VrZJ4yF8rDmKSH7wiGvspYrzikEck33kx0jf
aGGvpCGBKPirl2PBU5yeMlDZEu1l1oVhstC4R4o+EMurCj49xrELD7bpgsJqQULr
3pgUxGREyxH7VrFEsBCmh72dItPfcUd2pe1HjMYRrEidkrhUlw9K2qGeMO3DbpVv
hhIr8gAV6CNgFs1K1L81gChj1niD3rNtNaoSOHIyTKZkgUxURPmdvxaquRXDPoWL
56V9yjiTEO28vgLsOOBeglvX2pnrJdqTcPTbgd6qb6t7nfJHmGBU4h3K5H21rLH7
HICKXGQigyMLv3OZ0A9m+QBpx9PWeU4R3IyVK4Cw+DqnqO3Ukgk04bXpRoR8Zw93
o3yG1D+BeVTRw02/Cg0KBMKaytnf1sGayqpuy93lt8DRgvXOXxzDMVI/PKjIOvkT
NM710wEXU44M7NTKOooY6zb378Jh7zS0nvzY/pJVRLWwVvaZD9qFZDj49JKQe2dF
2GbAqvBiRb6grIn5jdwOdkBOstAA3J03D0egnSPm+kjC+xKTd555h4IausU6/j9S
EX75qUMbWErQxFbNMuB4c6VJA17y4aHTPYxtftHSBc/h5qu688c9okNP19eHe5gf
16inF19dsbt7J9wgLN0siihhyGIS3hg023wiet6qRcjqpbK5vgMQjxHe9Opy9bl0
dBzT4cinODp9CFOmkk+K3Jgb8LJDmVy7ULX9ogD5HzlQ12n+44QMdhek4MsypgV3
eKcJuH7zmRPG0vqI1uNaxIBxs1CNLFTrSROvmNtzWfTF36enhpr8gZV+vJnTtjRt
EpU9cm4h37LmcvQc8RJ2vdfx+FFZRM9NmJeWhDRQPyNJnCyoxfcczNKC8GWUKMFN
kqsrtI5PJ7pqWTtAlm1UJg0JElv1T2zXi9og8ngAUsKYv/Cr8DgGADp7QvwBQjBU
guJNZGwp6GkjgXjOflLZGT3FqvuI2sAdzYzeJkULondiS7/dVmIYqShJntJbn86I
FdRZFdbWMVlhyIYnltrgsDp08bwk6V6qjofwdmKpomYcZyY5IREoTZSgBkIAAwfd
0lcIJ+tbgVuT5hZg+umOp5VB6wQullVkESax80d+SRg4cv/8sHlPXIOhQQVZlHos
rG35AYSsszAMa0ap48Ax7Nxg69sShZuOrgx7ZQxQnFp09a+tbc0meoDjrisqSWhq
jVvpXwZYxH/6pAh7HCo2BUrEvDIageibvAZw12IXbg1X5/4ZXZFxJkNiTmZ2keI9
KQZmPuuBVu5YpykyMnLw4cgk8TjVki+WsUETpQ0NzFgiPVidkLKWQ/QmIqXNLCh+
7bbcegGVnl7UOh3tUFIck+16Yby8QBbtIomhDPBafbF+L0kd3a132MCJE9rEQdMd
jk1rxNlzOjj6ken6IQuXrOoEVZ5CUmEVaoNET6l83o2VR6CQ/50izlOIzuTpEUso
FrA4yqLNioFZCwAtT7Im6cKhudUvCFEGp1oXR6lqOrbL6tmt3+UIIUUchx7kdDAA
MN0K3zC2yWMbBAMHCl1weTNqVBMn6Cr+xnpE5obZacBH+TMCaTXcgBOwRv2VFMEw
GI+ebPJZyfwiVgdvxYb54QLiidd9om79SRszRYRRqczYvx8LH5Olud9ygP3nPb+x
B3yp+O5QlkMTRjACP8wJB4+sb6j2T6vMapn0pzdcDyoD5Qt7tjssyHdGvk0VMffM
/Q0DholpW5V+qyujC5siM4e09jCJaD0FaPvrbcMrdg/QkKnNGEru5vZq37Ezr2UU
2XCxmjziOGClHQTob4uSOABQ6O3SQqj/+I4gmjgbkWFLFrX3ID+nZSXL4LoT8dxm
3oMtYQlyLQkq+qZn04D/65VS0Dljh34GLcP01ToyYpcxT+xMZ/ZYVGkQDKY+toHH
09jFu3LwzsGfuiftx0zuPQuouz8Baf6rp72IFmYHoi75ewLwE30u5H06asQNLPW9
OPXWsHym+zXHOMN2bZPfY6AnJuegPXpVq1v3jkXda2NVurGxh6yZX74J9GFmgAed
ER+FzTQQkioOUJJN3iGZC7wm0joAbesig4puhW5LxqJwG/xGeaJeQ058HFoJv2fw
4w+W1+pzlXwRkuaUrCuu54gF/Q4N6AWQfHaPW53HhBoHvxfNOd31IngzBigTxP2z
5B9NLtNjo6kRpCbsGF2E4FHuOSDsBCvOHrZlKSxPNfOJ374TUxIWlZcOQuKaUGwC
94WrPRCeahNqWZaV3SOdyqIJyKr7GCHjCMXQzUBql6ohzGlov9MfFWAJRYOFwOqZ
EK2FZh5JjUO7Q5mrn9d7SP14Ov2rfTYR1REPzv4MzQ7tcowrDYj7GxMaPOEr80AW
alXtOPkgAGzdchT7aT5oWZV6Rk0oQguQfAPdnCVopzYeszpaem+BvP6gSp73nJqd
tbJyG0r35rRxouXhbCdCp52ZmKUfdoo3KZDVHOKaSzimIt6f20b9v8emM+L3WfjE
j61SXnX1T/FRoiY7k+VbfquJJ2DnnkoRL1AtaxVVir2MIBqQAUbfd/W2pU5fWO0S
cfZK5VlKDYfXgxLbr19s9rVaxWNbsplZAGEOIRenD5iP8jmave7IIJFQlBJL4/eO
/IRAzOZNpw0mN8pOZxfeSlYlenWEVOFHzJ36nKENKfDHPkpBK9txgsoDDamak6gc
/SQs1wiHxoPI7GJ75hrTrVN4kqOTf/LvsFzlmNO6K7L2fD3O06q9kTH+j2NZ19V6
kQsPotKZPUAwa7YcYqrxqHqPazW8566biMPSaDXIA5pFtDuq1b/K5edXZCF5d5sR
bH6TaWSA6/QVKAocUvAtArlhTWJhdjhzeAf5tIKGRRPisx9xhK3QznycEVfnrHJb
rIBQqBzpK6+0u4GtE+Ye5BEfoyhw1Xvqxei51JzEHQmKc/uOMB+TaApdejkqJgF5
a3wHNsFDzGwTGFkyGTBnRXZQq+iwi2nrmIxMyyXUrxLVbI4+L2Y6Pdm3iuKg5+XJ
RZ14Ie6rRocLJ65w7NpG+RgNqnj+kJgHc2fpfNs++Z9d9EkR2CAwE7GI96Rx1aUj
SxoHX8psSzXxnplEHbIgMmt9hgaApCIvP5QPbby6WepCD8Z1dMTenEbN+QUHwRMX
taDuqAiXqrbLO5/9kMvj711XBim+QpQtQE8GvxjkasCvvzIcdSa8ZLsYjQ/Mz6JP
oCcMaZXWrb40jFxOisri9ZAwfvGVllYw0qnjnh4IuOzl3LudFJ13NKF/Ss/Myu1k
PSyuVKvxSIlmyWxqpx1jeXlzoWKGgmuTwmmrRyaL3jnKGu4QP8oRQktxUgflX7kY
jFXs8AdXtNmmIwJbPIVxoS2KU3C7YpB/ww6F7m375i8zTMD1VgBHTkLR05TVL8iD
MysFGBIPUv9vDkalAQeD0+ByWx5MKWjvkhMvVoCsKYEfhP7U//pUxJQtcaM7JYAv
ywf+oWD4DgIhub5G+JiZjweNSP9dGUo0byI30SLGIiX0yltdnivNybl8Vrvl5PSs
2JExyHxkd3w9hQLh/I+C4nloaVQWHC87ulwgcXuXJ86AyElbaBm2pKbJpgpZ+Cs5
RlH8lZCDYqGwi8q2LUS86yirouQ7zQHF9O0h2ffoMpvxkhCDufiOiBAFwWnSDvE0
TdwkPr/lUZAfS7p3owK+IE6NtNgFvtiiS6hSoTWrnK1SrENJITP0iVXPab5A5p7r
VSzmduhj4ZfAMDw557EDazFezgksW9mQ2QVFexGkQm+HFq3rXAvPbyEGcni7tntv
O8egLZ32nwtJjXHqI3JcUvWPTxYL2IE32BeBTl2NgTPXeNLqlAfwt7IDqX3b+Vdj
YbcANlWxf/OetAXR8lj1c+AOOF2ClzCEPY3fdm57lINkrhTKemi0GM6aNzZnKPZD
eQU21AXm8/xlBgxcfO+/vih/GUSFL8rhMbSugxuuxV//kOW1i5MPqPA0bfdGOvBN
o42OYYGwHtqlQOlmMBIjBKskOdIqPgOAeCxAn7d+gg4ogHl+s+rR+orRq8E9x65p
2nc30a2xB4vVHU6sP5xNdGdZkqETcxZ5qKRh8ISUD4iZlu2q0iNvVfzixOKVyQAe
ZU/l2s1bVHj9ACiPy7QgpdJgYyolic5JdcQl79wDwVCU1aL5G0pG9UWmh1Dqm9dB
jxM4twzi6a0VoR13g094U/BuyREDblSAm5Yl1ARIbAzvVL+uENJ9U+uojKG/LJrN
+f6FZ3v1XULLyzYjQeEVLZMfh/aK16mAG8NBbFaIJb8IkgFaLTeNnxZYUJj6kqxS
ATmSZuX29pn8g09yRfZjGBq9H2erJnICaU05bpQJKhVu5oeGsvHxZVSn0bh5GlXd
l/MtY/lwKc7vkHqeRjYCxHtqjt5NRV/9k+ITeLHZTcBLYilGXw5zur+yAarn7IN+
5XVzyg7XptPQ/KM70U6oHLvah6mWslk8d4Y483mjlBVWBMmQTP9SFKvFagokFF18
JPmDhcEzhlqWzcTgrdm+zqpgcNkqbHpTMt8SWwJ/AygPDOMIE4HWF71lbKObI5cg
+oA2gjughSltBFmqiRbJDdjrvwjZgigScO+vClGsjsPnOCI0ukxNwHmWG+uA7anX
4lbEu9PoRYX8PMLwfBvHLuwOVL4ch4/064LLNyBU/6fEPuxDZwb0ZvKTE7SsW9t9
NBQSs+uMMbnb/72lBIlTS7BKm05FdLge/FKOyi7QLAHqxJ35ECqGFzQvta8mKwTF
PE/m0M+mhnieIOOiOKCdnopD15uDQHxyhQmjrDdfRcCiPJCh7ZVpNLOPBMzh6heA
BF9nKBxRWbG1adlN4UbNZJMlOu9ikxBY/pYDlpy/ZREMyZXcCDKtuDE03v6kH7ph
m6+0Psw6EzkejPLKEAFI9t0ut565WPIWUsagt38XRYU7Y3kyIh8Hz3F7hS1KDLkC
8n3lH5qKY/KqDdpEdBhTUc/0eymeZQXm4mxoBDuPHsBR/v/Z8apOcDJkDSQRqp9z
vIHuNCOxW08uQKcQZc9hTDnAR9y67huLaMM21avYjpK5JVmlio6OIADUzlNMnvGe
/u+CTMSSAbcBDNBtMarmERFePMK9TuV0URrqNPmJqLrhGGrje0Rt2QVOtOKE+Rzd
QCWirkNkl7qTAU5h+dvaOnLL/7/2lpgQ1bQAR+s+PcB3LpIC/55Pfo/q96K06PBb
IpoCme58AAEQi035e2vTVI4aRO3ZUwgMXcuxu4UXitZDgi3aIr28CY54MYyDB5XT
XmtNMD4b9VvuwNDNaY+W/l0z1yD6YJz8H+zMOUJDuY7GwHzQy4R8CfmWrQUYK9Fh
ThcENlujcrCioQcW84agrDseAK/xykNKi2JdJfi2Hq56ksFEayzQB/zGENsL01Qg
dLlVVKTWEm5gqQyAgIqFufd7V/DvoJvKEDAHKzhtN+oOReD8HSp+6LL6GQ0xbwK9
FR5ljsSBVuffIR7yuXqpQEAYmGngYHRcKsq2d3yYzH+YI4dICvC8PISmDYbsUupY
qVx5JI9WotLNgiOCRgaY9W+fF6fC+N19UnqV1BpAJTuL5kkSslAnVhm1odUVgz/2
JIn9NSi4MDeI05qQ6IJkS648RC6WyxDjXXUvOHkthRNZXjVKT+GRM6jbXeJgKPTc
f8keEKC3ytyrnU50uFY1x7HDUBSpaFrr25z8N2Nl8gQGHST0qXyNHcvqqNSuzx0p
5zhkR5fAzp18LosqQvN2m9I7jhN+pzUChRdE5PXfsFJjTBYIvoQ5Px4S6yKlPojv
8xoExt0C+DlI6OAn8FBRM+ZZsBx0Tb28fSOVrO7f/btsLHgzkE7uoQ/RA0c0WRbz
DdJs/glUZbc2mSiPJt9M9KA+3yr+N3ELNRii+dtPv53ubJIUSATpgWT1+3U5Ivg6
DQeAEQoYSrXKrlFk4mcOt2JD5sgdRHM/2Jxx7ax6bhoIPoqdYaI/23D1yX56tLl/
s+6L0p57niR6Q8LCKw0UnHjmePHbb0h+VikSBN4JHO7L3wrTslfVjnKdFGG7TZ0W
USWm13+01ePpX6vqr4QfqUqYl+78zInX72cpX0VtO/cOIlRV18BWqwUhIPIQdJgE
B1tD3idkMfC74W4aJCvIMofkJU9euQGQ37gKtdZGGa6B0r4AGggdoo/OCP4wgt4S
+NPei30i/V2lCiwWFtxOFzR5dmGg6Y8XXj07vin63/AOIS5hjFuQaBaJ4fRMfM6x
GSjwwGB7Fzcb/MftKSYApsKqsP/J7hPSPYlop8C2vTaLnjEQLZuPCEHml4g2F5p4
hsX11avLEf0b43F779Ujbf4LN5dJrVvdLPlNJQW7+b7UoPH4uvriEvye6THtnYki
Iby+KuLlwmD5JZL7J7x3nzndIN6hGJtA8jiundtjsa/YjDUmCRanQF1Fdyvol/3l
XXG4eaSVPqZ5cdk4dEOUsTje4TgEhYpYS4Vod7yq/b6mWIfx7xRDhlQCcs3nRaTF
v3ioBmT8d3QnoUj4c/wo2Bn/GvVQQdmp8DIcMZoSgxHRYuJBUlEkEPnyPSc6UevA
hc1zjuS3dwyygGX9iaRsms1zB6wFbPGa/asMyR9igc9LZD3daEUZm4oQAJd+F/5/
mmEwKTLDSukztCkaPK93SA8s50cNGFTaY2m67Am9N00GMCX0U1Z59kiqjJWgJeDv
YBvvKOpFUJRq0N7TCsGmrBJTRYEczxfNthY9dsSheh+R0b59Sf0u9pSvhIYyhsy1
WKmshLRmCzvJTiTkwrHLa9V4U9ARpAm/E2l83Jcd786EpKCkEFp55EfFqW1BLl8C
Luv01vwSydnOguEzz/cWOe6RKBZ4AWO1RXvn/yQEDb9xusnLnNCOu0yeXHdpC7Ho
DfxBv1ybXxotfsDO53OGqNMhdsoTfJ9cWzgjgZY9ZoLG1y/u94S0+joY/K7VrXgY
pOgTRpGL2+nk23yCsLTwj3lrYX0238VgSiXO7B9vZ0QGExjSmekZZmpyAlGtlkNx
yP/uc/7n2YTb7K6owxw51wNI0HROPxtdClowoHx9B7zZxxf5+uQ1bM2O5ytzK9Z6
3sMv/Q/KECgNaM52IcwSDYLzE5qVl+6XTQtKEDY19/+6AKgBen8SV/bX9g/ytOxC
jcjzLDft3lJgEwiOEN6/DMph6K+8RUhjOlmqCZzWI7qq5/JQ8HPBB9JnI2U21SKI
65h3kRLScBI2QGldkjQ5vvEhFMqXB8ww2XTu3rRAjujaIPzK5O31Yi30O+9QOrl5
am0jEKBm9WwItxdCMLd88dcCgjYts8uSEAJIoUw80R6MgsXEZLaooJUuGm3rLu9z
gAIYsLMWCxpi9ge+AIhxPlqtz0ZxZChixPNbLgfcpo7GpujJ8n5kD79FJXDnBvsh
B/v27N69TgFEviDtgRHcoPf0JNqTBNg9zo/kXjsrC1LSqL7PUogTW5e3zhFNnPJg
kpJ2XjIKYVYWJNa2japbv+cRcU2HGYPuU1voUw0ekYMKW7JvYCjmh5H4aGELrqav
qXfDK/ijCNe/fSRQC0PDXv5bhq583iMUWbAQk/UYbkfZN7f+Y6MjLBkoIvgW+CLK
qpdkim1dkYOkIpJgidWdSGtp5HBSgDroijewLA1nWIt1ZKNcY/wI6fac2LLgYnZu
mCt/PEU6i9SVsLnfvHqfkTw9QcM6MapJ7UvV0h1pyRNBFiE33MHuFib+PC+zFkzf
r8+01f1nFiBng1jOjtC5GBsZH2jlRXIeEv+hAShYE67U8K2B9AofUaVRUxEZUMLM
I08aM35+HjMZToG9NTqvZFLD1P5ACuFgSKGSDsjTDQKxecEMRkXfT5nU9gyim7qS
LhctnvoKZXj9KWOXLmyVo7wGzG3BnaiA+vzKHXZR8l48wtuRVvv62RxU5pKf4htq
ztl/62JBQjhR/0SaMd5H7bQ93WzViihvLVZgRHCBB3w4TBXqjuIyUG57w7tWztji
OUVz9Up+QwRFctT8Z/lLd6jRxmMb9uDZB4DmJyFJWUotnyYm21zOJex9VsrHV7CH
A+mMcatxrHp+qpP47pxMF2/4+sERo6++xFB9z8FEy4sOT3GVw8/ulkkn8o1KYNAx
FRubIGEyL3UX24WTFIFWj/nlCYRirEc5cu7M40Ap7UmwZyO5x2yxxZactegZK3KH
mBnhdviYNeK1UfRsMnkSIQ6ZPFIHNRaOqrpmkKV1bUnXZ4+hBYkcXbj7hn/iGVbu
4X9lQOENMI/XzJkFC/5N5b7mzYE/jdXbkE+yqBTzwwqHV544PlcddA3X6mvPXLM+
QJStMIf2bt5m2i7rslBPeSpU8TdZpyd0SqNO7v583UGELzyT8S+mYcMjsaf3BZNE
TlWLvp15SKVJFRyLCxBjsbSu2h2XElY8PH976Dg12xNCB+gECl7lo4hAZGbhHU1F
Lsmpf2naX2nmK1xqXrAkzVGxoo8ZlEEIMMSWGnY6N+MKgqNx8lCTWUt7kAe9Hpeb
MXq2YB7hLmJ3pR5qfu4QXtpTx7HD5ymi4OIrzyD42V7R77TYjQXb3RCaywx7DIBJ
1qv2qFvPD4jcdDkujmLfKNFU5rzM2DydTrZYmpieTo6MYiJ4jX/6fdLnQ6y+bsnW
t9t5B6SlnM8ZFNKDrSuSQleGLEGhYHnIMdqPsAJ5ZsQKyTEetR/W2hyh7QCX6V1Y
+eWvMKAT4b7RNfexbb9EWEJ9CfPyYt5qlUkvrlkMhrpKraUDFYdKu+CnJ8r0o2w8
P+nGt48UgzWimZAcEZdzHZPpnOn5QP9mvHLW5r1mK9MFVRJ6nBQOF9FM0RKrVLwM
eGP5ecD+hf7rtwXhavKw/i9oVy3IWc26wpXLEKx0O7GTmptIaKBEygcBkVDPVlvd
0sBOMCxDy7t9AfH2dgt5O63j3AvnQrkAV8ppxaXR54qK3M9rQckBpApIkHzGvYLe
0k7bDk10D9tl0KxIF77VbWjvuMuCSk4zesyGRNxS30GO5cZMKpp+EOmJqglU6nKP
KO2rMrSq8J2GWOxMPwhkcyhVxTYeMwoyqKLHDmQXpJebWtcmArz/0FXKp5RHiAG0
ToUPSurN6kuoLW/X5vmXUMjWabeGi//Vn3RYAF4SMWF1jRGyR1QK27XguovFVZ/X
d2IkvLB6ezFJ2/oXWHeC21f5oahkJMJSrMnN1WtlRf86+npXP0qYqKZV0U0YTlbe
wHCbDIecq4Wsa3EnwHep6eT1Lfgb7gJjM7S8mVOvqlnn6cVNBujx6eOv/tObgb5i
YYQNulJG9pi68dSx4CUqQjpcA7GTkLTgdakrZicpbNKjHA48djms5vIOQLE+hKlS
qM1IoNDrt/udQJjP7Uj3P0ugCUIZjmMr0cAopbwAb2SnlFBVzYHOaZ55rztMvDU7
x7aTXAj7HIOVS0QYYZgAtMReX3vG5/lVZ5e4rv2evkN3sB80yeqf0NFktcI33it5
ZqWPY4udAO4dG0akuXQDj/eUvY+WLl5j+1WyPN2WKHJ0kpIsvsYeGjtGycEWh4Bb
hlx2zlNA2U82bBgWOwOeRc4P3EI50Za03u0cSjGhWgDsUFKJGB7cv2tYJ2KSRySK
IILxiReSm/S4ZDFgP+SMh3jgPGWXIywjnOuARBae3I4uAn7ScDJ4O0YSG1QbLa8O
EYa+86r5odxSTS6Q4rJWaDKj6g10YWfVlezQ1kappIfZE9anU8/7KHc73TUAU0tO
HIVemBl5jdcBIJPrGA+KO1r31XngpVidH/Aj3SoMFkePTj/TOkn59/m8G8mgmysq
bZSe7MtfmDEfzRNvDBrQA2AgaNsS0CGD7DqOaIzLSLvoWx5fPuce3PQ6t6x4ThBm
XfixO6pGgSuiTJXjAA9yN0WFCsDPmuLh6qLvqAybk5vrmvKnsW7QjmuPJAXFMZ1Z
HBWOGVG4lOvXIq+bv2+NaKbXu945X2Y43gIMy98zB7/OeJwoIVGi9MNgEC5BRTr/
yclXjPuriHwGEDBKX679FY7tWxGoQZbIrvsAdpEEEIZhy1A5NPdbjyojJWVrSnGh
shO/WH96Cf1Sy8z2g/uHV++5TstoXnDxH1DSCGNDTmfwpUYS5GZ5ADMiAMQaiQ6s
MtIg28fBdxhbQZKjmpKm5Ls4FBQinDY+JTFbGN2UocAcrGsrZYOZk8Rp0CEnai+A
kIQlHYhYNundgRawpmaXixynXKR8UVPc1XyM8/zx1hCJA4zc6E1RF4KVie1kjGnN
Zgosg989TsiWIqYDRqhtYhkTdp5idE+zOGNuy0HIGnKuzujnJYywNvk8AkGMfjbS
S7/heVWVI2Gdjk9h+9WLkqmH2m0ahBL5wDcP213bs2Kf47ZlgqbzeMZvAQoPbTUK
pOLPEVk8DrTgQwEKjZTsmPrpnfW+oMFEV7hOzA81XJSRZlFDEk82lz3eoJLXF1wl
qK+Z7uuKOwyKmJmhYi0IfsC/XE6hGnw1CiGYwp022XyexDoI7VQaBPZ07NhGUCOJ
zhU8adhTKs7lW2Xfp9mcBCWhWN8y2UMQoGk1fBAmxDzpF8+veMbhd5sTM/GBvBWM
KRGHlCKwZjY+zdpmHe+WCJe3vEVCYASPNBa9AkJsvzdQQOAjsFR+ALlsUMMhMq58
G+XsEHEBFHMnPc9CgjYd+JvaPaydvXhD15xqZLXPXd0Ix0gZ4h/WJJ+nhADMIH2y
SVnbNLtobOsEvJ2dE2EDCHeI5AgU1fo03rQ0q2+ffRHur/qtR/ZUGSyU/7fepUwG
UjVp4SiqtqcdahuLLZmbGG//pjeNrVS+FJ0FWsJYHB8n58e4DyK0nGKerlqTiUUK
f3gCk2l0FJAM7OrX6bfvOV0ERwrYfAkacp+WHxi7F0JT0LyGW6nui7DMYh2HngRk
SxUEOcbgmIHBU7Qpa1hJJ3kWu6nt+N+nIb5O+1IYexeqLTMF6zRX/irQt5f/lRrp
qfexVHEgdCZcRm4uyS5YSxEGds4kt/lXQdtrHSwqjvbKKyK1AyXzBnnMcd73jDeg
QCoBcEByWJ91fWmuHrS2XV2zPwtbs8LYgeupbWlKV88iAOzBoo3b39tllhSrLJZG
pjSp71WVaaJutmXqt1rI7K08xQW7NE40he4+fVBy/NnMX1LFYQDndTb863KmGlid
6K0wVBF5F46XQtkBqoz8VVMiANprsQE8h8H/cSGi2OuBU0Bj0TiPmOUhlI2VlT7U
Jw6h2jQjopxNpztjaVVGjW6YBqTJQXwSWhDkt/g3zfntYg3R2ipO25MQPZNQ/f9A
P/LpY9CnPGM8qNRsxW09fCmxQzwnOKlCGw7FxWxDpaj7mLUxw9mVkNNkvdMMuvVB
WlP5NB6EpdlzWqSdrp2nM3kIpC7zfx0oPm+FV7XWINWsl0KktwTzjtnXtJCiiHwN
CPGAAMYyWptIgHbFosJ1PW7RJKGRyNrSCrV94ZSZZOdCrMoQUFD0fVx8WCUB6iOm
lOWyd/gkVlUzFmzFJ3zg+1JSAlTGDs57Ma3tmJSMRfW2g+zbscXO7QGxpE4G4438
+YCy5M5iooKHqcohHBNJ+48XueII+ADh9XwA+sX8qqeAmpnEh/Uyet4KfWtkrS0E
i3DmJBf4FWv5zqghmP1E9VCtBhOvN/Q8z73Imj+Ik0F06jgeNlfffKZ+O2prwx1f
UVXmCeM3sIbUpylnthOAwZ+qcYSZpn1es+tGZSFDgdc2QrW6rJbtygnm+B3KRzlN
gKz7m+dntEeePHAVIWLlHmgouisBE47NWQN+xPRAgb9mmb5T44oOY1RU8dF8iGX7
ZqsYVNBwPOSPOikAD4DfXKVHgBTh8alrcK8uQRZImK+v8r1agEbJZlaNKIat4lHu
tibIMlB+x6//NP7SWLZ+rDgr5v444iZa3hVKVSkNXb/HiwwKyBHdkkijtG3DdTNp
MTSea13bLkgyWRJqY3dAp5r73rn10JwHIKkXrVkTKx0vYq5MOiADzlReE62NckxV
VF7y7ybf1gOPFvGfF6rgutIeQ6PL5HT08nBbj4yYIkPhSQUEq+a9zP5eC76C4BR3
cPMr3Njbya5eJ+soQ3Dh9ubtRrGautb+mdzKASGEBIrbh6fFMYZIjV0psvGskRHs
uZJng0fUpchiAulKf64Dp7/oUTpZWJroXsIDtf1hPXrh/4J42Fc9poZkgO/DoJqK
b6Vekf+M6AMnbv81c2N/wUztGe4gRf5qFBVPCnJ3JB7y9D3vekChEmzYkjdNjwwr
U8vNydcHQIJjBV+i1spGFpXZsk9KNGIYT2Dab9iUlUp/xh1Sf0iD2ypn6wpZ9JUp
MDmYCyh5zUWMIx2iNkeIGKxSI1vQIQeiwLFoVg3icAqJiaYT2RVAcV/q9qaBWULA
dGdSWj+Co11elPiGhBxOAkZnEFVJj56rTzCekaoXseR3OMV1DDRXhKeyx2L/QyAY
xppebAljL7sVyS5T08NBZek1UAdtaU2b+jBPmR6yEOnThKMkIsgw+/Ad1Nde3EGZ
5B8GS7ANJ80IS4yBeup/ralzxNQt8+0ChApazmKLMeUIjGqd8HdBcQVVlEYJdRPh
FM/o3VOumMDkQrXJYzdKM372ou/1gt4VQHx9UoycHh2zJmwri4SQp2Wuvf9c0c4M
h/fpNlWNPrzklwcSmJRb2cpPMl/zUqnI9lHDYRAMexPg6AfiueuoJKWBjvcti88U
f4sbJ2FFW+0eICfAlUZpUaoB2/p+0AtiZQjHp5XANfUp3oELgvyQXlO8ZqheF9Im
Zm+LoHZNyVup/upBWQRn8eyzdEg1weY8Sk8tpaHYWhHemZYTwz7zZeuqJEtrQNqD
GEkRAJC5CYYf6C5AQnM6Gh9+b5e1I6TIzy5AAdcKSmSIRcgYi6N9acHtpbJ5Co6e
TpKkKos/B+KkIegXQHzPjFkgCTle4VKI0SDofqPEH8y1iMqAzE9QFQEG5bfiDrEM
YW6NCgnzYAYRpJQithGvCsk7wqQYcRGXRyigjBuPj+Qq2t/IODtdYx3KUXh21tRr
fAwGa5Jkp1lIhO1+odW+EJ0piBsItV4cW12MiiH9OlTVwIO/qyTGubLtU1rnBIW+
ObqZLF7o8aTFmaYDeVha/ShqW733ih7cYdBOK/dnrl6rXaWA3jytdqZ0VUeGE72Z
6c2VNI7xT0/X6nPnThm2Kl7+KOpebxgrTMeIeD+fGNbkp8dYM7tSF2P6HvDj80Pj
kRpW+ikVZYG/aDQ+fendwA+NtTI+UTtLordOXIyq+Zwqwla8TYvS+bAxdwVHZsio
qJnqrtPhfU+fLHkmp8WCVTvGMCUwg2cRV0sskz/B6mLrm28uLRSPM01Jv3tSY+fY
UZ5yUMj0wOud1DuDN5ZQ1enfBvrIONaIe8TFfK90ejYywJAUli5W5NhRqNiGpYXP
UQlbpFNXokJfmXxQfS/2otdF/jxig2IhGHy6/zYTZ7MczPYrZ7EUNuFtQj29rnJB
mBfmoAEjju/601WcOEFPlL9xmIUya1UYbfKvUTELbcHHFpzO/MoM/ySuvSetNxF3
aDPQvWnkVnAynn/Uhy8cesmYFJd3C19FZqZ2CBNMpPbD9bA/CtR2QMlwklYX9nn6
5/kU/czwC7pxIM11J03cE1nMtcRJl2q8iapyoSCvkb7xi110/hDauqwgfqyV8s/d
OT1j6QRWki3+/Bizllpnw1UCmZk918BNpLzpG3iHbQVxGgjBgREwwv9rJfIlXaKI
E8zqQmupfUKSkEeS/4bUoN7rSVUCWPkXkIrmafZjMW1XmnR/J0y6Uh4zaumEKjZr
sFI57lQqiSeLWpX8v8uZQ/tn0Ic7GmeyW3D+aCEUV8OKPhCA4kO13mapOLV5oQzp
OsAB2jI49L/piU1YYzYXauKAtdOBB2C3H2/eZq+MjHtQ7CahJNBZ9lhcDDKrpx0J
J/6mH/OvcGj0w0lL9TeXmPBhIljhDKMNYM6kibfQkZKLPopUxc+3EQmLfvfoA6tF
PIKGyDKbYC4RXQJhOxfDQzPJ80UezWjpdLj4O8QJ6f3qMRVmeCzlRa+Hkm0aeyO3
ZMkXbj6Ql4bAZl+YyCcw2GblF/Frl/CRjkCXi34gNMmvlWE8mXKN2jl7X9FeK4es
CnHlqEHKthjVnI8Tbb3IZvnwvH6GQeOO17fEbcvj97aDEwFQhT8hcwPyus/1aY0Q
uhrWBdseMeBKzYAwEANnVKRKhyHHFjAkrHs6dVqjkRsMd0E208FmiYrH8FFtJ5OT
C3aiIujdj10eiuBF4xYCZnOhWMczyl94v0gsBYK9hc5bnHWKoEyg0ojDiXvZXTZn
HEpJoZptoWB7hhQK5FOKKJHKCxDqZzDe8UA8gtdNoZsuQYQfDmDSUCMjTJH9AP0g
FAvuquz3YI1zQ5Ii78WdDt1BpK2Bf3hmNySn1GfOAX0tTzFV+jJWDZ615ZSZe8jM
kQepLmoL/8KMdJ+8sWunBv7ju7PQ5TcazcCV2buM6ok6RPFzBAq9f0ujLpwH2eMG
PFK/KCtxqZo70BnFmPYjAQEJLFZ6HZmtiKpPNo0MIdGpvsY9ofcMrApycQGd+2w+
hrv2wySVQxl9pA2LJog6oDOJTkgcUi7PZ8dwJYwAVHkpd59+oGxkacfSKL3P4GDk
X1Xq84yCjkPCL6tTRDfnzTAmjeljICSFEThcZEP8pgYZDS8CIz2sdBMbjaEFPnm3
pUvGq6Jfzc45g15zwkLZi7kkjjRSjQUVircGX/xzwoPheT2GfvjhjxsX1/QSE30e
FOrwwdOvfueQLC5BjCDLY1dCPMReU/2RjA+jzQXEyW2BEAyHqwHwGPuU7rweMho6
kQpUmcdLjc6gv7Mj1Ic5zwIjNurhdK3f7Hg93sifmvwGS2Nn5wWxMI/Y+3LtCU7C
VjM4NDKB14lZl791zVYpo5qaazi+GYc8MBENsSuRP6o6lS5VwwcQ39xp/bc6XM3q
mVkZx5XPZCjD4B4CkAEU2JdatMG7McFFP3lqhQjBm0cVoaraYAl4tZU5psYzKiti
6jJYksH1aljMDshJDwM7drOE+wlJP5kTk9S0lnLcq8dHIiUzspRZA72hLayhznQ5
YZVePlAb8I+aB2yY3JfHo8zYdr3GgJYkMkeGerfFQuOlUlIMP9ZVn1LWID1/aEkh
pe7sRby6C6XzylLTPSVtUxuES2CDH2JSmWtJZt6HOS3Zv2pSy7Lk/i0Nas6pZzJO
OX7M3poKsXR488QfdbJFj7kjUZpREF9LbhaDD/gEaqYxpqZqmfpA8tpmr/Izzegw
UxZ5gIel1z3ieTIZldOeBbUHClYZ451M9k6W+D/p625tDfOg8U7BRoPK/oVc4tG2
a2sAQ0TWeHhZmK/nFlHaFngMfR7ONlkcFcmeS/VTnKPu/fCqXx5AQZ4bq3Nv3Aeb
QAWE5KnNp1SVIAJXV7S8aOfGzaUuFABJKbx6uzFcZklZYIFlBDeFGc8gbfYtB9r8
gMvSjtsGf+DhVU5Jb81a/9y6pZCwLMjpFsvT5VB9jDfrJKOwmKvlBjj4YQ2oct5A
Vp2AIWvNindYBbi9wpD+nqgG7BFezze81HTxcZZKuBqf5cP7EolxMvduFE3oUTwF
Y+uQLIQQt8AkmB9oSbX9yiIcgLqqyjyNFre+VcoX8DjtgvANjrRM22n46QC89V37
bJYlhEZuklJu9BaiPa+NhWslsPVoVG2jtihgla+hjr4tZfLs1u/xL9OQQbug7s3O
tOq8smHx+i2k0y5wDVJyXlfko/mQAwCW9l/M+UAaGeR1qcwtkvgZehmM014/fYNK
ehXPFiLcgwfJkclpE2AwnV9xevvTp9n1aB3dTHPx0yMC/GMMwTI4pE+IOrlavlac
GpCbukcbXcSxP1Vwr4V5wODCKcE5FRP15KijAsVzEL3R09YzHPUFpt2BvGz4e+2g
oCFXJHZ2+NViymD65p14w628Vg5chIbtk1q6ruRTJ6RGZGHk0hDOVF9dJkf8qj8G
FiG1pzpw9G7i8JF7VZhXQutWJ/pJYMFkKjPPLTSYznaK82EtnILhxi0Wzio50GlU
WjA/Vb4hRKhry+VFhc7nIILW0ws61ezxI+rwpBibnimOLQKgZmpnCfKdFFab5Nyf
VOJzXm0XwDOh+vWKsRtthuTiPDiVbrM31Mgdm2xohBuxcx2mSQAfS0SlBHz80Zw3
Tkl/uwclzqJwqncAVzqa6OBE62mfcgs+Ch9Udi3fT03zFcEBHvp7iYW9R59236bS
LS2gNeCj97LxaWwWDdKPURVc40eicMBly542to66Cth6otYjeqJBOEJJxT/RBTbw
yo1fv/CRO91bauMeri5mdQ1wAAQu1EYDUpZnUyfGpGiQfqjLyD2VW5cspfbQffNr
YcdOg+tNkdNQvs36WZLbiMZC62wMTvgXe5q4dYn/mcZvLklHPnCF0sPrnb8VNpzj
qobEYZjeo/NFniFCxMoED7ve94UF/GFICCGLF1cxVUnG7L+UUAVFIo/A1OP8twiN
mWaBQejC6nA4kZsHnnswxbmqUqen8HBo97X1nfTWG1eIgxx1zqsNnwz7X/6qjZiE
JYg9UbzgKvaGt0wC4Di1rMWmvXTAB1vkVTW6Mvqk+dXynvt8MOEdROfFbfLU7g+9
I1E7u1+oXoHdxWkH94R4gQBr6tFegtLDHlrWTnt/rTLZM57CQ0rbrbbjHAg1zQr3
fu5cdEYlPu/vJicXITY8zV//yJaNXYQR34stJfpOmOl+FHznYfHB/z+CTlYmugoY
rZhntJfibgjt4SJhedJsGOM8bNwT320iebtOEyr2DMxi8a3d1TXN9d2eVr3zXzlw
uDLi2G1mVQxsN16+AuyE87ghjzZ+CDthBh+CmjwONcWFkHTkFoOUlaOExBx/vf89
PQ6d3AsfViLxxsoTa73O+D5HtUKWUOJ3c6g/v2zxkooz+HCx4x38w9eF382sKUMz
tgjNfaUO5iE0SI84WUHc08IT5ZK5UfcQAu8jGlAgb/8T+4LFmOLzof8CpWjwFMQU
zyJEHMCpxLDcW56LAaeG5yWPjHSe3pCOw2TOQvrcHZ4eG6e1RB19fG7TH2jquKV9
WmPm7HOP/9i3Oa6JvRz4s70zBXIlleWtV1Drxy809tpYUKGVGI6sUlXKf8+yi5az
4HDgIo1vZai8j8j3QnuCtN8sxgLX11eJ8NypDqPESC3GTUGus4O/kZmpkTVziLji
al4G9QyfuPNayoS9xL2V6IQQ9mplZQbWEbYwzBTk7pxj2JLwydwb0S1spkDKoJBj
gpm9SBQnF02VxT4i5hzPnW4p1PUXfQneY17n1P/1rFARgzxB0MOX4QYYVmq5wbBD
DGEGthtrTO4fb5SZXqDf4jRa8NJp4XU5SPPj8F2XVlRmZAPjoczEwZ3w4xp5GnSM
TLLCJt0QsoqXzJ2VPBVr6NdO9RA5p0YSfFgkN0V9cTUqGDdkTh+EfMxrZpXTGcXs
zDmMjxt22kIOUHJ3bSmiFk+dq8TqQerfUY/8KrHogXVQ35VaFabM0gwcX0iCLJuS
OrjZ0ToF9gR+4RQ43kGwn3Dk0iQUilUNMKofMPMiKBSg+CIAVe36+OCkRev8W6kU
sn13rrt1xs7WDuJ6+EZo8b4boTKtckB9e+y9fbDo/rBOQTNWBf8eDkLG54uS94t0
DUdtN2JgY1/s85V9uvCj8qhAwCcRrhZr1YiU3vG5+gZNUWjeGsQSbE2E+7Sr5IZ8
6IWeNUKnKaMJD9edhRJUuULlptNw+3W4FsFp3t+2VBdyb2H96zz8xnCYHeTAjry9
dncHa0zd7L0b7hMSiVh7a26lH2vBOk3urbzb7IhcQiztTCf1lhx5A0COlaRqf86X
olbE4HO5TAtHx1I/BcBXIHa5pUz1Ol8Unu4CnZFOON9qzzD9mXvCzMQ/nyyAZVDw
/nq58P19M+vVa5jlJLUOFJOG7O69bI9DbRmEdYnsehz4eRpSmQdp/rb0H3Mmhqtl
k0TKcDzj9wpLAKbR7KLmaFr5fRaMkci8sPqCIxoLySBss0nsxNjbDytBj9QVfFg0
1waAAtUUGMAfCGIuhpsIpsW8DjH7d3/xhY5hmJINrJKNLwnB5bWwqRQrVx/Ehq89
U5CizQL7/lJhgDoQOifY3LB+qBpW7hfKX44y1utlU9G6t1VJ5SqjR9fn/QWtSzRK
oeuYbuCFb9zct9zHEp8IMDlr9VtK+eRQQLmKq0fcxgKPyV9hHxs35ga5cWfIYHWq
g0vFJcEED1fKHKGIPbHrN52UxKdh2HauiIUYt4/r+C78rVEayg+REo/locN3Ed+K
rMCU+xwRBsRjVTRLJpUbLiZyZ6j3b1qMgFhrhFQmteJ1nWOyd1DYB22PVBfW+B0F
Duc8c36OaDD3gABhqbkrMvN9l0+1rqLgnPMeWrCeFF8bmRvjWkYuP2/GEZ706BMJ
wrJOavTRfTnR1p5Bq7K9TxJRae2Ehhw26gfiqHJ+z9emPpahi91DPUpenfGfl5n6
xd3BGZ2+d73eGG6U6A/3FlUdjczaOTFapnCKoXU8S95kGw/93j/uaNFVFBK0T9u+
cwBRAUHUfli4M7F2r1/5Wmsyfi0GVa0YKxXkagPtvY/oRfqlOSxfJfPK5x8T0LPV
sJN+FbszL2H1LQnpOMqbdsQcVP0KOQc8WIJPPuPLponJNFtDV8jaGzNiIbS+mXc6
iiMWB4xfm7W7BsvMjsAB/c9puOWEvG9RNJ/Zkw1p8Zx+9DWvcZnJMVAk0/ROR6Ud
4aDjHG3Iafw/R9Pth6LchvvzINqejfsohSTCIMOO3MUhCkAy4MuWel9lTrkX//WM
RJQcbiWqtdghCVpsOP1m3qv8E8ZD4hyD+OOkRdVNdGaQpgzkktieAjRTuY3B4QBF
fGI0FSX85y1ZpiYzADN91YvVmUfY1yoUpCuo2HLquz9XGOtLK8BJKzZdrrG0C8qr
NWcjQ6/NKNhwl32WE/VPRUg9xPC2mwYTZneZUicVoSEDaZDy97hIP752zFpkf7cE
GX9aUzCPo+ES8dR1Z2kkwPBifhsRanuyNP96Rjjh0UhBqVJFloglP7UtVtga96gk
THhQCJ36pJPfKxkXdkWc0L5FV6EAMXQvmk1nAEbQwe78mAkQKSZmGdIgL8F4LDaH
NnpdikAHyGJyvIfIg5WJYBFAlEvtiBSjvn9uXIek4Bo8q3Zaf7C9rKi3UhVVzpSC
K4q80bicB7qawEfNg8dsHaNs8vL0q1OIqIaGwdZ/bhI70i1AqmnQJ2QXXh++NJ6e
nwS6bOfgcYo9Bz4eCKLCUwkyevjSQenvrGUS1rHSxqgDkNR01VjSypWdLUQIJ/gy
yYTaQjZ+7v6evz3fVf4qe40SkW1jF3LwWPc1jHq5IiMDbOZ8kgSC6Q8PH9HhyIyM
PodQf5VGUtuc0v47EFxoOBn0k11PjZT+pa5Tt1kyQxHfG+uvYX0E3oT+HZzixNBo
1Tlq+4HM1U1D1JVx0CCIw4d2fpRohz3OcPkJGA1JGRzEPccpLqSgJvAIG53qqEi0
jNfXafZ2+PbMEOtzUVbmhEk41KqXMogy4WAScsSLO4pX0SxX4a3NxVlF9Wpw1c5u
cTV6G4rsB1O53GKMTON2nwhLZIaa5xmW0PcEJw6lFTnJcpRnDCQeUvL3vM6J55LV
LqFUMpscxuOJB0x7tVDPPMPyL+RrxtotietDjqz8gplkAffm16dxvU905Tf4L6lK
h8C1pxjXBzDeUtU8a0iEmdNY8iUXc33PMTULqlm/mUD2s508gTdJisHbiWjVlf4I
lrv+WU5cFJFpvrDnplWJ9dC7QBQdv7wWEgVgC9tvA1dACML3QLeTahoZv/aDVLbi
YRwxQX6KWwlNDluFEFvXo206oVLrFBF5K/7sq6L9Yv5CMPFN0Kmh1RqvcG59ZM0S
MBEnNhjlsAO8l55arrK8fHu4mD7HGqRombpCr+q1fZnVFSMcKR13oHUI60DAtjVp
gAANwa3yYMbZfEj4kpaz04C5sfKc7cF8S0Y11PVvxfrM5qv/9uRNZBJeTni8kW42
k2DpG5CRUaWrrhEdh2QLog51b4Q69V/nx7hSmymgsFuhXfNsgyEZQ3HoZwrNuRVq
NA0c6XXiDOZkIsKzb7sat05LwuoR5F/A2RO/AxQXc5ZJ5ACx/FAfKucNf3z2iE+4
nKCFdpqT7/qVxo6PoiibIVtO6Zmul4mB+Q+7sbZHmCdwcN00G7m4qUHZznPQzO4i
QSpJ1bVcT1Wc29lEfSGBoVwmbZEhTRtAIDMJJtbQkipP0UvtnGTwXtIAZrgwYAou
L+876/FqAaPcA3GMddp9LZP17CGQaiZxAfsntGEANxDyuKIeED2Edwr+EVM/fC7m
pkMTAdiBeeur/k489Dr1Gp8diq9FgQEQGdxvKNOof75SGMYAggIu9QaUH0BVY1VR
z52NugcLGaAbbEqnO7n0yHy9KNzcDqS+7t0pe529PNR/i+8prADTJMr2fvD9Jk7W
/M5yIQTO7BfM7xdLLxcyvS3ziJolI4ANP18+vcJ0BbwiRdntmPPq6wWAMhIH4tGB
gn3PErEhTDd88egF64z1172jq6/T10FGt2M5+m75ViogrTIcbtbg0HNRLbiQ89Q3
9mpAjrN4+7qWcCNdIWNQTfZvDNgFXmxg3sdIO8o6tpDtE6YAH77tdgBXH9si+vYD
/Q38k44EGKuXiIsWl/ssod9DdBeqyNh54YGzwMb6zKZPUvwN1/ocPEpgtc4p5yyN
O4Tos/+rLywnD18oukzXiec2jhAiYcljGY2PyXjgC7RD2nroBNMEuqAUgq4aSHdT
ktVNB61z+xuJYXW96fst8kKYhEqlFrgPTOs95eqZDvf/81TyWugLoFRkVMrBXwSe
OHjwh5JWeHthuFcquh75I1SGDpqonMrYuhWzen9CM34iDn6qWKsFaP6SrmHlVGqp
y6NIRNXSzWcav4w5K3c0RD5Ol/F0kg+swmAF2fSW7nhghiJprON14QWwbGpaMTWj
Eh8bTSY3tzUuVZH1LcD4676A3kK7gR2QQqn3tEULyX14vEsMuxu0xDCoCojPynWk
Etmrr4okJd1D2JTe9WzK5pA6hIGjZ4HrstcbfJu0l+XK+G1axpTUmIc5ZIVjOB8m
G0IINaTcq1IeM1eIm5bXjx4d2IprE/M5Meq+Ki8pFjDixoVKW8+pTZvgtctgJ3mN
xQMS7FLcH920E5M/mtyD62/sQXQSs9yDEF2uLXyjFKPJKgMN/L+cc5q6EsvExD2r
B8PoS9H2jdzXMogPW1LTUO54/pbv3clJ3C6YK09Q5C7G5LelV8Tts+M2hh8zzIyp
pU0mXX+7xTj8D766QDaS0jFGvwFSSs0OCoR+K9XeFiT8YNNqu+T+/Jj8YF/Q9Yce
W+sPJpamoCX2MxLHNaHsIHf+KSd+Tga8zOrnCM9ZnpYoBEhCC1mD6I3zh0hNAlpj
sflHNgak4JV4XzWY5iAkGDoyncCjHfBnoj1b8Cl6KUOHiQwHPZ9DxVvInKCHPu+6
7NFZRJJ5YStPg3MnLvuP3n4BiQgFQb+s1IZ9OUoMOYijpVInwhZna6niIn9OToXz
xGvkSBOJycMiJURFXtLJi0nC9nhC+JDOZfPgYSYcrXNk6fy5c0YcOKE2oprw/pry
mwUsek7ks8nOHTD7sr6YN3JbV9yW+wcdgGPTqOAgkiZ25g+oiGS3xhkIimymXlOA
5PSTY/LO6wJaZebwkBFch/lkf28+VCjosvk6HRGZbBGIEVSJ/fb5Ntaf+pg06gPU
e5DS/fWMD1PQaTH7oVST7iaoXBdj9NKmv398aW59qLYcW5EPEgux12htWpTqS8KY
LSvQxY3owDaawp0WxRVN2RY81GnrPTL6qx5AFNK0nKNHWC2iU9oSAv4AGy37Ay2/
pJ4lW1sQKf95SO+EIBRyI0yJayg/kYy/OR+Pm8ik+i2IvNnfIaiCBadQkL/ltL2E
uFOT8XriqVemkj7+h06Itd+qceagaWMiCNaSC1jiu6Al0myAwLL+sLdVXWNYEZpU
bR7xYqXe3pbpDuYk1dDhgpaGqpAdsLC2vo3aJWPujKHFUHOzne6dYoBRxkmunh4S
7XKzzmwXt5kCf60vR39jgaHiGl444fRKxGU17ZaOdhLyhYCuAW9ZfxQlWWVVfP+I
KG8TXWMLJZ9vdM2AIjtEmDHWySNXuDZnzuRhDUiTJWO4He5DPlkVEKqoRm4SZGHp
tg9j77CB8VoX8/wjZmZ7ifw8Av58tmPmSXMoDKiBpGF1rRZ00fprQ0Fv0Q4RJlaz
7Dm/hTKGSLxc2/ZNZG8/g3XeILyLVHsolgxdB6Kj6jsnV+dDBF4JjnY9mtLZSyBg
vn8HcjZ+Sit0LfB3zwyF4VFISVz37ED3TyyvGTuuAzjLHLoUxdJ3VcgsNewKv/To
8mhDJfSuFvfmxljU8ZOoIr6Rx6H2G9EhVRhTuMMikPRid27xvE+1tSU0zZLeUiXk
DwfKhIUQ1jXrv+z56/Z1ooB1DF7TtML9SFpGr8Y2m4cvZUN7N78giD+EPeLv0/G2
tmmU+RQHW3Q5d4xaKojE9e16yGC1Zau6kv1WGtMyJ2IHYIQBtJRPZtJMpSDnWTly
gSXkb5/EftwmSR6/pCTpfMmJODfyRElJj9lIgfT+IrzmPofnZttJv9tfvidboV2t
qC9Yf63nEGT2Iz6sDonzWkYM3ZCq80PUWcvxWHsY2wuHZaeNg8L/3APNjpHojy3+
ldpASW3XVo0e24FuHQCNMzhxvOrdeypRrNqoa4RcHgwRK142wq1mLb1KQDXqKgVK
blfJCdBTbvWhd3fajG9T12SIZt/BNAN5VO55+/Hl85NQ1sl9xu6bgWBtGf8pZllD
xWkuNB025OCrB1VKShJ+uRFZgXUzXAP1e+vYznsqM+nfCt49jf9yF17c2w2NeKXE
YAHDAOmX515BtOC4lEy0MCnr4/53xXnzvSbR+BR9aVoIky6CIXM+lL5UQhYUDTJv
whQ7RCgmV7OYWvJCwyvW1RN9SiPWuh0Q7pAGr+LgnYTKwjbL3QpOVIl8GYVScV+K
3IyfgwmwrJ9BZyAleiUlDZxt96naIE08oLdlvw61by+upB+uUkj9iP7IhikXDFhq
SMPIVBBxSg2CT4InhaVPmq92YaSH/Yew0cWfxKZIHb29wJFr9rqB2hFAnryqI+t+
JTJlrImV2jgF07kuxDL8dnmbML8NCkODoXrxvcJIs8090X9Z1AFgTpLTNdTrqjcr
cubmEDLszlSjF0em36T1hw0XG3SHOGloAKmAGKxTL/KbWeerScIUqVaUSe+5gc6R
MUJ7q5IcoqEphAD9lHQNunuF6nKgEgVWFeD9fZT4b2Q7ALYxj2k5uiAmsBpdhXje
RBVcoZVwLQdI9i76tJt6XrRWj0AvHlg36RfK5yn9DEzqikUulS19Syl8H3tE6i4w
rwGjadWY7uor4ydARPIr2SK5fGRCdZdYkI7UFBkX6CiMmqx/jrpUnpVDyt46RfeD
JdraN5NB9NR9ZqhJl+f8hhzgzUUuZqq2JBNy9Fsge0qxhIU+sosEwAopEeUfG2rp
irmNIY18zrvElBBux3F0OHko3+W3DD1+u7mSdqkHSQW7hGS1VPj5DMdS3zmezwqi
r3P+MuYk/afgdgbMXPIUaDU7tJ7TpXze2Ypi6wmczqV1oUm3fnfb6ZiCoun96AfH
p1kOghT60rKQFr7ARLs3aE6tqaYV6cnsIvLW1UZ7nI6n3x+a7N1CQakrtj7ENbqC
bHsJpUhoySiFWR4ijGwLHjxEFdQhtLB0c4skZqxNHEEk9Nxr0KODIIiIshqHLjjo
874oFa/bXD10RHGC4zOGQwI1Lir2wGJKXMluMd6Jltkz3ZciOX56fs5q+JNlH9rd
0tNp3bTqu0Br7KnbN5qNjk6WgQLPR1cYY2sV+vUrvvq3i4nXPX6PE28ZFnVp3nl7
yPItSiXjmqYqur+lIR5ZM4ZU26Otqu+jQDDkbCgx82gx0lUY1C5xvzecqJOzwPoe
HSak5bR/BJWB0dKOeiVERCqWH+8x6097ge0eDbx0rQQnfRMWxq4q6dlIiXwPPjyY
a+PaPhAMrY6upDRrw9kMh2tb5AJBpBdJFLG2G83hZihO0PcWrIgnYlotLhTq2Keu
Db0pIaVlPf4BcsDHxqL0mShw/Ct9XEHqXZ/UiyuYLjBo9NVS8h/aAjmmBrIM4bKL
SOTLj0ClqF180gJ98XLtnUeX+ba3D/8GaYJT3FzPPTwjO/w3bOjN1RY4QjCDuOEM
kB5LQ1RZ+9iGSc6RYitQO80MhGa8qSh7qBbPhvT+EHUbVUqQWjnZw+yC9GEbfOdI
tCp/1S3PWateQeWdGVsG9aPtrbmvwptrVpIlSWqUflaV04TUljAXoxc2BEtykZhW
bS+xPu4dz+xExujW7WBNW+Guj7ojRprQvqREvuueCQQpWSOqp2JGXYQz9V4VPJhF
+FZ19RWtQwOvMdlEwRX0Nmwv6pKq5xJfJ1Z7TBi+XBoORej1EeJz7cV6F7K//T0y
Ko6BlXsBeh50KhvrLT/7z8OTGnADwnW2Q1o2eJWduD2ZhLLM447pX3I5zYV28LR9
snB6Zvb12RQdJjej4rzOiyoLF1nDjsU53FGB9baeACN0sK0AVOHZQp9PWMFLt+IC
u1F7vUxxosFSSZ48xZ42K8kc84FXmGT70cOOR1yHFfKUV9qZybWM3J3lMPLEGnWo
0MWZZr3DKjvm4UuDlHtH4mv3K6NNH8E199xSKu5RqjOja84MupsH8d9sDq39Cw9P
F20nsU8NnMqM2cQ9gRFwBvc52I9WkD1jWw3a08Ek+aFbIRdK72/MHXXUUqkrbW56
JIjix4j/7a//YfKC7zUjyowzqqiwmvN1VfGFsBcdfNuQ1Msd+UAdGPjcTzsAcfNN
I7+zBIeOYD6M1sHMwYz9TsDvIjjMLWtLkpdbqWY1FER8wynkCymdcy3RJKrOcpCr
2Dp7Yo2aNw7RchEOgDttZ12groc44GRKahbFaRkg7VjCVblza/QI/uoiz06Zwb40
7KmHMLtmDIjZuE1onivwJnlzflBwmFPei2dALqLhvgUAheKCHYMXpb2SUAdcBGDz
GuEkpAU0BD+uVIJc3GUXNzKe7aH8vwdQGbfaDcCiG/s5Mdal/EArxZLj5wB/nC6h
a/727wAm85NOH8bODZMVTBXBkHPQbjb0DaUwOO37wBYj8XFKcCcqDHwBJSe7PfoT
AwnE1KFxV4mITra6nky7Z1Tb4cn+KEd143gir0ITEHW9y4xAnqN42a19UOlugZpe
B6NZvmL4sLaAirdKf7WUVeUt8ZegZdsUeZHmJBucP3nwkbOXbqk1dbzS7lpZGexc
/gXfNeGTx9zzAROng9USTgzmIivdGvYUaGA1nO1GgwHQwh/TugSo3kJcH1VYV1by
0G08mXXUgM556EZM+Fj4DuRncLs1qdOwkiuxWfEkejypcQF8H/Zc7xw4tZ/t8lrd
UmJmM9cE5sPNJ/fNqmWxsctx+VWgwF0//RoRA0NhfXP7QXPD4git9zEkT6jRFiEE
z3H5bahq7kR/NHDfyxnEY+CBsJMx/s+NO9MZ2ehsZXByOteGFy0J4Yc10pdLVRCj
lYeJFW2IpYOxlueqSFHahEorANq0hKwKmoOlsLrsRgIcdgaMvlWqDckeSWrfnetX
MNF2VKrFmkgTTH5nKVgTBU3jl8u0REmvDJEdWU0H3i+1PwGE8Yd4X9zrkixv4H5+
+a7FQ8odlFgl1hzpcudvl9NP30LIio12PMW8e3eA0K+nzu630vS0iYtBg+p8UNb9
Bhsv46gUhX4joP8ekCOr3LInPf+Pa/I+KuYZvM0FtYzHsNEs7bOyQdPztSaTajvH
DLw3pYIUt2X31G7X9ufMtoQgvLL05vjmMxUG1E71bZZlHw9ZydIUM961hCng3L/l
XeQMUtmqbMR97h5p3SYnyXTJpOSHW/WSixOEmW8V8ob7QrjqOyncRjILIF+1Of8J
Gt1WSp3MmJQTU3ZTIYntd0L2bxwtCaw9666cKD1w6JSaczEyBeWMhodEvL7Tx2bD
ecwv+sx2H3N1WYkgo4FVOJ2F/7C76B5Ynw45g3hiEXOzfLO9gq+AraomItsCdWox
mtBXSxXHO8qNJ2nhKK3DAoUPnkXMdyJ0YcGWo52gAYX+D4QPOneBg3JbYDFSyriB
+K8H9snnxCs+SSvaP8nLeo3xg3W42JUEwhZnEmcezK/vcMST+qTNS8b0SiyG1AID
Gh+BQvSDrMnxUjCgui83O3CoIWQYSUeoPY+GBl1QUBHhL6tfJovv2SmuEASxa3N2
1h46WfK4aaKsQ0cwoPts5a6Qz7wkUmlchbQFSSlUsn5mRZd+Vdi2jU/CmBl4bZpE
8vpvH7Jr4Xv9ycubmqNkbHOa6tQyozlv71K2nC+etpF+jJomGNhr9WQ5Mk1WkW7j
ZG5nZ+W2+IqEaCIzB08hFCVhcjzXY8ZdxKjzfdYqgojOwLdoJd9dkv2MV+8j+zbD
6C7llaxmWJq7C+m4QlGn28LLsCSZY6mORNtCRHRSyiITET/nrtHrijrXMt5d+NqY
3G1Ss7RYw2/RlEsOzrFikFcdD+XcOy+DQXHqT6xI3unRT1dGMXmEwzmojKWHyDZJ
xjwXRaHia5N/c7d1gy9OXhx15jryiqeiItRGFIIlPsMQ3NACfRGzHcr+FFC/vbwf
j/Jl1QlaOZqBkzqFvqewU6MrSJsljUY99xfdZiqP0yrRdM+XUJs9xRGSRBN/D60X
SHynvO7zjdQM21H64iVD4NN7fXcxT6g7MllatJ9JtOP1t2nzwi3mKQD3M4BSAbue
HMD2KYjV/mOWcPRIsN2rPMwefjkMN2l1JcwFNoiLCYIa5IzE4KwiZvnIWc2j3Xx4
+QwK3fkeWje0JR8XGBcP+SQ7L/A/ghSjdR71J41kYMiz9qWTRYE220+WOBG3/aqJ
U93RDFqdmHiIdAefIe/VFML/uQv8KYEaBySug1n9hiotDXAefNc4XwuFyQGnaozP
lkvn1McZt0L8mAR7OyZbcdN+1fTua8yWwUExZAIQKwVCuerGP+leZoGszNAV5eV8
6s4EIRVfxZnVrvzQ6D9Fo1gKxAvUiYs4tKeUjpdWitX50B/pOSaslQxiMkD31hJP
ml/Ivn+ZzH0X3495QqNN9Whb9EKl4FcibIWl9NzNz08qSHu0RRoLENb6O7nNESag
yXlotzmy6dcF4ynwmzJAxoZaTUvWMV1aBjLLY4FdN3KkGVANEv7hPM+HkmNSSzdJ
Dz/500GLuZfvgyUUZKSH6ocdJ1mMH31rfKwFVz5kVrZhx2kM/V52TmrTFxfmD1dJ
HLJm1f6AeK1qB9mkIlFVEZT3qeQuNyf/pY0AmkUm0iRrdHC1dLyMzj4fgX5oHrZX
1O6a2P5bEL7WHyRis5jlVzICeeWbAsZpD0UcrlfSQAHX4LTeNm2e5uTiVBirkTIR
2WJJ16lEOltVTBmzUyD6asf2AYFjgpjrtTT9ccy2Y3rs+ij41JOk5TxUsGvpBZrS
hNwOzb15MqmVkGPF9eln6GhClHdY7HYbuTKqbuSju/8Dr1bI7QncYpMG+F9iVAuu
V7OHeNhzScnrB4GzpyQkUEIAZ1v5seG9Z/AenJ5kurwYeZTnZAiHXN6bsWSzYDER
Uru9WCI+xpsJv6Z51p9vYWh5sm1T+5alhHIBoycqtyu9DuK8Msq/hV7B990oozFK
zodlytKSwctoP3MI24pNLgPkRzHG/2rCNPnqY5GpOdGEIZQLj3VeRwMWvgjYMjwY
75BVJqn+4hQ5OWWFiYqDcYVuk2C/kSRQf0/Mfl1k+ZFjvaxC98ZQxDCWuVMpxgJQ
hmBg9mnRzkYE+06XwOfVsr1FZxz1voY1N87BcyMbO1KfocPNw/i/4kBHB30j4Hr9
1ahNpgoZYiRSdBzPlZitw+smcL7ap182KsKOk6hDOHiD68YeHxV4QK/zpg8zzHqc
XIQarE+R9B2h1di3IYdQcqQzvJ07ji/6qWHmeEdodxW7J2nwlo5g7yeO02pcDJRI
tbI4jkfmTBKArSjJjbYvlJrdidFOoDTGZHUP+P/VRegb4rw9Iccp3PjXc2rh3ITx
ufNXF5Z3XZznxt2r3+FevL6WYYpyNtX0L5yk8wWSL8tsaUIWCHevuNRYwFHEfQ2t
aHPu8Sfu/1F1Yon+UQ1HLKfHNCY8RA+lNt+FlYQqToHqyMnBQ/Gua/RIU4NFX3Nx
UghorYqzfROaxBekEZ244UpAXtCCz3giZOnZs84qaSHFqocHlt0q/CRGY5OCF8zi
30hMWHCopFXEnFjkcAIVp6w2t3dsdLVgrNTrXjUJKV94/2QGw1KxZFOb8ot3Sler
GqOwd+Gb4BVZeUjey7n2gYE+Bk83pC8xvlBh9wL0oHKdfs5d7eRq9sLEQ4ErVQZv
O/s1wOGUv9ebt2dpC1mbYKDcNgHpRyBttBnD2lSI8lB/hGV59BSdGiM+XtfYqRYO
mHNVLgK3GJlEUQVHM1DLKP+wS9ZNqnGxgdFF/gKSRGQhW6jk2LqoTz26Pr8WUpLy
mQEO9Na46dAlo5/+fsH2XPY/QQXj0uYurpxjgX5Ma5WZKamd//dP+ixbTV/fCgz8
Ebu3uD5PehSwBX0l8u4Q6moc9FOEzQxK4VTNpJkAil4P1gcMbh/+sNI4WLrmS5A9
tvuIq8VXV2FP/r2VxVhu8VA7og5QrCAjXTQ29FdxVGb/YBIv6GTyoPQE9OTead+A
z0xSMO1iwtpd9GJVt1eXQkoP31tirSW/vgYM3b2wOLgUngq9igYtx0ur85WnJEtn
FFnRUK8jTMyh98X84bG97gL2C4R9hiHa9TCjeKIa36hm1BTEgdkBKlHfsmcVaHSQ
7TJDU4UBOxv3onWM5D8Qyd9d9tn78WXF+cWchWwfYefECcDdUv6aUz57oErV9+kF
QUG3oV6YcLlv1qzka/QVqvaoRYiWtGpCK57EcorO+U1f3fs14ZHWzZVQ8LTRbB81
YqxiWvUIKEb6Qcap6FKD0mx1AfClb9jYXMFLeVufVLBGOTXo+rfSyhQhSfJWdinZ
ythJlKxE6Zj97eKCuanYv1v6h6Zrjz5KLzbfszJtjCbpnxasVKP5qEVl4dwkCni0
cs5flumppW+iPaNcQO2IKKr3U/QKaTLM4Y9XlMZv15aL783ae1wlCDazfRWyisTM
puV/oeB/HTuc3pegABDgNOfGme2o/2T/yKxL2Phio9uRu5Y8Th5bu7vIuhEbynS+
qGPDxBWhZPmCHSHKlRKXAW1U0CJ+G/xj5Vemrw5ne6hF4l2wZa8tUIFyDfnPyx8c
IL7X9MXBpQZ3K5oHm+lN9FrPRLrESJQJACD7X1OhOB14F6sDxwuIoRIarFQ3hYaz
Nwi97JlGFSDnvconVtEntcd+/aCdTCUIGh8zCqnCz20TSO/h49fpqaCHbxwwVRuC
aSecNRB2YKRtI9kpcL0q8IVbny44qVhLn7fupUDwQeYG6D+ZO5fApVTBn//u0VSS
rEynrNDkTTfIvZet+jyQlfVKQtvltBtMSye6IEVVC0GRtoL06rnv7L9Vp0d4SPcl
hBPdAnPVcqF8FERS0oYcKDmxgQtZtXwiyL27j5Rt1s3yC2sVpB+OnkKp0ft2ydsE
HbFXAwUSUigpktoyX4Lm/S1wQ9WzX0SOdHvVyg969DClEc/mGKd+KKXFZ1UDZBrb
tWJYqWNd3O8pPs2h6Acqpdb0A+zWCW99S3NQNxZNhezLsXhkR90RazZaeh25PnmV
8lCrS+feGkL96yt5dexRAHyf9T4lYn85sgWRFOGcNGM/vrRtHp8hVYwW/SkinHkN
+KY/4yCCzoDF1XAVsoc6ZXO0FFUKMcrhlUNVU3Mizsxh/VueXbNUe+KOuZDkSJHY
SCEUEcgUJENWdszuA0Ed2AHMMv2udGGJ58uVH/hHSWQEJTCGUdSWZ7sDYZbCnQ8J
QiaPU1eTmWt08/AwwhNs2Kp5YfwlM4OnxEVdPr/U2oUbxPiOr6xeeIPnKIN8RrbP
O+0nuS57O+8hysgHHB0qBPueOWual/PmpLTiMYD7BtbWgbLZ9nC6KAk9PjydLdMn
OatfN+CWSOau9OqhzkLUuLtuvmvx+WRi1g7jKzAFra1p3aPJ+MzV3mF1csdAwxt+
22WTeuP6iJLPAF2QztOHY0idbO53t5iF90co1Rm4TRMzUAYc8kHTpq8LxeEHCvSx
yyIlgA733zEC68S0HWbsG8Esnh8UtCO5kX8k4X057/3GeZLl2C+yvf9oIvYmw73G
5gQCsS7dc7X2xUrj799aPusBpLfqBwK5Kc2IZlWfMgAYI+nmvngNv6n2VSgkfLI2
WdnIBhi0pi8p7rtDCnNIxx4itZdhMt/7qGl9lFkGibGCon6g/kdqEZ8OizBM4fR9
rQ4oSUgA7CYpZ4HiLPljcaGfrZ18dqIdpSUzD1MVaOauK4db7mOreHPPtOy/P4Yl
2LvNZE1hyzx77fu/RI3fm91FLmzOjLNZjOuR2t/y/hCUYSm2k5xUaK5RPAK+0duc
tiaEcmnmc21O3nBDSy7BNnIjQIoaifqf0aL+zNjqyoIzBlVM7fFd0qij8VVi+Q29
zoj/IO+FT1J+V/J71edu3SM2r+fLguZhY7NlxMlXM55uJ6b8h17eOCq/NtS9Y7PI
c/EqHwnhJdLYqombFa38yLzvgG/HL1L1luxbUHpZw+ZHI9sP3wV7kMBK2T5Noy2x
yBMjlVPNuJKOxfMCFVxd7cmAsuQ26r1h3pYOyd8HcJJgv9tdBOuju9IGhFrES3gM
G2NAGpG7uyF8KKaVhVAZGW6bDuJmuTsgTUSci0fjEi8Mns6iS53RvVg302+bLoPk
jFMJoKNRdIwwessc1fQ7OSAfbF2V5vkxYljdDCzCq+tR3s3hnKGyFC4NT3qzwFoF
aMuefYpyH0CYkANGjMHkb8xrJ/Iei8H1orRkXSuM66DzCvMB+cae2uk8D1V9h9Wc
rjgOBvrklJo+SR59CXnXA/C16jCg63gwKg51nTTDbFeYNYAOXTr08MQna0Lt4zUH
FmEyePntwSCObnwL9WfzgTxrDtJnRi8L+wxO6kNgIN69FYZ2m4W5J3OcxjdFpKuv
0ezxp4pRmvGrF2vWcPwBI0ICseezV3OEmSdSRv02vQE/hPQw6JQekCAtvkqMmNl7
n+JJz6MWe4VXEBVvaRecvHkdhcuPz9kRDkq0DxoVdGkbozaZmiLt48Bl0iVAgEx9
lWYGrhSjBDuirVeORi3c3PadY+fqKkM55ky6oCKaJSKkQyn8bzcdnmTFu0S3DS1C
y9cByTRWICjjV2J9mxxSoJPPwW7GnNyq9xT5et7CvyDrI7o8846rD6A3DeMAJMSj
DNQQj0IHqhjXr1GW8SpN3kr43a0Llr99ZNgZLmlmWZVPx46KOTKUXYtNIBa/u/6L
H81meAy4mK5rFx+lGHrRoQVOUPb6+kIPp6bpoheZrLgPpWiOwx5zh5wGLAX8PKGo
6xA2+/dErW11R2IhRpeeMBeurbOPIC0GsxEAFIrqduRc7IR2FEdIp7LH5/sqmWBi
TjrBjJoea0ofTgz6xJJOvW/+28foGTKKguwE6uKvRalN60c7pdYaXCZpIXPR6VkE
CeYJZ4HaGHLchFciwFyGXQolog12O931oI5gt4OJDnSeRQrBN2T5scHu2VQSeW3O
o/73NkGtRlYefFOcZom0UiL/oXvKHkcwGZwN721ha57WrjM5vIwBqP+7wFho/xcA
90KyWK+LkBrpn1XyhcvR5KTireeZDfTkTJsLTlphnvMhMVKuXJQ8fx3kENrTjV6X
nREeF+iy8LjlBmw3gEPPmvG3eHSpFce1V1i2ReaYin/bmo3lXZ+tKNr8Lo1ZoVNI
NmaYvmSZiZdJvx2fDHVIyBN+DpVG3ktOOs6oSDYocgUnXzGq6ru8WOoeIlBrBN7C
y3lCzBKAOyQUh+lfLkoQxbp07igtcmCXiM2LEzx/hQA8gSDAK+8B2kLgk4sH2b7z
m3b35sSQoFjy/mZC5Eu2Yuj9PVnMxjaCpPFqhaSB1VOPxh1pzn3mFIQSamW4fS6T
QrCX8vJl3Aj4XRZbGfgzKlcAYf6optjWf5bteOuRQJjZy6V7cESXAGBYtKd2GpG3
y6YTIUEdHUdEJv/KrmC8htnk1WUk4xQ6GbpAXzseY+5M9e1yFRGvXjHTsylNocEY
gbR7J1QrZNmZl+kbFjvKvspNQ6hq02eWXsqiyfU6TVtz6VVcDjE7k8xhi/JRkE9R
FZQJ0bfMdLURBEELS5LHjqdaplZ5PQjR69tDvPmjOv6Y/GlLkgoJZYp2g9bkifJX
op7lxs3jREUROw5xBsd0ddgE5IC/CVcP1foIWjTNt6lJ9roKvWzn5yvdZfSwavI2
D+9gP9AViRaqmBf5K76ykYrh/75VNKLu77ydiCM/UGe1k+xhoFryAqvDUpITiaSL
gk2+jTeoQ0Z0D7gbRHvsOrWRZB2/6HknoIfOklqxeyQVi4Fl/qXa1sRuRwur+dXi
MjsQcYNXOwKDSNKToUthlRAEc5NAH5UrR6P/yGdENemH3MfWGP6IUG4JudTlQZvM
tzh2HWB/16cQyQhjEGSjUZ3GQSMgHIEe356puNPlw0l6oVia9LJ1X1/MI/mWKRaY
OoQaQ5OzsuL5umFK4SPLe+EJWdqI6l3JouZdmOEpz9X2okQnT0tSBZktNZ4aOmwm
zFM70ILTWDNPtqDDn17ht9xn5G6POOtb+EC7n6xpdzRwMTPfcdUpzJJH9a4hSgad
Hi0sfkmltpA490TtqDPRL7JPDl9ib+5gUK1XgyYFI8whDr5Z1w4CpkMacLbhiRFC
PuxGLkNjfPCd1xvyHeLIxCTPQhePmYgDYnVTk8IGid+zfmIYnasHiMdtANOolXFu
0euiQ1IWVpD9IVJF2upq1e8VSgK4rmeE3Z04ALNpdXGm1cHEJcgfGtRYwI8PHUW+
ng8R5OmiEg2NKE/Ouco1Dn4PrRMmq5T3GJMPCfimKn2SWNB0t534h6yRY4BB9bVa
Ahuns5GyKGa/jdq7XaggOFD/uDAfDzSxsnPSNo2A+94cgA22LvWKkH29ekuWvOrN
gA62QEKZzReFdroMc7OX9bjITHDnj/1s034xJMznni/ZA6z20IrY7kiMfwVUbkSx
rYMTJAddEUOmWkCn5xG35N6vv2Se6dEfTQma2daVUM3mvnvQj/8ujvD765TfUkos
f6Cvwjw+PNNMAqAPWPEsuD8UGpKchLHx1rmsRoAbIbazEgmu6ErJ765Vw4N3D48Y
p6Fd+5jrZjG4MTS8nVDPNN0DNs1/6ugXZSPN2bXqutPSuvFfq+jl/JHjunGDGKNV
kdCCgPR+yoY1p77w5IRZzuUKahwltdojM2YSys7vwOxwMykg4jficTr0yRislE8E
TUlrME3Zj9BwZmXw6nbiYHb0iZ4i5gHSDOSZcVCOxL0KPy4MrVrDq60MoWOYWhgL
2E9IGfhuoN6wtR5Zp0YiTok9AP1c9ekRzFc2xCq9syIbxzPMgSjsYbUB05TQBIzh
pOJKm5D9lM4D6bLtxZMD5d2PVXP3Y4eaLaF7EsVC0x63fPKpL5DrUG7/NatS8NHj
cxNj19/nlvStI+OKTVDSUHz01TsH9CMx180p4PK2ToJL4m/EfZ0TmLaKuse3OiJX
uD6V5QCp8CAww7WC9RfsTeaEEwT1EvNvJPJ2vpbOfobuawho9JeMv+yxshgLuXz8
wSQbsMQQwzEYhv+jd88NmiJVRt4PZG/0Dgr7Li+4k3JZP98TXTuA6sdcCJs9nBw8
MA76vD4NW1+0wk2ZlpdE1iA+BKlhUaVYvHLS8xYnTNYZcPkDMq4cd6eBqxSfLpr6
v+RCUsXri49pjcMrZDl3Ngeq4YZYdxcRLODt0JKeR9AgSm98y0mX/vPSlCgzs/kw
xKdndxGWisE/wSbOTWUl/HPlxZQUyWl7xtrbEC4PCGiQZWkYa53Ql4Gg1D9bMoGG
F0DyWcOMSOVP8r5bf5NaWzCi2PEREB2FTSw1p5/nrrYJy51be6tSMwBimzD+Ec0C
m310LeDLM9rI9pcjw/c9/mYOy4uPCYazQduvg1FIDvhltmNeg0AQ4NT1Jv2YZs/8
RmmD3BNiNZybrr9rYbiUfYTLOtg48plWtkgm0ZudAICaPKExWUtl25JTJ1oR96fy
kxeG/W8IRplp45Bdu2ZxMuW260EpHHU/7m+DsNsMNoaquKqrh6icei4uq6otC/4b
iVQ4ZJAxBv12+o9AtX6QEH6efsxGbHlPLeYF7VLKXieaThncHqYYjrjGS5Fut+V5
F7K2eAJ408356i8vG6KG///2F6PHzIuNlFaEwgc1Mt89c7lAS36AhaP1PY9Uf2vv
M4IrUjJoYgOgY8oiJKG7GLV8yqaHFD3bgnXjhd7NUXR5VhZ109gM+laGsUwz0SZ9
jTeWsSa6rFMvCr7AgwTgDqqB9/3GztWjlHwwO4kYHliY7dxarMGqeqoOJH6UEyAG
ZFPG4NgANtyCd6ms2Tgt662+wGB9nD+l/doxSg4E/Qwa+lL3jszI7X/lcvGqkjLQ
0PhLlH7s+BPkxqmRtzD1i/Dh2++4XFU6EZ9fUJJijR1kcsAMZwKIP6MqHnDCq1OL
Ome7jB/8H/a2nn66QemmohCZ4kMxFZ4o7NrnNeDMKUThscxsG95iib1yEboSV5Iy
oDLLNs2SmriwwQqCk5+/ohqHAD4dA8YXL7EH5T/yqFqKt/OxA7LNAnIHMpfi/2UL
IXLAjhg89lvE2vAr1v76b4vg5zVu+KHyX2g1RWf4GDzA3Xih56DNVmWG0vX+jFuq
hl08eelH6mIoVMEza027KR+6R+NM7DbY5jkRjg2g1BW6XOO9nFgH/a7pbXJkPf0c
kA3p9WStPVUArn+KtaXx9SbG/HVx4Aie/vqIJ4EBlNne85Zoaw5PQo6jUHZCJq5c
IJ1u/6Sku/GRg/SzNU30tQy4hsfjL+92LovYxcOlnGjXTNA28ZxG6pj1DUz3VRZE
LyjftMLISJnYkjy1Vj1UtyaKe+54H9Nc979+cFfEkhtCOU5IJHubPZoqhLBRLqQG
1iw1i3Wu4fbB+JqlOeHqcuGV4lFOo27IpY90SEOKM6VUIWQtxBn1NTTp5rBoVawK
fwT7m7qduM/X2oWazf/HhgpTs74D53PC7Hh62ebkZVvwJVm5vAW7woIcaCjn13zr
ifFi5iCXGnwNtbf8d30shKShiOfozH3+SMjbTXxPxzE7HyZfZv970QjHFjoBtFLg
8efiyv1ivAiZdsQeMrjyzRgMLEH2He2p3HfcfH6DNwAMh/n5rj+NOJqPJgHOg23a
5bAGqfPmGdLn4NpfBtfvVCQVKTLqJDzXZGyjuQ/6OfhP/s9tHNqTLn6mbWs5Srgg
xCNTVu0cGYcIuWH0mN8ftBpkxeaC13jmyluzgUo4Bx5tYZiuoz7uIsc2G8jv/mF+
X4hIougzRIIJ3CDfttKr5ScRte5ygBkinRdZPXagXquqTuKE3PneZ4elTyM2eAzj
bBaXKEMdL3WE9SM4KfgZY/IBbFw2EVJCjY0/+sez3d2BzOMG8DJZFPqrVUX5s4UP
Ug9oT4XhN/FQKe/lGR9rDDjeXBHl85pRmeaV1aUYDcs8DdouIAqILBo1OQDpUUCJ
EGfaVWBjJ3fgDbDWu+UJhUe9VRtr9SpDyQ5aBcIGBmmyEiZ49o5WxuqhtYXi3qHh
32r3wHEbLo1ZK/M2UomqyPYxQyfdLXlp4Ym6F0XB+dRGOMkw+Wftlv2pA1HjFElV
ozdwa7VvN+nUvnQnkvxJ+6A1/144co4gCOEXK5Dc9c9u7O+baCGTIhqRuVEOD6jI
5E2Ze4Osx3Astg+fX5WPdOHdIKmv/OxXgh4mhXAtGnKsMaxhdLmaV0OvNdQGTEDn
D/TLuk82sFpn7zY1PhvaHbPGh5lzMMDyFhP175sEldXycHAvMDLW5rtTesxsgWhR
H9GORbxUqbdXECYHnGkv8o/Pexcaqm3FLkZYeCMA0Fw4l/kqCml/hx4LHnAAvpsh
D5UQt7wMCVaqEWtabD1VL/DpQGgDSLFMEJhsKNqJrXzrTnoxfKKpSULQY9QbTdKo
VG9jjdlSQuHA/5CoXgoMf8gUKfXqIkEIC1yRQSw9PO0CHD7IBy7XZ+JT02HeEnZt
CP6zYjzg98BQiXB9WYYQRXiIbvsXRWG0d94/pHISXh0fRg4l7FytvFTqDF5bkC0o
zrOxanbSctjvf1qKcyS/mqivDjuApSx49cfj+TP6AXUYWZ0DfD76vIYIwG7yUtO6
EFFDlRFnI5kiwmXwrBYX9ojagUKMvcOoGqHw8wZjkGQWLKewgxUoxmExsfK0/IvM
lHPtCdGPfJV6rYqMDULREEXgtFFFHYpg0dpMUeqjW6Dj8tDXMTbj0KdRiTUfc36H
uo85sbuZ5JhsHdmPwJBY/9M+etf+vRTBMnxSTU7Xnu0x4QqdmoQFsoKqZKsh4VY+
YnsKJq2Zc/t9EeTGnSxJbUGKBQtfWBWuB/H+oRgHtUhJuFecJTC0xkVQWoWpD0Ba
RSCiI9AKB8k46ZEneYzSXTra671uUlt7jN51BPTAo6N34ZqydsAOfN1D91U148HU
P3bnX/ndoR1D1VNEYBuCZw5P480WXrslTkWXGq5I3Q+QQvR6GoukNek93/P3tIvA
jLSSq/gVzKvPkhU2b4w0HeZbaWOr6RpAP1ddtUxslzAGss9OHbgNneSAhocTpWJP
ex1lD89dfwOZ/H1CURuf6Et8BzvLZ20UUOWChdmten69YqNpo5M9H5FSNlwHBgvc
tHd+z5R3sfQ5L8p0Vlifk+DG3uXWeg46/VChYqCXII6jP6rOrESzY+UvTGVZH7q1
rZxfcc1MmwI8IW5ht7Gms887kWrQQt0ZswZzgzeAiQLj5Lu65cI9LafZl62OXPNW
u8Bos5YhF8bSvBBI+EkvY5oXcpWmVqMAW/4RswwfpISxQF2NjTnx8sbvZpTmgF+N
Pw6v0GcjPv2o5z13fgCjTlmO/mSK6fuH/dRSbO6vNPx5xX6o8xr0ItSf4E8wT/wH
MFiVobwcEk3WTJOomnWd3p6Nal1WMkKkXvjQsZ1s+7pa3fmnrw13vf0g5B0NqkJ8
u3b1qYEk4kkMexfJZT82ooE8eFpqCv8tWkcj//UFLY1J+iGOvIGB1et0E6hq2yEs
Be/5CWZ4xGE/1IJk7qyzg30NnvMsHJE285ufDAvEM99B7yONi2rlQl1NF27vf5vs
4BjrWPMcnVloI0W2gVfBZ7JuVXyZTLeFHsutzuEjrU+l+5C7EMVd+RhcYenz8xut
eeHqtdoGoPlxNQgmiF8JNVbVcOPaX8voAy60r80+FqMKD4qr5KZ92aFmDp0a2sfh
RiKxVcwqXslvNa1SKeKpZC103yJgRNicZIGx8n/oueGAajVPHPfMWU5G8Kig1cbk
kY1PAxK5D2ASENKWb3HGItQwwdFxWsb5oMDbHGF8xDo04Y4SK5XabKghKlBdcMJK
GbgFadVq/2UZOIiQ3uXKkKryABUko/Ki9zcbLDBF+D0oQ//fYCXDT9Z23Oeo+c3/
F6BeeSND/fO7kHReAYGObn+/mpG448ZNLCSSo8ga0B6Pa9q36CGjoZpXvZP6XgKs
ET/fzwj9PJBZWBD26nzj48bpbOSSxtRs9x1vIa75BiVfuAjIouqlOsPg6rGLAf66
93Xc3ix2+0rEjs8i67fa48ryZAnI0eUHJU8AxhCij1/CqTiP4qRm8mRj2J6brkD0
JvFfwqs3W5HYOS7dKgzjpHNqzGIU0cjxLlr9tA4zOGYpx9HjA3aq42/OawScBIBv
IE2mprfHem4qjk44rwzhK3j6TSVgsi9Ih+LOc05OoBr1KQSu3N57ltexTySb5OPK
eBFsWZ7zvTWpRyUHwIoCwetUWUwzHs9OypohAUaPFaMs3J0Fq5gxnhRPLdI2PNR6
vZaqJOGWHq+UYZzhVAC04G093RMe5QhSojsknHMOvRRkTtO1pKlgm+B6hXVlPVa+
LAjPWJfn7Kb6p00YgavoSJinbU08KalHqGD8xO2cAXlIZEYdUuwm8p1UicKlzalT
VJ/rVgBlVmeUEnHV7YhWgMHZHj48RYj8yQF5YTQn2IjFTsP0etRlWHHHv3NmWz7l
Tp9q1kGL5fDTykEiNnoZkX53J4UZ3MKBGg8K/As/xhtVN5u//Ga+P7yLrjjkcItd
9d7XjzeUi8SGWjTvX6bQ1vtvjnJHMKq2XYfcxQjpoUxwvSsaU11H3AutbN7Xp07g
bIeLW3TaO4tTSY4y7+YigSgT0p+G6uEz90cx4A4MZQYoNoQZGXFMkNse3unPzebF
f3eth0tNxgQTPTv2nE7pRgIGT40qE6FNGiZhCY5VS9+vMQR7bxhJgV0fG+gdw76E
Peu9o3RYx3wUb5dJ17wrKj71m8rbnpJNoMx/uOLBMMLMe4HWn6O3Pfb+veGw7Qdy
jAoquHO5R4U7ijLYGO6WB5DUPlZcjTYVGqMDbs4SMYnE26O6ZblSDLWOckbF3lAO
+Rr14rc0elEwivvP5aP2UqmvykvnfgovOyOvRSfpJ0bC2cBbQCTQHA0Zvo8mcg2U
Pw+GfTIQEYEi+lc0sWQzZ5hR0i84kEi+2DbGzd7Q/WSijkgfqlffqvAonO5YalWt
1e42A6KzWhwXkeupXm2Pq1ozrhO7xRWokqx378+6SIrp804Q4IlRzrlQgYA6/jxo
en8sjQ23t3FEQBYEdbWEPNznNAfyCVf7YM4wfBcYo8sa6WmCssJ9hANO7oIvLRXY
V1+dpzeXGtOYbAlf9v7WBjXBc3MHCCvbKwiG9BhDaWl6cuMQ10gHZ7wzI9tFC7eK
UPLkrirOXGbF7DfvMGeTYWzYq2JjPrHHS9zS2rwYICybkX+59DC+7hs+jmOTLQeG
TpAAf0d4A5+mNNupzY7xVQVZEocccuVI1pfYira742Pw0FteB5HCbX0tWmpxya/f
FLE8Cl3aBmGgqHEEpnISSvx4fTWZ9BXDR7XiSsl4ottSTUZxt3yauhc7sAPPlJT4
cfeIXcB+npGf4BD0zKcuo17MBt+Q2RaPVpwO1YQtNpNU74yTYaVo330tBBICgUfa
6RL1AG0BVEPXdqN1TmbX6qyeGcrBvBocP2xK75X3T5akqFl6OEiByRyzMgKYdU3O
u1h6TyqKq2AZoZrY8js/FqQv9ybYUgACveCcZFgwyNVEjwMevZc3GTGXlcFDPgwU
TiuV4S4UqBjr1x3pyoMEPVJquu2gCBEtlpJuHgDLl/uhwwewCVQc4C2D+/WtTNGp
PvA0Zwj6uPmjrzyh+Mn9D2XQAc4UO7SfKKlbWi0KJGwuzBDDx8vd4dHOCF4hTt5a
LwSj9rNiJAbyhrT2umKycydL5OZW3ZanNbOILnl2mtq3u7OwYPJLZ5OabFyywiUg
KBXk5C9fpKG0+7xIrK/YazPoM9zZTy0OAyerJhYpsZEnuTuIpBc0KPadIz1lYxRI
jrokFTgEHtchOUUqKUB4lYleEahxdg6QkkJd+S2Gws5dJW/O+t1bi89GvAFz3iUw
1SkoYGl3SU/3Sg2ekNbOrgggV2bAuy51sPh8Vs3triqJ4OWFDraHd9LcGbbc+V3b
6xAa5fmU7t3mqJ6DUNYzr7V8Bx8NwQxQn9x/xbPNynFp+NnDdEG314IuyWyUT3do
ZOgeEJ7uxgHnk2qvpsVMrETjtawprNpdNIljOFxLPiNAHDJK8X0G5lBn8wjf3k93
wwxG2zsjtJDLn/q/pPObh/BO7R7DJo+WSZllMhLKmrQnxsvqLxAltwWesmHzB3YI
HqLdqLKSMkwqpBx0Hh7xy3EhcowycpQ6AX+XLBcToiRu3oFZx9fibWd8kBEVXQw+
H6M3CyzJMYxFXwbk6DuIxj7M0f7IpGJKfKZgL72RdH3rsnxYaJPoNEEugBDQxqwd
eYfLCT0Mek1bVGAMeAArJQ1m7Ul0I2Ogxe/D06RlDiG8dFugBbU4g21LQ89IMuEs
DePin2Eq2bQp4XinEt+z5ptXrnK1USPonTAomwRm1nx8g3RPBNaMLgg4a8tvqsFt
pi3S4U3f28muLjQe3sLNliWqi/d3u9wAJ6Yfp06s8th8++sOIvQFGGsRf+D5T2zt
6jXc18C/K8FI9uVaIG5EizJUGDY0uP2rv3a+gwVWKWdsCFrDwbBR3PBPuhetEimI
JsX8xVOlOOwv579+mM77WkFjqbMTUaBoV4GaraNlVGZkoZWwvwQXur0MhnNVunpm
LXpOv4QCFIYuKgjcB5tva5JFHhgbQhCaz9I2nyqhSb/ujT9OTcGLT+vM2FmxkW+x
LmmtM4faJ9kjNASbRl9ndlLoURNQ3ScOnkyd8vhRg7N7q8woSU/w/mzq6PQzG0lD
wPwjAo7VQ4ltgnJ1ilxvTGK7olZxsZntcs7VD0c+7wFNq/pnPy+FajWW4hjVcT2Y
pDoUPTrYEf4JwI/NgvbN4/1A/9WNUIDsJmDWURHoQXO19H0tdseKG5+R6tujnAPF
KeoylaF8oNE1Z82yt7Bh6gepdLcDnSPR+WB9O9gURTNA1Cn+StS1A+d0yq9J0gVU
ae60sEcFIZvzLDq5osvDJW9D5Sl6sfmj2L8Tb/fuIWTyFdsipcTRQg5ajsuY0GCx
u08TxQJQ4Rqhs9aqKXPhI24o7Nt9+Ky3GcEslwn51A2DCfbOXNYYGnNhvuudTGFB
VfKjcKiR+S/UdqBBcNV4VgYBCYJIT8DLJ6Shd1KGAn7EpqTM79qc0Bxyo0rAVQft
VBIQAjpWqUGM3yiutyQq6mg8Lx2tzhIn+C6crTVeayGYOBP3zEJuASxpRSiakgEz
rDFmqD3cKv5xy4zp+5NXb37mAYGerfgy7aEOGB9WuSRvGEWmuc7+Oqq9Vv0Q4toE
oAxj+YzXqsTDT6WgDhgj2VkI1t9kJh8AgXVVnERk2mqWtArGEINZHBh8hmA2Q0+p
83PCfeGQuRu+TYcEOHKrfZy1pi+SZNAh9Z1RCN956UcwpgkbgUY1ufXpRsJj78qB
Gt1zK7aDUcdHrlKk0f4Yk8Z31qbv1k1N6dOt/d1oR/JI2RYId5MwbMZK7wqrxKUn
mcuiaz3hGTzau9P+2ATP+ytA5NHX/Sx46oGkOD5CQAj6RNspbFsYxGClUqqQvh7d
+0k67momDXoQraDBsnNL0DhhagnO0/2Ai24roa7cuPANsR382KjVUrNuPVfEyKnd
+l1mcJL3TxknEj69rKlU9pkm9zPrN4KUtuL66y53Ajmp1Fk2FOlyMV40XBzL8yvX
HI0kPgVA91BjDO1b6WaROwnVUt8/PrfqFRZipIQCkttwLIk18PniFMh8JE7LcfaN
e+WSp6X9BrQD4OOC/vh/hmq0jhSfdijXkdsrOzIjD582UPZXQYFFdTL3vnWpB++M
9v6YVtFJYrIqlrbDAn3YeCBpe4iaHJCPMysIe2vkLBUnjENtvnMfRrDR2Rk9gQlj
QmfqoQMrZB3L8cJFV2mByynlzcn7Msr/17T/evnCFFBesypgnnOImHkmFS5Tb2o7
JgqmZ6vdGUoDFhzJ5M7EuGn8JxdUHqAkHsvEfZG3O3hhWPLCCJJtQtCwmGoDxZPQ
E/M/zSqDYg9f40UG7WpZEfHKTsp41k9Oiwlz7f3MvLh2k4vX9llbvRAvp9tPTEuR
aUOnDtEZg0sAHSTaBXVpNvxK+0J4DRGkdR1J2RscPXBJlfZfDsINROm3texQbCSs
U1iriL/SjoI4hWszPg20yNpYJ5t3lKJAv24/PCM3GQJ+BCGJqqBlSKpaJvX0NV/c
AAe0vQRa21v+BGoKBgtlkfiekWChwp4dIgQa5unmqZW5oXxU61Fth3wAWdmLf8lC
sG1ci85/eIXfb/Dv3uGvM1p31nDStM5I9wOQEVxK/oqYbJcI0GjLL+fbvypE8tHX
V0wgZBc8i/NH5ulZahA2XoIZFkIwM7J13XFXuvWNCQG67NEIaX8v+uK1ZFGqlEeF
21T5QjEPhvrS1Uen5gLhRLMdxu4r61yOq1IwsQR/wWu4nMBOYV1ZxKsT1KJZqzyG
sWJCk7CH3p3z+YTa0wbxiGlqmo8qV4QZyqXFeZRTTcdkxPdfw0G+tMKLdPREXRfE
w2R0hYVdvCEZCc0wjLBthzDGh/bSLNi3DeItHjHZvRZkSZqCNTtwt8UEnLyirJ5z
5mQfg2LuFWM3VLv5HFcDNk2X01Npi/BO5MgoYl1dWdwmQD8KH/qd022q38CCeUR1
52Lgn09mN3j1AoZpJ6DLkz2Sz6Mil+FrBD6ugNcM9jLpoPprPq+QwV+mQ5gA4rtS
qLzgUIH4WW6ebLB3v7D7KHxvhkRny0UIbayRGMJhhy5EZFelKU1v/N+70sjbvLTE
nNYaQpTrs5YpZXBLrJZAKod5qhdf0CbC/E/1VuBJIdb+GH2fXjmdgfhzQbN7fAdq
bD68oWnfznuL9Vdae38MOsyPiKcX6mcp33hqTzzrHoWzomeI3owjfgN7ITU/4Zq3
Qf8DlLZIJtBGa4ILIrl8YxXWngAwMqlgGbWFq5TGw96q3zNbFD9YUcGDKngnBrje
dj+nYfhHrvbILSM0PvifkTTxXqtzr+O25+zQz/C8GH8zz4TOZJPnxaxrTxNkP8JH
bbrIWIr4UzPngdsKd7oPWAa7SMWfCKH1lHKT/+hSR8tIB2+HxvHnkd5jfj8JeLp3
JJ0EHUqVCxVeDT1WontkldCiCiYrtxgRsjkzQaDN+4ek6s7UmqXjGOMCHnB2SNzK
EG+nexPlyk7OVlB3Kolso5RUBSNM+167oo+P8f1asDy68gDZeurn5rCyMn6DU5fO
raLroXSaxVLtHU6Azb+kvfrw0Efz0vwdj8MmUaCJcC1a+d/QWikxS5Jy8ckYQ7oD
3GDYmDMXjldT+RcYXEQeezsvNjFJz2qJJOKJ6NtRMzJkn8wmSsSV033v2g/0B5Ao
fj05wvDjlVmi+8cTYy2pQ6SY6uT3maC8oa/SEhiUVioiCxpJHg3ue9AkY94eW7dB
oqfw72GQ1WR989R2WAo5m8iOb7rp0/xqnFM7FpZUqOPcelLJDnB71t1Ho0XW7Bqg
ZkjN2SBlP2lR7ZiD+g6kxMdt8LaUoZffdoI9hWtTPpJP4dmyhe3R+0OUfrtG7gBo
5yAyeXsGhpxJUNPe4qKKENJMjMkU15W3Fmy/QiFShBYr948MuusGbpynJh6agoSp
BbQJVV5QQnr6F1iwsqD9QruIqj2dvuWBpOEN2TZFSuiHQuvSxq+ZTyYvQ6sWjyZa
sTY7SApKl+dLhcU3PkkgQTFxotr2KUJ6gx1ROBX0hlwVy2kzb/tvMPIxEHOzdq4V
epj9hNineGq5x/lrVwQHwFBePa+LrI6KyZYpeBQm2O8gLEvFBOCNVc0VBSaicCrR
evE44Gm16Jg+gOAbcqn/LzpGTTLNI1oowLNXhORrbvwrlQUNZBd2o8LezMvxzR9X
Dbzivmih5lYmx/UkG/FkPHIm5SKVe57FeOxHSviUKVDdzgYvzzvshGO5gFeuuEEm
HC2O6n/6yZ7evG5rRUhtlrVWCAIkxMFtjzXRI8fVtp4RJvPGfHMA+UgX66ZKcs+E
+cv7wZBCVCgge9748k9htUNzdJnNvaVrPDQHh899hgSe6PdyIC94h2bqLvaRGxbs
e00faxArt1PPsTgnvTbNp0NgMQoSAysN75TniF7xpDPhJ4YfsUZKVN7zHDW16Vl/
GzJVQX5GNQkDLld7I5eL0BPTfFXU47+wz5y6ZWNu/Jfctr6x8IAgca29lP7sb/yD
OsiMf2F+l+hF3X+cNnXcNOYiIMoMs1sug/EXJ0XC+tQQqS+soATpTqzE0L8IxtMd
ncOsxvXx64pbdXjOH7XqydVDFfIXGbWlK3u52Q/djNE8TzHRMJR8qr5InTL9G8Tx
eNbPw2rNhHr1TfrNY1n9fheK7m0domh5NhgQ5NFSuMXpVY7FSFJc6gzL6Dl62+4z
KAcCogs3b2UsVRYPtVy5sXdrB0cGASAOM/B3cGuNa/ExNtPbqvKpvJHxctXXCh4T
OGDD97vQD2wSh2lyMfo+hO2BG6vCOX3YX+1RbNp2iou00RVKh+YjuBB2NWbIef6I
cgjlZo7Qn5R3jymhXw6Sjj9AS778wWrwPP1OOmcYs8ijiPqkDdmO3NPoKL4Scw/S
qUj9lZppu2s+GCTC7Hw/xs1aeOqitSJX9+QUpioZBMacZSu7yRWnJiDDAZsnRJat
FoRiQyyL+ptpmnsMUZaabGjNmHQw4bn1/fh4W2CIDzeAbFIGsDvYC2JQ0dL7ho/C
9vhTSuj1rtmFW1EbhtAYaaZa7TC580btcT6eP023VV4Uh4K792qLllRufl8lnp4A
FdC7eb/wCAxEXrqD118/744j/+9goFLH46Vpz/JNX+8eWoonwT1NInwS+aUAR/d9
2g0J+JojQJKdcwGMC54UxsEMfO9cJhcKZid5mAhz5Leqqr92HynzVZoklijTKGM4
8Tsd/gOi7227vums/kvacViI1pExEbGNnewrOi40g3mGbRhVpPhhEJCNxlg7iGMe
ZP3zWqYcfMxR+9wpm16FaECH25d4qSR9tPs0xCcVCTeI72oip18H8KZvBwevKVJN
PQ6fE1ZrEdk2ATMlel5Sq47qibyGmESxbZhOfLbY7hIx5DwrS4ONjbjgE6/iCWOX
C3oSStUY3Oa23gvF3lO7hTHjMOaFMhCD/AKLsA2ocnxNoRKEmqGs0+RS8ZyIz45l
S5SjxUQRs3UNh1ga81lYNHn7EtSYxgMIDFlT+xPF2EMDslJir9rcRGVycv/DgqiK
1xldUna8rQHccVEAlI+i8/MwrKhAvHm1FvH/Psms2lv8ZSgOlvjKK0cnKuEockzm
P+t6cIKD0g8sjlXai+qMrQrW8MD32TlP4eA3eGr4rKWBhsRgsNq/wr5AcgMZ+bwC
mO/UT+4bwDIMquLj1Hels4YzIg3cC5tYd2hC/04/Ai7flf9/krV3iBzPe5PkuQcr
R0nUOkgSLI2tvZWvLis/HNNWiH7YpTdyAzeN1hm9UgykzfeA0lUr3grX2c4TPQwH
luo07nr0eqep4sj+JclSKvOownSXPbRnVh2rRNY3mTLJPimW+0YROoUp9yU9OsUd
NvttpTKxdngqD67SvMMwJhYXQOKiQE0pKp2jseznH4YtYebgssxOUqTlIJQOzPfg
eeNjGhSVrwbqye+UnHSG03NjqfndR6ZjrJrOr8VR+wZP4zIHzjWnKAlYL0+N2prC
S9TZPgBuid8aJv8n4ARgKzMX8DZtH9sYzyKprBHIIQvo1Zm6bxGkLptVkiff7BGn
Wy5Fp4kLX8B96rbecWOHvNCGcFdX0Baj9FYNvScRZeF8HVWQxOv3E3Fgen7jHQ/z
H96TAmjM8raxildZ9wZVtSA/G8RKKOB+5OF8psT8i6W9DGZQPfjfUan0tUqWuDKz
VO3nl+WSpW4QpkYA+k2hUClHdfl0wnf2g/A6G/y+LRhA+DMAaNVAme2EBi7QsvXi
MYax+LSt8A+6YiE8KBlGCzdMC8vo8b4gzM9S+WS1KYuiGq8ogrluyz9k40hqtBL8
Ep9xz+OF8mOuSMiU7drWnpZwP/x45OnOJegVtZdY+UygBWn/fXEYyCFxtkbP0FSo
46IhmrWUWvznwk7E7MyCRVzOQDmUNq46hgo2yAPjhbBNbrVhiEdZG2M29VoAnvc4
2H9FBMQfBMK5IXglhD6A+iKu8ExTybZ7cWcqkw2RdAhJt88Jo2NuQtD/edtNGWqf
yhXpeddFsjIFMihb/sRCRTGoOeGu92ON3QPaZ6PCBczXpBCNgbPUWitjKgvvz6Wa
++K7qR+VsSs6DrSzJH4qWyvkLdbxKpC2vpDI8ysaofaIMJXo8wZSNj8NhgC7xaKo
cthHigDrXRCgpBoQNrzA0SlraHwI2F8mFV7wIIch1fg7hQD3sQu0P3iPSBFs/rFS
vbihTUBqvH8sCDARPuy7igwyx808anD0CvNk4PrEfAXFRhpWeYqe3IVmJALn9BQS
VohXHI2IYR3TwAxVVcSZIiBOlbW4EjhOK8aRsi7fegYXbjO6opLMVxF62aAyzhcx
VV+0p1JdayQfYmpCuyGapMlKH9L0UMFbug27Y/NP/R+JTE4pFjyrIkewUioJETxH
kQpA+o3U9kCgvQrWUtMQbvtvug9oJmdq7XG5Q5A5uzkHQ9QiNb/6LUhAS8aocgzH
KEFtprBGOmwnX7RHY8J+72lTKj3X5QbsSCykBA+Toya/ZJr4GuAvD/skb5zzmTme
pHje/tP740KOdtb823eYSfzTBT1g7vzUuEOEitRWWw2Zvo3tgqwWuh3U+PTUrcsl
r3YZcktPXWSK+1LrV/FIYCAdVnOSk6pd1dYfqjYacH3AZq+VeDWDdl3SQRc4Ybtq
sSE3dRMbi4Ur1ZHfw91r+vLOw8WGOaMOy8k1scRs6NU5TleN/CBwiwQnyUlu/Zwq
76lpy/BuRXztuUkF5Yoh18d/dYYH7AqC2YtqH5UiqF7tBFcZUCC6x6PHko+PLOWd
qkLUdURBOD2mYIpl7r2YzOnow8/K5cn1nOPUiOuv4BKnO/mPAXpJA9T0LhroSxBK
GP9B8h1NezsGtUjUfZgA9ociOVpa43akN//FSw5kqS1DT9js0kkMyxlnQ3z+cMiX
IzNaUvmLkq9NkSnSp39II5ziXMafHpx9FrA1++LNydPdFsLic8ry/pRTJLmOA6dx
EPUoBItF7cZynitl3WOZAOBBjbMRUUDOr40vFhBCKTdwA4MnjuAw6kDL2iW/PHn6
2N2wLsJnUiooxkFmTJjY7HanopoeMb4beMNzw3UGl5tnUAyNVLnekV8jQDgktkWC
w7H4YHsPfvAb3huU+hfXLI8ZWsIujVTpgMRS3ngdbfqcDkMcd2oZlwoqcvrag1OS
vUAl9AzM+7JTtVOVY7aIe4xRLVlg1HwAu65Rt3FHB5UFBWezZhzDsI7/jbUwGpFP
WJ6YuA3Y6oQmf5g2rOhXMj4Vv7oVCVSF9aGoeHlB1teXm3YRUI7DzL+tZBYNyC61
MtPAKTnvInJXzmqqvIZ3us6o28JVRwUVpDPknMHjAivmIJgrsfNpZuaVBoM0Xvbz
4/UAb6eHV/gUuP4A7BKM0PeRgehJi3hpQ/QFqu6uA5CHIKAcJjasfaqE0uBR2H+J
zRIvYQcqZeAsecHvwMPs5o+QjUPjclCDQ6syGiehDidOGj6sTHV8h8XkLCvDSVV8
3dIKGr1ABwDJyXfWl4xxIp7GrIsnJvjZsaugU+IpuiGRmCSS413S6RHZKDAdfE/7
9/fbyVV+tCrk/YPWyb534fcJK4dWnrnNF/N2LoMmDK6Aq4gwtqH3zTL5qb5aPbPV
YxHyH0dv8ph5mXqmtGgaGLDUn+UrMx40aAOxtmkvSREBaWs13vMvEG39ZtMh3LrJ
1VcZuE9vP4Z3+wPrBted6Tiq04jmNO3DVTpfa4cWkmXDFO1KojLRio4rZnLHBHNX
PGRtLke5WGTdubYAOnyu+12K+7Nw8bnkUXKVkO4r4ZzaABve+Y9Fq8qHWOEjoJh+
DSdVsrwhP4Qq1cCaCf0RcYY3D48VHOUHP8ujLShHU294jWGoNtt6MmIKBMjTddk+
FfGzhX4KYmATLvYDDhBLSOJVmvKR0do1dWsfyoySgzBuzzQeJeU7cNH4ACa1GaVI
pPis37THwZeAzT7Em7+AWQQE5Hu/5L85657BDp2J975WZ/5TUY9ZIiYAix8uYxa/
vsvDHLL/H09nBNts1EJ61iDXTKO3HLHHYJACY0Hk4vr9iLZBKBT2+PZtBTB0hPW4
FnFnizmJDi0qUbldhLuFPT00h3lEo7g/VRLn7+VaPHyi0z8RPvePoRpvZAhOjx7Z
VHbUkU38x3EVsmdBjhymKnWvEHfWLp5uD25wTOdKhq/Y2kfEcdXiIUsuLVQzSfw8
Fpc5M/iWh9TmxKBP8W2gvKLoHWCoXYSTJwBBR//X6iOiUTOzIq60L/jXTxlPRgkX
xh/AXAHUw/j+GPoImmxqz1K3h/izfQLsUuQEMKJxDiG5MFkiUtunIMT9zskjKxO4
+vHW/p8BSxSLGGKxNbujTsh4lDeHU661zLwvKZvFjouDNkoZRMx78KLTiHGPM1mw
goR8UziUHetKKyr/CPPQgNjTKeTm8seXJIG8yIsH75Y8xRoZeXaRtsA3ncpMuUbe
ha/3oMVUCFUHThaZVpZuZQ9w5yqNu1KofQm6jMU17iVwHs7UNxn7YQPxxE/6saON
EOVXRsLJ9Pw3ovY8x7pfVZlajrYcDzryUuqQh82fEZPmqT3/RocnCR/3B6a/CgEo
zVR6VmE/f7rpfVJMaHZzl9n/KH3NKfkNlIUEHQ33GdD5vQil68/Fm/Auf+QPA0q2
5TweeR+Xl9HOcPqzfWFmlb6PwBxJ6RuK9pDxbYyoMAy4dLXOb/nR2+UGovieEfj4
6ddblQJcy4U5qWMbS7K2y9Phw1EdtopFOc4Z7BhFNw0FIt/wyJ0zLvnJ2T017RIC
C2U0ZRtCP6DtJElHcGnz+7kgsbr//CXl7DAxVH736mTlUzWrh25sBnHEjVRkaRSu
DdnjPsk7X09t4jfBNh5fTL5bLmKVCUgiqLScix8Vy4onwEOLNCrk7BI+QeBHRkyy
L02yCob3QmB71VhgwNln6punqSaXIBpf1mPnoz97Unkb5WgykJHO904meXxDzCSa
UKXioZ7jqHfAQzarybpC/5F2GEhyyL6D1AujQ83ROWHMK8Ggra1bNjxHVJLEMEx7
eVKn6Orv8fsfG8WuWivCLh/yNHHXoVl49Qpaddt/lfdPuMgpG8+ivgGigtUoOtjY
lqTi5htxI3cGqQ8fSlGmWsXVsZ901FSO9LT5IOplsq9OGmfsHkN3Ur0krH6u6Omw
BnNweNtThKFJgkHS1TCK5xR22YYau5dSZJvv3P+zC+3d7Wi5I0cPFzpuP77SRYWb
+qYQ0VMtz8VxHqAEwpd6hT2Pvx39Ruk2y4TeGUrJqMfJexq1dS3P7eteuhe1CMoA
KoytwWQfs9NkJJr2C1Pjlwgtv3n1EaBz1VROwaE+xKMBk2S7p/jid5eczLDrhzOD
a13poWUDovCf2XgacqjE0r7wVBGXyiW93mLukjpwMpS3uoE0hXJEiaeGYje8tP6W
3dek8vk1yGfOS5wmXjBuyQqOBXmc/uCo1ZXN9k9n6wiHanWu0xoExxw2NoGVq3HR
/iq06VsocUjLNfpffqoxzvvi1X3pCzFGT98ri70c5DfN+wnXcsUXOj43C/giUXYF
/3ftkULGvwvxNmAD25oWnM07uij2d6AOShArNsBXpnqevFMcCHZlkklCVIUpbmUO
yg8nQDmVqPEufL5rgFUV/pFcVc0u9c2I1ZOsH7uDYGuTJQ+Yaj5bMEZGbJ1EbiGm
DdJrhc3hVycTNGry5g9Y8dksPU/G5u/iXbgCg0zl2elC9s+mdc1l1JEko8eBG1Sy
nZYmAWBt8Uteczv5aqvSwMBgyglXsPSy1KA9oKIFyaboiGX9aqs6/EX6YHx+oFsR
cKUqoI+4QS8zEcASQYils1kKcTog0V8YUlVoiQ5YZnyJId41TXUNfpQ/lgeuodoS
vgofZcu18VcqvnRL/nA243e7Q/5xDY5q2D24JIrrUR3OVfIuQYoUBpyIGQ2aTV0T
DHV03LDk3C0m/9sVUfOzHMrOrWKO6oc9d+GuqFG+A5Zd0zokQk0KYxeiEGAPuSvH
epVjT5qZFZa0dFM4Fi2+gFbBXfficbeRbY3yoRv/Y8vsJJv4JSQnnvLN4i9LA3uA
aepXzP1Xjp5YCNg1VJu+mXlyEq4dYPsGoVIZ9QC4YyZWcb8OTNML272odB2Qyk24
j+feECAacS87ZAACOv+MiYe07ALDSlB9ybsHrux5dfXoKLoBxIBBlLR7ZQG+C3lB
X2yaYx4kIQZ5KNLx1nsezMXoGBdfCQ23/43IPCzgs6guVECpdCrR1Ynn9KqGZZTX
Nc8+l/ajWDXFmD2ppSR1i/PaYAp+x7tRgE0oxn1GwU9eTEXbQuOntWgU4ENajcYw
uF3vANQlTUaDZGW6Fe83TeFHFK6dhoa4aMpS62HO4nGXaE4Wd8eT3HEuHSY8uYsG
j/k8gFFSewK+VJVs6ddBpO/gmfdK4qsm/aghHPF4+LdsH8/bFUz3Txaoj/2SAkN4
DoPb+V4imt7PKdZ4QRWnTKgkAPQ3E9AhBOTHu2Qbjrx0uJxEltiU1ZqPJwd3VZuB
/BL4jBJySV25OoVtaZ2kG/fZP2EszOsy+MqOTJX4NQ0hm7e82JoJZph0OZeiQ6EK
bkXLJjmb+8YmWU/cvC0/O4JfLqAY6MXHJLFGt+Iqph81s9nGXD983l7zQ15iMYn1
Vow7tLhywl/DxYe5BWJfiFxE0aaTzq+5jEhHIyvcGyrjO9qybCPypf7Vmrca8vYp
w1GwPfTuTY/7CCElUQZE1H8kDLPMzu2Cmurhe732tWGMCrZw7yYch46Kf4EzyqEK
3NbfuDva3hy/9vAmZCubNKBX2cgcT9LL5azazucIxk9IzmrSeWOGKK0Me2bfNHRG
vlLiXQa6Da2cjWcTlh4r7d1hhd8j8tOTa0+KMfJ9uInJTO81mQ90qmFtq7j3vs9F
H6iO9HL+ucKli/+09ic34wYoffOOhWmeZjBcjZIGidO361TFJjcNIwolRYD88WhY
qlPMJlr0aBSW/MrG+a8z6JeZEcyoKCqLXGB+edtCRYwH0HjGQ7XP8Ri45OTFDmNb
YOeuDLFKYCT6ezCAJt1IutRHTwsniUpSBmFSbZtPR2NmIAkmnY02RyKbw9wja9MW
+kOSGt2rvBbYvp6KfkCi0q0WGZ8vqGv7GmjVMup5e+cuqDXNPl7p/JfVyT6hOfQ/
XSmvMq9TDvli7+CUJK98Qlp0IUFEYEUBfduo14JNQeNexGWZqfvC3KN/M7e5vVfJ
A2fFvd2tuopmQHAAphvSh85xJQIFLMGK4XTNvPaINhsI/aHajemWh33WQEMvGCVw
vHoYmVLJlypksgmgl3oxa7oDByvPMurUTaPJ46aQcOVI8iyJepYvs+J7l/Qsnipf
T7JI6w9J44ohCkbPKbKIA6n4lHeiqdlZIUZbxxERvtqSUhk1veVrx9r1zy589MSU
MgvvE+u6pkN0v5QmTQdmcqUWC08wcK6j6IsJjfs52eGDCBuKgfVSq2ABKqIyK3IX
J7doII8xfv2keCtp1sUEzXOAGu9ZqS/BOIZ65Zmr8hM1ypp26/yM0fbkpNhklUbg
isAUjLgRX2p8z2Po0z1mcUbWXRD5wtVZBkHlndMGxyf/RHEluj7wfbIZFVbcIXZ4
kxtUXd1q0QGWtflCT4j/E6/sPlKnOrikcPDFq8kzfvWuEjhfMFloNK1pE/J2FrSF
X6vL1Ju2Z7UHns+8uStxHrNBhwFpmKi/bIrQetSi8yuLb/pQPMamr4jB5Hdr5jHm
Abey1jKUidHUZ23+V8EMXKNR1i1oPnFFNef9xUusEegtTpPE8RYYprnRUPPmwqoW
8NuH0XcxuAczl6CGjYSBylO9lJTPqo592CxF6Mig7biXTVr89aoG8twjPt1m3f1A
WdAiRUel/4w1W9hVc4p2oRfpgYxh+a94H6DW+dwKgIGr0l8wr3lfCOig2/DLtRQD
gDYrmRJOMB/KUHr+Hsz/KsiP2krCcTLrP6rF6Bj8m2ntOScTKaqes8iCVhdLhrpE
WmfNU5Jf0eWnBFcv5+BOAkKXlKZebwrAEP3tlCqtXs6L95lXRiXdHam5nMBvbsdh
BICYIyM3g2xvuhtX/Sf/T6BDUV3bsE7Rgq30Q6TyyanXaMn34J0WPLrCF2kWyxVq
22XoW8os8iWf7o3vO0SpucVhupVCccucW00CHdTTuLSWdLMlsXi2ew+gBlr5hLot
jnaHjh79v8Gu/sp1hTPCHnT7OjpOtB96iNlQSct3/kn2qIaG0Km84BL60W09YWFO
HWpDWdQI1teGaMkAcqBtSBK94R/Z7RWS57mgk6DPk+lZclHrUUJcNxz66JVdNeUs
4RZtqBaQ80iJCjauDK4gCE0gTWSevoH9sBuapcoLPpQh85mqGSha/4Z7F+cHrRDT
+/ZimE5gmu1l/TMRe4jxtMLlPSwb09drxwnrHaimXST9zu5TO4LGLcxgCn4rlKBP
RcC3non6KZqU/tu3ZJpoB6wHACa+O3gDbJLDSi5lSAA3RfsdAZrMriRVb0C6ucPu
Xg1OH+3lBKdHh6GbC72EcSTbbLUnkI31xn9XOpQwIOxI5hpZrsxyhu/6aqak7I4D
8Bnbt1v2UNtvoQFmP3ej/a4dSdlt7COCkB4VepI6A61TFg40vzKjru4wPCylX0tO
cbr3uPzyk6GuVjBBiLrnYEU7gqSG7N+EQfUpqF2mRKha7qKnFerjxl345fM2mVnD
2QL7kg5PPWKM5Ht1p4VPD0szicNKWkcdpMkIRIhrX9Vd2pWTBNy8jJn+1nmnCbEo
byWBtch/zAyQ5uqm8W0Yt1oD3WoSyPvPr+nbcV7MNFj1BTFr/tgDnPjf+BskJdEi
08oScKkGw2LlMT7Ix30yT8qYuWYPWYYnueshO4R2+4g6rpo0fHPcoBUAruBxVEmg
BxpQHmQMPD/QOZdgwOrh5wXbMBJyG9NjnKXoYjXh/WHLGVR7b1LYZC9HWvoZDxVu
+XTACqUlEPyOSQ1sQHkXmaa9SgGKAVt7rY8jJZ3MKpZ0jXn4mG0WJUvdrwCKlZrP
963nnrEWUUmjLg4v1hP72i6slKKjAzrQD5FThGm4a/BjCYnAmnPVHaIGv7Rx2dyV
n+BgpNoPCPlucux2lQg9w9wTZViEN/AjnHjvYzSzXbaq6s/3OJTnsPMaJps8rKX5
dMvoy21mwju3LcqQjFY5TA2pq2Ej0OoFRgJALMJJu2MM+bsPGncHdsx1x/PF7Dty
40xGXeeRWXl21GNHkLGruoKnzqTiR01QrMiWYgJjTCypDkJ2Apv0/VPgeqxN3myq
67YrMnFbbbpIhVnhJfZZPHGWQFJfXOTXhjjVm6XHewjWHmyKXMPIA1Xl9bj1nBeA
tJ+7ceOmx3KpfrVKsw4Q0gl/dshdJUnaf7dnWc9Nycoo18ZQXu9nLAsG6OFa7kYk
DPGlV1y7y+YH9rE0sMpOKYPuS8MN+Fl8gDaUHB0aIEa+RIfwVGlLtlA5aiNcS0+S
+XZ2hJ/MX6q1SyNNPHjhsoqtexDUDhTJWEPa+8igSnIEnyPhlhFVDLytAvzbbElp
Ci5TmUncF0d8fSbDCbBGbvIwppTVNwuXwk4w8+/Gk5DHzGqNCK6WWNNtD03LTOGl
UY5eOwEAirVCiLC6TKWiXpExlvcclDobPdWknmio7WX+R7B7d+E8slfnEtTPVW5P
s2vikrePySnWE1t6w2Tw634VGETB5CBAMnyJ4UyUr/tCVvobdY2uI5ZFxS/ZJha9
UfMLQtAy+gx5IEKvZ1gibv+F1G/IaBY/FfM1KA4AUQEctW1pwCcgdallgx8dyv66
OE2x1oMN2IwOdLAHMVOtYJh8K9vT1ScY9NPrn/e/MAt2nO5Ex1aJF7EBEp+6sOKb
KU92aUWaToDukRCoaGMbb7ZQ44I2n059r1EgYgKUFQCCNIvDzLr7BDThBIBdZ4MQ
nMS7dfe8VMIL8IpnemE1Sxu9qmax1YSD42m6El9TTOAHgBWKhUNvvHYm16tiFIbB
098VkX5UpAMPuYwfhUMLKJn6KoEhIoKcIsoFAXdX5GA5I3G8a6ig4ws6Edqagh84
FuT1efuu2RTnatbJstWmrhoCpNYufDAUbGzQkkmsHAaLk8THkLjxflHwj8fpgtnj
7avi2dX2ZWpX9vZq2oXqYNzwR8NKywldQBLKVVaNb7t7JN07l84KkyafaYTxaJ97
Y3lNs/y0CvYZkViL0EMY1QH85vuBWnEPkdIurrF4a/3OORidx+i3VKa8aR6EEBwL
u4lLzndyDSO1KuRe4lyA026qWOB2DiIQgnH3Y4Ov9+8IpgBELfXLrEPm6IsZ+gD6
pmQ9/t2uwlg0zOSWOpol/Sy6c/zNKwvUmt7Mb06UrH8ooUVNXMQmHGQh6v63m52U
rShN3gKjqOrYhK6skj/6wJ3OfCcABgarP5S1Z4iD/Lkr7BCXXCx3xcV0PexiAGke
Cbgt5L8wvOtOIhss12I1AjtCREtRnGMsGt1Me7RXYZcJl8mvmyiv5owRINe9RcFR
K3iEI5+zNec3az4ca9OuKJqc5xld3OYHCfGyricUjXorOmjxJSv2RMySAzqpzTmS
mWVWwR3IMPqdo/Vh1Xw9+jwpX21QN10HWU2vLzbX1ci6LMtAmWFrpMScPVHtofVh
p2Nn+JcWFR6M9oJYHlaUo11+hUpzSN2UKkbXe18yJvJNKbKnaNllSR9njpcDNigV
4VI3+mA9q6cPepNqnuCaOn8q/vLS5uFE+jv2XjCOo5xt4qOb29X/QMenWDiFhfQl
ycDUcKLfkdMU3hGxtV57wvMdY0M9cU5kCiHFBemQzLCtoFLaNKrViPheeSYWVu0d
3vFIb870PBydwznBiwtfRQJvPmVpVQBqqaAY4V2mxaRMxyuh+V0CSWl/24dRaVxq
jCPl2ZKCqaXjxt020fK1UO1cYXL8NgpdSmKru6ByWsLyTuaCkJh1O057IbcAl988
bAjLxdqn7K54OVjKZzbg9G+G9S7PB9IkuDgpdqx23hPMZXprtEnqwpJGaKaMqS2h
MoHvxjIbipfM0W3zXraFTQCJPdTR/cuxJEocMWKSv8Ih7IOzGyEjbN4FTVnm3ZK9
3Wq0IWzfGWxckc2wf6QJ92effwdXqRPqC8p0dUiPyoiR1lAUZLCc2EXx9UgyFDnJ
P6KAw7JDekTxvfa56kbpQOIss6m+x2oh7cXZ8mURmdDeanK+50MUeyBrkOdGTIkL
TyiLg1QGBpwRoq+j/RgfLHeTNWD/5Ra0frwF2CfJqbvT8TTxE5KN4WTCVVxXd6vx
kASi2Y03G73d1T58C1TPshHqleIBelnnQoZzPrS+tj99dWckVWVfDZs85LWAG5FN
+5K99L7EuaJkMzWV6zA1FPaBCvZZYfADTqiegi7JOMYgQFh0KwKpLjpkgQEXzGou
J6vVCRqV6vRDXhFo96qjiGuViT36GnQNnXodaQjfBL/dF9rxpUhFQLa64z1PXdaq
9AqH8CEdQ+g71Zsbg//0UkpUewZQsF6c0thC11zLpYR7xNtJYIMGv5oKGoIkwDra
nbxBhif9Z5/3VWq3hPc5Lo5QkktkByDnt9nb1g3yCTO6lu7Ej+EC4DUiUpxsckh+
/xJQpKqu81DxVnlkIrrwcsv/1KX2qMR6lw2TwyYJUF2/V8pq8zzG+knr2qBPwPFk
9aeA9fZ9eCI8KKn0qVqk2uZ3kfx1VZO37UqDOep1QbzUzLcZ5EH9pb8F4T4QQWkY
eN4yeidhQZQg6BcOTnxc+S0tQAqRhxTND7xq3Nk7e4TaJd+xm9UmfSFro3sYNz3O
4a8J9O80KMUKPGyAulePgevVeJTlhYEZzrKAW8amD9oKCFr2u3dXGvLlfGWK6fTU
XWsBA7XfdwjVkhouS/HFjzpeuvvXIYHssAbchO3y+eikXaMz/BgBTy9neMhHnX4e
bV+G93znBAAAbZlNyk4G06J3zWVrkEsR3HdPMhQOI6AOOqFI2c5zr3yJHHTtmlza
epItQmur0oIVTDIsVeiJaHCr6I1b6gynn5KErKGjEjb2blAlge1pBk3hogQy4k26
7WCSL/x8ymx0nWZkK69c1Tx3T2NIJmhijZIzLNJppsdwdiOZU7PRmpaqSvm8zh6T
96seQjhwLQXjtB2L2yMSxO+8FYFXhn0XOQcyyNz+XM2OEXodLyf0CBZn7YblADDY
EYYW9GipnZF1KFySLGJkaFVHPWgvnCRRF6PZuPx2jPDhdc5JH5YndkqeAqlfzaca
Wa+xHdQeIptfoOve8nNgqfTtoyGWRaChseZwLL/RVrcCsnRl6D9qCJkGXDP4Vo5i
nh/Weq9qkEpWjpzJNzjd+u706K16xdDlQ1N1HzVYXzSiuq/nIU9httgpBVPGHpY6
ltEUi8+cdZL0sGFsLgz8hLg38gWDZS/H/8dEtCWchsr1x+POIDKQCV17ZTiAliKT
KHpWFMTC8+ut8o5ijBHB5UdLLKCmUb+jpmQ8u2joe1M106tETe4LLRFIyrDC8JXn
DzC9NOVcxoUDF+Z39pyzzUgP5HJ8b4eHhcauQKxitjz+5Y2bKBq8ADXlmUuiWMwx
fMFANFKdybecVJCnFACLpdFtTGht6AsQiDyZYxJbu55y+Lc5VW6j23AJyVtOn7c9
4cXBoCqnywbrx3rgwrjXJdz27oJymK+H94MEcWpb4f8vFBXl61LOoQmcgZ7Y2O+8
IcBr5XG9w6pamVAWfBxvcWSINKuld+C1/WG0HV16JNtOGtHYYsAktpCNqJ0Fk/E/
lo/YaPUw+ZqtD2PZK4zDgbTOWTYAuooA8k+ykOBLpjP8k0c4W9IlXOMdRWKjN5wo
JXPiDfdvUOB7vDvSHoJwsogyxeEUYIdB8zWbUQx73gTmvN0ZBaM77ojFYdluy5oA
Hn+wYZH5xbEeMqdTVMDrfV4N9F8F1v5A8HSKTKMk3r1GZNqR1KH69YRos/BFwsjT
98iY2eXO1dx4Ze+G110dd+Yoh8q0WSDVGHGbtpO6OUqwFYl0qK/5LqkKuwK3UYZN
GwebIFFre7oS4NPJPzbHLSvMlprooRdmqhUuFzjxCFOtFp3RE2jkbc7y/RituZct
ZhGlazdJdwAcO0RQiILVjU99xTEQV7f1zRAsCVHgUTwVZzowZtNZfrogI3BtUzyM
PV8pasrPwP+vWVUta1zdu2fTcVH6ei6ImrPhZ93siIX1hT/Q6RcZYNvTQDxZp1pg
uDfO9PHr1RlVbTsEt4OSt60frqoyPZWUliww2GZVTTIkPXunwcFTXKdx14A0aek0
xvKPgovaZReRHNnoJi8z7v8QIaPAkD807klFU5fVPwO0pvsd3Uqdx2ij1KW209QV
lHHcmNSzWfrpfWhxtXUifOSDRVGWVev198MTqAwqGDwCZ23RTPYgpluVOwu2HSJN
0kV+Dpo5aRJm3XIXbH+gFQBMmT0a1S1TBlr1OsmA45u5W/IuePGGQY4AumRsTBW8
wXkF44RSOoizJzvMHSxw8UbxDrDxBJk0RYBY17r+RYGRRpYznoU8/cOEkoQ4n4+1
YzdwxuCsGOHZk8MK1NiXgNrvQr4qT3w+26hpJis4Q3VwTMazaudrYlVt3IhWLqxX
2hweF8Qyi9XxfPxEfG3xjYJKgNuD9N7YsfM5j8+lFnbd9phWEL+4x7XjbcGo5Vm6
NZwqbZ435J6Y6//NCmL6I1hB1P0bfoAMKWolW2MjcRYdUoGrByXrUKvRgOd1YC8z
urTSE1IzyLTTar9BVRSeRB/VdvHdKNYGztBzg0Wm9FdFK6yGgQdc407ubqKUMx9U
wQ6AWJ3J5ecCChNfPHRSAFyrkxVaNxgTtlrXpQcUoOlrQ37SBet/JzyGh4eSvIXn
c0wx4d+KdEoYFPV2cxoWhb3RptDTc+2dgiTZEbR2mwgAbrxWPz/gcyNMC1ELmwde
b9Wxkx/xAC644gd2r3E25BW9znM2WrCbCZNFF4MfGxSS22t+3ciXo9RLvhPZBZbi
UL3yo+kqETLZI8NfckvzSlLSAkn8j21EHu+VEyKpHZ30XqHm8IUaSwX2vHUNunMt
0Hj2Bhtp1m5h6T8F9QSzQUemGfE7hW1BHouCgKWpWdDnTFBt6hEoWCAZ6z1EmjxX
0waHwM8AYIPP5RmWcVwlLHRz94PoAWWEtcMWXelIPy6uUTsIFYvs/wpnF2X54cAq
0eQRgcgscRMTme5nH1PHcx7vzw7nb5R6l8z7uORRUgeqesgL2YhDok0rtULmU1Q4
HP/4uqWGnReU4QeGuO+NEdfwJCn633HbHQzKWGaP+asUV4I5Bvh9vj+Q+l5RsdV2
QJqxqpLIjluuW0kpDUOo+VczC8MmqE4O4hn73Ic0wgc1AdWPB84BzTGWzdNJSh8X
rl4n/njYOrNQsEtqB8AO6J/B/9kYUg4eYWmNS3rV6m0Jpm3IVflzexot1gvGHYUP
JnMDs8fAkt9DxZGBpKrH9gykO4Q1AyeTGszzYq8CJr5CgSM1BORoVJ7XbutGZYzM
ZxwLEiH0n1v1NzxrMby3zzEj2zywQLVSvWHg9NUOHsrHBgc35jKdEetN9L+P0coF
CylgE6K24WSqzWkt9CFtCFpjAicepAO6LWcgJ6gO5CI5BLKwmQ9i/scT/oLBk4r6
W9SUvU0nLB31x7OL+Uyuaw5mb1ArHkxqZqrasiGm5ME0t2DwOZImTuqPbr0yrgPx
R5CsRk7PZS5yJrf5mRBXkwcZGdP1hd6ICP9gM2gQLxoPmojR0od+Zdyt+UxVlhMa
6CCx9QNJ6AYFSgIBOLNjK4HdvJPfkbTZusOqbGm9yhlDqaXgYNCvMYcj503okY5+
ifXBq1l2qTThgfzHkQfBSLb4ujlqrhOWAZrE1wEnv9Hbtay8EUeIMlr4IIXfGvXL
WUFdtoMshsB5xmbebb0JMomwDTExJflpiTpmmVUwz6z2/2Wn0QJIeaCIk8lIw3nf
wefna+bDLPcDefj82FRow5xL6mY9QjWpvQNXjjRJ2kEmHym3w0RJgFn7B0+6xIu/
0pDUylHSCju+8mEEH36wCKaceX4bNHFI+0IzxjkyqSllP5Tx9UsOSsa+q48UME2Y
y7Qp68WUu0VrBBzzM8hgtLJW1/rtRoDg5H1m/FLwST6T+jmC/F1SD9gdb0QHh7C6
dC7n1TaEuTmbeSiVZYaENbu3d1Iix/WeUDhEpSzF+WmPiPMk61MwBk2VzUQU7AQV
qTXgI9LmxqgonSdUBNZKxZJtX0EXuHqd3yFzQlaBwSqsHIACeXvT32v6kswc4nM0
ZJ4iRokY1VDO7u8MzQAFRHCkWt4lhxMh4wBw9rD1uwM4MSe1puvyBmyAVtwB57A1
pLBdcM9lDAWIXoEwTRfMW2Wsw47NhlxcG7c4MSQfq8ZFEIVj3DwFFGiG7QFw2FiD
vrU4/2XROBZdMeBxVbfafOU1SwaHvJsngypNKYokUDEoRzjY+05xbTRznqxp/6W+
gcqR6P3AmARFbiJpjDC+6QaJGb9Z6cqyFRivQxVC/KuacmSbQGwRUUGbkZjkNytC
JG4pUup7LrjMEtZqrDb/6uB/2YKwerwAmySd7/4wyswLsguX2LeofzinRrtbLVmS
EutW5tyx335bsQwaEZpOM0JLvVEngcDk9Iic14GPBLpDpDqY9YV3hf0499yFsp2q
Q3wVSWDAh4q/Ap5oxnMs+vMKUf7ZhQRNfBQZ2sODxp9OohVxXwCUiWjcv1Cx0/o+
6XfiLGhdG3yaqp2hpcE9weJyjo+td3lohswlRFaLj2eWn+4dSWoXwSCcn9YKKosY
Ce2zcbpuHGodzmu6Ao7lRj9gpKlHbRlmH4Dw9LVS0kf5iNfh+mqleoGthXIjdcXM
pFdv30WIHEHkkkQ39lPYTe9TZqbRwtwCsJppMDX9xKByYdMjieN4KLI0O/oKLvI9
VRwRF2Tt26rKo0eyg0ZVoNiHegMZpXGG0sUfRbZm3p37cEMdSp0HTAlX180cBMiq
82XqUwzmbVkHXYn8Dd+VQ5pbxvuixvgQocJW8k8HIE93eyLOolwlkpWkPKpFD5Uj
ScO1hZzTLCPYTz6h14+CEjpxyVwV7u2Me9eLS50YXbvScjLDNG3TvGbuYC0WpfMf
6KDf4/Xsw1ZGDuCId2p6DGzrl9DPY/qTP7fepmBj638IHSI3ks/XNsg4MdwgHFgR
NwzK4pKzgynJvr+xLqkrCxcAYT/iaO65Rkne3tpc7A6MyU7Eo78XBn+gO44uS1vz
XGNt0OD8FCekO/Wrsp8KHK+Uib1NGJhZLLOZCpYdwAjiXhUNf8s6oq+6W8gGqv4K
ri7SoNuWnQ4mCUYOpF6RfFE/6KeWCLJlkU8CvqSllk7t3ypi3tdEgn7rU+1pwcz3
LXwfwEQHvBTD1+HnlP4Cem4fTTnmAGSXXz6wrlD65mEPE3MujuG15cHIduzw8J6L
jjV8CBGi5VEfXdKm7BqsiZc1M6PXD3d/8SPKter2O2v1zTijM98YhIc9A4OHL/jw
z+Heyh6LTL6eoGhZKXC6Ydb8uImscAE9qiogj4XzaejcauL3/+dJHyNNzYrRYBg1
F9ahXY+EUmYBu0CO0kc03N2gDWjgnFB6WLuV1Tm7dbj3fMT0/bnYvj2WsiSTjzgu
0uky5GDLk4P+KRKEowBVELPTbE67wcnZnSUo/60JFfkYT/sHMgoDg+bZNrD7GwTA
Ai30fM0SklnzB8r2qmp3RwuvfmMBXPHgK7IcuNpJzqS2zFtpM/rwjF0s1MLqy6BC
OAEGMItCslPWc7eABQuS5QrWR39UnF8RbOMHT9ril/Nnmt+/TvZziT/w3+lgqpP9
5hvpPav3e2IxhyDRiLhHFUCVG5UHSn3HP3xb3saKp9t2CIULw6ogkL/pRYCna9EK
tHkpS89NG07bHnhVSrEJFV1DPS3wMAy4h2lHKL0ytNjb+qtntUKAY+Cy9SfoP6rc
ATvUmDjfDeHYnMD+D1LWSHY/jSpep8Fyie89+ENR2vN8XQM0Bde7w6KQCAmCXRb2
cb9OutprfLyg2FCU2LVTaVTB1n4zb8PqKxvaLoUD2cRMX3hbjXAZoBibH0Xw7aKp
Ek0PgNHmePH2M00z+6gPLoKgIfTk993UcFxtxyvH6mqU/+dZe2zBip3ZPE0FDCKZ
t7S36BmF0h+b056WOGI4HpjdqUukgr+qctkdiijxRYOMIKcLQ5chrwhhv6ANQYC6
PZt+x39Ra5RjBSMrkC/fR4HYRfvV+WJZiVnmEFwIZQXBKqvjCg0/J7b7c22fFV3n
3i4G/JsJNGoCOHC7QwMpH5z109UUHTsFBSrL94WSWzzLcFDnWjByrM1ak0H94DrI
36aVnThAqg2JdqLlk+FfkNHt88I0KcoSdQbIvjgcR97l3ndi5Fgajt2QDbSg+z1I
iHarrwvvcE69QmxxhxTdDebL4mmNYvgXdhNgn9DGIN53UjFnA4iju44qcGFN1wvh
3dm5l/x3JqZv6ZaG7Y2BAXLXwSydphy7x6UU7Fz9pWxkyq3UwWrWp+9xD8EY5LRL
+BG1FAPvdg6LkdrIIX2HFy5Pkpz1SB4ILe3E4aTPIOYI6vBEGcLpZCNagC+aXI8d
f3jBiVUJWLnZgQVzuipseiDlhRj6JJKBV51CgG9Hwq6p1vL+k7RqUOFOgan2drf1
7Z+ajNaeY2MH2LlL3po79WzbShKI4wAASueDSrhHPgUaEgJOwVYrYaJLR95AqCxL
t48K28Wf9Ezvw23R11pIjkd56kKCInB8lPamn8nABFjhILjuIyYJP1bvMo/zQJpl
Qd4kk3VUtGff+WvS3gJQnSaqzuXiUP9Q7oyDeZps4fUP18VWcVqLc9XWgBgd9HYA
Uau7sZRBDffzc/fQzWoLYdTjXGrJMzHrCUDrPzAZjcAuwzc7AK7puArXhmKbK7zE
9DmmrjpeYDXXvb85CKWJEeG/mwDarW4qMeYPFxXnWwujG1tsjGkfPGQGG85KVXSM
hFT1aT6llLf1UZFxRXRg9PE/tdIb/lguW57iP3P3FJZmfojWJtKxI8y1DOZBG4oS
aROrPYNlYDArKUdL1N8qLMESFS0rgq7cGjJN6/7DjIoVNpPpqizcwuSDR8xkGGRX
imfDBVY1RqzkFUDoZGkCUuTUuii4vC1sdliTlI4SaLD741idR/U8A5IXDQN2R96U
n4vWoSAZApAPLZ3icDwi14otOTOVPOl+CUVyV5MXJbcY9yvwKI8G6vtrZM1d4om1
kiYWRmoOB7fESEKnOoBlrKmKqh5pYw9g7kt50FPZGNO3mUHKJiPz2aj/VG10y956
7tVtCmSXNiwxz8Ic++e/H8uxtDKYCHVU1sTbfMvU+6RBq1W+kLDLSBHyN1nVoxas
DKHeR6PilNl5/U0Kfp+arf53D9ZxjbrwpXZYl3ZWsK5/KU5pBgN3j0DHglrsFwdS
jFRwdxCI1KkhQTzCoD8hVcwSvecwuHRxdjQoJSYI2bHxQ2fLt46gTCNEkgQNzeNg
TF2HsEV+vQba8gv6uOktBGYHH1fN0DAQVincNt7NplI2iiGjWBws05hkM4Bf7IY3
b6wfCRmVUUkyk/9Tu0Kol25OyiwPooQTwJUel/SFcS4KpiHW1U+Z4xKbxgQG+BWX
h0ILEtrtQy7vz9RWbdjvAdWR9jVSASHDSRFaOyvCiHNhI7BdG76K0ToUgEA6yoKl
wNppwn77Uf8eL8KKVSqPsULUEIM2O4A5wpGGTwtJfOiLP6Vjmqna4Q0kCGenwr4l
06qtnXrvA0Sfa4Cugh2MlQl6brzpgce5Ynr36mlWLs38DG1bj7BypuSUQHka3sAH
0RZHKMYGd4H31ZwGepdZcPDDMz6fG8MKMYax+uMsz0440rYG79aZqoUC8MI9kRuc
81Fgn51wlFg28XgJFbJFsY7mFTfH465nVE2Zu+rvk9jKpNsuHgDK/Vn5cF4nJHrV
MIF4nKmGr7i2hbUJo7PlDu1NPWEPKdCKaJZNmaVc9wZGWDYCfAH0cDZim9S7Gujc
`pragma protect end_protected
