
module mgt_atxpll_rst (
	clock,
	pll_powerdown,
	reset);	

	input		clock;
	output	[0:0]	pll_powerdown;
	input		reset;
endmodule
