library ieee;
use ieee.std_logic_1164.all;
--use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;
--! xilinx packages
library unisim;
use unisim.vcomponents.all;
--! system packages
use work.system_package.all;
use work.ipbus.all;
use work.wb_package.all;
use work.gbt_package.all;
use work.gtx_package.all;
use work.sram_package.all;
use work.fmc_package.all;
use work.system_pcie_package.all;
--! user packages
use work.user_package.all;
use work.user_sys_pcie_constans_package.all;

entity user_logic is
port
(
	--================================--
	-- USER MGT REFCLKs
	--================================--
   -- BANK_112(Q0):  
   clk125_1_p	                        : in	  std_logic;  		    
   clk125_1_n	                        : in	  std_logic;  		  
   cdce_out0_p	                        : in	  std_logic;  		  
   cdce_out0_n	                        : in	  std_logic; 		  
   -- BANK_113(Q1):                 
   fmc2_clk0_m2c_xpoint2_p	            : in	  std_logic;
   fmc2_clk0_m2c_xpoint2_n	            : in	  std_logic;
   cdce_out1_p	                        : in	  std_logic;       
   cdce_out1_n	                        : in	  std_logic;         
   -- BANK_114(Q2):                 
   pcie_clk_p	                        : in	  std_logic; 			  
   pcie_clk_n	                        : in	  std_logic;			  
   cdce_out2_p  	                     : in	  std_logic;			  
   cdce_out2_n  	                     : in	  std_logic;			  
   -- BANK_115(Q3):                 
   clk125_2_i                          : in	  std_logic;		      
   clk125_2_bufg_i                     : in	  std_logic;       
   fmc1_gbtclk1_m2c_p	               : in	  std_logic;     
   fmc1_gbtclk1_m2c_n	               : in	  std_logic;     
   -- BANK_116(Q4):                 
   fmc1_gbtclk0_m2c_p	               : in	  std_logic;	  
   fmc1_gbtclk0_m2c_n	               : in	  std_logic;	  
   cdce_out3_p	                        : in	  std_logic;		  
   cdce_out3_n	                        : in	  std_logic;		    
   --================================--
	-- USER FABRIC CLOCKS
	--================================--
	xpoint1_clk1_i                      : in	  std_logic;	      
   xpoint1_clk3_p	                     : in	  std_logic;		   
   xpoint1_clk3_n	                     : in	  std_logic;		   
   ------------------------------------  
   cdce_out4_p                         : in	  std_logic;                
   cdce_out4_n                         : in	  std_logic;              
   ------------------------------------
   amc_tclkb_o					            : out	  std_logic;
   ------------------------------------      
   fmc1_clk0_m2c_xpoint2_p	            : in	  std_logic;
   fmc1_clk0_m2c_xpoint2_n	            : in	  std_logic;
   fmc1_clk1_m2c_p		               : in	  std_logic;	
   fmc1_clk1_m2c_n		               : in	  std_logic;	
   fmc1_clk2_bidir_p		               : in	  std_logic;	
   fmc1_clk2_bidir_n		               : in	  std_logic;	
   fmc1_clk3_bidir_p		               : in	  std_logic;	
   fmc1_clk3_bidir_n		               : in	  std_logic;	
   ------------------------------------
   fmc2_clk1_m2c_p	                  : in	  std_logic;		
   fmc2_clk1_m2c_n	                  : in	  std_logic;		
	--================================--
	-- GBT PHASE MONITORING MGT REFCLK
	--================================--
   cdce_out0_gtxe1_o                   : out   std_logic;  		  
   cdce_out3_gtxe1_o                   : out   std_logic;  
	--================================--
	-- AMC PORTS
	--================================--
   amc_port_tx_p				            : out	  std_logic_vector(1 to 15);
	amc_port_tx_n				            : out	  std_logic_vector(1 to 15);
	amc_port_rx_p				            : in	  std_logic_vector(1 to 15);
	amc_port_rx_n				            : in	  std_logic_vector(1 to 15);
	------------------------------------
	amc_port_tx_out			            : out	  std_logic_vector(17 to 20);	
	amc_port_tx_in				            : in	  std_logic_vector(17 to 20);		
	amc_port_tx_de				            : out	  std_logic_vector(17 to 20);	
	amc_port_rx_out			            : out	  std_logic_vector(17 to 20);	
	amc_port_rx_in				            : in	  std_logic_vector(17 to 20);	
	amc_port_rx_de				            : out	  std_logic_vector(17 to 20);	
	--================================--
	-- SFP QUAD
	--================================--
	sfp_tx_p						            : out	  std_logic_vector(1 to 4);
	sfp_tx_n						            : out	  std_logic_vector(1 to 4);
	sfp_rx_p						            : in	  std_logic_vector(1 to 4);
	sfp_rx_n						            : in	  std_logic_vector(1 to 4);
	sfp_mod_abs					            : in	  std_logic_vector(1 to 4);		
	sfp_rxlos					            : in	  std_logic_vector(1 to 4);		
	sfp_txfault					            : in	  std_logic_vector(1 to 4);				
	--================================--
	-- FMC1
	--================================--
	fmc1_tx_p					            : out	  std_logic_vector(1 to 4);
	fmc1_tx_n                           : out	  std_logic_vector(1 to 4);
	fmc1_rx_p                           : in	  std_logic_vector(1 to 4);
	fmc1_rx_n                           : in	  std_logic_vector(1 to 4);
	------------------------------------
	fmc1_io_pin					            : inout fmc_io_pin_type;
	------------------------------------
	fmc1_clk_c2m_p				            : out	  std_logic_vector(0 to 1);
	fmc1_clk_c2m_n				            : out	  std_logic_vector(0 to 1);
	fmc1_present_l				            : in	  std_logic;
	--================================--
	-- FMC2
	--================================--
	fmc2_io_pin					            : inout fmc_io_pin_type;
	------------------------------------
	fmc2_clk_c2m_p				            : out	  std_logic_vector(0 to 1);
	fmc2_clk_c2m_n				            : out	  std_logic_vector(0 to 1);
	fmc2_present_l				            : in	  std_logic;
   --================================--      
	-- SYSTEM GBE   
	--================================--      
   sys_eth_amc_p1_tx_p		            : in	  std_logic;	
   sys_eth_amc_p1_tx_n		            : in	  std_logic;	
   sys_eth_amc_p1_rx_p		            : out	  std_logic;	
   sys_eth_amc_p1_rx_n		            : out	  std_logic;	
	------------------------------------
	user_mac_syncacqstatus_i            : in	  std_logic_vector(0 to 3);
	user_mac_serdes_locked_i            : in	  std_logic_vector(0 to 3);
	--================================--   										
	-- SYSTEM PCIe				   												
	--================================--   
   sys_pcie_mgt_refclk_o	            : out	  std_logic;	  
   user_sys_pcie_dma_clk_i             : in	  std_logic;	  
   ------------------------------------
	sys_pcie_amc_tx_p		               : in	  std_logic_vector(0 to 3);    
   sys_pcie_amc_tx_n		               : in	  std_logic_vector(0 to 3);    
   sys_pcie_amc_rx_p		               : out	  std_logic_vector(0 to 3);    
   sys_pcie_amc_rx_n		               : out	  std_logic_vector(0 to 3);    
   ------------------------------------
	user_sys_pcie_slv_o	               : out   R_slv_to_ezdma2;									   	
	user_sys_pcie_slv_i	               : in    R_slv_from_ezdma2; 	   						    
	user_sys_pcie_dma_o                 : out   R_userDma_to_ezdma2_array  (1 to 7);		   					
	user_sys_pcie_dma_i                 : in 	  R_userDma_from_ezdma2_array(1 to 7);		   	
	user_sys_pcie_int_o 	               : out   R_int_to_ezdma2;									   	
	user_sys_pcie_int_i 	               : in    R_int_from_ezdma2; 								    
	user_sys_pcie_cfg_i 	               : in	  R_cfg_from_ezdma2; 								   	
	--================================--
	-- SRAMs
	--================================--
	user_sram_control_o		            : out	  userSramControlR_array(1 to 2);
	user_sram_addr_o			            : out	  array_2x21bit;
	user_sram_wdata_o			            : out	  array_2x36bit;
	user_sram_rdata_i			            : in 	  array_2x36bit;
	--================================--               
	-- CLK CIRCUITRY              
	--================================--    
   fpga_clkout_o	  			            : out	  std_logic;	
   ------------------------------------
   sec_clk_o		                     : out	  std_logic;	
	------------------------------------
	user_cdce_locked_i			         : in	  std_logic;
	user_cdce_sel_o			            : out	  std_logic;
	user_cdce_sync_o			            : out	  std_logic;
	--================================--  
	-- USER BUS  
	--================================--       
	wb_miso_o				               : out	  wb_miso_bus_array(0 to number_of_wb_slaves-1);
	wb_mosi_i				               : in 	  wb_mosi_bus_array(0 to number_of_wb_slaves-1);
	------------------------------------
	ipb_clk_i				               : in 	  std_logic;
	ipb_miso_o			                  : out	  ipb_rbus_array(0 to number_of_ipb_slaves-1);
	ipb_mosi_i			                  : in 	  ipb_wbus_array(0 to number_of_ipb_slaves-1);   
   --================================--
	-- VARIOUS
	--================================--
   reset_i						            : in	  std_logic;	 
   ------------------------------------   
   sn			                           : in    std_logic_vector(7 downto 0);	   
   ------------------------------------   
   mac_addr_o 					            : out   std_logic_vector(47 downto 0);
   ip_addr_o					            : out   std_logic_vector(31 downto 0);
   ------------------------------------	
   user_v6_led_o                       : out	  std_logic_vector(1 to 2)
);                         	
end user_logic;
							
architecture user_logic_arch of user_logic is


   --##############################################################--
   --## Uncomment the following signal for PCIe extended fatpipe ##--
   --##############################################################--
   
-- signal clk125_1                  : out std_logic;


   --@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@--
   --@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@--
   --@@@@@@@@ PLACE YOUR DECLARATIONS BELOW THIS COMMENT @@@@@@@@@--
   --@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@--
   --@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@--


--	signal regs_from_ipb_regs	      : array_32x32bit;
--	signal regs_to_ipb_regs		      : array_32x32bit;
      
	signal regs_from_wb_regs	      : array_32x32bit;
	signal regs_to_wb_regs		      : array_32x32bit;


--@@@@@@@@@@@@@@@@@@@@@@--   
--@@@@@@@@@@@@@@@@@@@@@@--   
--@@@@@@@@@@@@@@@@@@@@@@--
begin-- ARCHITECTURE
--@@@@@@@@@@@@@@@@@@@@@@--                              
--@@@@@@@@@@@@@@@@@@@@@@--
--@@@@@@@@@@@@@@@@@@@@@@--


   --#############################--
   --## GLIB IP & MAC ADDRESSES ##--
   --#############################--

   ip_addr_o				       <= x"c0a8006f";      -- 192.168.0.111
   mac_addr_o 				       <= x"080030F10000";  -- 08:00:30:F1:00:00 


   --#############################################################--
   --#############################################################--
   --############### PCIe SERIAL LANES CONNECTION ################--
   --#############################################################--
   --#############################################################--

   --##########################--
   --## SYSTEM PCIe FAT PIPE ##--
   --##########################--

   sys_pcie_mgt_refclk_o      <= clk125_2_i;

   amc_port_tx_p(4 to 7)      <= sys_pcie_amc_tx_p;	      
   amc_port_tx_n(4 to 7)      <= sys_pcie_amc_tx_n;	
   sys_pcie_amc_rx_p	         <= amc_port_rx_p(4 to 7);
   sys_pcie_amc_rx_n	         <= amc_port_rx_n(4 to 7);


   --###################################--
   --## SYSTEM PCIe EXTENDED FAT PIPE ##--
   --###################################--

   --(Uncomment CLK125_1 in user_sys_pcie_mgt_refclk.ucf)

----=============================--
--	clk125_1_ibufds_gtxe1: ibufds_gtxe1 
----=============================--
--	port map ( i => clk125_1_p, ib => clk125_1_n, ceb => '0', o => clk125_1);
----=============================--

-- sys_pcie_mgt_refclk_o      <= clk125_1;

-- amc_port_tx_p(8 to 11)     <= sys_pcie_amc_tx_p;	      
-- amc_port_tx_n(8 to 11)     <= sys_pcie_amc_tx_n;	
-- sys_pcie_amc_rx_p	         <= amc_port_rx_p(8 to 11);
-- sys_pcie_amc_rx_n	         <= amc_port_rx_n(8 to 11);


   --@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@--
   --@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@--
   --@@@@@@@@@@@@ PLACE YOUR LOGIC BELOW THIS COMMENT @@@@@@@@@@@@--
   --@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@--
   --@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@--


   --------------------------------------------------------------------------	
   --------------------------------------------------------------------------
   -- The system ipbus fabric and/or the user ipbus/wishbone fabric can be --
   -- accessed by pcie through the ezdma2_ipbus_int module implemented in  --
   -- system (BAR0/BAR1 and DMA0 are used by this module).                 --
   --                                                                      --
   -- Note that the address in the pcie part does not match with the       --
   -- address in the ipbus/wishbone part. The purpose of this mismatch     --
   -- is to save pcie memory space.                                        --
   -- The addrEnc module of the ezdma2_ipbbus_int is in charge of this     --
   -- address conversion.                                                  --
   --------------------------------------------------------------------------
   --------------------------------------------------------------------------


-- --------------------------------------------------------------------------
-- -- This bank of registers (ipbus) can be accessed by ethernet of by pcie. 
-- --------------------------------------------------------------------------
--	ipb_regs: entity work.ipb_user_regs
--	port map
--	(
--		clk 					=> ipb_clk_i,
--		reset 				=> reset,
--		---------------	
--		ipbus_in 			=> ipb_mosi_i(user_ipb_regs),
--		ipbus_out 			=> ipb_miso_o(user_ipb_regs),
--		---------------	
--		regs_o 				=> regs_from_ipb_regs,
--		regs_i 				=> regs_to_ipb_regs
--	);
--
--	regs_to_ipb_regs(1) 	<= x"acafe01a";
--	regs_to_ipb_regs(2) 	<= x"acafe02a";
--	regs_to_ipb_regs(3) 	<= x"acafe03a";
--	regs_to_ipb_regs(15) <= regs_from_ipb_regs(16);
-- ----------------------------------------------


-----------------------------------------------------------------------------
-- This bank of registers (wishbone) can be accessed by ethernet of by pcie.
-----------------------------------------------------------------------------
wb_regs: entity work.wb_user_regs
port map
(
	wb_mosi				=> wb_mosi_i(user_wb_regs),
	wb_miso				=> wb_miso_o(user_wb_regs),
	---------------	
	regs_o				=> regs_from_wb_regs,
	regs_i				=> regs_to_wb_regs
);

regs_to_wb_regs(0) 	<= x"00112233";
regs_to_wb_regs(1) 	<= x"44556677";
regs_to_wb_regs(2) 	<= x"8899aabb";
regs_to_wb_regs(3) 	<= x"ccddeeff";   
regs_to_wb_regs(15) 	<= regs_from_wb_regs(16);
--------------------------------------------


------------------------------------------------
-- User pcie slave, dma and interruptions demo.
------------------------------------------------
pcie_demo: entity work.pcie_ezdma2_ref_design_wrapper
port map
(
	reset_i 				=> reset_i,
	pcie_clk_i 			=> user_sys_pcie_dma_clk_i,	
	---------------
	pcie_slv_o 			=> user_sys_pcie_slv_o,
	pcie_slv_i 			=> user_sys_pcie_slv_i,
	---------------
	pcie_dma_o 			=> user_sys_pcie_dma_o(DMA1 to DMA3),
	pcie_dma_i 			=> user_sys_pcie_dma_i(DMA1 to DMA3),
	---------------
	pcie_interrupt_o 	=> user_sys_pcie_int_o,
	pcie_interrupt_i 	=> user_sys_pcie_int_i,
	---------------
	pcie_cfg_i 			=> user_sys_pcie_cfg_i 				
);
--------------------------------------------


end user_logic_arch;