// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:05:38 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
BVsxdK9VGBpJFY3q0D7WVXUGK4C8VRxWgUcNtgjUa1aTvnLjhdCqyKFo0R44GIVr
FJ2XzW4kWux8Wl1BO6ysvfhxACn0JbcWtNdNvmdCCETtg7k1eI9ch9oZZ1GrP/Bx
I2LmD7aSRFtdJ4U7Gj6f9VhvlpiQ1UtedzoNnBnqmvc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 25664)
ph0NPKpTBRBexAfUDZMzATpIUweD8Tv3TQ0MXbNkqsmyxJLOHobqRbZhjFD0+aZS
N7ip5eQ+1PdR5iih9xqbvrtoi3QK/G7UqiRz50LV9JRlo8CyisTjBP+GnLDZUiJH
cZiL7fsTKgOvjBChMclwCXrO5KcDbLsqV50l9+XJqDDrOFz3hgBy4550DMgBPA0z
jod+qaW/X45SK4tidryF0N6sPg7lrTJzk2pG5H2yOnbysqGZcbuenb+Z/WNkaMJb
AW7CzAWRrPHe4A0rK+56zYiLUHQMH+rM+uu+gA8Mb86zFFken/z1QPCQcmCtyd4U
cvXWwVg44qSTshooKLfKsGGGtJPitUpMoWu00aKRXgGQcC2Y+YoL7/mZqRlmYeBT
7sLAxkL+qw/NY57CQy3CZkym6ojC5VLKaXdKb+glGr1d1gqd1/2an+XiaUzuvFDe
L937sz3ifg4AxRyETm3pjczsLOMkQZ0rGgTDBIY8yOx7k0JkxsTTIf89mIjN7MUo
+S8dTCo6T5h29+BaKOm2iYI4eOPVSdJKjDXIU11fu7h/9XJD1Fsy7T0vGZTrMLqI
FSe3ofDAiOPAW8exo6CymtGn4pB6wkGjURUcAA6tIbVSaIUvOEiN8PiBd8d35XGM
vM2guXE1KsTY2oHRHSiAn64AU6seF1W2MT+EWHOz7RG+L6VJTAPS8IiOpZ4CTO/Q
h5MXF0lnxiZrCXqBWmOA26UpoWmzlVcd8JpcsTLzUlFV+d9Jo23yZ0ucPOvQixMB
VRHwGdr0/b1/rZJgDOwlqSO9jUDrPQ6pexX6AZXIdY9X5DYkQkQtBqIdX8KifDtS
Ycx6kxwIJh3MSxnbEFOsGat4CvWyT2ZPh6jmLqgJdDjG93KzfRL06qqgijTad/6O
M79Mk1HMb8k2Nn4LvFnME1PGIDIGAXoovlJrJTUBr9aL0TKFwxOIxI0XIUISGZyP
KelvMWHYCOb2aXrZ1DrzN2Q/CbCfqiA2L9fKEWb/3Df+kKGuxp3mzrJ9yEmA5s2I
pd3eSpyKxDBrOXaV5jJAGti0FOE0jOti9BSd3nyATybRUGTUtkaFo1BO5NuxprNf
hn75A5lawV9APWuyBOzz8J8P5s+ymuqja4fTgOJmc3O3IQPCAfu0pwxflcRulgWO
C1VV/7Nk78bYlfzOs3hmfT8a5SECo//vdLInySCwc7GROR+piPjISTwCi+08gAMa
CLmk+1cnqxPkLijZ909PFibWEU+VtuineYG1huLFoZ9XhYl9+Io0Y40pxaafWh10
GbqvUy+OLTg/o2WRxci9a8AriiAtxNoRKDFY0Bti0BnjrrpD2DH0N1Rc7b5cdkCv
zP8HIo1Bga6Dw4mzLJCC0IMhNZtaGQTBW0m70PNViYrAS4QSsxv37PIGtDYvoha3
WX2GxJAn9TtABb/APLBr6QSfSxSXB3S7DoD7FaI0a8mHyU0Na0HrrnXhmZVjOIX8
7DTFXvLEqnOEFuD/rlw8SA/zVMCNsdbz/z1Q2n0e3yjEFNu02FvXxU80de5sy8D9
fSnu1OfIogCrbhmpdLdzYGT5igNCmmPYQVZf+2D3VuOYRuaHjFBHd071WAsw6JX4
91Wg5Z9BJN5Uz84mHYIgyzO4g5XBI3Ftx7pUmxj39KXcEaqccQ1DKBcCQemYidui
A973oFUYb9kmDhWUx2hZJXFrA4Wyi9TovOfKEnEw5C1i3FWg/KubkVFMWk2pghqW
HG5XcoXH0ETSZa+ZFkMKPooz5xFjtMfYL5Vc7SUqFG5iQ7CjNYRfU7mLqVGoJYP2
cOB1pvrBuop9PR6n/5leZ/y/eDCjr6NWNHsLCjCMmwPZQdMgY+7MdySs3Uqv7kr4
+nodVayiEN93uVC/LVIvuc15ywAbD+X9bqm/YUquQ2QnAI90b5XKKQI/Gjakx6gh
6Aaq5wMhcmZGSHAcQaQ3QHQNLJDIAZqk96A+Bji0fcyQgOitYN6SnYwZ+6x5G9yY
3rSW3COEVWpkK5dAIkWj7HgHNTRdVUUXioOswkgOmAG+b83ueCHPWxpNtYq0Z6gR
/yrfQtFgIOAxaqP1uV0Bp+C+E6bpJT43NMWaYHQ2zsXd95w4s0lRup8ayiV5yfKA
smBthfdsmrUFmUcdmftadR6SV4rpSsutjeXtGyRoW0W7bUKASa5JDmVQ7YQ93RQT
vxaTAPWG+ylduZKqerXGsnXzNFlTANTkHsL6dUEiEOLRVyaQrnKS2u6oGWbq1n0u
VGMhhLb3jD+klJcGHpeuvU0h3Z/Oci9cKO8BmPV+q2+DjmqIyMuSh+ww35QJrUlx
k46XD9RziGmUZKMMsoP887ixAf9EM3ERFNwdWDIc5u8uNOIo+Dp/sxVMnIidxm6Q
jQiA3sxDIpHkhx6L7dxSEQLjIiHx7Y5S2Sv/hsOAgR19526ODPRCatTQ/VYgA12o
eJ31pM4YPU6iA27ydQZ0MFEhPBgCTvbzVeAAuc8JDGk+Nn7sivAKr+TRjOT34hTU
gcjoWjdtNLoL0x5aBufD5WWUMvYu5UKyhZkmUPxDNAWOVwhqhXTAt8Hms57Jw0ns
Ea+d395q/4oOy4ta6Ap5kbtTZ9xq0uV81m/u82HmF/fwHjizx4Ru/Jyupq4q4mvh
KRmZER25ITK0zd3hTIXiGIylr+MicP2loE2Ed8ODQwJGz9EXtTrX2Z39FCZaqYE3
B7g34eHJeQafD0rxm4b4WV0UXaBO1MwMtG7niXospEsG7Ph7QY3cMJ7SCaLorNiI
C9QZVgosWuLPfSQUtNDOQ6Dz4ggxb6ywmaiA5cfUlYBd6Ne3/p7ppn1dw7EAO3D6
yEXC+JQTsiivdU+TYluCzFfJyOEgomBR6F+64hueOd6mLfbRVsVEvKZxcX2xaflt
7QMGWldFsc/wujqxhUK68ZNoFjicBdXPi/nlgFcx8DqdZrbVcYKlj4wl4YrIXDQ1
mHb3E8nDtEmNjk7OTRmjYP5mOpPhneDECR6++hN61xwZYeZttclxYdI1OjcxkcJO
DSZ6SHWH241HEykYNuGZdNt16yuSBJwNUM+6by1YyDQEsEl0uxRIeRFqEcuPhY+R
ot9qOQZNPk+nkfdvmiXOcs4MILOji/M3vjIYbJpIBoi5p6gSZ+6QjXq08LN2LCvt
ADMZwKk52FbfG+t7zRtLHIdRxisbbS+DfULHYUwGot1FiXsGE5jPEnOJasngy1aq
WjhyIbGXq1Ds7OHvu3JPxcY9McPm7EZeoGdsahGRpxrjpy5tVY69UgCrKNWyycQK
YLYtP7nuHRKDteTP2Ao23PO+ph3BVYS+U5oq4npvB4VgWfaDhGwVzwdO4YgzY4cQ
oNwPTbY/VgShhwJrMAO4j9dK+VhdFdrZN9XtX4ukCHi5ZdMG9+hHwdgd+aOTV/qv
3qbdC/ruQyFDLQ0zNwZ02/y/oQ312vdCHywSsZFjbxn52iW/h5FSJeNyxBTbKWpz
jCT/4jcDL7PuthkMNJ52vRb43UgjK9jzNCZXd9UHpBuXzcuUFfs3K0xGeWNIYuKW
7gckXYemkL9XnEaxouLjd9hcnSXg7doDbHNNZ7TpAO6kNX2yxrjX6sgLSW7eUqWM
+HHqTh3GSjB6ae9df6WCitN8X2bPTak4I6tZopqzUlVBeJnBjuuco3Ow3Yamil3q
g0m2OjCozz5mXVPa42E2QbeBuqbS6MyhhSqjdfOO7REIE2QfUqZXrcgDmqEmVN/R
053hk3/NfW7euRO1qo8wTqrwRc60cAfUXB3SdhUTAezbY/KVmV9igW+pjzThosz7
4Zca6RyIdtvxtiU6hjLgzWBGjmgbsLt+vmJBEY21Firyjk5CxuTatsUz0DXLL8Av
iI99ErS+X7Fk9fvd5zkue5d58F9arsQdxe59s4S+GR7WHLU720mbMxmZGs4ub/0C
mvAKluoHcosN7avSmG+x1FOCS+THb4tl8917aL/wffk9nJnQVEkaElfy3PFygZWm
aZGylZcKcDe5yVtWpo7qhJLgCaAKOdQW0yrug4fmyD2DUalpNTVKipqYgEvMtl1f
/iDrmWtBTfMT2otGo0PToaBBQ9yW/+XjxNHl5bpLyRp/VLdtq5z0r49vk1MUmVlR
ZrkSXyKt1E52UiOsYIxvdPJSW5NF9UHAHVaLzfeqyvnQ0FUIkFILxIQbIHGNl77A
YjccZGxCV6L/hqul+1CdPLbsBRpkL7fakQrtMSo+pjxlSVZOiYRIGeNUC+Ehq4IZ
AuxDQ9CztzoZi5/+TrHj2K3el0gAPdAbCV5dK6AU4we2i+zFGR+sqtb5h6bb8UQb
ePgNtn7BJ/q6C9ZvZtcTYKEDVp0l35J6oUoJsTWBM/u+B57rtqxdmq4YQ0vJGyZc
kjn85jsFKkYRvJWkNuSMBe1aeD/z/JMcIqZx1Ebqcjt3dy/PyNjabJUzf5h6h1Lf
vkNB3m3GDdTUkVzNNjG6mrqMKMMwM2DJtfhj/AAWtwNFkwWs2caLhb6UPHiVv+gE
1gVFX38FnFKLbyEsPUGytdotaBxy9c3mcWBUEGJzHFPI+JYmyhrHAY6hU2mTJcyH
T+Q4fV3P6s7yvwdxPR0bQ7bEHTE9uC6pUYEEMxBfXw7FweXkr1s8Puc/nAicIueQ
uZul/qm50xUj8GmrAfAECAokS+aca7a1M76630H34gzfJMu5FBMWnF01DlfH/F5Y
490VL3U59aYfQDbvFnQJGxWb02D97LHilxeQNNC0pppJpdKiz/d6qVLvSF4eEp5B
W9Q29KPQy98Lb9NiLhZqyLC/N047lKOVzM6UQ9I9W68Tq6lC1rDWSdN7rp2r7DcZ
pF4f6H0e82D6w/c1zpQYrWM18a/8RP1t240f5zqZYnGFoRd6VawZPJNiZSMW2+E5
wH+xVphtcwaTsnc4JzYVvd15hiSNajt2f66S6EXuesnjV+o3nbfMO8+3COmFNO48
HEpL3clapRG5OcM8nlLhPVAzOY0TpA/fEWcsmcGXOjNrPR+ydrgsmyeTIPKIy+Kx
yvU8gzPXdjpBCjOL+VPPHCgLcdB4GppP7sIl56UkDNrDrBZGwqzVSHLE60do/Fpp
MEyJPrayPtkUYNOWd3clfJWR3uBWI7GUnq9gCNz0Kcv77okkONMthAlFY+gdRdo8
KBiYf2wHaGE9h9MPNTpAsnkSZgh1ZRJNj3pRK2cJE5lKS0ARamwa2wyOJLXt7ONZ
fUNK4+ZlNBW1fH1AqzQC8b+i1ZeqjXJmqjtbyw7hGfRIgAIScPZB156cYJLh0sZN
OrPkwePvZuFGBzUIIUWpFM+3LDzBF4+PYNfiffNvHZatTAhs+NbWJx8ix367Jmtm
0pzbAcnPfeFft1341fT13BQa+aJwJ4O5TbP0CZmF4j7VITKZVFLZeABA4SmqVIrC
HF4Rxhz7gQtC4JdPBV+npTHfeHjDJlBwtMzv0qL4k+Ri21SCyEAP8R181dLhU3nT
/MiPK0tknmGP6F7WXX/NksU5G3VjYYBqVZTfrAvkP6s58FuxNxphCTJQxrnjub99
FGwmjcgVbXWVVdt3JHAMu7NzJERsMrkVS1BwRfTHC2sSVTTbVqNV+qEILTiH3sdf
XRP6DxFffERq+0L9coGfMeyZJaETV4D2skkf6UHKrFYSMGrnLdO6FIog7AMUMJUQ
L9BWUZffnj4CctFHIhL+jlv9Asq4+eZ1IhxHCpOidR6ozZYEA533kdcjPpfWj5bO
eAp5mKrfRcpsBr1Ck+oOGWSsHQyM+9EcaKp6+V6clJx3+XT7nAKup1pcNPGadhZh
TqHx9qKMbVNRC29OFM/YE95TIjql7LwWXcLi9X+tLmdw5cUuxvEx8uEV/0qaaj9p
i4Sp+1l6yLnXP3Jt0D5DPlzKQPVfuW1UlEAI5ECBK5x6BKYyUDNJd9Z6pcd36aux
ftBDzW91H1p9GgqRbZucogdNuQCD48ROi3h4Lbo5hdZVQxvPdh2QLaaIDHLDeUv/
x/ZJAVoL/LlzZY/BzDwj9QtVdRy6Agybp1injsPnGtbIBmo/cLEfh8tXga2UWqC9
HnMagDIMKe5plO58VsRrId8VidbbJCS7g11OvRoCt3MBByWyUsS6/HIOCfV838i0
76wwPp77ArDFs8/WJD6vjlBMYWjUxBqy1NZqhE5gRCNh0NDle9x//7oEacTnJsR3
wa32iJIllfsrmUk7hM/w8sTonnB8aXbPSmhmK2Yr4QK+EPmnqLArZt4hvnXgiVU7
2tylwdWIyRDEDqK7NNganRKtbFTKUA4ZRvldHNjh4NiTcQJ9C5QJ+7b9JD8Vp4KL
YU7nbMnBsHOUJ1wQgyzNVe2tSnFBDL4TZ92SGzNwKa2bcsb0yuYAuYI8BtNcp8Mp
SQEsqpWV7w/ZNY3UW/EWuxTwrW48fyof05LRI8Eg5VuBE+dRceJQeXhcLXHoDlkB
O3y+WDkS+827ecflY+Z9pLdm1co+Z/9QvfhBtSZvmRirQBOW2hlxFrtTicYtht/0
EjgfuSHStD7VO5Diz2sh7f/ps6477MA3dVpf/DEnWUIi84lEnqnj/fai9IJUxhgS
PbZljWeXHBIUQmr9p0DVsgT9s7LyCYvlGh08EyteRKxTMoG6SNbdInhpg0W4eo+h
tHgXhGMoxOjUrUTKLcKH9lyglG7Y7I+RWWwJ8kxhu4MTeBFYfupwPLe3RuMsb6Zh
Ir2WP5COrWHvhbLxeqH/i/0R3jpSd7jLOpOjUN6pGxsl9P5tgMQrdOlV9k0FTkm3
s3OeCQ7xq92GzsYmN82SGwamFGpbcKthbvR/otBT/+fkiWKmItJB855FT6D0HSUg
/U5pGNil6QWB53b1/sV1o6bUl5aXIdWjkQGwDmtsZrcWpUd3NSH7943V623fpzkv
KLtZekNIQ/O8xzNbmrzZUqLpBZEIPPYflg9R8L+wJhb40s7gph/mIIRu4fp3vs56
sEdgLjF0WCzbr/LLwxxupXWbGL3hwm36gizSFUnnCBJu4RMNLxzUPo9CTqwjb4lW
/o0yzi6pMBGpWO18Ufp+3c26TzRuaXLSRpjk7aMzTsxwfuepaKO9L5JwoA5O++8l
eDvukEgiWawWPjFO/y2Y+jXqrIe5IsG4WAmBcX5RNCDU7T6f+Yq8CHNAW20vibg2
eBt+RjwympxPJ6oipR4dgBFh7yCpcnVL8KN4Lb8mN5caZCFsWEeXdsTuP3SYVYWF
Hp89nDsRAJtyfb8sb1/mzh9IEPe4ZZzrxSd6KTiRQ5uSHjhpZZFxKYWWC0yO96BA
RGo51LW4rZi+cQ9lc5U8MLl44WULNd/CyM8lxNH8mjWr5xbfTpOQ6v0zQ1kSfh3i
r0oMYlgUeHwE2rmUIgwXSNRfza/BRixe9GBVBmlWNMPh7K5zFA+gs/XpyiKi30hZ
wrgX+vm4lgBhW2HjmQ6xO3qTpMzLDBsuWbJni3h/ADD0U0WW44tgutxdOcDWOBZY
2dKurcfMly6e+Zv3xmhO9etp1VQndoiVlhOgEgN9YTpdUVn2ZFQommPjx5nA37gU
6GgBX5MyGbpYUsyb2VHLIyoAP9QPVf0OkLsCqkmtri96GEAgoQy3qBJAvFMCeYf5
1TLSDs6C0atKgntzoWvZWsD6IetNJy9UWFAo666l+/UYAOW9r7VRNCAhKqewbZnl
IerUe8+Jsp790jrnlmlHJ0+DuLSJiuZ0pU7qQrJPqB0GozzKKjLrA+UkOxnX+9Fu
b6qt41jAhqHMzd2+KtDLeNS7z6RsYnLvbCuUMaFiFTp/juvcb064llWUBLwoauzN
7HjZibzx5Nb5xps60NaEJIdf8pf0w5ZXzsYyDiIm/GgxFqvlTYcUco5US38gyXfh
jGBnMRLrwMiYwoKDc1oO9+p9rK/pGALOFE3p4aSd8RedZ1o3tAThlVw26egzo/GA
RVN4h7n6ksUYa9ifsZhVURtFvbgwYYdbS/vqflSdfSOdCDRaiEdAthpwli1RDFwT
0pcBbB7EkjruST8NNjKXgej5T2fbcr61qmMQyJ5DFavAAKVNUnOX7uYrsjE1mysI
kfqe5JzyA47EkYypAF2iiX4DUVmlkYeGHra9BJJWffJCykjGtzy9qbhsdA3CuqSo
nLSRcJD6AqYc9mpVv5VG7McOW7bYyvv03CUKfHYUZCnTGfdq/2gGgiZymk+acsKo
9aegwzpuePG9ilj4RBpdNNTNPCU1sai0dYhYv7yv6u17Zh83Jmn8Yted/UIqLk7H
a2cjccpjKPRqQdF3RZmeT8xd5Ct4npHe5l1WSAOauc+6crBLtVg+e4gxuJ7VZH9g
W0W3nQFb8GpZBEsHM3emzriwk8ozLVHIdrrZ5T/NoclA04+8J0p274M4JC7DILvT
7gNqE48tJy9g7y7KeV9ydhBoxaT2YYgwp+Vk/ELBwn5Tfacm/ZvVJcPkh6ieH8uK
GE7Tyds63yuWxDAvZY3n9OWQ4Ijzcjhd1E9lUtdIxzgMbQRJDVCEbUyVMiv0NDvA
7Ffg8nTJ3gmv4G077nPHdxZ2fn7JVwtC+QFL1BWbUqZymaQZ+udUdW3HHNf7B+FO
EsnJ/5D7klneKkiyJ1PyK/ADLRb3aczZzBqRbp7JvsJia4C7v8rApx8OS1ff2wuI
X0kNgkr7wRi80gVJvB76089RveGtEgY221kg91CDYO1Cd3IzhP2Vi2tAt0uReYZt
NQvNNV/izVWukrnX/1/YpMZ1erShZAw36bZUCrfMbBQOUmas13/t4RJVfJEZ5Sg/
8EyLSP/3XFWRVo+Qw56lDC+P/4RQeo0W6okmv9GIn6EniYL+pDLqkSdDbmZqeQ6k
UZThrydd4P8SWgn4BOv8Ao+Z8m596wCsIISE8RA1e8j+WmNmCodEPKu2tW1MYla5
PYAbsdkV5TdplELfca5pXqaXJaG4okiRDiB4ogg66Pu1rYDGAa820lKKa5VotTzn
cWNaoApwgQZKzSNnhR/+ESG8Cq6SIuPejZVB2yShkzyRAajBUn3jiJ46IJBnDgPQ
BlWO2UBP+3I+erd555EGbyTIVbseVxLYs+0ggWhgxPw2My3U0GWZLjWsHFolewFO
+X3sz7Rv8YL5zZoDlR2elzhysjcqlPan0yyEdNgsliv9qLqif/wu8Upv9OFj3oON
METhD+dNzhE444w4hM0mDxRP2Kg9EQlI4QYTIBmHlveDidce2uxk0YWNnak4+bwu
vf0Nq/4vlZcLMYb0Zb5L+1tHsFjSfxpLw1kOgCcImT1l2AwWxvHZmrTRe5qTpBS7
LaTw0dyo4Uc/AY9ie23hDat/pDOG82gYDFmf68cfraB4V7tgFkxdWOCJ3vM24n3O
DfGZKZw4GI0AR0NORihyu6BupW1BGlovgxPjsFME2rkVB1vVLrynP9JNDX5m+mXg
H1J/lQfdKgygBqNs9Yyub1iR9kd7hiLIFxqlhDSb759/v0e/u13URVFNlxSEcxaX
E7xbvrILwZs7/yloPAz/A96R688pTZLWW2ru6rJ0Bg9NxYBtREKLkqxnX7W2zss3
2upgLD9R177Hy39yU1/w+27RNqyxeYIzG+Jqqd8Z1alQEyMsJeRqt3vVPNwI8W8n
KxxJIKZHrQphtKImiwSFQeqWhpCADpkKCMnjoWTRUV+1kydppTnzj8z3J63jtJX8
8211qkVDsBLsj/0hEmYWoQYANUBKYbKza/vSbrs9AFVa1gbLbrwdBnwBhQ7YrTJ6
yuN6gtPd6gnJ7wmLpYnjLDZf9tPZ4oOvqfrpqr5FtO5qIyjDVGjeS77fg8IlZw2X
vGFOc8ESgYNXtcelQdFVpDmBkvBawzOpMfnNaXsZ/K9hhufX0pzJ+teJfkn2dDZE
RrPJITHSq6YQ3GurwCHIps2EtS0FivwR5ExpE/hgCCT5rGUHCkTXDe1zAUj63p2l
p7W99bdBrCa1ysfIJ2C4aaIsguYco2I1Z8WLaU422XouB/pe+Ny+xCRyVoBBkOz/
+B9ksf262TiBflTF7YXANqD2uYJc+FHhsKSJSpIDI3m+xtwAvzZEMlikJAdQRmcT
mGSCP9sGEQAtRIgDd4HUIjYwUARxQ8/C77a+DxWqS+7fa86VG8QTwBw9AlL2lZ1N
UEnXPOD7kWmJ0mo0Agp64DSOgSGAabZbX0r/oc1AAQc6PS/bkyY1KSj9ceULq0Ri
jEKCUz7r4/lpuGS+PBqSpvoEA5OmGiENcgerg+LHE2ohejyA2fMycpbuZ9zX2Q0F
ygAk9e6LTxFak9fgU3SWglIduH/QT84dz/nkAJAsaQMOxYG7laODmqpykXsRkNY9
u/IVmZIJUIVoJU4eviCyIYGwikaWo285sKrUHnrjC3Cr0rTdfWsStB+kwVhCAlBS
xImtFs4rV+9QZcIRSow3LxFSuQysr+IUAzq4Y6FcOkbjs/zyXRC3NVo2FPR8lxbp
Y+t60sxBniCRe154pRRD3NpPDJ67n9AWHCyWIfdTVtITeMA0gj9XoA6Q76gIHUC5
GSGL8x8eDGnwBG7TdBUvd7DIjW0YTaBOyVBd35F3oaoYi85ahNiBf/CdOfwBeddE
us2HgG0fzDjHLj+rf4+i8VTeOXTCeak+H2GvX/e87mJf2+EeZpy2PzQtdTppPCwa
/xLFB4nSP8uIrBucg/l7xLKSnN7B1O8iq4gjHrtAezn/Xz49yXeF6Ws85gUl19DX
X7gxS2I8ipFovjfI14AQYB46TtqPONcGtb5pTLWwap9aS0fKhp+5uXeWw73lP957
0bWE5furVOItZLrcsnVyA/DuAvXBRRGvIiuoLTIYq8vavxc+NxbIFTbZBbmpyGXi
UpIa1+3KTH8Iy01bqIKh2u91XiucMN9MSOqmwtiShs9fNogRW7KTNRrt+G9Z8yOG
rO0X7rixDUxIr/hXkshxmJ/jgIADc2RsP/EhMq7jmQOLa9L7g5SbBCECkRQ4R3sg
BafTAvzkq867I2co8ii5O+sr7c9Qy8SaUMr4xffYVixNiRUhOZubpDmsFIlqUob8
R63YM3rPP8UrkTuO93fp8gLWe69ui89L0HQPTP16CMcC8M+LfYBU9KNQ/m0Pi+Yf
BuxrGsrowgIVb+M65bcrscn+AmwUwf2d/6ljcz4WiUG64AS87dcoRLUykMvB7fgg
lLw/tmUgiHBnIsZRNFzE/vQYv0lLq53XYF23uwVOAUnn+IA+I+Gqrto+oZNrgtL1
JpNLtod4YutSC+JfPG8r3tsTuiqfAcIjlUs9C0LR10WSg6Pmo+5pqTYkU77SHdIk
xc7xjKsapSQEIXhvQr8qprr5v6HP8/u9n/5e2OEHlcJg6t7XSHrsCm4xsTRgvWIq
MA1hjt6nxutdipEQE30+C1Q8R8ibp2Q/ndMtTr3I5wJ0eiMW6xH9zYfiotdAILPi
5TYyp/PFFjuxX9NfLG/CtN6h6I/yLwu6lje+fWCmnLuYC7gN+lftUTIPHwlmdNPA
G75XuMo0oGxKic4P+UGhxiF+mnjQptMsul+80NI2TV/UxwCuFw0BgVP2S8XWIiw9
Z81YT0qyU+h0421eUONA+uUaJK9urugMT6PHgob5ncuSqrEnM6VMv0A49d8+Xtfr
fS/fXU2U7a9drOWZ12WojvS7YT79uH5jhF7W79XijvvSf2REfHLVhfBUIlwqxemM
6mPDVGCLivSBFUIzByGmq8G+Lnog9UI18lIeKQ3sGFHfAiYbgQa3JTBQYtaOBBGl
evv0adbUHi85nhszGLC/n3JgDGXVx2dGbwrT49fI43Kqt7uHE1yICzw2bPLwkK/h
t/xcDDBc6Ff8BBzk8ps/MpLmNAfBxbRdjL/Oc/r/hpg5IDFDsQfwz7k11tWxI7u4
QmGiNZdYuvMnbKt5meOvWMTcUEZeHL289fh99vdzo5L+qaL06bQSy3moyw25HkbZ
+u12c1hjfbOvw2rzrZm1cO/pScIOhw1nm1dGT8tuVifSLmSXzv9FBAFw1uTzQTdl
OFzzT8sWCf39TVqwIFlJYKn++xT8JoKakUItgOXR0qqxnqtHfVnscmBWzsk7/zNT
GFQXYpafxkwbZZQIk7m1YOgXT6o9Saz7/HUc3VJn/sQdVT7Oy1ofziKyzKHtUZ3M
vJT/jJ4NQd5tBtY4Rxo46SjW7cJd3vF06XPFYXot7Py5pK7it9XCEJcBkxw+m5Gy
DDodiZP8p25xqMB56y+6Y9Y5ONZSDdKNqTLbgMQURN2hlIzT0/RQjJKjd9QvbG6j
CWpZW94QvJHVtTGhRVdY0B6hDt5M3aGjEf4vIsNexlAWY7Bem/Rfg4BIl+6CxR1z
n++3obwOKagGoWqh4twtZdA4srYzYKYE0559LjEHEUHTcsIk79NSxyDwFytRbPXU
ovYD1OhieVv2mC7QaaKHjO3YIah6SJbHOUWCoOzy0Z8e6tvQUIOtoDSBsRAMc0B6
MTtQ/dotwPmCFeuZqWNdx9NNbWUWDOXHqceAbAYOX1Fjny7vp2hgfEUZJOIBIaCQ
PwUfLfC8/+026ECGgxoOMccjV7xndhaZbN/qFpM6LFvPUDJVWpq78Gix3K0SxI0R
a/1oTtlfGSpzKZESSNep0I0YhZnO1rBy9qrtIq3fk9WzeycMqtdTwx9BMY7HNzZT
PcNmV1kPm0nRJKysFiRF/rnIlnV2WcSWIcXB+sRNk/5wfVX5htzqQZltoCidAa6J
KhWZXgIUlta1njO/7I85FYxn03qjBF/fBYtk48lUanYDPCDS6S4ibnSCEWe2Viag
MrFbICjs4L8sLexIZZp0NM9bnHo2c0rkjg5iZlaMn8qMK4dLNR7sXEJ3tcmRPM2R
Ah+nPVrRnmMWq/iT4oGu7hZORxnchYYBwO2sn43n1ziLFqnr6ic5EuwE8HMLe9K4
26ucDPvWMkNxWuMODSvoqb2elfdZuuQ4JBzeUL1Ba+pJMIbKPwDo8ufAzqk+OGhr
71DfdRPVeS45zDvDtkBECsh/jpcJnfUqHbWNRJF7DRFlXzznIWl7StMCwIG/Nh3E
Utb53vVz41fCjJMRqTrjfOiVsTsRXopZo6VBWtBELl2CY8thGQO+KUtDDXVbunfR
CTQc7YTswPZySkYdrgWTEiVAbmNv1R1ABWQ5VOXUzs72lR73yGHsyc4D3lx52WqI
8mluXb2TE7R5ODWymfp5CL3gmOWaaP/PRi0hlr+ILrY/22AminFBlIJo0ky0Y2Ws
MnYyXsyx7rcpwOzSfY8MCff9UwgILXyBbefLShDYo0ER1DkreWaxEQ3qKx0txUXl
j7gP/svK/FLP48oxol+CsBkPIdEEXw1l2hDI+OSg6ObznvMnkHrL7eXaCD5Tfe/c
tatgGErU0Wt0nbWV7g2V4GkBIzQMLgCrnmQwxxFFIC5nzwRtM/e0L1w1XASft87V
1AAebjPJuau++PXnJDJ6f+qM+nEYY3euV0haDCdprSDzqV30nvfeF9UHKg5UdcPH
BDsA/jvNQj8ip4Ihb7uy1W+bXOUsOcf4bcDcSXDQZ9X8FiNGtfTuw1XRbTLn4wdQ
8YHJ6E1doqh30oW9CHrjdJuhnup3a04hfSn5+iLU7PMCRkud1BT9BtLaTIYDDaKc
wqMC807GGJ5WkcUQBb4M9i8g/a2evbCKIgz306YfXQ2xir9ZVg3/44VbjgMkIdP5
uMTD0pxvBj7UTUaTPyfLR8WTlOBaGMZdhTgtpMZKQW0OPdVdKvwoxxKoQpyEJHSb
Ib8DKY+CsJAq76rOxEof6uyNBjYS0aiFXYHXtjYmD4hRvCPYWt0RzPipOU6lkXOJ
hqvSu/8HIqnKsQFxuphLqWNAPZQNW43BOFGv68APLkjndTrYjBuw/3qqjfbSDIT6
OXhWWamti0EC5EZl3pMb5zRLgCriqrglGRlgxXm4JbJo88Vd5VWfXQmn4CmeicPS
z4eH2sN7n0P/4gPSohGX3qJ8aTyV77uAdBMOxr4/ywjGFgFLb5gyZ8U2DQaCFeu1
BD5hmQtg6zi/p85/5By8/Ne09DIyJxZgIfH2n0DexgBfCw4gj06UFVkfuNmT2M5p
Vuo1EqPAVasYsgkY6Icsh44N00GcjEJjqXjIZ1AApBIjlEKubnB1gpxfKv6CBcno
69PxzE1AVmE4ERUJ+V3Xz2ssJ2NMTd7xxno70WI6QpKbLUO/aU7Sd1VMYOAzLpw+
Ll0ESH9YBxTWMyM48PGjPZ9A5xDqiq97M6a5U3pwb5j6H/kducdVy1MrjizLhA/M
zL/7OVgcOnh1lyTsQ5AMcRIymmpBBmQdOBMZ2m8MB3DGq0WwnQ65I9POWi5XQv14
fUI2QGNv+qd1anU1+ArpqkqStHam8+zCiu3+NzR7Y0HjrGiu2AvI9ixpNHEAIblX
EuuYPCDGv3wddK10uWbIiKMtJIS03hlCax0EVhzEVElLoWy/XEggW+cISKEnK4bq
wzv75pK5ekvUz9btGRL9J9UqfpUCOYfzojjG7LqsSYmNcyzkbRZyUzKIN4owSn6Y
eCFSdxIuLYKzxTEVi0mPQe5+5+eSDBrju173beDX+/wENN6JaKBySNeU39U7yr3Q
eHxi68ejdcNhvteZRoBYqmI07Q3y4/FaE1/bdj29yKNRkGWK0BSNmPAkAxpZxgYf
6qvukEwXFRDixh4CcWdNRZvtXE6ISRRpLyeWAHrridR1eK5/bUbFqaCs5TL12DYK
GKWfRcJ0zGu5z8lT0/A6GkjNNJ9whEYkqfQUUAdmDWE2i0En0Zp/b1i40maPqhKN
fPv7+J4P6bsjkfRXi5sl8hH/ROdRtagJBkw9crT6f35BuySQJ5inzjGi8PdeAQv9
HViNNYZAqC6CZCZRDoRKtvZ4stRBKkz+sGtQQZGh8jbi/kGCpHLYAqQ4+xufO/Dx
PfkTTNfa6cPeD+SCc/W1LthgDLxj8e68KmgCmfBhscp0ULt527MM9JbPSXVQ8+zq
RdG3dB8plCyDMlXzVwdTYd5iYz8NYRZSudNElGCQqs8ybSa3vxdDRlFMcOSIebHO
Aj8whKuZSNgKisJNsVWlrhFcjyyTEZnN+wAbXPti20NgW/sP/zHvd7JIbTRC1Tc2
BkEGyora3YT+mQ+ZdAR7z/rjyhw2KRXJqHe5BgNQFSRQ5BhCha+PgrpexwyQYQYd
21Joj1j5x6At9fMv5XLm76R3Z2Gi5s92u2jJBW/INoapNLDQrZXCmjsoSZKUaATx
aMc72RHlZE/EFpr7K64D3zwbMYFywaTHT+PEIG7soHZkKl13y4NvPr9Vyhhxt48k
2eDeY22RxBzs0sKCBi0Hs+ha1BWm8SveV3RNdE8A3xHhmnAmckrO8TUa39hukd/o
1AIXb4ukjcSO4H2wJz3anUz4RVKXJuRc4DURwThRwXETjnDj9dJaq7CWpJ667QCR
ljfCATV/6U9izJXYcheBJ/1KiZVEQKzq1AGyMa9w2BayeMXSvXzju/+cYXASxaZh
YalH18H1lBm9H77u83GfKgNuT9V3haUHDujBrrxBzKvSsSp7pN6lJUW3PDL9Vxxt
jTj/LfFXRFDP6/gAYJipZY65eCxh+PqZEOOcL8Au/x6RHgyQ92ASyqsFz53lUiZo
/p6+RA7T0KtskYTiSn5EX94Wj9Qqpy6eCB+i7nEbmpXY9sUC7fxmDgK4fNHjhU+m
okz238tVmYR5FS24nfyjMoc6b1RZfeI8LYGF61sqOod3Yqx/oa11lhn71c70bMIb
iMUYnxsLnMMsBR+TLzf7CO3uIJMeFS/DwEL4SXsx3rI2uVMP1vmBgtIUOK+PixwX
jXs6qqIg7Z+jlYHCe/J//3qnH7MLkxRm5uQUnY9RO2KhZNl2Mx6UOauN0qvfxGBv
GnG1TcPiJ5kaZIcqG3ry+FNMlwKnvc3qc+6MZDHxewzT92BlXiPt2AYiOUASfyRl
46yt/TMpwkvKkPpYV5gQpBSwpi5+4J+WVkCrVOXBSPJqU3vaU1CTglebNcbRCaVM
AcbQTFCCXpIGmt5Fkn4n2PBwQiwyewQ5xfY+UIOdsqOIALjlYoqaVIIFu4yoAzU2
gf0EgkstbKm4Bv6EyD7UIHjynT6ck5D5izwdhmMEOiCUsXO8aCohDCiaeRetQTXx
vcAoDrXuEpSUzxE2zgv7QmORNTY3YT+lAqw/TGuP/XqHLADIrBxEXsvukqidmCJk
3hhjGX8XT6tDXXoaHXopWCwb4W0bebEROaBNagrBmFFnRnfBTlgkoHzrgHiW04Cc
BhNSim4WCnqAh/gOzULlWUsx4+wpOpvVtYSbx/vAb5CX5hBZ3Av6eGx9Scb6ZJ1I
JicdadXXv5k+Rgd/rNsVfesgecmLlKikCNHexpCl5NF3tGx0iyGxE7IcJPVu+COA
uzUWN3mQQBCoWldW1lVtBW2VxB1A3jjJlA/LqGcLXvQjLuMNf2RmRdNXqR4FJ2tI
rgrb47bxPA06SzJTVBU2RH67mtQZvUJkQb2wYC8MGoY5tMuFShN7wVvgrXFEXpik
MrzagfXiMDGp+qSW1bMTLyrdaTbe4K6i+cYPIVbRniN3N/JKD3ECMXIXZ5llUT3l
4p6GYYb+Kx/3jcfyBfXQrD+QpPAB1HQgk6GSeFagILV9oBwaJfSbF5HaqiJIAuH/
aXPw6aRcr++Ee0Yip3RCsaXLFn4jtN39s31+A5je9xFWNRU1qa6MHg7mP2ooZYia
7X0NC30yNQvgnv1r3f7lUQVPL5r7AWNaQHX7630XP3NIdj03PYtxByn+OcWQ7BLp
t7CT01B7xcLJ89WSjUwLZFKy8kEv6V4L0lOtmuuAeb2S5ok5U1Zgmrgr1ONl4sbC
Vf4ZJV1kL3/rO0oRbZaZ/67xnBtbGpTfVOk2H9DnvdRr5ho3tLO6/eN1gqvmi8sD
WUT4oL/9ToxJRuB3cGRcQw/qm8qaZB08jW9oEY5+7RAx4QeiulfJWHEV5wVdjTNI
TOSHshyxPTxj4XH+vXG7yBuOB7DFV4OFKUVDdHkBM9Wl51rybxboTGlSeBjh+mVY
HtbGTH07qAewgJ0n1cC8dSBPkCrDPIoIXbpRkYx9onwJOYqLSeKKUmcZXfy9Rqvy
+0NvHo+C8KJ8cpGm6EkQrTRwVQdbfOpfwmQU00lhmr6jADxrOeWYxEdb6d0/pm7c
38AA8muTg2hALURKIYzLlgXhuLDRr7M72DCcaYIbkkAmV3pfvhJWt6ZMSxsgz2RU
/fw7ziA0UJzCHDnZZCZZfArIYclQoz/ykzNE+XvkynNCJdnD9fAv9hJr+uTHSvBe
sZ9LlEnLlDraceGxAdccfYkLRjpXomWjqzFtfSafbkUCet3GkSyuzi0PKVEudo+k
Zb4wfhxnA9fiEWQFXxf2zHh31oqSLocJWl9yIR2q5/aFqfpmqppPoAIR4XjXRyke
hfPWAVfqmROPqFNW/5V9G2mMY5ZViULYS/xm1WRyhKoOSThzPuvnqQe0mk5Vj9UY
0Ba3xJ7g9+fuzLi4vJmndf4sjVLJ7qAEcDw0g2MS/nclP+zdJfqHEbyfWG5fWY4m
ycC/aEmAsVb4x8yop5fiX7IP8NwKKcXI9Cjrqto0WUSHC+RM2W0LCSIV4waIg3+y
wR8J4PMMKwkxSANXoZMsIJkK78I9hCXDl2imSW+P7EtuRg9mj4g0yNuhZyNVhsWY
EWdPwmFLj9tc6yHqdcFFk90URTGxWbHTNjUHCf0fADIP8EQ90JuGHH/kDo7X92bq
81G1SU9D4NlgvndqFzqxxActUtjAoljSnd5N2g/jurG+/IeiMjrykWj4Haphg4BM
dMNCk18eqC+ZRKMK2HOnw4zNDujc82xOPTkG16juhAj7rEIBx9IQj7RHIiYjkS4d
wP3olznAaK2Pp8GuF2kj9LDsvPgDm/YgKTcwvqRNmx05GN6gNGm7ECx2nqCMU04H
iLC4HG+qyjcZbgan2/9trP00yFTvQ7QJPem/gG9C5B2N83E5qKJ+5gaifeO7Alqe
sLtv8+4BT/6oI7tDUyKOGxSeZKxE/Y+HQQ2QgmcK9KTI9BGK05JZ5D7UTg8TA8Qi
fT5hhhoalnnA+MbTqrvfXTz5mwRwj+G9Zdt4cUE7dS68cjB5Wv3MLmthsevUu7vY
9MvRrp0++wrm+Zcfad3trRE3jld1kqkYo+O+oBRz3jPtq1yJVFxACMpmCesJYVRX
5l980rYBdhUv6TOfhoa0/cYAK1AvlaYrvdTXBpEhz7jmBSSqft+EJVYzw2CTNO5j
inxmG04SjVjarw0i8V1Weyt0OJSM5HHyRpgVHR9M+Cxs9vA6wb46CvaXoB3Qfu6B
Aw5gKnkM6AdQjwAYcSprmfaP7PcbU/HH8v8GihWn7knZ4ZXGjyCPuCYK5kpkv13X
eNf0zxUTSnNOqZDaKaBmffknxJE2gQJZt8ZANbyH6Z36HAOozbNhr4/0ZLpMXGys
cEW55Gaa70f5s5I3nieeLOZRXZf8nm8okekI/eDjft/jUhnauWjF+fDxu9kyGKrs
iyuIPNMlqNfQj5d/LiiUbnCMXwKbUN/CngX6MTMeKuULwB9o6JfFAfkoJvE6ruAv
YrGZmVhNxgyCZ4DRp9Q9x1h62Si1wLnE6pzDRolxRWb8EDAcuxocFNIXOF2He1pf
KRJI9eLKC+A+HowC6MVTAKmoy5Ra9l6LMftNY9MVt8ge1lBBu6h3GVZ6GXJdNA0m
uKDFfqUhx9A+OlfZy5UVGvcQUg/DpGUWvkE4wl7Rf9B1xwJED8SGo+5rJ7Pxy+IL
/xLI9I2WierPRIjHTxkJYv9Oa58wkSbhfmY2DocnkGHKsFH2Rm8y8SkH0KLdqWBm
zOoZhm+Kj73KYjxWdrHpU7lBtHoOWEq8zBaEKGucVnX36nhlQj/pAmYdqRBqh21p
AAdSTHCbLSMU2XBm2M+SHSeoHnWF9tzd1cBuav19DoPxTZGrtIYU8F+9ymXS9Uw6
GzqZAzbFynGdLWFsfPJ4pVyI3yANhzBKIbxruiKOj6xt2cDJEnbv1P7+GuIHHtxo
OyVwsHbFvcIe7kmCRqkwJkDfoWjFUpTru3IfnXfpRwBEDfCMs8dRiGs8w49fSJcH
H6a7f/k+1Y0z3OhQCDJYd0E41y925UC1MWpdlDXHP0AlVMuVCvnq4BxcBvVGI6aZ
xOvY6geKS6drxDwzCMAiwVqt7HpoUsuQn8qltL0TXuLZadZAZc30pOLzliS6rL0J
49EDIBhfdN0r58hGXSMtMN1O1r9vTZoSWRb2UppkKF8Efwx6BXir7VZIDc7xdQD1
M2jwBm80tQ3seXhuIA6Fgz30CI+Ks4m7DfUpl+CgU1o0lNWwkQG5gg8E9948dIvE
EBz3wTYzfuO1wTCiFEcIZvfVxkIeZPzzuFk45o+53NcqTvcHY9RbRH/cy2GKIxeL
h7JA4Z0eik7kNdm5ORPHb6bm0+AimACnlvvubsTplRHmKhbCHSgrVTlWk/o49ijt
6gtMRZJM7uBVDh+YqcS06zlAXnoSOCsldSPyRCLO2tG43KPakUrgYljSdzhcz0ND
sCeo5zSSJA0C40qONw2pu2CigFdzmoYvU+J9FVP32aIMW/lj149wqeTvIQESjuMH
eRiWedEZuNzei/HbdsXSlm9fhleuBb1Pk0f53YgO8pqJPmPkp2iqBqsz30rEavAA
2/Ine+w6xqDC0uvy4ou8AD5U2Qgmn4Iu2c+MmGeDIk+s0/5nrOoNMquFWF/EUtW/
jqX6hNeIuUsMNlVtHSkT4/mi64oyxwRP3MKnAeHNurPMCYRAMFtGxhIHFzqSo3mQ
cOQDg7ufYQCBYOIlPbmJvk/A0LeWhFFVunpcwK3KewD+CMgD5MWZ2UUu6mcQV+yE
0TTcOkZgBi6D6G6u7OGCMOcJLfb6dO/XLLrwEwNRsxz+KIS2Hm1KEimLI1WWNC/8
Mz/Zl6q+aWd47gRcA0cFX6umr7Kj/uB6D2/wO/dx0erTMF1kQNalD2zlvDqsGfA8
gTcC2DhboMymMy6GQQtOS9nPqmoUSHTyEQxa3zK2sYNp3Aj/XkQVcFzPHLH63S8J
9OkA499TpDhPwFVUy0AVS9WspOb6PSWSNqE9ESIFat189M8qc1e9cCjtMbB9bb7M
UE3EFq4JXdtRRpy/fJxsFPFZkmxqRbc+DmARekwAVI9LUm0izY/zlWnVRu5XZ1ln
Nip0gd0qZOZMZ7ZWcB6zxfAxlqs//stn04C779FzX1nv7gRop4OxusXXyDtbgnY5
vFgbNbvnyBAyO1HBaW34eigYf2Ihc5CEppGs5wcQSY/1KWhz34MRrHiK254QXS0d
tFDfTqXmDnhGKr8PMqMfWfqG/LcLLSRSl9bJBXDgCDoZCPgWscH9BQBQCcLFoJy3
fXam1YPlTQFWYzkGoA8nUQxK6itoWritnW61Hvmj4Je/LYDsgCUZqdjTg+qCY2aY
xARQ+aU841iHkuMee9qAE0M1PX/nVRWbJ7Llme+YBRaY8ZSrhEcoTzaRwFJApmrZ
24JvZvlhZay+wLHIM+P/dsgjyHtyPBWbLN1vjnmLw/AqgOL8vivi/e1jglF8WO2X
pPESc34Ym7FC4Ug5erpH2QVX6paL+gT/0nTlJbuciESP86xoXAQpr5U7tPFGX0eu
pIT5hlW3k5Ns3oZFMFbr9QHNXCRh4V5hz0caasRwgSXTsbe4ADJXE5ErTJiwmQ58
Q5T/SEv91uNSi9OYxNki1Kf+677EDHIBtKGC5mYfMW58UvfblYOgC5d46PcOs3fV
JtFyK0xvPvKSsiX8zLt233PDseyW0VmzFcaRF4mZg7MjPVqEPuWFV7TA+3HaTMPc
MfB211XSRn4+egd0a0SUmQs/cV1jegjnkV7G9iv/ZojuhMLKhhXTOU0fBAK9622J
JhLPsAnlH8cF6+lCBpBya2hKFTgNkrHrHFgCS5Y5C8xYnji2r6A7jwVd/jLWZqLT
CI46yUVCxyne0JyirIemS/qMxhh1vbO1lH8yAZzo6tsHP2MmCPc9YdG0oyFA9SPu
iUbRqHverja7CdQkrO2jAq+MQDQgBqaCiSFcsLUHcHvCvvTlJfojG93yT6d01v30
z4vgi1O8FhlzpegaVvWEkIN9K7u3/7cRT0wkvFntM0P+qImUq3vXc6QqDAhNBdDk
+nvDLJpFgGid+uoSZUc0/33LnyNQfD+FZLwqy2bURC+EVB3WzEW81+S1LomoSToz
kRpXE9KbRqS+p3WyHzKkv70WmvEasEzLf5CeMYv/3Lkv84iH2mJwTP7VVz5s8fcC
NDA/fj7bIx/T6bl42EOJXm6JXCJ9xKHhGarOhMuaUVvQ5Ksy0OkxBivU9JCmjbxN
BTlNGgBX2Aq75aXqsHxuHVmsw8gZy0YAPZiR4aPxZxbb0P5x2UPX1sFhocNu3T04
14tF5U8mzD0k64AbuiDPxL29kgqtPlaTRzbCUoC0A/RXyWV8YBcpviyXoxsO8jft
DoOxeIFWJaBPoreuH8085ZJMORh59YEzxRaK6qFsCPe7h7WCVx9007MSrteOpim2
qiQbhm/MkUO78cq62lQsGGQxFnZRR0oGj5IqtT46M864Lr5U3kZE/MtB+Ol+5LG7
qvQjxGHdmjiXT8A5HiV6ojI5AbfdxhKXcwfl989cL/PIKPzIc19lHgdAuOSI0RCd
5SQENdEKyZJBjByoNsS8KAdg+TLnIxIRDHLbWd0LIhm2YKXsPlpHYHfmksTnCvH6
ejb9hvczUedJu+Ay4CL5C379SJGvoknJMzBHyGaXRPFo9XPruqEyAoalB/SNmm5/
EshCZUO873q9Uz/lZi/iGxFmPdLVUtPEriMBpmL04EKuBXsN6GwOYpF3jL/s7VVB
CBeIypcRpVpsrnzMH41+KMeMU9ebM1UfRTXyfY+m1Vfb9Dxl3wmmDn25yTGMGIJq
U3P+D7J+SKZ3hrnZvHcGRe251s4/N0QGAdko/A8AQqMtddKpZZuJoYT5ujHitnKk
btTxglBBoJIF11nr1Ib32/VJ8y4LgcMxImzKqNXD3P6ehXLMvKfR9L6eVJeqIkAy
qCKjMlkaor8KOhDUUlJsPqmrFqABOZJG0Ks0WyFspKzta9A31A7pLWf5x42TEUwq
26hhV4ELFSW5XOrhagp5T3zsbSJvZMdW5xUjZ0Cb9/Zc9bBkPt8BZrF2JXmVGERv
uqHgLWa4Y0JergFOt7m8OORxg3sEx2mOsZyncUJyynV4Auq4m4N16RQi7OX3tQTa
/reAy38eIOPcr1xjhmtLWeEpLgz4ytCweL241BGFeI4ydDchxnQ66covJqNIdVjD
OVrbeW5YJopmc3ZFwikLt/kpWYcOOzBbuskEdU2zbzeimbjHjR+m/J/JR32Avhn5
oWIKFayyD7kseYP9XDO3W08g9HxyJmkclPH8acj97ar/4FVIcw+1TWZDJWe1Q/PV
2wKeNQD0JByEoJCGC6GKkH/kQ0CDAsd3WAy1R5Ga3+CjPjpd+Lr7quEnf/lpOauR
72YF35JnKZNtVe0U26PLG+v8HupBOIJ7hqmsuFEmdQP74dwYrVFuxiTXU8R2guny
KD2ebjbLdg/SjghLP+mIrHY/p+IfH7Q7f06vIOMPvmcAuJDuY51CueZIeZE8o8WK
mlKNhK2DGHifEDz6kyu21HISmcB60caUIHgp7eIBoPA/xIL9jv/pVF2EBbuVoyac
+rvw/lsVgY8Hs/wAxBameDwZAhMGZ3fb/HbBt4WsstNPwWp439Dq4/vzvimXjYs8
yBp2kDUtWD40HF/VGLmX331a0Ms4K/oc+ewHhyr9PoKaSJbBLvY3Q+LTIeYUlw46
fqsXJdxLQZm9o+FT54K0w9wVUAq3AFQdZx3i9aeVL0xWVHUtF13dOOTBLaD6kkOa
umFwVavqoYK44fbZo0BCAo5WtTKuAbIcbnv4Dt4muy5onRGnG7u7D3QzFbsPnFfv
LHn4MOpN42YHoT0WXVKsK4BrPP0NLUTK5dSXUFcPIG6MB82EQuT3UxJGNyKZ3O8Y
/VuwwR+eSnQ2IIGsKruW0GZb+7o8wqvGUxgMsSn161Lq8254KCr7/RevBksH2bN3
RXkkeYK8wPAD2gjLidmZaHONZ8q70kXbQBT+tcQvgqIQ7bn6qBu3fIJf70HF0TWp
BHKIpLJZAUzyuRVV2SswLZ/SRrbnBv7cfaL/MwSnNIaK/ehVCcQXs1UV+LHTNOJE
TWy3cAl0HJ9dj2lfehLsQ5ectcV4Y3cIMT+9J4zcClBcWNARMp/3P/u6CsxKtZaP
dhuhjtEm4FfPU2/tJTcAQRz4oUGkQ1C90O9M1qKP9UymlfJSh8U4/xHnd4NwLoR/
VzvTeun1rEBJp6P4BqPQOGqonQgetOpeTPnLeWGKOQPL1JMplMoGgtq9DjJzKV7d
3vCfo0ucT/e9RJvtA3v6eeIhdGx7NwAd2A4l7eUD7BZdGhV4hvhFKChWgpFeEvOj
3h0XtQHtIxSj+3k5aj+G7kr9ofapKQH6YjONRv7PS5F2Kw9xb2AjisYyHzk57CY8
uiluaYBgcY4m2zCDcEg+hi3NDU5wY8XcKLfs/KZ0IZzd5HO9L8k68EhBh3Tq9MMt
TQLD+hsKulgGIv5QS+HoJyvcMrEd+mtL5pFAy+qNoZi4fPC1SpLNTSdqm+jvSnTV
hVKrWfv+l9ATmDKKWrBUFBriW4x77xekSitf8VmX5dsybiDlv0FojhDjflO+PRxW
CL3eiwX9CBJ/lfOI3LcBQISxA76mg9GCGrVMNuqqrIMZjgiSlxpg6uGLDMwpeHVu
3tTvw1mS0S77vYGvTRwq6t9hYXWaGe99bcDwp8snXk0O242WWWNd54WxWRU+8CUW
OZ/dj4A/NhB9D3Kl+gH8AgE/Vmz8wcZn+DjSeGA7boXq4Ycdfzr9siEloohksjiL
khan2FcQUGpCJujYEVVVW3Yuk9tNMwOEJrbAbx4uq6SCKqDcOTQnr1EFiI4Z2wd3
dQFb4tACz5kBuUAVdm3qIyzZmSJ+ANqgQVdoLzg8oETPSaaq2uhe/pFvilruDYwI
POLKVmNLb3UVLo+qNlI7LqJPPrK+IpoY7Dn6my1LDZ0DbAKk6fETlt1Ehng+Bwxd
aulj8Bs5GXu01ETCIzdlXtGzALl/O9HAH4BOsJp+W5TwfNcf+wZS+h+kV01HzxSE
a02v9iWyT3p8o3EAmlJZuD6jPR9Ob/yHmT5Q+BOZnoso7Vdz7wP7LAgaPFleXXQ6
HWIwwI2GzAxfZyuptF/3zPI6s36Yd/dpIUVztl7wNrxvE58Fn2RN/9Zcy74iv2bz
ITQhJtGnkEo5UwohzZSGTEXr1Ct8l74GKRGOyWeIHhXYNP4MBYZhq958XNO0bkN7
1r3zxtlRUnQDgNV2YK9HjjVIKxGot+TWNx21usWE+4qtFkGQBplGMH5vAOdsK8z9
5fhK+0uWTA3JiXQmqGZsQEH2ZJwI+zzbFgsZD8hkVlq2fAImOZz+9xJODUyQUWDZ
+jWGIbfIjs4F7ZUv3DKV6+NnBBiuD1WZsTkRhm9W7bMqfJhu+hUmKXFD9zS6OuBP
CcQsqzGvMZWwlSLHc+FlFnvbML4rt064nApAhaGyih4PpAapsjPC9Efk03Q6qYEp
dCsXJZ6BkcJv8ExaVg1Pl1aXwEBavTRoyDDAj7isE4YlmGk9gFRpvDSFKHnLMOZE
ZIXAK1NPbULnUBNdETqJK/+HGrXitS/Y8D5H7cuc/StHNReLYs9fLiq5C7VIBUbo
TRo+mIQz6d57q0QnH/C4tz9lBCClOxKe/e7vm59EeaawwMrjkyOKZ2pvkWVWg16T
SC8NW6kEw+HoxbBl3A/GuY4uqe+alS7p44kD2IivtfPzLajlUjkrNo8fsqWWWU0F
ngobZqPXKgUFBhEJm5cEi32Bt/FEK7yVYX1GIAQ/nIWQ3bqKotYoD1gICELTC9eC
nymjdBWBqwtey+Qzu2k2dpMc9E+U7V9DxymfPMqx4/2C+MATxk5xToTJq5Oq1ykE
jRA6IfvRzvUoamWmjCnKcpZIABU+mltT0M9zuFsKLqGHwJr0uEGF4byjzgcvyBbU
0iTZzYrQ69Y+rqCK80lqGq+IrZYMhCZx7monczqK/izb90B+zQ27P2MvfB/+Kgzz
K90WcCGJ81i3DO4pCpgDF8gi8ICIjRHOz4ZZZSviIhBwL8CmjT0rEFeH5ZAoXMcA
WLS6m+mmSHpnCvxgwJq6TLVCQo4G1cPlo+6FqrrU/ymar8GI2BpSYiF7RIPSqHMA
9gFiOxRyl0cgXU3FW8efECo2OTeA8FoKckC+Tbn9950h/8X82Aydti1AA2NLnld8
wri5FDxwVGz+2cVf1RzAirj8GuJ8pHlsGE2zbrnh+VgC63IiUHmITlx+njXReqRU
/Fj9oHehQGCEwgPOD2bKpXsZnEEw0BU/vsfxKFzcN9jIScI4cTkFNkWR/yfWl8q/
HZixkwU+8reShtIa84aT5QoltHvHFCnmTavPWzRp4ZA664zRjAktHRRLLjHhON7P
TLVG3CVAcuJBhRT0UNMOB5MlsP5OCmftDmcUowPP3ejbqMpJAGydEESmYeX0s6SO
iG2AyqKr38ODNInavwfru7d6cqUoXhm4LZHW8zHJ85e87LrW3OpR0dsMOSLiJXVD
rHg8X+b3heVj2Hd2M3MAusUOqKncGAbv5USBWdjd94xaotsoXJ/XT28M85U41cuZ
ueDWROKcugyaWIxB+iVghvrgkw3oH3M25c6cwnZMC9atD/PTA24KnHi2hJPdWMFn
EZ/J+4tECWe+3PmlpnQDdQbS+5Or7KZ4Os/XArkiTwrU6PuSMHKQA1dNOX4bsFI1
37G3a+tVtlFnSJvdcFiaL2xcv1ijQc2H9Vk0zPyoL/sGHMTEMJhhtnP0GZJ8dbaa
+YtKpuOxoQjX0SnPn3mKuHYysrlZmM2qXgJGxCzptS2Ia1QxkK5XEFl8+eVFK0zW
uCsaTBHPv3oIviuUr06LmeszKD7fz3PtdRYyMKbdafajskv/bI94m2eJrTyS87qs
0RYqdDEt+8Q+GAsuZ5cAFJ1wplFAbV+qRbOAYPwoWyFk3AeO7IVR0fyD3a0rxiCf
OqiMZo6Ef42LWt9zRBU9c0r9gXMs/NhBxLzhrjSrVi2JuzNXhCaOIoYmDT+hjCCl
oR7Oi9YGocYOtWRcG7lzGBzQ2O3+5mE/KcUOY30N3wsuEi6DqdgF5lheOQEXEKET
hAsJt46tpCMGeR33l3lCnrrml4e2P80KGPWG5lzG4Cgdlv2WifZ+fBbVC8v7Nd6p
hHgXgUAWZmX03XtpJF4qFP4oaGPsY4BcVwpXsBkuSbtmRNn+rcZChVyJyw81XOtu
42DqSJUMX8iI//YgrwkZOermrribeTEZe+aV/F1DnRgi6MLnSE2Y0KdyN6XZ+DDQ
YdMZe8rxJ2QhmXg4fifWOPN5Sd50U7JQWnThweUODPaeYzl+6lwoEEPhnY3J1u+4
jWo8v0EmYAeRTKDqHVxtsmNC2tRG/Qa4gMEUKxE1HHHT1b/c+edvogzVRDRMCsM0
FRQaCt/SQz5GjHTZcfaDpx0wce798fHJlJY4KFk+wsnYATgEDgf38owrKpFZKKPw
OkPLGWfhsn5OHVeVcMIq3mWNdoLFRfDvV0P9xf7ado1nC/o26rC5f5Vy4fXohf42
F38k/pcitEndfIXdpjFR4AxzjUhDU9VP7t8ZiwWH5xNmV92yJUIduRsQY7xKHcdZ
Ojyo49+ABjKoyFsQ5rQYVZn4Xmha3ImUkRNPrXb3HXaqcX/dY/YFgKlHKCg5CyBe
IKlINMtIRBdH7UKDVMlJ0ET41hVOiCORBDCzc/AHnPfpmzWofP/Kc7iO9p7Dyuvd
9wrELVF3tslM2l81qBUqIURC6nJE+KkIfktO2f5mzyrRon1TF0TQoh++t8fm/NQi
/7/8dABrImBF7GQgD6V7n7g8yoPl/jrozK3/H5ojPBMZY3Wg0ULY1zD1GPXggCCK
cs5qr1dySPYfn4akwmZcMBWi6Sbbu/TgNSxNpZS5ikRjXjri03ZeR25Ykack8PGa
+GcBOziYeXINHMcn/YGJ/jkv1P9RXQ6rImck+0ZN8AcmJSlcdk16Prum8lpUfXvn
c/skIk11TKuXX2g7hQ2Vu9B630D1g7+nh+ZU7W4jr0A4Ceag8qknzFZr8B/M+7uA
1YG37GO8iCrz722GvLu6KJZeHLKgkEGD7FChzGqJCwAmk6A+F9bow3FL9e348voZ
tBlQ34kfd5NAXCxk7X02yf6RqXdwomU1lq7dNjzEZSpOAdyihK8eOAN5DDGfF7BI
8DN7uKdfkjmZNaxlLmE5xjUWgfV9zl3xDX9yGm/pUWERK+g4Ff22eVHalYs+k//H
NFdXiUZQ5/F6SfenO5pUYaGyaERbaxrtbgYX57g1DbYzFRpNZSUMALPyKTIdYEO6
eBaMTNR/tJ3RMlVNIblSd//ItMc6FziqlrZ9oyOTssJqwt1J/PIDwftHufhClFGe
hZIvgF8R8K0yPLOaBuyGfGE27p2nde3RI8mtlsApisWVGr4NXryMfhiS7p5npNEU
x76ofPj0FeBeFuXhrcfhVKwAYo5kG+ILzYZfmCFweKkjlJj1wd3u9DmonlBcBIuz
ZDvbsGPjA2S1uKsyMhhsLG5tAyM6z5I+goJ46TjeS0p+leDZ8Yw7MwWUkxrf/How
jvnmr0Yzi4cxRR23ypvoYPj1b4wJlOwrddCl36tezfjrSDcL/2k8k9LRoKdbIH24
vhCku6NGUXdTfe2tv90ntgnfSAiUT/DUOiCXjpcPXiiWEgafPs6eODuUb06uPCq7
zgKal5ReSIV/K7HtwDJRqbOxSh2ZvKZvrKp0T76k5FFPIJNHa3FijN8SUaq79Ej0
11xHmybDHPeKIgeBL6lcfpGAo1Mcwnx7F3HlqmIdbCByfePXxS21CjrHFX4OeUct
xkyzq7PuVlW22E0rq+qaSzLP/lxCHbabWmC+JY+sTrfxFv7echVgU7giGRzaPZdv
pdtjsfC1HUHO8UH+LGkX3n14yEWqaxAlyiZ45V7Rp0ooLQCFq627LZf9Tk2tgMef
WxuPzwOt+5Yd8HRBeBfdbUC+tbhDTiV6bX4NkcEAlMSd2O9q5+xYjcvQqxg6d1KJ
/nvfDYolRXeQsLl4mnsSQZuBGRuBw2wgJnDyeS7//4nuIU9BivoE0MuG1IM5Ftxq
kfGJvDerzBwuO554+5ta68Nc52ixRBR2eiHWf8xE3tt4P2K3PadlJ7/iCYM/g7IR
qpVfpgOI+Pmpf20pl0+4gcdbmmoE606ZV2/Nhvzrw4l1iTIIDq6tqyetVXGQpluA
PGYWJQDtjGDXngQ9HtzL7bMMJmsVGrT9XGGVnimLPMhWE2aQV5fNBDSKef2oUFKw
DHgArngwKOKgzBGcTHWTHgrhv+01Kp0T6gpn1S70FPXVmC6nYJwsOY/ADAV9Yc8t
TOX01icFUETztqaJx1dMWiMvc6Hb21qcnSin/LLZSO7CWU46Hg8DZZXEkO7gu3WN
3dwVjf4KyjCUdnaU5JDSu2QcB/GT8RjOHDNzOkSrBD2PrLadstIqD2Ng4j+OqHUz
qQEQ/H/IROt85V1rcG68C+9EVSvaKQay+354CCIqK8RpkQoE9NYFb5jS45taA67X
QjZNvLFS0XKYpCjstfESi0psi5ubmPkIdXpwm8PxrC67oF9pOIMdcTp0Ew9w9EUn
xHbF+7kdNmbxSS7XhEeBUz2z8J93zqwbZS3vsCazxCva+DqiFFCLr4s9f1NmhLKZ
db2SXTJQa6r1nNeoPoNjhFxlUEQqt4UafJ4thqonGAJIKZ7vvJZz+EzUB/jPnCJx
+Jw080o7haYgaIF3+OQya84bejVPSNPXlZTtuPk+w3ezUSHmpiZyyx5HXLLPvX2E
brzBXJInXYg+PKx1ZRuk1M0aUzXPfCNlSB6s2bqqgniZiq5A/0UR5FnefSLkqyP/
9tEPY+Iop8lE/6Ok6lwjvH7wV/SBGeCaiO80KE6Gn5vdCwtJGp3SHI9rlwdul4Wv
TF1LdsbwSmKWVQqLxTKodR8oLEngy0JqVOaQmxvx9ohaO7X6Zi5SzeHllkzCURg3
rlh8M7zL2vbmAm2QHixyEfxxYm4rqOsr1+PRKGRBQKuU6ben1aWIDEobPPfTLs6W
GPbqvwQPvCM3hKtXbtTMkjfqlkxYySmH/J1fXJry80pzYkRRsRKxQw/obMluKRk5
4Hv7SP7AD/dH8PZY8+UFK7JJkbNflhCF6YsUL3x2A5br+UYJfZ6mvEudVHFaDq/e
yxg/d+35uZfBYrrsyEpPy2x4gCNPDa+fLhJ1tQ+jFmUTHLs+ilsU+8J0u3wGCS0D
nNUoDSJuWv9RGsGG8b7Zkt99V3uAJro1ypeoNHr3kbvNYIFd+BHmmTQyakDfBV7z
KQvoXn1YjT0EAVBCo3vDGaVo0XK3wBOQzZBPAebqwKZIo3UkYmPHZsdpiCgkmu8V
E3AVfHHjONuPIHdZzSjwelVl1+fEoo8FzgSgoTo7VeAWLAOUOET6a2FpiDv3LHe8
DqDH4NAT5rhEy77QcMUlu3KB9+A05KKVSE4PsHaf8GYqV+i6ChGz34h41bAjKpWl
3MR2SSgrSjz+Hvu12dKPD+f1VZcOyJdKfvnEv8IB9WtZ8S3a03US/Ob+Hfzz6xwK
fB1hVxjjyTZtRagxpfeAq9xUMDJlI978TsA9bDbnmWEl9yZXN9woUK8uylPDu4LI
NOAFf7y8VFhUZvBln0yfREj3jII5P1e5d7ExbGRxu95+kXgi/kQCJ56FypNc6Q74
w8hvctLYdyrTA+gGlmhicqJPC/p7B6S8xhNzGcEM32ls+x7oRjXqUqc2XVQwd8cv
yG6KJIKsnBTWA3V49F3FAzmjEzK/iOhQhOdtBKsTTp1187p3ti0REWuN1yA5HObO
1thQ39Gx12hfhoknDWYOMHIoXUOCgnVSVoIxGsDJNmGWdhflPhgcAiQAXGUnUusO
uZCYcTefH8XsjnE3XwvSN3BHSB9ejbK0LmMDhpsywch6nYKvHkXgUyavUJxhAkdL
dSEMJqizN1HaFluOpjx3+VI3TA0VDigBqK0fP0iYFBIyKL2t6BjU2gvDjS34V7ln
/jMGdCPl0e4UT2upGRzfW8eApd8pNs8RgEOxIRLzYa1LHhMQCiOFcFDbdhuM7dML
EjRdXzk2JMI4WQD71wpSyuoxIeWZTy4b/gKgGumNx40Jx9BmnhK7C376txVm0/zr
F/JgbUInU4pX4vPk4963OlvULF0iS6jTqppIWZmzZN+BO2famqHUVe4/wFmn/36E
PBvKUMMvIxepA87uUkFPln8do4j1F7QM1Cd6X1ySGOVSAN4mNVU0aRoCXDKcL/pn
dtVuGbg0IUZCxulfs1On2evYaPLxD5drjT0nsmHJQCGuJgg7/A9xVbchJojF4OP6
Vz5F032CK+7eE58vlLhp5jiK8fRJaKvUhJ3pALAsHiRSP4eEh9Pfv2Dsu8T1jYPr
F87EB24FdwR91tZ3UsbEbNuyPaQM+WB9oSRVBMfQILUuftwAs++DV0VQKPuQgt06
jqTSsTf1fkTH5yb9/YAKy6+VxCoj2UFu+s8xQJU/tyTZ8euZXzCYyf1qSCyRm7D0
acHZWxIPLwMbSBkzP9PA2qoG8ZlfuGdwXwsICWEH6GV7XNvmsEtVzrF0eLe9CENM
xi3L3MeqPmsgikSGSVR8rvF91odJNv5x3bLI16+sh6/DWjA+RONsLm1+PCq+p+BJ
OKSnEzmBnJxmkXJijjSoAWANl8u0kxubqT6V6MKt1iELJffNq6r40T6Nw1JgdORa
mR+0cuDCPV7mu89tHrGiioc5auMMAq7kQDE4oJpJ9uwr1Gh+GWpfZwf+UbP2ASoh
gb1i3Tz1lIwj0WwNF1QbN/Bxv5Av1GLtJ7ponLKclIl73G4c/Ql07s5xB+i17r2E
iqb8KRZ099k6NTQIYOZ29xrxIqr6PoUf/f2aEvqXhTDuB4fXeHFY7JHzhas/ZAS1
D9oSdIJ+zY1cpIhQ6wbhz46TaP3tb1zBGBQYU3DnHriL6oo5mor1MqdCmHT+0qen
xhIOwdZcOPyUVb9qOEIWI3J/IDcjHSdH3JPpNbufGOSumliwa4ZVRJGJlMzWPKF4
JtlDDB+i4GxAo6CfF5SgfejLa/EzSwG15V6ArutGwZ2pDJymHQVilztzZuSS1rWK
MIQJQl02qhcHZMLfE+pHRHywS5mH6p4HWbQzOxSAwKr9+NNY2lgsb1AtEJMJCMeL
Eyknucj35sP1pD1Vmfa9Do4S7GdZGjCRuwrqdecpE+QRXPmKrS2FmALPeWS0HDNi
2QCg8mtyX7VLEeW7WVEeeuI/fBD5EI4nJSmBy5mSA4jrbp04lgx3ncIDeA8A/wHL
G6pbrmgyUpZYrpbr2GhYTdpceAhPfUj44112zbcvci4fKF9FzncQU8OqRLr6Xh2c
V0cUFRk3i3Ij0QtKBos+9KC1gnNqnYHvZhPx1ikLVA7teyOOR+k7Ye0xONQhaI0k
oX4RTVU6cSyEdPCJKshQwktb+uTuYCJZrtTT7DrbTCRHYAlupf3BYxsW0qHWuZvJ
l4qQ7nTODkLmHvsAACL4jteYp3eL98cf7ZAQxQRchCoA9PSVK+l7Q8t6pQH7j+rp
9WvLNDDQshJ3j4enykQ47HoU3t03ytki55o35v5lCJstU2KEvSy5QD7hBpTYAGKO
HOcDVipcS+ygszsRk+049sm0cepy0kCi9hCbr2XhbchlXld4Za14mk2V9dCmXdaf
daFd3Y3QLMi/PpuWgoK+aUXF4zc0ftwhKhFkiCZGtLRMrI/UvQEMqTwVdTtBIiK1
+oKZvhEKCj0YZb85VIj1GCNsZ9POkE4NbpnrlsMu7ihGfaR/dnLME6tOddzvI7rY
mA+JGhTPzssLHgtmZoWmhDX4WjlcPkPyj5BQedqjxhRfn0Dq/yUkwT/nmZ2d7pqn
fYFgu6FBYxA8rpfl7pf0yZHlOFIKyJPxm9pPQuRsNm4TqElAK6eGrDc+vEt6rQX2
8VHB+6z9KJxrYDVmiw/IHBU33U1I5Ym+ViOyXlt3dESVF4C0rM77grUmuPwkdqnn
Rf94rZdSNZTIZswIXFkUh3l68BCNAzELN1Ap+g0QMveMJEFX+Cbt+sos+gl1r4/f
zgGjbJfLOf6V4tq8/jQKLHwslOM1ZpK2My/nSEvdkDVukwDhbC3nJ3lHcY5yLXgP
AtYmkBw2jybvlx1y1s/dISm0pV0SgeANcNA03qmDyaWEBxfmroOVQhpREVaw9iZU
PQ2ieNAmqxJ/PgEzizblGRR5ypEK6qEYwWhO26KGAS0MOip4B5NLi461iM0Pm77n
prU3p71NsFl7ClhBr/R4H8u9PymXbE8Cp4nlgVKNiyNSvgh9aymPcMODLSaF4F9m
ucg+WPDAAx3D2veCUxyxYMfcYa4Z+nCPntRkppF0CWQIHnhNR95rbvt7C28ze2+E
QPXSG0bn58Ek1hRCVy09GXbm0bc84NlZR9kLUJGDsmzOXfqBOgc/QLIkfh/B1E7d
yZny7hJ73cKwh019AKvCMMz2zx/9Iy1yOxHGfr5roFjehpA8qRRazA9ZqFwGHF46
b69uVVPHKGsFGX4N6LBUU8ljQFKmL0LKqsiywTOUj56JhBu0uua88ujGJ6gpH/1+
oW0GXdzLF0WvNvJf08TtDSB73fPvWkzBZteTllC0QHkSKGslN8mbYIIExOpi+S4L
TVImXPc870OHlH8FKiE0lkmqzjQhBC70urDwnMTToilc4an9pS/o3FwSQGlQNXZ5
Mt2K0R6ZZJjgCSciCp/TxCZ2+Yz955e/BJff/++l0aIOY0Eyxz3IdpFIS7O+bjqt
XSQZgjUvNSmrjjJDy420sfBUWAepXcrsA+DynmXKanvdGQj8wg5KvEnCU4DH36vs
Vmkzb/3ZInOsP6REZWErqtUGahJFihEFPBG+/kw2E2+jsMlDuxZyXlth9bo62bb4
EXWZ8MCrbQka/BcBgKp9hUbyx9xXl3LtFfwGgi3FSy5KkKJJKKIWElSyA+aH/JWX
sCvbK5UziwjtZ6jx3Cuh2rY4u7xuSEWDQOxaEithygVZFxO2WFd2amCQHLGEqyBa
Lz1YAvHmWPHxwgEtklDOFCwpH9hBgXigogr6TZ3WZGqdGiF0TyGXinIPX0+LrhHN
Mrbu66ggw6/ekZI4QEXzIDZJlZVqcNs0XVoIBPXhJRN5ouyKB/NcVMZ8jTJ/qy49
JFBVENgcn/+xVXBzHQCvVhLJ88iRKXjwbO2tHBU1dxBN4B+jYRXKY7bGLheDTeB8
E/2jxFkL++T1IBJp/Zu9tHWiIl9ChgSpR7/4HoqmvnJQfekU35rT51mJqDN3g4qq
MJxyj/a7HfgEGAxxmnzZDbzo6y7UdhozxhSotbxmu3aQNwMjssucnvwe3+Cq3tV4
V7Us7VaelOwMvzNQ0rFfoQKgrrfq129xJohj1TJIUyjjOwDbAp/DFsRQaD6SgctM
9Ff8TrbeRS8YxQoaSjOA8AIs6DwnDaqJNqz8kBWd9EkP7GA+i40UaDiLjmGhkgCI
Azm3uyeLu1TV+gS/OABgzj/FxtzJxuvM+jAYLR/q+DMzUwOl6RQrl3Jh23cQTD7g
wI1TxSW5/0/ziUai54G1qi2m+5pOUNLBZ/YUPmT5gg4ViUKhKIVDOzQLYFrhenEC
Sg1iePJ4mrguTcz3h8h+sJfmrdGrT6k+OZNFzPcnbJ/EhofAsJeyNkmBQxVFWhT5
Zx8wA8SXQHRSi1OSy2Bf+sj08Y1ARMhMgn8bBWUZGinHlKh/Bjlb1aaOxUHu80oE
30A8eNIPKT/yY9Zc4xpyyV7d1SDq0jNmxN1Z8q9/RuVsrfAOA9kGnETrx1WSpjrY
75IosGjrvZPaSvxbMtq8+i9c/CPA+JgpsVN9wae37XjQPkq/cU+VKOq2ODojJJUZ
3Pu7NOE2Q+VdUDeX2XAAJW4eznw37mr9F4kUppIs0d1dgTR/Lf3im/kKuxVNHB/e
teY98vE/ImHQ436WV0qDUoPHuludCLbncw0aShThOFXoOW+2WCNY0sIR3wjytdov
ifYahlI8kcSCAMU/LPAZCoE65T295MGvUv4uj3cjFWCG/n93/yzA7Ycv7dJ68PfU
eDTKJTg96HWsLFqxN73aQgrTjVspvpb9Jgo04cIkbZGwi5b2SEIouNYDwU+Lzicp
gLJIcpobVi1bxYd2T1ERhUd4GKlV3DAlc0u48GmgB5UCj/C7YcBi8XuOSnOz+vZ/
FSTXlIsLSvsa4jMMS6m4MoIbbHR1T5uFiqTu3X9gKE4vF94796hECAeWu60bG21b
6GeeUwoktJgu3tnob8MEM8wyHnfE37zdUxrONzKaP/c=
`pragma protect end_protected
