// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:05:34 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Ix2oxneRx/cw29KiDbD9+B3NtCk//UtkZ3NRo8Pl0Gdu+ThOJRsnC+wxOOjOYngA
DGIxL25J4nkSHiKemnV+d1i+LUFZ8SCsCahqFHW4eP7yBSAEv4NWyKg68Gzh5ERk
IPLq5y8cV7aunwtXbpdIoI27DVSVZO73yTjeArYqyMY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8160)
X/zxrUQbgm9qdRTgzxRp7l+4Quo9Q5Up0h7FPGji9CJq5pmYDGFT1wI91DeP6e4P
MzqHveCrrtLoWPFE7KmRya6WSUrQrJLROiv7xA8/hUNxS+BkeMWRJ5ZuNlYShHZa
TjzgaVvlXUxlg4q3QBnpsc2mBo8b2x6U8DLQ+zKKZ89/xYHe/ZfP9YAqUvDrNm+d
opuvmsv05J1618V43Q4Pt2Zri9wbvtHoabeqdL2iLgQmOL6yMkzw5HRE5cuwMxOx
hyloKTNb/wLtKvfs1ncOPi1MfYOcZ0D6pD7kJJKWPOsTOfp/KRoSrC0ozkdr50TX
49RniLSO2ZxSy/PE9o3Iy9xCAKrREi2TyO3Or4aicbz1oHy6gcKORJ+OWgGctxt1
RpS5ut4nT87h8NYXIITOvjztL3wfWXIu0VH0vGFiz9gKXI8Gy0uOy5HmdLPxphBc
mZKWNlNATmq+iICYIMt4K7I8WonFZSfqeJ6qe2FSfm96K0jehaD5N6Pt3Iv3dLz1
zaKVwLiGpWvoJ8AtT0HqvewkgbGzzukukSuh1ZFVeHFEHRPMIoB8+U+RgN2v9Krz
08c6lLkhmeJdKRChvS9nf1uw7X2MS1buGFoOUQSAK8RSUF8x60HE7q2whap3eKfU
bjrQOXPqAUJdQBt0fiCPibAGJdT+C8K6L3ixY9cAQ5Sb24hlN+L884TlLdMMwyx5
teD2lbHTkDqzAf6e1LoKJ2EVBgP65yK3QQyk3KkBDHbewa7Hx4HqJQNU7+CNiWEb
uVohL8q3zrF69zB4fhoOjF4OE6j/eWPhGKSJWwbJ7VWSWeI96xuE/l53Yr/9tObk
ySgw88g7MWc++pwFiOJVf+EgogL0Dkv0bne2GKBRCdyep+qj+e3vUHdybtSyWB6a
L27LiV1LmmnaqYMNPKWgfzPt0hWa4YaeS36tYcCR0pZYrWNKM33XYooJ2VMVz5ca
5Lu7ksY6zKllX6bM6O8Kc+UdFWhG4GJPKVWZi7ZRmkrQtmHIs33WUAp6bm44RwLN
Ope2XDWSItvMyVpPqoYTSbxVNLXy7X5H10N4h4r7YET7AsNC0vZXOr8/9mDYGKIQ
ycKTYaQR2k/9P9R7l4rtL0kaA3/8E80kcGB8B7XVIDMr+OczW4e5F+HkNoR7T8g5
niyD9jq/0hXZLiOt7NJ50TmGWUoZqd4iy/mE+/hI8qCUOxZ5W0ymnaXs8HKkHQjH
36CR4MFV8tXIW4hpiEmATCyaAiI2QrN0jeRLk1+jiUjDu+dNbXBqh09FcpvgDA8X
XJE/d59D7+EEx03W9OyH9mFOq05B9vTzdR9LvKp+ldVr1p1Oq1xWhYJpyOIreaPU
eAEUqcEBl8IX1DaBk/aVJFSnfRpGbYK6Rr7laWPRS3BNDcn3x4YYD/ES0tugc2SA
kk6BVMMybXrxwrYomoY+GU5gFWcJG3NRJl1Dhz0JA7ZKE/xoUR4FsDXRdhTv7Gck
QWeSIBKyVOhuQWkHxTLKqDoLMBY+481tH+qdtqUoNYYYMHh5jMF3Ind8+HbRTuFb
ALyjj4QJLYpx/kqHiUQ1EiyDnN4mjRDhso2fSDd5fpT4y35iRljC/CEspfB00cuY
und/lXxAm46VHz4GsYM9Fdr07WoATtp2dJSxj3r5eaj1Zu4BPIJGwVDkUdjmygvq
QnxZqt98BbIaLAL/4NrnBnRDzspJRJOWoeNR7oG4Wdjh063Ue1xfp/u609hFUqYq
/TSyqaqcmqc7XzlwbgvEw66eW57E+s/2g0JRT43KqL4Bpz/VG9mn6n9PlDjsZPz3
bnfKQYegQ9B6vmzb2DU5sCUy39gVPq8wP17TJXsCuwlJT1jbEF9IDF2CbZF++0T1
13P2Ab5tpKAzMddRmJs7JoMaH20OdZ7JDJaEpNoqjxFcNKrKrNjsjKWbDKiyMl0n
OkE1/9Si784Xz98PpMXarOALq4kgztPaxeLnBuRxrUh3g1ptlyzPudE7V19w/JAx
E/pP3WNVMeDjfg3g2gmUpcLLa7gJLBDBtvxAeoPE6v41oWMr68oqgoIU3UDX8+wE
QnJgf6rcZuH+ehyY8ln+h9H+fzjmX6lRUjyiOKdzsq+GeBHJaZyLviVPMO9Im5sT
1FOhY/XqykIGDrOXI0LpRev/YCQ/r8AU+IKCITbsl/QHiaBwxBoHDkptSwYthgAV
QJuka4nnXjV6PJG9Db0cW/MSeWkSOo99RQ/Wh8m+TOFssjSObOcv4iqYlMjlEIg3
2vEkD3gf1Bplv8eyVjMel6zstpGKnLFV2Z1ffJxie6pH6vlgDaI2BSjnRFSu8mE0
ktsoPjAuIcxYkcPDIGmNI14vUV//iDoa1i3ohQUtKn92KB02vrzp7KmnTDjwiShc
LzdwvlBdxjc4k1rFCsarJu2FtpdO2n5waIsWrldsCl1WIlBImkUMIo60fwST0AoZ
racB3jKgWHvbYJmQZbcJ54TlVnP5NvSDrVDUP4erD0dHGdbmka63d5aCmuDwBPE7
qX0Kw6H1UbVRTv0wuh4c8WlhNwDx1umoUBsTpCGfSY4GuP5fIxNHtdF8gjUd6bxk
jupWbqAIvdr1z+xXb6Srt390BsTFVcO1ZZcQSt5xBt29DDwR6S4H/I+Ab/qHRuqJ
ro6zsDTBmd9Y/DSyI2Q0M5JXPRvS8K18Mh59Jl3UWtO07iu3YtjMUXN7TUJu4IkZ
iCasY6Hn+JgZLscX4qpNCQNk0zgz3j819L38sGY6LxdeqrZVIbukI6LMZflhhqQo
0dDQJqsB0S/ru+JRGJM7SSw4qjSDZnNZYsd05CDzCDk8f6KDniU9DhDQU/PNuw7c
gJvh2MIvy106Dtggstw+QEeH3dm8kK0zjATo7UHPavLnFVgwB7GYQtcygTXAAO7c
QkthN36iELG+LQnDCtiz5EETiu6qP2Ude3xkNHk5ChNp9MgNg/CwmvzMaHew2iYw
CjWbN4tlOLhSkfdJeGuOtjAf1C48swHj8hq3sPyZPG7NaJiMttWUUpem9SvknI4/
9XizeSrbRCFnQMVpZmtl+Fvn+gJSY1k/9gxaA7dPEuKLR2de57YicBR4tdhXTz8U
MV5u04ZQa+qfdzSDzQclfhxPMTV+0ibEQZQU6kTnk60WomJG2PEJ9cvRTcKFcLU5
lnFlZAacaHLm6rS+Tm0nYOUpL1Q0XzA9DwgJ4VBi2C3vgGae3e7uow5nO9wsoJ12
VmVDojCQ/Eg+rxX6ZxUYm7fjJvsuxxsEhGX3TLv9GtQsveA9JVjlkf4aymzAvB+4
pJ+uOT41Z9aJ21G1jMrjyeyMpu47pJbUsN9TTJM7veofend4LEHzud6+95BSo0WU
2s5KvRyo/WFEZ1H4PFF9UPI49F+17VMstkGfu4+Zd4Js/0mhV1eDwoYc06p3Azdn
LCiV+W4xtRcL6MYwCGP4Qoh1JOztLxMbBfIZRjpcq/XIiXMd5Ot0czjVijNxgxN9
xzwCx2LRiu12PIXVF+JpExVhuUHE9MMKMoMzfdPApDEgXfaQuKzYB9yR2A8lHOGu
qI5wWiERi9Nl2M/rFaMDrLouyrZdTX8uVx6lLeiIUjI+8bU+oA/0qCvHJLJBzq6+
PS0JTgAP/dGqNL1N+G5b83Cr8dBbOkn+A5uEZF/NsXo97raGhczVIjvvMC6088vB
MHBN9le0D+lFnU3v1Pg9YDt+JKs9fg4Rs8p/xzPOQIfyCbei2jolpWFpE2SW0LPf
MTd4Ye2gKsE6o3dvOrUPKNU6S6EJDsgVJp+0Dt6XfGrT183mDQBl09AqDZQwsR2l
4hAan2Ytx5LCblqHa0d/9gie6RGyCuZ6log2e7cIT2lAl4H+tvW2YKX4ON+Uw0Ek
G65Oj08hiIOu2qzlrr0VpYVgtmJmbaZWwG+mtBfnShjBk8ZNkZ9Pi5zGSGLSO+xJ
gf++hIbimah6TltlmcYsiCBKR6IbUWxT6f7bciXaRgMx8RjcT5hoJY3TK43h34Ul
H6t5ip+6vJASQ7Ih3oNnhaXYAry4v+S0SkKsTcWdmiWdKxw9ST9842CjIyaIYhMp
zcAv/l/Ej4WYjQXOBBALRYJyj4f/N1Kh1qGcvm57cb5j/ZWjHf9UaDHUz7JP/0a+
sgipiUf5UnfrpZ0lyY2EanbL3i4CnMe2/RgCVR3svxmGcxpk4y5EWDBuS3QEJB7+
+eVUvm/EbTP1ODIyH4SLs1VHPY0AAgSnU5DHcwNgIB0y8koOgt2b9J4bY6TjBASz
vEeEgDM21bwxnocUbmT9xyY/J8serHXU/wjXqY/V0sHjfiZkKUnGrcRfCfqunNVv
FB+yu7I3LYhF1qtFp2AdpKExqlsxo04SS672OuO82k7fuGSUyBSvEZAkOU1nRXe0
PSQTdGJxlMN3Mij7ZlfYkYqq73LZI96Tego/dENs62M1bFomyhpx3R94d/aO5nzN
HH00SovKKM8+aAcAXxKGr2HdiFRxUeJd6JrzZqOplESD9CJZTDJXF9twjyH5FndR
HTVn3ABYLynV1y14oEtjTicJbxLmFbBx84Dl44n8epVCpo1+alCMJIOp5OmMXCM6
mzr4ofYnbgl7IQnw+0T6NEVvoMBB0p/H/pRb9d+wM/BlclLhWgaDwyOtmzyJvKTF
HSM8yNoyNMupa4jwNC3d8cabLvArhdxrmhoK7/Q1+iiBTguQWWK1I7HCyyRHEIxH
zt5q69tCZ4Ext6ewUvEkweKnFneZzURnDIEsRX1To9M++yHkXNGO9PQnOpx7a3Pn
6XlZ+NO3/0e2+gwpUYFVluF0VT7noN8M860Q+OPLdzz3hCos+amh6potPtE97cA3
0YEF77BTzEBFpBJIQkPIkajudOC2cX2C1JsOwFDzcqlLdCVVWhUMh/pal3mCEH6t
UhDrd2zjdRHYqnV/IgXxNy+dxss3VqD2HGqZ72ACmyvn5IEDHDnXS7UDwj6JbsWw
4lvzodmM/5UjQe0O80eKFQQVqOZrjlKq/OEHD3JiGbtFVtzg3RoNlFM7OkxMpZYB
QZKPgfuZkId2uJso03muW7ueXnfbrIghxJQFZUGK3TtIyWLm9ah84lYEsVYeJbk3
No3SPwOu5a0O/tTn1MyQHOMM4xItDTQX8w4PQhnQ/ralZkIjNM59cKNy/UwulmE3
ioOMcEU6QH+rxAe+YyiJVs5oYmc1+SYgawSIgVZQEnYRn/QnOyDQFxZGSqpfTcnx
iFn7qJnovb/4jLun4dgpLmgTkAzKyNLaQlPpVXqFX4p44nYgvOOd8nkwFWm/UOfR
RBvnLTMqVWZf7jgKcXDdaKzkNapXjnbag6mIwhvdAgoKuPSawHFA3KkLEWy15Jct
Narmo1LXo6xz4LmN+AiL+cmrM4U/O1Jk32yFNVFN655HDC4OF+ura6xDvABAik1a
aU/Q3X9s0dV+GNJ8spC1nTuz3LUeGgAK4JRuD+K7yLfBdMo5Jj206ujNPmj0248d
tq975CHgnV1YiZfmxjAS48stUqslsr+rnVRsXgsAyLBrimOr8kfIBmnBdZO1Kfbr
3qThuPk16Uxl/nePSJANKLQloELqHm07NtnilZadeRh28vqUfUA8ST3mYfkfZzZX
QgLlWVbG/xcWahqO9bPmeDzfVl+0zCBRuWccL+65GMRaTQLBZtHz1Y2SF16dTA6z
b0gxALGwjE/8Fhhl69blYuoY/frscsacUZ+g0b2wIRvKUHdvR6Zx+BYfHdfgYLVC
8CC+OCVKgCb8Weuniz/7jCIye5sooaxYTEzbhleyxckM0POhhXFEChbIhR0yxCGH
RysGN7f63Olj7sHKd0+EqAAhzon1/LRo2TmSr8+wBEi3ToDKTQQ0Ws10DMdnYQ0Z
98b3mBfCLnm4K1KXDrgA1TvqK5nRX6qVAjXc1QD9IwtEU7z56OLU3aGBFNcChE0v
f07aUF7sPNX6lNe1zxXzjIclIJ3scFrwrlaM4YANfoz73wlF2MQzY3MARijG9fPm
j0R/rh/NkoyV4Z/OBjWRqgGW57LOSe5ZQd3gfh50JOdzJ4gF+erQ4L8unWJrfrSK
VCVh5a21K5ZqJpyDQHUwyCbMbW5V5mZ1yPgah+IFz51gHly//RYb91X5B+5IWJhT
J8tAZjQlKNgqk8GEmWXUZm9RQa5GlbnynbR0+O1EiMR4Gqb8B7QsW+eBsyvMDV9d
Vmi791pUwF/UBivQZwqcKmCqlkFhQcaoKxayrd2PBunsjQwh/i4yXRrOjEzcX5s7
t4kGjXAjRhgGKq8TpGMjB5fDFk4rsFbACmAh7/AFJIeSx22f735cUVKQui/ldFXG
gIYLgXgNc4+dnjfKz3qsTvmuS56pTwC1VNobn3SHTxNp+Bt9MGCaSCdtt3dUrAun
Uyat4u+k4uq1O+Jj0EJ4ATjuaefyRJUbRGs/iN6Yl1KthUsRswZH7hCp3CrOC0Qh
EIggcef9b0U1NoYTjPtk5/uRw+6JT3otq+vL++rwm0XDcIqHKDvoLoQjMfRfyJIL
7MClM8iJ6xrVeydIfqHzaDZo2uap8rD4s9iusC1iKoiHdepZaWoTnrgNBKYtuXwA
0HiizA5BVCdwlTx5OAi3mBxdZg8yfmB/5DKvGFBy4GfzpLYfBsXjTeihLlB6qf11
BjS7MCfLY5CNxWbCm/Fy4iGXte8oaXIaDGd5skOJEywDjkJceG2S8IXOjOOWh9sj
a3Gra2XdYDcw7QXigV5t1kbxHKNUnxTxUN3uzA8fk+ayewp+HgbNUUFj43If6jNp
qDIm/t20C7YpiHII9np4aVYp69IvSPL2G6GDIWMsE/v3t1jBdb+PnC9ygj9Ebp+n
ghdLEWihUDRYV/CzoQWwDb9e02azyB4PK2wTbELVhZ4cT7bh9RZoRjH+71Zj4+U2
GrfMCglZsc7y+tY5IyN4zbjxuFUXYFAiO4sg1hU5GkZNZDLv8kekW8J68Y/2k053
FlCkWXgUlBMOZcMFGzh8EwLSLV1bdlnhFLhYUDf/3iBIsh6bM/5emq9+d8zEKR9v
hTSe936n0rNf54Kt1ZV8xGzEOksMzJe3cWZYyekb9ppmRh3V1Rw9Knp8c4ajVvAO
Fat7/YnyQ3xNx4Wztn5F9t02PYE83m7+SdBGBVdGgPWgHaSoNOrhdDUK6Ro+zaQB
Mj57ZEpLFlE8dgC7MWtf1gf1gCIFsJDb2YyRyN27+Mlw7KSNRq9qAAD73ci26ScW
aCUav07EUFJpyN4b/0nG1RWCdbEQCe9E++yXxu5EDlEvPtWEDIrOOHd4DyrZHRdM
rG9Q34InT/cXs6aUDiKbU9h/EN48Cp9/ZgP0PDnAIJUYTnOHdrwA7XG/w5gEC9Y2
E/oXZpm4o7w1GMRAupWzvv69OWpivpheINbXKvOpqG/EU9OoQVLFQr/U7Tq9SNrC
TAhg5ELi6blblIudZO8kABwwkBZZbOl7XWGCw5PnXIuNr1u1d+1JOuSNVAFoR2ep
mGJTneC1LoJHbYmdM7J3T3IiKHt13WGg+5kOViQwQ6m/3VAacKWrnU2x5vkMzwmv
EGxert/mCm7gxov2UP44+CFp49eZrQdO9W+YdVqX3p+LnYiuyVSaAy0eI5yDoMTV
7+rP+TArzbJ+TrHtPI4UUDFAy+yvhfFtHXnwuniVlcjyVTLrWVz0AmOEGaCWf7NM
k3OMKxPR/v24KRirEpzjg8UuQaDWe80e8SNSIPN8Kg4imHsn1w214AyiAB4a9icX
TTE3Tlh2ZuqSUXuvJLTtFYr/Z3ags5ihSUYNIOWe9gWHiWn9rTgKbNyYXf36B+Xr
wIu6h1xtlnld1K22i/e+pEITVTJfds177dZQtuB/LRuf2R6wvMDTYFaBei++97I6
xXvP/VHHfpRN3Rbp0Tyha90OyZ1zGq9kHBaVx2vK7L2dYS0ht7u5ASWbkkZrRxOL
ubGEepw11Y5CevLoIwr8rx0R5fu6co0uAF2kBdTyCZ7u6I04ttP0YlQaygWgMTRA
IST0cwEMaE2G+UJByN8xZA76azVk+1XyLGhfxTrryoEjkgWeqSkkFN3WV8VxaSaT
aU103mR9agOsCAJeck0yP0q66Cr+7HEYKJtzObwJgpS7hxBWQGOYk52MfC4Og7/b
du7cLmP/Mjz8pKR935oHn71EgmXwqUuLHuVIjtlVzUUhkGxjW8gvyJML7hbjAdUV
dLpzdTG48vJwNS/KhV7FQV0IJyuru7iyS62F6yJ5pGvynY+CDYedeIs5RgwrvVlN
oY7LmWESKc3Uw4xUsjbSznValvXrtdgi4DoBFFS/sp1Qi9H5NHVFbI2SQzIrbpTg
C6SrGEU1GiWGArqTMDp2CIn+7mB9SQ0X09hNPXz71m4giThjR+qxBYkva3TtJZFe
7XCwumLgrRySjjysgo2t7WbSCyHOGYLhDkZVoar4W/Q8s7IAorCOIubvP7pDXhuq
NiD220IlQwrcDN6x3O/R0nJ5mgNy0yc0M1sdk5LZd4Rrjs4kiqdOz0H3Pjwgy00W
tGMrXadEjkaYRoD8XfQtHgc9pZ6YP37gbVR9fngdEIhVy3S4Oy3zrVOvk60Sc8up
Feryl5bmvtwG7tCQy5dKyVQMHAs5akLn5U3UJ9+b6HFfUUUaN9PrdOI8qosXloAY
cYel5EGcWK4ctTbvGkxMXlpOne2vY7Lai/sdIapheeyFhL3sO4k1WG18VO7XqMXu
0bPDuEF5OUyErSqF5jULH4nF9yUsc4b0z9M35TJgUFbMHrFOBhQivCFpP5WYYbwG
X0dDBb980V5Wq8aGwFeOrAJUNOTUGCr7y4sXiJ/0vr6Bx89bW14o2lHxBU309oP0
SaRq0KKpwNks/NoiL0kvrdxf287Fwc7K8mM/hKVe0iepdsyn9+iaYvgWoiYbcS0/
6GOhegUUYacwqGvuS6qpFUhTWlBiTTFHsniecFayOIWGp4nGMwRy9nDpSKumC6yk
IHsa4ojnnkTDLnNd3oM9Bxrzw92gq52/ucw7WYVELg6+DzKNw1bEFKlnwiTSd/yU
VGEFdrzC88GOwjS3xbPPTvlrQky6pPn7SV81OHvhWZhJT/Mvuf7NQfEn4QYK7vIw
udnt7TCJMAZRTe2N0CXs+suh3tNrlUntGrQ2lSx88JTxhTp3fdoO42MdAn9yAn7M
+ojDxwliQVCi79ImuiO8bhk+RddV/Z9jsLJZ6lkZT5aVtwmbn1lrvVtxD9CMJVQY
dlt5tW0LkxR+wanaaeJkh2GX3l55P/jPiZ2CUn+hpnOZ4AHaGQTYiaHm92ZaW0VP
DQ+5UYx2FpuBkXg4GPk8jWy3ogt+975suhhkd9nwzoPxQ1pAx/rYeoxaI4hw+Qr4
C/982bxUveMBWt5GDnJZXcVX8wBaoMywmiX57ivkyf4WJ9jHn0P+SGhLfgU0HyoU
6vkAtRMFCkuYVbd00RbyreudIc+Pe7FaUlAD13FyGKfCouu7Us79pl/gXSLBV/9i
oIfJiObitvU8J1szVLSZaaHM6hakDyt4qyTL9Ivtmrc2LK3PB2USs6P+Rlm43bCY
sEtDQUqAPc5NON2m34eM/3rNK134iS3E4DUQmNe+F6d7oHxioGJF2Ejd9hzPmwLx
3eYIfNj3hH1KR9Hb0G0CabPx4xLDz0x06OrkNqX9ijN58tmADo75VGwh6VjBYFqk
8GX7UefKKWYS8Km83dPzWzMU29PeIgjZ5N0J0zoSJHax5Q9//VoqxR2gGzjA7uK1
V+D43um1ePou6867+sBmtClzCGIcubY/Hd/KYHOSW2jMqznMzwLIqfljlstOBPxL
Vj+oqtWnaiY+ezewnAlawsZaebryOW9jJ2TcZ8wPgaGMs8axxcS40jmB3OL0pAEp
ITWFp6o7ISIMhkw0d1VV62AlY6DxLm9jI5E4sWKnISZmdHN/qbndFAVjYoX2/1hz
uzT0cr6NV8+oMcCH7yDEtGrE4V7D8zypfnFeLEzlBNJYjCLF1MJD5vOu5o3FlJ/l
H/DFz/4s5NlbGk9uXLsBZ7AoTQwYT9126zmvqgZGc2L+vQ8pISIMxiyUGSwzVy2V
tNUdJ3EAG0YDChcLi/gAFkbvTpp86zG/5TcOKH0FhyUueRa1s+xNltxjZZB1vw9p
uPek+Yqj0C9I11LA8dS/Y2CqdtKEGJcKvDKOwT+yo/dXQxE+ru1TMOkj/SaInlcu
SsFRnEz3ASpWKon0IMVg1Zh1vNIyCdxvcXy/f2WJ2ibt3Zuih7oMfBKLEu+475eI
s3Ir+D9RNlNgaBds3pg52pgEhTCHFBFldMFapA2i/EWWuGImAM5mMG3jUclfxQQo
fr8/JYdCz6TrkWAUPPKDhuJTnAa6Zw821S2VDCx8SSAvgq7expARMNSFrNEDSx9q
4t1qwP+MR9GrZc1Vwqzt28+R0t1cizztSlOby9zbAh9w/TzAZMtuuQps7SpVk6SL
NtX5woR7R6XvJn9UgQ8mmPXvazIEwRb+SbNkZ5hN3zJR1xIcmbKA6NGM1KeMr6/1
YNkttdIPdvyOiJDAY1FeZEQC8w307PXCT05Y8jiXral6/l6AIpsuiHuE6pQ0HJgX
uTEq6uO8kuOoqEMDgoFlE/Th7AlqGZfAIVgGbzUA9RjUjFZBLl2AsCVUfUyE4GrZ
wPML/3NUcU07R59zhH6m5gLQ9ajYVOHN5Od7bC8vrfGrEVyEq3LB2ftD1Uzs+gKn
Jq8lJMSNMGtg4fNiEdcYE9JjOrRRAozjMzOZf30yLriBgIeol0nf01JAzxYngSRN
+Fa6iCjTOkxdQKdfKnnk/BB6m2gSy+uvSRw7UikArPIXXzP2RrObFvVFXvXGQ16b
anERWnYRwuJLTJZ5ZRd5Am6fsFObra4ZO2QTpaW6d24/VX6Lj9g+L0CiyHw751Nb
Vd9IJSvV3OtaIndLaj01WwKwW+Xf+H0rWOvA2q6FlMV5fpi0K7JwuT9GSljAsqxa
`pragma protect end_protected
