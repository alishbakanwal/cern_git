// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:02:09 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ZNqqrOgJ20sLmvn9RSgDdUJpN3soZd5mvuicl0MZY4yz4m4z6d9VgCh6fcpGAwCB
Ch/Poz3MU/Jif9wq0k/y84x+5KlZgNCvtKcPPuqshNoGrTICyA20EqxIxjnjygbR
1mOGHa8Edg8M5D3T6P7MiwbAu2xaflT0i19a37DKRk0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 12352)
es1pxAqWWWJEklnzeH96QQEFeYMLiOnsPgZeDZO91ibsQM4MGoNCT5cqtEKU0kUW
oWxC3MKjADH5+PT6XolQitTK22qP3i8snGNiWkQ0kq1POeeLEj+EfHNJMZhosOxa
wXulSgBIc71UyK/kjSL9kbhYxylDhQCBXXwOof+6QsyCMlhFU9z0LfB/TTjToFwC
AcvescIE48WpqzLr7geciroLi7VHrJeMINbodY4Owm0QNeaSRkzloohITXUvt07M
SWQN5aISVwS4TpGo0UDbIoDL/Bjo9Sm/Jnqhre7dKA5msJEEhOf03vFP23DhpwQ2
Z860fcIHE+jYNXNs9ji8ckVLu+/AexAbEXz0Cx32dgqRLRd6/0RbKstq7e/Vbxj/
BTHPevxJ9+28NEZoTWWcWiXzBRftETcONClrutd8r1BXXzVojrNNHj+NDFzAJg78
A5lheO99g+UFRcCLPIpui+o+Amls48g+k3FBlA8KivGJAyCNV70Icfw5JUEZ9uUC
oVHAC29QPpMwqAFo/azwVGKRaw/YomGM7LgwhPGwR6pY4EAd9NL1UaPHUHTMEZO9
yFUJAnofCdEd49g/ci3ehjLjb/dOu8ZuByEz+UOkdgh6EFBYmmqgAstKAd5QSaUT
zQugVvgzjpNIOqfq0gNt6ydmLkWtkavQvsfzGSoupW57PzZ6fo4FY78wEBqgasCu
fTXJMC4/6Wt8e0mMA25/VBR9BdFGBUBdzsdorUcnxGy6oy7mFkRnTH/zbTC2N2rf
M+TGJqWga4DVYD+t43s1E6Pg+gCB1lnx9JckwDnJqat5nh/T8hLJCM17Ok++AFAw
6gwwJhY8IhCtSO4+dmSBZlRgOg1KHu29xkjR8/Uy8pspRLNIfX92zMvI4RtWQIsY
3VKDRsNkMB8cmTyClDmctecCBagBKc9AYmDPelTGGrKVEL1qFSrTdx+qBJt7YwMC
iuVeOjHffXI0T+YT4MBmQfqt3n7vbq4qcqhGTizBQOhMGKBjzKmeL0XCOMFb0HHg
G1PRu6uG/jkiaz+jeZ2XlMHRr0JHJUMljdrWd7WEAq/haY+wLCGSQa0bylPxEcoe
VLCyygIEFdlUJFt8sHLuRjz0Xi/HsY140dQThl9Y92Sojv4/jdfKikl1/LcBgGTW
I4rLVhag2L2xB36c8g814JMt/3/B5IyUlLheQ60HkzzlqsyBmQk1ZOXMWT6zjTRc
SHxND03sLQZRyhc5T/6YfsF8CFtmS9xe12iAWiS7wTIDiINfdgtmatXD53umT4Nc
ed2hXdl043bCFxtMT21mglVuvQAyi9T0XxhUnjAM/OOLrNHxAsLEDsQPYSNaepPK
wdntq77kktCxIP7yYUNXHa1tiqI06ho83h8g3ObM4+NLgfDQIwV6EG/iksydEbtO
wfzvb3EJUIGzWS6xkt7zD/zhshoNbULflYmtuTJ6Y8IzSX/pQytYqQSYkYQo2jKW
p2Mi4KDR1kkb5lJXAT21lhIL6HveYFy0Fz8nGn0KyfiVrt4Txy5FbkLaPqeVZKrs
3Rv53VLEObzJQVPhEbPEV0ueF7rnEcTRApBvKwBrgBNv/QPYjHFL78He5BUwyGcO
q3WsrrOnSpnXnUWoN/3twKkLTGWGng5CpVB6UjZYacbTspKgGTZpDwOvFo3bbCkc
Bw/rLp97cRnczehOQEaYcB9n2mYNWVvQSVyre7tu5IUQvX9IYp3NpiiWZR8YFLM3
2+7gSnDlofc+VDgro7hw2ZQ8FiksjVSepwy3nCGeAKNcJorbOGLHia8az9sZhWMC
RoqmN8b72t9Wsh4HhtfIc94usf3uWsitrt0iABOlZ/3jIfwMsyNqmzPbhaHYq+b5
UMGWYAUo6z5u7PzKe86u8R1DgzCZ8zLvop/oW3htO0VKa7WIoDeNWTGDquQ/aTH1
PBUs6w2lSznVg6yrIjUGYaoJD8Huq7c99j1BlcUtjTvgqGkU9JPN29vAS3Xs34e1
H3nLeYjaZL4NiYFqo+zoJ85it7e+zvv1bD2iyfsLdf6IPOO/pWNWUvsx63p7UId3
x1IXDhVhNA7hyYTwdaTA0did5ndF0ARbwjlT0BR6RgWPXTRk0G8AgerrfKKjdzXs
j3g8S0qSuyTxedjMXk1jCvMTUTeU+KYV5oZ7anMya7S3UYjdmy2Hvm3WXLry2vYM
rfH3KuQCSEQ0TfYH3q60QYqKU+PV9NP8kDk9SmcWddOrWo4YgDS9XpPb8mrc3l1b
l/Wtf430N+ixPUoO4B2Jm0GP/lOrG2yTDqsVbfGF3FM2uEv1Uh8hqKou7plCX24k
3DYvZVFwdyg2zgkkUUQPK8YfDs+kVQdl4V78G1y/oo30nrbVK++RAk0A39/re0BN
xpB7wkCGgZwlev4/YVhMtK8iLmpAsBtYVT2bchOQAC39O1lPkP7LvNQhXFc4wQf5
6mxvSa4saATNbf6ehul4n7xWkXwSGbJ7ibldQb1Bl7E/Z4Mh/sFXL9BxJDykcPmd
twMZH7UON+0DIw95sua1Z+rVoEgP2QGoZkv8VU8KMnENw/R5wFgw/F+PvXONayiW
Cj6XOWrTuO8aDzndOEFfCyJ+bkrZCKmLg4Ra6IoRJ4nwCbEYnrrnDEwQQIePL6eg
r/wmngoB+TiQF+wOlm3O6zCPwWK2YRGnh1eIRdF/5Us4UHGrWymPJ0/EN1uaM00W
rFUo/uOoWVtPF4CwqdvK7h3p62HQu2T5bYnjs2DuESuoGaAZUs3MfQmQnnDHu1F8
rTT6rqGLNPP6EiuZH70kd1evA1dBOEZDWvVNljuPYULFEFhqASibsYgm+ncw3sjo
lWuySKbvNFMW0t1/CZuHqQzFWy0yJBNeKnX6OAzXDeZuDKnog+8EtMUiryZCzzMn
pFO35FlTOWJFurJlIRKM/oUpX3lZGmKRo2FK33mXjKPeOJks5+kZ3rcC2OBYUiSr
PNTLHBwWOXYtj04Vtnmn44VpVFc6gBxHqEskyRk2/LpX44grum98riDzxkQVtryc
P9bFD5yQ/k8A5bA1siQ1JQJvbgrSHbaXwEZoyZvTeJ7cQLSs9Y9UOq0Dye3uFcDn
+YasnqrvFODh+NOeLW1xLe5dVn8Tz3kATpW5Y/PAvS6VIkMLcQ6/u5pg08lcwkaS
QRpdzkh30M+7D3b7KevsXl2CVF5hxoXyYvpGxW63Lbj2dlHN1hi0utZl3+NxeGer
Q7CKps85RnrwP9EY7fiQqzKqw5VsFJBFBTbEWpdKaodnJxagWEOgPwMnHPdctfzM
FcjdI1kuiwzjCRCePJUaaTg4aneteT38gZf+DrWUtReIQTLCiO2JC9zV2vM0fHvN
3rVZvtUGlcHIiI8CXOkz04Zcga3+2qH5L+hnw65JUc/nGVgX/KF/L5Sgcg24K21Z
lehD5nZnNTSP863kv0QkVpDB33oNw9+zeRXtbicRE99YjpfskgNZsJpSjc7Z14HO
C+MaUApPXvy+c4Zh+gLDc9VN32perZZv0XC4qOSN/obWTbf6J9C1S/SuDNGNPzRb
6CiGOhEYwvYriKC4fFEJpZ9dW+hraf/M2JI3qOh8vu/nfynUQFcKc5FpjarRpjOd
1/oqoykD9BluxPhanYBBReuXPwAtHQFB3LX0y2h0qY4najxg3JRzh4bQUE9zYt6O
eilJUP3OZQN3N5XFcXK8UIxiqxIw9d9Nr/gadygMt65eF0945mJxdVnSDNiHE9EM
1RPQQJr6SSWPPYpKSYKvIQyE4Lc7tIA9wWcrDzDzioeaUZp/I5gpLdTX8lfxedRj
RsnWjNfqLw8gt2c5P64L0SgZGKvuCx0x/VoZLuaEDsD6+FucTNCu3CEXXaFsZcIl
UstLWN2gnRcYmMi0FYTS1Wv5u5vJhH9X9FPrUcdTQpYcmqnEBf4nJGFsIw18T7Fa
wEzm5BzRqucXk+qGUcjetZL7r6yYdpeROgUjZi5O44+onzdj60uvkH4PqLxNEhY/
yM+rsTdfp12GaN2MlCSlmDebKhz3RxSLA+Mn5EESDKbEggytdhO2Hl3t0FIrvobs
vRcdB0z5SNC2/iKK+gF7RZqrvhd6Di23S1CeAEqnZ36JdRqxtlBb+fLc26XQcByl
8zKOqUjqsCgs/zUPvVpXjPtB+lcxY2gPobFQbbANcnd3Gxbqzlae+uot0sBZ+OOw
W+pA89v2VewsbPEux6pz+hbu5NrSk0cqXBtm+YZzGrmvRgi0CS2OWtNTJDN8besd
1Sj/FFJiKWIAM0l7Yi/0NV2FFOxJqTgW4Eb+SlrwqrxgrHx5AnuDYowERZPl/4OZ
lUDM9PlCrE7lAy6v7JqenAM+5gzMPQZ5zbEeL6GQcUHOIPWxX/Tdv+/9epE8XFu3
3McgQqRLRoO03s/pEA0STzDWWLRi8/b4nhK0Udk6nHVheeQry6NO+kBpF9r2GkEM
su0lGrDVfbgiRf5lT6VOhjuVggQyU9aB9WPpvnf80SD2Z+GN6ECG5bzP0Cqj2G0s
qXsH/V7b7zSkgoyX7BgbNes1/EWHxy18CxkWXK8VTotUihjlyhaN0bPpLlWrwLjz
j0CeEeKzCGITmfMOdBJTLkQMZRkBcb0q6MSqbTjaFebJgC6b+TJFrLRQD9A7fRWt
sJ+boPP1/FTcBowP06hp6qMybDa6FC2gqOEvpVZByxoUV6UncZiOScShtAPG1iSj
9ZYzcbPRSSM/gElJt9ywB0+UMPtRQ4UiaaP3qs4hn69ang1/U5SImIoe//qPOWzv
Kq/1bn66c6wTYPoobuiY1utqgE/Djn9ym9MdLFkdvKa6/IpfrgGw+Wlk4PkvcYve
/XqZHxlZamc5n4B3sngYCVOni0YyTUEfvleYKSmThcEIC3oRNl5uyYjJX3SNAyHf
ADVG4un3FSGZwNepzh8rMD/iBSRY9duBCcWG9pHpcez1K6E5MrqGVmXDD+JtFSty
h+9H/PIIQ4nVU1nvTrtpncO+fbUXK2uqlp6TdXQ+7mCdXB3Z7zGqnDMmI0KBk7dD
oj5yjXpxyWmUYIum7tOuuH+YHuKM1lMeURGvqg1OBpVQoJIb5eQ4LIqF9dSYVgg/
CTf0aVf2ShBIXj+eXcw2fh1X6ilg0KXUqVZAdaGKJpLU1V9uBSFKcjsc96G+fbtB
fSw6TIz8mbnrLVOJ+SG8Y0agrCb7sIyAiiBwXuM3WMJjIUzilQpwoKV0s5giRC3k
B97dxiCqHJ9d2PKMWP9Svt2ybkYvQiEkKcFeQK3BwYBkrW3nNvISt2sYJXad8MCk
PgPtoMyrNylwmNCeZ34jRME5MwSJ5EbEqsN4yKBtuG0CVFavDK2ockFOsqeemVBr
fO/00r88ON4v4P2/OazFOUXdE/8my8SUnGMqWTxIk5B2AkO/99JDAFxUS+9GZe9P
JZRwzLD8IXN52rxlzOEYomyB+cvLO5nCSSOKdW43YVvz7L8JFrUu59/E6Tg2MVac
xrRdWMOv7XLsjgPSRhbKSjx3ghJzr/863Wx2rZacYn+2+IrqdWUHraWPVeV7Hn9g
vO2TFnsPaTd+yL8m9qb5jMXovVFW4vSC3FO+VPqiXxn8lKa24Fjy/duy5QaVfjzh
MmLc5E2QxWZX3VNYdSUDZzGyS6u96gqX3Dw2m6LF4fztm+qc0PGljgavliUUxj9O
U4Uoe1M36uK4dbpvTvxjLWqWzbKrW77x90V4YrEuszgvsfOFdQ8PoEp2wBUwyJJl
J45rl8mT9lTiGB1foc0P0Nl00dca8E3QkSPKnohMFOxsipKx/HNuLo572RVkS+CU
hcBPBEAgKg/ZHJ7VBlY1g4dmacCL4MLJZdNjRh5iQ62+/Z2ODEy+Wa55i3wtcPIt
ZxnZwqoOPAMRwueNfiSu3CO9v+dugcZ1TpJWNgTwT2F7l7PWL7+/Cv7fFCGc8//x
FHlczM7lEv2TFG4CM8FgN+Co2zNRo8svoeydr+rwt93/8vqtZmyeMCnKrfI05T5C
xXblcvhQodl3vJTkSemNpNlkl0AfUD46+A4Fo3GXDzZ0G2W7ILWA2oAkg5JY2K6Q
0QufGLhSJDs5pIBQXidZD7K5T/Wy6KN03FyhJE1yfz4tE1a1qp7envf75WpzuqXe
UgsBrLhQB+Hx8RadRD7sPm0yFovvWT53DIymQ5EjKwprJynEiq3MyL/irakkApjo
rR5niPaBBPXPUOP3FlgtmLe6wQSYeoB56cmhCfO0ybUQGhsckPh+Ekyaq05Sxymh
MMzPd+0q/NAZ1cj1rq5pu37P2noa2r9nfVpQfinkqbTHgdbs0+rNCD/GbItM6VpS
zpzm8YgxPrlZpsQA4Zy5GXC5pOZ1yVZ7PYVRoSTOwJcrMd7yHhHkiuUrECGs1uOa
DjhXl3okajAzhlMTedPK4t5Dz/5tqOSGxSm0WIidQos3BiyLJcFdaQzMrKZZPYky
6SMFj4+HWEzV1YZople3BDxtKNy7AMzmg0sOH6pxJd9pAWUZ7DoQe0lKGr1JX/52
G4BYbqbVH3MEhKEaY5Vrlh8rdBPMG7q8vpgZlIgxx7kviVvQ5xqiBVGpvO9yRRxd
zVlaXkyGlSvynGGck5d3ANMUWDeGg+M3vwstTvSc5y7SYNZKBdsTCnq140yBxCvD
0pXe1KU+ycs7U7wmX+8nbyvtK1KX+Ae0okfnZ7T8cDBO0EdsvrNcSsk8JAu4a+P3
pHlc1nA8s2Ib+BRpig4O16JE+6x5bsmtMuTML24w+xo1gAOnMg+MFmTodd064A4B
E46YWNJGJpIv0L/TzgEjo6D7hE4L6oogtb0T0GMu5wAMvm+5+w2ylJYpap8FOOQQ
WMDYKVKc4zaPuUHg86gwzx/TNOJ+7PMQyTj/2WmhXM8YjFXYR936+PgmKHvviA+4
j1u3Lq6MRLVQ+6dsmA3updQ6PyChvZWK9YVMHRMThbYiey5WRXOiCOysBdQ3F2h+
brPxJula1I8aUl2g0zdIMCDF6FA2plHp1iKp30YyPuIYHtyEEryEq1xfqopdjMlw
wtdDMWT1t4y+uMBHbvlrkQ5jXpxc+wmL+4KtyWwHkU69idr01d0y4AbHspLerNTk
3ubbfjyc1tk1y6k5HnKxuUzvJfgWWrZoPSgSOTcEJitgSDcC2cpZOHvql4wbCKVL
qbEik+eGFzvwcFF13KWBrcfaENfsFULCvncnD+ayukMuVHWd+RPQ6pt3eVnLnO+g
vzQ9/15BP07AxGCMSfSf7JijUEfm/CnTOhA0dI4mk4i9YXj6GC0JSouOb5hxA/q8
x/OBPZCaHYcQ8em4eX4RvmXzs1Oer38Wpme6ugU8B5cU76UVxQNI91HolPrtdn1V
ysSzkPc6JRfuSjYfF8fbMmdAjdNySh1p314ZYol2o9MWzdIw/D9wNQ+4t6b/cDdP
zG0C5a6qQhpE9mfSklxODRRnZS5BTLckgpEQ4H0bZSocbO4zB2iO4tkf/bf3zJi1
tclHKGpFPTtyYpEvUNaRyAXWJ3AY2oYLoxfWG8f4Dln9d5go7NVLmFU5Evos9gAY
3oiYmgIAnXh4Rcr3SiNuSihOT6S5vL7XIfIfY3ek+YG567q5DrkRLy8X/MJjksDp
8h9QedPIGvExNhgFgPhQEAlJIBknW/LK184hV8PwlODDDHERowcM1D+d78nYXYtE
VAHYjdEMzFfA2me80BQ7ucIPTPtbUt7Ph4zEwaDqqhVWIGj7J18feai8a9/ow+Ew
yMElyXwzDpq6IuQ2TMVoO++epKsiPvaIsVmJAPn3zv1LWV0Citnw/JKYy4AEDJIs
/RR48x3Lhe4v+8E2WG0h0lMaBqFcAYQUduTlbJvkPGfnrVA9MRJHyyG+mH4E4uAP
b3k3JJT8NtFuJdGfmhPcZ/3MQlPvBvdp8js+/gr7YcN3ZUrtKo4toakIlLeiOnDA
BOJSR50wx4Pg8uNmS0Nec5b0Yd6bIB4kf9JfdXnGsNlu8Cy2A+6i3m4LsLPyS9ny
rsuxL/OzzUp/oH/JQ117gYJ0Acvqj1zQyRc/5pJOawX8XLpXw6HmBO9DLIJlpWm8
LgfR8y2mw0riMo9EY5xZu94sOMH92Pg7j/UjmciZ57AhZ67vllp5fSMR18ZY3zIC
Bfn4VtDT915BD4UV2JruvrxrstcUHbC2/BRxeQ3BEnwi6qepF/03nasvBco7pkHh
1SDhyBWPm22n4tJccX0bXPuKqm8rtCcZyFe3N/uBH2aMPrvrO6cPADBLX/UoA+/y
wpLHCCYWJZMltOE29cGKE3xLve4IwDVvymypZFmIVOeP2Bkwh+xq4n2SQ4T5cjSe
eQ+f2LcSpISjlRrMCjnOTSTNAzj/iuq/+wRFJLemTlRPR/fOb8LyMD3nQcVtbdV6
QuYwO7QfbEirFBFQOHmVhUGMKmy3wWunb7T6MEJp17vLL/FModZf3EU1x7fQ47Ws
eir2RYakdSpPmktRBpKl4ap6PEZkqnl2HhgCMd19eBTZKN3EaB9bhEvSVKbZcQDC
hrST6fYenpUkY1pvxCUfsoCSBbyypiTOPN2Sn/jll6XBwe73os2+XJSyB14bFgzA
5ivF1bZPDiXgNDSd+SA+c9E3wjfS0Hqi/jPdTmGd9WpIlqju1jBKJ3CkRX24MLPI
OCQkSfsWzmlLuZ06RUSgZe5vfSvSB4FKSCyHWmUewzf8jbm0bxIyxV3L7fWAEI1B
blJxx2lthMSk+eAv384m1BRuHxdVCUqL+OLHV3igbGmw2yqItxi68sv0Dxblp2k/
6x9H6yAxTeLz2URVybZZ+BpA8RSVU/M7JZPSLsRwTvcuO5OodmSWtb8bxLj4TQlO
6iEmGCNU4XiUyozqgS4Dva+YJdAJFaE3IhZ//ieZwHrGX3+Dd1NOmJPK90eP/Hmz
o+eBZBtDKRbz2HGHiIIYFjr6clWAwUpYpNxQniF7YSUVSGpIyzE5KeHvhDRf7eAV
hyZ9/fRli/E5Qx5ZSNrlDaSnXo0L4eAyDSrZnT4311H34gXRP44X/gMuoGLAE1Fc
pPfPGwxgz1HFpfNKHjc6h73FjppXARGdIsr0n9NuIo2e0/zzj8QdqvVg4kkudXfa
UvqCAjF2g+PSHJfS70Aq0qW9OG7MTuqm/LFJh1/MyAdhfQc9g83SLB6R/fxpM0nM
y3y9iU9RTBynAmdiF2NnWOW7eXdwPFUGxt8lg96c2OmRKvJOL0Z5uKIahR09/Ysm
IYJbhBes7fWlk2rz0e2iqIc+r3j3pKL/b7Q3/23IN2dbVlk/kqLLTZfQPsAhep9O
4hWYbU8MnvTuZWMQytfXazQQuwnqcR9KJiAdunlpXVbqkKeVl+06qXfrAX7ld2u8
8N3EzjcNSm4AFH2+OsS+1MAv/LEJRVu5NhlpD4pQfiTzK/C/ouPKo57RKixxESYi
ly9D0ww4mscLFI7Gi8DLWf5LJ0Oq3oskGlvfc8y8dhPEGo5MjiaFx55XYTQF6jBZ
zAsbK0PK0Meb7gZN6X/3qaJ7lQy3T3ezdEPHG64LfFJDc40wgDpMoAs/mTm7fia1
LL7NCy+O/hQMrqNZtdY89LnlY7gb70tktcwzu2yKoJGmDxzFwxN5GhSrqqSsyMwZ
Yn4rZEpI7oD17X7w1lyCGVwxKLnSNKeDoNwymT1nSDxxaAxCR//vPsKGosy/9g8P
ulo/Jmuhs2nFmCcoaVXjadV+igiUKi0OnJh0sB9kQub6xnNKs59vi8uo8kEkHCFD
l/bI/LQof3rlvOc7j8jrr+cFjWmqf02J0gXtXmw89xuSttIG4o9w8VG8o0nFIiD3
CVgAczWYNZnopQyN/ovUgaxYGvg2eEpQ8xeMeN80X3eO7r2hPBUzOoGU1f+RCRP6
Adhehtsd29ZcRgJqNv3nKvLJ/doPnS0lz3kprm+7PwsO340ravq+3brYboiun00k
J62FFfijR9R0p0VyyKUudzz98+X43XTrtv1s05bnvEEUZEPVzUsPiu7u0FB4mFFu
ea62YXM3joOxajZv6OVUMcVG4WQOBU4qRb+3wGOGyPBN0BL4xWMHtRU31Dm8qvUk
HZ+fXc0tnSzgLDJHRzt3M5CB/LpE1amfTIk8pLS8VMwbWCrUSz0In1QpEndpzVF+
vcF1Zb+JajAtYiy6vFw6AzDVzNLuHYvT1SiqlpaaCHxD4tDq7NT1jLFE+9q9xINn
SZ7c9xyx0DT9LyRig4NbR/AoXEwSL+9DCgDYhTpfkTTMLKw6g59Lhh8sjmWOrZul
BRNEfLLxD7nYeKyATIYY0oE8n3GiNRMJtGEzimrHWB7+LHJr8rSB42h4K6HUFxYJ
BOtTmvT65iM5oNJRXG77AQS2N7taVurSmUIc6p2a7aifSCHdL9Lf7g2k03TVoorW
k0D1uHNgEKU2kTuhNPqk5GIHM6YsOKcKvsF6IEH6sO9D4vUDjdMViTeGSvDxyEz2
CYMMuc+qE8BGK8woJbq8XE9wCNVORuQWcoiHo/CUWIEz3b2UFFCzL74m7yNhVetq
HHPEkbWCscC6/C3Q2n+mfa53eEhZ017a/eTAusBusrkFW/y6eo0GTApRVWvSRaNW
nUp6X4R76yshmD/LZ+YeuXPJMwGBZodsbznJKm5XsxbM4YJodnHW4LB6bG1s5xvi
840aZPYr8pEsTCuRsmFFhoOVOc7sfeBoeTUEsXo2y4PFSrn0GY81GSx95Fz/ueyt
edZTfo3bstsTwNDMcpCJ1XD9g8/NphXmhv8ERRjr2d0nAg4og/u/aMURMYXrRd2/
SoGH0Nc+5E45iCKmo5w1nC66Rr8tcCORHPl0aEoZ9aMEVQ1+emg8c+m/Ynsb6Z5Z
Oa9b3FIHlhXv2ATa3xYe2nY2RiNlV0n8HdDBB3xrIW1qedYY44AZcHLkC3r2/X7i
PQikTBcq0hMdV0JQPOSzwnXMCJQFX2v8DUuaKOG7jIHRC2a5vq95fu1ap/WGhe3F
P6Dw2cmizs8SUIJtP1BJvCKf5ix+GnC+iPXvBzvuimdYBQWZYfJGV9+vupYkd2+w
bd1ZpkiNCEgT2LN7mg9OFmvw4Awzyh6OH8lKorS/8WJTsIqxUQuzVFZuBzOjOCwn
CEm+Oo0Wonl/5HkP1D+mLNzpGv7mXDO5VC7zcOXcnVLEnu8SAZknrKe2fpbkf7ZQ
kM0l9gp2fS94+Pm87lMFhFdlmStAUlHpGnV3qDT2FPFdzaUxTZdBhabp5nBhW7EB
n39sVJCnBf/mlDRKmlm+kZKbnA32EWmg6LcGazfb/rRfelXBTrmxWwMkbgpogHww
tpjlAQ36ZQPTTZHFAwQ5T27iLEZbyknFuBHkiXizmWSKgeghOx7Y1Qm+jL04k5Zb
qEkqOn/vgNk4H5QxpxbNH3a8aZFNNrn2a2IlIxJsiPw+IK1uqmSvcLXrTWvDVstg
rohNeYUfvpEsqhpToMvlzhFAEE2JFER1s3H9PnY0N4Wif+4R04LWBJ6/9wrLznqn
uNRRwCUWGjJu5JoOOpAzme2ujyS0qmclBG37d/sePiwNuw7Q/mceUqvVYwodJ3lk
6E5VmErw1H+FBsPVUD6Xyp0XLSyA9zTW1lXvX+uUfLOdmtq/Ol8apX26+KeYkgph
qYwGHeyBShFij9oI4Z0j066w4uIMTVudzzQKPjiPEdPWTPoa++AgpLkgK6boo8aL
mt+ikmugqV98QdkrC3D5FL2ZnrkZnlRNP4fTZHYveCr9oZ2PqIdeQ0OqqQ0/hfga
AIC15HJE3vxYohe0JISomlZ9omobl55eEh5rmkzcq5XZ0VSbV6OYPTNcFVfCk2jW
O9bdqvZjeCnlYjAbYmfOyInrN8J6x4vph4WY30ze7ucmQtNso4IoxHu17XcCAkOM
JZ8mTK0PpFXEqvTDy6LG3i1mUuOaVFcTQEKOObZJRugUbj4dmdQV/yj8+TeS5GRi
CcKdHoyCcNYvpFlHJ2vnOTWcQTvAD4D4Mth7rjJyF4L5Hh6ujBRGhAsB+PpaIAeK
dgPArq6NKzyUU/l7wG+s9xrCicl3Cj1z5j33CRX3xpgupZFcXIu5yQb9NfUyjbCM
z2r7h9Z4lYKBxxIBBn7mERnQ9B3xlOA37JEDk4vt9cjlzbl/C0re1QivMyjdJVka
lAKqlyZqlVyD3jhuT+Qx7VoKe3dXk86JQMH3BNy1Wbdkp6K1gzgpjiD7AEy1MnUC
rCqGXYfChXgqAESB8hofMnR+zkpp0ealnapgZpUlg1+r8/x73HA0yUEg2M6p9gZX
KGZXJPuHUs3yyjubd6bIpXfOuVdkhJQFXc+BMINzPey5gaJXYwy8chI9KulLMu0Y
yp/QRvs4l8HxcwLhgFF8hcq3wtQtGCvksXoJmbupgxtfPdsCL+L7CEdmpn24X3Wj
gQ8J1JJYCCAYu3DksfNjtM7TXk6zD4uxNiP0vH3m+wmUmQzw8hxlT3vWL3Ykj4h+
7c+U8y+2GlISNihBCdEZ82s6O6rPhHiq8TwDI5IGl0gmXYJIoAGSwsZEcnUbUnVB
F3oIW5qLB/sJRMpyNIpTyNpo2jlS7ZHc2DpSLWvjZG0Z09OMbk6U5ONVQE9WGbb/
2OIap9aG5T3i2HXLWP0BK1NyTgdsh6zPxOX61tQG2aMNlu8SRMT7zwx4NHREM/em
yRsR036QuZun1qD2QT/cYoCIxkqnxts+VEXkusdrFb96L8BJh6xbQUjQov84L4BE
DT4DiwFSFDG6bTx8/eQ1RiqoHgiWcdsyInmRaAS1/fTz2S0e98T+vkRncCBlZltY
lqAii7rCtqDEkzNr1GKLowBGjU9aCGTmEV78/YCGT1vLGOIoizZi+Qu6yTC4ZAIs
omA6nRyh18Wg65YUL7VnhFCNyeR0D9HpSC0rt0hSRsEdrWIKzxd/M5ITyp7OffCa
nu2ydlHcbNoeukgTB3mpTMHdOFxFVC/g2pCJAr3pxE1DNARTbDwqIUs1phrHbpZF
YnvhkNdFq2q/B2DoQEsKfkPWYf6lobg17H3tTODXOaKazdCPaFMWt1eaDCO9/wft
7RbNn0E3JfaqfjBLjaq2sR8a8mq/SxOgCdbwVEgtGk+jw+oozTfKU58AEbKauLdk
qIjWKY1Ysyv2MBDFVG/k5l9ZaxiAYBktR18XNbsp0V+EaFRlsam5yExcTAxBC+oc
HNhQvn2ByJJhSExlMSRXjEOR3+j257PDymYT9VHZ0LOPXYffPp+nlYiNZv8MeYlT
IfKJJv+DDuuTO277D5fSueCdyuBXqirSqabJtwrv8Pty3zP5xvxrORY7ByAqmTnp
iBqshZ/8iq4jC+eGnn3e6485IBBT2Mfr3SuvlobN9YErPvUnUprS7hX0KWd7z/mh
WFo9pxQohnafKQpq5AtinJA01SkGjZ0KO1Ygq9uSd5zJ1f91NOpunU8A66eMZAwi
3k59dIjKeHctT0Rwpx5cNsSHguVntlwnM1T57xJeWeaFaXJhFh2QwOh7QSbgygQU
DWOr4Ps2uq1FOp6+/XZSo4mhSvCIsWDGbG+V5+hQ0KIEj4HYJPeawLSlIU8lU0qo
pmfFeQjyekDN46nKm22S6kONdeouPj4X+tmZzjHw6ru4VScFs0BnKjjtZWCTCqcs
pt81RwlDaSjwWO1bve5vYkSVyf00Uy+cFoOMZ4fNky53GE8CL7Xw0h1nSG8JtprW
cREcC6u1BPg6yh9DrD8xXjS0mHDq5xgCJJrisCeFuHaVngsgTPCdSUbe/DMxLaoC
ARg9QdXmmh/tVgVsLnhDd/72lreUPuVKmelitwHgsu/CHRLmyEJ0gPy/yOz8H7H/
DWpm5LBdM0qIwEpdf8HvmRuGD8zOdFc6UgvFbDNN5TBkuQsGIPNX4aqn6FAHlE5M
rASjC9L3eu+26ioxtTRO6oCzSmOe0TlyuMy0FMPP8ZMQ7SBXKJ4tiWKUxX9YGCa/
GLrCfDhUQtajwTryaM2+l80hN4XM+W/uFq74V0ywxR8kFn4QLBRG57B2Rz5LANPN
tqYawwMX/VWcncz3dlKuvbf/yXTSJwPQ8LEAyqTi+dizJgdUHFcKQQVBcOstiZLn
PaQTX2MKiIcOBIoFALKFOPzyBL0KJm9xlsx9O+ScFGXxiX9kixCEvP9H6d68TXJB
/JFAHXy5LsY5+eVDT9V87JuSHd8iwR7U03/6EQBcLqGF7esujWg0rOzxJK0MSeyI
vJDSMX78Ex5VfwxNJwAHXn9z+HOTyQ9FGtbNPZjPdsNNzA69tiELPXR6bnm4Qpi8
raLBCWwMd49LbtXmKlsCLwRbjsETkA8C6C6s7ywD50XYSC4KxNTpp+CwvHXiOlFd
qBW8fx3dXYArWCa6cpJvbOli5BTchWNifU1KnWZG2n+/uxVwTOCPckwYoL6n2u9R
V6b7tuuKtmxOBj1+zalLD0fYMPqnuA6BT5yJJ7HD0oIGpbg15zgRSVwP7RD5MUtj
FGGfoKYwtxnGxj6zx6IJ1McEmL0YB0JV174ileV0ELzsMfsaJftLO5TT2eMxwrN6
EjhOdpEV/KKiDIQcggqXl2qdtSVorrnDEFr8xqnjQvhVvHRv26JSI9OCf1LJVY/W
5rcSqmGNvPdNurFoTo+HoyRXj1VuPnW7V2xO8yiRZ84wXJQq4v8EMvrqTGTgiGl+
lnrfHvx44stFMUylwwRzw+MwsGklxK+7v4XGUIC8IQ/jAbutg9G+TW+b8e/s5QYM
5w4VPWuMNGjcM3aQS6vCw0GiCUhGyamkIQQUxMJmo61mkOR4+544mtXNkhE8FBpI
wXMkOe53Yy9puZzn+GyStGKicGSerUlN8Qz20goWt/V50cOwJ0QC8mf7ukwh4FWr
p9uoi+xnBkcFljaIMGlQr+3M7zwQNyl80CNk++zmkjbn84S2lD0S76xwEs1bD3AW
nJ3spc81v3WT4EwQABnEcJ1IDwcK6TyNtP+WDhwvVlv4Bv3UuCLL+opP+x0y7yfE
3GapR5XEpzWs0jbKNXTFiT88wcQFAxkGrEaU/X/gHbm13pzCHCX2ZI2yPNsWFrl1
oAZAvPDjHNy7P/V9Z2TjPF0PSogofR+5UYRaT9tupngu7PTlH+6xfP17pMpK58r6
wWpF6jj+TmP4AAw+U6IOnLogwnK000zT+BWZwsXAvLbbvZi1hAmYEdqAOOh/T7G5
TbzIhro4zBnWbxxKsN5wWmV+8kqa/Ma362ALxYxfI7UeZ0eGIWMTVKm2lNvozYbq
Y4zf0sPcdpomOE/PeR2MHfE086bSoLRoXfeVkEQAtmEc9AdJSH6X2LzQlBB9aia9
owkA218wwwybT6vbGy3MrsHrfJQbFXsE6glcblETo6GxwpF6saWBe2rAFtVUuxKh
lzFAifoN2hyuUyJjAEQaMg9S5Pg7xvUjqMEjO3bX3qasu3W5Q++HGT8T0He96vI2
jlE1I3aXGgp/4NTjISwybdp8aZUdcWD+/iqw6gQiOvfF4sTVNcbTYoblNLOGnBuN
ZnPN7pfux3AfrvaefKSejefUwB1dmYC0OClE4jVZ6ezagnjgdszXVMu8H4jXkK33
PPa89rr3eShz2cBXaYCR7kHvRsaPsvfpcll8myrpSVoCwm10cWYSegUqY9t7tLdh
jd4OxVFFGtM5jtR5KyY8BlSeuLe/LO8kZVH15E8nJDA0ARhcw9wwb3nJI8sPOePI
eoSa5dy0NDtuvt6s+rvrG/l9k+pBmio4GzRaYBuG03bwIjlLd3sMy5jbVmX2Og1U
NC40TE+AziOX9ymV8AXz0w7Fs2ZB4KkxxsoTD8iAATzOLX9L7jhBaRKn1jGGZgaW
nC4UdJbtVAuyRaq5lY+EESI5dup6/iv/b5m7W7Rjrf7bb1hqB8vB6uy3+OeLpvMo
5XDs7YJF63GYgsC2xHPYnH3hLSp8AchoWgb5ZieTmPiOL6RDqUG30PpBiMaTuLwc
FTeqnPs/wVmk4yF07j5gSrQFMbF6dt8cXftbaStwSK4dpACV6AD7Q5hdzVAuKqXU
OBNVhkiaC0eD1neXx2NeiOC0CHxN8k1U+UrBhFwjrHMenhKafoUW5+BSuZIUO32r
oo+3yu6vrJS63yLtkIsl/XoHSHUDybryQ+jq21P1L9g9IkJ/yg3a3kUDnI7HkX9T
tOpl5NUT0F/v8DH/GcwQuicCKSShV93QVlEAXQsnuPgzXk5YvWTc1kLOfkT5dklA
K6qHLaHwZHtri8EScwTnGUBYnvIb2Izx/LSk0WE2zHjK/Vd2A+rcd6nzyw3Xi29T
hTJP11AOPkr/NiMkr++FcLJbfM2TJnBM7meFrv84AoLZCl/zMs5nNI4BWYW5MHdf
7ok3nvC16Y5DRiCI8QcQxcXNHZyjdWYOL0SFgDKt96O5ky0wKRrrD3ISvL/DZmOH
1Gs19aYw6mt6JraVGWA5wgUqZL418oaip7hOaL7m0cKRGjq+I6u1+JZeb1VcmLH9
2yoodX/gmwwgVQctXwYCVG5pCr1TTn6ulW+Cd74YuPck4szmA4/sONKca5mH/2PY
HRkzQS/USyRQ5J62ypAXH5fMhL6XLMVbW6oWUg7CgFTi/jl4Z1oHYaTsx7og6yFM
0EVoXIU7K5PXuVh34U6zWQ==
`pragma protect end_protected
