// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:05:33 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
IbzCxplyRuIrW1g1NLjJ0JRdy4InMDbGeMBxf7Hb+cGvlGyA+dQf5CaLzSgMg6/u
MCeV0G/uU4Gcihfpji4T3+T8q16OtvWsg6y1G9e2M3vg0sn6gfFyxyKlcfsSFIaJ
JvgAI3NSXsm8Nxe5KX4mCQoaw9QI0LLcqK9Hutudpgs=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 10976)
nmaZt8c855m1oZsfhx5XPHGxKlZhb5OdCzbYFKSBovgy78SdwveBPVF37RIq2ID0
1SPG3hu0O43wc1BjPwmFjyJUXLM+mVNBIMk0X2JGPVq1HyXw+PoxPU4AiJY4ev+7
9cHs2YPG6N6/dftHN7F3/Yxt01q9HisU3SXZdc3P/cNY9sdaQj0UAiFBzqvt4SWW
AeuCqnBOhmddqvilsWZGzLVM0DR+l3HTQjBQwY+Y7La3EEUfxXLoz8KTSZPBEzdd
uB6mt/pFXl+SW+PjcROW1HUarcNLijNEZA7bgMaKwnViswivIrrmn60fNY91eQ+D
vRKHZ9EtHZe/JZONuNKvHgUW9aEbJAVNt/qQE7m3L8rCRRIJUKHN4E8IbTl+34ny
HGwDkhpn4fsITSv7vmHPAAoe55bpWIg6X8+O5Dm1U5byjx+s2sNYrR558iPi7+Wm
BWl97XTJx+YCVKIbU+QCcFvSbsquPlZcBnBt8Dww+Vy0cGtwPzGexLqATMM9b6Vs
4666zNvPqolrApS4BJi7UJIqWxeW13a+nlpv9fuxHqplWO1Ty/x0uC5FuCin5BdW
PAZ4iIRPLoDBcrkQznt0bu/9/VjrTQt/+TneUs41Z2vJNlZ2Rvjg0OyL+BOKiQ1o
9Yw3DsHVXb4OZZ6EmT82pDcYJsqQ2qF6AA26Gg7uy3NMjaCbr8MdTPPuOCTAuC0u
SX4uA92c4dmW+Sl5mJMMVxgujHiJmvdA/SsiuxL4JO/Toa3VFq3F2E8IC31MNKCy
1/vSxr9JN1lznzf57tRqx0mzo6cK/ZLhrG7g1CLy325TAOgYo2WI/8AdSpCQE4vS
V0oqSB3ncua+I9kGUP3BpCH+OuAjMGMi863BZrkqEgTGt5H3yssQcjvl8YTDFnjg
Ws0QPfMRyEcCvv/My+l+cfkmbTPphsXTlKG+LZz9RzE6P9SLks1Zz5yYDR9gPuZL
NjqzVMtu7f/F0EY052fl4dpV/9+UnKK3334SO1cl+wX5lmQH8kL6PrcC6Hal3dNC
0jBwLwcY0oD+svOVY6s8qIhJRFLFs7XMO4FjsV/ENoxo3JaS1RucjbAGNU4ByDLo
56csgQO6hIb3nC4ksYK587OnYddM43VXttq/U8+klsph+rGdB0+5HXfXy5y2SUbE
NsxXX3tIYVCDDml3Oestk8ASn9KU5XEqWZyNGEJPIOaB1Fg4A+RS/dlr2RJhJgc+
m9ai8T5VavhKxsWOL7GWaLq4UgKrFDU3OpOy+S5k7Y4dVN/gsviavsnoW0TK4NNk
b2TftFAkCyP7tDgKOE0tyHRZEvGyrrSRD9TtPTGeXiYIGMcFvY3DwM42JioRye0X
wsA5iMnkxGLWG9CHsOPYlCUV4kO2xHa8SlujOqGU0Ul6ZrwXfSrSlUAreNXCTBD6
eGkM7DJd3gq/zmkNQ8hoj1qbeDQzdaxwQSzSLmcE5ZGH2HOy2C4F5yv1TCRz3vca
fEwBncczum4EQsvGsQn6DwtUuxvs51ftYii9nXKAfWzog3qJgt3DfnWpHaNyHfXK
8hpBJfYUIEepWwZFq+fXbHe5/U/eLxZBsvyUhwJHO7e70u7K45sfSw+ebARzUpXq
Hb8hEy2nL4I1zNw4ysv5LpKuVjhnxA9+teIFZli6TMyptV2dFs63ywz0ZMKQdOWr
MNHwwHg86zc7jVjNsFCEmDVhPJXoFFlbokaaFw4+ZIc03uK1DsXBwSMNkiBpolgc
wnP9uZwPhI8r7igAnoBqfKQ7TMDMKR11j8xXrF0Ay4uDjGhszU34UdK4BTZIlEaR
DLj/+gLIidVB6Qssb5ePemQeSgtXuuf/UQ16f2vDhPkNNWqSFyzrjn1LXNOU/DOs
Jp0i7ZihuZ0J/zcBZl2EbGSaoSmkk+AC4cHMWjjgK/chi31fSg8OroAHvVAdbtoB
4ryEqJCpf7yjanUYhYJjxM34vreHyYK3xlGCfyOo/pJVeB63u4PMrDn3U1qgVnTA
wZCYviIus9mNed/IbIhIrnrxgizxumgtpP9v5GM0KLIbN34BC/N5Q/5I/aWWHKDH
plI7n4NzJII7PHxNecWEcRaZpOxRhsAbsyS7kFVCAyWZrqlEmmwySzo289wHRvq3
juLU5/U4+oTtcQzjsiZi335EIiLjN+Zy3R9xbOGmJa+qC/+IgWigb6qD0apJtDY3
PsrJsIFwwC60/nxiMQMF/Cosg/pjdOvYt9oJWkXeQHQe2ENWLmlZEx2ulrBldyeT
HNEapyjxWL9aNkrxrjxtNZSByqiMaqG+Bih64hKJeN6KhLXA7nm/R4lhgQ/6Pjqj
mRbhfAVFWy0f6Uy+3tP4644TISVWyDic3x9fhBsz1EaTSQWIP6nZt8gH42u8pNEs
VwfU5nmJ71rHmI4i5kWDGZhYLvsEXug/ZENZXXQ3ACf3A5SZj8JHRIMGrNSDLH0V
lUN+a83M2oaDClDKGc6xIyauRlzgEGIDuGN8tHceXm97+pcdGOjoC9EmcMNBARqk
NEqQZN3GNl4f0K5stu5rBTaKH5IjCTwI7NWdrivScimxauTeBdoU0zgNaQ3kIrPc
3/H1DBcBqQX8bvOQxfQjXlJzidJlNRwjyn72GNU4lDQV/uKVp9q+IMS3nE2Zw2UW
o6s4PMS9PmwvdDNenIvkWRskU0ABbtKaKYf92ML9AZHhWrh7pglrPSUwLcezZPL5
8HFTD2DkcXwMF/QaUd36tfUBUO7ZxAg8boReQfT9W3Z/wzWiKIh/pc8vudmTeIUY
MSdrQEeLgp7bpuc/KddY6UIvKyKOrNxreGdvjFpi3U6ff092K52C/Vbu61Ee/9w4
nvTfZRwC7QQ9uW+d2w0qI5CKR5Vi4DetAjLlwQhmUCRw00b2L5l7WkfknSK9XEVz
i5JUsofTpTAR/jGIPfVdLfpaDPvf9MOuCcgEIDCsoOE8iux9L/4D28cJ239Vcx2V
ZLkgz+m8JTC0WpNnzgVA/CWLVUUQRM/VfnFenOspYZ2Qq9jPLz63cvT6fP2C1zLe
J1Tqy3A9nDit/+sAlAI0jqesnNDa8/pKA2qzNwF0g5dP++LxRFtwa3BKiLtL4JAA
CeLSDhAlzjTd2O40TwE/mjlInd7BQhb8ALCFyIylEEA4FSI97JQf/SBOWVTdKH2t
CBeEMQABwPj149aNMV9na3S9Rbija/z+YCY3grm0lPthk21WNN769s1aTSh6uK6J
ZrmNfXPkbfISJQWXQoqRrbL9gp3BeSldILWxgUkHo7CpunCVT+/qKaH2+3FhBYRE
w2W9BBqVcJXsc0dWKXW3kzSZn1e3nt0pb/UOvOUvCutKLFjAROwU6jiQ7ptI9GPj
psKsq2ytRhF+k38d9cyUEm0ImIuiNm00oM7DrlwD+GaMh9dglqY/bTxjAWjxqD+E
47xBO5/dNGE+fOKwxFJTZNNR8VexZGttha/1j9ZWxyNk1Y++OoCcfeoFjpiJfGWA
0CdPLMhd0ZscTrZbZ4HixGYJDdnVk0eDpPrUwMA+c3vlHBLECgV/Sx8ktCM33yMi
rW4Sw4GOYvuKHfs6D7EzpALHbnDnLM2B5VaIyYM8BY+B+oIgB+dr4geAd8WxIYZy
W5I+RWLrgywUiBwKhFdi+0X6zw2y84JVWdSLNbZ4IG8xB5EqEwsQxegkZrghm5e8
N2LMVk9gPxAX+cNjSdSFZwVC+30q+lFzfmVbNXVlVPABkt6+KG3fRZIGoeOGtXWB
lypczlT8evcagFcEsmJ/WgaW8t9vbd9giSz7ID03l6hcpWht8GDkUB5mATqic/B9
mN+U5K5WgQ8p7jOpmUHEKj5GjtUofvUTBgyyQU9hoy1UKsAFkjjqeVZdGgjhFJG+
RU2cSPyPujDBFdrd72+NLVa+IrSs1x0qWI+WOrOvBDhRZb/2wjak00YNouTsydPj
qgjdFZcsimQc37130ByFmHhTFdpBwqXWtGG5PXT58Phag/2hCTJJhAu4qIXup3Fi
xeMK/nj5UlcqhOd7gBqEhvJmdaGOBcZlyTZPLsDZXqnYqGWOiDeM2QyiU68zihtT
IC+JgGoaNbBUUgqc2iF3RfiayzEhGNV1fY/9+QUBV4axbGrx4z1UsuaTRcgBiqfU
WqdJx3DZtD/a/Vc9jA9NTEBnoVz8IB4G0C+XyoRNkgDX3zZj26r/LCDDPU0c+JOC
oUyxkaHuD2cJqrxznfO9lYbqmU4CvuHiHcgmqufQ+O70S9MHEXN6YhmNj8YwdACG
F9txTX2pEHp+qMOcOswfgjN1LbYJFDNxhUIdveG593T3Dv31FmnQ+5tarJZlgwfa
Q9hc9tN611gh7ugBxYSpXujEly9eI6yWur8X9QV/NK+f+fAcJoloiDtHcPNehit9
KXvbbQcu+AWmKP/BPnlw1P8eGiXiy/3z0Uy0RHNuocj9W0BjOOVIVaUXoUi/kA2P
4sC/YNV+qmqJn+EwpvnWZHS278TlfoNvJQW8lEyAjjoz3Yc0chHIJZOS2PPx0+Cl
LhiIqHT7k9hRYnUUxhKqEUbqnrH/S7x8rKa0YB7+2P894VIaHl136V70fq2dJY6Q
Lwzv1pC/NPZQT3G7Dpu9haTFsVTqqMRDFI60wfaJmwA2w89dGwrli/YhiBw7aaLd
fPUWgjSpGurkcsmTtHitwZ1P1y40tSpkH7HK7PFsTq5C6qnRlAMCRg4Xs9rDBy1/
26hZXHhntRWXBn/BfasOkt4ZrQtpJMAi9SZPen5zaJS3gjIIE9ssMPO8EZj4+7/R
+9M2JUGBGexT9WRhnoEfskDgo3s9tF56DnlkrKltsiGbRcvcdN4LjXmX8tsgkixe
em02bqe8cXmwQvfSX3cBg05e7jFVOLSR6hRBzSv+LaoVLG+O2PgHUymnTbvDuAFd
CAonvEwLlR+1kyEuH801cBbNyyHx6ANjWgKF1pRkPxBkiqcM2SH3QebFtM7AZ3Na
MMZKQOcP6FZQcYHYInHna58iVCbUk7MsP7222u1OZyMr8348NvOd3wHmVJDciB+c
nKRRCWxPE/nASC3CkbpwDhQyoWRcWwiD6SmcLS1Ve+tb65lWqrp3XmYFqJ154bCx
qx4PsqlDTWPXd1m7BDEcc1Z/TklRY/YtovBPQz6djoYz5CfJ2zaEF5sGebQJX4sR
2yv3N7aqHdmJz/B5sQIQTKtpNLNh6Kad7OxiLsdEITQ07/RL9C9pzwmZVXMUOejN
wkkDOYkphutQwH8lVRbgM2XcqhVOW12p6QfaSUbZ5BMnyYs5O3bGSNJCX2CJMOFQ
5sZDgZ+j7t1OwBatyh6Bd1PUinF9bicGbNFBCRvun7irLnnxYw5vxsVg7l7lUmbe
so7WdjKbAHPOxTrkWJ5Pz1X4YHY+mhiHlnOwZTM1dS3vicVah9G+87i6hfpBdJFc
vIYzllB16fRUU+21Ms+qDVYu/gcY7csiS8D6MZ1qpuDbSrEQtLBHKdM74w0GhuXA
462LXWZ+AZj43jA4GFVeudvCkwIqQNCYE2cxqXqmxucu/fbKuP3wvzJrHwS74Dgp
3DLorWNWuUcPfE90zoE3P+Ol+zKBSXM8poZSEhe8XAib0x4Ig0MGn/n9SBuR2++d
W4n8CMdNWc83HEHPYUfDSvTXYiYbVnYAGoSI67E/Kl1dICyAMkwdQF3bLksGlmZv
vF84E75lsEygxSQ63ln2ExIr/tbulPnVEqBPdMF2o08G7xASJZDbAecHP8ZL4dnW
FsEO9vjtkjMfrX6hle2dje0hCwHrW4kH0RlReCKujxqbmyVqnVIBqOTLk9uYpQir
ZlibZHQN0/685W0gv9glidbP4EMdKsYgB9n0N0h3feoF0CTe6v6a8JIBQLYibIUU
qTUT12u+CwiGMuRJW2iHJLXcD5Rc1YBzsLa90GT+UHkgm4myofFdK1A2oqjeNVtm
Mwg3ASaokLBifG3qhNF6auz1eiPym9Qg2bO790DZG3f/MfICF3iATf54zcH/+Izy
KtrXCrYXuMPbMDcJ5dFhnNPbOgJoy+2Y/BvXMux9wYlqhUENaQxnTlajNgS/+1ES
WoIi6TEEXsM6phUOs9UB5AZhq1WIVEiwnZnxnhhcX0j37U149FpLVfToVyHA3/WB
yLZ1qhx8UJNNGGLJeZqwzaoC6YJDms0Hm6zk3gwTWdxAKg86tbQIjZrnODwramoH
J/zD4dQIkPW15Boe9Z1KKQsm1YhPVZ1urdA01R4Z8gDs1ov6ydBX0zOXDKrAP57D
p3edxOw5sdFevkPWVYAhaScVCnvQkDHu4i+rxsHajGdyiAHL0PrGmk5AMk/1oCi0
moqMYQyQYQCMjeYEBYmxNi4+RGRN+E++aYCQirN09EZdiesTKGNmxesRwqDZ3I7c
oOFf4RO8Ph/Q6BkqWYSjpFv8hRSyhEvmhoVOhlygpyo1Tu/AmrQVCkaAe+eRH9lL
R7LiO8ZypwN0x6az9qUN9uYG1SIpYdhS02HAYhQncqYmVQZTmAt6muU4iaIDSMbB
mK3D5mooyUlz319nBE9ts3v7P+PudPxSHAN1BffhtF3NJ3SAfaeeQKjMoYtXYMWF
Tn6S29m8qCpzG/od5O7TvKRFkfPbPdKolrPtpVDXCD7VzlBSb8ZtZrgxij+p4Tvg
qKk5r2FTz5C3IJYic0kIIpKKVBp6/HaCMkSh+1S8GXdhF0hu54wtNHWW65G7wiy0
+inkhYIA5S309PiEQepTwtWit3ru5FAtKnx2wIhlXa8FWJEy2tp21cWACVZft1SM
4Rh8lomfg3Uw839Ec5c/SHvpMjo14g57mtt2iyIzzrssLJX0Ig2DbOalOJQvID/c
6RunxPC7UrKLaCSIlAW/UVWDdslzkuGy4DEpZHzhMDfaBfwis4sBINcrY87z/9aK
ceu6HscHX3ecoCNsFg19VLeI8sudUr7/METs0dW7RsbppQUtCAwv31ZC44JLhge3
C5/xN6ujzQauaor4lbQNqvP0blemeea6RAua7WSA31Xzi2QucgmNjhmv1BQMAOsX
AXgUvZl7anKxbJnFTRiej5r8MXyF+BT02meodo1u6neXzkD27Et3HVkjGL/C2nQ2
zapAxiP9t7+Ef2moF4u8SnAzm7u/e6ewebGtwqLY6p/WM7F7ntQ2eFLVB18FnYc/
10i1m9vOec4N4K0q7fpMTItbM3/xCDmmG17eTx1qz2Hl+ouixiep1jx68DJH+0tY
qDBmLCOiQOmKyL30ZCto3AOS3S3tZ7Oe/ezfE5R03zPMDrUzZqN+ga7/KNCMdJ6U
MZFngANdzmhM3UyWlr+u+wGJY0gAc6/l51jTB2ijThXENsNOwCyn2+KudUOhqOVU
qRXyT4YyGVRb30a+uT4ST8gqIMJDX8q+W4N7ai2cuo0ikczbgcJ41ExI62qkT2iV
snyquxZMHW8Z6LO0en395lL4JPB663yntYLjIwGkSHk1TwGyrTlZh8abosB2Rap6
9m2v4gNvsze0s9T7p0JEpH4nkobo2ZA0GzKYrVcfT8CklGCslixWmaUAZ6C0jxHT
J+C68JRsvTNJVmkhaU5r6T8QADqLPnFqvLQKFyYqzr2D3SFfJp4cJivMaqdc9W1b
MGUfvtfZ2Qt0xZd7Jzwzys3IdQR+0yb5i7Ak6EYJulkpjdkfe/7LOBbUhkDE+JSi
nQnK26HyNbD7/C53hKNtRUZhsMJZ+Jo2nsF8WbBnJkErwi/Vdm39zhwfpr7kpHFK
AgkrQDYrV1F4dfjnrmf0FnejGt9kxL+2FGIEq2YpdeW6ODrBwWwQyM8u08GklYHE
7kMa32K9OxqPPpFhAdw8NiYPXloes0hGa9Twf2JQI3+A3GiNAJCMrC0sqmQQuohM
HSlFPXY4ll6tcTFRQYppYgCjQ0g5U149QXe1fWp8OWb16ldghZQ2DXwcxWZrbBby
KpQr2P1rm4TrzYxbHTyLeBm0M36paF+qCN9ORZUEG2zXhzVAK2Y2BjbTUol2o5GN
RBz7ZkRXjiiJlCwFcQviy55/Vfz38r1hFxh4Hah6Av2+7GAHRE13EZaQxbJOToTz
SLR/OGCBNOD9h9rVQcwzWnlpV0PNQdQjj7serf24HIKobq3g9jR4NkkMYcSPhXk1
SSVsEOqiTJpkTZuCD2ToxSxXo/fqBO9AfcE0v3dzYLMfhGCbouXhgIHSUyG9Aqhc
FovN9aWDN/scwPAgdyj3jMBU5ktb3X5btzyxOb3VxFU3evtvzd3vd1kIUReSeS8o
0Q+kYCse0KJ5ndUWazXm5qipjgBq3NSVmHp379N/yPHCu6KkDSOHzUcaUj8u/Q/E
RLlbVS0B4zM6uALIrDMmPo+iBybJbJ7MG2RVX9cOV7cdSM4z/0si1w8mJubUHDSq
66g8ySC4llVnhI8ey33k+9ddifhJW+BPwFXvmC5zKDfSikzDmtZEho6+ASQtl8x7
DYFjWvkaH2gKGut5szkB484VSFUQQH2Tm59N8DoSKEeACUIVa0sUHeOIRszdCTdj
bXMI2JXhFqiEGHpLi/WxAgp0kMVj6HM2V0aPFmdeLvqCBQ6QzzZPsjD08nVA23tg
5b+W4N0zllSBI6DgBFWJZdWVgdyvKCQSlBrSpXx+ALP7QOKqEWAvr81sRUzDi5ib
XKwrHGNufr9+vpw0em4NvYVYVu4FsJJI4JXdeUFOoSSxjS01eiTNbFxAZosC1QdJ
5y02Ibx6TXCF4slKiXc2YG4+GlV4qKZuFfEWoXohk17I7oYOfEa/n90AY34gUp2B
Ahg1up6lG6wwLcoupW3JAPm2+qaBuTbiZDC0AlsqpXwMyG/fIlwunZ09HxjUZFEY
DmupcHlJkU/35q7+HYRQsNtTGmYV159jpebsZkzEdllK9ab6j3EEpU4OMCMP1tnW
MnKVB6M0GlIfDXl9FHYT5QXA3bbbxPf/YSPSzYCAauw3+w/XKwZ8Wi6/mo2bLxzn
EqXatBHDtkNhpGVc/ZafIfq/6nBpMHsYyfoJCvudHC2y20FKt2io8F7M8MgMclyd
4eILC8+onjuxSnq1K3yyth/S0T1z+V8xVquTbTdzwipY43WeXHHhNSAvsfb6yqyU
yhxr/KX3sy/DNcV4HAKx9+hyrsHR9R5nbOcQJ5JUEHlwOmgtSWpgO2hYyDZNUjTr
7YLL6kbO9RV5q3F2ayPh1UQwd81VNTbH+WHgrEFskjg9k6HtUbryPYrvYqlru0ih
dhrYuqVAHXqLt44by1aofVMLqgUZ/k4k4wIGyAqeaeu0BfXev93zAOgRg97bRlLt
RFz0hn3Zt1Gz50hLDzm2cw7X/ZBjfwHqpkPjxZManLT5NOw9DPQoXazKeRGUkt7m
uMUKvTnSbNcFRY1gbOyJeh0dgDgvmKG7H/OcV+mr22y5xlHyu3L7XuUqTBVoGq0T
vMdc7XzecUvR+fh0hTVYz6mPunYaoAy4pLGZSNtyQbFtE8koQ+NgSxCng8+unUQS
6jnJCXx3jfSYCdxaOiyNJt3szkP09hQEo2iBqxw5uiDcFPwBysiW4erNgJ5G/YRE
NDXDkvUSck82enFG9/ykpy0OBVu722QuLhiw+dU1GtyZM0PhBU7p65hvdlmIdBYD
KwTKBO83LB3KbZXor6TKu2HqhxVOnqOyUJ8Qv/gumFrs/fBQogHAqj7SB0uekKPZ
iS7qPhWkGIBor8nzZ64Js3dwQMk7jzcYXlUBerXKlO7299jCConsO26/LekFR9d4
e34TMWh9ArY2F+Ma0uWkYvURZJIri5fZ+EJrSTQgG9ptyAOF+/UEcoCte8WWB+Ys
wmd/etp9Kq46wExX1IQCKAVzi7dPoBIIQJuIMe5Yy2lMkjXw7NnqymWbGl4A/Sgs
toEdfiezE5I0guxQxBGZTcaxiIwywJ1yJfMwqeJrx/xJy3xO/0vUniUu9hTE3Ogi
y7Zsw+Rahkw5MpwmTTjsEUbiaFNHIIgbJr2bAlLVBtKZ3l23+5eGEfYJCRbVi95S
Feu2AJ7Mac5FLda9ZrJuejDjchASQyaAJ5EXx+JwHLuLIJXQRZvUM/RGVPMHKIK2
oH/LrWu5GzJRK/D/3TZJizBv9j7ujHPKknkBANgLDNF+CvvZvdFdfCm1kC9IJi2A
2jNA68jsE6EUlHd4vtHwu9PelBZN7Tv8F+N9xQwiDVo8gWPwV0dujB1+alGWd78O
oEQwjr0KLQbDfY/QIEW52BShpO+dRrxKFt7Q/TONVIT/9IIEMQ1sqaeQhT3ZpGHx
d5HVRT4Z0ApE4tOc55I/ePMZi0KtySutveDB/sWrJisqqr6Y8wliI5Lsy9NBwBAq
i5s9tzMGdy4ZunNfeJPSwESEHs/byTGfKYhS/dmtdouJcywq2K7VT3arPYW1P27V
d7xGPLZrJCOxpDPZTuEzbeOpvVKFDEy7w8ouwjXOXwUPBBf5513nY8N+wjh5JHmn
2KkJfGWc1/CN1shZS+mW9nrMhkAS1fzcvMgnFcVJecNhbggPpkyW8LJrT0uoEG5L
IOjAmwaHF0Bu/lZo60D3oEzCX3f6rLT4aFWje6NtT1X2PI4DfRXylbXQhO+9Xk6A
OYK8BTasoSuw2V2u/BO4A20rgPkzzH6d3NqEK9HWVfL23fuULOpR5Q9mxzqU4zGU
XngNgCLSnOndUWVYSgkhpS2dbxmmOj/oM+NgJGdNnPV4jZGw3LPUjR4jP76+0tVh
Ysy4aig8004Ho5cIM44fBiwqMWtpthJ182Phe661u44Ooro6C+2+Gmn2DnhkBTZ/
Fh8gwTYTuU6igIgdykdhYvmHuyIf2nRCsKOqNAoCMa9euE9FdTMwLGMpiZHrrIsQ
vslxWv3hDzscTwZbRJCBRNCRMQiyZhlKo0T8libfo6haKE5pMvYEu5AyFgdgKQcU
8U/7+CVPTfNq7XTB8ktYM7233sgS5LnvyX9Y5v9n/ZZa/ps2gafYe33WE92qElYi
hO2UQZ0y1t6sRE5aGqZy/MQtge28BZrYjNFBhn0h4j8LFFwT6BQwNFzaPD6KQ/IO
t+RqN2k7eK/Ktt9FlhpkryivHmS2dRYBG0FqdYAe4+ApgP9LYQl9SDFkDBDVlmkI
SzDYv10hAM5jJJgI/3StqUzXraFwFZ0zrqVdT2PC2DbbEjQJiHW9Q4jwY7BW0P0T
cczMHeGc9MFLZUNg1fsjBJwrXRhMa68JvEPCmd3nYWkfdYYif+visq7sVz8ZVxXJ
CXmbbEGAXJscxiC15Dvt1xjfjsMCPPIIEa2lFaRKpFaRQFAomS21rIkBEg6aqe15
4Iswscs+KxfGgWQhuU7eqj8YZNYh604vlzx+7HRIRgw72dWvn6mbVjQ/P+ArBvRE
8FCqzqXZFAP/AI9gRQ9sxm84qR6v027i/lU41f04n5WeZSf0kanzvpw29Di+Vckr
/QB5GuKuH8DowZxp+7daJVqakx5TMhfpM8lOmbt1WmCl5qHUc7Vi4D8exW2pQ9O3
Gwzlj9aj8ZXcV1fKnZLhaYEV4QFd6S2wfruS/zY5uESi7G9yKX/64j0MfXTNWNgX
mWc3OCKh+PsZO2flxXJuGc4bNj/0V4+ZtuMtUB50cmNF6jEiDnrTA1/w8ZZlpSz1
9CRsp2M9eyqHLzpO7yWg8rdYsWy/Gt1QESqQZbXYu7/AgIhc0rkkiY1NG3qPjl4O
228uihmmEn3jgqO99bvb5QNE5l42Fu72uvFTU/WHoMkWH6MXL8XLyX41feBJYRvw
Yf6Orv+jdToI1kD+64MeYm805/wWY4K9feWlUxuEUyFwbuVQcOv4AIcITdB1hXKX
VdsASUTiaZd88yKj5feCvJ8CmKsjSEbSxA/RsIWMGONRUOZXj6P9p/kCJYACNWE2
h4PXckZkWs+h+wsGO6gbI6/q0rQXxMHRMzS0MWi/HCy1s91Vp0NJlMM+WuODoPde
R8zCWBA4sub04vtC+r82oLtpj0SkPluqkybsjX6sZN4AqmqqKi/J+GlHMHnlcOBS
lRMPBNFxT12MZoE0ioyS71oDD6+n30g11yH++JrHWe0sC3GKQAizGc+7u3QX7mRO
fcNXH6mVE7yud55F7tMw57JFbpZaSmTb8ZuE1/3aD+LZfZettY2vbVH72x2pYUQv
2Ea+xte1vA+jyXbvKkN/kXmzDdxAdhBywzyA00zfHKo5oiSxetXHUlsxg8LyCrp6
dn9j9RMeSeAjPm4otliQUz5xaHjn6eoTn43ibm1YLJA1Kcb2joA2Rhgh79mKI9yY
wYZSK3BE0i4aH2X/tBtLaCKyMJCXGLJ6H+79ZckMRzjuEg/4bOsNmDi6EHre5l79
6YaOh/ANsZtXlpCVZslBf/j2YDyr6CHiAODVhXIdJyD3yRfDv3Gly7AcEWBiJBrr
35K12mZG1S6n2uEMaE2+71W7Dvyhg+F1vsErbt/tIz2FdlEAaCXECshNuIi3uhZA
yZMAY883lUYZCTpZT71yNyFOx5GIEbjDIBzW0+1veatclPfj/pLsQVL4Jg/sbUNk
8L3O4ACbtlLqBZEJhpkNnBtrIPU1LM6xOsBWMn8AnO5qxnaH8bBaZP9xllQW86bJ
J1+z5QgnlKNNGwpnTH4+lN2QjGirhfoS6zGi907Fu6r7qhGsSPQuuv4mtSbZCWqx
p+zwsegshNC7iV7GDKJKtqXhvs4LIc3mEjA16/nPueLxV3x32/cQghvUCrxWPzl2
4oASSQEYWVbl/VRqLFcBcUWBLHOrfD+RGZEjdUnph2NYEV3lS8J0NuCHzBfiL6nH
9Yuao0elhoV5FfoVTq8L0i4fzdl4lWcR2XQgXG038duJ73A4d/rJiDPjlh/0OjCj
X5vM+iGQIVGLFPhRPPKyuAuCjaKml2FnRxuktM/+El4XvWxOE9tP4zZR3He4bq8X
jVF/DCWJKH/KO7x0egNZeXRhOKnsCiVkkpcGP4Y/e5TsvRDyRt/nWnJeTfaWRCmN
shSZlcm06Esb2/SVmkMldq+7LjaPQW6SszVADRjNSxfW7yidOqq2mWkKiaQ1Ihop
HkUAQ5vVEbHAGBTdwyhisXlDWcROxkDvSRvKJLVOfrpuInKIT/utLdOoe99lLKMU
Hrcq1gR11e3gN6ySjpJol4/XhDgpaSbOgx5n2HsTJqF33T6t525gBrKHhtOVZ9L+
s8g4i0pW6/nhmnceMAMeiquYTGHElD6AHEeCmLg0+Oc+xOBR2U6dQHU74V83n4li
Xu4lTYO8Pn2Ng0b7SCBrwV67sZFVMtcrlC0Ak247tI+nbTDCQ/lHTDLzO7oG9GQE
Qb85n5dbv+eDB6rTEx/Kyj0+wkDLBnJSu/iRyCtfYsCl2w2DcVhuioi6wVeF61zq
pnsB7N4yc/jf3bJ9uM/p/fnEtdN17EKFGoriMMjFQ0IzcjNfdSKUMFz5mh4t9OKk
hnGp/IVb1TkbI42GE7eFO+Yh0x6iAzm19w/5OGM7Xb5M0ZOqlo45wf00p/1+EoHo
usvbLwkjoAF+4VisLfhKFKy31b8gCFMRCTfnZP6VZEp60wR8o3XqJ2Q65wHXt/uI
+lLi2Nk1RZlWEviFG9BE7HxWiH634jfo2f0NWmU2yb4SFxmqCg91SYKEnkgbLxEm
aMtaCpsWk1XU3S1I4oHbMjAULALAwKGShcFshrWuxF3AP5KMQQNtzEqsz4ad5T55
ZDDucPZ9ik5c8932QjSVU2SDsOaWnZXpUSCVJzVKI+0gpHtIYGEZfBgtGqixjbto
jTH3GYzS6eiJbF3TWCm7kjGsRWGI+EaHnBaj+lmjRy6OUy9opgQRbekqY9a6h2rC
3znVEc8iaYEfpW93AQy5ebF5TdSizUdpPuGCU/bg3w3XohfTcxoMYhSLUnmrw/vZ
v8OAa86dT4GWBll3QmWFfJN6kuJ+OR6wyFOrsSqiyXLZl0L+LwOcbnIku45LGiEZ
BJrtYiTS+kQmT2xMu9NksoO7l+TxDZVQ9sBw2pa39wEiFUlxvH/8zOYEW3+anDUB
Z6ug0IUidsp3RnJc2xQ69RpHy24Rd5ccF6ObD3bmDF9o4SMhKBY9sILfx6gsDwT0
it5IHbrmVcePDJELJ38GTrK1cvlBdxGPUJk2vKt+ZYJ2cBye87LYL44VQcn49Wl5
1j7QSER/NiNOScK95wmkc+y3ef9vyNG4Aw6ZqLU1igAuUv4CJhUo8/szYymzD+rR
j216X3D6acK5W59gBENSmmzcSoQ9VSuIT8tIJj/MpHLiFnEb8DvKnpP1AX2aKrqY
59QR1SKeB+1o+4ZmaRatec/zeIk9YXEV8NPLu6tbUdkObNbdlcsvCrqPjQV7u9cl
8x0z9sCngxF5Tx1yDxYsSCZMINTtEp8Dikh2s6tuUopG5/ydWh1kTuv6tSUzDQdF
9ODT3sA2KRbybgbwd1W95rL8Yndt+0fRYqwySjeDymsAsuQ2uKVvPnE/KVJZuVgV
75WkPsYMGUPA7RItavLg8eHElqpHOqm65UpgSOaL4yM5Sks0EAB/QnlgmBdC5tfE
XVKIWM9wrDWMcelra3zMLhOfW6L9Pzowf9wv6hoB6ztUvohHGJx1YVO7jailH5Sj
RbvWlZRsn/oRhR4Zns5sjYC+3yR65uWt/n6/O0gKvx4kjYNRCPtGM9J9mJiOaTgY
QlS53I3TSpnAyAH6wdULIhumbeqRM6sELEIRHyT2cpheC0DzmHDiRrp3Dl1XrsD9
xaNQJ2u+2bdjFdytQ7rvKsSuH6zImZuZPbfR3XdWebI=
`pragma protect end_protected
