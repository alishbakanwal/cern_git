// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:02:17 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
l6tr32RmLuGwf+ApL/4uUczZr6si6RKqguu2ccYJa4vLMCg30I+s26AxLdriv9PQ
9spfwCxl0EMwmMlmmTNCGk10rTak4WxzR0TkXQGfnz0jjIainGXhZJ6ZXY+V4mwj
oBXtnn7PvEehxhqwTSv4Dmn+/cnZsZc3CwnKH6WQ2V4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 20352)
5v9CQuuql2GkCQ/AQYD+LkpA5HHB9PYcqG2+Q4rrjt9OPwdfNFtwyxRXgSwkLFhQ
LqQaocofyzyXCa+AKfbt2XkZosXoapWNLoPqvQUxXJvzuz8dh15Qe1DTjbjJlGLe
T3sjggGxuDDburFSEPklFu8jLVVaiJC0sV/T6oApnuunxuYH/Y7RNyHqyYeg6jkU
sy/52MWpasR9gad4kL+itwsy7J5Ys7b3pO6vfmXnGVjjb4Pvr0bxKSrS6FAcR0UV
cBXN47fD+jZi4p62qjRlMUhE1XRh+PTipWFTiMGtUwe5477JXfpkLfHYFeScfkwW
I0Doct3/QBgJROX0MV8LYL2KNkl8gYZqbZTEiI/yqdq4skbAwlQPjBAZxP0sxrKx
IEqWzQYWaD89NPgtsResbp2yodycavA9yz96AxWUfNZ3bouF5PsuTDPldmyVPZkZ
nk81Ned2bkWHePNImmE1wGhLGxWTzSROkp7QqPB/CeOmaa4j8oRqsPXcxSrXVSqi
646K+WfdYK88+PLM/ueV1IPyZt1//tzAHQVsvp96tsBf7iWfRVMf4UoPrEEFTV/r
RE3U8k0ecckgqbJch/m2LUXEGfgcJpr9vBObN7S9js0KFJ7g0uLv6w+RGcEurC3u
Lei4EAwVU3l8lJnYfQ+7NQ67hKv2ziGnq6/K8Mok/B7ElUJd1Jeev4gq3KLgLXXy
fsWQrJ54rs2WbqUZQAZPkm+bR5sUKlkQ/uFoefz6gtOrcbRRtXFVuJdgrLxj7SXR
SZIuukjMbyHr++MuNzDxKhVsUvFPg3tjw6chX5I4W89VOQNaR1U1lulkomvwbNDl
id7dxTPV+2Tt8lV0UBNGScLnbxjxRxOOxTDxtotSlC/bYHTW35UqSpZEkelXmZJD
Z9OMt8z2eIbOnvv5D3gjAcVD+LKQ+xNotEaJSVyqqQ5dX17F39rsUcTfyp+gxMxP
x0umiz+RrIfr6x/IOPm3cyWOlVPwrG5BC5/+M8POEdwR2QyW/ni/Lw2FMb4LDmXr
RxadCM/T/ciCmJn+4ZB06Ib4Je4T4aVa/tkQxBlRRE8Yzd4/m+ZiWDbffOgI4tRX
PDRGk3uiEQmNkCvgmwiYJaXehrT+LKaFml9QycS0hIH+qX2RyxCp85ZmeVDGVOHq
Ivs01lPqKToC2Fa9Kp9RlVi/9KlB3f2f/eM3FeUPO8PKDJdog6zIiDo5mzFjmoiZ
jIsbZAMCkoBfQ4fR1rj2LTQw/gOg7Hvyb6IjLM5JLJZL473D46LleOC6c5PQBnFQ
400H0ssUXYIh+8QUfJ2vBNVDtqNHxPIhspvosOiYyKABH0YAtauDi+vBDK9EAZrz
ou/0/XyrdLKd4INCxm3srMwgDQfDJ52VePxJwX67uMIITNLwjwLQ1735gqEiMqVV
jYgA/3h6aQbpP971a//vcqLHhyabR/n6Il2V+xbj6JuqVXosuQr10//mMbrHQZtZ
Ib4PPsC8ex/ftEYM43weola/6K0pGrDYIQIMh3qP4rDPFJ5fK8rn/hcMkWitL76O
Lkqmv5RsoYd7oIHZ2fbRmHpYnV9JUP2irBkrddZEu2uNgtPs45Uil7XIpr6V40xj
hXAvVf5Et1oUNybCyIQ46BFE23k4WH3nmpeUJTTtr4uRYHdH/9/yDr0hI7fRElkT
qQ98lSeDWZZ7kDJCWPnlIoWbEF2EwAlxeEZgh35xFVa0onOsi/pVrsUKeNE03Wmb
vWwqzHtRhpn96qNpGhZWhPOmdO4W6yWTAJzHsu73qQpOBlK7IE+aaNEEVd88biCg
hKgz1sfAmN75iOAL9h1MHxPhe9L7CqdTTd2PBCBGflCnS2e1Ti/GbM+qEBQS9z1x
In8++2x10jNQRI3EVtoByyGcEcgLv8qfOw2o8kBm1/f/TX/0rlXlZDDhHjp6INWR
MKKCjOa0vDJ6IYjUYtROB4+syUFKSXYRxRGBQIqZpRMLSIdzGrVfeTg46NeVoulL
yHnQd1GLWPy2quF4e7zm9uINWpBrHiv5Px0CE0/EGViJRTC2Tmpqx0Q3WIGLLrrA
K+s61TDgDL2iphoYdXjdgZYtuMWeIMzSQ1hJtSh57noLHkWbyFFSSQpIppeSOV6L
D0WiyvsDqAq3FgcSec0rtbWXnWuERmOFrGYX+5LePSp34vG/bN2ismSISL9F9Gfy
ZABaUgXUB87T0jRMXd30Kkq3I7xbIxNsjWJuKIeYe8b64tLV5coPii5r7XJN0FUT
D2Cb1rFjWZye8lUb/+rzPTN/tvX/W5KlpNFa5be/+OJu31riTnZo5LMrZu88eS7O
zSh4ZJWY8Gpnaz16/eCltw1DAaO6mBTVMB1pWGCF3T9b7eWZqc6mn1pMvMyF7TLi
lbBnkrCuFng4bq/DWZM5S4l7uQGSaCSbYLdm1uftBfd56l3NBIcm4vVeJ1gFumOQ
knIPbCRGWr69vBewH/5rCPU7eIAUf4pF6nUmzfOTpH5n6gouTKvcbbVlQazxWftb
TJ4v9dlrK362QONiYusHt9n1oFqaXLYpyPwQZmbZCAYQmqnc1aDdlHDdkLKYFJ9o
AWVrKCjl+FLe0Yw7tCqsP2qc1CjJxW76Gs8UeEcUAgmVHkk7cwfgiPZE0+2dGqyL
s5sx3zqCEEC1q2sroW1YNLt/oZDUiYKkZOhucbkIzyl1m5irtopyb2i9PfRAGK7t
Uqts1VRu4YZZQGclDx4jFnkWqdTGpmJvhPc0HUtA2skatzLiPHPy808hgwHWBbfB
I8Wkq9xcrCGoAu84kXymkAR7ckXmfAmMEnnLhmtNQye3Wbu6llNvDi05IP3kEwJt
hkM13Ur5Vk1I8NzE520HxhBZ169YMCchp+EHgsshHvc+bycOpaaET/h2ZNFKaKgt
86LWkm47JZIriuWRuTQUhSqxZ2d7PyN202yje+iP3fxRE8dbAq5m5LR0plgHyXvi
TJuLaoAiZOeOwMXtZJVJfFpbhHEDUIMr3GtR075h00eOemNECv5jpf1SeW4DLznT
LqKMENnhY9ANoLONZLg+CZvCKzrDdPqUyg8w8novgihsv/Mfvw92/Ydthn4QQsKT
tEKZjwHaoQRBkoDW5QUoZ1YG73Mpdt5fA/X5ZV1vqkjmM7/wziZ0J0cRbqSn6s6d
Aty/vYGn9A+j/gJSiDk35TmMp+aC1wXt2tKl44lp5uajr+MBx4C/okcHzliq2D58
k5zmqid/oXD3Jh86i8+tLkKjipR3OhF1sEZxCRTTXYrsnc1dWCnhHp1Z63QDvEsT
HiquzxbXP5snHyN8XAD8hHLx1iKlLaohPq0m/lHSs4+u/iGBXRmLMk0mfRi0Jcm+
FECIEXmXoMtY7dvU7KCdUT7anJT7HQKunNy/w7W8jKT/ZVwhhIKPWWahxgTUO6Z/
sUQxczAw1/FiJaUOWLIJoW7lDf7rpHl/JAH+Cdpc0I/8qUJE1FRNLH+AFgUdm1ak
Awdv4opYq3uy5igR3mt+sEfWL45VW5ercT0hzhAymz/+soo5CKLvCa1D/0LS2sI2
yndosZClTy0NjRnbe/eLR1yRnYSPoIVbVuvfyei4jcgliv3mMIl/muVvG9lW1+K/
k+XFX+hSlig6QKw76HLKL9328SlMGjcjwSNTXzVL7WANUU6IORb2Rdt9VCHh6DCy
/8XkZCLEHGGiivzMmlVNXbeAy/lQKyvnr6/ZTrPn8tCtTN/0oNrbA8Ry7O3pJXg9
B2vXCzMvg9EQCHCk+8LnHKDctRP7hDhp6mzTDE4lpEV6Hz06LLu157uhT/eLrjkY
nCOojFXTwZd/pl8ydsERmvaZD0RPoIYAamc6cMV6AGX/2YmvPJdrGw31qDQM0rtV
zjQWR7EEPHN6mqYZa08sXx+X8/PeyaGHOI7XxZfY7c8KJoekkZJ60Kp9Ci8SoRvC
EtaAWwD6nERxAnT6+tIL85wBdkxoXao5IoNnbWVapXDtdMiscKI5qZ1WftWKz7Ex
NEN1ItfJLk47nyGlDUmqQKAAgYK5MmitWIHfEl64H4/8X0YhtcJR9wN2M5zMX4Y7
cUjBJOH9XoLnF1MlS1xLrFIB606HfNm4IekkTZdMASJO5HZLEpchscFFJuK07drZ
DG2z6L9LyfT9QJTcGRez56MUCPFbz9u4agH4aY6qvpu4CW5bSECvxfP+WqdBMGaI
wLMZAV8PIT+37Dh6J28Um9dpDcRjjiWDN2LqW5+hVbmQ/VJifDvDBZ2JShN60H+Y
DP0oHtwygu9y0EkRwqEmm2GlcFCVPrra91Uc6JSiOcY0OLD/cgzVQi6qsARJWU6H
HuPVS3W6IAWOlxCawiePTdQ13GuSseNNzIM3hv3m2D2Xb6KBAg3veK2fC/8QRZ2K
cX408b3DdIqVVQC2nt0Y98P0vS+1DNVYU1VGmiJJ2Pa0Ft47xVfV6+feYnwnW5lt
ejNcu6+UAn+9mPGT5OlqrArifnonfrODsZsLjRSO4vQqe/AJ5E4IIxlLbxUX9c74
+5hyKlI4va6xvaMsfaI999yLVy6LGYsGuCn31JKg/yfaQiWeA71Z+vZ86cADicik
YsVd/veqWTUFMIIQ4yXAZQgAvgae8L227GabBI+6O7c6zCPBzCtHtCaxUvYV1ZuX
4LQlJZgwJnkndESt+3AiuNDwQyrTDBNBNZT3Xzz12m5fCIJbyElPTfQuYLTX6W08
QU0pOHOY7mzneiKiLQzARTSgC0EAnBnoBnQltmCUw5Bnc3uN85G+LhSbOXI9teaH
D0u5pAnbhQFutxpzH/fScJaaK9eKRuoZaGCTjr3kbUkgjUbFeYVZ6K8Y19r8bZ2T
EKbRszEiW+5q1yt9luCVWsagCE+6V0fyo9o/j/AfQqUAaS1HnQGCzGaCuKq8eDUq
9G+NJR0WEf5OJFpbe82b648+tVMCIxdcVIIpZJxjXDrE+VDJ8TXmh2un4nA1EuWh
e53pgURKqlROzmBk6yvpfNnJX+lCR/ohhdSTThc73OrhEVm5NMyiigLdMHQHh0xs
veGjGsKKFLirIrFd/DZsiN9qqdnpP/fmebMR2pfAE/f6F9QbShlDkPAUGDQLLZIP
n3piqfpH+DxwSuzQF+xfE2iNyYzPBxhJyltKrzZzLriJMpiD/T4/wJ9Xu++dXnr3
r9nlzQBvF4JU/LJByIYaQRj7odV27212AW03H79L4rCZwiVXYbURmQjqvspqTR3e
qLzvMEur8tKrIf210klHSOoDsLKFHll2UC/3PU4wEoJI7LttIJdVxIN6mgT26Hju
u/iGxRb9VvZqAsAIAacuZFu4f9ymT/UM5Vp3VkJkiXRFSVzMsf7Ly2TXMM1BuzrJ
iY/lk34joW/IrX3Nqiiap9L1KM+uhvV9pNVieaRZjTfjkJls29AhVvjRaJJf/QLG
lO/80sLDnI6AF1nCJxgwKm5f6k2j6djDe9SZ7yWN4cdSWIsplx6/LJm/LxGFRTM9
IMKi6wpvRxA1f3gIb6k2k4VjlxNISb0fQkongwBHnpqqgs5H+/4FaDZ51fvdbdJP
MDBrM9p1ITocHfAss3TObQchmzceQD+PzWBNFUHfZLcFaFgYzYlELD6wiLl3OByA
ZKJ7ZS3kNveM888MnTXalNsHi815cidSl4kLkxzoXyyXM27/n7WsQ6G3BbqKfVef
cAqqcXFWMFsPNlU2Cj/JwPGOrgI5tTx/8Mha1ueHniTWNHZ03TdMbOKR3h7ySPGx
/CL+voeQ+hR+htHXbYius8yrAHVzjI11OGKchGQ2Y3lWf+lu7wmE3WinpnoItLUy
k6/sinl0yuVfZ3nyc9UVs5LgLqbddbMh8NhVnkuRNMVWiDgn/BQir3PpUJ0/qWxd
e2PSSfACo57KIbZVHDBfolDEeliEO7DyJ7eFRGQfoIO5nPrvYSAXl0v0RbNxUCVj
yrim8IaN3hsKYmGohZhgcMU1nfLt8BO+quWTZDrEjfzc3e091ob3AweIIhJO4BZ2
d1gZ+70KSXhdgvTn6F9pRVoF/iehNYYXz8ioRDRqvFyMcb6HH8KVcYjSU+PDLdU3
j4xme4odN2L6ppjunUlDSHYGDmI9qMNHPrrEw/tjJ8HZ7e4boA15P0NS2k2L9/IX
9l2Ru1NLIm8hpGM1bbWl06V8o/Q5GYEiKGv+K8cLXFPbBSjaH6ReBhzvDeeCIZH1
XKOfwVJAyIBZS8HU2hnBPWx1zUMzf5gINcgrCWyjmEjxC5mNXBkAhC4DXTGqCyYU
zUp/5clpI/NTqWlpCUyFXwOdQr6D/12bizVcp8AASAjTu2gQ9yfDCKT9U6ZglGiI
yKDdk9P60wDXjqiQfu5XJTMpL6+Qvj3fjd73O+hj9b1B5wyu4+ICo7I85LUceGN2
/fcqyrFyLG8TzwgBDQ/W8zFsca/g2WHKVvkLI7ZOMBGgaLTr/ylDSQPTndmOdCh/
iCwM/0Ub111/duqqc/CYya5ve5DsZvKyA7ZI0zPh8ed7kKySbGEVJAQ9fK1aZW7F
Sk2WLc3hgVTuY4A/eoHJKPKiAOEWRYdRU5hDd8Dcs89vJb55wEVvXVNDmmFups/I
SkZ+WgJRpXKgOJoRXLiIS+ntNIZtg/5QNu/qDikOO7pc2yeUSrs5d8vV6Ytmp3nm
J+g97GudCN6fh2KY8bbEuUtzwlCftZsNj9i/ZjxwSYQgkBVHi5Be5bYYIPWejwnv
jsTeAHAkVPW0WJL2QTedG0kEACQ4Qr4F8IxvFhSXbZFXLixijw8wo3EwlqFguhhs
DnW7sVve8WWiHawK/5UXqG0nqPvj5gjOUVElOnmHyreDJ3XjdxWD/KAwLWfB/Gk2
+7Axha7luun5CiPsg3sgXh7fUBSIofxqrYmHMTve4NVfTXFp3MLHrjwEbQFkxI3K
iYQdQ4x1UOfvfnwUGSpZi41IUC6QhB7Waql1i6JHBlaGiBSCMBu/g/Bf01483iX0
ojC+mK6K/Uf6eMJGrzcZ2AI4w3xB9R5ructPHGVoqOjPD3jIWhj0kmN3nY1fns0P
H13paC4yS2nc1IyUUz6qSkWyzI3WMAwGw3vV5p5UiMHxnXoM1Pw83uho+ejTbYnX
gDC5j5MNcYARx//pyKSxhhDzUFpcw63QraY05YTY9BzZngoPu1qhh6C5OO1nuIss
bO3O/pe4iMtsAJFwy1dvXNdvtOweJLn7b5Qca1hxdsSjEt4hc++RVZaQXts+Oxfo
fZn/rlOv6FC4rSalQcT2rCqLbpm/hkUrIYEr4KgVYZYwF1lIKzjR0g/YaByktEka
9bBVSK4FQa+enX+EgrXkXaDkiozPYZB2WBM05CTA5XWwHXVUUmIQf7tmkojF6rTI
DPrQ9vfMPcSC9XdvBaYcZoeII3HVgoFUhWbble5uI0jzVlktBXj6qIA0t/47/R3I
O5Elmv+kHgisoruStT7oMYO6qnmNF4ITJcmQcFB7I+HHdMsEXn2NeuYsci7vVS3W
TxbWXgyS4e3vCdaKlUYZoTiA/hTQE7uvqudaZYHvZp+cd5lxB2yH9V9z7a+Lu6lF
P9NKCpMvn01IKCbSyKamjrQbvahO94fwWqv/LrMLcLTBHUOKpltHHWTeOGW47ozb
Td3zghF540Bj11hsJTUPGWYA5W6bX1YUmKjEF0o0v7QtVo9UsekSGx5uHGDbLKFA
9tJfG1SGOeTEwHdHagMajLkDqSPtzdSA0Zh4s90/lAMCiayIyH1NSzvNAFw8Sm89
LiVMkZRUSrtDxDWiCmu4nhRVPGiyv/ROPQpAH2VIiSm8BnlHx/W3ogI4vaTND9R7
F50eGU/J0hipHXJSb0uzU4uvvsBZcBk+fwQoLEfB9i6Yl8b+qs2Tsh63SQSBhX1n
Lhm4Bvb10k/motIM9jMKrQaR0ond3lhuqSHsetKsQmoI3/YSA+TB1aEtfSOldYWN
nyVefIvkDzPVqOvIcGlREz8+gqjHrrgd9kfC/9WKajIHhDVO/FTpS6l0b8GLrrQQ
eGKVeZ2UXpp51Liy5IfBB9KNvDQ5gGpCjXNc+0vPHMNi5EW7saF+1NFj0wlbOWHM
88etgRCzaKW2y8FKBgCP93YKGWjsFEGZcsjB6cWx1MTjU8y9k1OtSESon9aePDr/
5ieAVJnEeMdgE/5MZeEVa+fprHElxG2i7MnHKnneOzrII2O8KNc1Gs8iYz3k9ZO5
5tWkl4jbRDLPmJHeVw/uHG1yScccI3DMm5fIAH5IyMgjnnyRyYAtU0anmaQzsSQr
twHFiXzdg3DTJIjZea0GWxwwV+yQqTgyScRyvuOi0M5nP4BumTBThkJfpfpqQs58
MPpRwa79PgsvcAR7GEZI40k4Dt7eXnaVLKTGAKyu3NZn6bS9X1L/A0JrRiJYYJDb
36YVWe9WuLDOUZomNec+nH5eI+jXtTqzQakFvy/h3y/LvQyuihyV7w8aiNrayNZ2
LsWkb+YO84nOHhY+ixj8861w5h6jgtlzZCVvN7HbWozQZKUjjEbRznty8gYWWO48
QcN4pAuxSJlBJjASPk+ouKrGeTmHbIddxKpDAgQx+wgKFTKj6igAfF19Y3utxy9J
DQqQ0oJ5PbIdgrmphU7QLH7As2FUpG+nCogu0J76YdJIuPBRpmRY+EQkKk9WarsX
nRvTgcndI2f9oYKNrBCIB8oe4f7c3pJNb3jYWACYyxpERTifUFOI0GKyfnoZ+2/C
bp1nPfYxqERBMVx2jalLCav8ozr3wMTUrcPbKyo0RWyk6Egfr7Lp+suYBqmmZD2U
XuV0YCRoKFkB7Rdu/oTVH5pj+fd58YwzRrT2UwNZYCU/U4AN2li453HERMr/ghI9
ddQ/U+G+uX692ALdhNHH5Ts5S7AfWS4BTVWnEnCwdXO44jDAgW4kvQiDSb+Ke+Rs
0YoWCsREyrv3X8zKVnmMHRQFHGmCxPA5NfqP8RsHYJ/fAY63BfMa7Rpw/a5n1kiL
k4N2Vw+8Wnti5XorJiY+8OOkpnwqAe2f4qmA58+CPRai7kE2RCtPpfN46IWTG2ng
z2hBP41PRdPEAuvWGR1Hidf+f2/pko/yi7HSJ7lalFdBE1mTMe9wZqQeWxM6nQug
CbgXEgDpWgrO8lxuhYIDt5U2WtVfB1CCLxQO3hWVlfqpEhVgDLPYP6MF5sSad3qt
jJ/9kpQE3JFcPoKFnyct6q1771D33M525G8uaRgoBUPCXsOsnbqcMVeQgEknbZC9
ozWBCMMy6kOo2N7nethEtLbnlCBfJvUt58KaQbJDyPN2BnlqzYN1VMovcBRSLFA/
Mjc3PlFM+eVr3tDXPOHXsuISBxWwIedyFmpSP/cc5asV+RYZq5sv4j5P3ZN88cCd
nVdw2dzmrXb6FGMGd5Nx1sDIXnI+SYGGlBFsu1CbE8t0crEcbvYWMfYp7uCWgYB4
C40N1mqiLX/IGLz0BaU3ogQvxghvPt3ncNwkUVHSxuB8KoHBY+w8gLbh5oQ9T1cJ
3sn1+vZ5Dlzpl2sC24ShAXxvrqwbXkPy8fiqCZWy2No0B3qSG/5jSBZUMXmFMi8w
JfiT5IVHytC/PCYupScTIt3g8Mtg/21U0ODICfLbRhLDPXGx5hCp95lcMguNiNls
aOw7QKINP2ZPEvrBUQT6fx1w9aTRcePTBscntMf6YniO184eijSEloreN+IEK40z
SK3pw44pHF5mVDRIJfZCF1s+TGge0h2+REqO4A17z89V+vZ/c02mD303wsAtXLsm
yasXp4Cyv/7oaUroeBZsNF5r39CFBW6M2PDmbteWxZyO/texT0mT+mfDje+hEAtE
nyeFdyyrwayS/Iy2FwR9tjuaS9rHxQHB29lO9HukAXFnT7wA9GxcjU/IQ1Qo92xc
QxsjcSa62t7msjuFw7vVrlzPpuahsa3yWGfccD+GVtH7PvyUfg372fdFpq7P6n8X
uHO92RhFM1MPONFptTQAUlO4lYFujYAV8tjC4MhCIFo1ZJew5z7YjpyiM85McXF2
CCPJG90c6j7b60vKKhr9vlkFI0HtRTIUnrLq+h4+22eLkmX0f8cX+O/FoX8Sos/m
XAv8mYZAfOmjNjqLxKdBmqfo/LA1ZoEMDNIRuIM4b+D59D3fmjSpoyjtjCLqK4fR
YZtHrYWTKwG50KbnGiF7NnFMtA0moJlXVGxafHJmTKySNL92psHNE2I11YHrtEP7
VeX3ECOKTyZryQ2jOEFTDOWY32m4uBJCIrpK8q5i/Ylda61ZbMkUS/LrUyN1ZU17
0oWS0+BCi/FtJyEasFibNIqnywVrJl4vpRMBewc/GV0sCy3eFlBZdisnSAUNfvCa
m7E2N+iA5BH/TIUxAca5/pVCxBWLRGT5TtGxnJ1hCvwWMWjsnGQKYt1wVJ8GdpQs
/xwfKmDz1sWCU8FvTdNsQB+L8wYVg53U+wUTAIPhi0XxhU+xIp5a2mGa9y4W2FRO
tIuJ9wZT2T4ExWucedfAKlaoRy8ecuWEKUQXu8N37Yg7aNLcZTns5vLa3fdkbYIt
nxcoy7TXW3skubysajm6+HkCyEDS9nZjAA9ILtwyQDIwt54h4TFkv/3nFK6x66KM
Eyrc59RPEqQXTIqqQ20SWjl4maYJxRkKuHc5gqiYczE34u5vvp9ifXSdAK5b/zl2
XaIoGjxKyKdCMOith1Kt/a5wHWREcusoWqQ7J+/I4UMXFcNe6W+ygIJmbOAXdNxL
t703Cop0f8RS1MShTm811TB5QKPMID/kU+KuRthFARoCVSz6LDuZZqBwKms2ZEFT
acBu19rggtkfEhcMbc1RcI5rmY3adgsQNa5dLGUObAa/uFLSaOR49Yr6pb3ltZfZ
85RFF+x18yDc2QyWTHETErMjdNNmqGtyah1/3puB0tL4+npfCZ3ySoBBS4QkdZxL
LMPwjaoxTYxeTYHeTq7XUecPyr1uXDG+whLd7VLjEYc8UBcJN+8qTVBya2jUo0Bf
6WkQBepr+jgP171wDODR82hfNh5l/sIGFU6JaxOw6tbZRA4Kne5wvYgJXH1UjfX9
Xa0Nt50smPtJr9VWWrZY2MzPI5EzWSF+DrnUyKVClc3xbgrLilGjsIZkFAGxV3Mv
Y1NTsbHP6oL/dU7nmQ/93U9Yw7933yiMIph0ECzkvSv9BHVMa99pYjNLd6V2EqkV
kB5YXi5lk8cKUf0iMIbdqbsxJc/LNmtifJfVJMdGqyxRVjQKggF/nYuVzssn5M8A
c4FslZ+nhV9Pg35nlcc2cRkGqG5MR3duZFfFwVdarApoxwa3LOcuVMtWKVxKOFOI
YhaIvhHkJ8NIIGhN2D8Tcc9fFheZmobCc4q+0RbQQF1L4K9xFlWBqOeIJT01thcL
vF0U2b04TW5fc9i+NiOcUbPNKZsCI9Oq6cmi59Px7fXu9pSk/bO2+wUmWy+abuzd
CyB/hjiYkVSRBLi0oUtTP7pzbkCgFhDF8l6VJ8SFzRm5974nKGVuMiHZuDTKfyvP
daemFhQp2XPG+w279UCXoVMkPqRuMoaga+z2z8wRGuM22pGpPHyngkKqUUAn+U4a
1X12UUCCTF003O2jO5SN2SU5D+c+MFave8DyOq6VeG+8sMmiTMqVx5SphP1zH8fD
SqloWQ9B0067Dz39Xz1AmJzNkNNIEVAvXdXL3lxD8CFFQ+4G8F+3P5FHXsG+9L4J
DKxGG08t46TPj+YoonbCrbtdfYE5OtCsXazfXNtuhzwb6KP66A/b3vX7dR7PGYUa
pu8sLa3FEOx8jSmtu6axwv3Tsl4m8ivSOTR8V5SBjw8v1smsHIw6CIT6HMjf5qj1
hkXcTkPGT1/TIeJsiS582+Uc0Tlwbhu5Oh/ghRGpu1qNuItJLyUjv6IIAuMfb0ms
aZJl82+C+aM3bfzkyNGR7+rpNgOInEi4omRleXB4LoH+VLWFEexYUj77IrLkWER9
GRfwrcN0WM8iXkn3mIaiiPvGM3CI9mysnuodTALclrLeSjaArZxIeFaeYj7lXwXV
2OwT+v+mlutqhjgjVzFPYUPXLw6OOkwavEw2dgQHKZ7Oqw36o9bjMLJhiW/F+p3i
Y/Yvjoo5D8LGVIZZI7EpwIYRHYH8SwTp/ujxCDkBTYgU7DtnBGcBVwPv+RPSYSN4
6T2e4wmTp8M6RU8k1+FR6QjWNz0a6jIBDM9Jsh6G+DPuDsZyZqCD2ClehZmtBV+t
VFXJ7tGRo8oKN7DqQsZ8f67usaCw9sI1e3S5dp311xWPqn4v0j98ZGaYQXDmB+6T
Z57BorWvSSFW4b0/ylEGhiO9eqXmNFSrrX7INoym/u5h3DEafRTrmaM45fSTpjzg
gyVc094Oa8SfYtf4RCKSNTqecC5NZzszfcd0GMx+N5NQtcpT/Mq+dodszSaxzqEp
7W1kyLtXe4hnv3w8DmUzOzUZnT1Dqt0TwK81zVff1ZVZ1YwkWho9GuUjmq67VZqD
lSSrK/51QiRAolDSFcu/lLj+3iq/lpJutf7du2kxhwdQKfZ7hGZTFMtEA6SMql//
ybvA8NBDOkgb3646IrknDtzSftH7hThsuROULKoqrDYKTZ4KQlZadFnQ3d0qUNF3
SR+7bitwcgZdPlMDkiHrqn8tAvHm6I/uTy94yB1u0i4sZrHHG2drKzZL3aJIMdKK
dIHjMYVIS3IKkaHtSytXCiSay4egxTl1we/K6ISbsfWn1ivJDbi/Y1+XFvX9Q/pb
6LB8W+lDI3T11FbsXEWCQOgOfSbM8fjnEpO3/4am3zkcvk1ubEPrN6cOSUwMmsW2
FGbw1WzghEZYM4ZwCNt3PjqNPYLYj2AkAHJnqFTQw3ggVCWnl+A1GpxmDCG7brqP
IbQUGG4N+PeFRoTo94uFo00BICi0yJdHgeV561X/4ApNHTeYysQRm5P1keMolTFn
qpy/mRu5bfGziemXeWyaoYMB9dbb1WPXTHK4x9f0Oz5aRfMKtu7YsnD93NmUQlbg
OMR2PTV4WWgJoO2kDKVIntoH+rh7qDezwBvJEyT9EsW6pOIxFOIGgsiBC8BRrm0Z
/O9L88tkN87W9jTu8wzLsYFehrAPPLzY18Sl43Nb8Xuexr2euXuDGi8KvfaQi6Ob
31YH/FTPj+ug1Y0YBOA0C9XULiumMDnroW102SNfmmh86CUUvFHWsyDT6iwmO5Dy
I2kf4SpA53WUzkrccRm50J9Ss5Z92W9SiBsUbYMBjvjip+PqDYoJswagfohsqwO5
gcVIflmhJ4LsjMlbvEKceRlJ/gvtOcQtF4mAvId/JqzEjSzwnqSypJJ7etI/qad3
TXKJRNB1bd2d7FVYNUzGWTKb+zbkflIOtg3tVRAgniGWh0qlYznOCV3HOVdeHgUN
cEdAQUg4b7NBLkuzQZ0ZTnhUyLq8UyhPzSt3iF5VokYrytEMhLPIy2ChN7zs2te5
MV/LY0wvgEKZsPal+34jQDlxfFGdMKNC7jp7+l1VLUNy05p1gAQjkrueQuWHRgHc
MzTq46b/3o9CVHhlUVjkvN4wqTzZWXcSY3CzAhV9c50LTjRbZbZgRsnU6wCgTC1G
i/mRkuAUniztGSxDxB+C9GqzM4jrCgtbbEPqewCjLon1waObWGyzPX0ZYxY49zge
otR6ZUbQ9BXjDvzFiL8rxUFXmrYw3/6ikcaEb1bVE6eZFzP4zzHzgfp3T2e09qy6
UMCxvgDirS1IunMi8aD3QJtbIKDtBhdh8nLfH9OcQLc6yGo8wfAMFAeIyQFsfErQ
lUP40/jkQ220nv7N4kNUdYTxJkTi40mOsAAQEKIH1tuL5VcM2tOT1ZQsv1N+WIkb
3cnRktKi8JKHykeon91pme+l3kWKL789/558EiN4LZOKJGJCxab8lj27uN5BimCo
PJCm33PoCsx9QfnBdFDR3ZhOqO4c1UsGjPoYvc2TBpttgapNn/sf2VwpppkF7pg4
672wfwlm/4tftDuTUdJqyWENQtXUcneM1PlF9uhOYGH3OjiYQIGwKy8YBbnLNTBk
hVh6t2TZ1PQVpUGLDqVsuinhh/NiMHwgoBwFyAOrZvqJSrAFZTeW7m1ix7vWqYxY
62Ut6jGzjNnBdGQqdrTsS3izFQOAoE614MKr7LO2brxhsgn9mKd9+F2wUWCCw+ZS
vcxXyt+zJ42Y9uefiduLwfimJfNBaxMRWMxw5TEBvOa0YOMwNv4Ah+Dp2KVG114a
+E0bKdHraQIXs1NNbWzjOBdMZBynkZsowB0OD8oCnzt9PKJ5xGdnC3RFs5adryoh
ZBWKWarviNEF8GEW2b3/bj2wWqQYtBWp41L+gz5ksHFBje1vZpaFA0OlU1H6Sugf
BXwJwZTFKawkuI7XwQpkbZSCcPzFQxsruyITjuYGe4mRq+Ox56lxrpPbxO+F0C7J
eI0uHggoqx66jFO48O76M1qZNQDaMV85E2y/4hW/5RI75uRuB33iQMrTZpyGSBLD
31Ec8V0+QMNZZ442kbKJTx1rR9XhPjUOSmKdphVAZnXRjOySLZtpOomDpyrtJ4Uy
9JFefrD3gw8q5d0jgNWujI6gzFLxAc5NYh+h7naj3qbyR3dSpTNIIMuKIpOcsYGc
l7nwcbJicLyTmFr9wE85KNRqAk/VYFStZA53kHPrNvftun9KvP9XS2W6vLbjKCR4
dX9Arw9xxF1CGLPiVumck8ypAFY6TePs1737yoGFQvky813iDlXTBTYvLXl3yyO5
WRWMm42Mejf9awalhIsEUoQkD0pcZZ6fA4WrhyscQi8gfxvvsgGxWKlXTDqV2jDU
t/PmozF8V9KvWUiy10d27eZqXQQUkp6gjD63J8tzbxvNfoR5k+1lmWLEUf8OBYJ4
JKH58HNZJFQFu8xCd4+ZeXPtfTeORnZro2hp/Ed6TelxuGANWgQb5QzvLc35TriS
JB/zYyWuUIxyTqIwnQdVzd7miu3I9b9G/GrwUVdIe2JhW/1s01K9x6h86GLeGA3/
saM/mo1qrg/eHU35bNqKda2KWDeJgU3abujFuA2/83QqBHa1n8cmLu37RqnutdWM
ohoOjtOCX0kjcgJ/66oxjcgUgnF+sYzV+8xK6wzBN0xLap3LvRz/Y8lqkU4PtRos
kvkKft9F2Odjgj0KVOXpIop1CZ1lyur3VueShcfK3MP6h3xLAv5clXp8+l7Zl6/V
45SOxIqJPwwz0Q2SCP3hxJtOfCUDvtKCKfBC7mbyzt4OJt1IarqvvAKZlBrgquhs
X3M+RscPTHsfcOsM0YW5YGsYaMKkkqQ4vhMVmzqQTJby0EWov36bGocbQOp3XuW0
7Um6A0x7b5/sAqxvvpaLdR0b4Jbfxay8KeDLsMEK0cSipt3QnjXajQa91eVNTg4i
Fzu5UwijhZa7b0xSGlORFnTcZnEz08e/wUq/ZdIUr1ku1P7Y14U/N7eLFBfqD0jI
5LQAcbS5+xP1SMfmyu2grIiyqd0K1ly4JBNoC3UYemZuG1OH4JRpNKiEB+94f9tq
SMy33YoSuczbqGC08JAfNkF66rIC2j/jDYy44hCMyZ0ViM4U0E/qQQvVv5sjhi+Z
l2fDe44m4u/WFPbIe1UTfydDFnZWz8vpp7s8J31/HuCEnNtYJsmyvL1K7nAgqqge
+loG62Satjqbt8eWqrFg1F0sEld7ZkbAzZUFDZ1TXoZ6LWA0TAwMkLUfkfwrbaj8
xz1KAkdM5ATCr1dVEymZtg9z0dYTQx/GsgHPYu7WhJOwGTTO2lKii4gslqc4s3yU
hW7xbFV9KiC0oGbz2Z6Nz9buCqYU5OwMTQleYDMBwOOaA/fivkvXtMSvBGA3dS8P
fnVLbC04PmDtpALxuTY8iApjuSJjG3m4hevAKOt63NlZhUEhDAxUUxUlLbgDYRCC
KHwagVhnIPoIXXQ5kVvd/WOoa9XxUUdDpjjcPPZo8qN218vSRhC7r/4aS7/zyxWD
by5lY/otQwiALhcKUnI1Y4CmdcE26OqCwXgUoNgiiPFHEBSyB3Hi4C8Nqs93T6mx
kkZd5p0YNKRPvkpuDKcaccGDMmq/wv2imwBqpKEo/oLKccfqQl0STDohY1SZAguC
TaYZWm0ExfEYewqMI0JQrnmzbCzBswpLIgYuhiI3o2jXLF7XSmAtV2RoVy7gfy/8
1so+xk75jfFewFrGGTvg1xJR6t8b9SDi/OwLVDkbLf4J4KqaFs6ZhzPzz2MTOPVy
cNCk4wKdxyqx+JE9THacrtZGj0Uqw3gGt1L8efmfKVdlJVIZ00BQX/FWqlcdwrzK
bj3IgvzmU55Uwr4NI8KGpmAMnZzspypQ0E3qza+DuQewcDDf8qDZ8T/ons+OwfI0
IBBajnTv7qTY4rhDYWkdOBCCT5Kv81VRzqGiihdtBWa7lRZPg8W4A97zOHGcyDsC
vZSlv4HoxFvppy3OaJV1DniXcD6q7AgB0RpolTeQSlY2JL9VfhZ+dpUwqICLFvKp
E+3VhGa++fTOM0c9RQvABuzswZldvtVsdHem9z6XPq+KhuUx1pVqyKddM9TZwCTe
YRnTgf4KDKhd96onrVwBJmJxNu7d4QKwewmYy2U7KOMEEnSaWTleElrrl53cdMqv
icvFevZHZY0m5iKUapUfBO/6m/TXQ/xJpM3OCm3Sbd1vTAKcHye32mYaNPmdQdtp
emmV0PVE1lYWfHbDl/dKC3nOwxN+uCRH74D9vj2wwEvUo2o+0V2b4NcxmgrRUeFC
NVNDvoNjY4Dsk8GQGThkKrSnbmDhvGHKg3+ugSUdf5t+BvyTyNri4Ez4qKgurjGP
SA/710Ra5T+YHryHnEPMx4Tk4ib3R2u87xoCy4x2LZgfxsiRUHjWkX599gj4gyse
/Fn+inP+dXP9DO5foexN2YKoCclgzd1/LXhR2JAXC/KcJqi5tXwAwCh2YAHoBzOU
v9X8YGWaze/JZ5jt8jYHc7CocAkYGl/DVvOi81y0vlAkzKFtXkNi7GMrsEexxJ+p
8En4acrVHKPoAu2/7Z6DCGhwzOtN2SxVLKu6WQxlLt9qqkiyKLSkdbAqVUgUL3Db
7bZttR3YEuC2ExFC71+m8Z0P8O/ojUepC8xaFcqn9A7Nsv1dRZNURcf46PeKX/wc
tDPDJSQRw/k8tMbLBIQEJe6bv2EgjTraJUFu0iLfnCOzPqcra0PurxDmSt5uyNxv
UHyteiejGy9KoXTAWq21/ropE1nvpI9pHSt389VldzWgYwGi/iFTSWwITXD/9KeG
459RmBYytSPa7NYvSBS0+CoLLaXUthU4oBZXR/HLXXjc+5fpeGm5T1H1bHycEP6I
YY/FPhCjUgYWf0y3M1z5wPav1dtYW0/Os5ZBTkpHwexKaqWaGisnx/tNQofcS77B
uyb99YYNA1vZtfgaeTJOYQr9WvQ/Gb0Gpok1heGYvC99cO1b6O3/e8L0xXM7rf8C
dkmeI5xzkdMVulvaRbkgPK1Rt9XpdPfW1Vr/xFhJu4R8sl9ieIgwNt02VNPMY+Dl
+BQ5gpPSpyQkkNJIPHvUmUsWyfTOPHbWWnO9TgPxyI6raukGpmsJjy4l77M9UUiU
QBjvLLjq24qXizP1ZlRKJPk0B+J3l5TgXa+yydpdPQ9DxjK39/ipEXZtErjeTBVO
XUUXZw6KDqgzzuyTt54FJKsxDLcXlxex3FEVT28NIsO+VrO4rHrTsUV3tsgJ+rVN
M28EgAfr691sMyl7HcjAm/C4LvjoeIgpbDASUveILbwg+PhoWnDtI9i6GR1cvv01
YPp/3WJKW2rSyb5LywOFyavMYs8I0al+/fuc80tR1jf5gXGeOcsmSSqRJhTGBk7z
e7BdPsmNm4R3puUN9nutPSumSiGdvVXQB8my7dWvoyifSEHkhQPw5bQ+3fldodBX
ZAo6CjasEa/X1tYdwyR+tWAgFzPL5k/y66EVWayFhwsfmXrJScjtncEu0n92kkt+
CBxzF0iIGPJoUxqhrc30Fw9pEYfg1STQquP+sY6XgErf9JJFac4QSiZmnn233mCV
pqc9NnxmfA2n+U148YkayASUlQo9aca8BawZwSyv5cyUl04WnZCyYiTJNeighIFz
MohYqaXwZ7KZiwvDcz5QMwwbS0BLu45MIMPOYRsCZSqqDwq6BrSMRiFad+uKgtNS
WgaxrR1wxF4nBPbMq1j2X5yOIzYXRVhQtc7JYLUZJ9Ui2OF0/UQH5Y2ZAf5ZDUWw
66VD336Aa8LoiVTuwvpxi6OBrTe4hfiCyri5qD2RrQru/GC1k8XJRjZDCm9aqE7x
JSUUmYXtL9+KANDp3kP5T0OjvEufm1hyAvgljcXiL4/C5mF/NLaYblwQuJy13rfs
KmC9yXOpw/p960Skb9356fHWfuehHvFWkuYeE3fusBGAyl60ZHsLBVIRO/fDU4TG
hYPwOOC2QPTWDpr9isLnM4ke7o0xCS7iJJq9HX7cEvuwFN3OOVayC2vpWmAndUqq
ll+Z0wbSk4VNqrRcOBfIJGbU5+S2pyP/mIcMN+iTWeNOX7Fbtmw7OxgtaREpEif9
ugA4WAIPkn22WwdvfvpiDhyzoWAlp74sK9lKJnDpmz3Fo6gA2IsHtiywLeB/OZ/U
unmeE9ZCSx5k7XyKFXJMZXARZ/xLTfl4kueVhzr1gS6b8uJjYtro9//+VUbKh558
ohSHLjBOQoLqsO77N2wpJqJFRiMIr35ynZmWlm7hXa68ugKGYbG+iPuJ2pJ332Lo
BP+5NriEy94SA4VTgGMp8Zk2t4zhPlkDOi9XlwPY8FnXKMcQBSWSsrKLiJlqll2u
9hWfHKFjlkGqCTuP1tTapuhEEXguDwVC6lN8R48wqnsfjgsJdwfKDjDRe0k2+0CS
vQsUWJmDnUcPdsoWm4LBpaOsxUovg/A8EkCAUL4QFmkzUZJEe86vbrcCs4iPsdHR
yAzqpwB+gRy14tsa4OKAOlBO3/KG3cUT6s+wg0NkqtPhPmFDPpgc8iHe94wiupT0
5VJr5cHLr7cOJ68JJOAm+40GM1Uyyx62x4LlzFk0jfDW44gnH5LDJx4eqU3yGUuQ
pIavE0ZdMT9Zl5yrrggQm3kQINydvLJVX7Xh3KH4AHht5h8amzLktsRNIY/Vsjbl
SX5AQiCxMGzYzWwd/WvABEYSKdVYYd9nQAZoem1lDGmPpkHWk3EXR9wQj0I2RFMV
ghf0QzAnJ/rrrmOqdnfbzOhjIgNDFZCzwbVr2CLVYHKVxITkX16yMCKEl4eoFXZQ
ownxcDuvbh0T+Ua0TkQ6ZCN5VfgZ2KwtbuShqFwPtoyyqO/h1KjSmimy+dkB0TdG
8dohIMKrIkC8KDpakxryXznksY6jzCRsbzVbV+HRnfuPNyJxtHQgS+w8xkOlYZkh
zRaM23IsSe6ynlmXglUsZec6eTTCy0XhS6orUpTuYFuU9fWfd9vIrCOwG7snVLQg
PgRnjLvm6sdmVajwolIIpx/zY0C+6xZUkYOWP28/Wi9ot/ofhurDGFh0Z0aODWSk
npK29K1LYZH7DMlYpdVMNaE6Q8vqm7s6uTATnDG+ENlyR6YUhTSHc89czKGGXeM/
xxOmSV6QnxwlU+1Sump4jgNWx66XeA9l//HB4+azd7mFPQEDVol2/MMEO0cLniFR
PqAXDaM92sxsK0cFdTQaKwtqPVu5IlN/wRyxf9IGe73iynYrN8ouTsYZ3pB+e5RG
fOEG9LPlW4ko5VUEmpQHTS4VKHuu+Spp2Xs9r3WysbbLNjecZOJC+fnMUdu2FSVR
9XJilp/W3Z678ccMVGyq5wmmmqOTxkC0NV2glg6kBsP4+UR4DrUwvCHmBGBaj/Gx
HsgrqD3nYsLIMEswakcv+4kworIWUXc1/crJ8otLOXg+TNyT/qL3Qpbuc7Y72vtV
rb4xZwEOc5KGlxxSLlfAaPtWXbQdk40dPYnJmZmoCHKY8Rig6d1j4JBj2rzDsgQH
JTGZdUgsz7ULY8T4d1lxAhgn76xWC8FgTyK1lRRUExYV7RNJSPievN9HQ6pvSjH1
FVlqZrdxcjne+tJ/98i1qvxiRTT1LmcKEaE8JDz9JOShemWBUHSd5CK52RPSi3vN
nfF9trQVuN0KcdqSUVgxzJ2/+T+PDHjmd9hCPkyLefu8M2v0uIz3B3VkzUO1r7pU
6ES4nio2JSTzVyjW2j1VN6RlJiNjycjtBRz1CSiCVrxXP1SHQfXSkjEh3uU676cT
2l7ZzJoa3JM2MEB6SVZG4M+vA8Jyll5M+jIzEoshZem1GB0AZwIIyADEodDoguEv
IoUd4rB+Cb7UkDs2AP1pYckbKQtlLgrn+fDgliJ/hja6rOxw944UZDpftmVG8N9Y
2I1UyAp0WxBjPsflZfoz2gwxzm6LuszqYX/g1RL38fP3azS1wMwRr/dE2zbqXAai
ZxNFNeGlECJtFeHpRhy1a6y6Pel0rvUCWY3wf4Jqzzhb3mU0UV9PK/bkFFtLR4mH
4tzK6DaJwrwCnefD2KmQPt7rwSGFlvSD1E7mDGxvR6SxkwhJol0VcWi8ouFkB7GV
6dMyGR0qSx2Xu+G25E0OW3cusfSQd64ksFPH+doD2oJ8ZiKd/5CUdnB29lM4hE7I
QFeIbHdDj9ZNDaWHhvg2ZOzBOnmkBjyNTA6diQ9aSY/aIGUX1Af53aVHjSFs8Ei3
34I0o2jkMRlBEsLelcR881LTf7oTa8nNk7tRLAlMiKqKDyAFxFo7C9rH3iu7qNX6
ouwLbAHc41ZfSO66vc/aXfHZoQE2Onv2SXpG9I4+AQ6rk7maMgguwI0if6i5AOYF
/AoPgmCW/z0FRPM4D5MCMEgwmA3pKDsYFgvGwcG/J7gtzA4578SDXByUMhQbWUZT
Od6mQHRFaNPvSVyMOnTa5NpT+jE9idKt13Yo/NJnmt5nucMJMdgHoCVJVqmzE6Yy
N7MuH83+6UlynZYLf2mBVBLlSVyREvGNhwWffWTrshOmWdA0xkitPcbMmUF6evJ0
t/kMJS7ZKpH37rsWytcbaT9CyrYuOfGbOdtl16RtAfX8FbeERdxdg2EPZEy7FatK
zDOB4dXQtoqyaSojAmsZb3DFkSMoyhxfFoKbu6h4wDelELvv6hOFF/BhxCwBRbdU
zI4GWfL/7gFnp3DSlb5DtMMClRmriET6UY8e9uX0So8JPL0QhiMgiHtCgg4ylQk4
aN7iLJMUBtVNXA5lXu62NCdka/wC3ohqgbRjzRfnfMK7bukZen8KmBgBVsJrdGK7
S9RrChm1TBfmN61jbH7niKgaLFZodJ/IdfoN4wCk5C3NlyfdwO4pQNlg4xnxdLEc
JYKZQ9C1pQVYal/mpYcvbOuuiEwRaYHAITWKUBmrXdBImjKA2WkA54bhNGQF7ZWf
dguDjhl0v2VGeaxxKa3SqIUh7XY3xPUUeacaFQpl8Y/8xsQdaJefuM2TJiUm41tj
4XdyoQuZkiqawP7rqKcKOXOBU1GQo9aSWRF0JmT61foBt7A6AKuGTD0hAQb5YH7v
ymUCGc9fNheDBpL/hmKMb7X+gVwzBDHZ5PWRrEfltlqVD4lABoClSNz5juRyROf5
UaOZ4s9tF6WehGcbdLqtS4mMhMzLQHtZtr4q6K2DVe4Wv4I2m/wWaDadZ/x+GReo
wPgWHF1wozFHOoIhYyI1YPiKhiGrIwDJucVHz8tAATZAC//CussF/Ns8aTfBVzmC
j+3s1wZj92kVlcO/hLLqDZHlg9/7ML9C3RdEvUtj7zl9SxfzZbcvjqb6wA2wRtci
PybWW2EIaETqCiKo7FSsCeRHmP0h9vwwCTA7yVYzopKQ3HfNDMTTyGX+jiQP9MMo
8kS1AzDnOI2dvIo8L6bxBzVcYvOfQ5UOFn2CT70ffQlwqnqucbQTWI0Ej/dGTLFj
xXX7zRP+CCZbkcAOiVrI7bvJ/v77TK2w9KXXVzpnXv5b01aGqn+y+oWpQSiYCwlz
4CHj7hq0w8oMnqlIuq7h0YDFFyHIfYRnf5yM/vodpLPspep5XxjVvIT/MEj0DD8W
l0hex5bUQrAl4EtuqobfCRpWxYrmj30PWq9ITOW85Lk4zQ1tGU2vDkNJYtHlavkq
HrgJRtXH8vIghNmcDfz4EyB3Bot/HpcjiYhaQVMJBOnLhF2WmLEjM2x1Murxwe+G
IZwSnODgmEcvtxJKQtmvWxgVIKVJ777bj014Z2OO6ZT2hSHBPS+scwCjBOp6B+8m
ZkchvL1KmKOaqI9IHbOFR3WTArXEoM5zZWj3gfQkrBGnjEwB3IncuyDhBwWXPW0e
mvUlD1Ek3mMNHiujfTbvElJYeQvkHN23CkSyAhVrZq+Ujdkflxrv5lm+52cnmRp6
Hfu1xfzirqqB5YEOeNOEy4FcCdlmAEkgUm2xrTb6N1lSBdxcj2mhA0Z+LJ9eoq4E
5M8D1pRiKV2MWP1xLxRIGqgF69wCbYFt5zHGhHAOuCPUXXV89p3sKPiXU0+fUKQb
THG9E/5YDOP+QAtuxG5+OBx7xYkAhK2s7xR13AJNhIqWuFbZ7hTNFJxi82XExX0s
DuGQScyvecwMzd5+tMVLrNsEvdyvAJcMnvzwHIFhebtKDwxYka2jI7/66nSu4Tpy
vlOyP3+w2fkG/jYLh3R7RV8079Kvna2etqpNxWpyvW49OpujQ0MuL80V/+mqKD0J
0QYhoJRaT+5VLXCsor9Tl44vUgtwD9DzlsKNxl7OKVxabwSTYZWETtsUjREtYGYz
VdlcbsIzjTsuxqnx7DfT1OtATQA43JbITE3kPJHi7fq1Y55mN/K82dMSbAsXdW5+
KgN1aA6WoclnzxO8gB5HVIiIYNd5LpNM59GBOOvw2k79qvgTRjwoO/m1uz+X1Vuq
hvuXbS2m99VWRkhH9ZHsigobLss4LoIOrhTBHQ3w+veCcNVPjZ+K8f8BrZL874yo
MkiSsKxu5jWugdBQnKNyOgjKLy/LyCd9vmS1osdmhR4wM7wnFaAah+l/Y3RyqnYi
wBbUI3g7jt45WvV0PpD5hKu0MTzcY3cda7jg2dF5GQFrANPQmK+gYm1fJBMs+ybl
ZNH5erH39OynaUpCuseaSzIy1xOpH281r2/RtzbOSYUkQgpoYfpkVolS3kTnnMMQ
h6Tb23V4aDmzf0cTsy9CGEMdM7HGXqz14UVBRHjIg6FaPLjDYa2bf6pV7aalbnN4
CLsHv3vuW6p1vd/P3HgyQ6mpR2SIPUjmD8SGE4i81SWvT1aOX+2XmcHUXygx0MT5
hppRa+O3NRjze14hnXALLeI7DQOG5LeArENKyIwzOc3zRRWeo1MGmmhvBd4mIJzh
lHuMJ2jwivaq5+Emn0Cy8TyKO5J6EC9Ljtqv/TMZdVLuFaKW25tBAvACU2EKYpOH
1P8g1Y3PMlA1ohwO+LnZHA0TLmDzkKZ/4MYTg06PCz7OD4/nqMR8WhdtkJL5dSGQ
of9A2DlX5r969DHTvF1B4d5wjfHwqoV9msSdo8gc2sryAOBOlBcW3VOHOlmwYQqU
9FiCvRFbpfYn6bpdFx/ZlwQscWYt5myfFGGhbPjkU3lchwtI6elatN2eLDS85B6S
VKluVeydNk/VaugX7l4B34LGBUzY2+w539qzmOxHQ3Cyx1qnvSRAHgq2ndKcay98
Ope08VTVbA/4Z8R0fAPoxnx4BJZTbUVQmTUwLG0wbcIEhx8/0JI66vJtxPIYKUjK
tGhExGfg5Q6H3lcT48NAusVLfPjZw+4Wg2RJxfh5dm3uHAgGsJYzDtYr+RwByPyt
cQnOd/XmuXZNo/TSMUBUu+oG6pZtguU/jhfKA7TASwhGbH+lc9u+SloU1Cmdru3W
ry5HJ0SlPG0jvkAYG3n8t0JpusvCjr9nGHr6n7n5usMoyqAM2tbZE4POLNDVysbI
x5twl37RUHGfj3enGlTG3UdB6Sm2Bkql/LGwL7wMGR9JXs1gLdn1gxUfo+xjl0xg
IA6G4z1w9rdVY9Gam9Z3XmvzxEjkJjcZ5yBLDuVcF8vZ/n1KDs3olKutPeGE3lVF
J2fCLDowhBkiBUC0nobjzeudbbAdNPoLImEBoZvDAcvqnbNGPoz0nrsd8gkwu/ux
gKC12/SiYC77eydF1EbrxbwjJDxtVopt02eUIzz9fFCI1eYo6tuUpgjg8ABPcQee
RHsArDbsLy8e5UrrzqPR5YkXvZp3Zx9wJj/78h2IKHrpoXVCjRuoBNrW05Ro9DqT
IQ/0JyF/vhoG+17bwa9Z+dF0SM43IQBCREds1Ot/1ZlME0nyDTC0iTlZXmMvLQJY
rWyCXbSv6wFlaVJhbgPfrUcMc9hXHyn1mtxAUP0cKBSS0eqDeKmDQLy5GRzEKp3V
v+Jmd9WHhCGViNGiVO35CIPpIOna3cj1HEaeYYgP+g5fCReMCpUF66qvzTEUbW64
6BSSpNsqV6JL0ZtFRYi3BqVN9eoltatkn+s7xNOjZ5wFGE8BufFOvoVCUotLQJu+
TgstvcVZFmtz+J2o+60pEX2XzKky7Kr1pLPgKBvs0TDAYzOa1i4cwpXAmXfG3VRy
MShBKFbDiQ21dJBGZvrahmdM9qfny1BSRSMxZXIkGMO7Cjf+TwBjcOlTrpCdM7/5
Mch3RSJbOUMlTQqijgXfvSFo4BZjNP8Pd42dzluEovJhcl+F0A8D5dWCIqSt3wbO
j6+9rCK1NaNhaLdYhvE+DO8ZsqklDX0BD+WM+FYP0hGI1DiJqFG14JugKZsoAaMn
FH2XdJjD7onVz2/WsZQIlOGe6b4125cVoOTrHPubV4ebyVSiUG6ZChdT1+R+85Qu
QHHpwZ2woT/BxUhvJRvDnqiwUAH0XMYLcziVBv9ikeJ4NVUtAuRzbQp7qM8kaHJU
eF38nY5JCq4IJVS+xkWNiuw/7EZvO91+j9aQmnJNO/Sy+HNu3blUfkBSNUpNiJad
LOYdjwLdZ+RyB2NHjOKZdE0//X5dcmWfwr3i23+qBKnH0lr8wP3WozEqyWEznd/H
481LHIoAJlUHV19GY/dHYpo0RHaNO0ZhmP6nMHHPxM84RhRH4J9Xy+yfAzgSsTbb
b4Smk/IG2xevslUo1uCs67qCTJiN2xqyQkNY/EzX6iY+2ZyBJOUDxs1qCVHiTQsx
8Pug9LBVUd1Zm91sP9QF2PdVHCccuJipSxYBCK9lBjQfC72RW+tiywAOQvZIn/lS
La3zdgMPnhcaJgzk05khT3W9jl9BFI9rTWXOns0B8zzanXiOrW4q9EV/V6ONOCa5
RBP7SkXYRrhLnJxOqapdwPIQLeAu0A1JnpESlI1RFsA4FkvsXxNs6KbfiDpVpMIG
ZiQvV6CaYHtTJG6xQA+9l6QXdwP4Riu+k+6AlrxySLM2oRfbl7qmfS+811qXdAjU
6NuRqu+859mtZHtQhISigQr1/xl5KbEK4XF+aLchQILHZIxz1kaAQyjVANMN/4JW
eT1unD8uIOPIRhMLhlU//sqMaVl/Hbm74mo6290wyeed4HKoQo77rOWf7yJyINlb
bIrijSsCyo5LD0QvfTkzM3bxWdSPRsnZh0p82Td5oJUcfG5m/lTLSwjIvkUTQ5vp
rkw+YvEg2O0yl0LobOE91QnGXgCBdW8wYB+blqHtcIaC00Svu95rFcNof58qLv47
9rU3rRIrG9obBCxGn7Np0mdzD/TbYZuv6udjJrRrIbLowFGF5Dx5W+lmfWsBVZmS
Noi9SNQVFFfyQFoXh4UE4lFa0ptECLnrUwF7vLR5IwpupWnIqTzAGax2mQlyPG1h
tVnEYdQWkw1xTPjKPnPna8IRqohilLP1+KLFyd4DtrcLf2gdL674OsTG06rg+UBc
vDu97b8nhlwGgyqS9n3YlFXoz46tmCWlM65pG/GNFDEQ7+DzRFGt/Lt7ggUGhA6P
CuVuaPu60039zGucPRbb0p9btZ8Ze/9/0+3ERBMxM4IG7fQ6yb8yEWmAIPWCPs3n
869aQyu1fzFzxFWkqSc2u/t6sEIXiptwWjQCNqYIatUIlO4jzm4lKTehx/SS7jA/
dkxT+N/0urM4/Wo+xbktOpJaGb3WYOQz5FRSN4FX0hBjy143zJfjjYV8Bstpz014
eYEh8oZ1wcsOkCItOpLeqHE8qpvhQvmXJQg3X+xeTjHzsshOG0UxRAKQmhXPowb4
eJzUoHeu/ieV7HxVVlVcEa4m6C61axlTfcLe0AAh5qXll3ao1DgZ+zIQW/bBFCVI
kX35lls7AwbRyo56aEGk8RsCY3t688n0Xej0aSUTrUgfQMmzIYjWczezF9+KW+k9
YwDULTSH+nbHyRmz8e2sKENj9z5qg8J69GvfqpkUhHjbq7hOWF/7O/tthNTtCTfs
y/CUBV6G1zIP8VMscv96RTrV+09jNxC8xNMRVFQQuR6/c8JJj7pF60CqFdJc49I5
k1l0Ph7s4CWuvOEDv8XKeRPps9K6kBOazxOzegmxncZKMDNccbsViyxgPBO+NGBp
s4AQtp9OBQBB1sKHR2F0c/+4B/Exf5tM8+cybktu4NtS2Z2sB8mNvt/F3vLfF+la
7iquMv9gj3W/TQUM51NaZU7B3Mf8I+2aim2x3SaaXoDmk7Akqeegz3Rfl+UULxHQ
awdP6JBAubVCSMZL7hwkprMbDA3HkAYmOHov6dbWtSmi8gPzT7p9/pQYt82BNgHb
G5ehyklBXUXi6LVeBBd6Kry9iPsdTmgYN7hY3XbPvxK13bLu/wA7GOw597hVgFX/
ks5k/mQTcV3B1aon+/g7dVeSeaSASnzVTewVhZ3qOXurXSF67UNKfhK9TZ+5p2sc
yFYEne5nDJDmMOAqV7Nh13Rpyyu1qIwcob9/Ex9Z4BefV/ObHa+DJGiqY/ZO9X1a
KyP0Jmt9InMe4Toa5zDXwFcvI4q5HCbqImqNvv4uSgPad+0thFubu7R/oqnEVL0s
kdarsCrDHsROtfdB7X1y2iytGFHyZ+Jmz2fpXOAswwsb6kYP9JKQ854eL6YLnQ9f
F5XjJqVZxXh6J07sbU/aGG1avpdEBkXy0UxYBqCLFOBSI6UD9bB+AZJmqVqykRTa
qsCm1sVaK3czKcRKF5YpvOqR2aQqqbL1GKiJejIO4XwkkLfZ4aL89A0/cqgFZtPa
xNqXd6LgAGxwKc7idnBVwwwQTfXzDr3/OlVXMdgA9XoSyleAavDmZSwc5UeCfunA
cFwtuypOEB6ldMcmT+9pFWyjijmN+Tf7z7LHTEvAhzawP9jR0eOi/Mvc4FIdiRLR
cEAJtKhtJwgOBDHgsuSiB4OL6uIX/c27OVuC7V1nW0H7wDOyT8z8F4IkXLlTFKIJ
4eFz+5+hhgh1eXQKmHw+ztl4anWDr4se5PS0l/GBUDyunhhx8KbPXHnBuRxu6Zzk
`pragma protect end_protected
