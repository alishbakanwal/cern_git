// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:05:42 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
XgwcN3gB3rvrs32KdH+hQLl1TiWjl2h/x6uZMgXy8BMRRn3DtNOwYC3Ij5hpipkH
ZNKgMNlphzssp5S0ubKJ4dylsmAT0pz/9ggr/xzdZFY+hl8ecc0AqiEyy8E8jZUK
SmDpzjmCjws9MET8y2Cxn93PP0Y7wvHuy3W+WM7V/8Y=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 16320)
VAb7drlcMVXM8VgmS0NLFAUhNEJi7kr1QEMnKbLNvzZKHqe2/xxt3Iz2AHHX9jZn
4IVzc7RtPF2h6yG8nECh/UHcQT2FmvBMP8eUrgsNHQqC4GQUjATN+eoBv67fRCzz
WNx/4c6Ipz8ZOyAXXFliLEgQBldrzUAxLgK4eMhyEPqLGnvVORXrGY6Ig+L0si6Z
ocwPPRa4Hy3MkO9412f/q8RK8u+YpZB6OHSpjExkjdweWns+577uSbh+ewjNIBML
4pyq/LweJver7x2uEZ8PfnAd50hrlGi6UAABu+EPn0/5J9uR1/Fb9EejN5Gnf+db
O04Lg+nIpqB/u7EZQnD/Y6dymZr/+WKz/TNqvKvBaUMmnhgHXfYdGabzEg/FVv0d
JBdqgGsQrFSuiHTRLb5vsvWOsC4cvtBP+u1X94Dtn7wIJoBTaNXU8UVPD/Pu8u+N
KvInJs2ooafelObH7cgsNf8XDA4KPfzFmYaQeprSZSbMztzc67im9dhqtfU1MbC2
XXE+wplGl+xCc8nQ6+RjLHotY19xgBi+StpdPhlH8Paby/S0Y0AOwMJs6eFjpjDv
1/Te22fVncSBr3pdatBfXsdHyJg07tace7jybB2/z15HVNbn29mSkZdfMivDaDzy
+3azmg2aIrBxBfcy6eGZcPTn2TiQkcuwSEicfG3I0kBDzpAVWYBTXQK2gobLY+xS
mZ2ct/7nQmtzQjxx3t29TKUOhQRmwzDaB38A968kIqNx7gToZo/fljQsow2b8AFE
NTgKigkS6QdL73USMu7IhghSrncqjGpSjwUWqhYzuK7U86YIEEc9xe6cozJZWrsD
TLx6Ydl13WryOYgaqAGX1zmV7T9oYHTZn77IgXI9bi7c5MoreQoqkoOG90zYJ2DT
6/mxT/BtoksSLu1+4yS5Ec5nEq67GDpNgvNMK8jwXSjicVp7JN8dvOX9A3F4TEcJ
zkj+ejen2Gatf/WRb2FsWpfIPFKDx5eMH8lOQzcLqqB4P72svFOIksa0Lsv3ahgj
Yu4Jp/h3ESUnrHfVMKqtrJx5Mi6Hqm2pKz798pbNIK89fUJsBGaubtqHJTelfTS3
xtK3m+zo7H4YbmQTBZpmEEikD287tIumOq9mKyVFV/bYoZjqTQhD+qhusEy1qByQ
clbKqcvj4kxQdnlRN3qoYIz+C1eKNGKjW2q05Jw3636gUfcg/yxPnx8/ZKHo3R9c
rIqu28IJFd/DwnoG+/HEm2gdbsLWQy0/9fnqPA6wsPvNp5NAZ1X4mwVwWcaCt4BN
0utgKoBRQ57lI44YFyRhwXH7bFwibDvz6d4HC/6okmApe/jBMkgwBLrK7LYy/rIe
P1/BIaFnhKDB2SItLqF30buH6eDLgigr3gPhGPA5GokXc1Crw8QexNAzRSOb31Ed
s/2hO5BD8XscwgaLy1eflN6hcIyi3SvIQxBmcJ8oTstTEGxpumbhID9wlytwWEvQ
4vWlVmjBe9Zao0jrEP7Inmu8dWbzBM0XWsEkGFNwcIaHlfWlCs8gWym8NNMP+Jrd
ffYPGv40ntybjiS66NSCK4sFzql3dHpB7unDNlg/k58TNB9FoRo8uoyEJPNTVvPZ
gF8Xq2vrPpuKRd52snoZqBlazFa55+fg04K50+cC7Q2YywRMR94bZL4Q21qdjxWM
lHoI7W0Ckwxp/VRxuILSDVv3H3YVndhpqqa/525nQf2xDx88TvnaadlkHWugpkmu
yXvfhL4Fi2poEPKlswAdJW9zCbobdOacnmLyWtEmRcaFX5Ifl8TpD1Iz9d5JcjR9
e+I3S4V2hq5wB0h7vthKIRyoolNdcWJM5PKaqfHw/5vUaiy7JSYogN9GoU8OXg4D
RCjSfb3M0n3udPPs9iyoVhxVLM9QcvlUtD0hmgosgkHoB89xxmsUAO/fWDJDTTgi
sw/G8rM0qHFd5yzZidzxWyMKkbCheh0bwvidXab7vHbWWKl21+ekvouta8xlUflV
KwBKGXinEbtQ7JOLnbxnYYTCR52fu+q0D1cuvWoapOAb26yt3DdFJqkbVEAXhE2D
iggMI9stWatcUe7B3gwO6i6afXFl+q2l0dRsJ2vmy+hxtkfxWhA1xl1/zCXfd/1z
HdxUF6f+yPxlEG5xcR7/6gAhP1D9LI1eIxiJnuzBB9mm1vaC8ZUVGW+GLFE6W81L
Mo7oyNwyU3uEtAv+QL0U/MmenzXgsmu065HS72VSi1kvkMw2KEx3ZiKQ+Cq5l1rs
y4T/nh/gPO7Z7fc5P1s3XPo9XtTrqfcKrBzcXvAyMZYWJlb9e1edujcVys/WBMpK
WgRYlr/fl7nhtBXNry90dQg5YWumD48GOMkItjkjdX09+QtYlvP7GH6B+Dynbsrj
nl3O1L8CAA4m92b4/lSY/j5B6lGNGKY4QY2Z9YHWIXX9Zw28mAYK1yQ6SPNFHspr
BHzM/Aq7y45sdBmvkjHPRu91aBF+I+i5TWL6k+HMdc1li2QAOB0aXLh80c4uhc4O
28Lg9CJM+QkQbkAfjQhSodzYb9Y8ouXIKDE+SGgcDLF0mJ35xBkvYeL9UnUztXep
Dfyi4r2FvAKFW1VhiUFMsn34Ni38NA9NxoqOcK/j1r1Wk72NdKwkzgoSFi162Jq7
PzUCWLxnDNWSeRyrx7Zi9cYirkMP+WAB5YbwLoTue3kVnHwPbBC8H/gUlKH+h3eV
Jbfr4aMZWkDqQdIPFkBryeJZTRAT/br2Ry+9D2sv1vN2F6KsruNdN+u540drTMZu
MxBANezZrMHTL3sY3EPeBCAm1stAo1KIU0XWb8pcwCIdi3gn5TMgkJABXjzzhO04
WIJsfreZlUg4TdJ9LB9YR8EuyArEg0AMdYHtkBj7DP2c3MczPauY/V1NeS+W8SAM
vTwXlUvrLFGVFKiTdc4Er1wdWhDJ0+FvQKLLk4VA6EJxNc/n96sD8XMMERUhlz4m
34y7qCCDfb5EFimDO/af+BupFsj0ACA1NnEYVQQ4FPectYGzhb4gGEvVTB4AmAHA
7sH4fBFhY1mae1pIFPyBDdXtTmLue/bALllNXDyZkssJ1EhrXJnpKYr+TehmOeFt
p99OoFfp8y3VknniDN5LyJQxKGMBm6zgyGhNt4jEsSs9WGmjsesNz+wzio1p8YDn
QFhK7kbDb1HTtg9TNtX79DYM3XoSZtNXyBxgx8v4HWZPaMl+96AyuEje3q2OVwEO
h13DCzH9nFwnnMHymhrx0tDY8VeEoDnFWkhIz87hmA2H6OCQZJrziXRaboT/VTEl
OlT82gwrWdOrEWbP6no45US6VGc8SUNy+nmNxRKk9SIzoM+kjjITpdHBxheenX87
sHsqluSusFZ3SddSCzVbnKwBAFqhQ0FigGv6Yhy85HhvyVTcrPIyP0yXkYkI/7bC
L+LftFRiI7rwHi9XplMvhlhJ5UUxgVDel/X+euBl2GAxHPGSPT5/7Ja0jelJ6lHU
Yz5JOb0T/gWXs0ivejPYvfuXbqUGsY5GzNo03zPCsx6v2vSGCA29+sDwRrT9mEU6
sSryYvE7/1z/8hO5ypmIjnUQYKoKVattwevR+ZJ70ZEZ63XkS5IPAq/f4kmC33mA
c29ti0uAmLOBK8v56L9IWJvab9+E+cNPwJmpjM78QB+WLJS8akDtEVNWjSD8JOkX
0iNWxyHfN3BLQf7PuVM6v3FZjvgQ9CEeq/jiq74xVDFOoX+TjR5PMVzjdiGeuoSu
e6VsyNj6cRbSCKzLJpPvMgjJcFDoqDyeAOOwTRpxq/R4n0Ygu0LNdWdok2rkLjlj
FOxhtPAQg8oqZuMJIRhpR7Hw1/Inte+XHklraRCnGr7+jG0p+1LEU+dzCPHwjnrS
mJ6yC4HVYDphpMFGvJj7KEYtK/W7Un3ObJrWGpVB3s3fI77QY5Z+0dEYPX2Vr/EL
eWOAkqOry6omKCDEFRUeyox3qM+0Pd/qnrUbJljdzwYXTtpXt1slrRXInfuRfDFh
Kn2ktkY+Bvqpq2tp1Y6TeUe2nVNXGBuD74SbofzY0EDD0DZktQesPjst+T4ll3VM
U1fEL8QVZrTvNj2T+m0ThP2kdB/V6wgUrorZM5PzQFqiu2/BxpOyMAuKkfSgyKCq
LPDKGttugctXRDAkOUMW6gIil4lvxlWPFTsaD9zpk2D6xkLR62S19X5Sue25ksGa
EzgSlyka+5pDFa/OFkP1FSTNytqaUTrxsbF7gQZO87rCwmfOfMJqVm7O+BrQ7ULr
n5cw5be1OjBAdWYTmw6c+n8ume2lswfTrqrHmHjp3o2/ouozESG1DnS4f6X+pWNO
78Y296i6Sq5tkpBjiE1zoNql/I2OqGxylXBm4t7WwETCM+cPct2feZCqiNQUO2mR
3njishmBqYahQKanYGg86cyfHczzI0IN60H2nJ3d6zPH6rOL++DnM4Ta+8wi90iH
mrBRGHiE+rf5kbmDdxa1NqfMAKJ6G43Bip28cQWnb2dGsgq+ip833+0LW4qdtz9C
v3GDnqalI0GDDyjd/u4R7Z6maDfwuWYqKKbVTEgKBGeSrvura5de8WbVzYKqDuTe
SppIHJtXXIubRDgdSIj2VelyDA5csFiuFoRMOZkRgqJnP7UgdBAm4zmjgQXg0vyH
nfpPGFnETUnHfpyBNz4qtKnTjUzL3RZ7afjAmm7eTRxCDdwqaYr0h3jW1hSBTN3x
u5Gl/dThriHYMc2Q9RqHS4cJQDjliRa0i21+Xspx6ugW0Cg3j9bnwlz4ZfR/BsUF
N3UMkhma7lReqWqY/EpVjFkiVDzwJVBBzsOrp5jAF5EEknkvXZtLbD4q1brKXhUm
eEXERQqZdLG+Lbfu05qHra/QqGPwmqlXVnZy0wM1P73ga5S9Lm4zgGnTemVmaVHf
V/GzmcD2WjULPStJMnYU0jcSDKXeT2iq5Hn+2toGI5Og3V/+XN4378I+HbbsIcEW
sibXjQ60IxdH+wRH79n28Viu5r+Z06hRSJegIIOtORUEYp2LXl94AK/jnD1Simmj
D+9CIzg4pR1ROiFNmf3OCgECEVdMMi3rL0USS6RUr2n9Dm5SzdLS47kVWE3tgx37
DMo6Iacta80PA4R1Dfc3T25cw8HYsPnHEWi8qb7sV7rgoTPmWH18zR7Cd7iTp8x4
xc3LGfD6qzMJJJNGkNLBKGYecx9ngW+xg6MdZyiAwan5FL4M7Y9pcBta3GUa6+CF
Dg6T7loPPby2qUeay+YHkye7i6Ntue3nIg3kcFMhwSVMUmAqHU5z/CvM12hqnhLc
eG83Ve1KyvbaCQD9Lj2hJ6R7vBwtKGaOvest1DOXq0+ZL4opfspx2fP/qBf7+5Hh
7W8Yebp7ck0a/BXdfyvJZVQzv2u+ec8o/00af5LQeVZRi6o8aKRlpi1ry8xbfUb5
ciPSePFKZ42+ncYJMyLd/ugEGc8qMdMbk1EyWhNCrYIpNolUPDViVT9rm1WW61yi
KrFZTk7XPeAILGZeEknpzugCUS9a7Qy7jVQ6Fz3MrGry//JKQxVJOMjjfcnRKqXx
GOd2cCTyn6qgI7ldMO8CFTfLmlIMY+VVFQV4vLuTUVwyTmmckvqUKlP+ocKiHSl6
rZwM0RZmTmDNOonpYW/Kt2ikdQst/gCnGp1Fzeqq8DH3SwcodLP/kDgC97uuhBsf
1fYycgu5iEEyqDj3GvKSTuf5RNl50RG8SOiBZG087PHHXwIgvomj8ATdKA7r0sir
XNWC2tPQ08+s4sC8/hJl27M79msS4HtI7Ipx44EfbYM2Pg2x+YYOZUFoecUqFsxI
Bd5qY4aWMyW6zRsiovPWH4oTpNAUeWDyiBL8tEAz8XQyzPsNRErOGbo3j9Rze7r3
jPLPkvo7zS5/u7e+0aF6R/vtGaYWNVZNBYRQu7SLAThImRM71AYF67jGvSkfsbSD
kJ3R0qiK91gNQGymqvR7+5pqDJkyfCywlhXsjY1IyZfXjyxqPxXu2SdthQksRaZC
Dl1dxyvj2qPnny50g/cSTAkDrCfWd1qlNj4eq/un7+RQ4cfisX/HTzrsJJERXM7y
DFj8yOQjAFQKjCZEJdkQOcezL2KfqRf9zblH60DuhzHct6ewWWixEXcK+dz0BCWd
HujlVkUAZ3Jx+23cCDDthqwQcIRaGnmCjXf1q+2F63o7qZmd8wJ8x499zoThqgmb
+OXXUHWP4fB7+moJbgenaW5tr2c8L6D2bB/nsRs9lo1D3PvuIciLSR8xA8A9l3CN
/kLT4blf9c3XGZKwXthWyv/6kMt0afL0l5Ooa+FpgqoIlJ2eUg/Zl7XrTD5/4BlD
j2ggludwy9gBbOKv3iwE3EUXKxYj4n9DJgYvgelyV3BbolQw79J219gTjDJSUofw
egg8hglsoU2vCKF7PXXGSwzoInY1fpn5Iq/AUtGiSjA4rHq6kh87uEJPf/OLDkUv
JHkfe1/QqpEudZf8hBdv9c1sJyXshiXkuQ4zFvms2QeOj8AgIGh5uP3Wso59tkkA
vFZaAkdMNwgLLjcek8p/cGFfriSLs+4e4VIERM51435OxDf8aCHe4Vy0YMuQJwBQ
s0pZdeQhddgZNLxmGBSxA0zcj7qGVqMmw1Kh9hjGWiaQiH0Nhz4pcmblKBJT0ABj
I0Hft9dd3T3lHcJeGLSzWJr5JowOhULd+g8+G5hxyszmu4hPiMoXQX3g1pkWJ4bR
8IHldlEOENOTg6KAqrHFCr6u1XcFOrvAgYY2SF/oWTuVEA8TJA4s3z/gGhBiRQlB
ZTdQucdupagTmObWh0fEEWk+reCQW8sMFGABSS2fwWHsCtd5Z7iBz55JpNPHx64y
Enu5T0yiDJqfJDUqGf7kY4q5r6jEGgfBr8r369c/jaGCrQv7vpa4rVTzFIgV6mdp
ac4ZEY8dR+83ZNAJQEjaGTGjMReZa0DRLJ8EuqqSenAey3MIsTd5iPqQHRSh8taf
e9XhQXeyoGDLxZZgEzFuEeOKln/WgZdN06/Cw1GDpqmObeOr1bTTs0HNzkev5+GZ
wb6rG76FlatdeUlvw1G69aSP7uC6IJu0XeOPBwwegTfFvQJIEa8fr5l/FfYhJfSG
cVenjDho9lkMR5vZTjzCAL/YrysO+Y+1iS7RkI+xAadbLEpufBSLmhuIRRAphW8l
c3GhUmMM8LlxkYLWtTw/tV30ktA09X7+jrxMcAniQlQnZFq5tT0ftOGc127onK9v
cG/yUW+V97DphuZGkkvXJjE2X5divCRlIdOkPnWNCjbYQ4Zv0fIAUFdLTKtniBNv
MNkuSjTfLmw1Hk1GqcVoKrUIKMXCbnZxjol+2m/GbIWOisyQgh3TUnQmWk1yXYlD
YvpXE1yaPXc/KpYTsU1aEyM2ySTkQUYRdGBe6h4Vz4DE8bsiuYzdVM5Pp2MnTya4
en5XrVSqsGbfi0yDH0FZJnhQaOCXTIlIziePYjl3+oqDs240ueN6715d33jcR5kE
K9swMj/RNL0h5PeNyTzLnkf77d5pBF9mWyTkhiYvus5EYfLexjX1PrQWIJZy4Din
LlQAajmVze4eidJlEgh9R3qAiOP2ONXwmQN8mcj7Ue4r3m2P6KmBVmE5/5qWQ7cf
ES4pcGc+rPFg6LfMDF6P763BvYUQ1b/GZ25lvO2AvasREbYnXXZs+JfiJrbFCWs5
XmfZNkKzAJHyAu42EXRUQON4SCUmYCOpv8Sjsm9aBuNjmnXh4jz6LhlPTYrfsEUm
3TyQDjY7sgVzn/DLVQUG+QrdNWHeHGSe1pfxwEEP4qHJIG8/SfPslsZ4kFXPsCWp
rrpLUVX7LhLelp+ZQ84MkNhJc0f/JPczoH0w/EeOn3lQoiU+NVe+8rEuBF+UdLuT
na8IOquhVrIYiZlTUKIuvRxL//jEpxpsXCyRnRwqR8TJrb/9Jh6wY3N6YR30fj5U
ZENsJq+q7QcBaLWHXFm7QEDEEc1IjhxrGkuzfgcIvjHkWUKCaR3AxbQEU47B+rnW
71jZUEfs1OuX1YadITtYcOu6itlXH+eHOGhcey1AEacVtnUDXpnTPOGa7N8E/m+A
6zpnB3iBZcz9JWWumVb9ZQgDXrkWyZ0gQbH0pW1FymP0/s23E0KG3V41OD5u4b46
FJQaNaAeMyyGZpTSSZK0bRPEwKHxuxU54wSmqwzFsMNDO/G18Raw3zMBvMrjFsq/
yTx6mbPWsTqcLRm5eV4BOOuHR8dpEDvy5++WxiTRkdv1eBOPjkOfhQQ8q5jtWgbt
Ou3jr0Wljv4GxfcuJT6SB+Gg0OI1l7xiQSeSZJfZ09yOlXnFzQhqVZ5Iy0+QDF3h
ym4IvI7dTxRVn3DafHjO/OtLuLDr6UXMiJINpszEaogjybNIfKS1mg0F5uZa7Llq
5+psXdjDS++kXyNFq2oJCC6edVSX70ztv/jAjneIsZcvFqdrOZzd4x3ylJ9RGhvZ
MKGZszEYI+rdqMJ770F44Obt7gekEkq//vZVsL1ty9DnN8xi9GKSMbQ3xWGu2gRL
j1a0IXnwi08foUsprCVTbAsviRtjV5P4dwiFdDPWAcFjllpw2reZZBphnXH5dkrj
a5jqYr4Z0HWDHl3GO3IKXy+y2J56Ed5LpWyQ/MtONYm/fSHMbHIExFgrKP2BrLnX
bo9PLwVt1L8xh4FaNXTKGPScYR7j+lJQt1bGJJmINCNYsW1UqryaofWONRtSJLVZ
CT9alsUH9wFq15A8798+hmYdTGoFWRT9qfglVGdbOsyHwyiCyGWV2E3lIyu82z3z
HP25HJ1W8OkBf9n9bmmcLmzZS2PS3k46kxDxDBpDVIFMOmmCUJBh+A4+S9Odzn6r
SffSiOrj7ezry1h7+ZsZ0F5jPNfYbPTP4GWM1k0MAeQKVl2t4gm2AHAB7tl7gHHM
DgeZcsr49Lhy9DjekahuAEz30NZgVi+faRT18pMW8OniIQD1r+6hhFsZY3eFaUQg
apyDEY7t91NAa5bMIXSo/+N0/WeJKvyd509LQTr6VZrsl55CPE+0xLpXXANiq/KR
i1+JlPSs0GEejAe/G2oVUnJnbgVyr2SvXD84k+CffAJvzoOr6TLguM3zH5tPq5AQ
fSyLVHV99favi1eHz3hUdt3oHqiWdUh1SRQDO/M/QO4FPzsv6PYDwxRyGCa8wJ2I
hBLicEKdof5HrFntaHP3AtDewvRslSXG/wmmIFzL7xfraWTtNZ4pVSulaX8I0N7N
5tOkMNu+X2qqFydZha6TgOUryXwxi67wBfuuafuiVSnoNKSpk1aei08G3w5gu5d5
AvP0GyoYolNs93aYnclNSK6/8J3O4wm/NZ6lebtb/BoBc9LUhEJEJIQo7TK10A+8
9fEw1b/sdVJHcVD+OVVEnJIOw8WX1Ey9UtYwCiyQppGKZGbY7xETBS2Nw135elhj
NoX+0QfVSR3VMfz9+ROSBhyjP7dpIsVQM8TzHWduUgOkMJ+6X11o/4I5cy5dY5oV
OxOIyfjmNjDHzrjW9OtVZBlPcScVX/RYXd/Bwm0P5HrQnXazsedrIaWg7tONJBiR
dER9JcMQCV2u+rCn4YVg32Jr588JvOqMfJKeKenKZLxTDSARMjv96AWnj6mvZDbD
keYBkp8mmSTL10sy5hCSGhuALKiHhjKHWTdTDWNwhusbe5Y+SHoIR0im0OtYmjD3
1eff9IceopL1ZxSepniO2PeAKB8jyuqUWyOWCwFX88tzqp+LjFyW/krTI+74J5pz
LrolYD/tkLGidhc8D9NasjoigmoUTrNxqpDJbZRYecgYdAqyIvuPeP98Xz4G+QGV
Z74OwSydcopzzC/0rpO7pZtAZJ1V28wId2UL8pdSnLJutgwXirLtIP3iGyvhKSIY
n6ewL67iVOSx1mnvysPNS0mpH6HxoTg8oWvRLY16asjG0iyAbQDq4oc1CefAAaMh
m6E28jjpF2iP4PDSPedLrwtt4f+ASdeBipbkT/APJ7JcdvBr54JZIzBaZwWFk3zD
m4+/QcAGGNVPCAK9E/Wu4Y8l2lAgHfpRayeRw15C51DeOuxdkeGrteo6b1tdQ12D
SKxGY0jCPd/FGosmwzcP8w+U4bcNobkyIpREFd/sIVqZhhr8BjpTt2fUC6A13Cxa
Vm2ghsupj9OAthHGjQCW6rkTVWLzahTMJ43e1N2If5WJiYxMb7Zcwb9jrx6kt32J
Kb4DVktDGAAZKU2J/A4WHch1mnQRIYIQcBk8EB7dgSZ3ADrbDVJKK7jcTbYAFOe9
tLoAQfI9McKU+UUoOdoABXeRC9ITKQKsVLpcRe8yfkbmamEOvRPBtkb5fKUOUiJu
J/+C6jYmhpwUrtmPALmsvI+Y++B0w7AUvFZkABSerIXQXbjXb4czZ+bjvUxMzVkC
62nRgS5dInCGwc+sAbqUDTcHGg0d3tULMSWoeOHqpHkhH0aD3/6vdIian4UzV7Lu
QR8n8CTuqiIgX4hXIng6T6wt3t1w4oR/2qXNLWtyXs3kURlOV5m2PVOsZlR9+3cr
uHAScWCrPXDQrAeXrk4/fqgj+sDPV1ELuBCPk29Lje2mctbu9jKyS1FkQDROsrSr
IOJNJ+BfjLOacaOvMpF2or6UG1v7zB1fifGICR3jv6j+0Zkz4AQOeCtB2rzahrYu
YJ8CTzSrVvXZbTGCw/1GWGgvAh+khTaq/hE8gqjvGYFtKnDz5Oz9GTc1/5zElUDd
mzGhuSU2IBxKAK9nyW8iMTZ+yxXsSsKJMidY08kWbYrgHvS9SwVnuKPO+C2vdfMl
XsfXwewQjOIn9t0JfuSMOC0UrDsjGcl0vsQfGBHrRzBkbhrtTMGIkR7w2e9otVNj
v6MdVlfkl6nhYqiZ8sQz6kJqxo2JBNoYs5mAwCS1TYlmRNIquURnbgcSPBehLvAW
zJoOZrqT8JmI79n7SmSLDu1b+U8f5GkGVPvqSfbhQ9cdsKQlBJBFS/pOVzVWtpMf
Y4LQ2o6cvnt9Zs2CHAJ7PZhXokp8gkCPgmKZUmiz+Uffu7Yq6kzKRE8t46uVCeyk
dAMHOjGEPPEuNS52JnVZbSorSr17njhcD2LzcnbiumpTdThESJ/GFvBAFAtx8wlx
x8ljlfQrophRgY4HkjUvi4CH9tW5F+qWc1WR3oHYT9htOReubSyg13wrSI8R9aAP
16ZHDSepRFPGvoOK5ZGN0OCfpuu4SfVSw6t5QnZaeR/ubq9mK0ebmM7PvuT502mV
YrVthAXulBzIz8URa6BCKHCX/8LSnpK4sJMIQ9t134WmS5KDIeVeasOvoUcIhsfu
TKn8Z3vvN7iYCPIhW48Z6U90ulV8wlux4MvUtFcwWi9wI2WbrI6Cm7fkqVpCDHC6
VAhVu3x5geoqXL6WjikB81C3XNkkyPtoP3DxZwdKbaiL4lO83/s6da5y7Wmt6Otn
kQXj1KPYZOhNap/tfZKfsGfcnVMDYVt4rdrVX+hPFraCJQgZQmqbR1M1PDZ/Jyzy
9EBc8DdpjJsPPE4s3RfQ892M7h6kdT5TDlGUJdIrmJWdhN81axwylWUiJGc64mPZ
BESTdIV6C/4QmAjs29BhB9OwDRsb6yL5I27P4ZqdVQW/nKVflZwMTP9p3XZOvrkK
t2TZpP/glnk2TnO6n1yHXiZ7TBVkIh0KMOoBVik+lC/Pga1M8KrfAAw1Rg3ZIxjj
N+/x58oivmvxwIIIOE8bKALdzKENaAy2OspUXGyDckjdf6MzISc7DUgw40EvA6jO
wlgPJwxc+yYXvPIz7qAUDdEUZYbAh2ZQTWtCRaHI0WRjKTmieU4CzIz4XRj/x0Id
e38cXsTagBVdNma7t6G4fZn04S9csuoW1pU1x5V7HzuXmfLBSki9ISy19E+sGg23
UbNsKGAakuc2FLHmkot+XkdN++03WlVkTh1NsC60Ly36Zel2k3Z8l326HkYKWOKB
9kdFqK2iGSsrNpXGMzYG3B69gTI+jpJZhyQmMPxLC5TiUZFiQr+ZVreYBVQZW6/H
to7ozjO7wqkMmwKL9LJbA8LLTw9N50sNENMu+0wQQQtL5QMvEvkcvExbP2qfWTxX
mlP4YsAXPeMzMk208kLXENX2TZqXaL2vMqdPiSreGhMeyo0Hk6Ac0odJqa0tWGUM
qH6OuuY0FPKTBYG3F9wzFWRq7rDEVBEfgQggqGgFtIAvqnAYmZ0cUj2vP4dhKtIz
ih+En1a2FvajZmz7y+/9mi+j5Zm2facbOvzcdqsaHshYWR3lbWpMjuNRJYPPUwv5
k7v2uHmx54S4nyYD5mHTE/dYwpgiQdvDmYYDWr4E2bUymKML3+nqBd9JHErez6ah
Fb1Tko2xB7TfNXg+FWumNG4Z9ILhRJVx8FdvI3Km9vekCSB4hRYZbMMStj2NKCSK
febHzfrGJznrizQ3QhuDr/zj0GHcD234OkMWcWqkX+esRkRz5MtuN3FD8T3iJ1SF
jsN8nQBU1v1kO+YUXDvcX2dX0cAqDiBOjGzRvfVdsuBYIdT9RXDLol6nBXChHrzB
Jbu/xRvj+Fs8UfmpoIV0+VnxvYA8ghbNVypbNuNbz0JGZc/5uCuXfEtuAifkP38S
LUc91SoLPe+fFGDyIUGZSHDHnACGB8dGKBoBSTmairfnudB4MjOcKC19QljI/ADC
ZFYqwkzbcrcyxe0PvL2Ht8QisKZ+8eHPPifphHJCtTqYcM0q35mV2PsK/kTGQvDZ
FiaJL85uzBg8fdloYqwo2ZgRBe32BKn3rsPqtWxonKm3Id+ks+UR62nfpN+Kb430
sFXEmBKK3NnONNhQ4XfWv2ogS6xy2usu1WlZI+sR0NAbE+W5U5Tf4Xx0xb1tQbZZ
x277r/tizBPP7b+QjMDIIoGm59Ns7MKmy0dzlTmAEUBrFh/8SVWvzWlG5Q9KRUZH
WjZ/C4jGOgH+NX+FzRY7jaGFCykizTxyDljO5npE7uwc1yX1u6rHvltr6Cw8QjGX
H9ZZGSwaSJ9ef/4jOfqbi5n7EBeHk69UXYSmDQ/mpd30TUJ28EnUet3R8ks7GP92
XLF1qje9VLwvukmAYWr40TpU2KC+tRwahbknLpSilXQnpj7YXv9LM+cw30TpIiuw
1Vz9RUgivVQWXCQ2tqvSo3DqnND6J/S/ODAnZClRZU+/GJIP/l0UfQpPVk5yu3Cb
Ds7Od4v59Y+i5CyGPwvrorTC9AIUT8QjDzjBAZaUGNijLd8iWzufRi+1kuV7yZNL
9RXyJL2OBuXk1afKkMMCmtu9N5b6qGKIhbWVDvH37Fa/75AoyeSYfBqcNnUk1/rn
b7xHbGY8o8wvvKlkrGKDjsu4PCo4Hz6K2kRXGEnlbK/tSgXFPL+KkO0i3usKXYVc
bm5p+ZJ3YYTyII8n5rGYat5NTYX2L+dGyfftfQBcx7qiXWMU1QTgFORyq2xqAUNs
8fc5JqVOtWtNdmGLur2xCZoAVKBgPjlKYDegicdPt4fV5CikMYjXw/XSD3ALgLu0
LBMT9FxTyr/8zR82T/U5ABfhGnhwcvOMybIybwwAtiSI/q7ID6KSx5imxdkbyrdS
/8vXRc+ds3+f3DBDEgwob/tpnwgRhf2egJExiGcuOOVjIJvSsYdDZd0QATQuN+w/
JGLRUJ4j4JC8h1X20WTQG0+fhW/9KlHFW+DL9uk4dU07rCtE6/HfhB4LsZhSqr9n
EgLT+jV7wSIuCUOAaaqFs2vYUFnMIrc3U9G+9DD+sjdaFQGJz/lVRW8ur7rODp6h
zQ2+56odm6nFkLOIpFdYR5TfmUdfwhH89MxDUbYqEpInoFu9TEA/86JzP30P83am
hmXKDKf5XMHB+74D/bKbKnHOpq96+woXYvqFXiUzFeqiXd5jnMIz7q2bcYLZ1wwa
CdDIiutgXw05u8WL3rAxL9uqarZwe81IYsBziEG2YUbcEyvsJlkuj/0K+AXn/C4/
nw6sf3ZhTc4QJdlMZCs+5Pz8e1J/8auNdH1lYjIaW7HV2zKLHEnWYRHmQ/TwSmvG
RT1ao8nZUotWL81ZVYO4yfOjYU0CRqfkSFVUP3jzzSrIXyMdaObfR3pIPAxqnhuP
cnVnBQJ8eUkq2MJCQrnopQW0wZkWIFX7n7Fvvxu5qZpz0rt+kQUDNC89Yg84/3uo
Dc3AmVupZAjqExmkM06ncjcC6D65C5rjhPWze+4wXg+sH7X/Accg/RklnUy6XXBi
R8aVuJHIXWudxCJO2akGDvkiG0glMsE4YH1/eUHbDUFHkdSHosl/DdVkQvRA5Vou
rNcFp36Eyd3fl9hO8fas0ppzuEzc16SLFyWNmT1dOEPlNexiBIf5YISOGwHMF8Kf
iwTVPVlg+fPWjeHPorBOgccgS6LWw+AhxqlimUNRdJatY9z2PNUGeutsZa6UjgdP
/DbkcZy41T6lTdT4uHcAgNJXpItpzKFphEev2bWidkCmj/OjfRYKM1aNLIsSIVQZ
oNsg+k/8OWWbY9JaQUb1XxxaVoinyUZW7Tab+7W1khLW2NYlFpM/Dn2+mT+zx4Bg
xhkLTzZ2e9LKInaN7fA2D1CWSGAzNAdMXU8A0gPcjhr6nERsxcWcKZ30KN+JnVxl
veCHFOW/KxuG4XQo3qZz94YAXb+svvhwmO2HTyc03RXky2l7Bcxb3F2CMJa0G/XE
hMZYpcQWSMbAsp8xIWW5xgYn/NVvjjErmc7N5yEB7SqeA2wb7ua4BgsyOZMcftcY
k5e9IkBpW5o4H9Ux4ipgbfn6R0cWx90IfqcGh2GqJSIN3zG3VJDoUkyanSxDK8ac
kxRzh8giTiVuUJ2PM/jntTcAtxcoTsN4Mc0DubPX8vq2iOz/1xKugf50fAaD1Bd1
Y3eKyo3n4qdM2nWjMFxb7ryWtbQzlmrhobbUoyEqcsQpntjfWPTutAp0s9c8mN3F
k53dU6JRRsIN9KLRnNbLVmhn1Rrkra/Dk1aHHLJIIUed1rDxLYU6T7KFaJsC8c/F
piExw0KnfBqx0ZwpGBweDLGUvgu7kbioglzeiuTveWptJEG+mCed3setLDU4+Mv9
TckLoEusKCbjlWesyo3Izo6PzBGX73dAVCThG4FCgD/bFw9rZtvDC4A+4SxwY4e+
6j4dvYhz5oiRsToXFVeu3K1Q6GXozDnL4A7plDuZBIRs4ZJ9roxBgbWY0l5MzQad
wXkr94WnVRtrqV8VXm+8rXC9nAxQhYB8jHrD+ErIZEJgTe9go1BB9AWSccbZV0Yo
RDSvWRmUynPbsxpnPTQZT/K/RIQrt5eS4mlsSAqtnP0gxCIAqiccAeWz0Hqx+kaM
xeK69zKidxdwVOFZjiVtRgaIJugO08lDNdaWTxStaOhlc7aK+0jjJRQB6vk9W7XP
IQhdxTlkaQ58KDLOqts8AEAgzXYWCTOE09gktNZiSmTEsr3qwc1jkzl/E6Vtq46i
QuFEne5oJue+qcMcTlHHbs1nt8+zwyQAsyYvx5apE/owEsn9DeigdameGxtW4n7s
qGUVBiNwd542ugr9a5v8NyvJE8eYjVZIwVw8zX7W9lzv8zTSDU1RPwpsgwGs57KX
kXx5sKIsVqfXJ4sWgplnJ9GA2tQ/a/Zc2JfByJjIUajaH4XWpNo2Mx3isGU6SYHq
OKgbvZBRzAh22al8UGFxyGlfssPylDd8Et7NSXyIXqPvxN7BAXThv0q9rCRk7UG9
fxLeX/hTZ0T2add4ZXPmnwOll/pO3Ca8xMZo0bpifKCOzHAddMqVqhY0puTu8fNz
LvafR2KxhZvJRRsBNp0eZhR0iBCAM+vWvyOhNtcLb8ePaOtQoJDpmxrT7I8M1itM
zjQP4+iFEiFrOirvC1tTZ39yMvmRWYV8UITDCr2BUtqBUCcF7GgSimSFtAc6IwvW
tpPUOabeSWkcXVHBjqaTUrxrT5GRR3HS5mXsp6lNvr7dtYhLm3C254wNQztx0MPc
DYgIPTbc+B72pI+ZacctPxZdHQzER1VsEOzuJbONMLNNUHji7PXm3NC7RsglU5RC
eC99JbSxYMab2Z0DCO5UR5zSNqUS76huNIzGaQSGBrnbmJ4hR+PgdwyOweEfFGUe
qe3oGECi7p5K+Lm2F81A5WJsD7xWZ/Qm1CEjwOwsMCpqD2jhjn8TxJFe/0/Svro2
uWnNZFT71RQyPlLdp35J4YorCjEvmqjJKtosf7EgLIaqvSqkb5ierZJjlHY28H2/
384j+ktrQrpdTU5k79WBXmVe84A+iZCs/CC3LRFM0mLkO/zXQ8DFUDZVGNX0sV0v
0+AxvUekK4FrWuBBlqEsiQQwTi9ZgUbp9mGyDxaLGSUnl+9RUU0cBgzChMPU23OX
3NAJzlCXhsbOc2wKYwREsd3+WSQDMrQgL/Crfx4LiFBrVzZ5MUejYyN9Om9XLyTF
HNolWb13FEYMdn1bikMoSQnUN2ACU97ViaNh5SoUslQ4Gf77GUmxtmnK5gIHeW13
/hmmC4NJDsVBbeLWXCPcCHx2bmmwtotiVfyUwAxaXATTna0LrLpIVjcOmOzgAwRb
RcMARZySvRRBiFddWnIytIzhx13BFPD75ztYpIhQWab0VCXoAMFKifWV/LMOQaFa
VnZcKHZNfg+Mz85+5ijWelobrM8B/nX97t1GvgyJEwV3F888dUqD2R39RmMNra1o
WXuSHgz1crDKarHleCxt5hgRJw3h0fgCj+pBCDfAqm1dnESqIuoXt/Nd0/eRKuZc
WTwFODCH2FwLzhZ5hVog5yIFYcClENjOVTTior55Yy3auNy48tCp+k5S1e4MKS5U
Et/1K6C748u8sE8bhc0Zhk4p3eD58LuEJHwFHLF5pbvst0/OpUl8KxKqVrXIH+t2
ZO1IlgiUVobzxBI2aF0VvEN3uw0XGdyV2tZbc8stwqzet4iolBCJNT23v6HVKvCI
DrwHvRsnzq/tlrd827ifvH/i1Kpesaji5cRr13XXpzXraExpqCWA3OlEJDQN2jtD
Jhx+eVbPnxap38EUD+33jbmnrspJC4l9rYZ0qu+GVaSaP/kQUKFiIYQ2wmwbHdbB
32/AAY/tN2312hFouXQuDOiIsEKRIpX3Tc9yjuSX3gAwfpcQl/HfoyR08N6MfRkt
fE9LWOTDkDDKDHqJ7/oBioYorAMHHPSpi2qfw+MQM95VapPdcu5paaLcmyT7g/Vh
vLzXMKl1TSOXukTUZ7F4XsM9/B4Bh7DxnJADylfJfFJ+c/gVrkdbVqdbCMX71Opn
Vkm3Y65pxQJ+rNmZ9iJ4fq+r1DtT//l1WYhpuXcUuOKYaB6HWLUb9P/eJaDBg59s
ODbdw0Oa14Pzfwo61yjQUwRCWqhuOIo75SqoelPTa17TNwomoSzHoZQYuknA3N/8
5dAbuVh6ux3JTJLqj1lCAQgVvisnJMFDGLYtA65TJw9yje3dMNGjT83uVBV8CEM+
HWcPEHR71Rx6UPJDCWrVkHO3Kbf//BEU8XtOAcq2Ms+ahuDmK3hqqIpxbWTNLUky
o/eylSXmfTQUeHBfgQXjh1u4d/PnqeVksfiV6fsVVYm54vCyc7cdDnwwv8zIn6sU
7KJ2uw4B0a0Jk3tD2kXoHfW2m5nGEIOkmILFjH1IvaHsnQ2cKmicGZlDYPhF6tOk
i5BAW+Uq5GPBgU8WYx2xAVdEQ7asogshS8C+TlG2wCJXGH+G2s8fGCWJOTTO0mln
QRAF39bhYfWoSkcQg+aDOFjYHoPNXf8+2ghqgzs5fGMbxAL7hV7xmvIXeH+4QkgK
RAlAGzgG/4kpHW6L6yg3X4TZqpxUBlMbQs9sMXTnyal+hpOeNOUtQfE0EnTgm9YG
ZKcftN9OPqIq7Gtc2pGMtSpU20ZZvo/PRCgKQLgdLKKGhXszg2jWPjpfjdwsT2oP
3vumC83QySbd4DIwQgl3APD3XgJDxMNeI6qY7p+hWKBqXduCjDVOJthiYw8qjDE7
BxitAvhr1PoSPyxXh6yByzH/EcGIUKSnfKfwnzVfh0o26F4VLDGeEbkHGDOnavSG
zH4kz1PjjE/lbK02KoqMjJOrJY0xYlr06PjgFFFaRdtVWNgLlN4nkAZEfxwBh8/W
L4XRiifU7FLoEhLTeHVxJgZnZ20i0oZ7XB7vki+qdEslyj9yLi0T6TAqyDpyLohN
KKvqiZwiuNQZuPRN9qXG8wXi/uuJvZKvKIno2q7wKsp2AyGss2/a8pSVmsP3HDGz
abLhM+c0tsLKZeY6KMpHAjCvTyPZX3l3zZR6i+wwiYVotRM3VEORxT45wO/964Py
QntRR7LNXzpMn39p2DHe+A+VdZv/2d3UeItkiKHAgLMHhNA+6Rg02CIgpsXRq3oO
gmBlg2gURDUJE0fE1MMOh/LihWjiSHD5MmqPc4n2+Zpb0M3nAdBbqgKsBryNHMEo
ZIiFo/+aqb1ktADfV+S7+367w15tSvF50e2KVLz61LBeIifO2dTts6mZvN2FXpoj
pYWz/Nlz1hUPlJmXGNckTBIBc84w3g+yZo1B42dnxvuAwKh4gc+Ef4+ump810EV2
60EAY85p7wUnQ8dePEEDutRCs9GyqASBnTTBGG3P3b9dsujtQstsoICoJsYJn/e0
yBazkHeVzLTGuGDXv+oKOrhM9nmoyGTWNR+z7+x6YyIh6eiWrExhbBeUHUpZ69qZ
kOZHDbUeQd/FnwHsyPiEu/eam7LCsjf6UcbpMOPrOsMTN9Jpg2YbgLMmDB5tK4EL
EVtGcQMa4VsIcnj6RK1Ujt4GKiKlToP+RkvfbmUPu/TDZnU8/HCAjVPHA5pJhBLL
P5l3asCCPF2nzQB7kMSNc6FZbSY3BFdDju1U4b8gyP7BjaAbQtaRwqgGv2+mvr1G
ib/G1C7lW3WOfmi8pjPp/pFoxX0GB+DH9YOTfvMfADPHPZ2hL/E0DthxbHLF8DiM
+tiD940Mv6wd0l6Da7UXgFZE/NTzOZvbfOGldGyxIEXyKG19Srq5bHxUvIVD+FAo
cf1batR0TRzs+SEV45pYLk999+0sByhPOUs4Q6tT6VNjwy17T6nPgBOSWcoxIogb
/gtY3qEStpOqRT8iQ07WycGNbGGMDQgwp4u6Edxy2JSEB4zR0QVR1RX59QvAGOkS
P1NgAsPCx8BUWViImf3CSHdJYUHVsPZve9EKSvda2uACelcCL0iR/C25JxTIq1Z9
sWsV/p4VBtgxCPiw++0X/10aG5jJj4Um4xpiomalTsj5pQRKNRB7EUPCtW9hNAPR
N1NXYUQGR2kYHZbkuwCFdrlEMQ4sXr3xcDn+YxPt8krMWcBMdie25tuBLRlJKEPH
Hvfv8GKhMgnsQWHYT2SmbdLgVie/WkDDshEjHru1JN1CgRPn3FN20Lw2g/RoMlfe
2VYxu+pRC2nJJFotiDn55K9KwqQrEbgOJ3uellxn+UHLUkbdS3LzZV18A5hYFlAD
O0pS4g7NX1HnwnJSM6rsViPGCMfbbwZbLJvAdPGfzefiVBxEPaikNf8W+R5WyRLl
ypuNpRR9+8Tvgo31ObhJexb8JN8sTthuxICJ5Oj31orh/mUzhukj3mYyRkqZb96D
o7VGfzxdnzdAm88gPdXkmKity15tU2jZn/l3sHpaWOvyRVQegibo+goQBo0PziA5
/5wtozMSLHv2bJLCn8iqDR8vvbXI2qU4QHCfZljxEjLNN9aqtymgWSteX6uONZlW
iXZpWBn/5AknnKfisZ9p/oJ4OCJRutbomXKNElATSLPpPt+EZ6MqSfGOdNWo4OqM
6PIfpaYwX74UTKptMqcbMsA/aH2NtgZid7VGw2u0WgWrpinUCr63KmzwYYAC8XGy
UGhkkRrWKRpB3GC2jD4nuQ4ns6VTl983cZdsuueiTEME6cJwaCogLCJPpqfc1Je2
h2a9RYsH4LShEhXcOwrykZWSfs2Kqzl1XRdhL3UFsJ8yqNbRYXmofCTG3GLnzryR
lWujCK3zwjJEYsu+oX+930b17JDQSeRtQ0k8975wyZkZTd8oxUv0b44DJDvVWx3Y
tRMn4d50e41UoNh1IB2DoMQgZ9KWF1qBdJA0lomi3y0QixstGuS6dpbPtptXvLrp
YaKoAMrv1+eg3Gabl666m+K2g3julfaD4y3dZT+vrnJ6qjc8bZYCXmypjXkQLatx
5ZcXtBdrRqN329juL4bSPV2ohXXhnY5uUfaZlmL3UJqYRw4qVBE4MrfF2TNyQklm
3kc3xT43ZDLMpjW9NF88Jqx2AuUPKZC8f78qGp5GljXZNKSOHDfWnDfIX26CvWBm
FDIxxqW1g7x+7NJvarELqzPujHXZCmrcPDSITw2k2KxxtjoVpA5JhuVOZ/3Uobnp
T33h8JYmfwUweTkfUOOTdzEXHcdqTFeVzTe5deJIu7sBw+CkRHf8PNBD+dzCVwoX
QSTFvi1FGTCthOdIDzMpSJybTiljIcjus5aOZh3byfXE0/3nMxesa4AHwZVm7TTn
w7GaXVj2LwZqLvL7oOVkQG6fqXcO0mPz2l66dDXWsCmAUuchMAqxhiLqAKkb45EF
FiCjtEwoHxqURGdExvAg9exlEk4VlNrOanrIVeJa/u3bel3ZUYWlr7v7KAPCoazp
JiEWUx9MzAx1hv3Liwfiiwib3BAElyOhpO4F6izoeI2x24J9CXIHcBwg/gTFgxz2
Z3FrQObzPfLWKVMAamQLSCs9kJ6G4MW8WsiztjFqOMITNFO9sKF6oI6Vul/KE5EC
hXNW/FfDMm1v03m4aBpWB2M+dC8ucDwMjwQmht62ajIULfzJpI35iVqbM1d/JKYS
qe3igiwWaVa5tzcZJ6+06jL+UvLK21CI7OcX56mO8bhQBQKylcLke0FSwGrfo+ZD
0uw7v9an8f2m2glA+MmmMRzdGy/cKQ9HNAwGDG8CZaxLr6Wq/3vEMVbe7D3cpvIS
DE6xy4TeQD1CuWt0HzqjT3MPF2EfmcxD5xwIYiedWAp2+ueA95xd6rDRhgEYSbbd
iMJNkNXv1bFqwEYXYLKkwUSodyrQ1M8SndCdtaLHr0dGZSAT+mRD//DOusdJolIo
NMn5stZmHya7SrfnJ0Yi278MRoLndbfieqOGwk17Z+x6ZHyXYD3z00SRXehn3An8
AfQTA/zIuvrpeA+CNSBPGL+LlY10F2ynoVJ6rGF3qocWLsEjMsaRCmCUpbkg7lmE
ns7dUWmUVnBHMLPGyPaWbtnNCQA4zWKLABjQ0rOS/D7KasOJLy/bWzeetzOT8vla
Aphvz09RL5KvwfBDZFdx/xG43kVicnn7gDGnpRz29u6x3cjYsYcGorKgv/mXVujZ
uQnA7+923CKP0g7QlIr4TlJ3Nngr7JecvcH3ZR7GWTO4sonQ3o+zhoSMvFRQQKHy
uEldjOilHAGKJfztZ6ay1rbr0LmGX3zxgch1UM1thAxAXfwdOVlZ9LvJN+4fKOto
fs7AyOwR7Ao7TyJAEDq3CuNuR0+ZM67lKsZSWD/02cYtOwumwDL4VC56YK/mIohv
SqpNhHLa6MxPE0InzhzX/iYtfttW5Mx2S/ZMv1wcB/fIVKV7sd9zXG/o7fl8pDAP
kIf+JRnqRn2s4TjctMfH54f9+Dvi58mt9SpV+00U/G7Uex46cP0gNiTDvuFY2K++
DBKpqHL/sksNBwbQaGfBL20eFsRMJmK821lBn12vqoExiPgirJMs7vf3LN52INSQ
LZC+sQIhmX40TFpSqGhnYHinjIQrtfRtB4+N1SPJocSZI+qumnTr07veAPTN6kWR
CI4MEowSj55V5N4IOTcCKg4YcSuXF/J9hFREBf32EXiMM7Lzi1EaXJ86RM9v+OSC
T88ulz/0dE65pAcNM7ecjR/JFX4PpGGTYdyOHx2hj4OjkR7as2FJwSCYfCsDHWAu
QV+2O3v0lsOLnhoScI1Hv2anhkEt+8/m7AF1/N3C8nriH0ck1oUchACjWTCh8OYO
`pragma protect end_protected
