// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:02:11 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
clun3U91AVJL1zfCCgXk3hwVWxetFs0taUEFCUJQSy+KlrmN3oN70CCDdtdQJlCx
X0NolgEmG/1fRt1hOFvJK0LjJOCO5puaU+hymolkF6t7gVV9hie7ja0L8o5efTBJ
lRbIqaj6FO9OKr3y5VmTvAglL1Wjgbaj1oZd2kPbf6E=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 13344)
VZlF+eG08yk7A9PiB4T1vliIwUoqBPsQU6swAIQloAH1+t4Ai5RTHutBSpQL0txT
UXdIwTIzwdpcR7BM+hdTiPyrw0q+48E2maCsymn06Ee/ZelYG93X1kCZ6FhoOlLa
vCQLy1sdwrxMAbSMkAiJZ8Psg4BOk/kQCksgQsHIg4f8oWAd5Dtn2HkEL8I+Hjey
Uag/PCznLFU9yWY67Etvk9aLMUHXbqWHSBrlJmkS5DaRunojWmuEy2h4Hn0x2kZ3
YoUHoL62W0L2KSU0DrJeOB93XDGuJs/uleCv25aZvFY222CNcT5jf+Kc7VU5ELn8
eqc6++Rcvz4eojaQW/A1MkEGOQ/mt75Pw7ozp4PRlHXBNDtyu/xNRWsTaW28Z/zs
idubBS1QSPc/eKP/DB6IEeoclDo83Nn6nq1QW/HI1Bx8+KMvmymplkDA21Bs0PWh
YWpV46TV4lv+v5lGZR8n8Ci8AkdelqGfzShgHfVE3nfn7in8JXUbC4NvDOfHsmL3
T3KQH6AmLWP9qMjOS5+I/Uax1M7uWfkYem7EQ9t3LtbsaH5nGgS3+nkwe1VYxdLS
Cd9PMAi5fYYuaVuMklWcGwy1miHRL2SGHkpwTmoTy9B/X8B9675a26/7jlGonzlJ
EiTIk3/FhvaO/m35B1fdRzsX/SAwb0V06DyqOscMgbkwgyYmu5vPgOxsH9dJGyk6
o7IeHFoDWfVfXhNx+LQCZ2Up17mNVj0Bnle6Q/sOijKYNbmjVCAZv5QYz0rZa05F
HTMG0rhLPn3AkJFOYfmmhSQ0Z3B2fzrcZ4heAlUIh38i62IE7HSM0nprzIRbJFtM
Acgcp4oHth/D0LTLjFiRyOyiLmOqrTrDhJ0yUFfCurikzA3kwyGT6mpe8cY9m4LV
usas3kZ0HA5hEev39RWP5vgUN8LdXKevlwrQgyIn9IUyJA+6GXVmYtuN22nmEMGT
rWOyd+uu295EpPtG91uhJOZJ90RxeDSKk7zQZkPMFoPEfqVdfKb5m+jjhTBqZIrK
wNi9jNzZLaTsKiW56/CuBKhdi48FnR6N+VePcRMLOCK88HWcJEOgL6VZq3fpEY4b
lp+Nx1O1rln70dws5yqOfJUzBMfQJ8sa8seVGuam+bAI/6D9R1PK3/2rGVrkmzBX
SqHQQNKD5a3sP5wc6uR0OnxBa1swT2S+/PdlJzUCE1ohYRGFYL8DifkXJUPEtk0L
PumB9bTZID9QFb9f/NDBtMMxnTjP0DeSlOyTfMWnnuyvxyHxy9zSNVGhO2zZj9hS
dV6+qHsiEm8FgRr1k0Icxi704G13rjuaKIQiFVpUK3MzNROhTkAJtMrcQ3MAQ/po
c1C/zVI78FzRUqZnsncBcoZXc8gPPuWOeWXcxtnZz0WB674LXSgi9VxD2jnzL6yq
yc8ck5lHEdU9KikB6PRPkNu6x80bJtfvmcWR2rUyhAAyOAYa4oMUojP+gnTDDdGS
ruxz4zCoItI3pXhXNVezY33e3j+QqJzQXKwtOCWX9YzDBfRq7UK22hWBIGWO4tVK
RqgNcjc/Pg8Xy38BINnhWhcX6Ae4R8e1dyrrsbTjS1EEfQp52ZL6LnVHUHAudTLP
lQM8Taihdaa71YR8vIDFuNmCe0w7c+P8VBPG11MQ+rN1m6Oq8g+y5e9wycFjpDho
qfEzD00rsswle3Eqzy5bM8v/If7bJhcgy2A1A65W/nEkfQn8srJAYOQCoRxuTN5V
NFh+0k5484vKmht1gPvSrJdLCGj/ZDiQGOhClyRy+I17ug5n1poSFo6aQp2x0m0z
k6FTUFuNIUhML9YTpUBPSD5Vfhjt9yqtztt+hr0MpKU7I49FvsQBHrxMdNoLrlNo
UQUqJ6tp6JgqQdcq0v3xEapxqNBqdeNkVXn9nDiJGqQUuynQsk99PMM8Jg5tQHUT
F5b7fzSkciLZ0CEhXbW9JGWVxBLIhPXcLbCevgnH7pMfK0xVHYfvpq/xk+vLUorJ
Q/0tC5+Ir4QoJLYMLDPhYZqu98uQ+aV+gL3Weqd6uwGjrf9/Vj7dLCmqZEcGATfk
q4J1PgZXWWN+B1m7FVhKOae/LSRuxdT5B6S1WQ/RyUb/ewNItyf/c4FcrEpREcrs
rLC2bpR+8W53e/Jp+6TDo+cg6VL6oilKyzTd2+jgmG4MG0i+RdWVMlMzt6OLIb5Y
ZggDzbq/WkBWIGQaS1VamP6BPL6q/rh/+wSVxqAFz8ABIrRYikoBUvrN4W8sPnrh
aTt6Z4Th6EfW5smz+181AsrhZuYpweohObVDZXd/D4TW7MPDC/eV9HQ7wDwggdVQ
pBVJDDRcI6moUfFVjDX9G+W/8mw+R7vOVCRPsqHmkUX3eZ0ddyVyamtSf4FC7/Wc
z8z7jYTuPOyD/F+P/xeUMVxxrU6WyQEpdxRsA7xYhQnVOAJ3AYWmr0T5HEhFofr3
jRJvd+mR+XA+uStBETq0Yw6kRRMmOUbtOVtuRui2p3vKOrruaU8ur2PScyiyKs5d
+JcE2g+VtCNGhgwAPVcnp9O4GNlWNed7lPFQj7KE+Igo+jcPG3S7hGwSYBYNMGiU
IqvcqEXm18ESquKR5IckiUDPWD21vS6rnqDdNa+fwBFThFq0Vw7Q+3pGkKSY6Wvq
SK0COC+7psiVIgLooC6BuUgCywovbiCnHgcrH1NNyfFgZ2GnxcV7p7BSsXzsuaj/
gYLoBeeVyccs5TD5bHcotRUAv7qNStHI75E2WQfowbrZbGhcPbvJkUI5ird1tOm+
6apHs7np8KkArYO4y9xGq949suBV09Bhmo9icm4erGYgBuwFs3RwTI0uRt9VB6k5
d2r0Tbxw+b0yPlm6d+GhHynwlfx+03eSgo9Iq2IJNEJaCaACTti9AuAvfbvJxVff
Nyr0pv/0ihgKwqqweMMqBlAYn1vsMCxMMFnMNRFk2o9rR45v44IFMbhpAiwn3TiA
CeV901vozrs5SnPB/Nvjfw04jcYLjf5OjW07p8gNktjvAOdOBZSOmnuhVGc2T3DS
K1/oYrmPVibHhx0wZWaiLWS2dt8DWlJDPGuUF5rZl0VGD9lKHFfuXA6og+b1otny
wAYUlHOEBjYwui+ojLgyxQVWEzVcmyB0gJk0CtEGVsosgup2ytkAAhWIBbHlGFZh
XOUxhqBjoi8CnsbG52B9vqs/+Yr9JO61gk68weGLJZeyzswP0P/JBhckFszEwONL
Om0xISHBXt/P7H7OK0ScG929WRspbkRsVk7YHSQIdvbk/ItuFbf0ox466ljpILwi
Z0xlRz/ZVIKojjt/+hjVXP2oO5H+sb/ySDpQ3M4bKpC/pFtFhkaJsTQhGgR/SShO
2do3cPpg56cg6LEg2VnkY6p9lB6Bru8n9ffs7EYLoJToPS02OkkpC5icR029RBG2
WL1WUE0nwS9imwRqKToESr1sMSKCq2KoeijcSyGnInq1Wq/8YGOBIUpgA/mY/Qxk
l9oZOD0cKVqSyHOcIVpsK2E1aTLldMGZl0itR5kARKSfUmYCLI7Jg0yYdPs1dOdE
KTT8LkgaXXcgc1zrP8ie5A6ISroob5ek5Ixq2xg1PH5o3jlMH7j35WGg44kOiJ5B
pNpDYY4HqGboJmSkh+J9WpvYWIQgYKE9yEDCx/ZS/M9dsP0Sg4O/eCbIbpsrV7yH
eqIeXkjCQ+CfpQyxvw6JoRx3KVcpz0/6LRPy6aPYfqs+khX0iRPD2DJ5mHdwATMr
J02/T8JV57vQoUnb1w1ViGDbdEOFoCmenDiwVMVW4lbYPH85CaFCsuFvgVhYCrJX
iN9fAkTNopui9JH3v2pGjSqQO2zU9QnPD+3JHfUjz6w9/lE0yYP6idRhh+3SCq45
SfAo0z7xQqfs6oUpTatqISDqdXMIxgwnJuyixMe5QdJK5bz4GDTKDzimPeIN0d4h
EXzD9PwpNBzgT2wYDLVVJTNHlRIF8iZRQz6Ms0oWm/44INwry6q2f8i8h9uYVe6K
b4Zda9UvJaElnb1EcyT7MW1rTa8LWdcMBEpEcnH/eN8bCb+tbY64ZCzDsyu9l94C
dS9YG7bMpAjJTc3qWceFG6pTSpczEazPmKXRe7YXMScw8yUw8U3tn/9vAy6gU0v0
dx+WhLReoXitWjyWD9ncWyA9rqas8sWoE1D9rykjZv37Uondxd7gNxu9PgO7fkwt
EEzzGLoHZmnhcZ4a6hi2N8xrqXiYgA7Y/lgLg/B1gUkG7IAQu1T7e0oByLtqh5PE
mG4U0r4qmO2xo8MyPyrGOZy9pgVBDMAKpHcdsQ+5GXNjcI014n2UZk+9UoX6K1fb
CbuUs6AV1sbzj0ekHvtYR8NqFtIhq4yKqO9EIbwilfruH5D1EBPxztVcvbtcwfrn
H8wjX8NstJQ9v9Zd+bxuV1LHOKXI0H1q2kME354zo5Uz8KsBIAoj4DcXE38dS3K7
barWsDXV1wqZfTkii0dO2YCL5Xje4Gdg3l2BeIumqMA5htQijjKeQA9HT0eATzeM
KfLES8VftVMd4jg60HngHRGq1J7Cuk4xsIcP1D1da99iRJKLa9+uhAC7XmS1EVIM
go+9hZ/PGreFax05cX8QmhI5NAqL6FnMh8D5H0ynB6cFfjDV2O/pqIOu+Xo26vIv
DccO8UriEYvpLjy1DAVN6GHIxzsecVRUBEUteya6P3icnHqVoDr663Qr55uA/lnM
rLb5Tp8OkFSeFq81wQJdqHYCgS6JyqCQtXlxiIovGh/ZX2pzvS0zM2ml0oO68nAZ
i2/m4962XKsBLhuFqH79eHntecU9ZgVUZ4WtXjuabdHggIeWkpkHzVJYMfqpzu+Q
5O484JJO/RZLHeeUx/maTkmrZo+Yf8jBHpX6voy6f5Y8WbKMJ14aZW+JDugLvHhq
prh0Fg6IAxAp02XRtZAwRdrQZQHW+UZET9i4OrniAQg7dgy+DhSZ5ljJh9yhwF5e
Mhfo5MYXVlR1YvMGTdqpH4YA7nt5dWpMRqILyoXeWjrXkl2//shypGkHa5luYP4x
F950yGyOotuUNZTey7XpTD3OfOX/0IfYPvqDbtA13JGjXdpDVvSIOicMQNl7pdOO
uNe4zgJEF/r8LXcDwLE3iCSPnWDN3BOPmRJ+JBOyb63uAtgF+lzkDPVE2JIRvNRC
5ua/fgrE2YeAQ5QZjAOHkwCN/1py6v9e5getOqMh4/vJUaXAVNZwYiq2vTmq6K2H
XLmCZRQ5tS8QJA5Nas6g2xIcd+ujSpVbLwP18lTfB6iWmpypBCc3aKJ9njfwlOOe
YFAeO4amnwHjv3h2uRX9okT7qufd43yS9lWuqAS+koIt4wfsk5w6967ewGx2dViD
QaZDpryPxKgGv18fvfDfE6MJMtFa6kd5LMYWeR3LOnpW9SieIe8PiZPb1WvlM+/D
lBbVtr71sz1JjbrWBgyoCG+X3zgIJDviI4zTxoy1BDyA4M/BO83Y2g0pwUiG6KZV
aQvtfHHLr0ozirJfBX2RzlwGqFfk6lofFgBacjlwlR1bBGL3dSWwyQipHCEAFhx8
YMpIqhReJ349Q66aGM4PC1JxeeMtSPNoHmOKPEDswoMgJRf9Rlpu7ntrD2WcjVqw
AQe9pcOZV7NVufUwbyHv/MQh73r2bSWMFypfQJ8lz8Wj87rXTAjqyfS6gngk8CgN
RoIuSSapUI2PkS1RjBLVKP39zW2+yrC4NjJA4s5YL5M+nr8Q9+Dp4pUCTG7OfrqJ
/MYqRr7r+zvQipof1t6R3VfNIWatgKgjiVFvghzNVRHUsILIM3u7s5OE+2mFgxg4
OBWXa2edp6sS3BY3ywh73+dLXTlVrUR6fEgZxZmiLaQxrpzd4T+AlMFBeP51aABU
i5N81vGG/DTPDdUGxOwofACIBpZyq69VzNxkvSJ/rV2IkxEEj7jkD+0huwDvyZWf
EnU43VH4hyklUaVcJohRbGWCvSeS8Zx3c1cIdt8B9mLOdZwZ0gaB9t/dtZuqf8Xb
bSbNxmJ6Lemj4y7OlxtorhegbQxULFPhbFbG/dAd7zN59dIzSZhg8G6P156P47x6
hyr6SvcloOArfoFVBPQj5PeUNMqywVFzQWqpMcQNpTKcxYku1iLOLVSSwwH5RPNC
rhlT3V5vRGr51BNIbGtYwaoEtmg4bLhpor2hU0Z4YG2IjMZCa30xpgkDXZ1OinKG
ReoQ2mVrz5P+Hkb/2Hny139kvLfZllhPc7FjIqSWX1VYlVEmO47VthH6WYYfrAsN
5VFwJMVbYQHznWPt1ZIv3gmyS/Uepjkff6+k2hCcjf9G+oUg22Iz9VcP29w5uTvA
JtFDrYgOfsoHPY0yrSqNTgDARDz6TcaZMdZlRbP9sWmVRFeegaHUOZmr1eyZTEd8
+Wk1d6cVBi93sxiqUpMxeuVBpH2it8dt4RMPl+pC4rxqFK2ttDXupeh0Y19zv4bI
o1/xp4imjmncRnMAO6d4/0lvtVodYP3Up/w3hXJWMjzhqXlYmMbIIv7q+geI1Mzq
mXvhnhYRY9ZS5LlJspnYt1MzJnpaq/zkE2evr/sg3PO4m3DTrSEVpmV+NROFdrO5
avGkTBPapepW6f+pYpyBP6bDXJoG80Ty1sD7TMUY2fgVtukQ99VpFGq8S3CQ8tEg
p7mDS1tuitG+EyIgWewxnPi9RzmqHkYdx97Aic/VEnYWjVFk26tOTihx52R5aTHw
VWSMexzN+qtRSm7ZuDN09+kq8X7wuwLCyCGQve69676XNGauic6/hyyt924E2wFD
Sq6BcX5aukMqj6zZCAcjmD7RieMhTBfskkEoDy0UPpFf9bgDr9ua07oVaBjRRmVe
XfMEShBm+ahGX09zcMkheDFsVSVrKXAENwAsLO3maOHoetrUfaN/00wxqycHmBLM
vlWKb1mxKWWgEKLAJW5dsKwTSHONTJFUPt+VXDWJI9X3d1yUDxqzdERGuwySBU83
4NEl2oOQJmbMTeeFzI2VAfuqKdaxBiqN+sqEBT0LPrCervuOqE2YzmhWyExBUHMN
OrtIccIEP/uUTr88bBJF0/arJ1PLemE0/qhwVq9AZDnUVltNdmKJN+m/CUK3jVO5
CHfqbyAQXKWenOnvLpUPNBubCWkYcaJ4c/Vx718L7C07bQuHcZcdI3fh69X78LcU
XCUfX9JO9wMHmndQRjTxMghCIs68hoR2darSZl0p/dp3tvU+11KVGwC0QoAuUt8N
yDB73Md3YBpLeT3ouhDy9WeMuMPhy7HP6Jk7mOyKGTLHhTrUwHxxw85fZg6BpV+v
p6r+4R6U9NLQnQXA35L+ONvUHnzXb3ULgFhTL70sLxJN9nRjK1g21PMp/cWehlcl
qpKqum/KUlzbPOWej6ottq9SPRZqSmSQ27vSvzn6ecQnZHUaQc8gdNOwLcU8tf5m
1eCRYPQoPGoUmpk3XlvIVgUXO/JrMuEzyNpCRrNj1aididXlwA63o3blGlKedaVp
Ris3MFk2Q+4Oua2Z+Ly5ybVlO4qThXYT2VcNrssTQgotlTfx2nzj9qGKkbsFpabr
e2dKheFtMk0rFNT9xoOuVrGI7sOSc4vGlX4zVPSRCEAOYrirCzy65UDdz830Diso
YcCHAV7r5LQYj6aEVqEClCs4LctPPJvIJE6fmD8CVQOq1gq2jCwXo9aTmJe2Yl3/
HZ52pmbREgGnM77BlE9ikdeka4l084nhKnryz4N/oRPo8s7DA7SuM0j+L0dK+m++
5zDoV/1jL0FiDUI/8+fPAyioHvEkDHaKsPlZ2njHE8xLjS8JloNP/1P41wPi/+Rj
oOS+1zqm3D7J2TsR4DAOcB1Eegpa49RNSOpaapMP7ApCLV9e3fmgyYdsZzDKTX2M
cyniiQulHwaoKOn+9bIS7V9Wkm+J/EQkrAyBgLZboAZagUR0JJVVc70QdBOoBCuM
u3GnHY2xZHiePJDZ6yuQVuWdw6Ev1Si0eSWhYD0yh89ZrvL877by8v3mtHb79tCC
Mjsi03VpLacW+Fm3DmFG/nkblfvrW/lVzwBrVZEMmXbIL6MBvdbCzVsYwKZ+5gRX
AnWy5z6siGeKoE1Seyvf8p0oZ9oii3SYGBOl2dQbvHWVR+g44TWi/sEsEON5qeNW
MxyUY5CmdwqgJGnFnRzkcnd3iJ6KbBWYin3CvRo1ywnkiz6LZBWKuf3U0CJSojQc
XiOP0uMjVl7/+/+oHyjr7o99v7NqHLfjIcxa/aUzq1tdH2ixDLsaavC8xWo+yLY3
eJkqLiORr7P+oyobEOmBlwA/N7XWFe3Yn3HthTLaWxagz97uafjoREuGBwwwDFlQ
UU0Wna6HBPHuDQ57j6tgLdR9le8wlj3Nulhj7x8AGrAW9V46GvkOAVTJ/nvgpGqe
jZC5ET+9Y7Lqt1KAZs7XaxIGmFv9OJ1m9T+Ch5iWVeRkeReHnwxr/XhbC5Ai5AXD
QLO+QDokFkabw9XkPcHzU1kjDUFWA7Qtbmwy6gnXfa0eVjOmJIr4cOsTH3aD8hqy
ooqSem1zUnBC3oMQjfIa0hJVIyWIK+AzfM/ErmEh3DBgdCWF6b5XnKvRN5D0qHKS
fQSNrzRjeId2RBZq3LurOhe0z6/u/fzNlLPz2O+k9orna1J6AWVTy8HqMf4nHVcB
kPrBd5QN/80wdL3B+uhQRe8caEOCKcMRtdYSPujAJZ3w2ajk/QpL0iTFB9mVO21o
iCEuocr71dGPhPF8DcZWBVBi+GrcYlsSS5R9KyElIUew2gm+IXyJqIWj/f+cbAJ/
OevY9zY2146lbssMH1pPLOynkZcXNv2LmM1jhPDoD0VHpc7nAZnSeGw/zV6SPQXr
KX2Odr7kHdGbNt4vV9Cby4R/LQj1TCbxl9uXygLVVnQLPNNINc6glg1uVTZ6jWKz
x3NbOhO2YSo7q/rb+raA0QxWUx29CvVW7oS18D/d6YmuWNCUAhQH13o/RfoMDiYL
3QMWDQ6MCpM22t6y34Xwi9BiGBFowr453kJM5lXNW8tWMO8iAP0yX+8kGqrRwvbG
IELm6nozcS7pcQ6F89DFBOer/DeaF4P2isxjAyOmGw6p+SgSdpoGdF7lQIjddPjy
jxJXJOAul8wG7g9jrgpLou80WS4929yYOUxiwpTnsRWpdF2tcQHQv9vwXj8PftjT
YcPh9/U51/X+11GrF4a7cHhrxNiXIMR8ZWymjxYk5LNkx4NrBlFKV7laedL123pv
mUh8sQUhHzbdG7sXlRTk9Oi2LBIn/9BWagEYNwZQI+SZKeUyfYSXpt9nxH+dRsFG
hGHJGjvhAINGkH8hgtoBcKeVynl/T2R4YyEoCxMLrvy28DIlGjkQdRxHHfXWYTXD
yrgB7lefzqVmWIxy3AXHsibiH6xCBsP6nhJIITidPmV118hSc/9RinG2Qgna4L4r
UNKwYtO/UX2EmJjrG2OA0MDRR+HcESJdS/fRIpQcw3F2WanV7+wZz/DJMgsWlCw+
yDRlGHpi9qGGu0WUhbONFDDeigy+zr7YZIvznsKiw6Fk+Z7TwtmC+8gW8oK7XXJG
0UX5BaKqwGgcPW/+mzPwCdbYpoJybtl4y5MEiqzbys5x5bm4M0//T9OBeF1ZSMcU
gCry8j/byYmyDVeW2ClviN/1jU+hdEL94K0tZuQSgwCO9G9ErxjLcBAxWDnd7CW9
wuEiM/D0liUOVB+VgR7bjHwIDszyrvE5AGbC4nNuG/sKuFgwe2+l/61SuZtE+nSO
HeQ2g0hWfxRnqnKeVQJEnM7/3S0oU08TLx/DjLjuqg2qHnoblLqbH773IXauepTp
dfhgwJXtA6Ep7WbTUywU4KVSUhQPh5NcShYEQj27G4tz/wp66OBEQxF9UQn9TqgX
JBNQrKXSQn3rm4EQCX46dV2zmf0/0zHZu05tkD082OQmjr2suR2SxOCbMbFhAkvR
5FZe+pTxeg2ZlSDhzjHaVaPYoCfitdlCbGPxcWdaXw7ZZicT2p/N4h4exn0/3YvP
j9uLmp20HRmDD5U0Ct02vQ150drhrhGxU3YLMFchDK4E4yYsRbtXVAj/GZCa6pZl
KSfihZ9rjyd8CgxvILfGmsCdrsCLjmCdZ4TQh6p95q688kFDzoAVTv1xBDQUh50g
2Nwm+fvQRx6ZcDWLXQ8LDF0JkcLKsxsjwHJ+oK+ShNe/8pO/XRAdHa/doYruJXjP
7bBbNo/lnZYItB0ho3I8vpXdsBeM3DIm+5CJuWAer0GK9Bp6X4PBX5DA+YzMp9P4
z2rSR7dOV5pY9KRCxPi7HwK5/EWHROi91Zg9d73+VFfWNNHge/a+Ia7kLrqhY9wg
Du9QO1OiRwcuDwWByNJd10QA2XXNSS1UajxnzgPD4fDvZ7MmCguMhKKaY0vUSOC9
nTz98FaO2e1tHjez6RUxwZ5k8IvlzF9iWpRtqinP4duJfDbMC2zKcb6LtwtabJ1M
U4d02khWqvl94o3i7IU3ZVWU2GJPqkIg9mJ/0la/K6GyxzIg6F8ga5jyCxoeXoTI
iok8EFhZ3jaX/81iUQ5RedTUslYP30hfDVFUef/tJUMdCFEZKIjfAOSQUNQ1KuG0
phVMuIYLb0r0rnAO3/aWMgMFYv3W8XX5uTP5RNJW1i3QIA61nPyQ/ybyCbiBARKS
vO2+DIIg2xdHyxwuopMJCcXfZWHnn55JNVK8NBTVL82UYT6k36pcgBh7XziMsUtW
ektBDNrAoq/6k9g/D1EVwj+6JggCIXe7dClpG7SC42A94i1mb/70CvmGxAFK+iBK
S2HDYJqq7/aFQmlbCwse7kjICnMjMhDFK2tHv7nsiC0DY5qkswjw4xn+HO4/R65X
3rkUKTbneZvbcbWowsgB/UIBVfajJLy2VeOrWPtMh5NFCq76kIjp6lG8fgCPfJ/d
8n2kmuIl3IK1LvO9kpsRQ+us6khezVzF9+wx8vbMCAL8t9n2PefI4vrqoYeFosen
lI/228WRmyO0WLVKOlPk3z2C0NGb11aqhlO5fJKk1qU10ior9Mm2P/FtgkCnqrab
E8xkAgu/r03p3gnd/u0l5TABmAl9GKN7gGY7r7RVx9rt6qKt8XeL1JY1FFIwBiG2
XulKZuYhC/bkg+XTwPqa5AfAVty37Vg0auJiFOQhtX8pd8Uahf/AgK+RMNo0bX02
IBixBI4uJLCycDHIJzcTW5famP1MJPsYr3Dk/QEC/vl5NuipwVaknoFpFV0KXRIq
POpxoEC2uaekdroMBcqVBhpX/NGl6cvPsQOeeSxikzi7JBL26IMazuRBoiySwKJT
AUpwHmafuuyi9ZEOkKsX+UdLsYktqpJ1nZMGLwX8KwUYQEKSErMvAtlRIFSG2Etw
ka1Df2Mw8LWwKsYIHqslW1Ewrsux7xc/eZoTvQgdBFarEQQVbgkENMm3K11CMxby
2y+KxjN8JL8kIkLgO24eOTWoCUA4eLWNea7peBENHSBNS313LNPDAlmqayRaQdm7
fs0yxUmNF+JBXGODA32E0Y7E5pBRIyDf6TZamPhuksFzyeiAaYZgBjsMkn5jtR6a
885kvieCP663NtyTKoVI7VtLAFXOwYqoJIUBq/NN073QjP/kgEdPkbgjloOZduzI
p9WG7fAixVp9g7/uZc/cUSGK+pgNoigRtxdt/rCDQ0c+cmqSMIwC+uBdNEGH4k5C
MASn1M/+wfbMyz6BCLKsor/g8ERXH0ePB9MR4Urk+TOMrb3zhRFk7rY15x++2YEK
5KZO7Sn639uN228RN3UzJuC/ibEC4f+w7Tn4sWOMrFzmAtJKn+EktGeRIcZWkthh
Q5m1pnlUtqyMNpnESCUCvi/me3eUoCU6itQSQqpE2V7g08QI258DbVv0lbUfwxEH
ED1TSa68jp7ir+lHMaHf0YkjEEZJiVnLLgREoQS02JFl+XwHLys6jKm+6NcXFazM
nriyG1DK/lCNh27jUvPQeUxZ2xQ9QTsNp15iswrDNqxWCQgf70j+bzJG/1G6J9o2
YmWSaXZDJQxWSpYUJMcmo2P/OXDJCJAWoDdIm1cVXOgyOkeD0SYjmJ2wH3efdAuN
MoBgf5HWhqldFR0ljbuqDSPpyiOnAgTKaFRT+63QZw4d0GsRy03az+1E9cGLP+fw
syIklqpQX/21y25ur/vaCLoIEqpIDtGs+xCziwBiwphiDvStkalgsscnHnOqVYW3
JaEdCvfZSW52BU6bb6KTXCzCZXwhmBldVGt+YlxMWVt4jLEo2x4OHshf6Xpnf7oe
RtPxhwMcBIlUSSrzp9o7+/nVBzHrg7Scz2rFV30zdl/mB5XvrZSTtaCa//k1tR20
pmVWDghG5fvDY8eSlaGzzYfp0Jo1DR1AgbUvf2lEjm/Pi6OzJxoFurevj2inwN+N
iOCCy2sWJBQwFLX+JnAy3mls75ZoRdACtATDXq+ejPhaaqkQC/Tu3XFPh0yQxXXb
1mORFDGdXWavzbtqm4OK157ZNV4/nhsr4AhEF1d06FN8U1fkPaa0j8+xSkjoD/Tf
9RsAohxMZqcVJaFOfxwPd26vUQqQaExJXzaag4ukwqZ/IErvy120G049RKWQrHHU
59nBCSoRSRq6RouYkubKrNxN0bA0WZ1lByRXeWuHEZB9Vp8Aj672Wc4/0kNDAyTT
dFULha0a05UHaV3AxQJBOiN86IqL7WJ0Nsta2ZUY3She4bqLRUkAsRbJx61pbai9
zYysj9/zNytSx3V3V/smMlSzT8PrcyYDAChlMXqZj+WEXeoFRz3gEbfJqS1K5Ypl
JOPw7eu7IRtPwrA3h+r5ko0r2Rs2bY7dt368thNmNnLMVo35Oq8XNmT28YbG7Dl8
UkSqr6cg/oYPGhUIcOecxr7sb337O+mi3d0iVZRtQsfMujk0muBg459+kh3JZJar
C3XzI4SsET9JPwNB1Y1bSwmoiIQlKK/7bLI/d5C2AhZb+EZuNMwVpRy6CR4sSR4t
JXl4U+Ea2SDY+4D5d8e5EUDrln1ZjU+CEE+p0sJuANA8mRyuLhQpxJmEIxvHdV6s
DT9oLq6N8rkBfbmIZjPBxVraIcMOpSNLVLn1BFhQsaNYtOkkx9r2VVN3jyQ5W5Ad
zScVKnjJxLeAecOjTTuNF3Vk0zrDGoQnfcif5kxIQkENtDB4tXIXmyvFg65z96oa
TmB6phqNLjR2U8wHkmXM+eVkW3Cb0CGmeHjtV5X39KlnNy6ESvbAwuOSHPiNSups
jQxuDJG0h3uCJ4FrVmtFnCo02GGw68wyhnYTV7CCzIcOuliRzpmMiAX2RGH+N/ma
wrqn9/6srqLKO1nlMQ5TolZmSah1HJueEFlTAAOhjAmssbVvwwd7v7MCY1fDWBfv
uxtfHqwUMySiTxRglq1MTdoVkjOMbxptixMrZ40qrPRpfVANezPDR1AKCC8UbBZv
gjmLiNQmqQ//Oe4a9i+se0uERIqi0IbfBf296hVDEkfgs8GbcEzrbDnHtfl/nCy3
KuUQMLebhMxtICm85nTkq/3faSFsfPeRsrP4eB/TWr8mSq9F4MzXCQ6jZ6mPbZ0m
Q+wbE9tVvoAdHISAhO9HUrzReB9gJ0WHv25jxuMHm69Vn7afW8D4f5XKx33zeEr7
LqZB6OFippTI3OwRORq5rZLAdW9CBe6vgYa7q9ghEmoERhAft/OTqIgfBmakNn50
wCe55lJP6cZSvgjAbuoGeiVty7if7XcZgMSn99gO3qpOg4HMGz56oIoC2hvTfqH3
G6uOonB8V07PiySe4P4vSzetqS0yf2hFvtwyjq0Ih/Z9Is29KLcd8tl8invLFt/w
aRFWOjEbsyvTBrGZIYY4z2pSw1/42KRXP9uKuR3d5JIh0hp37STuyebAK6ZAOhpw
9bwR6gVVC30dVSAd5oBTWmUAET7EKg5Z+2+fUC7Vsi2RXZBDhU2MEEed/fzSOxn5
YTTtriscMK0o3TvYf6WKOWceu1cIzqt8BRCwPrGEpFkiC/4bctgp8nP765jSbdlR
PwbTQlS+5Ex0j9I6ePbAL8tTJtnRiLfuq/Ys9sjhHHshR2SGLBVmmsGk+NWv6uhu
1zdgPWh3giHDyRn3X5Pw1j/yTRuMwAh6cEhHJGnwMmjmC+3q6oosTuMxzK1KSHQd
jwffYlFZZup0jowADmcxbTzcGKs7eEXGJ2WAH2MKt8q/nlC9SOFI6ANpMz4cldD0
BHeLg8vCBpfCByQBzdcMxWbGmTX3BHMyWwq/ewiVk+zj+2NRPZPjyyqYE2vdxwfL
WZh9Cx5otnEUNxXTDg4JLxI+5ESMUaFmNaD/bkJ2+UWtJ5gQQppmCR5jZCnq2FS3
anc5ofa5d/2z/Or2GnHUf22G5RVsl8d9TdftDbtoE/mv76zQYyVjfUXkrX9/Wr+f
D8cScIRdsjnSoeWCWYnbl65BqCmJt2WPQvBKG9mpb2uIMWD+bTtrpusGgi127ACB
J0fNhLXF1M2118Ij+khe7s7ah3bo/JoCOETalwxciKO5Ruiw9f+mcqId/rnmLo5y
uOLQKkhXNJpRs24DjZyYw1zar9lSKieW1o26N2wkqtKYu4gDGn99VlifeaIvZ5W/
XEmuPj+Qkj8Vc0RQTXz6y6CHqtl/pgnYOGzXq5Hr89hLtzLHZJ+J9x2fpphulQSK
pH6PT/eLDmHVEcB3EzhVkXbM9SowzRZ8Dcw+/6aOXLqm3Eta92C/Fnr/mitdYZAb
aH1gfY/Jhj1lQ5j88yCh3107Xk6FUHpo55vYuG6Xmz27KsEVw8jHHlk4eQB1VkEF
PzS3+/q4d4AvGiksx7lWMlAHdjEjTPN9sx45sOIF27u25VlN/PXVOW+X9Uet0p2N
HJNTM4VDeyGpFOatrcc0JKdo0VBciLKeEneM0LKvZIQG1X17o2Ot4FVdWc4NWyKw
OiiYZmC01bKtimuNSmHWP1vj5oh5QqBcAxR5f+P836P2QILckwRIzs3riIZScwVN
VcFeX8XT8U02NZ0QqaILulDvNZ4oItupKpoRklp3UHhBw/PkwlDugPXf7qOCZmGb
R4Or4ZhafrjuQxoSSwrRkFfvY2obKJ3L7LHT43XoMIoWlnoMYm5FrkgcDHGoLJUO
0Daan0MxPtZhDm3Chy4NTNRt+J+Z7PyYdO+4w4vosGJG7i1UU+ZYLm2jSVPugnpp
a0X15Bikfx7OJ8j0k6p5TmI55x1D2nq2AyMEe0JYotEBPzz1duaNYCFGhYf1kBJG
7+H6wVrZkOXMvxC74RbTT0iU2o6/Oq6sxpbJUpBttCFtZE29uuf2dxP3bhRnSY6y
XyYgzHEwxIN/tE4thlcFB6I+1ShBkMpLIagCe9T7/jmm62Guozh+nL1b8BM6o7KL
8+4JpE6aMeigCvyTBhxUlcyfkP1t4/m1OaIsc1rZAV2ANBlIxh4MChRycVBgms/Q
MGOxoSoTgihSzqKFd1KIcYPCA3/iKF2jhHpftCN/mAG8IrShs4LJ2xZD083rGkcu
HVZzZjDzQBNdXBebh1OmpAME6FkPUm1iRCvIGtuyvqPGiapvRkZ2X9LDDtWbY6Z2
HXX40PsnjsnrcogEsIBk/2pa8urd49KObvXMWwWJIE/MC9tNNb5oc19tt8yE+3WJ
LwAdfTkEkWk1QN5/oCk57c+VB2EKj12qhDBuiGReqP5iNXvhzcBGa51TCxiWfxIp
yDOCpoN1ysMJAkiLZTGpO7GaGA3zj/gdXE+VaaJqRDHcuEWjQhEfrITclMmqrbkK
OP0KXz9EKPCBVRW2qIHBytN7F/hOCW376dRIEnjuZ1iU7ZFgpDoQt8gRRe048mLJ
cUDdZuioqBuWKopePH5Fp3Xl9bQ81gZjiUyU01AfyxBwftUB344KFs4NX4vPAAZi
RnC3PqKZH66/lK7SOT0yLSZ5LbquGd2Kp2KW1XXE4vCzlhchhENOL9z3JQfMbpm8
sGujpjsChA982RGG3XOVU2uJBI9OS0KwDU/zUm8pKJo/4zJDzr4sRtu8BJhM3vlt
o6FJ8/hwI/XVWcZH8OK/hPb7rK4nT8yu4u5EqdJbQUZFtULOhSo6kOjMvLA0Jrhy
g8uCDzXw3fGwtQ08BIqBV6LuP6WliB+chvde5Zsp+fKNo0soN3+x1xsEhmL5Mjv/
2rWuTGjQ2qoT4O9GKuXl67PEaxla4P9SPzTNe95V0NPpInD6tJgt1H22DqPlsguJ
i5BAIpBHRzd+Z9GwNdl+IgTF4bwy1Z9B9DtsQsacsR8Goc0gqi/UgIDi/+DpMW6M
6n6rQVn1XlGK+9UTkl/RedTHvRDkN0YmxZqaMTioQjQvxZ0UhVGInVmRlKnZpV4O
fe0XjXztwtvgYnEaJwqB4C5DSN340yGutzA2hUUwoCTK8W9/GZabO6UdcFNeu4/7
seIcjGc4ufv1GC9cksoSt0I1Cl/2qgbsh+naQVCisn4OGpDevokjiQxZPLOEmVHY
upMDhuTxoqcWNy7dHThzuEVC2vtKeXnlupPTDO0A+312/rIBjnS3eXnu2EpzcJRo
YDUwoJvDBqZa6DNONVUFugo8g2XVgyChkEBq3ChyxSVuxUQoGpg79O3kBgWOBh8I
dh7pdwdI35Pr3Y6y4BhFv6pZ7BvIoaOcXH99UcnmRYuzV540foiQVOLxRi7HVz1/
358wQQOhdmvX5vfpkvnWDajkzxUUMXgeBUpnpvBgO4fdf+CFHzrRq4XTkMweYaEz
0Vccn7Fh5b8Lo3/dwWJnetEm0QOcYU7rROpy55gg46wLPvpoQ2Vy4LWwrm4Bj8VK
zsrH0oSNg/ZgzGQk5pyxtNJZp9VNHOCvt2CbSytjM1vh3ARXfM+DGLQ4Y1wVukOM
CDNJF0aC4K38CPMhZqO3Q8lHtSNmR/Z0TWAXcgkLla0l5IR35+RX1TrdT8spFIzu
XWvmrGIj/mooD/TZpDj9JKNlo3XlcSu8INkmwte33Hq/2xkNdRMc9Qwxyp45pkS/
K5U+v496PhWREbGYrUeJ8cwiCq4wxwy/EdHIvH4gMl8hMZWYLkUm6BOgC3HUgE8e
VO8opp1jsPqtzhV9t+zqJw2SKGwJ50AiUlf6LD7TZAY8Xv3hxRnicZDsHOTJr6Q8
bGntVfvqpCUHnSrgVXMPkbqN3Y3SNOacm3UZZGmIaEq/+wG3C+C+OhaunZ9j3l+9
TEoiNAuYlmWOkHJJy7pCU3+PkDfwdzTgPhlq+D4mfR25jcMPZHYr0XEcop7zTSGk
EE5XqZzUDl1fEVHPnO7IrAr60AJ/SsQsDmkjVAja4PddYZIgZ3FiYlsLnNG3tM3m
QEctaBNmhflRSSPko83N8I35GrMZh31vaZ/x8ltjSXgJclrtlTPmmNZMopNfpGxB
oXSG+MWudi3qJjC5wHD2dl2R0tfrpiT89YdyQLkLAjJEhAE4ACG1ZJkVMTRd/tWc
ux/kbkLA4aZlb8Is44Qtqm1dWL22Nrtj94nOXXMHfLYl8KVhq6kcl9Xwc8J+a2j9
XRrcYuvCiD2nK5MLHxe6bYUf6Ebv5rPRdHgncSFdtqj6lTKYnTt84ZYlXH7qwVp7
+JnZRdSWaMZ7ogju1Y890wHp5Y04StpDXQLm1UUYCnwOLM3Q4WGUwV/1qsRAisVr
hH7c6jikDVUQ9MY06r6E5SHLOJFTg4vrznAsMwvpA2AoJxHy11YYKZ7Uegr/ZPl+
0Q0822jVPoWpYhqzogUoCPR61DqIeisasb915Z5+krwgGzgEzABbs/CRxS9IzpZJ
6hwbYaOMx4MrSTpBAmIO8lwPesAPFZ1M43iJqxzaqdun0qTB6ovXwHVdQhwbasoZ
QRm17clc2d5G9CaPh43Sl4vJnIYwDqSeQx+lZulHyuUc8JBVNstPZRj2C6OUr2HU
Ydm/dV1SCVx4WgG7NPWDSXn6qEFM317GFZkKU2ifoT6/nZZpue+Itt9XT4p8wxVO
`pragma protect end_protected
