// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:05:37 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Ld4Tfl1cMOdgw585kkIIji0X52oi5HOIgpU4N3aAnltiTDY2lCvCk5clIi/QYSVP
YA+CoFSE0u+xHyH1YenSD3DNKiqUUP+VMQdHXkdF516ctlQ9ZecRdOfUU8nObsXu
OVp8aMXPhPhYkDd6KsieeWRC+sSLGZsp9KwPZDx/F9A=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11296)
suMo2/Ee9rU6JBG9J1PzOGt70EOeY4ptKg+DFnlmk5GFrPLkTQCpOAc0vRxrRoEM
hvwbeohJeE2X5Nfi7/s19mu+33rrDzT0eV6ZF6v6AY083S+ZBjK413OJCPls3B8v
lPLyV5fP4TedHa5hZBEIbR1xT6H0/SHEMr5q9GfgjMrW/9mij7bsLs+6febbRsIm
F8dFTCai+vytTBoiCKeSukudnbA5FNJFdzab2f6PAHd8OM7ncd70ZkHqV1me6Z9u
Q3P7xU7xJrOBhbniTibKeA7lx5VmkaqLjdMN24MBTYOWlB/UpoIwwPfCaoAH8zql
pP4pWiC27I5xqxacs1ulhPiASLm7y4LA5n0OQtTsOz6w/NkLC6TQQWYJp8feshOa
FkfHm+OEggso7RdYku/4PnSmSEyyfm+uGkokaxwBB4tSomp1Ec97rxZTgfEWHeZb
xepOON7MIWRkyfdt9pl1CRAzADEv8lv6CJ/6A/gWtDk2v7lcGoBpWiyo//TW9u5m
0udwQNDDY7PatZqQDDYs6ZD0MEBpY+jg29ku7OJLyYQpYEGzlDrz9jQV0GRDsVDO
gmtRrEFPC1SBfNyC2wAFRNNo58rl1ghTlKFOzxkeU/7KaZfdyQTGSL7j9vW7IOcG
3LgsXwo6J7nEhNg4deoR4aghoS4x8zTG/NmTQAi4gBLJzWPxQVpO92e7q55r2blJ
MsNAOj89oqeuTMp8zbxl71dLchS3D+W7Y/G/FkSn1oS6n9jdBFTvECw+bSzp3W6f
U5fXA28S2euPLJB/tEkCQjaaPzBefX13EeIdm9sncJ+t7gycgOTz9mQx/vGDAef3
PRSCBoTpqCeVq44p6Bu9pL17rzb+BsuYV3+7zKWW6fdNi4D4CpQibwTrR+LZMum2
RGDRaDZBRrVQgBcNlT3ZiRYWHvLjdzh7eoOOMbMvKinasoXvVjf6CNBamlGsLU/u
DZpEf2u4bes17limIA8iFjxGojfLU7gVX3Wqa0+4yPsT64e6VSXvz9+ViPBk4zxj
hrV6qwSioC1ALBmP7onQGLn2lZIIOB7oKKSp56QJNIVZXqZSJVY2imZMQUlU8bql
E0pFxBTLypzJaHmvRwbW4+5bDCjYiysEh82c2BDnAde/h3FeWd14v5v0/mW3lx0G
BvT2ekRfZvFPfUVMtdJrEs5/PZ2cEMBi3fWHI90xDE6NZgLy8SH9gY964QadS2u9
DwGXEEuOau48Wn61qL0RXymQ86BSD6ev6Gy642m+VoCNoGGerkS0ifxjI1y5NanB
1vXK2pbDwWxANLUzcfnfdUVEA00P/TL+HWChBCfK7EF8u0l+/kwWEKDrtyqhuQtp
ivbJmzvc+4eP+yrgW1LCG4/0YBm2lI9i3zRB0CWbEMhgN1ge4Ya4rrfXv3FvZNwH
PSWqxn5GTod4hblgbx4rNPGKhwxE0vK6qw68lfwXj3luqyeyskrGUofTgqn/xJJL
iLB/WEV0HKHi77/hHPDHFrobMdHAPRQZwe4MzUt3Bgv09Uh7js/IYyOmvs3S5IFG
NTkEoD43OfBaUqB3HlSKVNN7IRGwaJHiAN6JMjyZ+fOWdBAtSs7vaPUU8S6fycsw
hJJtEdGCMQ/QU1no4yQ2AOGrVZAXNAHKoCbhUt1V4q7GC3DkxyDqjWfuHN9Z+pYe
2Y//0nLwHFyamc5htGHapa2vKkHf/5sFBsMjfMoRObG8NLEPU/rIn6hKmIDeO5nX
+IgDGQfcReNDvoL7PUxNQItdmUtdcujaz2m5ZzcdJ63I4g4OUW3HxpNe/DzYhnvB
7Ex9MFF9EjMzSB15qd4j1fgRnJqQdl6mHqQ1MmSGVgt5Mi+/mz+aqe07Pa5EKGX1
OfFni8/3HeCN3YArocYngILrePt8niakLabAn8wkw8aPeRIlbeGBySKytFCpAThs
0xK3pfWwl5HKZZWzjEj+OwVyl1GJRRGytT2nTTzPyO6N2EJFPAPdHufr5LMu8F/W
WSqa2AsLtIw/ziyK9qm4eCVgNH/zunH9180Pkt1gcooDlzSNzeUhccpCPMmvV1Qq
RjTuH/daRiJMd6ekMrAjPlyeYO9gqMOtWnVevgc6Cu9Rh44sIL1chDb7vChadkJi
z24qaE0uL2HCdRuhqGlErqDeQpMzjvjoI87RyfmuAo6nqJd38gWW5or0CoUVGYKg
fzuAkI8uG+mfhKMg/iGL3UCYS/7LQuHTN6LjFLWq+IURXihRxSB0O5U+bPNGBgtQ
UjBxqmW3RhHx9Z83PNL+hL+vMEYHiTtB23T0xiI97NGUYapLTw+fTBWsNt/SS+nh
TkrGynpLd7BEkyetr7WA/ufvWGR0NAc4miINsxJ7sQJmQWV7Kly1lSqAOB25nZj+
V88zkh8JWNNxSNyhbQRX/mlspN2hsPxkN5m6g7DJrE6QmBhqHbf1/xN/LC3eDaCE
mXz0eFk+EreubEqhIEzcqzUDsnbrKCijImlKC8um4d1P+pJxBz9g9auRDysskyiM
IXPQhjhTa5c/qbZv5GGfKDc0rwFUFm30fppM31n3u13bfiGWh1ka9CLJbgl4UGxS
J9Eb45Lw0pa8GwMFQsjKPBlGuU0An6Y30SLiHuKrpIHOQyd/2yUXVUG8y0p1T6l+
EusfFDP/b9m5eyjH9EqRHDznPhjzkl289Arrykrh9b0nvb2GSY/3tSQJdXk9+SzI
GYRz42glt9+2ARnn/ttM34UDMyQ9IGB388cgBr4Pq7Wz/72GVS1oDe/rysudL9EK
6wKRmqwLNOu9iA7FXwFV0i1rGgG+LAQLq2Kk0PZldJO2dm9FBk9W/nQf5DvMkTNJ
NtmtZqVqeyiwrrgPXt4mnVMHAea9ZLw0cQqA6XJY3uLGpbYouFVF2HpkgvVlYm0+
W2hIbKkMFUh2718pDDws0Tx35BSgctU0Dnwull/ArZiJW5l+Pjf1dfGBwiOGi4Ec
n33MkG2Evz/9yZDaVRsjcZepTSbIsTdcvYCLqHf+kUhEh5/59CbumZDjjR/C8NbP
tLQF/afAs07folapfgvQ3ZslNfajqjQ+LocCTRuJ+sOytKSqEsdgo9EeW+hyh8M4
IiXJt7SYc/NlWUMTF7XzlqT2JbTZj/EbjkOPLYuGK5YTQ5n4Hv9WSw9bZ/krEepc
JIyjV8Ui0JW/cxnPS1k07y9XXZ4mA3+KMcSdUWj5de4omcjP4BFYQ5/hbSDfwwFe
hvOQKQVb++JVVCBFY0GRlyQKydwXJfyHwd5G3nMbN5Sn2s7/Sh6iXZ5exiB8fm+C
0uL0M96xyhNt0zGTe6uXjWM+jd6Y7o7oUah7YbMryxCuvk7QduRq0tjkgM733TlQ
+K+pQDDkpOVWAVPAYd0HMiNP9NvuTnHcCA5MZElq0cRXbFxV4IH5eokE9Jxqh9Z4
KmaiAlw75EQue1Z1CGx3WuFEdZPKDFo7tddQjUnSXl94gaBywUgxY24JqMSSz+v8
JMtF/BerN3O2i2T0aKNzdkMk13/fEb1+sAE4Gd6VbWBV3EKP7B/2RP3apwWufS8l
PWjkqqzY05U1Tg49AwqmG0XJJoCyYNMGt5LvfwWhUY4p2VUc386Eyn95EcK2auwD
biivgJVfRzMdtH3i0yS+gkjgzDm06s9XWTx2r7rgGdm0TjWvtvNZMkgoG3vZMzf0
LpPNbcJSK4RIK43i3LnEeXkcFmvxsfnQ1W95AzNN9oHopnwQWEdBiJxEUpHaPNdZ
y2xUh4vvewi4gxmRPfd/wLV1MWfEIn/odSYEgGyk0FbQWDp4pVSnVTvC8AWgY1un
sswjQorE60LduORFW+QAHMBdQiV1iRxXXpUoVHKGz7HOFdC70J2F0n65yc3SKjXc
frk4YljGpYUVyjA/uum6vvsuMD9+i91IaCEJR1JH1ZJkV42ZL2Hyz5yfyWa5XDIS
EEQHbq5z50lAckSxVrbFTxhoPrU800cyqLhXbjKzdgSLTZDv7tlkagNov7DsW96w
wZrGilKvQXxsGg/FNDFHP/ayC+R9LkFBRPrqYJFzu72/V11FXNbxFgXU4I28o0Ko
7oPyvfqt0f3UZfitlmnVgyKaQfjFY4pXFYI1M7fL5HzDBatP4yEBjfmW4DrG8ujI
NaDVlxV5uSCmdG22seEzTDqf5jHG5qAwiydS4oNHQ9STuR/2l48kHvn+iFsD0c09
FWdVJZhk4DOBf6S9Y/iqRt2gHxm29zZCPWOqbAwz1DyMH2195bXr3uJTRKzciW/I
7Nry76CgJuaddRXsV9h511r5C6RKlrSHD+0h7RZ6xYP/aCQ16/Rdt+jNS3Zmf7gd
tlAnYZdE+HuoEuO7/GntCKX3TSbxy0ljZBI3aOgMHqHqId2KwLjYHbQq741G8QK2
PeATf2G6ucv81xzM+qHWZuc/MmSXbKsOOuzQblUMKB2+wGTQuufs7msklucUiyog
MI2quYxsO0fGvSf1zlhwlDMPgRhaxWOFA/8oH2h12wJLNPE+Gbeq4p9lR5iLU6Wr
y1otVSv4bqjDf8zzzn7clVHwsD/wwNfT2uzcmLGWf5kaEuFEszBcTqvLYl4uPCLu
W9xPGSC7p7iAArKouHjDNWHrUGUqadhRQ5eGDoVxyP9a2viL9IEayJNgSc+eNSFN
Cc535CKkcaxI/82YTxSViaBZ+MpmR5KcKaHWvZm9tGsLV+lJB5+ezppsNtu+6LlQ
xSLpQY0wspEnq7zvQKYjcB6IRhbcTwlu+TG6ep537OIKrcr7h9CgnIXzNAHUREr4
5CziU4LLPdnQMtmZYVcrIx6CiQQjA1I4InPc17x8r6Pt1C09XJ2vyZKoqO1sQ1U7
Amrzcqdq/UaJGNM58aKu1kh24I+ht03fi9DxMz3RZiSqfiqdWNyJcwltEqNG6RB6
3fVH/dphjREkDR7c1w2B31GNM9dhBq06JVCr56hZw77VxcQ+14A4xjOvaIhBYFSZ
XEGFSVGmhesRrwgiD5LQgfnqAfvur/Cu8tQixbOMYpJhjYzEudYjy9yZmLb85nXC
tJ7OQ3UwBimyJM6AKmupcWPuzd5HsF8oYp307kipxMfxkPdWUyWzNhQSs0BuvQ3y
IgQWksrzgviWF6HjFe2r/kY8tz6w1JTm/phWVRFA6iKVCLkcR4OXlCY6BEfOChCt
+iGM2sU6mwnA3AQ0JBYMRnfFkv8p+7c3/jRTKtTiwu3vhlXMZXvP1KBOSwoOmrFV
tufFcEL+wzmoCZCPkA6qkTFVzc8E7lI27slRLafW/IV3LQIYc3xiL8TUltgf5qm4
C0GlUFsL615UbXoInEROXZn2B3VH8xbwz82/fQpacrgbqeQrUBejwiOnAuav3Ery
BmyhfVZIU4OJF/RDtjMmAV+mPJfJc+vfX8ObeI/biYEKgWsePzW89IL6fq7Rk8q1
4PiL1wDzO4jX6U5O534u9k27j/oS/54A3seyjQbzESpwE04dP8ltMAhkpGPXck16
i0DSjiqzWxg2s7Rr0/CMbgd/GlgH+w7U18koEcTNjTlWbEYWhS6y4ETENnAre8/9
JakWYbhtmFP5gLCRAfZa5N015lZJkS0tLaBF7jB3yXK3co/WYih+xq7YUCskx196
OF8lbrq6CqPSPceX6ExhSsjuOwEIMy+HKtRBlI3UsrgsrzYN+9Qrkl3Ho0GkJ5Wy
1/BUdYj2AANgVwcbG+r+swzX/Ecj/5G7AI2E2xWULEDZxe1fz30dgUmZSrwidPtd
xkz8sm3r3BLGDH3Ogbz9DBTcKApMumGqKpZTCMfuSMf6hOZyr5HZ4O+r5UOq7BLD
6AYmnqkD6CP+eHXIfrGlb9IrgE/eg1+lHyfOD3S0bpybSQ+NrMznkYm5Efd9NJ2F
nx/p2nPDUkvc7RwJRW13wbbdyUo6unIXuEzMMHbwM7xOJzmJbc5jivqx/bkZC0ao
wkM4Oqlx08VWODDSSFgkhebvqtauFrOY8vuKluyqxzm6cF8/SeW/FmYVwwixjMnl
ZGqqsgFgAJ788qermP5+RgAK/R3D1xgy57UGSnSBCy8D+bYhKnWcUu789SOp7av5
JOYRlrAy0+NsscG0EPLO2NzXC0DqlH1LSuFxNSR6t6ZaHP1pUXneu9DTL5pNnqgr
bo5KFsVFRBVDINPkL8bS+5vMsJxz5+ZcBYgensJ5lQkhlXEdsTP4ajhdYZLmpLct
CA3xvc7VeB7q2qTF78ZTr8WbMSZb2S34VeL9axs/PScTNoSqhV0AF0IvZ8owvnLw
MuUxw4p351CVBIur0U6adYTy9K+b81DRLzfCbTN/p97+P2ip6IJSUwF0GEIr8U7s
fRv9ZlHhoQ46MUWmvT7ZPa2KoVMXeubpDbE1VtGAWR3Zuf3KdIcsdisrAZBlTlz/
CXH8B0RGOBy/4MbRKvWB/auAVFbFukR2Gfik0djz9LfY/jNLyue6MnbxjUfUTKGX
NQfAWBzUqDTQ+DRm6C5LVyb2oRKZ6jYtIDRiqE74Hr9UdekKSAiQNaoCc2B94dWj
VlhhOfyZNSmwLRRAIzqZBMDjGujNCUAn9K+JZ3FZ3BTgcKWLhtErFlU/cNu7jMnm
8yvWPkNsGVAAdZ0deAvBLPmidTIfrNccl8j0oSOvbNYsZZsRK5T+yxb4L4JR7Q2D
5t3ekF5A+KwHxUdhJno7Su2ubhqOP8y36Ke7H3uG1MKEwMFXsTtrg+8vj/UqEnJI
7ZGsHvml4e2ZSz1f6GcgWQALj+PLZJjB4qmsl2A/M7mPffUBLo1xdYBqsxXAZ9EN
NlrgbDuv6zEeNq8pI5U2DUqV2PyDwFvuLIi6HUKj+7uX/HMsUIIZqnIyQVNcDbno
qmOLzQ86BjjeuIsrYHS4kV8nwHNCcCoqmzhMOKaGfMTtxHuYJKvNnoEsUYXmfpZW
4QeVl08XnWbVAt1YwW9RhEkxG+UGnIK8pj4kCO3jebFPiUwF3SwPsZ/xYDEx2XyT
zsTv9FLnchmEWJmaxSdBb1CLwFMdvYJAWtiu5KlV82T3tbcUy2Y9upEZE/57O/gy
e6SXBqE9r4eFMVP0zJ9Q5F9J7issXzDrzIwpzfbCxr7A4xIYstfi+0AVxNHm1tbH
tVjDdLU1Wq7z3UNjqMsDxmA6WrS9GRorE0PodZ5LaBRl3tTpqM7+7mr6fNUD54r8
yUN7Sd7dwvs3cMHnHz3SomdeeQLGp3Mf8SpCIYie1N0ZPsLuEBkFGiF25JoDMChb
gWm1yE6/xZmqkAJi5qzKZ8zX3ky5fXgIXbA85dtTuUYLN4FVaVdyZbHFMfXcWLms
jQ6JGb0coeg/G+iagoU6hfm8LrJwIIYNVRKufLbzDnvNhmZL9FEV1KE3g0mI7qyN
7VanlHtPkNnSeRRBNdAR5EEi57jfXLLErspQS1yN5YDVR7SkzTuRPynktxIjVYLo
HfPtpfD5VV2meufx1wQJf5AfBjjOzZxGzdxJMfZT3fXAT/FFjOWYdwLZPYww91Jb
5BV9TuCDHf677agrzw1zEtfjzbreUctK7ohJbClUBODkwt+XOdyY5LYF2K2ZvTje
YtQDF8W9V1ZvdbWIib9ICWnS5d4WQjDM667HgpT7fujfqMkF5mcbk1Wd1loigfRv
eIVS1VWsl/mKgSgJK9nghdiExBcgNXrlSC6Gl5CdfqaXNEcwy0KQYiEc9/BbZUCd
XTQXnn6aDq9ozQG/Jtu4uEDkyhGoXPE/ys3pIuU/qAAleCb+dEXviZPBd5C7gH13
Cjnpl0SvyoOSiTt1B9eDylH/oZOwfHiQ+TP91zd9b3HP4hfgUcG7n14fWi8HX6Ti
8UikrziWvFb/Jxy+cbbdnIqc7gefG682hNz6HtUoEMCban2cq1xNCGqyliCHM3jH
ICfm0Zr5TXQyzl86rXufSkPaheX18j6rRdto/R1oUVlqtcH/gsGhLi4I/Frclyd9
lDKG+YddEZZ2DCZ6o6YKEivw0n1TMxX7wU4mcf6bvK+n6OVrY5KS0kzGXM0TUfBP
aRCvc/iwoj21GLaHFRVYGquIKvxDfE2XOJXBYpGXrMIGncHZWPRI7OjojCXAhopJ
g24v4MjmY7RZzz0tWoDFha8t7bPqfOZhGNhqIlwZ9AVaKOkR/+LLRXVnKNmgiw54
ENgGCNSDRDcbItTR4N+RWR3uHzQtqdIpxD8hIZD9ucQGQQcAxgsnC7aPLaZ2msel
Jdn8pUkqA6zHBF9gPvp8JQ1/5Xxa46/LXS4SthsE8nVSmMj3/AZswZ+DfbpeYed3
00nF7q//n71xL0xi1wqxFej+Xp4IwaLICJjzZ5V+LCaJd90+YBIr2whe/5l3jJPp
EvF3rslX0XcVfP+wsMLpmsI4u+8o1zcwuvFQF89XJosioX0s7sIuqTOQh5XBsLbC
GgwjTxdnEDWT7PI0EslYjjuN4MvwnznA9c0joVqSxA/gl++kJqReFdyg7us+jx7Z
vqNHeOENOh4If8aWIivwDr2htIl+r0ZQdbbV6nnGrU6t4xPBxRFQ9xDcnEYHoEAq
kqjWsaKdhafZYNKyRanlozy8pD7ng6XzECkGR+0wouWZZT6/xvPPrs3bsbq8WeSp
DFdx9vxWc8Z0zL50nututq9VB0yzK5WoYiqpg988yZXmFSB6XljiDS3dtMlPHkRs
EYJoarS3w1VerZ8XYUhHcYl4rYyC1G6Eo4HX60cxA4FNhOZtLg58sNTRLW+0gK7D
fqAv8aWA7vfAUX+viTolCrKZph/olGjHmFaCNMXkota65hnI2pZz2iIsr5pcah5P
8imm0C36v5eJ2QbT0L6sbmlr2VmAqC+nljEnVYnRhSyFHBz7s7oAjSl/6KdrZf48
i1DCGANIzmje0ANdPUT1ALNApIAOCyJe8nw2ZjwZIlk0L2XeBd0z8PNaw4JU/G86
26hv2jygnnru/itTsuhAD2HXYKgYUG9j6HHJsH4KAnktCgevQ1rcddxK+z9mFezo
Mr+Mc1DzoGkVciBvVkmJNODq5Lx9ZLARv86rsBGAGHz965uy6LQIphvUiyjOYdl5
FQ/1bdJjpHfFCakRbJFi7GX8sQ/Mn9qkQbUUQf4L9Ev59Uo3B+Oghe802xwOgFBB
2GKP8S7V1IG0PSNARZ5XrQfgdA2T847jF3/xxrGt3ohqCWJwJkdKFnKQl7Rziknj
qsojVZvu1eXBd8zHA1jdkYUlQ2y07QufFwIfkTs9m71+qiAWgJIM8rLK1i4rM3xH
TCZQiMvaCspTztJGcLZMVOQ8e5mn9WG6czmDnSDHB5iu7TkuE89fxhfYX1Enp0al
kXvxStABjcXRR8w+Ug+GXb4Ppduz9dWhq5HalflyMNUni6Nux5IjeThxFjbQ8dpZ
rjVW05jNNPrtTYEG0LCXtvT4neO0kFnUCxfq9ZBx7N5santXa3kqJOyK6iHCBt86
rB5YBYqtBYHnFH3G3UdGUfiXiEaGm5u/UcfCSzHS1SjJniHoBaTOSu7/+xCEVr1f
CRVqv7f9j3E2aijWk5a75DG/0olh6XZZbl8gp4IlxXmuzHU44DONjgN1HqcbenVe
6stYfGM24ZHWYQuwEbrUxDRTcrzASsso87aABQ8kNVTGVjzWDemn4JiB3iXo6AQ7
TcNrL6efW+mJFY1jViZPJd+f9/GkvRRP6an5nbR+GX6TxW/RNV6CoIY7v5sdtfAD
KHWuFT4+Fbr4Tzhsnek9mAmPLuhYU9sgArUBD3s/mUswdACSiZopXkl1c4AtgflV
VgTZ/Z4qsB50c40QvvwI57ccLDEzcgYMCTFn1RaBXtWXcRyE9y/vqsCmjDRUWIlV
pR/uGnh24k7o6b+iYhXGJtsziz0IkSaK6xYyUBrow64WL1t7QSIxTcKdhG+kGv/7
zTG2vnu7k0+XbmjeWwcrCMfvUZOLugl0zFsT5OOh99n7sffxaQyKrohEP4ECay2z
nOyD7SWIn6XMfDk3iARMBCAKe6NMMS1UELn3DaSbcs0o1CcGxHU3uTLkXR2iPE9u
zp3zaVI9rUdJjzFGvnuP3A1HwB21D0pfDuY99PlZ75RdIqb5qpYCetngMLxRreXW
Y47XaYN9RMdPNnd7LL8tIb2rKLt6yD4t8j0qAbyPhRg/3ZZuqsliXBk12QSPQEEb
Nls0YX8TC7fSKTVQ+MlI8XVlEQC2d8yRn52Bfn2dumNY1qT+IAlpZwAeD036bVLs
ZDaG5IYX/ojDz/rGOCZdGtfG5nu2KCayF2ZIRCZ34nlwna+yV1fkYr/aRaSOCu3A
9EYdxgJA9lSWfXlnzZDgJdLniqdPk2sDZ/wVX3YWRJ+l12G/KMWvk+yNr4Iqc01f
I31tXDhKjsKCOehQ5tOXYJbyt9LkLb4MhN5g5xG+NmyKmo2p8gsqoZSL+1QX1V0h
xrxw4dT1qC94yQp7ytC5LmicvohxZwR80QNXW6wL94ZMdw/Ggyv6YfP3P4T7S/xI
bBGttmgcC9YqcNIvNFZsRscvhoS9j7yJHg61g0lPI2CwaVnnBPmwixJcYQD1vah0
sVqbqV7WkkjE+OPq+7XG9A4wpxsWPjD2RT9TUNhMlFhXq8F7bSYwi92LmCHt5dqI
Y3Ye1J5onwq59AZCzOw5cMv5M5QTuJQKuW0cASNHd1QdbMbjYUFZvqrplPsWh6fn
IAY9GfLW4yyF6lAd3D+21LzVs8a79b9GvsXnipy145L6ipPTHfWJD8hKy842ZdCa
dgpyF+crrjKTitgzVbpiXf4UnRMOKiFvSOPjOPUlA22NWvegzRXMrgu9YZsnbzmg
5573ae4cDpvbpH1fj18C5bEVsA/v8lVeNrIq6MKup/pAgXH+LSPdwGo+tYEDioML
Zr10zCsmnYHUobtHJmTU3gkpGQF7S2Inb33w4jop0or1AS4OEj2VlTV3NxDVpAs4
VUSldG08UiPugrMt/9XyMSKaiB5rWwTpBRgQ6e6D93Rdv3CsW4Aykxmr0bmFv6xy
md2P/0D78aXxr3R/N6xQ3MWz8rVQTCiPl3A0psUWQK1PE3l8pgS/pwt93iwyDDH7
hrMJMUvrFLHhcS0GtJsY3XmzgadFjOgC4YV+mNrSmEkKrxSV1TrAC1Otar+CFrH+
vI8qQA1wBpxE6UrGXEKD9/xQg4ZxYUCoc7bzeosCHCrWWdV+uO3RFA3MhObghvYN
j6T4+3Q2PJhZv7ob0Mhzw1at0SbDgjyyjtcTEdQQTHKikHmIeZevxC7F5/uPXcUU
bzZ+o+/8QdSft6T+hhBz97UbLouEVgpT2s7MVZmM8sRe6EGm0WB6hDWsdk4ToK/h
IN0REJJRLuWgRRCfDOOaLjWWye0uYuF/L2akAAjxV7h8bh7TPFBBrOd4teSVViGV
vhGVEVSyOBH4IOKFZhL4jhzTb5UKY2GtzE/P6ZeAGuhlQkKo+JKphwgFVZ+p5I8h
sxwiM/j2WeQzRWDEKWYWcXswfexKo+bw8lO5nXOojxjKBTlixA5xRaKrJYP30H1A
PzCwrpeYQw+Q95xLUnYPheoAKC8blMvlLoLqXGSJAtAwK2EXnRXEZ4r6h5Wj+cJN
VjPGSUWxJJWA+bLRNvzTaoyO26076ocmPwX+GCxB5dPR7weO/cpxCwCAUUDne8Z9
JjCv0DtJs5kx2XxV4Q4EbK7CzrJvSYzionElPZDDkeIzV82Ev5Mda7uqXQSS3QgS
869FwOoMQ4RpN5sMe/izN8tAkuHXbiwD9XpqOst4CR79V1+JIruJmowS9cUoP78j
Kj/cIlNeeuwVjNulEPYGGOQ9oFEQLhB+7WGkIUXhyTdsNeaYR1698tBLbgle4mPB
a/dDQaDtyF69hsgdvMaH4juyvs22AXLG2PDs2jnFKFo4gHusqIKljzT1dsJ/HBNa
DsS4dir9o444sT3eirTUV0qp9D2Sc2P/0OSVXRV/yzV1dPdmawlH9OyU2CLfoyOu
nhzj2Z2lKlLZP5TPeDqgf6u7oCjvhYnK3WLwh8PayZ9jmwF7qHSFWgtXe/9ixOeM
pJGTLnSkrcgZyFGmy7aOVaDCNJWfTEjfauqCHX/GPTOsuHRLpvSc4nVZ4lobfbpH
fq8orUTOks8/zGFV0Xiq/u722IkrbyvD5Tyy8GidZ+2jZYb5YGMBOn6cTCtHV2tA
K5jG8N6tguvmexmtRihs4PfAV/1w9Qzl179Zu1Aw390m/WvtKss0hW9wS3lEDnX+
BZkXTinmQf3J67P6ca2M0QBzQLKrkqGMJ4wys3mu2KULuYDLQnY7sy5COPSq0oBz
avsJVR49QOayJMa/XTLmGehB/ahDDLKNzJvb9N8Zp7a68L9qNQF45a09M/enYiJg
EZXrpQAIHHQ4V/EpsfD3d1/NBcbZV2e9QGNxcu+XkV1YuKCpOrl3Ua62zQK3/ScK
uh7ToDA48UI2WZ+a0JORD+P3EB1mAiUiKO2u56ccY/MuCkRg82r+HYoSWLL61HJs
3pJF1jhZ20SeGOxNSmk/VSYG8hLVAuysi3szUVz0dOY/ALB2B9gTbRsfjUHQPhAN
Qtpizwh5VfRuTZcnjNtiPhVQqcy1XKexblKSdgN37pY/nVFO5wj4r+vqAcVq2b4N
SZVNJaWOolwR86nZtT75TMt9TNlfjU9wrKDyKupt5uLNnCQ+24eitydY9mDU2wYz
QNUugL4wF9Y0QxmDkPzvTwc9ynXK+zmRyUhbNBfbS6Lrx2mM8/KNYCPadpIgjkox
p8shJSitrVp5pSavGXJJKZmLm2x5fzZUTnoHh2A3dIC+cUsM4VINaSAnYlpltPQT
BzJUhnqLhIkzCDXM3Yxv2W4AdIOEvQzF6y9qX5IdYA9jyuRkFHp4mHw2d2ScfOx3
bPGrGySNsFY79wRibppiPay/OKyMcSC9nVP8z1765WS3i2kEJlFWzUAKIubwAbjj
izHUZWDZbQ8FIv/NogW8El8wYrjmBXnXKlkC1TJUXOpOKgWlhOTqKky2SuHJpFvT
AalxfeRNHtqjcybQbyZQKoThPu3tC1NVr+01tJTscHP3SuYu/ryn1M+mByHbca1T
XrdcGfHQ2UUwVxlMHeZqgjsR3Sd5OGiPHH3rlhogHFj4DW8ov91Nra3mJlxJor0G
dv8i2zA+8j6McrtOpr7/IgZ8Szt6UVXTfEj3pE4lP31gAHmPDH7vU0rhe3W3vTHX
fY8Gzw6mLJ4rQDXi8cM4PYgOVPVzwRGUI7WicDk8U5j8YrjgzsVejnizMllh3Zxu
e3MqW5Ig9oXCli/Hy/NmVB1+cHlTVBueNGKK18HZQYsk/gMT1iZ2gk5Hhn5ZsarJ
pqWF1GYqlizXW+4yMKunJk19+gJMDpIZuMbgX+hBRI1y+OuCd3v6Q/k0hFt+t6sv
uzesmOeTUDHVjsvxMVm6gmGLVjHhso3wy9jL9wU05+xrGUL/21boQQav2tmtdI1b
LRhjMtv3EdnPGiTBNz7eyVZCJEGiP7ayJH0W10LWu3fuczApkEETV92GQ8NZDhj8
XCTqbcB9JWUQYhrK6RpWv433rN4RWvFqjmQxQBG4zLFxXbKiNom5XNBErl6905FM
ffXq2QGj7AY9WpxMngHh2JevBpGdZtzEerFZWQ7j50dn5AQxaZ2cioC+EBT9fpWI
+YRiHWgwV1OeyJm0U2snekbkNyCuOzZsOm6jF9lKm0ezaMie80ThpHHSTBaDKbI4
67cHF/8fzmh1PTK6NIC9Nk5xKP/v9Yk6zktRrZ1IDoPJWy61M97I1AaT4YfO2Ilc
dUrIjiGzkxMMXUWcELZ74VB+8wjzRO7nJQcxGDFaZZmE1b9ZmZNbc2VEXfJBQzU6
2VAZ+ru2sa4PivbXBKfmeKJxQVocL+Pg2v/cQ6MW5FZL8ciZ+TcXBUJQxfEiyOeh
x9GdqTKhnNNnO3+9zFZ3R6oMDQm7i045qpyAZIXBbMuJlmxhSV1/BjqFaKcFAEKv
H7SbPRMQT0XJV8y3W+OYpmVMThDFgaBxqBFOmFNcTn7kibrzJf2NA1G5HkDiwdCD
uYOwzTC3JMxwu2b0vfPJCSG+i9jBlqkwIUbi+TKReA9AwHt+2y7kFpLh6CIMiQLM
t5fE4tCNLxyZ8HqUIo1bxx33veshjuaFtshlMx4yxwg4hP4Iz5VEJnAit2VXv5gb
gBn7KNJBMlunc8KHNv8Rbfkivfh9+P7Jzt90IkhKOtkq2sIz9o62dW9K05UkOW7v
h9sn6aJNQUTfrP2P4fIfqB51Ur06t8z/XJyflheiTlRCLqU7eUhTb132EqLxb2mF
JWZ36de4pQHqSs7MkoJqwpJoEZrbdzjHYiU5pnzQCkgeC3cKCpXPEgQtkf7K7Kmk
jftVlYo4pAO8u3A1XtoImc0glWPWX8pcfQz5x7aX+0jMbInCh4krk8dyKzm76Skp
ajt1L+JYVt2qDUlFBGiKbayworUy5bt9QkZn6roueyMt8PGIllcJR7oVoe+B5EyG
zpa+4uPaWEIo80xiSIm7tFXIbEDkyHgsPnwXjOt7ckGnx1C0EGYJ9Rz05W4pDvwg
vhMa3MmIo1lAcrYOuYEhNItKWixIXz74GyiEIIy8RbrtgNPRNQNRUocKwqifBBXp
gfNwNbFSEqYZ/cO0er1JjuldRiBsEIM7tjFh6t3KyXYriDwBNPr5wTsnyK8XvIWA
Fj0oFHt5HbMe5VQtUJMo22Qg8NVL5tTl2uosPzVV+UP51oSfc32+rVWWX6Xs0V0O
upTa7SsQSnxZHJdoo7qgwzeIJj3klStuRlR/544aVnvNkBoyK/QCTy1I4HBVnTxZ
QtLKJAUrup0rig3RRY9ZC8q2gpREYYQeVzmvzKy3p70MYpZew0dJq9c70X8FulKC
Hych4nHC0FD/WrcRB8O+gn7e1PLLaObP2c0tn6Pt6JLRa5b43d9smK9XaBZ4QU0m
QVQ4duviXfGfCw0EQFDOqOnTZldoY+RhUosBkCHVj1F6PHnLlXRv4CGC/4mthbtk
0HoCamldoGrVKH9xRn91igusGV+iu3j8rQwSTkG/7Rp8R95CNxdWb5niJOoa2+ug
Ncdt43BybZDZVPiEkqtb2wQo++lJXDIzai6hUlSGHBgkwqf3mm/4AyG3SVAempFG
dXSOrZ0blyvkFsteyDbNvVHtBT6Xl9Ne8BsYGc4TArHbXoZvJbiQhrbd6i1EjJqG
H8zT0u/UhzMkbSceaTL1DA==
`pragma protect end_protected
