// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:02:16 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
fjlaroST+EdTrOcZhnzXbYfaceTlykDkx2GPrRHzGnUqDBEUDcK9kp8HxN7sOJLw
Xoli55pmxlp3SOqzcorG6ShotZoGsYvIIlkfrbrMDfLjgDEKHR+ay4Qu1d6K0Oal
x4q7QNVpzg0QlSEpRmiN1IBxmIm1MGXcN0Fp1WBETUA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 28816)
fS5PzCZR8FImxL2SyX5B2BFeXYP0O5SI5qGdTNKTMPEblg/5JQ9duWtrdzPAuBKP
uYsSZyTp48fUg7VPbl5w1OzqENQ+QnnDgez2pcvVGayQoFBI07bLevP6LqcJRpYu
xCUMNEXGKtMexX1QxtZ/bIe2n+kwJhvAbgwroXIIGMnT91CXKjzutAC1Xq3RDjnA
CylOWrP4V/2rXyfwDWA/7uRBc6pomptk8qN2ukM7tJX5kPv36dR7n1IS8ALhjSiE
P0wcQbTIucMXXu92YJCEyNYYWmiZ0UEJq5cTa1teMIy+Z4+3adOAyaIKFm4AJ4Kl
hBGGViP9FiKLGW5XPOKEaInXFbB5/6joAvGuddaNETrlajZv1Y6WWMOYiDHPQR0c
3toSWdoLLcaRagyr97UOODNZHpXysyDItmItd/VSGWccwQfsx6H9z77OcIA3XrAv
Mzs/QpIjH6g0sEkeALUyxpxeRwP9iyJdvaELKxIpNnEIGslq7EJfcQ5CO+lLo9ZL
CM3p1u3zMFtyugO4r+T5Q93ur/XRXJg/BJUO0RGbga3wNuQEW0VsL+DRXRoSMh2Q
OUD2UPwzJdRpmBlZQhcJjDXeo9rf4ucHhIKuiJltEHSTk2YoIrQ1dzhR8zLpFfpS
FEJYndjZHABW7Lbf7Yxnj0pe+5AwO3s5a0WDq2LFbSISKsjFeMWww3f1FCdkTLGm
CmIXrevwISdb+5aiFr9Sq0aqPxX20xDOZWvPECiw9Ld0YWvRqfqT/MI45KdWzE90
splIfQWG15x70AvlaRPFdVlyXPpnS+Lsn9/NYmUcUwVn3g19FDOAN9iG8+kQ11Fm
FeGMxiEltIFteXz2wPcu3v+w4emSA0bfwE4319zMsnlUFM1SFVPzWtKRMQ7dNDrf
0T2mrK+i8LVfSXViYnVqQweaboC/tY2c/zr0w2pgpDh/V2C6jLaYVWknowmxR2Z7
5Y41Gq9RpiLIBdPr3qXjt8CpsftGQF3tkF0tttcgsbyrKJxGaRQi4cixmNWL1URU
1qy2Z+KXLLoF+0AiiOR1fjCWG+d2898P4tXrqSh9Djpb8HjDz8pCYrno0EAQy/Cx
c57vYwcrRUKuereBxD79lwQfl9SBudj71wXVxAQonc3/v5g7mT7elHuqDwbQr3lR
TxFJ3nWIYwTOO9AJpIxZ8hFAQRjdUeieqmn1oCMSvghClPe4IpvHUB0fl7Qt04mS
emvrSOhgbHCzmVtiKA15IOS+JtnywCFNA/vES/toLbG7j2FB2ZMjxGSk0rs2xLxe
tpCrPNBVvsCPcKbf8KOTX7kglTCfBGdTvH9Awv3McLyNK2r0HTaveuX8umihYbVz
7kclmT1K1wJJWJRq7HXbaOI+PFj+RX6gh9c8BibQvH3H2ijxkjW3hsc8j419LnZj
IT7aGRV14hyJPjXi5JxbYGH3QGJd59r6L0UVORHbpfBljagjeBwmUqViO0y0BtPr
4zw8rmHeTk6UgcyM5gX3SoWYVMgTVAIEMSPR60JVTqWvMTqu5Qyte7D0JHKvLJEN
Uo5y/QVaorRXuTssOHLPyfDok0aNrAzFqodhazmAfmIGTNegMeBFeqfkBrQpOFJb
ya5VkBjp0ie4qH5hAqzOkNGMgJZEX9ZiH3ARiJgd9ZnAC80pmgHveRhYdbMYwDYr
UPygDZABBDuw805sbwjnj7mXkMrTr4tTfNLYqg2uYF9YQKihkMnowzGgzuxls+NF
/TjhzzYjCoRKcTwBZxHy6U9gViOnmTYE+icpxjHxZV8ZiFuC34gph1CIHak7tSOj
r9CybUPgnwWVriqbmj2EykaksU59Zp+g006gd2L6L59nL/WQMRE1mJbv2eLxussq
FeBUhcUKheQVqt+bsywOX0XhdbLsgDPwcvm1AoyhE2U6NxxbGm1e75OcEQbYILIK
NBVZR8lSFNTOP7C92lyzxUyGV0f4ltdnZxVp5Cqk2aoC9KarSERj1h4TrsH2L5is
udE1ouAntHSSW6SKjNqtMrOyX3OoGhubEBnrHMyQ5kbdcMnJJzzmjppzJR9dySG4
yzJsUVdJiaFwqaTKvoduF4ChPCxZhBm0AIzQMv6b+bCzO9LGK9/2CS7ZOWd6ZXtM
QBT5gAqmPTkGw7UKUChq1Sb4QQrqhtT1qIULfCPqBAMvMYSsoILVDxKbbIKIUumL
eoa7D79aqlcpy4QSTZPOCKH5SwbH1nP+4NnU0/O/rb7hGfX/Mad6NuZggoF/mu1h
j29nskjlonHW4e8U999VEE056JSJlbWzQzeM0KONkm8DMs1tPBSErDSe1h8d9Y4w
TzcucyZYrjgulBjsh7BqRfRON5t41BNsDsZO1b83JlEYw62JKax+3VTyRiAr5mI1
aI99N8dxJumRJqMVOsBo7fzVywBPhkInaA9kd4pv9OKXIm4AQdxdsF37V6qCYO8P
Z69lL+d6s0duuo+8GD2FUhYcX2UqUeAAhehUb/PHt+DuibqSW/6LkQpOCTmbtSPX
2Wt9WY7ZQKkOKUcxxVipbu2EAu1JY+heF0j6LHmRhLXkG5+Pj4GUIpet3p+fX8wd
EG02K1PsAaBjquDMu7ZsDvGF4dGGKuv++b3AvxO2o2GY0ji8+uRnIBot7yICuGDt
G5wTlxAlxJcwzMab6laId+mRrAmBh1IiG03KWu1gvXJdGhcMVl/zWcGWAaXH41Zy
KY0Cywunt8X6ZWb2oSMBRPqG7pXt6xRvZMKrbyQg5hNh7btui8DyQkDGLnGAu+ov
jpvlvWIUHBEwnVtJXWN3wKu3IC3g6mmwHOM0zDFhpzsq2wgOwMi2w5eFFarOsdgV
a+AhowrVLEd47IWUo1eJy+d9/HsssY2BK0Qo0Pei9Od4/l8eI60iyuiJIZQwYCWi
H4AsUTgitN4eMCGJPS3iG5n2Y+e80YvxnrhAPk5BTZvZXDRyNkVmkgs9xulJuPVN
+qTNEkjgpqCXMiVxAc8Q62R9KAZtAfJlOu6CI3vtZHC/+E1MqAFX1gDNaYyVfu51
i8aCtcSPC6tpZZ5D5maocfByFExKzadmGbNDMN1AJQ6BnKtIZte5fQrq6G2Xe3cX
nVx4t0R6r6f3ldoSi1fVrge623SzdPxbvyvKmRi9OYojrBloBgZgYZhvoEW4p/CJ
hFXT2Fc+ZmaNZrcIBWD0LfQJkhLKsVYi6MW1o48iKL7f0+IMZwb+x9ZcA2Oteliw
JdvtZSWVdxN8ztfaxPvNcDdLr1TDJaLTwD707AGEe8F7Hb3qWppYFA6WQk4WdMuv
1RYhnEV1KfLv1ikUHhewadCa0XnNVl+PyyuCJzKj43TZIpcwU4x20hhwoTHMB7Wn
/pBda6PKIaz2e71N8nZgDvdJlnj4TPGhBCNuhQx3CR+NwMGU0Dl9EFpul6id7oFK
a2B50XF4yh2koVWylmZPnNgbSQ9wftgQYPQ4E1j9J0vnNxg4WBzSMnQVOr74uK4g
eXQINJpAx3qXl5ZOLG2XV/XROxR71jOwABdhMuWr9IhwYvhmgTWNWceHnbWxgyxm
+2OiKFJTCGEiGMgLOlCmXsBs0W8AJ4+fygw2vH/ijfN8BKRD7UqcLyQwrH8OgneG
Vk3dRnmnxIM5XfT24tZtiX651EU89LGV/Lf+yo1vFA1E6y6gBn6ASRvGjdCi9mHP
OZlNzKa82W1x3+7YFLoVad/WLCrUQ3ZkdX9k7dr2it6fMciCy6JN0FOPPMETpNMQ
UFPq+NbspvaR+Qe+JakgQ33+ChjPB7HjbbxT+OYjREBHBu+V3yTWxwWhVSQ+Lt1g
uXJ3CdZybL0z+ddeyHv94KNMpa6rgEus0/tiPX0QVFk1uif6fn+NNyOuLPi0Fh0v
kzVxqs9rbzqR/BJRArNB/b5zFJmBlf7S1zhrGLSwkOzmExtDGIqcC9F8xst0qlEI
5JRcuSHPA2Uj+dDwi0v7I2kb989tiMORu7OyKQRTtwVoHHMbP+OquvBaqYvFWqZ9
17TeWl6GCVw5F/T34zn3kUR9Xzoue6Zv+6hpbRQWT4YMZ13pOXZv1CUUeFFvKZ6D
VPs5egcqBQdlMRbH4KOpN+r0S0/Kb/aHA8cVI4UbjnoC5daUKi0qzwVijJJE4XwU
cUHELAc0maDQ2I+QUCsGE7B+vZO5QGQszzW205XKuV1yFca2ISxmlswy4Gn3ZQD9
S0uJrAdmdA4J+xEg8BiuP5dHODTP9oQ0CV67VUZC5a0N5T+Jf0KTNwqCQRYNQCCe
RPQJiomF54Mj5+LaGvyNB7az+fFSpVrVH0wVWU45F7fK1U1Od+z2qWUm1yc4mKGL
miDJ+jl5uefH+fAaQKuyfjNctFCh2+RKDjZ437/FA8ayiHCxoqPgAgwswexNPnX/
B9UKjRSNbmdjnTnhzAqdSoAjRnk9OHRQkS0Zjr+wdbA2M5ZxfRyKii5L55UzPe/g
XpKY8b/6A5bXIxgRNa0sOP04ZZ1SLnhxvgKlEAxU2uqXQsrwX48KFzaaG1vSJhxN
82AVkajMzktLT3/TBzcnJ/K+aecWYhUiDxu6qpsWDqdCpOw9/cVIhVBXKl6Z3TVr
QNs5bYuSASn4kaPLsP52aEkV5TAs9LtrF/fcqVC66gdQ6Bv9llPQkCtGHJboTF2z
j8J7yZ6RGhW7FJSjMAf6SICZ5qSjcypogQbLf9bpHz3qAvssgdP7ayJwSw6VPGnP
U8+QxwSCRSO5hjVeVch3gdDfxr0Z9gqtdIMOQrQZBKkHyi5q0e7COntai/2Py04M
Tu50IDKdtyDdezgykakvaDWYt6Zi6q9ftjLBmrtpg9HfRouNJzpGZuuM9JYNmnE0
kSHnnfw2WkYgAPbbVUlH93k3YSyFma3aP19ghWsyrwhS8jbyVA4fFps1P/RRlVAp
lvkmSJF6w71Wsz/rWZP4UQj5ALY/r7OwT2XtEEbTOSVw7HsbI07cRExCGU2n6EKo
jO3bgqw5GzH7ajqt6bhatH9ORV3U7p8uTMzVrM9w5EPsHkGtSpulDaPzP6jC53JE
SsblxQjJxn9UrmlIkd/QfbmnoYgjDa/Cs2HZxR8xXZBYr+CBCvzm84o52IPICMdx
l1xhR/DDX1z3EZnkILKnsJ9KVzRJEiTD0Xx/9wZY9C96PGe6zzcFEcQffPuZ0lPM
hHadY1O//g/mZfx8hFsI6JxZIBzA6hui1R7FKQNA+CTtiCf6RD3cdiaAINnlWdNn
rCBNpR4QT9PMands3c3+kTOvZxnZPn5ML1NqxRT5FSXiT0s/oRaXbOjcEArxh6dI
BdQmajof0dEnDRdFz3gKC8wNdYCH7swErHLs08NP9lhGR6DyAa7a4jvw6TCW1Qw4
XqcuvzB0hHyrIFX9NIVMO4O4MjRShGJ68n+biwiv4MC/r5v2GRONzkVE902PVgY+
VIVsnem///vYgKT88PNAmTmvGMOjDFCB/7om7Vf+PA0VOMdYQ7wRv0wq3wXlP8Ki
SEArAon9oI3WS7P9nLzbtSTwpBjuQfVzo3CDvhNvoSlLU896GG36WFlzuqDdoFvH
k1l2F7+ohN6w3AWTh1LObz95MoQLqNdBHTWdZDZbtx6s8qD+uIkrzgDKYNA4LhpL
hHI1+XTpH90ieOJTutrV5SDHmUgil8e32n58x647agBfrFUUWdV5wd5KED5Mb+1+
0vuWBqEyr6MStCIrARUgBacgmMGJ0K9fFn2s2ewk1Gb9qWszcPsl5cddCXHwjOEJ
0Wf1w32EIJIC7O6ZbzbiEeByvrpt+UmApj3+L8fyoHUGMta03+PcGunTMA1CgLYX
Fxo7r2GhDqAdf6/nwHd3mVHkxgWoCpTmy4KGktUoXXokgJe+aHXCmm5V99LrEkvZ
q9awRka4mszlpb24hl6LfVuO0Cm5Y+SIkIFcnMyM/81Be79bnF+iRMbTpBLMDC+U
Urcf8yfuT6i4RlsECIi9GSouyI1oyZKJxslblGK46+YU6f1YjP6FhfslOdNKq5cJ
1fVgjZByUesyDeVE3tV8m6Ht/n35OG2aFZ5sePmF4khAOehMftVKWLGldjmHEstv
M0C1Li7oAAPFbu9Jmf1TA95/G0lzIg/vpj8/r4W8tvGv3LwgIJ+pS/3g43ZPXRb/
bFZLkPN66FWy7a33U6jB1bTRAREjyZVKqmGdsBgUdsZMeinQV2GM3u/2OPmS65W+
m3yd+AjcOEflArVi3+1mHih+gvZ7eU1h3EKtgXkMrzfIYbCoQfMSkIZ6os0zufi7
FHrOEaDfoc8PfJD35mv//LTOyg5O+ac5oCzYYPnjQKxjPDS7lEvCXMy9BqLvWAn3
z/MGUHMgrtCfuaHAEBu6YIpByXEoT3kGyxuStYCw4hLSATXYGdIJnzTaI48EIqJc
8i1txrcj1ehDhDR7GLCMSuwMzhYStgapFMbfnvxDHmgUKLlxq3ea7Mk9s00Kya6r
fqhU1ck3hwNAFHeDvIHNpfZW7zUebnMYvIPXJFh6ANE9Aoh92F/yD9ijwThMkfki
jSl86KeSPAPY6QYg0KpSifZfSQrtYX+RY/Wn9rPDlX2tl7G8/amm0FWpFa9xbnlY
xC2vcAUAGA5c0ylCTAueqdQjfXYDoHfVu7iCwFP90KHF/13AIa2KxWjqyA/nvWaE
rtLH672DoiU7nnVHhigwdutZ+/Rpk5oiR3M9xJCOxP1OG0PwIXpG/WUfrQ/Al+Se
yc6iaTvWzYDLVYthprotHu53cFKKP8b3p9DdQO3E923i9B9ibbzxq0mKgZRq6XjZ
HUpwgT0aU5P11SwrEsSfLxyYAOVdkEHMlbppJU2Id5+W2VnQhpFTZ2trHsYaAPcL
ROZvC4q8NWi7JXETB8yphpM3wCGRg9WRWtt5/fKTPWvLrKcDOJieTbd6+AzXC/i6
UKoh5x6u5dYyyKVimRSrmauB4sdr44GYkArD6hMa+8kaOfWs2535Ixi7QozHYY1/
DujL/peASZmSYHNZAFo4iG5kn9P2qEUSYf9E2jZNPB1p/58+m9T7nMvf9VhVmIly
aggB/CwQNu8XmGayt0NgV04tku1ZkGzqXIs2b/K3zZhSxLNuBInmZKoJt8QCE7im
MNa8bqo0yxc0WQUJ480gL2RrTO3i82617zEMOrM+m6ypDZRgZc6Y7Hi2OS4f0MlR
59ZEWDW5U8IgkLWA8JZJMNuf9MCBe3tj3Hh6TaCL6GYSKWA1D3Asb/sLqTKVGfJ+
8Kb4YPC9a5oni2aWQqpwaQ8uFFW/X51ORHgv1JqEKF9d8XhXaSFCr5roKz3W2Fo0
eS4qneztvMlxGasqyr0mAiun4nCjlOFxWuUKaSMdVSDNVV7pXdvVstBRGG4OkWBp
aY51CPYnRJ6aFFXzj4BDD7fSchvlCp7W+u+sQZW4oGlfKmwbhIhj7mfsjJhnHdVa
LpsbFKxbw6fUymdxO7GM4KjmKpqJ4stgHIoUayArzO0eJiuF/Zjw5poGuznilf5F
KKckj7z2h98P3KXfba0hFacIxkIn43tTDhIqdVqw0M/h2wxUTVzCyE6oiE0swbyY
Es7T8gg5wV985n0B/LC3ZBWwsvfJdvSgl5iEyfQi7YlO65ruraQ8510fvrpBNayd
Lh1rIfFCztRi7NJ1gnY2o6mXHj2+7lEO67NX+DoI2hursevZbGMtjcN/NtbDGLrz
l+SmIxFUC4fwD/h6gXQfzm9UsmChjH5GhDpszo9Pr10vkT1D4FWJziZpaLa+LEGl
81GCnMT8LW08IMxX7jyLXs2tAkk9k5yqIxmJYIdrFmThRhUTJRIrtW1oy6SqeKM0
yV+dfhVHma8tAcK7Fs3Ow/ZlZAB1pF/lmEQtg9wnFdrGckFN5fpkQWwDhfv1yxku
CHDBBZ7JVKd3VSzY/+CfnqQy1I2Py1mE5YZqGWXl64VofgzbAAgbIvwOEKUUQxTn
wj9796sy6wT89Xy4qDZux1F6XvlhNgd/kYe/gqwrtndmEs5npqLU/GSuWiCT7IaE
Um7UNQxJGiMQsiTxuHU1bCmz9bJsi+4q0kzsuOXa50Hq+Zcx2a/WqhNmpE4HPtR4
ejPWR6NPGBci05+klotOUeBl8KO5ENe1Q+Sh3bHd0jha2C+j1rmVfBvUvGrn9G76
HsXbpNl0ZhF9eYh+JhzpHAP+ma0NEbwFdB1Ns6oES5WRh+HibpwupeAlBMsrbIgy
WgpJzH+/L+KaFdz3nxuKy0h6RfvdeIpb3ujBLVbM4M/YGNH11FyzsRr+zjrvZmrv
YwzAG5XZaE+N7xIof5J83a4e5ZQFHhRXhXugLCOdZb+yMCUJoTMslxK2tm4tviLt
Dg69kwLghivgd9cCDZmYtN/SSM/EEcXGSioH2HFqr0pJ29dEH06MnSVIXTYg1h6K
TM8WF+kJeh8myGsLtdQo0tB6o7X0bRrKuKUh3HtOVfbTUq4TaH/uq4zR11mliAxl
jMl6JRc8PJ7MvkmJ377wmhDQqDObRYSvzCTtj+qzemvw4nwWKnLbn7NXm16TKOyk
l7xoHcuNCHw5N65kq4pVvDH94zr0+sfDj/bqEjEUtS+ZDdjkQZU5seo6UGmO81wf
NQxmLjBg1ot9U3Sc6LCkXaICVdjxpppoIgWUYFa9OFRhbVQyTz+BRE+atBx8RElU
Adc6qqe2PtpKB6pPNRC50nVBsGQyXbCUYsLldNNnyKCHHuGPf9DMqDSwrKBG5Qn4
U5+cWvYpdw0L0ByEgyMAWf60edSRRoOj/PotpPZ1vBm6ZZV16W6j1dcb7DBTu3T2
L9yQ+WsgOEl5h85HP8VFT4B2G5BewrOQi7trdURJnuR1KpGIg1ZDiOZzZh4zmW+z
iR8UnocjN2XiGF+7G10ZR16xUncY3iCVccnErosfml49I9eMUfPXAcTtmDMw4/2T
u0oyxyr9oJ090xnUk5CNmkQWArqBHT3LFz3WN6lsdX7WPMoanLKbR22hYi7r6zks
gFC1/OsE3jQju1b4e9WqCvY6s2bb5KKTT0WDBV/boFmNYYakOEA5IHMCUS/iGEwg
WYr0vMP9E5sJBmgO0uKJJ7CIDmZBOiKs6PEqMzi/cSFonMloAZEqJUk2SaEwbIjK
PBlbYvnK6HAlD3TIgOn+fiFYJDDL8XVI36Wu9LLGhfUeEdemumfyfUWlelH41nhN
YyVE7FcPR3bsaN50xHzgAbLguPkI5IG0YWls0nH3Gwvfx2lgmBq7ja8KzVqEcnFz
3HO/hoKMsVHNys1YcG4Qrlsb3lkmNw5nvijkMVjparOeF5FKvgcm7Xw2aKxajLSq
x7grWvq2yXVYWH0oem9vuEgQOCqNzPW+mfEosWwNKH2VBA6BUcuWrUgbfB0wOvNz
+AFcz5AcMP60Av7eBQehSugoecxD/YQQggs+PRABDbzAoW2azpbx+Ieb9Iz8l4qZ
WoOfnDv2jVy/venOyN3D8Utcz7ZQ+WE2VeRR3+Tx5gM8zP8SIDAZmMfLDZUoGKPs
dstkgT+aVQ4Fpsv9G59OF7D11/tklTA2lXajMKb1ddMhHeid/wn9GAZodaJpbeSR
DQxBXv1ubBhFObaVDnNFjTwlBqfzcn0MifE0YJZX6pi8dFsIocxpc6pgaAxmYre1
jVdOIl1oQ6rXrr0a7YHSO5wZppvYYIoqiboPpVrB5z5D30FWB9OFvlvuOEcJqwK2
3GQZqDsfYYTc6nsO93j5dJkDq5Gz/VgjHUqJ16pll0G8V7KRURiT1MKmflGNq6sG
YGVbGrJUNltf5zoH6b5lGDbD6kQsucSZzYj3oWGMhIMusiSSZIoMLcTIihaSPBTq
kv+9yzB4T1WehHehb+WG4ODnRy5ADNRJvfT1wdgsyA9JTXcg2BmyDuZ0K4D59K/5
VCRi90Wlv/2dAZ5pXwH+qUXILE/ZQfdv/IvcfEr84R1+wCbgEhqEqss4rkH28u4H
9Y2oZ4pL4TMqcaFeEG+MsRerIS9cMfLxbq1FiIpKzFAj01g11aE9WddBrt6Mu4It
nb+soYCZpD8+Z729zXLXLcEy01RhVABg8AXD41QdV1b6n+d+oF6xLPqJQC2nl0pL
KB1X0NhTapPmviAfXFlqL7MHokduKiQjJLJEwAF4v15eT07LbXhOgfLum39Q63K6
/jdjluvp4Oy+54VuiZoelMq4BEeQ/6MkePXKHFzLcAY5wu8DttzbgbOPU13tpglM
R0Gr9miZ3IbyEJL0UYgC88kmfbr8sFyBUfQy+1yFlWnMNeClr9EC3y5m4f1PA2B9
vkvZyb7XtH5l22dN2wyxsfr/biJJQMSH+Xz+BGjiaFKWiwMBGYnSjrg0No6BqIpP
uNwWf/z+aQ0w1LbcodQvqJDxVX0iCOc1pSF3VxeT0C4DCv47qGWp5lH4062L4P/K
4UpgMA2tK9/cTYl65NqvSONb8Eyw1xO9smk1YKhzMGtkY/BsVn3LoqUriL/PaCYc
WxDks3BMW1YxYxDW2/juqNE1+jkhmiBzhME/YBfzIwyAk4IOBBvQHJMoD9zHZ6ER
u1x6gWgr85FNsyjJ6ziU46z/oEVORgRtgpNlmXH1VzD7+t/o8O3HEpyOht1TO2dy
QEpZs3t6yyxWdA0wnCzHyeWKcRDTrXjA4u6Ojq/uNBsv6/VTNxpqwMrdobEgJeph
Ex37I22qAF/Wf7WQ6nlCzZm6K6d5a4L8lnDJ37J183ZdHc57TxdU8A2OQMy41Gax
sKxvFeoKIsotM+3gQVmXtt9KVaqhwQEsCyCMj3rB06x9wICh/AzX4ShwAin6wFlK
ZelPfPXjDDeo5O4cphJz3t2LjkwJYFpd1AMmgarOL7nZ6+layQVONPJChbaVplWn
LUQiL3NiKjtcQsKSAVZNhM+8vA7UnL+m0zJeMQN6c1RGZdkiaKxBFVnFpP7etpEQ
RfoBxeyzMS+684NeaEf/sr/1EFRySVsJf5e5F7Ng3DpYHQVCj3Bmfi4Nuf6bt+17
urKmePvz1cLuCHUFSnCbgenkkxIHtk4DnU9Z8aXoS/ZqzahYF1LfeRJJ/OuEIVuq
0mAMxfdczcHp5LC1vgi9kIn+yeJgqNGZSRqJpAAm9Vf9Pf/ynEyVsI0uZpITBM7A
sBA94lIJSGUWGU932+3LLyzHF6t79Dg9HLo/vt2Ox20JCIuoy67dhGGzb8/AmBJZ
aMS1AHoH1tWJ/R6kIF6R4MFggYDVbs1jq3YZDxx+re5TDDWBnDSHAPXIOF0Sz4Iz
9OBWg7kYhqHVBkw/seNs+06ZOqB2bozQYzWWRLiHivXKjJzPOZVeR236MUzzWx7n
CM9nUbkgoTwAe36NTCG33NafZKRjGmVuaXxHaExpEYp8X7iHu0JHFtt9e3t+ViOz
+vXKl6ns9VLeBpIvjmTrL+Ky1SJgiGlaVi13C7akpCWsKRCl12AkKmBsSrgNITwm
yAjDXEr8T1GT+oNIYEFQdo8uuBjINTr06OJ7/RTjoI9Hw7C1+UF4Xhiz68ZU5tX1
04Ai30q62QE4AyTRNClfZGI6FEoxXs1uuQ+w0m+SDgUaiWQAXa8Va+6hPIuWkD6p
qiTkMnjPPXmE4FFFiiISIO8SUKDl5zYUsX6TAa4gJcvlsK7jlx0byasnfmw3XFvm
/acK63wt1wQmxFXVOUvxH6E98xnLxoCg/aJNgQ6+zkAudn9QVT0YlUmZ867X4Sih
f8e/8K7OQ/IE/9TYl/a/Uv5564sdCSuMEdo1VVIGok+b5VkZcYW46s62uZfGzNGc
g7uXNbg/dBiouDug9ZITxlsW2P97PPg4Xfu+Z0jSeppoF47CS+EbW+eiPwGbfl1C
tULzInYWqVa9h4cdPP8LMP4888r7vtkDv1y7tk7WetXPzdnk5rCI2DD6MkhqpzPQ
KhWiJmaBkaFYP11n13HdWTPnD+iaMA9lq/CBjV3jLTIMqRr2TNr0xRI2zeAQ2aJe
MxE0bedezAJzfdzlA3EhlvMqyomaDjHRFsYNj78CGKpABxwpi+edqd9TBWyt9cRR
DIToEIw2r/s4Y+fKRAqFWQlJLIubYTZMkU3bfx/QJTUYrwaKLTjQeagcojk7/Zi9
KHwPGhH64Ww0BGS2rVcnnUrTBuoSuQTUnI/isaCXuBbXsNXadg3HaZ8OpcsRZxxJ
6Z1itrBecWcYpUC7mn74LLun/SOm0HpXiUonnmDRJHmc6NJAl3HkIszOiXbFYI1O
aWZlk/rQDFeNXbmTjUxZOYhYoOk9jChJZAjbCs9wz/KiW/KOECY16FoQQ8+ZhOMv
NQ7xsLVUrE8+hl5h7rXwuaE4LEW4HTUdHRRmMTqx6MkXdaL42/P6QDMGwbkO7bxp
fgj7HH25401nwnikdyNeu1BUJ0D/YefAiQrlbNfPru9mB/RzwKVhpyFf/I+brKQl
SgroTYvprD68lbC7SAiwEiKDWsxiTny52on3BDgc+oT7sg+SQcTjZR7YZdSnOQpL
ZSMjhv5b2H+1dMi+Hvk7Jkda3SkUG7A/oDCHIprFgAf2L+Fqfnxd7AqWJTaGApFT
9w6TGx5ZRisMGcix1Lb7bHitKk1pDzo/Nq1prZBSB74pNhL0rp0c9+m6w2WIlxzn
FW9gUkUQmKrSr/Bn3PEywLDx5EqSmuFzlv2fJc5cnYoXXrh7q/OBocy/C//7lWVB
HEKe6zUAdG0AAeupFDnmG2Ka1eVvywyI5C3FQGJMYoyozGaKUNOTgjEELWZ67Q1E
qnBgnqqedysQzAFCzNAZzUvHu/uj1BMwcWn+rfYa+khn9xDNeL1FJJ5gwK/xLjl7
Xe2iERWO+H0ZrPpcDFrQ9HEwPSnuGsOhlsPIjT/uHLyLJYVnfT6XhFNIDNAiwVsT
Z8zj3Jmsw2vTFVvyTRzfcVN8z/QIl2E41Q7+cD6Qet/lEBui63JlfQ2+xJ0H7mG8
y9xyrhbw0jAHee5ThpGwb8WisnyPvk+CSJsnjT0koaKXI5P0Ut1ua0ZBAIGdTRNn
wHJ8Ax7/xTdgEn0iBmAUZCelNj41OYu4j2JLr0O9NIQO2vOiWUKw9hF69AC8LT11
0DRtThtpZrWeIVIigAeMRQYDQspYjTMtn1tGnKe+JWqgKttR34WNe/ST+pJr5OtJ
9tYeePLGII1pkfdN+RQ3XIQaG7Jo5qW+qn7aMprMDpAZemm7cnqgIsOG+6jVVxv1
DrqOF4z8kU1EE2Cj/UqlfdFiC9ef/fDiUQoJdNRivOjrCYU/YyDyuGFKlF6d1mW1
OdpcVcpu0Ebfb+fp/4bj+qG0uYbKgn38u2qx/zW2mEFbkotLWEYDIc14JYW/u7vw
O/8LAXoZbF/vzvZ4MGqK/Fq0NFuQzytij6AAlqVs+sw7vqsyVtN2kmMXF63CyHWm
quXT03mZX95W3d6ewD2UD9rONFBzbgy5Fh2KrigvQDAhZr8Dan3Q9sD9KKTj+P+w
nuDA7Ca0VaFRejWKrrn4aFUuwvxlKYE2VItHMRGedbrg8bnAKw5OriHOvAbUD5Gc
zqFwVqYNIje6bUoxkFb2+T3aO/MLMMWaux3GvsBhobWTrjSEgA8okSleN/en8pns
t3FPPRDZflLg/5nlEV9hGXP6MIB37/jUXSwrRjXNM1j1KgGzoufznDzihrzUfqcJ
XP88/22MZ2ULxVRCf60dnxRCqfNBc28WdwFn4BqLVJbkCI9At4nN5JCWAs/1ZipB
M6ufOXVdwlh5RpDKGeW05EKxLdFR3LR38EFhKPpFGj0X3RmMiBHM94bIztk6ipIb
QWQDrEJQM7JtI27U0z/RhDq6dOTx2abCE/pCnORa97TN+1/zZKq2ck2ZYzc26L9P
KmpB5KZzIYtdjCUM1eseDaSf6sPfP9A5pm6v3ScIJ3wfmAqktBFCMU35u/P4MBqb
GlpR8J+9rRDpk9XiahaGg3Ezb6/iLXaEA0dr6LO/+Aakqczvd/jaR2soQ/SRYRpq
5LDYlTQfLw9r2m6lPDtt0WormN6az0rLLYtJzYTmnf7ZwZqg3L/Twx/JSsS9qHZ6
HQrVxpcgZSqXTsrsyvgMNdD+9HrjALuJ+NN59xRBYxy9DcVWv9HHTA70zi7mtsfg
b15r5SKdCTR856m0WilWo8q3m6oDanN1Wd5tqNEEBLZtEqAFTDFuKYnQcMhMfbtM
NikpdssvPa7rhhzngj29cdhy9DYPKQ86uoR25gkcRSnsZku1XeqsHuRCtSCEvEVe
P2FR/OCIzseBFU4hP24MtAPJgGBrMaIRmfOdqIRjNMIwtCmf93TpxLfEleeuNvSU
gJr/WfrxvbPjmhSUzrZWVOGs1u5UR+25W6oxnxl5Ix3EoHtGlbpHjygwiSfqO0J8
4yNnwK4Itvw9D4WGgEnSMIari/x+UjGOd/egOA4OmUDK+0N8n5RihNOOW+wZIvwR
MJuKVgJVVHYVzXR1kI4avXFTa8hsgTFEyqXgqLtsO/gifurIpd/TpY9NvCVVDCM7
KMJBPITaNt/uM4HR9NoY2n9hIUMQIuzWfdMazh4VhyggKuMQOSuQaFp3fdHRB6gI
qUjQ8sqydTwaQ5IsFQOQIK+o41cce/55/+80vg6KH1ZG+HJIVk0x5nLVtH5fEAm0
6VbZT71v5iHrORd0U/sgj65zRQ6mEkYGuA5PNovTR6kh1i7NYXckER+MPYXAU4Ds
/1icGU8Fjb4OvhR2RMzi/2S5pkMuO6uu/lzZvEmQGL4LncIxFXeLXotzPrNuKjWK
02w55/8QngcZaB9LkdjJ7A1rwRXGQwWcNLtD/DbofQpHx2V3PDd59SpAoR6LgPVC
MdP7Lj9b8Pdj71kEQKPvrenV6nzPC7PTotPLDCsxDmfVbfHap9+93MYA9UV1Jiiy
Cyf9duviSxC5CNZq9hjAJ0AvJ0r/sev8NqWQhDvo866wHw+Nx20xBAOsiLLAdceX
U34OainU6RSyJZZV2Rn7dnlihBwlPuLTiYRKfH4PNvxP47WpLzRxP8l7wACe/feI
LA2jOcn17Qt6yGIGaJHFiiidI2417h/lZx6h58ot26duXpUBH/NP2iO2+2paYgio
SnhO/ydkiJenZtmIZcpiWiplkXp3QZH4GkCDgYVDhYhOFoZGqhA+Q9nQlX4H/0gI
MCWU5xgRdGMpTAlwKnuPGGkj1Gj9FRSvmu6GImEQO7fHFuVEOB+4a4f6zCKIdAgm
XKs3aSj+MaXe1et0kRKPQrma9uKVrS6QOkhZUDPCurZG6WTEM60E3UbmxjUoYZqb
jZg2MHjxw2GaqKywaovDudnTy3DsT69xa0Jg7oHdGzhe+h88nlLgEzOckvcARA1+
UMmvhq52EULrB37zDEYY2XWFOtTzbl/c9gcX7M7WJP5J6bzYTpYPjr3JGqheGqze
rJ01kJWz5Z31EunRKXodvodeeeb7Qc/YMHdv32Yetv67YJNVdHqLsST7nXrQxAC+
G4KtOzkgZmIFUhlyefg2PyPrTlJY9lMv1AvEFH7R3oCrFrVzueHn2n74dVw1ze3K
F8Gosws/rHANhv9km5qXJb1Ey5VuaG8Bou7hfgJnWwYx/oxCojUB9NRi1igdrjNU
p/9Zu7rspAB8VPR2eebcZrPaYUFoB9RIH9X55V/5txZ1GMmMwodM3uo+XBgsXPdT
yzt7ht53EzkrzSHvkvSZi/qR7GCbtWyBNqGu8iKt/cReQl/YebZuHK9fWLs/q8Hv
/exdZNLoO6I038LQsdboaX+1CFX2Hxny+1sIVV9iuhUBMoRGG4IHg662hVWFFyLb
aHM85bSITKkC6EAZdWOlXqVN46k5iocjPxlNY6N5mgT3GAp/tCzRjhN1awPOtlyi
tn6rcqa+8qB7lzcslBBEsL7xqtAYY0FUO7hF06JqfWcwa6X15qXfWeA/3kl+NA17
M0trBQBwuaoQ4GrTh+GayUhmoAWOc7+byhuEw7GN5Muvi4IVjXGblxtRmIBzSCwM
RgxW5stQFM0WFbtZjrbhJ7/uDt5tw1BBKi5mU/9PTkFi3TNpmW59Wp6yQ+qhCtcP
9b4KBudyBbxjyap6w5JvtsiwHsR3dC3TFYhM1TUPOjF79LdTEYk/GZ8BiTjzgjxK
uKHpudA8Fl6jxYKWfybZxVG4tm9iVaycwdLO7MC3rf/BdL1lkc5oDJzXxjTMazyG
832eHkTkeUmW5xjkrNNhxK/YRx/r5PLOrOuN/pItt0/MWFx16WLpsRujYfy/YtM0
zHK7Bbpmoz9IKqqnCiagrnIN13uqFhuN1L8AJVERx/SoWlxufgDwtAxBzzIBwFIM
WPqyDuamll54zB/lIgIygo8fWd996ECAvTVPzBvYI4j/V2KRyiWFpPRlj9c2lTqP
laHNqFD+o9f1K3lmyWKW80MPeIQcWc8umAyX1gSWMOMnS9kIvaMFNvcsylBnqyX+
xs+F2shVmekP7BWrBoFqKumN0v+i9h9o1z/sj6wCZSwIswFTKmBXxqifhYxK3MG9
qtnLqkv468deqjXgJBc/EZMwAddwDNJnPlNAv4jfqzKSegkazObsRZ23K5St5jkt
56IEDMbnHE8MxtBCqlX1BCMZOMSfExQoLUy53qUXqjX+eRn2oUCpyvcwuDn/Exdh
z+ULU25JIlvkRcY9FntF6ygG7JfASLeu+y9FT0tRznF8YbqXb/gDsiO56rsuWBtA
HP5BEYk2JERY2S0zRJCYzXgQd17BNEjCvKc443Lmy+Zs9inLSGb7k/+E2ZlZ9MbS
IBSlX3HbmWtRWuTbkbgPA/t7cpRxtJFzBuFpek0Gke2rkmhlya1BQqCZvuzYr8OO
1FIhg+7+ejUsdTwqk3HVmMHfnXFnSkg9qIX10L6wSJ5QD0JIHUuu5qfT+3js/10y
83APk55mejcY6cvN4pT4ffI7+CZmNk3qlAnk6xM/TEBRGrYaqT8W7yjJjfD9mGWb
X9dhBT1sMz3i5ZMinTKGdLZ0sCoCx62jCkOgB6OO/kdPexxIJzm7AMOr9hEhwq+4
3pvJNhK0g6y64cOTERiSztimXSKJDJHWVZy3HlEasv9FFsEYUxc0K8k2Y+D6QPqC
ylVDOd0XOPW416U1v5WZDefMyGpwtfMa7TZiwVxznit0prEjZY3YHKmr+Tu1xOZV
9LB13S6Rei9wE1ITcRg0cGFfGFlPCJ/hIY2tmD0h65yXLPz2JQfTvrruHTZYIEQO
lhmwZEfpX+AGZKRu60NR4uEunSfG3EfOVZuqGtqtdXLSDUF/xEfSakgCps2Z2yQp
2IQhYhwGAgUVuWO1wE76tN2LFuR26mKCUi9M1Xw1uun/9IJTzg3Qv8A/ztISXWPG
WDgMl1hECACRMhVE2Ib946bwt45+o7Pn6EEuPixe1wOIoe6dVabU7234Dem0Rnp8
m3OzmGl1m92KtbsQfMLvKpwfZUMOpLoNvrTgK0uNI4xmCqjXUjsa253G1evk+pyc
r6MPyh0wioJFux1faplgUbva0SheQdU1DCyjYvgWBRqR0Br7Jm6OhZkPz9QsFiI8
2Dqo1YTRbWYw4dvKFAAi64lpV+wkO4e2EqAeK1ZwRYcDKfMs6P8KDnfADNWT4nBP
wjAvqb3y2kYBiOU+iCD2/MEg5bVMD3wkSHBDp6ciMg+C8Q1gbQgcNM0f3ggappsD
z6GK/WV63T/nAxzQTEmGBnCBunLKV+oqpmryWigNtEVN9oObbZi9q4OoKlcKfSgr
KxIh7mKNNBuuyfAjEqAF3un538TQ4+obByfwnfGO86ez3tsydXT/ARsqSWrTHA/c
T08PO43qL7tXg2/yi+FLbE46Lblc1qJC5jgO8XDmHWKTS04xC8xLIzmj82NIikpX
ROU386O6xEYAO0xxr/LslZDPPO8R4BZeXQ2knXEibUKv2KLaZfpqCvuxz94M41Ze
OQzQWiEfCpfT5frLGJU+PGBz/gDtSjJ+u+4XwZ6fRHcggM5Bq4wtxfxHp+W+LwXB
/8jmgPgkQlg42jw9ESAZAV7rP2c2M2zCUFkgfNrYEwMLfoFa1cavyjhVG21wR2XH
mzuRlluwyDOlDLQZkc/QUqfAn9nxMyKD7+/pPK+2MzIEA8N5WgYMM8x7g1VvKu2s
vpNXoKIO8G4DuuMMPixkGyiU8eWJ0Kg4D5m87LsOiy2Y3drv50BDXvVx5ONutJ9o
z9MHsDmjKIEdfqzL8Jfufx+pz8/jPC6jw++HSiHP5C0QN/fs1tmS8rbFCsrRwc9B
fRaa53BeN6qAuShdYPh7XljZ9slb1rED1hYeYW7pfmvODQYOIVPdjsCFv8CUmAJ/
2iz0H6AIASO0nq/UqOiEBg3Kf1mxv/U7axpFUKNjb+ykEb27nSeRTyDUxiLTPW9H
lIcqlPQJL7DcgQp9Dd3kMuJc0mkPMLfnhX6n2uU12AHPTPSwadwaLqjIHazNdmcc
KMYdME0EuGim8woFBSR+oW9qboiFsuXOP2bBy7Kx+aOMDAeBRPAQo9SeyMPZvUIk
hmknwg9o/kNDbhyKpF0V6sM7Mu5ViueL1Ey15WCXnIPEqqCzCNFhEct4serM1CFV
khoYnm8Ylna/p4BPcL3ZRh9mfzGUmAmjwZUNwryM4uvrf1UNsZkK3O6BRp2+pbVm
DHHKmcWR7Uo5Fr4c6P49sbSPhehcp03RYM1sqeD3kznlHaE23n7fPT3XyeDwu1E8
QDZhCgtk5wDuUtjoYwAy86As9wGVpiWKwGfpmKDEY+HqOiFZwWW5wbh821FVbeoY
CV4o+pRn8NnOxKmeuuLo+Qyc/BjQdPpyby+A3PfYebtQ7Af//G3jH56vpJJVOgGo
/LyxBPh1U5gqllT511cov+3fGdIZeD+rUdsf/lrvJ/ADOxlfzITZK7YhtEQOF5G9
0j13ZFny4wBtepotDugBhmrVX9ckIngYZFILv4Tq5um2hsmTBe4q9Z52yE/GPbP6
5Gvn7o31QxLqv9juC1t9YKROj//VC+C90nN/vaRTNU6VqwMzGvhdWRAr8mrQvL82
gh6F/BJ29Gbtaz7CoQ28UUhIWqtGB7xrUT7+F0gS8yakmiLt9Vd0vSNMJlxud70X
/f2XePj8wZObbcEexrd1tWkhGNPOq4cz3K4+EOQRUvoHHyzrXIten9vvgswFPItX
CvDgAwvWG4ngtj4ugQ3zmb3QJCV9r5uHLkj32hCtJ4U+UrHoiP3KUC6Mk9xtj2l0
bMxPAgl5phHJIvYKpnaHOGOCXbHtY54za+wkg744GigO2rzkxF4QT4HHmqTsd7sA
+55i094G3xFABk/kQY7u3EA2oe5gYLtb45GJEpLvHfDJO3DMPLC2F2z09izE4JkJ
H5669oSE07McuhaqwHZ6I4TzlY8Zw5RURpCs6cxE4IomD2LipgD5hXs6zPzMbGLP
ojcqv1VsZuVW3H9ytvqS1UQxELOp0/Elk2fXxW16TMHH6LP7sPCEsvrjJ8rfYXPy
YT1UZPU/kn1915ERApYgeNqicg8FR8s6NmNdkGsceCu8h+4fS4rotlNCkDuSOGZg
HhWmCWvC5Fak0vIRIrY7B9KXDGFTlrZJcZq/f62Y77aHy25etOap5z2ZpAfPO+hr
9ADRjsW/jmZCWelYXXMJGBGCHyvbotfwcxhignVyzqD6rwNu5p0yFxEv+Ngw2dr3
j9lj8nk2HSrtdWm51xP99TMmojnvSzQ9d/9aaAdu3nqiagYKml0fAM0bt1j0mDCU
+Mc16FA+tfm2vFZG0wf3fVoIRqePhN8yOeAyfPKHvnaAfxoz/Fqev2t/8X6Zlnnk
iFc1nX8PELvzFednjjWjEOCzhfeaeqQMP0Fdq15772OKpyzoJoQdyFRTniANuVVk
7z6ZQdNmx3sJ0zvziS35InrJPRVu6JUiGBCP9Fm4/3u184mxyIuJa9J5ZPWOlFvU
bTgycge/UdFojj4njl3cZUGMNEyBwpuwvbIKLvy204wgCEnXbGe4BQZ0wMAtuyst
EScnkVCzOnkwS2tYAaGvp4/kfbyCzlOKKjOAMx2hR/xxaC0Yozdt68mgknD7IZwD
aVelYD/TnPWdChpzDqIY1MvngPymV5tOFdQbpAv8upkIb/SKuyRlCDu8Vi5a8zzI
Q/m48EQSUu6IAMNPTweSYwgqzwdcZ9SfPWNLs9bnNMPv/iyK2BffaOJ4zuZLgh+g
HbSgwj/JyVCasMFzpiKVtnCCJx4wF4clcgVPlfpksTtZl0LL6qcHsB195PUPjND7
RKA1rDcWf9hCxLfQWyVHuC8Pr+uKFJqDFuOuNgPwLxMUJiHG+tWO818Fc3d7pTWa
cX1jV67iLUWKqAmWTxUVUrWTNOMplYx3HUux3HFDcvccCRyALwKVZzZj0+agU1U/
5roEaKNVGJlei+cb2IhdgMfNn2WqgMfME4JbN3rdp7C7cVEi+47BBFA5xUr2WaK5
fCcZRXxsTl1wKyP3x4t0duFbAG6SdqMJPKCAHMh8l2k2hy6XUJyYT9VqgNzh/OSz
fzOPn781V4qfnXk3CupTleGyBtEliWnSx8nz8OuZOzqLdP3ij0m/cpODT9yCeoET
2KH/yvciBuXk0Q0MdX27Q0rx6FVqOqYeGqCfvPOwFJsazP2F62UtUQ1wlVsM7wrz
LGZii3qUxLIX+rQK7b1U5wg66LT93aJZ4Slq8CewCHjzcPnLsgvhimyekr24Yo6J
5LlVeEhR3afDh6sfFK2jf5HiGYrAKYONRzSA1SKiL1NMnoRVhsJ2H/9mGPGU43tb
wbKK1TxO+df2Ka7S1HWNyGdWQ/G3uOhQx3akh+hlCJA/6a/PKI6c2xblMXgw+axM
+dfxMJxQM2qu4uf6vcghNCMcl2sJ6NwTL9SPvH2eoEQX7hhlmzFS3lsA542U5CJr
Ww5NBWFh6V0tpbQIcmWmqyniEth1c7QGGT0UtsWW2ooWwIqfsSjGUyYMKOE1rLNa
V5Zv6v9uCg5STv1Fsr3e9NvVhRNnhboJNSCON8hwkB7BFg2nmIzdFEQU413KKGWC
kz8RFGISIPk37SDG98ZuhTe/1LkCZG9QD0bqJG9Up1vp5W7Sd9myQd+Rzz4mFfII
gclHYNTOUmuCiShizg7xixnYbV2xlip99tSeiHH2v67A3UUF18Se75D3y3eCpQpu
Lep/p6xv9CxpBi5ahg1cBo+AqpPfIF8ur7ervJ5BBzpmmBaRMYorJrxme6molmbU
gOw6hX7kXNdeldD+40KZSTXrpXU/h7q8pELFLZVw5FPaZIRENs3m3MRAI50ev+fR
uxXvoimuH727xxhiGZaf46lKyz9/i4NzqLtKwcLR58XIGrcxnHolYHel4TddCgCt
0Uh2c/iiSMizMhI9x733K9o+4w5kYDP7WjfRwQGIF0wJa4wRurC8du6H02x5Rg6E
IREQDz6Q0yCwWWyHO2ht4zfIBk17znuMxi1oo5lB97HwyDwD8aSv5zJsY89vXTDc
+vf9hb5zv6y6oh1LC06RdS9NpVOrMF3Kt4GHKuILfr6xRbwwa3xJBig4vzx5G25K
dftO8oAfH9MCM86+PvY58i+mZM9XOdTK2oyNqLHm7TVMZsCXoU5R9sWN0LOKO3Bx
gZusFU9AWUTX1TOp+oUHKrPRfCqKlqrFDt6+U9Fqd0bZu6tTZTL+TWVDaGiId6oV
gBlBpZ0ZTkcr3XRM/KsVMIgIkd5t8YsrTGtch5Q+MSbbj+D5nqz8NlS+phpZ6zgW
Dq1M6S8SRbvJwd6LhLrstpnKA9nbx66e5hLOBoXXlx+7yG17CaA0I4niWTup0b17
aeoz+sRFQQsw0G3auPb4luuRIbhdr+x7zEje4KuLTknq+3599hoo44QMfwVX4O/7
cB6DPDrCfweQSZxxBCNF0NlWmWAl15IH9XZSz3I3LQaA8/Lqez3VwTGOlq28u9f5
SQ0knMp9xB3vNA7RJqfNCxU5GL7dh6/53ONSk6WF9pCAixWp+9NRh0fRO5qtcwnP
KwqTmv6Fgjikji1VL0luchFIwmrML5sntK5ZHMa1/i6p5mdkbRCGFLfRFC5w9WTl
SzkrhYsHExuZLnrLQ+yKmvto5XuF8Y+3mnWtnpD8EVU/tpX7z01CQ6YVwv8cYZyA
P/qTx0g1AUyrexgVAvrjmDC867mlG+/lCdsrhCoNp5UrWDMrb7G4i5JYQy9BmsvD
JbtKey1PwpJLm8fuaNZY7z4Oga2xaxWa3DY7VRPf13tlVdqYTfj6yHwY0yH0Ttaw
tsrtZq5htUqTIV8t6ZAk4tyvNRD9eJOgCI29bl5yXs/vFtNBhjG0RyFldl/KKgIF
FgpuKSxTsSQMhdWP1bMPsoWqpS7hFR+uXbgAecGSZvvfMTAv9eg+x9mEViW8eBVe
vSOaOYWku+1RH6H8GYvyjhas6wKI1GKy3k2x5lek5L1kK5nP5YxzuASZ8kZWx+cA
qD2+G9sdKDF5zrTd2YNCELdWsZW92mXLfvP5MTvhsydfhV3rmRr2Ojct6kqDx6by
8I8R0sjo5EMj9E/2RnVOSEP0GfcX5EvA4EL0C02zZxmEobIL2NeSzQVRJaB9Jyuu
Nexc9uY1GgcX55I412JGZGAiUd2E2mZ0GBWUMYcNEqmOXIVmj/JL+NNPTbCK+/qB
2aXq0rBe2RC+5WjL8puQZxS5wwAyGhwedE95KuTR6UJ5yfTTsfBnNvA+0OZce2yX
glZU8O6R35+CbJWHoHvJB0s1TncadyP5DrydHAficAPzhZ2y1IUOHilOuB2aIyjW
X+kbsnglGBwT2HZ/by+XwvOuipmsPnyihSdFYW/Q3I+FEupCAceeGzhrixVDr7xX
aCd83x+PgZdPVRn4dXw7ziFvuyNJMM5o7plBTqnxmZOxIzNES6zL5AxaVDH2SFP9
h4t0K11h8FN4yEBhxDeyPQ4+pvcdBCkT17yy+b57I9SXLUy76lYbpdpXJ6AVLUWY
tZDtyQlrm6MIxZhv97anPAF64vKhKz9hSo5vSxpuhnjPlkwMDnCNxr5I98mlvL7J
JKjwp0emCnRwODF0EEj1+1zApGPTdGgWQ5vJgEdWOzpe40327DdGNjvKry0+kQWP
Pgu9p0HWbfp/2jsdCPytyeWj+kmzZYj0euHh0xL4hbWzPRvCW4BvWP9LgoTuY7B4
dVtbf8OJUg8KlIXOnPPoic33N1QcsAyh6bkQaEElIlEBFmk1T8KwKF3qhu5IEv0S
qP3FTAw58r5cpdRN3lt2ccZqaLAxH5z/I3xkStOtQ3WTEm8UhBGZaGJtDNsZ9Bxx
Wo1RsB02JAoyLS8+7AZ3Ms0l7Dmz4dyJ1UbzlSUzN7tnHAaUKDkOdnOAB+QY51my
LSN8b3xP2q/hyRb1cqqkqBWTMEbFZkbYXAKF60tk0LqH53G9O77ck8OfiPc473qx
7SAPMBVAq+M99nHQu//lo5Y96B+yRzzJEPe7M/cWXrcrdb/uAAfW2mOoPsk9DbAG
GjI91Hf+/pSzUFR7JcMm5LbmPcfE5SFaOh/G0RbVpxIW+6GZV8OVvrrbz+v9JhM4
hUAUNmiap6lqSlNciilNl9bEkQVsjt33qz0JIgsxJFbbIOpBJdPBh6NeeVGUImXH
R0IRORWyTM+vFPcfBI+5qiGy0fHpsYtK0EqgA6mvmVx8LD/l5GE+3la2XLEh6VBm
bOqbAwSizEIDWAzwMW9K76EqNmfEVN3hfZXLd9Mb86e4jMuSMk1cdU83DueuObMG
sbH0Eit3QDxd5ZmxKLUHVdSKOOQTIezIEM0/BWa9QY7o6Md/w2e/cYqMHRY9QWhy
+p5e8E3Ob/G7ivTZAetGqwN+L3Vx4BWKN3w+QwzPPgIo2LE2nekJmBD0SxnFfe9B
T1G0y6pYtyfF7Tuk0MC24GLgMMrwtOB77o4fd3HvDOJXTBLZqLQeuEwOVKmOJnwg
RyVWEv40s/2Ov+13qZKnHCKvid38/Lu9+1OOzTjDGhpLZfReK7WpVro9qDxVMJHw
skTeiMsi76LdVL7TondU41gR/+3EtF8RhjHC/B0lhKNorUXyowMsgwu4fe33aLcX
mvQxMZI9SbYGgnDX1qh7UrawKY+ooSsYQLslnputzBF7ebJR113QJTJiGmJGy76N
ZpdFEL52Z6YikYPm/cadBeKLHUx9EwcEFXQeLUXwJ6FRxI7hMu9mLPwuZ77qurdO
prGzerbiZTFzdh+21YI2Vw41zX1nnV93sJcYDjG7ld0D+Ssjq6PnSJxj7E5lE5h3
ixuSeHyvaPUGnHxnSo0FWUHRUhoIuTCNdPJ1OYA9kU1MxxrZEeH/WxEky3UjRAf/
84cEjDerk+kTtAIh3IdQwsXGp0bbuIAfKwqjTcjOOSsseKrVTwju6G0RY+Z7QGnl
mkeG39kONobuOz8HT0+j5uBLB5dEJGlSFpMJmNYmECveF91LpxusuBGUf/AtNRSQ
11I+j+bw6X2AcR9kiFk15z8M60zj8pPFKLp9DjsTnP5Yltyf2IwKy6tkjpUYXm1R
ckpwUyj8YK37I9umDq+rBdAnUb6Y86PZWwQLUMikzJFDkxKB+Ip9pil/xxrwPhKy
Fn5jmQK0TPWmYFJGig+0eILSZFB/SbTP41E5af9SMWadAdYjqKu4bn3ylvP7TjXY
FqlofbwbRSN+xWYpb5CjfHX0EFcx+F4hFp0u6VJZ3ha8R+mXM2tZ7FcIsOyzgQ4U
ykAvzMynUzUyJ9wtbPEXlH/hl78g7u1/Cb6Wj/wkpTFXHBHBoChkFV+NCR1sMjo5
xCXlgf9pydbSv7BJ7flThGQdQQKvqlcEh66UKJVu8AcKMmICeYCYnq4pQgKG2hMU
/FVEuPFM7+9EpZ8mplyV10ZZyQKAvc8MROFE8mTKZacVj3jqcdMaoFUL5SF6rPZW
ub+Zz/XTVO+kVf4wxv2bjkS6pk+EANDVWPLRyagXOE/OTOWMLpfQQlyjumSzRYyr
F2NlgVrrxstzGhgbBjy+VexCl9glDVfvEfHufpeieg6aaG3wBp5o5CnBfIppC7mv
8ye6q2wnqea3og2BZiOjA36EHK0B380sxHQhxLF45WvHPgA/uFjDr3wp6m8fxLE5
Mg6Kwp21hfYS1/PDwHKDA5EOKB0OaDpZ/6Du3H2hE0r3kN6+rBXWt/VsHsp2/RSa
hhQ5wHAl/DX0TYhOuBc6vDfm11Ue5uy3VHsygd7dQC02yKHNnnLzDNk+PfH/G+IJ
T6xhnGXZO9aaFfPzi+M3BmttPoUuyoGrzQmiimNNulzrjK3J52yNMY9Z0y+A5V7Z
FiL1Qex9e7mDKPOOhe7Uc0S2Tgx37SVUWjlpc6uG0YpeVlJwLPkcTwtBzHeYI3vl
4ruyjdhLtjNEmmM6lALXUh06nh3lPDFZbiGw2TM2W8UiimD+Ng3mzU4p3oq3sEGF
ceFX+SY1iec2c4yVhB60NOUzPTkzTcLUmyqpOyv+npLT38u31JeBuIAo/dU0cXBi
ZRItABego9pFuPLwDQnLexHyUlUQodnpgz9vhInsBTq/w+dbMFRQvvjbGYVTJkwq
y38MVnImN3+IGALK6fl8X3VBicNlJyIDBumUIDC2Fyscdj6gdLJ1zS0qqgO44VOS
VrBmfYHXIT2fXb/yi4ZfgUkg9wXiB3f3++lv3OCma3Q4Fh3rRrP9UrEvswOiTQbt
Ms0EFAuQiucEs6qVuF0CXXmSBsLO1cgd9y+fV1rhQWX80LHMhxhsN1/oylNbNPXZ
xbhnL35IbwB4cQTBcRqC2jWio9zYGR9v9k50/tKP/wYRTxufTGkQruYbqjce3JMi
/600c1k7bQXl+VErvtC9/nQNuY4VDT0Q1TabUvb/HDZOtUdLmsxxFW6yditlBYnI
FrZUzcnj18+IBDM60mprQoXzxctpOg6WZ4b5YNshb98JHFRbk5OMklJ3mkY2kRC3
r+9T5AGcOh3E0cO0UA3UDjl8MXZ+6Ig7OgYyUSuV+qYbpSNj6WDe+nyvMFaauFWH
pcwZScJncz8/FIi+ybFnWRO/ws5roD7euNtrPypEa1Y6HWejBq1hmw6jrXMkIpGU
UN0Q43zxaeGYWVmY/i4sQlBjGLHLdkZUKWaoLNWSIFuPsQMbnluLdz3F9Lez+2md
/svReiwS8BhsZIpoNVGYv7ez8J3aNGPgD7niEIfxITs1uiKlgBS7N+iiKbp0SsGb
GbAdIfTdAmsbei5JQs/IVTZuDp1zOB1mZ/ZZPvHmNqNzN6Ewd4OhiYPfJD+HVh1m
qnuYsEP3nnDqt2kRcuPJCksCuWKmhKyX3+9dUHyGBVIvTJ4aLG68eOEV4kOtFBUA
VT9fyasF4v+Q41E3YYw36u0m29BDPUhkTPHgvrTFkQAuHwL05+f9AxarTHzR4X2a
iksnWQ1I1zRFFq69Xa58EV0TRjlaQpwPqXXUbQEbpG2oJHPuPS2gbazLarDMXeGe
5xe0660dAg9Tw9Za3ijTnp96nuF18Vzf1nG2DteMxri4UWW9CJnnbP8ZVY1TnROv
gsfDt1wX3hqKubE4B5F6hVZFDPO1oEr2yYwY6ZRPkCCc1DIFxPHgnd0sk9b3Goy+
uwAojJUDcwyGnJ5GH6hpBjE3ptHzYP2QyB9FEZI0Eoa0KaiWgz4yrLWKb2nhsVJa
aBStEKDui/haRkJcoj5Sgehof6RW6n/Oiy1A5GiYP+b3Z2AjXP/TOxq3A+u2W1eh
LLgbrmuFj8fA3knogJ588CA24JH3V9bMnhy66JZERbgXn/iQrROMXfTTbW8jFyXX
bY+s35Qfkud3TVo/bPRAaX56dq/HZnDb4lp4BoVZQMFgSevJSOY1WFzKvQCijhFJ
ecluADfmaDC0XPQvfMCrGQ899/SIZzE1RZN+eSuS9LNNhX/3b95SePSUILmCQyxH
zME6A+5N4kr5p5OuP3JEBdg5PuP1bQG1ZaOIBZK10MN8wYjQ4b56KEvxhepuC1w+
ash+Vb+bo2WN9JEGKS+uuHNV6MMH2WjdLoN1uT16+Kdfps2iGIP677KgwQAst7+N
rFHb7t7nAzhaUMuOe76lEd7TmhGCgUSh/ZVDZjKkOXytgq5h8TOtOR3+jyOwwdCd
THw+rJDDlf7MDDXLnAnEp/Mw+/dCYr0tGSAtITBfFLhQOW2jui3B1GPU3mdRDfiJ
JARGo67g438b+b/TbvtWB3VK62+sUyIbh4f7TCzwwhy8CU7e/VqLE719Y2/ZpSQk
cJuSS4XAuR1zy5RDoWnbYSrtuBxSLPIgRAVP3tkszYbkNF91rMi39t/g5VfleGrj
DKhvbGJIWD3d8R7hMZruyr+dSs56vCEEmdLBAJOXuKH7TNB3j939+nQ59nupOlel
wEnkI/uXSS6WdQOlIWD7BORukXwHrQculQ4vE2R3m2NJGEOQFrqZrDRAuCPGgC3W
6MQzHx6ryHKeQk39VEtsyKkHWluAR7Qab24vqwOXAS6ZvE/SfCvwVPvz/+HVyF+r
FaDs21hvDwQjCxbUnWi0zaZqdjRtC1YJ96eFpsMrC/gnjADOFm01l4Cdu0BlZ8Tk
sF56a+ZRNmtv3ILwLeLZv7Vz9NjgFeemlMkFlWY+apDE47NLNJ4cJTI62UN31dN+
BjmxLIHO4pxvkMfEhWXf79HU5JWZkhbt0yBJsl3dQJV6cSdVgBk3tgqAl20t1PXH
BfVhokdw3e3plt8qnRL27RIRuLjRsd2NZNYjkhPXC4u9iTPqaH5acjqR9a2keCJU
f9l5OwVk26ZGemUfTWpxO4sKlM1eJPbtuNU/J7su0akB4yWvKXUnd0Ztklx1vLXX
lsEOJeZvvx8Zi49M1r1M27HIJ3rJ61Nd0PGaTBI9qDxD4YUlLpZAJM1DrJBIbhCf
Ra+gvktsFJLxuzuA+dHB/FYPZxRZZ2803fCe4DQo4T3Ptel168wDR+iDOuhzsoAV
I5eY7KChwHY6DYbkgfC/ZTPboLnSy8HJcgjjYlPEPSSZjCjc9P+XhfDVmWHXIRxr
aitSrCx2Hkq6dotlb1WzPVDdQFbF/7+d3hNbqDAiAl18fBoPIpbfouw5NvGVexrI
IcTkEwS1jVLYG6ERuCFTzvQPS5oSbm8SoZN3S9rTatiGe43GFUUczg9GiIBOkS2q
87eBB/M4S8LphJZsN1gLSkkv+ztgsuMh3pd6FJ62GrLxH4kPp2vApZZDmHPOaG8p
3epSTJ+iIF+ivxA1Ra3RPvT/zBdEIWc3VqPGPJqqSh2zviSIks1c8N/Xb+QpEEL5
66Sw+PJbg6yXsZM8FqVL5GX83e8CQw23mqPe7kxLqVLofEkYSuPTxqjhf/pOhXex
gv2IYZGHSP94gCKcBtGJUssAct1C/r6aIDWfUxSpeF0vrt5M5PaELJMW9D1I3yuN
GBbuASMnUUkccecniRI8WFTmHGEMnQ+eRv4U5udQhRSSudu9MubdJZ0w0yPAhniM
0yD8quGGLNHuEV3lPO38ghxf3M5kUrboVVOsRRgDLoT0m74BZrrKDqaXkZYpsyJL
vPBd4q7IfdJr6OV0zwRpJncI4Q0lR1cmgv3xm8hbxSxCc958dw4q6as1dIGDRrOU
sNjiZw+CgOEEA5+5bBvpc3AtdAnjVtbRbXRON6X3nHhWFCF5wBwDpucO/EmQ8yli
Hl+wzjkaDlwoK0O38hAa30XeD3Fpx5C+WRONhC1GXDC9JfWhtzeKwm2C5iYZkBJ3
UNZJsmtGdsW4+dCdyR0TuxDny5GgHtGhq/EjxyOioEBbHHV9yEiq/osBFo1JwzqI
68/rmxvgcHNRtK98Voc77VUvwqQ/8fDQdheG95tIp+4PD5IqaNY8H7BWLhrDL0wJ
CLXpaYz5ZPxeIlFZdY5p/NDUaBXsukhcTZmFLS7qVtN/3TVZnSHaei8livDswe8S
RbiEMR+w29EdC0DZyfhluB1D2ctW8RFj5OMqMWRiyaIgwojCsGL8/K2jNjORXUf7
pDL38NWrcRVUWmUTIiTHk/ZJGGceenOhghy0ixVzwlA0Burf7YwoH4OMYdi7g6Fl
cC077/J/J12YrrnOeCSp5XiTJrxm+OIrrtvaEgB5AYSPtAjaDOjR+4KPZp8cWvMR
733j3sw9Zq8Z9WKSD4lvgiz7HDV7uE/cdejAHYXKoFd+gSA7RyJjbToH/WEQnE/V
zfhvgDP57ubTsgH2jjChdg+ZjqFGWk9bbxhoCfKF+7xk1Sdq0QFndTd7dXpptUo4
kcaA35tS8ImGW09kzKanJo1KXZMGw58uUpEAg8RECNnCkGWfBq3fGd4pF7C1F7+v
pa9QLxy7DxbjCXew/pJafTpd6HnxojUP51rvDaVlOhk+QMCErprNW7DC0xpvS9fy
EaeCuySzeIxs+YBnxrW5ammjRKTlc0HJ/pY1JMfBrEPgeUJivB4wWpcklE4zzpeO
b1osYFaazcV3cR0m+Ahec+BftWZ6DK3cr8wmeI8VOpgr4CQlONmnwDdkPby1pTMh
cNU7sy+c4B7BKT1DQ2yGQCQAwFyV7qsqDU8KROt0vECi+mDQpLSL2ihAVeksWJ7D
7EXWcnHEY2MFDf1PR8WN3zZtWKqn7Gbh/WNnmJNzht1xK7GwIPJNUoqNP51n/kr2
9c5bc0HbJcc4aqm6wzr1duoN6q+8E/nUAI9XPleOpphxfhUlFyZRkN1QKCj54GjS
EjLpQNopQdCYhNxZ09bW1Vj08U5lW6Or3fm1C7S+V1BqRcevhSURKNMemorud4eL
MGfQJRjiJRkTyCp4MQxCcthSo38zv6ltYGOzXqvWsaF//dixpBV8jQsnsC+mCxfE
MuVPoA1Gq0ZODoUrwdmKQI1EwjxRQ3wNOOpBewrxYZMiUzPnx1+M8L3hw3akLCNZ
hRY5xD0mfeh2jTaq4Wj33MUxHo3UJUQnCP6EcLHZ/jEGrlg/rkNPq4gUB+mmuar6
wSe7c14mQIdbmLJ4fH4xoXBhUK4btJiZfZXtDgC7OTQpn7JqDQIAa8qGq14l2nrl
Hc8TzDNW5OFXMOyRgyrJX8vAk8NTJtkBmDLlkAfmmqTS0tewlaDqfU/IikQKNfq2
LPSbYskw4N0Xi7BtaxOiZ1EOwarJDPoW7lajIqdSuVfplt2UibTrqab9ihOnLG5d
ZSPmHdeuz8P7U49yOZIHwkwaELsPKauBWju5dqiM48G7G6Acn9r7KPJ6MJ8xVuWz
6FMT8adnbUl78iNmkTiKaI+j851TYjsWYIhS8WaAFQz7vFDTxhlj5VhwUuhoZSrk
3Qp1781VcKS91O2aq16airoEjS3lBmU+c1yeU3io01h19p2n25UZorcE5sydfcWn
Mphs2Ywm4WMNTn/6PC3Mp29eeafwS61f3ofIsyhPn8vxqeoKnHhnNPNoYPKfRY9R
eIuhoWdHHa8u/DBN3xjw3ZE3dgZ14hjMxqFOrTjPJHqnr/zl/XAZbR5M/l2aeIFz
726Z+szpuOefhjVpWFh/2skvKAKHtk9TBf1pzgSUVtxO94d2l6KQD3q0RL8V9XCI
55GBsTxzXbZ01j4M5ZBIyFz8KI2f94rfZxjb/QzQvWt0ZmLICVfUTIf/FwMTUp2k
vq7Gq4CfAdIeqP/v39wW6NoME4nMJXmtGmFkNnB6JLLqowOKVzATyjeZwBUXQkIg
GA+2zQpI6Yh2f4GJh6jjJhz/7AtqFVzU5qKSf+UYmmvCU1RMgh216R1qesQ7c2oL
Z7CaEeODB7J9IP69yuKmawTpIn+W32RdnPMkydfgAinKurkjdXliV3yGXtUScdX/
p988aev630CFsqFEnMDQnRBcSRpGUgX8Fm4uEdfsPS9L9KIoNIKND+DXKvLoXdNA
G8TJ3FSlG2cpUlveVZLS9uvd1yMVLUZlnpQabhO+n97BA4fgzphJpA2Pagj/23JI
qXLcwM0eThqFR/wnQT+F238ePv9yTm7kD4EZYh2pgkfmTFWXQZuffAGy/sR0KcLg
ZGo2yAcNdUmZXlyLR+8WOOPV8bP+24ZB/s51jFsvO6jBYBWPRSW0CHyBA7q5JRAt
IA9kgM/W9LEzlr0bTkQu1RFSVEgAr+6taEjd9zDrjzLPrhOUVdrKTC7hTOMkfvCk
aWf6/mw6HH0gv6/3kwR0kiQEOt2wV81CleND2hojp+VXMZsJUQb759WeID4Yjrd0
5XmAToU5rjgwogQL/gYS77TbwIsFbp/BZYopTlOgbzIilKR29nn0NuNSV9LXDXQN
kN4oyp4fF5nXAt1FvGCn2ku9YIGvDJIXKWUYUYl3CVueUYf6tfxKwW7T571lcYkQ
abL1dXbn1XBdpHKcAqMbaHBFB7H+Z6NqxH4CtNBZTys1UvH2jVx5Px2moyR7JZHp
jMe3yC5yZU12ewFGwbBs0Ylcm9eHsk+3rMdxUJdNIlYTIexCosixZWLqJjTsNYVk
/xsO57/zXVEqh/6JJ0movdryzJupu7jNFPhy6Q/+sQMjqEsotC7pptb7c/TzRw+c
Yin2B+5a0aorsfRXgePfNjkXFdS8PdvHmZdkvUTpYeQXdCe+DGmEQP69V2ISg/BQ
NRx7mwJ9HZGz/GT6sbD+mHo934WkX9waCXCqEoDkr1R2eA2JKeo0jl46mez1T9RX
uHs/B02hWkpwqVAlqccAWdLbwUlNWFAbFKE7AdrPKuyzmRpsEnDomsMn+5hGEkBD
IXXeB69EphuzWHYcKzFc4usdyaSRNEHCmv+NMK/AklWkCYgq0V6EgvlcEH3idUE5
l2xn3e1QSmMJ/7k+++2o7kBa2wcj2GQ4u0cOZ4OUy5PK3CNnPgnQt01tUv9ckxTA
O27D2debNlQpHp9H/HmCHHi+ufr5m6odYHO1ySzEFBUx3hefo3WCCkCWDZb1rkYQ
RUl9+OPejA/LX0jNK3mDebGLu0VWuteNSMo/8TMSrWLhEdgBukhGGP58p0+oimw0
sWbeJwZjtdcL/V6Xq8OZi6eEQ5cgK7vUmFy/jCfaYsAu7QyJUI0HPmY6vbyqaO5X
lED7qFnFKW1aK/ZaIn1E+B2KWLoxoGrtAYtH+hU6KHPL8HhlrSg19I5/5SvfjscX
hPyvX57FZWP/iA8HWzFHRG4TWXwK+JNMi/ChH9XLq6BCpKLEa5WYLoudh87OEPqJ
WlPnPyZ6n7tUYIusTkT8j0beKkTTn3kLvvaXec3aLsqUGQTE4y47Y0x9vGEx7PLe
zItUmRMdOufUGo7wDYjprWi324Rvh7KnEfZLHZ3baDMcVVDI0gZ1bqtZteJiKulv
K9VmYxOusJSNiilV7jjAyFiZQC+ctpG1dwGXEqIOrhpTB9kBWpZ7g4cyk6En08Q6
Vus+Evbdo3QV7XR8VqWnw3noYtVsZOYjI6s0xD6x16CUa0KmizzajHaYiYeyWcrd
eQ4sH4cDgmnXRu22ZpEIizOpBmUcWQZwD3J7CTp2/r9pFUow6Rmg527jcROijZ95
JbCYTXH4d7J0fZYQyr2XmYhPFYdrK6SgepWowShBmaZMdJxTGdzxdDyOjF0Yz0pn
9YsL9I8mu7mrAxqZxKiHb6YvKGqBMWTNuNAKj6COjAaWQQ2oD5B9VEBGRa3sK7CA
DbqR6Pg1wv8xWwoX/V6n/Qx9GXK+USdq+5uLF9MqRmfpF9KUrXJiUIam3avhzths
CoZhFuOAy3RF64AmJfhflTL+igkjX6+g0fHmOCCFV/0HKmyAnb10mhzHUG3jTUYq
0dhVLY7gII9nRKICNg62tWxAxbkWCQ5Icy0Kur1ab8CqVctm0HMcuTMhk5L4OllV
az1Skdd9mWNHMcsFJ/uQLqlPVF5jtf2EvX9tLRKZdviP6XTruaGrgEnTEaLwPFHQ
trH5Q/V9N8W5lB9/jQTlqWRPrJNlyonlEHsh+2FiWYz2lf/kevwjBcMEuq825v8Y
QD9DUf9ynVi8JrnIbirKMViln2eYkWMh5k7+IBQee/40X7d90ENIcsHwBW4pXxTO
iuPZvY+mJEUqP//MGJU43njgnuq0OIK4h5MDapaVE/NVQB9x8p5SikL5wBpJ5ymn
6mHG+OwvynagHerwy8HWS/ZrWeaJP/S+9KrtiXr5vYDvicyPXQ555pp6ICvYkdR/
vhPFiXhUpKoWfgfkaRhMy5J0kMlo8HrGlw4XKjcxQ/g1y4Ms/coFqsNXnRe1UWSV
FL60uPvAOU33LFw7TXsB8PjeYPxQfXCrXtFSJjPwwrlwgeiBBZsYhvzbmwS9noa6
7OvQja+LD/MDHQ/iv5IeI8ftB9CF41Cpxr4b8MeW01WdJ6QHSqJvh0tB72XJ1In+
nqnjrSDtQBV5lQPXaovfPBByibEm1PTchvyJZG9LLD0HGPyH48R5/P15SGwHaDWM
KOZQySg3+d2ay37eTvsFojZuyexDXNfK/FDWqiu/EqkevxTM9DEeeYIrgJGVx/JW
apUe1eLe8FWJo3m43MY4R0o9NGXpcX7d4yzU1gFpRpDof4I4wwPcx/ySo0NUjPVn
gNlq/p5De1iDhZWKbYhu5hC0X/4FAlyaSL+kQmJN5bvu7bxqG9+mdeataNR90Nty
kvKe4YjUXJT6RZ8W4u5Rhz88MS3puCL3a8D/SjgccNQU0j3OLhIV6N8aRLoKpA8T
Nrvr2FrMvV3MJsJVv4wc9hrpUBRf1Wj0wP+GQgn5Y3hVEi1MMsN3vFksjxmcnH4K
/ydbHwcuZE4QSwM4v9qOSn3uBDQOOazKMFq0auuRMqrKfM2z6/9rN9uqIGtdKOvS
2r8YFmnyAQf54tpUIJeZu18cfVEbzlMO9E2ARN0RS5hKauDtfpdRF1tICjG00gxq
n7hXo2Otk1QNcIX1PPg4QlqiuD2yu3YHwCqQXfmuBFgVSa8KSrR+6qRumstlEct4
1K3uSgzRxFcvLIZ3+zvvXRts6o5P04wuhyFL+MnqZ4/xahXN13ymzqqRQzBp/wuu
AEXKC5KAgO25ktJ+Z/luUiLUxbfyAAslS8oqC5nBAIf5zY6emjjigd8HlBou5wzN
noQcjITrPfP4aBx1ap3KeOvNfd6hxMe+3Zi00PpYrUj2uSbk4xa6RNEIpN4oBhss
rbYFrQ6JZ9RYhup2m+sXBIHAB9fpHauLM+yMzRPCwx3DQLLUXPdqgthl2k3WYw8d
lnZRtSjURBtiPavZp9nn2wQVO+9b15DY0RJwapw66u8Hxdl4AA1OxRPZB1up5Kbj
6MwRSWLLRDZz4bcWDP/lI/isHZE6CdOXmjHHbAQPOENTLRf70GzxVvGHNBpe+HhH
Il31JFo9G8tjHxsyiwIweLZPybo7bKQekS5wQL4vgo1rGT2/c9zB2nQ0wAk1Ql1N
BIm/cOi2v9qdkUNEnB346n66mT7jxjVfWT9XBZEiuRecl03sQUmSoikmtcsjKZTZ
HYXAejC/6HsRf114+YnHqW0IpotJS7RvKb+U8KYuj6azIsp4SFxihlfeZ2zm9dg6
f9dwOY4rPpbwjr69G7MxltBMZNA4nO4nDMqXrtjvQhsd73M6cTfCqqwxrjbEbE3z
wAvFYsUaVwZ749r534YmXUgOukKA9XOboLPUaTnm7chVS3ldGYKt4pauCHXW/cxQ
oox9qKTz3roFNM6oLNuujztQ89wPhX/gkD3zaEtqyqEVsUGqkS9eOUHTLAK3XGw3
U6TXBt/wQSeOssq8xlrf/3xKRJF0/nDFOCuTOWGuabq8EBqtZs2mZfCEmK5fKPib
tUmn4dwT13CFPUTlDxlX31jowRI1HLLUpGtgje5+7jwNzW/F6NYuzMj2AjPOCH6V
rX6ffXGEKM6n4fVdz+DAF8UzCz5/i98jHcfQV9us/ZnA02RSIZVGS/x4ZnSk4z6M
aCG8SnbSp3I0NMcndyMBFh9waiQXaX7QVqwrkDNSk7pRR1oae/uFBBeUiKcPoAUy
v1V8/NyP/QWByPwskfVPYxt8sLqayocIHifAF64x4YkwMsV4+r61dcjGfPFGmH5d
tr/WlrxLAh7/s4iBgNsbyB/fBbsKzYIJVPyG3JDLA8qe+n7N/inqRDLfMrMbDC0k
Ode3nIpen/wmd4KOxV/+rpGK8Nd9+AKpodHNJCs6pnUo+owD5kCUmoRneuo7dbs9
llFNt1h0DcSEjb5iVv9EFfIByEVxQlvWw9gap0ZkFL2UXqC6jQQlm6l0KxtjNGh4
GqyD/Z0L7E6t1Ax9zYlJw8x15C0L4a21IXDHSLE2kXRdihn5P+9QtV4Etg1yJB3C
c7Kov6BGCG9suvd+acuHv6MIPma/7CrhN6nYTWajFgmIgmSCN5FPjYFm6I/CSWuk
pFDA0hK60HbdaLy/tC22apoOXMzhmC3ZoxjM1teWSs7coZIFJn2iPlgOn4Vl8D/D
f+ipOZYH+L1wJl2gFWIfV574fznm1iUIN09Hix63H5P1Z5vzvyqtwhtzZ2LtksOS
ZzKJMfOh2KqbWoA74YcMJb+FgFAi1ml1x5HTy6qKfAYiPhsPdJCBCBQwCf2eLlO2
0iu0Ko0s3+lKvfk239jl5m7X9ss2odIuyOp49xuLryXXgMteqzwToO2ltf0Yqvw2
qwKWyMxpUvnbGSCNaNunwv82Q2LazHzw/O5yZr51R8t9KKV5hvhkZsgfbwdxVXS0
mL3DcB/XlbU8vORZtjahxSGM4Lb4ZVJr6lgCLenhaofZIDM+/xyYHDjVMqle3yYs
ZFTDxNw3srN5AStSZHQST/h+T6x189z15fnRmVsVBgl9xSPxjmoFIPI2OVeQWxKd
h/0sTGUXFi0AcnngYRZoZmEZUZjefsVhFHQfNOPkn06kzKB3dRxv6y6AItpounQS
qqX13znb5LvERHg9fPYBVtG31+WoUd1P77SfvmZythCIQXxV/kgg8U3E3qax1ILp
+dOF3pHzQUn2TpfIlYj8K9hu0EMs7z5S8nhiwB4Cgoy6sriA7UNUulLK8e09czRL
yqTcn7AK3S55eOfSYFLBF+mRHnUu0MpNrsDeXFyPjrX7PDdw+n03yqM1+Yio59eu
Ju4v4ouymjHM3FBfy4Z/PQy+9RfrheO82PtQbjHnXmzKAsxbm3DUcDTRrNE1eKtq
N1fOvC6BeC1oyLMlld3NcH5zdqgSfPdcOQ3kKDskGnnnUt/46v8VksBBP6L2tneL
htxx6wcsAlgMfc0zYSzVHKgdjBFYvIbfAKl00jTVI7pN4qda+gBmQJGhQnVVOIN/
aS47hplTSjXenuEPhYeGOd1gLMFtRkrrruMTW3yfabMTIVLzcP0Ug41QKWSS8KYs
lvcxSVQLEWWk4oeqWoaZ/+1NMKsS7mvuFhYmrqceAOjlRgICKyXgR6CecCgmkyI5
Ah1HslrNBTeKMPqXvq8R+NEHCA8tgcojePDyde9ZMMeNJtBEHRNiUgqJJh/de4T+
G5Rf2nzoLLepqadCJ8m3iYXaPu45ajjv8filAp0IwD98Nm5u3KlcuPUCaT0YtEOU
6x0Xxe9YW9sH9mMJPCaXpzu70r9agjqX8lHHMHM9nS3bpxNgptUBFvUplWfGpaGx
/R9ETUxGA3/jWdxBCHd0laDaU/rmKZU07c+fu4yV+SuSej7Qc+vdUpx7BU6q0Rbw
kGHQChOfGHC3oczldmmnCZMh9mcGrPuvTT61lhLlRHmgUYNVCOT4CVPLcE1cedsf
324Tka+/vMSzkkajQyDNwmJegxhqaJ+VFhSTiQm+I7FzP2y8oBh/63E+i6fvjxrs
QNnD2RzPQkszFCGsZGnpm60xipyvpcIpCwYxUf7I/Y9uYGQHp8XaKMdqfoiYYu1Z
fV+SjmIJUdtvEFqL3ICYyWFWqcUxZuv2UB9CiqRY5VclBUmEMBERrE+yosYQCGDn
7Gv/cqlIsN/dFFNJHEQxYSmXZUVyobAQTqsXLWQfMPzfeMgZgsSCmqhWx1lBBlEh
gPlLj2knV+InjmxgpyZ1PHJv/KsP8JxXpRQf9rf1srUwPXqb10XxwwOX5c2SCZOH
36CLdfpzVruSJ2BsP9wrhMmgPBlP0bZ0IBwfs27JNiYD59v60+CT+oRtWEUC2Fez
7+6SxoRPmgTRbD9q2mf0A+whF+bjKIaiYpCIorDacXf5Zf5bq5pLnyqyHSqTJluY
GbhM73COIlLRU8Z/QfjMstNzjf/T0xHAEN8wuL0UJt0PgdRURyGoMKpvUkl7CEld
+ORIOelvv4cX0P8/N+cPfP6RNZQV8A95FqjHrHYt1SIKFlE+TZPsslMXcT0Ttn3Y
N5zw196+7CaqZtf+S3AxZZ89AjFp87b0OcrsMWFicTLbnh/W9QUQapu2FsAVgAj5
3YXRk+MNYVN8KBbo1PjkTjihXbcHH76+CNJDNdX0UycxlP2190R54uD6vIrlKQBB
0lZzrcOygTcLiH8atXq76SZUebH19RLLdT0vH/yu0WlGop+wa5QVwA6IXkO4rleG
bKPzzlLozZjeJw1i/+soT5CTtnURoLhdsRw2V9eSpHsQfIZi5JBOwP0jWEt7Gc7n
NTI8fbLvUIjJe5se5KbV9LBjtg/oNcGGYPlfMiQfUR9es9pRHXGWoAQkrkiAJA6v
Rq8v0dNlpQo1gm9aCUx4uQVn5m+3WqGf/xH6HydAlCNaLnTSW8jh3Xu/pCSlKl9h
lh5v7VP8Y3UmD1todnRp3b+PvgkXGe5aCBhXYl3+AKAztysGrHL4nzGD66D04sAs
WC8qdULGbsSzRRTFJd5QKi8ZsIraWOKrmWEtrbjqGPjLnjmqUC4Xoopjh7vwMM3d
i0ZsDCj6QchhpT+OR7vVBnJnQzjhVherROmwIcxLPzjvNettf8hkaVDUtLTTwStl
w5WPI6W6Ih1YvaVdJ4xYIESA0Bt5yUf/E+uvvHbUmkrIwLHt4yWm2rGe5W+dr+Xt
5vzF6C/Dq5GTNSu3LBNvqSBRNm0X4rpTAhnU4f1+mvSd5NtrkRK69NFhma/6IGwI
9GJrirgB9ZwV8MbY2WT7rWOBdvhWwLZLmquooYczfRc8e1eM4ftZx0PigDoHb+d2
pO0CKWg7/25EE96nS22egyFKDuWrXYGvXxpmCeqEwfBmMC93TOoDpgLLQgS4Jket
xBJjMSLJfw2rKFeal7HQPINdi5t69XiG3MQzRTmOil9+mqlKnUFlhbhxOfFF8pRT
2PHakzKW2gFNhICqbk2hJah2syvgBhtUoiNsYRC4c5voepGGM2WsllPtajL2fXha
LPYTaqj8bNIW1A/0JN5+EabZE+GZRKzQObp2bC/ojvAZf2KBHQQubRw6DltUAGcG
kWYIToxB+FPa+R335K4twmTUW9153r4mVQx3QtvjZ2eBsTy0h6oVGG3ga0rd+89U
k7++9Br84xBGAA0VZd9hTvsq6zVKDvldhGQE8/H2zTCH65WYaYLSUrUQ2ocb63Xi
EH8FzdTgmBirdwCSteVcz43LHY0Y+ZhgfRjuzazbmqYWv6OL4NfXX8JubvkGli+w
Wu7/nfG/AbVNGBUPNuV/TSs8C/Gwe94KaTquOBoZaZW7J9G+hP/FeIBcSMzQ4znc
e86AZf3/UglAzlbuJdW7jpYze8O8JOFAvdC3Q2xmZwJNdFWukftzl0q68eIWEvOV
yrpt9dV/b5wo5nYtqT26zXk8QZEJB2+gCv0CIgAUQx/vKkniTgeRVxl2Ilq8l9jA
o38OLB+LHYySzoFZj99iL79pLHLPmJzGbPJx4D/fJSjecLFeTlFNF5t/RwIbY5mK
ms/WL/F7yWJJL0our433Fcqz6lQBjGs1NtmpWjtjiUQ7xtzXCVlS8GT3pST4Set/
OtsY00Erc51/iCVwS3eCVA==
`pragma protect end_protected
