// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 13:57:50 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
b2uP+y+Lvz/I4pUQxW/2krai7bJqUS3c0QXtf4Zn2tjaEOzg5WHzOAXSfNyH72VN
ML/EJqYTve+9yrYoTjqaMGLpHMYQcGseUX2piqV9jSAJddiD7WWHE09OEQI3K16D
XtU4N8/7qUPTOFnBB/TBm8Gg74e4qoWGTyKuDOCYtkg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 4208)
1bDWETzVpHdB5/bQMISUTbaOpuv6wyZ+LMAoZbpeUZZ/PzYLPcOfQkj/FfpbNER/
zsOjLuq71/o9J76qF9UlilahHboQNco+hSXbE23kNBzNrXZLQVlPY16r7XuCjSsk
fn2MkzDdtgzQhLIlW83V5j2jq8QJRuUcb4TIos3CMBTQspp9pxCjGZrWeIf3Hui8
1/rKuIADFmxOVqcMO7I+RIR4VlqcJu8/OI54qSy5IeL+jo52Edz7STlyneaauGiF
W3IceCKM0IGwrFMQPheEhSp1FEOLtqo+9p1wWXKIHpOfvJ91NNub3Dplcu1c173k
ELrW9S+TtmYImLQVHiXLS4K5GtS64VJ6YmD1TfA/qTVCBDNXSlY3gpT58qV+FDzq
KOYBcAuvBN7AxuEUS4+XU2ojo2m1qJ2PAp3BRpIgbKdcdw7pgL+oRW/l22Oj9EHN
QRe6NT83S4rjdhbv30tr8qjrChnWR/B08kqBcmCYu1UqrOsAgWcykGrHq0yEDkgn
miMAlMqnstU19xwaSOz5NerC5+bTwb9kXC4kELwsl2b+RlYrUqtwdH8dPH/uMlty
GqsHp+APpO/8y0K23/H5Km5ItJPxiT7HgvyXvy30BUkraPJ8WHXm1e8zN7AJm/d9
KTfOUCc2IkdgywdfePlMg5bxksi0qAc7ueU7s4/cAw6MYi3IkaiApmnPP02QnkZg
dpysTaebVjmTGbb1mWznYkvgDFUX9Sluk3uwRxPbY1yeWSdMkZAmSOBTBhAx/Jfy
Q7uzEEYBo4xH+Eg5wfPhAMCoDd5aGo8HraWaY2JLxPQtQlqaaYARv4RptV+LHy0i
pUMK/2bHJmZW3TQYKKO9DIb3//us6/RWjZfSIQ0xpIJHQ1lvjHRLvFykm4FffSNG
zt5rwvBO6SrHePgMc8KFvJrtbVRirTr48LZU4rpaLJRdCJKXeqE5B64JwSsRBGfS
V2YbLx7na2T7+bym186bRMR2Z5wbrlKRffRPwcSbodw/kY1AJ6shTBPNrdk+AR76
GoCadzdeWU+XPkfxKTD+Mmp0J+5QndZg5Nyuo28XRs5EF5rFPCKjX9xmIb7kT5cS
sGwhRl4Nh5ASF1TDFtOL0cScM/yqgf6o3pWczQjo1qjL8iqsXWk9b5sRJs7f42QM
XqCYKVpJ4ODcv0nA6MBp2wYXjIpGUm9mrCdlV8/BXV4c+1n1OrSfWJn1PhF8/vsg
5swztBQJp1dCguyMl985DIhk6Jkpc+dz/EVpaoBPcesrrVWZ95d0MGOGmByXDLWT
0lOEkc3F4K5GXKcC8azdxwWk2GtG2eTun4M3KRHuhVOwcfs8e5uXbylblsq5gRZL
Argd1N+G1oqwLMit134YzLT+Tfk9ok/rLS4kTJYY26USTsZv8SCAiK/cwUM1oL+G
xIgmcYD+tSBTASNFxWbd6UYasJ77Tt+Xyu7hhK6TpeROSSQoHfGmgnfAbvucqYJm
ohef0iQjGwuMc23A6b8kTpWSslS3JCyYkJOfT4U2jn2omcaiEQxoEhBooV5j3JHf
s/Hmnh5lq3AIQDakW8odM+YlaPyn4bQOCRic7eDZG87HoFC/YOM3hvzfivSQw1MZ
QpkV1LuI1AOFZwPxLbkMc3xioJYrqPHK0c+qNb9ojeRwT9iEeqG589kdEsq12AB+
RCvbMkOi0eRPt4V5F7hi9IcA6wg2BeMlRWpW8pgyKCxyDU/UlEhgxTaI6LbvRH0B
DTkofeB1rQB2NbN8znIGJ/SU706O5RtBUj1iDff4crR0eYXxufVh+z9QqQArykUk
ISa0pZTlsWFvkkcGYjviAlj/altPy0xGHT9L9FB4cpohyIyx/VLS5FIDMBJEtyQM
bqVtsjFTS3yT9J4bqwNqiOylM6OD/M8/RwgrFsQdRmDUODw6QLz3xXNYOQW76CH1
3Mw/y/uB3dm1oKuYmNsnnUpIL+PNb+31ZSC/4KTNuIPKNFt0/LtCsOPOymdzO/j2
ci3LrTKTn4FAzC3IJ3/KusbYrajdTHrCPBHm0Gcai6vSKMgXUe24O7ciTioGfmOo
eX6BnQmXYk7ABWA1P+qIllhz6JLwngB2fhcdr42Dd5JCw16uw5j/KRZPHChjKc/U
xCBkWd8W5rPz7GlV9Sj6/XT9TuNsdyrGE4IqckY6BpacO/jNNHa65i6J6J0swbnG
1lEdUUbd0undNTmSBcZuhXVZZiLseiqPaNh+y1+6fYM7BBq1f3zXnYvh6dZbb8UP
bFeQzE4LKctzHAKPWon30mtgIY3+fuBazpWWQvp6Kk4MoBAQulHphte/zIl+AwiA
SAneuPu42gi0VxDQuBOZ7diFOYdPVtFsSF3tbGHcv1eXVIENEXtuIrXsSIB3QtIj
4y/HoCUuuBwWfD+KonXhh8QXP3BmAqNB4wJINWVYjoVVhPWWrTtIfQOpAnS5llae
sxp/TmfI8QYfaDdy+ByP4MHel+xX0p1Lna89y5CqU2KrfmUJhnPjvBebdmNXAKpx
cDR+zTvU30jLh5dIFqNYxSxWQ/Vj3U1vHK+IGXzu4cixvbZgzXsusGpGtJbDoZMf
MBJ6u3uajPf+NDn3xfv4M3YGbg1MAa5HnjdH6RtST7p3M4/qQsBjuSOuwa7RHPeN
LWNZkQMMnz/YjIUZBL+b/2FI8V3ZvxGeJYpP+mGz722kamd175tTQWUqVeXUA/2i
fwTBE1CrM8hChhGuUWQe3d8H1uTIyH5OumyWTMu0vkM9Mc+/+9aUM6azU+B3cuWR
euyZxTjGzb+xYxGmhTNyFwYncbRwVjBeMKJ9N5hw9mF1hg/3a442jEFZs9+37o0O
w6n55MIsFjuy4EUPr+7BF5vFT0wOkswPfmD7P6oUGgum/272hrBHBdRnBJuJR8wo
06kegHg0uUVgVnG7NFu8BfVWfUYGhFsLaErVuxN8XL/ZlZ05sMPw5Wir1l55lNVz
xzfjWOw6tUKlkhaAb1VdSxrCNECj0H8U+NSWSbxk6FfLKPaZosX+xvFANOdwri42
Uzg23M12JD0PWsuihswyIKLaOC0C3fIUONK3bdiDUhwhTxFBaKrkTlNLEpRvGGvj
a2VHqSHmzaEPKgCtQW87fxe2Nz5h33AVbQSLXBDQBDMzxcCcAhc4lM12zHHhj/J4
0/1udRB9wK90cxdWeAWcsYhou9KESQ4bEu7FP/5CJv++yji3p0mJlQ4Ls7HnoHYC
yvMRpLKuZ4qVabTEIR68eKUip7uPtp+4lM7lFelowAu/azx5n/iBJcyoJDWzEQ3I
ABsDStauT/eXHI+GATAAtY36z3jSVgT9+UQchJpQI1IUJbOGndlqDgwEv4lTpIwz
JA+JtRmsZf5NQnPJ/WhPvbJ79pHtSr+odyEeU8ChsHlKDOnamitfC3tqAmnWu2i9
/JCoXd4pmLFx/b1a9m6719m2Ss3d1bPB6rrwUl0+KqeScPeqs7mDOYtvBn3CQKqO
AYHzann2yUoEGqq1qg7MoXnqhwKeHSjIBkNWnLqBEwWTiVKOI1GXwHHEhpeOD/XZ
BMt44qsYe6s5pQ/+njaaDqT6zdpjwcHiu5aBOwFP4YN/oRSXfjFxIiVOqu+Q/wl7
I/KERDyzmLor2fbNWP/+OX2xBWFDoQgTnD8to84k/HTFNgau8utPgeLu7wkgrRSw
FAnJix62EouPn4B/P0G06T023Et3f15c4m/4tWp+1xjhUwo/gBMYjYtZ19pA5e94
CPv2GL5XD3fZe4QoY0FhLtlZkCvTBzMjGebfaC+TXX8uxPGAKrD5VCnYy45yYgiq
Obcbb0EU+HlOH3fCfQD2ESfurXExRuJuLLVyCDfslFc77W1AiOoMBdBqmz3QRbF4
shTTyhECUpaZkSHez78AHf66biohSBA1Q88iIlHGHZCth/wGcznEEcOM2EDxFUqc
9FnAD6ovgwNH/LUoqjytwEqIfH771tg2NLSN8RlKJh3OweFlo3t3MosxQM+/RT0G
SNxD5ldagAW+EVnq+R6lUHqOcDTlMzs6HQVBHOBp8+C4cRx/jP8TlSfFA4NA3ucF
vaNOG5zzbuWci/TJxEABYXAC67EU5fwQAKaV0auZCVcg3JVCX8kmMH4yEjqFSeyI
RqXIRphp/6TuvHDFcIWHCTjtl/KTOZIIC3uupjTTqKSh0ik0MCtHKCR0H8tO28hv
Qif2ALvcpzJCqDwCSxnpgunRSs3ZJIzHSRLsOZKHS7KWcxrfsrw4ucQ6M20P3epj
xXjpP4QmcvCW0L4hMJSlJyJNQJAxm9rqfUiV6Q8nWuclljAf/hVwIAQmCU95gGw+
cyqaSKQ8b0EFaLAAJEwBQCzmNIG+otWMekmYaF8jZZ+Yb2uIog7CD+xUQa8DuJqL
eO3PCBTsl6V9x3d7gpc3B1gdZJ3jOTsQHmis74hRdnwyCCJFFj42/F4LWOL6yl1R
TFDjD6Sq6QqnF/Ysm4YsEXdDeVzJ/TD+P+2ubyUtjI4qkQDvj6pTvrBSGWnNjWSc
WOvvJUKYnxKEF+mmn8ufRth5kWjyfHxJAILK/k9Flm9P15KIef/7fUh5Eirc2gkL
j66dwHLSeXvk2Ko1e/Szd4rg/zwpl+6nrveKi2R33rhmAK5DqRmXGj0N+vM3KrNA
+17ruLgz7VDqwoHv+6G3hArLZnQ5exGoG7ZUnqWx+X0tl90HSe7kECkIet3MVjZP
N9TrHlI627dC4CFXgjJIpvkBqK0LyjrP6WkqWm00owcg0djoWSFcUR/xYru6Dlrh
Bpe+JP+p+v84KPgs6HOPXR5Gi/TEPUX3oYJeHJtQU44GT+5nQDsuxCAARP2yCsNn
dryKuSuKcuNrC/+RsCZMh14AQ+jjabjolUzbVHfKne+vsqCC0RLzQt37GCmUvPVi
yTMwXgusBXopC2RbIZDt/aV19VAGVnHLv19lXqA1rX2nkNQQSQIb66ibgwSmKu7o
e7IqIr2L4SURLn82eP+JyeqErxP1BxFznGbn26G17NxdPNTygnczWR8Q/1D/d1yP
KfgtVLdYgoHUPG/Z4OApD0L5nicFtTJ+4Rheavzl91dd1Nq6t7Inib2FKaPwfg02
ymOr0L86axy894QaKUgydOpNBpXzjptpQ/sdlJTgO3ykIK/c6I0HFm8dZZXCE5DP
ZR7rUUcJ82Fnn63V1GfeSufxUqgJgUGhkWtIw0knJKSfS1nUbnnnDs8ModtteqTv
wVoHTu/cgHS0Ap4jMsHGe6DBv29cGbZG//dUusaDi/o8dineq8uELeHlxe8uQr8R
be6xgYJgSKgjfLFqKxSNTtkstqM19kohEVF/Swr2HQXz0T9HyoC701UMVYCyRujy
eY1i4qIcoT+NfjRFpcFX9s3QMoaxPCHicYT+rN4EHrS/J72wzC2/N9DRbQl3qu0S
RJIAX/E4ytnqJZEP025qHBSadp75oSwBJmEdSUzIClEaeFaCUaZs5Ch4Qvx6QY2V
ys4Qv60vJwEzIWv7A5o65sXWdUDscMb2+Y8v7X3yimBbmUHNkCv03Ve8rPYRWcbM
oXtlfSAbIaw0CnqJlq+bNyhdVWyEgTR0OwXieZd2yOvTIj3n+HLlGNdkBXlmL535
42M5gEC6+UFLBy+6gcdPQI/jSHR5EFzckZhfaK82QZU=
`pragma protect end_protected
