// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:02:16 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
PIYwMKNfcPi+HKCozgxvbc3N5x9pxKansQ6Mea7YxwEo8KnqX4UcCtWpkk43ViCd
EyO/RHdWhSnwos4zeWi7Qz8pWeWOVhcpbQw4H+lPT4VuUTAydFRCKrphFib79SpA
klURNyNu+ah1y6EaLrbzGkdhxEu7j/ZSwykyqmLU10U=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 195920)
uKKmTNvv9ARUAlnkdfQulfrX9ZVK6fdxKkMVCqSfM4hC5Pid6ubZmxG6YwOOIFaa
WGS8eZ1w8sSz4ChfS7Mp14K65JecDmLPmw8tEywiYWptMbx2DHHx57sKpPRPaw+O
HG04SP//nMt4oyyxZhCUACRVZwOOZj9QXLEuxwYmv7AXdO7yWSBLK0iFt5HdzV36
QHQMuDB9QkyG8rAQEpb1R+Yvouxi9T7zn9dWbJCd8vrWiF/EEv4Nw7Nz4ogwtrt4
4DeTqvzceD1iBfvuZ07ql9cPwEH6EP0kwVRFAODLNTEnoisJVKhxNPHMnJo9gx/h
y9vtGMwwsh+9rsvjoW9hV1aPwMX4BoTQ3tpROOskD7zyCjz9YutyomtmGc7y0FEe
/CDNYkdK6nvVNWb2fAUPgUqmZBc1zJAmW411QGU6rFdZg+L8a0VzvbvqFKjinwEr
vBkoXRfh3epxlHB0GBgd7y1HIIetay1v0dbTaRfMWObrdYCqVUZNevZ/DexuNjBm
r/x0wa3eu6CV4i+jVSIkgIvS5YsgGMZz5D78S4zfE5mlO6UEFJCSm7tYy0JnkHf9
ZavgJsG038kln6u0+RYuKhtDXA78Jj/PK/V0CV2kOed9UIRax3P9/WP/jixNO0I3
+KwbeT8CdyyyDCOWm48q//U7ZFul+Qm+/flnbazZvPEb4CY5w7I3MVIvkLZ6CGvr
hK7N/elwJOet2PQ4VCDYtM/k9SGsxozdAQS+x0yJpwzXgr0q4Ub6nYzVlAO4XaI2
QgyPXYZv0GWJso/Ke3ogdzQ9pcVcsR0gcFILVCUuIlcsoOsdjUE37qkkmCUCNSUV
s+Osih2Z8kbFQDjCyZotYtLRqQbMbdyBjj+CaUB8ahloIaWdUrN+BTKMuJXdCQMD
Q7ykqcQPtiPtE7KMjmTRJ2+LVVRYGSWLgm4Vah5AIB3YSepSlauQ0tOJ4QVCFLvS
7ABDm+Z+rc5tGlliAuy3iaAKAzCDSnjdmutbo8AMQcQtKf/BSpCJ6sAhAKaR9G9A
cdzGNkQs+SN3x6Uq5AME/STeVo2i4GXu30PuyS8MfHRGi15+mXn8YCOoQaMlz26W
ShMD/4IU02GC013lmwOjchpgNF515iSo4sYTeaeRmowujmCa1xE2dA5l6W6AP/7W
aKUdWC8jP0vjZCEKLnMOFVxqTbvdx4TnbZ/O74CxraczTS/ulyDn5l19b5l8dUFm
3bG0KCmuPPY3XhL3CWL5A0oyrFkgFyuse6QLsLwdZU/dWGgX2b8xdtUDTqxAK+SR
KuNDjvNtif5rz/zvuPKH4X5JqK7aQljZOUtMHosOvExZk8Ux53zLm3l6c+YeqLB8
a1vB5vtNAHqitMg3lzFwtS3o45lPH7SM2C2WQv7sCmWEyJ7rZ8euJVvTRQezUSj7
nkSzSX012b+Rytn/JZmuzOS57pfbJD3oR1vfycepkCKM/kysxYaEwT/YZHTpcWDN
u2dR2CqREuwxQSAGpswKvc6T29W8W31zUBsHG4lCkKiOidXxWfwKbOEJDZtAi1Oa
kjT2Hewu2GiaknMaxSvXyc22wtlhD65SXIAA9K0iUDslmr63Nzrapbpy5g7JLqaG
TX5Bzag8Sj1RIyotfu1ZUUEmSjomFtOwAyyRYl9djSu62m/eeNfnawxeDQem1GWq
PtbVWVaFLhsEGpEWxBW+5vDDBIOT7LuloX6OxsuY31CHvYBadW3TgsrvKV9iww8i
hoOTsu+esdL4uULV2/9ZpfT7QD99XLHTbtjmq2KUQuH7mB7U50RWLLLxF/irs55S
dnWOkv+2HvY2oiwCrowHDedmcQCrPiaJqZRDTYmPI6U6Emtm95ibXPaz769iqhSn
oJGzG8eqxpyhu2vFYP4dpx5CFfDeKEXS+YuM1UHeQpNKIFySTZa5zCwspJq975ft
DZBiVLczkg1J1Qnkw+eGUkRMuAyQ6P0v4TjCY/eSU8T4Cil5EAz98mrz6lRs+YsB
2Lz+ZvEUryBZnu/ntr4uVIZDb2vpInWm8LtnKrNTGvf23tCyw/jDiVqfbyifvgIP
rGEHNh9pll7Eg4ZraWmWd6HbGu9zjWoYGQgKbPWsC3fRVXLMLIU33tlG2sPSmEUg
IMP7elWZDr8Vhf2TeYc2cGDDrQ24zMLtfneaPSH1x2hVmIyeJwiNmR7wwYjpVNXI
UNcJTy/CBMONkzi/NvLVnQifHoQFi5nzVn4KtH1fnD6tG5E0qyKyN7/qxL2PiWd0
dV2XkyrId8uPFXDHgxfiR9yAGK5lNtthJuIM+MlD0tcRDAW6N+Qf0VCXwnWWayQa
O7Dj5uOQ6gEuyxJ3VO4t4aXfJc9saDPqTSAx/9rhPZB2+yEM4BhMt1O0MmCNKTfU
r15gt1nONUp57WHBkoNGTci8slsEczbnO/Len7HE1yODymt6DuN6BanSLRQ/RutI
Fh8hNGR8hiqP4/pXuukYw/r+eWVVw5ehNECC2uBhYx2pQEHRt6efwpC89QGcbiTv
o2qLdfLulFUpCZ+ppT/F5CpegnEqrx8jBS5HhzfpJIUQX8kMCWBON16zs60i2Brg
BFSOuFzgBgbAX/3215Zbuqg7nU47KjBZThN+RFN/E+331bi9uWVHgPpZZJ3YRYuK
T4u0FBDO+3OChlbW3YofeGrPs0DmP4SZyKoOcxXM7LxdLJkvOn+V8ZG4yZ1FaI7i
YdDsnDAPo/ekBfMF6i0a1Kwf9q2yGSC2mb0JIsR9hxiMeu6unNeswaFRm3ejbqWq
YSYEQreZK8a1BTh8glw5/DQ9wMEY7l0+77NW4U6y/+Yhe12Qc3HfmsZS/CyMazmO
J0MRaE766C7XGG9beDTSCcGdPAACDH2z936H63Gzz0KwcnIE0EYqx7eEP7/8bsAj
UK4nWipoZJduy9Hjuin9yvL5Od4JyRf6weH5UCE/XChsuov0svupJzeMLoWAS5I7
G8GHzbjr4FUEGWb1K6t6zBOcVT2mcWDEw5rtGry0jyr82QCiCYnyxQSMBpSYkm2q
n8ARt1ltxGJdeNO3Znd8uOfNAW1lmT8MMZtordS5rZRLG3IWO0R9wH3Cpab5a33R
DbAJDJ/NUB6DigAG61zYdKYlp9Kt3k2ie1/QrbJSaV8MWYiHZSk/0mF+KtWKtk3z
QYwprve0enNezBI7AFKlXbPYu4STJSQIMuCNYOpVXzLL6bbMAPc4qsegXcy0xR9P
3vxLs8pTNQ97a3lfVTvGVfy4978LzXs0aYORd7p0HqMxH2Vu0uGUYWvIgB/PvpX2
lTtUGmgJk72cg0PfPCNmZHqmkfm1KddFoxFwcaCOWTj/dVmh+rtUAvQvOEhqmDXr
2f8vEjZlhnrSozehC9T0d0cxebG7cly7mRN0l1j/82ltoisF3W10XwgdPyGopZ5W
3iINH9zKlwlqFH9oKrflN1QmjbBZ4EnlOlvjJE67dxhkzUaFown5YR3lBeA/LSHK
T4MxZz5KCBWXPxemgO3eihpqkWJ3PgZDKoWfRUoxHDTQmhh7PfInxW+IEp0IVC+a
wTcl7u12TgQ1yKcCEO1/28610xFvVEi/F+89JsK7akKFoEuH9tWUHOmMqV+DITjQ
zJ+IWOUja+G7twyLSd74NOuAMgrUPYZ8oHz1+Q58+UlurOqOIgOIxpzDOb3OTZy4
sX0biHAIYP+KdKQNQLaDCgCES+QDBtyAdxGNhMmHlNSU92WpVHSx/IVREvrbgKFG
Wv0rhJm3rgmcb81i8T1oeOXR7LTsdn4+bjm7qUHnvTKP5bCPRjp1nyjOsW1vc0ZV
mK2Nf+6lTcALY3YzpXoJN6N8Aq4gfs8BiRjT+oCHOMECIdzpnSWCipUK8qiXzzmb
df7xITioFprXdU/QmUmtg1N5yGS2uNGPsarC15S7riClI9Q4ZbPQvVyIRQIjBkJW
W99vem16eEDEOTTSmJm4el/ATge6AVV/wKTRDebLafZ8gB4Jd13HyyvOdjsGTURy
GHSM03RX8iVudgqn0XfLmpbJjw6GDr6QLsSYWn6fwLc0KL8Mn3uZSTuKAQyOhpix
MJd8FGfhaTt+VkBPvx+ES6e0VC0ML/eUgTjOwXRv2r+rhlQnyv1rYHMgTyIcwz0W
gVbfQzZRr0KDwJcYGQDL4XL9Cai6yyPMYMtcBVvOzeWmrwaWS95y47/z2Tq+OFKJ
GRkgFMfo03ZAkQEuQC2+hVZwmkv8DWAQDD6E5gzmyifO2NxY18ias4uOqkmpaK6m
Mx7gWYl8YYdIfb7zThr4srBezwsh9M/8aN5supCCA+gvHvrceqGRzgDWpZbgvvv5
vkKGa+3xSoJ5CsTBG4igTO+9ii3I35hGTc78hVZIkOZV+Ti1k3AvyIbnMkMHGPSc
dS/DOj8tg1ifjbWa6iAD7XfFEbps3kHOAB9qVZeULNlIIY476Zw+kPJAbN1RPS3F
11H7u6q3MBOzR6qZy5OQHjFvu3o4llmycpb7+R4St3/ZXDTy9gKkV9I8dLCK23ON
PdTPHg9El8YWMlbT+r/HypLIbaiCJ5niGcRxp6VoPu9j2H3mC2b+39iYpsa/wmW8
OMSfpkBEz/854DHSpToULfmdk8UgQdRPQ3zjvy6Q8hsY3OqWhpl/foo3Ccl6JB3B
YYXSSdM0l6kntkclPdXPEwgLfNP9QcMbYIWUvKe4RXT2uiGRay7M/+wlyuunv6yA
oRJLxK1HwaU8icCD3H/6xm1RFgChGUSJ3qzzrTuwIpA70+H0qEHdO3Du90NeSPqr
CuRhRgG0KnHMKbSTX9o052+kolceSiwjoCj5fZdrJUv7gO4K5N4WgoYppgUlPyTE
JNpj+s/xf9WL7Cueosr12rDll86UgLd5N9KX+Tm+W0n0B8kZRsAp44SQq/uol6xK
04Vy6Zkn03d4yRjrx/b/q4FAEAZxKz91ssNcU9zNQwX7cC7/Nq6SV3FVdokKUkIH
VdY4T0WCIqVcRfRtA/+3cUs8/+QqfMVJqSqjZUKfzGQjWYWyq4YEYQk31pcFq03b
030QN+7VMN5C8klOv0E+qgPSsYM46Fo0fm/Fw1piLuWhWopo/lKKx6SgS4d8CwWW
kLRxKsPSvl4tP82Ws1ZjZePuLR4I/N9NyHYAslt5pNZsjFK4/0d++drsH0PeTBk2
C1q+Tu6u+a6aCsUnE/MSKpwE8Ety+QyePtCUkGdb0Ultlf7IUTDZZ3BUhYv1R31M
kVrbB9FLLG9IQ+aigL9lC/nAqur+XXK1K2VM/uYYjS3cMgbfTL71Op32a/BacWF6
46bMXC6vdAJXUPEzBDQxCpjBPVdGjmknMv1YTsBMlNiH3fIAHlKq5B2s7pJk31TY
KgNT8SIcNdWuwnZ0FGCHSzmiN7+eshu9SyN89RZOjiOf7O3R3ZW2KJbQyz+vwffm
pPqdDcxDP2Brg3M+z6rM6YvUHK/aX1K24155Rx5qdNoZflTifTqu5BfJTullcJbB
Kuqqtmd0zkGjlIMKdbx7NucQiW4GQHD/wsVZ8yvU387Tr/TJqajzbM/D+LTCdsHR
CrkU9VFIar3aCjCQVhb2pB9B9bm7uu9gQCFAvhwaSeiOCAYgmfs++Ae1/AVPWlDd
7uK/cU3h+0glYoFYPvYi0AjujqccyncAdo1tbGRwOK0LhP2HVE9AwlilQ+XYEnC6
s4r2oXCGzK4IHrH5rbKstX6UB7kKs1urbePSrrIX63/3I1wt46EQbXuxPj+JN0WA
1typcliabsfyAcgB5JlSsIh/JsJABIdrEEs0v8W2SST7HXyQnd0RPrhc/zMO5cPo
DS2dg067e9nOwX0VscoJr6F7a2ltfHkc1W12TfXAnrMsYYU9kFx1Raj1pFiZ27HE
Cp1/LoBbjgYJXXsgopFsrNZk7DQDwQN/IKvXmlZGEutCNM/O2jPH8SUt8eL5Fxq2
Yxuw9BSaTz4jItJnnqZS1/YsgkDFW4vzCUPDjX2xYOYz9Ls3nFG6/OuyC3SIc61Q
p4+ok7TBld6lq4WXuDZnpt+HxGo8X2Na0kmMc73NXKGHkinMm+pTG8yNnBo0BV7z
TUWvfRdbl2hoofJQcpRgU7z7r3rEHZJfDQTInT3/pk8I7b2gLueB3m6TjNM1GB1f
CW5ib/KCpXbLQkkY/TBY/AXOcul/yDPTJOZThsoEIsxrGow80NbKg8CLhrr2Qcqv
h09QNJDwzqn5SbJS49M5eFgxqiGwUT6HD4vUtd1ly0daHarg1ESDeyGUAmbAUuXu
jGa9X2mr06QAEdHqgCFt2oYgOG1eBPcpr9DeQ5nvGw7a7lUNEmEREKWTieXRqXrq
wmmB0Gd9/5PCs3MN+CTYnoam7zGMEo8ADZVsxxYorh6t5AoipdoQhaaalSs2QXW4
Ub0eY5RaT0J4SYj5apF865UkhUHEXRGNUp0zNGBwMhIM8c7RGAEqEY851j1Apcy9
TY8VOeeAc4cX0vmGI40Pwh4Usea773mg+M4HEca7EloFpB6x+eNNiKJrjoe+GFgx
/Yv7R4mji5sfeY707HWj118nI6znj6yAE3G/eQUsR6QOqX5H5Zfmwqj7cONzc4nJ
8HmQkHv/m6KHZcUCu0x3UgO43swzS9aEORBiqDxVrvXuoUUl87FvdnJghUn8Ux0x
+YVhYUXmjlO3fWlHnO4S3V8dbMhwVSeQijM1CsGMGJmGDO6VvZUg/2VpxtVFrgvb
sV3Dx8U5VcJmBfq0FIoOckKhDd+pkuN0wdJMNx1TVaGsk4dcopDyWAxgzzL3Y4x2
x03qP+AdmvnoUYqNkERMiQ7wudL75HIHXovCeS8ew+j4rJPfxWIhODJ2wXt+QvGl
6t/GFEUs1FAPvRrEiOJt/rNTaY87ZPFw89XK39Nog6YSEZGsyVf4xGLvCyaYj2yT
AQnVl3qt6fgGaGWHjbDRurkgUoQFeRwlpbk/NtST/0yAnBwH1qAj+d7fnA7orkJP
Y1p/8mC5OyH4/qQGgFnyijxCHfv5lzpvx1SQRRygc2FjMfSSVfT4wRoVNDUADy57
TpqA+zGXCJXGRovae0KWWmVoEFRHollzJBaNiyRkEVhFNrGyoPxfkxuko/lUkERH
1KRo4I5k0G+YqD9Qp03f3zF3tkHv8neF6TUmqEATn068tdVboOAfdvQ2D4ZpdoSo
Yz3K+/V+8/WmRxoWy1yUuq9kowVcKY+umnwS61vlfk147RIJnF4VokZK8puztOmi
/myQhc2wno7lWFs1Jy6Gi7T9zPsRDVMr1XadBlQ3FXBdCA5dS8MH2kX+29b+yvwY
duFL2ZNmnxz41v7ZCkstPmfahOzBPVBcfNmYUil/Fx+NCZ1rdafcAf/TCwM4zo94
acFT2fU9tX/rHBx9Bnjwfw6/he9bM9gVm7NiGdAygYynhylyNHVeZeSKDh2IL1Ck
k5Unh9O7B4IpW+azEq0Vv1qM3mhCtTZhOgkcgi8R/Md4mccYtvSWAXIVNm3oNOYi
62nTAMZJpPYPFvtMYOdRhVIr3uXMfDutcQf2aFDMDK+1+7KdfK9N1ZlYnZHeXpSX
X8Ubowc2vVjiqr9wYpKYeYt+fLGhAl4aCv9UQ+3QiWCyYx5kpB42SJLhIc/tdV6p
CIQThEICMlEW5tXXGm87/USzp24Z2UOT841cUYDfhUnbA7CwrnXBwUmRTHNvwTip
t7KgpmMWSNndThztYdge66VN3Us+py5j+lf+v+FuLgq7ecqUIknenTIDr0wv03Cy
sLgKC8qHNMF3OXyVB/AzMH7Cj4/+E2lB9FsKFVwx0kzOfthEfZKCLGyATAPgoC7J
b4g93z92t19HZDRSQU2ZLuuW2tJzPwdu1ebtlpM3UHZoskeQ8k5HChz1Wbawdzxw
096tTv/P/aRtWKULlXGLt5h8D4mp0ZHgMpxN8AQKm5ziRBPLPgl0U1ldwWwoJXUq
2YaJf7Z4Y/tBgy+JkNlYa06RtFIE11CPgl1PMFDOxDi5rORTIdC7dMHCSaWDArQW
n/FBgs+NQOxu9h6tixtQbSyNQqThVMs3rcFTucIojeuhsv078kghTMyaAB0L+hUV
OpBp+l46DMeagBpkKu/c5Vy71+/Pksoz3VSBdi4rhsCJYQwAcSjPumSLMPAc0Wo5
cn2StDlI3vgiREftbPMtzNGLC2pgFDV09pDETA1e2nvcT0I9wCpbdi4eJ2WozYsX
ZgxYXUldauQg+bN7gho/H/5Ee0q25FyHBvdjm4TCrSHv8K7j3RPUNRusXIJhuO15
JZkWtmqGCbF22RWrZXArVUunZ3AqR+qjZdkr1LL5Pz6c2ONMeHnkoUaWHSTNy3od
kc13qCV/tJxH1Rgy07CT2b94k0q09p+9pqcQBgZDD0hYt1ogcm2aS1bl97kiJBun
S/8qbn9B4iHVMlSp+AN0TngBPFcSvPl6RR3IEYFnOpzdGHhBzN4AgCaqh5/JEUEh
SaTS6PQgp2okqezQb6vTYdv+ZwAKtfYUiLxaeK2WlLeEsDNzAoYRVA2nxr+aN2kx
lq+5Lz/aSq4SypfVQa1l4hWEZ5E3vV7oLypi5ccO6sOhkR8uUqqUgWMV2OKOGJ9F
9PuMzeWXn0S5b3XHLk8blEvDr40xW4X3cM3bBo/K2XpWm/Z3TuAKRPXTdwg8FkMa
eQNn9gwfz6LmE/Asny0El7EugHRtmcggQjS+/KVycFAPc3shbnuIdJFYlcgQnSTx
VL2wMPUa4KFph5kFqyENjZyYjHEEylZwhfyimvRgAFdMXm7zVLEo0PhRIacSRP4f
+2MKV6fA85zDoVcC6i5UZSeNqoX6L+NcwH+PM1rUjg9wblOfF26v3e4pF95Nzxvs
4+qaWTmhHW0wEuv5e5mjyTvvSWRYGckjQn7wjJSjVklUnIGJn4erU6XrrNqBVDlh
8PDVmFfVwYB1STfNNjHY+ophTKHFTL8wnpsBrt25YTCXy8qSNSKLftHLSJM4OxPl
kzcKcddufLgPEO5WY8mn3gPNdzdeA6Lc/ABF3S7Nkv3lxpAeqwF6ZNN4xgE1EF1x
vd11Q5Kw8p3W0wd9FwR6UZzsUDSr88x8SGPkdZIGj8vs8e52KuiA4JTp55+I/rdN
H3kXMPPEvPZrPR8yq9kVph9oqeja7ojAq60gcsOSkr2iaq0I09wFTwEkHcJKIbl3
RQnPWzdcz2ljaW8m0dGAkqEz/oNmZ//wGFxm/z4nswEqCMS0mZEjbrmpOsTgTWpc
JECGmhxmQaaAPv7l3kBpnnuoerkOEY1/FwmHZOmRs1OJGv/h+iywP+0Rwhn/MoXU
px91TVT4nngfvCpLBWCbbcT2USpIxQBm2r/pfsGsqe9EvEC6rLNGuXKNnGr9Utyp
oXF9/G7KrovI4RQxoR4KPFd42bKSo0DHMH5Vawwuesnd6+Bsxcbg4HPU6gDhn5Jc
TUEn3han4o7Dx2Ju4Z5fqQfC72l8eCfxRkVGtOP6LpRZgy6DMIchck3c5bUf0G8e
7PNWAuxgQYDKI5prRBWf4Dqw+/r2kojEL3iPG+ljXIjTjxyWp0INypr26Piy1YcO
5ZwEtnawj6qMDcCsfgZ/eiB+00BI48qmw0ihsQrKXiR6U+VQD40IjNLIkQ1eE9gA
6atHq41IvsfAna1UfRRGLexAG4Id2nOjJWYtDQD93hKl9BiOy41nudIJFMxaxwFl
GWWAIoThnJs+SeDmmi0eIemKnSqAZmPn3e05qZIwc5fGkV2wpqwlTmqX9r2P5VIo
+GznBLX2ySP72HHRaB1KUAP5aaYbjp1fzFbI91YP51tzkoGHM6Q9e7TouKE+ZZ3+
XouQRZ3U0r6Tr8EnhxTcU+G2lgN2R55KRcKkVVKjqImRsZa8E3Wn5dLEeAz4ydVk
2v2FJSfrj6G5hNcHNSf3x/Gr3YK2+1y2pyjmupHfyHeYPdkxOAtY4rtDIasFPdIP
8Fwb+4pYPPpOIgBwWfyrz1nNc4z6x6uz8OR9MxqG6iXEHR/MxzwUS+eISyrNWmsz
gLbquB9R9IZfftWr6W83wD9c9sP2QHeWWhRJSUp/pN7jl4rsVXYYHyhx6Qa7mMe8
ihsgXeFJM0cWOFp4QGogLsiNKlc2bFg8Jwzt0zBhtzu+2bhHJ8pQI+Wq6spj75Yq
CEPRLLfVnKLsuLFRVr0gbI51548MPGNTlEe2nKBU4jIkifwQKacD4ZPqM3+Gi9Zg
OuskIj8LULmdT3K2Y9N8D58hFngnN+6aakPy2x+z2or62M1e4d2SsCOzUo5ATXkY
SWBBTKJppOclEiVJlBfEW/WX4Y825nBF1fE/m4PZElq/aBeEfB1q5AhB2mEuqd6Z
KDU88+PsGVR4MoKWb+v7o68xnw4F5CkBiUYG0owzmOVWFYC0aMK5jRpBG79Swqi9
tnfrdECKeswWTl8Fl+IZBjEIej86eJNc1a107V6eReduauUMJV6fVVTqD+Zt3oOd
ReKAQ2H0/YPHSWVVnpvuPGlz/Qmojjkd+1qQkXzBdLwhhjLpYVCJk8F3ZpLI3sji
4MWvFtYkPhmMPrbsrioyTBhrgfSMNKG7huQDzeukcDNgWkCrdNsy1TDQ8GiVJQwi
OodQDqgyoWUX6yKqzBrW2jU4VVk9+JKkWh4x+FeGDNg6dGQHozsrKcGRN5IUoIMc
5tMGyzbl+AtpdRcTMrKb6Uj0+fUtpt+rEv8tCV7s8CJSTNlDNVguQOeM3psEINzc
OaOg6AcN3UdXvjp7D0y2Wg8qoxiLQROeJ/CWJK8nWSnv00nWUVmFOYd7BqMjHkWy
RJBKqwTrNxlztMaF0Ooq9CWKjTeJubdxDr9PhjLC/IYP3vcrq8kshrxVg5PsHMQ+
mUFVEAOKJtv++/ZauBdzJQvWxSUbU89IgX9EVXPEMq3N9LicFBgATNvBOi31Sra5
Vj+H7QgBomSv8z8knRnWfIyQisTgW+huoMgN9JYj9lpEBej0yi+mPLpBNwuYL7PS
HuOAlCR6UDNCBy3O6Kdyk/iKTVco8uh2gIlfYeh8mV6cPeIzzSJwiIuiBp+kzkGe
yzOzhZoopavzX8dJmFfzJvjmeTuHhnP2+SrJ1XBLylX5d/gIyX0u1wgyCnYb0dAM
J69+CI6EHcGPPcH9x+4NlwI0qB85kmvrxETYUZQNlkel2YFmt+GPywCIIp8NOiNO
mechvBTFm4vNqRik9k1bQHW9nm6gnjRKUccdr98hnttd2R6FgEXK6PPR1RORORwE
wxe7/o9JTBTy8WSfZtOQ1WfHQgYEJCMJVsQbzsQJTdPsgdpDJ1hUvIkx+HLNt9g9
QjP2MGOUuUr+tgk8i9EbyGY/4W01yy4/HYhip2K/rYcEqpBUeH8kHlnnp3iS23Pu
HrjBBO41gfx9qdtcSkhd6/cDFS8zMRjIu46T6xwHIGMqrlgB1ta1CVcz0zAVTEEb
Rx6rDz3vUoYTFTZJMHd+FiM1nTEkbp7Pl2KNp8uD7aZSmem/msEXQ/psyXiiXyjh
VrTvawNXyjJMT4rDx7BKhJ3T+N5bQZgMSxhaLogj/EKT4hBR6TniouSOaZF07Ws/
q1GJZkVEBOOVi//hEVlNXWPzmvJw1TQVFDy3IkxhdYBp2hSryXrAqqWTIwi8/xuc
GP8og4twL3rdK32464m5e3/KxIhF7phjoX380tRCNEjan0Pf0puDVjDzmXi74rzM
fZ+AS1IAaYEuZLQFnVWIgG1rBsW2yYRyGg/9QP/olVXQ9lCBH6td467n7cwAwZH2
2lXOHJF9/2FpW+fZVCAOm7UHU28RWX6TrmnL7HM/wEBm8R5+ZJXjXmJUyuAm/wTn
F1ydmr2EmIKPccST+RbQMEwmZuiPUZoFd/WuwwB2t060A1KQdU4z+b+wSrwDM1fP
57qF24CQoELxrHCfjr+twApRQt84O2L8BPwBedK/ttaKniXfPSHxbvXJ+JzaNFSL
50UOF8XF2DYJV8W4ZVdfFEw6B6Oljp0WAajeOHBP5ZsiBNs9Q/8Ej6qOnP+tEixU
4pvjb03q0v9yyuSbso6SjWiZWSqoPL7pA+mq+Uv8THhN4H/b+xaRT17nz+B7ShEG
cbmZmJlbsvC6MmKHpWBVsV9g/Ehn6h9p6vbrajUy0gxZM6NYm2ORsn2CZzE0k6uD
SEi2H4EhUcce+vpNQQNO/3Sqo3TQ3zpJ8+gonFSaUHr5SjanB5OeU7KdutQ10FVS
+cb+kdx8uzuMOn1rY8UQEMnrqLCU1gvjarJJVXr/Vt7ktuwuGPxxQ3e+Ai/Gg1Ry
v48RTJmjlhzqJ3e1nm1Z7h3OIAvqEjjkJT0oGNxH+umUTr8xkOTlC3BZ7XDEH2fw
qVGtAkDu8mZLas8EdonnqWgDkcZV9yTDotyxEVMxAF097mSjaUL+cPHZnMKLn417
0njAs9Kr5eKsd6XIuxVZllUceUCeqjbTxmnGdpUK9HtQCPq+kRa/XYoS+dYr6JHX
KwuYmip8gtfHZjNWyPErCflu+06WUvieHs5hS+hjZTR6J/ZIPZyICMVKLzp4lUrP
rxmJWRjGY5qknrKTGDlOFdZdLapxWA8PYXBACKmaqoLEUoOWP0N75M6kXoImnJtF
J/y9zS/nXyhkPcvRMsCvqZ147Qb+JOcCH4KuRZk/zaFbbwhsZb763as8OsYsL3sK
aCOxyH95urI1QjsN9VczfOaQlGHqXHnGq3Hx82mVGQFz0Y+k829pLYOqjrLMjjrV
H9MyxSRPrPe+u3fM7o5/7PU9JcwcAJ3eKxm3ZT2yzY7/zi8hAxLY9P8HRlQSl6Uy
e1733mw+sENljJkZHI69u/1QOIy8FncyVZhGjZayo+YXNWR43rNzQYMxd1EEuj24
S8KhcY+SYvF9PoKMavzp93eMcWuGuoonkql0uQMKQ0nQbGjtZNN+YkCvlMIyIvU5
+tWO0KXa7E2sICd49uf65EW/43T3OKcYGgbPmRDpGJghH47AnKpO+gijArJgeHpM
Pq99RX61lVOm6pYDHWAY7Yueg50WBsBtsSn2wqnmcObyHspZ0pImBTDATthq58kc
CIPQddPwYIuQ9hb1f2sBQw3IUV7QZ3OKadlE+ze6TEzrlQlcem1M4hpb2+xpzVVV
qHJKv/PQi3PUi134xo2cIsAdP62MThCymadvCIhYaeGlgu5xfme/bxpBLexhG28Z
N3PD5xml9rlGB6fRJjePMz8lwUJB9lmfx39Ha2bBAq300rxJ6q8ix/7WUicJKOw1
cNbh5dygAeob8aNFbuQnFCK5u5M5n9fE14SVQoJCtGkAQc7XoRx6unnZ7ks347M7
0LOaXPXJOa0ax3/CKxKDck7MvhX7+qOchJ8bLFTHrP4DVkeDaMU+dvXMVbQi+HJi
9G1J/0zxQH64hKM7TEJtqzQjrpvN0PnYa6fVKwONI81HksggaHqESui4Jvogj+EU
9SaNXsRWWsrzMxtBG4OIRdKSbIwOa3xTiyF7VdfNuTIJbfXi/71UOPxGaq8D0EIu
RV1Z4kefGMEQi65N6YGyMxRkzLNTSMkNtBxGDKGE8W2brZ7LWBrFCN+c8wT/NXh+
sntL1dmdyqbf4bC2BR3gfeh3+4Q2y/NtCCSUBiF5Vb1/3r8JNQfn91miISWOWNgp
6C6cWoc+iVH8oI8JdDi+i2HJOlSUYnY1DEhn4UpGAlnp4O9kARYGTZ9TG/vXx9hI
vs1wiqKvnaNRDP32z83zwB4Pm/Y0IqIyj3cXSQKYRHDG9maBtRQbPYsYZHWn6T/1
GfcH5Ke8HhTLS2CVB5ZCdmMY/e99/kJi0L57yW6tbno+9S002EvT6+box7vGwnzT
y598qpTVIhiuh6wzxDNv2kDu//r/cnON5VMPw3QktTFJ6e6dRZxclXVFZ4UXKJaL
31JcBW/r/HjIfxBZRTYINzmQ7aZqDP90RbwzwdFFVRMiEqygMukvkotgiw72S8Oi
2RS9lE/+P2SE5K+zvvNnVZtgojsaBRBwc9486Ib7uqMfLnL53rmSYbr6BV1fQAc1
/293f9ROCo4s6J6VQAbJ81XIuN793FaDT+pFIuKfle9NoWpqd1va/40qXDFbcx4J
m72wJweSf3mVk7FkgfNj+0t21z8bw/wazsF51/+nEBYSOfER8nYTFTfZBJhoPTr8
qpmRdzSBwgNbstk5BPH61MVqK3OYO5vWculMC18mzjlVFAbmnL48ic1u7hpY4VO/
C6FwN/fTglY3My0t3Yh5fXOhhTXhTj5QX53/aPMLTneLbYJs/tD9EcT1hS9mgE4s
fvGtYFqVIWHQ7R9mRd7dED+5jZ7kMcQxAWBQY9wwgk0DTprYJtfxXlPN7R8rqBkl
ZS1zOWbYDPHsLeIN7zM7MbuDHzgspOPZa5Kf8lzhQh/fdLNjM/qWX655HQz2ICf+
j1X2AmGgTR0ohoyU/bj34zC6/nEBwnyV21/KWzaIjvpM/nH8DPVL83MxIJfQOFFc
AZ01Bi8d1MR/4phaCbpeGBXb7e39ztLalsxjUiyI3nYnK6NMtod56+DTTTR/7rUp
hh5hJhWAdFHjIFt/oG2p03ySEoaTa5BaARkuz6CFEvEl4RnKbp+aNPAhfbFqNPgY
Lb88rQOPnjSSm/T/uzusXuYlAgQZZ4LRUdAukFQsZczMcpWWIgdsYMR/53NzaIVY
irpL3qbIu8vixaGm17jcmXTa0BLnBXWjthSkiLexXCO8xjQS6FPFo1p1UJlyYs8g
ri5ZNiv9OzLjD70HpsR9gCE0eJZWYARobo4QvmPOEMhcvKZW7aowAKlf7uS8aPtk
hicYYQkHNwS9pscXvklAVFg0LUpAQrspZI2y4onHWTPYxYHrvDAMsQz4DrfQN9HG
MnrLhHDdFghgVCgtzMwTLBEKZv7v3IBxWGhoLvzdlqSx4s11T5pODicCVNlDUtUr
KadTcfFNOVUHvxK1ve3958XS98/8iw6PcoHEOBWxgVkmjrI9O5/30RcO9XVIcUmK
XNOSHHiTdSy64Jmwugx+ydGIpQBTRw78yBvSEqoE9MtOZK6PbZLivG29aE4Xla57
AuUDBL18MPA8e7c1gpZ1Xy6YbAFORvLYAgIGd3hwWp78NwRpez1jgKUQisE9ivpm
JYgitz11trsi8+bJo3mjgZ42PY6EqaOS1hYbOwa1JZfz6lcHNHNA9sc3N3QHtEJY
fZydclq5y1j+qBo/6I+5eXUk7vwkRQrnlg+/zAsrwk1Nnw8EBMPN1YyYOmVd6r2d
LyX3Iv8hWbKdrpjaqlNyhKXW+a2Op22kki+PuPbc2nUGwxvdA1g3jvS6v0ngbM/X
QOFKTMEdSP8+xB4b8pHOCem6/yAmQ34OWD50Z+NB3cYhULEpf7TOwk2Uf9yn4uYY
fJHzrCSYCL07AoIK4biv0dtWuKD7uASfDKZC2ljBgguH7uV2KEMW56z+kxhCYewd
UDlhG1qlOeGLPTKHnwHkfvCOKQ1oeyB052DwZy7FoSrvsNvEFxLmKJ81rz1pSSmU
A7pOZmZChBKPtWgJsXzXl9DsDOcQO0APf2/uzCeXLr9FaR5/5NtekH/Rr34IyDUh
XVO6ymo17qfEv0OmPD0ZJT0T1xBBFiCd3VV5y/AqD7zFnaiVXlhUZu1Hzz/92LGU
Ev65Liy8sHW2uCJS/if/zNOWDmP21+bO/zoweWGoQWVdBIeaR4cEKCyNg84UvE7N
AF/5m7rmWcAFAXS19bcWJokddO0czokPTc9WeVAHYewEEopuxIR5ezqJZ1825ml9
Hr9w2+cQN67AMXPhhuWp/9G+5jynP7VzwCfw3IstK/O+WoUWUUGT6+WM+mNsGQDi
B1c0Pu7pBBXk8N5Hq5en/bEtw7S279wYXwsVQodrmP04CiR2p5VGqsA1VPE2Vfpj
XSamxoRZbX6PwgjrUM2kNzgYBcl+Qwkj1gbm+/LMVbC7h3/hmgZfbqx7g8QTu8sF
hlYoh/S7U3qx+44Oc6KDrJd3FBYMBGnsUpL++gOXvHsiUA0j2yeTuXRZOG1QkXQT
G8h95xlYxSCnMuiY6X/4JdbjRQ+Hj3s2h4Iz+KIl9hAZ1SqJ0wUX229ztPY+INGH
ae8ZhQicUC6L4oe9BotD3STIPACh+8ESz33OD7jnH/vZ99qBoh3dU6+KdSfiW3tH
LeC7z7He4T5KY0ZyOMa5mzvWG6tx/X926bFc8va8I52g/Hr+RMuRt7nXP+jMb21g
+tgu3xTKxB1lidggSPBpTyK6++AOorVcvE6UAZxmZyqLkAlmojq3he17miaIxe6u
dPWE80Jmg0dGyAa0Sp4YvrZBsZ8roUVgTy1MGk9wgeWBtfwgII+YQOXoY6m2meUP
VAic9jc76sXh6jP+AdMxFiJfOabsghesynIgvd6VEskCOempkDC+mSvMmSc/XnT+
f2ipmY/q6juvs+m+m5YyIslAe8TfgBkSRfJMaEwCMrhxBbQeorILXThg1HgOwIwv
GyNqrf32QyN9Wsz3N7pGQLMTVvmEH8hNb4fghVTSzgfkorQ0IxM9B4O1FOHBz8kB
ZgdwTr/4VibHZz3EcHpUfhGe51OGH4bfaUjV8T2YHs75Z9j9BmWfYPfsE6XWNGtm
b4Zs43O3Mw9PWmzdblKK6B8lcUfaXNM3CYISF5Ydn+EAPvRlTHqux3H2ksy5g5z5
m71aT3yPD4o1pAHsafsS02X+3s8Lg+TrplAf0ns3rpTvqvig4nl4iyrcFtgcI5W9
P+oWIQwqD0trI6hfKiWUzKszZdQegMGf6wUQhdhb3m5IN2pUbB7cWwvevoJnE5WJ
p2msRFxWoxPzHw+IL4Va63pu8y30n6A8diZoxBSwH4iO3BCqGeN2dRa1kvwhtA1k
C12KbIo9Dq1yQaNl5V/Vga0YgT8MZu8uSgKdvZygzi+/cWucjW1LOqmEiq50Rmt1
3oL0Rybw9X1ps7WjNSLopBcBjuD6IjkGjeHffFx8RPCK5R14dQEMnNVwWxUD/ezy
Idnld9VEoWQLzgE4hwjmJ7Y+fQCX2GzKYXswHV783QfLQj3J/gPpZQHkODDAGeKF
OBB2uVFIlnJh4hVC7WIw+h/AKZqouJVmqH13APqJZexT20HtlsmTlq3QlsS/siO4
HsTVQ3IVXD8rse/Yq3Mrfl6NVop2tHJF/v1DXnYwOwfxfmFUZkBpsfhJ2ICfoidr
qj/T1JOhGFx9oZPU5yNB8JpYfB8LYmBGMi4QkN4AULIA5jmM4KSqfzHZyiJqeLGy
fDTcB+j8UiyXv3P+XfGYe6AVw+qI9Y66bHXywDHJUds0YdzYr+zuwoJd0eWWl9Bo
VI/w8ly3TC7sneVGTAVUDT94NuTsJ0EZSdPYwNvBvcRAVc9ob6Koi7wxZpLq66B1
TqgjoOU/aKDzizBUP9a/Q8I0wCiKOP9r6CGFN98hh7ussdeI6SW56v1gV7nnPRJO
PuPObwUtGWH0AULDM/XeAWAq/LXJLwyV1uP2wET7F/o85+a86S4R+RZ8SWwwxUrL
lQdy2FPrE1jN7cz1fPPj5HN0ZOfB6QUPlJ/DUGOWWq1G9KF5z0YOyYuZl7vzTjp3
R/u2QuAVXx/VZkpuhMXGjzFCAy7X6jz3inWpX4aAjNtu3QwSPaZyyxajKrN5RyU+
Y85YVu+dMdw/4YDjFGPFbhiMSfe0BgykP+vnpNOz4c95NKanZkUvGS1zCBNyAQa7
mGcDhqbghI+/57nWWAM+jCbvCdN27BXjKItWiLmitUEDjYbN+9pjtVxN4aD98qcg
rLVl9Coj9T8VkfqnRFSBVwfYaEXLrBSOvK4Xr/gGP3CdFsuZFOA+xiABgC11nkd2
UC/88kyXqPtW8OvY9s/XRzOOy+kJgsIai66uFOzZ3ylCDVGgTEG49OJlagBvoCeV
3iDVNj5jYt2lRsDRV5T4OaEnsuTf6KAG19oSwvW0Nsy9t6mhOgv8IR5lWNJtEsO1
B+QdaoQyNsaY8zSehq3qyXmksF7x6QEuP1hFlEcCj0UhPidSGyVhSJ8F5g5QRYp6
1vWbRpX03QW6ps6vUNmrWMUKzKzc520mEu9oCvGizZ1wLCyRscPRoXAyizSDcBE1
pUsN6A/QGibuegfw39Pl4P8hTTqp+cj0wFh8/4vZYkVynqI8sjRhmnuo1vNx5V+j
Ke2hhj1tDOOqCa4q4PBPN8P47d2pSNQtHIK8Pt9LHQwcHstozCDHd2L+LdORRkzI
DXN1hXcvECUqOXxdz2RHnFhvLZqW6BWaJ6qo/+mhe8BqOPi7ufkZsockvaeVLFvA
ZZiJA1Yt8gzngiV9W75arJ20C9FBWhqDfbL79IjD7rDUSRO00eW0S1rYmD+Ze103
8gDeKY1+BbMdLpphZAK5dZRoHiHqJlbCY08uswH7OJ4J+RdNPwaCdtciwq8mL55H
B2eDl0ODhzvGpcGsfkAX1aT1TXZh1r7AvLM/0YIIU+ldUEBFuyMMAYd/5bi1ibo2
AFa+y81+YQD/5vWpHTs3s0B3TZW2MSzZxSg5gCUUnA7eAdQWlDaz8QYHns08Zye6
s+J2/iaOjYkiNIysYz7buPEHf3fhg5eXBs2b6eBNtnOHPQRrtiZvKXJ4Bekg8/R4
Z8bLKpFv8ZWCglPGCUHBLTP22tHpOeAVq3Uka6UPVaH2Fp4diaeS2HHf9Wm34nYK
m64f3bZeWf2haC3pRdL59+R8jGAlv8IhYm0VSKk3gZNHtb043dXYOabYguV2OFuz
yNNN+LgmSYus7xgPjxD4LGgdY/HAnhEP5YdzuTHgTIvLfFj/TI7f1H+LjUc03g9E
8d/cj1S8NQLCeyP5s0ktuwg6l5JFApcKTj7xlwm7SYH9wwYKT2TCpTs02MA/HwSM
BkQ8YYvM5WuTnkA5HXhBa0yj+FFdC27tgHNsrfycAF7hoqCJFFA9XO4abqQdhTLI
DcsXC5RnRQ5yaYiZxEIe0rRqLnzZEGDMWV4YqcuLKuInx8GjS2/X7Sn3Rx6QL4rz
sgEXYv4UOySoo1RUmTGl4QvPyuJo8l29TDU1mNOqoPxPdkl6wV/vHlhfo39uQofG
QKVJ+GJRrbFj/8qWw78Vce6U10YHbGVI4k6cSPDcvux4OgmrLXSIesWEepV4f/XN
2oVC3+NJ67GD/bo+GZcRLdghQTPhlg1HkVZdE86jqIhqgu7hUBv+hcQ8SV96vbTm
kjU/bpREaTDDqG0vzjDTixilwD1rkZuQobgs0WBQuzLIyfTXf0IjwAZw5tgWUuTB
MO1c3ZwfMZa7dSmSbcBoYZ/oQx2k73tnYPwYk81D3DQKBZOZ7eybAv0feHVCuLp0
RjEw2yABRD657gTSzMn6vxBbsfMqqUgAVGCc3FWCpL8s2tUC5sGwgGYKX1AxFkc2
MbLOY6DfYuu75zZKcY3UTlxX+ixZ1UUnFhBG2bO30cDM/O56p+ihckVZiiW89Zj4
4cZ7oaZvA2QIMewhmxS9uHQzQxIjS3IEmsZCj+s501G38S0309omDRbhsLm+AWkc
j9+jL6Utx2z4JsKWELuXB+Bo8zcN7S/5wMpeFu0kQFH19t1/5XwT2GIrcOljd5mF
+RoJETLav7ymbeAYRGmGsEG5UjEVnGIQQ9sfj6n0E7l/N1l2yafBNqv3inXuyVZR
Rq2QBUyT4zUbKc6E/fCncSr77V8arsdqGfzu1aUzbT+1Au29Qq/XQq4N+pc409cu
ifxvUvKsW4Vh/Ea184wBxSFDGPGsSe849vM/xIhwqqjJ2hJorW1UqDq/irE78wmR
2JB44eNR0QAZWYVr6rwuBhub54H+i00pZphHKydgUdJ20XSye8rfViurd/gBORUP
0zNOvH5sN9u6cCPC6kmidkr78eVuJ3kTylSHQP8bZDiDyrrrDCfbveZmpQRy4qgf
GZ0sk/zFU7+sVkiZZ5EY8X1lS9f9jCWt1gaaKR3Fd44NQS8wn+2q083OCapYc+qg
Y5tnzz0c1Dp1NtfdmaVfx7O7TM5Rwohw/8YQV+fUSYSGK1wdkhDkAYITFkitowv3
C4HsZue3o7y7xQoymirCKLxHfSmbeqgBD3MFi7qBGxmcsBvp+1rz7/0DDdIVeouU
6ECHkD7/cfpVr7ZRnb71j9EQFlXK0zPXOMbjM/hrEA4lw+PBXcYtjbJIGuWehMBx
bexBl1E+PiU8mmPAliQLPKZNp/ZFTM8u9hIYSNoIvARiMWvEgdd7w3GIyeRmXx1Z
JBuXn9/SoqvlP9SvIMZ6fG3jyeosAuC77l5tjibnkOxbHRa5ftC0kem3jQa+CNfC
+rIg9nCDIFEK3zNMMsXfR7IC8sqTm7l+52ot8IwphtWtV8i+spHGc0PiePm9opCT
yPLdCriQXfLCGnlAYjNMoOgwlLfkTGariQKSwHe4Hf3SpLd5tfsmArQwH3eQTuK3
8Cas1F9Nvt8lp04y38J98MIQNSM8PsQ356nwWfvzpaVr1Tu0MLj/GZmb7cQxTMvu
YkxU+OfqmvVXBwGR3KS/OFgZnSJB+Kn/t5nVSmJ4NI0sa0hYu2Gm0CNSL06OX0NI
Kk/rF2xvxp0Q5rWwS+a/7af2CJforgvx1pwRd3+uHLbfG3rnasTux9YbyGh8Bhhe
zDPLTW/P9qGaxMJesHB1qSm0KaJCmgi7gbcHoYbSfTzvsq/p42Zz87T3W5+wKOYP
OlfYf9Vk7jiq4sNkf0+M60AA+YzogcG2hB+zj2P1/bE+ZTB+DNFCKpTVayrTpsL9
LUjRxzM/vFQsP7xQkInE3Km1yJB45MKCTyzAlE4N/cJIo64jQx3WQXBzfoCLFtnh
c0KOl6qOhGepbUudgp0hKTi3K1BIOA91c3ufA1mwlSD6PLrc02n0pnXefZKuMtEW
tb1ux7GVHigy6DGXkyLj/7kIDM2hXKwA+46Fj5p6FgGiRAEnUFpEFiaVdhuVG4Sk
tmlejUdCX+ULwbOdQYmnqRB9TT+dP4b8fKLxHjVr6N8jwAvg6Igz1MrvtzWBmuzq
jIVb8SzHwrYjGXEN2gpU3MIWOVAYN6JxpH8OYIq7pPZhsxzNpDbR3El/GxZy9wg8
2ChRzYfDTM2CHasJuO1vwuG2l8Ey3JEfX6g+LiqxLT5bRqP3lnH/n/rZ0wO3gHDA
MNKwBzE7sgIskmAwAbDNcLF7nevFohtqrsLPxOWldmwKe8gaool19c9Pmn9h5ihM
0xpRzommt5RX6hg1Zo2cvBoFXSuGHUSvD1n5dxB+cK2W442jw7+Q5IBkQ1UH/P6X
zvml7GhJ/nu5EGmfCjfh7bbjMzGm74XZ1Noa4VjLdXrWQuLSa4n+YqkpN7JmlUv4
B3X8tJ2r/XTNRVrz4NU3SxyMOXLCRovD61Zi99MvzA4byGoV3I4LJctS7dZrgZ5E
iCLOAIcJbL4vhNrwIqZOLRB+EPffuc6mcBIcVAEUshR3FtTyBOlrDUE1zXiVVFYs
t18zNIuyijAQfk3BWoVEKV5zNCSskHCOVaQzs/y1+qByTdYnTvQ4z8XHCrbVKpbR
gxPUULnI3zF80CJDYe6wlkpa5HV5JgVXBkGSs6mA/BowfmmYGYw5ogwGx1YAsQY4
rrFrHWr8Cg1ucGgAYZ7fyP1Ojb9v115Lc5G+qlKJbJ41f5UNX0DuI/lQN5jRiNoK
Zcu3g77v3safnHqRZFM8xrBRL6fH3s7mDi8O9QDw94nr+zF8+NvW5Xqmh6i7QRcG
eeUjKV2HlYSFjLBQhP84koklreD0YnMH6/5Pzjqn+cqj8HUXOjiXGKd1p+icqF/7
7CRDxWEwqXsR7nKJ6tbGgEs7qlVusZcnCSXwEP8J6jjHelciEyxjVZCoSenrigVI
TlkYdE9zKDoQDnWahtdoAGX4buCIjwiSKwdyhYMXhzprFVeUrLk4peXHnP2J6ZdV
YJ8noorNWhOCerzMC6WlShakJh+Rugwtuoxe657df91BGTyrBr6pbWobRq8S5sec
V/N4E1UcBPIhsO6GuY2EU092wIQtGdgOID15pw9x1XwrZiTxxWlKS3El0ffj6Ahg
ZU3nm5A+UhwlLM5R7Gxm/U0zxyUxegArhjiAKHFY5WEo6I4JS+2Tx1UVy4xt6dT/
6MLGmFzOaitE3tLUV6IGvGQtyoRaj+o1AXnfIxDBdIArYw0IO2cOqeXtX4tZYjTy
x9+wOnPQa8i0407WsYjz/gg0BmoVh4Zm54lZHZ18Zxjg17az+C+ySabZ6gSG0bjZ
ogvNiYW0zT1eOyX9I0q6obVcM9l5ThLsIpoza2Ru/QHg+dZQD9+E7nbgwBeiYoZq
MWfqLVe4qK8U1xGN9OfFKqX9/VdkK1r2JcUFdUS0AOBlOzZ+NFI5YyEoKS6DwY82
azT/dW8NRGVCJbl+2QsRF40p14HYy+k6P//7hIHDjxK6P5sjchqM2TkrBw7hEf7e
sas9Dm+u0GH5/mMfXGamVGoUnVbLcGrDJXBhFlnO5yZArr7q0FX7+a0C59OHDXv6
ptRdPnWsnZocVjwkUtkHWEme10KxTktYL8paap7SQglJRrLJIdvmL2L8tQs+z+Gz
8EeZuz87ZT+AMbZG2H7/igYz+SSfMfGKQsrZ1sxA5LOFItur4dSaMorwy4GqhI69
K8+wBuzQTqTgTj4YT3D4tVX9FnUjpc3kwEACJIufJsg0v9FcAImqDyv6VSejfT25
mDkLx55j3/5RtX3vY0e5fjfgPQJGOFVIgRVuz+2zFngGrKCO+xr2x8zNLKexvAjm
IFzx+LrQL+9Rqyqj3mQogGCjBtmfSG95HkJ4YnoJmDNeMH97XUTTpAmK3pHm4H8t
FBtGqd99FWebyaZhqDlJJWGO+y3xlHrzjSA8SbQzrItqRohaxnIdVrK1F4IJPu7O
j8yPU7JNBD4tjzvSE3X5e5PPpVmTTB/WkUQ9r5U4olT3DiEqHRct0Iwo3/V2kiI6
OEU1zQvGKk2VDvh8ybilK6V27EfHNYbd7UWlyBN/Rv5bVJdgmRTOWY7LFmU/PckV
VuUVpV65YMEtS/FIXxSpIkQNyXQsGY/vfdp/TyVfAADY7n5ak1rWng7hEMlyvql3
ABRqCOhH0kbXdAjxYE2nibKMnYm2353+9AUuK1dU7q6a7S5L9Rv579p+VOejTZdK
ifBeIomun+p1mUvKdizdY/iFhI12fmanAwKHFBB+FYp/hwZtAYs94vHiWwH6fQnt
Sjlp+pk/mr+p2DsmgPuw6e7N9bZS4Agb/RDPrm6aOa+L5Rcwel3SOAocmCeqHZlC
dqfF6bq0Gy+//kG221zfPIdjpDe6q0/7wJHttVxq/5QliyxKPu6tdMHj17iT8NeG
fCQPHx1F3nkPqnvNac6eMhuo6/bhVEZCdEouDJFhFvBmo6IVmMAK59wO/6kXbNfq
KGSLGP9TwzlnO3s0AEMTg2Ts1lQHwXbGvZAiVGjBo0zBqycuI1273I/X1/tjfs97
xKWNs+UJGZ/wCs0/4YQY2F6U1e2DhvSsqtdBk6aabAXZhzmbi4AxA1vXkRRHlVMv
pBbJG2HHy0PXvBJsJAqSV5RE7IuPg1U4/oCV94ZuYRPIvqu8741uVhiUG5XHYZZl
TC8U8GnLTCTXdAHGAR4qFXhFVlJoWroqil12Sc5gEijnXPfs7tNDcR5flVdXJdrg
gV8ZX34HBq9H8AxAD2hwxQOJ2IOnZ0MWdGJaOuaV69iwvl615PhFCwzkdPZiOpid
my1zPnoW1E/AnxedDSYN2Z9dLrn+k5M5AIvUdUkFU0sHpbLfwiL/0ZqGG1dneJrr
x0o62Ucc0LEFlgtFWgo44qZmbJy3UMJOlJQJ80Q1R0E1zV3EqZAFPqJOEy1o65/N
0XXGeK6gANbKHCNnJVw+Y2GVBrbVNNrFRAY+jL6deGXB8HndzGr8xySOblEJ00ss
gOz7djcfPVWjj+g8acYSbsxwkCk+s36n1GLBRi1/9fc7G5pxpq05GEWEvGXLmkzj
NJcYPWjwxAgnTdBTI3/hs8WJn1VA4bXnC+OCMa7wHcT8pkZuutRlTAh5vzfMTavI
1ZGXVhZdy/xcNurfbI0Nf3606l2LkrWQW7G3gveIA789DNmGw2YIe9ohySLDTCEQ
RyFF0MMTsOHhlxFYpvKwibjwTWbvMPbTMTD2mqZJ1Y0Mf7/Vkz2JrUhi2jDA2/a/
XqcJ5+FL4w+M5j24RiwwIet+O/a8w0yzBghtUREjgFGCZGHqgchweSG2BRs/Gwrl
WTcCDcRA+i3t5raTAB7cIUKr1uJrRhxP9zCxoPRxUmviYRYHNvil9MGxFZJS3ymc
IGyOOw0G0zNDY2iFv+xGjYUD45d7nAienTMhVwfeXdfugAgYayyz8BTpfmqPqyBH
5F+ZkKEqZ+YT7kfwwQiSKY4EXgi4qKBlcycHvGOJxiamNO+4ECIvd/4hTxygVCmG
TJKbXa/t9OvzPVbdMC6Hf4nmMhAOo+5KtRj9VBK8Yhmi9LC5mAWL51ZWRVlVvyeN
UzULzkU/bqs2fVr1r8J+kgmr2Atq/ThncVFdC8DcuR0dityTz0HC3z3Ep1L3RDKx
1XLE2xo9GQx7z1t9rlLSzSkLKzmsXw2DQ2bs0CYnUCFx+X7LGu33keYYcuoOenIg
zPwsye88+UqWMd+2jkhbvEMpaLb4g56+FlJ9P1fIxRJ2ulBx/pTRqvvapEMPtXO9
fu3VI7AQkCv19zRzz3ayogHtB+vYVo+f2pWxI6qGJwglrMKLfDjvlF+IRty9mQWk
8FYOsW/uDdnDDWxLVPsDq9ISsM07nCbMLRJ+lLnixejcyYUwH9Bk/ZUYhIlocfi/
xy2il90tUSs7DRr/tfRF70YVmlO0j285cJ+SzniTHWt7WkbxQHtsMMgab6jhpJId
Xg5eKqjQ4ug8tSi3C2KFLge+Zhrqrs+RV2dSdi87FFwfCqPrwvM07HjCjBr1lt4t
BKHTxRIuFPF32v5x+f7esq/b/lE5j61hAl80z9bQA3hlOdlMQhgvim+agX9p6BAc
q7a+rWRUuJP5eO5aHruRiNS7Rr9Jd/eabQY08JUqUmV7Nkplx/AHiO9M9CUBda+t
wy8+0b6Y1qwX2OPPzc3srTjU+ZPD+LB+2ohiwZ8oV70ruXXHRcyDFQTo4WHnPoa2
z/JOF9xYX36BBDdAwXh2rXMsqb00GXiBaj5wNXEjYVOtdRw0g80UstwhWy/wCSyw
4LrN9hmFS3ij3p86qEkwBhtAcwa8dHxTu5cuoZ5rL1GCK8A3LiCffx6UasfaZiDJ
jSLauNT9x+aohuR4V+MuwplvkY+foFfbtg+236K8/7UnKt5jDiVHK014yhDHwrnf
K9nl0aqiP8uVTlWHXCxGkGJKYjDTtssHBiN+haYV3jU9Xi5xj8Zv7FfY+wNVvNVU
Y2DyTODwpqQd1f8tFGgBRwr0hMtKPJ2x7e9n4qN19OZ1bmEpET7+FzJsUb4k3iuG
TFQ8Vws87xALTK0VZlXhUGMzjfcY8T+sXXhr4gK24mywL/lLskKwQMOtysC/Kj46
88Nl3U+AWzZ10H2kvtx6oyp5nimRgdiDbzOGr/0Y1LaP9eoR/5ogv3GcYT+Hodcu
IX3n0xNLE+x6eUDZmfX7UbXoHvcT8ueGjTjONDxiBMV3s3yBwNSlCfYfd7E3jZEe
qp94062bq4nWMmohFWzuHqCW74LJdZ1BprxNuwKmUjLoPPy+063jXy61/5tlwIyg
IT/t73FO67URLfJ2QHKjfK9n6jqfXGzQTePyyTeSr80PvbbMxe+rUfV64nDpj0Fw
zomZ3SjoA3VFOdfJeGtrUQCgDSk5PvcVrEHS8k/SP7eY837r2zKFL4J818i7IIhM
+kaQC7zj8k0Zg40yY23RG4of4C7q4h374BJZZpU5RGWp+9WiCiEjHuOMqTPuJ7mP
dR01SMlBEXLuc/pLEzkkZssAsB95pudWPTPLrVKXSmgvu4Ayz/x0v6/Yb+hgocn8
ewzRU3Y8bCpZo68cNx12rreWV1iz1q0M7RtFb1CWEg1gJckPNtcDZyawJPcB5j/G
2GTL+rOIC0f9qhU0UKaryYWtvwRcsFoJZ2aEiz/JS1T9wDCO026oazGYOO0JQjp7
XWj3gemYzTr2jmF0n13ptnHgWQX/ePgWh+Aw+6AybmPY/jAkCFTmyuYjl1TKByOC
9cXEEmhORunJ0yRpeN12CcuIDkXklph1qbt+tqwnuvF8fIeEY5N8PhVRYryfBrfh
+NAEi+NZCGY/ZnkYPWbCoEkufUFOA0wPbKLCic7rdiJshoQT7yE5s54Huti/Hh4T
iIo0+pN6ju6p4hFFbmQqzHL7ApwzlG/uZaAn7HrVKHdA0qI24Mwala1qBZDOP+ih
z2WpbXVGlQJHlk7KpJ8buQ9HA5934kzennxagEyhG0Y8r6g6sRSWj0bTEAyKuQro
q1KHP/RaMW6WEPbvY+QDcqLZLn7xFKWOYIMYaV/+NJjBjmvNFFhG270HwcccoJDX
nL2KuXRrwaUjR96MVZk7NDyUuZsZHH39q+I0WhZrIXQ4OgVI5XEaGRHJBMH+ROn5
bJn+ty6rzYJVPCI5s532EYbpHMHyoMnuT9DJ3MVXnZuiQ0u+XZ64eEgKPGvjyX+d
xIQlYezCI1MzwVsuJfT4E4jdcDFdZRro9EXEM6nE/bL9zOJnLyS9j7/AMr6TPGnD
zFJN2uPvyhp2WmwefGG/I8ILWD0ZmXZg8L8vD4C3c0HYAV3mZsi1c1QocdweGbQN
b+XjQ6UyHU2b6cPWuiNPm/Ui62K9WTMYZV7049qRZscxgtOp12OvYOkfJE+kwQRd
dR61Q7iey5dc/YNSmjLEJkSzrTa9lZ9dpTZM9MTmJMaBfJH0PkPoJvg9ZIHvHuwI
2wg+g1I/nyyZDQ5KOylMfhkFCy6jgE3ie40wK7VnyJSYRSjyWs73HPSpzQSMh41Z
z4pabWlCIepr8U71fHINWw1L3uZzJh1a0SQjbcAiOWt5i2IyI+z7IgvqGxUHiGsA
M9ldHoL4cZJKBQP3NKvf1P/3/WYDiPqFio7WNPtYTLjqD+cDw3MFf9JqkaAb+uui
vprzLn8jgNwW//sBp8WBG2albInbb0rzPqaVurRYEqs+CHXOmH/OhSwExlqYBSBQ
MgjD2gCh2Z7Et1EKbGakdt1lYrNQAFbAblxdgFcI2RPvnNREMA+y5ZIdBVSWOm4o
Y7kkavwUUdzw4oQi2yW5dyyWINi+D9pf6VMiKprfmsoG5KBBYRHrq/uAoFH3J4+6
MXtpkb/IK4ms4RI1lx7vW/44ess6aIKO+SmfRslMQIYJUZ7mDHZGgcyZMQpISal5
oGN3o/Bd+Geianrqhl4QD8gvsVXJkRac+/7j5IXmo0hhkQi5pRC/5sIZSt2kqTTj
R+YE3y0+eYAWX7GirEY8YhAdqVauUyvQbG9lNNO8uy69rctUki342fDUGVsccu3w
vokM4grR6f8no2AtCFusKTfyLzR/ScNW+scOqxSsOHieQAURjAFLu0GKlf6TwmG1
pV7hPN4hdrbrXeDm1Ijuojf6DpLfxRU882rmYH6lScHiU3qIaV7m4ghs/R5VN7sM
glMOQ8Kk8Ep4xpAbGjToSgL08BN4hKVu5uHF1U5SCi8pbuOD5pe6PQLC7MA/twEg
UftYlVrZslEvb/UBYYUmVEv4FwryhTMZtIBgMf/Cx7b8akDaEUWhRSAGhIj2+8qL
SPXjvvIlrVXPYoiL0/1VyeLp8viSy+sWiUJwCv0z3xbsqPEUA2fr9etVZ3t1d5AO
ulzlMoqtguZcxloDCFZETa+pjRYCCxjBhKSaWSEfP1uIAskKTQw+NVSkTWQT/l2K
m5ymHk3D2jCsS/paHFbgHCMQRcoUM3nguiD2FQFQKXePAwPw5b8bj5u7UjEybUiN
jOEz+h6LbnFS2Sk9AF0Vzmw1K+S1RUXGhvULD335Ea91102ay5osUyWtPZr2OYVt
OCXyVU4RvfLnnmFgkQBqzKg2JZkuZY4Q1co0qYUxzv0qfQo8Cex//KuLx+sFARIq
IRacNjH2R5ZCdh7HkoaE5lvVDGxA9nn4Elvr7bblZYpIKrjwyeD0slSrCui2wm/c
WKE2ecLlymZsR7MDKYXo9OapJeI/lVfR8Cld6f7N0dltVJv7haMyzoEAfp22ZyaA
t+ehlHUoJ5m3D8EWr2/jBDoosS7fFGZIUfFFFjwu9Kxpll23K/Mai9BwpU8nJF6b
F1Mtbt2kkcltELncG8F7kNwPVOv51tfDmhz+MpF/PHhdQkjZ+4d2JXGlKUZB9KJu
3pXDxRlG2jb7Rczj41Qw8imKH0pWarZ7YsvoGZpQ4xJ9uaeAVnSatYn4IzhafPnn
qZsU3ZF7d47oUy+5fdUa3S7b/KSVUa0JJUNyPjhVPrW98QaFQFBCpEmD75RmNy5s
kw4+qhejSVMImJr0Tbx88ks+OLZDofy6sGePjqoamBc8RFjghhEjquiv2umw/kVC
o7lw0qNazXFStAlpwGqXg9VMMbGO2UbVT8Dlzb1wec8zNrgC8qtDOFH4/kb8X2VU
4o6fyAianhQzYz3MVkEIZSZ1lBFEFnYKu2G3yQGIS0cFp9++HLs7LozDxYP4PWqm
YOsV/TpYkE4tegb+wEAlikyV/ztFaVuFyojLUNp6WTNxhbdymyDT1IEcEf8W2Uum
E/kFXqYJZg6+usbPWMRPIt6lKgr1CjMZmBKGXIOxxz8mLHOLJMVezyk6n43BPUYQ
Qt1oc4Wkt+BnI0m9qSk41FBWWmQkUqknQGpVtL5g3oFgM2C1BZTM3eYc5FeoPFAw
HKHY1InYqhdjUatiyUXCEU7w5s9Hp3dRheqB573ZJjDbYcK1DuJGWrMJAemOxJeH
TV/55hnvTka2g/Jw8zIYMtVXdP1EYDBHX/05EZNCEebMro1lzw9GI+CibbtJvd+d
HW8U/uUNYnUMAp3ZTNLlvqopyNG70Qh/poOU5Ah4uk/9n/nQnjCspurhjnPyLSLP
L70vwFo19FdlD3Cbu7z0f55HnHdFiihs18IiyCF5yvsXP6xgRj8qVd/y6rF3LiDZ
oN1rvRCpMquryN1Y2FNE/1evixUR5pbF9RpwjLGKGZ5pYGdtDlyRUbr+9H1CoeeP
4jOGKVWhf161+L9P8f68nET+irGvWCU+qM6hJCaK7p4vNBMjGwlv+m/VMk8Cs1SE
nVAYLdZLo+B7PHadQ93tXmUCgmecGxPbhjLIBwwpFcuuM5dxIRxw8JcsLj/5XM37
PUWkcIahxdvhXDkKrXw7Iv6D8b/B3NxBz9WGZ4s++tFNxU7mhq2a6vFOFpTASzJR
EmdoYplmx5OuV/8e7SZgXnEbxiOvR1nW7HTtA7zvUk7uoQ1KIVVLy0XeECuiCEL+
/tJETIbCliDwLZsQjZkji0LTriVlJVDTspC3VcW8bVVDGrienJAqF6VH2unUvfts
yY1AOk5+naIOSY32jMviqZlpzhxHv90ofZB8+xFWj28txADsilxvEBiM5U0lPdyd
zgIXx7rVG/XkGPAkZ774OwLjamAh4c+FP6EVjwCAa6J41PgH58fP5mT/MATqOKW3
quTWC6B2W379MaGpkfvZqAm60qWiQ2PCZj0WHj9Rbn09kJRXxOY1n4130hFESWzY
QxMydh4Uw+FeI+7fz3swA0eb/CIfdaBXX5q7NIHKiy9bMgTevGWE2Ia5iTV6n7dk
8pPFVUUZgpWEyGHF/ieB9xO0APlusy+puNWRV92bgHZ4lcmAI93crxG7OFCSlkN7
tU6JvGUcbXOjLH+Zc3FESO2WWHChf7r+Q/Fluac271ssSSAYzss6lDPxydsuBOAN
m5jCQFgypz1XOHsdZO6sdqG/cDxhb22ohNF0preUhVYqTb4WbGFmizAnu3Yl7/TY
ZYf9B3vBKL+oQmseiA0DgSLAT+BcY9x511bI7apmmIatXpvyzQ5hKXHCmKYFk3bo
Gr9m5dSgYFl1QXRPbL+84ZV3iqN97FYlIcTR49o0tROA14CK2rj5Lw7DE2aTYbgK
ZNfT+2BhzcnEnwnlSnuDAi40vPuLtmMSAInxAasblFleTDvzTtAz4peyD7B4SYyC
OEfnFZMz0P1zFmX06s89u3wyOMF2Hml5oGjoxMD+OAsWwc6bp8+L36fo/lSbo9ny
V1P2Si+yNPmpPbEUCxrFkfoAcZU8Xm+3BX+1ptavj4hvGSDudYko9fUfV/zXlrpG
QpYo5QDe8Aohq7t1CkAR3dBiFkUZ3IKmNqW3NW5YoP/cNxR8xuf1b5OGCeFGRuSf
0TMXwc6AMvQ3ZLH8FmNmmlD7D/ESGDATSnFHXoOzZ5QMhI2PDkhlsZbVZubpn3JS
uugnHcLLT6ZG0aedoKnzm+CBl2hO6hxImh1bca+YIc+lvyBC+ZTZXJuLXdbSR3iU
3f4CE3GnwlYKRtulvK6Xs8bN+PIMdIu2HkWZKACjuNRC/lAe2yQ85r6waK5OUFK7
Zwyjr7Md/muZR6w00MSpAb20ywaeRYKhR9YpZxsKYr6tFZHMxPdVGCBBdAKDAYBI
VbJYhYOJ9qOIW/aUjeRy2zHbFt397VgHuwwik2NAcoNIPXsQA5FfqY619zMQbTBd
VmFrJhaKuMTg1Hmr/uSgXq0iIuvpp5yKlEu1C3hC2xw8YHYYIj1CoTfaEB5Vgtpj
xRB9XpwnqBy+K3xWptOSI5JkeeJ6RI7q0r0o2EIeOkTE+axnbc+5pxQ9BeNpJ2TS
L1Ol4to9dU/LrkuYXJ+UpTHSrKI1+/cSaOJ1v1SCLLNM5a3L4J3CKmUAA7kK38Pk
39HFWe+k0fCI4urfqjIter/yVcuVXNvGQh8+TRwlWcpLcTE+bN5cnRWMrMmcnCvL
1a6FSdv+tJYMs9iOgoPf+qbPSsmjoTVYjUgUNS0iRu4i20H9ROu/NI8p1EEhsW8G
Jqn9uEm9pjf0/r4E6eBQngBi/mlhc6feABknEK9/zV0xs+w12IegOtyTX6mzLFwT
5FjraAQKPBfbq7gX/P4tqZhMswpd53FFZ0jSVlLgHJJ2Jl48qHrn+PDmHQxkxyzh
EKw7ygq6E/1fE+tr0OClKtvI1U/VAIww1F1n+z4dlU2/0QUpsjWRB32biCDiIq0A
e30kSERbXlK3PuW2LYA0ofGsXpDlrkF1V6a3vDghqBljYBrYA1DVSEwFIlNIomkV
qyKihIx/6DYqyWaYh7KQRkmp/6uYVwUWXqyk75ELT0evx+q81it4KkIFGmuXEyRV
L1qG27/SHHQr9o3gSFlFIpDwtoyecZp7JIdvo0nVE3CKp/RMSK1Bidl8XoHjjUsn
EAgQbJ5uMzPVySVAYhe+vnWciBmJOEB1wILYagAKn3kQUabwQJRGCbJ+70onmVAz
mQWhNfsnN6Tk7HidIGSPrrv2+gh/ksDrz2A316ZfTq38PbGvxbVTJlyzSj2QqA6j
F7uMEskVoHSpE9DTqYGTzZQu2FAnk9TNSqcRI++LeZehg9+Pf3hjS6pSdUzhfGRy
RNtI9npjnninl/y/ZpqeBGGdbLZtg1Sm2muhs2geqW8Gwym007fCSF91RVlDfbx/
9MclZBXXFScZI4xN52C2wCCGVj45SbVTBHD3Aq+K4IpGVRkU289/6VBf552QImm4
nmAngix8Y85MKOIiyAQebYz6H9rA3yaCodmI9DmsTskin6ZxOsQx44cS/MJ8rr3r
Fg5VNpeHA7CVqjgSJorSoLFUPBfxG8SfIBoi5uOOLXpEO6q24YswBHzw5yy21/V9
4LbLJ5tVBUkEUzIqgwPrDgHscSMt4MFZ4jZIpMps0Ln1bahzYA8ij0qELOZ6PICZ
viS7c8KUDj44RiWatgesbO90bE3vglaVo0SwHobP5Dl36/DyPX8UXF1JNJB8fAuY
QD8WttqmK+ucnUHdPvzomD0UGXBHfs7J7pvgPG1csFIZV3tZyufZr1ah7Gw/FxsP
YlFgiw5daDaGiHGyNeqjx+uCFrELhw1VuBPI3GJlq9GOw7s8oa1DW24OGCPdaMYE
JWVZ0SlVtcRnjm60PuR8SZHL0oJUR5p42jkUba755IaeeIEfOSzk0m7qtD5Cw5FK
pPcb600Y0rAQHm2WjzzdzP16Hkp78aycS3JmGQyWm20CQx0APUif/vx/QIWkuRbj
N75xJct3rCXdra6Lk1RiqGQwun/ZVq4hhnR6TpN5O5PeWH7AEVLf02Y6+pRxwx5N
Tdm1UbhREG1hmZdmeTPjfjkRehb5xXtz/IevZwUKncm6kfhPl6VLY8oAjmckC4u8
W+oqUSTGYc9GLX7Cv+2LR0O65j5MR1WngryBovzupC1KeQXlBpfcOVtnV/AwkchK
JdX0Yx5JrwGGFIEkWDzy2GKhdK2ySKrv2bF1WEq3XChk297A6iTKxCxBJhxjy5H1
8nV+D1zzNXJtzDgKkxOed0mziUNzyBGFWgG3dZ1enf0gMO/Yolwn2Yo6OwrcveMo
2+UFhe3QFcOoLYxvob5+4eGbbupVQdg33uC7Jkb/78fSwpQSKKeNDx/R2cCEHTfl
AhRqz0kHUuWV3+0SNuRB3lRm1fdE9OGbedota6Rqbvh0F9Ml2EREePC4WxOeTM7Q
hWcFGxhJEWsmI9JSeQzOJGYyzZlcWyltyeydsbqceC5/nZW0YWaveQmYnrPBR137
sOmIMuJ/UN0tCJ4MlwPq6k9AUUN7bdrY828ZKodP0OK5boDJMX1hmlPnKSoBt3iZ
ybcd5l43P/1urhqwiO9FY5A+6XY+tyIwOaeVR5Bdbfn5TytV8fhG/qytAJvOFePk
4qJ3gPNyEaSXmFYt/KOHAGfEfJhhqMH/QFi677Byb9iuck1iQcUScbZIKsyAmW9D
Ii+47IDVwOhUKLFJqbHoTfHyh4w+u/njRBCruxyUQT8f1l9lY+LySQc9IF2vrMrY
+J0gOrQjrdQq8wtDXk5rp1NTIoizM+yTtOqK0EBaHnyasgY8Fjms54Kuahm05W3N
2xj4FvDoBPw6pO/ykHmzhInBTuhB/yTP6i94wu2wYaVtRoNp1zd/TnV1yoAPOGaM
xxCM7WEu6Dc/9oO/gxqHVZLI67IENTEVqODH4yD0olqItS7MwJ4dwI1htgiCm/ez
UEsQxqosOrAzL5GVNEgIet3FZ1XHpq7GEUKhB6N6NORPIEJJEO6IUFbCjH7QmAb6
PlKMoLHkj8icYYJx2x6fO7ljOTcTWpKa3tJ1nRkNNALg1xmJDZ1RMqeEDk7y+LiS
2y21TGf92acjNwUtU24fazLg+dFKsGYl4jVrMYeU8aCqya0y97IbdSVtkKr5IHwm
lz59vMhP+Q/G389yc/Xo4q0QrgzkNf+bIa7BycBzcgzs7/72xaDt+P8+gRkn2An6
ZdgDPp4NCYPn9oalR0y5T0aBRcR0atiJO+meEjvyRfy2ldIfSiYg2oPGwo+KdCf2
bWaez5AONilMW9ctiYnq7KL3JB9mjoaED521uyaAKKCD5OHP4YCEMp9zsmrneCM8
nLdOVx3YW586UP8Rf545od5tFJAFNWQFl0GpgOHttww6cqTT55CAjNqP7O6S3xeS
DOHW75EJAMILs/BHGMtOVIHracREWz7qVo8hhI/XrtSQHdNKxEo3kxl+l4D8hbFj
YqR0tSQMlb2lT9r2x3i/OURsX5auHfxK1ZbxDQLoLpAJ5BhBKmbccFyJyOxfFaU4
cV4B14gYfJH9tdIket2NMtLDCJfNRKGwwiyWVyrZYbf129pzT8pBB8s7gC71JHu9
Keq7cy9sb8CKKs/WDHegMp0MAVBFIHZxmtS7ECO4d0un9Px0dXpBFsgnmyKddyG/
7iKbKhicvNF/qHKhk3SzFgMk67EOfm3GRkLODIWR9+Kkyw6YgIk+LJLRhSrrRi6v
LoIHRjK361LG83owr73KEttHZgV1WX3vizG/DXQfFw3B4QVu0LcG9W5D+Ia4iTVn
YOs638SXffX2fDxqhaas7DdW6YoUnK1rdlXpsJ0naV/9NmN3WWhF92JhqDs0HaZU
b9Xlk4Ynv8cEZhXts0EWQHIOmXh0vKzlKvtYmgKmcamcrP6ryIIteHjrrkEutdEi
nHcXgExLGr0QbMelNT2xmZAq78D3fdTsZcX0dNfy/8exqWdpZkdDehiREVUnNxaV
Yg8imoIUYwrYkC5fV60nvpmKH+FIkV/8Q4ZStYeN8YhzItZArgbcCUsmcYjAxXCE
l3ilrN1dwzfQZwI8l/kVCkRSvC5lsbzMHcUTta6s50ynV44dcnvMCkfgRUsUzWKl
RpOeWHEnBp0piVGl0cG9AHMqOUVorevqBy0m/387YYy05Cvw1YsP3JhLANT46fXJ
E9XgUoTQws28Q8MjTqwZjySu2bsh6uVQm9sUQjN9lQCoYuDnMo+CyseFwbX6ZPI/
f8kMF2x0UmujDZd3+D0EYaVJkPhHGz3DWDBvU667ow7/20nIHkk2LNXPH+ec9RTg
79hhkXwLl38zVThpkHT1exZrSaoCXK5vWTv6Lz8scA+zK9eVP2VyCxjEMieV7Ju7
l6agBLM0Q6KMOfChlb2bjSWOGU/xHuKtOTa6T6WEFKQJyMdhc/Qm+vwiRnCr0caa
ziuM++aFd9lY/2SGm4HixezS6pv3Vta+rcbYU5l6+Rc2HxaFLaUyApd9t2roVQrP
6c9TrpUB9STHjxC/IKAF5BNMkXeyCxXDxSFMeqssR/WzhwbiD2gvooJdM58vvFWg
NG+TbXhadtXJO4rQ6ufoKtb4LC+LwLJJTCiAQ0ECidNCnCECceXkcNrVyag37ESf
PP1Exwzt/k+MxY0NpFdiWu7NDcWSuemOmV/DtrtLyUlyt/eyxf7BjeQ7z/NSNFPT
55pMJJG8ZowDTJfPrByQOwl9VJdeu6Xvl5OLfcqg//KR4h5gCx7bIkZXWcyaZRnb
+zS47SpMz6R5vcZcr6MhRBjO9aZY6zMr6NTdrXLnNtqEq7H6YtGzPmySZsxI8VBn
2eflwNmz/GeRtgZwFqrX0NjbcLEAU9lOKi5c10PW2XlyHlVyUp7nq1D/xbfWj4Q2
5q01VHbVRzo8KKIIu1vUZOoHmb8JaDdCHrcLgGUB3NlCKQxkIRhEyzxAVeNdPY4v
PpCInKUvqDvYRC+Ik7UMNDN8KPhiTvDebFZUWNCkFtICM2rRbpHGezQXXfF5oZxj
Tqw4SorFIdJ3AJlM9Bmqu//ezl2eF0lLJqa/VT29lrhaAfTqk/QgTURH7SdU4hIL
Ft/FR5K9X/3xEcr5rDxOvOYEO7fkIn+rsh5QxrRgDlPwOUL6RT/sY0yPImJ5yV1b
Od5dQMq03IplHLk52kXb3qzWI5/ismuzmMCKS9iug3jsIJymy5fwrn6VMmZVm2qp
vYldG3iSFlZQx5/aey6FGk+uop20wiCVBfpx4BpQV4sfybPFU0JGYadrThdF01w5
qaW4rdYcP7VKAqJsuhOZI+O0mCNvSFvl5pXMHj/Iw4Smw0aN7vP3kBCtdbJSDrW2
OiNK0ESJdWFkuxQyXojcJD8SHvWg6Ev8uHTEONm2TftmPn2Lj34yTv7+ptZbRNRa
H35JgUeEUBruqhhkJv/Ynf7Ibq1mLdBcwbPBWmnSEJw++md9MhUGQtCJNz80jPUs
0ASc1cs0YsY89/LB0JV8uFVEyN7LdtPh4z46dcJjqWhawJmGVpm3SiQo6G7zZ+ww
1ueUHICS337HTHn72lbuOynf8+RJwh3+NnczAK+36eB6O5NbTT7gEf8rOJ7tsSzA
NAs8Lvg9Cm+1/j25xm5GtObbn7KUeXb4w9ewomGmw972q2xCVT9N9eRrgD0MMW29
jicwiMpPEirD9crzkoBewmP96ZGAVuf7oJFxbkv9oBGA93vmU6hEiIlyl0jWKYj/
JQ+1CofEwT/7tLUF7htrfEUPgtbpYxzMaxNlRAQmTWR/hrPvEusCWP/oFV1tdXhY
yy/358ojOhwJtViWDMGdLfGMA1rwm1eGwEG1pSFQpwGmmrhM9nfHEErROD67NIvc
lYP+jUxzvbx2/gogmOq4J6Y7qc2XwAjm/d5H0pF+fCHyYrx8NYT1dseERCh8j6UE
K2KBeFrrnSlxP53EOP9GwsQZu+4xJ3RRZ9OimWXdNON1thdhRGYsO+Pk9m0cZw2P
51A4WJ73Bx+iTXaj/SJaLxIyMADMfnpnrwp9AMqs2EL9pPAy1MsN4sQs0vnKzDRs
hahLsVhtAjVU/05z6okiBMxKFRYUIT8jAxmAwiUbgaV76jRS6w2lIGNgvx9U7a+Q
/eSgD2uhcKBCSGAUHZCDvMJi9vdfnq718ThPO5vLTJnu1adtVJzckVA/V1Sg3eOB
E7QMKslFnMyXT9ieimD9w932XN9UnpTbq6DRJsQzFSfKqvRcCLT4KUXXeIydJ32+
R1cMY5THNPniJpnF8mLS8hYFM38av7cFpec8dUwGhkZCppgFZttwZRtyTxyssfQy
t/RMwt8AyXJaRIfke+juEeRZM8+lyBpTh/XtTiFOFm1CZyLkhlV5nvSWgXOR0dFW
U9So2mXiZQa6Rhtq7CWkFTMliOWlusnmkbyln3SQXsyWQnRNwo2wOYmJ1MoREL/E
v11NB/5/raTb41ufovZL8f+50CgRqNuN95AKbk5nbdpq7weIUZ6VSJBGnM2BalDQ
u+z+/cWtejHwlrl3jo6Xt+L5uab+r6ceaoK+zAbBM7OLMgG/Qf6DOodLGshbCOu7
RIDXNds7EakiLhqZlDqbB7BGdYxQj5betu0cIJb7Q+omLYtqpq45K98ATYcPvrQB
1l75/dmAaHYgmW20jlgdtiJxYUGFCFwflBBDAtYwyplsb/XS2Ntn3+jP1VFQNs0B
V/c9Cj/lkWNj7MGtPeCaR3Aw9lq2aFlkxaGGRaJu92eOSUiK9cZDo1a/SWE9luMF
LaY1GSyjPk+SpGlD84ePO14dbo2mWMkydmUqFQzzVERietEwu/BTqSYZJ3Hry78N
56XEDVzm4wK/OqkiVaMv/oJ3oWjpJ7YDor+9z/mKnn0qyKcUjwD/qOcCWQIUdueJ
DJ+MERGu78gVWqPvmWM5CAceEm9QyOmhhBiYB79dnIzWfFZdm3o+hfPmE9syoEWK
Cl6ngezaHP3xWG/hL/dPv7zgldsAnT3J2YGyCZHRSpfMcgYna7Zd9SHtGdSucymh
5d9cgUvVPdjXk0N5suVImHxwFSzs9ASgkS3KSkO9XTiFcHuOMKbJ69Dt/YlUv1uC
RqHfSwnWESY77bw+B+UDstcTyx7kdM1S+TA5Iivlwkco0341P0nPD0qctN6g08JZ
oCdzEqed0zQ++Jv+PA5vPKOglMy6K3JONpnggAy6Mnbcj9fitzRdLo/AhIOzWuhz
JCXYXKnOtObvK0NHcfQSz+5UZc+dXsj8DS7vwN1ZdGp3lADoSFnIgLmXJ/EUpBPd
iLMkRNnIIVkvYTE6UlID0QIgl6gPMiLTwWSL1aoAefOYQ4lQpXA63Nns9wzE3L2N
rF2Hy7uS1NU5nYFZ7/MnoNEf+5IFJdLBasTtGrVL2xlbyt5yW4xxiFsWlqES7JI0
GjSgZWhM03qoBGnustyGPc5pDdXrnmTYTohMTCiepvUOR7jljjhjJOprYgG6V5Cc
fzZsrlHfrCILhowucEYl6v3RRUwz0NAK13CZWxg6Q/ikhTzz1LEGL4bNqy9yKMbJ
oY+PE657Th80rkZvriM72xTATWsXGKdxJObaZe2Ex0C7YcHwWkANcsVH8zWPrk5H
YfyNNxiufQst2AIQ9SlY3rgaagAK/k3Q5Zw78XFThIj6Oa0Wg5ywnTaXZ26bWuOH
MIVt273Y4AHf/HVlFywdBvy9Qa8hbLZy3kQnYs80jbNNUm5jz7nch63ebCaMghdq
yzwlTt0ccWMQCbiNXcQfu4kn0S9i4+rQQSy68XBhZTya/Vl58sKZ9tN0F2llRX2L
sgwQL49miw8ZPjdI1Qx7B4WC1XDuyi+efE97ZCL/QU3Xq2oXxhBp0kAdhKB0LVQs
0zXCbBkLuigsKxTpiGFsY3bHX/JHynQdTiCDsJNcLmMeRcH83QZ52XZpM/x4pLv5
pFoANx1wsUoc/RFu3yvCXdnqgDJk56any8WGTP0eMs98viwGkdLhIHzApUESu3Ug
QHMNlL7tCtq8kYFmfbrlQLRsuS9rREJHhFrka79MvA+4O+2paTvbDBiVZAhsjZOS
SBWKujpkkpHWBVabmc4hvcdQY+3GKLLhGCjR2TgSEAczJWllvjyBq1B7ZdPPh/U2
nNVsGC6whiK6e1HBS7lIKvYkYqvNRfYV0jFsAGb8Zno4Zfw9vUusMxRmiZciY//Z
JbRMuUWll1jNYQRYMYtTEsP8omnnekkpUNddWj0Tco6Lpm4xqPiq6lli8hS3mIql
tMkNa72ng4cC6pJeZjEbarNqnyj27dTKkvQaqJ8kuRzgEcRJTC1UtYA0zyig3tL6
aEczgPGgql/prpHMGc+4kKRjXdFn26NkmPdCZmcIFOTDMY8QLzuMigNAbNrrAcyD
kvU9hsYAibGTj/mposRB6PcpxkX7puuYTQkf/KROhvf6XPY2vjiEVpX5QgbZAvsM
gimsOalhg3NjejgihNcCb+pJtcieU8zkQzNKhPkiVmFd4T5TMJLUInwWSW3rZp6y
iA81X6SbUM0CRwWgtgvl4O6mib6SbvBe3V/wEHo36aEUCpPi1cPC9MmTeJm26Jt1
rj7penN9r/Lb09bRrh6Vfpw93P0vl+w2lPZswVdsPlnU/u2kKKLMi7jw80FB8OC+
o81ADVnlrqC3lJsvnnUHpRYZ5WfrMLvdjrntnDRb5IGqqDhoSX0I+wSGFAspLDQw
oR9EqfZFZtMbjZo2rwNEOOn9a2adlAFzQnvoCFpHyKxEOnvs50c28mj4oBR56J6W
S6ZkV0AjFDnr63x7qGtZCgOYC3xex7L5LLsXHIefM/MRFRaO0BuJhN1gmmHGlh7D
CEm378uhscTgz0MBa8g0xahLXXjNSPcAwash7kIxMygUF8EcDUoSJMoSuxGd6Bl0
hhlS/ksbE/RjqsMEUNqlcDUdG14f4L7MsKaOMFiLiiX/XRvniPRl2Evi1h0FjENe
3GBHW6w5cnpzeKtXVxxIl5iGhd9wZM5gBUu0Ig4MX71NtlxPqRCax8bDLo4Wybvr
yxJ0mOQ3oc8mbAtKLWWQ7kGoF9f7XbZTZKfmZAC+V90rzFPo0N6JYZKbd+zXuDJS
BgXl4jFo31/v0OWnk1IsvfiSiUt35f3zhR5If3eprHGjg4M0MACTlXAC8H14lWb1
/m3KKdqEqhK6wPO35s1I8UQgi5N2GcOdYcbQgB4OgRHF2/Zof0s79Pb0xzmTj0lz
I/SWxLHdHFitAGYOsb3MjdZkFuvXJrduRZ12XHTgRRCGjBFTN2bTNqiXvQhPkCNB
T6qC42a0BKCh0LF/pF6HwWOwzPfaJ3bmNSlu/90/Z9OcIE7yoszCbBl6XkAc/fBO
49uNdr/e3lllBP3nkFUdKySqd9e98tWhhqDb8glabGSTghudVXxa7w2C0YBoYpue
DPvZBfc0rR9fJ0J7Bego1+HY9z7Fl4qB4lNNwmBuoTxMOUpRNZkDQcW1U717G3cq
1dBcbRqxvujd2aUDN2CdIT+HQ+57B6EpvrctKK6V/Zp7xNj1V/K6T97kxjlsyi9s
bD1pIfuuRzzzhpg+ZLsDsVny/XcbL6WLwAa5wlQ/+lHeLijnR7lclC40ZGZaOAUs
42OE5q8vQcrCp/HNTGY9zIFtwZVcL3gy1vEzKbxddPu8wFgpl2EdNYpVPuflitPH
dQI5fp5KJBV2xGwy/8yQuv9zLTSsXPjEgk4Yoi9VkXBFbcYrSbnzkiXn6pf9Ze4q
ybs5CBSs1Uh4OTOWZDVJ6/PGszwlfyntNi7yz35XwuyHXBTtqMfWgoJ2cp5b/R9m
MDiPLXY8AsdhCA7qH3vXUgw7RblxDkStt+zq67ki266fKlNAHyNLVdgerOCj5HPH
6C0kK3tpAhHDtUU2sAKvZ2iM3M/ldGbiobZniZOcFNBRk0iFy4Bho/YMzcuvgOIt
aDFQQeFxsD2/OVQ3KCguSwg9S9WwVnu8FnmT/QajnmFTN3IqJN8Gp5LlhjWaG/rV
j4sn4gK02ATyt3DMF5GWJkkBWme/MybIYZKlu/0uDFr7+2KDn7c5LFBbBB0hD1oj
AxvqROWUElnimVMC6OhyofOeajsZOYEUZoNlVcW3tFbUnhCVoZPiiboz4sY6Ead/
uVRftexR5gO4gmfvleNIqcbru2udwmLJN/NL6t0aTAyKnqSoyVFYfHkIyD/XKQgX
CcjE3zChq6Fn1PTl+0Cuklbcogf4cddaa/Zx5lDH20zKLnl2b6sJsYIz3I0++iuE
A1eA1lLVkM8RpnI0Qhazlsw7gvEEQgwB1qi3/ZiZdAaUgiiaRomOW2/3AO6JLHpj
Nqkd5O6CrPuq0PB0iDrfufnQPKKL9tw33fFXi9JCbXU8TT3cOMaDAISroqqcT5oo
ny67NE9sB0XqI4dCC9dTmjd5p05y23+4CW7jqkGiAh+SOrzItnR2Muwsi1S9Ujze
eqC4UQWgQVjNhwPjKEp0ZSronJNc9RVAc/uaKpJbUY1xDHBfaOY8aKuG9w2aWn+p
JRaWKGX2RtGUyKwQuFEA07sOLBstZdGUFpSzmnz/fEJ6Kg3+kdKS5SV+4Q7eqB71
48hPbGhzIERy7H1YS7M/nd7DSnxX46YHSb4/pRlsjPydqjUZrKxg1/TZgNf5ezpq
A81jA5z8g0LGp2Z6NvSvCeoDVakeGOR/4oC4sSIO36WvPcUKi0CVgXjmQLYfsBuH
dLpbLS5O4Teamg2+M4mUbVnXLE73t3G+UeNoucaM8SC1P810VBbKee9sSTOSPq0B
d+OTPF72v7WtsH45auM13HorDPhMbAkDCrfmLiJycXhl4oJ2eoSHE7YjwmYDBlAJ
/l1LY9rjIbqWmQ1NsTevIYwaT/SU1rGlkQZDGVqRAxSnPdALU8lbzGvfOjEMO7DH
ZLiPqsaVtBXQp/0qK1Kdui1dNsR9kNsg7Og8Eu7C6tyuLiRSl6w852andQHw2efP
Cpad93zS3Iwz/oaWKSAHy9Gqzw4bsi5nhFPmUJ20AeNBi3CNZTkUnpgNF7aifDHX
UlKFmjfnoNtftw/O6zv39aLJNHY9s4HSkgYhWwU6gPfWjZ7dO4RKKlNLq3ByGKlC
zxp7RF8GFdDupHkfAD83PJSpoJ5DrUOAaRKk8d/cJ75/kPEazwvYwNXpQeNL5ubt
/27cWQJetE2ihQb0eKl9yOQmOvrFJw1tIXJ9UEjeKhOQm4ow8J/VmtmeLSXjtGOH
sKKpNy5Oh/NOycS1y7GWBs7jUJWaUrI6N8ZqFIi4FVlXyHoCNLOSTVc0kN54oSJU
fFRXOp2JQ4dhiLSA394GDpe+Q7Vv+J9UzDpA4cknynT9xjB2Qwi2FnRq8I2JjZVX
BYKZ+mFA4v6Q7aDeShQsz548BWzNgQ6+kVaquCcfUC+nIDPXCaKlvCh5ThT3x2rR
iQFbqdEwPCJk12EjTF3cXRasolWIMMbv5gL5pb06Lmk1t87pV3OWaecLzV+/9lxS
EBywsLRGKuCzMn1PLqIM1KgL9I4rA5osw0gzhhbScHH6hIGmWvSBOxuM1Hp1SC2E
fKF+ZyrGf2XtkadIeRgGjyQG1QnpwQUpEN1sVk08JhzXaV0Tch25gjHFKMG3Cn7T
Gfs8dj4C851DpR0AFOwTsZv7t2ztgALLbXyG8y5aiwsJ9H4iD51/9g7wYjPMn2Lj
aIY6cAA6epSFQq1fwUVumyRU2OL1NUmTQx94adSGAhqp0QXZhQUPa7opX+XSTAsG
yeRzrYM2WK/NCy7G0WsdMo9HNK4l1++y+MxrHg8nVk+IAXahtC4eFWCTs2319Un5
VHSKqFRs9ifqSBAcY3pY50oLDIPrUxZFcg03ko3ZSIU61J13iLYAqHW+o7krV+ZP
z1cHE5eNJ7hSlIwOj6yiqq7X5RX1Lq6xD4liFL6bC/lHED3QEJVJGLPkxA1lInf0
LDvH+5xyNh8jPbJxJPQ7gWxZ1aSI35y2knxItPGyPC9Bzg1HWZP1mNWxs7Gvcj78
TL8Z6v0K8t8NMobTrS4EZQ22rQrSEacJwzUFkY8RjPEGGW31Mka36UxcXy1aCsNc
lcBAbMYfnZodAFklYD6rthOG9I9P++1C//xKCCO5OcByK0RA9H31Cnm9/PvPg5GB
yn5i4JNhAMOQ8gHfZOqZAOnHE6kGpuArlo3Pv8l7ny48a5hQBP2QHs24xAUoZHXi
Q33FdXStdWeU5dzAf78R+6t+tDOW+CyxWkasdBLWI2dpthHQwiIXlNl340BdxJov
KDa2LC7uAvbn6x7klbNWfXKdhivsRcZg34NeyQ3n4I94C9CwRtBuxl3mKs6qv+hM
12HnzR6H2H4eD7CQM+68NF4s+5m30fk/Jwg3EekUjcTL5ZEh8t4V7N3upegxMfPY
4FxFASC29Quq0crp2qHGBv/eVrtIpwuPsnXjda9USV6JCqg6HnpBxe3qH0zKqjyF
fQCYaZDGtYJvlk+NEnQKg+AqCLBVDEJ1D/WcVuPbHymbY0kKLgphrbOO7bMCTmwt
D3sLkhd3eDW8uJN52di7fIgOY7ynDzwBLVshcFEiTqCSMu7IU2B49bVsQ3Jm65/m
zR8D0g8sYNTKik/jQYvp2xEMABm9/dPkVvDFJscSgdOc+j+vr030WQWEtVU4DeoU
py4EcE55Us3tp43EDL6dMuS5ojb5P3/jRZAF6+X/BfMK6l24gUU5qiB1WexRbAVK
rZU40t5byl4wgo0Qy/F+0mxw4s7XjSbER2NBfhyGBTSjR0ZWuop+tJ1d1aKYrpXa
a2vmZeni43PNTPrFuU8h8FpnsQv3Co0ypZxh/MrE/slydkn9kt61NnVlhf/HCmX+
gZdeCYvLKN+SGVWEAbn3vjI+7xooodccHGxtjlPycI7wTmyNHc5aMG1C2diAwfds
kmwjsPudPThdBeMe5qq0642DakZxVCMCxfAlUM5bTGRB2rzldzLWksXCv1B4Q4Qu
NCMZCECVPlz9GekjqehDHTljKjwcN+tU07Kxvh7Tjigb8jvm+ktcMteMfZ6lvgyP
U1aLpjTxTeII5rb5ZR0wQtZu5AAqTYKIYB1e++uhaYm4nFp181k9zt75ziojb0Mm
e3WBnDAH2iqAxrz0Mk0LM9z9FmtPnRzcgxtz+FBX8j2QJCZTw6UgbZtOoUkdh93Z
SXA20Kpze9MTucTGQbzpgqbUqN8f8FUy9NvYLmVPhBjHladsCfsGO8RnPF5b+NRo
viHJ09KbC0AWqtnYpCF1JnM35ZKXQ41/UTh1/WedLa77b8brCJDNvyJsvbjzTNs2
31k2gJhlZXXlsuWLrXKCUPJ6fg1YetzVZZd/yfgNzaw4V/OfoOr2uCXmW87ZyQnV
BAGu2hUaCNaJkBBvSgXZvnYKQDx0+vZU9H0S4tXQXu1zGJKLSbit6NfZgoBNUo9h
FQh8hTEn9TYtjLjOE6KDz+ENig0qJ0VEvmU6gz4JYiZe4W4J5Ma5KiL72kPiVNC4
XwgDPO2GbKs+ePG8AD/AFhuB4N6ceHJL5L/tQISxsKeatlHhYEug112OTqZc1a4m
us+S5f4DzjGJTfDqLZR8U+wsTOo1RqIy377LXQ9LK+bD+wtDhLAA0D4yMyHCeGt9
Yk0NDCVFYEDzhy7ATzsHt/idc6BRSG6/Ux+Fq2bWJSSl5/jMumGAP3aZAfdTGLoL
lv+u/Cl6JMGfJTHC2rAHNmHLe2z2KEwMSUYGz6eA31PWsfsGn0HrB/cRNerhkdy+
uX3Q1MA5nYwqonzyLPHNn/ZktfyxC8OMhBbTYrPcE6d+IMZcepAv3eHnw9kMZN+9
90KHb4v99yywj6v751mSqhOp80hP7dJ0XqNblUBHZM7dFVYx6kgfG1uuW0rc3+9e
q51qHlKfgrp/gYySApZTmfPWPIR/MLE5afq6kf5rDxnYbFwsJS6P9lgDZyuxeLfA
M4eu42vp7hHUtMZG7Oiobphh7DosXfRE5uvhPn9NpD7U398J4iOrn98y5mMKsIQX
J5LLWpIeV7ITRsLJIgO2hg6vMwEzyCF+CiXB+bA30mR+FQJoB3iZdfoJeNuGzCUV
43aqGsB/YpH/H68GtigIyDSrk6f18YCLlYRpmbYGWr9u9BPZoHMrl9dPdabss8zE
qrSVlhuX98DPRp5TXqIGmVolyOF5rsetVFVHBs7ABBM12s7n01Xvs+xUQ0C0zLik
E992JWOcvYjDF5BNBCDSm46yEwlp5wESZzVkNsTZr/DQOk0vbeguY3FGcfrrkwA5
WPesSP91WtiUodAqwoW1k526d/QQR6KMIVZlpwbakxNClEcrtpYyi+/I0jOwckaJ
jVF7tqhoJL5dNJQolbx1fZUHjHTjHCxXLvDMCTqvi6hkI3so+Bi4wS9Fi0FQRcKS
gmrra9FoWXvY3YW9EfH2WV3h5YXCmLOivK1y1ny/KI5qE5OE6HO3fGgYxQiGB1Ba
N6wcFA4THdL6GEmjc/KDzn/Vk2nd1XQsu3tybwEVZytaJeBE2ACYkHc6bM0qh0BO
cRmLH2Ji+h4XFkVo4qdcvLcFAd6ekhs2f4yBkaEfDw5WzWjwF46JgPNT7vCCeMXA
RCogRqWMuDLGsw8CFFyn5FXuEsjeGbkxHvqxWF9qjMwO/3HVnUXczgFypkoyhWzL
Y5swsiMJNXXDhzcRHX5e8cgPyWkFzruXWOH3L1wYxz0Bcy/ZyOwwhZrKQwzxuzDg
pkWS7JKekCw9mCK0k0pcEXn8Gs9+ve9f+kThqCrYGoDDIdbwfMGk0vetmOuSu2xx
3B+YoEFMCr5Oj0+fb2x9iXHCsooD/gMb1Xxoq8IZQMqUIp4trlsN0hu23dJv2qtj
6SzagbR1dJGANEZwnPdUOyJ8uRUhM43/C5ZfUfsKZyXTSe5+Lpq3eX9VCm6QRLJI
k5UZNJicTX79WnHHBxjG8E0W594rQY6aOlqZmSrpzeUH5f6ItUfMf1xT3DAia5fb
65gaHLvqR7spAZg265rNohdwpj7jULNSju/wluhm5OYS2FUTTbqF7B6AX2+a0F+h
TpSwiGtlT/iIemFyrSRAi4xr6FMdT1HMa+fHMvYgyMmTFjCc7/f8zoCqNrJ+oS+P
FRnlRc8BCfSqo+nAxX1KSBjqu/HIb8WCLvpZCEZ2XMH0Dg5AYXDiQLUvXTOPXcOB
blfYYsTwiq11MhJ+fYHRuyVojXSi34igkL3JzJ3Z60q6rW1lpaasSYOxiWChgzxj
HuXdwHaHBb0mK84tBuhsVqxOPIWbZp30WYyVShrAyVUz1sSgS1TU3AU2g2zZhMNh
mr53z+lvl+w3q53Q3yA+c8Jns3wa01AOmmslVGzGP2JvMeJG/FFSE0mNw/O2dfDg
NEtOrhyfshEypvHlYebxvjviZwusUsSCF8UVEZXmTXNPoC9jbLFa6GCiJvFefGD0
bDJsSHkSo/cnuhn6q9kq8epDAtseid3PfkogkwyEELLeACctz0+GX5hBngYiUkNp
5pAdvDMoy4c+Kc/bYLCbxpdWAItEqyvAVlHznhW2IfT9V75IPJVWnKMbW6AbV3X6
EETVHtZhFmMP0Kftw7U5VWH8K/bJxda9TqVcEToc8ABfgp5AR2OIFs9WV/kirLmR
sIWB62XLhq0SfKTq404H/YM01IJD1UdrYGdmzPPuW4kaWq4i0Kk1hZyBCbtS3Yds
JJUF44fttJxK+EFPUuST6kNN9L0wUy3pUkYBcXI5i0Z+Ye9G9BV6GiPSMMaldkV7
7PiuS5QFo9XlTP5MI+i7AbpOy36K4eDNTfTRDgNgJbR7rp0hbDYNOb+7UPKr9qtx
9jNQVj0cqp9a82W5TqYqNo4iFS3XDfCwQUWqLR7bcBF2o5/O9t7HCDYRWO6B0dwb
M3qG46Qr2GcC1K8V5HVVt0ZDfAy8/Hces0FVc/XdxlctpE87/f8Lms2vIawMt/yu
w4zhqkRyPDo5q+hAaciHNICGuPg//D3BjEqtNQU4qVwehvUkdzZQ2b4c4bdCzNwI
8+Tkfn1WOjouoQRx0CrruNj5YaUrqY9gz9nDDifMENHBGr/h92C38qZpj8f2lgq4
tJH8Umv36JSyr8r/THuydRgorzo3QSGQ7HkNbTd5qqzMsmipHs0onjlQeGPV0jOJ
/6J8y2UZ793qSmq1iRbQ/XpZRydV7BD9l6ERHIIi62+UglqJRufefPSipe3nd0tX
QoLFhRnbUdyj562XOFYH1Eev1nznW1f44uoCKM49gMTs4IJpA6YMQe2Vnm1cizk6
VrR9ci0Ej0N29WfvyFGlfitTP+CgZr8F2E9m3tYZl7Pw99gx4F9US+w6r2ROI1Rh
u6yEkwQT2zoagpeJiY52tj8PdNO3ieESZHgxZw3rwVPgWbknWSQFR7Uu29DYH91F
cx5BybSf7A+2J7/xZTx6j6H8qQPnErCFWq2vu8DcAN3Bs7l6kX9RoVezErOD+Gw/
0htRClo2zwmhEmy4ezK8L6ukJjyCaqkvywHMidXfi0u3m5p37phtkE9EJAa2eNJo
DlS/QNyCD0JKg85GL5mMdfyfLRW48aRbeTnkTeshnJ1xbYK4VPPq1t22zJX2tWKc
QwnQdbNZ5lEoHdqSn8a2aK5a+hYqOT2AniwvU7cvYoOg3bjPJvEZF/RUo4FXlfCd
hGUQMNB/PpkDRzhzpJTgHLiwG1kdfVIFztOpN+LlCwuibOB52muBXLngRZ5LUkMN
PK3LFj5X8ZsFdNFYT1hX2aJ58qaNqcrCaPl6lITjDuEFfxyKF2NhE5o2u6fwMEnT
KyaGh2DkToRoNrvRvN31TVxsNuAgupFAQumVFf83oudGOcic5i7xekzITb3d56PF
VjG2u8VsnyEwjdE6EE5UDvhjJHYYZnOZwdLr75zJx+oZGCqFtU86bwBiISxGCQ2k
9I3JbWrLqSx3dhMRFNdU3RUjUAdKkoe0W4sIgnQLqlMvQCUMqDBCUx25KLcG4kLw
gTmPuDcqYVmVGpKC5xKb0BE2Mrx/ZmQNF/J2Y1vZ5cMOZhDV36BUohs2npNknjOo
2wGlw5SsBLAMTqylx4OfsgUbcyeySawgdygl/vLyq8Vm3pybamO862RWLZEyCOvU
C4B5Vpwv5tORlQpSTDiYsE7Apl5ZnkIPbbq2Ls1znQfUVNQ4XBCcsHWkNfExsM3w
W4uCDqpOMSLCa2P62i+K3D34GGYAjY4nxWAEhoxwcJvjz2u8UoGdMVsJYxeynFw+
uzqZFb2YsQ0YRvI6/uqFpYPaSqvW2EFRNnu7EqLtChEpbuNVa8imy0uVmsMwJSiK
4m86LGt6RHdPX1DiRhsbiQri0um2A5uHFyhU/EiLRqvQFVGqm1X76lF4s5IAtAz9
aJRArOdCHyJ77rIqhdku2bXJVHZSTRhmSV5nInmkCvPo0NBisfrvWWvN9EkmfJ5r
zQ0OzPPm7am2ZsTfn94DKR/knMwxTW3xYy9aGijrJqNorpuSuCoMjkIVjGr1Z3Ys
10yhNYCO0hHivtSnuX2r4U7t0PslVQorSBK1AucRknYllAxK/DRGIWkM4ZR6d2H0
C8xVArCyuOlc7XM3ynifwVXxPsNZ5qpJ1zv25Q8DWDFuZo2zULyG5EKvdvGWZ1qL
OTwkUf10z8IGDBQrI2hVKahGd79ptdyy8DwU1EYnC+gseWiy6sGdIpzsAiwOBlUZ
14JEdBiWT7X8MEa6QA3z8jhWXjNbBQS9BTNz7P71956wJ9Jo1qlR7/P2NXj9LCus
TP3AkJTDzkj6YnyV1TbI51JO+dF82EMY7/7NZ42P3NVmxNKJFpQRJIsRKUV3QdWK
PGbNILJ95EL+56IZKTOqPJqKAr5isKHb37dZqtOVPcCyDSpPdDZ57OIein23ubyc
qToYjdu+xxu37KfzzJd/wlkCUGI3qzmpprvrvKZ+4+qwNm9a93OTQ9AeXjN+t3oe
BDs0DZGxt1XQXp0V3uONXVii9O5RRBgxdLeX2OXHSkVrCiYA40NXso0j40etXnzp
Z2whfI49X0UfgzFto6VNVX6dWtR1CDjIHGfqk/d0nmCZpWAV6bU82vyHDhgMsb4A
fx3CQfNgzOjHkknSMVbUCOJTekWBrHzHFTwIyFn3gq7WAKwztjKZFibdfzjk7CXE
vMwZ9q/OyF+WBXohKowzm4Rz3O4RAwAG23jkPOxr428jn6TV85Hb/T7MB6YtKFib
ThWldOG3rWnmDTgRidULtP9SuRV4TTDcAtFrFRGJEVGhrdRFkgciVJuse1S0ZKvj
LlVPSt6+RXiTfK7d9cB5KXMpcGRMviwRr1P5R0UPksquJINSKpsoU8r+g2awye6Y
bk5GwfNCjU1WxLDXHvNLZDSp01E+E1zq36QlOxMcuWBtl/efNTk2vpKiZBRr5ENC
HVmpJoeXSov9txWD+jhri8ugzgmC/SSzz2j/tiM3pKUB+hX97g137H29MLiGYPDY
7Ndvm5VygGH3+E8ZzGWEX4V0HSFJ/Z/mwULDs9QAX2d8hKabzsxgtYzI32r0p8jJ
6O0wCTZfe8lS1+pZvUwXJ89ekie57b3kwRjN9M2SJkKvRZGGvwyBze6EsgKEx8MU
Q80k8p9/GCsYW0Xzbm7ahce2XaFNJmGU7/dwz6cy1rXiVyWWoETTARgeY/L+OQLp
woqbQDGipQHCWunJ01lFwNe/NKkP2/3xjlCzNFFkIMs+trRT4YH0w7mVEv4PR5nk
mLs9UGyUijubWcVbx87STFsCDf8do6oJdEL7Io1QQHFLvHlNXM1TFf6Ik8SGSDj3
Zeh+nwVrB1bqELS3rXQE7iTtKW9B/ZsKpsXSsm1SP1mfzsTB7xensa9pC5PmqPQd
jkV0cBaPtfTBBNAWI221TfFTJfU5IwgtPobtWDcoQInQ1mAyft0LG1n1y+TBSPbR
XK8m+x2XojYAJbRu6vq+H8l/AvMlvnxqDBtCJkUMm8oP7+GdetsB1cimOfPKS8I6
xhje8hrmqC+OZTlIatMDZCW/HLgzYEftLQiJTC5ImQyshx2xt0ObllABdTv4tSoa
xbmX8lAxtivSM6fxc8jtOSUr0RYFO4RGncYipCzEHVA2DwJeJv9zZqC/ORHrdI4/
G1/JDdTtTKIV3Sco2BFVJZFQ0crPUWaW/z0w0TqzxPkcFtGY8PF8vwLVgmlkP49e
CVqmMTrzw+Pyj/d7AziE1YCMRzTtv5u2QhcXNKFLOvQej1h1SsWVfu2Lbv7YuJsi
rw1XoSZbUFaqUfJAcC2Z70y4w33jAGprzs7MfFl/2u3ht7L1YVa9BBQMvsHP0PQA
2nkA6K+bjPRGiw1GZFsyFaXTCC4JZHq6twboEfg+IkPhOfTJqGiXo2Ow008lmMCG
RIwBu0EpzI6A4Nt3/pj93x3nRezClYfe5/Z2sfi8kW+qeViDmlSu9Bf6skPt2zGE
c0gBfopKozozURu/D7IlWnLv7qtGTKXJoBDOd19QoWpFMZbTa1qpOtYbqtPpNESL
drXihwaWNllpWVmfeE6HGS8Sp+ZalIi5pLBfF57oDMPFnkAuFqE/Kn4wgBMTLSLR
DvTxT7EYaLWtj6gCelEBxxggF/jIfdGb2N5xmKx+2utlBPuyPsv6p1tgGTd4RPez
ftD2tl9sUUyid6XWVUM8O1SAbugfwP5DIyF8c3SCKpd6rLzU8VyjJbDPN2pIo00w
bjg5168oSjY1AP1zKNrKyW/kSoX6y/FxvUr5QEg5f3GZndYYixe1fhpnmzMFv9lM
mMiM2TtML1ZUHBSP668U3gisyHgpQRYHhKXkk2eRtqFHBra2hsUZWvfPuF1zq56y
VQyWAmyXmes52OUAHW0SP+WkzucJxWwdfo1KOULbfZ1K6fEnRcMyjDS4BRGNCacr
uDuFXwUBBIGgW48zaaVk3GzVD7yZYurO1XaWhBq4dzjEBQ1u4ByvwGOmKCnoQyE3
AY0al3wucvBoGJeFdxGhGO16S7Mnjsa4mEhju+ErgVyt303J9+DLOxl7tvCa65Pe
rgimvqf2/pN6krG+Ll7wp2a7YKPpKhyY0VsaV/itDNPLh7ySNuCxNtSYlea/Tji7
MbVCnShcTwdNOabDsB4cuewMsyVMDN6GQrT3Z85HxqaDKV618volQYDo8MvVdtr4
UpXCWI9k9KUj782Veu3eu1Me48058x84uYZlq1LIFRuVXT71jwOcITv30vFxpDoW
AjoUDaCgbrMAURgn0lAsmLQwpYOCbPZn7uF0CWmmEbZsd55CCMaPZHvZ0CxthZo4
pHJZPPTENlf8yAKHmfWAjjVUVLdnq69XLkDo7mKeXwB+yIwClSIRh6uJNJ3o9jZa
JDWhnvOJxYXCbESR1ujEJSCw9yNk9ZdnqtQbOriLO1n9YTmAcGg1SwyGZHHcpzPB
Weimt37RjTxBwO83noCuMwRlYoaSQ+MAZKkgdIwhsfypW98PrFUvkWgV7kMTbJV7
oT7MG4Jt2hhtPagKiUiKlR0ZPDM5hB4msN4C/GlMdn/ZcMXiL8aiRAMNsdhfAcen
fmywnZIUwl91fsHBNKjLw+ZntHvWz7pM3eb+6yNptnsXaxEBCWCR7PneWQ6vdNPI
ER8HkPsewwrv6x/5SMYjCOfuQAV/4U38cFbknyT48PRZ4+KnJMNSwyWdR+m6gD7g
ofk0EjZrdPqp+91SeBzmWG3cYYZPpepk00a9hkNDdMHmOYiOWpbouNGJ3Z88lDHy
9IaaY9UTMAKyEwtJcgHywLXOeNRmMg39C3MZZ4pYzM4OuKWOwy5Y9KIrfZ9Obb+3
g/jpfHW9iSEg2nt19AXJVONTqd6HE9q4kFbg2OazrFmta4Qil4G/AfniCT4KW88j
GGHd23+EakVe9GmFATPtYOrJpAk4drX7K39wBflwDErhAEato5VbI066GWmL+eS1
bRmAGmTu0t1wQfZIbhte1AYSy4uPNT5ekJowqKOHr+yTj4chjd+H92nSuEqdqK1z
U3OcnziXVH6BlGoWkR6IjhePO3wgQ2NrrNVZxUVwnqxEU4rCPZ8mmDjc6GnW3YKQ
7LTIxyzLvaAoEMW+DYycFql78sOTw3tIEfUc1n0Gvn1onA8iFUjicOq2b5+dbfqa
8ZY1M85L6Jc0uocbKYNGG55m4OgLg1sIY8Y7mfNcfHWmG83baebxmbx7F1rMD2O+
AKbfhuIAg3xAcOeWsoPgAaIAaeSq8m4Onas++TrpKrv+8mQsIbXdUQSpyqzViNMN
W3DcwDMfU/g5Av4RG1+2sGg0dW0KYvyy+RgNhFQvnjZepk9km4c8fQ3jMzvGODKk
qYI8Hz5Jnnl9E+0905kLmqLnXyRv+AEYAvyCQVOjmHcamodRIA84urLW/xBE55ui
d0STN/LFIwzZmiKhwVASlb1BKPKX7weEGPeACJPTZfIzXY4QTaczufVGvGLkunyi
nPfxWAtiikZnjR9b/KrkrfoMKKZsvMz+9D6+C0nP9qTOFCKzFqN4Y9gdaaY9toS7
VemXwQGcXG3WDVKjz6NIGH6SsP74M3tn8vNPzJ/aoPhPlJhwUl87pxazwTlpjZYP
z4wcBzXkVYGs4AgwQnOnY0nlGLH0nznka4s3T4XjJpLxxzlVDeFfDrfTQRnkZo89
o5zUSM8gALoSlq7I9jSE1EOdZQ58eO7fOoN5XP5LbTTd4FzR6TcncoUQNg1n/bEj
lWXbfK1ykZDupC22hDTP7ktGVo4+LHs9DkSx3MCbOWgMU9R8lUWbglMrO0DPfJ+h
fCm/EQIgPXj1uULul2bv0yARwo3BR3LY/SUzIb/s2aPlYYrlJLK3P0SdNm4tTtLV
s/x8Zx7eKrFvX0FTvasllipCSd7BCNe0YRrtbPrKPu1I1b8bYJUGAWn4UNZ8+oKg
A+PDt1upJ8vPzYv1jdn+I+52rHMICrQb7MzENTb5/v9RWisFTTuvJ9lw747hE0zX
VV8OsNbelEtf9JUq4H9sGzsAixuZMyjqMW0ZX+Imh/bo61uApqoRE+hy4twiXCST
rUCZfI0WOsL0oEzOTqHh9/+Su0AyQYwklyR++NYj+t1Ptd5yEZMGxO1hwdXVxCAn
LBGIhOhDDIUPCHZgu6My2eK5jy7LZryREVkH+dU8xuWO8quZrVcdXXRocJv5lKrL
5UQZMwSs112OQz7mlmsg/qdxa/V8cma5QTKqH3SeqiZxpUj8EOI7rjPbFyz/E0Gm
29ib6KbSypykZCoUdcCKwlVUIhn8oP/2GpmMsDqPKXNRCNaIkR6FPKwnp1pzKJsa
hCi8QHMqC1BNEk9Nwp8UdV+SHSG3YisLDvLQcTnFtGcMHWsELe80HEYD2hWEDUcP
h0HOyWTKECvbyfk0rg1v3OqHoanEeR2LpsZz71zFmUFAK6wy0OqHxyyHs5JAg2Lx
TynhnVn2Wo2xY++gaCZwAw9hrS74uEFuRmzt7F13e8eNkY4VgBZhchSc94QndtcZ
VxSjLlR1f9EuHVW2p5tS6Tk717GdBV5FURldaMAsovuXgW9AqKHo8L7EhmkLK+mN
QtjpUJDDTHtujJpbmB+WLny18FqLS9UWuzrX8sSgpqvZiGMQ3zp5UuvOSz8SCxAM
goqD3gFg82U/yr2RFAaXUZam6Z9N9es6iTcemYhzhxeSCcK4o6VyV/LyqQvKaTul
Vf2/PvkPn/6eoI33jaH2nDWR7DsCDqFwyMcH/kgWJbYDU6aQNs1e7/XI4lAYNCep
Bp87KnXg9fCMIEkEeV0n/L/ca6/riIHy9Xhbawp1Vd1+UpPsJYrs/F0ln/565+pR
TJbkd9O33S9T9UkFmgV0Xic0W/ECEAkNqBRJVfJJMq5Z0kBUDE9tOsOxuSo7NQmZ
HE6kYhZZ1wC8XhH0I3sfFHb/pIWze/zybD7hzaMt1z+7JltDaUkSZC012161T60B
DJAqcqhyK8B+KMUVVJrQdrtiVssFFq25Kqf9DGsKd7ZM3Bqx9wCguYEmcQWLn9yq
89jFhBZ/DcTiJ4Qf8TMsK+jYLOSx+UV5SoJROVfgwKBkg1zn/UdI9Id8bhKto0lL
X1LrnOPwiX56wqZ6B/ON8BTGiNdV2g4v2Lt2kxwm9gdb/urV13jRgXV4wCUvieEL
QoLYPmLNrwNVYrG1KCwTqZZoMsarBIoEyskGJ0FxC05TWER6+reVRL3a4f4DVQ3+
r7XcyluUbfhyQXfJL26Sec5XfFCD9jumJqNvd/c6oaB7Y25f2VcidaVsYbK0mxwc
jBIwNwWMcFESYQ7gUKr4kY/SJhcqpc/dwlp7jCTuVP0F92B9QOWVPmjebxwTyhGt
BfOWvGnoKjALNSvHSajlnjVVNNl3B25bJOkC3x49M4z5Nkqq9wgSrUubV2gWBH5t
xHuvwfuyH8fqOE6iOdfT8vNpCB6iz3k/UAz35nStE0GOT+Xcv8Mkzqg/j6MMiH5Q
SNTTxqWNZu/B9jZcq1BbbEsc6aqYjzxdcvwDnd8FcYFWXFr4D/qDLssUf6l7Vd0b
Pja9c88xY4tqNni5905Zso4vtaT2Rbkzm14A+N3NYX2C6jEHEaY2cqUCDMo+LQHk
/kPh2BSWGr2+NGDovzk7iOfo7wx06XKbIx7r4C4OlnQ5SJncZ0sEybk/olFqGVC2
mnVRMcttHRYmd9iBbFBhqrgV3eTxsJAGUFhSMOKcwsEkCQv47EaUNe3LzgzS6L5i
O89hRbymJPdGnEZXHyTu1fVVRW/yhO5sjaZW1jzsi7IyJsDZYpS3NsERiwnDjEOA
iQYfFFrLzUcXAEy3BO3zsH7q6gJaO+UA/uTT6mFKbsxBZ3VqgZMGWuPUQ0cLMOzf
1Zw6BnN4AF2smhTfTPUM9Bfp9LeoSa7qUYoV4VUO8MYJVIeVnZNmUtE/vYMMuHBN
LeS2se3/BZL9wPvuVy9xT7e0G2SfkQdV+tIXR2sN7mIwAuPaCzMO5RN91MSwk0kT
/pC8n0GgG0zB2cxbdC0s4cCWQnVU9PFZJJmHoZnq5nNxDwwrLGP8i3YZs9s8fXQy
ffOyEMVl2BKkBH4LiBYyPZW31MRg0CalNjP0J9kRlioQ50OMbeO4cdIDaUj5XgYW
+qA8GNvbnPVl/U1PArqsKrm/R7SXMKmMRFDEKrvKNO0kLgCEyKpSBVUHFb6n2lxJ
irhheGFsknHsc/4zjUBenWeJN1Sb4s3U+uE2osKEcAlX8FN5vOrGMwKsmVTxwxoM
2A/ItYZp/hSYcLHax0bXz+NMxxaNazzcnBs54UpQD9hLpRN7INlXo+VSa/zk1nWv
Ri90+N+e73eS59G9k4RRfRcOelyBnPaC/MhU/Ctl8p1PC4c/EEBcRtrfbQYty4tt
U+BTXDzW7kx6HReiTg3r8yVR8lsyANthPsIMG4ngNfcjXBSilDZg3jqa7w41uetp
Xw0AoKimtal/hY+qd0XGQ++w5Ws794Y2l1iJO8mpXqylAJLMRN3wDuTiPvGlYmEg
v7SC9+LZ0SeQevbEVT2snu5k1IeTSoXFcNlRPUwzqp2d2CO5L88nsqQPzziM1O9n
pq4N85W5WedPXvP0SjLYUbvCXcH20P7ymg1jn6DzQ/BQiNObpTupzwzncQJfePVx
pHrTvaJ34vJELPfMi1xaCWtsdUI5WcL5q7p9QJcKYQWcJUzk0jUOZRaLtulXP45U
mCSt1l9mhYpzFsim+3Z4utztf/A8Zaccy9bZaazWE3v+iVFUJSNkdh59CSdK7JmJ
aquRbOGb101FznwbdiiwZMeifZkbu1dOv7A/13dT7czC6QgsBHozlUPr+5lNclTw
XwLuw6kyLNmLG1mEZG3yAAjbn++cpsCeVOKWwvMr7oZqL1nwuYhIN9LCfGop01mp
KBFvWKs9K/nNsmVt1Gz0ItdVxoQ+5Z/hlWdtw84xg2f/RShGNmmTIzlhL5l0OFj0
GNMN3KMZQsnHm7DPl9Tl7oMdkKZqFh9nzphyrk9PvjaqXKOS1uNXhlxH65nd0DSo
58f1I73se7vfzytjCu5E1Rq6Xgq755OgolbiF47sPXlVombh32ZtnrXzfBBS8eGd
3CsbVb9aOgE/xmxJ0PK/9jF4Qbx5Kv53PBMUqJCsr9v51Daz9OgiaY9q2Nb5WBRB
4GprsYmZwDlkBg/ie91uI6VkJgCQWm1gCpnqNIeJSb0v7Ido7Vohbv2m3R2U08kv
zUw91RDB8m7ccAC25XFXrMulpEUkdTqdegOYNtGjykcPExasVWy6RtncWLonMRlq
aUWRYe0tquabAUWltwXputKA614L41PPuUJVN0aRDgmRBmcA5gZklicGaQdL2TM0
MET72LSjdQYYbJKGn1yQYO8mvkU0EtoyW445Sj4AULJ0bcFWZ/OjvIJgDpZhuSPr
Ba9dN3L1Ex6K8tDC+K0ORCI0j8tjjoS1/XVxzmEyd71VhCiQKEpsT2ZloiFBvsI0
8kChZ+abHG8IWdKgx2RlxrXHdTTmpZyYabwY2ItJB6QVM41lRyqzOfW3Pdhgn3Hf
0pMX/fHUSZAxjNENyDYvJSwiP9ws6GvE8Aoins7/x/trIxPUdnZTpeuz/Jy+QDop
SSjYwQHN2yVSHwWFWRcxPcINZQHa/nNYFdhurxm3v+9wy9fAyLNQkDDSDXbyeaEb
Dvy6pn4RQozFJe74HmdJes5PQD27uhxtrVnPcg43Bf5nZ0nLGwfH77kzbIBHsPTA
13N6miUq2QaGLjJRkOqRTrs3rwqnXTsd76h5fMZFKmLwJAYYsi5f7mEN0r9RwlAf
eZP8lG9VzYAEb+95GcHw3YjN8SrgmUeMTgWIRcpA2SteDeDCVK0cKAxT0Rf+P5NP
r7IxMlm4iepDzJ8zBq2d1K2yDcQ7HmohQ5V1qjIEvKyT86dVvvh+x3UUNq4ji07z
Iu4r4756dyUQWhwT6czd3jsWGqC0BCWAAFrF/TYPZ59SCvrLFE/Ci3un3saLZiVS
OxLWS5DOAF3WI7DgbPlE3wTGOn2IwCPP9kBJh7Usgqe3CHhua5eHYPsZtw8RzCVg
+dlH/a1WRZngKchb5B/HxpqrQqASb1r8NDbJqXJNwtCy7x41vVGTCPVcaTbfxtrq
4Sr6CZRbfkxJ+Fo3Sqi6lclBvNmQvIArls03sdlLIYXK2arlueK3fHERCzkn2U2b
3MeDkYc1wCNM6kKhVh/bZF+7L9/v/oaFHl4hdENQgomjEiUJrrBK630aII6Bq1bf
OAO6xaWLLNsglKXe+Ow6JOx3Q9C3Emn0TeBm/GcQi3ibZjYiK4uWsKSQVBAWsT0q
wtwisuQWmYVdPM5j6RZGFYsVJNdB1Xrlqbq9dsCc/KJHoLku8oBlDDI3ggTVhUGm
x3UhDKqjayCpZf5qq59I3oVMIISpJprAOz/CVjDbo2o7PlNEX7DxIcCKwE4UUU17
F3DtbQaNR2EjqvIhWHK4AF+dNWg69y+wz04wdMR3j8yrZSvLci9vZ7tc8++hkUvy
9nU7OK44VrrC2GqdKK9bdylJ4q2SLyNGfdFPkaBT5WQ/4iukm00jCOFOsE45efqy
jrNKvp51Wfpk20FktS/DhE2c65a9BG/qZKkAXeBdlKEeD5v7Wj6zesDZhXC0oWEB
qSs0DpXwCGw3QVzHvamMv7zM+MkcgZKHw/CKB1MYT1jyeg5KUWXgpcgc8uvRgkeU
M9suHjzS2340OgooxreOgo934/shDK0S+5TxXmD6I0S3hSalqacMF2nIpCFUzq3h
DvfoeX+HnLp2kVM++6Lfn77kHQYb1oihR2RWnprklT8i6oY6KC3Js14/kxL18Ma2
d418gLHsC/ViZW7KN/TGMqH+DyKzaf336uDdxQXb9ej3b843L3qQy2tlpjPBEdjZ
hJdIpd9SyOWq91cNZmzKtdlIDLkhsqUolTYQWuta4JTfuXDlV9PZyGxg4X2LSaVu
ahrxx9tMJbPRHctQ/nIWebrBZvms4BUn1edkZlHi6a5pq7XZ2PYWluUyKKpBHRRl
4WUGWefClwKhWDIYdYPlCXX+5bHVF2MbeXJGn4eYlnNHN9/RB/I6/0zAGvXAHC+u
wGjUvBJ7oRx55izL2mbOz3/FSdSUxcfVlsh2jKYsBbIrTRInERpkxapK76ETKHWa
mPD/TUQQ5DVXB7vMtmi2o32p01Fk+Rde3QXbcKTHtF6TxhBALg842dbf6JiXZTgH
aaSD2Laoyfwkvtr908WrdIcx0Oxw8kmw+dT8Xgik2SRPIIxbqUljdqCtQrdcNTPo
4Olkl+neFm9f9kCC3Fyp6TbS/QK1bCcCEtu2zxD694EDFIlJZVjZcLw0pELSp0Pc
M5Mg+DviwbDzEJFYx1fdQNMW22b6U/4kXkVOuoliQZmJYjACGZ/KXt9SRgPKW868
LvGKHhQek908Y29I8/tPFjoB7AqCOhhQI3M/rXwJV5u8lY70fX++jX5BzQU96nZu
0IH3nJZ+JBFa9wlFGTq333Gd3/9ZMq7kPJxsW/1zcFJ/41dj9o2C9MSgajKWcTbt
MGREerpGu1EhNZhPDlTKeTcJSXeHYH5PPhxxayDWkv1pOhToRVLCiI3QN8pIvFP3
EAz0zc2/Ji8gcsXTflwghVurdrGZQK6SnoE9EtP8DUxnvOX8bTA2n8L4D9e5iUaC
ewOYzS6VN5oDnpcrnpAtS+QaeOojPvMVZfImHYo43ChgmkCFbDoTqpl0zxAgfk2g
EjZNwHco9o6tYJrcGxKnHCS1wocqruaCpSNxK5WOZ3OgMekZo+dn23iKkYGTTK73
6fLcRX7zfx5PCL3ScSJkYNTQsCg9hbhawBtgoVG6PzlHWV4Yq/tid8Wjb01nxhBA
cIBzV32N9QXV1sloYOu1swXg0LjB/sBhmWj1aLFy4uRULwr46KAOep5MgAY6mzQ4
2bUWcugKdofv4HO8ZRG6pxkyzY0AAUQIld6x3CDyRniuZXwMH7ltsLaT5x+ai/27
EK1uSeYz57of4O9o/weFHxxZxfTH91jPZNz0JH0v22E1aQvJwVu6ANf7T8o67lg1
Ucw+KYRSXxLEhjHRFnNN34sDgCn3GKfNlGwixB85fSiocbQ8AM9ySeDxUvmv9w3/
Gtif2Zc34xl1TTq+WCKS6h0dfc7LR6y5BW1lJtgq0YII9h0tShSo5DyIhXNI1tOM
o2Q4UD5S4t5LHkOavCjMX97NkqEccLUS8uMOqhrPRnXdPEYTXmkj1A4VHZYpc0JW
8hKZOnSdKKxDbnRItmq1THoCWUWzvO4i6T0Vxe5tXIEjZQb3wBndgTX3lDy7Bg2C
W9DfeYvLCOmTR6VrPr3i48aKYuPbIb6f+e97AjbqWYvlnudGOyZsTBCheg50cCzC
u29GWtieIy8ztTny0A4+LUf7V9c7G9NWshBFR5HkSqklf77WhAfc7gE3QZetLjbN
ocdRH5MABeXhmOYCpOsm89nQFQPc3RwyavbfskHNPesZmbXnrh4/MpFGe6KcKzvt
5KxZKgqiNMMZeVL1ggmwJOh3Otdho/nlCX+NNfVEhFUpwARilbzwFVouKJjg3rCi
L3Lxt+2K0D5dWhvsUWmgI+lcFWWA1PSose9T1UQ1isasTLxGZnAmh2nZbJM32Xjf
pTv3TBw8d07N0CAfpIgVIL/rjEToxrD5ZuB5g4Nmw0hmXdikBIGKJS6zEMRZYc9y
VDa0R5q4VJrY1C7SvJrdpA0l1j9YIA3UBXkf7klSSNaCPEsZ08byn1zK/eYdKESe
7ChnW6bDE58ojvAovU2f6h7bsQCwd2tfLyJ8IxBqQjCwfMA0WukLGpasXbeDmI4k
WXQPUhkL6yBosZxx7R0+aIKbnoM6qchC1Yq6Eb+Iiu/UOma3YjWn20WIIIA3DChc
Sp+RkKVFPaRoh9DCYKhP8rd5G2jz/r0KP2trWAUsLitkwixGWhlTclDIc2IX3Ycs
XfsigHALVLhddgz6/UzcYyw/+WY81f28zlm544Y5OZoFsjuJJtI96azkab4hOUmp
W8V+QQydAatnepFp4CHco3TRZSfLaHohhAVl6MFuVnpcofSG0D1Ab3cPBpxx9+RX
tHbuo+G+uEvoT1L/kL57qLYamLow0wpS0Hnt62XNuX/QEMVpAqzCo+HVV//lSvcN
Y3+Gmg+uvy6ANp9wAwIHbk4hGwZzkwsW//G+O+/xWwnDOA50opJBSYI8SfijKbJW
7b9VXiv8so1rN3bzo+ap0Hfu73btHSTAsVRnv/UhyueTvazl0UolPgcQpDpkri0q
hCSlYmd8c7/y9vOiVATZrbXVUgiRCzlP0hENQPoY5pd51aBNM1lsFjbdh4vDATe4
gOfeHL5i2n2wLlVxSJtKH6ux/BbOwHHpeO7thidrDfUIxJv8qaeJGapXQyKHh8zW
5FD6gGtHq2z5SbQiBN2LoAVbsV7/h8wrxxMPlZ2LflAOyn9ukxbFuLvPDaY8qvS0
Wu2DkKEtnxQld18d+cPWUCzyk1frE56CdsBKus4KFvKDaeX9ULasoYna9uKkzQz3
HG68pzsxtTAkQf6nzYBBdWoZCCB/YJ5e8idy6Cb+gklwfl+hUcElJsOMzG6ZUieH
WU9KzxSGuYdIwpOm8BTPr1i988wwiWV8I3On6A2wT5XAl7eAjNSLCQoODayWA656
vJNWZYRsYxu3sSmtRC20LbiNQLvMaYY1cBqKDYRODoB26scAh3tBEQwdyy0awSwm
jUmO25jQZvdQ8N+s2y7wnpzJjzfB/AbMCDUwlwN4Zv2ctoEll8XYdgQ3D2FH25sr
A6FJI4g5PYw9ogNxkM6dGiC++xRiAUIndSCVZXMj9l6myZ+C23vg5mi4sYb9EAe0
oEtYm6EXBPMRyO89frifVdLU/X52R0tPGp/boxKkgUM8ZAvXjSZLm8QGVR4xf6kf
qYoSsxaqFX47QjMtElxqG4pp63z9pTaXj9oNUkQav94ViO6UAY5+LRHqWXMTg2SN
mR57eaV6efzBjr6L0i1tvU8ExO+WZgzvSM15M0MTGMg7/MYYEKUaMPMUwYSKHEWL
Hhb6itEXffJrkOyUEfgRXUnJobuZjeRrSiy9vfT/CUSgz5hDwm8DCYOe3DONHGpR
VYNameC567LzUrN+JYaKL2zcr2UBUbFj8iJVe8fPxbT0h2H8jVZbWGeOTuIBMPPj
pBfD3bCqnpUpCm+SJejXlSLv5S0WENuvmwBp/xugZWZIalSoc8xIghOZ0iF2pVqn
a4ulhzKL9I1b/4rAAMDmPLEnPAJUvVKuuAXPd3jpinbCH7zN5q6L4f12GCy9axkI
97YFYn0A/xkiSMlf3aciHEbb3/pLfov1S5fV+rRIdrppXOtTaR8ll7SXa1gCimA7
yUWkjZzmZF6wA9/pIgSpLxys+IKTFqyK39xVyUMyacw0bie5rnCgZWHiMceOKGF9
AYKiLsQQLIIKVJ2yCgyQqdRIVkfzJBWbkadG5CtSsM0NQQRu0tC7Ya7vI2frAqKK
sM6/oil3pDoyIkyVMrjmYzzgzwQ0cgO5QI64ykZ8fpHe42B6iy/S5wYhT7IcQVC/
kItIVmiMhdiTPprKylp8SrPi+Xu5tI5iN8Hp/I7hpLYWtPKgk1QQj0CDQ9zpEcQ3
VCkm6c54iwCrmjVptEktriEY5TwzUHAUKKKkZLAheDMoZcuLxhowcAqUsWHvAM5S
rDYo4xltBwdcsPIgF7jdm56rdLMsmyQds+RA0MjHMzRF5EdksUrbAwDux+qtX8Lk
UhTGBApct9Liz31tfuYxoyCvR6DQxyVbdV1JLzqcFJiUrgl2Dn5iintXzfwtz7Hb
5AKC51tZBRSgbhPYhbDPJHLAvTKbYf3FJpdCKP+JAkvO9niUTFWDRJrvyord7mCb
FqziVBrNJuughyffDH6RyGhGrodwfFIiutksrixGxKtaAJoRXQD00Fbev/866QfK
ebjA8FSEXQH6QHeiheZwK2PUx5054OJ0Ey+3Ii4pxZO0NYTLHghPXvqajVsnkxu2
vATq/bkWE3qkP0LosmUU8C5qQKqcFnLDbdtTCIkJsgJ6Yt45KHW4T9ZRdHnY8NtJ
XAVcXAxbzh9z80bhMtVDobkRGmBCj7AQv70796eY274rz0CJoRU+x3E5YRvIx4/Y
7OmdHvAjkl1AOPtg+QL0y4jrU8BenH2GC679/xdgrrzJB66GXJi4HG/GRZqknCte
7o6cBcIAovULDXzJCE1ZIKWEW3ac3jFBaJNlNFDd4ZzSv0M92v4GfjN7gpzkEHj8
Qx/h5AALU5cIDY7nzbtNkcfLGgyyClfkjL/WVeEQU5sNxxhyb270fFvRMJFjhOPl
kIqw0TU0AJHCHWcBD+LmOgfsRjqsQ99L4IDpCwStUXn4JLZGbPiHmxCscDgI1Bj+
fkhwzfry4l71PQyVR9oNdZDYrRmucwNXRZvDxmc1xuNKp6Qc7UbRhxveLL23nihq
Vse1nRdV9tqtXN8N8vK87u7KUCxBuCdGxxq9XDYvaR9KeUjHxQnVKZY4yWIGdkng
g1zoSZhm5li+3kmsp7i1TTWhGdEWbvwd0JaPe9mbuDBcr42SgF8NKUs9O7t7zSnC
lVtb4xmMdgY8C3rLTNbOErvc9z4I22lgw5Zn7vUNWJN8GvsfK1b9i8CgxgF+9JUp
hgkWutFX6P3XokbbsKzGXobryYtwzF9o9UsHbXPRIwGWTPlQFa8uYvmjxlqQQ+d9
aPZpl4EWe6TwOW09lEEJSFW6hu9J5+6od3HHzRw5773XAkuZkwvfDWN65RT1t91h
mVbA18TlEX86Co7iWheRqbQcie+eEUcK0VzR7Uk7LBCaZMAORqHluzUlYVZLTJjo
3yr+HqvAuHatXSwcUMp/kGYE6JudDgaoftkSqzE/QBKP2hyspNxW8Pv+MN5dAmZl
zqnGxkWDLXjeup97OZqyUhVHbya/VwnttjLJO7oQhnDRDEm2T764G7jFzUZXpuTj
jI2PtJ20/VxdnzfnxtqnH64LFlKctcU+7aNOHCvzFle9JpRScYl9POqaYE73ie/v
MuJWOsOjlp1KIsux3X5taLGX9Kq0faWtvXTdKSEEGgWxF1LtFsl6YQEm7wSLX91d
z/Zpcsuok2qkgGCfDut5oOLy8RX5akp6UkibZsMayaWwvgtRDNqdlsz8MSxW4Chu
UFst+AX46d1+RZtJlSCa+zBQ9w7hKIq1mSl9DvbLzB5L6G+flxzGCKB64iEQUMNG
RM8FxRYhG3UfexL2R210WJYDCEUxTrdQW9CBD4ZoBZczNv5JJuovky4290uV3Avx
RgJMuE+n1dspiF4fUy7+aVT1FHlwbU3l8S9yfRW2LX6p74TEH4UtXR/qBlOQLcxl
yyMbA90ypKh5D6LSi9ZFYLuGUHBskDu/vlV75H8KUJG8wOy0/n4d+rhtNmzM8+A3
z4nOI5qGgrdlE3o9ju4MDKdlsSOc4KqUE+sSLzAetw1eVkJARyBtOnwva6AfHjf2
43ADcLEIezE8ivgrEA76W5BzFkdGtK34gWuRTT+Vx/BjeZl49Iyq7jD8jjOnouYN
tN8NBKtTSJl1iDGZsMfsUoTnpkgHxN+jXEnfaqpXZZWgb/cGZwhbFt53nGo3QmRm
SFJ72A2UnbELo/xp0pCtDIvk6ZzbULGe96cs0jO2GdWkrnYoKuR1ItmRPcfdzPAX
tLA+DBAgZBli142RmyxRriRUlvYks18thcaM6Ul0Vu8MjMvHvnHJBYLvTfzFPDta
vEcFPYNWyJGpvuyRV/cGEV6wKddjIBGH/vdZhfoneJxEmkVKcMrFxJtzjfpewmXv
FSE+fnNHm/eZOK57XOJR06N6FnmkrImfxEdONnx/WXhA4FonGbpH1WmzbOyzfJNe
jBk5RLnaSSxxX7XkCeLbS+uf7Jex+z0AVDu90N4wM0EhdCq+4QSHi1hSObxV61P7
0+rgdmrDgCVWNRlJ7Qf0TQ9TDRs59Ie5QucZBwQf0AFESEW/Y7FcNEzV/cYUSAkv
RyPu3yaRSA4/y7Iel+lWLrb+/Ze8X/Or0N+rimH/Ml2kBachcvmmb1DShpJDG9I/
S0Y/hz+Fyy6J2jJUmQF7iAbro+0QMWaeP6OEMTGQXs8LK/iblmGzeCr0PZ7pbMzl
yS7qVU9AkJMfiP8xdd6VY2pOnOCq2eeLs40sVE1orMHjnj4jZ3LvbtVelNuEakK0
sXf0F4n//lVaAubdIhygnVz0iSTGBMQaY251KqGfmJ5BvLFgKtCvCOccDOKnmymB
WOgG+diHIetqXUZsT0x/hy49z/CR+PBnwBFDwvjO9OYJ7FVnNIPDnN6BsYoi/3GO
P4BlJzfbZ3EBlUUxOXhsneC7P1qBlzuNff2Voy9jK1kpemoux0gr9fDAvaRxxjg6
926Hhn02syUvv6UO64Lvxw0ahvHOAiJVddkuqf0YRZdyAqvxGqIjo0erKBhAeAi5
RwhU3mU4peQ8yEw+Tq4yIP5hCxh+sBjyHELAe8gqdjlPpWPtcR8i7/tXFUoA0sjs
o77DEMc6fhiz6nZFENsWcvXJQhar+c4jzdTqcLrjhGY3XAQm3SdhZSbQ+iSOr7aK
dIj09OXCSww78f3q2FAb7FXwlFftj4cmuafvdxTwkJ2pJRUG9J67+SwSfNpIIEyh
SfN9gBIzZTc2wnN9wFHyKnFACbVkLUDZGyRYmnNhn3w5Dj8QysPMzRtuOywwE1nx
E/l5bobOjLg/059Wxr99OwKgq1/v6XacUqXRjBwLyBgyVSABXRDZaDrI+49OcJFl
F4ygLisaMK+DAhRMD6p8yDtCxls5WFHnkZTiSMnUZv7fkEmO26eW8NibI82uClCz
yxVn2/MHOw3sqiJjTc6f4vVr/uNwy9AsCYFz/NGZzZn+4Y3bQL4nk82A4b+BV6h6
uj7HlDEzGaAOl7ZaSMmDTjIBHchJTi0RJe1+UkJ82o9p1NU8ApiXFpVvLT24CWlm
n/72xT9jxohrMBPBL33iwsQNCA75AmUVVxDqtt9xZW97A7RMoY3PMrimgDHgJuys
SZozKSVj/bmsM6+VdtfRypdExcCo9xDTmexN9FjdW5BdO7YCq+fYsLMZFc9nwQts
L0y1JT+xHIaAI84L4xVRmE38zGzGsajHC4/HA3zS7sO1XqrYAgkbNfwg5CW+n08V
/IiT5QKY+2GprMyJDt76vD0m0gxBl+YlOgdxHbI7vQNm+YGqac+VYH6zkfpc4A+D
CVLNftuEOVjMdFbfQbxWEzCvJdX3vZWBUVOOOckjv2hkgZCOUjmcN6B9vh8CDUSJ
I1X7u86yrPTNNZTXkbT4nJ/sRQJilGHR/lwcoLJMXeF7YRAG2FFV2LMz0yDgXm0I
alW+8RarHOiFa+fJRL8qb6nlf3ejaZQEGF6MhNjWZfSHTzE/352OxybkrdoEvUUW
jO/gIoDC+lS3azTK0UciaJclMv/ppXa6SkS5Stn9Zhf18DfcRDgqpFoenIUrbIww
z2kgekLXhHb5tSUMzmg5PpHMcQqDyEZz+QG9pxYmXAPBSlzYx3KoAH/jN7AEbF6E
Qmos04F/SIriMQPKfDICslw2iLRUFnqoCGLjYS0KL0FYxqTYPJxHdd4bxcgXetfP
a1PkRJeJIsdnBTgPV43nCOeWsq2PX9nqlSiFZ7DX2t/VSxh5mriqR/0cjoxuTLI3
K595Co0vGLDn9IfVrWvIe6qsbjSd4WmXeC9k/RA0DsSnE1b5jjIwcKxQ9nAVKAmX
tIaS51YHXq/QWLHRq8g/iuYV1Ymr7yGdA3nJ6nWXDRHMB2/wNE/s/TktOZSRbYoy
k/wgT3K8S2XNAMBUqZdy6oEN9YZEQcuQK2VFTmRuKQQYvwVUywreDOjMLH9IonWK
pDX6mqwewSMEWpeMTmkDROGDyWU+VV+U5j+Y0bz499BaBx1uLJT6a0SdbQLew6z/
mwS+WSO764FomwsDca9pvXFCGqVxTrd4kNH+8OcMQtIhrQC+kopuERbYNdhbMScV
049vO6g1bsLabkO68zpUFdjGsoM03keJkuxJDqK4wEzbvWGw5ru4PdJRLQj9IEN5
C86HoRyIliDgUlsKlmPaTNSCigwKbQIq2QbpJfYo2W+XEmqETrsouZnSpLQhk5Af
uO9JKCbjQ6rxEESk8qDAV1+K1XiVtjgNoPBZy2WCb3REEjL19fYrEXX1+i+nAgUj
NJFmeOFocNE7alq8h8Y5WDr0expkwUCIl+rgp4WVSs1ha5Vr1mfrgfsvYESH807k
3TFjpEiyXwZEx5SC0DuHAGnBYKUR+wEdnAHkzSre4uefp0ghzXsdoThuLViO0dBm
FqMrNlmUlFp4FcC6ujWkqpEEv+NRwwc/elzkxJoyJGAd3RJc5PSO23u9J32U0uiH
zj8qptA+JG/HUeBpnjHBSkz9jdXzIOm6pBFCVdnegejfmZ5W8iwNabQFRSqz6d4c
YE96nBEnuHpvx48vhrnu0tASb/RFbU09Uhd5I9gMgIs5Fa2pf0hSqC4quWg3A/Mk
JlFYyprwJQlAX1GysKEPsH9ToEbvi9/+aE2GLrWBCccuWYeBq8re7SzI/8BXXuV2
h7QWa+bjAQBmXOhmD2goxUydKvzo1+xQQOnBuyd3QLxABmqvBk+BL4mzVZtB95su
e4TC5Yrr+uWdOAG18/PRrJRnel2W8U/Inpnx6ELVIltANl7j4SwhSXFq/GvsJHKe
sJMqTTSixnX7rw2QhTSkMiC9M7OkPRHoovqmHEr+aD95FHnIvBYxI6Auz9PyBK1B
5F8PfPbeyzn3WEMKBXATDxdZN2+j23gdjMBrlYo2h7x1UqZOXzRlrGtlGW9csyF2
i/jfVmgr76R91LEXCbwQX0ISxu0NEEUEVcTJ8z4Rruk3Z5qYwynamRATLTEyQdUd
x49mhngU9lpjEGOAr576cvKRs/Bg7wi0MBgIB6YG59FRf7IrGiB5jKzNvHEcZuQU
yCCgqov+WPsQTWiEC4V6jZnoMhX1btSbzyPKccoQ5GL5z2rQORGza+it3O5MCslU
JR1JRInqwO5AgUnQ/rfxk+C2ND9+Jj+SYr/8snKI9p3Do4JBcN0GFZXqUH+qcEtJ
YKZcdYuu38L6zB7qn+T0vVRuP7SvItNsMk9OG78wBOKVsAXEha2JTbKLyXTwy7sv
vyTgB+PrOUN+i9WXRYWoOyJm3/mx0Htl9w+/wCMLiAr0rHz5dJ0AIGC/iKz+bRXk
LaR2jpOdij7IWomhdf9RTjIqxRfdHFUpYjIBrLD4M1D2BzySlTkZl3Eic2bQvPDT
c9Ce62pPf/x+TYnaWM36xf5QVPKAcD0MB2+4vTKUA7TDkQoWtFABoI7LX9cl8nor
X81Z5vHX5C0sdThigQhylybaMbHyV+hVI0X0gRaV0vn4GujbxN9KYC8LQpvw+MBH
Kw/YT22Y8w9JezQbMglaeVBCoCtcesMPfXWi5ouYmKGgmkAT/fCasjZtL7FaceCn
DDTbWP5hFgHNzf3LZYyF2yA348J5j7KUl9fOWUUj6PXQodTyEN5N/YpweIBQzikO
rnEHGKQwlyg2kHSCv/8xOSADJlivpL6DA71b3G/6CEbUI8Uqp1SwmY4YK8K3kh/k
eTqgf3kj5h2zsGvVy5PXF3IwHM3YOlSnsYyDl+Jl55pI+pNdI3j0tFSGcWX7x2O9
KDt4Xv51sReL9AOM725QPz8PI8YlmsfK/8FJ5xTfwSl9Pu6YmPE/B2KpBikp4hBX
cnz11xmI+XhdTa6gNBlgKuLBY+hshTbhBn/B1cfRlx9mdj60kFcHRaknIcqxg/SQ
YDRMYNuOrCJEONVHQaK8L5reYexsX0cRzu8k23ot5LHmTTce8bFJIlZlrasdyAp4
YQQA4MT4WAMyyo4RKcoepkASxMpHIM9Ss4gkdLU2O9HqE7oTyRHipUs9NLmGLUYF
GnyjeblHzYIXvIwQYr8r2ZaUpqAZR/8NdeOpso8VKjBoKeKDPFAbfmdIHbuJGJe+
fyWtoQAeBRlkB0gEnFdDaffKWUgrclXVH4H92A/htTXNFnMVn1SDDRggsVSHIcgd
GyXjKv57wp/315cqm1q2BKxuI3Sgz28fwnlHlEpdzgNv+KxBzAgd7Z668ze6DHyN
hpXpVJ5r+mOWF2/fMoSr9J+xT0en0c/rftJtGntDpdIoUnmasFUj3/FWPTkvegT9
PbQwhVZQfza48QY/52Dn1izoElA2lHrmCNMWsnLMupWdunHszrrL3apwCG8PN7kB
QzON4HAxXT5CSD0/xfPm6CTztNZNg218W7Jhiyp+LEp/HxJK/tQWlh2D3/+F0ghC
RCedgbm6A6iYR/Axh9bi1dEEDC0cDNb7ymI8YJXYhOPzvCIGje5iBuUUglA2TzaZ
9Smc7WOfB4aI4JsvJG+wr+uLkbQeVtHgjGTDqn5XRRRukZtunBPI41a2MmZHOlKw
xjh9dK/LWhv3T4FXNm5hc54GKGRIDnTeHnXxJsAfj+vopNRLzcWxnSRg2utosZ10
t5flT5X6zDLSvnnMHTRH0kLeEwddw9jqMEozPIuf62Nw0SuFGxL7LQdgCPJJQ8YV
MGtczDoAdDPAQxMF572aGQ7KFYAWe1/4AknmwvgWtX42YgnfP9OCMddZWbUqmtkG
vKadpwRNsw2VeUcYE6hZ41iWJj5MJxeb7hlPU67DuN14PRLqS2vmiEm8PqOQktt2
j7Jxs78cH/G1B2WJ7xRZMD7mszYz14uG3OckNSzvJo+skEhImb9WvhJKp6MKU540
A7CgeFnibdARwHXP19nC24qoy1oMYtCquPDMI8cc4K/3qFEo+2opneqiiWDdUI0b
82ks/xrMs0sn+uoI9y4K99NHkx710LYuRusWiHZUGkd08/4Kg+Tg9y2D9mhE/15M
j5zP0Y+Mvo/FM18xaVHtTaZ6a2mnu/2WKk3VuLZHKsww0/yc9i6+I87eUqa9xlP5
56/cRWjYakrzbMkq2g3PnZm3eJZnozE1uouAlV02PS+HDA2LJrqhLborkMDxUkZ8
qiJ/zLAGG6z6dn319i/PiQTOkD1tawrBoaulUOnOGY/hIfhqW119XkKgDUWgOL5g
FVy/anQlHhoUHNFwbv4bm97Q34gBElL1JfBySNLn9G+rkop6HHRYUZawoh8zie/3
k5MqAvtwCPLIuWpjQjq9MEuDMObtbpl57/5oeYDDC1l7sHfQATaoYivxbPxtqYob
l3hcdPXPLrc5J+xP8mjsEwfsJWy575W0oNwyCb9XER9iUBR2gWbT3AvZGfrUhfPC
WELNPPaApKIceynTUnrXrPUB7Od667Nc2DCCJ8DDMmV7OzKDN2VMtIFlRgcY6RUF
G7rzLdTLzj5pf5xSXFK8kDzU1+vsyz0frMS4EPtihWF9T5f9p4mN6XL6lFDdVFOV
T0TR55dHel/J1N8Kq0x+MfQkGA8+0t9X+7PvdKh5bph3KdT28tlifdhipC0PaEE+
d60Q23fU6TKKTgn3IzGfRM94JraDbdbPW8YWzsEcgtEDcg/SEunFmfMnE63A2LMP
uL0lFcUDS8qvH2p+jB4O8D+GTprPbM611QPpPPU87K4hPRWKRBLTTaZOeL7JDzqo
TBZhSYc5WuyYztlR7Kt8VlURAXpF44nAyVj0t9dIc4oU3bUeD290Xw8xRgiP4Z0H
SEBXWhMJFYFvhanP8zO9oQRVROfciLphk0bcVaVGoh9yP3f1SG0ZiI7a+QMb2SgX
SS33bn/ERGLhY/hmGiskAETD8/IkPRjB4t6DXSZy084qVsLd2Xo2pVC+UspjAWya
eMPSLIq4eYNobtNgkABF59Vgcmo8ItIjAwWEuuYt/YmqXm5m/dsku0MWBBFjtRRW
Qm6TuOt6iu+sTMD1a+D5rG483En+hpUyzSWdIm+ccggge2G2+16czNEmpFJD8MMq
ryGcIg/f/H/NjpoMV9YTSvBHKhJ2wuqXztXrH88QpfyeAgZDil//B4JdwsXQwH0Z
PjS/A6axBo/StPojF6eqxOdMH6xUBTsXJ0aDW8i0DTvFzQ4/bErxubX4eOpYP0Aa
KZpZSEFW6cMrBqUjWkcl+LiyHFkmNayY3bbY8SBEra57BuLUMTZuJ0av1heDillU
5gKIKGrRI0RNKCqVa2g6/hlni8ocPCJMjLdypoO5UqOAgG/jR+1efjW3GbnUSEmf
LaNhavzM9xL6n3DKjRRZ4DyCRXcMCg5Unn0gIGO76An532TcFBSkW8DmwxSSZind
Jv4c1Va4WHA+2SXAyHIev3atkCxDnkTOLM9xOArTsOOxIckhLNDOdmZO+eqyFGqS
5w9VcixB9ETtGJv+eVGqdVqOss5TnxU8IznxDfFxa7+6YdEeRwauy5w4E+mZq4Jy
ead1MMz5EtY01r92ENd3yS+Ml2DtEdQG47XbpQ+DDIC0hEbl/K8qjoQUAn5zVa5Q
U5a1KkuWhJcE9TJOtmvGhoVLRXl5bra6cP0SUm8QC24ZrIKTLEZ9izXlrv4BE9/T
K4QPMzPtQ5Fi70eCcyAZ7DHmEkxO0EIRbvxuM6dnHmy1VmY8qOG+tDKnBpRdgbjx
v0w6tNOwja70vICmJS1KSVGMDzEtPkkhLxfxEKG3RZl01FA3mqXvboyH/4yiRqMd
qu2uYrI9z1D2KkZxq8sh1GrEw3hceRAVfSHV1s22Y0exdrZMC07x2kKoBaNKqCzN
s+bdwTuFe7kdf3g2C8aehy6RPrrq7I/v1M7eS+FW9inO2md7Fl47ZyBUy5lko2Qx
WH02NzTBBwW24MPx+CeN6+rey0jQ6P5473I5iT1XC7Oeg+grTcooCaNDSprQw+RA
FOAehkfDAvlS/xb7a1RLl90Mj5TvBxQFfgznbRzko/zPftsHpiZKunjrT/oCThSa
G9aLS9/jYMZo1BWzIxmCVwm54cS/OM8cuttNmWHaL0YTW/8ivAuypGls6AX5Ukyc
716Ys5YYu6tOarMO2uB8JLe3VQGT+tAtPbjnzt72G56aARa/HUEShh9saoRB72yL
BK7gC5MhbXLo6heeBlMauAE4NoSa/4jFB9hHjWJ8pRUFiqIMQ72JhJwwFLQRJQZT
9loJr1kXzTNjAz+BOUPnv9/Q1I93hny9+92QYmy9ywoWfPPNeDYVqdxhJudr3/Ac
8zvKwOm/i73STyaYoHx9iwtTuG9wde4xRcsRTkLarJmTygdKT5G+ucK3Apxoe+lR
wYtU1yLF37p74DNdBHGhZey3zKU281CPZDHv/NYCIuJuJhx+xQYAhUwI3DRXvruT
4LFXEATDNLIAg0Cqe5AF+EYRwvlbo1eLAtAnrUGh2CKTmdIQ0epWBqHtrgKGqupR
m4Yld60STzvDQ8ORirqdrpuEherE2Jrar9HWlsVw8Becz7G2tfZ9g4hMpsqgJS66
hVaCvHGQBRBRNsO+VMOlQN7tivNJg9ak5cj1N5HhGRlyIvTa829dC2mNV+iUwdyB
Q32mtlYoR9by+cgY5mDBhEEkTaKRX0W8oENFlEm5qJTGq4e0EMIJ3jm6bvhSMOJJ
TYGQKB4VBZKN08iMuU+scOMBgdmfOe0AayPw7sDafwG6b9r4u3Hs+tRTJHq/WtYj
22rudOtIZkXw/AprjsGIh8wNajIRfbWOcvQiOWxm0VdQocC/XbGKIE95s7T3SgyG
G/+pQ5Rb39kzLkGBpGI7/K/cktJGR1dqbeneozbZ7VwDca9GYdqBRRcaLxBr0G4T
N/jYKSCQUG6iFEr9NE17bh3eFtNQQpqCNp9XQxPfqsWtAEkWd2jGnQFkYhQU1rwK
oAi2YcZHA0vy9vyGGOdEUhH1I3rVoAQahCAbWitx97+ZWie94MWEr5iXG0Ne281M
nYXcCTATNiZBvYbEOIKsOOT+JBHoU6yU1+rcQzJuePz4zVF15ul3rLXtSwlzd1Vw
H1sx1SvoowBvGEovISTzu0q1YawG+XjgpCwYrlUAH+iAkA3KF2a+DJGVr6leSbii
I/OOmHi0w9yic6p9K4d5hT8YOp2r2H1G5HanJdw7hqVngkY/PnzAWS4WaA19393H
TxjQXbyy3fTS7ahvABtMIbU50HWrZN+iZa0EylpR7nEA9e4t6xTeRIptukrRnE8Q
03TTzfmO6jeWjP606/pw/K+SFPW5RjSxJ3WjYARSjJ9u3u37L6yURFU7inYH0x4l
IbJ1gDdkXL2vCtjfKMXrKM07xmtU6vrvrkntmyG9cwGpgKCtmYuz+ipnQf4D/bn0
KBNV74ugFehBWWKpE5QJJKqTibesRDr1/ki3DfLUNL0/yjltCxv4cQyZqdU/VmpA
EPNI4F3w/jxwzSLrESLc5XZGPCLnQ4bNy315x0tmECi6/9J/EnUaB2vYos1D9Vza
UCOkj3ieTG8WkSghb0KfqMX8DfjND+uk5MZNPKgrEMG2iLI0TY45ByfsGNC2LjUi
CUG/PeInCf7dCzh6cduD7eJ23eaovGXa0Hcr2VjFfU5lw6arDcwaeQT1yX+nO8xO
EFUf6fdy1nCGhMTFgEaEYklxBAUs0QwYka/xtogf1XYJvK9A2o3Kr/UZasADfdVq
v6iM4ywkL6jVdccVS9e1Nb4oBBwm7YADqmK17RGkRUEt26eOhHB5OWx2M/KRRW3y
DkmCuTsdm+nhuxeGYmXEB5eJK6A2VwZMZ6kxtYINcVOeRUe7KgbPIDLnrmnVxkDd
HcTp1AmdJ+E/9vT5CK8o6kmnsctdqyyYARCHCcHVW8UFSudzvQyA0spDKsZZjG2Y
ERoQDUKESV3Y+++kPUh4LUX8co2psUbxkjuMKdjpgC6SKsiZwOvsVlwlYOMXByZg
iVX6i9yLpOuxW8rRVtUNS30j12mREEWyTy7tBHJ5R50K9n6Y4zWl3AYBvgMDmAJv
2twM+/TBOqZIHNJ2hHwv4lpaA7kdNuqTSBEVr7u3dOyiptPSRVJOBmaYMiSjFMyD
1t/D9nu71UEEvkQkLrbGWI5gE4UKMVMQdojMbbGVr9CA1xVwdjixuCZ1cNoqc/1I
DRmgxbD1jRcbJkHSKUQ2HStYQlgd2uWiU//DMErSQuneJTjMN9O6+JUdf9/w8jYj
DS+QnF72QNs4oSmiMgNpyPrV1hd8HcryYNJUB++JTZJ31XzN3FqzcrRb3jqJ+wqT
ZtU1a2XDrbDCYuYgiwyuOMD34Y4guZAwJ3fRIwQ5xG6YyEYnTTv+aepBax20Vftm
6Wx2UbRX1MY+k4N4Ymy9iKlqG2q5pPH6ZN2uM9Lnb4EyY+fMJq/50A4FKIxyt5fm
+pHeXuI13aZ4qvPpXATFjmF8SG6+wBkEdjhiHnMSfRwaIuZV9SSoo+XyvJb4DMKn
JIQRslwNWK4GTp2KriZK3hZqRaJA+WN6BWp4fnF+NUWPrgwUDfTuDookfV5PjLg4
thHsRHYitHFVn/aiSeAMRnxiuBRYZQFk8JUej7sqxZWuGR+SKNP/3KEWyFSV2Hfj
gTh3W625m52eTPmHqtvAGTucuUlcDOF/IX3IasiiGHmbMI5rYTrwRZLkF0Lw8LEj
DdLuciaHS3JJfG7ORZ7BDXf308AvbrRxcm31gsVnPaJhMGp253sq0vdeskeSl2Rb
xl3/Vmfp2jj0cKBXTqqk0emqRBzloXOlUQtKZHz+al9recF+o6TcH+10mirThhrD
MsX9cSoIajP9+T0cCab+tG5ODGkuPQ5mFnNQoQaLnYnanURsf1ozVlbh09INm3mR
8PqRpRE5e6lipuFC705ljo2+QcJxxU8MYPVhvx2e8Tg2XQQ+5PzhNGNDkeJtJvj9
yTa0iIup+6cS02OpxUqdz4Mkf6RjO/nswI3SJ99D2ZNpyaJmUltoR6wK0J6GKT5/
gTUVRuyTSVe92fHhAKZ8AUm2Yi00/IChIHWC1kzLJHxL1VJ+m5iqTmvuMgrYBLe0
/gyM2AiRWkVhbtXhUYmlKfyTM/ZWWli5qwFlsPu1gkU2tA3Dqu+1Zdk25v2gXoeJ
HHxHLQbj5LhFn25N4CfDbidA040TEXXXn0OLE0oKrc1bw2ERkhdTrxvu/ztKQSIL
5MvQtrDXkZF0yHSMC1X/LOV9wDtybB0jGj7vRQiAPLSfOpmZgbcFMMxNPSaj6+y2
TffTcs8WeIy9Rzris8DwpilrKXx5Hp4qcTP24eUwHyo6/824xyFJRN4ONHTdjqky
GtA2svQKuK+hCXlp1J1lp6kw6sbKZYnPFLqLuWz+h55rAahf4QCanyzc6B8LHgd9
CIBAAdh+kgquok0U7TMPtc0++L5JCu1/PByn2BP3iTXP/a7nvBeKuYpitQwB02Cb
YWP3fsOv9WqLtRZDW0L4VzbfA8dBvN8Ig9pCG7ejvG7A6lPPVjNF9RGVHX0ajl7/
7tunvhhPbRWyZeowmlLkMYeYkKxt0ajN8+4Z5Hy27hjpTch24rtvwFvBcX4LuqBn
bQQx6N0wZ8ut8pqkDfk40h6yJAlTYQlo3y7N+7iqAZZao2Cr6NQ48Qw91DgHFb4q
xqOP72e2uIwoebYWbDGRTwxKZGHtcmLxbVL2qT7BBE6B5zWpSX/qHbZZNUe7JUzc
A2OG9Qu64nTk3EEWNA/FopkKYkdjy2cDVy4ReXO5ucvEghctK14eqO4f1+yYfOqe
9V6ZNJUyVxlkwx4upKNztKL1E1de3q4di6Q1HFxlUs1m10hnDLbxOpo5nqzRGSGx
m41cLpS+tJdIMyVyn6T6dQCmefzpLxQd6nfG7u8qfWV+FHB0B2TYRIKIO15GgkLY
036Pg5oTwmcgRnpFDywVMVCHbLM6JMFFhB5Om9IbugJxwbi2lK8jDIf3dhl9tZ0z
eW1fo9bK4L/J3jWR1xYZi2+z33XFow+p0zBW5zh2z6dzRKal0TqClBRgEQWnA6/G
Ou39lqvwVa8JsXRpjoyZwZDpDPHjdOEoHJmP17QNXW1kzyS2gBXeYHvb/96P6BPt
XIwfCNpVfbw3XVJdjVkW3XzuatEzS40myMxGIObR1erjQKKQZ8kuZS2Ej0DCsLXb
BbRwoWNxlwOYI1ZN0dmuiWgBSrCD6+wFmO5U1tf7BOdgtEMtFMq1D3cZJ8mHkX3H
fPzixzHPIbpqY0+MjbOBeD8gu7YLpNCnLnFI7+5R7DMm8f3bC7QdorD8diULOzcK
60tl6T1JiPfMI2v49hsk6amXFUxEW6oKgx2WhPYyMRDnKYe5tsMAV41D/cTt8Idf
gOJbWJxfL1Ov+7AMjgDzwFIm9zAyyYiuX+f815WW74sPdV+xbj2FrN7bolkV0nZ/
ubBEsM6dnzueySWQL5bkdaBv2XCUChh8RG8z2La0TxVXqa7BiuWevBR1p04GPamD
wqjicLd0aTvciFnTDHj3nGHwCU8XOuGG44q/TUyv8+7NcaLRgABbHkdCJjIgV0Ko
44aCnAm5DRJouZug1SyeuhK5vd9wKKKKAHFwAc/9j5aHNuwZyaamg7+yU7oC7FSv
HEhPO8RSfsKi/e2fd2pzGQbjrx3dGRqJIMLQu69NGZg+p7aBhG8BVmWr7UiN7clp
DytPtzv7ntAD2QelzOzc85YTA5kNDjsqUDVSjrEcfJf5Mt6DdFpAzRNHJKb1u6jP
See6kRIfYUGKV/pY205XF4CBYgRpz6Ao6H5ayCmRxAlkVI7OkhfLyePEdkgjm10X
6+BGpGOgPwPJfyNLrpjSa6vOmTn/AtnCBLcgHB1HAgeTCIdxLAy7vlC1Ol/RqI1m
fouurSNZ5p+tP/Vdohpd2wQzrAatNSyrtY8Fiu1I7DMgyeBfX8TJCuQUS8hNMLH1
k+ctTZNd+eJTak05egojvPpERivmmFB/9rYVzbP1rMd3vthO+bdPnx0f8mgk8Oul
mrSbo4rCGjV3IcdVoCGo/HXYizORm6IFTaXzGyY3xKI6lyUiXKHuzJ+EONNo6OLa
XyNCgGbij6c0miCC1hiAsB4GUHZ3UJqLzpOv+RaqWUrn4ex2F8uAU/uQGpXsjlCK
xK9jlr1gqB//UYM8mFQqbNkp+ayot4Du7YNkj+q1IJr0+tONLdNtruw3lY8VQs3I
36J4ziqXiu8/dwFwpkJgRymult1LlFEW9T3Vt67fa2jerPTsluxxhlkBTBxNGO1u
QjumoopARwJ1H8ysrxNxnrbo+SAvVTfMNLs9yypfnpSK9OeTkvpROXMAlB9Cfdks
xrL7iPHu18i+G9RGjy0MdXNdT4JDmVQ+yAZp2evpHZe0/WcQa/eF2Z+hoBHcVP7j
VVznrahUemDecYStyIPnYUN7TCdGWSTVozrGRhSTyPxawQv5/gCKcsQAeupLtBa3
2UJTJ1oEunmw7MNUntPhg3R+BHAP3Svq28WfLlfN7NtUtKeqtdeDkSu04Bt+th21
UFghq3jF4zEN1k0f/5fGqImXk1Sa0AWzlQLNnJSLjQEd8NVDBzpvDG58OE8sI8TI
aMq5nAg0Clp9DyrzRyu022TuBNugpymHGgrq4XFxmvBRK/jTFAMEQa3Q0SL5CtWg
T5HdgZaDlzBHNhL8tcF1S2HHyvYO9KPQ3IV0bLSYT8kFafZViU8vBycKaSdecU4Y
fow6Yvr5RGnviU5jFUoiKZ34j6Oyz81ZSEMOePW6LDjBmIWS6MSO8sI58hOvlwQp
0i7mzGL6GR83k6GwVqttGum7V1gdAPO4sUs5PFOIsQNN9s5jCuQiCtH0fiQFoCO/
9BO5punSj/9y1Bsax6zZ+qwb2ws9tBvQdi0nTonWbPJxnuI47UcWkOevJGZOwqWv
Yio+7CkKw1osr2VRsjA4SQdaM8Xi285vBWCqgVaEhtDTTeI72IfXnzLvDbA6cD4f
xMGhuQPLlIcHgyJwE/bLK19fxN9DWs0Qj3BJFvV1VM+bxqTm0E04vCgVg+4sFlAA
1EZrAHlMiOGZdJFmryyfj+inS4t57fdXFLLieGjGrrhx26QgRyAbHf61ic01JnVV
iXjfy3mufgGrt78AWlgVcE4e0H6C2neQ+F4nL2Hb9m1Za/qvXXMGriEkA8g9ENCw
B5KU/SZkBIhoXwOToq+AwxEH7KpU2LwK40cljiWR8q3cOySIKNRKL/IOx/DQVoBG
1WcKNzP2nTjgTyioXt3kc+t42yQVPyOGIGvHaIn0simKqoFpQoUP/hwe5ieQy5Va
L3i8pT9a6RX6Di4Z0M0vu9RisquE6Dx/9xF4pSoUOsjcbfi8/RGjA5XsOgGETkED
kyRhmm9pCDG9dR+cj10LEwMNZLJfr+OAwm/SQtH++4uuDX0zWjT6sVa9nIb0hQip
1Pjkr7qBNziWybNDvu2qXEKPb/4aQUx4HFf+rsIOYK3KfcGSvujW6kRKpdcbGlXJ
gaCyuP3PaOTfNuvX2EsZXh2FD5SFshbpiqTpypXc7k2o6dRYP6zuvYne/o1p1dSs
0f2u+DKpMzU51FkUlqb6N+yIL7K6eYg4HDnCKA1oewFjSgPnSQrsQlVF3nO+fdGw
j0iNFKbN883D/zW7f1HMfTFTDAtCQ4b8wQOBcLPfan3vhzWXsw7jJ9rwYVHybyje
asKWTiYwVzP2e5L7/W217BtzHUzfdXiqIegVCpYnJZUgRGHh3WVPJy+IF+QYM8TU
fPmotla/bCoqC6E4kXS+nxkkUV3MFlGLWPkHHam9SC1omF2UReaHeOMwx4Q5SRPa
5H/hMuhqf8sBtBOsXt2pjKw03Xz6QAJvE3i8YxPoKqKo/TKvrKXeuzczEWvHsDr3
s5CbAv8G2vtAKhwd21rhsy19uY3hAs+U4KefWW99Oj5LOJPYJZa6UL7VBADo6aSt
4W6c73e/nVwD+jAErfi7tAucMUb9xtOEwod4UaO6A79zfrq6nJ8EmTuBKcVgDhs7
jDPJOoeKemocQ/oIBI3l8MjTZhFrL20xRflq87wSvIgTAiFzVIE5QvMvyiMWEsbP
dG1LXLb9ZIBKH0p6Kl8jBUnL9QkVkDC+MowUi2MmWFLu+Ph2OJv/2R2BCdYs3BJh
Wt8M9NUlEJKdKgd3SLuThdNmTk5WUd2jpi2UgC9wqNajm63cLiULKkGPHEEOSyJl
wDzpR0F8PLFN2RT7mm62C5GuoAmrClOH8FEtalHrOIcMgmwhWnNEAI1k1Cn0CMGU
tw2EMv5xONfe8H5Dl+uSHUxZ/u0QuPMSdFPO9ZxkiC/hLgHdiNDW5zeblfnNY89/
NjXwRra1Ld5iZwFb9pgSTi6m/K98G6B4rM5KkMYOvZuteDZX6Dmhy3a0ebdWGJ+H
+VCiWIsNOMWwa6jW8IBTNYYpUDV/bBCXn9qdSB3uLh4XyBz4YnhWF5OeAU7oM9Gj
UIGsDdKm5SRGHv32/uhPhq/mwmsPQvc4PKIF7QYHF2PkIOPyU4cUyMfKPQrjd11N
BfKzUBV2zNUXiqBWSfEXfK+rSD/5BGEWUPW8t6yKI/jFBN5D/dCTzy5Bhsq6LOBo
kCVx7CAtV78i8Mt8CSoRLfJNiEXyZPHmOfNtBWOpblKzJpo+jIdKmKiiis05mX4e
/06Vb7HhIoZ6hGps1Q/ICKoQ9DqgjP+Q7wu7wbFQDky4K+ubksoo70s/AfeSSQPx
kqiJx5PqBbCiSvnjMU5XcisoloxmDQncIXNHTIG4MzfOB1hW3wPsC1/Q552YBOkY
DOsDQp9GDqQtqSh759L3fbpSx+rKMhnIauEwZhw6hX1tzEprmgtRa6Cgz8H8BkzX
/TlDL1k7RR411CES2Tyd7q8+pjBkprb6K6jqCiXR82/lrU1dEWMXYyGjWfWLCA5k
ZqCZfHdZ5rv7wcjMStrG1bgTuvm1BbMb/HZBk1ZGN87nkWUjd2WP35t15KFmlb6k
StzHMGYnfOkzoUiOilzFZBHCU2jdnWVteLimGHv6b6icHbwqXrFH/Y8tePOvsMJw
SgqerWIEGbJMgfvhk2Pe66I3qXZqIJd3DTwIDtpHqT1SQp4RGQigxT3Es5WwHAnD
c7HkY9FqAEFXmGPefgTmLjQNZAHUY1QbNPGH68VVAqxncJh0lT75iV4i9lcWoCok
7pbs3gnhmov7m6f8eHXup0mCkwtlhaCq7R2VTkRfFYuhTuIGsarJfhXN+S1Bmw2X
GWqEcIP0zz+B3q6y1ul/Ub3utgUxo9r+ZjobU062Bm2ufHHP86BFbyUEzV74wiM/
ErussDlAqFWabRn2QyXiub4UiGxI2py9Ryxlp2LNKK1/Rlt4jSa0k2pocFGnT2F5
JR+JIvGWySkRTeWDMFVchHoyogwBk7CyPQBEcfpq5yq0dXbR++cgCAAiLcEuRO2t
+oUYufA2XhdLGb13/bsne+x6ybaYFxtD42hWZzZNIFEdFW2ryWnuq2W/XlyHnvEy
KirfLZKsAPoD6PYJ78YjREDL78BltH1fT4niLpMwEAkuL4oP58OMXhz/20eC44iv
SGl1ic3X+rIh7EG0fbgQNFAnvjwnvpY+/VqF3ao0VKOEJ9IvoU1AvNHDtIBzSv6J
A9tUG+C6ZiubYpPVYD+4PLmj344COYM28sTuOSRfTPOPHWu1SM1aWZvzWgu88RjJ
F6KmEKfvEPM8s8YLIFlcNsMpX4TK2GmgY4JpPqYDragR0i+6yxivG0PQnZ+WL3cz
lUb+7uIT3Zw+KMXdf84fNzhsxi+yp8rlFSkuHV8Aq3WB4cCZjapL7iKMStvk3Bqo
rlp7l7QcstdMLGDd8KK3qRkdWKiQhX7GWFkP0qG/RdHKXOd5hnLzt8fhw6AFfg1M
p70yOTN/TPZJ/emxSCWVuk/ywTySRnqe4DdqAuNt9YbFSQ2STsMn17bSujoNOIBD
C0juL7SfwhQn++1umX3B6JYIAqmgQH4iJammW2znoP+maMg20sG9eym+3mzEieCZ
0CKjJP4ymezuxYX9/McKQhkdylbVxeb670roxuMuWMa7VpTXauXSF/gq0ztqFjLq
OBydJm12+4f3+IqTqwyGMYOD2xsHNghphtnLV6SUujRgCJENu4cf//0V30XtdFBc
8eewvXNcY/gGjYEVF3qFX0WFCk+Wl1wH4L/SBv1H7lnzMtbcD22haxa064LccBHc
Eg8BBDIYko6DHIUIo0xtiTWrcJW4Rzk3D4F0hp5N2e26niwXNYtqeZt6VIy9PKSv
l2nXjHwsILjCt4YSkI8LAK5KyOUFuGNAiD4fKi0Qroh78Sednjai20sDil65kcsA
E8E40qiyqTAqyVfJ08erFuim6apyxx3b8NErdjOA0KfuLE0of82HwSjxp223Z+sZ
hrpkFd+hEsp1nN3tQRlF37zQQAVMVwPWHjE1bWixQL9uu0/lRy07HrKLdF9pgO9j
Y7oXZ0jeo59B9UnfpL1K4U+R7jKu5sBGSrjrP0rpzzEzqScmMKW6m3ITU1WDfufY
3sks7pStq3cDe8kyW0cr5m2uwm0g+80lreqCMgaKwpCWeBzGpIiOSHwquy3LB5AO
TKutqkgQrRnP5hz2/5XdRr5Znls4Jcr/V4FcJ/fHHOZ8pmNyqA1+1UtStl7arDZu
MN+0PQzMHN29vS/2F9sEdVyc5/fc/hSZEiTA8ZAp+o4B33nydL9Q16FcfklWwU+J
gzYU96fA6HrB4Nyh/K9ZmlZsxS8iT/O0DesuyjQdRqi35lfJueyoLDW8/6h+Rth6
Ed2S5tgk0YbthXfV+r9Z0GuUNS/AulC5Kq/Xk3e3nEhWMrHzLA3ggK8D2vRxgOex
nzqgZOMvozX3vYFyyDnIsRftHCz1HouD67g4FYGRrSSGROZov/YT6rKIYgSgmafO
xo610QIRe5fML2RWRFoMBl2DgbMN0ZozycEPkhGqKsA5RDNxnTzlZUZHQ6qr615p
NpDc4H8ZEXesOjaeOkMeafts//56pRaSumVJuv/hbk8Djy3Atk7l0vvj4R3JCRWz
eczP4Mpwa4P6VxFx2hcUcoCl+EWwZ71iTut60ghWIzHGrZ2wYKV5JH2UZc1gaZk5
jJzsUgb76OnOaB1LJb994QXK/ewRPE5d9kf9FlTH0AbNZLzVGEF08ztgAhhUAs/P
lKeSZag78iV4NfiQ0ANEL94Fs0MD6eDFOAG9tsXzx5sMHhG05MgkYRetjN1Jrj/K
a5KPpLQ7vofMAlGxl2STMAVEXtz4hrMqH08Gn9yaUrTnPQl4L7u2WFCrrJBczFc+
6rFvMl7PdvEwJxMHzhLYhEvaBYC1yBIEe37RimiLzyvd96Icf5s1QS0xQg20FLrv
ferskrG/zswBvj5XqkFCLeV4YuVrqAaXSzAvS0qjzG4oVN8MNd8XzO86JLnzWrzK
FC7isnhrbgVqEeF8gUbkMb5UnerJGjfqQAhmedjm1UU/nz383V+Tx6/H6tn9J3iz
PqQfHvMjElhvQoIlO4LhkflRZgDvZaFrrHsl0sHpw4Bakq1y+inBsLTLM/YkzxHV
srMxOCqbVjXMNmJrzlmghKOhJpe3X5lHi37UdL9f1gYQ0BC1B2ioKgnPpj4Vk1Lw
203OS/jgYxBeUwYbulHwYBVOQJfMTgyCQ2pm535DvzQXj0SBoA1lfRRWr4Z4kePM
nXdK22GAvq/iC+Fk5orjx3iqjaWMnlOHHJD1W16Piefct7eOKh7E05hcFqYQscd3
u11q2ttRzPRbsqL6L8k4jh4DbXetr4oeFp3cEBCfMKXWpqwaXmSWepb0oFnAWDa2
RgYPgkpZCnubDL1mFvhAB3q8z6oBhOa6xclQgoY7pGCovt6xuHCORgRHpFLnJr0h
6wDIAi8QstQuDXCf8hRp2ikJXDfd7ReNVP6TAgsTBedo7oV5wRGM3b5M7kzx5IUF
05mL2rRZc6TbYSrBdgBAKTxPW9eHRZxnhls5GV6WUCeuSd5mdJsfIIHFb7wEl+jF
yF7c0wK7FNhi0gSEfUppp3t4kB1zACYKIOlu2SeWskq7TmLgx9gtJxpl9C7pGXGQ
1q/lcPxFN2xal+xa4WyTjwcWRLo6XNOQdxyahrUJG7ITIj/1xqySW3A+SHgUYvNj
Gr7SlkQSBBH9qfqQw9kv+f65PgL04gufHQC3oFlL8ih+Mh+JzMXdryjvkMkPbRVO
0JiQD519PTt4Y/AxkTORQKkdlrwymrRXTDYdlZ0dS/B/r4hGoTb/+7APQ2hErzlK
WqcTwH/3bZR7BzN+/hJZ3tGtJh2FVIcoSfu4/4bvPnI+HDwwFHiKGEj9RGcRdxjM
+QtoR8IJk+WSRX+vTwiNNppebZnobzVtiFT7M4B4BfEoWQISDJ0HadkZzqvLffty
n+jN8cvOCS+q6W3zoklmpimYfdQ8/I1aCtG5Ouyk4zD+ayIhqBK7L1a4aKPbquva
3IlJrsjlUqk6RdwAsY/n58BVYB2LwfX+eQefYRlDzF38NrPz4ECGq6+iO5jmsLHo
20AVAtovUFL9daOygI6KWXyyq2Tu7gYtZu8TKD8UMv53TeTuw8TV4n/Tncb6r5vx
qylT0a/RV/RA3NDmuxkkS+zAxsykk0oUubHCioNzO/hifvYd08Qw1kQMTUtDQPI0
jcMhtETH+vPL8kdWoz1M/btHsCEnsmORWG10YDqTxEPv0K+PtiyI74knsrMJG8FF
L0VaraMdZ8IFZwM447cgbGa92rvol3GEw7I4S0/euP7jqOxeUpTi/TYnZ5CCqjm/
aZois7otBVLj2XAWu690YB3bDEIIVDT2SBuMI1EalLugPc2jytsrUtIS+cERYwKh
r1OWYRUreS2boKgBS88JZlktVXQf36TuyDbWSha8b6aqaZZ2K1ZreNDxaxPm2gp+
lFiQ1WhkN3tefXaH/Rn2PsNPph9P5hy0h3JSQolvGS6m+uN+lP5XsvFOMYCDGbiN
fD/Bu4ocL7xS72DKQIogjcgrEsFo3QLJ1ugOGsLtfsIC3p8tGMtXySEROHzWzXXF
M7/6xJffOcfm3rUCdk4oPw5ZWRfZKfTO0UfPjdFwxpNIkMXZdkEkfy6oxsZoua1j
U1rlmpyw1Wm1GjupQ1TpyqtuMFZeVtLFXrBvcLrfFoN3sUIsA7PA5K932HvpPt9d
fZ+0/t2RO+lolTmcNyQXBhjY8OJMIXQp0zjxZ/O/hQCeFJElAabnBNnkCH4ifxw8
4m9JixyNi9UUpjY482s3qgsDlAvtNH+HC8obSXqWru4hDHA2lk3pgL4OlUSf4tFW
glsGyHg8UOn66s+yF3yveB6vYHCT9VR3ecLj7OtSZ1wzKnxTcVITJ7A9rXoardk8
hV0zb4YObF+RwkswFKMNJcLSbZGoclQwJJz81qQY30KKWDrnWvzb+HPLT8Hf34fh
OYJAFkyV++/J4qu28ln4JVDicZcmCHPVjY6poVrvcRjYhjcdSoEj8Y/VxvKBh7t+
hHN1hFIvzkkQMfBmfzVG7duP5s51Oxk6dpmmxxeYmxvFC61P6Td7ubi5CJIi3hV+
E/Gnv6RV9CsfndWKteKnj3KMwUPVNZhQmShRg/Ls1JRjG9tHp3W3QzEIBQkL0ae+
BNGPkOygNnaR+W5FsMt1uMgDYDX3wecarLnt0YzOUBbn16Ym+jjV/0ZWzOFLegnv
Fh1K50S/uSiY9OHexTCeCBkEtIZNXxUfJnkZVhOcizpuWphiXBmW05OcG/Qq4zTR
aWsuhYPejSB2RLyh1psjt+Kv7CkUBxP5c8VzWyqlepca93lv0LUeE/Wx4yfn769r
zq5QA2cC4Q9CMNRqauFV3iDDzMIJ00LDdaOBElET1yfuh7MIx/ENWUGMXFHE5ILs
q/MdA/uehdg8IyCFfr8GWOFFko4+dPZvSYJ23AsgNVOgZctoesYuAx5HIOUufiwB
of4lRB5uBOkn+6ZkGj7BBLjwU6kcQqU/BVNNOgoODZB+F0FoViXiGy59XY+ER+/L
l5IqIoWjI5I/BjIQ8yWAuZSmj5ZBWJDM3r9Gj1EsXemVuzEIci4Are4dpE/c5ir8
yUSdm0cz9rbMYlaHL5kXjvsJFebM9ItnpW1qixbxN0x1wUGe/WigmGKk5Vf1MsZD
auw+Xw7GeZkgNxN4NLs6YVQquEsBcBtKuyAhEvDUgh6cmARgrQufjDYZnRBwfaW9
QpBXi4p7tQQeAo6baNSmFJ0u1U8m5/CES9KasMVcjZGhUPvCstcMh2O0J/U19DAX
i9IG1lAcb697a3NMV3o3B9CRQjsArOoRzCjzP4b8CUZx86kkQE1Ipdr6/9O3lP9P
Ii5bCVirLRFiQfyxKFcyJ7ybQohIiaW3+KRUTvKzz6fw8Vk8zPOwZqafyMqmOSbE
zZVD3LJoK49uIFQos+E4cA8CldG/0c3RnX3MyrzOhu9+/t41yCuMjXbL3D6x2E1o
U1p1wQ4N38u1NS+rJDuK/TPpvhO44NEKWlsNWEFqXjssjcrALSrRkEpAcLF3JJoS
Us2kq0dgeHlHKt5glPYCU0ESurQ+JPdisgn10IlJJ/NJWCXGg+U2yBwd7YMw3TgI
TWUEWYdtHFyceahMsnzdoAFSq9aTZ1Ao690t7ogryj97vBiZH0BC6Blkrr2ETX0/
Jm/o8bwhBpZS3MutRzLvRSvPOv98bGcjuy3k/Rijwi0SVFD/V4E3Zo8UcciFPOkp
hKctWp5QQv1ysr++/xjh0c6uFDtlYM4zhPzkn5v6HF70Sf76FAHnWgX6jWgm5cBL
M28mOzfgMUfrPpMgSBEiSwr/kJaaja4fbU6l0NmicRQHGSTJepkRgvQ5af4Ojmmt
z4JgIkFHLUfUVdCP5S+nrqp6Nsg6X3wJFsEpK8Ll8tUa+2Kh5kLfX8VNyEBxHlJF
vqO58CoRn052QU+/B5iuJfurx6IW5z0e4qhqkwviZdSNe503j7X8vPxfe0qojcI7
rvZkVySg1KZckT1tPbuQdyoIXB1c+GO1jBPyXI9uEPWfAJDKC0qbhthotYmw/Nen
jLUEf3JhiyLq7r3G5cLvt/2l+kniW55k3LghCq4hk8I8/F+bFQMr3c4R8KhOfL0z
KXTKvVE8TfVN/0KOf5AYwhbocCQ4bbFcW2q2l70yN4IkIEEo4Oaxn9yC3oA6jBTU
EUVOrUCVrlDK/C5Ix8zQTG/C2g5KbSClsO0AoNZY/TtEjGH/FLr5KefQnsgN+82m
xGdZWL6Zk5FofuA1AbFtFCcV3KjP7v07Vp+F2AGn6h61rEIjyqEnplCIjwK1z4zu
+Q0Y+ewMMWCx3PUSRm+yq59t2bR6MWQG75BRK+jW939Jxb9OhJmjZCa+oJK1oqsN
/OXw8wXEkOQ2a3ls4Ka/b/mm9JZ85+cR7JVDyaVqi3so6rh3yi0vVTCrdTKkklYz
IimQqLQN+C+l+vcsz8JSCHvpqx+1MzKwahwnFKn2cNEm52Nyk5ALQ64fTeXK6qSj
1fIP7fbxzheRfGFnb0j5vJ2hXHHd/eWKtcmHXaBNEukfg54L6+coVhJDvrDIJbyJ
hU1JdhVRWAiYFIohwF8z3nmUEImqvgeekxSPYRyq0N8auk+kudr1f6cjJZawU1U8
Chq3ZegjgKgohkNtKoAcAAiJCJzsHLr+wq1TW0aP0jp5wYr7bvkkuLnBKIVt23TO
cDhk4jkEFuVUOlkp+9xolB3AmTfK7uNL94uvQ9ocCPHMSPnS4eHwBefeo+RUlwWR
a+BuXGtjxPSaPzfcmjyEzvhGX1v48b1M6RjW1y6J325mExZX7gF1UAEtM49uYlTE
SK/3G2Hou4Fs/QjEQJB7XIKlD+D1reTJ/f0nuwhUxTE5SFQCooamJc/y7wY1JbCk
aMajTHgpmJZ4ZDt/kkQ6uCdYPbOBO0R4IMVKdOC2vnGupBPQAZ9LZDqDU7Q0shc6
gN1nfPGBDpRJ/aJhEWL69gdt2utXsMDY9SjmRvmOWzQTIwln82pKvBG4noAuKVzH
f/1PWc4pVpj/iOKB0rW0QuvShkhtRDoPEcsB6DyVyJcOHBg/82t12IDrWFCJyqKr
nrtnpiqK31XVCKIIPIU8pMoQCy9IDm1fMZIRgPXA79LZ3RUxWgKDG6rce+6d2ip6
ULq33Hn8ybHKykWF4XP6n6P2E+qiXYVML0E0t0XA0bjUH10xDSKFdEglkm0ChPxn
tnkqW5pRc+f1hkukLwooZbIRX7kAkDorPhQ2yEr3Q5ASYuENANp+JGps291ruTlk
74hcAu6HXx7yalvhfhb/LsitgBY9z9997mM4dQIy1w12QhbGI4Pd5AoVohNMk6sy
DvmDg0O/fT7tIhYO4YOrOXXDFB6BO38Xkjne2YQp+f9nQVa8vAw6GV0+ZSiV2NKA
5G0lpiPsaWzZh7GNeDmdUp+H5wO2GPYjehknpBfVlkKI9uM9Su/HvlzPHEObMqHK
6OfGkH9RYNINLYo2Vs72fonVBPzF+xVaDpKMZM7Uju29OOJ4q7NE2NWUS1sbafXw
omPlkQ/kFmAxESIP8VmAFny8A1+8h516ORPkaQJf9yjzDdxJVkUxvWNsJy2Ticxr
FVbJ5t8F3wX+ROHp+Dt8kAWKmg93Is5dsdj2FcWXjTsgyBdLtNhNluH352Y7DYck
XEcX7zijzhOh/XTcA9WgHkmF8pvMpmD2CvC5jwDe3c+TwMl0c7ka3Tiogs8aqBNA
TKg+4QdCenwaaV/P7YlXW/1pTAiQ4Rjt1AQ1CIEJZZLPzs0w3uUmIPSyAU9rsKbF
v+ZRNZN4oG9kdXE+9QTEs3DoSywVgqOwatbMvI76WuuIfm0orbIRBNyeTpec3akZ
9Bvp4stHGfxf2FVfriPmkXudyYdtc3PvuCp9usiWljq9PwEOI9vbjhxyx2fgE77I
lVB+S+gqwIM2eq42l2JRi4on4whJrhWKIE7L1VlKajOqzCjyX7X/0GkVnJuUuPkE
94G/rfPxNsODOAeFyzggReFFd+/ldKMAu7mpCpFJcosA8hRyWWIaa1eQYD+nQBmo
pGqE0DifdiIJyfJiqI861CWDMmOq3YTiwWBRI+71tOAEAMoS5PNv/4qbGz0gMyDE
MnOMDEDvqyljJO/N6eQ9zpYnXDKExrYNeWydAE6Ek1SGbTPZLvo1jM0wzd8mgWDr
GUr1OePlNjfI7XbaVSyYBUuSxKKjLOSrQodrYCBoSTi9kMUeYeE7Se5111LVGrGs
QJN0xgD6AWVS6w4VBUpTmu0TeJFm3Rr3TaeMYXnY3+mJjYECH/G7jAnMc+cYDeF+
G5b/95ymbpPxgYYZ3jDVcUkjzF2tHEN4rOOd8cf5TN8G9FmEDKgeTt22Ey5r5cLs
GOzo3ibxDBP+OamVQ02EGVCLN/PkNnA2VzwPwUYtuBaXbU/i7U0EZLBzDsaB57ZM
8C1h7LiTxWq6kzuo3miwaAhrtfWNV0IX1KYLbl/PrKQ+lYcIkBJHYqFMqEMYrigl
scul9nvy8MKW+2WH7OaLj3nkC3Db9bBM7qx0kJyU19g3zpcCLSH1VmuBUqDEvuuJ
F/MQnRCrsuDaytQPCiocAtv6jdZ6hxaBGVVPAvgon6TiwjjV7X7ec8VVai94giby
RmtkxL3x5N4sARjA3YO7uTcJxDnVMs+q59vmjP4P+0YWx8zV8GQZinbAI7syrZf0
WspWUgseFSW93cl4wk2nnIFnWY22tcADmiq3dUXmUpSFdgD31G0NP2u7khMDDcIa
X5Awplv0wpV4tRQdsQOZ2K+HZu7Nb2GWkZi8rBnrjkGr/rJ+E67TNisjGkNH58Z8
vgPzWdnLoPB9nAq8M1NzsrcWOmJXUxevIRRk+5js+sS/oHuDTIot3NVXUoUvLKl2
w9nZ08gs+wxxWitFh1+196ls7EpnD0D5iERTfENqzSLwaeK0NLAIch8JhPNIaU5T
0AEPQY71FqnwNu9E0p+BCnpXxPxKAVDyBahZ7Q5ketcqZzFdUhW54+UvQjbTSO+J
JYryLFLoqeEzk1ElyeP00G4XY38JJoU036T4j5ET3Essr+4bLspBKEOG4oyzAcAl
qqaOZp7xR3EJz3R4mAiYYHMEsUkdOzEtmGumcj8tHS0oIBdX4KmL8u/DJMfu+5m2
naePG3EOKvrB2R1Waypyl4JKciN8uVGz/Mc79o/7bQbq+1rFaFwehUIP2EVqc7Sn
+Y6/w0yhh1wRJ0wQlS0AkyZkKNCybu8FGOWkcPtwzpvh2VDsCHKGPZtLHfqBOQ+f
LMyzJr5xOffZnnNIGebS/A09lruaAyIqO84Nm/R5k7z5DO0oF6qGST9o98BWVFD+
bC5r3o6f+Ba3efV0JCR/V41wtpaewoI2+I5b0KsjA3VJJd7JlFCuzwY6/6KrQLfq
JelzzLrEtRkV8WXUf/Umds7L2fs2TgfFvI2aAXniCa639axPW0fUrOk817NUwXvY
KvRF4USsysUqBC9XkISPHLaGfE0Q1vVYNKhz1rq3BS+aMTjWNtbaIxVodIypx9sZ
J60l0o6LFOCh3v9vOHEPn/Pet4YD8tyDuMQSw+yeGU2nmw4eKk6fPvmgaPtOkqn8
4wIriw4v25vRtctkOom0Gekgs9gqNY6YhtTyqABxKlit0PEQq7MioIaMCouDlkaX
Rh/H7TL64oQbvWvU6KvTYZ5hRZQYdLjaHzZmqeALvqR3XbR4PEdQR6DeNvJ9DfIL
d+yCEbJKHWVsGqMAdXpQauvr0VFiwH7H+puCmCe/xpfMTu/G7+MiLO8oFiK/ewK+
gQwGOvTq79yzAnYUyNiyYMim0rxWLoEB41w0f8vbTK804O+59b8Egk5aF439dmvQ
ITowwJrpNel63BGPNqGwR+snCnQNHECDyZa02tW6m6d7VFhHRA5sBqRaBmVVGQ2d
MwNw+PplpSR+C4tEgjQYcjWH1s86SW6QjNiToNs8r+W0dnkVdLARqwhexnvBLvVo
+jruSrWnhxYfIoxUqiBfweG3JSyIxCGVDrq9llx3lXE5FGfGwsP9aDRuaIA8qGrX
g/5prOqhsx1qSRydwNvfldJ5DnfQ1qkJJsFpo6RJHCotB75/ye8rsV/DlBbh4pMu
/o4FAJjylf98lIovdEzmKuhA3wDA4mUmXFSdEX8EVx3LfwOGkLlGUeyvi6Wuy5a6
ZqHXnar9erTBYBtxoBjxuxFRjrqN8hT1qzutkx8X0KKciOU009l0uXun96XW7yBE
ruktvsZlNv5Qntn3M9Bf4tvwxaU7zRAp5yJ4C7FnG/tmD+LeCGKEO/XZPOUO4lbS
vNWFG6WpQ1nZKdypsNUE00/lemU4aoVU8GALILCUbxNWWTSwenFy2Ao+24WCIUTt
qVXJiFh4jKRfgAXHzl7Ol8QKopVhr3NqeFN9OL2NOuBdb3nW9SfaemysQbCsrdQ0
YT9nyAurqqVzLgU5W1kCx/wJQsCOvdpdF9UU8Q9sCOOT67D3TYgm6f+icfgpptbs
LQzD1azi3zD0vNoiRwh4HLxBHgWmZ6Pm2K3CeM1uOJqjQdFoGJMAMaPEZfyTwZ/9
jzT7SRJy3zrDqs4zHU5LmxOZsxlHnlJw3YDnECP/1Lcy3IzURf92unxS5KdVX5un
XFS5GuAQl0peR126jGuzXMxnDQWkN9NTITzkjQwpvI2/27xhFVzDaQ1pC2EB8rVk
H3QQVYAxtY4MC3X6i5qoPugdyYE4TZXzTVPMNIBKjmQDXadA+qY5Hw1UivHUNX7X
4RIlH07km2LvUCthQt0Gd/coz90PtUf52/gnUyhdNrefcnKXMCWpRs4zT6VPXu8X
TyK5JXNl0KrgVW8lYQkAVU/E94K7nRFa72GiJZ2Ao1O5zZ72VSeYVzBaCCSR5E1R
dxSocOnLTpurUOwG/ccB9wCWPZ7+uUZsEdj2kxwX9XL+eu5lFxVQwjQn3Kgh/QVj
6sulDJYj7jjg4+WXD+FP46uZaW5QdufcphvgFqyoVDxnUOot5ExXRDylQEpU88wS
DN+x7Zjmknhp0diipGR93deeNe0QiraQE0e3dbJQu28NxBgPfBVMRcFJ9xpkCJLa
YCsRXfyFrdp/jOstMI0oajH1CTRcQAyE1wLNXzFKFuEidBKy+v9Nk6V4umB+jGA2
6H2CoSWU5x4eEP962UOsBRjDXgQzt0KBOW8fQII/SJaQ4D154vhqBWlmdyJNQpM8
fuwZdjOrF2zy2Ez5Qa7+wDuOiuMCq/jPIVtKhUCLeRo3scboViur7s/wqR1tp388
LhcuunyHwFFfwEcAD7Cmhwj2NaF+t+GbA7eFwo4iC43jROq0kWOCItYdEYttmXZz
i8j1elIJDTjzpLxupiHiG7Djco5Ev1XFR0A7f2BhzD+dbYjPlpdX7ETwFrDjymPe
J5h7jntaq7EkE03T+fuxCY7mdBAC5OZjNV15I3jz6wDGQ/gVur13n9OFO3s5Xd3w
lvqSeeR4d17262MgzOle6KrGJ26ZZ1YGbUNLU4Ocouq0dcj7l4RCdYkpS1EVhGyX
mEfWdAqOwNM7m9vY2fmLpgxELwXmjjLrYFnzyOEe1sj1QdLaV5K4h5LmjQHOBKNw
6zqVPW6G2EzUpk0TqxNtDtDmuutsfO8AArW3xq4FG+TCxbIbtwUFMBe9aWzSWBh1
y2k3Y1ZjACLyAYzb4gC9GUGBWBz/EX13mYeQ6owsd46hqrM0LxedNBjsF/tfAddK
+rsaHbFXJf4YWwQI7ZzAzxjvv0aQ+mianMlpi/N4SrRlJHCmWhs3mwwBR/IFe31M
PJbPI9JdTf9T05mtkqjncUOUJjCYncYVp+bHrTFOCEWo4uX16MFFKbOzEppC32vp
3y3Nk9yS8fi60HHIq+0mbfHdmrr8iB5szRVDETEYeSSlsv533S8FTNaNt1rUlLHU
q3uKSnWKOsUKX+9EZQHOex43+H3UvdVTiefPSoyM6lRtpQXLbuqGSZwG+Q5V1YV+
o8wEb+ASYw5t4GO2+RMyUHNnUGbepnVi4klKhcbKRz1N2rQ6EGvJaXfN17F4FajD
8EQwfYN1WREtl3VPviqnEryjqO9AsNzJFJeppahyi561XE20/Zjm3HtTPAhKqLvo
5ya3x694WitRVTUB3yHM9hmkQsRe9eQ8kXWpfy6VF+JWoFWYjb9uLwSaPcxMZFoT
hRd8qa8p1JXKeTrUCIxFrtsZiUIbVGmgycR0WNN/AoYtKxVtfePj7wy4PIsPYaIk
IJxayR+J+X3PLsiMvfCbdYcE2CRbfvw9q0rNs4XfMsqNYseKbdPtHZtyxwMV0VLh
0K2iX+hLk3IbybELY1XsK5zWqmAuhspp+kYr+aF50HPtHnV01pWhZCXSY13t9SjO
3Uf73pOSRmvQMpGwjXcH/f2Vx+AQ0EguNi+PKjsqm4PM3Mui0GSxUTDbqSPp91zH
7jYVZxhm+zCaKAAWHmpYpMlIcOsP36REBp888Ci3mEL7t1rA8EHNS/E+KDjKSlMI
fTjUQVm7XWhc3lmkBeQpIeHrGsWFg+GrxuWOBeVpvuApgrvn7TGIZ83aVxbu4ok5
Va9ARISSD4tI6y5xNQLxY089HstoFAjeEiyOw3wfZWxiSdoXewtMpjksgZPTRLHn
EZ/AVhdF4ljuST1PHBtz9+z8s8HtSGAiJU4tZ0gcCsQgTGoQox6mFqJNLZvCRZqf
fZmEhr+m9FgmyckGAv8T5ZdQ1jfrEqYJ5wtlIuXCQpaPr+dQUrEseex2PFAiB2Rb
5xG+2ey4xRPmiycUHlicsitRLcofpQdVZaF5pXDIRLY/0ZwaE2guqT78T75x/feB
MhU/+jwzQZibkxqmK8AHJGMj/gryF6XCg1bZ2W4NPrymKoywaxoeBC/62XP9BrkY
N/5zpRshsIV1C2ohlLY6IsTt0bGRBez7rnrIXpF8bfYGm6192d+kAN8Rnh2R/Eqr
e9nkVm+E7Uqn8NtWLbNVJanexC/dbqG8I4v+L5mP49cX5s5g/DewOqopPMjiiJl0
ZU0lgoKy3xEUE25iKDequsmo8Mm2JtEsngOTnOyQdqjV6Ci1t7keUlZ0bhg/jgpq
5AKmV22c1Tu50pkN0UqjpTLLjeWgiFp47lMlorciKsFJ3wmWlHswsHM3rv4QBrEQ
D23TRf9cAmIpxTv6r4xMTNekAMlTaHeevFuozfacgaTYWKlNLBRv7OtC6s6/MBbl
1iREtOPKEu/S84/wMMCmm45NFsd8YcMlA0MJqkRGarzlNC2/xi5jBdIehX+N155g
BAIapZ93q7gnA0DA7hXgT5fbh03e3FOicamG6o4u693E+hXiThJyCdCtINxBqZXA
wahb5kr9DsA0lK7Xj5zhxLyYi4SGJktSCjg4zLhvzRbx/P5kG7ECh6c0ELZkcU0n
odhXF0bHKk1Se03IM+NLuOfH+sLK5wLsCAUcXqdg94TIDr7RvA/iXs/et8wl26On
IxulUFxC+KhhHQk6RWlMWvL2atrDtzXViEQOAFs1yTU8SS5euCF0hEftbSD+iLUZ
+J/oaHIHUk3BfMvausEbzgWgoFsDJy31oEpVVqkRaaX7/uq7g15USOMZ8JRyxNE0
4AAfBVAvpM0oudxIudCFLvYEOomVtlVZoKIhfmbiBWPgbOm7h/pIdUwt1HPUlkMy
xbILvFJHUV0pH6X/rAY0Wo1n6oAfyTMWyzYZBXx3z7gVLgkKa+Ege6fDNHXF4Y2k
Lg6c3oHsW0SXD3Igxpl6Q1E34fW2du4B/4L21i6guUze9VBIRJZtrTdB5WRdNT/g
ZoP+QWtXst/aN3YdBbAv1Lc23A6Algypq4kIR7UwZnRPYmahE82TFsBOB1NLfAZX
DF9yG7B12EwTlcz4X43xMifqEa5Oaluswmyrp8PrWypDcA4t4T/LXEMCCH+U9X9L
IeHgZs7JQkH4NSoH9Mrp7hWYF5RgjFyn5gnBaF5kjcXuD4I9uZMuLw89yLp8yWgR
RWKCx532yhnVkL5pRik3aO1h+zkOdZnZUrSsbsKLme5fj/gkhoZpK9b1SgbLh+8D
+5Kk20HdBcx/t8LDLY4EbcitU4TCmYruEM3MzaOnqvl8Zbw3fBXTx5rihuqd0m4Y
jhAw82AVDTLmRLEPEvaaiXCVLkrdzc9/CL2/2kWj6U4Tx6rCIAQ93x33sTtR5Oj1
DjGPPXUdIuz/JMH0sEotoDpaO+LB4p8hemywb/jqtzUaPisOUnB07VcBpzREn1wJ
jhfNSG7blpdZ4ioHcZJ8h24J6ZTjHGSgdM/PbgYLuMgfHvD90Fh/cxIAI8i/4GxB
JeYRd0mi2ghxoEgbMDQrrWc7Flt09LlmfpTXAiQ7ThR7x+mYREf1cXer7+4RdLNa
Mta0+Cbz/obqo9SYdUcMe5KsQmJ4qWBe7dUwzBwq1X2GkEysBo6SSaAHl+c3dxZG
waGM3W0zActIhZ3imrjP+Mty+yKU8fAL9+GQTltF9ODl0mysjaSb2m6qWh26IHRE
QJfI2qkU1y3B+zcz4WLW8J/LuFBnlMQQaChcoQZvnMZOLfhD6LTLgmGgpO0KO8bb
Ap42h4QFH7elUNZoeoZp5a3EM/kBrrc2BSz1TGyxIvMYjhcXb8ugos+Vc+zFaoUu
Bu6+cX6d1EK3qKuQOp9dVWBz8oXqZRwvD9XMCB9Fh2EP+NeVCTV8z4PY9Mx2Pef5
+xjZG0ucp7J5NIn1RM2SnqqLduqxFNFUpdLWmxRnnMDRrKGk/VJicicq+YzJNGnC
FmrPtaoa2905yqZ2FT0Tpy7ZyouQof1O/Pe4xUVFLsXV6q1Ava9/x6xPGtmEXxjP
VR28VAa/LAgLXw30dXR+ReMWyhAZvEw0iFkiaHg2th6Wrc0WH/LJ8l+7RY/XeWPP
lh7kVcmyZLFzU0bRDNqMPt6lfYkyuHC/MZ24jntKb39DPxU++jGVlNZOfECdjfVy
4U4djnJBKcRbbsuEyOyDZEttvSLX25CFACjhZ9qpIhT94Ek00Y14dzTGl7/iQZdT
lzHncbZ2bt6DOdd7Y5l3gd5CowydZbtLxzLpTjoMYubDz0CC1b44Onlw9cDIj6TA
Phs38NPi0CQ2FHAY47M6AhwxbAXq56I2ojZkeBWOp8JhgVpeI0Zoxj74NxxtShdY
rL8L4g3/+5diX9/LDynn5fwWUEgo1oLehMNndW928AAK7PKY3aeNqjAA6VkQyWIv
W+SM0ti0DjXvWt/Q0KcXaZa3f3kXVAuvVTmMwuakSiTnm+Zvvdjc86xyFlhr6Udg
kJtblFqEDbYSpiuLpjM0675bHV/BFLioPyGNBY9iMwPF3BXQ1Jerj+Ae3bSxiKfy
Dcf3mF5PJADRvwRGt7W6qJUo3DrkAzhT+cuphCD2WgjeizimjppdssiIrd7j5ECt
t27zxq2Vb1KhHUye8IYj60Jf0BHm8iyIrmV1FPPps8D1BS1Ah2M5AtOzextMNK+l
fPQnkrFyfL4gO52J9M8CIO8FEJUhdCBCHXK0+3t8rZCP103dJb/dZSA4+CyzzHQG
j/uBkFeqM2luGYbvYofhPo/f9bSBjOGN3QVNYxmzOmCC2rsS/hcouD7M+/nV02Gn
YjIoc98weRlBaU7vl73lZlmQQF3xuOLLjD89nsl7kajwm1F8Z+MAJ2hOeYz7H4be
PQ2tdWmn/5Dt0kkDJwSu/3sai+r8rVJIJ4WcE0laOjCS6hfIykNzhEZYiUwKMm5y
+GU+ms7E+fn8Y/JblNDrsMb5qQR0A2aj/qtjiK0CGb4Y0JIaIfBBLggJShRErcK1
CU383M4vE17MtKuTnSwBpR/QbnvQUTkpEp14q9emz5qajboDbuhWEsuEnHTmJsWE
DGsg6OZJBY6luq6B3mCRC+iM1Cy1Bc4OYv4sJE2oyVzPILl2DarYREiDZ4SHkOCt
RFX5P0W5jkr2k9O8bR62P+8fJYRlQiGGsiRYFmJeKHROaOuiL9+fqAdqGwJ84Obj
i9bhQmnG7OD7zAZfx5LImobAXBArZgp3GpwYGBNK2Ywydbfz3Y5g0vifWdjKJZZp
PxGDxDMnizqS0G7yjRrmckPAozIzbUfhow/lJYHkYJ09Cmvl3NTe34s6X60TELKF
nrHUr8KSc6urcBkH9K9BGd7RtlclujIY6ZC2IuZo4wbbs3NoPqd+WKFAIdmuQ2NW
ed4CSgD2LjliDOF7I86VRAu2Fl5fX4a/eaIAqCUfl/f7Z897DI+mJUie2gXN0AY4
m4lT2SETw2/xN9yWat+/06lB8DCj745+9+AFw7x6eQZK3MKs85t02VINCx90qpUA
+xCQzpwPxytbcQK0CgtO6F+dWTK14sNTD/zNdB2vh2jLQWwSCi2jxngWqCJkLn8L
jSaAGQk7O6nOjAMPJnl/hAmVXw45SWs7agkXmjPnegXjMCT76G7T6d5U4C9ffNoR
ZmjhTwEbXlDk9H+YIdD4dkx3tftaVj1aXnZP7fKWSPWx+DfREWdgY7UjtQGqf+oB
gr8QzHfoFD9YbVAr3yOFOCKiI1zLaXMNtD+Meg5f8aKSNn3GJi44xU+Rf1jBQEjp
KRwRvUaHeahuK3h/bP1szqDEGfMvSPOQ9z4qU1PhscA5ffAzJBFI3LZtU4y2nTGh
ZdfKvhEL3nlEwEYAN7MsM0s3WRoNL/OD5wYZ2bur8vcVs6p1tXhkB5UgDGV4O4Lx
p99HZ6kT7A57ccTldP0+SxdYXlgh33Fre7fXE++UWWzcR9ruJO9KrCZ5JnT6bzoB
vyQrgOEBODCdQ1nnBMbdbbMkHZr6SmknO9w1YfT7D5PEfuzP3+/xiU0/2NIf1xOS
MVRW6DsOhLgJHMPM6syDEIE/zRxSh/YdQdxkeSlSIlPRYRfjiSy+jxBMWAR9Cvdb
wDjaM5+bzX6zCf9mADamwkCSacsSpCDcsOkOBkxmPouW4GmHFjN5fqPu5iqmHr0P
PzRYYEl/vCTE9u4JQiCf41PhSBDyKT5SPsJDrGvsIYnjKFT1PEieA51j0WQeToYe
9RpXanzF4JBfpeDWP7BdaWAKWg04OuJMHvi1tynxwa+tu/5Aul9z4ActAD97nzYf
OdKw70gu1e9W536kO5vEiUiACQIGM5x2vs/sdEWvFcGilfvfHs+C+g6Sp/wdm6mK
Pee2srid0QMYY3w79ndh+CtLxyU2QUGRd+Zexl0RnnXR3pB7vLGsSbB9rkrYPClS
qB1io7Dp7ch8nbU7OlbAM27qmSswJFeudjia0FYVCnmYWQRm4kqkW785Q/i2LQL5
EEe7tuPVQIeyghojYs9zuILVLwKY31nxoiUWGp0BP99P0VYOOFHOWJ1Du/VsHfpi
tA9DMvwqH9B3aANHkZafy26rzlcKopzg8Ko0l6+MEorIoTY3hyvFRa/PzvQQGcwj
YrdFagEP+AMjdQrCWVz4SRRiyCUIuRnoQHbQtSLiIx2egWw9aZlD3MfKC3jr0Lcv
W0So2YHnXJ9ttifyO7tjHgT0yX2k9cEYjUikxMogZrUehrflanihfAtfC9y8As++
G4M58ANNpf2VL1kwvcFLJV/aA/ttc9/2tQDFfaRR6Ds8WFJCySe25bI462t2EjYF
MrjT49DAjr1FWlq6fwRkKrIH4J5ziib9xNcJmWUWCAffdG2SkdnFU5YF7+7NONbF
HWuM7q+MN1V4767bwnE28sII+LMKyJuP8tVzTgkjcqn1Yi6hqLzE8mG/XTfXKVss
D/TWvtkyHJS7esY6rh/mIg8tYzlZXJjGl9a9WvUX2DGlKH1m464Udva5AUTf9gl8
dowpMRs6T0EfVgSNupOmkQlkJ96ZnIw+iguWnNjjklwHwtqCgek9HVJoo8ViCswx
edYO9e9s2xnmH0gOk6+C5mGVYbEdYAXIHjph4jS0vCrPsSnqGmZYVK146JIePlGc
yUXl/HqnWU6VEexgOIMd4o5cq1piVswuRPitq+Ewswauip0m0Pe3PcBhWX+KO+ly
jTAoQjSQp3jcfJ5AWfYXC7CT2Y2M2NjCtcIS9/+2vybhqVvwHQKe1lI7YLCBpVo7
XefIwf60DmUa1DjAx+5rJvhg6zppgjoJ26tzSTNer7YV3aTFmMQx1BXwYLdVBYzK
vF8gPzXg2AM5pvbfgSZmJ3l6L3vfzFSIEyh6FCMk21FkeMiZoLdSI8NM7F5riPRy
TYX851xtoJXTiaPdRm/sgxY+Nmfln/N0Fv21E+iDD8hYs2YsWn3mjdSJU0f7sptC
ntOIqbO2NUjcBAT5qtSjzDSlki0fTXvJHgThl36UhTxOAPHBTqSQBSvasBjUAL40
qLAdcUqylMUVy952RqrwfC5Xo35ERGlvvVEYO/oekoeuQgtjdh51zoFKddIL6ukE
TCPE9AUnZ25diNUoVlYg5ox2/6Xt3Mw/T1FxtXoJ6nD3J8oQ/PN9jrxlyk/CBugX
alGf58CsL38ehvjFVirXI88Kipz4Xr1u2gopjJjWsoSDjxq7qdn7vnGQVIYrT+23
WdEo/U9ck8NsZxAv0HTLfhVmn94FzfHlqnf6QMX1Sov5hkgU5ys6moWCqAmYZkGP
B/MtwXIipQxOn0513gUnzYIanDmd8UBdT4LHf7fK/wo3d7LxbpWkWLgfu7jOC4y4
id4IXPB5LYmX/Z1QBZI7kSCAxWjo1++OW3eosLH0a06BcJiRM87zUJM7aOC4896H
3w7Vu/3iJMiqwcXdONuIh+LemhRNrJpUQv1GrBGgcX9sx8nRA0EGCz4TqT3lQyda
K23T7AZuTqh8dYyXv7uLCnfxYoofPmUJnbg4IKEAX//lm0H+qHQuvQyl/a4P+MCb
4z6r2ixy/XMUbmAkyMxdcv41gQPx5NNezUmTtKuCbeqtGPqc57UafqkoRVD6zQc5
C4c3VQfbjUTrJtBKIQwX/jRCjDMJVtUloL1rGeDmzJy5P2soQjuKe746Z0WwayTr
CdBGWT4RjeKJ8sx0kMZflmh+cTOobThR7sQOkZ9rLr67yRApBgmDyJjd2+5R0dEq
Gi1mA7t7h7uWcKM3Iro5vJ06mRhHGw6LwywtAEZzwgFRBJlJWBi3p6gk37nWZ8R3
DzJA9Uouu4Eku8pBX9oLvs3NUGEXPjq8bgDmWRjsjCRi/XMX5/6IFrKxX9hM5VgS
ZouAtsaFXsVou66f6ZyDbKHOHLl6VIrvNBQHeThXsqdOEA5PH9H53PDTFpCQoftd
QJ+PfnAVS2/bdDZdCCFEEUh3Y1KSVWGiQZGpwkW69f1rf2n4qpQwfs8/xiV3mBcV
QmjSkaVrcslxLN8QlDKiaPEw8aK+k+ilz9L8y4ANyAIeWJEsaMlMTWzJ5dQTVI3s
Y1HDt18BUGADYATyoGvWaUor0lVimhLXIpxOi/FYeJtCTia+AUZu3Mq9G3W5jh/o
3wrqe5SsdBswnySy4fvLrPZl3UU93rvVrHjQ3S/t2j8+67eBPsSHuXB69DagWoDW
ScN0xV95A3Z2Wvmzl72cVtJnfGTKlYgVGvdhlUG3cvC/F5HoBYL8EHofK8ts2t1i
C3BGV9PLtz1WrmbpJjN3wha3XGATuLQAXq+iewQ7QMZx4HRlz2gYKjF0GcoTpIqy
sXdhkwda5hGcoAoZkm91wx9NzzhMlDmBvcmQbvZBDUKTBbgK0dby69li9F+texA3
8unKdIyn+63gCf8pcYQsZJs0hHdQypQFXjdnrbqql83yGKpOEwanbmNG73T0XwFg
ghlZsQj6UgsI72TZN77Kk6wqBgx6EWVbc0DEm68Uru0ddHlUgYdLfqiIDZ0ZEtE2
WBX71S4Ng5AcMp0oISjQx4Uz5HQkxLfzMHnfhbniY2nhijFTeQvFH9zKfWSjTdeg
o6mZ+vSKk21P2tlJiunFxzdBhwgUkon5wXLmHpUzyyVmOPAwVykCLDom+IqgfT6c
ZjY8p3yTE9b8LyCsYZy6we6UnM2Dvzj8uaBKbZC73SfRpw7TTRu0NYMW2cSz/rYG
SQ0c/mIhR5U4Bd668CcZNfIuficl6sD0rl1qvcmzhv9re41jABEQplrFAETE0Rz0
tSfnNAL6xvogeVo0xT2WkYSIBiDACFUMabIcw+CbP+TjyQXGoRsUNH6FCqhD+RLJ
637yyTfluy3IOl9yfQiNA9/WtrSBYyNTTX/crHoIygSB7JH1lKApl7HkOnxueorf
ZPccqpVGbmdYczn3jcm34Ii+/RABwAzndrsIa7/M14qIPoJI5SuoKvhVgfxMqh+u
DZ6fQx2dXExeEi/6DruR+gm8KU2TSVwZgg5xjaF4s8qcutlwOeWxlSpHefsMnGq0
47/kHlGdObUT3MBauLKzCYfDlIu+XjBtBVRDiVcc5zEM04hhbPk9Rmda08QiH8gO
LBZZFpDds68Q0olIEei+CrGQHLylPqkvXHuAjUzNhuNIiXE/5SzXYLr+ndlinrgl
Cj347nWaEgk8DNrn5ZaQ05JAoPho0qUiJXlxjWlbNoYO77Qz1MO9QJsTEKE2EUJT
+ZqbCq7xSU+msfZ+c2cQvZq5q8I9+KUdHu2jfBezgFmdrZNfXmoGaxcvbWUK9mbQ
1xqYZ/hSgW9FqIy3srn+JcZ9RbxSgL0Cq8fSV93XrIkSeL1GZu1WT1msCnXg29SY
ro3m2vJyE3qtBVfeATvgveEO0DWlS6LSPxbbRsCkRrCCbuGwiX6AIEDYZe3rnVzv
LfWRfPX9DA5vmN/YXEdlSx4pxyvGuZt87MkUdQv8pI9TtJUPknKKAWk3lcCL4wm6
LBu5rI2u2n5EGrBdwQtKl5bKnjiKJZPCNmuz9iDMHLm0V1F6n2kKBPGK6EDxiEtQ
Q0rMJcGuJI5yqE1VXj0hJg8sl54Actny+9gB7qJH2Moi7smQd+hC6t1Up5Eudefi
9jfeX0j5dxRuiRllZlF4AP7w2yf/J1O1fLbhj3fAPNg6OC93wdn9/c2FdkHleTDX
i6oCTPna56ZO7CbtQfigEgr3bP0cwxq5ckTBQ+avXTWHxmKUVgObAhnLhTRB3C8F
JulDWWjj36c8bcsNP2JoGyU+ELLOHt3Nnd0fNdAV//lp5wtxdi9jXGScyQpJNRhn
EdLxkJD4OOTMQ1cNll6IORB+6Z7CHJ5xFwvwdHMJYTuwrbsOZ2HmghXmdmRm+X5i
ZdIKOiahX1xUUCEDkqYQayZOeIHHVWob+oJga8pnn38b9uSfMWh1OLY0Q4F0Vmc/
X9Qir5O7e198qJs+guNJuO+5dhtJ/zz55xzsJDA8EAERY938LzV3lwPnyovm2zEX
X1bsQxSB7OdLWX4JPXVticUASYlAkqXN16CYLstJ8eo2gIVdRydDGkDXXDlWSzfu
Su+awxqKgVxRkr4nshWuHLv5TbABysRhj4MLquciY6Th0oWGU1zubILLmUdbeS/Y
4pVEqjj8eaqGrdoAiDElhjN74invD0o97pLsQC89WEb2MyzDt50/CIJDDWHQJcCs
vm0204uKM7nxHC7UJunVlLeOAuFcfZI2YZp4YF//eSUvQurU9ItXliIQTbfvqR2j
K7NCdvzzKOMibRZBO1TGiQ+BEAogtVUU+DqRXzEtcrVvXEDxeraVxGl/ivnBf4Yi
xyGc7MgYcj218UbrGKHzwoZtDxxrRqNy0+fb5cC4rz3gH/E4fAzq58uKFGpYbW67
9vO0fDBnJtwmxKnwBGviZ0wn+cu7wuzU4VDsK6jwYyr/bKo9mP94PVca7BV4sSXE
p4ZQ2tiCToP/Ctypxubou6jAhmtwkh8P7LbIgFnagxEN9lJ3YVE3A3HU8ZyNOxSR
WWg+SR7bHh9nUj2QM4/dygQVBK5YWLdbaHwIrif4/PT+N1llZ+6lhownLF7VRp0c
5OfJHDIz+BK+Xu/enTr6dJQeTeiQa3HXGnTLL3MeWInK5CFx56Jnz/V/4063QSM4
FED1bA7C9laixaywVgHhGfD9vhl3La67Gpx50JlxFpekvJBfHVqq0o011rkbnmAp
GRfITGo0350kr423fbqnsXVTDycqs5RdO7STuoGBLXpGjcaygQm8T3E6+BYl2JHE
2TO+Hfjco7UWwpNR4WHfhEXuZ4ldP4WFvfoPm7MvDKNYC2tu9fS1Zq0T3ofiOAzr
9/+qE4ejUrKPlEaTOJMvs9a7OJQ+GJqF+a6XHxp2PpvoC3z0Q4DV0vMe/x0vl5Ub
Z6wZ+Nd1lPnEokXu5GaAj/iKN194aFkgqwoNPBFV2znZBIcu+mYjjtbDgjYerp76
Bi/DQHL9MoreBg9jAkIIXwmfAzRdDvQ74bLckEMjv2ioKRoNWnLhDZ0tZtEGn5X9
WZkw7Vb4O0deCHz8rXG+X7TW7rtgC9yHO0/ALcGosOWb21RB5ww5eSwaOZWM1v2U
GciWW3AushluyZS5eFe4KaN1tc2JSOjJknxFaJR02l/ADpSNbqBmv2N450h6thEv
r46iWpX+ULqW0i2bvud6jcgHYDU6OxqUZ9XBq9bUZ5obrSckYSWnagiQugT4fxuI
AmX4g4YYytBGMC41ANXbvT8D051HUqZsdVyK2F507UiuhrzKTr4SJUefj5s7cbaQ
kwk4uzA5AFsk9r0u+O3JBpo+6WwavsO6xQXXgLUk6qhrI6HAPhSXUnpPuxATP/XM
XCeYwiyPxokGgc0C5CnMH3tF6aAWbtdWrB1SenGufAnrJvTJ1/6dPC1UQMO47JGo
fs+SjujvIvhQwEB9YUNk/Mo3JuKPLdH2Y8DM+3rieNOJcPPYnoVEroK1ODrciei2
2iOBxbFB4DhRNKK8OtB1IP1zhEESQ7SVyFQvK4ZvSAEGM5AX1Ux/8ys9/1uvvdsc
qlT5kfHVBVVzqpl/g9YKMw4+8LSFwf+l9sIycvcdpoFWItQ/eVKbrDpQdwnO9BwI
CcjOok1r/OyrTcfCLzeE/4NOGxl1abJ3i/dzuWmeYV6B4AriWIquIKX79hBme0vd
BibWQrbAmx0hGwUD0gOPjzI1hYHQylj/JMvZ5WZ5j0YixjFFQi7Noqt06F6VjJsL
LGYRpcbesLZVZNGvaB1kXC3zHOffbO2WZXKHIXvgjQ7NwkN3PhkQSaQG2+iSUv1e
bAw+2p82Zyql9HEmVLqmk3pQ6gcYuu55DOQqT1y+PSJ+/zeNsShT/z+NsOH3KPkx
XdJYrA/L3Rg6iHzlTx5QxPwW2Hmhym2NQcjlTbGcGWLjHPupFWgqKlXKjxVTk5JF
E5kuarnEAQ68fZtZEkJoFg5oC5XzF7m2xuZ8E4Ni8G+EFjVsBMLgsxLolgRYZdE0
xVNWYFcHRyOVqnpDtRTUFMMIC2aiqFTwmR3ccuHT8ZK9A+vrr5X2s3k8niddLa3V
MyqVBkp9/sgv3XM1IBBnfxA4m62+go3CAKmuY3AmuFvjcHPbfRlGGhflsSf4N5C/
hMEQIkQhGrmZub7t+OhRN2wijg9+TS5OQpqbuBLqvrzJuVqqCbUNO2NLWqM/Irzl
3vvU7KfF42c/sHcyWzZFeOguqgmHfbu4ilfr1/4kPWTNgXb4jBwa8q65ZsqR+W2H
csIlNgNYAzf4atzisCp8ZjIgRpH+x/MBcuInhl3HaSVd/i9hnf2O9542IVzmiNHx
NzjIe3H7I7yTzfdOl4XHWdcEa9zILXOIvzc+ODY4tJRuFYOsxIW1WyoElg3VRu48
bcW4r3vDKYJBqYwIBoXRkgcwf/Cs03fCgppRf0pOo0lMLiRZ7pgVaUCx8c22FvGh
IrDQM1Pyc6XtKQW3+iYKx/MyOQr8BBURt+XvbAYeCCj/AyyuWEyZYAejWYA4N8Dl
Wr1doVfRLHVnzN9n2klPecIRQ4H1f6Nno2Ty24TW3t8LmFAHTZnyRgbzia3tov1r
yPWVTyivUmJ7/QZ+6y/CH8vN6z4zxI57VKkTz8JZ/tTHlWJKyhHWiKz5mk5YCju4
DnRxh24uZigQxVSRDyOCHEswa1GtdrA/Chtf3bSvlqFlT/9TbcBmFCwuDDCA/WRh
Pv6cLX0BvATbEw6Sy8VBpc+FUNwnsqYH8ayyKvt6dFqQ2GCK3Q8mvL/M578r4yvM
xx5rC5EeQkyuTu8ZHwAZ60HhctKHsCE56GGmsvWF1yT6A+2t1x/m7uBT+YRluh+Y
ksidjeQn9f+0dMQFlDRel8XC1n3DOe3hP1/L/6k6kUbSr2/m/R1Q6uRHTiZl2Qij
LHXJsLM+pBHPOjLJrAoid4WETZVZQI38+eKGwrSSYF2539OMJL5EIdRs9k6NxTy7
yBk2S0IJWB1mCMED5WKyeeqI/SYJuAZlap+74ByCcPvWNraK2n9AMwgcRY7WgAFc
YpVtuF+R30n8jjoWqV0hJszG4pifyA2AkkVsHIE+ISp1dGyPBiQAFJIctEnNRK21
ImmKVmljWasBFPe2KwIPBMAhcpVDbN6pclgrV3BIoR/DVULMI0YL+oQKZAFcCGbD
YUo+o4lEiiDf6hSfUSpMTB9hYODLBCdGZWIAuYK/kyDh77MNiOeQgsihuKRiftQj
8MEPfFMQ1a2KjsbVAs/LDph+TvXuVHhTjTZjdU8waJX2dp7IIqNgatXYGHvp2O+d
LM+yS4wFQhjqtF9piC3rI7Dgb8y8OGC/NuMUZrKWP9s8KmN5crMr2/MUVCN5Wx4X
81z09U7Gojl6mtmqFl4EB45si1E1A4jbr3Oxa35vCUXEt/9I6oRXgzTfMqvqziPK
7h00q2Cb8j5hBZDjkMvz7F3czMGYmitU0drT3+wS8E2lsd4YyaTstwhesJzZimkg
qYEHcV4byHa3vOwEJSKvlJ4HZixGjAJAniW7C3tVtqzj2TwdJnaWkjVXm89nfX1F
whV7YSEC11wSRSUNpUQoIYSYvXSYKLkuj0fX0yniKd3eL0R0Jk3gZGifRTrCI8+z
62d529AqJLx4C9hrggtEwx+Y4OL/QziAfMoOVI6yYGpOWoyyvxveJouN+muWA+tq
UsN5G2QO8e5Ss3bdZF/Z9egvMqO4j1Hjhy7qL36AMHc0R7LTpTBT4RiaKfLf2GXw
kQbGCCOYvmDQT0W7S1x2emwqgpwz7EP/JxdA3e9Jjhy/Uv5DhoSx0oMvGa0zUXOe
g33fznYTAYeU7ep0N27suehjTjN6LqKu5LkteygZdJOAzSWaa4jH9x+ZNojrqi8x
OdDa62/PuswJjOBvVtqJsjDDwQEyvGirRQrv4+j9YR1E3h31vTOWzNtBnQAwu68m
4p+e9sVsYu24Hsrip3rvZ9QBvjtlI/umr2JtmxFN7kHJoBF6mIpBOlsqQl9x4mSw
3JNxMq/rF1ddCA3hbDnpWGV5JqxsfyhtDxHsyrBuMU75gc+Ui8fp+uEt8FVPOVTO
5DV/pB6vIn9nfMwlC5FLyhpCwv9LrTO3/w8mv/8FIUjnqg+lO7vQOrz74R3BoLdw
AIj0rbYMYYvJrIk0jeJdEy2TQu2K9M7o6hfujDhMmL1zrJk+TKp3UT2G8sZ75c07
25Z6/Xv4vjs6ULrkVwT36EjRLoDmeaZTnw2vhkd4PFhe1HpWjEEpQQt+XXTTfKWh
K2HkRcsxt0U9p6dN4iDwq1qg6m2IXudf/4WEkJU+8E0UfgigfSTA4w5XetxXZHDq
HY2YaZdP0wQsB5KmwQ4vmivXERx+tAALs/5o+3OF0DWo/Y2Cj7x+7egddTYkwo3z
boX8XD277T8g1IR+SoX8yC6LUnlf3NLawDAXzU+wJKcj1GrZf9M9b/fKAx1mrdZD
L9dI001d73Rd17Rs6i+aDxsF7O+ksorcX5Po1Ow+HXzW2YNB0tneD/wxh9gc7z8l
Or/+0JG0jXv5eMGOLFMr6ILJiKP6Z3Q/z1C/bwNoYj3vSzsKDdgJqHZa1iNQaGfd
dMUB4JNb/coc3DCSoHQMlPI5Gnq9A6jfVhzyXEXrFh/yvkbBJqGfDHd5w8vriPWS
ck2ORMrew06hBOtYQUyvpPzK/4E6ghLaFI3RYnhBLAjYdODQH2oeJ0NGDW0+TDy9
7hzrcd2Vw6aWqA2SdeqgThg5HsUcJI6m6AbAwDwrVY+Gih7BFr+YQqrDM67DZqMT
6vj8CuVR9Je6pAMsC2fvlBB3eG7Dm6El/qlHyh1kWLj16/5wpQpA35S+s20RVQQ4
lN8JsKwpovi20M+3N5NJPhMhrupFvF+87gdjUhA6Pfkup9khtJX9pwS49j/N+UYo
W/qisW2RN9Vsn5pPMmt2jV5t0LK1U+zsgSVMNKqrlW48psPTqzHWQkSYpYKVtQPL
SMsS9LUMi7VMEBOEorIvaDG6382eynkP94PzBm+mGKRkWA1hdDQzMIyKppPTLCVp
xy4nvRXa1bZAGDrY1lYyBndAuVi2d4QIuJIJIaJDs/C1VIup7q4RgXq/z35/Jwdm
VHU4DSJr1jlodFaUwfhWtoNnY08CuhSntgRHU2m5jrn7/ZIFabKSvKgNtDxwG1MV
YYMOys2KSTqyExdmIji3E1MtQeBjzhUvmoEFoCPWTAVsAfa0f8qmQByVfVteDmuN
yTRWw9zLlgusBSG4jI2cP33QfGZ8dj8mIz/FIl8OeapPb/aL6JxLVIEJQScB1rLN
q2LcG21Ih7RKlT4PIDpsJf0CctthkMROwKLDNhwLsdiSe5dUBqYTHiifC51MGtMD
4RwHW0xqZUOWrjCPpDpBF2MRupKBlweLK5UQz5g77V490gT2D9aUQPTmP+E+6f0S
LqfkcGvsmDzXvu/n+wd54fOegoazSGAbI2CZmUWcMjx2Uhjo+5VyYQWxDxn4cZCb
zeeaOHzO7cGyoBgjRpwX2EGkxAiVBXOJBV96svPN1Dmtv7PdeWDWM5gpx+JsChvB
jH/1DZ/jaWEAyWGQEyYZgH0RjQwfGQctXCMEmLzyH84/ha8ou1eLh7mbj5VPsr9e
yu8nVgE7hVoPCB55wt2LoyzO4UYK2r5gjqvq6J1/2flhix14892Wf/Q4KBVdjawp
bbfZkZRhYPqIDmw7mrqiWgkL8CCYaQgWUc2C2vOO83E6LH4zeVKOGESuJCDE/2cm
FwEQJXfWrv0PL/uwYNMUZ/Qnf6k0qYpN6LOM2TJCXvou7nPOUAiIH5IaC/N6RmJQ
FApf+Hhi/wguPs2a3TXk+Xp84FrR7jibfR3tuWLS3FAJinrcv8XWzWjWYZq45CIf
j6dphpkAOshqkdzZd04vhhKxwoLorrKH1Pug3kXy01U6SwEiPtvzlkiXA8yNfous
69LVjwPO6qGQT0G2DnChy2+uPGuhX4Qt5hTaUD9hjT3dAIbRCCD9N4RZnY+qMD2C
/G4Cj5LxDbop6iZ4rVREXwoiAAitd+dIu/+vKvQLbyRVy0yB7Efst3WNjPv5mtFj
Y1zs5BIXHC3t5APmLwDQJtYBx4/tZMEGK07iwRxUmAbAmJEsdmgICtTZOjeOcmOp
S9cJVtPkq0qX7jSXpSttkZJZtHCfzh5qgL1GHSbNazuXnoTGPTAvySwHRYnROgba
CeXLVTY8URWDn/Ix1LRJgctia2gQXqurcihFrvNLZ8UIzJs548DnhMiKvemvmk2X
yCNgZIxfzbmax8vi+IhvB+LkRJ38TxerkIm8Afq+D2SFXtxX+qtob4dBJB0WbAuq
reoAAD50GNxebESUmqAQfC16y5Jv/8Qm4W4D0uhVcbWQ9sSMoWeBF4JH6jYfKt3D
vG2N3rVHTfuEex5HBjXw5Sc9+9VtzCbBoXj/fb0BHlT6Uicj95b7QJE81zl8sGm9
HGNxqhq3kC1DmT0YNNtpf2ugc70aAwMlfot5OcqSqnGd4wVQEN945qfElnpWPMJS
eIG1T1VNxxnNYJ+aanDF2J0g82PJ3de0Ud3NNXiY7HGzv98YPAFkrF3cUnLJsX17
yB/r0FcAdBUH5C4F3xlr2igs6tcr6eYsdUcUm32nSgoI8c13dP8S6hcoV22sBgX7
8qI2ltd56sra2f2NJNsPSdisVn6LHc9pCCY+SI5ms48nG5ptK2jmkA23uSCoeylM
IrTIU7Vd+X6Zz1PfBGy5pdIErnFLK1aw70BUVgnp8r+5GtyEUSAqHFkxFJ3/LyRM
fOd9qivSuKN7aG/cpmNDaW+0He+VR3XRyodK0YIk1VS0DxooMSWydwce3NBaBm6+
JzVXVUc2dOoGSh5Fc3iSGLcSkvw2pjR78vNezNsZ8F3Z6ftV67yJrc9mLNDkgg/8
ZZSaaf0gQ0tJu4iX6tWncdtnoQYsdYdqOcgBsDLmBkQYeO7olmr3wNAi5U4oKzGb
ftPsnFfZmw5aQSDwckXmWvMXw5Rixy9Y1flfcAdTpR0ZoJuix5ceSMBiZX3uh3Pa
UaNZ1MVohbEBcLD2EaESg4APPBiz3NU5okJDwJ0vBwIsqw0GCPo46yOyhLt9l71L
bH61sRtPugNIYCvKMeD/YJiswmOHKuM49/OTk5gkb1n7eKnHhNzBvMRa4YaNC0xk
p0dVcHvacA9uh6JJFGs65sHuIT6z+wsUvitWAZYwrmSk3vRZ0dB3HPlvDPoREeHz
MEeyiGruacIS+ICM1pGgUR26MSjqh8mFF6rCQbDVyM3bQo5pGc8ydrCxctTTvzCz
YjErWcu7d4u4P45DexF95jmuiEsBDfwqhvrl2A3VFCy4986MOiFi/d9xGRoWXjju
wu+Rx+WrVDAlaMKfU0YO0uIb4lUrgNfHYmvOl+LTB7W6RxPelkkycDOCct+mKCMV
vS91W66UV7Kavx41lmMbTdAyzHE3ipugd1aABH2G2pj9x9eNe6fGWRTMuyfop/Ib
jrKpMDSe33VflcVISxHv5EqJ1fMcuKm5jh16o2ZkAUpTlXhYrg1cG1Yf370F49d6
TJ/BBNAcqQW95vZk2aa+0Ty6bm1WJ+tE2GjhVXRLTTR64XI8s6xeteJ8hKq52/KD
g6AV2tGEMvqLPMkPBjuF5inM/Z8k7vXWdBZ+Zc9gOxXngic1p1adMdhF4e2lEp1E
Kgi5YD/10WhQJ74ZVzHovhvegOD9dPKCkjQn80rWWUAZIksM4zS6enJ/ytzacZZ6
WlP3h9H+EC75UGS4g4PpC0wPDmnNpr+n3yHnSwwMbdPaOQFeRGXflQXGGxomnV1/
4ARaBpnOd2xWB1ms/xujJ+UgDB8dsXPtRPZPj2Sb2DDF5n8bBPbIKgHnMb9OwAdu
u3X0hFifHyZUb6f6RgNsj2igjvhZRKp6tm8dxFbb2oZ6O3/+d/NKgfISEwyakKPy
whMOE2O7Bn+OU75H1LPx2eHAzMWrDkb7A19VCEdr+5nGDbIRi9snN7hs/k+UIsBn
uUZt5CBYY8WWeC6nRdmAzNuGAXE706X8feBzMKvnbach+roNc3ktOFIPHw9NxRMU
NafhZPTSQudw2fV6WLyzP0oVN1Hx26GZPQna1MrKAESwZfOQc0rmmN3vRP7ZNeKZ
B3kJrfPe12nQpbUC8WfrZB5tSAT438w+J2JU4awwK3aFM9aZTHayVJBRh8S7A5gC
F3q/lDHMB/Ze1NaKPuGSF1SsR57QNZAP4EmCORgZFXL+uTq1DykiWBaOkI8J1qVX
kFOBnlat/Vh0mbJciiW/eGccWhpZxiGTpOP0x6jwNea3Gn7MPgGJ7DL9x+gydYNZ
kB1qO3ue6cstTdyUtPJ0eqKc/Y7jxPgmVxyE7wIS4klRgPnTDjEaQ1MZJ6e9Hesg
/345qBaGPllzbolFWaw6WZ38K/UK34YFj3owjMyEmG0LW1nHX/qvL8cf14TTXM8u
EnP3jsCmCCP9WFYoNXY1ihdSj0AoYicESoLS4jQHEp+RmyGKuBP9H4zZ91ZNGO6m
i6VVdO/oW4X8vjh0028KFGOKkK+ay6PPf/pS7H6LIHZPT7glXMqISrdOh32IL9+j
QbOy1dUWnppPIHO24GLBrNGfQmBFPDUPtqNAdX0X0ZhH1O7NS+ItsJtKC8VIxfGu
2eNxynFskesy9XuZb4cQEEmdgeRJEJbVrZEAxiRzl7sQ6CT8QbX5jug67gbFn/d2
y7W4c9qvcFxs5SAaKnKCeoXyq+5ycRlq6caXe9KAhN9LMh3tZQyZQN9l3etsuIzJ
IdJLNbnYkoTztXvWiUC2rhYwLU0sxjzggYfifcHf1Ph+9SAdHgaW4cCYGtMSYZTw
pyGVxVf+RzXYBl7uO8irH1kzwXeyWzvsaLeR6eMq/apeeNGLlknRK6LnhYo34Na/
02B/a03BPweoGiEBmaqry19kt9E+zpRXpSHqV7WgHKc2D3iE5gtwo+ys5UTlxDup
qJDOVydPo3+GpXArnvKPZfY3qDRzKWqUz60bSI25v2HV1NzABdz07WAXqYd2KW3V
5irBzlOrppXjZ4GDfqS1VfJLx8FQDdyZeg8GMQPwPXNc8k9zc+J12e0vj6LavPAf
YAiNF5L0bY2R4cjaS9nmjgs/qUwz5akFYQ9qHYPKgDF7/SgmZ3AFYMT2lUpIYnti
3Yf+aYLCRNIMkjE1iMwXjCyyuddiUJwhv/mtqUbcqdse/OMVh1emMD8uZvL/RWCn
ECQlviwMdnUYXGnAI/tXPnzTCanuW80EyW4MsyYszdEx00yz2kMHdBm+jGODAjUi
YhlOHKiMtbu/5BZr0w5E40yE1gjC2EkqylRJkmP4rQUK0Lx8v75ET0gHdwHGjd+X
jAvxSaVTk9V4/Kc+zb4k34/1eWvueoPqMV/TbZXn3MVZcp4fpPXIaJ2US0DvX3hX
zdAglm1ajdJlVBijlMctNZ7Iy6ntPWJjKfcG38NytD5gNkccA2VUmA/WLq+mczod
P1jAptwAGjCY5DysRx4P/sJMPF+cRBDhdqUKvnFZEzQYoXsrE7zRyLtlAFad2h9Q
W24oSPxz1cOhCJKH59tHLh+TwRU6qB928s10uhJolXWSEITJefqXSWlymzTujrY9
a9CjqybDJ32KCaxq+j+PXeLca/PexACyCXy5KC76HAUTuOKPWMyvRgr9bAMtZxrG
V/f2RmjyCccnfx8AUaV7skQJStutS8hrOJ7D4NyLMsvsfzaOrjTexRn6k63+0/oV
rRISpc5lwetM3EOEBJt/z9D5g1D2GxLZQBN/yFLH8BjJeGx7xQtht+VZZMZc85l8
FbCLRtn20ZcBxE2ybZzOJ8RdvVecYE4HHRtgz+SJ5UNU1tZBXffzlGE3/bHZbLT2
Q3QGMTlah8HVXiyNNP4aCzmsPS7kqcJGgWc+m1ZwBoCHEHsx6w8kLekhPugVRgBM
u+4F8f5o9GnEDZNTSIQm6qyV0iP+ofFIZR8WAddB7OOicrO5tjO9mC9SqIFmjeBC
KVaBCnQjYHS5fBgsJUkWEU2+036sg/XCZraNE3gydl46awe/M2P5G7iP1oJwCUhu
34UNE9avDjKRlBNGW3gjIaDP0Q0tr6q0kEHXpGalQm2tqxpeUhT3DqGoe+eb+79s
HbAyI5FWXzvqFetgX2dZ9J5qGLzYSUXYF1zT++ACU/zpgcOmQvfAA6xJ1L1qbEYD
/d6CnEKd7luT9QMIsJASSrMsVs46Bi5dbCzulvUl13DwofsPEZ20TpbDWxWgOJw6
I+3Xgyjm+pf/JY7816fu6ITzrXoIpxymBaeeW2q4O+5f4hClPVCaaNRMaTbWrhao
JmIGx7+XQKN+0pP4/WEk+Tz5qblz6rCVENBIYQkNoExMPpwvkanhl6NbKJoarwtW
brjHyO2vRpUBligcIQUmDWMcesoA/qiYXR39QMl2CuRN7shAWSavACEeUPemkNbH
RuqccMpRJMTPnHI2mFGj+JAcIF3KpbZYzrRnRisazYdrTWPecfRfQlZ52i9ETO9H
cGj9Qi999Hsy+S3SaB9MBQQ52FwUn14+7wpJNtmD0kO6/9aeAA7Vlv7AZhsX2xct
rwlsFh2fKInLrDdL+oVS3WBeTsRA7x0GEzXzwvRKBdkJhd4v7XvM+J2pOc8vYREJ
rThBpXjrMw4Jg+qgm5eUO7OribRd2N61Z8CwJPGNdLntkB5Vrf33SjN/6A4dqLFX
C0sOEqF+bOXYIpfH2ye3q7MdpGm9xGcQnPJ6Yd33W81HJeOLVBksasPdK/AByCHB
K5vEJ4nQ0zJ/IXnVNqjBIcUyGNc5XlPinS7ln0a1DJr65qlwp/blqgFTiSksvDyQ
AEoeV9mFUf8E6y8/Cz3wA+1X3eYkMSSwrarfuxnLE4QpOm6jMREhPh3MZFBMof3K
EZCH/z0VgTT8tm7yICeeMw3+tjTld0jA+2Bf4Pxn71u0ZhJJjzBdIcisSQlzXXC8
PlaxJD6+t4+DJxGd1uhQ6gwdcb9Q14cjXU+yzJvSyUvkq7U8nyCqTwJ71gjJ3hmU
feftnsTMDF1gK5idHd7AUsxXK/c41d+VhUbSsG8hXutmsCapzxyQsJAU1+2+jz+r
h05CX/W/vFRUCmfosnHL1thqc1xfHGH2NO3BFSECCoFIamcLjHngXx2Sq//6dFUa
bo/6TkkSgGHVrCwPVV1v62A5G/qp5Ia/UI8O38MaT9cfwNaFrD6ywGXG0zpZx2Ke
0t8mvyhCeZvPZ5SiiFH9gdx7JyQPuaWFc2oHivvpQo6DvRKkMokAfZBjTDZjBmJs
LLco0vsLXZb9+fuP8sf2JUgQtWnnXA0KHM1JlKon57xs5CtX2bnQ+5AUnSFJbdi7
rsSV/Ms49CBKuWOPSRLJyCNas3xV5UhdiEaITbZnspiAiUKlgl7ocFmZKVIpq8jj
i6c2MBMQ2B7YjQX9cNn2Zl0VaRvTDXccrTut67VmN/0XKgFF5ky7xVzyStKb2bKz
wzuma+11xZNRTvJsg1DdMcJ1UFu41aHJecX/9ccAmFPC87EwmdtTLbaENomeO0Q2
YUFiCi53MsDlLnXdUfaqDBySHT0QBvOFexJPav5+Jq2T1ZlHVA5MSBKk2ice+8Rd
avH+T2IS+bFaAyHnW1b87pTb2M5rffuM6tpA7s6djT4KZ268AbMd3eMw7e0z5OIV
sad5k+61Qc+xUOtHXuH+UoKBsKIbTJWi8GVD/AZzggxvHGfrTPJlTgTm34/xTVpo
ICi4Qy1qG09qQ0xZwD22+DnLLMe3sqOS696xKKsHMBAOaSM01/64TaMyvWhXGsjL
Pui5of4CSkUTK6COi535mfXprxrtFEq5oFT9FryRoOQTG3LKWDZggOqeQTQwym17
ybcZGgkRRV1C4Hxm0LiMqghb7Ic7pQ7DEnsRbgIvqzHlmUqEbLcfvbyBkGUNSCg8
PVaAThIHDr3v6o7XyYSU9EeOSmjBn9A+uhrTMiponp2Cg93KNu+RuqIimz1436La
OWsmKrke5Rb0O+Oz3JBz2+bs3z+MTM8EXaqrZwsPKjv/KWHjPkfKxBD/0uZFiMG2
6Z9mvXMRoD6fpVd6sQ0feytk9VlQJ2Hm0fLFX/Xo+PD7mhW9YAq2hi4tzFp2dmq4
EfD8HbiStGD4r5ai1GsMJIwveHVqnVS6mWKJgO/gz9WMybIWcjG/9SocHCVJkOZ/
r4gET/ojQiDR8RAJ5LDkd4HZy8PXyiLhEKyrQdBj3FBS8ZalFENwFwscSEnCEkM4
DrDMCDWRNBmu56z1j6U0UcaTTABBtTdgsf7+5XXox+LOs7qA3lIVXfBPhO3Sn2px
yShv2+19+NqBDtA9PXNKK5G7daVBQanZZSBpLw0tU41I/TXerDJVzqNbURtbPBz7
VRoBU9F7UXuXtli2O588pEsODa1R4+Hd25D2gwtgfr3+d9vvTcuBJGds2iLg3jvn
+C36XQZqpFpgHvUCadkhrZpqvdIF88zw2BtZ5ROR+bsqCS7oZcp/9aLHndVDwJAb
VfYSwL+UzbWwwA3LNzsrhOS//WaZl4jssdn8JMGamx+4sGFTyTwpRQXE4VXlzjcJ
eOZvlsi5H9csPnjTxWPxlZDWzo67lRv5unH9IDuDwntHxIBZzKe/eAzySzrp7FuJ
x2yE/iY0nzatL8aaSR6Da2ZGrCYsWb6PxecxXjekyZ05lauGpP1klAvI64Ib1vMS
NYEnRdjOIZBcazltZMUQ93jYjriN2+f2b+pvw/GhaLvirPp/sbvf9/sHqx3zj+J3
oqPuXzeBb8NAlmCmO8l1+c1fGR4FzQGWUlXPAOuNWbdvNJlnbQZueG81WyBE0lkS
cQy4ov/ZQqaJ9UxOn1bAzblSSpRsD09LDGu8x24PNlaWbJfN7QF4oAeivlby086D
J19tsPDTbKwPHkxkbf9wPZkLOUtk7TKABQs54JMSxd5HRG8qEzg8A072aoI4+uZh
6t037lB+W9DTzLjV41Mt4tRgur/DWpEhiJVsxQsHTFKLRvolZQixrKsdS5P/t/qJ
xrINEFUHhuU3RcqEtCToEvaFFhCsvoFGBgVehGLyhQeEvrNxG8SpNXw9crkaaTV8
SRPdYWj+I9dEvD1w6cBAHNDUxqfccTZ0xqf+E+aJe7JqXGAmTI4V1JkT1drh90C+
XzM8V2ie4cbHQFAMB/cCxGVDi7FlqEfNkybmw8tnRWWbdHS/lT9hfTPs1Qjz71Zs
7jvCmq+elctmVpEgr0Bc2wSE2WKKGQDVMUKlFOXeZtILO5biok7f6ha8RSEp22EB
LSWAtOZO3mxzxz/IT7OYes+wdHi1GYGchHLo+pnOU8mhW4bO84dd19+FIPF2Xjkf
9T5yE/02B/STb4mPiPfdodCLYlFNlbcSxc4LDOuTH8/G/GB8MfMO+qTqdyDN1vO0
k108vNFSU47XVzrvMxudbRiGqD8/aczrj1xmQn82dHWMg0mArPMeyzw3m8IWMLVx
UenR+rp2SjHzZwTkDmc/lOEX/JTBQL+0FveLCpgccl4D99OlS36/ZZsrkVHzIpjs
6JzfCJk8zbLkYaAdJ/OeUsmCG8FosyUkvS3oyb99UEvS3y36rRVwYAVUcmUXraiO
xsFioYOipK/f8v0hfZqHpW2O+KMisNSnjfk8AsmqdS9KJ9ZihzK4suUxwMAJPy7i
w4cUwxdkpGOQBt/8WJGbpIzOTK7LNJlFAs5+OkSBRmfctEK+WJXCvy4U2hifKems
7P79U7RjTKv3cG9mDH/72k8ZFOA2BFkbstFv/p78wgsA/hjyEbhvzfhfggVhb1Zw
2+2S7QWCzY3GBp2valCOJmJumag6UsTwm4IReJ85W4nHRLPfbItW6+Lr/99qY52g
2+2k2YmIUNDSRc+3Wnels55x3dlWtlgkosgdzdjoGXiCXyFqK7rQflvzXBScISkY
/UTYe8PN7eEIoxI1kPDbGHu7wHdy/ZRiBmd6hjrlFEhkNVo0BgsnZzExwMzxBZW4
ZUMeuVQSiSiH9NwGIB6Q7PnIftXpIdODBFoj1u0v/L3ArQbwMi+l4noWtKyS0cLL
7S/vKwz/7Tb8EvpEnnryzyJxdf625UiNLuNzLe266ZRdZiq10KpTTaubtzBF0iRW
/wr1aH4Miuqq3KAIbgBH4qXnIfHFnmbxd9pPPjzCJpc/JpyujNMkJZ8ji8tP92Wn
rnGPSfBs7ChJSVGyB9t7thXuPcRvM5nNgmNFSwGn8t1tQM4PjIl7ptWtI+MRtHp1
eI9ndhTB03sqgK9A6RMLIUTo6A2CUYSOv864nvJ0xMdbSrXdaIqov/Igw7q1hEN3
bA4D3UcPE5q8F/Z9JMmyE2v1+km/J9FrBQYLHTnAYlU9eiJFgoZQ4bUYPsvR83tV
PAUQKhnVPL0s79b8h5WBszbrpuoNmtuqwp8H7GmvQXHJWsJ6C7EOyY1Lgzk+GnsR
PBSW5aI2RxSYyFYeVzW7iiSTwMHkWXrtsiXdQgVRWfnZaSmmmlKhS8bOar7WRBJc
rBpikbMf5pD4oFbUKfCmB2IDTJxXsxKcWYxqhuNP6vo6rZu8UNstMq1PxK5LLll5
9cwtW663kI3hKabbMS13vWykoKLPe/QE3LEFJ9iQTQX5eCfLYcCJGLrDr6Xt3OsT
4OlL8ZqRuuZiYPfC/w8ElWSoLQSykFT+S3fvZ8hIASLOYG+xwfsAPWIBdwiIHhRJ
8zTCyf/sHQGIzOSlSGt+tutY0qtGdvud3yCB5fNI98eLKjajlV4YUMVnqjIc22up
FGA0gOhLjv0FbaytTTcz+hZ5X5EXD0ALl2QkBV3iFjjQ2TfNqHdFWTOzWU0baPN0
4Wd0yxlIIOQbc7ZASOFOwIt0xlNYmeLl+OkcvkYCu+kLne5OQYUvwKIeRj6kolEc
MF2BFcPVKLht8I/tx80Mi8AkaMdsYeSc0JjLC7NXTqKIKXPf0vI8/S3UJVdAQgFT
QhTyfEDyA9dDnGH17KwmR39pehOihJG3+I11goq4cO5TpdppQuYdhSHbVQ+6vaBY
HTxgemC75RJ4aFtltxfpnghTq2e7DhmT1FkwLGiWtomIhA2wBI2aOjHoXS/eiudC
QAJRWIZlGKqAhheNcOpAegBfyTh3VXG7g3zonO9IpCHYZoOdlNZmYgtxUVyej8ZZ
oRSEz+h7lQog+A+jPShmc6iTChbnrgnwe7u17AG3flcWLyLAoCmKCermIQYPZe5U
BCv8AJVmKrqlB2pV67KlKWl2a8khjEbwfGVkjRo+BnaD7gNoT2AgyjhLAHigs2xh
AykWkKWEOTavcii6Xy8KGSE4dUUjX+9soSxtchAwm5XpmDANaRoXFcpFcjiXKC10
/wSpsu0TdZKfktqAxat2PNPV56OsItohc3hJlcRHT/i4FLa93kR6/i1s6dlGMjqH
hcdY5WWeOimvnmVhMXymN3C5Gc+JuPrTXf084KJgJRLJnVSTUMHDtsucmYBX/+Xq
hzvrMpFAKos6slnqhtrJdDSvUN8tCOOc1ojTyryLpYmg5ew0Pgd2e9+eIJEHEosS
SLjUXGBBxEyxgFvTu/V5rJipVE8tpyDzRWQt90aXE5nOIWrfB+Z0ngiZqM9Q7kfp
ruMmRHuq4oE2BFvYtV0+weiuGZQ5bbCwMVhLRmXUwXaV1JWaKFRM0MbcDpty1uYf
UTIw5qDxi5mpKUkqqrPscXlyT3emccNuhHXbRMLXrJYDDvbi8JPvUyYF5/Ip/Vaz
pkNrZHw9/mJjaIRpt6OE5IzBxyhzIrjBUcX0FNXqG2X1techbkj4w8jyyjeApZ8t
ccHP6k0UBt6W9k2dDThkf/lOBNYGNT7sTE7K31dOQkwJVWpcmSluwiM43Ew+HYqB
wMmQ43qVSCrgwIoqO/ooFW+8XTUz3Aepn54eg0peu84MJy4vZeVzci1ha92EQ+py
mryrq8okk/1ojEKuwEVi731nNZXcVHGoU2gn2ktQ7RgTT+4ZdxILtE/BBVFaRAjP
xH+zTEm9/JDPU7lH2U0cvTKHEPSuLOEJatZ6/5k0TmgJJZXKui9qCP84uCFiMvnp
unHzJZ3PXD79HyyMOvzhaeC8WcrVW5X3cCS1EVyVRvV46ea+B12Wf00aIda3bevn
EdU9vDMqR+8HTAvDKuVFYF4I9x83AnosY1b4nbWpHXKWr6gm8nPDCB66W3F1GFS/
CjZgUk9FMLJqXRKwcKmDZQ22V3ofAw3Ye2gytwet5/2qQlAwTmsLLe69X7IeUsYN
4uVuENQCf+FgxhEpso02VxWA/H3S+C+JUPSJodlG097fOhrND1yl/Jg1pP2uQSdq
TY3FlpKT5T2l6/K487ApvrYnIYHFTTztOuiIzl+eVYkAbLIHB4dka8DH6iVwtSG8
/3/w0iCkueabUDOUU9+2OYo8/sbqWBh5Vhbdc8+pYuBPQCk6tWc19NZjIsOGYJZi
5Xxuj7bdMMXXuJ9b/jl/UNHziU5vqkFHvtU8hJ13PLQNY0xyPxB2m8MWs21/lQ2I
Drse5bSDbjAvuKjC9b+9nEIXJyhSBcsSDZqtYxV8uB5zdOaIRsUfTVk1cWk8Mv7F
fKVrq5Iqvyo4vUDXXjbHPBAHWl5UvnPfNdlA0G+FjaqYQR7ikvKIpG/hl6p9kNeJ
+KSggrLTOFPxQBoKpYUUlEliUi0j5QhO/PQsaSHN6Fvo2mrxK6XViwfz01xbMjvP
qL5hjurCyLQf7uGhGybsEyKPEwCwU4l/+ibuKRIukeRMz3RHvJWBkSU5ybJho/UZ
OP00CAbJmkKRAknh+XVklJ49DajJnic9TLjAA2wensDNL8+Rr51Xw5tkCUCEQE3q
WIZ2giYh7K15flwr/fwS6qKSDEixCxEYRVKIxD9E1o7fd796pQIgFAa2GhytqpRy
Dy5M9y6L2GN2TL52LUcFIlyT3U4Rll+ZeCMeBXBWI+tnO8NupoJq4Pnjt9+BUGkE
0OXS7fxAbnND9fTBAyWdz965xrII5QGMCw2M8y04abmdCw/emeyUUZDuwdlJ2KHU
7KeVXgLIHJwhZJa5fy3/vVw4j+dRGXvSe5SSh/JqDp3emKp/LgzvCrt/tSV5UXhe
WPOz6EFTl9dc7cypbT+LDGKvNfxSqtjgeZ5LU5VnvsbGdRMIY70ek0Ynx5xyisNp
Ix52kBzk/DT/YFZ8WK40f34TX9HECNlZRqT+ZKxeCS+GtL9WTchx1j+VFNHZGhiG
LWq9KtBOLLKCWlG2bPpP5jk0g6y9TqoYYpP5keCjhn4cs5/dWt1oX2YYjIqfPYOt
qUx4yOttcVuSCCAdCn79jZ2kMUmc8H2dpSp0MMbi/73a1sVPA8SL+Msp3Vq7cpUA
LQLpoIExEMyQmVDeHHZ8G5R9s4BmbSUPFTS7XgdWIiUetMq8WWRQZu1wrdtnv5XG
r317m8cOU+tSqeNfcsGJkJYHPUsiIOTY+5/v+7vXPFuWIXTSdh/MK8Koorci65PK
aA6WeqjND34+N4wv+JIWCSl3FIqMUEjKky01JhFDnXgZ2OREfV5sLPwDyi8UC+bG
LovLP7g6ggFrxTyb6jA624BFyN2EQTO+kjx1B/sAZHYOZpKkdoyvexSjH++s+vU9
WfNM5WxAtFrUjXGPz+CCPbKrgQ6Q9w09FdWfA81lL0WsdZGCFr9r1rEogj+9uNrk
SazMvc6YLwKANw1pY0t6G3dDLi6ppqkoyO58OEr/0ZtfZD8tI43H86ETeO7Jpczm
xrcjumpuvsS3TT7fVyw+AaTtBOKY5QBkrLfP/Y0Lbi207MkvAj1Oym56jbgZbBzU
H581Z3ZmNVNKv9xz43C3PiBdC9op4amA529pib6zL8fOOfbZ+CKTdWx7Ahua3Dpm
ki1JI0Fp7uvIyZ6sGzyeKOR7QYeYG7rK7/c/STkM9RQU6eaW0LSaVLiVIzgH/nvq
ZG59njmfRTPy6E3I26hYVy+wYClfgLfiX+zV9Vrtp1Xa19zK4FsdJotHr/i3rH2+
oXpLEHElGJT6QtU2xGwxYORs2gpA4/QACYiKWMi08EzhYXYugfT0mMDm1pWCCuyg
QxEeh91WBdesTlOPXewnOFjXvCx9uY1CIEyovyU0r5ZvT5+ByfSgPpxp3ppa3UCQ
0gypdTekG44L4Ow/pckxzdXHZz+QznUfez1nvFU/WZhe78n/ZpbtajzX6ik3ujY5
FTppMWalhWxKVCjT4Rsb2UTqyETHOd8nhMTtQJLiunyq+kUYzMp8V3m+kAj0mWH1
PFHi1Kaa7LZWZJj0da85DxiVo5ZXhaBWB9AVcTPy9SaU88/O0AovFfexFpTElZgD
tF4LBf0bfOUfET11CAKDrhkdLYd8VSRVZpUW6EAuVjGAaV0FNO6IX9t4FXzr4YDC
9Rslfo5sldz8FhLVDSbI8Q+zGObeMnaJclowNleEv1qt/XJOs7mJyrbYjMBNX+m+
HFZZ7DNwN2JImW77jJAHhX0IgTFLXu7PN3EsLLunkZ6rMmMwk1gLFUr610RTFaaw
wx+VDBQWYx8p2KamIOlf5INwITCZWJhrqNLEUtOdVM8d1L7ziUYoA44j0EqOogAK
vs6d7YksOvN34l4NBMxYwcmARtwrnWFcBMPzUQQIqiVJmZUgP7LijuuChoeL6r/+
pF2i5DNuFKkXxgQpXIwU04O9EaqgCp1FI2lN8kPaodBVr8SWCog/1RVxTgQ+C6r1
An6oRWfZ+dyIpyeasyAZKmEnKM/Eu4E5iLDea5j6685t5JLJGgaE7kdv+2fDppGP
n9E8HAEvewLcpsFVzliLxqdxL8gzCQVxRJ07Z9I1El7LOPk8Veyp3iF+g/YaJTWV
bz87lFl8vT3uHE0BpgfSM0LK9hK2JXri9eqRfWNOsiK6Z2z45ZAnISx8SbGXXYzB
rfmjXmJZN5CXJIJHoWrpmfIHASdnNI576VnVW6fTnA9yGQKT7HZkGjVUcw8ZmTYl
wH3VjnlstjK1FjBoG197AGQ8nUvCSFSZB4bGbP5FBuXK4jD8AW7rHcWn6SK3TGC3
ghkjqWiXOUv4qG6DhYYsm4M9KfcZNCr2bu7v6vNF54GWX0u/E3yKArJbp2arPSUR
1Zl6r1QnvholEtjAA40O7ijeCix2Bk2dsOLsnJz1ukoJ1TscDAfxkfOoA2xCIHQb
o7HBQ7F0paRZWfU7UZe2q+kc9TBu+xxQCX5gLm2eHw6uVomkdlh5xSoFrdRGo6V4
u/ouljRLmSbmireSOy8BO7jlymcuy0+pvW2JEtGzAsxVltMbmJOnbmv+xRq7ixtW
XsYf6lbZ80uTSg9suw46Bzds7mWlmdvKz2QgLfcFZci7njzAkQtsFJx2kR4mAv9n
40GzMJQIe8iVDkn4aGASyOg0DXLb0jqAWQVdR2UmjB1mwqehS/DCjbkxkp1QXBUs
mcpRzOhuTGo6BV54plUGYHUnHPCx4Dd8fZttuOlDpDNXSVfGHr3Jxa20TSvNSCKJ
skIdhIjeTgfd4+vKDuUEK0tr32LdIm+Pv2N+NQe7zOH5R/jqZaNeX1nPKJbOcVoT
dNczebV6uQnrP8E4t2SmO4jTZsCuRPIJlYruO+1uBoW4g7AcToF2z0ylPfzlSmXY
5bKBd11k3ZaONvgxqM1WpOnMG/IwHlTqzzy14YHZdRI/Edx3vNIjliYhn68uI1L/
Ay9opceegr2IFOhCwXwbKmZrIH/Ku5tRApTwHzSkiZ8ZXasUk+CdDYIRwu1qcWuO
K8jOurOr2oQFqMTjONWsTqsZhMSnoBlaNUV/E2z+T4NLh4UVIYcMmJkzBymJZcbH
TMzkwSmBZsSPFVQFYucBtm82wH/omUnPAf04BZk0Frs5K9lKiKB+LgLDKPNPXbsx
dE84H4A19TGgWJIqpvLu/Txla/DdJiDzTUXnW4lzlQHUYsmK/asUIy4/0mCbOaHW
LQYZTS+2wnCX56USl1dCegyFsLBYFkkoN3t4/Mswgwj6GfO7JM3mcQbnfMxYeI5Y
wl66jKcjlJEK3vimDKAr4ufIrW7bg0M0aWhkb8XzYn8hRa1rMTl1Q7OWrRQW/HTn
EcwjoS0YO9L+V+SZgz/ZFFHL7gDaBVvjhmC+r+zd5Y8xwrhDE8AbjSK9dTpMRZyn
NWr6V8o3JnKNq5RPmLl29e5oNSlgK5yYLElJgIKrtiYznfOzSnNqz6yQVHX5p9O9
pGnaLHMJcoTOT6FZrkBH2NVQTmCAhvAp37juOBlGBqNsLL6m6nMKjgqkys00k99x
C7j4//hJ1rAraMhxNVzT5KUmP05QJSb9UnbGA8xQe/omZHM0GcsQ/W7MFxc0iS30
utQSxpi6VQsD6W0KARnnwG1905h6aYZtmyNjvUCtjZIjwMLKtPSpEzkLHDTFA53p
lNkgK1KijBLyECnIdj3t1x35HhoRxS1GXbOguTBPTQGSvhiB/LkV+VOdwGhXFUfR
b1+U+6HXPbOGjyqASCO4uQ7yXMGCq3SiEL9fkJ3BijuWSSeEwFvKHbfdAGutZL5k
hpBkw+TRcHrD3xtaDWkBBVitIu01r7cixS3xQv/FlB4cY+jKQfFDTQklHLGNvKtp
IN1oiNRra06puvacynK5+6+9ZDSVWLjyMr39bAggXPDFMtMfr6SvmJHJUyDX/HEV
ZstBAibrOBtGkU6M83EVaShrG4Y1XWr7FDqhvPp1INCaFWEYOIIyqdHW5ojPnAGS
HQgY3jvPpafFa1AuBWZ3grGTZVXXFwDGzVxX5z8JUoxBHhYC8nI9eQe1f6H5PZWA
gHC5bOYub/cd42wkjF7wH2kYO6kBeglATrs2ezOjJedSsdk9vxhg7tRzADGf+rrK
jd59lEWGmqMSpLFcfxv1tmdhC+cemFoHYMAPFaRZexS4NY5EztKm8xdcqohoN7Mf
E+o1f/TywD5VIGhYOJkRsPUmQ+Kz0xAUc2R0pkzK4UYJycj1jknhU8SjFxifgHZ5
okCi7mzcEcRx/XkBO6VIX93w856QgH/KZegxheDIB3rU7V+RfFtzWT+uCoyiMdNF
cMyBDaG4AMOd3BR+lGLhXJRPENdq6XLmrhGzMOx0E8QmcG7HXTLed8zsbPkDwlar
PoEm9GkCozehcRZRS0bkKxMsd82yVRFGvURS7HmFjGWGSU9oQxPJ1s4LzndzOSdg
oxpsxAtAYt5aeZsNcFiwWTjNsacxDo8BUO5i3/zg2b1Qc+N0xIfelCMXZeoQY06n
BUgTqbcnvOui18hby/9M5S1FfuTkt+cRYyj5ZAG91ZrIyku8LqjEaLqKivFk3cHj
0C9LXw3M1cz13HFfZdTlROA0NgSn59a1vV1KsuQLcfehXvGfg2V6zc2ZxelWsORO
EjkVbBzC1Ln+q6hI23tqCodCMfkLZApTuYimRRVa1KJ3UZpzbiHS4G3CirdehyHd
lU7Acjr3apVRwDDVIXcJNA0+4yytNXwiIYZiC29VkxEWiSIbMYR8cmfCaBJnpw3b
p43ahpb7PWvRBHDNDLeUqTHCdPcOSmaLfa16XQbN4LSKTYY4z+5n9W2UbGPo8kQn
V+2lLieUDdZUa8b6oMPbZvlicJvf6iDBFGA9fdAwzpuYDK1KBL7RbOitzpB83iON
mWVabPTvPrLw5oxsdUXZL/ulP4AyiiuuHGOGgCPw/vkdfveV8t3xkmch69xyHB75
Q93ooxIFmh+u0zVvc1fxf6KUkgkogqD0exOJQ0paFhsQv71plOOwnJI8jrmUwe+B
cZnG8zXui8QvDTekO56OtJ3eN+ORg442hpDdsGGrv+n9XH+s9QW15OHBDjqkuZ2i
9j3Nhb/mnZFsP7OAxk/cMlkCEZEHTOeP8LRrijra26fDRUAnyxc7l1lBFecQAlLy
eR9JB5UyDH9Uu4HHsoIXjo7EqioZl8BlM0E441PhGZIC02KXhf3hz5LKwQJyYJTl
h6mTeYEt7+7Rus49QaJyLaFG8jVSRzCpgybBqv02io/ZCvUor1f9T3Gs7vnru1X6
d6Lat1M4HHwHO95kkfdRooBLnHRsFtJre0E/xlBz0WfwCwSpqNf+k9yuAaVBHUMK
EwuXDTZ1svMhsOYmrh9SF6l9UrOKi7SVLTOHEgXMTL182CEJRN5/wkt3oTYXebCo
v2GNO3kxWlxBD10FX9EAr6nVDmH7c2o+PIhWXyj8YKBSan7IQdaPsPthYgbD0Om/
/D9k09vGTcBZB2vUxDDMPqM7E6vn9seWTWIB1c7BXej4FlmKIxpbIAgXid0fkeN8
eIglYvXUNJoZgloEhWgQpcvKsq5XFuIMwV5WBH1nBnvfUSj8mwItk6ZHT2yfjxia
F5/4qMTdXSRK3hm9h9U0WcIr/Tx9156tejM17Ax8tSf/aobPXkl+Y+t5Ne1U9DEe
/ruy/TNHRomXqzreEdFSdbhxJnSO4H0SREhxCmCYHp7rVSj0m/xK/yigvBdduBJN
iLQAIZeIQ6GABKaSy30YVdq9iYKbqDHJRPQoZOVZZGM26DfiCV7paUqKFNCr8jPa
fp/RpWlGH7ypGNCAZgSWPVitoqBWVaE/BIlMGPyGWBMsy2ANnfgFvxVIFTIWi6Rs
JmPUtQ9jxZbCrBSL4pfsN73VnHR1erfFM2Rqvn+3D2rF3gmP9wC8dIzpEvBs/jOt
OGrT5qer1mZFRCfqFpUKjs/VYG4optnPw9R5KGiRkBaX4fHMf6jVbECFlWuINY2c
yvdlf0FYP4rN1r0+onaBBCU/u/eUMuK4CG4+c2bdg9HGFCeBeXWFltvADp+oJqBy
H2Wqg7PEqiW3glkawjJvwPa4ib61+rpG0rD2I+fIZS3vimMEVOH0ZrAG471LOKG4
C9SbQIMdZYzBu0C+BWJhuBKrycGYM5kFTT/AkNMQykdl/kbj3q0gTONnmHJ87osb
DipCN9ADcY7OM3Qp3/SbQqwFrKSr/KSbPMIVvm0SJBtR/Orfo0ff5QTTg94S3AqC
6u6tCZZroomWMx0S7qBrcqzQy58uODytoXJOSkFTNv60gina0cAYHk0VbrkXB7zu
zjxBFIYxc5QmFhKDdAoNZ5GHvKksU33gpE39ySFF6kTLlm5ZBR4mRkpdaaeDoE3z
EJtkO32kAPgEerVRMVbkh1wUDyG4YbbLpkzXM6pQv5BMudkCJDGwyuf10g+ymxyq
kFCaU0gKq6yE/Y6JdjSEpUWVC4XXLazqVo8aFERMbbAbiIXMkKsnw0HAgJWsiMEp
kTlcV1ZMZ9J/RZkT3bTqaBolM9+nrPRh9voMEhCLD6p/UnHzIswlbRpaZ3BCHGad
AKgmNi7AW3HSk0/9V8s9GbbfQSgWlFXqO8BOlMpo10a7fNerDZJixGql4LtMGwKw
2CK7d+flxfn5MOY4jPUXOtJkFzJsFLzN3bZ25voE9MBz2Gwig5qPNhxBDHg4abxt
yFKn9qNlZ7FSNIaI3JFZZh6UPs21evFACS91pWIb1bxE1xOOygS2fakwopyLeJiB
C0xL5t+DnvsB5q6BmkhlJLmxyss2P2bTWu3GXiJqKBXVsQBCsoSKKvzZqfueV7tc
mJlmBPvX3hVUUvkseb1CGQGxaxApSIikVyMtyRvpVbfZyczUv14jhFCjqpP0hDOH
0+IADQWKrJLUzdKq/74KGwaH1zxyevcMulza1mo4TwQ6gElATN7/JluRXcmXrleb
AH37Zp9EBdExLVAIpPVRuPPjSh5samv51FgKn72nXtgEwACmuoa1JdZeUnexYRgy
lSdsu03crltF4nEVj0+ZxhMKLh5vcDWucnGlxlkQddqYiJ1qaIAunbGI4To9JlTT
ZhTAAY9OiPUYRn/xv2DViY9TBJAANBnY3SP5EMBwCkKobQ0DRi/90FBf/nxb938r
FXiUwsQbtB19u9uOL+bkep6u1lfHrgvKLErcTHIZ+P6VVnIY0UNsqiEFUnw+PnbW
O4X4NSgVZkB1FsCERV2e1I8UAPMtcFmGipFfb/rgFspfetblzwwYGzQGqP/CLMhX
zgsLZfs2T77iqUtcH0/VXdmYBABD18Nn+RDLj9i3GEGsZiqpjMIwCofLHcM+PzHb
9TlrCrY+R1+TqZvPnqjAW64I9GNIxuQoV4F22QiyvoaN4SSfskYWp+tK9LU73qZx
8Upd3tfnBpiTfLyxVEez28GmVxm9OBGBCkYaCqa9S3azmjxhXmaZvk4Pl8REN1o+
aAZ+nNP6IkE4wFhM2rld7LIN5f34ScNFldZF2KXJbLc/LnnCtxXiB6zX1CLW2yPQ
7Yz9wOEBqOAC3DDciZAdVNVjRV4YtyrbvU+1JBl29y6ETl/80ikbtbBy+odbVdwZ
lNzEC/jZRmkAb5xXSGFiLWXdy8HSdBYE/ou+k/dC7VvUDgXPmru0ALWIHp23VRby
Qj7tVcDzlQzxM6wS3wXOryMp180AcaLJPsB8AaY71bUJw2H057JMEqMp3zsndFBJ
5/J609FFnzENPwdU8BrmRy5JTx1Nb0qVtcrnPNvZOP2zJydzwHZMK0fZqSbKOjQf
5Trg2lRuWgFwVo2VZOeYNnh6Q+OwTBLQ4v7VXLcCeyjpXbAHX/jZA9Zj8mfNU5sn
h6MXLpD5lKh5laElJzr64CZeWGTXJrx5BgBM6yVgtDOVjvj3qBmmkXHtwkagb/0j
oGoVNWmB7AJljC2/nPQIkb/fB6mdLgBQEyURe7xZu6LP4ZfZGgStPc02cL5J9i29
TQIzKhKEPmWQT5UFygQBUbgty28WaJ2k9mMxpDZlQQQry1Dfu5iFugqqvzhiejV4
miMCCm6AIxsLhMP8/vOgIZeMVZsxChYIV2Hh2jomgvHpGMMUwr00g8/qjh3HoPIe
7ZNt/hTH7XlJ4sSgNuU1RSD2phgFj7fhIan1uuhWWIEmIztdpx8MJ4U12kiW1twh
21JbQ6d9uIBa1bqgp5M904dHkk52u5yUePhmGxdTIgeoTOmijH+/8B8UrJRvMeC8
jSjunKIsXiP1kFKpIHLlzICUkgt8XqS/DdSKcjg/PaUbSQtAz3cdxI22dlPskpQW
42LaQoE3Gc3OJZ4k4A4sHsKf9IlxilokVWoxtw6Ia8vLsgFzwC9+jPF+5T68huAD
PmoGuAj+g7JkHWiHiNbMHBLJOh89qjBqI+uj/xZ0zBhn+BIRly5GynfxR+O28SUw
/UeN+b+IUlHwlzog6hnu76Lkwny+2TErESMdnRNBv+V3lWIu0lzZn2pyqbRmEItU
qje/YluKINl4QVBx1kbEDtbNc48slWn4j2smg4b4L9ZqQ46sz05VXjbLn9GP8ZZB
yOOxoTVkAW90nnQ+nWmMtUGj1MLhIWsWCmPUuAdHcFfwbkATiosKPVVh1yJN76qm
jJJJf0HBtABK6Clqq9pDbENQ1Wu6lu3hlnrbv5rVzlAFiBSEIrgWpN1sR7AoDWd0
19NWHtBset9HiwHh/KxjrHij4QjQbB3UKVRyVVnicuhNqPqjAe09tiI7hGW6FUvx
tRa6kPvT/0WtVPRIyqfEDwIYCuqZetFdSShYFUPHt7Zpa952Wtny8a2abwPbjRVz
SQjzX8SB89fRx8Zr76l9RgZj9wnitysqFvLL0509I3iRC5g1gd7eh3aCxEHmZp1E
yVlcdcp1J8+EQRTNLXYmLhEydBOhYQ6nJ91NEpS1DaoNVd6yRZVH2t5DxEoi1fUm
7Lt0A6cvPuYB4jXkfVN+9l+HYp4XzfFjl8AGVrGDA1v+XtI0Td4SMszycT6N69SF
cj13muXaW8RYAo/HtQwPuQgW4v7ZbO42t7M5T8cplpt1+5TLLtUMHl6dD6estLhw
thIX47TSLLHHlBM7VnMVi/k8JojTdSRP3xVvpCmxgRMQXVhzYYnZDRG3oLQ9+HV9
cHRHdI2CZu/LKs7J8NnXIZyZW+aMAmE2FL+24IUGJgNm3rYbwnEpTixMv36BVF1X
WcrtDKHnrKAAWTxVnl0yCuxgFBIw95GnHAc44qxe1egO9A0Xi+aOkApjdP6re96H
hhzal+MRhdn8LkhA7P7KvRyDYGwrrjqQ0iobQwWMt2VdxlsUt4pT8hlmWPotAUmM
nS6uDrsuS+C3bc+RDaKJkrXNkFuJcJTMROALzLp92zbxi2rMT7fGDHJalh6SO6rH
zEAox7nOF1qh7VHDmlHd/e8LBMe20+0bQCi+qQg2afaWDDB7s+MtpjlbvxDe1zim
W5O1wkpTlbi1jUqdWKaI0MMxIHYMRpWe8Wm1ogmbNBRBBH2FW0If7vqaqfNx9HzO
YC1U8ZYAZb1SUAqcxwPFoPRzofbVj1lPOv/yecPeJZfNUKk5KyfPWo8ZhPasExJK
47/c6g1QeGmXm3gFeR3JjXaPEolhmrPIA0y3RQ5ego4t2svfJYJb6nyrjGIhK/JU
hsWPX/gWIIxeMz+MuwI3gkTFrbR8Au1IT29XKA8Q9+zpk26z9Rv0cg+8vMWWHk9i
kbtFaEn4T+spN81n5sOyDWLXPLGlegE07fcfO8AU61wKC1l/6Ys03SbVc1Gu1N+A
wnnBFd3noJ0qNLpmoNoAeZC1VDtAy+2JTA0dAZBog6Bbx0m0Sl3H0yb7ysx4mgTS
kUvkrurbFn2lrblCPH+dBawxphYNQ9IH9mdOmparQig4MljZ1pXk9SCthFQfRnXD
ihRk6ybgPcIViXdvBARpthqj521N7GM7lfzsFtJVD0FEGHVGkLpUXEInhW9TCvlF
+JKQ2bNaTMzvuYDTh03rmT5aBRNXCW+31+K3xxzaHU4XYU/0Hc4vhIICWknuJX7n
RNA9WZWN91BK46iymlil93Ys22oOzdFAQf48LmqMD8VJkmsdQfh+vKXOkWcfvmvp
C333NdSRDxZgqy1nwcpXixfBx+3oixjUFVj8oLdnSYQhHe3w9WPQxDf+doDKVypm
cipG1cRnWbDuRWrhGZUHItssafx5HjqNgia8bqwPoSW4QHSYmzOzWGQOCA83a7YA
5K8+nohFmzeBlVt+z3agO2rO5h/zKR/yMOTKoYKXq45o4vp0f6IGyVy/9zDU0MpS
dHjYG1CV9lGK9aGdFt5S0EvvLcuATu8NRfW4IoidFYaN9Z2NtidZ1eAv+uSCJxsC
RRqEqDuKIDYtANn+iRo7ujdza4uIHWmMuwn8NUnoQAMxCJlk0x+n+o0LziX5Eghz
ChpOexmKVhrC2Q5nB9o8Vqk2lW3DLLMetNXhL2DR3+93g5zhHP8HxGMdyB0iJX/p
75mHrvTwhOm4HShQHtwOGkQdfWVQXMNpqzCCiTHVgjtsEKrDZpEaoqS/HLeX6YFl
kygiVJX7EkrU2khd6oqe4mVBE212plKtpPvw+b4CRyaceN+trLZalt5gEGuM5jIN
7ruN+lrlXkSn1iBr66+st4qXxwHwc0k+2lcUwiVWJV3GVb37J64G3HozagpGe+uQ
VbTVdh2Qc6a1oOx8BcJMNma8k7X8ZI+TYezc2Qhcide9Z++/ecFQC04a5AYXPbZM
oHWs1Zftqp8K8iS3qgQypAoATdHIAvDdO+2J0Rso4VoryaPWozbQJW5D9QURi+JF
pRgR+K6AZC9D8NbxShIw76APHWyMCGCEyD35xfJgOAgiDm/Jyx2vRP86rVBCu7kG
4kDd66mx7jTxIZWOwsAtJcs2jbhf/2QPh0FO4HTDSziI9VIe2K9rbH3fUjqSBQN2
AY4rw6Qeo+jpUSYpoWSktofgH6U+9506yefDPTJXJGCvIE3XCYHbb+WCxUhEcUkx
QIq9PUSj734QAiKpAgfwusLDIOss6pLhhpAADbdJGM7u/c38agHjiEXaZk8/PHqw
Wd8TN8WtwcRM0llN0JE1h0mNV03ATYIQGWzlLqsH/BpKQt7/fmtEoTy2xQ5Lv6UE
KE4czmugp9JLJucX08Sixpp2AHCSv1n3jT2QCwQlt48QY23D8WjNHeX/4ZM7MmiC
6/qUW9JAwmIPewkPm/5slN9fnizWvsHu3HKgvylkauT0f/CmN/xvKn+tgHBhnc0W
lK2KnKAb2Hg5M2iOIEM4W5ke41gpq8+XgaZ1T5puOxjoldWsNhfjzE66S2PkICCC
0c7VRPmV8SOYsYbF7wug9pGJ5DPEftT5cpdR5INisL2JSpCGtUv4JELcBHMJlFs9
07U5KRXy+AoF4tO+YzHAVyWsZn4C/fHmlxK9TGpleVAbTcDyeH+deQ6EmZaZvlTQ
3ocDQu4HXMPzUswm+47xy6+8QbFaSLCKA1BzaXywCSkUq5LQgREQogyPibbxyzXr
FoY263u4JYMNKa8AgW6SE7JCzSCf+KlgB1zVTWFjyLsUi1jAOhOUvmNogSaakMqt
5IaYzuF1DNcDWOZwjkJQchCh9qXDUkdTofbCTNP/QMRd4m4HnXTLDEtIOIxNU1B2
AkAWk/tACEQ+zuCRus4ZtxR58lqT2fjL1SyLSfX3sTFWIoaFEvMXwOGoESBjPzVn
09+3pTu+O2oY0UQvL3vtd0LgSKtp7FskfUbWcMriWjv0MgQqVTROlPAQP3scWhao
lvdGC91crBWwrEKoFZfRlQCwUTgkMOFJTGZxhnXv4xAQDqajqhNVOF7LZZHMek7H
ZMLniXGBm1WhuCLSgxiL+cBZ2PovwkzR/j8W0iygEbDHO3XEmYPkZAMQsZ1CQeq3
N094T3HVmD4W87dldTZU3XV6JNVk4jYNxKqY/EwlyKP/OMxUjUUhEKSkanrc+ha9
zCn4STxB9GRVt75Zof+5dcf97OcQnwI6kSxwhsPz6X6jA117T5r0ukLFBIX4HADb
Iwcdw3qi5XVg4Wvy6ovo4IFab/xJQEESq0kaBlObv+H4x3CPffTgtmYPfJrxZfe0
nbgfmX68FsvcRLCMC8kWVqO8aTAxxmueivq9z+st1Z6mccGJg6g3szSGE1O1QAPH
oHJmk0Lgcwiyhr1gsfJTrFbqi8c8qa77SrAt5WDUmWLYfvl0OO6tP7sj1BEi7uTu
110so3GnIuhCG1ry+QEg6C4wejfRb5Fysb+OEDphrHJehC2LSZ/AKLJwdmx052yx
4gyzJsTR2jWzWy28JwfGwcPTqxedGEZXd22bP5rAX4dhdvbdEcUrisrXThND03DZ
OUJN8e6PmuE682q+8wVvdXuLpc9hpRKGtwtz9YovvaHYzzKmzLjdngsUou0o0tqZ
AhXIAfHXGiHa57RmfZqCIOscPSf8gpiJv2Mbq8hqXOv7/skV6+vigY8UZnKQ2npH
WeE8isF7+cV2xsD9r/5ppCZtbRpfA2Iw9msi6MccTDQ47Jw3bI7YWljPB0g9t4Ao
+rX3iDrvo//8DPLB8ZObJNBM46TXgESlFMClr2zlQPQBMWvqzEmhyHdeu1AQrqX1
fxqG6but2TW/U73+ITdsfwgaWkKv1VB+AAl11m+fLUR3uNtDmxAHwRgwz+zAVxG4
H9OhY0XY0aTjCPO7sUszrVPI4+hr334X5vJu/P5xkYb0EmPWM0zzwfavPqsVFP4q
J50Q4U98hK0Uh26lU7wJ4Ya52U8B5CF81XpVKxdI5ka7az9I2b4tWaATmjgWinDM
YrKxFmBIGJOCpjAqCd/CA9ABTqbok7XPs9QxecjSguZXXrefFXA3wCVunwoWKaNZ
6nAkMkr7sF8fXcckvr6A3rbW81GmefSJLL0WS/aL/bfBYbknFBtUppIqFguyDBZu
HpUE+BbDZzEWtsdSEt96hdYteExlRwPSzA5mvVWo0APpxZbMPvctjJbfgFnCL6IS
xuVTQXWKOguePhpac3NUKxxUxdLigbfeH26Zux/Dtad1pfEvm1VpGMbkaRVf2m+d
TNZl4WBsg9zwRZFQ9PR9Wxo6L1sF6vJq1qaNPjm2J12TDmeBTJI6PRyeQXEplNJd
MOAbGH+7cQx5Xec2Gn7V6+0ek6+lIzJDYlNPgX1TgGqAC94+lt6HDTTJqRS8pMFw
mtLViqg2/3YVvySZpgu6x8DpUfsi5kNhT3Ml92QEBVYYtjPxNFdRgedFe3Lg+Xz4
6a5JntH6jcb5JPvUaOxwAt0YJSXE0T3G/m13EiShUFISOKX7wKrrlLBMrzNA4uM8
+ypID4JGdOA1wqU9J3JIJqge3/XsOj080cq5A6zPvZinn1gbj8CJq8HAwCKL7785
r9zghZF4g1OgZBxg5/SCflw6WzNQlqYcN6ztuS663j5Nd44Ciks/4YzrWvNoxbuY
v4StUYWAHT6cplKhNQb8KgQ0UZZZS3fyKqwuNEBOsmqkp07Xq2gm0YrCMiTBjzl9
cYg9TM86dj+NdS5qB1K9pzY6JHS+8gquc8dOHsPRDQrvYZU7o9Rwa0Ig/Oy66PVD
arQdjx9e/luWfilc19FhtyId4mF7MiVSEwlEwYTtKS6hwpQKF+uO55z+wCupgiGV
AZ5GCTrnazrr3XuVDWFxsenSNTAFGiG0XXsdqIqesPmUuy1L5x6/k5ByuOqm/zI0
UtlIjZFO3CtD8NgPikooILJENS2iDXOKOCdHfVyR1l2aXTL6poAc7c9z+/MtSy5F
kcctCgF+FZM2BVPBWQXgAoImG5BwGMFKMGWfyJSlo4el5o1T22yM+WUqnyrEqr8v
Zy9cTdhj2EjCm/ByjtQNa0csBPSTl91FN96nOcFSDlR/9a10oExyRSmnpC3dc/qO
im/qvRSnLi9z87O8+jEnE8lego2P/7yXsTwhcNCJa+DhbQph5ljszJ6b0aOqZYh/
vTCjuY9TgqgJLYyhPVf+QoxEeory/Rj78EdQhbewTXSM5vpts4h1AXHblyg4m1Ta
sy2aT0xaM3K3do/Job4d37cUUl9h9QHB0u40YJ/CRO/qqbQZYa1p5gisczpiJPGC
6aGWAVBXD6wqG15zpEfAIBeR92WucrMcjJ+RJo3M6ueRkqvjL2eMkbgpGD5bMzQ4
bmwrhrSWbxekFkAZ+NB7mx+h88ePL1GZLthIJDTTUElMweYPL7YE2CF4zYPKOEec
pVhyVDb7b9OJMDFbeH2TNqIM/ZOQL8hqIFQTqwn0brBJW1LFk4Bu9ecEAXz4QwN2
Joj/W5UM9RUyz3kSh/E0qedgjbseI6x/AaYNZEFsPCVCHP7bOKugt+t+GZ7dmN21
/XMlXICc2UmTjFBuvSnU0kX9fy/C/H869eAnr9jUDyJcMN/cXkBBctG0Cn9Vfnl9
er8BqawkQqyi7BCGIrnHM5tvoBdDbZmUzqczGM9joWbSDvRwbxd+FSvnDPDtu8Eo
IwTHEpGz+ZemYSkWdNVCFg8i7p85qXnHyvSDC0TGJm13/dTEKvxgPvdmmvTT1mD7
bOidwysT87047RCP0PYdeI8m0G13ynJdNEwufDlFSyUQRZSVOfIKJmyPahIFLnUa
8qzdzn4A+dqLDPtaO0xNq2A0DBfUa04oYSSib5YY+jqnG0dF4KZDymlVszFtu1QV
8bOE4Kaw4qLRCWbuTHEy35zH6w4tU/JAdI9m3VxXxVjZhEvmMPYio3M+/tv0D53L
GHGKu57ZIU3z4bIa3LzHUf4g71w/J8sJWsO9k4THm6Gt8CLa5RdNoZc9ONK/ztJN
EvMvPj/iezbwuBiXtu/4icPhy4ExCfSqvCOOUjgZnazQ3rIi9oTxD5AfINKz8Pud
NbDsjlm98cFj3WUGDwMQPhmZxVjuG4hPC5jBAa0m4WS4d2HBZUDUD66ycMeDn2QS
SWRKgiYf6tCYLVoj2zRBAoSpV/6eRTLPCGQR9hQCN1BpKKIGXvWmqJRTDte8YzNk
t9eLURagE9nQSZQtqPaTtxmuOWweYHN5y3cU0pax+N++f8DAVpQMsev7iH6/JegS
EzyCmWDQ788aa/QYXZ7s0KZ/60CKIJ/Mi+JzqYf8K8IcbpHgj+s0/uXUHUPFsHmn
ctk5QW2Wm7xboVLMpjafBvsSI1UEX6x5+bHA9qORAVrrBQQ+Za0/nUSJh6k/WXKC
0EDu2lpm3i06NgGl3s7JzYOh+UzHDZWx/A9Dei86wSTimrXcDnmlCOnZvswC8xBy
OEs30a17MLf9j5vcQ/H8xKx4r7H2eh+invhBBcrKdohdKTcCPLFSc9EH0/2AfaY+
m62r3SC9MqvpFwU5XK332OHKp8o0pjGhlm+VcGU81rUcQAiXUJsWm0TWAi0uPt8x
76L3V/rsoFbgIsPIP5WfsrEC7wPe79MQcrHHi3DNRTkURJ6fEwHKEQEWOzswCiUO
JO+BCq91hnQ54gMss39LazM3pYKYajMicoLtPYRPi1QReQIYstFYwoqR+opaNioE
YmozvblGT7ciIr/OwmomqVCGvEHQezZR+GqRjqylzNU/mRQpmGNavK6XPVYWGim2
HREUPjS3byHPyhQxdrbxJnTy6ZCa+jX1ZY86FlFEyldLhLJyxuq4Q03VjgWd97IS
3+guXriSVLKvZo8mj/3wrqJDv8+tP2lKr0BH3lCgaZGsVPl4wD6+R5uu9Lc+EBHD
CHRhdtqQ5+m9dC7IKy18LaETWS4uLk5lqC9Zr9RHGHkaUEUG0Wok2W4nG4jquqpc
fWXCEzHwgR5q2AWLBxDYbE92ZKtJzkQ0jiUPr4QEFm/5uJ9ub22CgSfANur6CS5I
ymEFSvsXUVnAK+qY1XhWpZL+XPqlOs1rOrfxLe2FDe9Sy6uKihu9cLx3EhqXR8D3
V0+j8ZJfjR4dG0+esZ860ABfuG6Omf2nS+cykPAV+Ni4RSh+ptBAeHkcoHVfYu6i
WATsj6z2QtpXrSUkHTCM9IZ21EsHTf1Yr8bS9m9doiQLFNhNkIZJ5ZtXsZGYSJmG
4dO38/bPzNKbLBqgczxBkOJXZk3kJtdqj3CF+9bcScledsJCDNNEIzdGA/a+grA8
EFcE7eTwf8t1tg+cw3jR/RKgSHfo0LKMPVb102w6aV6WqNN5M+UuaykCdERDMImX
K1cBaLroYKv1VLRlQCjxQWrtORBR/eQjy/ahV9JFnyJZ0nYFfQ2hTEHf8QZWI35V
nWKNSqi8MFp3QfmHtOM96MtquKKbpQddTbWNmPryhWNcXUueNXBZ2ATdDstQCBWi
39W9HrLcK+dNLZqw/sQk+z0mTLdNNKFzegpttXY1LNU3e78WHpqIaXHWrcKNC26E
xr5XFk/GzVA+X+EK9NE38XkNP+XUi90Nl0Q8G+COqvzSqIXGqJoIvCVPuoxT7s0l
j40Kg24BE4HfCrtpBWiSpnkGyPvg36dxkdz4es7R96Xx+y0m9sqjdjUeNjsuzqCj
ZPP4PNfvx+mBzrAbrmQbMXPzMgtlDjGtXqajyR4LYACMaxH3dKiVibLCDmTM+sKS
R7K3BWZaX0oX73sk+aFb98hRSzLRuCbvxAAcO9f82ctkzqmB2YLR/1uXtdgMPOK+
FXQ5Xf1IjgGcGLyh6cQ/ZL7ZsdeFDvjCdud4yzyOgccnFI6nQ3aG5/Bych0tOV7J
TbHFV1y45nLvIy2FxlvoeqnO9HKMaKZWnDiaMI+ftK08JvLGczne9DKdFFmo83Xc
6OuGRNEgFzXNUiK3Hc2F2L7jgXz0D9MK4kGD2aUH21xRLxClBoykIxqkjuuKsIj8
Sjfcku06QSnqQ1mEX1ytnSCf/pFb3kEER9pvojstWk6Iv4qXHFjIbGITZstEKTcg
rUmrrvUo9JgWtRFFo8WmBk+faQI44c0nNKrGdUQrbTdBe+jYe57O3z70c4riAEf/
uiZzkVQXotuE97uEx2JJ6cWRPOmdZh9+JYTdWjVrCHn1RD1pueGjcrC0JGSYrz16
bdM2dktMgH5LJfDuOCjrSrUOunRF627SBsi1rXsNCtDox6fyumg1MJRsJPGWisIC
aCBSPeiz3+KCZS3TIvpGw7LQT0YkqHNiPqhPvtT42diJSfTmolz2DwbRg3TQGyz0
rnz5HT11cs1V3NXn7xro6MJzmbrL7SRojXa6NCSXUyHJ4Sizaanjcvt/8sZ99cP1
OE880nYkI0hFGQBUy/W6LhtP5UV0uXHKLIm1FO970/gJkBICwmCKOESeBtA8mh1h
FKSmnL+Smze/93npchwHWr2eXvIRAbxYREXxCREp1ztqECD51OVO2rhKJo6Q9SqL
07jCMWFjudrrhQVKEU0AMoVlgqYadwbP2Xc0E89+3EqclqhzUX2MJ+pJFw/+3H4G
ScJXHN6Zgax8uGKLu8TrxcvWtzFIcN5aX+fcxF11LANg9pjHroeeW928ogNaLxZC
+OeTD2lQN0p4IqPAS9RrPbgowmDQbxyqyeLCgKnh3zSaQaHZR4UkX0ZrJ4b2grSv
BFYrYsShSolaukfEm28nwOJyhopgnDkgfqtpChqVt9BCl+1q/7U7sQJMNJlzNZ4s
eLLESIFKjCFT0v5m7niLJPQhjlMIAc3ZhXAsaDIr9Mi0qNE1yLQLqyB/14h3tzot
qjgPV+KcKUu5YPglolAND204USMMNs9ssBh1MDL60rbJRwpxGgL35rTCWxB+vrNb
OOhaSDIGADgfL39csNBO/F0/xKi7tIl+z61hqmw7J5P6opS8Bpm+HG7ohD5qoRBg
08eGDUEugm0mmHwh4T2/YL3IyBeM4TDEzKicqxqgDb7YC+WavZVNZsgOow2qcRVy
KVhNDZidqQC3dyg9jY9IjjjQKLjuotQKjsS/5G7FVlGDyGyQfvWvjEo/i2M1+02i
L90A0kaqMKggzYHto8MSa9zTvqVRKbZtJhXR8BorAl7UThg5QoM5p/n22ugT1hcq
ZkSZ4PfVqLcHatUvXUpnYlwmmUXbQ3yW523ELN4X6myaVbLAFTYgf8jZLkVqR+pf
FZgvKoSOsHY/Fj5Q3IUMSb14iyCihqpQh4O4QyTBoxT9hLGYRqsVy8DoqUJc0KdF
Lr8v0CSpaSMnr9s/X7H3uqDgibc4kZsE4P85nRCC9wMSYDZkTmQYYzsp+2mCtE7I
fj28534b6fr2N3pbkrTvGhDvj5wd7cNbcT/LvxkAv4Apv1xBGPCSmeGG0JUPed4t
7f/ftLctTse7ReUpu3KLKSaE5vArfbQ7/ELqIRKze+JRYgnry0bpL1sn0nQjKxWB
Rvc74aXkDKYVqqg+EFrHjhxenh200MEwnrzWY0Q06CRgIifDvRQ007KHb0E45cEY
Sx5mAOOdXWmqb/w1wupSFhlQrjeC6JSJPn0PWez5v0wJ6NmZ1adr+ySXeGW2vZrS
kxuLiCpw8NtMAeEySmJbIPzk5QpZ+IelH248HhOSZb8yTEj235ZUtJ3Th7muPvZQ
jY/h8Zyr6yHAcrYJ+4UblA6libm8MkyOJCwrP9SMslgwML4EBeaX+8eM8Lee/ExM
maY75hMzJsrAnQXZ/EUwTV61nrv4j5lghsl3oKozZCgCr3C/F8WJp4nUZE+S6aU6
+CsN/UVW1WsvwnbHsGtU6RyfW8+BN2mV7e/3blFXSBNkboXRb9e1E1p1FbiQ6UlN
4Lhwfr0JycNt97fYEppss/XvmYF7JhHdJiST7h0yf3O5pX1jzRIau8CUnqGVaZqu
mf24uVWEO5Tgu040BxS3+PgsdN1FSCfqdMbTYQHyXyuWV2mHBr6ZdeG935g8XtHs
s30eQSJOD9SJJLdIUKw9INeX+sjQmGQrtWKrQZvEDrqZawJwtmz7U0U/pLIg41bl
pTfQLKVLVfIRG82LV+QRrR+UvY6H1ZzkqWOXLC9ExeKFh6hk4/lkGNM6YQuAlJYR
+ylV2ej22GxvjxrB23+26NOijSO6OtkHVShOmujdP3Un10FPJSAeshLy/3PBD4gP
UTEkJ+XMmvlrTTYaLCBdDfdDNejDS3tYGG1isedrILFqZkRPN9M4yLPus7j2C0lp
Xx5wEO94I3GnD6jeX7AhuMA0VeuAX3c0eUdElcXqL/0EqvoFnR2HOL04ii0MlnFs
l+fSYETqUYNgIjC2BIpdzLhCr7LImJ9JCRWCZkyxTrqCXE7zx0XOcb9uW5NA78t9
nHBgNwunwWrp1Vq+TnMdCWGhXeRlxdkZSeJI5tFf2DBkW0q0UgosziHsrtrUh/1s
wFtPObaOOr7zCzXQoWupWaCFODWW7rzETk6vLeoNowmDl/at7EhK6KwU6VP1QuC/
oF4WhGLSE7QNWXRZWIXxebpJ4jm4iME32bd3czRu+BzJn52Vra1QdD/he5b/vJbm
QFqu61Pcp4H0Fqu5u3Wehf4ZB2kbn1dJWprT4ZShtA2G8Tz5DhAGcyzKuVReJP9s
yBXYFgqCI/h60KJAKhAotXg1dlu8FMeR5TsBYG7o0/8Lv2lrvBcFwsO7vM2FFLkx
iCeUaP6L1WO9R6I1cvz7IbjSIThY1eCrfur4aP3BtQnmsGRfc7KNBfAHEUKat6mu
KNhQDC9vaWjqPj6VT4EkuQRzbYz97GqwP1KZxl7/PVB3wqioHtcK5sozU3OEFwms
gv5JZlvCfN9RsB2Hh3Qlq2KTVRMtC75H9Qqnk0NNWTGwiARCOr3Lsh95R9T79NLH
jPNgwU5KTAm7pYnupqIaQt6SQPCm5xEksUzF6TXGSVVc8DXjyOe2dxMFqYw+NC+M
sUFM7MN9NUdqNT9hdVlzLWZ5QaaCExXoszQsLhNcnsZMddr3XZrRfEcanfZ11jWy
EDz6kAJKbNRDUnwtZ2Iy9zuAvkKI36fPyKBB9QshmSXQp4Hj5hgs0z+gJiPnXsIJ
Ceion14OsyxlqqVMSFlHC+uMZDe6aFH2wAk7Jrkxhb5g8tcnJTZOcsWEVcXdFeUc
v1sN7autrkgMkU29gwPukwOS9VJPjd9um4G7CgMZdA5q/UOp4jIUWsftidy5Lgjh
tVZg7RH0z65Lf/mOE9ctOqHxsGlZVlfuBbBuw5yS3rlmyaw0VXYD24jGsZRh7EWj
ZaDVLEKOgqAuufr8d2omhN4n67JEYUgGoFcAZsBenK3fWhlYta1qYd4EDIizab0C
e1O4F/rwSkyXae3uhijVvoazdr1Pb9jTpMbFuMx3+6lgTVhMDdEZuYzDONjAgsuP
CN6qhF4TdjFigM6m5EEBkL4j9Zyy6zBr/86dJSclCleCtr5xUTh8sa5uSYDrhtGx
Up1hSowA6uLI7k7cc74JluHa3ADN821+qpuna+EpsLfnoyK7oWOVZAeNV2tMtCEM
pjLfzPRiZvn6cUptlMRqCj9WFM2hRwjix/d0XDA7tjv2u5iHNUPKSQ7/0hDA3fHq
gs2yb/OtwdEOVMIjMcYd5WPQvyEB9jhU6mRIiXrvYTf4cOILB+i7vYNFrYZrwWzY
1458At9faElN8GMn9FES1rLSshL7GITS8iubQlJsivZDbgJ+63aDSc2b3l6XcNWP
Jy9h3LTRPSagJpYhiQEDhWWd/luybX1yXIy7KdbXkXQiUNndKRK+mhqUGijmK2Ce
U4LMVAgeh03DoUTPBcK8JfbgM+/TnyD+Z822lTu0DdeNHgKu5AKZoPC61vv47bRv
9MvzH0fSYL8X9hnomUkQEk4Tq2Ly3dWNvsd8e/+qBPlgltFvkV71jjMcH9Ah4BTk
W1U9VOI6xNSDs0smJRXEXufVZ3gg+R/wpmCED2HbvfgG31SR0nZPGIzujd+IukGj
8boFFZQ0A5ktO+PEgjmouyMJKub9RtTJk73zjSIa+RomB6JMujggx1JNF/xZSTP1
IeeDITn7wKr7bRq+wCpogr4iU3rYKkgxSf+tOT8JdtIi3hSsNUyfEwkzMYisQeW1
MS6Ty6OPx3G2Ygj5ZGpBKQSi0vxosLp5thjuWqzDrwW+yVr8ajROcsbAB/iU/rOL
Mv4Z6WUKXrjQlw62mPIs05v1zoLqqk8TcwnLaR5srCj0gLBzMIYyLE2fzI7v8FoJ
zBwtfXup8CvfkKb+xKMpozwSUXFF2dIYGXVRrsmAAqi+O1AM9nuhEy4rljOl9GV3
FmmkpdIlnKFxZhTFNbGKonGPxeperodl2jtJcSFSFKz9F7bu8ZtIoPuXESimb7K4
Yhgp+F2MmcE5kfZ859l0ieiQmc54Kjn+XeGHyzPgfKf2zP25hFQHh0wDL90dLeCA
d1IXH+M0VSWNyR6Kah5Moz7EH45apZumgb/lAaczeySbVl84vrv9MY8XffsFFcR+
clJYHIpPdpSqIiryuMQ8y88WZVQ0d6jlshqdX9edZIlLwwBIMj+Ne0FXxWugO6Jp
6OmtLg9LxrQ5NASqBUTU+XNQVE40Z8b3q8/RBPTomfwrbchihkiCtYte0ol+FM+Z
bwZSeES6P/EyY2g3bzJDZ69iu1MC76pRAIFRo00YqiH5Guxi4cdJKJO3wPGvOKwz
49k3lgVwUkw4MohZADKV6l1CkPgZ8/cRkubD/wE9RvK1+CQMtgUaqt+4HGjgsSHB
0UZjHqQcrIytlsMSGyJPTH4YQ8/OVYCN7dkUE4ZhCwTwLcohkNYUVS2wBcj3ndNg
kaXNbMbpPokxCWSgnTT8Wcs7XhV3ElOuBSOWkVJsIt64uh6pIdqNKZq58vwLpbSs
RIoqgN65KKR5RucHxhPwTAC+hz63wLoFuaxeOLVedL+ls9mmMjHCmjMMdizSe75U
ZsQ8qaK/q27eWDBR3yGEFUyYL2exiTrCPCCQTRZeUT6HP2BzY2w0DwDDfXgZJhPU
DYMnTvnEQ+iiMuruyr1/+e45q5wWm4MzPQd95Ly/fZEaopjCpjGyeVVL2luZFZ6Q
gjd9yIAhK6ujVUWLbr1d+bMHlYY2TnWEaENRRCc07AqXbMt6mWcqgPAIppzl69RN
LNfGrQe2piS0XHgP65HQycb9eXTCRcwXktjzZYbAbBKoUUTExllqMsEXCfM9jMVl
6hjbYC0DgXKfEBIxYU5Y6vhF1OgNfMfnCM6OIAqM1JM+cw5n+FQzLDivp/8T5D2x
vngI7IgrjrA9VFK80wK9EP4qVellaEJ4fUnu2qKVN8eDbiYfrrwcQvpvixI71ofD
kxtrF1jB4jtIv4+iLShC7ACScQoQO8NuF+x9uMQI4mVYTLhyF1NINj8DNtavCyrg
i4mzwIYwQfR+BkLClud115LGlL7yjmjVVbzkfVftjFTzsmXQ/KfKuCGCEAXjAk4R
9H6+qJoFUBab7QzknKtG4ep4Jb0cQW8dwgjUoATRdiqNdkql6/SQowBETpZndRnX
Knp7CrKsgD0PEz+8nNvXrXtikjAdWEAhDTnCll/2GLBKOlMaPMjXFlXKO2Fn0uG9
pGIrzwQefr+46NhJncexKmmTG4fgrj6zPcWzEzM4NHT2ig1ZtrclFj7M60udgMeY
Ex+zMX+L0rMj1KQu2wTmTf15TPAf6JMGVwJGe4JBIBZTS3T92QttaIEwkrJW8onn
RMdtEYPCJkXzb8Jtp59MvR9KoKP4amF87bV4/4e078wCmpajrd89oRIZKT9AtzmL
FDaiu5zdf9QGmcgKAinngXG56v9+KD6Pvp/UzsZ38nZWnCffjn96laW811i049zg
QhmMLpnfwg+ISRF1XWHJbzCnR1mv9NvIHsZqbrsvlHGNRmUplh2RHN2pZGX7rpxj
Rt9zwbEGrgJwXP3mKIY18aNXyFhOUdyBYb2IMASQ7xQLaWtKncxruJw14jGbie0p
C5toNvMti70Y9y9Oxvb6ZTIEqm2+owUnkNMkpLFB3Q4NCBAVKV61hINLQhJB3yTI
0uwv3C8VTrJqA+tYwNlQYuMgG8RwhLme+cqcn1visUI7ARdbUe/B1t+2ZY36oW4U
6CT6CBuwtWS7QTFFb/XROAza1v1IhlU4ZSctdu3hPQRWLBECnlUnyF3nPgl5VCsF
+xEtyqtDsr1MB/frKHNcpoxolGcgxLG06yRad7+L/uhmenmPyWxltxuCDNkBW5PS
MuX6q6Vn5jKypuE5VDwqHv2F7EKdbkAA1qTe6X9aAfI2byaHqEc8SJF6wT2SUkbp
hTMBT/rFbPL1dGekBX5BVBCbrJ6CNOzY6rOdOyzIcOsV91kbVh8psy3cmiEX/RQH
DoXDIxgLL0/GOTH2pXicaCQmviAsVkTyAVwgyTaXuzgsH9XzOac8z5YBDjagKlWF
QDrhHPjHhPOuS635p0l6ZgHk0k5ZsWpK7zI3VY+c2Vk8bhZPsMji/Uaaub/0w9cq
sNIArozDzQQ7201fMTRcT5+IzBAIDas9gicYN9sL15ZyrxsHAEhOtwxipdJQ4mpt
nCvfRFlK0mWQcR2e8iM1Y6x9pdTJnThiHRUmq4aIpxf8Masbf/XL4ia+ZzGWo79V
wLWBByjzKUceVVlad881TOsItTsiJMZkzFc4KRGoYyWYoc3EwRv6I3FVZyo8QaHE
Rp2L5aqPwfXMoFXb+eNnpv54ElcOBK2ZQOrCR7kOtzljony4R8Upx7ZNi46QVeEB
HSVyyRZ5sxbgB5L38uG0cRDGe3PWXcPqjfD9v7PkdQ9vfNJWPfgLYXFiAQLFAVMX
j1cKfduorz+SXd7ynFNcA9ltNpFRfWlwSGFc5r12heeuf78Fgpe29hOkO/mU7u37
5UJqKc0sgfXBctw5brWDsaTs9BeKrkSKdKrrRVOaiMwGiN2kGZPElLM7yHWEpRK6
huodqkPHefsOGdHhIZ1101VMU9QwfEdPUb2YZIgNW+U2e0/ezGhgla5aMNEtTFw/
XHPquEYuqNuCJjU2ZEjx0n0ojhIIi+ShENn1qj/odO4mGAQVCOpILCchaQRNqfh8
Rx2gR8j2pIs+kEiLlmPgmkn6V3A8+zbCVqyKAv0blZ/tj9neG5tjp+QhXvnj3Ys1
+EnZohcI5SpoOTMGBwXIe14AHpmEayXwTofdFtL+6waFgjjmZgGBkh32aedmkn+j
wzRTtGj3S/0klzyDx6vrkreGp/0U+zLX35CTVsaUr9WVN5oNQmTctJIPWW4RjCSp
1HSgsIUSJ32KEj43Cd4IA1kDNRnnRdM6HpO6JyfeTOcIS7o02XdPe+DbspmwLNmr
bMBNn05PhbDO4UsaK/S90RFQznZyrZZuvgTyyBIHwpbMAS8344FKROnjBVvDlvf5
lFVfFJTj/CTvoddzQhpXtsf8VOJHTDtyJ0BHgzDZdXfkSUpvOQpMjN6s06FZCL4n
06SE7YJMFgRwrYuG52Xj/Sdea2rTjvIJWH6ESXcPduI056KoYrGyK9aLCv9DkZW9
RdeI56XUBbhAx80ao2MQfW3PZWW2GAJ2zW/2UooAl7VgyNDbxupdBmGtbUtzTsr3
j8X9HVkSOLecwEkG7sYKndnQALqKpCCWs4DGK07oIoBOL3k2tEQ8sA0TsSntPo1d
WboqqbJWMI0sgoZ/Z2ImDgkRz90F1zy0d7ZBzTju7u+hTGYb+U1sI6WK+CHN06MY
/IY5cf7HnP9SVXbyA3tDX69RKTA5diUyx0rN4PG/75bln4Axp2vbj8fvsuhEGLzw
Se4Ia+pACp6LaXA5+q+O9WIwhinkYfr2SF8c/3VwRUXt5Ye3X8JH8Ro1ET5YVl/H
XCEX+Pic4JieS7BcmF5IwywPSrcT4aOySUcQ1A6ig2H0qlR2yr8/0tsuWW2biA9B
Dt+prTUL1bGojqr/0l97qgJ4zkZI8kSgNlLnZALeSVsYNtXsDuQsu2sdLEeQhfLK
gZLxffTCqZzmV/EdmycNLZj1xsjgxhCcldV/mFZFW3YqbvmBEZ52NGkCV3JrIcyO
B4T2JjkcIizM+J3LiL2OdjmTYBBJmDSMI5JCKatkjvKcbq82ROQXPXxUDr0U9gk8
E3wHmo1uG6RDdc8dHx5s+m7xMjmmrL35rhdEkkoh90GPm/9kkU3uR6huc0djUM29
HcN8ii+HHtLIGM/kNoNi78XrqZ/XWQwMY19lL/p2LGfwXZiaGJLjojKqVILy7g9i
WCn1kxWUYIaItGzGw7iwa6KW4t2E6HBfaNXg9WKumR/Re6NgyN6ifXHrsYjwTckG
M0PFVLgNNzTicxC2ybXSZFxuO+lny36LuUCiZ1sy5Y8+6YypjLQhqpJcn8bR7wVt
FBd1s/aGMuKk7r/p18QynP991viZu2Mj4z2Fd0La3D7Nb2Tn6r2SIT+Fr71ndbkN
02jyw0u/5ZzYoVUjAOEzUZa5DHwpKU+Y8fBRwI5y3Zj+g6dUaddakYVbHbw653Tz
MO0WRUhnQiwCyCMnSl+2NnhlC/6GHmyFgHBXlWMMyLycpysKwQ3sFrQzfZgflkOW
lpUiM03N6SJMoT9TSmZrDwTIPXzV/brGHjT7Sc6yooCn6cNkHSqzfG/Av1roNLtr
W5pdmOc2QQV3TVU2ZMwiG5RkQd9JPI1WpNUxm8j6ijjXcnU1V8S+dAKpWzV7GhKQ
gTN1/1I3DmTsERFni1JeDwr3sgtBHTSS3aW86yYd9a1jwIdzJE9jBH6tZ3zr7gFm
VBtkQIBwl8Zz57ITLT4QQYUOGruvDZjBYaVB5rEL6nnq4b8Br/p+uFJIo5rYI6u5
TWtEr97761kf6Nffk5SGBuIxzI1zrLigbWub7/v5/m2jz09fn29ZXnsa+Ogkq7tw
1l2DZpSAgmD7iqpNSfcf/RsMAOpkGQYXOr45a/VpVxKsQh5UF+e3mPNMjb55IJC6
o0ZOk9jwp81FInwnORTqC9VF6Brm4BRVSJxIITRcPJPq5cKfM18dDa6mau9tv+/E
iQmsCe3OrrE/2jIA/vtu3s1ejSTS4b52FHWxraJMd/iE1W9WuSyV+hlBXvGk5Lxy
Uk5mB3l3H7t7v66r7PlKM86J8aTdBeBFmCEYkIDPthEhPex4XeIJw4+cnzqyWxeM
FHtukCIO/C3xtpC1IXvvO64BV6ZOGEgZm8xlchJZEZIPce2wqUgTm+AdVxR17OXx
BwxV2A254BKjP2KUDqNBmqyZvctJcTKfhCG7K09jluJltl2zUCAVaShXJTTDVKiV
m6UVwPUHyHMYPTC01uZi7GwfucbZmTMC8gOGcc6H8afjehmnNytXInvB9/li/a30
NYH+L1THeH50W7rugkxgZFOskZOORh555iTX7zNHjhJGYzuUBv4uAqV3UDTk2icH
Cq/WsPoi0E1qDz48mBclD7CCLQeytergeLTRKLdW6mkfEL1DynlZNCVN1R4x16UW
gsntwfO3G1lsc9yNW2SP2KdbIvOoN4Pu3OisOb1Ie1kmjY4MmU8xbYs/IPMuVLOW
Sauj8dHhoU3ONB8xgziLA46omujXs5OiDRGnLpOdYl4Bb7sAfUJ1qiaOn8HutNw8
0YJcOC3eLcNXHzYQuyK7CxXPXzMaxyA4GJ5BfrKITH6NSN7+CiqKzRQNOC96TONr
5OPGm7JWWFA+YPaxLb1BZwYFU3u6obkI/beNQuGbkKTVv80VxpH7eOA5YSWyePw8
sjGIMXIKN9tI91xqLQ+bjlLJqcbnx5ib2KVd6wa9UQg2PmhvT5v+kZB6sT58Vuu4
Bh/bLEkt6oz24utYzbs3nbNjYh3vHPlrbNyqS4juamxFiirBUSJCR1lcUQo/Aozb
al0dV4jQefXFBJF/NmQmsLCEEqo2wfdHnm4LA1xaf5EjVDinsb2TbN/ldtEzyv4A
hgr0TPTZqUIg9XNfM7koYE9CK8p4KEW56QWT5/rkC5dZLy3Cpu06N0xwQTCIVeHw
w0rRNxLWchw4FZYwYw+8BnEOTWIauhUwqNvMxqTJbJDe+hLJxRIG5pYdWnMqQOdP
xdyXiiDOBMUC7HthhqGWBMqbsRRvuf/ICTZyotxA7KvBAvSKHZ83XkMCR8I3x0mi
eqhVaRZ8pnR1dp704N/ahPJTUmn3JFNZfIOmj6CVeZgkJOoznnmmjChdeszMV0Qw
1Mu+ZFUb7Ilb1ZygoEokyb4gVTPMv03Vf7Fw8X04BLR+D4rbm9va1zXesRKuL+fK
/etYlbVFmKkYO8TlUxGniwcLhqfcSZQM1mbYT6eU7wACZFtdfNrU3zUcRL3TYe0b
KBFoV53djS4psiJXBwf710cNyKesnJb57FiNHdpyAXZ45zqUZYP3KHnNV4svvZo7
A++7m6gMCbXPbaeQRgI9EqvydBkBLQbgVVV/ezKQEdB3w3MQxKGWBZGAZNYMwaia
b0WgfZPDbZs7XspiSKSl/+SVsECLo1L6fDbpK5eAcKNbujDmYonDSQ8Uu0ha0eA5
G+5xkuL3JWo/ESY8xesbowPB2oNmf9VXBuNTqqcOiYg83aq73xK/MOgsaTrl/f0+
aoNdA9tXzfz2HRWYhMGFHjS5acVZD6KGExQcsIJHkj3khPtRkOnP9pVXmpKyST53
CF93sufk+IyoqZfCATgNHvhWMR7YAYgTdoF/EXvsSIqbM3cjX3c2pN7439C50can
aztM/M7C3BLf0JlKmKvkRrmGUbogy0dGx8bYlXjG5Qk+GPSeZgZ5W4Doa9LUuMfu
Dq4j2Vb97X6Xm22DPlDGu0NBFljb7Cxys0SW/OMn5tqZaM1nA9+2SCPUbRMEK2MV
0OMUZCbSbHLhSG7NcLS81bvPUAW+qg3UjDpXSXHdr9PmmfANL8n3W5MPGENkkenM
JYXiAVCyFzrFGCrvPTIghQssYKFCU1hsVuRS0i6I4CoxoTc8MlTHNmYw1wr51CZv
iG8EkaetSLcHb33rFxBwsyx1Ufei82SkSbSlmb+o7KgU8h4xY28AUc9TkDtGh4cp
RPgjZlbNq9D+SzS17gJ9RGGdKeddSms2DAnAfu39fxHN+HriVQFeJF5d5RxSR7tM
fLx/nbkPHAvnrYmzHSC6jfAJhcvdZpre0vJ6Mt0yVPqsqMYl2tFaKUQO2GTl0DL/
9JIv7QGh7p8j9kQZfldxHnPSkx0FFgkRtn5jIOQ5kyhJXY98pN9oCZnRAYKdOaaN
M4y697+Sv4PQqq3rmCiYtWsOPaR1A9T3RRWBlwZyPUsvt/Nyn00X7NhhYHlROeK7
95VkOIiAu1oLnsk25AbaWzBf7LkzxB1ah+cmA273UuKPf/ovJ4T+44hL8ow2yqLm
lVHZ3xBzfYP9lE8gfWCdiMlwHlnAVuujn1dpuRJX2AmeZX/U9svJNbPo9R/t5yn7
zfyT+NhVjXgEIOe7g8nn5EHtca8Df9L2Clk1Oxej7+ojoJPyxmsjdomxrr1wTWfA
5bO17d65hGSeA379ET3JxAO+NsdSE//MI1Sl+4tx5F6u0c6K2UVxiEq+/3PwGZqb
p0ES0xH0eb9XcSwMsKhbYU49HhWdxTbVFp+4Lm8edUGOJemWcoEbO2/S9m5gqhkp
t81TmZG2w48KmdT6kdWVKcwIe2fyOwXVLKgz/s9Rk4joK2JEIFyl1v5Btrm9pNU/
WJeqjQS887sdDLbx8tqr2TpIPgJu8GA1dhaBt1ijwBDbtBH6dpeazRXXhBF5e2Wn
JKQMppAk694gUzjezbPMxHzJIpgfUyDvOZUW5gNxAY2m8J2/GC7LDZaNqqn5ZD9R
q3hcgSiB4H1NZiGaJAAfksjNwvTY6iyaQWrIiaHstxRvMEPsp3+ZVkVFEJEom+66
NVJkZ3Qkm2tjjwfenqCe65WBO0eCMMtkY3w7RedL/sgZ60kK3YjuK0Huib3GIUCN
GOpzSjxhJ3D68lVY1HfOm1QxCS2zUFqgu5aeWbm7Arl7KY0DtRbcsSKsN2A5DN/d
AG13e7luoxjnqgRbgXzjCYQ4/yQ/yhd7VFekj3BrrCq34yMaXdYU1izp5PSzPShj
DlXrv11b7b4PpER7c5coqe5PtRlaoGkFSzg7WgzyaxB623e5UpHEosnPQSd8tPjx
1gSsR6+Q1WDOxBVz23C6n10PHc3rZRpLkWOi4KT1Uron+ZQwV5vmszSMdiwyN0pa
NyM4+JaSJmgPGR586S+469DZUJOA+N0MoqTjVajd8xxO7ilgVdwJbiSbdKhqcIdP
nD+rEm9spjcVaqFGhc/cJWEUS4DoDoT+s/HOK6v5SLDMa+tsLvzLT/OO+Z1eSGdT
2fthDNQUu/BM4u5iT6H043w6kOE3vyC6Zwbz2E7I6WHJ6y6y9VRgkGfvlc4bfHwF
DEAl3MEKiXpFPp2z2hsYZzOYMJlCGG6W0d0ByaXzcFiLeHYkSNibzYwQDX69FPXJ
K2H1qfEHIgMgzrdBs0170r5gdyW4B8A+y7JU0Wzya4fMI/rAlipxOBnzT+J0fUWE
OeRaxq1be/Re8z9jgPrdIX3Xz6fAsVSJMQYiFnKdqIi3wqN7Jwb8hJbUfkVadwVp
HfmjepjP+LPh/CYDOlB5D1t+8RK6cCBAymhCuTZQarpUBtUV703X6d5jrSYAuNHK
U0N+kG6OIbB4OSvmX8+W/IZFlPEtobJ5LdemYLLLSrIJQA+31fbcjQQxfbuyx6v8
lVCMBSFLsR6Emhh8pNKC4WYwMFTZmIe/zQ2Pq7LMBxidAjDP8HwPfIDpejebAaVv
0P5s371/UHX6/GScgVtX7JHmE/HOWF2Lu+Qxdj5XDiJnui0S5ndpR4mdVSZy/QXl
qYbRHrMHSkS18kV8vpXQgCd3FlyjtmlYobR2GEKaFnvfyW8ArBe8vluJRprA/iZY
Axu+lLmerqGjAvcjM9Cd49/pumIoRp+2d0WQPXOJ2hQBMZQATL3u8ADzJCqBZIOu
udW5hJddmjvVOZhseDVZPqgsvsKrSy2vHHcbyqm8d60lO+kV1v4e2WYoELfbUrve
rRd7SQaJfnG5CMlMZC2eGaYF6hZkjzvrSMvgaHyn/+jzG7LieNQb2odBrIAOoFEu
eyxVjNujtrX/8PcgyqYfvpE44swutAI3rAaC/M/Qwd9IYjM5tRCatwaGX7BZy2cF
2HdqagOZbqBV8Mu5B0ifOSD9TisX2tHC2uJLt8i4IwqT+1SmixD93yuzB5UhxPH9
v3TKrsnGWPry7hdPEzDvnv6ePqBK0MNlERPMmhbK/XtLdoKjSE7B4uEZzjypa/8u
nMHfhppu1V8PFxgrOueACtxHI7MFvmrCaunIQbjLVMbDTHA4VGUOp+9EvPsbhLZ8
TYD1CqnAHkSh3DNylZmCORkzZDTSfiyFgaA0s5vHNDxTdvmHeTBs6eg9RNdOlgc5
OqFb46/ZbKOPC37qL1zkFwCLPKWDCEsITJC4vkZxQn5u/K/YF2+uIs2MBJ9B6m2x
Zzi+stO88eFXzj7b/p+EKT6AVrxF9HxqKj52JbtB1WKNjB99Kzm5ZA693q1Ica4t
H+gyFByzy9SBgknjaV0BSxMRP105wXQ7DF3ScKfHPOSzAQpFzQ4rvWsXot05F7sr
PO7jDVYX/S6NYZYhyV2AxQgnq6SsGuOfSgZrFYNkdVhlfbFwlZq+vndeCigNF5wp
guQcDrijMELBcmGUZSim02Qz6V8Tt578IA5GQRyn9b7spDMIzohO7BHj3nvslwcw
h3zJdccQfI8tAOMTaPgmgQjtsJpNh4eWfTw6V1TO2+MbS1/ePecQVqFD2FJItSW+
l2lIaXHmdZL3cm6ZWFx2dAyys3dm81C4Yz2oujB+94+WWGcy97Fa3xUUjjS22FnH
rnyxhObINorjcwW/Pg9siQZu6KhFh4zpk8aIHzbcsMTPqe/lH1Z2J37fNGM3v+8r
qPP/Sd456D4ElLWQzdfUP8+wo56cbe3KcpBhnyWiEylCLSuGOzoAggfqGfX1bmOr
Ok1U2ylEJoAu89tkLaWineu5mFKSY3RWV56c4FfB/I5D+ymnerrzzzpIPIkH5M4l
KWZAcenfkAkInizrUS4BoolaocjTnLsZf91MgiGtGArq7UdBUy/l2eatqY4H+lXs
UfWLwkzA1s+wpdNSs0ubi1droPT8NUcEYIMOgXMx4VBjQf+CtZFphrLjAdxUNuVg
0jcHg/wVN6UaEnQ01ArH/uCmylzsYZTsK/ujht7tepmFBX+jEth8fAkeWv3Xzawu
E/d7Uz37X8jC81lIOzb8YNUPfE8hxfsprejxOXNJ7HiqEs8aluurBm8BH0nmKuFM
CKbbiRypnPgLNyeLq+Bpd9Pmc1QqbZgj4Q9HFJgqxGVwBc/8LF/jRLkpEnefB+mu
V9uXjkciajZzj/WH1bB9s3hiBGOHkskauJrJVd3Hj+MdmfcOSp8AQA7GdwdyGhmL
4nA9pD8bG7AvVCXC9wq3mbIRcZ2zx/iGFbU1hXAxusUl1WCQiTJoUudcrDNuKkLt
dNy+k30Ja3mu3iXAtiQgXQ9xVWOzBrfMaUjAfdb2H6Jsa6Y0W3nL8unV/kDWqqfc
LgoV4PMU0J+2HLI3guMkc6h+LqRcYwQ+EbaDGavWzFJiJ14G4ZZHEfZ9VrHHomht
etZHDnnSfS5AZTieQoqmQX1xCHX2BXmy8LbUK0E8kFM23JwGVOU3TUlHf+mS7iqn
3dDUcOQNU1Ro/Y4122FGFuRSbUtAnd1rR0gDvJryT7hPgKnsXHfISsWUE6+91Eq7
WSFRID7xa2LnHYp/y9DCpK24qohyqi8oLUlC61Us/ru0iqu/j4rvnVZ8KfKz7t8c
e+nwggY1jF1PZ7diygLrD6mlSejSUVKCYA5nza+0affdKXVoqIMqHOEnLLlYrlVK
cL7pStNEXlXiiF2g9aRw2QRFcOoxNV4YGdl88VPkMf7RELCUvRJ3U1hKOy5VAFza
szGccTQ+RZAwP9/dmRRtjXW1CdXlEWGI1h3jVLghUzpCleGu0h6hi/5wvEYuA/3m
cAbEme9HGmlDxeyynCK2o0G+BqflTRnjA4JfnXOHWHP7olJH/J1JND5+8in0PQ48
7a+jn4EBFrc5Dt8oNiv9hWYmApPh4O9mIW7LBPQqxFBpCXlocyWoOT5VWZsJHzea
HZCnFqm+xq8uyywdL+Gltv4p57yh08UKBQSPqR8A8KCZNXzIvLVmu2jrcjISoyEF
df3dE/FWuWBG4EiY576NuLM0rDc3ks3mmDVxLb2y7I+mtmoZjPDZYVtGecfDIhzs
92NB6QWPqoakwDz2CfSpumlTMtzurYNp6+H7OuxL+KbXomMfc0EVZWJyUuJnGWS7
5LLcd+BTlmipuol4rWTdWKPNCP6NdUJH5aROP69XvmhYr7rKJAW5saL5WQEZ72/T
9Xn28hRCO4v6Af/LSEJCowDqPc66QbUHmvekbvz8t6Z9QnlJjEAlhyAlszrlGK+B
m4A6pr8iq9KWSwlbdoDN3leyU98pCAtpEt39YfRAJA1cNZ6Lzd7L0qK/LckH6UEA
GFpuCU/SlfpfvbaR5Hdls2P5Qz85dsJOYBDB7OpysAFvzTXsxXS5j0fqDSW9zHv+
8NXKxFMJAC/DzTcWfoOSnd4j+nV6K2Wxch89IENzK1No9CY8E1SmZVi35aEwddP8
wJjUPh64iSHSfGJ2S4D564iPZnB86zjbqXJAMHOm9Zqa8ej0shn5qI5unt5pzpLx
whSXNOpjXcTouY7M9x+VhJJTK0mR0M9FxSvpXs0GUgvYrYEy3Dak3sDhEbjW9HXh
6JSvx/RclkKh7Civwdarp639AnyNzkZxkdRBqllsKG86iZWVSrcABSYSUWBU6ZRw
7Ns5QKnU1auX84h8eXy1syHKC9SYGM32nv5hrgna6Cn+p9DMxUqj+0DagvmBoPAV
W+h8GNK9WzohdPtU7IhVrXG1FVGF3400V2d1bfDK/zQF64Y82ThByRDnMWqTMRG6
g9j9vqB3a82dTkBdY3uc6E1JVOl7NWMQ3xgMGcaXJl9JX9ED0gnOpQHwTfRMfrvp
rnf70CQWMwnoUU8UKwOxdARKiwUXJMM3GbWMzaDga+SapI981yUOtYl2pyNUQ6V5
nPqhIhXRpF1ROhPhnzcShjmE56atDdUcBzSmlpXqBTNGMn9rncplxKumCj3PFCmZ
/uyYejxzktd7PR5AdykxCUaUjKX9BgR0tjIxGkfQBrCoHk64w8Jf2Ywcq9QwxsZa
cdsZVe/Aon+Z1neUUcWGKeM0wOv5yQjhSD76n2PALJpsrlGq3qH/Blm9sSZ9zr6Q
0bkngs7dgCiLNzx8wHLTLyJnKW+szX4yPPkV20q9qPsfTg76nrbc+0v2JukTYShJ
8hP8SLt1hHXI5LPawH84MypiWuKHT1SksKOtjABPaLiWpOCKScbl72M85BHwcEAi
z4oD5iWe+IddKb58B2/ba5H+3DzRJ3i/qdJbz10uOig5jFbvqpMwhWz4GNDSdvLT
D2Jd+9K93gyI0X8OPsQJvWwN0k7/rifOhRbtH86Sv+5yW70CmbYxzGJaIevIBBAb
Tu73vwIgK1WjGMComgydw9Mazyqybr4SkTxfGf3n0lsKqCQkWOjH4pi8LUN2ZmNb
IIkHAOLcpYzhXYxmwnh4EAwyhe2iQLSKZV9hQ2fcMu3i3SUlFkOSP+gdHlVc2HTg
HPQoV6kwoi0OwV39t5cKLDlBqfiTntb2EroSvbN6cW11nGyE7wMvS6Njh4HPgEOp
ZUbsS+9V8KMxZkkqmQyGM1enpNvv1RtI6Xhneupx+QideGH2Wk+SBMPKnQkaQnSR
+xEADlaGAr0B3tFHVOZ9LzFf/bqaYYsyjjkJ93rfOWugw9uLwZ5/yYTfqUsJfEkx
a8J7imz8gN7hfLi8aTkKRQ76VUVXOFvb3Mmzjh/9vzprPkaEbM3aDeUhPFpa5QNk
jpTPRGQpJuc/qbVom5+ws2wC9BP8bpwrsu4oYXipfeaE+zThPjbhtW7gnYCBcmd0
ZEzWPj9Qy9i8Vgkp4/bjMmfo6ZnqKsBBSyeEwaZ9EjcXooNfyES/BzGDdYLt3nZ1
cedY5oWlHYIE+asx0n956woq/RlHAeiRmzdl1/s7NM2jEaJogWOlcJxn6FQX4Cyg
A/p7SlULEga5Y7ng9v8i5MxkphGYIn9gWKePeHN/bPuYOAID40jD7A1hyAASIfBy
ZVMIyWXti/+QB3Iy5vjEAl+RAla3cfyD9Jij5JEOHHnM28Gryf922Z8H4cGsnozJ
4x+bSyADhzZNO6vmL8LTvh5eURzhaBqwExM6/OKQbfrLHbUiE0QqVTovO+YWEu3n
iYAFcsz+fPGqmtd/JPMlgfw34beFvv5bn54/hPwOSn8YmZCee8UpGaLtIcF0ipEz
umuN8/57IbjNBecStsKC9f1lW4fiNAOlt4g8/v9SEhpcb55O6ba3TJpw0Ch6AGrR
JnN4CET+xOEMmnTDNYkX5CvVIvDD3ihbB60XjspG/xp6uct2bTmrn5D/9fcy4oWj
EeRrd9MvBOGqyzt1iXSlT5xDvgBaEr6qdGZKthP46GGbK3UCcEHQUO89Tj3Ks3Jf
AMkrpTi885/JgFUXTC7E5r0T5M4BIfzBoR/0ggDXAsmOLBErryOF1VlucXnxh6P7
BmAAPaIEjHs9Is0XtfSahU57U23c9Nd2c+DZvcH39OWxNvrjPu/zRb0YEMNwo2nr
Wyx0PK4GDnj09yBt4BoJMrxfGXblhn/LQTQfwd+TzpTkFFyad1CHa7qUpxMzBmOS
yiRZdVEEWkx6j3DBfhkQDc8j8mtXfG2yQelcG6k/yxfyd/ol1177T6xbZcjstU+S
27D0fmuwzWtd5+1V30TtQ6FhtLZE2JCldcOKiQggtHW/H+LsolbJ1nTINUuauZuM
x8zJ82SZtXUCPCTNc3C1ZCIv74kAcghQ7y/NFabuGS4duHr4/IBkL7DtVTR9kual
2IFyijfwMA38YxgZHF/+E36OxFODElU7XzdFPB4OtIWla1igkV6WXiQIRjGez20f
hkQEB2EnbMoS5gTJ4Oc4uI8iRB7+oYkWjmUDj6nCNjv4jx9sr1aqNub/dKKyf+9a
wWOBnx/kWT5NK5d8uQvQcsFQXyroOb6ZJEATndWHmXezqS6DgOitd87Mi2gs0ARL
QT3rOZalQtYguMd2jhAIvlkGCAy2mGxKfxmMnY7ZEVoRvMES2ZAZn1WXl+986CF2
FI8n/GKfuH+NDnYuyXeLJvhbTORRQC5qkK/uMqfICMO/IPzsOuiJMytF8yaLmkOg
BcrHYO5fIFhiKphn1iACf/qAyv8eh9eQatn80/PM4BB0FWb/I3m4mPkC0Mjfz+9/
COG7OCcnu07rjdEt3Q53UE+OPvSUQJF8ACypBzrF8uNsKazZ3Crl1pr8VG2Xqnrm
GLfUb0u90INRSJlGx4QiK7zCSoi1+QWUX8bGBIC4/h2uVszZIJ6Lb0DxjGQSy85g
+UywfPlcmUlKaupVX7vxLXT90SZnwezJEaCq2zs0arP4SQl+t8oMB+u4HF4tWyF8
moS69lzfaiBM7UX0xM1+sWgbrez84J5FWvWibngBrZAZZdxWBn64U1jrVRlEVla7
S9rEVc+dII3jzoNnw6AqXcdT9/MWi91WcvgGhwPG4ZBoZ6+t632fbL7tKst7BiT4
py8nrOjxGXn4y+EMsZax7x2p8jKTigIZGNgiAXwDkRjKdfnn34sT2VwHra/3AUdT
yN6AaeslE/z8m789mMp7UCDPNz3V7I5beMlkxwCE8UDOxBpcQJ+sXtN7okF3+PBT
I1zDqIhxu3NfoqEbhH49jpL4lOXagxlSnt8PNeENsGXQx4vf1os/1u400XLgAHr5
xysIGWrhunm4oJq1z3QIItI5B0qoKCjuDxKCJC70oClkWG5u/TZ27mfhkKYrBhCZ
TdZjDwHoVkRRBmHTrxSBlrGh+lk31jsANFW2ko06sQ+5nj3XNHoXpQoaV1HgJIUp
IYHVd0D87Shlgce2nR9Ass+EJBqGaABxrpmuIJdhZNfNqyUI6DGnQpj7EyxcJdnl
JqKY6d8DtbGOmO82fgI5GFA83UanpXH5OOi1CaP/YE+HJE7ZGINIU1R6oYLJpZuU
8jiU8bLzpdRkxtiG3gCQ5PUvSEP4PG8FcSzIF3TYxuAC584oC4S2Wph/VvcWeivN
eS7voQcuxS+oSRTJIcGRaS3zQokURfFgD/lFpY1D8VLrOwXp+QZc6H6bi4KJcryY
o9hwHf+q6GaEb/FvDMUgT48qPedhpHsM2/oGronkqx53s11YI2PLJcGU+qJfVLZt
1vXZ2vtwORAxIqB2GtqLzTYOfUBgjkyXHgaZJtc8vkLNMXjF4/xObNImWyx/Nasu
Q61X8RL9P0XOFBV6+mM9TTCFhWlY54BgkeYBx9fW45aUjne7Gx8aDMCG4x57KUyu
CteFchsMxu6vLNUUwRTUdmqQ/6YBtfEXNYMcwN6LutOyu0h3bpPG6xP+td6beU0M
awBfh5Cnu+sNo7P+0MuXR77Ye0lQ23oCFZ1gF+mMvw7q2g9BH1b0Fnx47AhIX4h3
ukwtBPq41SonMHbcpDzAI1k8D3Tlgc0KXTZGm+/pE1tWZNjRbvpexycy70fhdhTI
LS49JI6qDLh08apqyyJBk1GoycNj6F+r68AKJSs7XTZpVtNTY92WoJjeEyoGarWN
1buxu8fnGggbCfOLk5yRBkaui2Nc6W7ekRzX3CIlJEaOnyb3wUcqTgkzRpTYa5mf
d50g7MpbpKbpYATmdrFQlxcJXcbI/7II185nd+eO5Vkv588JQNgaPxbNzJ6T9hCG
O/vt4gBA1vFw+jMC8y8ZdIMVhg6vg8xRVplKfjF8ESNnSiJZEp1ccivS8eTAHhwT
VDVe/F3O7lkagb4TSXyT9ovk9E9Ek+Q2H6vq9TkiFcBxuD+K/Xm5GCWc6yu9SMzC
Ulur9PZa+oVR4Y+G0ou3nodzvrxc3bWbK9i2xoTFcHlGhQy5KimHFrWosacXVreI
y1D+utZgg6DH6OPOL3OPlORBSp6bPchrN7qyg2oMxYS5q1pqn0JUBBc/wszEt+VC
SM7x3l6KvOl6qlV5MsUCQpPDvvxvErfgpNczjD43I1dVQbYnlkHMd5nSV4WIrEjg
AQu3n3ZQZ8Gz0qPkDNO1fvxqeyS0vYPEHyPKPkGPWVLcFtph7A2J76QsOg9+lQi4
UfqIBIVCudl6pd7Vhhu/GpjgwnVz5jz8dhAEHugFh+utL90qn5cHxo0qbO4pn0EW
mXpfKx2WNWAl7u0bKxsyyZDjLCMgTtnjw4Gjtcju4/tsLcYMtcvcRzZMF6rOJG3i
9mi/UGLtnV53r7VkhcS2PxsgHoItDNW60H2o/04f3xr4DkZnkzHux6+Q1mDeRCQ+
z8SgByq4GvIQZZxYX9N03puoCBKoTco8kRT0xJ+h/ODZeANS+N/J+QGOuM2pqn6p
N2DnT0mPDiM6I01rkkh4ttqvyHCnR1HasYshNsVRQlwGb2uo3yhtUC5VgSTTug66
4H9DEluqjewEk7wnZKFt26Mz8RN23jr2JOxyWlqpiOzDA4wBePpcR1h/gd6W6RcL
lUltnTWVi1/kINBH6pXUCjGIH5fPfASOO5E88r3veo87WkwclT2WbVEXYeJhekOX
fUN3NgjWSbDwQglhBR3pOtgz9+/adVmNhGVE5H74h5nzfsp4cXWskSqOttXA3uER
rnugFJ4cFSxt4KAsdnE3D07cYO2uI+VphdE1q95ezf4LQJWglQqZgg/WqH+9m4Zr
eI97+WU+CJjwPy+wRAibzqiof8R7SN3t9JEJtzXgHyGr7GfExlMXqIa868iYsgPQ
J08CFHSiRrGQRu2Shjh+hYUETr0JXMYmp7Tz9Iw/CQQo6JvhkOfIwc9i5m9JmTIy
/oKnCi5Su3KH2CUj62lPt19IbgmePhhGGVakoq11EKyuQd2l8sD+G97fR8h0ILxB
QlOY960KmJKg9sPGbgUcjWyuuBiQszoQfzx9Am4sjSRHuqyEfR9MpZA1OnctWzoY
MjkR47/sd3bsnjh22zg9IoJ5I4KIgfbD9z474pMkFkV6SbwzTPA/ZWIFUf7KRvmO
uH0qQDska+Bm3OJ0+0K47gjdcGV6bz6HeK+ucCAezPtgxMyOVK76n9GOAh163h+P
tIHAZU0I2uK21AKw9qicnnJqhiqxjI808lptqR++ByYBQ1E4s9qMMVCFSf1czxYF
rG2377mgVAgcPG6om4HDyNWAzralEVfMnp9UmGpvkfSNhTFXSPwQrMsqxXk6dFvc
ny2Rd4TEkqCatZ4soL+R78AMjdwWrY9tZf+YLM7QgCkCPXjAR2c3rWZ0ZKqPBt8/
Lwp5yZIDXb4cVSgMc8j3DgTZIJMVSH/52+Hq8ReqaFs+t+cT+AUr+PMycgH3GB4E
4UpKtzERsXWNgob3/pvbN14uPE5G5cGUVa9rxyFJuMhgMHh/3vdX8SJo+Nzt+ON6
uPLqjPWbSQYBnoswanDqhboT2OypUcXhKE0s9IvkrrPh3LlOCAp/A7hQRlfChrUC
IG/JmJcnIVViro2RBZ/hZTzQACPPHihXbiWw6gaOaE/5kothTQiAYNsW+4jg2w5/
MyuqD7J2kzfOY1UuVJbppidY+8GaDRtc7j6GtoMCBaELqHzxbNJzinhR6jrdoeTC
mSU+cArKuUUngMhNc4T6dTDC2KMVMkM17dx+bilkXNbCdT3CwEh+zbEX6wG4UFem
+BiP+O0adUppDHZglUOOJExZdN848RW1p0tT7r7Ln2WQqSGSyZHdnFgSW3Ui+XqY
VYPg03l1aStvmTUMQ7VuTf9slVvh3zGhY9N1a2F6BB8Z2qdsa7hkbonuWrao8GUA
+dtNl7/j616b+RCHWhh9ZOTFgFUk7l9PiDdwBzgCtSLxpgULZBAe6Dcc85g6v7Vm
nKPxpTP9o8YL3hURVPXV3E6QwFRk55p2Q8xSSf/ZV3oPt76K7r+xJPvMHu+0AGJs
eFlNRxxx4fVLM89joBhc3HyRXlsw4+7ANfZGZ5/EKm91G4Ta5AI1RCV55V4uAC2Y
VNhEwhkUeI9ZZlEM/mTW1oGrZyfJBpR/kfQpfoM2MTG7SjEzkzAbJSs0Z82NbFrA
YvxG3HoJwr97RJTok/CLCShlEJBgJPFW5gaw4B0763aItgHgx/fXG+gbn+QocYau
WSkBEWz7v4kRP4y1xuDd4ISIfo38o7YPn55RyUIRmz2OC24P0lHPHpNz+pAadIed
xjy9Ago9NmpCdFFFBKmprF9NuHnWQqf7778j7c6onfB4AJAShx2hpI4O1ikbbybE
QA3iaUicbJLLJ0jXkHeioe/FyO/w6Guk2B7V8ndD9f38KgCugry9H+leiEzmewaR
OOMdQeH++w9vayOwyhED+Iwp5a2LvkUR8yam3UZtM+OMzBPA8e9BiYsnmmY0yOxS
/9skBv9xsoPRA8zI6By9FTIFzCH/D+gwhBjNRb4k7PprmeKQ3aysT3y1Qs+WfSmH
CxBvATNKQSWdU/UxtkjaKd2JodxaTr9PtSwImoO+b7JHN9kl1QKMYcr+sQhwwdPk
qxsNP6sOLG+ZQuDh7ni2lCvlZ4qgUUBakV4lVnuoylDPt0tY5NOrpNQJW4O5kFRF
aiDG0LGf6lLp8cg06+hdJv6q6Acr29bZOKuJiaRtN8WtPLoVmPJ7FP9ZlHJfPAKo
a9PUehVG9L1wcIxV0Kfq9GuXvBT9V/YaV3JHbB+2o4Hw2o81sV5ULhyV7JEdZKhM
IW0I72ml+vCQgoa/7uSX1SWDvoHClqBSRbSX5Owkh6fLzN6e4ojBQ8uMPJbvtQ3g
fd8QZ/l3ao42HK3a5kua/M0j50TLvoGQrbFlBbueJHLnKW5dcn+zhKZMRQFG4UMF
RiF0Ie0l3Pmo8OuTLGqmSnQBhOun+9i2PK8VuCgBJ8nukGHwjXeqqmDH0qd6p7U3
QGnhDH26fi3DyKn4CEq0RMvzDK4hFRn8zascIa1L71gnWZoSyRWBKa2+1XM3GheH
xzCsnEwf22EKwM80uXjnoqQSQrnq6DvgCT/6TB8TOIAFWczTRpKJ26BUujTSMOxp
JkWSPVecf1jOL+m0VO8gy6lfw4t5GvETWY+FxOKex4tb8ko3iYukM9vLJ8HXaJnc
67EuZVnWqAaB84LN8Pc1WTBwEXcMdwBQwiHdtrCH7scxEa4yck3w4UpODosagbVj
RRRMj0uhK8Yv6hbA8lZTguzWSSrer3KckhKqmo6pICt5C6pX92XkI8Kg3yYrFqLT
SKwFrWZl95HwsxQ5YdCWqzlG8qZ+/nJ0R+mwZj7DmbVDBrt8qrZhf3mDuj4Y4aEX
rhMxfVoNNqfgYc0hD5zS1mVqLP6lwsHNIuiM2irsZcSmnEN57BwK3i5aRqggGuoc
KpDkjMr9s8o1T8WOhn2lPJydd0QL636VlVqch3zvWGbo0m5kGh+e6UKIOxWntV6r
jmd74W8KH2CtLCwufSAEvk01TarstjQ6uocLtEsyPu35ePgR1q4ZhTXfboj0jRyR
jJEY6Mp2hHyAfyVwPnfMfepeKyeZ2GQd3w072HRuRHvjogaWTge27EeNc2XBqfFU
0no5DAPPCDiT3O0Ks+XzgfpXkLU3l8aoWJKy9wMuNV5QotQjuDk8Ijq5bXjabfso
vrSm0fFVcJ25rYcaiaS2l1io9F7lLF2BGRHsxR8FXV2GaMkG99jjHNLO5IBy+LGy
oHXmZOTdad+oM/hHvrM86+c3JZIFIi1X+jf9rR5gNMoJy5E5sgIP4UC59W6bKeF5
hNmpXPOSU91w/7d0EesISUbjVbmd6AWwz0WuSM13fmVWXgJ03h6e7C/Oc/S/UGok
7tby3HYZnjCIWgiiyofjDnskHpGjm3LO//rgeOb0X65bMJfLx/BIGN/l5WYBaJLg
9zGFpW1gAtL3S/ZcD4G4fSpIdhc61DPEnZzCQwZePnfKQ+IabEiaDweaC3w889cn
FeGyQHoaVEMkdPalAzzVJnJcOUROqNLov2Y/CZw2Xf6+DkUEdjfoMmTMsYNwThS+
xQ7JjfbHd+yvopw0mWT2dGFwCbVE+PNdkmybg9LAlPuQEFL2yvI+OWjY0IQpEnZm
JQkvg7/f8kCuAbXy+5QWL++bgqWYlaPlhtCfLXouACUumH8VhJFiky1Tv6RNCUBd
pns5lzwalFKy/QSNTy/ADuvdTiQ5PG5tHWMMdVEATEqQZdbg/qJq2R7wPcF58FNI
Omp9Jl7Q2NizWHIEYmoGZWr+D4NFcivgbhUrWPhMAjtJjzjzptee3jEqjfY1wjk3
YajVO+eMg2iLajIe5iNrTxfi5p18gh4s1PMVyRw5AH6n/CzzT5pZ7SIGCguNcIM2
sfdEXY4dsMD7xb7YVyJxgR6uHvGS5zQ+1AvqeRVJ2WwOZV6WPzR4dQFsEv/JIcpk
4+jEdHWojKl3H1AMVw+OEAs+9umG6oVuYGfezr4XfciXT/xtcmj5EXQNiod+PT47
0G7JLfkTOv7YMVr7G3kCoPw+rwxNwFLxJWliCCug0RlieiWWbmziPo6dFmTIHVqT
iE0jtgyc4VDheR2u0fbANKpra+BW9SICq7JuSeu16IFQPH/T9TCQnwIV+ovRd3nb
GXm0I/+Q8fZY14SnzppVSN6aW2fvEOCEO528jBdY8fNWRljrzfqUMyLjjJFQHndl
88JhJOyG1M39C7EaQhe4lnxGZJe+CLZzCSajmtmrWDRXBRM/P9W2VbwghGS3AZ5I
Y/tp0HvexhAt9qyazRlbA3lYYGAdkNoQrPcbWqnI/fwm3auOtGw0lM38m8AwFb33
qspU205VCeN19WtshB2ZPBOBY63P84t2/tPMJVAsymWtgRT2+s4PL+EQLjHNoNBG
p6puw4WgOruT820FKgddZPDNy568aYc7Ir3htlSgXEC/8i50JCGYzLQyReMVLApm
iTewCHJ24QcuEgSDnlrzvnUVcy4nhXw4Rsz2dNFpgT107cAWBvuRwQ+frNX28+Mm
Uq+zm4zGa28Qici/rGUoHTxyFSW84Djiqsjg34vlPEpX1iq6yfYhEIE+AT5KW7ku
0Gv/B4WIroEE+6goEBTQd8iNtvpFL8iKrsrAYszHBJBD/dd8bXcLaycxfCLsKMb+
JCNbZstcDmmN1JeNgD6iLCIIj3g9rzvGb392zgcJ/JYXSITyiTigqa01+PibRTl4
GdiHbF5w1VdUH/SPNxZ8aOcsCXs8Wh6mNkdRVKwTgYSCPTGYQpRTRm5exGHZsa3w
rkPLaGFkrF7UZJlCZgEf7AA6XLJGpgKSAgZxHI2pmZaXsEFhFXadhemH58j0TpaB
pg6TvMBXATVFDHAhWDQKd0+sLYXiOeMVAerr4b8ctktlRraoW9vB/WQNd3QFOfAo
sLhsGdcbSKUInU4hx/gWyTat0R5WW+FJF20lTBUtQ8flA9SaV04YUnA3twML04UU
/Sjio50w46L46uaDYdLLxFbf94k/X3lEI60vmcpCJIlsnbK99yM4mzY6nkoZ4RaM
fDAdB1A92IfxYpULFTqZpeBsp7SFlaweak8RIruCq+/xLbv7otFySGu8AD2xmjb5
jkV92axLRS8lzFf9isvL3R4JL92Lklz9ojIp8hO9SXfTg1XE18XmUPoNOBwTvCK/
wF7/CNbLP66fEEiryt4YnwjRBkUHVlOgr/vPPVy+YzVLOR5nQVXOjWEzIBugMVfN
QPal1llZS0kzHrofx0YdzHtzQxPXaGWH5chT89j5Kwp133L6hY/0YJsVuJWs+rN+
uy6QWO44oQqIJla0jPhariQa09X/k0hGHonetlbaizUcY0jIXwrqHJ3jG6ulhoDK
/RashnDOuLTw0691SxqRxP8OTf2pboL963NebV4E8V683yMNEG3oxVS5Nux2E+J3
DAG8f7afwP1EVuowi2AIsGWgScpkAHRUlGNcIubMJC8UCBlmEZkZPup6MtHStBcD
UxTKjnvNdsJgbMl0eot0AWURnMpul+EPo8XB1O0hlBuEiRNlpCWIw40IP2gM/qCB
omdxKBqO0oQ7HDqZ+CMNoT5ys3S161/lYTb3PBvmP6nIUoz4xT5JKp/Fulq4wQcL
UTNIFyFGHLFSwCeMAqogJNRgzNKEpPtFJ6ahHPpX7w1Tr4E2Hrj/ACn4iFZn993e
3xGtUHdriP6ZB6+zFCjXF1lYGrHDyKFSPm3zIHfFOeXNFFQKLH8tJUdmLjtH28sQ
74BfuSbaekJIgbdlZFspi2RIsohfyRqgaWG02vOe4OF+inJxAQpYGbVKZck8zqZ9
odtyfYOAqTR2JwDx87F0TwmNiYBPE8ytssEHsIXEMrMLyDTVAqXPmX/s40vmupXU
5/euZa55UuByMatLKUdut8XJwno+j4rULD3+tUNZGD06ngd/xQiu+SYqN+y8dIbP
bvJENXe1MAEevAHj6CnQuqCG+zw33T3KnjFEXoOivqXNPFM8yOnrfDTI5TimKGFY
tZ/IjbVjtkQbr8b1w8oUu+oxFToED8r2QoyI3LCuj7DodgUsCnJHLMWzZjxl0m/h
8ULZxGmo9Xs0G5Iu2VtFvqfGzFir4fXZ4BIFFo2Di3/oHL2hWKHemWp4P6fXSfL+
melvkL2z/lrNx7+7027rv5eJnkoU7heNjhVn+AGV/ae4mMPWr7wFP5smlM9o6jgm
NMBmv/jRlVjlB0sOtHc5t0We6ZQPgN1j76IAD0+Da2bMwZ0k9HFrxPWsRKKiaZ/i
NxRuxt1DZKJDeXk11g7bl4veAyEr4ZL4ipq5qTsOnBGEPNwe7P54oNgUKYDWYLV7
yZ7gy2GulFdzOr6A+DDBVxZ7XTdw4IStSi1lcDRKI5fCKEFmMVF/ZLeNi6kF16bs
/YZ+/1fl2VExJ5E2o4ZiFgIYeniei4PZfbxjRXzO0diCRlzMY2m2fWmNMVGJa1V2
GVq4qObvf8x56+yR1tewcxv8b3hOND3IxUJ1dwrioDqAYgsRGDbimWB36JvFotVM
fMkbcnUfcVOjMjmcjmjK4zZC0KPb3ZkO7sR6Glg9H3ugn5ptLPlCe4A5Apl+Or6B
KS0bSfpnKVp22MZaIhHJtNDTs04KmUcJkJi0cdBh0zmWbFqanXssJPqOeSIPGO28
LOgl5iqIawtHO48WfC3lowtBsTfINBm8e1acwDSS7Leyh8IELfTM54RcRxP7Sb+V
Xk5ysGePnW5bMStSClBYJKJ+vPSDhgrg1LKDYH7F2wOQTCfA8MQ3lc26DrKsYif8
4JcEM2UbKfvVCllaljiCNnKRULN7ME2wHY5TPGv4Bkh14Eki0E+nbjLxd1sGAhcw
BA9aa+ICpui4S4FDIRWN0LuK/xaUGu1WHKXXhvrpR9sLyZgZwfbZgUTM314CgnQL
tDJ8fATR522J49d0zzLm30e53AEP6Valao3Us+vL1UKlVLJ/MadBjuOSee6vqj15
uPEZs4yTtnN1l3BMfnsbrRGwQK1pDlhEPMslVoWCeAxeq8L/kbTVn+b7qd3xEeKc
z4WYSPe5MR2VnPqqDvm4pVa7YdXmYHikXHEzfOeD9TkJECKDw3mfMVN7803Ex8Yx
g7CS58/jwGdOJh+zFk2fQ7S7q8KuOaDB0D7JAakbonlU8L9psWWL8sajkhM2g/LK
xDVah1hiWMJ/EyvUoJVoy56whlB4Oug02LDdMaNkuT35/+xri+fTXV9zEQkGv8pu
ZSbgeUKte8AqxXSLRKJ0H1aqtjrX1DAWyzBlqpqhEIeyQTAmkl+vvhKMUAb63qRU
Ga80Y9W9r5Bm+OIhRMHM9HS+uGkEov2RFg1qEoT7MIp4EHm7vUN96OpperQpvxos
e2/QfYSo0mFgFuWThr3V7fxfdhoC3zl4Zl4EJ9NE/dzCI6IDY1/xObCURBlDKrJ2
AK7TYpO4P+3Jn6TUUHVKNOCCIReDiioNwCpSXBI+2wARFSMdFQZPYtuP/Ph5kBXx
nfP44J62GhcSG5zQnmbIr2Pay8+qT3NqwD/PGSGFn8Ms0IrpiWpnYvcsimKug1D1
uCp9Z5jw8tppR+IojA+/bg3tW3K28L/ACrAApMNM+Nf3oxy3qIt1hmVeXpOWKtmr
zArEc2c/7Wi1vudm+/bI0etCnzwz+NqRaEBglGFU7NnOY2umBXspMEsO2hO+Dqu7
8t/ZiM8ILaj1iBQ2HlgOTWEoIp0J+EvfGX+4ayeHwpDtpX8rCAP1IHmCGEiE5FhG
Ht1E1hc/7NAtyLqPrD4QVqJg9SAR46RmVr0BREjPUG+5BcrzUJUhPIoSyXIyZBAd
uGMAqI0F570L/nqNfKTFRv8ps8gT6+CflotSfXgHe0UB/x7Gqz74L3upeP/8p61q
optMgFFrSZix0UYubWpJkcjpoFDM8afPtnYAwzYvYKJNZILYSaczdomuybSlyhW2
k/qbDVCyUFOzSpbIcaNEuVB6jmZpWcLdG05kaLZartUD7aRHPEqQNsIwZ0/avZcY
rXcsE6kDl89Pi2kzGw1XC5/J1yK2LzL+ZAIPM+cVp0JQry9Bc/3/voz6eWE6WGIh
2NwnzmgIF5FxBTFmnOj0x4YrB0uDXOQ8kn63z7AFdMvR1oI+YJ5+q+G4hhHyV7hO
nbOP3OvtGhH8mvb+CGNm72JWvBGHwMQyc5/Mv1e7XW7QlTGPqhjnKd804KPEOTtz
44xqEgw9fnrgFj5b7e0CFRVgp624MXqlj9M4sb/rsVMFHI8XDlraibtHxJ0Q6chl
XRbIKPVJjiDNnqugFrmrDk06Wqj3TVcj/uPmX68KWmZRZbFpsvdRPQ3lsB2Hkgwe
I8XkZetOMqDA1OGUrf0nDN1G0CySpsJX2zYNLUCXS+HlcyMuROMsz7icPcd1HRbP
CXoRjkbZ3YQwS12Ne5uh/0KUbm2dngTSNPFhBWXIV//JaehIkeeQKlVGIX5dyd18
85dl8nAbATLZ7QU2TI4fkVZdxC3tETTId6cCF5wa6AADheXN8LgoF5ciSYjg5SBq
oPcJxltaOHM/EVxFeAFSoECa9HRJkvrYKjjhlUZ/ULTqXVqkJKKI4GoDvD7iqtVn
AMIXwRmb67c4f11dehFMPw/n5TnY67Os+s4XPk34kM+wO7qpBrZgs2GqR86pkqm9
hLUcjG6s8aXE27VkvncgdD1VTHGq3IaY5ObyJzGbFSgA/Rp/FEdFV5tNj0Jg5N80
bqEdJgZ31t6TVHk+WWbNLGwT4dcQ3gn95RWw+FLLifqJL/laxbAswxOfkzAYNsNo
wtpSL0sYjAFnvq5SNKIZwfrG8hH5hGTWJOiYxFfxB2uJhFgiK+bBErljKCpFi8Ng
F+IcSlTilK1zrcUbNRKbOidTOwVG9x965eQBmxj/YfXMOcZ51A3FHg5bpqmHdWcL
ubrbD0Obd+5wHjnlQF0LLzjs9ZSEPxy4cVrr8dgq80lbIxegU9rRzaZ8eKUgQhT5
x047WeXf/j2ptHH7pRXXWPYG1wWgDFTeniwSYuV+sBYlgrFj5o1SzDLx1NZdl/Jd
2xUkZAFuEjuqOFe4mgjSdkyk3hP5SzHqT4aEVqzD8IkKtPMz5+3G4QRmqWZPD9Zb
qlB5e7nEcHUrkgSjNGOaF/qmsu6sDwmQCsNweChk489ytNp2E2iqlQlQuP71dJe/
VRw9QyTYhSakeo0vjKRuV43IMbituExwG7yf5bVyMG//K7f1ihn+AJzaocr8LpvO
AqziGKvjDFQSCwMBu3d6KU0XxinArNhdU65kT3NcBaM4q2BihpUDj6e3GUvCsh7C
sFDWKAOu3qHMO8IBN7stn9fUGwUXHU5cIFSCJPee3Mt1cLP2M0YoSbOKoq1J8vMX
jgm4m8lMpoS9Va5oqIWnYQVFD8fabYaX7R3go3bDnkJPsdNin0dfDQEDqFdcdGhR
vWzTAbV2TVBHvvlhgAVzdk92QPeMmnxXMyoSd75p8m1KypXx9wVmHsOk02IdgeGS
fJ0gzgWAD09SLq+P1NETIkxPkzlxyycqbmz0/2uheT1Lp5gpA8xDdAp6RPjpUnsT
+5OKfl+XjDYwI9YlBmuhuTLl6EFTQNJJ66+F7OCt1oyezqFHgv2MKgFZHc/85ndI
YKZyVeiax70Xu4Zn961CY1laZ567P5bfFY9GPX1lYfc1D7r1gpLxmZB2WTri/lxc
lD3Zo8zK+dUt4htVIgjX84AJjSt8tNjLHzpYtj2q8GY2PkW60FG/FNpKNOX5ofkV
yJTTeJ4tZeFpukjUWYukk7VybGvjiG4Ux/D3xvFHqBEw1qB6KhsEPeNygQTNPliG
BvPWsJGbxTjbrunJP0yM0/ZpE7nXT6NW65vQiBnw0/dbXRTIuzOAGR1gZhusGfaz
VS6dZStpzzFOHIvAuMZBXSz6B3rQvfadB4B+aWci1PVsQQQF/Vu+Js+vDqhHTsxn
WpnpKihXhfcLu8rmZevRmsXNHzYK2bQO4khAQv/iYimr+vTKc5CImzBloKiNF28+
Dq3IEljzdiun3AMhUB7+fKvKxD8vJcj5i//2IAMrPV2Ir0R/T/btZh/8stKuGcoT
5t1QMSVwFnolwgCjYmrKlgzMQzsEkEErfnULMM7D2/RemCr2OB/QQ85Dojw84VSM
W2gMgtnuSSrNwejycif2tlu786mnzPfBO1bSBOzFWStci/VR6y4A0Wu9M5cGrAtA
B7SQQMGJ8Vgn9STvWrFcH+TKQAWJtsr1cR/PKbbgWhml3FPhMtTkaF+/VAHYDLwW
apgLwpIeUWofw+Oq+heQEz+NWdd0CbKhOtcrfSZ/jUhMH+6XSCArRL1LiRaUv0+0
kqZhL7gEHG0G5dFrRysNarSizRYSJ/RC0JGi/LYH16A2lnDkQvjWqqA2Jpmq4Fw4
c9p6OkdjSlKClPOzoqCO/QEgBc4nCnPyuGawDNlC4rkfObq8Pu3ZvR0Y+zNWWQt3
qWX6AKvltsIhxUgWGxHGBILhTY0/M7b8GblX5qZaUL4R7CElMi7Ote//WFJYLEE2
WdV+81498RzBIq7HuHncNdiFfuJW+yV/7GSzOAAIszTPPHZr0lLirXPZIPh/7IYo
BVqytXXBusCcyyvbcl+fw3BfTYcWuFhqPnSxEew061sDqaHONv++/+SMle+H/lYk
avhFOpoEU6anvfA3/caLrSqD8gx07f5+To2hdsaPohUGFtHKARCFCmYs6mVgJVDX
x6cZ86gNTNBkr/4pBFl8jCnyR6oY8lPDZk0H+Y6kC8CLTqd47wVMGic818/AYCBa
2NySnXZcbkaI3577P1JW4+YzGcfXUKEzfnTZFUxmzaclXeYPfvR4Cpluxao2RU6Q
uWNgBhLDqoMaHWnz1rNyutjNd5tgiX9Kia1V4QL877AnSYCD1k6Yo208eBUuZToK
LlX9bqJdOrjGWkrAtoP3oLTohrGwN3HtgRDTSc2IQm8MvVi/p6K1MGkAV6qdpICf
NtK3VsIw7FTSxpxyMfqcLgDKpXGu/yCkPVLbDnTL9men9pf3FHjJxEvySc6lMJXu
9qUhIX/pJSzYdj7WNrbjLqfh5XidJFiXMQEh7cuRn4k2meXwxdf1jG6LzWPcpIuh
A6bsXUbXdlBMQsTCsGCIv07+QbQ+jroaWy8DdlMoXb6++9GtwSiwHxKf0nsoFfzx
t4yT1kJk0mJt9iUjQ9i8Ci0q4OnOf8B8CNn4kG8ZYdNFDfCAE5MkDLHEh5ON/rm7
Cmqyz89vwxrfbht1iEnXMUhDYv9WhBrTziYbDYmYjx4yxTaZuS8/jQna3mpiQOK1
Z3SOBG91brNLJUM/TcUiuz0E40Px9MfchJt26trPJnEagePWay7FVd079BKbJsHV
6oqHD8sw+BEl7u6l8Im59fTyaeTw0aPImXkH0XJ8YIq/urbQkLPgXnnztZlv9MZK
Uu6FlBZkmzqEGXWYc5s6lz+bRKNDQBMT5d0/e8KCZFZg1WnbqVa+j75IHEXPTPpv
QAMU2Xa0d4evMYkSkLqj6RXi8Wm8CstibVGRFrxg4G8p5G0bCDOMlIQOLxcf3LO5
4FBHmhd08F6hwUzaLTjSOxGHzHa3g+1gIsv/co7KyP4b0WWNTCsSkF9vxMod1raV
k9U0tFiFOYJbBEof5CJpT8KR4vLkjxaw+KTKmaBnCnwqPqr/48/SSfUfji25TuHJ
oWeV8YiWpBKhWAc9ZpebxALs4sDqKm8nR9C7CtC4/ned+Tuku2apGReNQ+kD6aqB
hGroD4sMwgnUMfuc2hY/jYUyCeMKAHl9xBmo8FPRwcDkCzDN9+pKbUMbkSTTr/s2
9ppWW3L2DV9tJiQc1/iG30FKkEAMpxWPuk5O9XB9hgkU4Df/zJUJ8ub0XCT5D6Gl
uegqbD0Sdy+YU0Afa5KjnWAvCcnOaw8t24BMVf5TuwWAEhYBMCXHV7Iq87HDj0z3
6UsKTaURyb+2EsDAKmDbYWLrBljLJpcvIX8micWbgNN/l9TZ9A+AonNBfC6eOy7l
24GZ7JOsgi0AiklIkcKl6ezC5N/KV6JOUHlHiUfWBn++EUpPRVk7g02gYYFmlQ7d
uJVy0ff+VT0uAF7wd0GYM1VMgAUQa5RuhQAehvCjfhFW9B6uqqc6ArzFI6bSwyar
IpsjAhLn8Qh1+6IwjKJ0aZO/PJveVqadNjeZoYD70g/ZTGItMfvTqqMUcsngEXUz
Zx2owAtAYkkYQSjVk3/fmFIjIRGHa2QxUJse+iDXV+DpwBDft0g2HuvHW4fql2uF
zDNmypq4Pwkt8LG3ICYxyMrlXwFNRjn1CIduR6B5AY8BotbhMe8pee0NNqIl4AGK
mVlIR7xHu+Iq5r8viYtISArPwceFnOxpR/q5Z69HcgByy1+RQroUxClmawf2HjCS
57jjPbP2nebrxm6cvKvwanRhDIBQdrULHi5mwjq//8ibOLLvlyNDQrffzJ/x5fVY
PUqYYYdP8m5EKyM0WZfWpWmu5iAVXjMGJB14toB7YUEoQd/FHahqTT2yCzH4v687
uFyr/HpJQfozk8YmzmhRhoezwf9DFY31M5IrHxj7G2i1dCTCu41knXnbH0j6yMBO
eR0D09i8kpG4M5Ssi2k2Vd71ZrTtOHdyA+Va3ss/tzArzGTATcyD94Guqik1GTMU
udTegngk+6n0PZ2Ox+v2neME06G47h0MRe/z0Ie4lCP84ltNxsUN9w2Q7KqxrvB+
zK7tSBxR3Oybl7YeOaCuFoSXXyPLxMcHi8hT2Favu7grNbhy7q+lHXWoR3Nkf7XB
5Cv0U/u9LclmcaFh3cZCdyH9gRzFKTyf5Dn4tfYZaOeOylBOyq6G1I6/n80N7jtk
W8SNdMRVaMTLFeJbZRuhNkp9zN1ZtLyyGF8ti6ve9+6hJosBOcrXsodxRxa0bNZI
yYBZxG+R7Myg4l5m6jKTChAVIgs92g0z/6KRLZjQE4c76zYv7afhdBdH/CaL5uul
cQDKvS2cShqXNbacKiUQxMU4C7bHDqxg5XuiL8xeCPJFQLiv6iwS34BQXlfzWRXw
HtoiYEHJhJ5mmQpePoC7m3PGb4/GwmZIZLljo0DZ1qG6NOq3iwYQt52orzvyfwt+
xn+4UCJ/3eEZRcLKFNkSiRgjJ7w9xix6twkX/KrzC3ud53e4WsgkxTjrkGej00G7
FR/A7gmy6FPlA1EtUSN/AGsY2WHZN/2Rl28EruGSkQGtpD1N6+PcnBvNBUwPjx7s
l3J6yIzGCaAfl/ByOsz6bgZC3RboqZdFdR9lhk34s0q+3qOMOh6dvLDU/2Bm/TEf
Ee91Ss43eZfAnZFREY0PwoOESRt7j+A9SKKkAIHIANyi5lFgrJ/XvY98DEB5GLs6
a/wqtlhfEczaGirYn5rgH6LNxj6K3yjriFJRNUL51zTn2R4p1dEVnFlMforME68R
5Ni0a8dO2l/+UhcT2Hcl64gm6VSTK4hqOdeRW37y0duEgNepLviTHpncw8kTfsvu
rg0YRLsVgLwffEHdku46PY7EAuuA55VwW7VVOsC+xRChrqUXYqlKvOrM5kqz7Em3
7BC60uDSSyvRiGpzQbLmjroH5TZEKKeh0150cKzVBSl2EsXTT0cIgDdzNhB+bvTy
QaVabjHX8dfcaMT09hsRrn0HnmusOkter+GiWg9VaydEDpMJafkWOz5KHabTjrnu
0QqOCIW07XtsXQ0RVI9Om3WID4EV0CzrOlVvaFjXbeAEvUzPwgXI7Xlz04qm6S1J
xq0P1nn/iiwxXc4otf2f6Oj0WfjR9itkYGReKlVPWywuy5/LSmhFOK1rRWJ1QWLO
Ztpwkf1TYMQ0dcVyga/+imDybGiJEu1fhbAOmV/2Bo+P88bG0iUR75QF7ml5Btv2
81POl2DT0KGBXQAQ4Y5CNlwtJZL08s9d7OyHvBzHOb0yDGWcucwW+u95ZvTKzhce
GzRcm1SefRVIj72LIKVtsaR3nAZPImZbFZlW57HiMCp59dMtaGV2K/nNIK90fKdM
iwLtrz6tbdYBYb2RsrRuiJR0l9KgLHcb0JRViXAsX7xiGZDnwuMMyvRnceuC5WMh
HfKP/wuhIoXgI+CMEnmu78gC5qToNxjiuuUMIz9zR0Oo7prS6H8sFB4F6ivYO+hE
An7YeyXWyC4Gus2TdvRkb650PdXnvut/KALXwXuXIg7H0xvmlvWUQDnWSpWE12vy
xpTdySwGB7cji3fhpXtkjcKtYPS40tbsc1lGeZ2ZywZeopzQnyB3qFcecOIA0Xtu
ROUlZj+6xNlSIeGvMHNmEXWS6Myzkc7SXXLWbAcDtfUxGgLFWPCV9dMETqT09TuZ
iUPIIPB0cGz0IEWqHQoNF+z/I74I+I8/JYGhldx9TMYyhVaAJ0btiIx3WhvCy+1a
iMP7zQZg61aBq0PGyp7R50Od6g74fYNLUKQ/vgIjU6XmkvchBwcr0XuP/RB3jnMZ
eKVWDtaigYp+iQHtA8PH8RQdoQKoFi0/pd40kYt3hT/4fmpfUoYH9/yMzYcpYxrE
6MDZ5exQD9AEfnR5FDKkPBxGEbJtBoONBjSzBK9aPw+IDA5Mp/HaR1phWyXEw+P7
Ul/DTofKEuiZCKP1RFDcnqfsOajYJzeh9bdFRHUP2eyupcBuOnjgm+HaFuuqeYTI
6mppOc+xOIfgv4DcMo0wIwUcGPTghmsXB2ibCJu4Mf2aC3iol5DMYc9wvHgAifC9
utDWJpE794JGD+TrOZeznaZlZNXh7zntgOlARGwK8xgHjj6Y4MEO7qEWAciCsfNa
GmuFtLwV/TV73cTOvhpHp6D8sh03UR8rpCmJbbdpet3CwcFSq8XJdm/9uzED7hEn
Vcf30a5IWl5l9tcwZUcMAXVavHCjCcIoVezfNinXkCTv6lhyckIYH+0VrAcWksYg
2476Hw+1gqcrqTRfIIWe+rbSabt1O370dPSF4E92arzZ7EPDrfXO+Jbo/Co9tqFv
DxgzbEfY8g4q0pQJNPo4ynfJ+fEz1cV3d4Bpml52dtpQAlP5c5ZXefTH8XFgaj1y
+ubTmPRu2AKfma0TLzsoAZMah7ssAqxSJZtHjWUuKP/quBB3qm5iOU5s38U+KT7n
heNCDZQtauR1Hc0MkLEtKO7oxi1OqN5RF70eZPnUDm9tj5JF15JmvTXAbvixZkTn
FulPesoU7rZOx61lf+JlbGLoeZ3hYZ2wRNgRNLPSxCQr6lwjSK6C+j2kzkONz6Qy
/SwPiTfoI5pY6sXsyxv9UeMWGDe/yk7Uq4BvdqtvpEhyX0bHa4g6WUGQZuV1TVDQ
jNTp2JdmDLIjDRmc3LieiqYGnP9arlyYYXO1NeZYc/jF2M6mEsexuaVaoKXKCkKJ
HRYL6uNLGTi+EhgOotvUpel1giZs4jJt3QrtlHeCg79gmD7vkEQpfjk9d733nu/2
JsMfuN/b4v4ab9JmSIahnRi106HzWuiJI02oZOvy50xc8E9wrrkGyUbSosMaPtQY
WE6O4nbFx9kSHsIvNcPOWbM2xcGgYD6GoOFog3H0hVBP9eAsApwbLdOkeYg0eVXB
C3BFQpcD7pw193fohNT6L2AG7zs66TknDgLWdaKWQZzfzgORrMT/wusv8UNDTiRN
2Uj556ZiqNFbxjDehST9zfokMMg+/gw4tHbGgJZPw9yAX2FR+RirnAtjVzBDY22f
fyD1B/QO31O/yTFkASquWf4+Et53AAwVqvAMiSxq+EIOxSLe1P5fii1H3JjTsAK5
x7HekOqCQeZMin6oxIwr5a5YkjmQJrwNE6K5/bJxJu/08Y7E1w4JeonejPa9NkUk
RXa7zLtoxjMtv9UE5DLXODrhFv3byQf4JKGj4it6HQUyq7fDYZzROjyybiFPb5tn
edy6Ao89AkgKvfbc+DBeh5tcjFkR85GwXg49xjpFY0PYtRwv2t1N30TrXK4pOFMK
ICVsnJYbGP/6Pz614YBDeZcNJWqrmiOwNpwCIHImVkR2hXNhMwAOVIJD6hgbWdf0
bEr9U4uMWshpG9IqY0nkDhOHN3HVg/xTTfKlS7ELpXEPQDt/CpdxOOkh89YtGuOy
8VH3ZuGpdY714526DMppUMFe8q4lJzgk6mp1g3qaHOKesbhrTz+cOz9DKVTmuj+f
YrPjMcf5ck9SAudXPqSsOL4eWUUdBoV1YgZwGtMdgDRFIbatFn+HYnli6tT3zYkK
Q2aM0iK9IdSAFyyb8foQNnF/pNQ77lCn5vuUj9L676o7GFIBH8zuM+qI+vABsslh
68nIilrkBlDRkTICW6LE8vnOTUuFIKALbGt89WhSZwBrT41zLCYJvolUSB0hDzYA
ahxWex0ChJETsaQdVKl3qYxAqUYg6xdQ9OylGcDVcpBA15W3wd3p5mYFnz6tPwwb
mkD/5m6ShukCLXqhPUgTngO6z8e+xztrm9FvaA7R3HhrVVQLubShSxFI5T/dQ+lk
2NtX2GN0KD5KqB8BIacOdEI/sIQj+W+CKPO6E1FKN38QrmIYfQ1QC2tJ4Hk1RRYH
J7Qj8RAVsxdnzUnMqp8PGJgdQ1t8b1S2sUry8NJG+ufnVz6jLxVZGtez/s9/38LB
H9xasdoX+5S3bs5J/PtAfKfBLTprkmhle/KWR9QVH87ygSHIJU/a1W5LxhsCx5sE
0i/nqzlcfKy3kjKs+ZijnUL9kKBhQJ7PTLRqsld2R9wXQZbLXF9LIZSyTCF8/qYE
y/uK+OoAODMfRowrK7gjQX4EJvxUfoZ3izsjs8JORuF8vDTRJv2cTLx8oeYhkAKp
/I38HKEYeDdjwsLGFYyw3dy9OVyEia8FvElf24HbxowohctgOBQprCHk8U7PBAZG
3ZK0vrzyiLoJgE6/P5RnKZCbA52ukh5bFgct60f9UVesQmgfQ1QxGAg3365mx3XU
AQQDJANREDYYF92HThYLwvh9kkHjNSFg/xLtSMROCiBRHP9wpJTxR4evmvdWSDxE
0das2ypHn3M4gyQItAcUvfvJO/zXWilPtd9AFF78e5ybsxJAuVCQN7DuGGhBt+Gw
7PIdwfKqUgddbo3k51djSFVsldKzxGknWQ4NH/hOJh849pRqakvYq28vjbkD0wm/
dJk48RVAXngV8nxBMcevmz2S43T9xnJk0dGefDwF2LmC68DdcmdUlSQlvy5kyoRD
Nqh79YSI3X2xQCYP+W6Yuv50aixfyJRepcPJGOSJtDy+yNUlQHJ3N7PKTXcswOmw
9CTzQYGiAGHcFv1sFY0ekvXChJAGGXeQsUzHnWq6rHzKCgI7hRDdfL0shb+p0bCo
rCzBhbHYs9WxOSlfnvFq/2yoTa/P1ACAD2gM/jgWZpHeVfZIqHVlAhNp4aHTwXhC
bNWqeIfPIrIsHHZIT/30t0/gHYocvrdxNlxC7iuBHyH3tbR8gd7//nkoQdQ3/twP
HQ/S7O2w3V4ToXP492cTa7D1MZS8o2H0w0GTMAVd4hAw7dtzdUrJYTcd0K7uPPJX
GcuP4dDSX40ZrcribG7LVN997frM77GNVzPSmJ2j55wCBnBSvYHsVUNjTS6mN/F9
Hy80mgAza6/QR+mvOOsoHrxrPbHQI22yVPUpvSMJfJsUE9tzVaQxdLP9QujP4wRV
kSKWiwk2XfsdkvbOZG0I1kCr2ZUQomb6Lm9QaFeJQosPSHo92Bt/JDLHw4zsgM23
shL0ND8q4USimAmdQOg6Mqfi5KoEm/UbCFFtIXhM56FwxRKSWL+hnEgiPLRSyL3L
2707hASq8yH4HKhxeNFEzIptX8yY1k5vsAD+reoxqmjcroBcYtL1P+BvlZkdbYCK
Xr8rHHbT5N7q7h3lNzUYkMWgCpjH2GyXVVKJr6gOKxn+h7JZxxo8f1WiLfST0Jve
CZVi6hOdCifG4lZlvpObDqvl5LvZk7CONEMdHycBiEEzP1tiG2T2G+PRqFoGOcBP
BWPXSG1x4IrdGdJ27yPuD6I8dvdpy3hj9TvLWnVIr0lkzCYNCu58cSfS+Wa8VbBs
jwyct48ax98fD7YqUcz7h/s94hHWgiM7SCvlNf92PaYx8k4fRo7X+/mPqZUCdf8A
E27oTFtjo9nheJ23ju9F9jgExteW/Xg35x87oPK2tTrsMc7i1o1DyxH7/OWa3aIF
KCK8H2wBYaBR/tuqCAsMirWqsApVsET6znSvIT+4l16AVphPwSa1y0xYzqL0+FLd
52EnEyNzHG35uS95fnbnNWQZF3/dSb7cdUO8p1yyyyHa7Xje3tKW/I9gh2WEtDtF
jDBCZZjbcPfadSaySY2CZZ6zatrpjMvgdQ+JP0uuizCT9zndJL7+8CKu6tQXVHDs
fuelbyVJ0EnLHoWLA3RZGAytCWBc1uzAYlmfrrYGESQTC/nRWcAY5k7TB43Ml/FD
S8OKoJnTQaRlxGDsIaOEcWM6CfJF3ANUEZMbNftIUlHGoFRJ45mge1o8NFGBdJCm
2QLFxcpXYhUp/GupkRDK7AkF6pwJLRvKIThH77uT/l/MoxWwKOoFCf2JYKGULMa4
6v8kNpnzkSHC3CIDplVFU8ehuA7gwANaEiNVPbGTze3D4Iw7LUE5RSPaH9/VGAnu
qKAK3l7T5vjlS31QsRQsOO8aK/AF4EJq8u9C3EdQIuOznN777pxdAPF6Vruq+qTU
ez1DQHOF16xHNKVnQ1BMQPgmxkK8Si3LzsbyFypcatOgz1KqeJKMXRNXkfCAfj8o
Lj4SYCcCOFQn0LL/YIYP6L4JwBVjxJ6XUkz5DIrSuJLRpuJnobfKuAjfpXyyp4XX
ZCBqr+HUBM65jH5sh6eVywR7o4ssgBFPqVJJlB6gQWlnfk0JJhhVQ7lOeyzuDE/P
mMrkscMUVfwOjcdUrjoI6azParMgWCCmy4FZMVmtH4y6ObOjgZKxxWl77Q5YWJ8O
RlL0KmJcFBmbn2zD8Cns/EkRoxKkNCtCKDsGibx7LHOlqehafjZNp/4v95mhWlLS
/Ux43eY6f6AxCmGvpAx47Vxblj/UMpMNDtnnlInqx0ydHgaZXkJ99LTHlx6w02Hg
0ObT9cZZKKOBY4LPQz6cBRh6egHq7mmAie59ofr+daH3CJ97vKs1oJK6k3swX/fZ
reEStBUSw1rcVdjg2OejCsDQ/4Hus+pM1dpw/FDeN/7vHWaB4txPBvP7M5/q/K0v
bfkrGHO8VRLrIJU7oF8HuGWkVaKaVz2j8oEzje0RFl8Y8XaZL3+OdaYznRygcyl0
dipkxqHhnUs0uFcbPUMg090II8aRmoOVyVAbDi9wxVnspH0Np5xxDBZSKA9RQeGC
wUME2c2NuMmzR0QC9eheODLFSA8ToZBzSq0wv18DhA8fhpNUxa61kluI3AXkzo4J
Ab5p8rAG38kVybFhz2taaDP5C6euIqkBYFw+w/NAClZfOFv/N8CceWXnHhCN17xt
3r7WL3ohJmjAOV9LeZNUbcJ4wdlt8zad69s7BVmPw5ZyXGlbk2RMRHTeCjZdhsG3
T8HtVjJk03HMctrxmfAOO6YxvWQ1F+bsdyJBewCYdFVLjpRL3bL0CPUrBtjYFtty
PIZkV6UUWCJzn675YUujgYkExXf0MaTf9XQHR83PVN07hj0G0UtreKmZHIvetIXq
yYQav36l7CYzK4CEGtQIbRll/D1pUqG8A22p1Gz4c18YLsgbFCkjRA5KcSeTMksr
kmXrM7DP5wz0pPpj1awmukvuyYDsVYd9pGiHKcItLN8s5kZ+c29lv4pNEgrRLLWv
E98J9GTAX8NTr6L1eHDnBZti+OLj9ezTRSObQdh/o1Pkccm93J4cqCGNR4N7VZvt
15EaPgKSIGsKCXdZNVNznCMGTlWm95ndYgPOAeqdMUTbUB7j6ocid3ogq7qNeaVr
dKcUV+4Wj5sDFRDSvwDopzIYdwOhNZYfrZh3MWe0/n+kGhksAgc+aqjdWgX291HH
N5LfELT/rFHCkZWOF/GkM1eAmFvs+44rbxmXkHlg59tnzm3N0BRG04Fvmsx/21B2
0Td2oJ4tbiHkVHMQ/BumnTFKwAgYt7PNN09V2WcTakVKF9NzYxhZ/Dz8Valc93Kk
V1hKE1+YrOFRJnsHjKcxPLXrczQlQLSfLv685sipw4QioH/qxS2e5+Rhie9j1qK7
2jD5gdIIp0WE8222kmMKzotyS4QmH4h5T6cd6muj/P+CAFaBIUjIOxjHZBOmJfPX
OJWQPNZDY/bMCrBf2lBPyiWKGIGUoPgz26yt/xRugysdfiFc3yPkGygNndcXu1i/
68akbv5Cw9wwUMol3ATud9/BODUCtwWKgLERo0P2eINJ8KR8zhFIZNdSfc4gAHaD
7bpQkkGvV7kwrZgo1X52tTZzltvdifh8E9aYL0GIoEYREBQCm31t/giO7AznsGPT
5NBa3mMQbt3iCQGAsrWZFZiNX/mJAKupevg9/V//ht2R/4VTqAnymvcfQtqmZgo9
6aVJHxt2WiofeS0oO8MVKlgiWbSurtXg5U4uoyVV5GYJ+Y090L4RvxN/P/Z0Lr53
lNh4PyofWyvpLDu6Z/bg3p8tUdC+ts/bFt1i8TthEDGTMn6UJroKyF82aHP5i6az
XcWjEpomEX+xPH8PbtLOr14WiL3mVnYkYADJS7Lgc9F32JStQN0CL16jxYQjFYDY
GDpJn2wA4aGc59kCbq9A6v6QFPvqfQyQrLtFirJ8jKWGF7ugSGzmIKnAOFGnOgrf
e75kQs5pjeMfcLf0tyVPTvV+CdJ5IyDVfiJGdlKHD7F0SYF1sAlW2eEq1+c6K1Lz
eOd0r/O07Rwr7o79hRYSbENkVmGYm9K5HmmAuWuhXaj0mrPkjEdUcEei1IymRvYm
IrGhmiNZvpUqctZduqVAtCa/xLFd4+ss4P88PnGmmnjM/aecT5/hZKQya4+lJ2ai
FqczEoHA18oqZ4ZBk3A5jJ2Brhz7MvsluuNyuQGJtQzMnnsogB/82Q7OTBSzWVnu
gO89kQ8m8TAsu0v7DjDEHLqW4jY5t77HBOKK/vIkrnkRQLj2CZt9lOHIviE+wjrP
iguTij+JXQhfDLQrXd2geqyCjlqhokpS42zyGTsk3YJI2AgO3ZnswyF3axPjKiZS
Ah/kYz2vptQI/rqaG76USJr4jvl6HEnC0o3IDdrXcx/V0gFwoSHBNiK1i26GOjZc
w+6Tk1J5EOqVEGGGaUcFgeN0tmJWZszu/1k3dbh0lZErwD2/65hl1RCYXNm9psq1
rEiKF8eerjjgAIEvUBDxv9Zdz+SxekYMpXIS8Py/IEX4xn+3yV7vEbcPaNE6No95
/AC2WzXY0x8QYzQZLXbHhusAA1b2DV5t73sEr1OFer83EV+oU+kKRczGID1bT5oX
PYBC5MMknFgg/jiHWVGLmP/bM3D0jWihQa7qL8T4+ST1bHh+/zZ2A9I3Las2h4Bp
zV7UvpyPTheu+O/7CT6048RTWn7SBhhre7NSzsGsmonn7uGtYtOCiVkXNd6GTVXY
YdvTAXoWpIkXZTejyVmLJj5BGKIF8CH3TZh0YRvZzRU5C3+NqFZGm6/2F0IWzWHb
ObfstPdPtnQZlU6ZbexQLJyCnZR5zW0Qu7xUsqVSBKt2qFlLKsME2H6Zs23ESS9J
lxFwNMUOqTA1U46hHk1Jz4wr7shEO4ppTo3mOsq2f8Jka26SYuKW76WRKMmL/KcW
FNhxbAEAw4IEXsxNusGx12w0wWzDSYSe090TR2l6y7orF39xhrPGOD7YCmof3oZa
398z2X8nE5EnJeGeFUE/ILHm33TAC/Rom7dGm+lfMUFXlaDqbsomkOq+Y8sBWg+B
Kl4OKtxA5yCveM6FMIsnu/sWTc7PB2XmFk3mbl9JakJU/vCE5E3h7tUrcLigHxkq
gLcdu/Hc2NQXJwSiqu6tk1ua/BleyPwD9DvbBRdKJwE+/MsOsmLKTFNWabJiLcB/
rBngNhI79AKv7xJ8d+YRKgy2M5sOQ8Y7VLP3DW+HD6ksdLswS6aLKYQwTj8Ylhb1
Mw5lcC4WltJwA2uw0osSjLn/YiJeKaHzIBqOkKFyQ3Ld0cHNedL4/nntpS+6POqw
VI6QOqK9EarVKYe8AfC+lWqCEb3afSrkf0NRoVgL3cjULiV8KukfktG0ve06t6lD
FcegsozS40wq24kQVYuFzAW3N2TgRrV+bWbRqixbWc7+J/X8fQYq6mP05T96GJam
q1TydoqkolkoXaQS6+R6LHxjCaNg+MVXkr7xpYvWR0sJBMicDdz2DwmOGTTa+GX/
IUVH8aZtTMgfrM2D9dZ5QvktSrBRErBD1Igtk06pSunPK/GD/lvB9TfIZI7VuP1p
3wyB+jzGBuzSHhAk5ni1ncrMK1v792tP7lVLRFTR4+LnQvP+VogO4tsQIlKf4VBX
dWXsvkGsXZ3s0TW3hHB1LXteTN2IhkJ5Es0ZIWOxdTC6JgfPADtXsH7jYebaM4VT
noP+CgEHRl81pGJ3nN8qsoeO2f8TgVnKcw6rcqzqbvLgefVCFuGbyqdmcZRLTOFQ
gtnDr87+/guZdfGso0lcQTV2BZsrvZJCnPikmE3g7QP4PZxEe/OmwVkT4JuC/gqL
kHDzj9PFlMIh6dwTF1J058+kAOCmo5maVLsQMH4lS+4B9m67wRWtp8tFSEnXCJnJ
ZKVtCP5y+3RGg3h5fGL/g8bZTuQjpRHlno8fxju3BpZ0TgaN/qNrGbgI6iaF3egu
4SnDXsJ84tgH+MqJXjpg+0N0ZYuhM2zXrpkcdi156iOnk102SUrKOdjV69acse7l
V9LblRiEXvREZYmPbIik5QXIGdhCPqDz4FwJSt8ETmT/5JFMWlVDbVjrRXp0yje9
bh111zJ+HnQdRfWEjpY51wPyNJL0nGut0LjYjv6V1rerJyfw02ZY0TQMYkxf4NHG
P/+1gFnMPKt2+gvxWMg34pE6JCSyqB0SKrXNE2YFK+AdNxA3hQYvHMVzWDTEE9Cl
ILMUMh9Yuk/BdMhiR+b7LF1GrYMweP4xRmAybJctGrQQCH0vriuchHlc3Kt8Xbnr
vDYio402NOlvlGYR64SabaBYxNX+ZGWgTI9lx9l1DSEzuegpEbDJeTVSXC9MsuE6
SzJSUJLD18wQbRtGvLYcHblnJQgvWVpRbtzJHZqhx52/ZdCoeG8R5FUZp0mRihcT
+C9Lo7+1WLShK50XcZW2dIZMls3/IiOslY0kE7f3K0iftsVqBHGbbmOXt0wCXtf6
sv/BMZP3TNuSnj4vsfeDZgq7G782sp+MFPLIi9DuPpBxv6sDgUZZsN0tTVM6sQ1M
uCS/oCSfF7wnxuE9l3xyMNIVAfnziX+iA8xmQuVryBAkFs899ZS1VqVcTejyk1lg
Ad4ia3CeCHLlbgowR9e1PZ5/NMVidFH/Vwqxn/RzdHfrBJwcueRi1Rv52bmcsMKD
eoHbrdHsezmvuC+C6ggtz2VulMQ5w2zOzznRKJMQ+g6rBlujgFk4N+bOcoUehV4p
kV1AnKGVL8YK+kTDHliaKWxOFOGvzksgVAeX3LVfvi9TxlB3/G0UtlGiZLHgJqBW
iE+lNMkfdXXzYNuDYjY0ntfUcWfVtoR2sRFVFOvRrLteyqNsI+mmVrmt48dR3Gho
KDidQ5PHOWYUL+5tDrVFPaEDpXk1e8Q0BdDiCV4K+W4fes9zlaEBoWcYZmDMraR5
XlZLa0VW8WGgc+awZN/i2mG3XO9Z0b7oVrzydq1bEgpPTVJ+sYhAhZowW1ieWUY4
1QM2rok05my6ftf4s86anqaNBZ3Uk68jvUVKHKNxPsTQN+XcBi0nt1eR/02Ze5uT
yOiBzL3K2eFz0/j7JwxJtj2zWGxpxfk/0dVKkIwT1WBCjNv0RMCAi6+ngGgJYORS
sLNImoLf5UvU5qD5rPTzJtnrJAiMTgi13dsr5o8xYkeye66VwMs1pru4VxpUeKSs
JD5nqyilNuLFmGmmQzN6l0tg1qOKehAY7cDii4H/AY5l1bmkKQwE98xl1fQwMEKB
CmlFubLdkJt71sfFKoJhIYc2vZqTPIbL977mPAwSkRk+9rkyej09pZFhf/PHztH2
r//274Uj7vBruKNLXTeq3iRxlgL75UygacJnL4j6WS0rTnoJzobxQqA842EhYIcH
Pkbpk/pvjHVZn7C0JVTdipPPODRxFWRFQ+HJLV4TaHJq5HBxBgvVAsSzFIgofbHz
b5eAWAZZb2wH31Sbxze5AaSL1Q5gwPCprdHMUUfstjS3kkLXA6SHvaPMOrvT6LX8
L3bLdWeYtZZ2LIiv9KqihH6ulkFHl1L94SLCoxzPd+1anfzbF4RxID6y8i+k6jXd
fBkdkf2tuOtl+5XUNnfWPjSZscq0WDY7Bqlb6zVYxwDOdUB1EKqJ3pSgeQJmIxsT
OePbT6/wAmJ2Ohjtk6t3bHTYxBYwZfktJuhv2qpbRBCTVbw2xfOW4nCS5WEyLKIQ
dE4viADRg4pLQRB+5Oh8Q4hxkcoOMSo3tPohocf/LtKbLw2HyisHeeKVmcIMiGkh
JAiTq/Z2p/BAYomMbOl3KQZfTgoqO0Mv3M9OHC2TU/7ULix2gaPh5xM9/amXe9AU
ewJ274p2/QKGK1jgq51zZFSk2X6U5aCA1Td4rtgVtXaskbGUGJX6YCo3nVS6Regd
Ue6UBDvSyF/YUhLbg4AmDnhFlRrpZGfEKaaP7vlCPD8Mp+leIak9kaLFQ8UIiG2c
pKWoB6egahReTB8ZOdszSNb5uA+Nm5shAk+ipgMvcE7K/ML9Gkl59eHhq5BScV1G
bvlxTIuydfg10mz4GF7nJrrX54NRGD02DPmBb2lp8KszAcPXSnFwXglN2cQJGe8z
tEoWJxu4mk77C4/9rVV8FT5/dxV3FPnR4J97XNImSOagvBLclKTAisJUV7JCaR0I
A4rqU8LsQZ98RPsz5EbGfmkKikAefw736bPiM704lLpScThUKVU2hygqmx6x0P4E
R+/QSsz/8yVGnHI3m3Lqi5Qzi+MROazEyppahJhjxbgx0StymEzvR7mDTR/ivGCK
bQiZFvcv1SYSMtjB9uvOHZYlQzzHBjs/wcHlydFMblpeT67wWDNKhcgckE7zXcf3
l0P7TLgB22W3Z0Z95im63M8NstRk7Q+6mW9FEx6l2zC3j+lejRfAkrFLYOgrqI/Z
sF2LYmxvnMvrDVwDx6Dimxnxy7rY0lGRYIA1nhDpflzOeE5R/rKXFphu+P0/Cul0
RZfEoKLPpPjjp0Bt6KLZ0ocIJIo2j0KDb8vRm7jVF+DARyKhw3+8j4lYNhLYNRZh
ty6LU7p6o4eoMqiGd1snwaTe+h99gRmvf3MARYOlfRcl60HNgi+h7B9umhhgYgdw
VBb4/OPB7+b94WRygoduO5P3xtGpnmLKk5TnRJJbgbvTqlV3md+fiLbtTeH5Oy8N
+EJDUxkLBMOorB7svr6OyD7iPOZrJ5tKpNpxoma2IVCHDviShxBF7gocAieDG+dk
KkcN+x45zhwZfPw6xe3yB8yR4wrVpZ6Il2BuzEkbFUuwYFyBgnhsivtdpKaO479N
zoNgvVrNtckbqbumhBvjouPsO6s3PIkzV0Bbn3LK27vyFUD/3KQ4PHCsNjmRbazW
WZfPlfQX7+eHj5UCTo3HypHyDTQ4uu2+YJFNQShhSX0ReLe7kFbQk54kRHPrpTvr
+Y7xlZ5zLnEWhz1ilsWEBuSJ9PrtWkIPhW9tTyh0WYo2cGeMon/3ohRoxkf1Ko4t
3dWBJsucaqLagCEhwG08qoA3tm5Dn8E0620NQW/ruz8vc+c9bbFznuzjXyon6AnX
RmGaEdWaffDqsi66jr6BVvsgiOyc7O4eoqpHcUzBjz84qm0bm9eVeFaf0eVbeHal
rLw09TAomum1QpUqW7KDvcaryQ93LsyrplR8daloaw49e8pjEFmIn9ebgWsRtD/h
6fm4dkKdRO5d97ujtnVR5LxxXxUuAkNN+cMTuV5QCx3zl40kUDCFZFZiK+1Q25Nr
dJaAOisQA7o6qJENVtXhGFYcvxedsU64FP7oeOheJyZbik/2qb/UWQFJSS0XIyO5
3EYyJkG69UmaIL+l3kDeb3u85FT3MbAmBN4EmcK5B0Jkgq0n0Slb54L8ahzSHXQi
O2PMa/UExLhOn1MUVio+A9750Wk+UJrJbmCem/cXBl/18vsYymShwFm/bEMWfTst
0fSZOJyInITpTTOEa+u7jqGiwJSENYytZqXuXuU2wcdTX+WhTkI7LIGW7CvLqcRE
iuoSi3xXrtb11BqHTCXO5O2IZ/HrEkA2mce9JrqyDnjw4mt+gWtrT8rvCT778PCn
cueyw4sgCKkuOZMsqPFXWCLvvKZ1zLR+SOBqesB6M9e0RQl1TeoWD4duJ+CO8QhD
3eAiJ/SOqVEbA9LZDZfqt16HFdbDGo3wB6DCs4qIr8DqGo9ghSRD+Xh6w0aWP34+
HrTfZZNfsE1WWLFVmGSDQdBFmitqFFY4ddEzTt+G1e5Bt0bIGgMTtJdSVT6A60k1
NL7fUa4tgB9Zk1etUeRbLChJ06NoBoGFds339TR8+NPT+HyD79a5Vz/zJ9D8vmdt
M8u7lPWs3qT4L2/tXDqSLIkSDlgu+NyE+vS5TvK4NvKcPzvZA3b1mIGm4+t3/9o/
ucX2/e3qr34BkzvC/53IopKspSGV64tHS2JeeMNGQVOhvwDqTsRmwrxXi3fWpwHE
+XKUvmySspjDTebTrDoY768cytVVpl493zSKN2hBqNlmxiSxOTTUtTj7Iqk227f3
QwBZMV7itr8htycu1kHcxdsQhFkai3od9fGbJl/q7ARCnjQa+rey2nDdn9j5I/6h
OshgknGxtsL6eO1GbiFHR33V2jVIbObsGH4anJ/YavWLIFh38KSVf4G4zW0juhUK
MoJ+TPYKpsfxVIDXQ+sLemQ6RgvH6pcrYgWZzHEv2+wbb71zQK8fm7omjpcpYn//
hRkZGKs4Oe4yNmsDPNH7PwGrzJIi+Xdn4gr9TSBdSPK3+11Mhub94G+bVCZ154Hi
md0r4KLBmmAMs9TdScaYyrKVfTUpuZK+nhpP6W2U1NluTst9fh0cm8pvRnz5jrNi
o7gza2WqkOj+TBZ8qTYryqu59iINeWQR93wDB0012IOhvPD4eUz4+cx4ag7kg1FJ
Ehf9fp6yVSgkhnzr9I5VG1CAJe22vgaV76UkvImgtna+S3cak0P37aBSvZK5N/vA
1OMPLZwLiIyV/vtR/W5+uB0YvOQXSouDdyJu5bKwciSJr50VXs/yVSfRbi3xxnfz
az7xt+rJlD3B24Fg83NcRhHCbDr/fDoU73EVpOfLfIW0PF3Jj6xT1/+HkSD0rM1U
WLsKw3xV05bo4QLj9TqKgxAXAXsAyUenav42MnqeXgTyE/NCLG/36s7hh8CAYokl
vd7PFdwQ+X7rlmBywBniY9b7J0iff+f6HYv6sqggVC1eRLto1cbmpDk6aJSyyeCY
09/atjGp8jpvXTa2ugVB8aLQHBkAc52iT2HoQnr9SRXcb0bVhWCZJC5zqAzBEApX
CwVNzYxkkMffOQ8p5VTYPAAy3lb6yYwV7PFic3sM30XpU6JA1cTWKl2hgdVGNg0i
w2j++Qii0E3ZaQgdH3JCFyy68e1oRDHpDEUCi9sPgUEZpl8fO3aB8f+v1q+w8WDS
cC7FeI57CePQr9i6qUdMwu0Gk5vdxX8xTsIF9r4qMIVvqxtLzBZDHmRn+siee/pe
qh4VADB12fL/JQLTUM2eo8jfPITR+F+dcFffdAxAOAh08e1/tH6tXAMh0l1bAVdN
zLzR8QmgGS684W3GO9bYtzCPmrecj8zDYN21lCKAiaFKIa5qDr3lvSAJYTIh9ste
EC1CM7yeIZDCvt8Z8iOwL81+/wb4l6CI++gXLw9cUNI0O8rXPpkivsy2Dd8079mQ
FgKuZ4J5+jTt+wZKhwXCT8qQzQ4Ui2pUV5c39kmLxuN2LhBmcK+H921HsbxcbeQX
UpL2ZwnJUqRvnDX/LIIe6L89Hf3SX7KXEvh4UNfPeMdI39kxnEPvxTA+vU+mIqsy
0tpC5qSMLRiN7nHA+ocz0e2ped1Ocrd0yapOACEmPuyfHc6erjbOVTDf2mDLkmxN
bWPlKlfylAtmIvdM+ZWbxY0U2DJ+I8eZIlBIVC0r08aXWQX1xr4Wjza0ZHx2B+5l
Y8gKze4rDiMTKznMMB9wW3eu46QIr/JmwGZ41AG64TbLeTkdM4yYPswpMj/0eoLV
boRnC6jyglE7jq2q3qEZx468tEWFsSoOQ2BjukzP/JSRmvw1TsQBRSPQvtmelSLj
0CjFgJoffmMJm8jQSq8Eh0j+fRcIlQgcP8oT1nCUJXZPqYKTxLCekyVrOa5/8fOG
3n0Hrz94pnrRJxvMf2lY8XbW8zHqXH9vJuYVzgsvnxdear0anzX27TJiSxqBvl+t
LjnKoHf+5EiEXzSryeA7t7n36cMCKGQf056jkAKk3/mu9pme6qyniPzrfx00e48E
Jm0U40TfBYFWXep5z0ELVCNHqB2ixyLsqIBgEkiyXtEap4LysrTPzLf+eOycLPJk
nO3Jwvb2n3jDLGAdgOeaA4Cu7TdYRrh4xcINVAB79omFqE3EDWCnCHEZiTDvs+pn
nG5Qnt6FRwGyJIj5FL4JTadoBvY9drp0bRGMI8X8NwyFAqymMY8EoUd2egy/z47E
l6+NferT0vOID90M3y7+0U6HxaPphQiACmjw8PC7f2MY3ARoVHrfZPFjCnLHhtf9
Faxbrx+Lri6W4l8uLnLpGItdkk3eB9trn25GEyOjv/SOEOIaAyR+Q+ZxTtLQcwwk
x9tMOatlLK6K1ZMkuUX4/DtMN3i+pybWxk4+IVPm+fmR0iOWBjZW65gFWa3ZYMsL
r4qun1sq/G2c9QtoC8ZCbuReGzKyaUMyUAB7qkJQRN/KIXKT/Csz+qOPc8cOGINX
lNjS24ZR+1B4/i/47P1KVfpCuW1cNOHgFhXH909KPskLDHx7QB6tV2QL+/XzxAd1
Ki/iz1CC81KGkiZJ3LGizB9U7RvbYVtu6yIv9v/sesRPm7H8HhA3wIB5nWbCUYkl
JfWvlZ9KkheN0orXGTb9s2I/xvuE958RLfEmZzsw7CvB24qI/EKjGBi5+Pzv0j2U
169JJ3dgUEF9XN8pWio6mFl1WJWJfcMJs9UGazdZiCj29SbGDsxS0dtoDTc4gWT+
4xQFDCJmLE4Rd9HrXYPcJv0P4UGG+9tk6hLpwmMQMzvT1BnSzwPT+tI8XRM9nzhn
wbaU1kAvSAbS+bo/hvoCPdcUr625Z45KmWn8oDAFgUX0c8ypznrJME9lEQHuf4MQ
CTjIy5wGwV1qvvLPkKAK82f1PQ8biTZo/bY/pDfaAziHBMdqqHCoa4zaK2cHhIWs
w0V/gYocF9tghWoDZjqEnAGaCuG/JrmOHr0QIwIrKKlyPGhFIqZuR11dq5BmN0W7
QEG5yYqZTlI8F0Xp+mV4PAA4iDGPmPokQCOQgc6lln0XXxPSJNfQM8l9juTa4GKd
ByVq0RtnqOFP7EylLvOZGx+7mbJHN1/K7rDIEKVNvWy+dv9AJarBZ2UEvXzCMWw6
RAyx4pOGk3AOORBkKc1XUyykf3n/QH2WRQOmIzoC3VVERTzgJmHDZeF2mkE3TcQd
7rKXuaoEep2sK2EZC9ZmkCjzKPEpVgQ9X8XQBPL1U3EUCTAHwWWAwh2v155Al8EY
rf8fN1tBrepkQOh5Yju+9jeBAke5bdvmlarDpJeU9bJ+/xJAqeM9LHrAiiThdQXo
gBuPCQR9ZvMmhU7CkJ6TvRc1DZXCISDwTaKKN42Mxt012DLD8pAsxJvP03B8pX8Y
7i2hUn7AkjicMYU2qUtdB058t3KTlInSU4asZV2BQUOIfSJztgBXdTJheF12pWRa
negiNOVdWKY2ADKrFDaoGhSC4CUBtnK8mrm9aVgKXARwcmx0svgAc8LGCLTEMnMZ
3Fee+kUk6M3oAzvK474P8AIZEpgZTkh6wMwjemRIAAv8HB3GGo+Lh8tzHlMFqpTE
35zv17dBTC1mbbEJYvNniqRGv3AkqVu88i6tOHnQX92kHon025DAa9BWSNP8IuLC
ihxz1nICfejV4WfWHX0iXARjwSD1g7NETjQr0tu/L5XsozWW5plM28JXm0YzqGGw
tshwBNbxsSph1xUTi8L61DO1/ZLrCAeJKv9IUY3N1WfaCJkbOt0duXtsqwNbgr5v
FwuPndPvMnpxLaSX5eqxWwsxHKR/VyU15oAzhm2dPvBiMpNwCS+0vVkMxgmQJM1g
gXFnnFYGYLkC9vHqsGlsFPIB6JVo53SQ6cDIj/Z+zU+QMnVUReVY6Wyqo8d+Dm+R
9yvB1sikr62YZXjAYz3w/DhF4nk1REz14bYH3PQ9M7mcZ7FKgEY2gXe6Exqf1PyZ
D8PqxbkgPIvZAJIpaRUHM/2KAMGjC+16RpggDmGsSph50ZGnl4HpBIA8XCA8rfuB
gbES3WvFyJeUi8qq8j2BWzqVlBpSXtclxAe7Tsv+F7DUmIvIAcmKzhlF6tJXT4oJ
jZM43IKtFR20Kktqvv7DYbKXbfkA5jAbJZGcP+WfGaRkWsJ7r2nDuXoyOuOBdB1+
fso1pcZt5tbp7+r+/yj1CAT5CvNfDqorOVpWT8bOXX9j2knovhJRKsBelAoZrr4q
NiAghIPeAYxQ6eAkx0VpZRC02VPoQfDQPjOt6A3JcUSYjyxRmouqyJmUmtUsF9Fg
jvUQejBzalJDihvnxTKKkmBIGbhI2yVV+Yy9qUy9896OS8q0+4OYUEzIQ+sbF9VE
gZuM744rNLPPQsdP7tg2lfixjVfh7oVkaver4h5XEHAYmcF7jPtJhEzwFeVEkTAd
WqxjVw/6aYeNr8hEXtCcliUviiv0+LGU20fyaSxm9TUvV8624mT8+tgdtr+nSo9e
hmlnMuHdrb/Jh+dKqTENKt3/MLNsCbWZke7GQOpxi8Wnq3m3GNxFqC2BGQQ95Ynd
IAhvAKRHFjY5XOz7MuQF4UDNqoTnvbvjPr9a/jx94pw6MgZkWRAVWEPwiyF5udCr
AWtUPIzkU3sirOj/i/w1+VQnuqe81uPnXXgwjPoNiBQJe84SIpH5TnYqZ0cN8iQt
D4o7/u8xvlw2jnbJBxFTJOxXLDZWuCAAuz8dSjFevB7gvhp788oD3WORrlVF+Ut2
/pvYrFLYomDTXxnEgb136b7NLjHUsYU658Q/WssuvKIj4GHpG25Y846x9FzU/MDl
DajB+fjYlTK+vqqOpp7ZYsTfDgULwi+yc/j3DlDbzOVVYnvGYsB9LsfKZby9/hfp
CX1w41FxhoQJ/vbGtyK7kMRvKbZ+YvSkP7MFeb+dYrt/7kSqJbqSmBk2qNKl45oy
vWsSLlAnwwgCizUIHdgyJ2Lrda2mLpW+UsLVCyyBrQvSm1Am/dyfYOKO/3gibCwQ
3yTn0jqoOiVyuqVrBIWAB/GzvlEkL+r3ve6bU2WyUrIbOGCb51U7O4oofENLLaZf
Xz0oTpwsXRQ+PdKXgFefk47Tx/nwM7nTQ7bUc6LZaL2OyCuM7N/0pAGQSp1Cwjh3
zRZ3j9kOccFt9vQPr/ceb/T5UovU7y0NfWVI2tgJQG6KD7McvndjNaGv8UPpRdUy
ZJxj/ppFfc59Y+QGWkxUxzA/jeVWIHQEIgNBZ0muIdPPVTfQgmoeYKyeQMIzR3QP
5qmslC0UFg0QnVWKd9fdIMneZqYRTeZ8UFhCbDK9Lxru/j+EafwIBJl+IL0ZnYqG
PTAbk8rmA7XWyjRpJMYcD9itQo5fsMLMcTmJUhuAZVC6jlgyKzqrsyL6zSiWVwUd
S8G/ZHl5RDzny31qVt7czJeJeSs7rwupZrkS09KXYk7lgoNm6rchFclHIvIGuNIe
uAe4VJDmzK0Nh76YUZzCrCNQyvc8Fi7zNRynz2q4Og9RPFsLPbF+f8zlFiFgw1R7
xJKxZutpW1LdsrxzS0AhddhSnXjUNnC0kA4FSU60cisAnyzXO1g6NqfKYdVrelKr
RIe5x+X4Ba6Qd57fmENIJu5AwOLDCrGB2rwfRPdVbO4JPZ18Xkbfj/zoYCh7dP59
YSm8tE5M3aCVyv67V6bQ9xwu5Oi0ZJSnMXStJSRwrXIQBumQpXfA0pDrUxnjg6iO
2/MsidaBjj4kXDJB2RftOqELgRiUMXbqDA5pz3r3rGUfvnA8qUM7/GjVtWn/YK5t
npeCcytzC7GrmCscKT0Pi69Q6nHIEiGmBxZeplCJ4M1Ml7oHyKFpwuH7ojai8pip
wTQtqO1MEi+vSl8GokUW37lGqrd7sLkqxYre0hqvxFB+THtalHWKLoJX5GVs3u9Y
RUV1dPMNeDwCvHo3EUkgZKUFjKebps/wBCYDtW+uTw8nSV8bdb/py6hK4ak00oUW
2Dj5Qoi2lpgT0kwecDiZ/j/fqKoDqwBWQgD+oYjejGA7IMgyWoeGeS1vh1BZk8Vh
Vh2NUVRBL2sdqjp8colJ5VPZBmnqi9TatGAzHb7igLoT6tJ9ON36XHCYebu2Fs+6
hTR/PY+y9HjlTHZnMUEm+4qNBHYbWamGsREtLiw5dTK/ReLMLcesEZxZ5V7guRQm
RKABZ3HB/R/pgL8w67WYHelLLvoE9cOC3n/gKcCVyyEe7ODsUQI0kA1KFVj9AVyC
wwiKVfQIikA2qdkx4FwimkkrdT1lCOJVJ3rpjhvzmNoeztpxaJwqwh4SuXZqGHrz
NuqofolJk+fw5hDa0qWsO7Iu2copO+xVnoyX2iwOPc4k8pMyTf7A7MBjMHvcEkAf
ua1QKr1yMvWBvf3FfyS0c5/9N5XHIAoE3DuOc58OyLPq6E3vUDvBAcBbz4Bk4cIE
bnOZ5jwmqunul5sPwGStynCnKZ0ywU0OkkLlPdeZK0zS2chXhLYrNunVAjbETccT
ZAU0j8cmXtMpOgaUKcwDxiDOLQ9MFIEmV6l15S35ePg6SjHaIxO72bvsaWIZNhR6
KnNhsh1KyjuEMFB8T3u8r6tVL5WXxS88kKwWJjRqrjVLf3HHwv6xJKkqc5JQfUGk
yTSwUiVw7IyCgUHYrcrOfzuEvhlLxdY1c7mxN9FI75CVPNS5e8nfNgqK2Qr9eXTo
/D0CdUdQ0rtu56BRwhEoOF2ibTYA3OTwL2FsXmpNO2HR10jHR660J75UBhx97arH
khChNYGN3Z284ytiO28znisQcE6SGeFhrT/dj0xxza01TA2s4HsQppdQyVpOMb5G
NbiFZpehRd9aXD+YERPBXuE0Egiek6kRs6pMXq1v2LjIE5rd3/WO+UTzyZgKRfvS
VKu0cA5Ssa5X1mdIWiFfi3nVlwd/yN5RwFLMRH4J+i+FXFs/qyEsh3wybQfcTZ/b
mHnQZjhS+q7uM703CiM6E8nrcWiIllAe2LFZ047/ghtQuZijrz+CmU19x9Vvtej6
HxvatpMImn6QVvjHpxoHA/xys5vZYhOiImT7pPH/OB6yr6LJU3R9LjJTI4D2EbSW
8qNFJLkrFmP3LUMqveEY5p1Y+k6EO2WPVQnXiDPAjBqFqTj2iACfZm8FT5tu0lkt
ztH1S5J7ue6H95LBkIVoiBU5s3DBC2A/azFXUdVECBIt+7e0IKtxqTZl+hoQp521
o4q0iR7MgFqYI+DxW2jfjDwVYmbxQ6wITNSj5zhs493a4zxkpph0Kvxo6IgZni0W
XRQhWfUKKycby6sTZDQD/ZY9t4gpV2MVmA90WFFVgJGLxZEVHwilPjujJYhxNWNJ
Wx+hYBCbSpf8KfWpNfh7+qKO38b8xMkl3tbfe4/YwNGtoFyDOXsIPLWYs1WcGxb7
YsnFYeab+I29lJ4SkBRfIXFUiWqNV5wDp5QTVi31LSDrS4DA1EM7sjGS1kBWWtkb
NcvKNoGVFsQvUfH19f8mNLNCSp9PWIaLOP+yRXzLmbRL4GVwZ1NuFpImWnD9rwr3
oTPgZjUsI6o1gbg3R994DFsAIoM2whNnbNnIS/v6LSIfUDGPn2yM3Q4GcbiwKT2t
smvZwJEdfrN9qfsxcAzsg7J6ypKT7vRu8vC9WJF982FfjCDJ+9ss5FDD4f4vJk2d
xWj0nQe9JK0juRAHv5j1Mxe3Kdb0kmh5bwveglvx4ZZ7thFZcog7eCLCl+uxvUqy
teTSzysUotJt4XQpM45tlUr8Tbrot2NSkwkjhMeeDHvXd+OvfoQheDRJQjju5ezZ
umHSiaDhUWBQ5WeRPWDFSHPmMIqebk7m1ywcr0sATIVttt4en420vSfa1rflZI8m
aWAM03A8Bfu8sRodqH43NY7PwGNZOvPgf/kiFkaHhoZGZlBN4MBeqA90b1fTdX7a
oiO8MQtzrm1N7BDQ0h1hhgHiTl3VjBmvCzrrET09+cv+JDwAfAjn9EdGwZBrI75m
myDHkhh+t2+HXVI4Z6IfzwmfwlyfRWl/1VyEaMAWubA81rJ5OUbzmpJ6ECJC2Dty
LZDrJ7dTTTaQApyj6AUNxGD/3U2jkU81aJWZCrN2XBEiUX+xeMjLxJ3EHLV7olaM
Lk2mqqag18pF3pdkcybuCtdu7N7M7K3GS+J4K7mg1P3+1LGhxKLUzTJjq+P8WasS
OwxC2iF+q6ZXKuKqO7sGJaIY7h2oIYagaRBzBjeiJpITDUBMFVWN4OX17ayO1ukJ
AE7mIlcZohinZnNrt8E/0mJV9aGH/FMFgCqcaEGAn/eaV/irUR7DHZW+JbkBQjqC
9M2fHlrxwtFqmBfMFxtTHxzP+JSmL72JwY7ZqPpz/ku3pN1kDjekj2XyV/8DTN/w
I6xBW5NkX1tEdie4BZOgGY36ui0ICuUA7JpU8EPkoZrT034oYd19sp+ZfsYw24JE
31kaK+vd7pCEVzkHLazoTjj2t6hhDsaT5RrUTOnBcCAT9bNQ4PueWQsLwW8OmLI/
C0zGcpFwiye4Mas+nwd/TUHE7QyQbwxY7ZI96BDpIpzgLoGBmUz3tXDjsuPNwg1r
MKbqXCyPOv4caj3kqnKM+CwV/PTYkPolYSAeYwraVRwpCc22wEbl9j6f0PYMQnH4
tTxgEPvac9bRIvUE4SdzlVa8SM/rcIRz8typa9B5+T6rNTEb3JaoU7SomC6o8iv0
bFKTUgTKKZYc1tMZb/4uf79ThwAIovDJfVjzzQX0KARatV83hS4q0BdvLLr2PiG6
wB1xGv+caf6VOKjMc3iCLvtJNNd2ggurjGV9sgyvEunJz/dv5S4d4voE2MyJ6uiN
L77RpNi4omxi5/UylzZ2Jj77OdbMHrZW+Aq8cLX6nErf8oMzoasLjRZKS4BOMF8/
JJGY1cVBVf2nMRhCRhkedU67XQwvLO0voP2YYxMK2oyzTqzCOy3eiCNqLuUqYNbn
Fa5yVhtfTiCIhK1RJEAsk/nKHLVPwV6zY3k5vUD38yNQZO+GPv8j0V8WHrFnTP9l
+tVuj3H6VwMz1/50mVpvxhSJSSaErRidoWsHToh4akMBd/rNHghcv3Q0cfrRLTXI
LPIsC03QtAjEk0sTcuZ+ilxYdgwAA/7ExOGUEDzVgkcIzhIefGhrZO7edJdQJBrw
Mu/WNgW90Wm+VvP50pehmlnJIoKx408BDeADxdFQBdDe7O+aSZd9AMPmiZGHWSMr
stFgKRcVmmAznYmxETOjgUjMo3oLt02rU09FSUXVAkmfIIyiltePBDB7IAfHk4Y0
FaM8Rku7XNMQr4ypNJpHPZtkDbPzMxupW6Xxp9tq34vbCbRWUXalJjaIm5uoi013
U9QjIOJkeVB8TO5OKL67orGafFKjp743Fv64T3qfPAqgyuPmbxGkDRm5lnBvuunr
MjVEfefwLKG9hzOgkYc1DsADylLkmMtrgKySkHiRFgI0agOLDw4BRElxx7gRCIw6
9C0/V7FVA4NSoeL4x1Xzogbxmcvp+Lg5zjo818BY9eBV02ghNR9TioZ7ttIlFiiO
u2pPgnCU2F/cnR05TL5UsalSNoYRObWDgxloA56pzajwJOpwm/kTyFpiB2HGO7YY
GRdvoFiJvW4UJ8K3DndVy41l84mNTg/r2adXmd9ljLTXXS20HmcDqQAca/RncHM/
8HWMDQlOZzf8Pa0W8aZfVqbEhCDnLM6CLcC9yCy3l3hOaxAGoFUwGg40Ngt1qwTy
Blm8ieiiGEvs07SkrgWJCRTwemucJz0pRpR4Je5wFYWlcpoe1JVngi9X8Gj0rtv6
6I839lr8ASYSwy6qWBIbuAFz1GXGqWxUlgSFw5aT4ghi3nvJ/smenQK+3CQw3h1m
h/h7Y+hyG/zCqIzwHS0pokGQ2FLtRHDg+5eGVPDNvCjMxr263R3iU/BDYlxP02iC
uanAMdiklJI0I3WzoAI+Xz6md0CpUUsaESGpxtknKQBBVfEmkouZXYz36MoRszmg
y9rQu7su0lAP6YgWD8b0tWFt+429LrwWab30uPF+WddD/79FwUnZuBLsPSAmX/Fr
OxgNCsHkYUyKAG1TSlCTDQw2ziSCHQkwHelNruBmwOeyZJ/CIML8hSP9X0qwY9gw
Fqql8HDWmK3Bl+UUW5N1wT2yx8dN4aCKVKrSAjOPElPxQyPr5ISaKKK/xEbGetv6
aBGrIdwv/fW3ijrusaLrjxpU9EJu6zv1c0MV7pX6Uhp6Vts/Z3GHIOEZlDUuPkMV
iRwG7S1HXozNqaIwFsIuogg9Ns+V4RnstVkOVJEbIVvKjGFrTAJaE1lKi/cvn5L0
oWulWIDIV6XcM4e1/9jV34HHQk9fkibOQrTOUx7TPAt1QqU7uyUnC5ru7JqTJslN
QjdGZ3x0NyhNeyl2AWdX85gURZ/CS+ANJcP6NlPALLaYEOGwRZXiK6Fc3VTpYIgj
bmWGHIAiXSjkMl/j2lmlgsorF8M05eSROLz51s4R/vU94eL1p1wDMdS3AWDTGKuj
VONaC0s3EADpVNEWPaPFKzpKFPRMxiHVKwwQpeVnAiSx0T5eJepFl3UW1ERszS7R
a5zyUVgl2ylBl83PVkHFlzbVW5tL1trRKFVulCpvjtvJ6H1fv3jhiABI3M/fONeK
arBsHu3ffH6czrWi+j73Z8zW+PJTHCzBmeFCHEuUoTYXdu37DoedGMFB4Ahg+v/R
o6uYrNpfAtkMjnxt3a7W2auZbVSDfkCZuSmLL0I8MnnMQPA+f2LIqjxfYB2LGofM
ntC/zOG//s8t8heWdLd+jMpzMsACBkB1iNFAvgejVGRNMBR1yKc9bXfpJjK1j5HW
tEhgt4OpbIL6mrelgHjB7PgC1sovg6YU3UxpLU3wylsR5E5xb0aOzIZJ4qafsQw9
OC5y9Z2hicnDoSRFq5264Y8qsf9Y46uueGfiJj8TyliujM+Py9MfJzxdpAlm8J4a
K+HyyY+p4wNFfGqGISi7JbuY/6/22jlo2sfpiv8ugWB5vNx/lLa4HdOAYDujgwRk
Ej0YvROUKhvse1OEG/c97omzS1xRh7W3sz7LXxKTpcPQw5jWZC4iYQNdUheN+mJy
bchALqi7zaKQZQUjHeaX1cLb79761aJRP7xRpg3isdjCS2YyFNnAHWFCwGPPj+FJ
8OlPtMytTh7VUP6N1goKd8W5o2cfepSmS86gkCkT14raGbtVty3jRmYmQLtHhNth
G31mwx9kOx664NNFeQoeKwfI8kZUeBdQW/i9l69cQIgh5uXwLzAbYrnmvwTxI3EK
Dx1QgAtlloKGQA+BOhk27IiznHY1w2kRMA89buNaTUmu/pLVNFKYmgj1j2nU6BU6
FaG3wg/cFBFIJFYXAPR7wQWpKoD+Rd7tmXjesKreIyeo3Jb2wrPVLxRBu8TEOcL2
tHV8mENTK0PMK7Il5O0LlgUYBgkYCTk/LVbwcH0DkAdYdwUZAIJ9hJmS02DykQA+
NaaeLBvnQiDQPFJP3it1HFQGOgngmV13TfM9fzPDq4J2SAqanwXEGIHRuj1bpBAK
im1m/g2qtXOef0iAelq6NOEdcfKSCzi7tI8D2pT8i0riK3Ly9rh5TjQWGsNRVYg7
50K8Ib4EypsdSabIN5GcyoivdVO2xn304hLB43l2lq7deuo5FDSHqDgUdwjxPVBO
hMSQitnzVurpW3cq6i4hO+NdrlwoReD9eP7JWCWjAu69CdWClSun4xKWNvwrmGPo
5/AchpTjtEOpexh2VbI+OA+eadL9vKexjly7IcTyxkEEzvQBj86xtp2gA+Xa9hBz
weZ+2AiVsVT+nM43drOYkavLsbmFAt/9dW0xZ4iyCD7+sU0MpguIfCJ1JsKr3gO6
bLeFRQCNk7WIuvkKfLvjAjkx/fPoZErIRHnX3fRmGmlDBlFbpvQZHsQCfy7yTu7E
nb5zI3OE8v6KA/ViYIHhHFMSLOTJvw4CN+sUugSWAMyqZ5qtZQmjo+DuZcpt4Sf3
uCi9aufFzE98KVxcOpFlY6c6kKbvYxuauCgdJ2uGDDEQBFtdDmRvUB37fhE9PePq
Yv7Y6hw/c7OQlGFrd/dajhpyT5JYlcG06rQI1wh3i1jEgWTTxTkTNXCfOZFKUGH9
ZpLMBLYWqCU3aYOi/GXGATfPK9StJKQUZdwI9LsnK2cdzTXlIUIJQZYt3ltpk0LD
usmjqtgZz43z7D5f4d6CRGjay4uoadJmpgzItcqNCZ/OjPDbJdLPDMpQBC5+OmAR
cNmPiECRl3T3Vww/6NQEGf1wjjaH+jUyJ3hM7ABvIYJYUqXR/VK22stxGziv+5PG
ntVQuUOje5wiQGSHNYVwM6GIKHAwhrI3YrwI8Ns3Bs2Eh1M/+V8I46E4jiAU2Fq1
aDo15NfOYhUOMX1r/lM448pXIr2Fze4229VkLLqd8ypTNNkm7L17gOKaKFCB9TCJ
AzcMC0Bn8JDhjB/STK7BKvzC4W2at9FJS4vmkWv2XtlnIMgSwKkWXIWrq0+A8lmd
+XOOjLlRbc0Tx0TJKGbQB/dKRlSD2ApFOocZft8sPeTKeG0o8+vSnzky6llE/qp2
2i7rA1HE0s2QB3WR59iblrRGz/VQcMY17DxaHUJptE+F7ddAm2+wXjqEgVdeObNx
qMOGDcoz0uSwWRVQvglcfiortpkvGQI+WSkCRMHBNKWfwBf1KlIdFBKqADlw3BLC
+qiqeYncpuN6RgxxYSFgNwVboaqpzpO3gJaXdRbGs7nmBst2yabrYZGjotF+q5iN
X+ORfPSMYuNdbucE7joK5+gSRF7yFUPEdk8Q25NXq/LH0suTSX8L2tze+A/8AkQu
rLjZOr2tqixSMRGq8rTE3g4M98DRUhuBiKtlbmFMjjehcQxpl/KSmwAIwFmq8VCY
JBzBPRJn76dtQ6F2QrZzqBItCdPNneJk6zI1n61d7PpqiDF7puSJXvYVu/nfMJ/g
/TyZ8nD9MwM3xGzDlNb6q7gcitN00GQVWya15YKHV1z+noSwmmq8JgNr8+1mbsjW
e9nB8sM3I8hm6XAFeDVfsQS34pPS81ANyLJmm7D99yuv47fHCfRo9iykOZNxuwLR
5Colh1R1A4VLOB3hT+2uUXF1jgbI3vLrvPviTArRDezoZEA81IYXFHdn8EHzVldd
zSQdkxHKohEbq/27ElrYKisU8AFWRYPPI+d3pOJzwqV1MYd6SoaKjhSkRiAyJ5Y9
AoPqTMMhRavpKYz0XOTPq7nRo31FqP7tGgO0SdDyFA5awTgvXqdPSDlVWApJ/yzj
jLUXZ17Q2WnsOOII8TEILgExrk5qYn5HJKYqcqlTf6XnYaxoU0m+NN04yQ5pit3P
HxuIQ9De48K07b0H5z7H7Xf+94ZUX+T6tZ1Gb9gyvi0HygNBckSxaWorXrxdnwQp
iZ5G5+MBFIjwxmNCTk9q8+ef6cGD4xnaSjZhtU7iZzhUBBkso1l96avjQqK/GgDx
yzEaDED8Xg9yenn6cGIGAD1X2OSCZF5ifj98wimZsLg5H+8q7ryiBLc4lkAnTIDR
+w1SQMJmMmOvCmMB42buJvlRZYvckTdOxPkVpM0UI5VWPiiUvQbjVvuyZNM1PSc/
X50sfId0TROep8JxqR8GQyGwEyenV1sMTvJ1b0WKEovkLnttFqKjEYvrYY1+19nM
ob/kMwsqoa+lgK3X/LK97RbYpxG9wLlUBYJYvJYNE7ddMb4ZFd+Yy6Dd8PHR/DBo
Ke3uldPrvhQAyFuiueMWhQZUDxrsChboh7KAicGFYajLVvzRYNNVfwWAK3T3ioGS
d293jD5h5E5ATI2llWEC57sbsEPYKRGqj177+hPKV1v0JVvQP5qKIdbCy2tu5C1r
W03tu0n65lR14VMAMNI3oaMpHQinLgyAYJOjn0HckEyUV0KDgrNdSMOO0UwOt4wO
SoZspRV0OPvjYBFw1TxNTVHGUBV41A4Ouq1CTXD0GZxHzOXzlYUu6b0grts6130i
MdLyAcWPoo7afaAtR7Er4R4oXaU957QLN0OMU7kiCiVxYQwv8m3JgrQq6FShc1LJ
Qsa+Qmfezy93RXFDDQqJic0B2rNOsR8FRKEsfAnQ/1kpb5Ajsr+DleNSu94qYGUU
6UJYgEwe7Z2RrPqEnsZYk3+zCGepwCsWxcKROJFwu3CdvyEfYjHOlojKoj9klq9F
IHo85xAkBcQfE9ViUT2Lcj/sYNyTirfsaWirbux4X/PM5rfXuvdVhCftdDFgFaM/
BokDWmNNEj+KVzGAAe/jYBPLhkz1NetMi6u5bYjH1IcbTJGrS+dThTjJqjFJZdAh
C4tyyDN26lR2se0xFadhh4EjWVwEm5g3l9jYuGXQ2JxEjvkPRpXkBVqzcvyYXBDy
TxZkjtfUKwkq1zaqCZZivPVtpxg2R03wk2yZcfqpLOAUQLioKHvRNmBXn5X2V4oS
xp+0e5F4vDI5DWbG4zi6munbkes9bNVYCwcyshZp3fQd5K143e/1ZTTvgbATioVK
9m+1QDc7uCLJCmOFIhciJfSf15zhx6gjMqmMKFM4f5ii8JMbfmnhh0Wm9Jm7PGHt
6tBKLuxR505LRrYCLbWjLJ2MSbMEhHFObwKkhCDXn8WHPwkYXhOJBOwrN0QZDqI8
dRdVYLrYwY+2Bhgw/WSBUOsts0YzdxylNiEfZZC5pCPh3dtWvmS+cNOw5PerwEAJ
AmEy5xUXlrXQ6J2pYKnfYdfNtjuIffHCYuXtIYLlcb4lpSdy4w8aUw9eHg26Degs
QJMoJK1t/fRpqKR28RcOYgscPkAe15Q0ScGm9r5EmfgXxy0jLM+xoU8NntpB8laR
9Se+w6StZ7y58jrZUWD7RYsfoa66d45+qm28hMTBvD0xWvTashvsFZTp0gJctKIL
v9wtTyGW0tywmrpAYgymuWtc1C9k9tDlpUEU5CPLRFaD7kZNrKRDJYJIvkduCJ5y
UxNeC7aiuuGb1MKggHq+v3eqck2134AXGAyxSyEn4+IGz2X3NiZT3DceTPlBXIRJ
agTyL0/LLc+Br+KYtcAU+6PNAnHUpHf92uJxjAY0OAGAZ3wg7R93bPA5kmAEtsk3
Ot3wIhZ+iYX9NDDGrfTlCp2MLGKe8GF90q6lt+d/se9BOt2L0fNW/IIzXqaju2w5
6YzZtfNfgQ3lkOVzXqMJ5Oivv4XUYrVAFGxlSVKRPTIcq7b5CyiJSeZoGmDx41VI
7bWdftRYh8zMUgAAgAaYl/9g2TjJnj2n/8TtbEpTvN0A3LESSdep057sWnv2OeG8
sXi3tB1N6I2HSK13DCSRjCTB9mf+H4wW9sm0mrgEoiQdzARMzSFx+tGo6A2sOpKo
BUm9DpDkmVy0OqM++POrXZulud+3H5LEuWWM/vmyEss80N/c0MvgXf9h+MyEh/zV
aX6hJAq4W+Fny4//0ZPHtr0Phyw+ybYa9Rllg7qMh0sOmVOFxg693aUPPYiPo9P5
/RngaPRc6fVkbc95UJVOk71emxDQz3BFU7OaVQ7S52DdOsONkkRUGmPG1htRWKuE
M1Bzgewotfup3K9ohe6e8FSQFIBtUFM9y3UtvSIejsOXgl6HvFj7Pj7JtbMQFsi0
1kxmnSw/cRkgmwLodl3+2qBkG6GkZcbKxU//2WEBILVLbnm9xREAelPEiCsEdXmY
sMfgD9ds1l4cGBGkBhVvuwJgE3gDhZM9UQDyzo7fVcDBWCD5ZABstdBZ0LU+m+fl
UJEqU7IEUq9MmYq8r9hjJSbafEtzsmErkZtsZaSX5/+E52r2cGl6n0BXpN1TYnw7
p4Xbje33DWA5Pmb6dmISxMjHkVfB0i5mvFrSWIWwT9cmGqKOocQYKcPEwQhvMijL
NdnwXiJr8Ncgc7LZkjZP/9svVsDDpjK7SnjDj86ho4OcWVnWsRh3Oz+97gIsVvFy
rl0KmYJgvNOrVjvEQNrxwm/T/0cf0A8GUzg1EKOspDJo5qg8ca9hEc6QfsPiNUz+
YFEysXcuJIB+84Fe+0qhsJaTTyih1Lu5FY+ewPXS5Ap3GWDD+SyCF94js+AAXk0+
WTCdq5BwIoaJlDGRHjgkjpm9bCEdlw6kEYPej4g5N/1D330qsC5dbfWFyNtB76LN
GvTHKsgbi5iTSZnmWQnT8E7GNFdDIk5bsTcEi/PTRW240bCLX2Ro+pK7kwUugAOD
sWzkzQJCVWxQlaHzRciTw8no8qfXwzA4CCJFlw8g8SeXWhNW9YqcZJjOdOHoRXa9
FPQbLXvwl1KICFaY97gwRD+deh0bezO3qZKSLv6L5ypQMAf+MUNCf62UbFUT2j7D
cSR+LfN5+KbVj6frokkwzCjBhSqmtK25kK+NbJeostzzb/YYusi4JQjk9npnjkSE
dN7R3GM75w0UisfI6v44by5vKzvKPKwvQaV6jtM+wsS18GJL6UoODZp17FINGtF1
kqC65/Or7CwCiW930S5+vNISMiDNlYQxMpFDX0U4LFd8uEyl5/50ZA7kCDFUJLuy
0wKF2Mf9HeuxIiCMFn98iWACAm5K5bOyYKVRxISkmT8y5hndrWWEuhf/9V4rPx7E
jatLJSX1ldJeKbB6mzsjic0pdmRN0Vnd5i+gC2qXP3j+nyGU3LHLqKo4djnoJEWM
DWpkCM1N7rfefmrN6Db4OYKxv1cgsN1fsdnNGBZheu1SDZK/evd94pN8fb0aPx3P
GArnRPqz2mDHxDS/NqNDrrzxWWgbGbB6sBlp6P0ik2v2XhUJ+1FsG3It8cnPO0Zi
2u6VkdFg4ODqXB8zBlKjm9AdwrrxlPclo1eCGh0DLW5Yb1/AM/EqjxHt5ZaRh1GX
1wdLEhJPlUJ2W06GisCMLKGwEKXS8xk/4wsjhHyiLX6I7WxjkzmMGwkUcIxe6U4H
A6oli6A7YI359TRxMYl4+HWSdfI6uuEbaqIX2JSHkwgKzr5HhXtxUjaLJp/JZCTA
76HSd/dDBp3a6wrAMH84Ws0o1ABHChMLvv98apuAalIswAt5R70QWhsUNM9MEqDJ
mho+Hrak5F5fzrryNxmMNJoiMlqCg6+Oi9PEYvlLxZfzVNiyoXhhNL7CsVNOVln5
9tLLb+v56ssQNESmO//nYeWGldSHIURR2nEajK1++ihZ1Dg+LAktkaJ8Ua2H/Bid
qrfCoKvCIbf7I71Syao1E4KmOHCQY0rTzIPsSNvs2WpHBEjd2rrjlMgYgQI024Bs
rU8qvB5m4GJDZpf8Iw+ycks2lBYCkOcDy5Fz7Fc21T8zbIpAP6C73ziSDvEgCCjN
7pVTNFGqXnWlMFVDtiqtkNfBbU2oNR7mthcWHIN8qubH0Pr6+eWHoy+a8KeBBd8N
qEqpaZTq7MKW49q3w66FxTluuQU9tbcs73/zSpSsPA2ewkNqRhH3SBpKg3MT14O3
6PdSMnehpgYduuSOkAzFqiVeyHPhYVT5Ut31rarach6VAQXJ6pELIQJGWOoJREiG
C4FQAV9RTZZB1JkRKgUe/nORP1O7569wFpHr/qX7FXFyttuFciCuVcecDm2/J6tH
GdDPa0SrV/CfLeDjtnl3Fyt7f25C41VChcCgSksKDG4MNwTZEzFu9mP88CCT2OOZ
gGW0s7bxhll+Rhzle7tVGRPqrtHe9ltk22obTr2OcP+hT7LrvlNUIJmhhHstFnjE
bLc7KLxPXpNgI86xfT8sIpkc8r+bZdQFHGp10GP97uK64NfjRkLH0TmhYoUVXl8i
+UqOCssLuR61pBjxFVEHA5gpd2WEUr0HOw+anCEDll0DU6nSR9RkP5oaWNj876jI
OHZ9DBU+mLGDB8OSHH9kJsIbw35tzcPM7f4Qp2SfDIzzkDluf0CmzR9tTaCnVy3u
divf7+fXDjfuEcaDsCswD3LLRVv0NMDDjTgR8+93pntd8WSSe4tgMs35oMrp8qes
Xn8f3A+CF89AxuSPoXhUszmHqBRqc7IkQ6wIlMqkWKOJVB+6vyhMNM76UHHySlYg
K859hAggnnjLnTTeyko4kzdj5wKPK7vW3LoQ6IsUCffA8+mfmpIfpRPzAJtcq70a
joeui94hkCw+MuMxA4bBaSpo6gKyzkNLHhLW/sChyKYlphG0VWMd3ILxi2RFDrvx
J0g+A6AThogYZB1OtuhjefKux5yFnOXDKA0dM2DdQTll42F1KPnZ6729k2n43obp
T2v9qyFr7ElhwqqE0lWp/MR+upEg6lbJ1Mq+fMz8C9PMa3iakqy6SBOMV4o5M3tP
V4e/pDnwvDqxyd8mAIfn3sTJcyKsEaExFVYF3ENvQJd+HbPt/Cbyk+/NI2kPCL4P
7oExjWAOG4qwUKxLMa3ev+j0md8Glxd1aLgsowhzfYKkNCW89ys2jmcs/mFzbCSh
WMJ/W+zryenBiuKkz6Wd6jNeSQWyhmgT9uhEu+TwyA2PkVv3nXXyT7DXSIPnxdsE
5Ewd7S+sAFa+HQ3RTDOD3CEFtnwm2WGENQmPXgcsTy3SjbR7/pEBOGeeto1oNXcf
a1ogLzE18822/UcB0Y0Y9Z3SH4exTq2dufUPEZlP/0bAWiYtj39UNg+k7AJo6d+0
AqwjZVWhJBItqFR7FH5CeF0hKSk5qR/IRNglcOHk0gp+lzXgH3SUY85eWDAjGuHL
LlXQIamtNRJPiCFXRbKS8a/opVpUNO3uYjUavdH9Scer3+QLH3e6kt/DL/e48USi
fbLM3oRL/NBpmRyqaqzb3rIxR383kQGb+S9m6HcdOxhcdcsBqjmcun7yVFE8ddbP
9rSTlMSn67APKVPmzgI50ls4ATpgN6FWHN3dgEbK3raj4mP65ei6cdtki56Te6j7
DbXNrPNZ3ph3Wdj4a8+j6qsQU17bEzcm+vkYeEPFFi+1jcfQbqFULIxLV7Co2DqH
5s63vxloP5uHcAzI68jDZQaSBCSe0Urn1ia6bqNCJ8JIWcc0jTmeyacn4bBp9gAw
UE3LgV8JGclXmP3DUvfJOM2JzPgJz479kTIDLlBxbsxbB7e6YikXM3N49n1joeV5
8bFYTkIMBHMEO4y0uyBaK1ET0nCah/3HjPpxnfZCj8ZaouMRG6RCWYyFUM2bkfBM
yM8idS0QtDxVr4OmMMdkCh5683t4VvD3Q9X3RzwV/5pNVY85XnZvwYnEoDQNQONy
/09+os1GgyqijRuHg62QQLRtgk9F/TuxGK/vQ4WL5bY7kGnxbdRQcHzGn+AyFE1K
H2i5Okutqf1MJHmVdcG1uV7rthR1/jbpwCm+vMcIL+LnmeUFQGxdzeyNiofbaTc4
alz17EMB/xddNuBiNHJQUMVYfX28+N4vvP+nPAS73WOxI0cA5eiyVdFxhoCc3QRE
Uoc10gDb7kjpLZIPt6sfeBKD4opK19a0CaOHQkmVq001EreR+CRvTslx1BvN1Wyf
psYkSyBG9zwlOfA8On9bxNw+joo3RsMT4+0viDdVR4/4xsGXOuOHiBT3pyzEj6Al
b+lT2B+O3tmlGdCPmkMVqdB7hvdzmX7UFUC44CR6MWUTA5d4kaDg0sVPzjrynHJp
CyI1tmkJdwDuXooeCBCiq77jAF9WI/TZ0I80syTe2GroAfq3traAYAFdlNF+OglV
iTi+X+s1Y1CCkLivGZqDzsHR9ZFfgML3rsD+eeiKlNU0nI0o6yY5EYNeS7dilO/v
CVJvJMbi2KtZd+QNFlzGCXzxg1kIJkAfD2J1U5wj1UiA+IUGWsQNAoPWZtW+jEfX
ftFoC2NHQ2QkJQM3FppN5RikYHJLiBsHc3caeFHJQQONFukXxhhykDsdr+I7like
1e1b4BScpuM9LtrMIHDfVkjJftQNtqf3ebTawRdGUT8dtOKu7u2b/ZgBOFeKCl6o
FNR/yE8PEeKp/sUxKMZiYWbKCRotOCmvvdeFuOqfiOF/rRKXvk2AlP0TjrE/rx2E
TP+Rjj5+2TJX1zrbKUliyHODL5xTqbdZf15DUQfBOnM33l+FG3DHF4wC16YfuVGa
p6Ypxuh0R4HYlJcuBHmAK+T1BKsRCAGbYa7clvBcxy40IbP+hlXed4S51TXhPX+L
kmaUGk4lC0bLpTjOu0+vqna5Zi2GrT3AqjTJD/sIiAWlngrkGtY10bgJCGNnKN9/
npNRBSYMGGQZ6IThe+czo+WfSgvsHoKWnm+sqvdjsRSHi4iF8IObnrA18JREsY1t
WHLeszxO1x3db9kmCDoKM44tJ4sEm6s2FpLHyJ9w5qL5jzAgWXxqciDOCsreBAXl
4LmJoAsUo2lVybYgSA9Lhjga8Zh9nKo5fnxOmKMBU2yJGV4y5Sf+78LDVFfhtR3y
oh9hhfcIeFSohiCUgxrnVWatxHhM+J8tfqdzNdcT4F8UuXGxr6OyrQEoVVPwnIGp
GV5N/Ba3D3D5IotaIgqwpHxtGOqDUqRNgOHKSw1jnKLh1jB4Jif5V0jVNkKPcQrD
/eR3Q9DX7c091pSys3zhcmS1odZGpW30HUS3rOEvZ2k0+I/vEymFXR287FmiOFUK
mygVpeZsxpda7dGnSv8/HL9uX2iYxhcyf8I9tW2wnP1gL83WcS6O4Y7R+z0iDolE
k4xzRpE92/KGAjkGHq071dHb2+VSsIvvzKJYcQnbDw+UTGpZbSv+A8nvqbG3qUHo
XDTK160wkdC1Ivq9rldLuwFIIu7CBTwXTbVeUoQxxNbm/QJy4/MziNCw8nXOe/W9
9x83uiwdQJLZMaiRQrGS1nQGfDkep53NVQ3t3Ui91ATrTe/NmbdMSA6Wbne38IaV
WVpVuuqNS2PCY3NfYoRY+VBD2HagOZLnuwS+RjtSce43mXpR5iLpwjOSIXE87qaN
IexMCu7s+J5Y7+pW+hoplU0rAAekHkRdplrvCDnDZdo9FngUBdIYtHHOl1Q3Wh+D
RDeqyqkQucd7O8mfuFCc89cfsnYDLz0dAr3k67OfUTCvnRtC6HV4Tp7NWYGQ+PQj
OF95TsFQM1m83VmHwhLY9rBrfVbVqyKvn7gyfafEEoD6bncW6WHOf6kVUtRP+ytN
58sOTw+TNNCn5mMM8GzpJpynKiqXvLwOYmDaqyGdPXFeKAog8V1V6clJY6Ex5bxc
53XeeCoRXSLqh+Wq4NMpYY9mT4yEQPe29valOXalq/Rl9U5HpjKzNZXkWs/fx8/j
K3OvuNcRzio3T+j74N9d1qrs96DgJJxNNtJHy4FWPgctSige7lwtDnm1N9xNKiWd
PZORJQ+mXAA3JlmmuvaJYwRTsGf8WpD5kod7SrlnSI2QwYpxi7cKVZnT/E0b/XGB
LMg7h+ITBl2h3YoE+WYMS3AwsZRFaIklnsW5yAozB+CNRIcnL+MEx3l38ziO26pX
1y0L0lUehCM2EHb+CA8W1GXHi/FOa5A4xWIbtQjcrpAm15F+gLjO/q/dqh7rFnPa
5mayyNgrcLwV4sgy0jad7APU/VdwmYR7UT52GFAXwk5DRW8rhssSnhS09dchp6d9
jSCizvVxw5t+wdgqLcPT4NjFMRq5Nn/mewqrC9KyrC0/SoLfhWWIj/1K38o+EkVA
9LCV9ikrFAlgq3D7zj+L199H51p5JCPlgzWSk0MWec8H93uERIDWgWy9xbwGFEYr
eUzGqN32Co4F1OYhWlbhe0RtY/MxwRNdZKW/Yv/mRQoQeCAqzfoTl++piBZ9XEbq
g+ta6p6xOee4oo2O0okyuCh82I9/0tKMIp+NJ/Ehi5WiZ+9TZWv60T4oA+ZEeJuE
59e7oC1cVTCOCvsByTxlijUkqGcEutXjuGomi8lKg4+UsJMZOYK3qp9cFEy8Tsrh
VYSugZhqWJKuMwlrHO75zCf+0p02fDUtLuy60Z8Djv0rTRWIt6GcnHHcVoqw7UNR
3QMSXGx4rJtOk6oLGyRRfyqvjTp0vThTe4gz2nSaAmU1FO7Rq20vsm2Gb24d6ohN
U1JAprvqh0Dw8fOxxeNpELXwnN4GmInS/WWMfXllBYVIrZdLWAQIrjUSrXGdiyBO
G70XuUKCNkMBz9xo80kKxuvsfy+vrA1U6xVkg99fcD4Af+7HKZKlAoAMsmBcR3LE
Qe+QOUEHEVrOMZRdu50IB+RTMISo/kllu4DlMcSHzxLSE0JPQErGkXAAk4yo3dJo
HQdVCB8LFBPvCEgS8A5dt5YIVNNeqV18b90ZplsanDQk6y3C2sP1iIuO9Gd3aBgR
HXy0x5ZPB4EPI7Tx4ykrHnBZWQu2TXPaE7ln9OrREKKwMsmqBBo7fIWDi3ZfwkCu
5NpcbXmqNMfc9z4LLqYvzh9CXYJ2bhDYjj1ro9kUtxh2DpHyHesEig1a1A9ZDDJC
Tbk9OjLIvuMjlq+8MpOdGH4/xZgeqk750jqqWNr7FFRADIJi+mj6BLDJvzDEPvv/
4V982VaB+2cOqKOJpn7YsrnPMsaoIzytTkqq24pvaAazBTSLzzveakQj+MwZTjh5
h/eTi3OzPfw7ufZ64g+FYcgYZuSHOACOTYpsXFMezYyUI0eUwTin8eS4iWcN86F6
tXui7GWAW7TFTEX0Zi3yybmA1m/XQA6NAw5JfyUoYzn8ndK9mNtDpEiUeeINE5D6
DVAMxwLk59XxXfzuhIq2cZYlf6Ib3gshE2z5RvP7dswcbB5u6qAaBccE+sgqT27J
iJtHJUr9NrPxTKnmOMeIEZUlywn3Pwkubi1pRzgX5OqeftIt2fkWmJQWEq0Oi3TN
tKTXlTHvo78iqkDScWoIfVBuNm+D8+epG44CX7sA4G1Q6eW2dQFtS40wSEDGQ5vj
whRTclVjeUS3ANBBsrH96DQfhOw1WK3HQafd8o+glpPzPcPjMAngreq4Mo8q+fYF
yDMAB4YOhxhkndffVl4ll1hsDsKqAYc4Ojq0TERjt4E9lWpRowTdCg64oFOZuIru
m8oxGqf7I4XFrvKemXkvJNFNOByN0gWWsWyCTV2zIxT7ojQ+JVQVbfYQvF2thDek
F6Dpyw93bEtR9NYqvRnzUvjl2GihBWItbDWS/VawpLHXm/YfV6jj9jikf5PTNV4V
buvBVA0GvAoiL1i+RXmv81AHsWeKpfOWoWgOld2ItMzh9iRirLDr3gS+Luy38O36
HfJe9WykEwBH2Dt4Batr9qvEyDayMK+Vxz5nxwxXJGwtPx6o+PaQvG1i9CahyQyl
DCJuX8FogUrZEhNfmQPXOhLLCCcF6m8zchZ57EdwoSxx5Rk0Tb4QWKs+Y2vMvp8T
8tTCRQOQLbW3LHy5//o78moxOU/8ghyxJM17unQYsooQ4yExZ8Zq40vjvxCVuaIv
90sGB1wGmoevS5AMK2eePE8M2gm4oEtJVjmgAAVSiDPxHCwGTPqzmfJx2ORc/YJj
Uq9vXRnEEBhaTDSjUZU5Ayg9YDxXGESa4fl6JzvVu0lwKyFFXR1EPQH4XJ0aLb+2
Ls0EvsEKPcN/8C8WUykq3yW6O+K0XVewnnO7S7jKSqu+xcovqMRXjme9Pb58uY+u
jL1xtlzBQjyREf4OaMu1SkOc8XxQVsYQwJ8eGXVt9alwkImisYh8dokpQiX8VAEf
QnePeBvfqJuOlHlaus/RLYFEiJt13Us7+81cKGLEGyvG51xzFkrqd+KZvP1kcdj4
Xw6WOrQwe+CvfJxniLb3KORnyllTTaDx0IDSiO64HUGyFrw7VUP4/N/gO4Ia33/V
maa89g/5GFIXNvjELGIWogGXkO+WFT6x3TPStJXqsBSX5a0L4KglXX+I8gx4mzj+
PxAgKL9aH+3ZnL/OADR+JGSgn5foqPSRTUd2ktXVdhZKA6YKvrJTdzcIGvh198st
Ag+LKP/knOdcPPxWQ13AejH74mc22ScX06n8mkvQQDNR3wSTkuv2vwc2SXEN6aRs
Cclm1NgB+SP83kHYB6zOtUE1F+/rKz88OOEshNQ3/eM2H+xdkjC5VZTVlbu5aSNj
5FQHcXcPdSqKm68zUtp5jd3Salm7iLhQAz6p2QdOG84CXg5uvIgd+vNveqymygF4
02O6q30zy8TER8P0sjUHWQ7VRoLq9SjmItjs7dL4y8ywuN2HiuiANC/ahych6oKI
VWp8qYpbAPHekpkdYPiT0aUvaZLy6y5U07sOlqwHCcCM1de3w9XlNU1VvBDdeLb4
rDCMWEE8qaDCGsziOygItW9KQm02yk3HEpUuFtNR5pF4Yvon15WZF5T1WjpQfT6k
A0VslCJ+MAGsF7adbmgtPb6BhL6XCBj5Tk6alIYETRexPJQqTnLC+aqd/s/ewjjU
zIB3Xx4fM4Vr9FXtEyLI5GVsr6y00TK8bpto8Bj5FWnPGpnGF/fLjKwkFswd7r/O
t0QAzGIZD0vFK5Tjdm+Rmj/33l0hMsUucZs8LwI+kwUoIzz3Ur1a1tkKwYTPwT1G
lHv8GBjI9Maw4NhfTnV8wXBkFzik5Pa5qwudhV4GoMm/cP/lnkg/bvUlP655EZRo
pZRZm3lIrjCU3C/0dtIMaC8p/nPe36RDAW3gcpzvwnJgc3psiAmveYWappjtb1Wr
ng3tym6i+XwbNH3dJ3qMw24wlF2vcDbMP69IqayWuXY4QJoSPVlBxsi5WdPcMKNj
cHpbTRmRSVU9hU8sGRYw+I0+ghRufn0CFGn1AVziXye3K150gnBeTXKDqn4pw+IH
TsDBApDBpgfzZVhfziEzQr4lJ7P3t2/npP0DSigw5B7pHJxOn156cOr+ozuHARuU
jC6wbLpWUThBUTgEjBft7a7CbLY0zetgFnBmi5P+7Qb4KRMF1D7fPBzNtIQqLjKj
Jrd5YsFxwQI0+H06YK2WzuP2pOCcjjRPoYDL9ffanaXjQTFdLkPtlTDS97ss9lDM
Ge8yiDnvUoovd3/0auzQLx60P2EcovA/gYz1u2I7lIcSlg1lGkmRde8ftJyu/OOD
0dK3wXBc23mvHCr5oeKjFG6wmI7EDEv2Tppy41HAsHtWldyLArtzBQMaVKYX/M58
YfuUV55mDEPIdwHCKqjHK1Qo7h64dUu+Y/YwiosHLn1grEVVdHJqGn15qNigd9Nn
FTLbz1jlA+RgL2HcK0bTDj3aEE4Ioa9NddYZpj0X+XoRerHzWOXo2JgxA9t+PbHK
cdDqOwJO86LTlp3VJ0fixdNfTulyhT7LtowrZSUZ93hUOMctQFZvYqU0RvDrliYc
JTVSB2b1KVcRyKQI1aTIT7fhtKjsl2YPn95ZLFLImrY/xv2OWU5LCgkhK5DRRWnV
TGtJPIC8BVFFSVHVVZZYNL4kaZvdF7AemlAEY+7LEDLEnNOneBEtX8C2FQ+nhhIj
Y73ul2MT27EIl924K8yOTwmTAzeuNaMDn/zPZB3+XhljzYoKu4j7Nin3NmraEsUj
EsagJU8P4+epDgqQXR+VcYPv771G72u9loJeYXPr8FHsQpULJBl+PsawhZk+SUF2
OGhRnMt+yb39XVB+DLe3h6Cf7cS073e80V8x7SDwwU4oe7HuccHtABNMRWffLzT4
hDQ5mMK7dtteFq7hRe1wql7cP5ycvqkZfjDuresJ6N4PD2i6ooYLuOMH7WAfCck2
odG6r7S1+2wMQgUeDrOAP6uUIugwJBxNaWy8ilVEP7OYZm0AClN4vLeyk6/LmXxh
pgoqycSPgvD9yrPqmqCoEPAnI4Vu/xWnnzwfTKHZjAiu9TTx7GI1R5Y6n0lbc3Gt
KpK6ckLWWj/eJCAe+7CsApzm7NAY/IrTKQVl/frfaVZW5bzP70IJejPvInlPskhw
K8ZsZKyyK3y3y3wyT1BZATum7A8OzsGchgyS0qT8Ctsv5aQMjqEeJlwme7YRR4w6
nPZyhP+XycanmqWKTobuhD46Q7M8C4th2zgWaxU0h3kjM1zXBr8Oh0oCE4FDKha4
d2u6y3bvQx/84RmxfrpN2KSaVMvcsvLK7HUZNpoOhF1f67LNXkpaAMekv+KixXcv
ie9a9BuBS3EYDy46IxJ53fQYrzPudkeu/ku7qYe0/30STuJRuKjv1/9vuRCr/AKo
rbwqIq+mD33gfE1v/ZP/AnefSW/eQ3Ssg18m5MSf8flzZWnshEBYb/iTh0Mjv4x1
rlRli8nWB7iLtuugvBF1+PxOpvlRJnxEAWpBjbzIgGNqC9cWJNvGUenVO7+Ye8aq
MWWFvgLQKNim6epXBebgUqoiWFEFgj/BtFspJ3cQGu6/qb/YN7sIe1pprZNppjZu
lOGZ3zbsSJZ7mKTRs6YOCnoQNR2bsf30RwKyWrenMz6/zLt77UgMd6G6Ed/Mu7Aw
g6zYourZkAgu8DVzAuhYMzZhzSsMPirDq7moWaf/UKBybh1tsYVXTVczRiNqXWau
dj04lZGVfrYa1tBosDY/19LNjQboyjpoImdKeZMsCGTSDr+dEnmLfsZrJz3hnMx8
69GV3wNeah2Yj2Uvz75ICRq/XmdnQ2xiAEQnQBxglTqVzoPII0N8gOzAJ/OFRX7m
gF8BjrIy2tAHRbeK/7QugoDSD9aC9ZwUOB8ZZLoYu9Z8tPFzv2DLUj0Ehh265q2R
BRbEjpBxD19Jk9F2MfUqHy/9zAmMmXFJfvk3M5lW5bi+l+NbcveOjnTCm3Ay8GAL
WRn8tndGjTWGDhA5NM/oFblf9+ie+ac1ICQNWFg3r1yruvUycl1E1G36jqYO9h1E
OrkfI4KHgiRMlQqbygKYKNLNYwTy/Ye9Flo+JuAWFtIOtmdgVEapC6FnAloyxwBO
kPZOVR+Garm1zNFKVUE75GFhqXyJxeAE/gbJTtsR1oUfB31XuzQxHHEyazUJrhCK
q/In3IAKvrtuBE7AP1jBVSfFFvLkuCN0AGZmGpQD78bbQ1/ggDiPIjDSnTEfpR2Q
5dQ4ciMb4K89DrFNfYuhSbe6KP+V+QRSKNM/0v6+2GLNwDCKKULvpTJAqKlUmeWx
RYj/5WVeM4Qfl9t8WLSxXt0iBeCFuXrFBLkY2tZrs5GrN2/CnNYaIQup/Nsywrcr
1c7zOVk8K8f6TJNUObu9U0PXulZCsBkJwAX2xQ6H6+WffHPP1Vm8SbxUf7zc6R6K
VFrgPgBPUb+zGj7c2jB+ZCK+OxwuFQ3iDqoppPuOsVuaf0D4joFwXZZuh+1l4F/m
I+oFiylI3iPQ1sVNfXZ9/PQse5Xn0IqeWqODRz0t/aFNgyAHUlgteromxqf0DyoX
xROS4SnkNQSpFVVtu2m/vuwPqfnkHrHOUX7ocWitpdS+Eqwd85gQZ30K8iGnMmgP
9yxLJgI2s1vocb9sNPIlC66em8brbo0Pt9dEdFJNJ8On+isnYEcUyI+YNd5SkAOF
yXdIZWXa3ovpFueLpyZ2V7x7Yn0q80zHp2Az1aORyAa4yX8/QHyXsF0auomy2WDB
W5RqSMm2OJVInD+PlV6FqL3q55HHIPp+IcGEscq4qy36XWZg2Tj5N2iYyVxJa32v
6XM/xUZZqMHH1kj3jBx6JmRG8Oy67JW7ALhEqpeOvXYHQVA2icBf0Jy4sgfLzKk+
SS5CT6pr47IdqjaADZFTu9x32Dsrw2yZp3FqyOh+q6pVZWWX6HJb6bdlsVEdZEe0
LR+gh9zfsXmmeMtLgF4fIrSivVG6M9OQT0SPIUQgF4Foehhge/mNX8Dzjeh6wCM8
o944lrwLfEvXP2asBB6avFjHbJug4YmMRa0jOWuNbOocHq2B5cQ+oqxnSisRyt5a
HIYXUPccG576u71kCzTy8G38Q5DdfKRKEAVzS0HajLolTEKxGX1EXr+8RKzgnFzq
jGcrd+nw8IlRyC0Z7t2e5UWbM0MX6pLYnxw/djNnWppXLzG+IloHOJaICLAValNc
88rg7MUF0XTQQLtX2gWeTOhiX2HkbEF99rFPw9b1Q/Oi0F1/DrkfezAXJHlp1C3N
O6ghPq9tq7ppgfGEs2eE3w20P7eI90+bwaro/BEEzMU7nt0acBATU9y0Sr7dM3o3
5CTpTJ69gteZyGV5LVvuhp0umx4SC9hPmo9YAZt+WZcuKxtQaQN4Sz6sezWjgaZ7
KCKuHRHkcAQHJKFFmFsxREgaleT3R6ZeoIuwaTzyM2/0oyv61kfb3Glfd7MCn1ZR
hKviUFoHcFHuZUwEDhEZ6i0MyXVEhRBXpMb/Y8Onf9AxzSJSZ9NR/U7+hRwiJwQy
bhrxlotwAskDseUkCQLdU+JgJG/QxvcHqI7MeDap2Jyo44zJpZs9fOds++Sf9pFz
1jrtx9amwmgPLZSy5DvMakEH01jB9GfkiHASDI9mkN7xskJjOjI7pwGqKjkrr3Tp
ydsjjSzM0BALYuSH7OJWloepOhbi4GyVFUgA3LsMZXkZuY5f5l5vzR0PG3SgTYMj
kMR6kSVhUmuAeFAZOgSlC8WqgM6fXDqM7dZHkEdUWwNSDQ0MZ820CdOFlpCuihBi
aZ4VSkHyMspwinHDDAQdoaJDq5n7cdNG10Vc6WiPMsnxmMrRQB07O1Ks8eR7xchC
UJZ9cNEvEe0CBQ0SQdEXz4wc4x43yuBfznWXD095jY7jedSRPFUuZYagBSUlTtyW
XyEMABGwoI4sc80mfxYwp07c7RTuPGynkwoJoeIZf7uXWmHiS2TFdwDpDSJRH/1q
MfZRLd8+zZON4EVaqV2eVzJ/ZWomHB2a3N5xfwaqHzkr67T7WtiMjBBVFiJS8cwV
+GtcY0HB/55Onu/piLgUAALycDRuk99pl93qfV81eJgXH4D1VQRbhd56jn0gYod7
OsZPputzzwuGe0p1xP9+aXoBTvD2vII0EUTRkrrqq5FjLMaaukWwfJXZTOjl/abW
/YzTqR2vvDIO0UKl+8lKx5MunuPQN9vYzyFyoMUJu0yIm5Er+yvdRInXLp4CXOfN
6rL6QIZbM4YC0zClAaxor78XYpFH/KD0vYxhvd9JtXu6STwZYOWjGPpGOeEh7pdt
AMvMFUV16jREyZ9C7lT6EVeN/3G5wP5o5W12Mh9BKrFUluhItWl/tqPyGRvpi7hf
mrYZoaI3Z5XrRMcNqAfOiyQNhkp5xf9cFE/SbR8aMtzgozjaDaL3A++OxN8+aepM
KLnRk6Yigw/7binUZy19PaGl8Fvi3t3bxAwvB1awgPzgYYA6Hgg3A2m/flIK4Ryn
AOPcZZ3imoDSm7aKSP70mHZXtZzXRSJwim7ZVwbQikmu3AwKVFTUbSKosAygNPC/
ek5SmtvZmRJK7om/zaCt8fO+JVlIi4he5WGOoaig1qqZav/AHVX+Tz7mAxRjER/h
uJFVQRS5VYeK38Gg8MzSoKf1ZO4TXRB1rm6rgoh1YlYVKzRFLniXl/BMCa98aV4J
Sh8iL2NP3WML73Ohpye8jBpl7CaD5MAsgsSJ+WrywHDgw0C8LSv72taPmBBtdF0S
ehkjvt/CwuGPlvwsXLOcW+FzybvPbSsr0VOzBKrI1PHRlMDW0xPvGZPw8exGoxnA
awpo/dc3mpHF2F6UfvSJUlr88lnC8xHGwc+4bV+97WwIKmh6H7TiZ3tOgOY6wkaV
tHqj5vYv4BsKQN2FUazvFL/SSRNAWd6zjl6YihMusxi7ZdjayUtwet12tPVHKsxi
21vHAE3YfSVgmd5DrwqcCq4QU7KWGkkR8j36VsZHgsQO0Zjs0Q/YrQb26gFu2JCO
7dRhAqskXUwpGmj7t/8R9jdFDWLq2cAt3RIHTBn+37MNk+7A4W9QOYsGd/N68SBe
eFHTIsWSjRLgMXOyOqFCYI3zRJoBJd/tENT7ou9CWQansVeLC5ywgHaJfTyRh5lr
uco5DgvU12MzMsiRGykXTRDTswh0YPTsw4bYD9IFl9yjSa5MGlvCN5xDCwsWE0Qf
RU/b9tyNUa0PZqvWMytXBWPnBEbhXyCLZng1KRS6MieJEdibW6arz/6Gnj1J9hm2
IGktEEmFoPYHX8veY/YTkicG/OgEyDf3ScGOV1l2I4lknHSVULDtoKp/F1OyimhE
Ae8u8D0UPkIMKnWBr0TNzzWpol5Uc+59UxWJAWnSBzGML1fyVZy1KjBWFl5vrv7Y
VpmySF42AqS3Eg+2FxJEtEyRkPIpjbyCA+bXpe4vJMgqpLgVlbVLlFdpJgWgwWXZ
GABfQxKdlnajmZ28lj2a6b6hwGqcwXR7lI7pg46/f7v4dzSmUL8G9ScKm1AXRaOQ
C0EfTU7+HK43PribmF3lUTKJw3kLE5HElKYP2gBA0CImXt3xEYBbbNP9D+HTxXkn
ucclEAgNN8EdU1sSOmPm9X0AWycSqdbtmviSHZb+BO4t34j9pd8S3Dvnl30103+X
cL39BPW2IuCN2KhbXNTdnsHGvmjw20tgTTlZl3iXTJWMt7e7uKYOSSq8Jtr68Aae
gK+S4/OG1ETZX56ihEI5lBca+5sTaKl3hqtGB9z9bO/OMbxOzSBDkFded6tOp+1Y
F4uRHk2VvFRai8vCeBnEIsu7Kpps/16+nkx2ttVcxHZGERZ4callwwF146feAtso
l+vKCG1FHTTZp025Y4l16tEKZWQNpKtxEAHmSt3aF5j4RSsMDj4CyQAIB+9kbdco
GGEbW/M0R/hrt3/i22yAY00t2iYLQ7NUJmcaEeg7ozxljMU4srLUz4xAJ/jPjU1s
QmqQXZu5SUUbzmbYk1GXCsf5GoNIXjQfxDKCNRW+5kfUsFkqiJaKPzBGyJV+GMBh
auhe5e5BNkqLdmB4T8924k9c9//8dDka/tLdlMBYKqI9/YNZmpRT/CF3h8ZgkIm3
N0tnI8bdpZxpsKqX4jcGTJj29vezQAD8adokIjLW5HSkfqbxV1Hr7t0hu5dc18cu
boK5lX/jnvltyEIBRd9MytRaV1uUsZ7RH3osIYRn427qbrqV5hM3NFBnOQR1ohCa
R8hdIBW/Yy5Rk2SXLgQVeFzj3FVuHaTeX3pEj0eyiZ98yqqADy6vY62pu+a1lLIl
ZvoCbi6FVAUrczotwE2OJ87A4otfvwnSw07FShsYP/huuUeStKgmj9DAMdD2PrjY
SY98e86ViH4xueS33JmIxni2YBotqcbdQsoaHwQb3S9pDrZl120Yem2sUbUn+fHe
CBch7ofx6kjgd/1hE11wqT7MKhQgVoCTyZmRSyA+Wv78gK2cv0F9HTHUu7BifzUG
xMhEQtp3nvm8cDEaAA+0rOrKa/WCfR1+5x5VzE2fI+E4Mhoe7nswYj6vyDONWaC+
BgItEk2KG0CzEKCZG2VOO6GNukwrSH66EkyckktC8ynkwqaqzLJ/EVn65sC7XsqV
AQrCYNw6wYxHBMm3gJw695tkpAr8T8H+Zw3JIL66JXSED+YDDQCp7eM9HRqBu/sw
ML0mrW+Y2WXlR6BdBMMEhZp2Xb/2LuB1rNVX6ypWJxItBJ7kk42DXt6lDfKs9TWN
Gh+OX0dWoSg6OErwKIhvMdTTamEKORP/0hGlkU4BrbOtJn17H5Jjs+F2IP5+pPpW
mNWmyHOvwk5PwylP+u1xvAf78HPiL1l4UPcuAgL17VZIGuvSgjAbZx0GjNQcC5Sg
heR95RsfOL4WVk5Ss9Iw/Nmxz3aKZWlW2j5dQBWwxeYhU1FqukN2jM5wkq+60ul+
3F3VUj9gxmRrSKm1TIoTEvE8U3fAeNkg1h3f9nxD2qoVXqiOsMovKuLvAcLvOkMx
M0t4MFq0dHfLDxwe1JmFHcQhlNtSGosNAuAoPIRd6aBY/bAlOfqQMqKN16jVmZOG
DDT+liYmqb6FxwxIrIF6w6X9PMubFEbljIktqkAaw9bXuvaWODuLUf29oxhnRGP7
H1JV1yMLSw8LEK/syYpB++zChNbhFKwgUEDMC8SAOjFNZH/Novpea66fZMgeY2E3
WjLiwKVQx1jIYASoow3Ym2St/S7zzh9ki6KAopj2M0KpahHYZOElkUxLLM6ft3Ta
shl0+b3SyeVZ5I4c88T56LhTshxUINhRLewmdPoaljcQ4S9oHQDywnabEjtBYSSg
k1DL5gmU0ptUXmixuIR7hC5duYFSvZ2aMVj4rgs7bsHPh7i0fsVYExI7iqZfjLRM
vphly4jq98BFOepr8NQUoMIiuskvDr/ufEHCNciDUMc8ChvNyMSTM/z0E9nlzgvB
8vDHFdJz35UiyguFrzYFpgu1MLG5SYpO3631yHyKvYbrfY5fW7TKQGkSWUjtBrP9
P7bYjp+IN1uoTlEsFn3DkKuG5dXqYcBRiMc+HxtVISpAovs4JTWnWgBvY0OX8rXI
+DpWCbeP5D1po9OUr3LHzBrtYoC3pQ4V1ixvWSHNj6MAivwfJX1ZaTLrtoe6rQhF
EPMcVGbwJ0guFgZ+ZcXm03cl1x1I2CRv/v7vSQLbG7kvOLwmDL0C2thdZMrqN51R
JJqImgcCxRNvBrIRcUSqsiUeFmDIgEIc++D1UVqugiS8VMBPmV5chJj5FzaQhQdN
Pef3oOX+9SV8n/nAYVE1lPo5z1pV3iVOPCNW3UCKfNIUgQlXmNEZnYt/2y0mXUw6
u4+/J45IndvYEFE8ZLtP5tZ8etqrIeM9JW38L2+zWUfa5/6A/SfLpAlLUAEOToNc
VGPFSoXCK+uOnE9hsB/IgSMhVax4W5NdyhXou08hru4KXpHr3wYoQ0YPc+nzTXTa
UlbZDjc8gviaIjBIaykof83ONsMLIlGlvVg1Rzz5NQ4wlkRf+C0sy8I8ribgAeba
5iniZ1dxI5Hpf+pxROG0dfQDLQFNlWOrSwZ3VJn9YuivJ3RuCC3oRGKrFA1kjEtf
KQ+ot61VJTe5SzubiR38M7wM+N2MHOPm2bitN270KR0oSKOX9Qr1ZZacHHAxo3TV
GpGxTLfgtDd5KIcMoHf1aBqGO/Od/mWPhM45rFZ2Cwluu9TkpdlxSMKO/pd2Jmot
hz4ISSe2O4KKzE5ofbGQZH/qKzCfxC5eynmmL7wWRbfdpL88Wkcq68geET4o0yTD
YGXBkWosFAt/EHqvc+ks72V2xePOS1Ig8YOUAG9zH5y/S28y2LxY4lwAoZNGFNRC
jLen5rpSkW5PL4KXLfN1fuUEM095SsRiVXB3EiFAvuR+lJmdowIKpMoLM4zqJNkD
/0zF1uR4HQPPkiLH/+gVbS3NbZOQGQXz8ZBp+bag79m8YBLeDPq/LyrD4YEtQ4py
P+KEQc/qSeJKrAqSYkNuUntpKFsBrEO33rsKb8uUGE9nKiQqo/6Yko0r04dhto/g
Hbp1xr92+XymtuNHOk6Id2Qge6+SSFibPjsmsEijRAIfDZb/+n5dFqScQTZlqOsP
EHZxsmn9xkWk68KiSUk9BR1j/vmbj3L2jKToMpnkhjlfmfRJAZ9lVLib23z9NVBe
CDpq6xhnxIGnWwxGr/GfF1IVBUWTIUfsgyQXmWOsxl1GlI1zJ3Su2QbwLBq2FZ+E
B7JZVgaIvcOLLQLn5lY1LnTEjT1hey6elPh+/qfvgtrq2ePZVlSqu0HdMBBqIR4X
/+vMYDJP7Ud7gABIxbOACwvDNb/WdkhZ0VjVHjOqbik16fyEb1Auf73mtQ7qONn6
i3z1/bTQ8jnDK9QDFJ475ym+uduLm/AR2GofRdP5z3bB6kB7UbmaM7WBVu3tQi2d
WDr/5EE3fY2A6bUkjs7gATCyZX5ccZJZFyjCA8Pb2VbHXnE/DOTxOvG9rLgbyjCs
Q+yhPnsbZRg+l7jrNBW+Vwa8XBMujKpmO+SoI0Xur+vFPNqnaAAddwivIZnKbrBM
54c/IKqPRVqZxt42dggKM9d4WHnRRZV5oe8ZAXU0/lrIUEsY0HTUdRf2MTWjv2nG
cr6/d5RJC7FNpLjY2b0V0BcJ1nuAdXoLuEjhkg4e/ChyQ40sQypSBbYxe9Ala4iL
GIrjNdSchGw1j7Z/k8xqdWhoaYztaprNtjDvyMksY7B7UM938YuuJyIHmZ9tioqk
LO29tRGIulAGQM+MV2xxLUFY/Bmb99IWXopyjfJAqpZlP3O9QSoKb4D6d/qKc3uS
NNk9AHWUWj4UJ+eecIn/Cnl3xianUV5SgO/e+kBVy37gJkbBvJHFosyBshA8lwlz
qyGT2FPkmEyFaM57ixZXYmP/4hi2dKfDFor9Hg60qs4XVRMv7nTbyli0VGMuFoPp
1npekNhJNob+9HC7zxMvR3MzOIyT7cogWRlylamj1ftwzesI1iHC/iOXPhc6hnvq
zaAOyDyH73254NJa9xkqtoLXp39OHW9b1z8bacpFIIoUqdpFmmzXOMf3cyWwLP46
UijKEBxqVoq2FSNYT/nYlGltJyCLBVZNd0/qGyN0SIqfA6+Tvog3/56ZYp2TUZiN
jbLWd524OmJCLYYgHKtkfx3QXREoHTnY02IbBlp2YLScWjQaPYWq9oSgncAGdPn2
z8aTFE18r0tgHNNPg3xHUjq6WrIrWzEwGzcp3bLH+9L3XI5gXQnLJk9JnhIHtIwt
hp2kPN1CPZtgoc36SDLIeeMqIQU13sRhxzz/8SwXrYFFO1DczgoN1jI0WLYf579v
q41dvhJ/f1QD15T1oHmFDtZIb3s/1V00k+M0jWoeU9yKrTuIhZg4goa+eg5dEbGi
OuBtQsLHlWQlulL+BfQFOnhk1kS3UJ6Zw7RykyorHJrlwwqZItViHfUlgtovRn2Y
hk9OC8TVsklj8rADeZQlkDF71huKVFZKrr0rG9dajmIVHJY1ewb28E6Kwa+6+f2m
IXhB65x4Pg4uiCtBW5ev2XscItjI7fb0a6N9BxFResLWecfA8rIQnKTS8FNXTq6g
TqOUYDzD3PgzrsahaMVVcgd2/B0xdZTTV/CMxqdZ/cSsu/jsdWLMPozQjOzQ6e3Z
QvsbVfxlhYd2bcDp4J8vCowIfNFd8IXi+4ocwp0cPuPWcRMNlpXlBBJ94AeYNLMh
GGBx+vPNQTqY00Y2L8aYnRDlsAMYOCa/z32cIIfqslUyCM1SCtSD+aQyPRJ265yp
ouDkBMmQI1hmQ5PUBJKvCb7meSPhj/jJHTrN41HDGLcuHkdfgee8IwtcBa3w1w4I
Eow9MesE4bdMZXDroGU8Jh8UOSJKa0VvqL950+u9hkBPJWnMerKBdPO3uAv6pd4u
QeRpd0mgB9yxfXmc4pOd6h/ViBx7gOkUoxImkE1rsd9J7F9M4efIsoRehF4vgELV
QPpWDY7ZkRR7DCNnOvwi8SetFCez0oMGPAtKd5XAgnPcveNcFL0irLWnAFAVPJLW
qAFZpHYmJAxZ2AK+42dOLZUCOQfHyW9BLraQtTmK1EEDP5/5A+fpkAuMX+qM53OR
NXrv+CFSX0WGX0LyKjGxU6U8PYM2h51wmmnsyD03HhfTIJGUzq0FTf5sEnRzc4Ta
dFRomDv8PZn6cwpqbBMs0F0ZSnTXY46QyM/2xwmnj2G1zWv9TQLN/atLdo+KZWKi
qyimZgw9rbiQmaXntbRMWy4IPfcDiWsySDSr4Aatm5/NOVpQvxD5REkCA0xFXBWg
YbyVyQyeFivqT8Bk5eWgF/qlhDWNzpUN6fU9Q0ceijoATDq/8un2o0Lb0wuSj6xk
pfXtLpUVTBxfHieKp7QheGbiwJKakJBW2GtShqnjUaFzE/SXYlcjfADruk2f4sKg
vfkBSVxhnv5gnM6SrlRM9aHawxq+JNwLiOWNmpF9FtkhYcyNgGHcLRqvPMDIUKTI
eR/SF7B6tQcLztBkLznT87ZMdvvbDPmuW0Olyi2v3smILqF4USEM7L+zDFCEkC4X
V9BnuKHQ8m9PSc3nR9ES89TYTXRpOT1Q31Gv83aCxPPWaX3igkR1NbdfYIoyT++u
oyKbPe5UDyzSgG0AXMEe7bVRwHqnoGJ5fWiNaV1Bf7LON1xULNwejrd/gQqNE1tl
KBiKjtz712KHT8F85NiZWSDoICyTLQY3cuwSw0Ips7JSD8TCZHS5jrNvuf1Axm1d
PEYfQ487UjNk/jL3nFfLilDbKQZQQXziCaommETAHcCqKdBNwV36vxk4UyKcIe01
gM2Rq0Hup9ILl61rHPTV4T4QRrWSbdhNMiucsKKWRsY4XFnTL+4+VkTIENB3j6JB
QLVOCHfv+J7VDtm3kHMw3oWSEgE5p6kgx6z07y9raodAIrQvsckzND0OeF+udNS9
upVhGqdEkBsx8YD8R0Rr7YMsacD20yldxa/2WWx41rCnk4GBRCQ0XVOkaVn3KUJT
VtPkrJRcslIsPh9mdXHCzON75phCwavYeIE9wkJ2XTiKZzSNk8sDy2Q569jM6SLV
p8N+ZFbS6CDx4gQRcnXYWfHL5qLFtoCPTGjnf8nbSODrh5a2//voeTsyQfvAXBkc
vZNy0gyAWPl+LBCMlmf57Hgl6CqTfP+cNXmJFXQx3BF21pai35d9gRto8qXPC77Y
gC7zqnAonbuX7M+PSMvI//jVYqz8ykk1ibbo7WRPsHCijAgZjRK/5w9ZntAQNhu9
+LbHsISteuhXKyE7QPva0wQzeas2HEiA38MZnUIxOa0XTx3BnC335Fptwi9I6eCq
PHlVmxKVQnmQNSq12mE8LpYaHlAqgJ6YO4g/cFUw2hVpy2n+WPVHBLPklOPdI2pl
lHrp1HsQE3JM66tNAENKobC/23/M0ZeNS0OgnHx/CXAzXIkyP3Ve9DvrPdUaK9Yi
QqbXHFOdDdpM/1ucuLYgsCNTnykKbe/4aGT413nQrAuW7Zmma6LLAHBmEd4S3PkT
6UvjPrh+jAkUqai7q5WaiKUDhVlMVZETGdgq9x+sRj43kqfQSlS56PLvE8Z49cze
y1aaLcMog+XH+twWbIEoqlE/bzlI5dwoiP2cEzr04Z3JnIzC3Jb9x61hzxMQCnmT
aIuqqtwodaVZ7DfswDoLTW4C8Ujfq5+BpHQ0efwd2ExodCPi7cTA1d9+Ffd8LIc5
f4WOjKKfZqHAO+gylmLyYR/0acDQvOX7m+OvhqKvDdfq9alKzW1LdgNh9wnGMO0X
HZH4dLX9XY/bVWBi+3u2dJEmbnRoiKlOifitbp038/QBmvKSsZNpEwpoZxtzCUB2
JHXa0QvMYMPc+pGgMKwKHCsfEvUSD1xB9bgZaY78kGEtNSsv7L5rBf9d/hGEqqlB
N1Itaj1mBM0xkGniwKnzQo+e+c7E6tx24VX26xZGKGOnckq+6NMxGoazy3/viIe3
2ckwCCUt2LdWqd1K+CI77c0WyeKxXRXGZkh/9KUDVC4WupoEt/9IEb4V777vcQy/
wWympVBLDdEUql50zPktgloLnk5zYxAJC6ZpOuV7mzclxpOlA5OW1kKBhAQstcJw
2NgDcntz2RlqPpZQq9R//Fa9KCWHky0rx4H+bZmkcGbChCqrQzWCLGE3R0MXrLs3
UeVObbxSkrLo5mVCCEDLP/+yM5eWacCPHMGaUXDWmXuy+FFwgyPudkp4Axv23Sng
PDDp6721+eKQA2ajhgF3p4wAsM3s/D9IUUQICsp7ynPqvPIWgIUbKe/XwZiRzEUk
LIEYHZEcHbY0gjI7KwqM9CKPbXaNvDoAR+WD7Xfqx+utD1WjtfHwNgmS85psPFyb
8mGXc46c+YRxoSOESB8gK0cOciu8OOHqNznr+0PC5DnYyAg8Ixb5C2Gq0Cyzgp5k
W02k2s2Wxn6WUWi5m9N0TEVN4Na+XarWOO6NDxGAPHPkukg6wPgk3kn18W6VCE3H
ArosXFNvwlpReEBL+hv/8oxBw3LLQ0sP91nbb3X9vCc3BL/J5++X/n/IQtNFhoZY
FEMpAC/ofY50vFa+ZwvUXflSBFlte0C6T9xAUr+1ddNTc/r8zW3M6/jP/igjCoJ9
TkZEEZOqyWAnUNZV+fuinGTBB+JgljvDQJZyqa+zSU2yaCSCyAaBCR2UhZ3bVFNX
5wJRcQiFmz23GUCx1RQECfY8y9oiWYuuQjSl2lzAuG+BsRbFVr1vhvd/SiGoW6n0
k3uv5ekoRRPmWyU1kDSwRCnR4XXCv4pKYkOOY3UO6x0W7m58HIeKxHx6+vHU8nxs
VIzvNy2bNyDWJOejDVAakGFG7OKG2DqzER1vhcBzl8MQ5X58zG0jCSpXF+s1T+dv
KM+MRv2TQN+cfdGsLvpC5hIkyqiD5Z5n1nzpEg4AZxz9/d/EDndaE6QqhLz44nsT
1w/P8NRYrfgSPvPoMlD7gCtcLC0JyqXTLTHMNehPgEtR4/38Ftk8Bd5thwEhuQRa
ZFKyyrhTUl5zkE2JSGyzQJr0OXtUUjsM5/zXwjUmhTmfJrI7LbRtLtnGy8N18ORc
nYfX21wkl1tkLQCyAX6EAqEdjFKGGStwvEQRxSraCW5Z8cNgwaKuo3g8YwT58KYt
EQ5kUqJx/srsOr8BvcdP16DmAeLuLXabLl6IIIGKzTzudrlR6NskVYxTpky8nW9b
pPiHros5qqtonF1oE2VLg6FbCnz3bDh3GL/T92c6QWP3mffkkoG6JHdzjLouTnuy
q+XDV7nxLPszkVloKPBvytGbY30nk+OdqqDA6qTP08TB1Pb+GsxJFO5WfotBH3ol
q+wFHID37KUM2Xg35A1AS5cflePNWYS0E9juv8N2cX14TdO2JM7hOkE9/Jd2cfqw
nwPnuuRTcaOPIMeTLMLmXcQkVWxQ3ZMm+ol0biCs/aLCCN0xbfJj20zPjJs5fdxo
wUvBHdVkJOnw7/fm6fVnjraf7wdtjiLGrrMj7kKziMbn7zmjUxWpMZy66fs/GgWV
bTtHFnlBScQ6HfEsnu7F29fdVMqMMFHSKdg1xijYVcQvzVm2qkk7l9S5KalPOGQM
Ot30tFq0l+KWvYpOBvmIC33ZdxQBrWDwcaErDxv0iAnwgrdkGRPwxcpTQe+E/iIJ
YqaXDLxFe3Sla5yDiayv62LEG0LQeHdi/yVyCthOGb3IQdGFLD6RexuDzVCtDfuf
6s/htHYhP15wDkYiT3JXK86V61VygAaaxyJWZ50rmW3L+Q/6fe9bZjDZQ+f4gQ6C
mzItBXz9bH8csQsclSFi8/S3vtYV16z/5bdwhKNbJqhFQ7yf3rWmkro2HrNhLwWt
jFn7jvq8p7fuJLC5/nesfG88lrB1gB8f/Ees1cart8nO1YT17rpeVGEVvjoO1kP+
QBQj7he0YgwWYhSYnVLMOTcpvwAFsWRDxgNn10vsvTU0eM9vR+PdxRnxXs2e80rI
Y4jla2HXHqaOQVBsxXsgAIiKZBiCydVxGZ5xMIC0vtOkRp9xgdKM4tRtrFtkd9Kz
ekaP/cZa4eZZmLur77rDJcjnXHItkR1FXQ0miZcrrTkdVaJBZhxTelAJbOcqdZUF
1fCVc5cxkjs8pBYqe+mhjnE0x4pR+72xXHeaoXtZh0mKemarQSbIt5Hm2fWrpeQN
YI0BwiFwTLxkEUkxNbUoP/yULjCGnz48qiJ2Ms6BJbGWTjDeP8+ux6walxsF2gUQ
AIAAcsY0x4CbpQkE6OspFY3JFDk2SBnAmnMtEuCve+NCzQOs4hMN+vn6J6cqVWWR
LDQ8ZjOehu8ihMkFFjuKDeqOOcDTXi7nAvUkX69Uh6k/0eosGlPX7OQlHOpmSnGw
DnX2unBHK9ASdYGwusBTs48RVKWJ0aDHAVKrXU0U1LQoW8tBo0RHr4RlbZXHghYf
Ln6Xh+jqoyLgAky1s0WcSw+h7ai/DME1QjY2LL0Rl+OdqdlNs9yPME79kf1PLMhm
wdZ7rUqIxDuHNR9ad/9e9DEEZpPDCjKBPnzMOQn+k3MzirvTwBATcZTta5iRJHHx
QO7su1dejp6eq+yV8oR6ITmCwsdZ17A3McD+yr1sO5CkjCb2U/KtqB7DNCqXeJm3
AfSSvKloDNhmAOeQPqSKAytXrODWrGdbEMhM3iNp3ea6MhJP1gna9XpJDrZDNDBM
uMCiz7eWRjpbe9f8Ijn7rIpxVDq6j1oBYHjPpl08ik5GaO+TXrSdipUJULDs+b6P
Eob+Ou6EznXuDTJlo//B1qftcHRM/mkFlrNvXuguXwbwgAGiSbRh3ZqlZjyAfFux
IPzZZXBorT0chAGoxRE0/VrZO1b6NfKPSerJQ6crLNMNCfl9GjzKmhm8hozH/6Zq
cOeyTIZC8SU02FHIY4L+qTs3eYSOzr1/VROjV3q4q0OxC/sespj238yARrnBGa6u
0Rcuqa3J5gUtwJ/q6f9ZHEQQoapEKbchTcCT8ZkBFqgKPqs529obZZCY+h/Y1N1C
P2lFhtqMKkem+dQV2j2cVSL9Qoh8XGsDUIczeT4IVocentUVPxJSLYVBmFrxxEE8
A0boNdfKs/f3yKl8FbEmBZRFogZQxWW8kUiBG6/mDRzClay4DVMQWbvhXbSZVaeC
JDa2ZS0u+omAN/M3QW/AA7XGZBCy26vyGxjWf9D+XNvcu/rOqQxUkDQAF1Nv8czI
Zxese2i+rnsXy96f0qQv3KaKigzdyfw1i3/FJ9oZKvKUTAx7rn/A+v2NgjcMOj5h
dEDYhVDEBOLoFx+P9zhgw91oSMPxuZT/gGYLfo6UDUblUJw2lQ+N3b8pjMZvtLTr
5RXlVWtqIcHJ7VaaP2jtcnZlPDfwl4iKkjIIaWZwCwBXsyzXMV1OADqW0QxFDk/J
UtgttLyXxe14gzAksYuV/SkhrV2vkaB0+/eQYcEvyQLzT7APnYHC30UDIV8LiMxO
4f4Ltfy94vY0PmPryqot9hZPcxrIT+fF1si57K23D60TZ6ykHtDpxDl4r8dUYVpD
ae2gbU+oqMy/Y0rDiQnLPI2N09Fb+VV2I958HJHgbYgrzjyR2KIUv8tc1lUmPRob
QznF2sz3bEWJYY64O+JywHNY0PkFfQuzP23Fi3RZjVML7irAA9xRzHSW8c8sWULr
AnFWXg7/wM3Zfh6EqnJ6OV3hwXDNedI+XGrYyZYIF144gDZc5hvzxSiDUtZZwzhn
/EI0OjoVtZuix20UNWkZvlq046UiCCmmU3Jh8YvdBVx+bI3/9fyarQe3Uu/8zUW7
5+2/S7ht//kKK6tdMs6GqPmSOXNJIKEThjCVXGLXz//7+d/ojiPqbSkwZT+aMMF7
FTDWFGrv25TpBqeSkC2WQ6UjXRg1e889fgAXZIJTxrKP7sVJk1Ybl9Fv0r0JF5z0
DWXwwqWoMOy4e5NZnVJm35bFlSRUKiJOYDpBikl7d+QV64RGqUU2QGRxVKqdSjSF
FfCfJ6W3NWoI5hcQ90Mjg0d2E0SB4mAX4+kAs3RFRlzcEjJEvwv6r6tfatYOKeMm
KDS29SxAszCQvXFRDPVyelochG3TOKDY4n/KhMhqB6MOKLNRvLFIneEY4QeGEHSu
2wo/q7ETRdGNrjbL48Dr3J0S0jN5xHXijBPyEktjXG5rPrCiPiHuH6nQ5TaqdCpO
sxPsuSYjj5U1ds9KVuwW7uK2Je53EcvhGgIARlWocY+nuDmiy/ZxSSN3GG1brB13
FknYbQwTJwtp/O6Ry6IoIUp2dcnZ4F9UN7JQi5OIMzOn6kkTfml1Uac6WPlvESNt
kyIF8qaSmrxcCQAujY+WmAziN9hqci5d+4l/Iz41jkMryD/zpq4gvFkdnnHlQ0+9
INzO/TJ18VDjmjoBIMz/pfMf8s0lucji/QabzzP2zWTVsiY8D/masA/47cMV8NN6
d0DoZw/hl6c/lsCRxXbCA+mS+rsgLPS0hr55uKFXPLZU3seBjMW0pbcAVmrR0fHo
461Nqqwc4sjs/y3pl6NKbCylMMrDh/wA/kjvkrJ9VAtIg6H21cDdegvi6P3WUFQI
n4JtUo7YpL7skqslAsBd0pehsdpJ163EF16KY1Dlhq0mGzrjgJQACH60JLQ+ugq7
V5+AE6zBLTJBSsMMpQ7p+oktc1qgblItPwuW/ih0wVr1A/dBXWkumNsf5YDLFJKJ
w4JodV5JZzEDiYSmJ/BVAzXP35jqzYaopsIGdcZ976i4vZYom79dE2HqI6rAYY8r
DSwB+SxUI9Gt5aeRCFJNrSMv06pIUq/L9/uUwbSJlB+5jhOLYjj9eQoIhiEi1wNt
8/3LsB/S5EABhWoLCFIg4rpWydUMxWzSx7KzyndD5O4m3YXbaJbkDmpva2SfcGjf
8d252Dvqawiz9PxiVrNnwRQu5S/ruePu2IYihOqItRQGEkDIH+6oJ9SiWy9ycG5X
huOyd54bU7AJIEnDTwet5zzpXCfod98387cgQvAIU/AIwnbdt2Il6OOAEdjbZUIp
n3D/R6GWprVA1e34roz67tukgdPzfwSt69ITMdXnJTBN0/+eHasND1qyGRcPW7Um
xTZ+aAROHb7bmBvnMd3EdCJ64iWUXjOrtVPzcbhODoe2VqKcNO2893PlGRjHq45A
czuiYW0PAf08zocwdCNW0IAJ1OBG8+6VtglZJD1n8rZC7Z64Uopssa47IAmfgNr5
14nUt4fpIwfpjV/wFlLivQANMM0+FL2UwiXkSShFpouY9fnVMEevxWIvrGybo2M4
jnnYKHsfudPNvh6KSxrvtrgi2aNbx+4Okk5NyqSeWaNaNOgkl6iRioG4s9gA4Ymd
g7ioqfYVsVGuXEztMsUGvrP4vywbkpiEtAKrkpYSsGPiJXIj0eSfPUKNUN1NcuhE
9PgKbm7hNQqxAJCy9pGrM/lYgGAE5mJPZBaYohAzUL3DH7/kYQv1YJCDIvH8Z7tR
HOWE/n7R2zclByBiLcHZHj9GVPjZLCGVADUFOnzhLxk4qMKQSkyJjr1MNr/NdYCf
KtkMMs183cujsQGT9i0pemLvUQZ2S6EKeBmgYZ8D+EepbrAFLel3efGQ8UFRlsXx
gmgchYGpq9RA7dUl6R0kNxq57nuFkhnoaX9MG/A07Y68faMCVU8n/M4JtTcsofaJ
hCrvLFahEtETN4SCwZawP2AS7WXFbIetse6u2nsaSF9lOoZ6mIQywDc8jWJ7Dt5K
PzZFPu6+ABryvmd2TO6VPibWmns3UhiAly8qnAzlM6pwCL2MiZlnvLZvvvX+28+G
jXOSwzfAIUrqdbcUGE0w4qCdlwvkqlQHPzM62/z65rr3QFq8K8gANH8G5UhFEZwb
Iv2WVwELLfepsdzgofDTP05kYLydusVMIfNhXrMRkOuwFmPbiYC77/MbEYSjvGNU
VaMXP5px6EfMFY1uIURyqEKBVtdC9gVB+UUWK6fuQhLsW68mw69zxjnqsNnGM973
ksnwXVyyXYfLu4Y75oSriqUo4rWCqhuwKly7M0Dg1xvr934a9ws5POj7pImFClYW
ww0GFsCAnx3BzUIDmgNrbFL/keROiRSUwfKnvDPEnlfWJJ/twso6dF1d+d+orc3e
BmZM2KWmJfo7MLTlSNRD9uCKomtsaXI04/YY2739L/JCzao1bHOd6MgS+ac7DUH4
Sai1x6YAxiSRa9TREUjN3TAmF8KlPFjJWj1YxraoHtOWsNaEhE240iCC/YQcsuAe
Lu9hVCHFHF/B38mR4hRNnPb5jKcDkMtgLbZ8R2JZZlmk/y36EH3wkqyLHFLlMze0
tdRwzRdHr8XGQ7r5PpvnRWRVphN5DkJ+tYPblL4aOfhfUwCG/rAEq12hpYy3ejNP
Qx93QQEM4wAhAv5SvSuNKcjJrUICMQ63Xr5/nDtsNzvzvViqZvzHhke1nLmlYKbN
Zlk2tQ/LNUGpKR4rHQvP+DZU7dTBe3F8DWaitp5v/zz+L3YvU6HACDYqe3Ma7fVU
v+tJDIuZfoBmO0+cC78z22gcxb7P4iE8iOAoxXTsL4H5U51olmmYrgj1omsNyk9e
r/rpno5Dazb/s9k29KVQ/q+QvJUP6JIc9I+bXolJisV2xDWyPc5gi3jCvCWtVE7p
yyAPfW2aBlNFvbn4zXEliGp2leOCUmiyNtwc5GHylqVTvqAErZGTRPGkf6zAykhf
3AhyjJVb5+fnQYSPqEoXJgtO+ha06U7FHYOKndwdDmW9vmM2FeQMOu7NZR+yc5YM
cKbn59DZ5H8RDcGOyYErOx0ctLCNqheg9othOGneVv/H1yK9qoOjUsFRk8nFr0v4
wNnoKQ7YmbLv41iASZ2Xyz1dKZU9JwJkNW5pEkiYnC8nyEeAPZN6d0KgdOjF7M0s
tZY8eIv9JeZOUmx83cTLs/Yx8h+DMK8GVP95tqlFK8LGHhmDv1sUxOFJhnIqwf27
A5/fZvU31Yzfd3c3WdAYVMBuyF670RICpmCr1mOaZtmqG6ZhB5Ck0pe32c6pgLZt
HuEgytYucjk9bwPRZFr6peg+m6907TWUNtV+CO6h3Qxrp8TfuHJmzp2T910OQJOv
ZoNt7CJz4a6BzBQm8sk/txeZJleqLsu4GtCj+T37A1JdvTwTh1hN9jWoDDc/hzhA
M69GZPvuc1eUjtzaDO0LfhLs3fXS4Ah8MM6RtFDBVFO/rMhLjdy/x2oX4plh8kjW
mvT+JhwWSWkrLlhLbh/oXqZ0efF9Wx59Sn6wUgxi0AzpRv/fTq/rku0YHCrGKb+F
nMHpCGpO9fZ5+GhAHH6mtIt7eneYqqO7sE7WPUvmSpmNHe6SGWN6v4eIbVkS4E0+
VWRGvlCYC3wAI+yHQCwNihchgwAQ48f52Gy69sl1kG8ykd5fVO4Ou8DR/bhyfaGG
KnL+8X3bq/VMV+e05XdjSspkncN1iTBo8zmi1/0zpb5H7fLlwZ+zOeZiIFrYCV1O
I62YkcryBUR2M2A0z2Z3JI5QYhA44XZ188RKKe6GghxfqMWREsO7iLgdv3/yIZ4L
D+3nCBeMymsjyYgl1bTpjHp/M2U6hQQsRFY5Oi1fHm9CIFa3xipownV+e01ayvGd
N8s/W3vP8uxHbHr+AY0WmEANihCsYsLiy5SB0gHISFFCjpa2wW+sG0z4M6qq/O4h
Wm8ajzbqJG3PoQEBNJWUJKYr2riyhpEnZZDCCFsYN5n+7nTLEkpnAq+6mPZaavAb
8nhHLk05EbWGznv02SAdoEgGpmsbSe7Xxr5gxLxiHlZ6QQFLN4+i2oOfg9XxeqaF
t8B/ny9ga9Q9jp3WUH0qX3F0NIAm7D+Jsn7Ps8f1BFq7IjvjIWtG+yYXFojhuuWb
F4FfW4elbHgHkMR6oQnPtpWn4YUv4BaU7ZG1nNMoff6S+fYIMq3iV0q2djSa7l9t
MOgBLdQro39FtqHkrfAAxy4Wm5qiOCHOAnmRGjOVzgRzj+UrSSM3GHitJq9hRHVW
RsBeB3A6cLNaq8UsB1g1CpWwXKvhtMEB7nz/ogn+jVj/6utiwkh8BqC7a7OxafsY
FWo1vuUbMFFQUdO1WB4Almj1kKfYc1vNb7GSfMY4VIGMPC26lGzNlJktmZxQd2sZ
uZsup8LGnxVfnfkMv3LOpLg8nUkGc5EBO2y5wTSUktVa6a4Smyvzn3mthY/H6Rt3
p1ybHr5dVx5UBUe7QnIRX18oCpRWVUxZtUcF4qTfQoEJfrx3Xjjtav3GSPrZB9m4
bOnHxttW/4dztoKeLWSxpYIFJzwuFWjQfYM4afa4jldqFNMm0xSDm1f9yCh3ikxf
DFVcb24qgOblNW0siEL/lNmQBzZHOsoxiOE+LTabZ8cYdKDwT8wULS4E8anYU/hd
MueaQ07Sml5pq0D/Fs87BXusapawadMRFb7O+p6clVQ7wfGIfIBal2ZxPuUZmLv+
+2SC0UXWkmxYwDvYHyuxyFjnS1EbqggTsyRCznKP3fBcctaRi58GOzbXH+yko5pv
ZRHEpGRYuG7K7gBVVXkdlWDMy3XiA7xKtXSlyL7VWrzzA84Xv4l/QxLfhYvlZA/m
uvojuFTlsJ4yPjoOfE+gXRxUjhLE3r20O0iPlN/rXmcde7+f4dPbsN3AUHGfFaZF
GIkupRj7YHZvMSFNCh6S7+/+dp862iGi/lFxiL7Pz0kIXKua4k2oMpevaXzXLeej
0F3RNr5M+rB0g8o1r6vPmd7Xrp2SSNJVXSnpmKjyDPsU5hDpprsNgtWTaMrCO8cr
F4EFf5g4+fMnrmwT2NVboBhf96Bq7qEMHhdxg5f2EPArMFmgVlcaQ+p/eXS3VwF+
b7R30WU21m3mgGeA3pMzeBIwR3Fq7r2aBHkDWrj5vFRvoo5JQRPagdpkyDjCD4wc
XgfXtT/rRBdPOn6H2BrkXfoN+Cq8gfNDvyFS0l1pZ2RQX0i1p5mAE9nvuz3OzJuW
23/0aFJgnkCu5vrT/w/sSqROEFBzmj1zfjbmdnAk0qAlmYg0ePSoFtHhLdk1LgiL
qwE+6F/vFLIo/ubjMKQOOSGBH/EvTobomhuVrU9Ax4epGRWevFjKSBfmSuVTig1I
sNOao+DV9NYB5IKhu+GnBhSJMSdODZ6f17tGc12zO0/yKyiZalC/QqLDaB00ktPz
h2v3OA0pmmXqqnWidM5AW3/G5gC/l9Fz94+piFwYSUQct6OCD5oKJL8z56tiWyOi
V7fcEusFpr+m61dXDPHo9u24rWG/DBr/SaCOaWNyCfZFeujLCYpa3M606CVllXI+
bMsTOlr2vTUr7A1ZRwatSQI9tF6sDGwqoq8Ddr/5L3UQZwi0HtsZdWgYlJnsqHhC
PJfoDRu1q73ber72LBX339xmZVQF7kWI5xeznS2Ag9m7FO13lEHDoSjxWFz19Lud
etMwo3CVty5Fg3qRTUR9jIz4Urwwaa2z02CmPqJJe+QL7TmH9oIYlGIFk2Py+T+l
gouNmyvvw5+1JjZ2ECynOZH8e+IbcCz6ZfSrOPpi39qNhdPWg8y8UjL8wVy7SmON
Std8MSlCaHkOoocnGRBxlZKkrVwNLKzQSjnDJMb+FoFEhJ93kuc/hIXP+y6kRNec
tEPi3V1ArnlAB53ksxEbtLEkLHHzjMGwoi5Sf5mOmMG99veaSZlxExCFgap8GsQp
jjNgfbLzxGZ/IL+n/TrUVShPqdMMNoJtrlJZvLeNLSbQB4pj35IsxsIKsDslk12i
vN6C6RoDmNLPM4Sqm8Hl89m46+JE4IQXz1O56REcXVAED4r5jeAko/dni3fZi+zK
1FQZjAcU7OoE05fCirrRVeathQ6kozYyd9aSqyOK7bZyUZpxkCXomXY0duzx1ikh
gmkxmKLgZ9h0KN5bRg6XzfKhQHrc0rV6v6XeVCh/aSSg9XH22ECW2LghR6T4eOTd
5BhO32cpDk8KXwcJjbLdn2KtzI8RpGeRuaJZjLDNg0v8GUPvnnsoOnopN0VdX2ty
oaLV0NvAzoQMgtNaXdATPnJUhci39IGiQUuvxVpgKKFbthw0l6klT3ON2O0ei5RK
rperACaB+8d7AfxrJKzrGpJkD7QIg9wqMmvZ9jWbdZrvX2uIjq3CYRuPP4gBWO58
Rdp3CHe4Z5i1qx3uSZYfLIkF51yG9vrzIkKQ9eP9dYtb5y3GJSHJ4SnshK5aItDJ
SW7lyhfPATQwNJwB5BImqe7dFjiGRftgd5SzWfZ1i6rpsZzYj2lOznSiKwz4xkBP
qxPL2yE5r4aLXChqE5tSvbpL/qRBrBSVfO1xmkeNRn7TFM+sZL0JVz3lLpgSO2fq
+FDk7ByzLj8XRKm4Ch66BJNiq9tDUBvGW3QLFzDjPMu1vhXe3nH7Izx7SyQfkLXT
rXStTcSx/Bz6XGMfbkLMnfJmxLSdNbVYdZSPoPcB0WSH4CRZCDouGlfEfZcWOph6
VdqzahXEvOmPUWkMKSndWEfLhqP4/tyhhjxpP283PD75kvpzOj2nl08Pe4VnP4KZ
RYR3wVEYKfaRByQbYhcaWQWxy3a13IC36TPFg0lJEBahqeAQ+hekyioooVziKpcF
6L/bivfA+PlsIh0dqoeSvqkVijnnO/uWSjfi3J4ZScD4LiW9xSy1bg8yJ+BTFNaK
X8CmmKIHNSKwXbBH6/FTNU6WZZZyC1MfWuPJySykk7doWLCj8Xj4lRgeygpHqxgC
LCnyalSmmNcdp/ycOR1SnF6ZCg67HLAJMozKRHz/w1oo0MLJcY2iuKmuoKzP5wqs
Y+pvedeY0vArTz1CZW6UVW/tCyJS5VdOBOsBcCP2llDxyLONS1ezb01YDJvpdJSi
4IG+z29jJKp9t0iP0Ju0SLqZUhyLj25Rstij6P5cw92wuLxzmIUw83BhkjkppLe7
a2EGsD8CHTiD9wVFjh/E/hsCviXKqVP9JEyw2fTtJOK4TnnOlyFBwfJ8ibunP4Pm
PI2JKwb1hB+FDh6TGO6bWQV30AdDcfpvu6ulpHlwGtSOx2VwRAdcttJvy2PyTrZk
soI/BZflWlGGoZlsPB8q91ufaTTI9X6L2EA5gQMfyCiRIDaJO/ksc7FZvJscFlG9
IynSIBmMFTOlNjyWL7hfhEL8mG980GkOigE2R77JKkyFc3LqJBRmGzVqoxWyU/kH
JvuvWWzK0j6iOgFEUlZhjLyUVmWt3/2sWnwLlWe1A/fL40jPjRhb8tRxVF4Lp1Xt
fFdgvFo56MAqMq4xrRQ4jNOTCSg9hz2rLpoq+SD1TnYfuvRJGd3s97hsnXv9ysvU
+UQiyUHHfW/04euZqBQBdPlRfmkwuRVyLVAVoLz5FxocjXyCQQ/tucLhLnftPihZ
PWikuycoXNgqEsrnWARMkFS9EieqAIVRh5EmrEh8IGMXS9u84EbVXX8P16B4SMNG
ROXgzpj2wxUSHyGZT2gy04pm7uqT7lK2JB87724DkS0USodeYvYxfVIdjjiBTS+Q
q37i3QvkHVLneY2NPwt5jEdoJDTxs4maQy0gEywCu2+pRvc7aFQMyDkvjnTMhNM1
s7ZVjAjzD6gtukcqxcZfR+DmzqpLGCMv/39cxf7bsjnDWtMshNv9m9nwvMtYE9Az
7+7ep5Ps4WDdO1uhoAfVsq0vAPToS22qaKI19fCeEI0XYR0KjH3tWEAgknTLFSry
JiMvZJRdEbpDivIV8R/XeD2E7xT5zPlk0vJaR7bojAabwfnWudLE8IwM89KX9whV
/HklItDZXEhb9lFyHCv18T4QzHxnDTRBumL6iNqfxts5gmmY0Xp+CzhCfOH3rr1s
uHOo1Px2TBPWVcPtBXTFIRmdUMb3PqvlboulqkTh3DKwTZvO0EvAc3ZYFHXdQ6Qd
crlS5P8cBs4cPAWphGXAiyfo7b6BMXzOi0/eEAZb17mn4LvGV+guV9sVYpLj9vDW
HQ4DcPhx2PI9PrPxQ7xqltHDI1HtruQrPHBu+7TCI3egklYiXd1QhZnupXFHBGSk
fmS9lygCiP+kAHQVvLuP2XDI9S+0rIS75VHxHkKwluuuv2umwAgulSQYHuHvAsLO
tJ7KLymDE2g9sJoWUJuS18Dz8arrQQ6NgcPbSe+PLNqt4DYgEkQFiKXFIZoSOmLY
5uoAnxHCquT4vb9PBx7XELiaiQYuvVEEfTFmyP57fXeJWuKcfjgtTJ6urDhy1V9m
zx2BprRWapWvBFcxXvegeKctuPz8v+HHMuBNTFokPQfjn6JuWd8t/Y7eL7HwAmzk
o/V65EVIPyPY3UQ2NLBewU1n0JCvTLnpKp7c8kjx7OUpOmuqEiA1GxXQdBsG9QwY
FZiRLAjm9eBhaSyLJe9YhwrAY6yLqpYpFA76X45Wid9xpKfyb6hXjnJHT1RQ2o2o
Ox22VMpLUpEk3wez+8wz/vLLLYl+cg188zztW9IMaC+UwAAEHrtEIoEYZiYGFBhD
wFevURt9jkooT05UAJ2sxtmiRZxoUB59Z+RCHcYAUL3P4Sn1qPwpmwT81+rpn2sR
zKt+232zKJtUROtmPLVD3HpFr+4QPtZMYrtyfLK9igasI7vtdhqkPXe16Qu64JAo
4A+gtUv2GPi2Kqew0o3x0N8IsAzggkYby7xOao/wWEghcpr59mjcv7JuZhiTy4ud
iXIjsAn99pXk9rkdXn+/1BndHb4D3VxFLWtRv4lk8L278yz+YSKjwjHbXRxV4Nph
LPUPepH8TeLbLHAv90FDqj/dI0jUgzEcN3P27flnhKLV+AZ0DnaLi32fMXd3DF7u
gmLSGatjARcG2PMeOoBWvZzy6BUtJmTu/8KG3oXsnB5t4s91aoEcwCQI3TGzrSc/
wfxsK2bHHqixq+pUnjlWeFPPzw4CrBKXmcxNJKDjcv3rpeY4V4qWjgtqAOqotiw0
DPU6T+qxPQkwOF3A9uu0EE7xOkv7BZAUa91cuJ2e9F8EWtYSs2nMX8rXmT7YtZUK
TEvzZ/9gri1g7bbc/4CJVGdDwYdapOydjBGT3vpL0W/mjmMIhb9TG5jQ11DE7eSZ
JNp/DJ4j3URMrA6FhSzlgAtIbQ5AMJoxmJrQWp+T5wIruTH8WrRqwxGZXUIn+3XU
gbpHf5pMepdt5CWvW88TrZ4kHT5DP/xA5HeBDeFkpst5ULHzO3KumrShvxcxRKgl
dUw4x+4ImfwLtJVD2vRLLGv67HlU3s6FNrDRooAnS0zKiUceygzzAS+4TqY7Et5l
97ODr8OZtkZborJdVTiNguG7Y3jnNIuHH2yVx4MQHk9tqfOEtmlCD4FjQBgwRbWY
HMJ49MxpkYkK9MWkV26Cl/hBi6NjoJfumwgs2PBYcgv6EX5sh2FwLaWZGEhZrrC+
9gnZLy6kqCNZRnU2UvN/GyCAWd+ge5kxiMZkkvKe1iEbtzBYIJcMR81D8GGF/A7I
DkK3SI+8dESufi4DpdO4w1l3Eghg5NCnC5Pq7p1eInvfdKMT/K+q/NGUtRraXJaj
w3WJ7mP4ApL7xMipL3bOMeZnXWqF4kt1NKn9PQR8AfjZV9VWbfTYepP7cNXBJNG4
Iv/yqAeFf9tgkxA88ky4kDt5WBYkHM0xx2Uqz35buYFSN6Q7IB10rdTfj3GDKVgY
nj/igg8CN6QQ0P1k5hs+UxdW/SO0RACfQdZU+Hn1+qFBBn4vqMgsknfXuIyK6XB8
9wr1PQb/OP/R5GA3GHyCGcNMm5B1RriJewjq2V7kZVO28hq9c1PFfznTk7cX+PaR
MkNyLY044Ph6f2gIo0a1G7Nf97hx/x7mq5uYoS9VERB6SP6ozxocmGJcKUNGnrou
uZq9/MJHkZ/mvyeyRisf9PI4+PPrl2/viSthYmBJVgWPz7wOmabjm4V2sxZFVf//
AItKd94XOiTR7dPaxUktg+Pp/o+qh2Ft8NmgQY7fXgQ5SyRIHlqZMy28+YjX0LP5
1T5LoVo8jMiF/WRlOq/r1I1UJhLjI3vVXVH8hTw318OQTRnWq12yxLOYaoS2E7xD
efYDZOL4XB9EacdeFOz5Xh7ptc/+fxSt+wQtaZwMC2n2txipg+njSguvSauxt6qq
hIDfsM6MwxpnpJOSkW3yNXNA+f5k+oTTEO4AjHfFPMvWvZT7fiXBBedi9kHTJGBX
iMCltP0vPciGj/kk26vNYQiIwOmXYKeeJecSV1l9lA4PtfpY+4CowhwW+6toUS0k
hROM0tGiuOdTgnzO6GcU02cJM+8dx6GLzywASbXobin6bZlKwKpAZZmnm19epgau
Sm1XQQhW+gh+RP8TeTlHjJyhkLozkIcqIhVwc3y2a2HLMK/dxUmha46cumIlluqI
gBWhOANyxnLE0YjMZYODiknEkFcxXPXqsle95oNyt5YpLYiD2D/a9thFf6y52xRp
SlF4MATjwJ3UMpt6UbH90hi5FYGCwRYWRhzTK4y+5JZxdMSoblpwFoAKgSVWU23g
7gv9ddBC+ReKStkCQYbaCqa1SMWPTMaN4iYpAn0RjQtlfIUFZ811EIX47zFtDZY7
YQsjEwxp1wYRDaIQHErgSljfrWj8nH0eclP54AErPJM8Tr5twwQryiUJjA2232MX
2yFR6kEZ+k6KT+qBmIOqV4Pu7hucAnWv8BtNy7PbOzf1lNQGbgw+OXt0cwNPwPca
Eou66TEtxfGwAPS3ua3x84grulZyIJTzVF0VB9iJfQ23GBSB+6KkGbgFy0n3n6dK
XMXDzqx3uclMkc362vj5YsgWVGJb2WufmUzXzKTGkPE24dtLkpBJ+Br2e4t5Bslh
j3e5u7d8jK++Stm2N+YhAfQ/aE6Nx1smLjtPM6DgFhp7g1PcoeTiAIMacBCColP0
jVeISH+AUur60p9DJbFcyNn1QMFF1zvyr+qPLoo9AYzj4S6esZATVJtbC4ZDcvAf
8TUIiTCSc4WFIBXzUafXeZvQpZyAURS2du/N4X6UQnv4WiLksrtZZCkYWNjYANFm
0JZuGFy+nWWEwnsILaWM5mxdgLOR3qoLjZGLv3lDptIgqFlkClbaA2P0aEtgRwfw
PxGfZRu1SsW/Nk82jT6TYoyJjzBvSF8NaxLqeAw/r7AZ2r4y3OtqdNDdHTQJ9p86
qQdP6oMhVuZFSL/x8LN1AT+iJqv6y9HA0BAojKG2iOYbDGTw2lsvKU8JQyNxxKer
g74aLrF2mu4kvqmHZJwCnxuqgcppgPXu99Yxc71C4tD4Yd3kOyK8LzaYG4Bpt1UZ
mnNYtRP3EBlCQR8VsW27gejJe7o7VX5h2+rwFLoKyEuaPIFOnxyzR6LS+tpQchqx
CXOZz3UFQ8H2CbDc8LLJcMYae7d9mGF88ld0fk3zmwk25mt8IhxylJPfG8fQRWui
hmmMgWNmuAPDJ11VF7W9pXCWhyX8tZvc4xDNF98Gwyv31Sb51JeWG/aJ2PRbv8xv
lUfEfYDv8wJPjL/jRDoUvay4BHUkWexVWfVgliIZaWsucIJbtKEF7U5MO5XetsuN
GNTB/KQ6fGJztKkXaA1B4bUk7yOkEk8GDabc29Tc/hkUhKp15WO2YjD5uGZf4GVM
T9wL2R/nJ8tIP5D6zgN4fx+3jEVpGg2IKEkJaKXTDg6XuiAN0syFe7Klz8xnMqpI
+ymRys+DTyX8p4SDnsfos7pSxukhCQCT6y69Jb3Z0Zma4g634aEEvcj7sPcJWQ0f
BCWXrd6Hof1Fnmbcw4QRct+xlcX6d61T0UiQzOheJVGEvwxc8D8hzM9UYSXTqRYD
j/A7mdiaa+M1R4awCHTDgyA2+2HqtGWsLkhF7QM2fRrqEsElxsqK8tIosJ9mxCZw
Q7kKv5bz45G+zvoDlEtIFPwT59BO29a5nVST+ijlqga5AfOOuVQAGJX2BBIqWkpp
vrjiOVV6iv03fNRMGb9xiuMxjlYA37Tbo4c0puA9SF7F6+cgj5iHIZPly/OPMBvX
e+iVf58KtGaxHBNWbHl+fV2YjHWG1+x/8zW7D6wcbqr9JVNyvBcpm6T4bamnyI9N
8cqo5YcDzRRMZNGxIdTyHbJtFBzKYQ5rKbeusnRHBFYstraogB2urIgKGEG6qGD9
i9y1yAgBjAKFeBZnaeG8G/hpDOQGxHUz2LJP1Tb7gNS17/jpte6NXrl1P2bFuEYp
3luiBQ3kCEtn65lOLiN3c+kHZ7jCVSBfYIz4L+cZlmnxxsIdZjxyFSH+yjvy0i+b
YBA4F+1Q+cNH7gEIGb8Hpr6nmnfVLVA3TRd2rCcCn358O/nmQYjGkBByB6OiZFOE
qUQXI4dtNrF4Fx+rsoEOuaiuki11apPk4KLn/CX1hW+wXrB3iax9uEzyiBtzWv5s
Wb3x5jehcfx9wtzY4Fwpk0zYmhKmhnto24pikC8sJnSBhVveLkH1MzpV3yEU2czu
bRKi9GRHcpf4aoEiLRcDWFQlLDRMlvuF88GqsyMVjaSZlZWE3Xxo3yr0E5bsorcT
LLiN8JX0Jm/CHa+BIS5WVk6Mj74g7f1JOYV0Sj/JdwF/u/zlepBeTaMyBlu++fXC
fnHoDRIyjlpXD6cl0BJhoPvZGqPgh6znfy4p2JmUa5yboJsaFMx7UVttar6/YMNi
VTxJG0X7TetWtlmTfrSJu9hfsyw7c6iSETEygHkWjRj36IoOL8KD2JLhRCS9yRmK
pi2o5aofCK1kKjdaTVaIc3oItxt/2dbRdiiYKgYQxa4nosLs0oJtertDv7M7JU+s
J2kSCJwI8vmIthIzK8Kzj3kvrpV9C0MtXY0Aa+RrHGbrYevwwaBXeBTORH1LRTI5
w88cvXxRhx/AJaBXFj3GS+28iZ+0kZp5KwSRoydn5l/U5suYqnQETeqi90xpwuWr
Hjmv/7j/AlBh2QWUdMzwQmWc/2YuuF9eCx3CNuIcpXsjdr+esMFa8Qy3aDRL3Ccs
45PpTa1ssJ0GVqp/6hiW8x/u1QzNA/sPBwrMpvRAKfVk55CLZ7AL0iGCuOIXn1vO
KtVWMlJYZVhuVZWNoR3WXZ8J6BAoxFp3xD8oMoehchXG3QtjxU9QA/H7nrqEq5Oa
qX+0LtRlUTQn8wQ1A+wS0fi/v74sWlmKaHueO3vs66ouls68e3uPTfMaQbFnZbc6
SBkT7KWkhyc9O88MxPgKno0oxqo27M+nORKAF6Q5OqxJI98i+xPIAvaYCEbpSSDM
o3nQXOsjD4QaGDoKWg7Yx9zQxYyjfBTaH2HeiXqH2Z+TRZBhC9MzeDUeaCWTEluZ
XNyP8JN7XI++4NfHUlLthhQIT1TU5tOjIcAt21C7+EHPmEuS4yhcHadFYSlbVK5R
BRtBLeP7X4iD9CyTwVgCbf8IxDCibe7bZaHbhypcTLLtNqRwLhQRGhKibGMmQS3e
NA+srw19qKb0UBypYLrGq8C+sLBFEyKfYlz1vLDcXO/1iMocrsNTsP9oJuq/jAYk
CerRNeg0H9Nte01T3A4ig5zU2pwIJz/H/pQ2Zv8ftRULzXH/BdRPZbO2KgbUGC44
Zwj8metmAhF7Q1kQ7hF4HyYU3vYsqdpMC8AXGWys9fdCGgHv/S6Ilfy7u1ipl9s9
S3oABBjc1Xt4dpB0eCd6jTKVEtu0tIZQjOX/a7NGtF3FRz2TC++/nXK6IPrWdj6A
5PkYNxMoyTAIieJxeZrnDGzzjj1NaUazIsOhyEeRvhI9Udx+ZHKyb0LAsTFfCdTV
AfxcoWiAmrd8IcAQ6HYARvhE4b9wmm2ECWkDZ35HeHjzdrZ5+sFXluzstgosebK1
rlLbfLboLikqBxMKKMc36wUa3+858pzEALJ1wKuayayur9FFUR4c/NEopSmuswov
p9liFxyeSbCm+1cSX8Pu7tFEMT9NiYRmFAfakHJURcFSN98EXDmRMmSCIydmPZl2
SfTE1v9SDhrTvzz6o42bEr1HlXrfXzFGiERaKa77QDfbBP8MpU2Hm41fDG8H9HW1
IICGyN/CCAnY0+N9JjKjUeyeJaxNM98zGZRetFL3jervfntCWAkgrOXRLntJH7EN
x3ODarBSEaFAJZHoeRO2MGzRLvooGEMCltlyniqUGYzp1Wm0Mao2rLEjVWsAcKh1
sA0g9+w+vOTCKSp6iWMdWLbm7M4GwSKXZOf0iY/oNs+gDP6qsny39KgtzvOFJGhN
YN9mgoZk+0XJ2Rx5AP4H6r4NFHdHra6NuQgX4KqvL35IKcK8pHPnMXtA7b64qFht
KBaH7jPLFJk/PlmrXCHit0X8W6rk9zUFItz/iRbjBpgi5+5VbHVIN90V0+PyXCLM
UYN+3v99NYcDvcwv7ko3B/E6LaXIxT3BjBZKuEP3vy/PEz1uhGcSCo9JYrLeIPlD
usKn3I7NfI9ywsn2Wqj9w7CwkyOuH7Ueh95X8A8380d6Iew7vzWRCipv+HwLc6zW
LKxH/1JNOmJhB0KfYaApg43Ef+qs75fmXe+QsUicxP7UVWeVF9040JEUDfQM1u1r
Q1tBfPkiGddCEBQQ1Al/tG2re7VEoklQdgX7ULVN2c7lsQ2kpHQjmIup2NwU/xst
FGNYwtMJ2j5xfylnaw22lemVuCvJ7mTLdhIvBoK7e+7evOf1Ru2W+Bde/lxhjfJC
USaJxmW3lVaLxptjq0TQ+TcstXoT3q2Fjr8u6OkCjjXhbNq4VupjL5H0SE4OvXKB
5Pd+sdArDBI0LAsKwHa7Uhsksck0zjatejqganLz7hrZavzE2KyowEhz2bEA8XBH
rS6ymMNTuqxNgjNnyoc/f7HTRr+H8se7s3t8+4TKp2YLRqOPdZ7ttxkmTaAWd7Og
s8yZBRFgc0P/NKfc7BcUseGUyvFlmDSwJl52fSN4S75mZ0OWVtA4Kw6+5nASMgvC
bmecZkJN8ZRh857CPipxAgCRKscAYkW16mf7TXTNp5isF03AFJV4duR7apZkYBZH
g9gi6M5lDWMwOq5bDwybzloCZPaV0NSL6lEUyrmieCFwfV5BshbUZHRxzfqn1tPz
pFzRq1dpT3Y062udz1ailcJHeXSwDwUaL0aub0eiBVFBEL24Gd4LIs4LWgb9U6lf
z1k8574+50aAylbgjuoSFh/EjFidBMbyLbEDtprOWdZwQoMx2q7c7xYMEXJ132d9
dSdy9govPc8A85jLuIp+ZUdzTfoP/bxQGuWPylVEKYvk+SSiNu135gDN+xTsRD5K
WVaj2Lp8sLXiDhJoRL4vfJp+zffNzZwMHSwcAztaa2Tyj+nDFdJRELA0B0dYVB3N
aZ6qqQ0qnC5LNDVaTBSKpxb5mACY7beGkQX7m46EPV4KKLrD2Pjr+ANAod0rCFEl
rqU4ejE57YXviWDXw0Vlq3/mz4JN00zHOm0kVA5iXx90xLcwcEAPr9FKmBxGy7Db
1ZBeUk7fDgqsTAiefSxHAzkfncCI0XgIvC2NOFO7SQxcUpRAh3AIHa6YcVG9zDJU
07LgI6SLl7FQD/1rb9+6wSSf3MFtBQb9aoFRMJYpKm/PZw5yw57dXCNfWIC+FVVV
6mSa7lii7GGE83rGROaUEdLEJH5ZPCSvSeShOil1Q340DK/76jOFIs5voX4Sc2XN
2hGhetZ1fj617Uaq6fW8t6IYCN0JFyBZg5JrGYwaVSH1onnVa3cHCOXFx8mOUI80
FFT5n5WKo4ZVRnGshdwSxdgqDkG094X+/B7nyiAr+OVxQQekriIBZX62fMUasl8X
MlbWJ/in2ObSlPgflhShWwp0EuCNVpuRMf8EZo6zc+UqQbhr1HHnrChhuwAoWUXc
yyyLp/F2RmmBLNx+QjX3vQRZ+RsZfc66rpURrUD3GpoLzwwEL0RKjIUJpNl/oRso
zVvMeyNSIt0bFUb89kW+aCy12lkd/UwlwoNMpGL2fuXLG+Qw8DnVm2IIxL/UPvrK
mn1AM2YyYhDvxVPQQ9CLrZQZ0KnMy4BnjqpvgNZGOUGaH9gHZSLGvyVHmME5x8Y5
dqmS+NgcAHqVGVsYCmPvks/es8Vy+F7fh6IndtTdIv0AyrXwF5X4BAByY8Q65kHD
j0YVh9ivZIZIHrzxZpMOyJws3RmIsOlnu00XW4LIwUCH1D8Lfolvv1XX55P4JA9k
90NOtOT3uXcBBL3bUfLMppITvBkBlaEtcWHLp1wGmp4AiZjDsRF5M7H+xWtzzAm2
Isaa4tmw9KM8xPjYkHVHq8rPxtGJOpDZoIXeJ9e2RwdNGr3KzXGfPkU5EjfdBO/e
vGrrd0/j2f2t5ogAoGe9lwrIjnGBOu2g7xdtC5s9RXEioI6kqywGSOWLR1/d9HFX
Xt5s9eMoc8tf/uwMeEm76fwcTQUuKO35Om3AlayvtqDYcQMq1CZnAgkLTPInwspc
NyIBf/V2csnyLmC12fv+yvW4FuEtilB7Prn+aSWu3dlHdlH0fQ2oDl7u8BEThXpo
QTRpfZSbcGOsn2BR8FBLRIFQIcr8g4qGKkGyhX6mZ5YaWncwTwKXKMWMvsNtSs+/
BuFzW2m8qai+FLtge6LwvpwiDN9JtW6BKZTX790/0E1QxIGGslvjcb9PrD6B6IX5
g7Y5ZxdZyDOsXnC/ITCUuK/ck8h5ZmdgSvon1+hiyjlHIBgi5RZtGA8JFFnaqfs1
foBSROP0ryQDJ6JDnLnzqHnuv6Z6BCigH5N5eGoE9Ut59JGvWt255c5lY9I5AhgB
jC7XieK3ZY7MIy1VXVQC6JbaJsbGyXedjquAvh67TgkbNaYw8Uf/+YI03pq+2BbN
rIQKuiL7DRTyVoOMmyfN1ttTJ9853LGxteowWJ2QYuP4SMeQUSZV6Fo2oVLeMwy1
yuKrSy4z0t+NKZRzJKYfeh/U+gWZndfGPhG85BsAeVkuTNbT/j9neuhI8Eovf2xK
yLdyOAp17tzVqQ/PSspry3jPNbkWArVphwzBctewnOYScqQWRuBr80WUEYK7X1kb
F30ixyeQNSUz2YH3Q0dw6/WYwfC2vvMiu9UfCD4QdTjcJG53mrh6Lyik/jSzWLM8
TaIWHRieu20BZVHpv3cOOgFqPxc61Ey9Ys4wUvu8e2aXYN7EejVRgmE8DR50JqOe
2yp5xtEv88xdUfQsxwTS47DLPPfd3FjXephPyZzIOVpmiICuGZ8cu4nzM1swtyMb
yPvR9U+ukpDRpyRZhko/KvHBvoA7xz5s+G6XArVJw8QW9RZe4s18PHLJQ86d1RaU
gjgLxHmWBGAmDFk61zNhXwA+U+Y/sSYhF8H0lr74PRKkzEbJppzDsybgqezE8kCU
kC4a0VJimshaLYhJXlDkxi1ljaVEhmt9+6vRzHXLGen5FoSTSsneoQ2C6wu0NP0y
UeSRGOzKNSfycdRkp7wkB8qiaYkitCWvdmug0gsEXk0bCOYGdo1uy63orv+LETEY
9ImfA8CkICTxgnFpJMFPkz4kBKnrcxuIgJOC+Or1K/dI94TomWnFqb3t63zEBAPC
d7rOGmo6KnSFdj9jTzFOYJbsi6BL9jJ5EHWsF6JwWd6swWQIHZ/gfR2I38/YNKiV
EKdvCr6896k4WuzID4o4S1Eawg9eeUsYGzfj+n3qnxoU2xhONWvjUrEOGJv3VJDR
axsZUXLqTqZ2h/9izzGHKrwZsyruwN1nq2maCfzMido4l4MeixVD5ggIo8t9lrQU
dB2qPxI5LLTO5foSitpOVk2zy1LoViCvQXAzz9G/aoF3rc4+sNMcAq5xUE4GzGDx
b9DyMKQzTw+qX0FPqyqHaW7i8Uy2BTXNcElcPk5dkK7HXkaoZory2L2TLtjFGmJj
VnDartj1hpmkocrQPbitLodG/XoS0mhJDHKWamsld5HUD3Ja8x5mvMd4A0yC/WDp
+pTOYvCWaj80yy7wMSWEF/C3WqrZM7Rl/d2GNj+pc9JO1pSKlv5qGfwWxKAvvgM6
ERdBVKkIxTdCqGfcl12+8x4B2TdndCl1A/HYcMxnuJxpoK11rzOCW22ZlJGWBI2W
zkwj4Y3cqyNPmqxDMkvX9LfRNuhPgC/RVVgVrYRZUSquA5qPn1CazWUku6koTkd2
QT+I784hYor1DjNnhLNBDM9FARlKXWuExedKb3FIptbU+hK9KDiM/LVgPvoY2FWL
eDrHJL7ooveSJvuISsbTFaVN+WTA4EeFTj+KVutMUWFxwvOJvaokqnFaR1XP/2jN
IcXdQEmiRsd6WYs3wUlGCN2pQDM+akGYi2OXYkZW59dUV76pKKDd4+qHLE/eKgd5
GMZyzP7SFdnO2uobUxGbOj1Qo7OcR+jTYbA2RiHr8JLJHijBEjKZaeEer4Kb4BeK
jGe07UOlphk50f7aVuLzIGp04qDCiUYpb6/qYfgHphfbJdRU09wHMNKikl6JPsJ1
TuuIO01GE1+3gsCzQe8YaPCDDmxqUmyxKmsUuTvOL+HLVewRZrOuje19d7MsW1Nj
T2R5unpdNT2v5iEG2fa6izoq6YixO+T3eEuSTLH08ziR6x/+7GuJzixm3rAZxRMg
hObxjuaXM3g4vr88H0q7qmlrr18rweoCbyluXd9yf0wcGd3XbG1eAJNw5U9pkFbP
uY2QphGArVsWxk4/yfcmAnXzfFmxczluziOKBNoozIjOInSLcULIxQI1zgungF+Y
Q6MfTO2sZwNwW62PLgpipMPGtRP+92YbUvZhL+I8ahyZZYeV+upDWhxVJhNzwI+l
K3v6iU3SWwCGuFTySjuipl9X7nJErFZAetkmfHGyi4GsflqBkv1bHxgk1cYTUK2J
ImqDGZrMv3TNzMB8ViMHpHi2FCK8PEMHMRpI3OTV1rnkrnpMK6awe1QwmSrtb+Wq
VC9Gh/BlS008JTKWQRzIlLLVGdFzqXZuB+Ay9shajRjkGN28JIicOVnjfvFbRbeX
/xTK/YABKQ8XB9eADwCvL/n00OKakr2stxbBpM9lwQCRmHJ2ddBwl+wMSddxdC+P
ZjxLbq5D+kyzqG0Lhm0sVRSg9dDniv+cnEOVcBVxFTsrC0uycmuxBrdlPnEtHc+u
BGvrl0Go7s3OP0fz0ywcUB4QPLRLCGWDlYstfKfS1cWZqVVEOZ+sIMHcRn70sEq5
aYKyor8qA3JN+qaLwQZh16TDO0Ka1SJzZ66KIigiZY/CiMupcWRhn/WOd0o39K7G
197qUBv9WeMqK3gx7efuf4OE0K9xa77WayI40xvCy9/JTQrzz3PhM/ouVDOnNBJL
sPITxaaC1KZ0BX9tqnr86pW3kl3w5iIy54WP65ROkhPua26+vGftGWeoIZVlfrVR
8joIPJepWI76R2gUcuCWr6l9n3wy2h1BDxQNnGP2P4/BmcayKbJ5s+vXuTp8y713
z6WQQ4FLN9GmnfLeqG6w6hkJxnpQkIk8y4IeNTartUehAw7A3anuA9qCQfIStVMp
6/SCCYTAcnRS/9IfZPgmP+b3vcgOCQvNbS6y7KZ58U+vtJQAVXAOCck+r14Wm8Jn
49Mn0T4qoI53sEBGeLOFy/KLmE03kNcVRgEgmx5QuITMnwHwFhyw0pn+99s7KJDW
u6LpygILQUVT181rnczTUBXXPvtbUrXNKeEGynNU7H5K6zoG+Tk/7GpdevopxK7G
UMHNtsGkS0YLcudsL8r6Q1EDNxXsuDxkk1XZrK7EhI9K62Gnmt7nNCOOleeFl/HH
QqGjBDXX3MNEL/pluvgrLlbtvvlbZd8kIt29mf1ehPKoJU9+vytzSK5wvcLflQd1
KoOaQ6LFl7lAhzk9biZFp7RTYXhal2Y/sQVcO+Fjra6WDd7PHixjK/J/MWoShPFq
9cfUvEcFxsWURlgjQQwtIoHrCmqa6mIUId8/BRun/BlC4m0xDgUNzF1EPFL47l3l
jPGGV9r1I7K3bmQvDzZnYDNfbiBOVZxbS2AjQ6grbvKPZaLupgg2ElFq3YDBFOt6
ceN3ruttY23G9jImNIPuEXE8Gy9V3QeTa3ArVDtBDU4DST09LrEb3AGh/ghqEYTJ
dcjUuvXdyXoyySEiBau8W4W9Q9URieEFWYShMdLy/S6qTdS2U66HJH046wxmOjVD
Ztb29qYL5Zz/5NTB/eKil7qqmihWnINOjfCcdw4IA1CCQBAGPI2uE9dahzLkFP+f
vbhE6sI5R2zBSYddFUSRVBYqQckw5I7q/DTO5jPEKav/jU/gq1+8GORxMfumsoC4
yM6B7xMTJvUisIjkMtp0Sk8TAWc9Hz1TKn8ddeWWEXNgpB7zCuALoXrKyZRWPmyj
pCQASz1oniFIulm16PqoZdCpUL5I06QWtis8p+cATd6i/8e+DeIUcwlgOb4Sel9q
PcUL/mu4m35/PRJLYs8uhmemH70v0Da4nwDR1aJqNt4Yn16OnTRURFm5ICb5Xyu9
ueIyPfQVN1Z4TEfzCuPzh8QfbeWIWbuqEsKKW9L3PWMSLf4RyGdw2h3EiknCuuDa
ispmXVI/suTK7ewYv7p85sF8kKNc15mquU3ZsLXzy0O4Up56gC9ChoJDlW2J/aWt
Bk3CH/4dnhNMUWZ5WoCjqnD619CaRYBkWUCsWl5B3N0PR14/bYL5C0em0b8u4+NL
AxEWLCvRmsNvLslOEhCE1OJj8ebbXFJG7s7ySydwJeVXe0RXuedDsyeRHPhFcxU1
N16QmL/c1VxTEXO7WOiz4CjpieQZIsEpQS09PmLWUvt54OqRDIHIxMlW0PsOSphz
8gEtQYnnaBts/a3xbzZYPKIcuKEeE9SFrmW5F5rPzZWmvW1ulO8dgZWuQHOClFmZ
HxVz08H/baM+anglgxh/u/KfJgv5KRRWDlXJAHbqFNTLJg80K10t1+uE01uyYGpg
i5+6nvlffKvWBP+W8AJAnZuF92P18H3FnQnGgaraF8fLci9E+i7FLobJJEn8IX6Z
ZU7raNvHUqNyH/f5Q7XA/cL0oNVdKE/Qx3+GkiJxSsRfoBC7Gd+E6kC+qw9Ya5CW
FYZTHfKadG+Ue3dZWE+uYT0WGdKtx4+dN+Vi3VjUjbFTpz0vis8Egmwvx+3AggBu
OH4vwMva440kIfUz8R37op68JlKeY7TYPohakEDh20IIGi60u/lceUp00OEsCaU9
jpTYWbqVkjLDTzdhqDBxx5jm+9b5hQhbHnzo2KTFoSOwD6HZ+0v+XQR4M78+gWEB
A+oXwi8x7XIqi5HsVS5akihKQaL9cSdEujtlOBgSyq91roRUXOqG5OSLlEI87xnx
kYmgh75SWpYOKA5YTrXugXbwfijVH9lMApdoUNqNvOJbPgtuzI/+kQ/NDLjr4gA8
aQAGCwLT1d582pesog8a1CN0LxedNCzNV6Eu06nsKzZHeXm22Bzz8WQunFcfo0XU
mC++w4I9zU0H0BFz9w82wINdoEQjXm4rqP7l0EhTkknmK/wL6bv0tkNiUHK0e3pJ
68y2x9MmDK6s0OCi+cwcXAGVenBrdFaiSI+Ur/unT87ieTCmN6gopFsLwnFhakZM
tdjNE90PYo6Hp9SiUt5xk+VcFF6ZKu1IhObGN/7k7RmSIgYVHxWfpXpByGvKRbIa
MdRz4IHah7Tj2nUpAJwAVZO51PAz7QQHQ4kFI64L4RmG9sOArky3hDVlvrPeQSMZ
q7YWjgV18DD2Q/BWG3GjIHRLC20tAUic/gzA1VXzZ4q+NM0k/luv7vr//55qeOnl
vcqw1AboqcHFVPSV0fXgU8PDNXxdwIKpSg5AbrKht9L8KUvgn7CE+sB4tunhCC9t
ALp4zhtnnUHH2ypdPkmKLM1Nn6Y6p3RAdwjfCbsY0bKYKDOIvsSBJkQ94agKPiMj
l7K1s4vH7zy5AGavqB6mheajBc2Z+9eFJDhi/qKm+Jl949cidYsJFvZZcl5AmSve
duSa0AAll5wd2/ww8HeTHQns8ctVIWsKZQiX3OfKzfRxoOvVzWsXEMS5vPjmBF7x
NgnhoIWyucGgfarUFxEcqT+2ZByu+M+xSc72ZLXN/kL33THGFZ6tzlbRGQJYcyeW
eEVkvDk8ZHXN+CDVcFxRbE3yBmpmUUFRb7OGt3yZtSMs9iRB5i1MmN6BRSaMlN2N
liVwdndVI6G1TP7nMjXSjn+pNoMW7kHilwDng/N0EkujAWq6RiqUHWfOoT4mvi51
u6Ds7zi2af7CFeIZvS0CYh2xtYMbtlnDHRvyv4nHgX3dnvxNQ5w0ij7W4plu3QOq
8QickOOViFUKzUoEDDyGyefujlN5f00gKW55ZvNJ6O9olzuxmYqnwourelvpjnWM
iRzPWtV7E96rOvuW8aIdEDy0WqjIc1/EeXyfI3ZYkdSOyjOY6ckW4KvjC5ojKxpb
VKHPox35un659SBMB6dR3rsw2S4a0mq3oRNmxV+HaXvClZOywBexFV0NRtomclAo
EE6OcJEIhbNb9WYO0o+jKQ9YQqhJAi5QZ44MNNzqjKa4Lm4LHtiKMR8m6hS5pikw
0NNW+26S0RWzNvgOS2E6oBg50rFPp889dExOdNSq84zB6D5NlnHcYnXnWV13Mk9F
ARZBqAbMNWPoE7vdyvpsDQjSZRYRabGjColXsEOIiPvUz2c+VSJxYCcCgL24uauj
/R+1o72fwg+c/6y4sDZVY/CM3NvDjJakrCJkd9cx6vKL3TEd44MiB9968jmDRFLY
vJ3bFj4jUFfLJqTZ4HJ7cEA+LFDhAnTyc1hGYb9swSjlO0hKGFy9TolbTGsEp0hy
Oql1kw+IwyB5lDQZTD1W8Moxtu6wWygryY3S205ftrCn32iO0GR4y3VlBIq2XB/d
wjSIhfNOCxk6yTcMdrokSZef6ATHBfK028VUEJi5dtsDF2EjEvdO3mNPCgwJCsCh
xGlq3LNtAAsV6L5sQqDaNlbuZu3XVGQ4fRCxb46ky0ZFW7HLd5i4K4T+v2+IyS01
yzfsnBmEsA6U3VX2KL1yPpCFJg4Gg9VFBKfT1Guyvl1O4C1QnPf3pwLc0eIvKW33
sWalB9pHFXMsSFL5iPTX+aZ5EX89QgMDF9SLDxZiZIBijA2juaD0/sG/B95RDe1z
BThxr0c1b/T5fx5f+BmbAbouog5Z2q3ymir50ha4cildoXUxQ9dyx8NVSajAF9RY
zMUwWXqyAuNC9UEX1D0mxn3lo4IW1fyodp0DSxYXIGFcgjSY9J+RiSgQFKNukRgU
uPo28gxGi7sACz4tP1UfMqlHqvJFwONkHrF9CagOcZNi2N7awMBYfGfR92yALXRq
vkqgrhf25ISfrf6JiEps78Rh2lqiy2ls33odxXi5Ui3Yp9BTuIKF+0XQsn1zuczE
EOt5iu9Mg6rBu6HHPNe/PIlCnhnwtorNbwET/Z6jPjNYJ568CYrHWGQMKFRS+/Lw
gh66JTeTXoLBJRX/Fm5hR8scpsqFpuGmJaHHyduVrGg/i57gLgy9M6dpAMbx2Z+7
ksHdTu/DcYJlqyOUAbzkSdJmlDrUoCr4yk8cxgdzckBuMRZ1xD7syANs6hbSg2Pq
g2lJlSdPZ33jNdKGGLcOOz/LPfWW7CpOn/1GwOCcmpxD8XP8UrPv3H/nUw1dyH4B
uzYd8BnenoTgT5Uu3UQc5OHXUWDzCckhCrBbmAj8SHsCp5hXdDyu2tZ2lMAnzSDX
RmllgQFNbRmdnCODSpZZrb9sNOrbf7AXSc9Rt9R9VRl5K0l/d9LcFRJKZtRyY43R
gBMcAZUJn8+XR4jPUwgtPXumKXTBJumf9L0tarbvuoXskTRo5OX1XO9VfBqA0zAX
HjpDDJFxrzktuqjOvZ6oUoa4GyIl8McL5lNcyKBp5f4BdAXoKxR1d8WjGEr5W0q4
VUAhGFpZkdlyYpDSDju3y9hZL9P2lHgPUpwLrr6J6tHTPfPTNHME2o2B/pPYjjt4
aPH4Ez4SVuc+NqUj3IvTKGSyxFDgpC6MMemkbeMO5pkv316qUs3Hn2SIj9XteK9v
wtlX0ZJL60bY/QxACAFOnlr7upG2VZGsvA8SuPgQ6P8Jh7AjRx3IJYIjBSWIDWuN
MsWIhwTAB6tS4ONbC2UBF+ZfF++SUBBa3rUxALLhJrIze7E+MJtxns6ZOCZcU30E
84HYzed/wJ7rHvuiQY+uu5tvWWOpZKbD/Pb4nS5CAUqVp6ERR0pe2y0FhYxKimkI
EoTT5D7u9MUaJ/8i70f235CH1Dpg/n5Q+LtzjrDOwGEbK8UyeFAONqP0gQFfAWVd
DU8cft6gM59DoNct86QqctSGm1HrReuhmB9Ejj7FjullxQW6Rs+Kkss1pgG5MiFp
mTLHTccvYbgdCPDWHk5loaepAT42zPUfNA1byUWAsHu6mcHwn7llLdaXE7qpO3gt
KXWLqeehasnjGxsV6xMwB/hQVKbjCB6fTVnOBQ1vHn9+55L5lVCtI+CMdDf+/0qX
mLcCb8A+ZOLp+VMXhIj3GOhetccnV2TLTsCyuPL8kwlZAIIQPFto3XmkpdPNkFKB
hK9NptJvmOLwcqigx3LZb+ErphmSA4pSCDKi1ppXVnbDQ4kq0CZzSDQ+yTsYQlsF
7XMV0NBrD86mtfXf6mFQWCOyUp89BdEKXqjWDzBAnpO0DcLflswcGBBSzihrGzoV
Uq/+/+MZ+Ja3JIeQ5owbC0HHfJer6lZrnSFT7Vld49MiPTR+9lmHFdLRS2UiDGn8
hnsYRobk6fRUCAzT4YVPgmx7x/ipEpQFWeqfAJ6oy6jhLxABKEjxGOz1D/Qwkd0Q
Gcb21xFAhXHBEbCu4/YRDbPPGhp+WTHmbNL70Z76eL9Xiyiadh/eaeSTEVtj1a62
YyKPandsdG70lLeNm9ESGpppE5lMPAazwPx6LHDSNP0i0MAaDa+T0D/Dntgl72vy
El6RCKUbj/OnS41mAmhUT4u0Lafll7Ox9RkKSZeOu2MFFSDh4D+QjF8uQIKEigWI
jzkpfoZ6QJyOnB0d2GaFwMjAfR+O153BvmShJfyvPPr+7zFlOYXGumVw0zZy7Zya
L3rYUbGYX6ukWLah1uQC6EGyUNAEWloIeQKef1/QV4eZZPZn7RqQ6FLYZq+7bIX0
46q0aTJStZ45E09iEAMm9300LMX+IuDOMaGBtHxmCZM6AARdX5GkxK/aPfvaZH9q
3jFrmtiRS6btBrMYKX5nyWUnetsA66u6z9FFhJKa4144blvLaTq+sQYdE7zK4rLj
ly9XywEmsj1IYJLlhCcKDCL80PxnEBOl3zKD50dN9w60onlcc6YkOW6yHGASoGWp
uu8wZpwS9DjXwGtywrw+FA21hF1cKt3N0doGXTZB6tHuoGD3742tRR6quxxoLRJn
lKwtOBNBP6fWnpZdcBqlIV5LX6d06TgiLV2NHZFkFSPA95JeIfgTfwuCNsH4MFj8
EkdpoSvWZKkv7AfFAsJc/Pma293Z4gCmA+XhByssLQHVaimhu4S/djW16Rfw/pzP
Mq+WRx62KwVLHeboXt/NBn1EN7C0DK660dd2aiLeOC1VtrgmiyuC18TECcJ+e1wH
goBAKphj6KR2ZtMB+uV/m5Pt4N2SY+q3ZG61/b+ZFGG91TZMBQpdFK4t9VDiUcol
BFJQeFqhODpY5zMZ37LKar4LUU37oR5nf+80cPfJyDdM874blguaUO4aAHJjs/kT
hLAgP1vqF4CMfB3FHnXW5Epgu5MG0LDRlyW/60D7kNpK1HZl7WaUAZIy/WvK+vZo
L4HeofC49RdyST12RHiTDY0SFoMdGwrammKvxJPkSEWGAQV6F0gqagbHEs0Oxu+Z
Di3iSdW+kr5D0EKjd5u25qfyLcdgGszwlbBx7a29LgQEGUuufFs9wMC3B3zw/LF1
X6doAT6b9TyMd5tJ8hqwlUDUCVhe2pse5SDtQC+mORyl62blHHE5av2PF/YlHD22
ZZMv68qUynXueb5ib2ftWBFz5x1B7ezkcGmpd+dxeuagORmKVPZ/ZXomFEW0LyYC
GYSRyspAOk8JglGV0Etv6InYQ/mE7nlFi0AdxmHc8KxHVr4QDDgLJn/jiicLjjTc
cxAk6fIOOd47D2fovIm5fyjjIiZNwgrlww4NY1LRHQoRfyxAs1cPiWpMg1r6owQq
nWmG+euLfHMx+nRZTnHpX2rprhp2Mt5IeIH+gLNSVAizMbb9Dr0BTqP8ER8y/Oxl
agMVJwmSqBY90AzpU4ZxihXi7n9wa6jmj2XbG7sD0ozgLc19l0CkDNSIYDfIu8TU
cdYlCZ6mpeZEWN+nnKHfKx4TvoKcI6sG3YYthxMMqpq/r8ZJiMLdC6Ac3R8SEaL3
QMHqWP6p3B/t65vB+WdLIvmRq284scqlSVlJoJjT30FowT4c51sMl/zEIhbTXIOA
9tyL3vQhvu5JET2mynIpJTU3W/qj57dnD7XqVacCD+3izNYkPegsLegB3XZUIT2f
hqr1tNCw+2QVHcAhNLFFxsHUcMm41t4kjFpnz3g4toiNFzp7oBkijCKvTAfptvMK
NUOWlUIN5YTwUrFwGRVqgCWMxCayiRuC4cnkljV/BoY21O/Qo2p9oDmPGlqM+NSg
9ScVMTbX3w6BDOG1iFYL6q2zKLY8tc0QIbZE8en90Z6WF9L7F43+RY6+g6/r1tNM
dSuJkN0ZRGHXNcQ75Kpnyd7OMuaDLlrCUnndnTFkiGRbr/D++iDOWKMOIwcTDPct
86vI8LLxKz9tw6uewmANriwnQFoo8H5+klnLMQNM9NCTp/kT1iZdiN2CKZOz7Zeh
3m816AP+ZJrZ7tXSzwL1n1utppjPdA/KqofbzDhBhik8z4paygORSuJnPwyeu5Fb
N9sqX9jfTnXb+i82WVvUxD/0vpb3WX0vWEijCtWO4Yylh0N+H4z1sv7DPOat9HsN
IEkV4iSwCXap7C6DcsaEnGEbgd2KD+nqfuDwrbgfgZoaaFbWX1Ib8sEPn8JO82g9
MuGVIcegLWgOc7EghNlqL7xq4C1+/yHrJvkdHNIiQXBrz5ZuveXXl7zt1symnXTU
BkO8j6gNVIetqscw2riOdL+tKj+1GvjWisU6Bp0iQWRjv/K30NMhbbfpVM9tP/xf
WmprTf8KAYv/dXDHC+v9walgU7Ce4F2Qvk6ec1jt9E3BhPO16X04XgPBr/QSRpA4
QVBr+cbbXoADEoIk+RJbn2UFVtOjeJyCssN/Q8IzN2f8CZRMkyB3KeGHEJskcPAC
Sz8o0nyqI7XQROz3M49a9hrILZ9AaMRRHLxYyavVbiVCi8HE7H3LffyNX/Bt2Mdl
Q4cbTlf6sJ03tUZ67zSvFsx6JQPZdk/VZ2f3BrdqI6W/Qf5ZAssjCxJBvu3U45y0
2KxpZ5sVkahMT2OgowfACsz1ypFvO+pMWTZodsZztVFijfqfIOP4Zystk6CxzYKi
g4KW5QBitR8EmYf3gMPE2ZSLX5pH1nrvmBRyJhyV/7+3bPzpPfWv1OT289Wiq41h
hD/xwIGz1u3bCTJbPLaHRcek44Uv4/ph4li98MOKAi8nfBKNHncF66rIrID26IW2
8+ef9ExJetsWqjOy1bg6bVpgscWqbjakThAceR0QzuDnzqFEstO5crfJ8Zyh4q+8
HgbiIRqr9AcXELL5E67gwmjSnyWq+5ufl5haQ2IGni2r8r8L+lYG1LpZOj8HAt6o
yotwzr/MoLw/qNvhK+vLjuiTSRUdyjnWaaob7atdqt6X+qCdZD1BcB0oBKwJ5HeB
4fEu0CejcscEjxLY2YGF55rqynLexVPLZr/e9BzBuUtarHt44lHeYvj/9iosylkb
cqqPWiopGTv9gEk2O/TOi5Gq/rMDb2E1fzkinEiUcmlX+hrgtvgbQ2NCSzVsm8Zs
NKRv0LT4XEKKJPWW7qSxUjaBy8XgUGi5rOv+gyuGXOjYvftuTTMh1b8tMv2zjD69
ztUrIAbk6PL7nEY8imxWC4RuNwaq7yQKTI3bo5dVGE6D9FfnK9S2KHUEc0BK7S/d
15milj03OI3gl7PSygQFcC6sfBaXH6cl+GAbj+HKcKUGZKxzcg8zHFo4P6DlwxeT
qfHW44IaSCCnhxRUiwXVGKizXPgauntzmYA8D6ZnsMH/NnFFczaFwRFpQb6ikfSq
Z3s7+u3L5wP2awY3SvghIE+hm77xxRtjbcqztcpgmEPJaysH0HYjJz5DzyvaeStb
WivJK6fwZ3phvCuy1KpWkANn+6B2LqIS337BlhfY400aCBQfplFiCOuoLM3i4VO7
rVYIIqaizxjl58wkF3Rvdvyt1HXDPQexPJ1nn58tgCleyVRxgpgA0/vHQhGlVI/r
zfdUm2CP9c1IK5KLskBfuScyhRW97rRH33I0Ud+7jC/+GRkeDOG8eLax/k2Btd1w
BEM0+fTeZOXU8B3HxtbT2U9VrELl1AaAxCybctNy7n0lMet22c/MEY2c5AfIxSER
JYUwPBYrQnUHL5vVaxeyx84rUQIplP/+ZB/+8+gA1OgZOvqnKxMm5FvQlB1u/fsi
mwIGCO7lTHOsXVhMgBuSB7kSgJxmtk8gQHkdwj8sPRmvCed2w864lzJG3pyZ83EQ
db6hqlIj50EiIE6MK3QFXY4VKe/2nxfTPrEQrtfJmt76M52fy7n4i7bxHM09QF6C
R1jEpB2KRuxuVPqbBqKsRGt9XQhsvrZP4uxJU5vrOWLP/jlf3axR2g+id/jlrt07
9FRYGPKOnTrgbe1vqE+ugOhpinOcktd9sANb1V0N1S4H1bIjBFIvaBylYzdNAkhY
v8DmrMFonP+U1aFNS1h1J8ibQG1I6CH7jsM3mW0UNRUMJQe5PXo0KBWi5yi2NlTQ
bIqsuECFRMbNE29z7YqtnQi3ep3R9SLN+n+IkF3gT9V+f/8JQaErLviH5qP386Le
h1KWrMDdRmWCU1800h+co93dKQfwgy4kDRMH5SIiGv/cIBCYrmpGnCrbYx21wqBT
VYFJkFcJ9P3CqPqUYO6VKrIaODPhgS+dwjAnsqOMZcBRnHpE1cKb1GjAGSQpDi6D
8bA+3qXZ9NPKqzrWjeelk6HaKdXdd8cYOVgbyMy0pyomi9cy3KbJv7XRMb+n2l+t
fFUvQBpA64FGWRxmy2ZxzZFmAKGa3MQtRfUIa901LVKXORV3eenKwfkHQS7XsrrP
ZuucCSCjXB++ric8RGihP09n51Ie1bLUCattojfrE1cJoi5LYykP9HvP4uMJjR2F
gUbntPgfdj0VmYZcm3W0ISouovKEZ4jwTOAylzNHBMI8f1r32rf10BbqgiWBoaPp
dAAndPHFxOq1ngx4pzUxZFmsYxXhKY6D/MA4wysV9srk2eBVX4SFrFnHIt/mhnGu
5TH9LS6GWVTDTakVRv7g+0Dx9SCtr8lOltEnphFdLo67/ZsB+tVxNcLTTK6ABVay
8cfjKQCB35kxT9zTNp8a/CtE6IoD/CTkczDQkf5MSMZh4s3MOt286ChjOHX48mCP
BEKwPw4IIzeuwlL8Pl/glM2uwId7kPcwOul7LjO1e4lOoAXUXTqD2zW3xy46Iv2m
lP0G4p7YnpBcWn3U0pFMFvBJgXxQHOmwpom27oYICtJHmCo35UN+HKcBUTAhI/z+
rE+x4VqUwRMKuxLy/z5yGJ32NCW+PExdugtGHPPoewuWKtJKvleQDZ8lRzIgx0Bf
ypW49C/6NNSiFpMwOfsapCsZmy32+XLf7FY4Ca/vuIhRpmsfOopTmiSQho9ZUrTp
fmHetC2dpsqdkA1JmdZlNurIm9W9oVfLzGivzWUAPBQVDjqrNE4zeXAnqxU20WOh
gOLapU8VRBWGvxo5rZ4bxF4aPmYz4cc6tIOyPiyUXjMgQkLEIw5AsR+E/HLxwWF8
8e7FyhLwbqkoRWgLVW3UmqRQh8w5uNP6LicJuaWge9tM/0OypTbThmwLCMoZYjqO
ObQhXW2pQgh2t6aQsl6yFi5+Epr/Jg+sByx24reiUdMp7jRJgohUQ/z3akrxfREs
qL4ympoyGt0DYDeRmpeKaHNphVKRjMNrRyg7b7ZFjMQbl/3mV8uHPE8xatHgVcdI
X3N36F8Z6S8Hljns28/eQa0LMgbWHznDUBuN+nFxsydIpLs7HDAjdHjoUMZ0un4f
JY8zms3sAoDsrwDOO3arPlXHot6A6iRYCDcrCjaoSc5c0lsxQXMPPvjjW8oU/3BQ
7k/Iu2FCgCPdYQLWeBzTsCYOBWqYEEMQN2h3m6c0D1kSvvFaOYWHy7CImRfklurW
0AGI3Qp2Z4dnKeoHb4QrgKWN88FEK+ZG9k9iL6el+Ekbwha5e/4rHXiAuVFhwhEl
S5CcXcSCC00qLtCndzss60J055qIGFsAqR4O1JiNBZMeWl24Kh4rwmhWasuG9nty
IY25j6aolWaR5qUkUB8HDlU+vjyH3A7W+mDjXN1cS1uoo/YF/pqKpdWFwc+rrM56
5zE6ey0F0pFZX1VDTx36ZYEm8P9aTRd6U32Uj6Kn8AmeoQBhfy0gzeKpaN3Ua0xC
LM2zQurVN/stN/u667uOGZNA8S/U2N8kev+RXwXyENjXVZ1+XOIIFuaMabgosMBa
N4O4uOjvv+kH1MlOzoaY6wXbH9EOl766lG1Q9+Zya5wgA5sFCxAAZo23f584crmB
nX0Gp/OdwWJfhDqRc2Xi7o/aRpS5Gh5accFt4OTFSdWBWK/R99pPLZdW6APBVN10
cI3jWKFMoVHYGSgdanDHFmfKmXbuIQZAiXMxQJCbdsnAaVnwTT8Xw3dsjO4gHWHa
0KS6nku/4HYA0J6Qd0pqhHXpn0rBAsxto3bPRWPkXqB8HwWCieLOLJbeY4WQd6IZ
o5inlXwhXTz+ibb/mKaOYruSJd2EU2WOqlEavxVhGgAJYQtD3WAnitm0IhHXeRf4
Qm+MtXJo7fl7LLBe4LCh+yV4vfl9XnSoFmlkRPzUm1YskduN8nXXPwCbLmaxYhRx
aKzZX2Ucuc8w25K8jxn7YDM2ruIs7DxtR2tJR6NCpu+Ed2FiTbJBG3FKAuPnpKAe
1iXzkbEpwA7cGCZ1+th+ZYUeVhE6k2JcrrgR76DY8g0V+X1lwCyBePwCKNg26Qjk
D6So3gX3h1O9YpFvFxzEscexsNNAzNtrGG11mRuVbbEZHy8tlAyohbh9ZGR7c+C4
8c0WrYmylhQFeIY1pSZVNl7w2v1MBLjcNepeDdMgy0QSgORoW/Qbel9EykRSnjKo
7z0eYWuxcdoLc3mLPwiFb4NMTfrXCDI4ypUaApN4Be6GlhDNmVaT6jCihl0o4cEk
/xHNqL4eb4JtJUvEILyq2wwF7tWVy2Pzti3gbmcsp4vTwSADKVILkES0iueGDFOm
5Ivu9NmyY539l8FJiG+STvqkLhxShmHHkj/mEQvNsCseoGvIvaxM0Y8q+V/cZdLf
TcFK1uAHJnMdPBDjpiNtzuYccr3QgccgrSYIVDhdJAgYqrStWj+lJ+hITf2Tm0RP
fC9MleX7WswCnCu42+ozHPXhdxmlxc+uR1T82erYRYsHHQcxYYct7WKXPakT1b3W
4chixSxfu48Yq3zzugDV0s1LOuZbAUkJAcn4d90VjRj5sfqEUVm0UsupHSRAOYQN
YrRbV6+xispD8jiIx0uICEHK+wd7RmpkxFfIK0W3GAUXbevZTbQuvXVjJFAGeAG5
RhF1YvmF1d7qAzd03NBqQfbZ1KLLHMJQFRcEJO+5VLNiiXAc9bz6pmlZK34lZ2QZ
nYKkU9YRBm+GydQCp3ijBYFTHEkGw13uUGomsszhCmDutRbZ1HR+/Q7DQuHRxWZ3
NzcCe/pUysbpGWM+1cFGI2SAnwSCHnWars/4JiYWiWrOFCCIrwrz9nMq3MEHPjA3
v+PQwdYLnOLc9i2wvQRWnuuyKt22IasgL79vzEnYBYo1cx3YjFNOZ/rdDyitjGIW
LkfNA+1rrNvqCRvBxbr0SMdVYGgJhcfBtopnFXFlOVqjpjcvf2tIrHr+MUcoTwaB
aUey2wCE5eGhWbhrfCIcmR3zHFF/EjlJqhmTKafU9wd5Ua+BQzOGRo6pc0Go9pku
94FvcvbalZaxFVJmIzRnfYSdFehJ4ZDHU29xXKlAiSC9C8ni1Btl0/KYO0VtwJXj
ziKeSnGY2ZRdJCCDMRykUA9IkHLcexyaNERXfBddOM22zNGfZ6WNVEcdWTGOFSxe
p1tIRfq/Cxs0HC1ZDt/bN2jqJ2mFaSc/S3oiXu5SB3JsGQNXn2blcdXQKXyrIWpr
y4dnh3ByqrVZUJHCs23m19RiwsQDwRB6OJVe5lV6TnZXRMwcPF7hxlivZxdCaHGN
JT8b26Z5guEJ3abHF9Ip1oScWT5uGJLN0HbE/Brq94JaRKNGxMYR+z2IUyaqp5HN
sqHH0m65mePb5BSviODiupFmrfC2MLidQH6GV6kcQG/wEKptqW+6bm0i6HMnFmGR
I0InwPEbTnJs+YGhT6sSir8hlOB7EMijphtClKH/VmGhxMS0gZh6C+jRIHYI1jPT
NhK9TWHJvxQOzDSE2qI5lNBN9Ujm5fNwum4F+XWqGf6Hrzd14ruWdARHvTi3qavi
fBcHToFIF1rk65SFi3/C/XHcSHi9iGKfyW+eAy1EqyaW+sgeXj/wo0wykDX5Vbhj
yVZzW55jUvyUZ447zVX8rXOGmfLZcG7rpW9kQQtelL6Vtaz+qNnKIXbflyZCPIIE
dvWpZ18Va5QjvFQ/6G6re9sIHnB3qcglILRPAVPyTJN8M13lHTEMTrC991WCmtJe
ip9bVublngpscblcqnPxr6fmBA884IConPetlad5Ephyx4BgRaNddVil8Uu1IGmW
FQ8k/INmOmvBLI9RaYt8R0n0DWWqtYBYAg/wcybvOGnk1YU8EvdtUdVS2Cdu/a8N
vj1QzoSY6jtFPIJIaLu2JWteM7fK05cWUZjp77Jrh5JirXoMFOea/XOlVi4WdYaK
9EaaszhvC1yKjctJns+TNvI4fMP5l35DRxnudPlbY7ADG5B2KpXRwpV3Dw+jAxe/
/88mp/OqVm1doA96RfvVccbL5pbmAmMGwYsQTuytuYXeyPwm7avjIgkCdE16dQ19
h0P69k1I1tZk8bJxRIKtCAGGP/pMldhN1r7o5jGKsDAnsHnSeUI/lZwR3pEHCu7n
WmeEKZTJ6XeI/RzLRQZ4m9yp/P9nerrCiwnbh70YrDYZyZQ26he4HxvklQUPdb/T
6wVcYA/f9m62nZzcfrbwigScQ8paL8dW6RQ7zSB/P9HiLelgsEn4ZLUWPRJPqGGM
eHBlXc2pFq5abqlJ330XB6ifotYgdxI8R8/xNP+7A+1UmNgYZQmnC9y85K4JbuEm
wJBo0hQL2ToatCs5J0R7Y9bAB6M3nRXgcTqEzrWG1MEhwua5bLM6/mTQS9JbIb83
AoO+2x4E2CFBjbnc7nh0nMsNHkCnByXvELjBGyWn+s/phoiy3b2Z2xk42eWto5sw
4GRgIsEawaOAnlmOTrP5vrE99D7EF5LX14pRHe27XY3PPEqlwWvCxLrhwSozLKVQ
YiHvykV4T3u+0ss2A7aO3pnx8K8GRFULQvWxKgeQQ6Uu5Dd7PTZxujqUfxpI03g9
jAl40KgLiOAHkqcndYjq1MtHlnJcS5drFrev5c4+6b7RaRWY392Y0XSRbcEk4TbF
CltEXANCjXM3nb5CHKu88axIYjgL77pz0N2XIonR7RfMB8MD2siuM+39NuSbNH7V
XEtZdorVsciLMDL1N4zZR3I0rkDIZgea7pKKClIM2ekf7ntg5affZx/XmMQc2b06
lM/uQbNW9V52qYIGoYlVpbQXnnjrU3+PPGtbPiAy1YmMguli5XpMaP0NfTq6jWPe
9m+vfUfY9LWaqCIpSWnw+FbbvGkl//++QthKBqd2xSIj1VB4WtOj1EDAvS8MLgY6
ZqcHhzVB8EkV6Z2+Lo9WW4K+m5+99I5pHcwo++lugcxnwfSdnA8HzecsinV3eNzs
PBHzE4fsLZmoBRWM8FjzuNZe+TB5Y6ilwrEOztcO9+hGw4jVk1vIO/fpYgh7H4eI
MTcSlpgGvihkrH3PgG0ZXdelY98pFnXbHh0Gt7zWr6/TLtpt3AKcY2fYarlUf3PG
7s2yKNojxArKwzUEuSz6EBW/HLMIsjoD6f51eMo2ykpBC3c2+Z/iCvMuOPIFho7D
A/2pJKg9OZI7d5VhHxyA654fvHORs25tsf11V9r7/7PmUpURoicB7mwHDJq1ReFg
BZVDqkpYaZRfJ6NAYyeCDG+R03NY1zhlc9hw3EU3LeFNEZfZZg4ef+cVWjsveJjP
fzkjIjtaKGUXGtXiX8OynYgeT6t+l4Why9pWxMTi47Qa3OCv0d5XDgM/bXAZ6Ee1
f1EGxBlA+/TF6bJTrw5kGCA7hJHwWH9V/cEkoO5Prkwx/UFOC8rWoAROlhiDRoU/
vg1Ioxou64jPPRnMvIgKxNOzO/eHxV9rFHf/dHNGZCEuyWNTQ7gl8YnZ0mv/9VLR
fUNR9EKqFVycZH6L4S/usImD4t8vMzMb+IhK7zeQeBDcR6rbUaeX2W3rsFNbfjHg
7Jn6VgW/RXIZ0AYzAB4ekR5g6BXGy5m91d8atmRkchwYwngu950ogwJIypDwg7MI
nFV4ML6iFx6zl2QWtSmHWpEKbNJArCC+ij/znK1F/Aqy0qKIe7a8MrCVVT4cmYiG
ASiCKRSMpNhU8nwBCJemYgcI3wGtIgviU1e80qdCND8WJCI4LCwC8shjIpJAEycW
soy+E7t2xgmJgRKKU0SaCz6IivgrdoADmV0HFnsvhfQvgXyVLgaEda5CyxE2z5u6
yMALQ8yZj/QlQfXhokMA92nRFs/cp/cvSzkj5+kO/BtmvZP+GS+dD8T5nP9duiDb
t7Nq1A2MgKUOv1vLk0LutZEg1T7SVYQO0TvwzQSF6V8nPjSukP9mhufzW+tPczGy
P5PU4F7WNscqUQC/RVZ62/8Ies33GsWl4IVmRZYLcn4D7PgPndeIfpfjvEtljxDM
c5h5vqX/3wSFe4IC+lco2qHnX72E1JVnxNft5ajHvWgzYPipVTRymnUarXVMWRG9
Ixn18+Sj3e4kLl5coc/UNfLIClIB+GxLrXBHiiUMDmQkoi9liBsxfp/f6T9yCzzQ
WgwyJ24Jsex+A3KazMLjvT4G3lllEa8Vpe7MBtZGo9HkGlQQTkfLRrrOry5/xHiY
6EuSLTcVlcjKEAcbyEfVGIC+q63QhLqJAWl3lXzJ89xGufTUrO6u2PK7iKlzLM/Y
iUQzmRWowOpphvye4JrG0si8+nqDpc1w7Zgc0x8LYrKvLRgLUZWkIfy99igbRgnA
UzSrJhRFCQYSCjr+v90HvG0FWjPeDDIPdxa8meTMEmBRETLwarsIUzYFTJL+AHLJ
25mwpUbmPvnAzSi3BVCS2gfil/0H4kJ7CuME4iNIvPr1wrXDPqs+LSEPlbh61dks
OZdeQM/eZwBsVAPqqDW3EZZjJbF1v93RUGoHR/iKY3poQkfx3gs0xxM1fTLFTGv7
4pi19UCnxj9dzx6rHTv9/vnsha/8B3do+qmy63XEYYAlRwZJLcWcf7Ix408GDuJw
5bUjxpfJOCY+uwQsJpAxqYlSeiu3LxOqgYgshJBjXhVQPeS52mmNQMH+6vYFNXFE
qrmN7VFxdvIooc/FWk3ljEO9cLIThDKd+53Juz+nlmnhopKjgtOrioDhGO4HypwZ
BBSYz+hscdiTXPO+k7pr5dO6p0nyCGtOU3eK2hYmHGgxeVzmM3L1ACAWLqzQDSDD
GjDNqXfOPVRsj6gRbsqvjYHgak/ZL733mgROC8H/EJDU4iMwgwdNbayky/IOTDYT
T4wOjzvad+MVYNlzwi0W0weCVTBYIhrjj4taVcVj4mYcsdwHBEDfXYi4zdvD0Hkc
eigee9be37FiGQg3dFeILw9aftQmcJPkgAnvDiT+5FkzPjCEYV9hkY1bnU5I0UtW
ux5qQ/IIZVvHWK/XxRWkJ004ceJDh8qUVgj5Ssi3ljxZkTL1VSKf2tbGuyMk7GQX
mBVUjeGr61QMjbcF557IajZGaXHaDvdIawPMi0fr0IO8hBynAwqbCYRlSy2WD/et
NOkVZrV0L2n0q4nSlKCnHdBqFEmopR34tP7NwD/YAyqTr12oEhdRSGYUTIK3ySCr
2kR2bqZcvU/haB1+VRj4uohbtlngTC9D1Tf0LPfVdJqMKHDJni+dNF/3evI1tZhP
Ywa2YUGL959fXxe/+tNanUHZi3KzMrA9mWqKlzvseXN9yxW6gtaBsAWZuf0dfNVa
scdmCu3yXqK1jKqpiaBlMUz8dDpM/40Ruz0LiXicROV1j/V8AMBG8ENLnNWXjXLs
k/+FmZMEs/WeKogbuNCeFufTh0+SR+EebN+qdsVYq5UkP9dvLi2hS6a+ODOmLG3e
db5wSqhw8ClC9rPg7GwYmtCpjocr1xYw2023B7rzdcUAjycUX553MCDjBjbq+v8X
yeGcmIxxiZHxKOnSrTPYn5z/MpMgEYWYe1bKmzjMI7VQuD8Zhk9+j/UxlSneb7Ti
uyNuV6vSp6VKCFdVm5lBDOP3p6q0LZwE+W1q/eWBXX2gkqXMSBri50VfV6zyGh3q
s2xNgEcOguZszoozTbgsf0OtQvmR7ltYDIe1VzInCnvxQ3nPvkC6Xgef/7aGb7y7
B+MojpRdy9trKa7WnZaAo2rEFvrV8XRkVYwTKo4nPtTVaXPA6lmi74qayeaT6sbP
GjOVBVuyq1558Rk382KN4wlY4k0ExSHA2l3BG6M6zRc/AAB37ATatcTfOqvM+3+J
Z7BZN+UHGFCFmd8RoFnqG+9hR0dYax79/5Uy27ESCh9aHmkxcxykKcJG9MJuOPOb
PxEdxhWc/RBZOX/5LuEl56nbeCkLgMBStYgw+opz6lNRTOBXMdn7sojG8n0xvKTZ
1A4ihwoI2MFBRDzngLxFB5ItJr0VAKcP7Eq0LMnzdrNdFQCricYBg58up/P05Vuh
IocDmk0E3C89MXRAHdiHr0Lw4lNUcoG73jDridwTrxpQlfocB/XgzWH5heV7doMa
SyINaRGPgVSOX8+xb854tEE7V5Rqi6a/6smfDFAxclOK+XoANbKnVWRT8sNLUx99
zstfMn3Zs1WENX+7C8Kof9rSmhdJh9PRfxF/I5ZrEdK5r7RnA0qxeaTqmceke7r6
L6W4YvuO+NwJAvqrOiILYTeYf2CMsp8VLFhxwZrpMhoDjVdQpjUInqjkKrCS+CCs
08wQvH6oWbeVuImhh99aeGmnYf1yGg53H8C24fiAtsyUi6OyUOKVEhvu+uOqQ/x7
4QPoUWlzJxWGG/fmo7JduVPNl2dS37Qn/SrnCe8BZqzRciZXg2QOhwizRrCuRZRi
wnP8H3ttHVFtCxM6vPDcYBNYqP9RjzObV2GfDsvIBbL6PaS4IysqJJEOq+SY8t9M
YJ1B7KqlvYnhbSuao2HliDGTnQfH42hZEGEgo+u9bRMJ+02cMKaI5NvOi3Y5+AU0
LkZ/+c9V2t+imrAwhMYx9Jf6nazXyjGWBpaM+N+hPsECJcSvarQ4oZMYXDjsGK3q
5GBIhSlMhTjlRZ56wNbLKnLSsE2kKjAh8S3ebsJiJqe6Vc23j+fuK9Srm/poheZ0
o8wqdTZ64aW9lE7PxRJB/pcrlDw/0Epuffq2mF1gEiKrlJ/QCt+6K115o/sWGH3J
6UKHAzW+7l+zRs/cyzrXyVRWosWm2ZihLuyYiPIJhaHcJJyPSccMmNhNVBa4TLXY
breXCNqxeIvkXV8tbyYN5GT4fBPBCJm5HaedoNqR2wA9iDIQAB0SYmzQbUwDR7Js
/ff4XW2ctI0sDmW/SzLRaa2BSErC+DTXFHMiicKj9ablU2dDOp+wEoBHgEylcrnM
3OMU3AKMqHgnH1fAHVUnhQU0+ljvRYl95ZeA4eb1FYhnIJTL1lx4HriXCh4YJpTX
BDHvvHtCud0p4c6GKtTPT8x0rK1mOpW8gXIzz463KictiJ50WRA+h+EIokrvTFU6
gbhFXODUc03Y5+KyAJlRXPLgZ6S2dDzbGbbdoINj6l2irerbyM1ONj3kGIq9I9n6
QMth4l98DCvBAXfgKnGNwe98vW3M7H2RvjqLiVWzoeSE/RKPqmIXQOJRhg87HAqB
LcFur+VEqTMKVWD8+kBWkWevfCU5SQ4Z6QQCwjsLdAp6zMdAD/Y+hs8H6dp5vSIX
Vi0rckzk+PVnsaz7opOj6YkNBCVfgzMrceLZND/ViBvZAGIKRjwPTSUSv2gxhyUI
Y/v3z6fWZ5vdtDdurzDAwgD0PrZVfNrxBJTe+tLXWVLkzhArXK1XnukA5fTIJFYf
KZWYZiwGw4DwpgM6DvU1y3kUOM45VBfArpx6hg/d+IUUiSL89elwNFs5v09XbeUD
oOCR1xVOqvtKlntdU7LPo5payg5dza28rGa1adxyUVG+C3D93N3P2WWu2fNRYBh5
OqA7SSXtBJlljj8QRHq5VUsm7LxAjpDr5wswB+/3V3TAUeqq7WP7pqyM4d33+k/L
Vb/ipPmn8oL4Qg+y1U5NSjzDLAd3Rkk4Bs9E/jaZL+xIAZOS5k9SATGQiKPBhkr9
Fj2wVDrAdyfGeSnV17Uwto944bkhAGqWFVKwPKD1jz43NhXjWnkcdEXqgacpD6Lk
YpqcyNbF7mRd7gbEBIKMrhbR8pKkZ1RTPhL9Ey9/YK+NB1TJ1V/YRw0aP1hph1Ux
leHTk6mRaYRLJca6XYZ2MgZA8XtOQYOVaaM3P0tj+z5yJsuPPC4JCFPHMkuGRZdu
dG3KDIjtTqXOug/Ptp+MbQ8emNiZ0nEtPxUtDr7gxj4AoNcVoL0yjfNXZX2X4sme
udwzfOEnSrLO0GCHXDI5MkUaWWTXmeqhLW2bvTReXnjtPxCL2OmMu9H1WuTRGdRO
kS4qPs0hYm+B021vZJG7yFQBhesP8kRCdTJL1gdadUL35nbM2dH23wG5Tr+T8N1B
YQhY3CNHZHHg92DHR88i2bdGJeTE8jzKtax8yWm1PAqPx5CEiX2A7dF33V9UgjBY
0+weyH5JxsnejprWl63eSCFQ3FyxHLL6sZE0SdfVpMHsLcMIkr/4IshsCASrCY2e
hmolJrnWlulBVpNGYBV0M80Qp3VX9NvmGIyi0oMiI3n5ZBPLjr4dYRzm6NxS2J2W
uR6bcGB9lr3ZsegnGlAahc1hLPiGiwygR0aOPDmeahLaptIxVCDMmAi1AG8hooSt
U4UdANJc15OS9GhAtYkj/3U5LP0ml1pn2b+P849//tyXblLpTAh9nGIS7dEfeUuC
JD625yiRNOuonKFEXb7kDV7oFOQv7lRvTvZ2a7cukyZyBW5Jd9X1VEmWhSn7RWTA
i+v7o8IAeUA3MCZyvBW4Wnh4HKWESf3SDGIFS+NH+kiVPi77sVjfaCuqFQHluvXr
v8Xr+hhzYexmIu9/AEvcEj+tMJwVVFbeyD0Cy6zG9NZDZUUo95ugjZ0my9zkmj88
mI4STW22eVTiGJfXjSfmZGcM1pDjCf0nxaBq3ShqlXvEM61Z80t+LRSQJJgQWCT4
aFKPmf6O5fFsK7hmlwkUD7jxBEFxAuvCa7vt36sIVJkKXmVyYCeLHKOS9EJoQejj
4OP596qtYRNYEGZ3Knr5/o7egwZNKaDwjlMa3Q1t8QxwmIgz4rFc2naFrB0wY75R
+MLG0oP7nbURC2pbBDWwlZcNHKGrOm9EMVq9dfUOg7PMeF73xWbwFPkiKhcxBbo1
mhZVzPeOau2DCcQol04j9WyJv7b6Sz1R+z99/E3p9GKjrPjVoL5j/eMyavXFNYXI
jcNocN/fx4FBjhPmiTrP9liQt+vjsgkwkl4Jo6ga1bWfWIuoDv8AWS3jgZ3dOJmG
k+qiYfN+ReXhC4NJyH8x7Z93JPBNn8d9DlHpKEaAk77NTWPMrZ8TflfraZ/6KiPM
SQj8HQZrUnzTgM65ic2582fMTYZGX3FuzNwWwxZiLAuskxbSMFG5iGu5brtNBjln
YGhDzhMCcfMNs6P6c//i5XxXjCAsUYw8cZ4rtKNZi/fM+pYNOYbls1r0eHex2vTM
DHB1YsfW0x7WR+M/GSR51KYWx51vCICGAw7rNMH4VnFYivyyeblstqL7pcSYDouM
mSiA13esR72xsfnjCpl2SnI2ZgphDe/PTTDhqAw05/T6K3i++iOpp9fRN2RczKkK
NhEEmbInHBOKpLZf6oKB+X/qJLeK4iNAS0ur3LnwLhNxLTXGp2Q9VeLHe9F4Guso
goH/57QsL/3DJK31g+pSpT/hIFN6TzLwUKdp7JOAF6jsEJYIeejH19SpFFouGmTn
E+huW1xib0gPjKkmFd1YwBCosuQpFgBB6CxPK8++MF7lFQBUHuxnj+Z0If8Ts07K
h4ScJtwUMiIOSAZu05Wjp94EdIdvK3rhS7IBeB8WN40oWJUAnA4uKAC8688DyuEn
kwA97dEB5i1Z4BYRjcrlr+6Ka3CgKVJUxglUdDi4OBFpYH2hfc8ZW80h0QbtXl86
LyuDXuRLoaHpoAXv7kz6UFX4sDqhl8kgwJV+jfAQHN8yLhpe0caWoKYA77N7CHnP
FyCtoAFLmSsughVJA/r/ShsStlKAnILLHNfI0bFn/uXuZmj/yAwkq3Ws3tfEEg2Y
mXRCollZDjkSZFZfRgiTu9/CvoHxED0kNj6+2uYYa48t7efIwk3aVHjOfKQxvC5l
BDPZEdhVPDM+vz71nh6vQosBGnYAwSO19H3NVj900PeToMI1FVtjQqWKIaD/OlF5
hzBWP1Gc3x0g0qDfc7ApfjMfFAEch78YPwEMzCX8soJo678W0DItfrMJV6d1e+rK
hR1Myh+LVWepDsu2txhDDULwlRMIlPyY4dMeKrNUGl94r41MZTK4U/SdFPQtcL5U
y6dk+7GGRpa0edmLpXAABnQhjMBAa2OuVAYtw+rI4dZg6xyl0NH98deFK0/WB3nH
48OARY1ootfNCJAcSHI3WofPgxryRNbJHampyp7GxEgsRWbwpSGiAiLDF7AkCiBJ
KHF1qd6Xa/AawFmhitNVTnBxSMdbAchFGK+ADGR4MCQI1rVkBiXPgyUeovLqR+Fi
EYkMyTnM1UzASdue3SP66p2Ema/ClvDR05+NJyuEW5RJtIeZG7FrDM1rVATOKLFM
O1czt3VmxbEbXVSLU47ET1hUn5EZvlQmSUO/D5Wwd/zPzLh/tBrMqZ11jjLzelhK
3s/6Rc6H9Cab+t8+PeX3G/Hx93FqZAtcfIa/OvyKG/q8zY9G9rCoN9Bk7xPJtncE
eIEfeyEiqNBW5/cXfBENPlTaldRB7FStU2hEtNkuf1JiDKSWlxw7pkL19b8kazIc
h72r04SOu5/R4O35o0jEGQLVBR0+hBr5qRx5TypDRK1FbIjcXb0wFvb7GXjkKwoS
uMNWdjJepZ5WprBOkUQRTBrXM5vpEq0t7Z1oZDk60lr9ln8P4KWhOIFEKFOcqxAZ
zGnfvcpUzq/NhmBPP0GtNhlOCuw8HQNGzdKZ4Ogx2N1FAsMvZSXa6PxImXgxAfqe
c1zvzRj+1Z6aPqWncLfgJHkhqWvma9Dtv0p3Pl9yjxLZO2EYf04XFPnIIkwTZhyp
3W2SEoPe/r/9WBjEBAARd5948ooVhc01lwOLcoXPc8t6piT7oqg6m09iDRKB6oL+
XaanGveiwHiqCsSONpFnebty3zTMkrwFSkIk0VKUOBxXBECwVkNeeZycOWVk1riw
81XRXBRXIYA/MY7Az4RPSubwWHz8czudtXVPnA5mfNGtshYEFxKkV28j1a0GUvTX
dlZkLcBb1d2CwTVCYAUK5lfveQ/7tOKKey+jy3ELO7Me8UddWdtJzJHEctsRIhX/
22qpSalg/pWKnGxMb2kd+qrNPc0mTK28VBnqncStI3+hwvYdd+WOV2P1iriR+LdI
DY4cCDqJSR2LI91iUMrRMr3EJZknUBywwITFYQ/guM7eOlbwDootprkFS1PFJvDJ
f0ygFJYEHiUOfJ0K1DYZpXfQu9NSt3/wqsVrzkgkSxw3R4/ecS2R/nL/zKPoVm2U
5X3qoDZwnV0Ne+yK6F7QcU6G+dRulHhmcy+pNlJcHgKxyoNebmJeLj1H5bX7sVHg
LA5IgcX9mIgB4HLgyhiYrzPkHS7zRU3cBAR1XkHJoPg2JVeBCCRrHVLTmK/5IerI
/EYd5bJ1r1vEUoSj3jspRhbJU7qik7nHO/HOuRup8dJoTR8soQC2XEMspA1E/nXM
qJgy+F/nMglC4pd3/QgS5jZhJg+t3xq/0JR0EKgXIEpG0VrJxV+Ed+ZX4mynkDPq
rTpclnzkBHFrp7XgzAxparR7Oa7FZw20Q73mzuxo3bVRcLySw4d9Ll8oXFtdqQEK
4qhH2cKn7t4r+vxzjO3EEdnsJPtt4/kovDNCjmfcCMoqYCt7C+bqf8s4XLxBzQjq
KUPYNH26xWoEaLjObRpOVCGmr6f920MFV4IWc1VAPJs=
`pragma protect end_protected
