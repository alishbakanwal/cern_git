// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 14:01:22 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
VMxASLiUECaTKEW6xGdfjAFyxKxBnLPLZrOy6NOJKzGNVBNKkOQvMlNlywufF3fT
sToLeGLpBXFFugtpbgsyJ1yOHj1OaPTh6GjkwLTN+IWe0j1i94HsyNNDObo3F7tV
PiIzKvIF1KYGvW2UrnySIty4MszDaNmGCDnMz93bVxQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3600)
kCVqa1t3dmdC/EVX0D4CPcIYopPqmMM5hpQNqvcZoleiXTkTKC7tOktU5t8cf7v0
J03yCA3R482qpulnJTPPWQ77vkjJckmqdBtL2n9ZGmWzqSriDj9rVzQNj2ONhzzK
RuXRRjZroqj00hKSQvcspkNMAbmI2wyk223X3nh1ATkEw86YjlqNF25In1VBF9cS
530NbrXI6v1duTESy5+Uzuo1dzfLIFBubXGTnQccG169wHuqmLFSrRbXFkzTWmNa
wnF7O3hNvf44keZ5/2B7tlt8tt18+0fmyzyTW1RG5KOV/qZ1IfkjprxipFAUFuX/
Lqv3Us9Ud6bejBhWWoUDxaRdvsJIxmELDZmyiZdHBxLauWgh/hufSSn6YFHQuqxi
TW5cFt7GmPozqt6PS9DXHJ0JeX82/lNWrZyrQAUarTAq3jkJvi01Y9QZis2usw2G
ZpW3XCzqhq1X6dhiqmazXq5FNEvaGw86khGP1aczOpRF7YncOfGmlskz5lphWhyj
3qet5UNHgBYhUt/eUWjw8/jf2SGfePw5tGa+dUMOAspuV+83glLsuzeQ+kuSZW+Z
vCirj/wnhFjrnx3N9xkLlgQKdNL/6tcc6MClXiP0vr5tPfuz9mtj+zPbdvu1griq
Y5rX7p/ssB5fHrOBXhLODoqcBkGXgr0/XdNOCGAl6HqworEkNdzJK/RFA4AHoOJC
//9NapuAX/sdatMx34PFBsxHswmRtn2HpvzJ3oJIhHqGMTRXIsId1DhuD1RDxPOB
7Hzf9xWsw2+kncqBlxCbsuPIJjHYZAuJfXGo98RAgMb5n3PMNG3j/DxZTTYML8He
ammmfRv7WU8qODfeFzWm8NekSSDJQ3F1Y56Q3O8hMr8ir7KTuEZZ901LcC7Sf10A
0bQuqNCRDRzDdxZMvEP3mJduhuMdHhiSmzHdYP9RwLLga8MGnHfoeryIB/MS3ahN
vNYK3mw44wrjmX/KWRqHW4TkDIcqS7ENzIFNPdQTlJt5m9jcgrZEcRUfTDDfHfb2
GmUHAKgZMQfpWzdfbYu7jzKQan/WohXtOZmGIfFPtlxVdcn9+AXuhnK3qsHmiIAv
MfnTHQUywIu7KzKZekLtYpYRb2QfnWes2Vd5JD1t2mwuqYaeGdlvsI0YDZ1rilBk
ByeefKpl6exOsM33iwlOiQHL74irrOJ7yNtDifgeYpX/f+f/wPk7iiwUARs3SE7y
0blxB2SNNOjftChTSy5my9QybvxHIHckYeIbQLTs1jdFpuvvWWkFxZk58qOkRGKz
Hg6p7X8BQy5VQhz6Ihgc00arj66HbSKlNrqCugaxqRBsLEB1NE+SNmeJBgTHyf/y
xpthLwrZ6m7VfnVuLar7CjqwDpjPGK/80mvbtlXyqm1uWZZBKs6vaPNqNtw4jA9o
oKQrLsjfgEHFWhTsq+Btc6XgpAU2AQIU1LWqEcGDc5by5aza5IlD9+aZat8AyFQT
yerZ+4U7XkBVWv0AiIXG8Pchp2+vJi3sXSmB8VSw8x/5d7XR1Ef8G4nNWNOu0WGj
PHiTe3rHYNLUMilSoe/WynBRXCuaT5Gsq4SCA3qb+/hWE5LnXPqWthbDH0ovma/S
r5/fvC/6NGO9ISYwEfjI2lYWtBQXCJWJ4NRYlubmfXzJ8UZKy6PCJVLBfSs2MX8t
1bnnUMd8uKv9tLGfHQGflCvgHe9p6IQNUG7Bm02Pfh3ANhzW9jflLW7TAGEd0iUF
1cCNxR8u0sGf1QEpbmdq+TjjSCFpb+SS8Oo+ovTpGxcv1OhYJLQ/xSWcSDkmPm9K
D2yYXYpaVwT2gRnl/AhfhJJksJCVUSe2/ISuXlwY5turZewZ5A93s3hpBaKy7ZWR
zGsq2JLg51VMKI1aY6LRib0ile1MFVBiII8QP5DCuuJzMnk+OlbpCyd0jY15kTUJ
lJ27k6abBseJQg4ZksBl+5SuR8q2CpntqYtdaasVhFodaTBRRx9PcLOskQEX32Ke
a7neeXF1BZhX6ig5wcxQ3Uq48b6PzXuBrxevnOOgEBESJPumThyFyuC2iBjwP/LQ
ObJzbzJHmTPHaPXWy4LJRQ0E9B3n2bPG553X9/BnqN+P9C+lkjJXQca9R3DKv7sY
GZ05yxHKaDvNnLDnsXzVk8ic+7eKDilKnvDF65SBtYY8woL53H3s5HFjwDUepe4W
LDI4mJJmrZnlh46jaANhwsEMuaQ3QkAGY9NhMT16hiWZ/SZ8uHFzidelKf64ZiYU
QZC0fn5XKCZ5pTPuO1l6A4vG2o7ica4vREKtuvx5o3S6+C5LQM3Nfn3GEp8WGKPT
S8D7j23KtqpALqhOHELoJ4ekWwGbvZ2vSQY/ULsQwo+Mu+WQjtBQ+wHMeGT2j7JA
nSlAmrKAQWzNYb6ZZAqyaxe8uhuK0QzE73w0anelEPeyJxZfkDcUgEnVYNDBNBdU
xyvmoT/G7z4DNEsKF2Uokp/A3trflLgbC1ny93C4fTFlmeSUzwnHW2Xuao0wNCgz
DVsBygZNiilengTqBtNDwvtv/j1thqaQllV8g45EOwTipn9q0f6a8qdPb3POnzKx
aPZo1eiNENWX5RrH4hxe69KiqRmUOk2db4XJK/vQwRhedTwn14YH3qGRy37upRvl
F6DzZBWjzfwnZNHMJmxr0rYa+DygHsiTO+o5t0fVBzDT943DqoJYTfVHX5bCq/W4
a3Z76H1wjt0xEOVR/1ApbZVCNXOmsuhpOp6HQjyTVaAQLBx4AMYXOjIOUWUBUYZF
XZjCx41DLP4tRS7zNpWDHzADeKcWnWYnswwtNxyYiqDT35twbkBWduCjz5bCwUaq
nEsMcHhDz0Hfnqw9zND2XoEaMup4mtFMs+Zs/RQdxg/LOkpaKHg9brszDtb7mnrb
VLzu2oZBH6C8bMsTRBqSe3sgbhZV+2u2X58UinjM9PK94jomI+mrX4mJlD6e2REJ
XWfhBL/ilP51TuYrukY8VxLArduoNZTOVxVsP5P1NKS4a0SwyLVSMUxIQgwJUV7U
tc3inHiCY2Ug8vqavonKKF3BXCnd2ndVkI8+QIoOvnrBp8ZfszFZps9azhQdg43Z
5tzkxkNNeA+A9QcUfVxwibhRp43GTyn7ip5iMvSz+7enALEWirtzFwdIB4wZYtjX
xHGnIUkYHiL7QaIqk8/8HEz3BEgFRgT49ZIykX1QZ9iLAZZrvDQeeEuqDNc2kg97
chdTF9qvLAQghvZyTDffKDtyl5vARZ7+cCEVf5GogJ4LWC7dHHIddJIozdXNVd2H
tz0hRN3iQ+mXRTDgTXo0K8AefvWDAUKM8ly/LGnccobJWRp1JLsnAwWeusDNdyxW
xhGmF+ufSuJPkxq2TZiCfo71w3wvxqCEA8dBzKnmR3AgvbTp0xU9kN5sTsbOSGj0
S3JVYIqjU2FGWkYfajtUkW0OSBZ9OQ+5rWFSFMUDvouKOqHP8vZ+pvNBqBUrneJv
4UaZoqIG0OE+lGmk18SC2jPNEOUP/XaG7B+P3SWHXEdzSfOIHBuLdUqNrZ4UF8tI
CUmVII89YCkGB9tHwwecFjwZpmoTggNeO4BkUSTC+VhRG2OM4Nf2Q5AIJAojGzv0
i0ukbaSLpxYW5noVY0eya1O7k8icDDtyi4eB4KneZZ1wd/JmSaQL5d9J/0lgbbb+
3EJOEPZlAg8yo3ae2tWch91E7HA0pw4BUHWrpGintC/RrUxRe+71EACeEYJTzrNo
zzBzcsf8YaW+/ph3j6xoucN3lLyBayYTBptB89sVY03wRVTrjUb+xCguU1Gs5qAh
pHfK9jx21BhXjvGNYro6WeoKEyC4YePz71AoHNa3aWxG2KMwfjnWZbEtBjEn1xIG
yM1Hf6Hko4SAzypzK7IizpZrZnNgpcgOF53bzwmz5EHG3UTrWtXBGdCHunGYReBh
7n5H5eF8R5eIKdSjDdwmTCxENWU5zC5C3df0c7cjzNJJaPg0lti9l3cwiOXhWyKK
9rcefbarV1K5S0Rwr7wCrAlrRgR+uxbeYBnRWwdf50ow0af8oynrJXjeoJ/dIo+O
tOp4CyIM5pMmBw89LhSObs4MPcu0CxfuSnvULADlKrSMVwz+Yto6r9xwVhP3sQal
TanZjALIgvHcxhc+jGyscEhEiIO/hYKCgq2d5pJaGzL6tQv6J899GDGiyHDyfet0
nhIRcNyCXVJb1eDeOoC85nJOS2Syn2ErWFzgqM5oDVCYaTTEidPKJiH0FHk+mG0V
kureRCCCIP1XvvXj/ilJPQgLV2uKZ7v5AsjtYw1VxpTLBYnRxMyU/Y5n4qScg6vq
zwQtgX2WomIlW7SfFhEP58YPyqd8gqj5Ke+9aSQZr0f2+Vxp18R7OtJ3Qqo3e2mN
oBKjihLfmKQv8DzZvfF7y4xTSAi3NYzbrmQFnJNxq3gYRfpMePG7oGLha0HttjU/
nLltsUMHEr2qkkm3GfEmOsVvtCEWOTwo+VfI+eFFvrXBPUdkdz5YUBHfbNBFyY2N
mID5VZBLtHBXYsSrp1vjC1gru/Lx3CnIZxNBIq4h7yISev4OZeK2eZ4Qyp4cuNTq
Cyfm50uCZF1cfBQvNGuTnq7RPAaHuG7a2mMgZhsHW9wQi0ElpOMARaosbPai6Pmm
njk8gAOQh64m1SK9w+3V8NcB63OfNnAfkeLvFQKV4EfPhFkolFb2ka8jk6DhhsPV
/ctd+x5yn1MpZwW5GYQxvk154ssydXdFsv6V+/lRe16g8kfk4hn5rIXkJLGdkucz
Ev6CIEHOx+Y2bSAj6gKl05NYRmZVz0mgdPTmB8684uAlTxLIs8NHV5u0b6u28pVx
`pragma protect end_protected
