// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:02:15 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
p7gh9dHRhy7U9vjgycaHO41kwnwmkCy0sl/urz7/zaVZIsv3E9eUZNcaL9VQ6p+N
VuKEzP0HO+S5vObJrDdYhGSyYgdWBGsm9ApV+Dfas5ngNMU7zcnroG3P0I2lIht7
v9Fle9Dd4dB21n2ZH3Nx38tKhKDdEkwnLh5U19dBxMo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 27776)
Hz3p6g67NavfRdH8EDww66KGZ+tSFWhQuU69fW1PDEzbdoSA5uQi5ytxzl+kE4rl
WmeSOULzEnCz+tBaXCXG65IARD+HubpMw4nZuFywKHyk8Pjza5Nt5tRF9Os0MFrF
v8EI3sq8KphJ1J8UpUDuzwjyNWo8FXgg7+1rPqYtDYtiBrCH1iaoRW3uz7GmvH0K
MUx7JH2PyxPZvPrlIlQf80GT3VOHAPgzPHoTU+94pIy4WucfmAaYxC3aU3e8WZER
micZLZWxxmodExxnwSgbWyW4xJmYR12FHdLKiLPlNjHFCpwME/oONEcyLxtkbhZW
JrRkn7sfD37eAAmxQmGJxzMSs/f3viWDN8PgqZ5K1+1R4rDf/ldOxPaxNf3iD1w5
JihTV4M/25zOgoEqcEik/do5ktFZEzduLZm7/FcxJ7AQ6Q6X9njrC4GpkssfgzR7
Z+cKEG2pUKdP6kJeyqWVxSGQvbuaKtlXz7PKbiw47J5mKp8rkppXPpBrwuVMZdDQ
W1RVsefaqDk+duBUFEd2nEUav3UVtpBqGjoSHW0BtR2Y7abGDRiDHFcoiDYbrzfY
D58K6VOksuxE4jQ+JkryyaNyCA55E4LzC7pyHq3yhvMTXRQQbed7SaUdF8ySVXZw
2igylTOMriRrtJ7YDamHtC5VQaUT/l8hKMpRdJ3pL1EU7UcjBG/emWY8oOtgfWkj
EBV3jGGya//eQt4phHaWw2QK0NAm/KnnpLCPzhZ9HAx1u2s0SpUQ8BLozmGmDRVn
z6Kxa6Sp8iVsfeGfYji5wb0Ro8E5DEYILolofM6XE/sakmDq/hbZUZdIgWAeaKSd
Ux0MRYKV9vxqN/QsVkmgW923DAy0orgO88T8SwXbz66PRU7slUzo1ZyhYHWLmxpB
pNfufGPmJX0VjpDC/LjPf1gnBaTAmH/LBmSCqaSpTKajmOqkmypxJui/n/8mvPzZ
188Bb6Fir5gad5lMYXe9QmOUk/xSMZ16ZsPzxbgFIDIoYuFwi1x6EF5Pnv7vx6t2
PRkYPTp7xzKzankFyMblkN17DKzgMrf+VRHEfIxsnGI0Z8xiz/zxJ70TLm49p4+E
xTQtGqG5n+GmJGwvxzKcWkGW8ECrJ5x7rpsKd5QmmgRf4YbHYcnHneiGpJPEh5OC
umCQDfOLFkc8CqPd+39gfEkUJ2ZzjNSdMVhERg/AApYh0ElGzdZsvRS8RRmJz5CL
HfmcQIRA4W3WFtdhAmXjpRnYHLVhS5IJNTlBeQIyOz5zwEaplb2bA0GHZJf4sxB6
OM+5zsYYjC6JdsJqSXBS0l6W5snm+GBzcdybE7Bop1xDV8FGur6k8Z/7UxKi5/fo
D52vVNN9/FPsd42VZ2tCbFKgbvm/9qEtPSz5cfTU55sFxSIEhq/pjVZU0bR9uofh
Y1kSfSWkjb5KsNsGSBzn+KYeZe4XC0ODXO62RDAAbHwwz0ug6O5O6nE51lKE4IY4
NhIFQaQU+CQfg1fzRPp3g7K/zZmr06jKT2mpYGMRFUGQWG7MZgNRWZyRFpOmTggc
ZnVaEQesZoDt/Cx3VTVo0ZWSrM/Cy3RQCXl2wflPvgAy/AVA0vmRSt8WDzE3fkJ+
OSzaLvSp9u5l5hDHDGXa71I6d1+/cDFsQERTjd51tJrRvZpNltAFGo60yYeRUJne
WKyLkHKVmPfz+GsK+W0CECjMoOF2iZtHTPNm22HDlaQ+cxGOKOyfz8dyywrJl5xE
XRXClpAgN0fNPuop5Ix7PTNVpLCUkO7wWnG/XBfTT+2jJeplShNoo+ehd9px/WHz
DvaysYlh8Sh+AVEpcqP32dluDeCmBZApIAhMtpir6/8PdbFfl6L3MlRBiiWmIoa5
xoHKtod2FZLDuv8t/P3tlzwE8BdGUJszji7CU2My2U5I1hUiYVMyGKhSs6+dQ1zi
YvPyCUXVMlM9HkWnBPM3C2tbIE/N7cLcdsr+8abet1Mxg5MGHp4ijqGaHEdEHNb2
IcSFF8jb5BPwBnrBGw53AXC5sOqGfaUUmMKdNK1QPWR2bnh9IwqZr3c85mwxURqS
DowjJJ60Xj1uB3AINgQIGsCPrsgDTzOqpvGdeJM7wIjt4PKOk/xmNxLU92oRWdij
ITwWLw8tn/uLJILEhKxAPhDFKD6qvSTdAjdYyziV0UQi261zZYV9l4YQGAglGUOw
OS507pDOEPwHi+ku4YgxuRawF5yCXvsgofp3/EH1IUgLIGLCah+Tl/skeCeB03z6
+QemdF6lQytwk7pNgJQS3OGUoNTyTZCZQeCsCz3/zkjr6S7Dr1CuzSMWWPuAmLFg
YJQzg977hadNLBNkb+LmX8T889QigbmA3x8GMPuPffhM7g+RjQT/yXx8Qrm3pslX
FjLqxsJDp+5CRVx8Q9b2Gol3thkp8D4+GJrnCOlS7fjfF98BPclPpNRcZCJi0NCD
08Ccg/1KxOpR2xMEGG2JDs50D6Sh8jWTxeTQAWFXDwiCHAAs+JOuMrUMII8OI4fc
ISezhVQVh4ASDrNvWSmN5M+gJNWZljDbldXTDPIwqE0Pt2b+EdcQeqUP2Uu7ticu
wyWN3AHm/r18O0b8nw1a28J+wDLs2e8bvkt6EEYvfGzlTn5bvr0+zv5mu7vbKfx2
6BwQadf68btq+Jv6tPna5mTiIkH0YMNl/QLe0m6RB2spN2sahhEq5QIeUsW+4TJD
XV+uN7GRcMZaoMC8gU6sRBelIDq4l3aNuswHdOwTYOd66G9BK/TIOJCmg7DwxUAO
3uTpqRd8qHK6xX4EjrKfpf4JVpXbqPy1EA9Gj2H4eLOy6mSB9oxCj2u2vJ6WpMyo
K1k3NDenFlmM3fOhcoKc6ouyhvZcFN+8E3bWgvizzlkofnRwUfFLsXwe3ZkQ4qsE
uiCjVpNtXjLVjjE7ZDnhH3E4gtP4rtfqKiWyjhvCZziyomDdz548w1QP/RxXZE3+
wHYe4mHIfjmvcNd+2bUeTmJW9B1Svatb0AEcCkzoV0HIy2j4Jid04vr/bk6C2Ke0
qZrrcHPiJVWb3P0wmaHE9wTxJc1qScyJvZGAGwNkD5kHUBqj7odbgdXckwIU6/bi
9td6mf2bCjYKJq3aUdjYNK/NXT3JU20E6za85S66KvfEDyYTj4kqm3EUQLG6TA0G
l3vQTfvaN4XwTqgbT6898kcCGF7pv7t2N7r1IgEjD3h5Cr8w7H73aZkDxj+j73UO
7eQts/oULASjaiRupqT4fwelrXPjtx2b6l8EmizYWA0RBIKlOm4jHsCblBlK//r8
m5cumbe2X1OXJHKvHO9YZMpmmpdP0hZWJt+yDmliUbq3jCEm0ZJs6QoNsxHKMR5d
4+LOh9QQCIL76mXlZxiJnTkRqY7p18O7XlTv7PS2NsCr+Scnn1xE/meMqTKq2tS5
utjV4gLT86jzE6vXIWkwFp90v0eDePjCk00SHYj39j8rYH7n+2QemtYkSeaD/8cY
OiRKsOm7SU8xmYdGsC7qZ/IU7yJC9Z33uLXSIJgGW21BRU8oaAiGixJs6X6whXYs
0py5lYcfL1E6fYOrnqd74pYUuxAkT7LGjL1fzHXRyETlfjwAEwpG//F9yBlT8gpv
lDT12pcX0Rvhu8ZK9wndkw4yO5cqMHjBALvc/FDG/Qjhu5Tu5A1KBgx2XC/eHpos
hct0UoR+KD3kAq5kSVd+MqaVR6lJRuF3Sb+Z2dsNVS4T4G5RGme8cxk24bTFKCHb
iCXUoPPY+iP4ZyS1hOtlrjtIEavzS1QTQh2uKS+AXqjiLtfc3PBrHLAZHRtPzD4w
3lOqawbxQQptEp1cEBwXLp7ldnyPJDOJ67JLqTFrMXwwC0kLvdGbhBElH8RNWr6H
pcAUl9rBKDD2HhZTTCcZmG5RSaj+gLBnfrMvpmv3pp72K2ebbeFCh8EswaQsOQ/q
MSiMHKkjO6k0ICc8SRYIAx3Kf5UPs/YPKfsFVpH/xRffzbXQT24SgJqzW+M1EoJ8
YiOcQnb5ogyNosq82TFvv9Oa9qTK+CyzmC3A8e6yd1KrYt0DbupytxPbF4YZHPt7
31bIfamGfPsjHVY3Wj58IKmcyHPSqFI3E4smp6wzogjhl3ESxwMx2W2QfnipT+iu
VTHSnb3yafcndMwrwfsjRUTYC9L2T6MP2+EOsKbQ1cSI3ukaYddCgNxBhMVALwZj
qtOtKsT2/qBf67TVfkq3bBZieoG4wG34Glh+898lQQFesGARKBpGdILr8M9Xl8RA
uSjG3F+y45KX0mip9PRZpiULTuFNw9S5aRbErYQZgOCC00vHnUsfN8Qxq2bg9RCL
3da/ixDZ1w9rYeeExeG26GPc9+IAMEglWxiOEhqi9b3id1RSF7bwahu8xm0Fn4gR
+bkZ7yV6JeiSwGGZe/OiQGlamATUVzoeaEjw9lmIEZnrFzmX7X03xqWvf2u7y2wN
feUBL4d+BSv1YrNYf4D3fjfvNAut9jidIWiUxhkxsLlXFXSmo+95g6oTCBNDGP3Q
01Kre6m43itgWlrY2fG7W0G0WPoTAZIW+UBKp33fnGlTt4FS6qxwE/nRrDVuDsZf
isJfgppI46HR1vlcegbu9VgLF3E+CRsPEkpu++ynUjYhR6EqCUSKYWtWDap7uecZ
Ef5EXmDewKruI+VyuevU7MYlvG/De3XZLK4sZ51SHhGCAX2IdwHROzHh/aTaQtq+
PIA6OoTd9MEwHtS7F1M6aL8LTFQzud2TIJ6i4rN4XSXNd0Lygc17DN4sI3C7HqJr
FA7quj6KTYShz8UjNKdyZkZ28S1PDHDI9cDTSGoDuV1TrkSBGtEy/H//rPaE4Md7
eByq6fkSYUT1h4jkcoyoypaTaPGQ+/ec0S5bLOIgZkfKy9YG0RFeMfzwnI42epHl
xnEzDs/7T6Rs/xEhLPhpI1MLoxe/RN4ykirXlgomHkWK4wtyw27SVQRwYLVxi+N6
s3+xEDzuaLfXQpHbzaxCyE953xLD0h3fRww6ciZFYzH5X6U+FhUZlNRrYJVf1BKn
ZvuGvgNnyYK7eWiUzxyC3p2KoMdPJgn9fIYmH3wg0l8bPEQ+N3i58fllGXB2M/vz
4jQ3i39f8BH08OGGu6t0tFeFIjUpvy+R9IPVO4uzgTAavf5/HGwbFZZ00zist6Fg
eytaYCQJSbuqzjzklbKhIWN+hYFe1OnxNy+axVX/MrryJy9AS7CXEaTUEV57Pnrq
ei3c3mu1bPLAevPsMxSgC74TyqDaQivWjAHE9RbnPqi35gFCm0qJnNgL6127xeyL
8VO6qs9urDmjUcDupeOMWDB75Yzl6RfSlbOT9OY0bc07QVll4D9JLLs5lcHfdKoY
kfpmyAxlVFAwSeXeHPyk3nWQnvV73/V8K3VjJkZCnOStyJKdNH6wK1JU94jjj9g1
c/jvIiM2apehyIea8s4NeTQfWK6ITwShyUjwaB9dq7HIIjPM1lduX4e0QJzMA+WF
gRjCQ1PsBhl0e3cm6TGOzrmGlhh4srxzkeZE8CdlsV28xuwgYXepLa1dfzsT8Wgp
+Z06zwnW7Ul3oxQd2lGjEuHSXOT+wWxkosVQeL1pn0odbUnFhDac0Gg+JcN4pD5v
FbLWDF8+DsLTIHiT12p1X9X18PgFLjKTPmw3YRdRlAJSynZBGNsGEMaP5eu8gGsL
oQ9oQIEbdEmgCsjf7f1peJI5VgCWjcLYz6Hqi089+WZpIPw1At1tGKgTIso2TDqd
a7EKdGdjvAoXJZUBT24hQ6U9Q9eFMDh6aAsqNlOIXuaQ/Y/UO1aWZpL67jnB1kyU
RVaVVa2fOWrv/2rSgMf7SutPiiWV9KO5sbVCHpp8kQLlRwwvXETJ5N+tm1uSSVq+
+faolmlfmbTxXCjOvNxDtQ+W7ZwvzobMC9ioeaJARf45lToRSYb89RmfMM5Ooe4u
kLbaK22Wtgz2QPGAod+sMRZQmOyyLOJgmrb8hF051ZMiQfLaxgtnpMEnGDFIZzjK
JPvqpjxquAzUDqoQG+PAhmL0d1exlFeQcm8m36AyZXpiCALrQB8x7ThF+gL0uurt
EqsonUB07sdaHq/JKfj5aQA3qrWb+X9KWkJ5h2rYUjqqzJhyuW/Uc7QEu7dLrWLN
QJDnADQoAsa1P9+MQq65aaJkwa4TOGTEx8jLZNpn6h3K2UJuFOo+n4lrv2vjSsvg
CGv+uUCket1GpRRu4PMHCWIWVo2UsMqv5wdVfsnUUd6zo5s92tgNEBvbZylk2LsR
PXNlDLW5nsHbJkAbiFMNe/GDtBD1mHkIpoUEodasF8qBoHu9N7gD3vFyuNHrrN1n
esuJfXialbNaHde5ORQ1t93wsUn5cnz9VKsgnD+k4bKz7XV4mohXiAzLHcwneaZM
kCvtM4rpZUGrJpMt4Q23bIEQW3tnE3CB6d+8jpBzfDYd5mGPED20kqPZ1fa3zHjV
SbJt7LNxaZ3m8I9awbYjsXHrQ0w7hJLIY/sTQ4mY28WYTAValXTOSlwDZxb9NEBQ
dGG2xAscHVOsxWJ7LvU8hK2xVGJEP/0vqcwXvz5dJT+N3ZdKoAHmBYi9Dj8Kmdul
Bg+9dLVcdl4TQy2xjja78bC2tLiY5zETfeoA5C78uDolFVIJ7mBiRVw7ndzi+XQq
nKWQOxB/likyl9X/bSUjhinDU859e/qrIQf4pn5yI1lF5BavDXs49QNmGp9zhhFs
kGqbIGNguCbUiEKL9ioSVhRKKbSjVjOntfH7pUpLhhYULgExtf4IJehIE8VtET2X
Gc6/Lv0ZeE19XNabGZD1CXCGe4YYh21FyRk6/sa6fiZx0Die3Ny+xdVTDkIJt5Pd
NSIkNpZnz1AiWOG8VV/IYh2zDbJVtwjiabGbRWO3DAHOjO0kAkJoRIALJXFiN4cX
6d72ORYfoIt4j8kOEjqWm3PEwfR7mdlAu/w+loX/09l05UmYsMcMQdM9FViKW9ji
5kRTsOVmDpUw9LY0Fz7gnwVRgff8Aep1MNCWIY+SoYRfM1QDvS5u08pm1lZSNj2L
rZcN+d19XhTBoy9D0+tqXGg/QJEzzN6PM9IJ9+cJcqJ+TNjW8Z+H74Cbs/R7TkBz
0UIaDsC6Iws1zWZGvrrm59cUJ/rjTZKqiaNn+Mezv9W5PHwb4MdUyzYgYuz4/DPT
VuRN8e0HYJhD1+Ou3pEslgZT/UDbj8qCkyHkw8A4EWHSo6pYhqxhGlrOF4Fmunoa
3Mv4kjmjJ4FQLFWFRwXz0OiL3GnT+VrzPXydZfmGOAwmpsIEKROgoidSoAIOFs5D
dypKD9RX1Sy0Ao3KIfHCHl/KWWdnJTyXomL1iEe5gCXqqtyQL+42oinU6WtKrvrT
Mdjqs5B/BwVJE8kSGYBTfqEW1WZNP+SU5qeWw5ODTdvVk27DByQqcKdsowkH6tz1
T5pckXN56mpoT4OFJecjSPi2c12us894PRtQMReesDDB+I7yMnrRTEVcI367JhS0
37ze/RO2i5IiXM9B/YoWFL6XvQ5odJxPGoERTqFa/HXCfiHSiA0raGZw4GRbPgT5
A5Znk5musH0Vd/z8Tz+Qehbelw3H5S8rDiINXdxptYAEeld/HkU7WbKZ+7ou6zQK
2vtZMr3aNU64QjH4o2/6JErTJNzvnwF2fTOQqPXk81SEfd/dOEGtDQwfRDV4BkTg
iRYE/xSuxTYjvyCroaWGWBjhN0/4UicjVJXOno2VK3q7dx6v+U/Er2O/EVwOTt4W
T+kzDmE4t2wIgTJ3hdd7Wsn6e2OOPS4UxKUJnWkBFmPuplNHHv/I2wp8dQUmOVEG
Yt3WoWS2qn6FfhT5QvcWV/Ke34vx6Ukl8XJhgpevG30MIsnsUIxYLVxl73TQIiFc
bgX7UuiLaXRj6MpZOeufCTIElfDb53Rpm5UhNfaeffvXbmTVxSxe1TTcHzoBxbsy
7akMffbZNVA1+WO1zgD2RXSgpCvIOpuFaX66qNxfInnPo7j1vPP5/c5/XMIFFp0+
dPbmV4xoThWoWUAP8eoUzAPwBJYr6lBB/hpJHUODMnwndRfIYTPA34b2hRDtU58W
6F9cQJqDCiTVqNP+iZf1DZUOf8+nf+PRopjQkctxD8v3cQf7euMB51PvSdYHJKCt
s/YNFYS+OO2yYBEIy1+AtfS2aqqCCAdh4LrHRWymEWMRez5EY1mdqX5cJ5Gp/zkm
9t3iHTmWuLktprXIO8SkFqCZV8EV5oNTvwlDJFCVdqlT6p7JCHaTgkGY+jkYwTAy
kfpMxDdgq+hqVMKCBEtCeeMLf+ZEZzlZao1iCPVLQoxKnkGiARP+qaKIIX9SH9ZY
GtfkBZeUQxkQjJUG51r5fqCpZJ+LPVJVuUwNGDedR92q3fYY2zu71KeoqIkN2lgp
x64hfvdIlcLVj938yMDaK9/RdEn9/pcGhb0bDi8sxbZLbejNxVE4BUfBVFYgwIEU
itKL97G7h16G+4XEfwxJf5JBoTz4cZSlmHikuwHQyRytnOL6tYwXWJZ0X8UtSa6J
Nx93KN33mK/9je8ERt5l/IUSxwi4AaKY2yZP2PbPrF8+VzPaG+EupGGvEigPQ0WE
8ezx92yKaxgVSB3iy9dvBxQrDW36SOaHtK6/vCmiEanQlt1y4pVYXHlF+WFqhGQB
w5Kss02UGs0d9INz3KAyDZi5O6PO0+EcLk1iTqWVlMNtmoVaWUGV9B8FjVfF6Sl6
bu4Epi6AayvtQ1V+lGZS192AOQrLVEzfZOM1ESgbl24R7F804ztGG4AZlzy13q3n
Q1geNvzFdpEpYkqNAdNuWQCdMvUqCsC0Op1xJBj5T4EPpBY1tDfncjranLwdG5SY
JLictibUxBI/eUNapNqGJNNnA9CVol9qyVcr2V/0/90MybuITr1BgfmfCcXf9HVY
xeemiASA5UA8MbWnDmdQFnv7rHF7iw3+SUR4+CjOzkP1pKzD+KJoBowizHazLqc/
/QRZkBuZfHEI3UBcWm8S49/cq/qPa7+Vc+OkaIT98GD6oxQKBYjzqsxj462WAY03
0XlxiLHbBBv7vcMbHfWGrBdFzAKuRXtMIwjj0mmB4FRwdYH2Md7rtdNIWBH/P5+w
4vm5WZi2VdIdAVFy/5sf1X5jw1QUUjTVfhTWhotD4X30inw1LIUpUNGIPBEqCPDk
T945N0VGAsRGUQ90PYV+yluf9R5bqL/8QI1w70fiTTvgKo1L9WG8OCn/GSAOmOTi
e5wQU6HhTDZNSs/JPl0iN3SHZDE9ETVdwwjkSlJ502s8ttGSLbHm45l76Kpem40N
UADM4to93/BYNb5l6ANaTALiWYO+WLapSKTtLrjh/uqxUxp7Qij3PCepN8JQN3zN
+ZIGzEQu7RNE4g4C/6x+rHKpzK/XM29RIgDHeB4WvofLZ0HR5Rez5z/2mCdmXTrk
PL/y5FTuHtDw3o78/zMlARO+9KGp3SSdGzl3GrZ2t2C8cjgY8TuSTgErEvZjVvBC
EEqW0OZudfyDypbAGuP8J0fnpLwZ1/qfZL915JgbfutmUwDdFB+Lm/n0GeuiJ2rc
1VMZAqX6To+4iN+RdD8EzLlqKFgzk2bWaPNFe06X160f/mqXKW9p9T4iZZzP5b5s
/jHZ72FS30NFfn3UfqguDAvKv5hD/8HDWrRVjt+k+Jry/n0Zv/CkSR7RSeEBfEUQ
Um5t/MtzO11OuVPw7YaDAaNeQY9IsB7aJB/NbefNe/Spwd7wBiOpouGjN0kvvMkZ
OFfIGCZm8DjpAq7QSmE0lQ9xkiN9KdDkyEo3xgLErgBpP42jW8XELUWljFAgIIql
RQVs3JLiESbIuAGwM+t/uraNtbD/KOZFsyaHQDIaULrgZcBOzsZBstE5pFZ2Gh5o
lAEOaEWMgtrssSt1EkMUYpOUV1ijnDi06WIjTfsokgMxKCqHykFaFKBMEj7ytxnS
jjGGOD1LPbtwkJvMCDch3Ixt9H2VnpHReSSjPYH9DIUAoHBAxiEmUZlTrPB/JVKz
yCVTn0wz0jgSrlyl7jzqqgFQ/9K5kEGktNzDLZcig9EvyO2HBFs57I+7tHMRxM4d
lRR7ciXAvE9mZtQr2eOVeGxaw/iZj2+QrJ9BYUc5Nk0MLuKDdEbZgq+WihQHoeLK
DCJkVYsuTJarq3neO3PAW4BC7BHIk8ALURjnDLIKN5b/Tw7obUpPChPkofIp8gM+
dPtELMVWPVoRDClH7uqU24V2MrsJ9iY3v+f4L+MfMqJliIItg3jHC7Az75bLBkud
Us9CnyN2lz/iZI6VFto/X+q0d16xNJNvivYZfAQoy9v68QpXvDHqUNE6X644ZS+1
6sA9N7qmXejXC6llTAMpXaTrw5m9u4P46lyDZKxDMLDGtLX0Ls1RblZZLMIHm91i
QK2/J6Fio5gwxGuozuey+2nkHfE8ilJokZhebdNhheBnrWdzmH5wBAfRdfChZ9+U
VgA61ROqnD+FdkoiC2riprv+gcDvDW4oK9ygCsBT1bFOmy9KFF+aqtclXP80UTMe
8kEKXCb7jBSYkNgW/V6Q26Gz8o/broEWqzN+jkt3KXbEH61/03nwWe6IKPAo0Ply
Vv3NANCuJErb7oiLdE0DifjJrr00GPMzF65UwXsC1Gn4CmW6WKMqqMWitFUGdvzu
I0IffPhM5HSOPI3ViIuOHTH0i566FPisrPKqlLImvBD/lJAWLhmc6RD/ZbE2f3ZA
OvANtNK6hXqlJqh8UPCa50j1x2PBdg6qObKWL6dkQexB6CAxCeR8KaljAk87ygbK
u3jWQHuLjEXTIxJ1lXPgz08R98mhIGaxgdKl9rTBHbrf/+Di1f9brCiBl8sE2dMp
y8cSvIj9cUf5JJyqea/33gYBK8NE0FV3N6yH4XeISGKdvvqekhZpRWMHUZQtWzoY
PLQ7lnPvSnn2qgLFMrgpNepDcrNveZ7mfINSSWbprUJSkEvYysnt+4Ism47nzw3O
yUTLAYA1SWMHIqsKgvqokYXFCB87HhyQpwz1wgxIleCmfnBItZQ+uwHkCv1Lxdto
eF3Q4aua+PTKdW3MvK8SnTfRMkO1EmLWYsZYgpQMmMEwMO/o6Iyi0ywuX6AY9HI2
+AEZeBtgf8VaJLa/nJozgw8ZFmPdOXpwEHJ/iNsog82ItBQraZ+JBoLfjO4YQZyc
bFfVeT2BoqqHNsJEA13j46lL8MqRkbzYAS2ytv1q954+EGlzHLG+AtuzZW3ZT48b
0mPgx5kzOcOXwfIGP9zp3cJmYb99+kZLK3+w6LxD7WJi/+C+WDszcV/r1oKLtR3u
IVxsfTPeekefefr0Ct9Tp7XlGdbt7wqt1Wc0eqKMiCextlc3O4/OVZsPmXavyJSt
qm5//joauxEySATVkHTzRLTQQwbJcIQVJ4Q3HNt8CSqsGEB3lIMxLb3109vG6ocQ
gMTpVTfhovtUYVYVvG3idQKo7GcaGx0xuC9Ew2+qJ6mjWaLhn4EypbaRrxjnN2TM
SCSpt+3ukNfhW/oCPDo29HtAoAPt4aNxlTClgoC8JTpyhk4jPY08MWRlFwsKlZ4/
SKzkwpTbpch46QFs0xQgPpsKMX7asWe0EoMzs5Nfl/YEo+VVVp76myC9B87hjwpi
PSL3XZwl4JRQ8htN2LX7xUvclm7rl42DK5iL2Cll38XJPi5s1mVkjJpYrDpKri/k
Zf2jaFyacmC0LH1ALA3Zhdi6br//KPYvIIhChXMlaf0vjShX+rn0xYWxl4LC7Ytq
rUJyIT5muXhWJWlKicWrOP9xqy+xURCNUmguolgPeOSkrXvqe5F2c8fKa+3fgFjM
+AfcehtfZ2EegzS5wYOgfI82Uzgq22kqlMhz2G8yxZR6GqjfhlKtM7rR3OZicZFm
Nm8mbaHrXIu+9x1AhdJiTb2udC+DpbEFHXzPgJd5oq/egL5D7A4y7C45ICQWR7As
iowDUA1Pl6hbvyUZZfN8xK1eSyJ7Ee2LZftGg7fuH8wJD/6dQ+pO7sQjFThcrDsS
ZjA3gxzEoSypVG9nkIO/uT8PaqX1B4M9zRuidSfM9IidJeLKiXJaSC0cRmYXB3pt
UJuPVAnA4nPGP7g8qgn6jh4nBvDDqnKwcu4J419x+aaXRS4sUywXbJbW7E3EPBIV
WEq0Ke+8UiMpD1G1yzNxG5tpyWPo25aR4LEiDhUxfxCHafRhmGQVcKD8Ifb7J5F0
W6b1bbJsyChoMA9JPAkQnACK9yscGHJuMgnCCp1N6Deb2vKoF7YF3v/Y3E7PUxdL
kEVxWj0RnwXxyKC68HtUIQ7F9J6yuhfy6gipYV48l2d9R7MdPSQtWRSoJCz+ZXDT
fZtREuG08GamMf8an8hlZuOZob2N0GUmU01BXMFbKxQuJOVt9jZRAgP+Ts99jdrg
BHBs4AEkXis98EvSPsRB4PcDYSj3IXft9ILMU10uo0qpiq312Jy+djHDYQ0a1/tf
XKcgDzLF8dBx/2d3vI9q7O257I9n1XnUyCo8x2D1/++NeiO4wNgbzekROySM2DsJ
7GTQndxL0beuriySNZopKNjwzI4z9lf9V9YyFOO0yubHYzxYCbnh+UyGf3Ubdmke
7c4/eCsdlOs0tHjm5SSXjx+If6Er8RjuWTK1fcirCsXP8uig+DxDtJz3t4cQjaJS
TKVnlR+3AnFAszYOl6JyYzlhztwpJoS1N+fWX4b1zzZ9rVgU51OY8jR3G2GOvyWZ
SyL4GEGthxpB2e79fMlhHEh9IMBrRT1b9AGyXEIg5pFhz6YmytsHhH2jYEjghoDy
dDnhz4uT3UOKCCu/PjoYI+9chtsBuX/+9AQcon5ou9u8q6A+g/kmrvE1WKINe8sZ
b2exwKQvDSFToj28soYWkOFj8B6HpuuMNoZ9yanA6TktCGGNDAvK3CuDDsb3Pfd1
4cUeSwH+sFryJXStFgVxvWIQZpRrTmJEcHmkFcX3Re1+zj2gB8PKo5+K4CJuexS0
rjyPhI4U22giNoQ0QzoebSbzvlLmAB8ORnutxe5BuygmvojBy9LWYi+4F4soSBpU
duBGY2eOL0UC6+Dieab+cJg7Z5OME37qzGl0jaohmNCDaPg3xgDbSH2gOSMe8NxL
76jfEQqtZsbCbGxzxUAF1gDM5X8FB9hDqTAo8m8tMbSEyC+mJZ6Y5S2LN7VFP4Y8
Efkib57ovoRdc0J6ovpKTbsM5rtr6cDbKTcd0Qh67WmWviM5DOIqDOWTHt/AiGAG
5xMMWfZiiNDV6WhN5knoaq6PQLMAzbxHKhXmMSZ+wyO6Cbwf0BWebr+X1gt86Psh
Rwq4TrY85oxXfgGv+G6exDozUI76QLKiCcLiT8aV6KmNwlrpey+DbXed+DGu4KUe
DbccSx5lTUPGFIOX252RhIf2bJPmLm7ZQwnxJh0+buwMumQ8KdbAOtpNQxuuT6hX
AcpqHb+WZ07riZZUBPmZ3Xxq+m5kU703N5o0u6hitAwpfo0LuZCz9G4/zC3Gp/C6
I3y4hHgvoN4ekuaXueaIRIteKsy1drvKbuwdXAkEwtzHWeFxPtlc0w/ZcdLRoW7O
vUUwM9422+2/VthNN3NqzLqJNyrECPPQV/ccbvG0PTNHlbVhYvQmKpGXF6Nn9Iof
v1odQiIRAvIC9WASBP8rjPRPNpBDQYDgQpKccj6fcosPRaGuzVt/WPfTora2uhP3
W02zLTd6SwYadwtQ7igFStULW7NMFu8oFhjj/JFfLLProMnriyNYbL0VaVRlFdlE
sVUYfdJQrzdOxaEtQXQb0RG2h82GGLXQXmVZT+argzhyAFOC9WQ99ceke8OVlXOX
TN2xArXgqAh5GbE4Jkf2utq1POj1cmZpdaMUE7PZH+SFJSlCVapJQ7OI5U/Xs1vy
QNahk8sEIRGKmeN0HdMP0UNPWNdvpYotPMTGp5H8hzLxbm8iKZqZOKQzfZQc9ZMb
7jdFS1dcjOUn7sPtj/Jwa/xZVuV/f+ZWDDYJdogIWCyXzQUbr78h6REL4geERR2v
Vg5yQfEs1vN742utfv0DbsSlo5KJHmF23Ix4uDNgmfp9Zk4W5nUFmi6GT+DUpMPR
nsUOb7XeBEvkCx28W3qutSfvV1KLO1g+kRtQQ9EzP0LCPReB1WuNCIKwxb28ExhK
xexb7mTCOP1LyFKp10v8pmrNSl9KMGd2QMD4WJPSr/pdq7drpEmWvrRErDAy5LoD
LQH7NegQQ7DfgJtuPeS/Zsbh72SdC+aHulCk1BOjySsQlkhxh68iv/yGGWBkKOYP
yGEodRDLwSxklRvFyi/RrtLDQ5NxoRYITmDb1Kt4f+rjFv5DIcUM0qUCH3is+bFW
AZH2kS869yM3BREiDw7CAyZA6z8WNSK2h4DWqFRYt+dpv2u4T9f7DQhwJKs9Og45
ozaG7drGYNQQIg+g5Nb9x1PWZGX5ecM9Q4Bk6xgnPBgIkIpwsSRiNRgDE/Xh0in3
Mwj58jViZYaCoq+NhX6OhdEOwd2yQePXkv7PFGIDjhL++s1gSHdQPio9zO+VOUuO
/7p1MzsGhfLNAF2QbBe6Pg42RGlxpwpgOH/P5/4TvAOQxgtKNeNvZDIWXzwIL3pP
izeZeRdEFwVu6l7ILF7Pbr1pe6zEhLkRKT6VJzKDoEtYR4ZyUSxbX89kbhgBj8AM
V1iXB/9HfdMpbr++ATQNXHnrCtewvPQH+xjZXNJ/rBoEDXfgpp3BFwKK4md4JQKH
XbKDs0UdN+0NAv/p9wZ1HfxfnCNVLUzmMn5VlHPW04hsUzsxJzz+PLl5wM0odIEu
53GpC9bZVGu6C/gJICfCHAwwyKtTPCDkbSNvpFaq7QA2O60ccYvRpqbQmAAdrVfm
y3r1SiL05pA4kt3Up0XbB+e+0agt608qNg82qzC5j/ALIn9NCq+lpo8h09UNRlvf
cdojUcMZyCStN9swS+sJhY0F3CU3ZgZ9EGsSgF1f0MtVeydzHLaDbpS14L8oBWDU
JYPE8dHs99xVbtzGkLmu1Q7ZRPG8md0rpjLLDqNU09uD7xJKkVCp+nI0kCYktK0d
PKVy1/ZzOx2HCDuOZEl/JNo5Nn5pFOqwXkQwxcpWIJAzolxK6i7HPTpkGtQdk5sK
4hJkF/fLeGprSwu8mxWnf3RDoPNdUzTxHLPGARMgEtqKaD4K5fcpc2jyNmqkp64I
F4buCEpJwbUVSAUOn2fbsSbdB/thVyGqoljR0np/aljP1DtN4jvWUw58+J45RIQZ
HrV2rGSytDkbmteo4K4jM+AYKq+48lao6iHoHAK6nk2hgAwh5IOWXa66FFahE8cZ
g1RzWrb6tCrGX5Hcu4bRSI4z8tVc90KfCKtQHz9VU8MDOxADpMM4jcoxgyW/9U6Y
3aOIPuQLbsfpSeacGvsegvI2tlyQFCvAIUg7g/ZDgZF2tUJRhd4hDnyA2LdFbQMK
yPv4wHNygCbyH1YWpQzCFdNU11cya0WjYjRlfyVGPi5rCNjEqMLeN5GC4tk89q3V
Hu/wQmlyRvq9AxKct6UQ4H9+UegQooKFIl+iCSoosYV71AEidUBWWGxzeFQav9Kz
zSUBhHoTjTQNyy7pZxfsOlPUTkm3pR6WTYJjjlF5UReNpoVgqs/NLQK/II8LHRgT
WgwUECjkTHDq9a5L9hSl7UH0R6alNsVVVUyZI/epqsQCpXQloUfiZ+B7PpxRykaD
KewuxtyoDvgQefHzPp1wbNmI/DufmjjwHC/9hjy5OQDAtvAgle3p3BR9PXu1Mnxo
U0qMvXrl1As5+Tstsx1gCpKyhF7h21IC0BLhpiYDpwOO63a+4raYcx8T9o6Me7JM
Ce3MtH25jSakiAXYVebeI3Nm8lqTeMqrlYyywyLQFDcRLBKTVAq8YlwtCjXdD/eO
nCRCKujS24EPgiuiiAq1wzkYvT9YjCS97HpSGoAAdBefZ2PIJAGR1wJKv5YzYurq
7iffZs3iDQiYDosJzt/2EUREXMyWhSBkn3mhITJGF6BV4+9EifnKmwSHLbcDG7lx
hXoIyEV6aorgRh+K3gQXfBVkBDAGpdOc6iL2PdC+286JboWVG0+8qVJnvBnhbcco
bRNhFg02UdFbe1oR/rDBQpF6anSfBC/Cm5y0RTCaT833LxYbRKnpCKS88XwznVSq
kFFv5C91tqb2JdUvElMUWkI7h0Ij3foyiQ3apimV4R5qVVylZ6slayVdG1Amiu8E
NQsS2dJNg6oGrvBpgqFFVJ1xylyRILrM2nDRUl4vgmJBC7zXFy8eEM/QbchZM0ok
tbT5oJM3hFpLnbW5n8fZ9hhghh9N7i7B5rN8lQ3XnYB/VIA1JPCiNLZy44sUfM/X
DiFmpr2G6+AlVZyIDIGbB4HaYrowHUarFma7ORyuAgZXRV+UIwPkG2KTPDW1Fr9u
paz81LxWEf8W5vtP0ox2PohsBJeWRkTjLIY/FFuwRCRqSySJ9X34ZpyjwRWNlbfy
jEMRlh2z7dXxxKUYJHv+buNbpO64BHV6SGLp5t32OUC7fSS/fvaGKXg7L9dtoxJ3
QaBRNyGs6caYHOBZ8nb3qxCcdkEnSI922NV0+fWncEtRnTCJHXgNy6vQBkCQHOs5
yXmc713SxvQ1YiRFy0hmFGdua44mCCrPSFLgrbZS52sc4pI61a3Li9lSs7m/ho1A
dxyhkXVyVKzH1WkUhA3dXONUNIPmPu/b5M8kdWkjfPVEGBrRqBKtapN6kutEaiMF
1/Ogt9s7WKG559CFjyr6VMnUd8Ez29XUIfHSv3v6ZtclqmmHi/yuMZrknRuIpvWs
6N2ML8Hw3BLTG0nf3Mj6AwkhEsF1O2M2jDcL3fXjAFIb19fVJDmEUyaG8DFokf/F
eY7VFrmZIoyIb+3aL3x7vJUXvu2Ylj7hDa7yeH6e0ig8fm/YFRw30dReDoOdCv+k
GQy7nFIKaEYFIRmq3KhgAn0TwN7bIAfTiQ6ZbLbQJeUuYErs1hKtemGflsW/U5n6
YLYqmEDo6maeYPRr7J34PQ/3Y5L9/+O9jztt/rzRQ5M+frRzSZ0V/xZo97DvAJLb
47An9LXJ3k0en0+sb3RkQRPCTITS4mgPcNBIU8uOFaFeMqG2CHPHfx/pztVLAEAz
M4VQk2B3txeoJZTk/85MLt2+1zjzXtawwsVv+wsFplxxPbM3rwPK7+uffDMGF2Ay
t+9CdqNWguMvHh5xIKsM4Z6tTpSlMsWQYTY5chnccHb/rR6z1kUZRsArj23g0saC
mDBA05Z4JwDfVKqbQIfQRwixTYnjYMPDkoAtntu8AHtmVLGCwCTWpATRdZQ7U8Qf
bOvyZvNBa/xH4ccpwnBHTn8oZdwbov5/gzx/xeZpKLSjuQaFp6G3VDD4DO6I4zA3
jj0rjlW8cxW14BQKzYefOTu/ixE4gD+Ix/HsGDDYMd3RRBzVhthM84u07DqDxHIr
KG3kHltnwq6Hi74+V7B2XDCYZuMJE65RaLJNJlv43RjieAbq2UzMJWOsMX4BUxqb
/KMHID+2NwAZ2rblLOye2XqReGp1bI+ZiqgG7Smaj1zs/Qa1GocGkmkswFWGMleS
hvEAu9S+Hxanxy5rdYdkqZPlp/3nMrw7wSqInST2XoetpqQAk0XrjPhyPSLdJZkD
66Xp8wQiLM/PGN7ImpepkPNoEJG4Z/WgNCKOGagCUBWN/MSe0cIppU0gtBy8IwDa
VUVHp5wjcZ7fbUhKhyg9NjRmjR6RoLAlkMDx5/vsXNkPnzz1g+ddnymIg03schox
o5XQrxU/Qj4RNNAQ4aHPbXKap96JwgZId7D4JZw0tF8uG2ft265zV+wlfCBIJLXl
Az7/H+lHPkVrL1Mn0l7UGKPxupYk+jHKL11Jq8mcE4azWILncZL3fevPMEqhvB2X
ujZyz4LZ1rdHsecvKxnR+CGRZ7Tg8ZP5H/QEoCqPB3lEpSXBlWFrFFdPCc0G9K5B
f9r0ly5wjt2IEZGSN82Fa9kqjvfS2PFOqQAek0EW8AnVHWHIL39GCFFLg8k9/AEF
WnhAJngJcaywiZSfbCO6itPXm2iyH0ALa0M2FLrdz1vnSIkA0f8CG6phl5xTTomm
DcUvh+bY7OMQNnN78tWkFrQnvRqrm+W53kMf1Gih5u1uyC3yiJisZ5XsdFIyDKtR
08R7f27HSbFkhhSAKTfzCv5rewrC6axyH4o+Msqq0Y69B6nwV4KcKD4aNOOvh1qR
5DpV7ei1Ryk1cA0DP/OMZ/r5t1EnA9xcH1gk4gnrZqshkSG0c+vV9/67b4rRstaj
P3avsn6K/EPpfhqfJQg1nQNAsDzT33PBnMJoYgvu1DF0GFdi9PO5UTJgqtCfjY8K
Qx9L2rUeDS5/8gWOw9G1+n/aQdT6kS3kXsiB8Hq3hOzHEy75L3HWUykTpiW7bKw/
VfwQ1YUz7Q0nTnKSF6e3fHt96nZl4wXlruz0xDGX+RD2UKdMjh2jL3hiC31C8STX
g7s76k4I3RHnbicIvGMyzFsLIzNzKSkTWnGXKCOYwvw0ybzEEJ2J0+P1VySNo1Xt
iaiDtk/Be+E3k6qf2jHXCgPnTVDDYTLXoyCIBPNgJDDmlt4FcFKtztxDLyqBGFKB
vBBudhvOHgqewzi+pbOP5HwyZqqMCdAhEFdTu1UlZXCZnG2/U4LuVtWWPj9541Uz
h1elq/B5vFhFWJ78FEFaxbXxhah/xc59Q7OkBkTTNfyWogHp17sFYK3dM4f45/ot
2R9fRDynhRR71wCabb8nDbv855ET0T4u6kll45ORgDUlwazKOuBM40vVIXijriYZ
VAQd+XdxHi62Ha1nIKub/WV5/T4J+ovJhQR/+eM41T6r+vQKTmoDedg5QzzrrnU2
M5S+GCZfLzDMMAL5aYqrCYrEbzw9LPL8oMex0UuM0Y67/k/MTV1hAHUW/gv6XS8k
82PGlPh4cwytnq55cHVYMOba0nYjoLK0QVLPhJBYpUGK9RxNa+Xxc0U1VG8Uwafs
iQ2dCQghTzqrHunVy2TRM2Ro0YSwZwQT44k0F+SLoWQMwrujBegAAjT4ZDc7GW90
tOMG7U8TJYBRzmjM2jcntGZ/0cVMYDc0nxm25BNEzIv7ujN2vAMujA5aa51uHkCG
kRADMAA36dO40aQl4vUxdyBkxTZbgUrcVb1ezlfMyK8nuXx5dso5PUM6biG1iB9w
rL6R49seQqLRiVwO0ehOiltw1d4kUJ9iwJEtQNud5R7J1No3Acryav3fIIHJP6Ml
B3XCVJT6HpXV2s4hdFYMp0IKOUYoQZRnAZecKrmW9f2W3TkObgdshBT1Excly/LW
7RM7OCOjUFDE+/EltbSJ00fjGRtN2wfc7WT5vq6I0IcNJV/+JP57Vz0+Fhzo2nAx
mN2KJn/VNuIBvnPaZZOJ5cgBcs/TtUeUO8yrSeQ1/PN9QcS35YefiR1H5QJqmF55
fC7ooJEw6dQuZLYPaeIR9LlGvoE9/EmJiDQ+nCzi7J4Q6pp+84kM2h3CH5R95+Da
JmMO2xxCgLbx6i/bogK9ydxr5cAayAzjNqyAfbmFXUq0vGjgH8ecCRw3f6JNFAtX
UwomTQERSDW4zldehj3wyj8antnM+8ByNIwQ8bvTFE3MA+EUoNT/8He40LOuirWo
OC6mOCl35l+2Ttvcn2LCdvFNai36C7mXQYT2j2EaGkjqEeGzO0Ev6EVHz8b4fj3f
oyd7ExbBcjgGZGx8tIdk+rmEqoKnGtEbv0+/wr0TkGIrkpIjwX7WoIDm7OsKqLgR
OymhtiindKVbG1po7zoyh/+fA+iTj0klfV6qoXpG5iV9Dq9wPbzjj8t7NoNDeLU6
Anr7bV8YUNf7tQ5YXHy77LZwV6JE9E3GhOWsRWlj10W9hWZZUO7J/5jVmdkQf84a
0i4elI4bxkjehF7fCbYLUasWyFAcv/WG96rnK3FrjkZUH4VAt9ngiRnrTgvwUDVB
wUrqOSiOfNc4Wnf3tcmaGFJ7DvsZJzLHpFaD7Were1zH5vjggeBwlIA+bZO88MqY
mrGPn7sGYXx7jg+aJHOkW+7GmqPpuP9gbjdFG8uRUfj4iFle+TUpn6jZFXG7AjSb
JJydlY3EZObhCTKeeLBkBpoaZyCRSk9W13Pr5X+AHAbFZA6O9+bBvtqivj4/tej+
Q9k+LW8H5iofNi5knN45RifOxMJWYnZJk3QlIiVt22UaQUa3GQvsOA7dcMZg/LIS
qQXtZsakP3BDaiA5xbE+Fv99qS4Rw1+UOzGtUuXLOki9RGgXh3vUhf+Rk7DKkxom
ut5gTNBVhd/djI6XcQLnLKYC4p0Z6BR7KFcaOYHaTr9VD44/LuT5FCQGzC44SBdl
MlK/CDR6yiAZfJAuJWEL3H1vHbtwuuo9pfdilgNJz0VfGmCYjtcglWGv1UwW2iP2
rJsCTFgsqBBJqsGpd+SV05mgZYtny4Lo7vj3kNEgPXwfSHd8M0mpge+W/dh9KQCf
MMl8nFPfln04TGuCGcFrYODv4hbmiTuDULyiVwmbhY5B2mwh1US0jZ3thLq+R+hO
EKBj3ROaN/SyHGV+UM98AZGqcbt8Edm0ez9NkRaEdk8lNgay0jfIaoq9J/zDuCAM
SgXbUMsi8uwmyTHiJUEoBy705Cj8sDKZcQDH1znPz6/lXJEl5oTbcEQ4r3MM58mR
DfKTbHiI2wqj3MO1O7bp9T5mHxqb79mSD9JqG36UdS7dpnXxue3icBt2hqyH2tB+
0m/BAmYm8fKohrnYMt59XRaQRKNVJvfBjxIxmrjoe8VNOZ7Rf/M6VYgC3uK8cUuQ
rcYRXJNmqx1qDj/shwoCGsstLe3V38P10EEV985Le9cGo/G69YMc+VYKqEZAhXYA
vvVJDvnGENO/kWCaONITBuoksglhBgh3creWhGCYIwzG0i+kfuGQT74dfdJzk91L
P0BzPvkmLOMDV6TGtakeW1rmarfnJw+diIFN/75Ujst9zoKqLhmDL6OLqnx/7ymu
CM1JifCYZzLyyus/VdqpX40/zZ9ZhnqAByg0RPYoYlORsqffl3vZnikIedCBlbwk
LXWs28MY8zluxVlkM4+2j13Aw2X6dbZQrckoKEfLHkpcE33J1MRxEbbi6K1MFICt
srlVRdJLTS7k5/EFuDysHaoiEHso9Nnbe0ca3ZyjQKYhV5CmclrABSxi0Kd6lZbj
WNXPwpCNIyCeIBYdHHzHjyVJC6811VopIPufQGMGKEufE2zXz6c/X6PW2CPFy0xB
hAmSiB6eyQYW7D+XTzb/32zLKzi+5c1tBP0bAkX60igw9dKnASBKX4hWBiJW9RLT
uexXalOmaWO8sCJ2kpuN24hsy0bzTDhuc+wUGJGgCuCg/61Jai133ttWrSleOVka
HyYVbufZdXjiIww641r8HSrQ3tTWeqYrlJvMjvulmSNvc49XZnaXqIyvXL6jHuTO
R6PS2eQlRESD0w7e4PKGRLkN06FXJUeOg/hajjErTrsYuWeG3+MFeP9lV/92WaEK
2fXFDn+gtKIzVzdERrG0xD5hn3Df5AvNfEA1gc7ezt1hVH50CkFlZj1wdXE+2GKR
EwBYCbfDdMEev9k+/8/CNvLF4tDoLPN8j19GblTZKwejahk9qABLhxI9v4PNP6pr
mBjK0imPYIZgeQkuJ9++UTfJEOw/Yi/Ctl1y6ghddX0lTa5E6RPxne6O/WmjVxjU
v5N/xWUt2ofQ8gVc3xX8OHbE9rVpJX1/2S3ljtngYQgXF8I3td+3VzIU7G6KPYIZ
jgf458yMKqGAb8tOcFVoG+YktypYKk5LDl+w8LZzf4gC4oR0Lbl5dJdoHlPc7cvJ
8OSsKIoiJTnJAnv6N3DwZbMseDEFhgJRA/qGMK2/WtGIxLc6xB70Beet/WPFcUIX
WFFo9vysUD9m2f4ppIp1S+ZUU+nguZXpbxj10Tg3ceSroAkUttOMTJzggNrxvgTk
NhHsmVXiXwQSppIFeX1zU61XQx48Da9MGSYJYrUvy41PBja9mSdB4ETccui6Hf6v
XBogkLVYy7YOMZ8h6i+HbInbnAIRLLk+9DPr2XbXiLzzc5/wTA2h5bePxW/UNfs8
3U+qwKLUzp6UUIq3lE2pMa8VPbZ8qixoLfm75PVvjIaiy2IN5Xw4jRRlwwBvPCAK
1K1+EJ02Od3S+bBqn79m6sLsyqCOf3SILfMJ7T21NHna7ZJ5vjVs9hBJ6USHJyQ+
UbmTS87vHguliidFA8+ouO6Gx+JtKrmHXj2A6kAv1swPTxRydF/fUxGeJTxPBdPl
5ARlQ2J6Xfre4xy5AzoIBP6yrzgYBPv9Avka2JU/4w9jG/AO72W0zqswxH5eMdwN
wPQQmrkW1nx2DokCFPCrVFVIapKuG5rZO1mX0LRXpTwg+GVsTAXIxhv7klQXYHHo
Uts+JO6ogcGI/gWD3wo74H9LaG3d0L4S/wjzYXBSCovKOguj5p62FaT1r9qT0qx4
SsiVswwwOPaachvBKS1QsMJg7WYbE/VrPU3HprDPXH7Inu7zq4QM59Aq3gtzrqSE
9tyT+GxaQtfWTnjUtgIn2mc1pTxqOUFquRSSFz6xvrblZIdOjT1a8aE2SrDoOCPA
C07NhkRpDv8Usd1QAiddQav2dFwCpERGpS0CjUg/O5jzR7zyOw7Vw14gmHQV9HfX
6jxlgxAeL+T4ikFuwlT7Y9KY1AD7k/P90Hg6QCMu6+BtQH5hmjfDMHLYxpsYxbs9
BB4oEa49QqE6XqMHuz5DETX9DlDKKfvExUc6Gyku1F+5WqAQixdEyKFHNTqWT6rC
L2lk6JS/bHlA+ZtCKk0j8HeI69KaQEno34IOozQhHDmIW/jfh3H/NDraNP2c3gYW
+CutqVNpCd3RorXXvb4cIlhOQOkU6ybn+m2fdoMPxhDy6PkoRIwJUe0XcqzKdAFW
X41xstxD87aayIe7xxs6CoYB5KKV7/QnKdoxqHubqukzNQCNVev7Fp0MsA/ObOcs
dHHhjcco7iroPSz2gw1QIeVKMewKZ6TPQHdTq8hKL9EQjj+STK7tn98UROIJhBAt
fYM+Mx/TqPJCJdeI9Nv1Ec+rRFpAGJHRZr1Gbg1QyrWKNuS6EC6sdJT7FjtTMkeu
dgj79f1OsAgMscPQA1xREDMMoBX43t3t/UeRRc24kNEHdrJc7UJL37/ilMhg3bTN
4QBsWDKw9eRNO0LnTI9/ktx9YBF7Wvwah3uQmfHKCjAI9MY/hT7Y6IQOImOmsAXd
kkU8bUsMw7ytSKszxVsN//FQirrs+hQIvJSPnw8FgI+lpxBgczkeMOcorLHggB55
rUgMcbfNkjtArSre7k4SNT1JOzRhLlEybdUKmaJLYauG5W1hMLk0MqVspJfveKTB
sAhcq3DpCZeN+uuV8J+oUcDxuj8O3sBYMhtS7Ze3PEXgDcjdO5MFEc09nxWBxzE4
xqZN7DHBD9ispA9PB5/eT1wGOpCI4oII2EnM5QvumtMhQhIs5seIh+Oc7GrH7J1W
fcb5emKuwaVuUqNJ+o2b+QtDUIG2FCkRFhYFFxCPYi+zy/dAiDFpVa7U6PlJivkK
sgsEzDYq1eiHET+vI3hKZCNeThNtn5tR/NwTrr1kArPI/4Xesa7/HJVXTI11HFvy
J33j3mgwBlYsnx+C9pkzcp0lbcz8KIJmntPhRvh4ouTgY6+hcuFsBIcpbNUgP/fs
KHgIfQXV0Pfpz1SVVxUJ00JrC6zLJcMs2Lg9EUA/T/p/LopRrhNmuPpLo6NZJ5iB
mPK1fQGMymJ0SGsyBEcWab3HRzJ7ynkY1nCrTIMiGwbYIZPu7N4PM0KP5oSTdIWk
IC3c3aSxJlrdYVnZ7VIzYS7Q7yhYmWnOztdjswAr+MosRlnhYzuCnx0FwXCcfdab
ydroU89hqLHB1b+gTHSGQVLdJ/t/qb7SKlXjvH1hn85wMrE4x2Yd6p4OD5kXzJAI
q5QSt50pBFNNQM+dl0/hnWuyfUJUmEt6WhOuKkv2d8mOjN3LkNHI/LbZfXVCA0ZK
1wOVVpMxChpG7tbH4NxHB8ToEOe0ZVnxpT+RObGTXJCX2I5tvIHIdoMIGbbpDEq6
2lJ1WTnVm8efikzhZsTtA+dfb0lE4SASPzWHa7wlBKNcByzt9bh080iPIeuaVu2D
pHhUG8923xFhh6XJdMGNScseM4fe6dXiqQ9WATNg17d5UPMcC9BD1ECYG9ZrIBSX
+arlT3IofFPA0zyCAKnNoqogjdSlhaAct4DQQD5P6WWSqXc5vTMIjZqU1mUDXiUt
zy3wvdCVfL3Ouad2yNaC+1EvUa4JOmD5V05YOqq202CMq5ZQL75Ixsf4NeMHcuRA
KCrLl3X3Q/3pZxz5NBCMvknooJuAMyHIPw0Z8xQGzIiFIJg3BCd8Uzbqd7rEAcB3
TG4UaZLqDdQgAOnjOP909ODxnfyju9XR5JgiAPTJ+9x9J9nZe/qGbRvAL7jQHs6i
roZntmvGdjR2N2jpMFP9cOQFVtJ7uEk2tawAL+ELfyJeawDgW0vaj2joEO+GfKuQ
FzROd2JCMA9iYZVXn131K5UB4/nSHl7Sk+hBKSuIxz5OOj10XvP3/fr+5HOSrEmw
SAvQa68R0DnWpIp9GL0OHnuHnIiHNATwE8xLMfF4s7q+JtLTBgr4/FI+tT0vMndb
Z9H4j9FFfFAevQWJNXd+8f8xEdfdcOa4XaXwVFdL1yXL8RJ1xuaY5+zTpuhmqIEG
oyTp8JePcTD6hrggbh8MvXyX7PP/I3dhbUfiosdv4cMqovPoyw2WIuobIOyXVMHW
LZlEGMbVlebSWgPrPLZFfxFpccPUFwxHNBhtFOos5d66iG4mGQYEl1F4tlhZ+GVi
ipnvcieowCfhZcV7QSb5zQuRzwb4YP16cm2gJNtkiWcTFgjKD1mBli96oV6o5le0
8wjMwQftopWAiQdHLJNnLEGl20sCACYwekvo7SLJU9impmfOBMwA0EVH7jSVx8sF
Y5LUTAxCdKHEomDkyNNPKLomulqmJWURny+IdsWXu4qDVQhjwRiMulsW39+HovD0
ckAeylVHgmtn8Ot1oBtm/bnlYddynVceCIROco55yfkvFsEZ/psB6ibZEruBF0uR
q0PP6VtkqRp351GlU1JZ6VGc5kvJHkNratn+yTFWQKH+9EAE4yK5bgOwPDIS6nTD
f4HZ+nRamSpAiGCnxTKo4JeQIq8zirlT9kQrmdVVkbw6vB5t4BlfaAW8e1Ep1pWb
tIHBJu290Qukxl1ZlNxPxO9EFlXFb/wUH96kQic3uH8uRVVmTo4S6Kix+kVFxAaq
hNBHXJHdRhi7BhW115dfCIxvWY/vvd8hd+vz+xYgLYU+NIk9Ws3yVlFXl1dVFCNw
lvGDJ0f8GGGm96POSVwVzvsylqZwtpd92LJMYWgL+BD5kqwvMvaI20N2fzD0zgyB
+LFdbemAPKk5zLdba7vapDIy2LT+qMiInqXfKsgimzn2VYnoKJzEZG1cJCOzV3Dp
I07wsgj1dH3BjvNHUDYEgPMt6wDOPnSTI6uJk6zJyP7pyy2RSjcE8uW8qS3sqenV
4Xt38cVMFfJD43HVGDDwhFI437f3bYiDfqiR7NcZGkI9/SB0szRyFaDdkv061tqg
bzyFME7Gx2u8w64jAz/73oeIEvh1D+QWKIvvAK1eoZqvWr3uYdh7ezAE9m3awut8
xTT1avhUc5vo6mnhMgvAVTyG+glYJHhHIED5bVC+GtgFmplKi0Chju/UdzB2T77v
8VlmYxR9BbDJq1Nz7XvW2oakb4hp4YEJA3AZUJ5SgfdHlEoHya/KRWoPpTUWVlOt
79rMLmngws1u70UkRMKCz2c+AkhXZVxarEVjEvt3eqAlg+DJBtotcnqdSj1UPyhO
IodCYARgqYycD1sw/L7YzEm9SndJyDNgOEwX+9hmmAZrB4keZrOJeU0lJfcCCf2v
QkKpWx7+h4xSaCnwuhYP+D588kFKQR7M5PFHpnT237xyz6Lg3qjtoEPxVctLivpm
tCL68jWnBT6I7QJGqMftsKcv0R6cYVbkvHp+xC0mkDr5kmDKIVG1GW2jzNU7r8tx
yD3jWJc0srJcjMw9cesDYL0BIOV+a1l56rUXbZhcQE4mUCmjPSlUIPmiLLVhyCkR
KpxRx7n1s7DL1znH+4q6LJfOq1CZi4NdtDUjuKXYVBujXzIKliqAMq5aXQIN6WRn
Nm4hUS4kb0oe/XjpvptmMURiu1afxtGcjS74T+ZD0uBCvQpkJH9YkCsriPBsKIps
7tOyEd6Q0LL2BEXfw9p/eyuMPmrEXKJ9yue+fxOsh2K2+e0kmibz2tFv2p4/jrRB
IcksJUyP1W1GIAPIMXfeagiC9hqz9UmlnedUoPLquXUJwHjr4+qzf4eCUjNhoRWM
5fMXRXtfVbTNTfhI3waCG1CEEj7tIhNKH1je3ySxxLpAmxzWsIgIUfQo+/GQF1fl
O0UWBWHFoghuW3EZR8qkgeh0Dtdm9yviypGJA83zB5b8mwn+OMb/p7zTWUg/yJPr
E+upWQ/QfMrQMQMK5Ia29ClYonPImm4yt4juruOXs/KxePWrpfCOqZU5TvfYqmTo
TwGc+qmGufBVzkRrht237+Qkx+3rRPJZ0UNhXNexMKZeF0qqFQbwcox97/B+zcVm
r6/7VveZLcIoGlJIQm409dBLBranSwMFg2oS6l8u+5cQAYGPOb18T1GXHlHZrPse
b274ObBNt9jd6huOpKP6IDGawUEX0Q1YGpkwsTG+L8Nm8S1mLxL32qDFpTlqRzIi
MLcXngLJNf0T9FVwOi3Onb49bst9WprBzxPhXrS8pW7a7FpFiGYPShPsFgiAnawu
opTRptqqMQ616pPz/VuN6oLzV2YBMzKvNxDiBnPoJObuoDqtVQAKlMg0LEYIAD72
nfzEReRbMMXfPRYFdCEtfgVXxjqr1oz8cTVLwd2QT1YQHN/VpPzM/H1M9vPclpC1
Iu9PNQB3lhxUluoRD3MhfT+D8XsOQPRED0t8ByImgd6q2XWNQ63gYgbEyEJAQxez
QFhTuI719DkiyIS/D0HFuCkukrt0ynQ2iVpZ3ph+iHkwuHZ7zGiTyZ+NMlNMRDun
+17dC3iaI7kDBi1aOVxDHk3C/kC1KXVtcpKOG03LZbKLh1h2B3kuLEIQ9K7nNFfr
8jusdlNKhfBj6V4JFdTCYaIviGhDlcQvkNS7+2kXmt8tYn5QZpPCVqNIKoU5G/jK
Ixy/rPJM7xEwsXyZv3XzWmcGAygow9LR2HbmZACT3ALn7/q1zmhNfhxXSs5m/FH8
7BUQbCUjPjOI7EcA44E1DyEFpjT02VNVXRCKly1+gcEbTmeey8y5d5yg4RSkoIn2
G+hapzi7YZ3qqQAvBcQXggxsmpCX+z5Bo145EKoY1CB1ZfChYOOt4hGGEcKdLu4M
RBHrsRTvpzXQMc7/1LD3fdN8D8uBbHl5TOi9a7G7eR7nWSrMNcqnFO1xuBfLyu+r
rxRzDVviDwvaV0d7WCnBxN7P0gRI6S95JwVCcsag6MRbu2dCTYApxcIDpiVzojwM
iJPTZ+/ZyKmE209VpyZlLRBohN8roIooT9jzboXnDY6N4Dv+gdi6m8mGNdeI9TaB
r5F1nevUgWPCua2h0wn/HTEI9mIu9NNhqxbXzihmTuGZIFoIoi9y1LuqDUQMT4J5
xgkBEIeUbBaybCLtbGeMYOM/nsYtKh6rlNoOHxijMh5s+J2Wajn9ymeQra0vtz/y
aRmzA1oxghA7adaEkRB1J2lJOOoBQHwC3fb+cDe/WumLNNhI4GVEQ8xG2p3P+/4k
hMft95qJe0N45mrGk71k09ispGoMLkK7/hP0mDF64pMvi2KJmfqXq/qx2Q4Xv342
B82R2SRqm6QJoNBHPkbjsf2kRrfmO3IV6hE2uCQCpXqQN7+JuTkFCtV+zTQTp4L9
fjdSxFegp+i5+vfb7bvDxNFxqMKEX08aKnkRjpAZHDStStLKX3e9CYNX3DfO2Hq/
f7mOhOqps5EnY7evaftAbDIefdK1JWOu3mDcCqNTrzXhNu5qq/M/3YSwXyPVZ42S
cAro2ghT0c0m1NF4ijkZyztXDJeJP8kp7/nxYJDhTcqqHKplXSpTUS4h59ZXvaNk
yF2uZVGoiffc7ZAIue4LsyVZ6pyJwIjhL9wXZKkY3qxiWtYLecltK6NLdycX43G/
I1+XBtS9jQ56RQ5sqP10RobsCt3z1QQBWw+jnDx1yqXxoAwk86f3tPUmkBqf1oMw
/XMTB232oLO/COLo6dl8HQ2tgKIlWA1xI/sht3NSSV26w/H7sNZX3VM2YWEIo6sx
Qdepzd9vXhjugV+k16XAttVUwMw5eDJYYs7vrFx6Pl/oO6zwxbNmRxkOO8QCiK7G
IDscBalkd1abMrOLA2WatgNDAzaNavI97Wuxtvbx0NcFxtV3c3PNph5G9zRZOQVg
jNA+n/SK5oXbSiZMcE3hz43Rh7w6oX4/hEeKMYQAov1AcD3YScMCqDZQuQOow+nd
aieMl4dtoNeTxIdTIxXI0BOjzFC6WXZwFoGuD3qzDXGbBG5yFuAu22KZId6HN574
Kr5Cu8f17yM7FKdc6JHUdI2zOkM9d+KQyY0tqC4wvCmugJVqacoHozuGwCjNKHdY
yjT6wQtivSeZPot2vER4fKyTc68Y4hQflgl5mP+yXMWlbQtyrfWIzJsgreCMRRVc
0tMOXZNKk+elsDl1ghCHKBkr3l/nIBYyt3cydj6jW5LQj4xLJUBrDDE8i/1yn/R7
IqpxJMMIZtJuuoHmvCIh73ajuembkUP/YC0qh0HGrNhFZJPJC5TztxfCYcIIgZQV
iMIzDvPmAn566rXkbPcfntLOsvStWlLzZxaYg8qX1xAvOKiUyqZd8z7aWp7Ua5Qr
LKjyX3X2jyXDJbLeKXfMywKMdIx27CzROcmC9WkuDmt8PR5xejVg5lV3VR8m2Q4C
WYe9oaT8EXR3zpfa8rdYBoRPWdU55APXCEkDxM4OFbVRLm9MU3R8o5G/ljKFBc9P
7BXQrV9Wu0e5khbXdIshSRrFEJMscby7NCn/+C8wDjjs4QDXXLM0JXdU+RQWZOTY
ZxtvIfdPrWi/Rk2xdbiLdnmcwxH9vWXN8IHe1yz/xUJ/ahJItKVg0RJuTwj2b0rj
thJ5LTNT4MssZhpO8JTfbLi+oPpwOfdQU7iHxXZfUH0XTQ6sV1PLElmm7ZRZOg7j
GURdYV4FwlFgQOvj6T3NDFgXGw+++JpDPir6Fe1yiMTP2h/PvBmhmITliSUn6RCd
grurTtMt4q1KW3LP1yqWXgDNuQCvcQeW+UVOUHztmIo9Pse5Mmpykv7fwwIxfHhu
hr/2Fx7wC1e68mB4sjscIdzwUr8LXHjzbnn44LmQsrIOnoJ4ZZzMGbKVY7zDbtk0
zVcqF9BP+OEKnG5IbXS3FnDO8e/fhx+lPxDaza6RYvrMYdlc80lzEJNbZwZhkkte
aOC7QXOPqyMsvEzx7H3dRSR6n8hW2QGZfaLLJ4kyiGt2nZzaRfe6fePE/KClkV7L
heqek0Z+gAp9pxDeaquTms8kyHpqD5N9Heh8PiuKdkQedtnIJZzj/w1ocU5oiH5K
LAKV02OvfuYZBas9yNinEgCqs/iz2fk9tuQvD5HfcV6dx8jFxOmnMQw0jgh8Lx6Z
BF7OIvcszd3DzZIqCunSk3cHXyYQAkWCr50CwntqTN0f+R8ZFyuIJy8Ho1qtjFi9
LbWdIZJ6th2tnlXCvYRlElBD2m7JrvTHfIc2D0JP/NWl4JDd7jGi4YLiq5na2GBJ
tnNN8/AIoI4QP/99QgpHgOPmyw3Yj7ILCLFH/IkiYqQ9DD6qd8gk+tuMrejnQQ4R
6SSsnzXU/LEEpvUV38Uu37D93zigoyE040CO+jrQyHEy09P88SrVT4lLsKedOlVb
07VU686g8OwKBzZxzl+3BPQD6cgvuRVvgzbv7Sz+56dz/TcpW5IW6biKGzYDNLvX
G+V0EcWJYtYircrp541ODCn4AcewqbkGL0txiFJhIu5gsBsAxRK7XWbtvHG/arQw
9BNOl/YhV3ZdeTS1YDdgLTxKSUVn29EZHfCibQNZcG8NS73HO5tuLlCzET34jBvq
Jwhpg4BDUi6MTg1wJBz2rNkJyjyKLfqwCOHdBjU+SrZv9wCpVVmMgqj85NE2jhAX
EiVzwv8Ftv7vtC623avVMIKpZokF7CRigfmlYrhFH8m/p2qrAtvTjh5faSzw/oLJ
5R5dUy2dn9T+XmB58eHGJ7YX2jJ0UhZoxTgCY1dTFRbu54RwEgFHGNIwvXHCi+kS
O1bKCUkqgutIJywcf+VAPNTNUoelZSPCJqAsVRGpE8pK5hXZRWTSiaPvYO0/LYzO
TIlJ8/qP0tJ0cBkZ4tfOB5boRrb+MkmKrybyF2JxW84RNsIl/Qm2TyGdIVVUV2hF
ZLsRSDZp2hiG06atXudOUwtIf017c5U1D9lfmoJDsMhsdq6hbRIdidofiP/2CLJ0
3Ccf9JWFZKgEtCkekbahCUXSg2CLCpvvNLP4N57lqTqa/uplUj/f6LGrxbsR1zq7
qm2kdYqCttqtyWcDeYoW9S9QyrCKthC0/Lolw0JXPocHQhJ11YTmEzQp4gPu3EWe
xjvgiEtOgmsW2dMCiz7l7yJtAFbVo5XVpFHVLQ+SBJvIfABzeDHzlsSdJsYGqrIF
ru2wSPM8pMRVTNw4BlrB1DB2FpaiXpaHNWA56rk38eyM6yhT2wSBXG2rnqezLRi4
jQ4LG4Ec7/z34wcXIn4bFXAuzmLSeiW3voBAHrW1W8xuCJ7H78X+4W1bf6W3z0rx
7idszRgiGuSNVN39iVflyQyXRgvKBskkaL4yZKueg/V1jAr+jbeO263cVuvfcybb
uyDTzOM2u+5X9ODVg5KYlRa6p2B5Gd2mMaAcyUPR9h7lPcE40YfQXfy4rvySba31
J1AW231W0wdv+pBWoJX1Ewk99ezEtu9U44zqdZJY/l9S8ttvZE+jtcOJa4q28RzD
4BP9KwjATtfPnRi5Fsm+yiL7miZYhDFF8RNxbN7D9rdtSYcYKzT6PZR4l9kF4zHf
efejw+GybZaruazBPjQlnq6rFn6V9FTFTq1kz1IbqvhzDGUVsESNrEljVV3iu0tD
WvOYbwnrxMXUcIGQ5ogwnG2c/3XbKrDNlDr/PtLncgcvzNzvZQSX7FrmahflOQl+
RaPl/iEigGLeIDORpzXdzuDSVPtl1GxvrAAYf2LWu1EkSA+jdEFmGFNLzi5qasbZ
ojgHXKiNAfbeChOlcXmKeHjXNpQ6weaQC0roDN9wKy3due1llA6Ul9kw9l4j1zcj
IYBO8LBvAo2mcPnP6OzujSWxJSzyvDA1Ib+ivk5tnP76AVBUky6uo6tgu9nWOlMd
pf8drFsL3D7zoo43fZsdC/m+gDPa4DPk13YjTwxiYR+1lYkL4Xt9FuCNoqq4BuRY
C6Z/y+yn/4baZPJcYq8yRvpmXhISfLj2hSrBj5J8yVlDbBbl1MZ6ylvpdDPiemA6
RTQMtDWT++T7wRsz7g459TyYKuUiJ17RFEMpN5PvuY41Nt6P4W2yGbwv34iRe3yl
CXuYTKNPlz2MvwSFaUvOsLgqtAmsIyDqhwEK4DPI2SV9WrfTPI9bRukiA5J3TnPv
up4Dt58Adbj/SeQQeCjzpFsxRa4Cd45Zu0wWnxXEEfbx0hfvNJGx0M9nzZv9JQeZ
i1V7i/goHYubiLYyM5j+14cLjRs8OtDsh9G6Tn/740pUgsDnipXzdyXcrityrK0B
DDlV3boGRuaPSCnjah/kBrQ5yhFYQYiFd/QOrmB2j93/Fc/qLUu8FLyT3BP6p882
hlEMqLPDsPDX53wQNdm/JAxL746+upeCaDF+B1ruZ1ZFq1vRTS9nEkpqksOeYR7o
px0kQlEvoiaLMTL3rxQSgiPcVzcF1SattqzkGyoWIh22SA0kLVNHdxcfWk3csz+a
kG4Kq15OaTew9gn4nov5099ue1MpV/atQ6PUgwbLMY0Ao7qWbqbDtDlL8QFkz+F+
wEtJt7Yrbc9CGMR0pAr7cfviw47kzitvnkeit7QbK38ZQ5QFFR0v3azA/T9U5pif
1OF+imFgSaaJAtIX7mrpvZPZQsEHfmjOqhn0li1HzvwsPlHDNTTcC25Wv4r/Gk+A
5V9u1wuEO/BNxf1Wumc669LWWC3Xl4Zs3OI0TPrG04EdV/bZv77NDZeOh+MLxr7q
voGo/7DEfxd3ZGhKOnwCi/zIojJixlqo6LLj1e+QUXDE7k+TcRdoIZf4HNwcPLiB
TvY6u4K2YizdAHsiNdWCPfdkAeQ8f3a4QEZcah9w9Zf13G5OrmjrvK0byxL9QAI8
OK9w4ebrf04hNrSghocSKtyMvsXx6ef2O7BuKT9CB8eZUkBUkrFavZhA7ttDZbQg
SVP8W8O9iY7fZy0FNycgCxx6gci+Hemf5+X7HLWpkBKiZ5zutqBiaeosaq62hZ1n
SxI3CUwkeK+gky0Ck6UZlFyGHh8fYifqpBY8On2jJlf8F1sfq7BQi8EvnKDFqrvI
xD8tNrzSEVHXPnsWp76iB33swXDZBr6bzaLXFUVcLTeMKEwkkfs7QrFYsFURG4a/
KN3GqWA7yNH8ZO2bBTHT4RFfqwMJJPYxo6bzM+mu3WsktCv4sTm/AqVf9qUdklhL
WJRgYzPxVJJ0NJc35FLcaLMbsO7ClEBCIOADP8ZgRaNUuJCXKrUsiqQN9zcCeRJj
8UXLTAKToSmChEZSaK0YrWLXZWwIzxrsI6X/oVI5sBRsCnKi/EZH8UYWOJr4vui1
OTfGEVmETcu/itawAq/c51xxZh6Iqj/v+ZST5+kgv0CY5ymZ/yn9idbKu6Xg/VKV
U9SyaRWvbu1TX843ke5px6OOsfEDGpRH3ooDW6rwHgQ1mdY7zMOK/kw4uzizUClv
3WLUC78LeLRW/NX6sqIfAaP+f9Pb1jWNR3xaZsMO96kPmLkKVLrTiYhC/WfO0waB
B0nxIKWQW3Zp3GSkQmr7MVlxz6iNdFq5NFdpsEpFbzJT47BI7prxBM8MrMGodZBP
foa1DvtzRrxHTee9Gx9TI1EB7bXjazQJozsj/GesrVVUszRTQrQQ5Rt3mL1/Kv8y
PLg69YIFvmAOCC299pU5ggjoYdp5W/P+fKW16Yf4Mr5ot1bdtlZXJ4ZuPl1XzW81
QLfBaPOeAgt6ALQGyPkOFB2r/+54FwcxBfyIgS0q1JzBJ2IF8a8qL95CHnearifK
jXEOYp84e9XD4kj70CeWNkaYns427K06y9EuKlRmqRcqlf6zbyWqgL/9XVEoaBlp
Q8/iCzxXrO2LfNJnCvCYb3a/qt/qR4zP54dr4fAHsohxfxuLdX0OiHn7m0iwHr6O
dIRis8tlW7U76F3tWfCVeIgBJ1Z08TPIhVgr82lhLunhRiyFHYbeZ8hjljGLRHcn
OlEsSTaTGX9WAzTpEfN+B3MlvtgUtIln4raWUEfHMoDvU4D7RjVPQZOXZ4Tbx2Sc
v5IpcdOlHjsA9p8lXkSV5KSuNia/fU7f9JayOxg4enJ24bt6rUkT9HZt+UiEu9uU
youfyrgSGWTBOzXrDekFeQDvCKCzrW33h0GU4ziqDSBdinczrg/Z41Gq0FrTMy93
MU+U7bJxt8NSM0JfKAMlu+vgizOqWJpk3ULJ+tQw2VYdeq+JLbR2b3ZiMnbqrMHc
WWxUn94oeByVnr6HJR7j90TohK5FbhEBsUQ+JYyBDBo1DredVnfm81PRBa5EYxJU
pyt/wKlJt0uSK0ZyOTuAjfR7DK4FpsMxMYvB4NQSVj9bL/3h8akYZ/GFbL6Wc2jh
O7wAnfN5JkM0n7RD/mCN+sPDwbLXwqFr2vjwh3TBt645i9JVis3Z1hIriMd6wIAU
RG08sAfqlCPtej6XvazYqPG01sORGF0lgkMsxSHQNtQuUZwxGKZ026jxNZiYvlyv
v4C6rBl7gitiq97Rj6MT2IkgKlp4mMxiZFm6ONNl1BfNBulqyO/RYV8N7iHI3qtH
StltfNYjVFVKYAbALEokrehe1rogrYOPIxsuMs+aX7nYJ3jz9n0DrBepFO1KWd7l
10QymCQcc4TMI8b8Ng4GkM7YCYyWRV3mWHnbGLeVHjq2vgnTenU2HpJ5tOMTTPQr
J7ys13ifs5RfOF2n5BvP2d+9MRCjjozcNufhH3mk6lqPQhc5Uur7FTLCV5W8Q0Cs
PPy19eHKkR8VnYLgYsCeEDLzau+XhfKPrBPMm7vDyjRJZ5crQpaXxQjms9fMMKtQ
ZQxmHvcaQ3IWQN3HwwJkHb2WXyr5Uf9x+TmKnXs8yyAl3wEzm7uRVJoUDp1AIAO9
kopZhuVcXRV1FaCgCkxim9vtsMLWt/fy3f3lyOnkwggR00h4X85FyDEFgqeDgzec
53VEz3ZXvMYHLYoxJohEer1mYnISpnOGJnHMoiCJiLsrOLdOpzI78RetBIZMkIby
ealCk1aObv3xRy+YoHouF5eba3ikm7eloHxI8KVR8yDFAyWvAFovRS5AHcm9HyoA
3LF5Om9Iv5LqdF0MLYBuvcvbaU5ddBaGm9ExBTRiSHTUnLD7o5OclRRP0T7/rPly
a99ilMm2OHiF+G7BC5C1KXwRtwSWRgX5cjDyhm5ESlJodoX6LGpehdRldF9AtL6F
fDSzI8hTHuNXkFCm0UY1QjyV1GgiZgwuFEVjPfztv4uFTAEmki3Dzk0g9GjZay6w
p9B754TOPrSFUHW2o67jZ1NwN0TNcuXU0pbZKnXSK1PxaYs5CcpdWaOaQejPjec2
MwcRc1dbucYFY0mxciAgZ/OlUCaANiyhQoNUOW9Lj/ycsjA101YdeRW3A3N3Mo/g
68UWxuxuzXiTjNz19BnFC9FU45QgjWvsLaw64qiPghcLMU+2R4P5bf7OFRfRW2H1
w0pNfmBMIaN0WCTGRRYFCe8MhTmfq4w0sdnZDsF9iXG2FjlPacWQ8n5qwu4HRPMK
CByRPC+3MeFj8omUGCh314JAKUUoRmHuqrqS3t+Nmrrt0fmi+2Y7KbbtHI2NUbB5
xaIsD6yVO2J0Fh4muWI803cWqV1Jy+fBBSeMU0j03AIbwyYcZMmoT/NR9VWAfqAo
qGb3kgUCzojbhfPIatYYH4WKQrGh0s6Djl3wM24Fn1W+mc5iqDG7osEfudKpL9zZ
QbC0n9zvstmkbJYPhLyhKCst5OxIsPuLTPHl/CC+gkSD1mq97wFEtZtUZzcnIp0K
7KggjUJXfTASXMvST5Rw2p/zahEFovtHuykYoDBo7cAGA2oDJ05PTlT2Sg3pu5sl
sOjTQg7wyM6G/yIPo2FrKHy/quPodnQ63jKaK2+uqvwqtObwTtDsv5FO1ySELX+l
eMQwaqOm7cA9P4Nuk+Rh9Jzeol7I5K1zXJOpM4//tclVD42NZWWFF4/bpHQqNXpe
az2xJurmKUM/97ZWV8RbWvVMjXFpvdW99TQQZQE9Zw5kfiXLxIdYvwDEt8PJIn04
gQG6H6WMuC5DsUX7qggHBrhOwO76oZXY/7HzSFP1shtOO8hD0buJTx5yM12ZGH6U
PwaRFVS6RjKqfQFg+A5WdKzqXV07g82BijvCQczhGr36GWpUjUqwoiVsP6WlFWd5
GUg0wSZeX6Rm/J0bOfqb0QnLqomwHCRHs9H6S0CX0b2w0MM3GAiZ/0FB13gyOzYV
jPg8gMqIw97/MOMyJz5agu8jMv0diO1TSFS+fy41nwsTaila8AHAYZl57zuz3Llj
N4lt6iIPx58k3ERXoenAbqCzZvWvwYKZVhFmX8Yb52RSlvVxGKl5ycxZUR81FJHg
WdPKxa1LescyA/jQmKnm2HD7TcNtWwOABmIMnyVKiD3Njz2E7QAMTBpk36IcCI3B
oIvAQYGlERCnGo1NXzZ+ES0gO46VUKq0SAVjoZn9hH40nIoVgKebTCJYYH44QfgL
hcuPE2c24qmysu3cn/c5LnBQwtBXm/jFwByy7SwVhxGQx5fIaNazl3dAvQF2kVtJ
5iYQy0BwDPa6KOmdj9YmrgicUez4NvBN9fKw+co/+3FkHg0XNQKUMhYnfmWgmueE
tJRNlQf6UjrG3I8+EEgr7Z0/oNVeynyugsD//tMXbXQAE0GUCxW6ixabtPwT73z9
dvk/82LpoYeTakjKlKBV5vgmFAd6LsvMd1M1Twd1IbNANUvP6ct/bKB+AswZfnDn
hJzipxVczxkSfCKeGptRlBqLqWUgOHFEN+Pp4lfPSKd6lwPJDYXBCpe5ZB3Iz0RZ
rJBTarvPqARgg+fivob7WRS02QheBdhgoZdgkVwDJ+oLBMjjIi25+xY7JcdvNXF3
x/TsKN6xiBLgG6e3/1uHJV5Vf2N+h0TlMOwkyTeyvAY0SDedj23c5tEB/W0bHBdM
67vVyoE28SXPTFn0DUUqfzTShPgf5BZMOzqbVbwOVghRu3FU5jesTiMNewpe91XT
pI5mp5bLk+BgxnfWYTgD9Qr+7wJ1IcSI1KkosHWvOF0z0lnUPgEOprB/ck2KmgPl
i3NMMi9bYK09ZtwLjBwkeVRQF6fpsQ+pQfQ8aG48/tSEbUm2fziT+GjyBv6gro2i
U4Ony4Ms4olmkO3nfGPILokIOwl78ESj7IJQ/CScK4hNRVXBz2j2zCHqKpa0OCuI
PzfknFYvd7rza5CLBUj+8xzXaYuivw2C0J4dxHhvUf5f8V9i5VkryNVRCevdMguT
jnmGKNlo/x/IVoadlljVMAEa8U76KRg67ltkwbuiUIJr4juhYdcE/oRshPs+gAuU
2Bq6DFLQ1b8LAHUUwV4MRuqGca6QV0tFcZFXZs9PHbHN19ZCEdOe3ITTry2Ahn4U
UguYI5GeeYwadistR/XdLsV8U84qgzKpZdkjRQlUId6Oftt7NB/ARZiqMw8JcPYk
VNNfC7/4IKAeWCejLg0GDBHvBoA5vQkDtVMBXp8x1WqwcYgzHZTvu5q4HdkzrR7x
rhHKrHCTlJtgvnRHtDOr0Q9WtVNxdf3SeOpHuYqbAvVz32GG89ES/7jcXC5LPk14
D5KaImUTHjpvVN9sGgmA5fmJdy0Cd7LDYNlrHa6nPGDS4PTDt6F0X9VjPfcdfZz1
RW3LIMr3ocsjOvCCuBt3dOh28KaLxgmtCcrnwHTyBackXkesEmIExYagmAbnfvEN
jU/HFtEE72b+BOyfvjlvbHsrjrK4uvUpB0q8D2qvEVJbzHjvDHcBIgkQ3xQmpL31
QVBMB8EQGl6IHsmI3D7KYFUEl5Z9MvMV9c3CNnJgvaE=
`pragma protect end_protected
