// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:05:42 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
IBV/LSQB8qZG8SKV+iDKAtV93tk9l1wKCZj2tLiK0oidPHHey9D70wLW30oIeAIS
F9TUhss2olJNCbh4wfbngm6GyYeINLG5gqtc4FLMVnxuIlHMIXm4bdBfgV6YhtCm
+QTerVVgLG7cy9onvpi2zb1Ewe+SZFnZFYhg3oE7Zcw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11664)
LrJIALJAMXkTNmCt7QXUANv+lC5Ykdrb5M2YDJ2b0FBvEA3Rph6fTm76hjK1LnJj
7Dy7KiPRYiV4VO55Keco9VE4RgWdXOSC8QuNMea/MJjRqINDJX6pJA7qmJ9llJDt
ADZBW7ZbjWeyp27n9hxdmZv+vicm4MxwtjNr+bmw0EV/vUVDyHVlIt+kkYBjD0rj
Iyrm2J3lr5dw39nLcgQT9lBJKnqTNzfovGCRtU8uqDUC9joKcF5DFbIFKvrmOpuW
oUTSDO5wHrWEPp8GQaG/wIa3DP86DWic+/6QqHZ0AGf6DlkiQIfqMl/q0s03AMrw
7TOAQttFWrf05j42KoXcCzkbaS5IzmXU4y2Khk03Dp9KXtIzSGEuwatyThxVodiq
OP0iD1JwPQmLO5/8TZfrk4MlJ0hkitLkxnZT84x2BfkfUt3FIvPdcncB0l5CCXDQ
+eIOro1C3KqtPtECR9ICOQCeeVhtRysAiFzq/xgwH6S7nae5bjOoMihaGErVq2Eh
dK9fJJWaVaOp0JZJsl3BRmCf2FsQXTbrGUn6RteQMCvKrIG+NzadK7Jq+hEkk9p2
yKqQaP9KrbEBCTLT5FiITkoPzM+cDv5Yp3XS03edLyuNspMSFdIhJtQ+sLraZY8W
1xs+H4vbbiQDVPsfo8V2KQ7mv007nLrdt7yunX2bd8oSS4VW2m6XxcjFLrxPxyGm
kmkppAZSDa/rz2ADSI80UoB8aaYGL+NYiM02gS957317FTm2zR7DqmIz/5QxRUsq
HtM1tjhE5oYIfqx8z8EC2leeK+h0aIJ6sKkBYnAnq0XwmAieMpXd12LbdaOhHqwJ
cYno5b0KDNVIDfWRBEWplPjjvOEI3Kv02Z69EkrIBqdxCWE8cGoh6kHWinavYYNO
Ps+SmI+6z9eErPEfIDWjNBKYT6d1+2pHsI2OizynpMmik85vYi2Stt+EwrtByAvy
PG7ed56qNg+tNRg/2ItFYhnV1iDVEZqRbVZZUAOhv8DfPrHNnE/b6G2vWTN0yb3i
FJebuxRhyn0QfbTNMgp+PZfFxsitL1Ke/LWsm9ykIXOMojXprUzmqzoGgB71pioX
VRXDuuhkVss18TV3RHvIWA31m7sBFJF4ph/1wwVPBe9qi+neh0NMAvsoUE4p98de
fRYZAgUXWWXIOxBMADONKQbNfiHaaddTmOCcuI5LSaHxqqW691+Jwd4gpwMMIgZU
j76eEgFIWNgE7IA6lnfxUaFoC3r0D65dZ9QS0jDyZ6WL5oZjndTxDUcvpMz/DjXM
AYN/IBe7EhljDAlQOzonO5HhusNx6arhyXLbmYhKOixTFbwtrhTqQhU73pO4g79r
sQLpI5x8pkR1EZVJtFekG5ueuiM9YyZlKtn8zfvvCkkuM4kNPMi5A6+XZUWVeL3Y
j3FONAjym5fXpt+vY7fd4lgPoDLMlfFtTeB0tCeoowxP9J8Ash37Bz1mrUDJw/q2
F26rOanQkHekuu3JWZKhOeuTHAti34wVxy9/AmctWov3DzuMkJ+PSb+n5KlPEScE
VxJhaRP800XSaWoDLqGizf78SCv4E8rNF+NjBJqMklXCV7cqaZveJORO7KJe9GlN
ZtZWPkdzAn8Q2WPrJaVOKE+hIcxMKGTSEgJMPuEJN4fTrnZZlEQPXIEJvcxYXhN8
IaHCyVCDuvjdQZRpCtr93uLZphI9ZhA7wnSkqqTr5uBtfvVlLLDwbnL4mN9iEvCr
OaXKWaxJl9P7TUmphEgB/h8PaUbwkYqirNxXHxwuVLeETeY1TrMX1DoeqZaI+rsi
9j6uxqDcxgdoYGL4i1hR+Q1UvrxvsnAFrBfyoHhqoXSTGEBoEUCQj0yn5L9TAbYR
M45rBn2oCcHYXlMdyAv9q/RTMl4WptfFCNchRuV0LSb3wh/0sjnmA2SrEqDeDOTn
zD2ZMoIj2DG1/1vmDsJ+kO5bqn5vmmJSCXMl3781BQ2SbvJ+nWQWXGWePvC5yEeN
e/e8HAyb6gSL56oQpYYmTnKISJZfSrfCAf0N4Aziz9XGYtZOqzYmQD8i/EJBYNkn
5jKofSgXe4v6lvlW5rPLHJqCvZHLCYBHiKkKGaq6jSnxbx8eVZqfTl1291xDSFqB
qVR7dDaR7sbryqt0CpSwrGq+wI0M2tp+Zzqd+3ZgtKFmifQrQJhHyOQ7o6wWY1W2
MWN9yJyxNYmHNwo7tThbfgzSta+4v/cxPdTUu5ox750bkc5rTV+cr1acrRBUKubE
5Gj6b49PP0TVl8e9g1tBtLwyYU1Eq73jjnlgBhEyAf7bMBdhXSx/PsHbXYrnUQRQ
MeQlbVLDc8+iEtl47sZu1R1LItthAXmPlocU8kV5LKgDGKm6dthTExBr+aCNpMH8
fDw0iawjIZtUflkjzePDGaxOJYtKcVkuoXANJnlS0W5HEWec/yNtWtYnAGJMRlEa
NOinHiq8RHRh7yvr4v2AXNrJ+EtPj/MYzfLWSZLGxa8qqEyYbNVG6CZ2KypLq5zc
2SREY/TrKJDndCTVD6/fPjiGZhKv5ROUVxBaUj23+OHFkHev1qP0cbDtSiOogxDn
t+VQM1mLXWBfbpT5DOCUYe6qDyZhZ+F/1mV5hfCmmVKKkIhKJEffVxLA8z7AlLDW
JOTICClmwTNec26IRNVrmfPIrmaN2pgP4296/bxQnC5lMIkY26wPR2kkWDccSJjW
p8F8YKfDfDDxhjHB9zjjm2l6fC221V5ismFLUOlev47cP16Uc5yXuaBqQu5IzUK1
j4/UmYjUjUucHL6ZeUVcZcWQWWw/VKeIc7kt0mjIAR5Kg57HQ7uBLyWHjFPIzObL
S/7VcP4s6KhHYcy2pmf7IkyVhdJDxHS7hoi0iGxOuXDOamj2wrk9OwiAOhg7ZBFL
K+ld0EmWc1DkzVT/BQxh5jgNQ9uVGhw9G9DxctdWf7VJlqOl6vSQa7vPvGJMZDuN
WmOcH8N2J+921JwFCEJe2sTVn/KPIGh1QEZLAolAlqAzcSw41YC7BW2KH4Odl5Mw
OJMs1mUvgjzyzGS5d7qZvaLxYYP4gEfOE1FpPMdNA34g2+JT+RM4nF0RAOTOYVMp
kN1MsfJH8SfqQemVCnOvevk5p4He+GUMMQHQNG5Wz4JHE6SrDmqdN2IoCLjeM3R+
uE7o/37zuG7FCG/pr9fRwFERC6iyGql/ZUWfCVB1M5UT6ICihCz/RhGoq1zxOT1X
d44+6HlBbwLF1+AWjXEyJW7DnrWFHeFGcUTak0+lMsqArXDuh7rPlp3xINv9AvOw
Ecf1URkSuuYVbU8BHNYBHWOb87aSry+JeDX11vzfilbq2jpcWrqeJn3fQqXw3/C1
NISoqjlnj3qU7Tn1u9eHVQwLKLkU3PbWUyZQT6vNv1rqERKOwtRQMQ/cTLw6N9q3
42DqW7iwte/m/cL+ubBVp7ZrsB/ay9yxt/LcyrmNsNZNOCg0UKxcJr0rJ/5DWmrD
ETGg5dAzmkHrgcqQrtVoF8Z81AwBRkTzJlQDp0ITmQeOlI54Dak+aW6oHS9V7dbV
GtuTlI/lnusH722RaDkq8uJAQmf+mjWUdJNPUrMSEdovEYXw90z38JqJx3WrH3mK
xcDZ1Sp2RRppWBjG5gfjN95L/KMuM826N3+w8meBdzC8FftT2HWmTwOJaxpq3XOl
hbHfFdx7W1tCgX1z6y3JPXr2+x1toNCY+jEilbJfBo82SBUAkV56/N3ULoTnWDAN
M+WND88wUSLyg1i6OL8Hvwvm3tlnKEZ6L89u5awXaKOwOzVMdKul4wAoiKMcS4uq
BChmRxIRGGYosIQTB5A9JXuoyW9ie6Oygl1rtWr4i1n1xABDmSBKpCwvBdcF25ph
mPKqXmbhDhuR0bDxxe12lMJFLSo4a3oXcee4MMgpVs+f/eD2wyBw+NWkRkGGvdGs
uNAsOsqZJZUxDkATu9cSygRO3YKeZMtOlwY1p7fyep0hjbJaI0kaseS32AwPtQq5
mgmQ4e+vIWOs/bQM6cCWzHVd3faLVPB9TmgGDD/H+SopQsTw49cZoA3X12fsyfHc
qQr807dMjiCtT66qRGXKSakIpz4P2TbtinYYc47zcLD/ZhwFsUnUBZV34CozK1yO
4HLlYwcj56S/i2x972C1L0z4SF7VNxMdODvMNkpRUyF3UjFGUJ7kGhju1sU9V8gR
P5gvLhYy9EzSlFKCpcO7dssVj/q6yTXNEOL4XfXECTSzPBSo8GKUB3w4WX7FaB5/
qC/J/ua6dH9BB1ukyHBjCOS2Z/dJYOWg2CyhqvLtxQ/LLJKPG22048IU7D3rn3/n
gT1upc+UpPLMXSJMUSAhdJOfQMfEq/r0fL96sdvwdXB1G7L2gu6+wDpjlpl0O1Gw
qTEcbtobLCvQnJL1lOm7eqoT5fz7iIyE0ltSQPbunpqe5PS2RaY7NL475oci3SUL
2K02XeMsrOnLmkWXKy9O0b7mDcMmR+c5s9EnivZwXMS1IO/W8qw1tzA6q4fQtsnu
kbINmZdjmjkFy/GqALQ/d8gVJga+D8XNqnx54ICWDaKFm0MuOZ/PhXkZYFqT6lBr
6d7cY+GA4ySMetHXw1zK7WNPgV3CmvncqOt+36L0AKCutaA5ecg9xyP3oCdIkn4G
5MTUK/3SJ/QgZ3/sAQxC1am6x2ivVergQFMKemJqzutt+4gJWxWmfjDvs2bKXeqS
FP+uhAJV36pHG+wQ09vPfDVcYXLlxTJbr33Qg1jl52l4U9oIHRqWiqibZLbSlpQK
S5A296vzEoIlaTk84ns4KJpQBWxbPwMT9ZyNuFsdWiKlf6oWMgEyZXx/fbTovjYX
ccfC6U+GFxzWflM3wCT00n3pVjwttk89XavlX33IvhUfp2eMMa6wBlkgVfOJi/rN
CgrmnJkFvvNBKHj2fdsBSljapiNQUZQyNCIaYS0QMiUszvtoQX2zGqBwF1QBopAZ
U/CF+H4TiinFXdiKqILSE553zoOVCys1Z2PM0rjnh7eSTFj8nW//T2Eu/Qk3yzYE
lWt00cMCN/1Xrc7ch7FXr1pN6o5veZz3VUXGReDtcLeLYS254M+iy6vk0d9fThQZ
7aIlKxuq2rbBowmnkG7qzpow7uXhcg6JtTO52d08hoCvJ3uGfFR6Nw5QoC5hyOsm
ji+nJ7+F6/iQ9Ap2E9Oxa/4vI20eWbdh9ensQ/b/0sClIVR0PclpI97OM2oGENYm
/EwG52TRaKb51fXOTvfAlmtzIg6CqDSk5H0PPV5wAPDVPlWdM+HgK9V6XO1s5DTn
aJTwn5xqjecAJjgN3ZFgMwn67zhPb4+GtxX9GMAOB53OHPg/owxMDUsivNoRpgOI
VoGppkG1BNawEWUnd2muzhj4BZT+puVHF+K0ctol2CKBXvFtiYD6ISh/7SywNgp6
X7qoBYpp/p24ekDz8wFKVqlBZtQeKY9DvaqjRWy0E2rb1Rc0igTUZuhh1n54lFXC
iark3YcItSnB3uTb9DAZsCl8LoYcyQAVeUNxPHfLJpRrjxscn4/T8xvcLmKxXKGz
X+SiH5kYs0bN2LHqoGuExSaJcxOUwkdHUXWAJiw5E7jpNYCO43mxFtOF9cA5cEZT
W7OsZ+RSQjc2sBxQFXGGOSuumYTykIGYCua6LR+Z7dWA06QOVrfokh61VDEUbm2s
/QXOfn7jCe3znraat039g0xmNdjy6VYPWr4I9YM/uQejwIVPxptfm7EnC7SePQBb
NhZym7Ft1aXNDsGz150yKr7LfH/4Ejbq/d4w9h6l65qZErJL9+mRrf2UnktA/nSi
uDYbuuiOp8Dbp4waJjyRjX9RFm+iFE2FoRbBxI195xnSlGwMHlEx46NNTPa6uYPu
ONygC1zeXvtruFJyV8KGm/uCUhhuKUC0O963o2nwHUOMOdpiXadPJHtnp56YJGci
DJczO8bLm5mH21kapbDRW00ONZhQW7P5AYkA7uRsdMIX4baArwyE60/K0cqVovPE
qBGw4DsjJgl13S4Jacqf90BK5ZwIuO6mK3CQ9GLP8gf60LmLTmJ178QSx/rhm4+o
3iGb1a4bELhpNJsVaWrjL/e+MWsx+7mFVBPPFpCJ0PVAQS0nmsNXx1hRZWcPiguY
y9KXcWW28a+o538aKHT1kOkkYN6ch4GUlsD3CGc9GEQ/9i6/mdYQAMrMCduWK4c8
TbSnJ0VjEIS4kw4EJ06rZqRolEXjO7ODGMlZ+Z0iemw2W6owdvlkdf7seCcV+RrV
oV1NjC1u0E6PVuWvTTGnPGNHvEAzqoHlHSEr50l7PWbZJbcZwE3XWK9VFj+jYpSF
wT9VfgmEIffYb3JI/+b7lf+q693rz6jUJZKPvweQrymxa1KlgZ6bFHwO+I2olcgS
4t0ZXXG7MuwxXoJ7hnoA7cC7iruaLA55K9XDGlZ3DBrDl741CrAZ+2LRB6M0+zvu
gKXpIR8lKSV5KGtDIO9xFqrwFo/6LywsQu0wKABx8uzKK2WHap+MpM4vlI3vTBvj
C7icv3TpcAuEpGt5ww0iwbeAxFHc0nQqj7EZ2HKlaRWYNzz0sDL3M1X/WUsaP3Be
KwWepqNFBDBARzmBcfRjJl2KDXR8YHPYB9+yEIdT9xIfQhK73MnsxDhkEpKK5Tar
ARrUdSWsJ3CR5hkaXnMCeHOPMnTyh3sVb0LD96X4QkDkGnYl8Z0EQB1mbgYb5DHT
gnK2zFPN6c/FuYgnkf85UHsN5q6PSnXubSq87PIol4C6DWs53Ga6nDVsKvOawzwk
b1M9+E2YK4dekx2eJrjfXOfy6aB3nw9Tw3H85W1ZokIuExDcTjNjarpTys/IVFhm
TcGe179ioJYTEaWADG1GnKv28DCYqdeU7M/hj+/GlVktmZ8YwBuwqXPU6I7XJ0jQ
VCb+h8tbemtzV3AWvFpyG+OKLtCOK46/S4qEATXUJ5eDKwIqR1u9odwn9uk2TBuV
Sq6GfLDE8/1TN/FvwGqnl6pCxl4k5Ty00Kpf5CF5NZf4Gu3lFyq9qWPYKkYhhzK+
s0ifbM2WNFuBD2Tm7XwQsoxqarGLknbnEUOH7eEkrFJgfP6NMRGz8AM3rcgk+PSI
o519fwWkbkZyvCtWpoCabQbMevBC02CeG353Cn7m3PCi2t10vwuI5LmXGdaESLT/
g5QbggsoF43ww6WyXCjZ6pX7GPQNBqhTLGLHDTkv2aQzlNOyFRs7ZPCaEZuEGJNR
eLtlwnU8qugjwjbBsdcixIzC+ppmJ1UF2LMbFSguTWK4U/Z4VMlcjeJp4rMCCFuA
355xtHSKrUxjlMCpCMWFwRSw/dUBGV+bYUCbThuHEbE1lXJQEUazQUm5hFkTBDzQ
UD7R9cwZO/QFoLbNASOsbEIRxwRtPi/4B5u5GAX+idLIWiMEd53xQc57O+rgCcGR
GI87mDxaY08cUTsfM/rs4sds8PVeXl+TKZsI/2Z50gLqC2X7Vo6MCwB1leo2WfT1
vafrBoFNfCUSoFuDrJScbeoVoT91dyqRxrAe30Yx8y1V3nVtz6ALy9eRni0J+DgR
0hTGkJkttaKY2CtIe/iRPld0UyIVfYFEF+1X8yBB4wI5jhEheGWsR9/M8iK85KWs
ffHRB/dDoEEZkqxvznFXR/CyW2y6CfDlsEC8Y/WRyGqXmW38aLoUYlRXknZKMFhX
shoq8r+wwp5hAsXj1jsSYE4AJ8vbCp54OlTQXB1A6QjTyexZtZh4jJEkDBSgJqvj
aN3Gd81n/JsfntnG7RlBLwdavTxYNm0dGYyM85q/EuptODcoFHW+3HpBFJNT2Vh3
8KoNtxgQ/kWYlQRFXbUveZvr7p5GBHTNsJzwX86uWeWecF0jUyyz6tY37mWNcmND
yVBcBhT8ZA+dpg3UhHPxbnYZ0jL0mmI7PwTDl7E0OdrPUWsBhLnl2Jzg8n+TfmWf
/KTZyuEx4TrstF9nP511T06aHU17ZhG2viprCLVWNUliK7MTnwpZtXVOU5plIja7
RHv8qhaorPdB7eCHeU/s6sgX5MahumPQ43ITNg8mIOMc3LuIXda4pP8u1MZJZXVt
qgEgMEm6KnlNcX/R/AQHnreSCHbbN9dJOPm/PVLPON7Ljrf3AYNKFbcu/5Cp5t74
lJ4iRMbAuu9kgTkUDiAMrSxCUBKB98xHVA00j7ioIjln7CgcgR+WnOY6QesSU+TF
6EY5Pdv82Xz5C3/UdJOE4AGbGyulk/dD5BLeN7ip4BpmjPrni4rLuRbCeYhzU/j0
bzmzyFiE3Rcy4/SlWCQVX7IPDQ98HhrScz2hlozQzaN73yCLhFJmwuX9aZ4rNRwy
+FNSX4yhXXKsJ/dc1kho70xz0B/l1K7owBwSdkM5gco+10rq7ZYfQqfrzHLGH0c9
oGESaqgGxgtJFndOiXWbjh087KCQY3nW5QfQb+bTt1yqCHGHg0VUuOZTANxk1Z0H
Dszm39EQHJ7+xHrwYPwiYhzg96u1IkJv3HYzneMZoc1xNmnbFE4KjmlhL5j5BpiX
x7aHh1AXnp3yMrSlI12H70+WaBwgTkiaABJq8BNU4NgCXXfVBR4cdFc2el4bHSnf
oS+qaXC6286D4aJKsgPRtUE34jJ3OaZ4OURDsFfVgCAJdX2mHmk3Vv/qURq+uB96
J3uTG+rEf8vviMbsrt6R8GW2cpsyUioKayDxDZ8RQN1Cw39HpgpHj23Fpfc9MBqx
K3nMaL6ih8UBBpfqTQKkmQ39K5kFoRWyT3286dA9znoYbkd/lABfTZGU95IhQQVo
uCoY9p/HwRYdzUQPvzLko+L4GBu9ce0P47MV8IcDu5hPnQm9uNQNFpTK8pOehZeo
4VexcP16G5QkJbe2h1TfU7xWGznrvJUJ2u7AeWgEqbqdFb8opkunigbTPU6pN/V8
n6QMwEcD1Ikm4wM/QpR/JQmgIfdGYAZCCbtMiJck7hbj+/iglzvhki7Rmlco7Gdd
ucujbU0Vco77m3MNTgEnA81SB7+nmU9uprqEJ2QduUqo2M/lkCV6HcqvnrK90oo0
C2SdUcFt/8W6dyI0MRKm7nlu9dPAz9N9TfeltKbZHzYhlF3/ppw/piN1qfKevC9y
p3SXpGQOKKwDEDZ3OgBUoFhASu+29kwPkH+I5Ja3eyJhI3P9wr/5FVu5kmHPDIiU
kxFlDXxVZV81ggneVRQ30/u7pqLD2AnmBl9E6BU/0GgX/VLx5i6vVn/sVElXCaZL
MEoCUuCDhzsNjGjAxDIe6XqwE16StIOOJKMge9SZOHmtx5NVHLjNA7FT1B2XwyB2
SyHGifwrav6jUoOkMCgVxXFtBWVCNv2uwJlzi94GULXtVg/B+VadHqaJhSWPYAt1
8KQEed5o4xHk7vrE3nuYuGc/6uzPigVAQwREc981BeIMeWx1uG13OzEx4Dprtrju
9pmANoM7umJe2srJvHNvitMhMndLvVGVYiEFTgSES4QwYgmPnQtJNrTJZwcd8XpF
YhKDTkaDKM4WBxIYf/3xH8ZmWfweEbNNRFrKSvKe/T2csrcX2VFf5o38fwOD9kmN
xPl/JRC1owwLsyl5DYBzTaviEyx7Z7F+amEVhl+V15O7uVQCrXHKxa7hzXR2lTJi
jT1HHPADegKVOU7W5S6VxGQygWsODEQZwzx0Rzy6qVTsT0rNEnjfNFgdjojYPOE7
ajof2rZ1a0rS3x/qAWLDBcjk8xQxZqbYnpVQqxaum89l6p6WWiB2q3XjqpfqGrKW
JuTnqUI+UOsgSFXigXwfyRwmpt3MkA51Ijo3PBg6Gqnd3M2JVO46Q+c3RgsOjY3/
2mg70e+s3CVwjirh0fUIzreH6X0gw/QhSK0kxkrw04TopPChC9t/uU9PB68bBcUI
dvSZPu5zw7PlOC8VbZjorHn2+6Z7GtdXpjGh3X4qzZIFcrhEA3n7eP5BMdpoBk0f
Dh5mKrTrncfyGS3sj1JnemsnWhNQ/DR1Lx6Bx4mDgtptU+tEAmHyIXxwijc7++0D
QA3M+oB1bCEqxoNR2s/D2ZpoNOhPX2dd9l2s3kmRI29f9atlpacNhbURbaK9en4w
V1ey87rY/BvOrjKT1vp1F0gQUuBvsS5JXkBkvdoijq3bu3Y3WpDxfLKSPvHww6KY
cTjl/dexijpVRtav4BfgcyJWUIn7MJ/34c7Vsh4/f75Yips5YFfn1/YR3h6fqJxs
qcF9Kt0DEY+/oOfbHjIy6mJghwK18/zfCSffGcIVXId5hlbQ97qOloxVayz4syh8
Wr4slaVHcli3VRaTxS8smjSmRx+7OOvNqxAuJ/4SJ8Imlg1dTgvUeiJzBIy/OOt8
gv7ERnrHaNokDvIdJnW4NPNgZopqDR5fIPljnA/SQkE0/h0vm/IJMTWhH90+ADTA
TdlgJn6YDHe2u693rOTNpVTUxvcP12Bt8yek4YLlhDFItxS1doHN7R4gquMzA9nA
WDj1FCZaNBxbw0c+0wXbUkWHXpEO0ZUf4cPBvaKPd9Z/qUyjkxhhK9PPh35pCcES
HVKCka/fsKRJ6jXiRAgHrPF2Mw9/LsTFNu3l2FeNiXBslz+UiCgNi/RZiTIIy0aJ
bemgGgBW415Rir7GjCI6YVCBTPzksCikN6VuwaoWSVVNzmM53DujeUWFsl6lUvdp
dssCB8CnN65Rl40ekc97C65B/TW48fgCtt25ZrqYskh53iF9ZupelaE27KtZvJRO
hcmSf9/9hNIbRZ6+Px0fMPLgs/cS/fmhZbtZQKpGyrUTvB05mLsV73QVvONVIIL6
+HubxR/J9hiO3xUhjiEa+XCJxnnJXKQ6rx+xXBwwebUNoGj32Fs1vaeI6zwJuJ3L
HRvwC/e1+LwsRsj5yozrvKLfuqPT9oe8XRPgRagl3eHtfnsGfH4Bu8dNNn7qEC4Y
obxnTqaB1i8iTuqFeWrjcd889XlqsW9OZq8JJ8u/ZurRETCRg/h+d0ZFsZzDzE4z
RUUO9RPQLr+/8BzYNF7Jq8AsxxCpAMFz0HnydI0mm2q2Yf7urLJxEYzbzAX9cEPd
EfcFaNz44yV3wbINw1oyLEfxJ8gxyYJYymfAUF84Bo4acGGIjGdcfGQ+oCHGjQ9o
Twa+9PHACwLvwIIZGztctPoCM930qB2BDIIEMTe7xbNBlTTB4B37AsAeEhlj2+lC
Oj6R85ZGq3Sq/fCtQiFwqXasnjYha6uUM0dHEIY1zSVLIf/ZrZfBsuIAj6HANw8W
/rDXSc3xTyhvp3+pO28Nng7dtz+pf+X8rXTFMKZKX6rdL9fDTToozx72tt37cEGQ
Ws3AIGSVOcAtPaR6glztbbKDku9JBN3gH2PNRTCRc9vM94N0vmbg288h0ktL9vsu
6iwe91Ybyq94daV76+BXAjslpk6EaNZfrYqbHNhN5pt/RC33j1UX+cQ5Q9hLWo7q
AYWFNBraWG9xKEWL5LwIfRRRw8MKTgtUJmg3MY9yx7/YGXHRpZHVivma4pesJRvS
OtSJD1QW5bYD3WyNHGduErdHj5YG/SPzVlP2ifFvuNSUkcs4UNEb4UsDGiwEowia
31cuCwyTJZ4vNMbhsoh9IGcRVPVnTKAe4Pz3yw2HWZmNnDhxzzyzljCEMGijX0bd
R+h0L0GPUjbDd9zLs7uYcl5fFmymrxLtp3TWLlRSoyKy/dIKCpU+qLuw5xQDuPxj
svEMPCx63Di0HFevZEgxy27rkgWO1k3A+SNof+UpqTBdW1osITOv5LYh8yTv12iM
h95lncpXXgfWjqvQGVGIvKF0wz3GrjcqoEgVpMo6sBUdoyLeP9iyv2wBS3GpSusO
GuY/tiL0XestZ8unOlHhHITRi9bEOng5C1NPxUDK+gYXYOGtcRDFH9u5AqTIgRwu
a/2TR8ZrxH8xjQMDcUYlESOKlqbOumwmZjMoo2aNBJG57hlnxJssUBnWUGH6WSJz
xtbnWpM1iRBu9Or0EP4YWpiHM9hBF+MIrifM2AWYeYW9JkOd8Sw8dI158vwGB5q7
8zlegqUsZ5bjWP9owu5LdLHNWh3qUne8ak9AkojQHA4hl4KSg597ROhL+/Heu5SP
N7LnNX9iYADlKvYPbxKjHca9bNJmjCmR1PsSEBVjMnYsknOL/RegoxSYvn/Za1jW
0sTAVWGCppjzIFYXas1+EOZ56W4OOKx/cK0FnS+LXG/16C+eKdo1X8P275aH2mA0
SwZHZ6RWJvayC513XnTsTpiuAj6PE2U8fmfj8Om8qCq1Mn4L+C6CrpcykB28MY7P
1ImCZo2gi18RURFvRD4Am9dvIjbo3gLrI1iAPqw8O54/qfTXadxO0HolpqLKVTOQ
Dc0YqXRl6CGjMeuei6Y4mvvzF8AGPO2x7AdXfrKX5hir4/aGHTxumr6XzaWRzkB3
5oyMMudAm/vWsSCWKBNjGOVvMaZ3KpvbA3kC7yVZ6GHsjZNeFw6SYtesYpsL4Qbl
bg+acwx+Qtahgut5RveRAMTiQjzpBlqShk2VSne4hFEAjN8Rnv1/q2kBhod0NMOD
B6AyyR1RhQRz7Wi7hG5dg7mIHZhyz5QMWSyPXZ9igVX6mZXhpOWMXySHgEAvU7YQ
IstfjMEX8YUvrkDy9c/TqbtElljUuxLiMxWQckUCG4YVlFH1SqhwqDdHJWzyC4Oq
XAZsnptcdV50wp4wE7qdt017FyLi7ifuKBEStHFSL/64v2pTHRliwdGgelEUTfaZ
PZtZ3QsBBuFMyBHztWxLR3hJFCH/xnRhR3/5VraEtlBiHOI6xXrWAeYOFQsf7JZH
+AT4BSs4LiqGBcWSyaPSt+kY83W3NPHF9xNjAegE01GNwcB2bi2sHhFkNbcmN1gE
aaAc/Nqf822tVDyCpYElGks/x056n2IMkZ6j4RdTMLgdRk+sWbS+dKPyyHmgQjiv
j/f6s7VtNGGoig5azgHSJuvdmhP9BqYui25EJTcp/VGMIUegtI2fvvwPsxHJ7Tye
CbFDqiLQ7wOczOmHGDNiTXvHC/rrqqLemxjftW/EReHxAi6mhEdbSuCOrS9851h+
Z8QzxZXozKbjKtnz4AAeYmSQQeliwvMTS7jHz9iGqixAYcC8yqKh3AEa6FqVWdVK
PmcKmaAUvWqAcHCN45HjiypY2yDNg0fCDrWeS4Whem0K7mMlqZBSmxLvT+G3znhR
Lx1gxSovyAh8pEoWbpoSnw6K+s5K5i7gzZgqs8Ijk0wH8Z2LCmLdmcSmUVhylWPT
ewsDx2W52f0IZsUtHGxPjD1eNNY74WRbpTe9xUVh/KVlLWvwDP1DH6rezc2E7hyB
e/CyzBf04e+Fb6Q/dDqg8SBW87T/5Ly1/ISKwhPXpgC4kx3SJYbDjkO9K0Gl2uHK
QUb35l2WWvBajMd2PEsTU+jsMBLRErDoiZppWvXydO7UktQy0bHCsKIE6NVljQAf
jjAJ2QhQnZ+uD9Ocjs4pnRe18gp6vizxoN4C+XCWeMLCrrOQSjE3lv1FkpnNOWMP
xiGdl7DdAZIZQlZ2993xjgJnoeETBv7/1Ax7nZ5FhDciV9jdCMI3a56O5iVCmhyS
9e41T9Qe8ffGY2njNtw8mxHkll17u5/Kja7pXQ3a1ubyzm08lmSyS1osL0/7uTjU
j2oth6cNeCZdpFCsLueYIA28Kf9KP6D8IHVxNmSf0xpLBmqFdoYYOX132QdtcjTZ
5eaR9pDtQ5KnV7puJx9KafluoR3qVz2IJNDTJ97JP4PMy3qk0lUtHTEot3vh+gIa
hSVeV8fhKuohC5C9/8JM8HSkgKpObt7T9Fk1mVnTmyKzK/TGPOS3WkkhCWy3KZ0I
51m9ZS2TWel/9Ie/CLWBnQ918pCfUxn9g66Z220/ke8pdaVjCe76IL83yU5jJJuC
NSLUBvwKeBzQJdyvzvbeXZ11YxLb9LS3+6K/A0Ax2Y16exVbDGZ5lPpMCj+J1ItQ
Zas7Rfhpu6Emxx1g2eLyjJQ7Vmm2YEEHk4SNR2IyU6YLY+tvxI1jM2/m0p40LVmP
E1CH7+IcqHXw26ND85LG0zZ17pWKEhJ1yfmXPe30KQwJQSN+JKZupp+1yKZ/scOV
h5mxkQoZ5A6xsTF1RVhGq+F4h+xHa45zD9Qeek8V9AkuZ+nZ5ACU97m4hxBVg2Zp
E9ns4uebuOFlTM5Sb6fSbZxq2Y0vW8jIjKr0ucuHVkmc107066zcOIpJ+RIBKlPX
B4OthOsv3otZUmnSg+yFyJ7/uSrdKmY2CB4SnMbvHlm13G+3F05MFFHKG0SzpqZl
mN1TPSuKZ8u9QQ2sODpjcaSRuMqcfic5ucCPKP4yiS3qtJh6IWMe4RO2WgrPAq8a
FC3nTW1KwpfUcKIXh0Tc9a21RnsrhvEXLZtOqNRp56CuoUQ14gHh5jqJf5YNvC7i
wpKHgokNhRbIPDUJgBlYVNuaINzPEovHuPaI7rGX4U/McfRnDHZog284HU3/0VjA
l8WpJChUNIzNkDCKX4hLi4OJNGtObDcuw5KYpoGW9oZ2sNwAi8zOhgFXn+pv0DuP
h9uZpJtSCJC/RMmZAbncuHwBJqz3SRrvKn0Sctbpy7UgQwCbQvHXE/ClXaE04daD
Y7rV9kpxYz9kakP+W/SLiWtPAiCC4Zi8wTwXMsjnU+8+DO4sRhj4lgtOvJe9vES6
MCk+vJYHYWU1Un5mjK+ThSWuyHwUDhol5LJ/V27BwaPYa0KBzZx62jNxJ7jPXVKj
COsRgi13kIkps88VpmuWicuJF9tqct+QSVorqYwSa66D0YSbyhNsgiFa7LNTjaK0
ETsKV/fVd6R4Bzm5XZVyZBmstykuf7DGfdVY1XlN65zmKUYPrivIkbZtBR45fcpX
bm5VtDdljam3MpCJKtngJ+2jdEdE/EclEnfwKojuovO1ph6QDIinY4WueYbRzz3M
g67rUpIU48KE0Crl8lJRYmOKzMWagJ37Cq5OXpVOXmiWSCTP4MCjhLyFuxnQx5ud
FR+5ixIxAJUkTQD5YQOux0O+k989h+QCPuHWhpPIn6vA6P5RmQQaoPy62UXxPnQG
k6+niULqE8m/bpWVKCgGG7t6+wfbDWvAUVul+aWi8Ba6Y1dZFCzo003r4ZPE9N2H
9wjuMJqbS/5qMTNFCKwOf08d7Z6Pt8PTbMxBWzOiTIx+0DL/HajguHfT7QM3ftQe
IOiekr7NO7HyIeO5jIgqSuV8mYmFk4sFx+aDE9wg8XlAiiE2PIi9TzbwXppD8sf2
2RaoEROcNrJf5VENu7a2ADDNLYDn1TnKoTlabB39QzV7F/MYt9px2FvrzFVhSqJN
sf23YdkWhyAV1P2jlXMAZsL6JE+qUt/FoAyrHdUuIsWOGvtjjncwrsiax0UmGlQ1
F2rDjHb69Sao4RlKopmzofYrMfGqmF8dHygzohNUh1XoH0hqPauW5UbSoYC7+6yz
zGiV9McVgOdoR/lXTq9IRBKhr6ttdpgoBXbrcW9Mgpp6YsI9LZLQoLuV6EdB8ggo
g/rbL9k4ecfwV3PgRUgMh6OArKyylbxH66dI63PYVni7SgXVok4HNLEElY7z1gJh
9uhDoYrxrOruMbzrfB8ptoApjvyvnBmxD2yu3egl0CaYQ+T2C5eX5eJQJa6GOMQO
D0dWJQWTzHtQeibTWGDaT1m4D9jgZuMZngr9MmjeyTLMVteuR+ffYb8ZmTcmUWO0
`pragma protect end_protected
