// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 13:57:49 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
rGooeUqJww6dggldiq/NlWDs64h+Xhx051dT7Q4LJ0glm/g3zmImfk/C1C/deA2l
Vfk7rtQNsF7Ga4D4IfsWmOaFM6C4QEX69v/r64hCNOxR7NEVEwGej80ZZU16UgQH
L3x9w+2v47aGsxVQLOUtMEOHkTV70Xk14ozR0FGkIWw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 13344)
5f9iRA/NExNCaISoLrl7b57+IsylgdDBifHXipblZviGaYcVtFCJloZHxw6vGzmX
w+HuoZZN+YHm6DV7fJDClEqQ0DRqkbAy0bpGtsvLOGTeOHIHsXwxZ/UnIDBEBE67
35i1sOq7T+Y99HN+oTUotCWGYdReYY/JWUzsn5leZ7uGURAuHayKe/bcDfv5EMmR
ktYArxe7ln1p02cLcN2uMy3x49QXlsAlGwh7lTu3bwG38chxtzsO95XeR9pGBd3D
/aihf2RXrgIotf13xR5IyxU3JzyYu5Xy633SkQWNWauLNSSz4SZOsEPJzMYL1rca
ZKmrJ86OqvqlG0Lt02cCaUY2tlV8AEz3KnbH8TDkHBnZ7Ss+AY/wQZiRi6VXhghF
ykY3K8Sulo3Ie7qt0hU2Ays87X7s4L4a3ZG/BdF6k9k9l9Mz8bkQsMl6/cWvzaYA
IOCn5rmYDh3elL9TZav3rbzwtIXvfMwNzlkpXVIhMOb/3QJybJFL71joO4mFbCA4
RupooI+v7vcslJKEfirV0ecGpck0yaueYp4GHr0Y3z4dUNETt4prwIDkTKPfSLTH
Yy3yyqYy4N2oesWNWepp0pt72iDdtfnVC46mjtgoooeM97y3e4Of1BrlP4Ugc3Iq
79mW52xYrh934yX8Ss7wX73Tv7vRITnSuv0X9UWC8W7paozqvxmIEMoRwcQ0x/kS
pN7IRstzkIrX3kureEIYMDx+8MYyAv+YSdrpfzbms2PxTSm8LXPykyPkBHzJDJI9
GksT8HpaH5vq0RE6bEhgIg08WFwIzk/ke7ECg94Ro3lc4vV0h2mFA8qMHXFfHLXA
32v8ES67TQ7oW+2qUQF6HBnI2GAbs1ZZUDz2909CeHEwkf3PpbkVMu6t01XBUe7y
zLQEJRBkgXrRF3yXi5KUo5CwlcvCmBCgCPxbLW7wnlljOxVoSDBNYbtLnOKpNt6Z
5XNt5cC2vWYXImOoCeD2A6DgJRemQkUyrjEapZdVSHotKn5Nv373HQteva3VoPPg
z/XMmMkWr6Xc0hv8QD+c5xfe5qZO0NSdOYwlZCCBVBXtnqRp8vIr0d0A9gkzsGfE
WlieRH5aQT2Oy2pZtP4//CYHteTylRNI0DUOzZuV2NAShZEsSEtsumXFC9Wu8ErV
C4SExNz0PdgcMOX8Re/AaRbm41hYvSvRJW3z/YxVc9kRK6tg7WCH3cvEo/BzuX/e
8HMHnlWPxtYBSbX2DWbE26bxF2rU0u4ijLfw7kaetuc6O6k3RLqnmy6iwnhPftXC
lZmr7jQS41Jf3j0UYr3/yBDgEL2DPjNxfkUSwRPd5YiQml0j133IBJsO4/3xG5VA
Kl3HhXPi45Aw9RIWdTS56kWDjSfiRN/8KTycUfbRzfVffRM8hOKkWOUi6PyBEOzQ
/eoKLVXl3nDXC482g7rlYJs/aqIsRygoo96aqY3NuR6Jtw0ytNTSNSxVMghPJAGY
P6ZQK+bDC+HCLeyhHkbk3KzPx1GQzv5RKP/ttSlZAwWdKn4L518rySYbRMxZRkWS
bFt1CzyxBrospBhdnOr+pcR0QArFCM8GEKD2fCNl1u54eZa5E2GIlRIm+a78vown
rU4tYdZLL/6/kE5shXUN+gKdpaII+aEGUDn+xbzUdT7MK7YekPZ/lfzSdb8D2lr9
bEb+RRC0vrVB1RPAYEgA/pRToKtK8LMTVVvk5E4ubtv44dJS6v236o3+MApMFlk+
kuhIaKZ3fdARYlrD6+ThuZHG16vV4dqZLRGB9M9eXV63eZNCzxQIeSzwyihUDL2p
DLaUD0YAL3SAVER0C15savg/VXaxaFG/Lz+Q3jM/OgBGkOGAjjehRjrEuwkmbGVD
5tC06HxerqHZ1wNVjaOBKwfjvEjRGZYJJM+FKknxRIjmRXB4kz1QlB8xpFgCqdiS
YJw1+ISoQw5MNwDXbKmODp5bEVoYw5TtMchECj/TvapNKNQTFQBW+NWsQqrXUkWB
lKid3xrtWGYMh8J6UoRjRoWxv1W+2R4gqi1Os6Vn9vIF73+KC4FIwCPs2m0smZ9g
Ekk0oHa4szp7h5gZW18nBWLT2Z1PDtJnEf0r+YjmWHynvPvJ3bCwzLmHDy+9snyO
B2+QplWhJg6HBUSLOHbrrJz1f3vv1kZEwsPTpuELgRw/frqcLiQBqCfGa0FvF7dm
1Aw/RFiJGK63fFnd4kkEnKmCwqmS/NqUZqF3LOxpYB8GcnkOHJn3J7lncomNt9H6
Dd/xKcsC0NoCeq+8FSQ5yWypoqkFZjRkM8BI4+QBaz0623VEJzha6FOlrTXCWHd4
Kg8dyO0CUnf4wROyzCYB2IwX3fWCo9LElm9qGbEe0Fh6tgyH3IOpx7jRkZqvGUTW
h7+G7pOuWIQIg9KVXUwHl+M+8lZNo29yQfQsXuGi+CiFnQi4pwgBeSiFrbxdU1Gc
mKe7y8jHqtAuf2s9VnleeEzsOd9JDr+Sncvn0L4YZnth0UDnQDVg8pnsNC6CSYK9
YnSf1Z0H8FOvHPI5Okca8rhwYURVS+wTcXER+KEnijbwhFrgms/6RjZzpG8yofE6
Li3gVneDfHxv1sf83Dcy3wVsXVRC9ZGZsgovsltHWBblupRLzUps49jVS+SrnUvQ
ohYLL8aMhLNfynf658fEk21H4OxNHEllesG/xei5d3QqEGC8JWrXXD2rXzItq7B6
XgCmzvXDMYmcntuC7YkiH83PObszGCUvDpOu2o1hbbAmojcnM6Lyi+IK5r9Lm/Sp
00vOSbH6AQQeak3CiComVBl/hsfWwIh/22FGMwgXnIT6K4XwWStDa+hgCQEFohlR
GAKdQO3qiGncoGBxEGu+5O3kRtMz5eA1xsFoFWttT/4NsevAx/D/CyX0s/ldx/yR
GyOPF5X/qVP4ksnD/D74wVlD8d/LAhXpumQ5H6/VLxLhQprrJEUk4D0PF5NnBUb3
BPYlzquPTQ5HhzmSyqtwYv10vBSPAjyIDrzziV2GaqsCkIFxK0Q+zQhFR5welLan
Mf2wzs0QEQzD/u1SugnpK+2Pig5wOEo9sYgNvG4B7qVaYOmcL/T8ObP7JpkdB0Vy
b2OHEQ0Ep/FS+WALq0rCsHZpb0OtKniVWvjqBl2Z7w30OyrhjJPopWI1LvCePl47
+a860iX4GMmNL/Q6h277fH01I+Kdn3wQU+vg6atIXbeK5PqaUvX402oqnHXN5SfV
SrVsTFJU7sRlBnZ6xQjWMHj603Vq6jpyy0W+RZjFR2Izg3oJP4ASqly40Vss6Grz
xziGKpvfAgtSzOIMMnAiY7vIxJuw6Q0i7Bn9Ty6SoKxx5b79SQT+94IPbPI1HujK
juUc0F3uTTmheSV/tTpcStaEulwrfjtqIXTE5i1u2o2+sO7a0/IVTVpgbVtZZ2xF
Y33DjCDrVV9zjVzSbI+4b8YL21481K44VYy7P4w1O0bH/vJKmmbn+lJwLsyBVbMj
Xel/EoPetq84JNFcg1U9izG5AsB310KCLOM6j54zdzFF+PsEDFAE6D9UJrzJgzU8
AbSK2zOhBxSk73erXjCajHIv8BC+Dc0YAef/ng9n6GmSCN5/4q5dWbaYA1zlWSM8
FYnVh5o8Xt0rdz7oJCfA9n950Wl2bvetbPLZVgLjVe+ktz8J9pSXB2o4NBIMD4Ey
2vfxH7aUoVKinKXFSrzxedoAAEWjR1n8B0ky3AXeBKiHztP6J3w1ObTYBDR7nl1K
iOAFDV1ObTxZO86qI9ezmEh2XXQ6H5TH2vp/ZxF4G35aqctmMyGkpFiHyOeZpdKp
lebPFqrO25sdGcx5JRuzy2A9r81T+Suh6Zb3hPc/X38Y+brS1nP+bPuIw8p97y80
XuLEn/RTkhvNd6nWFMsmR4dz6cVk2MRn5q5Dz/vVGX1ZhG1juH3/nc6JrUyKwsjs
OdQZuB0+/bGo+KF+TstQzqsoU5/4Te//2U3QBnKs4vVQsDu7hHReo1cGZeUxJWpE
XpOkYdcwLYDr8UWlnGVTUiPSXSPWHLdFzM+sl0rRmbqeu3KRPyaKhh1O2sZHv9wJ
s+4GHSRqfX05doHChGFInPYZ7wNKMKVmZ7i3oN1PSa6eVYhFEMmX4C8zoIVq56h7
rneDisycq2ZA0Ao6Oh5FFmUiRMdppr6Q6fx+vxA4R4sFbvLTSK+nvybzdkK+jxva
TB0D9GPM9rx6OtHCnSKHZnyiqtzNDuBThHyrDvHt1+p1LStRJx7JMMWem5OQL7//
pCf2hKp7b1y9+7iMoiGrGiS3iI4GJSkZ3DoWqYr/zyfmaYWCMgJ/OXd6Sv1Zbphd
yY8E30bYyGnc9U35KIcHvptfbdq0WLMHm/CTLYxQQUIPIyD3lEyf1kWafvjWwkvm
Eb2ojbicD8mo436dFsKe/XnM2OC2oX1y+76CD9/3WLwE2OXctLvGneA87CDPt5w2
AtXCpYCZ5t+iKSiw6O7mySQC1OFQap1FIv85mVxo/F+E/Mk2/4ZNyN+vH4R9EjHW
yTDD9SH/FtHhRufQxL7ELl7hbfYnUDySBz2fwSZuWkDwdtEy1+F+cDTMSMBZL7PL
EYHye8FBv7BjSi0dpI+qwP41l+CgT07Axr0+BFS927IRJCB1lDeBrnO/0xaLdMzm
fQF2qnMBSucSlFdf0eZiFvLvp+xe8ilKRB3XwqO7w5a99OTTJu5tjhgS2voOQXYw
WZbOW7zeU5xD7r5pe9L/Hzm/RtAV3fiVyLXtbPJBXyM01lQz5W3BxS3+b3g7Fchx
lDbj3nvaGEw7fi7hs+9yMiU4HXaKa0q/lRGy0sJx6o7auP5oIaoStiisCIFXw2OF
a/jjrnmbFOcpgL+fqL+4U3RGfASSKfOc3nHjoAU54naxxiIXkO9+EzX75Ofij33g
YfQ8ZRMV/GnQ3yVj6p9+wZ+1dEF/OuyQpWhkivckLdsB2t4yvc2R4Y0RbhS/bKc5
Q89kIwR79c2gTRU1h/fmyqfWdl7ExTxX8E3sHGSmX5jsHDVs60y5E39Ed5xBrPyD
yqC4HhOQHUd2zQ2iF8Q4NsDPVePNpBOth8Xt3eZyxEP0hxksORo130DBsc7JVSR8
ODm5g5UTPcUP52t1jPLS9PestiZ65qYnhe1tQjNlk4vvcTzXDm1INNeZ6qO8dVzj
CDDXfCepf03v0bez1DSPbwtMyiIRZZZ52pFIJvRjk6gDU+dGgvGXg+uJ6l5q5gBQ
fxzSkio/QI9WRRPD/IAVHucCOp8uB96qsmZUXT/MAW13as7TS35pjcjXX1j6Dp2C
BD4kIsX7z+7+q6i3kvy7ALD0CrZOHzGTG4RVtE/sxy4KVnjCAZtV1yYNgQgBozhm
YYGNAQJZHfhCO3GQMrGb0i+Qamiswgb604jyD2YziNbMWnrwuXEnuGoUb5aRoNYO
3hiprIk6VDYNZK4lRiQD2LAznpXjpMFYUjxhJTQq6TSoma3DJcHQAYX7D0wCYVXe
Fs4TDCCOmNv+zr9AFhBW4EG/eDoTjoTJqtg8MyywdmEmqo9cN1iaNddk1m7WayJa
BFHhx8L65CCace68X9EoEhXxdM4GKTZ1NxJDB+oix/yvyNVLZvyLCChmcZdV6rY8
x7imiI8aJCtud0R3SbgQCc5I/enyI9l0qPxIewl0Fhgbx9buPs/4fbHSLtI6QpAE
lQlnJd8MsAGcfQTulykDIfk7gnUQtExtQxVKjnL2x7hRbhySBTYDcE031dD2hlsg
HBzejEmehkedmOaa517EtVaEugaD1o5TQcUxI1BPC9FEtzYadw9of4ou/fFgLLkA
xtPntxUt1gRvwtf6jclG3Hz4oqFQ6Z6V8QI2zdjcr6/Tqz1mD9SPzLjDeuMfpxw+
+kvxC/NgLcbcLm9zO0MOgpRsGhQ58ge8cMaJMfhC/ZoVT1kdQTXbT2yC0axcz9J2
viJ8ZUe5+gZ/EpXM/TV/NA5Yt1cf3XMHyz3iS5fZeCmOKPHm+h6gYC2U/Km03Ppk
mSDwHMAxPSvs0bkMwdAi3L3jtdEci4ErZhkAl696Rgm2XN1sFB9arwBpeacob93O
0p5QBzgPZzlF33rPy/ODcdNmR+NN8IHouEm0p+6x+SUEdCQ4j83KjYr9hH7GSpAZ
xyqr2N4BaMYHoVGjRW1GPIefra22e1kUSFkRjMuwygBWCBekjaUPQ9YQk7EOXvyo
sdAhFISk1IuNg04ujdF0spRx5Bsh+ivKa7Zmf9qowz1jsKmYd4i3ZOt84U+1Ieco
gcuvEpVr+sW96s/ATx7ibdTT5I2Yut/oB1m31lJXIwNkSu9dKdKyiTLdQzkNd6Yx
jfGyQtEwZq8v2atNl1DcWGE6vv2yx/sqDlFvbin6zY0xg7npbXQADHp91AxJPnvy
wy681sFogTI3haU+ERiO8eycaWIoklW+3SopysHvBG3TCwZF05lBZmkky2eNsekg
54SV6et8nd0skms5cu2XLfRvjwK410dp9slApLqNV9/j/X0XkwK5ivKig1oGJc2F
VZtQdJy/y7mG15eaGTbmqVd/0V7cybWLrb9z50r+4lqFAH7JskK/sXY5g7WkRh6A
ZMrQEfZiDj67Z1QFGVLsB4pt1DG7Zurx07MeL3KAsStt14nYTIkoHpxC/Q2VMjCW
vCHKMrStzkzGquIDZXeRl2IFkMDWdbFiW5T8kDbecf+E0iClQ6KESQX9W4puvYgu
jWz0jrbfJdvNDN4WS2t5DiCB2OPPsOVbvz/Da4lxEUPgdxkACZyiRiNhd+tNnqKr
0bZlPWKV1uy7OMRuvIwTkbRGCzFoYwl/s/Ry+FIP3vG1F57iI8+5ZhVjn/djDFR/
KltNgLyW7KILV4m+73Kv/eQNvItZjna9TBKnga5+kND3a8Ymw6uojLSWVtbwTD0b
zE9U+7LiKxT58wCQzJ8bNlJYwVwMnmm4EjtIB+QYzZKWxHDApYl3p6bT2EcctGXq
WPRcgck0eigCA6xMthSs/i9xZXCE9uepsn+AolLAmA91zQXrU7Qm72AvZ+NuUoWB
O1LbwbLM6h1afYAFmUsNOMBisAlZKtSmmQWfalCJcxyRooWtAmoIJkB0ygu3XSy/
I+o4qLwoAPXs/c+xFVWMM16FoUauSnu07Eyx+LKPxTtA9lYs3DM2eU5o5+rTJoGq
8CGmurMHR+biv189rOO+KGcg59QPSLW1fH1bnwsoPLav5pHF/dH8DUi1dND3Yor7
3vThm5oCKbVFDgRV11kgoRhPEh3bt9kvVoj0qKaq2nsu7c0DIHcsfs9OV308KktN
nkURwu6E+MX8dK6sVaXWj6jvnHBU8G/rPRHlzmPv7xyaOXt9EaQSneRtE8Yq5OmD
u0OEoV29/yG5Skrnaq/Fy8NponC2MBH25mbpyft3Nly8HoCFhekiIn01QA5RUEwn
laHcV571RVZOvmsPA9vAOk6iymyawavgY6O8jN47e6D000HEzByll+rCF73EE0RO
q8nwEmkJljor9LXMf1SzNpsbmINXkJ6ugs8HSK2hKwGsJLXSQ2P13L2Al+KCKSI5
8CDkxCkqxtjaJ3vwW6uMrOr/pVHxzX1pDJqhwW9NfxlhGQCs7ctUZJgWztDlDoRa
WLolkqoqMfSwH5bm0Vv+gC8jBA/AL/Iyt5nYTzMJ1gqCLy2bHNUixcaqEhDwxs7G
88fZBDMjKsarNsu9Nd7MS6hMpgIHt7/AwkeYEvv7W2HPUEFzChbUNuJ6K2ZB77Rg
LRGFkDHILgUigVfStCDRjB/xkQpO0agsq0tD09q2OreCNt1e1INnrCkuWC0ra9Dz
uWI+R86Me8ZUWx+sBNRNtDGti9p/SQ0LiMoomSJkOGuh+MjZTKthTgHH7l2T3Z8Q
VXMSAOBdbeNM3LOplCrzt5fR0WLw6+5qsXdlIscmgy3kl5FcUR5wrtfF8wq5gwfM
j9goOxy4L/ohwxSda9fjxutOHcaX9ux/ExlEBnOay5FC/E5xeXyGYzIakfYM3z3u
+ahv4afucReZ34s3qnY/D0uX5QHjLmZLMseVdTuSU3by8AXhBOaJoqGXn114yGLv
xZuu/pbNy58X6jIp/JdoLm02RDKl+D+RObI2s1XQILZOSCLZvrcpJkpTqTjmCmPv
kx0Acq0zpvzEuGR0nMx+675DfO0UGoiuABH4fgBe73y3rxhY5oBbrJkLmdCh9XPU
ehie+70WDRaW3FID7cDSR7ouG0Z+NOnE5y8i2/5lxtMzRL2TAYyKxf4fKTD5N4l2
52HCJNxl2iRUtS1PfLY9GtLkqrrVoEsUldUbrJ8MM+WL1peH1axZC1h1ATkmSUwH
QJTaVyJeCOCbTEMT+sV9vjx9sumCPx20SZ+TC42f7E4HfxCDK6gNJdsQa8Giwh1d
YqX2QVC/xjcMwv+m0ro+xRzsrcvqxVGoq0j+K/QKW3WSDGgyxKnm/0YLFmQhhYNQ
4MG3zoCBeSnaG6CeucJ/yQm2un25OA28uf8DVDatG2cDg7kc6IIJT8As9STqG/As
vtujFwX4moY44HYJhuQYSQfrQUxpbyuYbliGrkDt+lofMn8A3C//eqI7m4sA0PlT
T6/nQFstdpBghrCnUgq82iMJYpmbJyv3utHniB2FfbOF+lLtx2eXYi8QfpoognQQ
8f1PSZWiyxmZmWVzGN/yKW7JHwZkvyvYzz8H0wutvuao220cEq0LwAR9Xvc3pB8r
jDj4Rtkid8YiHn5bPFXBrOA6zF6QM6Njmgkmxr2AHLu9jDA5jZxezfS8et9+xck3
gDHF3QogxQW03GR9/W3jbX76oXHtTCrLlYBfuAFr0AoKoJPA2gY22gpRAhg4l4ON
vCuf8ZK9KtLSDBAM0GD7+EuulUaahqM1G2NYeseX1/3I9rN5E6pVO/RoOXE99QUZ
P8uwbr6F2rmR3cUq1R715gNgxQVxobviAXwnlLR9Wy/sT6eNh/2oYLa86Tagzkcw
jHiBnc7AIWnfOtpCkwtNu68PE0XQ/5mMjzPTpWk37rhVAn+uIv6tmnSMI/vYhAYw
V2I/QDa+6CWg/XhY6j8aULOyLjNUBtdoGGfzCWdYf5DZAr5cWUNgh/QuSrPTwkVp
RF4u8WJPuiBCfy0wJ2lACM5RNmCuRQd1vf6MZf7F+aCMHVnHGSEoyxwdMAb5T1tS
VUNRFTpLcU9ExDE8esp4LCm8YfpXAQPnBk7BCyPGNhn0q+EsIuCd/yiTEFffVPlX
63PtEblQe31Ptuo8JSBoY6/BMaCWDKTpicHxY5024/d0LZL//xh0pvyCA5X9cUHq
RZzsZjNKyfsdelXJtoMUMxol1sfhW+6BwS5LSjWf2XulIQDZFj0JW6Ck1EVlkZnx
dpgfvsx3BLB0eOiUukICi/CJqwm3kArUn+bOQx9kA8yAAeoPcgEUxP/6U3kzJMpv
5Abq/ddETQOdSgsO+JK16Avs1W04LfIyHkaCpXBB0aCgst7yNNILNpj4h7/R4Jry
wdHb5ZuAmnIXxPGoOzMJUh6fjkoOxuP6B18MeOl1JWhRG53+WB0EYxTyLr3C+LZS
6rm+/QzB2kxJKsAV+4QfvwXa/6O1i6VbH6yih6WAqvE1GA8k5+z+gsFIFGkxCRKr
XMlxJ8k2UkCL3rYpFKcrAlowk46/qfPDDOoL2XWf5bCKA5xdiqjvdjiUwS8SXso7
5pH8nLGxw2QnyYr8g+3x2EFupCguGGvFeaMXjzdmKB9I33v4iMsNRg4qM4/gIveK
inpHRvmZncSfp671sQqJlbqif9u6UtSx4cRV79S/pleAetiA+XtEWgtkkHX+j+/n
Z9HCbXzdD66u3gBHX6QDVHjIjydGR0ZW59q0ij9smaKw8PFjJ+LmHcc1UJIvDzwh
zTRFieNnOswZpxPMgceN8b030LjSY1bVs0KJaradFxmmx//DUduO18ZwvVzMs3fR
BJYkswvDMZywfGdVP1TvL24WA1eBUMM+W2rmHbktK0rCNB0DL5k7ASKkOhrWEWEC
aNn60TLNiaXtGk4/L0c4lUkKE313GZRc2wCX3vtLg02pEyiGiFVVLLO7ZHuTrdF6
GvkRdRU8tyeu6v/ZX0P6IVSghDrN2cHlKjB3FaTzMmLBE4qrCIJirESioqpTsgHI
UJ95KOAdwqR7qJHJzTX9e2D6S/SSf6qDxdhdmOoLoUStIiGMigW+rYlTQ+BV4opB
Sl9D9RPMzcvHJGBnKw7RWmOEhOCiN20y0tuZTpojNsNjXxbKGw31N5kjW6E0or6Z
eLL4i1cEO6Lc7WtQVnNX1nG9pwbsgrWiw2cPjt2VA9x5uZSFjPXs4j/HgjUbHmET
e5qxwz2DQXwo8UED8ZiCUZlCUIKDzp2ATmoI+GFkYEgkIqc9w4uX/f4peP5ut+mJ
jUyXBtE+/NGYNi3RGvXLje/TzLoMiXcZJ03bnPULQRvKTIIcFMcwmxHFxPJ82h1e
hJVIjJEZ/JO/ztLFBKSOrBypgcCbazP3oqQ32JdOKIfmBwY1JKTssVta0Z2NfKNG
VujGoEVdDkKkUwPfGS8jy0VoMYt2T8x81q9JfQg+LHoufFIclLDgGc2ecke+dt3w
Q504ozjEvaCBVGHliuwiGSY165OZLvc8XxbAibomc3eShWqbjuqY7GZ4Wkd9RPf1
PbMWp0ukbWgNcvAByAksSo4rLuiUt42ndaa1X80rVrNDf0MX3Pa4pTiEI0Wf1603
8H6Iz8OtaibuWGb0FPqof4f/rKT5KKCddcAgqVP6hG1vtIpIGCLmQlXaToj2VLcu
+uXLUNYyz5fXzwbwxxVSsk06cktnMYbICK+di14duYzEBUck5hS0lTcRZrXPHhwZ
2P7IDGr4vSyDRX6okbJ3xh5SUJZUunOgOMDjoa52x10sKe90+d8TgXlgsBVgMEA1
sPRV9oRPJJ/da5CtA6yJ81eq/SU/+wklDKZobwTrdU92lWQ5Fkg8LLVZ9I5T5bDS
AFAquMeKT6RwXY0Z1vUE6htvaCpBoPH23QVdINeRNZAitNCT6qvfZKNf2gTKfNuY
+7Qc28gQHoEBMxYeN2BEnB3dEjNq1+QR1KhK0+wR1ZiYIP2COARqlODwexBN/Edc
2BOAUdysOja1cRFgWcXGh7aGXqKb9LEdAEW6YkRIz6N8ROa1p/DHBnBoyamrDNBN
uKXGphsKo0Q8icIs8mHhK4DfTN+rAFNej7MveQdPzuixz0J6oLun8KBQVVDYDOQ1
pdc8orTrAjpQKz8Hp7Gb6qp4rpAqiu6R9fdMOzWk2prdZi476wbbUkk3DJSdvqCQ
NBGsdUUojkbf8cerML3rNUiuG2sN4GnP2i7zgfPk6cRlYeFEGqKff6i7dj9m9O0+
nUPXFl9qiV8KM2Cs5FkKFNISoUaSOkUzpG1Lj8kJ8xELspcKaGNf/sMKi/rI0SdL
/ddO6noLcncdahn1+SUyOr2oSv86UlD7ZsElNiP7LZbxSn78FUfsvRePaEKHAShc
/V2lvRzdqZbMgFxbD2CBX34ttk2/coIg0bp7cFVgO2rbZX4g0z8a6Wllv3zVg2W1
F3afvZKF6VMbkk5BbMCOBDoxQFt4S/9PJKPMP9o61FSfQcYanaUDkrjuEjJ0Ytgr
whF3ZCaRHVNkF/OFSBrz9GGOX2pFFU2NMzwYot7bdLLVbOAfOfHfe4GLzWe3ASg/
L1O/X2stz3cA9PN+ubGkjs27qm8/0dW1eT17k8wysiA7N2yA7eg7DnQrr6DGGFkA
veCDsSKnUcXvjkufxYTCVPDjjmsRjiFU+EcZ78x06zkNep1+ecAOc//18blisulx
Rh6P1BAv+cynaOCfl0ptgXTQF7qzdfL3eYFYKA0h9pDx3gFUlMFfefNnEdSjoJgE
V8FOWIi01T2MXnzDMcwhn2itFqhvFx6j8RIX1KZ0yliRT1tTDB6p3X3vphxl/VhK
lzEcg++xXh32ssxZqKF2LwTHkbFTeqfbMdR51eBzX0WlL/JXkLERn11AzHoVBdJe
K1rwaCOe0P0znaqFMVYlRP4ESifc6PRmu5oG/ZBIiSt2ZJkq1HBhlluR7//Ate/q
W4SSBlfpiy+06a0tpKvICgkLPW4uKxTg5Z4Ty9Rpaw1nVfXC2vxKtNvmr0mQTuMf
gyez6dta1HrNfV1jtjrG4k9PuOx2tFKN71hFRZsLUEJ1Rb2aTU2nzhgO9ubB030O
1KMTAf1aHaRuXTeEAsN7WTbZ3CGZBFk96yFBb+l8Pd3iIXOZb4Uu5t/yLRe9yIVl
zh+OlZftN0Oia3hZvdABO9QW3xQgvw+B64PVhpjrTPxKq3D4sVBKlaj3kxAVlxX7
9oeCWNX56+KJsM1cd6llqbwgWl/AC/vDQE00rLtXpmlNelAw6EFYfPIFnuqc0YZG
DTtPNxS2N35KtxJHw+lQh1jAPUequ5TyG5BKwUJpSS1Adcszua8Cs74VK7zvCuub
RqP+u3ojRnP1Bz+no0sMtBhR01tpdvMcfR6eIBge8qQZp2uV+H7MZSpi8F/wxcjK
ZK5Pu09LO2T8oRKrA+xxhT41fx4h5sigj5/gyKWwzVV6VsDb+Xo7ljXmYvqkBi+D
82Nmsyen81iZN5D+79V2RKotw5Ji/RAR7jvHFWjqYgxF3poAuA6yN3XURruwF9QR
rdb15yJP6hohOCPn9zYnkXmb69Vyi7mBin8Xy1+mpQBZGhW4/lfK6Bx8yl0IgVF6
HkGY9XdCYVLiHQKCkK+H5Q5gAth8sifvfYjBiA4H3+R1oA20bFLdzPsa19mjgnvt
b0Rz72AmV1SBkRXw0ZTqT1/yciAYLl0uwig9tCvQTwvF6pvVqZJjX7VXZq1CUfuQ
yvQflanNOLzbkyHS4CFTTYU4DsXvhzH5nBoFpxYH0syRGq0zlARQ3KyISsenCw9Z
wfXx2xhfH4liT2Fhvv4YSN9Q8YBBD+o3Zhutb3QxJ3zj3SMTpFnT+ulIA+J/apeB
uuINVxf+rE+mX7YsqEXKxyy3iYIuIf/3shEby2sz1PYIIa1W8Ce5674XbCICKpsl
AC8VVHb8PqfhMZiGwP9IgIBDOyr8Cm07X783PUr6pWWqkkq8FLJDn2sbjP87TnsO
tPOyW8K6+7DnpRnRLtelnk98tutTJsKx0FuOZgqICs4Z4+HfyN9Ah/2fCx8DbJ4b
qxmKHAdmHKxVqJnx8G6gwHLkIxlZPqkQo5iG0P1e3T0mF6ANS15IEMWpaPSHI9b9
vjHn5bLZKBjyeIrgWIphbok9JavGKrJcfsSZ60HdutrrCJwCoJB7ZIQcKUgrsl2H
6gCjrd3NDKIsTdNKo1LMIL5nUUa/z0mkX1c0x5316yYB2kVtARPcbwKGjNdAYFyt
hHmwG6rgy0S1HCvdW8qKvuSYr3Fc511D/LEC44G61GoJu6vPgTaBPPZK6uZNQqqU
/ds2i8nrUajfRvfpk8XfId+qH9xMLlYrsSPNrlWbkHf2Tr9vLz7xN6VaNDjjaR0E
5M1Ea3BAfkaaFl6eTxDHyf9Rzw9HE6Efns3E+6YbSGgNn9pflt4b0JReTU6ebvWr
9ILi+lonw7SDOLRkLbS507LqnZWC9jOMW8OuCrBYUuYZevdoXvKqMT8KDt9O+Kq6
Y7nwLge1i5KSMUfL3oPQyCiaiDZxxZOTPtb0j2H3iovFXKs+eu6kELo4FV7nzBFw
x2czH8Q7ItVVTBnRm3MQL8RuBmkq2VhEuw4m3eiarB1xu1suwh9hoBW5A0d1G/K/
no5chz8PSFi1+B40cT4k1jI0LJAf4kwNO3kZyDB64xxFMjPmFzKRJSgtMyr5bsXR
Rg5iWQ4fOSUi3f/2eo93dqBUJa/XuJtYF1Brs2x1P0BoayruaO1BJvIf/R3waDwl
F0tOWNxH8RCYEHh7JFIyEaelmHNBgRKX1PKp1OrdTjCJeQm/5XNwAhoXlODKqqIT
Zt9i/ptRO+xRrYwO49BBedAhK3sqxfBj6Bh7h2Svkav6BgQxW0KI6/ovBClkIgYk
ZPDb6IOjCynavdyq8JnjJeGYMGRq7HCs5KDqfFQ2d+9YzSmhJiZZadQS+z4G5Cyf
5xXs2ac8Mf7aQDgx14oOGdU2SHwbSUZyZ4den5q0IiuFUbfaU8sWPnFYgbP4Fs21
Xcq7hzGfiwuLCq0EbpkBqJq+goWCajdhdgUy64TvnN5p09jkKS5qJKCD1cLCBO9w
QOnlU6TS7PzLSMMLNBH8JddbcHpcttmGc7Wx5V+r8nz239X3oOq7Xy7CwpvENN9N
GVrfGo7IYVS+t7R1KHzdusK2+7xbTKXHhTWiUpaqG3Im9o6X8g16KIssmYqRWdJ8
5mWK42Sry9J9N4lB93OfOz03xAdpz6pKK3jHY5ORhiyQxZT0BF6TZ0i2Lk6IOMtJ
1RhePKeo6NElPRfebAiW87nHYO2LpezV95BQe79VBarg3+CSxz4wB7nnN/RjaeiG
qxIZ81nzF6X//rmL/eL2RaUfF2Ta9LDQq9Ch6ABLIV3onpMLHO68B7KFikKrJtgK
83pgOu687asZB8wpL6X05m4/mPGmXKqxBB810ivCKbUf1HfzSNSPz6r92/lz7ayN
uDTMO+oXM2F9DwLdiwc4n+jiOGHaGbPfHNzciw9a0oC5oqNlVqmOoWztDGU6Vanw
jU9n2BzYwDUR75ihktfoVeH+XtqsnM14wT+ViUG0jQQRshyluxpeMWxgTHNq8zq6
X1WyPVeE2EnUTdosEK8OPTCiJa7LRHXIxmtQP0tdK9K7tR9fY/Q2j5nXqneG/2Pd
RxYjw2a47iCmGh2L1HFc8riNQvLPOUEXSmzPVjqsEjBeYkXoLxBf09S3laaZ1xu3
0O4OdIwSHdNH7WoEiRwfDB1ZU0oC+7ukEBRRt+rktAwX4gYYem7nliUWkuG7DIF8
jrx6flIpE1CzxTHvCDwza98FzCPuSg9R8pYTjIKPD/Nj9dPg93QYLU+BkuSkH+Pw
WLiSBaajQp7dOuOM0MXPuqGkGxsjUqXqpfgA+pW2HOlo39GbdFrO6YmN+QujufwT
pK7R/0C+AsGk+d/7L86bLSQttIjDG3pq+TqV65YEHyjpqHm/JHaXUFsUonLarsQ4
aQSvv5kIRkLRP1gEsoIDtmOI9RphmxX85CLYTi4nafkhj1OA9p7GD2SbSsIFYEYB
mmWAzc7nWrL1u3kOkZ3n+LBceR+qOZQ+8Vl5U1W7LTKjKo23UIA58MEfomwp2S3g
HX+MJz9Kb3I2IBikxVKtDxlWmDr6WEkywe3euhsI54QGYT8TMAIG5kRNdAaPjueP
kq3WSjMfb2gTAdYbPLWPoJPtiOhxSX9uRvZ9O2WTnV8tE5uJETYwyW5jS6ewXweA
NzvuR2HIIO5saG+0aaNskJSl7lWe6BJ/fYNlzLGlVodoeVUF8ADpwXq8E6hawIoS
Fo49TQq/8CjPPhveUXL88mn2K1PKm1wW2NA2/7jDJvFKp0khV1W4dbzxmZa1YyEc
tFWZIpGEgjNu7G1p0UrptRwsNlnJFXE8e1/xIsUTL7jNE+AAxUJn1xyyXUYI9doo
mTZezTwKj8T082nhEHkBoeTss96wZb6f+r0ES3/txiVjYIMXoDOIuZWRhZCS0tMw
NA5NC+G5qiQDHnMDRC1/CMuPGmXHc7IDwxFzOb7mQUcrigh4WDJvTtZtxYllOxH9
BVTXq1xuoTXIZ3qaAvS3FfHbYNrbiZb4Q8Rmc7kjYkH3ZfJv2XHlxh7+0MNQ4VCr
QywoHcMXmiBoa30cWxYugCEgfnczsirV41FJQqanobQB1BxXADYytZhBYSN4M9jw
G2SLqoM07JlFLNstW5kSeZ8BVMB1tKQqYjEUFuFRxEphwQuWnwxdF1GY9Or+YG/K
wOVaRXRyY6uLmLzq1aChfo6juP177zEZbyucVEm2oCHCSdFtsJYFcSUfGCtZK+2F
uF3niU5rukregbC9YY1lrQYL1KMn3D+m1UiJvruTViimk2VmFAmUw1yMmeoUclrZ
ttYC3SzkjH1FSsooWMqPZcFcPmzmKTzb/iJ2ckhUPWLKkg2j72Z4SkR9c5Cxpv29
n8U21GMSjWKdTr4hQSyC1IRNxe6YdgxGjPEAlX9B9ocn1b1BgvAH3xLGBwfrdFY3
eJ50F/7f7lteuW6f73cfvSq91WaWVNOYzY3mltz+uPMk/k4+AB7w/B51cQhFgTFp
w+m1dJffGGIg86ZeGMM+9bB+Ff6er83SFa7wj/QZo1twQVrpiP+QJgF4mCUMkbbx
s1Y3IZBtrcr1gIj2rRRo1cn5kWaYi8C3YFEKKatQ7ccKCxl9FR/jY8Dn7NGfo7EO
1giNqSI4L56IZZfYuY8sadIvMwkmBlN1aN4W837ydMlIB/3TcQPUh+6UOX81TLNv
Cyq4rqCBm/Ernb2ULR4EZ75BWhUFH1oTk64kQF86U48ztJyVHZRc8amGRzuG2T/D
j2hmwxYL7p+fQI3gjosQo2aelqp9xN8COrpAbYTwQ5sInGjhGNVyX6sY8fs4gwa0
xmitj7kx3pmantxqV7lKm5h7vcaBj1c2oRUsitlZyaQVz/Wp4cb37ae/hkB5sB2Y
yKnjgZ72wwLfDr7uZ8qkNZnToSoVUwtHn3h+RO+yLElWaYL8GNSq/bFy/tKn4FKf
LFsTubQyWW5remmbpCEmJw1qxCCMFb7jFOKUPuVvyVnl2+ZcQd5sl7xy+em+maUq
OMnmmDq3XrBZItSdsQrk/DDR0waxKA5OOUGnY1P60eqNDwVdji5xilcW5CXHQBGa
krrNTK5YcmV2WEhLfPTSN8pnAYqhQFSHUB/b2NQ1I02F2tkMteFS5V8WGA/SXTT9
AVM5bgvUshyIrUDjr/x7ZWcqESjTqw1B+yVWrolg7C/xrrTphnelONmzpOWQVodU
4RHw3657LGATTGvm106eoXWddxPHvZ0pQpGW4FUIUQZBm418QQmnGs/qXNpeKsop
mZcgcNkmOkN7aVHY4r+Qsrj/7EJVkYYYKgkbXXVTICAGYDWv6kMZOE9seOIcF/HG
3ETuwncmAEFi+FlbOZ9+HaHsRFPglahr5rexzGWDPCaDvGoJZiXyVQz7CkcZtpNj
w0lVZs7Dp6YGKCmguZTbKC5aeOY6M56Phzy5GCEGEQyhw0LrImRG5BUjHR9dADp0
wtKW2Vs+8pUhWgakt94yPYlvcjegBBMktePZgeet+7ozNvlMQyO9n05M55Z9b+U4
r3V/7SrTl4f36VFHlYcg0Xltv1bwZ9SI9ri7EBDE8sZKdDKPwJbP8lBi4+aSfyL2
xzNaQT1scIAjTK3ER1rw/xumi9MFfhKK7Fx5EsL7lw/IoGBy6jmCwD8UpNIfzC/Y
gOXBxJlSAC2ie+PTJh1X8gObxVHGVQNluMeODPVB9R7ehtkP0e+R3ZdZ44OP8bu6
dkZvShwb8Rpc5zkywCt1DlRpSEzC1l4DeFiLZNF+OFP8t2JqpH8uNnik1HLaMDoJ
G1Weft3TV/u0ApBKrAZy5QwGZAaYrTwAJEFrij/1myKlfuYFq2bi4Hkh0Fhom1bW
eAb2dZZXqyeny2u4vRbvUoWiRunrM4UVDxdZbwVpDmGd7mZfljr8aKQoxyPwaFZZ
RlFZYHyJw9NMSaWIC8BLs7s9sqmYxkjJFeTlQPuUyZ1sIZSN9Yzq5rwIaMB7QU+d
nc3l+oJNN4F06gqrY72tEI8QdCD7vJWVo70qNoSJZIRRGH0h+xIOBqnb7BJ2N4j/
7+8B9MYq77tWdzi+GvLvbYmuFaFE51AulI1P/6UiF0CLEcX3hcyLnflVmZRpQKkM
oJqugZrC1VzCcHYQc49CHyLA5bL+tWPuQlzT3F+WKFc5JDXfiAxHJXgIarjZUHfo
3HyuDlft1RGurfnspJcCcwgwg8n721iXdp0dOX09jyXex/4Z2J6iLIyijiOnHpeD
`pragma protect end_protected
