// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 14:01:25 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
OQlyRgGuDDVpii239+icGryLtFRBa4X/Mm6iyCuAMUrq2zIOpRc+3kVIBXpdU4/8
9ZNwJpwVk0idgrRDcAy/GCHLyHewa58mceCYxSMg7ox+D/ow9aieY7hXp1Ajc292
V67bEeaxTGFdWP5Vz4z0j3o45tSWOBSEU65W02w2Pn4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 21616)
NxnBon2b29bf0UqsQorgrs1tYf7aysTLzyvSn5E4+ThSJxT5VjFZqujdFfBOSAFm
mRDffTWZ+ARqdbEn8lSTxLTkWdkOy532L4bYPLwLiBMJrAg0NqxbnDu5UlZdOPRK
2FMboY69GR5oEHvgNHgN20W+acvHHr2BoAHNXkCRwam4ZnPASBVqWcEyUb2FdnJT
6JBDJ9X8J20uVhKZjc4NPZBd/E/zJ/a8UJuYAbnTmUOvMGA8o5XD1tsNz+6BgXl5
v+ATkTUHB/yq//zLxffIH+hubp05rVaA+t27CRXeetFkxSHY3zdWqsvtQryoeUUU
3AvAbHLbdNTb5t5NRIyK0x553Dro5tNqR22aHQU1zSeSdxyoZFPU/xnRs5fHkQaT
DXuzcNgC3M38pxqQpo9r2hpmRT1+UG1F00Qtiv1+b2UmX2yCUVvTf+afZ/JikVQN
EyE6uEXWYRha10uqS3yKUz/rBG5rKxAClImqAxVa+SFk85gx41dfQZCXN365pT6q
Wis20L43skpnw8YdJBOlCTbNYjS57ZwWBhwEEqmkwfbYNaB1c/2xuocHYLBNrHQd
w7HXaRETbyEqR2eG/fcQhNyg4msK4z6RtipfyrI7WKEXXfanXJApxpOsxp+Qic9C
Fw/ntbepnlmwzIa8T+737ND/mZ5DrQ/q3oGLC9jw6WclAprWEMJMPVyWLvybEDxQ
eWQCwD0hn38v/qmmwgkeIOvGOhN9cgYuZ1U8ptBcV2s+SH+qjbaPgQG7EkeeHvyB
AWlprP5LpNlCPLSOHtq33mLGJ1cKF3t2T+jI3aBImbMOTuJqx257yKbOBdXQukf9
lJ3V1d+ew3L9XX9o/xcTFRb0zOkFGEFf9tWm4cYdQjQP39QvYJL2GZSm/kYBKSQr
kVL0ma+ycbihhizloEAerHQCKsOEpeFAh2U1BR+cn2C31g5aKMSgd0+6Z+GuShnT
5thsJVsAB8pU66BYMWwrruPLGNwwe1aVtUyBT47f3Qi2gEZOr0hhSGw5XYwd3rKZ
Q25nSXXadTxMlIKBJzanb77HI4Jw/+j4gpN3dCGSGVIhHamoeZfz58kWlgIHuH2Q
L1oEZWwioctMnk4yH5nQ1LyWNeRqBv1MsCh3Sx0OkI8Db/xkNCQb2qIwuWYfcfxp
xYezOcC1RP5ievyGpW0OfSRKDukl8giYeFR8FA61MFEjhad+2tK2c01gRZniXh30
oDg/6tNTKB5RbSw/kR3cpZXjBGOdeoLNW/gNGU8Kib+kr2nffIuGc6zppoXqTc32
baLJm0imJJQMwwpRQvGKHxo7mffxXPxnIw4OhfC59UDonOoWGxuPEqZE65kGpUKG
ONL5i112Dq6GADXtTZBGJ3hrbWAjZ8QtSdLeqYD6Smp2gfWWIIjrzjwR8LcNsVI1
2kCvLAqBnqgKQ3VMkNfqFn/8LDxadktrEhhZ1WIShJ6bzhnVrFy+v1dMTEO78+dX
a/36seddUjEswVxNyoPEuuYkDM6J+ayJPUuyN7uPi8+wSdvmh10TJm4wAUObZzZK
4ItqKEgPpfy58mwPH1BwIgGCxsK+HPB8x0PCbjvMeiYLim75ADDqfGaTFBYf7ijp
e72erzmN2xoQDOgb6VoX0ccAXWcLSQcqi5xuIALVPDGSEUxZKamWYNSOu31uzBXk
QYaSo+PTSrhaEI9wieGr3kr+gFNMZFI/35OZM9Hg1cM6wJWQdevUERZ3v/adlHoK
w6H+c9i8y/19oiuH47AwPaOmgBQ+hE7uhp1va6swZV+TDN+n4zmRlu3tsBg2IIkN
niklULthGuvBt8KM0YZEf6wHGcONBLIO8I1ADWEwktuMWpMVomT/zKcRVbQkU400
KuNH5A+SyXwy9AX0mxBbM/KCIE5VovJDyJLS3KpHaAJyT0hA2KN8xBnMOhWyzeno
9n+0f6+CwHV3xKY0dWuQJc3EpsPSryZ3PtxYq2l4TkWFR6VEtC1fmxUfzxXxS3us
WDfpPBbGBValAgYGe9vp6bThLu/msyga/PRX4aOz9kgdy4nJqGuPlLJZ0hthQJ56
By/3OPL8AxE1f8BvZCGL6TpE95U9ETGt9hEBuepPYveW//stsnUgxAe7b02xesZ7
9d9ITnELVVJsxC2j8uGnkXUJBfIHOyrin5KfVbqcPtUTT1Wz2BAjlvXlr63UgdB6
Smzn4OtDLraLgPpB3u4SphzcoW6HHWJEqVgo5SkjL8vylB7bSwL4IxMHbdaLJHVj
DtK9YPJh7rb8rKZEuIcesUaVCVHHjQURBKZeApfCtRQKQ1xWrkIzrA7fXDyjCNLj
sd24WyLBgeeDxmRyoKp4Xz3xvfkazYHw1le4/vUtGwWHqY3lNciKiOSb9Fie9ibE
+SZ1iQdgukeGeecFq1AQYQiVgCnl2XC5BVKVIyLeXYGMlBqABn7wnXfezqD1Eblb
woULbkkPbuQ/aE/0yKJqiTpT1F+Gj5kkzwbQ6JVdXt21yw1xK4HtUjU6/Pf4gfa0
2InFDNGYw49+2cMSgH3hXA/tvftYfkeVaCcu6MQxyWQOyy6hnHlshX6KR2jLbXC/
NjwF1z5jhIfjLAmEElgLZ71uJVD4oP3mvuZrf7/DXhEA8SNZKUXupTpyQtyKR0+B
x1WetA2LYgQkjiqwFQAwtspDv2iC7vfbcmKKixYtNf0TcaQHHbNVzJRSLe2MGJmA
F9w8D1dbYNubCQlVGsTxRiqgZfwTQdqtj0vG3LAGd3adQI+y9XK+IdE7b5/mYAcG
BT6M12+cbRIaWaCUgosRyz6Xm10/5TbBXzNRVtdC+QL0NiXdEi1Lv0QMVReaaLJP
1p1zPu6lPcp4vpY3Nzul5u3INkQCcAibOeFVffbqrAKIPbAhz3WWKiigsg83iloU
g5Vn5C14WJI7rEYcznjum414dRXR9iYtPQQgSa3Jc74v4HJshBYSg1mhsxQ0OuYG
OJEaAerTg6mFA1lOJZTL+wx79sRWnhaf/Yop/gwpLu1bH4ALCc+FWBoo0DnmS7Ub
lesA2AAg2IVIz0FZZ/mw/TNJxjih6bvFOeQ9ACZ/UJXFbi9H4w0Pg6+rn5yU8XDW
7RXBf3QBI6GxlHEkDb0ocjypTI1TlPS8Vtoz4r6ONvCe0TlHQKqRSP5dE2clZXJa
4xZP51Y6KqSPCqE91C7mks0DPhJnWHX9LFqjyLa70fkWgZW68kpUJKHB2Z7Vh9Y6
nsYTyBGJG6hotvxPfqybwgmqUeLBfdN8MlgS+c8As4Zg4LkdYLNlLlTripm2q/FG
2Z75QvRJ5URMIbVPmFvRTjqIujykzTUdJuHE57qR3INWw52+EjSjLZ0HGCOlVo8Q
8ijW2PtEPAZZX3RX30Y3OQpuCYfLMtJYSD/dlMpDDgD3cuY+HyS/jmUEbWj705N0
pgLEObcMwAahSZ13m0l/7cydz3aRyx6WlA75yUm1TSy610VEB9QR3YiXn/4TXJXW
Sv8ygoMDF3cA1mAmVeL8n6m1fvPXzd7JmgwGDq3S6+GjIv+NakCIcc+tgZ4ViJUz
J790JF652W2CIFMty3zTjQea6Pl1G2rxeYf6hoz+Kdhnm2tBW8kQvHD2B1x95EUy
18js2kicHqlcRNvvfdmP0J4Ij/29RJqtsrbEjqH2StGfSuR117dzOu6KxFigKZiG
57vYwnuzgZLjTJngJH9vNyVQaqyVP9BtQtC8PanFkmRj3dOGentKvlyPe8Oxo+2R
P3ithxkf8nIVWeTmGvapsGKBv2mxUSUStTpiXa8952QIU2wG9fYT/pYL5vUApSMG
t3nEejmOr+Io74eB22DBe38BGlGUFdwl0AWbZS7McDfVfP3TD8wJKNX6A9JxAuNv
C3cbN9P2RuWEUcglUWzFOB3BkXAcLCuIUFCqMntGmQUuwRVC2CaSWv2t89fr+8ax
jyoDGse+U/9DmlDkrHpGockyGytQz4PYQdUlMmtyc7LcQAiaCbElrkGScTSXScEJ
V3PV1ov7xFqZxBxTTRfO1tYUmfbyJriGulrwi9ZcXHt7E/2l8uBgMhZELXaZVWuN
1Kfekkt3iPiOwHUdNWzVCGo9hK8lKjg9Gh0lfG7tKRwD2ggyiaDhkT6bu9a9+OhF
H4jl/oFbqGjofyCuerHcOPWpbS62I5yqByXanaCGICdbUuV/6HPiAlM/Lbf5f2sG
BcZ9sX7r0NF45bQ9X06KEi3OGlcLsEf6Z2Mix73MrQU7HluCO3lOkV9jHlAKStwC
uzbJlAVa7EUJrIwQ1zsHOJkIIuu0rzgt3/EGfcOPqN8pKV60NmVnXYdb2fUSeVFt
uyFqhBjGIu10NiF92pcaoTl5oFF4fPcDx2X8nPOXZNreayLhag3pylfkN8PyRng0
xxn7emacJvpDDnZ1C4xcUJFCoM3/X26l6aIlg0r+Bgz1njmDGUBtEUIa4vSXpAPO
bmfMLpS665BOghYhGb3bhaV3UIY8Ua+r/SlplUDN0t7G1Zlg8ZGsvA4yawSaG1ax
RPBqY5oVCiLuiBd7dspw3vNJCHkwxrKAeNhEg+iJr/5gOj4IpP4Z9WW5LrJzvD4z
xYCj8rDS1A8ZbYQ2mARTVtW5OdY7nZK5CNAh6Nsv4LWsprWtpynJX0bhgppCEvTq
wAOOEAGb812yQ7D4fYTmmhWFGO+puVvXnXGHRMB4jc6XXRUpyUGxG0XMJ/cqvz0T
O49uirBMkGKuIuBRWIIiYLPdmJOW8l/N+1zsjXPRn6sx9A5ZksF0viHUi64EoYBO
73ewpzY1fPbLca8abRY8U/1ePeC7L/XZxTE1Op+ZjJhhnqv2q0ty14VoN9RyMz5i
eGj3DUecS2NYvhraPg7x8DLuJrRIwaT/NXccIraeugnGPiRvumbvSCtTUOqazype
dPTA+I5gIIeQLdiFLLlozNbibmfsQzq+KgrSSS83JX5ipsAkrmM5syxnKEFq/30F
OatkFYekiSDgrqoKEL5VXKyUHIu6+7vEfbxJkgr0cTMIxsFaIhV2qYMFj53UJzri
EZtzL/OkmuZ2AQFWDEsfsuQyplqI84xmymt2xmMvLFehLhTKCv0KUASqkee2en8y
sgGbUepZumPOvet1SGcviPhy3zgbGjqQdFROq9wBYZcwGAAwHTNNB8JtoCmsINg0
V9Wc+5kFiQ5aZJND01jT4p3rWEpY7UFabOcslG9FN1LsaAr8O+dO1Dm6r2QjQToB
zGdmRSopzHlfhG780r8HEwXL89GhSAWo+uDk+rJHLWmVWifM+McFt3Kd6czWovcy
8AfNMDB04U7ghd+mS/fEd1nubofpm9pSQfqiomWlG2NPfe6tJEyizKOI42Lvo1LB
mD4H1Do+zfuJMO4GcfhDXmrsy0k+xmMvSDfnDC+eZsqd4pY3RDTJ8B/lrcbnZ5G6
tA/1sc+guwZ0VyJtdYTw8lDEFzcfx4QgU1TuSyIb1jczHRnx8PA11tUnhiSXa4ZS
CnWRusiAEAgDzPN/5dsFH5+3u43AoAhxvKH+PVoT1tuAFPv3uRFFZm9rAI3DtVCh
HaTZIBgSSeRPKEX/SBIa/s11EPch7R/+djuJpG2AKogPAY5Exi3LZJECAEIOUfVf
uJ3+11WWEVvGYaXkQ1I1sWTYEa/78ugvALIH546iYfgnjhcDkmkFbNNxfJrE3a1V
xG/rjBuouEi1XoIaUSLU2pcUaC71+ew5VsJdK03DN2970vzo1UDtX/9jSbFwUW5h
ww2oqbmPjT+s0zDkszGMI/uDNcVfZ0eT06rn6QY1EjRgTmo075M9eJGaumXx6wCi
96sh84xEXdS4sB/pO660GksJEWQ43KpcGdoG9HrobWoDieEPya7XyDDWCx85ibkN
HHe37fIdzdRfY/advuUPkmozu+srVG++8eL2TobTSgQkus0PgYC0wEPLNBBUIQAW
ueA4GVQ5o/mxX4B/PRIKTkR3W0DbEzAChyVZ+lkGX8EN/Qac/kjM4AuZlItbxLnD
qZzBVvfgMhrRqnOZ4YIYpo2jj5SDGrIoKhy9tI1mUI05lLSiRzaVV5MH4n63aGlM
fQgE+oTNTGxPUBzkBD4HCMY+/FGcNSpKaDcG8BJTbsP8R050ei/Dr2comFj9vx9w
rTrlbCPpfpUZ92CG5x+v1W3sZJ47FfXn0M/nzVb6tbeNkfS7efAZZ0eKgTkUrsh5
t0BPZ0Gj94oBlsSMBOMOQ0YsE33TH553WnExbEzCOW5D8pk6p+g6jnysF2EkOg9O
7m9f6xkzQeEhTtIm9FHeXjOzZKZX9Z2owv0ZddyY206269EbaR/yxecqRB37+QUM
fYVob6eB1hdjzMzH6B6GY15SvpAflnDREZyAKIHszyE1UgIm8CgSF13036VBATcp
qRRP7UMLmgqPL8Tj4cOVJTJga5iNSd8wtdSioMQie3n0zj1xXFco+UQwyYOuySsF
G3HdGHgt/l6SX84AT2p1KV0cgBcfCNONaEcWXWHaGRB6/g44eP1EelaNe8lHQkDw
aVfk3kxLj8sIOiHCjs2I6Pnk6KmgBWWBpY9c6n9QrOc3C5jN6lAVd+AGzdlsqX43
OiVpZpBOUlT4AwE24909w1VUjcpGhPGcqI0viEcn9Cgz5ugeagFtqA4dpCGtdRN6
Ttu4NiwhFFbFhv376vjfcJVEwdzz7BRK+rbEbKtTjDgff6uUYr8RMatNeSeQ6B2p
g3f76MF46eXtUV2GLYtQ4cm2h7xgvMjaDW+zfFj4CVMqYHoKn9pY7Ujx0iZkvKX4
1o+u1ust6UInpsNupWud9fu1051JQAdda8s/Y2B1S3VtTKUjTpzUWwgNiM9mCKdP
Gx0Op5N0YWqbuyB4d6drOXR/3CzcfNVs/eKF/RAXS5Le1UJJHoc+EboL2c/YReYh
kX+lxZ5m1om23vIUjx4z1fwBkoK1yX27p6WT+K/GQwj0QAvU7b8MFfzAgH68Y4WK
KwcVtmZObt3wibGDviF7g3m9Ogk4MEc1imOmAXUG1y87aqmZUPtC3C9sKJ6xVta+
XhyQ/0L9cUPst1mi5lsSwvbb78HI4UPL/jHa8YlXUrL4oB/IoesDFtWGLpSHyuGX
6Xj2vCFYjuIQpjqKUCx12lHPw2ix1lX/pTuMTwEiLj0lkvb25jg3KZ1hy44kgWDT
MFoJJq3BgfVU7gTjp2pzZsly05FrCUp+R4TGJrxAfjXgq7q/sEc9KZ6o371xrPLd
bE+aAHqqvFi/O2Oio4bcwlM2QRt1mNPGtxt7RqztQTDB8IRLidMswvwSo9w1wjBt
+GWAvtz67hNPgtk+6IvrYKWboDNN3GXIxmGV7Y5wexQPQdxEdRj8DGBWJs9OARqa
BocylQJYHzsGfmuGw27jV/2MoxWuVylWzpwDBhX/HsShOWDX7aznOhVCePd5Ko28
TORu4bE3qbtTKD79Zo1E6CKOGy+17/w+6tqQFcej4r6bdu8FReVxTN4DUoUE7eRz
+kfWC9aGqcK/nJ6TmgakV5ORcEcqJm/HgOgxvHra/3m3lDgZrsQqWf93dedETQfO
0nSMdD84/TH9Jtbd0kJdq8EiEXcaCsG4KxrnndHM4LFO8Vd/V7f2xfdU+eeljB44
rLMfB2ZEF7QvZID3XrvUI4ELrfygXR0g7XjL88JaZTIaDB5HdF88XwvoZ1Grupyf
OLcjmciaZcRkUDqPfe1A79SGlLWtS6OgpqG3ZlM/lpcNlTXRPdpbo/rRUTPgJ6Rb
g9hSVnbqbyhwdo0E0a1WhQXXXMDvjDhFjL+xrfuitKrwRCRKFv9hBVKXM+j1klX0
3EYLWzSJfh3iAf4ovfK0SZbnfiCtXy8GfnrIrvWSpr/Q3DpNqGFzU+X59t0IE7my
BenSIfzYCZblVBXLvxC6yNQeLQlA7gnJp9eiE1W8yo4OOIC/xJb0IcCbCjJHlV3F
gcL1bH/KgBipwHn/jV2ucpI+f5x/ThT88D9ElSf8DquCQ3nZCc8iFXIrzGGKSz3F
taJ7ahfoAeUz4OOPjbnAJ9z+50qn06AAtl9wNL54PPxCFZgbchHIT0N69O60YTul
LmnlnMnq4lEksGsfYXvAu8sos92zNS45LJ956DZC6gG0Z8oncJfxfliPFBQRzy1y
itNcdpsDlAEl8e9xzpCM3MPnHBsgnANiTeTEITFknAN9ZS17t76Xg1xcJCcr85Eb
eCA3KYMaagQe9GE+o3Fw3I1ngM4Bc/bDmCq0hZrzJOs7tu3zhCLAPGrsVrsWOMAW
9KHuajN1uG6O8ZKe16wJzyBNiSnKkfby/6pbyTYZ+RyX5olQBmFwwQ8vXH94yc0T
eO5dNsr5xF1Qy4WQUp5tuOD1xtDd7Qne9UNvC8RRpvNY1NXrBg7g0U7T1gdXA0mJ
ORFMLgSBm7qpwpKYITERrGKsZWwiXg989t0g2i9NzslnRZIt/qrJC4Xnkkx7lxud
jI2ho9dIHIQMQ0B5wthIPm7QnNoa2M13jw0KtOBFZ6oCYf5c2DVVFlqHq0aAlkhT
oUL2/MdIuZlzZZ74OaTM94bjcASfvEpEOjEPshdB0aAi0OMVrsetk+Y03fSWAebp
z6mGuBvvp1QJh4mIMpv/QSdQtGJOc8vHemzsKjZpVNTOrlCN2Y/Z9IoGrWh0dfE3
1FnOf/JaSVwbScRnX7/aG/65gLO8kMkv8+Q71U8bsJGVm5QAzAm8fG5cjJ0WJjNq
GFiyEsnyE4t7jAZUF3qdmF90w1ATSxiDZyWh9R8iZzM9gE2b031VDKsQJ7BeLSyl
3TYTSyYIpaDrhLqjHa6UUUvuaOom8RASJODmVOfhQuI5QnF8Yofw+pilO2gMi6Jb
ZSzNfX/st2X8xtak4qUFRZ282wOvUFsgP40u1FuQCjRhmhMW+D7kQYfloCSMyngd
XRLMDxvCOalDHWY1Z8GA64SqDhEERUEqDA6KAwqYE3IZXplZmj8fzxqDWRsNV1Ib
G5wnSJM7wbhT2cMDlfvpo6kYoacKCO0isdGbpZiZBRr8FIu41nb7w4iEf+MvnL6U
F3zOCLin+u/6+V7e7alrYrORLKNMHi65hmp5qwvcLExeCGVbwoKcYVUygxGy0o2H
6tCrKxuQ6y51DRsd1I3n6gZPn8792mrmw2kg2vL5vX0h4xDgFj4MdTlY1t6z+bAE
GuF2yQ2FmoJFIPMiAOikHiR/Yzvym2u2+oZ6ZVyhZrUzUMlxLEaI9m9I9X0VLVHh
zEW1/vB1/k8R1wD34vrCrkvZtlXkjCwJENib90qTI0SqRcjHBa9AK57YNqcu+NVv
WYU7MiNkD9YPuLrjdLx2p50y7z/CJMIQzubFB+4bAsMuYfrAd6O9JgUlyAMuYNsh
XPpsnIr8+1DFcJk6CLT1XqINDuF86Rqc3E+N5YUZPMDt56ANNBLu9jVOffrXrxoK
qLrZNmUwjmvTFAP/rv45a9DghuIrXzOQhMBaY4bTMOmyDhRRu8UXOMi4kxHUbBbF
ctsgricbyTp+Ix70fyV1sQXxkNaI/ACIGyy3r62HoSzYr5XLwOoiTrwMQr5N38UX
QonbvpLyS/8vyuSmgGM+c9Gd1F+PV30244rqeiX6HrrDfPMflscak/iLAKZjFPm2
ov1ymrUCL2CCiv+Vqom2Dtuq4nABjUmORdTiRe41HkKmkx4fVd7mkjCizJPvUt2w
bnN+vIGE5KK0XuIvCCcjdb6xt25z/3cA8zP/TuHI4fZIRapipEBKvIVlS5S5pEBQ
mx7rSyYf8mFBixBn8W3mKb/BlQ9IIagUfjYTArMG/PryS+fR85ltqkz+mYo68Pzf
MJ6ydqNks6yqXwKGN8slNLSTe+xwhdGM1QIiosQkHXx6yg+a/KYLNSZpbrFe96Su
NlbYSkczxcnrmdWUQ86G62PIYj5oqicfeaRzzF6LuZluFKbP/RhRfxg/8RGpg6bN
FvGnk0QYBTFAplDD1bijQTQTQq1bLt3qat0sBsH9gAW+uoh+H5SCpwAAYigPiXGP
RoeUj80DUNo+cPFWIS0CUQu/zXKYuDA+3iNb/scPaz/nZNkAJtY0BWMYmxwtFwvi
6sMOvK2LTLlHo8U8LpE9aKEIq+oQB3ajqJs3Jue/oZfb+26P5WL0nEsU8UQC+SKR
dTYv1zfC6A0Z8zKLkjTdAB3iPnz9trHJ7TL9fvtnqc/0IIMNHds/J+gFbpg232kb
0IH6VGZiNtTNwWwPzWhhU3rWLDSINN5uxImsat/QOROjUlhrLqO9i1/ItI3mA8Di
gptHhnMFRINf0Uky5grLcrxVA+yq7X88k3QFXEzt32UfOsNZw0lkmWbags4EsGUZ
J9z4GGJbB3+6oBzPeYlttiihmAz3uf+QKVjv10yaHkKUK2RwVcsfotiN5UFdJ04+
CfwbnQy3WwQRFqGAft+LTjxAYZ6e3lSXpVW9f7n34K2/8GUOgvrGVok93AJ01u5D
80vtCMlEdTliCAVkVJ+MRCk4eKV+Y/vFOONgR3FQQhPV2THyfejH2FpH3633K/Xa
iJkyF6Q91w3Ak2ZjjvUAUGZWBWFyQgIibI4RF+cc9ZTHGbW1517x1zR717ERWIgJ
EWwJUMdG8S5GvO7C0lkff2t1F2brSCC3+h7u6tAWLfFRo2iuOXVTK5V5cqPx1/aR
TKgGElxe5eLKtgTlunjFAuA0se+Y4juySea+Vmd6jpPFyY/wCZOIG7IUNmzx/VDW
QYhZQvyfo+htifCr26LujFxZxv+ORJlvRmogiQjL6bCVFeGJpTJluDtVVJyPvN/+
Shwl2xo5uSjiLD73i9xOIPvIvzvv9xWkxgnrIDxOeMTRmN9xPIu3sMJZfbte6CIv
PeFapne9e5DO1nkDIHkmG0xh8dtC462OUc/BTn+c5xbmHl7qmUi5Kmd+wHSoXnRC
+lcM91rDJdsAFP7XnKInMAwo1b42NeMiRJLyn+841uw97Y+AW36KZkBCdcdsHGl1
B5ESSKO4Oqpw70FDjXdBGkL5ue0ddkiH5mro7dIPfiIHWRAdTyS7XS29UOfBtyEM
13oxt+IIICOo3Tlkc809WpLg3n0hMFZnGAy+nh1jO2Pc5p4UXOqXxXA8tpeAg6m/
VLIOAfCk6suC5tfffMNK7xesg8UUdCgoNodQ28zeKOygTeMupK6TVL3L9x8gZ4P4
q1xHNUnZIqRTdDqe8T32BYng9Fvq2Jxy648dsLGBwWlbtdXCpVpE34pr6y5ZAu89
vNeD8FGkV5cAJucd0LaPRmQRXEOyyWbM7HWEHv7ii5YCKRQ41cmASSUmA8EHF+jw
jMgc/Hed8uWdfsqUbksRPWGC2ptUVzgJWfmPdR2lPBgu4kehvoEMIJoQ9aCbMzMY
rhyYaDx5wz/VR9ILvj42tlOSPTe26iyppQvTE/s5vEYEBKaTuUkR6d1JHA/qn+X4
iSI8cFCMywCYRNXq35aWoKcobce9jGzavNFpL8qiFyHKyRh/nCmNXFVtoLVjfIKu
VsAIsrQIRDBGLiDSziY7/WYRCx2pZqYjqppZpWMyli/K4LwcRbv4U7/6o5eIRvlR
JbznRd+OMKsYqLXtcs39mpGiEd+ITEziOzR3RK8qAw34oUuQ08czsL47wmeVo3Al
HKUuu3mxzNiHNT4Wo29LjnUZD42kzwbtBsRbcqLBjsKhz5oP1lY9tC8RGW90ryY6
44RVmfPCC2jmFKncAVlPzxKEZUjy+hRPARAdaOZGaJQh+T7UqsnMtLHCPsAoEaw3
QdqcrRtZ+GzxZRmTDT3hbEPrL6/K0n6MThBFyyObN+VIPelR6f8wM21lOma/BLyr
KH6MlY0tozLGJNJz1ySw/Iwasb8m1GbgnQTYGT3Fztz7YBldaBqtQkZqzzJYhoUK
4rDeC20sxge9ZdhGJ5Vm84GwiqyADdLLic3FkDAe1GssKYvVlyU9rIjvP4iY2ONd
RUz/aHvSzRnXdbo0kVwdx8pHpyhYzufiDpn8jppdtrsr60ydn/FgNJ2lbg3XH0XX
a3PSO12Y7GKjoPti/kPUSFQBj03fptAGJ41Zh8/EIWOjxhr6hFwRvYBVTEjhnChs
68c/Qx7vRDRTbQ8EFCO1AU+NPI7FhUHJyjL1kSaAzQ8c2GVhzVTMCgDiP91owK8O
oAdHusm9bUmHxRBhX5PUUsnrABMr+wISx4elnn3be8/nbIayCjI8g6EsJF83Lk44
7goSS2qi0US614UAKw3YJg9+6xKKVM8yAj9G6mBQv5pbJfLYPth1+KSqw4DIo3+8
8olYPgdggto8pW7NrW+9u0pyEckskZ03qpefNxawO5ZVlpyf2FQj6I+xyxDLHYc+
/gfYy0LIHvjHuN0D8AYaaNmDvbcKGbu4GD+loe/42VnKRKSrrairY1xLcSCjTskE
ZmxOyit1N//4nh8l7NaQwNSM4Mc2nqPr4NooEHxniezqjDrNK5glK6hHtZEh2NB0
QY5XYN0EV2gkdhThoN2GFdQlgJFzNc2s/oMglwG7bvByAh94tDq8d7nvCWOcnH1Y
2RTW7y/nkaeEQYJEQdhuger2tAOIneN8bffbHNpEX8JoEv3QpQiFTDqKf6z4WcLg
WiOIJP/r5vHJHyXElF3Ifl4ceiMdZtX4Fuk/84dP8ixO4IRmJsEpOtrnpevdx9tt
gOVVh88MNCwE/jMjL5UaVi6pBdbtkKhpMHct5ZjsxsTMFyuX4gzoQBNv1M0MZnmT
TVZm+uZV1M8Hz7KREYXPFLDxhcHkRCNDXQfoAXTbLMHqFFGwSqi+oT7kDSnhwc9q
i2KVyuEtt7bOxkiO6s5gTR4XSa4MkUZXiIw7RJa7VQ/+qyQbzjFozhqPIfu5oIZv
YAE1wF+Inffx7YvfJvJ3SPVjSi/gKysx/g+oteJWz3M7L55TEyUQDufcFAHz5D0H
xH/trzBN2Jm1xg0x6QIk3aRHeLj/EHQNb6NQ8oh0Uc9yj1WYJTPBCBGyEoKGNpYN
Kitb1mEKRgjPIqbjmhdjWtNcjiOCWfGFhheE9X2kByCWFAfIekDCFxoMmScUTlQ7
hzu8pTmRpP6ilMvED+tFAs8IaJ2u+aayeoZso9cIlr8lr3iOc97Q4+zUx9ZLn/7h
llcmEiSLwI+DDRaxoS4EvrneK30vAbl/ZCIH0Y/rmJWxQKprKJVAWlMm+GPZosMV
RHJ9SUKGXeZAni5qoMq7PrHYa1vrdbcHdo0nTsVG++Yht/IIgw9Ps/pt3wKF+Pwd
qbG6v5IWOjTRBCRyWbpQYSSbvcMHkrMYwypGrW1pM7pMd78uINroRLuDTKzjTKLj
NqsAFUv90PH9IXI/6vaWlfIrGHM/5AbBu+qpHfYMhGM8720IQZRcmh2KuKt0AWDF
cAtcVre7u4nWZfGMhc52PHtLQh19D+o/ZZEna3kpJ4zuzTl1KRZWwj6+Dm50wZrI
bDo1RfpNsmvL6aoK5ZZW+nqaNiRYSv31kP+aS55ompMjZ7UGjizcO6PskejLuNmH
ZRHos1NT4gsXGS7kFR6YnAZFUBbKNr8vkx9fJUC4cudAzxqYOGNmqficUChnI2tS
yWjwCv02ChN7SFFDDz5/Ihayg/OxGHmE++JL2E9ve/sr7O6IlO7b434mxpk610Gf
kj+tXIiIT5CAGsu5IQvGG3VW906zdVndoVuQHlnUGtKDbNuJqtgbkoSXDrw4ee7e
2uyPH6lg0ozgwuTdg9+S0LUKsJp8EDlRnzRKRbZj4dxVpNkCp5kq33xG2ANzUma1
b7B4hD5eip1KppfOrlK+k+o8PihtKHak9og9n7sqQKG2VWNpSNHH4zyrcyDGj8Jx
vzTcRzRjp/QUxLZmvieu39/17IMx4qDYQ/uxUxx8tEmxIu6nPtMBaa1YI20P9VjE
5kX5mlCfIUQV3srIUUFRtaVuUwqUTn2VZNuDYOUIDwAzSEUoecqoO3MxVtTNvmAB
NhO8i3tggTQTQaZzTEw3/wz7ljJVnOBfDxMiPB/cCTw5aJKc0l9653rezuOSDdY9
2yYZ4CKkpilZlHP4X9rxv6WoRGw4xDEpl9LQcAg7fzdevWrC/LNrpED5YofFzMYW
0KVbqS047/A2ih7M0jMQDWRD7sHGaQGayek+1cUI/VJdcofGN28Hl4Gx02n9K86q
ULQXIZplMECCtrzJRK8Jq5xrCPhxgAKfRgjxAjNq6s3B38Khx4A0r6+hFH1AQshJ
HsDlIwwiteY2tbhQNBNF6DqEITPftY68/kQ+6Mv8ChEPIqqjQSe2mws0M6a3pbBc
0GRWWAg7yZmf/uFLOkLVDLZVPU2OhUuy8EfdnYE4w06hYSMbgcUbZxsbhHP2lT+e
ve2h13LUNl9UlX/C3txFNKiHFc9uoJxmAxo791jHrSwwTbx1JWSjXVWLlNqhE/zd
29r88JXLHUrwis9k1jeoAK2xSM74DMMlH+q3THYu+3lb5e4SUnl26M/ObnbSdoy2
bxqJ0H4ttmck/plTBu12Jw4KZxr44fkRWj0Cj+ZnKTy1LgGTCUk1q8BavXS3OtM3
OCH8ZxLRA9ckjspwpR8d5vZrltKt5/o02919e6S1paUmW1OuX2VPafWVavRbCBud
L5XkyFpmSVmXUwvtcdnpQcCtNrBlfY8NF8qIaN2Htnlv+VTEPqqd2zpfwHYusPcI
PuamVAz8PZbQAqdEhDwl4v7WDU248YU/qUNSmkqRoimv1BolcqjdWLPkekCE3i2z
BsXUd6yv8xTAIxvews8YXnWLTdTvzGW0/Yual0u1Qp613YODOihfaDyyfHfgl6Tb
Nqo+WeWmWWwamZq+45t4BbrfBBRI5qAwADxuyttUyCRfkGS0kW/KyPWQCPfPb72N
/beIHhYgmElSuwYSImMzzaT/TQpHBQFLjz+G25+C2QrqjXjhlAQ3+GNMcYXO1iY6
e5JVDcaanmcz1/uNSYi5K76Hzs8504ptrIZYpKxF/Uqfdof7BfcE9PF/psxcTF/R
ts0BQCj4gDdbo/IQTEC7WWHKM9gSpMw0GnnNzndkZVs8mrg6SQf6tHNePHkS6UGG
a2QAgHTsNxrCAGrJKAtvKDcFulUHUlSw4MsghEwoSi5UdrDncimCd+bbT/gq/kOc
I8JJ3oHVsimfXXUTttpb4/kD0H3Lzc6DOEiJKBKKCQe97s6UK+7uQCi/YuP10Bdm
MO7HCBw52dhdN6PFRwT/meaCXdKBPUQ7xI5MET9cMsBFVrZ8/8AtehBkjxW6AGs8
XvBf4zD9NJu9dEqpyQg7TXMCCBiQ4XCjT4AdkeYdiXo70gpRj8X9/e0JJc46pxkn
/2dHRgrliS/OUO3HEf8qmSAmz43k8xCxddGjt+DpfT9Dcmj1N4oE8DTMld/oi9LE
QVkQcCHPfjSSZuplSqaUjaDxJ3tpFZVdNnTuMF7D7KlspPBOI24AdMpI5OZhYAgC
QuKwZt11v8UlhOAh9LNvTW7J5YVCvTRn03ktvymbiSpqYvaL86KZ5X0dIuB+vs57
jpLuaywe5JrwMJdPVle+wEyTK/ZWO5hJrErLJbV33mh4/k9IaLsOF1qaqNUIcutX
BeNyr4sHaNd4zGWIqG/5ssdXcNnlJOyvIgndP6DdSpxIfxjj6eAp9uSDKHVjg4tt
ZQwiYzYVNoDo8xkShLUyfuWp3BatSgDuUJ06uCIUmjqYcbWiQmywmnxvvw0FPZQC
rl+W/e2vzvkWJGr7AVU9m2sHWw+F6xSgSUOUyxWfodUN9UjUZeYTxVBhmo3X9/p4
3GevfsDgKoS5SQEQws7mkxVHnT4SlrAYvkW4AuGPRakGYaLxElKpFRKX4A7fUlyC
nVYUGLZZGjRCCQJ++l+S9kzjhWJ54RIGlmcVjEZHFz0IeFkJqtL4pOERkJTXOdHZ
9EHxpp8glhOQI/hC3UOBJwjf14D6g1cUCw3O8Mge2vZ45XVYif0ODmtK9xIaCuDZ
Ef6E1B/HQOjb6ENB1FuWRvbKuyEPQHx465S5JmdI48qR/8a3CyGeguR5tt01g9+0
iem1Tu0w2B0scHawbscN6FwpstTjJtLH9FzTutSY91sUhEuPPNtHUTPWHyx43l70
RRCBtmivTIzEHJ/fLQrwzfbKoEoNYK7Tue2hE+ui13FD5iLobvK8PTpEESto9zLP
1EtGiQJlKH5PFkdXs+BQntzWCouUrgXMSVFyOqviwpIviptlW4QhgJMdcDGPv/S8
pWnMOZVNE7RzrdwgYniC1dTeMMfMPbyz/bYH9k13/vUwTzg/oo+7EW5c1ZwfKuXs
Vw2L9ep6M/cBfU7wAhbcjoYq54JDNj8ap7outQ+65Dxrdw5QFUCuZR/7umG0FlUJ
awHzjihm3VSC10LbpFU2nx9KrwdV8yVDoA8gbGXIRlFXTg+gJXW1CEemOH5Nofhf
bI4LBjQliptY6QsdGoL/xIG6vkrNSvmu4b9Oid05O2qxgRPl1tE6/1vR4b1XAK0p
jsMJ7WNO4p28BgibIC5RqhGjvwf91bTpV05IJ/JmZ26iW6Ev3KvJS9C7kKizg41Z
mquKAyJZXB6xTwRNu4uhrHHGHvegrKm6aKihzfo9Oeuo9Oj4uFrIN9KGnzhejzK7
CANjKAFjSLVt6919JMgJrrySh2MJqTOuSpfrlX8rtODPymN/4LlnvMDZESjjtQ5Z
qiV1+n5qpHUo94ImgpeOw3FlebIaO/GncaWNae+CQ9LIdQhBm1zBeWzJ8KOxdhnc
J4oS9nVjs6dZg3VGOZVoE7UG/p81Wtk/46m2NLxMAbbbnITK+i7TXZ+vnWGjF6on
P098FrmpzUnUkwR8/OX9iFTHsVB2WPNcR0xwrPe764lTYdpmWClXZyTVh3lxYohU
TdBWtJrKO73OounYFTK7rqQfWbl4ybr1kDdcLWZp9BnQobxwUTLxRsfN01EsWAuP
rNgmpQ3AEOMfT6OOUdh4HGF1biUdI1l7vSSk8fdgNnDLAWY9fL5Tk1kn/aGa1kCC
iXAvroBx2JTX7jd/QV/XKT6B7jGPyLHkv6uKNJl0kTsj3nlNASfuSyRixoPSaeO8
YFSLnDDYWUZFmjAEXu3FYtY+ryPZex1JP/kN6pK9Ipc8bfZWD1uB5ApPaUkie/j5
oPRr6aj0D59bfnc3mWOpHYg4bpbqzgIG2VBdRV9AjMDyCOi/vMxobaQPfwZAfB9M
WfTA88GBzs9m2SrqDRIhw3ixz6wNBEOo7WzUI+BSEOwYTHW1s/Z0vL+x30n3ud4A
r+s0WAhNZ0CGEA5wOOAYL3tdNrz1Tprep9d/SOccpdm3MebaXVCIrUrL9ekleTob
OcrZCHzXIZwiIdRO5U/0lKVkhbIc9F0O1I13ePWgaEiPQfBkh4O8vwE2oMTk8IWf
ufxmHXq4QcjbmO0a4NUg4fi+m1ocQFkWOEXL+pPfqiRRPpHxxexRla7jKyPw8S43
UMjEO88xBFNfL4670LNKP0ffBL7hbFWQV1Hbngauv2lQrvcJQspQIi9MT4nOXOO5
9/QCa4NdFH9CIxG07IpaE4hQA/0vW8YVDm+HGW4+QkpXJQnU/4BgdQ5RqJvaPSfJ
1sa/F/NA8OeOHwCQBxZjiiKE3V+89/De5BEEUJdz7bBLT77oh9RdgIFnZPLtpoBO
un+4cM2P0Z9XYYwcct3Cc7auG5ND5oAGLg6QnZTnvH8dT7r0JT4Gartto6lMYs10
o3yHeyyuODMba2rR9zWoG81QEO7Fd2WQw4khUt8bC1K10GIj89ZNsLZQqrnchC8o
xVEjAwiapLoRMu72f+8w9Q2j0JwG661x3ToaqswjIEYlRdve5Jst6UO7v9+gEhyO
DfqucylaFWMpQlxRn1biKd2lAofhvQLzmwTyFhsKfE0yKcDrl3T3CFKphlevGlBb
U+7PJryL4Ue+0aowGabdexTOfpHsr8Awa6i5jwKq0QmT28HSWXV47TwjDu9ce4Df
tcRvZFf3mjySLaCglXg8BkNieajZP5WjB4/TTUJ+Eaae1des9KjsSrzEfICC6vSM
TnXwviDFyzACqDa5zzIOZ9AOIC07bwoOYVxSdjq4vTstYsHiyUs4n2glJSeLdZRq
mPgfKDSQ+FxXoR7mjQ69sdErBFdFZyPP8t6/u2FoxTuFU2d+aFh3yHMakLteaRGr
N+Pw1rr8XAZwOtyA71W/DBwLyJUXoWzy+q8jkQQftRhU8KgiNz9rJYugFH8uGTCL
JxLPnjDy5nfplnpAa78Q5GONjO6RIEhgvqYRm5pJVPYw4ETypcVNtegOlkTBVF2P
snhBSny8LP/QcLMu2w9Ro3G+DMTATEtZqhPtLhkuRV3DQ0bhF9/odB3/80XLAYcs
ZjAqvdQL8FPVXnYuhVvn2XP6l3g7SciCiNDTEDwhgxif8ukb+XkCNkyHBoGi+lkO
t5ibePJ4F/UshJa4EzZyHxylMfJOMPlsgzYrCSfbx8Hc64dC15I5PDZeGkkGZfiT
EVLvRZMp5AlOBCGY9IkiTv/Cvv6DDO3t2OAh/m/vitnC5NllocSWE9M6XoyfjtYi
PDu/ZIuzYx4VmNH6piITne4AWwb0PTpTQ7dozbWQsGVkWNyvbTC7YKhoROc9P3Ww
OD5J/XfepsmmXdUfO1TBCjZYbOHkOg9rWOnVbZAVKjHl95BzyE6dN3xchGWXytlR
AHFQHD1YZk9xuJrfJ0OD9dxQxPlLVjSdZmlqL1ErpvT3hosCi0koVXYuKBwzDDlg
hkHaUMfJrtEQunY8Hhs2bsyvEdVQ1ogYECvgQqFeiakxggkqutYKQmeqRvu81WR9
9obIHNuO1hoh3gUdx2+svHUaQlBqbIemeXX4qq5UEt7Tvf3Y/zKXELnvi9s/tmJ2
XO9z2WcDAiNcAIRYvP/qiYLO/HiEziSRuEqjOeZPoTo6S4oaa6lhw88ITGYm+icR
HP3kNKeCqmQnoY7RSP8DvGJMXfzv+0pm65LKLqPtfwBHwi42Q9TQHW4fB6WW3haD
byfomhHnHcLCLBZJMgRp0/MPudM34iQ7n+5Yhqkk7D2v1RbHpMyWe+Ln1XiITGJK
v5njE1lSzzaNHgydtdfXhB7I7fJ7PuY8XnMo5cPtup/h5wkxAnhq3o8FA0wjZUYL
gilz01wd/Ll++cw339ySUEQr9v9pNt0L1TfJdAheOsUWZtKoJNE2Ym4WJfUxTn5p
FvvCup0Ff/WTH/NZ1Bq4kiNzNmYKKQNW54YJ1AkAeVNdFHxKjlPeIlup2yobSX2P
d9fQ2PTuHBIeLQWKAwME/gaGdBiTdVi+UjVX0nzI0gnIo5Ti3b3grRD7jGANbnuo
ASoiLNia9DaQyaIc0LmzwLduUUp2lCeRj5icGRay8bBZehp7X/R0rZKtTnNI6zQN
sSoy1923SRkghGXyaBQTbV96OOT9A6x2I1O61OEfRmYQy6eYIWV7WPQAFguxLvH4
uIublT3pqJBHIEjCk7Lys5maDIflAZqTlgzdEluoPDl1BWpfazTVcvY9qmN9Ul/D
DlvlnfWvI99twYo9IDnCINZomXD1ud/5CZToQa3Rwg7ayQB97VOWWSDbRz5Rp4Tk
UhGfvlDkatdaLBw1th1d42aRtC5aNbU23tKPP2pMLH0/oV9dL2cWonbJYV1cr0Mf
GFc61Nc0KqCJfdyegtqRVylCJdOyVPXQv7N1+aj7hwQ46s8si8c2KNZH1Joxq6bc
T+ldk49402lOtPeQQd6XVW4uaiWNbvI2IY3t1dBWHl6dwn4fMtO3wKhXUAGmsvTS
ms47tjoEOuPlTq2FTdwlT2NjFldc3GkyEvnKmeIKOMxK3uJ6tKxRb5FGNz7Z/Ptn
uJC5XHI/KGPpqMZO8hzN645xN2AnpBtn2NNTBZ3T+yrwUs7oTB01u4859c8uq1FH
OPU2vSKHRC17oTmjD3n8B0R5GymL4iRCIf4oyTqNlrdryp1AQzaZSEodg3PFpxPE
7qL0c41X0cEbkEFh2aa8QaEAZdt69tQrzcIbResDXR395NB0O7zRTUAdAVX0xfdt
1ZpiL5LPJvzbFcepI3Ncjypf9+679QumtE0P6yQ4fi8dKyeYk2obt3kVJPxdblPB
wTDgevHfscFl3LwEW5fd56uGZzPZaheNzGsO5WUYI+dhXOkvLpZ4b2rTgot+3Ok/
M4AKLnuDNCn+/bjHXprOk1+cBXyn/o8NaSAv/sDGYjxhAQW6CPUrqyznA0Ar+Zkh
SpwOBgvkxMszvriVg93BSNiFDzLvn5qObwWTuFtJuF8QVf4WxegwnSY4UcaW/38N
Bllhg8ftAnZNIn/tc+rAGTMqDhn73Cl2uf8XpFeYoTqn0pQ/pl9Ppd3B55niXMT6
38RpG4t9Wq2Y8kGu8MX/YocJCpVo0aDRl65pWOOQp3SJDcCI+EsBblRI7mrndxGk
oxH7BpaYKQ+1kkk/oV+0QGNbYT/q6HZh1no6YTf3OAVdrJ0rka6qlEmxfytG97nH
QvFK/TKiSqUKIX/JJfFQhha9LDBhxFb8IUOiU8mnTHR9rC4iH3FOdCmPYhL2dKln
qHciCvlL+outgYWO6i+yEtab9v23GUF80FUlqDA/7wFqnAPe7alFUy38mH+2uF9Q
Qdp6wwPfT/I6vCSAeWJu7agq8NKFuTN2o36cCG4WVBN5DUy+aDiolcovcn8Uro7D
v8Ct5XSxTv6Ao+/yJfFzJQcx5aypve5T+GArRHLPAxQQqyUtTqjfjShQ8rYo274a
9OCbC9jTI8UZxEn47lHk5gIGZjCbB97OeAPhGjfmD0EFuqnD7Zq3Ms5dBLuRDg8b
Zx0LyFw+nGxNFUXd8uoQ3VZHPyeeg4N71wKBv3UInnrMcXIpLwxsqVmHXu8/+N8o
vpdWF3yv/BoRQlPetreLMmXedtyK2Xtld6UVaa5lGTFp2ATVjRefXGf+yXNGNYTU
Ub1S9XxHTPgaGN1Dd2/7+We3nVYtktFT6gV/fUIcsKD3d8jGkqGWop7BXT2yh7ZN
xk0nziKbDmgiPRA+1FuscvXKsWx0jWAQFAhaJMhfG4EjQVGREwWVEkI8XVqhB4af
LRJkDim56WZ/o+B2VV58s17dFrXkFtC3oUeVvhbtjfxQ5H7dHkobku5be6HgDGal
aPcEjmKbcgLN2RZxHqaymg9pAw3Lo6O/AESa12W2R0Go0zJwYMTAo1UYlB/Nj/B+
8gZmYahtjeuMOIWcaoBZ7ZrF58Bgv8uxHSBO7q47MPvRy81d2HvLDt/ndcd05beK
i06QertTYHeFEHJ5iz0oHF2SJ6jtkw4juqyuI8FOCMtzobbEfomaMWPjdiyVu4H4
uOepwoxk+W87o8Xxuf0hAwOYNttfaXOGRHvULhYmSPK6vBzcye+7IP+mHf4yvW3W
J3J4jUudtZlljjy5jVJ5jJ0xJDMu+WYLGByx4JIYmqo1HnrfSDd8IUmBgGwE+GOI
e3qF+8bF+k1t4FRG2YzdrgncopQDRc6/SD3JeUBbkWHO+ssSjkOId9weuYUUu+a2
XO6+kQIe0GGlPyaRawfrPTLMho/BT7n/OWr1QP3VZKgwa8vPZuMYVOskvnumRTeA
i0Sv690dwTZoy5suWz5BEeynqLrmMiYYMZ1D+Oj4C2/27Qw5hbI6hnKbR15uMjrw
M1hFKyY4S8lHG552RuejSuHYammGiRQw/it9CgeUxd/HFET5F4lwnNt/dgoYdFnG
FzknToG+53HUlVG0zympkmYNhPLTWt0YkBEWPMk77bVu1INYl4gX/ch1nL4RudIr
Gt/tXMTBFhc6nMQVmr+gD5mvz/mgOvJv5HvBCn5jbZ+7f4VYAHZUglB6azYvnCnW
4dddTwj2Yj2A6pY4iNLrNrqqg/C9v72ruEuU9OmsuUjEb4UQ6UZva2vmc6+dd6r5
FXyvmn1Rxj1ZW5JbxiDzOrXLBMFknFrDwdbn2kBThNUuscC8ekYNI8K5bk5N3k4K
SL4qVem3GaUjrLnlmXpyWVilIdjHu4nBm4bS/uQacsb1+qo2QpEwi8qWG73wHk5n
IUuVvQAQh1eF1I8Fnz0ZJcdrwzVR7tC2eDZyiWeH0T4LcaF853eCy2g4TJbS6wpx
8pQkBmIgCZjblOGZ5z2KgFrchukxVhtGtE6pXW8IV/Zheqjzvm9zUphIUKWOMiam
uL7hjd7KSEbS18koSxgJWhx1ynLqqlQ8ADjwcZ3eq0vIh1dSoxdDZ055lRhfzVrS
HaKe0He0Fduu3ocTQpF4jfyyM3EZTaJ+EgqeIfDpig1+bslHgIndA18zQD9ebpS4
Jlx+DJI1KgMAtVjkZ+0Lyr8IaIXL3SAMTgm74kP2/uhy4GQnVtuonhRFGiUVYrHM
9cleoLS9muLvU00l33M4eWu+bCtF5diHBi3XtCcvvXvXedjMUOYWYg+YOnfXw1Sy
oRTHQsdoUCDAYsF66gU72djldbXKaZy/NCr4BhB/EFSPIxOBacfhMMIiYJAt3xSF
qqD0HnAq8hZ04dR7sjkvbukeRNYDsPxDqSpl9P1a2IXcpBK57StZJI0owfd1EbqE
MI89br9Jff3eY7yOIYYjcm5ljuYyzDoGj7AgveU32rajQ4wWbtqJel7cN8QY1lhW
qvtu2aC4duYhRH9+ebq6xTE9z213wGErHgHUKpzy5JqL/aScSdTJaaLV8bWNvLDi
W7qeGyuF1qmpeAGt7CVLcbmJxIZuexPpsN63/sS6GEI4Er4pUs3R6qJD9+ZtS3T0
fRZwz7JHjv6shfzV4RyjSxoVJgGCj8o2J8Mq6DxyNtK1oHErzpTLdLRGFRlA/hY1
hA56LjYs5tgVAApKWK35bB86OfDsMNTAqxlOdU4pJIOa+rOV5VAcSrYEgCDHmhNf
Dr3sZjvfMG5XxiUTQOzKNciYPXtbR9f+diJ3880lY4CwnvkJqdr/uXTSQV8O23YD
dYz7Ise0LwNQKDZqyvV/eYDX0J4xHJbLQo9hTBpgQsACzDyFbEEDb47D/70jbTP3
wLaeY1TNXOTrbloxePFxqkioNUEGOQBx7nEjlQ1TN/cD3gfhoWofsu/d/f9jgUaW
GUuseo9bqYblriXwFAzNyf/9oJzoOqpTW3+lhSyBKBoSnQV0MZ9tt1P1PsUgeUd0
Vn9FFZyNSYyyKzJO5JwZQt5nrTJcTYd3v9qNYDLDwz/Ejj84HFRnrVZwS8ZnD8Hh
lQBnhcXQSnRgr5BQD21P5mH5oU1+YpE14eXEeQ7nQCr8HCAL25NtVXNGgEMFCoFW
aWkbsZheRMmG/8cyz6s9iFxcKUO241ZUFjbwBe+C+2DOc6xXnL7Jp8qituu12A3y
teCyp491PeFdcs9xW/C5Wplaag+WrX64WWnRhzzofJSfF3UcEaYZkkCRQm+IbAIK
vTEHQI54oOGC5TRfzZpusqMdFDZY5gCDt+sFpoJ6hApEDF71lj8o5gKnfYyZySsL
wAfgApNle6mq5FT8TVyr4SaBjXAxKgQTKol0hojxjAXZcY+MyWSKXSB4xdE7owFP
uqsPKaLCAwFlYN9Viq/CIAoi5hZ5B/tG+RvjqIV4TSst0rLXW8IqIYpVHpBnHEaL
O5g2m8/GFM8Bzd5BjSO1qp1Rldi+KqQpOnQlQtuCZwAAlG+re+Rv0ITmlr6g5f9L
1BX3A/HQT0vHM0m01bY4wvarjV3fyBkpAappVSoeSLX+8TniNJV1j2uchC3blG40
pwbX3WvovnergLVnbnj643E5H/Jb4wXD3c6axsF4aygIuIZNUe8Y3HWPHyGt3XII
1yZc4mEo5yypwktE5yCIqD8xZLvAeKwYKG1Q94/04TUc2vX+0HSwqr6s/RZ5HW8S
vrjw0u0pK53xo2FYJLNJpt7T1YIe7HL5WXFpHlYZ6tbWiF/+daOfs7Ncusby2luF
G53tWFiOnqMVo/939CnEbd6jq4+lpsSpWF7sggag3HbikpQHgu94f+AcpA/cQZpm
Uewil7E7zDlpYMn6i4770qP9fav9GU2MA1Qnvy5LLVLNInwW7ChCSmgwrV2Kj2PZ
CAj0GntiDJk7ykohDKW1UGQHIt7KinUs28+uuf1NCsuXbaydSurfRYvw6e4+IPQK
p9MoCTIf/JYLNPmsJMAG82FDYFLCBlpdfmkXZkQUt+T8bzwCzitiic/XH1N4KGgR
NVvM3XrVAl2lzaM264UoRCb2GX48sOj4oAwysyyfBDnbZna+1sM1YaiSSG1xSbti
HrqBNvcv/5MStBanJM1i26BbsSK+kFMnBUASYw7YsX4/5QMBtpcOswff0GoGJzCL
sElAvRa9g5NGLnJlpNgBcswGCFoxaJPWzezxZqg2sXozVFVTSp7vaM+IEfL8WRQD
6IXmeAdmf2Qgy0wA+I64VNek7Lc2ILT6OuWbuCiCU42yVW9JJ6mzCt/HMqrHNp6A
KKkHW9EWl1dFQ8QAvVGWvwaA69pdmu8NykBHRzwR0NfiNM3us2pKl514Cmp5R0tz
f7KMvtT5uL1sRFGaNsEUPM9zlamwJBMmc3zm0HbwbMEGaMfJhx2b/VH4OTgzT/7N
efsTu22kazk/dG7gNNMRI9OKEgHlvZlavFBfFQ9WtuMRYz/2v+tIrui3gpLS94Q3
AFDkehShm6hB5RQEpRe5w59dhbF0E8X+mqLdwjSaXyDIy00h+6EFfqk4xM8nE+Tk
RC8I9816NXX4jnOO6MHCtoRMzeAMKUYCXg18nvoKh7ordN782WlFX2WpRuJjLhj7
pDsgtviaDPVYUFYqgphwaCCR7nW+4+5GmiiZ+duTtpiThmmfJ/sDPXs2ZWx12elU
F/2q83AhdZRt1X897SgQ021OQuWfSj5aRcER/X7ZSnxfkXWtUB6itrumIU9A8Jxc
NVj6VfUdMR+lCt19CMOVas5AxIE3vse8f9Rk9KlGOCrFjTzNHQmT77xro5Fw4Jg2
5O0bPV1P6o5IuVLTev7hTm/zpc3wTJxSaa0a/hIHx0JTshTowoSQHEvc5RHfH4eM
5RZA/qVBgnn41UVHqBHU5xzJnO+P+akYj2cShRQMUa00brd4mIK28rFrkB0jYcHW
9J+J/enUxgoPJa9eFJ/VRveNja7JGGpiJsft23CEEaxPTgHpKVueuB5xJZ4CdCFl
r+xylv4NwAnzmE94ezVucytAAtcnNNw92xdec/Ff5pQJ+MzRp1jItQie49+Vs1kO
mBEKtxFsGOzQqtyNGjnMHzjoh3cbs39KBX47pK8G3g4zZSeX5FqMX1a+Qo2EzcVg
wHzx7e/tnW5bzec7eWiCDkbD0ZtMuAIgamUNxnYX4lx7vNVtF+hgQabb/aLEzb6O
HbqNXJCJvS3vqsJpu76LCPUP9OP0x+rVhWRu9HDnOIfTJfQC/CTwP84lRIOD0QvQ
3oOSdiVIxK67AM6ee9we8BeCVHoHQ5frKLgCPIQ/OEbIFBqukM2E5v4zHwT1ypoL
W4jHyeLG2/95R86KzAxK6vXzlOUxG9dy2gsXFQLnGJnFrgl1vDzeSbxz+9J5EowJ
2r5aQ6oDlVFEO2jCFDsOXDtQhVKdU0ZPTlI9sj+YOgC8I5d5XelrnafAw/dtBDe/
iPX20tBQi/feDoKUi02ss5n98aH+FD0eFmAGm0W16KWlzt/KHWHmc0f+dp1APuV5
clynCahdQGvPL6ncJwuEHW/8mBH/fUqO/Yv58NAk5wM8ELwZ7lkjzvbu2qUeCFOo
Tu1lMFCrSGhWHJGucBIlubbybb+wAfCuXNmWTRU7JbID9gNAx+Av0sxCkCmYDNuQ
gaUnjnd1FuiSGePiQL2aezCx55bjJdErDVcVG/JzyvUv3P5OJG3cxdrykBEBsFZ/
U9j1S+PCEGALQu1DHeQ4A6+L8vyB87FMFgt9BHYUE5hUcfYbxlGUV3nyv/R1N09M
ffEkKY14ycY6HBw/NlWX1BWEe1cpYXAaDMvuKA21e8DbpejpKZ1v6fHUM9vmhy4z
NBq3qesJfm7vO4xe5UTYQ3ApbMItlbOi4CbbzWYoHEhln79kwDmKF+MWj4XSVEoX
84rVUo8GW2hpmKU3Y5/NPXJM4LBagUj27sH1B+JbTXHRhLdO2Zo/eDpf+CT9zpq3
TmG8v1rTFsaVwD8Z7dBMU1putu3SVvHKt3Iv7eUMcL64nZLPr3fkpsIpMktl4pAv
HabwKTVJy0/+K2rqrIIuZ86G0Qu2TtjE2JKgUyAPIOYMcnbrBFf3ZaMhQrVKPEW8
YFC1pXDMpSnGxMBEzGzNun4SJJhtl3yKApGWCSkt9Wp4FAma/Q84GJq1rGQUcwJP
G4d8qyyYL8PJqK3Yg6Wfzp8+SPmnIMcaBrXNElyIMf26wX0FlA5iQ7YHIpVJu9DU
p8Zo+eC/QPOALiZ7YyMMsQhOZgrKjwYWzS6gCMz2OTHfsrgNBmR9vLKFcDZMuNCJ
mHPFBQCEqNZuaJy4vv/6+JBKsp3jFjlzBCRDMt08jKaWrXF2/uZl2dCC2BLHqpcK
c7Jm8/HAQomFa7oGfNiY4VLHb1qvUMXdCDXKIfSH+Qmhy7peSUyxntQMaqVVkAaY
bebh9lNl+mhOew3QeJyXVgSunNJ5ogRXu7Aj9u5uZk0Lt1l3lQs5USjKZjC4gGWc
Ho4/e8go/IKAp5h29EpJytFN5aGPCx3DqG3Z0TwEakPHfdDvW5IOfDy8p9ZT03qe
XbfzLGVSdWtwGNpQWqdmh5gryoYZ02diXK7Eh2dslS7b+tPlaM6eRw2Tj9YgIune
ZW/ePkLv91R75OQnU89B6+m3YO2uAfiPa3qwE21U6IE/8KwjQH/Qstht/ezlm9Pv
xyViNmw44JqI1NJU4z/2rU3JH9j4Edvp+brtpy9WsHyhib4zk+b+7yUnoHsGB372
8R+Mv02sPcUZlv9oXY2X0Of5MqIEGiXV0JlXysfTzXzHygd4p4gn8tKzhhuBrIKk
M297x0Z61m+g5jE4Qr5WCWOWPVYKAE2d8O+TtZqNOTrMuqWBQ0Q6f7Os/vkm9LAs
9o2p7+OY0aAf9CLgAXU8AdOnF5+NJpwu29OH+lLriR40j+d3R3Cf1YQn/cwNwRqK
Nm5iQXlpPv+/t5o1gEwPd/mqCGNb+OGL3+wMGHOv1xS2Ncy1FcuWrIRKY04moOuv
/h2usBkUn/8Xl4Hr+RcHeXzTV9x/v5A8kBS/j+SLolAAQxVWMZq0/qlIe7YfGO/T
u0bFjfgp3mz1l9whITIKabR6FUowbON0lfu1kAZKPPeZ98ou5a+9Qo86sqEhL47J
O3uZFTuZA45cJwffb8S25pgu1Y8QPjA8CgYUyxsO0qpKSWb6Jg7LyDUa68zX2xxt
HrZoWrjUvvA5LRI5GWyfRXTT9Vy1G/Kn2aCkFPBAr6YGgKMV1KJBan16mHdE/ggR
Qb8YFMCqnD5RIKgj/9c/lFYedYF900XrkbqPau8Oy6dNEjrpdSdbnvAkMV9CMmXz
Ao14mzL0y4JDBEkNkz51wzvBH/0YoL+o8uZiHnHGBpqSfe5k/A3bxY9hcGKU+0Lb
xzWsng7reRDvxeFN/NwCttY/0dk6ygnU3ADeXo8lNH1qirMVJB/+nXfHo4s7EM93
z4zdmu/eojvyAHe7C2YVjS7YwxYW90nsrdv8dP9fo9qvWoxz3FHgUSYHWqUnHwDm
+OMsYEPf4RrvR6uqPzXOdZPfBeUzCIzW5ea3i6b6ITsVtYJbAWI5qvDETZwBzZFJ
vwbyxt7OU1I+yRLNsfcYiKD4Q3RUsm0bMzWdV5pvL2f/ONP/rTFGZQtCwQC61clI
NWsWeuBzhJ6aOkwwMH/oNz+L/O9nrhdcaDCKK6R6BmaoWRMerRljWZH/vDw7Eukt
hn4tF+Na6Q0dehNL2yk6HBi/Is/z3qDRM56d6yxMCXClHyUUg3j8ThH2CzYH4wYZ
MEyMXJosna07pcbm/uL6OrU1FX0LHHQUBfI1y3FEBGCDQWS+hHFI10G9XKg9BUkl
KgVnv8p8Kiv0Hej5VVAlkttESvmj5I8ChuMe1SBFNEO+xGpQRvNqVUN2HKuP+gyN
1YdSDiRfFm8wYo30LVi1l9QJ0/pNnhwvZJA7svJWmfQ8zWE4g8z0rMJ61EeGWvvL
pQU0PQN5iDAbYKJF4MeqgUWLmgXdTEnEBWqsNwzgx8ikxGNiwgWhsPDLkcwXtUqE
ndC4UzKsfPQLPDeBJr4SVF67Yw4E1M/FuiN9p59aQ/QlNdbFNXCc8mSrmcmRXN9X
snBLC5hy+DsGS09WHEmIvpEn1Rk1dfFkR+IpZs6gUSJBZYscypW3xhE+DIAzqkka
z2zzLzNNf5YRz73lr3bXgzSAKirp5Wzf/DkEKyjllpYBmYZLdiTuirtiKH+WepA9
/St8xKALVCYz7SGdgVvF+eGHb82TkKnewlgCy6KsvonNh4NDgYl1VimOu80gn8Z+
P8MQ0egNrvuvQ/fMxjiwitIJey5HKpoMAYDuk5kV71Dds4a3G0x1lLJLy7JDp+Q0
TOkETorPvWPMlvqNALgpuIDE/s1+td+Q7/b2ny8cCrhdAfAsjOjnA02U98oBUIIN
QtwIAmMfibXBscxogcI9/xrnwJc22BWefLJRfRMlkT7PUlD0stl+E5IBha6IFl3l
gCCVmG15IdM2CTnmLHE3znd8+zKMmKcF1lmnlX6qV+i3t3HV0o7DqCwP3c4/VDXA
FbmgiQW47lwXC3Q65cw3F6lI8s2QYS50Yajin0US3p3bPhRjUDOPeA6VoYMnfxim
YSQ27o0TZ+CX30uAtPdW9zPNxWD3s2ifln1PSA28WZVIjBKcfUY0zQhYZ3NoWq71
DPhB5+Jzj1WIpteqz6DNJBPgXGGjdk6tn/B0UJ0aBnk6CU/VJ4e908royO5OSx7N
1qbZuPU2AXOFi52J9040ntKEv6FGsqP5iO5jdTZ4HT5PljYIP6IUmR9YaKQpZygs
BHCDzOPB4GueO5NlkDGRHSPkeFGy9T8jJMNX/jh1cG5bfhgTkPahDrWxwdlpfroG
eY6L9KWMLSok+uMTfJnvQ2LQfu1uHlZmlxIHtm95wpO+JwHvu2EtunqmEo5CWF1L
X+l2ZmSOTaOKEYQ8SNLavg==
`pragma protect end_protected
