// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:05:38 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
c/K8CUQ7cnm90bcIZGHUGKKJ2SF70DIwIgn3Ml/jsfo57MyIIdt7CPR29SNVG9lw
otNDRg+UUkXoxi8vQgmthzxD9Qp2Zoo0kPUyL4SX/hsNBXZgmTC7yikv0LYD74SR
Zw+LXekqQtaokp7ylPh3RW8GyBCJ7Scohixg9BjOhUY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 15904)
Cpt3TI3Zh5DGczdKTixtIE4Fj3NFhkXWQ/RUVvszkajXb2CQwr2GDmmAcUPr89S2
6VmYjTwvKK8hF00nKkHWMsv5pztVariF6UixWGHuBIg1Ml9NeF5IjQJUAabgdhh7
53Zkkq5WiMfNXS/qEerqBjHySADg7VAbg2bYWGyKKXA3wsmz2u81q/SRAXzCiAnH
eqzvwcgQQXzxoiHI49tw3laO1z2lRBvqNvyfUpq0NobUSzq8PoQ1ilF/PyiOs93f
Am4sw6qJnbJ8PNTBJVUJ9IR5/nvs9S9mcgG/JP146p4IH5u6DmPUXdL113smKW7X
uhxLbYulnWLVPHJ7u5tz5SeYkCTPvYRpCqPvTVlkS41Gmc2tw7ZHELx/eTGANJgc
Ex9ev0rHg4T7GyIR+XYeaqUfJ2679RbiFSTzAF64BkVjlmE8mxSVZFsFDl72R9ed
2HPMRKaYBp+B5jpNVq9K03dHY+/IPD5xv6Re9AEFJlCzDahZrtDsOpB59o1GD/9q
zpZu40jOGa6fQQEos0WuHcnFrKCgSaE6ZRFjSzdyEyVh1szhr+sJYZycgnav64p7
FPHaLFMXctrhtiHzR6hXsPcOg/7GSBjv9db5tLupyojLUhpUtFcVgBjZHljUMP66
48vmRKipwiV+ckjrz+IHnNxIZLuJEJVKFbhHyji0/l0vSyiT5Go7fAn3+HWFiC29
B9XKd4RY/Fd7PHls6BdIcF1W7pc9MvRnExoZyu5MMDqYDbWhE4fO10mU49ESeMBy
3dIn5wNzPzaZFOxOMvow5CKHd8C+ape3Ra9hTExd4k1f2kudi2hrhDBt3K+hCRbn
MhJJOOhe1hoREa34ayEemXMHOktaoIfy5wZO+TT9enPffeHOovbixSzyNAK5Mfi8
cBjnfg1QrY0ytAOf4JkU/VfCZK+Q29oY7R3MvNAHev572GQ1I0YVmYrGEdSciVPE
/xpIHjcZ5u4Qri1wLOnW3dAaZoISPDmIsJpnrcYOx9P9RoL4PPt2iC0df3g+M2z7
wNPLLniuHtokGGMSK+Wdr04MW+6g/AbAJvlvWDG3KzSvovVwG6E7Uuv9b1u8xGHb
mT5auP4rfEpbb/zKkwOfyqas1i3JrOj21e9CSL6FX5PnmwMyvf7aERPem3WeoHTL
gC01SktqtIzjM4XfgKPVVm3YYnQFxOYoVRbbDSc7Q1t92XVX/qHaobc5xdiNCAqQ
4JGeP/SOoWsvh/otZNGrD4ncDopJs5I562ytNbPIxh1snjK/yNT6E9MQ9lBe7cnI
CZi3OGqIIuRLYwQiMBpjuGBYTGCqQd7WFeK1S7bzq9AvoovRojvFyFmgplDUp58v
hpDz2CSwbZHeKGmtkN7TffPdnaot65deSbq8iaxkwsSpQz79mVXL3jGzmcoIQiM+
TVV6pPSj41AhG08moyaBqjHqBYxC/RGKG2zTAC0izs8coFirLZdmbRS06agrvpZ9
HL89AYRoE/2OD8lA2Fr5TrbTDR3Q8P3RbfFKa7j1NyFujT/FhA7a6ABPBMPhxupb
M4fIchvKiqBpzntXczhG1PoSuoUgfWDu00NYhvj8MjB7/5C29WElJTriqH5GprYG
L7gWmltE5/A+adPPz7lh4IejcQt924nAvhow4frwZISYhUdi6665Q530yLZrloG5
/3uEADspBJNTe9HlNkNRy1x00KpbcnnwaGKJ3hJStuGw6qwKmB51x5r6041TAaAf
qoAPS4zDJCkCPDOTIUticx6CRzWLXLBXE0ygGTMNdJCGappD9kswQkOcBNwntIRo
0uONLxC7Ms2FFu/5SqlAjB/E/XZYJiK4TdR3O1XNR7jLfU6CpZoetAjyeVAls8lp
HlmkJLslIBDfXOPaxfTHk84nW+aycPRglFg8t9cCrj7doCO+WAWluOT9QL9ygpLe
pELJULk2XOCx+GN/ljHgbk5HrtGy8g4Fk2NhL6hUp86f5tXvmhl2pMIkW4GRpZRe
hPHrF59d9eJbHYV/RpDstiMdWNk9bzYqxDnKYFS3AqVWXULOaOJv1qKjhfz/KXP/
okf2c7Zoa5jlGzQMCAqvqe1f1EA+CW4xJo/6nN8P6hBYJi5hiMx6wwYqqYTkzKUF
GcKGlwBaTGz7R4caUb0yR1wRg9Kb1fuUpbKdGsYoBzrjU7qILJykH4NdgCjhYLKj
d4zvn12a3iznUlXRfY/MhH35YyDbig0v1hdsGSgLL2S9iqqUIjy3fqWdtaU6hA1w
02WqVrw+DzfaO9FyK95ry4SKOnUAC22mGmcg3VrMoesBJQnWZKUACOZXVbkeb8Kz
nz3p7k5HP0Q95TFkvsJmD0ehcP6LXjyuBH0cP62R8WFOkq3Pg7l1yHpwFosrID5S
i2fwl5UWRm6cY2+Jo71bJEWW+V7KF5ElHdBGyz8vcFgdviPvhi7IHF+nMyyIBEsS
Cxer5kd2u5LqmOpCmuw9UUmiV0R/t8UNYzaM48cOpS3vQDioR/wKmescx5vhPSTj
1TQzo1/6pLHZ9E3/ierrLTxSjgSBq0F/pcbn8SA+YhokJY3iSd+fIjn7/QBXFazW
jHJuhqqVUHkzUR1x50/YH0WPp1DkG6kElMNnREH4GvyFQzTLDx9OGO7XVKVQINMt
HC6SVLqt+1FwqkY0WJ8EWHIS5wzajlwfBRCu4U+yVPrziNrPT1BHtehEfexeo1ex
2OBpoWOHtsEoLcEtdxfHVYdFre7Q4D2KMEdZ2Il7RJyHmQ4G2jdtKQcnG8xaxC8l
yNnWsBFsoFdz+S7+rinQaa70KrRK5aH1D6BdMdYQrSmk2n0hvMtk9N5SrwKgcVo7
cXSo0ahKNWlzFfWlRU271XRlU7faJ4k7rmzk+a7OhdtS3U94KQiSpTgSF/9I1XF8
p8PRvreYYY5XMStrg69UWuK+w9INUsK1mDlc7GlZ8frA422Jj/8K4KfAD5kpwUPF
JfrXZ7qzKmjufHj6LX5lqzbIlKy/+wrlc2cMZl6rYqQsnWXR4lwWw8/2doGxH46b
91sL9rws3FSjw09ioN7Kjt2rue3621wCTYhLc5ZQsrxtylDXNtd4LiVKVDVJivD2
SlMvZvUvBhnqFHcZxmch0sZrMtEhG+pmZeT3fH4j61VN+EUS2zbaD803qhVubOPR
ZmquYNBoZgqAyFHeE/E8sht8E0UkT94JoVV+NyyghEzGFQO0SCmkmemMVwDH7ThP
4ZTJRHJoVGrPwvKNAfc3wrlwwMYM4lbVGcmVFDD26iGYQj+VJDjmiwlXm5V9VBbm
Mpl9aLTZAuTZADLq82RrRrqogxDzgLJJZg5kM8dgBmrMeeIOPN9ymEuQdrh6bQQu
qZXlSo3DOmSAPbOL0U9ZTojEgSkv6Xi430N5KKAUSq5bdcH900nl/VUtiov4Ummr
e4D1D0txdrcX/MRcCCfZwiVkgUwBkYsAddTbf8pw6h2OurEm1tEhxZ7icAvkjLQO
cmyhhcyPGnMeHmIHkRakwCl1pgl9AdIV7nhRQnSXBrgNJ5/I5uNDogr1veDEvzU4
UqxUGXIMBj6aCHYOeI3r09KqhRu9ZagKwn66EC604e3YmocP526jXVf8KFzphbDw
OPqgFHac4GNg/bSJEK310+GRme45mS2GLHcsq667DQ0dAE1Ywo5ZY5fto44l0klD
5U0URj7jXF3RweFjL9osBm0pvv9TyFkSIjkKPzgi8Kll/1Ws/D/Sjd4B9UckBFjX
DeSXNepy7Z4P9l/YuWX9CKn43VHxQLXHh+vv76n8CO4HFGhHVbdIytSGK4B99Afk
rU2waG/2R44HOsy21c6Ht2C13YzCIOgVAyEv6E5eBnjMRI6B03NBXRtJVUZw0yjj
PwqipEncatEAviKa7ScOjRvs5jP/R4qWPmTBI/ULh7oiPOzCrqgLeJnOrYpIL77t
wgm6mFGWCLOJFe2/sUmFI2hB3Hnk6PbfL1byFzqT5Kz0Nc+AGDRKitKDu92xlPRW
k8AQ+2wIHY7l2yKnLJ5TFSWQi3AZ0C3zhxRPa2cJ70pB/bBnw/HRC+L1SM3+YFWZ
pbiywR5gY86n8sCm88l6NZ7CEtNkpkgDjBcHZLX5ioQITl0gLnhkOWg5Fipa3xDu
YOhlBubOkR1hRAgTV2L3ivGKZ1e3hrWJxi3ZVwmpSWOLxBcD6C1HA+BpFneI7h4u
G4UzwkdwND+fYpRJRAaRd3rei+SNSFtEq+G/cPHapkfcmnJhjaD61viHtM9yJGuh
QQjALpo3C20etZ5e11i6ghgLrR07VuPfMExmhLiPP1Df5SftoQdICwi+lb5UerI8
NGYEHZ2k/g5tFRiCmmuc3gKS+3NlmDHaDiHOa0T7yyNWneDkq956skEO8ks11dBq
Jzz3R0+tdMRUSzPQpsdesAr4safY66eDaZ0cZmgIrF6C/ZdDU/whX8TWH5dD+waR
03SGATkaEs2D+gqXKpv3tZb2G2JiQmJVPIrxPYAyAiGvpaNuZQeiCjipnaoMmfgk
qXAMsjMeJCZm4ZDVGntXPq8vvWcoQNxFNMeujEsDFc5dNXglOZc0/yCE2mdArTEb
ABCM9a5kafM4GebmDPKYx9Cj47Qqp2Yn/fhv1hrOir6/pjP+73fkk+svfzmmzmBj
cMUcs0PYHjZy5zjzywLFyFocKoZPXXLKrgm+Ueo4ei7qvvkan/9C1S9FaMxqoJsE
Fjmnt6TXn2BC6pqNyamIU6TQLNGPxzf0g+IIYW6F3b/z+cg9nhw0LLMc069u28fp
GU2qLxyx0kLZxRaXagu3b4xprdZv5qMnHK30UsXWN9969QCr3y31r1F5qiZrlaku
+AHBhlDe5jtBdny/BbuuyVnClCccSxLHyEEoTytMQxS9c05pMBDD1A4ngqDXTYkS
yBov4DAHghZCscuOPbYHd3q5Fz6JKPax/TpBLJvQu5o2StKS0J+tAzK1IpPPfVzT
Vg2NcYNO+tPjGcqS3F7z6iVgELI78SLBZFy4vQ03xL5QV6ep1rxR4L3IVa7Mqt0X
IUOZNuPgPXk8dz539QhNI1TyKtXpztBccDs4NtqcxQj8mJ0YGvQnwDGRswjQNtr0
a/RW/J6jGBOjtGY93HeRWlh4mz0XuDzPh0LT17gE66fCPV3TNVC5vDSUxaOqD/OC
nJOjseBEIFxc456yGiXZEQqKcfqKeQSW5MWQNqklIpW7A9y1SY+eJfrL/qyinCBP
m5jUIP+PShRzVIw1TriDB+M+mJ4ZHap+6xV30lhZMh83NHFqE8L6T8lC1DBW318r
zgB5MDEJ+qzO+vutBQh8Y1qTNPbQ6OVCYC1EJiqWnOheSfDnahFz+GkpbPlLpVy/
GBnHVnGAZfKVnhNT+Br+FkZMA/20j88XE9LEKVk2qWH7aM/Yg0bP2JCP5p266Ju6
TmHBr+q2xi+Aib9U8zufuLO5eNl7gi4fJFRDY0Ma4uoJ+SGHRE8MNigyfvXSiLEL
/yVCnkXJRcGxrYjYsrZqVgD9dHVaC/Q0pi0ZUWz9qOahM4LrnjrlbDdzb9NwCgoJ
sigilh2YyqhBGV7TzYCEE7CtAhPFNS86t+4t9hwcoupeLP2sit+Q0YlGCIqxbYNy
6mOCjdJnxwG9KQBj0zCdSbU+GToCIz6AKOBUdSVLJwaOsUhJkOACbzE3ocd/dhnw
Zu8zdCTpxzocppI+6ZE0d6prwkanc0AKaSsw3FWQ0UU93p3k1EtgB8imbTHiQuQF
4E8U00jxD5REZcPs8r/uWVJDyaa4hxtygHvWcjXI/wnPBWpGTAa71oOzaAm2nb6r
O2aiYam0udLmBDMYTk9Shacg7ETrMI4M8+JMPtyABwBWs5r/chAglfrZHatEwv4X
FSD5tCCMwD6j6E5eRGKvNHU611TCUbXij/QdprhyNQN5NmcApZC0sty0UuUYJ+bf
kUu1nDJPH27VBWr5iczijeg5V3MTkLT5prXJDdG6CYXtEt4wpiHoiqDOwVB4/QGg
R6DsoIiOLVMKDiWzs8swVXA+d+jqn2UaRqAZJd+SaF2F5Yo2XNE0kqUIuPsKvbWp
yiZDA+SfJeH0WrRlEPujlCWIpbWvfCbgPQONs20KFnVhGVYPTMR9kDVZ7J4er6YX
cvWYRuJHmHr55DzvUktqEzEbmbzc8DvXHnC3tDsJuwBexN0I26apwLq6jItGgGNY
uJGR7d2d30THBJhrbnJrZVQLhq9xOK0Qx0ijuaXbp1v8DMRHnsoDoL/0wzJ8don8
2H328BffZOejXm3aFyce2ap5+KFy34fvrwVPPqjnPhCIE0/0tvXTw+Gx7/rU9zGg
1sQgy8b5+pJrO9QFDQeC0dJEplIpK74iXtEZVqteUPKldHGpsNwFo7Mb63pXRIUT
G7IZqdxQMQjxB5D55fsL0AqwSjYnr6FBd+UMxOnukxAPc9Z7ohyHRE7S4UKyShgu
HISkmLGgUdJJkluN8XhBNUZpyO94m7NB35LxtKLfo2PXdDQrh3MntqVTKeEnikoH
5Z3e81GucZKE2d6Zks7IuQraK3lbhINJfmSr1+2d9HMxbaz9lnA0E/2HE/O82BoD
D8K/PZ3Xz+o66P2DygWE7oa8T8v70aWCrPAbWC+63JkK4cKRU2m7BqNepTjx7Daq
ZrYYZg4TqFzsxaEy6Bky6SKr/kkNMgSQWdoGBicrNeOG65DHlZb4GL0X1+mKe0AE
UgJXBvwpt4HsSzqzUGsJN3siDUZKmRDUtzdpn6wd4Syr5HU3Gjg/131Xu8L04X/F
nhigl5DELDP5MkLG/RmcPA3SCdC57ng18HqbPEL5Ui8GxU/hwXlbathRx4BeuRzG
/2C5qPsEtYyT0kqXRmDGNzUT64MXeB7q+2gIlMMBVxZSn+zbfuhds8d0X37iJDIr
9LRGxhVXFRcB2bik7vl67CaS0mALTOqMgP+qn2FuPwBbz+7KVeEsRiZZq+RgwFtt
PK0TDyXifpLQU5sMR4kbi2R7IKYfiJ+C8VdhUarLP2rE2NBJcWNCdOFa2c+hwtR8
A1sA2NDSrrRQDee6W+EKBc5xkL+jz2DW9mvodk3FVZf5n76G8iVxxHk7fwjNrScW
8qZ80rjjpvTuOIu+hq8kuH6vgaDKadv6esY+6nCPU0NPXogh9qKGiL36rPOsLtLT
wwXILvVeUVaeYNJ4b3pxlVUXcieBM/gL88Z1P619qqqLe+zh28Lm0PR3E2IJGaCl
X348foCK7Tk/aEtlRGCLQfNlVzSjYjMKKSnBSB8jZA2vx0c+/zvaSsYah/o8VWAd
2hmf7MCwPTiItalDEdNzfKUAcTdUTe3/p69Ti70qZ0lskya4MBsHuqPSHF+IxeR2
jNKjhV/rXO3wt7VtCzfNK8FN4GdccS/TovGngpdIz3HGaC0wrS6+IlvMIby8ZbbA
2Mr78NUDF75OWsfiZdkn0ibqkwA9W4yjdRuZYviDklMkigKh1DcfKjkXXWfvs3Xy
sRuZCGVaDh8uQw8y4r/Y3HV59gkmLoknfXRDY8tYqzAfN7WJrk+aXM3TcxopR67b
g+gthud9ZwSa+dglUxg+UDZCE5QV7yS/0uaZ3L6yEtZ8FL6GCQCnwnAUcRitkIts
QBlnVzrCgWqglEGd9wSiMk5XFSFDTgWitGa3MJEhgoyfmtFm2EVM+Cfax3fOkky3
thRpVT3UoB024ndEXkop/Qm870L28Tn+7OHedqUCXyu/4avcKLco8JLKcUQAMNQC
m+8O9Ep/7P9R6u/5tyrn3Hg1qBxNoqDvXc7FJ9rOPBpRUCLN17gaJ+hvqzfwcL5z
lgCnWDhuGbx/r0IDLemoXAQSMpx/oYlkkw0hI7QXuB/aCDCeHY6zro9FL3JjLspq
yeMSujdimxmKR9jdj1VwzJdB/anNnvgAdUzwrLxHNk7S3WOBGiAnzKSQgmUliUij
0cOW4ROT8M9jw+Qpk9tryd+v0tlVrKDZhsNSvnAbtHfd59pC+3WF4HLA2rkU072C
yWGoxMqFBIagbquoJJ0CPobPNAg/jCUgW0cDV2oSqE1CLHQDp1ZnOby2VU1nupBG
0qXh2ZXcySVL5oKAkmBGa3l9WveT+M8XbliwsfGYbMDrWOl9Gh+7VpGZNRKEmSLC
E9qT393ZCDWJyFOC3MFuw2C4/F1sCdElhDT9m3wKC+O9KFLrEIuZpT7bIPLVUaq1
Vi/rlzV2qFjkWHxj1tqCCdGKEKftTPO4WpcvPwLw3xd/GT2VAcV+9udzhab/zLFG
D+b3y5WDc/noNwEYbOvgeiiqZhSFZ1MyZyoCyHAI8/qsJ4CqsSPflB8wncJKcB0P
IGljKhdOw+bCBeG35ti/g++TNjDuBaarRChsHZ4HskKXFwO3Go3je4JkWXZb0smI
U8o0OA8iazbvhPzTKamfU6bsl9NgbcIehv7ET+7qYBqTTh+TO15T6DlzM1Se7b7W
HrHM7iqDsGs3ex86pfXvZDHEi3yjCAyetVIE88/04FW/9gZq32LWavZx+BzKHfNu
7swSZybJUWJJ9NkGNgg7pyL30uW8FrjvcA8AGGd7O6PFWTlVDh+jfT7lgdaIpqyo
8fqS+AiIzCwBBKhjzJ+R6ZEubREHczhzdVq9ZBC998CQtrg5I3ZRLFq+d6w48O52
ySkc1HjvpQKbNzEP9IyRa7JATMhNRcA1mg7tIQIrvw/xxT4uck0xc1MeAEVITYFO
1/FBYVL3BqX6cfyQa9NEkdbn3KP2lBRXCY+xncpNbSr6ZxPhFLKUxa5tsiY9cmca
zy3MY+xIxjQP87Mju4N6uIVqjRWkfc64AAinCoU7pLGZSgs6XZ8mU6ZuyOQYgsOu
9XUhzm2ByoNseGeHg0QfemIBxLxT/TDvXV9awTLTsWbRX3xdAzimtMds7tlJS6g1
isOZuf8ki+T19sr0gktZzTJlFNtSQ+cuGpDtTb5nUoGJN+vB3BcW3uVwgo13bkNI
EujrTHNVc4vHdBkdCN0hi/5nuKBlF11ex7BwrU0cgYLSvHg/i4vavgK56h2ifyis
N3T6vq/mybm0jig75Iu0wAkMCqMToTSOmGFJIujHs4AVokE9LotHRYfilDA7JFVk
f/Cp7c7n5bJe47yezYGcNeVP50xh0DTQ3PMIz+tsikumzvdHIkLPiJOuuHAW5AWg
oBhn1o/rOuToAya2X5sUXQUQUf0drjJXvnsCiCtRE+k2mkBm5uD9J6Z4knm03Wn5
XQ/meTu7nEMp/lvbCcz8DMfiRnNPFa0D4n0VD3sJs7LEe4CJSTVj1a9JE55z66j3
X59Z4XPhQ2fHErh+B65emwfR7ldtkdojJiaiILOqDW3tJPHsmJBcLyIhbdeFgD5c
eRcVbM6nQ35jQz7g/U1lJuXGSqxfGhKtjZ+kXsqVdnKyUcqmrC6gZeLtxhssVPeC
HPrHJCfuwrwj94xWqOKkVrjY4MBSfB4nE23aZia3oAGRiWQ+OUq3LNKjgiPlB/Th
KKpeO/N2I7jnCtlN3ihqoYIb197Kj2ZYrpMd7xGzXX/vMTLLwMOaJMDQYXR54j/6
uV28kZ/FAKcs9RwuaBHZX3JHS5a9fMkqAapK8t9XeiThmSpV2Je/lCqG6FXWr/2T
r8zFNCsOwm5EdqQXt0Qn0JLqiYPel7g9G72BTaDqQnBqfE3f2au7sgWfIFFG0lq7
8YbPAK3Z9U24mlWXhMe3XAyO7T/zDWGmrhb9APZIAdqk2omuD63p0GPubWGdTgGr
yZvq9LZNoEb5TAPwD/+mEoR4ImFj5ehDGOmQ7y79muM3M7P8DsGl5KSc7lW/6sSm
rSO93JQbEoG4xKpU00eV2G65yBvcaznaccPsdVb8QXWeWirm6nG4Un+9Ub1vcUCC
tme3gcTlYoC06vucrraALPb30TZmJiTTIBQSsW9MjgevfsLDdi645cP1NXslKu/g
aRl0YeOQZvvUCs5vb+YEC5wVxnAsKI083shVFpG+c12fhnKix+wfS2c3cC7//k6z
i520k+SaekqyFGXmChlde+DMJ8HLSeaBJsvgit0/mWvww+2NnMUWnBJTTpqAnVqy
lYfXIOkXbZ8ZAjT4WZLCmspc4bAPe+MW6jMVfoSK/zOCXAGbA5bp1guzn5TtHhWJ
4/S6091jruyfPHDJyStbNh/fh2Z1j26tcsGxdk6lhoBApuzAkdHjge23ZsZ8myKQ
IJXg3sCC4/gKMocVCQfMRSIJbRfF+JXXATa+3WV6v7MaDgvf2S2hcPVoHxCv85Z2
zKocI1OST9EKLmbBeBINA4e+sBxOBbdmFvG8LMt639bl0OQIQcfP/pHGls6PPmvI
GoP9cUnmq4OBqLqI0N+5HbktZyZd59d132lG9Gba3F4hc+vOY4J05DKFxI1MjNzE
uel5S0Xwrc7w0uyTu3O6j6VPHW1EGfAP3gDSE8XeBpdey8wSTrY6/XSB7W5yET6P
U5bms7ibOvrZ3eblhjEnPUx3WHe30RiPBCLmeZB5kMvRdkFIkri4TqoNzsK4ui3f
Be1GEPjCINS7KYapDEAwUhjYsRtevLa/bmTW4cf7KyOHUM9OtcqHSlOI4NwNGjrL
XFWNehBlv/03CeRos7mDYpmeQw52XYT9eWgnlZy3vqjdCJbb/f9R/On/rFaM87t+
/3x0uCc0b8MBSjm0b4+Q+NmpRJ1rJzb1lN/8gkUW7xhDxFidMBD2YGhrvvu5JikJ
YGn6e7H37Yc7zcgKmCeiUSDtYXtl7HtkgstqHNnKECfGvT09d++DXqyx2qL2qLhj
lqTKFKrUmZLN7/b48SWAakVllCFhmd3qxErwn88sS80NE845n30bynpoM75tH585
u5bpeWGVwTI2jbDJSJQNGPXuzO7U/NTmlCezGYSncvA2bIaa0pjBXzR4LMXTZPZl
ktYTaifJN09tVb1au5rKgyRSunUe07eRuRwsfSnIwVUIGPJxc3k982s1Makme4rA
Jyv/QmOYmM3s6TM8g8WMm3FsmePo7y6kK5MPdAkJvhkXy2BUl7Lig32qZW3n9bZp
LqA4n//DWkbz0/04AuYc9MJQCTtokGNYLaQ9h0j90FWtfH7NzvLoiCGw45S8fjIs
4QTDyoLJTIf+pH8JbU5zOerTwJ94EoWNqcLHunHUY4uRtjEFZeI0r1mYs3MH6gsU
DB7gZIanRQj42T69xTGqGkYBduD9WcNuP8UlH8bbTSpyyHQ70v0ujSah/hvdDUj8
RM8CPWDSJF8xvf0t64cqbiuQcg25e4V00Q2l+ExwjYKT489pX+QE6RhHh1z4MFJJ
mmwh4WoYiZECvjT2pBhGchAGXwRgGksSHnYJpuUhYmpBbjEOu5kiO/ygsnGSAhq2
OKNhSja3WN1fvR0SZpD3vcTR3cmnRjGMmE0weQNBzxXCl6b7kYXdzeNbKz32F8Z8
sz/cS3O1svjVepPzuqEi2kZzJ9ThH5dW307gbZdBhralhhwtXJPhDEvQ1PA8NJgH
Qx+0n882Q32i8KTa+r6OLRi0O5JSGVq4CV7H0pXqjXv66/bsDqWzgBBIg+vEL1cF
3DKDvrbih6VfUs25mfhTR5ndjs2YRrn96ls2mGtTRxZ7EH0C0+sKMX07EghCh60J
MSD5CEP3YjhYbkMLaYSXMYESUmWoFBCYC5lwDERC8dxoWpZhyk5842a42HLYcFSY
JSywdoa/pKWtQRX8BiZIevrC7Rw7avOxUgFmOZkvuflMh0xxHr7nV2kfqZ5dT+4i
Y4Y94Kt+OdP1O5A0B8YAiXEWyfexCbYcaD1WNsJZ3eplo+82+qtf4CN7efUbrULP
iIMI3AH8qGDKZCex8iG0dimsUbXkD4aO8/n+AxrIc4bbBAOGeJg+sFVTlgboNpzj
NQGmctICSBu50wypne0SNEx6eXMtP5CyRaYtzJePBfRkNungnqraA9QOI7aoJFF3
dCbg4PMD2Nkvris4UzjBgv3Z13LkHdK+aNPNcKefD2jD07FK7Pf2p4o6IQndmNjx
jDtOm/4JfcN84/Q2UxBv9+/rJJLwQDmypTWf5/T9F5grFsOlR/NNgSWjmrAc7N4P
XD75eNz+sWWXQofu3t+lgFwpBf4X1vtQArjOFXEkaEpixgugzg49HjS9X5RjAl/b
3H79h6S+PYO8QvSAq6PZw+czADu9cN70jQqGxgnFiNrlBSjMNKeiLsaCqoHGeOiy
5XzxBunXnOyy2MVaGFWMYiTRQ5j9E4neYjYf3/pdCnoxggIQpzhFQU0Tgr+GnTDD
3/pkqzl9h7DqiYViyOuq+6JcZ5sT3a97aLx/raZ0FzfVnKOl14kwL1cJaO0oXV8l
plMh7gJIzIl9w+yBM2ZqULL3C/pRr3adPNsf9PMaRCHzp5NJekxrU5TByY2XoHe2
wxHgHSLyYhl1/EeNs/WePet3uhwv9ZhaJFLafQqbGDIvG/YfZecVWlQ7e5ldMAxo
NeFU4M3FxkT5EaIN2iM9OmUA1VmJQPLOvIEsjUVWvDICrTLnxmipyQlUxa1x9k2x
FgChycFoRe7miN9at4amRU4FimK06QOCRZWOuhZe4ksj1IEchBVT5zrCsaTSzywV
nZWE+/Qb5lFCmj6hgbBHc98Cqw7sypKwDBa8ZKHqzAdNALUHVzikWiOD91iWRav1
gF6vKgxLzTEw87iWeQYj9pynKv0ytm6oWXoM1/l/clotF+C2WMWqgMML3PjWKuq9
uaP0udBO10LU4cUPNz/vs5yWB0JBmMonwo+1H0PTRePK6c8oI11bOtU5lG7mE8Fh
z/ETltxNO5yqAGcBXv2uXRBoceMwgWHbScmdAqfH5CKWJjtmhdqoNzP+Dz/mUo4W
Fyonz94Hy1szwYLbLBoK+uZnimDMHX56uN9qfSyMas+/7rNwTCPie9t+t87zwgv8
Xr64DSYqIN2PAoCCLPb+kES/baP3KrmgukYKhBRwJOVX7SBZtxWbAF43MPVAPszh
SpdUycfDZQJhDjYpJTSAy2j2coLQhIyw3auPYDqHYFwyCrbhY9WKL2LtEgR6SIz6
NFjnLVcJk9Rbu7vI05WxJeWzi6wMIEHaB/ey+UO9rljEA9TvV8z8BwyQE+zCnuds
9LG+ti8X3FydAMYCNF1/eU4zUOmqAB/7ANc04tsdkJulHIvBG15Ll6nOaWenO7i+
CV9JPME27vpbRoBu5yt3gK1ExF7ccXncdxetBMlbOcUW3MOF7/U4MVihXfqBnTAC
cqTgTG9yIx5GOhm6MQQPTbBIoCjQmhDEluPeusLr2Rsg5HorT528Gso2JYiIORlZ
QrZFBkYfm8g5cAKA/LXyEa/kpNlGWOJ68Wfs7RmKC25lgerLUt7Ze9H0DoonlMvg
9myZgcySt93Yzoa942wXwMjPg1Htst6oli7lWuUL4/DjDjEDhwQX0Btw+2WjNXKU
gHQGWAk2fXOzcCtbA4FmubNj89S00/D2RQKMVxHp40aMmsGxVBCVOQj6NyPupaQW
NuyYXPvGS4teesUCjRoV2t5IOFFJWnlfwx2nfvZ7td62O/nZlVTXzBU9GXYijW9e
8JRhRJMkrD/WFuEfSsAjlzhkvpKfHrxVVrhiXUiq3S4UGCftFb9zN1yLd0c2qJMX
7OqOP7iiRgplyLTCi9lQymioPpySoagXdS3cvM/6XXB3A19uiz/LJJ4vh2WpKO8D
AM/+Jw+7j3/NmGGCpyAfVidkCnmMhg/3DsG3PTn4IRaXQuRpaz/s70QwSGjwhves
dBU+W76yXTHfua/oFKABEoSt1rqayzbNiFC1t6tFx3bIXby1vOM4YKIxacZyiDSI
borfZlE6QA0h7g7VmQCa704jxU28uTTuHkzQGVGJRc038a4CMt8Agij8Nn4PlKyM
8bycI7nzM+MTkUN440mvuZ9X6R+b09u8odEfjMYL+JcnUlfAxf1Eu6fX2q5cvOog
Ftk4FMA3amgtQbcRZwokCMjdp+E2x9hHW7UyP7aB0lSiOUjjnABt12gPRzWgjtFF
QNciPZz3CLRlWrJWz29ty7OiU26bxtT1fnUwv9o9zIZCKnLG2Ogi912kwuqd9bcq
0eAPJ7RWd4H3R6BpTOPAFZ9VDMKmMcAXLTV8GmEV2eSIV3tEeUq+ltiZJmkLHOm5
eHWUK7EPGNd3mk6pFhStjlYDELGZ37MOLo08LBlEbzEWfgaJkI9dc3JyqISJzFjt
IeYZhmqWiiVqd+C+PWKCr8iTknZC/FGfO439YwDip3SGTgB83r8J6sjAHmi8YUqt
IaxzsHenwvuR5xTbMrt6Km7yjNF4i9YMU6jN/KtJrfRk3R/BNGc3q0KcjdbeqrR1
UVSh8PEhbUfOtgjiTmbRew5q42jYhLC7ykKKAUuxedWJiDtOpEyoFiwWle5OcRpK
cwusg2QONWXuQI6TrjAYZnpPsavvJqRsqixwEyswp5daeawtP5UX2ZbwBDjchqy9
jO8Fp9EX/pdz+4vfgpW86CdyTGq/zUuPV06M4GwHXaDjiF/1sXPnom1kjCD0EZFF
jeNarG2NgqCXjjMR/z+EdOrPZPND014SgBxMbeHQGkKw4Wg4LabUsIiUTzveb4Ir
yAWxzi+npAP64RSJGGWP5Ecw4He4PVxUTyHpyGO3kTFIn6sXldEVuVHNj/OjXHjT
g92ENPOV97H8CXBdacZUDzZjwaHH/KzF+CSyo3xyKJb4DLHFBoeC18mPhVM++NQR
Dy6ClsWrV5Qo4cH+faLVxjYSBovZGFPI9XlGBpzD0f0k49HCbhoOFXpE4lorDa7N
xgzpwbt7+Tg6zCK32cFcF2FaA/FCGpkIxXdXGe4i8Ga0DLw7ktp500n5ZSuhKjM6
6PwHD+vjZLV9GkkFjvHEt1Q5GGjikdA8u48RSKv6PFP/+hYsgCWJJFQQP9GiAuI5
8PZbh49CcrB23Qr5s8ATbhlIYH51Hqob4+6ZxCcbBy3gHvgzsLcOcu/8ofE9SbtN
8bM/jBpR7D07wdustDQ5r4k/Xhpw0L0l5TYwpRVdGuU4uh1n/lxOVKA/sD4Ub5uw
Ycx9gk+VTyNB6rmsYpjr+a/bCVENS6hLtdkdENOj9J5+yGF7IhsCN3U5kmsBg+5c
cq8oFaNMXHzNdXyixsst4hcqgDuaIra5iocbGBZScXqr3uomD4mdsfauLM4TpIU8
WnnQZP28ZmxEk3Jgdr4C7wyMFuCaSt7BCR9zZ23QeTPatQzXKL3HEmCGiy3apTcI
0X5pOfrD40C6vjcyZaqWTDQ/EtkzjpFZvkhKMZki19fgZoJDrM9QunxV8WJ4s0Ck
rlVn+/ACL7CB1hp9lg8EZ+C2K2y311vm9Nse2ldr48xr4uOEZ8GtCCHbyShoc5Gr
+0/BuvAM1jgyVBo4jiYolLOeNJkh6Q8L6usacbsVv5B3Z2qIMAUUs3LHeS8p7f/r
BeM/2SBJxhbdCKnnmNzvHUBWQ33QPCyU8k6lUfGxvZOOZHx9R/m2lvOwG1DxvKFi
iJL5NsABvmii2mTTpkWMFUCRGf7ZZqveGg9rzC4YnUdo1SCdhobpHyVv2wIj16DN
fBUvbITz4goIRTYUmL7A4ljQkhkkJPpNJgZO13IDW7k/oZF1ThYkkzznCcfwEm/t
2YBdcPH5/FEte4ZSemA0S6bCBy/2ISk/NCkacA+ZyQOD0lylF7oVCAMXp87MxtlS
jsQ4G6pfAIplf7QVbiPb3CP1e4Q8zYr/k5f5t1T5X+6TH4+L0ZcnOV0wRDyCdWod
Ssw4XrrWtC05oJQLq3lLA+s2Sdmrsm7FD7Jwl8zXTqTKXfo0hETFJ5UDNacTlpaS
yAA2i3BXhxUsXbFyS4y/HO8PEmmfMAw4H3SKOXLueN7QsKx8+WGcDp8jBOl6ctyp
Qvg/ayD+nrzuQuYewf1uVMhKwHYWbMchCz5/XfaEx6d1qQCdQ5TSrXtc+x5WXGBh
aqGWETwahzeHqbZ2o6ekwfaY9GWxmuJ70emyO90c2et/t7rey2WI/DS6amOlXnah
oldFlu1n52f85KZ/d3ICkVLQHKqPfnQ815dB1uFMsSHOEAuTLgCjds1YQD1vqpKc
MOwHFNCLwJf/pKgqNBS5hy2VBAgONaN5TKwFbkVsWFA4XUx4rkK3tVyty4HQbfuq
EQ/s4yXvXmVKMHjfHmFy6WGD6dkmt2Tvi7RCwHigbzq8DXRVLBkSmVTRhXa+zLMe
OS9kJSll35ZKrJgDJPVS29lcDr413tLhTNdHn4YQU/izMNYGv1DP8ZQ0KzkXaQSB
Hs2XgBAGdaYU8M+vjISdWYDj9S/fz/ukQEaoWQBw/doCPHFO8IFsOorGRZCyWMoP
RBVHAP8K5/xXbNmXZwUv2qqaU91nfywhJcVhBV9VImhiCthiFQlmaw42hR90KK8o
nwehfFrNhYgLx9zU/QsSVH1kw4CWWqxqjAceNHebxw3WUeQmT2MN2ILmTApqw7An
plbImpxSs4nG+AtdzNGJl60FdekTIVkFEU/mEX2AG4kEM0Pc6+tGlIRLh7FlH7PQ
NEOUhkCAbv7kUI+Gy+Z+r763fAQM29eGL8geisMDkOw1MmEL8pDjqhbZiaaErttq
KP/H4m/stNExXagQewhZNrUzdkpIBgeT4PEfC9BPkx9ZU+nM4w4mXx0Qy4tTIU2T
Z2xqiw+TEN67L7LvBuzOcrs0ZuiXePppNGLR7PtpbSQcgVRdAHk2O7Uf9tDCwL39
vjJmdEh82H5tbLJUScr7tLCt6If4EVOwd/CM/6/JMFC5Jt6sxsum0HiuCNeyFJNX
35nSWkaQJNYLRMuwKxJ8mb8diZVtL6UbMn6jwAc2N3K/0yhCnPi5m8Y5dKW25Qfn
3POoEM72JsY1Xf2RsTo74uTV79VfUVeOFOJh/cEci9Qqr424a2ZFMfY2rVwibH/f
dqUyX9W+Inc55vaiUP975WDzdwer2/Ye9rUi/+gt85UL/CsGN9UCCqrkksulQlBf
lXQJ+/BfBBYnffM1k3hT262U1iuGOdaLYZC71jXwA4I+E6QgfWTegNLCi9DVyrrC
qq8CEDE7lGg45/yJGs2iJHGeZDe17QCKwIC8bHt6N5P4oNaWBIaL96JwsNGgXXdt
Zc+b/WX5IPoZwivGUllepKlCvrqfHuzWUR48zbr7gGIak7fDC0kJlQkZocy5mDwL
6u20L0MeCjyKGfnvU0dDmeyLRBMAuYHoGCg7RLLZEtSFxC8D2sBj1NEUmczvkJAv
jsTfGNu3V2MbA4P9it6Gpe2UheFo/+lYWmhsZk/4VsWAWKXLLrImcF564rBv4gFy
/n35Knkpx+a8UdqTXw5EUfCPj3dKTrPRJu9nZaGrnR7GBlkDAz7KNw3u1ZZtwOc4
zZn50caYTMNaNqhTeKRhgo+X3gegiuHoUvPOf8ejJEGpoPEd/kpnEjvTbgsTMK16
A3sAXZSJgRzoaYRS5XB3Knjr8AyXQwghDDSlOrGeBK3jvnii6aimIMtMaopHE1ai
RnQ7LD7A6rwkj1rb8X8Tdr7ygsiXJEkdX60rxmPpPvQipnWOoNfkdv2NQ0/SyPXG
n5J1y6EPaHEx4QxsOrHSvLbQ9TVDQrmpdt2LgbW1DvNasxgoyvyiLfT/OLNE4Fsq
0SuD67Y/J1V2osqIXqTu5kckJxxbCrZUXw/H5qwW10e8rFyPH0a18lAUPV7cJWh7
o1HZGut6NYrDwajg4XA/iCKfGeDYRFv7ZseqNQouhBYJspbfki1ztm6vl1Jibytx
dzzy0QSAU02bVDBhOBGfzhItJFiRFzJT/M65XyIPhE+1bhYIwqT5R2vtUwunvyL0
FzZGP1bz5DFoy3qiv68g93lzhV9fC/nUDijYWlwhaKP4oiHGtoiPUM6+4Gbor6+N
QiLsvt9OQYVSX0JAw7+aoWPIqDdZrLqtwYKy3DUJASMYahFsNfJiPJIpyksR2eY4
kcZh4JFHyEDWMlWZkPVvZlSUw5RQc1tnCwMA+J/bM8W0nDVgxYqiqGCWoYw+JLZI
+I2QuR8LtWi9FAZbR0zN4HN200vI0SALpiavuvkLajB+rmN6Lu1HV0KsEwZAbG7B
1ZNPA0732ZocGpmhu0h88LNTCZ8hsJeNHmcmwKwRJi5jG7dg1RdCgQaMwJYqSo6r
XfKu2esYHQx2nvY9xOLcRkyW5l21Lw0E1Jsnzia1aCx+MtCFA1MbdThO0IesbOa7
Cjf+fqWlQzcuJCfVCpHWTJ9F/BBf6672g93kCI0DxZ3kZC9kMAhouUBU2/TO59Pj
wduNU9c4NuUZesZbIPBWhljx9qBzx/oxVyO2FWeEH8Gk0hc0NgYubwAbADj/y7Wf
qam1FqEiaqhT7ICtvhU+SLLLDMG30Hg0iiEq0jeV2nVilTG4fAUvd6Dh2GekgzLB
OsNPw5VuXp0e93ZA0n2jOgBUL8kc0P4z/1+nTkcYe5NmuWwZhqmTdFcnjBin2/Q5
+mi2TwvlPQZPo6r4CUBai22Q+9dLZmN0B5M+t6gFFd223TKaFf+rJ1IUYZpA6Yix
hKMJvz5TF6/mFe+joC/hxrZOgEaOJx83XxDsyWLNJ9o7r4p9pGcYpe5xJrSip6Xx
I8IWxaG+cQxT8a92SMpc+jKlCMBZQs1wXZuT+V8KhJaxpO/Gvvp6Ww0FTHJsdsbB
iozy11t1bSG5zVf8zw4vzq4WgcisghIB/KMtPaP5ehp7+0t5x0wtcDso3Fw5Nbmc
yqPIIBL2+mxdtP5FQ5WZHiWXAnJCs3xKtLMWYtdW0nlOFARmQrN162R/7OMRc+hM
Ngv2wrzYniwu/0hrEJNlss9gWA+fijUNU6/8q3V/ZznU5ZnA6TLr679Mav4rWb8q
jXAwLEopVTqhw0vvgt+62pRzf+hmWJtT1bxqG1M9PY0x9WLLLHreri49u2uahcOT
HCaITCqZX3YNIDPTUiUsYrYIBjIwCu4cvulNUn1ryVtXA0TQcIGB/u9Bmlw3O2eN
v8B0koBzB8zKBEVrDq2OLayllP/uapSpDmhBGPZ7slOdKJxuylmcDuzNWF4wjhVD
Zit9yuYTZ/J1T1Z2XBjBRHVIFRQoG0jkmsC1Ww0e7n7iMdcBg3KOdIGgDJjHgPAx
wgqtd/fCifdbIO+Ly5Im8D31QTlrcUxI+DAo+07JWjMBT9T6UzbdjLV+UNpxUWBw
akGlkcVQ/EAIuPPZ0+bD2FGe1LjqtItVc3/XmeKaIEnN1SOrrvapgY26+/YMyt4j
kokj7kRIhCMwkCASrH/3wCKRZSUe1rtwMQxNmXgtfY+XZXZ6Z0RTLSyFcZ9xpLNM
EyoOlV2eLSJl6gUK2T5wa/YI/6zYjyhXurDOHMa3K75x5ywcEaSoRTuZoZdK1puQ
Ctop8Kt0ZKftQWH7UevBt6q+94nBIFPChHndrwUFt1nWfPC4ZtOrtz3Q9A9sIJIA
NyNtth95qD2mCzmYKdvA62IjS5s2wW0y3EL/3ulOxNE0W+MtW5QlbYUyBZtixMbq
TTtFnYd/je197jDS4jtkdFE8IwywYDZWU96qQtTta7iBWpL2KHKrvhzlH1CkAS5h
O36d+ZiIObDs5S3Y+mOY011p6QYivyBbB0iLAQ7NIJe75wNgcKVk4gJXPuUIdPMe
hh5zQEvZzvRa8yPoBvurItahp9SHlvArtJFUphg0JXEMDU4qBCdIqkKyEiaHvmuJ
IV1I+7fhnJ/Lh7dGyhKy3s0HEa7ixe59g4T7MGpBd9HqcFezHxvBDVfFSUU+/92L
2YZZMDceSiedNP97v5Uxms+/FFYbhXA2Zo1Enffl/kXB4gj3p4tYTFi7BFZwgDPQ
7D/9T9QOuD8ugTnKzFIXcqLh5R6mh06DROw1htSckziJ30q9oe/bk/9FNum6lYjz
3BmC5qKxf1vDXA5KmMau2iInOfXz9deQ/uMHNy1BFmX30LVd3nEHvGMcfudDo5qu
F91KlMrczpL725+72lvEO0qTSereWcIBNcSH+zIRMTIlKzsXhg0Hg5yL3KIe60F+
ft1tu3EB/bXKtJgkZxytcj7c8JfIwV4FUHl15GE0E7oBsZKrPpaStUJPRE7CIYIo
86UeBnpdqIU9gvkk+uBvYnwciIBRV+dvrgYclt+lFjQxp0OwTnD5Wol0kjpdiQmf
yD0aZF2OnA/w0E+o5z6/xwKdScgJOjMmQ7FL4RcQwMLH5jKnfH1AawNdpmmploCb
RE73kk95KaO8ji1utuIoyiKnO/q/vf8HwKqI+mKPd43M9z93sE1LoxQq6He0Rr0a
KpbHwJ9bwrHhPIj4eZWDaFFCAWfM/g/mghwomwn09z3jeBkE8lvy5uzP90t1HQSu
jow2+A/NapfPzrcQNgjSSl/Z9tEDz/ShnOFVVHq6It3wMx66ye2imfPrQ/PiQiPs
6oGIho9zOsz9rCHcFwzvWNVf2a4qEG5KxUPldfBeY3kizyz0wGDckDhHNocLk9lc
l3YC+JDIg1aX9D5LY0+kNyxO256p9smQVN05Yj2l+Qf4bhhDMsGHEr0OK3mEOd1H
A0AJ2rUi1ygQW+HfZZiL6EJPO+os9TTbP27eOkmB3yoKB1N+2uwrvjdY1Z+VQVJE
w+rW9SsxKwzUnNJlj85A6UG0Q2/nOc4YmG804HcB8Ce2BHEfmsDJPSVOb2y9jkyA
U4xK9b++zmQe9zjAxffWI8iYhFtWlz5SihzvnT9nPYkyjAKzGwJk3qSksM3P3CH3
ldhKShZGRr2KbvsGslO8cXRMEBhPt0jl7xmZEOZtpd1Z9VKT+wjkV/lxSQospNve
2OJ2sBStgS0nX7Ga32xxwL91xlTorAEaFPiEQsUJbjotB2GakP2bevB2qlbXGTJ2
G2tCuQcYbyo1pM0+QaZBdJlJfSj3yZkdzxGyeypWGIdCimb7TSEWqW+HC1j1or/S
VcwCHxnFLuq25i4pgvx/idVqzNBOll7rdePBNU0c6TqhnNVgDutB+MZrN2gwoFip
JqqCIENbKzcRm/ljy9d4ugSph7ZoF0AibTE8wvjuSEGROd3reebvdv+cnjAwVqvK
BtHLnmmmrcHULpS1yRfT8JrppEHs5NggV79yX8MymUcu+EaT8LPXvoIfWYS7XIo0
94O5eIubnCg2qZtiPUsqb2bYc7RK4BlLvpX+2e7uY2KzzzImYIZ0IhcEVj0t/Qw9
10dQ6DRllG/4EhLwUNDn0vfDXJfr659j2SpaEnkAEXxbtu1wKS4BEvbBFeGAXPQN
zUEcdJFBwUdlScIRtvw0fxLmyegpLwWb06oNaDzbCp60f986sunUZqSOwfKMbESr
5AvOGgzkKpl0jgNfFQjCLPWwiWfaKKL9fZRYuz7OrrU66FjvF2keRYx6T0trESGl
aTnx8sKQI39nyVg2FFjB5A==
`pragma protect end_protected
