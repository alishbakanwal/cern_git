// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:02:08 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
jlsrkHednv4t4WFxr0iqGZ7bQkiFXSOlKWbrxPICa0rYCPVugtka6tTGI1o75Yz4
ftejT+nkkqEs2BbMW8rviAeSggDuHIVkX02lTaVezxKMdfLW26AHwE5XqzUMxgCk
Sv2zm3r9gKZ820nrL5Z9VLOldgKGiWLXNws3kVydLzc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 71104)
r1rAuMKBTMm5x57LC/ukqC0JiyoUUdV5sau5JPC+bL4Dwuh2kaLF0oKzptN0Tm3+
MQfv8c/HLHJm3X3Xl3PgRiADhd8URnZ6ptx4EJdiJigf76EMMKOR9XNbKqia1WsQ
8oGIpJQURSWElktpRYIVNZo20tN0wmbj6SlDCbBeChs4bCUHSdTxMdJsGKNN5SeP
8MtRtT+QUKHeRbT8F0PilKVfyoccN0rUEA467SZx9fuFrq7YHafAONnxRikt0oOJ
0rGf8DQFWKeEzI50iupgc4SJcUNHv2AXe+levy6hgbJqdZV4tBdxq3LqvWvs3plG
VK/+ECWMTIYbRo5FjmMY0c25U2iBDI+7SeCmUeGZCADgqJRUNPVYlV8gY1ZoBJK7
ek4QdigcyU0vdrDE9bYd58QsXLzzySJZeWfvHb7JtqN620ABYstd0TLrbc1HOjNT
Tzmhc8hB0DtSnjdS1wAu2DL8kCoPLxLGXvDn/fqKDm5QefvOQeZUt5yIpr/XnJtW
mF4VuOUPUP/qfUNFs1T4yhlRZ0CoHHtr06muFFkv01zfEw5iqXqRLiHCaUi34tDH
08Ohwja3SrIfD786e2aqsn5WUNmZepfjybTxMOyJYg+GWP13vYyIhyT52XFuVnPC
REghuCc6ic9MVHsXh903UwA+aVBfUQUQgmEMqdiamxnlmY/+NYofSWfI8ZW8Ts/y
PsMxzLzj+YKLb5yoge92bs62VMhaEYJOp4V0HPBO+cl5Kf945paEeOZ9THjepYnC
rr8i2TQaBzorCD7/QucVJqZ6Q13BLMiu/0LD8dwwcBri3yuzEr2zWv7Thschl0Ic
b6FFQPAfgQL6tPFmmrOsf3TAiQIgvdVLZjiZZrpJD35AS3ZtvzmlKh5Q1ORbJK8/
ULgAF43oPXWlCiB/SIy04w7YRAl/UZpnjA86z6IK+oai4fyONhSIcMDaFdDQpbE4
3XBJfviZcS7zC+3B1DXfz8pbLWozk6Ll1vUj1dzehGflaQ+Lm/qdFRYxSsy0I4Gx
5CJSkpscq/HB2W5biEny7R1dzOnVI2z25Ga+cVww7f7RX66iFHlc/Ue/XH4jZb2A
VtEvfcMbTEzTL965jWQbSQg7GvCpIUGXzH/fmqa7jatD954MX2QgVl3IK9L/uaTo
2fTrFZWpNvFvCiFbb+G/w9kMhgkutwXSlCoLlBXB5gteoc5WgfwnfVqZ2WUtk6Ml
PmPuXiAnG82x/P1yfyjb56hcjmfCMm6AlusDDytIb/Xde+BWiazJiad+jrtEd7pE
3DFWXYpL7IOJW6L1yUBKdptYeYThVvV8GChMPFp+ZwRhoj6YWDnu6WNjkocE4JDf
tTKOAnVgspeGGIAxqC6uwkvXpQqnd4lXD8A/GxduP4tT0x/KfjGW9YBFNhOb6OlK
Zv7P0hinz206zNltyxIEsbkouEdDYlZbI4Uz3XohPsDRvtjCmzg0IWPOt84dnUpI
Jb7agNiRTToC+uu/q5YlvJi+5Fyf8UeJjy2LX40qUs2Xxtn13qMPXERPAHLP8SAm
kszRQvwQLRFkk/MHGW1WcH5W34JgWi1DYrPNNZ0xNZnwXDFEDi4G4Y2Nn7SdR6t4
XxqM1XPRGBL/tIxpl2l4Ka5RUAMO1RT2pef1ObeFLvgBK7mwarMnfHW470VG9+a7
wmLFvUyqA6rB91r1eDJW4TdWHvsta/4FUt1thHqk8IzQmrQZXl1xegCgvzoWWPQd
CiE7iA6GbprSKaR7TDillzuHy/a00UsPcoAH/xcc5RXALU0MB2nFuw3qwmf8lRNI
F6rzga/My5UW1nQVNkkDAS1bcEi17YwOSue1Uvg9Xq2BEGeBLtI8UzLpFM3Lg/QS
OtDgVxjinwchYD/MzcfZiW7QEy7gUyDZqLlyI2sUCyIoezoPLrZj1uSgHykT9ssc
ZJS14UO+8l206JVnphcHdlo0YxyzVvmFKrhl+zEY4xkVxR8+k1xwoFEsunnM62xa
bM8JKqOQB1geY9sqo+NsPDag3JsG0OjmLw9v0bTayVlsO+tc48CEYr/GHmMgSy0/
DOlZSSS0bMJiJXsjYPOl76/jUAsvBOGdsK14jEDug60hJrz5ULdoNdHDZW99Kp7I
b3g2B/p/ynT/WYLTM0qNUKZ0d+9my/RJmOOp5QJnMz1YNRnSXBnZwzYAhFOMJ7DN
UV1Pun5fhK0hI1ob6R9IqHrwkNs2KbaWQfdTqMqfEGGZnXp6UGmcuHfc5pOYUWYl
RRX30RXOrmJADGQDGDxqxzArWMJtWyt5xe/OeCbXuhhfpvizYJxcqV1XN02oi9kN
37MidiuhRXKxyvWyO8pNEUjYGV0cOuQGuBHc/AOySRrNrpOcPzu8HgzX+OGQg661
oq/aEiAHhVDSnJzRpXsQ7G2pcBZ9heb+XH6h5cyZoUveYVhwp5hoeEKSq9yyOTzA
Jn3Cy18QQXGnoGpo05Y/p3pkfjCG+bHua6wZvD6HJnl8jiStX1r6mPTVSh5us1HT
arxtJDN9AUV4VtUgHenbELBnXBTDwj50U3N84XogiFdfXo77kSku/z71UHBvRydt
LZZjkbdt012drjg0ajfcdjBvI4foOwLXE1zrlAI5fLpXm8sFIrcPK5h/6rhL+voH
TAzN/XYfcoCR6rMmOgSG2+RmLiaRzW3yLosWFhYHj+ycZwWNtDLHJQbJ1nh1psYA
w2KLgjCaoWEmdI4YTrQcTeBkH47Pe7S714YLYUeYLseknq1jOsIgWu1xFRFAEZpX
1NhihNp18jBQvrNy88BsHpf/3tlZMrGIhVwB9TdIwfz4zZ6KezvCHiZ/550BIMLr
IkrwG62WjAexqWu8Nm3MvTi2pZc3u5SpqXOuUtaiqXPQNapALbkb/TcGsnPk/8nw
F35h+tqJ7YlK/F5eag5mYLK92GqTlmIZ2dztjdgbPMhz1ZwvZdKu8GwK8N8XZvFd
2mga7tz1LDE0Rj5MHzWGcOq2LRKRqiC25LLTc6WujMgsusSrL7QGFsXTiV7yXsON
3VXYEjcz8Erm9L9GjEbqIlFUb6olidfdpA1HeYC0WasLQyI9KdkFHX61eC/f8jmS
+KmB6QvW9P+DMDV1td4iIhxzsVCS4/mf6hpEQlX5/p3utmXHipPeG60m3CoJ4Zav
eHQUXKzs0zKBgFN7wKEEhQYpzfpAjmnj2VOs68JTexjOJSaNZSrvzhzkCQWLIKLU
vR4b6AzikKR8/FeZV902amInsyAiXKrGZv39iNeWZ6AUXG6qFm0assq9EZRKtGnB
2wEJxwn/EU/hlyKHgo5Dd/wSex8Nq1HZHHBrMVKTI5ts4ulJ6ELgUMXLU+byl8oI
ft+Y44gJAOmCUJXxHHrjuflMVSte50IKJoJy6L2uWd3k6EvNwyzq5vjRglotv+ND
V86BQGT7L7A66Dl02Jsk44M88kL6lY4yt7KMVd6OojSwevXYY8w190Jy956tw4JJ
PZ7mfQt+KhoG2JS5jWaYM0g+X9LYjSGrJDVyotyCuyFHEqV77Vs+DOVQqdE+ybw6
hC/KZfvxtN8puofKcB8u+Hb8VIKE7qeV8KOfJrazFMoAx1NqdMEhfl+QjchQAVYQ
GSFsDs0otBwyRbvzABxVpejRGv6n8SbqMRi2a0WgxwSZ3YtqNgHwGuyYlwQ0nfze
S/1IMdbDK4qTG2AbKmTSdtWow1QEa3O+J3WjwfUoX3Fl3EwBqzvBoIukSoSZBRaB
KsGo+rpgCocg2cuS3UzJh8zPQx/Av/S+v4uN/IkxsmLVOGGz/SK1IkR5nWSPWaOA
VwBQOSzIzsMUhABKutuSjsOet+VTRvhyMFsTjJ3CVGK7bj0abZ3PCjuJ2oMLVAx2
hqTBuNlb6cK+6BUCT5OgzGXqgKbGaKSKXUaWRx5u1tyJFJv1vnZs9xgIryiqR4aC
w5d26aK/3qMWDiL1PXosPXtLx5mIkbj7bGjdRCPaFDMzzaMCUPHALHLMekksJx/6
SnyRdc5RJbThYDy9ddKFtfNmhtZun5Ayyym3EOq99s90vgwgwQdAtAwLcAx7iyB/
sql1qbzDf2IeiKKqFqTIv3whbkRAG7RDyRLj3/gTP+fDmBHIQrUBT/jnw57gYXBc
BrNgIewZ+A8mALDtptwRnUFH4ZCPygIwdVVykcWPcyrfzjOvtcfRJTxSjMCSyaNA
eiJ2N9NHuo9saJ194vpp3uruX0q7jxRYegMnzPaxSO57NSiTw4bVjqn3eMUZVKIM
/STvprLarAgw/HnV7z5EoAkJXlzpdsWcwGSJO9wZFviX4/pzrxMWT9vGUzjmF9/r
vPcxImYwBFvK2R7zoRhwE3AQAD6IijGaU7HPqiTc/R+PfU8yAKwZLFVU8qJmAqrV
OrewG5rlnEU3urK70UsNrtjlXY+HSooh3D7iZbI4lpb667rqtI2Jq+gJ8GrL2poh
Y9Acfeaf0/RY32Hu8sKnSXX32HtVHa2L7yhIP43bm52zIWRU5cElgekdp9hjfjG9
W5Hgy1ZDwNklZj4LPCefivrA+3nRSuBzhRetRi5WSio6kIF3Jd0o5SfMZI2Mww1P
ihHsvW8Ca/BiCndV+gp6U9eMujM4eD5JFQVxUAHwU62fs/tCW5aP3QQ0u0dylxbU
2/H9B0sn8KFjeJhwZ2pH43Ao7W2OkEXrxez3rAvUQviSXO+RovugegiPCbS/2CMk
AvHOdaOpQkRi/hVcE+fN/r8+ba8NfKpNxXTgXYTT7+pNP+M9MX3Qz1KA/tQQEPWJ
w6P773r2MP+sbvQ7HaWh0DOGGDuQD8B5NErrMWE/dAjUNw2I+sXu4tyF7KaZbxSk
GmmwtYqcP7oHWC+6nglORFWCiduzqvgjHt/QRUIqe9I7VtGE5rOr+bm5eN1jkLz4
qNpPXfSjcGAXZsJGVIvHM9NMTaPoJz+OrnBpXQ37dn3T1hjysMUvXlkb4csoFKt0
eg/3vqk4XueV7f4Q0ja/Goldgw+1vVPO0wIT1RPHy+UA9UmJ6hUyIQBkmgKr8Y88
tQhHi6Wfypw3Te0hxIdMFAKRodOzh0fCY3EmRQHK69+ncZoVqp2hSq/2hsKCbB7C
PSvYhBfb6bIPandtaYtO+tsasOGzbewAhun0uy4OLllbOIwFTDUV2cRTUO19/DEH
ginMcw3SDhLv2ysSUIbiPWwGVxwqx1Ys9x0ijeo29FkjBZUuOB57JW94LlzMhkRa
tC3vjgITz/HiZFyqEY+tjXmRwxFIAOOzXy8xs4Od8NpJ+6xBbvoeD6gtJ3AYjqO6
qEqBhX8lkiRtTl0DX4v+/+oxiEK3IXxiMNKCjD9cUVuntcnazr+dDgD1vsg5RquF
riVi0cVF9m8PPn9aY5mUyDIr97P+Ze4WEOtfFRLF15qBxvSBN/BqSJsckdNzKTUX
3eDD6ucUwUDsKnz10fDjfgFFMuLNiXrj3/K+JEXxgCe2WoazQDOX2AgnFwiASAsR
zUrLihqmoQL42wyHcB5/yTlB33jaGxrfNyINu1BZ6MR0BLPXppe7upBKCD0i6lBw
jxAmNBIN/lNgRUkUq1XCexN70JYq+k0TOtBrsZ1LeplaEljK35EIh/qC9z20yjN0
p8oNDRbx+yawlf81cxkUH7UZF8qeqGi8jCYsrINT3PsTUL8MHux/LtNI7U+1AB/l
Az33/gBbqN8w/089shSYcXruH+uV1iq60CUQvTVNA56JxTXt/A+SQYnrBR7+UsIa
hm2hoIT2/2tVkeljJlLu5XoLyEs09GYIT2iyIlaEzoPNbRgmo/BOso7uxgYAYvOg
iY8mnfbHmlt/Kh0NkF4jCnUtxDEzpOxZEl/DS7KsLqq/1+3TEIyjj588CPPtzTc9
BhqsBvHCldVJIzndPXB1U7PtW0X2ARQ50SMRNESYGFYs2W07agnVhpl0C9NoP+tB
E88+1B/1BTr708WFypRXfUaQzNaNcxLkDj2mBe2JtKShk7/5GXBKD3NF9p9oSrDY
2TO7vWTXiGJb8uA4U2Jc1R/XeNsPRcRqcUSzpJF7MnaFuCW9ksoWIhwRFO2bDBKU
ZXXIFIWs1SuOFHo82s0JBfB0sgulIFn8XUODz8N+OO8LOzAzRANlKakh66irtlxl
H15sAbyek12ndLNIlX0icGZkgeMZObfSkrhaNeB9p6dN0oaxdHHLyvcHuEzAmTaT
96O3pMgcCfmpIXZCcaZ8K5xiKUR+IemlyHuEhTDQ2IzBVt9tEQIQusU6AeNhQzK2
+HwbuDMvJMvG3lKcvdzGNEZdNi5TgQe50p4Em3B4Hlvgjomv60eGC4VSKLx13jBe
Wg3Q+ro/2qiBXmiyGPcq/QPzemZESTSMdttvMIG5tDIoAmm3jBxf1CCS9QEnS5ra
SAxQKndg2BwYqPClWSbCA+3kwapvkBNwgZrVcUM2W+3grAuLbbiVExuik4OfQHiB
u+z7YpD1cKaURI0BMZOQsipQbntjr75x4DmhAho45JasxTGoj0lHm1MCZbBqxpgA
z3qbgsH1UwNxnmKZYiF1HGOWYy43MKCTbbY76lk5GF0/sVmF0MtI5eu18f3PoBMr
QG0kRtgzoXHqgxeYwkTNsfTboxt4De/ghZyhlDdHvC6hDmF08Ss5gFgfuHdcpMwK
VvbahVAsdyHJrUY1z7RPhH/DUJqljvU8Te4/CAdB/wrJkqD9OpUSysFhdG3aBkHR
dwzOm3D+spCS4XENKqfOPmzBZNWq69AnflT8Jg2TZ3mI+Gigdrdy4dXi7eXo5+D1
BFCJ9FS6PqwFT0wzaIPV8aP93vgslalmF3vaRuMkE/jvYt49gaFUxwcR6VRelgq/
IlGhdi92dZ+Vgh/g5BWEUN/vpQcWrwrTssHwrouZtOLUIv4WLW27iWF+FUlcoHdt
EVbQ+33BdQmpxvxAbUEnKQniVBaT+J5IJXAgX6erBe/wlJbT1v7YKH4SvRQSG8ns
xkFrWIgpzWmn4Tw7DH8cCq7LPUG8tis8RLehYra3SmBFkqS2dK71AJtmVv/QM3z0
mpA+dggjwDGsBg5myz9Zuw+ZuFfCAxaEEsCoM7mP68HZCu6G6tWx7yS6+Ed7wbrM
eaHThRR2UBp9F/mT+/rcHeULZ1S9XWekL083oBVE8SU2UArRiGYCOwwxQhkMV+6J
V814gKpquRetsxIYxyDy4Yu4QDounjQYp7IV8urzmKE1mjHTpBSOIKEgGcd6yrRr
AzOUapEiCanoPlHTXSus/yB8g40IiZDzsyy3oBIzh5LnjhcMslxAZMYm3pHWR/uv
KWMTwbJHps4NJrgmYEhNQnzKqlXw3t9R84b3ExifZtzS3e2OHJj/3dt0gjSUAMFp
rcmuuVkdeGXQiUITyQc8LmtbTUShm/Qx6XUfvhFeUdKbcjQ8FXufTyVcV15p+COv
7XpcdGuV3N1C5SPTpoGk+Grs95B9rP+rm8h9P0iQ7A9Rg5gMPPiri+sUEcRohZ3J
zQwPzAUzGmWiCtLmvwjV2f1QFZRSz0ChrZYlTYXtqgCs6HzMfoJdgy15Vtr3z/Nu
5rtQopdiiHqU2kZasgLIKUFDJXO4FKWNsT8hg0sU4XEUsv/qK2pEPCevXcZefQFq
heQovimqXyt/jTj8Kk79EUZP3kdHkBlkj8dxQhioxKrkLDkjGSXc99s9kkIuwwD0
VTHRsxuovzftcYzwl/St+oTJfJepilyPwex1iALFpnllkgbSDuxRfLRLEl8ZJl7L
JNEASkLNmjqvzcPQWdm8Ew6s/eva5IHmaX+z1kc2slAZQs2tDbYzd9B3dlW3GScQ
6brm5NHI76sK+KShF1l7+30xKfJWhQuiB4EX8CXwDluwbKhgdjLw9i3+SGgtemqF
b3gVNYlHhis9ZVc6fQ60BSNuOl1fhiA3koQtRn3soC8wYVDrWXaQmcYfFITKLLI2
lH1R1Wu+bLC1/LP7uvBQKqEKBDM0Qoo5QBglTKs92x1COm+U9Eek16tpWXeafls1
0iJOZonS3IDc6gxQt5B3jriFTR6brtB3grBYyK7XaBvDlWSUXL3rmlLf4Agi7Kmk
huQz4XtfZOuaEsVGx6PFm5hRWXwCPMDfBGok89CknSmp9aHa6fSEbU+fZUb4y6CH
YjU495aealORdoxfxwASaBdhgWK395As6UXjI58H8nRzpQx1KFkKV8ayr0tewZLy
6mJxvxWsVXX+X1f2D+JWldS3P0yqLGMoMOiRkh15aCli5CIanIam6+yAarfXhXHw
euG6+cn0LhVmJ4gd33ZBGFURMutcJ4m/T+KJU3kXqOnicurFhsoU06ZKzTnKPnzv
Dp9aj/oNl5q5DjqlIGKuEyl86K6sAN2XGoPcyiqoCa+bM6mgYUe+ZVipoU06cT97
bBKGG73o1n0rdyOqK//fYn00t49Y7sUll4eMHRyixPlfoKDc9B3LvYzoPzZQmtgb
fZ9s4iGh/7bedFvJvO1p1p8J+iQGWOoqtPLxiHiz9milqaTvN8QsvGojcrj06c2K
Bf2+x4We1AN09knMIb4/G18Eu+MNRAtXWGJs19DHe5G+76HFGWZV06GES6+xLGdP
d2dw9bsITVC3rDDWzj22rIdOP7kGQou9Lx45OWMcihsmhC3yXYqpVSz/tu6H7w2R
U+4lJGcNxocIXeGTaMxXjbfRJ2q+fuN/6KiizkdngoNsCvcqQ94jq4oxzKqvqI/V
4KW8YclSsGhSLhTdn6l2xkq/NOGqBEMFObgOl0M+M1QfP43mwvQ70wjKp8MPL3cJ
oJg6VT0sEazzNSTAi4NjvFOvD62jSR9Qi0cpI9z+qvzfO94yaewXpmbH6k+toQyM
CxePvWRT/QpWoFdQVUqK6jKm/yVJCTVeuH4k2Wso8bKRS4Wcw020vt6j5GFrGXbX
eoT1sgdBMvpVgpeCDk+DbxYsjaBMTkrz5FTWuzOMqBSSMnfAFBzV66DYBbOTFQL/
JLFCaRdrekOtSm5FOAr3db471+0VVyoREhN+PE974RScpEBxc1BmktDkPCRFqrbK
FtXIefX/SIBviZMHETegCQ7XU9EFbfrHPsbqeg2CZXhYptvQ0Jeoha+dIomNeW46
ZI7/f/w1iKPj40WFxEeyMimRIJx+E+FCWddQTfI87ExRm4bnPsx6emYvcrDtRpp7
WIxDF+9xvGd+EBD3QFjdxptl7n86Ejs8rU0qXRpaxuwArWYL+I9/6EV1G+GkEpnS
ql0+Ek8gmIsOx+7VHTe4/ymNPiwbI8w8p8IXQsDpUT7axlpSBrlwC27OHN9eevjC
6ZqVXGW12KZnniiGA2PaKHLinjTnBQfHln9eZBnP5zThz1DZ+PUyTDOyItbbkGKo
03cO+h857HCCW+73ETn5nh0B08kMEl0fuMKzT2zcl/OwblRWYCoCOuDICt9nRzj/
TcZ/dS/nlVxXxCPZJwIlloM9SeOEkjm7op4R/ly5yia4NFJruiVLDF4bQrg1mQb6
ccgCiCeD/VbQUXVw+rQjC+DwITgSCKjjXe3qT+EXiFg/m+wEFxO2cIz52MmMkPIM
Wg02KhnF5oG0sxbMon7eZxAX7Ni30LmSICyaUra4txSQNwWcpTJcex8kSKsJD18+
6+8ssTDOZNHShg4r0rTeF1FdSLNrqGE+Q/Y3Nm8fYfJj2XTVibL3zKGC1+gVuzF7
unb9chPrjGopy4Y84xjlz+2ME9hGLk3YxiAJEpfYJ24V94QMTEtxSwL/x+P3ZdRA
Si98kAMHOfwJ87qZs83ihZK5QhA2Vw8EEtndvUPEhSO8hRwV7Q7F8Et6eb4dLBcl
XXR7q/STuZ/A+Dggqs1AKuEtS83xYiEieZVeI9UpnufAjRuiAF7B2XuyGVLcu7Q+
bP28twpohEUHAPbfJz+/ov42u9OtvhF85PoH65yYPxmueJHPvxI5PXNRkDs0dDNO
wFuoMRjr+o7opavr+6pIVQIMEKPaUg6LAWpN4fxWzJ3dSSFNvpFOiZpxqyfRYjO5
JPrO+QRHCeA/GDxOiAiGxnUh3ECfTcUfk4Gxo2D8CWX3+tUbED6eb2aEmkbQIHeZ
GZ6AQiiQLIcy4r/uzJ7APlgMFOZqVx5E65R4NfcuxAuBjUIUOGB0iaOFWB4qmeJd
YOE8FOt95DUENUb5T0sFt+spNpQa3j8Jpt4j5Dyfe510tCCroWryZUPDVUk+VL4L
AZJ7YID69TTZ4bAoJG13UQrSCC1D5RVWQBEmnwbq6TB2wlWdFMjWQ4tZjdfFK6Iq
VqrD8w/9u7CNsx7CsW9CEiziCX8pl519zRLYJRZnw/UUjQSeG9uj+ve81PZDM36R
b1dhVirbOaNqVuGVNOQJC9HmkNoGYrjcnXHCF0xw9/tYz1IaxJcsm0eIoXNDpH9v
1Vx9GFE+UrXOl/QHXleK07yjOJdziN34kxnZc8yj+bo8pbCVLt7wYl1xgZ/Sekgm
My467kYzu9eoM0qZG7a1MmdbqDChJHiDWWeZDK0pbTMuVHh85d7h+QI93wzUhbvs
5sTZlDTtaudMpe7g5r054lFe6hz6aeqhsVPpipQnDCL1LOOmjC1lbq46qoYCoVjJ
rqbputq4R207+JOq1AvRoV+eQYfoDANHXNtGq+9uqK9CDocOi8ofZAvYxRROAXSx
K32tCPbYerTt2clg9Pv4b8vWIpXx9RZuncw8PuZ4WzMG+bTp0RCFwEnKPe70QQaK
BVo5jvtQ5bmsAPkrj/2CBS4F5fSuCTr6pQYjBJFhITq8SfppbbxmoWx0IpC1lz4D
F8aVj5GckEFLEChvZIfOookiwjMQuEagc8Eet869tRRogrq/DfGeoOewYBypIjSa
0C+tXukVDJMchQquSUFPxUJIXDa6xOcQ5+r+QbjYrhtLxWSQiZzaPjz3/XZIxsQJ
n/vTPmLZ5e62ELYb81jECk80qh+yVDweEUxTWyVmImnARbWVah0iuayNHMR92C4i
pRGjA/rORSnxzOhyKqffXnd3mWnqKDIsfUH2ID7ucnc6ZSJrmvpSLEm1UgMJKg1H
32lFFHrKxO68iiw44i4wIFTx7basMYbG9+SyqyZZvOUH1oPfrGkw+9nVNAMl4d6e
L83CgaowbrzOP1P2tlPctpBsSnDcvXMc9vbfkQUSd9DXq6dnBSm4ESLKABwDckId
cAz+ePdlY+BVCilq3anKQnqQ8NX8SsGeCaLG8bDuakGTcO96wO6cq/sQ4NtyCijA
pv/qrrmIcEYRAw0zCGgG4t0AlhHc0ahv57SY7lNBL4eSdg0ZTcUM+TO0bYa6YnOZ
hmpbzqUEvcj9DLdKRrQzsy6VnaQ+7YOWadIFiKlnOPif/N8VMMzXkmopaA8wbx5E
x1A7twsPtn3oPMHh1aho4UpVNm6DmUwRUZHc/mMFnp04BUHaPF95JSB62dgtZ3TO
JDP3dGQj1t5GOjOAr0j5hhLbbo+ZsIzxTaP5viB68AJlbahbXu7maFgVGAn7+FMB
Znqji3ayNKUflRw6xzBaAtW1fcY9iug5nLf5A8RZf31FAm8v7gGN0LlPrh5l2kTR
oiveEnbqLEjIDiol7hsEKC+BBH15uaN+jStiY5W8tcs0HX0jrWpcQAKlHOGAzqIF
9W8DsO9/4Bouq0r0mvDPoYLl/bCNtiIyCxo9EfcpaO6Tyx93FZOqN5qZOJc1i3Jc
SEI5yg00i1mDEvjHD/rxlOeW2RMFi/ufVjNMN0ZBVO19uttLa1csry9oCITq2BOt
AypJYRYxwBUwJvkeM4y0UWIlP4dpJREk6IZJ8aPLJioYCD9b7MNdhyf7O1cy17HL
zPgjWNFlmjeJdo8WMhTS8nSF5OpeG+gTulynEcJbpwVvYQrKuLs1suD3UGLQn78v
tVxFh6Y0lg7TrREBruc/hxgs5L06JoGr5NXhT1St+9CbAOYwCbWRidomg2iQonb1
zzCmGVK/fPHaF8PIVfgidNn4m5AWze8dJDa5VVmigcyw/GzizfQ5h3d2UO+RLog5
hjTtQmRx0WMHJbmFgSqkf6eO8H+tMnvPBXpN8hltmbhRwu/JBBgIHuUZvC2Wz6oq
W8VnoOfNtKdYU/HQKtCQnkVJKILjz0qSYQEZbHcqgsA4ALewulx8GDgl+wJDYF33
/MeOdURhduDtNsV9cte5r20yVAPGMojkRfOGmra4m7nbtNuOuI4bpLrDbMII6oG8
nZyAdnH4Y6UNQdtq0z0WunRa6HxBy4JJOGerblRrNlRdNFHbFmtlaVq3BoOeD4g3
AlHrFfy3B70eZgt/W5GBGu6Z5wh4gY4eJAsr9hftqg3Rv27XcG/pB+NF+VZZeHRZ
e216N8zWiOf8w+RuAArNi1hYwv1EKNPBMUAkD9aegk2hEFKiK4hhk8/LqFt6B3o7
/gflEFv8uXr7aWm+VixcaLXL457tPtSNG8jF+PNXHO8FvSmMa9AOMAZMpwsCZ1Q5
90uPbjwb1KNyuqQHaP2CS2uXdlato9Ur7O7y+Vhi38JjMiCjw9AygMUhEu9Dv302
AXQg3HQje+0nKUANGd/6Gep7rl+n78NP68mSio7pa1RgEmFJnLW7uCrbIuSkoKY+
5EBTut9G9TgDVYuY2uSLFFMpytsDaFE5nHKmRoOBrADjOKZZqLEbv8pZxtgM9gM5
t88qGJVBBZBmsGic9lN7oOPzysG7Vfm+EjPPngJ8sItB3qSc+kl7yq2rk7jRxLvS
flEnvHKIx6P4ZHS9L/2uvow736KVUk5LtZ5Yd7R3SF64qNHnRJ+iwWBKqimssaco
m6wgFwEKZQuQriHpH8kSKSCNyFrJ9phz+qwcAFe5kSF+Wj6jeIUtQ2dX/9tLLvQa
7dtahyLTY1PDTKopYUuhX2DxLDMqdInbWWHWjJEmNnwZ9XKbl+Ow1FVEQB7yYqXc
5eoNaDAqSz7uWT3K70svY5s2WRd6npQGXU2FyDZD6wueusbilT/0DvIVXXWcgCIj
M2pICNNVW9sqXr1rJ+KDFfUvIwnX1aIYZtXNUgwmICfCfsT/XSJUMuzY+GtoNVFc
StNC/CgiaWI8FMYC32I6TR4e3j1c4tMNSCTLqCC9NtqI8IzvLJ7Q+KdVjrV5t2DE
wphbuMC2d5DJvUN7w1oqt2o7N374vdea0e1dTp/8NGZtAhGPxPK1/KHjt8rGVQK0
8YOxIGw3XGpUVu6+JndDPNdXBsYkD8qasCYVyjw7/zC8++bf+L5iy5lQC4wDb78k
RiL0GmT6hZq0EdALkCSfQiEYWL0aXWtpN2rFzFNZf+H/QbWN4CyymqPGawgfu0qx
Jzb6qGxn4mzmaceK4EbNJY8QYNpRDq8IcwLmIqcwikiH+O/28INLGzrqXZYiqlEC
KiCXMu675MP9rO57vLoFTQXO9fkxTia3ZtUhwPw6nWNo290Kf339+mnIFSvJ4Dcx
Up772EXAFK1HYyGK4IgMqSbfiQ4OuCUvsG1RbThWuTpYpYwKJsWX8QN5lZVA9mL2
5yR29ymEwAL72bG9+W28mI6s/nT30sKKy6djWQu7e/7QRpE/DNRPCZ+RsL1o0Bj5
I9jT7+xchUR+QzIAbDUZqS66RBQMEtz/q32w2LEut33VLxiGPZ+9Xz4NPjq/GPlx
KlbUISKp7HX9KdQoosLDti5vnl78aY82MRHa1hBtVkqlOWwlP/Gf2mHNePFlOc6c
yvY7zlvYhez6RnmfOT3gQ5P6OiKS/CEhflaaWeF38YtlxQqBAPgcktCfjDORDukQ
VzZmtUaOr0enXkVn9lU3JScR7b3gYju4/8HpWs9CBHejaxF0hVcQHiwqhpv5+cXX
VtWm1PrK4izenf6dmWwtjwapcBZsYcpTwvEL48Fcz89snTXcJCUV1nkA4mdp/ZjW
4qO/aPEo8f/z1QDtRWaJk7HHAGddwHQbOJAAK5bfUenoR4tC9+D2r3ovQKyar4p2
vNwJfzWTPxkqhQSKGCZpr5HlnUSTP/O6rZIjvI/qKj/cx4XUc1k0+pSJ3t3M/gf3
1upO8AuTngIG93t61BKFhs+VE/WayoBXgHQcPgRPxHQJQxtDBaQSgPH8xHLfJtjR
uc2Y28y2eUMOKMPRgIcn8eizSq16getEkVCYXmVdFo2Yw1SdLA6EKJEB8e7SfRwM
Us1TQUSehM2OuZuv+SpfVtH879iyKusYQCbg9WkcgBZobo49x0hYvSbAU2kO8Kr5
VRdb4yvo5oLIQfRWZb7d0gxazgXP/o2vOqkz3h3NvxBtaXIXiGw2ABqIaEfaHNo7
OWy6v339amkBWdLNMJ9Mx3mZ+WdVkPTzNo+U7TiNPYzlTcb90HnKNPSwCOvsIE0G
cik7HDK9WQfHS+ytkGTBr3lUrgozHfe0nvBQY2wlOlYcf/nLsueLW/O9ZRdm6Z0M
9tth4E4+r3ZiJox5wUBJy+ZNSSVROot7ERPDWKVisRZpPxeGwiUNRYFH0FiwPBla
VJfPoXVMVUuAdKpNl+7QPrGZhdv2t+1hP7dPiXvTKfFOjtqiy+UXU+EX/GefkUZD
CB/eEVG/Xw3d9KJTI6qlu/sDkAgpdyWvcEmGLuJLQmwsJE8PB8sDkYaJId+EHpgT
haDlktwSJrZEVb1yl67ell9R+LaiFkl34WIM+rD5S5hn5FAC9h8IzqGF0BM2nAjX
VjX7kb6wHEdcYreIWZNVdFrlTHqBD8lmT74lvobgYBUW+tJBzMWgCjqBWPXlzH1d
fQDdaphOpeQb9uFH42SDI9xIwBshU3IYHUarHrZ70rijoSH81lY5tVxnS5g5ebgE
j1TKVVP6khqXZTNk098hWzzv5Iu+EMsaZmtQAlKCP+Y9h9KpJand51IkO/4R0ANw
W+MZWaYIsC1DHwqtREjqxX2xZlIL/EP9X9N19AjGLtxYUZ/jLbLMTKoBR5CwEtZ4
uFaxi8Q5+yoYmysjdu+sP1KBV5N90ol4D2ByngG+GbWUCFJ8YOlBBFNpiZvZKjtq
BfCn8DKdwaIadKvAACntZqX0ocB1A/1B/qP0uunWh0nZOw+jBWc8AfxN+EGw5SxC
HZMao1EA/qVeE341GpY6dUfP1bTG/c+JRCzg2M2CC/SEVM70sev5+Wc8kaP7pK+r
sqfKcufMGjvkh42a1fEy2XzLDgOfuCdSqC+PC6map02Z7EOMvF1S4eWefYvBJJXr
l9YCdWDD4z62LvFR6f2nXiew/iG9ugRBBJ0rRW/cJrt/Dg03B6xIp7dSVkbrS8Lx
Pv6MR5JDwdPcstTo/RJu0VX5rIqoZjkiIT95+xNaPRv2CIutooztmZcqv2Z1cjf9
kfQ2NxDCL1q2iSqKEWuqt8HSCOkc2dDS3YV30pbCCrkVZXhNuLNLvgXueRYUrhLG
KI783PLHP3IHhGs0fACPWKOf677ImSBIYoUX1fky/GBANtgMn5j///90PCNEqkXq
/DfbZU9ztZsNb+Hy4VAM2019WLy2hTap0hX22RMv4GpVTWYdBY1bpBBvMNhCJb+3
Qv4pVCtDBVqVY04Li3boyOXzAzVq2bj8Cnw9wetRsiCz1hh8bwbzd9W34TvRLmN8
QitG6oAwMrfw2NyW21q7+UyjqmaBcsux4MSMpVXPEaotqiLmRUoXl0GmSU+gP/vj
4azMbvALvskYLif7oJ04ySjQRqqhx1lnZEXU6xN2JhXQDHJB4zEzdAgWmX95Z1Do
J+bzNNk/G8Hb3nTOLFQWb+N3VT2zPoroJMpJ8a9bBDkF8NW6fPfjkzW+3yHgnpnu
FbaA6cR+utbQeWE9HzzMWeJorUVM4S8BKOzVcsjxSV+Vfm8KjoPBaFsTRTrx7e6F
8MMsxeJSO16APZ4WEESvZmR/PxnEUTi3sHbrb/GrIeb7BCP/oum79CCZ/mTqVgyP
LVFfmfG3hHbVvVeDjeVlRXxWt7371EqCe9sMaIo8340iV7Aex5dO7jln5c3f9scM
2tMi2Vt3Fbd866+JoPNpTHSZ6vTp6NjXfD5cy/lzddOX8i9NRFjBoebewmzoqUjI
bkbHoQIv12fxLMUnYFZnEd2X6ywbQ7Ifs1mdQPbFwWTQXebJ7HWoINaIty8ocD2Q
j+CPqm4TX2ny6ryqXASv31Aj+SkCTg1zQmPXZ8Fqy7Xg0AQdbEqVxCRFGMYW4baL
QsS4rRPJKeSMIX0Fn7OAgTEIPW84UNsPz7/xtzsDG8u6+5276RsXshO7NCvBUoq3
bfxy+vIM2lvy5WaNiY1oa9z0w5Rt7rhwYUprw9FgDKpY4Z1Uq/PU2tWyv3bw/mS0
y+frE87cxOIv321nGRd+VdDJl269RPgAqvei5UzGTU2dWLCyqvpN5PMDq8CAcIaU
FVQQ1tlPva7mbbz8uQ1bs/FQiwkyhcNTTf7QGmYOrm+XnHBGaFngLrUhtaEWlHVH
vov4HeTmZmahoonWQ7nY+lMg6IY9HphltdVAhwNLR9QT9wYBxbQYZeEd+zxD9riM
CMHFFU4FNXgytoJwTEeDOdJdvrI62JT20B2qJ0M9BTbom6zN0tZAbdVEuC6dJwBW
jT4BdFl0VxKisj2zr5G9lk02VoMFIcOiYbpbithPNH6i4oszT+97J9MYWUiPe7Tj
j2yjTX7RG4f1c1PD0pWpl05/Virci2l6GXSvsqFFVU/qRUDrpPs7zE++VLkFylhq
LnNN5GCCXQoo8CKkkzaaAkoBk04xeWiEOXrOqSawYMXE8oDjWzWulmWj9ftlcgNS
Zdv7Iugnb+LPpMn/djObFdQZukF097FMIHcbaCcDV+vLTbpOcjbPC3R3p3DWKCWa
zsjPOBH+bLgDm0JaCO8cF6eutw5hCFSnZnAlUv5Joc0Kn08PiXc1pICQR4Id6oET
FauUxccgEstZoGzgkwHYZtv6YP3C9GcJgRV6dxVCzskfvkTmSqBTP1u1k7L+9Jwp
bbYfEc8NMszLxJxGWrbX7018JQwkcYHsOsViXbXcD2HySAUVkfxxWJN08ZQrSrui
AUoizOraEEz/WvXoOGcZQzPpQS1V3Wp9UBhyMmBV3uw1/Fb6RAlqWdVNbY/GZ7Mt
UZ11TLriuCrxwV9YjkR6gNIyRQ1NNgepvok4QG8OICKk+g7qXDv+R6ICTpg34Y4G
ZigLv0Axa40tX7BNayE1ryXSD3sIsI3JRI2VWTN4A9YvwEMC6oB3iqkPo0/4OaHA
daMqvqK0pJvryBlZD0BJgn7idTCYJo33t8h2VeNZ/H3JAE/kaVu+c9uJLzx2tP/C
W+za9+mZ0K4cIpGgriAX/kLlYH8CrtD4cydDC7PhQMOOP33OPvEsQbIUOcB7vyEA
PEpop/bl3K10cYiblbEmnAHJaLIA4SYEdj5scSS4VM7ltCM3npZnz5oTM3m3jt8s
eTvbjfqTni6UjYee5IWweo6bhmYued46Rme5gTr9uM90vNEFxUF0wCXapU0x992s
xykAKxHUD4JUHgL3FowvKBj1bgY9Glvm2wB4MB/NYSRaSFIN8OGb0mqlXNZ55k4R
fH6B7zM+pWGiTB29tXuxWc+GdQWap1mPqUSWMPdNU0QwcjgiNKgTnhvxCdclG0J/
aqrzdvndqaIY8tpjp7soguNKt2vQUVHHmd5/uZ5NaCCNDQ4jL5cCusDRQlZwkpec
g8fvt5wwehxNlnAL87/5X0eYm1g1TxqnOTm1WmDLSdP49y0lbOXHt7QAfje0gHjF
yXu4Q9/jduIqwgU2wxQQ1h0gic+ywymh4Ie46Tmsr/jzf0Y8r0RiBxzCOhL43663
D4bI4iU2ycz/WgiJscQl9aa9UHpdBtTf4KVQjzQm/mCaTREjoyCzJZHMPJqKIWXw
Z4eg8G1Bd4JEXaTl8Sj75U9pm3Ui9TKwzcIC6POOsKToLOexNoEy67J06JgV9kkJ
cxNQmZW0xUgHGu01clM4o3nxhce40KnS51AvdNaz9lVFvC2Uhz99ATujPSEP4UBg
flFmwYsIRRWa7MundmnwbEnEgJm/JmBKYn5iEF0rISc2n76tgjX8U+k9FIxZITcv
+t0Kojrj9O4ytJdBAQKypZ8qzdv6OcjdZb+ejtnIaF+BKAd/1ibQaLuHhNbvkkMF
NQJie3b2vUeS9rQ5vNxNIl3hdf39r+CXk20hjERjm0TQ2GbBrtKJ1FO7IdY+snsb
U5ZPFc5+1mjXHeGrnEjxqG/97uZcoIMuNfrfA8GfNhJ0KkmA03rGitS8nZZUGlw5
iM1qgp8sENVYGeGJm+nf8Sr9kjBGVe4CdlY3frRYgqD8Be4yEFPAWGrKpk+emF/l
99xqepAoKD20s8i0WRQ0PjEVZ2dKT4eQHFbmGMLcD00tz3EiPRvgOxAw6GPAeCvX
Gt7MzUNtc3wQ/AZmaAkxzf//jb9riHn3p7htljGhuWtXGv+/wuron46GBwFYWUxE
sux6jEl6xoLmQZUhkjoP+LsAnc3GzjsWJzgIIW4Li0T4EEvYPYA3SDWSQ0J0ANpC
r6SzTeBGrhgRZSfOimEge+YqG5OyfpEV7TiJ8DyxTttpcPV42F6w0OzyRkYpF5Mh
J5ifLyRp/clQy1x1ulGBbkMcN8IZWpWfrfaiyuz0hRBLL0X/eu96mai9HG3zXRes
fxbTcC28+PTbuETG9s/rxZOXh/hl9QoTenEpxqmzProrLeJHD4O4vO+TCma17X2i
aPBnwVzpts8ylALTx36PjCTSbw3BZpDqwKNK4TNm8XfhAc8p4jzAFQwLRizyvcpy
Wkj4mzrJXC51GxJFYVM/4FBTRf1nTgkmZvU6SSE6eQa6WsiHMjBZ/SNh2/YSN0ta
vukmbl4FEvO72dduC/Ycy9RcJgi3fyVB+QVWEyLczHzgrCxril5lLPDkEztqqTtS
MMFrN5LknfkOruSi6/AlSKtP7Xq3JgNuoBp3AgwrvX4sNqdXNlg6F7ANk2JyhFQF
F9RQYo/u4ZBqVCTBspwt799zxwHogZgvw23Hlt6OnWRK6gJD9a9JVXLfT348RyNJ
3T00OiwX3Rz2KrNwNYQ5ypty+hVJ+JjY37ZZFzXTk/fGO6YKAuWxQ+qWaohtQDzK
j0y/ymydPtzeSdOi1YS/hez7n6atQA/p4Com6k1Op1xxEB4Tk8tUuKjCXnevMBUR
6T7TxQiHFj3vLitJFJ9mUUbV3XW9E3rhm1R2tkH3H2TS6WeXPZO0ModV4BHvJjka
Mm78Wj9PY4pWcRWJ2g3ltqSYIwfxcz28Iq30meK+jEHCI/3FNp36VcK0+hCE60nz
2/GmFOUIbdp9887cPTbPC8BvPnrCjoGrgndEZaK3uEXK9hfAQRbsNCW7+PyXUafu
VSe1m+/GWfMdbjWRPUxReMTV670n6jIsYe0mn4UQpU6lxhhU+VWvrXSNmXC4m7YX
3ZcsuwiMEHbIBmcGQAnzD8M1XcBjHEeu3qX4EDJg+8IwMycTXBCs3PytesQPWW5W
w5e0++wfaAT5pcNxcc/Qk5LigI1n9qv0yAmjwI7rVBxd8TXhX/vFzaSkw9dMkT6h
iLYR3+4OTWzHue9p9DCX1rFmLIWu/4MdX9Jp5Xl8vuJeQxKx/vtYWte2akpAa6Lc
pTPbvEv9H56uq8X1Ni0Vs/5nS20rQXgCKBBOUzhGQNef909EPRoakZDeNzAKqs65
iMibd+No7NbG+k31FvtZANoJbv8afdgwp/XqOhHBDO8BzcQ6Tjuw060U0gdz5o8N
osOeliN00hKf8d16THqHkE9trtlRNfRIUB99mWKcfJOo1HNenkQ52Cl9+YsZeoK9
pDi3VyJIuPLYKk0985nzVCfSTJFp1haaO7gpBRS04iK8MqdZamb4orsmPu3VH3E6
q6MW/1oUVDB95mCR6oRHymKSJfjN4SE+gHFt9hEHyFl9BWCz2FpeBPTnoi8ONIqZ
nkJX7EEmp83UrNTGOfhVnTPLNnI+M1cHIpCbfVGV0BrhGyEgTglXPL0rL1T5I3Fx
/lkFqVsvjKVT7X8xfQe+0h7ibtb1U4ynTRJ3MYB8zVckNAqGQx1SEFLuWXvtCVAk
nj3LNCODnTBXrtQ7bU9iAq72ul6COrtjbL58Z3Cyv3XqqNCJcGf3q0Tnxb8W0Ppy
qtSEuO3oj8Xo6WX9UMBKYoSguW9iehIO9DJZezyL+fI5czjAY6127N6YF7Ddejps
HRzviTCY3MT6tfSy+waIE9Q2kxsV9Pyx8Vm0m3FlPW2wvHrv4AeeWP0ntN64PKHG
nDVrCduH+zMaBy7L/3sWfSuFzIRGpOeD8qawX/vH4xseUZfZXe9wz39enMSsIwRS
uBVmuvh4x0ZtxKFsDgUhzok5QngXcrQDsfH1bMYpstq5D6UYsT3IkUIl+VSt/mj+
RXH+KEy+E+MDggmBvugj5crAvHy/CMGoC0KIaI65ScnpStUMbF/tdhBerQa55sEZ
0UrUz9/vYn5ix9z0vJvWAFB7o4YDphDrIE+wUsepLnAsgk6pGdJhM3GIr3l7K0+Z
1roCq6R/QyMvm89CbMwQowiht7f8Beax0X72mg8CoO20/uR9aW3kmaiC5U7lLWfi
6454z4uIROV6R1iNrLIM3z/ufSLj9thlaS4DoTnU7Q/BOebbtQxmdK5fes3FHTny
0Y9uXYAWuOt/DooC95fNS2TZezi2CFYrtiDmnZljec4wpBKjD6aPQLttQfOzQH6q
J5GPz/PiY6cRUh6FQ7RgC0bkG8p+ued7x9bo6wUtu7kWrOrDS9uEDXcTsDppO3/U
4Xj4ggV7AkhAep4ip3ZUI4tHLg0fHAI6+f3+gDsOzlcrdrXMy/vzYZQzkfpOj/iH
NmeA5HXu2uYS5F0r9JmPOEKKo2G8auVbtbdpuQhKQo92fe21UoCjOY0KhmBIjHr4
tHIjGoosYcbnjJjAq3cvt2iWb/JU1+pUOsZvgg6CbL9EQQWYUMjT1z5iwhM22VUk
YX2Yks/viGh65lA7wzqWvyusp56LZqj3Q6qWndWeNNC5Y48MreIHqxVAjZlRqJaJ
6/8IxJtio9Kfti1LDlWqWI0zFdyZefsGaJ5ounyv6BUKbwre/f+4maoboEsYHRuB
v6P3ruEQxcw9EzRgAmtfsSAwZvmF1LL6OitzCIH/nBxgMvnsaTd1zx4S31euAUAL
ILExzWRtEQWAOL102sfjKULoewdlW2h/+IaNrIOvQEiHYZsGJ0A9iR+2ECDDdWvS
4AnLyK9aHiLc/s4KlxuJ/QAMTcucd+cFNtTFs6YUDOj76KlEBxBHTNXqjPFJI4+E
W0GCYf8MhLhF49f/Njq9zBbHlrtVsEYKkdnn8lWjl38asMQam6aM/NC/dOMXyUf3
LwADhnuSyNj45pMAIMMhZnyLUP+0yeOMZhuRPsGNuasjEPZTt+sMy+96jwxCF3tu
pFhhe+EpnGGoQ5zWFTMDnI6QsTuPj6mRGzszHU8dgsDwLL0/8Lylser8/XL4LakG
YiHzkmJ3iAjZX6JKxbcturZixG5xqnwafoWpTEupVq5dFP4kSJ7mpt3u7aTCThTM
9LkapT5x6sYsQtR4oC+DtGTT4seQOV3lvQou1kgmPTH4I8y3zkJxM0Wci7/+zH3K
2hd/2t/FSdf6IlBPCWgBLKuY2hdQwI3A0jZ5HA0vPHIC4v9waXHZMwf1/H8Zk5U6
+poPJj0YYiS4aObBRosQI6GsexhRpfPfmCRsIuU4j3sf851I0SMMADLouQMGo55y
3k/SVxviyV52tF0VwzrG/7uNnZp78IFZ5IApTe4dt/u5ZsHY+QU3Mlz4JlqC/yOh
0COQ6/AjFeL2wz1+4lisLHPIRVFg1axwarjjb78J9mwzH9ecwlXa3O0tCX5I+f2S
rLMT1XPPh6xCXyPak3j85fPUEdPvTQwibk859gaYN8M4WGe3QIk1l/8EzsUP1NAx
zHhSYhfeL4benKe3xxw1r+sVC8SawxFqzlKf771JZX6NUW1k71FIvhBVFU5vM0Cr
h9dZjxwqCN5MzNT9zm0o+ISIISsda/2RJu/XBai5lBHClvIGMooiwjtfGhylHP0q
TcX5+jY06FSkcW79REf53lLwTuzZvPgurVEGME9fSkiGk49mwe78CiP3Wi+nGX34
zmGGaMpBm2OFeCwafutb8UQKxTWoS1mHdTzfeEIjERhKQIJ6+jTDYaIvxIeItdWm
lbLsvnvGnljKh1jfXwbbxkmpN+49rC6w3rO/nNqpvY0yHDTTCS1AmYMqyPl0mMDe
8OP8pS8V9Xdi/J/sOcTblrXvUiJhxA8d6pGturLsltYIbrHhv8YwT3Cwj31dXMMH
hJE66Xbuv1t44uI6ZK+VyenaMgNAl92Au1RZQEuh3ABHoHBPGhRpfUBG7ZViVKgJ
RDXDh2pIcZXUAdO+xA6wdhnN8YVcByEvLrTes9Ea8CSCqQBMi7Wozi2W2Zdcw2vs
d3obxFifAPP99J3Albqx1dSAxUG3VYFG0WuM895Pdq+eFNEYxt7+4k0TrndZyKHp
khG7eK5JrybC0OxNBg68ph9Z1JuhijB9u5Eq3YBQ8SLOQ3G+rOVeTUd5bb8yYz4V
XD/7rCDPcU3IsJhRYEKBvY1lNThpurBMOAxgJLQaFiQM/NKKtv8cr2RfIyYRnNW8
V++SnKh6jSfBEkQVwmxNBtBoCX1WVKp/VkQKrZSO6GGCNxtdET2Dv3Kz5Y8ew8RB
PjY8BgRlHzM6DxpTyYzTj55pW0SNUA3oHt+dodpPQBQAnBPOK+ZoKpbjyG1rMtx9
j0UyrS1/bC/LhzsaP3WGW2a7kTO9Y//9NhuBEGlY3EpUImDsu9VjYVZ8PlijDVv/
LxAl0tflU/JDbmlRu9+zEe/Gq375hTlMCbWS/k4Dbf3gBC3soeoYJW0TcdQ6yoXf
9BduamqExjqkgultGnphe2v8+c5OrlzOvzn5zFoSlLquqjdK17KTqvTiu1Nr2Was
dmuzd9ggz4mYP6Tjk76AvWEA79h96Us51S6FMUltVpr7V27hhai5iG56GXewhmgx
zx+lEYYfRij3nvOIeojAA3FddHxRY0XRpWsR1jA0CyU8U1YE3tATkMNIlFPhvkZW
aIL2N5k/qeorPYckfpyGScITnHUz7HjQvd/wL8agsmwTbwQOwQTs+6AcURS6cKFi
XUDlfZ2vRYmnqRjbaE4i3Q93ZM8d18h2UbyR3wE0XuH1Ys65dE9rltjWsHRu2uIk
qLRQagrNLc/3R5/GIVp7xwJ5IytxrG4+xK1lyGK/PzoFPP3ODEFbxBXenMqt8GD4
gBf4ycOoMNYiCFBeCBazkpN28hQvuYLXALbn4ooj7M0FS8ZtsIQ4wkmD+SI8ub6j
Wt0xh9S6opFrhF0yJRcjPlDz/N3F9/r2m/6f206n3nic0Fvi8jagVTDE/WZoE/kK
ZMOdC27Hh1cGseM4wT9Bn/exCUgu0fEs7TaQjGmUTjignv3P4HSn9wePIr29vcxa
TjRs/ZXklZ4qLXCcxERGrnV553hvq0Yod+s4ZfruDI27aqoitNrmC/LogchvdCce
5KWOwfRTi8eS2aOnIz5+YjZ9GMHIoBPGZzl9Y7mHXa+pOZV2NYMwRBNcL2/wPskK
xd2MD9eyxeArygKmyFKrCN6cdQ9TGAf5soO4vuFiTagCttKPhLgSf8+l0laSPjdL
Jyzxbr06Exa2aSlzFw5zNzBNpHEDIha40eePzHu3pqE5lRNvp0ZyYmZDTysmUUxk
9DTzjDnFjx0gL9RZSWab9KUJodn34xMfPc3/m3KhKVpIhveFgazt5G6LQJXxX9Ui
3GtU86wUUMZ5QjeceLUPrvIAt2mIV3fABixqfhNaX6gHfLak3eP4nbKsw38HgvM8
Boa3uSBOxjIavbWKVjyFNddFs9JjLDwLO38/Tf60Kl0n98rTIUsRs+ejOHqrvsZD
RapS7NId+6Y7yVgsdb3CE9hEGl4wYuQPD2EOhfKg/oITWiZQLkbic8gilh1G58Ye
ukOcrB06kMpC1kUL3MomteuGwY6MFVg4VRWLPz1EcPOY0MutTN1zXcWE+VV7T9Dl
4LIHSmzYJK/euKTSyLqyLvrF6rsjykDN28VYm/3PCFq9e3KrEZpCWGRBxANwGlJo
VtZhlnGlMN5P1tEB8VUINlP34I58l8+wTnuwpLDJT0Zo7G7IuzH21py//UKuXXXC
mbBR9pnVI/2uz/6YTpZqxuzcqoWS6tMsBv7CfhL1O1dlgQHWJ7kMZxHAMTLWb2IB
fUy+ta5PgU8df9kTwJiUn03braUdf88eSB7VtFwisAH6eO1MQADdxduYWbzu4yE5
yi5biosCWpt5Ci8j2cr9f4ghUHs88PvgY7h3rBRk6q5t30CPJ7z/HwBf+NMDH5Ac
h4G8bJc5xvG4G3xgJvlXfQSoTshWkrNrDeJNIvpJkYpoz4T2czloZsrzU7YWUQ02
JXAKnyLBdZQc7fOLgFi6+2TloXt82nS2MxiHRWB2RSRQigZwJTQ7E2pQakU9YA5o
12gb8Ekjkd3Kt9kolvDHCIuVk+2Tca+2tgUGIIsLJQig3HU51jPjuAi+ZKthGqEN
uqZkCGH7IZr4Ow6iXXARM1mlYMYL3PGvswntuD/8JXHzsxn+MYwf9FmR7s4SLU1l
NmuL6TZCPVT1s+9H1P1Es7DwgnLe7eOXAkZnrd3trujeKv8qHX9o6a4xpFj/2oxn
D89GpHOygHutl2qUy+3KZ+bpm9EKkwrI9yJYYySqTQ9vYGvl/wfstUCktSgSShw0
QhEOjANzbHsoiJCy0yJb5Esgn4m2DBT28KuqoZ3S5/0Jx3b2C5Tncuj1ucffZeVI
NN4dJx5y+LwwBtGjzVwIXaFVbbf1lOund/nU7P5r7Yig8zQceIxDXd5tWhJh/1RH
R0Z9YitNUUAWXu7HAX9WjhQAN0tRqMWiQkqI84eW36ETUYRxi6MkQaa9iSPihrvy
zrWD3p0dHJTpNBbE4k10gqpFTuqhxRGF5PDZWW2A40MSgl787DED3fH2zpRtTN35
koekdWj32zfKGLNBMrozm5EO87eJPZHbVkvT9QPke87Nxm919e9oR8eW58iHjGlN
2GYOTWefJ6jfmoyShxvSwNCqUw9rPmNvfWlm2J6PQKB8aTiHcvxrcjLZfGYEspPn
ALkQKSvgi8pfKOp5bkJHGU5tv5qlT+gWKv5erRvIBmb8DNLZiqgt7p70iGm/LwXk
BjCGaC4tFdUuoEGgYzK02y9wMIIjiypN5iPrnn6oXFM9yL+e4SLjiQ2Wb1dYBk6q
aL4DMXzb6jBLkOoSC3+Ef6X5guv3nzrZ3BhfAxMPu+bjqCLfR0JTVg8k8y63qwIi
bRFjFFI4yELvRKBYlxsmIhsa2kelErH8nj68P+0cnQJLgf6tyRbm76Bst5ehOZI+
qAJR/xtr2zKkuPk3K6uws0IwsyEDTa39u7zPUSGt+nc1/s2aX8YXRgjwOPtUG7mN
SjZfPzNMs/oy6P3i//S/Y/OmFakw4xjVynpbmEXK0Jl9cqSCSfyaeLOrJBY201kn
FlyXAeS237YLzb1dS49A5b3h6IKDJZq7JqMmXDQyE3smyjEBGHZxg0cyAe5vQTAP
BtrV/NV8fgOZ9qjm0tUPcBV0BN/7+F+Yu4kjrlUdgRgyfo/mhIvFG0oyF22KsBpS
SHgTfbMw+3Gh4FW/w6STZ9tqMeBT2YplQrQys6E8IRCv/uJEzE2+LcZm6MrwMjvl
Mm8zy0vCnVk4i4svLNUhD4IEUJC0E8ig1NtxlrxCbpbo9mdJCFmU5ogMmHmUWliV
4LY+NBQoTbC4VoxlQOfWU+MoAXK007YvCxswZa4bptGCcCA791JC3pZPEp8gXEIE
HOZnwBWXRsE20ZHDzHwDl/g7ZCN6StNPbeeGIcP1/FZsOc6/Lgi5QtcoGfrSu4+6
TtETRMo7jDr6dE4Vx9N09hMdiSBFdQwSZCtuX3aH00pOv83ZZdlAJSZjK8gWkFzw
gO18aRp+xDygWKE1yWaAiJVQGvcfygQFjR6AaSMOykZ2bGWFXVvtyqqJL3G5t9kc
YJEmyZTv1os8iDocG/3Metj4wD6WuynbCEBSsNWoIKryoRzpScJo2t3ADZqe2m2r
owV9huoYElpPpTra5TN1OguiMr834/HGh7vln4esV/XxqSw3dA0jPoPeaYVtu7Ow
YCMfe9uQirx6tUaSPGP82YQ0YUm6wdH1Sg0JO4KHJ+1B7AQoCufBkGWyhoCQ7e3V
kyumijax+NyWGk775QuZUJtvNP1HLa5P/4l5mdfkdxTVbj2UXYW77UFDi9bP4Twq
7a31oppPzclPun3NY6CSqw7LBOhEtWncoty+bcrCJndXMZo2fMt2lA/MqpP+VVVO
6A4rAasgT4DKBXTjZyHef5GKw+YCnpfeYEOuMgMQ9lO6zyEUQWvGBZFTpUj8XdRl
/m/Rtp5VlFWHiO+0jrhcsni1yf19aaUWgUypN+N4q4stSoVPkyscAUQz1zc9rr3Z
n+YXVyHCfklJ76Gb9/wJdeL1emEjidZ3FkFLsWPrjXHUrTc3zdIHNgCEvfAX/ZYj
ZJbTkXrSIqraBDAqD/uU+8DAulCQfgOiKdQNAid8VzADpPuuAFRdNsNPBp/A60vb
RymBQ6QHPULfJxf3grk2oGxAvB7PhpFICU+rh2Ixkrndjctt0Z/kv6nEnsf5SySw
0MDycJNGvhhKeV7d+Y2c2bWFQ67yvkoHb1RqJe25huAk7wJii06LtifIxdvuHN3Q
fLTAJNa+XTk7JsVn6S4WGlt4pODRHSUt7vgWDEAVBazNy+10oF48pwIA/8jQOQ3r
i8lJKm3N/SOdlJBRPuRC0cJiux4lX3g49PHn1RyryhYhRJDN4qPXmipM+N6oG7XH
l3oTW6wV31VRpa7t1Q/uEXqCODC+Pa5YCEbdh5+X9k7htcHFOeSveLuTLcXe3o5U
EOyFKK9udBLzEOURFDx2zXlgXofKSx2bFDk+ypGEMD1WjlycVzAlii5Fh2cUrDET
vdYdMTskdEPAQOe3+HjfgTwlfRiwkIkODgz1NWUuPZGcSKXACAxd11t+Z+KSVl0O
RniDk/3noo+se5BLnUPtbHlQP6yL5XqYwJ6owS2ynp4zVlrgJS7glHHTOGtUiUSb
faI6TzkFt5ztVODuzpdLuu/8hMA6YJ1dKXOMicuYHsn1lAhpyORiNTrkFRpuvU0m
LWk9e/+4I29bgEvcmA1bVpKKaXDzA5aQSUhBYldiOr9IwwEkER/4CuhqHaJpm6ra
h9GbtZIFAVjwsem3NtrijZ3x1B+pX02XHlk8nY+PQYcqEtSkLa+4S0IyFgGSTglY
XkveI8/ekSa+K9yuuJPRibucZ0G/5zVJIn0UiZlk1OmwKEA0H0+XX9LdDmPDChMX
60dxy5UWf8E/7DN1d6hGjjkQcJB4SdowuFuaye1VIo4rk8ojcVx8OT2lrT19fd+6
B+IuD2stYSMnKJ3tzqsWoMe3wCxRKyowNmecEbm47XOH96T0eTKWv/42d6tiQA6+
ExPHSs4nkJEk8hGkzL6gVib2zBjjhiJ+kuIUnMYooPgh1GqOxw60YSPcrP8D/jil
HHqmgcs+GQSKzS3UZeLKoF+aLrQl1E2lPQjCpJm/P3scYaRF92tglJ0tKz7Byvbp
19eipA+OMpByheLaj9SxYqsnlC1lifkWEoBbXEUlWkLcvtR5d/1J4B8eY8grhmq2
llLtownHVmYQ2NBStEKi8UFbLj9ENyi4umQHQnF9rR28LeyklpF0XO6LWGqNrz4G
nt1r1Q/gB6eyxC+RBeJjNGWOYUS7GTP/lf/aNAbqyHickcMi3njkSuxSM6ysK7Mm
KkPOmAOTG/xwMHZj/ldTXD8bm4dFmmPCPKs/thCrozN0JTilV6QhAjLKs/ppiq4G
gA+Y8znVKLBzD3tWceNySbhsnNsGwDNwQJgonWYi6m9rYmkP5Twd9OqsOPZ+BNAy
N43ZMVrijKrux2Gb/9qo3pi53cdofvdE4+1/EGl0o5xcXSQpzD4KAJvLe+BNgL3r
GYHUFASeaCy6AqaKKMk9tAbbaPlQ0qHkrrxShtoK4rfBNwGzgFCp/jtmH9ACNb0F
nyOY2Ac9l1H92FoVWCLHpNbruFlHIgIOoIp3VtW9LM6eq7YUd65LPAZH4jOA0DN8
EYo9IvBRLq3ph+0ejGsWoCS98fzSmtuxUVgy7dktbsFqE85Hx7K94Ap0Rh53pmpw
zKX+BvYlHDsrKlspDB8/Y8j4SGS6KS8y2hQQd6TKfcMzdScXn3wxtpWnjBe4NwKw
PIwlZLMXpKFaci3w2+VUhEB1fQHe4gPaxfPhMR1QlZl6k9TsSQeSkQHXH2RkvcR+
fclM0sbwRmYwj+7arXmIG3Ls1JS42zNE+ch0dlffJpJ5U7Hs6lcRjBmELmHzaltF
wuCaoEL0YJ7TKm93YXWfu0KmrSmH0QA2lvZk8yRa5vnDhBnCpooQ2s89oY/7/U8m
F2VK7DigBrYuMFhDLrnU4c2SkZU6LpmClPvXU+NHquzEyGPwCrm6wxFLym/wzUWZ
fIv6tL7cdgarMV92XBXOrMJUowA583y5DtfsQkYTy1KeSonrxv1hEYF8pNcNAmpd
4Ea1MkvvUb4npgVEpFwGYL1D8WDSR2DuoFan5LW8MKYtrUn7fcvlx/J6+dJ1dmgf
sB0C207Hf4Wo/+UwSjPMEjBgNjts1msQflxzzRnetRrmGNinNymYBvKaFlzrilAY
rWqDiYMZEIDJpj50h4fZOUqTIOC6/n5Mhxkh8wEkw3OV+haQIBj2bzpYrc9XksHr
+TfTh+Lvtj+7Lksqc8CU3XD1ieK9TBWLZ6aUnVcbCDmpdzjosngWx8eQXWnxcSfa
HBAHGJ9DAeloN7AVQHwbGVl8SnOwohEgSsg0+AStKXW54gHqYMJ1/VnVFAbvL9s5
a6yqHckL/GQhQAUGmcTyMD+nBjnI3WWC+nGbXgYvESB4RY4X3ojjqsoiecbYmlv8
4XO9eiFtdMxWvNIPTccnr2/cIhyd8mOVh7rlF8kSZGSTwhMxEXXOgp70zPlXlTld
juRDCxw8OtAxeh2y2u4AWv8OUHOnMnAKA3bGfkyf1EsS6gMrooq/ABkPKFOnftV3
2rmlCcwp5A5X/1X9KX1f3A9m/STtcBQTLhvRBInB9yA7/kxZ4kz0qN3UTrqPDq4k
FJXRfV/dhJlKb43Pr0492HX2KrG5x/0HKHUxDAGV5LrSFPEqSwsThWI/rBr5lxT5
LRdKl+KADBLt7UOiPt+8U/Ltgs7NyJnbJSD+gk0IFXsaOXmbKIBo93zFmbu+sQt2
DDfLJSk8CH0NRCx30ihiYtsD9jJ8CdI71nGeBcQNEOzy5khWvImBZ5dLTlI+1UhL
ABxKNSmJrVa+sDPr//JSln45JGGWxbLdX8VueAHoHUx27NUL8TorZp5oSzHi7Od1
jT3TGlmOdtlddNFcPPUoCOf2q7RhzYP8rFamqBIkh+ZSUCsw3wlEynGYWYgpvtnO
ULfjJd0pcpvdH++bYm5VgiZ/1C0+Puy2GaBn8oHCqHI1IvXW72/Uqoje0lhb0i2U
WPafudP+zjHamTwaGvZPVV2JCI3/qot5TTWv0rIqIiLhdZM6N5AU9sBrFWK4auEP
vxrpBUmX4NtzjtIrNl4IoD7Wos/dWUA3P/XhL8+pyT1m9Dw8i3nA5y/EFTHWvNYN
RJYpe9wT83p1sHBs2QN/7wFfvJmk/ZUDvNuLdl8ZxpgC0n7zzAyG55RNVU30BEMJ
2Xvlo5P8jSwfvr/60sVvfAIFkQY57RIhFhslJro0xxYQ/XtVaRNEU4n3gK1AfhtU
+CKdloeu1B8cmqaEh2Za6k2Dcl1EgRaeFeNhKzbxq2RdeMl0vjvfACuJdtFE3OO0
0NGq82U8sFCkW01WjiqjNFaPnsu1UT2rqKZu58BCBAWev92Uykuyibf8c0edg4LG
iFLdI4c0TwKPt32o/+fYLJ+Vp03GBnaa6GBJfTCLYdCP7krXhIusMqq09y2nWGn9
TzjJM/D1TRVhoabK3RzRnnI428hwFn/daIMT3rxhh9Dso/cl0Qig9i6zc8i8Lm64
Q1SNFxP/Ooe61yvPyRwBdKOiB3o0w4Rn5RkTkLEel2ftyFmcEZh3NWf0ecUjZ6gU
V6xScdBlYJKxXMsIV9S5qhuq4W+LjdFnl49IVRSAvDrL03yJVuz4go/Bknp04VO4
2osJ95nwQRxp821zF9kz97Wwm/oGXjT+0zT/Ynu95jyXCV5SCimrVmbBk80P5Uks
twc63Uh6WWjjCVNHxdbSqJVyKypXYwGDFraAzT2LgKGJ8Wd+YkqxgB7vKb7lkTHB
lwfYW86bK/z6X3X/Z79nIkwPn6RCDdXFj+3VqdNlf58VmSiDbnsfBGfOU3ZpggX8
+xSRPINv2xaeR1935bZ194ItKY/JWUhTDo9Wr+akbQNz88J3xG+bB7S/FbD9Umwu
qg0i1cS189qZDzYy9GyFPjzs9LcxJeCMvPOMp3PhZd7lkmtgxOvMrkezZ2+8TObf
s7qE+wsWdmWQlC42LNUWiKWIy65gzJ03MTfG4N7+Pnm+zrMqJ4SFpW/oE1Hm5Fk8
7kPOXchvBQtUBEPmeTcIZHe0CYFVKsXpySgYqCs+jjNxYE0Ot6U+YmGZFiIYnIWU
7cO19Ax0GtnuCYTiv/nDCppsWGOBF76TKeD9R1++eJG2JG0U0K2Twn+Si1xMO7CZ
hVm1ZR8gcGdDWtVVzODOboXHGBf+P+lRmd5SRs704oyRkbaP7icyRmrpv7wPmW93
j6vTMA/o4wNUBM/6+OYQPmBBnH/X88g2rM1IYuMV4wH5PQJcKd7I9+7SUA8PQNQO
f8+VsoJiZnienGywwiYamA66aGkkCzkjJuN6mpSzR+Ohoh7a3kR8rdT+GvlqkNs+
SO9RTPJAUfT5IGbT5NCk6vLlCG75F/X6C7P3vaMIdjCKRA7RJCzkVUEFQLgMjTZR
fu2SyLZeP9e+hWQ9O05BElAX7kMwzD4be8k12kDEdvsl4l+d1n2jh6IPF/hrCCT1
MxucUJ0EsAOwBgjIdTLDNMtLnBGu/H9QDJHU00UN+Inl22hHNJfPogLmbbsm/ISS
W0oo0inSqrNS62WfUuACmIDBP8NNJ7YFt44ZRmEAbV7dJHPP1imBktXJMw5EjH/A
6wE7OdM7RK8WOY/4twco4udViIxytPa2m75gRAVueh19Q7pqlIs4EOw6cdXragoY
fwP/CEmKrepjTlDoNFC3kuAJuOuSVNED+zIoQXAynLPgNuGArPsKU+XAHH8aEIRj
DorWk6N9wDV3qNJu+1KYTLwfFPTndJ3z3/zNwBi4yWJ2oGbOzEmMaYGM9Ev1RxK0
2yMw2jUHXFKPnN7wiuhGkZWCrcfO4B97x8IibcWeRNpJUSMC3Tw7L4NVSPnOF/2n
EV1/PWI8iY2MFMl1yjejDG4wSLEbBe50GnbyiHlnSAAATLGsunIMJ4IVQjQkeIDe
EStCHRieAvBKL962xnnaM/dCcKEOPQNKPcaz0shhKZn3KzOdJl1h+ZrTKqEWEM2J
rHPIucGt04VsIgpS7eoXc/VjlTm8lsQG0k7Xt4EKZu2fZIhTLu3y+Gpl4rxFw2jS
Bc/qyySNnsp9DQQB/jF1tNtw6s83qVOvThD5RbmTUgVUyFpl9vYetvJIb7a93+jW
tyMk5YH5C03uUNV0P9ENxmpmY6DwZzS6z1T1MYBsGt/TxZr7OMxc+lyqUiEGDN85
5ETmpNA7UFHjJicMsnx0cdGFdS/1fXI4sTy1R04qvEgMfeJZqlwp9M0URikJC3H2
1A4y5Cq/yf/lWEldp9YzNkcrXJPui6MNT3Wz5ZfFgRdlljtpGXrYeJrdPcEX9SkK
XovqhqM5m8MkkyGs4UKtII4/8lqZFrLgl30SkvkVqFWn/PSCcmUrO2wU+FRLyCH0
Rj6+nGG0jczljQQy9utpVd1KxdFe6St40RTZkZq1VER/TbjeR1DLEX8VOZLpO0/L
19FIZcE4LixiAI0eM0W/X8YWcQGUsXx/LaTZ1skJso4Qq8R6k++tfddp7nodRovS
wOssE0D60NoZrAlKudoX3WlMyrDjGMTiTqnFBXWsw8atu/wNU9ZbBEdvb75oKy94
3zVkBP1Y+SWvmLvYrJMiDh0BM4B8ZLSVtEp+qPvz/ehadEWMlnvHY1ce8s8mzQAk
DCk7bYYiRkrq0YkoWJKNJkHyanPj15FtGuAbIlHIzgB9bABQ15I9s2XT3dq1nUab
gkunPuAuwJK41dN9acZRmSv8OcBnReL//ubeQPSg2MriDoABlHLbzyrv0YjM7yK1
sFXwkGlX0LEt1xkWeEYy096xViWBD4DaFm7bqHF2I9IlBn/Z1F5cSFZqsdqQzU4h
sIBgDeNzc/KiG7uIx5qxdEbBQ80EK+siIAJ+N9tKlkBLnVHsCjwV+g1aA4EgQnpa
XE3feOc2EmQcCb9mAnfejNdWCV/y/Dj1a9CLUSCvOjje4nZEw2g9251iAVuj6IJs
jJEp3JCRhEBGJ9CyPBnSM+SPFVWTlYYa4lUmHmfOwVwyM+/QWKlFlQs1sn7W+vy4
4ZxZOokeMWiuA5BCcRDK1a546mds1E9zlQqa+iz17G+i9hPR2miLCsx/hHl1Pqb0
NrOy/NWrz9rWtNXfj6aakpNf8L1+p06JfTjve6+SggudqWt1cMrPZ3L4QsFqRr1t
jDlZVMLeuEC9YdWENJZH+vD90ToGW4yq1ZwI5oaI16e3/LY3cmaMQ83vzR1ukpco
r9/jGRJf21hkWA88hbaYTs+lqwDYJLWSkVyM4FsxZJQpoGTiZ/zhH49Po4MdmAhw
WB57GckSXpz40qW3apOUve+a+cNjwfmmi/FvC3c+bqfH7tpdpjrItTbCxIxtsRTK
h12wpOM+QLlVKLg2SmpYNJNULu2T5MGSfvH616ARhDUzWEZ47T/8rP5IxK+JbSp/
ZRZYpjkOLmho43cXS8cEgIBlJ7VCRMkAplEXfgA7Hz4/4H6+2TPoQ0tI8gyjK/IE
5MKTSxE/78yQPd63dacUSP507ElcHU4Q9U0DxkPxgDMfSGKoCgmCAlxHr48/TYk0
SrHKtP+qAYJyhycqbL7HXirGxgLZrO7cc+n1XcnMKjdj32ud6W7bwRZ8viKB879F
hS0V6s0ahbAaNUBcwk3GQJ8vdkiI6cgMzbKiAwl+jXYrYOGJl9of1Yw6r7BU8V1m
dMOfQ56LQs7k74q+VJ00zuTvl/epNKQ7YFqhrzLrKrN/JFWfIeILkDER2UzT3xPC
j4K6/BqjyjBjqMnc4hO5G3oSm3dfiswnF6OURMBcBcZ8UOsPGTn55cE8IljH333l
ay94b7X5Boh288eDwpz5De0ZJiEtfaT3UDHHffAY4kp+YWhiATfZ7PKpNkgdbr4/
2Q+E33OxZofuNpilOnsa/8XP6BhkI2LcgbnCWJk9s57gLOFu6gd6MLMEcjc3MgGo
/8G7wiHEEkUaEKq1Dqv2BDTsSPwYpgU3AtnORGbn/F1jaV//ebQX6dnNNh3g3uNJ
Dj8K/O1mJKHApHkTYj9au9BvvqIhU82JxrqmGZR/l3P+ihGf5y3TbdV/vcGtuciS
O8+R4TtasBjfqngVctHn1y8uFoH3htL6A+cpaNw/Y1lFNMlK8I9eM5ydbOfZZGCv
D0lAexgnEERXG9p5VYOCd2ja/b0n6x3DsT4bNwn9PJxV8PSqQR5kOiJArVnhO/oj
/WUGPaC6zZDvHtqfiFSzUwIQEY5FyX4L6T4K7gd4LbKMBj8pTPH9Pz6OhDlUfXzm
IoCTjk2CYpBaT4F48YtYrm658Mx9LSUxikorKhDK2/8WuY2MoTcW/J607Jq6KF9y
pNJWFlL2dvZk8mj12xf2INHNbA/rEdyaY80mgJct/Qmj8gBAJO4ShPTGRpevzR/G
3rrq82sBPUVUZrlcQjNa9iFaCPLKkgCaPLe3hnozP4xaDGSNLFEVo8hz2Ef4zG8S
amo87ftHhpp2qEcENe1NmXwvXyc30qc7NA8vwiPdLpnrPaPzPEyyywqePitWKHJu
FJgkuYYZTqXvxQhJqT1XcKtm0OmWsOmVmspdCP4K55kfFF07336fTHaNv5O8za6S
BufIOsXC/OkzpTRdKbo31Nu8K5Yau+NIcAv8Fv665BNs6MHBSFovLgLaFtiVAVGm
bw4NGWr1lKxZ5DKm6C5x06fiOdkLsCyvJia5P5R9OFtWBM5evUEpPn/bR1giHhZ3
9NtXOYF/dW8Alsx7OoQtfZ/ws4OEhFlv3p2LTMfncmSLHOUJAx3Bm9kQlP/0vSQ8
DirRdFVXs2c5x+OnwVBVMovqUQCEsvH2Uycz9oUmqFDH2K+O7f1p6HNPSB5wEtTu
f2flkUwQ0LVmW3oOctBf7gY7AsvjMhHaCHXHZPZ6IJFcs1HMfzsDiSyoGAiOS7sO
04q14ZypINzeKHI8Cdly9zki6hiHAWXQpCY0VPStSa+L0cO+V27aljNnjUdP42Ux
yZf/rBFgbLbfRLGDkH1wMohOFv6/c2S5y7ykQMKP3YeTkiXyrM6U5wgvEGUxD5DK
q3GZZStnGTR82pE3D0GICoGTKJ7B/IsR30MZgxvoOVClL4SP8GQk++tcSSAumOPW
9JEyPa41yWnXsgQvmXyc/oqVHY3KucbHzU1pXAbkkqZA8mTFChgTV0DemlxmVKMC
l2yf9k//5VOnl3NTDfOVHsNZskU3asZQhIUR9xnlTdwrOzk2oyoQUmuyn9eE5gUy
9Oe6LoQjp85RUPVajAV8UsXrnREp6IHSDmz+nWrB44oDygq93x9+wSBCxeE+3bl5
GqZ92z0J4DFwo5hqCVYergjD5lJvp8VR1HLN+1bdTzLSpQW4mu+nq4fJBO25vEno
Kkm4wZXTYqMJAdLSI1rRjrgSdy+GKu9I1eCC0GySGiRYtqC/JTtQsgUGDOPIQJc4
EdutTD5LdIbvLkuV+5ZYQjIcjBSfDFXk9F6YVkYAhM9vvydjGa4jXO+By7hEafjG
VNacBH7s2hPkm37xVxxC17yuqtfdxp2ev87Qqx+hy0CCEurEkD2pqf46Np50zBlu
aCacQqjUSoGoWEmQRxssEQcYV4gZnxmNEqenSg/FYon17FdTym8mTvan1GX77wT6
39uRWOXSF8DwalvcW6yZnsQAd4XLv/DCMciCjUGjtCjwBWP2Zy2Oz9z2RTGTXjJ7
zr9AfItxg3EX6FtG33lXW9oEY09fhhTAaXR2XoM8ZskAsJ5ZKsvkN/d4j1hEmFWZ
pBjCb7ZKoliRGdLxp9aIhNq3Pa7wWp4tKAScDC5RWUC1Uks7bwnZ5X4xNzir68a7
c3N+xt+cpwmm1vNXq0d8vDy/csa6CRLrUhPG2twLmhIaI471OhCmGRJDulsJ5kHm
ZfEIY9Mv7c3ce+fLwFjg6gSm9ADxfolv/O1mMeHOqtXmnzI1QbYXkS++SNjhjKEK
FrLs3iKImwQj9h1mfLcAAY6K0FeMHYph7tOWqLNZT6abVW0khhtRoymc5WzaLE7n
64KasOsZ3b4nqzxZ2ThwzV/Ut2CXnUYVa6F3hHMzmaD3DwIerv1oVj2Zu/8Y608C
M+lEhddsH0mqQRfA715Hk/FgZAeJd7Lej99MyRwTS09S21CPKPnlzC9nJ+7riuKc
k90OWBUdLnD15JtxqAlA1M22F3Rn9q7mxBqIzq/UPXRk/Bx1YVjRJ1FNVPSKLwJw
inegztexGl/rERzXN0GaCxlspwdNmICBhi9l2thjC87e2RIBUijsugVdTeM1YtOD
vrnFSj7pRnCamKr8MziGMfDHIQGMt0BU8IYhBxffE1cIzcQeLaF5Y/p+z7d2Y4pP
fI16cjhFZ/2uZg4rtqH+mEpAymSt2bAPx6ExOBP5ORMs6/SnaZUAyHgPq3QETRQO
7yN/1/IZx6jW9bp62qJTxBMMo/q/QeNSo1dhvU8IMbJtaoXn/Vwya3Z7mR1P39Uq
na9sBuBeAGQTZF63XAlN/QIbGLMW0dQqiqCkWpJjOlfm18SutBRrXYRT1RfCWOgm
gW72rkETkSO7HCK1hYB1xoyE4e/epOQFNCG0dHQ5mYWiWHRzXEc8VGkspPmm7beA
KsQ+ytd/qffxTvnrgX0QgTIuOspljyRYpben70ooTTMs3OeD6GGLx9L/ZqhOe5rx
XNnKQu6scGYIfgIrxVzQmFG6wlGC6lkTcPQ732JUtULv1KYhA+p+0nl41BRVP9jw
3WLBMQmNqk4Wx2NlefRGVDKVsea4+VN1W6QlXUfmJizFtF26lgkqDg7hVW7RyZYd
Haxa77I16ikdNqYSUPBfPyufIK5391aSuO73NlAA6MVpZO3JOlDXzizoprg4s7FE
ylBsjDvXPRh/pMCwHGZS2i5VhVDlUHN+XwXn5FTKh4NapYjCtk80aS7b+LcgDzMm
fbn3uZ9mFs+M2qbSwJoSfMhtrlaDGn65zHJvbi+zxCbV8YuFS4NahwuMdpvqdElP
Iu6gPJVKXWVb4xrWkVlmrQD89jEsmdsiqJYaal+HX24lt38gvAse9KpjIMOtEIuq
7JfZUE9LmHyxZZhAy9lCyztdL+vgw5+WpGMVP/+fySnSfMGYHXyo7SmwEDxdoD+2
EunTaJ/akEz0US7UOjR+7hz4IX1eelNMguCRea24oV1lLK81/Vjhh0OJfLwTTX56
Z5NeF8WTVQ3tUFIYTC7HS1T+tWbrc6en5pbuZ3XFca0Le/JgOqU4eldRws4A3/Qa
Tw8+TSME3JbGDeasjpOIr/tQk6WCjva4JAj1bSLZr61NXY5NNVpoWNesDwAHjuI2
Hz93iXgUVXky0RCjV96ObXZ2rXU6LfWZp0R/I8QzILCipya2kxTc2CgmL/jO2uBN
qQp61TF0ct7rScymAVrkqW6D7oRngHBDXJtA3IcRG8ws1okWNH+zFNZXM1aNJzy0
6gnJ+Gqv34xko8fNY3CnqZf3zUjekdOQinIcBcx6YIAoi1RETNaYQ/qD1AmHCMaN
oCl1k5yTmbTBiA8CRrGLmpIJIjRhc7PxGgoFl8+i903rybxqP1Z/Dgzir1JOzDrH
a+Ev7IVN8AByoUEVRVG0nJvFVms+Sr+RB5wE7Eo+cKUa2cin4JCZXY4Gljvrgc9d
opl85r6NTuiAEner6fvUiANfNLrclJC9LazyjsB02C23QPZudj5PJoG9LDbSpug6
qbUXlpbTTAQh+UyyWvGewG81DIluAvYKIgzcd7heR0SoSU+4Ad2CevnhhIdbpVl0
YxTh8UIWeR6esWfgyMux62vVbnC8gt6vNDX3HSRAnBa2WMfvK8Hge6nNs4sBRb2r
jJEO6UhWk9TM0aRH0idwQLPlYtcxP17JttvHf9/cMaJe9sQ4OPcJOk0PKCeIX+Pr
fTkU6FnsTB3a1VPbesvssjQg5KviFuiMX5oXlo6GiNEi70GDK4YsIfkyoyjdUmie
u0ALUXNzgn9CNESO2DZrdEbGqidxwtHHLKoDYttpiTghHzX8QKXHC6D6M/cckZUY
P8D2gIYE1/IqCmqD48WOCTo9k3ZpOSvwRKiqZo++/hNMSE2rOFo3ACwQHGkmtRPG
W23A4fM62buhDLpSLdXI7MpMJ6iwriCL/GY6CFzMJkJ9gF9qmwB4QKSjlSHBo44s
ZnCXCgP5ufMWbjQs/vxZ3PJG1IC77fUQ3uwq6vLaRqeI1rxPCGYSc/9MOra2Jcmj
EQy8fBPp0vBJq1y3wvaD1TXR6R1BCQfdQhFgmRHoMhekNZPF4+alTxU9W+j6rVJr
ylQdIlJfiY6ER1f+VaT10dbDtwgc6Kdo33sgApCFsrrhkYfwCcAcmgW0TvWCJlMo
QW1f8srP/UB5hymgNPh7QX+oIl3bbzjALrZdXHuMhYXlbUow+6p4tnUFH4n98gM1
i8td05TX1KTmNRK4uz66N1qhXPke1eNm1WaZVGULe1Bw/SPuboB0PjnUC1EFiZfY
e3CXk4JlQANwKi3xL61QQt0hHS353/XgpRiHsy+LgpLOmjYtY164cxs/0oYj/30C
YrcUNDlG5hsJrrmLGlCs4KoLmszoPnhD3RoMJvmjr8/qAl94VPGbOlfgn7l49ce1
UXhdBaLCvbxM63jrTBqcWfXLIIMSTU5RSpwkm8PfTfC20Bjkrdp3f1nzfyw8Yqqn
z4OKXx/BQ7qILYiYIFI2c+8UMP+zyb59y9uXMNvsJOHon2PFOETf+J28PR1oT93d
RM/IzTxu1vxeMG/YIjse+7Ra072so+scO5RCynar0/nFRH5w2CtVAuQicKyWCCXl
7pcMy6/6CV2ilvWb/hFzpd4o56oX+nWigJQrop1TaceOSztTPo66l3G/qcO+RJsQ
lKRPj8VtXcNYkfM4HgpjwSusZAnskrx8q8NoJK5dNXWniSN+61ISqF1LMyNX+Alv
J9sA5EDQy+Gc+7NK+ZDzFdOvilL5DkZl33yCBHZTnupFTpIya2iVR5upVB342sAL
RmHGSYhJhzZx19uIqf9gW60MFB2pOtAsvgt/g7OGnAwMTxLIrB8ZPDaaM5UH6u07
FtR1OlszULbm5OwScla8plpd42vkQlNmY2nTiLxfIVGFMUtEytdOfckO5YbBCm50
toqpi2FIzvgggTgQbjfhHi70+tRGJW+tBEwg0ca58bvvzo2pyEdH3mWxA7J6+5Hk
uHNUc7Sv9kfTgq2yh7+MT71fputbE+r82FQr2Oq2FUv1HgOlXT0BUd/IXdXp8Z9M
lgqX/6JWCXzvM4gykzk+4oypQlMsmycozkADmE6HucWXTsXupr2AGdJ5XObcMhIS
Dvzq0u72GexeArqxJVnmzi4Hp6Lr8qlv+vNU/Ev0c56GYOrFQ+Y8Z29vzQ/5qOzw
lDgq6rjIsLtvxnsit0xyIscP9wr1MF56qxcEAk9lGC9VX7PPqBJGlQu1ijtoEBL/
VQyyIdMFOCxgv4NOMEB3wGdkavQF1+7hkPYMtIeBaZPbfNrz3CZjXXjA872gMXKJ
1TOCvTjRaZrMrp4t0Jx5mCXbGfN2C+o7zod5znseTq3u/tqKYYxEfOaRT5I9RCbT
c5/DqLB/PGgbCEvPwUMB3Pczr+AF5VgLTU0zPXV6gIU3O8ck9Qt9x8qfwDUwJJ68
v1EaMK0jyxCnQsU4QEgb010I/837w7RNGi0tWAsLhTrlNgUu+VqY1ybEgdJQEi3i
bQh8zese7IztkwQbWqzVuED5VwfSSKNr9Q7w+g1VinWQHYgkDPKgw4jDaiUCM8A1
3R0aqsPjL5rkS2IwipvoGU9EtY7D3cKsBPqbVD1D3EPd478qi34XpUoX8QZyYNSZ
hf7KrGon8yvfgX3OdMDASkSbkM6/mXSsE9qPsYXTnyT724Srw3ZSwJyPLVJDWyzO
JVT3wqSdYOvDjkVSSKKEX9bru0TtC3WT3Mc8cWqrPRQZoLaB895ArHramD4AWUV2
MKk5fIW7IMMBZ598G3pIvkgFHc4lmb4b/+ALCyIZvb0wMp94vqvFblNGMCEEAhg+
Q93J/GiCmo9bKCIy33Dje0ncT/uwQpSGkjZL+iVL1sHmjQPMT/pyGOwMq4tTZuZj
TJlDrs21nyZQJglbLtPoUOAm8X8tWr30TodHMwaeAMdvF3OL/99iZvVvuLaJaVYZ
GOURBS+EvPlITtb0Wj83kRtgMICTv99ojCDnHBmM0lrtDxr8jpiifE73QqPSxf/D
2HXFZIZ+4FjMsEolZBxvZWWQIiD43CXbw6NwJ8TZ1/MX9BhVFnTobcIdFM5Ywy6C
lUlts+WNZ9lu2KPUGFdP+rVMLbQFnP8wCIfQkcYIxkKQYOcK5x0DIM7DyVWyCwGi
PoKuzLhfoIJBe1kvauFU0Lqfc+nBJqL6i/zwyJb16zaB8D1mNvQQJe0EMPmoi7lN
VkJ4aBelIf84SJRRjn7/ob25DNjvd04Byg6OJU9GaEhX5kpxCxQot60bICg969uV
BRN3echxMqIC4r8W9GzFt/lSmCrm9MhQGix5bd5X8OrgYH6je7vlOIOBHgi0sgZB
urMygqRkwbczWnYmLpiwK8GySve5DPGBZubOmUK3fLaksE/njz7bRCyamjesMumd
7tlNC5LBZ4sdb6jWTa15Xej1PaNocME3XlE501IdUlrMGiY0dLOsdFZBiNeUhJQy
qoR2lIACQF0zsharbSJAjxuBtqy3s+F4jkEfoBv5ScmISHkcqEk+3XCFq86W5kZm
jKqf8w8Hap3l4KL+5kcP8ViiwG4JjL9A93JI6WhFtSCcW4D4ytorV1guhSsghshr
X6vSuKMPbReZi+tmB8TIKuzHgSLj0fO2TudX203TJgDevWlxN5b7nVT54BR74ClK
MM9SFdEL4NrHDnJBkIiRSVRKN6Trd+A6hdIJ7uGp/ZzHAgvxexHd2S9DNKwg43Fq
M6QKdNrGJYyE8/I96HPfBfqoDHUf3KBjJBTu8yKVLLEOLkfRULwnpfwJn9j33zV3
uZv1kEnG1aBuLS7xrecEEp/Zmp73I+lFZl3fLY1PytuKD8VFnBtQGuBa3AysHQNQ
HMITEix9tS+lprdPJpsEoIxJQyMptdi593OuiGnMy4SE6o89ZGC/LNGIIOzQpxt4
jggDBerFGFdHbR7oKhfkf1FPkKFdzJNIiM9xxr9A3osWQh5li+VdFwteTCfbuFfN
Dy0XJqWqYJQEqcadgfFvcQHw3g1Y0MzrXstgg4ipRVNzp86wfKXhdhCJfA/RdY3C
AHqowUgOQ4VAj8q1Axfif1QdFUixSpzAoomc9KuheqsdrtRDVj957t+k0FzAVkMJ
fs0o2KPczZgY3RRVWfQjUk0RGgm1n2QO7Nc1/pxi22M12m+Z9ka/IyMJV1vMM+c/
6BgusILtGJjx1b9IzDdvefqxPTP38RyOLd4tKRmArMy1lxb3FDUvR7RWXfSf6hRM
TJXZlDgNSh38KhF4ygLDSM6CivhDXN+prh0AdSdzHX0TR6Zp+7X8jSRVxEDW3uE4
K3H5fUeJUzUOw7evUuErUr9rMdSQs304pZE9oFVraNCrCEiXP3BrnImaelKDCWtp
yGWQg4PVLKiujN5hzsRKtHJplD3ihP6U0i6l/8+S89m9K9+4ciSn/lc05eNN/+Oo
bPfMZYbmjSgEOtL0c60jportZVJH2qyGwa0UALaByvEBtNLm3UNl9B6fF4q+huJS
YJVdZzc8YhgVpyHer3myOY63GE0g+9Cx8DAIyDM5MwxWjQXyBQOUSVXSqF5LZUCQ
wLI709U7kPyUZwInf5DHsDbEk4IDhtdSif/Usfhbj6nbkM8DxolgUkQZSbr1PfVY
b8a8BZrdVFrECCr3ueUyqSSAItnCXmmkcbnb7jZyxzwF8jHHv/B6YdM3r3OaNkUX
oYvLH0kRX3wl+7S+j2U/gla8L/PFC+fl4Sf2A5Yn/6vYNH8E5mrAiEtoitv2T+3t
jvn21A6lkqJQXCaMzuPen5mquBhACNX9DNpBKwfUGnhn3BC0yXhP2TiPVVAnMZNf
RvS+h3UiO5pRAj8HhIxP1GgnKDKX/Y48GjKa4zm0QO/+aE2Vgk4rH34LCcknvfS3
vhCm1cfsL1M924B8+tKhTgySQHFkiCYt02YMqJzKVdgFvnSMcMCa2mAiH4etzOoV
gdbBgfFwY5o8JakfIvleApo3XKCklHoihbn31IjIheMa42iLEo1pw7rzG/Xngyeo
vWR0zYY/u1VHvFVGEmGhZRKKuGTTOTioxao9Bi9MfuTllQcaqmPOrlK8Fbv0pURH
3cpPn96RDFUtSnVbypHYVVwmU6HJsjDTn4Qcjp3vPI/fmzD3b9Z3D4I4M0/dOiIc
0VP1SL9X56Z1lQiDOewpVdHtPQtIsMlf1nyfUPz7toEkPervUPuyLM6KdHYkp72Z
kHigRAos9xwPwJrCvxvdEt4ZaddTN/Lin+hfIvz0K9ypsCt7ufpJ+UZY13C0koXB
JcIh8YYpz5WjcKxJQNl1ln+IW2StLAeSyVN2eBNO8wAH7E6DhTaYZFSxhgJRBITK
BB+gMchlEHRhxmcnnkdYUwrCML36h6TGEtMXd0QA7r12KUHAQzYXqmMe4jljzxP0
J9uwgRZvRpIg0muG4Z/RCRbw1Scsw++QmP4hTYxiAzmhfxCHJ221ChfLZ2fbcV0p
cpBEs/NgUsiHAFy6xZHdsflII7ZTekADmy+Qq+i6wSuQZt28bpi5yGiujsIH36xm
9DwMKYP+FUPycjUVmmFOW7e+edy6KQfk0YTwoo9U+Sv/H8X+RNiGWJNyIQ6eGgEy
O7LogN/QTcX1sgqwGRz85Wyq+lIqb1rlvMefntx7jObqXqKRVkHpQs/C+UpvOmlb
o/ONoeVkhFg36ovcCsee0YMugzMg1LTReagf2QWnYlSaZ7INhX/OGkHf9sF9qAGl
Md1Axh1I0T4Rbs1kd1PGY8GvUfix1eAAtKvozGA94pKu2oHQpoYCCZNQnFdZzf4Q
Qf/mjNje4V2dqejMD9KOnY31rwkfR+dOvGQNWf2JJLxeN0IlvU92DC9alMSwtzTe
WZZ2ZuL+LRQWxV5xLFzzoROMGlrUGlXkyqFvFJOz8ifp/VHMOd4UR7eqHPdoGAbV
vvv0LYjiQ5c919SdzhM1/ymwITZE9gieO0OMSU/gmrArBGPVVjgDl0eluRdv76ny
n2OU02olfZB1MEOFUgcYs8CUXzd2z/qak63lNQ9bUcVR6KL9wtNa8cRVEn7FEsNM
L2LEiV1Rhig9uk9rxnqMiAHqRqmxW4KDaB86PF6PYQYiVdDPM6jEYvfswS1E6wYS
SI33gG3fCQnXYOI6fnwohW0Z0re68iBmM5mmC2B2auDtLxWtVTXcZWNRqcgPBKoM
DknJPphLqcGI3ZhyYQg+6lq1gAEokflWrbEgi5dz9EUw8/HfIfLXz2NkYUu7Hs1v
Mntl0acZJZxxfSV1ubSL+RyjPurfBa8kUgASot8rbDeOkcvMRTzavhAenUSYArJm
hmtaDWJ8jw2tHgujooAdLipegmAwLidntT3e/lhZqHdVlLVHSk/WQdHw4aP9LEHW
rIYlRx5xK71oxzlVDKvjlYB10JRGtYjJSe5YQDln9oWy58AulKgKnry1POPFjtLK
iTfF0bdzQjyP5bGfuifalWpWMINhnZ29oOW1d1bg43rpmjtnCYMkz1yNN4D9P9+z
T9tTSxaDIiXruvVZOQc9+3fRoviuRiZBGI5X6uBLfX2c40uVFKefGp4vAUHY7qE9
UIqr/iawVKwj5hULmuBizHcQdpYNkgo9ufuD60IHZ7L29ssej1Fa1Q2i26m2972Q
fE9bl8huP8ymhvmo1Pqsixv4rMWecSZssyPbJqcf976pJW29063sZSkpe53ozBg6
LxhZh4pvSwAY88lECHp8r0lUmy8mWqsVsdx92HMnC+8ofnKggG/xNTrxn5xEPxBf
80OJMA7pR4jTw+A90fABpKCUObd/pEVsL+MUGEAYKrEy9GviK8orlSD7BMxeBW8G
vp83HlT2VkmdGSaYnkCItaPqkzrxX51Fh23LD2por9Q16PTX9Y/Ohhyf88UlLF2P
iij08/YXpz4+RUN/lzdU3IAPPWHyzYY6dnkz/TpeVc+biP6g523PTaXPvIR9NjVS
PC/gh0BDOjDplfkNNxSUrLXl9+ySycqC9nNjow1ud/H76EvZEyE25r6Bwnhd4uTn
tlj4MLGoJazTdH9og7t6f22XTdc1RlH1tdTlY6H8e6I/WMCt3XPKnC9P61aaXcPB
+RRiyS7q1fpdbOv+jiX0DRbzhsoiwuaO65R3spp3rnkZaW2c4yaTNP+Wcl0fbcj+
8ZLuTcBVFdRtUiPn07db6qJMl01tAaDmBaCjX9vO/0qxFN/pdbzwzBuVTGB/oKvP
WiBgTxx3b0t/mc24OtA1apyzYsBLnW4a17j0jvHQnH+b8rZ0mrdZkhEQmzFPPd4Q
QLqCYkUzDYyoWfzOIcBvUv1aTENTbyjqen2Hqcs298FSoSYZ60Wi69Ykw6Fa21dW
BvZD7o5KHfzLAOJJqLddZISwXM8tEv8WmHrc9CEj+hSJIaVinWbe8omqGtkOB5LG
vhus4rPwu+W7xBuM9DcxhsfAQ8LIXSefRYRqFDrnS0yudymyA3OoGaprwhdE9DUI
UHMzvQpcP6/OFMrH5K8feWyPkMPgFltiFofOD1lJBv1jDevS41D75pavDJZ0i9Lv
WKBYgvRS1oZ5r7QSr2GKSR+AkS0OIdAcOU76gBMre+pZer2QHNljXiAyaC3rzkj3
w5uYoiff8OV+2b2ok+wS8RVLgrN/glBCIh0rKZ5rZgSess7IjC4dt1F5K4xjAMuA
6sCeK/XGxbAGRLPS2veLV/mgmn+xFSvCxYaRTVCmuCE1DJs5ICkCUztgliiRNl8X
FDqMUSZ0W8PR7cF6RTfUfa+t0Mw4zNC7jAYHfm1L8J/aBuNBjAIvJCMYmyZ2Dm6+
G+3vGL+yP5B5jQ88TJ/kYA67ynr8ZrDw+EXmjB91i+euyHYzlen8nOK1R+nWytJ3
yjjK+p1+E07wNllD71cPBY9xNsJHI14UQ4yz5Q6E1JOKm0MM99U+akMrAJJE+m8f
PIV1XuXR0ABULM/Z4utfd3v8aTUjLxs73DAOwuM4WtqcyspLPMghc0yMQ/zF9jKa
MssaCF2bqMSiqDzAOaBWTOjmquowRj/eD/hBPs6jR/ZTcRN3QdGErC12MuacTWjS
hxdPUB3f0WsomF0AqXLJ1IGMbpTmXdt5eZjgSGBr/wIctV5ED2UCNGT267UXHQCF
2rMU8fi3d2nkOe79j1XY7vhAhCVnccp3AWmij+LfakzD/Nt0tJ1jBrfyL1XJMaq8
+brnvZrMEo6A+u1pzNSqAW/qYRw2UfJtOdJ1PHD6JRc85dlk/nqyFsLEjjD91tmL
vquDPiH8eRTd5WC/MpGY3rm/la9pxl/hLxaOdNOIHucWM711bT4UwdmCJBtnsyvg
Bmxq6BeGzCF127PV/ErC49Z5QwaR7w5NewpPqQfiDs4Chz7t7sYKQ/CobnVT0Mud
DyQdvpPm505lJ8rxwUXZQydYSr0/c/fCJKwGIkVOJvc/i6WqRHY7hWK/BuBpbP8o
AwKY7N7wd4sieAymrF7JHSxQRLIGKl8fSjcHet4oEFMVuaQ4hMOak604NvVgajfq
5CkLKQ2Hm79E3hjOkmT2sQS4jlhXlW8JbFywh/Wy+aW3ZXHDf7DF3lafgQRcnEWK
goKEAePVeKTiqjtgmJ3nLnSJcTK0H/w0PAyha1S0aLXg/iJccJf6XqRqUK/RYSl6
mjWekniHQP511wt/otWKP4ezicuw4J45Slp4H8h0bIYknIp/KSRd2OHwdODYQeES
6jCtnvtKLH7v1ryk12Exkd88xnmiGI/k9g+fs2DUb4mah3QINTLo1Mu07nLTrxWQ
pHxX2Dv0slF1rGkT/iwzO1ZlI9gbQX+bre5TrHYn1ooBM90oN/A8Pj+mxswdBEd1
83MsxyHtf/YYL7WUXgwxPIdIxWfoQXG3mK178F14+Hf1iJ0E3IP+ALAPtaQDdyuD
1NjH1kWUeXTcElFS4ucPhd+7wbs3AkDirKB9tfusX9J9UJNJDrP1pP3DoPz0OS6o
eZsTeHrcR8nOBQ8ZNMRWCLNDE3eTQcJg8ZRlAv2wZdNQ2jxeDvFcUBHU5EXnFXGX
y71VgZnIXhdFr5kpcDwW3pGFm6AheqxzMkf0mLhJlZBS41W22pg+9L6/JfKuW97A
RUPb9VjUR5vGxKXu8HjFUE91lmeQEbQRBazLeFXfW38uhMoezwWiL+AnUthTCLoH
ErE62uWSMX9E1AvaPpLjuuMpLbdiIvj7vmBVj3Z6qHnnHNsUzNZgOmZO/kD82xEL
Qewb1kberiRl2/bNhHyVpw0SgFLkVDHaOdihsUB2hgTqILbBiQ+mVyRvQ1MfZVMf
D3EfEqIbT6o1adLhVrIIB4ba7lF/owS49bouPXXHGkhQgw1UcVdS4loZ4MUk/uTx
M0/zNbRqOLMvKDvdqvj90oF717RM6UvSAcp0j9Q6/yPd6g2opv5YpRsvj7lXQ7yx
jZp98gCbQOlX+vXpSnEGFNy5qrqDpDE/s8WfluIC/dEzojvIwftAGM/wmJwse3O8
oSsiRARn1L7VppL9T/tP2mJaBABpI+v1TAeyNx4fXUN/u2ETo4ysK8TuRS4we1VY
9raJv0hKIeXcWOBBic7A35vKRI8PdWJNjhCBEerSQMoEMOHBzuG6WDswMDE2ZkWq
yBN1QCAKH0msWjrrexqseawwyrZCVelAzKtc6JwutHp1kWVOOHZjq4FI6y9NndZ8
bm+Y4nJd+f0KEgnSpRrvQF579QWMjyVNbPStKTdKK59YIah2krdPHfru+/XxaxqH
zvLZbtN34AyBmFcObuYx7BK2qu5bzmXYRoD+fBcrqulaOsCGUMrsZmzG6D9Jo19s
NJyP5WF+K+V1I4TtxbRM7tlXriWsyGklNd3YejJh2/RITbQiNWPphblXbKIWBjcu
Xy6wBBXUz9nv+Aml03Oxyh7vFTOf9P6hKQy62az5hLfRFr/Ify2AtOlbntl5TPZz
gj4zNXyrA3lX+phtbFRQo4rOdDWdbfNAJc6bCFB2lmGsqU0kPqcBVgPNLWZLGPFP
ri73gJ+Blg0KeDRbvyHRqbPNp3UWPrMhGgsUOINkzXiMGu4A8FkfgHOCsOue9/Q4
NeegS64RL/B1DLJSRvqy2XGxF0QSttm+E7OP1Y5a1gElysbK3PX19HCArRpnYzKh
BNJQr+eL+HuJ1CaNmRW/qCfnPiGk+yxsRpRluWzcHg3VgyN4xljbWPW5YSWl3YPe
crixh5W1Nc+xi9In6N98t7Gijd5DLum7QKV56X5AqrV9fToWRJs6Hkqg2+ciV/UW
01BkQRJJCke7zKf0Gz4tn8+lluM6rFjqza5dpM7u1pz+aHO7oaPs+cF7LfkdYIHz
o+aqVrty8FNzWKNb4YlWJBoPXFiyhtkpmT8eNEU9lA3UVnszwEpFc2t8sUnDScNl
JmkJTwun57/xH+EYGuX7KZWVinFxnfcqx6IRzxaGWbdp6hBppp1dHeSqIkDtlBUY
gPqRr2KjfFsnc/q4ZFuFfhK+xZNKRNFoK8+AxGuRQu1lluqRI99HgxF9RUySD7PO
++bz1pDQiNS9U+ed9p0XugMA+iWAQAdefHM8hiFdvBRdaYdjgSIW0Jo/kbpbYP7x
jIy4bfXAiqJqzbsjBroie24LblaY9SHhvAYCWqqCl0Z/PpD7Kiz5o6DZxUNqEs+b
sb/1TL+eZT678qwqVHEDnADFtmQY2RS/jPW3d9cc/uWkDbd8n02FQn8T7MWCEIea
289yFiXcS/CaUJ+cwAcPz8mzfKP4do0iADc+ixwJyl+rFlqEOX6lk/rf3PtKfRbe
9BgxT3SymbODhPQ5nMm2r8D74xunymEsyzdurr6qUX14AwstxtYdKuGdkcBCnAdp
OT6eSZhHQpa1K6kSKnv660DFXoXAjl3yNTvssP4JdzxosyXU+h8COc8MbkKH6/Uv
hvWGrOKq3zARndNzNqpz6XLUNPATCbxZMWSJ7n27YqRyrT79dbbXKs3G1JVoQzSh
11ngdN14qg/8+eof0BUynsxZv4Cbfo+zyURSPmQRGVKu3GMndvJtooM/qPH0wtWo
SRllrlcQn+tKhYPVFlPR1piocnpCafYv3c0s5fU0oGS1c7600QoMF45RJ/S/yZ36
8hkQm0oB82VUrifbc8m2quzD9l7Ovs/zDMZFnseowr5WmbcEKFNhi+cWhR9E1/2R
subbI4JHELOv+RZ8HWbxEkW1WYwiKLqTgq/7hSBOL0AADAa1xYB9bMx+c8GGUfi7
meB6qY3UzU1aMy6AZxHldqCPieCGOkS/wymRrqMZdj3v0rAjv/D4Bwe5s23doNqm
iDuIktMlFPLlIy1RWA3bQhdORoVDkoxKq6GYK0lDbQqWEEOWNyZwwVCFIjjW9UFv
F13bP/lY/6W94ZUFo8zuDtnwBVlC4Eyem6RNgy0NuDGXLq0ePphCGovkeewovgiC
dgga2MG9wTFlT2sRY8or1XtLAlH3SIcywFweLx7KtQNZWEW9Vw1q6d02RG1xmH5N
KjMPur1EqFeM+tb11ivcc8BSe/nep7plXc2FYNTdWBpqplvpLu8KfNBDQ1UFg6F7
oWo/kzYGnyLAwg/0iQI7DJniB2uzzZRgc0bRElz56OfwMC6betNXVzegu9TZSNoz
lBAIsfckOdnc06mN11Fcx6xUDtSyZAxEJcXhKZgrBSLHRY87H7UIF8ir4oJl5wPj
+4yoF5pF4mYDt7Kf4l3D47JUvVmRfnxqGGOzrVZu6iEITbLBbMAL068eh4afPlC8
uR+1AN/auhxVrql6+r8CA9XBwpzHDA5N83sBTRBOly+00V9sIk1vnU6P6RJbNmWG
tMJ8kCGlkaDASY10EQ2EtjowzQdwckoBpQ73QEWClMSzmB3H8qH7wTsNUYmnTxcd
LeZ4QnCA1dhOKGt2QLidszbD6z7lquborIwuOUgMYVg6FIpZeVmpe2gxd/1yrmKQ
RqiH24ZQr+BQZFvR44QvFzMeRUqBBAsDAxb+SNdyH3IG2YNahFDDEJ6UbtGC3nzJ
e3C7y/SIEw9zOpdg7COQl2M01jDDew0s6ECr1ao+bsuKqRk2TWI4uQqiUiPZSUFN
V7MiJM+yYPNewexj5tx7Yvz54UVDpv7o6FoS13JzUzWGNmrpqXreLvmt041qR930
IblqovAPOrNuTCTibfpLo/jkniM+O6EiLiP5u90oXIUz3VVbSNVyXVewywLQIUyu
9i9M/Q4Vy/qqKik8Zk1XNwXOAz9Wmm+09OLW7xk5ksq0QNWhbfiZzYdEYZelD9kQ
BtMoN8UDXKw+0dWM6kkfdyom9F6ZVWoLhajQod2eVys7/rl57pg/bk4vggN+JzF+
t8YsQAwaBTCIhAzz4TruZCf0bfcTyvX2vlvBSLHIVpSAovAiTU38sj+zF/O6V64c
ffJuRJZuPOtlX7aVNFsOArCzwZYsc29qECBlaVdUAlvpyREHnQCCIdCyL9iAGs7/
MAkNE8BHNWVHiKmUgx30lvLRbqGMXVVjBK49afXlkjrg5HXrweD3yA3keZVEUlBt
t4JmW2KhGPzQR9C3QKObn0HWwu6aZYE+OCY8GZshSD4ihrlbOY9dYebxQcHxVxHK
LoPE9OBEins2TmBi5whT0mKN6Voaf+yufs/xS1BUoAO/+xqwDPXM0MBJuy096X7O
093Wc4Ww847ymOwnxziNgjBT/lfvBZ+VidOf97Rq6tnHKu13fK60UATmj/MV47YV
QKU95bESzhgUKnvpIRxmPdVQw8NKDKg8cZsfXCuqTKhJpYx/wSirfLTjV+3Y7h4w
XsLOegk5z9Cl5P1NrfLbOMBY+zZS7sWrtUSU5z0f8CLHhBE3gnyXjxauN3M3g7ha
EeHHUQB+hLQ1axTGxrGgdBgtXzT5ZwFvkSr3gEjmecd90v1RaDgqIXegFgBnVhho
12UzxARHIuD7Rg66dvxACUjNKCUsAwy6TgCWFvEIUxIsAZd29Y5JZe/l/g53o69i
+prOqt+iwFzZI7e84YL380YfpDHeHjlvUIZZMiwtpWxF+V9/NuVShN5ls8wBYljB
Q/6+lDX9lwlBPZCcCD51zeaq0tFS0WT6OCCHYIzqMpfi/Wh6MXOiEBNUZqktYOwE
+SpfxplR3W05neKgLsaClIwfLsVfv6xv6Vx0Y8L5n8rOy8hNOKdGZWTyUE6DV381
esnbfT8Fp6AJGIJgUSuXTNGWdcEo7Qn6sLLuVvJjrMvA2vVMDTmQERZPviuMpaYi
EsEW0tuFe3RwU8nLl5E/0pK4KVN58mbTnO1my8gbcnKNWW0/Ijh1xzQnmJOuCw6g
Nix0hk/bv3AIPSIMrXyjMl6RQRdc6YyDrWh6tvhDOjykxyEIjypW06fGr7QGwuk2
6mBUouNvwj2WJWd6wBUth08CL1kB5qjXvV97wLv7LhuFo/Ztn1YldxNXc+Dkwi1Z
NuetRN/vWQ67p1idEMZfci/66oHsZnULGEZUa3eoowiEWIhfDRYS9IZPYWTjab/P
nkU3lNmDRdO8qDd8zrwkhggbdw537jfYA9isdGOAyYclgnQ/q7GWV0zRIuViMuKG
cNZMXFMZI2ORIc6dVi2VUbEIm5AjZvnkFu+X7MZLchMc02mtVmJ6wF9yAbmgYOy0
H1IFZS7FZ7bOK6yl7H8O+ch9VRYTP6d7gjcoMCbl/kDzz4SCXOWjo5YRuyT1fnt9
xs4LJn2R77dL9UiTQC5CJBFZLwRCbe2JaqRa+nO2GXNLwzl40GjFITao9Ssu+ca4
ETc6B3kx4ef65yKWWfDSnX/hYVdthTiCmNFuap5zaVwiQfIs1s4f4ly6RiZ0lJ7H
hI9i+wGg7pxS2NrMBm0cjQa3vS3+XVRGGggWsEptK/M+qaIlB+SEUMKf2w1hhXhb
ZReIo2LxVO47x0k21uXCGAvf0hZysLNT4iN266fNQLirqquBbDEChdzcVZmR97bL
Tlk+vOq2hcWQjYkYqS9HqbnklKl/tSQV+qSKPbz6f8R48UK710hnQSe98hu4OL7+
PGlKmEjDpfVwlPXHAX4/YsNpcfQKB9Mex55aArDI5qkUQPmRAKN9h1POJrm853xD
uLgodB9OwygIEWsD7E0x0Xu5ufM3zU7kzGMOXDpS3TYW3iEcmTr1+rIFT1iGLtq9
MM3324Q/xkTC/HxHEej0qC0Ge72F21RNAnMfyhDjs8lZDZgzUCTPGMOVF5yfTON2
sL+FbY9rjRqavvART2MxPwvIgd8463DvMX1vUCIIaEKX5Bv5F0ZyyF/S9/+qa095
zn8Heoxf1DLA2XGi4U2nu1EItKHl7soEZQOFfMTqaPVyT9zb15N7wB8o5BWxz3M2
wHjBV2Mj0Ucg5MrJRntghyES/fni9OnOwu34kgkISC3juByIV+P64tiMsTWoY6F1
IwZPI9ch7kaWvHQF/DLYD5Q+wbQU9g+vMv4/wNKoKpYqvvjbip7U3Ba6CqJBcST1
kwskdc2hLl5JAILcUnHgGlKNFZa5N/KR1ACRZ80V4FJnAW1nAuErgvI546k93wb9
qPeo145FjA1sJaPZ0C//GG/FH+eZbVEkOkCLRdys5j9usAG506KeH8YJT1vripGw
lBc4Kll8epEw426Pjce+xuPZDqOPCDa/IactKqz/T9gGxROLCY17vyvG/ODoIVpK
58qmgLoKQvDcfu61UviI2SHwTfjZitesRS4f7upct35cHVW5w8fM2cpQR8gmDASa
FZAr0rspiBtraj1f/lVJ6n1fAMdYcnOp++3TRv/oiC90LzVV3/0Dl1TKGAj3UY2+
uhKrW7y7gSewRFgSGFmw+XUHlQRk/iNTnGuwPhe4FhnREmmQCTDay1LvJmIov3ge
AkpYGr5sONL1lvwv4OpQ+WJx36SCDhmW/cFdSNB5VS32iYM2BzsDQ3NEFbk3nFtx
tn7rKumFAmvsQBZDSjo+W8oeQ6hDyu33Xkwo0aHkMJXeQ/v8GbjDjDgTTsiPwv/7
7j2Ii7/F5D+gJhmT2YYx3peVp70h0ebOxI9wJXtV44o+hY/QcauESE0Dk+wfSkIp
D4bQpKGblooK7eendC6BnGqKpPMvIWPD+nsxwKIJZGZqD29obwTQ9xOl/b9qd/MP
99NaCT6ypZ14eJc5dP7CY6/29kiFpgeJO2oWji3rIBk4NiEfvqrPZ394802oUbrl
77kEzUh77orfth+AQMWMrqiNMVtl+v+Qg29QZ4tB2AcdzCXot3yVYV8gAFqW9LLA
wJJLLY0JU4EF8u+cpw8Pn+5BQ9oebNlIhXL0BmuhLZOD/djzy0JnPEV9N/c1BM83
5ysTEiJ+w58VowY4+ZAAb/OMm6lgPft8mum8Ls6jTNhYZGhqQYtrudoNg9TfVVqH
+ZJkWQutnMqzuJLlY0xqlek9CTQW6qeSmbjj1FKoTQmyRCmM15wxvaGV73p1N8Yy
Y8eysrt74etDT2xQe3L1DjecnVZEYQQe8i1jJgfXyJDGlKf7GrLduKM/tRUyKzsx
BNb5naWTErBVlSEnsLQ21DpWc9mhwhzDecp1xitkrL/hWhujC9O8QfZmAKoZyahh
ri6PtJc0OPnPntVL9v6upQlVnJVHQxIYDvZkmSmkqkNNXRCntjt8e51/ccYbPGSi
kw5pARVjR7sA7CYY6o0t3dGVmeM1CXEudOzhI9K2PX0bwhoILlvpo/nyZPqQ4EaA
9uxmUPyeBtnmH6uH9hGQdGRnhWCRH26hLi7BNrmly3NN7AGOzOYd98dtPry2/wbY
WDr2AErV7zSljERuPrxWosMIEtoEWuaoLtckJ4o2wO25fjgWBtCcWhvjhLhiULEW
MoZHAcL1n/Yc39xYf4oPtChisej6/TLyGDLNFfYp1bx34R96MPmGDRwmKaXeP1xP
r1f4ogj9ByUXunoJ2VXeppjRLiouOZrGL+FyZDmFPE1q/F5Ep3t8Qom9x7scNH20
Yc+ezaFYzqji0AuWlqyOisLUAHOrNd6xK8HGudJJAEZsyjwM/NtLBD9qNUJbWI4I
AXlNt2yz67WDrvtDoefga11L8m0AGosy4ObichSUDzFkd/3zCi8IkIFVd0kLtCwT
yZaC8hhXVjyjGlGnsSMK+tCZVITuUlHFaKUgMRDhX6W1OWR1/7h6xJXSXExk+xWM
J0ikovJWMdxP/bDXpEkPvd2Rdp3ZZTCre2A3lhVTJU4j1vZm8PS9NAusy8s9Nckn
jh+KcSqk1bRND+8Vw2duChTr81mHOgsz1XXRdZKgOHKMnJUGlReFRDon0dJHQbq1
Ef6Tq/FebDOJU1SodK6Zq7bSoItdhxi93vfgwxoysiUh7QK7CajTJVo5k14+qBnt
AbcadAQa3OH/4HevIROC+fOm/IBPcERmZBXAqnr+xEqqSqHAl+6/+7tz4uBtjxFP
Vs8raeNzHeQnpKXxE0bhY3Hb3KVm8WORR/5SkO+WF5uATL55p23DTUPB+dHmUSGX
UtHfLIOMt1Y8Oi2gp1g9A6bmvlJlkCH79yPp27nnC9fHJRg2YKdFigruBUypIJhU
pGst6qZM7cqlvJTv5QiraTVe/Mg2r6yZ17QxBnEm6R68LqXUzvleKTBhD2lUIUFl
s/wD+fvZXif3Z8H+UtAJ8S7nmji9ESAuNyTXto/09TGFc2UDbdR1DMM312fgacLZ
iIR1W/GGR9D15k0syheV0HiI3NAb7uYxADRtWzfMZraC8lSv/P04gnX4DBqhxla8
VACmymivzIvesFliefIUklLSOLM2EWX5sba7akX7sUwpu1Ph16J8SutXVGDjsGT3
idTNoyoaetDH+2y28d2frNCLxM0Gh6ZfUkECOWAnRWr7i4DGwZwNkrS/AboSy1cA
qS+FUVaR/EHwBV0WaTbK1CuiQkZgnf/Ahxb/bz9cyuf76O0bkW61C5NwfS/Y1sju
etWiqNoxx/AC9tIQuPxImvlnaLie68MkBKcjV/+hmVfuZVYZAzBjZGz9h3NCw+XI
v28CoDRkZ/pt3mSb7ozDysAmKFIyQOaTh99cs3CTHE0CKjXOR8zCeR6u9dW3nqVT
3BUY85F4Bp4QQoDsvS9F/zfcKZCltmqfXQ0Yu73YpX/KHiWBTuodsVwmOJ6twB9D
Dhhf9H8OVlB2D+krKW+pEP31MvCkqraT2+SAl5W6jIHMlb0A6is35mrQIrni7bMn
ONeqHU5odjVgC0ePWOIN44cAqxkY5QvAc0SKJs1em303SB0xC3efUqXqLEeSBK1x
WlrtEf9bJOmaVJ/WG8L4pbp1aW/X2jNNPRgETSFP6TC/oIDyAKZDiz9lhdKJ2RRl
aBYEEHfxcoh1aYXqoDgPgijEUD3sEpfGNB5NE02MRSxN8oLI4HEogM0AkA9mUuXg
67sBcoQ9bKVMOOgO3ClWmEj8eZVZkX4dCOfiSyChv0z5bW4KqyuO7gErdNCwTYti
t5/8hbSom85ImDsju/FTVXXtw3+HbWgeGTdd6ZgiOypICQ2vXVVmHXlOZapWeyFi
y6k8mAMMuuVB6SSDaos/sih1r/prsBJ9ieMOZA6jRjorrRU/bPZsd2/6JL0BJXiP
tnVkR4SowwXHStzJ75TOfkmj2BKE7bh/6ZctZsqolwzCBfbGXy+wYQyqsbUjfF2Q
fkGW9PJzMKp+sQpCmnSg5egoDjyxILL1rZL2EBlS55no0s6qraO8tLa8sgRWBo2k
fuprUis5Y6YH0ei3AV9Ld8souz4pYC7f9bUxjjqbs+ruuXwvyoul+RsP1ob923aq
V4ZLLkQaYS7I/O9LUQJh9qphRRfmzEKBbaaGvmKgBq0mPC3JnvYwWZ6I44VHgocq
NrkGt9D7Bh1g4Igtq38dElHN/BTaLDb+0z+ry/fJR/YOYGDaly/p6kgqp986l9fP
TL171RmtIVCQkmoISb7AyRXpOlW3qyjwUN/7poamyEnnfcVk2nTaol/njrV/YO0i
KJ6MNBGwm9oa6Fqm9NtI7+WraBbUA/CHkMmeUPhrqH2abHsFAZrBTpbLw2rTslMH
6hur3MLOH89JAetnCUvvv4z+zkc+go2CuDJTCo5jdPTy3pb8QU8hDRlDoV2EiOim
+Jc+6Z87O1u2I4dpCTCDFCiOGTY/qvRloxVhL+bl3uW4K9c4OFIlSf7g2r6ZtF+K
YGU5AHvmHY8+519R+gQzLZd7WtbV0J5Pi4pb7si06ssc/TZbDTzgxeSGPtZpWWzn
OLxKj013Q0qQy2wEJ2P3vMtxYJZ5N5Z55+V3S8hF0ZfUQKU6W5gG+7cjCM+GNj2T
/Fwj9W/JpClsEkHjVE47CQks4p3VToR884ibkYmVdqmoxOIcU+tngsQF0Y0Gdlxp
rl37bQEWycE1jecTNUMpdstqkU3yXW+dQ9/9GiZJtZ0rbatm//RXx8VcLjaIMExK
KIpmw8Vf49QsJ1AhqlkTJU3tJ6cvokTsCWs192jc7r8LRoUMvHiqhZzeUczj0Pqh
gSq8HmopVq1gMR0z9q774ShpEai97U6w30jLDc9t2S4cIEtPGioH1IRDLpEbLCjZ
EWR9GIKSxfMXJD/yo7QeKGFr+0HBAGrZ6qHB0huYZZ87AJ0nYwdwx3Hy6QjjrQuB
8ISvF7lxgA4dwB+PTtNKpPkilyfApDYhkxU7zi8prjv+Ui6Eo3PzcU1Ls+/tTIE6
AjTvJihhHT2Hd0Zao2/cNy+I38JGIIyDUYFL6JYU7zDT97LWFrC+D/Z+DbE8Tv8o
PzVVDIf9eeZ7eod0GmD9TZRm6+Xr7HXPLuT4eYInYGaj9SQcpoHh6c5bjJ+Y0zMy
9ja8jWG4QowMvoXtKSTv4CNetgLckJMYm5kA1O12+JZX9ixP/p091i/6HE2AkLha
HPawpjNfX8I93QP2CQ/RWBRAPksrbTNae+C1IBckB4UzuW20ILe5kml4UuBY0CDL
Ek3Y6Cb3r0KZarmHk0iqkaFL48aSKE9a4owModhH7l10KS0F87Ee6EgffRazt2Ku
cuGOGQrc++RdOXyXKZVWzREmY2CEMeSzPktaLIfPnG4LozQjZLmMTmwGiQS37tFU
YHlt7F3K7k9pmJzt5jZdSwpt4tA2jXb71CqVUo1KSRhozziBOGa9RF+qErfr+O9w
06m/Z7mkOrWqQkhxFuja+n1euDXPbWaFYN7h07InrusmRfvAgaF78/Pho+owpItP
yC+9JuWUYBl/1PjjxGmKEyOwf3NFf8yxZ8wgb9y9HxgzbFlmmoUzs6SusAtq/Q5X
Qs48chQqTCwyHwBPh8//MpKduC9s9medaUK1yG3aCOtGKUFzyFQaCPNJtcz9G6HW
jO/5+Jf/UQwn436uxN4xMinm2bz5JwvV/MJrlXBn/v80X8Tckjpp4xCeYjIoDNIl
uYKXoJzqTmNrHnG0xXRXrLBpJRotQQOq+l1b4Rnl1gBk9NCW4dr6KiLZA+R5ZM64
qYWbarQeFjmNemW3xefrRLsUYsA+k+cLLXmZmuoPBi8ATuCdxkUoNFI3gGjwnmuw
yRqv1bcsXKFpMAuqfUwmGKS3JgfmsPEWHu9Ppz476qRvFxmYoQ8eCmq5aW9teBmJ
RkN0SBUx48wvyD2UX1HEpAHuFdqQ7MwJgAX/9ouxQ+kvWj96p9puYDI6uNWF2R8q
1+KZuw/GsJpOD4oBMGHIwesPrXy0Pe8fUREdcWTTl7T14LPRZGqWHGDByvddA3LC
VE0pw2/QVrImXAAdzwBeoa1BiZoIW91v4hYf57B6YWMP8KyxALdI4+WwBrt3H70j
yZzLwX53kCj2K13Xs4ScDw1FX85SMXvfQZPu8RUynDyrkKNCHEV0zKlJySNHCTeq
YePwvx1vJuWOCWjdQc0aW4lQHOhlb8iTdLEm8vqBxAb3s2suN3WJzOqMg1239MNX
qYr+m4VX8kBq2JFn//eOWfQb3cdO8+oAP+BAekbWvE8imttcbGx957p5Y+9xp+vy
MOpdWfK/CEal4QqaLhHV71JHQ1cQQkKr1+Ds5qOXzRIk7rFT+Q5E07MQBi9z6WmC
UR+ytQV1wgTQjlPSqsHYMLBwtdYgJlxdd/cJqW3vM1MBn0tSze8Z6BqwPxCn0V1R
7IsmRa4clhA38MXd4WsO0eUKcraeZfRsHClL63BE4zI+0xPlTiyh+vdkbjjE2mVp
VQvL/NtH5ZjExrPdZWtdgEVf7xNmKPRvbTjUJIuXMkpLEKdJDdw7xkO902HOjQte
Hu+iwbXQVI5KuKsKz6pAMXRQqIfVY5Yfbvi36dMred/25aeOHJcZcxl3avaP7ZCF
1mPJaWyOdnojrlDcCt0Xfn3jW6GYrKctjTQdZJ4SJ2oIZjA+T/T83SuOKueAWGiU
GOa6T3ebLaeKl4WC+D1cZXII2LREXJAws4YSlf5yurnMua94fIwq0kxm7puXBCUt
FXppJd+GQllbZHASPAyXWd9MzxJGfUSVZfsaNZoGN56Prdvlmt5FyrGLr+UOLJgX
1eb4B/wIc6MpFZDCT1zhvYm+4uMgPm2lJVAM6anYr6ghtwHFUBAvY2syUg8TIn5Y
JyOVA7PQ0836/No8sujr5bxpbeoy4dUgJhDc/XpHcpbg39DTCwiGbOpEcAJXWNNd
msBNwXqMoZUJqY3ysnlx8DshdxSzTowIcv6D638GzNRrLY5EmSM7cm6iOzRUThZ6
UTKghqFbvzvFOELM9TEWkHYgzQtKgAdWCs7sKB8NZYmk7cvEO0E9i6mScMBEnps4
xLO6dYfqKRaqNfuflaPvlayRDaFqEahBb8zZ/2Eo2mKZhpnYRVItRSJmFywmi4aj
s5VIzUiLP5JIWNJt+r+OAWrOjskQTA7Wo9oAKSGXedB3yvQHUFNUPecIs3m5480C
wJVEZQMfJUKiXz8MhrkKvVChUx3g6bCGpCRjSSwDHcvkl/ns7GFwDccr+inlNOGA
YY8hzyErndUri4Exo808DlZcRlycIyAdhONsmV4bA2C+nt3etV/qdwR2nvsa7DVi
4cmo8Lxgd4INX+j8TQvwobQ4qhB9JwlVlhW1pf8c9l24v+paFHa/1ktPfq/sFj5v
X/4JL8ZiGPVhtMLEcr4VUfb7NnCa4PcFb35Ps4lVG0dGLK+pdhtDrnXEELAwkbmJ
5lE9Ei50VdZbysRHbkfpoHOM2qMBeSkLwQ+omQgLFslglm7D2ZKONbEuMZK8aMZ/
B/Khdt5iPqd/rqIGHW+z0MKql9IyLSRtBUl6COiv1iXaOxNL6f0oI4ljfXhvgtXB
YYpMZieLQ9XGaCw1MSN3qE/EVH9pXXlw96fu/qWZmeo8AGFAOxeFkXzZ/Q92Jd0V
GdzgHybY1PW9jEK8u1HkUpDwicJOaHTMPXZ7pQraW3sFb2LtakXYZQYUVIKZiS37
ws0CU3YKsPqtFxB1TWBea92QBJkEDZ4SMRm2hcuDeb2I+OaIzUywM1M7SmMmEvA9
oLMD6DySWQwT8arryxceZWy3XqUtxOhyM9QkFD6pc/okCwqlueUPYzLtLCQv0OIx
Q4t68lf9LtS4AP8m1Wj/Sw5jWvwUeFYWzIBfaGCXRuJ9oniw40aiMa9Tdles4MT6
QhA1P5alqrL0qI5BTHVcbJcYlLl8bbOKStbnI4aBKpn/28eS/iyql5D1ovIqnr/b
BAAZwZfPNPt+R62dt7HS48x3W+8m2Lr+h0rbyJDW+rMO2ivQ8kkJ/JEGJcBsZd9k
bfjGMVL5ir2HfIjrp1graYRLkaDrx7o1c1SOYXjot3mb3tmQSLlETc417CXZ9ixr
zULcpIXUUVhGBg4+80TuOxZXRALZgoTTP/ZlZiDVnK3Ayamf5ptE7+RPXJGswQUq
GCIKtkyQEmebJG5zs9EosHandR5NZIpLqdQ398xS5SY1egIo+8gh/4V6iM1zSpTO
VSNo6edcnzMBREleTSffUZm+U3BpjJa8UMYb3FfyniF+jN219/ZCJ+YrCf2vRJs4
Gl2m+DaP17NR2gmkLXF+ZlzCoip6rlv93xgwjhn41Y8dTpc9FP2+4qf9tcIzp6fg
OSWLwB6mzwR3Xpv8vCKtfOoLwAHOtuijz0v26TNZKcWBte1ytS6VXWZdSB7Yl/LL
6F9hCNKCkDpUbj30lxkxHUVMuQE0tfeMgCQ6qGlytZG6JnLq+Y2SsHNrI01VqjOg
4EAcczukxqV6sNlZjNoykEDsh5nSCTAWNYgYsn375TiNUye6eAQmQT1y24pgwtgz
VNKYcYV/E4ZWIVzGOAHiPTlLXdYW/hiz2ZyY2GxoQomAVO5CB30AqnFW4nQdl/O3
7UE8ToHBGgSviZFz/TcJtCVsPCJBpcIMid+iVV4udBONR2FBABHm2yeQnEGMkfNE
f/buAapYoqm5+udC00akMA4qM/FP1reoYE0y48zeI8a9U1U+bXyrgiEwMUMNp9A/
wjOH9feZlk1eiJqolV8w60yZohVSByJ6NmHHpf3RuYW8AGK/y7eFduuNBbpi7o/p
UkGa044BrIRHEhe//e9i5+nB3qfvZRGv7RtoKn3FihOIJtcwGBR0Ow7Y6PL1TGQa
5TiX0ca4W4dfg3AldLwTdcGRexdDr4+wiZOJN3cVsYfxLCXBXE1Rzlh/YkSj7iOq
ePEOzzT8Ut63N3oxyTD0MvYb5+bmY8hWkav94U411dosbdeSSPUFs6gMe47QOj6N
lyNDvWzTl2UWm244VNWCn62gWG+rozf2RnEFz8QAbH8ua8tPl3mvINBzC/CLH9Mj
OcXrM7ZSbEuko/0KjlZiBTL4sKJlT6Gn/mcBdUIgqfL/NCXcSLugEmdfAfnSN61F
KFZ/oEi94QEgjvi/f78bXdHZO9c2YrOGYdDuOks38Dqq6X+7lptM2U4QLPF7jGRI
FNXEvjfk0RVC60bdlBMnM166ZA98zuX86ldQNOQDkTz7CylsVP/hNG/QaeC5o1By
glOMO2ml59X4nFn87CwuHRw4BP8Yt1YIaAF1yAWxoEmirYylO6BOdVCWy+wq3Had
pF+ZHm5bHCm/BbtjvWW8G+xF9LRdAjJ8LiyRtfIUqB9Tc0tekkrcRHGyTc7+zFpX
nf+p1jXhjR8slPSZHWscSat/ZaLyuJzJu4ISFHJpubG3+woKs8LfhBkvdQOsz8Nr
J/qbOgZosGsZIZHAQnkAXRyERjxMA8yHf2WSOB3D7xBpEz2Q0arFp0bEj6QmeQXZ
KWOyLEViP1wrbz+1AMm2aIgOHQRjvlfmPVYN5+h8TgYXo+V+f1SgGAizaewdbn5u
5hc2AzwF9H96ezk0U4/4aN56ku/0SDDuo4Z7WmXeakIGwICRd7+J5ocXR7aiTGCG
NUWCDN7C9ccozZ4cwMMTx9s/jAJgTyAJhlZkdACieVH5IyRdt19a9Mv848hp6mpH
bTL1zCsVr7CdZ7MP1Cise5BDLiw3APIzXyMAnHY9dcFWBqH17X836MbL665Shlw1
55W8ZryjB/pHcdkiDbV+DWKGbIYE4+j1vXmULgU4tQTaFbSdlbSxhu7TCxGbwLI8
ptMHSVCQIqUdm5c+L8ugJKnFaE639IwQd8ex80A5O73EjFvtVB+/QYBMoj+F+luD
M+8oQagNfbXuftymCvtDHIRMQXlJ3jGqf7w6HM1RQ0a6rJE5NWUEBZkUsDSL3EqP
qQVQYekz+f7a2uWs4qGnxURL2fLaRr7ZGi6Syx3djtFNP4TJalwADh7boG9qb2sE
giCwc4rTqscruxBibxtxUHbRbRv0dqWycgWLN8hpwQC4trRnB5nKvOeYsh9ydQPG
4WXGxaSwLzZo6xDW2abh2hpzyAABC+a130s56Cln9muuObTItB+XP3p2XJXExqho
az8bNoZEvvKjI76WgWMfCfDnwiCzVNNb9CcJq/go1aYpBxW277aaCGQRPChLmsE1
kzGoNqZPDx8VnwFujYSTCyVA6FPuMdFE1FgriY3XpdTQBgHfyCP7PJDh4A0vv6s+
WGyC0Wx23SaCt4vXeVKBac9feytPde3hTzkloEJV1LloT2qctkrTfvKvF/+MtL22
pwyUJqfeAeimlbd8eYS4ICJVj+idJ11Pe+yeLbO8rJR72orV8YsPu7UawTWG1iuj
fy3IwyLVnWNpaUV25W3eglh6zMUcME0PaNya1iTKopwyRfG0+2tkclauTUTfZBfu
IBXpoaUx0Wl8zMfsj0tqDJg8PBJKnt4+XyXScv2Dg4DM730w7hcEc25WQ7w3JTqY
6SULDxjCOgtuigqwT1pJ3AOndMd6f+fVezE7Y4p9wtWwALREcUDoNrcE8jQABEmG
ioBGva4bE7wnoxhq7gpZgjFIOxuhC5PVykGwULuc5420N3C1dQBnLmbvMUHEgPcs
bShxg69/1P2tbShF3HEqMbACOSsEWfwZMhOIKnVyycoIrhsngkXmLOL9M7Zb/JIP
wX/ZRVelAcAH7KEJs9nDckCXb7/goI8vhewhFEBlYWwsfUBQQDx+oCaE/Hp2FphJ
kRBEgGJHWBD6QiDRz9I/XLR71f9KJcPnjxNtR6tZPMQDZmoHs8XfGGNSIOpD4UBf
43eesEwjB9ARLMdU5PUosnQ7u7HHaSvSxISBEyUKokW0ORQckXGdLG2HTNmULeMk
7/9Xnr34Q0OIoPDPrpenIagl0+z2nQR757PUKRBN1Dds8i0fwxyzbtsYAgVC0oxE
PT2MKtN9yiOeuhrErM4XKWWhQ+I0nOSz0xuTKRAQz9n7XJsTgaQ/nEqG4fu1Kozr
wPw2WbuYSFX0eec0kzCUr36VchwlxXg5x0u/6wipPfMmU9jcuKMCUVtJerw6QuAo
aDlOnUQrAeRUwa1V5RKMoyovkzpt+H7I7Cmm8REmx4ReEJClJejH69QGYvH50ZWA
sFiNzItb3Sgm47/qAhz8xoSEE3+X200J213YSGw3jqHvIzT0aArn+1FqGSIgNEZ4
4YdZR/Xqpd2Ey4oZvFm7rt2jpQ4ZY67DY6RJ9EJ1sg7NBWofR079i7vdtzvLnhxA
aWJsnjz9ajgdTSKw8WkPHcLrU47nKczpf0wd2U5Pm7dHKQzFAx/+bLfSJGby6Y5t
ajhR35pcarKdkJ5bCKuOrTstl5oqrIVN01DPPKsmqLDJINBxV7XlRmggQfaNbPy6
spEBMOk1IBxEY4nH6S89xFAnq3IEjLHDZnOWdwxArsmGOWwvVwwJT7LpYZ6rFsHN
01tUkEYUt7aq5WBVqv2QbU2yCOQrDvkp4qOQMYGYU8tL3FEfVGuwFlKAXZmjUdt7
X/TuC0OMnLJ0edakUpjASu7YF3aRDNzPzwANePH2NI4CxZvswDWaAI90vqCU/5sp
LUE7Rze9rEcyno/yg9OXFg62QyxsxsL83GuHRdYmyvSD6txAf7GBI4bSL0xDH3fG
T2lWagWAwIJLM+S8S421y+ycbZhqrTDdoiofbQ7qHuSZvcX3cblrFf4vqu1dUyE/
FCKSLi9guR2KjRv/mAc6fyep6T4aS1Rkj0PFaVahNIDuuIUWhJvjMOKg9iLlyQnk
lkaG0JlakFMCCp5+F6OJDE2Poi5zhu0kCNbGrgPQkgBTFQkameSO9naaku/QwP1T
zM1j6P9CiTa1OMmGfY1BOl6IY7fxFG/k7MvyJ7tiBIhEKs+G2htcMiNL6/rrJCgD
39SCfPLbHYP/M3B+s8PjJNiqAeaXghQkIVZppAW42KKMmqTIayo54iGfM/fzOJci
LxXUY3VYZLNk8EuV9OHJYipMK8zC6gJ0dvL8dOtNs25knvvdFaPf44LdbkeEXPcw
kUSKlrbhTRm8wmZT4fQ1ba5E/ITJg+fT6uz5Rvs/Utwd2FG7AHtjSRM7f/f1pucf
HckSvWDq6F/oghba9SYQrgX653aEM79oxBH9Zdr4AErbnkUfbdqEZ7kmp3EztWrJ
xSX0ETMHnyBMXH3eEBue/4guONUbSt6K8ogeLsrmWr6sGyL5MjSeq2sJ9L4e/Lav
sq5uu3/zF6wn3k1GHGRL8yD2igkffDFyeUxMJAxCorT5k2hYDhDr5oeRjEOPqohe
wlkn6n2ECgBQZq9LeiQ1+zwqFt5YvT6vby4wn/2/t1G/ugBPzQKkH9a8J8VMGzwi
/ba6e8Vw+kBs9Z1bSEc1imCXUAWe3IZ6ygPVc6dDYXS8/yWkfK7o4VkD4+j7zlNe
lC2dBn/ZvZ9JeACn+KvN4K2P4cHf6ckXzZ22z9qSWm+KxjAQQTqSPaWn8EK068qE
vQ+qg9NHYae0/2SqEwqYSFz3THYC1QsGVb1oEwU9iFWq0/4uUbKrCGzs/vpYN8vm
cfKR4yGTv14aNTwcYIyz4ybqlX2XiLYalUUOABGrUqAwgyTvXvRV2oGJRcwMq2bX
dt/AObYYeKiutwy/Te5eFM68wIMroFkFhsis2lVVV/55FBy86XPAQt/TXdJ3o/zA
1Q6Xj2C0VLiu07T2AUkTPKtTEk/RPiZYUds1d31jzCzJS7NLBVD2P2aQTW4MgCjM
uNQAcKiZu5RGJj0kdneQX+KBZhTHngbV7v1PbbATt7X8K2ssX67N4f3fx0e0SvNi
EKayHdZ/GwdekaI7D3AM9UGlYwpXMl6BfR/3XBlYDsc3kN6eHQn8V+E9fr22OPK4
3UFYS56i9SumDHv46EKBCvY08YaYZB2BCQzxy6XoxBdCZIgzDfjHAwfuSSBkwcw6
JoZeqOTZiqRzYFmnC5Fe1/Tkfi4SQSPmRk28q5kgbNUebY4+D4R2TfFmphVeHJXO
G8M+gVXWGVStgqmg2FnQL5joBvUPqL17WJhsTUP3Yd4AR3SFm7GDpuj/cokyKQOq
qVaPfu+0TiDRg39OzT77J+eAYGEDFA2y+sfmg4FippU5M3uhqPAuJj4awoJOIQme
1O5jL0UcYmVH5+3/064SMcxxCQYqudoQLG1CWXg8Wt34HfBtzmW9KTGc08Avjwub
ACALXHDqWB1QXGAu5IvTEXU9qe8Ms4cHkn89JXVHYTNAgaRP/ClF+vxpTvT4LHC0
fNhBJJ+7hjeg6isoWQMZ/1h3eKKKg37slVedHiJbjyGj5iAICRihoHN6mYnQ7i4l
uSOgzjnnVGnacSEQ1K3xKgYuu+6ltj2mBc2W8Y9+z3OvvlCGm/rtdk/YNL801IeA
9m6CVaFt9Ywm4Zsyb03jAnIOKFeEET0FZKP3FimRDoLq7ED8ZtbcCNEMYNKIfjOP
day35VEQVQxzGdK3gUvlXY5phHZnCx4ibOuLyTj6gMWyZjsMfnoymHcPBYEwXlg9
dN0y3TDBlhZDIUAoEsGyVjLxXsVgcZsTV6ACWHx6q6t/9ZsyCIvBBqDlDSKRZNFN
82ymB60scg+QiUwUjzoBWJLB9A7txNcit8JAq6AgoIBi+ydM9PxURdhIw5adVaX+
FPmPH8jqePTXATEdBPdJhOG094xXfSETGKGI2/njK9CiVNG6u8SzRhgydaSzIOFe
hfqa2eThELl/LOCZN+4vUR0JvXTLXC3xn/8NJt19OjbHK0YZB4fTXN6n0RBgcVnx
vHYNMDUjBLx2BsPGeiobMTA4CHBDL8u/lYT3VrJPIB0rLeuCIsqrP1tZVaNi/ByF
Gt4nJdq1oNXWsurk218oHWNSGDAi9GId6y0vgwTyk5ocfywv/t9EaXcDPYhJa3qh
BUAcd/Y9Ix1QNDcZBw0sMeNpXIvRiS4EzqK6cmYr0KSB3D1/d2+v27XCgW1sVomT
A0FPCaTuvwAdNs+zl16Vl974imUOt6BSiLCnlflevTmqjXVZYKMghyOD27okfby5
TtwVI5Eihqsc8dnHl3GElG/vW2sZcpTTV8l+W7r1LcEKPlGi4zcElLhTHo3OIDp1
0rO4Kt1s+gwmELqEawFRvQnGgNUFlf9lMUtkX2J0smGmlned9agt/VPfdx6hoD+L
67UF1lMnc/MoHujX/WdAU6bVmhRuR13RuJX45col3pktBMWvATcWojDHtB2aBMN+
ZGRD07CLRHjJzdzJvNYYaCV3B3wEfjL1UmfgzUU06l9taDHSramilAx7PH9WgSBw
XwvYyXri/B9t7qAF8Lrq8pL24zb0IfZHY79wLLSFe5Qdvtojw4oVsnw3uDomnyNJ
PK8Agmbqk5DvPR89/PBEsNcH9HlpLAbDJH/1KO4F49eYsumMG7qUIdqN4J1ltcoH
ZPtCN6YS49L8NTBWbeq9FH6+rwDw9qm2yyCtTyodpHBjL+7fq3nF6Wc1Hhc8dK/f
eHwfSr1ZIUfEalcQZUW19kK74rsW0qZiwNnapR3CRL3HHhOgPd/XF/cjiIbjgine
cer8xeOi/p7iNSOelOij2hgWqlS5ImdadWwDBc2qoZ5uXU3ZVhnt2gT/V4yqhzgc
yl63z8cMaPPBh3aKX32xpdN4Aw0PmN0/7i4eJKZLlVWv3MPTc/RQAH5sinFjNtf8
S8GOOZlnsuxU2A3CYPw8Gb3EVm5M6SMt4WtxdYZ7t4cbnimKwurngAo7vtFWZhX7
IOP1MvnQdysT/1h0dm94inoBBe3FptMbfsv3fitb51FWX5snEATGFbR+WqLkSE/F
chsAB+4zaTHg/rEPYmSDJMXVYtgf7dX7Lv2P1WaRhudriudbGtOgZNfil/wb84Ns
cdnOjU1obDec/pmhXD6p1A0qikdvNFBFGrBow+RVHwHtvCYhIUmFypBeX43g58j1
JIJYzF49Xjp5uRslwdwEdZgMuwPhpxTkIH7fBZzVMPIz+5CSaIXHaI7XrjiiQalN
7+nkt2BfS+9IyYBaYQ8vbPs4HLgPjdqCXaulL/+uP6iYNhYXInKCnsxvjaWcsGFx
YXTQ+MIbDuqfQJjeblo2uWVxmxJm6qXKd2tK/32F+IEFx2pErnT2zpEZn04fNgCh
ngPdXC947fskHOjNyF224xMzMcbiJuR7IFlNGHrRPzikE2y4TJHFiqwmoqzW/5nV
I0mUXUiq/+oYfL1menv3jhLeuKvtPc4JNO2wMCOzq1SevPiVn6jGKqMOXyAJ+QLd
mjRMVJQ6uqRawHsJVkdj+JjLK2HFhm3UCQT9K54rVdNLBzhcaHsoBuk1plgXB5FH
5+7I4k27UnQ3uOBGdup6HfpVb7ZrrFRMcHeMeqFI+deOckVUZ0HoEqDOIvCZ7Qid
dY9FB1+oLHOpPvi191h5rCiapgltfjtFoyV0yszB57gmIzjMTO3U9KlSJ4+Oxgc/
vIM4z53lXlr65e6ZFGFL11bGLjVMKelA+SbEdneJ+splZs6AnYPIMe4wYyE6BNyo
KXucQn93rod+U/VckTakpj0xBYBr68bqxF1rEckz97rCsY7PLqeyntnFPaYZ5IKS
kyfEQ4r/mNu/YbP4RMGMk/F3t3r0kYEiYlK9grrVmA3FTe5O6bzWyJWe+iNW+6QQ
OzesbovwEMBmkeGpI/UWjlcjReE9f7Kff4KVC6Vhc1I6/0GclD+cpFgiTxGBwgj0
Fw5Y1f8S19XQC2YhXwu+hTDb3oF61o2ZPJmRF2LQEMfdjOWXBlJfPQGV3dzi0zXL
c4aavumTltpjMgiSaNMtxSip1/0B5F4p5xWOQzT7pQuyjiERq3cDVIyXlmwhFSTL
Qifd5OLXH1GhQwGdH4YTxeuXUlD0pwyVsqopzTt9FKS/VGz+aTWrCfH+/OHOZzna
KX2CjHvtlOL9enDzHtVfGRjcRTH/Y271zZOMSx0uAMRDrMZi+Xqzj/XZHmIOB/fl
C9IYo6cXkjbcIDyleoB+NSUa89fdwGTipBc0eULeViIiCc3a4qpKhsHirIEJeYjV
lAQKf2rKUmARLN9Yd8FIkvNpQk+V3e4qoNmVdATDhhUwBoi0KCKvT+mtJnqDTsNV
QHlR9kz1QWlFM1rff8Pc6J74ugsFe2jjHGPppDnaIWSWHYpTxKmj6/t9zaXmxAYK
INkmQeRN/7Mgf0i0GiJzyhoW5V1MsbqmiyQ/BJ2Gmj9zgbbXfu4oF7c7wtJ2wLFc
C4onGm4JIvA/pfQj6fYwFa6HHZKLhirVEfegInqVTVPaEgP5++quZLgPc92IwjO7
5dyQwuf2sys+6P9/Hpxv6/8bHZnuKzyNRiDOH5hM+SeMMrJKlX2lCpxWyqtIsXLF
Z8Shml6ZYXlqYiWTF5W4n9NlsZ4O8bwQIr1F4DZVZgHLN6V1fHIy6/ye0d294CpK
GT8Rl6b2+px9BMF0ZbZMouWEorQZ6vd4SRjsUjllghiL6TZ65MMmgnThltWJTpxq
6rEVgFzfBOHHlj/KO/EVLOs5uBwywVSTuuq6tNq7fchzgHQ5Tsfy6dSw5T7PrVDI
1P3Ij4mX0Vah2xSVodSA+wGb2wR8H1nooxCnfqK3d/hSaSEGeZCurCNiLd6v/5lA
VGwuptNnjFQaWJKybeakgPTFpzplKoW4fUVH/MRGWzUPXCs3czv/pJqzdEGZOykT
qfu6JUiuM39xl/ShaqtXW2U55m+hdiO3ah/jcv7CDFcXeZPok0McQQSLyjD2L8Ji
EogtGqSEDzgkfsqOEG13rtxRkFY36WuL+Zw+mix82v5JEHD/Lymds5tQMqKNyj9Q
GCw+VX8ZytuZMJ6l7dDKlN+sr1sJQajkmse3Unae/3CIasNCGc8YQYU6kOhFzp+j
FWAiH+kqoozBYNLb9Gx7srDQ6pkJR8uMDWB41xpjM/5aReVpuZ76HIxuRs600abL
lrin1FaClJHtHFJJIblzGirapTdhYjMEeotxvWKf5aVchZlvGi16sjkeoaKfu6hZ
dZ10pW0WQC8dJLql7peZ2M3dDOfHKV2//Aen1Hw+6pOhJJcPZUaBDEpif2ewOOlp
N4RGhaOhj07R06CRQFDcrp1zOFFrpZJSeEnCxH8lt65hGPbTK/St1agdwF2i5wO7
H6ATahXxlP787jo+hYx+fwjx4h+g3L3vrIK/r6iEbr+6/+IsECVCEV7rp6mj9N3p
s6XWMwkvJCu3L/MlFzt5SuO3XtHHEMgExziaPDmRTTd7I4BXSRE9otmIbiDAOXJ4
+2MhedxwKjhLNkIVmcZ7DV0gRYYLxXGvyf3UPpO6Njb/pQCka0wNXWfDCMS/4Z84
nbQ9WlA6wb4q0SP62vZghMfS0jaV+eagMw5PS9ye2uPD+UfLhtI7/sHvOXSYgiRX
IwnR3yQ9zP5aG40cVk82kBgU6c5GVzurNzdLHfU/RpY2DUNPkTimJKr0oQmbzMq4
mcxlGfUJOnBFjqJ5m5j7OML6mTzJ2RI0UuwM199h+u0uiTUm3yNrd7bH/3IEqCJ/
ktzzwJIfM2WU51aPaiMI1jrg5ry3KC2hPv6Nj00w6JOO5w+BqfIZpcKvFva7P+79
3GXTGIbfl/TN6gTUArEpRReghLA9+Nz1X+L/dYjMeo8VPocSBAcIfSkD7rIAIWot
nDe4As9jiJzB+kACXUe1lNGsZiFqTUhH7trpNUhDt/zQe6QsTSRNNX4Cvy5uXQz5
FKuizEYx7DLseiwB4vaTK0b1HtaNPjUPX4XmRLcNob+2DEIYgeNIV+fZhvod28wq
gTSamds24Gll6CGuxEKad/eYuBNydiLtS3x7Le1zEuJOvQyqvuuxnkehgH3lElyy
OkPxG4tN1qrB6xLHy6jLVuVyHLm0qu3CWw2HJhmGDDJXSaB9Lt3m6j/TWt+dZEEA
zp/LY/t9Hf+3i8nzdiiuXJEfQ92m6Ae74T4XD8Kq+J81oI1FltRiK+F40WDuFpxT
KLPUbkTM70IpWxKejCgQu960EsPTDnUw/+kwGFsO9OURTa89WLYBUAL7WcyIfp6o
8n/EKXbCjxBumwNgYm8TMPtsdBFuAchnLA/e+PpHQgQcpQdq0AxRMuX/UG8/1UsO
er6VqIyVV8lWBO14HY9AjNWgcFTkazNwi49200j6v6PBtcbuwzsGQ5oiM7E9jnIC
KTiytue/OJEe2Q2ZQc9bFTMAQg8iGKjnxgNlX4RW3JrG2FyPhoRSC3j9pChfyAwA
m5pI/eQ55w9/x3YHkdhIe512P9RZs1n/78TPWwbAO1/Oj4Hkh8gKlVXAYA20a84B
YclePAYqG6zdKDgoOf0JXP4sjB/vuqTEHZpJePjoQKQeY27DM0gCp3Z3SGfyF+68
QLL/f4zI/aeY5lylVQ6qm7eamUHIMlVLg4SA5PSNvgsxJHVehxygYXm7tKGvGre6
EzS9Fo7MysNiqYSwt+0TCFrUkzA0PODXuF+Vqvfxj6ylLYdBpBfcCfQASeGz9f2k
O6eQZCtACies8PyD+kXxnD1bKjbAMhGRTf2vhu6YYHBIjaysO4vRJX9ip2Qej0Zz
fHeixIFjBwMHS41vArQBxY4B5TgCj5gTMlFr/fKB/C818FVlylP4qFjXAzRdz+sJ
IBvW8W2VJZmz9veRfxEu1B9WqaJqindHSe7pJGBi5CH48w8q2/ZfdrKwajjQb06W
fuytcnpbxDRaJJlgWPuQiYMBH8x/RmaD/d2kBfKhEU+O3TP10HR0a6lWuFweDQm7
Yw4hW9bFKRENAxeUmI2xbT2e/zDiWaz+X6rqMx6znsa67i575btQLdJyMgNVinqK
F8UIcZy9RgasW1NtFZJvPMRyDQ3HZa1xyyCxrBxh1XHKnnFTJHS+RHBFBsrhkVtL
1Vn9Ef6FIyzheZpviqtL+CMw4XsmvsvRMgSZLA3xW71NKN9hIIwnPFqoQv8/pWRU
d1pOfeRIrH5Xvhuh23MbR0t6lPWLf99Q/oQFXwv23lcFCysqyeaBAgN1X0KpebvJ
ah4ZYyq2zZG/A58MMr76W8/ioOfg+ysg4cp2aQwD9PSFBjAL8Zvo2uNEnaSh9KYG
p0C70hnXrD9munwZga8K6d+9c4vh/iRlhRFohHRNLnqmbkPBAV86bjoydJKyGTst
EZjlshnRj5GMuSIxG6ci8OZ4cLs6hLq8blaqO0wlrQQln+3k/E+HS69teOKbwrKt
45QeQ9cXWueeE9MJaMjkdSOy4LsHR6Uy7CcT5mcNRdGbz/kmkszMYqYY6BTRJ9p7
Hq3/MHLxjYokiJynmZ9Ev38DqWt70WM0S3OtikC2yBrAqWvLKJKT0OyyJA+bDAhc
D8ulYQwTO+vszV7GAs3eYwabHUp7aU0aRckH7hTr9UuiD2Uj65Kv8uI97qq5MVfp
qOkMC/EKT41y1a9iqIeF0KQRsmq6RhOc8GZfyor3BeLT/bVI2sKvgNkWS6WUqljv
lG2USuSayJyzKSUPkvm1k0UKzH/wjq1/sccbd772OQW/xnlkxWXN5N4MuFaWxrSS
d26ztS1Ht7quiLVLNprWqbwHen0iHC/945PwG/E+MKKp+a6fPAoBbE6E/3G2PnEv
ow2FwAU8LH5cw9yK4LgBCYgqfgdui7a/BRkng0HNyuunhRxQr6qsV8gESrwg0ZDc
GRKujusFfaf+s0CNR333mAICeTX682EdW43vKTZAC7Od3T1nTHQO1RbxYDuKwaaU
8vJz8lRYcbjZJIx/ci6QYtyAb24ZYs/ULkLLwD1LjmqGhWrQmgcJZRugBetDFGDR
yn0CVyh6nT3+14CrqHyG+jDA86sgMaWvCq0gsE0YQcx0/fXmTT9LEcpiqruTMulQ
f5LCx4HstsBN8iTkd9muQ2Fon3D7bDykeizEifGtfOYChbHK0zL1JY5oEpyomToo
soyD3zH5LE9kROFQl+099ZNyuZy4DxioVgOXP9Jumtn5EGdzh7JPjUMPgxiNf2T5
Xha/4JEAHlOR+z2SJ9DH9oU3Vj0yaThW2foyZ0zRB2pBlmF96u6HM2Ktbr8bUJub
V/Q6rGEmvA3gvXDS1LBeEs9IdW+D16r0gmrJyPeYLtbSFQHsTyV4Jhn2LtcQKJdc
I5tSB3JLllNFYgdu2belnt/VKYQ+fL8HUhxlD71CupbsAKFaTwI6AgLvaCH/rViv
MGyVHkq3WysUqUvPDAagSEBQ47J10He3dH4SbOE25MS8vWMwQEVwOZL/dqHE4KrL
bfQJFCBdLJO7HNYBP+U0alOAlvfgfvJC1jKv2E7TdW55gpb0X2myOwjCUioGzDDA
8lAx9wPt96VKWMwL2pvTl/w8bOxA/tKO4snxqh4RztKphuGp1yc/hYsdpeydEURs
6hXFhWdEzmwd5oEVKs7qsGuSSOBgOpXcX/1tuVBEEesY81YaKgPOYYY/uwYj5/6P
I6VLjfNjsxSQgHz3T1Y03Fz6686nfDC+tjcQ0Mdq/na2MpiAmI7SYAFpD9WkGzH3
fhvL+JM670BfkmMrBcPFTu9wHjmlpnpG/JR24ikXoHBOlsLsSFATR04Q2Egp4Dtu
Sd6uxF4MooTWV2uVOLg78B9IXuWjgkSOiQf+HpwdYwr27Bsak9vq7wfDGCBRrrFZ
yI4n/4AXqjuh3Gc6P63KrGvAlCW9FL/pcrTICJY/LiCkgJ3N9evulNOYCGM6EUzb
puaX+3A2Hhy9+pbxRaXp90ITrkLN8BzSkbvqOBp+7lz6vo0kD0L8s1zlG2OwlJ+0
1G9SG+GJR0AbNsDMspKUcR/eLlZa7pZa64cFCcn+PucFxBMbQiAHKHVnES4rZ9Aq
UQqaeN1A3T6YW9e8A4dTM1CSj+izLdlR6smUobbCz3BAlhFWh44ob0Gfm5qi+/SA
I8MarKMA9flVMP3XTgC064MdzXPxXqb2fpjTQT/KbarIjFsCLd21JkMJFW7B6Y2s
kSFLSbuQMAEd6TeHvwY5o+aRpQMr3Vc4UTUXoggWcG7wMs11jRUvhm4p1J48iPib
eTqYNURG/ZSYubVEUjg7mdUQ1si898EQrzyk1hD3ex9d9giSOg+o/CBB9gs0G691
/aB+/1irMtHApetg1XuY6gDHYvWrsYXCOv2VC3B8p/N8a5EHdropMHjVvdrZzR2s
CIxkHaAloVeiA0wJgbj3NArS+EAWIZWr3BwG6M8LhfJwF4luXD1ln6ozCvuFFXuD
GWGAM9/HoTwnPlFB+xUh+UUxZWF6BuJE+/qUCNCvDcO1UyJHDKw0RB/rByW//V9X
H7c584wiLsSH6Fv49U+AEW2YcEEWp8vVESQNYIGmaUZKyJNqjNrPsFy7f4PgsJ6p
rrIJitNZ0cFgh3ytJqwDZek01XMeTcANXzR4RH7EP+qwxGLiq6J2CCyn6F0HZTHB
9+g+tlOi7kOZZ8PIQWG0M+h/F2eLHje9u+BUgIBOgvPFcDTv6k8U5Ovk9YxYfgwj
M/Kyj3RtTVklliJe21ybUevsdjgj8HusJpkrF/9TMD7jpksurCvV27nIM7otaGEI
4vxOyuXIfXae/2i7nZFlzAU/7jY2BvsyicqJodtF18Asm5pP3MiWxovFSRAXIOE9
cHt8SJPx4+NgUce8PQdapBSvzBEO7O782418R44XvuL1M6yvpUWbxnfWZpve3eM5
4UZB0S0Zfp6NbtWJOwWLA1XwXDXDCkLYPukJsbtsajYuNWHH69sFLj20xKj6uYXb
gjpRgiohsvFLW/mqQOUVitpEMA3EGEYlgVke6NeXHQPE12IzQooetujqNbvX2qy3
u0eXPX3gZWDX3S6yPsr7qFm2oEiK7kaM4T3mEXunjt5Sy/qOCONy0Epxp/X3NC9q
Imzy4hvWyHc/8o+rIvGTu9VYL5Br9Udbl2nndYqOyUlB4vl7dsDaI8zi6v5+Ghy3
SX451+37mtY1JnLcnpKWXW6Z3guZJoGpfgsDqJojScBVGOjSqjJgFspdNA9XwjdL
35tMAySbGfWG7MYE4NYbX8hzet5zFgMc1rlVUTj20QeroDgd65RASfrxe0Zhmzu8
A7N1cK8gw+fvMgNowd12bJTQV7Jrd2gCMUb5PZu/1H0px1dtEFrG5j2qNKBfcpFN
b23SlDV8jHMjsMyVq6S1LBXWWcwSSHCl+fPwHWMVazQk5jbSRKK9AFRqaIltqUX2
7AqpAGe2pDiDHvHrzkdvNvcVbSRcPuNYi2Rn5NhRKiGAQMY+SfE5ndFdMjkzMQwN
w4zjqSy7IRe8i0Wq9/JCN69tNDOL6R7a6rDuew1Q/VUO1SzVrn/9DiVDde/BrTfr
5iFfrV+furhCaFaJnfybEWAloTX25Z2Cf0Nbl1Z29YBOik+ro+KKZA8lRbIf+fZH
R4wLprJ39zVdxWSfsN+bXYvdLbRT8C8/cr233xNJyg5LySxK26btebjGovWiuMKb
ClTaSGVw0DJwvOhkHKKqHmw7J6DWVEEbjpYM0IKk0Tx/w9b3BDxyEZ4sUpDlsz9C
aiD4Zu1aS6wWIuxLHSkEu7tOPGcOtsGNJKkrvkKuXaTFmC/6P9Hmhc2f+5oXvX2M
nWXKYi7uRGnUlly6smYTI6JqWAMzJRzhZBqMJSP/Yi5Cvr3obJiQmdKNMoAmL4zM
0+gsLk9K5VpICjUAKk5fi/CGJMy/u0J84W5bLCrOTUNp6wE04VJxVuW2iC6cyMCQ
Bxiky9Ox1vjdaX2+sF2vafitVa4iguojARXZmOJGhy3ONs820Kuv2zcu6HzZCd9d
x4N/ItSqBpYr2GMkEHCjMOBHLz6BAPH7AXm2D427qU6TOc1CdR8Pp1Lzaf/RV8y/
avDG8Kqy2cHfgHmJ+mUInAzKGFDzVXPHuxwtM6KoKVGT9HABuYq1Itr9snD9MmLV
B6bhJFVPaPi/dfZX0l6Z/K9AiaMVk5hqYNhj5DR37fL08fP9+xXSgWZx1XyzU3zx
648wRsXA573fXMOPzI0D0np7B6bm3gWketVjFGeQV5BVK7HEPtjQkv88EFjbZvEV
c/GWqa1YSImaWF4zpNHPenPZ0dWKrf6cOYRKB0h6pSeM1QkIQr+X9sBfJWZOwLyN
ya6/Fgy1vcG/p5gmjwhj+W8JIBIzM9xTu060vdxoEQeYEcOxeozCYNpbpYHRiPJm
TxPoc1Jv4x+jaCob6iY2OQGnPdone0MbuSyTOuJ+afCaIyDSNqST5DNjD7BGXg1l
yOpN/haMWkPfvGIHNAMLgCopzJtDB7oyfhlZzbh5jUdca36b5lvumTC3y+tLxkOp
Exq7AcGz5xXRQNPoj9tJDHCtkYG39ib5u3MQ2LCkimYxvzKZeqHvlVtrRmDS3+jT
496iVZHHU54rPhkbTrMPLksuVQmSi4cFG7m/qXWuoxbHlulKKC3KGMWpE2j7l4mY
1pL7MZVEq6V//tRJH0o8MOb7r5tDQpj9YbvoytB5G+46QxF4AT59N3EdjYJc4pOS
Do7dq54lsUq4d/VMtPrrj9EOxO2hXj3o6l8QHIOWhv8qVf++afWqEMyBIVBynldT
FzjD9C9MrYejpwKYDaqnLQSIpCppUZJHBzUw4lsTzfnfcHKGLYk/h6HFM2jPLYLh
OwuOnOUjlk5G2y5s+Hdz7PAty3nmAm/zGrtdJawX2bEuZzhv1SlADushUbYSs+3r
w0oG9bJgY9wsRA/uCf9L7RubqE3UrAVaow9O486ASxt4wq72V4QJYhmREka+eFNU
fI7iqEKEhzY+AcospcSaB/iidxNu0wVPaEDDLm7NEb5023eB8RBnN3kemP1Dh/oS
UzYlexL5EJ7noR4Ql01FGOBJNVAjylLHj+m+AoWs/BK+GCHJGIqK6M7YLashLGoN
nEoYedtXDupO+r/D+5KTnQfB7bptcCWlLGcUITFjfFiQ2CJhNCofakQ9ibu35b9c
ML8ax8pidZiyFaIWnolz7B/WsQdhYmlzQ91fPQzeFuMTo3vxRDTJtxxvmJT/vvxb
Vqc4/vFUjyQbC9J+WhUf+2SuwlYrzEoNYIJ6msCcz2axQzEOOe3h/5LQ6wJr9UkK
B3CgtUKl/a67n577tXpn++Rl0hSpPCKwWsJgztD6/epLYboI4uPoGPMu0dPA6lNK
kkpExfe+kky3povSJkyisRnpSSJFyDsWB+sHPfoVBoKQj65duTEOSlHlfex5wARI
JmAWm0yt9uD9xZNBu5NX6xnC/gmTBLH3Mm8iuYJJiOzOklRgonDUcDBztUfhgFNr
iTtQY97dA0GpVr9h3sIsyRG0MuOegMOZvLrFytdWG8c+mxkNL4f0XWN8LWh2TwKW
qm4VLWszj+7hDYPtJcrYI6vyrycLuwECY54Tx2dkNwME5+qLIlhJCXnePtFZrAnQ
9pHvyZ79K4KIDA1W5LIraXdjEbKz9FieCActV/RyPPi5t+MddryYt5LRtQOsC4mN
R6xvr+XB/zmXY9EsEhJM8B/lA3HdvQ3bQl4JaaUlvGkTE+827OtW68serpzRzGzc
EGBxjqjcy/uYdhHQ/aAp6wa9DGzDfX/YJXKPk8vbLIgqh0tYuFsuFtcFX4Pc1aKN
c0H6uPmGg5gqGnXAGBLvyyJdJogfHWZtKOpFNRHmLJHXk00u1zYmhVBz8UkNwKsL
OWlRuS54mMaU7AP6kF6zVeJG6XeMpNz263+Jbsg/rmuUmX+vQ9pDWlrk+y7381Ib
trXI3BmxVFgGv5spWahD7GD4DwvZeSo3a+hYP6D/Ca9gQa3DwDj6TkORM+5xyj4I
uxatyhlvH1vLRoTU97195CuTEmv8Xln1yhKtvjHm5sz7Abvu+X3DKvQPHkYPAJrl
KCKxkj17X59/7Kuw9U97oYi6FrVEhnSpr6ZgLdYepGWP7pVlosgmxHX3XkBr47SL
sM8BzT0HBsqs7OXeRYRusHwgyZG5n+xw17lTwoTNSJlqtIlqy1+X3clYLzVTQZR1
/hOOI6zSt6zUJIAGbV5dNr6RCVDjKsy2cLxFiFWAxX8spNPbRuWU3MoxgjCb4cwf
dFoYZbenIiWhXloUDej4e4tlmWATn22uk7e40l97JkUi+BWCfSO8lik7TdyEciqZ
cnK31u5v/uh4u9fzFm+mEdMA39j9PPHZrxAOvL+YZmy5a+H3HAHmrdwmh4omc9Cj
C920+GKRbk7ZiTpRZB3SWYJ1qAqE3Lq5C75rj+5iJJ6z7CvM5a973W9AMopGqfrS
97+jIcvQmhVD68Rb3SKmkQgKIW+WAHliiLQmB9hr/rnCIkw1HYZ9GIU5izN1fnmn
hIWwRdWnYUIGMPA0mW/AuVik+aasoVKAFZMVGKYIadjmbzVRCDcwmCUNpv/ZvSBg
y+T/s8ryACAA9GPMf3DMreeom2+Ia7ZJrOV65RYVKiMgIyN0MiiljfeUO5R/wI+y
BuT0SiKUKsggrJ5e2omzJrNf8uMDLF5lIIRmeG4kYhEAcqh2uSZsI/0aLE1dr4uT
4xw/uUE98GRyx5M07Hlakr5KTD8AlDCGzfVrwx2O/UOaAVf3H7NJXakhMvQVO5yN
KIMq+R8AfXgn8h+6A0NYZQk14E85Wu9XTFXxIzFqTF1/N9oqqt5l+vHLWpm/9wsi
hLAzCOxNCdcPzlB7pJ4dWuInnXJUXBgCOMqGVShBTu1KkkGURJnVGjM3nxDiHgIM
O+OsmNq/MAPnGH9qXxxcNzkkq5nA/uR5AjIrz9OMVcrGJl+nycIpPuBtywgDocfc
7nB4xWZVzPARQsJxBHsA0rrdVs3PoUTPFlN21hZb0DYktrqqCns6Gdhzo5cJ3b7x
L80QNZ4ReUlfn61zXy1pfkzhjFKDPDNMRQ2lkP3i1vJgh4HZOpU7nATzt2jP1tSo
kopdb4kJFvKzTCMcuF6yAiDbTZ/HclJXkblft/fRQZZVIztIU9uu+UKx8aU0/mRw
ZYkZigFJdFTnc5VAieBsv8eHWI8OrwtfOnKs9Uze0gPyrTrQkE4oHTsLVAIy3yCD
kzyNIuE1QuGS6Yoa9rFBG/5Iia+fpa/taKVgm96o5ozYQ9G9v6OySSflFsYGXCkZ
rRaWfmbG9TFLV8tJE23GCC4idKOIEAQVl7rQgjL2otJ7/844kmwHnj9qjHZU1KbL
owoK4oKPhoLz5K/Rn0tmbH1kOJZgFWqkDXWNzbJIi52KvwpLRnX8qbLDrRLwZ+PJ
CkVNFA0dCZxkIN+UjOJRUJ2a7igOkjSzeroMzmJXNaWr53FcXAJMettfeI2pz/5M
mDj/BYwp8wZoon4AuUs0MCMMJsFD8xHR76LJkvccQZoiF5kSvq+lQnsNAiC/PJ/A
N5zzd6haRd6E0B/1oLlssnGkXwOhKtybPNhe4ttQOxZwS6cDqj/qvhIENKD/Jeem
us6o0YIqvNV1uLqGRibVAuIC394j7jJX7+w+tdmfL82v9Afp5/RFzlE5WaVmLyYg
EBRl6Mg6BoIWxlVV+vW8JhIHWrhMdm2T5HS+XXZQJSoewfH9Cr6GYhFMKz39/reG
lPvnp02Z7NTiVhbtXXMc7JengdOQjvbFIsvkp3nxawKKCWhmTYb6ZEsxrWp2G/lE
s/pBLXbNzt54QYktIBegJXmuOCNh4ke068+OMY/avJtDx41t9DKSOdO+jswMZ1xi
qfh/6swtvUJfJ41hNlU02PG02m822qpVE2PbKygC8jmEqcPB/YvCO63JenGna7sU
X1Pm1DnlpZktQ6g+Bx7cTcHjSPxZNS2YyuG06n82CeywxBbl+jRANn50hNEgUtcf
JXKTNKTkuMYLnvYQbPGk6/niPoZUekf203f5bZLISMGtfcAtiwC2zJ8nHjH2kubQ
Fw+X4eLDiafWvPc5Mwtk+0PyqHJk1IcmFym34sdQ2cHYo+khox/9hm2tDeXDyzTs
n4/xlQdCggyHt0k9tShSqSXPDzyDU2tdWPpcvjcrtjFWibvZlLoTinUTGvxg1423
Z/Cn16l1KhXPBfRxIf+hc6OVTrujKSFn9HHnd2eqK6cYdDzSbdwoHNjiprsZ2dc1
6FzFaTHY1wkLn2b93BkvPx3Bvc+GN8c0jH9gpRHWTOymKkq8hJbzE+meLZWyvuEi
ntsvKkpmKwR/aiiFyRN0VYgJKtMXmhTT4D6KFl9gSMtAXRAohfmViXofV/1dj9K9
5YkodTaNcE/qTXvc05wFqF0PB+0vfHmskxqqUoGmC8PvMsOcgOMdi4M0TdYpO2oU
lMk4RKfN8GU6Pg2zB+L9QFDvDQqVirN1Gau4yx0Xo26TXoA1OAc3BSWH3Lq682ro
/+R9i/cowjwPky9Sh7hefEemz0D3pzdFjmIYlIiXiVe1FqX+o5qQmhDQqOp1Ro0T
cQf4m63JgUfbH1V+l/X9rgFhmZGla2MR+pkFMeAv5bmAJ6KtvP9YMvy8ofchSQQp
bgwSxBnqtaU6ahSlkXYuxtkv8MJszXBV56bohxCjdY5BOVI2tMXQQzZqgao1yKD3
n6AXqZ6yGuVccEz/nPyjZJnB+Ht0b82Pdica/qQYvcZkpTZfHnzdN79Tm47LfW/m
gcEiubGok72zpWamZ1hwlWx1meis+zbKN9QwlReLcTB6LM2dAwLqadjLh5yIDpCx
OK+LWmT3CbCEWexJNfd/GNKnAaQl4RHxdJl3iIOy4mVRLOmJP5t2PDIYdpVNsLpN
o8CFOVzjsWKbnTGJhT3zmEnuQYeehVRzdk86iF7Y95XgXxrq/ovrIJ01VbpMwa2/
52WLyIWtfPaOFHGWmEqRY054y9qQzp6rPhS4dhwJbejJiV0S6FdU38wJ3ShA/hk4
jui6qRLQyCzdVwhHmtjjWZYq7tmeReOSlCJVl0dragNdslmtqLZ/EZe940z/rC5R
8K3QE5gTShAr5hbma2CFbQH5HExqJysh8L3POI//LgZ/OmJEHXuhsRWU4Ch/sXDO
TlR42SrwBembTNVl7Jm/VD23VeX0nR4vTN7hrmy9RkuO0BgYyfE15BJp5HspIwKe
1NqCPctLiGAXHJ8H26Rys0NuodEV0N1Jmmps2OCTCUgsMs1/b/e8cvJxkL8XQs6w
x5A/tYwOVlXVjQR2bLfb2g3QFnrGWzgQl2RgdBTqhRIXRZDU1PzPNnHsv4DocJ3Y
YVDOf2ixCyXhR0LXO2omk04W2uO8LdC1sU463pzFALHo3Bley4XTxKMl5D5uSDOq
1eMk+thj5jv6W9dwUUVI5DrXEJ3QpD3oXMhoxgPl5edX0qx3igSc470DeWzVgYqD
HDIYtk6zeKgzPFqpzxsWruXR4KgDmAM/kLXtwIwjLpGJARbIOCdNJ4KYgsRthed/
JGiGko8+9CoZoG58boP+2UbQlQ0p60TqAiCZSyLTXqMU4ZyqSI82Gs1zItRIMIPw
c3b8amdZ4Y4zGnxnB907xtYZ74F7ZK5XeoMX30aL7bs16EkSiONDBVkFK/0D/PCf
Mnop+935ySBMOStKPVWcegoMr/X7h1+X8fIXpcUsfcaK+Chd5Xbok8MepyyJLvDy
Hso5r8hstLF9JtuwVvUaUlmKfiRE4O9nvVWd3hF9PKszW9utzz9sLkmG6Hx7LzJY
UD5urWes1aLZ3iwMI/Qjh2Ci0XsyTsm1YsnrRsNLU6g4xUyr92ORq5pNLEQSr3Q4
7luIB1TDAcByglRDZD1oTCcsyyAJRSVvD2MsjeQEUKp9WgeoS9DaqE+I2zF3Hg/7
m4C5Gf4F2EXScIM1JRgtIwWw2SL8iIh/iW9e1HJ7WFklvTJT0cgURIWOOmVEP5Ng
II9m5WO6YsG7nNDrTznVLp102KRjOhdRad/JQCOTKlHV+jlIlWNJU1JPXMLTqeyJ
J7ubxgilqYWkCMHixuWEyx1Xx5pKEUvzofNJQyQv04S/rGs24gCjh6+vjQPgUBMz
n2HLed0KEUdFUxIWPH9p4FS2VJUEf6KKakieKFBSx1qgwBttqoVADueTXVE/CTL/
FIR+bCGejxWC55/839bnoin5q6Adc5qq5Fu2D8t+/6xca4kRnFZdLWpfq6tGPIvi
3S7f2sRNEksOkYVBRLxdywLOx61fs8WA7HrTQ1YpGn3e3xKaI5M2jx17IvyhqP18
QjA6kZLUzIxdKQc3jyYHxhDKiNxPKdQkethJBFNSj/e23kojwB99yxPeBzPOKBO7
ev6jRzx6mmMijCMLnVq3Bpn/b9uUIbLT2IG2nKEU2aIKk9+eZucIertBhtval5Xf
PPpDS7pzt6I8ESL51/4a9NafEa7A6NhsHY+rsxS4mYQsp2kLGIx4VAOQS9u9s+CT
tRk/KWiQjCrrIwqftEQ9j9sURmk8Y87CU5zCMZKSg/IqhelusX/alUxP1K7W/IwJ
iwV7fNdWg1D9W4YL//dM59bxL3EmHeLLCfBVXg+8WviZ1lXrWeGEFvyHYpJ7zi5W
e78wZ0MNtRYqD2WVLITX4h74NI+gBkDWDNtHLS8iRvYxqxot/TxHZX5NyFcWvdZy
VSIBo+QVRnSQ6OYx840rllLSxAFgSJgetzJG/8eoNvYdu5X3rCEke/8JJLHAj+SD
9QMMSypEu0JcbPA2Jb5HsXw2jdQsu5o64Ujz1B8sxp7H2/jW3i84PeYF+Sv71Fkr
C5L8HeX6t14waLCLcexTYZi4BtN5mpOC/yyNT5UqpIOLZG+UQjJeo7Qr8n7E7G+S
Lv9v7yUe7c/KmUa4yUXf69Z9QELXt7+gOF8SFDF4GUaaffgcger/2F03iQsj4tyT
RY1NIotrYBgENEluJizFKw8c1qkzaIbNrN8nZEnUNToKNCe/gS+zMx5FkGPMDAW0
jVlXjaZWrYhlar90Jdev1LiHq8jjbJhOGqg5h08jUqQ1wv5pS+TU80xlqvN3uJub
nuzwq0RoBkfRM/r+QNiPZws69SBlBXjLKolFe/y9mTlkZwANBWt4Eo6ZQ7ASyJCu
kt8VGVHl/M3feQBWJv/PG3UeyWkEGvEZ2tRi5DyJAK9ew+yCKYQUDNxysuq2xkfI
1UGR8yhVL3vMuIvr9SqB/8a3Lt26rpBJ2k9zv4IhTjqd7h5wx4x3Qtl2dDNmh86i
m3l4TaFJxzpyRxuGW392X9Xhkg5zJy2G338kT5LbkD9bFlm8sVX1TVvT+TpD/RIg
NbvnZU/VsZN6bGoMH45wIfg6r7c2qOsj/pN0QOnkstg2OQaQaWZiSvPFQbQMnz9D
FJM5/HQytNNGEVlX6R5QPk8nIM96Spm2NE+CkZHF6iYFAlcoXoxPre5XuRjcyiPU
dGvkw77PVB3m8LJbuvx8NqxRMtWuHyXcMPhDOWEiSCJeFY7hhV1vdrxzyj0kU15q
Oe4bsIeNSTiGuGaBFOKJqlwJQSwWcDaiE6xUGcw3CFEY3QAG9kfxMTPV7uRPcjHC
BytD8+NadjRR4HjgukwC4BOhzq8C8Tr4V4e6GbE/ngoAsXQjSAGBDlQEjmmYgDhA
9k+7xlt2G1TFzUHpes/YsBIwO7O6SpWZ8Kx1Xg2BiSR9HoyPtvHjUg2ObouSwlZn
WNtN5BdrHHuZQS99SsW7dhxQki24tcEpkETBdIJkDeKGxdwWMomzq9fC2VJiqCfD
p0/PAO0tT4z+xJA7BsuBCm73U0M1TDvuW0v8Wv//689J2zwBjphqrGRpkYWG3Qfl
SiMoUO8/VTxcGenreBaujGTmrhdEnrgEjA3/ojxkhK0F5AfnNxJfGfbNj/74OovQ
n/Bt3GddAkI+eMvbbPZY0ORnNxLDJLucEtkU74pFRHRmmwtbBvS/yBm4lGBg3fSr
UMZVlz9+m2Ma78w3e1aoG0o/4S9h0x0bhpADV1ZCF8y9j6wUmIgfRkRPkt23nZEY
JN8oSVhlQ1nmW1bGl+h2CVIKwmUPA7HRhuvXhNhLKniVBjpO1OHDEKlnihUKeIbQ
SX4jjIlG6VTqI6B64TFzrWs9IsebqJC4o83fOwaDTDm3SjqS4HszNcD8KbAo6VVT
j0C97crPuGlSk8DyUEPKcotYy62krIzL8MWi5GaORnPdR0Aua8KduIQ+W+nVgsXX
wF3gELZT+obyhzo0v5P5H5BjpETgsn532818VkpjLfjA3e4ujbV+n5os0F47r3Ng
HWQI64nQFiaTQALW1HPMvXSLsW6SdUaoOOOsUyLCZR+zZGrSZ0aajWwTlfGrSo8a
4bqEvPm2uxcJqEEz6UBgieTE8oQBIGpFjfddLjE9PvcHYY3CylBJ2yJRrroyqwyH
RgPvt3Q6sHJCSyoFPzXmn2GA1548Ok0I+Xgdg8Rww7PoAZpZ7jqh66WGo3502JuH
3KOuyMEcj2u/aKIyURb+BDkCDejKN5nTkPLfpddW/+pxATBPeRn48cUz5CLgMZwx
FUZbuuur7+1pqMOuHsCz6xFPNiyohMefkwEcNqTf//upy6+iNlDdg5wRDDg8wo5J
IB0Hnpw+SQtUvmg1WS5cHg1teD5tJ1Q40iyTCRWmZx68bveGVX0ymv2e9GNTBGsE
//Ir29pLii1cWRaMBrJQzh2g9S7jljsR5HV91trsswjEgFkhyV5LRIq27rCb+gQN
NufBqlL1OX6KPmtAOafQ2IyuyF8Bo5xJmADWeXQ/jAHzKL5gU6rGMd+HJehGNyJa
1bJqQuzISUnpR0xQxB7qv4HYWDii+jgCHVU8SKLHW94y9URUdHJkFpTaKYrGaeO9
g3mHHrT+sOzS3ubbU1l1JHglc+Gir2AIBgYpEXkkN/zhAMCmZJ0QZpCaSxSxPb/a
3NEYJ1iB+BMj9Cu46a7dVtVy6NZ4zMD1PS0rZQDdhLA+dAvYdf/BU2/h/KuG84PN
sKTLQ9JeGcly0GFQmB22kQubq+iqm13XrLz2e6FKBaKl2gmiYeQmmyGx6n/TSUHh
xWknF3+3tlrH/L8ZE+QVeUqnB3x2rBEQE7nbUVhZujkCiadHEEpKiS2u74vpxAXF
8/fJBdUtTiaUTfbIR7/MQUHYjPAhNYB2tC6Et6r9Fl9ADSPkMNbv6xBPamXQqhB5
Pgj6Zpj14qJ+/1woSU4cTTSH7a2TYwPtt6F3pAPB2Q09KaiP0E50CMCQdFPXSZFv
2H4RR6Zjvd0tK7oFF/y0NT4peH3zMTvMvoZEXKfGyLgMKvE5WNWL2JJFwikmgKdQ
v9qxrLvKrhe+iMRqVmzC1m5bGg9S4EYmMPHb8EbNddL1IDnC7NLRS9ySYvuOWgp4
7o9pOsXDpDmHJVMPx7lrNkEz+oZ/+pRDiluu8P40XC7oF3qw/QnYjT70uzM+WHSz
7/YyOXswH4C6NSuZv9g4TgbB7FPz28BQ4B6pZPCg2+nfQLh/7wtW5u6ihRTFP3Xw
4YeacGZn6zaK2/xhPmwn7OEEz6bWjMcT9SqaZcZRpsDVvcX0iE2bL04jPO32am2o
gu/vLL7QDdHbKqtzq1eOmy3/Ji2Cvot4MkXmDFlkgixKh2G/Cw+esLrGWLcpkHlb
W/n+kQBaMjqUwNFqAJMI8s7rnR72bI+DjzkfF/yDNExTMo041B7ex1T+oANlOEw/
NLkNXA2BYZkHZGsqS7SycNwg9M/ZTY5fANIUL2y69AhdfOlqcWixKdTWezzJ0HPp
sBn2WfH/IrnL3gMxlFgXu/k56H5/q89NVO4cQ3N7ueyjqbiiaDPldcJqhvbRmi6R
gZiYM/Dn6UYgaFYHDyZIJuxm+h/P3kluhE5P30pf+NuZGwaFgxkFItTZBdNZhLPo
dgFnPh8Ow19skTEneBC3CQ9b2SpYR7uTju58dR7tiC6WVuZ7nvjaxKsCesIaE4BO
p0x3HpM3zjoV5mUSHuYs8n2r3581sBJJRt/N0A391KRYxtPkqek2YUvySv3FJ9WL
vR6fSY/fkE8vQyfa5r+WXiaZtRK3oy4S+EI+LOKdU1kN6uz6a9jjle7fOzmSNXmL
czTGS3ibc5i7AkofFlb5QGGlS3yhkHLeAdc0Xd0BTSgDDjewRJ4sPAuQPeggNjLD
AvbNbu+86z94Qf4qwQULJWjOnTsyhfk8yyXVUZC0CK3JHtHlDQUZFraxaEOZLadl
S3xjMlEeuNT+sFWJunlWTWrdG6AvTX1YM5ztyB2dMET4/e+bXjSiFRPA71qmKAif
d7Auc9XiVWAAxgN7tsblpQu3RgVSCD4OhFJl8gU+lpz3DjSGgZABojfZErmHwidm
Hsa84t/3pF6S8ykg0PJyTl5BUvG2ym8P2Gyh4iUUC3R+A4HZdWvrkAhDh9JWX0Es
0pikYrA+aw56KnS0v+0rv6kgKaUoGWI1Ab7j41FOjRynFfmFH9fCsjWwJ3KDu3/n
CtQhE8ryArLf5X1PhRZdujTVzW57Dx4dQ+ML9HQ7Y3Q8I+R8q9cHcEncsMAi737b
wF809DMkNh6KaS1JPl7Ov3Jfy3KVl2ADfvAF8kvEq/sQ/v3wDS7+SV3RzgP1sRPB
4DPTJ3csmyBLX8BZm/QbrvlAPaw2k750sVt5znJObdpXZZkxZ9Y8+b40+bZjW3sx
YT6RKICjA1qbWnum1WqcC/YUJmFKS0rsBNqt7jjc5/DejbeN7hMWQjzuL0GHsOxZ
03lYbocVUV9uYGZmmxcxrCt+BOnmEfE5kG2zFoVpdHuJBSL9xAXiYdqSqIPIdR0p
XKQpiAH0qCQceXIGbGnyw6FeA+eE7E5JHQtrBuZXMrFu6ol0mpqHss6HeyZiaO0/
2HggEV4FQ7rWnjtECMuE0+xAZ2NL0s3vHXhPmWG8gtW89PiNqY1PINUymwu8tdkh
ZUSY5d+oqd5xAyasdgigIbrsjcXSe6CvpHGwbwTfBGeghWCzvfW04xwzRUa6jyQA
aqEcuwolt/yaaoQ1QL2dE/dul+lU4C+ZzlgqbjP5cuPI+awSWKjJlkkAr5u1ulIv
0llEkTM17ZkO+kkfYKoe+vZwLhIaqCj4y9+O0ekQabq+59rrZUFyH4LrTl6hpPi4
HPRQAha1VV69YaC1eJdRoZt6xkwpVBLHy75SkRnGFynUuwBA6TeUAFVpvAVdSETB
5RVTXIyK5/tCBTQSc3Fobqzx4+plWxuIIKR7vTRVZuobNmmQHRq7eKFUcwoUvq8M
MblQl2VxbmIbn9JkKPql2M3MMfQWBik7dqCsezgre+vje9Grc/72E37Sd/TwBssz
YBjyY9UwdEQb69vFl83SCFULQLwu5Km41MUmPTi7Nq+7010jOV3FYhVOI4HIrPbG
pxYsF+wBMgO0nU8TjvVfrE8HDMLOCyMpK0jsLu/lsFyDqLbj3krYWsryFiYQewOS
/nX+o9U9g145fzaaob8xmV3NwzXMBlUib0ZLjtqJx9V+kQHJT7Dzwo26ZXZH/6vq
9BGXkR+pMpwegjXCT66n4cA6nLrjWAqo5l+Xsg14pyOcIe02Ac1fO9PHYMY7zp/e
oTYk7UtQbZoOeDv92AZPnLM9K7fChbY8WODEhx8X8Dsl3oUJaYY6eP8rx9DYAtBn
k8BOCyOMlAbTiF2wsHLNFa/AwS4Bi9r5sjrcwyKiG210SeeqIrjrt/dTKloHYBDo
drk+SVGlRctBFqlLusX3uSkRgNnRe2M92u2pqvBgPA2dbg47LZWTf8bxKbzhPujo
TJ+ss05r7ni/JuUvjtC9WmFmFWhrpLQFK5Z4PVPiY8o8qlgcbTUjtE0FvYPPZflq
myFTUpqBZZd/58GBiq7gpZg2Yp4nv7+ZkACvQdqfKT6m6mJsS9edNyJqR7GviVH0
cf3TOwSnunc0k5BQ2d2zPUybEavkbcXXxN+WipH0fvg9hwnxw2QjHFDvfUjjE73W
VU5kXERtLtIspi/dPyfbLwY1V7lpfHBWAyfApm5hBWniTLpA4QohcE0EPw8fGS7d
dgAh1GbB+0XIsornwRUcRlH2s3z3qlxkSP8TjKfJnMHvwOzVzuIJcdqEScS9+Lxb
g3XYJOkZ9Qv1gC0TDzLOYLas24QACypAGAzZRUiP/NgO8r/6Mn2a0kFBvqqyqII/
l9qvVNpyd5kOKAaSG4jepkFpQ3wP5vk/aUtQuW1iL3HNW8Ew/6g3Cpn+JQs/zZPb
04w1kWtWA1vXOrtxs59KlDLixoFsm4Gn8hl5/PlKJxu5gZWsu+F5BhATvwcpf75R
5SbnO+2liWlLmC7FdsW76PkiXBoSHEU0C2887+QiZvHhqV2ZN0GXDS+YsgKQ6dGt
Eq7rNC8yg0G8zoVxZWsy6dBILRSOmyiVHelaulVD6lCwlx3OiT59Yqk2PPcK5gJL
QZIi1F8VtMe4KbsIiViZK2qN6orh7hzRtmsSwRA/H0BgkXuXM2+FkgmsZy85yyVh
39ZiR2PfwOX0mIrt66ABPrarZoOBryCdxhle1Mk2Z6DM/ZHmywqjcpn3eAO68niu
jODv6s83wruv8Lju18Rd3fouXJntVBAoECxw8UEgsOvBVKGK58U6hlbH3q3SFHHU
9hcH3KBhI300oT28hxeZaII2x/frAkFOEpE0zHe8sFwvseJA1IMHo6QVZStX3vqX
O235ZzlcflEXGebCIDjhPd2OZn5R39deZwx5gtar/h8/8faEJGJVrZYJZKSqZbvc
Q8u2ffFeASRXShLGH+CZ48+Ja6EbqZYKPkNUfTpXf5K8R89H53LzyJ9dOf0MbNuZ
ARzkfjeCi09wSdGaT/wPr4qtIno5VdABILr5ONHmq1IkWcAuZA49pSKWC3Dy8cJZ
I5RKELlFEngbcOr0ZFCTJoijoRxSsjacEJNkYHbTIN2iqCaCvxcvvhniuYbICdaD
JbZls0ktacYGe9qNiJLGEUX5EsGfe9zQriodf+yGHO12t45N4DK74JOb2Qofvdlo
pg7lcjflLXShYfg43+/ySI6bXbGCPCmym8NpWGk8uS4/yve5awlteTpINyQX4Hff
7FiDjI9mAC3Y1IoNr9fEAg2vOSphxeaAw4mZ4OA2/qylkAICr1ZKBXA4G5nzwhbC
69XwK2OFr++E/wjkNz26tdATkThVR+VFQzHtvRa/eerkkmOgOZcC+Pq7RxA0/7Zn
Ia4y0YstN3EyV8k/CAGCylVIkTJukPU92lFEEt4JZhHUYA+oddTz4rQJuZAvCaNF
06lZPD5FKfxILlaBrQSVj9MfMrPov192M9sgStBWgWjimfXbp0HuC4f/bvvScjH8
+WC2YGII7mnAQp3Swp63db0TSi09arNwa/fDNvlQoKW7bPN2J2cFcpQd/uhufP6l
Fj+u7ho/LusXGKds4vM4QUn4MQBGKMH1QpiWF5zEzlAH+G1jHuNaBlagqnjHFEJl
xpLZ8UcNLFMkf3fRdjjGsIUJH5MKt5RNwXlNztxVH2/csZCJMcEmwT5HrIMffFNy
q7XpTDsyRbLnckiKAFkE/PW2CI+cu9I8c3MGTNOEnUpWSHLLJL9aSGgGP/Goz9d4
epGmhZddnkMbYdqazTdwOO/JCocze68rc67UJJzeKIXQXdLeccg2a4xlP6lxe8Im
s6GJdFB1T/GkGCQhAomSAFvnil8UgvMB16VoicmNJfLEv7lCCQDjWl3JH1/Vztpp
DojPBLzNowwDc0MgfbPQn189Q8BMFBj4DzykQ94tlO9GeV8Xxrb/rLKMaOuAelFH
4jlGOtMbzgxuI/6CyHkXfWFRn31TnRzmP93qLZQh7diB7Ctkpf+fiQ9hVMGd4zKU
jynTn1D6Y/6bu1pHhehX/BY5JbhWhvzQXGaiwOicrA/e0XfcR7zP9hQUq8ytZyfu
nkzX5Iay0oSwAKLIQelhn63tKeSqCWkd//0BCJ6z4M+7UsXPSjn9yavbT79oR8IO
a2RBGBdoNG3j4Z2Ru3FriS0lp7gzMU+vUDPb0pGF+l999bBot8sQl5Y3tTpyHHl1
lN/c91S1l0rPxBKJ+C0k0rNzlOccwVZ15o37eIJc7+2e/J49ujZMULvO+ZS3g8zn
cmBoclwn5evDHP9Pm6nD1BGpc3WTRs7XRXefa7zLC47Rub+4cmiQvBt04bo2z3SB
Ig/hPh1Rhp28xCnqr64voXPQwwhP7Wn487AdfcZCAUxsgSCbtf1qz7w0q8rSY3HE
xLxBZlSW2RIRGb0jXeqK/msKKKLdWSG62l0q1x4xGrudSShSxWIQ6bfOXh1yr5bA
2u+jvlrKMbCInnLJwMSBkciozmHPsWOQDQZ1LASoLyHbmVGhdEQkASkL+eyqzOy9
p0wcJqOpPCQv+VdqBPOxNdvMcgEiYCzPMsDcCMa0TxHTa47B/lruz7RkWwqDSorf
/rciTxf70M7ExjVVKcA7hMMVAU7uucybh8aesRSaTDOsZN2ubnGG8ROW3Nd4gG1R
YPsB3ZskMdc9LKZd04Pb/k7OhDmkmBBEWdMfWO+V9r2RrPex/uiDtWpRJLSyl4yv
ZeeG5a6eI7Cy138Lt6RobMoFL2M01qIvxA+/PqrSGtvT2VtV8rf2UEMQRvDcRGqL
bvBr8yp3GL5QyWn12NTr9PC5kbNiGULDXunl7DxCX/Qdwv3ZpUrIsFYvGs+9/QyK
kQZI6FD5rKw9ZvglBL7nahYX2Vpk9lmR1cAeIVdmOaM1jxCozi213Bp9aAeiUwgy
WcF74ciDQbjQT5hGX6Ae0LK2MFTAtJCAdJ6wHILKp8oZO1cq43nQ0y7LXLxuKOVu
9DIb8WTczSi3ad2CbyfSJL+dRsRNtkpvEyaMtL76PNzeDGhFLsxLZYaCmGBOjSvm
cyFha5Uja5LRXT/EJxcBxJc6O2ENDppfdjCONUDqPXRXbxh1Ij6AiPzn8VcVpqCQ
sMetrSoDXuEUsTbLPASnYbEbZ7UI/B81WXGGnsEs4Uk7xw68NuEN3JhGgoBh343X
Uz2Rry9tUJn9+B5QmU2DVP7plU4kTpDnFoul2MlTbDDv/t6GodovR9RCqC2KEPVi
gPd08xZWhTqiCMioL8DrraiiCzH8GrN3t/xeNECRHDSo/jX1OGx9SzEypOlAZyxW
GzEW/Cv8a3JKzvOVmQHvfSpfABsRJdPJ7PHYrNYc5UtkVRl3OqeIPB+uVnrOqh/h
Db2zAF2fOlYsLLZLRkW4GZUGBsTzCsi7klxqltHRvbDROSZJZp7jX/L2NkLYgrAk
nHC2SwtcgIhQjTTB5tqEi0BK7O3Eh2LYtPiHEs3zU8i23LJbf/68pa0IWkXuEQlh
1D749QGkthu4zfAXgXysUiDmncziCGGX42UNJZLlJIR/ZjICNzqL09IpaT5EZ0u9
9leL2i30ZZlE40h6hK8xcL+q/QKLDh17WHBTgAngouMz4MF0G4LZHDwOXIzXzOGN
Te7WFGjClspL6ihFfKvmSnak7rffFvYf1vXcGAMIOcsxjtjxkm53r877ipxt5B24
55neWMsxIAsjCqRnifC8C8Aa7rNDoEBm5hzdm+S8m9WQwdOjcAI64SsVFg7Ip5H0
piOJv6AtjUQ3cWb3mvt5ZB2/0Gv2fDKdWefdNwkr3suUIeWTUHwVH3+MrcQU3Bv0
P2aucSAai70Q+6OJT/QOTH/5wjC96sjb5fU7XWAE1ZnaTti4qYG5672x6vzakoDY
G9kpm2JBcI6MuKKWODd/WlmOUasdYSab2uz9jffYBTwtBkbfLjdqLkSvYaESloBe
FUaCTj6AcxFoR+iX83ePLLQh4g0+Jy9a4wf+j1jLvpJjqRoEEJg9HfpaOvdWBezm
QcttFObG849x0kHxvHRYapjQhPlASvKqv40L9sULRAg65z3ixilCVI/z2YOi2faw
mIJcxZwLsS3UaLELO5CYN7o095hu92ymw4Yyg507fsjxyHHlst8gYnqf5jmbnqXo
1BF2PcRTZ2BeM83r0BIQFU+iZyBKS2o5+xHtsqwca5fGS2Wihy7Fs1eAegmW/EU/
LMRwYMX7EsxZzV0oP4A4B3Q7cLaMCjA91QU5XFAd7gNMjHLqjajAya5QTxpltlyy
gToygJ4ZjQc2iCq1qWvlvjS1v12KsmLspCKDBvFN5ygSvV+9OJRO8I8ztQXfhWRc
zLHERFT73E2lhM3SfHxpC7MLXZdk/SJYAAIXkSRz9QeexS1nUIp0XFRRbu+h0yK6
AcLeHRUp1FyTvdyf5WM0mTE5U80dLd2jhswN14YA9xWSihvpfi2OC21NoBh3j/6E
MrxnnWaywKyE4Uc1srGgkxZnrvEH4l1xqSl6joAgdOLHt1Eojhcsd5LEoQD148rQ
WwIXg4v1ErvT3OBOpSGS+i8PQ/qlIBDL3dDVhMVwHptX7EHVbWXYsQdiboWViy6S
sgQstIezTqAUYLIH1htRggYf6A+iXGWL7CAqoVPBMuJVSD07CepQ8TexH+2aq+9L
CnuWu+xasD8VUfCc6MxmrTJtDpEUUqd7XAIRXUlESahmxc8zJH1VYXHKRN6c5LrZ
qjARIGi6aqnpF33EHsXabUTzEMtieY/b/3+qo8PNnsg/s5dara8dDz2UQj8kHYNy
AAwAXS3p0Xv6KMlAHVZENWEaRzVzgaHEZLRqvXYazMB0SuzjOGgbn5yjatpn/qse
y+V1CVppByxP5lBI2aPfcVu0ZSdxBPvNEzl8W7qtxG8PaG6dLz4yAr4itJHCg6j6
m2eIvxdOqfDKYMRmXmpkWmI67OGfaYHgOOHHNbXMbmxNN2u/m7o9pPyLDxPeraPB
7vDn9Xo/TkPZvKeijpt/U9OgFr7JrNBVvfY6wxlsHEKE1C0PvOXmTEbU2xLszRSM
6mlhsDATcMhvJiyGz15F+RH5jJRAdbVjgRIjSGKHwrKYGk1Fiz4RZzUx1bE3qvIz
p2ZSsNpiRYwzNgS/u0FhfEiQ+tuOdgAv3c8jsxIdUhGlEgNMH4hwBSxQQHJW31qq
XxMdhtAWGsUFMXXsLZAkgJiUZSbtXh3JD5kESj6zPalru8X1B3/OPtu5n9ZaUQvh
5caRHQRMxG20RQ4UebM57ZMwRDzjv3hHGU6n3VNZN4a/sKNREObR1sBpNWa/m7xs
NSljchDrfxnyPv2wbJrSW1U4FWICKpnBt0QzHfYn5bxbbq0ImAJTVTpvfwFi17Fr
+ao+x7R0sVsulmzSB+dMAEeEAVvMm590AfTf2e2fCBrpN4ULQnc5jsthwXTMEUFe
E5zy9hQtBYI/tEN9cEsCH6G9t/MvA09X/6gxW33kLkgzAOghX/7f/o6GkLVK8mYh
uGuULscJ5/hiDKVn1x0pMQuMLcScZ3bYDZNNboJeA/U8KX98UcxlffxG0hOUKqRi
pxcTMorOHntNu1cq9wYktNr80f+Ti/wLOZ92YeJVv7lkMzJ+xYykroznWAUmeKhG
NganaQbXZDHK/lUVYnJ/ZlTQ/RdFzHZcKzexTPXjLY+tkhqFOzCwGcOv9hsnAo8m
cLgOgZt0Qi2lfsg8BmZr4qni9TOWWVyangqVV+2Sj/p/GS1EBNW7zyCpYsS7YICP
/9VPdxXXFSdBr9gvBc7UKtdSKljGhpQ7dyMfAzJNWxPWfByzGRYUR5kI2jy4G+Pg
dKJ+IqD3L3wkWZaHwKtdntmWuEduDU4jxS5XEKd6kI09lr1xFm/xkp/yHNN062eu
J6RtLG+BUHPaaQeCnMQ5yAUIGHt0UM0r40LhPVydG9dGBnZQXB5eEv8AyIyE6gY4
3o+nTTr5W1S1bOZg3J9ONEjveRVvjbQTIXQjgItJMyh0crxsMM9e4NmjDpwj+SXt
/BdPQm8A3t7BMqYrARtPmphDyp5mwiKm2ZY/tKGBjWL+TUv2oq8d2Y6/IaqZWCzH
OJejJN0dkO0N2cPSC8JYjiwEW/jTUefSkqx+LvjGksFJN7ZIQQqcZDHr9+lzEnGE
RvRHWC8OGy+P5JSqsGbxz9fEKwM++Yb0v9ZAG8FpMF4w4jZEi39Cv6x0ov9FXGh5
5sx5QPhfgOezGd/zpkguY4jIkS+U7osjOeSOxdl2SkwaDhQvNQB+lSHM00fQ/o6m
tLHw4F09xHar1WrQB+IPx7UCewM+N390zEeqJkq4dWzYMbE/oLDzs8sX8s/FIpbQ
WgF2wuENXl9Rxd+Gq6uUYxQ5mDXb3ZWIg7HZXXJrXN2ywAoSaJa3ic26t1k3Po4p
nSwppG5FQ3jb4urBL6DH3DYCb4rPU7nY6LQTguaUs8XgIuNa95PZ5gM1tiCarSs7
rSxN9d6NHBoB8Nmv3tLAZg3a5deD+thKC0vvjHZs84jjaqjrJgZy2wB0eqbMrxI+
4AiDPYGShFuZ4d1IskGARQzmA82Cn1nM1yoS2onIssi7sfAEOD/pdBJzXHr/040v
5rPMEOIlfrdpl+0vhiaBsyuKy8ScfdCTIGOKnscfmO5uma1Xh1fvcfnY/8w100SQ
pBrk9mEbBvmu5YP0CAt1ZAY1JCQrIPYwatHilnmQxJMARBzBCaTeYY/AWTuwYEjZ
orgJApIa2oARoVl3fWtG2+VIGEkvBJDmGXwaOcJB3DwYeIs6uV6wldk9YZHS/arf
/NHu03gDzyizto4EdfJr/opvAxuI1PS+MN7rP0zZvmMNX/P7erZjMSMriFgrPru7
imkzIzT5T81rfCtDJqyNLpUkIcbHm8V07JKpiUP5z0svPmPGwDP5xPIZMIYFZDG0
nu56riazs+Qr6/NzXGq+sTwRASSv2XrT8hs4tvBIeipyUO+4L8Gv2/aX28cKMXz1
JQ7nWCIyiAxYWT9TgLsWr/BIljPu3cUoYj3lDlThxRgvy2vihgwLkfKofwlnHaA3
r+Xz3yIRh2heo87b6Uz2EAyD9je4eCOFI4yYDRMErdwQhvaEd94eVvqXByTiT7qO
VID9JUyhLKyQEi2zFyLTU/CrUwwbKupt5c+XNwI53JYD5jEXETVqKdF7VfF46tK/
zCDbmM2jnYvL0GPNQOpNKtQvnR4Wjxs+xXetf5fe59eAYb7RujAmeqLJq79cj8H6
tqp7p12lU5+xxetdzZBq7jTsRf2QNTHV2Q2UWZBYDxCAujWbSm0R7qeHx9Jh+Dwd
W/VdTOUHEJbkOfvQ8skSb1Ry4hUva8mzjvvQtD7RGLSiqlhn5JkA6w2gToU8cOP8
tQ3PEKcNtjH30HX9+Tj1DKjAi3tXVIiuonuYNZp3GHF4hF/n0ksHIktsMhiF8Lc9
7YH5WO1E/PZ2Qn0PwZI4lG2Bgt1IpBtvxfJafUOx0ZZz86tCPyVXKGE3UKshrUe0
blZHuzNVPjE0pGdXia5mkkub+SDpi8q2OAG16zZPnB6XrFgICQo46G8BTgYmc86J
uGnMbPVY94MYmak2a8D3YOglIEnHhPqiyjWU0NFeDMsbptj4ldGuDm8Md+UqX5a3
0mKpud38T0+vnuqp6Ff/plLOCYYVpce5cpUQ/lt+39M+thlYviYNVEg51yfXRSPt
1EPb/I6W6T3JDAV6IFCh7zloeXBNUQ4Jcx5rwIBVI4SxS6FSWQhKlhYkjrgos66u
dC2rMV63sDTuLwhIhEel5z/2lpK9Ou0NCcXHk5LHnUoSIDAm5GnYTtvneXDp+XCj
u5uaZ/5SUTeTi3kSbes/NRP/OBwvFBe+1hgqDo7aiDajnQ1H5yD5V9O4cOVhXo+w
TSvzS8kv4aCYJjJKrPg9My2aIBhwD25j3Nc9oMz9Ahi5NiXJspipTTEq6CrtUcOO
U6qT4lqLboIQE9PpBYTC2niDuB5qNlXIlIVWey2G68U2xF/fGvDl0AOU1gFukHXO
yYNB2P4ymluPcQhClxQIb+W3TTKz9Bad9+fWCXj01lZ+qTu6ELyogFLko6CsgW7X
tvl8dwCAsa8QlvdhjHeDb6annHpFWZAgJfwNYwaE81/nsgFf+qQnqdkY7oRSjfXU
9EHQaG8ndH/wGLMffKfMGEagy5qMircBZNiOWa1fognp9iL60LZfkyJpdPbqwacr
Q0Nqo29ObY1YQyR5gsWqHh1mTPA8iHiMAHqMa3sA36aNBYQ2AqlDdTjmfmoGlCFC
WsiYDo3aP50AxDrIYvRN9hJK/glR0Le0LqUmUhJb2n7dl0x0APccU2tVXA9MZ7/9
DPXOiwSBPcjtDen5qQdEnedSSNTCfoIMOOpTUwGBxtcDVCaAoJr1o/NmywEcConb
xvXAjyTcvReaOI5cMK6r7OdZL4sYjKcrKAnvAaC/F4hj5HKN7VPeo3spI3F7Twgg
WKEJV2ExbhTZRBf+Nu4NVXEYFwGuS8YVRQ/IUzAD+KV5tqkZR9fW/Iy2jJj+TAQ/
jHl0nsCOdgdJxQfcEf4cQEYHMgoXjZ6x1FfhLIxmWJCkJtIWO2xTkePhKSETRKfN
Lvk2NmskKqr0s4zttz2aPXQvM4PBygtk5WN4zu5ygcQd4sL9dXaQFdJB6QyfvRjF
OYWr2uoEM5DF8ikIjPE1tkpkpjZDOZkRIZtWJTRioAwz4QQGzGDMCFGmjNo+DbZc
Iuv+fvQz6QPBhTbDy7/aG/LPUjX4MjO6sAsQ5jTVP5nB5s9WUBLjgfnQkTKZfceC
KzbJSKaW/HarCgcU3UX80J6D8ZggyWdMhOeOaj7UbVVPXN+cN5xLTAA7g4lWf7xf
NDcG0g2z/IjYx5iBjqn2jNPxfWIB4q28E8SqxVQigi2mYH4QR5cylzBM3iEc5LMu
ky/Y5v4/q+pmqndvA54fhXeKv9Igck7DD4f+TlKiRZtz+h1k06v3+FBsfzIEFcyq
z3+ILv7fxIqYdxUonNh31G4hA0wIWxHFlWsRaGl3SV0aKOUh+SX/FbSKTKYUA7ri
eijS/FlDYRJuKm1H1A2ODgy1tXw2z6if4j10yc+daU4JLugXaQcSdY2nyDFHaygH
CkSgTcikF04OZH5RVS9mKWJ5bWJvF8C6CaUAUmmA/3ZvnrNqfVhKytJnr0UStutN
Ohwad8KY3JISeZNLt8vkA5KZTz5SNJX39YcTObAE0UJ32rc7NwoBd9ymfS9E9R4f
AIvmejOeAZFiUzknF8TT/FScYVj7XubkXasC+NCqmu8Msuc5mM3tYGrOEXLeoJb+
2x+oH8tsgnzkrWJ8CfAcQ5hA/VsJyt/UciE1lGvI/xVhJkc4q6AbB+a3TfwnRGnD
NI/FTLhCWC320tFreskj11oM9vfMrBjxl/c0KG7pNp+xgeNZnjgoUJLN7PWZn4wD
ub6gqX50AmbWWs56mQxWE1dMIOYB2W18TVkAAqLsoQ8Y14+W9OLtd5MVMtPxVly7
Qc09he2+hf9cMN6M4EI7WwOgMNeNjbpX1R9L9HI/KWvPCxJrvdafIGw3UI0vM6hE
+MABJok1WAFxvs2A7sXpEvgi8uq0odcCmVdnL1eWN1Wpwcp4HKFqQy3HF4y0I+we
Of0M52rNvTt+JiKjMxLUyVTIjOUN/uxr6Wk6buqovQpZOvipkyGaF6A1CKu4yBQM
M59iBRCgFWpTpGCBRdG2hsqKMj+BVC+JwT6wCP/F4tAdTPyQDJ0J0tqyjMhu78nC
IKH5f0c0YFDsRoFxvXk94Rd7JjF4Xn05bg6hxH7vRM4Ennpl6a/+/ot8jZ5Bs6HS
75Ko7MWXFfDEd1/AF3URyCVhlZkf7o5A8ybwTfs61Oz8oRc8yChVpNjEMBehDheq
FMg/Y4RTmTEAa8f69w3mqp6sb3yzZjzQmqxlTB3CZ1RjCIzTwf6HRZc0Ic+qVY3O
DtEfGRP8snNLZkRT8FK2x6gwtatt1p0ran0npzRmtC4LSzi6Hn2AkZ/09RRNRjOO
1Jo53lSkxkN3eFEia/yqU+soJMxUnY1EFVuMDTppsRZmND3wgwMwex8b3KnhaU9l
YPXJhOhvjsXbdD7d721h3T3tmrkClf/D/05xYxzAAO5n5DxRDDTrWOhm4XjgzMc8
GsbECrpMd8tgp6ArEjMcKrKw2KCtnUY/G0lma9M71PvrcWQ2c63/cS+MEdhqpmbd
vau5NKP7uKi6pwRK2ENYXTM9ql1AYNkR/l83/RQchHpLANQNgnSopR8+696MHvrt
ad0wWIMzCQKHEluHVuE64TDRCqmBcqI9I6l4CH3j68gB+L/U/FllzKvO8gFQfkiO
4BrNSpNgsWTjGZtH8/zbEqRsQI4oXtS0HmN1gDHjkxZkOlXJGIxbSEoYZDg7togz
XucbOW7pY79q5/qcIWYTGrxfKAc/5vCKAopqXPZvBqSgtUV8ntIdlb3yqTTyr5u0
O7tMf9YwVk1jgddPf05uXObNGsvvfbLBKBdq81oft16m/LP3RRFxwNLQoHEAowgN
9BQBpEYu8PB2fuhvtxDziQ==
`pragma protect end_protected
