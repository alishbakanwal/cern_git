// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:05:34 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
pLFSaTZPgO20env9earoD8wYpIL/P2fgdN46GFk7jKXQdLfejaKLX3MbezxxnrFO
n6j2TfUASDDuH6xcZZDnFcEt9Cj+uOoR4vxtxKsQlu8w9IVwvB40lh8Pxe46FULX
TDudZfmcXRasWAJUQ7H3PqBtT5L+ZJYicAfn4f7aHjo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 17280)
LqbxtkPvMwuUmFeOmMoP5cZpn3o14HU92Ql7I3fMpfOJoTSnZ4bdkwqkelx2IZsc
m9Vl7qC2eG6iaaaQTKweEIW0l9bL+lXm0IHGCbA4xrPekSWueJCHCQYcWasGxOkt
EkMABgVR46tVGaZquRbnnrGwnc2+Ka8HKD1iokUmYXEccPuIqxqC5oR1vtPcRKnc
gUZCcwDiKAntQaZsnr1f0hm5Qm41iTAGn6AqsMDtVTdMibXewSEPw/Vn8fZZKe5f
oxhgASlVNDW6BOt+FEWQoibGqKwXDsdGKa3szZStNJrNnp6tsi5Bk+edAuekbYdQ
BNiyb/NVrM7VxTUiIjXj7q2wk2aCFsojlgrZejXl8WTEn0L8iekjVaQ/aq5t5Y50
Rm9cH0M4+ikiG7880hQlEjcjtOhV+7zWDPQh3a1grNJR5qljtGKTxmjsRky9/vtx
796Yqhhqk8fPXShqS6Psm8cElS1y6rJVm/mKAkne0YEqsnpT/VPmMaf8t2PUgLdv
paxvMTZRluQQN5kmoPahrfDlVQHkifcS280Cut1WBV5X1gyGp+pKCkybcoam+kyk
ZK4Gk97yrSwKhIJ8cXEJCWNWNhPpRjWvkTO0y4Lh5itdsaU1VTIqRg+FCMYo1om0
8YsiZCs40Avu0QU4EwUN0ODS6VQ1uh6wjEpvjpeOG0PbbAmNwcmwFpwAB3o2zHjh
xW5mp/3lkKW+DvMyMSVBk1jbMntjMURQsIMM1gb+L+p1b/cI1RkQLmTjpQQ3Bs9P
xS1haYn4kZbKhN5Y/lVXJyP0p/0WUS3vM/RKPMp/iu6q9cLy6zthrCzYj26DvZno
PaHZVP4zwPzPZkI7td9jdPFrzPM4WYh6aHCma6ISleTJLm/W6hhjsRR/sBQyouFK
I1hAhDsEC7jJsybrUc5DF2GNDBIYT6Arkr0+lQ2kMlkiCbvB2agT15dOqRqM7D8W
0Jpw+I2+UjCyaaCMv819LcdD11oBbx5SM9VNiNs2RYJYJNMK4aYBgEcyJ3XV4tvo
pMI5Kpvfuv5qNapwu8waNda/pduNQmResWl2FAIHLY711jLGmZ/OyxUPRWfwjsjl
qbX52++cg4PDxroJazLFsn4dWZbMrYuEcaQnrTGSAjHb9i6n29JNtz7ROJZymqKC
YGSlGaGmXrgRqWx3dv8Ngd/FYLoXXr7x23AOnGSIno+SGgG31wN1IbRIO5Vs76jZ
7Uvgjb+0EkKV+sYiEq2mN94IJRN22uM8/xrVFror16H0/YL5PLTS58EXZWr5tbk7
TjqPJRNJ8I/w7TJfj+dYV1jPpCLI/A+OL6iUUsRkdv0GdYo4/f6Y9zIWbuGYXPmp
hPARmNPRRkpN4TgCaTkE7tSKQ8UVZgwugnfuA7v8WtstmHC+Tfp78RC+U1faS4jr
P1OkapHRnjJnbZKqUpVO91kqOs30aZwo1GPvSBkc74mBkO1AASH5def6t4i5F0M7
4VRUh8kejHdK5jPu87hDvGXTAo6TRGIk1NKwn8qjY6nSfxEX2bnpi9AAF2Nx51KZ
FMofqrx/XFVrMMGnHFDYaWTPjgWJgocG7cluHTEELwpBWu6P1Wnam0LzAT6Txtdu
cR/hfiRptSiM0NRzYN4C+naCVSQBo7FourIZ1sa2oObJrS6ldXZtJoRX0TUoP10L
u4L7uPV4d7cJZK6e7v/QfyLXQkypMmqdxhQz2ofB+ezY3+a3A/58Ha31YXTCpY8n
i0Y7igeLIvAmFOmnic2mVdojHSwRUeMaMHZUBJVJb80kw+NcuTkSlSNyfMiLwroY
DEYw3h6GlKZTCvubQeLYH96JiO/bejPbTNjQEKTrYYLOk4iwg8g+3DqpyoxiHR08
fUf0IoP2/AKeDmZ+EuRODeVg46ta8Aq9wdu9iXHJvLP4MSmS5HoxrSZVmkT14MDZ
+Zbqjs0GA9lcY0M2QXHDGsJHGZQOVSzR1TGkDTRW+ha01PIVgTn3u3p3jcwDRHnC
IfVmH6eHz+XIbQp8U9VqYaLa9n1GXCF4DUQjU2WtTnjpt1zuEVzpbuY9x2fuVSYA
2TrYCEMUxhvUr2ER4Rsh6g/NohgorqB2is/RSdlARv7ivK5FXAKhkn8ks62XmRxs
/yZ4BEs72HfCS+P8P0YDNLLCD1AG49o8LQkloq0PWBRJTzosOr7POFl9bBgOBWA7
YZePb2+/1/amSWF16PzEeoSan1da2ohgxo1ribcBLgOdtnjjBHypbBCt+NfrkNWN
ONIa+qLailOlefBg7AiFIaLYDUdKLQUdvLsnuddNpYnqE85G2Ek3b5l2+SPmVGmc
wBwsi2FfS4NNFJyJxqJVfwGqqaWPlQBvdzCKa7WTdleGb3wmviLS1kk5sv++FF1j
pgHr1A2DBxEiKNIffDEPw2KPIC/EDjH5NOWCC8vDnGkwEXO53A98Z64xNR3KLJHf
Secfn4SeR3siOH3zS0Bj6KMXPki6gqxW76XJY9IvFK7RNd0bsfMA89pDpq72roea
e+9kwO4riO8/DdBMKxZwCUvE7da+ieosLwyGsKeFtV9ADNpavl+ZhkH4WAyRsHqD
SV+sE0PPbJGuRVGMpx/dD/1cG9BtezogXNEhsTXb3pNG8HHt4guU9e8rv04cVjhj
azkaDckIOaCCxXhvJ7G+4SQA8HLKBbVce4WhXLzZo2yPBk+9DrUm0amdCXs2mGfI
KdFBBBLI8NWpUs9Cv7tRqeL4hkJTG67kQ3jjXrdnU+KuTe884eM7UYtCae091/D/
eDAMEnSU5sj6t6s39oRBLgv/wy+5EOZFzGMNeQuhkVgec21nxk+KLFClybiLZh+Y
g4FKF3nhtVqxgpCNjIzadKMazOol7Ev9MAHJmISICKCm4TUeJ0waXosFr5nzZDBp
0bt2JMyXMYoQOoZ6POBBpWQ31iFQCJV2ejfGeSwIrn7RDGif+POppltEYFly08Mo
BNLO83bONNumf+f+33EhxqTzebezXIrRKBY+pQRMPU7oIow8j5QFbYB4PZqyqpU9
AypHaj95N05UXA/D2km138ZnSVqdJCMTBFk5Ikxb7pnXzzdgH7bAPONz73JmaMKL
Su2Zq8hrE5Y5ez7BEwzEzNlmziO2lG5jMjws2M9ZUOg86OKNpq0IPx1fujf/QNbL
Wt8jYNrzD7vBXFmeI3+B7Tj7glGuhNYx25MXieZxyn0axZxPzruw0eOhsAljX/Uw
meEohT/iU0AvtYwYITMHQ9mkCzQ1w2nb0b2Yh9azJ/7Tu5khvFvPpvhKV5RXPA5I
rYUfgvXu+hUk2VzPWurMGId0+bQxUj51A6/XsBSz0U8tnSp40Ag+a79yewNj5WdF
CkXYHZLTocLeHT8/k0WiXM24MbF4m/QI+DXxnT63wtd/FcpuR8H74prBnWkcUoyk
vCbNQ0LJewe8LKsKLySsCZsOxVjhE1LKC8jIYOs2G1zA581Bk0ZKkmPT6J8+8W9T
0urql39lFonkhKOyFLIsi6kfyK6LiAO9OrHT79h94OdwjjBYzcQh2kB/MrQ8FIPK
Ru/jNa4gFt1eksj6XWUyNZmvUOD8lt0nYP31SLAD/prLgEcOcOIFlhLEAlWIPLMr
WUPBX6yzDX4RIQvVOjm5T+FFE6Zk6C/yEgL8Y5ALSGkSxsknOsWRdoBuLa+hzDEm
Qs/pA/H/fXkh7HyQo/IM2tqrI41PrmoaUq53jt3dizopkZb96IhIOC2WMCHe0RHc
aCtgN+aiS/U+MJln2VhqygygQycgnRDk4WqS3VT5MuH/tWi/igQl0BZI3GnUSsHA
BiPSMRT8vXNa2cWthBqI+pYQ7fdllEO3LOPsNNltR+mo7Igmkubrps2MWx5TW1dh
/KFOVzxGvPzsMMGwLKjYM3P1y2War4WNxZRjUPoaonAVYPA+Jpicyxn0KFYqsWOQ
4E17q349SfIL7waHaXTAigy5incDOTqru+PRy9TtyRQNejWQXmZC3ycE7hSb8NcX
mlsYRgJ0TZC+Jj1zWcIZKjGqiiAVGzbYwttq2GE2EAWRDNwY4C8+6Xw3dGgKZWpf
Ky/s2Vn2kgXHG6N+os5U5V9rud0xpviqd6RjOh1/QU9msF9vZo0jBHnAzkfwXtsY
ZR6JaiQVMNHEjmK0FLlNBLdCzI8z3DtIX/sr8a9NEDDobWanSSHvhzHP3mDitb98
ORh4jX72jZh5HoszyHF3lUbknYmeKvXr4njbYD1uA3cGhX0vVj0vgGl1kVuWIO6A
zINKhNgw0a5THZASt8alcdFSToriLSM8OlBsOfUqOFyNGu4BHoTH93a9LqDhivle
nAAV6osi0fN9Ggeqi7R1GTk+TOS5aybi0JNcj7UCmgW59W9T5WaiigGH0dAPR/Z0
y9LQhatXIyRrfw4x+6S+LpWJwDP8+cts81QW7YHP4wx9Z0rhwcrYX+uodHZptqFO
8luPnYeREk4UfTJCcPbFwhngcrLfv9iNRNfJy6b1p43h/20w+E66cDEJLYPS3xDJ
KEPZO2XhLJUFSmz8a2eg9QA4Dpflbdj/2hss7aqLBo0fJqm+gOHgxT7OOCRaB1ln
P+2D/26cTnTHIdM2ruPX3kq5E0iX+KPh1y5Xm/twHPuX/HpLuva/umapYKKv/AlY
Jw0HP01a1O9+/A8R6RUNiurwpK3pwrz+j4YrS0v3bGCzFrBg60VzWpmiwRFL5y16
Q3sLYD7kZ5ZSaIX6ko0WbZwjOfM0QLdeSAwmhiJpsH5Heh5fjMXfnocac3ImetaT
ZQuoLRvID7O2Xzzq2OvJ1cacm1tXfQgPR5rBC+l1jrzYDMvNpxmvlLP3SPdpWJ4l
Evpic651a/wWdr9N9zZkjssgTeULfkL9Vb2w8W0tMI6exqimHn4URmWTuCPbgdzW
Op+GzGvhthFILvCz3lpOluVzXMPDb5R7ouRb0BuTy/X2qwyYsO0yg6pm8nFK/6cw
iVPUHuq3cpTxG9weA3tlrnS8vzWSrZh83eS59gfHImTp3b5Icm/t1s2TJN9WisYa
YE6QK0rHKx+KN3/zeww6m3FejpYgQ+mHFq8qBwIGgzsK3d2Ylu45ONUWH47/pJP3
HA7nITpJpE2guUBTsCmQ3YqpNeo44ME2ZgZDx65DkHfh0pCEcDk60lM0jyVs92XW
pmUGGBFED9WTXsPAqrtM5Df8vn9Y2ibl7mMGPnMzCGwD7keTvncuyVz5w864xiwV
qJx6JiUmGaDLJ1/pt05V3Gkj5F+U7SQ75/UR76xkWSG1doiUpHJHuANlr9dVan8a
eO3bD4xmq5q3zFHsHrwNs/lLkfmOlhi6uQBRNKzjnIRv/nMO+nqZ5T2QDd3qli47
0VW71o5+zKGz+6FjWhYiDM03SmrNXg8ynFVTl9WprrMawFgj42kNI60DwZEDGxsw
F3t/SulEPbiiNgQ4ufw+DEs6eJHM7p+GZNi1+1EUIRVfAxVPJ3EgGZqfTkuw3QBH
zo+ICqJLhGtkSXhuQRK64xZBBjcB4tsSAu+7mHMqLROYiVZjRC6FFJIXZ5VDbgy3
vjMIr6sCu/5vV7AQRtN3pysDVaLG1uxpurLSpSv9O+9f/YR/ey1Aku2ev54jvwyL
jsoeCO2s9srgGbOPI5i/PgNZ74pZbPJQ3mcBPL8jcDNiCk/Yy4Bvavq6TgSw0Q2A
8taYnhXryPJGCc7YqU8WKr1srlrrpRXwod7vB6ADzq5Fc0wb08S61pXYsTjjpPJD
UqShsS4bjd7yAwloB315EMDtxLoCiJ2prLdd7wXp637wviEcQlCR83/xNxNt2as6
ySkBGxqhv7TgLnMCaJvwQnTATZ8alThinyOTIspQ6oeBe6ZidR03zIdxXfo8Ul9E
hGXgF+1qGWnB1m+VcpaIRC9BSoUAGIc+P4qeeCgivoQGPAlp9bxcDPDohCpTo+Tv
cAxouOJPBhRoD5jvNC/TqU3c7Srx2uq3+nMRbyXSrXKWDhYrRY0DXRP8XPmv0wky
8HSZXH8bngrsAAC/EV10+hQHp2Tt85GP33nDhjAr0FOU/cK0I8wypPFi/nXM6bGK
qKYDnDHVAPfhpcQQRBU4OlXmhSFytGAQnArXT4083JwRJnwa5klRcdq6wswxL3Jy
KAylcBkNOGndxeXWj66BaDg4RRkYZlGoat3B2fpEVsn5Yrci/KVPK2w14VGvXvK1
ZPX8sVqC1YDE9Y+qQWvFjN6P2FgUqrngpgWFcQuZVngWJTgAPXFyVgswLijUVlAE
E0pQvBZCh2XP6H6X6r7MVXMqTWUGw89BSRyK7PEyCrYMtZ8nZ9V/57/+1ypTWFkm
ConmvygLaxG/Pt6b7xPJ9Zk7CFhpLKtfSQeZB6KAgrKD97lW9aD/dMRK24FIeT5l
df3BNPYd+/t/pAHa5of4NCrikhdQZpznflC89pkayj0hCGTqQg1BwR77iHVLUguK
Py5IxPQGLOkOjYB8A5REVYEwWWgQr/ElOhycS6P5qdCUwWrgmGnNOXE3Kz/YVGKo
bjTeozwDCY68FeM4o7m6KMzEV2t05L9aVr7xGMttRCpeVRXIsptezYHC6f5xqnN/
ctnoHaA6G+PyuC+XLhDSgunXe+8e6ZV9B1j075C1h0GA3wtey9ELThyiD/oXFIRM
1u0bZoEWGSjs+4ifoNZSEUvtmVH4GW6c77PjL5fVOoKQjAeVIjTPuPutAN5M55dl
ZT9PrtPIfqLg7UcAsDosulsRUuN1lWMuPG4G+DDZ+smihGDQ4j7KoSPbmYZ0JK0g
VuyqbPvjfdFI3rIiPCwG4mfoEacRLcpDtcy7xLla3rZrvbIRjJ0VD4Q99tnDgkaZ
zQhCRqkm2BBqHin69YQ9QAPZnnOX6ogDfHrrk//ZJ96lDXNk8dzNYoO8JTKT1zJJ
6gi+9zg8+g/HEJNXDw6jhPb8cYBc/CCP+rutTMXgZB5PYBsnxkXwAgBbpZvZw2sS
ufDbB/Nqv7XZhKXo+ZdJKSpEDEFnJ1ulc9v9Px7yxTyXely/CcBD7ByKfvGSzXd3
ucBWNK06Q1titOUZjwxaynHZr5nlIxxotYepKk6ZUtQs+Qu130nmF8iabJPD4wOC
JZ/f1WULlQzVeMu1tnmvjotTEUfGHXpx3FQUMrhgEkh3uvxO/8swWEZ/Vk5rytQL
a5M7UuwQOZsSD1uIB4jSRWd4GPqKiaLqw5x9yo7Ps0BWI/YSsbN86Siyagm4w1Hi
7KaS+nTCAW4ciHbcNjF5h+eyMQrT3ADO71kIM5EfThbbBMTAZ30zz+shXrXx63Pc
FQDiagTnFzZiyO7t6BsS6KaquDi9kOMto1bo7OiQ1xavQAPEYaOAkJeqgc75xKD5
AJ/YMGzKnyiEYyKsdVV2SC62PwSKDADzlmd5weMtBi1AER0CYkkPiMvQgKZESQyW
z2Vddyhei5qbmartySYt7vV3OuWqzNyHRdK1kAqvsaUiAzKLldk1mIecQ36q398v
eebTWMH1UenUZLPDtqNfE2tW0JYvcrPJVvEAM8kjFO7WVZL96oJifXf25XKFEHMM
kewhhfavKZ7iGs7vS4eJ8NZRqQ6wF4ZHTLecIVuNpndAh6tlOyYLgXJbntMuc3PR
c8NB79OojogiobGcI+C9+cGPxQ2TkceU5D4l4XUdNLE7sCj7j1gWKzr+8c/2CKFd
36hAkoO3ciPdRIwfW6ZO5520KsiSdXmgYFKc121S+lw23GAJfgZBfag8Khw8L15K
Z5uigNZtq3FVrBcHRSgOWeow+ldZJ2/KKZHF1Tq0XaLL7c9CE8LL7Nv6h1wXmVoH
GORP82jIznAaf4BnUEnh0NtDXNKdyPCBFCuxW8NJZUv42JX3yHG3y8MH9SkNn38B
z+ON1PfD/U3sJ1iQcMkW1AM9jRRiduZDMbL1+sN1VpPkfdD+cxtNUFst84FVxzBN
S9mx6ucsfr6eOFLT2Nt0Z9iZ9n+pL4+PUXpxoM8LmHpXkeKbHsz0ZaJ1sCuV5Fug
9rh4uMlt7XBM4GdxgDZQF3QHXC6QZIrRabP5Ed22PCN0Ts/++rQTbFE8elzSbbm9
z7nEqXGvVQxZifW0xkYXnEX0zFjoi/408asICYdZQK245/mvjFR2opj4FUlxXztU
b2UcE8fUpnoIdmu66IXCHwcbGUFRDhSTFE6az0BySxt2cepySmI2Gp+KPdbhXvwd
sza2qn10DWPxyT1oa9eblgLX8kGfBjqtE+h6QaEq+hDlyq/34peg01UYMT2TuIlP
MlzuRJQXu3e5MeYc9P9SJGIRDc1q/52oRlMjXN5rgttoe2himcmimZSyTJGErLdU
nQz6PdjJ3b16OOtfLrFoqPwZCU45ct/b6KXiQThpgewN1E+2C/BxMmfYhu9aEvDj
L8fY8Bc0U5DYlQApqM69v/fCg0dN9tTFU0mjyzThOYq8N5H4tmy4GwMyek3HB1Sa
iIlHYnbL5oPub/xfnCuz4TfHrH8umawse+eqxON2xYUJ+VGNzOnxce2GGu5JNgRT
Jn6t1mq6519XXyqpg+PdfEsfzjygOc0Oj93qTHSRY9AopgymGM6SdCAFRSHYZXFJ
4wpO7HXK8B5jWLh71DY8uEgQ019BUegE8KN7cuca61M1rzxBTDH9y7XbQE0u6T6V
vcX/U83/5EWvG3EhZjZJ+KMK2wPJcbvPjxJJZxT45UW2TXK3Bo33wWxxAXyL097+
PfAINR4f1Fcx1yyresE/CwZ6iTvgxBPjEjxzBEqVKixPJTZz8Bc2gjlUuSubowdN
Oo6JOlmpocQiISfPqHrjpFngR91jWvyc0YsQ9PqIA1IAJR5nAzAYi1ROLJa+NREf
P2KBRH1wlh1ZN8U3p+Gy1jXPu5wmovHmLY0y+uSyJkYdkQuzD4F4SUfi489K0amP
TzhrltQ6ijCNOYN2GoED/WIwIp2sSXVD/kwSIO4hZBhPM1OooJ0QQSSHYJ0c/6ZZ
jgHQaD19nTAeU0NvVXFhmINLD4NVD6edZArG2oubE+qpGddxODr6IZfpwHEPBxYP
PvjHR75+2MXJaO/OB2rfb6joMg4ZdBtMYv9z4/gX5MIYdJsHgWSgzXnitYOONHLi
llAgt0IpMHwn0dDlN8wTqFI/G+3a3+N97gWXULNCI5q1cv6Hrev5aySK6FS6Fwjg
1gLhrq24de7nKylBRFgJhWw7GVlaieer+ABSploGx2Awo1qi/VjEi09US+t8SZtI
x1gvAqLCP+i1fDvoC3CNOvR1UruGUOpbAf4KUbHobMYrzUCXXT5sMrOZN+OISUZP
6qIwnYyngjt5Ly7Zf1KzoOnavSy3InTO9VzZ970iwxsg3qjS/vWES5x+QFhoO9/p
qjIliZmu0PJ8ASLKWK2q9Nc/kXPzvCIa8AM1647y8bT6Zp9nLhIj2JzKU6srMkSL
t69MQTTh5+TTmgc1aNKl4GrcR9gWeoTlPbthB05Ml6jPYr6ZHSFZJxrzF+i1rFXq
t8li1QcbsUzEI340dkZxuIfjuxK9AjU6b/jGelA02LrqCRQkFHstZrAxOvW0cHt4
qipsyU/nHT5P1IDdp9jpySi2Yq3pD8FYSCprhNmUPdxtIOjWSdWSJ5QtQsNP1Cts
aRyL91tmNzGdsO0DuDStoeRyRy51SaR1EVy6LuvMA/xZ4gC0enWezQZY6R3Os8qf
EsRgEi0KMroTx4E12XgR/kMlQ/cESu0zzQkpUSIX0C3dHXq2ChASiA9UdbV/QLO6
yql4+VnRZciIFIbPHQsO06ZF47lEuRyOBrUit2gPAXJEMOXfTBbx2q0deImg6MPX
6fNHhiGUHMdtjKL5NtlaCg0STRn3XmwLpRviaaBJX24tWfHcx1nqN3YFSoZRHYsx
MdAEhpoNrHcNSC2yoca8xPKcJRK6aGNcJaK2iI1aDKQVJzCx5vXcXJ0NtVCXZAZa
VUYdAXZZgg8z35nKuPfVBbqhScC3RJ1XerFEnNbJWy8ITFJx/m703FqW+2C3Q6V1
x3HQ/r5222xIHOCheDvhZ1Avcen89tms5B3Opgwp0XT0ViK4cEvqeiwbuuQkrs0M
hp4Kk4PzBG4c8LPZjXZfMG7O+WDzSs6bf6XHLQg0lprSHqKo+Ho6bTGo0ld7LF2j
rC7RF8a6AX+hzSSW8Eg3iEiavQkZUx00MhvsHCbqoCdgj7lKQ4X0KDYcJ0CWx1Qj
dMsva2fyEetxWOJnRavDNtJ/F85vUU1QEAvobZLsvEd1pcOfxLVzRdFcSLK2C5UW
mXJW2LQiocjTQw9EF98WF/TnxsSdDYOu8lVUl6CLbN93WcD9vOaVv9fabhHU3jE4
v7SGFJRiNgWAX7MeTZHW6fDCGfC6/N4QWc+5KDwBdxxoCDwZIVhSlIJ9mFQG53Sb
XYRnDHM+jQy4lQe2CY2JhTl0Ncjv2HRnB+7yaR8Ga8f48QDkBOTRItkzkikjeKgU
QYiGcsi6Hfs9BlqLH0UF6hcolzV99dv9XdeFK5moWsFqQdYKW5ft4husadHAP5ON
N+OqinB3Zja4VkY4t9tS738AF1H+Cqq5aPs6ceyt4GDy5rN1+1CMAMnRO5AwqKJs
BLcNtF5ToVwIiWpCmlsg+u+AGlCXqnYjOhF/xrREl94kdirSbn0oUn/a9l6iJ7bO
dmoQXNVBxrM46M0f8bTUfEdV0r6oY0tJkRyneOiXarGFR+wu4D9hwRoczSZGMNbm
aHPpCXQ4PowJHjJPuyIfs2XCTon7vmfiAbu8i3PZ4aMQ0UQIqDueyK0wA0Tf9biq
haePlrbFlbx30eovRiDZfkiRDtdQesd7iPRRfB6S17jpwj3wmjdD1fM9dLgUlbr2
uTuUcXqvm8F7m9Zc8M7664ExaVBttRaNTxNeA51Yeu75xS55vdWbE5uwmU2yUwu0
LQrqnKhBXYOTo3/Yrwjc1jIgpA64/IwtVQkZI1773rigWUcvZd5OLgDP1yteJrFc
+BhIAVn7Z43tg2w7goo4YuGdbX0u9cReYxSXEAsJ70wlVRbA5eJiN/MgRBZSs7Ov
Qu5+AC12vGGLV1xz2dfwcUQUWHUvXozzTtm4hXzhvQbEVApLddx1zcLI7HRBEIdc
5aE2W/7jhkCQgXLDSw/CHz/vJedz40e/M+0JNQ5sVYbuOvKzh35VyT42XisTjqST
TNHv+SH+ToCYOvE0yBjn5k1LBpb3isUZMlwucXcW8wV7qnoqHd5ArbtWjhuI0wQC
5jC3L60fmSOLXkkqh3HUxGJ7kMXdMpZj7r7gWeDujPbm+munbq2YSVEvUMud9Da8
MzriORHrQqpqo2r9yPbjxNK7Lm4CfozBq38dQ2xSHPn2ZzVxIsLJpdBKdo08N62A
3EhxOgOQRTXaZIrSFla7RfNyZtFuT6udEH1xsF+kD91042WR16E74gDLzbn6uAXk
U33DKA4kNyqiNtZ2LnqsUE6sekr4PYmHBGAmZ9zhlZetZitO8NOMXB+uJKYAwv5/
cVzdkXIen60ODoZsotKpjkeej57kmXPnpmx2cvRf/B57x1QWQL+1ZY1Xn33vdJSQ
WGHW6KTLHRfnwzU0kshBoxkjhoEfZJ67iMQGLxmcgupb+T4hc8jBR3co1ZwduVeF
HQvt8hRtt+3SN9EMnRU0rQVhsNkceau/PnJxg9d5S9TesTWu4b5w6uKEZ0dFRckF
WuRvHFIx1H0xzbGhxLBHHRuelshdkx0Wkge4sG34kvshshuZOqIthnlRVTXOyfcP
qdoFg/97YszjHjThzsA/UKbyyJtmewzGsu3D/rA/wDyJBdkcdRQXP+/U8FDNgxkN
hJqzEgDZDVZwTW042JHUvu8xYiwwAv3phVfDNk7zglAXylu4GfHbNATxu6NdeSsD
ZC5UocgqEiCD296r7on188epn1lKDwrJjaEs1+zhfCWzZPL8OL4V1bVMS2HEs2lb
CveiSqgYAQcLw0BOHyH5EZxYc1Yag9QzpGGN0XXugk8zy49onII9UtgBmf6/OO9K
+7oYNFyBIHj8DVKYgPXQthrbuduISAfS30ThwzfaeVprdIzGVRNkvoryh3C0JWoa
SZHI2/EX4slxPHOy/eqD/2JQ99W6tde+St2msO/e1mpvkniBsBc52blkXgSVgWmj
tCviVUS5JxMAIXJFqIIt8ZbD+Nm70+QB66BI9QwPPiwTpMSwt9RjaGnQQWosNJt2
liZhX3oXM/kME5T6KBPARzL/p1rnh6oCdory0UJVZil2jlG2UhbDTCAUERCSzmIn
yczuI1YdEubmfCkDrHH0WV+2kCTY+rAWOoeGZXyTYhGRFMHAyY576KFDE624MzAV
5eLzDuJzVTKBza7biKeopcbaeVUO5A47cXNGCSOqNF9JlyPIu9SLRWh5EyH3SNzS
fvSnFwWt8h+Tj09PTklfGK+nb7zPgv9tAEnqQfssIRsMJO0sHzKl92ETjvQ7Ev81
1FhfhLx+GV1HmiF4qhlGTmUP1I76obZLFlT1GTvaTlrWKa4+xMlZ0eMdqC65WJbT
oLyy1szHvjlqZ2dazfjlgeOTGBVZKy987ojCYHTWV5vaMeiZgLC1EfkhqbNQ3y+U
b4YqPym0d+PJjnB/pubiKw6pkAjav1PG0N9pjdHwsBMI6PABiS4BMlH554otoh4n
1HcwqKuNfvG6k4h+Nc2O+RrbySkvDnFfz31YE2oaUZtro87KjAOwgxlRyY2XMTaG
OlW77FdYi/N0CfSrdusV63VSsKGhmeNpEFeix0Q97vHFqlX2fODERKY7Ihxk+QRK
xpcFXsMnVopVFWQv6Fmy42FzjPR/bLoZM9JkQ/dmk0jK4HUOHHLf4H+gR4OctoYa
xiFZMc3WsoA8opjSqu/2KvdL9FyaF5Kdwg7GjaVLGcmgyCA5mgQltfQTBi7f9NqO
yfENG9AdzUdjfrUZP3zM0lx9yJSvL2x8aR5MJJhkNolUZmc0UI0qjH/fNPT+G/py
82KN4xZ4AENeTHVAY2JKXSTMZdWHoCcy/qi39Jxi/sYFso6l8rAPMH67IfAFf/2K
sRS4AaGi8CVDa2sXuhPyu26dzz9S9ducShA/tV7OGE+6pYnJmtrKj9BVGkbqN3Nv
91tChh+XI80OUyiLqPwNEtcJl9no5RRduRecngZb0uRom86WDyj5fGtuRH5wwD4J
viOd3HU5WC7++1gCMGo3yTx4xnz8JO0Qot0/wQLYSqhzujGCXR6ss/olMNXnFhZR
zoEfpYyy0aDzII3tDXN0/4d3cxu22wY9nJDhglKFjvU7M7xL2R8z24cHFrEdk9eD
8eJOiO/wTXS7CUDmvUALZiXf8tfzemcUMemuBgBP4zUOwdSHvR0Q418+mlU1LuOT
cjjodnoukElfdFq/qtZZEp5n/IohJSVY+xH3lR+aUXbST5lY2zUSNFh7Bc2V2d2C
mrMFbv6yzrvsiU360AEuyXtGZyAEzVxWN6wH8PTPiiqxI3/F5B07XXDlOo6wEVgS
hPQCJ4m+ofNtozmfrk0FxoeshB2nhlFvX9yZr7Bqefk1FAzmzogPG7FEUmRPaIh8
nmcMBeo5q7hNuzoCbtyH/2sI50LXmdWMfns8yg0LB0UbDEtahIv2rOUFWs0b+xl6
EKjc1YsnvJKxM7TKrTIRIKc/Xy/zXySR0vUSFm6iLwUTOdRJznQ0tK4nGj8EjvNU
YdPjTIcYxO3FXHa5INV2qteQmDoK3bKqWCCW2/wamoqaQvzxD2uW82MZ+r9UpcZN
Xh62PDSdImcV8QDJRr86Wx+qYyUnsAKqXp91CvxDe5SWMWGz3ek1I6ldTENSeZn4
7LQ7s77dJHAMjCqD4H2E5NQa444t17hCvJI7thDFfApqKqAaRY+XCRmBGoRTl8Hc
oJMbw/eTHxZqJIXvU9y6fKSDXvAVjhLytKkR1U+UwwdOFW1cy7cO8mDKoL6VuYqR
l4nxXQdsimVOJZH9AnDtqm4DISi8wV0QCYYZnAefzxxcry2nUxGC7eJ8ZlPgJNxi
RKeQcI33l2OPGSf1v4FDyB4LOEXWCtKly2bPqjMdUZGI+VMIMQpS0SGM2xwS4zHR
+oV/ivZR4IHZyJySSog5Jv8ZAANkyT4Lv/A06ZxZpKWSEzGfY1cwWLlKwfS/OdSP
+Yf+Cc/+IvnrfuscLH3Dyeo6phIWHsbVZm9qlxkBh0uSATt3YibxDWdlJ0Zdb4Ds
vU7tCJwGqeX1n2Hsi9FaCuDHsbc/C019CDhOb1xQSecp56BVtoqMR8RzkyEW3Stx
2GdoFQUohIKvIfWq7H9xXS/pyRqm06v0LkCr1ZGwzkchm9IYRoah1lSC+LN39xR5
pQacbwp77HcdF5DdExBC7g716b5jJNC/LF7VmQGTp0Kq9VLHIy8w8wHqpQC3DTlp
pfVefvfa2X+rJdb3u9Cxgvy7+TAs8cSqOLGTO2iWSM11w/0yUTD7vK71NDOW+eRY
F4jrD5OPCjwlUd4nbSF2y8C2TycDGH25aI1pVAP3a2Y5G+NxNmRfZj1gG2VT1x8g
22jd+zx4qcycYQ5ctbj9RN2A3xRyp6YbrZJxl9bGGBbQ0HQq3JQWSHwS/VY1J7pG
Z5eJxTl8+raIpESqyc8dHgSUV6mNT6NKnbjQK14EHGI7M7pXAsGD0oSASdAYzNHN
uSvBc/G9naaczOk8zvZOxSbL/uLcyW9CQw+h7VD0rQRUYVhEayJzwsveUklnS0lf
UYG7Q0JCRS8cwjGxfLVMpTAoXC+mwIO+IzoGmmswDaXJJ1iyDtoLYU8vquOu/mtf
cs+KnnPHKOy/pJskQMaGqKtkAv8FcrXCMMJnXcqyVIq1WYddnPPKe/Q1MsciOQJ+
QsHkUujhzJTQehmVNpS3C6CjZv+yy/vt3CL61Kgp+902dY1G5fptkebUB/Cq9VnF
pU4FRYEF98VIiHAZFn0R3Y+7CYFDRqMK3aowBZyWlmVFkXyTNCUIC+Cu9NVL05YO
CeMHxiBjxGy/fWTAsRo7uxbLm+UvtUyda2sm2VWdOzJEstCe1UY++qsYU7pjIxWI
1CKntgRR3qev6nU5hMXFHMDp3JR5egRsCwzht2mncX1NLQfvtTNA9J1c992EFRnX
bKqio8TscBFAn7kPCZH5aySS+9G4XBIHPr0hE2ob66ecFXUywXGDQSwwNinxswWL
8bEsbVB8Rl/fr6vn442GDnP25HwlutUvynsphJ2839QH1oh/n/aMlFSf1hCfH3rI
EFubNZJkjY2ff+txwaVfSSwWrJ4Cg4FZLvu8RvtUvAK4DHyrBe94W9+JKkn/sWUC
lMh/wYM/hDdHSfUs2POo3z7VK9Q8Doq/bvHyeiwb5lskNE1ZVXolgKnP46wyPI22
tjspCza8BBuChJI+rHB6kDOg4JRK/kHUK49/jtVWmkHWyOOPffVb4wEhjd/rzoqT
5gyJbFpqlQuXFX1DYtbeOjjgK7xmOjJy2h8qX0bnF5dr1Pul8qPdWPjhQXOjRvXp
EvVUtMpjFaSTjotg09QrnfMzjehd4dNnj9bSIDXjZ3Dxm6ylvL4OA4rS+kuKyGpq
w32txqd+A/aSMzulfg6SKyPmSEeDTNRe8SlViwioexq7HdIMItsubS9m9Jc16TX+
m7/HdPBn88DrfhKzvxHJwHtb4lPGY8e47Ojxw/foxHM3MKZ2rGm/J0FA3Jo5gAYL
IMc913DREuF923JB0jTLvzxHF9Cig8F23rZSpmk+sT+1LqyanV8dRhAM+IV6hUWd
PNTKiviz5YhZ7Vuk/gOpMh4XtJg9GpKTkfRAyIOVix2MZ4S+pcelmFOeL3gzTP2K
Fum80ImvodKKj8S/dB1yQ+US8T5IO7MMsGAj8GO16ZN3oPR3t5+X1tVuufHV50H+
yOvb6bXDmmvcq+o/AfUJhKOU2Q0k661Q0kSVXJxF2JBGjuVpodugu7X+bn3eD1Uw
OIffgBHJNQ/xbFd6MUHNgi49KtaWZ2LWGv4ywLd9G2IQjI6gye6OVPa9iEuC5TqA
u3UCPFnseNVKDACSMktfoTi3vyx5juoEumQ+HPyFLjax+Gmg6UfZX+LIEjL32Eu7
2ysGRHkUf0s+zItMAaLCtyByHvOwhHJfc65vbhtryjhhwZ/QTiE7dRcskZoI6uon
tQ3dzJqJDDdMJ6I3o4bxIO5N5Xt61hGCB7s0J25wLWRyJMPYeCmgcVj0BYlgti6v
tWJgMjoALEOSstSRoozj7CC4MIQjlCL+wL/xI4IrW0ov1RfvXOAIUjlrsL5rJKZE
a6fsMCRQNFgM1eGUWY8KOt+DMmF/jLFkgmNnpdoA9E4XYWgVBCJ7HoRWP+NSshuU
06Yp/UyAkjM9A5qfkHmI+DQgOVCl2u14qB9vz+eGa3YqPSY9xnoCdKEHxc1kkBXT
7IB6UiNx+hdzvqGtl7KuETXQ4HbEKFZ8G3Si8a1navhILk7visU579+uxxWWq3Lt
Bl80KolKtqAdRzEqqzhBd3yiZISyFtf9P2TTNRkY6oZ+PnLsr+RX8lWqFvA9qWQ1
cBFP4jK7EJJGgN2hD4MFpMt9TjWT8Qbw7NYNc8Fh6OAfPSgXV8FPDxF0Im3j15jn
r/7Sj98lSLxw9tdwlsjwb5JmEU15kH5zYJvcPdJXyVeAlSQjGVK0iRQOOzWG2MIn
SX31PvmlSGHoijFpskBAX2CPTHCk7DZOPnqqEo/NmMQ6U1atP6Yu37Vt737crZRg
xw2Wis7BLN5/rnwDUOLhnLXO1wy5rr88dpOr+0NBAFqvesXAmuF22SIgnVoshmtE
IiJybx1YyblyfeuYbJL8R+0hc0a0OnW0cuEl+3IZ8voQPv5sviSsKmG0AaSc3p6v
MaFY4qwh6dvtmYxJbjMhJ2/w2n4Waw4imDqavEOGeqKbEnu2Aw36GN2C+dRpObPX
yFHn/5JFgyQnuoedt9wzExaKsNVnZYIstZbpT11yARxqAkzph8uEnCtF8iEGTDFX
imibtRptH/OPoqkKqmqU3msMxnf1qcWPRJO3VqpqjcJ8cyitAqV1ptRQd5BoYnac
UQjdQ+PMx6aTbbasG8vbrKuXisGazhGM7a+VGI30AeMYpMG9vUTYjThP0F5nmS17
Ak/Nm/36B7sAmXs3EJl4hT1DTjab4sK7wQCBMYbvwqME7tt8+lFgEGCglWYIpuN9
ZtSrdk9Lm9jJby7i6+v1F04yeWiqHUo3n/6nD1MsSwSFc/0QopItnd5ZOELDAvyg
ULdD/iGubG8bCQMsC4EZpc7q+SXAFVQBPni46NTu+j+dapn2FDhT1qPwIYg5u+i6
cx3O2toBHSCLJJfU29FrZIvdY6P5bEXhVzQibyCQtInAmgcAP0pGFyf1Kh7iFnTb
rSAoLDGwalThb+MJUJN/A5HJ2hFQWQEwqHpa0oAWust41aPV41zp6ZB0WgJCOCqA
6UA3RACcRKn14numfKojshefygxusIW2YbzSy9dPAKLeZwGKxEurVonwVjyNZX1k
TIwQPPbBpq+szC3taQJzUXF1skremzqf5cBSeh5/Aqh/vxblM7y6q+DTbvm/I2du
3qO8t/Dip8nQHLdJwWAY771iaAzunZxYZZBoSagCiA0c8W2Z0HQeHrMqb23RIKh5
lUPuS1r1dCJecNEZF7cWlxXKgfNNfyUiGtCDiWkR+hj9stDUREAuAMwHbmrzOy4A
/48q67lpFcmjZKKAg/cooxkjcwYSGWqapu1OL5AxuFpWNuuRl8c6VKwwrLa0x5jP
pRqVRLJyMASgbMnyZByf7PKJBGQwzZ0ViPy9MRiI/FSq7EEQSxKHVyxUc7JxvlZ1
k8ci6aIQez0DuzPoqnwn8/Ad4f2XNP3aKDq8p5c7Ygf7S71e9XXCejcmGcqFREQk
ImKydS3iMp6OLF3giqO27mGA2gisVcXgmnUGKYEEdDVQIfd2ZEJlfL3ynOSHTH6b
sIP5ioF1cE40O+QzlahI3eTn5g65tEcFrcs+CHXpxRznxIe4wdkUmpqVlfaC8vvt
/eDIk4eUq06Ts4BgmY9sJSCGFlR1O0aeG+JLWJoS5ahlgeqrmBaFtXKC/GqgTY0q
1S+IBacfJ3dEd6cKSreTzrrzJIyi508uPxJAgjvoLi9Y8TRCahgVw/SZvs66D+IT
z4Wo+1ViHc4g43O7brYyHwM7t9knAIQ0WgoddrvQyVmng1MpSrti/CNLlNsbmRZF
v0tNfkZJ7mtZKoxSqkDQIH87r4uYPKFV+seA6uVJ9MuprsLfIi69m7gxhQY9hKOb
rOpLxvrdfVFzhEbZLEpM1QNs73cBw/qUq0BUFU7JW1RpMKNWoHKQfyUTFAXXukiy
ZlsvtYHb34C/71PCgfeDw4kR+aRjWRaY9EJKXqtZanQjaYZmfbxtGF2//nMQFZpO
jT0RYf5A5Ad86XrVdCLzP+85huM/Euz5e9yxHcnLy8HN4qQ9P9EC5a51w4A4DDmr
/CvJ19sbDyvczX6Ox9tlahDQhTlXJ1bSUTpl3T4mv+EQAGZuVP6ypqG6UIy4+8vj
2sHHSYxNgik8AmVJH4Rkb5PZf+ijR1dGYquCyr0v7rPKcHn4XseWJ160PzR0B9NH
+w73MGptI0jeyzoW8EI2IrI7O4ylFaOMqVWPs/PmiLRE0C4YU8UdrxAKrNIfGiUf
dMALcCKXSw23/0JFCLeIA0/yGNsA6Zs4Xx3Sb1MLLGouiqEVPiuJEzuZOg2bHUSG
6oUwQfUfv6542ix7oYqnQcQye3KdwkqgQAgw3lJuj8ny9hNMFzdyudR/96e2EEy+
cWqXUqhORTKNKG2WogFSc4MlibHQbPpi5NL0xz4PEj2wGwW7afTfnmAa6iOZ0ObQ
IDTmMWyJGeFFgnPLpGMiaxe6hZhWKMoEURLRjeeK7BxJh1dAvIwSXwI8FP+QHa8X
fsH5+LbSQhoysK1ZzsY73enKcvCTdkgc7MEgJFuKatVHoPc/wfmtM7FLtZ0J1Qpj
2bG2cTVFbWSll68BL+XdA+a7w1rV6TTk/1AzZZzzo+qQKFjZiz5CmWZYADmb+gjl
oMOI/snjmk6BCSh1sWEF2K6k9Q7pmQ9VCEI4CDsvks3Q2Q6Ixr5em2PkUk9w33hk
fpci8tNaLAjub2gc19A4mid6kYgOplNk/Loe5FkLu/yYJs+MTqYRyD3VTPdG0USF
n+TSk+J5X5F3wrqLLPVf0mvy5wE9EMu6cMX5ZW/2e0vFtVTWT/+hwJ4uwuKqt62/
Bcetl6qzLIRidEvm7tPCxY/kxclNEOUpk+x8pR6VJnMQFz/O5vuUwCE+KZl3jA13
FvgvFzdOZSctiWK/iZ1Zf5ZvxAE7ZePlnG3L02P2ixXC+6P9GtS5/YIvmiws1Q8m
KI8panPEsC1U2XLlcD3lS/3CUSYCFcw/1DvO2CiH5Rd+Ics9MXTSueBpeZms3LJm
Lc140QImOwBbIhV7GE3D0EfRd/UbM8ZJGwG2CmTcNmYASAIsSxzG+6oyIF4mcLQ+
Bcco8v5TqWty3J+4P7thwVqFcZBQu7wL6jcUuS9/cXYeRCwXDpLy4EI6QSYmHOuL
ysOH8wLgszQ1ikmOCe6A25rzJ002N+vxxlSM8jtGny8BaBWXsrNqXvhbxVoiBBoU
rZKB2iRcbVLh4ELW6L4x+aU8ur+jcPvqRrsejTKAugaY9LSYG2uvIhoPkU6GysWq
LKpsGuLn3fJmY+f0qxeU/342M4MjCafIBG79HU3/1X9zok3MNQiXKSQSpIXQPWcK
hrdtrU80g/WHGVU6j4o/VS6aHZsA7beOAUv7FAjQozk+bsjv6NIVGsuSW479eaFW
GclWNlxB/OE+18o810yNHnAX4B8r7g2mO/keK5/ObpWtbVfflrwaFlY0Vo/WObQq
XJiQyXijPFJSOB0cH8GH6MiawCGamLRgDDLlYFYbh/w1EpgHT10SvBHbgtq/Q96K
VQehplJhaRGbVHl/8yi4u2pACmqqHFxeAslfDQIhVupuwmUYPLy7+Cdsj7Zz+pG/
nPv2T91WrLFReWxOqZXmKmZfl9cB4rEFX8BkNKEP6pf9Mrfbdd1hDzn+acM6Wfr/
1d7CloNLdBvkCfQFyPefypPmdsdp2YBpPanZzW0PC8hlMfsJPIWX4YkSogC1rJRJ
vfGVXSfKlxFl+O3YXoqK3VcTCJtJORqJ7CEnLwOTkEgmcwM2qnCVBKTwGJ3j87ir
Hpa8zNpKgMDihq89OQt4GQ4zG6MeMGezPt7M2yEWZ6dDF0eSnuW44jCQbNcF5H3N
h0pNSZaasghmLLUcmNXexjGl8b7LsiLwPiKkEc2FtVcjBg5M+2lUDBJKgXRATUag
NDEFUqQfc1H8U8mgwcr6sT3OnF4cPrf4x1MwKRWkND+5/T8+27lpPfFS/ep0m13E
E9qLFI0jWnWOq1q+LGDDXS8R+TpF7LfoTcK1dRC+SvVXDEK/GX9cAeQRuPmE1LQ4
KjAYiuRbFUK0IAUrlU+x08E6YOg5q+hRt7BIXSDbqs1SP7B0xURNFOPM16JWQdw2
WZRQjHis2N5WNpZ0yot8OG59jnYGlNrpjGQLMSwSttsgb2Iz57ClRCYq/n5md8CW
2JHspzOUY2OCLbKM5QtLxCRLLwtoFDsCHraDbf644Oq8JEO71/LsEZOG4QAWOgDR
RBFHxet1vMXrcFo8Sr5sv5vgPVTeBJXqPMzalg/0nZKsFkRZ0nqfrqf2xQvdpfAy
a5ZafUQDi96ADpubDUFRqmW3PyZ2NIrKGzNrsEsJ9k0qqssmhkuuuX0ZDZp9KLDR
/HQspfQVTcUKNXviZiTXMClGXhFmGlpReml1cPhYDOAyn1xR/rb6IgT8gfL+A0ir
YAjUrVLRqwur1rU65J1kzzh52FBmHaZRr0XDRAq3Q9XUAPgw9Ovya/OGIszeUYPN
NsVhoqjAxPV6UsCtuNeGsckplB6RKxuolyhP1Vi7xuKoio2pmd6dZ54X2N3XxnuC
vREYTRGiEgidHPAekYt2kxKx/or5QLVmUhUb96MUKXOKcJ7dsWK7qUatDemEfPcN
VtQOvyiOzzieBlB4yxlkfKB8uvLf/WRKtb2O3ZrfK4f7eD3oynx+SE9X2t8naDgg
+2T0O25rkJxzIEldUyfyUQsaT6IndZTZbfWQ5qk4zLbdJoIeKhEL7CBBChFX9+j+
7XGQZ0gCcDmx4V1iFuFxawWGM4vnTPmRFl2lCXrK/z7exXZT0qis7UxaXgWo4Vjx
dR1le/VJleH4Iyyp+IjuAGU8/+jAirSYY25iSczpE4nCa/KQIM7aT5in14Bicx/B
uk3ztkkmv0uO0ShPiPT+p79AAi415w1GvCmEnbyRGxfGKa/hRPAXJnh+H30tiTUX
6S3LcL5vKV8QQKGtASY2UvVW69POj8WrzVKSzwozuIqAXpckheZhAhK4UO3EeaMg
6Nc0JH8MD3m1awamZc9ZyFt7hXTEJwu8oWT1SvkdMCx5ns1wTFDQqrPIl6PQ2kKB
j31KpXLrRraDdkkkSqS6TSJ4hSjeyad22hLQ7goK5TWxDZ3FONURvPLnTPjtSDPI
mQm9gwJtJPuzSbPr3oAOdOMlo932SmauvQN0a48n4x41N46e87/2uHzBXzii/YoQ
Efjw+yhZhIovp0w8Gdm9H7bGfmxOCOmERp/sQBzuxoTP2l1puNnjVkXbPR1QgqfM
HHxuZDIzRfp45Cvva5aLUMnMej+3M5kVeQYS/gx4ILFc3o4WXo2AFLWHTmXNa1ci
xev2EU3sRRVBW9zyfsx6S3+A3KHA6UG6q1IHK30qohHREJcYDsIAmBP4ZRTqjWzw
yB1f1/LbNM910my/6gjQzXt4C63PRILQcgjQgBlnSGoQk2CD8x7lF+4zLWTP1wS8
xakmgKL9g1aIlX2AsgO+rTs+90x2ZhGlUsExzcvPKzsvJpf5aMHsgYO9O++IaUMT
OKhCz5YyKyUHs24bCD7CmvCmuued6fsqzWgpIggisdynkrSytw2vCj1gpNQ/Mo4O
1iCK1DPa0Elho6Ufs9b/pOdCINT+HQeTSJ9N7s61ddlG2ePoLx0zlJTE6G758Jh5
eNgkwPAY6LvKiPBk/XpQzRLS78LA/V+Zwary6C32O/f5E2vOdJkGp4ctOBoBJEC8
yZwEYpAa/YrE5waqxR9k0hoNZvANQwaZ6SRdLHwUPHdkMjcysaVJbm33Bt98M3+r
eOM1l8DtExmEa0dlcLpMP6lzX/HqqLccw0a3nLjZE1nBwgqGcGS8mub/8X1rJdhs
zpLZgjazbcBZxIwRjFS497gFGrrBb3ZsfZvav8SDvyULUA7I2txnxQLKrp7CLAIe
CEA6jXNJZeEoHok79Djo+SAeDAYLARbefTR7jKbzcMje+/Rd6ovS1Z0g6a370ihw
eckbB09ICeQmmELbyl18I3Z9WijpiTVZ/lKCLnQYqXXayM6MYVojaRuTEQY1nH8x
HNtfL2InygaZjZyS23TYtLeoYzUPLcI0RbcpxUTS7yQYx1bpZ5mf4kohzEvdWURa
Io8mCCYwiDa/vpYOTfalOqn7eFViDiTrvjKV5wOFNFhQOf1VEKI6D5vPW13YWeB5
iDpP/NWsaSeTb31fD1YvKncq8FT7X6BDtkzhKcaRY/zFxp4oRy0T1O8t5jYbT1qc
UPd7lxYDLsUgQeKsgzlRYgv9qAITH6apSgcNp9cx04ecMxaoHd6o92oU53BrCINb
l2UXZIYAg1pFhrmlTYfrkX+YmDq4Eqmtmg3BXhymUXFV5o6gx3ifzSJD7kD8vSZC
4Z85w+juqXhTCmd3OCjvtwZeC4LlE2GUB7HJMaxV7AEUf5zl9iDO2Dq85/MejsDv
Butrac+2pcfqlJkNF3t8GpP/oFU2USvmximLHims5oE+GhRU+Xys0U3iP0oGGZXw
hJhJzKfxe+b2aUsVYfeJ1b65cFTqFMjfXlqNlels1Excg3MnbJ7gT+NQvdVqIKMh
hV1iTRRavhF4BkQ4gEwfa/SjjGOyY3/Ia/LdAa1I3Nj3+t0jbtldP520RCDeagix
hzuvmDyDyQMvpKOmc7ZrtEzEyt39HEtBj52FIqM0WIDhwBGhXlzKUKJzBVESk3Pk
FrFR3TKCmYysmH5evQoeYCK394P6p8IRTVeKGoqrH81uaoF/g+cxm8zwqABZeyMC
/Q+aaegV0n08B18dJGm7vKiYbt34Xyt04cvVSYKkmqnqibNDJAlmijZUUNS7qq5a
`pragma protect end_protected
