// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 14:01:28 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
cV0wl0j0jrBfaGAglnDn4y3vgT4POvZA0DpU1TCCGbnoKPiyjRjqh3+KF0ZkgCXa
1QYOrkZFI87Rn1Gde07S6P/70pcIgpuIGqkok6bAixzCAKC0ECdjDpEvi/fT1NHJ
Xv1zmqSsFj6R3KvtZx3+ifiyom7YOt4zD9sX26Njrrs=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 10976)
S5R6dyXEOkgPe7y+qJlHlSFAFtmYZdEPidOtttkit2kS46YTuEjmy2dQJWoF/Qnd
pgrTsC3jb53RhStlI5Zh9khLAYsnNUopRyhl4X/pbM+c1mQE2/COvX2cNUNQkAec
p9uK0g7UPtDwFB7IbVpa4/ntZ2BJ6F1Dl6ccrqCkybZvnMhF/yBg4Yi7f8rrKCKY
75Ec9+EPLnesm0VebGsw02k/kfrtrad6xzs5KDtAbgKtwYmNTVHUeee9axXcEOOc
+OUY5utwG9a1fisN6mIu3+Y1OI6/qUoaJoQa8M2xYnBFS5qXpXyK1sepwKx5jIgd
A65q3IR1qwiUBMl6gOJ12rEylZq8AfxgPiHj6n2Nd+qAE/HKDu2/eu306n1GdlbS
tSHKG5oSZX/EvEqdfhMNwmenzlpd2/2LZV85TsrdezcXH9jU2TtDTPDKdqMbA8uO
F63i9DxJBSCRiBDBdP1SWfbwmXCImz161NyYMa5nCaAoNbx43KA4sEgcSa/d5aP5
uPC/y+apMvJM7Xf3IjfdufkNzj6imZWwLbOTjf2X+TJAnDM4wxzz7uNJnR1p0vtO
4HaoR4NO1x//w/TXz+ks688F8Pt/5JRedgFmH4Pgljfdgcd1L0AgFNlCZKV6F52D
j1UVA/ik9rlxRR1xGElM92PGYScAKDYjtSwXEwvrG4a07GfBD5lrOEHtKOl4i6lO
xvA1q86PcY2VaPdLeyxjFw+h3COFP2NKNt0VeKXIlt5CJbZLRqToYX6Qjcn6AHcn
xwQNQZZVo72jcHdACQs5LHdHpYcAgppNgzhkCj3UheOYkss887L2rWpdfo7Zh6I2
g13oZkmJ59phiO3FFE9g1twDpAa5ZDpy1tuHzuAfgn8ftC7Vi1YGLohn5x63KnGJ
TfK+1WztFMYkyl29N+nFmB8jwfIuXYr3WRC94gfMTloqfBHwJyqMXZP6qHbFNE/F
PaX2CdnEijBSSG6VkOtsf6shqwpCA41ltbQaGyafQjzNnilr5m7vhEBJtyUCxF1h
37sHl6bJHrQP1AtLyf3OIpe2Pz6W5EuHhDifJEd128pjBfCQLWD12jElIRwkzkVW
LY5sk3AEm1Gfues717aLFQmMEimPfTYlrM4PT0CyGUylHPGcecl9hbrIBmTWKXNV
go8/FywHoWpmdUiaJ16VllfAm9QLHe3JY+/iQ1dAmIldPtTe7G3pz9BLZtAleRiH
X6V/+2w31/FI2ybgTi2ZlKGn+icHC0edErN3Lv9X0+wqUloG5NRGuFQBH3wcbXkL
mHRXfRn8t/F+dhUfCSd5SosO6TCmIrkvFuczz0HGqmlcDPQ4M+Fbb23wqXc/SXoL
y65GNJ9i+ded7LtVQVBsPsozWaxRgLDbHZMXiLGqMTtsUWWPhBH8qDjKeRG5e1e+
tEgpRWzfoWhutqkx2RZ88AQntQuPYpK5z9ktg/LBWwEXYOhq3Lgf2yjx+vRTk2cf
uWfzMucF/TIMoCAwtSA8C8lQ9Kg4kbuiQ2sCI5ngpiyNSNaDJ/AzRBzwBb2j6jvP
B+2SyZ34cg1AeV18vrR0V9sR/w2fWcDSppnbsRXcQm5nGuDzg+RMhvscRoBbDyVJ
FoFzn3cuy3i9zSRCrR6klnNPfP+gAHmT1k28yvP7cGSowvvaoS1BATDjY5crF+Se
6EytU14pOnCYaE40iya21Or9T3Hx7uF9rhPnZ1n0a5WqFflZKGb3ksPZgU0D0XiL
i6qwQh+abjRORMIKUjlvtDsZSHhwj43hirz0j40wgTL3kGfH8eVRnlMr6TpobCkH
xNaP+1t1O88vJtFmjIZGNmuIXFzHEUW7WS8/LqiG1qdkyk9Z0SLDPIHnoMfA52pb
0nWIqDMY460biFndR508wcIHkcDyorpmfVWyQHFEMHFNb80Vc7LPeWUsDGHepc1u
r5B2EF0z9/Mfa0ah3aVXd9u9UUt4JxTd0D/VOy/Ah8nRX+CYklCbVJHhdVnIxIdz
RIksFHXcmnG1fOWQhg9FsjtQlTxrNt5pQyTC4WXv/MAV4RQmEhfh0RB5wKlWJyNS
VxBTRQ3kkFoN/Q/b5Ey85fj8pbJtsnvryZOQbBkyKgKsUmLwljqMTp1a57MkUTNR
iYZd2/u0HeDAMo3EIijRozZoSBq0HepHc8F26cTORap/uMTceo1HGUPoPNFzaIIa
r1p9LgWEXo8UUaXqk1uj1zsioPu4oUmwhWU/ylCiCSMdnJT3VtJWyqgJRob0v6Ij
mPJ01inNVIiwjPAvgizOUdPLEKAJP9HpZ0Bx8iOUlTU27v8gCku4Ur+3jWWF9gAs
j4gT0eXPG4Z2XBMFdBoqr+iR6y0lJLBdNi+yVCXWxqENqPtFnNPbyn74osx2UncI
iWbmTNDGWBezAhvCaOQ/9L8cytk0cgovWumJk7ME1ELLKGIV8oSv90x6O9phj4Af
fVO160pJd6b+fyAYAIqyc0K2wlsVUNZV7w2RYAwbDa/hvkYLH9k8R/wcWRPLj4Ex
GKbtmsgZ4qfP92U8GKOumSb94jT807iTLqcaoylCUz5WmVzwL/0/qeUKzc2oCF3l
0lmttV5elIANvSrPXaWRpeW71QB0uE2n60/u6koJcs6U1ZZse86DHQLctubS29fP
DaQiXHk0Z6lLPbNSZGSs+5SuGkSP/3XABmMesEtORhVH+da/o8+IAa9juFqhu7Ek
e3wIIR1Y9kBgLdnkUOLmjziKwz/C1yR1C3RV30uei3+XbIytomL0kVwj+3ki6C4N
LhY+kBtUKL/39Ifp7IrML72LZK20BjovDpD79r8AjIfCHv0FdW9tfoId/F1fpm/s
26UHF2d438XXNLr75qrt6I8QwU2DElLHNxUnxsKA7sOt4vPBZHyPHMQpX6sYOB48
amDFtpfR16TF8F+fpZ+HP3gqDEkq1Bq9x7MNo0Y9R1IZewaDajz3QhkmYijIb1Gt
dWrO2gIw3KxIHh2VunvKZjaJskX37y+XkIFCa59+fmQCWGDBPJ59F2V5Hz/XWNT0
XIAtt0OGmB7YPcHBpNIku+QszHxqYPe8gPQmLT07cVxhemuz0oJA6z3JtwmnSUFN
qb8UrB4o7BvnwYQOH1TMDL/XT/fmKofdUQf30VVINuylbOLIQDo6Xq0LhQIcAcT0
NBhPuRpL0/4B9qYe+H05iSYfkA3fUHxS6lIp6SwvzaxZ3Yyo7tinJTT00o07Oo2S
9qWmSZZz7ifXuozkhiSt3Lry4VsIFy6b9ExTJsVVxFW+iFKvMQtiKn3iHDby0ntq
ZqEGz+InehYWuBlqlZxMFDUfPZ8vbUY/oIgZ8IlBCZaKixYoB04slUYSQ0LAQi1Y
hsg+z0paCNpxqwm+xtVy5c3+yYJ+K7i9cq+M84BBGHOBjgrwhyAYFVU7PaylJAtL
M0g3Ms+icMaTRC3akZzjuXGXz/LwxOIlNoun4eUhd2w5ejTqFPJwH3kyK1WxFTMf
fx5+n9f3zDneZR0iPe6f9KE84pQp+uoPFlwciQyI4JLLOH1OObn1TP1JqJC7LTS4
I8tPr4p1/pvl9aJBL3FZsHTarxYPqkMbg+Lt8MBKsKzqypReDS35X5lQJjWFedqN
FgXsxc6SpT7KHyUN4Q+Es3KTRcpjBlvwDYY0RSr2vYDMtcDerIrLvjvaqST7RK97
Zrisbc93822+rktIa3k4Ch7yA/R0Vw9bEq1/TfmrgJ2RODb6wv5vsKqhggyCbdf7
ZAmPq0U4UE9V4n8oiaqLPcT+/EuKaeV5NOmB/LX98L/3PaznyJ/pD3OaaG070kmQ
nNATi2p6e1zC0ZViG44dD/esKMUE1naJEo9AoMm9hx4qPivBDsTs7tsztWUeU9Jp
b1VlcRCLzZrjeHCkX2XBCHiSP/VFclrQ7sM0lKZMp/U6jMwvYIYmriMjz6f4DWrx
ZD6pfnOJ49jw1haazpsuQQSICy8juvGaIjamK3sUzbFt3AA67R53bAq4QW+3quEJ
sAKWqbl1iu8gT95/Z5Io62fTdcZsuFgEpa7zneyBZsMM7oa8Xlrs+i8PGooeS6IQ
wyjzYfgzngex+aBK/wOU6JyHfBcbaMMOp2pO3n0G+1k3bQyeDhT+XvUe4lAJ8yeF
EZHLfz/U+ggguIhsQ7GgOiI5u0D2/5oHOOlMZ+w/fgGPAEeKm9TmBxKsQvB3ffJr
5neuEr+TF3x+rds9+mrjFnmtsaia5/0l6UG67ENTfk3aLTdggdnIEAn3GNGm4qPg
vkj0rPja0FmjVnAAO0gwOj6/W+NonVfYjUFF4fXZcCRVwfNQjA2ylmyu9qILw/if
HUrs2Ow5b+TkCFVuYqh/mkwfyRnACmUL9sB56NUQBfEeKLL+BYTqmtVqmyfIyPCr
q3NHdQFDaQtRCpui4IDCqX8anifISaa5CZzasmlpBqkTLvNe3+VXckKjDGjl2Ri/
2KqzZfIbpeKxm3Z7GZbuArK8JHp0JL5BwMVEf5tYF5y9rFtN3JXBzd4mNBa/9qkS
Z2npZPUHs7+9XXfq4CwMTTTF19+puUS1w2UkwKZB54xSx2Z4aOwUa6i79r2HwHz2
sqPZJK8U+ngN3Aj8+HFdOJ5AqL0chmFMi3JgDuLKwzRfYNbkty1tLeHaIVHjlCD+
qog8dmYs5FAj5oe/T99+H7+x5iT0rtOAvtDq4CzXWg7g4eBkA1ZWW7JHx7p14qH3
NtCsOa1tPidLMx4KdXqlglYKVmHy7tIt5PLfv094JSqufGZSapEGNyAT9BM4jOLN
oP0w2Z9aW0RJFBUjT83NY0bpuCmrabVzuwxOPLhHwUvT3jxxEm5SXTRg8L9TlbuR
TPim7iKIDfHgrkC1BwzhpgCWIIdX7204Ye6c3NAQPqv/AOmUrHmj7t+VeKvHlmcx
v7mVOSEkJspYmN98te2ta+war6BFoVMPfHHkOocNC+J21sd6OnRpMHZAeiCZOl29
Ve0JLBZgg4Cta4buq+R7+puguCBNgr/nAFUaMMw1ko0EEXP3Kyqb2CjOjIqGarYj
P9AzGaeybHtO5QeWcwJBJf7sUIyJQCN5bKLbqWnwbdEyXPcpBrBXlbGayr1UwReE
Hkt8C/XX14sjgj1aHvGrQlhaqvgwD4+unVSwoKNnLMJyFflv20Pek500f4HMizEx
15rwR4+BEUoVpzqk92nh0LiSHH5bcOMSVfTw6mOhyvguS5tQknRM6vjXKF7Iz8gr
tlXw92mKV1sQ0uC/G67bxNdsVjtyFKECYTBdVL/0ilb7HzWu5FqVU+JI0KatYtrx
fY+4ip2Nj64J1sKnyQB8l5Vr99QQKNKG31wg6nKbKjnAFxUvwjGIXwRoQyiSP0Wp
OaPhhR59TmsxL+rcMihSN9CsY5N4+FSifaSTkPEiFvqKzHvlQpuKdBhrw7qH5jIF
+Kji2bo0xkaAlEnKfnNTc05I1C9QHgbxwVLDMrBoMGZGDwiHcFDjhCPGcAu3TAIH
dhaECouHPzEowCH7JHIOBsFKeEiBM1rcoAntTXtoR5uCTeW4jCzFvuyhMU1M1+5c
j2c44rUewJMzz2awzd2eFB4J+/OnHHkApABgjuKB8Xs1r4io+14AVb6YFIlcQiGL
UYHS7kaPQCqb6heq4AoKshPzr57rjr9Us9QSGsKBiPgQBbG0m4ltC40tXOtGLRS+
qKaJEZy9I367HTDQFXx7Dlo3dfxCD1MqBTCU0fk/1+5DPzdKbRdKKn1XNLxzuVq/
WSO1rf3a6tjqV31fb6sge2v30eTvUeB+pX4cA6yraRt92F1xBv+4vUI9nbQhFTSh
cEvbyYGy0+HhgCrccIcBI1Dgfd8ZO0vJGG+lBNa/9C5LwL5HdN+/WfvZlYc8FOoF
CRHDRabx/zwJ9f4lP8mPYJS+Tv5WohQpyafTV3r7zrcUX96lQ40piamPGIvQhz2/
7Vc9dT9cQDcsqldK4BD04cbUUrZk7x5g2VceeSfPRVK8XP0+NnhAM93o/MyxduXi
fYUEC2NiD5AXKF6AuqVH1VS2T+oA4j/rtv2BP/QuC3DRALjZDATS34tuc8imzFRY
GYqUH24q8fTnbHnwk4jz0nn5hvNOQBnaL1wR/Tq9LSSoU3XSIg2J3t4PGoYnkXT3
xBgQQ7cIGEx1PpkXietAkwDmrxIj2S1xpLZDuL6olE2KjXiHZYmKVSuXsqUNO8U4
cUPU+GzgyJTLR4piZSkos9sVbJf3a3I77xWHznC4D8121nTlaoHMm6oprHpmRqY8
zBBHG7gwo1tF/0zTLf21aAvJ1MlumOZDyWPiJZ4kuml/qtDB/v7QP8M+pFjRrrxH
9E9C3h80DyTUu+/V+yZsR5ED5tN5CJIi77qSmvTpd3Nmx15WfsquIrFUGhGO6Wz8
vDbMYK7HvSeVpu0VQjDRFoc3AvE8kHgaWXzWvSPlAbZCTW29qH89CzUSvyzi0TWa
zLL/OaDSq5TwxkEaKtu1FlxTNDnEvU/IQKW+ZkCVm71iYqbUg0SK7UlXpu6YHiNb
BX5/uEqP6E0bkJalaeuQG4Z/pkwLmjLeeBGdbWRsCRFqUoEL+rFOP8xfQ5tl69w6
9RxTBs3l7OgLDt1+Bao5uMsNIpPASZSHr+hMPml3Z1OKUJU8G+75UDgLOl6+0/PI
R4C1s2rVpXj+fBy+HDD00Q5aje5zlJd9Fkldv4hECd3p/n7ERmW2kIRsQGH2X1Mq
naeqT6397kUKmIP5aMJJsb+4BpisObIWdaIkltHuuxAY2RqXD76E1i140fgvZxlh
Dmw65tS41lIALthlbacSrvNddpu+abXFiDl/8E78OYh6CiUb0rbB0jdYlZxcsbG5
Bj3rc2NvTL5yJctAzHyMZRxHaHqnVi95oLQ5xfBWR70EdbPF8qjIW8GuYrS449gh
D62IrMP1AZRrcolfWNl7HJfvX8ctcTTIM7nMcHrRhu+xXbSu2SXuDIWK+8ybAUXk
Q4HdbYzWoS2UhZnA0MOizWbVjYxz2PRHjnggPAr7rlUMGdC07CSN1LYormjDSuSo
iRNAbkmIYfP8/TM+K9kz3mN/2B2erj1th7XQ3Cp19eFCY9BmvwnjG3b/KxypPVG+
wWk8bAhnk5UKgMSv7FtkpzG9WdRkQZ8s9TmtQcmkD/xFxFkWwM7oB9x409shlzXa
jPtFgP8VpVx3J3mrvQ3YgD8V3i2OyTt9SmOvihxcDvfg1nqB4VlPc7aiAxGv6w7z
Ip/+xB9bsA4xKNUWcPzPiIJM08Nr2FynYnjNDdN0kye+FyGRVCVu/r1vTmZB2mcx
fRZI/twbL2Y6Ti/nyWpnflxsdWobeCWJ61e83cycK2TV/tmhPYPtHRyhT+LYM96B
PgvAGINHhP2n6WA3aOQRxM6rmjCVuA/2o7HLp6dmqSH2dX2FFy3GMsjtn3Ju9ImP
gdrym1OkaE6FBR27xWzxsXm/zchHa/Gz9vqwKIxyK53TjssbVyRdUbMHuS3sSSKn
izJnO17BY2kJIRHvvcGrzAX24pGIjjh4WT1waRIcDHpLfK1ywDUQ+4l5Vyalsfmp
hnDwmflC2rDuwrlE1vo/+646aKot9/EBLt+MZ+XC6QrVoTl3UFi3uU4LfTlFdvFR
w5m/YiFN/JjnS3xZB1iLKb4hLDGlhwrqfe/39MwvC4WKqanARuzdi+S8j4xqfps1
Jv8TPMa+1NZLwDPVeLPtq6BM4+9XOQFcqY1NN4DqvZnttPLE9lfSDmOZNXuKJ3vN
Rr1eVtuo9rM0s6UKCVN/dceiU2DQi5dPKXRJWFjKr1bofo3c5EW1LUOwUs5scZec
M6dN7NveLJlc7gPSb0S7e5HpaeA3fVX325yfaIkA+5GaH6tQ4JHKIDbCOdxXk/R+
OucyzTDT55c9uPRZ9H+CQBWEtEbDs751c7PFtNOwo3wghDqPrWBtz/Q2TkdW4Cmd
wEAwRxNtIPXj64887m1nSKYFWxeDC/h35V8+dPCZHQxdPp9XJGrkKCHdCWu3Ca9z
ShHMuFJhzzIkk8iUgf5ahNz6pknAOZay5jfJr6ieBzKe0bmPqax4S7PasO3SjPD7
REs+1B0XzRHqglgwfzogXbPG8ydgJRmYy12acO+6wp+KEYOBOr0EgVE6mp8aOGZP
xiZL7JCxMR9a5U4KRri6c2Tby4UJbHg/GA2+v1LkYSFe3PqP3WvJEWzj460N+hdA
MeDUuMRel7ibSuCvcXyvkfO/ByHFH/LKUQ0/jEkEsrXeLDT5Bm3s3hkWvZYjPFHP
R7BeZUL03Nw7/xdrjErGe/7lxt+lLPdtN6SFAcjToAVUK+LGdSvM7QeMtkwsp0Hb
CmC4MW5jxfB4Y1Efu0bjkhnRGkuj1w73290XlPcJSWhhoyeUA+CRJsnU3BoglCuT
Zl/1sPTBP+ScEK3vy+TNdz1Q4WBWeRCbMYag8xjBsILRgxSUUT+94aWD1DAKupZJ
NUGTo0j1mqZfNtDcfCFlyfHi9tJV4iRecktwGObpukD7suc8TDn0cp+C4YcujWX8
ISXuYDnMS89h48gA5kbYzS/Vd89fdtijuQ2W94XlkOn1d3QLaeKpNVns0AS+Pu3s
yQkLU49vuJGzhn4azJb0fLaHLyUGOYRZUDO/hCUn3qnVO9lDx77eER/gkmdEAePt
S83Zc/RENO0gYCcVAEBMIEn4VsiMs/NnPDsgql2+jI9vy6vMiBx+SuNsFy/a6g/y
CYqpkNQVib/k7jYUrSpWxG8DQucuDDbAK6J7a0WV8yCmcZ2mtRvohJ4yZoHT4+vJ
6wBM5E3IvknxfsC0b900M/SzQZ/B8AcZss/oZl2E1mmazprCK+sen39e1X9hMOi2
Eyw4c5mjUL+dJHcfGtZ1nErOiANTIQdpBSpXgOUD3pN3lP0uqk5VoHJB+6Sw8WXG
M4vUK72ygDSrco9Ob5t2b2jbZZ4yq53E5Wi4UOukhYDyMypy62WxTvpgWb/RxkkO
7TR4+SsArWgCyUYD9ievseyvqUWHr6IV99Lml3mDw1y+Cilj0whY6dYaFjg7XFdg
XUKirvb/RCDe1NiJ5FmbHLv6ylevu1fh3fEu5/h3EFLOYIPaicmVNQyIV0rrn5rX
5ORRmOazP6uLUxZaumXwBRFkYSgYncUpO2QkDP5eKgX58BjC1UPIDQKLuBnb6uZK
7aWbEDI53oZJHMje3BCa6SmseGrr1q2QXbjXlQCa75a9h7VTqG5z1NRIpaJXcUvk
KcwPlwkffn8Y+NDniyraN1BEFpl+L5uhQ6cmC7FJNsOK1lRlysayThZ2L30xRC9c
Lmmlc9uYw2P+lIYbo5KajyvMZNlaL2rUu2iPyaKLDiWymBzEekZw0ul7OGGaapCW
CsLyDIrSxpCzP+k8v77KUSYtdPsUJKUbKlG/e+5aC3fseOOhztzdI2X746Htjrtl
Y2hKPUsVn5WmYW+Cq4LHuvXz9jDJXqEdL48ydl3L1KYIaKmuZpNRfU4YBkctCJoW
vpdvw74BRHP9IadCsui59GUKuDQ8yKOnyJ6irrJViEPkZUltfduX8KVqsbpNAtKd
KqNosZ6Fpi4+i/jNSnMvS8j3ps1y/0vNKua0bl9TENZzMA5umJ0otSGU3PqeAOK2
DHW1lsu9eh3kxgwzdpvv20ZyYsGqc3jFWfx4hHiJZT9MvRGer21EAUzLr6wlMMIo
nBWRsfYTU/dUuXynhP29ZPP6fXePPKoo5ZYauks9YWzmqr6eEEjZLSlZqsQdErcJ
IMuJg4K7Mk9tAXSbvWCpbbyFrAlzuKWcb7ikG12pzc2BSTEcO8O8dDAoPrJQx/ha
IKd0IJWLPDVxj+U1W1v5DxbTqaGsFUsezMj9o8WYuJyF1BuuGhYACRqrShUeNxRj
AxtYU6oOhrAm7iNdp/2y31nGHwWHPKcPP0vVmuv1A410fga0RqgxwT7Cj1AmVC/c
yxvCxic/G5RbJaTflmLQ9N1bLwMzilj+1Jm4RzAng4lKXM6tkFOzLA9UowZamGJt
oiwDLfXlK/1FuSqgawaKeydTlI+zp9QxOF8unJTqDJmuVPVnAUinMYhy8VMGMqAA
Tj8oNSzLcUO8yyk6KEsOlt1aJZo4pnvHyH93fAsdqZxKFT3o2EKee8HTXZ7IkI6C
mLwIwg6L07ruEtO8HawYf3AaBH4dCWk6+4uCEzcVNKZMYaN/7TUBXxSHQTr6x2BA
w6HyN889smp/STAlQ3G6LNUHFRlqcSNufLWAY3vY/Ptn4frUEp3RUspaOBUvCv8M
Cl0WfAvwJo7LlqAbpSbXDhIxvpT88XVwrH21I0/TzeP61ouQPV3zNXbd+p+eWEYB
BWNC/mEWpQaId7o7/590kdqMQc6iBSVxZuwhg6HYQbXADxbAUcjeGvRFu7E7fgG5
Tg37PhyYhU0/nt8y+tdN8Kd/6dfgzrWhhpFXY+oUyTF9AfnHs4bH4cO3ZnSkahwq
Bk+2cnEIGtFfm8/GpdUN5SMfMUepzLfE2ezhbLZP64h8e64YvHOijjUeZ2s4Is/H
97tcuVEueb3lnehSo9U+lIV3+W9zllEk1Kn+nz6+p9LGZRz9k1U+dKPWKf9sBjHz
RSSFe6G9qkiedQMaaUh0tfn2HZWh3OY1v1dSFfudMVcjz+c1th4S8BzKTgNJIQ1n
MAuZpGXZs7eUZMPQKSB/iYaxuI/8U5QiXagVhwm36jJxOCSWN0WW6OBC0bApWeI+
X6kBK7ijpNgfDig5zHkwEawxPM1uIo+SjKZPyRGvpmduteY+E7WJ9/L3z0S4sHqU
kuiD7jxSqTovSbWi0tKbnDPzq+rLhu4G7sxmjKnYPVW8DGEPK9aa4P7CwhmcWgUc
glmNUrne91GyNzjzM7wOC7OmzZr26V6ZX9PjUnC0YeToiP2w0A10b59LVvIIFQ66
WC/6jlweI7IXKAM3bTb+MnViyZZtzL7CuCghXXqXDXJTNt+KAcfynQfdD6UqpswS
Br4L4w8S5Jxe60O9jbhYu4nVslcPleTkjj/d08SvLwAW8ygrDKK1aUEP/BKJcBL9
8GVF6LonQ5YK/tSKvJDUP1zPN1bD7EGoYLWaug/1ADrr3ArD8zVoLcTz0SLP3NcJ
WgV50Ih++DmiUWEaUr2V3e/+/8jfDznl2ui0OLAYPGpFgElfCareH2U/jdR52Ytl
xGyqdBsr9epmoRczVsCI40a9YTeYIb6CFDQeOL5APn5xIP2fS3cauAZ4xKif2JNN
r4Yiz//PClJl+GkyWNvW12wNouXrfzdVFxfX3ZRTjXe8VaOOY1h+OpieV6NRiERk
LE/Vrr9YJvD/e2/RRqsi9aOlgjsHULxVl1su7X/E+TAKreVM/v30Mo6VwhC/Ea8e
588sg59gdUL3NqbIhESfSnjD9BdD4fGP0mEg+SHh2SS7jfO2q8ks115HBUMIJW7X
MZBMkXl2yFB7Z18Z/Tlwg5L0a4WNji3woxwfcCJ8p26WVUz9H8XtDQGe02fbZhgt
yipmRBLj1S4okB1iut+fIyf7lmzMhtPJs0L0twia6U1ygjYNyfj0tLqFc0k4CCe5
3oGCxeWN6nFGm8tQJFWmtrIKXIylQriKFMSdPqRYdDwo2+3a9gWMmJSvfOZRlX1Y
I+hNF43Up5STfpu2k9jGHqZguyP9h93jMEJCdi5gWMN25iWBNtiAu+H9u9/sOwyZ
uYXmgDb8V6mJnpi1g6MNi6Erdn7+dEajo/8a9FCy2gHRB1GTUU4B5KPTNWzpX02+
m59WM6sMOJjcbS2Yy2oJHsao1BFbRJDyHX67uPUYO5a6p0LeV4y8CcDxJLQ2lm0V
wvqQK84nfJM6Rb+KHAQPdu1Ds4u9g+F7Spnj4PZq4byb+S6IlnASuwVJzJWmiGqY
7XMZknIPGNyyAz//L6n7C4IsiHqdnovY0bnV3J0WfT57qBCMpAd+InpdyAdG8Ard
VUnWfqejr2Ak93hW4g0czqVN3RGh/mi5dxskEIUpE2fATcdBXvZdb9GWxCNu3A1p
/ytD3gtK6hNaIaiBqODWIZLDUBAZl9Ix7heQQhjHgjIpirk9vEcmh9CdnHtbjvga
wr3/f+moxk5aZiai8gbXEvF4e7KCWaceqdeESzuEDPP3VbFWPEgdWmYwRvQF83BM
3/cT/Ji9BwBjfflDAL0oeMI43DMNcQP6+m0+CelI8ITY8St7XjUY1uruCeLIlZnF
k+NQGx+gb4tQ1u/zEiEqJlJQuRDSaD57+I6T5lz3d+YoU0oTW9UZxpScsPL2gpCo
XQCjhnn8FvUewTYhVIOhgCCUy0Y6RKuB7Hal+EjTF3swreONiLKx6F4tbYjE+yD4
AdQDempIpGl2pFymKmpPaEA83hSVo/yyP/41iTInp2OPvuKnE6LIfQrf/m1AaNfs
WV2JFnxgUmaqMozboCJiToVO6IdX1e2r13SSbgL4lDo0LHZeQpRcRujjrqfGmEQY
owXQdm3jlCq+1g2vMwZYu/yYNLuo06Zjlm/Wldt0qdFylBqWZZK8y+TLgWgzf2bH
+n3+1xf4Nf21sndLqlqX2XLSU4W7LcZ6GQ1OdVBFe/hC5kEEtFZK6S8dONNDuMVx
Lhf+fxPhdHaTIUpPgT6FmaKlwH33sqA/QuE6orKFt6lHzaUq/GPnXCAVjMFCBi3b
NCpEmzfDtobTZVd0hz8w+0R+CkRHhGWqXslTGp4sSU2XPopWUDPEIVviIVafMkvo
VTvJ9Z5x9cR1SuxlsFbv9VPEt5li8/jdDDJgPqleilXypPFVlwx1EC4UxAq8CPqQ
dWyaubg2DS078LHfxMxrxizJbsG/8zC7erjBSlqjIeNi3zVkS6S7hvls5zhVZ2vj
qUNpZ8PrZOiLaran028vUPZHQf8MFPHCIlDQOxCdob3Ytha0RMvHpmKwymhsqFfe
JDUz9w1niRBsRl+dKVBjkxCmOocYk6iMxXKeTuhEP/7JiGcMOlhc06UxTBYdthPV
phb9reUEKXT7REx7hoecZR9HQcR/ENDZcDywzHLmfBJBApOrn2qSqcazKiHHbOyH
q0uWvQhXxO2/q5a1y4R24h5ho5CmOOug8+/JajU6hRLmMr2BHMsHRzcwD9tETKvl
kUNWrAH/5ArYFB0FMRFLCV8C3HJO3JcT6QsngU0S5U62JYHz3dsW8JMoPhFjLIz1
usEHe5WjNeRfpOCGZb1HGOfhsj/aV50z8HrMpcYhDwE1hPovAuwZGZGmQ0/OvCD5
ddD/w8us6dyATG5dFR4s4RcvJ5YKHElFZgU9mfCIt7rWqVpM6zNvWetpMb/rxf5N
aTKmczJrrQc4f845Ku3RJYUHIuvHbZ/pRDg3+t4RsyIBfcidpFbmCQKWR6epYjnt
wshkiTNl1lxLEQsJy83U5wx5h6VaOIkvKykcdHwu4CFGBoZlLfc6IkaF4xT8JPTQ
2WpwSmvhCW1Clp1WPJLwmmQohP11SblVaimRL4RU21FcHxrz2j4m1+HHKDmi3rjE
ztCMRpd+dtJdROwka7PCr2MAHum593n1dXWJhHr/zHvJ2l/1HdzbXCWrtopKLiTa
qNPHHsCmGifsVY8q1yIXci5e+f+BY+ve91m89y+WTUh8NaBBG5t9j9g2+MJBqSxC
tr79ujWjp4DIQ2qelxjdWCDGxM588odNYDDLoW25/UrJmp5r31I/amjwm1zGoqK3
FB6j4z1qNgQ/pjwgoykjyD0fSZk8AwGBuqPjzu1YqS4T56DcyO8F+5njEGNNOE3F
YuRKbmbW8J6G8r8WRULPROCHozwheyb24lwkVI7XfZlh+KN4HItRly3NvH8Yxr+6
gyWY326E8+zcWu3hPlE8V42dip78FbM4lp+Dx4xs4bfh0i3cxKT8aM7PdrR6Holu
5Cn088CS4IdHyGQmlKKNIsqInUReu5Cvy+ICSfTdwkokMUm0P3kPvcLSoH79+M08
/+HS8sax5/aqGpXJw3vKhpiW/Dg4cHBPz5hRU/3BGZnuBrLKShNFm4MVLTZ4f07G
UQDoGgxZCBS6Y1PJF11R9Pr033Oa1v5fbamSXXw4QgdGxHY7Qe9D/EOoWVMl/niQ
8A0eRfHG6uf3F3yeFKCl5/QrpvPf4J2eOiJoU1IVDIl/kA+4XIBkynrTBy5r3smE
EW0sibVCvLD1qoQdiUv3u6l6e5quFNhAfFSY1d8SFECWkRtXkOxI8z+oeKM0M1SE
GXX3QTy8Plj61Kcu/XedugULbgZZgH0QvOweQLE/q7TEGPWYrKsWwmenDDxOweTN
HRZJg3HnHN1OQcxN4PL2poYN5+2CkV4Fgi976N1AiVSbWDGgg/awk018gXI8KR39
T9dpQq+r+dw/eWKKNrZdc8fEk5U6Vftvj10Lia8pFuuVmq+m531ddR2T2IZR2vBu
oQmc1rI1rxcjtyud3U+7G6hqgnN4hz2oNPkQIsR8rx6CQpiDr6r7PXzg9NYuc7R8
tLav+WGD0iG5zrkAR0gd3UmtHztKeZiwN+ak4AWqH8HzO4QyPhALkkYwvySNYajK
8qtVSnLNnPhiULyIPEa3o2Re9HeAYmjB0ytGjQ9E/SJourHNZNZ2biJ4V2sZsjie
8TpacssWEup498p45cuvYukuOejQWp39hs5QhaYea3DTJSvxRtLKfpv0yBkqaArO
mu9JuXbrJ2mHT+caLPaeXLxK5PfrpYYC5+5Obwew7OIJZWqL/wUe2YVSLmD6KUUz
WbSn/J8P3o5tJqMnCxzME8dJCFKUpH/LUHqfioxn884=
`pragma protect end_protected
